`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
sS6PDlWNj3aRpfheCtq9XuSk2h5AnQWKgRE3rSmBMs2lRuxjgo/7pddzlmIzOeKw
LaFdkzc+dUc6qHwqDdM9cXXGLAPeJWqnUbholDA4cfqCsVnFybzWYILFEn5anJ+h
lNsLwtFYrKboHgBNcr3cKaVb9jsvDPSeC6YH9VrZBkc=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 59872), data_block
sStt1XBEjXIc4MfOyCyitFQyrobQ8Uv58/lNPaj7IY+cbbjiQG6qrZ0yhE+/ljdI
8fM9X7buwsHYJffXg8qVTCshmZHbDX4jElD9hr/dcxTEHs2+hskGrno0DRFioqat
UOnrN0ApI0lSosTwgho3mZ0LyF7RUsEBPVMLbd+OcCJEOURAeWAPpzs4WuBBmEog
r1xCZLppfFeL+6vOMg/HvQ3zJO5ZF3BtrJRfrRzTTV/Jp+K2cwjbSA+QeS0fhIr9
5OutIn7EbTvbWOyLl8b/wuZMy4WJ3k33aUdgQPUgO0rEYbW9hkv8aQsq4SLHOPW/
nK1wYZzBzhXY3CWnJPVeh+Us/1WRUz7nvyiP4J/MpvH7D0wCIFtP470TMNHxdGW9
zzmjwV12V6HYUEJ6pw9vKJ39Xr4lb9+Q/Dvs39YkY1TPPh8kNENyIpxkIq3yLqm4
fX8i6iybLudtKHmiofc2iJQ4n/MkL1Ikt6yklNvHO+pjTVL4EJQ3soqxq5dXYlzX
k7d2TiFH4HxfphMJyC4KkLzZxMvO4/9oyD234hPEwOJdfRwS9AS+NlDgMzs6GW46
xo5N+7njBwYJT7HZEBmANLAvJj6/nja+gikx7yJeu46VPfqtAGxPPkEL/8TyV13V
QXFkAULs8nMqLKB9kAKrQlAsfkJbaFDLht93VoDbSTI8d2io+YLDe1pPzF8OG64M
Topoe25z7rMITlRAGP+VWcWfqTZ7u0WWs84qk7zYmPlXYPTwGlgUQprjPjx3ZjeT
xZlYRX/ximmE5awQL8s/s6NSAu5hYUXyEdAjXd7NQVYOF6LRXctcmRcjGtCwHKae
5trHp7CBtJE6NuqCCcWUvmkIIkoWMXgwUaVjC2a+7YOtBFtXmRGykfUiK9XgRAtl
t8Og47BkG3rgECBA+I2gXaEsdIEcR1QlE7jJUCmxf+oHEn3coz2AOVFk4iuSnSFh
edfFRBvQlIQ8mifkwK+zt00snfjN3/8BTjiOVh4WZoCOX1D2FjMjzJVtz2bVGKvG
BCx0YCt7ex5gPy4Sm4niq2rMsTJGl3zr+NH9IPjDeMhLHgs7b/3lj6J1isDUCUXe
sHHY7DXxs5juNwABGkUyXS0ADbfVsdAXKRwrwQ5sehYLEKCyQ8FPSs5xLwy3ChM9
aRpL0HwzVtNn3Gvu/JRD4Tc8NV2DkhZxIaBc/SZiLyWFdleeMHIpKwHF8lJEYWZp
nV4RxJj0h2mUtsrMHnCKX3DwjAx4Yv5hsDuhUNG0FIl3CUjwGT52SOo4Fcshyutf
FvSRy2t3gAnoBmM0hxNEXkLMxeagwQCuSzKCpBGy+CjkSyJhCFYrd+wdSuhIlVne
QHngk6Et/L/sVxaUrc4Mk43PsR0bJ7b0Erc0P7bRXVI8CNcrl0TY5DDGKSaVaQcw
vp+QHmLyk17r7j9x/QXWew/mbNZpK5KsaH/i9Pzpl1PyDjurfc3lgnUSdJTYbAi3
5ClrCC9tKV8zheFUoTaMtSGLj0b6W9hxQpcTeyMHUlIUpEtiIuS1Sl4W3nZj+e3I
boIIaMyowDOa/dTIIONBpjU9b/PmqF+xR6r+66GH64fsc5XSWo0NXqOxchebRqhR
5T2KWzHXGYcLUh5UGnaihCSq97bDTab7B8S8kd/YerPAFzmNDzivsAFAXkQ7X9hJ
kg/mWHk1V0IGNV8syN5KX/LkX9yr/pziILcgEqcEmPytXGiV3GE6P3//LdR3MYkA
6BfewvLweegOgR6XJfPGnoapyJKtfgkxJxk1MTNL+1RJaY0d4XYPr0T5Zren+FPU
VQ0XHLOCFkcAz6IZryEelHP0YJCf/oLfsGdizaYHJGBynhF3QA7ZP/v6VECua8tM
x+jHL/9TEGTyHFQdpGj6XqI3OPnio7Gnq4fukduk6aGN8M1/gL36afX0noGkjy+V
WG1vT5ryE8tIIfEEji31M26Fc+BKLt4yp3yQYGK55LN6d5mV6KZFiyDbgTkCNMBm
3rGgY0cOViA65AV7L7tnHPj9k1FfYvWTWad1UZW0FKG2XQ4vZCiNJrh22/fttUJy
+Qufd65uoBL0FLryqs58ux3hwZXb03TbkL1s6h21Nxuu3uBYZZb4sLMDCbpZR8mr
lVJc9lCjOsfcnqS/FokQn+VgHIMHXuHlb5g0Gok54wR2GBnvVy5odqVYbNEVwFeM
ET50uLCIqsoQQq91S5E9ifp1vRmsVzmM4adyI3JorOU/EokbYHkTqQ82Rc8fM828
E3SH7PH69/HOxowfcwnBowOFn0ZWYgV3kXqimevH3mbPpkjneYVyU83sig/IFlbH
o6/MdT3WnQq8wvMI8aeWyrjE2efgRkTr9JTt1XQMu4DRoV87T9HUQw7nn8ccNAOd
hV34tBLhWeM+AP7oohMRospYC7a0IJc0O9IHaoSpD4yMUdro9ZDSueutzqrh1Il7
DiEX7PeutvHCuljclC9sS+L34EWgl3dP3hwP5JKvzDXF1bzdqLGBolx9k9NKRx5E
OpXLa0bnX+zrp95P/ZAum3nwrTd0g9qnsTYhl91+EFKf/+zct4PS3MF5g9orCDYy
SQo6+nUwW3jd3q5aJjCbaGSwIuVbFdDsfF8vv26ZJwYdkrHLIwD9leXa1V0W4FIo
+uUm4GQ0ZwBiWfv/HhOtizv3x8QVRjnKEfRUmvFsDMAZY24/Jk6hyxn0hAUp303S
IY1u1WpfuFWnkD2c3+udWqt6ndHJ0PkDkk38leAMSATS+aqiFLu7DBRcctziSSVD
L5thY4OzVK6FD1ulW4QLNwpGMxK2O4w437gkiiJrWeTfewdnB3dG/eiPkihrn+b5
zbZ42Ofqg8yExQNf+OKbfymZM27eGL3RCrz4adnIYlCM4tbR5uw90dD7jaWMYPD9
r1/m3qDAMPHV8GwC8mD0r6Dk1AnLSulWyVkokrlkaWyijiaUbkh7nLf+lX73WkeX
EbyZkthgUkn6u4I45KSH55Ykn0HPHnuJq6hXHhuTbwNHdWcSpkaRu4SvvoWgH7v7
/hfPZyKEWk/tB0GXn0+tHok1spNhJ3SC9ATUduinQLbU3rPd2BuIZFKA64jjA7W3
3qnlc6fkUe588iB2qKkV6ImwK/1OViGtbRYg4maJLYHdrlURCgSaRyp/5JRt8DHD
DNhQdqo5v27FndWt7uirAFHGGIsspm1ZfMn7H4K6y7dEJBnipWxTV508Z5XdUAVO
o9nY9DUHvLIsYf1YNaB7SFXf78tUnQ/tI4rVpfOKKwWlTyLSBJK7tbAmpg3GrIIN
uR/2Z18NnlLII+kLdyAaMjYYe9Wd5Z+CBOVrtLxpMRu+cacwAtOAjCcJTiOouF/v
UhybQx3DZ4hwuPC4VoEAbc7HBEsQvXiYctJy5EZ9JaoDt2zI3QvLMzSENci9bPBZ
F3Knrw+oqqOqu9FplQAYNFEp3nhGFD5r9+oLl8B8TTONGuyJG+dCioIGvsII8odQ
V91FgxeBk3KDlO0JRboCyMZvp+/E10u+IX5ja3mV61d2iX3ua2KAQ1VVEbBTW+FD
sFEiIOpF5xGGPLiOHPpAp2RfQQmiYV/MOyqywpyNyxn+epT+Mk0cvNl4gPDCWzr9
8qTdOWzpJi18EDV+4317YdN8mJ8gRq2nFR0CzBGOWDY+18vOHVr9E1J51LPx9sRn
DSKos7Uz52GHzW20bfYHlW/VKTG1+7cWl8moeKU/+exDa+eOIQvz41VmrURQhKC2
RfFW47trMhwXiG+Txw0RnpvO9xWKc/rh3NqLnm2o2FtawuxGhA2r8qnGF13Jod6C
RnFGRs4pvaU1Ik+3DJE3890LuP4NYMyXnqX4qFel9kr5QyNHzIRObRRWf8Z7r8A1
MyFo56FY5xb/HbxZrUAKXQSIHUSopvmaGgCPlIc1nTakgFCSQ0/6OOfvWO0Acm7C
pV8+hkKJmm32Obl6N8eYaz9YN+jYm6esCrqx2B33XG+z3yjfncJnYjcXlFM/Q5UB
dCI4p8g9/MI+0YkZhaaAYqf8yc83kjd/ocQQETZgR30CS2be8Vny0wJIQZPd1fAm
AtWewlK/7b5gNuzCesXER/VqqIa19n1lik2IG+nEmstexPt8AhPp78hyz+ppNyCH
DsLDwWCSx/ZJBE7yaCUYIuhkpE995L8XZ8lQP66GO/XIvrDCLCBj2mHUp3CIQahB
fwohq0kA1R+WngK1CdrpogiziekUvC/EypkuzPxHgYU/WdWPwiYkVvDN0lSMl+US
pMXPBEQ+z0iTP1kCN0TB9QK3X34DdcIWnc122yOtJtqY6hZyC6ygZfb/xJWryzRd
v/eV6M9Vm1n+/DJIIZJOgLBZuN592dTT9yNovF/tW7jY3R4XAk1613RzcSn+b7N7
BReMQx9Pu2ZDRfFDjjhQSNFZvrLYVYrC5zjC99l7EI+RjcAf/QfPIaJu6NWkw3yU
tRbckGlwQNa3bZ7f8Y6SK5gHGiQxR8a8x3EeKvHzqNcGGGrr/TZ62mBd3ScQvwn8
H+sUwqctsGyLtd9VPETKXFVQraJN5ovSe0mRpAWHhPS9gm98sBAE53Md3f0fEwyx
ni5Y+TAYCspf2/EQ+TzWR1DK+KuGkc9dqmnsOJJTCVWVApgCKu7aWvRJSZahOnQV
9ucz5m9t0bU4YKYwPMb/OYKaBc4CdPuz7FMU1VEgdhv+Igkq5nSqu+z8vOEdMNN4
QxjguJ/sgpOTa6PaMNFGePJo46xF3/GMf6IkQ6jyQQQrH/kTSUGiZEXsCdhII2KN
rleFq800DgzVOzjfSjgxERjhPgmDOpEn+tbkEetfrOyihyg2IhA5ifp9i1SFgJa0
yGGwN0IoBHX1c+p1LejMpeqJJa8HkLxGnKokT5IUUVkiT2W/iXXHpIuSdO4OxfzY
dD7cMSppg9GyEfR0nM1oJSELZHp60zNn186TIWxh/vEtxxng6Yvddk7G6V7uMCv6
PHfHP65Gcm6y6Rjx1PwuKJ/teVrtXsrAh7gvmcwHmbJsb02vtRBo3CcZrFlN+qBj
oGuZZrQuelIVQQBR2rBLvag9ktjvibOzfsRGOKKt3cKUq3Uw6SJiltQ9iuepCIPC
7qUFzm2Je/Dz7aa0IcZiJ9ys7H4FS05QslnbE/frM8fYgZm17HVHtE4rixQkIYuL
mw4tItSPeXWQv4hAk0pTwHFmvFAxly5op7XNhaPbKn1s8G85poRiZRmRAKnzVSeB
0PKLEmcsDaHY6gBHs+ZQoBBbHsjHUWpnqRSwgBzWofDGS4thZCvx3zeIDpmarzFq
vZ6IY6iiA2aQbBMILizmvZem1+3fnVkjDNhhxXiZjbYLNT3uIQAkbr5A1cxS5KCX
3TGaTtu4BxU7b2i1cGwv206J90yM7HTOajKaiNKQ1z7oi4u5B77o4jNbTuLEYi9X
6VuPyX08fPIcFqbEpmKMI0JOB1EhGrTJVVlom/yi18T4+CiNJUgbJ0lH10RNtNC7
YQavcD5JKjo31pEQfyLSXAGP2P4vG56cm/u/5Q3iqt5terc71EMlwAiBAsURANqS
zbYRsKp5f3m/UhZIxLbvR2MUBOnYs46JpJomr8H66g/advkwgWad2V+Dg//mnWdu
uLACBGwFMvWpIZPbkH4XklhckulSY3M8uv1kQGokmV3N0lA1Unvux2KiAFsLDdxb
pJNUltK6QALzyGcCTbS5qLsrv95BAdx875kjiUb8c/h5SnhAckuA0VVOZjIOcrEU
L/UAaWv/k40CkpyD0Fijf6cpcQJCU0pwlUdUEtZWQY+u/7XHo+DEnnWos/sqUAuB
ab/j579ge25RJuucATjCNgU3D3hfoHEcyjjrQW6kY8u5K7H3fsLzUmhexQncC9sT
LdtNJ4ncAcRKgXZwBFje5f0AuI7kDwKDRmtMqrEqjuidedeViZt9ER8t4D4RGxn5
q2boTUQZTbclf3ed5a+6jX56aE0gHxHdiBI4UXTkvEb2lykQw63QMtZYCgcX2xwX
uVdiYqjGpsOYQu9FJXabemlKALi7OIl51w3Xk+zVMZ8Y8z3xpc9wbJoeuF+7ubrg
6WDPumAc5h3dztErxnULBLWVvV28YGkgJ74P2Ep+8DoRZ65n4+tH7Z2CdhsfUZWQ
iCtdW6kBH+0cGoz3M0pfT7yBjgnlJmd9a/fQftUHZg8fMIhBoebndF7Qi7C1qa2d
dUrH3Gps+Wuel+N2HS7XWzETMN73pICmG9g8UZqZTZO/K/qAZmpnTpNvdxj85KrX
tKs7WJkIh5yrsrT4lflykqpuOx3NA7voo0W7o8uAbbBg37zrI8yCj952stJ1efQ+
npWWdCMi7OPEsVsZEE9pQa1UZLwLmRjFSgE6pig/z+BcsT2N0hTHW7zNpJ0W4yHp
2pOrExrjW5A3J4M0PoZPewJhV89jdnJbUyJ35/miPxCCtJKQ+9ROVrOHaGDnFYXJ
/dRQKVD11wHqZSeai3iwEaBlDOkaSLeXqwwbFQVhrE3WpWRs0+16SEF4SxEF1Dq4
k1AF0a5nMAeiL0gAfd1KDXJznEHnaKCo1pgnlHR4kniIWfCD5sMYKAkhoQ35HH46
+mVLzyP3osjseU/joI2wMuGM0+yGo73kOOT4K8Yd0WdRy2Uc/9+VG7XgkqH/+0y8
5UMjtvFnvzjoZKkHB+5QCRNScvz3Ep7hdbj6B8AL3CtBT+z4H8XEA6ov9V8n0yp+
5E/KFKi3sdIA2IGUDeTiAOclZeajiofZWOi5yGe9eLihWbGZQ8kZc3s3B6+1EYl7
vH7vvNqFPKl9wWIhLYXStEjnCqyb2aUNKF2Iey6AhTNTEO1pKOBMoZpwl4qe+/9y
nPj+9otgbJpkJuPcLWkZQcLxOPlPAkSFsL66Aash46cfY8K43ZXU9yHF9Vmb3zKz
gKk1fAVG3Rxf499DbfGXNpIkQ6Wt83z4gsL/2LljkmHrMHqxQpZWxAyrXn3a/cJr
AkVhxpPUwIbe6qCfJT5PeJ3teLY3JGxX2kFobwk5xwTiHPdD+EF2yv8pkIupe9pQ
U3x8SZx3rNFuqVLKexNduDTSnNQn+n6+rgbCvjoRzvYVh/8LZT4UJD+Cb35qFZnN
LMrp5f2EMrXZDvdmGhA1YR52JczSb8PZP2O4IL1P8n/kCq3yFpo2WU651p7lS4DQ
iijScIrGB7qIMciVBm9iMVio5TFCKd/Ilog4u6nkFNhkUTA5Bkj16lWViu8SZiTn
N11IkqE8B/cxjTPsVBLuKmajZ3uKcpLnruBKjj8WxRlv5lilKer+M41girxHk2Hx
OG2dsTy5/Wkr2yD0JGqymfKBBFlKTfRyD04vGnPv7DNUI/2MEaDv4YwgtcDAYyvq
N3KvIfojBnGUfIZvbBVPuNCJkhTtWFI53dIsPt4Z/K0FBHaPXx2iXDTYxa+4iAgA
rhIR3eTzurpiAXB+8MeMekq2/vF6Tfscze22iQQydVdCyWWpKRbnYemoriO32QUx
flpkTzh6FOmHcyWAu6+xuL1KA+FIrUjnT3lSlAOiQcLnXxeS2wIQkcdM8J5CJAlO
FFFRKrmy3uu80UXjcht6/BpG5mVfs5E9RsVxpu1qadXF9sOdfQa0p3URDyMiJo1O
epa23Fbsln08q5et/rb5uLccyPFnG0X2qEt3irQC0Sg2xeVmhwvdWcc+bKXydU9t
1N28A00pYu8knOYruWrIjdXyvn3z3pXOn21WK+SQIZKkkOqb+G2Yee43TXP4yqYi
cfvm84pCajkZHaA2szVjGO3PZjNZ6f+ARVPpb7+jI8yqkl4DTQF0hJGua1m3HC/f
MsPbC+F3hrmjpIGs3R0keIo2KQksegThrHGvJhqG0TPjbSzrNLMRWPj4TibHE3Kz
2XpDzWdCN1/Gc8ZdEfgjZ8KTVhZiSowtGW2sHpLo2Y5PtBzOLMHmFgVHrNHQrq35
DduSjWPGnja2lHRjDGyPXNX7BdWadt8zxAJH1+QeytdmTgDEh83e4pXWNZxWBj3Y
LJb/SHOrjfNbA1fPHjY1ieivUR3WxrvbL59iysCJ2SIN1Jzw9uP4diQV5UtM4pFe
i77+SqhPuMe4dQEXH6wrBzPZPLhkxqBlVpvapcLUThib1WqH/GkwIHfh0r3HUmaW
GsxI9Dw3Hgzx0z9NiwCsIJUKGkcyyPpGNwKAo7VRJ1MmEL4U5j3Bvhnha8aGhEWp
BaMe8ynpGp3oBJnVjGx3q5soWmS+eat8Lr60oZgXgre1ltapv/GoWfiAQmNG11ap
8CsQ8kbtco/3/Tk0nIgCRfWRTNeBI7hQJYKAMUJP2goI9uWufkJVngcGqk4LCUIl
2mIrubO0yBQrD927FghfB+kOTtUobCp6fJ6Jg/TsKZoY038ig1OOF2T62S0yI1aF
kt5BNvAPZVwuyzHGjJgeROgK4e5LMvvMSXnC56xwmMFZS6vwhqqQ/CFO4xUV5mdZ
SfXvwRfxvJKvqxf+NJESaclYvJUH3boLg6y2xLD76fjAY/uOZ56G3Zrn1p93zu/D
bIf7jU4+g6xVSGQQXB3K12LXK80Ja38mIa5x1WgkGyP6gaulIjP5TVKjqxlQOoRv
NatjSK/t+vio36LSIQYs05kUUZct3dXfKh5gQLnfMmBKU7UMXTye0uKghcMz6Jl5
Gmv11u1G3Nvi037L1exMh6D93c9e8+oRaRTSGLY9IFCKmEnuI72OkeGhKpIMwnbk
xqGWvSggPzVawlNSej+Y/loZwYbPNt7NJFg8hyKAPO1zsVrvxxZya7rhQiH/pLsK
KNRrfkaTOgQHLGNiWJRfqtiZu4ny8C4u6mvhC3N693e/DKS1EArpaVjTnd/Y/aSQ
8heBQwFHGUan1nvev3KEs7uqe1yoKPXZV/hL7fwOJPW4K8Ygra95TZnCJOYduE2d
voGI/wLIdNr9RY6WbSp8LZr2yqAczVpzdr1IL/upyUVraggMX+mKYwbY9zLiAk6v
s02e3YC5vHpaBaaLNSr6ofzKohh3IgjrbXnAn24ZORsQQk2KLmvwGvEsl8a2eIF5
Z3GKRT3KfloRM7RdMBT2Y6j7gW3yqyM3yC1keSFw6tWVHobYF/fLv50GlCXzemcx
1IqbYFoHJ8OzIJvM6oj7hVoIK+dK80v2jdSKAsuzh/Jvv/GtJwR1fnOQlwHYFcJL
XeYTo5ww1GKXBDHFlvw41BIndS+7CIZh1ClETTbGYzYFPWm9DnfVfnAef2Qx8sAH
fLyiLFe/+M6XEsi4e07GG1F4wX2zV39GfGWq12oo3GfQ26lLjbO26C9M3bNkPe8h
M40FijG732W2Mpr80sl3jBF9No+qyXTBT8yPlWtHcnMlkgs/ji+6cxd0F+zVbaiC
bQQufdMUMCtkxacCftWrMq09mvhoo1DvUrJgaDGaPAKqVIRTWbtYv6wMzyHzGMxo
jutYKIg5RYLi88ir8XeFzBeXwKjV2RB2H4c2LXgX86yLG9IlUgMVUA/H+FexX58b
gVoJ2oKmPHJmN+BwSWCMBIuL3vnTayBncnyxErAokPXcC3PGV/P7sZ4FdRWkrnYI
XhkerZPO5mtWCyf+s1LPB4qEo/cdyVHNvI2qiCiCg2/wyPHx0gVE4RHM/8mnPdWn
Q/hx1MQ8COZQa6Pe88Crwy9iLt5+e284vQXWoSo7JERS/yd1zv3NNoJPH50gdovb
WlzMRvAYxmKm4yTE/xyWPXtlvRiGeeI89r1MgApN9ZucToM7TgjWIbVc62inuh/a
X+Gg6geBJ7Ody9q/lBVpmwWB2FGQ/pFhl8NuJigBPrywnDyC+WlvVE2F/tQFV31F
QfCWL7/FWvz10X8DoPpfMODswaRg2bSCk4xdtu+Od052zqxJbyALd8jx+9g2thmE
FLJRlGSFgcABNb5HqmslTLf3TNW4IiA2ZX6mlvz3T4m69Tv4jji/juBY27orLtOA
edygao98kYQAJ5ha2U7BtdUGtiORpp7+B3S+2wV7NaOuwiIodzSKnzjX2qdDw+DK
Wv+wv9j7sO1khjpOVJOjQCmXKvSViBaL79/hu21b8twiWZaAJo2X94sFmGGVG37O
x6JD6LFNrGSFlpY+baTmv6rDxE6cICL+i5otIMJ8tQ7idsZ9HxbZHa2m/nmJt7+4
UVpIXn1lmlnYRsfa1Ecg4Q+M3vMsgAthkkYFUbX/AdENWCXzB7qRn2mcsoM02h16
+u3eDOAjlabpYgaBB7q1FQR81LOVU2cYO26XHupvLc3STzajaT2gMoXZg4bgKcbe
ZFeD7P8+vO3S/skmyHl4bxGoNz/zIyx9UfEvtEkZ9q+t/qGOX2Qtj7Ro6kYAZUuk
hX8xHmRGM6iyBEkTU7yYgtoOuRdP+nrITNydpMGNTQ2s9QXre/blxYJ+38+NXie6
WQovmJqfmIXtjLqXIGqA2fka0xYOsWie1jAPGL0BrIpMjTyjKEg1u3qxNrJAQwHO
buXU/Y22gp6iNs/SohTFs0XkyDhejlnHytCwiYwhMXzuVyg6gUsxdNHi2bc0Tpp1
VWqnOKd32tj010UVXPdbqZGdWc1VF0KXtiwQfYCX7RDCLxuxrIERkf1blWL9RI46
hmQGBcDz7F82vL/hpEEb/FgvN+X0MfG/QahWWEpFRvAsAUtFQPlBMKCFYXSkETrz
q9Pe75XHlS8uQzK7uZQ5WBpkU6Za3Z26TZTxqx2964RL4C9liuf4tOF/e6UC8kIe
d/szjsBujGVabUGWuZNyWIhu4F/O5ZpnYfLsFaKVwNi3zagTSTvFQk6zTqZMnikK
0eX/7xGnMMQgIrxjbCBxkjhi3R2vgmHUOPqbJPa4CbZJs2+ay30kxtYXywZ1BH9D
PLM4XBd9szN90iYiYwjcP/9DmG+Fm3OiQZBhYhszqgBlXbj405tipdC2562AEypZ
iYXLXeS/en/2iiaQCIWcAWKAGW8QBxmgqMUdP96I3KIqpkxOxbPpjeW/H0uCGMHh
4cbVRc7S1S8NhtSDiYB/sWLDFnZcwPBXfFKrmLQ3RPD5ts0FcXKhHUlWG8f2QKDL
/cBUNUABkLN5Q8cPzGXlT6fT76uwN+Co3b0D4j14nHCLPF2pFNJ1meImX6VyPrWG
QuBE1HgiJ5ngB+I5FUFibIojuPWP0SqbXDvWkb/UrP8pjQ91+RwyuRo/GpnsEerX
myZ1EOMoorklpXq5IAmO+qiTZ1wjrtie0ZFBc6DdhpmilhRkRqzXKH9pQcOCE5xI
fz1Dux7sGiyvCp9gwxJ+ANApxivA3QMrIHDU4Kaa7TgGYB3Ebdfa1ibM/7gFrqmk
pYDNt9ukDkF8qAKe6zfK+Vs/5qW3qs2MykHYzg8rLYajyWGBdUkzmLucDU0daSDd
DEqGVHk+Eqbrv3QFtPJQA4IB/WhTiY/17NR95W69S//0L9auAJ6YkdW2LhINgK1z
C0YhWCxQXHYIaIErntgqYHhvkSC6xRVSGm20/bAPdb/8DCq6ecbOQH8YLPt+Rn92
6XFcl50rPES34CvOH53L7RSEfHto5nMjhalPprs5+OTKK6vOKqOnKCZzj/msq/6P
XeNE0oSxYZiDJ59vTXGVtc3ROO8bFoEhdAPuF1DAW0nAh/MGJVhS92i6SPWYm1Mp
pSCBHfqCSP86wuO6lOW69rXn4r5oG9bfTi9IFkZirXatN4mE0jiT5fA68zKHclXB
Ys6cXXbFsAE3YqnTMw1yXY+9K6LCVKsKG1AiPV5xzpsWAG4vryKeUHK0pzb1zRt+
wBovY3XqhKi/BYhN3o3qG8/Ixw76vcT3ssaOJvICuVw3ty6UJcFBTcz7w1vkX3KI
4O2ryVewDo5mJqzBykv6nENUPAJ20Dex0hWS+RL8myoR7N1iYA6i1ILo6g26r0uB
zc6kUIcX8DCgkxi38sKzsZSYB8Z62hdGA6a9HXLMWrdlQ+OWdmfG7jqh4TAMUJu+
y05nEEB8wqhd+2GkdpFPt4IOmggW3wX5knN/loC39eEZ9fBT0mT8iFt983180UE9
/D29pY82Phwtr9tM8nQkYP60TzqQZH6SaNWeKFh5G7ojs0UPJYgLY17zIyq+qdMF
4oqiJwnW9RIvqI7io7zgSflXen4I027bE32v4wwxxjKVRmFvlgsRj0p5sjqEeCIl
k5l090RQoPoCRkjEFhshMaOBsWmAgY5TD4+U/ka3cmp33aXKcwSYf1qpKMTfYP13
unbWtrtU/FyJMvVePRJzVNquf2e6WRHMDZL6ifnXvRb9Ay1dT/W+W1a86lHaSyUa
8mMrdgAvjDahBTUHhfLGR89m3MijulqrBu/EYriEcHy9gPzR3YG5CGyourffbksk
xI/W5vxYoHJ9xPnhXwtXC2ybNkxABJKqxNAHdaRdqVYoAue2/GDsPRPLUvzImANI
rJ+OUrqoQRKb7wj+O5ruK5QEgIaCmBoH5lNSuXc20mfCKzhShXPRn8owBykh4MpH
HCUd/ewnreuvKeM+IxaPQyLybW3HwNfjflPibFHu1VtO+b/oYvXK1lM2ckw4FYfU
QRCMGAlOfpRN6YBhw0eTRW1fy9Hhfz3XsWH1oMz9QaMrWyLrwO8aaglRs8NySxaI
+NOA6j3DWbNvZMFxxyAflBJkOflGNNXTeXRcYXCnbp3EHN+LpQj7+o5lHS1D6UEs
rZghOdJDW2rt2zfGVm6q8ZQ2awd1f6SEhQtHroU70PxbVAFZ5U5auOQLCORf+6Ic
c6rNssARyzP+bQ/GBLSq3n0gI5GVaiV11TagrCnozg/fAyn5b5gG8sJPAVTbQXYO
1TLFuP8uU42ubYMfPjSacKL0wJhVUcSlbLJky6/wgfjla9r7nX5k0u7gzplhnwA/
GUPKiX74pKDAtLLPxq60TmYkkyQBtVKbPSHJoL/ZYUf1JCW1sKembQOXp3ssVMfQ
3N9S98CHSdgjW3kbTz+483vQgMrSnIw1Zj5LQvtCMSHt89UDaxKKKWiMHieL2wIN
NnFKCPrXJjofA40crWzegThxT5W4TRVLhRYafd88BSA3/Jng9yIraB4KzE3wQgf9
iXvSSxgiUbEDYHyd48p7auuEfkIpyXV3XqHiqqgaWuregW9BhPa0sxxKUBa6LwvP
SUqjeX5kc5hnZJSj8G8/cBCdKUohP51CuiZ0T0yL3aQc2AmbukCcfWV4X2OyZTY5
iV9GCp5dJRNI3/I8yXTBLvthGbuoExNdFTFk6lqpYhnf8YKBsw7MrbpTbidtBW/U
AOrIimvZLHueWbuiPDqbSL2MRFp4+Sf4UGCTIBE8LDdJrxIUbnnWs3NZp+1P3iU9
hmWUDc1jeuToakDaY4je9Vq7PRnOWy2aAYe5F/ZVFMRTrdtGdy83NyV6RJ+b7dyM
/7yu4ODLIM40bm1t4DADvQUhMVkI+F/Op9+vxR8Go3jeOErYOsJJqbO2sNqL+Wk3
rdQ8RQ3iiAzPMUdH19mZbANbeIZnxjtxJzO3bQNZvyf0UeOZlFBTip79HvWwCuWc
2qWGQ5zOutwjp1h43gFhh+UuDwzrwbsFMiWeuEswLsE6gIDJOvbtSUs0KaBjb72L
A+IoI0I5QkBmxXfgC1i5NNDfXCxY0Kl2SN5WXxsLJrhBGBEkRZoqRwcqwk2CuuwN
RNvanKJpaKkd/D6EE+cC30AwAs+BeDQ9of4tPKZndejdO5Ez6sIGWEbrR33BJiL9
8ZHqxWhYVv8SzMmuQwU5JDZzdInDbHYynKRK5WwLBCf7XL3fInwu2nmImQixDXZP
VKz3yuuAPF+gnZC/UU8Uy0Me9BBR+xqkpIojVqdiIAtlh9EzpqgBk0+eWlSfKdAu
Z6h9HDENAcx1wne5db7giIFf/o14y7t9p9Wxp4s+8avtjoby86zcn4rp43trcKQF
LMzWEfQLs5hyphmgsXuyvhIMY2ZsPOiZZOjuAHlFYAfmhImAqZe3+Vxnvx05H7ci
MhkCocisEXvgO/2J652Mxf8kRzYsfOX4VSL1LF/YS3Y9hzDfVC2bT9COpjLSS7nH
0NdlpkihdESY5GVT/0OOa5s5QULojGLcuUMJKUAzhFCS1EvP9xViibOzvhIj1pVc
Og5IqqaWvqc7Spget45V8UKVi7RhqWJ4Nmyst6PXlizequ8Toz807AjO8XIDcjdK
iq05HdYXEa6J2jiBuFxSLJyTCdDIQhFoGIxlqdrel58XwAhxP/P2dlQQW6SOQOm0
zV1r/akerz2G9J+DbTvyyXE+YzPDlBwdMjGtqI2wzBjMQT++cX1YIMRKAUoQ+qRn
t/RKijxKIzzZbIb60HOwwxeG6zAkpS6v+siuUHqhoaYH7VpO3LPMCUiYF+8TlngR
H3zeCy8UtV2dLlaXN4vtLiGRHE/2eJktLZkoWJjTfwRvONAyWyJgKVM6yEp7xZOH
jZWst+O2BJB/kV3Y+JtMlgfmSI8jsnx6m0QnDHbp/m1/pk5rtfDHB68B1eox3Md5
exOyTxOvoZFmsFI0+v2gGrXDnoF8UzQWSaE6pL4TIIWoXNOUvV/aIrXDtleVmijR
j9PrD37LTKXoW9lhV4TvxuddVVk28K0Vk9D2Byi9OXiMf5HagdFX3qCtOyxDR1KZ
4y1KzPnZ4NwUnXRtcBC936eATzuZ15w9nTxIeyqkzcffOo4ma9Csk4olrquTgbeE
TBZFPghdFwodtzry23aSlURezV94xstzuvCnWueLCQxT8XK37P+rr+vBgUIuLs0n
ZNbWxvCPxgiKyLjDXPO2Y70Zetr1Tde/8niJkCZTS920CvdMxUuXr33CZN4nAo2v
H+Kzn81jUslQTGKZRu3UR3TQX6Uuv3qeW4co5w1BhRgaO2Me8Nms/cBV9KIv615R
qY+fOaxkVqKGW2qMbRWZbGRuzm+iil0SMaW5Fw7vemiDYYvsGlbJQhbhUAEPLPbM
oiQqwk9mwPkvsV51/BHRUFr47QfPL9qz2ZvRXv5bJiovvtTStH4hQ+a2JceUsmji
k3i1u9weAVdgOSpGTTZbTVa1Gj+MPZi5ZtQgroj4aJbzVig+9nAFq1k684SG+w6z
L45mVtUaMjS8YF8hrpmFZP1lDypuCa0rtVyDKA1AN9akdRoXg/FzrOZIoy/dvfy0
Tys3CxSkJ1/TeETOLOKxEsG9pcwNZeu7D8O4+Gkw3SxY6YtrUbzFJiPzGdsCxnWz
rTwsR1XH8bOFqkYEUrPGS86VaiuHdXd7lhlYuNe0HzodS+t9x0Nl1zlkLPEZOXRU
ySaE4wgEWZK3qwUYXWdIHub3j43DqLT37yfAoSO2m+uBjN0tKi3iv8xR3S2K6keV
ZpdYN+U5AomZnq8hCy5fzAy1f9RUoqiH1XxJnEwm5I7AI/VRVslIE9U837NOx0pt
nzZW1A1c3Dfx1WleW1yu1/5DF5YeWIayBgX0OlzaDAu30Eb5zH0YiMqv3uc31NCu
mpGomWISBGPsmMdcMWlNMe2qeAnlx+WR4q2N/WJEsdc4d7/ow+D22Rik1krPjZ/y
/+1PvtCzoQEyciawkXP8mAb64TqNPN+R/+F+1lZn6HrgvOJBMM8K3MFoU2PMj/lR
t8YcmkQ621AnjX/dLAJsU/KGIAAIyDkmzHPDSLEATQvpeVY2K2ssdPjUvNOiVeP4
2yHEN/ulqFzu49Nt/PcvjEABn7fFmwXeXydYA0fDwCsZS9rbWI05BbX6bbXZIkU2
huFEH5RADc+pUMJ1RC1t4rGE0JKYK2R8LeAeJFK/Vxq9vb/yci+GEGbQt2f7QrEE
lZs2xJc2fVe4O0dA7iYvnfiCbl2Ul+RZzTJSkYY67GzEsp5rpE/pattx1s7ttKI+
lpMymJN06YSjYXLn313rVqEoPOjkeW15tCK9oIHHv892CjoVmH2srlhz12GtZVFo
uCAAWbr0xxnAXHR9P8V0gZ5sLmYI1GvLNXaoYPX8tmAUDZvGrvuabYPatFJQL1U0
buen9uRcazMgR/AARskkZFZjwcSNBz4wEhtCy0JHByQFCpdvZvSwbf3PIRLlb9dg
UXypdiHyqaU4fHBFfVZPUJ71e9jsUdvwSYDAGNjU31aNf5nzoVW+eWATYihkFsxt
C/0ChJezJ+a3vzfj1KXO/QhcTRu9dao6pEBeDJsKX7fMBLpOBPwH4PtyLX89prBq
6953as4Zxs1bGw/OVSEZ4vapWoFs4lDxPUVqgFRW8nZIrlXbY4+8sEliFWof4CrN
EjgI/utnlxtoIQj8SzS0ya1PzOjpFC5vqq0qg9XUfULJkDX/PRpKsb9LGPo76iGc
9+eowsAxP2aW9GAWlQL7/szgKF0/fXIirqOBck6qyJPtQJkSdcee5s4iKEz0H7pl
9wCvG/PnRrzSX487N+pYk1HowPoBmq27B/LvUzLI/ncmbvHgJsN3CoSXNdPaZqtq
qNuRe1Ldw2a/FOtjxk4OyKZXKBO9ncW3RDAFmXXK++W/njwHKYzOvCr9w4oVKcgE
onmC7Fbhk/mlBwk9cOLI6v1UKmJRAOgSJCOggJshOHiHnegMzjMnhXroM8UT2jIn
IiEBMMh5aysXw5fHcnU5wkd3ucWFC5/By8mxwbSqrAjA3mOYh4DfXkP7N/ipZ53X
zfi33jFoB1MRUCbBtpbuDJ/Rw7afKaZgSV6AWu33ZgxtMLVU6XmuJmWCLaPu1rCH
vf5voStgLMkITsX0khSxQt+o/OS6oYrlzFujEmMWrKwMvN3Vw0DQQSrhhFumrywB
w40abgamH6U9tBchctRVqsYiQsVOjF79gBvj0uALKptgI9YQ+TBXkT2t72kzsQMr
/vzbhpddjd2CgVIsDLexWQSV25GBYGVX4tx/KB4dxwDr/a9zN3aT74se516unDYH
sBYXgJ2xl+6ouReY8rvfIw5Jaws3AnVFzcj20uiotsc7GWCz784XlutD18jRCTII
ra/63wI66fpK94QhimM4ecqDSxMdgSfwdYtelRqliZJ1nDfs3gdPgUpmUTM3XyUq
XDXfXtKJKRzXtVLpe8ZqUDQz+6cqTZAPrsH39LSGZfuP99OxUiZAC/LbsJpBLplo
8H7QtGy4RP7ZnTN9G1h2IKrRiaikGarGHtMz0Q8CGoEdIKQYA1lr2d6xeWdyPblK
V39ixAc+qI0cgiWDhu+N1Bd11EQC2Kpr3P3/osbxCoLDCSVQ28vNCf6LpyvmbPon
VL3+rMAGflDrjeynrdE12nr5wRkarqR1njar9GmNnwfGCQ0+1nG1r2fGaTDWVSuq
QczrTLgrcCywu1jvbJtog4/wx2fg3O8+JLUOfnHR/FCVUfKbcbQtuQBtlHHMeREg
bHrkYO+aug572JzdhsOu7gOCKC4Wcw+BmkFusLVBtn93IubvTISCsReTj8xZ4pPE
bHr6ue/NrLnt/uh5Olo6VE6PGnECKwU4QD4oYINibvE7TakguIKGEG99goiWDUzl
Om+O/TCB9TW+ek55jRXflJAV6kU/eLMHXuD2rPYd6PjgWTjT1TXsw898yrrcNFMU
ZIS+20DluxCtRDJaZ6ggQh8TzH2rKjIA7DSgsnS7tJzUTDWYrUlKw2Uu+BhwblZK
0L0hDwOCcgjmvkRhz7NyixymO5ZjUeK3KQlHlckM5oHOLK5+hcRmJ9Qznr+H8s6/
6SRjQulK9Ej3Jmpqnuw9d6o7d1jq6UCxuxdLLVmNaX3IwE2sKBGV+IT4KJB0sK18
LqJR4fqbatKfVSc1XkUVYA6eJjcuBvA5AJMYZY7v9pOfSinTUiD3DDBYb3SRcE9L
A3aDNHlRasgs76acgYeVGV08ybdR1PweNv/jz9/uBCTkaZR25OIkHZia+U4ea490
sDX11NifW/pOfBtJ1M/89i6ItZoMC74qI8WMXz31Sf79Xdkqaf5TheK+hq9u4kV6
idcXPhTS5MsbCgkJA5pORbE5/l6zXl0fwDtxENJIlYJv6c6iBCDR4ZdpQzsivF1+
NSM+bJHY2B6YZ+03O9IP/jZhfqAYaW63+Hr4pOQ+6nIDSoBOBaBZ+xkLfxlr/hYl
bQ9BJ2GNIpd0r051HuwmGb1k/gxTAcbl8G+fsrMMQ9S8JuXdVOP8whqR7GgEj2AH
PyLsuA7rwVMtQ8IrzCa1hvtLPBBXR5HWrE6f73v/shcfZ3PmThD9pHyUJQiWyFNG
TtFDz94mZoY2Ys8pfODi/YjERBiKn9/Pdgfo1BjXDnyRvTdryJF8orYuiad1ukSI
dL5ja+kIiEzmmJ7lJXw79vPrMwlW2AonfZ3ozsJITmNwgFM63CsRdd2PIkChldT4
MWwza7mHbqA0fMqJqiGEBHzLu5CUTe8qNgRq61Liqdz6JJX0ee5T0iX2ppDrIfY4
DEsy6aAoOLcyT1Of1S9eq9zU3DAFdccoj2Hb4F0iWOsxxBn2lR5Lf8FnBMiLX6bp
94o0ZlCO7/zBd4Q1VssAv2Aouz4koDttuK61pmDuYn8KecQBknml5Na8D/+MGi5Q
Y3IzhZkdYVsAuqmFHN/bXN96fqLgR2zanaUa7WhvE/oju21O7AvOfZa9beHMFKxX
bQkTB4QFejS6WcrbkYZewn21GN+5YfdCOyiOQ8cQ+8b14LyLOjdpsPn1cttQNCRl
9QyVHJCAWaY6D0kl+bo0z/Bm6wMxU3spCxIVGuviCzX8pKl6Z/Yqt49iL43Vzlfj
Owtrrr27Ewgks5d4Jz7Sc4YgCRYQrxS2r76OSn5/NQ22A32n6LDSM1YB6XCJsSRW
5Zph655Tid0nyuXZ7QY7846t7ozB9kReUw3N6+GW3Zxzith53xsWTqcIxX3mDp66
OMVhhARfCImn1Yg2LM3MuMKNQH0/qIVB1F6UXpeMnIIzclEYrotMSeDv1vdLsLfn
kg3RhXBTFiDch8H6K43MUYTHNfo+Qir4kMUtjDcRO3YsjsAKdcjOo+Q//ExJEovg
CeUZ3XB+MyiIMH+pqwiZxE936+DeLLD4wLEdjAXPEOR0j0Q+2hiS/54BGZi50wlv
iBA4RQmnkpgKOtENipet3PEY7x5M2fKRCbp+8r5HrN61PkWx/mYZzUF83JvQLJfW
9/JvEH2xpju/M9eXgu9PYMSNMgp4X9uW3f2rcCzno0BKhe8ra/moDm+PkmrWRny1
5m8796eUbdwwUxMhRwc6T1fwuLwuRJHDChRyk4Axu1Op1aXDFCDKG/a4PV1Ck4ZZ
pFq1fJ3w1q9UibuUV7gZ06rUFvYvknZ0uNZLkdUzSgeBIb0icRuRq3oivl1QbwJp
6wMeZ2QqDH2twVQY73xb2b2xScKn26jTAxolgtkcl3K0J5uXlPX4Yg6AnhnrhsKg
hg7S23IQpZH1tuYIal9qifXCIuesq/EjGLNEveo4rtZ/dSEJM3UBf/hnDFsA+lwv
dxzrjeiwxGbKhm38qJo2pniYg/2X0zPLv4rr4tPbit6fzK61VWYfIyI4W/MTxtj+
S+QD3bI8eN3bGGR6vKdTmQ7nBojBu+wjKvue1hx7h8Wh8bENQnTXqHsXyqFmRNKE
FdgG7jUpAblcZOniWK3xvGztBL+FbXSv++m5FuVboHrJfIhTc27FgM7QOlEjldcs
bS5P4pnR2IKnfobuauOqJfshwrab8unpxX8OIPD7Ww9+1UmjmaPtGun7fMZFqzCw
kUDNL90gxvMIfRhu+QlOWckX4unsymGwSKQOBI2rkYjMCRHhaQFsM3emSfY2WueK
/ZnvR86KO+s0Y9KEZxx3t0RZ+54W8vn+X/KnD7ec4pyLRj/tBxi2LoloSvX8S0T8
Rs2UK04CjAvfqFfC7TdQupMJObw/t0U+1mBn6tbsS8Mzr9YKbx+0HmgsAGYCoEHK
Vq6uAH5sWYnatHYT3IUO3QDtYVLRc93hXuerOGSK/86vsSpZXEa0t/BIkvW9AE9e
O1sfCGKB1ILLCIupqxD9QJk9m5gd56A0AE17bGgj99vww/LJER9vk78jtBUQy3UG
y83a65bAkERZyryBvm6Eet51aH9xRGoxBrgRCZxiRZ6uowzIOdMsxLiAOy7q8dml
5ZkFY8yvCubyRy87u/HV9OEVE3kiIxsGUniLvwMJjcemFMMY5//X4XqV5sajtm11
f+bv1Yb3sQBBiEU85oczGRdT2GuSsy+Vn1gl1XrNys2rPWYZKfQuCBor7LJSuWUY
wmIFGIoamSTuMR62lG+NHyEJ8k7sySvm79+I1dY/xBEp7Av0qVTEwH6CNiuKrQAo
TUJQmvZtOQjyGEnytFVBA+beKV8wvkDW469VZZXaWy2Y0s7GkEtksyBuS7JmmfOo
v2YFLGG9WQBcxV0mFwSfj8fFo5p+8Pyklv9CEOt5FivI1j4feRzU/f/e0dfwqIR4
TbJhZaVjKhvOsCvvn6mmBwvX/5yOrT/bw6d27ljPNABjbRQmOAD+BE+gK2VclmyX
g/VQQHzefYcfdvW5FcxPAn8RiQeh+a3OQg6JwCGQ6TibKiVGYqFc0njYztB/UBj8
+1e/uwxm+nqRwfnNltkUETUpn87n5rwUipTBf3wShNknmwQTkwrK4/rfs82XwF7a
nkvAJds+Dj2OKn4yhnBlQCRPF22//PluwJMDUA6HgwULrFMplpLjFVMqOzMAxja+
+52WU111oPek5nwhBrRagkwGOReVlTQ8Ab9+EhL4OZBYmB69g630kZecFPLMtX/h
n5YJT0c4mn+QVrM0EMXF/dvfy58ytYqHfcTi/ebhDb9CYnKZEGqTt44Qfe/2vYIi
wNbQWcwbj7MHYYYm279iIDlgCZmEb/ChcSAmM+VKL9zUM3XHOz4eCMFzzjaKAZCP
pfiEWeExpU3178J+E0bega2pEsi190h70vurlXdT3sqCbDaJHQTgM/4OWe/pPUYe
yPN/yXGHAvL+3PvQKVhRSb7LBGxZ/u1ICbNXqEklWf40IEZcMiWRT0gec61xive4
x3Fy2x6o0OjyNqKOrZBLrv4Aq4uiNEtoBunZO8CPvTDLl1tI2Tc5u5PO02BUq7u7
GeeIgRPg6VTqSZAGvTcmciaFR+S1Ac0MStxgRIpwOUgVZtBiIBENy/KU4aQV+6Yk
uPQkf0Lqb3VxthzGXeGbJ6irujxUmJzy9grQetCPjwnYc+TLFmmZ/Mi91Kry0K8N
NNJrBZpWUgSK3LttvJy7Xitvk7ywT7Y/aGyrV/tH1RHej3fwPiBXIdQjXSuo9HMr
sjt6tgtKJLnlnNOC1YzWIFPPODn0F1N/gfhwcyVEjl3jJf8rNPG8RDHAubAwi/8i
bQHaSLNsU5t9w4hsALqYl192BJYmwo32CzJ10fRcsfV0wIY3PE5MeQnyl0ClWl95
CN70VVkhebP7HuPBugF05UiGFYy/l7ONJzfZV7pDXbbEZRPsemaFef0H/jpCMaqN
rVDFR/JG+ip2adtxkCk5TNNG5BAy5pqNFwsNBYwmXcx90a1+/gApdYTOvO9HQepc
HPvkAh+XQTdwKWXxWmbLMPC/UfhB1oM8NY32hinf3BLdojujWt+ne+I+C9jYyjKd
mTv/wwOgS/vfWQs7tp+4iTEM9IWIKRfutwK4heeMjah2Xnsk0g/MMZC0NTIlQs4w
DsyfcCdHekWk9kj/toUo2fIcmxDnTyJZc44pAzRv7SkBUQGlTbClIxE++Z6PEmbx
iWgRvxJQ3lAnwnbSZQHbZcZfXgC2K54SjxMJ56OdBNh9JLw3W/uDkrs1P7olsg3C
uJ4xV99q4BaTQiHwPnQvgv2y7z/p6ZAC3C8wDUpoX9Zg+vpBVG+0xNjBmm6/j8Rz
z17AD63ZgbmC+KiFOHbla6ELz4OvxSO0oQoJ0yQZ9bYALhjmSUB6MSgKl6dB+8YT
YyTH/qbbcP6WXnTJRYX/NS4znrUSNmW700JGynXefrLR0HcgK1z6cDk6zJhlXcPv
aPfdbjwqiSmkttYBnHwsKY2ZAyUTv1+Dba569f1jVZWiTrgmK+RRa/zAcmVzw1uJ
3iatExKYKw7msim4Ibw6h109h17nPXjQBfj4hVI7EATMq3yjUFhu2gJDYUuVlnlY
Y0G4R2Wilvrskz7e3uNWFjjEVWYjXZNUngfpyhhud+ssX1SYKceilH0o4QAy0/lU
SCqvzByihzxs3EN5+xe8LjP34fZgHmv3whu/202iCnw/EmfbvaLEUOLrlB+0yYRS
zwjMW6xYbd5/mvpIyyUu4KsXw1BkIviNiswouGFrc23GjR3Tj9dDnmFAhccb1xv+
aFxp59+uG8vlNZl8DTzHdWnKyCWcIw6lirkJqenVAHdyadjy/fqrHaxYXb3j1ElO
Aj9vTOuOabDXB4YchKUVJFcLgf3arak3nk6w/WVFcP0h78khT7Y0uvmo8mLUcYn/
LhyWmOEhadPo7HHefgM9F3DZznGheAuGDSUoaYzBttQs2u2w0HEvBCU0xkzv++Zw
FZw6zYIU9YOYnK/qjkOKb5QpTRNTZHO6eQuXilfVKSUCyVqPijzF+2dUGeohBT9e
DCsrvZEs9Gk0Zs5dhCEiceMF4gwbZrW5EvLta5B4UF5L0lQHhUuZGKNCi7KKQa0c
TR2VOsEUDzOqXiKL1urwqIkPyp9/sPn3dxyGVNIymj5lOhx70fGAKEZiRCsDk+Q5
0CIsYCK8I0rvmMQvHUlf40cFkvMPKYqEc/duD7W79ysMojyWG6kqfU8u+ZgvpM9E
vjuCYZBv9bCFMmJSqwUZBeZMEk0nVO2N38YCW8YQPIgm5aukRYuwXTW7ZW3WkV8C
v1d0nG6bmXliQYh4T6og29kS/eniIyV4QJ6bt44HDgL/foCOnX0uhWHczkhMv6EY
+CH/PsW6M4kERfbSGWzI2fJ1eUNXwdfcBcMTG5OfHyyBEsgvYFbQqOtvAL1RhJTx
RCdSl5iTBBCbsTTZ1k+0TlTR0lrSe55W5g3xy55ObXCgnwwNHYARmfNRfiVi0diL
Gw80pI/H29AvnHNmQaFZYoCsBwo0dQ8C9GgmY1bvbNXM8X35SewI4us2vv/cAHnY
vZsAhn/ZdRNIP7BIVWg9GBJNpPWV3oyJSSUOufQJxoqjtpXCLWAvcbLJpsZ+ySh0
Qw0EcPf0lfnYrajyIcrwAuXY3PyUM24akHNSv6BicpNhGlBA3tksngWzsYUuYSfD
0ZzT43hZS2ONJ0OS6jEkG/LuteHmTi0OTR/kMovejGmswbtN8/nkzXorNt+0IMNk
XHQtq21Wtq0UPTKnm27/zD5ua2Cmc0YOq9HXSBG8K4RC5ptsUUcaMvhSCeKphj+m
xCNipplHKjaClEMiP4XqTw/dY2uZsPGI4fWncs/jebeomgVDoFQAIeJ+d0wVdQD5
Uq7N+9e3a44JkjdgPOodheivf+lmsqEvlObLMhM5IncFQRW6H0UY4eW880kaXZ05
sh2PxtwMTSDyP2aUNV7x2W3n9dP/E4X8XZOdbmwXcT+2G1589BbO8RJ+u/hTh5BU
QaSqDcFMewL93TVMjt9bGC5mck0jK9HVwRpR3E7ebEN5+67xVPWIdGyWYkyiP7zg
KggeJqrlqJYTRGK7egBdLDLh8IDCwjJWnRbp3f9zbW+KbmbpDVFsFFYUdZB/6Hk7
RxOEbII+Depvp8AwOOm5P8av2MrO5X2paqpKBBFiIDMkw7TTwgX5xDjeOXyDYheD
USt2BLyoW7c3s89Qo9Wk0JdlucBTt25EtP3SgFHcy/8t/bZ3uiK9pY47oMA1/9sM
QE095psppUN0E6W/QZCVmIsO/Z91/4/9EHWPg+33dM5z4vROw4WBjFFh7iuIjYVR
ct9cS+BEQbyvzG1I14XdA41TKrys3SkowOU88fnXZGLQVLgNBRuEFOak8JX+UO1h
yxbLDOKgTzeOFmL7e7Xlby8Ctvl9xOl5ZQ3DMVhHNOBudN88kwJryOVcktzouH5w
4AOjQXcETUPv5iUB2l8YT1U0lYVYtqZWuUtObzAipxM+4K4DPXo7BJ22mifCoLKP
6AktJ3hLuUhNOECFKWHd0fjZChdgL7pROkYq/Zu1N+MgZVzBubTDGkxRcYXaJr5j
bNx4vNDdZCEu/62wZs9CvElLQ+W2DcJvcYs3zfHN8/i4yvjTDlPcXrebsnlTQk+J
0Jzwlcdu2tOpXNjee6oSGROWTRKV6dQZ/EJqmJTmwINyyDyg4fmVFzw4bf1Ons4/
DYajzbwd2MzBmywanU5QA1xmRzucAmimCC0NC3PqMKLqdQBhl8kS0YRrc4p7PWYk
ByiOlV9hdrmKFdBYuZ0jDJR8Kxnr+hPoqnJavcyjDoosr6XYVC/rlUP2pkthSxHp
Mosps4rkepZ7IIJI/9VjpVuRr8vMZQ+AbgBTOxUZxQJVrseuSU72iaF29NY1pCEy
f/KbJ3P77fYLEmPcB2lZBMUB7oqhrUhOLkLjnZMf8aGyVnNkxFOp+0t4rxpdfKCa
DhwXXd3cb2EZ3cKXYqPcJeLZ7CnhKT4pbbUmxzHWBK3L2y6gkxqodi0v4Mm5eq9X
5oMzLB9Ntb1oCGtjExfnfGiulF0T90h6kWJWwyReIIKJAOlUYZZxdovTZTy3idcf
tHbaAOGmxp2KfSu/L+7Gyz/9jFUk+2XuRFc0ZlA5e71vUOv4gw7vY+eQ5uhJ2h9G
CdB7Ida/m5+h0pZnegboWIhwkeZEgQTS9zWpy9xEjoKq8gkWq767CVVXy8yfp3sK
zI4IYvQ28+P0NeC4d5InZl5Jh+NwubboqEH84FFm4gTqZH4A221fqdIg2jzns0un
pvnjAiS9dfRwlLhMeg4k9EI5g5B+p3J75JVC05ZZ4S+sGvoqfMb2qlFkigY30pfj
8kxY5/ITb83I50gBtvu5qvzdj81UmU+wHJv25pi66C8KDBqgbzHAfozu1UUMxj6e
n/gxODhtG5Xak9wIpZEqFG17YIM0okiYISIw1YzF9xLiYrA5hWkLsCW+gwPSnLie
Z56toEknmBMkPtzVvO4HeS9OnMdbXCGpGRchHEHicrpCblKoLos3pg+OJvhBjg9g
5YFl87tn6HrJ6/Rt/++SkXV37ZSznEikDdHdFqkyyHpBp/jJeag1hzlE7+edO1Zv
2FslLJ6lJeXbhHnSje/qmSJT8+gnUNhoXzwZHcBtxjRVYF+QbUinEGuBtSOLua7d
E+vHaD5Aymzdw1G4Es5wLUKa5igam+US1WvSgXNt/jo5OEtHqYeTxSYhbDzzXgz7
f95YIxRXzoykyP4Dzh7zXZLs9EtSfTzAhssXskGjyA8wzsOPcyjHgBJzFRgL2/vW
dseEFLXJUtNZxgwK6nFpDa5ACMP99WKNhJowb/6IaYFLBYZMx1pw8HV9GIWFsCi1
pKlQlH/tYF+G//2UWn9FakAwOZHuUW98S9/CArbhAkN5Eg/8oN6jCoOAI1kx+0Lx
USppdiMzLEEq2J9VhisA4a5sg9oxXRNd17cFCNAeT+dOMBvW7Wxfkk++BtA+WWb+
22ITz3lMxwh5RDZOkZP1KPTaIPA9352g5im/g4eXxDDwyb/Js+lwZ6thjp3SIaDr
nTOjpK8/Rj76gvqVtJi3ptBpEn6GbiwwePH12WT7seDi0ERF0qguJbvQPwL7HTO8
h9fMllrNlMnNvDinxHn7GoGsaoPxmp3LqTbQJi5T6f0VMEAm/kD0BTaIV8sHYmkb
7/tb4IfCRKW5qwROXfNvvUWtwuWbcS6EfEyhtXvdHBkC43h+RrgAiOoKcPnm0WG+
bwYmxKFjILdffl2Gt/iiASkLcBbqk4ZFShOCn2ZE5lQZQJ3S/aNgo3Pl0f/45BK+
Td5LesCYGdrtYK6A9EIs4VWESIrBjP/c5RKMrSnXCQhPMp/hmLy0sH24Khp8WCvX
SmXu2izjLJwAgN2q/7X96X0xdyFhir5ecekeogpQvZd8oX7+ZElfnd6lHTpsjLEi
knkVifJOcKeH8zp9FF0S3ZrbFw5M2Ezpp0hSWAfA3DbumyiComriOpsHdFVaVmRC
mNvo2tRn6p6Vy+WOlUpA5OcKrnQ/V9tgOF2sAPY46v+7kPGEnFNGlMsNR0S7CTF8
+Zp0rZ0JVjhhzLtMot36mYKjIzKGmntOS97sEP0GA/eo54frM6Bb0uGTi+OIx3G1
qs63p3iYw8xQHJ5RmS1SaCh9O9q6FW2tuSosguEWV0+rz8KPn21UWjR5HWm0588j
+Y5kvidK13B/6VFM3B/bBQI2Y+dXmLbdqEeBfRIOGrWYTA8RUAcULaCEToXJqPSX
0iAi8eZeDFHcOFNOwuyKZbfvR95fxMUEriZIrIFFmfLc2v1U+Tvwvg0s+XkZ5Csb
fY4yMUoDOfOok40EmOAmEiNYrmTtvzzwLJItHsjyxjrRdzBBZY48JVPA2XJ+q0kk
GsiclesauVF7o0m6pNj7y6fS1jntGDM/xok8gKAZhd05qEVHMV/4bnk8hzggvBTs
IjVAGLk5LULeY05AQwUkZSHYUbmpEG4JDR2Km+jIThJD57BTUY4litrrT4LV/4GN
xKET0+/QCmHKPetsX7kExpHvfcmCIYUkSzQ0JlxcTaAg6fH+Es5QmtjhIYuwLz62
73Anv8zYyXzH9lazGjEacgOKNmkJxjVvA37HN+ahQB+tAfB1ZlLqbw1LjISaxoKY
pxlio87EjKpQqugymH8qp3/Qd3qcexXolBwBt5OX9t6fKbz7GVcBsBQNkzS4YNGG
8tUkS+8BW5lkPB5Gnp0P9Aa998d80QsAJots3B7KMwHopJJjvor5ctTq8blgV5a7
9OPohUjaBZbJrtwKd38ijNQCl9nbJttSeFlNd3DjxTYOEC1n2Nj7gltLgBg689WW
Q5y+YNN7oL9HXuEvOUsfOu5WtQlWHCh+5PY88tm41fvqAXnbkTnOQDytcwPBn5CR
Pnk1lYcXMXGh9Rqah/FLlk5z7vWun1fOvjAh8r1F6P6JQXRNig2bVtlryPp3kvSV
o5PzJTRBX8sWaa2xTX4jEvdcVz86rTTbwPCVgGbr9ang5ewrcOD/MamE9DRrT0vL
yIrouWWTQVtz6CvjNE8OkLgKgrrnVn/Qjj1e3rED2Flw6hSNjmOvfEafIH9ce5mN
ytxUd2rkOuVNo9abnS/HBP1kVgyL55NcerkUUkggKjsYH+tSwaHVZq6E5zsTRQc4
Oeza5y0mApVGcjwrcsIL0/UWvbGO4t1YQn0pQe3JPjwSBO3SIyrMinsOegsN/E8F
jzg98THYgnRTFA7i+66rUYE2heB2G6kU6rQ2XMJ8+m3mqCTDRzTyhe1GGjlxX9mK
pQeZUZ+DqnvXNrFBsSvtC0n0b8F12GPZ16Kh91OJl3WNz56Lw84mNZIHgUN+8oYJ
IKoqAUy/6tFptZvmhQXYt645TdWbEWxcK4q4Gf2x60YuO8+l4Mu9xYm5N0I86hvD
CLLOwvCAtfvfUaCl/ZXI32GsCdw1IhikzkrGPUH1eOLA32+h1zqF++i6n4dHC2R5
FNj7OWP/cLPKFe65wfuVJE7hKomoOIByTLq9+RxQAMeIajtfj5TonKuh7/cWMMXY
h0qRNk/enBEgheI5NQf4u958EpscoFmGWQ/9jZtrRqsgMy3z7+MJWQCk9/AptaFH
Sq5NbJ37q/JScw90ID97pvSnhQpXt7iczjyid9FdkmWTTZBXFzQK59cnLLK14LOp
xARdKqQz2i6PWuC2rYwgcxYMsOb1pRkqsst6s14Qs/zguuRw+0eDh05ZaKqpN6pe
J1HDdSTzdXVNglzT4oEFGkP/YqjOz2YuBgKqfgRPM952SvGIvtBB8XPqz0x6fu3O
kj2ClsJ+OBey0mBWQjM5316TjYRiobBcF2qduLR6Emi/Pz7Q7/ogsQkm/EPyuXyM
gqMQBD6H5/6qRVRkoBZXTVzK4gqiqa7ph/OWtQVV1P1bWf3yyOTnqdm3WnH6tZrq
eDM9m6jz5sc0rBB0XaLF+C+8TQ7VjOGp6HUVFlc+orUNTYLZNXk4WH4BBxWJWCfn
tdzckEqsGdW+/L5VILNr+/em330d0JBsCj2Czq9Ehu8hLfC9IGBmO4GvRLoID3vK
ct1sszlMcZlqFwcPuBZZv4XEga1KPjGDiN4/sACdr8Fo+ADQo9aFvDAYgQSf/nsB
wGN9JdG3524kTmbYIF0LjJZlc8kckMOBbBuU0TlWFAB8VYY/67ZqNm6eTFEBbC06
6W6JUpOrFlWEwRxz+P+xB1HWbR7ZjZ//KwTWJNIxo5CiI1p7sLdnNGApUgD4jW/v
4STQb+V2aRT/SvrUVAR0Z+jDPlHtxxMQ+7Me8TpC83nT04bAqq8heEbj6gtgHrVV
oHe/mKNi4j6YkmmiZUoaESxAygGk0JL5DQvGXpXtxBY53lKFDVFcep62P/IrrOE5
14KO16KPIM7xD3xCNQ+DbheEEfkeTTmPTcBpi74Ee0nYM+CNlKmOIrdMWx5DAOD6
n9vN5WKgDe1f7fqrL2KWQtjSTgqPDL9CrZehi5ZB0q2inyzxJpfM+V2T+2ZPDR9Y
+2l1KCmhOg76vZ7C0PlpAENlo+jFWnLGmbFmjww6If0rpJPXIcTJ2ajfmg9OLO7W
GJL2/+vIYRMJyxfs7vFQ++xao73z5svV88umyc3fCQnPJROVCf+AbQdX5b0PbdO9
0/GM3lh4qjy9GvyyAVyikTgr9BfOT+OoD2tgxJOJ5oU5oNJ5/SJf+bBHEDUL/JOH
0cAjuZlH4rtnwLWmZSjv+JxaVKlHePtZfZyd98u1KoI/GrYyfFIdNBgsqkwoGrdr
fgmkEMO04+z5HSdATIPr3kLbj/A+1XJ5aetbAxw2bx526Bh9BeauQoOxVfsXWtQz
e8LOQIRAZgapUi1UhhVf4NWIlFbxXvdoI7er6IUCBrhnFuhotKvodP5ERw/BKEqQ
1EyXHJvoKqox7IAY0Hnl9zAwjsXNDbRLGd3PMId/vyYDKBd1HnAabeDVmeDC/XRr
jAq9SrckzxY1kDaUd1jhrZJQZ6ja9dd9ZF+R6L7OhHj+OuI0qzgPm4syxwE0XOkJ
frWB4y+oD5Os4KM5qQxwSmox6OjeTLN7V7DAGnHNmk4cUxR9PPhfFFLqM3wKzRuX
PYZjLu71jjBbxkOrHz8XW6gn7toXdE5uLydaUkoIbTFj8IkanWN3rN8n5lao245R
pZlFhV+IDoguJ1tszv7i2dvohg0B4t67CDMZMpAuxC728pt6P7H3mxRjvoAdTDNV
HEYXBPVAAYHKjrW7MRmMySvUfVky5Dck125XkW8sMO/2R57FFWdWaBYXZXwZ5LkF
TYrvRRdfEqC1Fv07A1UHV9Yj6nssRmQmNnkxaoELTe1/RQfk2kIcVzvHVVQ0Jpk/
juAIHFdspmxMYt+arGgA2N5/szLcYF7tPyMTtzI9j+A8EI6sVWLbtQ1761LpacBf
pc3T3/g03uSDUCxeDAQHyLbgFWA62qb5lUUQKGcGP3eJlDkkxM1MLf8a3vrgLcDf
5ofgnp26KC77VDoB6XK0VYn/kNRzanM+N2vptts6S3S71H9mHhbyYiN/0Isp+MF1
+P5OZQ+S+2afHb7jgRI2/tEDZqqqhyD8gharbvXW9zZTA5fvF2JKFwta8CjlvNt5
63986SzIYw68rjHf0qqYvhm06lR2ssxGZ78MJ2hH1+sGBuvnVMAvX3sjvdZngBQa
YA0g1JkTo+dHi8m7kVAXzvNO1xuMmIfTNYbLi8w1O/LBrhvTzOpY5NTL+fim/CuE
hIOPr6Kt9lnR47ZcqxzrYmmBAgS8SW8+9zkgQVBcgRiIkdDq0ukHcVkKO6WRXK1r
Oq8qZgjG4s098ye9MhmMDaV0UrNaE2IaNhdOnDF5D+00VmME6+6PB6XGDI7pOUOy
8J6oRWdOwMiiUu0YJvxqKY6pjAhDvSbI97mkexHL9dm+mBCbVF/CK3Oxpc7F521j
sOUZAkHa5TZvSISE6cXa4nSgc3TeSSGDkl+j0Mo7dqvyh8UaiJM1I7mYJetYVcuO
uMmD7TdoBD4Q6QjakkTuR5yfBEtU1hZaQyW7XKd79PQYHcOkrdkUxU5cbL0pae7D
+xeXL+/mEJ6AVzKI6E7oZxIiO/9SMYZ7RYf9iK0wZsngVOIxZAorLma8RPAEikjM
/LVov6jfHOcxd9xjXYjpuAIBE6gz7/tjpP1srvx446sN7pQUSrZOQXQd6PfnaW8U
FCMwT1PHSgq0SldfAa4rmj+xR9bqBfIkwRFyqkaxRKT4PTT3OMNXrnLgKJG6kSFN
UbBVy5oWLHlhrFPUGwQvAulh5oTJaqBC9qJcpdf6jItlyRJRuHc7kP2YrDtvQiMG
CElwO4EJK/Kle741tQ+zPUAfe/KIcxpM50FjA7MFPjL0O7IIrhlocfPNwaitqK6I
bxfx4O9FLl+NUKOt8ZsaS2+KP6cekPb6zWtanIWZLDm992OekeHOp7SOUzZxH619
n2FSqlxscobbZjO6rxu4gTM25qaUzlnvfg2WiJsggDWjUvEZlrBBPsb0GZ45TbMZ
tZebnO+deOrhujEQ3XQP587seUXZpXh+VTSWeI+EdKQImdT2IF3I+K0z6/LV9KSH
343SPUWUxBZdQ6ayr6XocPtVoC7yFh3VG/oYUGBC47DVdq+vp5zvgpW5V8wta913
Q7mzrpiqMJreGHnVUKQhBnRINf6fEQau9Jqgl+MafKL9WTTe5VrZRpayfPR1Z8QT
hD+wNoFln+Sb86aYDMYH4Pi8tD8R/6UI3fVNqvoBRbvDErzl4YiWnVFhOUnSrvtk
wueciLpY5uXpJYfMPUX8kAAcDcWRxxqa3G5dknk2UWiAzciERl18CrZJOr/9NBkO
5jakyAvfEUNoqGwL1Bh66UiK9fZsvVm+9qxhyQXrAAVSlx8iJJhUqFMxFv/tF0JC
NSnpNn07ToaiVxG/R2qNvCthpUUAxIKo1xZokYCoGp6GKiYL6YGk4q7Ly8i2dz7/
pELZ75/C+Q/El+hFUiPHNJhJPlSFxXchc4zqfHcsDj7OSoEQS7xvOvlq+z5MRRe3
NPELvFn3pKYFeHNhOTBfKJHNj3QvMTUam6kru16oFr7IrIjRjDKGYELHSoQVe5+c
eIB6YwmjPnLU+vB99IhCfoefOgmYqXnx1QWbLndiHYM21+1icf0huNbbYLLQ61Wc
w2cqSaqW0Uhjx069iwk1Icp1wMmAkaPiiwEdvyK/DDmZNgRkXEfxjHygXkm2mtIR
/E0Y5RkiKOJdjItrB44VyIiDrvt2kxZHf2lxEcqA+/D10Ispa90h2NPUm//DCQhn
QPorcdgEyfoODdGb+kVY8Ji/uMXCs9bj/XWX32al9l13/sUqdDsXAIH/kbch4UUp
Enm0Juyl8G585LpM/kifq5TACofmaP1Y6+o/y6QnwEQpHwe2oVTIwQqCK6jHWkxb
nEO2JD34glIULDm0n0N19OD387S4Ks7y8KnRy5vl8e7CiyFcYvKFw0Rz3nmHm4yA
3Ub8RZfi8ZNRRuaVfhh5kUhvn2FM2WtiBXliiivs+MyMEtskR4NQY5/47le9oWt6
Cgb7ppRgnPHWutsgQ4qmnT2pAzqZ2iBkkhvsn09JAoV/x75CRnAL7iYyGSb3AMMa
PMXEXuFJjWlDohR7PekerjzQ2gChlzm6f52HkQ/1GwT/KjweRMk75XDzJthOq6C9
609UiXvhETCfCHdslTGQ1CcjerZFF9NZ0ZqoSYNybXyEDd4AUgySpPwXUJ3cZtnI
slS7ypTyaH8Ns5S3W/Yf33+zOH6A8kgPpRUHREpssQht13kE0R2DLpx5ZyJdOiXd
GXW0iSHFuNlds6yq+TsD8ypincWp2vZTvEkcyyEiG/eyHIKQ8/E2LiAlRX5V9C3f
2/gM7IfgFTcv2rsF0URB012nANCatGwoF63M86osTGLZrtIXXwFT3b25//D2FS8J
Pu/LX3i09blMvIqxyePJLFJBsCpsEjQkJM4OyJzdvfg/3WaZ17fNghTZsGICpoYc
ivAVuv/NOHMgsmK4HrGHdTJrzBCbsB9byYvaaeiSWCU5j6TYKnx8rdIdzzWOqI3A
h6GGau1PoKBoBgHZQdCSzIoWN+hwoy1ZSxQwp7YBLt1bFJ4aN5A2Mpdtp7Ke7kF3
lkr6pF6gsIxT3Abj+2zBuMmwG72+Wn8fB+TFr6vzy+4vXmKWZmQTfkWv/sn7KyIv
eHvi4mrvLnIKW1uoGmr8LvkiW0til+SGRg3fsqP3QH+WY2ue4XnrbtdqQJwfvO31
wA6esi9KIQS8nLGZGdTREpVgk10pPZ5yBkZLVx7UdqYa4VovumDImthbkT5z5G9M
RoyEIKtcelUQ2h1sZArUT00vuQycq2yfAKnQYvcn/ko1YVMa4tz+4kKs8DKrjZqi
r7qaRIAiRv6zSrS+aFcXYpYjxCoCVEMMBgfsUyeV+oq6KDC1TM5QXAPqgUjbw3Jw
4ccwWcL1fLMAJZGZVx6jDVxx35DoosPqu/bryvx8s0SYxp97IUupq/rmhL4YGcYY
lDu+GBgEH8lIBGzutIKdhfqCG2LBMv/wYuCt5LmM+ByWh2GbG4nYrhQ0uZe92VLE
+zPMz/OHymV1MxdyJ35El8PNojZfFCVz9NV6ov0b8Fd8Ulsds2fyUrGmzEfTJwad
Zvb2rofPz0NsPQyjiA+8gsBTQgWzRNOVZyNcoTaWNhaBKYJTq+yBityANdCWQE5M
orVjJTvjZVfUYASYIkgCILyCfhGXuHVbTL8hwdxm/utsrlhdr0LYUfb5NWq9Rgor
ULpteh41F1P1YRD9dPu/CO7aZtky6Cr33kg3C5RwWLj2C+bM+k8wX+5qlCcSlDXs
Y4za5g6JPD47oex06EwV4g1xWb8ifpUK60WTEVSROzMMu9EAKJGFsSLm524ItE89
+eofJujXo7ywko7UkkCXqSZChsEY/Y2EsMXpOmD5JNKeH8Bec3wm0m6CYN8XJsEq
20Uc1eFN1sCthfrut95pGX/rtO84thXv3KvEvUWsPcrUk6YKt1Td+ogJAYT+YDmG
f3KOtoodiZY6uoh+R61nFVXUYy8JKx55WybYB36V8kNkiNIiuLP9Oy0487e7igNP
qtGWlVRG6rO3WUrUlXvCVLfU1DoixDHAak2UlI17T//CQAub4yjURn63Y+iAfZcX
RI0NuHG0ZXxxzjV4C5HiDqXgCGg7Kyc+BuxS5njQoTK0VVxWppirmE+JHuiFTmDu
SDg0uPwKro8kiWu2eQ0VfS/aq+b+ASMSd7CiRdVtIN1TSCe58IkwARfGSfQa0YgB
krByKrUNJ9JmU6P8vTdGIJdUTjliODXy1frwFsfW4i313yAUHKIB8XemZ3GluhNo
udGnMakVN02vaNdR8SWlxQCcy/+icNQQ/z3q3sCkH25NxVa/nVXKhM5IO4fuTZrO
I/g2+zGMyTru+XJwtPgQCf6Gk4VeQGh8cfRNheZ38xDrwK/V+I3WvL9bCIB1SIOF
B0MsgEqo0ke2zlDjHEiklmB30kdpS0E71dUsOpnYmjvJSCKHO3g2N01kcCEHgS2+
w18TB8GfcU5vojShHtCldYIKmsf60Ic+XhaKDPhqcgp8pxjaUHB28LXOdqroPExu
8vg3ZepUM5ia0xylKxetVBTqltaEjJYDgdwzyeFyOA3HiBfUv7TQewATDHVHxDAj
CLkN0Anc7YaunC8z2BZW0TPRZewCnndV301Xsg8Lv5mo+HZ5qXy/70IG62qkvJL7
tlTvBx/gDG3L2mUNP2s3j8KN/wS23+gpOmyHW6Twy4QtwPsuZAHD6+1h/Ib6k8KM
sloE1zjOM3LSPlqc5HCHCM7uyO5FuOPAeQ8RvRdZ8XoIlGQCaEhOO9vWMR/SiALU
pmGL8+RwfoAgDL9mFC5IIw3bWo5tFo5ihaXWLkW5kUNKvDpNoQxaAScCzwpj1PPl
iYmtP2upwPlS19p2gU/1XEUVYobj2ggE+1TKzZVeDoBBJNA5yESbQXG0QWbiG85z
ve6FI4upHio82Ls9rH96FnjtDK+2jARmDGfn+2+ZbHk90Uvf3wmTL/prdiWvTGJp
e/PZSx3UFo/IeIeErZKNPfn0zDNddC1uB7CF/HutsePzT1+cNFvm7wSbOLjJ7P4H
Uuhy21ik1uBWv/zMefZ3ndaNHgq+yH4HEg8yC2+fcEPNeSDyzcu/FdLiuQk6fwyr
31G9k6K+FFSGNpqJgqKr7bHzUrwyUjzcaewj055XMSOXf6ALz3MkUPd5eoBUsECp
gdTQ1eyY5X6YOM5jJ6iApLl+2G9fR0ARbdJKnksMoHQ6LBrAquJZhPDSJnAAlCxr
31AW9PVlAjLq+UIH34CBIkXLhLelMvjmin43iMZR1IqnrRjM4aYF5hxMCM+I8VJz
8RAh5JTQoqL2RhtVG0+IUnQ+iCcVThICQq+deEd2y9CS2nLJobw+y4rdPmevNg40
Pkcrz9Kre/kVPOYwYnPibwC9take7XRV5TBfBmAlvSqKj4fB3PtKH4YbDPC37CB6
WKh9xhmoosGJ75G/Hoo1nYlpJ6pw2P7xg54FFeH1gkTuy7kPGVUxEgKTrlHFmwQI
6kEXMDvhNdNiU3+JUBUtoZFmXgp3Dwd9O5cJpkM2Z7540QZ4TDEIDvn9gXgvAL3+
P3lL8C4yeYxmZdwSzTCx63t4r0BI18JVc8Q8v7S5dkCmnKkpmGDWEhCxH3uQJgTb
E8ekZUuigzSp7dYSzeAgpt5k1BAX4wRW2zVLnbRe/RnAa9qpKEZ2ombHJh0iovn1
xXR+CFMm2bB0Zjacz0YFYf8vpNP42Dg1NE8P0kK4YpjjK1r5oYak/7Zs3PkD1dX8
vjWJv92DRnPzEzq9ZSAmJJEuWWdh27FfGoycUDIPI8Z1AgV5tA/TpoNfrBmkFyq/
LcEYpizm2HKHlyLPjklc7JLnkh8FrCd/PDeb3GupnD0lOb0DbsA3N425iPgk0K6W
bAKaBHMwTUscgPCQ+hJ+KXnc7wwP6ImFep03LGiG9PB94BwwV6imo2zoby1oEiKH
OWCBoG3VGLED4l933xm4iBvl/7/6ww6LmucnTNeP6JG9hm0Dg3giRQyHGWGI9PI2
eWBL550xPny9CfrPY2IYuxY5Znxe2XEQ1sI5tHJkI6nTY3cO4YNC5oKK4kCYLWhk
fUIvEwT+DcsTI5Ix9gnxAF8jNtk0dMxTSbUFrRH1agA1rtsT1yi/ETbX+pIugaW4
bSx5O+osg8N5u8GShguyYWZHBVl0CRtLAQfxuzup1t6poChPCIfyzRTE2igmI4BJ
RCEcC+jbkMtNeZ+rHZDVpkMK0tR6VlziGxxRfD/6+uy5Rzw4K8yAC50dYxNM33Fa
uq7QUICgI1U8GDuSXRUV6+/MNaCsfya7oP5T6Xu1RAE74CSGsGAkO5k6Hobbqs6H
QOnTg8z7udKpvkv+odxWKR8fcBpYGBfoYNBbwnptOlWDBU8zBWYGo8ZYPidiRDd9
HBYBuLp1NGr3sNyxn9RlGKA4Hy4G+qqj0dAYurwG+gkVxRrvw/nDF1TnXdCFOfcY
add1dmht/hvH9sZSaSN/dmxVojqIvjT/62FHHs/D7fa/db9lDi4JIslxPcLlNBgD
NzHFbHLuDLZIsc2XnZFc7WXbpkp3C/ZiogkfeGNIBYhXWeXGxM1yTeb+yGdu4d+A
b5BE1zmZKb/Gl1ZHOwc6LpLlhsCM6DJumMgMcQRRbH50WCoj4Vu2KohRmq+QJ0FY
YJnpE3Sonso7cVw3DwPSQVbdH4g5LJf0YksS+xSLtU/DovKR80REhzyxXX0uRgl6
TDR+KTR3TEeKlze3Sy7vI5TKB7n6pUWlTAILaKor/N4irQU65bc9+aAXWuNpnEXZ
rwXM8TZOAMJATYXVAY6aystenYFBcW6F+SeBWUZ76R0x7GH8hw3LgTDsrexwd+Vv
TazTQN5cyK/g4qcqF55N5wyV7aFxAXD0BLT5lmt3Or7hmuRIUCGN/Thef+JiChEg
O8eNX8Jb8mwUfJPLVxXQj8GgSl4uHJMNVpWAVHnaNNcZ+pAO5X7MZeSmnEcJR/rb
ONHd/+I9bTyVig+cyOaFtd3TMWFZuWzjQraMiLhsftTVeRnGZcyt56Xb1bXaDAhb
yUK6MSfnqe3H1OwnSlM13gxjqxMEEw8G1A85j7S39uD5M93g33zHg1Cqi2R8BTBm
PkxfxbyJLz5qpm0GhYXxaP9yVeZNkIAiZfeO/dJAL6TjYSbVpvkxnq9vEukEMbam
OMCmR5S9751pqlsXQJ5ZqItgImCzbfHnMbhEneu9A7WfhK3jPgOY5TodymqXfa4N
uPOx0Ky9exohSJFBADmMJiKAy1Am9XvEWfD36mEA++drkmupv6yjWgY62q6qDNPN
k5ogu9IF2NLqxs6judn3vwNRp14XSPgT5WrwuYrcRX4l1d+qYHqbWLDINWzQQaSd
vYLIxU83TDIhnrxLpemrMkFUsdGIynHgkmvSOypzpobTh62jl2yybfEOFc4z7gEO
LFLKChVQsQ3FhuxHs29hm1ktyf4k1qvK/Mp5zK6yiMBDDXY/G7MFqiJGiZO26Azk
wyCz9t8zGBI1xTSy0Dvr4mfkzqc+3pasASI251fIdk7xV4n1KoPhxfFgvgFGFZIZ
QzejeH3TIleTqmtg6nhgp9iwtcTQLMh4QkijyuxR/kNCObtUCetzgpSme+pkhW2I
Z35nZ0MKHXec5NXY3/dOlarZlEnrAZEvmMWaVMWCbaFZ52siteJAFjFllx2ZHXZj
0Rw7xJhn8EgJvEugOJUNco5CbPcs/dYpm5bpYBu9BD7WX5QWBxtCUB0Ujcq6Sx1S
9/diMPKZsiD4Yh8i6ENOcP2WbnIcuxKRq5Q6Q0tKa88v+YBSudk/SiC6WmI3S0Bv
eRWnsA/kW2VwC+WyUKn9tGNk6gQYRrfn4oK/iVUTrhycfhB3szXHCDpRLD4iywAJ
SiaMZYCIR3IzithkovBY6m2J5SzqZwdPm3ubEnSAJTvTRsPGUpWY/pvhiEipVplZ
+UQTZ+vMjUbLQmwBYgatEpa9eOA7NLDKE2xRgXwSzQX5lhoVwHue3quVNmHs2Rld
MkkfgMJ3DiIGj+6V4xvsRl9uGrUybmr2oEESG3m6RN316uSiOwyaJBzL+lrqn7gr
g/2NZVO/nZHU3+ZXTGHy0nQm7SfbanK92jW6UHv2ZXXt5bPszLmOxeKsJlH5BIs+
ZQsrvPX+/4NV+7kZYkMBtqDV+5i2lMLN6PMH4jixEdjvLX3RPp4fIb0sShMNFBnP
Fs5ScdJcLmML+uvj4PuKUIIUVvDolmofF6HYsRr0UcItjV8FTS40IpGymGufVSDN
kZLr1po4tuZiSfUz9H2FTbEzOKplkrKIcq1+fu+Ix0GP+cZRGULo1OADFe+wzfnb
0AL5mGh+RB2aYxqAaM+liyAwr6wCPxfIkMHLYO46Sqsg3lC/h21H2Z9BDFDxEgmP
cxCHgfUugirM6poLG6muhn7E+wVMVGIwHW+JEyyXg31sY9dVa5c/vJPX07njeHkB
RjllAERSS9GmrTjHAznl0Jdg8kN1AUUeb9ALwIe5NBL1hseqz7HVTEcnkkjCXpYu
9wrpXVl2guzWLuZ5ymJfjfy5G4U9T2Pf5PU3AUYaO8XvpydrLosqbRgjeTZUoM52
MZnY3O2JA0ISZgV9qds21WKbFlMLLOoRbkYQHTVycsDgZA5uhN1cMrTDGUqSOsB7
NxCYAjxi2JN23q6Ie7Wd9gCCL042u4WnPCyQShAvrs6zXb1QQ4+OVnbCm6RlE71D
HzS5bgn4jX+OTXtgE0R2BW7h8v/r/4UVFk6JR12ybAA1/VMTQxclrwM5nCzsJnrm
AS6kb7Cp6IPgNO6hbAN2tThUch80RBnSNJ5TYM7bf9Isqo5L2lyNRCV8hPM2/8Ta
DCKmGrg6llnKnjLQoZA1hE6S+WUZOInxMFp6Tew74YShYpmUSFe9oUilvXbtaArf
NrGgrTjroDpc0C32wEPM6pgiF6JP1evE72z82teEnb5CXe9tE1DNDB0ZhAh8XNTJ
LqYs9KmridwMcNBwoh+BUVx3MeCRQ3q2Ip0D4qIJibX7IuAoG+KIDWwsXZPmxdfg
afXHDNn/mQxICINAxYDSBXfnECYqw1cCiu05O1kwc2T6/YhQhc7K0cjRXJeucV0N
lRVQyG1QYMswnDwDXWgmPGvvJaEOIy2j7J7kHFkeqOQcGyRY/1HSCvIvve93P5Ay
kduVjLM9M1SSsSZ3LUVrfW0Z0t2kPx3nubjsrvc49ypu9H8Bz15DASD2VrH8slxC
wdFa7boNXy89Om2D3T+YA8Y4uImFrSe4/3faKzBRImDgkN8XrbhQ6bZX8Y+GBNsE
b6LyZefIlLzGK2Nzav6+/XhpeWP9/1p9hJfEAZH7s6+tGFVXUPgxGxmRsXh+gmXn
KVJ/Bx3NF9MvRADjuSJMR/rvfbsAI0W9739pdok8pWeay+RfcIxsQZ7Ya+iQ64im
CB6guCCzojHr/+KEd6qhCGEuADdWbz5Ce3vCaOwEYsjZJB0G4HTli6vec1VusvxY
9U15BawZUGfYy6w/W6mLqnyLq/O5RRnEb15avWi0UFkRn8LTYLfDYYjk3cpvPpxx
CHDztB/xJffVP9UlgEXw45BP/XG7Rcl56P7evSnVPGFFrDQ/On0ZsZ3yo1cWyPI5
yG/EpsOAiR61KPNlolCRzpx0CFPbyMtV82BnozZD+Nkd4ep5awLWSPvJwJZZv+rU
eku0OFCHpPJVeVAFvVwnGPJWriEJgq0eYcIZO4uk642w3fA+aOhY4PuiJ3ZykNm8
n+vZbdD7zw0E/G8g7LQoevCcRSAc46fLf+9lvfM3nxOOCH8riB7EobEazfmPD2xi
kOZmhoNM/v2iLLi3+ZFhekdbaYuNeoCYHH10k7qVVR8FqpM8XGt4qeGxv912oeff
uLg+PqJEA/vOPp8c+zw7nZ4AY6AijOxcVri8K2IZspuHTKq5xHd90SBOMg0yNjvo
6L8WQJ7DXTAcaqxk3/GZSKgHNv48avyTZ+l1gfwVUaqdk6EV4Lvr1xHS+6yIW+vc
VUpPGXv8qI94ixOFW8GN4V+DZ5l6b5XN9WHCyJ26vEBIm32stt3lhPUqgOIQ9/i1
VGYxsQWU9K067mq6f7U8rRGGN9gtIk2cYaFCl1RLciHESdQeiJwAAlYSbxAJY5SR
DGIzksi1Ti5lsJKl5U9ctBLbMTJkOP7HfoSYdBkY3mjEJXZgDEH94opP/dgp2MUC
fWDN1OfbUj3UAnF+UFp7RmERhgj77mXvd9amQC9E8UhkOVjc7E2KSQ8tqcdPnEXT
z/ZfvmD/GCC3f/HfiJisRwRkOmlJ6mtlNMpksV2M5fpkugS8HWlJr83sXYiAmSMl
HVKIAyOHjLHm+Wmw7c5/GvffN7Dk/C+jZuIGxLCdnrTOfFJqh3uxmSwxwP2cb15R
8WUZyNmRE4YcuXgBe24zpqGmYpo64EczlXaY2MMR8Obs8CYJQuC08WqlhTalwO0Z
y4WtBOq1pSIW49rUl+X+9afpZM/Gq8vb55/7zEZRsw7lM8thWnREywWtnHjZODRl
5qVVMjqyR4lJafT1mwEbRju0A5tloOlo9XyuwRSNJPMono0VVaO+Rq/u/YLJO4kR
6oB/xrzAkWRIspiigH194XWNEENcDaXeKYblRF5Dn8kuhNUYrju+q9IUj091kGQS
uuMjD0PQaVgzRqYSam59IiqXvLZehpg6UIClHBs6JGQJEM7OYZXf9hUL65otFX+R
SeuV1Q7oHIFrWGfgkdj2iZqrQ9oWkYVX2QF9QauLiLKc7egeAgqLkvND0vEVDDOX
/q+Ifv2AuNfneK0FH4IKRJBAqRSp8NCCwEzKYWe6JvYcgXhkxBvbfzUa4pxHHATn
TNV4IPN9BFintocoMzmt+MuOk62Q0sT82YhoGZjUknZ5W4oxaqVq0kk3gy7Anr/m
dEV+rw+q2Jfujb5XY9Sa2umlSUI2mrn9/TW9RWBvmBUFrHgH6fWVOvqCKvPAq7r+
pu8kIARawLVhP0UrVOvc1TJeDUJb1sZi8qGwHNXWEACmbkVHrkAMRswbqH6AlBT6
SkC2XdiDd/XRCfpGrftZUoI5OHPws6oXXIG/B0IgRbdyhb1EG3CMkHigxkq7Zbts
yG+KKYHi6Mn5pgJsBsBjhjHL8I4+9Au0yEnFkUg08DEkONfPfjO6niOuOKaHh6u5
M9Sl5hKS82sQv8eylkAGg8uA/6NZuucVTG7wea0Cxr/ii2gfyYmcjEcRdk8gkb+q
m13BfuQ0ZlLbjuAjVv66JGFef9RsnY9GJjv+Irr+uv7mud6SB9hUxXfmDxrVJwgG
YVD1h/PUnlphOyCEMgHeKxULgm/j6OTdoD2xCV5F5VnxWxN2aHmVrLJ0JiPNQzso
m8fD49f+HFwl3Fbkxmk3IVQ4209U01+dFZ8uLvPdiL9tHNrndJrGvqqS3/4wfexk
CBgGq+BnRsFY331LGtMe5cpV2bkrp99VAZd/twhmxLV2kpmjRqMDfdssm8Z42jUB
k3jeM1p42PZwJPheiN2RzvuhZ1NmEc1IJ8eFhzMLJXMvGwlk2QUSTFA8yHq7qfTk
+N704OX1s9ISq9ub2WAyjH42ZQ3jgX+viDCupZxdeIApItjKsVeMbBX3pAEKkuBV
3+GmOhuUuxgLzzwo68Lv0Mh1REbJITYqo1TwUOR4TBf027MmI5gHvSp4iTdrM4R4
xiwrOJ+W5kInBF+BxbPguN5ZxNnB28c8kNHrcnS5eBfU9qgfwlYUQcOMLW2Yzs1i
7rARu/QIJ15hDkic2HFuVTZuuFEFU50Kbk7EyfvY1/0c1A3q2GDtnJzFDGold51b
LIuH9M3SRBqaL/C3+tdsv6gAJAMm+gO92wmX34TavaSowhoelgPGoLmvaWZaeZTP
m1SjL1X3bKYkZcVUdKzdKO3378Ec/SzVCnfIKWlaAVgk+0HikpdwPDq5OUzGUoT3
+TnbX3cL0tR3R8ol6CJjeVJJbCHQmBt7pv0armlAiEkGyEKLb8CKG6LcZJfk05AI
QQtTH9VSoJgamn5M8ML7RPLnfSg9zRcbRTEnhPDYKt0bKBIMr9GdO1LJzvUCe4iZ
AYOxQmNLe/reQmSpownfUTZakb00R39McaL9IML8Jj5Id0RNrhhP1Li4RQeUF6Fd
ms5RV55o4pDTEZtDbg4vesMNhzAEpsesCiLvC3qWxC+7cztwEwHjtpUeFWwh1N1K
TNgo3YeUbfL6802CQdoq2jdr5ZcggBm5HSUY17O8g4gvIRvFL9qJCVoBGmRyPVbF
RYX2IEIywV1A4IBRBrr7BeHI7wnvkzSFSTMMBrKex5hJGazOmOg4pgE28v0zw4sn
dm2c+PJc2qxe+3CZ9+R3vVURoqmnXZaUnVhXrI1JWzUFi3FgvoRGli9fEL9WetnI
yWO3bvcDarFBpGWGtxAKOaAdFINVhMdc3MSIRJUb0poVRKPkSe5rEPEgBf0MC+NS
Gj8sF9NmBqnod+dkdqZTG/bKQCFdML3oypIDVhqeIVU2YXwl9C/R8Mkfp5EWcEZ0
zvOIWc7DmxT5+RcXVStrPVGLEa1D1B5Na/nYKyW56cCRW4TMPma+14mqB2a+s+m+
sr4XiAQlwBIKrfAr7cO1m8UURVi/h7tZmYIMTOgWm1WVSg+WvMTQjDUDM7eKqv2p
kWnCR4mZbBObCG+1v+u0T3VyXAWapzEDibVR1IsgE+VFsQprUN98c+5YqSeuAOqT
1T7fTXtlac7xEx62IoMQewACuOvS5S00B5MsD47gQUyok+g1A/shnEhEY8h2wPNh
ZwNjYcsZ6CsTGEQBnjwT4qFYZJsjd1NpY0ZFns/Qv6q888h9bkILwqcdMd1uH431
idWEl8YecyNajMMet7j4vsQ2AZ3wlmr7Ke76m6H25IwxSBHKWLwuAnh6xTHaxZxX
Mxk3wckq+g9EHiASbwHl/5/YImkps69AwdJiMVuuiCTlVLThU1Bj9ji++SgKj1IO
ZY1pZN/AgsxiTJsRfVQLa6up+1qwIfQ+JxQ365DP7lehfy8osYf+LGTkqeRL6vgM
U5e0FUaihLgecK4yKg3Zmo0c0ravD2LTD2qbr/31NvQ0fRYSyzaecO3t3Isn5W5N
JVo007n3N13LdBwhFMOua02R3gGdgZIZvp/5jIhZ3G7Fu3TpnEgxzrvR8thPvE8p
U9M2zO2c2e7/Ixg+TZrOe0VEw4Fgq0WTwLsfmq7Nnjeu4oXbA32CBQv/Wmava7kB
Hy10iYjEEGw214yJGva4KUa+QZPCwXpmsO1xLH7ry7VnCebAL2j8KnkGRXdjS0Ff
XMDqCDNSjmrUREYWCKDEFtwOutaqgHRXNqX1JniaKFmMV4GQlx7pvd1qYaxSpDFh
D+T5tOQv/prWU/DXk+MPtfMgW+4v5v1oQ1iXCdf9gMtwRuqZOdFecf11KivMP9DZ
WNAPd2DF1zv0cdvE7T8Bj8ZI/y9IhJn5xPuD3Z62HdmvQTvLTHW0ZZkyqCQ54VsS
w5EoJRY4bK/zav+7GUW8usuXFpH2kNcM2DGJ4B/25PpghLoW48T4qVN9K38+fUeS
VnCdMe8Bdsbh/dvYJQV1vZXJShnqp7ZizircwzZxktDiNUQuVkLwFi+QOLu292In
kO6qInWz5ip0G1tsSvQpQf5MZk//qEDnMNebOJgfa1g3MoTu3vC4QWHdB61T9FW0
/2WyJZE5OrjWHfmfuilhtKIxIGhAskW5wYkrXKRQU6EhxMs31attTgs584Utsnwx
qhzv4BlYIDBfn/YUD3szNPOAYyAA67WQs95DJq+V1Avz21/DnmJ59V2d93DYBKCK
kHAJbx6/dMS/sg2xG8woYVhwQIfExS/IOEu7/6UZEi6jEBHy6YiT3hVCBrXPRkrU
Fs4GbCuNMX8hzbHLGQongAvYou40FoQy+Uqv+hOLkCevbvKItQ5OnZKpm+kxYWKx
danxQ8wRKLVojNhM2yHQB63kSXJQ/oXFozs5iPRBVr/1RD99DiaEUiJjeUEGQnjp
GxA/ABCdnfsHBlbsaxKtoGJHDbBHJbmuptEeky6uj3JL81752ZXhH2TjvDmvna/5
FORMcCSexhDdhW4eqgxPxbzHs7i78hQswnu/8pNLUdlCEsnEq060txQPo3FNj4WQ
WaDSA3xtBPXN1G8+y2MjzOgy24mWhzGRbOxk/XY+795J3jacCMv4fj0LYDe2jPJp
zJ/MIuPPWzXUyV/q3a1ONuFzLEvtuqAkRhC6u5D6tbxc2JIuXJ/8j/jtMybg3L0A
OsKbCONpS/ufn5RoYy9EyJ0655RUuBNeZ5dvXvAe2BKS+UCT+co1TGXf8r2UbgYh
yFrY1GeVZAFB7ERP6QrNWiAT+dwFMRl4oQkNig3HvZIpPBMPQtv7JnY05LXPAO8x
YjWz7g5nSlJvuae+XxfWoNUikPl+h2bO6nfI3aNMi6AygnB30+oXVhrrszDDh1Kn
QDLiUVIotc4DKUTF0zACbna5lXJggx1NOZ3il/wJhT/ReWzZ2z8XXQaIJ4JzRwjq
FU9EgIIjmSXjkXLPDoI3JGbISt+BJdcRSHmuEIsAhCoSu3Fzj1ZpnlSe4xCqeiVZ
+YC8J2nUTMrqlaaecLe/MevO197HFpdziaGbPhPqNzID+q6DpHEOtZU8WYzsn1YT
BKCedq9uT7GIZ0erqK4vdbhbfEVZAJpGUNI8UhkJjPhXUNQUR3KRFUnbpTbH9sgu
U+Fenv7mODE2beEZuKSE1V5VLrHQjqPrEcgRkj3c4tMgVnNzZSb4P2PTXZMwa7lD
j6HTi6sT7qGOWShfJdX7GGV81HcyYMRlBa2Q4nt/Gs0a4PSUsjRZnkdO/R77C4Xr
tVWdi7cVLRvazPxF6nQNLdgxAgWw30CfdIY7iSYOiPEBR9jIfZUU7WZF38Pb7SlU
2BeLMXzHQcMXmR83iiTGi6ILYk2MEIbXvcvQCqyps0uyN72ZWDHWq13qEQfMxemB
mKFpzDWCgliytsNS+r1c1+A0CyVwd9mIBDbmt5/InPYavEP7lIjrsG9KGdoXN3x2
EpFfOTvzYUlRG9snOKIzm2ql0GdPdudN32cVK2oSV6dAu4ICCPnoRrkZp+yTjdJc
MqwbyMHsDWv6OqldbSkrP8haNPyO8shef/iGFESymj//GP2pdI1Qk0bYe7THS4Qd
BruNqfrAXbw/yJsgaecPQMKCl+Yo981Ti8XXulpCVoMLPuMWOLp7h3xpZZwRausF
iBDpmDkstpwkWePePxxEuwSOUM98/ABQ0aAUYpptH3S97jkOYfBIDGn/O5QmtzUG
i1I5Y9yKfZfABSJFnHGRWMRoslrpPhu111HKCMaHZsMc0QdY2idHhWBcsnsP/a5A
XB+TfZ2q1vJj9R/xGOrTufo1kmIPqfRnKBXHFjemguIyxoNII5x6HWaYEQKWr9+q
D4XhA3wLOz/kIw4y0OmrDbQCYaedsdOZCc+6vQ1mH4yJxl/nkS/ZJqeQCWgXUido
UIOkk1qWw/RrgvDyCXX158d72cF9C8spu1bEmcwjm815Kss09bNcAecpvyVgkZt0
uSdSGx7uIc9qRxk4C/OAzBIgu/MWhn6ej6Z94DTpPrjM7PGxw8Sx0Q3dXuCE5/6s
EBjDtFbgSNqQuKAD81g7lOPNOnoxcEM9S3fLtZwz/xs1Wrffwg6aLd/IjREq4n1I
37ZPiNbG4LWU27PBwGoYLwS1N3L+vOGbyCkpMjiOfHkn3mGR7LxFSj1EcTZQxwNp
g7JTzVIYT4r7Wz+1Dw+x1cNTZUWJUmgLBOaz4QD8VyQ1Z8kITokdokwSArVCmFnw
KkLMws2n9eFHmUYq7R7QHYNEf2ChcoR4DjctGdDiWajjxS4kMEWDRDt3bL0z3QjD
ArI4w8yVrh362RXC00Y5qnD+GUGVri6h8qDaixElaG35XG1SGCcpV0bqBV+eDsHi
RyMoCLcldSglkE/5b+ckJx/b0GRQ+5vWaLn1dD4mc/5j153R/b7eFIe7HbDXDjnQ
P9ZT72xRioYkFPlHj+8kbU96rIi8zE67mRSySc01uEQythhnaJbQJphwmGc74qv+
giLYKraZTLOJDL9+t9ixPpwjsl0/X1Ytgx42fNgRo1ky4KzIWHMhTw83MIQzBfvQ
H0e4KFKGAtMNDttie7suzbSq9rILkveIJoPRE6ariZH7FpEnFxkpWC663mMSAXbK
Qz4dYtqyoX1m8vnXyfOkcvgpZ3TZDX1RzBEhHX9gkkekzXWYCGeultYjo4pUOTX+
xZPiGWm+uXY6NHBx954Gz8+M39Ljyb7VUxkku81vx1aXzh/AF+TpFsgNDqiMaBbB
7B9TGHKhiPdefA/KcpFx2D+ZJknk2ot1W/7EvIISOkOC9ENEB8SSeh2i8o1S/uVO
fwModbDHJTkeMshKBt1k1fBymT2NgOGu1hLyBOABDkboAiE34NAIpPEIC2G0J3d+
tJf94PBe7wSZLFiIJIomtDjjO9Tchsz+kMZeii2dIL+Wrac28TFpizvZYYwoef3g
r142hUFmsg+NE5IiSi8V7wevteMt7Ai0DC0/ROP65V6+Yi/IOPQ7Y0+l60pw/IXp
MBGRANuuLPkwInaMGavw/61XBaG10BnYvY33RVUTor+C8NNBdfpZs/3vIkA/D+ut
yXwi/9fTP2JuRxYhDiRz6dcQQMyumBAvCDQ37P8ipt6wgqwUynL7OiFrWsrO479b
FjgBuziPrco68/34CdjznwRnWicHmvYM8GQTFOeQ3ieLTLa0N16KGipMiYbV4fu2
bRO/t9b8TIRW0WQ3tL3qoR9IDLun8uynb4eBPUf1AJxydRZu9qtE9irPUHA3Qeq3
haQ08n9Cfw/y5BT2SLyC3okRtOl0xOv9GS4Hl4BGJCAprzGq7vABTYGE5xy7lrPW
osFtfMceE1w0JMXGj9ViQnfzphfU7NcYyc3k3xZFxxrZg7pLWnI2c4vHI1nj3KJ7
3QHqnX+0RWS7BfD3v8WdAcKXjC5/9NWoxnscsPqf9pavOxdvIUMzsGkTCmh0DGF9
S5SQ1ILRd9HagG+QF85aSPoXGIIDs9fWpZxBkTcdUv1SEUniOj1Vwzq3x5zpKfcI
9BYm3AT8nJJjKe02wF3WDPX+dJC6NvKvhffFaeUxJnY4x49ZUiA6q7QU+ZGxbuOv
1Z7ujD6z4SPf4DKdn/yDRVZ9BHWMOGdNFon2p7ipu25lr/osLUeM95W79+WFfqNm
9JWq5LEOoRKkBHvjAr6NyW8xUddaqj9/fOs8OF2co5tlRxgtjXsLO/Z1n+tNyE1u
fXicESv/yT6JnOjZvlNM0S4LfIFKrtcG4XOmxtIw9mknczgQlt+wzqO1Gg6JuE71
4C4HspFFgoaAIsOFkYHXAcOWOj3DGvptb8R2LxhOJFU9BynMcGFkA5htbdDIeYy0
uRtlQ0D8Ae2BSYB9bD7rvSDTFUyLV07p7BHiIlkZlb7Tmh5Sm1qjxskMSGTCOFml
zQ87OR5TqVSWzi6Qya6SXDD79hABVLcZEd8oXK5Rv3TPpgIEw6YjqxMuzcXfoD8/
KHMwwV/A8IQBS5ThSGJxsG1BBDzxnUO5N9/AZQIhRLNEO6GqCKkbLZQbYuIy0lqM
2DNwEJXYqPkTdsNEkZPejc1edwPNi5HWscK5LePFGp9ozTbtJv/rQZ7IyNnG4mji
CpEqdpZ0L3mbfZsDK8RBjKg24m4h2q4v0nOikdE6f/C+tPOjsD7v5AO7kTMb3ojw
rbuH3ZlABoyKoUteSw/II2TMuAmtJL4oey5YNbqEepoFbF8qyGw5HvifQqf1fBhP
BtC+3WKVujzOSeUT/AioCTn3d+5t0tgy9oR76qnairUi0KEQaT/IlgSkGFdXnyBX
H9YCerbkfRBiA3+Z028uCVD02+UfACAQtLbOUir7vyV0KQXqx91/3jFdJ3a2G44y
orTeK990hyDiqV6TbfWz4rB5HvIx87fMoCpNdA1CRKlHBuu2K4w8HTKOn7PPFUuJ
56CQ42qLkIDlxIPbFtSjnf1wvA+FJNs+8zhdyjfb3KULqmNhlTOKyz+nEnC8q9pv
djGyTzhLVF9Q/hvJdK6X9AfCN3SgUPwW73RRxPfGb4LqwPQzFoutqz28jetR+5mV
tSGi7Xxe3ZiDXj+N37vRZEzV4t4G8x/VGGxT24iVnojAtFaEfyHG1F5AkWEGD9AO
zuDouaBfvjK1GH4U1SbLzOS4Jtm6YPlsupWt+c/gdpyG0G6TPYIK1kVNHtZj/5k7
1LgccG5GwIEqmHTr+HKIYHthTZvxXkO9bMzrGwabZeaEe9lCcfmsl3hQqSqpgwzH
T9YUbRnsOn4nCj7yHF13v6i36TXZNfIObTd9qY1Kcsjr0MUoP0P+SkudDZiBWLs7
pI9SuKn698v+dHRyczVvsltXJyXgCW1YHbFMmHFjQsPgwphtZW+LVsqPNOoJ1dA4
4YJPdkZ3OlTLkOItXRLG8j/lKFLvHWrf6L1MfZMnmdTgjDVeC+lvoBfSZe60rq4m
1L4RH3fkuX306GBEMLIYC4YFS0G+AfZsQIqFrdmht09ljqXB3L/TLoJR9GzDwbH3
V4mzTMK3mcxTbbKg8xdYADYy78B3dZVaAkwSFRTCYmHfkqtAsK6FkTYTzPiRJHKE
GVbzRnkXRCdjFY8Oflm8wCa4y+HlUXRT9+y6PQPTTIh1dJwvHkUcrqYh6giRflfN
OlwEKJ5cRRuReAKpqZZm8yvJ4LksMOm7Ups3qLBVZbTzvvSyBS77Kz8cf2gtEnC3
WNfP1aOHMdAyEUKWyQN425Y7Fok8mhqp5B0SE969vU30WOxePIr+Kr8mEcHKMblm
ZJyBeCsqwV0Xi3+tdyDnnFZEx/E+zCpD8DRVT5hrcw9sSuBxqWyHSV6faLloMkBR
gtIpwD6YEfHszeaJAGJn4WbL5gegtbMPoje62wxP053L8nUC6pVSL0uwJD+BAu5e
tMw0N5zKvhLwH6pIZauH/iFxsFKStl+ext4yiOhHK4rn2LJowlqQrqflAn0dkYTv
jbhBFPjMIVX2/5ReiWvEaa0aooPPNPmvKqKyEqI1MaNLkGWoXT++wTI96dD7Su3e
2636B3tikLELI+DzVZLlQKKLIipOIL+XwcB9Rn9QhLo5AJI6bJmSmzpMjj6CCmVV
1bSJSkPrOxa4vsrA+m/FV7Bi2QBB2s9nbuH4Ci/N/ul6E4g63t2V9IMC6g0epwn3
4BrVGvaW5pYNTq+E9aTLCDucnID0T6E1T+cfEBPxpHJ0piBp7KMXdQdXSsx6SEKA
YuFL0GgEX089aYxw1kP+TwmIR0KOzPJPg9RYZMAWoqVwqsI+0bB8r7VfdpOUEtNK
D0oQUgyAkyu4qoZYlMnajVeS86ZrH/m3c1NxPskr5ewY56cT//m6a7jRqoEuFRym
3H2gJ0pRTPVgulKsjItrhl956Ldf2z7bUi6g93S358uvoB0DI/8FKHyKpf+v954F
LcPvnAgaX9Os7143N5h1Y6rO6yCjv3bGJN3HcubvkRfblCotiHzeflFLQ4NIx5jk
+CIOTZTJQc1rII0twqNijSrPghmqsCLZSWHpepUost77b1zKt8TVuzAId29ZCcvw
O3LZkJb2ctixbfjOEfih8gHJudAz25p6ZN9JvQkCgd46POCEJ1ML8Coqv8vp+VV0
7DbbxEtgCNFBT+hb2GqdtusuH2hH45pjgjt6f9XLi5SJqYCKzkFfKJ610L5WYmPw
uJIcuALZN7/ou8le+Q7x9yHQNia8gqZauXVdhJwye0612wMYLdBizcgaVOwwAcZR
L/lLSRGk7HHvxW/2oTBajTwD1vXESOhjhztuXLccBp8FWMLhmgK0lxifuEGbPwok
1COINf/pGCFY7i5JFBv8wvan9yerc+HGlpD+opGCX/rUWPHmpIhScwcJ518wjvyi
pudPK+SzkfZmgPL5iNnNwC/KQZLpJdZ1q64H0wDGp1TVVdBID8+NB1DXPG4wlZ8E
f3zVNbODbL0nwxBsjsgzc0Z+Bs4JE/+22NHjOL1/h85giR9BORIvF0qF5PKFV1Qo
59imQY6nxDj5rgzcWUEQC2u8Zw7jsDFz5Tu8kbqv7tT2U+nYOQs1fyF51EtvF5eT
vSNkz+JFAQyYPiPyJadWGQYpWuFM/g1r37Qe9SVXs1JxF5AkbbgwY/ZS/K75L493
lf8EYvQlwa2cUSRK75dmt7WfOTqIFarEF+c84QT9aUUAZO4ynKULV+Kiq29/9b0T
+1wq8TB5wYVLPjNHrgj5BSbsV9IeCzV0qG6xKezcJvDKEDBL5sMgENGAmwAr99J4
KHX1SdG2fDlbcb5MnvZVOYLC9yEeioq+QJiCRyKNRv95u2JZNzDbkGKevRW0I/1g
eZS0dK4rkeR+nwaR1ABzYXA2ex9Wqx1R65cHibIkjPWg6HMPIvbEFFhsZpEkXEVW
4qK0HL4yNyy2xWPRG4bs6bRYcS0yL/2tLc6t7W9X4yYys2+DW2lf+E3aO9+NTO5Q
+tITh3L/bVC3HP2qnHg8T7eDj8tEg122rPx+qVt1kL5CB62OtAys2pDg3+3X3x3t
5Gne5B1t8ur1VldTqrMCAWMcYIqA5IcgBiQomu8hCt7T0WrYy+spMf40vSWy9k4+
DWXV4Frj49xeEiqbEGiCy7nxHfrGu/NEN0hdTio0eDvZVNyQIj39AMZnWYhavgSo
9pu/4BMHMEf0ocayX3hKcxFbDbUxWdOrElz5ajRAsYALMihpyyMP0KFF0kPiV55t
BYNfw2D5zd41AHAKWW4Q0hc0/LyJ4Sz1bCFfR+WAIsgDO7B7ovP1+S59mN3qp7ig
gWys8phnS1C5VHyV1HcqpPqrYcRaCSI5B2Bjq+lk6v2C4uJdGbxf028QqNswUpIi
zYKIa0vUOrFgCRCAjWOM2rPkKZ/wqmj11VDkyzclllPVXTzEYxvMEMIBQhDeg4zc
NPUXZTAQ/fGEMAWrPBCVTzCMDNC8yGeqxEYd8A3IBAARKrBeJxpKUgfXFmxNI/t8
sEvjxL5L2/Jej0Fv41P6DGST7ijAXc4hPFuDaELhGmJ7XwzLTlHz7wzhrlIL3FKQ
kSS+5ZPjsDiyRHsUcriFZvDK9ZBFRLJL0+ee7XcgemXSqRVgwT0ShTn6wCvVg6XZ
jVzb5f2rzOEEk+8ON4SozaObnq6FKRQ+xhWK/acpKlrYg4+tPk1XxO59uqhPC29e
KgAlw/PSB8oSrpGTjZXXFMWyV3pQ74eUFeyS2Kuw6m7dedq4evqQNodprWuCdBuL
uv1G0IfaFv7zha+tlnChW3IjCRhi1AFjlEuwh3eExRTQ4mMwTRtLn1WNupZ6CHGm
6c7LaGHvR0j3ario8go0+V3rNyg7zv7xIk7NI2gEFxI1Cgeq81N4+N+APwzMXgWa
5yY8uh4MDhYfZay9aRdmWgvTWLt0P/xsajBvdUwvdz9oWrO4u4hEEyzensWRpEHM
cs04ulpY2IW7x5SihcrV4LPHPl35kUNQDYapcayhMB7rCn95JcN+2i8bhj0KVk2c
1Ze64rUYtTjsBHb7VcEdDzkN23OrcLz644+DVR6gwpVeDdxO/uKJAUDFQhS9IwD0
vZXTrJAoDVPq0zbqsVTh2NhtBx+PKhMol1wGQdvjQQynd2dgXKv/ek7tuobs9rl8
hLYmJVr3R4tajpUFwN1vkG08u+D6XFXjQNCzNrXeY4GRUpLy5hsCghQrRPkUEtOF
z70TRPZXOV4cgvcBH0TAkMLvvifNaaqqwGccf8u1D7IxqREs5mChJN6Acz/84xun
8iTe/XMj2xpsGX8hJfhARg6AZtYy5Ri7cPK7oK8zJSHfi0q2FlMKupeFFabqzooU
nwuDT6deiV91ps9VqY9/LU7C1T6L1k7hhdeiCs1wz7hilB8ImhMvxJxya9VnFstS
Rmjepnzx6tzsO2jdFiy4RNoiCUhCSIv9Bic0QFtz8zwEEK+AFVdDAfPMbOoKfrjh
AESVqBC9KdYKYN4UdPBdWS2AmJz+qK8vbG7iRTs0RvyFwhySU8uBZwfIWQy8+wwL
pCzZ9jTwbqdPB1aeZZH0nUnzwzBFID8NNRCeDCDLzejhbgqgA/nyoz78nqhlMh5y
vJvaGRFqB3dkPmz6x7d8/me0rvn7wbPe3cTwvxscvohlJo1AYhVC6JwQ0ihKCK8D
EgnKZOHTUzR77s4sN+Mv3qEuhySc2fTIlWlQo8TVHMZK9/q3V5vsJKKNTZGFTMIS
4F4+J4wgkil13mqhVdx+qFFm68f43utfHdV8BVHXgLxifnIh/jAHGjYAtBHZ8x7F
98chSUwKlCt/l2NwN9WSt4o3yNICwT5DsmqtweeobcDhskOzYWwODPSEfRTTdsuo
geLgw+4f3POiXYJJoDkJ0XOC+jYl4kWMZbK+ItRUS34pjzRnaygHGvwUDpig091B
vMYvY+kbB263/HMAYlX04NMDmMZCy0R1/zPBo98DeT/43I294yhDHi5hUSzYRqDT
7y7GYDEgi6l+bSreg9Uhx0OnoZ25k0fYu86fBJuEjFMsm+lnw/xHSGezoeKr5yJx
qPHeSa23gTUTE/OuC3iSkRSmhEr4AZ7veqM+q/mvFYhAyi3B8LxNFNd7smb1Upof
1cl/Ph5V/Z1zs9bhnZ+WECZ99X7210gvxcfjIITf+yNTyIXyPIKakUE5ROzJU2bl
U+2/raGMxl9IJDe/Ms5GWygnhFebNQYYRt3MCXftdJVqG4XyCQm14SFiyOUf5QNC
OlLeR/ivFxy/nRZTaJMXd7rhWfYQsxdfAOw4SJ7SFDhngZufF9LoGLI6KkFRHbbF
Z8pWR+Qatak0BoNwl5Tw30yDxnEf90LnxtX4uN7eqiOEZo4IV1V5jF5D4DLdg71n
Jmtmh2Bpzc8fLN+7Yc7CKrdZjD3/Tg5+MigrPT/BdPjrqxdK6qKjUFB6RkKPMnTx
JshTYGkeHlgW/XWJ8j3lywSD49KNBY1KBK9ZzG3BUU6lfo7Hs6Dmq2OvRy/jH+DA
mlDNzTWBNUkxtnwfBE1csSOQqpZgXxN05kTLRPtuzLOV3pMLKYgJmMe4+fpXN9IK
MnP/Sx8UtkvTJYzR2rrDJc1OS0YX3xoZ4cJS8ke+FVObt120/uGYdqveUBAmOlGZ
rTU2qVm26WEl2D4WZT7vruKDEbGjcFRFSYkJM7rq9LUaicfS4zmYh0jD/JAaT4xh
boOqqhWeH3XyN5fuA5SvEPxvVvRv2Kn4b4O/s1IacI5Yb2Hey4O+AEUVJQr0bwMK
WdYcEAuztoh4pqyM0NuYXAYeW3Sa5rkI0XIlD+TWG5ZxbNk4tzp9mW0NDT5j3Euu
m982TDKrv7x5R03S6RUWm85nexRiZB6ou0gqAse5IU3N1oCgYNjxF3g40+JS31Y5
GD0p+5Kq2bdwrTA5ZI3YjzJJ30d+QA0LLun7k6SrZIenwX/tJxNQJCeMF41LGzDJ
tugH+fRgqqCN+OHkcpaTe0QhnAByejsauSv0tP2xuPJcpa2zwEZEGIJD2QG9Hgks
qB4yRJ1GcB7Zd+68mDHHM0empvvdVImefPUgfI1EL7W8VhmkhL6GSnv5AxjrlzNt
msYp29oEfQ+iazezFND8qxptNklm5aAxLKv0ufQlk/f62CG9ThHBI5S8LeWY5U9X
MwkM3lA+BJdZEvGLxTnHGmPnkLBvasno9C7aETEvs6KrmwseM3xyxPsI4j3tWTEr
BK7+sEU2uIm5nr56qou/L8PfjuX31uAoff8d4rYATmEZbDoOFU9vWXoWSQcuwZxT
/85yWMC+Qz4FqOGpdYLds/lPp3YgKb49X/qW5eQC5J3RQiJSurw4MGYF7to0K4We
jea9tEk7KxbwUk2fwdBycMqzo98FhZE/nh3SRUUzGNka3icLrFYc5UYRUC1afDps
9Ri5zwVkA1VoEiBfrYkdiGnNhX1fqbcNucDYUOH0xGcQl4Ot/YozAb0XLUPiLAXt
2z8IL1aJYPl7R1mCuoNu3remwbxueLhfjHaEzX2JMr66oUJVCyTnxGEZqg49PqPs
pula24wAIGKBl1eky4+WghFTXw0zbn0XBI1q2ZhA48WCue5U/oC7wbZX+JCeYr9w
W9YuRYXqEP/4sLEZV8WYawtrMaNv5qiQyAYfpnoPzPAQ98UrWhd23X0ka5jN7zfu
frDDZzxjjxEqKc9yanBrPjJrgLZ79RQvhXCnQTaeFxRUQEhx5EDV40jvypw+YZMD
ZMig1FNlAxnEjorLEj1DbWMzcI7QswBaJS2GxdISU2mSD7si6Xnk+eUE33kCuU1w
z70RnE0AvHZD4ekJBe9jhh8VoVMXbHkmH2AM3EwNYTNWTAsd9ziEZCR8RQ41uWiO
XWqra5mxxFiWLSn/9H99cvD7G/j7LLifFtrpo5AdRZpUlrScWGFeL/76EJkU1dWb
T8wIE5TPLnOpDYfK7Xk36/kjc6KMtzskNSE206SnTQNlFOz/l8kgoR197aflZtMX
nQjziN+Iccaapxq6VShX3vFHDdIkRLaKGYli4tM9N6M0T6qVkV5OKoKIa1vw3XCX
aa7Q1MTlmbLWczB5In59TbRzwzN6lut0RqNlaueFB14gLF3NRgV2KqZchmsZLFkR
Rv6got2oXgxDT0fH/K15Kce9kKTP3VZKt1wSYz/o/zkm6faAYQbqtu38gr3K4pch
DUIm5uvcyLteOi5ZcHZ+bDXg3wPpEc0MqyBra8v89Lh5SAvs81uv+eG7Zf0uWay+
3MlX8/VNgpB49+EIW0tHVJgKjbhcGQ5lbEIDNktjDnvZt8OyG19OCw0uJyW28jcL
LzeDZZuwAiTORkMgJRIZCilr5IHjYwiQBFo37prUatgyawZ8zeHwHk8YXH6Ah1wb
PD3vNZ7xhaSSXaYK3UIrxR7svG73kGU6LwCETu07QpSZIHzDQE8WZD6X+sLRLAkx
tumHh6U2n53QLOhrP28ZRz133a129wUXWFYtWqlC38ib/qc4YfrV3PkxXUc1Jy7E
g4qdkiXCG6nyDiNtSq0aGzeHFWr2wpHdiYGSF8dqrixRzf8ymYe3s4cKHqIOHZnD
IFQ1MLZLBTuG7M+QfEAijKb9S40aSKzsLhXhCYLCDVJMsdL3K7VNquCN0n70F7J5
/29U3LhQflduyortErj4gCJ+uYidaXE3U9rbaHzO9G/ePR1+nVl3Qzt2jeMownNA
R1tVsWKfjwNnZL8q5AMwac7/7G0Px4ocvkeea1yhhCLAqdnppVC0rYidMadClBZ5
ZEw0qRnu/1Io9S1TPWBwxLjIxpRTO6qBXgPzywsu6RCeNCgLYkMtPWZ1m/XFqKku
uMQ2zeBJg4dI8YJTtJtBOa+zGhV0FHCeYrvLpKIlav7c8Nd1dfwriykADAz8Xe9U
ZZ5tJ6L9MPwL99QKf6e972AV5zQaMcjnrC96ZzbAtaJu7NzNIorXB3EDFlligIIS
T6hf3yjBsUVzrq0zVesTlZDQHxk7KfrTFPMMso4SZ1m/JL0NOOF3Nx3+x6pSo514
OJSU4WtWUBctdmo5ubJfAlsy/HcKDntYlLhcr0t4Xzz7toKf9y2Ae2yB8oD25q3n
fBjSJg+odkG+627GNIPADBxU5iVyCVqtW2byyyXuQ4g8Y2scIi0mY1WhrAHzEgPQ
0u1IxkxCxr3k/OyNqMkkQ4qjGtdj2a4qQO+HYeVtwml+YHzhNcCDzi36ATu0/L7i
jORB+qKIzb3XZI1nDlsZwVXm3yIOXXPvNpC//vwGBUJwOqT/1G8086/7W8raLB7C
jFTf6FEHm7i3LG1BV9HQhQzRsTJbNpfdNESv4GOxT4D6qOFFqs+KqwFLkEsHn3UX
cTGxXojgPK611sjKRCyoJEQw+okVcvBzAT8BDU5g4ulD5cgH4yDtxUoGYokjC8wC
5eAV9feYX94AnMSB5OCU0WgJBfgmOfNyg/umBWXWu9oBfxSMoSF0tucr2yz03Kyv
TlOCn5/uKbIGaa6k4RO+ix4YNPkolH0PR8amCHEZ//fgrrOHRBs6wG0Oweuf14Ur
S7wad9LmU2yjGMBgABYV+zP+3brQr7dSRNjngxarAYhFrEc//RwBn2treRiJ+oLq
LSCXSFbLuf+v33oNhy2Ye6fy4nBdrQrQY3tAZsnF+4tajYcmO52r/9BSdtXPe4Yk
S8qDzkKarQjKY2tdhJgFEB7TnIesjgf6urfgAvn/xyw96ke4T7edpIt+f7cz959T
p4GsiqMtF5YE2WXPCht1uj0Bq/lgncpvAQS5TlBsYShQVgOvsDaowsJe1n88jdHC
WB/PFDo8AfsDsCB/joeYyarWuNx6IY60S+SQaToDWFvWmHoVOvlPpkronrNAzYzw
9wdG0vCSPzOcmn38GLJi4Nt0Fv96nxQbeg6tFFqtg8bKlQAOXK3wGxzMZ42v51CY
oK2Ndp1STI/1Yo5yzDY+rEWoEWZr1SJKX+JJLvVqWFpU9OHfWdnCje1NLrm1u6Fk
b73CQWAr+ULLCr22J+Bikw2nYF9TRzkrEep9/sX0sLVaqQ9nC8F+DNEhDZo+rwtd
pwMJZwZ+fa1kfnKfNCZ9s5MWLJLb/hiiHOLSEeBJ7HJCM7gOXKOShxHzJexWHvIo
Lz0iYom/J7df7rX/Gx666JdqgJ439394P0OJqlHdgGwmasp5pwTCdk5Q+peNM+CQ
XDAbc7LYzSYCKuSvzkGTsdHvVlvm/wR8Il01Fysjx+c/CcocoHGgyOcg4oxsKgu2
nqbR24FPH+xkvLbzZYKVDu0fvbKMyq8VSyT0tTZ536n4lv7pjJKpdQ7PvbMghPgW
0IIRRkES68G7yVqBcHyP40KlGMKX7RCpSgb4Rnzp9kXQiz3tBebmESPwa+Ws6Phn
r5JQ/sM5lIcQSsjqAkKxQK/RPmztBo639mmwO7kFR9efcQF6MPKOAZjSqFlcse99
7/Ov1IYOoqVUQWBunVVTij073gqz0JTryTsAJVFmH3FisaL+pOpJ9BZzYOX4LY+p
1q897oLX8RoYxz+yasXjp5jXcDGDP35S7QQ4xJV6jzWIwddTA64OkxNB1yJKTVwH
Q6u9/NlHBCQDb0c52zX4AfG+Dlusk0kclJd/EOSri77lULZpp/M34fLKvOt+dj1K
cbMgZHOY7DS+63/ji+Cl4LO0wH0UToXe95pjYsFTWjHqne8qFjW9f+DgWRmSHp2r
EkY+aJMWi5ky4efw6Czx1XxGBwbyhUNqhztsUKayv5wG/B6wK+ZkjLLAc1k1zJZ4
/1EQuf4RgOskI0TTUA8YG4L2wuEVc+Yiz0EEeSZvsbDhHqmg+xZZ3CdT4+ny7Q0f
XQfE4opGCzd3nTfD4DfiM+dK0HJWHRV5rfxF+8fmrNrY6WNyrawXFKsy8rApbGgI
9L4mT/mIi2EtNbZh8uf3jkxfCC72scIBbX+uZjs4/2PG+PHeoog4Hgu6fqraZamH
hKBhxp+WcfEgBXabuHg+Le4cbYTW3N1YLCnrJhgpdWuggNtgdZvwx84gO9ugUSDO
L6gc6OBkZ2F3Dc45U3vPX/9+WsP21nVI5g5Tdn34a6hRInfWLy9uc0ZW+MMrd+Yf
7TSbjiTLqqG0+rSFBJhZ4C4P5RpCtGCP82Y9U/gvF6pjA7Kx5O9QmUewSpXl3a8F
FK7RAz/8MPdHMq7A9uGhr0K8itg5TK30YgMJPAgg+uIpwH5tbwwzvSRlgu10mOPW
37msdJVINC0lRsGnawbHXJb6FePpPKflyQqILkih/i44+xsDPv6AjQXU7rZ8B4fm
6dCoG34GPa9OxDXnO+upVEI4FsdP0y1dltwWM7Rdj/j0xOg3u689c+aJ4ZjmEUQd
ArQgZ6b+7K02SWUDdPuRQ/lRroUr3Ejd2zsIzQOp9Loq9E67TQnbY2AHC1GVPoxd
UvrecEo2CLSo7yx43po5IScPFCAMzRkQrxS0Qp+jsZAa/miwyXKkRb/5z+US5CuB
B6jcfecU7D0p7sfeeiIu4KtLJ0uwShoBVmJYQG+cUi6YAjn1icZVKo88Uu5cXNAY
4bCIRiels5ib68C83QCy97S8cwzQThbua732Xouszy78YxHukhNvL9/G08yPtbhA
8Q3FWruCHzPjpYqyiPa8psY0lmFBJGXKM/aLTUSY+MO3WqlgyHuIl72JGrPUKwdt
eg1TMQOgYCybdl6RsnIVZC/WKNUFx2LvH9tfxkjWuthvDgvUQVdEh5Jhbs02aPVz
qYMMJFTkK5SPqmDl82AqHtwrVnp1m/IiyDfCLutJhaUwi3j2JHGSBz3rN6NCmmfe
RI0lCy3gs+G081DNs9cJwDd8bVyDemh6uEwIzHuq2FfQG4wfyVhsSDX+OpoFFIKn
k7apJse1CcZwplcK2ixjRz9kc5V9KY+WqveqzklCGb4T6jlIJdmdxW4sW6FQ6X2r
WUlKYeley7vaPEfJBRZlqtjBd/P2OKkWi78bMRKmn/ala2cbn2wzxzHo+CpXBHXz
beqiSGPfy82DhJ6nd1a39VmBIJiQ+vwmtGvidTKk0JqUtEsZvvzTHW9O7r39XMoM
dasK52dFdtW5TFw0sP6D06Wzq7QlzXVGXIAB9kpOTNJD3a31gJJFGzS8zYBM6qdr
Csq9U0x3VPXKc1crBbmbto5tB+iXjIyNo2Ko0PGMtSPdg6LfzhZizYF7rei2XSJP
j0pNHhbe8UuljZBNURLgPQ30GWJu1AvAbOAD+kYYlJeGKtMzyWxsMyOebQCnJzIU
E0qbkDrLG80cvtW7B0aMu5wysVIDw1UJUIFLdS6OpRZt+W1Eu+wv1kEY7dUwx58x
Jza85R/FrmB0XjSSxFVGuVWlOsp0dbZMkrKBuSKIuRcBRuo2yednZkcMD0q5+dbq
5T95bOcYWrHk7LpbcvTrajzF4K6vffN/5BZCdHDSpaQjAskl6b4iNeB0vH3TOL1v
ijskzKn2OiWIxjBaSZCcV2wWFJYkBoYvmN5QLcivVusJqu1446l48kYAMQD5OZq1
63EFmx5OXQ/G/MuYq3Nx1RM1EF0vEMwTeFNwxo1E6dWVpzZIhTovxP4T5U5Boi3q
rsEA6E249kTjRejH3IG5+IggoStSZol1GmOlmYKDp/gh7cc+l3AZ0xVG5JJahZNn
yXNBuSlvgYzCBDwWPjqAJXhVSm9pMtNnw3s4hvMDmS5Vm+xmv4E5272TS1S/b3uw
t1R0EZyl+3FX2J5iEOOnZtbIwYL5jOYqPdSjsjEKKW63/B10006NaNliDW6QcQvK
J10QI4bm9hxbgfznBvACfJ4kj86wc8zPwoHHjWoyt/qUAOSBmXmp4o3aCBf5K7A8
IQAZTfuCEiFzNuQbz8TwEwrFx3qt9QoYC4cvQq83ea0wx6g4FyqcBL9KWu1WFqNv
sx4156g1tb3uXVgHGGIktInAEHHbBrLSiwBlqdtGbjH6Owm0iZiddqKLd6mo1W8E
yNIL7V/5GKTBnnfRbQbqs34WLU+7oWoa4F8WqS14VKRrOulAB57iYbD2H2kAmztw
A9dzXa3ilP0GG07dKMLAdU9UB41+0BPs/t1lcl+J7OmXzErk7+KR4kGYKc3hniqj
YGTu2I41fARVuT7O6RoNn8X0LzxMmnz5e8ZjVW6/C2pQf2W6Zlya2fSBxNPdOdj5
kwlhII3NPnE2trgsADrwgCNOWTmDEHrgK8lPwJlrNJ4uLJBWmvGByZeI/YPAml+d
/QIWE7GNoTSvCBQWqTWIqxMU4YvpnhgaZQ9Hpci6O76hW9ldO7TnWBTYpG5XtA8+
tRTjMNRrXSrVIIcMKysp7IQwig0FQLh1cZiE7MP5HrndVzQFfG4apQIfsMYxQVLc
rrOxcX/Mpj/UwXYCSe3ULBy0je5xq5ZSG68KKlPNekjPfBdR5VRd+Uw5USjI3pW7
q7W+iVCdDu0cWSJqN+CDICp9P3MRhOS2sxD0SI9Co8HLfyJ/I3zcdGVYjf3RBEdV
g/zDu8oHMNCWV3ZLV79Gp95slyVYa4zB3+m777aeTsOUBO0l21QNPpZ/QYqDWMT3
CQVVwEoCKSOpshMs8CurVnP5KT6HS0R8SkAyE+0z3AYAIhXpWti/MDn3sXYI8Ii7
qMm0uuAgMjxJgS8AkgHpL1zunqgzDr7ojtI3W10yapeY6jtmn3TqEFxoTCQyIVOJ
RUHOPaR73bYPnMcnRtpMhym8OaAiHpxj6ts0AV3PQFEV9XGmgXtPzLWXNdxEvVkz
Oi4eK2GeYnUENnqhEmtbTuoJoKes9u4gNM8Ds9Q9gs8PnH+eO2XuZ+Ea2T3FwaXf
1f7fWTq2BmKybUtGYq5cx2z+jWdXK0K/KZ6zyRkXK0zT7Y613+I6Q4/iR+SnGY2r
3zx56OiK9/XiXSFS7X3tRSACe4+QRTSVTTN3Iv1+/bkfPrI69scqo7zRd3tn0+Uk
oScxYZuLmCY/muYJQEeFqJegAiHuEOxPSN5Ssntkw9BI1kWxJ+yCDL1WofleAw1h
8HHQBtUZm69j5/MOl47aboFqYOHqc/HKuVvnKaDw+qTcWWm4Oc3N/0PHaMUQ8fm7
WpWQX0J3KYz8dAds+p0zOBSipqofNR5bbrErdxMKIuzLkdKWVxS+EBIh654OB90t
yh1S5UsRLo87Vl+9KZkqqpCJAsnQ/6yZ+ssxpNeJTH0vcVES4AvkUN0I7HP6ziju
MfWk3camco8gk+pDVt/ZcU4TUnADkxWYhE/xBA8zWzPAC+rd25FrO2sG71JmfNY3
UtMpYKDmiawhJxzY3muce9NNjG/kDg1Nnz6H1wmPBCoB8GdZ2QexkIX8mdmysTig
ZR8DPRmBzVD53DNS9rTrc2wQOTx4Yd1LTZ+B3qq2pZPsG0SK2rkD2KU121LrEM4R
nZ/HKB0Ua0gSk3B/N6ZqvW9S9gHAxhcnhx1y4kRmmjiWPNi2ZMXTKVtBMNMcm13U
oQcSaifC4EyHyYbQHCzaGfAEbkYdXeRFIOLr5yPxbaJ7BghaUVN5b1Ktp/4tkKnJ
F+m3WSf78kt8R/Zyd7fT2nbjtqC/lwvIE/2HZI8levAWvKEAghzvvCsV3TXp/o7C
+SUyAhXx7WdQR/lt27fVoLpZy6I2ihB+ZySQlFbgiyP2vbev27CDFzvJjadoWO0M
FZNxcMkSUgbP05OiBuqTk4LzQrjtO9j1aNkkPF2L8qAyiMvp+QhpCuBAj9lNLpwq
lL+FmifSJLlKS7tqIQdJQysiU2myCOFUHZBVQmDsTVS8FSuPpVlZu/aEo+vQablg
2IImZhkwI00nea0tIpeBfeCTT66/RZKuk6eWCJfPtCA4LP59L7V/hC4bnW4A9UPs
hCleVU7dXLMFsymNgsI/L6+QURmWZnKZ3wcCooUB6QqYvleC1gih7Id4l3EwF1V/
5mMuqUseFwbEjny4DVS2Y5VPgyw3Bm8X4wq8nEfSrzPMqygth/MZRY/zu4zPlLgW
KPzYICdLK0S3mEu6Jprpjlmc0Nj0rJsDsL20hfI+dPXaR8hZmlj6nUtcsRv15IIW
R0SeHkeVr/7Bd8QcQfdNLkoigAocgd2DpYibwkFsqPzshlqTkkO5dsnaOaeTQbiM
pVUMbHxj47+YIZ53V7fOd0d2e6II57LI1UTtdoLUgVqnFj5S6I++L55wjYhYd+iA
sDZKVQrrP7bCOJ7TTOQhPohVUVIbLhp/jV8QIAU6uN6wYQFeX7oZVTJKNbBrGl2v
qzTUXBZ3bUg+fNAwv4RxkvOwYZVFvw+jIdL7H4TJ9OC6Wc1l3OJFPAzPC47hdPvy
oIebjXkmbxwkMMOg8Oy5ybs4P31iDp6CixNlrehlQt5HWwFpH7QjOb6vmYUeVoFg
xGC9cJsdjJKhVMG6Qt5KtdjZqy44jz/YM3h4Wulx0tXpoCa6P4ZZoHk4UTFijlIN
yDFUvIRNw4CjsWG99+VcPGxGbNfBUX6wx0zKNGZFCDQs3TjkgfAf+B2RkXKcbJLi
/vbsqUxvMqGGLquOA1rsAB24I/TkCc8rG1aKB/Nf3D8HTHo8QxVOlqbuq0Esoe2H
6X7xO69NuAxF6WOftdG/kjPPDxIXspUug4aWY73JaF8hkroAS7h0YP8tmcXHQAT1
vSXYjZTiEC+gnOr/KDGcMdM92Casc6lss39lQHIQPj1tirGNnsoQPVFR6oiZE1sw
txer6Zkt0IY8PN5Pu5TFsI92LYAz+2Ra/7FqhntcvS9RlbXEr3wqx7Dps7eQ80NT
0WdyVNUYfXpa6yuOwIRz7lR+4NDEI55z2RteTQuYrl0KIm3BHbdX3ivDtdmypS9g
QgBFxzGTiwig0LTpXMhhLFusyqslAHpFc5CX8VrAZPjjX0oaJDEujef/3ET17MlT
LVxccm7IEmKFCX0cBuCTZ5kUl/oDBq33ahQ69jGLRgbrRn1wORQno910IOfDM5rr
I5pEvo4fzkGdJmkv1UgeqpB5cBnWnxSPaXhJVZi9V1q8Id9ZO62Ib0O/sNoyCluZ
hmdDq5IhClMVKoZsGQsZCd31V7mjjUYRA6sM6NARgUqZFvOATioTDjUzS15TTan6
A7vbZVEnvhyle7kHXx2CwrPuPPuSfP/6lL2nKFoRgYQ8UEVM6+ApiaaVR7x5su07
GTtvIh2iSbY7kesTW9FjiC+tMvNP72bhJpy3e/aRq+7ewA9ifgj3O4Gy9IQ06MQD
y6CISknvyHFCR2UdZ4ejSR+8OrBqzpDP0/NIZmL2N723gfL2gZQOjFDX3BAgnwIb
vGe2ZxrEz5+zyx5mNf6eAgPXlhUtOjFNVZQ8l/vp4zdT0VSiSzOnS1n79wC68QpM
tO4mJAl2yWtk/kTJsWCtAoZfzl1HgwscPtXchCC6+whGW+W5n0p7VuY/NI+8JhdB
nUmpeVya2wFWnZIya+RMeiLqUubIWWXjp6/hb4V4/osE1jQPlqMj5BvFWwagOojC
l6fvr8mSHYKUeUJFP0nFO4uYAQQVkbyDn7eDaZJOr6+4B+Nlap7C1yFHhH/+z7Ur
45UNzM6MuEN2b33FxoZIINLjcxsVQH+ZCH7RNC4DZ7byQ6xQmVbu8XUUmmWBBaEB
D1YSt0wSG5TifydoIxQhfj2FKLyLBnsosfzjb3B8NLpEw5ASJAQh9m4Ck7WNcE8h
j1ikgUkrJ4SAf2cwRE182zFlhs02VvK+J/GWeS53+p3cGS04tMinjYa7oYOiDFZQ
FMwZhrGzSdJTb27iPooNo0bDQqADMrz2qpT5r0NpKO8a6FZMJOZbHmjWFI36sZFX
e/O/UEyusNl/a0mdAzkk3pR0CZSdLvX9MsotjYy9wDYCV327oVMb10ocwCrWkaS5
FUvKgIx3TOAEkLUsmsbwrFO15elGIeVeGufQCryvUD1pl4LKsvVkGvcqBBS3zdDy
ej0gIZg5rhOC6ItUggNxmIkzdYLbqQILMpgW3CBJo31MCXxScR6XqfFry8yQwXfY
YuKyGYhLlCm8WLHgzFQf+Y2D4d3SdGETx8fsTPgBOcL4wLZ4wdz/ahyTw5kCLiUe
0bqAo7sG/GGBAcSMFRkZrWABGU8lcDC9+3XIeWSI2XBK0GBB5Cq2omCKFCYLEneW
QJNG8s4SVhdUQ9+02PJe9Jl9UqPd3aGwbTh3fyMpEFuZg2NR0Pr2Q5+ThuJObbaU
GhT394Ze92cyS/S8SaCNRCWRxlGaINhxZjjM3BVky2TMZlATgQ4KxAbWmlA5LDwa
7WP7NMKcRLO64cuarNna2IvHeTTuYV8ohDq/vfml7zPh961yC+R2iFDBnV/2jMl6
eveJQz9DolTkxguoOh79pZueO6iVCUU+/QTJQBqAvreQp9Fw3/BGR3ntgkjhl78C
gkM0XX94mYB90n0TMtrNJtOLhFoMfdtQh5sPlYWewjb0wJd/SxHT2PdboOs4V18h
PWAC41+T/VY2uTVj0USVKz2aioUxyriPAJoRPfTUTZYK0oQXWoLe9VrbCSwadgf7
Iw2x+Pv7zre5/tURajIEawMMaK9c9CkU9fg5GLO1BA4hI0APoPCb0NIcd7XWA/Y8
QCXlc2GT7b+JjfS/Dfxpu5JMQ+C6iaTSqIjtwFjYmoA0umgJo9diBll5KZV97jdb
Z2w26mfzl83SJuFtkk0fY6PgtwunOaB2aNOhhIUcvpT8OnMmD8bWQr7lpGwdIXmZ
TYwhuSUEWYf28NaRAQ2GL5C24f2RMsVqRdom75K8/5SYh442fx8RBtZwxkS3l8ku
2PHuZ77t2FEaATn92Bq5/1b0hJsbSylpGL0CNjPdrrLH10pcWvT/kqoSbIObTw9X
GVhMyzAgreJDYeZ9pGU8LJMmHLrEOL51iWk+2XtZSI7nV4z0ufIgH0ttJswkqLB6
GylfhxA8nUV9mBBfAwkGF/Ok2VM56uclgMLmA540os2fS6kpbbKWWZVpLwU7a2gA
ZDcedDavpgpatxZft3KqLwfoqH3iy+rnQT0RBsMiQm9o7I5rRgadLhd/QLmxj0Oy
WaoA4ndlBnyPdhLPaed8hZs/t2u9LPfFVb0ixNdJ+qh6mXvPKIxCjmUnYxNUelQR
pXrNE5U5h7ypqm7VYmweP2Q2XjaWTlxxk38qfjnI9S8Y8SXgkWzt7+ZOmo+RwAvd
4fNWvfBqpejSGc6IG1nqYWH/bZhyYzD/iXP39f1c/eW31HE5bg79UzdSiepefJVZ
3zRz9rcicMZQL8q40vWuW1/w9yx/gMqr2j1N9eqnOUjRbJzhSMejrlK0PzFqeQNW
avhSrF7Ky9r6fz3C0sa941qgXzXDZAwDBHPLhNZfJQD8FBSu6ynMJGXmNICwGMNQ
QAZx/68OodIUEOSjtbXrMFUq+PuosR1K6ADB4ohjpHH/AxaMCKsY+ZFsPYqCiifp
mPbViqHFbDijw22UXoccUIW8HtHQxay5B6KbgfndlsTqTh7A8mfcLu6ffe/Q9oKi
FRVAdc3yla5zjLVOEyhoU6HTD+dSTk8Ax169Sse8/vyqMsZSRnrEMOjDgIkGT+TB
B+DTNDUW38J1ymCbvzYSKJFPBXbzO5S9Kj1QEIhNCwqjPdYlK/rcj4hKHOUMqg1q
hb2zJu+XMxZfaNAgVb/jgbBxed52ksb8KW8dFepWo2sbXEd0OE4fzEplseTNwKs/
K3GmS53GvCvbUBPfo18LiYiC3sknf5GOCRHV82hHFal497ArXgys5XMWTwQ3MhFu
QYYLg7ThzmNMO4kC9/GmAHN9KgbiuBVYngPkHmJE3lJC2cS8CpoaGptw/uEvMKIT
NzwUw9sGdfOvxc2aPyZaEoN2wVWsmoGhQKGXeOB/eXYTdogz2+pvvMgMrRxGQCyH
1xnxnj+hH+JvLqiE2B4F6UXonG9MdJgAT5srOrpDU9DNEvF1EPdziZBlqCzOADDB
x/ISdkooDfLLwB3nbgtHrJI3E1TugTsBTzce8g5X+eH7QQsLIwpd62DlN5DnuUaj
xYPLBTUYGJLKAFvshDN5/glW3ffGxPuzD5VxaK7WNbAx3OoMKnjWq4SKr4nzbaBG
9cRU7l1ETuF/qp5jKTep9HnWZCL3kN/A3EbJJa+93Kl53CPKUUtjQyHS57KP4QwI
UuAg5wzZahi5vyHdFm03q6UzlS2d0LIBbzSbcOVY4hZ36UXSFw8Z1PARSP3LuxBx
+4r4gpkfadx48hlxMp4PVYoiWHa3dH7x+5YZ1ou982KIt61KnTZ74QqS7owSTGoq
QO1/8OBSgyvlDD5UdxtvhfpG5QcVvTX/nDYWlDuiwW2ui0uc3/slgcs/bcuX9nYV
Y/9G9j602aNz8wpwMZfJ/XXjisdSY4mQcXdxDPNboXfHCNl9dfQD/ZimtzqpTQlb
Mmr9v+AzFBM+jOWmUWhwMeqUXS+BTqlwV/SJqcI2Im/gK45pk+0i4B498FCuGTxD
BBEs4q2DC6jHXOTta6VWTPZ+1scaxkKmyyd5hF6yBD8nRsI/o4ki1F1hnnbt1AW+
ZOWr11jBYxbJ8kfcgT9sfVbKfYa4h3E+ivKDKmbIW17HTmgoGs1Bt9EPps0lgDtq
qE33j8mK1p3GfpVEW41HbgOq8FPzJRhBw2MK5MkcZvRyJ+Nd9ULRUQbojVRHIxEY
unyxZ6wEsu9XIs9DGFSxbGn+uEFbTh/XF5Qrlfh7L9pqlU+DUgvLg5DlN9/bE4iH
JfypNO6djtBBBAyNJLBEFL0KE0JQCPexpo8PDXMF45dRCAfgddSbOYrMxfBOBTFz
y36ssWO0rQh4V3C8CzoZq8vKWOzJ7OTn0SDo7ZpzMb4LYsEQ3aTw1DrV3TtABimq
JEGAOfPbxR7FFCKbCQ4aEyh6nrhzg5FUGREKIOqWBjQzeXX12wTv6jFU/0Ijsx3B
fuTu5K956WqmPm8Tw3kpXTw8HLChwg9cpqG2qNwu49p04PgjAPGPaDVPbDzH4Fys
GjaWtroCX4M2m4IMrEScl6RYshSr2s5Vg6Ve/bAMNrSW9FSypdRJbk68F3PlNmNk
+unPQLocBsuoQ4LgZKjcqCl7Hh+JandjqOGk3wkcnpe/3XfeKVbVWmVACq7HvgAx
fkQxVYtF6UOVW40VSHytccXgFTR6+/wI+duQmVyAznEuq6Vb5uEjKR0Aco0ycq/+
gdYhbxCB4EJfbkS8xcvPgqZ9m9MBOKKIyaqbwY+tD4nfxiM5olGYk/uyILgkSONZ
bJTy8LbC1VuW9G0J8usFbPRc8KKd+T/0xOwylosAOX3ZfPbyioxhQoIBBsFkXE8c
Br6Itsq9J82Ttqww9skZLQ9p/3wd/RoIlZblUh8IFqWMDCY8jkAMUJ4FSRDFFDIa
aWdBFDrhVg2v8e575Mlq2lRhI6qED/idlsKQoOu3fh+twDNkPDIve5DsHJl1t1On
YXSmcAyVJx5a7FGRUMjT3oPYy9toid+GrrvpwfNAL1QAiYZE4/VfTDo1FT6gbGT+
2eaG8My6jh+cPfDZi9/YaOAANE0JcSH45flvjrxhu1dQN0yqioChfQ6nPIpLYLjh
3+4T3JM7xYoMJWSXzH/XfRAH1smKRbfENRJ+aNuHVwuPlWDJCLaZNIBAh1Ir4GYJ
fM+L/ODBz5+i8CH1rUzpi/jFYCW0Uk2OFOISpihRp7CftxGH1REeF5oLSdXV4G8g
6E/YEILcK/PuYXYo4l51dGxXeuGbKlPrkjBIxfvSrqArosmgoVS0QnxFrvL9oxdZ
B/8+h9V82QIl+qjEJpx3B48f8N4Bg9C0cpEdJnJkFT1x+SAZW83blsN6e80yRdTz
g4+VV7lYrtqeYfdlEk5Bk2MuV1343coulyFS2XhCEZ6ep1pXe8h0h3fAe8Je+re/
TzDpqCYnlF8u7V8WjhZ+nbT9/P0UBb7IdQOPMIH3cyVKYgKheFUlD68aaq9rUHFb
/Zur0uIN0rnqk7VCcqC7aNCYsM2TxP7VXgS07fZquilQENgolFXav23Q7TJ1m6SD
p9SayKo1LX2H0gasL+gJt5ksq3eEgRL3yEhAal3NhDSPzhmts/GQJrvoLOgIzGyq
4ustB1aqr87XObTdNbq0okQFi0JQbvgavfkC7Xdbs2yVPxFLlJCPWz9rXF3BtY5R
FvZdBAyD9oXiqxqFoUUZ3tEcgFuxot0lKMkgi9ShO12jF1hpygzUtc94EV9ASIZw
N5bnyj7asvFLl8O5sfk87O6w306tL/bffrFS9oIOgtzjl/48Z52062MV1DZaFVo2
e+jJxtjX9Iw8QP86FxGnC+ovc4LBV1+J1MLNxXO35vl9JJMEvAFnMWuN+CZzVgc6
grm5//EcYihdkcfR6QU6HgV1CELtuAv/4g+oy+WF5n5dE5ZpMwvHN6RY9K8ZhgEQ
AFDfM7m9wpTZIkh9Sa54xcyYHZvtdt93plpXXg0tUCwU+uOtoNbjJJ7Os69UKxjz
UhlfucYuynfe5JvtIutoITHRqVTw3n+e4YFyaDLIjkBL7b1YVZX6njrqkogqW8t9
WdOxIoWu412z1x5K5BlVB+jt92mpNPWvn3Sll7JXhw7aBgkiDz5HaLzefZlNDk32
VWe2fa+6sKmiKti5U/35OBXZc+n7OndH26k2MNb5y1QIYWcfscaplapkM72YiC6V
s2tokP8AQMGL22JIRAfVRbDHqo7jTn0IL5YKmzm24rKxo4rNnNmUeJcCW33lEbv6
OEu3O6mOsHzS1AK3RZd9apFy7KEPQw6OqAa/IWyZBa9roq90/goAIubf/TG8Btmi
R3TL7rZ0fU3jbPlz6U0WHnhqbBnBtTgVmUkKGurMLNXAzdh3buo8cxW4VXyi6oyJ
/LNLopVonEN87CMb1Jf77bOxTrKM1mWJYCXkRVlDquZGxqPIdm1TyruebaB33X4/
KVo+YZ8nG5OQJM/aU53X2BGqzpCEPOV5MuTcZr4YZTolxe940Czp54RO2hSmLxql
owBqY6g6TdVp4XOdyG4FgDlHOhFVFO82nTJBJSBaRoID3Hq1r0PNcFK2xKymvFKS
tt3vhLH+s98CZeEJxw943yCa+R6Vd7mBXXFoi4LDc0vxH0pZgAt8gKGbi+Kql8zc
4Q1nmB/cYYnCHXj979x2tgcUmB9WJvMQhSR7t2vo+bIiRSwsILHo3eFmhXeFycCh
HDt1Flv+g93/+u+3dybJnFaeY/3clEr3N+UjFY6G46B2bmy+D7uZAF9ZcXXfMUiQ
hS9THjVaQYVq3qmohG06ur4h3TXQtzqE2trgqjTvgFx7TfynazNWwZYpYpNCVSq0
ZvpuuTzTX2VHpDPj2b5xZ61+2K3qnN8UO6kbFc9I+cZ1sWkFuyVs3bKJcC8bt8Vy
kbYZ3fEwSjCaP26T1PGopJg4vPn7vVFkpEFzBt6phgKwkSNTgHRpzHDx95Q5crZV
BUzP/IuKB11bAMfK7yAmfwrD0RbMiiw6Clghv0o4jGsWUxmK9rP2ZiPdCbl4Z5TT
Cp6EqhO6vmEvnSKSVIgi97dXKOJzLrY7iHbzkSKiNCy2VirbovSmMwMQgXnuhWXD
CmONGCOysq6JYKbZ6aCdFAepLS0WOIzPKxrl8EgZkVmPZAj4aqvslxkuHYOuhNA8
LmiJR1m1JKg0oZEe74BB0U/Zt0BXdZjyc3bnFUy2t7o7GBmctT2zPPldeKtEsntC
YgSnPodzhlaPWoSiwuz6IREbmhassPkE7pbMUCR7cGP6i2JfnlEgmwv9Nu69+Z+F
I61etCMI0Zwvfqldk79Px8DTagO7MkKy2QWnmdbDxRjdBxMctoIlI8ZS/huRdjBO
Msnx/T7ayrQ5jGKkjkz7BymcSAKiEz9O0SZqhj51ORvlepXOwdD5BIK8GSU82+mp
mr1qtnM9xA+19WLCBQ5kV6A2/jB1hGge23VRHUn0IFs2Oext1H46pPgFRYWrAIpK
uJertBbyPwIXLwn9tuDeijqfF4Zk6rIRyBtejB8tOSCjluKTI+fdgrU2RgNpyLbX
RjQDmGVMtyWFkiSfi1pEd507u8umdE2SjqmGdsXJav3Ay8po0m9ycN39ktt7pY44
NBjjGlI/rLryllDSa0ivBhm2Rwg7BiYbvH2O+zhQsaKMMt2aHg0hkwIOMADI+KuF
+ahkmXMecDhhxzVh4EDV9K3gsw1bEEaOC48r5PPsS3tuu52FXp/z+JZWqWxJEOjL
Hv/A18aFj61ItBms146y1qwRmPrax2TFXdn72Squ2bQnquXtDHkvP3jv+h73TrPF
9qdBDmq9R9NJeqzcruP5lA5wV+NZ3U25ErpbGO05Z/Mvd6ZnUsACOU9Nl+/PDiui
hc2hjoeJs6kIMD1xzT0HT74aU0IY169oTuATt/Gve5t1OZ85z1ZyHs+13qMQBrZm
V0ixJkwRWdd50+/aCmCLevhlCNt54zST9j90ts1yeEwg1EgYFhTxVd0HJftifmxS
JOKa4V53lLRdBqFel1g6pr9Njg10O87S9mgu0XM6uLpXtllD0QyLG/IYh6ettHvm
O5c8sKXF77QPC99A0JRh5R75QzhSeQYHQzGP4ACFbMv1VOCXpA0jLNfUFtKYZWXZ
yXIgTlV6zNFN6kSGkyKLIQo5+EyNQyfAgGbUVkzV/AvKV9M+7z7b5uwcs5yP/pYM
nEvlhxZ9vkS09BYrCEHG0pEFI1lxeCotdexza9wIdlyihlGpaI4jJWefn/JyfZmt
S/AdA+kMtiBg+R2gFXqV+NFAgY81Txi/+IWiQNmmqAZXyTgRIMePudBbwQV8g9+u
VIr8dSMbOCIibGxQV60jTld5QmDI4FMJZ/NxvnFUNcqU4hzQJw+S1M/PWXyMSblV
5UJyQYyQTFEc38kfR6F0+oXb4WE1pgCYka/hJRbX54PwyBXL7YJNdFtC9uqMEG4P
FooaKvVvkco+qB8Ea/nXXSUWRsO63DFXC5NXVeM3ZCxrPdXo/9tEJraQBkGKf4kH
SL2vFH7VT250nON/Dh4UMGgJkreD1LAt67G3yIIJ2EFdhIue/9UPtqxWiZP3NuKD
YdNKZ09FmHiin3j/SC81uLpee4TBn9ysiBg9aqhKOFM4QDx50kRwILFVkj6WDQiO
4dkeHSL1ivtXm7YZDstR7OoAqRD0BulihnuGMjmR6JHfC17iS+/dzK/G1tAORuKI
TrEP0IpWeKfrr7v5iTtRQK3GTESYyy7jXdNX7MaxUi2vGXQNHBLcGO1vYUcZDS57
YYESSq+03RxzxDBEsDCJtm1mEqPGE657PklZNBZ6nJYHUKW8t/j9EaywYjejLYAz
UTqOtVZPFAAdp956T6R039lbwuLSRqP3uLalbSJ7AEzzr8aQYD33NO4yq/czUTYl
SDANmwalWOw5RSaH2XHX5L2P2G14jlaRXR1FqW/bSjZzCCXqz438uP2xRw9Ct7dR
5gBGJrudlzqUwqyOR9T3qQpvW9xHJfq6fx8Vw9HzE0AE3JD55K5mKgkvCfjjhHqh
IV03yOMmwETHTFA+oU2QRNIj/G2qPni0vCs1MrGSyHy1xaIJC0lQAm8uuLFa0Q4L
4K1y94YG/AUzyZs2BCc/rwDjzWQ0ODl+j+/iqmEaZxu4QpV829i0dH+60HK1oR2p
F7yzQ1/2j9l4Il3jDlSoynLjOcdu6lC3bk/4cWJo1Ym6jQzCxlqsPTzoLIauhKR1
8mcZ+rsyZLufjKcBZvnQo7eIMs1AXmqN/JsOTksg/8a0G6CTrbdxp1pmUI6fACtO
ljUIVv+RaeHHTyLIK+xZuYYXXHCBGdXawB/LkoAR0XshWhQx56xMtgzN0z5rVSeY
fleDtnwXGxX+MrrrZ95v61Ha2jKEJ/eTFW6lJ6Czegrf0iPCgSg+um8m/VzGpW/D
RIdtr9ryT0PfU4gmuJVXhNown7DJTzcWZs9nfGt2EgqiWtDOJYdU2gUnSDhNLWtb
aAXR7jtpMJjUM9sCHlVdXHMysIPLnHVYX7aonXTGmLXiQ2X4uPonwLlkxfwuFS9c
LxVaUVhIPmqflTIMRUlD8SquEESwgrQXyce19nvCjNtGW3RFx/5RqM+40rO1KTu3
QAWGxdX1SAv6gElRkZfNLltH2fwrnDkkiPXY7L8quRCy4XRwcz7u6uSVmKfHVc2C
VBARGAxFjSdPLG46U3cIGwQbOMBEBvrurn+3ZBeOUcjSpDy9ZiEJ3pshUl9YRWfn
vA+ehP2LP5rzw7dT0ue1wjw3Z8/NLLNnvyLjehAl4wiSJc7mfb2UvBibao+UJrZ7
YCtgWy6dpIqRobQHaz6xUwEsQUbjtdC82qujXmiE6E9HL/TDB9jHpbLiVInV7MzQ
zbw72lW0fPYiun1d0Cl3LU0tkUsDLMKfqv1Ipew5LvpkhLpIFltdyOiYvQQ1oaI5
UrnH84RYuhQVBRotTwR6/b6Ob67Ko3AiDGxloeycUHicQ0B36pIUXSPiIjucuB9j
OF7ozil8D0hP+dRCXa4+EcxOga4WfBPiO8MtT+rKP1Wu25GthJAVd/exU3cJ7l8I
6x9yNrUIQpYVGRjkacsyiNXM09Ijt5HwOxj5mRPGQXz2ahJ03Us9LfSIIe6plxTU
dr501VtoR3aOkbiU2MY0sYDydqEuLF3xEQjI8mRZ/J5ZzKvSuKleX5sytUPaWQT3
UoPgIRmh8D5u5oOKOXtFFM56VznNSd/xKKnfqhvWjTnsMSviNw73Je9p8o7TQedM
qOlji6aT/DEmESbdT9YBXkON0MzKUW1ZyWJc1cuLWvDWpEVDNV7hVGCeipyj6oD0
Efc6eXZCUCoTGaFSmMsPdJ9bfkv6B7wR3wn0pvrgjMOwXQPmYbID7qokihrqp995
+e6Dwv4/3fC4JSj3GqEf2Dg3R6Fcj9rG4JRvfhx0xnmBfNrjjqtF8u5N7leQXDWs
tTjeWy9p/u463qJyrWUknymW4pLpHfjVrEC/ObqgDDvprEAwHirzt74h7lw3lZjx
1T8i7I0m1tUdeO0pjODC/j/nENj34LQILv0KaCCPOFgup0VHm35pO9HK92dXxwds
kj69O/cn4LugmVtQ7VKGu1zbZ+a+ZldrONS9Xx+FBaGGqpgAXDsyXucW6DQPtBJ1
8XZ/5DysNVrx1axBi2hZ8AfcTZFREWl3XOSjGEhFcQA2p9/qmuEzmrUxcB4fabzy
PTJHFGDRj63XIvWcIVbNjnw+PTuQQ98DUY7TvGVu6ujPowMZIrhPMHKwo8FhifwN
HiP4vd+lNYl1w6Az57nrJw05lHdcvmUoWydpP/Gjdig23IEhf5dYZiqH15b+zRgZ
XsF32YOXOA1mGUE5Boqo8q7BRoZAyKC/JbEKbh/kB97DQpGrTm8MOgA87GgmRZrh
ZU7D7WpMOvhU4fwIzgeH5b2Ztz6c7owkzfEzzg9faD5Babgr2t/RpzBVfjqA7HTl
Eav9BmDAfmQNKN2JZyEogvdMm2AEQ3O+jCIV0kA1s/1FKmdZJFq7Bqur4RqjOjnW
kZemqyIn+BkQYR+QrtyBFHi93Bi5gw520skESjn2+rskXDzewN3to7pewsvsHmps
J8MKywsgVh7wdfhfhyQAHDs+tyiAvQjk2TexBpTyconfWupLwnAlHaDA4PWmFzue
S9lylOQBvgLjEqjaY4+VxvqjzuX6QeKjx2kWrH/f/BLkPfATbLG75JHQD8D962sK
3eescd+0tF5K7h7VAyq9dj+I00SFUvXV9D4JioKUM2A6ksK0K8BsV/G20gNJEtCW
L/IhPI1T8PRT5I0HsCnrUHmqz8pISfQ9FmORuWN18UlUTeMhPNcZW/thtXGNJiAG
Ihr7oTZzE1AZP9W9ya4N1YZMHrBymz7VGjnwbEPjzF6KyfhFbckxX7okQjHR4Cm1
6b7/gmPEcEEba7WdltTLULr0brnUnI9yh5b9m/plU30FoST+kP6Ss8QlX0AUCHDH
GHeFoJ6Yj4ihgsPMJE9HG10tT6SFxMD/Fsi2ycZ/hsed4+DDd38q7rdnS3HpFbri
6edYBgEO2azB2/vxEGp6BEMXJgE0LtbMJFLVfAtWKtZjoWnoxBr9dQ9mwsqvO0Tb
bRP1/soADfDWGALl6DsHphi9n9ZRwmAyH/J9WYHTRUr3uzprAln27782l4iGvKbB
oQXNm7hsDTey4TKGzpAX6ouJMTPem1ZxXh9sj1l56tF+hZE8eMqh6aDhAH06k6GV
X03667DnDGPjRAX5yNN/b6uxtzT1Ywap8SyEqNSfbPJS9SnFBFyiy9pywluupdVC
C8ZEkILIODU01JnpXH5be8GhAtTTqG4RlpLczypkXK1jsPpw3REa7TwV/dhvmBGZ
dno4XCZI3m8aNFegARsQ9fvlQMztCbt70zvlXKh/oqpUMSennWReKhx3sCd2XPDl
gcM0ZXngS2toElZFffSl1VvKgKeU5RRIez4lkKcyGq3Ac2B35PkwjJvpoHR8LHjA
DSBMAXp95NPhqF+0NFuQFXSnPGzI2bgBGj3c7Rehons0Qv/nx9dcvFjudZH8uisB
vwd2XxmDMVw2tiEItcqD5Vo7rN0uPZlEmfnuKwiBGfDCIEwovTg3MSx33CsTtcZC
OqGoSkbJ9HxtqVY1lzOpxY+Ew2kWUy2gOcezrwq1viMfXcUwCRIL7SbOotgMNwIo
hGxOrct/wu+hqVSDF7m3foaXaQKOB1IS6Nz8sSaq+uoDytArqM9FRWg9SpAsPsbt
urwShdEOCeyKI3Jm7/xJCXX7kbZB7UjEFi8ap/i0Rmn/dY5Qy+2zoiVwvCZ+GpUJ
h+tcSe27yi+u8cmxE9s2gtVi+x/JEO8zAeclLejbSpngTAAV5LErBury13ZAORwQ
bWlXVM1veQ9YU39W0AUwBbxURwCJcE46GhubuEmuCzFCmlrCnpPiT8iHHOcfrQMr
LuQnjfGW8ylr7vW8LOKA2kNqDwFeUrOYfWsIxvFoaJgK3/g3gsQ/x7b4EQSwlhkk
Y1OvLR9qe5B/20Pbr+d1tBxizuzloBTkO10bLwA/rhnu/dBEyk1iSbdtELK+y+VN
argXBE4hwMpYZ4G2r8IdTc40MRoSoOWK+UtIn9rx4m34Yk8pUHRmFwyeJyGl/bb5
gZ3NUlw2A2xk/l4CiKDrk1pq0lBiX2qDEb2N7143Y2lpuAaQiTAgxEdBBEoWoqsu
/gmPU/MdqfAQoWQKIegAETFqv3Av8cXPdBTMYB+x6iIdI8PIjbsRa5mmfUINrpLV
SmypATw2pfmi9tJlbykB9flzbHWV02pWHRdKk3nabLdp6QQ0ECyJkrcfQKNwwEwv
pAVto9NsoInoQ3xCjU2TsNwezjX3gjWFJx0tLKJmHQtQ9cNv2munYQR1LjR5UgUE
iYEpz8YPdSeZs+sJFqtntpUK3HHGPBN4IKozrdk86/T91DXluLSPjEsRzH3KS5U5
oqT3TSD0LbJ1sxGIqzLJhm69LnAT1Roz7bikiofjV40BZCJj1ZOyikmsmsv2xtA7
dEsei3hClNKBfnWQelR+1RDkO310EscABK3zmDQ50ef5zX4XnCACfytDGB2owjad
1xzpoyMCwwoQqB7UE542Sy0U2sbAZU01DkouCVGIolq04WcoIyZNNS76LpNSW1XK
EoZhbF2x1wwK04tWLVdPoa0mDv5diY3SoXaNzuAG/a1vNBjUwSmoErfQpLfJgjky
Ux57c62GABaDBMLtfUCy5XMnz8XznxQPaDWqhu3lPWO/3NyVx97kHRyN+ODz/f1B
Alb2ZneWoToKwFTOj1H6BC7M8fdm639cbBH9xsBNdpGyp9vCcEVWor83t0wKpS82
CxpLXfzeyVj2k2wGcuUubHLKH67JBcCGcWzc1afO+W67tHcig1nYiNl/KlvQdghH
DfxqmV+VIe6egXyElRB54XBA0ATCDwiPi2NZwwQ4A2vhWez9vafkVSfTxilo650p
jrVYsdmnTtF1dMxjxDBI34/KyIaXgu6pmaJ4aIyKIP++6LiKr/9Wu3eaCIDBleLi
yQGfs+5MlODj+4mbnUypmDvFh8ckC+oC4//2Q/FZ4NVf30cNSYLzfxjvYPShjDTS
uGvCDPpky1hL68x/hCwQqDetAl7Z49CLGilIpFe51drjiU92usoNM93uqB5U3ZLZ
46XRYG+pQLza29epcin5CEEE6OWCUt4gQbuQ43MQCB7OX1r3fcuqparDW+hVcfX2
MEWVRkhGauiXBoQsQh67yCk4Av1XgNYUAuUgbo1XlNUq065v5/DrmDymXKC9l5Qe
SELIqUCmXIthBuZNKqR7rYmnws1qkpekzTFikgi3qzj1aE5kTUTXhuel4IE81RlH
9TZXw+nY0RzX+/A6a+Xn5DruLmSgVZ5y/wYPrO1T35nzE453lSBDIIp0lbPKtRHn
piPn8zHMYrUIT2mJXDMgB7EY26Mnsnpwe3XiRRndJuMrKVUk6QK3w8S6aTxJn/6y
r3em1rSaK5IfLyR0tVDJGJ7xHZgpdBLIDDBza+P8QuyWCcQqqb/IuY3nrob1Yi1f
hN1W50FQ/omwox8vwJbdvFEbezHgIZg6aAM5tCKWcJI3Y/Z824WW6DyRDaO2GBO2
mbPZR2Tm3nLLJqlMZaGyy73TEO/NGlza/PJsOYsroqcwQZ2C0VywVxwH1JmsxMX/
9Pc2InpKvJVbJ0g5k63rGoK1XRHgACGkZzGNf6zcjcT9mmY85TwWDvOBf5Fx4skb
trAjK/kQ69uASizvsxEOyGlVSw42v6q34etOSh46mIQFnhD5jrY9ybARXvWvntNt
reCuMAxPSFqhE9P9jiiwPxwT3X6SaU4tZ6LljGxJZdL7Xae61pQFgFWivsWLM8G9
0PFAEZ4jeFh1NHws1aRgDpsWz9kUUJCZAd9d32qDpO8Z8hKkf0YW51MKgnHcjIn8
RZY1sUvk+dBZ+73dc7JGTk5xgzPmdj1HQrW9tW6Eu7pyEg+UFSX8JE2jhpzP+jQ0
3+GNTzF7QDL5xy33L43aKUSGTpytDgbJJfjoAyObUSiR9ch+ly8D4cEo2CQLpMKb
nNnyZxbvLM6+IdoBbiGxhumNyTodz+dJL4sgY6xe9wtANJC9J42Hk9EdVbGYU6so
hEYBVowsTPHDIOsqvELsM3ykyM0OT/mmZRj30C6FsYwzWVmC90WW+mXRumpt9btD
OgR8HZ/cddvIcX39HcNRyRUQLT5EStuLFERH7XD3G4zXfRMj9OXgRp7Lac3e1sRl
j8+JbF3+6BLr3lM6XKtzSKU7Stm6akqLUqWgjPFLST3PGntZDijXb1UZ45PgOT6v
LOSI7ADbfHoVkLLW+4uSleEd1XMcDUr3y8MQEDu0gWuqWDOzUmRrlVscKBnCqc9m
ZOoV+7X687uzU5Kt6Gb9oAVlzpiJRY8zJtqBArdVm5HOwWSg/EUfnG/WU5r79c9p
zG0X2ojsCydu/hJhfLCK3E1iutvE9Diy7ZTkK0e8HzQ8mKQFekMKA/QCM4aUwmwR
BCCwgMFyzElm61C1gPYIgiVzPZhgunsO2JyeFXhZrZzvIRLrvDjpZrljhlCTWopZ
ikD04yqP/3jxsZrch1jsHZ6xk/Z3goLs8DQvcu9k2zaO+dWsd9JeAEBZas8uNpK5
ToCaenP4naVHP+s7Ua7fxQyBGseKltTUcShV2EhBa9fnhyaoVQ7QBxdxUduyK+81
opHJsouACf8P7NDuwbtuKyPlyJhxJs6IV7hSsO6P0D4a4u0pwj836CaqmsGE1pRT
FaLpyozJFaYjfBbVwp9is8FylNxb3/vZ3rmASLRoZ7XdFlM6/+ckK2AGXWJoVFcg
X6IhdKMRlj6gKHkiUfRU4LQ8xtfviIHRISmCbO6rRmmwraxzP7WMOdUc08LiysU5
/Qm9EEIAG9w3YutPX91OaQ/6GLjFGwV6zE2SuZXwqajOlSmNsSvF3D7Jq7wSk6Vs
isMPSHlC5QuJhwrlZw1sn5an1Fm+S2eZdo6Y0XpwLAARiI6H6mqSycJFwglLc3/u
SIwqehFDEb/DZjTLFKpuIkd5rljHKpDuYWf5siK6f/HTk+yd9/Y8lHiSYk4EtzgC
MH5mVC+yG1kUoreT9gXODbJYlOjXfT6QlLFzM9INLeoYymkOoL2JI0s8lHH5yTfo
abWunJ+yOEIBdYSYAusBVIPAUuzqFmNBpr19+Llz7AssCvw3aytj5KYN6al0jKVd
Z05VsDCjmH5b5RSOZCTeCTrIYwWhHRc2ugx1+qK1p36WhpV7rMtoSByqZFv6/JP1
8ugIy0pIukRxLf6oFb+f7UXL4JIrpdgLIFi2ivZtS+R4TnlsWBuwDkgaXcrRJbaA
hiF4ikBPlt84jFWvj48rdGX4TrgQ9UEX0oiQZXI2UMEs/2KB+zAWioAFXtNVkGDk
5fcSdkO/cLm2YmZAmn4txYpPq+nOgRPV552tP446d/dlr6c3BPiNQqhYVE5PyUXF
DOMDqNRGfWDdDB4DOUCzD13OY1mLWC5OZSD4kmB0rezLaFmQKZ59K5gCF0AadVIJ
9eVBo6fAjWEp1ww8vT6tnBiyD/Fe1tj228L03wjy4m6bC22Nm3omb5gmJxjdxxJB
xgai4eg4izDSKjG9hBSNZqZ3bEWzI+3XTjQWqgi8yUtFjqjiwwlioXLcZmOLQW/F
z3XF4YT0MQcU2TawWVEa+LhHrtxKmO8BKQnCBYV18paP91+3LlCYoP31BRVWBjcp
HOSPALABG+R/wE6ct7BJwQUmYYCZ2sqhL3ToTnOEcXqv02hGDJ84nFuYnm9WOtG7
CM9P8vrgO5XuCDbzBOB2m+o1l7o7Ti0zy/gQYfqZPW5weQt6xykYwMfHpmYVry+O
6argdAkockupHLWLp3bW635jhlmK339BUbxt7sGONCfhm5gbl0B0MW4tKaHHy02P
aZivksZwBXzHdHKqOP/3d337F32Hx+yZhnSts/cNhm2Xdok0WrtZNtrZnPZleX4Y
T2CnkheyIMQYb/e//NUq0LNE4aGi3S4C4+/rl65AVxmyju+FEOfGo9GAUrpE5Ir0
uCFDUO5x5rF+3XONGCingskmSz+Ut2mW3dZZ5QjhW+69O5F6QM93xwVmQpibVzV5
m/wJXI9zdgKOy5bm0g95nCrEghHAYBMcOgEfueat2iexDmZzeCz5+bVbhSmKbjip
BwFMUWwJjnemkQELBDfn4iN3aBpiSe4aFD0xVTzc8YHMOg/kvAQkDPDYWVscCGWW
U0dGCfIo1e+c9yAak0B9R58jGX4NuTM/drSZzuihD1nS8did4dkt/jx+52a6FbdT
YfDloesIsrqC8oGZhE6vDn7tXqwrrEeT78hIk2jRIzOxr4PhP6oj+DS2VrhlLU/M
0ywlctK5JaWVBEPcdszCyNb9pSCSOwD2B51vMjn+ExfD33kQCJDdOwSjfJMIl8rT
nbMgNKMfqNIcFjKUpmW+HukDmHHddM1iyMJHuO6DzFPxlOz/y932aihawcI5Et1X
WX2e4S74G70KOAEPMw2L/leB24H64lhi6QOed3aPzVqLEM0RQtt29iLK8O4Gf7Y5
yfLI+RsjjoStEbjQ9Zn8uhCjdKKITZtaO68HTY++oHgYkBCMVyX25BXULaSqeNvy
drsmZjiacKai9UmVAa3SttrmZxoH3U13mG9xNJkD5PUd/zwQkgT//RYB0B67MSW/
xR2s2z50AAWGlAol4gW0s1yDhg/3HsLjS3vy+1LGvBnyGtfzhpM7KdV9HZQsgCau
bWIE7l5CZBmb06JegiLnAdYBRhm63Bd+4H0qCvBMD5ppsgcVCDbYEdSxfFqdOpJ4
2Kkt63975CBWLGA8Y6ogF34Ydvxve45nfu9rusDfuJiO8HtEnO6Divlj7uJJDNGg
OoR/aU4uZDJvAbtdtUKJBiDC/hCYBrFoY/GOZR3tPk4uQinsk6VzTw0eBNYl1dZN
hYwqKtPhYT3stVOS4vFh0ycCbs2IcXnCbb94TdS0eF5Swd/JiGCnx4H00N/uofRb
jcx4hjipgQzOG/A9w4RFrdNxUAOy6MUWCe3wkeJYuXlZnx/LuQN5R0Y4TLv2wPh6
E0BV61mfVbZqX/1F9+NhhC1MqFWCZByinLzKjPdazOvzk21W1FBnRlP1SXz106Vn
78ZupRH7+bPv/UezaN6RzRH3x1or2XgIDQD213v69DmTwQKp52AZYtUP82ewgOSF
GwCJopThshVmMM8OldmGZ1rU0TL4ONhOGpMlrKwP300/QunhfgBiRqqg2hAAvwZr
r62+6NyGJPyp+6CfaVpizUeNIYHttW7yETJ8YMClUon3BwRdiwYEwQKz45XhgKwb
GUneOXoefIHboO4n5+YAx/f068da3PtHbwvJUUZ9gbrJiJIG/rHfepJKE5JfJG1N
UmpnLFbjU9BPqQOOYIo2wRYRBVs+Iw3BsgZaOCqDfkFjh79oVYGU9KxIrzwSt+st
9EpW7WaNt535w13ts6kCzPg2AIDaVDm+cCTWUR0iwk33qVuH7MBoLqjftNsJGQBx
hbkasteRuoFNxQRecQhlBoMGkwEe43l1Js5J1GNkIvEuvdLmUllBbZ87hFWWs2DB
TXwkJcesPpdAqcaLTaxDOr5N9rMrAQme978A23U3BqKSP6MRuvZcaUjpEP0YK6n+
/IqxDbrVS8GO+3RALVwISPSss+oLbMXMrEiRDP+uI1hoRbLk/QcxyVzpI7qSuS9X
RnhWFCc/FfgpCEJJ3BCbNH8PdErJjohKmhQvqqFLs5LavZgCT8ul6hMkO6Pg6Zdb
8Wgv7tSlpdW0PlB/M89NbBl38+IAT5Qap8fOjB5DxuE1Ii6tkdNLWnyLvFt1WOKK
MXzh0f/AbCi5AxfMlnL49eXIWil7Mf5tMjthopwu8AlhkW4nRMmGu5xW3Ay/QLs9
OAeagitXd5nUmD8+miroKrRO/czTabX55CHvBnhEP5AVV3UoOer5cu3g/Xs1ULIj
JaS/euBJgd3YtCaKxNhkZGmYiSQI1QsWUFCHhZ1Ts6plKxCdzcOpEPrKJ0XwA+5c
7QHo5FxmFqjGLF/bhSSfK3lkemD3la3wWAdZ0pXZZMLkZwachMZhBti403SHN1e0
CgIl0vqFtk4ZgdoeY7Cc+uIrZVvrUsujFJ5GVJ1yWYRM8Ct0O9+fYePomI+ghUoQ
Kt8ZT7qA7QLc+56M/KA0FiftH1w5cu9dt6vNbu0KyHYT4hOR7d0FnxhJ96fVLtYV
W6BkwBxOeEMHiFoWXMNwlhuFWfo4GKxRNHrpQJje8lIERXMq/P7BgdepnuIMCXjD
LL97jv2xoA2FEzQYOS9XJVwSTCFJGc4y/7880GWbkeL8z9tRaiTiQ8noseaFqUic
JmKnTVbEy0Nr7ia4R/avAd6/vKCwfx8C9g7BJwexLcxtsHKPeigsThQpoA0rB1zN
RIe4myBMYKt1oqYhz6+lzedeOJF0YptZhLKj0yPzk1Kz1jx2UC8+dNEZ0FekPNCW
H7vci/f2ZxuK+QjkL34YyJz8uOW9cIEHNMmJ2dKXdMiT+eqC12D+Z/qza+W1Db8f
WW0yBjVdn0JkIsFtq4dEpbD02oem/AgMxk+9tgYqj71KwpCrh9CfCeTqmw1b1q+0
UtUCQ1SqEBqNLl/3oOeivy/I83+5U6M2lk3eENAn0nlnLCkO/QaxHohyBQizkQEZ
rClFN9Mu2fhGkvihVbyYkbqcE2g7TenV6t2S0JYJxvddSnMYotu3KpyuHbwUgTor
OD6zimNh6brsPZU0vUCokF+s4Ou9B2awty1sfs3l0dCq5rN2MNtz26Tz7yEYf+ii
fAWhdOXppFRH9ldB52UrgojxihGi6yXsHXH+7n+Hgoea/gwNYiTmMct2w4nO1aTh
AIOIXOjk9ERmi03OB6qeJaq+ncnYTZ0LORRSEPydB5K6Z2J/9uS8gYW/k6tsnzIL
qj1tqv8sB4q+Q5DoFAVfjA==
`pragma protect end_protected
