// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
IurOGJKO4MxU2/xkSRXpZ/7sdhLSMNpuIgOlbUdG5s/FZhyCqRsIfjC5GjxncYY1rC37kPRV8pqg
Zy4mIacP4qDib6H3947t/3skgFd8cPMMpaUJ/+WIy/T8NQ1+bf11iLFSDDH/+r48VXNh97jjX7lY
AS08rRDUMtC69Wxe34CIapdY+YHsnBXlbnhVA6hFvTg4zocDIhZXR3kgBo8qby9MxpYDPd+N4Qpt
tjsipxF6zL7eTYRAQCLP4jzs1MuDA+YKgVvdHBqxw5fj8zbVGf2UzeliLytQ/yDcE+OMZm4b6ysK
NOvx1kdi0V4OA8SFj8URiZUxKVNZyBZ+/pMyTw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 37104)
ldPCqx7xwwXWiqpi2/OX9fHYv2RYgHfnFrKwwGVcGL0d9jpaJV+HOMnqXJWf3JhoMlrNor04qDm5
TGyqgX3c38fTDqPmAv2+JQT4Mbmp/tSDVDg+8SYsdhviP0fiOoSRhwtKE5LeRmnz52OGCH24osw+
ZKXZT5a7IDeECmZnYJV3p6hZJdkCoWAZK9Jh7qTfKgfshqUTgKMk0mXSthpxthO5mJKW5WcvJEqJ
KDn7eny0ma7plCRZr7dcIwwlU6bHj4XmQfjwkbW6sbjGyAWyA41MGsQcv80ihtkS2jqgDJHLNuqI
3hgW1nbSWvxIWbs/xa03FslhopypNc1LfZSWtCjqA0Y1S7qNxfvirTqPZ2mILaQ3rSHjX+F0uuqh
S+VLQ1+I34uJDt5ZgJXOIoz5r2qMkERiikxU/DZF14vc2qaFpBOMyw2KquI/fJk9klLmU4GBrbRk
5JjOHkQE1+0IthKEKhm41qNeXvm48l1Kh3iyNIZYgbMc7fdwFao5uzgv9FKN7nAO8Zy46nGB/JnZ
8zxJBQ35BY+t8izlIzRc53VSdAhoEaQ5fPd4PXw2Wg/lsFE4Ixi5TYs3q6oFJtmglQ9Sg5r4wgg4
iPRLrgyfk5U4s8oWEmuSUB8UuN81GkQhcYw2vwSUmlg+SdGik5o2JdQNU+roFeQ90AVOvqzjLgZ/
YJSzR/SN5G+0WDDD/L2gHri3+g96xGhcvVj8osfX2fmiXo0LLTjoJnu4JlUO97S7SIbsY8Ll5jz+
aaxd6IMO8quasrLO9RxcCI+WcTyAWjZf/e65j+xVxS6Xe7Bs3UjhJhVhXp2/p/cJsT84adBhfVs9
1gQWyIXtcEdOCCIjay7t1X03LMjq8Hv6Pp7lq8UDhIVXqGJ+OP7DpedFOgjt8W76HWZlmNn/TmBL
earC7WRHO7nkktJtaXT/k5znBXOGnOkQLIIVmaSl//14ZBTiyo/UqGz4yY8RSHwH6UYKbYEeA+CT
zNloVFRl6aBQOOUdcg2xS5wbK0tyAzKNmEr3r+Vx26WD0bjSmdNV/9h/Gubh9ZInrypwdu0yEj9v
h6sMKdSBlm7fAgV2taFU7wt80MpsjcjLP2x8NHenadK5F7TTzX90cHDZAjUvxRAU3mwxxuiSsWBt
BbV6mRmvonz07EVfBowniiVPFgYeVL+Eb0Z/OELP8aW0MCSOkmUJ/1pLKbukuVt+JIqPmTFXhVVG
PzJwQiHSp6IWWSyDAkvLlUotbnGAX5awV04I54u9Od5rLnLzJLhGwKGsgEX+VdlqkYkLTbZXiLbH
IN6P7C2XQBjG8dOgXsPXlQe6jQanjWIpKmIFg1gSuuLycDA3Lds8EjY3jgaCnDf99VKK8Tety4u0
OyrBy6unFtsDzoCB1z4eq2BbnZFKRM+EfWA6uE7yVb0Ha1Y4zggr187VeY2R1+Tyjg4D1NETbQUt
3B1bKtq/RMdSfBZa281W63ky/sKOYBrMQQ92+UMFRSFu0E/HE7mh2v+QFXXVNQH/D0eZFICbo1BF
GHUwEM4wtg7PyOm0GkbJgJkbFTVEHl/9DfvArOxYsGCTJV/bIfxIKsNeRn7nWw8WLe1jnz2UXBDX
0HNknoovm98OKW8zZBZB1aGKaPeGceXBeqJWvzTofVfaPpYyzxWLZyUGbYGEwsWene/L5/7ea5bw
ZWBw7XL8e9SrQJCvwQd2GURg8tS1rePYjFbTsTcgK+ZR1u+FpRz5tkUmU+eXHimxcIzIIQedFEkP
idtD7eVPNwvNZJiB2DZvRfZj/fcY3V7R7Uz6G0n24XoKjChCUOItJ5cQ/79WNofvyjMoT8IaeIXK
XCI3aC5+stinADFI/Kn7UfFgKIoTdKgq8XLliqAYfPB8M+NJogxqEi4jEKu81Q3xj8/HXDuZF2bV
5aznAJJXIZRlLXwjcKnmz5G30jgKfI52XIQAKsuo3WE1seJ/e8auyeHy5WJxmO2GqP5NRCGXg4g8
V3WFGvCuqgoEKzQ+ErbrfZUJM9mgic8kgA7zrE20rt5ZIFBwny+nS6MVlCA9DYmtQtY+Ankv+vb0
WrcZlsqB/UIZK+jzX5BTFVT4+VJFI1Wm89GXZqLezQMYEHP5XG/6ImIbN8v8vmpLvPkJt947G0s6
T7WaNSDaQ1cyKv4s9xuh2lsTYKxaLp/L3T3+MpmtPW1OClmbtzddW+wtEMt0ABWa+BJDPb+5VD+l
/RERqALn35sx5wFuKy8uM3OpNtL8nrjXh/sFlOsQmoJvJKLGPlKo05uR928lknvNBHlUo8fT6ImZ
f8FcxHqtGjPD0Cw+Me1o+tgI5deDhSBU6zeCPrhsQ3zZmMhfiWI5X62plFTOYNmSq+Lz0Zo86ykK
yEsRu6CwGJlLo8JKFhfe6dnED3bdMftIPQKOjIy52+HqS73eWNCUj2RYFKgHNtuCJ4njAuXZRG0C
e8uAE0LH+nYjjAMx2z3BuyUd+QqactRU6UMmFBlj9AKlDY2ol0QFTCZP9Jqxr7EDaHnrtvBijCyg
Y0w2YpHNKXuDyd3zGQW2ZIQW2gYeY3raxg2MnQXe1KWUMmfnx5uK5pODNOjks61y6+TPJINIdPdh
94HUbCSgKPkyn1+yRD7WN75D3uRu7MFya4pggjHcDIKiUUJMPIDb5zaANrg7KN+c+HJdlb9yi2cm
7aHIE+UgleKlYxVketJxS4pDzoeKmWrq0kFJdtHosfuchDO9OfVd3tEgcz0mIlkZI/jEoUpMp5WO
F94m1mZNfqMMp1qTQ+i+I++6e9X8aPd9ZGbGj1t6bxElwakdXyvCruTmvkNwHyVdlm5EU0hfz+Q9
rlsnuCyU78RV098I8bHyR0qO3QXfbYB6RL6OtwyL3w0nok2AoWbzzLJ08yVHIcHFuMLX6ae4E911
DflXK7raOPJwPeoVhYRwUjPLV52zllTTPkUPiiznIRjvsKJueC16aogXofQVRF7kiw2caD4JIYsK
OLdG9JjQH42jwnD4otenrRyb5gsd8zscU6h9fudZqRLHes6Xd0Sr5BHwr14MN/ym3248JkGUJ7Vu
YHSaYZcwDF5ZFWZGzL/td3C9AEmnxZ8s/H7wDPStMY6Pzlwo83HXhSF5MdieJSZGDDN4/fTy3Zgp
iJQHknh8fmQqgaUXqDW1EQVS4gWXd2DhlcPVoAaYcZ+6bqNIH5tpwMGc+eAcjBvD5uyOPyzzSqHf
N7X8cq+aQSwlvtf94gP60k7jLrPA9birPByS+/G3f2wNHCj+RvzGhXvbFsh5RuBjt1HlsLxpz5Bp
8X7NEkqhbJ6ejbsnbXCJpRSVbvHLZbkST46opA2UTIlvFyw8/9x8vsm+4lkj1Zgm9TJJVUuaWoyp
eLfhStIAL8MPZnjEXnfd9Ybzv75MfhDC/YCh6TMv97eOyJW/OvQQ50sScQCCVEfSCnHmMyhTfvyi
IO8GVhrsOn/j6Kx5NxHAG3fOSF43+aqmuEWRYXzrB9LRh/MZnLcZR3UjcVrcOQEkcTfE/o2WswSl
V/+xfa60E6g4VGRr14O8/xUU9n57oTIcb/WNXfQRPsdUgZWEzi8I3N7XqmhBw+slb8lgq/bYiTIS
aQL+pAg0dBtA1uvGx8uFRekXsQSBajy7RP4LTnLMYPhsdbjBEfOMi1ECaq9YkI80r0cPg9RQN7WD
M81I7aZsd0yE7TO1+Ka1T3jBjzmq4wm5OQdh5D17+5Lz6rgJmpHYcTrdPc30CQ7/G7fp89g0Vytr
ccQelgUrAUcWmjNo5PHG2+dYYuie8gV4DcRekreyndnN+GT7zAkXSrlXMe57FTeOUp16yO80LRpn
B/2qxcKpa3kVvTcuuK3GkU3LBy0SkH6SfUNzI33ua/5zgdZHENjDBz6mV6sNZyMEUeXdTgQ7hajr
uZm14XL7dD6x4NPPdOY8/rrpHGJsg1vbhpwaQwjx+zkQ6LtvselSlM9fveoElsVgTM9l8IxyyGGF
NiS9xbuEsp0ffTmCJKC46zY6zk4E7gdE7G7uZ1LDW9KzFwbuYSY5/0o/HwvTmTVoxMwuwZOt5wk7
1PSQZZgkHSBS757iTo3+TMx6is5mC9RcPNxWtEtDt6Xj8h2fZ9Xm/zs8YMYgXsdkEytBXgALk/Sz
h/PMubIZ8oyA+z6ZiaP6LnoChLOTEEba45EIcuG8eSBLcgR3PPGOSAg60bryGy4qk+cmQNpiKGTt
OsoJ0Uy6rDR9hq+/KdrfJBDrNkCVp2S0ulFadhtzz1hW43Ru/06ZiyYo6kCtAzUI4uygnstCePhY
leLtQGgKyeubB8YK95y/RSekzJvQvo5tDg3NEEaHUZLfuDDAV0ME2/h/kArYdI2FAhOsWerNRSNO
9X980AP2QJTPXWooKDA7qdD721A3W8FSzvFm/z3bII4WcwApaEOS5/AgDEAfxfsVWMrP7/P54Z7H
JTE4KkS9I7fqgXJIS/9019k/1erE/g2f3o7ktEGwUiDCDs6e/oqkti1cG9r7KizGf5nzpPOC+Aj6
F3vmPBQVzb75h5zjJRxLXDG5kRl1/Znre129b0gQAMTJ6jQyanzwVHOgIvA0uwlW5ylq8UVaiaOs
/FXDzo/hBZwlSv+w5s72vagb/85oiSUhZ4p+Bz4BBbe7u95O/Rs1XoKJp6jUXDc3fau4a1cC4OuH
SOxq6LzKXuBPy3Odz3a32hrvrvK46GbyxykeBkmPG+DD2aNcPkd5reRZHcbajTUMUJThsPac74lA
+EGC8sv4cNcdhMQ4JrGQHmJGwPTCcxgsJXp4LbWYzc+vQ81pJFV++ODM4zWmi2Ub7FDyim/kTpJf
GOantZuVWy7HNR3ZAmLcile9tsBYxt5NjxIAqP9srJX5bNXiV28rKBIs5cH6AHoQqQbJVG0xekGH
CT1HpgBBw3frHwzOWVThF0q2HNjbYrq4SksV8toAJcyiL5IsIa8XLVhaT83Fp+Bu5ikscESNlYGX
qz5QiJi3Ad4EgZjzhAffr9R5Q0M6kB7EBRoaDeS3nCUEMCfwljYeaDrOhaHAtCT9ynyojJ23MI4N
svheDfqNskXfp2iqKnOD98kstGjN+Z5LL5W/a9iic5uWv5hl4clDgTWkW7/6Tp5wXh91teb3aHe3
/uky7h589vq7+uzRHQHbHGnvU9ylN1MV4q8MCpJ5QN/qIOUnfHxaE9aYnlv9PqBOtr5PGsDpcat9
E6WN7IBLg1GmYd9/u+ie8dKRDTiMQBltlRul6/5fR/kTRZicxXI8af357D7QFfoXjwKrRTHClWtp
qCB5zpxtdn1HNYU5ZSgrMk8zm/VGNcgnFbDhSxw2TkRkiF/ZnXKDlteXiQXYkWo5LowUmv9KFafQ
yQiIP69uXhPqwvuQ3uDBUfOvHkJxzCglCy/+oAmf+1/BwlrNUZoYZQXrOJw0oaOO5XrEW/av/WNp
VXaD2qFbkyS1lC36/Wzsv3iqMewxq0QcsG0zoSTbei7xlGqXsuxvcErAongJZGqc6VHVObKO6Bhp
ej2LsYckc0xZF2F23d2AdXt/vF1mowOknOAD4rDUqFK5NGOd7GP4cwfI1SzslofZjhZESunvIRkH
EGe6OcIQs+YyWcnGjQSOBXlc/9H2xaE3i4cLHPQPTu+D9DUx6D/o/roHasqSzFzbcMDTTKK6CPJu
0OJDxzv7wRNZscKl9YgohZtVxVcZPisWRaKMerxbaaQ1egA9l44NltEKiBmxiRSCDuhB9k2gwPa/
Sng9MtTkw+jRNtk/bKlmhuqLQ34XaocxwrWMBmAJPWSbpUvUUIX+nxvlzFN5TiWxYH4TmzHXdjwN
eXlBmB988D/ToPZnjj5OlHedwCdy+vFr706W3E87atSXt690h5Btthq9ELK3UPCGJtj0zJECf4GY
lkWsDJoDuGjCiaBHJpLHn533Gsex3Z5IxUa9Ae/uMiQi/kmydhxwiM74oY81iGL/bkhKaw0E6Cso
7rCJ0SuWc/J1lxgIzQvGln7SnwbQ8jrG6OryAEVBJCKlCtRC9axNekrp9cnXzsNE9JxWheFm8jdL
QDdCBTczs//+dv+GmTuxBcMjqeycgU00Zf/pSg4nUP4TdqG8Lg14y5732lzJZ6EXZ0FmFXUrp4u4
47XH6L8XUmOuDnpTrCrBYTJKl0AmIgT2/CfMkhpPtrLPZFKQng0Y3aSsUs4CkTvEOA4W4emn/rNN
UpZ/JgQrbB5NauP5Mc/z8Ju3RDz+VMtIWCQLlkjau40RNusAxe4OQbqGoN9NfBJXau6SgBKqPwm8
n804uMA82SpNr2YJ6pmeJLSraCAWYTiI8Xz9i7Dy2WwY/GNvMt/oC9O04Q034cbDxl/uTjk9sGO5
1TiHdE4rA+BrVPydCE0aT0zzYBATUc7315vB+v7IMuXM3uIPQxhvx6NWdUzMhdo2VyqRq9DByO7F
fbJKOPRY1k2P3HGcavk7cEDtDFhcbRR5l7MRXdoszT9pR8H+GSUcJv4iAgc1APzIsy6j8DFJlkdM
1YHxuTPOx+xxwye7BNGP6P/bM4335a3mEiO1kRDJ8jlLfY3UozJ+CK+ZUrDoHzfQAQKcfVDqOhvA
Ds7yvVU8vMHXu0ILRj2dmR5QymbEH+Trfj7SSAELPukTURWdX2HwOgDHjD1C+bjmWBQdQg6mybUy
4RPgu0j0xcAK0h/GpqAMpNwtmz8I1I8bJ1erb+9BKHnWLxHIF3YGMXAQ23wXgk3Ir+k6Ygpngk0b
uUxXqKwpTmgT4tzDfxuRZwwgblR9rWL9nENWYExP3eOJEnVz6+N0IleJwdWutO/O9J13LT5NsmrO
orRLDHh9HfhxisKNjRy2pEC5ndiSmp9Qrr7ynLKZjPfp+U+2U1mq7oH74FtV3uBBfHI0CcOglYfo
FK+ZpNywHe7P6Wi5ydQUvvJVPZjHn4ZQ/JyKxxEkamCNEVrwOvVYoRxPbUrIVE1rfSvuxT+sTRda
FABHEz8hQHzF4Kg/nmkZWUuZyObb/FQfgyUjdd5JbbqfvBA7Gme9QJrjMczjwx9omE3B80POU762
VulWPl/JGSIfr60FdqPwEylt5XOfl5yQdR1D30YugBooagLMtHU/YdvsUuXQUXMPRyMD3se7KEkC
CVI4kad3SX3LnPls7TxHXCkQw1jc9PR+TVeCV+ZLzFMaABhAiwGZhh74inpsRkQ7fUtFNi3o6Pvq
bQ31nnm08H3mK0TNUdhD+awpYsy3nJoabDKRmJ6Go7qGiRPJV8HiqdrVQw9UK9dvdrXV+H8vTwar
IB1VcokdTlthk36axKb+BDw+CkFJxvf2yNH3yWYPE9U1glJdyRQH0C8wJf/JvvASqgYbvRRVJY2R
eaGB8gOiHZAZuWm2FCoXkvBVn6hGZMEWv9nr5iZbKtweTHwyWWW6OHSTNn1J63VL1hulVKi1nx9l
JxZBRvKbtR2FQaOuUZLZ5tUP69k5yCADm1oly9PhLDasaAAAczC4zB4F1SD5UQm/pRcAMphxQ9HZ
p/Ft92PKmSWxixOlyyh/LNcxeo5cLFzLUpN3qxiTeRNxFSfioi8B/DPuYAzr9je+KK3TYoMSoNRw
Sz7mg/qT51BAtXJGI+9x32IDxv7hamVeBAIc0vNwv2kOIIcHcViuqZw4cjoA+noVBjlJ5dJYgecG
hwddHWeVDEl9/+1D9fKhZ1g267qGn8lL6mtwDHZQu0M30OOabVUVIXzNTGzIBmqN1mJJ1p2/wv5f
2CzJ6bG/Ppas2YiBHCQbEXrKJ/pIqn0u47rLaLNx41EA2X7JkVbIVhYXavrWOg7/IVctcemy4pKX
X15Jv0urvyenu00dQumgfsz7psxmQpJj2Hsce0TpCJIgQpThc4yBwAkTNXKqewwzJKzUnZW/o/Nw
Z0Wn1hsvT90ZbN1hoLbvcS2pqMlZfwc9YFmlir00+yVii9lsdeoR31JML5AZ2igMxcJ5dg4xQwdI
Md8bO+nWezmMuaqAtBJFdzAU+G9JyNqw5ZX2ATLgbVeQF7zM2OZD9/kxyUXX5jGBe4UQUbOa8oqP
omel3/y3HQSnmjPmODd5eZjOiFVvtkKeGg59IMA6WLmytup1Zf1vNDZdpJjyWNGNM6/eYqnu2vN0
XcqqZGM5PteelPo3MNVguB2Ylyp+Ia5jaimPwNPVQFJf4N9FCcIq45U8T36o5DimbjUNdJzP4gCA
dfbK8khE+tRUewOnaglaVNdnvOYBBA0aO6K+xgvfaZGKrUeEV/pYT57/i12iJNxJ0XaapLbCsUn0
u3Xes4sS/5tcf8pC0BDfTBJdXa6uHqnrhRUDe+eJ5IsCQxmfXj/VD8IISrNnRV1urrPWYSENHlML
QroRvOHEUq9MXkTZSZbf3XeuhSzgpQ93v3LaxujWKHQgU/5N1w5ISgzA5IF18y4QDJohNs18OH6r
PwSFkuyzFmkBoloNCy7rX4mVjxHhVnk0DTE0+lufeoaMEWOUSkxNu6Ixn309KkbDpKOESqnKg0XJ
8B7pIsRfRIihDJKODz0BIoarv77hYEJCob2395kQVkz03DG4AoHOVyqTsu4sWAkahmlIxnbVedh7
MPs2vjcri0G5aj/pwUHvVSx9T1RyZI+0xHWwkWpG2W1qZLZMhhpCDEa64vfZxIajpvl9cgwZ1lpm
mj78KXvNcdjfk6YajsJL95phPGmBnAOtB/IL5BoxoUDoi0Vl+sBZkqo+pDy1BkAsdY746Y7z3Kk2
PWK62AWbe/xJjvnM7vmZBv0OIXd2mOMSfGvf7fz1vzijLfPaCUE7hmEYYnEoqdwhvjER7Hj7YnIs
1H0wvJRqglJd5yQZz8egDE0+w6ZszMm2AcqGsQwAMJNvXp4hc+Q4CZVCItXkXfrAA7JN5QHalxpA
wA2VApO5p6+4itqJ5p43zRL5zMn1w5fk4hVDMu/3e6gTQhMntTFHqG0XaY6PN2D3LVqlX0ARazK7
t08lVKAt8vVRIlXmfCBc23SRWsjHi8Cie87Jb3op6VEiChqchw+tdntszA2qKBbBJiSQ7JQoUw9c
SNmZSS91ASUTfZZbHX5472gmp/HIQJ2OSg0qPQwLSDD9j58VVqkQ2tJjBbTQtN1q20CIS9M+inFs
7fMU2o4xNMjtUZijh1xeDX95LdBSzz1xZUznhOIAWq7e1Wdm4PuYgfgP8n2yAVQNBhRLVDNvt7oi
5ZAOqrBdKhUh7+0Q3Cv1GuCqrn475YEnmxsuOdxJ7KOeESQ3ygtuAQn7Kwp97cd+iPWMdbpOdVie
3kIv82fbA3Qu7OkksCc3Dk6ZaVov+aBHe2eeFtkV5Ewk2mugX3sdRW+YDIEqfU/628N+zxkvIjTY
Vs1+BMplSK38Ugri1Vcx1lpIC5mi6EbF+nY0rjLgjmcRC3vn60u6ZN0EGrNPT0paKQzvym9rK7ek
tMqswaKlyBpTLYgBFobj7I7pqVX6HuKsJDOXfwkjKvWg7TyP8WyMVGvt09R3lLdcDU9Skhvye780
/D3SbFQZl1h9HToeqtmclOgE+UY9zi94XXYRhmwhXCxOJjP3721rmY5YcO2tTmVHKJrRvGmpo5vN
FK1xa7XjJRWi2A0EnQDODJgK/oAsVccXHqf08vpAatIR2+6BdWzwSC9pFVka0ctswZefXo5fFBPT
JJcpDJSV6O17hxlH4NLzGqw1FcnL9aNLYHqBMXN9+edLTXBEv5MmCtnK9E+OGdtiHm4yx6aBEy5k
46BQgubn7k41ZIR3sgh1E1FPCtdSA6ttyPVR1iCaWuevlTg7eMtDJPQtFSK+mfunSzvRiBDCRnxz
sTLBQswbs1kCkiJDh7mjH/Pmd+R7HxiCzMY7hkknRJ0ngmt+E63l1xlzbBXF+m+DWL4o7ZAZ5TE2
QuBWVVKbpMr1P1y9KJs2fZ3y2MZdCbUmbdnu+nFyFyi7htKRYfy+YrbzcRDCdyk9kVPRf9dAc3x3
N/bLXRiJAwwfqUFdcl236PRPoaEXerVYZDV+ivUChDH5x5eyR5GsjGy/4bYfCl2FRo4yZ6r7WuVu
RxACET65b34wiInbE2Fie7y+076dbUxu1EYDwqbGevsgL8OoNOIqFelBkDi26oQJYCZTiQ7wLcJl
n7YUJlysH/bwNYi3Dfc77l48tggLZpzGA2e3/ajkHKiL4GdYyE9vdecbMP5ghbx59Z+pH06wwkWe
KL93ESO36co3rL0YsHBJrAqKr1vfH/F66fBCSGn9VKF3hGU4L9/7l9RFE3mfG5TO7BD88nlgkm4z
4OCgsKPgO1eNjzDsm6aDkxy2q+dPJn+tC3jq1r0fzdT5W1XIIcEpPBkf2pc1tN0surfDgQuLOZU9
IewN8aDrgROlQ2pGzeF5yNgO8ks3d/p2klzqhbSy7Fvr+/gbCbValukUxvnt8ZKRGM1hhy+1tv9E
AfB6qk0pqcT2R2eZFTcdLfwf+ifqxBHOvAugr6FZ4Xfn/AZI+nD8F+qyX2pvbqGJarbTohf2P9dm
eOOyNIberRjZEsLtNoN6licAzpQ0SBrrnYzZ+HGgDpROlOzO6L6iwB0QhDbb53zAxj3AsHPIWoPC
pqdCLLL8/0esAtpfHy9WraWWIpGs+lmD2/9GVXe4I2OZ14U20REHqB3lNmRZpibJp+uWDwTuZR/i
W0oIBGt03Qi2j/DEzPHcRxzzE+2sLdU2wtB/P237iDCkTNL0TynHhyakYdVqj35VbuajeGtix0Ke
mgZYa7EVVNNYRCMbuX4tpRoODnUseHD4ewE6S3Eef0GMjS2bYkfstdackIdKvHBMpdz8DRyqnA9Y
xIZvTQR3LtIFClnAeFXLyLUDPjaecsr1X2VWXUUAtAhIHURP3UosZ0+/OKQ+Bdvj3HFXNMhqRE1d
MXy8SvhQZJVQYf5FWNFA2+6V9ardUXewKfMPnjVHfUi6Ds1T92ImuSGrC77A6ygXLG4DyrBVBDej
iNpRj5vpcTXMtrvyqHfjWa0SK76HzBywGWA8vN8JBvbXxSNczbRn56d9aYSv0UT45H0mKGy+Kb87
1YUvTAqE03LVX8J1ohqj3SVvmlX6d0bh0XP6parwHEeQtPy5nEQqFU+dkwqtqoVosC/DGt9qrA1g
Yh3ZbrLocMkQeyU6NEq7utF2O3YGyi/wthwNZSSJbW68FbZYY9heBRlNVybvMv6DhJ9iozRmmRC3
LywRb5o3YKzlHAuAWSsjP/suz9pjwfCVg/MQr8dzALT+xSzaqQikNJyzda1p7rnP7BzP4p+Gog8w
1J1v7Q0ABCRussyvRCuJsvilnOa19Hy/uGFO06tzGZJ188NxIl0Nd53oaT8hlP3eQa1cUF/03odd
2B8ptENr1sNEz+O3BgurB3VMbk5trwo6N0eDgoHM1L8jaiQnpBpNQMd0lmgHW226h2uNRUOh3d4o
5oNgJtRwomwEWeULdbB3A1NphVdXA+tDp7hNpihAWmXhX6+GhseD5MaGnvJ9x0wwuyZ2AypoDN5K
v4PqOYW4PkN8rA+/v27jCxbNy66AUyfVtqlLk2YIFcFrRZDpSfXVKzeaducX5vwWRdbF1j0pk/oW
1gb2aG4BKufVFP1WhznQdoY8lLvm4Wtn5trvZTYlmpB88cpf+TKLyA2Myedv2WJJr+aYjd0esLBC
BPL5pHu9yDgVPaOihM+0/hdsEh47PChdng2A79dapQSsxdz7C0zk1dQViD6mUJCuVKg9IAz+twzE
6/NOTxDBhWBHG0UXjUv/ALW7DOSbjcrk4zDONzDhhULKjerNjW0fynLOSm1w8n5gUI2fkv+KmR4H
qU+wocRubcxB9CLNZayHS890fD8vqpnKFAELkag6QfToy32ox8IHNy5Q1yK01H1xWvvKBg28Nj1i
o2m4aO/F2RiA5MS05eAxKlKG/HWqOI2Lg8ETcuWYujvLliHeyD6bQy7uvaMlgTSbvWztGDeJvqE7
nfwLc9o0zHAN1alOTnmp7XYgoliDNPJF3JBMzhoh2pDcaVYvHkrpeNkVNqQLK1q5DR7Jgfz7sd+l
UExSH9avUejTN2wJgqQ3GGvm6041zzPqwHvib+b4O2Cp0+54qDL/8nLG6T4dv+ZsPIqwAu9WdLJE
pF5Ka8Tx3C9UWn1DZ5L57XSh4w8SGFl4e8XI4P6Ufh6z0JJ6r4uM1ni1Cd/djqXw+wFcmIYuVAEP
J9DejS4MzpYtxuBdkFMxoKSVVa8PoKmusJq9ZOyhFeT4zUJdq3x82rwWprdCDqmAMjDf3RNdFs7K
Ao47mNd9lnA9qdzHffmCITkgEMcYhcIiFf/1tgz1n3zw9fyLRocybMYt2tawuSFk3BCRsysHmVzG
0HuAFAGhrZ8DLx32WQ54I2tH5r1mJhKpbZus6RmjFv1ASjQGgH/lLkWC0BqSIMQ04FVuERZm1kWQ
yqviWLmf5CxGR5hsvBIp1QBqwDw12jK1QB6o4vPhEz4rOt+ZRFr0y7ZY5hmD2y7y/eI2/YdXDa9S
nCEqW7zW57nyLLopllm5AEASly0sGG73ec9Pq/LDyEhDJkrkAkqqXEPW4TVPDGGT9irNqljBWK3Q
a9LLQ5xW1BJklfr+XhAEfe0UFBcL+CswHUWZEq5ma+IJPdbW4QR6sCqreIivBbdzKFJCpOndxlgf
xF6yLBq9ri/3owJesmV7EUmIe9OItOAsvNol2LUi+CROxhoqVpQZ0CU5iaVIGkQnJA95VKUO0Of3
3TtGJRFmbXFNxgUym7ib0V9/OSR5+8xI6tTJoDvqTPSHsDUrAp63GQrpAH6km1GA+jkVAN92VBdm
2J0LgV9nyuZQvNeX9h19SjoMZcSv026lSb69fBr5NaNi3bXvrcqDwZqJSERxDo5u6/C5wfV8CGtQ
4D28G7ez0514250fpIpmYHHTEDBF0sHIAq5Qb+e/gBO4YRAocdwH/zP135I0n5sbK0j4J9f7cHZ6
Ic38K0DVgHhst75hwC+AUJ8CgMWpcaCW4fDAS8g8HpxOCv1tDPafFtAXa5vPITfndIp9Tj/xuU3U
G3VzBuhSawGWDgviVimRlosRlwyXZqnufV+s98O5B+ulPxFYPmLiM6fdHU9es4hDVlpp/D1n4xnC
eeVF3jnUPvlPup0dW1/GHrGQ9/REM4whur9iKQ4mVPKPaLb2M6/Y4gzZjRRFsBeT3iG8NwMbzMuO
B8iDIN3rGwSxTSp0viOkMGZEXn9OWdb+qNXftc+LkxGfGXY/tXtNvagRLeQxwDbkttJDTscMytl/
3rCpJ9rx00p7xbWRYCrwACLPZiJm7hqlVs10DHv6X0d/41EL52MJlS1MUFqbH3VFSghVqyZiXNIm
zKhmGDgWlNhiJ/OaowDZKNgiFnzY1SrC1PJR08pT1mKOlkEukpKXhzJXG92GdIxwvLz7N0AOiF+z
1O3WytrumSavhT4GJ254/bnnBVt4mTbGZw84G8mWXqEwXyi0KSAPNgpYfSmSyS5mPuMgEiWU3MMu
t0EnNoX37yYR6wctXiDAPSUqKX8dSsbXzQ56z6W0zmbOsF71aYwYa6TStyPC4/5ERJmMHt9o9q1M
7u2XjJBXXSPIe59H76x8Nnk7a1yudk5EzjA/O7YJ7J8Y31Z3PpYnfb663U0j2gq8hrYqtZpA5IQq
wbapwvjrxFvhXfEp0Wb2ckZImM5zaORfHncpHSBmndKKgk1JJ30cSYhFdlxn7hHgF92sjMN0vdd6
N+sUIlSzT5SPQR3K+004tZ5zQoYa+6dPsmDftVY1sOPo57FD5i1t1ow8rR5fGL/KzHMKmNbCCZZo
KwtehlcdWQ8VJ/nxQH+6RKgjorZxFr3Tiec3iV1F3ZX9Vyna+a1nWPR/N81A0OfenK1IVt+LX1bI
ccspRdcSHCC3Z3xNPM9Lkds27f0VaUksRUfVmny1Y4/UdqvXuoKpFCFAmHY2S4nzKqZ6dpuHhWUI
OMXvPGhMUlyJcJAEmcs13cOipF/+lzUMxrAng3eJAnbrcSzpoe4H33XMbLUBrDURFCurf0cZG0qw
aWHPbL9FXHlAGqCOcET2PPmA8oCQC4JHBc62j7gtWvUD9+FuiHk5d/RBVbeQHx9WVntjbNaWXp0E
+oUI7jlQUtf+8HVe1itJykjmCLRXmU7xW7iH0IaM7cx50UQhWOfJVZimnTlZAP5O7SlAhprkV2KZ
vf8TW6s7n/W5ckwa2//rRh4EHDs3WrwSVNuVMkqZGzKz6AIc2XkrFt4rS31lHyo8fO6jYYShn9Hf
s8jPp2LqM2hRQx5uQStmgrzX+F31fwEd5sHiglyFSPZ+pE5BLtFanVoFcO/kmqbVS+a1ebukPsAr
SQKYJG7WGiIk1qz0UPeZqt+lsy/Pn8zlHCnqmdAKefeHcxNJLAhKSBDDQL3tBZti633BnKPvfAdp
oX6yICWTxda51NcXQ9XNXrNfPwWGMGt4jMHdzdaDSvzLhe0OVIi/yqSEqKT/yMXqommG2mIZ2TU/
rS59OtJKjKkoWHPw9tte0e86JjsJ/a/Ur8ICCA2XvaWd9Tb/XSnwCyju0HY84kwCrW7F/eT0rnw9
x6vop9alaiXWQmpfhq1ttYEvkq/3bIlSuS5424znuRbO4X4v2hBEUralDsXKraOPbqWA7jXc/GnS
pjuXsCWRS1ZQkblFrSoep5DtkWhmvfcYNpKDf/FQThtq9UvHTJa13VlXVbNgf//jNo+gTzYWtQS4
hn05Lo3KbhzNmVWocw62nGi7Uck9e8rgEcPZA0rcsjX1tcnPOa3vQRtoi0XEARA0snvukUebyOtM
or/9xuNP2OG9luQKXEC0elP8R+2Le43hqeAm/JmFNO/qWZ9K7qN5fXSep+Ulz3s4+D83ZWqtmdQI
PKjBjSKanySKCLopuq/7UzyVkRdQo9MLsirZCPNrAkLK2GFl3SRklXteIS9kfm9pQsSP8Azyqdfr
khZFkH9qlIjg7sm6TwZI/u0eYxgRH1g64Ds4h+B6+ayKHvWEAWYxrBwTM9MQfp+WjfBHbb7ZhjZI
hvi+MdnUdtt852nV3PpbFXUQM4yCIbpG6SMSd30+9bgbrzyPYvZACGrnLuJ62+tWTl6MJKKiT87V
DRHdTCjbTzP1TmwUI/P4DlZfOxXseBvXdbhqjOgz1SU6SRy7P/hhTPGsTz2Mtgccoqbi5UkJItWN
o88PNHtxisxrEcjdC/OvHu/kGkuH2rVkAAo68/6Corm3/eiGkjcTmiZWOLXojDmAD5vWl3etZqdS
GT5zkEjTHSeolr7HlGz31iL+nGzVZdot7l8Shr6Vqu/M4IqVLxafdotOexemzNPF/hqfTrugdob9
iYjrJh10LcFcWU5xYgZ50RJxToIIGyykpg56wIFp7tg1uo+hMxfFf950ygk/pPh7/1g05hEaRN26
SvNfHX4tMeN8Y9wHJXeRub4lqTUmjc99CJug5nPHbimQZ9glfiDuzYMy6sKJcEoxxqdh4590GS2E
7yS9LTZUNwhz7suDi5xxaTKm62Iz9RqIXn3yA2CkWkS1a1R2GB/71DHsbrc6X6+QqZzxvJhyuzWb
9MJk9BrvDB1/Xs60pC9UtmMxON6B6eDqywOKCIXOK35/CVJvDp0AGmyx7K+nDDRKRSWnAQPp/C3u
jequ3/ZKH1ZYY0k0RWUaapW8PEgejbSQvD6U5do+/u/3jVAjT4jMXPrG0vfbpa0DlP983IGmyUMs
60XBdEC/AQlFNvW1OvH1Z3gRX1tr3H8praXQvqstmwOGTPOGa16BdMf+yGgKLm4q2ki0OOgkSDWx
hmRG5MYzgLBO3rvsdDlyahvYSwNSsb7uXEh4CvaHMFOPTZwNOcKIYoeaFEQ1RbySZaX+eY5SMbPD
/Vg5lcaRRExwI6c7RofuU0OmSd8RJGbjaUylaC8bPDPbV4/glTnefVztAsjyxDBD8uwjrkONGcTk
tMmgF7f4kny5rz0/+AZqZ1Ap0VUp3iiDMQgpAfTNK9XrNb8f/mKcs0u+oN6SOKK41zTLpAXW0Doo
xfDTOnSvIxhEu8KFjMek97oranrR8qsKT41z1GZcN6IVvb9aPauuXIytnplkw8UTTna8gXSPqdja
pvCuUIPNb1MbDmAUTBDdSCv1kLcyhzgPJKiPE9kwNS6DUhIT2r2wAXdjfX80ZssmB1LgtvqYH/xl
GHIeninByz1G1h40T9Rx910yY3xC5hqLvVTIB4sAJnbtA3+1JnzVpssZNE+R0Cv0yIZ9UxeWgu8A
+8/y4+RILrBPkYohUnL4WbG63NtBtz7utJ8rX5SkeVcGNz2C3LrFvRDHf7frN6BjqjsVipeVQ38c
n36roRA7SEHRJNXnYfh1WJOHSsiSGtgJNsvNgIZeI1M4PwNWQhh0/DBANvyfeDKdcn5xwdL3gc63
xAP2bF6rSCGZf7ctv/Y79Qalt0xMNJnuOmwGIH3W3Pcbh9TUefgWmLixTsy1M0x7khbX3vnffdS5
9O5+jC1eTFbtL7O1v/vukN9rZk82LyvOGEN5w8WZkZiFr2AeXAA1U7eZDapoJHgDbjABh+Afd2RD
RDZ3l1FsfioqB1oTD7pcFNXrrE19MDYynyYKJO8rIJG6A0uTVL8yThVJrKgRKDcsN3ZiPmJlGveA
9fmA1VxgpmU4J8UA2vdCP5MpSu9VT2vT/U/r17x3t0xIuZhgNchC/j3rKAzjHVRDnhT2+1Ybn2fd
Etqh/79+NE2hwOWzLcPlmL6Xi/n+PE7+wKISJURUD7RXbhNCL6an+Gx5moABLm7nxeJBckSgeODJ
K9JcTqGk+sqSzNCHA0Ets6GdgB7pAohrInK3qPjeseuiwuV8fJTnt4xGqMfEURitOFbVt7T8THwk
/zj41d6fv1oGJ//g7wFEq+dctPWnr4kCyGkXPw38soF/udgI6D5tYS0dpx0Lyu/xkF5K39VlV0ak
4n4Hi2akzA0lSTj7hk9xl0ZMyB5iLxJyXfOBxvxFaMkWjPEzuLUc2ED81KWoMuU/H3Z5IG5eEKy9
TB2GfOogwqfULQ3046YBqJslPswjzuqjJV2i/kf1IRiBROlrJJFt87y/rtM738jXBftmLPkBQfMr
lOQH6wC2oYpWwRw6m6EZVdJxBFlqFtyMKtJZALEUq2e+PAxE3wkrl82FTuBtBpJluTXDUKm2gXGx
xK7bU//sz1QYbisIi/+PckDxIsu59mI+76o15ObjoKVhfMhcFKNm+NSTxWDqQkKIO7vXj5AKKT/e
RBRNaqgQlwz7nrAIPhPUnPMIbB84D45xgVES1vJHO8G0qDmzLtSTG4pPQ6T+efgl+NzoKgrb4qo1
/e/O419Rsd1ISYazOAGqhfNEHyHZNIiXAS60xxV8Gfn97/BVZiCr2CETX2q6UzUVCB+wsnUm8PKh
kn8hdqZJ85Dp7q1NzZFIVK6dEKLZjHbROB/H6gVoALD72Wr+Z65KDZJkEHMuZd6T/r43J3rRB7iB
bBFAC3zCSMETCnAjchMSx4BxvQcjdW1bQBRdx42Ix7k/0f/QxFPfgL1cGX2vo5ka72WeZCpGyZWI
5erRx3ETrAqkn4C1dL+0n9DzAGqo9Mi5HQq09gMoIMh+j3AxYGSn7dDe6PQemVOO3IT/D3eZ63oD
tTxE69MNn/EyCbib0JFTPTcNwhJkBTZT4x1wSlWdoJ1v4KjasCim6GIhJMRa/JtQbYFBkAumajSs
JvO4AhWUIXVEV96Jx20trJYlP2eQw48YfCluLHogQZ+JJqCcta5G740YqK70lGzyrRvVjTpBqYoD
srR6XoFUCW0OuqulMRCLil+31AkfZIPiuOkfKOvGtwXIu2SuhvXkaP7/8uFK+R6U5AEZNJHqUFah
x1cBcYYnHL3wqoKc0ezQmHnpGfKgUpRlDEXb1wwh2sZdn90d5YPOGBohb0xFIBetxOSFlhVvfqCO
zPWmyJokk6eLXeMvTkaVYlqUaAej3/t3VjLjZn1Kl1VSYiXB0I/QH21SLNG5LE5oBbLWhf7FliGS
IGD5HpxE6JJjto3F2u/VGmy34nSFZOAJPekixUOi9Mt3uW4tJNXvliaEOU3WYk9TDnczk258kQWJ
vYwvw/J5uJXdZEvV3TDglSmGOhag9fMq8XXzz1r67z/sCHZysjUXNB54i19zseB+6ljFDxEkHsg4
AmK6+Qgz3wqn4O3cl20vkIdAobW/sm+Z9xhaGqi0q4IKPKAXdDjU7xhv3aeqeBqzfxgqydpEFwxP
DX8DYZ/7L4dsIDgtanFjJG0KOhKs0tpcm4bv32Zjva/U06CeMTvt1ywe+/Qd5pqNAthJOWhLZA+l
IS18C4qtkllHnhVAaXiMQEQ2iiU6Cx7Y5aDZFMfQbULr952ocOg4m7WeTZ20euoUcValCjclDj9Q
NoC900XvUJWFBlKTJTmp/IpG/G89QB0ZrfzkrpqzQb//BJAvvGBOGMpPm7zZ5QJMZGv46NpSkIqE
4DW8vytOc4bD2BAm0+VO1wT8WPqw7bBjyEMbFyG2Wke/dbQx8WKM06TUVwiAEjXzwkexSYqnQxEW
Mjv6wmSywoU3PGPpGRMwdEO71OsAvQ3byasheIc0NtmbTS352HCPoPoqFlqIuJE7F4iMq+Nlildx
Ini140lqG5CvHkFppPEEUYN9xZeuc5z5jpPWZHUqC9qVy7IVjk/2vzNc6GLMt6XBmPkGR5mR7iav
LXMgos3GLvlqxqtkT5ndPmWKIHnVVsEvJLd86ZLqaVRQUJaxm1zTFLtThe0tYub5qFf/45/PNcMr
O2weP5eFH2eAwpQ72Bz9XbLK8m0RhWE9PG6W7WkFZ6umMECY+quvCKTkHn9x3mRuo3tg+8I6XFdq
e41nWDbNnjv0dtR9JoRh7Y7Q5WidXwu5K4BjLaTVcAVkq4SjoFbEgxlzFK0KCnWqsQWntaejm/4+
/8s5f/xGTD2KrlkfBcYE0evkbgZyidUPShZc3XXxxFSn3boXLdGdIcsqE0kSz5qOrNzfNVziG0Vz
uGJuqD5dUBu4USew4LJyEPu5VC/n5so0KkoWLt0VeZxRHDk4cTh0E2WTbixqACo0W94npTkI9fzh
BcmqwRfp6MA88BH5J0uq+LIgNrR8j76TkYxRWzHbfOvLndCmysB92p6cRm3ju/1bK1KbvzNOV3kt
ZVlv9gqWrpV3ynvZ7roRhgFdZmIj9SXxB5WPpX2ys1OS3h9wzGr2OVTaBumqGWu+wf5qsY+PPU4T
2F4F6+67MqVW5ePHeiGr9LqkbP3DKEEw3j6+YdeT9+GIcjp5A43nV/IWwkYgy562kJsSYl3mSlJX
y5Pnp5/hNQyC4Qm5cxVttdG6BKf2+jF/dYcnWoKx3oWzcqlNxW3mkqze9gUWXb8VEwhlFDPrbV1z
acuMYI70Kb/ox5UdfxC11LeWD5/2bHdHiFOj/yj0ycY8XFxv1AbUjfIaFBOUFgp2UXW6cPu3MGZH
m4wjuZreVb2neQQmP+vBD8A8ejiGW3zIfQt1Cvh1sDFmHVaYLrrTxEUiFkWl4o/oYwJGg/E1jagW
uxyxstYkgHMfGK2KgmWFpag4MD6lBhK28LPHTW4NFm4l5B6z5dmoN4s7DjYBg9ONOiYBN8uEJQuC
zlPnGP9HWS/OJr6m+E0Ul4uE1B5UkyV46n8oV8ID9We7/irh3JtGC46a1sZw1pmpTvk51muKkp60
c2m8CfGM+if3vwE6XtrSWWh4xPKFnsL46o5k7LvnOMxR1LyzBex/zaWiIdgem+bwpcl4LioN9G97
6ko5qAAgYJbRfbivzwQxTi3WaS4ZsHaXBlD8fUK5Hhx3EpTgJ2oSQloT1d30HE1SAhuIHoL6iAEj
wHu74/0sP1UUd1KLBtsNS2ZzrSZgB1iweP802v1rucz43uZmz48n+GTDSWfjZ8nCenxj2lhSyb1K
IQF+4Cegdj4fp121iD8vClIEND9K8970vFOGAzclzu7Jd88aT0JqvAaeBf3MEEtzlloPnzjuzyg+
EK8boHJ8fy9O3Ai/+vMZedz94hhaPyZ5IBqcZJdFPhNypowhfQHqhyEmOQd5YooJyjPOg1/f/27S
habEvFP5JpgJnGp+91mZocfvWrLF3wBqZ1AhK2Us26biLJI8aovBICvb/sGIHpyJ6JxuKk7vTb7s
g0agqeyL4O5EENh1uvTNevbf6ygnkDaBOf78GYDgxVpKI42oRF3OcfZ6jMw76Y86C4YdThiKUSE6
5YAz1qZFWcMTKJXH1naJCC/idrabnx9JhtMJN/rshsVucK8R6vC6fXjHCUnsWbOuWCY6/uIA/e5n
hZNVUSj8G1SylaSICpeH53r0ROqsqDo/Xe1kN9/7cowWbL588RXsTfg3Iw+h1BS68TzPcP7sn4F3
2twG5QAY6oH0vBK4T2ctXH5pQMrOEWqU1AaQ3OBDd4FcQ09u6Q6A3iOn6Lq50a2sgYwt17/Ihf+o
QypUufMzJ9u+Fg7IwTH95CudMGj5MuUM49ndwGxNdv50bytS0QzN7E8r95XEb6qGj2ZhZaCdrgeD
LCg1nXbX4z8r7XFTShIsIwykR27cvReNzMUFOL0MxPOiebKoy5TRt2+BOKufA4J8toHk6lXyg0xx
vtJh6t5hdrvmwz7AhDEEd9+TvHQG5LNryjJG590CQOyRKHQE32ktYhrC/vqIuH7EnXBRppixb06B
N0yCDisuEO5Y3MO1oo1bFpL+AvML6gkuT5arbPr8wxcUuwdP9b/iLFH8TUQ5tFn8n16w0bx5ftFa
sdM2bwuKPFhcoU45zKV4zLMJ9drLyJD6DkiYtFwLW5RnEvumH8lt9dq3kizsALfW6yqAnfmeR5FA
V+j7fa/DR0hPfBNFRxCBBN6JRhMYoNG4ewhpVElOeQPCZ94LkTHMLcg5hdon3c1g8iGM0Oo97Uma
YEaPr4maSIyLUlKf6h7R8uBX6PV0C8uMU9Ku6y2jQ8D/oRhfQ1+zHB8MjcC5aHGX+zudfWWeA8Su
RfFwuevYByPIvVCxLaX5g2MGNXGqBi/BsI0AMod9Dp2hyqvfOpDni23bgQvJ21DpXiz4wNB0BxsA
fYb+hRJnWSRek2MwmJjgL5KeoW8dqmUOqw/oqMGj+X/98CRRU3dGsQuBZPeH5dQ8CKgc3Oj2hD5D
MHI8ZIXR/2cUEIN1vzT9eGH5G2hvtSkKPX6SHQuDXAS4uRYc7E6ARVWD88/lc7cAkk2zMqHUbhh4
6uvhID/460EQzd+gDhJsd3z6POB3S0Lb6fNejtR5jcjuOfFt4LaPSldM3IRNfkYCOCQ+p52hJ3tG
bLpsTiO8XBHVm0bTOt5ANLR4KSZDjHi/1fdAscp3/U5ZuPosbWDhe2R+gNbJBPcyIkLMg3Tn593+
49VXW8J/UWZMrjP9r0OK2kuymk9ReyWxe5bDv+8xKNhp2Q9SPVT8kHrfXIF5oFwKltISAe4jGLhp
SaOnksS4IOvm6jMj1mrjGmUQHKFjJH6SONrgH3L081LH+XCEfcBlkNoL3fAp2ORitj8MoqdLHrfB
hrvdv1G8xNdv8rn31nznF7nMeSPbofn7IRuuLNWvJWZ0r1VsWUl8p6tKVSGZrNIEHcRGMSbcDUch
AQS5gXfCCacUz24X7omUCrmmeQurIdM5phM11kxwnCSZEYp/B4iZIuhOcXiePqa/ZoA364ZLlH8j
4oZjlMLMyWcGeiVfah3JdN3dYgUFLBIIDfqmhuByz17RxpgZN/QvAEByrEgl0acgDoIX0ru8Y613
/E9KE/N5Nmhh8fLvjdNUmvpuVHuIaNaa7x4dnCgH1qQrJFTDjB7r7Umf8bilZdA322g5PpLJTCen
TlME7PCJWuK3c0goMBvs/dYMuJhUSPQ7e7ctVOgXSooSiVYidi5/PvLHIr2WLbjJA8kFjWRpQlh0
uZ5dg5DzGk9Vw8ho9fGfZOh6z/vRba0ro8gyLnC8dkfYGGr7DiQCPdcPgy4of5trhr541Tfzk2/W
Zs3k8m+sZIb6rWuvXxMWQf6OwuvIxgdtbumxLKGM+862rxKetxAr6Qmp60XGeTTQgAHFRvj4uPDb
C6XuSYVXLx+x5kpDAmtRc+tMzCgqTWnG3pWZCtin1ttefvlMFYqqFXLlj/6uQJNJiFsTGCpxWLR7
C9krlvFudSt9GLBlRYbcObIswIp7tRFfsiiTqwDmvHFFddWvU4Xo6BjUotL6dgV4Qg5doAVQfo7u
DuvsxVSiF3KaxKVZetMRoFuAnWz/JXrIn9+xZoqLL5iug+ouAy1wFcNF6lEj7wbV0yJsIl8p9Gtm
uDvblZdMcjSNiZ0q0y8QuHQOMAVif2whi+Lqd+Rb4jMR1rwMhhSov91zffA43+Ts4AgAHlYGBDKs
GwU2Y2wrYzCDGkNWdGLJwoLikKwFituDSu5B0xhzCKvTQviZsPAA9N+Mkll7j76HzdRl3GfWqjkb
3yzJtkfTqdcAVBfjkckfH9TJFoEwC4A333XuLgbfdnJ2nphGtUIMFtykuYiWNSocv0WOOnJAya86
17Ls1837wJmql5qI2owTOgPSyxt4tDo5sZcMixkJ91PQPqfymvitScoGPrchNewLEkWO1iOul8Qe
8orCPKZMr4ZCvcCSEE7AaMIr1Zz0LS/4Gh7dzZpRAS0F8aWrWKrnWGQZYUddfr6R0II+JBdpFST9
I4dV952ee40zx7AA62IrVbc9W9dK4lUtqdsFJM28DgIMdvAeJ40By1fWfp7HBFjKLLFwQES0oqD5
Ga5WfevdCggr8G6qycAXwhRCY15JJRDALZWKSnFZzLp39wcvt3a/NHNwNtRFzrdUp989RFAr1+I3
9+mXGxd/okUyO02A8WaN4tnUHQcUOKv2g1pPYLgZBJmPcfhH/xQeWilhj58dEjTtFZkrpuTi6z1c
m1bHjws8VCxwgPD7CdUTAmAIAmXz0OKIuSQIXfB14mOCRxABcl0HKgRrCf7arXTPqEGflyEX8eiT
DIUxrK7kg+IQtsysyEnc2wiOKH59wA9YUaqfWvBb9SFhbQ4k4rcCjNZIGJNWfienl6bVaHCD7ROY
R+p1SwMoqqx17KR5eg4To9PZ6p2gbqGD0usRnhowP7f/5EP052p/JmPv7gpU6/Q8JLLv4TRxtI6O
Bd4L/Wtbeh/zX/dzN81Cv0Ms1O9cz1w94wl3m4e/TJ+np0rq2XmZ3Y1tCXjMoksyvz20EBuIZyIV
Dfp7v5wKrxoPPpgHV+hwRqd6oHRNnJFH8EusBMhZqnxLDO9ZzKukmt+Bvx3DwCAXMSgqQoKmqifx
85KJMjRvojLaez7rIaUY2qfygwhDrZP4QnQO0iEpyvhsAqGJ5Y1Yzerq7KkJa5BX5ELCK7wwf6Qw
iqmaS5RY1qVpxkMvK9q0Z3ojutVgvu5EoIchukELrNXwUWnBgcBFTYDehBmxxuVs8q4CH7m60y4u
ehtqwBd/9NU1VOxQDoR7aKGAiFXLvdEb3b0R1lxHptOJYyPfPsYSIifQuk582feHyAFzHiHeZ9hI
ig5DPUCyEv1/cZNClMdeCAS9oFLmPUH2PaAWfIz9+C+b6KovutJz/QvnQHIDHIemUNtCLcNwWeNT
Mix1EUY+yXhWjWMDiT5/yMS4ptU1MoTJg0kmoSDCvLCu+BAXVl8Is1DfCXkOV8LkUD3IeWOHuQds
kKwe65v15IoDa4hzdep+p5b7LwiI+jRGY3L0sG7P4Df4GZ3O0ZGiG2bqiBNVEchrWnNQ3IbjkgY+
d2V+6zkYrffTakpZo30ig+uHdNDGKbUn9ANPjCqYLcCpzxSKmfFuKH8EOvAp9d5Zy+yGNA+YXTl5
LclHTY3pL9kQBQICvPTmUTH90ye+WAmMPphe9g/S5e+SIJRAY5b8PpPBkokUWd8wh50TNVi/SYzI
5QBleFZERHY4UyHf0b+JVC7ZsykRFgFbp03G2sHKV8krCq6goC+0fWXDyTQsnURt9vGhKaVdP97U
KsCerhxkE3xOKBzd//7aGTl6nRgVCyd4zKFxpe2coOtiCNXl1P7svH3W6KouyDMhgLhmHMvwpmrO
dLhBuPsd9EINUiCyGqbNvpVvZ8OBbDdsWRHKx3OukFA0T6CENbUKVR480SIk8qzn7r7xqEr7oiYe
YXTmtI9Am614CONYTPjn+KwbzAWyjlBvI6qnPhSEz19jyjLUru9Yk6lEmc392G7tssDb+16DpE82
PkJjU3oPj6Gf54x2gDo4ZZmGzHibuLNr9veUEvX5INs++6/7dnsb56YlWCEnWLsF+uuLw2KCBSed
B8QumMJ74JUbYxXsRoYNJtqdoeehsmcY40vclsOd7J4J6vActPP14b1jAGVt/O1dnWsWGbKdczkf
g3dYtnLB4CFF4HFTuX8n25J9JO4JrJB9NK/DbsbOjSTTLpD9Ohh5VCteSZ0qOJjcxrjC5H90q2iV
LA9ljDwsOqSnlkoGGoSlcb09w0iGaWPFUfBACRlv/OyEL5McB5nWLHO4a7VgR/6E7uWr3ufFqo4e
EOIIZ9EJ8djeIzMuAi/NTtBZrD2MmATBDwFlgEzPxWI86vWPyPCSguqLoKr6czMcpU1xG17pvjKV
3jyg4FI6ePmTfypGeKljRXWiqezDN2pNMWZuhI0CoMDcsGMfy6rVdzwh2Z78QDncymlao25zfjxJ
2KdJiMA0ALRxeZj/5Y1zSvUTE0zVr9xViPC2lUnSMBMCnyqWdOa5eOlDQ6NV7dMRfFMF4L1vgwgu
hEQodIGUun8ncDhijM046fW1ULYGWjgyQSnNjNd8p4/YuECony1XBsrP553fYBGG9bZSU/Utn3cV
ahqOnQxafc+isOimC/TLO9noBZq9Tth7LbZyr3Wa1YqZbLZoFopOZhQ5YjLMxQ0GAyuoVeL5iPkP
mf1tiqOg1nmHdoCasudGfbM4C2g5MEhnTHFzcLqE+SxhMbjh6KWMtyXSmxsKt8WzAd1wi/G2IPTU
oOc4M0ZuzzJLSba5woI3RmI3iayj6L6N0jNB8EuD6vjLLzeAbYXGdjGftu93mOBaAGnanHfEjwL3
x9+GQ6njuBUxEBxXwSymhjwgwkQbGtu12/FZeaMrQ0YDUK1G9PQ8x6C0QuIcQny5qYrGTDoAoPC2
l93VwfvwcLf05XuOHATtoWl8zqROWzB8O+4l+NIWGWTX8Qei4Z75lsHSYyfXS/SrcP5lgjm6Tllg
F575ZHrD365LiAGXnzZV5YHw0OcQbqdc4EGK4OcYuIJ17oB3FtMMbADgF+I+2+l+JYD3vj7yxBX3
TCBQI6EW6+tglPrVwSo+HgoIcNooz57BYoJv5tmEdfqH1iV3yqGh1ftrN+CdWjsnYuc4HvTrrWXz
y7oVewBit+175CHKb2o/94pM68D2iPoG9poeQIiZ/gj1bPcRBDKXaoUYKFxs2eIEDOsQMlIuR071
EGmlm6psHveIHgAIDa8nVUeaq8s5dFzFN+4muSbv9qMXpM3/fODDA6v7EJIPY3IXAxJLd3LpUeLR
keWrHgae3PyD3I9Lsc5Tu2AXk5SYlYr7q67KEE8AGbM3kpP3dvUDvL2+5E3Cd800ctVkZYQ7YkY1
HZ8RiUKMjodXKvOicLvtQlUe74mY2n7MBHcIaMeAPw1rVVP9cuNlhNIcelUW9nrPu+kFhwyjH+ka
8XrJbDt5fGYixUJzkgsfMKqt7w0I+VM/ZJQzrveQkWgELJDsYHFiNZvy/6NA4ao9i/Hq+p7ZMS/z
JI36U+sLCCbkmwcVvfsoKB7PIenL1GUExH+Kvx+FEuq655T1NfHh8bP1LLNkHA1ejDrJijsGd80r
nI8H59XyEi4ftwSEuHgbO2432gNw8jS0xSpXOPR5oq00ImWpaNceaJnpnRT9QlzpXWQyrTWgGpcW
BOT9rFPKi7LSCA5CFQMsho6GkMFgNWuRNFu2BIvdE0DZXrv8H3y7JM6owqZ9OOcIM51Qw52srntd
tEf26QmZoVV+UtX+2FozlfrzcDT2bGZD7nntXGti78HqDlVFlcjm2W0RoqTqV02o8NBu340cXYsY
2kaSboxbXsFYRDh6OmFYH3I6v5yBnLdUPMKbRfCJVjjh9ocT/uLgK9BUK7O/4FMBt/c25Fw044Vv
9QQ/IUkB8tnHUmZ3jBBLynB1RNoCBGvT05ye0Z8MTX7J8R7V0PH4XN4EPtMDTJVu/Dxf1zd044Kp
+U/79mlAxJ3Mvcvp09XMz2Qk1ddnVcsBL9CfDF6KfSTJVNNNWQnjT4NuMirGmObJ2fhpBPedP4WE
feWIyNw+leLM3DikitsdkQ4ofMwIgfaX3VV/2+0VKnfTgWpnrhscCDf21L4PhWWzEkS1s5/Y9tJO
/aAG9FN9qFk/fToH6NAsmFPKtfIJTJsANuw7TcEjHpZ3elXPEW1nEw+pjWz+EnmVh+H9zV7FO2Qq
sG+0WEk0uTW5P5MrUeHxSsRUEwQFZlE15jLhawGrtyPrVvLCXaBHqG8498hZ1tB1oKwKpsQr8GaH
q2caDffsbaHyPsS5uIjW9FZ8Uwz1VS4TWf0DcEBeZ504DnI0XTw0mQ7l2oQjdHDLSbFIz8lmb+qK
lWDFG+bgbsOYbehxtDZ32uqsANvNPgD6TvzajHXcLX+xAzJSeEdE7aOcnB7d/F93q/qJRwo18+qd
CCbfD4qg1v+VrZFsXhG438NgSAX0/TEpsCA4TBan/wyTGSkm5QrB3EeMepiusXyBN/6d13jTTNP/
f2RoEFFN+snWuOXd/+GewjVsxAP5kxcCOQOCp19Aw8avbbu3gNTCY20re5XbeIe0zaTE9dbVcAsf
Pk2kwVqChrpNHiLpDC0ut0bnysYtUcNBMPnrIm+MuTUgcKYt9pTDN0rNIlB02HVzEoSxuPEDOQsp
K8c5T/Id0jx8dF5o9H8sycUwlE3sB6d5TmGRzr7vJ55Zdqx7Y1yq1hBa9k/Cp4OKvonqdgOr138M
y6rDyorbN2Ossfs7yf0sNrkxM3dSrQyoPKgMjk6dsGgsLwD3MJpKQZNF+QNosh6zHdSy1ZvEh5sP
E9OYWUEq07hVxqdVdM2nD08/V1L5xR+tx1SfGU2zD1s3hhv2TZI61x5at6y34ESnk104JDEl5WDa
KyUYc4cB50APjZSTkxVbHXgjuJlF1+QcHRffI1czc9TNFm1XDVA6XbzP/HmQ+6WHgif4CvIdUI8U
hBqD/ZFeKG6qy+tJqw4eoANcULeZQrt1yLd2hqWqxdNT467gX19nDk/Agd9dbNKqj5qqkJFGnMGK
/FJjpo66Xev3Wrr/6jOM1AumXBFTo8mZjxqYpfDFV9SUVMCmjBofQp0WnP5uE6DXsE4NvsKyHtSJ
K+Z+SkM5m/M9xO9TfUS9gV4Z6loH5+5Oy0RFfXpg9cp44b0QfJknyWMbdPy/Adhf/ALFYEwsq8GA
M+V9mWponlBLKw833G3Cwcl6vztY3Eqdlytnb91GLgCdN2n3NoLWtdTUMv7o618lxZBkfgo9RqVP
awl/0xH8YfQbelyG/0UY8S3yrtMroba44L7hsU4nPCf+NVW39DDwxNReb5m/9F4kVomUHjaULbdR
kPNZPrpA5co+0bh2a/5Or966LTo+GHyeY7wmcHdEpq9t8+xo6bJZmADBYkMijD5ATBoPOHyqEVJ9
Ws+iaK2ha6HV3YwLRiwAlaRraJfxAziraVdPQOPY7+clRSqawp1hPSJFeSt7g2AWQ7LF/SHrUeay
R4gQC4neFLTg5VvbxwOfXzFGYawQYi4m3gHVOTeYISIZQqrjCemqy3WJHIwqGMp28dqby2082OiW
Ru2gR5IuQxLcU6MQX7Q+T8sNXWRHLuY/mZMPcN86D6R+TTDWYicdVp+jpxF/bOWhucgMU4Bu+moM
bdLqVpLlxUR/4eDXxdjzYuTAm2MRRp61BjDvs9KIcC/DNf8oOk5eEVU5s/Xdmz6raIB15SQHZM9s
BwsLJi0V1w8nnuWWTfsSFkG6tvgQhMEAJzLg09ApDW35txHEhdF9JWRan1va6Et/we/fRYs5QF28
eA7Jr3ISZ63fpwiqvZAVTkerKQq7hcvAc/WwoYMNSqYAjsz8SzxEZq18/GAw+GPgV1ZEK6ALuQaf
5KIxI9nqjsE8RGaH7KQtSsyjAP9SxlB0asbVAocCdrJ6sfRMWk0hmtVotad40xJqrcBNYDiiFoNv
iQD8eYPXporZMLv9+JfbjbHAWcoszXlIUEY/V26YhNe8FA6Fms/Jsmv8zSD/QRP9I6r2YoDrCjlI
dMSqFSa3+dDZOA+eQsTDC2FiY9wZ6LkNV4VIKnOz6IegM8GLtnh94tErQsBLeOUzPgSq/oEGNXlh
v9nqC1BHi8fYXZwsaonAR4n6t5H5XqLiRhgn/YgDXx4aWNZF6G9bIB+gXIDMnvASywvPdFHH2+ih
4gAN20pd2oa7E3ThL1ul9h34UgyMB/82J+ULSfWNe//eQqtRGzGuqbizaok9cuO72EjOVzPBTZ2f
ims9/CGRctJHz1UqoiJonz6lSJSWsMSB3XUs7phnszHsf26puQ6Fxv3vewDbuyv8T1eTicbDRMq0
BAfhfEQhp7/TVyCGlSQ3YupOxnYMW77qrVQz7DXEMRfRtHtXqQckrG7qFQXMFiaORJWzz0sFFGeC
NPpDffewRQVkEuLgC7BFAmb2SxhPvt7qjd8a1K7oR+a27Suum9WBw5a5qAZsnhnM/8bJDj27Pjir
dDqR8sMFNKCeV1Mr1gPJj9pcQts5yXZIuIDb/Y3zG1+XYO3hSqdSqviK/AQbhz6A6sEaXqKPrltQ
7egbR7MXsDu8yPdfESCwiPgHPtxXaUH21SWBt2vtwC+DpEA+uybipsRBW+ePpDLFngmkowNrsnPe
wsv+2IzjfSkEMU4sgK2balrgDwFZyJMUs4VxanQIR0Kw/f7Jys0FO7Vbxbz7hv+u3sihqfvHrWSr
xmg/8v0IkTtKDLFlPxCyEI64NGR7cmSNQtK3aqTet+8E0k+j8NpGtm0RMtXbche/wSMpYHjPmCkv
JoR69iP/Q0qjR/P0HCJxSvk5dm6kYOSNTJEeI6pvBYE5nuWl6WKkGhDBZaKrLkIMEt036zQT1jdN
BUfMquL6YF8zNmsndw5C6OeAbawhYm2ynrNEaZm0MB+pkLZvhEmrCVTbzA6unfUvR6p0PIPCkeC/
q6YGvX5Xay3Yx4+xE6DwzKwD7yX135DNAbdD7SpwlPcOPPIrP1YOF/F5gbDMbiPGIVn8dw+UC7Um
pZx4KBao27TF/e+aVHmOcydgBehlen7kjm1uCHlatjTdxvjJUQNq95SupBoKpRGPa42MG3/HSuvd
Va/6h0zFn8T6scKztUcWVaUXKoJ2qIiUv6LV7D+/AkGCzbS1H4L3Klfghor9bIdoYJL8IdYK+5gN
VJ3Ze6nSabqKeG7gLwhIHaYATwm+Vrzt69btLPjNei/0VIetN2f5YEaZE50jaCyTET+a/6rwUYRj
VmOMMYPFCfLKMjvF9pz3QqYMJ04TOzfc4aoTVkcVvLMsLKpGrzt0djj//RM1MrbMwcHSl8nQtaaQ
ZLXwKXaKbZq5e1pwzsArycAfH0H/d3JuMuCQOs+aFFtktDVZmHOXRZeptfeyfd1S3TPLFODxeb5O
7qCct6cD+ZkdxHLEufDJi9A2zfPPy9sTUybcvMv6NSpLvOIiDSJIKJKQgsDNcY+Hdpjrj4FHtFQn
mYvk16aD9KHbcEd8ej8Zb9eyy7FURAkDX/jtVdhYBT4fcbJ/AKnF/rvN9ucLF8Npwj02/mH6zBBB
EltdfIC6JZ8kkW1Gz/3zJ1CHkxYjRYdCfZ/K7XZRH2Z0Vpx/Lkq+4kQeSasBnJoRaf5Io9Y+Ke0t
QK+KVpM3j8kcFbkS5dbtKu8vwtAxO7nYjDFhrtgqjVoqtfdUgBhbVIp7Ha8EDFIbI1ck6oxmatLM
FVr36SSuDu5rdRfjvzT3dNoxWGp8uXQ3WHHcqY7+W0NFg95JGCJwZR2vKgUTas+fGd8LgKa/MhTI
2ojvWKqTKD6BbeGKWQwZJvaec9Bd2rP6lZ24vk6BRmQ6MMgqIi/NdynfB2Zyw4mqdr+Hc0qKjUoi
uLg6SfsTkbfDwMertXRCEVLOedCNqqtKEsJHQihR40LvEiugGN+uRTlQQEwKK1UCl3RZg0FKTTCF
l6d9eoCxcTnACTM0hqNe0WlXhP59os+szmEOsyDUFbaGLZ4FeCrr9brbzqmIOw8AHCCH53xu4VMZ
p5hq9A41HMoystPmTlAGgFAipTc1JAz56SnuhPS+5z2lnmBkJIllwuO4DCETWPbjCCAq94SP/6tV
Y0kqTclGOVLBOAE7IFQGgVeZYSMQ09y/rJvrXRLb14KigXSVhIc2RlKZGwGD/qWO+NFj9rUoJp12
ib8S+oCkqjSUdm8Ur8Gs2R6WyGyV1uNaXyIKu1xCA/3xk3YcTItDK3Yo8b7AnLJ1KOlTpGGpKmV4
UYMyl0MO/vcACBldyV4cFuqkaONeMcVpJlQst5yXKQqcRRX+BAAyKzB+EtEsAXdcum2YiAhYY402
UExIerpdrPyoT+mckHSryq2viAzGGkkht9OLxNLSIVklbSHMfjXOCj3NcmVjdG7VzQXeJvo7FmKu
rgir59lIQutTeyEqDRn05gC/4FcddwzG66lYihnaM+QdpDk3Zi+vaHmZZgVwicfgtT6qwij19St1
Gpvaqmo3FE+GXfN215MSdUETxFgjGkn34U2pUCtIl+kGp5+BJXvBuOVRMS1veHaOLYy1AM1hPz1R
cf1Y2IKQPtkn5QU487oddugZUTrMk7VNWg0rZ9aM2VAWasonkavV0f/3rjxmFAe6Sz+D7G1L+KFz
X9Uh/qQ02JY95XWteH+yjatPuWh4Ig4T20Ukr3ml2WvXTKEhYRFa1x/xdIxKxLS3gGcyy2wz7gan
41yi+EGeaSrV+uThYT1Pq4QXsvztCJZNhdi2cHt6WOnVm1hLx6huVpO5SHjcd4PTLRLO0XM6X8N/
RW2xZLl1Ruw0JDA8cV9LUMlUHEvUFwHvdopB3g5oBaLJ/x+o6k2ALW2VQOc0IgPEAVqNToDZZDKR
koM4Ap8pJgBxpFYYSxizJoPMmMVUJjlrbtZ+pb5wCBUcwaP1KDlvlWQ7wGYh0t/b/O95O2EsZrma
SKiPlZgSJgar0X4p+boQJEjwYpgU7IJ1sEyVqS8qv52nsCFOatYASfs8vE+fo0PC76wSs/B6txJm
AQpEwYmxJFws/aUNBWdetjcW6Z4GKJDlJJ01aDHSWdb1LUOtTIKvbGqWk+a5lOhjwiZQNDmqL69e
WoLrPh3jKX9jSax2k0AjjAgPu+14zJGmqPz1vS+jDAhWN0JSfVn1D9Iq9F8LdgYTTp2QpVjow+3K
6FLfi62zjF0YmG8ZSod2dVqjIegEjK809KwQJc+NNoemLPfzzJoQbWj0FaWwIAYz7j7II21FL2EJ
/2x59xx8vpaczaJRtC12EaDD7o/YVT0TuYrt65z0dwEszhB7vyszp0q9xLU9JYJV1IhcSDy0rVm5
7gIbfgKn5McRNGNX6PltWSNZ/Uueifd6yLUjMlRJB5PiTqUNFDV2iCdY5pXaj7DrQg17nGWKtLL5
JEHya0LCDCU6iua4jNW/0eKCqzLuwEaMTA448WkNnuGtJl2MgN/rgSdgk9Xbsp4U14opXeB5yDP1
RFdUy6ol0AsJVjlts60FrWSJEdGG+TPbLIi7c3YuDwMxE6It0fwPpMDbUR+Yz2UqStQeI+J5Fu8v
Ent9qRQ4HPPg8/ScH59R2Ds/JSlNR/r3C6fDKoQ1RDSmqIgJTOWS+J/h2ZulGK5ws9i2LCI0BcoH
F9FJQoUfw3fUaPbOGZh5jPPfLAaG50GPuihFmyBExG5nCKvpppRmysNeaQZSJ3t6NkS/j9RnWVwy
+Fq9Kx2mmUzda0mDT/T4TXSdV6dY5yo87tNKUJndOytDFOWlWk7RVpGX7NrfveJ7MfJPUSvoSz40
3hQukk68FXTM4AvXU2JHzay4lpnrAgVjdnurWvKH0w3JLdhy9awv0LtYWYC58D+PxRrL+IAIDoMz
R53UDF16kGqQMdVkRbbySnDtHO1WMWA2hbpFB6vF0+uQnd+TRvT4hBmgi31wM4H1KCMyFVNtB+gH
2HzC+sfVRx1qhbthS0HKij867WiUXRTUTtALhgOFdX610cjdNppKeah5/KWgGlMvcCHUfn+K5PEF
x0XcYpYFpmmHR4neRgFRx0CTad7vGtFGoOaVexkOI44qDaRbgGr3LgBtGUv0A31y2psvrIBfTzOL
ucqZRf73wEwIQtKhizXq7t8lXfL9CrAe2qC++RW7InMUUkTxHjYOF+xan+VQ74EkvDCAWox+1XZ/
zp/4nWr2xCTyzbjcgwvuKZUtskKTtMGZmj/Kvz4ASexxqZcZ/x1oymbsJG19Sw9F6dwVH06Ej7HY
FpZkGs4VKhPLasWSmQp4j0vVaWRt4FypTM6fsqGFWBJltZm09KyWddh5c6qeEIBdr7jxf+ykp3/h
zgA9VTE6qDOUDed/44O0NT4hyCq3kSBb6afwMxbHtrO/azgYh/x/6YHGsNXsDmthBgIkzrEOzhur
d10y/Cwuzbq6OryqN0v1qKIXZ9rb8QavylZWxTxDd5oBgTsN6r9xREzQBpqDpAC4MyZyFDhe62sd
fU9DD6bqxN5KkGybER+qHUgm0cNBzB7j5NaIJ04OBs0bYiB9G0n+lx/b+oBlRm7vmJ9Gzppjen7Y
oSLKCZC4QaT941KvuhuuQ9YsDOcy9nG0ctOeB98FQupujhCS6Xa7ZYKUJvUN04LGoA18JiKpHzrQ
Tu/nIu1oh9oPpJt6rlfFjvqVdLNmz5Ul4wE5pbNjmzGwBPf60Ood3MztlE+6jBZbAzHQ5lLlmOEM
lcYjBqWacIhxJQQgA51bnGi3+j/YksNPQklbo9OP/XpJvF0qUTAQtZmc4ABzgxP6KR9Dr2UGlWiK
uXQdpEiwL2tm6j1o3nl5FMcLB8B0FkBBe6JC0MEaXz7ls/yt5ggXt6PRJJ8HYK/qO9Mc2OUbzSVD
3NbKEH6RZuz0uS8z7BefGGA/1fIF+ARw/+HsW8VkZvuh8EBqc1pK5qf6kHyUirzK8JcfY1V5KyR3
NhYp6L+ZGAMc42cVLg67nLFCiCtakG0eBPSHzbrSobwOaZHICFLHhPxOmBKWhAACLJ531qZQC48d
tGqlJTYSnyT/Krt+by5nz4Qf4L5EOdiKnfJdfxP1Y018Hq+yBRQIHOdgCs9ytgoKI1r3k1oeP+lF
1Y2Y2qDrSnKXgvX8PtncAX4MQ0ywEPltdKftrsGaILrIaPT4v3x0CdEQKLUMxai0uw84Dqlnv/mb
AAbZga1ug6/hDRdsbrVYcZzHH8P7ceSzyTiUfuG/zEEQRo92ywOD1Vm7mKk9yxDb0tNqWpWRgedh
XGzH4znHeWPL55QzPDXhpF9D8b43vPiUtcEcnVRmuWds6mT4G9YN7l3xk7A6jJsRkk5iDicRPVof
H776uPMETBl/FRSndaZDLVbhEEZ+CX3GMAeX8wD0qZ0OGSIsfyIi7pVKS99nzn2zS7tUrYWt3SIM
Njs431tDmzK2zyRFGe9VD43UM/bDwUZFVaAGA6DtFV8Q6yqSviZQyl4dqe8YyGH2yeuZo4LqNPsp
LXQAYzpt4IV7KrfcN00+jCFzpzRyx7epWGPaU0QiRJ2N0qg7aCwa4d8abNcrFUI90/sGwCn+U7T3
5xJLv4azSWjPRJBWLktLeeyuP+cID2skkU9UBFUJx0OlP0K5ZNI9GOS5BFqJ/DvxJ11UY8+awZan
SqIo4QLQfIyCcdpe1MhJmUmJnscjYVRkUVx/Avqj9WrU3JYUx9HyzKJb2N9u0vbex3ILGg/GxW0T
7iBtdxb8FB1FCrc4IstbvnrvnYNFCBH0dh111giyaYospTKcCS3SyNZjNF0AbGZDgMVr2u4q8eZR
JAq5NKRd+d5m2WMcaDWhixH7fvDAGrYRJlnrjlj0hNkaLm9i7wunUBpEk06yI6erOR57B6SgFi3y
T/wDua7SXpgre48r8bu8Wi/mh9v1BV7VKOvBYJsvhyiEqkpqocgD7kD6sssffFu8YgvrG2A7dgIs
B1oi1bT5krw7DXFbhrY+VaqlMiKK7V9E1tV9lY4nk5q6evokH48wXoNCnJ6Y/kydNaMsfSuq+Zrb
2vt8n1rUDa7KuxbbaeqkbsLIw0JJD8xGYWbT3o7fYypYiD/QkkB3tWCFPVtf943xF57Yz0ZY4hx4
h2TCPVy568VksC3Jo0/cFgif+rnr8hiBLbG95GFc2o61jdI7HQazrcMsJYtp8ePKadBFWdN90lv5
r4WJVhH8KZaKumNn+fgojhJpTHbGRlpdHjoOByfGx90Hwwd7gjuNaqvOFME9fViXD3ukbFCNAfnF
vzMPNl5/wF7AbCVeMMFa7TVUYqZko67r+yCYs0tw/g01+3lhuruzjPf6syPYzDnzLRd0o8zHldoG
A835qPB2cnWT5pkByCyVGp3NIFSx5lyduV3RE4DIO4M0oyiFGO0du5IRg6QEWZJRYvrUK6iIVR6k
nUJKNnfbYnYvhLcivPfevyaz1h38WW8M6SeqQmUuVgDVTAvKEIqR2i+SP/RoDyU8aAYD7Ro/Jba1
1cGa6MavwQ4Iu4mkBtbB3rbfRZRJ47nUO1WJoUjw3MbWbZknZ/cOk7gkA++6+PTt902js7QSvx2H
bPRtlKLRNhACF1vi9L0GEPKnor4A+5Tug/6hnEW00eCGLGkTnBnV27d8R7xkA7HQkvagvtt5yZj1
ztU9ZJqC7oCJoeLCbxCwnKHMKGYqgkP1vvLm3t2+VdVP/wO1j1SpLAtmJ5qX4Hcf4ZShX5ZCfwpH
xEAmx3PJvanTv5cfBu8oU/aw6JdL+FAmO/9jkbbG4gfQM7sYPKrPMvSjZjZwHPPsEol0SqODnJZn
zHwOHBnl8PhMnO83r/DG9tjF2v0pWuEUPXYd2torUCmq6+1AXDlQ89dDbhurztXwXphSjsk+0ErK
eqNQjFzmPrhAAKgcJ1yLhr8m9P3GnEPo2v38faHMtWHrrf9EevU7fW/YpO4bdU78v9BNWffKtzv8
JVhRp6NSPiOmcMdHJwNB+U8CiHledwjKNNf/+qot5SVma2xPMcJPLVddLqfIkCUNp0lrUNFdQ/+P
tS5edp+iBf5OLC9QEJGvsCqwaCRrhgff5E3xmjKaTAFDeFceeXpCGaWwx6oVZ4eWzBC5dv2J5qff
0q0yEk/oOCRQYNx/XIqZHyQv4kU6ZLc8qgll2h0TToDL8btQ5Awr/W1TpK7wThItQblMqK6EeJEj
Ov1dBvk27w7YfFfxP3tnYEzaIyDCVsxck1o+/YFH+urggO3gmvdQ2bQLlhSv1QYi4W8uFyuY/fYr
QRFNXM95lMmtDNlzeJPg31W875i8vzBrVaFqb9KWsPhE8CI5Dmajext2oc6O53V6CjyAUc4ktRpN
2IHdvQ+AouIgWyuPnBq0kmIzPpcIVEh0n0eWXIAHYIb4Ne/C5eE6uxtUXQS2bXPMc1m4R7rlo/y8
OLo3y79pUoALppX/nSdoqpVo27fTn9ZqsbX1+eUY+RmOheAYK97c3E14YYjh39ABlK+0ZkAY1tg6
et3pXKsXSsGY9nf8I4Z8ceqoaUEWczj3+8YQ3uaGZk8AzmoHDuDtJhL4BumW9bk37xsRW35/VKgN
NAIrQ+tTUMJz/xmqaVQIbRW/05lKeTPVOcv4j0xE+b+zJtvSj6VWLuVOxRkyqisGAwPmSkQZkSpw
x0OSqP5k5BZUW59aU0GVXm1x3gqwlfzTKbpiB5AJmnXMxanqBDl5iVLijhbxeY6tjJCZ/RwNCWZq
4Eh36S8AU59fpQONWfK2ijvnoTGs2ZcmwpWSRgA/BaaD2qicQkTaREnp39U+WNN0rLeRVoW1zln5
6iDX/OrcOHNlin2g5VGUK/54mFKA9OubexhirstbtulOB0z7GRSnPLH6rrY74RY5rNluud/QTuYB
MaXcGaxJRDwwRjY7Z/CN7KKhrvisYaJInPJ5HeMPouKBTcSbXmL7iaXlVDb4JFNssP0qVPdUwzwB
FQWopnnt+ySeN5wSkXEn5asgs10TqnTuI6fesqS0M0+uaCJ1RkO1bRYZgy++J4Ukr41Xh53SMd3N
3FinaXWD7mFGdGc8N8SoC8xCWw5+TCwAjUsLfCjn7+xqMGUK4sUTbX4Iyw9nwc6gzp601ar5TbIW
kdGwwxXTG/BQ50mK5zsjFD5btSzhbztAyIc2JjMx9Ie5+RO+UEZb4ot1lx5adTMaN829vzSEyRqM
cHaBZU0bPTCjpX2+2fWkXG76JJ5i9RecdqOBAK+jqzuziuF+WXGBXZfLhV3J0RkbQCAbeAKxphtL
KzYBETT2VQlLMlDKCtjoVyYPkwci78Bq/Nvj9re4xcG4MP9bTBSsMMpl6IKehfEif4M5FvpFDwOP
7pgjy5Twc/lTF5PuoaCy+5Emr/H++XfJOQBug5i+bVbLxFFGdyX1IpOWBm9MNKuoDJoFOBEB43LI
3R2HY6aIqh9OqVCuyCWFv29qLqj78haAKPxRZZq9G9rNsqGEMliTBbxivJFSmrNFVDMfYlxSlPHj
X/EW35/Oi263e/tV7Gwg/a6q+MzipoPJoxFRDugwAQT8V32DVcNP5+zGAanbF5JzR/Y8Z+pMNeoi
9Cvy0/Na0Vlci3StBO/NS/SMOk3Ya32cw1NJIiSVA5IFiolugWpUcurdXro7ZnTTtfZ8Sk/vfSDE
uvRLLhND8iMmCKPdGksD1SZwCmyqZ8pWbbgv6YCCzNxSdobxt9i2W2V9alCHCgm944rhlrBoDjNT
ldv0LmNP9gKDsMvoGPQoUfBDX790hUB+7FXl8zysQOECFoWezBNOoZgFCGBo7pWGCFdswiz7uyC+
qUR88/qLZrJLEf8LbZQLyS3obBPvoap2/0ZmGAuzD/PJHG9r9RVU62AmgsRnlJ+b8EPq2JA4BdJW
aHqqdQ5hlFtmnB3gzEM5zGHNytVLrmEUbMtNDENtEK1WYmCIp8GBtS5m47CZfa2PmgMnlenpSmta
Vu9dQ4aSQY93QAobGb5zfxaEYsgd2FK33rhCqRsEnNLaVwoIwDncuYaEVJcdm2oaA2fyLePAC13t
hxABigT4tABKBw3zvlDSvj4KJ/dY8DYPWcJJeDuc5QFCSbXcNEDrs9FJ7b70ErqmX9YZLfdXL5j6
ED3XWy1xZV6cnOuGlCNILK1jQ1s363tIGMu+yTskS+VikCB/No27AnbLpziY/A6he1FrH/2ZgPr+
ZYCNz6Qvo5nZXygjpfvIhCaqGkmLMk8IRDScsWpTw/XIwK07ZOGvBOjpmaj6+a1xt6+oHyWy0LIg
tOmN/nXlbxZQfLPJuM/9EaDUSiOp5r2wRT1eOWwsTqWtm6XYBo1p/gKWDNhjJgBzez477iFsIbVg
wuey0jIiM5X+t6lv95E2edjVUU8OvMM7ZNAlA5tdsvTBmKKu7ytIktZTnStRu0IobBY562qvtevY
w7l/jAkukmF2FzuzHnM0UgMj6TUdwnGcfupENtLf0qYY78I6ulYjjoJSenWEENOCveqp8DxPiTAg
Yen3fQS15flZuNLbrKZiFvlksP8Zu2qaSJJ/sV0oS52IXuSjXQEw0ugmB/43orkxvRcrx4q5s7lT
mL55etapQ0b4lh/XrpL/hVit/VI/veBkCfelBC/JbCbGZPC6Tj3OzFn3SMrvQReal9upj8no1vi1
wy4FQkL6PMySifS3aYvg6wknCHfn5O6nvcJdCmL9AarKQsfS1IzuNj1ujGhjcGdeX7t7fz7yyRkX
qrw+rW4uqd4nBKQDWp1dKuPBJmQ90roI9k0/5efA/ODfiVZn2nusNAfkhiqKxBhSus/u/k8i6pR0
NMwWNcO2pG9Kamt9dYFU4zwLDvFONOPhWG00hwez1kJEOO/JrIWWrOUrzx8q//Hjch4peHHpBFsy
xhH8f2seTdduAj/Bl8qgNzzFqEHrYSGs+dBaGCRvprPR/O+Mn8e1UCTSm1Rn4anG4rSxtSvxUNEs
nCUTYzaNa/mwLUv4ZCA1x9sUiJkJffqSugmtkEPv3D2UImVI68vgZbkTfion3mpFCAo/pKBVq4vc
32/uFUqVhdmWM6i4oTILK/0Y84QoRd4V8O5yz5C0SOXfQ/fjIlJszxhKVSDcnVXtTxR34Vpkdp7U
BCFPpvoivQB5/JId0m43+obuBAPBDPHb0r+d5YrCOZNItRwHXu+OyeUkVUqAqc0Ica4H3PbpnDRY
rW25WqKvJXf6EIO4x/VxuLiIgE482lQRvDo73byn8bmY1OL1tbJYXLsv3JIUDPbbq5G/qOkCJO57
uOkRQIC87OQTf467/oERLOc0aDMA7sqFo6wJwG7cORcnEoVKUiNkqCWOfAduFelM7AfAPHpnV2Sg
3lSFsuvzTZatynbe5L8APc5DAcuSR2Bh8dGimAPWpVYs9IIjLzUk3t+dvmQ3vziWVW5poV3aTqRS
E4qqawUO08G4iOY8fpdmxI2nk/k6o4kByjYBJqMOzA59LJuol7bozWyEu2sWQ1sPAvW1I8nZG2DK
ZaiZIlbnUgDIc/gUJnSjw1Y28iMj30hN8nQD/VvwQBykSc74J6vz6KckzRUnh0MLcJNZu83sAGnl
sgJrmZLANfpOhV4EDCKEyPK4GIX7kUEQKC1Z8sVb9SC2+oRaR5pceqBzV3siStHi30T3b36ZuzKb
J4g+IspQd+sQl38Fanjl5KiwR8pxh6JnBc6BED1maPnFd6aWShbMKuM1i1ER+mELg5duarqQNvqu
wDoSPvtFIA5082G/pprosPXlaOkAQqMNcd9yy8OhHpBtSorQ1ZcNir7SQSPPzjhs+1ca7QgKVze1
7qj3vU1dDvxFo+Cv+LuLeY5z9ZiSSeVjyCOd5+aXCOTojqVDQ0Inm7rgKC8DUYcMf9kMl2n3xHUH
MK4okt4bkKkPC7GmndtcjhrnEn2FGMNWl6ZGU7ooH0wVy36nFyYEst8oUphqhnpRiO1ba9fSG4rU
jLm03xpRkyJxiRseKISunfWn+0JusLCri63xjNkZlDN84A/ZTib6Ktrg0IYEZ+GFE2MIyHX6uOlu
mNa39ugMpzAb0FGekEdWImIPP0wdLw46w2rsiOENwXknc8GdM0g/qr6mDhCQVc8Kz6ovB0gsNBSq
ZSUj6GbRTX93ELGvYjijdp6OWVEcKPZj48NZgLVF96d/PMWB8wemPtxxursWzViePHp81mCryvkG
KM4cYnXXeniEw1Lqop+AMtQFx2GW3o5hW/K1G33qQn18fZxYk8pdaZtd+GkJN0abgv8URWJewt6x
R1jMm3pAk2tZGrfFn9GwJcENTU3/yThqGdvEG9Q2FbPhHVF9RPzEx/A7ukGW5tQkeIAsYNrOt2ck
PrxsKI47TRSATW5aJaVvdRd5IR2urwBtzYAfPx+jBNRZq3hseMEgtWvtxdqBaYlQEEciK+f+DgxU
QvIHdGBtOZtyi3dvQz+UOwMZAyfC+sNQh+6IlU9ngBcyR7Bi6NcuR+uUmGGgqj5POedm005/2rMD
346S4GczxuRL+qcplDTnN454dy4QLUWzaBPAQAPKqCyqmF/ge1yloJWUA7dpLyw3OKf/RMRuAYT4
vQLRGN99XdtM01H+pp4GglbWxfGuDalZ+1FeA3zFg2Vt8+OG+IHpqieuPN8ee0dYlGGzE0GZcrmz
XaHKrknJbelridbI75FDRSqQhAusTGZPzE/v0O38ULmvoqmJfvNC7sTC1EONAgWgDWJ5SZh6jtpi
U5NN4LXUKZI39xdCJdTU0hSYWxWxEi44o8SvjJoHH7Mqp2GZ9Tr9tbtemUIN6seAgaRjVqqQegUW
AHqjHvm8G1JpyOLpfnhp4VrkO6V4zxfTSb6P5pq5Qws0UfKKrlWyv1TO6qQmiieT4mkzGfzcDx5Y
2Ofpc8xY7ZfZ1W9SADOIa9v7tnTSss4db+gvxkHp2XHIBQcdpy6/t4aErHms5eNFQpgTfxiZAYHT
ilirqxqNDJAHbxIHzFx12aXKuk9Eepa/+jxPbkS9sufHuobDjvmfbB0cVty+kWupYI7SxmEEluUI
dZEoS+wO+TJUhQjWOTidGoY8hnGPwYcpwuESsmr6UGtvt7q+Q+fAA4V6akI64zY36dAp0DJnT4dU
WrrjceidkGAreZ0mVcq/Ws2ERkkLAHMzbefE5I3ndrz4M9fWd9gU/irMbc+Y0LAmff1F6siBCJvY
djdqxe6t2WqfWCuDgeQEN02w89VQhqz6ezhmDqnYSIr4syGTLlgP0SGabk1CTOCkQ9xhKgtz6Ozo
tBPLA76mUlVsAFJkKdtxwHNOEqQ1Drszmo/777MT4/EK1cuD1fQOC/uhQzmfKr2PbXyXCI2Dy7US
l0T7C1j+c0yUrtgC05yXoj/GKqsGRGmhrnJlFIot5WnujNwNRgC/+fem8ioaw+jfJjAC46f0Wupn
QPo7ogBE8DLONIiK6hgwbAGntF18h98+z/quVBdkTLDMIzkjCC6pCvNlG55dheokX05j5ZvBnOJC
UPCdoDcH0T8KqwIWw6w/kA7SJBHqn2+n9bWqWcU2LEhMqt5rso89IAxtQjymRk44b5ZxgbFjTD8l
W+kVuYxZ7vzsym2ZznUzuMgFeFH05l6Ik0IjjQXkefq4Y2+BOoolMUNOvzMo6eJd1PeKxxkGlcKC
3shfcVyRc2RC6gVxwxVAK4gcNMso2mtQzhALSVK9tfS/TjecqktBMaOREJP7YZPEXnQZUGUT7El6
9FM7DfGbG10LEEvjLI81LOsKwepQJshFZlXNSLm2aJdjeUHgJuK8Q1jMM8SpCOC2zSo6QTuSeea6
Nx4e/xyghDNJpNfRI0kFAzagu1yDMvfj0wFAevAigFqk+gVNLy4oVMp2eTbACGhY75LxnHrBlwuS
qrwh3ZGYvD/R5XQbCZufOtVxWweNS62s/91W+EvgfYXlCKoGSWzbPE6PuJWzP8kjd4w2a2QqGB9j
O6vYeVq/NpEh2Axu47YMOoS7uZLxWmb1u4H8xBmTH6I+oxGK84pnoUxIdFbwPedxyF1HNHt1qOzx
DQTyhpc+Gq8MGigC7MRyCNIacDOUZX65+Q+NCtdfnz1DgtZGXGyhWfXe8JxEI2qf+jxTzmpR49Xk
wShCg4imJKwgUP8NypT/snNNiGj15HoZv4Wrl8zwn6nD7igccTVjsgcKz8Km4Pn0kV3iJPEGyiyE
wMXpAjEYJoxZNqMWep4Ggwbe85H41erWDF8x7Hk/bzb0JUH+4/cBajZ/ayjST1IjqLt6FlUtbxxH
EdzeQW6D+VARJEWTi9mqCWiMpjYa6RAi0oydediClBxuCMSzi3HEC4j7FH252LtMSgSfP3i1MMLq
9JCt7AsBRF8djApWGqazLYXUU2rcNQSEmbcc5P8r/ARbNYbNg7nqSjs6KD3rePbxVrLYUeOu0+UL
qVVfeAQplqX6+HFIsKgmFe2XQlW/6OUFxnU93QP6NkO+PoqfuXMII6dwbeopyxvntUMtnX2IzkwZ
LfTLFOQDVVFAu5RwR6Spo9iUs3rC6CNwF2aNX9jd4iIwT4DGLp8PDaXEVnA5FMEBQg8HxQ7t8b/B
04GV1oxFUXiA3YX53gzTEvPLwWTneLz29TBLo54ZQ1XouCBxsjCKG/GE4ic2lRnUDO61bM1ftbww
q08v7/7ew0ReUYTOp0yiO1AFwiSsBIC2NgLAmS1eVGxc/L6q2E54gVkjR4nYCPUepv4DkTxlruYz
sbQlhlpKf4HFXivHdpF66Mi6miXAShVgUIMY8xTr/P2CJTPfHLL3OOzEnw/bHQAqN+jsoYYmiqcw
RPMIVRDdLmnuObJYoZOqGYgPy1in4Ursk4u1nvqljI2lXLsOXO/Y5aN7bRcwpu7Od/2IOKrChn93
8Y+PVlHEsUjvVApCFVNqAiH0Wfrl6xSwmS9SYg3u+xO1Ol2p3Zbzw2dgLSbJxk8S/CbB5QFEvyVo
v63luIjyj3E/EI4jOG5licgx97R3gU4WTidBLZk5YXkW4HJobZ+JVA6XV5UnkrPBVGSsxbMg5kPk
ZouHykep9x4dhU9WHPlNSKEliN9JAvnALgz0m5MhlYYtthzOGcdYbZKMw2NFtADXfgNe5PYVDy8q
jfLlotsgJXbaI0st9yoJbrMA0CvHgqTb6nPWevYvL9A3iJMqAHJeSSc4nSQ+BHUBoX7b0mlyO2Yk
VSLCwMAjIbcMGXJSEtzcRRmg11jdRMs0nRVHh9m3V6QRT9t5TCo4wCo9nCl4pyJWJz3kUhcyOY6z
QCCSFHbrNYTDwv8kx11KPBzZHluUatrYgtqeYdjdR9+ZcalOMgSXQwCdqNMpp8nEZOpW9Je7GDBj
7jTyir/72nJjKoOmuMbbTilUgqYzvP2babj9u87u6lkBeknNkKGdU3U+mX0nD5eKz9LECwCpZZ/z
a4PiNPkjkRlJYWYFtvMgxQuYymlDtnCxJVoqhtbj0k7tsOIhNfLhK8TJ8Mr8HgXTbkAtoukjoMaS
0hAinvwD4l6JzSUKgZ78M6aQBWVX2eX5gdAa+fv96R7AOF6d8CYBIFqkBBZl3c92QeAytJuGCTJV
4hvjGbmZYE4vt6mJpq2p4mUpvrmfxISyAjPOBGFjnzBpwtMjBIW4J7GUgSWtzjl/yOm0Yo0WLEJE
VD1g5BdVzZXJL9rUvqFs6M8k/t3hRNY5scsfQgM47rDG+AboyUuHZ1vZS7YJHqpr5PGQOzxN4sp7
av3diCQIZH/ZEfBzZE6R1ORQ5xdlH26rP/niCfS0t2E3HzywnLQhrgns6gcyvpcNxaAZhmN2i8l1
CNKamYlX2/nmfi9+Hr+7cfBuUFqQKj5Q4FvqmsLp7wmE3qOEtojmnO15T+CdgwEZwIGDOFa4tGsf
qJKhCVG8iQbLjvI+L3fbcIvxsx/o5QcajN0SJS5ojsynKLGSA4EuHYMY5SAz5M3fvivwWzolrdjy
LscuKwtAkNu6ln6CixiGRI87q9pCkjLosUnGqPWP3xlE28OAPsW8Urf+LQA4Ztc9NPYHo/iqilkM
/JrRxVY/RiySy4HxizqRpx4SlOuW18DWkQ9PBvTv8l0PpeywMZ93HOGKbeGvojgDDYvMmCHtA8UW
76RZofjb4GIRfOzz4ZgjFER8VsM6OlppcHKl0dHSj2+aO141qFwXIxXR5j2ycrb3McTOCABsVFxj
nMu5SO6xijHEStCAdUMSL4liNt78NhnL29yiQ2XW4toxvQXxLywa2YSWwnQYCCY7SlpH0v9F/Mkh
rXNFJ6SIdwyfX5PVen+xr0ePXdGOhouVR5SVwXrt9NGSOVKzXWB9mu/aOAqW6Q8et7jInFlzNYB0
vN1VKqee5XbgjPSnkc/PY7Ooo0C2ZXzKGNS5vz//7oCzS9mygAjfzHq3UgIhnxJqfANdN1yotiaQ
xmWcs/wUrOecmRAO/k+19YG5V8dgsq6mopne3D+1RGlrD7VQLw6brnN95a+9z60rcP97rLihdd5R
sIwwyA+sclXkCjyFiU0L9wL8wsBB+H5ILnkvsHP1CkLo3QBNn++vUC/+P6ORbdcv3nzBT3QyZ5EK
lT3U7/5pfGBtsLZu43myRTG0U5bvYEbliqfWsQn0dZOAZBrTkYPGKsqPMmypUKKJEvyvnzqVWG9d
lg3rzCVurjrqcGozUhhqAscY5klChg6ibBxGMWvp5lVrmmfAdyEMes54zZ3OtAk8ZJ3QFFAcFjzX
j3XYVM/TJMRXFdD2EMLKLL6wuPeaHr3bpiHt0baZMf9e5FiOrbC2UwAAqM9YFP5xyv86VjNEIEE+
U1U7JkuIE/RCmgvNf5TVCYKYKgdMhQy9qb+RgBIdzB7i0bT1STG8htvOfNNeqfLUljcj6bC+RxkP
4ibzm1ELVrol3vooQniC6LwzFVUJHrCRnHlXYoh3ttRrFKmidq9CJejp0vbjBDLKZ32iDL1CT2rJ
omCnqrFiyGjs2gEjPYj5Ev9gt1NoueDSO+DBDAq4Cruq/quUfSNHevaJ3ud7cD1u87t3u3O7t3St
ooH2N468n0hgHy1OkmMwrve4EEBXduzS7Yl5CqfUtLPpbZ8Z1PRW3vfvXlDG3sXF1WR0V510Q/yj
T9nMui94zrIzsI3sLE9JL2GwYzKZ6Mnz9qhz0c6m/LxxBac5mfNLMRjoIkkVGcZ2XYMoVi3KFRjT
6GEM1FJbY35SfDwh2p7qm10i67PFNrrzA7qddN4iOFvoYUtSCRsfSylej/Ef2NCjyRyT75ia27KV
iguqX2rgax+YxVxkqNQ9ewEOODIRU8n4q3E4onYwsjpp/ijZmJjFs54bOtIg7XTOFka/Txb9xes6
Fev/plOGfdx/OZLAyOntTMAt3a0Aulcfnhg4GMk6TxD3kXDMTrsiGX/dqvZBRexxEQQPiN7s4V48
AIcRFmeRB7dQ5gu5363C4nrtDlcZ3k1uzU+a6P8HwRzK/0T0ZzyDw3vOr9zQCQJ+5CM72GIQwDBS
5KyWfuURwTQcKeO9a2Td0u/djUdP3SX7CJ04S2lXWriWlK4oHXO2CRol6+wBrYI4Pt8h387L+mu4
XWDX/GKdwduW2v0mkYAKfe+Ndf06+wN8YNZOOFLfpB8TJDsqePWBJxA3ZX8G7toNEFLEjlInivpc
TWWy2Eu6Ww8sz4/tDoHqN4C0o4Eohx879Lyz+nqP1L5fptOA8cHzl0ttOEXppOZQoRsa8ZM2CExu
PEm2NrPQWCzMdEZS4U6kZm+LVLtd3Av//mlTPe7ROUC6kiVfGCGTFalpqYo1nRkBLGwcBDBT19L8
5Pa2p94pwvmYbe/EEdIrnjjERYDhmimbEdqmVNsesDiDg3ykdt83nODjqPjzGReoRw0Z5iJ1IhYi
UA7blZnnyq2p0LZA1xNszcKimEcTFamS4qhT+omymvAXGJCW21B2xPZ9L0FsrNg5ntMAKeyraKDI
V6KLmZTrBSi2kEYiiWWLL5HM9roIwbIPq/QTcbJGVXZhgmQuh9ly2fFFwKOqKTW2BmmNX8Y5mzCX
Gvo+/ZyA+xnKIDcfE5Q2sXt9XShhbbiEMbjikWRFnZvAbzpYHuHsmB1VOwll1Usmgbqmptl7+b1Q
yMr6lox+Dcelcq05mdd5p499j/1EMu3lGWZedyYCZy9JVmOW/KJ+kIuiiq0wqTiqz5RRZJDFLS0k
ALZcNuC8yN1c254xzKYxSGM/4jQXUj2blAHIwLlrI6bK4pz9DrUhsTD47l9r7xEAw8BTQkry2Dt9
BITSxcRbbgjbznVmPzMAShe0vXO14nFMkgopRl6SvUDNehoooIl8RCqnaQptXsYKxXucoALrbdW7
rmrt1xAS9LpSHgUQ1jMo8HTjHakyAKpa7PjiFxjsQG1wmMzJPbQaKaQzIJnKJgDaBUWuGoNr9xK1
gyzN617iLqxJikL4r3vt922dLNPW0mDwrDkU7F7RI5bvM+kzImkGVdPJgtuIb1vwmqu/Ysr3NI3+
wg12Z93kAIX/pOLh6RdRuJ50uRZHQqh7s+yKecgQZbXxBGgE+NbcQexWxLIluS/T0/HAo6MLw+15
9Eyor2EaCmfsBAksjcq60w9dj28u2CScMad8DkljwNOipKABseoHop16EN4jI79ERaGotYOLYUN2
/anzn69j588TlkHD316u3YMNNmi2XAAI8+JZVlGZnRGqPyZoH6LGXmbS4FG3wPLjL3g2WS9EQkGR
y6RFKez0Vx3ciUrsZzXetGcUZbF7Kh5P3lG3l0dVxwvhGAgztKVdz6V4JugHfRkX7ERi/P7Dp2/d
Y/7y6xunI/IW0UGwIPIJKB91XxtoM37dWvTvXX/FkSjgV6r/4nutHLt+oJ6XpsKCdcU+h6EHS6Fu
VHiA3OVfAbpoVAJqfQIcj97YYBfjkN6zbesiwZv5MZjIq+tgeZ73ADZlK1zZZR698QcYiL31lvXb
90cbvkXvK6YQHgcTc6F6QYtRfe1KIvkSD1zOiUXFkN3W6fFe69ZmRAJ9CIxkQ2hsq4X087FDfhmj
9T04u3j+YvgsACMKgN1xntpTNrfbG7QLdX8RIo/a3/DplDXeMtFYlusUgN017RuXi7o8HynRJA9v
P214vb9mwXyoS6IMqWZm5fZW/DseAp6ty2j481BJRFv0ycvBTbz+RAxgsn1XM1HhFi0YDqQVw/Fv
scA8CyXwxIrtOm9MSAdZzFENSwZb5Ov6OKq+i767aDafyF0plDWNsGfieMMn3pXJ/r2uBbxNiKrY
NcnBFrkCa5eHJajI9/IcOJEA2LaiGYRSAvnaurXRZukDnNT+V5GSDyGUNr5SoEK2xrr8W2enc4Fd
Z6PPGmhMdLtnivyNAr5r204RAg9Wp+1Udnj00+STIszMgptjr0Sd/ZwI831rScCMmIipRftQr0Vd
CXwBJtVTZ0HY6I9pfBmN/tkT5r2Jxd8Y0Ce2JKJjqzABxnp6sfQT+P6n1KBDe8zJ81FWTLhv0N3D
HOV7Q2QYWK+TEn/hdZn8uz34Y4rGvG34MmyiNgsF0QCe/OHu252Lp0rWj2IloTXvzaUHRsLhbXqy
lIMGFvlVf/jqRHABjZEyr74JT6V3w7WK7zSTQlzugCino7fmgiulqw2cN+O6p/bXVtGalQT5jUYs
C3e4i7v52fS/EHeXa0E72AxbXFn0EBHD68npOJPuRwkXB1+4s46TVHrsBSCooUEj67X6TuAzf3ox
Lws3YdZnLxVHV1iBLi3PRnYBkONXxghiMUfIpLR4IWOTmxjI07/BQ+Svbo6qLD7SZSVy3CodGs9S
Cg0Tb3xJ6AZmn8o3ZiK02OY+b7kHk4wme1WR7vFVSdyJdYs5jLttK8csutIVBBnuFz2SJJ08QSm/
E3rdv3OINRWAfYTTyv7lTN3OEVqkl4O7RCs5+UGKi6qne7BvfArVXSGE5nSnVWRdeXEesMnwyZwp
AOfiWXXrWgKHBpx9JjgW9/EBdy3HXjVXvvMRENBdIA1fbAMKM0Dl9V+xAAI6FNvOIJjciuCwtiIS
bx0P//IzRetduWIHJ50ZS57Sp4PdL9UjUQeX1ExLDrqdY+h6MfxtZmz3qW7unnMUZYnHYYyd9tYl
fba3HvehLk3lyMzba3Vgvy791QIO7n87xMUKmAIkDI6prI7gF4dwpvHJJ9M0nuZg8uonu4TqaAl5
VrjVhiyCAl1I0h5lQmjI+eEuh59cL9URy/1hsf7ChiGsl/LGYB3HCjSKvPq+BSKYXI70nUBsGyGB
Dcyut3dWlyjqWZdfrO+bl0PetWV0G62mOjk0p1WodKCRSjsYfceyGs1dIRresyKVAqLmyFs9iNeH
G5Wa/fEUX9MsGjmBonB5lTYtuYsjKcV6ySeePi0MR62SNgxHGIbh7ivwkjJrSCpDE0qUpQBhlB8L
EtTllZkSaXhGDXrmJjtMTyU1lyk3R3Uad6fK6FyozshN2mpCHYdBGisZ4cwRiZ3vmaFqPaIeRz0R
qnVrHoVeYKKHvj68NPHwBSEWiHu64jvnstH52NHhpLGSI2k/yaumdc0Co5PUEz2FQKmA8l0ktboV
PWaZdTwnp8S0IGdAW5THUUxWUcySq1/DCrIXJ16Qdegq/SXmEgLj0AiPjW9P0t//Z00Vq4vvsjll
9qWoLu7vBQSRbS09xeYfEhaw0ioDyI6/zYxEb0haqNTBdRsSZ7uXhvZLTCocnptJvzwlHLL9rxWF
iTVwJo5mdM0YbnrJCH8xju3+pJ9ik0wBZHjVxLfLPiDG0bzBkgrB60m3nqVXyVe3ELWsyJ3Jtfph
6WR++TdZ1MfnkzDlEeCOl0VK6jYkNzVcF7QJ/AG1AMhAB4EnnplM9FoV441HzdghJtidnaXvc3ID
MmiKaK8lGhvI3FfKAh2Gc6ScXBsLgXiplnmGejDbBM1zZH83/LaQc4P4c+9yVHiEXrD2vevsjPpj
JKzYbT2PJmO+68RR9BewIFshAnWAQ9n9POKeAN1iEASr6OimcWW11vDJX9Sqq5UZZiYu0WEJtxH3
pL+sfJHPsMa9oycqvztuBn3juEXDiVaSUYLB8/uvY7mdyHoJXdq3KFxojXDTNcS/jT0UQ5PVdxZV
aXWyjRuPircouTadM0n13xKtIPOQ01/b3m0O473USsF+XMAJy3dn6fTg5xFIf1onphPjrJ/a5c0K
V6GXcDZ9PxDtN1C1XntlowXMWxWb4viWMR+ILvyGsYGYNBL9tdzVCoWiJxpZjlm22Js6koZ+Ay09
uycezOAwZNq6AdNzxJpzh3THwgsNl++8ZS6rbWE8ARWjb7hXbnFo32soMx+Xx/9990hhRprqbboM
8FP9HIgbKoIzb7Fch3d4feXV4xjjk/Q3P3aLTcrtTF+WiFG9b/jZMPv8IirhBuNbLx1VHq1NGaOG
ZzD4/q2FmUpdjUoWgeqtk1HUdTUvOkeQ1dMTY7rsMBd3P4HbF2FYNIoTgtH03pOzGVPUuIkSrs6u
Fy62iFS1hYVvONhuZLLgKNLm1oNWuaiTn5HQ7Nu8Foe8WyigAyHLxtJSMkKsGLKQyon93vzipfNp
Zh+4/oj7NzNb1NXwLKOaOG5Zay/ijkwkaGsI2JQnIU7QgpnAvWutPaP8/xGfDLTyzkr2QXjAPK1X
TjZ4tPvB0o8Ysh5rvj5XlglAukX+FbgYHMvxeyM+txRjghrjHyS+GTv+fq8t6d65Pej7QQX8bAXk
gZ5h0tDxOMuu0I1gAGwGTxWZoFuSYuSy1/8ULW1szdWJkdFHAXLbP+WrMY8MZy3Aw957bGRVZ369
X8cUL4HehFda/Ep880QvDDv9yQWQhHKdHsbq/x9fvowxlHZG1pilT01NApZ1zWi2ZEyXjDd4jMDr
etQTfvH5n9hwH1wzlpGD7pHow+qUyyP+kCMqlbU6s/+mxlrEK4f+Tp6e+lPjwZAba9AlPPjRSInL
q2Q4Ciu09/PGLPwruOJHU90hYvS6eAQNoSPxeeX2wvF4Bsl8PcBqIKxtX9tQLsc/gCxbEaCKY2zO
w5IyHzWG+JJINq6QI8JxAqfKo8sbCr6e6NCS+D1n/6BYVrB1emOCdf9115xXVWQJqkFyZJKcQvWt
zjsuNVrNAkhQiWdFjTHpFDGRiYrWHfr68/CI4Yvy9y9CH1NjqS7Hl7YBffiGaQDFMqrn6mlqqd75
t0Ao6RmdQP5t2oPqLDFmD1aYlbdztt+FTwftTHAAcpGIf2li/qzsaEX5h4dmKzgfYpkgqipmQ8Y1
ACZtjvcx3p1e1qF3wasBEIiQRepLPe+ZfNEB0CGnAnBjNqQN10TNBeOvnLn0j+TN6zYAh1++jvnk
wH3l4kzIA1G2DrzyQVIg/AL0nRjEgmm9MM0uRcxSdhB2pXcPIlQKBLcMHtxYCSjwTvYtZ9V7X2Lt
3oeGq4CLsbNOBEE7qe0FBqNRs3a534MBnOL0nAjBAcJqN4STZ2BEekA+rtVI7UJH7+dxmFjBfxF2
ePM9TfmP7rhsGTHH/nGgrslnfpxy349BL9M1FuAGq4zQlp92nMlplaVA36XJFapIbrUE2NTHjIUn
62JV1zi/wXGIG1qWzt00pIYnOUpWV+AKhhaB6REhQkc4V1V4USkpSkygIUN8/goBRZcEUhzfbKtQ
z+qZki9pOO9Pn3xJ4m5t75x0kg/pcZkV9h0LQgMN0DP4zG2MBDqgltgxU02jo7WZa2g1IkTY
`pragma protect end_protected
