// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
horS3RvYVDPpHDMfVmpBDjDr7WmX4JlmHd1bPA+tEJ/EZBY6igGwDAHD9KlH
iAXNnNwk/xj6nQbe8hCG1+MoBKCglEoPcKRaxPf5NIpZy8NtWXH52i2VfMH5
3PGbxQqa1vr4Xt45T45ifyAnxZEVFCY5tveYaQJICwGArm7T5+5sPQUwxQwB
mlUk2SyYTq4judZXaJrCqOQRO+kGaKywBpkVu2C9ECjqP3BIKlNtSrflvhjc
Adzu44vWWAD50aBrnc8OG6hqw/D1Et5KVY1mbFDnPUNxQrmPbwOdUZZfBfzO
XkkjMFpWIO+gsrxSpWH+hNywsoYfqd9bM/87To399w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XtOSvuIDzF+q7RLKMwiHeLuirKZW4UTvGkbpKeK6GBEacoEiTDXubdzjqqSo
OZ+PxJe+oWfZ2Dp2ZJoOWxhNQ6kUU7wi3ztPIIl70L9+KoTm4YMOH737nCGI
hOEC/XEpEsfdApRECivn4Q9rSY2tcBciZcy401ZvJJMCTfrFY671AdHfA1fD
Vh0YoH/f+TfgfBjg299kK6ZbQabZlglxOS/HCi3BruXWvC5nQkTfm8txIwJc
76xJC2rCsxZRHsPw0l9lgec2Dz4eG7+E5i4N0B/yO6ViHzxx1dvYaM5pRJlR
h6bYby47Mqd7/brTUb3Z6ozND2mbo0HcipLcJhuMhQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pR8I2sQZpR2b/Im3Be6TSDzKkGV2JuYMMSntl8lif1PeSolPx2VFX6T5lb06
hSI44CaD8WW5PEh7udOIGV3afN9hpYcKjdn+pd6/en/QPvvMR74eLUUTF974
K+R34Bh397AG/yaw9lfxraj7J3NquUXm91vR+FXhrhCU2fPPM1MrBheLqYAa
xskj6DF/6kbUvoEgrfTfUnAtQZjpYKq3IBtygZ7LJoIVOXWVIuGbFNu+NTfW
nIMCLH9MqJHz3uEzCIyr90VRlDljISsStfb9TuxkLNlzJsqHyRjM7FLnuw+o
syjr+zNSetQsg5k9a45fVSNOcivdQDCSya9Sb8Xxuw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
slTrcinLtsoeteGz00sjemlgQ3XqRYLWjNfdypK//dksoHVDgV99u+BXG+3b
NQtObqj9IDmGmQRBGFUIBwKIhG4WJrMy3EStqYacKdEfW4qOkavE9P7qCLOp
Kb7oUj13JeVHAnBdHEbSPxQgOq284D4rQWfhWjcMGefg7g5XGB8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NKvq9aNAO4s84ad0uccjva6MbNB7aa8iakh52Kko4FKgdhsCXjtYZfFTo66g
M1It/sQsQPbKajDkTgh43NFZ1VftWBB++B+HyA4KL4VnG0k8kqYIqWu8W9Qn
cVsJr7q6qxbzVvlY70VwZ65XGVMYS7Rd+cRWheoMwJ0E7/2GomFYLec2ADHr
Rt2wgADloM8jqXU+DjZyqT2bzSpPbkYdoaUQlqPDeDBVbILpYFKkcELUpafr
qFzcU3uw4OAylrTXbTHo/qrzYL2ApJEJezDZZd8XOfS7sRxhRXOF0iMNrABR
R/+hfmPrc9Qa8El86E63tCBwRdKJImW/TLhF8IG3VoLP0o5gk78XSQMDUoQi
E9ItWERug3rmrxMlpaVqQq6NMmt0TigiDOnIi7+xUeDG87Jm5E3UI6wUC0re
C99NdyQ69aVB1M4kDpxkx719iCFdd36UQb4OxJzll/kxUumm2RBkGjlbAFhn
5Qlql4KcaWGyid95zsGS5Z9v22w2FBpH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DNLvH4pDSaWCeVEEAZqqOmIduf/leO/Uu11Pxog9U5xf1fRXJq2UEBPMHE6d
WVz5ZwMsz+sjSbLAKd/NmyBs5ZSC/T251qFR+cS1NbyJoyJDFzIpzzj33nwN
plFjzmIgdY81M4PLe5C8ZfEBPFO/RllNQFrpvj9w7eCA02IrkwU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ReFjxQqXzG1JG46zxRLMZjxNomRgMoFzWo13qctFIXYKs2lQs+pkED8nPkWA
M238BNiryS5aAti/r32B8ILGq/EXEtMpAzq/S8ZacELUZFUORfgI4Tkkm7wH
03Ssq0GEQuMjpJ61OAyjNitdxOVacFc0imSMVxOpMMnNDhjTxwI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8880)
`pragma protect data_block
AFgysYGhcxgU/pLfQk3nZcfOnoZ9M0sbD6YSN7AVAVJKe+OVZoWr7QNN3cZD
68kPKN2c5hh5BLQDhG0iGJHLkj4ikCZIRMSzeA86jmzYJTnE4mNl9OAzy2Nm
IXbOFEGk5IXk2mutardSU9YA5aei3CKest7+ECuouJdYtzF8SEGTiicer5IE
izz1H/XxQQW2TsOCljguer0R16amwaQXDhPS4q8IF2qcTou+RwgD62tcnGe1
+IG0lX+P+kUy0pUv7Kibe1lq3tT0P15bMN6WJE5LM3lO+1rQkUh+xsYlm5hB
txhshEq1WcN4GUFartgSikVvg74NTWDrrV2Z/GUvdMiJ86cUN0g0NLWt4GXe
1IQcK3U3GU6Pz2HiNR7An3snzL/wiIP8b9EZM8I+fXAmWR2eIaZou5ENIW/K
k2uC7ZOaUIPpYhEEKxIJBfuffT6uo0Sv1O2TnRTw3wykRFs8EJ1TzAQtUMpd
MGfhS1ld8eoZ4hru+p4UYT8UJqngxcgbzZUvo1jlvppHw/gcE8gUzGJYSrc5
SSWldMP4XTZiW2RNGrEJ0WlNJS9YNfmOJagi2LpVofk9Lj6mEOs3TQANjh0X
5N0flrgH0m+aS/GIdMscfW/9yMdyUh9fHTkb1kUUKayX27dKlrEoCZCfk/Bd
oxdICrxt6SH0l/4x2bDg81JcKWu0ke7xZjKqhUaeiZmiGjzdpEKqz9oWDP94
AZ5zsQPqNt8Vh5pqhKDzhxcR/qoB/gnH0x2rzQNoSGZ7ybeUOU7rd+2h542t
m3u2x8C43m5JOPH8YF9HK74QPx3V0QlrjOj7aWazTsoGqTk7DKrdQbE5ate6
myGbCFk1ZiKBb/x91GlRajlJ9l4dHM3MsK2gQ8Ig3oCrcOVqrRk/MkyyFDr8
JjWH/DQPpzi1tGMVJ0rtplfUskFOMseA/5wf05aAE5BwUQb6HkJRi7R/4Doa
TnRTm7KgJTmi0yd9FGN0/UfqMxl70wLVc8Eu2fvRrdiEtRylN+7ynk0ErUe+
zOK0+VT4X/1yGpfcfu93NHKLvuTKjN2IagLeGOpLukKEwWxdpmJXdNgTFGA8
ofx0lqbr7ix2LthhHiVKYP3ciK5st2pBi2wgET6WeN+AO+xaKqcoJcB3Fkcy
FzG9RFgs66gHVJV5h32AJEJjuoeusyGIldK3pLNysrg4MZ/HeZbdOhxAtaJ4
9/CGPq12hyQJQMEOBbwIXw8bhyVp/EpXqOo0HABHjmbnNRkJvZkEkCl24FC5
rXtIvOE+7jDwIHsYN6ceTJUgQx5wezBb9IYsjhVHWWVhVBtnwwsmLhkf0DMl
3vboiVJcR3kjyV3d3Z97TUPJp9pEsaOspjpf43OfwcVX0QBVFd3StWgRWVB+
yehWC3YQaORaD7ZZvZuAhs3eQjL7qfIokXSQnl1QMckuTBsLOFxhadOht20V
DZBzUhq+4Bw30fuutxwaM+jpTSwEP3lXbIGV8PUz4WbmhlAUsJ/cXBFNFYaa
ntt66pFHsgMzOfrt/qmBxyaryz7+nyV2oM1tRMcpxCQ9loj7mshy7jlUfdgm
qI23tUwyiDsSkeKznfPjLGTv2xpoqEAt6BnRtt099LpZuGN3jyL3p16BV5nl
RCmUXI1B/Xtwz5Ot5BLuDQzmK8I72MS3aD15C13Ub75aFoJ9cOwr5mBOXmW9
ieZCFmbtz8wtw5OChibMeM/OrgufANQT/xjYkJ+2bvK6QUXunmkKL1hY4yhC
sX/nDcbjAQmTP43QiFTFXntytzO+O5duA6Xqun7Ul+nxT4htgN97kuDChkce
k0yTZ/FEm5ggW0CA1VOQxQ6+pM0jfG+IgQlRm/CYKU+HnKNghvliuQaIp0DT
bAJzgt5UH0RcqrXOtKQffJ/EVbwn9fP9ZF7NYaLtKGuYsqStGdS2i673y9i3
g8oFoLH12i1KRfMohsnce/jEjVe/2hq7xCsO1+eAy1k2QHAUc/mCpN9rCgSx
7jLz+cu2mbTam0rcChEDWm/k4/LhfqKW5lf+DXH1LUn8VvcfKRnmmjwY1lnn
Su+q8NFg3a9+h3JJF2IjxvYxR5YUWfrFnooFwqDJPfFxNpC1TqbHFB3zL/FW
fNJb3ayOEtT2hZQm+fQp466/6vca+aAnOdNBxWCeu64pYB3AFq2sZwLSSUcC
ZNUMuDOyqgQ9Wj5gAhgArWskKDNmeVd1X0+unBnDxgjub0szbxru5UyMCODx
QE2SYMuq8MuwgO1g05vvK1Sn36246w03Lk+oT4ODcUTQB7nX2908Q/x7kCgb
SwMjS6TeRHPiSqJqTKmYxhsPYidIrmXpXHc9YcX7gsJtZd2d5EX5nOdR8Hsq
eZ+oRo870j5HvGug09Bj9ZODq5PbeMFhowQgcfV3sH+F6Gjk5S/n2h60FcfV
u2Jnf+7Tj+NnioPutsyruAPf5m5NH36/OY9BljbsgivbcUX6dJ9cl2SI2rdk
OoFPHg2muxswiCzkuaWCudbIScKVpLAYJ4gEmWBoiU5XLYz954ksDHf1merY
uMLmQZHkeQEDRJbFHt23UtqUXJIRtdam4TCr9Tk4D/Fpixox1PvasG+ao+/d
qesh51UeaxIyMdSwPnRUac79RLkkLDV2KBRLvJqcjdrL2A/tcPxLmZZMJHFN
8vBcfL/P+fpNmfxNhodV5YTOhprZH7S9d3HJ4Vi8k9BlOe++392sElySC16g
S1YhGel/Y0V3+IXWAWDKClgbqycgVQd5ok+cLKZcVGhSNQ7Ksb4KCFAIEEoD
Q91PQjsJTkIOHFLgFu5fLiXK/NRJ0uFNyCYYYnILnFduLLXwk38+D+HKqdKq
oTC7m5Uofp10xFbWYhNlqcqdMi0fw8S9uc1jzeAikj/PYnHNvbJvVhwP0NSW
3KXa+aWLCAvsxzqCaqTpdNbkwYTU0qSDhxqsBUWZbgHEWZXiufMg2IdCXDxD
T5ZEWtktEInr09zCwOC2uuYcnOXqpD27g+rVnCc9O02xbi9ua/l9cTViQWTr
gh2ljARd+xfid9kTPKvT+M306laNESl8sUMyhCz3BliPa5791HrYoPYzgEd6
I7DeKMr4QpPhOJLR8QVzX7SNCqpQtgFnN5cAhNDha/rzGhcwZd94J7WbIE7b
M0VKSGSgflmZjEPCUXgQGFn3tKeTcdPjjfRNHtFa/Z9jyHkCPMavLidDEgWn
G+sAzkLWmeWimeFIeuQNWqiEaV9E2Oz7LpDhq7iquj7BBT13cNa0OvdoDavo
vTBRtuNVege+LvHk8sqHcgvNrQ5+m8hDXaYHV+ZtK7EKJr5TtT9EhxJYy7d4
UWQaYvx4bynuCi/g9kwQTOGVw7L5tUnqNat35/bWiFgTnMS+xe0HjL0MtbKK
Q8i2nC/q7/gFGEXr1RHHofDBZXRF1vDZjXpUtNNf6tvfNpPEBcwd+Vqfz+ws
nSmbYRJYHZjhrl5VmWxBP2+PTS+RAhtHAi9/nOQ8LsxJMTe4R1zWbHpOgiv/
bibU2lAfUF+I3aH3wUBp/UW34PifAVJ/rkBNzfhKowtfumUG8bHmImEf420q
ey4Ln08lT24/5p2I2WdtbbnShfW9O+rM+Nc2zKaDarkk+018PK+Vzm5DdFHY
abE75NYnMDt2lmI3vEqXJqqMf7rkUZ08hEa5LSjcETC/Vqm/FAmAy8KbGw9T
Yw26Cz44lVYGKuDlo9SLzrOqu13FPZYKA4Ffb67W1/37Bdl/KMRXJ/PKa32I
NTuOI2fIMBZiy14Fq3w3K/6YZhnCABbN7hz3nUE0g/xmrGTcWK+SwbsTV/k3
gUD448MwmS+yud/m63KBbhZ+a27/xRE2O/Y3klKfLmzf/y2V+UIDd79Ody3k
84RKPAKCHrLkjfJebzpZA/wBBU5Hv9Vs78ESAhd56QrVs0KQlyP+ofR4bEi4
SmRAC35TGu1c1PfaJydJ/1TYnRHpnbGhNPIz5mEyXeNrYgSYqHlaukaIfbnr
3AvC3uv3MQOzMBvBhazDfigUwzuC/1ccRhP4RUmhoMCyxEq+EN8fw9Uj7jaY
0AfyH9V0sQZRs1bpz53rBhhDO+2kzOVcXjlCJdC3Z5H37Cl/6LTjc41t3Eac
gS/xj2j0CJ3bLwhos5QHHziutk130xnBTAREJARnLPc8OqlExT6T0cNdeUAo
7tmRjYgOWrdJw2bZgbzJfP9VaUO/bLog+3IQnJfP6RgLUe1YDMz8YFddQmTC
9HMlu53s1dCS3vPadNm2/GBpVFJ6Zby0r/FpGsW+3oJ9o4AsqBWL6R1oLT+H
Fg1nMuyi4nNut9AjEKyIQxY+lPeQqOtI1xRQ/xiq9UxdwdK67nJ4Zy0HooVo
Fiw7Nb2Q5SItcJ/iEoQVzLnqklWB2RDnLCJCDV9n12g1nC0UMa2bjj8OqmAv
ZNMF8X/DV9Ib6MxNSP8HAndeVVHO9jkATht2g96hHOaLzsKgqQdotKZRRFHr
yGEwmCz23+vpzwa7Hkvi2T4WnkSLNpQAatjs6F5emn2nXCe1kxbqM7jYXdAZ
MYGY+/2FLfvjP3MST9pJ22hgh3DiVEJ1ZiElm6zztOj9jixGut5KtDgWncJs
qX8a09w6834XAg6uZ6bj3hzkFJTZ0epP5qRS7PRKcUPB8ny/zLvOw/AnX8xs
DtkmU1q9t8N5nF3wXvx45smSPR/4VDGhwKwYZdUzPBgFVHePE4J+xQDcCm41
MvobBHKc+dV+tmCyRY7Ej4vbsH82xaPHvdO6N+YnrzfAub3OXV5wT7hPJZzs
Sri3tOKSCYmcD7BocaYglnYRt+34M0bwMz5lhImQy1vg3XbUuHroKyxwXBHC
+pA+fbxwgxBrP+zWctYO7dTAfrw9cSD7fNcL2OtBYtpFqr8Ep7DipegWW7B8
QMkvxa/+rRzUl1L04PfU5+Nyug+FbOJmKSm7pcf7DY2eTGseiV8HTxL36yfv
LOWWuppltSs3xgP+89xY14dyTlVPa2k0asQZ629/q7J58tmITdFky+ZOPSrl
Or/XUqeVBdUGX71C+UpoCvv6DHKVIpMoW+kVdOd4IkOnDjXRpnwd6oChYQtq
FnlOw7AoAwGx0/ML2C/YMJ7FU9tB8u8xR5vuUPc9K8CJkTmP1H0pAHxCbzfG
Xz9UUbOaICo/blqX0bSHqoDa3Or5cocq+wlaqmd79FzrdmCI7g6wp4JXD/qv
Q/Kut1Xe8e4t2hglE4GAd+gDN3if86OTA7OPWDkeve2SF6D6JM7Moz4FaoCO
OPx58dBSAnvGDLOiDWN1d2wH3rL4K3nbFj4fH2v7E4DH47v26K30S41Xu7aS
rtyrTkCjJg7axh2Yu1GRJFrJNaPq4FOUt37nDZEZePmg+hOy+uTOVMOFbyP4
Hh371F8arFa5ebIbBlzZuoV0y/DPzGRYVWs0Dk1yrB7ua+xWNDI3xLcvOAKs
g7tN5e2NKVSNMSfzTBADJbdlkahTGJ5I9sgGNdgdw1WhAkZ+5XiT3zDhdShI
cVWARTT13ndqsavNmb58pbxCFx0wl+eyYT2r+8qQgTRD+2BI8dKySUcLJB8l
MfhTyoSMgTHv78I8Og5qP/V1nYEjJFuzeYJdAZATVWXuVMN/AGK0Yw/Lede/
IGVtitxsODkeWJTJ4CbNOy8m6cajS+sClwNcl5UREl3XJPP/6uaKZtvebZBa
wqzuaatqYfU3k+aDgKRfJtKIVGRTxpGJQ+0xL0Yu7wG5eUOca+/yrWD09aOT
m4i9rR+Yp7Tr9FNJWw3WjlKD6ZoWuaTFCh6O1A2v4GjC2gRSqn0H8nyLreVz
FbJx1mlYTYouuNFJL7TYKeruUoLcQJc3Zna2ec+NcRt0yMEZJMvq6ZN+T76G
ncvD9GlHzpHpmJs1hmgCv9ve/mUdH9iWV9Gp1fureeTPSk0AX559KDzD0Y5U
XtrO1yBA0qKF6NU0XXsovedthme1GRN6jI1AV/QTwxUKYDZBap/5N7PgAmy6
lEMIwI/qB6CeF2UNrbJYM/flrJDIG6x6eFL6BJiuSO7nZEcZHV/muSzg7WLA
SJMXfVTswwMeq5XEFiRA+RBFJbj+9Dq1VjOtcJ3brXJOAt96YdXzUEqq8oP5
YIZphQo2hmN072MsH0UJ7TKJ5XbxAGo0eo8gTGkelc3v5lukbMTEvB3h9nvr
euu7fK5mZ6n8jPsiDBY6KucAmAyn8m6trzX4N50q7QF1JNmi8bcEJVl/TEkN
8QLr5oGA+hZAk260YpTTyzgueC10+Ep+VGFG1jDERKy2U+oyJk+0VXXNaarN
V+3I5mJ9gTn4Vq8YUGjsyV5fnX9i0578CZSHPa1txgO/J9mN34BlLt8VzY9n
HRjm7d/KWbsUuh+LXK73wQb0gsw+JyteKn62oS7JY6pxIUfJpMXF3LpxW2dl
gP4yobh5cTN7QF+CgddcWI/HWn3z76UvXkrbE6+UtLSP87Exb9erLviofO7F
ZSOZfmEnz9L7OcGi7tKe1G4KqXpCW4q/PggcmOqRsHjhj/TsROWt6/6ozV8g
yTvyfWmRRoTMIKj2jMR51Y3uprmgS6RXBg6FKnliLIfCTSmc3IrDB0JP/0h9
75Sj3F7mUqRCq/LNQ07IiC+iRdUsNMXfx3povEYvjK2tAkAKepqHBRM0gmvy
YCc3wzgPi/pb8kplHDaYfvIg3O51m7rDuCBOfHTXTZ4XeYcBtKBQexRNTdK4
JZ49fKt0AwuRaWOe3I5xmJAanZO+eQgBFyUzh6eeeJBUvwuUxxS4FMWGTR2R
lPLlStmmmsboXvtiNQXLEt7tz2soWjo5EBacAl9wDbK7AO9eIeCxVK/e9GvN
dXkUP77NaQhU72UNsZjIW6vfPKBi464j3rYJBHF95znuAou5Q3qnsKV470m7
0pni1Ie+dDejwmaC/ZusZNV0uJUMKTcz7QeCXZ2PbHNrXASbSzFgyqFhfbuc
f68fj7wpH0+YXlFJIs3zyHCNC2GxZeHE7G6unUm0vTpvOA+WNyzUGEVcPbMB
Ylt7gx5CTCTpaKS4L3cptzNnLbZIJuVS3OXilWf7kDqDVQvWEbzPmNYZmQGB
woS1mHLXxCfQN6ZK2rOMcuFM7RWUFDem6S6sv9qY5ZQh2Ta9LQ3tL//5ppvN
9jyW3gZZDSMq5bRkTK1E4lnojQ/+KUGPMgtF85S1Gg7kDfKsj5Bb0ds9nKJE
jCP4K4aGDr36lStosqFa2Ag7omWqFfN2O+tsPcnQcHofJVax8GJhPvwCozjM
yJrK5KsYZ7JmXuQOxom8g5uUppDU63cdkGQxElkSe2SwRGDHNiK+uNjbLXz6
wnvSZRKqT5kYKZOKqK+IQLdj1HsShLGRgJCpphqr+lodGdz83ycFp2SCHt6u
eQXRMdynvHi8gJFyYnZ4nRdgXBEx0lhGw58To0FiKbJUUeTeos6cdQig255M
5iJ1b7UXi53LFOLgKHHAkyaEeE8sboc/e3/ZS3/v1dU5fGdPYWdQ2iAW1Xkp
TO+YM3lQgKZo+pJF/c1mof3gqbYHGeU++MnR2smk5ciJnkVWyF+aj/KjnaC4
BFZN9ujNWl8oQRm3uK3SR+96cGOl5lS7c8XFOyFzN5/nOEs6JTKOgNo/vard
fH+PDpFigb0Ej19CC3s17nGl6VXAc7VXRB3RXrQ+56GsNDUs7oSvTfsakPp0
IouiABkk52/ifUrB2JPlRv+zcBfc8YNMWhlHuxUcX7ytptYOZug1N66dyk/7
QOSq4zrilGehlnSqyTUUEUz5SM/nsZ6iWDeI1YTZ4G153tsUO6mLAw+1Djdw
EnpFUWbkONhM846Tuww0IhQ4wiSgTixSgtiSGcW0WVrpEdo/f4AMp183oh8b
3nYv0VcB2RVAnq9/ugMEopJgBoNBzx6lzu5CgG4qSzkazGfKhHo9CnJObFlT
UD9K8U5eNMizilnU4rLMl7qWwFMVI3lcVVvc6O6+zPELCUyklOIZgU1O7D0i
kI/dk4wqqW++5OOXnKCKkaojbqMmj8pcEfAR52T0BCNS8eW+1w8pt3IlO8Ml
nDFaIp6dKKDLOaI9EanRyIworkhy3hE8xdDRbjXANf5xXK07tfcdV0AQHr0J
QnX6EUIPOnkwVV8klEwAw+B8uVUjqmQ2he2m0icb3IpVrMCEeP9npdlbCeFb
YhjYWNgzoc8762sfNXT6VgVZiFn69xxfn5UVGDrMuV9YoitOeymkmj9fLSbS
PSG2IYTyTuwK0mWOG3keaAbCk6+ulsSfH577/pVamNpuvxPkaIRbTxem19BG
u+bVToFoqmULPM14cn+9qzLdW7aJAI0MdYAEj27jTIVOec/eowWBNvX7HJDD
34t6DNciO+Tl2y66ZWY60+te77m2E7dVtSq00OjbaqcFmRZbwne9lEuJvZrJ
YcXOJSGVQ6RTr54TsamjmqDH4lxCLGO7iD0k3phcqdVAoGyegfxa0SAjo/Rw
q+cqs3MLjscxw8vcegwyJX+4wFjeH+6M8VeaLEG3P9PqfOGM4OsWPxhT7DYl
EgVJNX1s+WG6oOPRUD80V71yrcwOkpnU3aQ3ILjFNT/Lb2JKTNlVPfLaqYay
xElEMS39c5zcfWp3TXteVFmH82EeTD5F8Q3R4x0N3znRX5+MiccRv8R1NlxG
L6eWK9sl64eaNj7rurRdABjEvnQ8AD0nhptsXcQ5H39iExx9oA3rJN0c9hOY
Ga4kRdxd1+ZbFHQcI3n65Jp8MTm1QolY+ioHUDwsQZC4pyjrqYTwD9O/lCBS
2jrHwUKKdCl6S/O5ouDlFnTI3PkPdmVHC0p8/zCyZjRsdvHtHi+9mXC2HQfx
B7OCInTm4LkVXhy9pYiJ5pKXkm/WVlq8p3nkQHnFp7EFYM11jZc7lSf9sYWr
3WS5/YoE7rFGKsrSgw8BzbvPKM+7RfUaLNY3KefqCOguG1ii7Y2XvC3qMhfZ
o6f7e8PXWP6TD5OuxbV6UqhzQzQvWiwRBqN5u699aJBOabcms8QGkU9kwcZi
7Uw0A7pkTGxxOm9QZ/1TMwoiMIbL9cdCGv0V8HPi2f9aFxmNEe3EItNfXDxi
Nxe4B4ZZG0qfPxbopdpLO4R2tsyM39YWhwG/JUEMs64pndZ41ouxd4DXcuaL
qe0A9jOUVnnWroysLpLC5k1CS6Oj+x7NUWQGT5/wloJDkNb6IQciXPRE1I0b
UgreMrSJExONQV8dMHA+Xjeu6sMxlxfMXmvSvmeLz5tUIrDoOSC2CzGpZnVB
Nq/oiL8vsdRxBrjUIzCWa5/yCrNkjESCZYY/wi8YtAxrOjS6CWbOgHjr7ocH
aaomG+yOnMjZDNR9xBuwTT9gPGqBK5nUNdup2BVaByjpatfwjvO1YCLlG8Fb
D8my+fHC2yQSaURFM33HevI2EGJMXC8n3sOowOdufuPlZfb/+2R6VpumiWlX
jTtZ2rjndrP6namQxqgobSVLMtxqRkMOMzXZvDJGzScFP9l6fAFD/azOGCKL
IyKLvCUD9ULMvWZJfoIqEuWJnT6bXONBmddrcQvoWqoG0KmSO+2UjTX48P9j
JSrr+7jk31nMpBY/NGDL+lFDLvxoECMvc+7ddhyQgvmd2w3CwzUxd1zB8ixy
Dh/u+N7X7h8bD7RJObS+17jL42NbQ796hpavun283YT42MhBhyfXXvA2XWzP
hRX8xCEEHnl4MghYSM85UHhEHxcR09ZuUObFbCU9BftlLC7lBJo9PWCmk3qp
K0Hq4KuA7x/Px3SigNPhfjlHdDksgwL9bTa//0t0sZ+pv9K6JzwlHXZddBDW
usYNP4Jp36O1zc9ZeUTV2kve9n4UwrT9P9GC1ERzCMDtUfot00h6okhGjgZq
eo+wvygyBhu8ktrk+VIRT8p6dAY919ML80xBgFCXJb6gC9ADcO80dMA+tn11
OSAbEL8TbgBAwNzElFcmOd63Fg0dKQxSmIXXz+Uld08FU0rPXl4FpLlqQlV+
7CF671J1WmrIRpnRm2IVPHjQ+br92ubZg/EnM6ASL4iInZRf1AVRfsKOZeea
40XmmZYTpisD7u7B8mE7oUaAnHpCY9RBIXrJUDTN5W+bC84oEymzo4Y9CgxV
PoGO/XqFk8kc/aOBt+IXW94p1RStF+o4AWjeHl6Q2jCxY2xb77ySg72M3jat
isjbQkZGlQV/GegWqOx0fE3x03ZV7kTlkGRCeI2x0/MqcKnAezX9EjSZuTbo
hSmxI52pi5h0GtZJPzS5mKKHki4IrtoVdEnOPI0C7g0GG1ynE57xII1b/GkO
+HvAazGIqOTL/NnhtptN/7cBnUscpKQLyJAKbuXQ0aeUloNNk2KaQZyejgNQ
QmAn+x6O+4gmkxQ2A7A8SI9snxmLg5HLdSiAhNhUF/87e+aEsg+oRpKmh+hJ
Ww+g+SBWQ+EomP8WLjWaKhnsIEI3wsr59QJuVHLS1C2w1N9Xcw3CBFv0T2in
zVgBk4yh82Mgkl6gDse8x8APAZKyGMO9OqjBcruYpJGMiIug1KJ/exUdvmHk
GS5+lZv3cEPSwMhH4+DkBkgroBeIU/TAT6MWSSASJuxLPCdoRuFhz0Ex5o7l
zA+n0HcLoA53kFUgkHM7azzWXXAo2Rg2GCB6VoSE/GDoS3YN/DdPdgz+taN+
D/cvXmPUstht9jlZzQ7nJV++yVfTS0W1aKtf3KZEjhwJx2AQTf9NSyW3vW9Y
GLj+u/M8A7BqEXkEyqYwNFo2aGCqq3iTLE5jenOm1c0iG2taeti0NBzGDar9
rzqLObhg/JhF6A//MB0qO6bVAgxmcV7BlfofUH9mXR0KG3bGyuiyv+mPDfuu
S21DJ9y11dlHwlB9vWe0zQs4kjhPog9/1ZpBofWCVZV5p/pejbFY4nl+fZt0
oNC7JBlHkDCw5m2fQSgikiRRAwj0giWTDAQb2N/s7gYMUtIqLJBWUHv+xWaP
+RPSbewB6Hj0ShphxGyHZZ0hHYO7j5VyM5m5QHqqCPeB5AP8cmdMPEbrF0Ba
4Q66Mj7nUebobsKJ3IFbHmd1S7IZimGrjLlnwM9UDQD/+UVMsyLY+c/h0eHy
cBFznMfeh7H6tpx3dcvJ4FgqxXkwrGEKOGp2QN4mqMEvxwEPL/eUDp8Fdj0Z
9RoTc6RipbKC0rohX1qc/5sYr9xeD8n1oFwD2wJwK5X5G5nOHuF5iSAPRbC8
kTLFh+ic8gB5InliUoh11MFr/l6au4r0YOyZSzSCMDVi1FHSf5ien9RFAVUf
0OXFdGxbC2fkY1hHetflj6Il+lhUkSyQj1zGY3r/kPLNjZbI0pL4rpSsYPD4
tGt1Lkhfi+7eMjmWXcWRp9/H7VBgABI00xM6q4yLF80vdZ6yQsf8A7vqJnwx
auogJSyxhOZEnhTLHIwvUhrM0eZEbUqCb5VdG540mveoeSuuzQuuoTh3Q0HM
+tGB4BI7r3PvvgLf1XPft1V9Qel3Nx4k1VvX/6AE8/yxO3GZTCGmP6mUVbhp
i+oDMUYavtxIgjx0YxQgeAQpXeH7FD2G5ZEIMJi+wzHRC7ZVtANr0ymYofjM
S/xtTIEjhy9WL0lmrSztqO/NOgbINRw76P+KzLMWE1ZB3PQjZDXE4ZXkeVpZ
3u9YkKakFofY4NHDsUXxcfuEdwarzmF4KdQh0p5mxjXr6wLsuAMaOC5+jNa0
PcpBvyrJghFm+Vzq9AkL4hKz8gceFZ9/Nv17+V7OYwinAvhUfgXQFFgKJGyW
pEdyog7nVY3mczK93ZreONf1RO2tN+mtVx+78eebJNwVygKlP6/ebd1U+Gbd
FLNwrqKztR4+KqZtBTGMOtOQglsdcbXAzDhWg8GA0rSRxXnspuZBVhXT+jWp
uuDhg8kIwQmVRnXiPK2g107DpLJ3AXbJxznrI+QwfnPaEs/T/R5GdsIQ3IAD
V3Ut70Hxr0rzQVGCI2mJ

`pragma protect end_protected
