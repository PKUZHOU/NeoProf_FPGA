// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UVYa+FjBH+Iiou8biNVG7e0ot+n5gqZ7nq0wF5yYrmc98h5vSdnaoaKRQH1h
J39xQefAdVVIAMeZkG1ROk54YMniFdGIjPrifq2tKrkisdFBhIUENHjVbzQG
8De0QaTMbvkRCPK4YvFMOptzCkZFBOF5XcJMLHaRpRKWWj7S84ec5hosP4aU
rcFf2f/xJG6nGMcONlvTCLghC1O5cc7h0HEvauSsUQqI/L3ViLlT3f4bclML
u/BOKdjMZGVzWhl9It69ijviOOHlSR23Au2SrqSCKow6nUAQKKRPOdCz6caS
O7UXzV2vTzlbbEdeDfGGvEEltLfcku/0lj2EHZyf/Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UjNVzNym7xln5wVWi8vZhuLbUEGmZ4QBXUq+gFNCU4lNa9qFWosK85qFbbd5
bocY8bLdddTytgqv22P8hrllgpl7ngKla6Hu+gvouOHE2eSWzJhsWGhFbwuQ
OvpO4XhKhspa9g/UwvB7yiCiOHDNK3Bk5AOJRJTlYZXwJ0MuNmE2vceZXt3C
i5nzvhenBbaAqX1eRRDEdnvduKGDKpTB16UQpclcM97VkfDv1/mCNJ10bOSG
RDV0rF1kvL+opfYjSQ8yukpivljy6Rh3Zvz2HCAcMW2Z1EgSUUXaljg9wu5i
sdRRqEebf4mxqA2rI0R5QOX+XWLokMbzt8V6qcbsIg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iJBjdrw2Hn9H4gQ/lnf+v/8+cvavpjmmrXkLApxlg4g/ikC4EwJXZiW73N/I
shPM7N1HhB5yvhbHRrW1XCb3KXUWGKOk3BhqNO0v6hu1tYZwtwn118Jv5sUO
IwENuUJCHeXX4UqQX+rWA9fi57BKuDmdzXDOPYpOBD9lzm8NG8STU3Q6HM2Q
ukyQEtHUHvFidezNf+2uflWPsjQZx0KPA6LAIPSekfRZCdN9qwezP96EBzcP
jwmBkw+TO4Q+jk6Gwsd6nTe8CURRs64ZMLdSJDi7kMzvDGEhJrM2+KBELuvh
thmwAAYfIrF5v3ORuresHxbTsmCAQfx5loEIFVoe/Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZUxLkwdL6GD6DSmrKY1PM8mvn/bNgVZwDXcKyPnIA9+zV70k99YQtu70Vyn4
bN6OtHXXJdCItXEru+VHjCSVQPJcbADsFUWGKCdXpz2VYQSjhwHQsuYZilmQ
qBUT2wvDcKxORGDkqqc9pTH0dr0Z0ZB8SHqsbJspn6YfG/mn0dY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Lk8+31uoC2r7MUAJFJOB15bQ5BwJMVSuLE6IkvXan5URdqF/60aBjrN6BkZM
9gzow51H4XPJQHKQP2ccuC9Xax1p8AyrGMF9jMW06dOIUod/p4IhL4U5nqQc
GZ33ZhSQXwTx3jHqVaIQ9GMSN+XBjrY6qK/cVMfAuxxYk1j8mb89AGWeH3YI
GsL3VfS1Pm3lg16eGqGQV4FSAhTx99l4FqIiAAOTTMAyNcN0UjGTgQur1eh1
g5Z6nGwBVDtvLgRHIL+RRxJJB4Fe07V7sZtohJbD8SN2gPOx/ZZ96zkVw2vZ
evtdlN26PDrsjvRPGKLn+uXXEdFRxL6P8yliJ5IeO6XwpRVgOPDMjdWgLU4Q
MVppZ3FDs2JTGA3nI1zeBYYxWIQ+qSIltS74VjKCuMcUZ4IlarXQgz8S8ig2
VAeWzDHtLO8NW7oNL21/rgeoPu3nMbU9Q+sLZ8saOjAT+aK1UDb7eYH8TDb2
sqSZUwEk53f8pkJYHhWmYSYtdVByhReH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h0FgNqPpauAnf5ev92CZaALithzjFBRchqcgNX96vV2S0dIPp7GHRLJwc2zm
XzxhQYtW7pC7Of6RjnqD4TT6HnQST4AUOfqMsRcfN20dG3zobYJDRjxZ6kgw
GttPxibVzIJxrPH3URJRz6QwtpL7lhiFrPSCzOiXz2u7QTY1H5E=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PXrZHp1vgBpQvTV1oHfkj/L+5785Gn+sCbuqBkx1uDc90zYsskCe/sDoUEkT
Il2J7o6WET+6MoGW3RA/vOt4IskPhmXDQZVScsQE1TYZ9uAizdV3qgwwlYr1
sHwJlYR+F1j1a4qEdKreIbjERe3461oLSU4hWeKQ3mPnu2oJisU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14704)
`pragma protect data_block
8m/TU2M2poMh/FWsX/fVomndXsX/K5wqlAEP8L4SfK2dx+JRWRwsfKFqkN+d
sHDm8Mf7YtPqsQ9hTxdqnIlumUehI8ON+eT9SdNiSiGeN6bZqOQJaGvg/bi1
8dP7fcqazotq5326nhdGQ4u/KjFAHfWWVO6y8oNDPej7BBBt4yu49pkFWIXL
ryr2e98gsRZ2FKuuo/J5kDXVakTA2rWsIejRFynJnlmoq5kDz4tDJcVsbRhH
Z2oTwvrWlSPuNzIZ2Py8jRm3TIPA9E0EzSj4a5sA14akpj63Exc/uBajwSFR
ro0xXDAArn0CYKNEt2QKfBucMcp3S8Arr9tgDKPsb8vqRS2E0ZSv1mJsqHjm
sKCeM+sFEwxPjh4V9aXfvAt0PjCVJwXkXKN0UsLe2Reh8ZFz0aKjqhOo+LF1
Au1k7Q6dYbylVEqKIWKIlfHXzvdHCQyJcgwp3VR+oS/7mEat4VJQGnr1ZNrZ
B46a8cAmzdVR6BChOQicMkcOzpnD/KXd86u21uxS64MztSQAmkFlTy6gO1Em
6eTGMaoM5Zf75Au7BGcLhdkvBMk41gvgG97ucp8tpk2f5C+OS4FryJMlD4nq
1GswLTYVXoWvCMrVRxq5Ws7Ou72NgeHDP+q4cymhyylutIpQ+p167hJr0/5l
qL3obnZ+AExaecT4HvXF0Ii6myZ8xKLNSJoRsmmnfiMqo1w8Zd9ld2VUd7ph
ZErG1QbxTbblG8CnOvotlJhAwM2W6vATlrvzFiJELDnrnqlxlVKGvcDHxIE+
k4HzRrBmD+DD/RAPFlaB1ifKoLKoaVewV3+vHiALehibKTispkNow2G0AkIR
81Za+56KgCOxP7QS8VCYY8T9oPcJ/svIAU5fhv6Zd1zXdfVeJCqDovcOPBPP
sK4tP/hBHyAMqKwbrFli0fWmK6HYyr2bJ2bd+MVA3aF5/nG2mw8FsDHa7SZI
nvVzXO8vS5MpZqsTlv4fNtl2QW2G3UXtr2on7eqmlt7U0HGSoDMTzweRaE4f
HzSRWBPtvyIXfIEiqDiJN6UMfRhGGfHornGGAHsnNFugg5UNucFIEzpvuIEY
PJbIER9YQXWVdy634Z6PHkHtWHSP+qxmV+voHXxjmGOaPsfnD+SzMKMBp7wH
KPtGXJBZhm8UIF1zHHKKMkA1lG9BwSsOYXBMwd5xzx43WR48PMH6Mq9wvZos
b+WhD8738wmFIDElw4uXN4tB4Co916Q3GFK5dAuYmjaOX5qraqeN7Vgf8l4w
BAlOyg+nj4CZWbMPHhONlEc79tiqjcR44U4o2y8+EmmFSEaSqH5Fp1v7iC2O
WUnC+y3nTUrF3SLJaD8luCuA39oIoMWA4MVIHjTHI1CuUKio3wlGhNgK5Awi
RjGds7TbvmGROWbQJOM2sFmZGBcuTlR4N9q6pLChj062tw6HgwrHGH6bZSRx
zoMgPUrjBSRhxkIGONh2JThWY9PPmCs8KefWFvKJH3JCszFJuh4Cd9ge/SLg
9cjxRoNCtGIIWoabDVwkufN+qDk/sOKyhotY90Sd2apRTeU2ax/FroW7YqVQ
dVaSsC2RwwDplPsM/7PNt81i3sIVZ9qHAh2aObBcaWYJ4wIRG9u25BQXGXrs
JuAyD9n72INsSXokiwLvlHLmDSEEWuz7hy5UxKzXpT/i73eUU8afgavFLzWP
IKmK73qkVbsIqE7ZRadXwghI+KJYiHIHdpqiNQwZUbotdpbEPYniHklyitmu
GwB0OK/4HF6JxQkUvztGWj/CJswMD+oEOH+E/4lRbhCVzqe1VodtH5Zigcyn
14eDlNwct4Xul57Ff6lv4488N8kEhz2rhh030VcVeDoVyGHFAJPNgUTT+05h
+XWuIN2QyrRTlvkPynR2IZ1l3dDKDN+mcBh743u10ZWTIT/tq+ZhD1XMRu9J
8AtayuMyCypyL8DO+m9CxRhxdspusZ1M9MoczQxjhC2rsuflVjCMorFw23lk
hVW+ZzQzcelUHOXlY0lxCTfInBugF5nbB6bnK8tCV9jCPfEwDH6GLry077/8
epx1Id6Laew1Dp2i5iErjsqf07CUoC7TrmSN5In850/DAl8ORrIy8pcr493g
MrKpJQ6uw7EQ99fingKhuJEiYbiZJnPn9epyq1+uPAZQBCpguDKjzkwIhOyL
8i6bgUcKDTYJfjaYX5Dy+owR6JExP73C+25Ba1fU25Q92HDbaTIwgggNVrtn
H5ZphdEdpMapQux4vbb5nhNxmKwpMpKKA0uuGt5dJTDXtduIKxSVqYDs967D
jhhZeIZFyIHiEgC2ZQDWaV8fcy2QgnifddRVD1kpzLVkhRf2W3dWG0qUxnbQ
bYh1GBlnfDFCMaOFj1kuSaa+OGhTSok8jgnOmpRRBU/ijpaA2ehNi23oM3D2
nT0Z5lFyMJwnyMcNM9YJx/WBOvswUcz+bkWpjJhLAG0OvkmdqhkCsK9CkuQC
Dp2cRPUedHBDng+SVQPvINxhii1zvc6Eq+67lDH/w3/TNyq6I34NJKMGIrkt
8CXr89GUQ1foQRiY4BqhAGIWGyAxlWsvhb45JgqCvDjHaM9Mi4s8/6DKONsp
HhQVryIjF5nrddz6gKGFpY5iGJ5D1QsbsurdWD5UijB/VbQYO1oAsEcVchky
apAQLdE2sKl1kQEGHKorDydi5OcJT3RaoOTSD5/lMC8JqZeqkyfOPkYNktf6
wNwBNvGfoXD14i6chlgmRbgn9GobKGrm7UvLsys2S6qB8Iu2vW+5cy6oPA1K
olCH6+kRmuO/YQ+Y8NJpfBMY8q9mkzEBiyuxrXlmucOKgp7FoNIy7YR1PU+C
EWC51z2MdNJfKU9NKQlQML7n0d1a2AFRZmpgmSXAeFYhN257KRIT9HhMjetf
7lVJYGzzTsqSeeu+Wr33Rf+5X6hC39ykrI1tvShpnBrnUVB47NLUov/Pj5Z4
ZkyD8kRBjfz6ZX9Eyd8hwP1RT8rRJg+O9PJk3FUpluZmMp7MtQ68uOvCJhfr
GZm2uiqaSSMQcsKTXGaBkMsHdjaBrbg45Oq3u+Cq/fXE2sU/FBA3OecrEAmq
8pT4gAlvJ2/VbGX/4o2h43zwCVFUsVG/8A8sPHaTNGMPeehlOCq0WpRGVT88
8LHYBsv7us7fTHl9E2MpyCIFHKq804p6mVw2HdDyEqKZckkH283UrYkwmwqC
hnhVIGOv+8EJXj/J408TBgHAfDtgErGHcxcTMyqzCd1Ovdj8pN8xuWsmum4T
/6va4hTJXWygKoIBO02DfN3w76lksoog3gaACBDIa1VsQIn62u68XhUmDYXM
C0HhXc7EBTUVrHWZs7cEcgR21QDOznw6qK5/RgW25xyyKZIYz/cqmTmWrlM4
Tytv2tac5LljPRlKmo9brPsL0/ITxncXVWKrNrvwD3zHIurRfWUuaBiy47EH
bmbgJfP6F5AoXlOkxOd579BW0oZjQRDzOfmBOI+ZPt57Q3gYlh553ey3anV+
toztOparfO3UXla/ubIgUJZmvKjdLh1UiBGR7weepqlvgWuWt8Dx0OChYlqJ
6LADHgF0WcxKVSVNg9nAA5z1d+HV9ECoZoLKAbeYNASRVKwhwR9IxG4Jf/Ly
KHHMX1KXPiLYvudf7Yn7ZHM+nKMvysB/S7JAFq+I6w7ifKflsg5NmUIvtGHw
XlRDSgZp2072s9t6dEKX2xtb/V3OWhWUhW+cKCE/WuzHB9jUnrzXJUXkwt4T
cQmflE56ySfQ8x/oGvYnBVpvksluevQur6zgaDQb+yfuA6ieYTi3EGo3WYzt
XvsUC2y2Debvikw6Ga6ao/Tdcfsg+JAiFUNCfgqnKWm0KuUiablH9Qcj7gOW
nZKoYGEp167KrUIOFO3xre3XjQ5aRqarxf663q+5rouRgNbJ83XqWDeqMv9u
TLn0Xy8n2zDMsdjMRwdE3vI4C7+clrhFTDJZE+gyRA+LcgYWBLAPl90vPxdX
WlHhtZZmHLwUIiZjFvWSrWZJl+09ep0I1U0PhhdQLGBVhOYpT+Rla0UmhYuZ
+0skwloTUykYFKEHC1u7Vf0XD7SQPDpuFxQNr7l0rbkBXJ/d2LOnyQUL9IAv
lxfnxnD/sK5H/JPiK8PQ+fuKHNnfJmjvW0IcS0yYr9B9bYFSNjohsJjc1hN0
4tjSEd20nXVRmCZOzB2GdXE7u1hgfKbRie5fVaTelerakLidwPiyVZE69jPs
K/oc8PCaxUkHnqHADtR31EdOcUDCqzb/IjlrUdyVlnwtBzo2eTCQnyugkKMX
uPib2cpxPTPAvcp2SRWFIXSqWRiQfVy7glYEVxmrDM1MeNYJh4q8+djALRLb
rfIoUN/liU3nezwPR4MPopbIJeNT29NGoihIMITRZFFHuNyAfLRJIzj90qlx
L3opn9nlsR4wiPO9avqQjpIj4RDIb00akAZGkgLOTXMkmzFI6tMtcihdRrcd
QQ6HWzq/FOBZRx7hjx1K9jjTETy3hGvzLixFJbDbX5hiZQUlwrzpoqYe2tiE
b8ZzDW+lMG0H7JwmU/etbohdh0J0QuUHQa5yjtedmTOd5SNT2DoPKrrBM99z
fQ8DH+LSP8c0FPND3o1oNB/gbo8l2CU0PCFRl4LQJT49kAczlVexxbiKmhWX
GVAmaCw+nFwoyYHWcHhGVRyi9zNyYiT8cKgc0T9LNJdjXDpTkr66FpEARhdI
QAnArtl4ITIJOjklDAbSawTcirs534SFNPEsVIJ6WeumDRDnPhfpoTqVSJCf
uYMho9Wi6K3J0AkzaXdcVONTHicsst8Q2shcrDOvp2E+JsEAOm1sCRulZxX3
QQXFtU3F7so61VaJw1K/+9oTq6Moq97loDfzRaFHLMpNGQxSfjr2tfmFFH9p
5FvjnubF/6tszdPsOdTzeE+GPSpXlZXYFVMLhPeBop65JeR06ODEgYqOsTTx
9xY7knPFVulbhsj8+nP+lcLI4rmtFPEV2YqW/sZqvsJJt9dhmBC3bvK4307G
7do8tFvcQV+ybUuagEtiJEHcKQxoLn8g5+HpLnk5Tyz4c5SzjuQvkCJw2Sb4
XPsy0nFIKS0HjBKriBSX+PyKjY3NE3lDYm8O/Ect5ZPRHzrvQG4xPsRnv5F2
uU5CSx8/lw9pEWuxpVwYOxOOMVW9atVCOjC1QqNP0t803FXw9Huf0BI6OUjC
k+mmBS1eB6UbESYhamQ20bZUyErAP71f1FpUZUsFZElCt8WNbOAerOYNho3f
FZ8tjtvT534h9PxR9sFLJeDOh+6hjROLVT3z0McADvnjSvyS2/g8lXrdehR0
xpPzjsnCE8/QbxBU3CujnMEFCiFS6Bnmr2Fjbn4kCHcKBQb0kNRPGkkvElD3
sZCzUTTf3NbRFOkhpwpkvBRNnqelUkOOvT//tmIP8jMq7/8MmokT66PAnxJz
PjtUPvsTV7vzPExZ++lVCeAaoV6yr/Ae7tenWpwE6np3xI24Fr22Y3oVvIVF
D4IO6p1dXYUwAV7ndzLt+DwabtlzZmnbTTAs+oWlfORHyebCgRr0wWg7OB2e
1vJf2zgZHSLOzg8iapAFhvvJh5PZdwCmGy3UMbRlnCKznhZcuYPXwQKiWAse
CIaLGdLDOvLfgqVOhnW3deG9ILcbnBFPszXV82sVptXItB+9l7XWCSMpa9la
YcR6XbruoGrthza1qvHUJDIgIeTi9gixDzrJ0HOqMaNJc7ob7YQeUwOK+rwr
xvy5iNwxKx8jXKH/znN4jNMu3MPnHw3mZcxaCOyE/CK+R+oTdBf87Yin6ut1
EspSk09C79AhEq3eyWiQldGaRGsF5S1Ci97AU75puoy26Iz6wOGLZXy+U+tn
nzhMkrzSbHKeZWZmhgiHyaBweJl/sT5KgwRJylX5tDXELyIvsXkntIoAy+Yk
apJNdMXq+qQtl6zKnNofd6+rtuc+eG2cNcyuEDTPlYUuiq7B/FQo+QcznOuq
9Il+gV1lAjKZ4YXoSeY0psRr6eU5eYX/YF+ksazBB8YFoxFf2rojOBkJ6Sji
6VyQ3ubfYVsWmrDShmDzxJQFqdMCc8ef4q/+JPiBRb1ushyrvNRJbWwNkBDU
vBEbLVeB/Ok4d0ZXtVwIIgS2YFaep3alYa0soIeaaXELCYQ9G2+duMD4gSn6
5eqY5EIIEfrU3NzAefVFEPmKyFu9gyljxu0c3URL+CPw9brIrhSi5fXXjQ0g
NAYvLLepYUBSHvsc1xODYaag7s+C06wUr//LAnk2IuXSLUKktVPDnRgW5TN5
KfLbQhCYRRP+qvqBkTlqheQYzDEG0OC+ke9GYyHAxcPAaMv76I9PnKfSLaY7
2q9udPVk+yQXeN2sRhT936TgI7DSIeRgKQvtytl9J6TqpAcANiMTFKMJh8wM
yBvwWwL7b20G60IT673+fA92+U+0O6JSWJrzxBG9VXHVK1dT+mZ6xRn16rEn
nUm0RVNlXlREayr4lcytNa9GKBWBLdj16mfw2gqoknBMxmFC1jnFgp32tUj5
GSFF/5Cx8hFteH1i5gf6bHDOZBJzceLC96fwJJRF5KaNtA8LQQsuKNPM+Kvc
U1a5W6+sbMbDa4hMHC95qOOFMzPu0sk2wr6whHMhu9OLEQlC8zaRU9yRuwdo
Me5Zgikv1PI5HWHkbUdvHHNlVP2iNHPj8RLcWFHMKIltf95G2rS6Zm2QM5bN
buULls4uJ2zjp3d8bynxzzvN4KlWkOgqnmwxrZf0NNT87hj+6liX0Gjg/Ex2
rtjA+86c8+2AJWhBiUlcV+iXuNNc8K2eo6VIky18fqA1Ug8SA4P71BurvVWz
rkmWBG3hjuZCDkSQooZTZVb7Gh5ESVABfh5ZF7BuVvG9f/pxMqMaTpWJdW/R
OBxuYWrWEw3ucuRaTEgKdICf7gypvMDIsgdTRNPVIspvpXgtLxkcDS1rNqLE
C6Idbk8bpu48uZ6Mg2i2ARDOrvOiuvI3g6FEp7Mi1OmeZU78Yj5eYbRpV/jO
kHybmKwO0LQhpcLtu2Ob+Qdhan4oRiLrsZt8QaKLZ8sfDuYuYvnFyIjWLgTX
fia8VhNQQ9zNt3/UOO5lrwtlWsf8vHFd47Vv3ExazvOdklIDDtA0+UCYMPz9
nfZwxW+2GQrl4s0AfwYQDU7X4ebmv36SdXC9y2THMcm3r+Hd2NAzqO8b9AAn
HY1Ky8Hk2UcUUlTi0rcSJzdQ1bWgET+4coVW11/a2Dq7yXCnHmoEmgVwBdso
lHmJKpwIFGIYxcbXoIIcvqJQ5PNczl+zqTDozwCDAULZDnv6uVDQK6QAIHGn
Ow6N6a1DEFAeuGD0a5McvVPQZ3zR1keNt/uGtfu+xWqGMNMOkF3UMZZ8drX+
ar4vfn/lGLQtZq1dgjBrtgSJBjbbfp6qgZEWD/kxxiBJ3Ftpx2ALpO3umjQH
R/GxItki2FkVzSotPa6U+o56jY0eJp54sSqKyNbAhuFuVkEPW2rdTzA8Benq
pkABXIXuHd61yNt90FFEPV5eW19Pppth0q5GnFkoUcv3p+u2tNvy2UMfs97I
O2NADWshpJq1HYUnIS3+NtFWcu4MwZEPr53K2n/pR323OQoSFhWFNCfyuL2g
CnVHAZFMhox3Jd3ueRTP/4l+LC72XcFLI2EJ7GzpjvAfGg8QAwzd+zueV0l1
Y/AWtV2YJrjdu909gxaVTla+yAYQmlDE+3znhbMiLkwdsx7wlP6iPQhQ8GP3
W8azqtdtk8Sy3I5tsek1OfnnkbcOdc1P4Wa8QAnQSDLz7FIEdF9Jkhkdxx6z
VS7+OccYYT6kVa04Z5dPYk/q2SX7d8qPqdX/QtH/oB1ou7sEvhnOl+B2J4gF
XGl/IIw8DJQXaM8cUE8kVuLdZ0h7yWpKLUL7cIEORiaK69CuTb2JQqtrjk5a
183Nqkp9NbmPUBzEVK6eb8F5o9F5tQpTMV6q+WpAX4Eko9+jYhTUhfTpaH+O
CyZR1popoloulukKZkZPiSksig+m28JfFzjOlBEmUkxjqgufHEb4wj1QFr3R
qBdAilAJjf9yiJ7vmZvEnEd0UXxuh5Wyp+UTAl1WjMDk8AhpJ92HXS+PVmn4
gpbMKSo1nQv8ktHivAxrIpOq3zAdG5qQgJwIGvIQPoW9neSzvdYc2TeH8d2a
vb86DDbdg7fE7bIvRFzf0VGZZlQm0GzeGREUbehBwwuMIh5PS1tkeUZ3kTjV
hF60nRtiTH+b2UQwxot9yNW5SxWL2qkzNpjnZn7gMoLo0gLoG63lYJXfpgMJ
kyqsmQkYLxf5dXlByKKVoLfziC1RWw6Jur8qhg0ugdZX4OAEIA47YtWO2g1t
SdUdX7nS1/M/h7Uk/V1JXVLQLPIQPHQhlejatK2tW692NorSA7FmQ7aPWMlD
jSTalY2UE9KUqoL0PpgYQ48DZQ/G+L5x6qkIaW9n9Hi1W2MsG2HI03kB307d
htBfgi9iUSdHKUizEkBMF8ZziidkzYOHL2tukdF8FjYnpIVnqsEIzqQxFzwl
NSRLkso6zCSRZMhTg1D9tgKBN+cT6sP8IBPH1nSUH5NiOhM8/uxazbEPE6Bs
TXYQAedu57qFQFCyc7yj72Q70awXZ9iK27QFA03JKS5gG3wrKjnZ4XYYaoKm
qulE+UBqlmB2Qg3lSWBFPPtgkCESp7TLdosRtUurzhrppTXkwt09tY6us1QR
FqtMTVmmDxxGWV7pq1x+wN5lB4DzWI50/BXn65nCkblx64zDyEJYBbbf0Zia
EVNY6+3x/V2cxg05CKFwBNH1Id0OLR/d6Na+P3eZGh2M5PBRlnH7D5ShLvhb
bSQH5J2VXRndrk+pX9z+Vkgrwavf0UOgIwOGL9Ioz5Y01aqoOY8xVm2CyS8a
G/jGPoBvhN3MEv1w357ymSaEJeK+nm95Jh2ryk/+2SSyHzthyX7d3I8Cefgy
EjMKERiq5LBJcXGjLeXYLJ2TFBlou0sf9SOtVCc2tVZ76QGq3jjnFAyQjB+q
/XJMZp1Ag3u1jHewwzhLXQiDceYBZZAmrNrD8UwWGosxxqxkQtAIzjqumZZm
NlFK0dAf4uwPuAYD+AlJHFPu0TZkh3kloDWZ3vFfjYh6grfpqrcPCOtmVCpk
3UXza9ADH90RX/21C2jQPnaJIDYW1XrazdZO14mnd4vwNFjn+F3XYs8mDspM
DgSQu2qfAFAyifzXf+4YgJCBIOfgZxWvTqduP15XwX2f5ewE0clmq0mZRLMc
ZOOxaiis6xxhDmrUtdUhj2u+tC+WnF3aHVxEkc6n/5sZXrrFZMcdX0/NMZ2S
v0xVPToqPHqOyweFE4iT21b2JNhwmYq+F50/AJK6Tompk99mTQwp3xfEexjq
AGP6nFZ0LY0L2M5IstSYOoR3hNiiKaA+PZU7LhOlxYT1NIocvNol11d0SLq/
WxzxmQtYzRbM9Ns+6DhS7NApUSrEAVaGmbDt1/ZRaLe4xDwghbxE0SNd4q37
Yr9g9Oa8c5L0+Dcwn0qUkvInQXGshZ0sKRAuPzR17oWmBdfQkIKyj2fvkczs
+CU7oNnxc27YyZVA3uuxmRQC3auOg8rA1/5XAl12PLF9Sh3mguegfdbzIFKh
d/3qNDwKmw7HToylWtQjs/XH3Tiz8wgCpG4gXdCa8C9gkn/6DbM/TlgOx1Sm
lDmcaJg8ecsBgej0yTWum2AvU6GzBf2GWanPJtao8nSA5TwqiSGxyV4KLzne
zL3B2zOm6FOY7bK7WX72BXYAmOuiX1uHfEIB1bWn4Y49YqtYVYGqP5dTVcLx
qXRN9xw+oxVzKi3YMeEQmrtRBsRnHAFV+ifqVkuLMYZyu+RmWybIcDhR3mZY
mLca4acuu2Ty/yXrtWaqlVP043kXObzcpl1pVHmghlXJJnJGwo8gJ4nBarld
QWhKeaUoypc19b4lUIJW7EZVxrIdYc6Ze+NHmoYCctne+yLMTfHuXHJ3qTnv
5Ydb+aVo3F2V58G3pob006dO53Kj4okLw7KkX2AvJQRGOWw1yEF4vmsPQ1CS
jCh+DxupZ5O0OJfqvTKNqhuw0x6HbykUHcUpI5ie/LQGKIwHe3TxZR2Gv65U
HnOk+6fZprG0SEvTG/BC6XaUR4vrYf15cQifkprjvosBC8UBnsNlAUyJTIoo
EWpAHDZOU1LXZfCxRhyaP2E0ON1aiuR6dq7wJ251BOOoc52rL+pmv58tT8jQ
Fnf9ccBdDEI4OBhI08t1CXEySTge86QXibUcMFo8OiUwQeviHJR0IGsYD4JN
RrjrW+cZEQItduJ7t6zygldZKEQqDqbhDa95Os3tKn5GeViA6kuAoKh+ozpF
vItOEbNg4gh46FeufP/F2GzEMm/MWL8wfj9O2+eeV8QfZGt56X37uPirCHcd
wQWl9deCzgfaZFPRsV8HAkyPa0fxLYwWN+Iq7OVt1J9aJf23XDl4NIJF6Smp
vfpsi6teaA29FiIvYFmRywo/dkeio7tyPJU1OVRIYSKg2j0c8hqC89i7OZOY
rVc8JA43mjZJpYtPVlvhCYktKAR5E1v6DtB9nALlHbf0+dq3ffR7FjPhapab
8JnEbEARri3B+ym75RzlraBdFRGgf9JXPzGJS6N0HYtgfm1u61ckW7VG8b62
nmQSUrmhMZkUNCNwHKuFMSjNvVcM6e1QahL99IPSs/H04JkXfTGynhTo7fJU
cvRvlJHpxsraCvipfFjERl8nYSwRQ3BSWsl4Fs0/LZv3IcSQXwjRtBnp6RvP
G5nO4WPuvXMi74NhwisuYtS7M60ikHcEZEYU6uDzkwtrnHiDLDUKnnftkNSs
Iw9i1MERnTlbEI4avI3APnByTEMkIi7PF8viesGnhNhjoxv4A1QbL/xfXjT5
35nn+KDM0Yq5Jqj4RY7vN669SKDfxRD5bNYId8cbeRSKg2QRbKjgxtKeOyn+
4w8KH81SCkgy+zgr2mUWuW3QgGsONqf9tpmt7Q5VVsEz2CoKIxYmHUrAKur+
qJtZnz1Oy6zP26nkvv9kHXTlIirmrq2ilkCREmlYFj7L+rIsYxr6PjdFALw7
KLwMG+vn5fi96GTzX1z35YIdmjZjILeJwVE63IhZivRl3MUKBLWf84g8kHDk
9g6TBd/ip2WV1RDdQzXMj9JCzy+TIB2edrIbDxeI3Jc2NnH9eTuZyDCjStYf
5kUjRC7DdktWhDPTcLnFsIdemlDzftgFG608/cbHDaNc9ThuTkFfAKYx3Wbg
dIjhq9JbH1zsyDuZ/UcPxfrEakNtufmXRX3pMM0XwXzl8zrnTq+88T3x2oP+
i6BJ+9pFeP0Yw29RhhUdSnyfnZ6SDHNszz/ePDNsh2i07ll96VXxNHYaiCp2
PL7xZFqeak6Okn0G7DsnDSoMGYrYDq4cbflyLxOml2WZGZBgBrIMCNb5PBJw
qlPwPrrOS099nrx4RGk1WHSlD943M+RRoLzPl0/j6u9WDkymNAJ5p9HICxxi
ScJRQ8IusvHMS3aLFHNORtsUJjl6rSQZ8qnlBvkNuDwcLegnl5ZnrP6prDjT
1tjuNKhO8Kmrck5AKah8mv5okNbshFYnx7XX1GKsSKS1vFrQq5qYQTCpCNCc
VNgp8HkbR2ry9T+mM4LgZWVQVegx8mNu/pMAEjyCw19cCEL9V+eeYD18/y5Z
YOOfqmd1VzTmxYGXdGmrlafRRzTmEF4Rt/ATHSn/xHYtMbuePzFscw8y1B5c
Opc8VLm9upz5wH0fpTe7bFPMQpT8ZzwvcBI/TFT/+aVl8K2F/6kXjhMF0D/F
duop9l4vglHwGWJnATJGp2QuQRd89c5ofN9Pqdjnd8c5iD+LWxPgR/dhIcdf
IMomkWCnrDjFhjvYnZhFMKp0Ig8tXzVDKIbaPpCdiRJwElxQewNNyP2kj+N0
ldwkiCl6UfU3MeWuisFyXetrx2cjm0sb29uEPDnJjmE3Nt6VBcpiGHoDTePB
2SLQq/m45yrBuv6/P6hyfSgBNL/vqdRdXIqHVE47DtlQsot6LRPuPkKwulEq
EvHYAbrrCeHz+MuaFqpo/xv/QqJxik82eJE9/trJrf2svC6N8H8aYp+DHjhP
TL1/AJKHgDy3lJDan46cNUgSBV2jkQn5i9foTnCSfWFbp2P6TMzxY3gRLJB7
Ie18k15dVsuXsYtZgjnP3eSeFa/BETXunumHaIGiDdyuLvX0IqYKUrQLp4dQ
qqk1m9H5mIX4SDM/gbIvgyfyxogovcuyd3dVLzbzTaLvcGxBJqX2PacfDvjh
4vunQaUIhhurMnkZb+n3860YwPcNa80pYaWgPWCwFLkybmXZUNYtZ1aOMLJn
m0/65JbaPiFMvstvMTq2Sjui3c2KfHoJtdXHNioTvPi4PUN/v6VHjyjLtBmi
VdOfDPtN6cbQg5GC+OIw2PXATyhu4SG+a4ExEB+VxifaFA5UJfjLhGZpAPF0
zcM0I0dgdNRkKLUExqQCMHzTcRrUbvt/wh0pgN/Sq/b+nyst7bkw3BAawiL6
h86htkCKgXn54TxhUWBi7aqkhwXEenQHMnULEsNk+d2kTmFlVEBDJsPmXvrM
B8y1wQdFbdI2fix8GTyw3O43EBIny7/RV7G+iflv/BcyEaexi7ZNUJNBmq4I
qNi+ublzQkddNRyXQVt1w/5M1zTvcMRRkx/5gB26lNCgPam/2cJWxcsd8IEC
2Q6Hz33CgjAZCfakKcXadnb1MK1FljuhZvzkk02NT9cVDiGtrzhoWKYALj6p
Fi/CzBlp7AJWkwev4MH4lMGNuqSzQV51BQHg3Kjo1tvipEDiSvLpjhAGHeW3
DJsCpjCFME3cEKBpqDxqd3Mxbkw2hHWANwcyRn10AJsbOKXBWCKITPH1NJsZ
TJY6Zk/vfwWgocfP4DuvoBdbZE+zvE3I5HAqxMt/Z4miyEmcLa/0hYJ7DtoQ
b/jzYhVz/rwtgHjHsxlpvpOZgJbRWAkqvDhstJAbcrXgQ3JYzHHVuc26V16S
tFfi49E+Kqp3kbcK9fs4GH+tD/eeKxvBMch+hd1LN+fLjKlememhMxPNcof0
pGX/D/wYTkwqdjSb7TQusTcg9UqAAKLjhT5vqR2loaTg9aMujBQL1OVYW6Sj
iqv3pGfwoojgB5uqdTuLKJ53c3dWSgdhZg0YRggCKM77OGkgtMq6au2IcD3/
v63/LEKpFxhfi/ONUFAevuY+OaWw83RtbWOZuQgwzIujJcfu12NA9WnmmtVU
YSPP87we8rPPr2XN8m+TXACgnAsjI6V2SwPk4Uoa0Ae/iGjlZ/+sG5IE5n/j
lfja3r/TZHbOZc2iHZ0wF+VWGKVjQUqFQIBHTffNhNok4rFTPhA+sYLKrZ39
NLKJMY/IO1G2GIk02T8ZA99Ub6L8AcWkAUR0TV6RYOsyl9eYjzx0GQLKp4rk
iIvXQetLFkHRbpm0CPNgL/1u+WHcQXvI0PFa79W3KYydOS0Ah9I2k6s9sZF1
PK+e0XCvy41bXJHQG75uDDLS+KYTrjdh1niDTzLInb90uo8aK7hW2VLCva1S
T1oqYs9YXkRChDVFQ9lcOG9BASWARJv0O5ZsWPpubsvRhbJg2a9GrQwpgnuL
vF8ziwTKLoaKSkiM08e7Wyeu/PcVzY7+xzElGKK1v8QP3R8W+b925zjRNCd6
uMrpdkShOmxZslBeiTomQZKVT5KQ/Td5ITBRhR5sK8i4lric4Grd/IsUfpB+
oqby4eqTCeGHE9A2pAaGazO6chtXMpxE19ACM4aJZqzexa2sOtbaFLnU1HgZ
dtHUdF0XM2trWQ8RyrjDHvk4bo1rFq9hShvWUuCUWxSBnQWVZ2EyHAI0qKYq
1d8zfDQkZf37/K57X5aRoNkhLcDOp/SUrp9/b2FiXGCZf4H2qLRzIhfKcQLK
Uv8q7Fpzf46fKIECcKFRwEi+fpnR1C5fH5ge4d3KHuATu7ySp7qRaoumLe0u
jqW8Q1h/ek3ApTrHfQ12Gu9uAjb527Aj+eMNN0CesSlbNrFFRsm2p/ZYn/kY
74ojpFjBo38VTnl5XsknvnE+GyCFocdAeApFyQ+MvtUaTXnWkzl7uLXlwi0x
Cpfu3TPXAXGDBP0gwTnxDtskrpXeETe1fauR2swDc0KwlDKbQ2/hRumDGdoe
LqCWgK067FVkd+dGB+/GBQWeE08my1qetFZZEHbkJe0M8viJpGXNDKYHVIh+
bIqW0j6c80S0vhI+1ECBmFC2R7NbMTZWLwFb9qurtJA/nmzgH363K/txomGf
okkrKlAHGmlckqaXfILsaUvXzjHHU1OYikjwhDc4cFj3sEDQqZ1HHu9YHLqB
Z4GTfTvAOyvMmhp3N1wu4dZBfY7qc/jP+zIWXcU2pmEhV0Vs6foG3li47xba
YR2j3pYNTxeA5sIexbqKOAMBwH1qXxSUAt4iVXl/aI0eXZBEVMSklnIU1gx8
qRNTt/scM4Se29LdKL9hRwcu33RolYsrsLTakP1ANprKj7S4Zr4OIoL0MgWa
Q7rqKlxPF69t2jBlSVGJk44uJIwEOXaWPSFdqNZzBiTzv0+mrkz4GvjtZCNv
KBqRZMwC7V9x4vJnLy2/G47i5Kby6AI3Ocmmp/ypJ/WPMID68rYtQcnMzPTF
MhcAZNGuKTG3q6Qd+FDwJ5E9CkZtbiXePU+/4l2/l9dL+Fg9pBtZvOQ7FLba
SLU/lHOpY6Q8kII+H7JSJAXrRWYIuH9z0seRaWsrpILGRlizoiblz/2FPa/M
I7BvtTUC4aKtqh84PKBUKwLlRebTSreGyPS84ulqoCq2uRLpRwFBOSCl2ss5
5hAcbV1sLg4cmwgZ49BmFD5PUIsbOiCXoOvJkghf3v3HiyjRTJaUaQ0GZ3dM
hUUBwsvWhn2qQQrWvxUtBrXAowoO6xygBTbiU2QSYqGwBs9iQ/EyYLFmNEtp
ylpxtUR/5IojOaOtuoGOCX7TOfxZBPVe8xlpr8vT+2WgZrVqfEYbGDt3cYA6
72j+xCEbGniqQsauwg5jykWUsvwy2boOj7IKlwJge7QAUbfI52BrSbB9Bogt
DGQaxSxjd4jHl2/71aGDeXckFgRc3aKw+djgUgiXplEVsdxk6uPC2ZUPYldY
eZPThbb6V1GFpuIJuBYWx7Pb2y6AFhzLud/DNGvtmuo432pjfdtXRTFWhA3Y
0xiS/Nn3avfuKkbctoLowaNBIETtlfZtaWX4KrxoRiue1wGjsKEzYcR12tV9
Cf2SPpyb7qN7+uUDSve6vzVVnwWV/K8UqZclRYru/wdtUipBp8zNKCX7rb5g
H2jw3ZXmHMaIGw2AqjhWev6WAsHq4CurtJIO02UTYZClPkSiAN7y4AMEyWgO
VoFBOgAkUGOb2o22GwOy8iWymGziRlq+7e92Onob6bGXMKmISqlSQ9f+GVRd
LOIVvmiGxBDb7s83DkKjahMpy8YXAsTJ3cePTA2jagyP6wU/vSEunh55/F60
pbaenK2ZQ2B+rO8xyAfx2GrbGeUvcpYp9aMcINH6cFYcm61dmWjryLaN3YaQ
C/0+aVOYJc9y1dq7qA60UkIDC6qcmfFWB1iStmI73qsnSA/PXxseYprMTghh
DMA6w32drHCFbG1Q6sjsa8cjMGzDJr85IpWBWhj2Hi2VnnwRgoic2zdcjClm
ttmm2rS7SIgMDE6EVJApSMLCFLnwbS+cXiBCrBe3gYZKK8j7W3czbPv0vNLb
sZ4bkHH1aLCoeJbpd2VuMo+ucgM9kaTjHqz1E24hAcPuzyTuoEMi3AXYu5x5
p6cMYEhJNVzLpUYm6x5j/tqW8Vx/e6BWrEnkkjo9H0C1a1E/UKmERXxGRbXL
Yz15I/HBZRQMvQuoCE3eoYBUF8VuUnh3x9NAGMnATeWBVMH/ssBjn1vN8+rD
DjrlXEf6TLQ5Ywq6kXrj9lCwPJYoJMHYoXYFfh0tsp0z2tQecjotZ7nN5XOx
Fb/hCTPwl+xoiqXLZc8vIGc13699ciU3lTlFYHKlyBfv8zRHPw1NKJFg9dhJ
UTPgK7Cj5WjL1cl9kK1EbSngzsLAilgyApBxvZeiee8jVu4oJZvUHRiuHLff
8T0PyLH4yisTT9WF+qOhBj2YujoK6wT3Q1vw9GcyZKpNnwc6jhlasYzLvTnn
nUcts5/4WYQqQOrNCVRlgyepv+w2BkZOZXll9zBUAv702ozWJxbf+BJwVM9l
+X564Juky0kmN4lZ/RgoD812EgAp3L9kl4V5jl3x7OrQkBX0O/aipBaxWpWa
9LhSYUdaDtO8XCbLeG2mhdSywK917l3pOnKDbFQljdx3iEXa6Td6qoCduzpt
vVlUqb2uaV/hYlS3RpSFfF2RJW4RaodRDzAa7oYlMkHTz2isDi2VGDE8SPjN
wDqvXnZm9hH8UTL/aixAQ/WM4cQ7GTxyvVHtYpy9IA+GQup0PwmjS0O04med
lPWsCI2IitSMM8YgZeHIbbAjwmeNC2RDrze194JKnCV8OYamndvvht+zyAji
ywPUkSTm3dpdFU1hDOmMNtqUF4yD8eyDNcGTUVhr8zumYB2AxIns1F6NWKYL
34kyad8Tf4ijoLp7tHtxhByjrqUjyo0M4oAhnW2hItpnCfivx9AQw4qpH6QB
iJi8jIyaoNvHVvSkZ6un0Xa0X40HQa2RLQq/h15YY4oV52+ZBxVFf4io4bnR
Ang3yJzG4i6SYRLd6Luyn1t9trtIcTRwWcA2jvc6vgtGI4MgDhPpIGYPn3V9
fNzAFyHc45MUmG6oTrLsdTMEXv5Sem+LM+Zezra8GKNTuNpxCPgwZZAYClx/
TxgXZKXBmqAn1eNHJ1sT4xG0HA2Akfu2fSuwAs7M+1YB3tqw8dI3UbPP5Ms9
ajGoiO2wFUjBhIrZPGctotc53/yizfWAMpu4SkiNHWQ4MSYBAIhbZrv5GEjH
+dmQVM6yczwh9va8qqmIIJoE4h5jKKzBP2WSkjo22nwwKHafOxckfJhKirO1
RWWmy98IvkYfDOPc3vhHPYNuhldMDJvjk2rd7WZcd4xn2mRG8XdrOKu/1OYX
qUu8dY39xSIOLi7ppj1aM0CSWtN3XMd8IB9z8ObcV+XqGqm/TUTT8FvFbu4g
iaeazDbrdSrZMdbnTjEl70nIAagQfHpIozZraRnXGqPTBBLphzDd6brIRm46
r+dOzbfqoKzGpFKstyI1jrW6rXhCMNquITwHJmhlrIT0M6H0fWecddz2S8ZM
Zw8Rn5DyDSDS8vUqWcxAvf/JKCMUA8Q94Rg8dNp1ivM4HvgoTCnEsF8aZ+5P
d+PDQx7a58cvRSWracIh1Dx5yqGbUrvom6CXRPZ2Tt5Q9V6zKdsRFbQUDSPz
y6eQTJxB+R+C+ztobOca5XmSJ3/DwFIO+74xDPOZ0xpX7iR73xO7Dv/L2Gqs
0yy0xiot5enuTAA/cDbMhJ9KVRgnxqIrj4MXl5KnfKiSs24P1IMQL3rDrjRj
uz88fNGP7uFElJFbEXR0gGPaI5gKqjlSzRlD3tSMn3r7QDmkxMozsq5s++Bb
pVqv9X/Wjf/i88j3JVDdM7DOyW1JntUc2aog/G5lUMaLKXDU6aIjywoppKV0
KVPg4VDyzzYXFNJsB6YA19TLMBIVAp+Nd1sRR9RP/TaPxw4MkCwVO3ljj0o/
HvzYFxORhi4lBNDXzI465MAxSX1YjLuxADPYE4hZjENs7mnxxi80QJEnBPfm
GHV0xfWQ/fo39xSzTty3WJOSSx+AJS1ccCfHLhtI9u7meoO4BRZOjQ+AnMaS
GwESlbhyhKGYwHIJnEqFdvanyVf5RmUlbERxyLNslKnk6ZMd3KjNRL3FER6J
wzYa+X26RUopUUxdX3+o71Yt9YR7PspVCwN90wGQCKPjmt7sW3aTYUQwB8XS
+dg43sseDX2f70EZDlmTAvmDOMr8ywl26HU896XCaQMh4P2Kx3nU9aA26P4x
Z0uinVchnddsV0ztF2FlLGebP6LjbmAjsdgYmvQrttGRDLOD2Ez0955+U/4Q
hHCGggXIXjWEZ+K5iWat6xTX69eKvt2sByNMXOgqD6bO3cHVq5WY7qGxThYW
+e67BBPoE1+9scLO+VZgOc/iC0Q40x4F37p02Gm3NVlIr3n39gYx72GzKlSJ
OIogM+Z9X/8XdfM3NOY11FfV8wWl0lfAGWh7EtA6eywep0UmN/J4bAWaSe2M
Z2MHYM1E2jz55Bg114HPm5FcJ2pSlS9APUH8/TQZ29bQDZR4sCAqlvNDqdha
w88PTWB58mgS64c7Etg6iY2XFQW3Z88D932iOt0FKgQ4W9kMwUfcK0ZUftpn
Fbp6fLSQdZKVzWJWg8FFszHAnvq6dfibz0QlMMQjK4qNXWdnKK05oy6FlaVL
YTv5zP5OKmLp+iksL3akFTSA2nso9+m0OxhjQwU5Q3Gjgx+JR/+saJoO41m9
dwVsCpPl14W5DxC7B0dfD1/AJheQ/zaJjHxeNyyn0bE9A5qvrTkkfnZCFj7n
JPKWQA0id8h3V1FiQJlBdIhFap0T6I4hOWBCi4WPb/53+dkO/RA4ZSMGRfG2
9yraMnNLvlynd+bMrOandmOIHOgogX/3KBBTLD6VdnjqIOgXt6C1QYgd9x17
+1neYVYaDC3Ulgv/xdC+sVMeMSMDr51m2kv0kQ5vYreuS06NGDg5gw0gQI8w
/E3PlWyxLn8YIEXj4TXogrs8iJaaYJCwxtK7UwJ31u7W/HBEuOz/mJUHBXkA
7hzzBtiMDOKj3F7WHP+z2ogGN4PmUwOUCbC9dTrxIy37ZyW2NyECQfG2Fjaq
pUIXbv7z1xC4o8j5ns7QLYtkBuLxfytFHST3/MjvBz7mDDxCFxobjsFFEUpA
gKQT1bnc9qhWiQr4DZVRgnui5mvGt0Os0iDqPey3u2M1LCUvzzoggBzB67S9
nKvj95UvpdKTMvjIKQORiRM6JEqegODklFFOaVl59WDrO1mefbkvQ4Y5XNQw
WaEELjpSh9oUKgmcf+nLO3Q1ClGH3r/HPfYm98D0D8uLHoh4BDVPH5LraqcR
N7tR5sj/K46lIg5vU11KoFoB/xR8utEasYSGelkbDBHyqXF7Ck6hMy0PI+bZ
mQS7xguNMZA4cusBFQ7K3FNGT2obCQV20wQH0V+YHXbxGC9h7rD3DnCU7aNG
jU3xKIAUqqU0Bw7ANs+lJUKGc2tUEJ2ZMdaXL/DmDrUSIbYeGrmVCNR7+e+H
PkKEnZlMGOIkmy4ql/XjNPYzmI28hR4BL8LoymSbolRFNnGGJRxg+igm7mvN
QwDDKgyiuCYWyK8IeW1G0Lhfw3LQ0KCZvE98WZ7YoncX6jVGdJc4x858438r
kCnnCo/D1uz1ORauRj18lI5LjVTwzbvlr/8he4+xL/Qp4kxe4/OD8Nv4fHxh
I9qiLctWybC+jRPY3lZpxCHQI/SvaxQrRhKeD0OUwdDlnyhpuElgRT66HjS4
96zFmpiM2GAbawwvmBTOAmtF3gpbMe3JvYT0FFfez/nGOMZLa958g02S3S9t
z7DsOXZB4lnfmD8u5O5huvOsN/sZ5z/jFQaTWRPVDgjlMQnH74Lyq/3pNIl+
icdntUIh2mjEFHwK3Z/IwfEOElLdfPOq55Ui9IfuVQs6hlN7kk0L6aw+gm+x
CbYzdt5Hwctfx/exLISiM575VcQp51tPIu64NoW5J+TKGwiRm4XW6y3Xz8BI
5IRx8xNDC4iAQfOWEpRS4RCfX9INyHu/m7xPoaWSmJ8pvQ==

`pragma protect end_protected
