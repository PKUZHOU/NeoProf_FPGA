// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
LIs4rFeyeyzCVaDaL+3Cr3bTspzicQrpSmwckbCP/pZCxWBqqCZSQEs3Qrb2E9/1
qcxjl6UvYVj03RHULlHyXr336t4uTfpzZ66NHHf/Bz8tMYxNrxMlPMEfSE/N3At2
9gastvwTibUbdm16zaqjp0MPapZy9Tfu7DpFGAxpNRI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 22160 )
`pragma protect data_block
Bs0TVJCCe61bpmQHzRr5UcsQpFECEEA+Y6Rj+TYIU/IBJT48P3lxJYiqJKvxYz8v
HP+F2O+59ELv0AmRNWUnIWnGyurPAcmVx2ywlPKUruDogMeC7YvGmdpmwF7i56pB
SpGLfiPUU0gqAqxF7nNhoK68sRnplIketkRu1WQudU+zr6j5Z8KQG0DQwxwB95iC
xq65mrqdEaTs3squImD1TokliI52imKyUvOU4hruELcI3MJKnpRWfLX3+tKukdU3
rgt8tFqSA1ErFrt79x2WO3QzCQ4ygUwpYOeieFTbOHfzRbHRkL1ZJ2gX6EkAJkxm
XN9O6SdZQSA1H9VMpaxp3K0T3zHbM4Ypbhc9uZ6akQDX1YMd7G/fXYcLb40QCPDs
QANzrbhOXWZRtqGHvEZZi9PyTLJJs+/BMO+AMb+1bo8BaYzIHsdTY9ByaKnzCtQr
JTrbAZ5fcwaf8aP9wM6FfiUel+n53JpmZcj34nzcqztI+u1NjptEB4fEWcE7WM00
wnJ4xRlDhhupFRcX5VAL5/ZCta0t+9MLNLJLXOWo40l2wv/by2M9OOH+Sow5Es1K
kEmvma9vmE2dz6JE6SuYvEoVaZIUXv8z/s1uJ7MVpaleRUDZQfy0g3jYcUd6ox0L
6sB4dSTwImeSE6NlOWMt3SI9Fx4jdfvEfYcml7/OK260rPyDcm0SOYB2tSLXLiDR
DhxYj3TcX0MepzOj39lOtm5eZxiQ2QdBb74iD6abfRt8EeVi0MDtH2d0LuyfrecQ
/PZTiOTY59G+O4SB3JuV+WHkkCg50aH6UDNRdl2TNZ1Da42yNigFqApXTlVCoVkg
VlNq6m/BogByMH/H/2Oq8U3Vc1AVQLIVn3QpMwYUHGtVL42VR9gtVUXpNl6LHkt4
10cbtGbN0wL5n2GUQSjEijYH5F6s+VSbOnVRaE1lMFxOxwDUd7wNRJUKVjv2j38m
pg2BmC6OCZKOgiJ+Kvm2jZC5vgFRCDkHldqYto1QzMLJdqgTtAVEvGuW6JBaplqJ
FpoClPZfoixVyO3s+FuWfCb3pnTiZJjDzbRYOt8YzIItyiF68IFElbnIM2qvjhhK
cWyVXQtSka3RnsLKQ25PmTtmcTiLAsW6aftGLcbhHa6g4HpGSCUsCHxlMulPTtJs
JQq+9TBzIORyYr93uS2zIF4aK+gHlJWSiBnFaMbWFdSoaF/YxsARleFrOQJQLZ0I
tLS6rBz7bo/NmtJdelpGyZoyzzei20/C49BJgi4e39AZBehzWOjElsuoJGLsSIGO
/HfmtWY+LoxEwuRt/yOQzzXcY7yeWTvnjZyQtxHDejPSnBUvZy8t02TJ7lEkVq7q
JXqla7l9LewwSST0xidocAKXWmwNiOx0WiExOYKIA7oU9qKsWoJdHvHDn4RUPu8L
1+iciu2OJr5AbGgCVGCGR+m597goTo8h6grl9mSlhT/swaQnXiigggxfqSetrHUS
9dbN3HTSxmW9cY5KvtUBvVg36h6H+K5rDcNdXVf1UTy6AR+yqZZNuP8cz5fWfTRm
xJN1nt4lobLU9P4/XGrzW1F9CAIK1qUtJtNyvze7OeCIUWc3aSYedgyudUn9hsPf
6e1M5rS6yQ24CAm4d2WMKjlYiBR/7Txby9+ezaU+UmbPcFKYUKD5qenwTVHi5/vn
OnFhD0SiG2PIhNKLE3LObhUxLyS7Q+oY9hzuyEeXAF5RIxnn/8Z8HwqZgsTfSomv
LC3k7fG7wJ7SIBF5c5TcVFI0IVu+wbMiZiYyiltWLGmrrBC8kRO9P4XULrTKhQZE
KqGSkQ8sCZt5F0Hs8Qumh3thUBw5Tx3Kf7pQPKw0+HlUSQd6v+0xUdDGRNeLcs3e
NWOMFwc7r2JXmw0pQ+SiqGL6vn5eSc2rt7amAZsnEQEbzNeBwLqFxPZamdjiScHl
cEG44fDUuynHivZeYcBzJbwOy5RB8l+w0YdnybIK4Y+0NXrbj01mrcFW26ku3prX
8ICYEqCBg7Y26kke+K1cOOqr1EompvH3Gm9G1q04XHZz4c+/hGJm6rVH7gBq2MCf
du93Jx4sINCTGa6PvOQ/zkF+PQCN6QT+vsGQhM2ATTBDuQjPRtT2m3/D3sikFzgB
HGQajwCCNF47vk7Q+T8ne6NA65QGD/HASVez+68+wOAmrqCPHCRGBh0G23/7kz86
y54In/NyWBAhKjFE+M5LvWqZalS2KYsB4lLjd9Lta/ZWhT/h8ZPFICxoDntBX24U
er4Pam7RJxcappBvA7v6erZ+TMCTGySw7952PoTjOsnXsc8VnDZbYAdf8RCzRg+s
BsG74ahIFLbfvTwoZWoUF8ZSkUBh3EdoFdlrMqIzjbyhn6a7xyUh3U6SdbeEfevy
sIxuPfyYWUrmQJa2B4WrgPZiz/x0uRu+v4/bbnvreVZM1PSCGcNOqO8/2qXyk65T
C8L+l77ykOTVyDpMwC1kIMLCGH67L2MfYCNTEs4ybzFm39PD3nC74suMZy/U+rvy
uHzIEDQiO6SxyvY8TSDqoJ00UAVJsDFdbvgIQ49euGgwd5gdrSR3k5LfV+96ZxL3
dMaLWa4S24l06/3TV/MdTj4tYVgpEqtSyYYGIrIyclLSkxqX7LvidKXk9TwknJTU
vra3+FyG2rsZOJm2qlfzr8DfQ3WWY4FZQmHH4vQQCzPgeM1xQebCdZiMw/UopOtm
qInKDYRqdB5vtP3CcUDnP7TFjC+o9mflozKhX4M38wdFIETRwNapUiBra05MAWNW
wfVR3mLNhXWzIXT5Ddk7AcfshIKEEX6fzhS3gbysLNXRAbu7ZubU3YgULA08jxrh
OvzSr7ZRyoeJlRoxAoA5SzENjV9TkS1Lek44OoCtNFN/N8Hh8IpsXd9zK/kP2GQV
85JtbvNolG+s2oBsh4b7wzFJLEPbHef+75/YIAiBHFunGyjFVLCJm0hOCuY8Q0tu
NhqKldm57KaxAYT1Ebevo/7P3wcWPFHaxGpmabhVzcJaZRAUJih6RnE921QIvGFe
obNvf0LuEhPDEICnQYN3NhYyNpkBfHZUVRhmFkXPu0rhLMHbyG9pF/ZEefSaEf6L
qoggWUP+ym9irUejSFBV50qizIeTBzQ3pEBk5y40R73oUBkD9OCCeApW9CWTQz4p
9JszZzLbGx1YvzpAFZz38C+d4gp0utGepeG7W4gDlbbYWqNVRG4RxBYWQ0jJteNT
UqdZqydBXFTuRVenT3XZnXL4rkEJoBQfZcXX+KZckODEMS6tMN+RnaudwkIKkHgG
yAMmyqegQzzSEM9zQhULzUxEs3C0tb3hHZtYFH1kEyS1fik1noShuGGNlrtgjYQn
ogyGBTB2uyjuxx/Av5sfS7cAa7rnfG1eK1r1Gm7lBYu8/4Qm+0aaUS/iXr1Ehd3b
STzw9qxtnKD4bycokPYiFqU+tKoWVsPCygUwDuAP6VERImJ+a1dKrg+yI3zc25q/
uItJfEedyJrRoCap7LwIxEWx7FdjXZ93nYhJuBKBuOCaoDlzMDS4so5bk+jb6Th0
sqEK87GaJuZO62c7uyn6sofViClBnMxDzP20ZSM7pgTU/1G1mrgpswHhrYoJG5lk
c1gdk9EUgspYQme4pG0AoYGEVgH1zFaarFeWZcN/v7WJe5beM/PW3Xz05si4ARY0
h4EerdilSBG6xo78yNsOAQwO5aOty2SdB5fVknyiWcGZv4WM6OpyiI2EAxBmKYTn
w6e11ewuKJ7nJXiunplh5GkFCZpMLWJVAozYWCqFf623D5Ey3W5dhCe9HRwyTIqj
5ctldpbgwbN3H5Jngfqderh/1qDq8gPmmR40QLQ/s55hLV3pqFlCfMoPDKe9++dJ
EwqHYTqfdGHpO1aeuQWqrUXkip5AYhGcPqf+jS2GaOYDfzpFVm1TBQWV6DJMPlZb
Jj9pCB/tJfm/L7U7B9GYbhIXGLU/Pz/z3Ki3PzbIlHgeVrZF1aYdhujFofp0ExfF
MvU8v6yOYF8It0RO4iY9pyemollNn9Ho86tg9OxuT67lGNXz6CypIPq3BcPGuBjo
cDqZBCjupsnRubXPKT1UVnnol2e2IQWRFqQrg+1c+GND4OTNwwsgIFwWoGe6bsdc
se7iHxF0QO5l4MJMMU77n6dhp1JGcyy/s2M+TS+ipn1hWV3nbLnfaXdMoXCK1Gni
Mml2O8X8w8I2V2KjJo+ZFe0T1LqUjawCq90hxfnUAq37JTzIlzpmOnNW5TWVgqN9
1nDxhhUcSJzd61qwOzNLMTrzy5owmaHPGV32cpx6GfvRdjwyu/jfV5j1NqgzYi7W
YRemPWwg0oXL+EyJi5hAnU5pCmAYmOgKT9mJ+kPyDrlWi4uYb8AKyH0a4jYN4hzU
7GD5SrIcGVPs0tfvVDvwv5IovIF+RcgyEFw9yniD4BgblGAxHkhfSvLYoSswQTrO
K7j299AfUC8nqeMepthm21GrqiSlroz/R3OvuEuFeTlHfgwduB36FY0dkSJPLD56
HuTmQv/n/AJPlmwwOJjyq16wm0RnGm/aqjRU/5r6TXeNQEM+fSiyAZ+wyF251yfe
r2jW3yFMYCSb02f7oDJO0RWUxdFUw4d1D9TeZe5ufaBne35mvQz52o3mUT5TFPtT
7O7O/n0Stm2TN9VSK75rducjDGPIGfzFtyMTnQ566gn/667BuQb0psHn0psmbJMO
PNsO0OsQOHgLBD0Z/uiQTWgoyqqePMWbbSmU74AB7ChJgebm3bzV4mWX3telUHDX
G0mfY4Fgo5EcjBNxQHZ1VViKE5edEFAZvxqtm294s7Ce7+FNzzdkMdTRxiIq3XIj
lIV1sFE1aQt4nHI9d5RHdSNi5GrOYrNQlhPbsu8gKXbcXHoDSvbNXOMgBNlDidBS
RqO8TtnCYJZqdiVhck4vQpwH0HoOH2s0mu6HNeEWXzo6jhozhl0XOzo5FIVw9iNF
JMXUFapuofW4fARglPzPDPMjmAI8koo2McO5wOG7ULX707K6O6xBhaVerBp3G9ZL
W+BI5pNkZdIkylpbDmnPqsN6K+GdYRcLrzeGs7sglnlyZ0T197T+zHzTbNnQX7+b
VMs0dgINfbtrtKR5ZJwe8M1kphNjGdFmWm1wkqqBePH0AHcHG14f9kpbrCOCFSLV
N75nXOsYeylDersRjCiCh3MZWnP9IYgQVp1ZCAJpfWHe7ESgDwbV9IBmGjgafo3m
fbNz8DcivCsQf821br5RO1Sfgskx5iraLe7mmX6Z/lHZVkk5j8ZcQOnqj232aZUy
+IYxz+h/x4ICdVFKHiteU10yf83zSwz/t9ndGRy901pXjGrUON+nN55wmXZsSkhp
IUuIqyCCVgNmYa26IYzy/SPHz2ox5aV54FyiOGGrr/pByetxlw4HdwwnnX956bfJ
zOZ6136Y3SL0wR+SBYCyHTk1OHjqFoMABAjjR68OveaJ7tmLHBC8yPDWClIsjCh1
gN143ImOFGEsxRQgNZ8poLddOwPB9o9nYHjUP2Sjsabx53eDh0xx5sFL0jsSk0qx
ft8/lCYHiwhPKc9Zrvb4S8gu/fQcR6T3rsysdoS4jCA0QXQZ1plvPxaMW3whapnu
7Lv7atoBBvb6IkXnCSDrxnEW5CwVi8PsarJHPqYari7P3a3l0VeN8RlnZz8QUFDS
M7yHq4aObr2RUF1tJw4HfArl9uodvCcBcsHpjo4JVfifOvZPiQzAZ+4Dqz2mOmkq
us+JA+BCDR9WHy+2ys5PcszcOaw8JVFBtoqP4qktncuWYbs4VSE8bbr3nAAY0Fzb
CSmvyBRs8B13VFJOdolLBHUBbkXiFwdIDrKE6fzaxQ+Is6chyof9fNs74v67cyIl
E1Hiaeo6e8XtNTV5EghGzMBvH+s+qlVC8/iDj1K+/heHwOjdnF6E4YKC7zImkjcF
hoYdjWA7fKZEz1VpAg/vErdx44ANtZUXYuBp11W2XnDFu1aaJfLvoJMdrH9VTJgP
RSFo9Se+FJXZ3/CpsUQW2KZWDH5uEQebnLoHMqlHVhdomT1apIjmcotL2Yu9vayK
K9qDHAHfj9PSiZhZg54BUU+656dzPZNSdwM4RarlkGvlRfOdadoD26uRdxj0yN8m
TB5xf7YgdREa6dtRq2cEABPFOUnln0EbBMALI1IsaRNx3tPSTNCGvyBwiVqjD3Kx
/Py+3d720oj9Q6iF5bdsitrmxQVcffDXmi9Xt6JYxkJZmc2Y8g5m1ZjrELcCswyk
a0qCOlU+aNlykp38WygSHxlZuJJ7OEPt4V3ZG5j7Ze/0iFaNY3CqN/yws3/sVtjB
GoM9P+O9q99P4tu386/i1n4KC/7/pk2Crd2n6gh3cLW/P9REqwJkPmsRrsVgeAsj
ovl8oIgQfHi1WkRxU18tVwrFh9dSW+9YmIuqBYTV0HWHumfEI39lCe/1k3q2GGp/
V2ho4QeGcJsAskcbJoC1zUITnJ7EgcvQVbICe4k+alPmrPsxhtP9ySMS2p0+w/Oq
etFAVGCwqCBzCYeP3dWfxWd+XCxqtmLJ52Gjj/g0ymMz0nwEIuoSMX66N54Y/WVq
/sLqB/v8BEBjBVzzR0yU6pv3AXZHfs3V+hOUnq6+9ZO7hL3Y2TMvrsJ8xyBZG0On
7ZyB9ZtQhvKWeDWyaj0zqVtfOV+tL6ON+nswmssVlEeTY0hFtfyNm7hE8LrUNPNA
ePw8nXZMlXnBCMN+nHKsE297p7tT+FDc2tKRtHBnUEkO+jXTlOPIVJZdbf26YWHm
do1l9rgjhtIOtP+KEReYdXhlnjzNYk35GWXJWENWGu9zRIe7YBhn+q0YBOXk1S6a
xhIk3oL5r7VRrJCTnFQwgl3McrnIfApF49lCws4ZNLVGTn1g/7zIpANQtW+z1dy6
DbzF98d1p9UevmOI31ZkCFpoY8IA+Fy+aax2AOCtpSdbmhpAeCxos2xLxyhBeZ9R
FiEAlS9WQNG+fpepME5NydOR9pdHDbd+N/7pHevmbZ7H1ngnQmtaxCzrTTcjnFtZ
C3xcApogNUXKBTMCduPm4PLD3b7Ceb/nUvSvcNr8dsmsAdtZHspHrA0n5eN/5sA1
6Fu2f4hLNxGbOoZCOs0RP4/P0am79ncMD0bv1/mgz3LZBe6aNP4qtCIZK3D7qKeB
OzmNshJZT4uQZt72FohrATGpkYueb/lpvYje3zhz2ArwaPbfMcDYO7G14AKMEjaH
H56aadugNfljrM2d8JyBXmxnjOft3kw/GygfvcOUYgjnOMJx/3UaCKIsRM2AIA8I
/ncAkoRZNqshRCZYhY82bQ5C3LtbLemrYaF14NSJgYc5KsWAEKtiwObxaQIoS06V
t/tS07gB3Bgs96p/OuVs5YTGt9ytyriPiYwJ4LEZKCDFKReKpGht3tXV0Nhktcn4
/YsklvmJRVw8hhLl0K9jf6P7WiBhg0zZSouCjvgk0/D/i+rx59UoAN9XD2s/r7Gg
9tBuTXnfiUwXHLs4eGVRygJRPpqkO97S7cSD6cbhBkSnMd1+Pk+/3jfkv/NfJULH
+yeFXFC0ChLjZq4PpiLMC/WO8KUlvun8fNfIjl44DU643nxaPfKj2YmUS3f3ZAiQ
p+Ve8AB75dpe2Yb2ckq9EbyEQiLIBAI9If0c3UuUCh6e3nStBi/FCOZmj6cSswc+
Y9vYfcBsDZ5OgdITWcm3HMtA8t6a0QnHz2RQfyrEzGqEa64Gl/YzF8/Wv0z8Vu4i
VmN6XCtPK9L1jEGzCVHHJTJpjAk8VmPgMjsfEV8C0ICFdgzGRfufaIrLODpqn0pC
rau/T78zSf8Nsy5jSLIbkfdv3ASzrvubpLwbLGVFOtrrxIxb8eHTUHHT+LByjdPg
vr7CF35AUqeqURNCFIPC/LvITiZIEkjwxuY+H6hDxaLZimva/hmnLgBrH/00HOOw
rc3+2Amc/UZVIUaGe7+4o5tWXr8JxvhrnxHqoKu8oBBzIST2ap2yXOrSXIEqprXH
22jDoRyaGYCkqP85/AszYXi8C5c02zzgvCDArb1FQ0VZRpJhv+9pFQiqXEOMTlmD
ONNwJXbDoeW1e2cLYrCtT1cAGkLVaMCMylLzAGXcChfMGLgfy2yj6D24GPKmPhBg
/74Tyb8/vTy8shKSLD8KSGMFqpVXXGMEjGDIMkOWOQV5BVrUfvJS+OSYjhtfzQBA
DLnMjarU0voBgq+51v1BNUHmlc9xJlO6nOlG+cwnZXkWYUX+bkzwv2N7zCSo2V/j
+G0UJSeOLAbQga+zlQwDHdrJDxTA6i3fw3rbrvAIdOFocgnBsLWwctBtNTQ7bNjt
vAU0ItM6rpIg6X+PVbX7e0evUCanhdJ4aCK4BXoXnT3v/wVHn7K2ULVb7Jq3kSfU
95PYxN0+nhnxw7Y6OgZiThTy2nSJWhE9yvqVWBpCjVhC+FAJouIpTB6zeILnJHOX
hoGd4/+6I3uCujQvqO0d5F2VxFWmSULahuPOJ0m1qNC8nNXLOaY+/q/n/ciUEsln
LOvfOB64jN8GGZGeTWNjOb4qStmqcWzEoThzbDm3uerZsS1YqSLpjxGW5V0TibxS
z9Y4IR2IoXAvItVT94l8oTySY/ahEcxcsM/dliMcrfE7TMmBzT4tsJQTIdy7K1ch
exUh4sBT2jkt2adXZUZVkCzlMxsoCsJlBRA3fbgNy7LGGQc4/oso28ZSJScUhJSF
1RhaVVpByQvfE+uPsdj4TZN+JyuLKYHzLpYUsP/lUu40FT5rn8BzxNzuv1mqRtJm
5ST2uOFdOXelmS1keIsiO/2U9AKhYQRVNKfeAnCEnqLc6RKTHr5imHM4/RbyugGG
Qnuk4wfm4VRojJv3oaA4LrVZTN26+qgR02Eg1Pup+E5jrT5V4CSqfIJGarOfWdr5
1oT9nmV8QKOM/rKCRJjZhmzWw9tkGds+us7J6cp6bUJwt10ibTWOvO8B4m0buUsG
CeBRzJBtdJte4d3EWm+ZmWXYsVSPGBn0YSqQI96bdFUnHOpngjMDI41zuyAKlgu+
t/WDLJRq4DmGmDY3ZcdW3pZetl7HE/9GGtUIdzran8ltomjQwgn+LKtBDZevhe9h
nCuJ/Z37riV8YoZY8vphFlA54oB6jPKfHv64dpPK6d3J+khMSjyNd5jI69LAzJuJ
lW//oJQz+W8nDFMGokmpDxgOoNqtrPwcJ2PFKdHghM41zKLagRS3btnAWhsnjh7M
QlDXmveoQHL0W9+IuYRVSTs9iEgnhBdUNOhcNm0nCq/RWXXs5gFOj32dYMerHYvP
931N4HZ+X9NBQM6miiCttZ0fJDiKANsCwORA540DYGHjbo2sW8kplFlNLbxJ/6Lo
f+3ocDwFAURFXpcJLuS8KlQcLnS5opUyJ66RJfhdDY0DIhH/JXgE9Dlbd+DFWtpC
KL6qFhPn/6hZmbjI50Y0f8LTKPMQCjm7Bwl/R62AzOhExqKgJcVe3kjpKyz5jMam
xjKdAdSyUOPeHc7hceqXs6O2qtDNJ9WkDazoMlNzg2qcCaaSdeBJ6TrARKocc31P
hl6UkGjrtwc/g7oo4svkfWRlDgDTGRAipWiTtNTjmpZoPdplLWXf/mNpncjRU7Vg
0m5XylRQvG6+g1x8K99DZTndhhn6tGJEXZR7jIZ//yam/pBifZ+jB09YTL0hDovH
uhJu3BUZmSN2HwZMQzCGD34U/hB2rxdeeJeKpTA1+6egsRCfYHbtY5Xz/8cdl+MU
w9A4aG27jXMIzpRItnA6wIY3cz9jOAmPXDdNInZGWUGeKpbBQUQxCfq/wqqBfuji
72WVqUkaD70Is9ouw8ed1/SlM69QsO4IfhAbB9IiemJOcJ/wXjgbmY/0TF4+Xtcu
x2c4oQt/GpR6qsbVdbuzhbkPnD0EaBYDlBZblOoLtz349NOwy8RiRqF81FwAx1gf
flIFpZv5eY4W++PK4HfiN/nKwGj+YYDp+Eqb6Uf4e4AwVYAgKj2ueQCfB0lO9lai
EiPPIbnWKnXgw6yEcFkaD080GUGb9JiQM3VkHnhbWazp+CT+QGv1kmmIQd48z9KS
tfNa7WRR+DgPeGLs3Q+cJXuTJVXZLAesGdxmMUAd4MojeySZhIs2CvlUNmCqxFsM
EC5fW7YZYlYIqwtlcCPV+WTyTASa65FVGIzisSv5pkVTZx7v0snRZ33elAGskJVx
/aXvCPGeR/CCx9pj4j15ATfLgai5cy5+kB64B/7IjKt4DsDIpcO3Tfpxw3HdixGc
LVpc1M9T1SAPOVF6beso+qVgWGSMyvvRtyV8pM8q0sTXznFg0WgSRnzWmtG8Ytj4
bDNGxRY4+roNfF1ilmhAsxb1+ES9tLMF1S/HO6bvjYRxlew2Ltb8DJFMdfHXMcbr
wWhE3gdRuu8CSKA1saHZcfJ+BCwpjjOzb5k8cciU7SCzQbUAdyTGVQlfmg9YtGHY
+ljrpiyeAO/IoSixARyT0qBHJWx5cfKxhf2nKAWLy8SlqC5XRSuIM+q/OKwCeyC3
kx+DwVuGWSDA+GNQfUJQdypMTYVe/rfN8pMSoTab3cUdXvkZozIrMtCTVZFScf2i
9frwWIwsad1F+tYPHI0ItNLV/kg42pvl8nW090JAOCqiG65/iAQ+VjeQkzlbsUUj
J6ldRynCU9ThNYO/YV1U82ehmqILHCiMykETIuONxzBo+2I44oHvtsmbpmAgu9Rf
Lm89m/UJF2bblRvOB/cZj1a1BNafyelxbkTeISM3PfPxpKaaqffvcZqwugOt5Wau
ntrnzRc68xvJO8ocUVW8M1iLlOcMo1EXDESDbqCHi3brcg8fASzkF8/0iQjiX07F
2X9FG1bSzxJPawuxEHzZ6zZ3ybRjYDU8NpQ4PKK/9kdO4Nh02QAlmKqZf7/j9AeG
P88MmPmtmBdo5Zc60lnZpbw0Ydj0OVgzoNlUFCkwDw6eNf4679hdNpNqEpjzAM3r
JtVQF1cDuY5lBKukMPsZFOKyNJEbRTH4F2HEC2AQ+YDEBWsRjI6CFqlCie5+Ea/Y
fZvtyilBLkbaEFc3PPoxfGmdowpw4VfvAIozrHUUzcvWTyWbIYviYuuT/jzBAZqf
Y+8uB2ONPCCJCmFipRsP5INRx8DcOO3qNq/uIM2fwopK44oEB1fYvR/2nND4vnZm
YS2hFFB/iDy5u+jBGXAnSrrx1pThmzq81NI5wsvhfh4EaoL612f6P9HW6sQ/FhwU
DNjxKLb7GUdr1VXEG3s+faGZFIjajiS4Ctt/StIEwA6btGy7IMpf32QD9Mr3yGHS
ksgtIVfBDEKvQiJ609t/D9AdNyXXKXhgHVcUQx8mUW5yR+Y56SMJhLW3KpTbwpUE
rxOWT48QpNFTUw2TsqNVAuj2SubA/U/rKXV0DYbNejesvve59JHpNuh49k3D7R2L
rw+Oco9Gq/A1RzmI0g36uouk6/WDJj6AdACo9xuJ9uhyiSSOzu33gllFSQT9AxaX
tIu4udX+Ut+jtheww50Hrvay3tfsq/vOq0jR6EHSMGK3gs6sWNwpxtkMzw7UHi7I
NQGv97l6jonm0x+vtOpvN2rW10J/T+t0Zwb27d2PV5ojO9zzcSsdeyabBtllMfcY
gbmqHXisfz/v4H21HqIfLg+M8iA7F57lm/pPWT67fT4GhvW1Sl3MErMfWEUaNy9X
4LUKC/PKNyTy9ycWcCeGGieLIL88kpet9CUB8rihQSq1ShgwHmZKQaYQkjL+WToS
p/Iw0SzWV4XVoMktYHxPkYoMzaB//nZ1NprYEgk++ixMBDHdSwR0ECRDuyYDoUvI
Kb6ArRpdthO/kAFXUkr7jRMN6bdGnBwIGOFCOhdWp5bslNgGjWtlZSIAYYMDmESh
XNdVkqANVMqQzaulC2HrLWm83Fd/Tkt1gAQBVwve2hZ/mLOYE9XQyBGJepc3gawV
BXXekliExszFPVNznBIdrJBFYErMC0Gh7jQYZ0ZUEgVi/BYnoF04s7D6U1zwB2qJ
dDFKRnD8ReMU7Ht9i4RapJ+G4EO3K3zWeTWKc/FsLw2LEeVPuzdSybjzG3LrsDPi
B8LUWAC+M1t++Y3Vc8NcPGjjcC/8p/8xJx7l2piNvrgUeSi8YwRGhwAGxxk/MxMI
ZxK7Cb0q6v+ZNw4BMqZW97Z75GVszaumIeZzeqZMzV05or/Qxc4b8qfP/p/nhsKT
w8RrIIK2ieaKB22batiyQYGftzaghW09Mnqh3mfVq8yeZ2jG8r4A2GGlfEeCZsK4
Ea9kYy7hgb7MDoWd8JwXT9hw2xTvMz0Ca7koOXnuTz/mDO5UIK7YM70wxs9gx/1x
tccIXn2EjoFWc5kkIwGWFbMYKc+uVlyDqXvl3molch7cklBcXS+g7ICjAf9rEMcx
H3hdoRikHrP87wYhYfVaiapkY2xXJD4NS8pqTlUhlzAhrBGsjCV0BQuNnOF+ItVH
HIonezApsSBmP8REjpo9b1CGwhjFHUPMd9aYg/LjWo1KTKbYMF55RdJbAmzQBRra
ZOql7GZfMneFRVjkUK/CbTPp/UnXaNHAfoaw3cSaxmjHk+TViMCItc5NcnapOYYj
U7zcP/mwmkKCJytE1O804pCAU4x0W9KHgi/AIxWKBTofZ4o5PGc+3jVz0JUAkQGx
dxDkc4tnh6yl1TBtywfs+rEcDlIbsWRXf+WcXI/HJPHdsaEKzOUouSw0aJoweZKG
ortQdeFUbZJhhjsIstxmpy8bbSFPAjc106MbKocV1aLui/45BUe5M9NYC7XPw+QC
akQp61mrSC6goIBaI6Q7JOKJKgtKfF3tylZfZ40BiUHrEoAL6ROHKCfJyD8gQao4
xrBmtUmJH4UwFG3Qpqp/IP+bYEiPsnBSjQES7VQSg1g28F0F7n6h2U0ojAMaEnyI
eP9zfcVJgpwQ6A2TFC84h3og9aoei7qfnoZ0twohDqkNa/INJVgLyTNV9OhB3Ckg
FT3unNqdtYo9FGYLgzDOkEgaAtZ4CkAFw9DkrtqfXNIV0I6DBP5TzYER/UXGqURO
mFlOnPb2rHf07OnosKa69iIp6DFudUUM7VjCn5SfLM30vtHhz64MO89IXHIYI8ys
hiZ196zDaFPs/j8cpvFmN7B3E4o9AF7s1BefjVa+rYMMI1hSfaQw08t5E5bPVixD
VJyDBfAqz/M3pcvP+J0R/RJBuT4TeFPYbzEHVw4jhbIiKbFy3UosrrRKUR3ItyUH
QLWbrICtcSb4iSGcQO8Y8LpuR8SwT93uNg1d5ieq4nn9NcjPdRO+9Z1aW/QLaVeK
28Eb0VeTR7SCViK/t5vrX1S2vRVsNZq+UcD9ghg0fjW8+c7DVcTF/m8Y+tLI0EG6
uVtd1TPmOuggwCnhUXESqsjh+uSegA7hHoZzZPn4EkgtshxuDV0zZz1nXF35G0Gr
ORumzKa1al89aQNIQHOzwDhHKS15jB0eWxeizdqPRxfxg9t0y/jZSwe5wSnf185A
Jee5AA0QjvVzy1OV/fsMrzpwR8vX/tQH5ZyqQmNM6zlY1DCr0KCpS/3STUoPicfI
HMQiXVZgBAmHimKQ/TtOuJ4l7nO2UqHBjioCuyoBe50ded7VP8qS4ZDPLNUY7TmT
lCyWCcTVVW+s+R5NIS+YkbKjGgt7b8K/reNv8XQdM1HUWw6iODIV9sbZVssG3h5x
XwP9/H0+yW5St1V2W9uzJhySQ1SFZjvEJYkb9EDp1qImtdEHJzIEifWvT9osF4LS
trubYEC261w+dLFy9G6vYX0DfhdPRzMJjk94e/4v6k0tluAy4PeDFLugKrchn7Kw
Q5Kn6XOJ0wUdvq+Q+C8fbDh4Iyt1LkRutdASdJzGyaBa6ACV8VXId23Ck6UV6eM+
PPluEemDj+hmnSSHLbhCGk1hhyDYoF6VoR5cVckzWGjEaqnaETDMN9SldzyNZ5Sa
2il2mNqGibWtKFrot4fqvaJ4sgRhVHWrSz0t+np0oWnNPKhIL6MzG9hpcJQpmFcY
ldzck9uMF3nzN4tAoi0MNc0uWt+nS55WIpL4JxL+uXfxQQAZ3HhsURg4qtrrjHin
QktQwL0YZy1eXtCvRmiPnOUIiIJ0arWZZSNXl2cBkD4xoDpRNxTuLWIma8625tBR
ZyCjQArjcGCOn+oCUwzkyEH0Osfo0ZAJ1+DK78UTU/iO5EUg9TdFJrOslGebFEQI
JgNRG7K5ZaM5uf7+i0hP5LAxyW7ah/MERzBdlJIzjk3x1gYFVi0r3veKKEtrG3sz
ee9zKRyIwweqXcux042y0IyaWa6FffAO4ztZx+/684oO8V7JeiFAP7NZGj1IijUN
d4RDY6JX+VmsToxVt77/bQJPRke+xnmBLGnw+ppN1aRQdqtss/wu6VEADEZIiYI+
QEcypTs7b8TvIvfZsJ8+xBEojJHBxewtshM0vs6tDs7/HeME1td28o3JWxLsYI0A
gcF7s21qs9NdYOgpjGiS3J7TfNoZ8uPzTS6DkSPVB+xlZ3fAvMnXy72ImQtYLMYE
ouhoZmCwpGHmDbQt7R6f7aJ473E4UuDcX/Ar+Hoye6j21J+R5Ki6bmedce8fK08e
s/6nsh1Vgcmm6srTBYnTeo+42ox9D01qLFGfwn1Zbts7fymbtTa7A+qv5GXLa6b/
/QXCXEMJ7MgWaw+xbj5QmN8fg5WYZ6rUHzVugip4CNHrP2ed6n/Qd6U0lM+5TrAP
EdBuSy1jqf/Jh0VYVY4o3nC6xkUwlgHmgrpaIBmo9wgQJzwobzZgrFWbLZNrLPgC
pmtXkbtbwEO0kzjcvHKT2pSV5z0wSaFCaCF99pOkcbqthmPJxDNjYlAqI/JbaQxL
eNf+GrmfW80kUL81V9mWkh45NCpT6rmQwM9ZBdmRdijUjx4xiedz6rT8bCQCaCip
yjK0pDQ1l9+FLcrJqZzat7wM1IIEAxjdK38hQBlzH2RgRqR1Qy0Pu8w3VSAHQQOj
Ytnx79dwE1LitjseYirzPnKJjsPjdviDqIQR9mb8xVfg5FQtECkQVryAGwVUrJrA
Nhq2Nu2O9FRlxUIVGJPYQyMm+fJgbl92qq9OWurvRs8L3CaVgQcy+FOQj4gmWF/9
r2THIUBH/Vtl9aX4D5XBaeY/J7Vrqj/nk9F8RxPhZMbJJHVWlkHyjATGVZAgKxRj
dHrdF0LktRLC4WbnRvr4LmnVX0h8+waOEkiJTKllJsGLIgTfeGVvsoIhpMAv1eVp
JszUZfpeaAV1H8oRgeBwS6vqAH5PeUWNu3szWgFFHJlksjOq/lrxxOLc51xAth3Z
aRlfWXMjF2fqEkJ3ImC2aRSYJe3+XJJ/1sFkbZt+WLyphYtSaBnC0SwuXWqReLfr
e5HfRhg48V9fGaVtUnvUov4JcfNEeGqJCkSb1OcvOiKZsj9S5hCXuSEMPREEfd6C
EzKvVFIrMU0P917iD4F9K0YWRNlf05n0rQHQHDfpNRIlOL5KURXmn7lOAAKIifEt
n955e8W+g11IcqUPCKHoAcDMI8jNigammNT5uJx3z62+7wFGq0g8u5VDxNvq2S9d
fXNafFbTsnsgSe0TKM4pvfuzqatZbdR8b3gXBh8mFEWsAZsbwLnL2WoMhexaRsbz
pc3AxUBka9uRtGBlWI1392B8Q3bp/qd6QLRcCswZC91myXtv6ZWtEuOJPhdBCTD9
5Mn/Vj796ErLRzXnOV7WqbVYA6I1qJSEITjNM5OZSIzflHyVmQAlKiz+nJ749Ibl
+cFhdzbzTG69ZbM3JXq0JrwcNhDEndqPpHP5Ach+V7x7J4KYpn9bG/LdDYIjaCST
eHAEh+RexRr/cEhZEuIc8HVdcU2rppEUXeds8tPHE69WVFCNBVVbQqbvbPCHsv9w
XG+xroMN2yVuFMhQjgCe+8dgfzAhiwMgj69JNujOH1tl1Ot3VJlNiurkWb//EUJp
MYs2wP+ZEtgzGkgHGw2P6MM/o1xkbS18Nn81lTb32vTW9tYZWYzQp1uZ0/gGwyLn
ZErQEsy58zQnEDxc0/S4pX+aC4Shj/F7hlUi9k2viyexWaHDpXu9HzYdF/vcLXJ9
oboI557EbIWM9RGX5XNHWe+JF0kpGpue8MCMxaVDu4uN4YiwqRjmHGmOlIMjDY35
rD97rYKqNJCPgmmKHPh035c9F4nUyIldnkTfEn2Ap0zArFcBQZVe6zNKdzC0myhx
b470Byt7ByV77QoerBxeW7LUv0OlaPQr6dFwgqSnCDKgXv2FDgbVD9ulL6s2XADa
F8E7lwIn9pkAfDnRyfItc3uixSysvGi0Ul93tRRq+al/TdsY6xl5zRez1xxXVlnU
4QaMt4zCvOF8jNpYCmMfIcObZw3358cW+JIPnzFedF/hihxjpHLGeQTWGR7cI+Wu
mxNZ3VJ26UWvszWBNmoqvnkTLF0zjsX/Ss+eJAoDruA8dOOOD52AwIcUUgauPvzI
UaGransXU3caSPlaJ3t0fPzsrrZbT4gDDxp9eUwbcomxpE1v+hzVsWWPGSsMlsl+
DSk2K40MmCa4Z/INYePe73TJ9mLyvz99ZA1NSiS9dRlGlDBlo6rjCvOvLvRbN/Qe
UVCu1G1TXpn/66UhZGpsW5iOJ89zenanXk89mFBsZdxQ3edHgNITjYALThj6/mrp
9bQfdJiRemBJXwftHp64MM2WtfOnNZqZKFJia3ap78WwFovLPGMIG8y2Jv87/U9K
loNWofd5Exqo/8H6JDh99P0MMDiLr5BJGxuixQTPAR8nNTNEoRrACuZj850rEet8
w9I7aaYD/3xr7XQuyiyEtzcVtgowx8dbX9fgdTK3YIlS0z1IC9ZX/aHEMr/FoKV+
38KheRXyMWPQhalQsCgDa7duy0/BBb9Syhgrru5Zl+GSpiAvX+xjSMHFfk28vFVl
7cuKwQeCshOaLE7mZq5VUn8YGlYL4wihvamRfBQ6rYRIo9IMBnY47jfgKUx/tADt
iQrNgmi26y4oLYdgC6SvWZ8ISveWajTxIwxW5UIIMQ73kt07B1WBDC0QYGKiLX1i
Y9/a8fZAC+fLHXucVQX2k5Lm0dSl+Ruu5fsYG3w5BfFvv4Mn0JEAmQKVOEL3jg4o
Pe9Tqu1R/mlTnnAME7sbCXMkRxV2IV6MiKX4Y5dfHdlA6jT7LAIiKhH5/jRdQKkn
ox6CmzyN9FoZ+m8xzyC0oqQbWH6yeMfL3qD42Sux/7ZZtjukZIWUwPxD0IqRG/2C
5rFBYktlGMGSwmwcZb7jfmDwxK+AP2rl6fuaknL/Cw4YvrNDO1NMiMPw3gFtBgtP
CZngqkcW/BrXuv1857QSuww+rbHXZIUBlLbwp3duzMDVPzg3aCrNfK1RbzghippF
7BfqzuibmMhMVwAg8Lh/xX/2bf5wBgfDPa6wO4GWKN0T0ehGI79Z8py3yFgSg4xn
/GLlnppLDzRdJtmIXw7DbAJqxZSd+sP2Hs5f8b5T4E3DLYyAt4fNcqxxdVpTith7
mAJPtHvagvtuKgyyIU/2ImxZ3wMYe6udlb2v69oO7BDGBDaMGzpNSKPLNCapkOfP
RW4LAK8Rp+/Ie3k0XtdqsRdqz1KKT5Kju5WwPyjpb7ggVRLGhNs7KyTtZorVleps
0kEDC3jiL4zwgcL+WGv/R+jEsctzCulx4Q8Q7iF0n4n0S5s0PassI0QT/mPNN3Q5
wdp5XYlNU6FsLe/cv6HffWwzmjHVMTSONoDyKSCI5CAsF+HDdxhp/1stsmiAQSco
NL3RVaY8XUXJuYlmWuGzsTIp+8nT/AGzhQZ+SWKVuMHnnrqOZhH7UOwPtebBF44Z
YqDYywQiq8aFRMJoU1Fj68TmpaO/c9ObYt34AOcYkNU+FCdCF4kKs4Fu90BlHA95
SkCXaia4j4+b0CBroGomtxqnxvAAzYsHphmEIgsGoZ6JttpkVP7xQV5jxj6KBFqy
8ngw22uo9c1bWCEoyCPxnfbzZIoVjFzEgQXypnmvFhF9S4TC70lbrN1bUtjhLZhq
CYL8hsBXEdc+5lkCUHgtURnTNB+AwU92Ps6qJG9cM+qrCwTkwir+aeQiOss2UG5d
HRmRl2j0z0+YisXVz5DuuPzZci2TJbvizhmAd+c/5/xWtlhBVkVU6Qy97TKxekbv
JagO/70lGMjYUROurL+9PQfqb8lG2X7Ob9fpQ5DNQSvlJcr/+jv7WbmNAC4Fol2t
xobYYMI3RE6w9m8ENySnxJNT1fdHHDD4EPAyKkynAIlhcqyTdr/INL0JxRCBQxcy
ZLkiwQiJU+y3pGeXpegvdJ6s6BS1qKbvrJwfEKxPpeT7o6jJCjW5md3bhNkFSWcq
6gPzO76lriAGD26e3X/0lGOlfttXzND3jQQ8401yBnJvkIIIJz95T0OpRTuEYxwZ
h2xmbftbuDeLzQtgunjiIPteguAmNt0g9og8rLm9OffqDnhKyk91T68AU5tCcl53
KQxPGOzuVyCBjRvIBnfkBQMflO9tdfFQHlPluXPc3pp6BX6WYYGwnBcsVTFMihIV
+yCNLXkXuG9P6E60J+vBxZNTu1wJ0OJHukE9PTu01syVJMOMzSfq+1f6VFJUGHtT
wY6F6YIW5VRsK87k36S2ITp5w8pDzLpI/feG8uTCokksFkctIDkWvuORjMPPnetd
ZTed22DRiNdbVv06m+mcw3rOOzkaJYb/P+cqMS5TNrehkm7xWqCuUiwHIgtBsIbh
XylARWVDPweY1Qhu5COCbSz/SIij/PCfu68LcA/rO0i0PofOzmUN66lWMFrPo5Nc
prWdDJkwP4cyQZcuKudFN6ye451uIcCNcZJ/gRiKhgZiOB/zFUegrqz8aF1/sKL0
9Gkwlq7dTvVbzbVJjldiAtbwVXoLxWo5EzY/c7cjaKL51XkJ8KrsoKeAs6nkU6wU
oU+SAotUPSZph23BAXoDKn+VHG5LfNOe94FFlp+kctwwlOmQskyHEuDVSlGgnebx
87GGcU1HkDpbqVj0vLp/reyC4Uv5bYupavfTUixJm0mM6kPXL76r3TixQ3C4WfUH
W+I/rG9+PTwZRNQgZthqkcZVsiT75x05xS3W0V8SrdT8Hq1ssRc/jZI3yVp+7RgG
Z7gp6QqLDWgbbQ9spaNpi52+WNNBiV3r2bHZXT6/CYBOfDQOfA3eGUE4z26Q2+KZ
KyvBciJBaZXNHL6pAeU1JZ26+9Ec/ER34fbQIl19WZw85VvCn0TJvxuH/BMSr7tf
j0GIO0D2Wh05bzl+GHJOFdSvl+uoKzhijeg29gCq9iDZAbioG4T12ao0kR9gWaae
LAuFbgL2251whBoj0O+DfxhkIk1Q1egS4qaC+ICZQWr0bgquC2i4G2tEH79WWM6E
UIrF4MvOQ9iMFNji074AeS0o/GaMwaKx4XpjVQfFhkadKqGoZSeO7dSO4mtBHRXj
TK/LUuJQkJN/wnkPcZC56IAKrUX5MzU6eQEeIznHMmUkSZQFEBs9eTWLcr4ITbI6
hpX6kZvqfwfIMqw9yXGX3EWSCqA84GExKvBXZ4H27Nny8IkVl8z37GtdBHxLfHI+
qNrc8nO1zFr9YTpAURCUPaDwNZ81YfDanqdNfvIQs+nN6+XJ667uIbI1RvwfUSsa
5ZB6PPMKXaUHpEqT0EeSOeT9AvbAnfMVLuhmPCZrudn/DaxVhnam18T/rSdjlSPd
Vc78kEBtFq+BqpIxME8+WSElsMjTnSvVr3+gilaPRMNtNgQExyF2ytPKAwYeFQr2
81+P96cC9stoyu2SPeRufg+j/eyieXGI/HwdZi8PzcNctudOAEbqp9sVePrVORDw
ihuMNp9PFUUte/wjaJNUt13cFzYnqr+RbJVLzCNgxSNfeggoW5nkK5U84JyWeZOj
1S72j8ETsmPckhEfXpY7KkhX5kXZofkFmdVJXLcO4ccwqCSkEnarTsw9P33233y+
lI9VXUG2Tu6IsIomA/hPNlDtoZLrWJsR5mYniBFli/NW8Hvo2Dh8if5vjl9/gzLf
BjTgOrHKjhg082+KD59adHeheonZhZSYqsIphYToDgKggWBImecoDnjq2T27rW+o
qs8SkNzAe2QuMmccezwXxYkJtraw4truU0tlyq/cirTQq2W9SiRm2AB3HMKinZjb
covHsTnFgknXjsH4Y4iaTKHUqLiHsmIhD4YujeCt8kqFBPhxpk2odhEUmgyT/eJq
csRswnsXRLGxuwzDgD1mlE2e8+xvTJf8SnUCjoMsr81TjhqKZXB3hhGBEI3sD/Jl
HHXvP45D6MpGr57N3K5dRmss8Iivk75/vuTAyyJMJmuHQf09s4Hzc+o5P8C7n3Sf
vspYRXcd+qNrQyNi/o9LbjqWriYgwekvQZ2L24n50ijqx4SMWTzw0S5R+TtzP7bi
65wSYGt06eMDBKkMcGZeD6A1epkQynckCXZxTgaDtEM/4I3WNnkHR2oGj5OTlWW6
A8ka7GTOR3+TP2eXaa1WxDS93o786Jv2p3rEOvKoLmBxSO/GQCIRrCmKsoHxt46h
q2rueIYVN5W/nG06nQtw8sfZ7kgvREzcBlcDv0KaZho/UCtnIkdC1grBKh3eQz8u
k0FFHZnpwdz0cl02J5Dlznviq8b4sITHZEEreukC0zBkPa5vPG3gZccxmzeU8WMG
exTB7chwVcQA+C2ebJC7g2BUmUCFPYKUij5aKW0E7G1gGrFQxKTAWaZdDj5Psk+7
o+0vybLUGrIerEA1uqolHvLwpuHLEJo8WE1gv9CP18X2VbnMVZ4R4be/+YoUKtl/
Hr+yALHMrsEAKhBCRYoMdatHFACy2yJ3v3tMVPCnWfZOY8+53THi2/CYp5MlcqN/
dO2B5BHCzPl8pFZYZfUyIyMFASndPZxLJJhBgH/whWjNEgZhs/EKHV0ms79aFWED
kSdhlR3cyE8Ifnnqmj7hIT9OEueVHf7EJU4UUFwj8tgFxxvAlSlazknDIV+L2fu4
XsU5JCJVElIuLYC0xay7QW60Q1Q5PXakULsdF9vvomKjfBuyi1an9dbbAKC9BaGZ
OOj6tkvuVt1lSOGmcI3JjKcxD676zK4SGM8u6dYxmT9Ya9zPZvhDdzOQZDV9nazm
RMxd/WprlIWwmcGIYA0P84QxQi4QnOC1gJUQduU4fc2oaxm73pNXu5qySSqXi0dW
rF9mQCFdPV/ycqFfQfryb089Vk55OA3rk0CyH1uQ9LJzZ9z+zHp7g+CM2U3JhVuI
Z6+rTWZ8OvZM0psT6M5u6CCvI65owl8BA/D7s4hsMozob0IFTqxzQyaGwuOInZsd
HHUKQDV7RKpT2RbhC+8xfSEE1VostrKpZvff/XUdldNAJSCQ3UtsOM+T/JT1rMXY
vtqXa5+Ae79MXCb/driBvzmvKzgkphJiRhj/na1zK1C6eviz4laM/gqgyI2cEdwl
EdVWnWKQO++8GQOhup1eL6WL2eF/CKDb50hgHKoFBJeoMLaLYn65NJDk/cINU7h6
c7TIZBP2JqrqXkiL1w3eLc3DBEbW2+71JJIZMkp1tS1X3g2PsY/I9EtvZcHQHRZk
0ilhqMTjmYaWwCKgIf5zUCUllNfDFNLQQRGgNlGwtCEO/R2xSZRIsgnCupvg5pAa
/PX94OhyDCb1E4HJxmqJrz/cSXuF+K8KyuPaU44EurE4q1b3Cy0dLxfWnTB/n61R
57jP9qezzNAj+fWKHJzBZqqKVLFHWe28z72QuhRP5ydfdccffSWV1Z/VGmX2uIs8
HRYi3kkp8jF4ceIz96APKkKAgFIDh/pdhfVvlDzmq30jdzvS62DMs3VKDaMNzSkE
jzX1Yp7HH+BKgvBuvlh1MA2xFtAoNINqqB5ylzwlnR7817lpIKrwUJGhG2udm8Js
I02nAi6o0JQZoBgbUrottwKJeNMd1dbYU6Qgx6nBMsbnaDGcV++iXm488IdPaFni
JNqlSXOXiuGz6rZyBCMovP8FOLwjz8P1+mL10MzaDS6fpyVke1AqLCFm4oJziYOv
FyR+D8OB51PA2StjIcjzXmFljFUyJJN8eFBkMi+qZoCR4J2OnplNYqvgoq+yOWEq
Ad2pGiG2GMFcfHx0I9y3tuzleJmPvSX82gMLGjS8TYaozgywy258bRRO/vr6NpSO
1EHFrOj549PNGTVrXYOeI+bRC19V67Wsfvo5FnCsd0POMMX4zazQfhXK11+K4QCZ
YXzuPBCxKzOP373TxZ3ysnCUuElWollGI2HNUyAnpHzlKI90S5sy12mungCZoQC0
uu4vClFKy8IYTcrEDskiQ5D4Pn4TrePDgouwJBnxO/plu33MG8Ql52VJu+5jSq7x
hpCE1lP13euM3fxTQMb41RJyHu/4PILYZg0v+rTu+sovYOREOy8UwyDjrya96Cow
GWi1OUo4dUN/5wWrtDd7fggw5o0QomLfxa57EvucOR5zMN+8HAKAEj3L/Dzru6mU
kQLi3y4cHdmFCQXpAvZJQUAPErG8O4YlgkKyd2mczUuJ+GBdIDOU1A/5UsdZDIUL
axSijEpLPhlMgOtxdAipmxDgU35v4PthUBo7x1O4pJx2koO7yFZhjxpKs5K8cSLX
HFd3OVT1DOItsmA6ydOgFw1shSncPKRegLUIDr+PUCxSV8Q8d9PgjGpIDtgWIRiY
vECL9ouCf5A138FjkhDJuq3bQ2Prv0lrX6f60l1ZWJOlOeAWi8TrMlh6sHpb4PV/
xqoTquoSRx7Tql9usQl4DGj1Y1jrBDAvdAwBvav/ti2mUKmyB7FYmvrljU6pbi/R
cNRtQlKF+PgNmXL5YCHYREp3Q1LzVCVBYdU7Mog+5PIIdElwbq4bkS4P2+sliz33
F6UM7i3VqUA0l+7PcIEcqXoEnSlg7gNLAOJ88MgSUGxt4jImJH+ajpJg7CmJVEID
9537pA8BxJXtwjOBt/eyx8nB7xxeukAIQaiaHh2Zj0Ir39cNcIPiOL333vheLhIc
HcCmuOUOTxVFxkA2eE2W9knLWGCOKR6GqF3GxOWkFu5VrdbA71hHCAl8npLBbGwt
qRo3NeAjsnx6a7TlqXYbctYJTEVXTbSJ1vIBf8+CdeY8W29zGKShIJegixDcb6EU
3ms4fDHHkcMcz2fQDbSm38rAQt0aE8lP9TEpnd7brHB85RVqJSiGsFY3v8ZzrPft
Dyot2+JJH9E93nuxegQK41xi/BrnyEzRG/xk3JoTs5V0382GXTl1gLbxjxSDwC7w
bZu4NfZFqPXvRjlIQQkh+I4VuV+irmh+32LMjRTHNaQkLZoOsYyCn8bo/ajTcxTG
qUr08LcpAgaoyKDWYOrrChtQtwbK+TY46MH7L/s9PSPCPIDzZrIu5Qbxphw8OTGA
8fSw1YY9gVYY29nSSVAXWUYOkcT87/VmZl1b/YYPFRWjaVuwry9klIvSDC9SsfjD
CUgiS5le2jBamA+jyJiN09lBQgXPPjt9LbbcQxw6ydw8OcbXLLcV3nG9VdNjocmV
+DdiCd/jZosjjybhmG9NFmSomDvqIy0qXu4MT69trGSWLAMtpT4dLeKgeAi5YvlE
0XohTEg8w4mdhwF+2XwD+TUpocuqdZXEy9wrd02LFv6Yns7qI9QWi9vMRjt9uSYM
AT9eAEgtXFSYdfPE1SxacKy/44ilHeV1m6lIDo5SYTDAGeE9wcamocjZhVytDVp3
we+KkR7lh34kWjWEh/wZQTgh2nQgtBxmsyZxgPJyNO5MpDKQTi3JKhujIsWoV2xv
lJq9mYTaRn17qkmH/J34Ek9I3bM5EFgsCFwXMYtexyS8Hn4AMj949SUIkoZ8rYt7
Q+OrCPo2ddZcSkLPEhXGqJZmKp638BroreqDp2Mc1EEH/HgSmcKLs3mcX3XW6d1K
eK8KKAZ2haUkQ19HcRLSHWDDglrfIbkr3C1k2vpgxj/NV5quFDSK6RGeNTd8Cw5+
9SCFQOWLjaZsCi8duetFU0skHPP/hCcPY/Sq8yarrksBpY1Us6AimvD7AQVhIOID
+uLBGS8YyR+ksOqnAlPqK5Z/hFgoih6NVJP3OCYIhnE+aF+18LF7JviD9Oj83ksr
bxeN347Wme+alsOU1evItCiEN+gqxs34qeXlNpMdSH2900KPXIH3oT2vimarNq8P
+KvwGtCBPtLYo9FxurxNFpSlxbzSw4ECHkZMG11ZZaxsRxlJqOP6J+0jaQ6TUVmd
qLulJqtbk+k+ECPnvfD35ObLQPyPKtnPy+U410wljOzNhtQmzz8RzXBgRHs3TBnj
+vE51QklLTjZod1/tMEanci8xT7xW7B5pP7lk0eXTB9eciJ2YR5N6oZRouagE6My
0w0ttlziHG3X9qUAMXVn/167/iSQyL2wCk1wlc+c7UVDmxZ8zvz5J09kJMUB8mxD
V1KXwxH6xXizEFwLw3XX+bAUAj79ELGEZ0PLp+olzs80oKkvLbicH/wEoQK1JHfS
hSzpIfMKzE5k5kHQ786pG3F8Y/oFzUoT79YZkzf3S1wqgxXJnMsdGn5TYPWuvSON
IBCUq9fkw1MhN9pbi05EC+g9J/qoz+cpgW6Gg81A0c0Ps6EEK4t1fStKv8BWvpGS
qAlcNRCxccwFdd0OHXUBnPno/BtJ5YO7LUewNmHaY/6c2Q3w5sCCufoAZ+6z7+lf
rNPvYnVdVYLPEWD66zkGWOxSXzJR0R15r8RpBqKsYlsbE2dojaWSuvPJnnARe/su
tmIggwYiV/nMNrNZfO/hejUNeCQJqqRGTNmsvtK95OX+TrSIB3X27Iswb117a/7s
zVFIMvnh890Z9ad/Vtt1niWluEaL5cgpeOAjKx3xQhlvVDPohu7oSyLdTa34VXIk
EWWycdglFBlERMAu7aOrl0vtmMR4BYfXBHLEnYiok3W/2oUvycuqaIsO/L1J6TqY
WE0wXrul/ENpDEcMc/B7LGcuQu57i7REE6HjtUf+C1v+2dBFjRHtyyCEq11hhokF
S2JbY2aE+82AxVH1YqxYKHXX14XxHxts0/V6JXT4zV8uBe2Y1epE7wgFu1kA0wzK
1xTRA0yKqlDHfcr5FoNShK5/3ex+wuIKJ2mUQKObWCmdQOFlABm10pD9u8Y11gH2
xjjQJzZaia7yMAnZzDvIAmRcFGnAakn00MFojjL4zywDCjY622Lxqua5/8BTzUZp
J/n6j+CL7gRAjApJp0AbZHSFLvYvDilhvS3zLk1FsS7r4/r1xjC0NUAlB3moz7UL
1dapUWYenQiRvsMZcGq1xtkCKDemBj6QI9mdI1aCAYvKp2ftIa8FUlw6egOBaADe
gV6NdBsURJbyazpqDQ0rRV3blPNHNh+ABTj23PNA0mHCJ4Fq5NFJ+8kqiL4TCB6O
/zAi/K1yTZobDZrtkxHohWYAECS166h2hUHuT7NsgexxOEimm7dLHI8ImwpePc1J
EYbUS7F8Nr2MNQBj8swbUUWN26IMzTB5Du8cVeV0j3N49/fSFBjJtNjAcgbuFMc6
0lS7BzLU/8edbJr0hEZyPZfB89FCbKfs1NtnM1qw6iZuWA2nt0tt68/N2IzGhM/W
4IVbpRWrQAifV8C/pbqKwUmeQ8uRDtzVErJz6dQw9fUXQa8gypmAs6zhNvqJ/F/R
nVR1EFto9cEQHk5Ya+kR/xfueGU6c9crYte700DSzzLSLmdtN7WTrAfhobNON/Ee
ya5fTWN6ufRP8wNFfypkwYATE4irbSHUGp/LN+BYCeobR/8WSIiLKG6iAyoCf+77
+tIPFBgAX8V5hptVRQQwd4068OB/39Y73qi27ovZ+tmfile5uy7eBp9Ynk+j6KNq
UBIWlCcOzK0zj5/rgyRe4OKP5NfkiYgMzof0NU2aCWJnMIPfHDpQ+Io6MUks4ecj
36m9CQO1COJ6Q1uoyrgDoCQWl/8iH83utjAcrbfeTohjaN+PjsE73VcRXJ6x206n
wa4uEI8ztwz+RjPcG6D59NMyfTXxdfS0UerHAhUFupnjsI/B4wkxzfnt1SDdxQc6
adznzYuoykB4ZiNn5/iNMNj7Q1DxIoBAxgPgkg2ceex3rKItxAelw++hWzywjhUN
9HY9cAe8Zr/iJMBvoeIWRw9jRNQE889cUSBgP7xer5GILDp5i8aaP1Vl/o9rYKbW
55qu9mh+xUNVdwmWwcqZw6x/YemFB3L/ujgXOi5oRXrmhiu5w2Tscek4uOyvf69L
+XQDynXKzmV5zX4n1NoY3wAZsTUc9EcgncAbtqkFVb89WXySjBBUsvMV6su0rKAn
PY2axRVCRfnf4aQZpLs4L2W3foqs2ee1sr/tJ8s4YiJ6rCy5ra1HrfY9vfz+vtfr
qfGhU+VxePhKCq9/3QMqdXhCtY1TOjXjxfVmJT6dL7FAUOqIsn6+Az2UiStI7Jhm
ey8HppCx5cP+DcUdU13PrAzunWGBDSk2R95DpHtg5Nng47qH7M16FQA3JIQLc50G
ZSEi/RRO4zdYxAivtYOoi7KIWYRR/PXCUisdIdMkvK2s4OV17o0WDddmaUCxbojP
eCkWMqPZEPMit8GXk0ti+q/Mi4bunu5E0lCqwGXjgparYhKS2Ryp+ut+zZUBwmjo
eazEXWKJyDYhfJ7x1WJBSDUqe1kOqfPxRPAj8u3bcP1VEV5GuP/A7o+oht4WrPwS
GiO0o7E+4eYSFGjiYQpa2262LCwMFi4CWAISzZiivImXG/VKSHY1p9uuju5Ophpx
Vw7qKwr5dBCJ6dnuGLId5TjS0fFvWvHm/efQAmPUjiBGa9GIzPIzLergw4HrJ38m
1hXDAXxK53KCOCaQ1lNgaYuA00JlUtRD+iCrC73VuLvYWPN3F0dXcw2VlhzheSru
26p1PcXXievTfouWCFuTvPkjkLdIAGmwSb2rpYBUhNMItpFuIVPt7hc5DIg7CSYz
GALHKWFomfcXTEEOil1p0mJltyUwf9qus6OGQAi5DwrdZk0cjwdZ8Let1gBjLa2w
jhyrmWAj5RDFTpXVnia+h0iKbYMIPTdu0RsEguu2p0KNNuFrLBSk/yMNzUrsxTuL
p5epSpO4OItXdsufGKdUCK8Ok04Mnw1um0+7BH6RSekel3xpFVqu5/nDfsU162Oe
jUqqtnfePye+KWnmieCdONkQpRZhVLnT1n+z2golg+3XzObuv0etC8PInLsi8w87
7d7OoZzuWrFcZ55Q45i0ToUtJyIee95puB9plyUYGa3nBH4v9x80EEWWAYziWSJo
xRLfOab/pquGHhZ2mi8rvgVRyCOyX0Roh0jwR8vdkph5lCsDUTkhmb0w8XMbXywf
LniZTQQcqVRHolkrK47FNrd+azmmsvqL0qWJHfoNIFugWBV+alQxaZHXpS9FlrBv
SXMTJAMoAgUN4T6TQ2nhd/crDd4zB5Bci3fmBXPvxrgba/Yo13Fcif7WOXDJ6ZNt
G+o4Uv4bqXVAvnAX82zGmchzm4kxnaO2JL9l2aGsMcnYjYb0foulJDUGrFsF4xGz
5WA50au3ZyDM5dKed4oprG9YJM/leQ1Z1dyK65UYGsjIhsUC4wY3BLLpeGAI5H8P
qT2UO4gcKIEaHlTCpKkgPO6sND6KObsbaxY97SGX+xdjvuqRZXdga8i3BfWJ2TM3
P4WUUbKCPA6/fej/4UoNwGAyXqFfF6H31jOTzylcyH7mOyiH5FaksmUJOsuEixZN
KGaDblfjEkOj71N/Sei7S8kd82Aqf7VZDiv/2+KWVPngSy6v0GCXVhWDHuZaLkah
EBvfHAeA0BnUrPgjyyBC+G07AB3T2B27TpAWLHX3eVvHEaAwLjiaTvAlnDboSdaE
uatcOc9pCVuXQQxIH/WCiuSxXf8gXk8rZlI6VwufD5Gg4aaoRbo31m4cTJJ8Ifu5
rM4pZDA2X6cTjua3JnBreECwWEqWFxd27YAYm75x+pcxyaPFS6zHAS9RCltWIMlw
CDbSARCMvJpmIKvlRDifi1EtJ9oGPjHDgstnUi7JEQDYINPnwx6s3I6RKirgQkKf
M1g3zgqySve5DUQ4DZdl7JYEm/9/CU3g38cfDfIDdg6TR4+iAxy5uToo6uUSTK+u
giGcFL4k0ZtwOiwqlZ2aIUS4djsoLw5xh1CoY/sOa2VfOfg0tKgDsZfmYC2eBbha
9fQfkyQl4DqyFcinHf6CO157TvCmqKMqjXXw79D8kY5U2tu1OiyuS53gVtx95OpS
w03lD8sXA+DsKG4jJKed5a4Dvhme0bvMZvfn/LK+KeyAZM6K3V8qipfaCUcPPGKv
3iG3O3s6lvSK5sj/004iEyUAerE/KDU03nxTpDwNzTUD3BIHgHmidD0mp7cy/kbs
mlH1dRs5sW3HeC4vvL11Eo/Zj15r2cLaV2536iVzhMEqsq8+qSqiukTCq9pNHKct
1XnbcGIJYnw19+DvZXqXO1AGEOq+ff+3PY2sEsIXjam0/jeN4OkfUBTOCPhvhCYN
5x+aMMu35z8lQcO5trDPm5I1/xERrkTLBN4n+1bgdaZepfT2oaosJqjg3TsQMGss
ThiZxYHiqMt5p/+C2NelB2Rm/PR7qM+nrE6KvGi1dSu48wZ/C4NNOOeyDCnCSE2t
PoXhCiWDsmdFD4JDuZc8tPRdSB3vMMCdERfDE+qxwxFox2+UqoH5r9EQDaeBaKS+
Gtlvn0I5xEYAn7XhwbygSn01LY8xC0+mAGnKvqAAW9Tb3BTEUaZhawqUkX1ivjwt
UmNP0gO646E335odFYJcBJRZZhKVrS18g7RMr+snW91PmgsZQ+RuxEBUWWfLZFe6
Ki7iWZb9twH5B/5dj+dxRHXn6MHVH+5B82Sjt9wigjc46/je+ElgBB1Led3Mtnmc
GO5WIrOPiimAVGlIyF32grGjuIWBkyOZZxNVasfmQHdvCENqWt9A5/UVSYTQigRa
8jodwTWSFGqizYKqGCeuEUQaz96MHS8U0WTIxdvO5sq9/aL9f86CF/GPhHBkvOOC
5TmTBQOHGtPC4wyGtZ2tLO2KfT9pdvtIpbwa1iHOvx9J0ankqJUBxP27EU5vSBJ5
0w4fpZqqlYvlrqRWCZnjO1XWLL3IXrE0DnHW48uIkyTGvM0hAbQIQtUWDnySXf4n
+Y8evj83QzClO7AlJ58Z8PZPiN3HsbB2j1EYR0gUl9nA+31Mnl9Q9W8yDKTj+BpZ
CQvVQhKNS4QjlVB8702XTqfcQjlHyAKLXqs+bNRBnbzrNK9n75VT7GPfzXjUI7kG
Ry01V4uZffCY9hWfBsDEOR1oaerB+xeCg2rrbCGpkgPqDqve/5yeToK34ZJbQCDW
/JnZQBmd1gFCIRq36TuPolBmsFm9NkkknYNQYxsqSbt1L5l4qlZxfl3lOoLTnHGS
RYJ/4YL1xayESA1bPSg7ITgCt/AwVh0hMntjTRAebdVm8nrl5qqburpInCAYU1mE
pouuJ7Pd7I7Su8FvSSbODpug9GX8n2fEhePcyGIvXCAHZg1DfvIU2bGcKWiGDc1u
Ns6QICshxKDl/R5Ims4wE81AMvaLTTtDboGeKmd3MWsk1IFqgm94a1P3VglB4j5s
015710zFuvjbxOugynZvUyUAHSUX/AxWqjrz44CZftEI7AbwYCk7aWPj4Dui9kbY
iesrlTDBVcnETG3MD0iS7qdSm88WeKINpb8mRL1fiZtGC0PLfbC1Dtcr55xDGXxG
bmlG6tT4XsTK5AqvAh3MkcoZhHUwJ9jt1b3mEEh+P0R5JSMjYirbgD9yIJ3ZL8Yh
/eOv/B/CZTXFkiLsi1IFwJgcVqTaG7uZHpMmdqkJWYo=

`pragma protect end_protected
