// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
1kaueJjd2u2UvYMacyvdg+a11hAP9sUucnb0sgCGtoQIvQ/T8scVXXdNc4Y/x7mm+Ls/FM6gO4EC
DkKDj8NUMjlnCTe9ts0uUJbK26QZs0Pvgjz9nVOox/2WU3bR2BNQvqpcVgfmUe68qwqmSsR1ZKtH
6DP9vsOHoYuNNieaeTMmjfks/D8+R0je/eMIyNZB+h+IvQRF+4uX+Ve+aY+pjaGXEuJT2pqIi7R9
50TPPMGy5jjRpiSmNLZ8PxvyUhE9RkMzmimtSIw+XXvmQ2y39xGFb0dkxKo1qDQEcUY+aZhnk1+3
bwE94sDuo/I/XUm4rgBCjSXGVC4vGm7vjW/obQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9536)
LAesEUIqYa5UH84lOGqpl8fwYddKRNng/B3UxsvKMztzIrJNn+0i/BXyXQ61VnIh3/Ja8ekEPCxz
90HWSpwzLiwbwM2bxFNALQ5D1JScHuq/fFGDDn0vayZaryyE/cBW5GgCwE7ZaMMKYnOvtF6Glh47
mscuMrM/AQj1NIaauREoqL1jD2G5QINGSVtMO3qNnfcVO8KXzokHcH2x+f1tyKD11CXW7APO7M3w
BR1BKqu+4Y2xXt5sYz2yktCUs48d23kDoALaGVyQIBhmOJ2fExbzWtr0X2XGINjXPFUWYqRdURvE
QFX8UCVUKc4ygfHZXhtxiYh/rIeWiNEobmP21MzBiWq0W0qzVrzbhIcNm5d7MEfWoWQiQoc29G/o
s/gj+OOTVR5/sdkHtKuhe3eo/aBuuyG/d3rBkU957E38xWkMbprzp1oi4wJmJvJSrTrXb17LVya8
3+ym4Fkg5k7DLRn69JoCQAdq7LwYsRD9cHxU98sNBzDcyO52pNg8kYpXJut01viMWtiR47I03RFK
me0wzjD3cC64AAIt9VUo92mn55MVnyslpayiQ9TYYre4tV9/0vzzBZVbY0AQ0GcRFeF83NtGjWDA
peB7qo+8nav8cNy132SVD1Uip3vmCsXR35+cNV4ih2afwWxVK9RqDp/b0Ekyr55/Pglt9mvYvAA7
Uqz6uAuJ4zzKNcOjxiWrncT9FsbQ5up+v6BqpnmQjeE+KoYNj5PIr6EunR0+a0STv03cH/RLWw9P
qYOZCg1ifKxrXKos2Xljk5UbhJ55VBnJhsYDhkmxx97fCSBpM2ZZea/p4GlW/9Q/z/2lt/jWWlcE
HYhiYKxlnGVC3TTX8nNEG0OkOC0KswB7r48jcWkkbVqAQ0z9P96fX1ba8tUIw9jOIkcZExVC0bbH
EUxQ6r6XgcKyw6y08sGT+/6J/VNfFySsDjQqkLKeXj4R6x2gqr+REPjSb1Wuq0cClNq1E+qBbaFq
/nY5pvclAR3EIMrZqVv9TYxriR/Q1Ec+GT9qwUWrsnqhnHvDGjL8mBp07065VHi79gLOeqzNIcT8
Ava1cX0nnu1U6SKzwmL85hqxd3MRFLniwU5JCn1oSZJo8NRa79selOiftqI46+7absljAOty2oKp
flGpzcRg0T/76epBQ4YlWWStG97X4M0q2Vh5gfR1bg83SWg/jO3Si2Oaba4EaeelTvrVqSBrSbki
CIRL1jP78s48RN0DMis4kfrXi6knSXYkpX23Jc5DAoVid8h9c8EPAyBVYk2LSET/beEZa7JCzg2V
EhbIcAr4RFDteFjf8h5TbHQN/AHfdnwfXqATH4ReUVIef4JX8+oz6e3wzh6aUPn2Yx5cLltF7bgv
ElF7aVAOa5FZJGnW/PrVSCWhyU57mm21AD0j1cBm5eRnxh+pR4HySIygRijdwFl9hY1sS8NH8dKl
xWuobIb6s+3KO/Wsa0WAmK9AEuIA4N5X/JdbTZsEIbDHFs4twhNJv8WP5z7ZY+MDFk05W2JLA3SY
7eiAlmsTXRYq4cmShslw6K/U4ESVktZhKVaI7iVr45us0TLPxrrCHuOyzFpT+SX8xDh1twVPkx6J
scG1Tbo0TJ8duuTFst+HFwkJcmkiXAFlJGipsyMChvfH6rycwCbrRKJVzoGR18zXTsNVBsENsedF
sTK66HifWbvrcwJnPn6cRtRjKXH7pKPbjh4E5GR/zApIJkgQyhU/IAmlBK50tFWyZvcP4MLql6V/
Kql2Yd/+EnkpShq7ovfR+vy+QFqOXwOviRKBa37xs6VAthOBTgiKciOBdecnPHjzdoTq9/cVyH67
BQeKxvJsTEfsNpRk+j5BpwZG2pcMaoFx2rzWDAJXyllXHYksWxtx8mAzYAT5BW7HyPRQjGNb9kwB
a6o85zkGbdzcbIDzIa0dk/jurwJoi51lSVJ2B7rso5WgS9GS5zuqre6Rju2rvTjebazuJ9iR1/RY
tzCo/fADXGUsNPiDxCA4PzYRXe/DTLocOSNgAmA8wgghRD9HL+V44TNVNnZQT+fo2106OH3Q2LVj
1NpfBL8pVysv0OP1xj4e4RUAAP9IAwtG9tK36Y1oQfMnG/rnE3BvWtP7iwDWMmArG/6KU4i/sM9S
Pjcgjgvk7cMeE8Yn+Y/Nb3338BwI4lC9dYufhK0DBiDfgaG2UOYuroD6XC3tYEHkyQzjropq1ALN
sStCM1GhJL/AZipce6WYxQRw4lkaK6Km4WGv/gjn5Kn5nsMbYmDlhpvSJikm8OAZYMN/+g7Lc11T
Rsa6j6IUFmObPciXTIAjAavaaCcOd6InYj3jeVwNbdaF0FWF2SDA7GmCjnNndDFUWZrXt2QL6RMm
OWQ8RKR90E+SrIaz332UnI/6G3iC76O5CukWdiU2em5FrILIr745MYp5Uh0allQ9M7xVnrYoeTDi
4gLV9HQhB9s4C6Qiu8/u3b4XSaaFGqQz+4cBIw1KFjkRHvsgKe2Cby2b2YrGCZERIUKsAJOjvhqe
s8+2dTIW9A2trzIFfFKyN1ZEAG9FIrVS4vv0LNPVc0TO7NmyvHqkark0ONlAzCAylm2pRuxOqpcJ
jqHK4FaABKMxexRFJvazku/6F5hFnCHYng3mE89oGtzYFGd06DwhsQGKu+owzGWur0FnuRpmTxS+
pirw96YJmWiAC1MnpujsRWXEm1aQH/4XP/YMlELdFAPmyG+VPz7glJPPmD7dYUuTNRRZn/b/zJ9y
1Xy9XkU0AF1xhgX9dBd4VgyM72hcgNLFw6Gf+aPNpN4daPGegL3UzhVKumQks4RoTT5ZHNF9BhFE
i3f09W2OlTZeTnHT2jD1jcO8gO6N5hfUnoEtTb7pJChW7WI4G8FlF9QRH9kFWIrQFvIJ+cOOmHXX
hsH/RMWqGdke4sdABASPfO9EA6ZyhkXqvzlIqh+WJm0blS1hpHkJRFIImNpyWUWqcTJrpsxcJAOP
O1oJWIjaAGLCyAe79Qt6DpFQZ9U45JXuBP6PeDiMCx53o/3n7pFRa0zJEVT5u1YOvumWwYmISdmx
/PbXLivyIVMABCppzAVz0QtE+KYNGYXDADAphU/mn+3nwAxGxQycP0Mza+cQXxEUl4FI7lvD/s11
xkzo0g2wadl2aDcy7qtmc8mvxjVXPqtBcfWOMC6LfJ/TsLjRhwpXxub5V8UHwTdS/Nn9K+AccK0o
rn7981BbNUTMK7AMBDHwNeN1tlvVl+L5cQ19vheYejPhU/xm/cJFHuhR7yHwdM0s8autIqx+4JSy
h0am5zJj1Xqhsem+SmjNjWRjspQlfpZHD7nVQ8Op5XxAT4O0/ZB6EonlDrW9iZ97bwFVwceQBq8B
sNv7g5oRYRGt90ffQjvSHVQyI9ls6UJCs5jeRhtkkykSu6mkFoMEARmdmQl6tcfZ50GaxLZdUxHN
582q4wR8c1db3P4n1Wm2v7/bdtY2hzxqPIOO+8G6gg4mmeqmpFBnkySKndeCrvyycOcG+voH1UxL
+SQFIorzAbopAhCh+75Q2VCQE94gE7IumYb7XVEsrRyKGmt3WYVaMBvC4iqJu7AcEoEJ3ne+FslU
/y66jACXXASNJdCRKcKq6wtCf3euYBJS0su3fLpqRD3H34x9b3osAm/TaJk6W1oWKNTK+Iu/eziC
Ekw0rNlJamroBc6t/tkWc4joH6apiGVvKwyW+MS+ZYbOut2rJ5/jNP4OEVdVf07oFcDX7D6tCEDF
Y9ZLn8OU2uucd8pfq/ZI7GKGbGxgNZvdcYdYfE8MIEWA7A17THoMsG11uQAbejJHyZ//7lp79y+q
FhfVtVBGKqC5Ax9Y6Bmhyz7oGzk88ub0C6V4Q6RPd1fFmPelcwFyTgqORbirQh7ScffmBxkOdAga
bUR600S4C/Cms/5apC0DxcNWcQxBVVIjKctSfBOZ4kpGs9TVx3XGeRXb4t5m3+R4wl80A4yxnJMd
X/FSm7g+yED2zQ3BvaGzFum22wpHWUPStvVdbqMkwzQ5Dg3yezoHehkYE824azBIqT2A+6Vi93zQ
ovSQMKcO+bFlPw5wnPPz3jps04wy5MukeLijvBhqSFCE1Ho441LORByQPKxmV0ROIi7Jq7HFunb0
UyrkLxOAao3BwCEPlv6iYUIZu4qveR5Ndbgw4PkjfPpKZKJ5DkI7z4+YIBwhsZiNSE1R9Z7nIev6
hWFwfBhlCYhrD9iT9p0i+jKaQmVGu/NyvIO0Wj6Zp+vkKHVeXyRCDIYM/er1oP2V7NuAjqbpcnm/
6q6CfrqT95xCGVeBWcqB0Q8/XrwapOk6iFiz5CuvpSavjo9TtYfNDPVDd7aCJ9dPsAy68+MsoFeF
ZBq37gV6BGv8GTu5g9txWJMv+PqcXxAhSIWhBEU/oPvfphXMzn38PwWX8bLyHA5n1vgsh6h7GClC
Gux/T5uW+rIiD/XA96StTWlyjZiVbv7NWMuCQENnrAGWlmXgnt92JBvAGLmebDOfIn9IcVeESDKD
lcFjzt/obxkXrzwtd6FQsPXSjSvpXiEWwq2+Ax0xdVxsmxybGTZCl73YEHUZMJh/I3jex9TsG3Xc
57OyQWCFehbv8FCaXgPtdB7I/xPSPe98YAnYu+Z8p+D5rAijxQjrX5Q4I4ZBj7Uqf8CL3cmA1dUJ
6WQIWqB/c/7oav9tg6l6f7Qx/cWI6Ut9rkLQCDfMXXy2MIY18POpkEI2+ZVchTKLdmTXOvAJsvHF
2grOTA9M/Adpl7L5lglmjrZ7RoTVqxm8p8iT8WZ4pSsCcX5z7wOCrqa9B71eCgP3yt36oy70eyo6
VKrXEthBOTEXRbSyZwyODzEw+r9P39wQS/FPD8RVEZ8AIBeFtNdZ8CntcIGWQ8c5NXupIfV5w5aH
6KgYwAHpRNVff1XqCYgeENtEM5gRJSuDu/NUwLRFmjQrdc06wHeu3Sz+lrFOB6LirFYSygvngMF/
ZQzuQHICy8ck+FwyeNilK9FrkSvBIXfOCcMptjRZoJICKgraBUR+9oDHgKd1wDtn+GlAUeRoZFvZ
zIAx8eWDACZ7S2mFIZlbb5e0lqBdgKwhZScRInx4tlqsgjB45N7QytEInPva0gwIOjelT1BmCUfg
ItE0WZthxWKRQeQGqJv4unZ680c9GF7wt52R6YdUu2WWHad+mCYSW+x/p1t5CPBnmac9gWV1RMqP
IguuOzYoT4TCh9E/sJsn7jhz27lsgOAV5PaHOblVC7RHX9ezcfsV3qQDU2iWgJpkhOX/rOhP12Du
mnvc0h5bjscB+7T18miIDCUZjKIB1MCtydPAbJq3NnMlQFYFyoC9kN0ArJ5cufsW/FF5kX8YuLH1
uMzRUSaTisrFQ617xbhlJogIeIXXJ72oYpV6TkVMM1KFuLLmk5FKa6UJR3+KbMOU1XETtpP/gFli
BZ4GMBHNz9vNDzspnsDBWgBngyt2puccdEwawy9GqedPV3dR9hY3RYVrVYAxJ6AGjT5s/UEN83he
C4LDvOwIdi7txE5wxy15KIP9iqWIQX/2mvGFROoRAly0CPbHYBZuYUGaKNjTO7/DcBNCSb0j33A1
RWQQG24NuT5clbKUQ4/IrABe6iaZAT+Jf+T0S0CGxdx7LD6NQKQRuD+ajnPF4qPHFsCGsuTQhQE8
2D0NNGfT7WY+iCYeKE1V28tKj+1kYbPb8GBmyAN8i4/4nVLt66QIb3pQVWmJ2Xlkg3DFnAJUGT5v
joOhhMadi6n3lUt7BCwSxGYf2GpZse7FQzU/3PKV7D04qJzHJv3aahy0tsrx8fG5SP0O8x/YPnv+
Qd0K6//tusIvUW2Er/OlAYW5geAbYuCAoRnRLX0MzpiULlhGn/xhr+TyZzFb0SDFD8rM3r8BW9/h
tGvsvi6wJVhK27jp38iGwtJrXHgXPDmMHEL7BV2r2IFCoDZ6uy2grENNVvDQ55yYqJc0+DCwFLyP
Pyg9yinZrwy5uAlWxGZRKad14Ti0L3PxpFRdxGTjriRwLA+BWHFyru20UB/nDhamuOrZXuSuPoAy
UH3cuaDBIgF9eX9MntbCqN9NOH9PvZPvWWKPEIKYYOZNPmQsYCPPqWbyJsfRk9v2W7wAlBapstMc
1HnpmO95Gu+mHTOd7Td3Qw5DGWwAsfsTyk7z3DuaKy5oYDYMVLhRofDeNoNvmNGmdAB9rBUq3xBk
K+7vShAfiCc/LB2Fph5nvqU7SJVQ2ER1K48Ur0qTolc3bSjwNO5jENDn24SQATzh1g03n3ejz7hN
jXN8uAkXOPclAV+0qky2ot5PLLVmCKk2J+YOCm/L0TI08Ky0RSg2XuIbbDU2sWjJ8ZgXgpCTE7A4
PiUcjLau5mB3Sj6zzJYKH12phtjthf4HwoK38H0VAqVDwgnJ/6EyD3kwQ2ar29wGV1oRGD9Nhmop
HUuaTABF5UQi5MxqxN/O0QitBMn3lwAWp4j3bUt6iQ27ZYMwSXG8dBgsfOT/H0vYUqbFtXdJB2sC
70j/eciqXvlKW/K7LdiRgsdy4J7aHTrLEafMywqDpMC1EcXDukPAXHQ8zI+Yh5CCga8fbD1+wtMT
yhEO5EmvAlwAjNtVdwgcjAQoscv1WX6nwEFiTnMeAc/ASdwnh3WFfJ3FS8oziB+CLzScvQbSHNfK
vX0fXEYmxNYLKpqjJdiA2bZY49Z2aD+6hu/wcFsafAsQ0kqiXwxxlWVvr3Ck5/RQYgSIEjgRKq7v
dOlkkfs6an+BTrF7OFXeAtZspm+ZEcb4sqeFz1CUvdUNGv+so6QKqHByLHKCPH60pX7pByPDXNtQ
Ols5Lq5x540xro3AQm8/m43m5P7Qqgus8O5yFQM/U/RpafijA5rhTS1Ewg3O9yuIiVx7fNrfoe6b
VO1l5Q7Au9JIc3sJWI3ebae2RTGtK8IFefwOtREn8rwh1aPnuUc1ezlyKZdFHcEAesnT1McXOOgh
JFZQAG9t1Tzs+2Q12jRGoJmPD8tKQNrubJKTaB6I2lGzos2AzHlFMi5epGEufyKvtC/ECr1lQjrG
1QH+r0brhfUsJF4wTjIwXWf3jglgOnjnVmiMcP/FREhZBH6Bu+Qewt40rGvDz4g2BXhyMRNzcinG
UiXURlFsaqkpc583Y5N0LumKICoKFJKgLk3s8SaHlmkG7uTiKSjG9TZ48PnIxEjR5sZf6m2FJ4sO
UM9XIzwrDaRceAxFrmTWQQSo+D4jUrTjUuz5ESk+4bp3UtNnY9TqiuVkfxks9HhUIAodURPPoNQF
EY6r/t4tBl/IHW6ZyuvcJ5hEiYxotYCHze/DDTvsuzn06f4+Y9lq/5MS3BspD1i150YL4/AU7nPJ
08R8ktH83NUiFpf7FP5vYr1W1e4CjGcc4q9scKl9LG7bMAeuJvyKKbspbW8tAkwzUTlNpzrf78WB
2fslkpglcEuy07zBNKh+kd2gvcU1yg4ZdapRQC1qoLPwtA5bcbXDOdZslq2IerpuVrbtbA0Yd+G6
ugZrn1EOlk+XOewMbBnyFcKKpMR89Vqes9BiKiglLUXNNny+hdnUBbiZqTrosb03CxHd7gkDy5O9
/yW4XDu2ll+hrK2FELJkGyInWNhZ0kNBZ3QWle4xtw1czGndtH5xycQkM3cjHJq5e6m1mAWJk3yB
32rEwQ7Zjm4XkLAwUPW7mQ30cDKN5cu1HOUUjp/WOZ++UkHaqp4SLa1W8zy+cWVlhK7YzMyt4SPE
TcfyjkS3Azybn3WhzvdNUL4iGrv1Ok3rggDify6d6hbU0TvjT2jk4MQVFUDJt8tvZSAmtjoPj8K0
w9QkEjTvh4DEcpycktcW9T4AakoF2SAOhIc004FUedoBhuIPz4pH9udBRBkveTSkxZ2TsIPsUk5C
UjbL/LvI5ngR4+vVY295vqTqLYShCXHr0aLyuy/usUv9TKpEQVlfFUwev8wNRj16ydP+GuZyd9iA
8wPGM/y3IFP7pJ3FmUHI1V7jJIATbLR2oAtveVbaapdtEY6KWYwzfhR04jKXatpity47fjIMIyAP
doGIEV6Sfu2MYnwBrMNLz6V7h2IC/Zu60njBUfP3jgwsPFbjdqE8Q2VEwOIo1m3sfuZUlfPasede
//nH/WRZWBEuxLLTKgE5bF9ldDbztYJFRbwhWPCLIJ0z4VWLTJ7tAPx1FtZTFajshmodCtHTBQJh
jhPFZ9IwIDc/vUPDu2PX+xWtr4UbH0gp046YQwpLr0DLUQtqsx03kdgb/Q+ydTiS3KR5PCebNDCQ
0zcyRdZAsmp5CisPaQzyyQKMsDEgL60xH/99wLtROh2H+v5CIEm2NgpoCMlBfQYOhxFrDE2wmaii
85lKZxdioFCkQLo/vEOeilnZr1LAw8Eo7b70XGXQGQuk0RWqknLU4h7lCUz7yMRUa1/ekMFOu6pq
uLZ48B5GSL7L/K6Xg3hn7pdUBd7psGQzoZ05BDoxbiszmhLx3O4b8g1y5RuZaugnlhcA4zEAq2/c
VQ/P/VM0+jEMOQdTsrgmUCJJ1Cz8/r5gRZ1elSGHDQYMOvpUA0MRS16Du15kLzF7XJOr17IU/Hh3
LWfpYw5qMwy/8upDWdnd7BJkhuCZaA9pYApK4uZmYlcWziGstan1yD8f/niB017X3WrFjJZMRsEl
vBOLf3lliNj8ffo0jmcGCFMuUD3k45M4WgSGyRgEFUW4m9s9Pl18Fzsnuenr7A0jc7UkavVe8dSu
vA80jD+6KldYdJhxezTjkZvhqSyeo/6Ngu98xuFUvA+5RFWJWWuTBkuv3mulLt0mVvS824ecOP/K
q/F1AN2LhHd85pAsC5ARl8jQa5sqKONyOgLDDuFDZmduPIjlViHNpcOUrcwxcwvsNliGcw0iHMu3
1hKXIViJ1WYlCZyr/E5DpGBojqEv15lBq8N6MrtAqPwmzmOeDi0sLOW35JDam+tpadHu0JoPe0d2
Nvr46DU2QyCOOjDunS/+vitTPzWTGRZ15dpksDs1XQNRphCwrqI30JwN87vEmArQ0H9xg8QKAxyj
B0V99FsKq7nwYQUc2DuW6u90P4iA7WDwo9gDFCQPYQlcBAkwdq+EL7I6MtNdQRBjdIuHD/JuNszw
9dLcULfDCAnUbqQMGee4i4vWwPGy9poC8KN5k2Rk1vyIcm8pYMIjh1JFlFWoOh28sKXbNMpWu4zB
AjSVvGC0vSzdduQzrwm1kpPV/nFVBpeXH6WL1RE/ghuKFTNZbKuSK/li1SfE+TWRQRSq8iK7RGDt
oH+/bbvtqez/4AyVp845Ipbiqiqy80sYBhBiIzZKzQU0DZSQiuGnQTvU88QeS8M1Lvjaeq1mGdEG
/voJD4yiImyELVUAUqJ0FHJGc/e6/sZ3maYMDjvWz7pjfsd/rOVfrtZup6ReUVYtLzvE82PVOLDQ
eoruGu2SGp76MTYI/1JWq08LmbJLn+ndNJwrGXxsaea35gz4KUhsUIOT4nGQwmeG2WOPXgnoh6/Y
pDhXLBbrrnVHXAg6hzAlG0VCeN04q6NU9VdjM+CSQe9H3RSt6coOmMbbISWLehGSkTprbEs4s3uz
AXpEswKl2uPa1BogETmiOFAtLuH3H1jGGipVeuEHn2Pz8bYHd01KazdSjBh52xw//GR7JrStbKOT
Si8//Y2XXaR8lmmzqgL/xi705SPugg9lGWRgYtoUdn1snBOeQsmEfS86YTgsamrBWOnbDaHIRsXy
8M1QKcPaNZKFexn5MVDZbhwM2I53Gh0VAPPyD40ModW+YfaEextZltwBQNrqU/lSU69mI2uqzXXl
IeLYX4IrCzaqlGPDLBZScg+3CKJDSADzb3q6sR+n6SaDZ1yd7Q/y0mhSC1lZ+NZNPwILArOhjjQ9
Et/Ghl+YQxm0t7GCdSpH6g+8XgN3q3ZkRo3idQLf1AMqL5fPMjADVzSuPr4Ling+xqh9n2UO3Ora
Pwb0r5OxSbuP5jrzURooz4/uSC46othgV9SXFVEWAdtTXNcRHmCDHFBAbmoS2nXi1/cVAgTuGn9G
XNW03lMmJi7AtJWwobpmSHCCGtNUPT9dg66zZIv2fRVVE5ThhqWe+Ee4CwbsNRlHIdAa3Y4Zl9CA
7RwsbcsncW55pH1Rq5xKf1eQiY+DtQWwzWCiZSak1kz9Z+seNaXAlUPVjSPg52j9pAO3KO6bIfY2
9RdaOJ7Hm3pGghaMR1tn3FdQZmcVH3YuwKeJQlsZbNX1V5oYHkN03lTi0W9eMuPoGogOBed+0D4W
bzIYKQeL+2ztCxfZyZc6+RIWIBSooOjToQkukCo7Su/FBClhbaJRNovhTGe0T+4W9nFqwB9G9mDJ
marwr1y3xJ5KKxH2DvCROczY300qiQw6Bv+evk9/YnnWqVTh7LXLIePkpGK3axc+y9c7I4NLMcCC
ffh6akidsp5A/7a4uZzNve3s2bi69xnMliRdlYLdk7aZB7aadAQqITu3s6g1tctrV+ZHpZBDEPg/
MY1oKfTkUw+NS5lB7QxgMlDoB9o50oknz9RS1THHPQqLX2/+qWRKMLu8mRjEjHzdJHszxhCksu/z
Xr1XIWZt4BYiavE4ctI2nfni1g4icLl74GKbVUBbWOd0F9s8FR4PhZ2qVrQ2D42Enofo6m5Gj37W
dCHQNSnBhA0fCcqAFagEUL24IbA3EbEMolfHp6MI136KS2biaqyGbCd5HoEx7PhL/8DP7Y7SSXK3
sFP5Rp+m9wmg55rcZy3VwMEB9vcBrO5Gq14kDi7b9oZDtTDhrBQyN4qQyTPW9WEFU/A6HsZktlNm
iBkqlmAAc/YQfPKQnKAV3Q4L93+hvof2cmhFGNTAxj1RSiYCZCu2FZMWMw+M6sJIkSGJo/4KVojj
uW7sX9N+B+36HTiRBPggCci7auDT5N7Xc/4tk82SMZL2YshG8914j+7aANpqNopVNcn7p9DhYTYt
5l/hLJTg+nudhEKisu9J4DxXqU62itgoHKACQgoSiJABVWaTNg4z3LWHkXZjQJOSoEDgNB0GzHfM
5/MrZrkN2rhygaQWu2hKaPgzb36/xVl2iBGIAWBl2gCTEpsTnuqmuf1xfjFff3OX5fouQHkrJIcR
zbpLFBmW+ZJO+/nGtwtsdLAKZDG3jZ4e91dW2WCFYRe0Z7pbX95fmlLR+4Gg28FOpxiX1cbAcw8Z
FGdc/PgX+IjEoddh3ZnBfN91UdGVIO7/9EsHUMkfErOCKMdmwjIRcCyEGmUlVrxgxIHlVGYsopDD
LfahcOqz+kLiAB4xjMvUn5t0kehrpcVPRr/ZlFN9k2+3c71n1eSrN7S97+ybQzb3pMdIMEPYmQaA
9A3padG8mELcoEu6uaq3nI15A0eiVTRxrnp/vUW354sKF9dG5P9Ji8qRsKL7s4rH5qN5D4DKL7tQ
tn8q36yD/lozjgxwbQH0Xn5JjXkVcX4CwIEZchcrTrIMvEJG5gSKOpeY+E5/xUDaNHBOzY9SUCnA
ObTmnQaU/ocRnhgsNBRIEEAuhHrhowH6uPAa9AQBI4YiNXzNtNXPrq9u32x4braLQm21ZDxGw6Zg
dJyftjeMuzoKCEVsIyLPeqAR56EzXJog/b2PnK8FjKu7Q/x+1qis0mrTqoqVUc5+2Cc4yfAB2k1C
FuJKYiltgZZdsBCsv2w92446NtUmj2b10gSDwEGzG0HFRK1MoQgSPS3KDugE0grVhsM8u9YcPCbW
9HmcqIF1T6mkTyre4x+iZymVK2yZ6E23uVNK8yHG9Vodao/Rnyvu+FnUAO640A2MozNtqYIiKM1f
ahTOqjnk4n+m51iOE6jF370KP0Lq+TYDoOc6LG7LLsVgi0DwUZimAVZQA9HHukKsupy4cGc6ImOU
2EYg7M1rG24SoMG2IXutsRXFdsu7RlNqd+2+OytAq5diyt7ZkOMQzRO1N6+R8euVTHRScTiiRDve
Iwp4z4kRw4x6s4f62waq3huaXemR7WbciXd7tRJjmQPKcpOOqJn7NYrTHexrH7KN7SdY0pyheToh
/OpC6+1bVIOVeFMqSogXzsQHxehjjdL2RYf/E35ai/zQNLVHRPwyO2eMv8VCvtaGQewPyOtYsn1v
uwWyciChY4E2ewfLMgqa1dBOudp00MeAUpQqCGfbWMZ6Sp3Cafq/yLQIjU76oPvoFL/cyAFiEKFK
kxdhcljTXFDlAc355a57H6ACzq+eZ0GHobtQ7ZQTcLhxJfqM++PF5phiiXiE+1IouqB6F0rOB6ZC
0eU4B6u2E9Ob8rAPUpaK5EPJhrcbZqpxXPappPjjG57U4X/UZ6/NYOU/oAmLD2SP+mRCEPm8WUKh
S6IKHj2DCTtwGtQ6kn8eGlCd9qRzsyppaizZTWDVwdoZusZlurb8nsgvMxtl9uahn/v55mh7No1P
5Z/0cb8KBnk96+ZqPZRk2ibrS/7am6CnXxy8gx++wcYKpUd2kNLI+nMXOQyUCm8aSNegPkvjShph
qUvi/0FTXJDC1Ee3GUTHeXGDnI1OX4hrWkrbdr30MlGjAeS2mKmIB8Mdlkr/mNjk23LLVhxV/d28
Dhr5I9sO/fIqkT5xzY9nqXatqoaQGFgx05gOZQRBGOQKBLeJWfrjV4xfk4VfkF2l+o1ZY5w1W36S
dfLm7hUMYMpjo8A3w97kpboY/AstRmrm1LBFUnL4w7xOCyBum80ckvPybQDCd7o1PCXUw9o5bL41
tqedcaQK2p90QjQKPj3zHqDf7EMHJSm6t6xmLS7X4C/TM5Q/wEWY+O6U//YjM/CGM2Je4y697T2t
77g2vrGVFWJXKD+vaZldAPY=
`pragma protect end_protected
