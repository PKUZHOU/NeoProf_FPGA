// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
mO0QOJz1/j/mliDHKH6HBcOhZz+Kg5GeKatNLhZJ5DbFKrJNX3/mHrAac/tl88/DjQC+0e5FVSeQ
tUF83GUmqkXwCBafUFTNr3gwBA0n5rWeiKnIVeNTigS0YUqliZ0vzlfA0ouzHUb9foDAKeMpgdRQ
d6KBOBqYqhoYvMLeWLGVzmN8f6XnDBbui2qjA1LwkNiHcEtpFLWOneKo1AJ1L5FAL6v+jyUUjkFe
N+ZkqW0G8gfzV10y4M38rDfDbjyX6k31vdOiw30HOWD7EZnbARHEL3LDYMMnNT33/V0ZQsw8xUMI
8Fl3gAkINjo+NW+Pcn4coEI09e8wGkuS6Oaz9g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7376)
yhPRsIiV9vvfGa0ZvW3bHXcupOzTuXLwncuto71UAfOHW2J77vkLlRO1ltpVU97C5N2PFxiPVsO/
40ta43j+SRZ+TXbu3aAdoQ/Rl1hd+mjg7e+Vsh+pWTj41qupqv6EtFGyeizybChk8K7u/R9j3P+3
cbCS6Bvvdi0Jz2Vw7cG6AbV3RiyEDgBguvoHinIvtKtRApsZ7PwmKdrf2R0+nWakXZ3NFumIQAL5
GOcW6nmLIsmWdBdpP+ifwFWCmG7FUou9+jFOMlH7qqNlRrQ/qTD1xhIWrcK0DAMD0iJptX2CdgrM
ZvRpT5A6ENqbdL63BipTo/a/6gWd922HTScJcaE8bd13QFPZfK5X3OVYUdxHzw0RrMWLGmBuH6mm
/ISUv02NcE7F44HDjRfnTFoYnpRovuNxoLmSHbJvZtKwsZ6+pHWSPbmaYt5qcsmqX5IKLATzMmLI
928D543fruChfmNAj0QBBHXlCG/j0tJJDv872F1IGcwQa3SRWCZP6R5AA5gUi1NfsXpTwvnRiZZ8
vLw8s/rAHC8sZ/YASpd1QuRTBuL+oE9iVN9+1/kwuEhGnmA02I3U/UtFpRVjrXpUtG1LmCme9Ss5
+eMLGPU+0xJLbeI/9pmdm6JKTKMg+4GuoHAVDqE7BbvSYTKxsXIjmY6AMLpxTZlQSanQRA5oA+0C
XFd7Tj8Fmry84dfB6DzqN6PXV6bTtdYRKBx6ItIGu5N0ZfvKWhjvmcbd/RJ6y76O/aT3OfW8A5IR
VxpxAXBBUdx7TiTqQZV2yScJwTNz4CuB6UoKlbPLGoiLS1pNE8PITeKOAQl0bgferOhqCL3eJW0m
bbFcjk5ygU6++2nsBgxB8NJh5YJ62aUbq5VUOCWpxaieIZ+4SiJ4MH3FlqJrrgfRTErEijRNuxmt
HWdimwmrRESOw+L6qodYCblbfm0YakeZ+Cyz3LTFTgGQH0dbEvmxDKrgy8jXQPkP2NsNY0BbxvdH
b06Q41O0tMAs8eQlRgq4iSAXBZcyo1MXNyQSJx+zklQxF5ReZ6JLBvEPZ3qRJ5g+qDEH7BG5V7iO
TZG+coKEOfc/WFnLsQpxI3R70ifhx+h5n1aGdfbsb/pMbLkRMGeaQgnWGwRopKhyrGFnAWG7Wt1D
JGnxKDQkw0Ee2gGNRBCJqDCx/rZbWQztg7cBFxrn2Qse/qvNGA1zFJ2hERAlwl405CL10a2Ww01+
JJ3p56F1qDRtO2QXOGBf2WowjqQZglE1uo8mX1GHFhJAlND3v3okZY2weuOykkTz187fShIlInBY
af1krIO1PgsGWRDNFlSJV/0bDPtR7yLeukErLeUj4FsKY4nevKIVgHGiAs1wGxI3I0M7K51DSaCf
cp3o+8EKm+tqCO32U1JMQyjkS2LLm3h89o720/2mey+Z4bil3/xy4zi/5zXK8IJ3Zj591Lqu7t/S
T4QzIRIqI2R/jxSnO2Xejp2dp1l+jDE9EBMtXoIwEpUgO08jj+NmckV8Mbhd4W387g3Ik4Klcgr0
oA7KoguMNnoBGTUotD0xW5WfpqWF7niEl77UJs2FcA/w5yKngFQtlc3MLWXKn8EKKr737X8BGR3k
bKJFh89lt48/zULOUI8/OKI1GxsyUVALXHF6YVgFlcPhVAHy1KF1YaaUUs2Up4sTGwXALR3Nga/f
jYYfp3d12DTAS627FVkeeUCoESzl7/P4woqT8C/oTvGSz8D4oWsZBI5OokYt5XaBnORIE1AiVoVd
6PYoqzDzZe8dWNmRa6fBtVjRaJlZo1JY+PC7Kn/N1Xwj4smfd5MczK90EbTZ6P1pcYJ6plIXRcXA
V+gD1UBeIQWAJF2h0CX+eBU2zf/07ImSCGlubpGh53AF1BSQatC9FP2WGCG1EBPJJy2XNb42oFUM
GxJNOOH4jBp1xzN6tBkBbN/ZMQFS2u01LNBaMEHRKbguM68WWXDnRIfJmMu18eS4rRjkNAec5XvS
Yv81hM2W8C6d069PgVVVfFvH55ALGDvQjNDx0OrVEFV0iPIG89XGpSFwQMZpTIe47MOmJc8O8Z2C
CfSZKrfZzAfgx2U7/YC6y7E4e6Hp0sdV8ApYOmdy2nr8Kbgy2x5WjUV2aikRCNUjIiPpJTj38DJY
MkZjOBaYoeZwD6nFevbT8gDdghC75HUMuwxz+MK+ys3pvx/fYq4FyoTwTEWdkxmEL/EhewwsaKYs
8yH2w5jbsyDQ75Pj4YFsrV05NAK6AvkAl2PhmkM1Lwi8YM1OdV9Ngi46aFeTMfe53XxBfldDVFze
nFEGCuow5xhC/t9D5tIERZ31SS0+B5ld2Lm2ydcSoBhTnXzBoVMQ44UJu37BCAeas62jirNnm2EZ
ya+wNRgqxnxAEaFB8er3yrYPR5QCJmk5I48eOxkLlf0ZQ8k4LGUTFxVlBhA5zdJlbzG4v6RDVfO7
EvTw5KnFdmIPAgwUMsf9WCtrP046gRmyqferTvafQr3iFjgBwLY9ZARCMQdQ9p2pfSRUWpdqIHxF
IN/EJtIN79Au6cLm+cVOdl735RP3xYZEq9zRT/HMSIF31qRHTwBHrGuTXTg/tpz2jximkKE8yBU5
OYo92hu4erO5vkXrC3f6ZXghThObe4XQG3C+AF4HAFRHDo8ByJucjcF5XoIwQ8BB4k1b5Pai1JYR
qRvpLsEjF8kEJ7oRXGJO9zW7lTUqf+nd6K5UfJXBkcZ+lMWu9AwWEh/jixtcmdQp9XHw9vRPe+4t
rkAhJNYfiNN8KZ0zbFf/6P3Z01zRcrhk6kv8vj4m+tp9g+fqG2xYBYuNkOEENrz50AqyooO+fnPm
LwgRkqIT6m/a8lkwVq/Ze2OWlgI16KxqHAlq/gtd+WBrdHteW6zhBXxWHJvjnCir1xKKamJnXvdH
orAgy2TtkDsfMAzGJ5THFcX7cXCvEaeyAlp41wmrIxtWb65/iaO1rt6zJvmDyJ2zgU2JWWndMdiK
/NmI8wPILxlcOYI4FGGQe22Y7RyebvqBqwXzka78HyMiXZPXwuxzmaYwBCxGLU5TchcIJjxTN/Cm
0yIhtSwY0d9eRqteS2N9ONUHvUmLkGcOMfKcMB9cRTT+Q9M9K4HXgHnLghv9OcN8PYuJSbYSkP2i
yznuyGLPpGW4yZGn+qME/VlosuY5jainGXqIy2XSxm6CDI6Q3gFiGQEr8PBcIz6c54pp1wUUy062
wCT9E/Th5RdYWqspPKVVn80xUSdBQJt+pKB/UBYXr2J7bRBqHsS1NOKXjYzsNqKoQ5QJ40oZ6exK
e16S1A1ukHUT8om3hG83ha0EaZYTudSXUtxzHAoYlm56pd6gGOVhq9HYbQKTyhl7a7lWuShj85ph
kwxoRMHSB3i7MVRTgvFW7mrn7V+ItHJOThPINQRghyw0anc0OMLwtQVSzhhWB4dGNKdH2D0q12Qj
yKyBCKuGJqBxCESTpnPLiMgtU0ylWejAwmO8Zgw3HvFCzB/yAXNMelj0MFD8B/ywhJQ34+rvNohM
tlZ5IMyGuzImO/qbakmkyDPGW22oj22pJ3/23VnOGX1Lp7qVunLSGC1tnNWaJz/BlGfAzT2VMXNt
BnDB3t/IzVthz75C1GNWTl7uBps0tUroCzHeIzBMGveApt62A/tjlTrIBHRpk6Cflr54TZPXVWdg
oUPwq6REopuvp2Ox2ne0lak4f14saOHckUYfdGBWiM0nJWSpuVen9ovZcGv2gDSRzLkLYm+Qub/f
iko11kKT+4Tkd2OsTig8qQMGEFVRHBLoSNrEZRakffkHMQb6dKGoA2LU3LitkwRSWcOFxSTJ979S
E/1SD3K0mMV43IdW4Pm606IVesSfgJ4nVudL8Mql25peXnFw9zLlqLxqGX0WrvBaMDcGi/fzx5dC
rCSijQ0T89Yquv17uU6SZxCXmfHPyEymCxD+q6Vmk5VfDmqJv9s4P624+vK3msSl41vsJVOfCddV
+rqx8N99D9uw49jsEJpO0Tiei4mMRxmHhxjEVrOTpb0M9lhfSur/9yZ76+TwlKYUlKMLTJTBBJIw
FL1Bz1pF1oKEROONZft6Kamd8hWcv2rNxGG7ITZSGNWluTZ8l1cCjnzGGvbbefJvWgxMMBKtPx46
9gkmT2Dqc6gANoaeep3V4vIkekNCh944y0UY3/oOwBJIYvZfxLwzzoIpB8SkM/bgc9J6i/1o28QV
QpgvxmJPqxMDUQJXIJdLwUkRq3QLsl3w6N9pCT0Rk/J8XVVRxK6DgPMtqpHwiNzGsohDrQ1k35iP
X3qH3XqU1kdvJivAvWrr8DPfdF5k9d5KXnL0DvxtME3v2ZhTd6i91Ky+WgycjNP0Kp48cXmFNOXI
4oB1xgHd+kAbSdqSZCNskkK0c1DJQPt7NYYeGdgiHbteUhdGViMiB0FcDk9hTWmAXioS94zZoxs1
WWX6T4V1xNi7Edg8fr02bP3rU2n8Gd/aSVb6z2PjFaGMDuBng+a3upt3udECeZ4u54p/Q+yNlhbE
XEzwVgcrCKku8tHM9B4Zcgrvdr9q7AVdtEumxbcOdIXWLIke1LGYIxx3KEHXsl2vGn66WPVMjGwE
Zvq4sVo/vaZ/z5ThblnMu6YDS2vnOFO4p9BS7g/9f2GVUNOkQeFVZl/mCrSfD11rWLUKrJyrJ8xp
ydJLuN7ZhjaYEBflKQ/Zaxr65/SKpkKkWAd1PIlPo5VVU8UoijvuYMpgjsxFUj1IAj0hxZIiJMGh
AatDUjPkBaotKbJJGMVFis9c2ONMSGnlkjb+92UueF8m3uFJgT2sp6MXlqO09sOsiSp+6kbwEjji
Mvl+P1+feIj2K9if33YoPqtxBeeGxioylejEcEKKWxAMWmS45cYV13bYAnEuUfUQcOvH5ZEFzSWu
ioA37yHk1cMUr/WAlFt7P8/+F4YoUVE2cLVhlLkrbuFzTelwqj4O3DML3GMtt7cgnWNojyo6f8hD
PzsfBpjjhh+W9ixfdhk88OOEeJjD2vHGUiGkkoRUukPJxhMSIHkT0Q14pdZkllpIigAUkiPdexlv
C5vC40wuAGC0cEes/MioH4Yj9PcCkA78rBppw4im+YfJSymUrVAgrARmPczvuw7XalBfAly83xwr
GR9XtCfNrVa8Z6H62EeF1XyK+gaUC7YhpLZEaxd7koirJpsfHWfJWgVHNmJ1FdqjmMETGUtheIPb
zEzaehBE1XvYFAcoAfePClCGvXM5w0lekoifzKa7k56HUmUPQlODL+N4JHiCKfa1cJ9IvTfKiRQn
whVwOBdcSIDHs6qWRUdDzUwzDSEdbprihFEk0WKT/1SPjoqy3l1FzR/z0vRsBcLeek6Htulab6jX
c1yA4aLb7slhEubnILnWG0vHgHno9y22A5r7+mPwP4Q1KqV9WOKkab/MWK4Dge88ATPiF2bvlmUe
fA6YymtqTm4ikQWI+2Qa4MtOWC3LYn/zygHZUJBMj2LUlhYM5GTov59cUOsk8H8Z02WTmWKKRTNT
ZgSe68f7aRsLwgX84aYf2GV4IQEPaEc0cKMNdmx1KDaljALQgc43FSNPVijB2ovH4MPNaIVp41SM
2yKi0J6cK5+ZoBpPv5KowAiaD4qYfvQyl0mIKMj2DrzpsPI2BIXfdyOrpoIsTRDV/j1epjDcEhl+
kIG7Pum/L7sBHsTnVLeqbxP0gkAGjYd0wpFrWei2NislinSXGJcVOt3d+XAUla+acgh3osH3Kq26
6GKf7NSHSF1kHMCX2LxhigqtQszhJvIKRAyDHVgx1K0dsv7QozefAxtP00ta4/Th+HnyPGjReMIy
uTMSEQCZ5IvaaTpOe4GoR1GT1HsqQ469RsmWdl08kT+P/WgYyrlkN+JT/oz4XKaxOzCo2Lbrlc7H
f34r8SLuUTBCRpa/n2FuELhAJQr2m57CUzUNh6PD3INA35gs/IWZ4HxCYuKUFSg0uzqXr4DtgyxK
+VcG46qEvDEeiHAa7M3N/1E9pr7X/mLks0uGMv6ZEZ0d0sB4iwg/kosfxMjxZse7F6TAIL6NMttZ
rOXcF3VBzXCRNdNm8Yfc7AQ5jsVmHPpWSJik1yBBOefltQ4eVatXVePqP1MTy3Da+Qhzq7H7OwF4
S/SZJRy14x8NN17jCictLh5+gaDnMOzY7Jqx6NvAnl151XlekfhnqHsNzH/s5PSaOwtaZFZgVSJa
h3K0MaH2h0TEru7MiZ3uNfkC2/bxBmfYxbiVd/omJ/e+SaExTcV8/6boJjKO+aNOcdVz8MPage5b
biR5f/IJDSo0/taWNuqQrREgZFo67WOJhKIfc28KQzCejhtp3dVMvnKCwrOv/6MaOsE0nJzjVeAx
/CYl+wGFUW/dSYltoR8gxJ/0qE1xPBU7V398TdJ6SW02qgWhY8am6uqXc4rXv/WKhvBWRYEVOdNz
QxPJo1S+b3N4LVEq8Qnfhnso82UDKtgeu8Q2iBFIQZTK1QOfUQ2IPjHNLQ0dJm7JDLtsrXWzgwXm
yMmQ/LQDdtRuZRF63JvKSGC+afu/lZHo+kf0lrH9iAQTcemoXalw1yQHu40/Tosz/k0y9noc3jWl
c03udoXuzkdg5OC6V/UTn+akpe9s6NC1vyqGzlN6ABjY8xxkLeNQvYatC3p9A3BwAMS7DdIMKYvG
DAumYfRJaRvUILnSE4CfrV/ThJ6nvZ13SAzmStjrYybAtRTkci3s0AaLmW92MnKW1TYQDDUDt3kL
g+Ok7hJJX/VMVnsoZdl/ltnCBy/B6E0xqawGuXzlvqKx3C14I2o+6QVCsJyZpx3OmRXp57qKwqy5
C6nxBH9Cj3jXI6jnD9rp08ReFgvXKSB+PU/ZVzidaQryKYWf5ZdbmFXrdE2Ak1VnCN5lStCvjuXP
OB4z+3Is3LoshdGut1ZzSP2Vk23yFDMH7So0jqTcmRL+XjrWMcBsMVQyeXZcceccwqUTnGq/rwfl
C00SgJVO68QVuUWwCx3gZjxfaLwuIP62RNsAZLtMTjaLRG6jx8uBrJfEf/BRsJe9I9DeO25SQNW8
r4MchRJICzZHGbBHXSn0BVmn5KfuUCcoE7Xx2poAtPlkquRxrZQSLPxmShSv/g89zVjsItAzDpuZ
0Vm5SPgmtfbkYi+EhDYYpuFu4IV+6RBa0s/rNh2Jp/kX0WTvCy4H8ZZiLjSq+BtOBOaJqb2nOA6Y
Sp1u27acY8NQFyqhDHKWEEm0WlQDe95qFrizwViEDcl6yFODHgYU0uQzAlbuIvsMENN1h7fc4EKr
GMzsDSoDjsYr32CSHpggo6pf1qJhJa95c5+FAkoCtpB2fYsU5Fye3O+eQlrL4xXNy7MPuYhBn/8h
pSUnK3k54379cNuLurEjTnvyPgUpnUPfCGPbrym/F216vqZH2bzHSpDqITvPPNFP6h35CC62mMtB
vp82bkamsr/X8ezCuiTH5OlOrY9nNmEEDgvLLbX54qd/LwoQuL1YUy9idZ7ltY+jQbeLCYY/Ehji
ruJEoho7rU8Barzz5JGdxBa/gP24IW9Efnad+GrRxeeD9BjFFdnSsLbo/BzbBcVgFmAZtGPKw3F0
XgCkdkA1bzaxQIFg3aMU9+zyuZbIgk1ICCZ2SRphH0JNu3CATHyUvbt0nSxwgQCj4fUp2aVax0rV
T/D+GteE7jddA/SkjevgZZ6r0Xy0RFALZCprEIHcg2E/sxw+V7APX6IzUaIeL7NxzMInmFrnGAul
B5Hm5kdyFwlu3bij90P6rbTnlBm+YKaFWCcggOnrhRJPcL7ZosTXSJy/iO5PNtU43Qk79S4dYlrL
Pu23QGd+J4YbbDXTmJbjpKYUb77NXFvIKppZuXi1Aonn2TMaUwwU6myYDeYpN98GDXRxOJuwbKU/
eb+X/qjz+Kpirzp4lfOSZDZnkM+qxA0vXE+DqJmipmurs06j4TnnAj89ACdqOeG3Hg1N3gZB3kLy
4RqaOxqjJCNcqnkdx1BlLRM/1UUx05/nOi1qAuLUJHjPpQf9O0SkVt8kAdn/3IHZ+lZbyG++9eYB
veOYrRtF+KS3HNOzTn5lM6Hkkt7gBHXCTl0EwN3w8vJXJnGU0QAq2mjFjSuEI3opfnxgxxtYTSWz
YbJoB/yWTh7By5uSMhQk+kUaHuZS9k/cPssTGVqe/ZLfdqCXhxWAUayTcdhyXxkINYtGgAaau6kI
3UXIv1I2d3XPakrgQ1u6ICrbUn5a2r8CvIj6wiaiDWIyJdgT/Yhsp+5ECV45exTL/vWJev9jhRyj
kfCVoSf831i2f8+fi7P/aBs0zvON4mokzQqlzitmHc3+GbW5kpi/s1Vb4XrAQY6X50iEfNtFH31G
JQ4WHhjClNhc5drgNpE3HSQeMaDeMTlo6GcnW1FZLl1+7PPtiGUZHTayLWx6qGenYQB4mFOtIWCt
JCyf6ZO52idAEII9K5clKM6MCuG3sWJYj4UbPfTteKQK8RaHCV9c0bzKPbvzlhaig2XHfDT5LPAw
HHseAvI6APmQZr5oMihGEBrtGXf7VC2CqJBBzU2A7V0oct52jZdOhOK9RBFbITOsWQDiEuQWimTc
DiIJeW/xmeSQ1Tn6N0dRLHZan2kwh1h3C56Kd2lxo74PnJoetJvKOpXoqcwaIgtsm7W4SQR4kYJv
XF+zirKOv2rex87+4efSKo5HW/pJ4JO3+qa3yVkszL6kpPPK5+JvssvGXX72l5o5OEJLQajLYMiE
kDr6FcQsl1W2a5td+pnlLFMSiwBOenDGmnkAowapBJOaM4aLrSSCmRiG1mrvKEfGwPywqhc8pfPJ
Ykn/2K6k3i2KTGLrpbnQVApmzhppIE4slmzMZK7bT56A01KEck6fIZmnP4mESAkOPXM7MM+4eGlJ
JOreRBPTbN9ZR2IaKGLhO+8soWYhemf+cp63pmImjZIXOSnvF1TAjQFoKqXo9j/bTIF9pDf9CqUY
UU7yoZayJZbAQSd99Uz6Mk8TkICCfK/NGNGxjmMPvfoYuJaE+AqEjPt8a5zkUlnLvSy7nAy+jTkQ
VUSkYFhfN5SIGgZAKJbNXUnyJJNeKG9dJrPE5/cLKG5JKX2nXNu6FZV3+fi2yq8Jz3aKQVoo04rY
C3Q8bA5vBopjtb0oUynlcm+BKRpumhpQhW6aGhtauKb/hH70keGJSpmxm3E4SJnOWG83NhBVHQVs
Itj4pJbJkMt5rKz5Y4pWwqLNEhMLl/zz+65YBu+JNIot6lxO11+f+v9UkTbU+hNDoWpdQDzYzPOG
055J+NXwTmXxjRynNMUeT2asGR4+E1Pc7LQKtunyckGtr7tA9WUoIdeujbtG4DFRsOlhp4+226e9
flDdcLy0F0cU/8RPPnCjreL/iTD6sZs/X7NF992YBgneaqLADNbaICbuue9dr3HRFmcx48LT1OwG
bQo0nmQ40bbQoy3Eef9aP+jhI2IttxDPqk4AxFtYRKnMkOFQvFgnlL7gCEajVjLrynz/VrbZyR4a
ee3KiV5+o04PL8UBzOYrspigj/aiJGmb70HxATmzALa7PEeez9CBV+Hut60Mk6pMt8kx5fZk0ty6
ZW2yjUooNIqIj4a6sVEeTZ7lULfyvir+yK2t4RD6VYAMS4CnSJ1FuE0B0SFvWg8pELnhl+36VWZZ
K6TZBrj8kvjX5P86tdYX4kqXhj00TLUGFGOYXxXiyCRnrwjwGsP/8a37DrPqItVB47wSecCj1Jv0
/BYa602ZD44+Lr36WaGLpeAWLD5zmgHgFiZZe83uhV2i9PqFCm8teo0anHKzKqxtCLSSjkO0Y2Xn
4KMCfg9+pYXQSacqaYPvq1SncAOi5PYN3Rp2hiV/VRuO/1N/YU8hVkIgmUjreQqhEwS2LixzNXgR
vNXEky3Orz01InqdNrWq69RYJy5lK80=
`pragma protect end_protected
