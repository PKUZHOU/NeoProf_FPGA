`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
i0UUuIZxXkJUeTcelY98UZ+Imy32z0/czxApx7XUZ6JYBVcNwUH8uVZMmuz0szN+
w159AnbCbZtjsIknbZQgkNDJ0jzIYrpSL8F4xeowNpHw/yS2IFf+MUYI9/zBPzbI
qqQL2dfXh4rz3I1fiMpPTYvH5AlMrrGTzaajvrO0bno=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 7472), data_block
OlmnGIZU3Ae/3o/j8TPVpU/5GBi7LRjJR5vboyXcsarwAZrYM8QOHauomr7vn11M
sQ78/V5vw6SDSkhXuJ1fACTsoQ0zB3YRcBTSv1QdTMIIAteE2vwGY+H16a8zFtx4
fkEP6mcfcBINVhZZ1uqrljIxF/LJq4lFPK8jGjaqkEJZMFEZQL3q6cDJtYGOraRk
e2Eyh40F8CT0A86b2dfE9xvQKUsL7T96Z/WH4COu9AehX/bu+Q2QPqqi21UbB4h0
kIqOumJ8M5anLxhI5mLmTc6TZvUiGH2MP2toIh9Rtsbu0CJIoXmgYWH5z9nuuvQc
9lCXRHsLe6/JYEQRBq+xhQDG1KW4/MedKrrGX3iwq7b61ZOgnNLq07XixM/O5vMO
qrMO0t3eK8jsxfo5fHvcJwByux7a9zR4rjan+FjhNDQNPU0tET4LN2KbRWSLAjgQ
2perQdpUwBu2smRL7isJfQ3sVYG5aEntWjlC/3k1Shb/E2S/zzhyKMLBifal0qkA
2H6vy24tW8w3t5CggC0N9fsCHrWQChAONueIcOL3GdgaZmowy9PCgtNRphuoXAWz
ilUxXrS+VpBJkg4cnas2ZyKukD1bAuXwFJTC+9BLk562Y2AZotlawnhGuK8o+0xX
aWkU1BbiIijL3aaHCJus8PgoAub+5A4bItS/8zt/AiQTqtc9Bc7aOtUVQ8Oqhcgm
x+0H1+OGk8Nm6AFaT4iEUq0ePUus30GrQV9Smk55iuk+ieaJ7ZT/IJDjTLgypc32
34yylsslJjxo2NtB0ncX14E1nKmJOWHAjxst78bcnLxsL7kGQnQqEjn00vMnFqr/
negruyZ09qCAD/0HGShhDuNn66f5uR4YU94XFpUHLH6Y/yjWteWxcYpkMF6ZsPmE
auoLQ5OpzHAx1AmP6QtPoPp8QAqol0PmvxXH6hgeT1aH6BMyUEujzDk6okE36BFC
GVpvO9FLZm/AjIFPa9S6UjaKnrGhuFBmDaryn3kPp5NFfIAkXjoriP4PSfg51t0d
Ybv9wELx7P1Ajd6P9cliPWbqZ0aJMOwcza4I1gkBqMFj7FoPUWbl02mCfDzrtpC9
06S7Y+LCYzPKny17PFmkWCKTVUTDdkzyv3LsWRc6rinKL9s0CWp7cJ4yVcyLZWoa
E906ikEN7St7iYSwvpGQ38lFdm8RUf7VmbsCDZE9hvR53wirSZKkZcGdt5WpreGR
qmyNXNHprWKcAjikoEDjr//3fALQxbz+wvCwV9lVxINriw3NiipHHCgztt3/JHtY
vCcG3FcRFfDMZWeWDk6HKV8jaj0mRgY1QPFN39YcNInPYI9ei7hNT3BagDMvvUpZ
bgmA+baq1jxug7krtaXOniZ21LLXxIPPCNmt/KIVLQ/3TZcONt7DCSZHg1q1CRJq
jrK7L6aHSPze+IjCywmdpMrzeeWZ7A3hif9fLyS99ciCZ7kmHCKWS5tI5IQpLjNC
lfIpF4A/bPA72/5sanKknMrNYHf0WWuh/echy/5XX962vcXPETdVS1ATguJu+The
QSG3ztEnys9od70H/Qj2wgyfTlTWzjxjbgVpPTKgR6q0Rxljw/vZ9H8tzymY43Zr
QRGxEqeZvMmcg+1tMb56CEhiWd9r6IJ7Z1/lpOQmzFyuWkIrkPk2DPZ/bwCytqmC
9hOlX07gu2XT9WwntYVRNBe/a6S2+QG+6OhquuN+osqo/UI4uh4GEE7V2QoSsR4L
bRvEQyN4V2N2vbtIjHvPFs+X+F8bBhAoDdyqQmlIbgubR1ezPPwTz3U9WOiTTP3E
EVoocWlyfFz1oH24+ymYm2FXA7ANYxaa/Ip1JeLCRvhFAF29BwYFdpFYkOay3zdA
uT0xGXofTaM9aG4UT0SMPLg7E0544WxKu04ZkVe1bjqLUBuFr7aj6J4oKjtaRuUe
uamNmwkQXzGb6fMNKh+L75uL141zTb17VwPD8XXMCekQ5QLF0yaqWmdHFW++qmjZ
tzhhsZMDW84ctoIZWWDpvmjhtb5UPfwhkHRa+B182g66+BtS+iNU13VyuYS+udm9
9wIxN8BZVc5sCrn7YxsKCvwvsq/QyBRfJ6/m3BmuVzobg4nGWxhB3ddVRalgH0Dm
awN+vpxZxgW9IyxYXsA1m7xzxhOXXJGeaTJFevJzVRVyZ874SzNBk16xhoBFF2nW
b8Fh3nN0gOexdZ88Uz9nhfCQem0unXBiuV3VjvS1MUt4dAZP2AApv8LmH8GxBwjv
p+JU3V1QYjOjeqsKb8LOhfq7mD7IhTWGfeIfKfa9lZUN+l81PfNrhUGSWMNj1ynO
BgXOugabX298cNtEERTngLAEcT+4zXZXUOXb32klX5Xwdj4HA4n5b4CzMeEks3yl
O/O+N6yHhETz0P+Mxwxo20FVExK2QpdMBMEDAMBBxyI90IZG3rCmoT3KfLCks3zR
flal6s14Lu+dwfsWXaQHH1LDm5nBb9hkLTbHuIu2kTFm2og5znEo0N5Bow8eWtIV
cSfQfQvOAkGLUTC5WNk9uuZnFobiDbpOXvOLGp7ilXS8qlaBUIQ0+G2HQ6S7BB6s
z/l9J3jnreQzgV2evNjO6ENBnksTpyyJwjwfwLUx2an1HF6L9Fy7hyFMbLcdBfqY
AaRq8QycUIz9ebQFEqbMx5n5nH5NdApJgXvZjWzDVaZZbsuxvn92FYb9MRqF/wCB
iQRuL+rCNeTggXE2VbRKmsoKHBmYnf45skivemIwIfGxiiqaEPyHpWYunzoLYoRQ
eUQABPAaBRAomryZHOu2BqtnoiVGSGjIQOfFjnXfBqXA0CdqHUxVn1MHRbmpef2X
N/mUqxtyOmQ4ZV6WZBIcuizfx/Zw0JFV8UDgJ4bU+/KG2rLu0WsjGnwkYEwD2x6I
vwMFt03Iw3MV9UUoax3ZICvDbwzYpwJcEznu8+6mnbkJARr3t+YMocyegKzikfY5
oOl7941nKKyNNJk2XfOi/jCMDx59N+9SLTGe1f/CpYv0eYbktaYb0DMyM3O1qmsm
jLbI78XY/vecERiAKdx71i2CqxQnQOjm/350Rp2wFI4DsiPUnsZuf1gspoRbOEeF
hXsyqYhDY99N1iZMO2FyQcqB88CHHMgIz1jI5XBoM7If8+7t1C04U6y1K7cdQbGo
RwCCvnRi5Y6FsbKeRbvduYRqXvBiI1YJVGvLaz5+XGLsWlnicdKK0kRSJ1kESSAy
QkPeuKaU36q3vR6XC5BGAaZEZs7+8t1q1cDQNKKVPtYjjTjAUqZgrWqenSYwTs68
2RvUd81P6EUrPrJ58IiwPRt1XZn8VX8AjpXbEXR1KO920bbb4VZnvUH0eh9XFtYx
xkBjjHYQcf6pKQIcobfa7G3z3FD1+Z5t3ipkvaPgVSj4n9r0Q5xrjXj4Kj/9ck5z
6VLhujbQPvR9eC2ubHCEOom84t0BAOdKnlHLbn6WXCSqgBr6q4q1Zx/Xd6phVVgn
viO5B5T/9a/4oK19dFRYdZUTEdXhu5rrkS0ILUmP23dsD3K4o6/U1bJYDdHssdyb
SY0aLIVXQzpHBS/W6pauzxvV8kVtpeggXF9f952KIfRrI0HTesVhtQywwp0sabcl
oKgYyTuvXQ1BCDXGVJLjgRrYcCbzva+ivoTlOkSMRXxETlggBylPbL6Xa34H+hDX
Rt6AKUoiCnsLOqzVLxvf/GwjVe4sZhrdQVRZ2fqKLJ+DyR1iH2VuKIIomK7WkHDM
+sc1K1YY9tusH19z3PkCkbPnwnCJXn8x6LSX5bqPC2EYNQ84kfLm2sUnR5tQi0Qt
T07xjJpryJB4apnFOKiFxyftOi0v89petzdkM3eiY6Dqit4BiFbxTuD+ZA+w0xps
CSJNzqqdcaiqsUdRZz+oCSsew8BbffWMpuJtkAmFEMbnUN5/Kg/2OrqpZk5Ot7lR
+HwQjtL0LDrzgHWTPmCi48+mJkLZxdVMxZhWz28MQ3QwDqc1Sixh3tbN75+yv7Hz
BezldiU297DJZGoCfYTOpMeKczK4MeqiqLrWhywNoxcdLgNcFL9dqPH3jXw4t2Fa
g6TC8+ZE5bT+EIbcMK8ki9xWXJdeWLFnXqsQRb5i6PZuwNUh01heMrETKqCsHV7C
oCFaJm3s0XPf4dME+9tfgbielZOxJArH4nMmxzxnAKy028FJfv/ggWY8mSaXoFKN
Humndv/TeapBtPTETOVbCW7XFQYRBPU+/LTxwQNDZVoEGt9ix9kGYXZsn3lBzO5Y
GSlHeet1dTtZce0IQ84u2/eRe+3bY+j1g/+4+6trSW26WoLKpjRcv/WcPebHPGuv
8KfXCK/Za6hDvtUluDkOcY5m/Xy2GacmwlDwR6uaI+NBiu/bHFU6TXfTuhcjEXwH
90sWc0iA0MBNPd2Vjl6aJ7S3/KMzePvx1v0Rv8knzAwHbiPqF7UmYprrC5F62Vo2
hO4NGFsiUp+T3J9Zak0k+v8B1XW+60F313wZkZyegFBLnOzF5zcedQ1HqabeiHB3
5KjpRmUFCRSbfgQTeIps+46aUAk5Ht1M5hpM/eMvKSTikw/YWrMcX2WPge+a/zGG
rOC6FOwiAwFU+/RRk0WOjEldsDw3qJ29Efbre7TUtJTYKpUjtIEi34nOiDJbHZ3l
PYq/5LdDHoRlXJfBUw9MzgntO4x3V3vwVsRRw4COT19EKtAxUALPov7YAtOprSAu
0c+E1YD9T5aB1Axf9Kb35jnsgAtKeI2tA4j/q2fCGykRwqBSUp/cNEenNVxael2w
psP5UPexB6djlviMgoHpMbBq7Kxw105BsiskJdNsBLFX1HREgMn9kp3KvZ/9KtnI
jeiwPheaLXpje0+JP6DmNl+VLXpiNeb++TtyUPPCXhd0P6sqDO9NvAMEgqVwsknU
xXOuxm6Bke8i4WWSXB+yQAKP9ZoEJr7LqxgQ1k/rQvsJJVqB7Ku2ws5U4HxP2Kcd
tAWOBA+oxM8nnolpUIvDhhav6b40sRk3M993EcoAnMA5LdaQ3dTbYZ88sUqNrcfm
RqLm9wTPQUaBMiurNemCglXQX0aLa7uVZdfPNgiXWBnyY4nhNdM4H82TGceDwV2F
9L73V1r6pGQVfZYUlHZDyEYWuS7yjsJ2vKMF530aTnEpF3wQqljJbVs1+nO5ULUO
P72HV0/tP/VUBh74ghv5GIS2Q+6wA8DmCrJ6NyGE+1YqHe+m4Zq900kf4oRSU63X
Oq4/D0ekHnVKtrTbcP0ztSl4MfXmUNu/KmrWemt35Lr6VPzFkhhoeHVULjc5QZhO
AsR3lEJqJ+iLzllny+Fn1D8hF1jdjkFO/wf7oYIRLFbOJb1uisOeGYKZMjNdvsQ/
FKvjp9ES/iNaQ9c1PVV0uS5NR6Lv9A/gm4VmAnlT/oRYP3ll+M2FMnC3xhRnVUDN
LDjfVDejk67Y4qPhToXc2rQ3Wp+JfWIglkv3jn3H/0vV0xCWP1Aofb/pfchzjEWx
yG9IMsYrF5dnkF01uejAl/3zasSSY2SZGqOe3TfiU+zlxUxso23i2Kwk5DFX7bu8
NsYUGKL/rrS8hIsKGNcvODNOWs8Jx5T4NtsnGAjZAESF8WXVOH1/yJxJ3Ru4Pb2s
WDI+dvvIDNGqpCZS+obOi3G64bzI/Ij9t6dn7wHlBlMTcAXvWHbJEB1RvM4jlLTI
uJMZr4B6P/pqF4hqX9qcFrgIShclpLqLhiFQ9ydgrS4L6tpyg21YBXjTDdjHlaYl
8wmfaJwHVge+T3V2802kAYjwbsN2/dcHm2ij1LUxytL2OZ4Fa6YSagm35OF+eijT
SBJcJU0RqnzUgw58PVeyr3p1zbI4yLMMIA7Bh8gaAI7M0OvX1TZdx34mXpA7p5/x
P3xmUYS+OQj4JCJ7rEaNyuy7eCoRJNfjJAowF1JRtzkiAUrfnPQK8ZyE38kQoVSC
0aUpPpqvq/dR5rO6UIdoUjXsSjF9Mjsuokopw/MEEidPX57vU6xerNysJw64mB8H
ZievGsa3fx2ZEHJlyzujQwO1vW/V96tZ2ZU5UZ6O5O8gsSr9WtzHzGO45ayvInj4
XMPRRRCWybNBOLPKZHd7qDIvzQGvnMRLcR8DYedDjhJtvUW5NvV89NbRhDYXH+AI
6XVDjife/2wpvSd/BBj26mlbigcy0+/Ho/ETc8obXIDHN6CoZH1ZYHsieDu84ZY+
U1022Y8ZhlLJJ2wgDfaKYzYYb7rSJh3EMm5uvfFBlvpr+OPHZRygWmCLWh5SrzsE
jAw9CIIvMwWQYOGO4IOYA+wojje7J/XVua4sCjR+IRhw2eAtui4KQi/+pKj2IhsS
St2KFh82+U4iY9fg9K4a7QigkhyEBn6Ozb1G2YraxUaj+02WtuK1sL4z2DbFGr/7
bqvC6QIzNleY4/RTxP0wHKfeT9iA7XD2YWZ5OiFjLNBGiEfD0+YJM7trNqR15zGd
5CZueIOn/ZWTTUF1MgZ1jDXJQT8qJjz1iUekMfY4n2VVMpU5elaf1cAg2naBSPMm
jzfu+EWFWwwWZZdfmkpoO+6xyZXgCOR3qMvZDs6/adDR+m3awKzPJzJT8kQFXV4m
krnxQZqESZlJsYl4rrUJQeCczKF9mddNXsR8bJvsP4f20nuhPJEqpQ/ufcbXSKMX
p1daai9DlJX/ZJmpgAmep+s+GgTYt5BB85thQv3f3U6apyNQPXJy/+qXPpEFvN7d
f6Ez+38fmxcmbur9wmAAJYKQPgpj5obKfXpx9UQHpFp4laG3x1OJaGLh++53rWlg
Xo6mqRjWxeeMXECbkNoLcI9Gm3Imbk7KyibKmoomdEMt/BZsKH9ahxGg/2HHIcox
qb8POk/QNILNuYTYODpYrIqrI1WIMWcBVEa6Ux3KmSUj5lduuTfznzenFDWIsouE
RFlKArOCvTgDSFpdajgMaORNN7Np2X4bn5Ira0vJrB25cutZjs+gcRJjw+xRkQJw
SKWxRf7Y17cQot9NYeResfEP3EauDlvSwRvIoqNvBSXymc/cj1Uut+6hCEuTiUGW
cFMQTUz5mMDTDKEGB6flUH91eUUaBfTDDqCjYJoatcIOt14TUls1oOtjZOjGlVzK
0J0tVcDqEZdSJgYnffar82usuZaEuJmAl1pJwjAavrIXrqpr+Neo7rjVZacUmXC4
H/erqBTx00F+wbkBwDFymUsZzRlDhs8lsIszHe1qpRd15xp4HPEx/TpFlU28OR4J
zqJ/qf7Xv48QD1DVzzH7dzMbT81XAzF3Rzq+4dvta4gr35fi7fnMYPjBzpMt4B2q
VurDPgO1mV2/dv7EWAhvoHaizUeHzLydtsa0LGJSRNwwRCWLEECcZzk8yRxfOB9s
KWoBdFhLuednxKOg8crCzWVOefGNRvlcyuCDNoNS0jjzqmGK9P2Yo4ff03Hr80RL
ccwQFaTOuqeLN5Bx7WHsHKbo6xeHTREt0wEOdHXtIwE0ISY631RN5nKJO1ZcPEKg
f+uivlL6dGSQWZm2/LLybuACVmyZ2CMCrMk992Js5IjfHPB8JlWXMmpEsxv7MBAX
EnmfFXB1fIBqqAWWwVtx0Ixz6cuT6VNXmxsLnPWwJ+udmnyGtYsY/qq4UOhqCaIO
em7QWlXif2vdp989c1ioIAW1BeG2wnTnxJwbibT/USTaGvqk1vfhehzV3huRG9MF
azVsE5BZ+g9FfmFogk3jy/hDNTskxC2YYzn3z2vIpcaH7IWIONMCDaDKR3pn7jHB
Hh0KUssyqWeMTB8J/cLiRYVmw3LwyOJEmKkHpnCX1rPuTNfZt2uu/kofsh1+pdbd
YPWhJKXg0OI6B82+oJTPUasUlmRo4fEHas7Cm+LMrwnzp/41cA+OpuFrbgLhygRx
nuv3TKijUv0DACZH2M9AkR6In+b5IngPzGBtg+CK7WZ0Vm5r0K5dbm0Sr4/hlbcb
ntrlyVOeZAKh8FzK1JyQTwSdlw0TKt2e0SZf0TNWglElnI4d3exFT9AM43Ot/NHu
1YnSDghhjaYlQezdsVEEIW2ViDt4/PCq6T+RTEmSbZi2ZsstolPz9L800aSjl6rv
p1YRT6q9RDIjaa32SVdMoDNRDXPuCqKXiyHkFlRpndnOziOK2xzQK/OHlLhcWCPt
5nkfiiuO6fX9rTkz1u/1M7ZuypQc4e85TmTJFSzz76oNX/OQcjNbRnH9kUAvuZrb
YjhCBVbPByJqS8kC/tTSZKSQN2dQyZ0V8zqV3oEHW5eiHUjyz+jatxuv4OLgshvy
dKVdhZCEnlpvjttLrcGOwYVO1m7P+YmUpAs2Nj7PgrbE3RvGAeyQRbCRWrXlUod3
ShLtppoBcvKS1+wxohGIHeSNo+jfn52mLB1hTqkIzytafnjUW+YdmH22jA8TrqHO
hEebj4oa+Tlne/miVg+nArqrMI+Gb23iT9xk5NBA3DhDeVUqoZJv5L8oYRppvNPA
FHSGT3I+s4rBakTi+LfGNS6v2jper03bLrFZHfqIrw6kPWgGMtaj1T9MDq61n5+o
FbgdvjJnjLUNrw4Y8kgUjHQ0oV32akJD9VuMGc+v5FXMXK3fULVUJ0xpekjZNmre
7hHmUDwkeWzIpVCJ7OnkNC28itKnY2u/hFsa1YY/UwfSbpU0ZthNBraoDAmS7ig/
xGmTwlv4DhJpLIk2WO5EcdL7V3emvvxNwD8DuUjynvOM+WLFu/A6VSSkUUv9DGoO
G0JPktUTojrQ3uuI0tRRexv9d4DHBuUVNmUxsHNOXMp63w1jFwfQMXcqdfW97zeY
L4CzDRweVLIV8bKZcoqiZcNi3PMUOWaam3c95AB3HAOjtz7oqu85Q3P5Ahhd7dba
EDabW/6h2LCCILP4YmHeRRVZJ42R5FutMAcdp2N9BepNy52vCWsllypnLBNO3/r3
DksM1Qw2NsqGs7fsQnYiPuMSU4WCN5OBnPxdd5gpKeakPf0hwZ1+S2E/XadBjQXj
7+Ql+7K8ONrnf+0ltZvaUxW6aqnDFEiBihafYK/pR+nFgajkhcnnD2Hqtpy6xrPj
t8i1g0xERffCu5xKeMEp/PcoyipZKitwHtZzq/36xOfBAZULn/RY6kJIapnYVdsP
ZJJe0vtwoSeXb7qP6Ny3uHURS3VaBy7pJW0xbbQPHJIBSHhUjXcY/9bdS73JEiGa
Ybhq4lFK0Ps/q1FbrMzP74BtdKteapMlE9OmI6TyWOMgkP1BJ/536+ksdTLVk0D9
FA2PWzDIgnRhLkIvhff6mh461INN/jc6a3fcLyyMDfNLmOef/s6GCWdESFSPW5TD
1XhiRJ7D2C+DMHj6oUDyciHt2ilZ4NgRKCpGkgZbUIu4QYG6IEWJ5PyZjaU+qMXR
Bjf5maaPUDVjciQEBZcfhOEkYHSCpoQxkYa2614JrUA5m5YSEXu19zfBPpeuWDGk
9rrGOXhK3wx0W12R/PtqNBx25Zdg+0CvLyqM38ZjAi7Td+J7IklP55z0K2MjC4fR
Ev6Qv8OCEvFZH3v3XNtFY1tA/Ptjc5ILarIvMJg3pS9D6qCVrxIc1/X1cRcNeQdn
rudkmv6HXoOVROVWlEcn40afok6dwMF+1DsDnpu1v8IgKga3B5EBmy1BtLx2S8U5
WqOyWf2Z8NB5Lae/2hSs4g5TOSVFHn0IsDKbxqW7ZlKmUW/Y6ZJ8y2f9OLdZkOUJ
qyV6bRdz0wytwE0rQkdnEIKXcd/EegdDQXZ3DQFGU2bD6HvRkh5V129X+xdNHSXh
8JB57C4wl4hAiVRjQ3FEB8ZjhVxz751esf+FB1lh+Tx3vA6Rm5IuMKqozfHB8PHR
K//3RNlUg9bVFSX6XbpFiOfITUKS0st7TK8JSC6r1YKj8N3ygAEIPRa1giV2zp8b
lsIaCmXti/Pc93dyds4M1W7E3VogQbsgGsV53HqwgxfXKTuU5Icp31N3PZAeb0ZM
wkmk/10Z3tq5owXFse4aT7AbUR5s79T7z+wmyyVFW1xeQfchtIZuAks/Sv2k/Bw+
JbZLtdWaswR8za/Yu04rBO9m6TGAxAh+fA0+TofFTTo=
`pragma protect end_protected
