// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
KEsJ4xvTG1flTUL7Ow/AtOF/NJHJmWj/Dh+NVcOBRxp9oxgpxZVSEzzentivf15t
spoSNM+7V71dCdQSktl9vaXmNaFfoOen7fmg48p5BEfSBz5qamszG31SDja5OAIV
XIOef3ZAhoBcYCIHoLyYeYHqgZ1wsOyioDj5nHr2tzU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 4608 )
`pragma protect data_block
mV92H2QtVkmV2wixTF4KO+FJzSu4iIuOp/c1yAYq+zgWuGFDP6orGPxMRSrdepc3
6u0MTW27fYoDZhJR9XVQvjbUKw0n4ZmzdnmMSOiXDQKlm3/38iTnJ10c4fh1zlLD
AcfLam3oAqOg8EjChj/rolqFOeYAoKJEI17CSdfaEDBNS7nmY5bP9lqVpRcZQ+2R
4UMwE1ZMNOVHoQN6DDvXRBBJmZpW2GSNPH4N7YYc2pbvLhcuXaGrb2z1wcaFBmJb
o/EmGFLO6m/SdgEahKHevEpbsvSaLy8a0Tor+7TuSXO3Rp6B7PhZgSUmRQn26OdP
EHtjBreicfC5Uuk56QGoUmeeC7fgkhfLvkfJmqKJwCU3/EqspLPfIJ6NpiLzE6T3
1EZK3VVRmXZg3LzVSTwxzr3wZmcGUo0oIwMpueAeAnsgGEkYipbi8kg5Ck7fQETV
yszVFskKhX/bqCw00q++do6mAJ8tc4Uw75HTiYXjTbfHL7TXLdynB0vYHlbM6lo4
oVvvX7nZ2e53G2vQJMprYGKnZFQ9pM1c8fOrCRP5KWDSoWf6uDe8t6uM0Qb8zBZx
Zi/7fdcQg6tjdPyc2lLmyOVMq9t5xxMjLxqMNGd2Uf0oWAFkWau9qeJWBty5Bq3b
C1BBOdP2hz6QPJwl1R3rmPvTSFJlBJ8G9Zrnskx5ZGlaSLTTLSzawEbjvOlnWvMM
6TsB41APKHbGmQSZU3lNbO/BLeE7aZzc581laygZqcvI0EGh6emQk15bYKm1Z9oo
8YqFgYRGCe5fFl9+UBL5OrCnyKfKfVPFVjbggGp7Tnf5BFAKLxnDYKmgCAm7lWmh
I7I3Z3SA/gZnKKcUGUs199mcEMxbK1xICm8wPjlqM46rk9qSxjmvCGJoFDegJ0wq
f3R/9r+lhtb/nmVz4rWyn7d858NpwXleV4gjyQreUitK5nglwszmCKnUMe6tUdCh
fBE4Jg8fccf4S76hyCoh9wLU9eijmdMpGO436SZenp8g2obxIEkkftNsM80nbRCK
5ZhZ4iNSYxClOvkBwVVXau859RphD9Cm0qsnNxdh+jycu2DesF6jRgt9EdF8Flhw
0d7eU+Z5Nd6ix0YY3llSgMsStDY4c0wHDjmHSVsj/eEL61zLG1/6ZkOi4nOPoZu3
sLsp9wI1zZpxeKsnH79zUJ2jLln2yjjrlwXyCWA5t4d48eJyq0NLYczJk9IrdBR0
cdpXGNmRdM91AylevAO2pug3LoJTe5ucr0vRfte4XEunSuvDg26kzk9ebf4VaXAe
jr81fyIsE9PzdnsGumxRZbeITEfvYSa8yqfARGpuzfYt6ohzXSDzvVKJkaXkgrXB
eXFkgppZC6w5/XSHZvZi1MCyXGXgQRSUS+jGMTELJz2O/5U3/OvKizOAUXzNX2UN
YhVXl+VrmJWYp69Nd+dZvJyWIi6K2OEIcGle27wWLCrKGQlwmzwkLH2fZxVQScz5
0AS57Y7x+RtiefwYdlPhqlrspLB8IuavSXh30rJlccQoG+i7SZaRzJiupS/YL9aM
pF1Tz8hR5zKyR7DNWWuK9EtgQtmKWLPzduokiJWhjeu04K6QnZbVlLLLGMJRst3t
So/EESPCn0s7wu9EPBpzH2dK+zM6tsqhU4fB5zOEavI3/2gof1w78Yj8BbPBmvCh
1YcyuZ9+ikxbl3ew1W4IWhSVmdpMEAaGfausAYOZPzDIAEkzNbwHXbwHKLsKYA8g
vmpXbwrlxA3q3dXd4RU9+hjQe4HGly8w+mjS9b7PwFbQ3RfHsaS4Jv+2bJeZa6e8
JRuRXu/4QEtB5KVaUxV2Hq0uJrY2yV5x0IDRd+xXM/DCLaXcTy3QZJOsqfLL/oXd
VpwwErfDU70Eb/rR5oVSxtzj/nQw2BRYvgl2SuPMGGsqwAnieU9krvMM4MslOLFs
9pLmZZkE8PE2HoqurtXhhEWhmCU12XYDkarNuI2+6DWxxsyuycKqXAUWytA9MN/G
KXX8OqUdykqKSgqCQvCWZMNOHMb54BeXO59ZEqld3QvUivEcTnMM77Q+FXC2gk/6
CG2ItqdGsuPMNjMT8FybkFsYqOIGQNtkreMvS8NyUFlXN4Wgapj9I3a5RYS4Ktr7
QcbBn6tJoPFOJbWcQZvX0C/g+Ob3aStHB3jHJ09RyyEf6vQSyOOTokUrOwt/qC5j
I5Nwr0TDn+wY4DZ1ScNRtqNPMw3xrDID6jWK/pHwqOmzBUN6rI1OBewwSq0M5xnJ
n5eGi5Mq0GPTAvggXCaSsxWbEA6/Ma5RxskxXK+L4rBX5SyRH4zupxjqAYOc66Wf
pBJbwxFAovfvEbY8ud1YiCC1OSCSaIqxHQt1/hT56cOocDtWTHWwK8EGeACZw9Gd
0F00JU8YnmJY0FEunt8gRpypWMTcIkEmX5Z4RMph0YcBoWzmBD1aL6f7PaEHitBW
w/L41JfvMoJVuSvwyP3iTe80uSRLxbz/F4nsd41ni6GKYcpOqQdUQKVuPk70lyNF
WuvO1JZcjBKrrUpO6KHPLBEIhdCwFaeYIP+2EAsORgKCI9qZwPJ4cWa1tqD3qmkH
FF1NRjr3ocZGsKbqHIT5QsbpB2ZShV/eE47FboH45jAW96Rk87kM32yP3oxCWAt2
Y6fwaeIjZkWJod0BkaWuQ7WpeBNGd5vhe9e3QiBNQjQO3QrIdLpuv75r40a80dc6
PVByzl/n+wZPIsm4Gp5sAS9VHrgkxxJ7JM+Tf3PnAhALTjXsaa7aFXyQr5wtFwfY
WWAd8ZJwxyQi+H1StSibAfBKlDGtlNunDmXTRlIspVRrr1NgN+sbnlB8yt3YVGs7
tRlO8kWdIQprjuT8n+vnR1jaavuGFzQp8LvTH83akpMVekthzLCtUVFImQ8ksZ0K
hVe1SQ/6WQzyF5cMKw50l9/WpR31jHrStWeAq5wxNNz9NTauIoHtV/Wgf3d6UMiL
4PRN+b91OcUzyeckkGBVKwn1JGTUtf+SDsGcNZfmoG0cuqt3vnr60IpleOAxLIpN
6Pv7Z3phIcPpqCiSxN2c8ijPe9JY5Ogx7xEW2mtPCwe/La4salD+IE5QDzFCEM7f
BgtPr5LS8hy0RjB+7u/1lj+i1T3UuwQtvfGhmjtv+GwoFoaUzhCKTz1f9TfaQ3lZ
vWKxuozzNWBrzhf2ZpVquKg6H+x9WFj7bhbqTMLjQL0iEfTPBwjpv54daqyiEeOw
M1QIXW10T/1hcgPD1KZmc5uGvfDRoF+hnm754y2TqsE6RAEUOrskhk9tRx2L+mp+
VFkKYAX6LRnuPD7nALXN3wBmVYVK16yLxBRznmXkUPKj2LqB9K2FepV9rEm9/mWT
+L+Ca06hMoCHXTYauKfeTZ88eqHHOnC2BICWPvhdbfs++ySmQgwpVT5hZ1iWmF1K
K0D0A+hM/mReZyxl+4siaqdznTB2KxiyigBnNowSFuTbnsT7EpQsXt4G8igaeVko
J6rpQ3Vnq35XPdd776kZKBsuoG2ViEzEvpPy7BRXNkyJifPgT/O98iRsSSv0+2WK
J5VISPIO1gKzx34b1sYhptyebICx39IjjLnLhorE0CmJ9yrjG9vvI99mPSaaoQmL
s8G2fLZAUMyDzi59t6srW7Gvv9mig+75fWJ2uzGjDxMbWRhXC4/O1YK/ghUxouOX
+GZkgIa0nWoTYcW3yjm/CmjA9AW6dt8/IGnFOy+AYlSw6qLyGrQmz6BfoOGlBSWf
RyvGrg8cMCEPp5L1kn++X1K9VddXaVO55JXQVTCv+a/N65deCC3GLA8salIE9LhV
PLl5hGZE4odCtFfIu31vWEZLNBZjJrA/rjrJBbeSIkFlfuwuEfLIH0nVYRab3xmP
30DkGFX/3BKK1k6mOJJGXpV0spQ5e1ZLnWm72Cbdv4Jpa7ydveRta9uYuIpEfGt6
7l08zCXzvLDakYs5psz5CNTum1H/X84wss9pX3Da++U1BijZ5VGyLfHtVuSnPH5C
XM74L8qKjDhQjNVT+3FlU7ZWqXoFHw88Gk4Oy6FXXTqKNGYrnmLi62XWfn5d1PBN
iBbOjbuMpZmfTZzguE2Fe3OBIlUldzi2iEg3s+6llyL7WD4PtFhrC+MZmm1vYO2l
ufFd2q7+wQktxc4MLtfiyR/kRKGzNpx480SdNmN/uTdpBPaJDP6n2SqaSYiMH7p9
/xXTDtj15lQK3dniqJRuTEexJctNDeXCBy/PSdE1DFTPJye32APCVivJ5+YymDKW
gURwcejgYo9m20lovVdBMNhy9jgEgcQcsCP5im5qnlqBKKJf2IRHAV9KANJ9Phyk
xa4nOoY6XNVurj9C4KP8XTeF+8xDcPS3mE3yshTORZYDwWQUxJhERkyuPDCJtgze
t1EkZD1kLyb8ZVo30Ueju01koBGbPzFRQj//p5nRpvE/zB0PUPgQ6HArkCShZ/i6
82ZTEaasi0EZOUfAJRpkMLRgPWdQe9QZFR03GE4X0Gm84hfdn5g8INsclSHT4o8f
yrD5FDyg8wqfYZGnxdyyuvCWYxBtHs585WDGsWKMHiQTfi1WL40gkqH/UUiJC+CT
NZOKKT0bQZcmDgqztKkxMwGJi2CJn5+P8n8YPoiVrDFTifMk/ZowuHvFdiSuQhax
B8X6HewnybgUSwnh5X//EvZu1FBH4RgsGzfJ9aufaLWuIRjs/fkqfROxiewblRr/
+33ijcwNwjiRmhGlVpLbErvqy8bNFcJrKLa2YAVj1y73Wq3KaIp65BkmY/OA1lDK
xgDu1YSko4E2sGwt/YV/VFw+VOZ4yffdHARKRHnANoW3lsfnsvLkYaKoDAdeevk6
m7qjGKsR6eNVhR8NsyJHmNJmuh6h9FMQekuPCC+IaaQog4HO+OVvl1QahdnCC536
Tv7j0Cy62mo0JiA/GF8b6wTX6zDZuEQdTLzIU8Lcu/Ac39/Bsi8KRUYTyaJXMPwH
5anpbD0VVANjmXXNJkC6NjL2nwmXgzpm0j2MLXi57Jmgg1O1OT9hxsEMsTUsDPLz
Lxoa/acVC4VkOLB4szoX6U9IfVnjwUQWF/+OJ5Jmk+RwtCZEUPf/7cYqsygfhTui
a03wuZrS1W/9S4Vq+ZninZK+V0NKgs7kFOmxP3h37aNLvwzU5H8NWOaDNhQv1+lq
sWXOBGYDaqnfXw9jJnswDSrkHwNxgraOiVCRpbg/q2DzjOJHXlG0ibAa0WVn1sd7
PqgE0DXFGadM8Rg6Yrx2TOhx3vea81i5XeAamQgQ24el4m3Ps4CL29M7Wd71mtS4
JFKWlAodo04wIeUaDyHudbrwQtNlsDuWHTeocAy4VFbReFZR0QKJNBmyuzRfUvMk
M/C36g52G8oP1DOvfHLj86pPIb/NqYptDU7Xnyzg/IQut4rIscCpdGCJ4nGB4te7
UI5HqtDsKQzBYylz9kGQJsKj3S72xrEOgyecgSoJ0KIpkE9/4sZom3Fq7LC8aWOU
ee+qiK6vHq0mEuKZiSmzwqaPJg9HLpXqu6/YFb8Xc0JYZ15FLAP8X2yd8DrEaNF3
E/lVFM071SnizPFxK5Di4b6xBtacKsiwGHz7vk+ePQ6eIIOI5G7R7eMdX8vNiXkB
jq7jS9ddz2DQoNDhcoTO1GL4w11MIxmNwZbMac/goYjw6jKMyvFXwar9gzWXyUaS
H/mU5uwTVdP2Geh+uImOoECESWqwmc26NyPSAIvDlHFJgryqNJ47QdSKVJrD0bVK
zJsXq0+gIWiBk+LT7IA33JCz855juhmwFBp2En2tAsAzd+uTL5gN1HpVtk/62Imx
DDVUFIcCVkE5XWVGQeR6CVVwqe2n2PXKW0ZK47B/KwVRW1VwiIdBMZ9piXWIdV01
EKfJgApp4cOIT9NOWiIS4CMpK80Ej3lcU210BI4pMxHLPiL57+4ROy1TsMVge7Nm
SXzkpyUiNTF0AYiKgwFggzPuSyPBs5ZedOYU3gaD/T1ZeaybCCyKFJFUW2mZC/Zq
JMBL8TLHhuzeGE1Qs4Az1niKA83vL0L/th97u2sMLGTGbkrw+igLF4vsJQE7hqP0
QtWGj7qS+fHEReEe4DRII62uDLgbBnrZzsCt2RifLBvF0JkseLoXjkLAtjCmgQyT
FMMJMQGU7vsnG+r/PhNzugInDbm7hATxb2i8rRS4uwUyXZ+hZ/9TrDzn7/KvjV6s

`pragma protect end_protected
