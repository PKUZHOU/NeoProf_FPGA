// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XXr+dtXtK2fDXinLG+G/XQ0UmjezWronum3ZebD/4P8wc0oY+bhjtrr60oP5
WKueaIIFli1ng+x+yoGdwfssJgI9dAvAuub5Z6xOyly2DYVhJYg6uhGPg5n5
PF+AlFARpJRLq+Iv8d4Qqnkk88n7OfRHNXc+TVe0hJA9e6Lh7nwKoNgeSNqS
VGCEw9W1U12N+TDvnHHyI2VzKGxk5H2fBhRMlXQZZPzASYzx1UIHCUU5BfHL
Y1IXXuSvuEZLUz2caNHZaUlUXIuI29zAvF4V3bLFqljxiBCrP41ZKRduT0Zo
9ClpPIKgzdwvfFXeSBff1fOtn18PxQjbEDDMl8441w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Qht29MlqDdUXBlyP4TVwCyW5WR+A8o64Me5ScXMgrpF5CUMSfqvUp8M+ts2t
hQ5ilduuU2R5LEUgpY4tjLUjn+AQhkyaOTy/d/Toet+KWucKsQnfqXKr0gB9
Qk4xFU1QyBVtGnQnrbsIotmV/mOczccIM8Rqwj+a/4P7DyFige2CmFXT/Isg
xhYd6Zy5KQVsT8RAyLOJKrkDIU8mT/xLUQfUgF9LMw8r2cI6z3Y/dm5VM4gV
WMi1G6fI/3LxwtmzfX4T+jKVmvHBw94J9AAuoZwsGTNhh78XJehD95o+Wl5U
gxfuJEJd2phK/ePuT/XzSJPiLf+/4rXfjPo/Sn3Gpw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oRoi1LQtQeEamA7tWr6HTEsunhNWdDhYPGtkgbbcfpILa3ded6Ynz+c5irBN
RpO5Lu5z2aGEK/kpx+aFRE2sL7BMvsiawLQabOIactz3kWd6gjOjtZ9VtYSP
GC8NQ37RMPh6WjLCUuC5HbAWRH52uvkDW2Ruzj2q6QslrnvsvUV8sNt/jIYq
lwDM6E+xY3W4Xp7M6w2l3+Tr3IPLYV64velSN0K9xq0c4THaGwT8J3ijEaqq
19XNxRSpcrEtkznOtfXI8oLE/Jcm9fh1VqmO6ggQI6U7/HnZQLcMJhQASC71
1Wqik+jTpPyrV+VkieDcZj1IQTrBrhFe1F+jEJhtRw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MkMYV4XOTo6vKoheN+bm+TqoDgaL4InkJoS9kKzSVm4KRgxVG512EQKIIENj
lPddcZXNlYMSZyk7kWx4QjtwuOjwvspnvkBO5NiFCF6JXThCJ6nSubl9Vw29
Ts8J0humkoK+Ag99C14mXlbDZgATIsn3Dj/U4Xt6auW5L23uW8E=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
G/JlYCKMgUppqVaKJ9t2+TchZaG6N0YZOa8QYzNuwDhD14YvtLhaHnz0NKTs
O6gMwEbrOsqi0A2jtn4w85MXyvRKXbc1N5nPnKBCE7cmqfk3YyQrme5baEEA
SIwDikbMadml0nU2J4uTLNsigvTEEmapB/oYNbB7AivgpUBSM0u+TZdxsn9m
Tvbov30iMykeGZN0UBmL1JJORGe12u9nwZZaExVfEK/QBu9IQagCmwzrOHAP
foc4ZsdcXFxUYxFzS1e8C8bXalC3MjmMy/xNtIh9DXwlgsG1bhIGZ/vpe1df
Lhxo78m8dkibv2vrIrc+Y8VPHoX1HewAF2RzJSWe7hQZ0HuSIU4g1OZdNW6w
A9QMYQ4Brxj/E3ZpYO1fuHq9QC7oUjBDavgCT2v0FDWVyJt301a5mFMgsKbB
6+jLRfTXzXhA+1cEnX+G8JIoFS2/wC0wNlDyX3+MtuGWxCednb8p9CvXqGZW
C1OFllb/CMOpDPJK6kWjkz5UKgaXCPKa


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eK7Lfq4zbPl62bB/CMr7nOVJkPxOmI4THJFPsBwwOUMLIdjOGnhpoyYfU9hH
VrgX7Ixkcm0RJoNVksI/8EeB+SzTyLi3TODOoHyaB9S/+uW4JgByuR5T/d9/
j86GtwnBKLyDfY2vDpODN0r1DOR/GnnmTYuhE4iSRlKVMJlNkug=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uigFUkfMXFlma//fYTn+Pk7Ykf1gB1kEh4QSquSf7fVW714FGAXv//FZJYhH
Na6vcA0RMdGiD4C65YqB5VkslSbtyh4O1Y5aMGVReNItkginO8UB4LmiPMr+
LfFHUXk1uFL9rvoOhhj71CK1Z5X1IUAKlhpHdNY4k7L8jrfX6/U=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2496304)
`pragma protect data_block
DKxKItIz774zAINTuKsWK4SKaSZp+8nrwBUmjKShEeTRpGrO1pF2+oGUMoBz
POATK8Di/kFONlE0JjkpLORmTbavNmOinyPtng70oRnIfouWTHNvxsApeh9S
Fzrah1nfGJm4lD8G4p5XgbqbrX2U7FuvhCSJiyPDy5SRYyrn/BKTEsboV9Ox
zpW2GznmMwRhGfTqQJb6nSNYAsmaZvmn+6rcGmAVCLup/0Uehhl33+Ti+oTW
fjp8+311j60yix1QqHeLTruQq1Gune5QP1egRVCdpbdETb3dvOoXi6EmMJj7
Ihs0Xatw0qLlpmHnvOcyX6Sd9s4XzUypgQERknSFy6O1+L9endweOJT872Qh
H8I4kq2UQJZELLRQ4bWwS5etumc0BUfE3RoY5RzACBcOVqyh3i5RuGRsZCmd
EVLPZLQ0dC9opt5jwXS8jGLesAKY4c1Spng2UIy0T7HL6oqH25CgZ/qSRJFI
WvUg9Zh8gwavOWIRZzS7ijD9cGQ4NOSmS90SpIm1fv35Op9/mpHTTTcskZok
d+zFTySO8RffFjsQ9O/BU8XF+UxEDHB9XhTDoGwYr+wSNkcvO0jrENCV9v7K
ot7Q+pPc3hrVZNvU2PqA5smvqOYisOQydYSNDxLRAnS/G+pl90MiTOwdsCkS
xna1KuzJTprih529F+AkJ/0OZrMa/so4jv153rrqj1p5HvK2f7Bw6792uCtT
zyJP4ME8DTcuG6xfeReMkEsOoyLOYFCZvwGV11jtSvm5BMq4FjxCzett2BIk
mTSV58TTMv1FKH4RZ3WDR22zp46oAKbZ5Ur7bsGV4ldm2a37/hT1HJbfw9/L
fJhcJzXdGAaZ+2OWhUYkkw9/qwuSm/CILlDJUbxgswwkoKCQeOo+6ogJ3tUb
YbSAprg8nZuuwVqQ5fJUQqnxfuR3yLEd0CvJswAtlvHtOdeAui3q9BFNeflM
V8zLAGNGCeddumW7s+17skBr7vNYH4jC9Wb4+ugDAg9cxggtSxxAbGxc4oTj
8VejOBO0779JW5+Fk4mBosz4Vs3Z4+UgWjSLOMhrL92ia5GuSttT15G3JLAx
3WYAPjv+GWt+a9UeGpCRdP8Nbe2bFcmm3g73xJno3p7el0AizGDrBv6GZ83V
78tCyRJ7zWlHkdzXP14pRrs1gSjRKU0oIuq+2jRvp7APjlIaShhZao27ZPXD
8Ti5DXtK6H5iKKzr4rJkBqRbJnxHn+tbpJP9cs4yxyutC+M08NHnU+lqKqYw
pfZC3onvn7MJZr3kVM75AUKzZqxzHO/7cNR/wl2PjCV6UqVE/rHEqPRkg8QV
h+hbgrz7kwUFW8Hej3qSQ5AiKScRW8OQMdGmij5P1t9SXcplACyWKE+6nuUd
b0FF2S+aqF6qUUA5cIiIgqCnwGCL+Egs+dCGgzjxVv5QgseEU0IaptKMOC1Y
1LG6GsJte8bYseeoPWvXzfdkUxD80a0cqlt6MD+O4w8LwxSlC6sG/CpvIUe/
Blv5JSRsgqTuo9oYwYDm7oi3VolXDvSGsW0OElk+RH2G+xE1AxW6lyXUTekM
ts92ekzjFxTx4yOUcmUGdD+qG7TiCUCEB5+hhpGfCPKLb7x8bLGHtXZlYO0J
+TkbCkBRDrY/SlvuxHXeReainy1Htu2B+rPQI4DiHJtAbvdqyY/WT4LADGmD
p1XzDEDhdIjS7Bia3hSoBI+btTR0q9pBqzfd/3IveXUGrra6OlqKiAzwdZ0v
o76pvM8poCVrwaiOHIe8an3XLZ4XHkxIgJZg6fgOuoUtSTJoMaBh2bwBcvbX
tXUhGg7ZK0Q2Ap4T3fa6S+0sphlfLt0n9oKXbRfIhAov6ImSrjozjQfYr3QE
vXxSFkaFQjv5lake776WB6OZOq8PJYwwgIXL9y8JctMQuHiZOt0B0JFNAsoI
NKl3kzHOMh4J3PnIOjVw2QF0C3JF+FlSeBtmZYmeHpCLDci5XWAcQZb7V++I
gpjXsnPbFKaKC3sATNXVHPYbr5b7dWiNxCme3Hax7FYGrpp2djYJFlmzj85W
Oj/UF43NvtqEoR6EofgxdMrAyBr4wR3qocGjF9pUUJcAXm2FVVhCrjxi4lry
Qinl9jMRrN35JkeMzzmvrYS67+e7HXr4wWtZ3XxEpK2Oi2BPNRpYQkROyt5P
/9E2KnXOdKaiHe47DHxG7bF4ZiRkvrd7hoZGs6Pa+nEtQXlWVNdHXcKgLc2c
9UIpho+9dtOtQw8YnRAUdIOK2DC3XPL6yArZqsW/gEAUyXgllbyzGbwhq/AW
+h70AjQ1ndFQ0aMY9dz7ZCug0ITobneNONOOYBnZICrQTZQKBCeEC0YnAboP
DW+GIZDuLY7jmF+Q4/4TuQD92SFLs/5o0josxngQBvSoBz1FwmJFUsDyWFNq
f5Eyl37joYrtXL9gSWDqWLYeG0hgnD7dVMOsnNao+hS0r+QvqYOBdvy5sDcy
voUrGALbXTHoFBTC26eoHygg6t67Oh25HPkoaAmHmf5jk4QOm/7JhjKCHHdT
e2pxnpATCQX7RQCYqPVNx9La7PddS3bfRDjQ7Pr7ABPgGyZ+nMVOKeTAyvEZ
s4MNfXs8JOCVbqdEDZyCgR7z07P8X2luAaeXdlndLoIPOcKJ7LWb/bYj4Brz
U3CuVoWUoQBqq46FGFF/Forzp4aDPkQ0NLAkiT8pQ4rP2AepYXaR3FkDtRZU
piy+sizWT2IHEENikqzE+TwTwCtTsGtUla/XhMaPj9UXWJPWQHvNayw1SI8/
dlJwBRIAxfJnAZnKkZbcc8FjsCQARn70FG1BkeBjzd6OG3FKv3A75EpKVeE1
QTTpmDANMqRssEXGSMnHD45exol/2/RUjdZnGKr+567MUkkOurPzgnVn7p7u
vfZUaXvfKe7VE/F/pWGP29R4aNUP11Qc+wJskX5dWyM811r/RCi5PVKl9vIC
ptIGAOMUuJNgbyPn3xj0qjvVVlrSiK2u16gDequ1Ud6cBLN7byCBMf8Xk4x1
mzG4ZGHKdMHgPv3fmOHdWF79wNmT6hKB2kYMmAsPdgy77p+Ornmg0XUBvDr+
p43jcLOF7kXOspuSNcKShI5kxNMfFQxD7ptC/8qMoZ5rTJ9xYcNSgU3naCHl
SDZBxoMzGag0b3S7TWnc877XMEeTrFaH51zxP3a8qq7cLBenVELnI/1pght/
v5cXxY9ZZ5/kCincBboXf60hqBc/QTXNtCTfHnG0JNZr1rkr8CiEPMzPuJjs
efMV/b9CItryZKLf/yGTzjl2H/8heWvmxujiw1UAgxiVmpOrIiLGihkSXEJ+
9hgWketZpqN6xhT1jFySa2VnPCXHZjwiYQkprumQdZQ/3/IBQj4w0m1R8Tnp
r8dnjCH14w1VHKcnkXBDVQYXbK/eqiWF7Eu3DpVkmeFwmU/6YGP+wDLRxX7k
iCzKCnGQrIggb3VkCW/Zj6IkTFplmb1Ed5ScZXGQSzep5ARcGOk4lZt/s8Pr
AfumKM9+3OmXqw17pQkpk3e4VkdH9Y2nJTnuuH0M/P2+ocEbmk6faMvmnsXH
kJJIviBlZZXWVo9f/e7eduxhajZBd1mcvPeYiSxdAvRWEn8thTX3YQNuGglS
JPVOQYtQNoW8Ira4X3a/Xj+Qguon3iOrQEENmbQXpQuG+tPmFJThy9q8FNp9
dORLXouZiLE38h0/ozYuJeZv8G2N9KClFUCc13QpptEWoViC3XiWEsDDWO3t
QEcq8ATpUMVukSkk31Xaj/qKyjKJia++9dbFq133eaF1YXH5PDHN7ayU5DVz
gGKz9YtYGxalibIPY9c6yeybvpsx0xaXPWees3JYXKoj76xaQQIv9mvgeecb
tJ1GNjUW1q/RfarLXonf2JTF8WRWWh/rtfg/zL3+wyrex31dA02UkYeFGME3
5Fa+EDI9h4+MZ0Llk/PMK9ofZnQumh9D/0eYgYv4cADis7IFUJZuWvdLF+Nf
1oeZXZoH3QWQb+hGXkYIMS7mRLpOzi7GuydZyjKUbv9M9C6/GYr7Jnl+4EZd
+ejkMo217wHE2CLm7V6yThx6YMKQPW/eig0I9b5nRRwKvcGoO/+wvFaRsBvi
wzudrkebaBl7H2KOm/hdln++jFxohF2NKj3jbBd21ab3Onss7wbD7CCz8RKt
7xLVYeST3JEqxUCQpqxZLwp5ZnpRsYotb0AJOeQf6kr1oh963JuQONjvmVa4
daDiRUkFy2q7q1bzzuqx7p0ioTVjEE7SPiNMi6e1nNdljUVMI1SZ+PvzvhGz
tL4Uz/4WgVcm/4Qy+Zkm8V1Xn3jGKtezzTcJR8ZzheYGKrTe/O6VrtSAGSwd
+fGEGtzRsumASAvdOJxOfwhPjusjkTsRsvdRxbboDCt5QkPSuO5wXGHF3pF4
IvX1zzWs4cCzn+39I09K0/uKjoX3Pt7tLbr1pU2z4yglq9JAC/9LeIWZkZrE
fwq+tH5oLOFwumorlq/XcCOal6Z95ZIuF24m6MMtvAfL8JDSzewUt2zmtKFp
sVQZdvrwQ/62iz+fzKQcZsoa99PfK4edJxM2b6NNQUx61bfKma4E+1zoCWd/
LcHBIPgZtaPj+orFjgOjvwDAciqBgfWFowTNlibj8ViC9WlomCKXxZnlOw+a
QBYHipMEDH7VWrjJETjT5GRo5Ws5dOkQn1u6F3CsMwn7uSSBDvzOrDZwVu5A
JT9J+EbmotyE/+fKX/ZJMG+5LpZtVZs4slRrV3nw8HRaRWNmqCtd7TdIdBvc
Thj0lazW05S8pPuOIR6Ab3aLzxOPWo3trkGkEjbdPUxrSDShSlCq3us4O3OO
hMacEj1quvlwlcBXSmGApy2I+Eq+3n/1gJyraYxY9rWRESaJEqw2BPKZ5MMM
wkKWIvVT7afH1Nh5BM+BmqY0u02HJ4kEzunZ1oUDYZ6TS/VUDTlFFwxS5RO8
zgyYfrxWgfo1G6+UhQG9y0iWYsa4oNdl65hznoxSt8/v2FJBMsPdFbZgOAkT
FelK8PsTLy3+QwNFaT/RNr5ehoqtJT0ZQ47DfWyENIJQY5yljwlRmj5hua+K
Csv3A9nvkX1BS8ewkLehAlECoJbkKukRs8IeqtRFJ1XzO60ibwbLvLTcXit2
ldxKz5VfzITFMLBgZc6zZzKqqeVcbN7Hf7Z+EPjBkNR6gtmPV5MZ83QY9XLW
cHTRt0DoV0D1AKc33Ug906n7LI2qKW+BboLahlF91xXat0nXS6FmwyyCC1EQ
iCC7CoCa3v1sZ5FPG6t6mH8ihgnBx53xuwq+20Uz97T//1z7amiFlNRYyuxT
eSZMUbMJh4ks2s8MdQeEZCMUpqvuod9/sph8+QQJxWkRuCsLvn472jKqJzqa
nfWQfxHRjKe4edOt0zngILM9cG++om5hXgjdE70DFO9u5NETbLkd8v5dClOr
qbQiZz+XhZj/uWyUhZrEA24IXShJpPFERDCWkbyUtft7jcsFL+dx4tq3VfeB
BVAoJRdn7aeqTsGyRMDW3lErt3VHQs5DKzJ+24ilcFpX0CCoSHfnvXu5vo2F
sqBRJIWfSA82/ifCjxd2XlquoMK/gk782vB05evCqTF9o3/8hyAO5bh9tZRl
KRWrkUw002PTmjY963FQzqQ0JOOLVkBA1eganBmPUNO9Qd5O/0BB9iFuxkhC
ovN+S7B4XztUdE3/qKR8jyWi88Y6nFv+/Y6OIy/sA5mF/BTilsHIYeEXKJ32
XRkhxQUwr0w3pDP11hmg/j8PtWvTD+m3wl7PkSx1wAIv1dg30Ad9AZgMg734
ypRgqJiukL3oByuwL+C9haV6d9+bsLIKdTtyk43SdrHY+CBwzdOHErAfA40N
h2awDPJTzwinVQzcPDmpCEmg9vVJiQ8OqN4dS6jz8R27Y6ITQHZfZcg+0N0t
Y/ch+xI5tzpozduf6tMjQZ2EsFzKm4eo9qyuMloSVSh35Ay0YbA2SalaebVg
9BH+VrIFN52s0vo3H9fl1RAmc0cgdxh4LHecZsNfVF9E7zEfQugdGCs+eE4S
h0MLpk7otM5iiLp3dPUJ/WlI/5qLLTCqEkIYJXrvBg7G9IjvW5kehDZzCWUi
kOACRs6hEEcnz1r3VKuIgmS2UDA2jCo6oJ/3yGzmKSCa1Mwp+Kzd3USpFGqj
S3MJ7CECRLqAjOi4KzG4JOeHH+M1p3uUyCVztiTpPK9jsp/pi/wpRaxvDF+O
59aElI0QG+XYU3y0uHvyCCzxERpSYZ30XiGci1/9+BN/3Und+IZiWbiJLT72
mN+fYwDXYuewjlrSGy7ILRzcpEriUyzEhWq+v/5VOzqp4amp1xUcSZBFn/24
VXE4D4ucXvSGt+iJg3WW+0leV8fKx3imP9r1x1thgg84h3xjlEdNw/6BJtqa
QfLQ/ZFvtPE4X6JV6iCGqEQZaMgerJWWH3h0v5VbkYxigO7BvN1ui91XeSGi
02IbuqmBG8wNocXMgSylwhVyjCA7Bl3QmNWFCZRNn3T5tYIDgZX2GaINi3lQ
hWljwlVYVMvWnsGuyPmwf11EkWelFyIF+qBtorseDYXhejbJSsqRPk/idm5R
r8ax3nCyJqdkQr0dgS8KeDijWvWVHEvhmydCNdQ4B7Sonyyd1rWPLX+6fGbw
ZCBnWHzHcCghCR1r07k76IROg2EdpAmui+t+HWBiLs3d02zieiCjkIaY1NLG
YI7tV8shBW7O3G2+utrRe7SBUS/MywaB62SittYQOrcQTB9+5Cg3E1TgUFqF
g1T3pYJUopU5/GhNfa9XTbqX60HgzS18Pe/ty/7L5KFsl6I55cjisXWrDueZ
nDFAdEoMqiSGzlPUy6OqgF+TsmiUgdl2nONxYao4qPSGYjioEdp6fEgU35sa
k2s2HW3bVKZGxiqv3N9Il6Bee+t1bM/dxugB+mnNc9vRfaHpJHbicwkqE6JO
GrXpOAK426e0RPeyJ4z9KpuQMLU7JaDG9v3eY1/M07bKp4tP6RwV1dC55QQ2
fdFHJFjm+U1RkJE8J8gr8WXcVbPGrHAZtiNENngo5H5EN37i6J9FDAsqzjV2
A3N582NZGP1c/njcN0NT0V/VMhbJuwznKFuFscTndbn0WXOUmoi4i1Vb4Qqr
apUKFRTrkLytBVHRRm3vH/w6nHPLPwepw+OX+VXgBftgetm1OO98Y7xKnWUj
bPuvKjSEFtImeZibf94s3MMRWT0Ak8RFXqPXO/LSfedNYzuwlXBrMYbUMj11
MUakmyu6qMhv7dm+PdEvLqISTq4UCEjDIjhm0Ob/BGh9agUe+jRQq+PkT3Zt
gBJHVduV2virlvW2ii+7138WwHHejxJzDLpvJ1fDqrxTmmYgu57XnJk34dCa
7J2vCc+hKQZE1D9ku1nUFyjTG+0PVmFR8WIi/QjWAemMGEqGSZ3roXjqckgk
ej5UpA5g7FHbBxMODrayYLxdQETX9gwORhsLJ7pFHIRNYEIylgGcHc76XDsV
7dAZlNUbbgE7gzi2nyYplj77YJXk2HGOwX4nK+fWqgEsee1wE5eRQbhwQv5t
1AQwRs6IXUG75dV13N/fwMSqm2ILu+5DWx7EJ4AVM6ZYqFKOFDcUeB7ZxFl0
1xMdlleOQiV99YNLtpX50Tmswp1zBaPoSQYe6vPUzBsJ1eLYWIQN0XlDdfvd
F+oYKFEN8dwIRs22GOWKu/4kDr6rxL92ZlThiGope9pvc1FO23rRbeRzyrm7
beu+JNE1mq1j0QhDAnXgZ03+sGhy9jSgZpch9VU+7MOuC4EAK/8TweH6tz1N
yF+IGBmrLWUTgw1Cr5KCK0PRywqFNpPBMkxupbOTxY2Vd1D2zawHT15B0Eah
CsCNv+bTCxv38EW33wczR0JUfiypHgCUUYpYGUjkJDGQ7UAG07dFmFe1qf/M
nv3YbO7M/EN70PwDKbsB9w9Ob2RU4kJ+5rPfFI0RghchDbWqI9IqoPzgFOTY
WLFsDaxPu6dvk4SyYCBadjtchaSDjFxryRbmvV1jfOqTGBptlikdRWLbFL5t
tGkfgGjNpzd0/BEgrSMyDJL7JSljofEFiSgOpMye0ll1jZc83HkP2AkXdnQE
vP0I3exN1hPrRVLzZ39gjFniqORzdaPfVMQ10BmWa88hrLXxLXAbK9fWeLgT
dteXrzXAR4yIYYVo5v3qrucr9pVS8N+itmLX8xwrmzhHNpIShAUTRxoBftzc
SV4z4Go14Gz1hCxVmeBii6C3xdkscW3ckdTugEBOrjfMVu5wmnZBYBKNnUOf
oQ06jq0KkrRiqap4PCf7NtDI8R+/Dv95ytH4q4GZrdRa5cO+q+0oXznens3E
XOAb9DpEjTiSGCSsVl7SFqYaDB25Lhv4hCdDR2X7Gxgo2YVH15pU+BCNC37x
bLr32xkKbUpGOahZjPlcxB7BoqToLOFVLNOB6wX7LFEruqkyhMmDwEVf9IG9
vdlpQ2+qQ1swsb63vkticakNqscqWKLgNEwQoIJkX1Ay5YOpjb9u2ECD97XZ
JPKOVemkxeo8Xs9rcdSw/AHKphxPjdKQgrnidTYtvUTdNQotgE8KYspY1LVX
W86uUbWkSc2oNeY0fxzdIU0M//mv3XiTlzPt7AKq6yMeB2vNxZtz9GmOjhgz
snS3ap8oHdTKyVJLnYpBtfmvb8XuqUEVSpN8GAmLtJneXcT93y0pn1VK7sg+
43bez+kFyugauEAZRBhb2XNGReQvPhDP/71HBnnF9yg5mhMaQkge8WVF1uYf
LO79/pDNuiKs21X/QwyqIFqNHNEsZ3alF5FW/aCSX0/RmfPG1IbIpLTj1fqr
oroPG83uiR5wgcv02tMrcmplfSBIp2lqu6ciCmpE2mmkosG4dyH79NEsLcaB
Dskx18mrmga+X/pvO3T3r31FKt5+nbzdSH28N1ei8BPLdxEpdSAhq1+c/A+m
Gogh+4I5jF51TLiZrt00+wMosqD01vKunH7xUtHWE15Tx2gdrL4SbNglYb96
4qWbS1npOrRkICVvohZcbNoTJksIQ6dh+mYs2YJiyppXFIIPx/PG0PiolWke
2JTFITasm1kaOELjaNznnqw1uVZDRQCBGH57KyRk2Hdmc2ulUBSCdrh1GRSJ
wYkOBvGH05s6CPrHx0hslkX5+Ri7z2MjVvlChk0bJ4qALuTDAD1z+FEsbcOk
M3j2VhPX08IfiYklI1ZlxDbNbBxGXEGa9B6n8KoYbGosXyMagnjT8XG+9f2N
cq7dAQ0oARtkA3J/Nlcm+HamTdXENiMtqPdOXrrTWfkFvoLio4mNxyNfJZHu
fpuNV9YvEDkLaooododtvMonkOYa27ZfMtAAJ5ko2Vk2oiGtEHPzr58Ig+di
1nKRU4CS34dY0xOdGqOWMcRftEskl3XLIuGU65PAu56quMMlbt9IP2F4eff5
AunuQQ9jURseDWRK3ZeuVx/9OetQHJ4LCmlyldirMDuFYRwgWhmudSKS1Pcw
VlVCl/NBj6aLw84nlwwwbB204qIZQ+orD6q/+CI9hyoc006mqiCdPlOwv2/f
1kf5meCRBnYBaV4ti4jXhuPURBuT4dvKvZEpGziPU/y36sVmUxYZnpnjACy5
QcdLtGvep+cR4I3TZWcAqBJzHM34w6dPjnsWMNisCT/b9AxiYoMN3x3gBznH
QsiOnI5LAEp1tgXzYyUUA+/Dce+UxEQfh6opf8GX3qdQC0tRT0y39pcGlvhd
V/oj36oslPd1R13mgCMaoaE9MGcrG2QzMPsp3UJ0T1pQSDaJ7eSP2qyz2KdW
U+Xy1ZhRYIqKFb38ppR9P5PB3KMK3QEGfmZodU4+CjUg8tnc7UszqLNQaEWJ
DQPaiv9YYVJZWWWJrlJY2K1A7DUORoTtntitaT/DX0A1ZQRBLhh9oG1ACdp/
HGVgs6LNPgz9Dg3H8lp+vEy4WqdqWEOu2giXS79JnjtNSa9TaY1c2T6erRvq
PkH4vXaZU10KUEMuIFGq4HNKVPX4dJ9EFRwN41yGFvRqtkdD9He+Q3akGAj0
MOOksh0mWZ1tZCzI74+pOOrgtBgtzRojtfSJJBRXkTcnhr/4ExKD0TIr3PSk
lGrCDkL1713VnFPzjmPqs+q0N/JbGMfG6fRk64OBTUaA7HnBxo0lL7r65vGJ
Ycr2h9SQwocivBkfwDFJi+Orouy59QbaKVf+0fe343ddcIBeKT5Un6/Wc8Ek
JbjIfG6ywj8juGuKjBSBc/KvjL3YhDUhF9guZM338JnrWJnCvPNoV7yNjOu6
f7e3dkxZBTDyr3smkYypMUg39kl/Vf0ltv56Fi6zczwprW3xpEXu8geETNjq
Fn3xrHeC2Z7Fi2CA2TCqQYjUC5KnS12rGYVyhj5AOI1Q9ALnlJ/RMgErI8v6
fMiv0uw5TBq7L1eTjHfOi3OUqiZhyUTFoPoqkHjCncAG2FJOHYBSemcAg1DY
Aquqi/j1M+DHfUYzzCRkelDDIeQnRKRlzfCP+fn09vT+4rZcMclrndNCr3Wv
BtRseOnBVdgAO4pIAEqLQJ+iLDT0LG5bCPl2YAEjwjr88JOnmWpPIvC9KDnR
iQpCksr8nTZW5E2STt7LkdKd89gme0qjActOyq8ziHK6FLP78GiBsR0zoy9m
NnW7NPAp0SLK88kAiS25QLc0zSEqihq/kxs4U2mqxo5PZcsNGGmgXlBHw6MB
POJgJrk9ZyvATtoz0RV+22To6kUgxNSTgd/KYCSWj2iIJ79Ej1DQGMLQM24L
iJjWz4Ab66FtV7KSUevcstKqIE2dc6Hs/Bij1dPW4sIT1UPmhwT/63LB91BO
+wLkw0ZyVIE6BDmIEmlM2RNBV6+PCBdo+EePdeDWog1vg8gZUfdVrAILE8Kc
CYS5IkuGwHcx+B6IZsdpOdOpFjNKQaOIZDoSgBlbXHTfJ7qPQPYiJb0fyaDI
Xn9idRvF1F8sEUAfnicBjvunMsRkNP1BfYy71GK8kd/89gYWSfNHgKsJrGIg
LMAnK9xiRU7wOYWWAUv1qXddgrNW51DSGsH3B5DPV0vb0P/4iP7h0dDtuOcr
XEtwQEhuWp7KXSOg4FYSdhmQsG5tK2kkvN4QUb+GdaQnficcdbDhF9T4D7Sj
RZlFlT7THJ+Sub14D/iWzhRb2Qa0sH2g9kS6AlSLJgvCG9fFNoM6uVlbgIfT
E11j14yVL4/8OMe7y9Dn1QCSFzZjrDiPhkEoRFKrmL/Us7oRzTW7rR1YTUSv
oFrXZTJe9XKcYMVDDNK6iqLi8GXkXkNzcgELReqbF/En+rWjisDuq+MiEraZ
ycV5DeLgqfDPtDbAJD8mhXwPr2ld3kx0dN3RishNxquBLy3Ola63X+/zQNl8
C5Pjup+LwH1FqDG7vRPgSbiFUNg51wNoBvZC4+86/JRCe4A5eUXmSmjRWM/9
fnNSahPbQrEqgSiGqAWci/yAZ0ui+k80ZKn+BpufJGn+IgI8XcgshLebKuh/
B2YVosw5xdezA3eEZnHSHU9QnRTu22DV7aPB8afuGZhmUpoClpUmTtjoJpI1
G304Ao55XaZovW5PfufhkyWAzUuVKoH5DFf/vhK0OHSRMedUFmqTdidG+qfv
obQ9yFCa+uNzLmg1iC/PnIMYTnJBUtR8cJUa+5GSx1I0if+RyfhikPVrd+Eb
utx6rPTA5m58lZWNWaP5WkbqZUWCpz93/Eco4RK7A3qaOAW7kw4gHktz7NPO
Zngi3zLqViDY1pNC5J66BlR0iZwXuJkb3y+l+OVA9WcTcEGKUZe0t+58727t
tiEgLZxT31hosRy2i23gE2YIqMj8sL17qJG9MumcCEKMzs5u1MDgPyCB7La4
ixsly6s5KA3bkmrxckx6VCj6Df4hGedGBdkbk80nmhRsM5S7ZACoF2+XHtdN
ymnGOhJSQrnsQ+Hn5x265MDcSLcVkz2he/N2QNmPhEJVd/qqXifHzg/ndJzL
A2OGPi6WNAI/NO1OK46QIaqV2K9P9R/Bqi/BWhFxaVp494JlPT8SlwlHD3/S
jz7Z2f3ac81S8BqF0n7DNy2pY6wrU2NBLeUDrym05F1CGcMS2YGJPN9jawIk
1FwaAz5Q8nmTF2tYI/UReq1EX3f758S2FAc3IILFRPvRlRO7tr2PYlOiZnIN
mMA4qnie3EwDLfKNFDBzWs9a4ORX6x2WSRzp5MM5aLvVmgsD8QED35iUl6c9
MNy7SMqSIobxDw9k2Y4zSoS/vpqzNiIF78eaXRprhe/hc6/0h6fk2BIc+x/q
6HOhRkhcLn1uEYyBCc6BTQndtXIy3OazX7FTvZQ1i+fFHcascLK4Lr/NOdIr
9U03/XFSwW7Q2huixP4XTwVJtcHdX5rnyaZkyAJR8VJHqFKYSizADQrcNIxv
GYc8/Lmi6oZSLcagzyCgkKsKtcPACJ1U3u0Q6wmSZ8b8ie7sKCxOixVknkTj
VhMiJIQ8DVKQHPESMBPtJP6PrVZ2sEBKwwFKGRZu/jomuCVGpBjCF6VR7uZ6
uZIv9Tx+8wc9dOB8Htnta5/Y2Su2VTcmw+bHxSQ+nnVabZFnvFBieyqEKqzi
gGNQedQE9sb+P205QTKmRR/WhgJrvdl6DmQUv094FEhCc3eFrKcEp8kncVMM
Q+kShjMb9b3WFchf6q91IofCH86MPvHdQX+j/xesR0FwacVCThP3Q6TTonL8
OpLF3pll+gaNZmmtPb3xdNCBRHGKwDONMxlfmtNTcNpos7q7sJLRKCKjxxdC
FGIQmQ3r4vjSTY4+mUSEMq/EKEN0tiLhNjvHG0zPuCyG/6qCvzIkDHFEC8bv
se1m55NkzPlr8ZkWA5y5f8MF6NqNet8YF+qDT7fDLiQXrp1mBOglng25R2nx
vLQvwb1DYMisfEmRsN067zNJvneet51/ceOXzkfkhKMhLvDIab+uiuOhjpFT
E3cdk8PRBValqXx/Yi/Md52+N91EjMvxSFlvFe+8TXyMfNyy0+iLrLzt9SaZ
+pfS7BriCulb00hL7yS/LhNuXY70GwfmFeiqVc4ECjOONq1RO11rtYbtEx+/
i0z6mFYZ08TOQl1SCPmvHptJJ4zxaK3E1ysnnJLv+UE+1eTnN7on2RT9Nej3
zHG26OvnrGxW/Vi4zmYozPfaOnUDobawdBjTyoLNVHdqjaJYrWb/UQHfrR3O
cmOFNCZjeMVyxQtR2ZAaW1FhQlpm7Bio4/3Io7e0SIl8/2LuRFhDvjnQD3SY
95p2fYOd0QAdjzx2BKXf2BsEZHltoAEfAxnRf8Ao19nWRJ5e98OR3vKvOeR6
vPKJKRJdGuasxaIUi4Yu+XFrYZR3HJKPd4QB2HMzOc5hcnkcFzoXTnzb8E1f
ixpyfN3yCL7TdXguIUMS5wj5UPf/mmluVf+XE50/caRnaBBr5P0BpQKCIjJf
S1lpEAfsw8z35fY5ENZZ/oIkRVMDvwZ4DkdOr+eMxSV8w+sqaHqOGY9qD4U/
ja5Oa1xgqsGcToWa4KwORYDqO1gxI85nXckHIiTPLlbGT6/svwI1QbryKE9a
HeLJIM5HdKBM1p37nSwzNAl2KCpr3QwJ5UZdnOTgEvnvA/MvNuMznK3vDUu+
Tvre3MyBKg5NP5VO7y+OIFtNW94tpNkG4vgw8N0rN7BurZoc3SYJwHdOI9qS
3UrG6BByUwDQiTGi84LvZB6ciDftzxNHwd620PlSmLCYZaqos9hpxeoaCRxf
Agm+YUocn3vNjRlCPvwqANUqBdpLQaWBPVF/gG4oTqO0OEGJ2j9bRpNZOx8h
RpfMYarYThdpcGMcLc9qPj1hkb2Ij9cuywQIwtyTQnpkJjuOIejVZv5mPcIg
IME+OxBc/681SE8yq8m/ICh9VweYiSOqJWjCl1LMCBWDJwjY1F2gU6CdbdjL
iP2MCB09MZ9qwl41C1OSKyUYIoeZEmnqoS0goF98OG170m66rFMjZRUoxsyn
OqhuyCM9nhwInsNUu6Mx0575RkMvspcvTRgZ+EByzdt91ussA0F6Ib4VXQD+
MECY4ffciBejSh2MfTb4yge8ta1L/trJpIoTnlVlOaHIm9QoaNHVNEsIZcRS
qYdTflX8J5yDow6Kt7rGsD79P37ucU0qeFmnGi+7WTU3rY0IpixiIfuailWU
ojqwqSdbpaTK6W0KyXa1D8CyRaRcpyu7NYmeKJraDBJJSoPHLU4OhvsyOV4W
pSQyzdagtERtfkK18XNR+OhY/KMN9km5fvxNklYG39PVYiBLYbLdlY9IxMbl
SHpO5Ugthee0eRDwpG7Weo5KQ9nq+bgbl6UlZjq5Ae433AlCpnn39J0mdsCU
nrbCNQWan6gAXInXMkm+vClZk2W+zi4Pdbdn1Lk+SzN+PO1pVpLZ6g7tfPB6
uNsFGnoqngeewiAcmM3teEs2GzDyHOuk1iz/pcsKcdHwvDFiRdwOlHu6EuL+
H7e6YRFambP/U/Zu+JECYdH5u9mAUzEMMWeyD0wOsJO5/cTeOTEbXzpxySPd
BgBOYnzFlNvqYFTcLd/xuBc6bFDkNFII2ui4sYkfEM2roqWAQKqJHi+cgspV
6HVGvNjHe4qGVHNAA2Ib0YAr/Wzr94lZYeuMXa3UWj66sCWZYXzBgBJzD6Iw
JwUEvG/A7rN8MBuYzArx3XFhXwgZnIZgbzcQ58l7o+cXTueNKIvRpidmD/RR
T24wwbOz+hWCB3mUhhfMivg57jIPwOyxL1S0qzlYSJ6vcQIZF8jaMAVg9fJj
PwUkgS0hscn/CkmPl/lXrntq5vtIDekHZcQdguvoynu0/2/3L376WeZDCmpz
DXITgpL72URufzeXjd7DfJsfmL1PKGcbi6rkvSxbviMbp3JM6qUKhQFCsVmc
Vn6DtW8uxPNWtQit/ftEC8yjvXsUetVdn94WdYEhOz2BWzEZDWsh6OzxOZUC
rq+2cEejL31sdZzdppMLGTy8dnDAkxPwdc5fgLQwHlxUP+JdwSTitxT0iOm5
nlsscD3lGUIFv8z/J7h+eys6vXzXynr40cS305DlQwTSGSJBXO0x1Y6C6UJ7
8K/z+K5yFPsZLAsxpYv+yBn8ZfXRsGn41mu8xQBYuEVEAWZ4rinffZq/wMhV
Se3PWw3ANprxl5bzO/qESmm3EC5YyU++c98LkUQBlQNdU9tXmbPaFCp/XS8Y
dxcwijSVsJvHIyrHyJSLdIPNJ1ugxLBxU7ENNqsnTJM8h4JLoEMc13oY6wm2
c+IMoC2Uu/SRdAsbTQDFsJupXk8nTAe74UmEUrv/DlOM+yiJRtK4VZr1J8By
6vMoXiyDs8NPKOI6kjFdpPdzgihT2ncAIR3Nz9OCHznybyd4qZSAghReogXL
YS59SuGK1VX/hcbtLcSbmmhfKHTxqDkfVg35T4N0ridxktY4DmE2Xk1OaVYK
cZ8Ls+hI6OS4HMxKM/0i+Ji5myMQmpr1cAoq+yH+o5qy0OVp6w6dBMJPt7h6
pEpA8Z9hbz5Rkcx43z+53020mANlLWt5rJQd9i/jXLEtZoUDF1AvWA+BpWz0
32lAGGA95VqBw+7/mxoHAim4oTx2yp2pf4qeegnE2CsIwXPaZhyg9746HgqH
V/KGU9ckWhZnycV69S6gEF9UOe78dNGzDNjVD7e42+6IZEQcwD36Exx6+0Ci
mUQD1M7LWlYeBGFRJztkRl/FBgmvWXKuJpAxY6uZEBYhIWX5OfCz/ladpLz9
KKnJG3x6jytmAkMYZuRFfzD5uF3Lg+/An0AtiK/asa7W3vnrvujjLLDvnN+m
yySWdjgAM8hv5Qu0itFbkEFjthBNHIg8txOZHI40wAsmgSWSZ/LSjA775vMb
2DslsNWvmPnL85X6JPZiHGXNPZi2hvwXJ7axxxeLHcQj0SI/2aP0EPNnqD1Z
hlkVlnA37lnU9Z5PytAlXfc8ICwXcKnOiVFHWImSUB+kN6YZGKv6JCis4o00
gPLqGij7Bi5J/6rr6rkNMTUkomaVwanf0ilNUof9sexLS3WTVSuXYHhxn5EJ
9MOgRwvSM3QWuh4zzLcnNUXAvRbBiJp/3cOGYLTlYuLa3TPWm68nJuZ5TS1p
00Wm6rBJVytLnuUUfDqGqSas+i5EFaoUb6i8WSxvW6Kode0TvuxUBYfzoNZF
BVQNfKOuVuCqTassrV6tQ9qDzzV4EPE09rtVYTwyBATpzKI+LbJheC885yaT
lQxrzYml42ag+VMP6Fpv6KO+IiayYKSOAH5fs6w2u+7dXwVANoA9PhPzqCka
8lQMUW9SPMKT0wQF6Z/McoPa/NkfsUf2vwQLSv6bv8aTpP5YtsEOwPNEFZtH
e/7iF8hc50v6x3KQ6Gqms7Vn/0RB+fBFbRszpGu8SDBzRl7hplgYP2slQzB5
gh1OFaCT79AziOHAyJFmqBk8j/5oiVFl/Bl4+PoUOMA9PSoGOPFaDzdLlsJQ
uLSLuCnc860Kyyu9CQic4Krr7U3svd3HlRPtBScZxO3liWTWkpSzJWvdMRVS
3JkHutoA2oM7qbFCo8c3iNQcYhHs6pR5Nfo2lha+ZsU/yrX1fkZ+CHMNQUcH
NBJ7Wjh6OSFd/aXehBvk8rMl/8OObK1nFUSXLAJ3QuqseF6GbOuoZIFq1xEl
yNvZ9hFHCdjNZG1gn2BEc1X/rIh4xsMIhOaYHa/wAtEb+rYrXcf0OxfQYqAC
xd2Co6RVcja/XqNY26FbZprxVkZqJs6viCEAJkLJOBX7JxvpD+QwfjhDNywr
QH/RCgXQgbMHSv67qFoTJvPNRPKJMG3UbTOd3bO4O+iQFNzDBCDTkv29I5An
ttr/B3Hn+E4c8mcp3Ap14AtEvMw6za6TSoOkNjDq0pezAJJ/fDBZKAL4fLL0
AE8SVXdled9kAhHXhz/Sl5lrAjKMEt/hxDDCH95ZzoDrOGrLKwpp1nuZ5d6M
oVXT7UgDHI08N1jF7cY3TokH4EXGErEgsi3vHNuHIUux5W/q8x4uqnRHucoK
Hu2RSsmaX5LbvT1C068iJtoskEGSJqxqz9IKgDgTWaWbzXeWbxHrh/eSBlcc
EDvPd+nNezvSGEj87B7UnK+GvRxyBmGUUzAKsjerOuU96T67TWkUVekD0rbt
rzGhyTvc9gucHuIbiUy5MfHTYgqotUDASaAkjG6REJSjW3ZVfzDEmEFaEW8h
eHmX86X1/KZyaGxQtQu3ZNrhKzLbNgtt/jOo8O3TBMfpBaoIbmiv1iKvZUTW
nKvZ/P7BhwUhVbFLco1toiRflIHtCE1kOisSVV34CeVaNeL/9OYqC9B/GrE0
XTp1bqHz9f5J8eFkDJ5TD5FOMBzPZPxlRhMGUzxP1SEfCdKkb6LlLulTMvfD
HoP78kVVb8Bh7OTWxTk9YKWJpUrGN/zSXpUTgHpY0zwK950+AQCFLR4fakfY
dg2SXZjtvCi9dyElFfmbYAjEQVSwxWbdJgJ50BmHe6Jf+vIELNTeOEoyMDpw
fD/dj5QjMt2Oa+2NsfnMfWHhNKoYvZJz41jC71fKyB37GnKuFPL6R/rOVhoV
3mRFdx8pLy8XxoaHPrzuJkQVHcmVpN1fEApCWgUSm055wkel/t8nRQPM/Bo2
eKfYyXfJrclKRTr3RExD7sdnFa3VONBty0lzGoxbsZas+zxegAji3KnM56iq
3L28WawJP/nVBE/OWbkdR29P18SKqUBETBf9fF5GXNl9k89l7dG9fKRtZkju
8SZXy9dvi5p3FU4wxuZcVdCO0H7uoGSXRp9dIimXr5Rd8MxA3lN46LmerVcY
IR/hlqAlTuYOtMxe8dEcK3EzK7hBISSdhDI1Km/b0rN92Ho0aDto+2JR8cZs
zpD6K5gaVH3Pjntkd/uQDbfnczT6X9mDmA95M9QU/kHqK4kQfO8hWKfxHA2p
XC3zc2kUdiW0ilv0mYL6rOtyK4U68zde6xUeEKgWlVGqvo5/6d63bhMhdwzH
jhs9qGvJBbDkCn7o6Ot3Zjsz1Jj/HY03RzsDyjrFRozRRihCW+0HBRq0rddg
o41TCYV3i6Xn8lFd2E7I3FF+GlDCTPiV4WuaS0I6YBjo17gy27OIbfztbzuH
cqg7yAiGnWJXk3f6zf8ijikiMWn1eAozOoRpgtKhDcYdghKlDwe/SeHvbRrt
UXQs1Clv91XDct2b/qPQyNQURv4jHvaRVbCfZkmXo5PmI5w+cyhHXgFYXvZz
/ZEUK2MH6bKGZNe5OdNFxMaEzLjLsZQz18oEvzvIaArEzhOhID9EwPA6BFn1
sbF5gk32cR0xfyh7Rbh/0GaFPPFiz/JC/+RaPVVMhtAT71CDCQkCwjkHWAGb
YriKyGEbYMrveqzC7sVE5qzHNnKD9+/mht4ht2L5fC1aBLqje3ToucFVLk3O
2mZ45zVdOEu/L+ZvbUN+xXpIGq10AWYzZpbfg86WjsgDjhU8JE9iP0j+AhM9
QAvlKzPNi2WxiYSD9uqT4/g5qnnY+Oo4kFzMRrXGQo09exovVOe7CNO7oX6y
HN+DS8YRsh/4hWAnkiIiv+5cVo+ScGJCk6uwyrvDU3YD2bzitOvxc02rEA1+
p+p0nSecWjBm9/mmkZXoDdaQ8d2vD0YoA64IKRfJkdSUumQje+XJiGuN9YKs
YXGNDmqNC++FUi8env5bhW2X29cGjx/kjTyYNAZEIVXpa3l566yfq8XONW9P
mju85ZlQmYaKFeGl36TL96ZzkdusKZ7heYZXbssc0foVJ+1Z7kNzqEXYVzB6
fALDlh+KMXVEoZiGuROQRlEx0Z2CAsELLl6seQyRR0UhYejZDJ8zn801Ze5Z
i9e76Rsd14SYYlM837yNt11Cb+4rxis1C9ZjqFtStIdiv9Lrjwaf9wCLByjC
einOao83diqZ2V+7EB1ULnuPnA3z5zaxSWa1Hva1nXNxS3yYZTUT9VJOZIMJ
UhQEIIUykOz51Ez8S6rVNPOhMLn7/BckLPoo+RZ2SYidf7MsCp/ayC1UJvY1
7GiNQjcM5JX4XqQhMWSO+bWpc+8/vtQ6iUU8t63rEZ1TdMnkS1daci7HxKhR
4mIsE0q/erIaLCn72pKBGAhCFzQG1tLNHl3G3mWpexPi68mHFyXxo6rKxyU/
NYY2ZhMjHaOsiW+MGh66yrOf12GelAvGayleywYJi8ssMObSKSl46NnmvO03
Xo2AID3IJWX8ayq016aau+8YONps6TRXGIPoT29PE4CCf7rM9ynp1XsQQuqh
53Q7M0yxJN1OD7rEJrP8mGt5b2wNhAVuf89mlBOcy9usmGIPDI6Vxi/1BTag
A7FHdjSF/3zUME+MvEPI4HCeIpeUHXXwRoMueIVeuNX+GGL617bq8CSJRSC5
cfPo74IRkdjo6uLmNfmzgJSYT+WzxeblyWc5T3LcliGrEUVTLIuNT0K1+VZ7
Rjh8yqB60Hm7vjfiFhz1bKvvzPYwjLI6H52fFhlFxjRkAuzl7d6Lc7iC9cZT
0Im5sfImpaKJZgK+H/RKQBLKQMeYQZeNWBL9c3roggjudYL0EG3BLANi/MFH
is7/NOJbcgiqtXklbHknWUM7gSoOfiX3cKyO6NculP9h4kWgZEW0XZYjZc12
P97D2uoHGj1DvLn9qP3UV5dJSD2EhQLv9/hz67YfsI0Lswyi/oARU5qDpS7F
mnhv9d9DVnJ1z7j6dZwIx3c0NWdcXn+E+5zsjfTCBTnK3t/fIW9aaQ/I8nbJ
S/2ypbivmp6AixbapuU1MHZJA4wO4P29orDNkwLs4PJmEYCXoggKVkb4Bx+E
VMjpA1jqp615RRtgyLnij814/4JzONbVY25YhEt0aq9hPqM4OYf2Gp0/4kCd
zyaaTzl9u/md8VDIX8qgajUtNLnksT4ay28pmRXfXItE88oYXqP+Vg7ETZdi
HCQ9jne1mwjqKaZ6tuMXFKJntFv4yvajy7AhFTcEC2rnzeQPaqrFdhrmP228
xpEFA17X/wT/kkyV+LIJxRi/DT6OubnM+K0tBf2rNHMNFLpDzxljzp4ciGbY
I/caoJT6mokxv6laxWzctt3J92xacKPVky04UHfgwHZCAMhBG+JQtU5WEAln
0cMAliuon2p+YWNfUlQ81/eJEOcz8OimuKvqM2j3AEhNCRO1XzPTdjI+HSBB
L8TvggRy+BE3VYqrOl1H9O4FPZFz+Dv8Z5uOzisbVFkcF4mdqhwpRzJXmWOc
41/jngFLOovqtZl/FZPnLMIKWlVk1B9wUvb8aq01UWlMRq1216Y+7+uhpsS5
tHc35R5iowyJQPZQHmx4C+pq6kyUfgLtqEYxIE3BiMAd2xyKU3HtEg455NYG
fi1YMO4w7v4414oQIx2235+jDr/bihJmsVpS0vbXT/Vqy6EDCpB5nfgezyp0
tfRLbeEILlbKe1IjqfxMXilpCbzxx4Fpvig/61gO6T3HmS1ytUvltUJsZem9
OCxwZRLFVxCGsD4eaOg+EJac/bFE1K6+Aarf6FoK9v3RoJXjZIXVP+vSJbiu
yNtcDtyNz6o9ta1OwM6HsNQO3MlaW3ms8e6gpaCHSXXvj8Abpt8mLvCPUM9U
TUZnol/4NMjuqZDFMo9qpCpMNj1KCSCv9WlZQm/MsM7AJWkd96zrLHN+02yF
i6Icy4AZZsCMjvGzrT8/aJHik0lfSCGcOxTPfTY7kwbQmTK5BkQb8XHVwMOq
SILvwMvnPZlaMhScEK2ADJBBRZ+q31WPvG3bs0pQiHV5HmYytx5uoOnGXXtx
WDcDqRTniMLSp1kUGJpsQk1UIKhVIk1Z2OoPsdSQbSynyVkr7RXmZiNQ1e0N
Nuixr1gzqT8JDVJR/LJAMW+xmqVEYM4zQ3WpPaBAgyIWHoIdJW5qZKenXp6d
62f6e+rsVzfkGCnRUKb3hoxCqqBoQc3DO+xWVceosDmlUF7jqJtgAAL08xdu
/aWPzjC/YsY+xcxb856uoCoBSwozyKoJuTGlUNIiD64tlpXC7JNUPX3X9gnl
xG9QyZzmkRQ6AI6H8ABUqkZ4e9jt5zQnc88xv6CtfAzm7DfacXq/pw+F2zkn
EFfcCXRnREP+OCulm8s5RcV64o7qH4QTimjifAhD3WGXXD/BRRKb869QoIDg
5R/wZedxu5eNrlhSuGON1rOe1n1od43rDGJUBRH8oQZ1SiekGdaE0H0nztn5
krsdeKGaZiZNM1iHBO3gk7zpbqvl6LnsvcTYGgDGtD9xY0mGhbvfPL6LGGCE
Az4USVi/lchecnoPttnnDsGdlzq7ZMwsZpJTuN8cC37GBHvsJNsPY2Wcipj6
c8FQIT+OZV+dAXncBi10Ar4uvR85L2jv5lDS9RFGgqyZN04930FrDiBLyoZC
HzP8aWMCWN8YWAbYK5xnG2wbSo3/ihn3ngTOlkIT3mj7lOiEujUzlWd/PR3i
F7yXj+yh2EvQw1Edlt89uEK2SKJndm+QCyST8sN5mGyg1eJbmApoTEXEiW22
hx0HEv+a+J7QNI4hDNFj/hEeIwB9KgMdTAtFztpxFGJa6/lKnZL+3nkNvX07
wknPnplx8WTIU58QqvGkuE8ZaIciJCeihlKvEv439//hfhf85L96ZzqUzAfi
m1FUdKYiU/+sdHDIUaNMSX0sAB0KNyk/o26k3poSfJ/tCx1LKbXxd9BuQpdN
nb5m6UFIbrvdbJwLMASVp8rzqiFSxCsMqiTHj9p1w9v7S933/Jhd24nbY1Dz
RFW4U6ljNAhx+lETHMZ+pXndnihWG0wZC5+7fglIDf83/8JxN7Uehj7IIPm2
xELfH6bc8KRDKN3KStwkVd3IfN3LOqXjHyURxjcrdqdV/BbCvVIwyJPktQDN
03NnOp1xmZ0siIR86KHQoKbNs3S7XObPq9FVuBntfIjbQJq22Z5yygxIr7JK
O5z87nO4+PXR7G7prnQ3JzUnX0SE0JhboPznid5ZknNxwk6WRc9RJdfhhQNo
+fJ717cNhQBr39Smhd1G+RBtfvhQpK43+yhvdj1OGgeLwaPxJNnxrHAscISQ
YuJGnJ3ww3RPhjo5DxzFZjp3bJa+BfMu0bX4GNd8c9iNT5pCei7daAJEtRgI
0awx5s2rO3yUrQ9gWBHAWBS0bZmUEpkjNVlZn7HhUz/+C5LdvF73/Q3Gdtf1
m9lxZnw57hlLW6g0B7hkmDEF++BSgnlp50B/NNcOP+WbsznME+vhWtKWuLsl
frISaIpMTwSHJTi7Ew3MWhbJB+Taj069vuIc5dBfYlgdERDKdHjC9gkqV/Kj
Qo9nu3Y9hylnvXhJwxw4999Ujl5V3kM7JFQ7Bx+WyWI8PQpwJXbRCRqc/5dW
iMhUXwOP2T63KmtMIXL/bZG37F2CLPp2RWt6goxlB2Bdb7XV8nIGSYLBHIDT
AD+nIyrQ6eoyChYpDi7IiBjwozO1PCOu1DSw2dTydtsGSCs+Z0C7SFAmAxvD
7x3PIIaRzLXqfx7TjFLL4b/AIaE23/DjeaUupWH2qvhaDfF0y5H1IgoaHasK
dba1sMQzwfyGFqzRdX4bvMhrUeYaET2EUU6KikST+Gs+rblNo/PvEa4ryqgQ
JpJc6k2i9ZIF8uNSoL+ZUdxoBWcDwi0ez4upHpEPVNPen1ZhX2eVBM3RHyYL
XjRUWxm6xaOKpA3bobT5j0TJtv7y0Sn1s9qKZ+1eyez5Rbb9jDWBnxrOuyl+
yZHny257A4L61wgFZMlMVA0f26Wtj7CDVKTpSCbkRbLo67/cvWc7hvHuMCIS
EN5SVhEdtK1ZG6unPekIbMxedIqmGfjyI2MTTZUpHJUTeV9JHtJt8mxqT/E/
ecQeWxj4TFFZB/8JOfJvHnYFcJWV9aElbDmRN/+t0jO7lXLy5p6fBuPEGb8V
OEjgdWfkAVtFzfnGergJcU+KPMyrLysrlFXPJgv11yWz7uFOsZmm3ezqJhdM
Jp7tCFhTIRG5gFTO+ynMIzMJRJJb7Bwk/0K+O4TDJSyJj3HPrsUnmJn7r5zV
Lp9ARD7Rx6qnTtKJ+9shq4TYFK0MyapC68TI+vN1EG2st9KjFHextEvtP02g
yDC28SsM7F2AE85hgkuhcaY/JTeOrV8nmtGWeSEMxoDFWQdr0Z3+d8/JWe/F
hMZpwqGLi3aBGgGQwYb+D/1CW5b4iGHrgJQB6OQqKABmMUC7f7GxKZ9gJUvO
sbniDprGhw3s+rYyMRv5zXOTltRwEj/66/FoE2Jg+ucKmXB4w+sJ6QC2T0pk
D/O3po67G/hPNoNWACtPxLluBpB7kqPl2tjtipfdiQEU2s8ffaVd2vGZF99d
DUoadxE8AX5vf/ECIFkjedgx1BXeGPVy/Y/qqOwjApMDq/R8sdVw9lvDNfnM
siYKIih1o6BMLDh7FJjCWwk5Lpbd/hvd+wnVmJjcTxszvreI2Za9nyFl7CF0
ctGv6a+TwcqhgopT6sESjI1YH/tlqT2LdA8U8nGDcIwMblmtz3naCmCFW34S
O8aEoE0ISgKtfEYyjd1uyd8g5n2XNMRYauD1AEKMlbugTFK/qeTAREbPbs6t
2goI1OOj0hlvaFaGP3jFtImxnFfFF82d8gOMCsLdtHyJATuTfjVHHlDX01zW
JrbOSBsa5z7uyaWarzjLgkcU4xUqqBSPb1lzsG3twtx8O64/onkHcV7fbN/R
pI8fYuNl9QtI2VJxhiZfus3E9Ob+zPtGkj7h2c6UDBz3LHjyNcjBBUSFakMu
M4QSM9yzvS4MDEn4ShxYlqxyA8xqX3wTQUbS2BDa83GAD0cww2lEX3ZYqtXm
UHEysXKVB/w1sdZgCovqZUur/5MsfHEhiYhZ7YNl5SQ+jBT283ULPAO8ztE1
+3CD1CQ9xlfJemkYyH3l8dW2XhBgrb5prRPDDDJpuh+emwJwyfwFbXpvl1Lu
KYizF6/azadRHFChXLWCRZxDg4RyXlyjLU6c09Vq5w/7BpAZvP9BG0YezVEw
AuaLNiVz0+ZUVoDMJFYZNrtraMiSV6JGZD2zaQYGO+Hz1s8eNr2I8ArIjxya
16dz/RXNTgsNXbT1qU6ra627ruhd8Hhg/vSTT+cvvPM78XbOxIsIMK9wvNYd
FYF4qZR4wXBBtH6l2KMOEwPptkVd2cf+hHNUDiLq5Ckt4fF9v8Mfv80wWEnj
3HYp5glIPDD4ji5UN94x0qYOxH9DMp0KY8BRVQqUBj2o3JCSr0mM2Sg4uME0
PFV99vts+ADGpMeRDK0VcAHSmIg1fNc294kGklx/QOqGA6jTeI4ePY+XUPy8
ccaagL3A+O8CmE5SvGUA5H6PuzC5GuDWZ20Ilxp/jOK+sNOmjJhd7o2gcyfn
WjKbwN318P5O4n7pOMgFC/JuOaAix2LRhQCP8FZfm5V5V2ePaJ1bypwzn/lf
2QE5gPfkfLCMzI3UFsmPxbq15A6NMznyeg1XrRZ8xE/oLnADq1Yz0s+JUL3D
+DliKyCHqAlPWy/JRLXvnfq6QtEfafA1V82XTToMC24Zev4mRyyoXAGHgzNu
5q97VbvaGSA6RGviRtBMhSCA8VPqIRG6eGI+DAw6+DPqu9+V/eIGRMuGNdhH
hQ3c11jT4zWrYJz/s363V48+fGRxg6vRkj11b0OGYRGTCk0WAYl+7kg44s+k
rNv0CPy4eRmfPmjK/IShcchV8C5VmBK0JHSgAm271zBBVx8M2PT8FSvI532N
/68ZYZPUK2S04fDO67z3p7b+5NPqMSP0ZAZQ1++DOYnroWZeqsRhCmuPvy7r
07xyDkHs1enTEfW0kniP4dm0DT/pXx0q9XiLyZjy+p7vkf7JwSHn5Nwkz0OC
PNXLDnzlhDpRd6du8VbtGiQsWlr8LyXMJJwAX5HX/xph8UfOU2rvjt+RlHxb
C9fdts7m5yIeH590ur1QYFB6/eStnVuok35FQoM0ErS6FOE9LnstXHArKx9w
BOaLlaJNqUr4op9HEuiFZctF3ZO0huR9AFURzLOW0fvDM1VMCq3Ruh3t1T16
THj3RxkIBZ73J4XmBGbh8bSuhhSJ/fHuWWib9cL7Dt/PI8Hkt+a7VpeA+Voy
zo0QvOM6WR8neiXpQGL0Lv5kJYS9jh9GVrMOW3HgVnAvSwjusYSxHrV5IfWH
wGI1sGzHrFTdokBEbv+ABGBlxHOy3+moKWErjARColkrZmpfwiUOabbdqDUT
iKl1zL9tJ20LOHn0VE926ooI5EmMCFnI4q0oiM9OktBkj2R9SC/rEooOipLb
ppts1+bByQzwmoXqsRT8ctwQyHJ/CoJLhLAqhB7ao7hrEN4kx+IzQurSFh/X
Vd1azuaRH0w7PGZteVo7TFGnvUILkei5zgVu+xxYYLGMa7U9S+bLE00v/V5g
p50Fmuzs3pXOVIKnbPNDK+dz9xBcrE4KQw7CsKKc8frptR8EnVwIoG+YOXYB
peJhE2ck6XjVs/W5O//2IAu9xkKsqDp35UEE4Qzc4/zpNXAn/Irey6cyT9u+
jzlYdxiE/hZm3tl9qeMLGzOQykX1TMlj8jVqLEq5fgRRVg6AaYA67qtGC6uc
/NrDXDTzcnoEpOPzXaoxX8Gm6foTmwN5iGx3GzpKxuajwNIvxoTn6lxNURqc
KFTB3BtRjgs/6RpkJEs5yL/DpsW2ilsuKvMdC1AJiujlF2C6tj2Vo4MdjYmJ
HoezimeafRtBLuhOcwUO/RlAMMQdDElEGdIsICeUPU8r2Hm6uAxEalpCIW12
HaPnB2FEXEwsEHnGUrXk48o73SMRWN4B1lJvXNYEVFYnD880wY3OfSV+lmCz
jbJGSaU/a8nXVGdiAAMbfSqYpje+Wnd6XhcqtwI2qKEq6f3VYgpUQx4/2yLF
jDRoo439pL9DLpR/Efb9tWGSA6adigz/7fU+kvQA2pcykmcIV0uvqJAv7wzo
wlHKy6PbHQyKoQP4FvlZMGdKevmISAgMkH618i6Y1ABP9euUMdSDL1INdEC3
+wrtcmjZuCMzOjFE6lmFq1lhjraVSjd5WV1MYFkh96ngr4/HGlcaaXDR07Tq
x4qZyUak1L/mKKeJK+0i1cHgksgMejUC2rmMO5tjQE6T2jGkUVUMGJ+YHe4L
Np/77TGY5hLxgJudCYSECpNLaPXSdw3crE8kkqmcdJ7sn4Ay7Sd7TKbgSnKJ
F2Ytxc1J/NC/x4saZr96YOFrORRgecAhBbw37aWWIhc31ZogpZAMHCkEmDWI
ItHapWTqrb0oODWC3boq4Pdxd41kYdOMHAa9O2KrpLOIsL8Zt9Eh64uIwv/7
bARm69wiNQC/h1n9G5tL8W2Qg6OyuR9aXegGWaZLVrrSnVM0QpanufbOgsrR
ZqPM6+VH/LVwIiz4YFvr0byGVxNY1TdJBbklGB0U46AAeGOc3xg1egHIMiVq
xs3D7Uyi1YpbNn4bEsKfsKaCVFS7lPEhrS587DU4v45y2yhYZV0ZRsyFYKNR
92tnrKLq0VqG6aCoq61pptF+8wgbdVTdDTGoOPkaSJ6v/DW26bQHM9rGexag
0dj/KVd3uEKF4inMJM46k9VJ9D3y4UL5USgoAD6+sCsvBP9Mc4mAwLXpB9FK
v7z0x9v/ZWdT/ZLoUc2GfOcgj+RIRg4YJg1N3DQD5cuD7Jxb2G8OcK8aMG7F
Jllx7Csq3hQN1LqJASZyuYY5Ux24FuijSZK9DWaeyp3H8f/DhjFOSf0Lxzue
9s638iDck3VAOQkvgpzfTKXXZ28nKcXNMFWRfGZAgaMbQPguGQQU6bzcTU6r
Zz4immrK6py+FU6QWEt+xkt4gKTW3c78ghZgt1RPcQNh2wVBZIiMLgSPfx9t
LokZIWJAVJtAQpBEtiyAiIOZGzXhciZPEvKEFsZx7/Qd/Km3DyasfI2417ok
ZDKSF9Xe+naXYjZ61ncwaxNU+Ab2ANFB3Qhvuy4fJSfMqmEZh2ksFmWOU0q0
wLwLNnOYxz/pRm9WnDguHBptXpB9qvMcoB8yv18BSWlNMxtU1qqg/6w0vlIQ
bhGpfYMokmPHShNve9DlN46/qbDGlUWty2X5ocmPKZAlIG+isx5JQogA2/DY
DK+zvRSoWYAfOFAu7IzQcdoK1kmkQlmkPIJsIUREaw7qB6h3OfklmgF8sTdx
hjdWEqV07B4fTOBG1eLe4CXyCiRYkNqdxwvHUT8E6R8R/+US8NpApn4yYF3n
WfHggnA5Fl5eCso9yaGZ6LOjOArA8e/wPjVB7DobF6cQ8o6k+zhsmMzsn1fY
aM98HEmRw7tx3Mhl/CpkP2/qMAaVRXDXSgeqreU9HAfT8fZGU9dT3LnmC3Vn
vh9PMSOOxi0eNuXcxM8xyvGDaPNzkHw0mhLE1oL6aymLR4CEleu1rupouvey
CB/0/YRnwCbI5CpuTsoC95SHdoyAxn0RWn+Evpc9ZKKyU+HN+bLR3xknHqKO
RGdr1lYWPqhYUryFlE0w1dwdVQN6K4koGF/n14/KqtgTwC25WvzVnGrsEg4y
5jfKSdMPYtpBPJbOO14BpEH69SlkDZHUHI3B5OeeYTjGr02yFTQQ4oEvjza8
z85Yl0ecMj3YvOdfuAEIqdJlE7PCOa3qjLOt4qy15mtfp7AlSjyJA2eaO1MQ
Auui4TIkp/94W8EqMChOcCjK/3kpLZ8zBHimWW0hb331MHxSq3kWbLWtWn8X
INU1bhBrTzuT08rNE0e2ZztJqfeRi5n9pPjFR/T7PWGUXBTFw1sLAjnamdVT
oB1uvm1FyAqC29ycN3wffnKGpKFgMYnO0KMqqktqGjybaCDzXCLbnnMQ91q+
zHxJaiHjHfwaGe9nMeoOwKKr3wPk0WzhS3N0tIIR8GVeHz3V69m5vlV0AH/Z
G88J9dkErHfhE49pKhZ8GdESL8P3kwLnUFTQDjpjjYF5Xkt+kFXt58fZYjkZ
Ix7xkKA913w910tZ95NElkV0VfeVPv+ddFCN3oX4c/38HWIFzyMJX/mV/kca
WaO7jZaEnBxNHTsB7NnZHwTk/3qP6379WhfHwUB3WIPt72syAVhTQZMtJlp0
Q+ENR22Mau5c0gwKd6tiW9NFijLCFQpu+bOMIDULV0hlsvkdse0D5RZXrv/o
HHoIPmnuX/oVFpOkBnpyIP2iorhz9xSOpcNPMif56dAJYKcX8ySvpQubw2+B
GpFeU3ls89akb0KDxYJ0LwNvkzb30XqoKzOXzr4awugwHIIFmOGqMs3DfQBG
7NYc00kbuDg3o1DRxmiTFe7o7Jpl1b2ae20pA4pBs2A3SWEClPZAirew2FS5
H/lQl+WHrkz783dtOI23E6gZ64q4CAXNX34BcWl3g+G3Mp6LXYUkAN3p1xJy
Nlcm1QtKlIIvmvLtqvux1/y2YpCkLGSRZKUbCxCfH6aDdVqL7iwUPToRlnKF
kSiu2YYgsRfIjdLp2kuNVfbgRjhQSCExaRks+WEHWoPCfXP4p6cTStem+RQU
2QZJNI/lpluSY13O+dg9SV5U71ONyPCJY4E6DJ9lLQ5fIHRYO3liLHZOFxtP
EuwTFNBj/u3UZBiUNz8USe1XskDAhBXK2IDl76FXOePQShWMOxlVu6109bpU
mnoxmDK+TW+kT6ac8SBPgQTOECdURMRBE3JLZvYWVYYnyVnjGBacZ6LEMn1e
BGz03rzqPLMb67+Q4IIz2xPYW+Dlu3Ju9fvtSS3x8iSNkL0OKwMoMtSmnLYn
PES05eqnwFk41Y8qMprS3Dr5eFX5XnzoqAFHYiDRIK9toVw0eB1ovZCaSBek
uSjsP0XTE8hy0Fd6DX2L7mZ/KuPHetXK3YB1lbHdyXprJ9jfLRmd0bQedIhl
ak/BNgrNESxSQgeAp2vOpUYQcd1MGMWUJJRRMsjjFAQyqac/2VerjwoJ3c/Z
ypATQPS6416lR4EBZ5NRjHv5P2DaeqBfccrW3q4uKTHDYY6n2kt8hoOvqwPO
2b0UuGwD12dapA3M2lSRbn2iZ8LQQ5zQ1KX9sTyTWRBJibA2W6pkx3T5UUHg
txMgQ+LyWsLilE06FaqjAXMelAPVrsHr9BY3q6QEGydKeemc06HCUdZG3LKu
ODna0Gdnw8I2eF2ra/8xA7Ya/sNWJmHjnT6aSoJmpnTFay6TfggGKoZhklV5
I6i5rZm/QubR+BYmE/gQKNF3U1xJ5Yveo8YUu2WFuD7YX5pCxPACRA/eBdyf
u+wqPxJD3UgM9tv0++6Pj3AAUuRs0+n6pSsj+viWPBIJ7tnM6IpXylIGChHz
d8U1CRIQRJZP5iEygk+HUz2MBk8dj9X/uOXlr2d52/bBRb+PZaj9+DZMX1BH
I2sQ59AH5/mT3OCs8m1shkGL5kNA2+T8zeMTu4sTocIMS+LONjbBRpdaF0va
dgJiMRlKSJmW53sjHCa7lzv86iqgH/t/Y5ou3Wu4wbMw+LffUmvNVQZ0/iX5
xJzNJmHAvhz3v5eeKhafVA6AXMC62Nulp743kW04N8jF2aCw2RKoomoR6i/e
oRSBoepeqx1IIbRb2iLlyFKqhBERwMcD5yMjjtD63/X2S9QcMNAWSecSuTzB
UER59nhFLZ4vK6Yi1XqYYcKc9Fszn7dWOzKEL1iPodgmtKZPbk+Y8RDnk4ww
VFhp69NU+ZjPfTAxfaVwrofM3G761MsKdvAyAdhsEjPso9TOIp85+i1jKqQa
+PkDiS7m9/KzsU8qxORQx+4OfL4WubF2V6m1chrV8+uj13AhMypE0/OFjvXl
HtEw4TlaNUGxg66cz+Nx+lIJnWe5LWW3C5h+MCmR8LapiTCd130moajfmBuG
P4dYiuCU+YNDDPlvG3sDfZxtsfS0TpTLlCceOpIR0R+Ha9rrYtcJ5Ro4QrMH
hatJqa6nyrxitKiM1VxD2/r0361+QqKKwUiE1LGlG/s3SfluBpe44nZxTyGy
R9FWHVpW15xoQfE9IgwSSq4lJGME49L3J3XqtNj/bLJCASx5HDt5Hz3piSOS
1biCUB9jn+shI+pGuFvxU7NUqlogeKyOuYsRDqnq/pnhkGoSuW/nlk6v0Jex
cGEIS9zHCnnaU7rilOEOharJLcmFt/t+G+GV3rt2kM+RCG1OzeKPhzRVDclG
FPTRybw5JNAPfuSOIWhl/Egs38oHH1WGY7fZgCqIg9QTVFg9/uM9Jlz/YlbG
Wh5x3sD1bBkQS87n0GbvSHWaISDL5MECdSaziXxSJYlli5RBMTByVg0dSzQl
LCAYi4UQIaVOSBWaEibWk1Nm9r+2Xs37Xlrt8+wbeWkJc1sLDPEZv96X4hqQ
rUVLKVyxA5STYT1mzPj9Rniqn5Cblx5QsslCQwouVo2bGrW1SK/XMiLarWOJ
/c2hBcHd7dCzC83aU3C8t77sGZ2qYETwYoMOFIHjGHrTQ9YKDcLv1MJBTLOc
Cukn8L6qna8Buox9zfh5a4CBO5hwmbYJd7fCpbst97ThmSCirjzOo0/FfTEX
86LBWv+YO+mdmIUcMEvQJ4mqyIQW/nZQCnFU6MH4zQPegH/DM/k9s4CwjoqG
kbod9lXZPnMxFm3dOCofjpaWDAoyiU4sgHiE6kdaFlDwnDHjRqrPBedJLr03
jkrbPFE8fX5/z/GXRLOpiBQuYJs+xen0NKYZN7Uqz0r7jh14F/bBbQwxUP7/
WAl5FzGbsVl8Ky6q3T91U55IkcHaZd5JbMu/zroisUouxtBtUyIgFfg8EWfo
Ji3H7Y1pKz0Ri4kYR2mOGDk/X/BPvrLINOHR9GMO4OdEd5ah3UWLyMO/o9SO
5nkpgLeSP0GvMUqbU69kOcG7c4Grx2uYMs6btp5q3D5Kt19oWN6LwVv4buz7
nVuI5gfVvhM1zvY+Lrx41s2jV9OLNs58lg9fJ/L/f+Vu6CJ2tuVVrUtiosLy
NhzohJ8QGlT4MH2qf6Wp+pMaVGV00BmZkJadp/dujMn+WZ/s1eokmlmRkZwo
+CZRJUI1Pl7jf8Q0hKuQZEp/wmfPiNTPxTHDhFCjY/dgAGPwI9VFwYu0ijFA
M50m7pacuKtLCVBW30wr54huJskSvzZKVLT4RZuwk4U2dyIhoCaYIgual2yd
Aq3TK6n0KVToWReh1OmABkVQ8B6hgFX2bPrR+4ckAsP6D7Oy27HK7JLYhVJ/
BN+3Ac1mpgRcJg4yKB2JEqI04TDN3BookdLY1bC4iyBXToT/qmJCd+T1yoq+
quiD5WPSBjX/HIkbJACLEINQwq/MoOwfFCzFZXKufEOSpk76C9Pjm3Dp1RJB
60YvjmId86eOvMeQ9cCIGSzTdEnPBjfAe0QT1xijQtqjaFWmo7Upvpcnt4Te
48IKEEN8QoLpop8HejH/mI34jCHXQci6N3i/e7YqpGz8LqVuj121Ywinky2v
aOGeBcFhRMmCCFNS69uyg0JOVGsEGjNNm6pIHJ9nrwmoYT8TcCK4qmz389IO
PtDrEWlkZFTvQ8gJ71NxQVzzdmtXP49yfTUhtHmrT3Mtsow0QgRnsTSzyuHM
q4YFsBOKwNdg3m5fAgy17b48OdNQVsIkQ8r8zu6W90uncAbvcYCbdUv3ASJq
2P8xtkgWuBSmZffah10nuFw+haDY97rKcjlJygMKyHHUJJ85EG/TAC0yaDSD
pi9kPR1l2tVDiP7wawc8VoJ4NYS7ep8TOk+96lgz5TQ6LSRfk0McHY4TmiA3
+r/YRV0Mo2kErKk3x0+bs5CKbfhawvVjAG9pQIzZ0KErVOkuu4LyaWqFlGuo
qqm2/HCqV66nEyQXfeJwLIhYIAN2Y1BuYxq9a4ZwCHm1p2mxZIEKoKsfKRAx
b5tx4+xgZvPMZ4Jhz4fDcUJ7dw1PlDmp1gegTUkEmnlK6jW78XX3alj84xDS
NxasxrFG3HlLiy7dlBwN1uyIkPIt5d8aBbm+imZKRPHFP6YfsGfaCRi/SIFB
1uRf7KMIy75iW3NIpQIftKx5UwMp/w4kYQi/SGpnZ5vTwZBk6dfWAWwKGY/Q
pS8i9c8wfYAY/Eij7u7Vi1bhx2Pvciyl9NR48Ol6RJxINlkCK45yW5zGySJe
TzLKmU0A/2cvnsK5cd52I8VPuZOzTzgxJwunwEu6DniGt4hU7e5VBRLraqW+
ZWhPCR7H1TNgYKzBmOPKFXNVIfBc5cD7ZH5dnKjmP0wYyjlcQxDPE3c/6Vx+
iCIbKu7+0k76f5yRT+R/pIyLoiqCJyMEa1OLH7+lUDJzAfwvzSzKUwnHEGMH
izD7UtmM67B3inbOGyyGe6R1igr1UILxmjitRXVXdRuV0sjdC/TTgiP7hwq7
K2jlZ0bHG2YIKZHUqZgyIEynxW8PSWUCYe+1bA9MppXJNos+XxAa+cozsM6F
jOs8fVn/NAWY9qMc4wI2nAv34wb2pPQCt/B/9iNaaUXG+StINqUniSrK0eOX
OwKiubnSQaRRGNkOHFsINO/DU6IbNPX70hbxJEIO7SsW0YX6iBmBIp9W7krG
6NcVdcbNhrtmPf7ZXSej5ScOihoyrrzi1xkjymUTrfx2g56pjdLnXOvy910m
NEkIiUV/Nptv4VnrYM9nJUd9KMGkxtFcWcoykDWRus5HmAkJ5aMjO4ZNOKJH
UkQf9/7LKNOPOLF9YvoA4d6KrMhL5Ysaa/gTTlrfzmr05Ut74u29I+cyqueo
L5/NAzuLOV/IO15/V6YjfbVY7a9X/VFCHHf1zMLD7qXyb/zp2yGizUj7vH/l
TiyoLt3BoQVM/nJkPZ9Am8rBLG2yFngMK4WpofgDwgstvdD577iHCLUgCfUt
FFSmfS4Z1CAbJ0nlAhiA8QkKehoyROyE+9RTKAzKEyceGB8p/tz38KArBb7I
IITzPPnfY9xUco5MFXHwI8pdh1vQUK4YK/8BHa8LxCbigVe+dW6/mj/K84rX
jt+b/lsAuO7BPBnzlvZ0Te/9hcpVgQRW8aNuvXWCe6ACIIEq3kuajDawkLxK
i5TrrmEOfa8siRZOhf6TqN86d3NEWMMVCaa7XOwcKZTd3JDmr8cM67NK6VuX
VG4KVOgot/KEkZtEuKLdCgUZ0aUfwb83Dq1oKDIfV9GAikRYiwks88PJk+MZ
xq6qlPcJxiD2zI0MPlH0aeEXb9l+RJG3NmMkDi3dtrF/XHD/lGDaKpKj1Lsd
O7H8nX0NPbojT7VLV78JCDIcXfOn1B9jV6kH8Am0c82uGujrcci3IWw6cq6k
5bddfEaxkNKqdJNt81icgRnERZ7pdxTQlUKg3a5bUtXCWnpsaOJhmcLTnM/j
HC+OJrgWUoW9lpED3pieUTuT3MbMUyIkLSeDvGAnCdnDBWb6L3YNKpNL+tkl
C7xEkYRleywijywr8pbMnyI9Kiy8GOuaOCqmZuDDLXGQDL5w2Vip0sNiMb7c
wIjlbTxkway3+rYbPo8tEy4PwjSaRdZ7K549HvGJy+Ka41G5SlmOl8/PSTRi
A5M0XvT5TculnlqC05kgGkAnQ4l/NJjsUzsAQKXjUjjLKnkUmNgVxRZ1JMkx
yUHJVyevzwl2m2k4ay4eUOFhTiRLHqR1rg7Er3Q7YmA18jzzJ4WXNSf/is6m
/P/qh3DB7uthzmsnKP8pyvesk6AIWskBTd+YkXnpSC+hFwpszLzJg4TXXNgP
9RxHjDvTKucDpRCBAIMTv2AzgEf+nCCdWhga5by6x6iJI3sJfe0P92CPvZwL
8BlUpCA9TxWnrCjCzwLE57aHp1RKKwyQtXNfnevWjPcmqWBvB1GB4cen/TYJ
lZXIaXW+YsIePZL003Q4VLxyIfcqOVmLlAuwlwJYUU6EajlKmWW8zDpu78lr
J1cy/d3DvFeRyDq+13rFrenoEm1FCkmDwS1tAgZ4LLDqhrPNJvZF4MKvsqa3
mXqQOijqiR/nDMPbXLOwpVc35ieEX/a664GNXNztS9jMzI/Mvs3SKEwGURYc
sbCy7heSrnE6yRqgDY/S+/zob2Zpi95a+TVq7/J/7tq9DcPIauLjar4IKnYi
jocd1axxvVNe1zUZYCBDFZy69dxfjhUzVSPScHhrxXLy/nBy6P85hoQ5Uf7h
p4SIHertssoIrlMHI+xLV68nUw63aM61qkqEwa1p3tNh5EVzraC52pLpRe1I
cciCoJFJM9pE2xwTI4FLn0PTw7uDGpCuiORSL7wXhXJ9ai33eWEM20sj3HPb
meZmNqkaR0WCjng8TkWqO9iG1cWGHslIYnSXF/0fc7tO59SJP3Js4SJf9UF3
CQIADweCvyOkKD3Bb9P+A1MG8aKEbBqc8OhkFtHxw5a9+u4BqciH3UmIjQYv
lMcA1x2/sAuy6ogtwZBjZGDSr9Lw9RKi9VmC53XST+q7kTNdpPQrUrP46D8Z
4GcHDbRJPQcSnpgkcpcvFzzGe+Vj74teOP8QWOspHtxLJY7p/UG5xhzc4SAp
cFsr4vX6PJmURoETJXSBX15rohCqla3BGmx0IJKGsv8cgqzsTOSUShOzw0a3
kPQVd8HlskWGTOuScts75tOOaERp9KXCpdHGDsU2xW86leK+fzXn8Y0oInSV
qV1uJ/S5m6IvRl5F62Ai4WexBrsIu+MS9fdOn8bApZkQv1F2MknN3o0GZlJO
/OoMvQGBYgnCHKgn+7okm3gPqtYTviH/jwv2qhIS9uYo3i+UONFeZWFoyngs
ixD4y94orwGtzRjZ8R8M9477WZsEbiXM6NbaPVcmTezVI+kwqgwbamhOTXKY
+rMak+paa8M9y+mWi5tI7fntNmD1rdH9GbySDDnjNRYTRsv5QV3J9tImaL7X
dXE5vfmV3PBrZrV3ytUoJXUwMRNlcdbpBxYIng2aiIMloUbfIgiKXHurorsb
uMKe22HHlpzICLbI1djFLtZal6DOhQ2meUaWHbLqxMluNVoRP6LXmLvLlFBp
RJVpTQmLAuzgeRh8OkhrgyBnhVAN77K0tp8e0zNeDwTGOr7+RVCziscpi8Po
BF//WPtGMyqGQt7eF7VUZ1yrU4YhQyn88o77RmygD6O0dr7MuZe5xplYej8C
AjRDqun9xhYSnQyx0UE6BcmHn4mkHroI5hWl8HpM3D9soDoV4LXLGR9QXcqY
HaJ/4f7HyIGQ+mJxw+pNUVGNk5kMsuBnlFIfUcX/068dNoSHuPYdKW/rcU73
KRnj8TYeREzvHia1q76ESvchZ7+kGSrgwR8TiY4Jd3QyL20bkGBCa+bzX1Nf
IFBtKTn+oz/epXqlHELFQzwxojcwevRit6Cu9NO3L+BUo9wQzA04WxBn9i3+
c1SbJjBxAgcea4jKUFMAA5oLP8CNwGMu59siIL1euGJqKXs2rfVRwncqWa4t
TcTN+KkrbtPkeH0buOieodI/GOWrYE/cGNa1Gbl7ZoBlrlX9nFqFhCHjAtOF
wonBpOEBeBKcZcluPNERnPa1ISChrWoQcrUSd+3QgYTMNyy6NtNYzAQa1/mY
EWmHXPtt1UO+627ODN/YV7EJ4DCAgCCRxkGhOrQ9DPlD8Go99KUPYvBUZ0zX
PYPRrIlnYuBSliEhJSY14Q6GQynH5F9LNVgEwKrXDKVLosyJfUCVDQA8BI7/
/nKi++4/tMFzm6HgkLBZmb3uqmjzdUxv/5Eq75b0Qtm7QBEicesXhiGYvTnO
vLXwo6+IPNOJntTKSnk+1wTDTP/h2/wDCtKPiZTx/Q545ZlgsdbsLaHNBfL5
eMok4+mq4N0wKNPefIkWK7xKKlqQ8ikMBcueOESU2nb5lp0wCWJiAq+NIqfg
MKvppMVWkQ1w91hA1r/J4P2AJXfghXoA62m22qpI0HuAeLHZjXktkvyOsw5s
6/ysrsLEVo2gn8TagmCX0sfiH2gdjdwM2MubT+yzJ/nD8Uc6NfxtKYw7Bj9y
niqa84cV5BAKBwc/2lF8W+NzNn6ZnhRQi0F6XHbdtbKwsxSmk75/nopBbCKV
N1c6GNn/fhyC/fmCyBVmYld+WCzVrTQbtHYQ8WZizz4cBGXlJZcjlm3aRH7e
cIx9Ju5IJTnzM25lgGzw0a5KG9QBq9LajvfDLkRR6H6DQVpp1C7gYptIvsFt
Xj+C3pYAa1gWSDCor/dsZv8W2WObPxmS3DmR9GrBsgeiD44P+eQOisnEcgRF
TTeSyIlr2N+Dpat6lMtYT9qQt72Ya7TKpi8a0Glk3Jg93i+1Fr5Ab/DDh+yV
evuJoeSZAPTVXexgNGbjyY8GDdvgDWFxlnYQYUff9hTfaeSd6+7L15o1rufC
17J/5YJxt/aNbsHUbwpo/6/1HLUwrUjVjQypCeIHEZT6qD5kA6z7DFtKDw6n
c/BO2AxWBaY3tHShpCKRuwPyos3vtm6U0bqMD5FKM/ix3+OKQ2VZNoDiQky9
N88NFW26KJac2Q7vQD8rvzEDffiJaHv0uYCBomHRwkbbcilA1BPdMDtVOA1o
sCFAmrXvW7EX4YFnSHQHqvvPc2Oy0ALNTmFh5O2NOo4vlkjqnK1uTqFyws5c
vag606mD0cXFznEQSJCYJR9r7+ghAwvzRUs+o3awa/9jdPAvMVQFzTDnHg0l
QflWF3s39FHzrK+FTO+KQni+loSUnoSptmw20EhJqUVLDxKyX7JyLqcrjgGz
hSpMXeWbzu96y5p/1tjl0EoDcqmOodUiQ/IKUHMJWEUqPYmRGLYSATjQfCxx
p3bcSNaxHxnVnvLyw+TCXCT4jiWlkTwwjUNcn5wMpsDQ+8E1Eob7pBctmco7
Jv4PLkP4C9CNIwcO6RtApes0SNRF7wqUxJR1kNRFjGJYIOBM0VUUqhRx1tLN
9h78kysxj6CmBk4lL4Ak9UoKpHsZzKF5+ceICvEq8O5ghADtaZzctyT25biV
47Lb+V4MAKJ8BFth+Dz3V5WbUkNrK/tYk3X52CIaPToQ6PovZVhPfDYN2h5s
bZPgFgh/arDMNYBKW3MONapoU+yGpaZ0/tG5381M5FeRTeiNVYy4mzYwP42R
8jzC4LiJnQaB8ajQFh9evSYTIVClagHzFSxSNnCrwtvkZeaZZsPklagiqkHM
kP9VVuD9cosV1uugd8j+CDE+wOZOl5ZGCBrZ8kK14qRI8I9ft38+HgsR/us0
ksyBCjaHdv+J5QbSD7erBJVeBLJyGik/7TsJfnUlOIAXI3q14lQsGw+izLAt
6VdtQyZ1jd4R0U149Y6wExtiUWYvI/ECveUFdRvshLTVSxupB+0XkWk1w6hN
Br9mMSCzYGfhrKx2LFglyFxtt4VOBmCN4P5QMV0YlI/wU1bju0D/3g9kanB4
0nVYoJfCCG20vcGjqCmIfblOIZ9s4YxyiVOpSMEqe+YyUmvQvVGfBgIiyExW
CS640i/6RQHyOkTk2g0JK+kJ4adV3EIzo3+IVDi7WP/HvTQiuDzo4pbX8OTL
bdfvxhiLE0slPP0pPQt/8Usr4CmXud1Bz/xZUwBx0wRcZ8qphmZ4y6fwkmB0
Vj67XmOaDcUWbZCXKq0QuM51OrzSR/MA7x2NxpzlDuVQYw+BR7oIt3iI106e
8ChlwVdQgYqWVP/N06NAgmU119C57JMxQMDphi6hor9i4fTd/xNR9RXqGcDJ
vGEzgUqh8wEiftvZPfk+INvAfPG+jbQbUg3DX94azdv48WY2fxsRKWvrJ28k
fZkkYptkWGbQaqgCR52yVi9RgtEAO821oZ2kPlVYoQNrjf8V+B6qk7dVuoxZ
BCLHI0qL8ztp0HqUJdrMetgZJUlKkhqAf61f+Smcs2QdCDS3/MEgC0IXbV1n
Dc/j6xIC9WANK2URxQ7ztXueTCxepjd1T7gZjKua4EyX16hbqxYcwqlIn+Nq
om7tkyDlZG/Mjg3OuvXlRbYrzdD/PLRv6nyYVWW6pMZGyIwKOFc5SgTPI4ba
6RHNIZADrtdMf0JXOmPHFT4jPNZ0a7OYIE+ekqAcTIwFISJ5PaRCVVFb3QIa
TGwBFrB4dJ1Yo2q2zM0smtcU8I8UPHGS/WWUwgkflq4Jy3g9tispDt5nL1iY
3oRmy+2cxjGQMos2YeJpiahAq+tXnQSwygDMOpZigmXu5s1Q+c3ICMarUbMu
oQnq76I04Dzu8Xw+dG7y336as7hAHWpwFDhCJ6gY3HlAsaBRE2q4qtkzLPm2
Bnb+PcOaojTBuP8BzN00QNSn+ZetHQBCQapYbiI5DpF+Ap+2nF7nJX1AydZB
2LlVhekiVLeiFt8sRVY4i55Jd2M8UyqAfiU9gloU1BrrtBZDNlEgZGdvnVHH
Z4/8B2RVWK+F6QIpKCi/RpkJIfEwpXgBvo1jiAAw/mEH4ZOVO+aLyNaHHtFF
0Wtt7geU+6t51WlQ1K5BYzFhzEdQr57A23kt1D+48DN6hPQbJI8XdAky2Dya
sQ/h5K8vQTpq6xXORWy1FVrm1seVuDXyh3bJGcGVUuixwPSPfKHEGDLSYbYL
zFWGlE508KeJgeHzfJaPlV+keON/iXYyuWy2CgX+WJbhy/HLjRl5aQUC4KRY
PviciHe/3E+9M2aPfHUhTmHZvcq8SqmHQaL7ZuIa7ZghdotNUZT1KyongRcC
5+RpUQPL/upAVW2SNcsxbwm8ZR0PRNqoLnW+PzINvxBNdZ11QuAYrrXYJLRm
ccPvXQMu2egv6/5IEiQuv8jawv+lUcj9JVtkA2+eeyaFw1kSlqRkAxQZ4PAd
TiaoDSTJQrbQNwFne+ugkme+TMIeZ5Tiy7NgIFusIvbSQbHH3nu5w67PO3y5
PAigROAzEgx13kk7ioilHTfxHX+B2CM85uU7CW5hnSu2aYKYOHs5kxcnyILl
ILUyYIEY1oxEXJNvuKIgucjFp4SOzRrv6i+x8aUyioQYXfwUGygNoKqnFXnV
uUO2GRxJ+oFMOUm6s6VHZTTuPtkv+AJOEWu+zR5I74ff3xa2KKcUtx72Kror
TAF/4cc1g7BQXk9GGSMq77habgtEBuaiGMMKO6Swgl3LfxQ23HF5AxUBV/xV
OCPp8olyvlTkJsfASiovV4TlTyq9chXBCeiF0ZBcqwVtX3Gs/j7V459wO6MY
e4SB2+iGs71Nk1VMK5dn28+fGqi8uyigbtPWIawO/jrGf6UGRJzCcjjx0pt0
b/4/zM2gqVfBvHUX/05s9YpQoUWN5NNx21yvZZhQjxt/e+alC3RhLs2LdriI
oulj0s7n7iPbIY4Jef3Qa6PgkPw6SpvjVAzWKTckY2G6rIJ5BR5NgPc+4Qys
JT072j7wr7idfeHduRx7txpr68lnAejZnbhN0u2/FtXJ4uuJxxi/IC5ZzqHO
sCgHb1QWSM5HqJPWHKrv8fwJSQyQ7WXPFptjVltnZwQZ+VKKx90jLGWYC/rp
zmd90W3j1FHJw+FL+bIz/ifpa2KsN80fU/8j4jhRVLBrWNMyfPMsQxAMhOa7
glzLx0lDqMwZg2iqpBioQBC+oasQXZt2ZXsLA8BmFkro16DuZIsDnsXB5eUa
1jk/rfTly7Tcdl+bdhcnpci/K4c1CRPXPrLsi7ad/g0JZadnsmRJSeYklvbg
DVvTmQTC9qxkfskSHbluyOwZ/xdSHQ9hdiWk4Q4Lw8KQXR6rYsyU7Lr9Q/9Z
N+swMUFXrkcJDFpiXdNl+wSPqWRM+AW9vr1BpTpcFf7mP0wXBVeH6iaujpQ9
7XKHHSn69Tj5FSudQulRxpQybnfP3NU7Y+h7ZmRa6TZyOUe5+y9NfjKm+xhk
pp7P96HL118n/nIMQykKyuwi+CgJstm2VMR1hAPnaD+WR5i2303upo/bNDDy
Jw7qykich/khUAgid4K0nNZ/wxHTaPgRmaMxHeedZiJlrb25dQXm49SQSrY6
fjMZjAQHT4aXa1LrC9ojR6Ep+XWFcvj5JlFB/Z1wS7rk27yIUse4nnnSmjZ7
2q8UdrbUumHKKU9Qm9QsV/v1ZIAWE1O9hQiwBsA+dP8m7WBX9eLtX2xgzo5W
WPwOjakv0zoI54MckrU7f+YuHQ9QsDMMmYppR0nMwH4kf3ny0X0DCtbTGWws
kg5SPv5h0Pi1hhRzV/joyUK2UdgINAydTIjZN0rDvsHYCKkRzP6VW1ATb5ZG
ww6Y2aCIgATIFECmmlbkD0kKvxEJW3bCB5kGz8YmfPIiB9R2MU8K83GotYHJ
6/xMwG0RzrfeV858ydCsG7cmLKFQPzpO3Dtv22M3X6e/fGbkGLPoIx5s8iO8
Czm4ortinj3r6UItt/o4nACYDDTqJEcuTxBog531jTDDq9BfcLutEwvLs3eL
M173CAZ016OjGUAoE/uuD5DYsLEaUQEkW96bw9CzWz1LOUpjbKwGwdju4Bnk
gJ5JSJXFTBKXdp1FSr+N4ojuYt9FUDiRHMB0hyYznTSOzGkOqza9p1zek78K
tltq4Xge40PIA9w3z5tO5yeIk11cAi8Kz3MWhVPUY1aVzh8L2btz7qsjVW/+
tcYnZOeaiNrz5dQ1zD+qf3jfHHo8QMFvVCZuhOTllJ/oNYXiJMkIfUo6/47e
GkKd/rzKNSDu24QcdNKpwHQboYDhoJ9/seyTcR0cI9wPDzG4po9Yj6gEmpel
i/27s79G5AJ/AEDBHheQDlswYqgwidSuGemfuyiYKqcLpFueauwcHniI5ia3
NIa3ow4P3qh+dlwPuOJ36TshoLSez/n36skMXBAtwz6gYhJeFTISlBgNyclT
Ns7qOUp0roD8IP001Wo5CwNgYkQVAlqMCYAGFv3oIF6uh7zGeFKFmAzka3pK
7lAssrEnZ+3imTOEcA+rORj7X3L0xUi1pERiavTfk0Lbz61wfQbJGZpl86th
oMdZd8RiZTJxtAvU0GzjK3RyLOKaj2h8iPf73RpPYdnfmsYRNh+vrLwqxyo9
ZHWPLMvHh+diJ7EC36rs5YXXCLlAr67+AT5/QFvpuJ0fZwzS0Swg5ygRJdZc
yPwkAisxShbB8vbEzBVIx5P7EBrqrzyWj+Xwo3YCn0QeqnvTYUaHAUsm470m
PmXTTySdolV23B5EV+VGlbYL8Gf0dJ/PJxU02VHdI2ImyXyAxfL+LB+/K+/g
zcccOn40KYaiYpjYc7hiuabQLWA2CDlk5LLq0DWpJ+Rr4RBluVGMUAdTeLFw
rGoey4yeBEd5WcRloAYwGTBo4waXD25BEJ0IA961/ZVRDy++NLEB32dZHIpy
atIw/+upjJb6HP1FcMcoY7uh3hRJOO0rF5o/5wEOStaiyXkRaN7fQy1DxiGo
eX92YHCHfGp+gVWfB34OfNobVPY8AFsbTfbXLnSsv2jzti5wdmj2+SG8RW53
+9YS0qmRHMgSJrXP08VkucSyMM8yZsU4qRgarLXfLXxjpPgoolM5smNs0DvX
vT6k5/u00tSSZiTAVUau+lqV4R5npWuXMf9D6F6PBPtZ5nuOZBGZzzIW2uqO
X/of033p3vQghIhoB9n6S0fiA28iPn0YmK1jivfYjWzMUfK1Hzz0lkYCvcQg
Fc1QcjsM1/HesangyezNiIHvl9p2wNRATV8oVfpjFI4Kk5FdRE4GniS9MtrA
jMXnYfjp6U8MVGkChFCLfO5wsgtL7mnacxHJKUUV4btpB4LOC8jg60xmlOtH
Tc9mwIiZfjOG+5jO0SCQtMBW5kjTAFhoKDZ3QYoiGF2TdDwBEA7gPNCzttdT
SmE9as1DIVlrmp2ZhCMsRwESZcaPfeSBxE3bnDizmiqITsyETz8ROPlhnjn0
M6C+Q+Vfs0WIvJBkDz3PVfqrsl1rL+5vto70t6WsY2/3lCK/0LfzspGeIO2W
RVyCwS7b92IA415vTxJ1EnuTVIvMXo3xH4yqo9LiWsFl51lNBCnw05CH/OEQ
7/dZu0cWOmdnKWNc/PPByJpeV/AVIhk+CavIZsBWGt2CopIIdDt6wzCeLZMO
mre1U323Hxf2wZwlxFD07uPBaTxg901ylMW46i/fYLVEo0IJK82sywh5ylOL
RdVoQMryJdckDKs0sbYSfwUc70QoNY2YUHUnI4M6SON9DeR5YMzvOaSDhFfg
flb4RWn+SnjHUxg40F7uFtEg8mh0toN9wx6+tPivIGrpQ56XLqmndS1ffsy6
yIpDLUwEUjebzjF81IcY5rdRS+25YMHAIYyTV0vgYmhaIF/g164kKho6EHWN
LJZkYIsOn50ZVxOYU1vydZb8rPmRz5fChJEOZDLQNvr8/sDqGj6nPKh4ndM/
/Nfe1dkg0YQD8BOnWyEgrvrVRJSjm4dNVUYRZmAV2OfHFgJyB0+7QGQtphjE
g87f6QKRWakQmfhEJ3YZeka7StXUMHLkSpLpjoBYmf82QjlAjBkpttAzGoAN
vcZhdP3CqBBGBJIQsD9tT3quGqw2uEbTGV0CQMBi/35UUXM8OOYPr76nODs8
jgNFxHZ6497l1QFaZbP5Vvw5yr4gZ87GQpojZyCyMSve8BrTKRS+40w9VvGq
pIMMsKtS9yCTi753F2aC7x9Lc1bEimH0WHHjdbsXgjXgSnvssyZTBptYkfu8
eeg8wvq9oQM1YfK4jLe5xllLpN1/ls1kOpmvAavTQc643R2zId8WwmgdhiPO
yP5M6OrmJJ4nCrZzTqdY0DUYL8LmxvE/oDjxuvVb04Y7PuywpVqbHx1XfZ3W
jX8lwVDEXx3LsuMh9lk9X/RbU9HgG3fF2/LtcyY7bmZjenPU4H8vqx1ara6Z
ttKiY8C0tC8yJ/AquHvTegR+dcH0zQbTuq++Bn7MVeRJYDNbEgmV3yMoauk7
lNuMOwdJxIFOuE21o8uPgpLo8mQFkDoTISQhLL/ImsohdA6rf2iRHdXAx1JU
FvjFArl8UOnIT5crB4ObEjZPk25ILF3+TCX1WL4x5D/hvZXviUZqRV1c/XZv
E66k1RKOGcyvGKA3ihyQJyQSIFdLIOTG9AxgPAIQL7gxcFMLMkIDe9WYUb+5
0rJYRaF0kpfRnOM7jsnpYS6o7oFCDDtuQmD3WFmJGu3PW+74BxhBsrGgZLNn
xuVdIZ3CMNzD+ZgUtvxweH94PBeFeO5A6TR0mg+hugQ7RpkU6zb18HzrI8Uy
oWb7nn2h86czYZ6Hs7cAI2BZ9ZUtXRz+g2rjnme+VMoc+2G1n8t5NCp+soX4
etADQJEpaL22WRz5BX0cwh28iGdB6fUvi07xgTiXUJHjgkh0BCu+UZVpMJf2
YvsHP2DgbDeQqtr5EVUbrE/fH6By0JWDldBXLYxdLk/6oWDXk4bTwI0yqWnU
gGgGO9V6GmEFSSnS9jAFi/BGG4H4Q3jIP9mDj8Qg2R9DeKaU7RqhJsB4L9o2
gaJYlzQZC79vv+L7PDnf81NjZaoaMclNat3NisoH4XTwxfdEzcTrtwYt6ukG
dKn1N62xjwazFpfJlsXaQYKuKE/co+xsEptUb007yk130S6WIAfqUAQFVS2N
B3G/kWKT1BNI4W4E3SukGtpe6ZipoBtOqLr1NT6yyCoaFRFhhB1ozfjacEJ2
zhB66YcliQu86QMUtq2Luuz88SYEViy2sYom00nP177ek6H9uKl9G5RATOlF
ZWIS6zpfEIiRxYkGK4wwa9YFTLc543NH+uKgvyZbMthHh0ZnigfacCinpE6U
PewVOX0YsinYkXCFsvc/rSHZvr2Ok5oAgbLZKoJjGXmOTykY/0i8ctHInvou
ztXziJ5NGaLcDhF3iznEWD9u1Wzz9VuqKZTnBF3Vpzm7jbQrzyPM4hWlDWDF
xXohxdUC+NKxh0OGlEYB/L1RsuM7H4yrH4zd5oyu9tIxwo+3Mc9pCCP65L04
HnAK8N2knAa4mRuPnfe4tz9BencNYmLQhM/ndoRWrYAEal4/9cFLxTWODCKU
jzN1Em2cUEqXRyUt3iq6mJVQ9LMPjebcUlBGWZedHCkKCcCGsIqFheNzuWi3
voNJS4R3CpzGW2XWYWUGIml7QxBrxe8E6JtLv9zUnHhk88oLyt4QSZXLFCUC
bdEslg4uX4iJ5btDeigz4bYllBm5O9sGokwoRc8hgnFfotgyeo2TeOg8NRQu
uL4Xm6p2PQ8tC8T6lrlL3KssR7yUeqh+b6ola2yEOSqVPihEU61zh5M5cQqm
LpyQ4hd7TYp3dSB8y3Kp3QGBRmuHQpQqMk4E8FbGcpugGkLu6kbDWhKxoAIF
HSpIRb/Jo+aV0POIl7UGQWYZl/JrU+KkTHTG8iU2T8RWoX1nh4qXQFBgsdJV
OcHkvy8Bpd9u2TyAsP/joAT7JqzhTUmYwq/Ov5DjLjQOevKZdqrrqqcU1Q+R
2gb1vgHaKfxmeEY1bdk7lZtaXiKRcVeXGXozDMmxDL4F1AWnu7/ZnRQug/1Z
Y4puJIl+V/cSO6ewt9zFHo4gPc7ga2eXcMcnA0lonobIE3n+LwTMQD1hnweB
4FhMp+1xEE+R3cwHr8PBdDam6eefgz45PdtkBcGybbfvM9P07j8PgGX14BTG
OyAnUVMdtb2BGF89N2IgSWqR2kon4KKEE1ep65pxLlFZqiWnJ9WI9u3plvLE
SvnNKeTZj9Fz7s6GJspXInOyidBjj23V3c5Nr5KDj397vUSFllpq2ooLZ0V2
CO+Bs7bPdSW2uAkh8N4t4j0UItGOlUWGSDRwbSq3unD4Sk/J/EcDYo8wphw+
jhPlf5c7+pkzssFLUy87WPipTvSRqnDjSKqkzqFMlDBesRrdyctFiw0geZ6E
gs69eyTzYzcQdvfPQTg38gAU4GuImDiqqxHFBANPruTR+vIFA5yokj2M6v+7
S0JestRTTThNVDqtBi7QVXQ0Qc6f62FgFUkVU2NX5Yp3yVwPT4pwSoibXmUQ
D1RgfIS0SU2IJLUQCBjYjk4LJvNWmtxb2skxXlrWvV3+n2MPGEtPuArYiGEy
5Et/nyAvV7aAlWJa/cihVA2vNPYW1sJZ+38fcysnDQsKhcjUJ1fjUWAH+89M
vKcbDO3NRcV1iAxneVx1mx4AoBmKz1EdH5uOWibspGLK7IIWv8oezGi7ppxt
xpZlq49KQUD0rSldS28Pp6HKta+SqScNfsddmFv2TROQqT1FGU/8kkmH4j7U
YqH+0vjobmm8+GxQPt1AKa6c3HbxDH8aZ/ynwZCOzzSIYjnug9LOhEBjkcNs
OqOOaoZyu5vd0CywmZK2W/SOzauAeZHuERQXKoWlq+EZUCYEQnQjSv+is5tz
FWYnajqf8ycXvu6v/BUKf+BysooLlp/grNxTqLsheYbLDl8jrhEwmYidKj4N
zJGB/88XkTUwLt9Ykr50WS9tkFB8P9DWYuUP8IF7Y2BIuYGp3km0asi1cj+t
A9Kmh29beiejopTG9WQVpO9Q12heJRN06sYe1JEPfuzibiCqQ8cuiUrdk4cA
KO3tbknofg2lsYcL2sUziovbuW1fA1H0KjMmK1bXk7atShHAIuacm3SGH8f2
t1xr7o7QXCzmbCk3dGCFXqiNbi4a5ql1aUKSp9Lz/NGIneyfwJTU5sGixe/O
8g1V6tUSY197ciG6HDmVZyJOCxdnS3gEV0f3zzEXBvTpJ6quE14BKseIv/9d
Xb5qcLlzrI6093wOaS/3fobpkcaQW0pSEA3UPlOqotkrAFL8SraN6P54yZzc
eUGS9l9nmZjk/YgaTRmj4U9t7L3yfNV85C6aQGIrqDoDC/23W3VCDvEhtX0B
yTdr8o1C27pRI8NNf9JeDKGsGpfSSmxVRgTtp1hb/zbWqoJCNrTqOY1gLmWy
nTxG82k65mMj0U9JMZARmPBepQO73pVt+PnnxR+CV4oJFQA8PqeABqEpqVUM
ieHDnkw9Igs1iW72KphtLqgnqm9VIq+KyhXKpe9gvyKc61fIvo8NuRS3b1Ls
jfV6nfh7E6C9bZJTt6Z4JOFYzi/owHqLkkAJiikFDFUmvDBAptQRroZlTooD
oNvVyxWY6lx3K3E2MTBEmqVuUtrjedLLDpHWHgom3qPx73klyqeUAaqLmgpN
AOz+/62Uj57leSuTNz7GcMzAc/5TX3E0UwbbclyY7OihkR7GjWju0xlWpHN9
kkur+ereT0em1Z2q2PwCIQZDwK0kmJ6l7l2H3l+7DwzGXCUWlYC2S5iAx3NL
Vq8Gg6hBEeRLxMRknf7KbujTZUPuoqwNPKzfMvAWZwAzUNi0wVN99ShL3NlF
W25Ou7VdSQXQSI/HBx2ihkEULDKo4KsZjz5rZ8pMsPREBqOsP1QPMQ2zjwvj
ZX0HcYCCPIBfrjLV/K7rHAs71uuK2fJZV9Jn/W/+r6GNWihiruxMQpir2jby
5IDTybuuV8csHzsWTuEfTTK9Nao8cU0s4o4DLuL9zAojLr2gsBbEqEgwpN6G
43YBOmHzbTVVuUzO9ulDzB0L1Vf7vzf0KHPbv3VKIR3+zx577g05mDeLxfJp
5Zn9wk/b41qWDYVph/vx3mNgTSRxLnR/ZMcFkATknlhOin0aehoscX4L4ZZl
FG13PzKrMPxDQnhE4h/MczTpPC1IpSGm0szjnCbPeYjvNFgCKbG99FuUe9F6
R1noC3VwGyOFXP/Laq5+DRcl9IeaO9q9/cjFLatp8sGyFRbnxZg73u/qnuj8
m3fA+oCqpVwfriGgYmiPb0Tnnc6VP/UpSPkcrH2XgeWXfd/bBHo84y6o5Ky1
+MBpU5G4kVUQ3W1MNprHPyBhBaJmcEY54pbBV3ssK5Zw0EmHExAQIhRx1xmr
k+oICAs3ShVWVb3dU76lenpj9lB0FernE0TqL4+qmQnJHPbloM1/2dY5EwtA
jcUqFC978671uuUURy5t2srs/0nohbGC3SZm+3vWI6Aos6PSchfaC1pfAUUZ
5kUCYdnu1hM7WT0TFHwW+8KuDbKtDLimHpLx9nF8E1+hRUd06VWhHIhrJF+C
M5td5qyGFQoxwmds3MrOxt3SQ6R/he8DP/DNhpon5pf/pnLUZT7gzFgLDv+T
RAG9pUPcS13jvEQYraqbwX4ySzb/F0AvFvXK/HjOUd4CFXA6ntyV7A/udCFq
hsnAW1UWTBjoVIOSj+Ix7oBSQhjhVtK6I4fWphfVwWs6jMnqJjMdpH6IaObH
snZAkbRWZ8GxyCG79fjP1e2Y6CyK8EjPKN2mcEvjie+7SvHHigUxJp6oPTG6
LLnArGUk7XzjTcLphexmyaqC/bstcFK9ANaXlQDZ0a7aVvnT9q0luxymcKFr
AXE7HEwUIi4fX6uCOde3ub+5Ge/h5ilFNBIflP7yqu2z/Jdm7VlEc2SgPPUt
qIUhsrEX5fGtri6KVfp3P8yxQeZZuQLZpkRbDdwRIv/So7q9BHk4U9MrZRlC
M4HyNgyB0PlXAkhwHM2f8cx2B6qjpmAltHcK4zINTTJPo+0AOb9NhKpK8Sx/
nmT77Vtungvo4jj3Nyv9I4QBZLsg12Gh7f4eN1tcjAZPN+Ad+Sl9bBq8INka
LDE2K/ijgmI8UTaYbk1EluArGAw+lNsUHtv3DczB0DT0X0aoxyChqa4saAuY
XkXtOe/1ahs68FdYW09xfWEbf61Y9orauv2OULlrlxPnrDjVOBQDRgtDv3em
PDvodymLBAFwrxgXE9ngzQsXWCLnvaEZnucKGU6ulQ0EjpcIjB3zClVmKCRt
VWGm//y3C8itBDMr3FvrPLmbghFL/4nB4qCNtzmH4Kco3WQSSpmKNmyzRAf6
CE8gWCq3QXR7GNmOXvNvEHblutVXNWbGwX93rKNMp0gsrgHrnAHtVVQX6NeU
FKCdrDBHnCq4a4a5FVnS1YipiWHX6B0VLDEJ8cxYhA8hPIezmcIGRqH7BVE3
BfAe2ZOVnKnBS2F5w/FBigBEo8CX7ELN0oT73b/iECY1FAeCOyh2m87b3GI3
8ZACUdNtfvy8t4is08N3/q7ngoDA9opG+O9yfhhnrmuWr70VaY3MtyGdoomX
9xs1Uo1J0SxdslZrtAXeZI/JThOAxM8Ss4I221gyk/IStbr2zYFkfs2FyKq0
ZeCWR3K6IP3PNF1K40hvJn5SBPQTnue+HFiGEWFCroEXuKQlxidcMXvA9GGA
RHwW4bgBEB4mw3+ML6rdNEwflI1Juvm08dVEWdvxEGNDtwuCZADQtbrH1+QC
++29LoEmyilsI7EpMfiTJ7C7IIBQCe0oma1Yq59vlOk+TRD1yPq9FyBgGJCX
JX79a6DrDJQu2r8KX9YNNXXEwjxCAYTSiUKGJOcdb/PNa4/ZiT+hDP3OdVOQ
ncKuxy4iq03ktsk4jtGvR7yef8w1xebhv6jM4nsDrYGSOmGy72uVptCkQQ/h
Gv0WgOFJC6okdwa3/KNoy3tGkDFLW1aa+YMX3lfJssDMIkmAqsDoFYSH6yAn
h4tug7ZzuLdIhjAtrNblVCmeykP6ktNptTjQWGRN2F67xLaOyjoQtk2JfSau
55ZXOXu0soJp2J4wT5Kb1IZcDy0VO1GK5PfVziQxC3TthuRsbSa9Tgiugjzq
l2YyDTBnwwWsTVn46xOOKCnXgNkUXEG13s5TDm5fZ/46Vy21U2fEHRGyydZE
vroOQhU1Ksz9MMv+NQo1SeDoW4Ptp8gBbQXumi5yDo62nrQFJQXqn/4DApKO
7U3xjxGHgC4s3FW4p1MTwKf815CY0CVhnmpLAurnC1v80erfkrRJYkRHAd1Y
X6MR4M5yMz1uDw6HUZkvb0/5KLzoM3CN8QxYClDRPr174htIWubSEe7DsiSK
PpFMD3Thyh6CnVSilOeveqMu+W6I7/O+MtQx5amCqWmAEiqJ/D0z6t31o8+j
tIT4ZMx3WbpdZSsKBSH0TXmVfhu7iiRR9tb1ZrYG4xCl3VSeLaRen8Tiak7h
xZVT2UfqZloIImT4m1Dty2ESSLjyDgpKi7QcZCO1tdz+GG7U18Vet5inQtvi
STeRFJ2TPZQtVamB0U+ovVwAHQ3NlNf8L1cNxkJvYoQ9/ENlQegSxbXtL6h0
NX8xD0I9ghUAWPjRAC9yo6bx6cdLSCI0QpBbmU6nvtDLW1FCFYeN7jceBhyG
5Gsjl3adrPniosK5zPUbPCr60qFay/9KtW26qatJ01G6F3r3zUcVitZdaMFv
8x8vMOeNu3ECZnVL1ESqMFRDV6shxOETDQ+XZeK37GOhh+9eKszV04izRUGA
ASPnaGrpeMzMNcOBM2TV+TU42wIICwZDCbT1hOPMGBoqX6TTHfiWbApaAqXz
S4PO+wQFqHCHMaisonI0uqXVzBRUNaDztutjrw/3rYKyVhTXO8JV2ZraSSBE
40wjgRgnsHZfTNK0MLDzkHY2HyMxieIrgIPQAjgTxL6MmTv8JV1TmltzIzy7
P429klFk57+W7AjH9HZk/pskUZIic2W2UJvhFgEjUtBPKy5OT/cXiYlXyl6r
tw80OVFmr5HsFCO5HUai5E52VanS4ZXWvqlDGB2NjZmnC+C0krP7z5Yba8Ut
64rC7KiydHfN/Bx8jSUxMQTbf0MqSZicdVGYxdLTVmyV5KhMZo9IPTyyFXg0
qqUNAy8liPOnmvz6atcKIimUFgSg35+8IWArJRqp0ctVVVLGQ+aoQur3tNUn
xWEKQErQIaHBH3S6JxNb+80C0Iouv0BnYT7U0zJ1ufwxwZo8WQfG0WSexxWE
QqgGSNRfyJdJpcPa2frWrp2APaS7y6O8OvmV6SyCEiiTXRurLFEKg4qYkdiI
X7fx2MKMxZ+aLhy38hvSzpfsUGv2VcH8zlFzkXkaVIezMThRxPDHsQB0PXd+
A2/xJv0NbyLRSMyTngXIljG0n9xp6CwAC3o/hxgM5NRk+K4hTCS5F2EOOv8V
5jskZgcW7SPyufqTB9vkt5vMogsXY5NefaepnSalJsfMXD/qSEWhOu2VawTj
saNsYdowYNnwnTp4R+pb4LZ5bDVzwwaL2fSDQxR5ucHe9YFfT/OwRJ3q6d5H
1R7zrabPBqx/q2+Oj8a3f++QQAPlCV33oYbwOXKmTx5WNNCDjKOZlsnaFFqg
ZBpvMI8poBxdtATeyDuPGpkfXxTPOaaEfoOtiQ9PUv3Q/YmV9T4V4dY+BqN7
VO9XhD5tKS58pzabvCaKvggN06vgddACCvMDqTfwR0u4BkVe93Brb/38xg8/
YjdyINhUMWA5hLJPNXR6rW18jmxq2Lko4bd3w2vChzcRHp6R/XGKYAWEvWgV
//+LGUw/ih2KtImT4oEsCJ/0G47gcBMeeF+RybsEQdT0OIlOvZjzc17DM/Jq
GRjCWV6Au1TnTW+2EU/HjCY4LyzLW/h/PvhCXKeW7MgmjvX/zneyPWi4GKc7
QakwdCiT8A8Mf4x+kghnPO4Uyb8TejmUSdBj23QkJ6cCf8fAdVSTi/iX76cH
qqjAHrCunf3cHXtXuWVRaa/i3I8KQ+DZ7ZZ+eFLhUIiW3aTtxKXiQ9Avq53o
Z3FmspDPaq3D0FZT9aeTKzU6VaKyxGpW94tlB6A/J3T69SGFbD1o6tzLegt3
S2Bjf8gA3ZUw7doUeSmggDrguYcTPQGC13R5yTF/L5T0fyP4Z8zaqoZRQYP3
4olu0gWB9RM3NEbpq+TfRCjB9uwGqxHFfvGVDN1Zvechm/Z5wuku3prcZQTU
nuB24P956sEk29RtiqAwBIFQ/cpzyVB9/NqJn726YZ6FIbwwmowJao7n95ww
yiMfDCIHeGlzYGiMcUPWuKe4bNj4SAT3BiLWhxYMG1IvpX73R3qEPkvyewq6
BlPfygkolerJgkB06P9fMnGXLjL4MvKY7EJYcaMsW9vmXSLlc2ef9/3uvSq3
hq4UsLB+JpljARqJzCOScixYWIKs3SQOYi6vGe8q8gq3vMrYmmKJbyvOAkVk
F+3TiLjwCPFSf+kHKtaSk9iW7CniglCTsYAKykkDzmF7+E9WqvqxBZSlINkF
MkbE0eMYPiCyzk4pI15moxlAVeDyJ86PLhX5raGOHKoqvElblyffFHx0wVnl
Rl85AFpaUBJXPL6c9xOtJhmWeQKHqXYHSXUUzEG1UzONwdgKgHywvuAuf3hC
3VfcnMjbw00RfUuK95Iz1IZvxxuQaKa6vracwoEwC6JS+ZizaveOWYl1R+Zi
mgfpvBs6FJwsLXOhFHzFMb3Vm6OEshjNc0qQQ/a8M4TN8i22Dw6+yRwC2gIG
0zrstM+2jMqgZ6G+QYHEqjzNQxsVbTsaROyGQiJUof4ejw4IGDcbELk1cREi
4ypxAkdxHMMRakQQ5FpwF5IhjurGDTnTUNelIcKOn+i+n0vVg0scfcYGjQWk
E9f0r05yzLyfKtO3FusjBtNZ9gqWaFF8QxNI62d8/TnPVo1i1UlJHuKpaLyG
NraovWTp2TzqPaPkYUqOa1xx2j8zZk/qfEy6rIIEVS6nUfL9+e+VZowIhpef
d0TU14Z2PYUJiRDPkSPmtPdmMD3Bs4yLOuvlNngXmtxFMQH5udzAZUTfdnfx
ximV5EoZxJrbYZ3TVObcdnoC6e4fc5iUrtEXaB0ay6yQYHBjFdmOsybxdt0O
6e9tUchoq7YEM4b+1gOkW4Y/S5ewyhcV3C3FcDg4w5ecwj3YpOede5ddhhCc
lTTrc4Q0QCQo97DecUptmZzU4pUgC3GgVWAZ8SyBW0tJ5/3uPm3kQN875vNW
I+usBIrnWbn5x8E3cCVLgboGaP8ozOT1S6v2U8opu3z+45QRoehilMJVzEO6
qbxFfD+T3knysj7FKEyxSPwxaT0I6N/yF5U8lecAJ+a+W1/x++s+CUAbMXw1
XllPDgPJ5YMwGQnZPApVxy5qhOVsdPERvcUOq1V5cDDF3/CiOy9QogUKSaZr
iVFHWNhBoe8p9PhYhQfdQm14yVd+dDe3ZD9rVQlVSdCjeYCYPUQMQ265fLVr
iZ/molS+1Qc6noP9JPmfTUqVPwe5E8AP34KCjNpWgoy/ueLe7fZp2bvyBNT8
U5pV5jzb/NRXBew7eYUCxzUBnEFIOnyO/9+z2nBO5nOtxwgFbEmZox37LWuk
qQempx3ZkSJ9pYPkfCYfeA48d4VR70Am2ibhJ4E81Kbmk9QSVTIpKuYs5ORi
d07ai6dKqQvP/WKYKIpZkgwQAi94sniCknoPby+XxZzVnaEgOSzluvyrml8/
iVi4jc2GrtPFGyHV5UvQ1Z7rTIa8j9C5b7sA4q4XBQsmTfaUzEVJObV+slxg
EGqF9SmUs0yDtkhvW0CDr1oM9Ktykqmb+Jw9JpB7upxpOnnX4D0TkS4R4eWn
BkI8ofgClXejY7LFRAGXjdx7wFEZwvtT7tUF7mQ/UDLu7kxILBpsWp3CWxLb
ebHS4gBg1G/LTvlT+HPggp3njy6GgZAp3eGnHqjnv5m/cBJUmiWcpa9fmW3t
JAL4sbqcz5AUY0isdRMyDxvgW/IMUsVEbPIQJsObU3suhlKbotyJxROMc4WK
XsE6LTUJPhNy1kGfoPoHIhl/gvx6ll1UbZoWYxfgWIukPYR/gol11HjAELLK
WULoHkqcuRamr+2CPj6+3CoqMyyezQlJRmOa1FwUQXfkGgSpDVT6cIFj+laG
zLXOzBC5lLhSKFeRIWcLYY1vbNx/JFZebDYlYCmWmVqM+DLq+uBauOqVwaaQ
G+ElAzbj5xRz/JJA+D+aIZ7KXIA/sZAJcCO95rkM5Bao5gO4Owy/9ICTNVkf
zqT4Mok9q1BwzYvGz5eKJ8VMhagnepaU1zPyDz2/y+0gdMPsWz1SPoKS1bPN
icbMuAAwigrvQOvBL66lqWrs0fPQSXPLN5u3A/a5HfUeW5rMfHTBsSQ1OqEY
mlSLPcVJoWwrYKuI18F1UOgQzbE/YfSaN+oduyP5etqm2BDwUsKExKwtnrnv
/RHBmt7At/yT+TfIWu4S/0f322mJK6BT67y8iUbIr0ozxtCzUFa9YXUd0kRz
trKzSP74uAUhLpdx9Npz1AxzGt5DYGQPgRNuyIXZnGt6y1xgSNrqMF2JT4nH
qsAOIBye8eWiBaHWGyYFPrevO9UINu4qBRrHA7McFLrtZfP5ZlQnyGXRbraQ
bz4X2xifGxRqCvcpGsekoLWi2mvwFWX5D2bESM1Mk9OdPp07BR5GzY26JEXL
LNxkt9LqzlSvFguOI4TxEwusdZcNp1YuoXROQfB+sj5L8H6iyNQjkTZN3wI1
xeIzOA3fWhSeAHV/aMYrit0n41+tlfBYzCQgHUit+4p6+aGFUu0/D9mJl1JF
N60iSZuuK3Ef0byXG1LwTkB9F//eWM2DAvV/1hb6i2lewsARt8ObsYXiHrQU
uGYgUAImSZfg+YH71iwcMWsPTbKvTP2y588Qg0c7JXYiVYw5B7+4HegqBviA
Rm7/IVHHEuq+KnJlTNxEobs8DI1skHjywLl6L4IeNDuk0giwkKQg14xpkbb2
LTrzE6cbyCnSYq/WIRR29h/Yhx8yiSG21JVID5MbMuAydZNphR4u+O6rST61
ec2WwMGC4eteegV1UvQAWJyS0iIXr0gYd0jsTA5r6a/9i1ImV7/KlbEQ5x7R
blnS2Fo1lccUos5G1bI0jFR0yY15ayXeZ0V8j2f/p+zCGiRqyKFZzyGAwkb7
45RvxRt9y9MWxu8jCby1QacDbh14pvjFA7B3n8qhdQ2/5+LgoWiBw2rJG2+H
vh56uJ0AKZLAoxltMNeqGql4M3YgUeGLaUMWUvTErj3VNTd82/Vg2Phtbef0
SB8xgD8fyKs801m6GsVzrhO3tDrtH4OE5GA1zTgZLll/dINf+cP6XMDKwBZX
pU8aggwXKOhehj0v9CIzz+2JAXrcXPzlqMucG3wl5DWTFDGbxhrL+hUwOKHt
hjQkpEqyZYzKjCnp83yyJQMEd+TsJ2QfxZBJKO6tGPaNIF5S7bIAgqEwCTXX
XTRI/U7mFtJT4vqRtyNsbYSgXuA+LI/JB9rW0WCbEDwKdr0/vcA6tvexZJQg
Ecwi7UOIUeHqSNFsrILryWRW9ciQXDTaqMTxsval57B8hNANWjYdLrOlyhbe
67np+q7gsgV1d8VTAlF5JCZSXCTz7jL2jnuguJHr4AB4uB2zqch9AfIHN0JC
uDLBCWjPzxFNCkPUc9gfYGV9rxFk4rCDzvoHgkAJa6Vr2pfHvxK+EJ3hBQrd
XL4wyc/rZPzth6z04hpLiedUJt4tnNTwsP9VtHLfbF8nRu1WBD2mjXKymngS
g8/saeKQqTo2A8as5WYTApOGPaStvPaexo0x8ZjQo85foKuGBN9S/PXSqq2Z
hBeyZKXcGwflI75Ifff5mIuDKEpnFFN6Y+/pdmz/It1ZVqb1F1vLXmjHYysi
VfDC/Ui0vQ4cUiJMOLRtGNrUc5KnCjUZ4kMqRP5BSWEQPiaORGoFGeMj5Qlt
QM1/MSLzV28fLVps6JXTX3vZ8Vr48tsHmqoteDaeoHQ3XIBUKqQwJLB15ya/
YsKn+XEgh1K+PJMAsJQq0gFPceKFRNnExUYfgOfHXWcpsjmBYDuxGlWZ3fZ7
46nRyd70lSsJCAOXmrlvgwAyFgrEla9JuJ0ysUxf3cqM/q1RYAF8GREzenxr
MAG0vos0LB6ocqjzvqCvf4gRfo45XWcPhWi5cRH274fF+WMb3fmqSuQNY6gK
FvpZVwyh34zG1OrvgarutGFy3AhoYecJbQb+odQzp+4UlrEelHtdwUssVAm2
VEH6WqZ8LxxXils9EYkm1mCczRUUi57B+vcnlCiaswQcQPgHMJJ6pNJRmsLz
HG4Ss6ZG/ZHP1+it05XElq5qb/cWdRrTLtymyRxZQK5BzQ/dXH7qWrvIN4fb
duT8F+9J8NiUK+s6GaLS7SLotB2+l9glfljJHqKw5UMYiNP/PmnCJI2xkwMk
JNYHe/40hlhdI420Wy+T1nt+TVxgLRUm9GnjuphUK+0fWM+5PuoKUadEJps5
M5keBBY163YEuzj1u206ZEL5bIEG572H/ipVfYSjbJWZf5AwND83wM6DIbPw
AwGu/utb9U81Hf1S3bJEpnIcHuGKuCGiYomnBfqkCvT6KIu1Wzw09tB2VfTs
ovT+3zvh7wRFi/o+ExpZWaLDQuKkFvyi2oUc8pZxE+1FBn8vpubQWv9MY8px
39VorU+tGjpIUdhL3zSOUnfoJfvXEs84gBOI8qSlSOhGvFgA6brNcSKHDxx+
TLcG4LdOZByTaF7Q9PcJ2DYNq7sLWBoICPJFvg/SVp6vqGaESH3121L9Iw4b
S3C6K7bZOqJmTzWSySAmDBIslfXxQ1IEanm5vzMLON3qnkMXqzdhlMFXhICf
EF8lk2uHRGQWu6/30pcRxKLyIp/jj1ZKMj5mv7RG+hhxr1YBM40/WZsOulyV
n1OrFM6wn2IEFSmIDyjbnXckqXl4r900geq4QPGKKMAmrEzj5luFSvESVwK8
7RrH0gB8OId05qHATycAahVUQSBC5FNJz/cdaS6BvSkWktuXfqSfA/6xXbC1
5kZukmE36YcnMLk3JBLG7uaaRDrvoBiZXzW6R9rKHLgfeqKEazBsA6NOg1NT
NwcVSvy7zWccTJrFdI7YvAuyV2dgGEOHHyfbHS6KHz/qwNQbJMtUfmJAXS6M
yIaiAkBy+Ibz24DUe1ziiYXn+UD+BTwaPSxUF3qZoSo0/9tKuwTMgF1P1ngC
ASFbOEJBE5GF+YorDnJWA2m90OuONjP0SF4D2szoHl5WtZCUuVN+CKERRLNX
+WrWnEDj7x9Yc6QRvjoKxcyR6jCTCj91HXPtAB0qSvNg0/Tvb5ZZi27fwUnU
/pMJlxgMKOj2n2cE7MRcz6MOyr5X+/Ts4M9hGGaYZ2L/BWZN/uZnoMIGVn4C
IbxPzR2HNq+43akP57HDAsc5xisNW1htQJlFA87CB3l5MhNusQeNjqDYYrUP
p5bzp6pwMEdTufCaDJDoiaQW8SP04l+kpzTXB1O7wdNkZAn4bfxkqRm69CBT
lOjURKoB7V2DGdoAxNl9aGLtqFTElIFYTXycvfIVjiapSbdFeG0P01zZtoc4
PUbHzm2aRsK8VlKzYAufhcbroArqY1LoEhft0+p+GyaPkoKPf1MQEKQUV78K
sG4zmPRtA9Ucr8VfQsa+w9qeSRK8H1gOKOeAkVbl4EpkmY8zo6317bhkvpCo
P8Z2SkOKiEsmQyPtc/1bNok0XBFoDu9Dly0zzBSs11CeOHFyhdBUq4VSl6bm
6CunwizBkEBxWBVvj1erFn3rd4n/mCF9ducD63GyJDzoJZdfw20D6iAYgIyC
2pEqWSNT5KwcO5v8KgJYx0flfexvsehrKLQNT6LHFF8HJ3AEKfMwFYmKiBwX
HjBoM0nB0wV5u/DAOnVRlH0oQ66TyzxqEjCfS67y1lpfcmvJd0CO8sGkz4M7
MnMjsApSp9OUpXrVid0s3KjXm6Br9OzaJtWX1dpYO/rc5LMaznAzLcL/jOP+
2oH4WjMemFcEUxA7ZNEwpDrz6u46nwJlWI0w22H3L4BIsO6rHf/jty43GbCL
wIqhKlbFC6h10k1BaMAZOAJdG60OrBggphnoiV8WxocS023S3LvSlX6AJbbB
FO0ZTkhAUCZhRsqNFQ/y+Qanmz/3WGCQeq7cG8XeEdHw80rYRMd9CzSldMiy
uUynNF5pIqcxHou6ahTUnEldxQj+Vd/O35qGR0ZYjL5dBWDKvDlD9F5H579+
b9A1mTM5s07hfMZVkOFc71jfZWVHHzLOx0FbeUryrvEfIFTnLm4mFtc7OT6m
mkj9k8pGIww4oFj/x6tlAeiEpeJGW5wIvKE6t+0BfXpMriUg/IxkGZKDw3AM
pvOqitinVyolOp4hVwMZn+FUle+WqUqBNA+3nbHjr6pVdkK8V3lrSkqFiWj5
Jd+dj77XvRfUr/jAW7NZtT2ryt9gP534NGLsJDzBoGU/ak94Rami+BZOunUQ
5EzXo+jU6XZ/t/2U5S2RkRNFVDER9qvLq+McURk+5wM0GQosyI4SAD/cNw8j
dNSbQy2HVidGtHSKprVQY6Ae6M9pObZX4EdrSC2YvghZJkpqIGJmpdARe7tV
fgCraIcfi5bq5kvjbjTN/5R4eVNdWwD3nf74mcd8wwyC27TwIjPIVO6vaxXR
9n4crOsosI6ZzlTcNJmMjIoaZyd8JxdMsMQtn2iB8wucql50x/RQDiMB8jKj
hDldMWTTkag2yGYj86c3RAex73W+4v4U2Qa3dIJeOYFJy9gb4/uViul9PhyC
3Nd0HokCRRBwz1LV9DSpDIJ7YcCgYzveJNSCclt9Q6XWKWZ79/VoOZ8+nxzA
fb0mSP7WmJAXFL0YqlbQOLH/YMxRvqEO6lK21EsFhzONQYKkMEP6y94YHjTb
qphEB7k38rBERUVQkMZcr9gnwPTa+UYT5YvJLuFZyOVVi4NdlCytdxAs+rDk
/q5IOOl/ErnfStBPmQ3Ls3CCLLxG5247vOqbWZaG51OhFPNj70cyMLV8Vj0L
mN2nzVK+mq5dcT/MaT8iK7XGDl8TRllPk0JWGQYNaXuS99/d5CE19lpjPBnz
449gPFnXpA6djjY+j/59DjeLB2B8fohT4IiMaFwKSvpUyMXWstmmYxF0X+LF
mpIrjHeAuGGn5md+NnrSg3M0PXqEsdQWYdBzk2CD9cehW3YToF40ZQt1FXEA
n9eYxbprkugtfHdlzdzQqqUgT4G/k8ymZ5WplzFOJI4jNMDEiPeChsDfR9jS
Laou1cKydR5skBXhCNegSVpRMqD4BhFzBA0Tnh20K7Zm9L2UEMoacO+lc0o0
a8izP1hY5rgRFrFeeso3X+d/MP94zM3MCZl2zKzlOBSspDtVdU+qEY0I8K7j
PULO/RDoWRfmMkjSTj0ILtSdH155ssIkxRhvg8B3h6eDWWvoNsK/TwCimXNL
YTNIwdmy4ztAWI0symdTNi9t67M4vjxrXkQhaE818i3J6rMmiEbd9OKVW1bK
lXNB7/DgtKA54HFvdihPwUUXRxEd+0QK9nNWSqr1GG1gGm9s76JBvP9DCMlO
byLGguU0uiuaR1aImVQQm+/ZhZaCKPeJSZB00zVD5+HwvkoDpEYUegzb36+p
ITKQ1yOoX0QrpGKSZlT+x8nDTcFx7sj0Nj4GVhKtRn2XnatJsUIgroIveRJn
lXd4t2Mek14iZVhnCJzO/yYudM9paTGHoq/sXxI3Npgy15HW4J+CkQOkrHND
ANezU0PGeouAzyiVZvhervmBoZYaGcQ0fse4IO1TYRFj1hXWVW7UewY+/7ww
EMujBykhuwcrEQ7kR4Xp7akJ8EKjgh8HbaTiRUIVo8wBEG+eFiQ5VPE5KD77
X5dnamt8Gds0Fe/8AmJ1vHx646t1SwBGKYjOzxW7nIhSxql+pks/8SAQKNVO
z1UWiGXiR0AL9ATaED6ySqa/BB/uoDe/zmxATlk6UMBRwSTNpCjbnHopz0SJ
rzs8hLazqcj1swnutZu7k+aaOr4ZM64oJWhGKMhTu4/rUX96zEGaypB3NB4Z
b9ziU2PYwewXUc+zB8MwzNnH3TNix9eRdHj1+OqSswJmHTP6O/M9bGBQD84u
wbew8vu3C3FgCsQD8FeUSkI6HTdy2IluAZe2OpAd76Sc1ZWAAg39Jex+Lp8z
IJGmtWoHNj74Lfr5/+WK/bQax9RgZ8UsFycxNhVfQiPCkX7/HkfWictDyibl
86rj7qhZB3F8MpFzI3wXPk/G5ebZtLfnKaRBe9LOJanVcP//cYuYhWICDsMK
UWTwvWptxogoXRCNQh7W0EPEmsyNjhymVTiAvXxD5HedS6Gb94C/XYybTA8L
aa0sbVr+O8VVpO5coQ6VZG9frIRGqUNPmTCz7H3q1XViXYTSIPam4KDKaBPJ
XHDZhkF8TiR5HpKCET/F7ea0FBbyM+HhctUVhVPjt9Pz3pxNuaHDZjm2rIFf
zNvrR3DLOl7KaL1n6+LTgWTgXTvFA9lJOpB7gY5YIR7uDTeqGM5hyy33c83l
jKID0moAxVEKdZ2hAqcTGoPyplplrqQsktnUBq9uf6z8FJ01ojozd8MuGIz5
D/DXihKaB2alwJAtIcvXNnE++BLJmPMC/HHSwCJjdNZKsmd28cUtpdw9zJIT
NUgBr7xkR8DGiMKaX4Ubzu7r/bRaGaIS034RhAQV+7zeY5GW4f7MksRTMtmF
w7xfPuF9Fg/Y1P0JY9MwRefAloGYE5FsEXOXuoE7bOB1PRIiy3cI1wDF6wrv
Jnsj9oH/x2yay/A0mdqZbhvJV9FU7MOEgFVA3ORGyRg13UmS5bz1CEpXo1Vs
DGAbQK0iFqCbsCfftAGmXpWIYAGVq+HtF34PnitMeviI0fjbx4QKv3cF5CUj
3MTyz8DVkt38Ei4cFNn2vzvwtmFiSkPEGyAa4BtX6/JubMSTfE6C8p3AROVK
m7gvGTNtSI/5ZUuQE2jndOH05JgZXSTTSxx77EklDtPnaq81snOuJztKQtEz
y+A7kHvv60BWy7Ip6YP7r9opgxvsTd3+gRElJwu8202lGcVEU6H1u6T5+i2R
z4dVA5sX36dri5j2vdXzn2Gw67fB3pitbG3lKOIyihBXoQJVLHRru0s+QBv0
AGkqPnHLtqhKeY1gbuuMPz6/mV4TLDdI+Mja5s/7C33GbzF8hHo4dPCL37EH
6xHUckoluVWtyUcTBBFjgsT18oIwDK7K1T1Qu4gGvcfDkfTHQkTqlsRgAos9
XhHURhBeizbaf49uV5Sz+sAbiKkvo7XtuOTMgy2ibRcozGuY13D7+bAXiF8y
oUIdGYFH6MFD4/vC4pKKxTH6gTizex0PFnJZZS0it4ciE9vyjnyL/6gj3Ied
M92hAlogzDepEfZ/ACKjGhiJ9rSp6d7Cc1rWu2a6pYXD5BRdV9Z3hdSKzSPM
3TnS0qAhI7CAcX3C1j6KEzECuEjaxSF4NpHvY+kb1DYGDyVohKvTioPL8zuI
0gTdOc1XqQ28uUkq8vibgMSpvLgMPlg74oLih/Tktf1L5x4VikbHk5It4fsK
hLfd2iCxIIyChw2rbI6YZZrL05HHsH2S7LBQjG+VP2UsunDEftXTLewq80+K
6+JvfNd3kIrl+hIdXpql0y+36mxsh5Ee9uBdGhYrN4o7ahmuuLf1qVByMVI3
P6rgiOLrDbDUUm2mhNkv7rmMHFLFe0v8M02MG8U6Jnsa0V+zuW0UrKWqDK05
ZUI4oRhAG066M+pWzVOUWYymoguAogUNlA3RXUGBrAlnLUnZ2bhGTNZ1mT6s
iq3jfi9Omvwt9njS0qBJZmZaZWjJP1qm1hXwT/yEWC4HdGTPSrLUegaihbTG
Irqi3JFlbvSA+/jH++X8jMgUE5P393sG2guRiwioQOdsEU8FTsa0gRxIFrKX
08QdobIzBskzQT/gstpZ3JCe00JCKvk8kN/lzpPiFSsx3Mem4AooqCZA+gQp
Sp5K3t5euhSlla8PwTl2adU2r8qLyBTcmelLsjR815nEKuiLxsMjLoBnNll3
dH0K6MB/B4BzQ0wGp3lwTjlMa8uKxTXjOWa1YQiTsWIPVHVx7B5E4VjmQ+Al
CGi3K/H3Sp/Kn+KR6eBl3zTsmf0JSKaimCyi2O4FG5c0pVocedhQrUzBShNv
cpyKptPCH+UIxA7hLcocRINGdOXi2qvcZbVBzDnKaHtSZ4KQJgyvUGRtOwxU
kYtIxJyQ51CPoHNV50wC55GJxqSFJyYT6lANbJprjhJkbczBfwvjHF8kjOLp
/lUJh1AdZBeG96w9jRI5C/IkY4PjLB4AIZkHgfhCNLR1fHzf+bnCc8cn9XME
QkC3eGXuce03iuax3VjscaLdpw/NKI9lCtFOYvvsp/MKBgqTA5H9R/RdraZ4
2TUliD3ER7i4rpPX2WWtjCo/zL/iJOvdxRWJ8BmB6zspM/INnAV4hbUbZ3dN
/t4QWsLWhAEdXd7/ORWy6dKTH4AtD7FqD8tHxk+Ge19Y7STeTgYwrbIigzdv
2cGaB5LLIIFUZVsiXxM3zrTMCNm58riNjP1YA9S7vvd6xMDT4leiTbk/ukYK
A6Sj3zwnfh6fXC0uPFfeL/jRdmKA5/Po6Abxqv0NEueJ+2J1RwxyM3CbPesu
ii3VL/tDcKbsVLo6fT3vwRgCaKkQdOEm6eFzILy3OU0o+vbBmT8qgBIxBvxG
1yOEzlcNqJAIAZQFrEAFtdXSItm82x/M4x0t5OtfAyLJ2bg/oy+ZMvuY7pUk
1deD04mvvDbSKuhqV+4kfFLsOvGS+Sg1KdYMKrWs16P0LxR9sp2KKqArlnWF
7I9EOYbKSYMbFxbkG91CtgdN2kTEROPFLyGB/Xz81/GLQaxwjpc1T6GA1nhR
+Kn/yYkqGrGMkEYhiWk8GJs2fK9YZV9HxEtHt2nQY+5HwqiC9Jd5tpjFiUBJ
0Wss/fvqlIZzRXmqF4Cn1JyWiL/nmimn0QvIvlzSxyYgTa764HIrD5E+endS
5pkKXHljDO2rhBtbx0DW7fxik4Bifd3bd+qCkKb9yylCpeqo2oqUc4MMy8LP
12Plagdnq0n1Bsvl9xFO8EVBZ7KCVGwDthGINUOGli/9P2l35Ft0UrTGfEgE
wbtQ7SAYef83TtahsCy4C1Jio8Mn5ipQX4VYzvter1RlZWijYSEuorHP6w8j
7LQTSv+HSAttY7jhwDLWcipHRsI7IM/dCLyLopzh34Q7EoAEhf47KsGFTXAe
o22e4K6EL96r/b2/bkaMB0kyhYXUqegdpp/HxE2gNr9Knt+Z+ET366m9uq0m
Ztv0JgtU5j9ShSe0Dr3CaW7h3eveZX5PXq21XiXmuSQqVqSr5oAvI6jOQSBQ
4jdnGVS68Y8yzjz5yRW1206mKmauoYZ5vOFPgoY/Jr1m6uh2EfsfqaFobNCl
FmBGnfmpGlw46cyTok477P/c6kho0JxaQEPBdomR722qQGT9GEZ/ZD3lmDzZ
BlJe+JssfppUBObxMEpVWH3ULhpij5WCWQGmufqYLR6tivzjBdQvRRpsUOfn
XVkBkk4zj7kuhrvCKM6bTFLPaCRAGkG7TwoWRKopS3u8nw6/R13v+Ipm/ZvN
9IamTMtkE8zX5Qt8v7Ejk3/OUjNqz8A48ohdEsYzmguQD1uF9zYO6lAMVXnO
mIGaxi93fbP4GLY4k2MnLTUW/DYH8hzH94rTanTNQAlvQMc8ntvqAFos/Y5M
ypK9hW1vikF8lvmquvlVhufZX6mwwlm9dTsxIbnCNK053OQEEZUMeaVn5H3v
D5RY/3esvyFEksRP1UX3NpdYHIZGnROBAEa5HPOLlhJbxu8Ax2+HsexBWbQ5
ypLT5DMHZfb6fnGGMoweSGIQWXKkbHcqpRssCvOgCLqYsTSHwdd2HsYrUxb3
8+j5h2g2G1yeW0coU5UY+OqS+MRDj0EzmU00RKryt1KuXsODks4jbqo/k3ik
LtHTk3zQSW8ImwQTqzwDW1Peapsa0pkZSO/CFiNq9zux7GKghuA/lubwprwn
odZrXwHMth2VS5ZBjwaUkVJZI3bFwB1ipa2tEvBM0/uIfT0n/h01Zx0Yd/Fe
Xn0XlClvvY9diRCOtDFwZcOljCLL4/MA+o++0ThcPytGhmYeBsneB/41epdN
3AY6IFJMVqTSCF6zG+USf2V3lxABp0rc4LtsyytOjBkr9OJ79mfAr2HJuL17
7GeGsXz5/Q91S/j814w7n4vZhQxF34Sp3Fmgx/zGMO8IL/Vi619lFL/AMpQo
TNfII8sljy+xyhpK4kNajy0tIOhs5Cuozk1FjsuudWEmc40QNhgcomQoYkvJ
J2a7GX1JoZh9RcozkNctSaVZPhm+NpcDvyYvNETlJU+dt1JLEVT3U71ZvcGq
1IYo09sF8xXdjuU+jafMHkqbskoMaIbfGmgHHwVzcNG/v4BqfN6jJCSWLGh5
5c41aTTkzXDYhN1TsY7SLWeknL1QmWvRGjlb5wOzmRHQZhfMuTujKdiS00NK
AgJbAjOdkB3NbQCyZ3a35bXLaPfg4p3XPVzpFHK6KiFNZpssFWTomuSFL8/1
ZnERMFLq3C6r4/6IJJQC6WvGpAl2/+jrecIUHoakkON5Bm/dBnykej05zj+o
ZxficWSXwe6F/b+zLnKaFeCSYG1Hc2CYV98vAmF/kCuoC9eXUfNlyjMPGBrt
iWqp7DSXY0tEwlrinLeSPXd3n0IkDrWh1VpWN92xrhvfAdX9rk4CJhrXDB2t
5BhQZKIfZVlYFl/zRGRNWirTz/pyf/PwSw2YgoutbqHgqBb+28EY9o0n+fy4
NLDgB/Zvh598W8acLSCcRGGD7XsRS0RiXpsoXn78xqgARFRuE3vHBWMXEUKG
N1I/Fpx4yQcPB4bsRhlre+s9+Tb49lFMIIgCUqI7+2ZjFWR65Ycr86S/778W
uoGZ3nEk6993MTdAvT/Xwt8R89wDGzNtCpuMySqpB3H314OrcG55sD1kk9uR
kslZySRtFWOFs2lGwkfZ5hdoyYdpTPx12lykEcgQpBSx8pnA3WZGvOmDCwyP
rDQUh0syoQp4zSmBtNDX6t4DZwMKe6HKr4mCNRbxvTPP+pWpjqzEjX9I7u3H
Hz8IynHdW/8GjltyZPBlSWX1ijFgERzuJfj9WcCxQNb4nZxaaB2IacGwUD+G
Uq2iyYXDyx7uFJbpbLKpW2Qaw3Z+wTyhqIlRFMS2LzOayfiEDi5xV+055HCt
OSmQyNhQ25W7r1ZxVExE15YrL5PYlY+MKTthTkUy30BRyoM19MJ/7F3pgr6/
RAM8AOIrnQoEE1qyOdCUNQAHkwGwu8YjRFNW6F54Y2DrrxlIf/wj72abQieH
vJFD+5UlMXqjLop1Xx/IHQVFOnP/B4ZnMLxq/aWr+yY/B6YYK+yPaz3MG/q6
BDIEVy6MkqVovGpNKnCguE4kjZaiKZfoMNKwEqX8RTzx+qiBX/zCpFEt24MU
j98URkT5zF8/YyWLCfe5fBuzdgRX19RXh2lLYCrWPx5njXcSDlmj3WeKp0eH
X8KoZOS4gVcke7skRqzHZ+cj13aPYROxKT+So1VsQA8cYDx93IuCZGP9R9Zb
WEYO6jRAqP17cEeqyD/Oghtdf20g7vESA0akhyh0598bNZi+Q7Rw4Sr+D8jL
dh29x+icCTqv3HATChcKa7xHA5VMH1P6pHCDwzDKk25F6c0xwesxqiQ63xZT
qV9gYLGQReBne2ukbIRnSCAVUcRbU65mNgOt3idYEKvE1akWOND55zz1YvRR
TW+t5PQbOqfQIgUVhMQLbwelfqHQHB9DMKL390CIj6SMbp/vypAAdIP8J3Om
Dze8/2qixYaESGtwPkVskLmdbV8Quu/OsiEuCcqQAc5mwXC7otUsSNCp7NxV
qf86qBSgoU7QT4PxWoIcHHD2+2EGeB0FfYH8c1e6GlVH78rweALL8CeUAd3m
9/ytsbxiTfOLNxM6S+WQIDDD8FYqa+F+oGRfGd/eJQjTNAp3RcLxISobDdBH
4D8b1xxK6cVn1e9eERkUhKlqVUfJolyjoElU/2lo6ivFwtW7ciUWhoufK2TQ
PE3I8FMOJOL+P/RsKzZt9r9EIw1z+g+nfyVCRR8sdCvE50+xnUQF7u4SwZCc
8rWYJaP20RKm3EwYYNWYF8Q3b02HdTfh0imqpZzADG9JFB/ZKLdMnMkiUfzi
mocRSlaICIWqeMwh9JGi9PwP3e6nKtpUheI5LcxKB/dQ88NAqQiurv6aAnQC
ENuWY4cMuV1pDsokvDkwlNK5cHUn/JkHIBkdQJlUlldg+ymIxyy/zDYY1YR9
NYjkcVnpKFTHrzw0cyrZ0CqAXcS3Yz5xGHFLRXGn7MvtGhWjqnKp3j2080CD
TtgmFrtvU8FcTov0PHgdfVaGkwOyAt14QISHFnlz/c++T7TatHE66wJSIkbk
8HkGj53AbfGBTl1x/ZdUd2kh4rXSSPwLz6+K+bJa4XMbl17nzd0H4GLMKB/m
jOwEzgknp/Xyczph2bZPFjaZ1GvOGNTC8xBkdD6dJYrupfgPbo3tLFAO4dBm
g50haNYMIwFWxkKBA1h7txfyuhdtMJeWiBoFfMfh4VIJVTV80kogDe8PyLCo
O3PlZoIEo9U3OI7EQ2k2Vz2xV2P+Xt7vKw12i7wmGjASJiovDb9C6GQf9udp
FVAHjL249euJII2Wt1OeDbKCdnROkq1fSG9URImkQ1pk5lna5vRTFL4ow7lF
mcaqtlIYA4JMnbmteBrmDB87x8guCs30y8Xrmw8p7nc2D42UZ0Z40Qy4NzcT
2BzKZaST46Cp5QRf8yeocN4qsDm4WsZeT87jW7icRjPjNiY4U2KF4YGIe8Ae
cDCZs5ZRMoyLlbSWLb+Lv7jcfnP583h59P3AX/7oQGkhgnqMgGxdJ/WVTpzu
o8pjhp9hpiFdbFzFeBbhfjsrYZLnghxHQRq1Tz/j6oDLbHUEagYoPzqAkX7Q
xwwk6SJJ5+2hrkd4o8dknVaBTv49lih5pEc47K//afLweTTDbZ6WV7QUvUag
MEUzvRSuIp+091ZqfwZX+msdc1OcS7et6bpGixRN4mTtSFJJwkAQLtbc/EzF
Rm+yxVv2NL9ckgrwrzvBOhyNYD0X/we6Ckcr4X3crlXTuR1W1mt1wk+LBpAa
siCgwNn+v40CROZ/1Bsb9w98FVJnTLaS7rmh58PJ4sXdnun7W+iJllviNw6c
jVA8GfCH62aRGhtzSiEcg5CokcewSj0OTQcGeNqLvWFcaEfU3Hp+IUGXU/7c
XaqSHKgEbEdN4uMnD1NF0alEueD9Q2R4V0iB4SPZaumVhuKHpRFqZxfyR6J+
YpdqkDR3fq11RHUMoheXH4o5iKtIM7EpdWFhKryw0L1rl6lW5zTX5BY7sNs/
fwEZwxlvGkYWnBL3mwgS//be/ejxqLCIeN7H40xG3ZZdBx4vth+T1MUVJrvB
K5aDAmWHDmEVRiYl9R7U1vvEYJazDrwKgxx0a3C0/jul9FfhW/GSbULfxTga
btjQ2pIrYYGRxA8WUzowq3PD1FmUes6zBDkgAhBbacEydwykdGhisLurtjf4
PprgQoirtE49UNaHDIiN6zCQaQgMo00yDZbu8NjI5MoE6kJPjx1d3gBYAwX4
+RfdTRCicFICLmZwHoIXbRYGnYbUn+YIAHIXGhOyxOrFfUjAkocx3roz+upH
q/JYQvW/PyTpEVJCawJuw5eR5kz+ijW0nEDEK6RDP1PCeReaRFurhLOJfn6t
4iQxyOzmxC5b/qVNquBaWHzks4Y/GqXKwmowadkinB5q3EMPgeY7kzmkogU5
KXir7CAZWq+Vt/CB6ympshjiBrAQg3hgZFhZRivlYDlKvRlu/5YJp1VqgdJm
Qnve5mERsFd0HsVH0RFZnvSs9tTF+WjEepCSqyq16BcTWbAIvVcMN3xLqZDH
e6dHGPcMp9PveRMTrLI89vGDDouOIR6i7k1HfkF3P0EzyeNWZTnKyaURr/Ol
C5eEBiWGRR6ZcRQOORwvWGMA2RrfpbSer37y4BxBbeDr+vnHLNbkvUTO+CMP
boKpeL1/Gk65xd3fecqNkIUv5if2z0Ek524RqmaxMs11WYQEsoH/rW2MmTMV
UuMLPlVkVRKHqY4cgGC1KDSVEHNeka0D53M2P8qm1MX1QudbZNP3ycJwxP0U
uqFl24FXeZa0/dpqRrqBblf/CPsGbINo8eYQwpmCCytYwj75wzXZ7xA3jiBl
ozJK4J/qQAXv1XT7nxzM/qHbuq9WBwx1AYLEopchuG04SHr98ylrMxIDmc2W
LvAOQSivIuRI8Ps7vc8JltynL6MzgwmeKE/hegL65xov41iMtuXveHPu9Uzx
WDapYXrG1g+UwVALCwhW4jawEQdkCqDMGK4Qs2VnmbjfiF9/YBL8JPwzJWoJ
rqK+ainetIqI3Zd1ZGHT1bXEtc8biZ5vdrlK3xlVHyJ3cTisVgeOgFzILGRt
GD4ez0pjT9Hm5H8rtTEp6iIrQsEE7Iy2awdLys+1J05V3dgl6FiErRnhXVcj
4HmfmhEblcmJxmm2peLy0ytm4jpgYQdXGgjku3QMAS8HUh8azzeDAi2ncFdD
BoRLKxvVzXckNWEzR4UZuGc+ypMUmaAeueJ8d1JyTapKZ8aLQKWnK/1FwBfT
fsA6uuRzzovpSpSIee8KGHrAceC/hhQPvCxqFqbmHq3DYUwMh4eZzU1IwT1d
blCYrBNhh7+HxHG50HjQ1LVSfMVRDWHliON2OXERR/pGzJKw5ErDKMdwrbVR
Kcv9TqgK7lsZN5e4Ft8+IDIEFO4bi/FjWMTnKohCRWxhhNMnNpZt1YrOmBA9
tdP706fNxT2VnvKkWy0D0Av3q2QIagMojAFEBVpuH0bTUXEqsBaomZYx1UPL
7O9fZh6vbdaoqCvntrC9fN8/g35Zri+hLm4Vo4fwqxTWRiOTy5RUFPsrm28Y
3FONDPF4pe62SmS49ZRMP9Cu7jIHC/6XFOjUoGTGYjtF771inxrI8p5czEjA
wr1d9ivF/Yiqnk5VNS0ESz2Geu88CA4PAcPd0Vcs8GAlylHLF3TEAHORSspE
wmn+9EVsYSYbksBDt4ku2fTicM0ViTp9lutwC7lEVrLOZgLxczom+gJRQqkP
ev/oAkxPI8NEexzOST1BU/fMlqlCT9R1E1DPUE5jSd5pB+hNVUGkyeA3sLp5
Ufc7qPHqiMWDiltoWqZ0+pb1RO4L2cw8YX78MEeK8WIgoJfuS1erV3Pbg9y+
Y6eMa6dQ73csQAe+SHMVISvnP69zgK5OlZYHNc2HSIn9wy6zdqCgLWPbLi0l
B+MT5JfmIUdvLxBG9h6SWi2yr+oy6yAPSKgx/MNMJs7WG6HRtsF4Rt7RaeAS
IysPlyuHvNzUaRnmJuz3qViPh89LZ7FAP6VHkYzk+THBN/px1nBEOLXmbWWW
bLtqAG0Hwn9+RY8hL3wrhqnRL58OAa617ZShcINMuooqPzulIBTBT/EWEGiP
CPQ6ezkYwG9ddyA9MksN5EoDSExvC8dwXOYHLr8hrmXL1XD0o8kNeVBSWxMz
WDMEyqUaTkBRUcMZnu7eRvVBBUnPSKOiS64jLy1RRKuPem4fboCQlBczKzVr
UtBoE69dU7C0cnsyp7jsd7NZZXDZkauUlBuQogG2eW6gm7/JcJsPudVqjveU
Cpr6UX7N5VvdBpDIJPM6VG/iMtuf/5DRqhAQUC7LFGSrf5hi61FAB92ojkOC
r1owMjsbpa9CpecgBBgopGT1izuCDlG0fvCA8iN+6KPHsuvzUFkyvpVk+FDh
2gTxsEZRzSXJ8q/AI6JO8Adttk8yCZitqO1n7xeajg9Oq1o5a7IVAOj9e6Jp
YSBP3EwFtwFF6v0Wst4lGKBoARwBEvzFfVZRLJlhraxB2fXObB+/AMIcdcBq
VWuw7270rB/kq1BlCI9zeWCtkLkhmN6nVxBj/IsWtITVnDHQV77YTFDu6sEC
Pq09QBEi5b4KjZpG7lCkD7Xax/rc998NSrEXG1UDA/ozLrub9iJocq0Prtft
2ByOPCdDny3IjDmyHuVqlxlBxOnIqq5hULbQXo1CHOMNpk/SZpmxFrJmeUCC
XQRCJggiFocq40NoZga2IOZhFOP1/xCgdFG7y/kgNRYDb1WbwIwN3odeaEzv
Pjb5CJx9SK8OLEGEnODZBvZ+A7k0YScyMvJ5Awnn+mOWeokHDLfjK/uTJDER
/i0af5UVjTtBQJ1AyuBoiPpmmrPBfZJtr5clJCnDIvBzxmezcKb3svaB7F5o
99Dj8RWCF4ACeIBtYDgnkqMBU5I12VTo2sGZCoiyg5oa2RJlVOvzx+P+iXMF
IdXK2RHPDxaxN3n+tz+ZIIe4Hao9U2pvm/Pdz0zDeTxhGMbEFJSNFhHc5ofG
0QSVLW9Xg3cAFiIyiGGxK2T7Fi6utXH1Mj/Xvfrw+ESm+/ngRczhOyc6abYK
fbjq6Hc202KGPvxJIf8wu3+zUVaxesrqZxxNTAHFA1MoppcXqmvlhe+gCy5X
2aoD/rz6S7chNwxlN/9YbY4S1WKI5XzHWH8LgxBCBXzwrvDrvgFM9PlsnFoa
7ascKifK/33ZYZZOxf2dnv8YOnjM5DNsHaue9NlkL781V2msK1jjITsBVXk8
pYMj12PMWUJ2qBgMTLfj32c6+DnCGaITKECx2SidngnhjxuhvCp3ah6q3jcN
dknkBAXhtyJAhbeAhppkp2rvID7+08frIHpL5Ml1QAUvToJgkCTsNVGLrg7n
HfRL8Q9mheHeF+20TROSK1W6z/46LBnA6n/8JHLGOWTATlH7/L1KPflbzvyI
8bABTsMibZ0tREjbIe+aB4KLPuSOHHA1dGpfLSlSSlwaKd0LgyaBzZ2VjrYj
6CoHKq037rDo0psK5UzxSpX3ZQzUSISHvzp27D7sdDkqUw+vMXTgyGMwR2DD
wrV3Ss2YhtiTxcFGXORC5InoASrGFnfoYRqQ7aIeJtIEQclGiwVPkLWCeyNY
idoznFP9nR1+eMhtmuMNooqV5Op9u6NidsLhmuKPTaJAdcf5izY75xxkbUgN
SZdFL8ZJLjbPDoldi6G46zQ35vOxm4K9YWonlyBX8RF66mmDfUx0FXt54AGU
BGg2Rc0c0VVrr8mcpmE2J58Q0SUpCyHh4Vz9vR3NzPZeuahqex5ZAQ++sJ2m
6xO6CY6tkfteIT1AWUrQBdLhH0nucGOnyB1hVUm/rjMtZGiXglDXWE14ty0n
s9Iq0lT08i5kh6cU3e6ahuYfapM4yzxJSYMWjrVbQ8+uorgkvuT0sbuROLYi
WIfXkq153mJZZVfJPlhFUzI6nM6UXLanMBCQ56eWs+CcYq0ptW9e8/uNXc7e
7/eIy2prOy4m3JVglHMBygQ2C2i9g70bGh9MMqwk+RUS3PMbqcm+Nnn0GouM
2W1Fbt8HiJykePU4jPu/hVh4ei+XJdRso55b7w4W5jPQn7gHmw9yel7CrJd+
nrFkzpVkP0cZ+TRJoi5Mlmn/HZwgeF9SFJpxVfi1Bhf/Meh3jUnCso7tGqao
I5Z+J+HNswUhj/CYzGOygxIv4bdGN5YsX8P+5x7jDASivhuZczDZ16ZvRhYl
fPlLgEz6kQNBupLArC1j+ZxHJQTFWEl2I3o1dJplw8LWoSdNo+3Nxp5k1muF
NPY7Rg2KBPjoJxDoPOo3UNcR019FXIG3XYFSoLeJspTKeT+PsaVp0/sCfE1c
At6BFAiKiiqQhXKImPxI5wec9dcsLxXo+xq7Vb2e3T0jIXPYjCPP6HRzBafY
CZtybVuXfszfkawpV2nB8Je6Scy3NZyTuqv7d37J6pG9YMiCm6/RfdGF3uNr
Jc5YDQ+z4bqb93otTt8QG8pL4IbLb9Xtdas5F4H8dphqmzXMyCo5SZ3Wx2IN
ogPrMrPv9bDfhqctip3/kDZnlxKIrO1zFpIJnKJEkTUxiw+DkpPXv5tGY8VT
KfhPhIDHUgt5+CtD4D3o9fQGu+qflKH2p4lM4VfOGNG1JsycNZ/JwCYqk3wL
YPAFbpOZKAHRjaGHQML1Yv9hyF15LfuG0S2BaLXrg7YZ7Q2416BwVYqoyYwW
hIm2lPIa68BawiO8O0AO2hknuUlGYRrFN26f3yorGEZ0UKxoXd8xNCsIxMOX
RvsfYUjniAuHm6tSSKmkKXnbpndgH7uJkcvhgu67tln1OrWDfiQCqvo/pcn3
jBNN1qZcLvruBSXaxFLYtIPQljbqkUUdYKTzWV3pRBm5/fv5dy4SMZSEOz0l
9496vjUnUa2+vXXuDkoSF6giDHvnI+YXdLBp/j2zdlKOkJE+OObRC72HnJYj
vFiNrzCjbbR8gMJlYY+9cTRbXcFY3WJhN+6JrfYwEzrLMnJkPEnJyF9Afw4O
16T/EfuQ09MUlpZ7W45bvCW6alnbY7fCVgqEzShoWxnGtZWekd+zSqseau1r
lGF3/i4y4BL63gyrhGx3pb/gZrSzht0Fu1RTgdPs12OUseHB5sy9gUnWPTSQ
NWUvHT1fClRwTEgBAJRa13SGxzNZJatQ4GiUmBSAvY/KvP8zgzzrK2z5eJoS
BSq+4V2P3asGnlxYawBsmgxAdsiKxoVEwz7GQOw5BSSFjMw1Rj3Gjmiyct2U
YyDkMJfmSAbKVty1bFmnS7iv1tWyt5zXKjUrXYG3qpwdr1ZibGZ9cRT8UBo5
U6pZShSzDMdqCSj81FmiWwcn29bTdQ+3jaUcH3JGnrsh7NU9NNSuZm9flAqs
MiZx8niL6EDjv+3eHy+FVT2WNRFsgA4hxiZBw0Ewmds5tYJUG30xPvPrlJbl
xfLLahvs+W2GZzeYNYpFhiTAFk/OnMHjLQujZVTOwDhOdft0G+QfeRvp8X45
8FaPDxf97PdBLotys4QltnFYk/eLna2fZjXyPrAX45iRlh3DPDhriUe8H4mF
9uWzteCdR5eos9hTYjBWTRlMXX2us78rpI/3tgEwhCZ9SoRUJWZ0w/CI9n/7
9/RG9mQj+bRhEPRgo+GKXwNs9wTDhntsOD3OR+Wjpw4Eh6jnw11NQ1C/UnMi
K3ompC5d4vcwW8e38Y5+W0sNl3TNzEScban+Qq8ZSZ4c9pGhLxElNO5b6/Ee
A/SIbPV9IbxQjd5w6RC4XOxTNEZe3CLbe1s9RBJlnZTnwB4poeUVSGq7Tz+N
nZOEt/8DF4yI61QAQPpi4FshRE3svkQn9NEZz/3gowPsVhiok12zv1WWe8Hg
EhAp+zNJDgkKFXi7Wyb2+sfjKalZd734SuPS2kOgZgluEBLhjEu0t6QpWys/
SqXH43Jd2sy8osTmFcxr6WxO9WmdUTUjrvKt+0BYxWzm58e1aS9uZh+oz19f
yZYf88dScEaSFl93EE3jcFCTQJuJDl9SHvSodvpTcZA25mYt0ODt+EGnE5b+
WGih2hSM+5OcXWNu2+YES8YW+nGa9+CliM9OqBQKRXsJyU6EclRVXAibNGPP
A2rNVKU55Et8UTx8o9LprK+W3ICIQOCIk+lVSkmceqKVmFBj1kisPHZpBk/0
MdL4Bp+qVv99HQczTTd78aKFy4wPW19kQMGiMDG9uFi9I/kn/LIOTmQCUX/F
08eUgN/4zZElBAjvQqUGRl704ydbiClln1/fTNhMKvL9Y7NkTI+fOGqJlIVd
mTpDWrO3H3sT1BQUpzeZLspE4T6/h8ecQzNjvdfLWcAeQkuCsZA0RFaiQcKQ
CLIaonlrscoQqmYFq1tflHxsr3BFe6nA/n/SUQ7jD0R8HdTyv0kxyCJ3yCJG
iOn9h/LjLNwZyFvAsT5xr7XSKtb1zAF2ppKhQIFuYCYiEixOf4zQbIynad7c
K/q3sM7jrSpCsblaQHJERxkbNNCMZyjtRZZjnu761WUvwyq2QeO6Hzu05xqQ
c3S1Go3OjyICdYnBZw5nW+C9n9dNQi7657O5K/6H4KVjdD8fzlzuBh3H9Mvg
XRZwRzS9TTgtj3T9AIF1YtlJ1D1cSJYcBGrtnsCz6ab8QGdB0NPvHx4qA76u
TU+qVELp0LyQxyw3QHR0BIA1cw8qUYNFwDtnvelVYetxYGsByTaNwsamLnLy
rHPgTmB7XKSuPLLyPnhyRSMvL9PWWUssCuJ7tJ0PYSuMQ3S9pQU8iOqe1kpo
2/Hmp1Le86fOuTrvz7fCdM3HOZMotMNdlNrGfjPgPSLqxtZlBGRWKspsHj9S
86q0ED6k4Sw9txrAnAFx4uOk7HptKejs9JMI4ccnAhHETGgUzK7fAOtz7294
SWJwqez8wlYu5zoo8YsMJuuANw3fDWCP7/BPbQTI+FY8alRQbwMwchvCNaCr
FMbOU17VSqNcB0kIbR1j4DZe/XCqQ53WWBxzqdZeYlHD5Xe45zgVGOC0DXQ8
0Nnmv/H2e9KkSuyutJ6kN3lL8UvfPdtNaN2KBOWpzZ9WYAp8kfGMF7N4V/Ng
+xSzaovvHsM6IH9WXxDBKKxWBGxp+WQLCP+FZB3T+cBYCbhvNLIECI/pso7k
+H+6pF5ybWbMSD/9b/M11RifV3BSPehV40y+XPSQYNYP2tJaBLsTsxnBzbu8
tisoZHKwAmubjlT7zk1HU7641jFMeVWCyuJrhJia5U/1kRihawlWSgDsbsDf
Anh4fsKJTTdILIS/lZ1+WG0xe7cyZ4ACAXYc5fU+8ANF3utMdSso2cqHaCby
fmECo/g//u3LN0Wai3IPwSf/C6ePFWgYSNT/0qgKNQz41gFm66W1k67dkP6J
rWh2GtYoDATFPrlVxt72HO1iV5Khvlsc8IUG1SUR1Ap2t89JMwbQgY8maTQ7
/4C7RRAr927U2YDkbrXwqK1qWkelCseTaxD1fKABFxpqqdVk86WUJ4FRoms9
wKcHXCWp8wZreXgpN2ulPy3zmVVwjyV310hb+RZmUCE34CccCUvIaH7ppUJj
NHxoOs6Tj0xr+3Fm2BBq1zGcxbyIa2tbaBEchhUe8TENO8F/TU4XXanJTzk4
oDFCMpwzvDKVSF780yfMG3+bEgzZCY+5lySqHOKuzglYo+sLJBdrC38D37ZD
+ZV2ixRjHw/MU24nGkKV7Pz5F65SedJF+f8faA53vjSIEvDC3ufsUOiICO87
J3WTRFr/NsCHIEBuzWd4B0ECdNlJ6ZfAr5DVdLArmEdXLVXAAjlBd8lY4ZG4
/DXKfsuE+lNfhlQSaA7nWKnjzb8mGuoirqzBInHALpeANWOlVPhm1Np7IXHx
7u7x88xc6CIcvpdPqgbzsxZEISmRBs7wNg6Yp61TXYo7TWO47lTZzOr1wYYG
HhGmjol7twNbFLQs2Qy6c9TMaNWTUy8GNpEWEf9fdjg9fqbvKhYp3JUaiicC
08QbcrHiFDEJNT8wfVgrjjavY4OJqAw30u1eZe9Mil7edxf0jdWMDszMSd7E
k44WCOy7CsUFyjCBFSKNju1sxgYpW5FREwXUSwxxhhLomeVBrWMxw2N2XmGk
FvGJ+ja+rTkEyPp/qKmQ+7UQWjTCS1DLuZ6Q4KwGjzLExyHdYeZqtcz4Oli9
nhOIEypmFa51+OQJ2pA728lq+Sjw6Zzx2F2ngCMOapvt8uvLrn/odz2FADNB
DdHNPUHKKYpgSCkZtuYK9FP2SFLp1Xa7O4ZhCsTC133jp8zMxn+A3RjHuVg6
uZptlYHN1W/hhXtdRGGdr9/aIBHXxGO7sryYb1fB4EjwmgwgJYFBlqCYFK0Z
vERlFWrFqC0KPYltGbbTpwyRcwSChrA0GzaoE8QgmH6tDwy7rbOgcicjSA+u
Tnys0YXjgDr5UITtrOLRAil+n+2evPsxD5NM4tkiO5FFEl3BhDWhaxgjAFYs
FsldMtgbG88a+Gi9uudkn4HlmrGLduiDlK1IujUpnjVPRq0wSpCoGCJs6xsL
b4STSio2tyhrqvCeD0TUPG540H+nD7sI1rVa32XtgwRj99hZyH2WtOp1jGw4
HG9LP1qFU/h63lQKiCzuk3dHcOqXMxIx5NKsedryeJr0YKGxeAgAlx90rrsg
MeY7g6UelIyd4PDtXgrgAVIi4Fyr+P4ynu1scaXd0mIy2sm9rgedRFvkWPhY
fZ75i/cAsi/XNKry2hDJSbhcmddqMt3s9qQqImlD6FhByKCltRGLDwoE6Gcv
ew8T/wzM96JYMxTFLsp8nWFJFS1NaPu02p/VMe/5So0KuTVnweN0nWgqeF5Q
vgO3PNeZrKb2Phs0k6zd28YerQfN9mX15vzC6Z00S2kOr0t4Rv7iSSqtZIiB
GxlN2ECOCv84DtkpMCN44bmCGeJC0gtwovRIuMBOIoat779hyo9mrZQcvIx0
lSB/XF1KFXMcg0+3BQNObI8ZISWpfllNCSn7QHDI5X3UfrhljTa4uOx74fhG
3OsM/Ma23XHEhlHBrKeDyATjdoXqdnqHb6ng/2CYJz+y7WkOQf5gwIbJ9PD3
MSaXivDWHv9If7bur2l+StVG8FR72Sc4AKY9u0G/HqCJoZWbd0FuZdxQh2dv
+T+2uApgvW8M4F6qOodwmsRpZsHdMVszJqvpmTikmcsyvtd1BChKhFxumo/E
XJSd9rmyVsn7lv5KJhSiFWzOlMLao7OEIP/I3h9ew9aUf/3zCfBo2hl4UUDn
+UiIeC30ToxH6l9GfXrAF1xq0ZsbzrV7Zu6NFnvNzuY2PQL9ENallhjTWkf9
hsN4nQX2q0K0P+2z/4O4YPs6uc1kvOiZyC5fLDS8rFEYJaxcz+h8IOLdmo3V
GxXmsrRtvZA0rF0u19DmQ7X7ioqyAJ/T2HOLnHArfd36ddTkrXJASK5ROUAg
GuSNdh2DhA1bXERV9pDBP0EImJH+UBJwMFmTG5Teh/5ufXWV2Ko8HfcvUUqy
y4Y2hIkLA8sIIRJ1yn7MxUEk7SWm2rKmMzABCXfdjR4XoYgt72wE5UFl9SAL
VW89je9oD/AnngYnw32Yjom3QOC9cE1tEHvNv4oQDMRfj3uYJXcjbTrJsMeX
NOQt/lcaJ6IB53jfBmtgXL3vwuPFEVFFU9I0/6rjLM8cNQQd8kfaSkzDgv0k
EEQwxoyc/7GTHFEVJx1QKXvd8NTd/YYvea/NbwtmlUbZmZ5L18GrYOX5hedd
vHeBAzThe+7dh9ryqO0WujOA5ROQH8uNdx3bUhB+Yp0yRqgpsZxm16Aqgn0q
K03hb8K+VVh1IoZNpw2YzVUzgSIVGN4Z4m2uC/7XKe5f0V0M9V8wluh/BKud
ETF9jXiipSMtO/D76jFvWqPR8dBAMx+1n+QmMj7WVaKx7Fklrw7/RQ7fut4D
/64V6S947/zCuozo3WDRg3wIpn4v9CpRxeWH409tQFyZxrjj7721h7DK0kxE
71u67JNoIhlUvB7d0YxviPJZUmk3zXgLMHSf8nEItWWRE6r66JWswflwqZRu
qLMy22hgohKKueBDuHhpzVHxReTBe08hgGN7+0gKg0hXM8IQ5CaNIHkaTsC2
TUC0A7VlwmO2sgZ3XAo/i+iNSLbtF1GmTxY/lsfit2bnTJnuPXcKBQnvCvoF
/YJaD/HWKOBWb3FDoyO+TGOO7ggRFwtgSeWfj3QBZjoKBjg8pOw5iWirRm1f
lhrRsqKoU2lR4cNlWCKJn+bM/vuWjtOs5yM1gtPVz+ZFYbUXJTro2TgZwEXU
jrSclqIl03xbcjBnzGdh9Dh2b9l59HrysqyvT/NFSm7G5dsZlSSHPcBWS+kj
Pe6YRGqRzbDCGj7Efxjl8ly50hh7D789+EViatyC9KsAcsN6WuvZOQGFJCTP
TOeVbZLR7trlQLQa1CFBZxe93UoBcFluepmpsvrAhviRPv4zvz5zJhl76yJW
k9G/AyGk4EEXWv4oVBN12KcNY/mUXkKRsu6imum9fecoVwvjJJW/M+1OqAv8
haxkq2MRJY3/KX9W6IMsvkYfZ98wHaBm9pIIWqApZ1SD4uSmDU2TGBlq9NBe
q0Tz0t5j6iqTqhzctwnhphFKPBWQG+Z+th4vUuI6cYexGbBA7p2BamXE0i7E
MDu2nrF3RqMbPadtH4a2aLLTId2QWHmDsEqddcGb2bVbkcdwPI0lkIPsU1br
E/5rejJGjEfv/rw8yoQPR4hGxiStJLK6uXkHrt6flAxZFOqzuA9/XJYQ3lT/
4AlhctrAYq0aOSumT2L2vwb/nJPS5YCDfSw6llV6T1CkPDa4MvPY86JUhWqZ
hJ80bPZwB+rtW5PH2FcsNgLnp87hVr7n1aeAehASINNPVsMHz2qy9yS1C5M2
iao9IQqNzrS4jSBkLX+Drcp3F9vC37/pR+IChsMMlICrVckUGadfAvi/SyDI
c3V6UOkirw4nCc5MhTtCgWg2FQthvarYkc5yvQQmi86FT3gY6LvDskcdP8CD
m1jj1ygs9sleoSFceAlyV9Vx7k1PL5qTaHtGYhkFmFqAQJ3o9P57UiP8Ks9m
LMJoDUBRTyArMm+9xqpOZDaSS6bdahb7A0R75by3nq5nPN39PBCyDsnEdk5M
bORKR7LXjclsu03WiuzbbTzUH4oL4nLSV+6t8ZWNLmRPoew0+y37E9zAft8c
BKUxKffwaaMLRzU8XQZ3E8rT+ZzN0FhYk6chgJZqP7T34VvOkCAmqTbdf/iy
FALnH28jXNxh8SQwkBZv08MP3ShdA/4IxnQrzlCpHmsnlHbHtcQIenO8/yQG
mxXohW96it/+p7Pmx4XVHNHUiOWPyP5LURKdl1v0TtHzFVKv4YJlbjbK4LR2
z7hX6VNXOs+/IHji7RYNuLkZu8TsMPuCbWNet1PL6okp3rbyz2CwjNhHjQKB
ctmI7QMafLn8kOiLI8Mor4LOyFYGVg7MHeTQ1iNxXUo/b3fSAvgkef3SOqMT
NXm/Ybg3N1HB2TPi4D+a3KBUiFUDK0RoNkrjrtZjKOn3vD5SC+55kZgiEMcf
78CyS4BXmMUxxlcMz8lsh3w4tiQhKW5vYyYRTnACiCKg0rL+I5exf+/7xKe4
Fsz4+bQteLpqC82Bo94B1qxxHfRGlCkurkgg57ORw9DsiF4WqxDJ2UKZRkU5
XPCDgmL1eaxDlalRJiU+PR/cZE7MKM7ymPuatDRsK8IjOkuvYlOxRq2xCyQZ
1vc0y+4GoxdjAWh9xb/cQBicaFGxiSzM+Ls/TQOvZh3kdXLqfi+EDMyNE/GF
O9g82epm28or9zK89SBd1g3cgcoVEYdGqzkdXq6ZxFXse6XYEeYG+YeNy5DJ
KxSQ06LxzOsprvmVJiMpnv+vmGdtEG76QwtKvUqdQPlkLDfN9ZFb4CKT1p6E
FNvKqa5J0XijCRMswlcLHPoGOoCApnb31CeWxHoQ+R6X08TCNbReFjJb5zLb
ULVrERTkuJvbewC4TfmGr3qAc5oZDRXGWJongztgY683mL7vIQGROyO5I0T5
pBc6MvBMhM0qJQVWoBLpikZULEO2FoH1S+EEZdIbGUQ5rgvzTIDvlUtok060
ry1Kfv9rsxEJzyMVQ3vkK2v2TGWNYnOvyv4l2zk61XxJCzQnOlqc4Qhcbc3X
SuIqdUBatKfvtj2LFiUGqLgI4Njp0kp+i7p7lIrxi+T7ED7yU6NkviF9uyWu
YgaYypb28kMEse6+O8bl2lpc2/LVo3re2xy+oyRvNV+p4rJuRnSn0bp6IJTO
siawI2IVKnD2jneYr9XYsMoRsWsk6718heNdSukZM+ngqehtH73Ww6ba1peG
f2H+3b7AtsFC9R/LH3oBhosQhN7vnoCM4qSlsjWd2YXKIR0F2KICqSrJzJ2l
tB7hpzBAmLvHf1LuUMFK6Yflhj9kWr4OBKuWfNYiwRT3WKa9j00amo+TDZb4
tFYI0ItreyFzT1sWdnVIpcSs8obyCxtot6Gmoo1ifqMEyag/BP+YepSYQz+W
a1hR5pOm5bUCRybvSJOoYKmzVmonx0MJMu/nUpTTroJscAZYsr0cGsGze2Z2
Bc6YOZ4FBcqh57Utqf5eO3TyYdMxnjfdYY7p/lMNfoIu8c9QMbZGylTlvxpx
cffFC2S71PX+pGD3GJ3I2vAOxlrD4rlpFI/nHTAaCYmuUHcdcQ94CAYqLhlK
9IjbZhRptwizjwcWTH7dvWRNx1kNtkyFwi5qI7kYzKVCTM3iPC6FUDW+N5hb
OpfD1RBVxXnqnWmfOH79b49wbOQy2Yqe0BMsNMDH5Lxrii5r4Jx3iA/2WVNt
lEQyLr+IUlmLk+5cZnQpZ7Q97SyO2HU2Zsw6EIaxFwrTdE1z9uumVtzAITfc
YGwtqnKSWjglzIivMyRkUkmE4cYc+3E5Cv7qjpWUSStErpgyF2ENB+IhI5Zx
d6+VrmdVWxgCKhJqj8sLJqVN5KhyUZYhmPDy4zmx4mApH21eJO53hYYTrKgX
bLTHyHaPNLktAeqSky9Q0D4FmdOdhzxrxvSIdWzWIh3UDphJvarRFRxgkmgu
NOAWs1QAKebyqCXMSLGSYHhmfAdj7V0qWlugcixvUoBeNxuNgmCBjjq8xU+W
LPZLANjBAfJMRvsfj1+4WFwZJA76hfK4600dSpnYYoW1lug/uWHGjgCymvb5
5ddUli0FsQXKV+ZfhLUEyG5OLA8klZgkM9JPE3Q35nyXUfvAFGmVTvxSbzpm
dCbtuUFk0RtYmEVVWG9lASsjglIUW5F3i4WEA71wbRi32YujcRO7SXeG1FW1
efNd8X+mBIexH7/iy5ynD35/NJ5Q/zxGVZhyKlz1rwEzvMWs/hGajIm+T7Jl
1txjeMaicB/iovJRbGijjfR0h0kKvW0Uyp0BXUb5SgkOqoloSbRB9QkyeOvn
/bgWS97gRoFyVjMC4xIA8SQzjihI5iLNM2ox4UCGbLpOZfaVUJxuS7fOJKOc
VO3In0tgDyYbZcAJ+4TSCMxAQdS0e4Xlc9kjHqDSorsiXOS7RieWWQadMKru
CnQRut1oFqsUBJZ1eirKbnvtNtjoKnh+q7CtYfa8BPzl/laz4p56dvSsZYC3
yYxz1XIO6CHxcXqCuOK/FTHzWMgETmBqMo89737TFv8nsEjTBFhdJpEdo73r
1tr31WIvpi/g6mGw4uN0+/uI2RyNr3R4AGVRjrDQ60QBzBWwjyZtqjJDrFmp
WxPy3Gx3kIUM5+QbPfgxjL08paLqLpbfkwViB6nGH9yhx9lCTA4/8pm35FpH
xsqdNQlI0482rEkmWmfy6C4vNW+ZhbQ/vu8OkHMGW6z+oTLKPIeqfqnyc7FG
NCZTbMriYzJMHw4NCAYDlSjgOTUWXlN2aEoz4l2IwcUlCkLT0E1ln9aNgoMC
NstD8HpTS9J0Am6LaNFt/2UpieL2pHqkkg2vYrRHZcQckVkQCeS3pxLZeFmA
7a889O4CJK4HzsADoSHz5HDTL8B1GH5ANrdupGN3mmb/ePEBfMveuBtZFFp6
hF14QWk6OEVvSgABSq2ELchUvFvH0J9CQWhr3PPUu41p7qkuwueKCCgO2qbk
M3eShflGgCefWunJw2oxDDpFMex9Ro0f0+/1ij+NEA2YKegm76UUjCLq4sxb
ZzHVtmosCl/G12ZAkAUhBnXYioShXRywuUOyWRrP2uvZcwhfv5YtgGsaUOBF
bMar0nLNzX2qbDBs9DnFn3WwY380dirkMYPgyXTsB9U3DjCo27WWso0X23yS
78rUl66NuDJyr2RBFB6XOhb/IlbMmit5+I6YF7uGk1dJurQ5RyJZfHV5D7/U
ezuLP4MeSG52JnLbcOqtqR9ARly/PJE5UsyUyPwG6rkJsPqf1gYeLshr9S34
8M3i8vbqCSOLiRhDuXkHtBXAAzHvZHBlKJ5MT+FbbbiSFuX3/7s/q6Qqgei8
CfG1wThXxOOA4bMcJiD+2/0sDfHYFyWiI6n0wYmMvqEI4wL99+NzvohORj94
3sywRR8NwSXwn+GhRFzvanuWkAysQt/c06w0heVVpN4umLqMT8DBTNSjdGKX
Iqyj7PK+U0ITpk2vU1pPltjQ5ApBiHg89l4FbM+fquPZJ0kYY+y8NW26fz76
GbPiZmWbxEyg0IuwbCNLRen7mFwNgHvGsrqpEYkMOcYa7VsY+rWs8wZW3t4f
9bHLtOIiZSy1voJYwQePg2UzrO/mr6gr9dUKishtKiqTAYoyUO4ZC/nFeXjy
wNn31EgfG8/K/TH9ma8/RDu1zMBav6sbSJug6ApIXG3zepZPR9ls22tMOq2s
9k3j0AqWY3vEg1V91yvT0nO7dsMhN2oP9N0LLd6f/Yv7DBg0Xhwyb9zwYNL6
2bWAX0r1Jwd48kfuwbUPjXOexkKC4cn+ntqqtE0ocge35J1bc0fAE7DYZgDF
8jrl0Q6pRbbVjggX3b0WfktGcY4Puxr9sk9us/uJCv5Vk+TVZawXZuflncEX
cOoNEjEgeRMyOaBBrOM/N1FQ6+c+BWDRGO5OZ4phI5qwdgDiRrx1qaxYWH1s
jySsTxA8glbQiCsDW3E6Alyl0k2EeMtfCHQmfcBkwphufjbv9CQ/4FstbBhe
iHrjMy/uY10sctqEw7m0+/lISYC8sWnpph6uHj9h+omTWrVEGST+JqVwMi7t
zbNyZLMC1sf3ZvM1lHme/v9LtH831EXm8XoDLqT/Cpdo1im52QPrBQ+1vVe6
ofjuQ2bqfm4OeeVFmQMXTNehJkb/oCRM42u051/GQmtev8BVMc92CGm5vKhC
7Wpbw9PHUPiKSJZkCzUQGT28vK90kvEagNrPv0W2yG4zGDYeldGCXrP2tF3z
1duQequeoG1Irg+NqJpIxLRhfQNPKj0hbsllqd0KtiIm4WItNiHhB3KzjfQ5
6aZcKorWIicr2y7kNtHxWYTFfumKSDCs5q0zG+AST4NyJR7pmQxedmtceVQJ
5MWRxLM+kJE/D01XNuDH+PJHvKc83qNrJfoddUcByq5pz49UcRKAd+EWkrPG
0t7K8PUdj7XWrSYnMEY2J4GlRObaDgswMGc96+hv+d+29JEehB27LWwcArOw
ZWb8SQQJe/PovvmcKLPuCuxZwITVZrFGX2yGpAMmOkjvEd9+27G6AQu/rmJB
WMDEDWu5lWrY0q/ZgjMSB7eNn4Kmyh9oF28ic3q/35Lb3zd87S8njdGCbY28
3ra2EwvzAMbJdtLrvAWjosyB/4xwkqalyE9llf2MoBR3Wi7ldJyKcbID6Ehe
SZn+RxNMbXTjvAYR2FoZn+fF34TQJiohNgZIILCDkHDmCJkj21E57FRqtnFC
0QQ1cM8iAB7+tdghdR1e9707M/1fMrWCGvhFpHm4JbjltRsJGI4dwXKHHOYp
80n1jlqpWl8xVV+UkYLj34XZIl+ZfxgLcs1/yOOsELEn9AdeWyPkn1m4ugeW
IdGpg5sb1X6On0ft4TlBEQgugrYe3a7IQ5mXyFKO23ysgwDmBcm62O8+kmTN
YGi0xAEZUgrT3gMBOLY6pkYzuOq4X4pi4V6L3w8EdirEbQj3lypSKDKPHiG/
ApzAaVc9HnZXXmf/IcZWqJUXoheBHIo0C88ofIV2hgV2BnzmoARtEREB2nME
04IS/NyHEYwHImgN0GOAkFxLD5Put1ANYYLA1W2nnL/iunvz+HdOm7NfpxFh
kfjORJJODnJ12THswVwcq1gUOdQJA0MbzMwDYj3qxaUITaM28pDXJeXUGle7
XhTxGsUpVB2aVcH4r/GDoCUS13dvrLgNcBPz1XweOZT4NlsnrIVqR49YsE2c
uCIuPb6KWVlWQL3v6tCCLPyikvichbaRU3Xz+nAA9XvbCJ6C1ZYEc3NGH5Vv
J0pTcmj4WxmYHAhojm2LmNhIXxzY1QwxKgxbmtQ4ONrEVpk546X7ejsMpj4g
mT09jaPTZdg2tmIHkbeLI/5qZNzUMk2zfo4L/XtWchaI0KnqpmmBt7UMofMx
JrZ2q8xLD0C5eVrcDlko3pKLj1nMWQViUzb59MZsnJFPzUbt83O7Xjg1FtaE
EWTOFBN7dglRwaplpDBNxHbi+zAReUl0Env63r50u0oYKhXkRjTjTZQkYm+Y
JDCiGfVIAiKovsDEsHo/r8kClaxXsh0gZoY96FLZ4ZTUzrH0Vq6DTacMdNAO
T3lo8lpgI++nwyZUrC79pFG7JNwd9AQeUlMc8msDjZn4lOan+wx0lKMrQJNF
Wd4nOKggji1vQzqxKfu63N1G2GDfk7ctcht3jUfIBcJpZn1M4CrW5gmX8c6F
ExDn3NvtCCW4LSranHkPnfRbHCUo2QiDLqXAM3LmVvS2/+dwll4R35SsS4EZ
fHYVxCHnkXWTiUKCOMDp9ehQOc95oDK8RSOQMY+GoAmgXlpto2JuBdijpQPW
svKWg1DAh9jNw0w5un8AZakzGQur83pWrs0hwAyPkfK1iuADbSsC3bik0wG3
C26sfr6Y+g/FPiQZgDIMJmAE8vPfbFyOVshTGTu3k0AnT8MeQJ48VKLCoRU9
CDqmtIJNIRVXq3knJHpP636HeGp2/wTdm6JsY6JRGMySBZl7QKYHRNtZS0L4
L2XdJMGlJ12YnTmoZuGPUlq0nUdDbNI+pDFgGC7A9zeinudTuIs1xH1sMKSv
Q1qKgRq5OMr09WBQxkXO2g/aft0NLAudxS43owlzLoH7Nzhc2XuaAkcTiDAZ
60urBxiakQOpEUY/CKOlmfzWUovaRTi0EcudljAEHSaUCccmyawMA78kil3N
MeG+IM1Y4U+NdZ7KJOYRcISbrEZ+i7G6YEWdlAOgUlZT4mRch4eeOtslNzcj
DkOlXxVvHa1k6Uvg8mbWiRgL8ho/1ooZ+CS07CfYj95iRvisBxTr5JoxOSDw
VkjkOC1VKZ58WguetG4DFa1jeXDp8cHSfLEoElT2rhReau07MnI2n5+4PBg1
YWQCsP9tyc8evzLAPwGXOmxjlV/cy+udQO9qP3qCnvnbyw1C9c20xfdUJsqO
T43QfxN7jSebQ8sGqNNTFAsdKR1EDpLVET1/i+DwejE77GfEr9h/cppW8Gcj
wx5Q+VQaKJTGMxu3JDHPYQCTmI79MfeZQrwN7xiXbWwUrmWbuOoF+nCwSRfY
/415uBNu9+SGwpAsz1/N5kYqiQ9/5fA62Tl3VOO1dphxhAx4DVT42+/dkfcM
xj8mQ1A2BMdwIv5oSVZe2EXAxfxmKXA4qrRccoB/6laImCeOAC308tzybX0b
9KkpqJzZzwPJ790Y4p5Mi129gsFL016oB9dXMhU50zV0WXLzG8ohfIJqQM9q
d9n5w8xBhJ97+FQTu+aHdpZYopPnHfTfOLMxqTURE8NJPAHnzVJSIj/hjDOg
fxrF96OukFFmPXBmdmBiQiZwG1RGmhmJN7xuT+7yU2RASb6dIQ5XlmJJyZp6
aMtdkih7BZIFBn7iS0QHbwW/S80vtFs2tt8X9/wplFO1ESISPPP+9dhe9C39
aJEloKCYrqs9Ls8hvpKlB1wfJ6BYdrImHLlKd1k0Xu9XKzm+iLYyCapQawQU
teffMBPhQl3h42lMnLkLAPeSMWTUWXQTljrwc9j/ZBXGD18XOmi9CLBXxNRl
lnaXj8yzUd7XZvhq/hNUIFHGEvw3ztK/7/BAOe6QeeWD05mrBAXjgLDDMg5b
szM8HejSfPN7Dyxmjp9C9Ygs8C9b2FRFmU/31nVuB9MQVXmVw7JwN5NOMS0d
RUqFMKCiYApNHfMLsJWoJbbSqHb1LTCRPM05WT4yvfrkkEGE+eEswkhNYjJX
uoBEmAQf33uktsa75q2bIBbPLgjfeSPt8djXFXG/HXm52wLJjDGIUZT6fAT0
+6ryHMXeUBUbNYgvU6BvDz+/3KK6K1sYfkK3zLriS6hz5sPa+f91Hf94NCs2
kxwd5uWhqNcrc8a3cZVy3dMl6FrW3ESMw4BpUh20ImnTQWWpIUPrr8m0C25N
GC+tgw7/zoDl/Pgjg+kbBfzHVpNfGSbcjFrnUHFI4/VaYo0X/QGYDkG+c1Pp
0029/V3tgZBKfTeHq5cxUXyj8X6a8CXxLAV+CUHWTjuNRtAgrkXdVurIXxsn
0HSyuFaJ/jYgModzRI4TS6xhoCHFsyVV4TiU1L0foxlK0DuZbJZZG4MSYmBi
BurzzNwjws3hTxu2ncKBqMMGaSp0fV2eUob9ghamrNUTJU3ZOqMQMIZKwH6R
1XN2RxpF0W4HySZ6hDkXsumSPSR8LsY3dVVQN0aEdgk8JbNwy17x37crw22Y
oC7OIdhDfLacU02WyH/2kqSC02TDvX212c4NamrZOGFOR2yLUYJw+04+be/e
SF9OU1z/tDdXj8lf2eDuWLR9A32CzDrLtBwLxkz6uGSBI05LPNqx54arUsft
9AuvT3m18RYsjO7CDOxadiLB8WiFesvycQqYb+yu17ZY61pbR0CWUDpyErB+
MUYfuE68syDdAQlalLccmE1Wq4dSQemgkg4hHfPTHOya+TPONOXQ8HkZlJzo
/Fwg3epR5phQ8e18pgggftXQlTvUfMnaNRmyUrepSD6KaF3ONeVatICIzqgO
4F91HUmSC3W60g5YF3ofD34kEI2K8ioZ/pmTQq4y7F85n6WGT6wqsgzKISmo
dIpRQNZyRJloPcRbre0dO8TsW0BPQF7NXJuFjuVgaFL13zAn6gGjQouHrNLS
nQpKcZPv6lInwaMkDMaen28XEi5jIjnWntNJ9k+H5sTpAgaNBo1pZFE2er5j
KanklxfcUnmCSzju+1AIi90zVAv4AZsxDxKNNTrmlc5xR/n62iR/4jtRFL5F
sMT46RZtSEXgc/x2/yFrTdZenppZfypTTLnrBdeAGpc14SW5uM1B1ic02coO
PnGqua/q+Oxt9MIDQ43ws3GgwTT39+Q0npNtiAZUlHAvzGxBGZw8CyMRpofK
NvODgrXaWBJ9aj6CI/W4bEpxwxtJPS4Y8NnHAGZZiA6vXbEEiAfWz6lvMk7c
Y2ieuoL8mah9+i9O5WIVRbqhWeOzjQJnY1nhPvYKuHMKYKrCzlryhVLqGROT
b9EowWEdA4UXsw/ilh4X9uZzYYaoYZ6wjqhJEoZB/+zWww3ePmWs3IiBIeos
2ObYzyOv19me95yh0B2ozC37MU4hdrXDVH0Dd7gfIR0HlfrOUmbdmfC12iCp
85Ah/WqNbSJXXjyx/Mn0QU7vPJ80+AByvfhni8Ir1m5LHoj8Jfe5Y1vThxLh
/0rfPps4aGa4PTKtHltIA/JWryKNaZlkTug4eNdf/SPhTbqxVI5LL05CkNh2
hV+7jFF5q7Hzf6AMTlmuM7uf43JJ1Ih6TVAMehgGeh3sxdpj3SCIvvP/5xxG
NOiURN8nmdxzO4XGQkv4AO45nFdiVWtgZH9fzIxHudx0O16q7ls9NJdo0sy0
+TT3NSrCq5Liymvu+VEtZOh5kNzDyp45LDKIctTpzBHUpZeF87jFiux86zQg
ydrCwwURFBwBH6bF8B20jSpCc1YqRSnZz7ETtyJ7ElRwRGlJ+jqC7YZIeMf6
KwGGh3rrYMQ3/jyfM1SlB4CImX6TlFV/9uLlcuJIVeoJ2gBFbfuYelndkrzM
2KTjkja+Hg4tLVPDX8Hy9TMERJ6Q9uentxn6JwIbhmvM9O8CKDZyalhHt36G
iWlH7DuG6icdonrMxWQixVPhhdoHTm6hf22ussl0P4fje6LBmdOBOUr4uOC6
X96UcewQhOuu0A69xPaaPAIsBvCGoo0ngevmt6oM752v0Prq3MxPKJAqtXxh
uqbqZrHUBCdLjIHfE4n1K03L2VdLwHgYuMRpNDxDYcSxcGhvFnHD/zsg8BSs
se+QGT0pDe8pIs/HuG7nhejUSyjdWH7zqfFl4S6wXBV2hkfaAHRLDPG/kVCf
XSsNc7miV5mYHwfuOQHatN8O4kvvQ5D10N4wmjDLt+8p2e8ypGoi7Yl0wKmH
Kq9yk51hjBxJz1lqczbFfZqfn24YMopkDTMWYjpO+FwxZrFCRld9I31Xnxe2
smX49f9CdzoZ0OKJDnxO0k1FGDdF9E3szteGgTnNo23vGjzrQOV1lnu0i9q1
2hQroMgbw3XcPs1tnqzxDERkHeAhXC9NpWNNWByb1w3CsyY9BDWxsgEhZGmv
GejRAvSrquw+dJTPjCiQ/RXR3Ym/7H5R9uxZM7dQIxVGVHJTG8EZXvRYTlIp
T96SnSOuwy2XIXHNDgK2wWmOlgTRfoFM/bnOC+baA82iibq+zDe3lLP6115Q
hAHOsrTbuT9KTPz9MrFepLr4EMbq8m68uf5BL/tBkHHTZVzm2LsRhzSxVOft
ctRnDAhSQiSZnpJCLfarM6NfWqF3PPJhLYWzmlT2IGsBsy2nmAp+DMR+1Kqd
C07CRmhEsp2GTC5NTmFiGW2o6J4Pcl37lPfZDqtQYs3hkDtRtZUfV7UbXMMD
KYKfAaV38aVlJko2H5NSegaj3taihgaf82msnf3Lr3O3EtUrOd+jCtewTUmV
LPvLO1MuXxE0m9cYLujV1bwHc92ZTkn7z5X96est4kO4uHqTd2oFE7raezGW
s4uX6b9wFZ61A0gWE0+GlvbRpV6FPu2aPK4JvIplvQACj3T9tIrjryRzxUJ6
uijMQ/OkbgbqwlBC9furz8XnQEs4QUBHLAVhIGvL6lnSzbHBSiroNiira054
SuiMWKo8UnGmwCEEtLxzYhaAr+5/bPm0PyfFRE1FS6h1pukSptARpFViKfnp
yIq3WhZpRe3vBW8mwNQJpGbKNA6qlGwxdtLpk8y5jWv8cWbUARFur+9eVBDM
5Vt15v7bbtBiQctBYckj3Kg3MSn53HI53B5NxOVfhOTVqKSXY7k0HuS2kM8A
aKXVsxxKuJr7jc5kWJrVO2XY7d7a+P1NyC+EiwYXg5FdGWL+QIvDidhGEZnN
5kqzjsxNjzzczUSSBggg/Y8NWumgtloSDiTwPKv6kYbWBKEB7FU7hb2JXImr
PNye4v4Kx4dy+rSuc6vILsqrI4xYJKFrwJzPwpcYNWDcQKsplxkOZg7At95E
HFv4clGHy9HC2RwpHvqpwqQkIkAPE2rn8+rD1FzkoflDhqgfS38xnsDbxy/j
zK+oH2NUZGOhBQHRCjlmy0y3fRtIyh3IeFBbQ2aMnNRx6UXgmq4eaISDGtEr
BjAonng3cXiI2XcHtvHHB90EcHCd6gTqIG7QZCEbxDPkdAa063w35J3/wcPo
RaRvMJ79mwiLrcx6Ipx4UVdzuJhvlRNyBIfSjo67aBf4A1Afgl5KAuqaV+qY
KeuiuWIqrbhBU0H/OVCXoRLHTUy5jbdxRXjOfpoYjvJ8KXCxW8/jqDsGQfp+
HEU+DMfr9nnVj2IiMjRBISPzPW18lIROvwiG7QfQMgkIxWzTQCKX1UVOnHOB
kciz7tlRtA1ejYMWTS1NOKtDXkqNR7fcKrNXoWPlTQJ2rbSMBP+rRfSR8c+L
QLgyOniut84vQmJSZXpULCRcSqLASTNe3R60zH0FpFLn0b2q8oPgb0no1Rqu
gGnRHtq0F0haq8ykDzsew6SB4N8CO6wtZzVyX1wQIn/STdLECGBbdmExN0J2
IjftH1RmRFgKX8fTQ9YpNoGZ+g9F+LgW0oacWs58yu/wV5PdQ15xd9ex00wB
jD3HZcT5d7rmTKRzsPgNun5kFNSI2meTVg9+t5lK7mU0uG0qDSNoyolEuLBm
pnSTWN+9BIBREl0d06eYx/Bjj32zYLFV1CnZRx54iZHk4ysAmku9jIPy+pKW
55OHHbfjfyP9soWyUeDYLxevX5soao2F6g2vSCxAGiWmOHTftiVKsxm//8hO
1xlJTRVUiCSsHLqRu9QD+/JR4bgjel+ZLJeeQArL/NVqhp+kFqCfKqEL6DFG
B8ac5MEwcrOCX3f3J+z8SoHalnTbYhjlNnmsFkyHlH7rcsoLXLzFJtx9w2it
+aEZiN2FwNr9A7toNzoGdkMQnGQ6Wo4tohPPWpSwfD6z4psQiJrx75Zike/L
Fbdx5kvP1pai3/yf08qBUOpK5xoF+kUaix8PsuEuzWHrIRpC6vO1uxiKy8Ov
jLFG0PkdUjmeZFRbj6YRz3P4CNpLqjpRhZzvhlCwYh64cW2mP96yAoK0pcd2
IBHBIcIuNM8p5yZwNbOwKtkIanT1lqzvVbOrSoYpynPWx+gaChVXrV8wKf5u
uZ6mlXLo/u4YHiICvzGsfJ+aa6YIOD3R/KxCPCR/gArwa3HjzCqisW9pdfD7
eazmOMih6tOfz+5jTnXZ1HRbiK0FM4waGQn62Utq2GPCw2yoNkFqoHNuWG0c
D4nXnAlFbAlN5Y5Oso4lVtayvf42Xgl6yqb+8cUPAkgwXLrwgqR9vyKFe7pr
8At8TtQqvIygX7tyVR4wgBJHXdOLSCM5a4BgjogreCXzunVJlw/lY2QhRKv7
tFvQ1usoKp3siPFLpF1JByetzFLPh4V4EILohODV6IEr67PUuc6edhtOFEsT
el2I9NxArMNB1eRpRuha6NMODhnHJabRVifG6PVDMqekt321XH3r0IeBgYka
hqCe1+DYEUZcfDsvgDg+CearXELQYYMvj2wzFCEKc5Nd8J1ddMnryBGtZXHk
MNZh4C4UffPuY39Fjy50SuRacWxCxkfoCjWfqmqdu/QL0Y2IN/NFfFKqfLn/
/g23aM7FTYTKcPdBT9mhcQ/8SH5vQUZ/JwXFAKmqAQPmRv2I72JMIRjxSbvo
PuL6mMopyniUrfVQitQ/jbRTJDTqAXQVeLZ8gnwCo7oETn0i5hW9QL7o7qOM
9x/t1qRLA/E2/3G+dp1YWCdFiVlFcfNDI9gdebgHedCO2feDQLzK5VlJCzD/
gkAPcq6ykknVupaNWvhkFoy1MT7cbtv77ZUVVhfb2ySWyDOL3y101FfKTtIv
3eBaSxmAvlqqGUBCTj25f4FEMhuqFP584qSsdpiTqmrMeOzXlTMJ5l4stMTS
Q6Nbacq/9kuA9S7q3hGe9Tt39U9Yi8aHhh+zTr2JNcW69egUWZtG9M6iTExz
lCrD941/Rou/WAnTJdWGv9QHlSDwasbV6691JttVUxkrKvAqnJx0NVozdOR7
COEG6Eg7/CsKTqrVZm9OrFEMocIztBVHfTpUCepjlrE4xVxDQ/3ph4t1RWXV
wDv8iZKr1vh036ycVezKX1mS8nS4fE/2S/Qe3LUNhJztqByAxAGhvJS/SVID
3h/V6ZcVl/6/YG51793Id+cLtC3GP43sJERBbpff6Ehav+P5EeUl/SmDvpKV
wVZHhBgU+T5b2/+Xk1hbIhIEYZCrTH/dhGdiTUmDa+WOX2Y98s3ldmb174Oa
CdVH5tHcdGI+edR9XCYH6jd6Fa8Us42K32cDiDxMRudcxavLw8WyzMkXSryo
cCk1dQeHnp1Ueqv1AYlQzIdpnCL8ipV0+/lIqntk67XPMbSMNn5AtbNQVBva
QVyB0e9E2rW7F1Ky26BJ8HXWEZ2q+/Er4Z/t06934tB5G7W7rUaRd2r/VCqp
qfq3k5ZVoVWEM2JrfXjgEoDgmgQVHIXukd+lYOMKehZVyEBqsYDh7WdGrEue
BgFZBP9a1SoUkB6C4k/8LNYbkDm5FM7Ub0a5rDLb5m2045c8lnLd0ndyK6Yi
BgkdZNeAiIKOAjJsbTbjm1s6ZYY93Hxq/tYyA/WNPHjvxwbMpgmiEHzzx75U
uf4eCyBjPPJwk8sYAWYYPcKWAmYV3x+6zke8mguOP483uFuHGm4TVHivqFrE
ej7Z01NcDqreyNwba+rr7s+C8ZelzBQpdH5QdZJuMfNPbqS8KINKVxAsPnMv
b3J641vFt5RpdR3xzejbZxj5DnitovUDnrktXTXLApmemPrLKROUUjykHqBD
lW7YGiY2dd0Y35Q6Bx05yirISpCaomcm0qIDY3N0YxfNy0tshw6PFJP0WdFC
/7FrQGztseUfF5FBWZpedsk/KoGhhUjHv5CHjBA8niWPREeqa2K5k+Kd5xpC
c2+PKl7zaxVZ33yNDqkh+bfrd74dtdAgD7L4e+bz/Ai28B0jYJ1ezra71+ut
rRRsa/T3SHUcuDbfsBH21iCwmO17IuOr20Dlv1i1ea4+QNrojn7R7XbVgKKC
1K7KTShwv5qD5gCNBHF+pFkXOM/PDN7NiGWBCAIfaJZE/Kvvdn+Zh+revEa7
DioRmAQ1IzeEtuSQEKxtZYZbKOxnYR/TBS4kMdl/Kb0gPEdqfy7Rinwn+x8E
tIJbEjTzOIKyZOJQBhs5mMNexMGi2dyBsBb9x1HpNOGT6ngx9hFkZMCYTr0q
ovigKMJP2FGhE+FJD7WMCQGrSoOlRHcSbrxYJnfYYXB1qoZpLrYgjAO0xzlA
VZqGy+e0dt29LW9vZjyrTxY/fuX/ChLN3AFroPFuHlQKRNd3ljD5LCbwhzoZ
GIG33VMiVh9rRAXWfs+vgU7KUaGsV87MQUIKlHzvuR2utScCV0YX61Y7tO1P
V6denJDehjTHhbFxENkvOO8Hw6043uLKwPkE5BivQxXxXLSBAsrkSJTn2C8p
jMTPzG2XVAZZwbbfHwM2Bi4KIzewseZifRK1FI5eYNmKbowDyDhlfAmhPQGa
mn/5v/pm4ukNUG5ja+ATZQHlOJu4u3XUezpg8RhPGFlKgb3x+OxEVig0wvlr
Op4tiF8xIXRgZ9Szz0kwvmveJalNhemZqotNCCvLK1XMMKedb2MiXEWZ/FE3
CW4GgyEw46ZENdk2syColoiHh5kwQE6f4PAZG91QGMuFm+oOJlb4zS5iEGhj
14NXDuJDATMNdi1ThU0Pa1EXByWcjPRg2U77k2W1cHYvCgb5Th6hZ7ozfdUA
tQ4uBidOGEOWTaQiQ7VsGJWVXqjXK2gTUXdr2w0Fi4oW/dSKPTDGqsmm833D
8bgdPWaLXcumtRN946EgSECLF5TEm8j89eFZXCQh6CvZ72wvhdg3DtuVyuEp
hH+87UM/mr4LurMf3F8kjyKioP5OHYZoZpcCCieagOZVdVpe+BGWMw+N1VhO
j/uWQOffNnBDpcZoT/TTwmZzy9sZ8AlNU10VzLa91CTTHEhOQh1XExUVVEas
SHahKqVzhlmNpfBw+F2kjrTBm8hcSAjgOlb5zLr5EXG6PFHXwXnqGO6nuXzR
ng9GFG+aHJKj3Cvs4BM9MOLSnAhBh0IqPN1TWha6GR4GEcyRcmW4A5zhusDb
LWI9Qi8OwgkRozmNzcRJPeqtUpffVV9wGG/cXUj96+MG+OSyNFgJaoyeEcMs
ZfgVBc2GBm7dRM+rzxmBVbRKfHYHySir3paHuuCGgI6+S2HfcmAuTHCblQWl
yQAKK3MwiruZtQRyEaewjjDz5MD/3oGOFgjjn4h1FvVO19bPz/K+4CXCcewo
ly/d/jbg7WjvPDHtmwUlgspiWCQRH1NpK84UaZ7w6vG1f9BEpVKIOAd6hBnh
Glvi5oYV3VzO7QdIo0PyTfz2SLajo125LZ2zkazAAN0/ctHq6i3gO2BC2NQH
g2sU9cd4QLyvZCS0s/zo53d1EFIexdp92PIZHrt8auUE23DzbCPovo+2yjrz
uBXvhRZvm0ev2Flxbx4dMQVsEpgpgR49z0TZ3sbwSXGE/vX+Og53A5x/m5s7
NjsXH14tiZ9Far2C5Smc/BWiZpK4sLSyhfKqDHKIjSJ5ACmuBtcu9FVSDdiv
wgGqcrJ0MJ+oaP86hvTVApcnC3pZVXu1U78XzJk6Lcw8+DlvFB1oZuoZTRUD
j5dZajPNef2e7w3C2ADIBFE6MlzLAAKSV0Li+AYYOuJ20YMbJNDBJvpNN8ZV
WtnDjrP1JLRNORZXCH1wwrC0RrWnciQHP7pJw1uwRJINzWHikQSVe9n3uwC1
NCXz8FOd99o2kFaKKUq639x6oRysx7Wcbw8KZZd2s+cvY2Ck7KbbBcjg4PB3
caGUQZgJzjDw+qTstd9Tx1VVf5nlGRcxRU6VWaRzrdZ+fXWr0Xj6G2bE/oEG
yOlFar6FYuD4XWh1QOnkFjoCW7bvsy/XKZf3RsfswSyxKObzF6Wt7ZJ5/41R
ICykWtocXM3spnKHMpIzhN0TsgckHRe3QZRSEzbl97w10qd516RU8BPbLx9u
PNahSP2zaz7dEbd47jtrAGws+Szgm8AVUWV5gC7nA7eWTxdI6A7q7MxvUqsM
3LwmLG59SJzYYvOXQC+uDyWGZyvw8S6tJBsSoViCoH/SVn4QfXqEibccauci
+60R4Iyzl7WpI2Ip4qqG+g7nlw2QYjSwqU0LduMC55S8DZ5M32SI2FTyCqQp
hqDeoFAvtMch8CUVv9tpg+MCnAFi7IkUSSVAAS+/dvbRUM5f6WdXNcPkimOA
nl7bbpKnGz+L3sUxTvLz3fhsagin6pJpRpPChNvJ+hAUadyUoTAzE5eFF9Xl
Q+enHR6WocM1rUFdccHA/5TV11pO6of1CVsEtxo8eHcQc/IuuC7BJqzg1RoW
42JYSsUy2gvt4PpsBngvuLVL+jYWvY98m5YJ6kpW7WAvlxsZFvMZq6af/5WP
ts/jZ4iX2gajq3Jz2tGKoSWO48Jwz/H6uTVqOtVkPuAm1HJsVeOLT2nVigh3
sXMKEv40BY5YDFklEzxfQ5xHGeSIxqyW7W8HgctSWPDvDOuz3lDJUH3lNBsF
qBwZAkf7XtQc8f92fstE3MwpXGCIc/4/9wkUQL4lrO1BdIPU62VgEwalYNo/
uUCWj6x2EwO/n4tjB/NaOlbbED8wWlCzaI54G/6Yvkud41PtzKLpX6PgCMNF
Hp17hntTV3IVwoL0rujSbP5RFvbfIqpoGKAvFRaIQ6nfCjRnvgCRF9aUNHM8
9srcSbgV7+Z2HXOsnhy60jok72CtLOtWAn+z3aE/v5eV87nXC6IeL/Uq2kdG
lAtYejHxiqTYc98999t7XKTa+XQNpptEwGtm7OSi3UO1pWKWpr5NVydp1G3A
zI/wpKJ9Op7pXcGrcVED+25tR7MKO2i0CsPIIMD4+LffY2EGWdOgs3t3Uuj6
OXrNDJ+6pKKTm8IARbkfsmCTMkICFNPnyTV58KdXSc4jnGxHdQljPwy76+zS
p7kiPMDhOEgyAfL2xW7tlgIdGWBc4v+brjmvGuQxOMm6su4pqYW0ZFuTrQ/8
NsizPsDnbcL1Ph/Wi4G3w5fWQBPQ4GGGrgF3iElSIPd/ZvlEiL5AXpbJ8pw9
E5XPJXBwt1ucPtpvvonBLQikb0FhKwAYc/buY6mgcwcDDoe7+/dIXOWzdxC8
fFrRbYUANnmb07CfrRjEFFmMuNi8FyBz4av9ngbdcAD/RnxKIu+soHQU6yZj
eoK8J5//3vzOYX3sEJ5GtJPkzYpY6uIP9mzzzboKly29Ud7eD6T+rNXLzUlo
9eJN8WQYWwERlITm1bffuBMV0vvFjbaj2GaA6BiWvoI0yCyn1uZIhIk7qq3M
6/JLN2Z7e+hZosa8s2FG4sYRhpcZxOKHN3Jj4eEXTftlUmnc5KSUzEP63IFw
6JQMsedfCGRQ+Kzja9aSrk07BTCtt0uNGG0EDo944qaBlCeea0VdfctYsqga
sdoVuDuVXti0ZBIkH/IAPJUd0wqOfa9/M4jdRGE8E5n3Ik7162KRrRTDAxUY
lEClHxksSjVpmt7fHOFO4QYGYF6VemukvBIjWUm5hsr3I4RC+o3Vb0uKF88d
zySFhgytQVk7i6ztTGYG2Q1aDXkwyGNFNBvTLjtKgCx9OmGrcDEiKlkjPuD8
Xaunk3V+OUjadXW3teBCL1dUmsGur0WwZuZp3QXrXehik+QDXEy2nx5xkRoa
BzN89+faK0CFu7zpPH0QNQHqSB8WRRlm/Jx3BhId967Lot/OOgj33ivfe707
nFXGBBRH4YISfP0u3s5phscxRr8jGWieqKf0/Igy1zuVrWH00ElsBimCudys
AP9YYKeFEOhcTgTpCZtLMkE5ZbG2D/n6UN6NvCQXnkqVfhqMTKAwGjvSFZXP
ZnaoFfZaNj07wdgDSgm0rcexGMtw5xO/dvLubZN8v5TsN4azyE3pCxmbKefW
n2u+kZMDuh9d6nKuJ0/wN/GStp6libbkovWSbGRLlILtHuXOrh3obd2oZNvd
f2nJKBbP+i852bJXnhCw0UNsoqVEr1qzNVn1gruIe5cmn8iM7citfTOsI85b
bRD+aVhlJac0jdH0FJoBVR1IiFfWWGbMRZusnDE+N02pyH9unjjpbJq96f7E
zskPNnWwSmXn3DnqWvncxuAlbsIR51a48ckTuaqBdnjBPWcfOBzjQyXegRxp
+xI+WVtrhn8mVjIJFRnYAn19OMUqNEzxrOz4JbnAfYdfAzqVrFXFk5Yevboh
GeNHaIoixqmfTkH5q4elLeO7EMaAtT8wDSoToY28U44KwlwVrMnEl8OBWXlJ
RjrbDaJCI3Qtis1YRp9HjdtOQMYWclqDKdakXETm7Rm/0xWSD7HPjDgd7aSF
wizKkHlDWfGA5BBYf14dWYiCSD//ZY39A4jy8OhoSrhHj/YKck/ryzyrxpzo
of4QJUe7nSacNz7GppqNRPtw0gucmuBrHRHQcwdKtp3PYe4s0fimTLQk0qCA
nWXAmlKm853pZ2FTT4tvqH/epQifwwxc9IlS1RM9pv1E9WXldtNcQ47DUmbq
GzaTsoUI+SVJlxYvybFAc/gNJuI2PCwOGNKtR3T9LIFt1ZB4WcyH0iWt7hSX
vB0E2n6BYqKq1F9TVvprPWT+PwQMFs5z8PTpY1sxyx/go56bJHga4iGsrOhz
VcBQYHqJfUaP07l07EKxMsVlVzJ+hjj8QKeyvs2YtZGFYUybst3S075QOFm4
UYLjBNVAXtuOqUav7xqH2IGOLo1eG1A5qrbOJpWFbIzNEopb/SAeWfNWLXcP
DVW2q4F5q83ii7hmUbVSUEZQVVqffxIg+uuHwZXT9ApsPnIDoDM8IQghzr9c
9S4UGUcH761z3uzLFTR+sIuNX5G8uj6bVFrwyTrFVz7P03ha1NEngmwda9xI
rGtRL/WDsjnCNwfLLYHA2kSvSrOvsqhHzmo+4sQjtNj1b9kAB1nE76F2ODUw
lCN/vpYbhqNXobHgNHYoHHhGeqBHiRGdSRHOifHs7wD72lJotxn07i5gEwXK
dCc+MjyOqOX1Dpmsz9L5g5mETPzSuwUFIZr2YMVQDR1oozmnHZWtdWEjsgjS
wgAngblXg1BZH4S19wfZfFkg6zOyUruTK51FecACS3lxidzxZOvQZ+l22KWS
XtnPbJvYnoKmtOTbIPfqhPcg7qwuRixqHe4krQl3dR3sGYi74wPcMgTQMZru
M+Y/Z2Hmss/IrcYSrxqt/ptSkJyqrPjCly8cBFECO1pk6maQD1loQvrU07SY
E0pM7XcRpljy7cS5Mu9kc0nwQY+tlpyp9rBM/iCuneIGirFoHorsazKCBgXk
zx5QBg+rJm/K6vq/6//NdgD+QBgP27U70RjUyA8SL7jiJhmicw7CJKkwVFjC
yB2krTHhBWAZzy5ZcvOoA8fB2FihrdeJELd+YwPyntokqqHMWrpJGFlPw02S
HURK9s4HZCLOq+wgsQ2/eRZMop1xl4KuTo7ZHanLOvWiZfV/um+G0THR/QOq
gA/rBLFBVeoFnjciMA6JwOodbIBXdiF6+8t8A1Q8CjCHxX56cunmEV7+mjvE
5zjnIcMg8yHd7JBC9HLL2fKWXceAPPMkPZIig2Gmqo58yX+/2YEbFKo3YBgJ
H0SoOb6dTJx1AHv+8FBcR+tlqe15AuGn3pu3R8xQlIIpGoNxh1hxOcsXflcI
LRmr2HtY6KpBmCqtmxW2H7/2+u+d1399VFKOtZO8et9XIQeautc+IX6kT1xC
tNn8+UFfyr8jlBLoqFxXMbr2rIaXg4BAOJGim8PXwCunPosbIxa8rpn6TXRK
dnYgP75C5/NaP3StmKgA60L+/wRw6jUglSiE6wtqN+URZfiGKuYzsKg792xf
clbAKh3VVdrtslVEVowwMqD+f9Mh+QRvA6MKPGXms/t7Iogj4J39QRlIdsCu
xezz8alRD7478DHbAL5COymXU4J8bRxYe+6wMpRvxunCihk4T1dFSZntOp0u
mQvNgqQGj0FGDwS/5UlxYK6wKqUCjIjiJxV391oRf/iC9axzMw2RQXf92LMi
oJgpzXywox5edBrOyHG46vzLTNH4E9dXPcVd3N0VEn/VTsKEBK45APpk8f+F
oH9K6TwrlHn9jxVSXTYp6RlLT0si5b9nuKmnuN0lKGhX/rzVeoq+oux1CKtN
Gv4uiZu57hLkBq58SD1GKDdI4NOMrAJXH5Dqr76/9dW+7vM4Zo4+YUKH+M7H
FaI9kejY/hp98tPErdkuXShTJFcSUYyC4tw1s2vN2zNK95PaShSMxgfMwZDg
wVcNpH1fjXVdis4U25jaMZ6owk9CrolvnGQzAsw+hDoiwOpg22B5XgPArDlG
1tb9upZ9vnchLKO24+b4so2IiSBSaQi7AE0FyisRfAtvXchzCesDizshbdQQ
zuvmT0T8v/XvwY0sC9gcDbvyUfJPgrpUaWZZWs94gi2nmqprk6XQMcJcRvk7
rNqZB912fuJ8ZUPhGWktbwKyhrCDHc4eHxA5U7sLp3gL8o/HzrlzXs3yG39L
D4yMds1p07PZVVmOp0jd9f2pRlSV/G41mOmYlijbtCC9NQJ2KXDgHtsHxNHr
wStopTxsonLaS8xA6xCgeld21fX4fGM2b6HbIRN++P/jvgaAn9ADSqoixjd9
QwGknIePNiXWL7xG1tTxKGTQt2rjNm6VYVPEIzvl9YuQwobqK0N0MdfiQl8p
WIIZBBHjYICOiBd0/56JzAUOt9+wBia0RVq+r4yqxwtEWL5U8+eb3piBH83p
U+7FrTyT1Dk5FsfqN7Nmi4gclGU8W9yw6ZfPQfRsOp0gzCRZb43qNkKNkwXH
9TDmx8FJ1TOwaxaoAKWFGrQul063cW0wiWxSJEbTGc1wCYrqwCxoIUps3SWw
j6/+E1muiq+zN7WRzfzZcBrDdzrsuE4zsrCQS6XGAKlfNKMEP/hLHh5n3IkJ
31oAhMNmUxK5Rowj0qndpHp6whZ2wk07hYFv1/SWjAuesgHvszDWNFvDyhz+
RwYWtoZmHCNdPS7/yI0mSopepNaiZ+IXc+Hr4XfwOjkHvZrvLY6g+oYIE/sX
V2e7z+7oWTg0Nm7EwFTKT7eisJeEC/5H3922Ojkc4tbv4VGApc7VIdw0agJF
1IbAenZc5zNRhuBM/UdQ8Za6jvHvCU6EA2lqzIKsEBS1UU0fdqEE/S1eLPVQ
aCokGnLImTuzcVJQaany4DOvadnfMJP2X3TO2dpXdqPrP8IKL9ezASQnBWPj
5zSwvPAbCwU4hxiysq547rZ/q0ZaKPC29ebsr7XCCqkDlyWVn0MQ7xWc3cJe
6OP+JQKrWjqAuiV9dkAhTqoZJNPIEZlRqAmWg+IKidvvAnwPbhQvC8UBRh/7
nfRXtseSegUoNq7STQeGLU2GQF2r2GpXDHLvjrL3j4omdeOYWgZkxiYeaGio
2FdIeZrDVe70txRhbRYuK4LbFL/bCxiUgPwetc0Cfd2g6uCWi4rbAJ/53elG
cfvfGFNQYdKO/V5+2AXDBRqrMJrRr4hLBza643uraQfIMwrat7J/x+YzCvtd
9QGzIDvUlArPnh3RQDo1IBroZeTYkcCgGrIl/l7FyaswpT6YUN2eTJ5GkE2i
eipVBVMQOtWLUZ42V9xT9fnl0VcoaisjEnel0hqLAH3xSLlWOPBFvTMCvZ+M
dzDaJPxDVV0dWi5N3T/6yIsRIwzosnoturKONMX62aAzC33+l325OAalrmDy
nI/1D08wwPzyf1DAGm2MzaD2IDDwIGGaREtmUOJN5Yi9U8hO+Nve7Hg7Wyks
B6ZgF5dBXeWLimHSjD6UY1AM4S+yLE0/bcG/tTgVK1Z/UawIbekOpQk7RKnK
iz7V098Jg0aGQgkDXZSCR6EfsxqEFh5m0HodhEKERTWqBFLWQhep3GGkDnWK
Lri6zuGAYDOgKwGBdjKFm/7QG/vf+7NenjsOTCwzf5RPLEm9IBZymWIyn9yW
xlG2wVHczXZtSYdPn/BvS1LbenChu1hg8xqLISJYvpbq0rzk/slc5uNnAr5c
p9XLhVsZI+iyb+T7ZR1m/o38zZWQWlVVzmM/cxxph+XWl/3tUw+QP9Yr6m0u
E1TeTAGp5rjU+Anz7YGjEqB0BnZEu6KsOrYaQPZ7A6OYQpCM+lO6PUVgtV2d
5Wr88Ao90gVJvQfGnDgmWzCV5kX3T0FVbdEROIyqgy8zr/XY7SVTEKDrHmZQ
Tsb5y4a84Nx2nPlRVlhkoGLzOYWsHmeexbURpW8UsdYlsv3lTuGnOF/dcIRX
TfiBRe18yhr363KhIknXgVT9hT/TswP7eoQYfL4ZbyXmQs86NQt/AMeuKF+A
TWtB8+GOB4qhleNZwCisBy7wx/IGNo98wZrR0T4J6kY21JY9nqWBzjfA2gBQ
56LNZjY5NPGVLKV4CcVHNOMcMHxhTmRU6eRmyKe1pQDMYB96ZuQEo1ab6P5T
Ksn4U80eiUK85sHESVM74MURPzZtJrxdaLc9/gt3KnCgPxq5zjhfhczzhg1N
jSmMc9567SHGZ0h8/Y3g4+UF6ktmmy/hjv5HFX/EkjMb65fSc07rsJTOxAEW
Mro04Cmb7QcH32WFXey409lUqRCCScG5PK2i7IZVawnatW/OdqDhazF39iWG
Yh8DTXBco2Mn4Y3p/ISs+C2yq9OXmWnpd6faZSQHJzwfw8vo5liTl4R2r9tH
DaSFSecFaltc5GnFPxbufgHMlFzCLoT0oeVoQ5NSGapZ3Qm3CNovvutMq/+G
4EAP5OEqkZoowjuVEuXyCR8qfgfSgQzcYvoUsLIbP2TCJLMFkhOdssIchaMB
xxoDBQ0HAdZi+q6MBbNWIvEbjwSZuw+eedhPhtRIUklAdnldULXyr2flk5n+
572Ep5enkN9a2PPzSbr5wwBwCCklCwtBU570ocSTRmIJ6YCpoWXWrbUdh00d
F5ZxmYg4Wmw2j3HWr80JVMkdT9LjPvbxg75vH51JEnB2yd1uAZMHuhAVzIKG
VIX+SF/4elXEpbI1SpKvxBpaRIEeuN/xDgzd60npatfI6yTTwIqsGPU53clx
2AyWfQKYJl1VruvKSbTK2oWRAOOciYoQ4ZiIPIqCKS9icFxWoKXIsrBX2LyA
5ISrdKG3hDg8Vr3LRF/nR5Te5n1klOYBjrqsc5290Fhz/NnkmraEYyTgk38P
KPYfiZl0Qzt+mQg4wOcNlbQgpIxCjVmlYan3OLeA4TZbkb0b2iwCcPci8i1l
yi5mqs670BVLHX20BLNjVhQy6nDUsSZef5yAg2N1Pom2DqKu/TO1CS6yYc0p
xvkMAsBFMhUpFh6Zo4YMKO7/ue4ldtpJHbY9OCLVUbaGj8TXuOW8IX6fIWM2
ExCiiwqAjJEEaD98FyJpLgcaQQpEVjNx+WW2WgDdkSIUH3vJRB77oGKPk3YY
KAuv+Y4tY/cvPqyeihZV0lOllFjQ4I1rK6LzrIKPlVpwvrX1Wg++uPWxNHD1
kVGtas0dh5c1Nvr/tSy9HuNA+6mDoQZrBolh9R0k6USbqsKgyMvHvAzRpKju
5u8524O6/JqMaK/ZRCTg7ItCwYrRzicgn311WS3FzeAVYXbYF9ol5mYEF7rK
12D2HNe6nilrxWBrzGQKVHBQApPfLFsaLHyADfxWHldpG3BWP9XGPqVDveRt
XfjBjPkBuo373qJWrU2Jld9hVCIV2T8+7Ievva417FkbuiwGySGBCZkQWonX
lQfINBo3hb2tDFJBHnMjPeGabnSGjF+2uo2UDGoYnSStE28lyovpu6AWAHav
gMdN9l99VMr1oVXOitjwHHpaGEJE18Gy2wzQ042h/evKJk1t7p1c0PgDjm39
ksE6tVXvY+Qp1Vnr07Ki2rGEyLdvtwmRiksvzdNunGrF1kD2/8XmjhpGOjyY
Kg2WJ+PbqIycj4+2PYMwP0Px4DVvxz+/JSCe6xUKa6a+/P8UVR1dRCcUub8Z
bHpay+7D2XrcjM3yFjJ9QswD7mE8ryn47oxSgJin1cPbocppV7GyEkDN6WJC
U/3i4Hrufu26/9TB5cYEZEi9iDwCu6Q7mef5o4BAvM7joLOhjebb/MpIF1Aw
EVjkmezfbI7M3NQZ0m9JRFkG1G5+umcayUTGiVgQPIWW7qW6O19vSwsYXKjE
GPQPGTOi2FVu1n2CE9w2GnYDayVDis+Gxv8ClTswG+ooPuu5xXYanRMzKEsy
1EoFDT242YdGLuFC9cH1Hr59z36MlJNd/HbokM6W3K4CjRnp4D0/rytepVFL
g+N6wNDfq9MzbEPcIx+bLzaM/6P02hA1B1VOqQjkFl1d/K1IOhK67Ea6vsZE
Jb9asihBCuenEqS/PGaSgdhH110piMRdsqJYEH91LRLRgvRGr6zftqsaMB6h
sfwZUhnkVMZUU73cLuPhWGDcZzTT+PJcELdaD0rZiVmBQk/5pQP7WWsPHzVW
3XoMnpk13l7S/Wk91m0hTV09FWtGMagVeAk9/Joed0lu/J5LQPdl5TnMphD3
czJQ8d73arixEE0v3ZHXlUbJtDBdREPhg89DjIR6g+zLQg5qW0qyeFzgFMfQ
e8+xSt+O336D0CxBuRuLmfNOetWpOfNB63lFwAQl8mIBVnBj52j/EzNc3szY
hty0pqpmDf2mJ9SpxCLyT/1rL6KX+pCYYPOfW1TsEIcGUTqACG9wzcJFtWIC
sPpODVK5sC2GKph/GHdzy79hAYLSZcboEV2M2RDSEwf7y/QgSTrTtaYiTQDY
CezZ6YKAVsQEhtW0LxuSS5gudh8ytIQLT9tobraRVqPlkW8C6P0K+ZszMpBb
ixS6FJ7ZuGfR/A+VlGs/ygLvS0YPfBYC2nr2IId+diuUJbr7jcC+jI3zIIZL
BgSwUuWhggRVyX+YEzK2pxUT6c69PQWG3i9Tr6VnEF1vWCCven8xHovE1Vzl
Qbz1vFdKEqpDTASWYOZFfTkaSxM5bU+SAd9V227ZCoA2Y6iP52B4B7ZLlu2z
ziazVdh8z9RgdivspuzGM7psRWZ3uddueMZwQpltMhUFjVOfRoL+IdBafJTA
f+UcWte7xeDSRlfYfUQuqKB0ODfG4muUzEK1Wer2yUR/Lp+tCutddzlTpKoE
3ajlprSf87eznduBieA8lhjN8hl0wwa1UF0hQ0gzllN/OLiYxhZiI5EbWLNj
MVoBK6P5+Pc6ezq0/j3VpeSfEb7O0V0FmUr2GvUru7TJowX7P9Eo0moSm3tH
79hjTqTlRuu+pBJxj4FN8/nSWy9lFVKk43a7lYZ/V3Npuy1SW08dR7eDAHMW
9Udn6tYXK72H04hvKs7/YzJqPmwfHF7F4i3ew5ywjJkRhAXyA2Ilwi8ywci3
6eE5OHe70tFNxjoFnc51S+JMx5AQVRQHO4E3mjB0jp9t1Y3YwKGanQyuyaIt
F9Co/qKaSX7BHMMc2vgIof1jYeFlKpAzej1kto00qhPIp7J/NSNsuT1KbmfQ
AMMuVMLsHsuUZp9yYrJAPqFF0IA1PHcXO6xEJHfX056btx6t865l4+SCnHmA
VeKHnbMNGDon1tPvL6HwpJO57w7PfFD8Vg17l57ru7mfm5nvt7QhxxCGe/2b
avJYx0mScBZU8J7QT319oxYPKJvwidh4Z8fxiURh23WNnTROASH/lq5pqMUk
j7OrKRbr4U2MOs30P32nCIS8oTttRBICNlPzRSNjqY6xAtD8++jsQ48BSP/a
AaHflAiruTtxv5VktIHN/KDFY0Qn8gRdqJh8rKGl4zF6rZ4c5V58sxp7G6Y4
UbWrx4+0MNgOQLgM30Iy/tFCCb8qisejuCkMGyjANeGNlmCOnCUcKSskSUqA
oTDTFrUgNp2thBqJUNMLLNIgyM7KOi1uCpkAKrHqiTBpyMTFpk3LaD+Et7c4
Mbsq8T/uR2BPQsjdzoxsXDBPO3wAYB9olUZw9+tyY8b2FNp3FePJPPeveTdd
wNNE0AeMAv7E2QomdDz+jelSG6cWaJQFdXySJUKQOSUkSb1Py4ySsQ7kISO1
YrAYElINehoQCJ/JwTTQmecuZbqveWZQban72/09b2SXE0ZFxVUuu2738cYC
MLvZhf0ES6T5Eq5F3/I63vFfKThDA+rHEe64atvHyz88Y3pPaSMizLIu8hY2
wfBoAnXxbA8+x5jV/JzEWKy7c91HHWDwqbuZAINh919crBscMoA0cU4M9AfE
GMiOgIb9VhWvEx0IS6GlecuXjjcJLkHTJBed+k2CGKeJ6oOHYfBqslJgco9d
OmAgJYRlWFrky79EcL3Oc9nOAqxH4qh85ULOrp/vvBgLae77XPqBm85iPpEj
pTbLCOpdPSsU6+DMDz2awIUvkU0WsuO/UQVipzF9ZTcjbo84rqKcdVMv+xRr
Tmat95S9ys/Yr40BC5TqgHqN22g9PWH8vICeiEvP/27dVeG+wo5g1zq6+IjT
Wey4icb8j/Qvytg8Mn5CbSLZ/l01m+rxDdnchjVH1YHsQd2wGzuDEJjwys8G
l1n0/fjEcLOeEf2w7kUc93BxySXNOujn0m5k2LDBKvS+KAaUCi8EKQuUWn2B
1Dgy4e4BnDNB9djaRjs9HEcfvw6eNrNhIId7j6oe0G9VOb/WNyqFfL18SDOs
+xH9c0Y5vOGmz9s04fgKdPiel74Um4z9M1CuTRw+x5k/L+YvLWAe18Haswvz
LXgaktafxg0bBhVmWrhtoUCOEf+3ka2bDQOTsGu4a21bDeHj9aG+mV5yobIu
kXbLQxWF5kY3oPhVlJv619261l/7ucrB/e8KlsjXMTcVflYNULoh4PCe9mMT
kKsRROtb5cPWSVxqh0X5LPHan72E922PyqgZgYMgpmAdwJH1VScUy2Xcao5g
bNAVuQe02C3mcOZ7C903oMiE0FHmuz0Qyw2lzbMycCU3LM5tCi/Crt+TTAlq
KH70roAaFOJaZ30ohIfWGoXHWjx1YHJhwvNCxTEkRyMrEYfW42FTpJSpJgms
H/8cIPNRhjUr0LKao1HMhW5HtIcqHgvKLG4BOBPbWqXFm8hJTVyikdENtany
T8zXG1AtrEnDeuFDV5b+ToJYre9M8rd2p+d+VnFrMzE/7BzDiaSDQy6KCuJa
UftSwRrXK3M++CPSc7P3sdFFfcGzgFJW11IKFPV+bh+MNVpTm1YuXMrdvZHn
h1nC+oaaSxQssDRfjkbS9WyqlZe62DT8Q5rUTY8KZXCh+yKgnzPWybETVsz7
tJL1nE6MBVd1Zv4Vg5RnLNJMGf21GP71CFBAgnWzm5mWaEvLaBVepfBOpThG
AZlfQwGx0lk5zP7IG2RuxEb1aK0X8UolIQ925C7O1DlTbh61z7kv5ipIs+C8
axzhSKj6PjMobMHXr481S0ZsZPK5PjxPLu2ZkXaV0Sd99qewDbfBXossud9f
ACZFa2YGQ/lJLuVVzMH/TGksUolP22ohgnNoAjnFC8v4nUDwkBzEORd2VDdX
zbIOF9bS8pf2Z5I56sOb/1IzrUCMnUkpecj9MwFkOkhBjnxXGXVCzPQrxnwI
nTBDZmnUL/JFYS+kBt3dUBWXpTIBJJu/HU+uSMdxFG6Ns3UnOXSI28zE3bYi
n+k5FUgOhUj9gZyA6z7/lYAniOK1Mzi26dUmPrF/ggAvQSJ1IPtXn5sUW8yc
9Wo25DzhRBFc4If+NyPTAz4blCyArwiTZeYed400qdcI1SRau3ijv13dLSVh
OxMp2ONw/Dlhe+uudopbsIsXBE4Q6NMbHgDGfN47P0G38+ZdaJWNZuBtJwMi
5O7BS5TmrpVLPKwQNIet8B8YZ8FEoQPZ+wW3DGGy8KR4VZJ9SNuoucJhNlVp
4sRwxnL/6loim0AU1wB8/gGdjseBNHr8nGpoTvX/soMIF98mQO60MPuOgO0a
pR6pSWM2hMUur4OjKtPvVJe0bTnDUwu9ETB42ef1IIAGEU5CxUqm5FVsu2L8
uSmvyM+50SHhQQpm0Pi2BtL6ADtefEd6/5HTtK0XWVDmuHZ6J1vVr3Mz+CP+
hSYy4xdBqMkvHgwNr2wcv1Byc0aWG6DM3W6JZOVkwNqaqgXeYOXoK2iqwYrt
cXLLy7DCD7YF6zmHVq+5pLwvqZan1Q3npZomotudjjV4u35zSVPlOAvYbId/
Pv7152ZjeeSuCQ5qnaBkSOUxgk+m9e0+7g/mQI+U3gWUrOmBfTF1mwxM80IB
rv86ROiM5W5X0skmAafvyFPnuO/XdttTp6lJDNgsVT4um7aguEcwlS5MvgDt
O0SDN+nSoZRPWjUd7MoaZbWYPn94jhdNNJHy0MP4Hz7CSOO8k7wo0xR6P/fc
nx1zdxBwd9B/tYSg7bOndudbv1/fwIur2ycb5dkhLgto8NbvjldXsaemO4mo
YpQVuO6VSWzTE8hehUWLEzI7GP3n2hO2rtokBHOLfQxuR69xRkjLRdNIGSRD
0oA7D50O8QkpQO5sEoYRE9XASN+ZvWO2a4uysI0GOE83ikX4gLw/z4J10QdJ
AmEY00mtkFkixXu2NXGwXuBipKvR/et5N6BlkmDvqRSzqXwRedwlqp0D+wKX
/8j2G5bdo2cPFz0xnQzdATjE2/vZ6ZUAM+Re1MyiidQPSEKTY3bw5g5eomBb
Pmv9jNe0ARQFaMT/+okw618lYn7IVWythkwwQttXuLKthMarYl7F97GxjmYz
3ec4FPOEc0KF8Ffbd/lHH0CDH+yGldDtWxZaLElKGF+py/JvcGD7BXs9py0M
wwYp4JE7UZk0kW3XexRMYHsD6DtG11cEPV9QpGT8gxEU9ZhsklU71oHmSYvQ
1ps3/ww3nItniUWX7yZBMGSJLvEyLJOH7o1KYHejsWVcTn4FAJ8z4HqbaCV+
qwOfwzHsnEFZlj66MajjtvHiWzY810HCTJLISxgDL+hL2dEpFE4Zf0R9qSNv
fUCZ29v76zykORNB6rjf0i37OF96S4Yj6x8enz+Qu+s0TT80qHmwDQtRJTF2
ASxDDCLTB+yaFd5CLAKYhUSg1j4atq/ja5H/OR23KblpA17LvXBairkj0BE6
52P9Y271D1VsPmgBvdZMfGdmTXcu4Bft8/rIxliI3qIKbHLIfgL3//z4RowY
jpcARNv6sv68s9R/WyjDUuO09JRAjuO/tvCGvNXYvIEA3FAAc7pOq6H4ZG7s
eosKQnHh+bCGNOJwDDJKGK+ynV53IqY5/cynuAb0pvhXj61eMj5cpPwUVS6p
rK9jT/j85e8g2kxOtEfq7A1+qyGaoxKX9ZHRXN9e2JDGaTB5D2agO5hIwzXq
ubtB2QFEXnmkm8PGrMEMCXBm4Ov9XaaBi++Dh18fJW3V8bm7pB+3DFr7cvu5
4RQA+WXQQw6n2FWLvCUCDcaPIBosv6DtfU1DxyaTczmd9eHAJq9/k84waCj7
WDItjRdyFNe7Ds/icFuDR+eXXSY5TWtXObhiv1p3JlAQpA+a530CrH8fIc8T
aZbORRD4ZgOrMOmR4fnN6ER8AHqMCbiYZtYWkszndpv1cNt9MeP01uE+xjiT
/Ft4N9T2mv/6YX7j5RXhkZ43UXY11/fT5GNcJhRpJc0Bf65mGEv/YERZHgqB
GeaPP5btzRCOeq4XNaFe1VyhebSrAFCj3Fv8xJcTvk+fFdtYuFSJ4feAytQ6
B2h3FiS1L3xEB6syFLQGdpqdDR/HpKV6psvXCBv+m+GphYzPS581YVUWHTtQ
wtLPqoDYACICJdeKkv6d0+1D9DRVqy/5owYZj9tlMinoRDcqIJQj6PcVxFI4
QdFhpmrI1fVCj0Hm7pmDQ4jUwNiICi+RzTlT9zXwOp0NMC8kSWmmRAVxzrac
zn30mHquUjY2ElQBP9ps/tiRcnaIR0vTsyydQ+Ypwf4Rr7povSVq3DRAQ+xY
aCjko6iID3+U6Luk7bZIyPWMDMB6RRetBa55EK0CppOIMdQIEfy7HcG2ZhF3
tYiGOgGk9oZ+32BSUbaEWom8XKsGLLUq+1gNxEXpCfDmCg+pXsbK2w7gMx9V
IORnridXaqdrEsZHSoIFDc0/oTUPR7UlzKiciCYqMGlO0p/3egTfAluqyTjk
tWzXgjMkxQvE756S3HRmR/19jApIEUwXXxLeqGh05iAMUFUaWXHZ78g14ovD
Mn0LsIruQ29As92MICtO9zY+idSQM8dMJfWywtkukkelBy30lkEK8hYycAHh
2edlNNJjSXunBM19eVQtw4as2iF0n7EmTDgcfGSk9SsQ97rCS6qt2JS6cSaM
tkPHsTs7sSq6C3k9E/CyeOi7ujTuPyJTRjM1FP/qkSeZ8mcqFSXwWPwmCGgh
+r+BBj/lQTm3gip+fRyZXXB2P0InGnJBPTW0OKSLhlVZFWr6yAnE2E0xzKV9
GmBdKN8NhXymha2F0/CU+SQBYE62aAjmZzxjZ9L2uayMMFpdVk7NXWavVV71
Mc1svONhKYtN08qdubVxAqlB9EuwN0iFaHulI2H2rg6kGgLBYTUlilGxVPZt
krl11mFtUqj0KzZ08Rex4C4yZeyYkkCrFsN6MNL24Euj8JTpc+FG63+C9A97
MS2NMw4+KcOYt2PF9o8Eevbz65+WTBSZGhcy5Uuh45r1d1bZHrjNT2QruFMX
F1rCRRSDVv9o47yomjYIwDy9LYm8DNTV+2tTwSZ07/58nU2Wq8bqN5NjvDqL
iT75cO9yhN+meQjOdgjLGm//Li28KZ61PG1z9lNUPL9769dgxVOFg1WDUGx/
e6lUxxAsGLTO61XNYILTWeCdTGG+8VYOBVOGTyHqp6ht/KxJAgfApT1aiQRr
dhK8RO99Sz3NFo4eQROSsEExxt8tHhnMnfjBVj7xuXm+ItFxHgmlDa1KwPdM
lxVcc37TOPc8nusKr/aWel2/f6m4RsVTZfI8qMi9mCBqjLsVqxExzoPPos3U
0JGp+WdANWIs2aKanb5JaiYzbW+0iK4Kv4eyiM1149Pp+kxd0khwKxHC6zIV
4BMUSQ2mY2QP0k0s3dBvywvX/ZiOGOB/g/v5DaoiMa3eW7TYordgKwIYqfJB
Mn7zO9xVoAKWp8HiTOt+U0a+IoMc5UEU/tHSEoLbRE/VsY/MklbD4WiZQ+Vh
E8twi2Rh5++RExU0Ju7sR/D8+8uN7AQ0Ob8IuNQeelOoWbykW3tcV5u7HQku
YGxF1I8lLOQ6hTMswnvGUHmVekp/O3izucEt9spwZmrsMsZSsEXgYp124GH+
RQO9qWsrlTQOUCY+9tOxSjur2KeiFyi7FnlMCzNfZOSqcVgy434JDT7VhaOW
xwJPWJv3Vvr5oqJ452aDEDBLkg7CQKTjSlKQR5+Tu99HoiUQGnStyfZFKhYz
LAR2syAW6BBDcmrCxzjMFTXNGR8NNDc7OqbSOJ2b7FAcv6yGpXmul93XGNFE
x29E0Og1emXLahoR65DpcZURGLuLG/8ydZtZ4UQY09MPlRSzbmVyDxh2gOtk
FP+MUQIaBvy/OAQ4NxFdb1nE2/ny94hxf5yMhGwwO77uslK/zuaBj5EHXKOn
rEwIA1jNyuQN7w2nx95+x109j2CXmAOLV1lfJtonVO/LE7G8CHCXyFgxjETl
X+MyEmDzOxoHBfIi8T5qCXKwVV8Fpzhv0YkCcSvEMWy722IJcJy3/mze4CYz
prvncGAqDWzOGvGVuprNoPE0mxgC38B7BRNdjLT9Ngfe9gH3256XMOoqY5le
rZVMqf+2YmqjgKTrRLpCliGughMoAYYMDZn23PGjf0i16QFEGvb68dWJ+ymj
+720H/3KM3DnQTYhzyOj0lZZGPgAYoTFXLtbdk2xqhoU7r2Cplprp8vro7Y+
YU4icym00TaKMlmUJuj726BLhJeIkb/hLrM/mT+jy/9gDy9f3wPD1C62vC1l
qnEsnbxa84Zl5lBfAXp7LeTWGjB83zze2N9eIMwsdPSZ7lbmJiI+lFdb9Sdx
aIY5p82OKb7ZtfeO1XWi3aCRs7gt1iaTWxT+oyah2mNW4AqUNQgN7C5fBsrG
Jx6bPoI3G8thj0KI+iMdB3CGUtAYk2uCDdqIgaS0K/QBQlcNfQRxSNpsd3Mz
Ews0MKLYxaCt1HPQORDDrNoJJ183a3ZQ9lCviDxoOg9T/rI2ClPAYmS1X6E2
SDcKXu8cMjOFzKQAhZk0Cx+3VWI7aLYS8SQ/I9ipaot+7Aqa+vF5g6hZFbKM
1fvIIcCjJfMYUH2vDvGPJ2GwNCJfh2euFvFaAtlwPGLywDwjdE4yFlftkHTU
olVGVJJdtYAcB1n/S9rWIyexuGi5mKhefL5/VJbKDbOE2btqyaMmdSWIwCpH
AyLC0eiHcYqn4SfcL+5cIpiZ7RXAz21QT+3WXlgor8lq2gkkVH5OSfPWE/YS
h+f0YkNNVfO21cn/s27r1z8u3IwKCSQDXXVgI+XYk+Riwr5XS+UeHoS7s91G
6mioesXxvLTTbm6DUkPSjxDpqA2nZI9WpiBoOXgY9S9kXjKkC7uRm2V/vt5F
g1yH5QYo9lFe5wit4OsOeM5qEqFFnYB4n1gVlm3QMFvWI1Z2O43gQvTbejuc
mI/ur2mtLJ+k5ZpMto+im7Q/WftkFZN/WFE42b066ntwyzF3uKfdV/psSEkz
guNNpMr53X6r0dwN1XWPu/SRU6M5bmWuynm4XZqA8nYIoDJq9zfejXjgd7Fu
2siwNzlUWb3zBVGvW7R4Hsz944vBYdngabvqomOSAKqicz8nzeaZqS41uV43
2tQO46gFF1kxPMpFudBO5PQxVAnu6x/nEoKLdTHKqu05CeO1f40vw1aCCPl0
aWtVYlAeirms2jSzBKxihtUzVor49wHUwq+Ri7eaO6p0QqMMlKvwGdADb7PR
4bOnIksP+sMfwYgFw8Ayitv+9RmhEq6h8f+0rEgje1phxlb8kViM9i7jqO8J
EDgbSbIcgnNMMfWV+0tWfQOIz1/wuKqNW4+zy5ZoJJ7QBaYTJGKTvS+SoF0H
ArOjwbHS0sTLFypuPQNuTc69hBl4k0D6Fai64dmTlXt49T1prqYnuJ8RcOnD
L1vyn+8xOF70pFMmHZsvZMCA+i4XczeHWoBEQ/JyBjlwEwZVW4VqiOS8hp6P
g0pLsQGddKLxUY/5qjGrlQrnUqbVWJgUJjvOaWEQuCFLV5VG9wn58gfdk1jA
vjUEV9VfHWWnlUitymGn3sra79ybPxkryDt8yPrDZVnaWjrPMbDpu50hh5Dc
H1tJqE90WoDzW3nxJiy6/epT6evXvhBqUwvLqmpNXg+hE0bmIhAnaNhB7EBY
u85xzTeZedu6idDStXSqzPk9ssLDpY3OBhOtKjaN7H725IHAgAnFkiuDpUXe
LVBpc8fqzQIydUqqwXFras+fnwLaFn82d4pVb8Jc4paHFN/cYkmNNI+/er6H
DLypf1AlX0AI/9SkPAzWJokEMnUJqV3yV8LlzEWp2JPC/iKpQeB7YCvsihdZ
2O+CZ4Q/pjV1fxzpYyLf5rkDw4Q2VmUgRrV+dG9Djw1jjfhDtMCIr7Lqcvmc
vgJfmI1L3TY9E5tq2TuK7ewufFC8In5mHCH2HBKQSfQTWGsXJ0OdWyHEI8MR
0lSybvf4v8Ca3kXsDANemrV4n7UKqJOznLJzfVJeRzYkwWI6HMmWQiGQP687
OJIzm1InOMyThBrGZV46tXaztEIdbqRfl1UjloRjBOdKLrx4yV7YTHvQEHSY
0xZ4nSrEcvZFoo1U3SnVisH6acvy8JbK3v+N/skDR7LBPq+967O7axA/C+Nk
WU/O/qEeif+n+p0PNC18oRuTSBEwhphtrSa53HHWM5Wj488uFH+crLsLfp63
PilOtbR70h/vfdZiwaw9ho3u/vGmpxUJRsNB4ZUmVy7CXnHSd56722nK6gyj
DsHiFnxU3zfihm+LcWOC9wZW4vdxyD95IORGFaLbPQByfDL0GSc+kGLIt+fQ
7EHN8il69fXdFks5bYh3tzW5biO43dyMhIV0PIvGPQ88UStqRJ5maMH8tlLt
R7t6JdNEEsfejaJIheGzw8UzZKRGolyFLhJIWkMnEJxhfK+nEcHyKcep8QWK
IyCz65TGr7sUYeLMoNLbLRC3T5kM2H0p5O0jdlfgXKTrkzZIuubKyYdIAA+z
OWUVUZAfumCNdkdN5eAeDx8RpMMdLhY9DbZEYOvp0JBfZY7HXWjdJarAWQbe
xsKo02kKRCohmZoJrCVue6kXTGLxsSQbmEK7M2gFW0yiBvtcgpPz8gVKWWkb
ARp2oGJODn3Z0hquIc7BA/ulVvu/IHOP/1nfu0dj/D4s0ISh3NfRncDji3Ak
xEC8+XRPqa3Q3tH/syF25JPNl4TW55Q0BtI1q8dgJt+nfT+agirxC1y7wB5w
pJeL6Bp8qhA5jkM24QSs2SPWkFrZZHuCG+evDLMjSv5z6rSgVyGFn1j7itdW
P/0GN1GFB9CUQsCwmPgj7QWlYkTC1D7GSGMgT4tU5xqnHSad4+nUUGZWqxU9
cVERTI0D+CvMUM5t1yUju99YgckGJUj/1uagBKs3cv9wwVYvxdA30qiCYtRd
vQo1FqeqZE4mN6Q7vSMJqtXsS0YYcOgpT8rDCO3lejWVkIlvObIt+yYyONg0
CCRag7rPfL4VQzW5A1mENLFbv7JoMpjqLk20nDWmCKfad21ChAn+fANFgmKf
jqymtlfg/MG3QZVKuGlwEQ3eBbmvbf47yxAyHg/0LiX5VQKdIeBJ2z1YfYKY
q2tn2b0MTCVtR4ZKewwGwus3cL7SPDUpDuqISYWFm7A9RBuoCtrNY7h9S2Yt
U8EuYHiOIk2+owuZvuZ5wdkkUQZ59DZvnsN7bo9ZSwPWR1KD/LCO1ODF+5vs
QHA4FRHLO3ZQn1GXDBj6mtc1hWr6W1b0Mw4x1MyTg02ZVQ7wmn8ccwzZIHBy
cP68X0xjmhHT0Fk+Yw7ZgQfNgqQgHuuknrjNrtU2fk7GA2SMdTosGDknatja
edSUAFu4Yj3dFdj79VESXz6ipzPzKNbll8EiK5FFEC8UlxjQ3fLOo2KOxuDj
Uh6xTIKn/0otiEa5H6xFdWuE2B5eob4EwQfDSCmPqc6ZsRSCA3qrHWuI8Obo
uS3FU5J9Aka0Mka4NSojP1fZYrEdymUyoL2WeFeVQTDbPqx+77+zb6VCbHca
QQgCc5PK6ZUrY+AgeA3py4hrkwL9M9enjKY4x7GSKcXW2cg5dYOOqkZ0CAY0
xNfdy1DJ3x7bn9QyH+tfRF3G7kKQzmsREniuzC0sf26sh/T139Jud8b1Dr0r
4DFjecZ8IvlXQNOseNdAOrdCuJcLrwKyGnD+kavnBHyrYeHl/KXZnY+/x/PA
/c2hUhB6SrO6ZDXIoUpakJHGKBQjexIuA6KtvH/QwkzNpLmunKRNeG0WgA5a
5jmurU45Kpy3gAcaSZo3WnxILB5B2BsDbbIUz4N7H5FkRufLQzYt7YjpoT14
VuPppRTdskckuT/gkV6ll4wVKr/OPE0QBXTyiM+ha5Nk9hI+H/EBzEcoC2rs
Qk41HTX0su60adjoivWJnd8aPuXA7cMoea0e3z7eX5LOgcfBk3E6F/yI3nWJ
pZkcmAXcVyLOi6TtRiedCotN6yhBUlBwl4rY2ZWuVPu/FXQU/+0ptJsEMi55
sbohEZJSXq0gqBzHnbruh26vWMbsx42i50p6rQkgaiMS3zZmoBwzg3kRr+Zw
OMfVYIH1PLe6jLPp3dWsQ9KDHmeQ3cPLY9KNezKhRk72s4Pgb+I7TlTfbeYl
vOt3ILNpile2F85PGAmMevp3ODDj0BmQtOvdGnED2wOGCFwCL2zJLFyoHRBZ
n9QcDHdvq6uO50WqgsBr9CbcBQBW3W5LFtK/Xe74+2khXbMYlVsho3uS4+nh
9u+jPQxRNz/ANk+lBZ4Az28jUImu4yuKQwJ7e6conTq/SfyzfsMIO4Sok74p
wfh63UjyM0iDdNeY8LBUtXjI/UYTpftgkJ1Qn5kJFS89tWbeZuJ3p6WdVrI0
FSGkp6sXHD/5VtAr8WUMkm/fCBYmAkHcELydKt1SMzvVQNJ7XgdlOyY7yhHg
BH4+/YEhLtI/Yvhm2ljhhFbzuwW4Q9MGKh9pk0lE0T3Es2JXRBfZorF7x0OB
ALzJadpDeEbjq75AtnQ6tJLDVPjoOIwOWmu70tn9yzJ/h6ttmOj91FWZLrBn
0gZhx9GeCaPcHwhl4rofAgZcP3FNW1LzYG+JCD3VPDCurypQ4Mb8IPmaxjWa
5jBSYLHhNgTXSb3mZKGMsBN24nhNc9ahJNimfrnbolWKEhc7oCFSnD+nHQUZ
AcTnz057UBm1XjLiunCcBJEo/MyDEPIKQWsSEj9yCUG27wPz9mgnDlVxoWL1
Cw0/4icm1XbMflbXpQA7PKPeLJHBZSELB8c47uV/8dCn25/8yAJlxfCJ2TS7
RppdQ2M0kNlqk4AeK4oBHV9pEbKdK0me5bAaBEN5eje1EopWVKvouyuVa68q
Ab8A7z+WtQpNlHLMeO3uFqWST5axaPviZnl16BlFCkLd6Wb7Ml3i381ZUsxU
aDst+NUNpdHTpE0qJD56nfuA9TNxTZn0DAwqGyPoMavpGoHaRi688rezN8pi
WgkeLe/bkYykLAAwbyW8vOlmQDUOZwGct0SeKeGfZvKlJu5fTw2K9DMdyjyT
dGja8TFWCOvcyZVIPd+msTGtjpFT8VgziUWNjee6/zURAxtrEC1Hcfzskpg4
DjaEvgXR7cItWaD6m/bFVthXxhC+BywLyRcRkEL6feags0sKomTEpJ/gP0Ye
PRAChaYyoe1emoUPekKC3/njeAWUemZJ/Z2nPdaWAVzzvPTsdCy1U8P3GJjc
u6kBFE0/mlPaBKlvRrBSmoGM9CuUrf0g6DjF9w8JFrMU/OGbUuPSuxw4Vtw9
vTNbdQhRFigHC9Cm1Tr5imvoWpWx7EbaIS0HcHIJNxTfrpzx9BazfUo9flMn
LpVrqDT+lvuHTRJQHW57aqosCkihmGTjOx73ZJBjYbd4ZZjrsUfLGOSpbfel
XMFgAhjNQ+L2ZSr3nT7F1dcBl2dRtJ1KrnSMKLplos5GdFK48jlHwOFylHls
4nXqolBoMifHiFXsxQOBJvjn/m40+uqG7F1V9BDRk1wAfS0qDrPVonDQuRZ3
Yp8xvLnV2in6+Pkq8OzlCIX/GL40wbfkGg2t4XdALxCcwhqumx+5eIs4j00f
aCdUd/5Dh6ElmLLSLV4E2fVyyTMPj9FAUSrZbFgo1d6z1HJw7yqOCAxF0a0K
16mUbkFN3dZIX1p3mkL91WUjq0z3Zo+fRqmHN0FQ53MSggLWdXIe2bHpqJUc
ASowtnlUDkT3hqpR0yfVewoajfaH09krC8DoOqF0zC4jf5YfjwjmPMEh+igK
Frtb0E7Oo7XiPN2rX4/BhnEXT/3gY3upQar5Jftw9BxA+BFhzjwnozdGW2jf
BJU2s8NCoGW5Wi90T7NF2Yq/7B2gygGUuAhdXgChJnV0rDDeRCet7hgM37YH
zDyHsQK/NiaTO/yYpzCgCjZtE5WVP+GDl7R04Z/txholAVbEBJxWaFZG5hU8
6qeMJsRA9g/F6vF6XIlVWiAEy/gyf/prObWoxhky9XaYHK7qZn2YEAZ/y2Z4
PW5uJTWnm718Oqw+3oRJEwDCjwb2JIO9BidOI03lF43CNRLyeSwp5npvt+2g
bOkDulSYztm2Au6JV5v+nIGSEBM/Czqh3FgGW/vwTjrBQR8TtSswiF/p7eIU
Gockwo4sDS0OmTnfpp7uQ3B3b+LgA7KzA0ffAMCkq297gm2d8WpWPipJi/Gf
9wTyr9554yuD38I7si90Br4LzWD/cXRK1r016QVOeId6avx04Za3Udignepa
fi62OgoVtMyNXzovYQauZ/dYLV+uytwYpweuOSUzmCElznXw4Xhf79GzQbqt
BEY586nbAxwL8azAN64thWN2IU9qt5GSeS3GUhZYqfYyxEe/8bvIzS7Dgw8d
RORR+MTZIUHEQ2ZH9xloYZYtPdUXsvG7ptsfPz18kyyu2UEh7XDkgTfJzftH
VevUo9djx8T/gH06+FXhPa4O7o6QLZlKAmNAFHH8jKqyGmRGZKYltQwgkHwS
8vBl4HEQcoma4cVuFLlE+OPBTEDKxh6FSQX5vWUnBdG/9F+SuEGxGfMFQJaZ
g6AOFlmX+KJVetwtu/cCjjKmjtEnLk/qzsllFeImOfq/Np3pvpaouK9MeR3O
1IoAQDjZNGwydvWvP0TrFBm4iYdvhUXIIzg185JdBXL3git6eq28mDGOwfcG
jlU6QhD+0Lx9e3+8IVIfDKllFK5hz9smcKYLw+Eo0Ht4MZsF4Ol66zYUvfT7
mMCbCCJOZr/DTW/J2riosZH6bs8xMILksZIJ0WoiyRISuNfI9IqHC30RU2Yv
arIbhwU51lyRRD2F+pMrbPwZsxsBPOWN93LjsjkuNtXr3yJzSrn6OBXJWMeg
P3dIUbGhlrhhrdjOwkz4lp9doJKQirCuBlmDgixPcJAFRn7zaWolrPsbpVuJ
CZAzaHNX7IF1aoFaHV1bWhP3a7D+aW9GU8XSU0xM9g5KboTh870/aHyl0piZ
mUeoCuiIbbFbDX8y/rX/s90Rles9eipPlOPlzAbuLmD5aayNhDi+JAL34fEQ
GUeLjZgjdlNAY5lt6uKWGeWGnCgJPxViV4FtKdD7O8KurYE6sZZJvwMpM8Of
rpz8ispEfRAAgRLMMdSpsqwtBPEh/vlW9WM68fp05qm9wUkTadVVL+oxl1Mt
yvHiyW0uV0911Q+lbkSN7IGy4nTyvsxaX0PiwKacEmcCGSmoZicTJOHDVv9P
vd0yzYgUNwmD4TeGqc0iuZMShOY83EzRCORKCZAglwUezNMXShyEVzshxsmi
gzAaN7rnoDC1J+mPaZd1j+kyoP1bslnmNnB/7ohe2Zj/K6ao4Q6h3nutLnDl
ezXS9WSBQ2/OVXOOIuk3QwwZywTQ+98iZlJfBoNfrfck9KrKosTBekLskbmb
38MzNJuTQNUTznhl0e1vu5s3qnvSj3zMOgfvEsvswhtNWrUaNOiZeDb5098k
qWLEXGnrpt27OauY2qEytrdkUmXC1Rd6nSzvzH+y7I41AQl6BAFM3DzHWWHG
9PBJWyvw/RdBBUqfD2qm0bh6HuNggzNPUCygEyY4IgH9oGg+kCNmpeftbSmY
oRYk/Ib1dWkDp8rSoNHWpPkybWqD2QfE0I/Mc6Bv2vA02Hf90Bwc3RbC7j4r
b6BFD0X2B8BybZ/lMP8zvGLfB9EOX+IFJjviGxDRpBpWP89UgpSU4SNSXXtk
aIrh7fgIpHm8/O4kxlJADGOZvVAX1PDjnRN7e8s7jAoBf6CIWlHYsBRkaAZl
OaXbLGp7wxkNllX85S7bk/8qZUEzW2GNNh1jObIHB1iZUGH1DS54xFa/GP/k
01B6uFWJH9rRi3IW0qfeE2AogLas7NlgUzFhfskJoqVYxsJcjIch+EDjiwSK
O8/OicJdAV4v2tS9x7Pssmq+mv9NtDS9XC8hbKLTODTe+W8b9PmNvsFvTrqg
UKfM72fx8jIMrO6TU8Yzk8ycWb6/Yd4lb1hqOC4ISz2s0Siih+Gu/Uv/aiVp
OizXxbz6KzIx5bLi6f7J2xuKg+7doITc4eqAHKIpElPcbBJNv5BkQPv0hw+g
oPoQhcB9XseCtAzGqDn01j8ks/VEJgI5IC28qNazwAuc3IzewjLzkMoZEkHI
r2tofrJ7HyKHh5n8ShZsVMBD4yZ13a4PpwdfIZWycUeUfIHM9bhsebDjQCEN
FyovEMfEZmTNYAWGgTx7Xxf4RKsEx6UWtL9vEZc8qUc2W/VvQaqm68NSrDIM
aHPsE6fWty2LRbledtSEGUcaspvsaqNUoWjq+h9SaPo6Bk+AvUNS+hP/NY18
11pHNunZaOYkOXPD+usIxdM5mfJPyALA4dRu6HFRoKHdL+yHYLPTYr+q7u4I
392AmR+F72zosW0/7l3Pnyf32PdqprFwEIHjVy/tZp+oIKZMulEPnCpJSyyH
j8ScQugvXZtk7A2SuFTE5IpJ2SI8eGkkSEPZcy+tJVJRuBb2fZRXJBjBOr8S
8z7WK23aUexoyS7RPMGmDH+PYrEC/HcQAo3Zf/00oQvS3x99zjM93D0YI77B
Xa8XUjWQBAD+0FvIbVuHe6Xo/EN8KgirfuwYuVoD0LMcn4C47sstcYwsnTzp
PoU0VLx5qcy6c8H52geKgQ9d1A+qnjqmABWUztm3KhQMo6dTj1IckNPdcgre
AstXFJvs9ovGB+x4EsEXEBsEfN8szpvtxVlfqkhBfEKczlsbufhwhxdIFxtJ
jYWLs5wM/HzDdruleNa+SWklX2oVNKjCADJs8v+lDUm05xg4gVNmZrugpRKq
IuhN9epPT5+Z9+vVhAqJ5BnTDs9ToxfrIvFQ/JmF3UmDc2wlETTa3L3BmT2P
tob4P2r6Vwy4eAZQssZW6/ItPaA6HJg0+oYtGyko3vNaEIxaYT2h04AoziYt
4RCfP6uupx/IWSGjkCaIEoK0uMJ9Cqf6IVwH8U013T8xyYrsPzxKKpmcSW1X
csRDgVMtzb/cQa2788hHB4XkfgiUFCYupPI1xmmTWiRPlyP8rcJddgnD8EpS
t1/bt6t5Oyl6a3vk+MD2jNI4gGYKUmMnzNHFQiyCHC6iOScsoSdcGuinvd/U
jl/Ge5DmRks3ey8mNKDrwRk83zmi84FoFaxMFkQy1jD14/5JxSPhjAh73SwT
54ARfFv8aptmiGspdAQ6jHdhyLlMkhKLUL8dx1iRxeEyD0wdpLr4K1nQbJTm
r5l+V6iuzv7Q8EFc2QNwXfPkfFSx2y4iCPPjP9/S8/aZdvXoc+ZRNz9kcxfP
k9tl5SfdrDAUF9V3btppYzbHCGlVnfFkf6VBb9a2rArIU1FaPDRjoaKrpVlz
NsjGFF/U12ftY/2uWTItxw80PMcCtRKGSLb17462boCgxaVjcEyaUNQb7kRR
kBk+ql2DWzmmhXG8w3xsWY7njlc1ui44PQTUasy0aIDE7pOKy6LBPZk8Ehtc
E5b+RbEwTFzbLcvHKKAWp/IJ97IuM8R4ncT7rXfnGul7ICrU+Y5HQQkUURS7
vc8KQyLjH/WR6AaqSdosNyjhGHlwaBcyZm5UThxJ3yZUSithIPG8auhQNL0r
KJ2gEN8FWtZP5vqvNAm557JYSfwlPlz/6bqDRk5cTU5gctptpj92ONU9IHI5
mSbErdz+8+HL2/T9THHLrpcEI6AvNI4K/pXZ5yOanqUQj8qn304mVIbS8/EY
OSZU5GSfLxNpIcc9Mmd/FoIbPDU5Ekmph5tidAbgf5nN27L0jmLZ3AkXBA9j
PR+aF6VblLwEyH5vQgaM5oiBNPUahUO7qKlRvYAbIJnusGz7im8TNhUcdKvg
WzlU5V4bKq3bMyxY5em+8JIVLEZhoU1Y+RgP5JeEXNQWazy7CBktAGFYkZnz
nNWtYhNT1jiwLsmrNN2FZVgaobPxWF61dXeMoGv28tKCVfcbaxb/0uyqZwcv
G0ILx8TCd0uNTLCFeXlInph42db5IZpIxe24vY/OT51V59YCPBjG8WnLaT9e
iLsz+Z/EB/x2OhSBq2MHnMSTwqN9xe/25nScTJO7Dwcol1wnZS0VpiKPoixu
h2gwelSx2h7Ls2mhDWCqTeNt/m4IStMmTz5lFC1KLaBqZFGN2GdX9El1BBzO
ibnB2HX56SasT1bVpVdGGqN+i+0DNQvrBq7PNmrlQFG4i/daC4hi4F+PFUXG
/WEUSvGw2ZrSeVT9klhZxXx6w7Hh9EfB5rn6KQSR9hQpkL+bLaNYrvww6Nof
5c/6S0z8rgHHHZjKt5Ro9T4GXOgvrEfgTcfK4/P2EzeAHuLsKE/yOwXtZlLO
d87sP+oxOTrTFxdb7YNQIiWn5PwKJGbbqoaLoSBeQ6ztXJBZ0/ACH27XdJsK
kvItZp8Vv7ELCODy0zbzYd8Fqqv2uq/SXgEtSFVdgm9qR9Hz5zNvVibGxrv+
Wx0Nj8f8E+iRWKivPSA5PqT3TLJbSLkRwHsKur0VPPBku7DC0vOzccHwgiDl
K6AWfl3pi1XWqJNkudwwylpCb4Woj0Jqoc1cs7+2qFvJUFoMpau+YSvuXO+2
86zYwJxGzqOK1285CibKaor6niOM8ezAMvgVlcxe4fDMdtUYPOyQBUJh87cI
KWVUXUjMNQA34dnAY8xudQFuwo11d6WAURp4PJROkrZo15p7dm6ZloBxm9Ju
dFI4qxo9N3BoHns4sAhge+wK5IWu9XaiA4dggH1wa7U7C6scmREVsQUwK17O
/o7RHFYfc9dw5R7Eia/fcS6+V2I9vfCVGVJft8dkdbrO2ErymUmMoltva3QM
di4QhTdJsg8+gULU5j8K3ghK3dthuCJgF0O9o0P4Kgr/4jfp8dU/fT4jgVnD
GJlqiIc1KhNCA0ULmjriLcvcViNbUzejD9GAgLp0yC9TkoYUiraWpWZdzIZA
J+8sNzFUjgLbmblx02zGR0AeLlGg5r7yiRaW3elMMXvOjwX/Kn/glAHW2gXs
lUb0WQv6pTkyVO9Gf4r/jE8KEg5grHGzZ5EhCChscY+47/Bre1lxVfL1IQ77
h2iuCaeVwXwH99wJ2V6rdJKytuVXgTkfS8paNyR9Dsi5Bjg8ZRDCudslPxiy
YHTih8A7QxGDw512OteRJLo1G8erNVGCcnd/ITkPM2gvo47q4NLjCKlk4qar
GnK26pHe0LVHwLcJlLS0Z+jO66Lni35ZtCEWx7NdIgSQglTMEtcvRYWwaXaZ
yXz1tOmmG0SoKVbvRjL6O/B6T6ld7oCkMyHvcd/uvzeJFxFNguChSRW673K9
OBY7IkJr81LfOYalAsTxLfGhtXtA6XlmEonjjF/jMZALzQHg//l5VfcgDmL6
kD8O0eeUQk4bcROclulJVYNSakQLaOxIzzSYP2mDrDn6zcrp+0NcpiaByN/n
/5KGiiMvruF/fzlCdhKJWyzl8jsZyOg9ii5ocGNO9aUCqF/eGX9NRecjLuoA
1bdUhyF6fPKs0dyseI2aV2A+Cxjo+18d5/boK55ziYgZe2dho6q55ccUdeOC
lopSuqN5uHPFr+qMj2OyIrZ4ns3n7bPIWAeXWc7MzPgzTTUZ3fjRSgmxLJ6L
iBJm8sNtFacoFKJGKMzVgcQnbWTk3sIKGUQ3tUTAyfXoLKS7tPCGEVSd+DCl
5X62PzsoXU4ad+srcv6bVcwc7+7LqgBDX5zAcomM3U1PYxBGe0OqRaL3fJWy
w+E9rWsLmd9ejiiI7sIK6vtF2ErL91hITVWZMYNxvQ2Y1+IUHO8NSJ+5/NpN
pWSkqswDSMNOYOA6thcnIi+OjSScui6Q5e/QzGmejoPo80Grmw+CXiicxYXV
X4bFsUwHuUQ7FOpraKCBIlgbGHf1716aOzIvzlcGnJCZWfN77AUf75WKkiLC
Jr4MwgVOn/rnesAjDtVtvdJtT2HHThFA3Je45CUIPA/9Um30QQb2H+ndFCZC
iI+JmG+VT3xRoreCuef9jsRg24qEp6y1cyV9lg5J1ej9VMbdjicHcF7OOr1H
yQ0+u9iUl0O2zIyff4ThNIymWj1BTnfUvlfLb42GlSd3TMM5hZKlS/G30LFa
EX8SSGFH6JWeTlTPwJCYDcrCtn3p6ae0OOzIqMTPBtH75LHknTfyQE13d7cv
d59uQyXmqC64GcHbICuvEOuUVs0/TodV9AWNXgiGJQO24jvp59NLxQdtXJoi
QEBu1Zt48gOPy6vBuxxFFpH2nE3WNsimbaMSuBJK5uMBybHRAvvkxwgwnM4k
RgOkknUyhSUgj2DW6y3JF/6pDdXoD0c9WN0xEKU4EnNJcM24Ta9jjHChS2Vk
Tjtf8iqt6CNFgrfUVuggu6Muq8tM/U6YuoSd2fp0WE/XVLVDRI1rlMeOK3IS
MtpnubsDGW2TO8Avn6/Y5QDD0JnqjieV5xKVdHmkrXNoxwm3ToZRKoi5vUf8
lDw0aCsfL+pZHkHGJfTs8SCJzpmfEEnhhoS9LvtF/9LOS5jatwR8fqxebIyM
qqLg4HZKpGNqRKjCrM1EPkq2ckOFef93notmqIkrq4e2Cpndh84ticPMcMQV
a1LGAz7qf/p50IlvUYo97E4FXjFRGSaSTKAfPDNr+k9WcCz6a94brVf56ydM
XP6ORu6Rl6DYC1+tME6z3vrSIkiGHlq+XvLsNr2NLvTc7MLG5tkXgz4IV6e1
LrWrbrXy1ArLM5I0NUApiJrJlD7Pq91vXCYgzqBDfEdlzkbKsPbsgJEA4J/5
x30HBqLkVRj5PTxcej4/yR6atuM/38GeFYrq2Xuyh845ltq0EqSpezT5iPzI
pKlRhi66foYlzbzw+2fLxtwkrDukpssGwuarcIdwWwtk53nkXdlWQTJWrPC5
YNkNvfbT2PRVlSzQNlffzwanp4bXLTJ1uKGFlZvAjTWZGRRJ/f0EFdC1W5p+
VjGkNlVEnI+V29GnEmkWAurgCxY/I1uRLNXUW3Cr9wAS8vrjE5oM8MS02uo8
z/JKJxzDj55duGWPgkPDbiaZTDLmKLzjFw2FeAgFrGFClNzH6ItM40pGCp5e
37V38kUbtAfMiDCk3LTvUXaMJZ+mWm9dyx5sgSu+qSrf2aWtVzzDBuT8zfys
gQVz+ygTvrL+r5ThrckmVCwBrqv6G8ZRgtA7V0smn1I5MD5c58aD86a0/9nD
0nEA7FBe5Kuq5I7PCbUpv3RmYq4YK/gW3XT1sr2rG2X8L/nXhXvTHybALPdK
H2DH1qhtfgqEsP4GP17Gr9SqsWEDWnT7UlBA240N7nqQF99fnBrwSWgWXFoJ
T/OkwbWDfwkw9O7bVTD+O/fx31GDcy/FKECQrsumpdx8FisRWduFG4KH7Cbi
G9jLj/36tQhd/VWITGYiMZmQsWJWG4NHstRMhAg6AxtGsRNtwDMsi/cUkrk8
BPkdOMtpdopdwDAg13Q3W8nXLf/oDBOoC6uH7DdPP0SAfsO77fR7DAQrMHhS
EVedxxYyRuCzAVIUl4XoG7Sm3h0TNfn7IclIkT37eP5lOknixKGOl9KvUEjg
rBGAiL1jc0g9MdjtLN0+Q1vCMiPwBOTSxGso6S0ymBIVg3Ol9VO8Us79cYiy
ZErHoEN9J0Q5mldiH2fOu/fPXhCwYHNThKCpwlWS07solSJFh+QD06qVqsYb
KnQEln0yHMhbHyzVm+QaQOlJqDFZsDSpxTEgWxmchiAvRx1Fj/26mL4AIAxz
9kM2VFVNGF+1utFfZqsBhMIueg/8BQzAR6W3mxg/Oz0611zbz2UyLpXV/FBb
3N6WhJ0FtSwwKpLH89IzIBW8PJ465MRCdqGSFP43/PaOXiYV8orrFXByprvj
eGorX+J4VnqsCBBjXrFAmtcJNyhe9bHxoQaT3dGGk1XNCscGrX7Uhb+GPfIe
VzkCoFiQ4Rr7ehFdtZ3hNSGkYBcjcIoWBa9SBzQOFBr9emHO38MORNr/jONA
RyS3I1CWTHrkcPrro/o+FyYhr2pAkNn8FiBnpRC1G5aEzBQPOcWKB9uzAXHl
DV2MfrfyDad1HC3PKzxOjv0dphuCLqQqpnAnHLvjc/I3i8qRGa0SKcG1Yxsu
nvL5/H3IFaOTI5OUlyL3svtxR5v1/ByNwfwHr0nRgTVYka+LopOHHwOG009N
b05Qwo6zoOIkNxugXglMgMj4/yyqrkJ1IM+oltkaMk4F5AIpOJbDmVePE6wX
u2nJYgPPZ6f48yZMICu/lblsfOPfcRng+IhTLlVwe0BXosE8nDD1ew9QZDcF
uPjhvB54GgoIrYTovnc8DVY6EhmvhEfa+wztAM+IhotMvWP7DnrkufcWqpra
AoqwTu6DgX0shlHQjJVvWZs/Q5rJuSNcCxkqAqgHETPorB3arA7/qd5AezEt
IURh9StFsPauPKFjr/Ow4YcSsdy9ee2VgW9CPZ7WJKt+Ty9mhPItaO4ycHz8
BrE/F51B4sUm7eVOXR0TFcuEYmnPP8jKtEnLfgAOBF0jf+9wS0pmZ+BXMjn+
IE8k/UVozxXVx/YCh5bQ5BYIpVrqnTfRrKAIIpWYOAyVy1Ie+52JGcWLAcLn
cAOJyLxRcseVu6jO7OfvRJvC+FwyWysduQRkCyCNe653N0xU7fxVzknO7/Ad
YH1UvLES3HXXLs2jrXXCqjqVC0iIfQ/zfyTIM25OobnuX0XqtHdDPdPlcCzb
mjXf5G/J+4U5yUIIO9NFDGkPW7x90W4qb0Nb1hJNX0duVdmGiU0zs0DEqJyw
xMk1HP0+B3UQRM3wVlBBgOpU/y4UkeaxOHfsBc4yts1qsP7gLJILpgk1da9B
r5KK8xaUDmiJuF0XKo72rmAn2572Fu3FyqBC/UV1DVwaHsFTYSaRZvgJ9djV
NNqK/nrlaqlxoU6BEj7v323EmDtHAZwfJqQxr5q3QBQgKB42nKLXx7XY8fzV
FR4ej8UgF337SrIkJtXvNc7NhKstSKBTe8WFEOEVr1EJHTaS73Tf0xKZ9OP8
HafnVvt16hYrnUsX1Sf/Uqkm0nPEL19AGXXc4BCZvYEcw9oMt1nFk/cBbw1h
c1+O8zWh1XDkSBF3/mjr4yacRNxFAae8ga1e3HSE8r8emZqTDXOquMivRHaP
5+Ij8QaY5+G8H+6eL53MQ9KEXM+VNS++HHE1dYaN/FwybMxZlAuQ3pmJy+8r
ibeXwo8be8oZbKtqFJpPnlmRIpsXZRB1J8i29fBiREkE0x+KvKjWaR1xul98
j7vKvIGvQq/Le+D197HKCbp42VWOfigglx0hU0HAgIABR6+fDSzI1FKIxtUU
EZm+/locIRk6cOPY5saLtirJSBFAGx3mZsKuS5wLJXY9+jj9x0LvW4RVEt6t
jDAnmyNDU9qbep+AxPF04+V161U2kwv6W3QXh0OVirVV4grFH8ERLJZGva/x
oJSLQfHgXQHvroOLYwNE+UHRnU3IY7QonY0L5YVYfqkkdsrt9cx33yQOgPug
+9L9IC3hhAcsIZ4bJ+JIevyTCJLXyHU/vrfwzQZ4PEiKqCYOlwViF6T5SsFc
ls+jWDZcl/tSCRI+NgdQiw3HvmTitNR/g8xANpXm/CMGgO3zJy5zpe3/DPoG
wtvigP0i3/v2kCP0KH5bliEH0hoSpUF4JuZu2pOkw9SPDo1/Pp0QDhj7WB2Q
/4yplIgbtpP+qayZQuQ1cfbuzGyN4KITqzxIkEME/rmWszLwewSnDraZ7f30
y/vXysn6rNN5ZDZkM3cNmslt9J1b6GLXBSFflWkzSDEJK9WYMmKi2gRuYxV4
voIU3SC/Vs0WLuGxsuy+85EQcOpKkhT4TK0Bz0UT8nfgP+/WGbcEBapmCO+f
X+3zDImHe3NfsYJc2hL6rNQvHfHOUL/Y8fmhs/NpqaHLD8UZ0BQs/HfLsOp/
4hSnUdzrGx2VyEXML7HSclsJAx5toIpErGGPeDJ7P4bxTWgEoG9EKgvwdlK6
NufcnzCNKFN4TIlmQsHcRbJnuxfomT8/6oHg5VK6NzLNx4O7l33YpMePA55z
f9QTVhPlKudKuoALZOTC1EaAdxt82Cai7sCAKURO+QuklVK9ct4Up9RsSQOG
o2IaY8cAJVLEJVoF0wn3zGc4VP0AbJphZXYhH/9R3p9j5ek+pCaOT3sKEeSx
8yhmnuVOu3j4FBhjI3mjr42d8dk7Riq2KE5FDtSBKE7mq8kXQV+5VT7Ep2gh
QEdTt3d6FSWFblq7eCvdljXEjanJkRgiYmpKzZs+frAyMGS6XA5dW+ASNaw2
a7OWh8GayOBHWZ/yF0i6zIx2cXQTgYbstkviTTyJM/zfc/6dz6Afrxxelo3X
FnZI/LQ5xX4Wjyu887Oi1tsOGcU8i+p6lZ9nST5tcWwfp49aM8MyOgZfLEx9
8yt+g6A0mMhfV6/HK8fCbYn5imYpKtMe4U9KEOoMM5/ClGMYhXzkKmVM3/0A
s/rEY1RARTPaAcyjoJ3NbG0NOCKhI4VMU0RQPxlgmnPaQ15TvgOND7VIbAeW
I3CMSO9ubnajSUKXAAxOToC66rGthsCHEAFTT0WkOFPWtE1BOAlxfJeR8LSS
t8SFK6CLsQgxjLnicsxDEcz29jBgWl1GjMfAA7LLB75niCVil43lf3Y85O+G
+DbKJQ9VHQO5JnI3mjXznctLkggkxXmhDRx6qNAe38Mb9wQZaamfvmg/bG4+
6JvL6D0g2yqE2dOj79QTlarH4qEuu/RASa6I/wjaz9uDjO0vuh700mMTzGXj
gk06xVaFVxtWT6ZDfMOZ+EMrZoZ9KsROt6hqfJ6IjFiEqJu+pSyUU632v1NZ
iCTpN4V5Ghsn7517sNEEy0lfgUHeIn529ghaapNotSHo5BdxQh6zNMgOJMCE
3CL1oazWrbvnmO8m7ibs4jTfqv410OwCe5FwVzzuRWqvejB++3Bl1vsIIgny
/VB2/1vqGVGzVTt0hhLp870iBpHN0mmNUswRLsQrea4pTXCQ8vpKcqVAGL0e
TdFVGkGmmm+Ye7eypRhwh+7Jo/f5Cw4hrC4O3MQr+rk9XJ7rYzHZURkqQ0yv
4LbMBDhxngbCYYMVpXEthWFMJs9B8NRaRnVAzDVB9JQt5kwx/pjYxJCAa/lV
ItsYWx6w7SvOLQ5OKl+QTy4VhyTvs4LlXOw0NjEJ/HSHn9KAkU+k/jpF9dY/
wiQY0jcJaEJ5P1JudnCuu3d+6QfEDvf3vumNZ/PqDfoDg595gIfIFjb0lKVf
rg5elR0bT0x3oKXurXt0s0GRX01F7i3ovB5bIzR/zvA3OOvl6/MYCbnJpcgn
N8w2kMa9Z68ZlFWb1pxbosiX4FCZu2aZ5EoTFTWem+k5uKx4h3izZf80SBFT
09mr7PnNHMMVzp3VFwLIu4caWFDe4hfseLZtNXHZ8KIcIMXHZLqLVvMfM5Sk
Q1D/wKexW/PUbGClffOxZoCBB9mvFgTzxpugBVmYbzY1jYosR8z7/nK3mq3z
DGb++SDme/J/l5k8Qjjj4zqozgPaLUtOjjiBa8ri2eXRwPgc957y6rXNO80G
6kDsAhCjV1Cpltj139TSovXCFks14G/XPkt/HLXeoHI4n2ZRI9q7fcWKMo/W
oxO+K7hFKj6jYHhlteZSMKYvHvo5eWeJ2I97mNEw3InD/qfUrVyefiHbFhz6
A3Gsv74RDl02qWt1Yzu1huM2kSxar+HVmWNICpfqHR/eZ/p3duYZeAtsbyaV
3ULJobamWB/ek6LucP79ILoI5h9XZvUT9hIOWOWDrAqigUTNCjH+sPUq/kne
nQErAp1iq6q3whOBx0fcu+rzpONZDCNKCrG5NH2prlvMQYfE9ewf+hpXrG3h
coQ0VwRHEbIiCnqshfWTpOgfKjIjPz9b45IS56gsXcmjt5WkpGS8wa+b3XtR
3kTGjG1RQB0GJ65SHl0pUGo881LEgCVBwD6CqcedmN1H7tjNFqiqX6A18try
nkcsCud3oH8fjVnMztzyHedhGUiRDgLQYJaM9aaV7IcutsRAyOXsYPfG2FZB
t6rCSEGyFlO41ykirri0DxGKXZPcFzNkWaNjQB4Wcj+/s3QUbxyxfJLNs3zY
4SxhzaVh/Fns4fa6fYIO0l52z74blx+LvXIMds4G2PzPwbk9q8JnpTolNwkT
HUcrONuyhsaaECoBSPQHhq6BMKL0r+XxzvNH3EU8bn5Mw2E22LtVCjquOYXO
6bOLjyoLRlwA0408OoDO5/OMrPPueoqwU6nd5bgL1NZqQ4iSVtJHjkIbXkZ2
HR7GDIh8ESFmtXR2ca79aniOomByEPFbt96ARwdZbt9FuV6JKQNVtuRGfyg/
hUbbRBdCM9g7AZYIZnmp5t6ylSt/DwlI/RCQS6370HuIVafGBIPy2LPhzCAd
CBM6it5b9xVNdeJv+8C+/KhGVVXv/eW9S7lcbuhzxEEhVS6t9TlgAZjlZnUg
9PdylIbkG/iTs1tBCY0h7f7V+/jzk7ZgUSjQnT/QcapxbwMYwB6UbGr9HDvQ
UlCYfFrkfxCfc0XF3qoKBzqF9CfAc2Y010HiWrXO6GNxx8bdC9ZwVybe8jjV
w8aDRFINNdAn0p3yg82Dv2YXswCQCFKEejcI1EMAZCxXetFkc+U6Lz3f9Zdc
rKUOWoAh05UUf3i5QbEHpUVoL52mhojtuAlVAfmm7R20d/iXnxy3D4cJJzN1
06W5oSGpmh6yiyo/M/enyvVjg5nnR89X4gsu72AmtZd+wsqD3Zf1r6rZ8eqi
mC19k/p+/7sQm20plh1LbriVfXd8+Kh/gsUXNdIvowAVJALR17sqJUcoqNgH
R6lzDWHyRw1abPmCropIW/m0DZRCn0YLyouUuIKFF4cyI/EeHQA3SsjwcRxa
LLHKgxPYGbIZ9/xjjb8DUdIOQ46Dp43bpmElaP15L3b6XC1r3mOn7ZvnIN8S
a2kkC+KAjcKPFMsMQWb9j0nM43flncOeGNPx7oFm+9bobhwP1J4p1/5+QNNp
yTmjCJLvDkoTdMMTMw3ZwAA9rncSgxrAsRGB/6nM9ygzZkBek7T14jSga2Ig
MVpGbPt1DfADM+Xj/QNf8Iuy068pPQSllp/dZL0TD4jyw/AgHY2MJCZqbB0a
sWxSM2ZYRiLSaubqUB07sV/bS6FBbVGJ++g8muaQBto9mlNLTqE7K/WiVAaS
XZnLgTzlM0Au27MOZZtLOnCpLfTgpWPw8uCKlq8j0OvkwJnCbGbFBF3uFhS2
06OgNpNccbOFVvDLBp5wpsI9QSMinEK37PGTe86OkyXr2SjjkR7HzrCLrdLR
CqrmiMZTRLZTDk7IJSwY6TqVMTgDgrgYXep2VIq3nfDUME7wkVXre6ratjXj
/1ROyKqxrK/t1hR5B9ed0ax2aOO79BB6Xo+t28IJ7SVNDv/69d+FcQ+wEQAy
KmxMRggW+YWCDqMLJcLNLvU7KvFGHsdUD8XYdij15O9oNWRA+tSBm2tElHBO
6Kx3ubUNkTIJymD7i80dCkygRR39zLutya16rjXJX8YuRbqVrzKE9q9bVn4w
50LGKARi8eRCtQNH1VsoZ/wOD2ZkHuOmz9kFPTyUC1Xfr3tXHMXbwRmQa0t0
mbxPQqdSHPq7nqpLEsUH3ae+74N0+A2So/IEsMqtC7hkUrTnWREIoBnMvXeU
U33z5piNQBi1BMSWVQjo6bwzAcjVxd/5YfiH5Fh/rSlQ1wOb/eWnX/UOyQu4
ALUJN9ZpMFzp01b89QOELw3/towNaq7/91Oo8OnRZulKE7ggaKZXnNvM+5J0
wEMqqkPgPBe0ryBK73nJJEapcgoYkFcRQ34LXmJuPFlpDs4KK4MrX29WKS8z
MCetjg4tEP94kZihHia6SOvzVMJ0RqZHvIu0iqHkP9CUp10i0nVigLFPM+l5
Y3G/tBX5n+fbWBUKJgVOhJfayCAR8Hn/lnUMJyZxZxFrXxTg/nimpaPo27Bu
dLOqiNJHHTxavyB0W0ZrMMKRE2nRlmZ781vWe1Hl40HoN1x/jlGZRRzc5Oa/
O5VZ+9pJMG3t3YQ4Yb5l8uUgpMf/p8H728nvg6QKyGPSfH38c2qlbqMzGKSx
gWKaDrV+XR15MXhWfk63AxcC6TB/VmLZsVmkawNp6STx7L1p3A0fsT5mGXw8
FXuFMjSAuIsYUijjQ/E4WXu0N33YB+yElC8gbvAEmPex/f9+/8WYK//WHQG7
mXt/xIDHQL/HvpMJuK6bw+1X/oSjKwgEYjBFgryqWArecdnNNz7OUWjTD1Zf
FLs4GF/lPl6NgroBHkw9o9Ffy7/IDtU2qqg87jKDVqbc6siEOAU7QclUroNI
mh+RdWvdGSChOVYrvP3HYzPSbG+2Ftu19mkb1SiijHIilsF0sXoOy8yR1H2W
jbsEGO1ALh9AW/PlaYLooYT3sr8LrcJvRLyDCD3PcpWxme6kSjLrmM8o4Vse
mFQZzJbDWKrwnuVLHFkGfvLW9IaBOUbyD3pVQ8jSDcOB/dRBjPJm/HJrN3oF
nmY0ddG130tGbYJrs8IfhjEUG8VK0XkldumuRcoYwNKNHZ7y11zRP3qE/LjL
gDPfbcFIrkU60CfJijNxlm6juZFvidVBtz/oIYRW7NSN0fqgFF/5nN2CP9r1
o/0creoeeS3y0ZOdsE+4fsVZ0KoWLl/q8OFnEjd4qviJDb8eZw87S0BT2MiE
AFUposchxMjeUf8R8QHtm61hO2fiUHA4YACH/FXScHpiMc0/ih5HHk96CQkp
tik/u2hOGX/H0dlOPWocNC7atO0yc93f/dd7Y/pmqgQAjaTg/QEDeSIND/WE
pG856bs6rwIAI3RkD4zMgWZfSnthfALg3eRD29o4G/3aXtaPct70w23spkXs
2f/MeXDI9drtbFHsauRXjshEHvwYf0RD2a1mP8ylulm9J7OXj4cTUA46xBIO
Zyf2CPfnWpk6bimnOQQfJIFsyFq2rkLZyf380D7AlMUw800mHk88M7DKfYmd
Hodz8oXXnM4AofT9uY1JliHIOOFzboVxSa+H/TOZGlXObCIqBm/KiXv9ahRt
Bc9TM7fQUWiUwexO6j7d//Ot2pD7//EwOQdvZQuWzJOM3mV5IwOLczvi95JU
PUEUYer0rETqHXA4/uWBxwiB07F5Y5TRTO6Cht2O0Th8qrcnjeoRC8/L2ndA
q6K+E3siR0Fie4PS0C3a3QXuCIBstokabhdj9VBnUAom8uXhwzmzFWqZbUbO
/A6Ni/WP8HLVIqzX9Jm5KmFfyqiTWlQGF0EfJo9wKKc5t+9oXb5fyceCe4TK
nUiAQx4e2ETfYFvxqoI7IHXT/M7Dc+S+reXAhlC3536tW0b/lNzpoy9kpxd3
qv+axqTe5FmBgVNsLhbb0TcvrQmmMnieMwZcTIUuiqSwVNLreqXhvy2I1xrO
ML89pA1kTmRywjUxizkeodX+mrFngIEF+szfmRrySV1xsiH+FG6mSPpH5saN
a7T7FVYIXBkY7Fc+Ekqyr+FJrIgQU4Er+XChsiupV/vqqAEApLFn5kZ2nAOM
eLqX/SrSdRS4ykc+TeQODTw/fS/uX+Twf94+NRfX2/d6jR+2KohYWqGW2/Qr
pyXznb3MlGGq9VbIRLSSrM2ysT9BvpYtso4X2/r166kDpQlL41Vs2ko0bgFU
Y17uC0m9v+bVbWkBoLO5Ng3xKDb2JbaSYYIyYW9KGgEP68pFABQs6428kFT5
45waG+3bTxhwURNf9qqI41KwXdJWaSqzu8loaTKfXluGsI5hX02dfnHCHrqu
OjSkS8d2QM+BUchRMo+ZWCJHaPNeFkcQ/5HLlqqwLFk3IauOEfdXvy/iW8OT
z8EnATOsO3P6ju/reviaNPJxfRRW8GLmq4Awyl9wEs9ywI7KlLylbnJsa/p7
WeGdCPrjwsuh26+2QIkL/UR300lVjQQFpwrSO9rBu0cSLPs3gs8Z+Cj7alSb
1kO5zl0LrjE8kgKyXxOakhv2j3y01Oiwyah41EdSnF7/NtMJSNnBezUbJFUE
NXZM5lQfrwuH0kRcx0mG25A71UPwlvGwU+w2YCTdSnPqHvhwt/x0Cao+8Fw0
qBImWuv/QVghIEpN3YEXIgr1AK6Hh7EnpYlmlLmsR+G2psYRl3Zb1JpaRiFo
lvKAo6EEz2rMxgt5A6/M6yCNSP/YjW17zwiBt06a+xFuBqjx7LiO3ZK9U0zP
D39Mb2jr+LCyVHFsV3y3rCL0V2hvp+4rKDnOqFb4/eqVqa2LQmBbpH1AYkPu
mmi6/JNgdaLzbM7/CeQ8As4okRQV+mu/V3co4c3xhU/2YxELG3L/8aEY5GzM
QBuLhyNNGM5/aGOxakowuZzTdFwYwCEt/wL5EqUVvwQO22r2OegVtQq1TFCd
2i++gB/+MyZYltCmxN+bjKnSfonubGx+SGlKWt0hLF5Lk7kgwMZlab/xFcDt
yRoOa0XBaXWMdC8PC/iGoYckb8x7hHIzND5h0O+M6mGJXEMVt9EbTRFXT9Yp
rSSe08iSxAC/GkOmxw2s88jnjKgOaPeUhlCcLe7sD9j2GieV8F7t6KHLrxSl
O/xjRyFoIyyIlKgfWk8cMoE9QY5i5VgQEJByMRHHStYNTsvElzCP/BiBMHQp
lDUFy2GF+hvLq/6azNbKcb7qWyBUmfBGZG0V+ti/8xayB1MmTtuTyuJwa0Te
pgF4OYzIzRb4ybDV3HzYEn8PfCDjROCrx/ESF7nlDu9b2sO/JkjYFxSEKetk
rUc/YuLz40FjAoq0w7xa7aWD2GrzA2MYLh3hMgNBrmhAV0/Qqzwrhczjtxiq
Nj4efKCYQj16VKtxdf76O3QMatNBuUObcXI9YVm7W2Tr50wi8DvHZpyQzT7Y
k8SwVdSvCA8ZgpB3nbtrS24bFkv65rrtLmpi3zIKAah2RQKP/rUNrC8adoth
QIYI/KHpLHNzy1ChE87YLQwVr2g/3cn6XzGhpxyWJd63W4ggRBYSpqpWkxfS
KwaxIFc0GyOrooAyQ4pD0XfEIzy9DV0lB3n4+CvzoViCHNWUygf2uMx/1mqF
DR/C+SqlHuUp+Yx2WGjEVezmvVQPz5X++6pfuATPzJQAGdcjv3whhU7vVOwz
Y8oD8hxTUBoZvJuq+E7aQmJWXQIu/CsqRbmWya99yAzRx2ilTu/NFmldhP8o
Lu1u9tELIIgvavObeFZl/VGmvQ6uYtPLNnGDWDU96dBiaPT4aFApNBlwMnzA
I/KKuAhfe72ps8RsqjLVIDvxHCiO3frp4ITYrokv43FDCRk/DBMwGyaj27c2
ecMNIyH4WAYMUfPB4YwdD529meo8dbEC9i2gjJBBLpvCUnyELZsOrVXeBT2V
au4e4I+bM08Zgw0wsqtBWGSSOI12iZ+IZEAT06uIKZLUgezo/AZ2VTIh8PMe
RMw4SH+VG10pkdgXjPyHPP4RXP8pqgiy5mI46jveFlgR0fzcPwR33srR779/
jXK/v20UHCvBfl+oC7cMvihzVpmfWRAEs9nHrvmetneWzrr9LfQIONtdJIyk
w2HwwpZ+J1L3nuFrprF/wuSQwgdGgXBiWZEo4ckEbIOPqjJ87FdX38LsbTTF
JPtc0zggqFirJJsqO6e+RdmRtjSsGm8SpyHv+SMjt1KxXTFWVQ2ub9itIW2G
seDB/qypluc+10qS115jwkCUU7CvmKPQohmliPPU8LuvD8YXP1ZXfp1spBWw
Z0un6pOlncdAY7Zd8Jm9WfWSMztir9J2mEUtftZrvalcX4uAIVPGff9+clH9
IE6PhoCfwL7ySkIwCLGke/4SYDRUBRi6fDO7M5Ka6n+SnQ3NQnCmH0GWcjHm
FXiwbmGwQH67qIZCuatpDeeTSlFAKZsdXTpMxqN6xzhZB8wpMnmvpSsix5nj
+r9NY1QR3qOQXD+E9Udu3AEH2VFA7ja2v5C/8DQkw88IzlhuvkQF98/zLoEt
ak1qVyDA+SKd+lcgbnZIOj4ur/vM6RJsCJ/xom/h+8zaiy/QEDyfSZVEOQls
1ge9xnuiV+6ykh39Romuk8SYQjyhV1X9rQQL6LBFD/KDEKePcII0Hi6AiTyv
PvHHOU8HpVUOh2CmdzHE9+H2WKd2xTQH81HNlp4HP71ijJP9S/sPArorCHpn
UeWKB5amybKMVQyKvqngfbauOXGWyEIlD4dl+Cv/uJQ5iwbidGE2pDSToJxi
DQvxH5Qj26UGIUneENZTGXgKuDmMjUncSNtuagMJe5Gf+2pjjr6Xa97ASpzA
ygHlugQIYGR1RVSUJOP6chV/jI7WBwA3xNPKGNTvcrz/zEr5thbu12sEEWvI
1DkUGr6OgZkyNJiNWtsc88PvIez9sEM3SQGeGCEJgo0axEHi7qkXcUASic7b
0tAVChlDdIXfZ8QdS3rDjn22kTGFwCpyIYIPu6JTas5PF8EyKjpDW7/ly8qh
eWcwUhQKBM06YmqkDSylZIegGFBxaVSBj/ub4QmvnjTUzZj7bou5v6RPDB7x
n88p+jjh6J8xrKy6DC1pwjlAYCWrrnIY7B+HM7+/BjeRSBwO8sIPmImvRMXc
Ydj/UU5hLR1P9nQ20GpxG10C8qQ9QaEJYHjgtNaYe7H+jqf+i9WsjzKCZwkf
8Jdznzrqsqm8aHKxJZXpCtSFpFqJmZJowxOQm5+EsGRhGKIZxWwkWaGLj42f
QQf9fpI1rvTOK/fAgDhFICkt4hhIcQVfdAD0dJ4lOa8oZ74thAFqd2isbtTQ
03YQ2Bu7mk6BLwTOx4keVAW4OuASm5dmC86fcsIxLoJJNFI4abRfL/YzTJ5h
3Ob+TWL9lF2RHKFa7BWGNdoA/ZuxNiys76KoZfKhAM9WUqZK08FfKHebCbBX
P2hnCgb1VMusY/YpQFPKnTB8N+5LQ47g0xYldY8KwGxSmMdbKWi801TqmCHx
Wicu6u03fH6Bljpav/oqGRxELvMECk77SdFZtg2SZGBjgioy/E79RVPjBKRt
CKRnJBfKxn3lr6i99stTzer5FKq/t+c7ZVnyWsiuC9G/IueEthsuE/BMHBQx
Fz4UDqeEO4Xyf//JmE9Ag+hn8bgR7D+hnINhZBn05Bn9QSQUUAMUhXh8wmOO
/vM7E3Cu4v97uEHJRGaOWWSBijX0vKY/JRyDu9rNs3OhBzDltbfG469ZrRHR
U2qeNM30uVICrdrubDybu7pOufx1ZBgPm9YkS698+XuNyjkTwotsY1/UFlZQ
3Gs6MEeFzdFUfuwcep4oyW9QzHZrcbN3d5ITAJ9+h+e+OL40ln95nYr4TEOM
4Is+gYhmGT49PWYV39KDfgFSXvpk5uD8wmt92fu8rwsgJEHb9heaCe3ztHWP
NmQuNK6dTVw/T+Q4QTP79UERHA66jZJUKY8jSPXEjh4dOC9E4WbPOpKJQv7C
DERmcvTYX0F8VoViubwzTOQm0nLF/xMT2TfHaD8kDN7VgjnuA01yT+MfJM0j
5Y+YO8bldRRGLFv17AhUjn6asqEIbry6Avek0IRJXg1i8YMC9nAvF5aLF2b/
jYY4BWj+PeBlzVZNk4WsSJ3khfamBKt6AdtMSSUov2k+75aw/muzimkKw70d
kkavTM1tmqZQb1GXjVpNC0am2HzTpf4tt01rCZZDgBtQWelMqo8ogp3Zb/OH
bgK2ZgKwX9qG2+3oYet/XqFhgdD5aReyqf/2rN8jTzfQrBO6dpceKOeQ/17V
WLrYOfkjhVIUBYp+SlOps39eDWweoIxB+UJekJiI2gXEDBzXHgR2kn+/snqN
5xkhd+8b4TNcn2mEgET9APusOdoPo2zJznCYRjSD1UulgppS6eKp+Vzgs+dk
i29IiiTfkCOWyySMYTg1Zb4lTooV2bEkKdlehDRj1mGSrqlolBGDHVQYBIpC
vk3BvQeIj60pd5tPBc3HaNN9tpJaIXhrAZhdTWvQFHNvoSRPea5EifKkj9a3
VyPstnpz9kfbzfe4lVeoUpWYMiIPm5JXZxpOlbfvXL/owCVvT4uroGx/oW+q
tsTS6FDxadbvg06M/zosD4HWinyR+yVOfTUTpS410XWDphMQvEhvVm7sLkRV
P3fkrLm6kEPHnZH4pKL5urNL9xS0B2EgipzOH9sekML41ulMKJj+jWjjOjtx
0iFQtHXoSLLqRVhTpZjdMUyxCEOAVlRhgpkEbqxJB5gsiGsPFru2uHNZKJph
IVF0Eho6+5O4JhjKox6QkbJ4g9XC+nWdUg7yDxKfHD6y963Wi4DN1X5mDTyc
sCrmkNCpBSb7sjcSpfJvvNlnVUO8DbC/BLCCDoPL1GLIQzFAIgPWYIEjydV9
5QAam8QkJdUi7RDm/Ly9mOFLx5BNNJEAk7JvuWqwmNg67zgKOU9akS8Iv7Ou
w36f/neBBKTSR6s8EWBCKH0hoBidCAhHyN/Vbaw3GB7HlZeB4DCcBgghRWQD
QMWUuxw2Aks437e0I2icGbtSg06qYceRXaEotIY2KZElU+DEh/VQ1PtVkD2L
CFBkrwTR07aPh6a+dZyfK5zM9qY7FL5bD/FJh/+rR0lDgyOyp2zS6buPwSWp
hfe/Kn2NcUfnrDanoQdKMHRVwWp/laO102DLvm/RAFYR+BMMUpL7m3hnxNTx
XU1gXseblhRRWBM+TBQFVB7oE2rZvzEszJyuvQr+BZfvnb2yXWMWsd5wrz6t
PPM2tEVtDbyWcV3Dr4LkTJkiX31SKYf59YzzzqvQjpyNavDwBRqp/cVT3mSc
c4efFcr5wUZH3GCu1SYTsst6Xq6654Sh/Jcm/AR84vJPAyJbd1QyCZF+AwE2
pb1Jr45tt1+8FSbJp6yZAV815A/GWhDbmt7XRrsKQ1RD2PQdvkocsr4QfvzU
mwRiyiL6X5S/GsWgVfiTi8/eTlWlyeO5WwPuLLWIDfsrP8ehwDrUK3SpV8x6
AWRTmkDG5j6WOuXOmH3eSfGx1wgxUuvmxKfJS85/Jf1ruBEwDyomIVzKlMcT
+QLx7T6ChT5ZIQmlYMDLmvgbPj3Vc0qEn2bHGAxaur0j9t7yOuSXFgMlnlFR
rmGJUbx5nHMTxzGfXuOE1KvxUx1PhwV1SN4skbzWX95mrFAvmEAsHJeAZrpP
Vg3mr8MN5k+nL6jKcMivKpP1WLpIeBXHm2Z+k/TMzRVqs58h5WGOHJeLBXgp
Yxxj+Ej8LqohVu2uJJ+VimeN8fQelhw0OT1OTcMTPhnjwZS/vROgM1xDAiIp
axadCxWsORo3E6tjndwtVlY36eldfI2th8a9dGQH2PtMUeXEjeWZwCpYYbD6
QSWUtZWxht6bBmJbmNNOEK36eCVu0rN1qEd9OoxybyxnsLQzzEP9FeyzujYi
9J47GeBa9g+lSYRZJiMwyCXTfB+SHpvvpjY+jGB3tkOf/zpCxHdzb1FyRqrf
XeCpWQClHny/kitH9C9NO60ccOeGwT9gkG8btdlyrfrBzBbJhGvlEsheQNtJ
ksxFh5ER9feC1SRWdF1U131LXs7M0NBnfpwIVsqhnJ5Wwy/eq5xqgyGi/dD9
/m61jpmKQ70jMNzqwmAjxLY41aFdY2q477O3wXUKPC4OLcqduFroF6awx21e
xPcml76XB88oonvZ7sygi2C4rN0re6Ukq8a+E3QArMLnqJ+6K0tLCYJdrzOz
eeSQrnVRwDokTKWHrHiw/gNiPN/MTX6gbVYu4EO7vngUewSrcKwHA4cUYrYZ
4rzcNxanDMnvfDvGw2gBl9Pu72vCT6sMjTw9/eyNZ7qS1+TJr5AyDbcQlULP
viSJ4KrDX0UAjdMURvJs55Lim0MD082xuaQLXp8UXqPpI+J+bDM1pbaGBShn
4qv48bUqWFQQqObh31pl++wdSEzwhZ3t05Lr774ZZ6Ws76bRUZjfeqT6tbye
3UbmNZ4go5nglFVnSwKX4qw/gFBcu+G5mmwjITRaAt13rrG6VIXmVm6IDnlT
FnypXZZ5JYZ2AHUUEIvMPic5s7dozw42EDrcUMNbOKPBmspgFRNi8VvoNIRQ
nS2DkXx+N3C22cUvp5obkl7Rzq9xZuw+xpey9SuNrsIaT9917SQrFgU+A39Q
H8HLlDGDocUOnCoZ6n48/JCAzjoNHKZRknMtgfAYJ4qMj0pTdRwP98pD74Hj
pJSdJWQmWABSYrstSB5eo2KMvrajHl1BfuB6/k0+/0T8F6+9VJrKoeaALtto
PI6HihOoJlE5xASdwwqoacctTJMJg/KMik0GLINPQI6IWb0onRDYG36v5jAY
b/6dMM4JnKBRhC604+B/EnpIAdiUPMPjNrPzj5zW1+wEg2IKsKnZtW4++0eQ
qg0rnkaXmqV/Ek1Tq2e/s2xFstYOf1F8+8udV9qMR8YVaomowk0rDm+hS48y
pcz1lcFjEeGVvFj3yXmv8EHPk/14zATCJ3Vw1yTCj6URr74jAJF6kVx5Jol2
Ix2mJbJWgxiUts7Lejz3UxFqfZUKQbpUHbH3JN+Inpb4HU4QklVVvJEHaPAi
EuzqoYG3/KCPYY+OeDf+GTe/5FRD1wXrQSOZHnoxjNRDNnPNQGD9qFRowa2R
T+4W1dK/Xud7SmZAEdRP0M/5l5SzPsgmJ/UgseIWjOEdK7T+df+Fl4igXOKl
XCV0Lj5T57+bFVh7pMiho9zGqRsXxQZUuE5l+1zROg+Eqx8HT6xx4US4EaZL
tBXivZzEAgw/r6dC44ohsjYECHSiCyymTRTeST4LICxUjAshrCsk/XFOifmh
Arr4xGrxom0OXgNYABhygecbKzuY6dnhZVn/ejaSd1ku5MhPD6KPr8Ty+SQ6
A28aqoEdSx3Abg8SsEbRPHfWQI8BjmBLDJXOIzkRVI/vdP8xoRJ6QkQJaVsL
RhBQ+UdB/tcoc2kewS6qEmto04z+qFlO8WiWdL3XvOdmdA3fX3SmUYNoX7oV
mErSGJ+xa3plQOqQ7HTiR9ylgeutSndIT3nEOZVa/EWBwfHDdClXu+euqorr
InyVSvHpl6/EKvhyGqn+5Fc+lvM+XByGUTgHMjKWqAWXFcAssDiLuuy0QGy4
iULMgMMCHSoBvw2z8qu55BN5Nb24wCgzHet42uwxUYjCbjhJPO1oHhDVkOot
NtUpYuxs+sgHUJZ6l9NNFhQbUaGtSQVn7w6XAFzWQmW7blzEzPTgRR75v/0i
8RCN2UfdlfOgaV3T2JZr8PBguIQq1UjZ6t8IFFRP4Kk93Z/YioVLOwpvzIFa
MUoPqcFBkQv20jCmjhxoGxfjDSqTTpdS7+5JZZ8X8Zvfqkxcpksb3/jexUmB
IIIR2u8q3gCkupUXCc/QWby8VKUHiz6qGvn7dp9guYkAkNqKY2qSxjUvJTIu
R0CxAPEJx7Z5SlARGhhGuf4thcAQds8YtKiGK4PoF9HJPyjI19giXCRFi3bx
f3gVGrJ5V5C/HbgHjfqRk0IXPkEHJJ69H40Xw3mhk9Zvan63IbRDuKjg51iP
nblXColCAc2PPhXDONxVNb/HhmBn5oI+MtWVO3i933QIIVA/9AlaAPUkc7hk
5GsijW0pJ1zoTJ59ayD8mk4eGCfNJUuDV28DX9rWP8VcIROqXl4Nfxs7iL6C
I7S4qpb54m7wPJ3GxwY2JPuwdn93cfWBdoyxAW1njgtbyIDZ4ZSUL/p1lZBw
dvnT/HxpsnExd+yFx2/5x5DhJcfe5OfbnadrRE81d/FZV4BovgWS46phA03o
jIogS7B/Q3zGmozITf8bZJMgD6BeV/2MgjpqGIyhW9qsC3mw+hCty3IwQW/H
eAjPInXR6+2PGxC3p70IuE1uCJcJZpJbzu8dabbp4MgD4XuEagrE8UyH5tRd
BQhOAzBrMZzkGxCoCwCAO37aETeeA5t8jVfhs3ptjDCJkaTKrV7AAPFcMo0c
gXt0oE8YTNULdsvSz/KgnTodBpMQtJNL8n2ZX1oy7Vl/ie/IOMBMhW2oPwY8
iDoF+jlSNV1p/wmzwLbxU43oVGFHxvJQQzw3uaRr5f8cV3QuKwCdScojSlG+
IQfu6cCZJOMn8A2EVY5Eq5But41s4hs8hoxhFh0Z92xnc0i4azq2dwCiXswe
k0AvjpsMcGvWIY0xadviGQL9BvPESbZGCaK8XRSi2vaEsIT01alorBtGU1gC
Ds5uzGhT7+e2BH8R0FS49hK/SvVndG2t8JDrQUcOizn5Jc4HaTPT/+toKA5i
pNmVJ+kLlXEref4tpXlI0aRMDK7joV4UHsi+XO3G6kQhCZIEN5u1c4LrFirU
PD0N5h5ObpOFcImeGwcvMimFQlcQNNNPpwWYEs3hcYoEA9IyGrdieQUuPHhf
Yrh9iQRQwfLqRreNuEtV8BZafmgcdDRbnHUk62DHo9JmQGdvaO9YYSTs/hfl
J2FxUB9y5iohs16dIxAHAMR4LhRMBi1QXRZ0etFih+Han/tkEVqf2bl+NwKF
Sme/mgH6AsrcL9Sn2ajhXuJRedCU2zhGuX6A3FnPOwFS5I2WiJqycowuYi8h
FVwB0JoIdOhQolE5UgoDv0nQbUwrs0ZlarNYDAj+BhFLkaDIHJ6mpQhNxY9A
EtkZWnBxP4fNHwmSeW6zqCAf50uJhd/5vJrYCNFsk++vsJfYS2JcoG7VyjkZ
pVGnNte3O4o8ePE1CHsO17kVucMVGWkUGAFAw9IppRI/gh2GsR8B5C4e28HW
52ZN6rVWH/FajQpF+GTTlc6gQMLkDomC3Nh6e0QNcf0f9PeSYn7kvQ94ZmPe
BKP1+iqelrOejVXDSnVdVk1aMU1jI80LNciW5hKrbp6iNPgsPL2zttKNx1X5
Ro/i/F6z/u5Wr50BGJ2Y5xuKnAd/WZEwbSpveH4TQc4TrCAoGIRqLLRFPdbl
I7g/hlHK79UqNm2PvDViDRHRJT37HHbn6W8LYAK5jJW92aj0IHCeqhnJlCfy
SXj00DpFFxBG1cAf4hP9hfDwtfGRRbv2FkixOv3mAq2dpdwAISctVPjRxPwe
BsWq+PmX1V+XW/+7PMm3JnBfHYVTmFtgibincsCnkSs7dEIir9SgvvhPvuef
2CIjvDcjSpvZzPfwg7nCW1O3jdwZGrrkveo/DuTd4H8i+Ov1g5wx9H5g/e+P
YnwQ0ikCzowkHoI5xuWODGMtim97P6AdqPcfdSaj2A997AzORRB5+5cZTqA7
hWkKzSY1GvnAwAg+IFB4Am/1mX18jsS1w2wUOm0d/cIwe/9pCr+oZOgOF294
T+RYOCS0j2QFpKZTyBAxGI9Y+ixHyoMBJfDQ+bu/Q3Etm3SdKKAi4j0n1S7C
u5AhH7oYo2tP3iF7uVhnahk1nq43TbOKDJAfFa5FkkmnwafGJUCYtEHA8T/h
yjxt1z6oXlPJuhivSsHMeac03ya0S7EzNZOLBAEO0mhy46eGUE3/NqjfQqNS
47Hsnn3paOmoJtTqrTQ/cP7PvG3D8N9Hqi6XYE7n9RYJ0/CxA89ypP7k96Uu
E+I/XhtJ5rfTfXKzI1Cfv6BGD095exwyjQsig/hQtkFW4AmHCZnMs7yJO7kG
GJddduoexxwGJIQsT5pomhVpyteoZGRYMH4qW9DTBd+ixUpNtQtin1QEPwWy
u2AvgF5zWzkU72+n4q91HntFOmDEEqF5ZV+FMdx/uXw7IAlRj3Eqf78ZzfiS
qD8NVMbfRraMiz+vhbxtSJbAhOA1N7c6RLoDmj76qDJkeZjBwTC36bxKl9VU
9HHj8Jtt6i7woIF791AnZ9meGcQUNWA7UVrWC/V2wCW5sGYR3OoDncGbg4fw
hR82MJeB2e+wZXfzQxGOMpjO46789exFEzw+zORQGm8I0NmASwDkTe+6trC8
yx0OGLJrAsHWZi+loYI3i6GCmwyjFuMj1dO2vmP/Ao//MS3tDBi+e4QUHQ36
tOpT0wk0mMtrLQC2bCBBTG444zJTdw8QuU27CTrZQi1jOuZ99RE80S11yilb
bYsplXXQMhh9R4gfYIdoVXMjX/upu0RP9ANolX6SlUb+oG6shwLZe8l3qVde
/Z41MQJJLdMb5IWCon5O3rU0sEfCnqeZYm+1Gigx0A4EQ8m31JqRHrMq2dba
JdKOOWkey1lA16rhpq65Ux85UIjzF1F5sCrRb4zyzCxn4BjztjNaeBgUK62l
oR2RerRl6bkN3pqU5LLNlBM7rYfSXSe/HLIXHBMFoZtjcXPL/k/zwP7eNHAI
J9YCYbuXZhPh7BHF6+CLLbEZgtRpTtfrE838prwMASmydSvwvt0Qvl1s8bs5
znUIa8UHxAFbEk4r2OmWd0XCx78PRrkrO5IgMRcQhnaZMuRUjOCAQLx6t5AA
bvJFIoFOKUIPryX8ve/m4XsQc5uFiUlXgUYFPlNf+2oX6Bm+KpiPtBp5sdgG
RyWAHMy6om7MPJoETsE3uWZw/hg5NazsaIUJT3XoRKNC+KJJYEAoDo0Zyxhb
1mg2Z3+GcwbQShVWc/AvpWdqdWbXbKrQHWJZBaWP4M1Cn9uKTsXJT/8ZdOD5
TGbsLeaTvxhAjB4/fzOPTXPycPShKyt1T+tZWCQ5vSszPlRer8qrCKSrBsaD
VIvpQ/NAu+kYwFHxdPqmy+J5xq7J/n8JR2tKc53o7ZyIMJITSCi6TPE7K5u6
wVg6hTH5/1kUD6H0CIhFa5EeX1AUISYqCZ7LEdpWDuAflJcWLjqym7F9grKe
VF7IuBEqupEBeLnX3Pt6/s3G0gJ1o9CvUzAbqh+Ar1AN+qQvHaxcrle4ROIn
GfrHDEmBiKCPti4bZQc5EALh9Q1XJ2+fdZFBijLehwQh4dcNUfNwGZbIXNVu
+qiIZ8VD1NkR97LJRzjZsOjFh3l8F9okMbP5Ol675Rqj2kh1afYkRUXFAgNa
uhEhxqJU0vy2wLK/lIxo5gB5P7fr9Uuj0jyyAjRKFNS/Upd+o7LgXJq72Lu0
Mv/DfYgzTuOuTWIFpVyBJ3KuSdrs1Wmr0/pd7/jZj+DGtdFPwK0MIKPscXmb
96vgP0CkPcBJjjMN+MKxxjOnd1wI4zXkI0bo9Hg20W9dK8N5aguf0sQ0k74T
M6v6AfT33G475MDK+pek02AW79UIA1LBoc35L/n6lUN2jDo8GZ1ZjLtTu7uU
QL79+JJj6VzgjoYrCk0/cIqJHupmK7p2ll0z+CqiwwE44he+vv6qG+pv7WYd
PNKLk972A4VeFn4Tw174zUOIiV8ojbn7PzZZ0QJuScguleRb3yCu/avywlPF
/Da0EiRjyY1iewcBVhCRjbkyMG19p3/WXcltGuZ9tA2td3lBN36WrADid3AS
NuUiBmAPXHpaQodxXx4GSKXgNeapELTvF72T8Z+3J81sSL7O1jEZy3EebM/U
ZR0A5kixLm3OTznia1F6jDgx0bs+wnjsuCsN7ETMPSH25T7FTIxoo0ia/bi6
vroNc8N1iS4TosLPt6PezR6stWR2K9jBnm+cIRU+khSKgMK3uyqt71kgXDLV
tkXopgI8r+W3EtKUkq8z0yvnfwnnDQdorjyINvsZVf3hten6VOYEZCS0o5eU
0P+SueRWepNQB5mTT6/S9koaS0X+9tIauMC6CeItocLx9rNOg2f+g3EyQXAI
gEIxh8PBBhfXTgIIs6B9dQOk2szuDoV+Xb9P16lQr4KaV+1XCV1cO3GQNsOd
GPY7Q4PfADZ2tEEuupaO99Bb+P39pwkqtU2BLPOErPp1YIRSTgs8Z6g5rKrn
pvtDiV67iNAMC+kI/MXb9uEk8miUTed9u2ErsKIu4IZ6a3C3YxkDWyUtRYTC
QPFjvirDSR1kuk9VXlFhrncDydjPjwVOBJyDtBX0hYTD5JcSjq1dA5KbvrV3
WFmd7RTwpsYHPtp9Vcet5/uEaVuU67FHm21vbKerr4qfmi6cUuFFg+YvpLHa
vDTyIHeZxuPwheGaSmIvko4Pbf0l/YHwEczMNt8zbZOwwMpD0hwwcAqCGoWn
csSBSIJGrckQutYNZtdmi6MMlHEp1yRUHgcLLseteh+Tnp1Jp6r6jR+2rQZ/
+Qi6z5rdUBeFKfNZuMc0B7+wYuN3mIFzBpXIOKLoK+ZUzyAx6qDDOF6reOzF
IW4ZCbLn0JoSEX7e46lVle8WxreVilWNmybputuOilCs0y8utr14x2hfujqk
f8fljEh356GQEdgmJJ76IuTuLlmI69pA3kxQjGoZCPGKzenTegEVhRTLr8v1
hAgXXR7t9HBdJxEFkMjdZOd8Fx7YbIoIs1aF+El8VZ1s1LZa81UemysN7zAh
rSJCdP//VXCckhftS4SRXM4FqNwOWcAQ2sYgEDRdpNiOvD3XMQRf7VwR0gUq
leUKMa7cPYXumCKls/J9ch3tlyn9FC0ridOWHvpNWyCygcY3USKso/nj+1FJ
+hyE2NzdC2nUDHFfn+Nu5RLDjxfCsIBEbFHU/1aCqc4EJ0ztD3UsYUyvFWqE
vWA0jA9FAu+BPs45H+lktwHcT2KGs6YKKXDavqGa++ZRscBLT/8TIeskNZDy
JrEG7srSbqmNCABdoJzNF0PNH6gJ0Hvf7aCwQFktSZW0OyCSKx//g3oFDWLM
KhTLGMBeKLaWqkRozr6pOV8fURNWqg84hQb1DwVpdO0A2hEaIKx4pOKMtbHl
/I/jNVQn1GQ9OLDnlsIwjjPZ1hmxhr4J+11t5sCHrsDSTlRvU6P0cWfb0kFi
7n5K1hFJKGp0aYCG1XNRQEPg4Au/3hU8eQSzy/mrEVM9Fk8TOGF80cgL4sGh
XJaygvcBN5mbq2jmePlkUXFEkzWvx8KLEMa2456XLr4BOK1ihWBMnzKT2mLB
GgLTkLkEPuHwKJ9fCLAqzrDFjjT0OPkion/csKbRdn6VaorRcuofwYJrau9g
5P7rgCFUcMYCoei0z2U6GnyTvZC9tzBGyzv8Bm1EIT+VuiqlzKCdgltlJ+oF
wp37r5tEmbEHewKseZ3aPkCzCmhei3JFwQGqt1qAws1NNG0fR4CGeXCn2iqe
EH309nXs0YwQvbpNMsA/nPpvxVTcz3kzK8hvh5FMz46RsCPWblYjfxSnhpHb
fDD2ObW8ypqEMl0uA9kyN7JbP3i+46S2YP/xcucwLJNXhqpBPuMaCPGaT7SO
cSrnsXxnVIZIKd3fOco48S4OE5Ncgwp/mnsCxMu35VxXH2fS+TIS1ZsBsV80
TDL0fx1wpkLVpcZK9JRmVJuJT2GhVoYVdRnbY4B3nKyXIcLNK1Rzrq7etnT/
Gq/85mGpvwXgoNu+nzSkbnQl19OkKgVL4tp/aiDTNvklYOYkqnGQAVy1L8kW
VFDEbgsGW5dvLL7avfQrW28PypbCH+O9Lz+PARdQ1o3GJ13relqf1mDZInY3
WnYg+nXCpzYeXbgoidqan0CD7mTF7DKDiIArE3DXBSPU7OH/2WREyxEve/cU
gfqE0fxrjIcDbIYkLKa2kn5FwaXjuAnfD+KLFxvteXPqlJj0fZ6vfaVL9xsE
bolDbf5+4r3eLlkr54KCy3tK4IA0ogVmg2nK2ZamI1SIH/5TUVtXB+Lm1tAk
YvWbquphsSmAkUGylD4327viPHbVRPcoSM1BeRP21+yvfymU0gfiydVaF0E7
Tl0cJNd0OeZ6fw7mMmbBKd62G4i/lAwwSrFUasauelZ9xySE5bdShMNYgKfO
EWFmP/R1g9NdkCCyD6gfJI/ThZl26ufpA9g/BhHhnkESeqS7nCas55tTFcXN
MV/r5up56g2v+RaUILmF0baNRlvROO3xm7vCe3HCEdm9txaRGiqUG1Jj5FL+
gHt86L6DxQj7lnAjBl15AXNylZrQCzfKvIw9YomP5mkwtsFQD2lbW1UB7MrQ
Jm+b5sfBxSJXQltA9n4+XZ/mKP1ASNWhaLNxRtg7UcHx2gA5XNu0gMOSRN7S
VicU5RUMtcDe/ZbisJrqc1VR5WAjscGbZ3xmT90watA0krFhF9B1EgZnCVE2
5nmfTM/3ZNnlJuRUBJZMbYPtWP1vFLi36qx/RsFoKi6kwzcbIT8qvRNx+JlH
MW13hV0MX4bsu7o8aHOJKMnHq2kBExlZLYbV+DwZMRVtF5Qfbej6Lj7cXs7D
vt+wy/502kDzWa2hAjsgASc0EvVKh7N7HeWx397p47vJmMCvPYANgLJcpnBl
8cLxRX9CJkxtTU+rWWYGuGcd3rhn/Z7xPPyuUaX6JXihkgPBKKLgNgLixvbE
XI04ReOAtLyGZaGu/NWQxEmUDfoUBzqbTC0aaQqdXiO65fddT3wMtGgq5BNu
23GagjzbKMQVMsa8Cu6Jj38aTcVOb/UneHWi6yPiACfU/nNMqhDuJv3MvhBA
FJcI+izMJuogpxZ10/2Y0qn1TnNPZhEryCjsatEuH6O3rzEUUrRp7UVJZXmq
+kxfrladPFiEfEMriW9Vd9NI8CTMdVqu2TPvTSm9sjy0f67OTVPhHy2a2BU5
XHZYSTWvidabudnQjai5YJTy7Qkajdn0UcYpEVaor/v3BP1Q9+6XHs9cM8u9
0PB5EgxG/UnGE/MJa4rHWTqZrHhzNSFtP0BuRuArA4lntKYs6zk/SORlu/X8
nt3GRQxAt7yFaQURcDztpr6EAZ9a5aH+zYjCGDUXmGuQZ/mwqgkCvivd1+tx
WrZ3AQsK+PDcd4LejbPlQ2Yz3H9v3RPHCxLy7j9Fx9syt7KU+t80HZfRBFny
Qk08XcUh+wafej4MRZpTJA59J/2qnJFIhYKAzIbXjMBxc9IktutVDpnH0vtk
yKjhqOhL6GK08ImAImTU2dEJA2WBdzAK78hVRHjANxFQskzXrAgB7mo02+we
v0vs6zmbmhPy3IlsQxbZptXj0vhB3qpYWPrZWgxwYJTW/DBJRT41BcCsnsa9
ZxbQfUhZAWlec+eii2GciawtVRL2lsJkqW13nucx1nQHlNkcOvqmOzDUaGq5
uuZZtVTW6yT2c2p67Tv0KFeLb3xlKdFs8J5Mditlz2wMjmceOFeGMROfmhDm
kHn+90hfpIg5jdF88ShgbsvRATP5Ru2Xc+iMfnn6zWrwbg/2xfQzzgohhvow
m/GeitbfnqIlX3dAWZvURBfr1EvaOeu8oAGzLn+cTVYCBQ9MMtQD3DzpU3GO
/cV3teUMDlpV6cgNi5x4gqUN+do/lMc/kp5TxkrqEYnxRU9ORr5IwgTiYjER
FYdnG/UPKreagCWFspyX4BccNRibH+6TGAJCd13Er8AqkloeiiYQsgD7fV/b
wQ0kMhnciik9xl5RnrWWQA2AnpvdoWvNdB9CHZjojHdRp+vME4IYuWmaOup2
i3BYocZinla35byCPL7wEQYgHC2GraLmQH/S5TnhyQZl7y+MhRkK4QrNu8SO
JO00jcP5hwRn9xDzUcZDtc9m5AcwSthvj9zT/rGmrENpluCjCWNz8trs/O+d
LcoBYlMKw2aZndVGuvegGujBa3LNhPVQ/tXQZI8g31d7En1oqDrm+zpD8FKj
LEpsYZQZqUzfRgIip5/BenNRFeUJQ9HaRBV/boeM9+wvnD2Wj/rdSOP71P8D
kS44lZSg45KEvcFROretUKEayf1H0eexyoCksZ6pPiXHjkEYUmAtPgkGA8Lr
SNXqka0wp8sX5QCuhxysI5nawGla9MxRjB5RprjEOVPZLCH0y/Ux8LYqeZJF
R3LPGpJ5GJjlVnn4ka/deevgaHPoqOB3t5XG4SLnXdeN73NCXPsOqxa4BcCy
0hO8zHM2j54NFOt+OxY8Nz3g8Bt4bLX4to5rW4/qvi1RE9QkC5yiGVowD6O/
b8pN6qcR5EXLUvtv8T2oJiv8cNLSzQ4KaUcwCdBqmzpIFMRyQiZ9MlRZdNQg
ktdxeeT7EEaiOzQ3rcbB4J3ZYRzqAJeJoB7LGOGCkm1oPr3TeDbZdVFPaA0/
OYoXcJAi7ndsCXzFtg+6WYzRmPZPve3fCRIOaZp8DGH77XDyFayXIQ+kwtBv
+mZWpN5O4KZ4kneRJYZZiHZjrms6Ryv5VVOC/E7XlLpGXH1Q//bIF6krNLIx
eNo3OJtoeMeQ+LPZC9aksBtqLFE2hiZ8NyU97IdquenX8CTibRdopz6yB36l
iejVKF4+Nlq0PAr7m2bNGTHtJoCEEhFcB3SI3Z8bxvXMNMu/6y55P1xk5ljT
EBY+rHDB03m7spUjkfa3Shp7koEXi6ILV7dmyclc/sF5bWqYSZkZQjHNUq3V
rFX2HokmHCqAk07gkO3abFhIrgvFRgv34/Nm6uIDmOE48YgyF1aPX1pt9g0L
inGAWZV4eyo4AlOwndcLVzkvspH9dtO/CH8ZYzi1++N1ER1ZNpYHKkaq3KX2
8RuHDBFWmJpoPNlXiFIuj53bIGHz1J4QJs6aAZwWdOgcOCky0kFEKaiftCdz
aHoyAtQ4eqCy8r+Gm/SHXiqXXMIWrbsZFJUUI7xH2R7nbN992x22HQl/22uW
/ZgLBVYXZVRoSScSNO1ktBzXac54Lr/zj6vYm0apa3JeQXUv3cdX7ZbrjfKW
/vpfwEd4Pw9ATSK96e2AiDUltvDpcBGI2Dg/4/eh7GZiq9n9nCxQ1xMSDaeU
UtpXgufaPTA4zxXLLV6YfCbQOYngQ0nrsyq8oObP9pkdbHjVuOahuLbpbNqB
YaVMkBTN+M8EIWn4OUcwYV2Jx6+ocD8r2gLwJ2hPrXl/bqD/ltdbAB/bXTtl
RfiIbkEnhAM7hFN4OCidobc2ZQC7jOwNwS8c0fwtUMoTeLNax4A/QIxlXsrO
H84lhjJpSks21lHuax1r72Z6HKH1t/pdUtKEzZfEg2Ct5PGuSjuKxk5BEuH6
NMn8rpiUuu4p0AaWoIHUUgp/99NTQh/v7lH7dPumh6TuxrcGWZ4RyhZ844Ei
ywVM2ytBLcWdcxLxGa3n271Yp0r2UM7d50ktlaENImYRJNDERoZDeecEUMPO
TtulHCAoSNRbgh1NuPpRSOOS3DY8HY7yNsYvzFL9snNLt+7giA++73aY5omS
82uNPIB9MMOlKucnGFP9RnChxEZHrSS/wuShG9a6EIAZX8zwXMsZalFq/tNF
pUoEFVK94SuymwAF+CEYe8+MQVYs652UQomiYLnmZpziw338nM1HGyAQRWuh
7OvAo/f/rllbzxXcboMM5EvRv+frCa/4sdBIDMaj08UEH2O8lUoL0yXAf3a8
WlGI2Yx0KgUE+/62p737fkfQmN+lzsMrLItqWPws/WWiY1fANp/MfiRef6kr
cYY3HSQwYKnqg9DnZpaG8RN4sWu81SOcyr/UkjOkrhdqAGl6e+JeL1xIqJ9V
ksZmD9I1Km8QbpL5G7IR/4vntF80og39Xc+vJiHKd/YPaLC3rl2TIpbX6t+s
RVh8v0Uuba2dfoezyul3KN08btr8d9gnj/kRtyg38bdsOrx9DlbZViZ0ARI3
KyutejS+kXuy+5fozzlvs51Wg1w2p+OEWGzLP5KeTzu1HRZMhXYrD9eTmw1i
Y3JhDtjn2RRauf2KZj61Nla0jYuzhXOhEgogYGUjwJyKZvG8JsItkehKS0ue
dJePJ+mafg8n08VXki3MLnlVFl0srhw6pyNfRhVowQ5kXS74Of2Ki3rPILwu
Xovzp1Coavyz2hXeOJOu0a6dh7wCSq+WNJbQ9LSHjhS06ZZ0GvtNofADdIky
gW94/kghZy8QTd//Q/cYVz5rBuxxd8sjAV6OKt51qMAiqvzkuwpr+1ocoMlS
ToAATDXDYCeI2wld/EoLKtWpLm6Zo5BOrBIKbChtCNwpFU6tFKjPYi0a6M/x
4X/OhxhxcP7CZR/SOMPNI5jgSatbYZUBwpo7/ZtUdzhym143nooAUhRyxLzx
eQVyePbna4tuXXMh+v7C3U2rWc9H2RCbKE5HHu64PfESyLjEye+YnqxmnhOm
3k6loss+X5mOcEPFcbyCFlw3kCbZeeX/5SUti2XtDdVTJWBKSoOGro022CHu
LDos/6VYqAFTD7Ye+iCI3GTxry3NuJuZlDEr+q4PLPYlJBgrHCVnYEnFUPgM
QjWS10tBWgafdBnyy1ETINidwW2mmcxMue+U7OngfMHj5NIOxzF8m+qHm/U4
XeNOXXgoMkH76CsQMZKvLDik26IRqZUntN81mgm8M3GE6YUhS8QAWE4MXs/Z
vyfcEZo/2ZhAMaXaSSeoPeNM4i2El33AC5ydJl95inoPeO2sJdfLLJJiSnsO
SCJpS8ErgKWeWiUCwZbbdY0mqkDWFeIPSxvxcQ0Y3dFOWu8mcx9P2H6fEJxn
4/QSH9RLFv9nOyqE24GvqPZ5IaE9A3oSvRkoxHhiY4Y9OMZ0yTN8xry558Sq
fWbghYbhOWZ4A2alicHqzkOwx4aZ8p8m9IS4PDuCfs9BV7FOJQpvqYXUEFOt
hxUXDyTT+ElzDDn5/1b/zhYxgdHwLDNNDYchHHYzSZCM9YY5dF7ErGDOOLwO
DQgWfzrTz2VSLmqfJclh6oTQl3u4wZCjcOAAcG452YvVqoE6Q1XgGcsFII3I
8EBVbAxyyQfHdowV1jQKYmDBsPrT0UXXXQCHn2a2HOi04KDpwBP+ZLFh/4mO
SfyCYNOMZaXQC5/gAr+Oyi8zPfBZqIdhtL+dO6wZq5/DYsICik4R/wi8Kh5f
/3TnHfzs9dwIO6xHEZ9nnlcr2n7i5We/kEdpeRdSWLqjl4qh3zE3At0X7zSG
RGPKYlo6lBdlHydqNJ7ZepZyxd0lBm/0p//YvT+M6zEcnhBkg0BVEfoY83tT
fhSOtt/FXYzqOccPBhvxYzMLAtwEeHjXdTDpv7ajFUxxWAnBW3m86Slh7lh5
E6KhSCoi9HPNG6cCRUQ6YmJL5vaqvj2AU0voxXokenaY5qvvQkBh7UQDEIVX
nAku5Bx92rbvczQ2yd7s+YMhwYcLtRsszWmQM3KcTOFosrKcK/jEn3sXKcUM
QtRPt74XsC3/LuBxtvfxdMd2eIfTaCqoHvhg5ejXlfy9y1E42uOs9sbdtPsQ
Nhg6jpsbqLMAYb+Upjd+uXBF2RVOtg98Ckx5+cvI6CFp6LnU8ACiGN+Nbv3l
By2UyaWEEVq6r45vfTyHTa3jv4axAiqSl6dNorlgApVO1y0VlKlsNeC/con/
pXgwfaIZfgWNXSBRHLIvO30YN+MD892g3RSMUXGBlK6nWqtGBFJoTUtQFpTY
VX+Y+OZ1io/fG1hxmxRgaSrNE6J6Qof+8Q50wCmkZ96ZJw28ZM2hOuE/WkQ+
+cq8iLggCd3eQbVumA2ZIc6DWnLY5WWHeFHQaq7bCUSDlnCDk0orHoKiXmzn
ip/ndDXrBtGmEBiMPYeXOEdOBhLorARtFp+YxP35GJ6tOLbea3z08GD9SHhM
2AEg4q8vSRMjrI1lvnmX584qjjlSuA2MQAwpa0dbFoCYH/7i9ACCFGWGqVxY
z/YAu1dJ4H3uVjLcdYT/k8GOGEzZEoCTaZ1aumF8aEqdKA4fmIPm5jCaMS5d
RmWxlkjWaNemsyxFEv6iTH6mJwZa6ukJ5yleVQ477YBKU1ero/fQEDV8Og/u
8mRuhGMn+wKdrSzA1DJP3oDsUiTInAUHafuYBmXIMn7keT3q4N4Md44YGDx3
gHrt8iQ3jrpXPK50QacDAan+/DnF8GhPzNnfNE5jBmHlFA68gp58qxElfcL+
Egb/cDuVaB+QXPbwc6qGlv2gMQQmSLX7AfsGMjuJCighVI+siYDk00nwQjhn
8ZeCXb6vaf13fHfVzujI9kmYXh4/Nf+v8P7hRUDVcCOiIaDIPoxqJQ7CMJL6
R3//Xybk4ktV6QcKYZb3laLtWhyRWpt5BG5t7HcPaJj0nqhplbVyD2aq3W8/
+qKJsS7UdFzrt3ywH88q2IXqRxfd8iSprccvL7FCEpIG1kh+R5QcUiN2OerQ
44OXsk5YGusbEVyE4bcM/RHj6yB3kiYO9ovjBVCl3U/KxmPXzEaWJowMTUkG
XZ+np1IkjuEDv8ieqKFBkf/p8JDn0+dc8lbp+G0oE0iagAyrT/sDU/eQsgbr
lwCmq7OP8OoC1Z73qoMOiyi4lVN3JC1Kq07mjmr1jTzuhaJ9vL+K+ZT+2G/h
R4FTz4EEgmwTJqsNKNLTy8WSVHunQ4Ed3qI2JO0x249008jKR45ly0hOXUKP
nh6Yg2puEwiG5jYdpbVLwlkEwc7wPxfTXdHMs5RV+YOyHS/5efg+BjXc4zJK
6Y0/yK9I10B9J+8knZJPxfOJTE11X76n5GQEflwndVV+M2Pw3h22rcF6HVz6
R8ljA9nt4BEZEttzXXc2aOWTGtcZjNQzGpRZgljwcD4tFNSl8g+7t1jrw86w
GBQ1u8qpmYLMQeGN4HC1BINFMX2Zr+5BWJpag4y7J7z7kYgwFtLD/D6lHwYK
ObLm7KahdohU0LrUYT8eD+txK2ApaELTw/AFmtOu2mtnqdzzRrSzuFMkoJnO
NnQrdJqPtIlprG/8Rq3ykvlrsknRPwPedKdhPu8YaSLWA83uTHwuRaNjqz+R
hX2QVpLK6oXgYHvVImKUGf1Dgbl31cUE9i+0qS8PeJmcqlnkQMVYDj+tFpKt
USroODdZJ16GgREALwknk4aTE/wumw/ZH0RSityUrutk0XRYwO3uHcIsjAGf
zY0ymzNWi7RxMv/oQXDHiWWPsgFX0brndSACNitxqFLREagff75s9RZVb68c
tEnviVSe5mFExSpv1GxWs0+OXdvX3OQoNMB0ZHTv0CTLuIP4Akj9CS5N/h7v
TmqtdRMKIKf2Xgs3fj+fzXZlIAgVSbgLFhOHHCq+B5hK5sKbYGqgwhOT1vBt
nIkYk3XdUu1kDlu/rqNcdusxR2lJdz6rctUI74iAZrNnz5hU5QvZS584CRr9
FZFaLitOtt/JqteT/dj7BMJbNGfFObWkJ4i+3B6PZSX1+KRjvyclmrETZ9sI
EKfUTgAZV+pCDxtvC64i0ZiS8DuiXJ2g5bEOpzdtks63zzUbzxY4jj9gL1/y
7Si7AInvuMfc35N1PK7vB1PETUVn3KAxsz41VpJ9N0EIlYPUPW++Dp1xsQwO
EiaW/gkAt4nam4/Jc66Ss659TOzRhqEN0El6ZnwdZhq2OiYV4HtHH17LiDKI
KT9AFVJjFz6yNoUerlwZKZaUtiG9TZv6lM2+I1SJZzNfp0z9lGR/VucmkbQV
rpz88/1eySuYsNhMla9awfLWbjzbY7ENyhgvCwMUkuvDDsX8K6LSWaKudgbz
LJngdz2h5YklUT5RBpw/AcBxZ9A0brrPwxNFhFbDYlDMK/xfosqa8CfwVMcE
B3sWrjkla0meq3d4ICFafNZbNBGQdapJq0UlKGs0jicU+WEA8ULRSFk9AlKr
kRMCq50s711EXxTCaA8KtN6MWtOGcOPlgdT3sAdaQ7KqwEt+8UsBZHey27uA
RmcU54IVslPkEra+tPDyJ9IsQu9FdjEpJeUc0Nr/F4fI0nwO0Yy+ztTrodiJ
l12i0PdgMcEaU1xR5OdA5prllP4RwnkPKxoHesEHL0NT3W+dqqkY1RjP0lPS
RZ8BHr3T46yeYS+I2XMXfWgHLLyaqD2iNRrv32UHAIUtCy/ncpi1LyQTLb8E
qfWbPVJqIrDjweq82ciTq3bSLFyxgZPa2jMy5n6rV5ZpPX0llmFALEVfG74M
hoTaDrwf7/OUYFc8YVUCDy2Weyy+nk2GXPAitZb0w0UBrqjS+06iONvOKwMB
28ChGxrFPbwzlIoClcYDayZuYGuX9NDov0brrTIm2Zohv0NHeniiKT04EI//
ion3g8Dxj5AoYhdJ74CUMNR+7We9uRsg/bLZ5NxeqXM1fuVj3CsMCi9zR8uN
e6NxeUvoJqzV8Hw9Cv9doxWmTUXj7wBWy1pL647q8nwr1ER6RijgzQtUHB6S
VGvYLWmqRnMq3C50FuOtC7TtW9mS0y1Et0qAHf4CrSGfIaMpsNivJOh1EqLm
irazDaa1GVAf2E0eA995HNKqKfJYmPraBYmQEXxoNXVYOWi9yDWwsdeaxy0I
jPnZdwtBuvIvuRs2zbrmxLPtFJp+Iz9xJOpY0tNctGUb8rfFhX/Hto9O2tqd
eVD+dOn6+u2aYwYS3yVuyJNLeemexxSJ/6CT86t0KVvPkBSqwdK1aqOEKFeg
p2d+aC3gdgPRzBedqgH8pymDOTj37SgPCAJBqurgtn8BDifRU6a5ugdvE9tg
qEleB8Da9GRBAIq75wSNs5xWR4gOkJ/Q22mzMbCIqIqUM3vXZSNjRbHBysF5
cY9EFJ2/wO1H8CWVGt5wvbH+dX2marwF4Mx4uuM/o2eWB0zJbkQlRe/vPhcH
otPFd4ZP1AJtdjZFb5lHtKDz6avtOG0flhXKjkXIZ7Cn/DiwqFW7NTBu4BiM
3ERZviUSrcYmWG0XIcibbADxihrpi8wTiNFAGIJX0PyUCzAt9hqsnvYapgCR
XJ0CtxJ15kYyyjFt2n76RDSUVczhN3BStiyqM7VjtrArSlK2dkQfkbSLQxFq
/8DP/s9kE7QTG8HRS+Epj8UMMUopLR/hXEdbbZa7sVvR1Hfa0yk+G4q1z28k
nc9YTFGDOXX/bAAJYawZx88YGJpB1w1b/WsOUg/QVWm718Sr83+rvXbSa6cO
5ZXoDaaNCnFiaWM7jYBt2BET08l5VeYbiksD0fnvaLe+k9XgdUgo3zIyL28I
c2mYvlNU6kwQaHZrIomGjT4XTbejXANCkmML++M886OP3TOtSrB1fVmCSmC9
two5i4QwO+FHS7v0YOezE7YwbLdwCjgPFJvejrmxeLss8fTFYTRbhzBcbNFb
NMNc5ZQrhjK9fSxzJMRgB+VHX/97OHHTAFh+Vzm5DGN0zlg2sWdSyssPpVXi
/hzOf0IMoMM8K0WD7urmAQuHeGo8zIddi/QHFxJc89iK8jETHnd810bC0R5/
ecqUJaLU7S/wVs+NIWqdiWjieJYRxpxWxZ5s7WoDAEygMrjMZrf3/fJRs45K
UjehKugRxubyyBWy/qO0lEadQOidl8AMncoEZrgDH5h9Rt2ZqQ4eoW8rX6FD
B//5ypdJcDOUI7TawuFPuVEulw0JaseBCpiQ8KqXHFJ69I2iczGVJ9W3IPV3
jnApDE14cJT76jAW8FfE89V1xmDqQIv3lomMsjcnXw/+SA/+FbbS11FOYjdZ
hFZSaQ6/KO0HNvlYg9tgxhFJ5cP+YHpWTHKKOFMQmvGs7NIpscX2zfuKxQSh
O8RMOz1scfgN36sOqEaamhVXkkmEkOEamQZ1gNYgSHGIM5ev1GqPnozX8pp+
r77SK3zEEMVl0yduxc0J/p3SEzVtqT+UJKWwJ9yBR1m/yW0f3ZjVgKsJ3Vjl
rGfGwmG1gFthq3DaW3hqooYD71KXfID72NUWOM57NQ22VSkZvEJrukj7oGe9
i1RFqAsamnbjitdKO84oirVf2UUuYtAvW+qzDoml1yKeETYdJk/K/aXQl3MB
oXmyG4Egkq+yGLmn4It7xNgqeZUXaAGSmDlv42oxPbZZvln0EafA9DsSFDTG
EOQl/feEB2fXOGoEgsBHtfmyYNNjGysTKspzz1Ta0PVD694kvgW71M+YDLXC
CQrOKpOhJ1zHVokT5Fn2/19y6wxsI/f4ewLhIxaEjFkKMIlBiKJHGekpF2Q5
VUdarXSTlqCjHDKwhKeejjf5tv6cPDHuZG3gsvTAJfajoAPnU5wwiR3L0jVd
FnnHy6wdU+Y/qofmsQRVJtyeLKfIE/bLS27wUPikDBJNlSAICxEC2I1dsZkJ
bTMTCH+4VNGJP02tcA1QhjStlwPO4rLZKZz9BqipyzGKqJM+YDx7m6oR+pSv
6QvlG/1jTBkwBEkajlaWAaMw/C7mkyzDYKYb826wk2geCrYRv98iu+kTeIup
aatKEzz1MAmNbyaBk+OmW9aoPlOE5E7wg6bqGYdTz9WyRYYSRtyS+3CDdokF
Z3KvyDwK6PpHOVpQ82wMtqi+pGEQDj2dY9nxOSLkGvkY49SI4+oQRAvAQtx4
8NrDumXLU5FGCUBwdzzqlys40NW67jcdjsxY6erTFSVdsutUGEc6vYCv9UuN
GQPPaUHsQueeJmaS+/Im0Fs8i0+mAfkUH0sxFObnnb9gfyZgNX4Sh4BcTDpX
C8ENTPIMGPM1xe3IFfnqKBsRzNV7NJD7O2aV+y1ZYgFZYMej9/LCmw2h7ZaI
cRmDPoD1bhPTXwUURNLBHjlW482cyujZr5rNNJolHhbqQJSZmtXp3gDJYDPO
SpIHCdh2nRdw+qcZN9m1YsH2bZ99iaow+dPAyZMbkgBbniDkQRcFyVw7jyD9
6zXOEdBOCHYIwj+yjPFzizHggekRkE0C8ROOHruu7QAfHSmt2x+d6f4NK39W
7NybPTwGetARvfodKzDls7czpXnZzvW6HRmjR2CUQZlbxvOfoiTucASCa47L
jKLK1seezrurAy/mfvmbZmpq4ZE3V/tJB1fFpegePMUg5HojGJu/vKQJ+0qR
xKNF1deOOedw85YUg+bqRXm1uVmzq51vesDMl6XFWtOBgaEiBEgjUDbY/6wp
I6w9Q+yW0DlSoZanZeNL6tGUyoj/GtBakX0H2pSatcbZpwmWkobPq2tsYo3L
9TNX6i5FrTABlmjPQrGGQOSLmdSdYexoQMwwvwvEsTsvEqWrCkV1UJ70tv4l
LTkAoc71sdnN3Yclf0JGcIJQ6ovmvNG6DBUea3tzMsizuxL7Gyp8F5/uuFrD
7/AiFXmEfrfy8dAepA0r2/EiwaCX6L3fDpom7AzVIvHx2M+iTL1RdSqmzGuv
usv7/dWnU2R8a6EPK4XqG1PQVkRo2yQ4y5GwgqN+N+9q67VvaFbb78pM2Zze
DxXYQE3cSboQbCZYSmaBznsz83khrOocRmalJYPT+D9HGXDE85oIOVGj3Le2
qmUXP9Mndw9UGm1R39XU3eMY2rs2rQXFEBjgKazkTps8ewYrgoiWaFMnayqQ
gXp6GCgSHn22Qe4SYx36GQGjHl7OcNFLDnXIwJHecQwhzSUAQwQqMBcqoRbJ
nGKpkC1b/Ht3AdlarsHTeaVOHvq7jDpUxrsW13LU02zFQBJNTZZCpErkVvLa
WWmc3X+ZzY76QnCjBh+/P+oykLJ/KkxQpiDXIjBf5Y473xn4gvIQ+PHdihuI
tiTjZaIsg4sSwF5UrtKyk+iCDR70pnxh4UmRptO1Vl6M1YG+yr4vuaJnYdOo
hs/ialyx0zO6KZRwStfS7lLk2Nshp4ctcoBF4IXWhZZa0+nqnWvUHex+oSUM
C2QeBziQMV12Un3+PbUnULVEkfllNcW2lNtTou1RgkV05XDxBhRIXmx/84Vp
yY5vCKWfSCl933lHMpeUa4cFgEJv/4ThCj+/jRhcTThjNwH5fGZCpc5UDmHS
/4uptC0YPYXwL4czn0y1fQUQbC22NMewdftrAOBPwaDk4/30s2y3BkpMZa+a
H8zG4gYKs4Xa//q2n6z568EV8FV5vNtqGzHCEPJvgink/t/y1HtdiX0FQkTT
nVNJzvlzsYcX5Y20hV+UWFKPpex7ZDCLuwPOcnB+Pn4bWAZSO59/7UG4tnlM
kA5rHskuelDX9s3KzWgNGA0/UEzQoI6D1vl0moteee2pIESal37jbsV+4oID
OAtVVW3OlHMK9m3PmOmCM9M0xdrEIG7s082ZfTjwZKji3NolelToOPv7vT6o
r0Ul+LTUOorAgD1QUAf11Pb6gpVeTzhOM4+dalo5LCtFySLwWQs/eP/kvmV2
3yvFuzOutEeRPX1/ovnLfOF9+h3nkN+kus4eC3myVmcVz1zQaWNenQmhgJpy
6cjA3McSBKjfKInQbgysPJ3u9A9/AoJAX5D9nP9dUhlxnVxJSyVO7mmY3mmf
4eEUJg0NUKjdh2juvDEeulp83celprzOCYwiNMR8EZvLCY9VC5rZmHEWMdoi
oizBrBhvgrWasgwfh3/dn/gHjvb/YljPLO58CTcJ/QUPHn0c3AzyUAJ0BjEp
L3r8eQEfxQMBukgV8Xg3dzF39MW8dwbjd8S7czxgZEZXWHjB6Qc/taHj1hrO
j02HnXZ8kuM+9WYGzlTToEQVdyS+ZnH8nvD9Nhuio++t7HOR6WcSuBJdKuHo
8gXqVT0KLoXlHsjI1/2sJV9pN1t1qS3JZrvL7byYgRTqC923pCUrod7Jh+ur
UlFcJQ3R3PLD++BWbUxZ0AqVWbbpx2XxqvxyJGviNSvi+b8pe6NXqwcEyfaJ
EufmRviytucmCgChQ089KQ4tsbIQGKr+/g2AN9KoT4YtuMCoihb4G/GFpjpG
01ZIbD3s81molo9BqiN/Os01Tx+vpmAyrNgaSbXcdW7vso4Pus8TTMl3FTtW
5FG2AI1gVXyji9WDTfIIB7+MlhAUzT1YmqCG/T7ehQE4m5gyi4TIP6BBIfxj
URexH8gCz5xZfDcB555LMvhueRDITocSP0al54kgVd7Noo5+KHsqX82UqyDI
0XbFstVSAWogeToPKjsaKHY6lbUzbX4i1kuDnmec/R+OxR+Teg7gakc8s083
/eIThoqnzK0poHg1fm56GT9xq50OjA8sWmyASoFRg3M7P2gwANAmJjU1Fv/a
uzvIre7icoXgcbl2uUJrCcJRrupoxm3/ixXdtpKT9sDT00k7qiiUquLl2pSt
VLvhY0hsTlV3HAWZkI0HNX8qjGe7oZasGBFWU77MHjDGoQaZWIv1yJI68DC7
vrRm3N3+dODrlD/WybpmvFDAa09fuP0X4ldqT4RGQ8/npNgb8Y/qVlfUwJj8
rNLFxhws2kRGcp1HK30OIvXEellGUMWagY8bI3wZXOrPddZgSBl/HGEQWCzy
tR/9qwIwH7E5DexPt+ljcMIq4potb2hfsNr4PiQTpEPgpiKs75cJ2UrOhfMV
sv/gqu0Gy3RMbRHpMz1qoL3AIz3wRMieFzEyfdXyd1nE26tzCJupkTDUZ70V
TwVzcpljFXk0djIX1l9Tyu6fqyaU9hsJ4yd5OtEkvBlCbxF+S1v/khp78B3U
JtWMVNAalV55950PWhV7uLfLdMXn2dK1RaDFAYA6M8XqcV+FssflApqLa4i2
DXru72eEIepsf7/Op5eG0NZf5JGQYhx2fNo7vXnAmSptoeC69BvCzM8QrBLq
5ZWpks0fFtTMxMF9m6bQMIGrS91DZY6yuzdnXNbb2JsTd4c8TZ4NTs0Vqrlt
HIBWW1wEhEjmBgxpYtSus4eyH4j/I0wJVmF1oDehesOL+8yeosSRCuohDkat
3Y1NKWah/kOMy9uEsMWt8zyRVdJ0A1YVhFNcRPKc+dEKSJVdMgQT+W2Vum0o
qM4ptLHCpKKcBWgF3adXG1IeN/pVu2/hBu93ZO6tw1fb4aUBg3TYYtZj+/Y4
r1uRcUZvRoy9N5nC3wUM2JP4h5xKQfu0W5DK9Y4uo3eqXozXyP97Mt0MDFVI
qKKfZRcsRnsPivNzWhB0KOAUX1UFGm0Fl2VXcpr5QeddtBTYiyH/gUPI0d3q
mZ4lVkaL9gJXefRZb0YADJxhmI+CoNxft5XcJ4mu0n3Md3RmStLPQ756T4tk
EcA7u46aGSNxOc0l3tiBnbzqQI+/8X8y7x57TXp3hoSWMAF/RG3Egxf2ymcj
+OmY6N70Vkmmvz9d5rohcuXBa8IbANu0jMejjNZ5UpWUtxEF66th2cPbg8uM
cijlfj8LNvWcflip+xra35olse66CaR9ZaLM6dKDL7X7cL490OWju6kQ7A19
RXHKo8JvRrl7I3QrxEoH/tvAfvIOHbQYVkLBwypeFBtvjij9CZ7a/0MAB+s2
p2cPxPSSggKwTSymEk3gKiVk206wPLoqJqFa5777G2mF4FnY2KMttgoDvFCf
rU5cNOsG68z4pwyXLLZbugi3orNFWs+V7lK1XaHJSVPfwy9hiFe/2sFJXdkq
g+WzwGm3JDxB8TwOKmGFKNgPcn9HYDcNAZnRTXYsdI/UFkxNtA6B1+u+6Sg7
I/D+uf8uSO37YbfQ/Bapv5daCnpOlWMtVt2UD0j/3pPXmczYA3EjYDrcthmP
W6p7dnZE28aaj0UJXigVO46XGvD/i40vC9Nx6vhffxA+oS+HcSnM6ISlPhgI
QLstn9Z+dioHu3xLijMZeBqGVJvkBwnKOxl8sSoaKtof6Xj1JjnEnPHvlkwo
obixz4yfwi2fALYvZuFKDTI06GfBJqJc4Z/6lq74qljNy0H4OjgsNUSx8KJL
gultngMeB5+Ix7H8IcWgQEwd4Nb0FzOtcs+H+6VfyJhCDZ/48hSqe0TXA4HO
FryUjcloiwUA94trNEBmVe47ZmNdhYjHQyA533GDnC2okIx/IZ+2Rc4ymsAM
S9MhCB5an8MudLFeVVzoBaXNK/wCGz0gLe1d3KNt9XbdUVbKc6jaLE16Ka9v
K3JAd/PZ0OoBhfS11njJWyRyPSzJbySVQybgQgddWhJhihp94UfXmCIImcwP
nLU3koVSzSwUtRWn1R/VlU92MLt+h9Hy0+1/ZuyyUztfTt0mq3ybVaSYz0yN
CXBogiFZvkGjejRXHhvLOp2ocHRSquM5T1Kk/KpuQDEjd3UgL+oF1DGp/kTr
nE9MOdSGSDPkVqscr+RMfo5q2W9N61/A4ReQ2uUyWdJvbyH3QJyVy8aDQxBB
cNXGVElwnbICuX1x/JF64mGcrcXqktAs/R0ItC7eVy6yRowBg2OuPl9zJiFV
gSHFIcozhzTGuFZdN9OxonpHJIa6rHHItqziBElm+9wLcabZRhuReu/2Q2BV
i1jGRI3HZSBf7Zff9SY8DqOz0T5Bzes6bgW56bG/AGs4JDqvBIK6vIce4jBU
6eZ05toKUIuG+XYVRUtVLr2sRvHOcU9u03u4PuiezFImrOkyLhpgF0BL0S7M
XmVS43u42+G5mb+M8eS5UyyLegYkgswUHIEpDkM+5BWYqvxjX0+kdE2kwhtq
zeugGof1gNffYWb1kuJud4ZlJcJ+6i4qIcSJzZ5DDDUJD2MZIjN7ggX1DUKl
71BmDUGM4Qi26ed+nOsoR5XJRSPt96f0dNr/IWbrAhPaun7d6vEuZvnUfJIH
e5kRQtaJqlMu1F1WMYcVhC/sPAGSg5pm0rEcgD5n/KQFLWj2FXmE9FvfsyIz
eGIQW8Zh/N7qxYjVelUeS6R5/gOK6aWPkGcwhifwTtuxVz7mauO1A/F+W5jO
PEJluTofglXTXjkrrEgjrEh94LPBN1J1tODf2xZOiCcuGMATVwDHen57A+g0
tNhz0wxiJ0F0FIc61kTApBnTfa6C0mmEXd8gCCVvuWGCfXKY2bgA64ovDj1o
/WIHGK/rMDa+j4BfJSc/CGH/ivGjulzHGCVN+y4QwurPKJw8XSQjWzybRKgV
S3mUnoJmZnyWofaJ3sZR0eCdfeMGPBJq6Pegk2o08TOAYHckqGGbLChX3gUE
iUVQaJb/jSI7F/hrdTmgQELU5wjeSc/qkGxjDa6G99wBVu/OsHsnmfPgBdCo
8T6NnZngRUcDAJLJ9ZI992Kl8caHJZvtUO50dEqHhmzp7ym/GbPuF5X7IXwY
s0yiQU8VzlkboMy9HAV8zPUHeYFSHkSwD9j+7kBfqRmNbqU/9Ih9ub4IbumH
R7RyXadRt/e+Tj6n5pUIFX16dEEU6WJpA0gB86LarT9IxnEXVvm/SGSZDblr
vWm1nqOEI8Se0MjKoI8NhP19+IOts0PDmjhZDsv5v/37maeUim92mgFDPOav
NX00VDAq15GkSmcv+PTe1dHrEP0Ls5sxpnXWkwKG+5yFG4YwmTWrZOzkFd1J
1izp0+kHElb3foa2BjcxJWD5w7H4+jAEjqtlUCOQS/8JW+KFGEwjIMXgRnIo
EiTyTSisY5Bx5UO7zhBUo4XceyKNAYbDiK593Mh0/j7l3Wm8jHV2+rCidLzA
r4qoMMJFAWOdJT1Hbp5JhYKccLnw0SCDOql02VkCZUbRcx08B14ae9uLrABU
8dXVKSczL9PiDak9vsnb88UWEga9wEtqbwvwylBBer//3NousiCzrEyK/kWp
7f5an4MU/jcZRdImEQ25gvnHhlugxMD8E8dIHG6KrnscvuGjwz9zkNrDM0J2
HKEPclKZWEwqoYR+npBd/CvsT8Zl3hgQZ8Dw24/eL4rEjcnUm5N0Y+BVJZhU
o+nLg4bdWSqMMHmM3mmjKk2KGaO7c3wrkZ1a183CRuwhEpOXj0/qOWw9oIhh
yf3XU2psxSj4dy8Zc8A3W8NVAoglND7uyKPDrOortGg+Y2HjgVo7Ib5pVqq3
dhYQCKYxpBIawB3WvaaevHNV2PD/9Ig2GouReXE66OK2Pb5vcDW29ez/noKk
1TDQRNbIVAO/jZ+27g3EbpupcCA5y9EwFR0WCSvwWrCfABwC9+URQ3F5vfF8
glLuqjALqooP3SEagZtrVs8n1Yt4k9v6jMATVwrTLM4oka3oV8SidMS77/s3
748PyOfHyrcUQiFhEDwmZi9NzhKm3ODArONQnn1komcNOSR+1pSlAjuOFsAr
GXl70A/i7nH87i1SbyqiyjmyabuQC3mz5eWm/dRfolNWg+l4517+l2KX6joh
XjrasURT/4HsuvCQReGDN860qslyXctlAlxsAONgaQd0GF69CWHvv2aiTt6M
dRSTcPeVyCnzR8Dww6t5L2nfbnnqiKPBd9aKm8iYoZdK+nOXCXypSQWcegJ4
8MYKJHn8n+F0YonhUhaa/ybmxXFvS75dV1fFfRxK5bxM4EKuQLULrZ9PGMZG
RYjsZ2ZPNxe60AdAK7JNlvDg3wlHpfEuDq8ViU/v7OtJKG4FPMF36YARm7i/
T4+vaSsEtlYRiDnBuSLAfFpXbcvbPFE8CN3+CoKAshcrkn1lOz7QV2vrcC+z
xYDhe7Sg0RKz7juJL0SmyrfuXgKq1Q/YzieOXEuWqr5815w7Xy1mcyB1ylxE
m3kVFs4xBf1Ygmt8Z5pXAvOSBa7xp4Zk7F6C3IeDYbB7IhpCvMLJM4p86vyK
VhXpmKhDUX8FtsZpPeaxNCen8ItjsNegJjvtH5W/MO7sDlj0CNuskbaHu5QL
ueOSvWJ1/p1JOIWKZLTTFllR83wkbNPGZN19D8VFnyuvlPJTB1YDc56y+zkU
lKJP26GtltfcuvxzB99y6vLbRzskJUhZqnRjIWewEQCB4vHBUhHabC2Lv094
ccvfHVvC2CjQKZs+bU6+ByoHD7mdX8foo+mvrTZzgVN3UGIi/OkZUivnX5p4
+KGCjuZK9u6jqYw24eXvvUGGU30LpG72otXrDssE/G/CjgP2ok+s+JkuqIAV
GhH2nghtq+SDS6ralJMo7eF0/yysqe2bh37OubCDHLTSSuIOL+hYpAShH3XT
rLZj5PpxlpLjjkOvfCm8n27dak3cA8t6xiYxRAQVV1zxDukBbpIPOrjquReS
hUF8TUDAAu749XuImo+RJbsD2Bf2I50oYmwHze87vp2b8W7AAO5xpjr0UP6C
p4Rka0NJCmpO+A47LbPwjFtBsVvm3mDZ9+3bGtsVVUUJyGrg7pk9+bUlsJ+Z
zo6w3pDzSM2Q68+Egr04+vQYbsK6UBbVoqGC2Ea3qdGEiVzru7AtWEt8ztll
4V7IJj3PLlwwWOqO/mqyg8n20UiG9vX+zWpokZPdOufq9lCF85923zt8eO6L
Z6zbCBDxGfSkJf+spZxkWZzz12jWfLOiosXicSLhQq3kzjLAAlTbxhpAnbCM
mZI3XlUuR91R+2VVzbBE3xT1qILTQQgcOAUK+ueOZ6UpadFANmCTQ/tEkgiN
jhnaC2eIuMQ7ycdKj6GOlzUt3jfPqBkBszD7Gxm+C0h1NyxQ+sWlRcq4ONMz
5vWKTOlbK12hpBTFHSH18AR9Mo7cyXjntoK2Rq8S6rX0tzkfyu4MLzSDkE91
g2o90fBqPxW850GEUQUXAfMdRuiDyaXPW/3F1+cY2KKOiossY64uUXUdylB5
bjYrfxNG/42HrO6A5Ha9H4K4528H90OXk9R9XVnVxmtLDa4KucQNRqJhq3UO
tUYRAWm0RULBuE5q7irx4EolAIZDbemKmBXKA8CBmAIUuUnDoEeql42xyvkg
bgFV7LmWLnX0oU43j9He4khYCZC2Gk6nO3uhTuMwCvQrOKmmhUK7AYGcKZ+8
LdFwks4kMXCa7mb+BOlaTb0kiF26J8IRKl11mePyQwKL19GXW0SNU0wckt1i
RX8pF3qg/wpQijUB7JKvsJVgmBKxfJWjHn6D9pWBAE4vVnaaH5l3gdxFH8Lx
LevniTi4qpEKHfjskPllB3YBqlbQSWSP9e0fpQjjOgorLnnKOuN1mxVhbkVb
9za6YqOf73xZjcIA7VqwJo/kTOAp79SJ7xg9pVv5G8QVYbs+yTB09cCT3/+Y
8YBEdwNK5JvSgLv+P7Wiq6hTOK3DkjCZqrhWohKg5XJsWoHdoNGCkoq0up7w
+UPkRhkpkHbbavCk3gLc7GPHlF3oHqd5SqOifOWcYBdWJH6874LVzOkoaJ6h
naRpdwsEUAwc86sCpvPGWvluk7h9fCrYhcfFUJaH/5pepfvyCyyjtT/bGoun
4rspK3ismpzH4+uTADoa+mslXn5k8hyLZgEq3Z7B7k/zDrT+xqMFv+XSM3wF
p7i0sUaf7uO/tFB9py3TQ0hdwrNoI9UrT4Qon4Z8Mz76oTOu/n/rxBK5MJIa
+AQ1tVTD1XqQpgmSgx1SIJQBJKfZId4CRavGJwoAzS0Q8r0SqAadfsDtDFCs
lFm6aPK4wqWseAFupAzrdHcfYtHC+6PxUF5jNwd53907rsb7HEr2enExGQdH
v9EilDRrvM/QBvJ7eaxw1JHL6KZ49FJERficScb+7EEh/JkXPKgzN5LSmu0q
CxnI8TmoEv6SOu7S5WwdjbOCu4rMaErzAAnFpgdsN3Nf1HHM5ScgzANrOSDf
HTfMKvMBkdmiJy5mLNEfinCzv4ZZ9OktECWyxMdJXSh41kMuAFgh3NOYbduy
ThhQQvdLf/RtrVwsYL9CBpZyoKjsp2gq8wbowDQdI3GCJOqQ7Odp7EHrPW0u
gzgpqjVtgiNgJFMne/GimpmgIU8hezyJfyl1oiV/6PbqgUEorOZklsXSaoDZ
d7tiLxVyTVPwLYqZwQz6s48JzGaO6J7QNhedzeV1eIzSD0BRjSJPNQBeaw1s
IjhsVL1vPPhki1ohqEW/0IOsjWKeGVCWkM5+eVpY/1i9VFPlVoWMJyW97PWJ
AZowvP2i92JCTQEplwrR46BTItaOF3VjKwC++UVvAwMKicZe2hODAdYOwOnI
VTooAmY6t1psHPKj8fttrsAuyO/twus/zOgUKCUe/eCJpnJ1aNSqLwp3sswA
gIwlkJ1FfQilwQY6LWGGa0hegr8l1mPLfIexCJ787VQ0ON45BGVK/E4McfML
iZmWVAKO8DeSALICsiDLvXx5OESpfIaaDK2by/zh7+BNgHrgJzz8Rdn89S5T
SjnFelmiNIcyMhAdcUqYi0L/6W47EjuprgM4Y9USOvxVybsKQO2h9EMDIpUv
h4NJ1/bJKlDV+KHHMx3V4ZWpj1oOGvFVABnz9aWRAxBVk/AF9t9zGbRaTz38
cM9yfuhRXjyX2BujPWwAJx4E4b4gCkjhZrX5Z2TJjZS7c/2iG+m4l41g6EPo
kPdK+uXyiL0VjKwKAYyMsFA2sT5nZieYIl2YGXMqVI2UMV9xJ0f+Js/X/1Zf
whPXoe+toKBQs3KCq00F3F9Km1WnTUV+9FzzGkDhbOdg34u4RLYaa6w5A3Dn
f9vSxGFx9uLengFKSHLup2LUSFX0Uh6HaeeX9fR65zFErlUZB/4Cc+xDbgi7
+pLRKP/FY/yRFU2uLd7vxXAl3TTxaNIDl7LJh4TjYqwBGNoBsrHxR/FzyLvT
8z7XiB4pQXsFD14k8H0wIQnZ5x+7iEy+ad1yoEjTfXLooM4EGaA6wVVvrYFh
oCBF2wkft1M8kNLgTm4P5wKllo6vkqCtFA635oh+l0zagC2tF2UvVboYEmq/
hkmGSrRQfhhE/EhhhpU9tu3JLSfgsy3s5r8cMmlHZxe9y/4etNT1D/InitC6
xrw4DzpWLQdI87NkR4DyD67mxQOYJKJF3l1YVSAhPDs64DQMVhU8GXkXp2bu
2vv2aCOkCr/Mj+g+Kjfffv2j+1H4P5qO48/DNGiuYzfup1h0HusU6TDZe9PE
V+Lo9ok65MOT0d5JiIjzzmB06z3+4sig83ClnfkiDIz/iG/p1SXp3I++S3Wj
yxTV1nLzdcINc8V9tcdik6Rcf9O3Tij1dAjpkvxV75lYvusYUDuQCvhFVYoP
apo+lKy9Z+Rx4u1ov1B6Xg6LixWLw/zEfSMhp/1bREM4qQoOaedJ4IBgnkdQ
KYXFXa7Ithtsf2kZj56hRJlLBZXBvjC1Jd5sjnDWEgZSbPLrHk1IjwrsMcgc
Nkvb9r2cT8oWCpntZW6qA1IOQhmiiSsUH+Z5fYS2GiSpw6iPmmFtFgGtTx2K
i1SvOQzHFih2bjWDs2YiC3Uw7oCTPWhMadQNo+00Rnbuc2pl88fLHBeu1c23
F6HaxCO2JEXIKZSGfASUhauTm8kmBwJM1vVlQKMOnrFhHTIqHBCL7M3sRQJ+
mzjch7i9No0mJ64b+XDgsoMYjn6j/iUaSoePa2ILRrL2oV0GVxschlHjX9+A
8V+b0sB36qsa151G5LCfFF5SF5EHfaizh66D3o7g0+/M2IzrxYJHm6R2jRh6
cNM1Pb6vHwIolcZhINuHbtW2dg+6GVUhASC2XEaHCu82tAcTX1BwMOH7DFoV
ZHh+4MTYH94nHV/4IDtXeXoW4XIZxPiF5F0+4opbB4dJND4fsSPc2XIYfT0T
Et5jqkPllXrbAk5d3P5+7GhV2gzOk1oDdQWusJjeD2gphqLWb5kDWzkldSWQ
7Y3kIRG23stq/kQCw5dl5fG86MF4p6y374Cg83QRsWzwmz1dGmX2sZLFAU6l
+Hw3CT2kp6EidhfJ+y0DSjX8zwUczBJSA9ZyuecRpufG5gPtnacO7GDzN29B
j77VaKiUZie5B/byb3fo++qqRbemqb4PzkJFHTFLmjScf1P71hGzm1jspAVv
aWKA5VwIriurgfcg4vqwy2rGiIWoHgu2tfx4O+z0VNtptqH+cvE7yInhjbSq
ALbkGwocFDbJzUprCR4XE2Zr73mDf/gFfnlHxcAa2rpLzUlfAvYAiXwnj05i
+0UpFVDBMpR6G97Q+xGE748Mj5FSv8ErF4trts5+CAA4M31TlIRA/NBIgDaz
8lO40xzWaK93keNyE8vdFhC86TjX/7ASWZTwfS0KgxikKuJW3o3S7fnELhJw
MjGTzf/lWCiJ5kgATWQZgShl6bCjgjfrX+BCRhjJV13B95TnHLsrWtvFBMDP
9/2J40xtlMGhcP+3n+idZ+k2fcjM46+nWoimQKbaGG3cVyJI0N/WTiWBIFQ5
N/QY7gKs/s03i9PnMchNnsGrIriThxIBYvV0+Qw0ER6Ctuv2hrjCPKP/rOMO
fentng80DgEir3OIKBWvBnIqA7IrmiybQ95k6b3fghFVSCTnYLj6skintGdE
4ww1hzvp4MUuG6pDZsmlgI3V3zzRc5yv9/WhxpOaFNpVs4vIi8SpiIRAx+Yw
CsPJ+AEZeNXuFvaNOPZzp9Apct5lC+I4n1A511zbKk7a99k0S7KW4RaSKkV3
iTlQAa0f1S33gg+Sz2ZnLq/XK92KcxVWz2ngrEFJDL507C1jR0Gk7yDBWqnS
zhh+yexA/yLGLAddgFHf3Qr+tiUp4rg7N2W0fTddBSS1DNAq2f9kTEgbLDkh
pJnnfmt3bNfmZctkqnryCrF11FZHxx6k1jS93uBT/PuGphiRF6P1jl5qCyN1
lCtWhC2JLIkMEAWgF9BNdg3K9KfHAEKn5a5zFEF4ODw95r5IOzmIVZIftho1
fWaUFS6czgTW2ClD+rwF9bLWPGXg0LJI491NvNixPxi1Gq85+lpn3/sPsllR
57Lx1PC6g5Xf8CTm0WZY+WHk9vpog8+ueIxM+PpuK8AeE1hV6apHvN9uKc14
MSElbNPPhTCom02eZx88AQRLuIWJQR8UyVUhv+3mbSeJL/rTW1yX1lP+pm9d
WX7h+z1sdg0FPv/GgT9EE5Az1BkFoHP0/SHmeXSs3AJyhIGV7bkkY6xxDwSl
z4E81/1bK0Uk/XBUU/n0H6Fiu1WxMATPr8CCA82ba5d3qONjzf3Ah4Dfgr/C
0JQGcgoGuH2DesqE2++Zgygq1uW3gWA/WObc4Oi17LPZnYFDYqsIsRFhLnif
ub2SSyH830iFbsgYs6hNqZqGd2SoW7MBers+/qTS6MEj1l2FpZp2H3MRc15V
ZxMjQlpPDCz5UeA2OmuVrckHeERzXaVA0UYSlrEktkIPjttWKgib46OMsw+C
E+C76ctyWNRUuUpIwbcrnLZQrbBcyaQqtxKgR96/ZnwB5fjkzIUTz0l0EjE6
w3ESJb2+q6sAVV0nTbe9e+R2L2d3QSDEOpORLKhbJmGgcsWX+IGtAxI42GyB
aqAWJxHU8RC5tu9a2LdXLhajeT9r8zXTB0v0vx+tGkJOW8ssIOlh856tz+lW
b1g4d6g5LYrjJ/xgvd4+N2RnGLL0vlKiDf5I5oL/EDMEs+YWMXja1veXo+s5
lRt9NMwjVDeDv74U9fS/ldB82SlDu7M/Y33frndqlmYlABCamZhkY4W9TG1Y
YnL4mnpqKgdoJxu4spYEG6asOm2jmJ2fnJbprWGu56GLpkqzgv4La2PeX/nz
v01S6WCvAgu4Rz1X5oyVM2mowgF4mm1Mmp2AiE5OcWsWGW9t/GMh59nFYUf5
nwXhpjKXC5k+4FTr2aExh6IOH2NjxgUhWSAAxz0kzdxAg7EUjBRbZLE/daUh
sPmrP1wiJ+9MGFRKSDnnQLrLj/GA3/O4tC65V88TtlKZDfdR0NboPa/AGbz2
m/ULjso6NTw8Lt75CEZrj/1yvDKaAKT1OZK8fyrqljATmxRXDznSWgAEshuG
N8HTNLtzuiX0kOGSW4WDKoZBEu7aRwutj2BF9FXe3mw6kM4c5V51SaqkGp2M
sntMbg7AUbC4s52mIKpJ3Gu3P5dKWwnk3vdP9KnRPOoC5SdS/crDWks+LxRQ
qHLtCSOPRZ4FF7SYGboXFosuHruRyBeOl1FOt+AI7giOTlmth0Z2pPuKmtFE
murneCAQVefrVKhw8MycqgeLulriQiDCZpwp6wvtHiJvmQL0PRKEmicMbED9
imvQww8RRwroc+1MEhwbX/+Qv1YYD8KIJcSsH480+3RO8j/XT7vnxRbGIeU1
C0j8cY8MY93HYzf6VGDzyrldCdvYCjnVfDZCjQT91fJU3okBX0j05JKYQE4P
dn21y1MrWefIWix/sVf780Dw9e/Y9yfei9Rp9fYJLvr1LeNNwimWXuWqoIG3
3Gw1BqXMQ6MjMDmLMtnee5fJWR4IErLRCNCnSheH1Nsl9izp/vFBQQjazQsy
2lVJyurAA73OuyBiC5kc/L6yGHsPFjfS9Io4qBsQInEKAcNNMRmQhJXyXq6s
DGRfal0UL4cFrym7MuxMrlLJ9CMLpI9K3ygfgjyqfsbpvL7gonktlaq1kA7T
DZd+3doo4rlW4XTo9al3ouMOH9NbeMQqhnb0MjSUvLvwNMDc4OgUaTo/TSNF
cGIGlvzPohOzGveGTtYBZARRObM1t06FEtBCp/hbmzQ8v8LW84+53rRZViEc
cHa3nKfk9gGd1hPyDel5jcp+4m4J3iUUXFwfSPwhzle5krCBGhjedAjuOswO
2kzR++j165f10JpM2m5lPXk5Xfbg/u8j0VgWdurLrU99OvPOzf2URjrU/D61
Zx67IujhfKp8Kb4+HOHZP40cYHQ6sMlPjGDvP2vho8S4gZ/VWAZpmnBVSB0x
VFDOmKgQzm4fOy4y/62ZJU9GJXeqJ7vcfEB26NAPYC/jip3ZGF1Z55VMpuqk
nlaTHuoNlC1KtOvVwLE3/nMSTu6gyz1xC6LtvU/eesl7JALhmU5lq93ZFl8c
XStW9EOwRGjDq1ZhRSbG0sGJXXPgcb3cgPlH2HV/BFcgKNOugUQVYgS1YZVx
gvwCInISZm++sgezT0wWaLOjbucDOdsk1GjEk+WP/lMOoBh0nqCi956m5PNE
0rdx00386OXthaHIM2zM3Q69n+6nBUjS+S2ftwLkNIsJdSBga4qJwVvl4peo
CCIBt2SlJ7mZqLy/wKNyIJEvF1lzEs81RwoxgfInPVpRwxwde9EaH9iQIObT
nPT89rPS7+W8EifluL/70apKMhcmyeaA4OdzIEq7GcG+H/XMh8K95bZyYx9B
jTo0ezGLs588gqtPoMmmRZokZmv93TaBQc6hD4BPsQXG83LFH6fw//M2phb2
cfpSAafBqP0jBBhz7LNbK82T69EwdDrIDj3T3LPdYRy3ZNohzStblZG/hQFW
fnFWSI6I6Do15yvFFyUsGtaTIfPf6S1BtB1KGfQjCIHFWrsxYLCIx1S9OtYC
JzbLPWdaq1qg5H29MC7h8BHLAEh/9psxwK46NDtMQJvt8qaf3QYlrdBU0Zup
xwseZNmAWo2B3Au6MuIGQI326wOrccz9M5RY+J5iCQlHA+ru/M9OVqRqcUsy
V1UmAw5bt14C/Jd5UOD1hFc6DmLHkIj6WF/GhPP+qdqOJXgOmhYDwsKnkwel
HzKeWJqWL7dDaNURODJ69KbBuHM1XmvvNDePmoky4KrSQI8IFkMfrw4pmI7W
FqcDzER8u2ks+4vRg4rnO4deLKri4dzaSXebvxMX7/5ku2ItpiE+TuzrBpFr
IWaxbQA819zpTTSFm3D0t9rEWRiK46fi9GWrEHaenGYm+KPzB1CEaEXYXgMl
ijF06Fakh2V/y/RLAv/gg+lTXpJvr3MEQRf7Us5vea2Q36ch38Qif2/hbicQ
FYoZOxrXz4xKyNlwMxI2MtyWj77AG/E/FazL7soX3OjXHfVxj6yveSOZ4+qi
2whLauYk8LDlJXeZv5ngHWHcAMdB7FcLAx8Ouzse0VlK04lVboT4fOcSLhnm
LzT0Vb3T3YHrYRNq0V/TUr65YIZtPagM/+nRBDTD32yst25LUEW7/HhSC41n
SRCj5x+PSO533MIqLuJ615JlsRBvuNtp1gik1hi1fM0fjk0gWlLHiMMJwimW
X8G7U3ddk9n3jETnG1y6ckfmzJrlDaTsMy7Oj8BOVfrMG8ljrWNRTYAVEVhj
L2Hlnb851izDB3Ambqacdn4/I2snUZD1F5Mkz1Lzbgx+QoxX8FMcPl27S4fR
srEDAV1H4cim+2si8KS4W20wCsDrouIiNg0hPKwEIXspn8xAmtN7eT7/GDJf
Ri2AFxIiNMBCuMTPhwKigQMSByecMNVBq9aGj0xPKgAzI59pu+WRkh1SFPkE
xvTIvRDx1GxfJqHtg0l4sRSOKxTY3KkTEXIo2l9ftyR2d2mHtufjHlkaW5B8
GaJhS6C5SD4J/hVL7tQe9fMJwUDcrZ9w9Us4kE20RCcPFVgG/qW6LxpBGguA
eVSmPjNl6WIc+2zv7avr5mEyeAt+19W0GmblVBiOUwDJ6bdnkknIk7OJIRqN
Jfi3t35quCLThJMO9zUDW9PLNOVkO8sLAyk9G7cdMAg55Oyas7B+Zy53iogt
VOo3EnzJk3fQ0/NKQuzn5oi2igoF87f6O0MnHkAuiCVeE12NUUDL/QCXX9yz
zoGYJxDxtHScOmjC4HfQcSQGIebqo6RRKcYsHKcrCcooNiFgVuB93e3cf27z
dnAB8oYsYC2gqmMWef4xnvJAOHKozZxtFdtUUp9q6/yJl2UtzaTmxYa4ha5N
ODz9dqcpe4tH2ESGEGe27022AijD6BU3zBLL3vFlZ2ifa2rgc0tTM99Og0Xl
4/stqc7G0Kj6uR+Y+vmLSPssFuCBH81+psI50gwfCFR+mIFZyBzTsINpbs5K
Z4zDC2CAAyqNQyN8IrD6ne8KuAt9tMlXfId7T6aLT/GSgmOHvnb4DscSL96Q
99zt4qAZVguaHODgK7Mlbrd7NE7TW5CFYCa/EYgV9X7sH2io1EQOvlEpBZL6
UCUOmX93QmTrSBkQT/fEWOlMJq9VjvM8sKmiVGF40t06oE4qTjSb8Mv4vvbr
tXeoDZVNDgBiaPZROF7+cFV1O+rrJNpqUAt4PpoTpQhVsIuRmJyIG3Liqm3J
8iEd2AHdOM2tKE1GYSj1hlM9ak07O9cFJgz0vFE6QWmIuylAUqsRmXK0DQMK
Yw+sl+y2/XNmRGLgMltb2C+zSpiFOT8n6kF/GI9SRZ+arNS9RZzcdc7UccBj
xp5L9jQgylgIWF21itG9enZN8czKcFrNzn05AgLOrMngJ6uX24Mw6bf0pzJQ
XHYutpaAy7sbNQsIvyowWNfNlqjdOgBluoTDf2t5fKlTR/P7pfdXfO6CbsX3
AJgYqmsAUsN0FGWxJpC88IK9sHI5D1vGp1kJ8xFqeq/Dc43ORb/Uok0K+vhw
aC1d6hyv9x2smEWB9qCkwfpwzRm8KntsVIUzx9Ikobq+E3QuXWzCKJqCq5M2
BGqq0+5NzvVC/+a0md/ZUe7qVknuXR9pCHvf4Pl8U1RyAGfcTL+hS03qnbNw
NlOLovT1dNLdtr6wjgswal/KJ8k6x4YoasAklm8aqZ0+4L9LHIANvY32NZ2m
Iitpol0rIzaZ0n6xcyHMRhZrjIy/8RCm0kgWeAvsjOOjf5C4nNRYtUH/lA/V
xVIrev/dFVTOmS2NPaXy5/PkbW8Q3BR3PYEJWaIZaE1t80C4NzhGi9oO7dT0
31EN08/AmGAV218XuEyoj4hqRt/6qf4umVysKRkGjAQJk0DIIOvzZb38PY+g
+A8p2Vbwpdr8YfjJN2nC9c7HV+3GX6lxqv7PWwSSbpXI2alu1sf9fzlmxJrK
ALpA++obGUSpiAAp5+P7win59DJA1N18Ub9a9w/Q/29LdWGguJkviTEMKtYO
bCHPMneD9ceNkSzioppm333irlaVS51sEwYjQYSK/oWo2QrD+rLuEYpaaC2Z
Ki36IWRjWsiS6CsrkVNV1iynu3wzDir1lZi3FDv/W7IycN4ruC214MZJvJcb
8wrv0QmZ5jxXtbvMAE2flW/5XjjBqwJu2geT9fDNlZOsWd5C9tPt9U7gGolg
7EymfIoHbx7DHmcPUjeHqmlwURCWDSlYi7aF0g36fEg14KZTXOdqXRQYwldN
+HTLxR9Iz/DoTdITO/trVmsJ4EuWJfeUU8Xt5rrdHpM6naBTsydGbAtmebRP
VoE1zmm3N3Dsp4VP8Jn1EC8xG4XkVYkJiJiygRecqBCnGNUG1qHlVUqCMkcq
0wjE8y9pTqvInACa5xJLnegqxqppT6baAQXx667C0GOtnbRQ6CivIXnyJrxV
m7xbRG2o5oaiRh9X9X3yJ3hsIEi1QVXcg4WzJEbsCbqhAw+gLJqvfKx1Z34H
ONNt1lYiYK9PSUaVikqBEsklVp3ApAuHWHyCFsEtWZcZXjk70YHuYeaEouC7
VWe60ZUuAHcttcKg2ZpRQvLBjp0dXJHNnUt+31H3oiSeBcOoj75Ooc68mFl+
sc5P3PDmnal2Pakjd8kFqeA0lFD4vg/Noge3bzKY6yqBf3FKVzuIfkzBCQjW
aUQNUlwSNiSVFELEkphpEVjQ/MLNMm4IADjapr6Mr83soyobFyZc5rvSCbDU
PXwYE+gTNXUWf/7obCklsggjR1TIyZq87KvZupvFWg2+HXgKnWjfoQhzCMJp
Vaqf8Q85iFWP6fpNKdDIJlPNwYk3XHb490Kb2iFE8rO0EB9hqzw6+TdMsYJO
jBcWC/u5fBGCUAiXvbsuLLkyKAResvU/w56fXiQ75IVv5dubsXfm1V87Uksy
tIMRomECOj7vPBt2TDraX3VVf0UM7ChaYy0ktTbD72OtIjbxhggnoZ5xrwiM
B28TeKpYL9QA3rX4wtltOMThdqlGsuBQPds3ND81Teax7FkyqV0C2tBZ+K/T
e4+Z6Vo12Eg6BZPWUHbAakeneOUnjaW5P4O255J5SEookHpmOkP76NdCdTZF
0/uNgQCOrni1qnajDgXri9R7qn2P52pc3TDv1URP+VD87tO1ChLrnr5l6ZVh
Xyv7PAOXKXKCNwD91J6eASWcIkPdxqgCnJr1yU+6zyKudgErzdYSVG2NR0p9
DJIropGJQInOFjjTlcc5w9IBnZUwqvTNFHDLJtV10Jk0SBx4D1zrXayZ1AfH
LrFLtY/sbvz8z6WKf7eAy/j4qoqf5hZR6sx3+j2uhchkG2MXu+JO8Znopmc3
fdCN0LshNRJhK6/zB7GeABHz3WMkgFlwP/mq9X8MnutS54sKwVimLx0mZLJK
mqNceL1Jnz2Ig0h6F4o1kwE80XuEcCrfcffcN7bRBihCFdi1Mmi9CzC6sbIh
nwiW3u/6IiA8z1T3G60bRTysqCYV44nPjw73C8lNqHekcuvySCbFwXOJvXaS
wqsbYnNnEr90i6xgQsdl9XhFifhHFa0PDEgZ7wXwB/8OGQWgrjkQpOcpagdX
+Nn59aZgsn4DtHGmQ1oh5A6rUYwtVftoIKooRBd+VCI0WGwY5rajpkWOrsEs
Eo+8JiIhJYI4HHkKBknubghqwOsPmB+KFAgfAsILtldhSghLb82R/gMfXufz
tXx5YSXPCYw10NLr6e9xYMuk6rgCtGc1cv5RGbKN+JHvHLt/PAKsHVChxODr
IuzZodpHjAaXV0yF8cEQhRmr+bxMJXbUpmDOOeJv23k9qP5Vv6MZ88BUMh4i
qjXYffnBDLQK89xqYR4L3tIrIHh0TwupxocOOEaO0heMwsLOX8VMcVm7/ar2
vSTyHzx57beCF3DyELN+Jjat/fx+t02vHiwPhT61OUOR6ihkGQHUpRYDuSiM
dxaFqXWGsu5c7yMygfpNFqs3UdqKeKvmzT46pO37+xZfXJkmmfE+Jduuc6Qk
Yejx3eV39LAgGAxIO2kyTLbx8V/kMQRy86o9ReJ2BigMw+FHAzf7UVkKgyCs
yJaLfNJzX4X0+DLWiEavA+XcZESGT++IZ6br5nlxbiD3r52DJErTxkc5Bddi
J6gixVeHS/nYCqr4M9LA9wVr0G6qajj2841zJkhLKWy05KF++oUSqMkXTUe2
7kfMkRYjhM1pOWJugAS1MlnqRnv0x8Gy736HLXqyisdjJVyEWUu3gAgmUOTR
etI8mdI5xBx3GH80CDFBUzpvtnEtHvLvCfBoWeBkZ8Fv/OrTkpyIR3bPzUCJ
UlAvyhstmp1somVF6VHLJ8pxJUUGDK6e5uo4FGg0KeiFEXMiMM/WfE/2/Q/S
duia3eLvI0QohLYFKn4e4X/s7/rnYJmkWyZOEJgjirA2j6WT+bj4+NDf7WJ8
e7bEVbhmPdB8yJa5anuY2xszrgijrfuN9UCUQLCD08Z5IL2jPngeQqg56hT8
Tojs7SQO+ZoGut+CWXsRzrySE6HhKV3bsB/rqEhi3CG2e4piqk1dHWeBVd1J
Pn5BAGG49sRDy4RhCxtri4aPr2FxyuM8OzFGky7f17huYbd7amXSp+b2+V9K
1UR5KAW7I6ow5r+GVnFNvnEE3OMIAqA4n6vqEla7/5bqVYsi8brAO1570734
EpE/QnO1izrahlGWVv12lPR9dFA3uAcHgtJhFU68YpyEtP0b/+hsCFWuiuPF
t/GY0NK9jn7ePQat31oDX+pCryLqXxrOMbyw/iq7lyJI5hwW09B0ELxLkCwe
5407d1oabzz92cJal/yLMIdvfikS2wTlCT5Ww/ZLefCoDf1fooFbVykG7bF1
Ka4rabw5d/grSumg9CU4rLEYLSz+lN4auwGfuzU26LzkIo7/H+OnZnvfL6CI
6VcHGcY9epV6ICpyz9WTONCA/DzU8whUpuj9fBf0F33BeBI6R1ImJjDfJgzX
z4OPVV9PxZX8GLnxrNKOUPh62P+va/szFdCCqY4yKQl2/o/oZ7LBGBr039bA
+cq+/hELGPI/5GHLFUQbRNvNPVsprvJa+kXLgN4riXnIHK323Xi3LiVQTNHE
BNE7ovwgz7ek+adYAcLGThjIJgRZenavN6JUPNLy1AZKKyOb71GfAXJm1HeA
SoBO2loA+NnSLbved8uwuXVWYuIfpYfKq4tN5zvGXJD1P+WMiOJUnCu1YS99
1mipBLSCi5fgpxR8WHHXbacfptu4Nd4xhT3SP+wVDKPJLmPXsYFYuBmfxmeY
TyrSlvXElws7mlTZFXtOgjCnaSeHg2yIr1Sh6aN01LozV1Dz1JESMvJXBvJY
xcPRc2jvIoM2p2USxvkKeIXMfEOQRktIJYplKjAm3P6jh5j2fTrn73lXQLF/
N5CRInLl7DcG2OXvLpf7oH/Ki13Z/+v7qw35ALOq3jCLjL/hK8aflJcR0wWA
Thrn5zcgotSE1ih+X03QNzcGA/bzZOM8H9SOPW9Dms96xdrv/uKH9F6cJqGH
cGfgl4RLJ7wCI+07jiIKGVNTdXYELnWx25+kWXlddDIY5JhtQWKWDlS+LBS8
yAndVLegMwrOWUKFBlQdZVTAiHQbbzsRISXK0JeQwUxaZYVYzrqQZ/C5gnlY
3NNqLPF+yLKuysWk1kTCGoeHdwMxAnSfqfLhtDpZCnvrahQT8S1GycUJYZvz
ZBqi6zKqwiWKtHBR75Ny5cTcyRap7yaZ7D2nF8MwNiC4pOG9MclEPG9aXbMh
Bfe3SWahPqkCF08KTzwMxV3nuRuwL2MEYgvwWmdyGab0fuIpl6IgxqxivTwE
I47eH738mkvbOM3+K5mEvkfVgNge6yJLa/wzd5K0ucrlY4SQLPxlq/B1HTXJ
REOGYYRlK/IPvy57lynjEj26edSLb7o7fQKttRZzNkpEm1I/u6fPaU0mmnqE
0+fDtCyOAqn70yCstT7xVsKf3A94enini3SXSgt+ZHeXBi+2PBnNx45tHraX
1dVKVfxB1v/WBYlvAwhPP5CgccRpAgatpalsgA5dUmQy0iZUQh2Fd8k/gte7
v4fU0G/n4+ByBaw0ESJEh2fwUdhAzoJiaXXb53PQAFdejSdUIlatgf+lFH0t
AB2HK1I/j2oekOVkHHTrvLUDCSNxME2NGn0XjtFGjeOd1KXJCXx4ePSux92C
BR4VPg7tztKlJPEOwwHNojYEMj9NWeKPr1KV4YU8HM+Pi5Hyn3bUqdTJNDwx
NzDl/XETL06RgtQXrnPB9HeLbvkvlqP4M2jiRMGrVmyA4NYmajGnRJhrwZHL
rllrgX3WrB2i5rLu8e9MHvzZ5zS0VFkbC58qp+RY9VGfAEMvcmEKXYh8MpvQ
OxgGs8oMdDTgDV+vxQonJZ7t63dVFch036+gXsQlFVq6TC2ozkaWdfRnZPum
3cohA7CT73jORIn59QU2HDW/BXrr0AusXIGiDVtY9tYKDTpBSCQOlp+zQepu
oWuSqKWvcpJQkB8aDXyOedBd7Lo+qJiXcEVuVZTUx9VtIuvdCHQOMKfjao9O
DlL9cqIwI5xNoCcIFvTaYNik6+Uv/nCJ8/OWdYoKvC4nSJHDcntS72kE58eo
w3NCUpXDuBxWtNVzZaieD45es0EDN89XMYuaEWt4TMO4FbVQlRlMXGQwgzye
WaxH0jlVRm/voCJTVFVqkHSFt/WeL5QGOMLM21HovPuA9m00OTP7VjY4Hecq
fk1wMqzO31qZt5MylQtv7lbBf/4KGu+LkFTYQ6DHIiC+2d9IA69r9aHQXpZf
ZF0wZ8ZQpiph7V+VVGV8QcBu4Lehr+M/0a1IoNjaM0G2go2YuBTPqG77cEMO
81N6yN+EURlGKHCiPhDozIjri8HWDf9nCFmDXd/rr8Mab0gYPFr/lOGNsPR6
insJZY658bwFjoUiDL5nymYQ+upcOJ9XNTTRA4QwW1D9NZPzPvlsIvHDDUSo
erAeUQtou1yniFMn2BZZJSuv6wGJezgACLY/0gyKoutmYRBx1/b5GgJtYvJ0
YuEybluoCoVNiqWCNDcovC4irqq8bXnfRmTxCS9T1mPXxboWQv4NkhmrKyO2
jCTeGNc2kbiK0idpW6OCSBAkgota86AJuV1wwPq2IZv7BBM7K7yk8Oc9iZ6+
TO8CAGk0sz1aA6YCY4cSXw/Xtfl/D6GuA3r4LsuQTVXnqlBDLEpylfmJr9Gh
l4iZ36kYdLT5dRtZXWUttiCrGT3OjbBnWDOtyiZo+BpnYR/t6DN/rh+a1zrq
8e2cTFBVyWehb07oo2BgkxUW0XBM9s0EqSbrWUID8nddD+nVc1FL74JZ+rOh
cggFInwfrFyV+wvJP+uuhH4CGJc7O7XmClMfaj8ewDlFOZPyzZK8ThEqDlZ8
gR9BGN3MEAoLYs2Xp2KFDsL8tAcIk3zx6Yjg4ES/encid4Vc0oBMP5R7rQZq
BixbRcT1cYnflyOM4X0pY4ByZK1mqy4Ek7m8C7i/LNdc0gBWyJsYUf3IkxSx
Z+PNf2YUVIT8LLDZGcOjGsUVSPSkEhO6nADXbRXEgf4AYDCxLhQgVF1uqn//
GDogtOgycYWu9YLLIBj+qg5emoxJZ1AxEFgRI4XBi1MZMrnB6gZT6SW5ERIg
kufuFBCxBL0ccCc395ks9r/BGstMQtB3zF8eqs49Yy/0yM6UdWWlgYXh9cZV
3zPXREE8ZPrbPz34HChWgR5jCpDD5terkiiF12wGZ/mdJOH8SjmHeGMSCxkK
KGIqlAO9Znd2CnoGmNKZyIiR9s2jL33gRnAEM13sKY3Sd/tLUalk5j8DFyzV
KXInZmyxb4e51HpG7MphyuwaTRxrRAZ8mEB/PM6Api2Q66Qb/TO35vaAjx05
SCkOhYZCD7tXuRzmVnZ3LjnBaptvGWR66EPkBNxTPvSpwu5onDdw06IVT+Gv
GdjhnEndfgYxadhG+A1SzHF/RhVTuvaSJgHO6VdmpGPfBKvmyHetZnNvr0HF
cmgyied0DvyRiRS59KuuwII9yQhZMCC0OQhDuBwqvppYgIJcZSN5uRutoZsn
mx5UJ5+HH/LxNPoIOYS8hO02yhfIA4FhV0wBJ2nOHrycTL9RevGn5ez3EGUV
k3PS8COaPv20OTwqWS/6GtJrNVPCHWk7UbWwmBMbAGJhlAa3u5ipsUJ7nDOO
zjDCANseti4Q2LiSfgcbYwiBiO+BSz5UPpM30lvu4JQvBTeeaFZ3KKFsXThY
CcaBBuz2Rb/HY2Xt1k02dco9+bu1JBhB9I8Jd79ad0Z+zK1pYJka+PXOL8ET
M3d6UHihc0z+di5LtEJb9drzTEBwoOfpRwBkBB69P+TxdeAxkF2eH5rq/BuD
+1SxWuGn/LdMzn+FnAMIvrSCHP6AMU2UhzIb+09KP4/BZ8dr+napKxSOqgAV
DjpTr6cEkgwuz1NIOYP73KNJ/vk16DcqYl0Og4XalX20OAAtnoMxXYPCKu1j
Uwho/Ly9eFEHCsD3KoQOM34Kjcpf+CoC1lcGVHW9q/nsNWEVdhRDSWVd2xpU
OQ5/g7pGafqZT2/T5Cz9jrCwt5tbAkd22v2KkvypqYnbccgWJU0jVYRGXreI
pEZcQlh9HcyeUN6wGB8ocpKXFCXgdgG4gkleuh0+mdih8CkKzNu2FPj/TFdu
BIPWl2xnnqasVSjCESPkCu5W843Qj07GiQeybMzhgxwERP9JHRm8A6lF2RwW
Csar6vGg+meepZruYRLPhJcr9daSHahNAr+4zgu0paZjfuheE84q0H0QJEGT
kiSeMFuFVEKJ3xmkfCbhobgxUm8K62txTT24jrHfjm5vLk6FHB8hABB/AKgo
bsQ9Uq8UDPmtnzovVdVY7057lMH9Egy2SLGVS+tENBhnMH7wZjQ2rbK8NgeR
ocPUmQBoltW1m50yTll/62LPOXzszBavxn8EyoYCcWM+yV750CRmTvBagHMs
y88rwy1bh32fII+2v8UJdzTv+rIQXKSAY4CkgQdm1djcn0RZNPozZlLKgDkw
IKOrE54BhDGry7mcHkYq87wkTcz33gs9xaoa/a7DWD+zIVKU+1SqZhspW/5n
w5V7s6UTmbFppPjQm6Wu+V9ZEbnnKHKgoTMZQFHTy7w7Ccjl/dZTlAth+c4D
KfKbit7CsqLKY5LglRatEuWS8Nn7GVhenlx42/FJJR700gaCII0reFnJ7Ib5
Tuwmj49OpHhfcuqcuxTRu5M13WbxtHrhwlsRtWoGLR5AJcbD2nJvBNoKljrA
Rhk+yumng0d2UmVg8gsDI/cuRj/LgIuTiuGC+Q49gMHehg+iqhgDaFqkvbVp
5cgIOAjZ59QqMN+4yCGSOxKnNZehlu5j1CIIEoXX04/J5CUBDiLYvMFvKOv9
UR/faG/T5OIIYNe9vND06Nk/cAP+7D0rRKS1Q7n7JjBHAiE2kBj2gh3HCsEw
takicbQ+Q/Gp+zJwKqLBtm8IAeaWV6fsWmXVzUTFFCvzUE4dIot7pxlXMDRh
gcBJ/aZ4Y1iFBQjxi+08DmHQeoISJXfDucuYJUPCj5tQqRFkr/Y4uUIf4VQ5
YVwTcHlGqlkGonNmcvOPtMtmKx+2E5R/s0daCRLKDRKotqGeqMD1FyFMRybO
8lIYD1YCRk7hgZEA2KZAgm+uip8P/xng4GKz6w2yqW+gvn7psf32LUdsRgsW
ix+AEjYJct+NXW96kJYqZsPNvkcvHkf6nBSZdqslH2XTBGKZv0Q3lSlhFNrb
eHVPi7VuOn0TLfehGqnmBlb27ZhTFD5MWJ5DGITh4G0ctGVGyqcyOrqZFPSz
8QSffaIn1yixWgWBfWjF6HBVGplKN9nJSQDjbNIo3HrVr1vLeKMPUu8K3ZZz
dP7hSN9dRfOGi5VaDFD04mVJV/6gU4X+ti4cbTUTOVYLQmqc7bXQlJxy9fl2
NJwzNMsUC5GaUeVZLL+7oKqNoQFXFOdElTmxXV63+/G1K9vpnq3McL/pOORz
R4Q5upq5HbXWd1SDVAfXCGZZsrKPxvQi2Yaxs6b5WAxesYouCPsEZOl/abF6
wbYo0e3lw2X3cOcbrqTkpyktzTjNb9SdiTY6ohbzAbf7DvHiWoboLip92JiF
o9EohJ3grh4sbCrDyzSi3wFD8/W7JSYd3Xdu8l5LZ/fZGT1bYFXunfcUyWrW
Fq6YD0k5kWoYVyzFkp87NhClFaIbSDImCUYAgSf9i3E/+BkNLGEkaYd+1MjN
MyQItoxwpHMUCDvnan3ngZQTI85Fpu1+zEt+wrB3b7CzBgxkLLj8oYLeNXmx
1pzghIKW58hFUXMIHLauaXbmgF2AVU3Gr34klOv6WA4zjFurMf7G0JBLcN5O
RMVQocTrzYtVSFxLXKjQ5m/i6ZdtW7Xq8AHasFoA+oJ4bbndNdjYYadz1yGv
24Zcx7gA7JzZdK0Shrw8nKI0KPO6g8HW2rOiYx3j+lLkKY/rCgFwTPyNxhOp
PLuxk3oOnE2nu2OINP4oXJmk8zKxWAPkPeTYb/OHeVu13X04mSBdIY9VueBn
ZP6wdSVIFLh91Q37bGztHqjzxPfvS6/Se/KdLmos9JAb1jHLJEHDN37dFftH
XFOy2dOSE6w/8qUgPGtUA7UxrqcA4SC1ImDCiAhZOUMztAu7RlMQDtw8PNgG
8Q+Isy9EyPIuJoOj3WpprzGS/4GFmKY1zq4x+2EsRG1mgWKN+X/o7f7qKq2A
XazNoFuzsKRznNC22ycizyNd7fnb49uzaRM+zXmcCGDdjOCT2rJyf3UM+Sz5
v62SZjltIUEv4+0ZlSfkOck23T8Vdb19gouw0HYs2OnLEHhYEHlA4lwj5lBv
/hk1vwU78EHE896WqNxpjSj6bZZRC460Xxv6aqTt9cZRMvmqI8fAThCOoyfM
glAagPFWN7jZO8M8W5VahK+/HDuR4X4Nv5arotV4wSfP6bdlDnFW20lhejlk
hr533ykjfGTA0QcXVLKnCP03j/bVuAxucEGBQ+kOWy6AEPa6yNA+xPT3IC80
Q3/qK/l+/E2POcJugVlVIcTwYd/P4wFA1ogFqdOjJ2Uv00TpgMthRwsXoNLY
nIcWKhNnixmko/+ZwUlFx97zSbFg0HyD5hKGWQuwxOUHFhkEHi8JaLRnipJS
+lKkJdv5rQRcyeJ128kMKpqY3OenY6Xy0go32VdZf8Fk9VTcUPMqphT5/3cN
dWo2yXjUME1JO9OYkBtqTgAKh/zPpN0XfzyOFczrTFRDigp5kDGJaIIgFe4I
cTi8vybZsDl81So1IIAQN5rhPsWzQQTcL6E7A6X/EIX2OpZyRV5oF4w8hGZQ
8LqAY6SyiygzWxaHsVJbuMpPrc2FTduWYxylzdu3M5igbCc62VVE+kFEuw0M
/oThiW79V/zTc82DwhNVATIB/FulmckvVxI4zANYc+WrsDhFPeQiyfSuP6hx
WXLNVdeiOuO/KIJMATO1sTDHm/xSmPky9eQ5MFVpCK7kveuzHRnp66MZRmqQ
LK+wCKx1dIFGDcwIJdiFqT2JptE15BHS1rBaKUO3LtLZZxZtGj4JkyO2PRJx
duCeFhWNnkMnAF9hteG0AS/uRrshTf6ZTWkRGnjRAZOqf25oCPDtoIgh3+99
bMRM9Z00d2/7DQKf6z1RJOO0TFO6/2Z7/2o3+pB4M8pwt8TTZ5U1+UXf4yvv
EUic2EGU1Mde9eRTBnlWL0In8cpvkm+UC7s4mmuew7KZClymHIvynkomBoAY
PaeeLURWq/d91Ma7OWPuxPTDPRTm06Qo8M86ErS8AdOfNm0pGuEPVKZ3Ipbb
wm7GsTofR/rZhjdomcdefDrHPWKmTRT2lkQ46xfIKSa2S8NlJ5l9BdOOCUq1
jttlsgEQ7sZjmVZ1nsHd0PB1ALX7pNf8+YzfrXD9mNyxtyq0m5jXaZLkPnRy
nL1VFAZYqm7P2Eu0JPdf5zx6ddj5mWdKGLyqcJpsoDlWdz/2AOIZphjNuBQK
33FjQ5X6l7qKpKIU5zRWlMUzX99lulwX/OlyHHbeWF23LQIpP1BxlbAJMBeh
u/DnAg3Ljdnj/Hyd8AmFN75wjRSQkeXdaZnfhZMa9Srs8dkcRdzbmNJsCLhx
iax2RLwHF6n5uRZ4MQ1wZr0FzloaKiQ7NjBbH7BlsGcTXpijgXuN4ayFRD4e
58Q02EYiWjZ3a5pCRTFvFP8hxpIopErjQB3qcT0j4Q7nkJPe6PKgpVEUwxuf
yb8YBxyQEy5hB1xxNQtfLdTe8M2RT+kVFdg5ZUpelZBvpPRb/YQHMXaIt6Ed
G71Q7IAwu15yKys17/JBHkaKtZrdfNRW+9AN6qHAu5Pl6bnIVnxjx8ymc1T/
WsbrNy1awA69OuaXq6Wx+LdYngUy6ZTGbt/9dtLA2yfBbfyMl7sTz/XFP2bt
A2o+dmbpl7TDHJx760ePXhcaVWWM5K/hSN1PlG/PTw4mCuF7ZeTlRa+BwV3Z
241c8GCvyLs4G+XI0Ke1znHnNqpIcPUyO4pgCxFlWzJUKOb4w0U+fFhjjaJp
ilTmPdiZtVUbbau9Fp8adv3XNjQ5h4HYkjVgOPbC1RohO4dsSLVOaRFu9nWX
U31RE8CqC+OKXZ3BFcUyRyZX5MjIsYC2GXNUyk0YihEcxBmZFq5kp7PEX+vK
oE7XNpIqFSP0avGeu9IifLWpQqtU3HX5z5J853TY+Xec0pvKfUMg8p/SCVtv
JHIDE5nwY/RRcuOlsLk+6SIgWXh5vUA+DBFh4YLk7O9q3WRpMpVOWZueSHX3
4QHyLdhB4N+/6e6I2qrWgMeSfV1DbNmykmNVHXr9jypKclA2oUwat1eGXNe/
i/dvD6geqB3cup8cPRhaXn3vv1X+7lMT7LxQQFyAaqNeDn7VC/69zrnLwkJB
Z5GItEZ1FkK77FuxaRL/3qGOumvyo5yjxpeAmqMOyCgH6LPjAH0QahrnNdwS
TegXPrfRvjOxw69rQXzd8DwvcJydJYzi2VBkSUay0uOazX2LXR5yKfhJj0/o
B+t3ZKbNsVRG8W3HigzdacCaNmZYlLnsKKB1Arx41KRUEKopGbu2AOsn9CVh
bUoi2/nCqWF9Js7U7CpeZbSgxpseUTlQ7mo4Hk8otpduJXPgoeEBLJ+ihBrv
ORMhSolZuRNgcgp/HkfGpddlv99nvC9U1K5D3fslTkWckcyi/xY0OsM0bwnV
PeR6KDHl3c9UOf8Z2JF/rnFj2RrOwgoXoCaYDojQ6ReR9Nvss/0SqYj4zB9C
j0UaNBTSabWwbRW7ITAjJOYLCz0QotmI5HEsmmmORrO7CfUb6S9m7BlNDhu/
USpUF5BzygJpZPFuC0mlvqNCHmaHLr3vmJxrngV8ByZNr8nWiBFkEFJHYgPp
U5IX7ftErWuvELpAoyZTKd5Gv4yTx05H2Wu64+CJHgxbtoSHZMRPq6XZd02+
0MW3EAWlIIpVgnKQaI167I6Sn/AfRdLgiWn4PLChaPQ/CCQ5XLVWKX72zFNn
HZUA286e9MOWmrebcBYCu9+TLcOMjHgRnzBQRzuOmo3XENGv/9U066Lx5ING
6EgNMe3HUPbBC40/PomqLrlLs+V07svYM98cMLBySTxPzjG8Um9FMvXus5hp
g9ITWdNQugHJhTD449yulfcM+nvuTiHql5UZW0+gtP1+z81Dx0N8Md+uY8Lk
w5gj96ZQ8sc7mzWM5/8rdcHGfC9+nEgRL8YYtYmI+dkG46O0XUBd7JdL+QXF
9Hajhb0K1sk30SvKuH7Cqr2nzBXt9B7tAL/JIFo2c0aiE746Myu6IP8jlRdj
U3HG5o1xn5ArDcceC1xTB3oJM+ihh8x15r5+OYcm2qScbyAQpTMJ1rawNSbM
/tWeBmINT1aVkjcvYbvsHU4Hi79td7m6Hd/8l6s95dzYvYVfMpeQ/0yDljJv
JhZRhMYX7ghiVn7zrRO88Jor1M1pLseYUHtFlCPhOhYEhiyCsqpFu7bUGqZc
uHCAHinrdaEw9bgi98A8ZHKp/KaWcoS7KyIU1YXxq5dYNlXzjQGQ+H3ZR70W
sBJduPActEoKRlM6xx36NPMJa9UxyJpyCXN8M6upRXDzoVGTCXwjkzFDBInN
k+m3SNQL26NQ5Zjin0IJAT7l8OrrlLZgOi/sdTIS36sktBbqgvZZbAucQC26
V9F3OY0qEu4GSrj+JwM4CFYZdVU/qLwjz0k8Nmm9XXhl/UTA0UJWuIHu1ruf
w6uHKv1lDGA0prZltrbtE6BQTJK+cOcJoodV5MOdIZAqXgA28GkmJlcO0wgK
jAD4/5f/48td6oKxItuP7C9Vu3La8KpJe3K6TxEmZy2muPlaZdY5LVQTMouy
i24T20ArYVd2D0bs6CJstp6FuHK8KXp3spYIIYCewqv8dwiQVmb1twW/vYSW
bAfmHUDmuzVOmh+4emnwDLKhrSEwMkYq+a33ZzAFTbSUE2DBEuPcxF3S8/gv
S425KoWW1+JJ6wNwNPBbjnOiT0MP6vIeNj82LxKoxtHbYUx24fr/2fAvj+vk
fPHKhxDe1l+RLoIhDxuAARvgrfifPWBnihYH18wNNwnYBo/n061Lk69oUpQK
dcwCWxgsDYp+O7s8nP8KODdmPbU5rNF1IdtjUN0v1/e+ViWpZLukFTQ3SepQ
/XVPYbyFLOBpw/UPPvQiStgzCMfhw0l04Iys3vNpnn3eWJQsC7vIphuzD+QK
PisoxRNLfoBgt1K7VYMCBIxONck+UABnKBXMGNObr+OD6o1yO2oa6OOAKphB
i5FevlMPfu9lS9v4a4AJj3mhlTkDLaypE5jg84X2wUpGm0DkR6WfLXEZXWar
xzxqMdA7yU2nYV/4vlPo6h6pMQ1khFUaymgxOK5SDEYDerXRVJnZ5HWjP14N
w+BctVq2CEvUJ9gXQbi+Z7QvEp10QhSGavkDvVKVvs+/zqyfXI3DTVdwfBG1
OKwTbEvJGPoFHEuiukhlGhlBURAspD9yW/bgI3CBYhbSVXEFLW6P0od3XgeU
TnJWWzyWAfbOmauUOS0flCrsWD53y6dLIv8Qkyh5gfs08wsqkOrsuzxIH3Iw
qTjM7IKhx0ORYyeV9P+Y7JPHuSt8SGz+/7JmCXam7a0wlcoSU+8pHAJfmYsc
nYFYM5Lhovih5myXLPrQXlGdK3NdaJQq7POc7jCVBPpKzvKx06rj2fnj5GT1
e52SVPRx2GyPIqZ/Yu7urKHZN2EJi5QSU6txze4YeM2Wz+M1JL568rPaFhBc
2GdHWMGF58hkLlFtL4uSDFG5W+7jQC0qVSQcQ7e8kiZjebbRy9YorTHzyI3p
Ai1QASIZIQHn3Q3w9PtnYATYOdj/fSHSFZvACfNmFh1Uhf1r3IAxmVUdl7cU
eY5DUNE3WR3tzRERTOxh6BlzBiQtC1x7oMLynnlrZItIOTBGxECyHdpj0Iwi
jMKIoVQBvIp0PNmmvKACMmtMiEZpJr/kxNSfvjyI/nIDn7Ai5jXxS4FFrJ4V
VGsB5HqSi8fg9mx3fP6ema9CB2oiVx+nhnF85x5EPYcz6tuuAw8r2CKwVjJ7
65Lbivlex16jgmJgLAnkkh8HHjwWNGu6GQgub8kB6XndG3MfTFympKT6q0ut
rwrnsqmBLMO3xS/So5By2R08sPhy3PkPCGMiAbdozPHiGD1drCPRbClILYfs
xc7psZ5iSK+4uLbH26ZQ9rOJFTsyde6vvT4HLdyHboJYVEIBlMJgwMuL+UEo
3iEoEBlIeqqA9ryhlZjuRGCHBST6MVIQ69q7VXKrxUKOVq6eJKJP65aSW1QH
OP5A+yXNc9Ym7j4XE6NzaflRNLF12YzZvQEeBHhZZEW4cTAgHVDXBW2/a7Dn
1k0FMyX/Sedy14t0XS7HH+sTSV8nMN09J+zKnVImEReD1mebK8NeMsOT5dn9
L4Za/9lj6z2N4HtYrhQS8Vzm5K9O27XWou767FEVbGKZ9F3poaDjKh5t7zd3
PmN0Dzi3/WiyCQz4P58T4UuCt6f5yz8AjrOTl6ACjV13DCqR7e9xqYxF7fGt
/Sv6R/deSQA+Ipg7EE2b4/kESe9OPAuwt1ttZxbyXIcusl0f2KTx0S2+bnOz
+M7WkWP8qqCcZD8vA7qXrnxrt6eGH7RFz974hKiN27bvX/DDvjLXaZT7uO3C
kTiUDxTyaQO3YYL42SCHReM8zt7zKslkmvZH90iLAlmNxQZaYfgF7vh/sNu4
1IjKQJE+5Vm7mZAHnLXNd5BUQlmnpjAymWEfUs7T+t2U1LYW/hGMIXxCeCxF
dN4PJA1BjiweZgb2EnPSiMJzen5xAsKGAlKMlc86asTBDOK7fU5bb0xYnGd6
eU9QZqqveC47T1f/1z1iWHmnZxI4+raB7VkEakcgE9NOW82hcUMMSfpRZvRA
aUGPVOEhfwBq2gt9sXUFTNKQ3+OgbggL7DkS7r7xEz5BUs458F53OoVNKKZs
ryE50CahfYHAuSrtxn11/zaSZaBzbaeVL2wAPOiFV3pKZ80zg+JrHa6UlPoo
7GgpD+S0O2KPtmr46LcXU685kP+yexAfqIgoWmCBqd/pWxXE6L8bCJrQF3Ra
fQvu0EQizsrs29yayHDEUmMfWtrDyZ1DRUjX48XAAS0SnouAxmUbRt9UmpFF
S/G5M5q0MRrY8Zdro2AlnEzO7bX2FJag2cvFc+sg+QGBDD4h7AP9DyesOrGU
Y+maF/04yj9Hza69Xie7Cb8rTORFoeSs+6vIfzo5gSwvc+6fowFdoWg4ZmMi
8JqZbzHFQ6islLIMOIOAj+y8vnJrUR5/98Fgel/V+jDoNfEoabZ9bgUiC+4C
6ntaDEEmUiwU5oEcgIgXtuXRR4nKaCm4Ql41R5vyaB5aurxnJyuLxLtiPR4H
3EW/jmKb3fbFblT2pyGwEXYwfEZSJWqkBOq74Ly9ZrNAPhvL6+w3dF0dRuhW
5CWfLM7728cJPGDN1wNlLme3kdChGG6PiRK11UGyd7MgPyjtSfLtN9Ak9b60
CVUuJlklJ+jsapr2G2naDOlE+3OPQMge4KQRI5JYypFfE2psi/uFm8oV/mUz
sWk20WbyxQ9MPYzxU41OqnbOnp6VDbQSJllW15VRqHIRr+grPs7X/e+fs71G
2iRUvBFFBkJZ3TtkzMLcFMxdSP2HucFHHbSiX/R1zEhDBoMX1sRVk3DVz2G4
pNoDMbPDN5vEmuOgQpDhostKyvu7DFFw1X7QDye78UK0e36iCaEknvSLXeG/
TNqSnHRofJ+1ZqB/Zdp4B5MCONOkpJnF8aEax0hbc+BITms9s8Z/0O5RZFJn
UeVWFjQDjG1KA1GeZl59/FHPFCiFhEcjcCMgC8IZjvbcIWdoO/a6K/stSGXO
xvsMKH9UOCXWZ4VgRMp5fXqTn18MsgqX8Rl50fikBrtCQSQJMDMojW1Ezz43
PVRqytjetUfu515C08M35PheLwDo8y5rvoBCiiaFID6nr0WbcvTJWMX8cMzI
4gqy4nnEKMmh70Tdc127faT/vcOaKjnxTv5juL1scBJCz/dc6k5SI/qbzV6C
UEnv/FZJfhhsRZHzNZbXUTXU1e1ZXnW2PfNko+STZp7H3tunIYYxQ7eNrnFt
FBSjp3Y5+Ysr5Xh6DQeEdcdktjFNGWvy+0joqiHIYvdi5F4JcN2IY5PdP5Ba
sJN14VwzSWqlDIwYkXmNAMkhXHdPmsJjnxF4mR6D56arXlfzxPhGYlocHDqG
/wldM7WB3znDBUfEwiwspdNqMdtKl7Fp3+ozo/zxZNPVZR7G6WPXe1Vi6u3a
P+Rl+KdkAZ4cMh9XAi90wBkTCY+1kk4+yF1tUOyoTA9GD+90XC2XRVBTf8XF
u82+LRsBAvMFJHsyYiy6c1tO9IFGA+YLpikx2+/7Euicfwh4q/tPBcDAWOHY
y+M60NTH/9KmY2f3g1zwoAi0Bsq/qRsKDELyoh9xGHClu0Ete7Aj+PULXV0W
di9QI6Rw6STXlAcLuaExHiO/32XMJEo3oxxqlSwGy+fU+XDOc8dOPH+H/uBS
ZtOH97l897mBqhBJn97dg6UOwGfFPvsBJk6Q2zGfRutHG3s8U2Np2P5inpnz
9mdkIUR9vQGdyB+t2DKpqABDOO2ULPimFVjOHPcn+m8Su6zXOvR9UYw6JB4f
dNvK5SrIi5Pk4mrnCP/BTbAVwiz1u1ssGaHjEsrWirGoywHxbbQEoXrbMMIZ
kzhGSbiDjErkc0eODx5xHymE93wHO7zNucDBRqXJlmALOvOXjvFEom0XVAoA
XUtHEwrssZjfJqvwuE6mXlogwT2bQSQV1b/4zTyL+Y2thceJHlxLwNPiSrKM
BFTWHeWl1QOcRu6bFOEUzaslss4BrzWihaO0LdqSTcD2eRZHzH2+PpTayqre
dQ8V3XfR72jTgobBzujDkoIDJP4HN5M18VtH8m2H6+7F4O7Dmsb6+/TZSp3L
Upjn+Q2nGYNWQn+ZzOAwmWOFItiw2gbZ0UYmDSnsFdwckOnf0m1bty0HAWg0
l3zgRi5KZCb1SwFO8FQVyR7KyB36Uvm7HL3SB+gpGQkmsLVC/1IAtABxBVlM
6qBM21EPMHpxPeb5IWnE/fal4yObwEu1xMzTHUDdKKs5dnwK6d/LluocMnSx
7GJU2FGkF5MH8yZ+8HQCoZjf5LKQLZ5RkRIbiweI8ASspsigQTHB7F/IDYxR
lfnzYLK/A1HHuUWv0mHW+oAbgh+gMNhYTR+AOp3nOGpDQjdXvY/zjAMXl2ZW
ioqmqFGdDt7H5eW4LL0MxW3WJJ7MxQCqUB+bEaCnOkrpk17nQ3Gd6so1OxoT
AMHJLxwR2ANWM+4qg+e+OastscuPXlcZvsqZ3qFHpbzzXO1OcJcWPSh7yjyC
2EzSGLkt6vP0Qf4iuaNLbUVXTtsdZzi+xYyGo5kbO8WFj1hUv584Lvr/8C9B
5ELxg4kGKBV9QF+7yUdaVKVDXZTfS/TxaICN0ndvkhgqhKLVSgG19eM060aT
0kiKq/u6F8+Sdcx9521FQn5P3gJ9+y/bRV/iV/TxgxzrDnubrDT8a9DiM3ss
Cnm27UNXPybT68lGtg2x2ew1+mX3EAuHnIa8iP56LheNBq65xuAfWn/z4lKV
oS3lQJMEsxq5yEZzM+C04OqtoY/wA5QZfyPQgNEVyymeDB4htnK1RM8FQ7Cm
54C/IlIjxugQIcqVC55b8GhSex6mPRNn9YMyxS2oUjOGovPaGiVvKJSncKIc
nG0eJrO28Ht0t9TdsFLmTAT94B9YJ+J8M51ntQf37J2aWaHWD7eRysBbOFMU
qNFlggRB9HtUZWzRJN1j+Yk1I/+X1UWS2VlZxERtHHWv5To7HIA5fj4T3aPv
7s3KekYmbP+CTMGCkdvp6Nc65E/mA0QIaib4zoQvvPzxXkJShcKKl6+OrmMH
Y4eoEX0svjr8/XOMKT7R+69posecrT/s3XxVTKH7Xs3C65f/z3oBRsFe23JM
00Or86MlIEbwIlrP54DS79QlirTol8cI+4Wv0WNOsYt/dtiMyZahOCaY551H
md6A/k95249d8SwTTPJWDc2oge1ugvRdoQYdre62ENqUfzGDcSMJYy7Wn7ed
1TJtyIPagUp+GJvVQyBB0ydE+Uzsmuek51a5twBOYf2eqoBNidx9/me2xNj3
moL/CVLszveuxNp65KzP2bWcFw134unYQ2ZUjeZFN7rFPcbAlWMKBcyRZsIm
s/wr71unPaCb3iUHO2SqfsvBwtNK+rog/z0wG12KK1CJs9H4iiYQTqfY3OUh
Fj9WL1+Y37jCLC3db8jF004Flf3frcD6cVfS+mxlvuznLRO8kE0uyhF2P9nE
cghOn/gFl4dbUkAqxB9GtnB/Ylt0L3VWQbpKa4S2tl/OWa7p6IadYoZFJLZM
Jjegcg7ZkNWxSp2XvBJfQxAUYQy56TzXS6dnXcO6gxJZfFSXA1U2NMZuTo6Y
PpYvDEy6YnGYmYXP5J2LHMZj65kn1ug6UQFMKM8Md9vBZ4MZycN2sc23uHb7
GWHT+R6dyqNlgK5wPUCmrwrSbSmvEbQaeFbmdros1KPl9MhWOuBE7iMaA/Ix
YcLZeVpAxJw4aBIpBtW/4SuV7V6GEsrG+uiCO/5GH9UZEZ3l3Vl0niuRgGCV
7ZYSK8i2m92Y4wb/vmsvMnjtN/C0EkgKr+B0Pm3v3yaxldtBloYEW5PSBCNJ
RkaMvh2u0SezL85/KjwRBbTiaX/AT9Lux6aQSjHNJb0nt3BRnL7vQzwp+kGC
dQ/xzhVzVasoJ6nZHm7D80oJzaaVAJ1di8S2IjXbsLGPgeYe7OHv+/PED6qM
FCE2IRdq5qvCXPqnyHBYNhXgNkEJmVmg5p+X8qivO8R6tRpcZ97hMU3wTYOp
HR/m4duRKIbkyNHPDGIdjXGj9biK5LwvIbsVqt8Uef9o4CzDo891/7y0/y7X
/CHNfFK4rr2/45XD44XR7DzokvAvR2wSt15p224mahmJQpPAM3sxOaogtN9E
4XVlEokXWKmxK6gel93jRWhMF11cbEUMxriGb51giWuUgEDe8qeh3s0cQMPd
3tK8bXPMtGNdNVUhd2P7tU/sBoF0IG1CRVlcQ+wCij3UTgqlRbc0Nbm83Y2W
XaqtMN5EgQyRye9AtbqRsIj8c0PS49/pZp/ZjfXD84n9hJgGtDnS+dhrj6Bs
MOFgLxR0Gp4N0yd2Xbu0nE0hkHlJOL5iTKaUoDJ3Yp1xc8pl84fNsTOU040p
GZe5LE2Wah03VjMGVCtiqKLn37KkxhXiGn9n/3JHavkKpyizG4s+ybnEqZZL
jpbEpcpQt6IQWkwLA6l9JPkDmmombmV7HmScZ08XBDQVM0jxT7XUXHSfLHxJ
ZAZFrDse8V8ycrxRPXRFFI3D5gSvGlf0DBSchXQ3rulV/WF0SzICp3B0ZS8h
pt+8/bWXFzBa2Fpm3UJRntuC7WB/0jLxfs08BqgPaW/GTioIhiCdz3lzbzDX
awa1WO4KyK7YDDkoUY6EdM7aEugfDwVIZA6tnIDBKFRO7IvC8gEWbcnl2PPx
UtiSA/i5TJ0+3z3Rmh8r7rLBxSUTuXHC6Ixpg9gIw8wH34tq8Ok/UTdb4SeX
YVNmG65C0l3FDA7+lpWSEINJMII5ik7C5Pna1z5+DyGJuNBylgobC4SPt1YP
CuZeOZcyj+/osDsaei3Qb+/KlVzbb1vUSwlO98XEIG52UVs8FaVxeL1Dz2Ns
kbg1Vj6NhpoXVGa8geZNC+bumOFF2yyfiDw9C862u7LGgWTET32zE5Jk1xmi
TMSfHGlFtZ+sFITBDTixqOHShFkq4pNOFMbyLVrOdOtIIraitVcGrYN3IC0Q
BKHWg1ii96KZsfMiH74sSjx+bN/+2Vaf8ZEsKTS0x3hV9DQ67YP456L3juNr
Egw6Ui6vINXpbIdEcn850aYdkMY9CRdGFXbk7I1hAvRLcF0H8Fjqm+19BMvc
wiskqOqCVduRz/VkzjWBILo6Z4M6vArO59S6D2t6UWg0z6aUWBf/mAvd7gyu
ZHi64Tk+8R+WHXSKVOhiv/v2Sw3+0Age2SCrvaBBOc8xGCl5wO/NKXRtvyNc
KWv+xSVRV+axbQGDN6A20Hxar3IiRVVyWQjK/e1+VMRC6Fk4CMcpR3xM1jsS
LIj9DQ11FluuYlME+lsgKSXULyiyKDYvR/4PKUDYi73Xvb0Jc97W39gpMxwO
/rkK9uVtabnC/uMtA2VfrkJjxAnn12SYSHyKkS+l6F7f8mdpuHjrhvRUQKpd
QmNYsSoM2XJHwebcqDmi0dbBEazzgrC31FwAkc8Sj3I9PUsN3hPBxo3mdaSo
InNzJrndUr71awvzhzuSbthDk+IAs1FUNUt45mZbZDxXo81kbNU7PuyzGHco
giuwConTUQbKp4A1zZbBo5LmTRhh0itsdTr8aXqXdpFmLeYM9Tp0WoAU3UF3
Y34o+s79wy/GkHBNSTiS49BetPCAdag2fZGJzQqJam8hnrinlvdr+J9BnkA3
Lb5zQM1lR5mT8xzcvLuQuFdZWQ4KpnYr8L8z1F1yv0lFWVFzdPXc7UthNqLG
CusG91Do3FQtL6jl65A0nV8muyhr5wYfIKYD9QX2FdYR7ZpbDQ6UtgWbYhnW
gVEgfvRxat0KxQ1jt9MYgpi7dBiQx8VeLqGK/cJO1SjpXRRDPQrBENLP+ijN
oMLzaVU+AI1X9o8aHLqLWTdc84kH9GvRpqlp6SkJkHQTGRApL4LqhhLsBcOE
dsNcf7wqgIaQp/dnHwpgB6Nd7yXExn0NbPpkvwANvu2QZOUEzECBx6zYk0FO
LAKmdsPK9p6PKzZKYhjK2ZvWOLZt6kxanZ533r/JzxgBNicfKbRUngz1sjv3
jWJI9jSvIly+hSsHFA/I8VHr2kJA3ulk0AMojyPRTrKcmuiX06xitoXThpfs
Gzr2H9yiJcvsDW+kdOugjlI+jfi7g8cs+nT8u1kzxN5IhCpRVrb+lgTNP/JV
GY1rRvClJjafyUs5ERKodzb/0Ey27kakKddEWZeAcFtmBJXVlctMaNfK8Mr/
d7w0PeFjfjcoX3IcOjU1AnHCdFR/20bGpy3/xlaLjC2em3xJY907GGIksZQH
+X+AUXybBn0tRkg+5StKC5jIRGCrs4FVFlQR1RkOOuz4Gzu8tYZNJ4dhthQl
zyu7+VXbDM4+sB/0Fb67f56s6Mg3RYpflcsVANdR0Pt1aKNpa1ym/3Jpf60n
udpU3K6YT7M1Qpm3dXyB6wVJ4MD7+YIxCSyDGiYOWGsuWEkyoF/Yp+VeT81u
BYvwGB4qxzT3qKD200TCDBkiTiPg4hGI9nJ+IJe/BaICZ5f/lpwVnnhcWgTg
tnRI+HoA88ZwELGfSz0yWC6lSOeGCPq08UqXXAZ/zzP7qqRUJyp5A8opC13/
JdX774Hp3MvYeVJMiPU1ELGmIHFVtifTl9UvlRQqYxFRk6jsdhMFIZNT6sL2
+M/qzHzjfGDa5Yjie//lpmCTdIM52AfBYH8ieFHaxVAerkGQ1QP61QarG4+q
H5lfHUG1yCRnlctJLtVy+rU9dNZ78/BJOI2gfuphYdgpkQkD6Qt9mUAFhAje
Jzp1vItJR8JFXgVIiL5weADmqTrAJNoo0kpXu9jo2zDGv/4sAzCsl1IehAQW
jM2X3u8V24HrTf2rt3m8efjpy9247XLjcBjK2XRF659D0kqapoUeC4rqX6I+
UuwOicHNRgd4nU673/OaZfmsRDpAHiHwsoQeE7/meertgrEWlEj5tGI4vr7Y
khC3Povgv4kdOa9haQxjUscqaCnYQ8X1ddGamcT9yD//wUMMq23jtEPIsV71
7+zc/7HEIxkir2AhMh6Az5l3RUNZOx6KFKBJdxAbmMsoWjiZD0e/ePq2JirW
7HeLOMb0Nek1XXdQ2Ixqa3pJ0a6qY0/wbpqZ+VQTL39QgtIO46jAJIPURAP/
Ab4zTC2P3M6k3cV0ytDtraPWS4DqcccMZ+ew0AKqnj6XbWI0yby2fjLxf1Mq
B7Q2pvSsoGTvq3mP7CexrefOToiBWNMulgLItyvkpVmFIEmmuXLot8/F2O8B
ZM6hRWguGTEJaB7830ZfHpxY3TCqt4ipxMQaacEiUYzm5O0gZU/sANs6r/GE
sK5o7zKqnGxwyWalbbbHmMhFYOGoBf08kdRKoQ2VegR/KFUZULH+9QB7Zhwb
XZUhsU7bnLCaAklESEBTiilBlmLt/oC4GOOK3TsNiZIymXal6qjVg71CqG+I
LL48G7ab9ARI4KccKAzlhQP4k4JAAkK2l0Le9Wpz3sMc5t5Wu1BOF/ii7nt6
w6VgJz7u89UAZDk7ZzRk8g63tZj/pTAdIgwwac1kZyB157o9ADRA1VT/w7hu
ypUhOqBajnhHj7ojv/HidlrGOfTj/WzAfhr5kCQMeDeJt23GwEo3JkbmuNqg
r0ZXr6Sb2jLG9k1jP1qzsYh/71CjL5vfafMQLl7VL9ioJXS4XBhuUQYr8sGI
/GjYJbFzKSlWaVanRDfRfmLnvKI9+wLoDEXiGZXAe2i07TMGW5AshCHkyuC5
ZyuRRMrg4/Twkh49d3CH2io0ziRj2C/Ox+LTQTVGy4EU0DRwJ4kK5rJ40QgA
z+ew/wCPHejU51OxAoXkp3RVQ/i9CzdbKkNyrAhdwt11Y5JiRtqItf/jHU79
Ab3i/ZRdiFeWwuR6ZN1whbusQi6fgsNN2ODCPBFiEmXgOb3xn+03A3IrvEtd
TzIJUcc/bT203hxZoU5PemUYtBA79AIkNcXWkW1CEzY3rUIMQr9Jta28h4Yi
865kv1G4VKf8fpRqy2WIIMCd094Ragek1pZ0AJX+JnvBs0cLQas1HntWwCSM
7DV8y1+p6sHEAumgHH9f2qrvw7hLQn2ERBplUfPBILUe3CcVJuOmkC/BWmss
Du5gj9rP6Z9ZXI20mrx1hO/uxKbpaOxqCjyOF1yDVFkzwwL/z3RELh5EASuh
8WfzYTo+QlXJQjvXcrpFR4FSMfBBshpzs/D6ak9LWAFXVc9/yTNKWnN+VvZO
r7DkYBbP1ZsqMh+YNpdnOiNd1f32/A3dmZP+q64ep7Nip3nST3SUBz/UJcLx
x5NLXE2qiXLlIKWcX94AmLaTyshlFs3OdhRlZoLOCnvKbsMdLmjGieIKqj5B
MyEEEQXLB6iwF8QdXl2KxiffW/gyULMnCm6RHYMPrGqiinhw+icI/CbBgn2l
CwaYQNDh2gb0BYd4dFN8GDER0VHnP4AsIZs3KmQgdakVJy5fboPFYFl3U5D5
VHhxroDqs9Yvu24V2yC4CTPVpM/OD25a4w7zUl1Te0i4JRuwtGp6CgrLb+yb
QsTtXG9qqtbyCR5z0IhalECMpeEdmeVc4x/yca6t13nGVfCMe+Pf1ygpprU8
1bgDs5eJUXUq8CBqM0zY9GSwbl5IUJhgHMnAOt8tzmOv+LoLNrWBH1+0363B
P9BZ9B+UbH9fv+5dQZGDUIaYI7sACOKaE9moVCmifUHlfMbhJ5w2eMeuWWnU
DTjgWT48MjGv//QB/2a9hf+s0Oi5yOh9f/ppC2YjV9DligP/bCCZsfFC5Yij
str5GWpRYaGGaw+jXpusCyOkHHshja+nZuIA7UYcuEknE56y0x6Vyp6XpJ/4
Y+Q9lDiCy9bZXKdQVEf7PgTiD7fxSL0HygGHPZEhAtIfLruJpta29Me5aw97
OcZ5omZixUmJafDKGgbslTCfaQb1ISN0DpWhCp3Tk2mWcb0C424cFozM3waf
B0wl7xTc4YS4DNxFHwlC0kWM/Z49Fpn1/DtaiPg42TY73gb4Cnt+1Y2QbW3i
WM0ZuyZtME0ar4P0fB1Gmbi7mrylust+BspM6TF/Mp08AvYZjc/09ZRHOQR7
nlDIxPcOuapOHQ0lPtXxi/q4qHv0NCfDn4o0VvE57YDaDu+Vv4Iuc2xP2EHA
dkkgUOQGfTomYyxpSUPQL6ZoVZOkSx6JCFZSI1f7LoKB1s0l4K/ZGBb1j/Rx
YyUzg2211qmMG/chznZL0oQPsFD6e+hNgUJLjxP9mZBb+pM0kBj6sYqEy1k2
ZSKD2shg+KidP3HKTX0oE+j0kO3igVeTuGJZAgGHMa8B68pKAhfk0hD6OFKr
x+5/huXpl+KsDhCC8NUQVUBa/g3FwaB1cTeTSsrCTzWLsg9+wot69uvAgOJ2
T3iNprdilrBrmGN+YP+sAWliqe6Z9twZ2yZ8Y1wbdksvUKjcL+J664uwItdM
+9RGV0CP2yDgRNvP40gMlIP/iqfiW0yg16vNJuiGXnlw5kcQhnIJ49xs34Ii
KdzP7ot+MtZbiQkUivJQnovYv58/IrKU9Re04Hryxe+B92TpILOavQSUNI+F
2rVNaonryTBWbaGGXZB75vd6JqOu037DYIgtidT/6ua4l8ek23PLEeyUV6yh
ABlvZEUslpMXvn6SqzXsMPjMiFbyhpBF4LI6nJqwhPLWxv8CNnvTDemU1wZZ
FHOMBUCg0EB5jdd4YNlpC2dCVEFSxCO/H5FKhZ63lb8QGE7XyJ4YlJoFpA7P
QnYAsxEW2+ASCD2hiMmX90vxiABe0Ym7nqA8diG4WfspAzQlzi5IJDFWrFI6
HNJ/gErB1L+cxFZRCiBr6uXgKw2De7qmTZ28oh5+aEpehdsEzs4O4DlQ7aPg
SJ832aHv4FhfVLbs4GUwKHLml23Tv5kZGydqm4AhNPCGcvPd45J5x9HJKbjj
UMg1ejcqS7nsR+eOUIEXPUDUD7nIPL3la3HiVmmk6zjIyGhoWDC5d7TqccbH
Qa9qVZqQfK0wfaWXMwva81lXqyMn322Z13LwS6TU+mdgYivJmTDEuAtfnFkA
HxMVTPmQoqd9i2oeaZOGlTobexd+DogSVtb4wNVYMp/PhUVqVmWE9/8Tz2lv
votcmXgV99heQsuwxLl/q+fwwKFy/DWOI67sSfIbfFtvhS8Rt0/QYYXJ/LmE
+Eu2VPktnT6nOetLLtOrMj4L5forqgMe4m/FdtGpwcBW7gAQMdljVMXlsbys
RklPaGVi4YtR7UVMRkc3O7Lh0eeX13Ga8Mga9v7QCG4q4cYc8KmXQRJPtXXS
CW8L40ZxmWPe1rlcA6mmLpt16Z7paPrwuTpKnYly29RFrJQAhMtUOGIDQWuO
ku3h2sRAjsrl1mB4gUmUhQTERfrkbBzP5cvhOSAqq4Lgf9YoVny2EbeQmJLN
xnZT2Prvf/6y95rX/DSL+aX0IvidWOFSWpwzJIlyUZV/mKi3hjW3ieeba99y
xansP+IZ1MSv4eAkK18ZIYYaI+Sw2H9gutntpBhKeZS2TCtIpg+b2tpSwK+B
FIEwU1/8ZETmqTERp8r5TVBUXfsEbxLnjzbnRh/Zb3/C/L45n7NuMlVrh8p4
DRRhGObBJtvZik3izFp2j8LwyzZxp9W3F6ZKRtPQrmTL745OGS1rJrzbfIWc
gIyi3B2d/GGt+Y9+UolpAVCYyNPo8ZO+CIil+n1/U2EDef3XI/HfrE1E0qbu
F6uHqjoWPc1y2RybOVXlZTQQCpQwrLQWiQm6qOY7tDmq2Jc8LltTegRg0C0u
Shpx2zw5lzjgN/EkSxzMWTWvfvQxXOwlPnZSOaHJfjhnJmUUpig4w3b/0Wil
ZAjmQXFuk2jntmqzf6vDuYAXrzsE77e17J8T9c0Faf8YD+3/GRrUBQoEL5E8
H+xZrNFGcj7uYkF6t03/rxMOPyoYN8X77D4AVeAt5UrilJVIi2yw6+MQ0eRg
ljmio3yyxcpzot0lcV6ciuVKUonPhgA+NGRurCmioG/JK478qXufiOYyUPxN
V1p2jyiBHSpqXKAtU7+AO0jkCHLVgdly8a3RnAhaEgMEqhL1929REvzVVLBK
tCqTEyfpS6kszGBSqlPMzFpsAIBsOXfWKaE/+Mbpq5Plo67FdbgtCTq+YL+N
gYUHnevHRpNOq7GZ0gR1ilMx/aovhWM0SXtekMe9Yv8K3ZVOJzPdatQKHmSd
gLYqm8VFoKuaaUNTD82qpBPxh4oM+/bpGbtY42vlz6zZfhkbV99jRRymPvJr
anMrc7dSwGhO0fOqF1H/vPdeOubtnRbOLumtJpKnr5OwfkCou6x9kJL94w0i
ILHAGZBBy5/GCStxUJ0H0UzptgQzHU44zXovhgRNiubV10y5CW1uIOs98H/Z
k9MfjdD2sQqZBfCJe+pshScj94FUrfXQYfAcw87drRcNwOyuM2nVbmPC8feX
ahmGDUt1ToD9re/lGiOrXT2wLONfsB7gl8T3dNOCj8YQseGHkVL1+Eq5sdFp
zM00kqJl+zXcczO9ltygACI9/p3yjyxev+CB4Z/cPfR6vzsdhfsnzV/KCVMp
h2o3V3I4sGLYRnVnxkCiqAvFmC5CRnuL54XcLNN7M6QHo9lLPJJ1+EuV/s+u
D0EC6dDRBm6A66NUsl8atpt7jxQ5xghmpFqkeJtPFnXZG8DxsdTeGV9LQs6o
t79SbV4O3BkgiAeaPSa2epQDd8knwTHfB4T2SSPl/2IoqxnY/5lMpKKn82GS
V8Oc7twWD5XrtmmszQfWbWn3oDguqplY1UhiyQlpctyaPE6sNf+lbGYvQS5q
OjBpILgb1iNYLgB+1VZIqo9meIvduYo+MHae3QHHyH+SOR7NefFMi3kSRQrU
UH1674rh0zr1uKPek7kG/vd1aRTRzwUGwkB8N4d/WD1EA9c4l6/COYWWdVxU
NuRUWOvk1hAl3jKaX2Lur+FliXAX45wY/9JrOi6jpfiWAvWBdh8xpeWacM7i
AdUdOopfwHZ9gpNfuLRndrtTaLUSx+IlePcIn1Fa9fO0w5kTCGsseivQ/0Ug
vJ+F0dIGPyW2yiX0b+3SMFMcFhGMp50RB9zazGomCzpJgFs1lBKSDVibxS+A
hibayCsTH/oZ4SmCB1aaOPDZIPa10Re7cSJbJrQWOkfLj2DsYFfjwVrI5wOg
WCB6eNcVfLs1sdF8ASkco23KmN1kEyt/ztdj2IPbTPUYWi5pSR0KIA1K9FlU
Uq7ZTaWXP9EEtncPKOgjsxM4yvPDNO4SkARSvIj5E93BdvIHPhzoflqjV0Sm
Bp/n98+CsZ4scmGXfI7TLOXyWabDKpp0TzyGzkzKBIeJlJg77PbVvRxuMlqx
g5ngTn9Dham2bmRry1RIVrNGNLsoC4CZybTK+o5YRoNrBKGOFZSRbhgFxgaB
/WL7TayUmt4ag3aHpYAGK7AiSElGtgv7+dn3iY/LVuRejYI02umpf8+VKtRS
szhOsz5Lsn9newhiusBRvniYJ2Fq/4VJDGi5/B+b+GBy0Qs3UegMAqOZllkE
3M2ANTWxHq6ptr4sGnI/+y9plf2aQQKezNRzldKXnvx5DICJiozPrDco3GkJ
/xZ7O5FKqMitJiWFBV9K6wln+m6hWngZPE1P50YTFxYo08IoR8uh7jcBFnlB
oBPLa+KxaBKqjvO3IthVIqhtfMouUXA8kT4+j7JCMoiMmNDydvZHAc2ApfxF
wK0W1v043mePi0Z1CLpStRN4nKTfQJSuwt5d7Msh01tt6Wnz5com/88vrSQV
XsUWTUE7Q7ewU4mLVH+cuyySm4AWa0LpxxUv8VfVCkxpxz09i8Nd/OmKUhbn
7AC8d6g3wcMD14gWPWpxm4DZUD2Ci5LBuXKxjUu0mh2iF94WCnNZvx8Pexua
SioX/rpxNXir0thfJ5+YrsuJ7WxiLavwodVz1GS45JVKqWN6Iu6oJzV26y+m
Nwuc2jwIEG/RK+7LS77QYmtccQB1T2fF8QJqg08h4e/2Dj5Ogwn/LbYuirMT
3y1+sV0gWIT/WRQ910pzG1fSb+VeD0+qQn6pG/1VX5saoZbb3XHS8VG+Qq0u
+ySVa4RQc0JWRzhFO3ZRV9AM32wOJqqtQ7gu9ucjd6nNDb+HZN6hiDRK5zFR
zEv9n5DeuiaXxebcGnBugPrKlnv6AMVpRlg3ZTA0reTsmQW1vd5VLD41o/gn
qkuoWE2SnNs7HFrhln16FsQbVo/qnG7wcBm742XHHokztOzBt6Q/wGIG0qOo
naRQGeSE3NbqNt4eJ+TlCWI2wXNJbwrAvFlX1utmmCLjGPTG7Q05owoxvQsE
9USwLhnw5nMagaYqOsWTI3aNzqEzYHlqjku+4KRyR8XVzu5U5cw9uw6MOdH1
3PHEhe/P2TPPFCf8EPcV8wPHKFMwlx1qtBe4RPPcpM/u0LGbBIWFBfJI8LIb
Zf4Kids2KAc+PV/wzJxSWFPDDHOgepurKB07aveTyPiRx+RMuent21TmbRXR
hClvBrQ/MA2uZBstHNEWEcbyYZU5g4pRi76N16P+PbRZTqHdX9vWU8S4ZOb+
5tLUO/50GPhouTalxqaKcD9HVanCCP+eI7k+90RIN4PrVZN277Fw+ezNHhlr
Pw4mDIyUD/kfTXNu6EpaCkNa93mSZHS7/lp9BEVphwehmxBfJQ+yq870Culr
54rT9JQwM20174ZuRIiRACkF6rtBfZ8kH3Otp4b7epRyKSBofj6AV6BKYsPu
xGltcC8njpfjR0Qm2lQZBzMxugL9pShnwhP9XVYybgNAG1pT3lOkAzXx+R/J
AxifDwHNafQ6rgGT8U/RZUFnXj438jfFNhbzFFori7BKr+iQag563IyUcMe2
NnS86ox7I1m0cDYvei85ebGjpQuJ13YTTm52tZHP3X6XMI08Fgagpkoom0gC
bhvve1Dt/Ab1qtJpwvTKtegL2+Dr46i3OJOFT+GPPUQC45nsN6wsZYXoxJ5+
newU1TBw5sS5XNz/9/YIX9lAJYUiKaZl3XO81ghn3t1GUhIxsVUY3iTEZ5g/
OS3QADOFo9+CGU3SpAay3oTxqZfrWF21i4crYqWpLYVZeZSVcYiC0wDbKwZz
AO9nuQHUj1AMcHqpdsYY2GVFijlhWljMulKVxIBUDSMFEmpD/734eHyFsYPj
QK4q/qhvX752dLuexT53YeY3nflN1W+P4k+jPqvQHX/i4RZjxu66Dtwk49hJ
+A9Zm/BFnJX+UqaaFcqaqWTC8K2g/RWG/h8peuMznMkbeQaIQgjvosfrCJGy
SCjYIHDUiCuf4B/vGUJX9jRAS6OCauUb8CVWpU5Qw89u0s/pYsDRtaWxvM0V
s45u9gIHa9rpn20gdvwDdibSom+anFzEtB5OYwaATVohicdo81yeEirCoPUS
zzYGTjEmzxCm5oir3GHhpnrozRoWdynk7fPXtPtMir/4chnTgAJnYEXo7HC5
ym3ynYSnftKVJIWZh/xECDI+09BxA3LX8NENp5EVx4HcuWPasWCxOHliZ4uU
5qIwtfu1TSzuQZlGtLrw+3V+UbrpGZ41KfMUVcUbTcESZnfW8DIaRXSrWbFh
K1SbSVDN8VNGP1ErIyX9vLryRtHA4lIPbDLD0RuDZgsuX+NO2YxmjX2gLYUM
HgwDWS/Yr9JY0nkObqy2i9ZbC6dnRVm43eWoliyztRDFVVkZOWFE/df5gKpw
WcwFqhLvq9FrOZID88eqnJjIneFwFpImsBj5go1CXmnPDIHIvMfPNkfmfude
yv7Aa7GCnukxsDO7/YOmV+PFb5c1rn4wqZ8XZ03ta4FUG5bfznSImZ762YP0
z5voh8aDr1yGt2JAXIsGNzFJ9GDjnJ9LslHvuGpZxfTYWZio3Y1ufCKFr5jv
1IKJVNHSrly/bpbmaCbRm8SIrE+dXOSxjOFVnWLJOSwHtWlkKfDhyv9LpZAg
BpTptz4v8kyljVZc6fz0Rt0z2GurFG+Dx7QP8jjlO31SYFUG3baqQ9Vgkgcs
PvuskUMRVHR1cIvmOINDPUx/Kqf25KG9uXpGrrLWNRNdfQHc58GgmBMYMYXK
TvC36rH6s+cDJnlJlW8ajsvrJW5QipV/wdEFULQlvmEg9sJskcdHuNT2yGS0
W4QJDPsfvcA6E9dFLdde4MtLuKt7t6zslyhLGXAmjW12fgbGN7OgiTKz5KFP
2D6K10EwZMQxFjrH54TfjMZ48dlA8nJY+zGF6bCljDtY8ev5nfdhTlTIwzJq
fToP5Rc6YqYTSwai80RUiwMF5ERjJ7SPW8U4n5AxDthpS6wKSAAUJDKspz/P
HPnvHNxttAfDzKMw5dTL+hou1tVES0/8X2EYCEOz4X0Of4CY5qp1z2dfWwlr
t9SPX1r5rqiEt2gzY5McUy3jZw4x69f48NU5fkpZuFIXlKPKXYefoUoDh/mu
eRqcAMHd2wzTWCRsQStcMM2WibrOGSN62TFjZNhx1H0Rw5OBAHjOjLnecgiX
KJSU6xzG/LFZPqfGoyf4YHvW03IRd0wTgy1C/FI8GyF6nCNeTpscSOlsSMFA
T2MkXaNXvAl06322me+G31c8+c+C5cyPKFKxqUEvCSkSUad8CFYIJtjFVX2E
dp/wxLSe2tLU/o7d3Cx8f816oo4U9Sj/G9n850QoHJ7+LygOLrX13QEm4Kmp
uAOY8URjV1uopDHvzKL6q1uxiGibOfTcyskN3kzBG5TbKn86zDyIIWxym7+v
vtHHi1uBBE1FcvznHDPI19jEuR2luzy7Th3knHBlCwIKVGTzIqXa37TMFnMQ
yFuSWEE5IZkStmCyvvx1d5C1kdOFeY02njikfpRVudQNxCpFlm7cOZzMPu2I
RnYwRTXg6w6Uz4LOuPMN1bUEnuDygKNKxN5HE+sMyfITacKyYH1Xo1Nu6QZm
8EXqbBrlDhLNloLZ5XryI5IGU2L0qGIB2mXpmazZW1tUksYd7DwWR6Z4fZDZ
Eqi6jqav+9LnY346z6oMgw6KgOuudYU519bbUvzUKaol8LTYt8RYypMIBz4A
U1ZNxAKwVKll0Cl635hCYC80I9BEQnmZskIPtQIDgZjOJEHCqN8LytG1kmij
HI+anS2Omnosy8m0BLtE+qXeVVLKhZ1PTZeS8/ArXuOj1hAe6kXkdk4NL4AU
5eDsBEDbFuY8SbUobEmkweRxhjadXPKefHPo3N2s0o0nBqQe3Soa7gvKs/0U
sYd+qhG35neQpMuiZD7zt0mtphsMavan6z7B9tYZaYoO/uEGrUzEnU6s/ucV
4LwE5DOPl6p/qgCk15r5i1bzXiJhRiWIyN14DwNo877OT9nYDWVjDY14OEOY
T5rD3DddpNsBO20DvLeF0BdnowqG3r+nH2dP5gm8SNU/Dfuxqk9zLSqiNRCl
J6sDvJViNHypLUZZZxFyku0vJsi5Ok3RWoWOK4iHCoUPAngoln9pyZxQgp3z
NUy9TX4spSBxomsLD8sDhf5HJliQOlk1a5Pay7gVvIyBCHOfzYV3waIr19Zx
aN7DaTiJiDjyE1gTS3WUHD0jWXb1hyN4j+W3v4UyJuN50kYqikZ8cxDZLHoE
TYTUoLT/xor9e72a30Zp4V9h43qgT8xmnsX35j7DLo3eDS9EmiqBgucxspvu
hINa0EJcRPFLXAV3aAt2d+2CsYyIZamaXDRMB7rmKeO8rS4U7prUJafQ2+g5
9Viy6vqxzX5SMAEcf62pUCXwYU9/349hKgo1bmvAnY8EQayzvNOFfpaR3Ecf
1dyDJNlLZeHhe9lD6W8HJMQbIwGRhPxs+y26sAalK1/ik2Jt2S5aeCu5Nzo2
pCubemm5ZsdeUoxdy3eL7VMxyDBfoCtzBLK3bGnyIYRmqBhGQ0apo3X0oBVd
xHKEIUEvS0ssv7zYjshtEHaAvKP40IYkrSfXu/B8Jgw3qQoyzWVExhJzU3Kf
uKQ+XnlH4Oyc85DuCEnt8aysjNvP3Fg4sp55nquh3OJHtN45AMe4gNjJxTu8
Tr2VhxfQzEecL2FGN54Slfoy3/VWT9T2gVd4JK+f/fV+WMIQhMNapSH7108l
j6l2KvWF72r3N9HdfwwEcLWhVmFvJABPbdhGhl8eoatllmBNPUVOUQc3QObV
vu7lcXIE8+Mx62e4c+ygsKqI5WAgWpq//B/FkPy3b5oft8aNs7orCiq+KpWv
S+Dma+5bMo4aNS4ejEmqukoz8YjfooLpzXYxqRmdWVJYkFZ4icFRhsNJuZ8h
Zg4gCKoK6wfiphAmN6RqLkni7H/HP03cqWCzxallXfnq/TcEoyBalJEQLacg
oQnwActrKndu0jl6NfO+Lrk6N25BK5vu4wJc68CRBH0H2XJU4ZHt36EqsnzU
mu4sB0atc1RA5vzQebRcUsCt8xSGTV/iADRCSxDK+C91w7f5tvmGwto2XQts
ATdX6tiYKoun2e6bpsnPKcdVWYO/bwI+IQ+r7Iw5MOQ+WKzgHYzVYs/fgm3p
muWQlOcl0WL9quzwpi9aCuAWkUAlM3OwCvWlUr4rB0n3kv4/rTjT3v9bGmS6
w+V31OeLRx2OTcFNzkCRpmzgS6zw7MzHzXNcgMTXb6jHFmAzbBO3zyn8N/v3
mSSMl3TFKOknc8m5lOCcED3PEJbyBdJWp84sfS6rmb60QJCYYQ3hwsJONI+S
MYmfc8HnSXKAv9al1n+i1d7jw2UEe5ZR99o0v3y55BkjVoqk2aMBEXClze1a
3rSVQYxR9V/piaeSD1tRxCkMEYBLuV+2I2cqnEyfW1hNhapIFUCCStrrcdnp
ZrQd3cP760Y7b9zQAONF9XYxubOS6QAyv0bXa4cl6fc+MI3+iOveqAAg4HJV
qX6lmf0RQL+uWX78jUCCV0cJnQNkGrRoid4j0c37NJW9H2CMX0wiRVU0Xmj4
8Gq22aHsFMPHKcbCQTGuHDBZVORN7tdYF/JPBuf6r/uO7lTFz119p+TWwVKU
KfCRvwJOXq0FbQDCYXZWDkNCvvf4YoatCHvQpt4IeJ+nJMtr4KcZk9XeFVz5
Dji0I2s5FHjxuRVKmME6kvbJKL8SPlWKCut89v7/Er5fE/I8rYeQom1OxczS
hRIWY7yyR4QpnKp5CYBC92JbsGXYQIezK5LWa3CoAqQGNVodXf2l1QL786Xm
m/coqeTFfsKCdc0rGpgM/3Cxqm0KvJap+HuHE4OtfJHzpofu6LXyFIR0LwQP
dAOM8jCQWzqwRe6b6JQraDL34EAOz7WPWx/lSxVB1mqZhyao+Uo1VgGRmyUg
+xq2r86dn98yaR1tbsHZNFKgtFDl2Bgl7b5IiUDnvxaXwDsPXb0BC5y66W+T
A/4HfvO/xX5PVJQ6eRiI6s+d2HVPJzHlKoinSNaIcFKaxQU6/dtkpnOs06AW
BGwX0E993Ls1vkMXkPcjueCZL7uljeN3rMPKJ7p18ld9PvVfueZehaAAj8CJ
c7/RxCZ6oc7Yu2HHyV5j+62Hp+tzFi/gJpRNneoeUTLR3QT4VPEnzN4vYFia
cDGirgK767QvOOAA6IPGv7XlQ0hawoBhv62/WromCrKsC655EY9a+eKp7TeD
YWxuUn25jBoMz1Kd1qBOSKnzmzgtsECgskd24mXz5BgpTBHADCHX//aZzlcn
oZfsT8P/0FyvwLAFJwj9Yz62iL7qrJtl6WWx5V9PuqVelkd/MWAaKW/pzVm0
bEDlLtS8IL98R9diFIWoTRWBB+bmrrVgw8JwA6O0mvGZZywPf0m6RY1DzE6g
v/gFQNnztUKJo/wBvxtW29RkHT3kKA7g2m3JY26q6gKpZ3pn/wgUorj7j8rU
kFUIB+17aUAG3HPs8r9Iqj5A6fwMIQkDxcb3nLrhwqOlh3Btyv8NujvbGjrb
KLIcNZLwyuOE4cxmnzpJ5J7Ovlm31p3IMOtgIYDKSVOk/TBQhRONm1OTk+Dd
QMV1pct1JNIY9lIn28qo7O70usjhZS8mFOIDtL6tE8XFFoofOeWh2SkK+xSN
PfSHrmPIYIU/M7uKrE0DQ0aTmRxdRZClA83omvCWTuWbFNBKfFpAbo0Sdtvf
j3yB1rMg7mAXMFEq1mgYAnAvLAjGk1H3AEBAgmyZqBOQSOtejm0kqbus4u6Z
cK857F6DndRQ5jQwO88P6qz3z5YGr3Ah+H3tUYEblMywtzp1IxIb+Cuqsecu
KsP/nu4O0GesSmafZtE9LQoTweKjB63sp2s3GMFbe0smahe5KSjkMHpNkjJS
5tPHdGVMGeurA0XtObq9FXBwGTIrbej6gR4XXoKPnZJDPQqhYTYvD/6IAG+A
psm3LMAxRDx5XIDVNGjcoBKtzUI9loXJaqm+z3YqQrOMsG6/S9bzNsEbjlkU
PaCMF5BvLa1UAV0mWs9O3U+R/Hk9jDkUcxyXmm8ALOspitnKE+XH0FQ4uurZ
4dbxuKhFhBpfL55P9b+ha4S6R6MkAaTX7pBpedbWvDGgUSXjOvK4GYsFt5Zj
8AFY2uFDqP4TnOxnpstFkVbnsxC2gkNG4y1kG3yVmKwUvdO2bdcfbEnhl+oF
om5G3QOxqqIkoM/IaqEG/aWOalycqOi491Fh8CWtC77NRipcm0PdkKo8mGRP
8+11MBSHcaO3ApYQIT/o+n5z9hlZM9NPOcvuH/AlqUzeBo2iBMtnYmiP0t3D
gunqEHNPer8NXdNzhRyOvPO8lm0pNRr9uOcs/ZM1O50uMqySfkU+yK1vCVIE
QaUugY3BL/yohtaQpY94mCwAFnjJyfJYE9FpujqEUgi8qLiiIWsrHUEYR1p1
POoaAvpzVS3XY29DJKxkmAwpK68QcghNGpg8+Aasl4vT6vt8p2mg8KeJaX1d
IBYXHhgYGzetbxwiZ7SgF7mhbfBTb0Iyqa90SCkMbTMZBNMtzLOnMm2VnNOJ
UzpHXIOk+M77MOrdb6dW+FtnCDrrMZagg0Tkrqy4gqKr3rAdNfkDCMhwOEwQ
xWMAwTKdZchx20PfRpHisMCl7iWN50O49JU1KkKFkKEu4G2K9h7kfhDTPL+n
e8BvPfrNZQNlADbWO0CScTZb7rNkrmcX9jOWaMwtaMZ/8eLn7alJtl6BrHkT
Jg/FjuuilDm+0z0Sn12o8vvn7TtnqflErBCkP/fHaTX1QfuJGV6FkOdkpcq4
Z+jw8biri1e55VDjwseGZ7pAhm1nVcqgWncffE0wCt6Loue80Unh9EHSKElG
SLIC8yFLTRz8J04w35ybvPz7cY3cOgy+zySGvU/9dfoSqbRm4ZGmD+wFmjYB
Lga+bknZPigNw+Accavp0phXT48RWcLA7U0VSY58DwwemRP50WEiyKjySpw4
7rB6ciq7rNCmwSPniuvnnYq66dC6JnsNsXik4/SFGoZUtg81HOcDKTmfrK5m
ardGHqoBIrar3/eA1VfCknLuQoSS32+uHoNexGvewB4EXTMiuw38t1sBLc6u
Zxl9pDTC7fSMLkA1u4+bnLFxFGlTq+Y2l9Ki6+TOUhgyaGlkC/l/gepimKeg
ze6vrH8SiFV3SHCr56Ymr1/lNBtKl4/BBkOQNkgaS+ig8Bl0kfry/WG7XhyM
cMrC2PC3Y2AUhwPVTzfGezq9ytB59z6PBzR+1wm61iqazjIFskpjZ3GLImOR
h9FLtai/WYNsO2pQMgd8nY2D0RccS0oY34frfOeSJ1A2hKhVhaGpi/wctZwC
9QFz7Wh3e2dG6ORLvNbQhrF0T9Tnc1RNTBwO9klmdKRRyOvX7jBR7Z9kJec6
Tutg9q7w34EdwW4b8kLp6fUUh00dXzkqoG8/oyDNgIa6SsOdHoOgrHmY6uxw
d8a5FLBQJTATknVLdWOvqrxJkAQviNkCkOCuz7qJlp0ifzr3swEm745H/Ane
m72pU0KvOA0dNryx1Og0vOd+ao47HXBkEYzszlFNr2zE8e1GdRX3SMdlqLat
BJRE9RLpzfSqUWrS3U0+ODHwHaPY8IJu6nAXPmWRUIG9oYGgGQbWIVs4L07M
S7Yp1Y183mkqLUBOpYz2uIM88pEIIAW/uVUz/2QzNEPbsg22q7cInXRcHAD1
JCrn5mq4+3T5n1VBD9nyWBgnU7El8WGwIOmRCbUWlkfS+4GAUGcxNnKjSHL4
4+A6PQioML2P6eF7yPHZRRN0mf9PAl5IYBXlI3xiHG74xBrZLjV9AGL/EkGh
e837E3TNbjpi6hM9poa26c83PRCG3d0rI5nJADs3Yh1zpTdf9stCrp1kiR36
qnN7Vv6QN+gtpCNgncia5ptr0JAixn8bn/UFQBLJAUtpc1jJGPlCLVwv7l3H
v9jMYj/m3hkZEB1/V4b8/rNt8moeIe6+XPtnntJ+Qr2t05n1PmGSbUa3EAVz
9ckcYJMCBHoU1MPcl6MoVbLzMbbXMNbcdjD90vSc4aQjhZgUKk8bdJo4n7Gy
Lhysa0I7KIj4z85pNQvN/kfyrZy/BGI5drVAMLu6YusqnuGHCbCa1VIcHmdz
aU9jqYO/jfMBokufo9S3HCJ+sC9A4P0wsSSXfhWPmpdI4BFlRZYaFacOElMm
Y57mk70I9/DBaVJk16VhtfqmQMiYHfbOv3NTsmJ8vU6xslctz4H71l9UEjI6
DKcbgPUafWqzZK7ENWLzCi40sfOxjVy79fzHonT29uRJHZZnjdFxlN3Ik6Zs
2Qg/jcmAR1TEvXfW0PL+nyOq7ivbYKq/Nebg8hPyvtz0OK+0yuvPoImgm4aK
9DgaBP+C9s6X1MPXGH8WTXqILQ/wOKKqUEiBB0STSWMm49PoLW5psxBkjP0a
WFyxur5Bsnc6pK+yX2LVbJfqeFbGRCpR3a+AaU2r/qVotSA5Yy+T0mbJBw0d
gzfu7ATqefhQdSC409OD64eKTQm9gjctDr7hGBMNx8c6xR0WM3nX8GZFhL2q
+eOQzUeNkgCv5aAopvQ+QV14shOvqViUDw1F+mQv9ymApB6m0SWNSC1vZhxA
n1vreXw5pGhyXIbFT0LNerJMEgtdHfRnEZr4EGL7+ot94/cGpnmGVizjzQPO
hLjMq4EDSyeNh5twLaERF1mRK5R+NfLWngPylrUfPYPz5qoq6Nk3iMl0YWpB
bF/kGeAWwYpPxUnuKXstVVkZo7SDmOMaFH8vZP8S7RvV4M/QbYZDbmhdNnwU
w6YD3JMXD2QiQVN4wFnM8JaLs65yNd9XE9qB0uXTknwPdqA1U+tCBI1YWc2h
uXbEh7uZKxHEOL9PLhvH/7PO8EDKnoX7UGkWXK9+ESvOcA1xQYejj+7lJ1Iu
Fx80XmpknlYVvDQBLDfOu6xFAe/UF4Uv1cT6s2l+gxM7cCnVeO9uzgo3FagV
CezCmvgEMjFT7gyvPgpDA94YqSJfvuZAu4KUTpE/spLB594ZzkPhn20DOqcM
LxwNTp7HWAKvYj7uzu6Mo9wWWJyrvI3gVkOowsFo21tyYfa3TafvI8215k3s
/6vpnUXKByUG4oEnMmAm91/cpg0PUSKN6/qRVU4pc3eAr/SYMpXKnGQ2naXs
INmfrwMtt3XpDzhtrMP2VtWH6Lv/nxaB7i5PzvsCa3KDveNszFmnfH6yq4Zy
hal6C55JnX0Dk5kbf5BzExusjuCPhW3S6Sb/RkStM/ckjV53BIQVjYeazI71
RMEEXfWzAe4h9YlsnSYzenc4uGR9d535f6Fzt6iypIJ095SPWZe49VDUnKqw
QetsSq1OQwowcCsqkdrkNIdofjgV47nqMsOp8mlArYcfFgQ+Kxc9qMTarK3+
yxMvR0D0ba/wN+zYtBPqwqjLzzrM7BE9ewVjfJqwz7XBWNlxSyRSz3F2koem
5HBO+umgOXyWu5rvRAkcUNTYSZpBggEf55C+X3sQ/r+z09UeZYIo/+34pWQe
leQf1FRK2lotB6z+cRJ+Yif1O1lQBim3ZlUCEBnmqZz7zHg4mgWToSfIdfiC
JpXWfFW/x75G1y2gu8mqdFgNndNytyw6evvzx6sS4EKf99dx6541URzxnCwf
kx/Utc5jKoFRxjF8o5PTK9e1KH7aSyuRbgeR+QtHit7rVNnXdkoWeR8PIrNG
7NjcxAsl/JOyUcV0XgCuAQCzhqFYlK2RsEpHCTvaG//NB34g3U4PvEWPt+3U
it9KvBpg3tV39OqGjqWu18d1PEvb9T3Efj3DIZcogLD72LxBVLZnUKg7He7y
+h8W22ElBf1oOJ0Fz4gaQkCDRZsAYn2FggF0veucMpwx7kcoPi/CVS6IbP08
92c+DETPlgErQoCm6tGSWWwPKuiNVnIBhZnLvekKDHdLqQaTVCY7BbCB5JU9
rZlgaTh29u01zWLRff8NBhDYZLGamIfoOXg7YBBs6xCeC5rZyLhzHNi1PVeD
fLf9m2vSDdafJ1UpLavDYZ/xA/3MC9EC7foAZJjUrxRKSSlVq1DZjPn7iLRY
SGLV70X+KTyMMVwDzwz8/3bB2NdxHg0b5IGyz2UHoBySGPmDlkaaTyC+3csL
AH6Kb6o2YMqNMVUKHGUKDmLwU/HLS5EDsdfmBbdWYjtSVbeaH7Pq3RiUygX0
5zmK4NtM2mgq/fL+Fzm+gOIZqlPJCm01k0Pge5f6Tl0slCAbrRzeZCFbFIT6
j/QAquzR+3jWJgoY2QmAn1At0T9Z/Ul/i9hiE2ZKoBx71ZyTt6f0PrcMGybE
2+gGyxurYhOXrZErAOvCrT/2XBGjNNMFU/mY8Uj+Z1nKSeDnFrnxO/Yr7u7b
PV+tsAldW9K92vMyzA9zOU4Nq4Khd9GJy9wvFzguUyFdB7C1j944c2h8KRN/
GbBbzeLOHYC4g4s13O9/odm9yZ3g0e8OsFo5rRZQmbIjp3jwMiRoeYACYnrw
mJellbeW6/3eQHHltWi0G0jVLclc/0jqkL8+V8ptUBNwSEtvF/DZXtzEFpLa
KaH1jSpHHJytZ10IsIzXoiMAt4/XKmfMYHtckFwkW3JJwVyc8rAx0E50R+zV
AZTQQnev7il+1SLyVVhkdF2qnZuoS0eqvfFYzZBKAWSIas6s6bxFcKOu/fie
0cxLVYpX8rDvy0D/c8zHwF2k9zyu0G50QQFk7oaTU2LvYV9/UFDJuQ6CaAke
6bZzHFV8hHebZiTq1vYVTXT4GRAcWtaYMVYYcbsk2Aa7llITzdf+PuEACThZ
mQr3pubX58bfu1Jkmqyiib9x/4p2W9/BvkLlbKc3e6gcl5L9nJ3F7KE+62Mr
dYVlV5jpGaOMtfltBRK7HX4VO++VzXXBwg+i8rGdVFEvCdJumJ0eorNUqys8
DEKYx50DH6cZtr6ckX+t89FVDSxSk992gt55yLfMVUPe3TYdkk7S1+0SI7ip
9mi4sFNFEw/iGI8YAiEZXhExHUKoYyN74L6f4JBKJBTVfMhMkcSn7Nh8NP3/
zPR1zOTXvoMCLCuJKXYgvuNTeX8tT5SPHPEqg9QPcKq4hiwTTv9lmtXUEqZu
ODFvYQo3fj+isVnZwJ3yW/dtF1PCnK1Niw/SWS22FxIek6cGXy5ssae1rt5i
A//5+bzEG/AysHOZFCeFOdTWPbUj35Dit8xuQ3X70KyQgRgTpNR4g5+/YmjZ
7xKcfHsUkrzxeKjHjvsbaWWNkPc70/3RCAJT6S/OWQXSqdFp0TKe1jZP2oCV
efwolRzTIBBKs2tv7fgUJCHL02BMuJsy1AvJE40q31xj5s+phrOP0OUxfxQI
VB55HtZp2sb946NsMUn1j3ff9a0BFqjhBNBQ98bpAskMY37gAbGoOFUhVNIJ
Eiap9x+u/Byb4L7B/F5y+DgJ/pxqQEnNU/+ecr05+7rdRtgiW0sy9y6O/uuZ
KDNhfMC6pcOaMv64kvfWAic+CiQv+mAQiQafNKpLZVWuxsxIk5KAmxdjyMKN
4DSQIjl0OAHMwwZQmqBFMQ8xH8KvbalLgKfw3xl5SRqfvdliOIv6iMA9rwrW
ADaDm63t/lJY925wBK+ewqeeuFYTH9tUI0mQvG6bnG29cU2RKHd8aJOcPChR
1vmdqxlisiMOCs0u3i4nVD94s1ET1XVPyQkG7+2r14VTPCpQUzWutI7Tiov5
55ZJdzksk1eXYxkcUHXUcc8sb0Y/hvqis2JWpA6qUfaHAkQOAi9/Cmb66hkB
zBdCe3KUL8ucEA+gduqHctzt4D2SSWn2MII8hWJyBRbrGUP6HPwaF1ws2xuv
byjhDUJuvIpmJ1I8OF1Dyk+rxOM5iOQ7kWxr/1G1I9z1wogTQ81NvUk+A9JC
7Elra0lIdvgsN1IkottX7wI4jJ0k/xR3lccEJ2dQaL63jEIPsL61lQd6v4w5
ZIeC6hHBtB51iXB2eGCkmNOhQo2/Tjtauc+iVS+kUfF6L8VL6Z4uy0KVpZvX
i2wgKKJiRzZaEbk9X/3tCWVltJ3u3Uhgq7A4i/2JZ7VgXVnUVSN1pZDb88rn
q7uFLINJFBWIuEDZhs33cBVOWVeRCnChFt/lYGNMtLYBY2wJFRqCMHGPXKmN
/DZ6yveS/uD1E8xsHrLFyXpGs/hJvRo5h1EZ+PDirbUwNfTlAByMwm9b0Kgp
RvCx9XS65HxqvscTEKzambfQ6yeTGnBM3cW5s3yRR5opdmZE+d9BvmQHjiZR
DzxZNfTQbwEN83mr2Ty8nCjGavcC49hUTVB/Mz4kLTn7KuDxEhSsUtC8b/2I
/sd1EIUFhd6vP9RXMB7bRa/CKUqQ1eJ/3iOnpbCf4PhD+J229t1bDTwMkPpW
lGVP+0Szb1uPCM2eaHred4QN3vAUmAvZJn9erJTkpsT1BnreuUYHowRMqQzB
X/KAjK67QJbuclnfFp8rl+8MIIN9PHQpGs0yNo3sUe0I9qirTsctKG901o0t
DSrN2XBccd+U1d5AWGe71GPYh53xPyMJRFGr0oTFXytX8CfciX4DVGxpwt3e
PeZqJdDgLxBUPZ3wdnNkX/k+TIcZudOTbyUDFVSXeOau3sygKISADLvCflmZ
cGC9JT118oOwAzQLmlJJuTOR4oHkZo97r1zU6T3Q8IoV5Vq7nKDhNqvpdZf1
xhFvVtj+Lb+HfLmG8hohjw8BnsVPeh+rnfHLC7atvXBnvsJWyy09QAcv2ts9
MpaGWOkEB0/MJ5o4lTRWBeSxkI6iigmPXqFCMQtBI23mQNQHEsK9ckPKzrJF
QdQFR+t+z9Kf3Weck1XJKIqTMmPgye2UnMzGpRbnBXcuvF1OWCXTsSYxGwfj
33ULyh/CqopFyN0QNV2CdL3vZuIIgA15whSVKxjJd2vs7SZGZZbrMUlSQZEG
2Ju+q7Uo+BrW+D7xWbcC9l4EJcyoytJL8abT3jJ1aKcE9QsdsnBDgwChb2Gt
ylasON/rts9i/oW+Buzl0F6jw5tA/1cy5YUauQqVhejszucSujWDIRUovQdv
R/sRAxynCmFoh7Uaobm5OwOZF3VDVCzO+EH/WygOVz+CAFevuCsLnqyEunbY
jBINtrOhU1oQYwKIuCF38zDbwXroYeya2dirIxJNND5bpTYxRhBtbzt1QjC4
8hLrCtKoZxpAghDuwqGMBFAb/PLhWoucJx79nXI9i/8xA5yj7MFmDqZflnqk
4BiW48zvAwUG5pH2ZYXzohAk/OXIP7cn4Ntgmn8U4EiPjeOczT4pGw2dbDXS
q8HE2Y9sM3SdX+1q5ps/iA8O8qtGJDAp5/Vy/XW/e4Etrql2dbK1+ghfoRdp
wlL68rOQzqfd8NUayfmiPv9YUjSyDzI6e+qRl024suH3+ycsh+4reE7p40Sn
YOiCSPYUphV9qqq/F38vUgEDwYa9j/cVYta0S/66O/IInztnbzuhXe1nXVjv
9k3ozYq9aviLpjd9pkrcpdA3247rb9JWFE3NneJSjP/O/WypRPkgS9TFPWvD
3GLouVefXZpuuBU6sWiL/5iffovthe94MwOOUU7Flt97aTx1sU42Oz2qfOpC
DwGGFsGv6BPy4ZR57CdgBC44s9MdH/YJhiwwrxOf2A7vnWYBK+LTmfZ2Op7d
FzqKBAH6jvJ4c5mQSLyZlHHO2ABH8yN+db58bxsFciOClWDv5b5tWtJ5mSAq
LkLSAr9UIexQGbd0b/EwqWk+9hs7jPuuPAPoKgXh8fVQxlQFw4Uojb0YvfMr
Eyn8X+vAkoMUUNpOqJcdQncO7ATuq6jQjTw71favYjHT9Mgaax6WQLFBlnJ2
xfK6yUaa0uccn6q/DOl6th5JsmmHKW7kZxKqQV+gc9et/Uf2NXWuIwDVy/mH
dIl3GSH7wE2+t3Hm+pgHfXERTAAca3I1bsckAXcOCw2Ej0/gSbc/DRceQA9B
DQe5DMs5ZRaPSYBXhl87UMtO8TVTpwfC3h4z5RB1jkV2I/cuTuZI+UdLwnHq
F8WAZyfDUx/I/9H7cxAvkAiEgQM/YIw5rxoDcLvEYqzVu/Xx0SNGO+TpjLw/
ZCxU7a3u7a1zztpCNbciD8Sp+cJsP0cuRaRqGJCJNCzufD8rmVlQtZHLNG/D
MhaNCSClNQaJ4IjqxXuHq2NttSC8W5vAV0PEVrn8/4ICS8RRrX6oWXjq7rHF
GkiYJH1nx0XH87Dii1ZyKDS30SrQJLHK2oTq7PCb+JjEqHToa7vcuHhfzjfV
ISRPI8Kxq1GldPjsyGaRf7iiJ1qHZx32f6S12FfCEDHGne2LVF/5GtZi1RkH
XSv3B+czWE6GSDTjQuCgUN0amidcaSvGUSO6zsSRXnOzHOXtA+6bDVOQfeVt
jHlOlQVtHdJ+GwzGdW0GJuz0oiwo86CGCl1OXzumkAbDZnUVYSfYwTiVx4at
W9MhhPOie1C0XsVktMXiLdYDK/PgHaFWW961d5uB+NqDlrq4BqgEiaakwiml
0WrIZhkBiUPEZmnFq0oVh4HzP1cJWb2XGhBd+nw0KfWBUqX3nnqef7q9DpKX
tbbkJfy824OiNy+SychNZYBdCp0G95MneSSrhfrttqPR2lSHchNgnDC0/5j2
WQWM/s9pRmI96GC5+X8AsrwSmg9l6q90wEia3xhCHb8l3tCKVZYHWVHALVoL
0R3WQ85WL3nxq8/GwFQGPxsqwLw0o5qCmCILBRaOhbv97mSD5ySK53DS/3A5
Y2EKhKPVrosjzpbnEOxFU5PylLnrbdetaJ2sNdMhLj1GiDrABEcl5j06+5IO
MAd2qQ087lXBuvG4WcIuIHtwdc5I655D6i/YI/gnOBQ+m4Pmx7JTSxpx+O8n
2WU2AB326j3ValhAys44aDVSvDyu/EJ1TgIRIVQ5QqC1H1xVovRpXts9LAtv
acIHq+sHZT51HIg4dssDbyf/oYPqxTxquFuv4VwpauGAbI3gNX4D0nooC7SZ
WC+40Uv2ai4JCiaUht26LBshgEXhNomXBWij3b2msGUAq/+JeoSy26wT8sPR
CJZJgGPZSA/OthLhsXWvW0uY6Uzo4U4GxgchdKvRsa4EVawNMoq7bbMT2PvI
SxMFvFTQRU5UnMhAINFwDuHHIGbbNYwOmabgC12UtoEtmNvzY1lePUypYOfa
1aQLxCSy+AaUH4agCgOZvLrvp0MFEOHiKaXklvgqb0agKfsZJDRef8ri7sZh
2f5ilmdzmB/OyBCC6gA9ossasVMvA1hXWIMoK44LAUU0AHOd9LTBLC+x+uBG
AQ2VhI3U5laOALxBfQIVp88qbIbIjI2W3MFRfMwyTT1yXHCOQbWdRHvOkCUx
4ans4eAR7eMeHC/ZhAceqVUYSgc/jtzVp4UEEhRzOuUQDaXIKYy5GJ2gXtFR
BbFL0uate0Dt27c6AhiJeI4pWmhFim8I/Ie+6QedlVWI5od6aaUV3i6GY+Zu
R8htT3Cl4BxNm2PFtkQvFjLPXjZB9J4/pKKyhIO/aAFNGe4TW0BJaMsX/d7u
Ikpyrg6D2IJgB7b5gl3cJf6L9F7ujvCwligQLwAN95+xdWi3pnTyvuPxGq26
u7BPGXq4BlExTVn7aei26NYRyT2IqlLbO2AP4u49oMKMlcpx7L6ykwX3Atxs
zNyJLQWH26+bMKKVY/SrUmNBUPivC8A+SLTolR1OK0X60Zb9naYjxjRdZgVK
V+eOOQChfZOvOmL+9qHeEMOWeNyBd4oLmOulRVVuWNxsIK5GzJXRGMuDZpg0
7Or5rIrfV0ZPg7td6AFDEwEWWKR1Y/9lWV85pvUG1TSXc6xzTvujKQ/zTkPm
Ofcp2D6K3L4k07ZLa+igSJivfg4LTG910ygDLUYwklbAoyP1wYhwp4V18e1c
KDZvJVX2XfAxzozx7vMcYabzZpmDryTtzFgVJ0NW0IFqgij92fM6MNd0vc/y
arI5Z74Fld+S+iYwoc0Th5IxoijlTv+f6QeOOl0f2empZYukYnQcXmJ3uL86
0xJToRM5kJnR0xfABGtsGCWXj23KP10R5cBylcpA3pNNyRQCdHoPTskMfwHw
kWzc4s0b7/mabrUmruvqq85wVPCt9PgGOT+vak+QhpDawnaonmG82jMkgBoy
4/X4H4tfY7r3Udth5T3GyKNW4tHO5c22BL8s6YdxXk3vSQuMvu1wvPIfPZJs
f54/kQAH1KlzxSfpJDkAGoappFLTIK3NrEeKhUF6OXiDn49X5aM0zk8PhwyY
YkN2XnLdrtPUcin47XXuzgCmc5ZN5B+x+KN2ur5vsfB9mek9kqHNH831J9bo
84+LHsh5TtE/fn5P2OWCfM3hjKT9rxqV0yqVDi8wBjNahfJHqCd/QCPkQsbS
JZviy3Bg6y1DkqKZPedsPx9A0k6eOO9boYLGSsCLlEMfHtBxB75BBkrcPAIQ
FKqOnB5cuUajN30rcQGBbG7I+Zs29eoS8er9DdcWv1ffTKsaqMB4vjIxgNkH
3xc+q+bfLKKaWjSGVHQm9jr2bpsLUi++GOIDb36MNASOC8WV22hUxqg+uW5i
/f3bFyyIGYmMnTftYHRtRRBJqShTniOthxgTP88H3OmE3KVLNi8147IaHvGX
KkcTVRvoUVkTPb7Mj4HknkzzIw5/3lbPpbwu+X4e2JBG5AckFmhOAORuCVBM
P1Jt2Y1I/1Y6PrpMrMHMsh0xblbNNRqEKY+gADk4sRAmdLn+8/CMvQxbLDh5
AUp6At3u5HT5vTPldekTkN9kPwq+jOQullUldx9r1FGdFZGTvGWtHDhd8sX0
wmUAvgaF89Im19BV8JoEoSjiamNif34i797O4VxPGeGDS6ETxTfM1ENrVYBC
9OqUuKKhqXl9rvH0c5h1QitUwih2PeKc0lNsxv77M3c28kMWYWfTwwPHelRP
MTEAIuFvXCmNbeFaaXEZheaQHg8GqazLWWd5SQhqIsooqAvh8Zwe16r98twx
ii5laPe+m19LnLlQsO35nNtwPjP0KCIgNXXVlwolWiWinRe3Q1fjURMMWi+j
klHoGUZ+6Dnh2ecZLd+W8Cdz6mVEEru/MujEl1c9lcvp1ezGc9mqYkyZ4cND
N0YrhPFfDuFIPp9Ss6fNj07oXNViKXVUX+r4TehtPRLkTezhJUe3hi+UtTeN
+5/Yl7sKXszHCl8oaArArZIEi4wMp8SQHmIl2RvGRBubeZQaL5PsxLdKLIt+
3XlBGcikahK77ksHux6dCeZnMM7PqHEWb7hHA7ZEYzyy/ZN+HFvlMoi7KdMo
BiiGIbnSJ1gdn3bl4ARC5a9RwkGowsu2B1T5WiAyXnVNJ0C83HgKH2GohqL7
EXdRBDyTuO0KWahXVvyW5kecNzck+bACbZkD36wviZE+7qw2Wls/HI/D7hlD
ConfnaNU4TEBgcFAqMBn8DkY53ng+fw2aBQHBLr4Ik+NWZgLIjD7aq9D6WIJ
GarB7PqcB/AoR0fb4a8O2K+PeoiEqrIt8su3647E2fbQ+Dh+BDTfarJMuxa3
L9rGLdy/3q7KGUYKQuhdRxe58sSSEodo45H1HCT+VDBjDcXfpyl6Kr1+q4iF
9QITMVrwhdMprFE1QiTN56E8S9wUSEdz7/PRk92IHVf7ItAuzBahkXr1nKkI
paIkjxgk/CpXJ7BXQfWyUEsUM/rSMeKKO/l1HFnvr8mnhnArkzgNysq/6ASS
xtXtk4HahwRHD1dYJs2uCVprUdpBAQ4nwUmoSSCp9hxey9NJG+uwd4ssoHum
ZQSKS/3yLaMoEZT7zP9Ajr/kyXXEEVfCa5PEeAUWMECwFSjETUm/hnkpRlKY
U8pQcdGrxvBJIHioKQMpDeQlj7wtTyWu3OdBKWPViX/Rsyl4+vQvoRjia5nU
bOwrVY96Gb/XFuTdVrWplEjHLM+33ADFmPkkIxB8wndGpy4DT5dRLjBNzqd9
ACUmIgo7ULGAPWKXrOQTa/y+2FUow8ITBeM5SwhI9gpNXvfDjw6Joxij7Mqj
iFkPH3plphcQu0g+fOpo8uMDLGGXguBpytBTAThVZwQFIhU6Gku5nfkBbKds
FN9EBpwSDR5CmO3lCFVypZvKztYj7COYCVTI+FhZkkRSPiBfEQJX28KbWKEH
S2iNjrzMq4CIuc6wjfPPEFVN4RH75mHar0CU1Hx4PJTSseog4zgK9gHdHm8V
PKYyj8nO5RTvDcSwh8gXaRVOESJTnjFLnaSjgSE3NIoeltUkvgJ8arVHTTj0
K3qkkherSDFHQyZtn5BAxoI8NrRN3Ky3lCXuDd8lI6q/+mqnwu9+t2kDEh/o
4cVIk2ARXS9C5dMktCnRwsWrLTgmEImSjr5Yrgq59aqFTuoKenYoKmbQ4wEi
oI36KWSy9kcq7ZL/s02L74WSyp2+H8hqOAmFC4617L5Dgt4qcrDlJZh6se87
ib7eEOrDZk3T76Z6+WMHBck+CNkhdk//TuAxBlTUYI6TCYY3e08qOF88tYiG
OC9jOO9JPTxuxxneKKNvCa2MJ5131XIniqYmEO631AUlQjtmf96m1JDsfU4+
t3Cl9+rCmCkweR5nvyeJYVRTn1qG7R45mhS/vznl1/jd9SsRxYp8+8Xm21+v
FIX68cW61Dp/JrTJL53mf9+HAK/PRfxNFtcJEgGWGmZDqmrFi2ef70eFtQNu
KaWZ/jA3DjA3qWcsdypm5/3Nht5hbR4tvuUsgKdQbSJLYx2j3PqAdGL13IYb
RPVzlQj+mQ+QW2aGUzvfHzL5EXIDox7vZcKld/awl1ctAcfFIFVqDcNRYNoS
Y961mVaE319mNeFPAromSvb18i4vThb0myo7Nkp6AFBw04IfPM/v5I0XFdVM
F3vKpeokoez9AGFn/HWn9BJJ1OImId8juqHu0w60hYSIco3Wxua60CDDs/11
x6fcUlxrjeEPF5W5d9yjCQsCOZRTmG2XEjwbXyd3IiyphU0gJXSo0QQPi6UK
kqA67f++pD8aidIeUeQLO6jRYLykZS0GGBm/k9MIkPFg/n67WEbxrVxrW9uy
eDI2e+nqIkbL8e9dt0P2iav0/CbcnOwwVLSKnNy33uDMZGqt+wr2FVzyN5Y5
ywmvUbOaAR7yC41xAnNp7UP+1AjAJ9lqQS2fv8n0wTyNoSFNKj9ajYXaYURj
qMlsZf19EE1aGk88mAbjOMR04JKoHFKW5gih1b9EJsbGWmULZrobGukGEHAT
hfmhOqRtHQPvCb1TtR6PcgiL5VPCxN5J7hcmolEqXk+Vgdgc+TgZLLFZD2A+
jbNR9Wi6vy17vBAeZwKB0TkadpWURPoMqZxNYzNNG5GIdX5/5n+wvvPI+3Xl
3WK/bJZgyAxOCbxRANFtTmuOH7uyZFdrSVZcUnquzJCM/p3lNIqMyVcHpOOJ
W0w1GVUapmHWLUI42ilN0N0bpmosoNcIaVprFWxNZI++q1zj0RaGbK86s2Mg
mb7ONnt53RuXIeWnVCtXy9Dnwg+STnCoiVS06PMCFvgAkScHM1vZ2Rk2EZn8
ZLEd4cZnb/8kZ+f0otQ0Arboh9WPwLHL+q87tPWJC7RgDgUC5xnB28PxQD0p
yUYGax1Rf8Vclw64q8CY492ifcUNLQXT3GYxVxppCgKhEiqV0x8N7be1eIS1
YCv2ILsze7JGL3proEpPFnnsBkdTwpSS6yOFOdubmqxFy72esx+qcMm03g1J
e+Vcpx8xg0IepRMUfNVBRDkl5ulAsAQcLldKsU58zQck+zXIpphs8hpXGMYI
plcF1MoCBWPu+ehVk4amablslGbYqOtN/BnHZ5tIsY3/YSpBLp1GShgGgeKI
dnPyWF8h3TlYf5AgciQh/YbsMD+ORqp9eELwRbgSRxxLCWiYBPzDaizd3lQL
w8wuZuueDRIvNIUMP9FDsucyPkaavcKIl8rGD+oqnsImeTKKEz+CZ11itxjY
/4DGvPYoJkXbjanp0SBoef2Wy+HT0qzu/e9Vs1WBDL2B4dgD4IBTUX1W2vn6
4IR1gujEzaRe/sfY/psdHm8cupNW/t6WceadGhFjlZh6b8Y8G304zn+PM2u3
qfTMQej8CejVvlY8BCLtd0RnYoS41h3E0j3S81kzw1b65Ip4+l4w9LaB1Iek
t6RGO3gVX3FO4iThcKQeHp/ELdurBEzL7ljipXRPaXWY/l62FaA1MjsOLbNB
6++k4HSFkKqP9kY3Dais0NKG/Tn+KUcre8U3baqaS3gJcrr/vPkGfalmNau3
hRt71GTHeyxfXv6vuh1X5MLY2TKNip38Oq4jIYjdpXoNyMoDjnhZyheKCcTs
w9QdL09zUwhBaFbibrPw1RSifKDDq5ZQRH4rtT0awnOh2oISCjjdBqGtAMEt
TFt9wrmjZPGc1pZq3JAgceV52JvtYSRVq84vKOrcIAi5SjuGA+0lrOGJEmM+
9XF1qt8HPWET7lV5guVS25imqNsC883+FuaBYek5/hpteDLhMx/8yzXdsHuu
kiofDneoUGgRwIq34X59zAMStd9KpZGv7G8HqgfWw4CTYL7r1gvFMNlI2xDP
E/k/Zk3z4Bf5+ENOG8zPclgYE9SVz2Fl6mzesaV8X2g7qs5rHjs1DLs/rwjo
Akd1MKH+INxxBRXWtvNYCBOStco02dMSQBbaknNegR+SOfYAhrhDP3IYIBOi
DEWgcVszPbrb3EEylH7SwEXp/Xkpo45amNfDNMUEpzMX9ADq6xgPC3tDWMdn
DnHX1AZX4FSPyzOtPIonCNq+0FbIb9C22ShI4NdwsNmV7Nrdj1KehP1CPXvN
82OM6u+nSoseugVUgkDRDMFxgNwTu6tZYV88paGIBTYzLZocb7MmrD8rM4IR
jL4br1ae/3SwigCfLKpZemCEqEhEaQ1FXPbPBj1p5YwbnlcmfIt16laWLf9c
EjZzmzjrRq3+awZFwzUTSX/J0213EWw0s0Hy5mculfXRAXgIJQTnQdYCGI5D
hACglT+N9cU3ibeHB53ACYmUO6g4x1g24YPCr9GmpPdpfcmyhxqve9uSu2zm
UspypDdujmHn6ymxEIGPdEIB+a6s83fFZkXDaGAXNZcJEsr4XtniaDnl4J3n
6oZkgTVrMp5D+R/3VIXYkCpzso1j0NoontGeKI8Qt/DSwi7U+jalqll5WrFw
9ufOFPCvcUqAw6MkwwVezF8l7EkYBYUmjlou8egvRF+ImHsI1FsJ+JTRVfoT
HV/iVbo2dKLXx4S9iXC0sheZpnNhcwMEowFvcEeKPOxwQ+Fp4hmT5ExY9DrP
PlelWtXhO0Le/JlDZAO7qCMrZ43O6Hf+PjqchX+UBLRHMyoXFzR32h9wT17l
fDKe9qmOsGXi2uoVr9P+D8WF9fS9CL+SOuWsol4IzvD/Wv9Mo5wzWHqyUb5j
ixg6xFSWGNnAoBAc2lwq0KrDaSrZV8qQPjkuk2HXQ1msoplebw7OpjcbaahX
SLcOsqhJEljHFxOntbb8RQYY4Q4qS8Pl0OGLLAjfAHljRNkvsedsrtgniV1k
FyMV7gRJ9nl6MJffPDFNl3k2n/AZkJ9UJpcrbkZazD9MOU4b0QTQ9Ejk9elq
Tytbbqcn9T+odMLssxHD3atcBq4a7lSPQ/nVFxciBKlGG1L77uFQ0hk0qCai
fVRFytn7iPrsEhcppwDW7YpPIqPvcooI4v1SFqYdLRXLfGW83hGJfmNytTvd
G2mMruh0a9L5338r7uK0Od14nTYQxhhH28BQsVDAFq3KUIztpaGONNL+Vm/N
xCoSLvLExCHpLy0QNq5Z7/E+EOulgspfD2Feh1LV2mF4wIcmDzpb9QEiixI9
kyXV1Swk9FjSO3jDZNlI+WXXIGO5bJ4N3eKSicH7unX8sEDAB4QKbAUdiQeP
NG6oZU6ezC7PB6mEi8EfBQCJvz2OzbNdBdtwCkugaooPbJLCZfKRWSB0YvCq
XeBr/RnzMTZBFWVW+iqywAtQAda/PuydcBCcuRpu6BXbYqSOLnIZgf4NX8yJ
Qs7jymsLnPcSYk4aqhT9Jc68mGL+ChyDTG1NJ9CsSTG/VcQw5J8fO934gJc1
s1HCp8WtfOdSP+/5lEwMQwQTQOPywzc2BL/75kPcwZlZHVu9M+rFxsF0YChc
f1PJ/0Nje3mrhtlGG7FssYLPo4WXYbNn8Y9vjPztUOpd1daGMxyxFoRrbXVF
lOvkUa0cq+s02qaPdI3P1Ff+EvXtGp6Svq8DesNkToLyy7w1CAbd+iClUrcz
1T5AWvphv2LpJuqje+lGsFMDjFGvlt4hx2Jm9c4OMmfaCWExYQn9jD0KM04q
tFUsx9/Y/ivr0Vna22LMp6gQ0JDBZ+B/w8jvVABzVeJSFheD80qhe8gSSt9N
ZVK7WUfNge+yCAc7s9pJa+msXo+oXqr07Oh/E7ZpZzyxY8nYL3l0MHbAVg6U
epRoGomN5mX8j3Z+tghUjx2YyXVuKx12yrBfPNBVQUdjhY7/9jj0MlYamTpu
571EOwwa81a0HI1N2sEYD5GvQWksQd0NtbLtDVvLp1WEuDcwr3iyfGQCQx+H
UTBrAKwf0kYaAAbA3YeGa1zISGNCZRObSoJsfQH61PrdEsOvlQgTf8DqstsX
X6iow2Wm+IIROStTK/NHVtMfL8BWSAjK3izyL6LbxGtHR3l6ZbhkZDgIQiny
l2tUdFfiy2JuohCfcItla8oFQF0DylfzPZiTuSq1N/dYGrQQzWmtZGdjt0tL
nOj1bljiNOKc+hUo90miqe6VDzMtrwuVP9h3fz68lyNBO4WhC22XQZVj9C13
NL9PQXU++7MvWtIyhb26x527P707h9E0THbDlkqHGh9/YkISjym4At6MEFnd
LP+E3pr4/rxGWdjSA7lkqe0fkNNHcE8HRPXDk4fAJzY3boae0An0zoDAc89I
n5baX4gN6clhPRGm8CB+EUAuaEaWK3YB9mGzpFN/rrXvJdX8XVxrC0dM1m6I
X7uCksmzkimnaB6CJqTZdroEDGpDI+W+9eVOKp/4q997fJhnzlAH4fBHqGt4
u/oh3068TfChtaaRntQBfmSLJyjSJXjEhY4NS/POQRJ6vNBey7bjg7/dyIxe
jsw4U3hZYyTXswOt2K+bw5p79Hcsc3YZqpcowJ54KSAEp8Mm5LeoXikMv88/
j7G3E3YGUmg3GwQ5R82FcjqnvK6BwZ7m6mSZTLh2/u5PD3EbH0yovF1YjaAQ
YzzxASLfZXyPSE8Gpiks8p93Der9zLpUrLswYxlEeslvw1y1KV8apd91ZWON
bqlY4rjMmgESWIfblBo0Axh4YFZ4kCUkQZjUEYzcw4IgSJsPpwfeVN3YjZrR
oEtMdZHOSp+9uts19HIhwsols3r/ic9l/WLo/KdTbwsGF26XTiAbSnFHCt0t
swASMAZ8o0fSdZT54GPNbfVR4Qjl2WtKoquXSJnGixNyVVkIhbPdl47aTWoA
c1Sq0YYCvR1a6n2EUFG3dPnCBo3GtO7s88V+zYHajlWcooYrr8n2b85OBAv+
923KxkdGSVo8ZTyOjVtv58bWtYQI5TeViDkhh3E/kDb+otSQz2a/0A7jt4B1
YJN29mRDEPpDVX0t+o9t0mftq3SWRwmrlquvwI+I7hYcEMl1E8NquIMyougG
VNXhP5LmLxFTCujH//NBHN/RBek2zWRIGonaUiPlFGvlHePmQApoBw1ZxHSE
SvecBB+/JPTtb/U2AAyyVdt6kkxktjECcrFT0uTg37QxSKGajRapFDri3S0N
BirTYcqojXVBOQTQlYrdxdtpfutSHubV12KT6o+oxDbWNAmDJvccPTKeOHCB
b6SpYfeI5l3jJ6rnrPWcxD4W2D8jUqM3kYOmEu/kDyGf/Dnb7j2ptmxKV9QP
Jun73z90rjnp0BEATbig1mbcM8kR5BergRwPnKj+IWFFu/srMI607kCQbFRE
LnP5F5LYumTgjBz2Z3R9yIIV3bUBSASQuFsE6dOzPYDhRnLyOeVrBqGz91aV
TWSWGX1kG6jiwqI6q6vfibDTGgjZxIrhKkcUAv5uOgjhUXFyGfrMm0Lms2Ja
mhqPepSWYCu1fe0XWTSxZ0N4To/ChkqDuWKqLPGUJ6Q1mfxAIBkIXQniJ95Q
EsGJx1vKWIsWdPq58RFDrmVPdAQhH7qT3w8UUtmbCOG5euw5DVDSW4tzBEfA
HPWaTO2Upzg7EPtdW0jfNzktoxwGvmVx7HtdosSg1kC5IW/UsUDUExUlsZ79
kBKusMj+YXzPZo4m5GeABT1onWIwRKyEMfPEPYVA1M9H6J8X2lGZZjmsLALM
RjGF117lVqoehuyOLFilUUIqPeTlX47dy6Kd/GzBANewe+liNPbgPI6jvVOJ
DvzzA8PILkA27Z4UdRgfWuANqNvXbcyIBRj8grKXcSU8Tpdh4x5DTf2sCYeT
6UCtXDVzi663fm7LFIm5aK7vv6M6JZUo629NkRFYEsMPLyOh07eQd06sE3Mm
puq+Myeo6GiFcnSSmBLYVn4SMWy1Zn4pEvQh6iGHZyPBNwPYT4uKcWqP5LgP
5euERCYOMlWmUs+3Uq1/N23AL933Eaa6cfTWUcItrkdQ2aK1/FfWC5y3fRqp
g3DuWvbyG3ej+xr+ukSPI7bKvT8kCcHhr91XBd8dK10+XZplkAJT8QaMwspJ
jIgPtY9C0FRFjtcEMkZLJ0jwGer5ztmZ+UN0Z73Jp1rUMBLGbOYNUxevb4NE
dKqwyhbEE83HUKvsr8OnWfSeAq64V+UZHQ9NQFCnoMmPowoZQ5imtHNWxD+M
N7uODmGJrODwPAH5iwxymqFFVbq6R4d4XSJagfAXc1OO2Q1LYAHnjR4ggIJ9
4jGelBWvNFfwxh4W3iwhxsaqKzaqcytH3CEhp5d7rakF83Pu5h68ilT5ANNI
YcY6UBayG6WP1iuUGL0oq8lT3tZMi5i797Ie1T+usKDMyYLzq7wD/mEQt4sI
P/D1kP0yTI6ifNDhFNWYwnvgjxz3XVlcP2UVHiIKIG5VpboPVXnxfEudBLt/
aMsRYTMKy9wnqxn749fHEQMHj3bt2yhXwtsnVrbAwEcU1ivTSltxuR0U+w1V
D7w1ftcHT9ZD6BqjUuOD/SrpdRSkspmekvF02FhGTIv8T5xYu6eXSXStn26l
/kRVACLRlDmqPw+D6T5dJo3qteCQVJfeid5zCc9KK3Q9Ro5vTEukuFSez7sh
5qv/EB2NcCgxn2XscOD39PO9OZg2ZMq9CtlAuhOtXXI2JCq2Q+fxT4E50l0T
YMYYBFoPo5JHHzolpyxc155yG9IiD3KpjJ5youOn0alXDlHIhZc/KhY4J+9k
H8iWZc3jyhPW2gv5tETGY6R+LHgOpE29S8dk8ecQkQFQoiHO6ixe3zmWAuwk
Ou34SXdtQBr2Ir5la9HqCTBBbV1ni3qEaipcdr4RSpiXOOSKiTUyMWlPH9sA
YBAv5nR9PoMPIUSBDD0UCBb1UUrWgWirWN48sWyl6XNBfIWVH19Wd3XybaQR
yC9cTLN+Y1Qj1TuT/AuKn9lHuQQEj1XzTXLIjfA9l6UqZ2jk7o7ZydbFwY2f
zIMYXdI183qPuw0jYbj3GJeE2grVhM7X7DLT7fmMvCHZVyaUZ/66KCZAqJAH
T2THzP+GNsEYFJQyUYqOxe4EAxdZFFifvSkIQDT7zQT3uFbfeK0YOpahK1xW
5bWjf+myhikpv5xyFWO8p0qicxRI00ERP/hI1XAVUn8y+eHi/ZMeAZTbr5Yu
P+IKO4vclqBO3Eonk4xTV3mHzSZXpLB8mFo7iMtaqEqzqro4Mgk1ua55yjc0
WRtEsyXxGZxas+TLCb3svslYUXknCF2b0rVxXIfPzWyC/0305JWSMdbKfKCY
B8tPAtRBtcIkewvC4n/RH+qpHwK+aw4DiSagcVM+z1qjjJ0Xzv1jbUwZBD2S
qWFoB5W27vcsaBkgJTbJf6XySvpVQqFc7UXzj80/WkzsHrR9iX2FgK/zklBB
v67wAYHpHZJca8t6DFs+6irQhQQaHjgMHa0zmM+sRopQHwGtJRofcCGWn3hh
V54zG/K1paK4BLOq0WZge5i9RnaY7muy9JRnrdYa1d1+hiYeyl1H+PWyKKGk
j5WGhZAuI8I18xHLAGaC/5IBbnmipAEe1N0AT79UCfXyJRT+6M9vR9fLMCvD
dUAZ9zgDfRLOZtSpTfEyADjZgxB385iMo0lAyXckMPcx/1/36nNgm8+/Xad0
yRjmMPvH/bELkUFWZVE9UVdg8t6c+YckvwtcN6NicJF7ccxQIC/lTECZl9p4
SbGuNYUGSDPQ2YrqRybp+babAcrqB0GxnrfrQRhj+pVexVVKYyuIscIUbd3P
WLh1kw8FDVHnxqwzTj88S7ae74zsTE/hsmuQiuTXTlgGA4lqfi6yhqdcTJtV
RpxXEoiqqnTmywaCfd3uzySRqs2NPfh52G00TCvEmX1h/BqqwKM20aCCVXAA
9jOt6AomjWWuzbwrQsamBsfjQo3bcavNqmCHCBgOHW/yWZfFPjijpQEBzrQq
bJEuKxJEk84FBJju4DbhIy5h+bsHvHgvOfxK+tAI+iCKloZ0f3P+Tp/vIOzR
ulSJh06NxuwlVUAtUDjpo5/2U5ixtKIOqxoHB+/L/nFKYSH93IEsFaSKe8pw
mZokH2aEgZpcCg0jXTqdL7eVQNuw4JC160hknxwhvlUygu/Nbr5Brh6coX0J
mHUvjOIgDE3n34oZn6e2DzypS56llZhMMdWDFzf5iZ5gFH7jxr5hGpT76Ig5
Y2Nb5N4YbuyOWkYUntnAM99z91bUrx32XoNsg3By6wQWJB1adGCYRYH06EkM
VljvHXjtOUHHYKQbNNcyyiYcV5UprgI/5uoQkFERD2vI/XL8Q7jT2WdcxUyi
CqOtmeAzggzd0zZuq24kPw6VCfEGDkjqxS/51xCU47nytuBhNLfQSYouJnVj
S9xAZC+qBuHtP4wFHG07DBGrmDhkxB3WQRv9XEpkjLOJs1pbtTlVgd4Ui6Iq
/9pYRST7z8DgYTisS86kP6jZagc5eC5VP0yH9cchFkkonuAUSQGJzBt88I4O
mq8QlNl8gwYytuYAjMN6+VdfVMHHIOln6nuJCbNIczIuvE2E64AUXkv+9lA1
76LBScp6EA0jvKrV9aKOorKd1oaDcb9r4ZJTXdaAygEEKUu6He1pV7Yizu5J
uqXoGU8pvc4T8dxVsXlJpTstju4mIAZSP1z1GHPqnNAPvo9AABNjbgFnGLXz
qnc17UBKR9TrYGiqiWm4Tp+xd5UrYQyu5boeTheSMQTEGnZT35vd+3Qp9+FV
Ac5T134lwWzWgF5kSMUZr1WyWfs4Dl7QkrqKIQX+4XBxTCVVb4xqSqVjSP7G
yt36up8UsJjiBIKjgz2tg/g5rPljU0PsvswFuX+YRnCYPpG1X2QxkhYQT+tz
hh5xN/w8KImPqFhsDUTQHdaA6xfdQThNEp/q77J+QutFZUXbbzTnv0nF9ghF
tAaqy3seKi0W3qaIcus1p3buF0j/tKyIAnLR4NPaR2+ecF/0JTPebswp1EUx
H5cU65Hai5dDFOUNmzj9VY+MymOxaSBxEVxhrp5tm04upQqcR0IKG+poYIyt
fJVLJrvQDiO4ZmEckuGU5eDYbMeRQV5Vw5KP/4ueRbwBhEo0iZ25Y1jU5Uk+
LYGiPSi5IoMT6dGFSqxNR5B1Z+r7ivuwACxIRyPdVTMF8BvtpNEQotnRnxMc
4dYxpAa616jLeNlLYf2f381+VOkJ1e55jCahUNs9aaZTVSE5zIqjo8dwr/lH
fFyVaM8xDGkL8sDju6/DJH2UHA499ylOiHltvDDi/Yg3FAL9fn6wDg133Wqp
3UUH3hfihMfL/CFYaeqwveQjiwAK14y1IjlPpKxZyWX3BkxuljWv/ZWsPmp8
Rr2JJubtBx9yhS7E3iUiaq7dj9Ox4ljkRQVpPBm0F4zLELX3P6Ss5Zb9LvzU
V9ppnuck5YSRDOk3Vz7pro6Q71ZRci2qQ4lm8wM473fytFR6hyY1kU0F98N+
wdeaHRiJc1fy/x3N96XHMXpxqMUI67pi6ZxCSm4+q8eobXsbpNdJFK/UhjFU
wIO71xPPtgI4vaRqVVEpGJOGfK1r2H2FqsFFziI8Aqf1LhU8az9imZRln6Rs
N5vozuPmCpkyBr2DtF3ob09JLdLxUrDoqtawCLAeX6OG/UJbBvE1EY2fgXrc
ebAdT6i86dNDnC3WtvG/w8qcG1Bvf8nHcqKWwCTqvWzSxfZbofJaOALxfRWl
Yg7fsHxK9vjqAZGYwzb2t7M/bZgIAH6hDrqhBMG5A4Jtw1rlHFVqyMEbedm9
RM5p6/fgvx3bmMKUiBYiwy1PqBKJC3UrzsrdEIkmkO/3bZW+MWj/cNzbwtfx
91YetCQYPpqUiGetyUO5zS9pjwik8yND8/1rU90sdxK7u+/eJG9ayUaNPKFZ
HaBbzp2vAVAlN+X6j87tEksC802R15FdMnUipA8G8BUhVhcltTw4eqjyIIK3
GHAyExR9W4YA4r3jduSPvXsA82SBZzV3I9/5OZjzjwcTiSnZBSz9oYZFDav9
B5VGjp7bT1vocdjLhMWcQ9zmL35AIcOfU9xg3F21O8oSTHypPjG7yp51mwiw
o+KHDPUSApV7Ica5k4vY+TnzBc+hNlE0e2AdMm7cyBxddD7MECTAewldeZLS
T+4CYrHL5EDaO4WZ40OQTiBdWNnKyFrnflxsUOrliir6aTHTTF/1IV3bAhJ5
A8KUBeeFjhEGTy/zx1D/05pcEGUT/bk1pDz8/9dwVqwrjKFb25XQwZBbvTOz
W1AM6Y70MohdsUnZo3xzxLsb7UUIT209RPrGAX8ScVjfCdu9Y87fYO2nwKI3
1xfUwPFnn5aFt83+D7MJ1//Nb7L4ffIHK9T92CRfL1WRih2XDFylmRWe3s+w
vlw6UY/LAlwO35N2mtJTJMWcsWhFgxQ6D2kQ1JRQq9XeY3uyhyoOgDGC/9wr
iRoK90TCSXJkcIE0kVNhozzGo3eBuos+Q48iBWlQ13oKkPhCmpUOwJuQMy7J
SABZ6pG8uAabSkqGoonAGWux7x4tfDP9L71xcME/lcy7FuhwQmN4UctfNzgx
WUmK2k2bd86ijaXxygxj9khnfvArPs6hf8y0hPLyTlsLI4bE1oUv3HN1lYoh
2lynUdF+HDjDeJklkeUsmNMwdAP80Eo4r647RmdWprTppntnqlaBYhHRLW9F
GNRJ0N7qJrfqc4iuc1XQNtEKIUypurnAzxMDTU/9//4RiDukBQGb2A6Z6i6I
qMIhUvY1FlbSeT0sxIh5YBTi/VyfDAsnD41jw5RzZR4nJVitUfnoRxNrDYAd
J3JJZPxOt7O0onj5aIPlM9ZrunY7HDyFtGywvo07R9P6/497m4+do0h5tSVb
XXta/8Okg5EJcLX3ztJLsALDtzGqvANLbZgFJFK9Q3PeXftZmy76p6FiPQ1/
OvoC2g15gIaqVwKcQOqGtGTUhUETXvMJ9nKBBNR2e+zFcThyMh2Sc+Pctlzh
xJkiPOAgTTrZGMAJ2r05ihlB7TY6/+JWONnk71DGAeVmPEucb758lYHP4BYD
td3b29DBWaipq7UhWZezu01J8vkSpN+Zl/9WUJnhr0kJvd5SajaY72pfISqM
dTsT33CU83HJTEuvCeso+nYF71JV3unouH4KjKCQo7EjjOn6rL5xuwQcVc21
RFrKLDGRj4GpBgQkrcmuw0dQOgLLj3AFRWzV9hhwQ9ZP4E4sWC0PwwTRXtO3
FMJY8RE2CGh1a0BaDkccG/e93OEmvD4pr+R7ZVcYq6HmRdwOuQbAatFyZX50
7jmVrUDyXjD26oR4rpnbQvw3E6UjZK+gLGB3dkmFVKV2qaT3sWrqNkXSedU7
Xi2gDn8ZK+wLg0B8PZ8KFJI9HrW3GtmM18WHbCe7Aa6Gss+8+y9BISMxMNHl
kFHwOIBJo/L4QnBEHcewAMPrKAUcsa+q7SuFiwrPOjQOL4zSuoi+S9Xb3EMQ
bXtkLEsRf/wn/NlKYWp8Hcw6GoITcujxck07bahfQOYHzaLgUYMh8nC5md/Y
xExgx8JhFms5v1rVaKQtPo+btzBWEa26FbuWDNX02MEI3EgpkWVToBSpC0rr
fK/dT9zsAxkQIUmkQd9eFFN4CnpN/v/tS+BwG+Al1e4WTwbcif1S8kOWVmOG
GFfRXepjjQSrw8egNb9vzMT1ZlH+Ufamf+BMX++TyrTy/fVcxCQgGP2rGXxT
vMdy12lGZjyN3Xfv0+oObqERxVyjoYd001Do2bS6Yd6ATOXEO1CgFhKZek+A
YOAfc73+RW7VEXu6qyigNhdnOlWBJAd2UUaTNK493wFk+jIRXQRCpYIzhvqr
nBTGuWsENO1gZX59HJ2ub9j6tNcdLqQUjE0ltvsKf/AnIlAB70a+wXdCVOAW
ZYeI2wwlEe4MS7NRMerj+zJiep4+3dQvDWrUELGHXDgekWTqc5sMCETjuFlT
Gno7pNuYu9F/POsiFcYnYiNEFpp4m2glj9i2ggcWCltngLJfggNpBBYVehn8
ssUxbBqjk9+j8s59H1PSGp/Cb35Grl39FE91pLKrO5RbMu9znsjkFZHgvnPF
f9pCy2KyUuDJUGabe65gNgLLmjjl+g0jYyXRLtSQ0+UGcMIGq5U53zBtmR3C
B7jUvMJNWswEQi/H7yT8WB+RYX3vDRSaQJOaJEGZ48bDhdLKO6ww67ap8gAn
XoT92bsJIcrHCAbrcp25E2fTKHjMuj8+yyTifYaLKN9p2yfyicls7HCFGM9L
nu6EBkuAObDj1xLC76IgIWP5+riQN/WY+GkExXlmHNmx9G9mec9SkKHEcTdm
VxQJ3cUUBKRQRlJiVf6KvscxJswpdafWwTzD3SEtA87wcu6omKqE/Li+Q4qA
NRpyNYiJ4l3C6qJuLDQJLqcujvNChpXOUyrTcHtoQlMF8xbYFOPcLLVcmO22
iAjcpqMrn+u4XcCtEptokGItEQKOD/5NPdcPz2S/A4+i/4iYTTUbg9VIuE7M
RJUHlmHKjWYOsRHM77IVBsg9ZA+O84udy18fGU4HKAP6BioondE/wdpQYyUa
mWl6DDq5oQhC4OQx+IFjERPcYNgTVN3YOcHYXyxLTMdJZ3i5bYzvfPq/z3o2
gDSy/lsL12PHWZnbQWr5zKU1wVdmzqfoBjXqThwBs6hBlF72TE03NsdgQTkl
+grLyqJUOrzyx48Xyg/8VzMMwkntGIk1AyC32EHAMIq/YE2gFCPk4yYnydRN
eBSKaSmXaKNU4kWDT06Z/+BAGDTe/sjdtdXSduN6hylkpp1JcNBE3Cq7Fnkd
1r+JNt3hM7wzvEIUfR6zXT5xjjZ0fE6Z7wcUeZjXPkk99G5dCkQ2i+lW4w6r
uEVC/4+pyL5cx2Rsmolzjoj1Tyg3Z96bEaSJ1TwcBv4AgXXsbSSxGAuzDCx2
0s3JOvKrYwpdHlVAYO43X5mfpoqneBv2mF77w+11T53xCLNHyL4lzhibGpY+
B/wWMkbZewrTbLbkuSVp6iYSfL8WpHEBYKHpbSxo/m3wDBypE/F+AgPVq0RY
fYNg3RgT5VVfofw69geYD1BCsVS87IPekYEWECFKKR4ulb4VH8sbFulKOYdw
DHBKmMH2ZgKOdK7fSxfL+s+S5CZlkctkZVkHvk3l/PxdE45zlKDRpPx2kGx6
76b5MlXUbtBO6pv6rOmxRxq+CoJWoNH2DRx4Cj/xjK322iu2fNFsmVx0mR0W
0kpyk7gKgQDbB3XPvlZ58JE14geJwPSyXFimsGRMw8kYIs/BDRU5Y5uzmZ34
Kbz7bUhxnb0Im95WLlOCTXe0wGrX+QhXpwY8toQDvEXAxIyHwuIb/JoF6Bg+
Y+0pXmHOwQaewRfHsISiS9q20ARHIao/xkqH1B3beX5EhYY8dvtLH7wSFp4i
KOG84PyKjkArvLcYSAsn3aEu6MPp2Ruf67HvPzTx+DiH4xnCu8/fDsQN4C5T
2WaFYlSKD7Xkwb9/RmIrqacMxDWQKtaiTp1JIvdCeiUFjn7Lu1suTaJQfasx
zrkR6ms+WC3xYjwWr310psuDQsWGz2v7vw7utSpN8nv0TIFeG92tUQEpayMN
hUqGXG7gu8LFfoUmWv/+67iekCVPe6B68ygTWMYFIMXAf7DwD1DEcruDaoSm
iAzEtAq1z2YSNUd4h9Hqfx/nltKeevBUUywKlMILLAvoqC2ZxhOl+3Bl7ryt
9FH7Tv6SO3WP9Gf1fApFLuGTJklWJMLP2nopR7vJ/ozqcQ/vmTGTeE4MmgXi
cLgY1ErZaP6cTuFSqt8/YlS965FWlr+SHMsiIXrubnYkW1eVDnWnAPsnx1Xp
QeLBYeXkWs5+7LGtKOjsYcNs6AKAE6ef6TPe/6RNntDWYTnb3AfSSghjrYhC
o2Tnm8rQExqBXoh2V1aWhh8+WznW30Ifmv3vSrVs3K3+mDksadd62lfXAMIX
9RGvEMLgaHzhfkW4PXHY4NzCuRYZDHZtfwJrKvQGLoeqqp27norm4PmV2cfA
zrqLjUf5I79TInxh/xKqz29TZiz4iuZsFEzvuabxzoNsKE95/W5YjnIhd8Vw
dhM7vftqaaTQOADJAdopYJqq5TZdOYScd/H+jKGyu6QGKvcKXTUfF8EXZ0wf
KgxKkXFqLbGswxt/YEK5OLuoCOkR0z5gRY8MQOf0mAe9Qg3zD/r7fEon3+76
dD65hJukk6FE7+NAexHG6Csrjnc7B5+p2KQWwHL0NgyWA35/KrFIArOb2a38
n33osy8upemmGUorRpxj6fjzaH9JGjMGTX1XtHPTJy3Hxs7rAQxq4GeLBKCM
TEjWmDG1eFJj/LC5xFO56P/FhR9FQ4OF8zmmrIBXZnhA1eMYn2PjYjTD0bAs
32Rg0CMDURj48t9VrSJ8RmwnlWoKcEYD422aHMV/XbsrguP66aefDwzW+GOo
scrn1S38Am65iRBZrBz3kqsmn3dFwkzZx59YongMkG4pAw8UgE3Bv6F1LUH5
VvcAzQQadOzCKoHfdt6fyjQ6eAdungDx3slWPuRhAU8c51uXI6yM5m+sufQh
RzkQ09h4vIo00RXM/fr+R/D/A0nNX55Lff4KnkzdetXefm1rmQIgBWTyWs2O
KYBPVxo1V0KddqdvM/ldvDKjZHwE8ZrIlSoMTQItAk1QLEMKXbTbjJE+hrrD
JA59UMUKJA6pOwwcTTvwK7ywns8Riqp89ytZqlZ7CNQ9oO2jLMhhk/R1ajtS
LboLlmpxrnwh76xHpV9Syv3R7GDlPk0fHUGW6bwuHa6D1yvndeBwDgGjTCzp
TBlm5PO0TkEmcbAWqMagZsHgIPnd1KlGxwbYcY3fBWN2/GwdHotRVGynMVwC
T8mYvm+wd5uDd2iUWN7cmKTKZPxSgfi9iaJMwl0pvXds4oRSaJ0061f63fwT
T/Lo9FQHfVrhCHEL20TBmQcX5o/2CLJyRyYdKhv5yDUOeUyQT3x5vHvvuw6H
XlRnAwICm9kc4rZP+vC+GKjHypjFtjHH49PqwYpYnXu/u0IgOQpTxGX8iF7Y
GcCejL4TgAi77AwGyDRWrINxKWCaXC6t+l0TVTcuM6AoA2scUYD2YYt9U8e6
Fh5ENY1oslFA44JZLL+ycH8Mi2+Z3h1FvecZQrzO2xOo8HWdKZ57P4NKtIiU
hlqDHoX9DahcsyIBgc6vAZaS8TeM2REMRGP1C/vzusnIycVuCy6Jyeu4s22o
mtT5DY/nXa1q1TNNRhENpNZTPga+o2kvsPcNNNNOghHLpuVYoUFg0UVwnrJn
IHG0yfD6WA6I6Nzk9BeUEfhjgdfX9ErAqJuHf72Yqn6DsB/q4fO77VWKbe4V
HmlhbKcZoA7oUSWfW+90VuQkIYVtq8M6pMoYZ2stDgJsXmSbdfZXar4Jngk6
SHEZZoRC+49Vobi9gZSg2uWHxYLKX6+XcEg2LVR0m2wGbyEMPRbkhR9mTZfU
087vvFEqCcSG6mz66cOxvEyklt2BAPuvGhKYe2v4oCIjgTLL630f98bM0KBQ
gAvKM5EY8jiq9SiyMyFdsTSHxRjL/jhCMxtIfuALdQJ1xUNnYwpq9LT8Op74
IpgP5uPRbDtMKFVSy0uOEI45rwcSEBFDa2Y8KsEEtvp3BX+QI68NMRm48AdD
DMTB4m2YDPIXGuuUVeziCe+hXKiLs4hMkKbWzUehIIw9JZj8EoSygTrvUo1E
LjdCXwswwe0QSAi181snz6XN6pz7mhc29c+l3d2unLAbUNKo/VX++VP7SHvu
ilv0neji2BT+VoOsFzBjMwje2aj2sdct/tzDGppn2nj83WLTQb1imhiswXFA
7vm7ADyqcho2uaOkmd/PtKE1JKjqglFa5x/ef/cU+wSN02xqB8SYW4N/UhIG
VLRkIb/MNGo+OXOjO4w1MxZwnZqNV1rXOL59liFE1WxqzNL91eAFjGM0ACyN
xUy2xKSxz5rwBkDob4D6cAR4TPZgyMfy1wJ/lR3tPp3gccPNyv4Ze5xAfIxj
9LrIkpAyXp484s5Zi5n3VlQabfEorWA2O3Wm5321PtVkpxQoTW0f53Nh4LcL
UaNpqgB40vLz2w5wo3FjJ/nWO88cnzBVgYJMH1RH5u4Z69XG79KyFuQ6tMzg
3Yabuyqf9BAfAlXmRscHoxkDhISNhCQR/jE0n4oWMPTO5SpX9PsU0EHiW7hL
YRMf5AwiSBa6yqhWZMtwPFEUJnNJgqVIzoqLX+EvqyUewDq026uWLKFcU5JX
u1OaAeQHuBokIZBHRdJr4MzvpFEYWoQwSi6k+Fz3DoiFto5vkqzu+wPOFDF/
N/QtdOFbycFCzteoMatS8lpFrtf1zXvWAvqKQHSB9l1pcNSJw0OGBdObz//s
8rQ45jWHRV/H7INgQel97+foiie+UczXxPWAsd+4hlyMihQS0D5rXnZB55u1
t06kEl1jvUpHEHYl3mbezgKKlLdUshJTC53eCQ3y4m1a/EDVNDj3xhkvm17l
E8wnbZcoxbHv+JHOped+qQf2IH2ksqZEQz9R0Ft4roQSbzYf2fyCTH/cX3/V
7d2c+fll3IqopiNP31UO9YUcAQlMAKFW/lSUeGzfEjiDWqMXzkyImmRe05Os
ieeWqznrhz9GG7CIGVrmAVYOaskQRJe17OnwZUb7jnExTu7lQVvrvqmme0z8
EsHNzqghmuMgXaRGsJiSkeYXTpMaphhMeQNnwApMf5odfQov7wG8MX6UK/r8
lpvuSqffEuzmmtGahZpJVfNML+tKt+TKjYsH7LjPPwZ0hA/8kTNlNWDGwIjF
t/ZPPMdNxfotmNReejdc6kdJOkWb/DpQjlmGSzq5aDWasAJqFed4wF1UhhJM
aN42DZv6A8RCu3w1L//9oNX2tSHAynrk4ahTwJEWBaR33ZpGHJC4GHlBqCAT
TZukrPqgjnN5Oe5iucWbDN8LqxtAGx0RJcLYjci9rjN8gtEt2BrARhmZblD7
6wrc+firbVYE+K3G2xar18EATFTz1Rb/f2yk2WmBMP3YMHEk8n41/d1VOT56
Nq5z1fRtSaqsKT4fJmF4oOIR/Ad530MDi17DSrzkhp+NZSF/B5lKZebPsbQZ
/qjEJ2c1Iluzr7qbZneYErKs6s6+QvIXfnwVatkM4JINJgpXFI496592xviV
2jcMEW51ji7HnUE4BmamJiaRZBCiM92Q9EePF66bxWXcrr7sv6j70rarRNjB
70T5CBO3Gv7aNB75+g9jo+vO0CwBtqmkrG0XZKTUuH4pECT3xB/rqODD1EWe
9STrV2CbMX0oH++VHZb6E9iyO2PFjbDRyjmVwDHCKGdjo/oWEg0+cianujZ6
HKfAM3tze5te8IKWLYtH4koUqVnViu+WixsvNfoaMPNf9d/Imh+AWBAoqaw3
UdaiwCVUTDahCd3pypEakMjkQ62mNJWiq52ccoq6lMITh8JMqYKk50xNXFTA
lXznZha/OH+5fZ3IMHzblT8JqaC6LOfYGmT9SQV7MWqABQMwk9wv4aJp1Si8
kG6M4X2QEHsO8HpN3Zlk0e8lIO17JeXLV6EaoO4vEhMmCYPb6ak4YUM9C5IA
GgCIv/e+X+XW+Z3JOc3r8ScoFg7Nk4joB5myjAHmxYm1IBQueJ0eeSbkOU46
Qxktsjp5rv7YqXJfshj885Ad1lkaXIe7xHK0p1XBjC3wkWOjxpDNviNHlLR2
qvFKxVcbszcfyOOuT2vOwmBHh0UXrRk2dWMoo9htQbp2wbCX8rXFojE9x5pE
2E6R77NhbwR3eNBxMhNn3TjKjY005Tj2HJFV4mMFqmcXlzvZ79qU9BQgCp7d
oGXnCSyLoMZTBey3PvFMv7fGThA50exlG4OYXEbx4A4w4Ze0tg85R0ZMslKO
dcvvmOiaI2GAGSiEsl/in/Cw2uGIZbH/qpAxyrRtJeYBoM7K9NzEgIYkVLs8
wLgf7kVBa9yRQ6CnmKSjWonjKWUFxyTicmUK9+PcLkL7oLxo3gp4hOxvrPlS
Xx8jw84/AkEyyK2SRlGnJrCZBgcynSc4yqPwjRkmx9+NMrXa2FY/z0n4Vu5p
iUqGPfbwdJxstVysarnIMUT/PKvmX0UDleKoW1Uw3ymjyLxEmjxOj3N2wSB4
C6N8bZhdnRG5PwIMe7tj3Shp9EI7BFH+/ovKHM5PUdMJpBqy5aOqg3ElojSc
4tyh09TxYFM4gmYTqAJpS3To1CZ05brtCwEyK8qZHpeEiPlo4/+9xOFMPRZq
y3S/P0c6KedhzYaOx8wHQrWyZ7K1FWQOl0zSGMtZEUm7tUOMof5bmAmu27tY
ywJ+jxwwWgx4m57kTj/c5afZhIRPRDGRrzGWhNeTl9vNKn2jpvvf8GEIAhvz
+oT+s43+NRfAB7abNIHozHPNOaC21g5CvMuq60iQNs6VK8TejAMu4XGClIzw
LJPZWFP6L6b/vTYtTWqNYDRTPzWQryVvLT+tCauaFW5zxucn1c+CiBjkgtrc
q9UXcy2T7RJIB4erEwq7cfsV04zjTm/zsrQ8Ia6M4UkobXZqncVacEpKPo6L
/8Fs7POYqE/wwKpbfzL2b7bgW0fM/VdS2HAAlrEzLJ38jw41OgaXl/mhD4k7
MtQxlmH96WwU4I5X983q7d3CKK4HURtgrTDS5v84CSxiwUIyjaHCPeJ+Ow61
kIP07xkZop6YVxnfLYJX7JQnFySZSYSCvwt9pxPKjsBsM/pcZdfs765IeJmP
EQ3FJ/gNdX3etUVLNWNJsncdwsA+eajqRSv7kfvmFjPJ6FUx6/9q1YqprM/T
TsvL2bBQ5tEk0qlSHDME7i/nhJ6xNJBzlRl3ITQy4dzNxBFczbUUEHpa/4R+
4e09hpvTHpSJ4WVr+Ax/a4UNNDWb6tcvTjkC//ofUn3YJIZ/kLMtxF0UdqwB
ThZfLSNK7rWuP1cAvAg3qAVoYVO0SHWb7pH8hCeUHdifEBdUcujeDiD2VDbe
b81QTsyehsceKkN7WldZe1KWBXqew4sNoM1xqsQPGpJYP6/6bfcuosW7qMQZ
UtcBSxUX6+Z91MqVVklMaXtYHsx6fSQJI6rcrx3YFzaHTIdP01IxB2dWp6Ks
m6tCD5v1ab5YV+BiWcquGZvXPd9y6PbJ6EJjMpag7Hs/dT7aSTm6Xv8/4Dmn
h983rSvInAxknaoK890db6gFAffJxBGz2BhSoO7HHbiA2+qPTzlr3Q8dohKX
5fYJc64RaL1iz5n7Sb4kt1C3uHj7CICYOergAxkJb56xLJJ0JfZkPXVyGGJv
K5l9MRtkO6IlqUVCz5XBCNaGxe09LVCJawkrIHWXQOYOjReT7s21MEiXeQmA
ScFWdSIbzNACFHlgdjTOt+HmzvLpDfdp3x+7Rv9sRnkmO+RP4e+uQ7SCKttm
tagJhawuHuyXUowmVU6jlFgZzo9bYhKi3fTKrJK0wsJcp0VaYYvdM4kbUV+Y
AN4YkHcV0dpr9UBKsZk9wuFKavJ4TnRjtKELWA5RdhrCtpHPAtwQgMlXpd6p
dmQKz+NHGbFkCfZrvfLLTigqUtrE+gBNJi5do3VTKqvTxeSjQqBjQRTne2rC
8ILt/EdkXf3VPle6sugIOy062oit8kWTgl11sb2LJ5qKxwoD35VNPr4aazxe
4vQ6TY3gJUKMlZ4xGPiye0ryCYuSjegykrF23pLDjKc6Cg+eHErOR77uRnv3
X2/tzK3U69noRUQBbEnUb7v3+386djiybLU0msy4w0lPXnobo8szR25BFzq3
leHXmQkhYPemcROKCDvFlDKNsaIgmqk3+i3+JCYLSpOTXe/4XHEkr/Fzgg7b
jGzsmlUnnhvIowBKXCIvIgKRkbtIYRZ5mBG6veYYZkai8YweUlxCMmtePXz1
nJylttq94sBIysTfDZpvuFltiB5Xc5Yq7Hkyag43DVjdRwLOMqp7JCIg9kzC
RG/z0+u+Knw5WavK2t/9s4fW163hX1nnJTLjZviZOM/eqKFqnLCQq78rwbLF
JkKCMFxYEKJEamILplckKuISmIw82tjGnRszNcChKhYKRDDLtBKq8DEtT1vW
xCxBScPTx46Bb1AUvEewskwKewfSRTRKVaoA8CxTetO/e6Pq7HrhMYZW0+1j
T+M1pIK6RPjMSqB5rlBRKLe/dt7uqTtS9fgu33q+5pJ+nVk3rykeN/qpfW2Z
dS0ncohjXSCoI5q214t2fdSgSpg8gI12YzjbqlxyKKRpV8PXzQwPDCNiI79P
hAuWf5EtS9X41L+dm9J2v3lKZUNwuvkKvn5JJp53mIuunVTO/Qq5ALMXPMrO
Yy7sKJ2DYLRcWB2lnnhwb4f8XEaEpDeELIPXXiAN7NBMDV4/NLfRsfpAiBwL
ivPVGJXheHScIeVLw5NIRkQ9gkVQo6doF4zuF4rRih9P17FqcPeX2G7Je5MR
GvR2wC6HoXoUlDqg/bOV+hbcpfZZDOi5ufhHLbj29Y1l1RK1gXQ6kDCY9h3f
yiVoSd5pgLeHmxYZQnRLqU/ojIRagB5jLGxY7u5XAMlK9fT39wLjb23veCgM
1QWVjToteKvhb2zieFVgriVtM04CRFYhf8W+BQK1PZyDXFD2tqJbDl9BWQyp
KH5Lwy9u53Bg+MGvFmipp3GEDeRvta7sPFbbO1nYJp7oYOTlHVm4di0gbtB/
ASA1/zp5a48sxnIx2XzbxZWfx4PJQDNDDI+VSyiQCTffkDOJu0eyiAAKyi1a
YxDdDF9vrLWUgxbGqmaXGrpJm3vfOIAIqz7isYO+1jkg6OuFaCv6Yemej1cp
pF83JIU+4LZVx5Fh59NaYLmLKEd0zX2fxghPICYa2x0ahls+scjdbAoupNm8
Bvcf1sGcOUFVFbC35SSh1wMUDYnf/LZk4MSpk4Y8ojRcxXnzhppEUh9/FJJ+
opaDkeRiJnBTnxaSOfGBfy51dBiqI8GW4JgpggwfweMZLIVL6WGEAwPiM+p2
SoI8LcaAADRj4RWSGXg8boAIIRLAswl0f4snw6ACjIBorTEnQ8u99GWtGprl
7NCd2/xD3zTP6LUkUvdVGaBSEcPGKF3aZw8Hnonc97wXE0xWatshG4Rf5bnq
gYsT3OejEcSQzShNC0JBCXtBOJv0xtrOOW0TQNXGC3jMXJDFeiFmHcpcfEO+
YCi9l1q7aD2prcwi2BRYTJgL+8SGueZCxyS0fcl51Yg0fXRDevkmGmiKFmB1
lhpkAehVzP9SBBfv3d3GhHUL08pmOWBH+X0GZNXdzqDF7GLqIrKVwZBGNsiH
xdEs24VnCdek7YKOfx7d+gnRzeeV1TloReV1mGcDMms5mXv0znel6T5pO/KA
3M/Z+ewdgBdouIQkbUZeRcmDGuy8kdxF3ZODmM+8cXbMLgNFocMNrb8bjrTK
s5coMf4ncEDWpGiG7+bqT8j8B8fo/CD1rAemlzkotkmr8od5KjV1tK9akJ69
IJF2NUzFV6dD10bveFHkubcur4Tp8v1PSHbdqKqgHoOSVYu1ZaS8fM1lJCkZ
MXXEUyr0JdD8pQLwzL+E3sfvdvfEA092opX3e66tJOTzkVLODvpJBerk4YrF
Cn8LYDu8Z3zgtXActwtv7XymgHlIax6yg/r41AvsIOG7QGxSHcrjFu5/a/Wl
7iFJxzkVW6bVz04XbrW/++XKECcSoeuy+lzXh+kAnXArQt/dp5mYM58jz5+q
1QFYVEExni32kkCGvYi7GcPUTd3L2ZPcje9jBpmlJfCLzoJDQgCdM1bhbIXG
QaryOwbFM2fGj6Gq+FlLV05uJVmFRDHjaJOZ0TPyB4GyYxMcCclLMs4cX9k3
GpjB835Kfd+YpBcmadrnfqw+ym6l4Fta8oTTLkX5E64U5uEv8XaLzOIUe9M2
PSaZoDCXBVOwKPmMu7/4+i9BS0csH3hmLOs+8L35ngWHXHGUOFFveOkV96Iz
c5OPctMxvB+0QPBgACTviDX8b52jsjOL7MWOROTtGnfBL5HW4TSe5tDz5hlZ
U6UP7KJFablwhXPUiyRq29s0Ul+X+J3SfuQQAK+xeHfMlM9KmbxBNXzoIWZc
kqFaHfwLs2Aq0mjj8uy7TdG8583+AMnNlUcN12rYHn/uirA+Qntp3QOHAGOw
XAxThO8QAjKyiyNxk+Z/yjXG01jBpjX+9cNYSq2rWqcoEdVA8PCGH5V5ktQI
Y0QMlRY2F7mYDWhMIBkt6n4cxsmtkNt83PxkdltIEQefuyBVRYsMwFYP5DJg
i9i1G+tVdkJhbIsbS9QLW6+HcOG8Sj+7s7x6iHDFym7r3njKzHikqCqwuMx9
4Pd3SJBkEtLNow9M11oFrFPDE9IM7LmUpnp8XaqfLeF//GvLW9X2iOCXSCaX
vs+cOVBKTXr9nRclYkkIPXVfEYAZW+k1GLnqS/HTtkicjQigZ8Fhl9X2nekH
W69Y3op201oxnYPcqBZBAxIS3toHmoDOPHonlRu28YedQERnNXCOD7NQ7XzI
QzbFkjPY/N6B00fk24hhy9hR1YsN/EjOX5kAzK5u5LPmkFYHnNuJ5YgSC2dk
PhL6VfdrfFa5BPFe+q/bhxnTRfCvPKCpUuxVmEkpFPQEqA/fi9E0Mdiw+dsN
hPVjlqmtZpOFtyGAGFJmTW9P1OJiK4fB7pWn9j+VurQRcEQR4VZVu7ihTazm
I5mW6+mVz0RoczLzev9Bgb9vfLI/fnSiaGD6T8e4hTmhUYo/Gje3SbMzoJFD
qpbG6DJ5Gcbti0mnBaHwrFtTmWLPBV+3BSMpqEvPMEKTRrRG7jlCKoK4YlnX
henB/oBSTJg3vnuYLoJ6fQ8RoIyzJspfMcaiWx5RZZH7y6S8wnGSe/c/ANRx
7REPbhfABtfkkgRA2rFKXj/Qb0AChV6e+Ex6+bmNG1BhTju/7U8u/qDSk5PU
UmgBvsozHS7wBdDejGXIpIWArKkSgTM6UO4YwYjxPbCoNsEPturPfW7l5cQV
ZlaSN6/RiFaodw8r9+yHBQbEtu01cWK2QajmG5ca9hEPr04hhPrk9UjVGKeJ
UlJ23kuZDYguZ1BMl4yyTOtwTUOZwvNcIlyWIeM9xrNtt+TDFisF8dO/GEdl
EXvos9XdJ6b7LpPIiE/5bH9XC56xmvdyT7c7+GSfolXMM6krzeJ8Yhk9g+Ot
GZi13l4btHebh/ZMzx8RmBh1AQrHBZcDhFkOHbjHIBPWMsBNBAeT76zTrl9u
XSZTWEa93vnmwT496Cs//1LIcr8MWBBjKfZYgdidZYlSeUoHlNXQjUAoHdjp
OUBVZNup06z1eU2OQ/Pc6BviSBoIMlC4tfmMeaOOIHjrsMhW2btv+gXhx7So
abX14T+O7dD7iDFJ1l0TWbxyVpp0/cKeIcOi02pt95JAfHuouqyJaz4tx2Dx
RLpBtGI9Huybl4/l9wmEHiRBoL76DuXsep61x2lw/X2Krl9bLgDfYbCEttQI
oEHqQOtx3OGVOsgcj3GcQdSP8ESsKayas2SYSGkTkn3XiQfpFW2JHyDUV6Kw
M49jXQfCVuyLGZh0BctJjsw18EskuOtnW5U89+y2q+NTBVXM2U4TlWUvoFN1
J84SoVt/Z4lcXoA8woPgINK23EDI8FmXSyithvSmQ5weZ6xTSFHcC55lFaHe
gvQPb+3gQahaxI5McGNY3+TK/QXyYDiCcxhVBA/3knuo704BGlktXGXxQbjB
wVEIgthmwldh4EHOx4hZZOscZnqugtooWPZkVohCYqlz88xtIXlMaU2u/6LA
yqs59EoTfKz10/qvgArbtXfUGSm1leY1X7TYahz3Nm/ZeI7tWuIlnj3jKD70
7iEWkKtLAokouE2sH1CFxmAp9RgAoqMzm4nWrI4jkQP5NUlOUqkRQ30wzXlu
96btECB76J/gQwuoVpmpLYyTXUzcYfGCVxHtCSms0iIYjSzD/1k1vRo/GN5U
yLOnapimwHoxSNReyAfqfJqzustbWfgOv4VoxRTFzUphBoyA0Qixgv26dlz6
00hqxyY6SbEpahWQHcfk9U+PpGu0O8AnLMYoMlwP1+8rFNLOJjb63iQU9Nkc
ZKDQP3+GcOHCn9zcbpacyc58Cf0zVO/MbOkqNyDzdBW2LskoIloNCGxdUjhP
rL7d3CTSTF3snwvXoS88OvQ1MwDI9YZM2aDsZDdTiRrpAId2CyYa6RfY2z2l
EGj2yoruNDH55NaZ6t/jocUKUTeaDYZHLVApteM6OVI/KkjRrPGNwRA/w/U/
QghL4Xl97wqxIROVG8HPfyC/ZbShliW/2QCHDyqLBIPJ36SVQLxwBA03NMue
Ok0+8GXAgEgi2Yu4VqlMn3PjO97bM0w/lQQkQbzZMqxmvaDGtPthkBSbMvVm
1XXeFBcRCJ8qosXCCnYv9YscKfWd9JaJPlUP0wjbdrpsW36mHZizb1M5ZzhM
2bQeOdaQ+UYQdOx1YiHdjDgaCIhUfu5hhVBiGvPD+9hOMS0sZj0J3/Q01e02
27NO6zosXcD/pawZhxLF2W2vQG35vE5f6W16CFmo09WivYKGE1MNgl3G6X0/
NZ0NdLDwR/N/gjJJk9DYfwl6rBTWk0C77IPAvpp6H+jA/0p2P/dsdxltc/Jr
fRFb8WFdkbzMryGZzaCZTDlq6I9mf0l/XtaYQUPDEFhLldIe02Lc306CNh6T
OMwIvdSWLzw+5oWIWIsClOanuCmdvphEa2l+KVHTDnSgovsSqoEOLRuiy1+r
VqsalaUPDGYnauM9VjNle+IdMzxxJcCTTeuYg3C6wNRMOas18aSXkPB/f0ng
7s/CzjDXmiW2GGooVwudBFipgNft8Yj6NQ0UsSJBMlG/pOqJtBIVj7KUJW3Y
ISJT4Fefx91/opDYhD3i57J4ie0bBMf/K4UNaCNm3hTbu0ivogQtz28AP7XB
OyiW2HcbbSt1FCazzm32O2cr6EuaD0UxSWgmIDgtKf+E2hHi3WlDxKMbWAv9
xYBNPtHkoX7xAqwNMj+fERjwXy0PGYjHYvwA+UpPNUHJygNwGrX4Tz+qNl8s
iy8PNsr8ifRZUZEmDTkexu9AHUtKfgi0aC9I1OVsn4gzweGayoe5irPs4rMv
HOKmjHHHDHOQxKtCwx93ip31TLQ/C+DnA9p0O15bE0tlFG6dQ8Tg+Q7bjvCm
1BlHPyU3ZkmhsvEX/8CKADQrSQZmWWgj5IPvLEWEpfXz0PTYnKZhUjquQ7A8
fi9XRZLJZkl1cGOPVFIshOHzqK7PUNvOIQqqAD73u3uYmmaOUv53y2qOCwsg
9RAySOiHbv4uOxIX6Rze3PTtVkF3Ofz51D/Hb+uEqbqrVpCaKp1JS/1wEq8/
Tfh4MAT/95245Vm4evwoBufoGsJxtSaD6wOdWRP+v205VSo8zzTJYsVzV87t
DxgwLgi3TTJWVq0EufIlj+Aqkjrd28UC0vwuPlFiMTiCV/uZ9F4B2Ka64WtV
Lp3tfXPgCTUvIk6MV5JAO0kH1ZPRZnksE90Z4P7N3ka4Xd0lKb6bWkATuu+e
dlFkY04AndWPpTWdwNI3MbBsBLdfRmihO5/C405zVdZm7oXLtzqgV/8RPzuy
Tv3n1zDJy2edqCtcZVXgEfQB3brHhcRFfwAkujEviBS0ejwZpN737NDi84pM
M+mqSu9sMuc6fpM/heL9BrODsJBNW8kkwXM1vhdr246A7pyayYgbCqhpTxcB
xSxVYpvRtU7XTYXCPqsJbobzvF0I+vKiRujphnfr664pWQURiYdGtRf1rQQn
Rs7LsUMM9GxhJAgBukoKnnA9f7QovuMo525UxwrJShlShh3JXreLr6pzEtB7
Zuj5Eo/UfIHld+KMzC7Pah0y+bx26lYAkBr0uXVFpSFyyogW4q7avyQi3qaw
P8foSIY77i4H85T015KSHgyTllmhBngs2sKYgnUoQkzZsu0CAiUvNHc6utUW
mAAD8MNab5cZhCOY9hfFkgJyKiJ1T3TpayUFz0CWEGmYcsaG5x7IjoQREorr
BGJlxQi5tMUt5gZHkF60fYxLB/CzH/nsm/ym35ZgfL7FhvGemM5uapRNspUc
F9GCq4ptL7JD11Tvsd7wHdnH2k1Z8uDQC6QccOKp6yrp7Hc2L+GlGl0mgpzS
FKzWfYgOQP9sypbQew627fmQYZ8GMDAvcUgKWm+P2F7maXLK8e9gTGHwhiJK
BybB+jJyYcRVME5BWv6qryO8l+0gioKwAOanSd5r3cp7w1A9S+5Nf8wMf5o8
s523UOA7hUzgSd7bDQ5V3VBXqKWdEWm1gb/eQTDe2FD2MrXicowm9n9E4Yi2
98R8l2Yct9hp2qni/1310KisfJend015WWWfSMH4tS1MAf1zD1Zt7jBxx27U
4Xe8p/oIpfa2yofGklP+wYI1z0Sb5O7WWq0y9UWyyqLDk2HiIzbFBOa5cYl6
E+zwz+ZAf66LcpVf6QVSIMT98+cmtT/k/uPXFSiycv0ycNzQveU687qRyFvW
Zbb0xttteFFlzCUvq4JHGtlb4tNRL9+NMQDODhxdRtXnlc54FgcEFwlxdiSf
PNtUHW2bng4I3U/ehW1n/5NQsihg08x1IGSzg8+BsBZcd2FSVQc/mm0qY/0U
dCW9Jxh3iI28qnS0/W1lBUTCjkkm6NgtFEkdrfRJ6nbuFUHjhx53U0v16Nu1
aZeMmHDtxygslg6u+5UYG2jFP3BrgBJT3E2nRx5M+WQU7UlJj6MrrvWTqnIt
u0cYrmBInW2MzHGb9qYFBwPe+9dK2LKTxAym1Dkrer5Kt0V7WFhq9eo+HvpM
/LZwpvfaNsjsT/xoWLzHlkTebtKK+OqWgNB0cUYT7XFirpa0ax8H2wwybE1v
PNDi07V50NQWEI3veADHBDNDXIjiQ/vDzVGYG1c5Mb1w9B0Vlp6EsseMB927
hcw1ImNe26enFXX+bagg9y+NdJMC+GOK6lwb6eaga96DozlWT/VsXH/VSQAu
2NSPPuWphA7ibkgwGWw8AO+OK48BVTY25JpPvkpKeM5X6y3g1aid8Tvrzrut
ldyN3c7zJGnTSiWJOxVBKJfipEtdXu9TzFm7wHeVmAa/ED+MFC/xTf5H7ezr
X1ocr4FanSNYAFCJPNMyfGtjkg/j359uJ4CGK6k6P09Mqy4sA6qHevgPEJsv
ln44Cp55H4gAe0ScGrEJvYIA5hpqSsnknU10ir/fPvdO3ZPHUB+FrWl5XErs
UReMokWVkyRvH6BC9oS0JKs5OrflyfP4OVOf0N8/pdG3eFPUjQJ9piuqc3Et
MQy0q0oRT789GcAvTixu7t96YQTN1hiPJ7YGU5FVHKcX95FWZukJRUvvmkde
9k+2y+NsbPdAf5kPFcYlcfjxbgjU3b3e1Plge5Hx66x+meUE9upqM1DHN9tb
N4OyP2D1taeFiIljqloq39G7U4xtKvsWRAk+49jjRDAf724qOEggF4Px/Qhh
YkelPnTdePPfAVa9qIs22xnPZZ387h2bZW1JcfzlyztQfizasGjR+LcYXoZT
WUhqFQaOi5i1/+Nwba/3jPURespq8V4tDMmFwuWM3E0W4JAXP/pquC3IfDev
IB4hoaZ/SoNdvkkAAel0TrVA/QkbYaWeze17KQ/DZsKR4KhvUDMoHsHzT1ek
17pI4e1E3pGVac4VDzlU6JWfwzpc3yZ7FiuZzJwuJ+DzN0AChLiQdpHqg1IU
6LLg212QoKY1UGO3/Iivik7lGKeR/lF0LwSHw3y7wJNMAEDg5XGlSKQINJnQ
WsKn4NwC35zAu/w6UMBDifDRXRmSF/VBy6UjGqdePIvcfNbGEMcE5xCuZt02
RxKMkT5WITBk8KfOVvfrusrzKgMdF0r8PFPwHwNBJ1sn6AoFIDAYEoLoHGU8
OA2yZnaLn/rCbMre8t8u2KBq7APlgFNIJs79KthS/FPlDTGmBwB4USbIuVUq
pM17XBwNyiDtI47W1pOQmxO0V7wLtyTveygQHHiiLuWvP5JoXNtYtf0PxV/M
hPwgTQhtA7Pir5bo9Ni77JJZuR7oXCCzPRnQSER3mmPijvgWVL9MRJ6bszn1
7fma9UIr8T3PEXPMoK+E7ngJLGAiJhEaOb51XSR+baqpHpFGoHfICV9M3LMP
GfJrbmsg/8XtTFt0Da1KnYsZ+usWg3MmGHi9ug+S19f2p/3pDNH1wlR/y12E
ddk6HPDELm6hRnPr50a2NCH4SAQlWg1p89CUm66h9nCBdri7chrBaJq4EVmg
hsGGPd4GBosGQPgsB/gbt8JLGEXnrwriu5DAAYi41J+6vrcIA5HyDXQV+1hz
7TqudttrP21z2AFV4s9ZMaPahnUhlHDXOlNmb1aLfDKT0i85I33gJEds/+rX
czANqNQnC3YJSsZ8E97KR1sjblxTRouvb5TOItlx8znCaMlAB4SMTTQR7twS
eW08xciPEeb86XYgpdXRjGkszlh4SKlNwUgaM/c87zImSCjp3/rtUUH/xP5n
lvEIF7QktAIxxCVIYXHGJi522a4nhHfJzmu4Lq4YOax8L1ZBT2FwcSOgtCH7
flEHo+6YU7l3b+UT5s2tQBgpKNGV6h52DK9gKitqueriSK8xuhpOQUUCj+aM
ktY+dzbUx+z51TFCjgy7BsldIrRVYQ/nE5WMSkSGOuc2s9KeKkai3TUXnofI
LNmf14dCrSq8nuyU8rANyrbgvFttrm2Pvjmhcq7QJ1bU5W46jnWOlsYCTpFA
hP+x36A6KAWpKxeA002acrAzKBxmX8R0WWs/5WSJX2L3OSuAXTMm5dOX79gp
cBilr552GTJouMCrJ8S3D3P7dtWNaL0w8WTwsEkUZZW6ogDmkA5AF2RPsMOG
0lp2nQsGfXrbJyoNDbkwqAQqTU9FyObAZCyXirGEaDjSnSd4+ZSb7OBD3FFS
l5Cdvocl8vsqLJtF0u7jeXOHsjCI3TsM7F4X82gOAY1pt7+SbGDC1ZL6Zl+p
iO0tyENmQ/Nh/0iDqkAJOB9MietmDKMBHnY5SNvijaaamkao9vw4CbWk8z+V
365yRwSLsIOzxDudeuDhCbvvkDNVQqGZ2t9LIymkg4Q4IAEWo5QICfXG1ADD
yatOkHX3WrcZyuKcVXItM1Z0XqKpr5d53rHKzHxMZN//d5c5kAZcw/MIJT7c
DRulGRTRbVdvVJSYGPPe6drfADDGo3ZNpHuxKplF3Gkg2/pjpl76nRGZCkQN
OPxAZoIHZl1lT+7M6zCGp0ftxEVpjmGgSG9lJrc7YFOe6Hqam1errhca1fgH
FqsqcKEQPJrV+n/MdCSemgBTIQG1D6HoxwzEAByzX+eX82xIZrd5Ww1O8P1m
10i7DVJdoJL6bMb5K4zE1wjqvFq86JdnBLWZJcIPnZwgKPXdYuJDvj4Tc7Wb
ZAA8zjD0pTrlHAP5nPWG/Xtd+t46j6XMQJjaSyckTQWjxtZhlq30yco3H8HM
XLcSC4qKI/aQFV5cblyi5218cvESBfNHJVmg0SCOc7/yB2VZ4R2WHyMuI+qe
T9thcXYfRN+aFrzGZyx6DextKoDMPbp1IY0pdp37CLGTRgzX6FTCV8GYnulw
ZVP7O+lW4C+SJM9YXHqYoFUZHbytII8aVDLbzDdz+wp9Gw67s3JDMwYEcLGy
m3bwmxHRuOUjZglzgQCM6RJR69J7+j0p06qyU+BmaHWm3vNqa0AMJwh1Fp9d
vePGPESJQfeWl3tgs6mJZreKorCeWUc/gR7T/dSG/1LeRZLILbE6D7mLi1T2
PkuDxqDmhL/3zxQnhox3ZfCbR7skrVdYaI94Tiz0Fb6Lxp/EmNIob11W7jP9
KMiTSCp8JCKEOwNsUGFWP6cKZ3hrk2rA0JDLG4a2680+12694zt4H2bYav8Z
xgJ1m0kvkFOLCyn/4wE2qbB1y0rQqt3JDHA0NrT2oX5zf3ezrIKNxi2LACZ6
gEqBYfelQaCw0U/nrr/R9nxT2BaUdCU/Yt8pHoa4StTGaWWVPgV+uytv+9Qj
au7Hg/WiN0rbVKbtQQgYNG/9+oY+nltuuR6xk0oiFNI4hSemuNOguCz2lI1z
gg7DU7I0Fk31CmV6eU25Xv8lfsM2IjZnmkjRBsq9vt0Hmt+WHHQ4CZHuCmLs
FWKKcprLKhst+xRk+CBASi0u5MfompIokhlHkva66m7BQTiaEs0nWnPseeY3
aiTJ+4FWbmTeyc+lFtGoLVsfnBwc+5ACksxJzcuHgnbOdHQlLCHUy70nHckK
WGKBz/0c6YADVrr82B5YmeU8tTdfvTVtQmkd9DQpQfZK53H749RM9pmExmGc
SGzi7pHK6XJAFYc7x6EPSzM3bkOrN1rf+BstD0e15KbxgVOkvQaIEHnuHiUi
YDAIwjplN6ehRLeFkuCgU/hhWacSU6iKAsvaTd5P3YOJsp3hyS1Ph2ePhmxV
L8JWy5DFRqdPGwhkiKIaOql7Kx0r6bve4VCK9dJSnB1ilcw9Nay7dqUXl4oz
PvsSZCSzR092zvWaw9cM9lL6pJzV+0EPPpmBr0lEZAaSVstwBZOiRRMvVaMg
Ek8K9l0I2eKuwlOhvY+AlCC1/iSfq4sFHq+T6dL49EQoOLrsb57fM+WXYPRf
7ZxEvWDOnetCwRqjIEAtakJ/xwus1duXzj0GTjuLZGWhbizdDK/D8X1Y/rPd
Gv6lrG/bHc03xg1lpcVfzNN0Pxs8wMkhlRHiNWJyIWSgvfjXmmtp2fb/wrer
8ZZpMLYy75uhIjtcBkdFihJ+1wUn2jUneiXx96biNLgtQWOlZlav9DGMk61j
uXL0298UHRN3XNViCBnwEAhCyRXrMdOAY1C29s5OjiEgFJx0Srsk4g6WdUEE
OfyVfxhihaUj2NY3jK5HcAQcgUrySCCEtgpZRWpOpeEbbTrq84WuXkGm360v
vm8AoKpRRYY4WBWKV487NdcTaDz3aOiWqRBRnI6batl0UgZFXMXpVTlg8+ae
gg+sgi2eQIAmYNGI3VQKv2YAa1G8GCj1mgcNnpDu8xgvhRoKIae/2KkoEx8o
PdylGxhdV78ScjKkb2LhboMoNFIdGZImYknarFTRoOR9+eJqB3wUnF49a42Q
8ewjsRS+AjgFaspqDUigcIjhkfeRyh/wGxz3Gm3IUNKcntBM/jkAATr0FaCE
fLHh3V5dSIePJewTflUZ3prW82DG88teFVLbBsEdOIY1/TlU0+W/9bv8yya6
oFledFWEZ4q3rVfOPG+T/rIj2PKcW6qzZfz8aDYVVB0EKCjDE/BoNWKy3ZF6
fVKvNosIk/Sl+/IIr1kydeNUApPGhNfDrHHUYbSUzpNbz3Cl8IJxv8xxEvzX
oDN4Fv+9uAvRBkf3hYzmyIYjg4kCI60X68NRds78v3nHgFCgoDVQ7VpN20FK
+fBdT+pUqI9fV1WIz8J0Zq/LXJrwnDg8WhAV8H7ii60BwwGLE+aKzWvqnLDB
CS2ZhuHKoEprQpu9/geY23FEpXCyDOzHyhvTb/jNv4ObGvMH7xnBni0PGSYS
Bqx7Z8+QvsSfS/g+f49M5LN6UjVOhsU1Vot1higxWhlMq5Wnv8ZMAlTruxsA
J6e8TX6mEeawzVy4txtqb8np8KbX1VOlS83h0AbC97J1LWjMy5+bknEIYG9w
EazF5rnjEUkY5DwBigKt0LxJiVSIwBkKURCvEgUXn1FRFauveIOBnciDXVQf
eH9WrAkRdIEtU6+rIR0KVO8p9sjE31pcI05i4ogqWZ9zY0HdzpQJ2JIK7t2V
2JGUGSf5hF+f6iU0mSo9uD/Rh+ZBAq8mTB+rCGI05lxFxVlR2RJLw7I4eFdY
0epzR7h6RdX98YWfNnulrL7GzGfDghSQCbn0ozZmjtmYFdwat98g1Q/Y3NC1
KMx9DTVAR4/HaMKks7l+oS+uwnakKMHaYCTtgWJTXHORcUNw6+vsemhJSbcR
h1KwwclJpLOid/C6gIdrGoKw9MDrexdfA5IB5IPd9W5+JAQq5XohG271E2o4
sBFltWX1YURhIWOCKtHhfykBCyITdD0XFDvT35BlhTb7Uw1W99SlWtI8Y6sY
HrmKOym8tAC3C/azz0QP3vmVXvnzqEw3Oq8azEKBjAkrahB2oJbrdcDQdssJ
xQ0k4N/rDzkx3zOMtXVsfkTulH0nmlB7QOGKqsOR49Qy+XApX/P98Q7ynzKg
Di84xFkv+sp+Xj2uNwoHOzVnoenv1/Z9K26+PzThktHcB+5CjBv1yl60bAeO
o2ck4ihAGGJ2F4EL1JUaql8PFyYiScU3kqD5r11N3+jw2kAomoUhN04yDvyf
R8FrtXHcA3PvX57dVcaTetQ+Yu/+4rW8p0xue8TujQprdFIeBDK8RNJQLnNR
Skd9hUaaHPJzROB5NBipM6WdJSNxBpgBCGgDlgECMkoxogtwNfsRPeCpMeVC
r35ULTfng3zqM1mdDC1mSQSVUTlp4L/OxYbC3UCg/zkyVh3lx/Rzy+FqIZD7
Qd5A+0tGNRAJF84o3iDvJYvgj0sUBxSUsRYUXik48sRA0+CiEfhgYKCDEQbx
eEgjbOO85W8+JeRiZyVPlkcj+cRAfJe49jSrdyJCE/P2ED4Zd9IUaaDoBdgS
2Nf1wafP7LGaQSaBuZuiv3jtOU3C7uaQvx784LFbV5Uw+M4Gz71FQE2Kxp8r
ctYDnv+mjDst3T87oLZ+UGsJsFnPD0AozGVKPJvP0GwJOD+y2LJyXsb9O3Lt
1Xy/bMwGWVSWZTt+BvyvOifbq15RVf8HiiD6EvEBVVbzhYNJ2FkxZDg4xsT+
shAIwqif0N2sB1g7Beihl0PQuuEkLF0r1AgAFfF1wb+FuZqQmzBElN8qyxrt
Pmf+CmxAokogcV5+wIMRmLMkPTkfTO14c/Y8I9JrK7i7lHpeeaxC2Mi1IUDQ
muvaqsqoufiOwSeEC7UQfVUot5EhXhitostACdPngozrmUB5FAKovceDyXSj
dGGx0WQO6espxUaWbwQAWKUd9ZMaSI9ns65uI36jWNW762AGH/sCWsDSpEWv
mFO6yH7lMczDr1IspJ+YZbPSfU89/1Co8r9YQvheIxJ6e+aZByKJUDQ9267y
NV1NJUeRvbV+D+wBM90EaIK2ttFS3c4PpCONc4RGyOApqKDt119kbmssaqXX
R4ZRCdhE7T2INXOmrPhKzC6mn3WjPnbDL6wCUlrQAiybNTlH6AyPTCLuC2Dj
uzur8loZYysn2nC2r7a8A4Il9Ec189D9jqLYZU/fwe067MN6XcvmwZD8Fm0v
d/QbNWp0d+EmcQTbhe3NPNqOK8upSXgpydAk9mL6LF3542ciPxkgYd5yiHNf
6s7D8Pu/e3VHg4OPIXi0QZMGLkCZhKQIdJ+TBX7+pgScnNhiHa9WeYm/GICD
uMDoyM3xOh0m3yPfTq35X2fPPt28zSzx5ANdDWyzuR9yfL62yrGTtoIaJwTT
vXN61kmQrb8hqWs5l7izkXtwc1pL0Z8bnmqjiHODNnb66PX7ePbnZAkwaji9
VhWDMCyKGwkmsSsCziAMy20SrTUg1Ko6czo1sagJi3LXgVFV0PCml9hpZBiT
VPdcdJ3nA4XJU4D3CZ/7AqGqsluA3YU2Smd3N8XuNkxRKIkTVu0vZ6PEQqtH
bA3cUXMJA+32AYNWCvqmV9PQ2mm1Kg7aIRD9iBhQHLM+0vZZsjFduieh1ddJ
UveONqhDGP3Qgqe92ow6YKwnkWXpz3VcxWvKrJgC1hVOcOwJ8qDxNblv3YuO
Xog/uQYrKAy+jhzmgLzgFSTJ9dp17fPDjZq77fe1kUJQfT4BbZmIrXvYOApg
YtJVWL/kd/vNLG+uqyysrv3B1FZhKYALsy3dI8a8YNSFTsVY2FnEm43MTjJY
i7y5+CbAZf/+GPKlZPHhWGofqspJ2KwMw3+t+diszLa90DknNgtZi9WJ5uEJ
U5er1ScCGpXQ6T4iZaaPdrLPl0peA0kTjyrRRgLwU0cl7dJTWZOZ3k/qudNN
hA3Rll/U0J0UZAAvuiikhRdVlEBXpushQ+JDyYYrHYjvgf0DlWQ3vZu03Pwv
v6QLcK6Cf97cbPWdquwV6XtmjJZOQju5vRu3yoHjIHDEXJweryRQAujiL4v+
Iqv/6ua2I5X54MHdytuVUx5tTp4pb+n7SWRuBVo/T35i4Yrz1Ei+SCyJMKSd
nQclOG5qDDz9OLAoIr+fA5QuqCkHY6idfq+zgiQ/kXsdnj2JPP+QcypPITuy
Ayn4qUyUJnNxmAPiTwVixenhO/amxr0sna0oYN7ZaOexyXKo89pzHzgNqYIi
R8eS/t1M+c7FWw4z+pwrYYmwov1mwQnswbzgQF9fLPKuFDbTSCEOLJ3aZy/P
A9yzyh+vlcyjAR4BJW3QQExdvr0FIk+L0Cxw0VyPvcMC/1IEgVpz0AaD6x5/
dbbss7kDh7ChWaItLRkxxwpbyelSDYiXulXOqDTAcgL+AfpvK6eNtSzR0MDE
HIihXrTE583+CmhGHCBa14giF49CYj8lzdMSo1VDoLewo4yrjwEmdzBZcYI4
CSr2wMsjXc0lMqejWqb1eU/KVz5C/iMlgVFzC4yasdK7jdNJcB4O76V5IN98
i7KEfTBbp6O/+fJoEjXTfNDPBD+XlsckCgOeg0VNUGUvIuVo/0DEiodsyTcp
kvfcb+8HbvjX0NCGAf3ejHsDSE5/TZFJCklna2x2uhYoGAtyGEsDbGkwqQio
qT9rMqX4MbD1nDdmcLy0xkjk80LSRVz1tBX82ylSwqJjp9To19H4uasJAZLq
UWd7ZXlDOsyc3lxnhCXa9p9ZBXJ3y+KnETzx+cj2uLSBrITAFtDDS0YJnC5s
DOw4Dr/tDijTZm9yHcTrsjpRUjMIPDf2V7hUpFjAPrF5ZmyWo50eIAUnDJ+P
Esu3BmFJ2cnzDQEpNbPR6ceLqQahhLlR1bMhVyXBLupcyE4l406ocfEAvlUU
6IdpS10MFbzRXocZsRBagiBdnL9rpl4sqYuZuUGDS0kG4aIuknTnaX7eSR/R
COgKw7ZaN+GoQlkv886LQmxE8VXhYViw5uXnAsySPthGOD0D1AKK74uocKwB
S1uScg633o13exKUgmtKmEOoOddtlKOXnIRT9E6aQ60ZW7BFtyYadWtsfb5G
JIfzyNHVcVm4Axn/u8pDZjIg52vawTcDpETRSdEMTmco19jiBaaB9KFVg0vu
t/tcIRMSfNF/6ff06LXYFHlXgOYChMaSlutD13kI957vHontCa0y0McXVbQb
zPte4Qym0TtEYUECSGInkbrPq/lH3SkWEFKRz35h0QB+MzS/FmYR13VYNXVP
YEQL/4G7D8zEfdMwHnlKq5f3B2WS6Xt1Bb7bgWZdoqOe0qaxeOV/xtQvsQQ5
+2ax3JmMMC1cIHoDvop4955GcQ45gmuvCFZSMaCj4qc6KA5BtKpwSqwhf3ve
6rB4HeWNDt2V6demdly6glccHLkNxPHRxowl5W9Z52UUOzZ45NDLA8bVD+Vf
6KwdAHDouhfXfI9JaLh8Xd2V4BB6H6j1u67LnXpsZp3h1g5R6BcZ9x2rDtk0
4uEpz++va8hCBHJmCweOJL8ZP0sD5lQvSXnH2XbnId4RVMrqeDhMK5rBGg1F
NjaCDpPcILYI7CVUznI7EQoyUSnauraX/SmnCe0Vd3KBJvrRzJ65zax2l51w
hoymh/gU3HS6FHjCzLhEHkhMqJw12weJfz9GiJDQLMK14qvL2V762kKYmXcz
tCfBgCmtguX6oeSYJnbSWMWZ0j0YebgREhhC6iyflgh0b3CG8Fn6WNPEXksJ
cTieWZrotzzNOQRbyGytRMAG+tVOGd14jalKZpnxaruLfvDB4aS02EjojHhE
sGlWMOiXit1z4watSf0AMhjaM2ZwDR2YamIy/BNl4DjLUDQRasG0P73Vxs49
zY8kzCeScMr/MqO1BzyWQQOPtYKtR6cJZKcX/O/xCc0IfTA5rOTJXKIVqHvF
JEiSD/59QyTlkn+tJ6I8nMKgkUqV7FkxEOkoqNX/Kdqjj30H7QTI2lVK3sIG
CALDJ/zHzqCugkTbteUj4sg5p0Tm6/4TPoqhMe8OpROG9/WIn2xet+KbHNY0
Czn94j1TY45MAj85fKYg+BVG/Xk1MZd2ddzwTbs8ElC6PMG2hGdfcKVLNY0w
2lwGxQZ+MxQUY5Ij08IjUjfBEvvGQccsUkwtFhqiM7uu9dw+aABrfRbTNgRF
B0nbLZtLp2rGA0aAVNpJ+dGpaUWemY8PorLFjR4ehfPvgxpXqNr917Q5Slfv
LFzldgB9meDszPGMjgysWN6oFShz8hLAG0429dejgbY3YyZt4EH4t1XlINgM
PmfBAeaHUPYU5clFriXXBqAvzjvybCtyEIX2hL594oD6inAmLrY0Og/ld0UE
de4NeQPRA73lPx0Z/Nq1kIkVKjplPomk4sRC2KsnTDJbkwLaHcI+8AT3+2bU
0rlvouMX+Iq75wtroHUs4bdOKamcfV7TAJSaLNqjYlNEnUo0aWtaKttP0dgq
SUsn1Ymk9AVCiMCs6sS9d2KarCdgj1wfn5+wR8IviB7r/qS/lJm/xmjXlquB
tP6u/u4lyjbtZcx6fCJDKyJSyKXGLl0fgAvKkkqeyoUC64xg0RZwF6SBxyNu
sCFYAEe+pUuIoMSQO85JOgHVbdnsFhREOuH1B4/lCw/Ac3nb3O7Nig2UMd01
pveNWAgoaBer/2eMOGwLsBuBPjdJxB98bNAt/gIy+dnND0DMV4Amg435DlvM
4SO+C6uoaPgxuyDutlm/2hz+1HIVfTbZnn72PRPhCZJ3C9lkbGd2LYzy0VHG
Wl6fD3psJI+S+90yZQysKMonamVs3/gOksWkKyJmcqsyp97Bx2u6v2hy6tZ3
nBbABnzLXGuoFS+SU184lJXQO70izqtgql38cqBS6DeXUPbd6nigCn1crwdg
K2VR7Y2bDFQtjFDScBLtmX6bImu05EdKSz7cjlYi6KiKXk5wNmUDFat9l9/K
ApKlGafi13/frAsoASC54wI2UMOaEv6eHU5OmAd99hr55czhtsveOzuPT/I8
L9oWEk6HOjO4hT5X0NjLeKsbzn7V+/c+8P8meeWdRD6UB686uXwx7gi+OeDT
a4NPssovCUgzibPcs9TBNcI3VLZHYSHXbItI30lV6qRuDutFnWfwMiw1tLvn
OUqNXvQrBLbvygg1kqbnyv+CsiauqVx7r0Bdzz73b3tL1hCtMfAkIEw2b2dT
lCJstdvqT3m4koloJCTqeoR8TBg73FmdV0WyJpT7rN2WnL7dcSmtfchhS04A
qfdKIRfNA8mz3jt1pkokAVrC1rniVN8uJsXxmhma83FWc9f0+Z4Zci4fMj9G
Dl2zPDZwyTmSJpMd3DwrYfRCzbHCyX+YlZ67Y1G5goPxSJxTpXa8Ue04u3ma
02H7WL/mNBpyvQVfQDFouOjzms8RH3qjvONOi1hKLIPEzdZad1rzTZW8AsbF
NWYtD0F5QGZRQSUkOR5RzvJa1bM+cwg/giCwepIcTVrjS2C5pUd5OWeE56Dv
5iIQR9ShEMepGLFIDrMvWJoVrQJ/jy+G10vzVsQvlUcbzBcTcCPy2SfVGCp2
HDEHZ/NbX2iaTV9GMyGAMktAwRwPnwUj33Oto6M+10nPWlbym65wH7kVU2Yx
Dr4+jbqQXxhP0+N/C69GWZEwar3ypC87TPMtRUaNq9F9WuhsyPvy2sFjnQhq
AsCAqs3ZXg7tHidhg+Nw7gcEzoZq4iWlfkiAb4yuUQRfMXrHd8IkLrHMPXJd
MfoqDjh06auutDSiJHXt6O2jWu2J6FEDvdieslSg9qMx8n3WbdUuWiXXTCta
WSwTDgvHDyMJlei4FPXjgE0X6TgaegYnLmr10plhe5jj1OI2esr8uQGO456X
D8hywEWqsvqdkA3ZyJtbG89yWhIMT1j6n0eq5B5EX8ZN/muvGCw8GeldEbC7
pof/88c37N10LnIn6lwheb6/WCP5kJa0N8qerVP8CCqlJaZ3gnqS2+I3Do/w
5sAf2orMdqKjmgg7t18bM9aG29hAvz+79hVwwR51ZGbGOF4UHdESbBumopAQ
mCkVY6P4BlGs8pOVUjixf1aUGXhtdRrMa6xrGybomwpdRh1tAWtEGzgu/nLG
BYy6a8AFiKg/1HtfdJsjBGo3R30kb26a3kJhpiDsWaBfTrQ8ATph6cttvvF3
7QRFCzE9hSmhe36HUjt0xO/TR3SMmCkeglZurPtOvdWsDnbmBXkgh5fQjFAl
m7vHOctZRG447rrCyxYsqwmrD6SvwwuiAinWzg+fHz4uUqe9dL8CqC+q9QEU
lEx/t8XFirdpyCo7qewC4PgoDdP17lxkf7/32ewCRZLFROhuB9uSHjOQpS5B
ZitgBWgpgk+iFrZ98aFtnYikv53A8ilU3+7yMSnzi4PR19oJGr57RN32zM/j
EUb6icdSZE8jZC1P9I8FRCjH0XlEZCCx6a6U1iqpOXl20dZsTx5tB/YsFqjt
ogzKcOUuDA8cKtJRr5JdrFMtxXbH4x+uFhPldz0BPHIXvo0f8CLDubeEXdYd
hhq3KQp+Hh97wxUqz4hwi6AQQ612BsowTD8NO3p1WDRTTWgpLEzkIlj08WEZ
mYXV5EmUdDfeS4MRTG04l+wXT9XA3FPOESoZEohyqyRLGmsIfU+icYpGzEq3
E4x7fit9DGHbPBQ5lpfHGtEpRiR/sSieoVkBqOCGy1bVSzDD3J22CynWHBqp
pUtPp+Mbu0rIUs75Oq1ixrB9KSr9u0gpmHLomWn26spnXsH2WYB0UltrYRCk
oLQUEjSzXFn/6ppZSAFuvVJP/xYW33afrNu6/BKm44R/Y/TxsLA+Xcy2gJx6
0yaZJGPvd+0+tJ8LcUoB60g5Rv3y828Na2is0Y9s5Exs0dXYxI0DMJVR5//n
5+1u+ftQo4oCrZvbXGugrYDGsy8OPk5es0D6MMe0s8mGD9MvUfyBC0WQ/Y8m
T/nf7DsfleT4ZX9mUNIPSPCK47xeUrRihrZ/e3jVdoQiRN+ynGNSAqvjrXtH
5iF+mjgsW6B/jNF/MzZD18MzxGB5Bw3Hsz/kJv8S4V68RLwxNUSst3ZKhCM/
6ZJoYV8gGzAyINiO56miN/Kj9qYUrqvKtNXVNXC6eREYkTk7JaGYqDZlv5yD
2dYmSSFNB4SqT8oro2KDkCdpsfO6lbtuSPTVV1qAm2NJv2aPRsm28/M5xMWY
7fNxo+1H7NXnv2zkThsUj7FSe2ef+p8tC8/pWM2ACzcbTwNBq4gKVOn4bvLF
bj1hjRIa7VPFDkUrij2/RI8f4OL5km1LYHdvU7z5icemdjvekyxIPH+ouSMA
gVE9KAIuNS52iwo2qRfHMepmJ7s0HiQSHzupkvcvcnVRyPmoPqY3I+NmeDnx
8+bd1uVrNEntPNIMwvNG/oPIDF0qIBCgRgIvl9ICuWkv4bWt3xNmLboXw693
auafJaorQ8QyeR8LfydM90mzHWsFse9NYbrzkgkcG+L5+MpxjWVFlg65GUY3
NICflUf+zrPXNQ5+fVwAoxpy7XL9Xa1pFtFOFrj66gYDDUnpFWXfB17VuL6y
x6umvV5MCbevg0pAiW34rMQguZ/nedu7mgQP08SzbLJPr9OtQGKE+fbZm3hd
6zG9VkRahGPt1ByKwEVap8PTVDgXqxfLVmtw71c4KNQHFPISy5+Q3LxdGYzI
z+IgMABwyMmDsMAbRSOO9XTGcDam3qJjKTIXUgaE7n5b0eExQaygsR/V24QS
HFf8uELyhRVnXUYP1CHfO4vm1j6hOlos5aV14CfO18YPzx73uRU2RL0F53rZ
UpTrEcLLrvUlLZP0Y6AENaJ6IY9I3lfn0bt6v6rxsI2LT6yPrfns36+uxkEc
M52XAJ8qxNUnvum6ojr0ahCUKdSiokSybNlWg/TGHTY9r2Q1q7QUvjQ5fs9y
04hssmXqZodKEyI07J8rE7Plblya+eMutZfceTU7LZH3zqzLRQ4cZTw8P36J
mOUseFMrCP3Mi6ouP9m15JYDVgD3Kq1WX7lLrQCvO52/yzrrra4/gB6/zQ4n
m7cg3UvtEP85BdXH1RlBTcJB/6pNPzUNjY4EFOruhl1RY4YP/NYwh7Qtq9VF
T5rGzddHsICAOrBj3KeiAuuZskTysS3L+hzhWIPSJh8wopNEjja63/sOL2H+
5tA3d1HfNYygLQo1BmtpGzVHbdzzfllZk0roQZ45oX4UVgVk7HG+1e4GHV8K
VK6XKhTLsqYmwwownvS2MKGlC7qpoFXVVdhehWnHQlPvkRCz9WVtTywhPIYw
KKcWjXkanVnihNiu8N/C6upNHL5Efyt2nDqt+pLYCAoG6pIzK8tVOi3tq8C0
fDCkimHHzYGtDzMMojKFD7SzttsgGBaoguJX08JYCpH8TtQcsQN5RPmL2z+9
TStnJi5sPP1zzF8nACRA2SLdXxkMu0PwYeTYxLDizfeQ6r7OMpbCgOctIwmc
1xHuLzke4zeOrHxjZZPepEam1FPIzz5mRlbDgz2w3+G5f0kYjrfP/klrDnS7
lO6msyObnrqahZmC7UUPFdxzuuXqMUYJJjIazIzGfXN9aHKPJMfE2/+AXVUT
MTAiifu7ZrwYHs9RlXmoSFtdPKRpTxgVUr6KzEKCbu/Vo3EnGvg6+K/MxNol
6J4OPMaqdnWO3RZIM+WGJUpZo3C791X1etXE4IPdn7lhe0suhzqsJG20UB81
5MksPL06R7ABj/cjS++1c89oxwI3/OWkInjwf5NELd0qINidL8YQ680KpfZ7
D3dodbA/uAU72q+fXRcQSuihdm70/UUuoKxYScf3ojP4SPEcdGoOIKQugwO9
UA2O/NWzkc06T55CVJ7jCWSYeBn0vs4t2/VZGK8KVrZn9vYtURd7POERGWeI
5q3T3y6bbQTHQ/PwfltkCgYgnZQtDck+aYe6WqvLh9hzJGWrQTGs0xChAX1r
iAJhO5tNdoNEWbaOken5RBoYamwFoQo9KrFzSV8GV0hsx3zFHLFQyng+oS5R
RvaZ45ttYIPxtqo/Zz1j33pKaLmzVDXZm6Eg9TYiVYohL2h8498enuuL3oo/
PKF2e+x+umJMQIfUAXnXBAYtUf/kbOPlzxdG8Nk4XvvZ2NOllnPaIX+BCpJM
OT5dafrEMaiiSxMP2Q4YsDFXxxQylfy/5lY18R2f4pYmwCuoHLjHnJSlsHoV
/Oa08fPhrTx3dLLFmVin2XrwOtYmxCFOCj5Y6su+JJVm2A/HVsjedmab/eqz
5rRf1kEMswdNDPDrn1pjQdHRg16OGpK7Cmr3AkhzYGbxdkoxueT25WzGCRsf
jqu7DQKg2qa6nBmfF/tnLSeoqWTWIq/3nAzh/bhqgpY8uSOe6/H3XylJ5gym
B+t6VjKYCaUxb1mxo3DeSTL5RimX8k295CqK4shzY2Rh1IgHcp4QQZpis47K
aLSSwTmy4tfauzuyJuQWY0upHXj4L21hJeXufLIUN5yqlvcnwuBLDxHUOws9
Ah4bLayzPNk22vmGXAI+UZSEYH5savptQbC2yC7Me5ECemBi417T62KO3t7h
JNKDXi7Rw7WQzCxWfoESm6MPsSjK6uJ7biomAIi4uv1ntcEYZiEg7NFmslln
uIZ3edUu/YAku7rPoShPwjcGkhhlf4oa4ACPUh0GkBnxHdAcFlnxteRAiDd7
0+8KZKoGex0ThGP3JO8ZKbkegQhuSlqqtRbSWJlhYmaUS9HZjK04EkSGijWi
5RvjWF7+8Z0mXRwXsKIfZFvtylKxW9vg8XlV0eAzip/iADQxL7KJ5351UH9Z
UoXzLuiaxMrWkvg9IIVLmedh0eAA+A/aVE1wOGgX6r9G33EnzMQydcFV33Ul
cU7I1QCVUFJ015EaA0XTEgNnFk6CnIMwE3Rv13o2Rr0L5+oYjXcCMusgG8lv
63uQib2AlEi0XNj3mE3Uq7w1xF8/7M9D2cjKV/z2x+x2yMSoimu6xYq7MTpT
mt7QPU2o3LVMRrrrIBE56PguRzXWxJhRUTIVSsKD4Of4h4ne8W2n1Jt5WvgY
1zG+1W9Z1/HWJ0Qof/4URru7T7+/FTNVoEz+rlnebAPYxzyXTf6dQDw57nf8
Q0Yovp5vc1+O2LWMlvL7bgPWhBYzQQG4TNqt/TXDlSeB2C+WiH+3Lq4hJW61
emRHczszteuVrr4sgo3JeP1mbGqpoBPGKt0dt5XJthmwbHj/61ob6vX01ks1
x7v3XnNLnOFrvlg13JAfNjk5MVn9svkJG5YQ0THS3hHFShvWTbkDpfYzepzX
pRNbBSXURna+gLE7nWnsFJv+Swk5n+K7zFzEl23ZAyaz2IrnOYzZWTIax6Wd
D1ErTry2wikUq/L8WmTM1HuTDvOfRHZK8jpHwO/tM6gAeZLU/ZN2L8rkcxk9
B5IzCmrX0SLOIvdXjOOOfVgeVc0yOdn+wl56zCrvoObz4R9TlYjOLIcYRlg8
Etsyu1bgXBmjrajzf9I5rtysR9Ph8eV2p8bMKbBlYZd+D6vFAkO8vlMvW8fD
2248mGKttxiv7T+HxW8s1PjfP4wvdLdGlDk2N3XDbUMbz3LdhA/Jxj/Pa1eT
N/KkbSsR+Hq8ovBJkax+CZOQ2P2HVmz93/Oe1PM3R4uvlr1waTXb7xE4eKxd
XLlhw86EVbKAw+mhpKj0iCCDrUunZxJ/Hd8cVByH/BzJKJfWdTLgGGWzDuH5
xtKC3T2mWKCK+zDbwOCXXvh3Wxx5PFQe+15ldrSfD06aQ2NEzTpG5X9jmyg+
TdRV+gfR76wRYO4SJvE4x3Luqo9PUQUziPC9pkD4JK3VMZS2H09HwjFiIYvg
xSZDsqZLt2j7La/cpvxkYGWwWRDXC+fLvs8Pg711VvquqxI2VR1TWTYeBoK/
ceE8jkzMaRt3w9jHPAUsiKnErDvWKW8DuABQP10zgr4kFp71AwvS0tOi0Lt7
WxWE+iUfSvy4nii2yTel4BMPgGZOCd7Kj0fmc0Hx53IQTVSPCs9LoNMIRfib
34K494oRr6WVtJxJ3MvK+ujq0+zjuuYpinrCr+fb+TXN1Lxq/eH4A0ZKttl/
HVO/zSHS4UfQhU+oshDpGWcOpdOWwPmIEqyvjw6j4YAHki8lbT7ISghVxbjp
OE/SExcJVOgmhVZi913lBaI4pWzz0Nr1j6BOkCIEFP0Ip93i+8N4rGN1PnIg
4mBpV8p/dAAu3ACDmTnQQjJlMLljd93ZUHH75nb2z+eqQ8QPtY/dPTA2jwpw
nGp6IJCrSumuSzHYY7IiOOEnHcDZeeVHvrSZs8X/BAmyhJJYQ/JbdTJxq118
aHx1voj3+S9lkYBsIoQWd+1JUV0HnTtKUISHvX3u+UFdKEPCw0RfV4MwOthw
ZCVasUbNzfrKiEmsREsiygTPOtnITGI63BXKXsAuan0kSUf/PWBzfXJg7i9C
2l5dzOgQJy90gda7d37BU6oO8VpvCdiRbfIJMpnPaBJ0UJtg674GP2rKZrSe
lKZfLVxRWridil5Upg8XMLmFU+ySGWrA0Ky+rl4Dpyr0PJdbCfv3GM4PlKPz
nKT2quiSeG9H4nfSmeHFDKV6tBeQY0IUyyDr5x6A8s+6gkJfL9gX0TOvDd69
ARAoSv1EC1pi2cZL3dO9csm34ve3SjiDDKCM8jwTbSuf6jGHHJ8L/6x/GvPi
yg4ecThgHbq57Mfr3PaOiYAlMzz869xfVNCZ2wNMe/E1/Kx4tjMz966NXuox
DxDesuL/G9VqF66Dy7+Fm8H11xdQlnFshOT9zIvLcyYG7/zwhVCrME06Bjnf
6IQnj/wX6RgS3RaI9zM+NjWWtRD6qxUjEp9ekl3LyaZX89AB7OnQSPTCr6Lv
kwY+hA387uCOrL3Ir9/Yt+RtT/6sj8NNO2+z9gOwbG0qnAcS4JkZ3yiKYqzW
iLdHSR2qvNfoWV2fQw3GFscQQqyJFVmF5GTeCMHwrxV7HHZ/5/B/2AS5GM+L
buS1KffxqAafDuFdMNow6ohGYP3vrIkJkkRiWZ8XLuJnXbyW/oQIoGlz2eZH
Ik6Glip0xqx+okoCe2VsfIKrmlHuAHrczj8H+r9Mo/1YtDnSqdn8055wJkff
ueNf6gxZMhuMUq5P2zZ0E5lnXWPy6eFixofn2dM7ydczx4IwHK9/NrElM1xO
/N73fkJvdfJvPB1BctqbUVPqvb9yf5wT2loPnwo00RtCD3CcDuk9PVULjK6s
54wMvo6QbQt4HVt4r4tzuP/O2+C+Fs8QoFEqYZxUs8TI6zS7v7qaEpt79eHj
rAj2drk9Fi5rhEhVi+eWPZrh1+JJLtGAwxvNF6GfzKDzyWYC2NBlRU4vH8bv
/M/qWl4lgDvpjfyos/SpfUmU4V9gIJFAWYOi1kaPM7GC4q8Naonoqu7OlCX1
OFUljJHP1u0o/WujzngqNIm8mvEwoQNs66h4zrzta86v++eaY5OlYoyWCGdE
QlI4GlAq94kRcG0AsXz5cc1U7gIpAeXc84hWJ/Fxqs7RW8guOCi9uKFyK/1M
3dgp94Oim5xSzS3qcCiykUSZTfwYMBX87O/lH1LWAZKiWRSZvfkFVPg/vZpZ
x7pdiuNoEyMLcs+qSzDhDwBnTYFFNVD0WZmKEB6czTf2onyDNKVvXbXTIzQZ
cB2oe2Uq3Vl9kQ9MJgCFw5PEhFZvKWwoS1jQcd5rlsmF3EODVs40OpBtCjxV
8jRbPXKyiUM/03D1Be0/o/lGSJVMIzUmt6GmubGDXuTjEgvLO0ZQXvPllGq7
60xQLzcxFnwaP4sYk3cvsGZxhFtv06QVhUc8DCztOdZQmRZXiHh7ymMuLv9O
x1k5st85nhqNGepGsyo5blAt/pah5DXGRZOYl0mAHK+Jt0/bbpw2zZ7ptBRF
A9YZSYFDT7z9fBPliNTDGICzaacvlA/8qFCW19OiZJMw5prFYS6zQJYkitXY
RuiP0lsDZuKFpDzdYpqTWx66XpQp/mQqTO8Owign5Nx/D+9bEgwfE2JLqKAP
nxiPtqoOQIBOP9fXPMpEoVNGMhhX2xx5PTmjC5LJVSbU49nsr+Pop6eWjIDk
BWPtGwxa8MeWLDE/BLpsPFYyNJN8ORQlVkAbqggY+BE3jHoaW4wpG9NdaNQ9
MEZ3FZtZ2hl/D36victsRlDuTljHJTqswO22v+RVVCOxcoiisd5t0fypPoNd
4NxcdaXu97sEOqqoxFULoOzDz0IfVrSGRl1qLSpbYXod68tvtmBHyksqnXKY
a09pW5ALbJ/CsrK90bUwSvVWYFNAEWqeBrK+QpYs473o2xXFyOjQYl0U2P5i
CRd9r9ZuqLw8od6Srq4/qySB5fGoBY12j12JfhNY+2hxXXRJtIBAHS5I6HJT
pyXBDznSBzAFrI9ZgxUHfn7N4ZUinl02gpFQHX6GdVi7hkaAu7PA7rsPMMAl
PSOxwvL6Bl9SvyxPynW5TmzWTudXERRt36uQB0K5QYPlm4g+IRCZFyZP1Lm5
wrNZeiKprLlzhxTdXePyQRj43P/IFWmFAwK0/gLJQXkGRvZFj1quDGCUtTdr
5y8SYZ8o6gz78Zy0B/+bt7uPXqJ7Tb27DwacVQ+MdGr9tnB8OmBLM0f7FmK3
lTN0yfuRlSRhXO9fT09SsGgL/F6qAqurgBKpGTnDO55bX18iTkzZqhmlHZdI
m636HvlTJHf3efGpRIwmWsgB8928pjEBX0FcH9m7liwZtl/XvcDjmvtXkEud
jVmx8/bWIjArSpGRjOUJGf8khYrdDwgNZBIBEmAbMZBtw8R8PlR4Ucn+VUlq
953dY8dA6p6evUdbx/ehywRF4ACmlEJQejoT0HHmFP0iAB7oTKwf9dihvV96
Dl6ws82Sj6EcucV8JJ5gr4dJfxwq1O7BeFNz5/fdDyhllvA/ZBMBlVcoV5hZ
gj3NSWHXBV5V1J+uoyv3k5wIHgGJwvWhjDIhJocCCQEM9olLjiGD5F29joQZ
DGozRG6t+orvPecs3MAsosV8ByIgGNuGn4AFoJ/6gBnh3HeCaeSHM84cM/7g
wHviCk6c9ulD18lsrgOECSbrSMnyi73XBTf6Z6ATxVzxD8avJLeOAbQkDw2/
fUt5VAHiYKfzKSmLbSsU9rfhYSBZP3h/wM25JII/v5Ff1TMcU5vMLiAkGT6p
VpuxBn/XpEIgEVbjDktzgRIDVlzhjDSmyXfiAxi6H0D5uYAcoUmm4WvcYF90
X5mh2TwbjLGwCLmBpJRXMviWG1maWYP3sE2f9fV/g+daBB3bXoUo0cA6kMWP
LTObpDKI4riWE2k/kksziWKAUOjPIz/o0LVHNMGs38qFBOjITIuIwS52PMNm
rKUFmJv4AXAkbFdt8KjkRY0DdPKmTxT3KyQc99CVK9KPoiN6i1VifTK10VTO
cFo898gMPYsCHGxSNqt13QsQLkPM3N0EmDRY+rGniYDUhaJVJQ7OhpI+DRIj
8OWVsScuvF7ttUVO1c7b21UaYOiC2O1bFJIMygmbg7SJlk4WaB6ZH+q3mPgi
4KsFcQdgCWRRgW1FZfUwRBKJXeXLndrymHuiALoLe/eTPQeMCw7rg7mAkCpK
Lpw0vr9YCqhPZ58H5kmJX/aYLqmSKVA1dtW6iWRgV0yzd79ncoahfSGWvxiO
VvKQo8x4zceoV1eLN4WAiTxHEV96C+gh8bIocpf34MaelwZIdF6qMtanIrXm
VmAT2hnvUsPlBk08Vf5G1Pyen/MsJx6D9bNbBJhzjCueBQ+qg2cngfnIotA6
xTsDIa9HYMtqWGn0no8eU2RIdKNiCtvYXkzE1B3mXpa1+LO1Hr4IRFHuQXHB
zzw+uwvcoattdlpHDo1iZJS4DinmEdaJ7Ld28OQvTflUs/PktBB3EKFsjnSM
+9wGlVAzBZ7QUWfQkoRvq6/c5UMjdK7KdQGiTfIH9bnh34xz77kFYKQa9zMY
lWrfZqBHFfwrtqZSLj/EY+XMHjsZ7dDUhsvpg9d7DTIJkfiD7aK2zIi1S4kr
3K6H24UIlzWsMejTMTqv1IMefAjc+HiIt8qwNXiOiGBF/riIKMp9gw9DCinY
fS8Q9dbmmSpsiz+riGGKQUOqyYiZjyIpB4wZsoeGwiEN7IAfSBDv/58jY56R
9EKjtZ8aBMO/7/WOr8KSYutdchprC0wdwUdoTFNNi9uVIVf/8ADTN8cvu2YS
0XGi4tP1hG48UXbxuvWb5FLwrqEIJgIEmAyHCdjBPWLAjox48kXr3X/Y8SMS
ILI6IQ9YKXgTHwviErmU9Wp/vKze+2pprgSSwrhz1HTBEDLyEAUYyEi7ae+t
wm/AjfCyGWJmERcykU0fN46XK2Vy9Z16SYlvGZ/yQShQ4FCi6Soz6x3yT7GQ
wDlubh0PJ4lxq3pWvTVuNbJeK1NXKMLJuh0rBHNT+8nQUioU7hGXWux6Q4Au
p1cJ0MMgVjiQzE36UW+bHW/207PHbQ/af9dKRiBef1BOTZHK3pBdWvgIxI/4
TYnT40PAtv01MoYrpNDg1ROySj1rP+7F5rxxsvfn96ZRosb7iIFnYoPkIe42
mYgobcOu5NPpj24BnJUbKDhZsfFGbhWnjqJBDZM5losaWukCk4iDH3hAWnRc
Zx2Exk3tb3SDgNZ/lSm6T9EmQwWe6pxkLZFtLMd+QjEjKB4qpjQrTGFysjIP
JTghhUjoGkreVF5aRxyQGIZMJpiKU89sKrskI1LJCx1koNrZ6nKyJC+61UvE
z/YZTdLeDRQO4K5fIWw3EnMZtj2i+qEExlyGRmCnjneKZca8TUOh59TcpHMB
1C3Y7cBYKEBqvYhB4x8Y4+dfa5PbTgW44nWoaGWS3VW4/pJYuzE5wo4/lNef
86+0ZTEzmMv6gAYvQs+bioVP83UtAs/5SE403fMbdU9gSlYnkyDUkTRX/XNB
Z7QyAldVMmPQIpiKpd6KDOoayJxNXr3CkSpJpJ2wgas8hygjP+JwIv1edH9m
RvUVP4DD76O21O4sNgb0P8EvSxohAn6j5y36elLtXry9ogT5C2kJolkVCudx
pXG+PKN9WdMT68J2VavlDYMEaiqOeMr9aCsxP524TQk2m4vfJr/NLdWKyyPa
E8HOipZWzaBjFa3VrYbkYEku16bntFO8k3TqB/Pn/GFtohcIoqRt/kpwWpJk
jMPH9Uf8MrA0mj9fYW0hbqrBIXEDSdnGUMqDFDWL4DW6Y5Snk+28qKA4hysR
AqC2bLwN6Z/aMfAo4SoCNn12dpDnjUkZlSUDni/84HmMlB0SIAE0nvzOhWjL
RgymNi8f4AxB2AlNdlxXNMFS7poGIN/tDhXGbUXub8i10NmgWMBF69ZB3B0E
W/Tb8JMptVdZCvQIoLh7Pb7pCUlvN6oEHLtDDyJK7QFHJSakjO9vDqx4Vkqt
QKqlzrTfrITvUmvShsP1iKJmEDkYcUet6TA6eGl8WELoqPRu8haVTnae+oAy
UdtkjAQ/KIOnrBAvE8XDbpsyiENnb3RA9DqQHZEk+RGXvehlaK1qp/afvpam
lS3nvlmrFsz0bz4n4s9dTzuPjGIiAi6H2cjF8OAGw3CGYq1IpMhkN2RYHdrs
K8bKmzeTq3dUkEvp3MQN5bJC3zWR0VCviRJUcgfydmg0WaycGmK4nv3sk5XK
xJNz1GdMzX6yplJJMZyQJheHxZM86J+6VpqtdkiidX5dUroOFqjXvOAGHj4d
Oq9sj4RW7n5MJww3C3lm9v/8LRSICNAzdqpYVyvmJmQUzvCWzRrDg62m8haP
u7zCl01kq1ZLpTx4WTEOqiwTdOcouqN4M1voKR+jwmkQvMNxApAIDCpq0NnD
qDA7kmW0jI7stWe1HLMwGH9u3uhUHzfcVWBIw8R+T/o9ZqzhAwKVE7wmz5ZM
gcPIPBj02GpHjeny80GVuikq6umDuJ/phzQPZvfuJbjlaF6dW7Hi+5OpidA+
2sJ8ghbbE523ShO9Z8C+n69qxwOnM3auUEXmqnVWH6jRBV7d0hew6LqzY6S5
8i+hbaZ6VYvtCN8mnhtLjsixcOD9gOuQeq9ETAjQXeFuKt2lcjU0fHz61cUD
uPoatC+CslX/LuKiey0Q7vZZYBMjzIYpvnwMEvtVUv2eKvRpsdhixqkWi7pN
oC6738kc/edNzZYaYvGPktnvjii13yiJ8gkNU3daZVE6TVHfzYnCEOMfyAC+
t/XRgygZV4LQ/mtmV1Q7fBEBHdRQU3UF/4gfpSvb66YmP7+LDwqUgX4b6G98
TBH/VsCcSQXibqjwUz2kIqwTSpvzt/eLxVKGnIbXqN6refUvRTCqwwG7VrbK
JVBzvBvUx/JUS5CVjG2Npd9XmVqD9UyZNK/txCUXeyVRnvwrMT78qFvVl2Au
W3WTCVFBzRQqBbKgkjzQpjjdwiYIxgjWB38r9a4UqX8IxqsO+atDREWrDHPQ
xD1AzaKmXGqCPY9dppJhXEoAbFdPxR2LtbWjd6aMdbTAUM0/iZAl14MAAu80
8ppisln4GHuc5BjSMgRg82auXayZdWK6rPORb7Vbh1MUmm6DB1KXBekxyRPe
iCNPHXOwvbFzjdSLjLTRxcFGgA1JyV4+12Kp4A5xnmXps7VRkc2ddBb3J8f6
eC07dvVSavi27yFegeyMSGKFW0dAvL5Nu9NJrvxO12FPt28IPGUkHtX3wgN0
yV38rT/bGsSqqyBck+x7z5tAqfcoxyaXmruvzrp9IofzTA3BMrpVrZfyE5yG
WvAR2YqFm6OHHKhE5fvrlBaCd92t/nNPcYQHZQWbYzKaPTKwzoBfFZ/7d0o4
aWOAbRSvTi4QMWiNCWTS2WE4p2+9o2egxWnR7hEQ67tvrNNpW3qwnjAZNEMY
gbMispdw9pMtLbpUFSE4XYNt5CozFF7Fe7HZo6Xk4YhzccLaMrO1r6lVZvjb
Jjgd9SM8U9Q6vcY91V9FtrEiBbi8Xav/j1nYpLyqgGxxqu1gTJqTZfzMujio
QWwYCij32rP9AqqurKGWgGxjvShYD0cvhO5TeXtnzDjt9u/FDE9mE/a/yb43
rwOT+4xlpl1CLGsEesOscf5+MDuCwhdqqFSrqt8mXwA8kzMa/vu847/dfsoQ
APUznFLtkaCm7UIkNi+brCOuDm2a4gTu3eOxjfAG/45Qj6/dXrg7S09FtHtX
+FwXJImTD3QMxzh26Kg8J4t+HazPdphLWp0rLGcWPQMycsz8uBdezJSvo6wh
pTb9VtHRfBM+5WJJKuky9c3nEcPhD7L5WokmXJVhJNQr+1MZ6sqWl57t8+q5
rkelv3bP91v+6hV7SKV6LQLQ50avfjS/cL2pbi4UGICB9VmO/gylQo25um/q
6KNUiX3FQdwjlXmrEIcJsSN3rjKwWTDEQo4Zi6+cdIeDAYuO6TGC/1ijQQr4
QisH0Gc6ppn1TQ+L90KcXj1JInstHy/Vf1sP4ZtryLsfdwiuviv3XuijSNDW
PghJ2ViD2fMD9gbVW/vplx1Ju81lYmnXaMSekyY0hG+cMVQeOy+oaTYDwyiy
YL5XlIiY7IDQiJIQTeQ8flhP/eh83+Kmvj6w5gc7QgNXYOgORKP04FPPpFiQ
xNslQ+CWCI6BEohq3kuXPxYWFnnsXLtGIhhquIYlgyXEP8bxfZD0jUvw8rdZ
GpxA1wIaXxTF1BUzp3+kMvAlj5znk19aS0d6+GxRFLL0FEqV9Xt/HLIXojfx
tW/yqEg40osLMq06i2Zr+t7NjTvoMhLc2X6Pwg6HQj1IbHbv3KtSE/058XJc
UySGefQ9YuEK8J5jD2+uCdtjMomYJWCQuXFAaohCNJMY5tLK4rXeAw/DBPJf
MiLVITX07MO5PVBY71vJPCN3LzM8wM1utQ2uPgcoyGb0PuaYPBSBsfJCClja
0bYmY0gjd2R6wejZ8N1RTezKgsM6ObIlMEVqyJF+df1eBFTlmlaOyAHS09ei
69YEGU+A2RYXwLwrMuLONOVWt3I5vjfgR3us57+0pmBsnzqni32eKnbDJWGS
xroQxcCa8MU7MJtYwe8blsSgA9bCebKm3Eyz+yNO9vYOuZORxzfyHeSTaoKs
frDMtZ/rroIUTs20epPhN3Y7jhVfuIXkdJjxjFsic7qWd05gukWfu2tfFfeT
+UsIOpWugoAm5XbD3mRPj2Wq0EostF/WC7eMFUctI//opLFqjQ12CvigDEKw
liN+4hjnU6ngssep2oHQ9MbmFt18BxaMw42GmL5sQuKfeTeEPjqBwvmpvYxx
FBXb9m0bCJnHVq/BW8DELK8PZI3TPwNW3nF4/T2rUpGyGYoLKgal00ZEKrOk
MyF1U9fhw4PaithI9D5Vku271/hoI9qc95F6HhHyZpgRigD1QQty0cyC1A/i
6B+zx3lRWrw7Lm3+9AcRNXc31Iy8C9CSI3QiUZkeotQfMm68yO82m+6KmexY
3P0+EtJ4cqQMSn8IwCBnNKJ2cjSr1gcj8XoFhWTawrWXE9zH89/CxwZhWkwj
8V6uD8hwNpzzzxuQNeWdnIg4IEx0iVWne/p7w4BMv5itpexLNr0l3o9ysxe+
pp8I7bhHxZrLHZYAXYGW0DOqPXjmgLqk+K4el6FdbyzhLIO79rdVQ3khYdhg
PfIgMm1JBwb8AvKoh2pNeFdRoywhxc9ORotCl+ds0OJONOfi5mskkofiMyPq
G+lJBEzIHDjz6ycOIsXLaJrRvpzfdu+hsClxgPb585vbsXX/R8gysicjx5mE
1NVRH1erSfxhQnzOsBG8UqiiN6wC72LMz7RxpTzYeY1KKjR841iW9K8lT6qX
2uUyErtBqBcviGaQH/BOEULb22sqxCgBP+kn80wl98kLKgZCxfMqZ8oiJhNv
cAUaGf6IldnW8T8awO3uR+Md3GQ18OPH+x+kQ8tgKGEgmj0BC7ax8rdnlPg2
lAWo143uvuIXIqlN06sCt90o49Iw6D+cFq49RPxsrvEhcxJYdqNrKj6iUDXn
OxDkcBJL8fJKcAdEZPAWcFd2Yb/8GlKtJptW2mRUlplf2vTCU4293Iyjxnkf
MXl6Sd/5MygT3x7Ng+Y3lxn1wam3jq79nFXVuZAwuVT2PYyMjMVBq67RHXFf
ZKMCKZ4U1OXVB6c8gymM75pdS+XlzcRQbfm5FOWc4jy2uybadBcWWoS/ZFYf
flxK/fjIHbXee3sHF2TtquL3hqvuo3zyKltSgZsy7170i6UPeplONcBhMOKd
dK1VUrRvyN1gMealSKuFY1o60Cw/LSzeIgIj194Ec6NejOBcyu31vOisZT2A
0yM1GqeIuoSMagES6ZJg8tuYm3i+vK2mREgkxpD/WsbwMF1Pz8LGrsbT08wF
+RYJW15AZEADPrZK2MUnVPlpG/1zVm6jcz5vYoBCKciRlz+TjQdfmxmC43Is
J7sDOVaBNyj9vGRzGPmfpoXUvRbOF/+oGcKgYlGXWp0rXA7+hLynzBa3tAGP
+Ke7bfB98IdtNlrvzsBR1qH0GxSwiC1IlkzTzqd6EyVwxHhuEK7+2eYgLCMa
2BYVnLHrmqUsu/AVJJihKzpCMhvYvHFBlE2k4p69N7DFgZyzvTPHXDK07bbh
1RMtKZmZfEO89Oi6XBZaZdPqp5vPr1NB7jzzcSPmwjlKGG/9NnRTygJ0P8n/
WWxsSXA+Ob2tXNhQq8hz1zKnjkZrKWLwiH2yR72vvUID3thyeRO3uA3QboNv
63PU0/X9qW6uJpMhRKn7fkbF9j2kg2Ppf8MlKBFMwq5i102tv7NGNxEzZUOp
JumWUnaEFV3LXsN9K0L1OxNJwUnc3+BU1nuCdACDGYJqa6O6mGWndg/FxYAi
VwbwgX0ty6xLcOf5xx/XfNQR6tJ9ac4YcZ6rk6r2uAvCQ2NqLng6oy2pyGm8
k/fSLhM1pRPfMmcWPUSncZ9Nmdjf3PRjTPYP+DBFr59Y5Wt25y9QpG97wr+0
qZXwg20eYEUzORC5dVXfxCt+7rCYtBZFGJk3JWMHh4+klBvNJAHyON74e309
mXM2V26MBh/C4P/kjHacpIyuK/JygBq+uxeq+3ugpZZQ2cYvpGhBFARYtY1W
1THSpVxsMK+8WUXbLNlkToJg6d1TA74+a0BQ714augZRC65nAbujt8PYRIH6
ytx0zE7S5XxQcYA70SKT0hhhm2Bs0jiJ+NJBfY2Wpugfd0KW6qz7fCmRSE9l
XiKRQ1YxPFS6EZEE0ElLfo5q4qy9wmDJA/UDmhCM8fnx9mHIq+zpHNBGUjPH
OEF6Qe4UGu4mIy/8n/1yZKSE+f5rs4p9BnUVd304Svi4f7C9svfITfHWZ9Z6
rtqawbTMiwp3fJiCCjXHEG2StcLQ3+bc93jmtRToMePy8yW7n9y5puxIbuT6
1a3Ke2llwflrLlbCJLx3jhoEv6olWE0in3/1TmqxTp/2I9KcMuCM4A10YZD3
ezHrEES0GX6PoiC3DRK6Q78bJNCl6p+1TQ8rchu+souHZAS3z3mgjk11SGgv
+3t0V8dfGwr4nIRfpWnYXchtkVlQbI2nyzuF++LBO227AXCvV1SPuEQGhP+m
8cikrFKRuOj4ZO10Y42bbB2QXXTvTrJC9+LmoLen782YnFxk4NcF0LS+JQhm
Lu9oAmZ23HGNkc51RU1JFaHJiVBNpN+MxkxFi2/XyfagT7QruDxB32a8QyC3
EZsVmjlZF/LZrUybln4GgE9LvtRAPq6mdV/32eSiK6vRWOf0uIKZRm4GR3ZI
LjVO0JG9JXeLLs5+xP/z+0uHY6uBVVAFZ3RoN6LxbEdiBfgqdR+uDQYLFmEW
MFzhmwaAVrLA96sY0ikrETC6Sd93XcvrydBCmHD8D06+KgB4CtBo+9fRXPeE
zJuutIrL4j9WYBBbCNDLDE+cJLHhZNSyeiFvW1djtiLnIsgRsJQ/JZw94F5t
y9d+xIdK7f8HeOFaRd5BEtOmCtoCt1Avm4TQN5S9pGWgXt89BeJ2wnPHr6Ks
Y7sMcqq8xylMfazOdtBIXWmQnJV/nz0tNVX7O5u0gKG1hBigycVWLlUldi6D
pxcliGk03yz13kiCU+ZY/VPoQyQfSZVcFsKaIRj/4aQ8bmqPKFp66pVfGqU2
YY+7MgOxfvRogR634X2yvchNddGniZlksHz4gPvSnRub3+rfFJazJe6Kt1AM
/C1po9vCREDEx54nUGKEbFYH56XzQWO9trbIOEzM1lv4qn9AchicIPUKoKH0
04B+mjHvFrDjZNbmdiEV+iliWqWjNxtta7bByurTqCOAXQQGnutTX0Px/sLj
QC14N4hpbVIpacRsNNJFPt05zZIXsJILsX5nqL53buXy8qvYqsN7CrOLR0u3
VLfhjFrUbQGXga/rh7IBBCaHEEX0/bP8MlgQtnMmombMHW8mrm6yWuGXSwdm
6blRJxIMpnaPk4yTZWM0p4VFLigg7wby9YlzLoPJYN1D5BSWDWVI4RGLWv1r
Mz33ExWz2v9E7CTEf6emnFz5AGbvbS7qbCsS6x75oGNdDVMwYN9h8FsVTWip
JpIDJ3EjcVMASOfSWDeRfhAxjYLXR8KiQfhqxFswPoXhIOQyajpNhQGYl7Zv
qLNjIJDG7ir9h2pHdTyj+3jDjDdrJgSr/4n1kF7gELe4HUoNuWVTnEPdAVfj
/CwYKocxZYegkwm8X5UZlUbSnKXJOQLzu+DLVKuhTEuW2jIQMYODsyjVn8+9
Yzbsz5/mA5maAhdQBKiOVG74IMNNMaGzWmeg+kPrhtGbvkjWjn03NwcAH6gN
1MuVyGpJXfhxjaPnkrKLIR0cE3aS19JCVmrOvT2dD35bNqFQDh2/Z/icsmV/
2j4DAYukqtgZSAvdX8Ui0uqf27fukxavnBUXipN1OL3uphjmZNZFGltS0KU5
co3NMn/Hln4v34kmgzAEqyumpn7ypC94lDleiFMqDryOM8HAVsI2vBM4j8rk
AWo/S2+qA98+RC240u7XGjTFaBhb3y6zu8xT+kxSJa85UpTJO08GcA4ietyI
nC8jtb+aDSeHgn6xKN1trFSonlsN+jf1LN134vTAahuV9POIrIHBuQnb6C8K
CKxLgBVPXz4cJPVoXveMRprmXb7d7vhfon4DbawcPAFg9Ko0wxyVWvnn45Jr
ZNDi/1inArCbgiAKL4RAbarkDAuPtGfgV69H7bhwQFVXzglVS4Xv4zLQpMfz
vh27hgYI/3u41u5AKpwVvHrmjOfwtOWmb3OJ7G1wd01ZOcOAb9JT7O+VE1FC
m2yvdkbp9v7hE0xcbJ8kdeHAB3Z3ghTqeB8EBh3JLKSW2t9dsrpE6pf7RNU1
czvwaXteSD1TCp0+vBtlfFNciW3e+lUHJLm2lK68nzW/w/Vgl71+rnbZBFqT
IeRiRWFdvCcd2Zwunksl9nsFLezlgxzoMhjm0hicCoPg+/ev0J5jGW/5Iy4Y
LB0J4N/JYcPQSh3s50Vu51j8ZOBdKBSIkLKDYnJLzyqxc+7VKrrfaD2v5HO4
lI7EQqdIkhFg5aOSo+4MPK/GzjeuukuQ2jo14l4j7IpVJYJdVFcB9RbhIHGb
JyeYiozvUEyHO3AWOMCiBM9nZ15Ab92pd99ZcluzVy0SaQRc3jpk/m/qHI2x
p+5vCABGcz+tmASUGTmqsnZbyaUhQUwakSwZfdCjmN2YEqQRwA/6efe3QxsW
vPz8JcCLOfyFN8gwr063I7ugCo0FBjSIhT3AfN2PicNSUB6JEGm/kgyv5LVG
bcLnRA81cRKzuwiIC0stHpfF13KEEOAZoV8qmbTCxUEaQO76lqgVcCfzUfsY
Pnge6icX/aXGyFnoVzdKObzB8gAHtuYocmOuTI/kF9abPKwK6bVS5ddFXQ3r
/QLPs6LLjq6dIbLQraaKLPBUJPkodSWbUtN44BWzeBkfk2Z8cfUeDy2IpYd9
4HmgctcIjyw5RIx7X7tp3vXSayp8L7eGwFDe5A9hXnFk3cdVnt3v3ydOcOSy
j0zJJFWWGml2Zy9DhkMD4EpsG9KWYV0FufuUv9Ys2xZUljKlCUtxPG1OHdTn
mA7Mz04ZPwBfWdvCPPC7/HeXozUIdeEjsc5XVh3Sf7Ry0NbXkSh7N/j+cXPr
vPs5PhAC7hcQJ5wiXfqRLb9fw3B6vVaGa/1DahHbTA76Vw08Vb2Haj9uwzx6
c9DYUz8M1eQgZkt/+rXvczxKBOt6rh8wagseqgql79J3Lx2/0Q5HlhQ26FG/
5BrlwL8FI/xERKf4jOcDRjpQeerixg93KQG+lfPqVUIrQBygHc1c0eUrUmfE
eAtJ/pon92YeGa8nRPDelfH3mQpFGwaOgLrwiWoLjamucdXrKJsPK4gbbwkY
cMuQ3vBywpDu9R98mT4t078LqV1dxqxH2lG0Ob05ZenZqNjp35XPLMAQrMfb
BbrFYw9WQo1Fn9tNeH3ekgSEqIWybcWPnQnBw1qWa1UBINpw7DEhO/YFCnge
fI3+SFW1XqOYkBBXUK04pztP+e2tDZEUMsbLAkkovr/LoeW4fTifmjJEWna6
Z8SKrdje1j4L5qmmW1775eOjR+1fKkrnbTJcS0sOljFyrqbf/OCHA6wYRMm8
NvAoG5J8ULUtZASogTlW16xSTPXf1ldUtOOQ+eHKbh9xD7AVPZD/V7vupLqv
aZGMDgARohNI2XPtTExkXKOstKQ+SJ13utEZspzCRIS072c7WWi97wwGQPbV
7zHa22Yhe80eJ94CiejJL3uMnFf9amJZvtpC00XeMMS7L/w3Bq+j3BOINOWw
Kv/ihBP7yjSCmMZVuqg7Vzmwdk39c6E5dbt1WiGM42EZPAQ/Xck+xgV2QWDU
Sx5jf8pqLIyhOUbcoiWHFQ8YTbcCTUGUHvbgNKDGyjs5xq9MVmIxfBtacA9U
+vYH1N8Rh5lcWZ96IwDPBC0/XUzu/MMa10bCUvLANs+Yp6I4Y9dkhRyjZyYU
/jywL5WTeqravzn1eZlGXVpFA+G0mtJurRyCMk7CxBeKQCvGcXUYwympFOnX
YbXq3VCNOa6mA8sdSQ9FCStvc3f9pBV0Wn9bN8Hliv+TQv01ax6pwZ7JzvcV
h+zUvxZ1Z3Yxqs11FKQRywQjXRH7Vkvf8Ofy1I/EsHMbeeD+sdvKSWtZYZ4i
FE6tyT9nT3ae7qN3h+YvCAGg4d5/9jQt/cPs+a/FB0cbGrSRIhYb+kLC3DpP
6kBAIDkxQqTTXyJueTFsSXdM3z+egLhkzJU5/UXOin5A/kfW11dfzBOtl+xF
zjynY0AwGl3rmY/WFUQc35ZSC90NaNJ98yqMSRpM6me0zCd2ONbUOa7M+k7Y
nkJQ3NRiqJ1d6wEfFf1K/06LQsGSgWRbGJWbzlXUdpF7m0CcCEWafCjR0SpL
2AAv8KbI7ah/DOZfbtv0Y+mIivyINysl1NTtwRpVepa8oxKi04Uw6EfxkM1f
pmPutFQbrUNN2jddNXX0F6MQ15kSuy5dW/arXldUiEjQ4s6x6Fwauy1SbJxj
9jthIxp9wvidtG10A3WTuZZMpRIKrnWZSMh3ghBvAnYfBcLCTIs64f8CyOwo
Bfzf8QqNUA7t/ILw64n18HY1cA0C9ZWNXri+SJ3V8Z9hSzmd7jyFu+Q+9vTn
+GhpkJypNmmkYQfJnnIj39yc2dykd/1lYF5ECDQFVs673LGc4eyNotQNXWlP
9Q/TGsNIxfkUiwZg1XlMsVDi/lPczhOTsafw4eGnIDVcSb1Dxa1A1odQ7OwW
+//CHvSD47HGBrH8A9yxwLl2vbfa8+rIEuq741u/h28X2/SypISoN6Rasv6U
TDKIhzcYnDvcDE8SpI8gHcz99xBFpoM0CLulNPTBf3dSrz/r4CgRcDAwLnOq
3bdwn9VnjuVwyQBgsAx0nvGoJaOMPoRWpd/qe6ayCB5x1la9amleC+vaWO/C
kxzB7w4HqPYHp/QqeC2kIdJnI2HgBnKSSkZIY4a4I/UysfPCx+jUSSVbkORf
n+iD80EB8V8zWKVMcZyYNXinvT4ecnOWHUlp4FwllUIRN79eMl9Wq/y+xFjO
pAGFAa+A1f3P7qltNALDBq3Fdex0An1a9cKXOGQkzYdStcWhSdgMV4Ld8wi6
AG3ZJ4ZStt42w9uW4ZkUz0MwC8gwI042dUAbn8wOlLl7SIcULnoBuaW3VlCf
YXyaeslfhuSBbQg/c+aAP8tDGWLbqjsF3Hgyl6eHtgYzrC9/rozC3OEh2G19
R6+n0gZK6LsY54nSC7VZff6epg5JabLgVXZ6I+PjAxck7rCPvjL2p6pJY5Fr
Wpqhtf4+xGCpibcntW6AQodpqYP3g+wwNVdAoZYhexhwipxP8LVZMz04x3Aq
IiDwXYSeML62gbYHS8So4h+p4ak15cWvCmFx6PKAC6GLadUHaxQfNcuxiHi2
XGHUPXrEw6RKkOQjQ87qjGMJhY+SN6GFXmU59eSFY6OMXQKORrvk2dtap1mg
0OK+KIElWh0fCU2mw6dNjE9Lw3HUOT+9u+e3Qt1MDaHCva0Bny0OlL9N48Lm
hQzmmWwc4/PcmZnS36790MukKv5KLIEyLS2grwfAN9K48DUTia5qvoF71JYj
WqkeRCFbsfK+VhY+ugDYFla+y8Kni6dO2LlhR+PL3CW9MQsI427QH+BhdjON
imtilf+nu3vYzFKIi46gdXh7a9kv5nErPHzG8pVa2gzhcu8/50P7OTZ9AaK2
pSscbPpJPsuTePs9sOcnHInLWjhXdjrbYZ+Y5yaU6IA/ORgsrPp330qLucgJ
FifLSV5XUCyw8PsbKkGoXOaHmprd1L/U/YhvKRB8ePHOkCZeTPDukb7rmG6B
CIc9jfSGChAc/qCAtRKhImWgizQNbh4JWdbvec9q3YFtspk6diM0xcwKRL02
9kZRVw4F+LEfk+AONVmoN+vWCckFiynAS3vNGadH/aFq/x6+0LdE2lgerXKq
8A+k9hVhAT9FSf1WBwvm5VSDYZnlkEt5jHmWo3JuRlpcAT71NFgsMZRmV+cC
sn1Ajn+jCCOiojWEmPoLTPztFTUL/eIQ2cRWRIU1KivTL02eB28St1HJZNny
hfEMP0LsabviqEHCMvLq9CocfhpyCXaeLPennO1mF2yF1MIIL42IyjMh03/t
qOttV+hz1Y+qXddY349UDiy/Tf2YzeUI/FS11AC3RUdmiH0qnTIM14Ve+ta2
25l1KsXn/e7GdvoPhgZdJ1fUYkMEEt1SXjE6myyYzjQwl1OJQtMIzqicVSDL
KDKh/WMGP1pp4tIjS8aSJ6KKid7NSRMUSIjJIOaMA0tMcSA1988kXux+q8Pz
CSdwaflWfBOxlOgZK18I6kjT7Qujdg0koKDqDaGslMP2UKHd9t3oOtemxZ0k
6qn0s5fpx4k3eMpuNU6PNcQF2mdcg/cIWyKbQvykLYIGkhvTOrjIQ1CxfLyK
V+jX3Ia8hiMOkHuYR00+B2EGoGoHxpXNSNiMOcZ77Q4VmTqWmtBwfS+Mt69h
XZ7yex9kwTkOZYIWbqS5KcIJc16kmf8a+QQqZRyfg3h/vymNMl4/tDuZq02M
PeqgGaYyOOOsx9tiZ9HjCN/Mxww0pJrCuwOgKmPDVQ0FgNbs3UZ8dAug/SnA
gU49mtwifeGVmYcDtlPYH0mkS4NZWohhQe0eSR1DR+bDH1zKuxLARnP6cpdp
QR2ydvYo4+62MH6syRipMPt15Omd8QQL+Xbqf7jWQz8RpZInsIfT/ebzdcD+
LVRIZrq8UBDzKTfeUQ8AtlxdFY4ieLxQKTOt0UXLDVn//Hu2bHh/A0QM4GWT
xGNz2SRb56WnCamQL03u/uRHkouxW0hDZq/pO38bkQjzF0DR8+Bhtx7EOcM8
3CDo80Akx3X5dcGSZMbjDiK/xwPQ8bn3K3nGFwAXy+xtipHOs1uZiAiwIv08
0qy1OvcUZwwlfUFjoB98h0WaedRosQkcwTApcJ+c175VS4XA1pxlFjJc4g/0
58kPfgd95Q0NyszSf6ow8ZqMRRftLtbkcCi5La4/8LTDwtCIZ/eXYHGD6Rna
Pz0M3RdSAemoiQNz3+vHRc6JBDbgYOoZafJ+Imnok37mqbGj7wmBBfmYew3Y
Qaaqw7eWtCMKo6zrOgWVRMrT9A1cFDcPFckhKWAwbh6EBwQjkmQ4vGsrI6/c
CSj40Pr3UNHIsTFZ6lvbKgq8EJAyaHpPh0tYJKIGG5USVPIwRW3QvmqGnrhS
hlBuA4bGGikzu8lRBYAeOMCmbdgwsmRXWwquGnxyr2ubQ9QUK+3+RqWX5Cqs
OB2OlL3yfvHFcLe5V7u7CiMpIJa0POXAkJHXUyDPbtOUKuodI27wd1pcB0nP
AIMFXjrEnR+oOP63qjGgDZl9cI6DMS0TuoRJGLVWPl6P4J93qvdMCSvQ6RHm
QV06IErGGJjI8ImzAvvTJYAiwtg9pfArrkjuXoDM2OOyX/d+9mb8YJhUl3Fb
Ld6gFNf5m9sYCVGnrqd6NDHEc0qnqslt3WZifBKhRYOkgWMkjaf+ofR17X1X
6ymu7x93gzy+b4af8ui2iCqWvPlxpUF+vo8K6ppBtZsJ94/4/bFKRZAc1HbX
+vQ6aroz0AbHZGEnUSHJUUkkNWXSwhlz5wNk+VQ7wgLYbmImM9EHQr8Ui8Z9
8cPhXWdZy3MjEdznWzGwaj9l4r8C8hBC0dcWrRoGK4eMdxRqtaTadjQLR4A5
nGu5QTDSxNGPwqB+hN+i2DKBZUGzqqH2h45e/7inPs05IvMEsgnyNvyLkWWL
udflw4D4JcfsxcFJU1oW0Qvt2sc8FzKEr8pjVXlivqjOqu3Q+GRDa+6i+0Dg
rX88JQHVJmv4MVvYzhnOXoU8Cec+84fmLUTXp/jDqDwqmL1NLG2tos3bTIkB
bYK0D6UjoaryOCJ9ugGmiHVy8Y87d27wbch3t7fwVViwIkCuznj1Yiyy5Rmp
fVNxlspDAeVRup60Tow7FJgDKitOdw6m5vTowFmpQus4qME3kE692rE00apg
QvdJ4tQh/zqVfySqSyq20lppzT2teiOSGfVmPnqglGHB6ibvsLeLhyd/+TB4
eAL/wJRDO5hPdqSYvJnoj01tXX/fVWDP5ZJyR+o2pBfVY5mmK2ybD2N3bI4u
KVJqLB0D1eFDNP1N0dsVUdZ0jwIZTKgo38HD5E9e5qLHVY66LoHOCggug4ZA
bvjrmrB05cMGIfUVGrA2IvxUlDCmJCWXeLM+HsJS5yOK3HiIRtA4UJ8Mqv9k
FFFDmz+nf5xQ2Sz6SAeBKPa7afQBy06Jo8gid8e7RKBL2LSUfSBWiXase58k
+rhmyr0y2tdUWfFb7E9U4fCLUlkUWKQulb8aaTFagSOhWT1vo9TTcIkZzOLi
lQ4SNfwZxzySRI1HcQDre9/7ZLD1muRY7x3Ixj6A2cDV5BWLGVuMOyncptQb
K6oF46DvjZTPnY/2hSPtFFYr4ihJVE597FDOshzkjKWHK+171+PhjfZrVrXQ
6+dNRzjIxdgjzgPBksccsc+Wba+mJBlFefh9iGuQ43r75Ldg1OnG3piz+cIZ
aZ36nIHQhaMP62fvr6Dom7N9LcNFy8o569S2KIzfKIlwv/L3QwWn0loJzC+n
G3eNsMmoIVN6iiu7gpB8RFZeYUvtMbDhq8nAS+mmigDcGI2F1TyGd7WX/8UX
ErKMKjcOPa/Cyx7nQ6UBz/Ug2HLJtoFGC7wsWqt3VilV/ZPfaaLCULRmalV6
yIkyRmALQ5aTesJ/WVOXff9bszyZK1Ry49wWVO857RELwfuNIt97i7426LgP
rq1mzzUN9XsR7ejT4pfKh3fYUiJLeoSnKrl3q8fjri07ZoXZLz63ic4euigf
So4Sd1toFTJP2UUxhCn/I4BhEBHtc8gRP9zKwXr+cCY7WeVg186vZ+p0DCEU
KGsGNMj+5gpt4RMiyncNPEmpkJXOTHmfln63982Dgp4SOe+NKn0fjPrzBH4N
NEFhRCOLFtYgxl6hKsvnFDFYldqxphuyBsWZCgCcmv6Vel8W5snMiLXZaktd
G+2jgi8zuDP/xfeZiOoSKHQ6iwLEqWWI1C9AXinWAQ5pP+xAotO0hK5sTcgH
uOj82dNBtaBxwRCYuzx+3ijKCC4dsJzsxSLU7qANH9RV98hJ5YIL6iMqEE3m
LJHmQ4xasiQ9eNy5SM0I95obKyIhGLBsgJacQnETDsFW8HrxL646mPkFTdYw
QQxkMqJYdieDcyJqfSnTvIm+lVIdcFpW8y4vWOMm1Ylm386qaL5O+x5YuYEe
vPTDHCMIAS9r0fUiFcmdmqKfhaXGo9miI0zm/yvkLGYG2p2QXQmJkTuGW4QN
yRdES7Y5WHRUSQw83VRGFVOPzHusnfWBzwQW68sZH+rUpDpCZ7PDkPpsWKGu
zBAkFR3tcUwl6GW3AujwxObKe5Xz8hqaTq3uoAS8T4IHeMtaxh9OkI3b12k6
FH9cagVBq1rL0gNmUARmSjBvDZGRsygvLUvZYuMCboTfjtkNYahX04TZco16
Pnd2pJiPDOPGXGHs+RiEiWFjGzwv4Qzeb2oIE50ZzejRqlagmypS/VeIo+oK
CPTUFTE6x4LDNPmNRZINtEpnjzkapELGbuVQvJ/pnWTrHO91nMNH/+soW3hG
Ix/bDj6HZAD32pTdOSD1hvwQsabxIj2bRLjqrudgJRD6GS3S3T2dN0peCEaN
L8HVIxtz4AWOEvHhvasUUMSuqoXleBq3lEN17sEmpwz8752kXILJ5SHB1Ry8
tH0S4yqWV4vLfj/o9vOwZP5w0f5wPbH+lsUaRB0AZBR9mepxiNtteGcteoj0
HPAjg+BlECqE4O+zDuElq52UkAZQ2aiQa3M4MlWc/MGbh/Q4Ty1NY952LIrQ
cZ9kmtWv3XXiTffdf/QYeKkWjjqzdPnQWx6sHfpaFgIaDN+nfEq1Ru+2LKag
QGOTuPgfC7G8P+EiNXbZhO2RawPgdt/X2YNWSfubS242GHozZ1KKtdo7BmLX
vVFhrfgKknwoDoojNfd6xGAN4EA0rsmt5xEB2ljRrid+BHD0uhLDljTb/bfX
3KeY5qjwsWuEmyytUKrR1OqOtk1/+EIFynVnD43ApRt74OLLCj1ICWTPxbf4
FE9uCQwN4pvJjPRhIi6Zg66MawI/iv03Vy2MvH3Oea21RsKKAao281JsPudp
UxanhPop5XzkWHqJKVtN3UxpxYZDGirg0BEaxYcNttryPDUB9BgHg5j7zAJI
mzai391o9285hKG7vrZDHKPD3UVd0pioSUGaR1qEutSYzpgJlRJUFbmH2e4o
hYf563KQ/mXSKU8BkejLlhcWAqbuY9DGgJCbF2mpwiYGUtON7eVBc8ecNxqZ
ktLDQL6Skxib8WVgYE6NBcDeja0+2ZQw6MPb8gsIZsWgg9NjtGFnTK1XO4H9
n0H1MTkdzVZbHWa2RVW6eobrqoukDOS6zbJoxyVbnu4oZZpValPkLaJ6X0fu
Q2z4NE0h6GWOQxFVzePmSqxGB8KOC8DSql+anBx4lE2noGRgugL38MyHwTLT
VVYRBTEVxHGfGUMQ17SSE1okUmLI9HP5WclJ2sw1/dVeGAGzC67FMBot6p4I
mf+gWF2dca/NcWlvCduUFCMlc1fBhJTtiSYMJaRqc4z5aorkI/NCMKWbSdDY
U8yubmYEbXslqwhnVh1XbYowzJXZs11+hjnFbjGWuDoiylg5g7hi1QRTLGN6
on8vQpUitni+GFeY1lsUPo2Os2quTULO06jZgBsdZF5vNH+vQDfDNED81uwl
G6p87NPekKEPHrf0hgiTeoYSs2Hw+TL0sKu6urvUT1kg/RW2ne+0kZ9cukGr
OzKsSBpr0uGIhgqEo5rvSWOcxPdnsnHM1jJNO4MvQU1sRs0prDSj0zldA7Q4
1riE8gJkC4OLJ5/U+/9Q+LAu/s1h9dUtGsOOYZC04vML3lHgdcltTpE7KV9j
BgK1DqDZfACVwxW3+WI9gOpwMZR2YF+XtB2IT7HL+6nfYOcP/lXFo2CEUGW+
dF2b1st4ERF1nDir6g1+aquLnuKhb5nKL0gkCx1a+k9z526DzathKvBTxTNk
hFNjKkxcfPrd+TuMak6YlR7WKGDGVvFHffXbePx3MyBkrP0G3/EXbmmWABKh
pt8XpChZMJENGyOGZZOq/Hterbwug9WMNAlPq/6nLRZqFNIm5lHrjcGL8Gxc
tdlQ83QQ8UMmB7maBg4i2MJlk+5pHs0DxBxcBQCx8WT3+/r/fa0yIzcnOrVl
vCKIB4nZTF9U1zSHGuQFZ0qPyn0i7BQ0iZPjuUXZaXqDsI1pkNoh0+z6JVDE
gOIhPfD6093wKRiR7nhc7BUoh59221IPr60Ml1NQgu1b9hFCb0haNwPHq9Rk
rP4l/Pfpic3lpXJEdNAWzLGNZX/ywfzzAK8one07IKcUs1KdtpAvymliXD6B
fuM7qCA7la0cZXVPnxVY3CLX8D97d2gqLjN+C5vZYIvZItgOS4F0AmUK3QO/
TzgTl8Jyod1ZOYP7RsRR26SKmZIL5++EzhwDJrBqMpBzw8qc2VEPRJ8huc7i
v+V7ysbv2hqHwFvk/6xxj91XmBH0sDlJA0TrfxTbOJXM73aOCO6UIAjEIl27
tTNFIlx0+4r1O7zQSMm9/M4yjmmeDI7NTqKbquT4iIfR/oSas09rPBmUz/Aj
0+jofnCw9zAK7kzGN5cuIko/n78/Qn3BeGHqtRKcfAy5ibQ+0PDhO6eO+x4n
ugpV8clU9h8fn65lSNwawZ0TRVGO7NWkrW6xmrtdVgUXAQLumzIcLXbxowjM
7HUFRYssotbkOHtCe8FHeqpvgKfgJCPzSKq0i+abE5KZmHBOmbVkyQOXlrTf
uMuYbnh8TW/8LEEMM/lEknsCaOFgLTpxVmwEZJ6O8KiAgtPXYEDLNtuzhCe3
XpDlxY/GN+DrDJJSxoIo0mmLjA5Fajek5d7A8dcCk8BHzJwmsYPCGe8Q5l/9
Oc4NFk7yjqZIyHB8Y0k4ZB0aKxEz3zZWgv6yp9zQetJbrVOOm37Anko4Mpzc
PJKvbubu1l45bUcK+uWcVdKELmUgMreRWhwj7Y18RptMUwwgiy8Kvy4zbP4q
QUSHWy3cEL46BgqZajJquCV28jJ7q2sgvJkC/Z+zzpLQDMF6mFXavvG3cwTx
4bTqdAwgXlv1Otv+X/srthuh3CC3hUl4OvSJnGehKSBWiGIQr/CATOlSSYyC
vZgZOm+GdxkBarMNUXskC3lTvbDrfyQOGiW8AId0FKYdMAobVJxtuMqXCaZL
qvx6QJcN1Fo+cXrMteDKPywzj2ljDAulYSx0M3dqICYHAE/jw/P72U0EC6iN
RiDd/YdL9/sOEgm7cGguPbA2CvRaGNqyyarYs5NnXrSyCdgUrVh+uhDC9ch2
01iNtbvyB98RYQyxDHSOWWDLwZx3UJWqeHBgOO2jClPFGQzxWe5kzEIzN48p
8/Q4QQCo5BME+OtW/HzlueZnZYKlNoe2MSewH+QZeVBPJGHe0ax/j6CN8p8G
mBnBHQclkUciZUcmedGZKAV/Sg0WEEbNrNZfojC5oH50yfb5EsTSY3/Ho3cn
k88b7ACsSb10g+WsblT/QLzCfBecrKMXu2JFg8y3K2H9x1DerlPqTUrtpUfB
2Z+ApJB/npVVxtqoN1LDF0KcxegqWIPYyBe65YPnPkPrkay/kG8wr+v3VTES
PU0Mhi+sCMBxQpdZ3LJgyoAnMC3jOlGFU0URRzGpv4ttV8Y4rdtApKOoHiBg
6/jGqx1v2+K6MzvDx6L0IUQQJG6ce6bycpoT/Fa9f1a31utKqlRD8czQn5N2
R4iZzDe/C4m38H4OghsT0d0I6MX8Fqgs4jUVwHDB79ywjVOi0gZzD1jVp3Is
WcePZCm97utdQvp/UVMtSgosO6/2+AEqY37k/BXEpTMxw32cpIWJqxWHZl9P
8GYYwhmStRDJ+YOrw897rRSjmDVL4lbL/nqG846X/ga9xIU3zqqQPahCNk3D
c4+QJEHGB+ufM4oLw4PuMdgYu0gDcibUy66/VPv7CzgpPQkQi+xqRztEP+/Q
Om/MlLn6+vta8eopZqL26qpy8n5O7VPMAG+kFhvslHqw/zFZauHQoAHY1NT8
9U5DC1rk+vZSEYSxqwLeEZ64ykSUBD775NCYHCl4lkGiohPbK2kwOp5OvUR8
laAGNA5hFyUsycPZZ9bqgsHI9ulA9ld9yRfWHzjFmS8689fvM/DVsMQ+PiX8
zxSqMMRVC0KYRxPl/oXnDjt+XbY2Cd7ud//8XMfWz/lyQdWW22/8P6G2G+N5
qSmbsZ/JCRD8L3WAhBJkwIiC+9+CetgGHlmhOURul4FmrCCTThSyvEscow3i
sAN8viJsGcVdaymOcrSmq2gWPA6k1nH31oiH2WbTOtiosyLWqvEpDhNZJe/K
dA6YKghcqPB0sIXYhjmbp2OgJHmnU8JgRwlB/0XSNeMy/2N5aN97B6D3Vs9Q
j4HCo7r53Sj0Xc6u8giy/KBklRO8OBCSAxJsg3a5iwCq+CWfcp5Z8PXofZ56
ITa1dYiwnLWxvGaLyj39IHGzqYrSS4Kuh0/oFzxxgmEgkN4R3lcWgAdtg3by
PNu6nqUU638/aQXk6jL7+B6uPCxL/ep20pce9poklViK4hdMYvQaQRbQWCWf
j0D1IRwgigPqcRMBZXj6iMVp4oik8MD3af9RGGlPNGRF8JwtZONG7W3tY7JX
qHdzlIUwCAE19Zs/wuFpMeJnf7xVk+l4IOiA8RqtO/4fl84PaiK7atzpVkyD
VFnkMDT83TEbZaKuwcD3XMsa/nFd/hizs+gbrnrLv3cYGYEO9Pcvtwz8BeaA
AKqnJkfnqFOYnwHy5YXemzYhJ+3MVXjFH1Lo5rUmZ0uQZW65dj1/0rgerVfl
DU5CcgfENiNOYlB0QpmdcrcZbdl+KyClPo4Xuy5QPjCHwLH8WlD9bWMlIsTF
YsJ3xMeBx8wPQsueXbs/Xbse5/wPuOZN/FP0af5OAnm7pVyP4zAgT/6ZPTtT
e5g9kIrvX7V+dOYTu0x28SfJPQX4CDlswkyM0tqYTQ9bJZh7o0+QJrMl3H4W
ZBP4FM+YBkgKVQf8XXNXNeN5yc2uQVa1F2zSFZTzcAXAK1FHtIpywEmq3lLu
4CfyiTJ7QdDZhaqochn7F49/+xzshrWAXmyRVU5YGNypXkZ9WUcQDyw77PFz
itJ5JVCnEzs3uiGuXWSgOsP5mcAy4v/kqntjNJWvIY/+6AHf2S/OaMinGZ81
p5zzuJGcpf14GOq9EHgXNhXgLm8GUv6W3ZtCYvDtEDN1SVZtzWQlsEW1If68
o4ozwD9fPmSUY2MzPxUSGrJ66BceEj8v/39P9Hx5PevoqdaMy/wPpTiz2nGk
DJIItD4Qvnanqxm79skSNFSMlhji6yqoe0s8WElKoEj14BFWdQuIDRELjvgd
wvIja05ts/3BGAALqrPX+Ml8tFMZWxjIu5bzWvtqLMpTeOOjDrOx4o9pBc7l
YpCnbg8AITLIAkyEYVs9wgtXX2qAP7jYo4Eloqq2aXxS2AiKP/RSg5/4aUpk
bOvmjwIZCR+IYXUepK2k/2o996prDxSuG/mbqZsjm+V/f3eWAKf1zXvj1KnJ
Pf+qK326vgkglFTJ2/OpE4Y2wlsaBH5vQksQrWeEqyNNAXNU33Clb9xEQGDE
Ku3G/WApIfpCNL2pjREIgwu7KAf2nZq4xsQrkjOcCagBSsJRAmo2DSJjAG6N
k128T8kS/3ABYwTOcECzSe4Ni1kiqEO/T4zlVTkewO66TCkCAriOZGBlMZ99
DI5mdi1jtqjUxHfkgPWdp5n9oPc8A8oCctTuFND6u9xpnwI2PkSapoHYSdSg
Fce7lBCwHxnsSyA02pMIyDL0JXWYNTlws6LUIEWKnx8CZJRTUGhT1NaI/jaT
cYnS0vi6tS7I0lNAYI+s+CS+9fr09BnILSxHoXc/XsVjXse4gC+UpNbKtiC4
UuWOmLfflpW2QfCEPRo9HFiv7+4WojpDAHhHGKLh088VujCuuS1go/qskvPL
2IN/CMgc823ErrOAdWJ582p5UxD+qSVPuyWRwFU4SGyIYSVmw2MVk1odb2d4
tOab7O/nTzKQNvm3vnxZ21b2JFjpRsBfHxPMBvyE6NntKUCc+OYYq9BT2vni
5pAUVi4fyuRXTTJJUaZHM4kg59AtCdJqJTTJ3/wOSv6J7AjTGilEnroXFjK6
896GolLh/eW6WfLUQZMPU+xMHc4PJJZExeZznhLAJt2UBvYQ4owZ0KP0ysnu
nKzAvUTzosQ8RayTtVMiMx1GAv2oMGROb+oeZn1rRUsqIoctVwig56bjZjm9
liP5LBn0BvWwkAqzKgXDAoVgp8/szbRETywhynfsTRmXDHhqo9Wg+sM6bS8S
WtwOIg+/mCd8Hp5eMhlTGZ6qpGm4KE8zm7cAlQVhZZjXnaUI0NwMbv6LkxEf
3C/8WxAHqfGthMA3qszbi6dmle3XeUugGBghBQTj37vKJG9e9hs8KG2iWhK5
3COVn2QZgKx4o1Q1orcO31M7ll+RwMzcd9WAXd8RzRoj5gxjlHN/SrpjSQSK
6nO/ROwktnLG6Hpu891YhZwXA84D8RReqqHFx82G7F5mKkiJcEwhQ3Ni6elx
Jn1dkReHtbonKgKznxDfuzFwmYtPlaHq4fTDnyWXUE79y/Fp5sIfRwgxMyOB
VWXWanW+V2Xojyty30rvedtkMHVLOfBBU10bibAb4TpiWs+JW3ZErkCHGwq/
iq9MqfQEifgAC/91RoEwPd9KkF+Bz/XDB3N28x0FcljIMbrHj0Ph+2jYbhwT
ckOFXAs6RyNHDLYx/VGHVswivV5ogRFgh0SbNaODA5TJnEABQUCoqrxqMlFm
GM/I2mV/7/XsbFWo2eS1gblRGnIBosFEnQCTJTF8TmRvwcW6Yph6WraltrKZ
JYmN8oUUFXQfxAOmyH3mQV9bu3rHkmK1b1ZM/Ykxhk/1iMe5KcjaqSVVQcSo
UOf3C9gEn+QAJkVD2AKBRuINGEAvL8YjKwES0yjz/Eb/YBhrVauEoP8BpRm5
PCvhwbr4kAOW505LzA/ymnEVvuW3TsqH2Ao+IXSmtxf3YhTOlCckjiPkNVN3
8yikk7JenOcSeocOb0e016tLqWbD4VBCRKWnwxHkw1242jeb/REoZXkdUWHH
814QjVq0ZZd7Mp2cYTEos2nyT5qRDxu0JJXlg56HIO0q64eMP4V7N23vt2gx
37Q+uPdqCfE4uUaGbFrrVoft9bNRl/8audPTg8F68dC4+8Hra5spZhNwdwcn
pnqsIpY5uCxeF/1W+OP3AMzee/+1/LiuiAT7HoO3TIkAHnDhBkk3lToQ8prd
fteSXCHx3/NT2HD2wLo2FcKK2NWN4tyWkHnNisq1rqtZQ+D5YGHJBQnXe0Fa
dYTHLsyMKNb7VNQTBSAVcM52XMHxioqa1VcqdAdqgEDg84nL1n4Oc4oot+U2
nMx8xtC4NNhtDGKu+1SUqYgVtpBP9oE76q+naPavEhNk4z8KViOU4LERK1uF
onaHVnEt+wtsZTxGImchFj7dLxhBkEQdSyPxbGIxABA2CRHtRY7f9W9fW0b+
BtZzw/1XMqOIZu6pwWTQfTowaFEGA1vB6csDsPMlQ1rcW0PWyQ5g822wnzqJ
S+CLdoxj7RKxB4sfzzaKLeK05d9JQTAOjSpNX7Ih5FG+CMmQ/NiRT2hT5SH5
zGykEZrSa8MRYXTG79DAj77Hvs08CcuF9uA+FmmFcK0sdhKtQ1umJG6ZTdwc
9AmWHJrM7qJL/Ou8blS6ADxOklJ20eouu18oqMFCaXBIqs9LoaTEkufyazlk
78abF0aZXStkQWXo6xTWNg2nIc2a4HSsPYDPJpdWkhNH1Z3DlRqmU1VOsvaM
Df8NJ1DgNKLSbm+rjuJYwHFj1rAH2/08u4b4fT7bB/pW3JrLduhxjxC+VjSJ
b8i11CZsJ+kN9Ioo0vnqxXvoEamc+70+PxnfwTP/aDmab9gASinNVZd/Tj0H
orRU8ys8MZEfodxVuX1BoSo3JPN1ti3xgkqrVmK+o0Q35rHVL4+2IMDLfZLQ
QlNxYZNfgYh78algzatyyw8b0k7MmCFUZtolhSeUW64qapZ2hlC9ejYNmNM1
MARsdALRpRRLe6eSI3pBnjY9MLOckzTVX9iXMqr6iuYLqgtQFF+sz3QYJSf5
NLCwPX6y0FJm9zBWnH/g0JaBa6MOvpHEh4h2KnxNqd+VpmuLQnBv1g3wzkr/
RMB5txr7bclxKOH2tYPl443okNOMRESSNM7TMGXnOe3PzrhlvJvXHb7Lk3q0
nhAa+FK/dmKMQ6UbNG9C39YQWBP9hJjAo2pa5zJ+bFOGEb5Gvw6ja/gBWaVe
piOwdpBfMLyiLRBZ+y5dLkuWLjZIffIXuCw7nrP+q1/HC5NpoZrdwmm9qSEy
ko2aF9244uchgv+JT84GRvpB6GZl0Isdmkf8al/JNNNI8Y9k8txCTU1PapYq
XMF/DhqncM3JlZt0HJ9aCis8vUXxTlqOYfWnN1d8geaB/lbYDIMtkzivil8X
5cpeSxtJ+ODb7uRRDEf3bwjWV86kOE7ckAYDvAnBkicvZN7fAoaHfOXC2TC8
6/tjyWFVXLxLi5Yo09/Ratmt83UH9TY8zfgBHN9GsotoqpglUs04aX7x8hOs
5OIYeCrVsERevE3IenwN3Itn22QmvGXoexMR6BxWphDLm53DRm2NTHsdnztP
nARGmVWcZyJ9xPqji4Uxuif9u2D+cmCMrgLGUezJ0sai544Dki+X4IsitkzZ
T6WVydJNidBqcs33EYuVlaec4gPKusnw0z87kcvgqWob14pnnHXqTtsd7x1M
WnF3XrXH58wm1UEQnAprRYK0tzKYnHC1jE2F/FHEs8Qu4nC+gdInLnjavSQA
l5Jc2c+X0KD6qL+IiRpX7IToQNym9G/4NJCvpE4qAd8GXpj/8HPr6SfUTZgv
z/JRdkhHGyJ97q3wgdjoekvY3qzw/TH6Uf0qONIBcC+XUAyUmmKq6HqP5+xp
gPWkAHWTJm9jXB+ALGM4POWlJvY50nSFwxB4eH3czjSHhgGrLdp7m5L0tKlS
jf9pb1k52qJkjYSFclPOFE1vZlT4Go5xPzEhSk4TX/GcmhDqIjTrqP3hfwCd
A59MBTaUkqOAjup3K8x+DxIJRnC9QGD3ovE93cUykwFZLaEZMs8pgFxcg1ja
OjUA79GdLE6Zzm/tsBeptF2KtQCOHsIRrudcD70foiY1ipBH1TODuO7ZW/Ax
oJAJNo7JsRXLbAyvyvLbd9QtVMNo35iNCRXxgfyDtbyw9UIlTrHrLR59d/9I
AISGYoN1/9lOdU4taGKGgw3F5KQu1GYxRGQJ3aI/maPX30UXhBQqLiPT0js8
mBXbZNXMOuDwN6yXw5QMxsxn/V5QcJnWZhUpYkMgyVlqF6kpgGCvZh8Vh7gY
9YT+sT+aE/3uwVzRrS4nCe7NUAV6MNAgEk8pxT2LWdrRnaG5Oqq+ckh/XJDl
Zi5V6a3oR9963mv7eDF40NkGYKxOUra9UZbn4W8gAGJ9NkST4yts0Wo1ViNc
uAFKgaEgPFmkzwZzCTKVfHojKVQ5EbIasAftbBJLsYABdtnQz0ZmDYwSGSU3
SaDikfs76uPeyKoiI/zstrOc79zZsDr5V49mJt4ka5/TqEAs1baWXJcxVpMX
2uE3hXWXV6koI7i9AxYM6g0bCX9UHDwKF9x78aw2dUzQB81Hfq4ecZFi11Ex
HtM03YPVv9wCeMc0CbCC8U9nrlPm97NA1FAz7wJnqloyhBKL2l/So9ZwR7MR
0E9RJ1o9ubYz2xS/mRJqA2cahO+ZGoVJloRsf/gkGXVhlM1s+/5LiauLTD2I
8C+FO9UY70f5t760yHXfr58LeZOWaFvD7fRn/bireG3TW249z1kr1Ff2VrwX
PB8qU+ElL1FVrfR2ENOrGHON+1zwuHofr8IKbGEC+vBUkG8ZnCyO6IOhvLl3
XQ0H8oxDmTAEpvOFrMXdrmWPjceuUP+NsDU/rtj7y7LA7P6aqGgfUmT6YyB8
JVYZnklE3dcRJehtQ2og+bS7KvLXLPtP+HZDENmfbQwy3v/z6n5iNmx5obns
DV30gNNF5whPDSBRJha+aVKDS1EUBnYN4iN1rRWIvFNTVAbxkrXxXTBja/Qq
LeWcX/sE//E+LoGSUI3M4R/iI9ZJFejyr0O+id3MoiVCXAHbSXF50wgssR8H
gVMNSy3OrLlEGCuWbK+1Uz5595prpuoWz6BrlyXP1FB7qM1QM2/bnmVJUIHq
J46FnvSWato+yoGJNk5faVbMrGXdZhj9IpmizvTcenQ8f9Trp0y/dHrOh7nk
z6VtjPOBh3IzanR3vbN8wc47eI7sqnZZGx1WtS9Ts7hjzKX2YnrAgnYnDhBw
6B3hXPJiO+RaIXOwgevEYgKa8Bog1tP2XJ1yFN2N4RmPqMZUG77xjuKTDRrW
2XbkR6PHvPKA4TzssdLi23lIz5+n/4XoIBDLwW0Lj3P4cbjt+9SKUwOcM6CP
R+zJkdBcQi346iK7AhuayoyfoJwR4ipZDI2UzLDjMojAyh0iBKnA10r+Ndo2
AJDlSxoWJ9SZIT3/BBJamgRO/xD7m1DaYfSHvMd779jkGh8DPgRChYq8BllT
Sp1H1dtjw44tv5keoiSGA9nr61pPKjjxnCeEEMYUynUxEiRMguDL/EyP//6M
/+miJ7bUjHUYjdROWOiPoSSmdvlAVFk7GsjeLmOL8si8r5Fu8ioxAOVjp9qI
sHP0qPEm5L8CO+5Log0weddIuY9ZNympGlTmTyUF5khWkQ++vvH2dm6Qn12q
22nhxpYP8D8MqbzohBUPZmci/xla8S3hWbBn1CqIKIDDVAtibHFoPGGlsM26
fnXx+dj99T72mi+QtX+Qu/qumeVf4FkpTq853qP9qZth/cmcIMX/NrPJZD96
jR2yVHC4dIKAYhGkQbOgzXW2q8gWhIX7n5Ucrug0tWtyLKTS8MMH80w/n+zf
vKkxF/2/HDgYbqtat1riHtqbIEn6d8e5eJlZDUZXZR8cXkX4jQiXgalrqy3p
bHRoPSCAmSfoYWwQ3c7TrrZvF+NzO/XHZlNZ+p/wwew5oVeUuKso8HkVSVIi
03p6JIupGsoXTwYqWkqMeyDuyvtxclVMMF6qiTSPzowWRexzqymM09JPbfKW
6CyaxAifYxtZhkiwv/TrmmF/5yOp0XOydGINFyH/kbLcNxs2AQcwBrhn67EH
hutbzW0qGuLvfMW/D/vMsZicnOEYYXhRyPJ0ejT0pTLfRijbfziAvnGUykC9
ePZEQV+OYgKyitemvM9sLnvJD1L+jaBhRuKiJ8QYYEgPoV1rdS9iwU7UcGpg
amxy6HCozaVR8oDVrdNBcAaecBb05sb+NgE7qslzYiA+QkXmzaOlZrSW0vZK
U2DEeA5foCFafvNZiEMRB/r7kKugJUyCmLknu+qtQ/v3QFksFgvDDcuxENIY
jrrYtl5/H+ehBzYFw8xydp0Sky/cVOPDsfLIbV83IBZaosrMCE6JOsRJpEfK
qpQMOVno9ns3GwqPCkve1OiD8FmIcfzzC57IUO4/h3c2Un66/XpW4CIIG/ob
7KTZNIOL/sbIJZf1tH7Jj28R4O8UpKkT4FDcrIBCsxw1Ms+Gjx96WXCqt96R
hsB7ecB3ZRQIc1jo9Mbgy5NUHydt1Aztp5JRKcqZkkuBjEuQ/PDh2xetHrF1
EpGmRz8wYURzj+GO0YpKt4AKDfDh53yQ+oRmAmpyNUGWODV3ANsbit+wevgK
mNWNjRYfqYvgLExhu2M4PXwNkctni0tWAN4zq6qVWQLNzebXzXMNLRiOCfdg
8Ua8BnZpYCBqTeLkh0tOXbOiT+0SOL+JXtENm34OX6RXuPBBcxcg9+ryGMUZ
wqm9czuPBSVgifaHPZYTsBY35a6l2xZaO39RQsSCFLm7CMSQoOOCCvf2gK/y
NfpqXOtZTLlVyuuKLoC8ZLWqTBAkB+ijyVSX9NYRCbw/LFDtZqDuEwAieUvr
kmClY5DA7Z4hDaJjSbw7TJhLqIsVYIu5d0/37ovx+3jwOfekmnIkwekQ+XXo
piND0E/Zmirk3MQkx/Bvn3Qnleh5CzB00EsjPrc7vmOGPfQtyfaki96zD1av
lIZoMaDAQ/EhJF76MA49po4CAxbjqR2jYA6M4LxdbS9iYszgNR2mROtQpTp2
Vgmfd2P42B/WnLaHwNazXGp8FbfT5311OShh9EeNzhXSqr+O3ZSnzd42mqCe
qZj6p0Nau8BE7TVluHC4rZK56T4qDdJ6NvrxGKdujX2oXSjGJd2lc2XdC2CX
rUZvY/57CngIWQTTr216/Hw05/A4zEJn1PBTwDySBc82CDrjxq6w43jOv5I5
3RokZjkkZ4y49tMYoEkYH8j/rBcT2QupSAjtKRgSm8tkLSfaBJK4e3bweg5C
W3WpLy91t4/eg9AyKnw3OivgEYTmqq+ZYHbN6ZhNZi0ApIUemovPuJZ1SCOs
/dAdBAoxsaz2Aq6aAAFt4XaCjQU//JLYhJkzG4OhtYAhSc7Wo46BB9zkWa6s
quvwDxfEqRJ0yQsNOSpJDddfKB3ebiWCl79EsUuTFGZnje1p+4hbcESigBV9
4S2tPYZ9/H76ZLK764WoZd1zvnt2eT7crfWPUp+kvraRZIUo1ItkF1JeWLbE
/miuKzILJHqT6bhQEaBdtVcSQbn8Oyu+1hjiR2uDkcuNeNGUiZxy9M2h7buM
NMjkDbOEqM1rDjPIFcfAaOH4CEx4iPV48WKpURYXFIT2fWTAmGz6wqmmlJ3Z
qtIw3MhDDKk7vxosd+qUXPMvqFe2q5tLjASy0GpkcWbMgjN1GN1972eQB3rQ
wTpOY3hk/fVkTqVroB0MrtoFuoxg1wg4qkEQow6iX55VoRTwIKtvUPTyY864
7YsypsqNcI/yXFzCZ9YZ9vyAdMHGgWA8zv0HYYibtI+ldV6GSG/9RDeDqgV9
Lv+0A7x1zjIRJE3+KQL2O0b9k7Hem5O7I2Sz34REinf70R20JrEyv82AJprm
NKpLN/XjstycfI1W1aqDzrfLMvsISfXjA+gDX68ixyDH4STmPiD5qvofLtw8
Q3ZDkg3WkRl2xrbvnp9k05oswV12K+H2HfYVdXBU6VQwhBl4urPtpBG5+14g
C+jtiXUrl2tmIsCpTto0w4sZb2kFDrEROlLYvekch7Z4Zg34bE1yRxDH3lgo
zHrYXn1rN7D7UxQ6U5akw06VTJ7+TQQC4vrRHfC20KYJ09L8ShiH7ksyBW9C
oz6Th3PUcClnrErbkjBTe0LriDuS3W+rV7VjcZxDFHyo2tdaD8IzEj+jFZ/X
+1yzPUsqMYJHig6R4xuB5QNhrDBXr+lJp23lnnaSOdj2qDBwqAlju27nSou9
5sHlOY3+dW3V1ZNKYgfznSnQnWzgrmEHZd9TfsROqYbvcZne0n/OWeBGybpf
iw966HZEdeoEo9x1Mf/KByRpUsn1ZOfje5tT8LJOhcZXVuZvd2chZMQ7OQcI
8Z55kZv9u5bM/7xbAqcxDedqN2ryaZR0zOnaVytXtb7M0iFLMVgRiJg3qihs
xSKhdcwmM9+iyc8UxhsIFk60NePcmclc1RMrVePys+r2vrWvUFHxcvZt/iTn
ljR0NkAT8fmjuo6kSOHJo4yBsvoK3UMIlPm8RawTIEWDREGmOQ/Ekhm1DO+3
zYOWr9R1YIviIGFRxSxBAVcHOMwfA268G49YcuSiGm40bsQ+Kv5ArStSpkOJ
AK60bCmVhL2cczDyMzRAC0B2EH1RSC25bA43tqgCOo+1dr28PDG3Uj6m7tVs
ysMmkUw9DnqTvVjFV/QJTqylqyexDbmC48ZM5bbjAsfdVb5Qz/b5Mp2ai3eI
LUVugiWXnnTXmA3wYe2bUXcgG/4gXP0zUhD9XDWCYXWSvpQfIB1Tk7jaPpI1
Nq6+UG9XvKQro17RHHFxSb1GuhnFodoaRgLtA9yi/8yeb1QffS4MLuq99H8/
0Hq5cT0nW+e7WYCmB1SnjsaAR0svH+/4QX9K4RSsoH4NxhWNg3NFWWhg251K
bUOm+U4ZNnO2dAJkGSgGX1h/NpCLMR2tL7UcWdo/WX7I+80WUrcSm1Mq1dvL
7CKAfZ/O/wYiQQZIPzK7vPyk7vwQQB3HoFTyjyqV/pjPBoIq2A0usl485157
m/GteeqRDybISRbuacXRofM2BFoPYzSEr0bVpbVI/txiJQ40hMomcfGqFNgP
geYdS1kYzzMKI524y8y8SEG58j7Zk8gEUpTJTvoQZy6sYZC14qHXv3if+uvY
i5vz3KIP76FNZpqWZeqNecE0vIY9NiiwW6BahIXOWLj7mvVKvZ1Bk5n8OS0m
stnnv4shgTwpEC05im9czoHGeeFdgTZcbTL1X9JiAIEg0CkoHsI+LdWXZoYM
VkLhsxxIjVil+i4GPOwIyZ1LEQieGFZokStSHM/Gtn4U5XLP5fLrwqIGdkc4
e6RzJx5W70x0D11VQmm08mirsgVlPzYolNkbNmE9feEoongkuKhUV4R06+lR
k7wGOQpBvzSw2FZTVo/JrZIDccqA/hgHlkRnCEkwY/J34OGGm2s+mRMXq7TL
YNGNHYz/+JnRS2nI2rFalY+XKfBCMXA37N8ZBJQ5mAUxMIbII8fYOKNRRiPx
8eSNbE6Xs5NjPfxexz/uwHbL7Yk5+GEQVMjLg2aMVBIsr+Yp+ka/K0GY542e
z2cz4UWNAF6odGOgdihv5aPRa6M94kkzuipC/WB5jtNzzPHIkITHgnFdFXcw
RX9lUKkscGHJCJweHyv+nUpHKFMlN3CRBGu5Xs/sWX69w0vnRbV0wQ+2AyDN
pDEN+3SnkSvkv9NaACF6x7GWiKxfnRPNeyNDTakznTQYrXvbp39Qcv5qap6M
JI9R9uD8Y8AY5Tf7pJeyTprUKpjSjT6uxFPLcoGeWO94lqrclXCqkUyqRAXL
N96q8KBtkT+OdeW0HbCm+JI8Fhm1wAcoY71tSwHLw8VQscYyei4UJJDjeEzV
RG7v7B4snTCAUbZ+5dAQybw03cnXw1jNRvSdAutVYInXU7JHUNP2P1JIlKpH
+8+N8mZYI4hvWd/WAmwSW4fTKrk8U3c6/B0tLAMtEdqy2jNJHmdewS/DBs02
/9gZbkfpVvlDun9PBeQm+UveAN05G49vVS4J2hGHhXGlVaiKmqrVdIXX89CX
KD7+H+dvp5wa0Y5gn4GwQ0Dj7rmMReR9ZdJQMNTavLTFZ6Cu3SwGU090L5Ui
OiL0b3d9rNoHsn2gTaeUlLBLOYaYRgNUzYvrcSVw+KsmiWxWEvDJlCEIdzcI
eWLnUi/qBquutxgfz9hj+2pAmF/jsAqsY8i2xfuT/YEYQboxkn4bas2ClnPa
0xNoWnAcd8ysXni1IW8c/RGwiSKMNFU5jikzgygfp3cQokfyYwBHIjjmbZEX
cmpdKXlVDpWU56yg6ITcyPuboRp74cKKuKimgWzcfYPQblrmNqCvteD7L9gy
I88aUum1y4+0up7JHlvHKUZDZY6JtyBKmk5eEx5g38SZ+osr/BW3Cej3o6N4
ThPRaAWySbQz6e6I21Cnvetly1Lxn/qhwCUNaG4/CAiYvA9/MqX6GwMgeqwm
y9ISu299o+P9Hj5SdcphWmfFfIrLGItA0MCTqY0SgizvnT6cqXiNCS+w4Ka3
lGT2ERsrQ26LheYWPokKSOkhbr79hgEv2udYSZdnYw6Yu2QX3PPxlGw1Ee+T
g4j9/I0Ob+xcFbyVjsYB8LuPflcfWNNvZZ6O9I1JxINzVx9gnNEPX8kTeXca
7x0G9U5880Mpeqb1rR6MVQI0vILcTGlXjy+wyXDd1ouNnZiBuWVBqPq+yoex
2O3yOkYD9izU21KqYdAV/xdYB2xLqiftx5lUA9z4AMIMtAy8sataDPG8TuNo
8gSih3aKBQdX0L1JQjvixNTy8C4fntgqi2fSd4HD4EeBfyZwyUybGni2S+rj
9QEJxqnam4mFZECZ9QMBwx/K1/RWPG/8loITExhxgRzhnKhCWxvsT6pGWFwJ
xH3BTQtWpiMf8iPEDuStwhsmys9hCE0quXuZTPrjpKW2e33O4PWglN4EoUNM
PK2aM48yL2vmrzy/fK9oklbIxVo3USWiyf+l+WTeX5FXth9S81tZEcC3feoo
P77q4yfbOo63/0txkKS0svnUtcZGrG6R5f6p7ef0Bhl86VdeEOQ/jQ8mkqU2
PAclWwznPOPKXHFG/141edWLeCOw23MrFDRb4vKdTFZtEl/aacYgPsuNkjWk
HG/5CSQyG/I836kYDP1kaoB9J5qWpwU7l65d8etGl3XGKa+rSNQ96rN61bZd
fovJACqFz7EEMH2AHIQlXZPwJNilUvugfThn1Wv6Qr0Qr2DGKlAru8r3C9Q4
XqrEIWMpRiwBGAC5yp3wTwo5UbxR6Ab/3mmhjdMNWr1WGGVtelBonNBYS+XX
buhWtfUnbIa11f9uVtawZLnCq1RZbxRepwMzYAwgMBzqCHmTedDR5mLX0c3q
wSkU2Klb7CpyPvfGduLxmadpKnmPf5m0MTgdyAcdwgjif04+7EflZX5kwD1B
WiUrSZlO9w2BbMSt2g5oTutVmlnSV9cOKaSRo8PP9fZseS+7eK4v1vrvP+M8
8QA1BrYzISAjv3xp0ofE8MZjWHLeT5kjM4vhfxe0BOn6jbVkOr2+qKlx2Drz
K01A2o+eN+HtHxOEAHUB6p2Ffug6VJzhFqRJHBGefSRHyYFXFn5GR8K0aWcZ
ORsOjGfsupb+/GHUZT/bOLfX8GyJRy06jjp6Ed5hxENoEh6VV/sguz6TDdBb
F+QWKLAL4AjbY6AKV8DDlHnNQQnjo70S1khsDG2EuBsx26Xto4tyATCx8ZKk
/WzzvYZ+4XbQs7sP5R4IoQoOh+gkI7gMOe0MUKygp0wjhDiIUk8OrYeGR0cU
y6seWj2+o98mPesxmqoNsxu/3CXx4Q182fYImPlYyGnfvWEd8Rh+l7N1VAXl
yTmzvX3bRbRzRfLNncu2YqB1YCcPJUfpGQQ7WP1HPfAXfnj1GUlugiWD0W0r
Ocnb43iANh+3hdZ8+LczciO/u+rQu/gjtzkKzyBDCCLAvuubdkQFAmGlIvoS
n6gM1lBSY5JR7LC1sPUd9nVFzNZQzKN+3CiDapZHJbsG79MxW+WDB+z2H1z0
3vhh10gOtlgAfFmxwZTzPSVZqBSSQNBo/Fmt6SH9C+PsJy4wRITVcFX91rah
9BAsO8vZh+70G8If5Pehc+zRCN5O3Qq068yQEM9P0dGyvdxhI5RAnPYspx6n
WhCh9SrF5SQcWlF6XJHGJP3w4w4YUG0JLyBcBxb4MkOrCYGbqL+rhOCCrtGE
AixsmtELf16ehfixxJASALpTM2ily9VAQv+n7DU1bHFFB62f8tAGayox4OFd
Uxj2mRjZ5nlWiqeAnDWtXy4GXgFbrEyw3Il0fkWHGS5x8eBnJ8VBa1Jcdjcm
PL6JCvJuAAbe33764J8i5VnWAoH5krcEJ8zR3xG6IsTGVkGefF/gkTa6OZLf
IuHOiSTsIZX4XLdztQV6OqP/gyCTY33XkbhTp+Fx2MaYhMloz8IW4UUHh7u4
KW83t2jkF0aZJUDp5ZiLKGkTHKcLJS/4e5XUZqSjq5t2H4EZ3frBO6+iZmgk
yz2wIVpuZnJ/kRtKqubrdKS+eQKXOXhhHyG5HyP+RuCuLJbv8f6OlPrmB9aL
+3Ly0wZx4BJaDyhv10j9jHrZvPkemflouHnESYjUAVLpJIlnujADyVLrc0Wc
3laT89kQ/GLvdzM/IwoH3FnivvIUdh5zTG0P436588L/5SmAZVGR3+QDfMAB
V++Y/vzbR5d175eGJxivzLLBoW6PpAAafspsHnh8Xv2ht3IXVbK0TyyUlTeJ
PM8x3FC54+TVFN4quG5EBuQRNa2iR5YEbzij/ZtFdH2HmRMAcc02WxrOIRhE
H92bNDDKiURrrCw9a9WYzNfHXEv6Y/r0opPFXkWGasDmgJIYEwxS5VEDu5V9
sMuGmNjY+GWZZPNkZgUEwEfxFec8GTBNBSQ8WZmIDDtHnJDrPm/RtZ2oUjmc
MUelWCwLw36I5TCbvGqg818Tz1pmdlSCSiHLD19rpvwu5SpmElN6AvcbR0fq
vbSGuIE3U9U8si6bGANtULjQ89jqZi+4L4M5cx/6V1tkthS+WxJug5/lPkJ/
SJtJ4rXqK0S3GbtsBti+Ozopv0gstTaratyT8BV2DzwFeNX2y2w21g+fI83S
x4bG74sk1rnQTcb7XkkdtN9d9s5jhdQ5TAMwuWBciNBcAya7pcjm4SiD3Ng1
LDEupYwFIXdv8xyf/8z7qNCgBC8QQCkC2ukgDjZX15DAUKCzarD3SlwmhKxp
F9Fg6TnDR9lYd7STqbZAr+sucnXtSlfwqQ0I6JWH0cJlkFl9j6HNeLnnWKyg
kcnJMGHt6ZKQ3fZxqfA87HFWWnNG6DC4j10ayud0qJY0y4MabnX3MIKJDNeJ
lnxLIjxon9u6PODK+7eZiHHth+laDOvVOc1AzulWyOXtv2EVmC9GxWUfwkGm
/BVzpPypC5iogUGeHCdLaMFhCnYwUGshP70Xd3HcmCVyy4464soL9tznTAar
J6hjiFfiTxJAUkDEo7kKpY0B5y3+gG57iRlDWEVArYBcJArz+Ymw+QcK+mUk
NPYsnIhT/NJMUlVQp0a6XLvKJRLX/d6eLgkbSnILpABojATKjrGsAQWZB4sV
Q9VbbecYoyvHARAFK1at7l01R6S0lEnqaBujI3H7F9OHholdQsxAaeP80axD
93VlnRcEZWJaHnHwg3rX2Ir5pe/Np3T/XGmhCoeXvxMxdVSqZ547AMDY3Waa
3+qrLtwXRpjpKJ46SNmhOE8x61EWiPEKOYlvqgLYDrZmDT2sS2G32h2FFTq5
QURyFmXwljJLlu84iFnB77Z0rYZ7kUfzC1afuj5K3BWoLl0yG8ejirbmVeSB
4lNGG72prxdBx1YjIiIbhCTeqKUkbC2HzkO1PyZqT4hYV5CYF8gC4hHPOwA/
Y8mr+eX/WzU8Spl4xL2Z4MLSCAcBBW+o8wLccitXPV1VwtuSS8d5nwq9juAB
j5m2I5r00LKvpcPm7TkuSEQK7EC58GmBkKXG+78YcRz5Bf/6uT/g/BLti8r1
EEGfWTyr1sTTd439DwO+n/KndpzpGtwVwaUdI2Ao7eHxiUaMXQFdtGZy2k7L
SHePkULsHKsIH1AyW/gdlNqhIxkltjtmWBynJRzZ4xBJ4ndDV55pi8Sl61p0
Of2rhkD/z2yIQpd7VODiErABSIIOjX2F4cIThplw/oSGfjyqvWXZ3hS9MpRQ
KpPr5aycVa3brSrorV2nAtnpXQSLyBIn2O/q/gKx9/wIesdkYkfj4AQMM67g
cREbMBxjjOAWmvg8d2fKEEEhlCjCG/NroNwzPKD0ATuIFT+w6+DF04Y++cYX
S4vlGs2zOCYGqw/j1AYvkQytwypVXOrQ+NcnXD3ksD1FgEjJdnaqICUb4YnJ
RH5A1TFk9pGcHTvfMpghhImzx2XahNNB+1Z7ahevvlta4KatFy+F6yNTazLo
rHVJSy0C2SdZ64vjCy7k1AIupUDDZGxWdxD3RJ/Ez/H6EwMs0FeHPck4dsYR
alprvOCn0Xd1WiXjYTOIOSRc8fiC9FHXxezBEizxSjzE596sJtq3cpOueAfB
mzDtj1xRQo79E2sRhxZYCRpG3Y8oVTYzZo/C+1mFs5jlTTfdiGMXoyIpCcxb
xuNMZCpobIjGJldnFPV4kq5wyxL5Ajh6l1leDsndTOiNSvDdA8YSC8dtQRuV
jwFWo5Jqt1TFv/LeoxWu6+CdkqadA8mXybMuo5nvwCIB+A79vNNP1m7183oX
pRj9flAQe+S2EcaT8cSCL9BQkQMJNbNL4FaSDicT0DGh8h+j14/jvIPbVOM8
M2qHo/FXKXgS/TVMn5Vtm+RBJxuwR4MiYlpnTCve9dSXanPYLER8Mhx69pfc
K1huB3/IWUhQ69SxPSC6EQFwsiQfgFzUQq22I6iQTVMJecDe8KvbX0P1NPMK
7Nl8Qrtur738a3SCE3lalHXFj6ThGbB1/aSNYnP01nXflPlrujW1dpBEWug+
EDnOES/sszKoLjU8PE01/1GJa1Ou8wb5QS4HHdwEem5G0hVFRYhin7JSbCHT
0fYGySwthDsL8x35atrAvKNQ4djMKU2v+lAY1RVmGiEZj+ssizvivi/dpelx
ktMQ907zEINDu9iAgnz+B3ExcUL8PmUjnv0hUwQNwahZpVUk14H0MeKFnqw1
Oz7JzVChlRogBWN/yDl6qZSeSY1qdNZ0DLphur1+yGpluqSNMhLkHNAVYPrs
foYjfQM8qUPG8dH16ewreiOJFmo17nBvWQCMrImB99c0sb55R/WK3FOFVsVl
wQ20ZV14jOzTlBiM75g/C/Q3qrslrRrRC0ReoiwT64bZt5EZr78lzGoWQIGH
6XrPPYs0b5H7+lRrVdzKWL72FigT2T4Wb13lDduECvTId/bDqMbUFdgq0Aw3
Xo/TiOowrP5eWKD2rI4mVp1hoilhQ0R+VhWBu6tBJXIFpywsxetVVR5yMmFP
MtWHZbgl4/DEnqPd9WPuvW+tzV6G69Jf4L4rLNSAd9jYC/59rH8c0wrU8+T9
9vNwnmYCeXMqu4t3bk4YzhrTzAScxUmzoPOo1kWOFi7jPVUP4/fzqaZlFDGB
K9Zc4fS4iayOp+viD15wzgF2PUDo+5XBrfrZvCJZgHS1BADFCadmY3Fw/Byc
wBBX8Gj/e6AvdPKLiAM38SfwApkeXKgF/tY2dt+mNnVTJOGe0pMaiRlqKbTx
wRHOfiBIyb+WxZZrSoi8E/L7vea7hoPulx5pHPhNWgB3NhQP8OSvm5A/Xkym
Pz/sMfjZ219xM8HdIQiMaMHayXVptZD4AEmHk4kTCXFOQMBrR2ur3+bvz/PT
qKmcTfVvpX9tqTCJ/u0P/758Gc/k15g/WBP4G3FBzqgTHNC1bBXQk+G7hEay
cnSOXFyLgtqor36vU8+RYpA3XEQGV3O/2zSu4PrinII/OGIJiV3Hk/6SdTKe
OQ5ZZGHYS8QN0PI2CrDLQAbAC6396t50c8eJvXQhaqpzjMwPltVidRB4C/F5
6YW6FABPRdxlAFdLTe8S9hQW1RHNrZILKW9hPGFm1uhP5UuFypxQMJmTqGft
IVN4ocdp8MLfXejumrBvxEeqzp9appcCb7ezKNP4qZAHcKTJSrvL4ZyRmD96
Mc3KgeuNP1ErQga30Ok6juFtbGvCh4NlYb4wtktPGeAbaP/hq8Yb0vjTJ/HI
5pR04gR1oIum0h8JzF42kTZqNWYkJXfrdSvN5qW+LXgZs4GlKs9QtAHgJucE
aJHa6vLJdcwkq3/Gcnki4dJbOkc8kwFLH9foXF6kyasDohwdCBzdVRraZ/zX
i3Qd4Yu0auDck6kMQFXcDGd1/QASaArHZvfewvc/MBK1As2cNB9Firha/Mbk
DYm2Ushupn4j7sabb5sfOooRK63AJXtDMQUcZbvgwpUxOx5wGWy8nq6cLbjZ
U93OvsFRHn7ipUSnBqJrSzliXY0fFThB35d3RxnxwQspVTZRj4ZbJ4nyXeFX
UzoTWKugQd+jwmT15ZAVOnV9utrptBSmD+oArpPXYgjG38AAifsJs9FPXr+J
OuYFXTyQZA/d/9VvC/uW9LkDiT/PQVQZ8jnJ1sJeqAvGoD0bzgg4ovaJ+Wsj
/4F1X/n0PHv5luHkj5HgRpLvziLqDB6CvLBX+lKEI+lKhync31vPw2j6su0f
EQm/a/D58JrS1/2SDwO1NBswggJWxj4dxuw+u0uI57zjV6ncC1Up8E0BqrYQ
x8lnwzAk7ryn+GZjXAhpaBrO4IHujsSGPmYilT2ZI7/M8sLdvTKIT6BRNsTM
Cu/HHeBeEqO44Hvo5M2he7PP33kvnhmYV2oev6NKanP7TcnvycjbNMVEZOEJ
e4erKqSiuRUg3wV0nub2DIErD38y7oh87Tb+pZyh1pjn4eAvFQG9QACKEyRK
+g+bHJtE5kUQrIsfJQS0UY+Ok++kHHkg/3c/rN8SpYofnexA5b714IT0iKgt
M46cm1db5umvktUkqvIivyUFsR8hFZPJLzJflmjqGk2N7XJ3sklilrZPDzZ8
0puUOYQwtJULVYEEAY3QalYR3wwgJFNBxTfMYEsOFYJbMPtFI1FVTIwSEopu
CD2bHjxqc1csahQPcXTuj2TJpdFPh95X1PYh3tJieNPJ3R+hjg7kHbxm6G9Z
HiK3PKn7xxKITmXzaY1lLS7H6LWx0gons6oNIphi0fuWWlyVIfM5B/gn6Rhj
iszCAUnUEiR60vlrbGYTaFpo/macMSwMohLe8Kl6btC9ZiIX/OgJAzPxsPuQ
bbxcFpsOBpJHZjcWe/PzjHz7ZDQLhBw/aCJBcP+HqDAJ4yRMmFyyPO60XrMA
ecODd9wOZoL//BYHgYg0a5UE/tdGmEFsdjaeZFbNjb7WowEv6VBjKVntnncn
wRn9eAu1Ag3NZ6C7fyKANkYSE6FDVvFckRsgrrpxcXC34y5+9q5679mHNgEN
6gXPTwvz6IZugGTo5jj2Y61rnn+uMDUhkpzqsC2tlxwUhprxsJ7XjCmoC+P8
rc5FXhGmbUylQYMZfTxygWpnm4XZ3lD2eGWLqAjSTi6EgciD8HGLMkNuXfoG
H+zCDwo4quDiL/WnpV5j46QMy8wXMzGvDUALXHgNm6MdYAd6Cw2j6a2YMcQy
86+5A67lf+aS7AiKflZm62HB1ALy4DWho/cPwf//KCKoUkQf1f8/pDVjgp+b
knW60szF/e8KVGBQJnA0lglKSPaPE2FFYMyKfBVYguQixAWQXN6GpdrP87Rp
JMaY2Dwlcuq11MpTuRD7Xgr8B4+yTlYxI0zYeD3l0ibqql9VgkZ2k8ubpFdJ
DGqUcFezEQdSE6NcgprBH6CEkvNg2/ta3hJr+JCSV5X6NNiA/VgRiroxGDtd
7Wx3Hmu5sCZut2ky26HAevpp6c+v9Hj0xQ9GxvgMfmk8AR21WdJYC/r5J7PR
FPgoZIG0M1mptZHtrcFmSUjx+9Zf86MSFXUQIvEppJZ6LzDlsjB9jmg41QMP
OlpnkHK1oVqqKBRfh+L7ZHTzYqO3ActjU5X6ATIXc1cKOfM8JScuzxyYJzgC
VSlrZNovrbq3ivXmswTvzpNEj4/6IDADGA5N/qcKHAXFF6UqTkGtHg5aPHXX
p3cxs113W7XKNE5h0io80TS319/+2GX6cs4iR5CcTCsEcp7jrwAP/m6PRWeJ
QpsVgD7KBjSchZXI4wwe6Gf3NEj58HneiTLut2k4mEQJcu8p+oNClT2VjPLU
3XM5cOpf9jLRQPnggLnN1UnnRRzubGSwlxwk7uo4AtAhLaMwjgr7r/b+ec5a
Qejs29hgeY3/xV6UcO/MC4T06YkxzeJM9wC5mwLv6N7mcOnEtaVh0xrBi6b4
s1oBMNdPtU3fsG0uFpt9g19Dcp7Cm9aFxTYoBvz+YWs3ERdT/r/Q7mxWrIic
/G11PZ8JwLAPYH3WDGQdMUob9X8lHqNGPFGxIH5Wc4ZXim4094/7ptGkNTzk
yv8jSn3llVOgLdyPb67P95Us/uHawCZP3ATMAk0RFBdGC35i51ZxXLhgNXiY
C0aFPQz/SmIxAbjg0I8D9iwsHc695vIOzXs2NK077OJCclX/xbPe+Z3hZeEx
3C4SR9Jg9tglUE5kTS54KSl7YqU3btx0fyMbOehZv2VIeo4MVlu/sJxM+4VF
w0VaGA8hio9KmoUr36G4MZj0b2eYnBmkmLCejdZDQFNDCCShaaLTHv51DBbZ
zRJ8V7MLu8Ut2Q43fT8b/kHH8aMM8gNXE2QzjmWx73ErP4rzS5dE1zMahZCv
wl8MlBJUw/fI5OxVLQTjEs8vgOdeB8lN2rU1F1dDN6rHRymJd4NXa48G4kFp
0/QvF7PsLeP4nCEe3mSPaYpCDiOIAfwEE1Mwog03lmy7F9Ugd3FLesLfymJD
O4chcJOHDYqzmuSGqw8mrQ+S7OfbZolingajdEqVwxiTEyhBRF2wwxDFana+
rvMM5mP47YADaUARXokRtefR9HMYxQ5R//fJZgoDg/pAQLjMRxhDyRgWQCKR
9PKjIBH+28p7UyDr+qwz0mOsHpvmev+ffOl5HfFLDsswpdH3wvrSi0TLn2DU
C6B49JZ1Yx5n6v7O/Eg5axTLQOofik8tiEOIxszvPC/GCEFEs/ydS/Rnmn4S
XTLljcZaAB1BMj6K3Shq7Uv36p1/zUS9BhwgXCJv8fG6j+3AkuoSB42SW7Kq
lQW9ZrYbICAFkbs2sBBz5+XRXPw3OMyk/cnk4/DEmfIYckAvikr3eyIxpycl
sHIWQcW+en1G0ap01UqR/2SboYDY/Xn+p+4vmpJdm0XO1ymr9A1lyw2foo5c
pIAbk0kY3QhuF1XqY80yEo93uQ6Np+ELCCQFaXoens6ix0ZpT2Nl+tjSij6o
Qi3a8EBzKrRFgU0uVGj/I5NJTeS9zRthQLRHdPlo2aRd1igOvAmZ/Jou0EVA
mAbSqvZNCShdCcl+LXuZqfoCJxjxvUDbzAcC2fdycLSFXzyBS1paS0JrhZ15
CB2h7VbFSj3jOyNdfkxNrUZMWfJNeXu7n8gIMp0WJwLbAQeKEcnBz9uCsNRY
iDd2532WyOJ4zncXrFgfeL7okdUfMjKAQsr5wq/Pl5SfPOFlKRITqPqiZe0I
NEoG7Mf2CbtWq1DJceIjwOfIq62j/BAybjK8sARvI5x1VmobpQ2kmylqd43x
VxALrwLkSF7wHeU3s1e1w/caQ6JO6q5DsJ3Z682NF1PIPE7eMTFukCc7Wku8
ROpTDrFRJjSz+E+SEeOyd8LmWQ5gb3Cc9sa0NYiMyOalNYra36T68XfICkSS
VayARmuoDRpgRIxxJqw1Xl/6JZYIlP5PPFZ5sKHgkZxDbM6UxlEx5QGkAhLG
Ief3jD/MwxmOKZ1xW6p+g7aA5TXgnyfDeqX3xdR8hoteteMh1BDRSDs7bu0X
hERcAovePHPGCN/6w7UlHyKof0mpg8H5cl7JPw0s7ONmO9AzxduJKJdvy6J9
Y2v4wfZKNI0M/Lbuqivjg+5ZTqBj4rz7rfFqUXQOekL/sLa84NHmHrV92E6x
hHrzW1nbbALG6t1gNelSM8AxZk3nkBJ0dHb1NzDudW2WFLU7Rufys8pD4YxZ
nLXc1AKiU63AKpOvXoUTvYtLvjU+7qjOB1ZUxtrNU+qVVIY5tOFCzcC9YBGB
GGjvZfy45YjdMBg1le0NKryl8KVC5dsq97zoLT/CbXpa1mugXPW8wrPMuIR5
o5RUyMMC4ZasTLAHE48LZJ6gSy495Ak9kGZhUfhcw5rhJ5UY3nJbnWYQnqS5
cONE3/QTE4g82hVVQmbxvISLtbUA+8K93kXVibVUtbwEC6g8ExdabE3x8QEQ
omX/6+yaZpB1+D17OT4qJt1/ga/vuloU0YVhKjYcXtbvxbCICoYYki+yydEM
IN5c32ojk9PqJYtTOlsPabu0/gYQ6Jh4J7skODSMKdU0+DDnlBnsfTKaEb4V
jn5tdcyvAEfuasR3UgMDMziDHYkSg6f450TBLYQppKEeky3I1Nmz7mqDdH8a
+UlhPeVs3YD1jhqWJcOl2I+x+b1x3Wc3/2cMDxmE4kupRYHOo0ffF30XXyTq
zG3rQWz51HEAehhVTvUyJAwcFIoEctkaKoVWKxpUYVXpKLikBbI6t0gpjxPV
Hfcr/tBNyC8hugTkUev8RwrPT55C5cmXzxkBix8iF4TPyGtqQMYvSsbP3Eno
SoJWEQAS395OU6zGOhrw5rBQ90w8umTovmkjNaW6GRgLx/WFwTwUF+An3OGG
gfbxhcWvfHKeuiNfbezhgsyCx5UM90/KUNKtzWohffTWYaRPzockJaOV60ft
/gVjgUNywmDkp3wVK1rjVtPxKceOmQc/D6dRikpEv9Fy3PvdbjiTwzlEu2wI
eBt+FFYUe9OTipCrBLYh8nZE+I4G29P3mTbxN3ORW0i+9YUXQ/7u5gF6rCUo
hB/QAidLE1ISGFmD3WdiYj1Sua5meRH94q3JRCTlkaJYL+RB5tLr6MTGPw+R
BtOUujJLFlUI52vpn9V376viQoIDbcEy9st6K6m4u4nrrTt1DNFJGdeb5ATU
XCia13gWwrkLTcEq7xP5ihpQg3Y8XGQduyz4opSphS4/oNFU6Ts52nUNmcXI
Q9jHRMVZj/TEUSTKaWaDe/dJvlco/rZ6UrjGc7lEyt46WSNdhO/OLQqHgIiJ
Mx9p7kZN2nkZwaKbmlsmUH12wne2GMs2HJNJA8vZwnVQC3pBd6GRNVKeaC7Y
XU8Y0f7ge30gOLjnJw4qvsWYHFTJBEF0L2D0AppN1gOyMqchBs7E2B22fH81
VLpndw8KR4LyQ3qDS4+QhBaMcTujlv8i1P/dFK4+3eLkpmpGKfImRJcXlPEL
emJb1FXmW24DwonnbQ41jXQw/FVW2KmTYHPzrnfbzEserkwkkqzmFZjmz+XX
Fl4afVD346SfIPIBkaoYz/QcAIGMf6Te+l+Sts+w1DhJRrAdVJWo29EbwKxc
siVJ1D+sCo0AyPc69IklLkfTGezPPpmbTZ7sK9KDhdZQeDmkPwrWdDG5SlRn
QGjSBzv0d2TLcWgxG5fFBAcJCN4WgHwC+rVOGZFJXDrNvrlaPzifDCXBP8x1
6C2f4eFjQj5FANq7Z5zCtkBHP3Pt0BvpIscDMyzfZbPYf+5NfxYxhVt6VCV+
fEyqxFrFe/FK1NUz++jBgAkwkL9nx06cN1+qhq5ld6McXyLIRPaNZBMYOsiW
GZH6FixsTh9AA666BGfM1tGdoxI/xlXVzHbweUe47X0FF24H4Id40T71KOEE
TTXEtMgQFUu/pJ5I6Q/A2AisE7JN8YBSnHjonwKBZTgb6ZsZ0kKTuWbFNWqw
LMFJ3aKEQXUSXx9069DAKOG0yGo2SzguR9hMlM7cVm1IYvqWwzH/M8V+rWqZ
1BwyaEnrQyuPKGmrWIZoNYmhXeiCDpYyFka6bLk9M9JWro0MKNTpfU0yl2lh
P8Hqucf/EUrsuquFj666qrcOmQYASY5HTZBqxzW0KJbYqpNyke9aEDCE8OaR
9Wx4DY3EWM8gH4h4HX1nlG/Rq2mUN9RqvsFWecRlSTaab3T26hLLxt5mUEjw
kwPu8isWJDURiWO2zqqwWRcd/+eSKIBeJ14pjYYUCiOncZUUOKoIXFKnWfI0
0rVJ9987AsN439S8OlBRxeXHC/YUwIZmN6bX51ct1xbgExKNzy1iBBW8ruYD
CE0OV17MYzgbfbQw0/CH3aGtvQgDMw6stXrZfmCdKg88GddpKr75VWqIBvjs
1XM5B05m2zcawluFcWpPhTftoI32NpPyAiD4V0YM710z3PA/a8zxUxe8j0Z1
P5CSzNTbgDC5LlgDxa59STKoRd4R7Czz4JMjZGrHEFHx9QcL7/zESG4zz907
qjevTzCJg7aRiJI47HUrF6t1z94INpNFjMtqvUFgm0Di8uFu4+LvkH9CmTn2
M4h5fHUobjvO/w/czyyMHpqF29UFzm4He61apmY7lUqajd6mI7jM5tfQJWjG
gTcX7yrk7acnr1FfbgXWJloIzNZGYZZjQ+KR+fxhkYm7aN/RQaKI93TcO0N7
VLXozDZR1UN8wDQwHjuod0FEI1Xi82wrxpxr+GelsCaDc35QMMHEqVUM3fGn
h4dc2MPxfDLBBNr64TQNTUxLZcct8glwoNmsl8v7A0ZKHtKN8ZMg19NJty7B
rJ/WaUEMiKlZbF+yP5Wc2kfVV835EuKXAOXEUmstMBSF3BIrbed00DhABZ+T
DrxLD/tsaKaZIZ9t2GdBfIEFFl1REjDkQBhEaJHJqlu6eK2mdvrFCSELBLkt
ODLMRk7w7z8wYtkMy91BnX+kDBDoBNnW3OYq5mWnn6q1DNXYGhLBH5heyM44
Iq3z1iix6ie00O+bx7drMOebqlfzUrnbYUYvG8AMvJWiPCiuT+tcXl+VNlZQ
+e1CVHhyWtD0bJTxITD7LY9jz8XDq5JCShSvVj2OCWBp36g4NIkbsU78MQWC
fXPRR3n5bxb+q0mj+IGgHlMzjonxh62mXaIgU05gu36PoNPtRkTvLibtSrqJ
OsfMhp3sBy7gZyAsTOKeBVHZjYnK/9oQ1Kz31qbbyDmdvSInzp7D1YYmulm9
Uy0rrEAXbBvyKQF3WjU8U78XYeexOGt9jAMc0B/qv6/I4v4wmUgTWe22hzRh
cdvG1dsi/dPMJANOSO7617IqqrL2JFyY3tLx7kLMUbU9kQcnDauuGdji2OAd
MSczB+UQ+P6eSb7zAiGzJRCXh68PHaHlvEIYHT6r+ffHhZ08orCItvqiPp/R
I/TzYmUNosO2h1DBHrBDhO27E+vB+xQZZZRAnZavwaruAaKG2Q/fI1eKvSgL
dR4+jKmOBNuWE6Y+gZuCCeWlWHsX0dhbcn8mptCtCvvnSZbRMysz/ct2PF2E
x1psREsbJPC2TgSuitow8UvucEjagDm/WVX9xBtmZAM+dcwwqeMOt9lb6wd9
RTF3Xh2rtRi58d0kQsSWsxxwdhUt0gt8xnX66Jx0H3KiXwzudR1q0WSRetgs
q+jopjSZmLifRFjwLrtPIL1Mu6toD5VD44wXMv9VuvTZdaJRHQTzHfA/qyzM
8VmmKtRmR8rlidR2PtC7IvQrY4wCaW+JTaYYl0Fy7KQzFJy6eieWFLP6sdwu
rLjhQ6SG4ZKMqlKwchDT62EziBdOJDcBddairKsUFZyj+YOnKFCC874hoi2A
x53Ha0IMEAYJIlWaSe62volJ8otFBG5j29LJUBFiTw8Rsk7htQNN4asnTBLG
psL/FvdQxA5ZTpWVU3Tu1R+EFYn87oxtlLDbt+8Bq38+/Qj21JakW4N0esAq
czdq3OIyGfSfB2gJH4+CEswJXsao/4Vwiv8Xr4gSz3dqxAFNphev8jahLH37
B0zBrn+VTdeX+y0fRKH/Vmj9YRC95l2i3FuKMkZ3vK9AOKdG5ANPpjU6v80x
nkpfLePCmN/GBI6YppfcMKj4loQHs5qlo/M8tKV4sOwaNU3IMACqUzpBNAey
4qjZ4xuvEsUO3sx6hbrJIaPnON+bkKieU40MG4IYi1fn7c3fssmN/ZeJxJBs
h+roRHw39Xhr6m2iiuJygLEhLrm3naEbtKvM2Fd4z0IhM+RUrCdywUS6xuiC
7hzGpRUuq3/UAsMWpzZyaF/ICRhN0NNngmRHeuJlRik4P1in8qhZUqxbDxWT
FyJ3rgylULU5TT9qtEG72J0wUQ8lJklPT5JvwG1i/DwdZhbfJ/s7elbD2t9s
rZ9iI+Vwq2vdK5MjZ7ZVSjqRHQEahE9dNKLuPVLTcjG/Db7drQzvo9XuAk9x
ssxMhnJs3IX494SWYDXMdB3Inb6/cblW0nEmO3Ohveglfini7hsAcPgeKDgP
Uhg1P0cfgS5T9PbGeSGdsZVnMf3EEuqwgLjJl71+ICq9Tv0IdsH+kkfovwcd
hDxulDnwyYEBa2YiaHzhf+bMsRemJyRttlQMPTA6H10QDWsd3xR8fIv9RgZi
yJIQ/Huaj9TFoXMrnvAnxVru2+GYyclcvb4Khy0ThetEcDD/qbMqvM9YDK0Y
wyM25cgx8VrHOMG4UV+j4HGgyaRoMNCTxh8OD5gCF/GRMe8Da+vIRXOL3DUL
WZ7ctGrHccgvga0P6n30sTwvwxLpNhnEiPdmefHGtJiRf0SIpgx3l+Krt+Fd
xBn8hiRIfzSWdWc9aqFNif0tIgvknQ8Ikv9LKlVt+kYA15TSleoY0dtVgCyX
4S2JvV3YvlQcvokFf7+jhE1e9aVGtTdKGOVQ/prbU7spNEde3ApZEtgY9xUn
dAuBFETeNgr+N+J2DeLhlnWJFANxTiW85Nuyr/5pRfK20TZYGg7+8rXfm4u/
lL0JrHWch3z1WF8AR6KC+UZQp8gH0CLXhRn/EYHE8RMeFUYJDCPzQqoESmzm
89JXPvD5Pnb2YexOhTv2sTz3+LVb431UxiXCNPLzSCwGKuWh6waiS0szuLWt
tr0d5+REQ4WtlY0DJHlPL3TGLQk/aTnTtQjObY2Egv21I6SDYmSSYYwMHFnP
1TlI1XRXxnCiZE2pSBbAOuF2HtfS72sLOw20ERaPrn0VOIg1cYcYiNVchCPS
vQUZ2StooRnSej3Nsx75NEDW9GSBMcFISmy39z/xTotnJpPlDzds2lIyfqas
Uk7YTI1qObNN/UgUSSqQjP08MPzJYL3pRpSStR6nGCy0W3cPC/OLHKd70Uwv
7e3K4IibJEwanoJ74XgPgLHshKCF3egIYSNgBqN3MKpFhU5Y4xTL1HW8kPKE
nf8malxOAL7kOGfwrx80VpcdBRxYwa3FGGeEi/dpW7F4haJLUipZEEEkwp3h
JKw+pe5snWn3EOU0c9KMSjYe7Y6Y0KyRml3yHELJDtRWCTZP6ehkhJ1SWQJ9
3yItn9pnYyNCGzMgQwb8MPcEBfwayFzFgEhEDevQxb9Mnp4wCWy1zyrswxOo
YHlonOBVACqU5r9DZm/djRbvrMTt/iYbjxRmm7u4yf7ls0xy6mbWN73rY6Ab
gTvbxUwRc8Rv8JsF3DMkGC0/G9DK5hL1r5STOka9rfBZmJ4D2v+Z6WLljN6b
hhv3pmPwzSdl6j236kbzuSNNdVcmWUUurI4HFAd4IRyDW8pGOLruZGCOO939
x+5qEAIIRUXLuarXeDTh254cd2FFH+VETWwJ5wd53Zgex2QzcnT9ddGdQfsC
ARAUU0V+FZ0/QAWJm9CWgP5dWYrkPxCZP6a3Z58YnWMvDNbXmEA9INj5Wk+q
2m9fDu5x2zWXbXneBLhQRLN3sXe5jdCVKhPWe8684BhcF2arNtsdeuDdFxbJ
Pkqi6ONGBcu0vcgxYGVNEsku4N/PeMjufNQYUyZX1xoBNW/fUKvgtrFdo2Ei
dqmdV3ey0YqbIcQYIAkIdfIDN84/gfEIIQwl8mkngPPyMdybYUk0TWalVpa/
GtYxPoj0q0pIcDtwm2WFtPvLpRsgXzqWpZ7uB00j5PS9gyRR8JpPwWeWn5me
+G9uHeoOhksbYR+I97r19tnIeU/pxzaY+quVuYBlX1kzVCjhFsbhXbnz78av
EIYf5uBvTh/olxQob/eaT8DY1VIOj/eJ3W4c21pLeRqPC6u/f9391K9INTaO
6pg31z3XELZWo2f3w6rB8ZMZwbaQJQsUwiLnmdpyhGBHDhDytpTLRONvBX1d
z0NNkYIkHw5p5c5xmK2z13PywEpVyY7n8FQ7baddp1IZMGhgtJA7GI/FMnb3
fGv2J7tvVMbcyshGOBCIB5DkGrmhcrZ5Jlbe+JPZjC3k4UNQAqzUhKu10tVf
UCRScyoLqvFCKAvgFYZQtaRFXHIWV2qwqTYdmmQgAXnUC6tc8vPE+D7f7oSk
8HniPhNU+G+VmUVfltswHWTGpBcRC0SYYobl8KkSbG9sJvu9xmZuAVzDL21u
AQyerXODtkFelC9BMiy5dGSkwMW+qxnINJpCjUnKdaL1TFEkL57ojpJR2s3G
eg0672InUeQMn+4uUQwYZawfgsg88PEbh4/zsseRCsWKWQ8tJpGOlNWo4tXb
wZwEwtcbqSwej4vZ/jH4KhiwGxILGbGzpwh525CPv9LiVIUvGIhw24EBpaUx
baKkZpVldH5KkqXjiohnnIWLYRdoxz1UmXghorAkZ3P+JebYqQW9j4MR+vGi
AKP6/0blfIfXMN3VyLMNLUdaCc2mJ2ZEYg/zHPGsR2PMXa5Stt5m9/QlFN/d
j59YkMFDElmoL2nPlNJtSALK9iUI/Q2y3S2KwJ80R5CnMCeF71WYcNcEEYZE
YchL+tGbT8uxGFQQbC2snnI1VgsbXEmBPGVoxGNok7Wm3YE+N5Amg22R+ECk
3ZVxB62nUo3SFYaetVhMnJvU3xuVjWKKqP8hexzA0M0kQVuXGyEFkrmlvM64
4Mh6Ib7GT5KdfFHXPdiDfaS8+BpWN9n6UtqhpQ5qgnqCTtZ27l5I8G+3S9X0
LOL11ipR+YD6ai4QQDmeXReDppHsukHcGG21OK9OK/ajesoWuxQM6QBa/3t6
Wp5vOKsn5ouBmlS2V6BE16Coz7dKTvRqk49Vug3W0J/9KV/FjmSU0KGZvn8N
lluhbgs96WLh1Cm+aAb4BfdIEHBQG4rHw0p3XGDzf7q4oa/cicUQoYqOhJ5l
/35K3215luJYvpDSPD8XML6qStwBeQAIAyvbjh3f/LxnxoU8UVBSj+UV9lsG
MxRyuFIuZs1dkgT8cXiufABMo96zD0PZ4bPgRw+xQ0lDXkqI6k8ZYQ9FztZn
1RnRTp7r3W0NbBuCciw567QsTDjY0+nDIlPvolNQ3Go8tayf7pxV0bn2Xg2U
8nMbyCfLjOc3hCpIEKm/0ufh+YlUzDQbSjaL/EV+Gz6ry0Zl9MXqglRB5Be9
gdZgkDSIXb4I4+T9z0ngJr4qqNzoH98CJfFrpnU4HBirUYVAlMft7zjZwG8I
X5YLieo4OJn2J3i5f+NSdGH5x67uUcQKrhtsfIhKgbZ5QTXPLrwWc1FHdAWf
vG/9gAnsp1fXV0FObAD2mPcPuE1iw5jnldwXFmssRExa7hAeQadunKsUBnx+
JJqA5/cUcC4Qi9DTlNsByoJBAfh6pwKhKSqApGYXwwaQv0B7TJ/o+bIZP0Xp
MbSYzPOLRtuJ45SqQ+ZLrROs9p1gxwTXt0sdf34f1eyHp703qODgtdc04nb1
5BFu9mqR0ZC+/RLFS1CQW9aPmdku+rxsYXmJFKHNsrpVXYoatg0L2AGJk3uK
Ht3rVOk2rLxBwMCAj9jwZPm7/rJvpOmzBZRn0LJCK1noeRLtlUFhQp8cWvWL
Uz3Eio6q4pRqxr6EAtnlYEzAGtSijnmmSSx254LQjMXkkPGv3VXfQ0u/11b3
5ZuUr/KAc9eQ8YRspeD/PEfGNIRVgdFaKueXebgBmJ7aJnKEzOG156Qdty/n
fyGKmUPzqAz/bN63eJ+IruIoqYIPAVGBANsAR4zZw9Ftr+j1D93K0kzTAQ7m
oCk4jQp/qUJkCMgz8Pui6K71HTO9qBJ6e09aY+o5LASwqGxTZkHxJKMlL9Mw
5hLUPauhQ/UV9sPC+XAdQcaB3OSKLKYrs74+3vAG+Vq9eDWL3ZJB5XuQJQiM
QVkdDT6tSG7pxPWLZgU2JSA2aejL9TXGN2x/tXmV51jJogprWRnjvAh3pzmm
rn5brj0SdVVr9MjWfR1z3/5mvDTOfvNaFJZSRmsg8LMLyO6o1QvxX1p8oRpf
YLDhYfVa89ZVUOwpuA5eaL1qfIuX0BfONSqoWLbm0XyPyzoEFztkJlbiJJVE
rpd7t0r8ja+Az/5YZr7kfRqSt5mdt0O4lvcEcmaBmbCZpx9/Nvgcmz7CNDvJ
9GaVOS8JkVZzAylQmHSDha00bjmn2tClxfaV/dUOiUrwUmOpnHjeocUcDLxI
WbW7W7ZvTpC1AiUsJ2xdU+M76LahxOlVUM8JluhTQcapYfUzjrO+Muj0RA14
N8cfAmyr/+hfIb7dgZZQhShQv/XYwgn4FwlyG1ioWnpp2CTjDTrXxTFL7hRk
OpCvzkCz3AWSmWmbET/u4kFtDDOOqTVFJLY/W2p2GjsZEkf9usJTPmYV7w4m
QuFQwr/FSV5cWRC2RHR9fXUknTeiMgK2MJTWP2D/7ewYX3EBRtxWKNT6VLbl
GMUdKCuieCl/gFinsrhsRhDuDxb8IzI5nfA4V74DgI8ic+ckGrnp7ITh6YKf
/iA/8q04JtSfFvherb91W5HlH9OPSTf7KelIhlh5nTXFiMyP/MQyKp1tlnW3
aR3JO51IOUPyh1nNBrzFmBu40ReGwtMW1CgGElgMyGcO37w36+FU6lcuibVx
VWJJosc3c4RngzXJZETi0ei7TUeYsi+GiTJZ5Wk1U3hU2n+0u2wC503H6Dr8
7SAkl8aDiYtPTU3CiI+qUQor12rxX+Ui3MizhhWHfvT4aSCIy5Jz1Gpq1/rk
BfE+XTjiZ4rC+doukxrRRHlkfBbP6DuQl5ktLxpWPcIbH+zxUQRk+KNwgbS/
hjRYD0Ww7TPJgIFis0TdBI52/k/OieJednJtQR6TtSBA6tg/BltUI0V6nEDn
IjUCLyRCNyOp8wZPxD2Am2fInrmcr0sdOShUD8/Bhu/kADpJHARqKeG4lE+H
ypA9umZ8YLJCVltM+MEALyXp4ODmbbsa02CTDRiSa5dYlReJQIEvuor1KxDj
MZOv2wJQfCm4tI/CVH0ZxFggeYjZCzLaMKe+HDgwt3NfcM2ToS5rIXwopUB5
EwAwGaJkfTSO4guwSd6YihTu+xHZfU3qx9QKHkUQsLcOe7uAjXys+BrSwOyq
ydMsCwrgRTeP8BuZzNp/3pGVrEBFG9hjkT4qxCjAjR862ebtK8F7p2mjrkJ8
BDYTF8ypc0lE9uwgVF1mY0uwgpWhg32k44ew61cqAlgjKH0V3JsMf0y3P8qy
BjcKuYDrrqZK0M0+KcS9/pblA4qPfCL/qnXom6pbVGf2D+4AU5wuOsEZsNJb
3DfLgUdpUVImaY7UXwY92CaJ/nLWg0DiQYcx+DFE9aeteoTp6gBIrdGJP1hC
cdNFBrCEkYVx9Wz0obTMDtdNnmRhbvfyi/yP2dIGBQuihN3a5+Q4jOQgmnwA
ErKB9ZK419fXNIOWW9NNJbsuTTQjJB3w2dPkDuJ9bRqnnzvTd854PvSikpgN
Xy+ywGqJyXzWtifIAIUOt8lWcj6eGFvrHf9JANP7yAzQIFiY2VQr1ZhCgmMx
x/aZFuyVlQ3mqkV2waO1BFpmr5BAoZDkg5Fg5Lq5raF6vQgB32ITXhg+T+O6
SEepCbCB5+VN+6lr5TSYoSsqlXP6+QgP9EpXPtsio45Ek/mkylOePDx879GA
3XfZ8zFzyyzINoAYjFxWKoXxbvWTFmg5rJ0gFojq8u/diVBsbE8j4q9G15hO
IE1WrbmwlcgUVBGbKtifTPB1jkaxaC0QxDtM+wHk0X2xyH29iUvKSO0IfZ8X
czvdB1kOBo19BLuGHHzeG+uOnN3Vax4kOfFsecE6hnaLH1gcnvswHCFBQIk4
slhZEqi7c72cahzdHCdEoM1rzVj84O9dRr7TXzXUatThfanm9KtLaVWWeSje
ZmtmEU1e5ms3TIvcSTGYqGuDXsladw8FmF9lV0iL2OXF3tgfGqDb2kLq/eI0
O7+j1UxuDtv/WpFUxsBKQYdkJ/wVwMSr7FDCsawtUZyOYsu0BjbTuGoDVKI2
HkE/4qappSHXrV2F+wds0XVf0r3vR1H+1pKQo4mD5JpVCxCBYDSv67bZ8+4I
y95PQv3TsYBK+IM2qtX8QKqT9ZhkxC3cV4Eqlw1Cv1PK+Tw4+lGTspSsIEHJ
7xCUXDgBupkR4ztiPjY81PCaX3NCxF0csJxvHkAFyNNijul40/W6RRCuJwGo
FrbGhovgoqIQvpKZUypG59AoJyszxYTHvWpdfS30aH0P3pR7AlLGyoXjaAiq
JukU9AY6hxEBxTaCW+BFKx3ALTVxUNRIn7dd4CryX631fhs7ZiBDh5rMSqOU
yhsnhEHGB84q4//+PHArT9FXU8etLKrMBkc26sYsfGAVqEcPpar4pf+WoPYn
UHmbW6jZwIIPySDaAT4HIlvR/6KCEAGRjrSsdKOB3BbQO+Xnoz7O4ZnsRwwd
vY7WlPopYhK9BJ/lzyE25AnmD6gpMjViQST81RC3JHH7UpVXQd4r7Drqq1Tr
CTzPCGIsCqo0Fy2fE0sitkKIkJNcZluAf/UotpnHxpP7nrLizAEGNDLRFbzg
7YSdcdFnKimBy4aPctQLjuwceqSXEW5cuT2WiZa5EoiVQ3oVeDWn+4536EcM
3jQwTWdWj4y+nSYfSBbzIzWa4LTZEyAq/GwoWwBTbq2R+6s2YiGL9fg6vigr
F7tWBUqWEQvPV78ITeFA7k3ziJW2R2QFSIxQp/Kkg0BHY0/UZHeNEicadkHU
nX5LYkaKHAriuySMAnZpSWzx8LRMUhzybNoj1ju7UhFiEoMBMER6o7E8A4Z3
Ba0fn6hmr3cxhJ+eldbt/YI+QvWQOOSeWz0wR3EfqBBjmoTxIHEqXxWG2KIK
AbCI1I7CvNG4vuPD7ojUWPXco273AwTNDsL61SrofEsLQUt29Hac4377hJra
X+K97dXJ46jSCULoFw86xGOvB/ApjAH+fXQmkgg/K7eN+NIxzAFBZSpeM/lP
hg02Cfp/08//jiUddnnp7zzX0MQDb3SwFEDd2bec2CTa9dK7h/omqjVgVPVi
uNv3Hoc1HL7wWGbE7ZulY2pKnzZqmZG6v0fndfsSaHK92rifCU5/FJqgd5Z6
FNY96rpVLY/99MsOMGiiaLRUc/t7pc8G0PnRAyoOuPkIYjETlZ07aJe723HW
Gpfrynu2N2lBGumREKRSU0PKsqsEHIocujhHys8CuCUWh4SyatxpMNgy4fX8
zm+4YHoRSrTGhnK6qvvx6VGqlr00I3KvY7f4rbMomSYbcUqv4AbVl+lc6nEw
UfTopegwYLB15NdTUXF7rJLWfSBnhre9MwKz3kPA935APWJjs/mo7KOoo05o
dxGW1SKsOKtgSuP5GFfL1s3K6Cc+VILwOs4I9vGEGpAb3SLvc9WRxFD7hr2D
HGpVnwbMlDRNuBpYc3GOR62MJVZqySAowNlFmpHh3zx8cnFCSMAE7yHtbB0+
yboJ+5+KwKgy7dgb0FoTegRfl/wmwS2yNBTobES+yg3uR0KEor+hqhz+7R/F
5vBaZLYQCYvjBsVxta2+N335FCgrqZrJ27576YleyPWmJ7d2RM78JOd/mlbG
ZgKyWE1gWct11IBIcmYQEcNOX6R2kWWEaEbcNqV2wZHkIaI3rq81vVOEAJu1
T88T5+yQTFpIN6ytFEsmmkH36ytOAkIchRr1QHcw9O1KRHIESUvZRJPKPPy+
6qDlnq6H35dVc2ZYAJrsz4Ama39cMg6Qm1DRiRDLnuGhBYLNNeA+x5MAsbAS
AzoNQx2U6zxKjbr0yOhy8gVncRiSvyjs2h4Zi1kIcbqkxJX1Qhn/+kDtNkNY
tkOIL+aFdHZIO47BGPNGBdGHoTA/NIg4U/hEqhO/JHEoEQ43EiFyYEC3c+Z5
WkY2w84YOozcHuNZXYD6ZqGf0WcFPx7hG99fQl9wRUDc66TbxD66I88ASICz
2dWep3bSN+k0u3x/BEWiQ61IPXN1v1HGZsoJT5aUDO6pytrD6d5VwaX8S0ad
uXoOuQN8cu1xffEfKrVzFwxfL7BMwNEXskYRebxfq5p8oQpUYfO/g0ibDhAZ
KUfEBT+/rcxW4gxlpE4G5+BTcTUuMdPdyWlwb1FpX1jInYoxhc6cIxPKlOP7
zNX7JtRKdHnpfkmwX1ggkGUfSS9P9Gx9WLiKZ1oNKlE+VcpnTeWWouaFo1d7
OhHC1C+odhu/exztEj6r6HlmDKnU95KqeuOF+4H54j98G6P8BZ0x46XkYzmL
18EBGUuI56snY4WJCUXjqk3oQz6KoRjIOSRSVywpFU5e0FFKNv1+XoBjVEEr
Wvltyg0DePM0Zs/BtZK6S+4BUWoMqDxYBl3be6hme0O0amzx9+VGRGow7K0R
rVoFkT4AMqWLbaQhDyre4Oe7XmB/uTz8yNtgd8aDMQ4rnj3SOqptkhBfMY+T
Oi7YJ5n9Ghs4Kgjknspvrl/pJdzXz5dMF28OrjuaIOvPmoeiPMQXJN+KJeEh
LbesArlEZtSIrmKrUgkKKvfPOXL/o1NiseVOnb0A2n25vcq/dAGeIMwArZ30
BoWt73WlY06Dj9ZgcD6ty+OJTCaNUhXtPyBa7aSmGwPNQWkW7OkdAAewzEuT
wksc5lKL2DCKEHW6wQ/oER3Yz6N5szq3vsYfcLy+Zp3E4PVFIRDacExIQQ4T
AIG6tfUrOfBLEkn0NBsQbg0+CfJes8yQPgOSG6lBwCeor6NR+zPnwYAlSWKA
vlsbS4SI0KlkeyebCaL2RkB5ve0xAuxZt5e0Cjxm5l5euAnFe/KXIpBkl1NW
2zCF9vw/DYTJZyRmTvSS88JSGblEQcO7aCcQvrlk6xyDzcvwmLak9z40blx3
mj1865gMl+pTGkPyxM3vax3ZEheA7jErbamZm1GSYAnMypWRC3u86zCR1UDj
fOLUJssyRmMZlezHZGQgKcPqx4GUQyGpNnCUbcg5g5xkTApgDrRTEh4wiTKr
IMRxwutdcD+g0XFqTCtMse7Q5pqvwCwnB34yrB8KfoQ6nxYgMor5Fe162PlO
0F/qD0ihSxxNh+6Ahw/GOgYjswnxoBnflCq9bddDA9VtUjuykT+Lb6QZMDOs
GzNM0Q/JZgyB8bIkKOUQfsGVCdIABXA9vIqub+mTillun6IMFjM1S9bzDA7g
DViy8F2X14mieGDSM7qA0HW8Vs0o5VQ8lbNa9YgSr31PBkpTedpYnqQMwnl5
6Lv4HgNE52QM+4+zLjysdZYXt85/XOD/QhXbKcI8kSbarUOlHnQf4HHdXW1f
uO07ngu/9iFLXuBYuEqi4+IdbWq6DObOHC/Gj5cJKuVgBuPS9nZscAFYEsdo
cnFfTvX6mpCzTLK2/UCMacyWisSaK/yaEGb1G9Z3KLzpVROJq2B5VGWN4yE2
WwUmx4xnjcWoLdqScm95fePhQrre43iLJJw/f4xoG9T7ihWgg9y/4OrOQ1A2
M6xQyzLpAcsLhLCOyf3jLzPIGLQB/1wREwxkBVSHgsnFvqMejktGpINP204V
qh39x3dcfJ7GuFlZ1O7bZ+lNy81Ne1UVGHrK/Fp1x/MsSjYy3J7NbmXTgAf9
OykjeNAbnQG/8UJTgC29dWJ4ovq1sckq6khvte5oUucxCqiTA7XUt64n52Q4
0sC3P90jfyk9YbXrg6huoJUxx3/Jxu7ccEPN9q8lzQmJtBRM67k+rtKQ/GPD
xVIg48JU2zmsFGULYpUNxe43rQZXp8fl/UEH5BzAB0OY5o2lVq4epqtlBU+A
VUyLdT3av7hS3p1tlKQ0ZpPETjKQSaHzPvtLVCGiuArxvnQjJFScIZIkc3Uy
m7R51oznzUgbJZEmOndNXIFl/hALapthGM9XZ/73clm/+RO2cTsfs/QMInpt
eFPGfTmeZnzfrC3sQt0VXgqfJWgJ++sSqurJLi160I4cVYfWs5M5a8bPJxxp
v6VcViNZ87D6t2xxpEKcMEWT5j6Qn5S0k0bih/MRoKgfCNzllHNAlpcZghfM
cfnki4POqmhpJASzcmxnHWd8Pr5gTOEBitfQC/tvr3h7Xp4qMC7cNED/D+Qd
Dh8ifeNVG+sbfAadC7VgyOe8CveNR9I5ls6mRUKIcskFuBQrd0GcE136P2AW
n2vnnv8unzTO5eb1/9/GIVfTUljTdSukeK3IOLs21ThrO2S2s3yWTSgw35fE
IKpXyWEMFT75cy1eWaHVbe6KEmXPevvkHa3aYO9wZgUd9codMBrB8huvb2F/
jdsBcGtJgdm3zffhvxGaIvf+CfitcPZumFmXwo0tF3UIEHGnglScO9Ux2t3B
2DUB+mrrqL5s14RtJloWgfHCXSNuxerbChihR0lk/8aivRG01pL5+savXzoz
6gR0iNK8OC6Vc2jFBMS7zKXhsD8evAcrwyo8d+Jc/hsZ7I1/hN/XQS2CHHlV
bdrDBafndGukM2zbqBce7jh6JTJmVsVyR5gYb/wq9ds7tleomW7b4PUNhPZd
R+jmF6T6W/Rz1+6MYFSzRyYKfFTSCmoOfY0YQLq4OZXZNBFsWWZMKwNKDSIz
CHXMVFU57kQNaMnhESitrY+ZCKohI1DIfZKe5672HoJT/hPYciov/YtvdMOf
0zF1E3Pt8/TdO5AAshFLSDhv7XXpW024PrT9NRSels0NW1ixvE9yNnBd0TM9
du5eIICYkliocUnZXHDDGc623p4d8IQjZrsm8QKWSIe3sX4joXUoJqMP6NrN
8ldL8hueFTO5sfu6yaJFAEIm4kb7Tw627MM8w8zsmFxhNlYbpHvJJqdlisbq
CtMLu+jfee4Cc9z8dDAoy2GVydDcZrqylHdClwRFcl2vXbY0VsR++HfyoYLr
gbgEFOWIry/6cZxiG4L5oQzdJYwmLg4WTOm0sDnqe4UYcugJzdIyItbWUue5
hM3D0onFinBNlRLsXAbk41MOEiKoatvHpWNC1ZlfvDALkLxt3Tg2mfhkgToh
e53vfLgaeNtiOZv5HonIl4PtSVQRRwB3LGLNoJLtUntw8vyQcruR3/mA53uM
sgqatm0moWXq4sWTpx3fwbsqtZvNUZ/CSYw3kHQXHxQq20gPlBUdv1XoihMD
18Yq/cDT/5rhIjVl+txMcyGq6SvmrRwBXvVLFEwk7Ft1PQFT8pQPHOf3mcOr
58Xw4q52/ujddisyU4Da7zSFGBzD+4OJMiFODwkW/+r+giRxDqvsdtJzjUVo
KFa1IEcuaVLoN/uU4MtPqdOB6LMCgDmu5K9MtzZoP8eqHJheRnY8TG5nBfIS
+ihO1c/NEeTe1uZXvbD5xHyb32SNo0Psoq+o9U4ZQafCF2o6wGNgKQqG0OR7
SDRP4oIIciXgF9L349HF1FheTvRT0djRPjL7AN6GOcOFIx+ZsrV46/ZEvxtO
GohRWDrh2nDnmHqZcyt5PanqF84hb+4x839GAHvducOZmIwluMOiijlIPZHA
P0IYkm9GTX67GgUIJqTF/XtKvWzA5X7cQcWTRkZBSFA9o35sT7ya1MFAk/DH
wcN8MrNmQC48fqz4f9FozVf0IQUvnC6T6W1KAk95Ax+9v5J5VWls3iBZ+3iL
7hxhAMxxYTlfritNnf7UDXEhzjkXTYpUf62TKyYxEthA22pbredwhAB1zFox
ynkeXhoxsyE1XEk5MyA42K33hTRAUni+pw++NFPXiqrRzN+OLILssdyOxOCE
g6XBESpCboQomQzvOnuz2wwMW1II/nDcKruegEmD0Q2TbNhu80C1pw5helaY
cGX4HyEBoTs+3hICHzSH54wztn78ya8i0MM3ZFJ0uOfEUllrO0G+/BXFY8UK
NDFQKcPMhkPam6He5jV9WLa9m/KU4bG5/2jEnioMZJWllZmr0FCnMb5S4fZ3
COPScdMtS2CJqzY893+6AQwZlkB79SxrChpxbRkMHkrdUQgqtS08JSKvZKne
ZWCAeSJxG53CME3hUzMANsDOlQ1hgkuZBd9WNlN1ga2OXeJLPAdui7HV1ioU
km307xiUdJDvgFIcXvDlyEdiEKj+7UM5OzXkuTu+JHqRdwapPg9h1TahmSrJ
h5bY+iCSPQjR/Oayl++J+tLrlfN9Cg6Js0hgKfcn6hyjkBHBVx4iVuisNEsc
cu2FX0qEsITEtATAEP4Acou3r6JJDWMJMDaZzIJfhzTwY8v2mXrzLXyTf7n1
IgZrwF5khSRA8XkPnVHZB8C5mQAp2/8ItJ/2dPD2gkhvdVHjIdy4iRcKnR7Q
pQeulZzXVA37Z1eQitlO3iQfnYTLuG1WUhEg0Zm31zbesMpREl8e/AptaORN
TonY4xfHL5SXl4cl5Lmeu3wkbzBAaxQ1RdwhhFoIoUPsrCK7MFp9RGobKuL7
O2mO6akOXGImIpTVN5kuh0MQeQUBnVmtJRDwR4Zh26b6/hLCsyylXu76Rqqq
eHz2k/B+VrzJt1hj3+4co9hxXub6Flcb4gj5BRYOpO5G+Ydsjt+QRLRm7W/D
nqZpElkjApxZlI6ZmVe4vcDWAS3u0ljdyDxFGGjD0h/neQvkDbbmOwXW8G5x
b13EE8vOU9odX220QUQVS0DhQ7zXe5HbmcmHebSpSR7dlYIigipgfjqLh8hA
ogMVguPqlbja2NB5sbpf/adWMKLGiwOIyIfdIUq4wLchykkG8Cd/a+80b5D8
1GrCkpV9LygA0UPDXrjhKkl1ppr4DKqJ+vx4/0y0jivT6EyBbUDtZpHZ+RUX
JKGeVW1KMLNo1yLQBGBRhpyv+kMhaCl9AuxZGiUq5Zx0+QZYO48UIDkn/qns
y1k93ZbE56rMPuBl312Ot1HpNwQtNRsFjCuDRUAujyWEUVAMeHhfeK/+xPmP
jVwR93+xYW1wHwB2YSz7AdnmSlaD5irtDcJF6FvbabyhO7df4vZoQYM2dLIw
rtZaLd1689cEuCOBKi4+cN19M1oAFTQWWJ3xJ2o3mPQWtcv49ciElFnvop35
Xa+h9jxWgONeN8uG9haZWsRYmnJce1NJ/61FlXWqfyAztOYnRpNVDA7umSd/
nCuLGf7dABGHjFQjG2PWHxCEyultzV7rMNDPFh2Kl5sJAwpiJAnLokLmJ1RV
TC6sHnU3V8d2i5vSDnGdD+xqHa4GfYths7crU+EVyGt/qwEEsM24YyEyA7Fp
dywL8LVdHp5fh2ZlQyRc/q+Lf1yDj90p1wqRQpUXawmlzZWloxMImeFUH1eN
f3wpx3u9lqtE8l2w/knE/nFfvmuuP0GaTeEwO7kdd++BR5aVSPfioWOe8phj
BfCxHEVmk+JPwOmdFRfg6JvHgmFJ15WXfBvCsUEUNv8kfuoyBnmG7YVvGRWU
Myqv29jralKSXn2/o5sE2K/4PkMxN8xI1UsR1PaWgtB53FivthcFhefCzmeu
W1NX1dLKadQN3dTV1ySgdsH8niUo1nN/AG7qaPUuqVMrqH2LPTWUiTglPO4n
4cRGgrx2lTw0sbG1zLG6ok98G2moe8/tNSGp0uiTZ4iYCCs1delMrp/NIgjj
5Ng2kbAI0PXP8lwAhv+ptAOUwO4gF8MXtT4ZAZdmHs5vdK2j3RvGIXuuT93i
mTFFbhc9hvsbepwJJs+8ntboCcqdlId4yhlaV565lgIgtDMrV7I2Bmk8T41Z
bJ1ypBUM1HYqM6liD5Yudlx3UD1QfErP3N5vJWK5KuXFw7enVQfe2CeXpoPG
I3wfvVtqF8gaXPTcMlgmJOFG/88w0playxNrd3A1uZ9aG8cmwaWBFY8oyG9N
VFScrzkSm9BiCvYCP7h36fmHLVZrfEEZRu+3HpZxO7TH29qg/6LfGWjvvi7H
k6wHeho7IeYb7Wa0cA7AldQr/a8TyxELknbt5u5nNJvs0tcOEC6jmwSWnXt3
5qZ4b1DyB4Sp0oAvQDB0PC7Z2nBe9GoxJD3LHPKoVmq2BVKBHpymQbud4I5K
8LBenEJCZhDrj6rRU7EmMAOgs9BsN9kZr78LzYVg6iFw9bTf8A1so8+/0sDP
pSozA0Qf1L2ljbmqCbfsA225DyOimniCrg18mHujJMqfvI/dN4u64obSF/EK
GnnEaR8tay15NEQZvy1SjFEDn0jjcB5xX/XU7mViuTDGANDg8BzWktPrqTvK
donJA28rCZngTn5t5LTZPQbTYJZUKG3E+m70wSd4vRL7AyIQfUrB0aU2SA48
q+UQ4dXajTGdRpQ9lqQR7+xxnh2O0vaSZEHh3OH0nUbQ0HUbPGQg8Kl9stA0
F7rYpDSxTKsGcuHitSCvriBYKoVeoDwC/OmHz70Q32j4crXgS7XxP3dJF5UT
LdWLNvT9SqxoVd2i6G4OiWGuugu0Lf5PIlNHtF167g4BfyV8Q5q3IAm+9r0R
rev8T79dZDXpQJi5tXJjnFzAAfrMnkG42R/51Yl6v1QXG0OyNmGNgqED69IZ
XZAjsaifH4NsDiDqFncGJrUR0WXIbZ88vWfDUZij3QrnzJh0qk7dqKYzDJKZ
rbIac+7a8QX4mHsac/NXBr+GTunuQ160luYcAkZT+63VXjQbvC4zC+5GVA/T
YzXwXV1UIk7qDMYyK4OLwP1M4o13XMdPdiGA6ATmG9SfAeeqXAnEaHf2OoK4
G9PDkX5sE9g3VIdBaoFcndPj2ABb8GJdH6NZpaEnKODM7x2AZlwhN/N9fQD1
EQvJIOULUcMA+FopOyUQSfvOrwAmWTvmZg2Y/a47DbWZq45U7uXmv+zlxmwD
mI+fMlVICNpm52a0rY47tyejN62LmJmJL9/1tKoMnP69+lEJ3bb5hVmMwq6f
ab9X5i7h1qrtH4/6se/61gc/DG24qVDvIxeN2/8LfoWgTEyZcEAjOPyIN9VA
wgNho7ytdVhCFtmk4om9HejUje0S6gcxvxQTn3685sTwFtk+igo8SK1JS3P2
CL/rzICp+XQEhhA5mUVk59zH5TyNAEHLZKXQqYrELkc9ybSRZCU/GeSApr2d
RGt4nHxG7p2SzZX4vchKO4386S0Le7xxAH3mg8cXSDmI+9SWukaj+MkC9tZA
ye4UK13Jxis4E5OzImZaKK7EKp00TmalOSw+m2dTG1XJFQIFtAbio76TmYnh
+bLsQ7jiqiUH8Yv4VFx6DPkpUzZqnFW5rjBCpo80LH3NOu837Ca80Aco8Z9G
5LnMog1BexYvKDAQmFXAlEchJKmgW9EmEbFaTHURWMEK3fDnb+PSqyw9PDMj
JccXR0a4y3hRWokjPiUgsb+QoNbl4IFt59spXfqhLN/3vf1OSw3d2ofei0d1
YS/sYPj+zLU1Kp7sDGBs8fgm64jcGk7zsdUcZxbda46o4vjAsozfVN23/25a
PGTM0JX5imj+qCltaz1HVMRtIp5KDSQA5vtN2TrFPNP7cHstBz9fMvJRCW2i
nT/AihBLIZ8bJQN93D4aPGvMbIiJ5G3tr/QqQOfeuozBTP/pcg4qrCqDNd5x
as5NfXKVSDnQCIL3oUb4iLgJKJ5AdFx2lZWHbTu/yIrrC8gTy9/xoRp0nP3p
aa/7Tfik9e6EhRSudRBrlNs2dJ4ccXo0edQzO9BE0PYwri49BJOlkbe8cS5F
dXMMSbnFr8OkFTMku0CIntjXVpVyZEx69JewW42VOGVQPVtIKnLS9did2JS9
SesYYawq6K5xfpkOkikW2PC94wcf/07f6J7Lah9IQWl5QT5T7hoW+QY4tTr1
AsjPhjV1gMxLge/9i4mPBix12SZfRFeGwSX50RheatrsztEh+ZfXnxunAc7N
MAZ75l7eIMHrt7q3pDzWj++R0Jy81dCLaUf3xbJTazv6yqyfM7miQ5ByEB1r
fVGMWWWDBalQPOnm28Wban9B8wsJHLhPXnclrdFQjrTdYucIwjk/TFW7OMEZ
PFG+0Di5FjQO49FxcCVbWEfoz7sNU5zT4oEQxbifV/UD+yJv6p4xLNJjsm3G
PFAnE4EmJhzDMy3oBXC17Dfd+xrmfRNAmJtCHtVk5HR+YFmMKdix17KLtQne
r+uWUZ+oUBI9yObQ0Xytuw5cEhRBJkC9ledan0KR0DTjwBSmonRrO/wuHn0+
4HU+BUvzz/R59Tihbe4Fi2qndTCAtlbno1LV/uRhqGfli01lqWWpueCvdOTR
z5CZugAMrbsXvyfFdCjsYPkg9FXWvvLsczEmpt/kcMBkfJvFct8xVoP3HawW
DX8hhBxuO1FYO6J78nKN+aPGBcZzvrcDf/INCIkNhilEIp6na3AAV51LE5yW
ZpJisDYLB11tPyTVF+nQsSpl0eiekpRhRWlLE4ueNnqwVK7uFfJ+oChbflr+
Zi0KbmLRcQcZXSGAZpFaWI/oWDK0R8COchLTT+5ItuiPx0LNFWi9iHWtkUGQ
5uUJbAwdvDfAiAPdZnEiKWlDOYl7hKkre9kME99IkF1+XlV6ctlV7B0IELsw
EoRCFLIT3hbivlcFMRbR+CEigDbNHK4wnO8YIk4YhBmf1Qy9iOn3HVYx1MLY
j9L/ECzpidnzYpDdT+z2L086B1anj3QZJl0cETY7EZoCpwmFt+WpsaLgniSH
QfQ0zu2rDZDYG2o/DTtuzQK48hHMo6ChIoDjsxTgTEZp4HkiP9wZDjUdeBvI
K1yfdXjb4aMqgxTPwWQBloNTPqAJ00rRxBE/ICKHS+pNAgru7TOWBpCYGqnu
8lrowXP1Detre9iPlE+lEGbE/cDueFB5HXZOQRHCpckrtvpjsSI87fBetna0
UWFuM2x7sRG60YY8UnU1Q20+myXDMB3wAIojBE7kknAKo76GNAdzN/HO/sDx
WTk7Ellf4V6DANO5a16DHp0tebVe53Vqmei2a5DfbMA6vrmIRu2xpz+knAXi
oQBRU2FiTmm9p2G/7sYN2ZL4yizNeGGkII27OqDqamV/Y+K49cH+8IPSWgwS
2i2oKQAH2q98lFuCzjcaVY74QSwcz0Knz6DIuYzjGPnOJoP7HUgAB/pjtmPr
aOH7Bnt7gX48eLOLpfgA8KOdVbx0HmHKpWbdoM0ZaIPWN/qgXSSo9/bBj/NE
u9FULRmfwIm4AlNd/O4vaJhcBPLN6H18VZzZNge5vif78rR/AgQpkQbk4jUU
lOgeOnR+pJI6X8Cu5vLBSMo7hlPHf7PZ9BzAMtl+nL2gX72KIe3BholfLF0J
ro+XjuZGnrmjdwrTmntHbaU6CErd6QqYTghGKaXeb6LwRF9aBX0kGiWOuVGm
i2KBV8tQ/FcNhghp/gLFEzyx2fWJO8tFFPLak+YlIEmIKnBjkGNxOCX4tNyo
AIF31AaSIkZldcq7rtHgHBBZs8zCpe7ismc4jH4ubAoUsBW1LQSCdvVck89d
oYAmqmmirW1VWeOZb68Otiduaeun/GOG7HIMxaOqGLbE5sCtELeRJYS2p43N
r8H1yL5Ko9DPENeLZRjyQJOB5cd7LXSuVM2gJiwuq7ba2B1v3BxtNkmJkO/M
jI4pKn+tTpgT6MyFaSoGgXMMnwFrYHkDafRXkjjoSrLGJNlqCdZae/uUGNjj
jLC8w6PNEAojSsVLG7uht9SVzYBW2dV0x+s0C+iY8Pkrk/qKEVGIgpUO4a0P
1cyfyUpOa1Qr4hcjFOMQWqVHeJE4FeSOWaIOOGRC0So3ZTXUA7yFTUfjO9Cy
VPtblVQKrC1di/28236kftRP+6n2uy0mbOwGjH45UF4j4n6sxxcnOKcRNLTE
P4icB6Lvw4WVfxzsOBFNZLdKf+4SnDLMTPAgdS2Pmau0qSQpPwhk9QCc5LBL
NM8uMhhChHKTdn1IjwHNQEvwdU5pklISZfwSMLcH8GYPNnV3k7ZgiNBjctWr
kw9VwMI1CwikRj6q5rsGLxXweMUoFHdGb+kWepG0amruNvKchSGIXToNz6j8
BNTdSo/RckzalJbR+p4/bx5U5NZsqjasVOq4ZncnI+sxwhvBLG7tPcquiQ+K
NKTbFYoOSVAsnZNVN4ANLqYfJUWZkV30D/eNbk/fKKoVscL5CCLF/7zkWgKv
OuWaIbYKetBNARywa/cs+Ryn2fr5+SoXD3RSilU5coTG4sh/eobdgWoftWG4
9yPD04LdNUmC0WCbW+Ard2hiDu1a70cKexv/YCJsdFUbcjM/b4Xb4zVJgVpW
85CHFnsHy2Dr+cGqwEIu58IP/Rp69W1VgoNMxXbdfp2M8LF3oWWq6pDeKu23
noONq4usx4w61vowafosOnHHaruPHhDUuxdrLizVuwEpLwJHIc5vr9BCBiLO
rbu6JiEIMDzZ741s6fMeTsg8pnsglj5Jft+akLkegikf5VjMhatjaJcCXrJJ
ZKCc9sprmRDW/Vxvaft7tTFZjJL+RIj5YGw0dxLf8FY7X4DyMU0XmalkNbx9
TnkNStnEudp6ROT9pq+9SmopVjT9cjokP7ZpaYrLoRELHID8G/OC2uHVX5PJ
3YWNp2hE8WoVZ0JQnmEeSWUN/xTYM6xXpDQlg5EKB4h4JSWcYpWYgVxQRbav
S/2UbV8glGnE67wOrAU5hIIjho/2Izry3TF0mQZ18f1k5Cz7fAa7g1e1XWS4
y7Qqm1/kBghWZ6w41o5J5Ox/pQlFWnEHsnRG4ApBlR42yGmZ+pOq2Fi/Q4ZV
121Lord6mErGCrTMt7OSjmR3RqyBgp6yE8QBofCdsrnElYKNneOpLyJNDseK
hSJEFk2s/hXNdGgCkdWlXwAjVDrLX87HWvJHW0V6iP2+AxdHmTRnsMFFUHgu
Wbhp3V5798UExvwg7JqzISIRTWUhxoFDFXlZtcitIsDwfqjaVt9k72P/0A3T
FoZYA5YdDwg4iHYw4erxZ8KTK5kCkb5Q8kfCWlFIYTZbfabRhW1SR9bOOdWJ
wEY2+3aWqCsAwf8ANO8Xk1MOGN/qd8kg0YZoZOp3I2uwtGBUhZa5RQeYDKcG
oguBwT2S79j9qRXVOs0ntX3nHSZEk2IXKoa0Tzf1WOf1047QfLa94ROI2TBR
aaGe1LVVVBLLMYdUIunYcH9PSIt3iiIcdJybRS+uEksogaD5RF1qvBKOE/bp
CZFvbkFBBYmni7yy2M9eWi09UNcP0h/5IkA3PX1wbUY0t3DqmqwZC++YU+HQ
q8AOnkJGM+TIVT67uzbrKo6yaNsPKgps9sxKVYMsk5VA7EyH7cCjd1N1Rdbo
UmCejk9WEb8XaLycoI/QI6TxRhKxmG+Fgzw4/Y3Zf7vJq5soLJ0IEavMa4o1
gkbl+D3jUndcyb7HHGCRUpxjiYGHJ5Eq/ebMoS7AxBtSSQAQMk4HnStOInzw
OPHwyFQBk5/qezHKDkdaxj2NaK6HiGHva15XZdeSkXBim+XZaq/Jkzu/LQcY
PWBlTUL/yCMW2Eu45hRWh0gMWooOGEkbxMy7jBp4WZUFaZ3yYBAaKu13/GV7
4ORqV2HYJ5qLO5kL+ctUOoOm/+PfcRjPDi+SK0UhDmUq9hVnNjd7qvdjkhq/
QnLfIXqSEBqU/pSSNWSclqqSeyvR/0BWkwxekFQQi9UgR2mYvuQPnKkuNiOH
ilaJyQlRA0YhNJ6fytwg2dZ6HVPhbiOkPVRGcK6txjjAeJgfHUnpkMP2HKY7
WVe9Ti7TXApWBNZcYvLaATtDEcmfCXX+OWxUGyKLUjRCfiZKytAV9Aka/Lze
woCCSREXd6qKVqGzPOw68F+kDTlDnfmE39Rjbd18TjyaT7kGbRwEM8JJGVdS
TGP0OMLBJTTWK0PJH5JTEBNqv7OnkV7IrPDI2Ryce2R2PUOKWq80XeS/lx8f
FYrPsJXB2Fhz5hlGm/2p+UlzWQL3HnuS8jA3g5pOJlSwAQuB+lJaC6l/S6I5
GJ3fdi8aZJTvHIGaO8Xn7HRWdvr0XtVZZ1udKbe8OI0C8qyFxR7guiswlNfr
W0cZTvH6CitVgfujXrEvJlIZVCo1I6DegXCJ3ZclE52fa+jF38Mgjp9MDH7U
H5w6Qu/1GBHXulktMiCEWVEybO5EONPYuPhAn3c25+uJ5C0fihFKqGsofMe3
o1S1CnZAY7Q2f+jUyqWlyootcyBajXCI632v2nKUHgcUZoQFoVjEYK1VPR/1
RwxkimUdyrT39/K+46P5jdAtu8wza9M7S6H3l5+RRpOHbhWeQOOc3eQR1KPF
BGqr+VX4RXP3U1ssl4fZ+DwPjF9KLAEwx954ik72j6tYzW4B3yYm8pfxXEvJ
3jPvoqvCIb0xShNotoMDALDXtSphz9S5srXJwLLM8Suzl+8nBO4a28HDOByQ
EQ/DWJsYaz8dHbGXL82wyhxKSgMDOh7isXMy4AVCx8QndF9NPbCPexlvRhcC
jcjJ6Je8o2D+p+qLWV4zGwD8cnnc2kT2qCtwvKNeLT5qjWQkEkAlETGY5CMP
b+LUGinB+XsCsaywSuEXP9FQX2BGEegm4NGWHtLfg6RnRq95dVA3LESLjXmE
DLrSSkYoUAl5LzPDJGMdgOYV3cDqtSrhj1eonjMcrI0RGhpkpu80sFx8yRL3
wtH4JUnhvmq0SCBdYtdTrpAVKekFOu63fAvaSvjbPx57R9NN9LJkQxSt8rGO
EC/tqYF9GCb4HHaq8x3SC2z9cJTWOgV/0GKhviG6IJ+dQCpEuoAOvWKYsaB2
UrhMOrRl4WQxySyAV668UMuISQVW1ptQWfGp4muooEqgvkGubm3ecODb+Ej4
NRIFxJ0dQZhXB0e23wPxHWeRH6uQhYL3b4Aw5riVPYClpax20Mha6/YxAr5u
lEbYZQ/xMUwh14Ful/hUlMA+R7RzeD3vDrU8Tt6zbvFdOKMJ931PaGE2wliC
H0zIjlgA8fEYm1bdgnA7JAzc0n2Yq+fbIsdh3NO8LZkSw81NllABlPaKDyQW
7+spwiV1NyBK4EtEsQ3FsDvliFmU683hrBhf7H8F5zXAv6QPE3jgb2sd2XhC
Bb5qlYYahmVvWA6tLuW3qjD2WDO/YXyGqFi4+YIN0L3UvyUCcABs1Yc+zvHv
Q5JVBOWVK2CcJwL8qmR1LPKZCXz8qrb5823Vyo5XvdeBJrtNNaKqhZUthcwQ
/YS7N4Nq4AxB5uJ+PMJ1vT8nQvRo9Wv6BhrD+2V8KV2e8WaJ686S1OJ4eAer
fIhBAqfMw0N0ARvh1xg4s6blQnr2aAtr0a3KwWo0uFA7Z/LmUaQJ3S5w66QY
PgqYnANwlzz/q0Oa/UOEl/uQXXa4gX/1haKWr1O8KSJV3eOM723Q+A37bLRq
e6nUiAvtsfBnSTMeEtbUCDhalshRw9NQSYv0d0p78IEsVpMQvvypECMY8gBd
crxwFbWxUsLqpY0NpIPeluPIBHUBTmD5XP/3Cb4o7OmdqMi+JDdoNT8eMFAT
7Y1A7naveKqi0yHmUuIxCY5ilAy0grjA1acvx/l4VhDCr2MxLsYQJP1/HXLE
dXFJwvn7vA39LT2dFxEWhsuZT/mzcCb1yRX35X0YvfwYlALtHGODgbpvgIFy
DKjJqP5dOz5B8YAP3Te3GYRvMQIzd3YGi+lGcfbVrnvjyu4BAG63UDaHHqIr
ozwXxSOxi50T8sTlIKUbuMmIlfdp7aCFEgETrrvXA0T2qT/Ny9ENJgUTTW23
ohL4btjuzmM0iEw/v6h0QcMrU8/PDMNOtBIxYzYJmWUoZAjAc84og+YNTgLm
A2SpVyfoE3otsZkxwh3NznsrSY38n/y449BCnqijOpqKCQRzDnfkZi9ks5CX
zpvf66dumAl8SOYO8xmF5KKz3Cs7XTE3Xh1sv+IEMKgx2XrJpmwosUeVXuYF
J8UjDGvI+XrFQpAzebRubbootQWKvhI21JWUQsh4XV0fDP2FTkVd4ax/Z2Y+
Iz1jL8QTwtq3wxIO9KEd6abzYt7JLSuiTmzwVhuskHkclBjQ2FqqpTGjSXCU
VtQdS4mvIBP0KtfTwkX22YW7izo0Gea22u97DvbVEZAf8DISB0udGvZ9d7cG
3YrGVY2FiPETW7XKNaZS4xJjLvbhhb529+XWonqMZ1hP4IuZHVlSL+FpymXg
WB/qtvHPeKZA31NXynaaL0x/QqgJecJMLKP5no3PCUPMxrBcimd/QKS8VQiP
djhSQuYAlsLyrYhcOHCmXrZ5AVmELOY7ac73WFuxQc4/LdREKuT6o3a+nQ2j
kL4YbbwDz0IyxANU2NkjOLLIA903/Y7yWRvBv9dktVQZ8EDO6fs5rt+x7aMp
B+eTN7zuERNPpDw6ogJnCrfDrSK0f/ZE0MPDWT5OsBXYq7y9MgCfpY7QzGxZ
/Sk6YFziCE2oZr4myM5JEFP7HqeJ0qYWp/twOawI1zeJ5CJXbko6Nrj5vxNC
u+GrLQ0bRKP1DvEDH1S2l17Gw8CXw2UHWKaWp/EzrXbrTnBe4MiJedxWqX1F
+sweLHrYMt7f09FdvbW3rrwAA1rqjvrSyIj8EVrN9o54cTgf3k5WjmNuBkM3
WD2SHeHDrjD7RKvIu5fPLn/yJJBh+90qp3HUB1i9ido11ChP+H5bVQOwPJl1
nA7rG3xQzcNATizUT0zDl9/wKZWA3wq+ru26rAOgtVmislm0lq6d9ZsqjDCj
idanAAx4iOsKojOy+Ue4jh6raCZ88ZnneM/LsTwXG6PGA1p0/o83wnWCN1tV
BeccxisFmx5TVq8G7LXfPIaTtESGlgHflCKNSdVqJiSWDnxRc9nbwO3RqB0Q
6rKgkXWmfWx9sG8pv4E3nLx1hp9JTst9Od4+qmfMdsIiSYrk9fvrMaET31+r
67MH3N7+XBOx8sKMNsAUAFO/as2pfOHGN6BrLBCvItix7/f7d6lMWUPJP7JX
SQKJu9rVCxUZjA9i0+hwgqqzIs8bhVpsCyGfpCJUHi34ctshm0GKOxhs2cnV
8NWkp07jQM7/KvtMCtBOH7pRQRrqp8WFfrI989Ox+ZygbMSlSKAkXwnsUVez
RvbB0jDq8fbd3R6qFjiTm1VCPgZLc4Y0HuUfam62OxJnhK1pwKDd4D3NsV89
XIhzwewLuinlErFcNrtYmtLyYH4/0R0pzrn/oPVDm1wVbc2nohfAezFBw22y
HAezbvtgKSJna4H2t304FbcU8nd++z5L6TqOeS2pYSzYt/ipaYGj3zanGwEI
3CFjDqvCO4vv4POj7/HT7zLQN5LKG+haXMUT5NtOK5jnlezzwh8ObUnaQb00
+YvFns7rM7Jj9fnei/F6hQ37GDX0Qcr7Nk5oNE38BNI0SiU7/VsPkDHeIIXH
zBsTnytOuc+dSLYHNedVepsgmo/zfvzpiDjlxarQK4k70f4S3gm0UASckqfS
qBNXz+1Er+9RPuwpjcvMynJSMZSGkPuJ65Ij7T3Gdd7GYu4dP4XaaSyVD9gE
DpwQ7IddTctUJ5YAs5aBP86nEGN/JcJIJ+OEDYIIFxKGT3lHMWUY89n9zsgg
l5D/efr2G7aBcAj+nFCo3o2FS+E/RU4HEnPFUfgMTnD6m8s5et/0AuGlbPav
o92fx+O+xQEdvrsiIXco6f/XqXpy9AbKLPewkWTd9KAH/HoFQeoW9sjGJfr4
68l3Xhj5MRhg9rsUNoPwgFBkfPTmgERvIHH46JIJR1f5cctUMxZMyjzCGTRV
XlYxRAdVC4BhZ3UJsHO75gA1EYAd3+ijyP3zZ7SvDE0sctGhSHf3RGVutR/7
VbWqjB4HoFNAnSMrQwpNLDXPMFoZui5luC7cNV1GnPt7OEi5mzb1FHSeyAaw
2S5PDWOEWv3x1oy/lKAunA0Z2dGScSBz+6OED8fUXl8Bs6PIoQEx2DDFeNWh
iSltzVT/jNbRravW+RaDXODV3CzZ8i0ArDZVJBafINPhdz+irSOzpef2+26O
N20TYIlSvQC9rUNNM8p8MHqDvlR2pw8CfBL5dGp4M+s+gMieR7RRiHGg1WOo
VX3OtbjhL0Lp6+2rXhSGOAcQ7jUSUixOv8UfvdBUmhEjIKA/DuyTlr/RYksi
aYwbpErd8rwdUq5PlVfQeUuD6KuawjthseiTSBqOWjhLOc0ikIuldm5HYndv
Qz/g9Hs67zVsPhtSIthOMHckguEcUlBgnW3fDu/Ua0YvgCwE8OBcF9uUkigk
EXil5C97TkUYqxn8x5EjlslUW8k+h/z1Fj4UGmojZgWY8VjC3+5TpghNKFwF
cNJ8ZO/9QvMOz+NYGs3xnkdTDws417FdgjBWukmt0cvjTqDKGIDn2YVWHaeF
QgvMLR1Y42sE6YelKkygyNgpXS8HiLVt2tinf/LFOqJ+kTTVpv3n9rrKdxF4
7TPp/g69BqxNQP9qH38I+sbzr9LgCrkiY+TlPEs4FMW0jklflwpVxZNeQWKx
lZhu25PXS3RhPiWUpR8V9eutVa5JufrnOG5zax+tuGju6ZQKKPdMyTZwZid+
jraIdFTwgBxwLNmeu5ldR0OYi2sG1//4k3YGHa2KIqRpGZtUNJFLgk8ySYRB
iTmhibXg4Y2hjKNxdKRj9ffCtaTC2gUwHJQSZlVrOpNuRl6+/fmTMD44ddkf
g28Wojj2NFOvIGhUdcEVn3arYZo6Uoz3CSuhjO4wSjzxU7HdJgPkpjVqRvt4
NSktlMgQoQm0DRiPaNDpgSzYptlJsOuTidCqW5S+D9dcyfRyB65zCYfIohhY
hzwTNKldKY1i7NAAOVO5NgMIeQXgz1Z+Zt9soZMOV9pkHEY9IPjC3QWEZgeu
+eJvbEDC1AknqjMhukOhDXccEDCGYzx7R1YhSHVT/07/H+L+/c00faZASLa4
rQ00m7ZGUpvzmXd+DBHa4KcE6u4b23f5fght38/XBHFXBwN3EuU33ReSM6lD
ixcfotxPLKfH+WwBgDrQICO4q2M1me5rilLYi/d/xFZdI+82yL2UNRgFR8aq
KooNmSFypucyXXGUGo4zSiKBywxhEw+VzsBy6yyAJvqnj96ytnRnDjyQfKU/
pPrB1nME+kYcg0rTfbj11dWklcoUNV2Je54L821M1DTNhiXHKg+0rbhsFiWy
esvwOBuj3fpdIlL+eQ1PdIyI3qllh7iDKxUTWAhUvi631GKQmb8UXuV1sFJy
jpz2E0z/ntek6ZNR0ug3poI9wN1fFzFqeefOy+Uf3AQighivWlVtz/0eHuXQ
7hNP15dYqaD/aqeeIisAxAFS9u2Rh51aayjxd8m5HCm3y0Fgqzjm+JdtZbkM
NrniyqsKOL45iyl4lJPfSk7/DLigqIN0gefEH0UzSAYCmtYkFJ8wr5qvnCOO
y39hZfaYYrG8HomQg19Ypn1S4GbIhXGR3xr0LPFVmJqMZZa02QwU0g8WUZz1
q+1wwaOBmSWzBIacBjO2xIJAd9i9xPX5aO9XX644EVFCISc4fi1eJBc+M8qP
8dXfF7M34v6lH2mTFX60H+GmsCiW9LcnkgW6cGIliImbStqDXcPFyvhvPrgP
sJfKX6e+umIlxvO2jxQMb7sGF9EbW+QIs3rvKy7HjyrQZ+Is6aauEHPWAFMy
9ad++l4WcwTl3IJe9DTMnAHxcRoeJdVutfzWEXgdU+LMNSpVJgxRd474TxdF
XcE72DPtugE6JRR9vXaBdWImfhko1rQMU4+Uc89BW6omDRftMKGpJO7vbEJ7
4G00FROXQOmr46vcNfv2sadDo9986+myS7QCdFkm2Oe4n/YNPN6JMBokao5k
8euGgorf2aXvXpeq8j9E3+la13HSAWY2F1KMFRf8LNxnHNEdvEPk26qDwY2N
qD8Z9y99+X/CfqOoquIWUwg/+FXLd62NGLfA9p0YomxvTN3hLu+/UcuyagJR
m7BOb9qqx0rYA1bMPgAbTS5qQscJe/t+3w5uS0Uodj5h5Np21HeZHtn4dDV5
GC00kt7IsrvOnVktk5MfJxERHTpmFrKrX5OTS30DaiCpz1f8fTjFCrSGBN5m
d3JhsQex3s0tTkrKzYBbFLgQLGdqE6yxEVqp5406Cs4ftT/LMLz2Ytpn5dLE
mtbYlcLc12DTFQ/WePTfb5QM8dblJRIbTsEBZCUXOdUXc4NRy/7KEDHFPJNc
IQSucNvze3jDnungthtKUTb7DQFWS7OH6wynuKy+p2PieTh8C9LWsJ8M13p4
FJCZJYDUzFmVvg5mI2Y+3oGZ6JtCwuHBvmJe4fZ0P4otjy+e8SU7W7qYxsFC
yrsPSldZyNhKts7MYXMyxzcKJYBkWLfoV9+Td88ilr3HcM4U4aWORJtbn8Kp
3FG9j8LnB8NHjYFA22q2o27FdP7a50cKt7HJvlvKzn9R7YHifPuvxuPnn51o
RNSzKOtgFImdQMT+QXcZtyXT4gt/zjYw6ZGp1d7JLawzYHym7feg2dPkAID9
PMauvpmveH/G6ybeEKPPel+YpixWtogIMC1WADx3znR1fQJ2ZFjSMbK6+oPz
57LhjDYfHkVDiqOtWnoJ1eqKYvBDhssz2za+XVHQTtNj8q49GyJDDmmkyY2T
7ep1KT3fTcFEmP4fxEA4qM5vKyjrADtTGpSksiZbu8J4QhrLO0WbZIFlJEjD
DDq3ZMzEZbpDHd0VXvU5rJF615T1d6pXZtRo/FIcH9FGsvY88j1jp9zjhEZy
gHQoZQ7d78dqvLL00DC4YaqKPHidc7wEkS4LDS5Sd120vKzOA4OGsfkx8keN
j0qA5N9U9oNXM3P5sOvlVcT9Rvdlnsn5WlcLg53d8aSkrQnScpJw4Rk4Mv41
pCF+6Iz9XW3esniFXDjcIfP+JW7ckOQvQZ29or8ucvFcQeQx2BURbtu6DDh9
iTOUTTcqjZMj6aMfWndD8nyygy3nUGwbHU42Q3p1C3LL7wpmfpTEM6rwyFFi
ApfaHR/2qhWbarwvse9cD9oIPKroOSMK0YB2Hrikt1sEVbhhyk3aX2K+tToO
0u7HI6iDyDWzNvoOqDZ3N3cd+0R00G79NGd03N5oDSlsHrHDtNxUDP5W8q5o
seQ5+stE4UMv6IBRYsjbD9NlAddzApnzqMpEdWdgwpPeHVc6sVnziOapttJt
SGvBf8keU7ou8Uy9lW/I5DNZ1pt7hfZqxuSjMxUm7i83CRMoem3qWIKkLQ39
KOO/ZNJm3BV4qQfVYbwMMWJxGSF+oWTL5PntBNFpTc83nK5ctkCrfkMNkN2S
+G5aYwtS7k81ikd1boL2cjDR0tNN4oJwGvR418kMz8yWUjantj7KS1w3RrEa
pfTQW1DfqJRSNPkcW+QKOcbjzC3O++HoSTdwg5guoblnUleRkNSAPQHs9SDx
JD1tCrGz1SCOmnQ0IkdX4KYhKZdwLpf8cPCJbN7kgJ+iGXY5nj5xtW0GYNNS
XZgP5ep4F5+0HHsg/v0unHog2ac4apnRBp4e2RkxonTiw+ZpEQ8uW48wFQlJ
CqRVk9l4FwRaVBmfqezJX2bTG2ycnMFDy1PJxE/ePVMg7Uvkw1OaWiu2Hb48
IDv54YNoF8Fjzg3oYg/oqlQ8s3vtEeJ2CKCA8OiWdJT/3UPFlOCq2ULGiGhW
TnMu5otRpL5RLiWHbqWA7LDpcA0khaLS+uqAKu4UJGTxHHeZcgoK6iuAmljq
chGSC67qXrGLpNnCoK5oI5NXQ3/AwFRUc1sPBjwDViiQygcvlI0uO52b+7ca
6djwS0p4RdAiinhXo1gVqxiceAxIai+jxJ3EVt2hEgkQIsvdWYa1j3NdrBVI
lq14bPA1soRdoF6sD9fAr7BK0pd4uhC9RMMZvEFOQeiw/d9swSUTl2MUWJU0
3jonasYlYnIIt0UishqS/NCpsH8uQIBEwlikM1/bA9gPje4QTdesoSZ9XsVJ
fadMwrkFN7SD5GT2UIm3LBz4qGhMqwA642aV2rqAsGn+qsE6Oes2iJsebWIG
lFmr4ycJVYuWDb1qGN+HiTwQfgA/4KaUuUQEGe5LkHYx93l1/o9PK7pcqf7b
gx0qEEfzUvUXG0LB634UaMBSxBdgbxvD4TzL0xxFnLw3yAfKu6tAFEbLYKU6
0woM0xYL5VRnG+EDeJlb2Y2JvvWN2jjIOJHvSdpewRj46rSR5XoEW9LnWSHK
tyeeWPGke09CI5T7gRK7u3jf8BpDds+LYuphXjBhunm+KbOLA/ceA4mvV4AA
78d5kvygOGWDNU4Q7MDB1gKYVC2RfNoNts4CPpU8Ak6dYu8uUh/U17xvj8S9
xDi6kRU3W8UlsPLJNgr+5WkWRsMKb/U8VFMMoum69GG8obbWjeftIoFywhrc
k9fHgqzVZ7vCCGoY/3w2onGeP68Vv6tM56vw3W+ONgtUJ3IA7QBYzHxpWl1A
Q0j1yTDYGoe9WHdMVB8ySwvHduUJt5v8Fn2i0VUVdlEQ9kV3HNGo+UkceoFQ
6p/Lr6FSTq7jjYEwP3HT7qtMtWAy0LzhOQwXWZLTJkRTEjoVN0X9Mk2uzDX1
IX4rUvX4lx8T7qqI3ouQGfq6vfVm/5hnGBWvLHZnenn7/w2AhTvf6EPYBhFG
Up8Nt5hTdQucetnK8lG/0qZhETuRclopBarGF0U+Gb0/NzmSJFO47RqY+tzL
RyCO6SmXcUV5+pei+gw3QodouUb8JXHMP1wCK6NfBnKYOTxMbvN04cyyEd3E
6unkca9/fvTLlXI29rBLN/C9s3Cz5FxLNSw4MILDCelUvd8sMlM8BtVZ74uD
4nOBzIfJrqgup+jZ3OxH9S5ZtYXohbveiM1ZGKzPkEfQBPBiWnoGxNmYKe1K
jvp9wYxtiFa6at2mKUrSqjV0hr92tEaA349+v91xAAejYoXi7JGC9qJY+rx3
Nst65dh2icJW+G0MNITr0Nlb4VpU2u0mRsH0yYntQpIMs0Hp16JvODefGJyl
SPzBbswttu0fweHF6O8zscvC4/bk3/W5+jfzpHwYKjvPIGkKexjYTDYGJ5ax
81Q3bhuoXWTyWUy0/KOJ7mAUqVB7HX0P7a3Vu+/jOptARur2zE6knhS61OOY
n+rvi2OeWBgaPuS4eDV1MZXh3AljU/TB7BxJnXoBP1wDiM7rpSe+JVv2uY0s
gpXYZDxIMve6rc76pKmR3PdlIttz2Jp4rLgZZDnTjE1tUilBnPi7c4xcfj5B
TPBvl3VSxfLwCWj+idFWYE/prQGoVRQaOyqGIiw3dCXwBP5Py3xO60BLgvU3
WoTwKCrtUwG9iW/STgR0sxbpLo29M9rJNzFAV2pZilxkJPAEsuGY4rvhS6Po
0/RCxclRCPQVpUvA10EeMSYFomvIii40fVLhi+hA423/jGuOTz9sqO0FzSEQ
YiSP4K+pSLsLIrC5hK+RwC+ghO11qPNwiHwt+ycMzVMs2KwTxRePWfXJdGX1
pimbyb1UflVfTXPaP5FaSC7mIUdXptF3UhsKB89Q08Uj9vzjGZBmM2O2PW2W
EmRqOLRMwip/bnKhqvbrWdCruM9Y5n90NPRb6LaTn4rXmfBzlxLt5vi6tJKZ
mefZXdMDGiCJsr+PpkbX9tWepryvJuaKhpsVTdDvLqaJpEBGGwCrcTjw+7Q3
PROJnCS/M/ByvwwQXwBmNs73l1QnHqGyQ8muwzharmz3lnJnH8zeibSvG/CP
APVnLE4RBbABfwbDwFAvjXcOKmbx0j40xDZg46w1P5GRDhJloJ+93XArcKa2
a/lwOwneDH8ptQsixmjJ22BkJrCSugtJraXWMjYfyuQhg0ImuCvldD5DYSLU
qEq/Y8E/qN3r+m0OVLzPI4jL7Q4obD2NISKJqji/CrAKDhVPy24RPFcyehkk
ah2jiVvRN6miXQR4zWGr/Djw2KA0PVKGTNGCQ733emXnM7fO7SF2wtGzUczJ
j0Sv1QbtK6FcWWMHpE67zBRvtV+tql/a0vGRdrPy90lWkVM16DN7BTIIkozA
s2inbf9aCIAgqGnso6JqpBtJ589Qqrfn2eSX3Ky7B4LwLV2VwG2iSwnw0fZI
JIYHZoE8Nt8MbPmvHUt7zpiHHyJ62/yHCFgV/N935UNWgPINiUY44m0ctK1q
j0/mktgoXoiaujR5mi9av0Kt8EvaRUq26mxG+OQH8ONCA8Ogv5lkuTbszyAq
JuxvpocAbPsEeKSWrYeRhxQz97/XkTUg8rc4+FQs2gyitfwuK2EeQIQ1hLo4
MTod/CKvps5SmvpoVYbm+rm/cGZBJ5VZ19vQAQly+H5rkgsFopVLjkDX5Ha4
nXuC0yqw1E9zzfyFWxhEELbzSu6/0XO5sSRUlYVIxS4NJNgEYQtQSvgRD1MQ
ImcevoeXjIVLxAxkYthtQASr4brqagLkGiBwlMktRfFIvJdmOq2lsKiSI6L3
YzEt/eIizkjODpgq0EraVIBXZBj4pSZ668NcZwKkBMuMqRJlHMfRTeJLkOOH
2JwAyXqb9guXBcFtKSQIrNVAAahCiUEvLyuPz8036zxrP6WgIc+Vb8ktUPXo
wkwBfArwCoMfFN9QY7LShirQDSBNWQC+gptUXRoJyL4nE9n+EpznLyH529py
h2Sx4KyN77U6rKfs63QsSC+7Afc+X6GnrPEXlerACYnXMjDbV7AoDVc72X8S
6VgOgfBmuIGhEuw5eSYXIUYnFu3ZD/BFkdLpMznaxQtvxLb2mjkPCNdV9He7
jOck7pVa0xooxIwH2ZL48I/D51JHO4L/ZWnew5jYyYmRZqcEf1bpTx3K7Jfh
B2JjmDR3oYwTn/nn6S2eTxcmlZxArVatru2ua18ekw8L38y/7xomQNmIPbQ4
2XVYnMnAyjg0jaOEiIns08kKdRg1Jw02ZdaUuFxRZPdhZiuFXxY0QCa6Qlvg
/eG6+JSjh0he9Vr2ObFif3nZv/dxbpp43I/cx9HSuCts/4CMWFB+ewBpPEdd
TetsRSprFyFMSf2d8VcSP97Go06e1Emwhh2NL46Wt1Ca4O75nUWzf/updsgu
mWPzKDF/vzmG5XYoZ25URq6UE54N95x3ZOgkcWgsrJgaDBxGEzYwpyv3UuJI
oKTSfaKwvd1MP8+yZJjGNm003EvbVeny0E5Mp70jC8J35EhAF4zmxLX6tDGa
5kUJbGRP3FSfmHIsF8TPTzCtFvJsu2wN7alu/Mqe3vC/EsSMaWg0WK5kFm4e
v/q3OuBhXYLkS+NfVdIIIaS+o6z1yNJoGzVTku+CBZ57P6J7XpPc3fMvtLu3
wHsaXQ4yfuqQmFYnMw2iqWnJsQj5w7kODp1KEUxDT0ybLJ2SXPAz6FkfRo/t
Tw7WwVwxbbqIzalPdgdToQHacXP5+ufdI+rhq/jBPzkRNQ5L3oD1vRWuF+F8
5GTV86oA/tAMZtQ63MtAnMlNgOqlNTtXT5TaiL66Zx+4FA8qnk1TxS1HRCR6
dq7Q6K9i5HG4Bfe1zbYBxgCzflJyAqAA27vUYBAQFa5LWP9aCA+DqEfQLpxU
A19YKa5jBY8UWRKktN0HTXcoIC+zFy84AJXJwkvohVQLPdfYPVh2V3Cm+SBw
GBl3vTvx9eo8m/ualBH+sS/pfFi+kCVIPdoMSUjSF7/616W9C52FsFPKwW5/
ukm96R/rElNHYqQN7UIY6paF0DnkJI/wfCDycZt2/bMAnnzPfC3qnriRnGET
tKq5g1GQDnz0RJBhDfl9PFUhH7QqsGnwZrRFb6iS+HP9kUJZddzGhyIBAjzB
QqX0MxlluT7ElJ9iTTsEfcSzWuQndQZ8uIngXcgvGOPpNj1PkPsRSa4VBOoO
Y/KDWdls1n47T4XoMZfBD+PByEbmyhp0yJRr7vmFcxqG+KXGrR02Yl7NBW7N
ZqvjoR4VVdoPyZcqzPTY/0s+j/58Bnkg0vzgygiga86PhmCd4UKYJ6zYn50F
e4hIkzGBI4GVRzcl/weS5JqBWkagTRfdeQVhJpm3ocFKsFAWaONjFE8qIjlS
m6aiMc5rDTHln0Flv2meRtO9ta9/cglfpDBJrHVKXmc1txKlUxUU5giZQCjr
5O/6LZDLaIcmaoimBSyToKUHKEjZI2aOgYqyArT0WcodfPo5UhLWG9mx/MPY
QzM9Zb/+u+lgKUVt7z7tudHfRoj3YzZhVlCV00ZKEZAz8+ZZnHocNdiD5CTW
Q+0F912S8FvwCMEoPuRvLz8fkGXkxWblBWYu3Dtu7PDzwMAMQg/QUSsTepZH
+seeAKKxSAHRBK/g/SUw8yAkqvAYPPN51nMKl+tDntGjLiKM88bqCHHzRRx6
5bo0mg9bCSOA9aJzIxFWjukzfavl5YF6rMHspp1rmAJFE8Bgo3pF7drTpRug
JjSsGhtDewM+ufJpaqWsKxxQFkrCRplJbZr5K6W8qKgvb7IZyOOGX4qtpoCh
I2cGmRij0cfE9EFCPU7622S5tqJB32MUcWGXYtWedHAJ8yxUo07ah+VGQgEZ
f147INsf7QpURokZrgOIIDW8yI/dHy5sz69yJGC2XZMDFN6kgCki88lpTaXc
ww3yokv2s2utXEHMMqsbPHE+FSHaNODfsHg4DeraHwGDaufkaB4fGXuNGsbc
nuMuXme+PVFfDy9qcW7tfHqSiGU71Yolsk7Y0Ns/dpmxJ/umaq0X0tlVTPAd
BxL8J00dl7rQve24b/OmsKkXLntT3kVwtGVyBwMNmlKTcNcwi0vN9cETOvIm
zSMSjU2hprRByj9F1kRgm4+1U379PTrEWFtC2AbPcCMU0us4K5MhCzDRQWUy
eZdPcxMrpMM6jGJGvbIE0PM34mhWi2UbP7Khv59xFQW1KgOkj+XVBFYIWj37
W5cARF3OL9Sjv8nLNp7Sh8+iTyHcDGWWeUkXDUwaPNUpc6/TGmVkU8W3kMOA
6n9B76k5anaq0pB+jDBlxYr58+6ou9lE3tinHKlN8LVpm657QngkWrkHzewM
X6vvNWqzAmhVd2cRplaM6G0mMI01Ka7y87GzwYD92G1rEBJW70oUJW7AwaJq
Tlf+RuM+v7sJw11DyyU8G7owpyRDWfA3dYIuF5NFJjXIVQR1wnA7zixJp7SC
xnapuqaePzf3KyKA5sYCWz/x92uEY7ya25PEWQgnwmjEMIOji1j2fOthWQPt
FlRT4PO4Dpo6/WOn78saH6+BA8zmfAeofRA5LAQbprNNcqg4u+gpCpmzr1Lq
cj7Qq9s7dP+H5CK6poVEh8q7xRmepLL81sVZdP/qIku52H/HnlZCwQ7bP4pK
compev+FTr4wc5QzISr1NbNCyOeAKwuYuNE0iGNsWsWeZJ7OU4L9A04JlUds
Z7gKcRXy7Wqz/c4sDFdXTcW5Bi6rEVK/AWAPQtDtQ/mOH3+U3Tg9vmBTJ631
w6FgjTUjvaV/Z4+82kkWCjqw+9Ld1ER2bKyNB9jCyWCXzdk+e0QjkcxVVrLa
Y6ntAVrxqguobuzMWV9hzoPjQEauVfYZLw3N0I2bsEmzddIkErYYEIcEROUM
8PxmpSIFHLZLIJb0SwocaB6foEk4zpQg1xFPFP+PuO5gDfvWDdJg74iAI2Xo
RGp2I7Sgie8l3c/+7azKusKN6XKHeq2Gec4k09JspOsMK5e2ZHQCuH9qJSpg
4EwcSUeils60aDtJJSWXLxnTvfsnbmhV+tlt+WJb8fNpOisap8tyoIKctuBo
tmXGYR8CfSUSvnkAWLpDKIit4RSHmynzv55be7lSFScHLjjqjuZdd3EAzoso
dNBmPWzmyvkxA0C7bYh1nCmCXj8AYVWrq1MdqKH1UivrCSXs1q9OVivc9fKg
y7kFcROfIYKrkXfv5w6fOQ8KFA+azmh8iHmG8FK9+4Ui6Vf59cbfla86QSGP
sN9FGqnX8MNO+n7hnvy4jsGQTYmvBS33gYwnEyGwFOQqMMSioHEM+1mZUiFs
jNdNTGQEi9qlYi6LDZ5QEv1+37PXf8HQYh7I9lHfqDrnYvDrYPP1KZjQebzU
CoUCRr+0LTSR1Eli8GzMAu759B9EXXO5vehZkUaesfsfHXkgqXeOv7ttOY00
+L016kZiyBDU13CMoviMyS2BHnZeK+eSzL51n8xbqcw+Q4J+QRgj58S8mev2
AgYVLwrK+OpTLr2VmW6CWe64xwsxdzpUWJKOVN5m4S8eHFfw2y3duIJT6SIb
X6WGkYkz+UHCQzujTV9NpvzRdSN4uopRAEzxu2Kppsu/0ZQuTtc8Y84e38HI
LsHauMNn7eHR35TeyheZMfwdalPQhFaFbBM1q/wnTHPlTtw5ndj5EwpMm+35
35MJphpf66Eu038JGr+28kgm8J9YREvlH/1OMQzdhNiDl2uKViCIbAEq1olu
Q2Vz0QLwDBFzCRSp+yAZOQJDChUn6aw95qzLQSpiXpDb7NPLOwcmFHsI84pA
C5lh3ZYBTlzoHNDLKOniBfSz5KoVGhXxbAhu7OLp6H3bZ+1p5cpAiKSDHp2y
PHro5EODkfC99927HUEt3iy/0LBWlmyG3iPH7Gem58WuKrZhYoY+PokJ1Y0H
66pTYVP5ZD0Po3NoSmrWlDSQhygrx64/1rI+Pxew3IAphLTHjQq+Q3Gag+N0
rGAzLiQ6zoJLBoFH2Bi5hSPNKY8UyOg7xwbbj9WuqGC0TSRgl9WgBDsJhdwp
7cMYH5X0GwAAbXLU87QmYqKyxswfmBeHUteJK63omRSH9gMwhHuaYEByKBBT
DC3JroRFNI8Sa18mp11ybqgQ81fue0OJjw12CXGw6Cfr0QEONzHQik8jekxj
vHxPrlZjPRrdfW6ljPGmwueyoQEIGd7v2ptuvpw2DjJA/1ZsOyfZ+bwh160V
asC9kufjVGlpXRJOfm2ss6B3i3AY5b00gnjLicjUKwsa9r5sxUp3mMQFMvpq
/se9ebPsTXWrsUhAo737/SvtdrMkUUS4mIRIhfYGee9AKBaIi2YdSUjdOE1o
CvdHEqR2KeklG/mnLC4pJr5wMHZz5R7Vnf23OyKEkJ+DpcImx5BjiCUmBddK
uKFX1vg9Dhu0kRc+WYT3jpMBcsbClzweZR5fRgUw1xrLIVfCDbHvphqTEU1c
qg+HcP1dg+470K1d3myUCNJZ4+33DXvnt2MWrxzOdZYSROI5gov3gYUdlRcN
l6RIFt61GpdTg6tFqgc6V0gu8+9IGQQvei/N+x9NgSE66wpBpO5kXBQzQOFI
fLNoR5NV1okbT60G/llnQYAVLF1emN8N2BKv4CCHUcjgwV0wPM9n5+ZlLKVU
gW8VhC9KMcSOnlYnyXgDZeUdbVKlaxfNVgahXj2FZn9KV2ViFWsjfZGO111r
wnEiJmAyBHqSSVj4Z5UqSXzTi1b6diEKGi0cw6ssy4ntmMdZ23XkjJsSU9W8
w8ct/wnd4kxpa86UseWj0u+0fqyBpqCPIQp+j7oOTI8UVsQoJSPsQ0fZWl3S
nDVmQR+oWZf2m+cmwcjAHkdHdt/q5Ee+hNn0iten2ZOLMLC6kfWXoXlLusMm
rwlDjllYvRb9/EMtQxPd/h7VCg1NkmUM4qUklbBX/9FSClSyjrNDJzYqA96a
KdG4tgBy60rggVDm3IOqwvNyp3WAaiDiAUmZOcuPEL0Vd5JSB01MGT4IVl75
X9a++9TQs2cy01+sCZdrEQILQnmvNKFhCzGRSUtFBnDLv7zfLe4UVYmalXsN
fdVaqYE2LTkv5Kx93mDvLJyZfOz6Bc+XrzNP+G+RIy3tbzkvRFKPYUWDiXRB
4AR5NJbGWwXOAZtadRnxUJnpFRICXHIe8D4LZlLT7/+/Lue0XlslBKoMzmqJ
dMxcFhlepwRqV9ySDaZyNCd2fOavppbfD0m9t+LLZRwUoA9IhUYNkqSYHh9W
oLpMjnyMJGHP7HcYDOpVoRlTyf1UL27VZrmZ3M+n5UmnHj+Vd7MQTVWBpXuZ
kZlHKAg+FbMzX6jPkoTAFfDAICtm3Qo/S6sA2nzfEpbMbpY86nRG/vNsrtXo
/8s5nXEZm31twwMlGRY9it79s2oeU9O62SASAsQwi7qCFNzOUpzevDOKgSBg
Q45QCmvBEwA8qx3dDFxSwWZjYywKuzCCXKLIc0vICsbSqdMd5DWe258QNlTD
VDpEZM2RhuUqR0ClsMWatlkNKt8uXZFfK90lb2pa1M+frEjrfBxbMTioav2x
DwzeGE5cMufLz8nQ4JgMb7Ff8G5jk46hPg/ebChdKnluw1HbrA1IEKjYVUsa
7W64zvMt8+bDOGnc2BHvxxJE9lrkGvsrion9Pn3JlK0/CeLW1n3PgZc8FNMb
qb7NeVgdptEb1ILB8k1U5ilwme8727wGlnPOcMujua9RCugs4WsBqkjwsO7b
r56C7k3GthfYFaQJCYc//JNoqxEwX1VQ8t3XdnnPIn3nctAG5hZNYZVDm8Yo
g7MVoir4cNz92I/GYDvgxaDDjI81LS7hQgRhCD20BBs+sstbxhCXWU8eisjg
PhdICEr/+VteyS/zqz0NHNYScGwIH795YKQNuHTs7fS7oSSByqaqnzlyOxA4
HJK3ouT9osdkBY5J9B55RC1EPWEJ5yXgeUklEJCZHrOjoVdx3ABz8P/kobdB
ucs8ActoLMH5bThyQq1WCVavtIKzTNn4Ot3eGIITjRpO++j+xh0KLYe8iy/o
FWmVFIM9MnkeF7sYT7MFJf//olxDBhYXtso75gzQgQz6d4qv5S/hmDACKZQ4
Q3pIG44/7Lctn4Q/jCZQDy2Ze9Uu7rX2wcrO+kmnSCZF6P55vjsiU3of1def
/2qidwAOciQ7B+exNe7Gr/Wfg9jkUBk03alg6HAPZCUZzfw1Mkd9sWhYwNFA
JmVm5PT0VAlNEaKPWSCFiAleCmThookOXpkcL8CPq2ZtmCoqULhQwTetznpI
KEjfVyutv7OG1/nIeWJ/evOeqGZ2JasxN0+YykMJERoJwLtBzgoLdB6O+AE0
cR9GgbFymGpL+7TRecDRNvu6XX2tQuruLOxlbYk9MHx24nTKw6SAKf4adslx
fPuMV2Qy1Bp2VbME+kbxd5uVssThwm/RAMOpS6ZFc2XIBGY8fxQR7YmIGzsE
5rh6CH7wCRQHIge6Srbn3yqo7AV/7eoqmgznU7vqpCgPbMNE6+UcHf1X/mz2
MDwyB9et2zCCd28OKaFAhrXNnM8UApJK/f4X3+WZZcY7nlwcmSJHmtSARqU5
8+1+rZN6mo5Qr+nBjD+WPMppz065zq/sazx9DOpkhxA7fq8pPOFHU9IZ3zik
l1fcxzSfORid8ViK7i76thiHtmSQfyR8mi9bQefBMLJ4tHZ2WNcDuAcBznF0
BQMO3wj76UiHFJmt8MWq9qJjTkxWdKf2yU1kqXyuFXQJPGWlJC76vs1FYE7m
U8vzhHhpiFxbtSRxUVNSfkI0ag8+oB82mLsXTyk7SgOrr+lPDKur8VVtGeY1
jtnaXcX6W9u9GXHXg23Mh4Md609/E4aeafSYR3DFj8L6apOR6O9NkbwR3jLN
4JiVBmm34GQVN+qVpDMROxx5xkCHRt+WXJwbSrO73HkVbBpRnCYU6uCgHSXE
ProgME7vPbA+XPoZv5AdFcwp3Fo0SuCl4gRxu/lZbM6bHW+KsVawfjfbYoGw
hqfz8cvXZKt4vgLt8SOx4fB7JzoBbZV0gbKvrmmjLlpE1q/fryy+NKN8166d
qKjOSonO3iT3uup0rPPcKpkeXHBocEzH0b6W6NdDLC5Q1mMcl2c7ZCb7y0+d
6fkUz6VoFaMJQ4MTYmAEUJbDr94mte0iYk9Cn/oexC3NSX0trjWW71YK008Y
OH7KUhsDrZs9JXPK5sU5+pGNg6ptoD+Zy2wgLoX2x2ignWu2jwiY6wATNGdx
dgGTOu8jJQ3FBwaMZrXCHSGmZ/WRjLPoxf8kVPQVg9heUm3LDBmF971SyinN
VkWDRfnR5CasP5c2vOvRBb0qpnga/QHOrcHmbyTM72GBH8/F0a+rVHr/ecZ9
liZv5z9ZbgR2u1FEyg1yxeCoBCVBrCfuHEsEUstjj86tqQUBOEqr9tsIOaz/
Sk+UebmYcciNgtHjvkGCxSK1hEwXGlHSu2sc57DLve6Wdo0RoZBwewZSaq6k
9MSmE9ZoyKgpy9wLy/0/l7X6hNW1YUNyleQ316bnDgnzvCUUxyigegdguCfe
e5Z3hJD3kej5OpoynOI31h9m8GcK1hYpCckk2CIVsFUhtDik5S9c0/6AU1dc
Idc1GmM4ZcPsIxN9hp9uFIPgx9PkWzaWH3HCgVVxKU84eCSs2TB0JLus9w8H
1EXUJ44zUxGynhQo7mMNIPbEbra6nFWdgtusP+YBKDECBUynw6ygt9w2Zrln
h1MzSrGOsTSeu1mIq8mPrm+oIdUGI2q77/DE0bjYedmv7DRIoCoVW88BueeC
svvjcKGjwmJGStyQGIM79m8DSjXHDgxMgstSUlMJMsiAR1M35EMXWz5pwOn3
VNh6IWAuW7OwEqPFtzxoIev8IKya6mokRIrUYQRii6LFw8f3cB1VIdpDT5o4
5QDyvcbgSRdEvZgTTHFT+EHtTNAxgO8PUNxHFuJt4tqClNS0Vz7kdx/1lzqZ
jPrg2mJ6bceclYaaVR6WTLmTEIdP1cahwc0L9RMJ+oNpkg8h+piKguY4hkHS
YL54PSNb1zRYCTYS1rV5td3jikZITgObXBn6TH301FJ8ogYGflFUn2rwYEOK
sFlH7O5h3RW/mGJT+za3SifwYJzmnYpQcnlJNf0KUbZFjIpuwdGiED3L/rp0
eXPtCQR5OFc8p/2mJ/0Uzl1Va9cnNV+hjbESZjGnz/97mes6QtzPz2r9sIj1
2VqB8NrdNaXbtY04DHtvqGAWnG/ArEpdNC/j9HFqP7mGZZj1RXAcPbXtZpzx
ilXUDcerDlBrKxphXCHZHBLoKaGV4eFNtufAijidnujslf0JcGlAwYSz8BLw
mtl5SGtG5eHOIZnSfwemsUnw4Bfp1k35vf8lbTfDNet0owDdLuMYWpx7TIyN
ANyFC9MxJOTy2UIzjQUeetnkfBspYVqY8XasBt7McX8ujtPVSFGM/WmENgQI
I2gH+PmujXEGKdfKfIwVCpgzjHG05VkmCUuEGNZY6gJv4Z4mSaCGSggdauIx
RN21Gg38FRI4Qe5lJw2PMeNYTGOpR/SCpCkR4Bw1lyiVFrE+40Qfs/OW7sC6
Qv3KvzhroQlkqGVDHzthMXUHTQE4PTxBO4Cx4HUpFbQCKO+yDOLGuZ1cyLvb
gmELFPbaJAV8ZRcBEJApcPp6JmQjvSozmHz6Y+EFQj3AEMEoNTv0qIodavUV
T13VYcE8aX/yjfvWat+CahUl6+x8HjDTgZXGqtIE+u9/Kk8UA4Z8kXs7Oeq6
h27rQKZD4MTrEKtLaOnLN2jZq9pNAXeP8+zba1maowEcT4S1Z7eaW9wjVsMe
8uUXHbLwXpxyS1Hk858giyzpvMhpHfjqWI0tRxM3iBJLXYn9trgkyddoFMEH
aDDwSqbDszLE82xa9EkG/PftP5dCoprecwbi3n3ssHWliiQfGZ0gOf2E+/XN
BiPKd6hoyBsWwG/JiYi1WVEnLvTx5AWJ7oto/JYvymGlsk1AWqaENdzd/EXw
+lbK9N4M6iNRUokEQkNyv0QCodxhBOmKph+KMzcNU2+D6ACwDAaYwwBVGzCI
6QnVDr/qPpVgDmW89ZwKx0pE/EchRaFzPxbN3xmDPIwtQBX7Iv/bek3AcLFJ
XS0Q0nHSn6p2CN+KUgRKmI786mAReCr+IBlqEzTmUUftm/iK0lLal6np6ejs
PAIySwlRJSxeNKz1ZKQT7DLTBytd5w4LX12iQ0nxVcpKvDLNwFQu7wYZMA2p
yHy603PiKVheqmWQY2FjBR/Eo3WYXByTFo0F4UmvGn5yh9T0hECd27alqxDS
v0KrK59viQXF0ZHkjsZJRSldQ2AhjTpCybk1CH/9CkI0M5jhr/ZuL8KXffbU
qJCBDvfcZ8agrUqePzYn6Jql6iy5F/Ky2SK+AvnMVdkyW+4QiIwoFJom1GA7
STTdQPj4D+eY6uJsdzxKN6ZAqonxhOVt/K4RBpEcM8DrS5cXKnaEJUqIqH6D
wqAXcWhscEgvhGhqW0XOtnwHqUKxpWEB/Kp9dVA3YQi8ZUuqUtAhg26zp3Hm
0PMCgzXA+rofp1NwPeS/b14z18ZUc8gethZb6eUoUhhUrrEWiaVmZdzJSUNn
wfJjllKDJAlPVP6z2zXuog5EoMEhVZhbXloyQdg2kS81bpYa+N0RQ2hdLIK1
2keBwYnf7bFPUIOEuxlWHmJk92zd/0ZA350zCBHWDrfOlkd+J+uSJMZwNT/m
Q56I64WShOoy3OGHk3lPTnySg3nZ3DjQgybtacDQRxAg/HCo9NopLvReELVQ
FuAqSBEJx8AX/DQI1PJPT2evndEVHOQq6FHfyXTKRtfxn8VIdqbdU2DmVqV3
P9f7OX14MoSGqr/v0qoPiSa6krJAm7ppPYMd2Isk7IGr+YjxKPX7yB3msUxw
YmWQmi+FvrNpVlS33Zu/04aaP11lWLSHxY8f8ZsFMT1hMQpdKMQPtL7h5zhC
5yYiQYWHBl9DJCRL+kjRXFV/XnVUaQxrPa8r1al/e+rkJudQn75tMNAa41wD
OAPCncQVuoNcMXONiJ1X6UKerxiysrI+sgETr0e3bvF1v/6yE55Vx5kHeNkB
u5hgpmt5Xo6/aI8rsEYAi7xOk/AVZX2fQruWl9Br5yEgBkinnQotfNHqEjyd
JItvMqf39T+vO33LxIV2cdKR+eCm6RkLxLCNFfZjY7hscHLCNgOa6Hysh+iz
qf2jZz2aFVvqRvYsLsfluTzWl87G+QPEUMezgRyxY8+1ak9vN4x1TldJktOv
UGK9+yq9YngJ8S/CbfJ8YKe05p24R/Nfw6aAdzd+Tq7fGbKSrZU9E/8QrgpK
fLBONByonYCkxnBff2ufiS0dU/oGRXxCO3gPeysTVK/RFOpkrTWI1QXLSXli
R7JsVTGCEXEk36tbFRqoVB9MIq7Ug2v4piQAHRYPlfEqOLVT9q5EHNTqEt4b
S5PtNGBjwdvaW8hkA0SqL8/p5uTuDb3BtVsL6zYKRybqEn8WfvMFnFXLpffS
RTSjUd2JphoDy3/+bKGYVTNNF6WENtQueiTDU4/uQdy3FkfhqkfgNdOnP9hw
949FsaCYxrRbFgsQd1kHaQITqJ5jBEGUI/PsVn+Xoy0zFgML8NE8y5dOIcIT
jUDcm0i36DlslcPj28d7hg2D2UUfNU3yn0JCDlboLXGDsdnwwW5XNEKRi6Ho
ZVrRuegZo+etLdmrVez3aqdsXUeFa0OkxdlxZptCx4ev+m7DOSp6DLoOJsAk
aaKUKQ4QADoklBH3x14Kf4KxMTF2ofVv469iEbHBb2aP6iFLp7Bv3tfXZ5Mm
EjuxCNmGRGL0TSXMjbjGWChBBBvewqSmJdk1s1Uwq/UBbAKJldjvy73UItk/
BZP0X1MFJXvC7pyw0SnoIufT0TrL4j19fBASuQ7RNgwXyIsdGqVMB6PR+Emp
PmF6Ami4CT1pt4HzUMWXBvmRIfjX7/qhDLhb4ZcABDhlgta0zwp5cmljrRds
mPCD2aJX7kUEtvT4cGsRQGWMe6EfINS35OeHrJvj+wt6CWZdcam33fiHCEl0
nbwPG5nGLs6ljilD87oLJjxc5Dh0eWbC1TvaEjgZwLQ8ZR0BoKxiV/zCYrvL
vRbF+/ylGgmBnrSjCMWklyIeVCgv26NlNeTjc1C0i1yThq37dm3RgEw2Dac2
OwJX6/TZwnH4nsllwRnoGSuL4haZmEau0ZkjePdV1YJY9DPbpo0Zl3NH52jj
BenZAtxJu8cdM7c9M8GSv/V9nLRRZcRi+DEFGncb7ok4CZVWVS9Pkx/Na0vA
ZDqLO8lRFBr20pQizSmfkL/4TWxHZPCuH4DSWO9y4uytu5oOZcyUlIHvfAZg
ry6moRySPhzmMKZRbukIh23IrUtUJjNWYDar/ZQCwLBegFmssqZZHlHOJwRq
on4TDAj0DGsVT93X9aCDdH0PrqgCcDFmonND+ZvltUqXDKJU+FyGdcrDtvmk
ez3Wfzc99AQN1VsrJS66wiyRvhHBOI9bbQb7bNtFc3P4EIGBGD+/VxfIBQq1
BsGQO0GDsTefQNw+5z1TbJRNCw7G66pnYejFqqxDwAIvYSaIWJRrii3oHYb7
J5sYm1AYnqcI5MFTsAAsQ9H5Si9Zq8AAiuYPIjNiHK20NqQ3/VMQdvd/WvRe
V8h+7nEv4DstbAvzF5Qtz/zhzhIx4zfAp7lOTUL0vshlcjzgMWd3wHtqHL2p
HQJyRduBIfs0YTi5IpvfR3mx/zSRXN4EsE0w+Rr5P8iqOIRuFLfltA7iIR+f
bmFtGIwByBHpfVv297PW9u2JusI4Fsj8EagbvplZfolDjQ01V/y7WL8ngmoR
HsEG+BIl6hja06X+afDpewdppmVZsg5Pi5ssxCU1EoSE/dkTCW07quL9pz6h
0utDHiGCX5Ls5i2VORaYcFdVzc5wFqdhVoVMIt2CM3JY1JB+S5H6uGci+GKg
hzSeAAHJ0+3hi78h0M7zuvY5hY9Y0tEGPLM0hLTxtg6FBJB7W5Dd3kfNdi5A
KZqAKIv2qrELV1VWtvkXV/8kdAvNcjQN1e6y0O7BBBcBDAASTmvrITOfYzl/
Jo3dqLYttGhFrz/X15oO8o5WUYwMePszrZliqqfeSFdUpHWTiMSvcpIzO1H9
xfIXqOsYzo9IJLcHy+1Qaqwh9Ksw8nmx1b/Z3fAagC1hkhygWa4QBI/txA72
oVHLpIpGphLCkWLH+ErueqshK/B1r2RRX4fIlPtL6Bb+iCnRVN48d4E2I8S7
qkXW4F6NwV5OB4psCmMlpyuSW30W3rpvs1YpOn04GPPtf/1hS3zgj8GD8tu0
8ikUEWj2SNum56EWjPjIiwZ0S42vcS7tO+QOZ6jXt88WvZCXt6j0I9tTFmvb
8fUuFXfnYgxCljeJc4s4+njCpwPlqvIRq90l6AsLVwtwBAaw1S7jnMA17sRc
LcEhON+YSLwbN9WPk7S1hGFbHhVLRQnrqK/sOotJDkhqz77c2t2T+s1VbgWg
UVxxGqUIbbvKban4lZ2czLBKfTjmrghmFiH+7p6+yYI+9NgNM/qX/LpVZ8Bb
72NyuS+WyykQ1mYUi5JG/oOsApapPRIW2fhTgDVAF3GLNfij0a4+IMKtHe5d
fhBRVAKQjUPhCRH8YTurNW1it+PFFVAuo7A8H8rcgjHFW5iTzjhUEVGZg+uE
Fet4VlTn6RDom6dmbFgt8Ap4edzZrZO8wHcSy9K4o+DcklBnLMz/YVlwWvTD
qMLD8sX11hxTQcczNz7o3LfUu2mRUj67EGVrIvWzmFF3u0bLTgtFUusklBpe
m+kiR1IDMnK1M4XNFoFSqyWdCHVQeLS7iurlo8VX8rNeo43pzVvgf3osUvnr
5pQXx6T+TXpYR2SWAv0SlJtW9ErBYU1xrzRsDBh2laSt1zc5Lc+m+hn8mF+i
dcRSggb1lebz9w74W4+a9qnZwPj+eC77x11SMEXsB02Ct4ayVIIB6Yjl9Fqq
xz4rP3t7ffwAZlTcBnqEcjm5KcrK+jdNETPBp9t88a7+S615tPCBZ2j19Y04
ANkXYYbhqDDv6Cp5TtnnBWzZnC8KbW+7EknwTb1SK8PS+Gj5aVAONvUKuwxe
997T3N93/FH0tKxXTW9d18htSnMK39QbEZhSgDcn02PR8qZGltyjnveGMvoO
qp/xB0aF0nXb72sozN5KKRblNYZoPFobnK6efV0pPm5gGV4v1/hi2Vi1us/w
nVxB0Us55zQ+uJgJZGKQrifpZfPPSZgHQs0xpJQLjnOYJg0Zu1ncKTRPVhT/
jKVegFKo8nImqShcIwqW7xomfFWnO65Avqeqb9l7b5ErKsdFMnz0jBtookAz
UGbMQACaYhAlzrZqhK8xNGeczzc7kmJhMR8Ol4R5D0KIiSRlPe10z6C0zRb7
ejEZy4CFDe/MHnpCaNo/A7ni/8L8M76Jl8/UQTrytETtqatqQv6MRiYfa2Wd
Fz/OHxjl6ujVEyO+gD0uPk0lpTbYh23dmlfHZVy89785HAsPj4ZsN+eR7O4d
s37i17QGjjdrWhz3eFQGcOB5arM9dyLuNaQZ0jAi/NUPdu0vG+f5O5FIJXSr
9aoPjO2+VDrpJO1ls94smaiyhcXI7ebUtaCnRMZAvNV5ZvUtyB4bqLo+kM95
xS/OggG0Blhymko0v9rEZc6bS0gkr2vkimocXMv8nJwCnjhjHUwOFFdgqCA0
72nGudbJmDpIipcM1i6S1V8O7RhzZXNzx+ekUFMIwYXF8QaMUilU54Ps7tRQ
npBoN0e/ajn9baR0woFylx5Q+31ohq9DA9Fxu3FmiDfESCS2dZEub8KBv68c
VD3AkYS+jS5PUrfU9+a9dRGOkm3cvzD1OItLLA6yld9ACWsQnW2Jx9a5jO3n
2A04XgmKbOrX40s0Eufvf5taQlOxuEZZ2ck7FeuOGizCiuJcKW/5ARH4Jbaw
7zkBP30VviEWj4U8EvuDUN5i62YzdoRgZbt42xNh68tKuX5ek+PLT5iOoHvm
8J472ECj08yTxatB2PsZHgQZggLu9C6eJC8BtmY+5GLWG6JFb0K4w26ZZiBg
lNn/rjE69VBvPPhBJ3aZkJrcW4iWgVVVQ5g/gNLwYW8pjXq8JiD4kvTQgQcR
1k0v64uDYfL8vdBxCsNLxMFJP44u7bY4dL4hcP5pp90QUgAhD1uQbJCHPQPd
yvNeW47eMmMd6UNF+lGhA+aMd605dhz56yddR7IheoJCiCGZeAuIgsTtj+Su
9P6oLd56JMpoV5736QUuquzzmhc4qazk/mrHEXptImMXlcYPSiMtxcGOmE44
hHvTWymkxeaVk54YNjAgfF2a1DDkqwXtfTCLP+ldoONwM3s6M3Mocsgyqer3
aafXAto1KP/ECGFUN0ivjAf00OE3MtUMwhxnoFW6DtFn5sg2fJGb4RZyVgFM
dVZh14paeGUM/FQZDdkjpBr2WIk/8EdtFvHLM9fSquD8UvDJyGurM1DOuf9p
mGOdMp/DpqNn8subOHInrTSuJOxcYYw4aP+DqXzYrV3vMwwKiUzAcXzKcqra
IKqzvCfomV4gurnb3TV8YqyxTQ09P/it4Ozqz4nh+xqJHfHgdR66poBGZMyV
z/RvDgJOlejWPJZvrnhjd2VGzeGjLYtD4E/QUgLzFBNFKqe0eg9LgYuV7dHM
fjs33CeGMg03WpzXsBGz3aw9xzb1lIBnIIqyWzLz3siRKvUO3gBYJ2ebDYBB
u1j2JKGS1DogfGQ8PqXHlUlO0P7DkZNLUSdGRMPfsUTBxsCTpUl/F9EhzNr5
/1hR/rxxIQNW2iEs3gpGoHWvYm0mPqLggwVpl22HDSD6cvAwCY4QWVzCjlDg
tluvp6rXsLtjF+0cUVHt9eyl/c8sCFvFYiQPFp6SgISS7UQDI9tTRnroP8W1
0+8P8Cf1dmkggDDKTpzz+EZf6YJEEo6tJwyCd3Wt2f9Z8pOEJTW3JE3m9uwg
dHMT+IdH+bYrWAddMrSBq+GENmfOCXqptPUSFfPDbRBC2Qtq2QBOOx8OuYdN
udfYlxYtww0WEqCm1Dxy05117VtuWi7GTi0tO+ZFSSumneYr0uHBQ1dOArJX
bDrt9Uakh69efAkTbXQpw2VkZBO+4XIlqTKaeM6qevhr0gUAt8UQARhwnl4m
5CYkGVO9pGFhIiI2DWazLZz1ZiVCOwGENUHzgxEoVwI/wVUY4n910vsYoHhg
MdB6KMHxtwY+DmFrlkfvmFr6kfbzi2+4V8NGVomh/KwYugJDA+yKfg1lYabn
cDimux6vq6wZJJ//XzkO40BBsKtkTYbeYQS3RctcQXYIImPmpCZ8bCeK+b6Z
661e2Hbs81DLQv6XQSlHnAEY6AVu5Zq0/fS+iL3qBrEHJBg4g6V2HXy7y7Ck
ZOAKxvxia9N0y6/9XgTJBvH8eeBJPOMl4nwOTPgfyCX6kS5zmQJW9nnpVNal
3F1KKJXfJ4DGnDHoa9ZyuHQrYuhZuWFGpIpT1GC+SLyzBIFIMiiV2UNlHoQG
UQnWha1XPTp7r1a4ivzHRkr18IULG6d4mlHoyiBJVBX5zjMMy+kR17fuV9P7
/W3KHEfbN0o4KmIB1xWWTXZ3CDplr0W6HwcE97Xy8JbNjHCTtQmDpXHgFmCK
SFgePx2DzDJLEYvczoFfGkumQuNYQBb089+Vm+4cIRIEwlSif1c8ORXfwxvL
2sxYPcYDi0h6eXtTireNbwBtiawOWYlVnYVuTewFVKDu/Fne4zzNIIEOKsd7
/0LfUNleyyg76ZPybmdEz12cgKeX6nldF4sz+Y4nzXLojnJeBDLlyHaFQEod
Zo7c/RBhzMqcwclH/nKa6n2/uoAUK1SKI8l+eyPinPquyUxjt0EnoSojNIz5
ohnnzgCzZ81civRYGTWiwdIahhpNWY+eD2jmu5AhnVEFEW+PHfGV+W7w0AMs
MsjuEL6O8f4tHOYhWzUS0ocVjHSDQXU3s9+WVAgJV4PPtQ2sYY78aJwroGly
Xi89cPWP3qpOe2lE3Fdd91ai3YhRyI6lIW5+r/KBJK4kSQPwbHbLztRdmIQm
JKocLm1VvTzv+PVUeqsXEzmMocCv3swbYdV3xJVNZGhDBrzsIg612uE2zhVx
BmOwDrDiZ/4wyCitEJIcLCmoI1GCQXTTOf8k2jgMZVbjs/tQS19r9TGj1v1p
fGYiHLVNRVRhEbNWw4NvQ1ECwWPmrjFUdHiFRsg6YGpneoAFB8YEx/EsYnHh
9GGPQbANlN2nyuHCTOxCsfWfFTT7FcCjDVGzvFur3kBMPQZ8/vdUfWYJmFKM
3VKqcNNUbsXKIBYJ79Bar597cyHnIZfotcp8rpsEQeWxjP61UjTubcjt2oiL
wN5edl+0nKO6Tn1xmOcjw09QJ7dTO2mhxjfhy0cgnqy5BdGrdlcmtnGRtkYS
gOHHPHPsmdM/Dk+R+Td1YvEpeSp9Oi7i97MiPwGBEATy716BUPUkrShpEW/m
anxPZQTcw4ka05AHWKMx8xf1AERc+YvQD6MGmzRpy6mw9PVmOtwDfDIf5Dmq
r722VakoISC8TQK1hy4IKuTrf7cNseO4ACTO2M6B5S2HDqCvZwAzRjklB1pj
LSYAXtT4SjgbDjCdgV83DlQdUSFPkD49LkeSfHaztLyD+WtOQP4mRXh3xfNM
17kURrvuTOAc0NtDwPFvbVf2jRRJS6K6vGLfpsvz8OxD0TfS2ASGxsBefo0a
X/xUbf2yxLAEycChRQy+Afs262b048gAVCIOFJVg2ZHdzTCKYPzdI8StPUDk
VEMljasi4Do7rWvIV+zE9BnZlIPCY+Tqa9SNpK80n+xpOuMcQWMtacl/+5HO
mii738LKupYr939Pte5IgMOn0SzQ6Vrz/CcO+8vHjAOwzIB6cjw5CgGiqG2u
nFPX6KhvyOZlF1u5wTnNE/oizfwAjOZk3CVk2eKyvjYlE81o07mmgHLgyffe
Odg/WtxyLXUUGkphVOSrS89CiHM1uP3X+I/UAt5dH9KuPEoV+zl67HDuWq9z
i93ewhOIiIjTwS1w2pzpfTcHYUbmpKqYITDyvsMpEsNCE5CaORPt3Ulnpjr/
y/T7y32rzu+lnJ3n4LefCjjjsirkWRXGHEm40WsCgEB+GrFx3NTlC+uiVNpo
K9aMULfd+yfxEGBsz5hIHO8SITPaY5Q9QxQP1F1trXCuI4l9OOb5V/bsC/iV
CJCp/hoY2lOmiNUiflMw36H/YkmQxzKkJj/tVBL36K7T6FBdFh8MkAlSheKy
7N8+e7dbI1m030mc0gov2PrCu7I+ZHID78HuIu7y72PA/eMTsWYKoNFu6mCP
3cUg8it70s5cbPa3lDBvp/e+h5a9E5bKyhhHTJRGnuRZEBEn1mn++VVmn8pg
+L9ytm/jVNUY+cH9lUN4qqvhLNFn9pZc5tw4jfKzYLOjYkt5FuScH/YQQp55
RJuIVOyvVdUkEIWi4ugpD300rQyIzAF+YV2WWol1Hpp7q/lp+GNHE0qUu8sP
4m9thk7uIzaqTA1vNNYlJdBn9SwRDOF/d2RHqY+EAirYl+WrkGUUbt2mZZsP
vb9RbABOXBBvyvvtFtaPaM9pCylRsnAZcjFCupFuE4MbCwnnZpDNc7RdF+Xi
g2tQ98pErxxltPdcGosW7NRYdcVOiB+g5tFlaxWKAvn3EqfP9Wlaz/WIH3tO
bWNodslyxMV16mAQVnUqlZVbeLjyBptgzS7NGbeh6lqJgHmyrG0BgEQOhgxG
yNtfPVJsWlxw/Mv/gjrAF/o760aB8ARVJucp3+INRHf1+XzwMZuFs+6QQofz
56Gy1WZ1hzLn6bROYtUhiKefpplqZFUGIe0W0+Ep4CfZ2xOTYzZ3uoFuLvq5
wq/Dei5QD3EyGWwmkkRrbmsQbjsoOJZVhp77UQRymuoFqhI2B9TZwWcz6v1B
nv8z253YgDlfCq0t8q47TCaNs1lqwlikIbcrDX1SRAD/tW0UR9ElFuEnYeY3
uyMP98ip737qi+WJl+IS2Y72y6N+6Wi0kwbRRdHC5N9nWwRryVVlbfXkeLNL
8hEgu5b5Rd+W36g59sbH6VZbYC6iffrgTnXqmaKikebbGU1l+ieCJ9mArtGZ
NUO8SsCh9gqpoueZDfI61xyCe9dXscg4IDe+FaL2VQlz3eSk4Z08EtA2Y4tJ
FUbB70H+UwdeqNDXlRC/u/70J+B0QwD6Ljp50Q7bOuIH5r3xtz7pjxW1OL5K
Z8yGaefs0mvaK9Af/7G2KbN+wQSnzTLTNCkyWdQz0GfTIVfdIhuIhqhn65be
gFoc+n2KhNKBmaLLkkhP+4w3AwinmM2MNhUM3atV9qBq+GOBNYJU4Q/ojCZb
HQdcoysuuBZMWokYRWJZvAvwP8WPpB3t91RSDj7Cfy/dsDHyyzJt+aO/Hcz0
ZP0ANeGSFwT/0zli+XstM4Yj43PvPtCSkfIqbv8+2ROxal2AJjBs7mqRf36A
/E/12H1FJIz2dRFtPgpHDOsBySr5uOrAENWZ9oxFkCS8Lj5i/bp4SZ+zocyM
ddWXRbxLofECD6PbsP7SXk53Z+4QtTh4q9NgGak4i8soXP1xUppgPiKZCcUj
GjXKRGPHPpaCvEa6HoJBeDsLUFbdiIairxnvjOyn70bqeGwZiYB5wS+BdJjA
iUw2bfIo7kwdfyOceL+gxHt+XdIOYn5KSgx4UoGB0mESzXNA64O/ZOS/vsku
a6Zu9MzUNvY93cEqMPT4BE1svgvFsj6DVswVMc6TBFITNwnwJSH33Aa0IuwI
vWrsoSYTxh1Q7qTtLMiSdtwLkMkJQZwQuk6WfYkyHqvI8fMVbmKLDuVc+lvj
XUDt04H63uMInJha9gl2g5EMH9shT8gOBWPIWk5B+VURs90MoOPQAA4Dg6++
WltKouaqbmd21/K8yAW/odRZSAVuoAdpIBGWO4bxIJIM95pctpA2npWexNf5
YvlL7WjOz2+Nb/xxf4FraLej2jCdVCe6wbX9IlSKjyTYganx3XGwAhrI0AR6
mV+TC4yTMQuX1QUAtnFyo7tb9TIdy+TBrXypJWuocpVRftuvuvUr/EEcB6XW
KcqfggAwu1A0qQkkLXMsCkeey0k/spZrwdBMbeLO/6gsbakkg0vFN9jFBjGi
jpfQGGkhKWzYc7GQvDSrw0p8wdSPGTbxeKSd290IK82G6OaIa+Gi5CwRMD7H
o7ZFbWiEMAGmDIxs6kkMkoQGLaSY/rJ7O9NQZusMoxc1OtSOJ6tbv2GmNq2t
2nJkBnD7Qk9ejJBNWab+vHnRkBUrVmh5D+j8rJ18QE7P3JNQTAhaomerjWc1
T01F/9K4GYEaSa2ukBN+LZIObW+wj+CghuDCI1hO8OAMp4H7X/pUlTfYUhLi
a14uq8seE4S14SY06MsG6sM9W/AHbyU3DVcLxK7gyCEgE/gLB20/cNrFUb6k
BhfxVVr+PRVLSBTPddLNcICQCQ/f9F0gCWvPoh/1FPqoBOHftwbNxe0Ep4LP
QekGppt9GXll4V1g8OrcF4AS/a2PYH6+kpEXR+q4Z428wYB80MgnTK2mnSTm
Wn2EZM72fsxwPNokbmeKN0j7VOAScvDWx60Td+e2AHmEMX7zPurp62vjC2sb
8pVcJAflD5kSSjAIaAVY56HpgdxdGWEa6rsSVjCwyUyT6eMFCLS8SL23Zp2V
I0NlSL5xCxZDS913q2l84jf2KyNak7S0DUMGyXm+PhHoyvhLSsC7jpwnM68S
wLrRhM4UrCTk7/nNiEz3KUOXZD9K1fT6KYaq9onl6DvbgokcmUE9jaj697Jh
ovQsouO4XvnmZhCSMIAmVUgyGHLR+LJ7HaRtm3kIav22MorcJUCTvrfL+K+E
Dr9ZnY9seSNQcJvX0oercuZ+59rXrO5CkSYKeUUeoz/5z6v5ALjgdtHi7J6O
UZYcIeHYrOFUpPqP3UTsxPmOBXsbVxersu55XkrgIKQ2NmzXcYBHQdPBJImQ
QyUE5G763UAkAFqTrgRYJx6p/Tb0IPgmqHm885ldeLDcC44zLJd3he6mD7Ql
utoz42c462C7Un03nIzVuT39FbRm9BB31wOnKwAgDZLyuboH7E4PtfOFaEQr
SH0dba1xaLpcmg3Z4DeQWur2owBgDruFyTHchcyeAHlJPucT1P8KKB4bxL3b
y/qOYPJsJONc/8dAvLlsomEPep6PUbv5cAGAA2zxn4d3ib4WBpaqfc7lceLQ
S5R7OEObX1WESfbdZKHFUvXXb5DCF24LegQ5k4DU4TYzosa35WnUeTXXBUPx
IR6NCAuvxE3QuSP4m1LEEr2UyQrEyUnEDyShbrb+EMagtbDzh8dbHSZepCLz
btVUWAIxa5Z/4Hxg6koIMGoZDiZWAFW2olT7YwCemAYlSh+049MtrULPg4gx
5oja7TsqDYooGahHHGWWiuW1AO46polkLcyoG4CeKLKUfvG66yIY7bzbi3dv
0MGLDMPqk4zNorWkzidEd46paQcXzyUuQGIk76+PXrDq182o3A12/vkIsA60
nJvrJE9zFXz04QFTTec9EfvaAFYtlWXibEIBFINZwL6fmdBPM9qjEMQKra2P
fAyKlFYg8ft/qdS6DKF26joVsAXCER+2AtIeNL98YG2estlr5NN3Fooh4ifG
LWZ7UCsrLeTHWW4MtbnN7EdDaGmE42Ardpa9WO67tuM7G0ExfaVsO/1nuaB+
W3h9E35C99dkzBlaHtorR+KRBHCjyHEXL5/V3cbZlxGK560MSEPYyk0aj4E9
QEDgSoT8yLNBDfP0R732NgjcqY9ChPM0eP5l+t2hBHVv8HMel5yqkmVn60x8
/WkF8KCzysseLcb4oRK8qyBQTkWxIg1/0j6THZchxDPOouYPmZv5rabaFlFS
HlZomiUAQinbJVGIdwAXTJkUbE3IKhCvqcYMATlkomKpIacIP6JYnwVtgQjo
gV4/OlO81FH1ze9aw+WqIQ/3hmC90EWWZz3fCAhYOZdarmwkacASgcxrXeG/
CLkRuusZ6/ax7LmYLGYDG6QJSM74n2MGO2f6eI9MnnR7lqZRZObXbo+SDacK
iDfJLiPnLkQv7+WZanpWAlaVEULH5dysieKuRaoA2xmUA1w6QuBgwQH/upNr
poo/9J2dp7mrs7by/VswN5Ki1RBYVyJTjbwHow7eSQiAaFmt8ZSpxxlWaFwI
74u6+QVe3w/f2+e9h8CGo21/Q8iFQ4gptz2Mw70VPEwDPzZDX2EqdpvQsg6e
mhs7Jn2BmVKRL+veDAR0x+MF+OjQczOOcHXQ3H+kzRNOyIJiQZePx+TgpDeA
tZammn5VX5z5Hf3jfzMHC1fjkWRcXEk6kITNx6Vg4M9Ss2XvRnlWBJ4UJPNd
3z0qiAS/MITYvaRHJRbiIe8L4oTJyjFFwMQNbZ1GNYL807OdRESV9u7DAXTz
lhQVrwqlhoamYkcwsGvv6bkjKO+vhMf46hPM4/G8wDMSNMQdFqJJ8wDsKsTZ
LZWu32eRV5A25jMmEjLkTYr+FTnO8A5ACt2rqmhCXY1HV+GNLp1Im2lB/xHo
A+KofMso3Hh83zywhsIX8alQL2nsaHLasPwff0s3IInsRPi3v9sMuxmI2TtS
3N7Bm4cniLHgK0UW78XurPoofnVjG/J+Ohs45lhPFt+1NMWQ2Ocsh++dvdrW
+71OPAjyKLzKne6TzB+CAa4Sq7g+91HZhhsytZvRGPFPc1nPvON1cIn0sDUc
pK41GDnQ4ETNKO5KLVY0lZlQFdLEnOrSw9QMuoLPCI0yt1a2guoPDRwPVaNd
yDpCR5yX+KLSsbXe82C+l0W+ChRJaKqWIWnthDErk1X2RPbXhA4FWBsoUwa8
KVhygf+3arJbayNOC0WkYdnYdUsg7vbsxJuz86Y6d44YFkXlzGSHFlGMa3nb
HTJLbgiSoyT64zsO8/ow+tYXSuOcHdYUWf7RbPisDUdQULasLjt99Zk4BW3q
hpwPlFidb/ujPq7SRo3Af6ZJxLenaIVJBcBOUK8SURHH4BWcmM8/8cl1/tPf
NHiWizBQYoa5CtXk0y+SgWpdp8kQUCnfATOpevaIABanurj1jgY3hTJlV7O3
/hQFqzI3eCjW65HZ97niW4fpbOaTtOreIIOAZ8kL1kx5is1vCPCFFjZQaWsb
kY6aenCQdp6GpRUuF+RjeMfhj9gxYKyPBNeh+DzdjvSimf+9MFJdgyu5k+3U
C0xbP/TuL474i6RoPYyxhTNKX6NEQiJNUXraMlq2e12s/rIy8nj2uUc4Q6cU
ZTBUB8zUYzaod/NiRasfawfN8DhAnL0SvNjOysqSznM2a2hMn5+Ftc1yWKIK
wU9gvx39UpS++PXIwSsMJGZeqIcUpMczqXp4PsBVRW4B6dNAuwxvSy4qBJdh
hWEXJnXuiqJT0ow+Iuvzn/1h2bz2DvOLqZBm7oi0Qf3zwmDuP8RBkWRlAZhh
r/p2VleH5Izp1iQjb5lqJn2ud6VfVhA5CM652T0Odg4Qm15Ckb09cfckRByO
W0iguep/fqWcxLGhZih4dc3liJVb7VW5KZj5zYD1Pl6Apl+PL5XTHtrNrm5P
+SpG31Yj65pbwXeWh774VSw0oOmJ4GU7EBMJzJnSWzEfTxjaYy4DDnXv6J9c
dYSoz8mgVUOPRkTwRVxnUCpn9geM2ZUk0A2xoYzQMfxpkDRPRfyjSoOuhP5V
o+Kcezf9S0wI4fJ3Q2m3CmP+ZJDhyrDAgtO3e8ULdSt91HaJO7G9Z/AFaZxX
G+0GbU+O+1r/sbubxRH7NjGaN5qawAg0mLltwrF1UcfgIgg1TjGkt72ScCFT
p/n1exAC9Ek+RgBuX6+g0fc3DeABRwER07paEX31rLkfC4fYvhSSXXExHxB+
6AfBEJrZ1DCtyj0N+Wm4YTqrFXZpUt6qjMVBXJA5Gm1G0Iqb8HwOXJD+IWfL
3Uf0+Iq6wWlrTqIb/3C9aPUkZ6NcXGR3jpf59UpABxNXcgB8wQIeBXcuSJq2
3FvDlGSGZC/jbSxsR7Kz7tfmMus88F3tkncHLkBKNF1pIbjj6ez/wheQFlHi
mVikTyJs2MWNGwybOShpY4pQ7qTeKjnWwFCYxcHPitT9fxajswA51bfdyd57
QFRA3hEGdmeHbm/8haAdUMJnfDQCx2DDhpwtdJjZgNldWAeCsb+XPm16SJZ6
OPZ6fODrQURPCuMpcALKUAl2d8v3Wh9mc8/CpOQzZiyQUWmxgDCF8mWcrD6l
51Zqu7U+G2uwkeGSHF2mAPlOyhS1ybciSHW5UNdpKpjIsqTjbGBmbhIdNIpp
DRaFHuDfV0TwW7KKW69gW/FgKZJFut6wzjkhCZStP8KaXylAuVDWwW/R1R6o
BQFnFeUSt9Eom2Az+i80O+0+bRfHbqRQInduByvE0tzgR90BZMuO7u9FTSz7
evdcQtDzu+/CSnstrjM32aVVZ1U2b7O+vToiNIV7WniWoEd6DBIPBNcsf3HX
CEffQPKvJqrBcyt9RXjkIH3hp57DPTsYs3eXqPN6HUD+HyTIwtfFhPpjW700
icz6VWejm7O8uuU+WZQUKxCzMgnd+eA/KcwbYvlvQD58vY4u6wQhcyIZdVUG
JQu38EvF160lude0IY1uinJkzI9u+sBdCgfA5uIxh5F/7cmt+dPiwMTHHuKx
7vm0lsBqRFt0DdMWXt2rlVxQUHFt4YjPoVee3QmwQDi9G6np4gSi/clzGyWK
tgysxoHjHI2bf52/B+oqsOEBTedXgitn7Ikx4ire4tSrpZE1U9fYucDncpUc
yEQ+NpGk9qpr5BrrewxRzy2cFVfzX31Nzx1QhkKy085cfQKPheL900PhMqa4
iH6JcZuz67oc/Hdo0/khB3128x1Na6djkc07d488LfetO3pjajXydftdACrd
Cd10dOmC3nJzQFVuHnXvTZcGKdltN+Fkj+WHlZEIvf5g6jregQHN2tmgoAnT
/wzI6d9cmYG/2MPMEBsbLIO/rt1vlhMR38zKgFdRHIkcSJQSW2TDZ/utvaQS
sGVgjoxIkXMCMMAQMQdQCs/1EbqNs81Q0YmTNFKDqDQIjRZyu4+X3lQ1Ggnl
8CVf0SLsRvWMX+V7qj2INTQFkpuKS4Y/+u9E9pyngez8ISjPSBhEjSQMvciR
x5y/Y73o8qwp3NPJdJXNYNuW2x4RUjr75TtVTmRDIqe2+XtXBrHZxHslDWYZ
XBP45qktxh39tm3ezBtAToCtgitecjgOmYcbWDc4XBN/5LvSy7YKbVWgjJLX
wcrFRu0XxgQ5n89hnx2N8b70PIwPgevSsuwmWTmmgPccGO9TYGGGCqRFQ8l5
gFl6r/wrWUkMBNY6S+TN+N3HotKb+TC1HKCwk2XN22Sy7mHqhSssZJvHgPUl
mnR3d68NsEHOgN73bhPVEORI26BOcoUOVYeXpZUNeMI3lMx7a0Jdkf0TGoJc
z3mRdpIOy7XZ4upKpuqhgtZQKTNIjcng/YHAXqQPY5T/U/VpKflYrBelup+k
hp0ZgqzryAcnWT+K6gb7ff/uu33hFK45MMxjC265wFbxPEm2i1oK7Sc+nS4D
TQXubVSbS6e+NubkA1HASSqVjQ0fhQhZRstiMqjuQk4Rgb0GDZeeqltZJrNQ
06d31cXo3Ayg4UUTur3yoTiCxRD6ZPasfos/SCE/MePBKlgqsmn8HbzCjHDC
lxVRBdc6I5Urk1P8XPUkJaZwwGvszYReiK3eYhG13pz9nabRau4yVxonWeQO
+lVi784jarj6klutjJ3xspoiLkI4Io7BNPaUdQ+JmBi5guI9iKGtJTYStm2A
ItY73DEdrApIcdty5HPz0W9N9WbxegKaQlXz6ZRP5ztNxbcEVsB2BbLVrgqD
QbMRPo0Cw1SJ0SEV8CjxvqSY2jQgbP6rezR7kBSixpOXOl+6LheG0IhO6B+x
r+z0yjMiUJp/l5SDwzZwoDpvhIaUN1R9o20QHC/kGZjsmaOv0o0sa/fQOVPo
4mIndIaW4l1cNO2wtRMXo0UPAIrlGwA02KvlBGLrHTz8CmJgAKYs8jtY3lid
SgxgvwihqSAdXsi12z5swYx5fdhi2Eof2rSBbAayQrClELlla160VjK/V3/T
G1GujFI+TcQJcA7Uw/1Vowy+midsvuSK3GCp8E/YxUd4aGzcYpLbJu8Hj7yt
oH7zrqK/cTyJzd4/CilJhsgSOaB9ma7dWmSgBjIQmBbv1o6oW19YToDXzr8Q
XdtVzkxGdjdi0GPrFcoa9nt26TlgyYm4JIVpeC+9/W4RwkzQmj9FebiNcbkm
E2Q14iRYdWaqturxUHUJMUS727DNg1Rudqvj03v/2uvsf4pkt84NIS/nSSEu
A3qum1rWCROo0AMYnmeQxw25ylJp40sr7Y/81EAwmbCCT5bzGtDlTmIfixVM
xm2CV6wAFZkzm/jUlxRNUjACjdbK0PZ7mDEvt6YIhgQ0tCt9fy7mjeaiNMRP
hxiRnMmhxjt4zuZ4Un8wTcNrHkk6x2Fzh+xQ66lw8n3qH0Zf9hFdpf5Ev0wv
SDpTTQ/Gp2TeJjtpwIT8zsHpZGwKSCMFY9NzaMuZZC93vzFiGNGwdQoh5c0t
ghvG/xTHWLS9JIQrYy4Lvsd0PQbgoHYParyPULTrveNrMU5jn+dxQDfI5gZn
FqfavA8g+/vrNdAMCvTVTtqbZpplgW1cBEajvkhdjR9O9V1WH+Wyu4Wgx+Qi
KqpOgw+7TCU07Ysb8WghLaUcH1QYDc8fJNNWC/CGpAP0uVKlwZ8JUjF8tBjC
9eDhu+msC94VkUP46ZNjXoQQ0Rn/oYah+Q+KZVc2iTdwEc8rVhso/w5NNdRL
rqEgAlaY71n+fAa3R+SLs2yqY8fkbHBJwkn+eVJxxc5ZSym8SqSQrPPIYncD
DUYPLKseMCf0R7aOg7V1Ud+oRpvqyAeO9rpr2gygVhAHNTAqN6lH6U5tIMIG
gBzOlYgXSFCqiN+pIyyLriTfyVL9unwDFWgPi0JJI942kslJz5DuLrziS34r
mf09fNqqCHfNHnUlAJQoIrhSd2+7njPb/YdZEijWz2amMDq/Hbrwyu36D8Dm
pjuE/STqvxf8snQPoaYS8nzyJu0oNS0tydnE9ugY0UxdtLSg4F7LTfIYXhN8
7sj4j0GWNHpNzTxSLhfZurj5VhwbwnxoPB9JdJGc358wsxLF5h6VtX/0y0g8
AkFC+5fWfoOSTS8eCgQK1/mGJ7QqeySRW7ewrHUFhkJ5hKrRBJJpweivw3gM
8OYRAGaSnxZvVmUpeZdZ2n98vUqOpaQbp/0B0pfLXIaKlGERs7tahHjJXYSL
NvI+K11k2AqwVGy+1zQY8X6GbWHBpdoFZwEEg6W3NTjVXZ6CJLswwh24mGt1
nnbjudW6Yxx2aqL5SZEtIa+c198Fbe3KpIcPmYIWxGhFvrVimGZxv+hWFlwU
nmon6TmIom6RBHeCyKsxmGLaNsPf9kQc5wb7y3bTzccgvozoI40kBaxgAfpf
OXpC4BO10oEGTt7zWduq7IgJosdPb8Ivw0hd6IVWafDk0PoVeC6NqGlS0TUt
iCCDjniF1yP9WebWpLRqF6T2VKvNR9R8DqZOx3CskfInO130npEbCCyXgw7Q
ms3CkOBRDuHBaSqSlF9v2QOd93asSjSJrYbkVGgMSjPd2SsbvYq8p5y7tr3A
SJO1gXTCAcONZYS2UXLj7tyNU8MT4X/zlW26kODXw0u00PaB0Sdk4Rla5y1q
Q0OWlVzhdD+9oSrUD0n6VOdj/Sp6vNEbVVqQaRe3fetvThsDeWa3XDqyLg5Z
SU3BBdE9Yxp3riOUQvGqqDIacNQMFn0IxnNA1fNqhrwXz2bMv/ic1Xg1cVcr
36JwE+PqXYApOMDAm3Pt2fENptesx2Czrprelvf+ro+AFE7Tcq40mPQBKBsw
3oFgtw7lh1/mKg1Dzvm7Gq/Dh4K9xFijTIwJqzAUxFw2z1i4Pz1oV+5atXO6
xHF4EWG9zpDJiQk6S/Tum7D8ou6otdeiR5GccPEM1hseP7IiZv4eKi2FrzP4
4yzmRJtVmQsZNFD/sXc/L21uEttwk81lF+g4c28/hfLLQsaTwUwZSP9/I+T7
xpwJ/bIAMORUQ/JbEukEBDGqb9UR88WB8Arzn0LD8q7blNuHJrEbJl7sDdWE
Kfl8I0exuHNhfzivybXOkMZbwfM51OJgiXpjckjqHI4xog2McSK2LvtL51vs
4ftHApP1sr4j7U0CRyRSwGMlgcaKaJZx74M77LccpWFGRoLUqo0cpEJP5JP2
1UBsRqHBSQtJu4wj4Z5xYW7uyhb8U0fhX91t/VXkZKHgmpzG6R4MfmjQuaF/
OkiGQo1COki4BQSgAAo6S3XpUPx/Iwx/t18DvMBrbBTHQW149h2PrWpej7zg
7cKDRlfA/Z7ijh/8CA2m2JSG28m6ORap39VYopKx1dI8Bz0KdrdZlbUeMDqB
EoYGkodfeCvY0mR2vQkwfLGH6yyAT/Lwr1S3Lau+j7iuHCChUohodzfwBOvG
PnaeQ2xL4ElV2DMDQx+CNdmoOLENG0DFD3BpwVd/hRNddLDZrMFi9VfKU4xP
hNFSyqOKArKlhnfSQ3bMWowUQsklpyOwd/OKjdPWQCglqk2BuaU7aQ1MNsYG
SmhRdOQuZz4fMnUXgLSb/5Opxf6uLVz5ke/dHm+jQw66iGwSkNiaY00yHBao
baDivI0rDNAwDEoOZVTgUKxiSJqYiglXrIwwBBHOBkqld3kLnUU9Q/6JPjqF
7qlNL6ODkk7gDyLHsn38uZY+/1ZVtdYBYkKWznJPNIoQ5J+VoyysMSzD5yl1
FRNU+8yzmjgxdwQantvYZRlHXBzcLoHiNfqdhxrRmBMyLL19MljYpSI4cjiI
fB1FoI7NJPlQTcuacXafxlKr4MtCJ26hzgIW+JqSYNLSrqTxIWv9pwG2Z/3p
F2zMlRbHxzB1Ya/J7/ZkA9aS80b4CXbl8sixtciI0wCWQ1adaV6EYokPIREP
EB0W7Ys6kn0p44OnY1UExcA7qcfngQTsJhn+tWQwzrLPGDBnSiVZ8IJZ9Fcz
KQU5CorAsF1ZRmO2m2Jm6Fapf58dDaMVo8pJP4yTDXwbROIXjGl4oNoeLNuz
OpZZFaQtLbHlyvrOlo/9taGbBTntTGtOhL4AYEtWgLLtFtG+deZ6a4CKdVIn
p+em1dqL7ZdkxY60RbQVjPRW+EFRLlqKYFfzqpXyWJaZs4Ugm2wApitsd2oE
ItKHs539/aC/FhfRadF+uhWlh21XWSZUtB6G6C9nuibOG9sHdUK2XnjsMnKE
hR7b+/GwWr+J0I/aqSiU+UFZc+6Y2aXHddk1FNC0kAFComkRhVwOhydiRvD7
eGIvGfQlzNK+9R6sxwmlKAoaD67XQszHNJQet0+7a3gyjF+7RPTkBCMsI61R
oleLrKXPv2D55jHCOUuZsGhcNxoppqUK8mkRMmbZTrlSd3tXbx0xsyy2ITwS
s1vhOHR8aMjlExFbn7BXEy6jd5I81mCuPs9vY4Gufp60yStP6VR/KeuKecLT
NqBYriSm35UUJwoEymhqvTp1wYUVlkV4LGhPnRF3ietB4zFhYjRfZDcasHJm
5WrqHgC/KYJPExdTd8vTX/UWDByn3w68lI/rYK9v+7qwmeyUE2szfiFVB4b+
ln+F63w/LWWaAaSxOr77g5uH4cYD8vzCVNxMr5hEEADcJpnlyTqiQlwz4AaH
Pfam4ffTtWhrqrNS/ZPGjeSSE9/wy578f5M/EVvdCY81Jy47SGsAESGCZubZ
qlzWBWHZVaNcKNd4B6pqG9uZeaz9ANki5sWnWD79E6f2MA7AEqlWiEhl20fC
Pf0mhkvadBiEpJYsIJe3x89vBkITnMs+kCRep/vuXpHtNVo/MHy64JcSMWnl
p+EonjWbix/yzBdTHK7XKp9owe4q/FnekyWocQn5pBDVyEi4bXJXucinl9dG
m6JbhdzlqpVrhFc85YSpuZxaTV6gfTyUthbD90XqFP+kiOO25pRZNbOQ9/NZ
um1OkLlniZTqF8s6nE5g5caMae6/P6mbb7EbW8z6uGbNCRlEEMmAkKqoSRJP
XMq2JbJc6mtzbXla2UOzK1AiF7aQVVhNQT3DyckEpwlOpxMTWRw3/mYr0N1f
RgfLddA3CiTIq6yC+BMBfYNWO6faak9dLN+83RMJrik/gp140wRr76M2LLdW
gtq1YC/X8/r/2IpqT42h4Hgy8NRbzY19YQhQRB2D0y5TqvF+2IaCFAEFDVat
KQBax+9bO8vZgvy3YKYaMcqx6ILi7YdG+BIV26i8bVgRf5ntzjGN6bQz9RRJ
Nw7fjDQ3Qgv+HWyGXFZjghNWK5J9sIpzDuPGHPvKFTqN5JWDvO0kBG17S7F0
+M9Wbc3fTuevj7QcDvI3LklgLDexpYlpj75lc8XtOZ3I++FeCFhyYdXDU+ZW
/67UIhMMyHSQSO4SSJAnwFldCh40BW5rggRsGxY6Q2YvU4b/hraaDXAvMraN
o4wVPTmWe0HBe1wjwZwm6Ddx4PAEtMkxuQsbGmHulzVPiqBQ6hH9qhPkxYQh
l4FZ5gmHSLbhwFZfBSBCXdisJie+hBT1BwUkILGOJ2ENxXZoWS/+xexaHdPI
z2uC1fHZenWRq1ECWujXxtOxNvk89jm38aNfgOCQnjfNFaaITgm7FpKCfyf+
FbD385jRWTH21KlL4dLZFDXI8hKil58vCIHOEe12ENVoCJOtm4w3CWiSrHRv
/tZHS44v/E/Kvx+CLT9reVnQZf1F3KrmReHdjrOMph9hMtnmvcLWeM//y419
Ma+CrMPu7g0bMiTU/YnSpoLWhgWNhayx+RTN+AP/TaXJl3YS+qaRmQHZrLV7
r4TKyodTtt4HANFdnaMx6b6XB0tT7dQxq5uTxghInpr0rnbZZNYVJDgkjKYW
mDTCBeyNf2p3V/PCjjXif4R5M/Wq+ulkVoqlMdvHuXDl0FM0p8SeMudy03Zt
1BjLlMrr827A6JnLyyyXHoJ+CoB1abqPZiAeANzQokKQS1Wz1u5XJU6vVgJR
wgIKcKALBeD6duEzImjpxn8aNKHJz3X1bZ/NKr+CAoyA4MDUHrelMbonjQyN
TkMQGvz0QFET0n8TRpd2GJ9sHCalzUIHv/umFIJQBvewNP0OZULX9uQnt7ST
ty5rgb+lNqipkG5qZ7Q5aNqPtRkSnfNuHabRt0Q8HzJ2eERDaG0d445XMdlt
ChBoz2jgV30kPP2teWUQnEE++yg4SC4h/nM8LEYmsFHio98LFlr1D7LYxUia
lr3bx2BRbGDaKhhBESkg5syExb6RQW7mYusM2vuOvfDWooy9YQm5BiHMlSRv
dBIsrV1l/ttOTcyHoG8XbUAUCh8LrU/cjGLqodycWdHPwOK+bp6zRHA56UcH
ExGiUgUrM5Y/9G0Uw2GAKBMXPA4gz/cacdViGXa7b7M146QAj5t3tclzMxv3
XNFvLSCQIaO+Rp46ramAYkfchARVO0YwjnYVip1QLFJvycYHRDMJp2ZqBbBn
PlGAnXxGH3ZgdaAnKz5eX5F29O5mbhPi3+jNFkfK98l9zr68ff8xZXhl+xIF
JSXGDkc7AWSbBD7yekA4Wj/CtVbbOFqs6jHj/rB4oY6Y4cEQ9oeHYDo14R98
UUXiWBF7UU8dP51fU+cKGN865Bphy/DN3B+LTzx07ap8RWjdcPM534lM8Oqr
1C3+INAOqQEgGv8rgJJQcC3qk/fgWLdTqEQIP9X7jwtB3OL7Ex842APKjj8I
zPFzJcxK59weFZKmeiaEuzQgJkHgDZ2qseR37eyigGiDAKkoyXCxBmoDXTWv
Qu7RwzCuY2+WRbWHlm4URQ4xU7SBMfBfwUHM09YEvRD5zibP7RAfDLRFPfr7
GYtyD+WbDGL4aCIZs9r90Sc3lUB2mmK77U0nVK2HZPXwdDqe0wksu3ri/fka
eOpOZ/ARlGxHbLRqT2mis4KAy0ruO/a72+cY27h/8VFILQhuGKG6f4Ddr4if
GnPajYGwfaL+q4iO4BuTeOyraQe46+Nvl1pQkM7toZ1UtLrMU12rpL6+odsN
SIdTisYcwFFEy8fY3YYwgRscoO9rCxDhr049k+1+WTYCK6pyjEUlG0G2w2Cn
tMdwsljgPqAbqkDM8/yncN3SSM0EHkTMuCCQzZiVRw7RpMsj2PbUziJJ1iLX
PimxeTEaXaaxkiymMif/MX7PZ/BvuPXsuE9rngDFP6ekV3Lcr9OD3NfidY4y
Xm/LZzp0exXkPFrp28heDEyX0mcvINxdOG/HiqXiT81VJVC9/Y0vmXPQWK2x
5sZpIaQf3jsOtcAs99hZ8HZTjpa8K6sPaZslpBoBanN/3GQToUSsVxjGvq5R
e2zmVgqvnDnpBIW1D+KILBMC/3lJzxNMsAmYvovWRzsjMvd4mtajgRIM5QAs
gY47pWEmDZP4VEzVz3dlUJqCH7oesYM6Mhnogx3tX+vAfgrbV/PtwdFvf7xF
3VpBPw5iCXajNTBPl+o9s1WoW1BjVE9cUUrTIOV/nj8fjyYQDl8W1jD2Xs20
F3BqDdxJoaMJf+D+gWyeKlHkKC0Nfb5psx6As1swpqlwwY7OVnSa/AZdkN69
IzBHXE+OYrEmO52ykWOYWKawFtiwb/xzYuyhN99YQGu9MM55ws8lceHnQpFB
Fpzvlt28vg1utK463hPdy9WOPIydGQoFw5QPua43s8q9ePwjuOfLDUugLXMs
pEcyFPbFzxlpQEojNpGCYz5nM4iFUmvjfwMaoh8hOA06ltdeNVwDsk4ICP5m
uE4QMC96dMv+SMZkucxkuEfQ+wguNupbEm16DTROXORYP6QiufD4+LS9hBQc
s8rVh1kN6E9B0wtOWVvZCNvcr64rxDsrpdpvf2d8sWXwusYv31xPxbZV9O3q
Y/qwubXw8g+RrZIdG4zQPX5Pd2VuyDo+9AodY9S/Tdw4vip7A3U565Lb5VER
nsTD28qeWazm89N9E19Bjv8AnMHEGVwbOgdp6ir1guBg9wfrB+gGutEJBMzv
OCliNXfpYa6xJtdVkxdNO1IMaScUzx6aGdmbYivs7c3e29sweUuVrrzTkbhf
fmRSX8WOKNLZ6aHgGig/RF3dxSolNdcih+jfRVMItcI++/MdoWH90VUWs6H0
DI6r7Br2nRvTqReNElmvg2lWZWG7GD7i6rYjwQry60MBktYBULkA+YpVB4BZ
Ll64ZRzB4NmEjxorZ71sx8SZ7lfWTgZMRUmJ02b0j+Zho+W4RveeZ3KtXC2i
8ceSBhBXnwCMpmiLznxGALLVAdaLQmBzf6/eg4gIKhQZWD3rIPpK1nqurCJN
2U8FnRQWGMOu/GpcY8PEOZ4pKxmllmzDAtRrAzyILo8eax/rTZFENXRyxBTf
0dub0dt7/UBQzg+3x1zETVglq6BjDslD1i+9pbjYuoVTg6XQ8E9yRAVVz8CP
5CVx8vQezrV0Die+YyPkC58tcY/f4PLFJchsVmWbxXEaH6YkFMzoPUWtOzNX
NZAkjw6R4IXn/3CpES2IrFgth9wamJmJbaBqQblwbUdFHGnXDZXjksUptvuM
tQaTz/Y91YTImiVigwWloy/un/22f2hJKNstVOfvDWkuaA9Sz7NZKm7CErbp
2k7IrUe9InEmPGqfz1U/oc/JgdLLY07y6V/LgR5bqwVTf9SZD5LTDPgZWQ6G
UpKsxadW1P4ei+JBTv9K75siTH2uGhSqUYgVIwJ2tj+KfCjqUk2HADdUBp6S
sPtBiq4lst408N2WYus9lNcQ4kB+Tu+P3h7LylyfBpuATfT2lcp1KGx0ZIG5
fe99hwOyscn1vObN1FeAfzvC1G7e9DmlMmyGrx+qZ0i/bNslVdqncD6xgD8J
3WWUIIXjL1/YyePxAaaURKF908co40JerVqWXPNk+ypXaAh7ZyKCCMcfGXhE
Xt8n4hyXMeGEizJhGXunK+TQpPCQCXdPro/3yV8/T02DMLGdbDAx+O2aCRzO
R8Nx+S8kibwRLysvcPItuUUYyheJIJ6+pSQHSVTpGShCktQTqhqIE+mf9ItF
VCKAYjVuW53jZdx774LfhdiqGQYZ3gyDgh6PawWWK5AexoQ+h+r1C1ykXjfY
FoQ9GMhs04a8v2zEvqBHj5qUgO1IXFDlnDfFRg0+Fv6uMYeTgnicuTGcye5j
BDeetrbIOvTn1gIWuwZIkc3J8VbvHTnWobgeAJSxLKKiZNgnIkxD2OIqxArI
LnIFkKJGvA/Nj0nrvRO0lRuHuSwmgl3lsfO0IFKx6CM82ZF06FRgTEg2oj8l
iBalAjEOIdT+o4brPevyq6gHT7TEvdnk/viab9irBRS0dLaUk71tWjWF+IMq
Ayfr8eR26JbKUhYJ3IEpMLCs/BKF47Qim+1fwRIoDkkhQXoT82ojyA7JhIIB
0wlXopv2TSHhzlQXHnnGrjFAX9EzSXXf06Vw9g6Qftyh2bDbp0TW7dH0DVvy
qWhl15BUUMr82khpYTKOZ1R2TZ4thUo8LsrrsjklnXtKZuXNSORMKf0PrJg9
DHN2S4g9Mxk6fT/fIGQtbv88ARkd4Jt6ieptB7u5lbFxWB97nPAtlHhQnqB7
qQYgOsI/Jo6MxtqXaUYOytUllPj3XhCfztVAztZVmB0w2BL1vhpxIt7deRmE
xVmwmAZhpNy/2TuXeLkgWOU1i7wuUMOb0drCWa25oZHIR8M77tvRL3WVplRc
ar3UhriE2EJF1Bsfh6vWt2+ipfeHhRACNwF7avdZ2bDdxLNr60Ahp7WhmOPs
acKbVVJ/MwjdJHV+Ztyc13T/t6ZL8vdsv4JWwzuzicjxIf32CaOxrbQ75l+p
7Uy8dVxFE8uL1zrTwQoFNlLJQjxkBKOvHKIgeS6JfbxkR04HdKj7IC06UX/c
VlqQHDIf9jJSw2U/xylD1C2Jr9qfj3rVqJcE0HlCJvFOekJ18fWlZkqwIHBh
8P9HunQnrIzRKFiBJ0YPlN1GIphc5yz1xK+zOkjOkzhoWByWDT8PgYntyZyp
4pAJFJQuDPI/kMcAWn/CeTvLWD2vJUGcrtB7cYjgF396z2YtCl5QEgJoINDX
VjZ7N6Kk69evhr0LuyT52VwOsUk386XYXVBmXFKfeyglMki6Fh7YzmEqF6D8
/MICc2J5XoXXVxFY6xKEOIZBO3arDhOryiWqrX4ePcxckc65fqGNPGFAB314
hbQ1Yao6H1D2GFplrDmPN/T8GYxfm9RcunlGYUQjugH+LmBW2vp1H4zgo+4W
dn6GZEZkSyazLouAVV68m6/J5pjpoytDPfmfhULhQxqpM8Ys6Hn1QnREqa/0
NwBUu5n89cQ1wW/W4OgAlcv82/TPGVeTOAetXvSCdd+x6G6b0Fy0+TXN4ioj
Lc8FnILzuJGVS3CmFL7qhpaPGE4ZK2/2SwPz/QN2yTu7/jsVa4o1IKCNOhpl
4zdsM87y3583PkvY0OReFGszLyxR9QDVMmpJqhmLUaoV9Z3T1iGsh8yraF5V
l2ADEj0X+EjMpyXt0Z8770O2Oz64MXbGN/brbni+mgzHIqJoelRoWmBq3o5G
tCMXfr2gLAcJqgP9UIkDV+btf3OmVimwFQDDacpA++8oDMkuJf+K+7uzl+8w
fn7TS4jlQP48sH8BXP25t8TMUS3TIOmZyCha2VGeNV3CZxbyE/r2KVrajvuk
WyLz2mGy2+sAOG05pOtHCJlanRK8KtlzJLwcWoxm6Bfk20vyBsaZH1sc9Hnr
/aqwJCequM0LHnf/SAZ2YMZmCOk05bF0bnUhZRPiN3n8VbAJAVhp8Vwzpyb4
KPeiILxpj5bvSStZnf1YNKw76veGyweBspYd5jzURJD3cxYBgymF0ec/GpRF
4cGMU/8dmuBrkP3zs57K3SAgbI4p0Yyp3+rn4FcdDe6CtcTSOcNkiSy0bRLX
VK5pgFXbSjsjS/O4uUlmZdsm5sSuWgtTq5hWWq+acvnslB+axBhjV9hoUQkl
SOuX5ZhH2pHG0gXZ0nzcTvzxy3hEa72ehZEihgFmatNLGLJbK3jGOVRvdwg+
zr9/VyQKi4x5UAicejWP0m8ZlK5d+fRSkBZsk0MOAhv+7LWMLv7mHnJxtWXB
b9CZuvXjTiBnKL9HNWHinBfyz7Ibt8ov5wzblTAXulunR0Bjw5zvigrH8599
/9vANDGpWmva1tcD6uCc4Arimqx1kpRdPJ1IEpiHjJVzIE+6Mw2tqHhtn12h
2ElVTdYTw+nbRljaT/YJjLGfxAo0LQJY8k43mpTdkc9PrHeMruy71Tw5CroP
rSitUswlEPQ2r+c0HQihvaEZyRRJxm3ssdJUgHiwFafFB/W81y4fYkc+tO9J
D8xoPKkNOhARFpfzmD2R3j4d3n7dNBOb2qbBe36COquI9IGRUtCegAI9hRJn
QRKzpr2uFq+/t17mQ5bzty+5iW2ABb7HRuo9cwGWq9qlGwynN91fnGlInin+
+oVwdOSmvtNzDPMZJoXqz20MbyRGuYQvs8s4Iye/1RDQOR7gBjepbfBXesjx
w4NIZ7hk/B1E66kOoQqAsqi8kJLbVYW8jew2kuWfYxSxUXX6C9d3+R+w4c1/
tcPk1Q9lYKLORWAgIhEh7m1yf0t4RnQvhRIU48+gS1iy4vc1IObYC4dkNVSK
ahKyGoznmigCR/vYCjhcxkzJ8472+NuVw45z+meCMVbvXACerpVZDvy0mUv/
nOYdcEAzOtA51WBmpYhUYTGRe2uqgqXiAGnhjxG4Pv84cXdqIg0o8iwAt9M6
ogWgr8+DkYVmEYi53WdmIxRRHIkxXBiHXja8hQ4VnISScPrgpQpn2jjvr/bU
rXhjxUj/xCYPCItiYYetWHsAbe8LIbhD6j9z9IVe2GPQoxt0OLfuXSY+6+82
9BlakkUsM99Oopxb8a7NGWfb3MQgivjq2aBChZNunBsNqQzLuQRCg5Ymmk3K
0kpTzkEgIdWRXQ6ObbvFBDvyNQQfDsjLOfwTpiUZV1CPDDcOnR6H6iz8TyOm
/poI441ibSqsmNSqEaIrF6fT/E6WdTwHWvcTGVgXihBkYRJofwQxLwF+tKuv
Rfh7xwKT1X19n9DlSM3IlMTPUrbcqSeSV0bje+EUEqiRjA101gKrsgH7A4nn
82DI6gtZO3N7C9NWroFxUgkd9+ZxiAtZvULLO5EmyAz9RpBI73Aey3hgsMwc
rmap9UCK4x9udxmXW068rRLY2LKYsNw+0NuP/rGOfdO1GurzsZEWC1B6LnfH
67kEahBT7548HeKYWwMmTottPeI1iM6IN0idu7FUktqW6eoCjk8/fXs0cSPw
rG4bnNz9MkS+U7ldDoE9f8iaTc5dJNKsWfN/oEHp7IjRmSlNWmRo1kn6WSa8
Ur2f3IxOQ+VEYlDWqCe0f1ROY12Uxh6oQFB3vEUnVRF60uxgiJ+J+khSQzDE
TZQ1GEnw155WbG/5/gm67gJSR9+1JswpLJL/x9ztlKIE7jiutsmpMD5Ri93v
q61AYQTvW4a+oOtPRbVufhxpgeEUAB/TSLSFO6NzX4Lab+2KkTZcCgFsu01d
gvB6adnZ28BOCPDd6XLDjGaEOnOBrFXWyxekErN87QYXvHTWTnnjRvICuENL
AA9LWKXZ12eFbfXK7nkTdRCsWKJOi4Uv+2yTjo2DAa3fOLOjoWOMhBQ4dYBH
9YnDz2ekHZy4Jliug66vPrucVEwfPSKk5/zjETZHZQifjpe65OrFxvw8WX3I
0MtUNkbWrRpZcNdk1BGma/2LQ5tesUEfTVM4uUA0i/cSW/JlC0AjBCxNKQ2C
kFdblf5+S8F8S0A7Xuhf2SuLa/ZhMs0qfoHS53NG4LgxR4AQ96dbW9UrfyZ1
MS3G7VBOdi2pAks4kvYyNATZJOhgrVS/QSbdr3lnZRnMNNlCZJq7I9JTTETn
gaxyN5UlmWoLmp+o4SRTxCzgZdXy8Sjg4STpMEeik4FxMZp9h/dS6ugB9xAZ
3y6MgciBxzHkDpNMMnAxM5mFIYP46yN3sXWZkIpTQVQZvq9o2FuxLBBNMU3j
Xq3rX8+eNg7FvzdA2L3f5bIP7084zPN72EHPJa69+cZh5rIPRTu42nG4LnLp
dyrpEjE/BA+r0aYYcjkztD3anilumcJrEeD1yBWmeiWdv0RanoPTifRWyhOM
ojFH7nqVjgLV++rWi5DTb9QCl00uJ4RmBp+7vFSrLBs1WtVveGm6cX8G3t0g
vZ4fZcreFJqspYv0O0JlJ4SvN7FdMBpOWKqWuMz5UE+Jg+7N8gSWGRmIYc7B
Io5pvInJRz/bH+eofVzNDexyL4O1Atn6coZtbOGjPggeDd6By3n5O+nYxtBV
MiTo0bPZTeQUWxp4MlBuw8BC4N7LRU7X+wZa9CKoFhsGGtKh+YNpBiJlXOQZ
x5PK0PrTnxvfaTnq+UZgPswhbCsAKNl9SXbFAZGbjxQS/YDugwblGQQxZMpT
oDU0IY+SO1gvjHDCshd5ZvTzjjYiptrdm7PHXSOoCXOa/doWRFnP5OQhyXhn
Z7KUu7De9XingpKn9KthbzhG7wZ4X7RqSNBvrOxX+vB+MOS4oKXOy5OvXPDZ
gsd+sq4W4iPsjvzJ4JXdMZj+2x2Z4QKW+JENiguh/UVxwLdoOirhAvtcq8+Z
vNRSb1YqWlMh/C/HdFTVP9JkkwTwQYrldLDWx7DXRejoUwndYDht2UCWvCWa
dLjs7RR5FLDHoOp8egsPS4WjYJSU7n2D7iMORKAUs+U95zfGsmYcaNL9iwnb
y/r/0o0rAUbpD4euIxZN4RDyHKDwqVDKlMwFHYnZPcSesWuAWtgI79k/VsGi
C5DYOtajuvDW2xaauyhwYPzvYOrIyn+vIpHCjFdi+1y3mai+LaHJn1TAOAKj
E8F7TUxWHHRfyldD9iJIej28YUxduj3oraap9LrBG52FOXgqq1Fl3qIsga2I
grFazHgjUqzyFu5WVvjJNq04OozgD4MflU8FYYcfCw1AMEaxL3578k7pFv7E
ugX8OawIeiF1RbTYFM0NJ1T1zsA8QoQxlCqGt7Io0daPEX36vo4w+JIbodb4
U5O+HT8T43BvXNcmhanmM7KYE0uHeljExwSNe3crbYGh4LHUqw6W2z7el9NJ
4aQBX5Bj2MFeaUVgI3N5cwHLOgggeDQJwkiPCgPMxyBcoii1v1EEugh38OvW
/vWDENU0ATtazVSXyN1z9U655JGddFpJClo2fForhIv+fxmAsuYpfChzVA7g
3ZfNdP4P1N7pLwoJPbB6/yWquP1BfRmmIxhny2JX6yYpjOX9ncfULU5sbMzH
LdVeneuRDUIbTztcXcoVzJweXjYfNsGlibc+Wx/8NYJyuwbrdneF1N+1fGXx
qvV16HlRM1NkAhA3GWu+o4Rht7anaohhP2idz26qBzLC258yPYDVJjEW8BQJ
NtoTf4t5p1LnYWqwmYkeSlfkjx8p7O1GCvmOBgQpM1ee7TCdocyFTdymD84b
/deVXByZQtp9MT27dGtfSlZsZ7sq/8/Kl0PyjFaXw7laRb2ox9E2AVEnT0zY
GVsiQ8ENmtBAr9vtB8AEnTV5BaYeS/TY/CZB4RP6H5k6XKY7GANNGYtyg6Uc
tlVLgDZVt55cX9mIbFw2VAPLjxf0u5IrzEN7a1oNktomfsz5AbaV4HwgoGuA
CTIx5fer/9uqq5zJSVptUNqIyHWCBFIfnPyPoAWguUXlpWBtvHpX4QuYYGNG
2GKHjnHfEJizM/EGWU42XVptay5Ve9q4hDG1AcMWzem2H2+TrCaUT/VKHgwd
H6tELGw7lNLN55A54n/TNoBzD/ShZjlK0tY3eS9KkwkFjHmzdBALpmOiN0Dp
npiDsMIZfVptZpdnyTIQg5aT/Gb9z+s7h1Ly4DbsL99OFWykBGkouFj00i6f
xDZoNwmAykSiN7gK97BGfmPkk13nlRm+kigzmfprLC2RhqdLBoUFP/v3glAh
oQWNagzxyE9o0Bj7Xk2YwUBe2nDXNxm+CyFAf0V89jX2vy8ib12kHp56M0zr
Z/nphmI2D97esQ3EEEgp+wAHalKWLwPwibxiwMFSw1QjxHkIPeX9uzggfAIP
NJ9FBtDWRw4h0DoHznKywVjlKdN60GVBI/h6eDF3G+28kJWppEfWfHlxq01A
YOQtIr07YlpIMy16vZgl7Gcum5eoOt4lp8oOmCHgQuf38BMqN0a8etNJX38z
tdLg55vgnXvAAfbiqEUOfjTapb66wmWh018H3dMECxIpyW2G9lAqtsZfx2U2
ziDyn48xk/cfzWhjJjH3AIQIE7gSDjEu6aQPSouwnyp+nBnwJPOp6fEwOCgk
oKpuhMDooATsXLUbJXHKJIGF8+qB0pUoFVlqUhIr5gM6fFtRMbhdFiGd8tAt
tcQnbEdhR2OiJlGXh/lzXrbh1WM1xRrhf2LIIgp9UyaR2kgv6bKQNL59MXWM
3hfMpBVbErwHRFIstNd7Dx/IqJoUXnxEBA+5dsESRglnJ9xNY0/dqQshZ/Ce
vL5E2F3yaILZ0gGvRIHI2zECXagUfbEzB2capaiKyUe05r4dbXsR+blTGr8B
vfftsW9lVJO3a2Y0v2MmoPykRw0v2/s0Na82Q+4TtIxVfc0+gXnGAvFezftP
E1HqRUJ70hE5wVwY5SR66zBqBasdZtEAk4MoZHrUCC0QFS0BgJP4VM0+TLab
w3thRCQ0XuSgT9NjkE5BTcQjAt7koh7Yc3LQ3Imha+ix27vCjkfMaa0PxQW7
gDnfS9bJ1MVA8GuB1HiPEwqTEV0P18nXNfB2QSxYpj2xTqfhAsTApCAN+a9i
2kwnWDZPcp7r+PzaMbdoJ7BcfWNRlnJ7jqmOwKyQF4pqBhUH3QCuDAXw8IFU
Shn2FqhPrrF5mgP0HHBvNEyk0JhJjZT+8Vw5oCVMalGR3DkqL/9iW11D+bNI
LrJmWdhuu2BJXeFM9ZWiMXq3PTY12IWKMhCEoCoFxbB+wjgn/c88gk6HeJyM
yb8hyVau+1SO86N5rOOKQpLILya9Z74bZOITErjGHVlnqioBga3x6BB1Urzr
WiNBaEbUZYXTI0PX4vIZPvCBDleTrmZ6rgrA7RWayNJBoppNrtRc1eB0RgcL
fEpe47Vu+fEcFN+r4F0d+w5xAcb9XmIbjatjzcqZS3EEQuM0VGXMIdGaqsAh
g3HLhnuyxOJGXJswF+8jsxDjHbq35TZwD4VG3n2WgQvzSyuwd8dWtlGVGgCE
ASkaDjdZhaWukOtvyT3xmiKWXA3yLXh29dr0rtAm9AiR8Eu//Iu0Ox1KZAme
ngy995FwiLL1HiQ32+2QZznJfQMJ2lb7R1MNFjO8V69QbKInCbmHesvaMwnA
RzDt6sPNng6T7EP1ECqjlexzYOfbxcu6Jt0xg2CQmu6oJpNjIsI7hUjnWYqK
Np/oJXt/y28UXOZbc3zCnDprQOFpTc/7H3ZBBHkUGyK7yevUGCTXhAXkvMAN
Yswne1q+E1KLeIoIpD6ImyvqxKkIFQ4WpecUoyiUYyFQApDJE21EkkekJENG
hNCyR9lKM3y3+5g9DjVSETDh/AMCrocabEuYJJ0V5CU/DdvgA917eFByAGPk
AEB71G49iYtZfH1hMmeTT3KoYCJ3U505l8y72HYcNdQZrrB763kADTIZ1QQu
tevyDEs4rxfuoPzKrSBCYwAg0KYs7/eI6OuYuhMdat+rC4krlALzeef9sB4v
lAXobAdkQVZh79XEbcymoMbt9KQ+BtquUlnP4/ii0GW03us2iW+/w9VhFIga
p/20FKocMtES8tXHdqy4+G2CYlLr7CR0DFQKDYEzGq5Jgybmr9n1LyJjlGZk
A1/lbI2WhE+/KEVU8xnMp+Q7eTNx9p/QGwNM6u7BeLSnvMH+iQTnIa/zuNs6
2VDa9tjDrC23qK8hdtMg7L/dO+atAR6QhEXt6A6V6J18jhVwL4M9m5cAIG+u
tb0doJPmaZt6OarS+0tIoO7tBJJPKR/nlbA+rOZRCTa9Zuw+RxVSm0/B6Zo/
WQQ1wiig3g1PeNX5efBjCgwlkZJeUKZlsqjngvxTB7kmiZqMVFW3dqaqraXt
Q1LaPnI5sKtUSlvPlU60yB6i9Supvi7HBp46Dqg65QRxb2ce+ZCkU24ypEA0
8qwTEM4sGCbkyuoQL+5QgrXb3mjGwbMJQ8jG1UEBd3z+s3hTrNWHoQQelsp3
DwNu6Rf+679Z+x4cM3YzbjBJfCo6SdNjlOX2DOSIDVZY7+YxIUlHjK3cUGmn
i6AFoo7reLo2kftBqpwgmzOuShksBUn6+fa/gAyaa4R7ATDrQj3TF6JgNY35
9c0UE1ylUf0rSLxSH8P7FrGj1SHsipEZTnwlucZJ4yH1JVT0RFuKxwhZC5eu
IZtC8GUBlGkG9gzXbVSS93J4d7Rma7TtsTuljdhs82sBqMsLGkFt1cw5PnXJ
Vg+Pl2N9vURtIGfdt/ulEDG7fJtElR4fx1gsSa0hkzhWBWvyMPpxwnPh6LyT
2GzpUSy0rZh7+ZO4HuZExztWbxZZSFXoSGR5mxyLY/jdBkM18nePwtO3huWq
wphcEkGt7PVRqOvk61uGOr+Z9N64nIyljqVRqixtwUSU/QNkd6Tu9kRGb0o/
8RAoDOOb1a3qNfkwTFlt+dUyGxAAmLcwvGtvPjYAWImvVV2VuD0Vud06UDOc
hZhsv+pnjSd5O3f9hW4GhSvy3M9Bf+FtpHuVRUSqFI4HYhDECiKrLMz8c2qZ
hujpxHDkVkal5fdHFnFKjwgUieQiSRZYLb8KWbwLwlWZBdmK7bMPmZiR0ras
lateSzc9Dvsm5WZw8bFaFWCw7LSRgy8FkpZjfx91qqhahSGGNchrga26FxjC
veCtpGKQYcs5DwYw8U3dmon4ZfNuljzjE4ZtOCm1cGOKDloqAhlBf7tPP0Qr
s6NzSHldMPTbzlHGw/PAE9kLHsw2kzzg2jWZrwdcuV+90ZxwqifxDP4kZhTU
H85OGJPuPNgd2lbo4JnCKXZg10VLFU+bXSOh/mHg6zfNUpD1fbZnIOExVmA2
A6LCgUdsKx3lKGaAPaiUR8QSlwgdzLpQhf2L9nk6fC/iuDbYhVxgKPwIv8lc
I7Sq7NJfChdH3k53F5/CakZiTJ43tOUDaVX8apDa44AvKjI6Cc0ghN204ipB
OISlOS9LbhmAuD92FkZR5dTwwRhOOXkXZkdPRza6pau5jPWB4mM/q0bN3MG1
yu1VbUHemTmhXCPQQ/2IuQsbTPfM4PBJFAg4LiapbeHilSBTejZF33+AR5Rj
Llx2lMNXHrwZ6JFEogL3m3AqWk9g86FvznlVtkecGQ9iffX2s41hIes0i9gd
yqnAJmUzxGJZrOBo2h4VELOY03peCiM03NV8kVH8bW1aNIG1gfjB0Es4Q/Ko
NJXUEUQJsAEqgK1xjCz3WAyXNJqgD58d+Jho77hvzHX/YS8fjhjD4s5KNFPz
XMQhaFdOxf01ktKoIuLMAaifxt5iS2grlxDOCc1RW4XZB+7/Pn7ZbV4mPtfJ
tgRhem89+rX0VqWLRQhaa5FWpSBS7giHZvWrZ+lgQqcSzikOi0FpH+NELGMA
ASVb+v7H3YjQr/NqojY0F7Iq9YFhEY8a1qwWTCVr035VbVMPomvmzJSWbdVw
5sSj9Ue//vXEGoX0ELDaW4TSSPtskUlLdIG4rVIqOpreDypRY4G/Or+vfoRu
xSLQZ5uHqSugF7JP4W7EOfJSiPzHDDauXRdBravE62bQFpdE67R7fPhMCFSt
DBWCgB31EJZV8WJVi/9YJ1N5UvWpJGF5ZRBUhUNg++qNXv703cfhBejzPyiS
gKtdsK7MXOmzpVKN6C9PAbvoW7Cn6En4i19pDnjTKKwn/Od1thg5he5m0dFS
7Jfvh4LOunu3shJ0pqBbUhBPny4OHR287X4CCfh3R7tlJ5KM0Z7ay9nu344a
sM/GbxIYGnrwcu0qnEdg3sFgA8BbTUj/RJ2tVyA0XBtTSVFE/r7HBaop6twH
KFimR4C76rTSfpzmYAPrs6wzXQUkYSOuTbXdZXlEHbqCKw6VYG1q92hF05kS
WAEYZNdtAbOm5315aE+ZgugzSTYmBPcbYn3avLA6c5krEM/UJWPdM9PWyI56
uy4g0s00WSwBUk0ahiff0jAnwo+uXp7r0CBF5Vt1twxHlKrndk+Jv6CVLWbO
CQOIzuPh2U/sVhVk2MOpTqEyfKNNkHGSs5ep0HoIaHmODXQm4agw/5bjHKx0
uTupdLRnB8LIgQuyxbpo8IbRDTsu480X90O9Gwb2Zkl7POsUqg1KTM9/LVLz
XALZFop7SOgUBBHPiji7Avc7LvGvStw4v95fe86gP3ymZf3Q7iL9TR0A+pJW
4bZ44cZ5R+SidHtGAk6m2zLs4GUrAzR8+XljSfOEDIs5niiSXS64ugKUXrT5
pTS5NT+ZJOswB/sA1votzat/olOE1FgqShVqngPFM+MHvdaZJ4zk+w9YZvO7
yKIE/CmasAuAwswbXr6roJGxis5XitXrsDRKFk/2B3aXNeJDAfYbJbGvGIjI
OhzZ0HfU4dSBRp78h5ml0WIBfeISmckwQio0Y0L/hfWx0Jtb6Fz2/dpYnb+E
pBx9Yz2tc9DP6rk9zbFL3utGW+ivuc/hrEgkJH/SqxLJ4Xrs+K4KerVgH/Bp
7o8OWAEPsee1wQdpBo/XhZQ3dWvhad/SR71q5VB+kJshBX9WEfsom3lEkCVW
51nFZxEQSkZvUHhGb+nO/0x1vNxhV6Z1nPFdB4a0P/XRdAWpY0Hr8MMtq7wx
Iavz9P8hoKmiAd2G6/Q+gB5UX0beA2IHSVcZvO/D55G6NWfdUmI3WKKLiUD9
A9ZrJ/JltzFSBJgwtl6gCzY9rxIhPXxJEW/nbbrkG2dBdb/Cuo0LzAKPKGOt
xLM7k3eApQAy4tWON3r5ncBz8Sn//XmcOQCqFcKJ+8GuGfhIRzB8MQxz7Fo2
IpOxMEIMwmoeoSV1y5pNk2pUw9afAQtOpdu/91OwAgVJoYqp0VhJHkWyHEVT
uy18ltLe2HE8QoGBBb4SYywFhYBoExlPHP1ButYCErnMsPhKlOSRNhrrilru
zGvIsrCJqdUXaPS4tuXyGNVmH26XpM6Hbdt3xRoleJGUO6Dz2Lih/aO8/g1M
In+iDoR+YXIpskNJPfmzKO6AnvhJiB9QvgiR1AswWToWeHaNlX++sclTiBWJ
4Zdx0dnZvA1d8ML8ol1k2iQ8yenCM13h0jSuDWtnxGDWPNd9TLrS9MAYq2rd
R1PnFUbcbvz9483NAhAflLaxmkpyyOjTlchyyNm+0V7ZOG5YWgqOmSsxFJC1
t8EvumZA7XgzmqChXZJ+M32DHlj2zYRzS30V+0w/g0H9W7ohVHXaJjxgLtUK
r4jDfbkT6DGMJ5AOLGSl43GnpmFdhtHv5+l1zQ1nwR5HgrZ57vEM8kC921Wh
KBirz0Pu/nt+Qud6qJC8QJ9d8n6LTRYXIVQ3KiA+ouSzyWZLFEx9/Ypvf3qS
3XNHIdgH1IDptcC4Pct3rjjmflobYfq/7kqt7P9aCqg1+EetxxxMl/twjemz
tPvL2a8gB60bRpG+0Jt9EK2PjSznsE5L2dkj0Hmbnh/3yWZZOiV+xl7HyEPS
befipkLIr08QoaqofyniDfvjxds+m6BbmFFFEjR5/OF5z1u/njNW+Yd002Rk
zb/XdQ1bGohQNb5qe09oW+WDShxXZMvKGB00mEXxXmC8vIciK3wbwCihi/30
WsrFhQQAV0T1utpJvDZPFEhRB+t9otjL8ILh2YYU1amyRzvyn6Wm7NpnFYFA
MFeq2uQWRAhw+pyTPGSHcDPz802O64xSfA+jnHk/7DoQaHuOzNKSr//Pgn8K
v3kJTXgw+nIsu84zygiM06JVbYdu/H+JVjyy0plIjX3aX0BcDvS0z5tVk04B
kCsboUCRPI9wLaDsNn5gfavoxQO4PyoDIDeH3sXhjYNJBJ4PHxMwCO73usrz
ySZeDrXzDNCrVn97pToz+NZBJdxysLh9jegEeic94QLPqf1+u/nJXRseZncH
KL9G4k9sD4bgZNJ5kSnd7vdkaYBD2OLnRx7NKpSBHn6e+tUvKDuKJD8psDbl
c1X0N4ERzRePEJmMxN4PCHP1r05QtcOkSEDv/CHbboqw/1qjGi0w0iculx9c
UL27GbruQl2kxA9dMV1tjbvUCo37zLf9IXjBwBF7kLzj5ufg4/MbgJxa9RR/
XhGFzOYKTaPr2Cyk569D3ChczqFnkd5nEiRgnXqb8IeDM9h54VdTr/Mt9gtr
NbiXeHAyN7ugyR2Yc5v0nG68wceXXjW3158Of4Gf5gbAgNqJS9GGyl/SISdf
QKTw0fH0jH9dZFmH8XZH5vMeV7b0w+rQq1XARqhCD/AsYFxf6e9/Eypet/xw
3ZwjsunkK07SFMpvkZXf8qgEpuncDOYj/Qnfi0zCPNTgT/cmPdW+9AVvy1CS
TFFfbXc22dFnJQ827y+L8RRB4voJk7j32A4CjOvI6Asn7tvM6Drq3te/KMkN
yk1ZlV48PrF9VnT43nN/gbkjCUMNdfVwO8rKSuT+UmCckzzOe3t/j0WWa7ni
pUNE1VFC1beauP1J25hkjlPClFznq0aP5xTSvf2hcrRYdaGPRfB+fRB2TqqB
ZA+A7Txp0XULaJsprll17AW8C4waGtDKtQlrhIDp2jfo1H+r1eigELWWg0kc
Fpnd9KxAZGF+75hl0Ycs42j0F4xmuFFuOFOg6hQ62NJ24ILZX5zzWshsfPON
+X0j85eczorSJaK4kS4QHhMnuFzoBDI1fvSA64VAfwZK7hpd/zPFXKPQzt5+
+WrdZPJcQ4BVeAwq4m7lFdcO4LFXlfe1MUqP8nmlfD1dDPaC16L71R8ZA/3Z
pg4T3Kd+hZnM8VAdBoCYa61EN2COxXax1lRFbjm/OGfNFvXAVsAvjQU/ShmJ
FW7puXfByBylyRwzFLFHs1PJ6iOWe9UGywlub44bvzwfeyM/X6wtGBrSP9T2
3pXOEBi+WrXN5+Y2fyqbISmfpIyajm61tKkKN4RiYgmEYyjWeDjln77gNl7B
xYXw7ux3wch3R1EIyQOKZPeXVLlp2TzAOQyzuktj60pCLOJRGdJyV9TVZZXQ
bkZ73uDSa2w8jkks/aMNeChaENshODW6zTCsWzqPBmUE3pMpRzuHuveubyIE
9n3blFwevF85iN8ZAFZz4FDHQSJFddFwOQSIWMXAo5iLiNrrA3sJXM1Q2BS9
DQTIfCtwB05Il+C/oEyrvh44ED2byZUAWeBruZHIaht71ZHAmzDQ8Ulk3UTL
PxcQ08tNikpgL26e0sTtx/g1C54N7bA3NeNgczBxwTUWULKv4+EAX54nEfU3
T3ZR/wgelV+d+oMLxtkULumvOJB/UqUdBrMW02GPviVjhCL6JeieWHABpMhF
itNYvOSKzc5cJwqClw3fNBMkhqPy4uu1JEWXFiqQdAsh1Ak254iCg7/SoFyD
ohSFAvbQpU09m/S8/zNu4hf9mJPq0VUWTshnIJ3CjGQMIYjI/F1tbtRcXIpS
qWUzPOnh6S6/kRbD9rVt4BDZ4qPKgKj2Nl8NCOCRQS/nt7WSl2H9K5qCUp+Q
ZDypk7E5kY2yTP3cJlqGyQA+oUFxB7q6RogmWHTHF6MGhfy5S//PsGULOuwl
J4Ys4kHer2u2vM5253lMzwK5RqJ90I2RyDeanYJ5ggc6N4kdF7xmLQ42n8jA
UCgNcWiGQE3XfznmU9vaYZbd7TNf2xdavLM1BukEsIP64rpd1P9VieWMcj5Q
2nieMCOGI5z2e/ROc/t33/j5wbTEzhLl2YwiLT9wYa7bYGZn/a89ZXZneqtM
96SSmUMp3L3lROQyI4KL5zCyiCNtJsU2w6AHRt2tBm7rtL4R33TfgVGZgt1G
OHPdB7Ws9qheMY9+VrAF0dGF1Luq+LZdd4OCVkcRDN+wKGweXidkhteSrf1w
K8HRrTZ3vPe9SbgfRVVLt0eRtkWS2eTK1iOv1wsNyshAV9pVWoHN+bHbACGx
kmKutWh/4tqWLT1/JwprrnG+aKbFU9hbU4trDvGMlS1mHxatmAVjOsGXr72H
85+c9PDGbaohg8W2iB/eA4go1utA4T2mEY1xrZpzITc7VDtG35Xo5/NxzLoZ
zxmMcbjq6ifXk9Sxf8oqc050f5n9/HGcPW2iGZ/tK6E/h8S71CIipd5P/1wo
ELi1PhbWUGlRJloSVINPEkVZKlzzodHe9s8c/GrOurccRrQnK7L30Fapaiy7
umfd/D3fFoVpf/hs4yDe0DuJzIXf05iNa+xngBf8BXqZ1lHGAKqgNLi/CDSK
lvO+CIu3SHUO3eyttKVrZ5n2PdU4cxzMJP8e/rIeN2c37IlikuRP6Jwd2oQz
o7HYvYHL11H9ieA2JM8RC7zexCX48p3KHY3fxB77N8eM6rGPBbaUyQlMcrMR
qSZKeii4lgfQlUMn0OcQMSPXRuz0e2cl6ZSbryUb3TGAKWOTBSpdKmjj67qh
nUnwgwBpbaQYYrhKF7tOan/QiYP9ghpIuUa/X4VpxnhxkmbHidfqq9bWFw0E
faF++P9IszQoaY7rUU0EECd7R54JEmJOnFzt8owGaOzk4zkEL/8EcvumKWuN
Ux1xkgK05UR7Wgy2IFlIe6qMxJuoYpUauKZDCvcIKyfBLL+ET3927FSh/44X
RDDepVSmkGXAg3Fvya1H3je+d7q9eEQRlYdkBX5VNTNGKhPKsu9QEk/EhAMq
0MrlCLBB+oW0ECvvoEuVyjqqTV7UiwotUUKcQzSugeLzLapANCPuNSdmqQ/G
8SRQjn+ZuWx6/9a8s4HbOTvqoyirGqrS/segC6oRvoMXQYaz5IXTNww+ioh9
OtLxwoSUVeKIE/ANdIG/AmtCDQ/SedI7bpYomqV6J3P9939oC7TefDqtoMP3
aOOZrndH2X07hsezz1jmSogghmaqSwDn7fIslUpsiGm/3j1EgQoUePSUPZog
KmKTU3vODmG3o4uVuvGZ2yiwqbDZfAFkKUWxnmxbTnmHyjk4pAy4k2K9bJXD
OAQ72EHmxC+Ao8OuqnsSuFcw2BJ7/Ll89aLLRlxU7z8BRiHQ6fTAXvLGZv/r
HclSZH2yvNyy231i+6jBQsO3B5zUf9RBit4ZszNBr2pNqy8dP0OTVvJ0SYrb
a2aA1sCJpOM5PLvqfIShL+H94IcSXVdiUykwaVykt50/GVd3xpBmVV3BcYiX
jjyb9V+Jp59VkgDoyxZBYSPON+3pCTYfsc9bdGb2hWBiNXZJ5FO94BXi+8g5
asX/oEQw45kE3JUYJPclMKoc1vXT9St8yDSHCx8yYM686mTjETIBApZwmKYe
6rv2pyGy5uKHdhHbwekRyLehoFr1bLRDaPbaHDFj5G5WA0FycFPKqAjiDITB
fxM28RhNZPLEzEsTMHydJIXy4f8QRAc9HX7ZdD1t59ZrN98DiMe6smOaNEBV
I7RE6VDL3FqmbGMgD/qSFauE6NbM2FWHfhzWyBeRVhoin+Q6QUETQb/0AieZ
rMsNeqpT6z6vbA5MHKStltLPS4yvtJPF8aL8RSX7AohRyqVKf1VEv5z9CNvr
0YQ4mmVP5jj0h7QLeJaSeANdTXO4P5pAHe7mEKhGfp7cJujecutRiwcY2HrE
d5OTussuCFF8/RW1txux5a5iYoWaOEkBfN1f83J0Gy4NFUJu17Kq3JsjaDsc
w9XLmK7eekJ70P96QKfWO0J2VU5CJ2FtM1ttx5nX/LuCRX24GO8t4lfbS069
yzj8/kD8ecnKQFct/uoiwL/lBsk5pJp/IFDvYXGa4xlZO1JhowNj4DwZ6Dfu
tJdekK+1UASm8kW2p2n8xs//4Xhzi9ezo/ylmuUN1FKov2cgMKgPfODzyN73
ZZjRgBDMdZc1ue3fNoBv5fijBDzc4VvWSyTzH2aTIx1IXAlJMWDY+NsLnee3
5Oy8nkmem1fP97nfFdrKffopwW+K1Mzb2pwjrdyjyjKhtB9tgJvWtVEO+pf4
io8uqwVInMnZiiw3iKujduTBhcxMQpM6aqOpFT2rgzEp9LWNbPeuF2MWHfQ9
M0OTg6sna0I7tFDmbMZDUZvZZWlCPUMs0md4dXu9zBbkNQi8OEBKqF/6i/v5
Ugbazf/xd1e150jkL4pbP+V0xBswe1CJry+NmouPqHvK5I8hdVBfI98tWz3F
SCvdxVAtZEihcqw6XScIdOsRWA+OP1A8bRUHFPy2l9fVpxEYa3a71WdfnDeT
GvOyMVH/T9T1lJlShjLdu/AZsbhUx3kziWAwyAEDZQYbNHmWsSvm7Eq39IBH
+8y/OLOKiqgckM02KYYMHqaN3GaweFf26nRntBKMaM2hJ+Xx3CvwxBtpm90G
3kKt0G3AKANKrYLuaaiMEyEewfqVl77OtjFNvBn3HmS3gGaEJGhhfeBS5+au
r3WXX9hxnOj0K3Mml7rRBG0mw1I07vEgwoXZpMnrCgJ7E+uQXGgrmU/5G5cg
/wDroYuHKEQVhBRjfycjVE0enwLcBxA7s5f3cDuOqxUZbxGDDCl1yzpsTMFO
n0KE3KThgEQGO9RVGW39k2ekIq4GECVzT2+wbw2Lhn2uPktvC7LCYOajLciu
lwXlQ9wbDpTnam8BpnnKAREfdPEsTVsuldeakQKjVZx5n0Obeq6aK/tj1lpv
twLChG6SbQ0nVZ6E5AOeLty1W4bWow79KUergGFaPsPzRF/cj4GQF5/KE1K+
Rug7HOUZmq8ZBqn3ZBCrGREeuqvNGdbekoStI33x8/jQ2eWGO05HZnHlfKSe
poM5nrQP+ZLPT775qgWfgUklcbW+oAKLm0ts72Ax7TxRMx82LR6BMFczRMui
WQGUWObxvuKmWNPxmxk/YBzWlbR2xHDjUE3bN/g1iA5B1VKAxm9jbYgZfgJF
f/YjxCJi3fY7vFZfpnc8OGSnoLqoMMNSZ0FejQtN3/h1WEoH/055xuO93xCt
wkaC5yD5uUe9p0oK8M5hdJJJxPxOD2XDvtjjKPjyUcfQZuLPCpaMQbtRjN+W
jXfC/Lhq2XND1yG812PcglmhFuvEzcIo6Lpdnf2o880IS0UfrcXu+ID7PDZM
f+LIU+mbnUOeF3D8Y8dyUx/2yaDohv9fvmoBExAUXt5VERPL+5CAkYaqCO6S
34aJKb9goIK0A7shNpVNyZPSyiPmJX1uvrT0M5IajgfVDBzcBp1uHt2sqL2L
U9reN/odXkDeb/Z68uxsMnyiw7M5yLSpJXWwVPT+pczMwCQkr0g9YvP2Z15Z
26Qd2sZ8+WKMIN2rIZZXBCMcYGGsxTW+JywyDrVOn4f6dA99jf7OhcOGLWui
NfBLGp6lg1d3aBCUAh2f/+dXBDnfbAie3qVLReo8z9lRZ8doCPCP1dTCfMdd
o2PaxWab/LVWHDTkgY1hDdwEhqmL5W7dv+7g9rCjnfwZx207TqLxUkeC6EWa
iuajk8BpAGSaZUwvhaQ1GVJhOwHdN38FkwxPF0dMVKepB4YH2tjdehLwJB+r
oIqUPlvrffjWaj8j0AT0CY+w5Jux7IRh2lj6brKYQyDAXekHfNKNJD1NTaOk
/ZfcZQZ3jwar58RWDANQDsyQ/EnEKYNhlNda8nOuVB3+1HcKjCWdXpyd8jfn
9FvGhw27N9abU5ec+67HTsYdiCi1ikzBTR0P83dyUJq6F+mAWA+kAgzZo9++
Lou1HTIFpZMG5n1EtyLUgpVxiaouxl6JgICz6kejIztcbaSO7E0/AT4Ak3Pa
KLtSDfrwkr/quS3XoCG+5e985RdXq3PVj3a0R7R86x5/rKPmk/ih1JCPGJFb
Ngs57WOu/BzkzitJBpUPXA2Tv8ABWKswdlonVzAukuC63Y92DgkpoyOyLiED
G2jNM4h0CGyUK/25sf6M3FdcbT0IOgccUxe+/PvjG5NOv3XlILd0aIjwKRyK
iSOeXr6cQvouNwHwxe9qD5hcuEp0sRYLNVl73grPzTxHaPzODrzufT/asw+9
gdKV2FPYqFfndMOdgxfKlWS3fFT2MKKnDr4KdOQGZOks7/V2KZjoMhcLzF8x
zPUK+22Uidt3epxchPAGhZ3PLVUcbXZUSgYYHyCfBraard4i9GXr/AUFLtP8
ny8h7EKa3mEw2ABEw0p/lZ74WQb1LbswGlHGtHpxjYD0w3gdqSka2Rfl2Yxe
gkAGoBFl9zNn6SVrTmH7mIPXHNytITkMG6Z+Bg74tx5ji5dGaPNGWLjjgUDW
f/qjawt8amBoEHGPyEKp/6nu1E8uwrwk1jYJ6/HjMwLSXAIEFJDgNtO/bRiO
Yl5dkKJdLtWptBjaUs3RHPqmIEWoLvp3mL8FOKpbD9SNJs9G68x0VIwTDhgX
msHQoc2ktJgbpolTa9xdPHdhtKxqq5JwzGjUA55MziFfb/88q1Ic0kQJp6MM
HIRmn/0G0LOcPZjaXZdDukFcaSjjC2GUayMqz/ersTgwAPIpr55QY/oEGYs+
q5zkGs6RDBkRyR6lWMkkWPJcV8BPz3pECiVtfs2rHyp0aqiyN4f2+c+wkQjA
pH3aGoY+uhSVQ0Y1lYZQs3rujnZxs7IeZqdotc507QqfklL2Ii+5Rc8jnWrQ
E68Nm/+9kv0D25TPQE6qsZFqE5IJcO7iI4QtqJLtiNcO1pwCxN7LKUeeJCXd
H3rxT8dmQaBxPPmBqSsXalnTarHIWSyeIdIEIV0rKDwe26snIs4W9exrbgRk
AaD/p9ykxIovBw4RM2jpoRYN5SbYlmllmJGDcQHTP3xjOz2zWznuULAmwpMx
vQ7WEvBBvwwWXB8tamYD7N7mOVkQvW/oZTO9vES5i1Mip6R5Eycs50IhvitJ
MEx0qBHmXpddlHS7l1wDpxQ1ht+Byv9VbvZOa0EH8xxWCulIVjKDZ7SaMCD8
W0U34XbEljEAnml0ed5Zse1BNTXTXX4IGllpYCzjqPHF+CaiIcYAner9lP7q
luzac2AnyGsZImW1EVpmt+ZpJNDFwV1CnC2LOZE+JxdyDImrIrS0vNLyWHRI
A3+52YqQj0F215EZ2JyVAqJNExMffHP35t846wADGBfTHTFWTe5sZM4JGdlB
RqILtDHadcNceDEip4mdfwzV4K1ud85YpiuCjXlMhswN2S442STyRZKcOq2N
V+EqXkyxptH2bJ0zr8QDfsRE69njjd4Xco2PhY40QVj8GB/dLH8Ldivq2NOy
s3OeZnKXb9F6ddpXhxii6ZEFraTQBPquxQ+S8HBOWTaQ7smFJAhAmWtlVa32
QNFX73LuPtw68kEHCP40Bls6F009vd09Dtq3iIi5RKtmgf+8GNEHpBmgTNn2
HKgy4SXjLSOLaQqK1KQVsyMMZVKAVpDkS549VVQqrqAik6Q8fdS/24w/FrQs
Y+jdwyvKcc846KyoZMHJO+K5rCu8c+AOqfkqPwNx6H3MLTMPvnPdXg0tCwzz
wrT/GTGRk3lRhOc0lvvtQsdjo8ZKKR2ks5/CmEbM2NzjK2TV2zzo0/WnIBMZ
OcpgMNobB6NhT9IQORfPm4zsxZOT7tLfF3hzHDySWH1pH/F3dynqmYIu+01I
/drYRK5hbus7wm0oXw/sUA+CBsElMPP6L2kE32gofHZa2YnoQIMqtCyjjFf7
eywm3PycERQUJ221LN3yZ/AxSSx5iG7nzkuzYiIimmhFEAUXP3df4dOSFlHg
v127It+Du5ZZ0a33MnexTnbwbz2dkrlkYu5ULCVTDNX1rUZqvFtTP0etuTB2
uEm+MWu9ik2wJqV8FGWp1K9QPI6R0FmHwERV6s2s3o48+WoYvqeVwj3gQhGk
tKEaI6xIieCdanpZIg4aEnfbdMqHLWBjZzsySspMA3dtal0mhytBJue71dJN
+N3Q4/7DH4qb4mkQ5kkaUgY857b64drkdbXt3460CbL01t5b6t9O0s76zCeo
vzXxjlYaDZWu53u4QS+H9neACyW6Cye13aZXayNcoBjgkEjIL4LfCXYA7eEH
zo8UHQ+P+8FeLI3BiBANQV/HAS6u7Glg5uxEqMu517WYfvnnKD6y/lBv1j+v
wU3I1FAtx6Gk+3CosnfFvdEGvY5R8sXMqMCvCZgP/+4MAjzMLex/KMmHxbc1
GfLtKxtGSkCmyRca/AcGRm1FrWyKFk4qoIkqpvZmMZ+ZrGfo7puYlpHsAzHk
PokoXxSQQEPeCj3oQkO9Jz92MItDG0KO/ltkbFu14zeVDtmWYfRZ+1MjflL8
thVqVFdAzqBYNOfVtvf1pN6kSIuOvzf5nXHW9jNw6vy13vFkBR+8y0Lq1k9A
qin5h5RspwaJo7S6FPAocIV0h92e6dyuWuIFVXKmCjFv1xj7qB4tvhw9RBI4
vWJpSVCmmKhau8SYuE0/KxyeBEaYJpMGmU5i/8ZzUL7Fb1ZwtVbh4z0KAX/Q
a+aJNN2uQ2hBKwN42681M6PQps7THxNLcHAlS0dGLODFylMjL8g/XbAAoMXu
s0gNaHE/mx0poFKh7067bRbngRpWai7snkCDFtha907x6AiR5TzxpPo8NKiy
4Wk5bgo5rgUOcnsbXeFpp/H+luWPcD9hfYktg6aHznvVM0A4uz5cdKTRo+T/
zEZ/8E+VU63wei6PHdh82YFmbRtlPJyqW083diTue7YthBs6ZgG6PZiGgkXb
9wmF+XO0rZXy6rP7EQK6gBKIIHi0hzWcwgtBoUJDddl25xvfyU8T3AQYusz0
knDlLTdiv7Att4tCe8lWVah41zCn+LI8OLlASXtmGQV/eySR/PHF7d1VL5AN
O8H/MWMl5CcpL70H6GInCq1RHU4zicYWoifNk8/LDfjaMSK3tvMi0/L5UowO
InnFxpFqf1KUQoeSXkK2zXlgSDmisbZpunwFEVed02esum9ZePQ/0wJ0Lj22
zuoNnLVTGdIHV7Y+9C9ZfVbPwEj5ERiaBsIKcCF0nxhW6uwQEwkJEOey3oDA
2blctYQB7+TeolET7wqnuANDb0cA4T5crPhT058Qo9gI0iUVsT0ILWuYCetO
J1VEij1fvEXqFkbjYLe9ytNgeThS2eoBaktBKSZrBJJdFFFjg3K4wGfcy2+r
dP6Fm0mcRzrOuixthXbIL+mJsMt67WJ4CWhQ4nzpvQUzn3+tqpiXuKqV+Gue
jZ+bw0UQcEb+5Yv/vCILaqPSTbhF++4RIiw5nlLa3j8+S3Jgtx4O7JP1L99p
93V7tr6a3+r5FWDvzajQYElHQGh7U0rgyiC/JgALqlm6zv6CmFmYJRXzgk3F
K+X5wj+JcU9vPHT7tNVo2wXJahbKGFjfpAAPWC4yal29X/C/mSntF8Gsk7Dt
ePAt1Ijiar+ylnyYPYgtrY8EyXdVmsQg3pr9G1aCZ2fVBl7iXkJnhsz1jKFv
aEsI1NdlEf7O6GeBd/pxtq/3btwUsI1XD6K6MFz9bLh+d3lmUC4kbRNcNS/v
6UVNyo4TVXFLiqkX/WVPtSbj6ccUPB3p05meTFdSTOudK04RC28zpja69Oxk
3zxVGxro6piOkZ3SQeOpnjJc9zGUzbumh4YfcZoWGjPjSt2aedLpVBi/ulM+
orx9Wwnp/32AEmCoM7x+qftIk6d8DXQtP5sWHWPzAJM3bG/X3Lt4sLrAcj3V
S1QTKjxf69H82N+UZizik0lifLVDupPuJlUDJCaOynjtqNDoWAF+tFu07hVk
qmWy4ptZgxlkOhvgdGmV+LtQdrKSnz5/lxsl7bd67dMX+MVvuYzOhxhgTIdJ
eXCKPm66c47kADWHVwSP9MgT5RiyOau6lXGuhl5jY6RI2Ii4Az0Owv3Y3RuT
/h4oo16sACF9xBX+FREbtHEVoXnPlxt3+hsxr/9YFF7d26zGG5MjrpL5jWVo
9eL9h2jrn4ifGIbo8v9X7wYEvAWbt7Qr5uJ107+2TLkegg6cb3j2OIKdVMBf
a5343FKFXQDtHPKR6jgANwIGg2QS9q52gzBVAZ5CEtk0tSVlitfYVIiOOGTe
cXVPNEfoxUg03pkDLpXSKJuHspf7CxE86sn60mwQFLugRrimhSCI+XVbMIeX
C0fDyMldcIMwxN/jfaUD9oYgWzcKBSdx4HVeta2+polhlg7NIjPBK/R/ABf+
07bj4LJKM8d1OvrbunLLFeH6GJzBQnlcmSIY9O/hl5Iyuk8P+jt3HVAE45eG
tAnScGGUQU5oiRVUm4+gFuZfOyl886uiL1VDk2oj758i4Ta9u1oR/q8LOvPb
1+hrwbINZG4UzDVTPixAYSNBz5OtDL48y0eEneHzEDF7gTIjhdgdhpxoPtsg
Ak5gqgat/j/EX3u5Xnuz3iHuf1rWh1285k0ycDMtLQoKOYJcm5j5/+ZUrVC1
XA4robqH3e7w2ef/HNBNSPK8lpXZ2QGqNPAKIzMYp46pjDYcer+qkxWZHWaV
DvjEQKFJQD6ceqVVasbmR6HhDtN2hCktMINi3+ekx/OCVQhz1DTkomMx4GCT
VR+vyojUJZcvduCnxEjC5l7Pune9A82UAmgtpSxjR+AUYiKIGc48WlJC792H
+ZEMRsj4/bqAffC4IrCYKrgqGvm2Va94FSSmM1FRt/5RvBL7hMKv56lHORqv
HKBPka54IG9GwQUp+8uAP6SmTx8qNKoLsoAGgyhmp3lGYfjeOysWkpZymKZW
HoP9quqGIYin4yvT7wydlg1cgSWyNWmWzmb/G+PHMRrQHuwJDPEpxoFVqpbN
Mtl3lF0/fqXwf1sWXSiCD++bMB5i3GP38NjrH+3HEYGdikgD0YKHeOtldq0l
F+u22Ly3aZIiqprYtQRjDjCz9Iw4hrHTX5T9h7nUhfCixPvhmZdePsg1Y1oJ
yEjyZdSqlkyvScyw5JFaxwuAuxIlx5Uv1tL6XQUxgrqG9KOBP5mBaq6lTfxr
iZ2yj3EaLzGy6rWufNmV853w1aK3kiLkDo0jnF0JhcJjKRDBki2W7wCcRrqg
+qK+mNirxplz3vhBAC+Gpwm6qTp8mvYXlWJ5qekn1fs9M+fYVeacl0OhBsWs
gYom5Q3wRNatFHO/tZLQuyX97/QJpL4s9vMZ+rDPFhhRobgDy5/dWT9+8Y4k
JoceVyUFF+IdnzQ/aYQ8wRn4ronm2LtWu5gIXO1Yu1IVNi9OQX+Y73IQG8xF
bC5Fn/9LD4ku/tSEt0QLtg+moNenfKA4u6dTdJaD7dLYdIeUlyQAmbl/dtTD
ysFP1T/i3IpuGM/8M4Ux5B8MBbvH08I24tPHEXCaqBtLBPKSDBD1hx7ERkzx
+ht7SXthz2oVCuncD0EI7zzxWAoIqyz71gV4xC+cKrhg2Fv8DiNQQfTb+GIt
5cI2TeljLaabfLfoQZDQg2kFFzjAwrbEOgM4SSsVhTBkTuW+BChqig99l3xT
dAnPRtumlcSIncbwXou01h0R9tp25JmrUfaQ+QTcAeQJ3Qn3WIH9IJl5jr2L
LuvNrSYb4NDTm+aZbhOP04B26hlC/tm0C5Et3kVppD2+uIy3Ut/KSMIPFVe4
yIk7k748v3Q0ieT94RwM/ADhmDWmvbXGMS/ru24x3++rAypILgZcHPannuaG
/WsqZnevmoIXbhLCwjncYZfe2UHbyk/uzR2JgNVVKsiCz8C7ujw30BTAo+Yj
966gADkJObS+UcvdfMlrD/vXEXJp8OhD6Y4SXJ3yh48ma1s5P1Lhfs16Gus+
e1aLPli3DQDYEznjCPPf2QvmemWR130B4xB7Tvs4V4XQPls85JTA8vXu3M83
g0iU7j/3s5QD0/uZ1GqwGuEtQf52jiC2h7zVk9GktbOnlmttGInn/28Tejv6
F4RP+gBh2XBtW21Ou5oi4sZO0D9rZduVRQIkFewuYxkF3SXbSaAKDnfBn8c3
9cnDulvOvgCJgXH0ojJa5wCu8dhjDLa1XUhBNPaoV+fCj5bqwjaSEsD91KV2
BG5KdQNPaYihFESRKl4Ylozch964jz8AngXtZNaM61NQKvzt+Y9zpMwM/iIQ
TgQgIkIc9c0YegjULTOgrqw10KWwU10n4Nu1fQd+9wBMGnEWo4tWa89/fdhi
Pp3IUmWJMCCARuucd7Ra35Zb8O9MmUH0If5woMcQb/5XrD8TC7QCeCNg1aOm
MvKtBWa6zaAzifXoxVj+XpeYhaF9mYQ9Hl6nqrfVuKAX3PEJtZj2onuvdG2I
2ZF7z5ZUeLVKxVteUmm+JZXcOgG/r9S774KGyHfiKEBuTU8CsfaGChZNBvB2
wLAAQ0dv66EP70ispVuzWfqhNAWdTU1qbGpHlKYgaJ+OVS+f/5zyPQ0OpK3e
zxgt9fLMtZ/ImXbw0sY6FYpiNbkNxHhuw4RMlApTWK0Ub633Cm9z+33Naqli
nZcBtZM+CNYJo7j8QMga+t5TljdJ5fPCUfrWhkF544jYZDHWh5+FXA/hU1fv
L6pdHOJv5Dg8Yt4d6NvVHQDcIfA+kotzW3UxZk6kJRzXWzFdUR/diGxx3qev
D+aYajWDVHU0JDDonLAmIj51OAcPLFg14UppNMoMP/LZsh5pTtq7ZtLNCST9
PTcEhOPxK7s29w2j2YLNfgcOlB8XJaWfclLJMVK68JUx4TwEjpQh6jf/Of/8
bFUxAp4o8oirSS3U79kl2pHIy+gyVYyH4t9A29ScLyZwXIhyONa4zJ/abarO
GwHAnbDstRFnxlrviMeb8YkCKVRSBjLtLvO1UPHyt6VuFEeGS3hy5Haue+dp
AJVaImhAW9EXzp+sO61ptU5AS5WFXFaszbB2aKrPLisNrbQjdQGp9jdl/Gst
R2trp/TA3S6z8Wo7YWl9biI+G0aCKsFSC5lhxKJjGKI/fT/OxI60566nhbfp
ymmLVCLYrW2CYuKdwsVAZDEA0m/jgJC+LJlkIE3vwIGs6GKsv+ENcSbiy6E4
5fCJNoQwC8vH/cyjI/db7evmJZ5L4nzNMG62f66/vqeLc55wjzq/jarrevdg
iCacSxhOMpwExllkqw/1I46Kskvw0+lZVcgFAxtwYff0gyPruk8UXyr9YbX9
rcAs4VbQlClXhJjk6jTfgPxL9C/QZ0huWX8qI39STvLpnAkWMtoefAIZhKsB
XYaHCY45CaYHJAUWpdDixtF4eAkGFQ1UmKey5RqWHiYTJ7DDRs92vjTOSu1C
r5gMBwKsIH4qRjSakA7yayxlSbUkfXOnR1HeMf3laRyjDuo34Ql26H03f3/3
eOQnC1KhjqypziV1sXWKeZNz28ONLPicTrEiFYZLfZDwOFu9tNHlMl+0Wq+G
mc0JOybkGBsFwXx9NbnOEXXenIkTMkMXEecly7L6CDQmCdqyfoOIaO76BTof
fdpy1l0s4tpGoAbsNoo/+UxeX2vYKZwZ1bSn6pkKpGe5U2xN42JWDSa+Pomv
p4S3YzuPEA/JNZqmfJV+gQD92gycTipwStHHl1lm9Vn1I3OqZZuFgrhwVMZr
W1fdQ8YGPtYy9FWKJILUBZVWTNlEuQ2E1se22vu/phqy3ozgTZVtCcw96ouM
rrDZcvQfX+PvoMi3FCifDQy6AqqGJ/7c2KVD4RdpWUWdg/hQMYh0Wfwxi9iV
TlFkYeYBub8BefsSuqmOEGzeMfwiZ9A4ayi9rZtFV3Er8E3z56yvWUnanoqn
y0OxOy8w3aXz9+bXdmudjEw6x9MBsX2r94WqkaHlfhoix5n0Gy92JABqVzHk
WDBw17Q73BjzhGcxxI6zRexiJrubc06E0AUi3O8JUNLv476nevF1jgPfCwo3
KPPC9qD+0pA0OZLJaixkze2vABZ6dToCEoXL3Eb13U2pG1h8HRm+wveSb1i+
Ap9KRYK26DrkVqU54k0j2bmfawZ1wfxM3O9p0iuyo11r3cw9tgvOekfXAY9o
oVgit6vgNOVSa2SPeP5r3pIiQjEYcilT9YLLSDM837vvj1YigdnRe51usf/Z
ADTrr8xfRwWQcL2T8hr2o6iUp10BwJnP657GWS/sZMDMeWjpsMZ0Gli0LdMy
y2PNkJeqD9H/T+gmmk3e8KNR+tIHznZ4dt8CJcgSzbpby36OeJxH3KeyJ6aU
HpyBg0MXhOMfLAyf7sJlQPRVwGRsp2J+LrJra4NgxDAmgLdntCGoCgtg0hyG
SBvffC3nFxCQZY76wBhDtwMdz5t7y4B9neBG+lJ0f9K3k34K33CVoHoq03ru
8jSmrmoFH05gHjfU0xJTZoT6JO2fBMEPqiM1Wi6VrZkPpCIS3nphDZKEWwk5
oeouCjovy7SUVyXGCHxzuCSmNgA8AHZbGek0wWzUcOqCpOuR6ZlYvv/2mj/5
gLqNG4WmvVlutGoDc0L6nfO8VfuCtkOxpO4PxIXgo69SnAt3CcriUTpqLONS
qfXoIjH6NtJQZx5mfAv9GkZALyaeqhsoftXVTz59HJ/YZNtBvgsrYzHyH/v7
3+ugVqQkWmVI/xw+tPApQOtJ+tH4VZjJQlKlIssPZotjJxBFWCiGU5PDu+3H
FxaFO5a6cWC5eP0s7R1VJwmdX+MMBcjJEkIbpGZwfGMbvQ8Tj4XUZg0EQ8hu
xPD6XP4tysVl+S4RVi9VZEOctdgTCyPuCfOxFTb/r+UowNlpwYvvS6TP2ccq
hcCKamarHzuqUHenG/0vS3Z1LB36nmsbS7ujIZgUN79NtzGdjvATrAOwzCD6
TETFVNfEZrp/Anui+Sx3jAADDP3PlBdu4dCaVTY7UA4vUctxUT5ZJ54BsGuo
ncsKi0+Eq580jecYNhOaQedUfVUmPwDjLYQDAoR8gICoX76WmlEM5hPd3GiN
s4tiTJlBjX2JZx2dRIfXFm34uHZZ2mNLmFR1Vbm0mMjZRL6+xwKtXpgkJrVq
KvHdGKq+geIFWrc1Z0vlwZ2wJTKClBtkfeh12WR8ED78oqhHzLFn1tAaOvQ5
NjFS1q3WXY8E4GgFjt/IWEKDbEfjRHD3zXAGYbfmVHPsAPdeFSRTr/COJV2I
Hyk5QleoGkvEkRFAkigABUBvQn4HB/CN9ht+elF40rQJNaYkzHh0sy7Ywyi9
b2VhasvZOLIWcMWkplk3RZh6sTmXoyNezIB6ohkGnfyrpO1b1nv0ZooAPKZy
pB7/w0rpVO3M9xLufacunM64gnbmyseZcaBJyUhaW7Wg83uxJZqoMholH13S
861NhGTHhlIxV57Lbc5MOUXlTXQuzePun16bTn0IvdyKjM3xVlBXX75isS39
coJAuAnZmzubEVteOE+L7/vsPxmQ4rk9Mk2+8fPVX/3JsJ6nAOdidYXzuRmI
5sWyemRo1R5WgZm2Bot+HOhITJHgRx4eK057NemA1lgXqv9rW1oS4BMnO9bO
y7ojw9mqH9rPKsou/T0Vf9iHhB1GrGl5M6gl2B3BerVzJv0NiSUq+bUmsb0E
rrTuUnvpixsD5wiQCpj6kAQBiD+nBrwBEhIR0eMVSpRlw2vHXbanYV3c3Ir5
28jeKeudvD0Ns5+ecKpq7wUU7H6fVblARIfuS2yyddaGVG9jw7kohoODOkVf
qgOkGSuHWMWtttX83NcEFCE4c9mD9AbHdwxsxcnubKyP1h/WBdiNHK+BdKzF
6VvmK1l4TEmnD8fxRjfJVbmzmSrl/YHzngZ0rNaV2j4PGneTN56Z+KjAphQI
5qE0QNb78cjUKGikvdsV0R36eTkolQHXsV+GW4qMhSprKi6h5mcnIUV/wW/L
fADB6EZOxEzlD7Cuz2Ue5aGgzzgdENn92QbkyS/j0YKM2NLIdesC9gvKNTHC
7LEdEqY4EXiKYjxhZy5Hgn0EImpWxxnplibzIvYLb+pHHtqendVzUbfFMc6e
WZYtob7gaPoe19g7V3DtNsGX+kf46KhKJLm62gax/aJN8Zwz+bdKV8pRpDos
V0P8QZHRhclxMcHft1H+lvxcWW6l1TNxT6VARJ3tyZj8LyEws8MSc6i+apFx
m0YakW6Q7artatN4GB2J5M1+j/FxueJP2s1eOyaIscOJfXiBGFPLfuLt3DmP
ddXZho5JzWYUk+5Gbg/iWHp3hpoTtykcIJQr+5XmiFeuEvme58Sbn/q4QnBW
Yz22bA0HQfCFWzmf6fcwYgahmFuK0VUaAjC5C3CqZyaH17ez8exurCxXUhQs
2Nc1P5IazZ/bWrwRVY12PDt+YVrH93MThmgosfUfFLHnc9VpCOXepZjD36xd
oSfr0gOALEp4L7CJxMmfI6hszEALrOxt/OJHW9SAhB73lU43XZNEULkBbwUu
Of9BLvTX3vc+5roPIqjPD6EbiZjws6HRJz4sjkUh2fLYpm18XLjs8Nze2lHP
8bf17sLjALaXczCD5tPMMcYxJzZz+DHx7uQUSNmqQO1BQ1UAXzoy8Lrv4OOP
WRwPsYsPzbj1bo5Z35mEyNuomC8GDedX5+fpQrUM+fazIn8/5TmeFaAo7zoo
OXymfu0VBL2hVqMcDeKYcgU8i/c2Atf8wthMb7r5d8rp1bnj6jbXcs6Xx2cH
l5zfvXelewzC7i8iEckvRQlxeZ599yVVyPRFwVusXzSwBhOz+zsHaZ0nkWs0
j7H0oD+KA813ptPoT5ZprkW71ZidtfeNUoF+9WYYaFimP5cRuWqNW43R0iXc
AT+Y0LyypMdv7fWq3GR+E8bvh/8tviOv1M1iZiby1r6EBGWFY0V3Xx1PybVF
DwWJAvbKk4jlu9ox3+vriPpXCA/u/BEG/9P1C+E5L/BEtbHhAVMwciUiPm8B
BRRO+YdjWCbhuy9v/IOn8/u9JadDlbQgc643d4FH8ocssg9O/MM+lKrnfgig
SUz4jN8QgZOVBzhdztxDpwmsuBO2UmXhC4+xtCno9Aq57jIhvAD+uGcdOxds
o4x/JiHInaUAGU5u6IB8l5vsomgahNtpC2PhTaYWm9xfT1zP+MT21PaPxRu+
rYUVOVM6eRB4FdNd0jFsAE6F4/NGIuv1Y74lcmL4etigBvCLze5ook635kDw
Mlk7SrM7wPhWRXhcIio0cKiHuETHJcyaiKSSTX4xv3BiN76qJhnxE/Ls24O7
PlevmNAYgc5Drcbdenn75FKErMoAMSd9OFY2O0cttfOhrktPitGZRQikFckU
8Si3QeRVTq3CScoLGoqoRE3lpYhoZqWdJH/pe87mFW0j3U9aJF1d94M5l4Sa
32Smuq8b5gGkFDxNiSWYVht2GeMFPeHevnQ6ComNl3jF4zZ7iiBPj2JVmaR9
odSmY6d8g2MRPEmSnRNamMq5rrpuzou4Wd+jqHu5s5P6lnPk2RhU/DM77dI5
LCB57+FzdPoc0bGxlOj6NZFNsVY4mPzC/hNSxG90EmDCIsNaKpYZ1yy3MWzC
rwjKvQ39YVYkrbr7+VwyMCxsmHbqD5jEaoeUJgoDuoHc22WX6RxKS5OsL4da
SOmFH3tWkCtKUob7B+dEuwo53un741flVosLO725GAOfoy8QXQtcvdvqCxml
mmgfNglsf9W+hU0BYidBHPy3TtKZIKIEFptwqQNZ1NqiPYB2BqHqFNm1YhSC
qu6LfgB0Sz6b9xAZTw2eu7sSprbOsOWTmQLiLELsd3o5QWmYRhrSI8W+alX0
UgsWYWqPxqRNaEONu/KjnoO2T4LT+ifUY7TXJ5UPp/6320PgYIwdHyoHQ3U6
z7FGEljUgFowoS/vXv4ybYby3b1E6/wV31uyLEKYtx+kT2RdgG4L9Il5PSmv
ktBgEyrwY1uC+bx8iDyMSI2SrCbO+e4M6HrIoMwloXxxn5cI85GvsXF5oYaj
hGD55jGpycs1L7cHlCgV5fUx+SZ+88eo9jHjwGm1BNum6w/OFEm5uSCuA3HA
heLFVp94Shifu4u8LHLGvo9pphefN6o332g6aFpQ0CP+lyUhrsMaZ6mcJOAh
qoqA6Tu2q6pBTSQ7tMSsxY2/Hyd4D0rzAa8joGFSKXWkarlg33s2h9/RjG4N
Vwyqv7HrJMdlPzx9MTL5DpdFKBpAFMbFnsRSiZ3vMXevNmlSnd48pdTqHiLd
wG0S367BWCvYtYM2RoR2whjfMibHlhMXgijClmKnHLtp7QzYzi2nh1m/bqe/
kFW+g/9mR8utE4NRGi8zvlG5bGIO03DmGnFEzjsnw4N5AZsogg5OQVe/wwZ1
tOo0/AU12qSBoIVdq8wP2uriMZ2l42O3RUN5Vm/sPKx2cSfaT/lLt2INwK0W
DvLvBcpPSObVuzUkRUK8NSlltbtgZmqYboow8RkK4WXhqBWMNLfJbkjQ37+j
ow6GCHuHMoe0Gvvu48mc9Pa5sSiHLRwpNWKjwb9jix8lplfvhaxxi7YUwM4j
2dMq0R/BkpH9xQecv43IJt+AU75Cbvy61rbh86UMMaub7lvJTMbt44inlQnY
zwAlKIIJIxJrCqhp2H383a6fMLTIGzrU/qGuDF7u1+7dCIavh+kSLPL8CCju
CnItNkDU3WFbtg7+Xsd+S2zjimjHFTQVp2FjpZHV8Tn3DHTYMf2kUuoTn0wl
6fI1FUQmaDS+YdrpqeAgvUdM6uAcsTX1wD6JpYyNRHRMy/hWUa6ZrpQKXyN/
meTTpc05KeyuL8mjtVdmOADDyYkVT7Q/tBSjJeqGOicfz0XRFvkHdO48D5vJ
/vhuht0nk1maYZA/ah4f5es/vA4SPXpkNaOg8fQW3pB0unURz1iofmbOFbSw
vFnPvdpJiwPSe2RXvDcufu9FyhfsbUP2xRyFXmt+0e2vqQlH3Cx7BP0xBkwd
I4XL+Ig2zFfIn5nIvy9kJvRhho9OwUu+Km1NZmOR2DsetLvCbD1IV36Q7y0x
IkBTzOlscYhnCi5/xGdDe6ezQZyqrp3K2tklVbzpOeu0pflrnxXCVlnFzEAB
jAiM4P1afJ0YhavadxWqpp5rugjiV0ZQgsqbLapnFFnXLuSxPXzDlo/Teck4
Z4P9ytk2KSa8n+hnYOci1+StpFu8tGtn7XwRooR93K+qVCdoFsiHPRUQ5W8m
RueMxKDClt5jmYl+xuw5YpoS+gkG3OqKVpvN1cYe8IWS+h3kXaVHAnoYmrcd
m4VwdLPQSsMWGvpjj1jq2su9QcaqEEs6BZFpMxsy6NhiKm9mQxQHHW+/Ft0k
Qwi1tdeKcG0NEOCvbAmvIRF14rPYbP9PbMGkrINfM/Pqqb7wBgGHJm6oMPAY
axutDB90X9GQ9B4SSl0wLBnYmsNmYyhYf/6Qebx50GwSJNaABZ7eWpqokb8Q
3nGTBPGGhybwVR6w8CSu9mysW1UeTlhMqE5BvBHsu9Uo9691annBwv6D3MuG
2RtIivM+eJ/3PT2wswsb2bEYM/GwMWhAoVRfUuMR4GM+cZQB3Rhqk87aeP7q
qhNi7PPMyKNyab5f05cQYY/mhWZrswQBkXKhozz12fubMZdvMxKgG2k9Ksy7
FKdC/JKOs7B+7ph94JU+NCiTp/dka8U4GNdSV/W1eW8YFWPL1nn3nzDIw3PS
CY1mtdPgxCkJR4VDdZe8KpNp93pkDyfMkulHOT4709TSA9IGRQCYM7EQfuJo
7kFMqLGGOFqock68preo/kt+v46lPH6sM1uy/nY3xN5PVNcgVQUTMPtYktqG
nRXZI5k0zaCzDmgdzesdDOvq9JbuafHGRWlQ+CDWjCKLRr6vqoo+9FBHPLT2
MDVdeLSyZhxJ+wKAWdqj3YlOfkqIBNJ9ffjO26cBVGN36ghHtNRoSG0R12Fz
fTy8noFxSPm644yygCrykxT89cOwxf68gMfB1Lj00XM811AJpbQTyI3Ed1a2
UdDNFgGMXxHjXbzdidB62XceXFbb+38zkbRKLU1FbDwft24GmupCuqV+x+VQ
/UzQWtzMZD7U67DOWORnN0BFMfjv3SbV4O28XgzHVtnJDXohwm94A5a7GV9u
hRFedqXzIhlIBH8cMiD4ltRdOnfggmKeELmcxeq0VdP4rDSJxZPzzVoA9J7T
Pag/aokS55OKmYmT1KHq0+wOZd97LyeAZ8tI0zBUdce7/aXSGDynMMRfIX8r
LzSOMpuJuntoe69aKynQlgRBWFFptDqq0iqy/Ucs3i87MCX7hy5hICyQKItM
j/USo8r/vvZAZqtHH6uRAGDCYq9A6sHo5iLd+xhOZunnNTqBoIjiX1sHx4tN
I+R8z6hDz77L0NUYUdSyzCbLC8MT0LRyYPJdbaQxj/YgRT/tOk0uvuDi7XCg
ISSih8UWDr1LoE7GukOU9Bg7nltnxs/xHr7VbSHNb5Wz5cia2o2Fgz/zIC+u
0+L4EH1OLevRLHBSagySB7B40QVg46mj12otmAg/4ufzE8wiA1moB5c5yaF8
CBWLwkPSmT9RY8uxe9cc3jWFizk4YxBz7JnoFXsXXVC99OnXuCRCGb5wB0w+
FDBPj5bIjnt5do4VqYrM0spnuBR12nV9YsLjAqPSYwf0qo2+WAsAAX0/YhNs
JHwnrB7eCtIIZBkYzOh9WxXceEFZyaczox69xp1ytTBQolS7fUuBoodCeFPi
+Nk7p2KIRPgA4skSZaGKIHF+G6/AApD2lamLCK4C36BczUcxP4f/0cmDCaDs
Sq7trfx5sJwUAuk45CmGneeUqkBGFY7wIwkwhtiZzxNliuG8Qz9t2x4ZZ3ps
8vjew2CX8p9gQsA7lOPCq+AB/0VFe38s2ye5nb2zFB5pq7DhTsqCgVfkwoON
Dfojbuzam2wDaxIgPdJ/tm1hv2oSL9AfIlTmdbZ+wfE4deyLrgqaEpF0UOd7
jLtUkaQQyMSZMgnc4NlLP5TX+7YWKHbmwjF/Lcc71GlUAyGOYsCMSKadrkh6
XHLEKUDlTT4S5lfum6ZzuVSj4HtMhVTGbI1FIo7hdXy5vFJ8Zne27bCfZ3Gt
p30P7ygR4njTM0HxfAVIbdEVb4HfsIPkY/DjFa8AqQQl2vPU82jItWc6YJLG
vi/XadD6W4PkE2vw195c/7w9wrIHoJgrI/QHGBuJt77HuW6CSy0xk+mCgMQp
f3uf39B1ARxBoz91wqr0CrnIK85Pis4YpoC+UG5PM2n4wAybzOnjW+Z0Fc5U
qfuOuc9Ln21rZvLGgYXbJnV9E2QD/itm873q/fIcfQdKKggn2CVbAPIy06aa
+EaNQ1GZ+xIUd4Wl0jnC5c23Yy9UbZ5W1kllUZST0G4Atiyddl942Zas0UvU
Skj2H1u6xcIyb1Ku1Y3/AL3Ehpw80lnvESQbrOA5QQ94TCA/+2YDANNn2ob9
n5owoo8xYZ4nkZqk19OA7ss7imltd+N1OS6GpX9n1zgWnowADn2kd+lCjxF5
PcaOvDd+jEQtcuNaBO3vWpxR3AhWNa7jDfmFh/TMc92xgfMLbHxEnwrjera+
CcEgk1uYGf50wIb6/XXEE7NLuXttrWKSLAKoS1YuAb0P39DWKlGCSI3aPIvM
SEseLBLOsriVi1Rag0cPxRKzTydXsixbUa754wJQwQTgXQlNxXz9UQ4kenyI
hdXhTBCdRUiZkW9OjZ0fKRLjOfEj9BkmqAUtwRMuxVSqnomX6Bku02OpOX9s
vNtAAXAOXEyc1HkiISzAAyLE07FbVHkyUmUfCcbepPvITJZnHobY0wiwl6wt
hnadDZ65ObrqvZvgJacYMO3A/GGu2c6zZGxt+aL974EWBF12oQK82n6+qXt5
ua5C6pLTWgFT8oIV+jQpodXLTGEWY9IHuPiwrUjIer337/iTiSWf2htGCFIJ
bLW2nI2cyS8woYv4G6MtnwyxznN2G/6ZpUi5fEAQXLJDAUPNS7+EI8zSrfX2
2nokDv7Db0ItEHHd3CZhns3NtthP2TDnVLMpyOyiJbG9IRAsHesn/XbxdbhJ
1If3n1v6UqiyfUD4JXL5ZDd/f2py1iHPRSAHPSSRKbT3INjWxzcQGm2AyXeA
uraDKFCAMymaeIr3a/TywACtUTYs1Bi28nfkUc8SDGYEanGg+1NicUw3bpq3
cvs5lOGRTnLhpNOc/qdxsX0WasxBYU/p9HTlIC/vbzv7Te5ckV10jf7C4t0W
o+/m0NFGvcyvGUmGAAdb18AgGpv4hmk1lXfXocHcVMebHbBxKTpMG+wqPlCS
1LjA23WfOn7xSEykIDVFbGR+bKupf/GJkZBwRoxSZfCAZp11E5hz9DmNbEb9
dMWJyza6yQEc+A7AKiN53r68IrxJgAGB3dMeSKg5rfVEs91Mu+ivV5PIytMq
0NDn2XcSYICUCU18LZWeWZh83K2zjZ7NMuCwY2jHLx1BqWn0GnGanMtQgeBh
+g6wOrvIhQdla2xU7LeDNBjlhzosgDThCQZgCVVRBu/t+tUbvat3ViKVka6n
g2eK6e+n9B3MmgKOXtLixxlJmCPT4Bl6rX6Mp1WKG2NE/NnvAIm6eDWWTaPV
iwZTDrBMBhgF6738ExSQ86Ig0M0+N/bPbwwwhH6iZpg1kabrrzXEXX99Bdfx
a7gkvtUXUhh8YIgcr0ONZCarGmYtelTcL/vLi1QmlJZePlsdl9l4JN3PsgIp
PVue1/I7IIiFXJj7GM0/OGyTwaJFb0VMvZkEBtQ3OJ0cGJG+g8BaNV0jylCz
WLoBaNrn9ZvTirFEJx8U+TK4ucLeQkfjpFdK5Qso2SwPguCALyo7TaWlxLSd
4u2KazJik9zrDIaotUaw5OHz7cbbWArnzXy916YsqRqrbYo/uDl0zsqibarV
SAfk/n5/kq5jFyh3Gr/TlWZyASFEGMVMKC3eMEsJfoDyTUdU5MzaniJc0/xo
EgD+xRS4+pc5AGi7lH/hjt7DPmliInyjzGTRolEPQY8LX59f+I3HQzBXRy+N
lh9DAY+5XgIB0RnguevYAIsnTexy2fb8p89c3O6XhO3K7zYmtuUgUnlVmy27
pN/SnJfxyuqbnsETeGUXTm2kuCwnTwJRiAwxOmGJE0DmThi87H1bYmsaMOQz
Hyh+Hb5aTHQDuOzzIS/pWmxCnv4Lg5uwCyX/dVGcDzJY4WdtDpyR6Crez/dr
MmyWOJtSoBwhbz/0CvewdZ9N59azsIzzTez4GGx22Ce8OUXPNr5r8v+yA335
ZQiCGKLNxvLuI27qZF+MDNMS7qXICbU6iU4/tmzP24Wl7+hVxmnGx7SkkKHH
A1GJmlcKwDfDj9+qsjNbtKYgoNNnmzUw3nj3SjtKk8lQV6ov2wZBehy6Mb3F
yi2Zm2hayYLWOBw4OF+aqm0fnzY2U69Q/YSd7y+fOo3I24ufCEhx51e1J5Qz
pjxrJtoZQSHaeZkPPYzUAbfBCX+VOZBQK5T0ZWO9yJzBnqMv8h3tGJ8OZxUp
dTms61m1Py2YAIyQZ75G/LePg7Jl1Jb51NWk1XWpdpqnAyHRaqw0ZJnra+Dl
osAn/aZcFzkq4VyOtbw0/ScY+qf62kXAa/nI0hNKka3qRuWT/043ZfyCTj8T
aHd+uM0UoamlFWikKryquZqOIZoAiIYmRHC1OV2YP5VhPt8rIC0ovGUCFfZc
BiBXv1WoYnM1BvTG8DCpZd9I99W2UvAN2hhZSiX0ddeZ7MoE0Sbhp1LJR9tk
eLeMv0jM1DBNKcvE12vDvpwbM+yJfsyCRTYprZGW9AihAYXs41+3Hhes/eBF
KYr7TxICGiIIa8bkveF1KMW3zre2W/Vc4jjwmRLK4EgRxzlI/iMjs4Ma70yy
xd1huak0u5S6m5jgAdw7fgi9xZGUOPI1DubXxdgTLU1AZw5fD75pvhc6RKVI
wHJW3LgVbJKyV+Mqz1XTvNPMmBXHq97oSRzOkdFAkaI4GG1RcVv8QiB7g0Sn
YVw3JWMixPPiLifHAW7PMMeMCbRIyCkK57W09f/Xhl5GtReDMmdagDPC3C9S
btDaRkbeZkByb6chB4cAiwAwmHu59WU2uIgsGEX28DyTZXA1gClG/ZelAZUw
0a0V1PGzsHcMIYGaUAXE5Pqz05/gFLkyIwAJKo0WEdEuMNfWAcbkeBJXLNg4
zccWHHPn+WiSPOAm6OLNrmNsT4SMZDi+bPQm2eQP2LSgX7wy+MA3t0fd9dtR
ZAb5ToQGjbdk4BHlY91dltMwmIM2KK36UtHLT5r3vNYkqWUoAZfBzIfs+zov
3XpYHVj2WjKWOuHodJUT8tbbcND+7qODiVJ5lSS3tcPZgGHFbHZWL62egp7U
orO3QC1AZ/saXW7E1962MN1rHl/EEVY70A6Ni5lhJSNQUV5MUeUCb7IWwSmR
MEUBwgribuNwCHJ6yTHReiK4zN08VmkupN2Dyc+LTLgm9LhopslmHhSdDweY
3nfnkumWm2h7XY/9no5ZFYUzQdJsFEKFUoWcvmxbhLB/NkZpV3Ll8yXGp1FN
d4scp24hS9lprXOhPz1yF3qAM6EWhsw4bPdsklezoZN8q/xk4J5aBlez4+7h
HXoSl7T6TzJw93stFyfC58VMG/B6/0LAZEGKVQGb8XsclT2THqhyQmujEEoj
P3L34cdEp9sBpMKZvaB7KBrHs3GF8G3yivsiCyqM7JDz+0rhtT2C7IynMU/p
rE68CipARjiYcnPLo/+EYvE63Hp1I9HTzBIs+PIMq8PPc3OtZYSRiTU7Wu5H
GxXm5hLbc+QefGOZKxPlNV7mJ0qSDyw3zVtN0yYlohJmJvByMzAOO3z5qQiR
qUE9SzGK/TLnYdUW61BdxLtlxSDxVgTgcWBBPyZ/YetS2zkwB/gFy5Twnf0P
f/ie/13lnkgMc33c5ISrawbK4yd6LwCtppEqA2QtJ5ws25/fwfrDuHtNC24N
xcq8PcgzYHcN4AqqjMFXtL1chNnTV93NXEAJp74Rl4Te3eR7Hf/dBbZQ1Q1G
NEaK6Pjw6PRnMGDn0KlxyYUZqSsZZFfjt5/F+tq44WqYVJicmpFrCCkafEII
qgIlIhQTmfFGyuA9zQdjUPs9uUY97/7zeV0IKsMXonZwgpqZULqLNPIfW0E7
lPHtbcmIXSxpnne09M6lF+gniZZEkyJZIz3HtE4kq0idhFO9hPwHIKrJw3v8
WTSdaUKqrhHkYe9ccOgnOlMNdUpinF/239jd4ngPxpncJA12ZLC9YIxFj3tO
EVfyl6DXn5e/Wh8U6cy275cTnb2EJm/Ewi+SDMRWrRr8h58AzQRcwQE5AdV3
p46mXgleaJSioYuOZWPB4xq7v9uGY6qYPWFfyQ4CdKaclOearMcl+lgkZy8s
SCGDU92yb6YbKW4dS08k6d7In8IQ3TXQWYM+anJv8DFAWGxhC2Bs1QrPW/ay
hmIbFAVLE2Gw4JMw+8paZQzgbXbh8/rCi4xT4+tBuVzTu8TNlevK+YJPB17u
w44VTDZOcUtu5owV5F0dJux+h7ta4B6nc0kZPckYcU4mbDEk4nQka2DLpU/Q
nJfYE9EcQUHeKuAmyIjhgWue2VJBSoq5nZr7Ptw44993t/MdBNbBzuodZwC0
zOko6qTkbMSJum/6/GFVXJ1Nez9gS5rjlPLR0K3qLUm4BPixY1r8WX8F3fYt
pdGzBcwVL5BQFRNFgW0eSlAoA8p05Ux3HJHn+hIKX0ef/QuP6ox4BA9iC2no
m5oD+l38gKINrW3a6adDfKeJD5jMIPyFwPnUeDQfz/jM0Xrxflu8RgBi3BYM
ZGKUAfoP4rdVyAMACBIGi6bOzI0P0yrtk6Uzr3OtD2HSzr+ct8m0opM0Ioqi
/2aegjP08GnzfGN6p7bWIUsPVbuVfG6OmUZeSdcamI3d9auB1wUylczzfzHl
sDhmt08AJo6vkqAGT+9j9qzhh+IZcVZtI3+LQu/th2UI6sid6ynoXSPf7P0m
dOZ+vuOzET5duZlsRWUNhEep8uWJ18yp+LfQduL84ERnsVV/8YQAcX0kOS+7
eAf/Bq4IqwFB1isQGGoM77x7W3Yhb1jwcvB3Yz50x6aA3cK8Vk2uGd7guX0a
5UyYfgQ0cHdVw3na1lBPCQezHUzQm1NzDTRlCvub0VRpi8jhhxeltG6SjGIA
BmvocVBu982v8/+xA1XiFt3fZVA+gq80Q2u1sNw7+yzExM/J/jVI5Y+aSZ5n
fldUf0Xwueey8AeO6IuEe8egNCFSSX/lurlGVimjNTG3eBbMpgV7qev00Dz4
0Yxa/S1ke12+j7HUQnJruuW7t2asPRfPtvzUrYAHaz7F5zZkD+1wo30fu9d6
xgtqlf5/YQQ1qbDfFBCBad0cqZLKg4cNC9bPiT7vp5F8iC0wT8yDVkcynKgZ
2nS5K4jhvg3QmYEo/qjzEvQAfGHFmJrDr78nNxLmyWi/yvQvHUz7XNrP4jtu
8f/Mver/OWYYFBv2tHTpeplUgfdZ3HbtyjrIJvDCJWTBksb5Jugm/X3Zd7rp
JQ06WXFrEo/yebiQ0CddjI/lpk0f491rD9dhDk0GygggDBbFkxyZTWzWHXXy
gGalpAVgTC8Ble9SwKKiiLke+Ifsu5LR8sINwbd+fYQtmppnwXBUtgPSebE2
dtVvg7CvoTzot1g+DA1qdPfuqXRJ5PKMEQWg0NVyrshMrUCcCOqa6ojbcds3
rs4NUC66/plFENj9eOD8SpJImZJoYyiJi0X1oWQne0YmuxGijVBUkg6Q8HR8
aDEJMKk+Jb/gHffJW2u/ktZwgDeqFdTDKSykEVdakSIqrKxMzjjl8tn+K/kJ
/IeGCAP00U9Y8sKWEn0+UvhPJ9N49Ehjj+Y8hK89s7vfXlycOWDIVdpG5N98
TA1edmcnY/jT8asq4qTTWkoapNjr5yschqUNykNvA7pCy4qa9Zk5FxbfaBLa
yogU/bhcyocco4vWrIjlaRMZYMsS4OB7MEkiws+0AKlry7C0bkYwF6woQtRw
hYF8U5y8PUPkO/Il7ErvYDw/yAsMRcJScf24pN7q4QPZuQ3qAR6zjmX5x/Og
h36YNLACvH7rsjMmClgVkZ35OF9VXuOL54g+Wol84/k1cX6uB13PO2iFGTGW
9T0kxYrHM579XS8vfLpcvI84rT6nKz6soTX2MSOpMDiPmOoM/4r1a//kcfAC
R3AStnXASsYzit2tbo0WmY7vF4BCDBlHTDyhvaqrK4UmEM5YjS0UdQcOngjQ
Sq3ppX8nSFqvdgQtRT6vzFZFQuIGfCf47xFAUTKjLz82YF5DpKg50WYfXf5G
VUxA8pupgvgLm2IAB4QAA9wiUBVbW78dbwypDpy7Me50Uvjlrc9ALuWHkReF
3OUaff+p5JvYm3vrrniu3Sfs/vAJaOOs9SJYL6gc4bPLdFoYjaR/FWJS5z2u
Q8P2WJ2DSEYdLZVP3bF3r+Z9EnXrzS/1i6IB9zIzp9qhYQk3mLH99FgCadla
dPsk5+h+ykIx3fR645SoIt0CrBnZK6VIainw/v4bMNBTK+NbBWL0a4YvhagG
AGJaeMEKEsAfGc3xfk83GAFKGEC6/vNJmkaEFNRwPuoAUAetjdYzXky2em9g
AIbRhJi8ghHUYztitDmMa9AiUs8wBGL9H7Fhh5Mf6qi8LbMuAEXGr7NJUpFo
apSICmFz7LLp+hXh1f3CFH3zMkXBxeLpgmgw7xQ43dYHPHN2PVQDGkRCvKAa
A3I60l2oA0CqO8M16rIbK89FknYk0Qq254oXkjtgUerQ3/peQuVKkPlkjtOO
s5vfzf4vVcg4abOky8f59/NqlnFFQ1kTk//qX7NmuwHO5uYSiKe9Xua8pwXp
7rRTP1Z7vIKrWM4on+ZKGNqt1aXk3GnbLcyqDcif7n91IWtdYc3TThtTqRIF
RviA1P96NyLFEklqaHHb+rLFzIC64oZjrkt+phs6INmBNDCU79QaX8uPTDCl
WLhM86CFKS7C0tkAFO3Bum6OUUHm637f/oF7jhLfegrplr+BsfWSZ7yJI+Lg
kE8Kpg2ptuDVrI9VTlzQsIYzWT0vr4JO1pwTk0FBep5BMUYmHItyV1Zw/e0i
CvxAtc2+enZHg1Q+Ml0txIc6PCEdLyCR7yVr6qOxPYewXp44QdP1I8wgbr+b
CupuH2Qe2PbL11DQk+fHgGzQe6fEwNvI1oomMK6fq2AC6uUbwDF6D9gM8wfN
IUArO1apksvVSgM86FfnVfc4RSyo8TH/yOkGnN5826K7ZR+ndrxPycaMDPGx
hzG34JO+J70jFFgpwN6k0fqrqTFWDKGwRs4jEJy1GiZg8KLPCrQAQQNPI+S5
vFAtGG8PYTCxiLsoDx22EQmgm7lP3triHF5uikd+GqrNL/pfIWRCiOqwIXby
K+zUFGdqEnCTfOv2TxueruhrNZdsidJCASfS+/fwLCthQG+DpLDTGGsYdm2t
hVYyno1sQjRUrTX1lREK7oM1ZeHaJZKDHcFr2DTPou7neyCC11QanB+WGeav
rHRqzWjsT3TVvHl7fX+6f0WiNZ9nZRi9E3V2y9Xoubm8T7Klec+KDGaIMRgJ
pq8YzSvYBFQwsdJVgEH1uW0rZwJcdq9TiU/E1CWml1OAv4CcynmdK6u+c7DU
/VfEJT6OHvsBtaUxis8zk5ZBKja72MW+zoyB45H9pyxzEjgDsQZPUHvP8tCi
C4ZYskSYXQoRmQCL0mRYiaNFkhFVXqX4bPRasMHLDdspEY6LvF4HPZIhVMAk
jmDYj+4YVCx1dWdr+T5rF/zfrUgT6Ck0RKhqlFys8wIgvfTYSXf+GSbX1z/U
fmBN11ogoS4irhV7OpU8EiMyDrRTMJzDD2WDszMVgoTy7P485QET2e6ViRp7
BXSWzINlATEhMBDEy4VfRcUN3pukLljXQMlFubV1/Rv4741WEIuvxkPhHFTg
kPCpabmx7StP4BdMp0AnRTGorfOmFUWuJ4U7GqjCSf9VeXeYLhilJ1GtxDSj
eyPTQnPX5NmzZbirf2Cic6/YSds0EpwcU4pzpSfI+fjeNTVcNajxYwoLXyHa
BWuVOruyl0hhY/QGrVRUp4odb37SH/vyMcCuu/P7l8FC36kE8IbeEn+GarXK
+SdKZiNcm1gdMnl6jjR6PO+CcKFFo41099cMnZOmKTxpZ8rVecuKBpYUJ/Hg
omL2O+WnE2pU6D+aTgPt3XKzzksgKSU0bB6BWIkZicrHVoQ9aXd8IoSZM2Ko
mhvw1Eoy8HjJG4PuR7mtAz4FPAJSHDsfCY1ueIj0CRtZvbNYy90QVI+N273I
HcXXhnL9129fvDPcW5TXtAQpxZJPbIIijDGv5kb5zOB7vizoJYQDYDj0WmDz
dY6GbqTAyhXSzUARDibb8mC4Gxgf1yV8qGtJx2GxkDRRzK+SjaVTLD2FUjGZ
7h4LQaONvklBkg/x9pB43BJrMWOYEORgpEi1yQ53j5qU4qs65Jt7y0rHRjHM
8Fy76gsZvJrZON6LBnnTu8zgpTn+z00Ox1hbeBFBcSfsQE5Iv5rP5HZjewTb
UxNN+rgdy92nO1T5cW3+rOfAFrgw+sOaV4Q0lxRLS+HVF0f8xkWAOXEn4wDl
r2PUNWIzW2Y9R7ykNBQAfD5PXaineSlBBoAVoi6oY47KMRKeG8P6cu9CZ7x6
MtgYv/axaMbeYOg+QcyVzg4BBMm1YAaYvZhhxyd/lVy/P8HmqmYDtdciGm+y
mRWdyO6bFmQqdKNKdvGzNrQ0lV8lvqYzHXNRUWDguIiYAV65EhV/YQWTT3q+
G3rE9L20NsjIv629v9qg/TCyboWzu3+KLckkcby8DNtRSppY9LxCNtMrgrPz
If/5kitC0fvVG5wLTomLanpf4qj/obe6nfSBQ5hXTr9kEVYFXMbhMJxCakQA
Ie4Fb9M3PgFWt6FV6qaXJzzVoMsEMx9OhGFzn70PAMa+55f3E+y8Kav77SGi
jNc6D0OiBQQ/By2nYnZ3KeTYo8UMiF4zgZQYah16Gckx1Lj7HLNmHsGBALxb
txD+ntUT2Mp6kEKloTWx+HC79TL/sb3jPFftOOGQqt3/YNoy1W3+grTtsoBz
RIUDHxU62gBFLp/SjuhleJVv34+0wahvj7zfYZ/+q6yUAFqOlHJdgIJ6UIZN
q9NwToGRS+aFihvVe89ajSgQY1irAz23M8HeZCCfaQQsztX90SWyAnGbhiV7
dck6de/Tqn7M8FbMUXQ9AGWwEH0kNKNpbe2nuNE36ezsRF5xN20aIGYHVYCv
TzHZCl6Dm2pdIEym5Rzvse1S0ydyjfv5Rnq5tfMNXXBHyJFKVmW5GfKihwrl
VdM7zVUlnhzd0zM6hzQm2YlToc3jyJezaTvrVQxpPOW4F3UNDBGCN/jG7cZ6
+yTA+5X4cAhXlY4kIESAEK1w5ev2XxtLxGu3we+ch2CbteSu774qXm3yG50i
2RWAaafwDmN6Y1hR0cWC7axLbx6Apkn6OyPF+1RsUe226rK5TMagf2P9Pn7i
NRsSE1JhzsLhyE+0ebCzXQ54c61YQ8ryRJLJNnxf2tMnB4LJL04ANP7tGOpS
0Cla4BjE/o73HZ47JD/pQr9MBPKUtGXu6SEaNqg2onMe7o9pxo6gyNvQtdAf
/TSIh8uUDnv+MFZdbtC6etLmAtYWCH7waYg8XxrzjI8g5aRQeOGkO4SODwdP
L11xbDBbslRy5orNhT9hxNmXxDPAXy20qPxR8EfpBqKsTCGBepWLdAYXcziy
ee5B+CrFxfrgBYdZDoQlrZGc3FuFRX42W3++fMxNuK93/xH9dgC5rraalNwT
bc30HgS8HYGz5JutP2vI3uoO7qBMBLqpTVhlB7C+yEZPgG/8SvHab2eTd9db
PB8/MWT9zmKfq6UkFf4YYY7ecsmBB5I0ZtXe0Jixii4zpbmfSfftq7EWU06D
tj2Zxc9lNDYonienD2+mJuWAVefQGon3YPw8kOIVB04m4PNs18CHNcKcUBXV
vDCC/MaZleiSJIPxAyRuPDnkJGtYQLVMQYp9h6GQOFCUfUZgBGx4VzePGhsu
y1ezpv6dun6MrQh5hB1iV+8FKdJ8ihlGf/faZP6zcghazNQLBS9PlxIfrWBP
NCbZMXp+WDU++QV9JBlTqE1P4wrHq3bz+kfD4pwE1Aanna0Z7wxSRwxuvfH0
moJ6Q/3bYTyr20cZ9FNSz1A86Dy2DCgdwOS2k2zBGsTUS/a32VQa/Fb+EVCt
YPLd0Ca/Aay5I9iz6IU/TLoEfJHLGGxsp3qhg0+YjjJmBFmuA0BRDMISH/je
7t82TKqLJDMwmgRtfsBUDvNw2oq4DRure8B0464guWEhoU/d1v28P0YmFFIy
+w9LqJpDrjz3LlIBodFtzEtCR3mBEVbotruf+gZpcu9+VPXLwWS8H2sTP7K2
8cO8G8xtxkkIfrcXEPi5ytJ3UBzbbqZ3MXQ93X3qtGGqh+lBkgt9Vkx5333a
uTW/WntbRiqkkFwDrB2LBW9FtE3F3BkclnpQhHRgoZ/mwrx2FCbU6SCG5RcU
fdVtmkFEPTDaTS4nwl+k8wk8TT67rm7+CS2BXzzitLORyY0PrJBV5V8C8jeY
fjm5C/9l1ErJxWfyI4tQwrAzs6w/ehDRDd7eslyI+4wuXoOUZ6pRe/eyJGvS
p263klkz3vVA3yskbaCYrwY/SYuVY9WzlIRs30TLSTWDmO2uCbsm4N+FwK6n
DqA+L9JpG1f4wMtOwLIhX80D8PRcdqqsdeViLpmqo62mOnK+M6aoTZXtddlJ
fMGzGZQF3n3UlscLdTJ7rol9d+REc+owBhLkJ0CRjCHo/SMSQKsiZAUosZyw
Mc2Rb/hwRER0gn8jGc6KLhHjdx0U+T0WdxdYTK7tL02j/jYvHFu58GfFcYQg
iMPaJY2pPYsyD0vrzy6aOBcaBStKG+zGaS8rpm6QVkyUqiYzgtgen2TNVEtJ
IzZU7Sml6aCnAbKkxp4zvN1asxJgVC4R2870Xq4xXPbWQ3aiki3rspPgLzkm
sbidAfltTZB1mw9QGr+ubfOLoHKNYNJw/QLjV6418bB0nTTFl8DWldGBk94S
kJ9HPUzs7e9HZ2ncSMpq5BdlPvalZ+VlMLXnkES/Ea7hgdQYlpowyzly32Bo
HVWFApSnoO+kcBdagqqPbgvsk+QCv9Tl9FIrBaXF6wDzquD++NxgQ2XNVFwP
emxkh154qb7xFRjwaClF6VyuhxTZTYZW2+v09eMn4R2s9KB28RjmVRypQyiy
w9+Jvgcfqc0nNGfO5nwuoBjnPzvktwCftfirIIDiJDoSWj1LZB8mJvragsEC
sVw6baLIXl6D/M7Y1DHDImVY5W9YNA2AbQkdBoKY4FSepyElXKuvrURxhoYF
8yEb7uF4pFdHuMsZONwNkmCNWEaObqHLM/VjXmZvcNLRq6J31yL6alCCFK8r
MQXEw0l48rsOCDcM73dFJxn6TWYWXMLEvcsDRTFvOct7N//YmzRqahl7UmXV
0467cpd95y+7wRH071D0SyKaQuYZg6gX3jyy10iopDm7NpzCQVfA6C3d0KhI
hKjJhjU9gV+Lf3FYSH6CoMyFeZ9yBrRn2e/hlCRaC7ueQVJ5LKDKfDF+3vpg
Zb93orHtHhXPFHMsuby+LJC0t+y2U/AcdFNBdCzqTmHKNj0r+PC4z4hFD8mc
5pELvL5TH8Qm38HIHn5sr+FDk+VLz3OtmCekdbOMuO98DndHALmfyABk73qC
DcjciA+xvnSPCOY0Q8ghtHxsgXOeBSmpEDPtqncMBmqTKwZzrpDX1tNywSCm
RbzV6hyLlS+mrT+P6pZAiERlL20wdsbBXOklk/k8ITMCs6BAAUt7LhnnEhjK
agGCuNeHuxMcIdoj3W5wSyvAVxrd/wST5JELpA2hRCd7fqXQYACvfV5dYXf3
SJzRmWdYudycuyYNtbtgQ8UoRpM5fCe/LyAeda/1vfPIrFN6x61GkvnnHVHu
ahU9vCFoiflR9lsm/8Ks+VPA8DkvUwNW59CzJVvvjBU6ExKAT3hNQphzpDPA
QDvxnxmLACyhO8XQgGp5ruIdLZV93h3A7TxN0Qh/2TH/WOcyHqVlaGnnfwSG
Y2Z5NZqaPKTh/GbRlGRyYQ2iPHydxFl/I8DRSzkg3yn8EDRjJ0+AU/ClvzgZ
a6EGhSzTL0+xf6dWgzvvjsc1k/bNzKKHbigY2JK6Sy++1YpJ+rroI8CPs1Zw
EDg5Ncp4bjOqU1vzb6V7sM+a5cC4Aj4IY6FjE+gyAQ9H//LC9Tw7SDztTQVj
38JwsTvF/LtsIcp+1zs8wm2ZxgggkCATEk/nicAp3SRgaU0KiYiRave4P9W/
Y1ImFFboVpc8fh+/9miNzpz+WalrUuBqMOyUEAlEq+/g2Yv9SwFimZYvm5tp
AlEY0GT/dFdugJ5Rsgq0fPhI4VvUB9lUO5BD6rPBb8wkFN/nfJVJhsyNSB8e
Cj0DDzxwAvxVWxkXYdpK6KqFk65DAfcVy7iYLcP95SODhcuGXD729KqD7/Tf
jYhvtHhXlmWHwa54LBxmfzzP2H1ipC/pQtNujYFQWEg4l3XqjSFLZGVMCAmT
Z8QHjEWcp2d4F+rQOEajfGin2cOMjCe9zeOhIQ94rB3e/6YrtAn6+2vQyKVe
nz1gC2AZoQvJ9BLbepYa70SwTLfoKJmbxR0oM1TlUjPIVUVpBjegJwXYLLxD
YaleU3z7lC5sAUi8OVJ7sDT+TaBL9MkAtcDyn48y32IqD7zNk+De00kwIy/g
8e8Yhut2PRt9HMGxWEGjJWJuoip15jR/YVeGWviJC1OsTRHZIe/MVuuoc5L5
o3VHPxI7FMBo+STLISCnDaoVnWUBJI5x3MDkFedQakaNPpeNVjiX3G6rhpRo
P79CO3k1pFEr4NGM5A4zqVar5DDzIZ5crZz6AX9Zr0jU6xHnbv7kyyjuOW9C
V6FYI2fds99pR5mA/giz9Ho473nC9GrfMsHcBsNSDSjpNMEur1RY6xtmpPX6
iaIgU71Od5sfIYxli72hG1L/UVhzDoEIEqsxloeIxYQJA3P89WxbKMU4p3bo
LXvhr7XkutdKFxyLvG5uoMuc06L4XDSUmPHmhZTysV8KXL65bplz0B4ty6Fp
1HnQhYugDMgj04ZP2ac8vXtNqoHMC//3MHnU2c7Iy6JCZu3oH8L+wWx4O+Gd
sYiI1Ca8xK+7ScRxfkxh4NPOEj04MxStljKZvqT9wyyolMdR6wn0JCZfGxgB
alJDk/K3JWWcha2bW+liS3DIszSIoSn9ro6akdot7fuu9YtgkIkx4yw40op3
T5uMMgNHO4Q5xobSZAL0HzLc/uxM5Usk3LNLBCcb6gJlIOe6efk4ab7mX/ic
RWOguyOHGQIVBLU7AcYG9xe4myNwUpIm2WG4pTIrBE9JcCgNc4rLNu0voqwU
lgqKXxUHzA/oFRCmwBgof138+13qRSns7Tk6U6PbmhLJxkDV6U02TeVV4VNW
8DlF1LK+BCz5Kg21y/+lr18OByUT24fFlSG+Ffe5F4AhQfoRI0OOv8Jbt9qj
LEFrv+Ry+ibsURF5Ch0JRBFXx7pE2fQk+PCCLDPoVWwVO9X2xQthUUJ8XcTP
y9RqnAjf/b56kzXVQQjCW45dggfcM1La74EtUpEjQwTi1VBvBoZSy5fVxyp9
WU8KGOMZEapbOXBj66q+e2uIfw3bZ2DsUcjLlfodLnEW39sJxT8zvRVxpw0R
IUopBI7Jb7rom6ysO033Rgtsoeq3MvBrWLxsPFpDYDNIKHVl1mJk4R2xpRCD
sHZTyjwWfQdSb16CpfssSnOr9ICwndqHLdTOGQ3v//evOX7nUHLUWwLrXvAF
uMfPEFYkkepH+2MLbNFBdO5AK85g9qgDPYL0ZzjlLVWLfL1ukHhL0zwe43KO
AbuzVl9mzqvDdPtnq08Q8F4A2vrrEsV3VYJCmlg8Lz0SqsfW/xqN0pD6YlUn
0AiVXgLMirAA/thcxfzQ0QJD3ABwHQwqo3j1zvOVqxyDtHY41RhRehNN2sG9
WUTcZhvW7v9yRUYFa8WAqn2lQoH5OYR/dlCMopKkdXtEPxMq6knO8q/Z2dLW
5M5r5uI1VX0FR/oZ/vv+N9aU5Rwp2AWTGeulkWcJuNZF9cN0ZIQ7rCt7zVtN
sW9yvHFzuOEu2skuSWooiBDM4qA5rTGYtIw/IwwYwsAdMegSjcPp5NpDEqQe
ZbOiqqYu4cjQcuZlyh9fnsEfCVQrSXbUhS+6Tt6/6XlPe/CxIrtdCw7cbS/Z
OdXkp8DLIW29tZvYvkDAtelZh51jYg/lSJ42iIIe2qlDVDNR4DLODP9zzJfq
ZxlRq9N0XEtS2O8Gek7gWmu6NitWnmLRQCxN1a8rJxYkCZGmkzEt8Bd/w4nS
XqN4CC98eevp1RnuxjIf4o0YYjELVi2+lAKE5QpcfNwIDs29gwSYjV4egq4E
N9OdWvCAOCLtUm+DrpH+BlS/G/Gkx9Pkq6+A9mofMaOSGyeYPaklAUXqzvdn
gIVEZdnxg+SI/MDDp4xSROaQjbxfyWrZMDELc4fEC/bna3xix5WyrYcvPvhF
pLzSYQfX8OyGf1eZaGRyK2ojS3jzXmvTqu7mjzXznWDkhY21NKbvyGTK2OLW
JxwyUbX7HVYYw+usUCfIYiiqj4hlz9Cjr9KhQxhv3ujULpEqQMO7+EE46mEN
54TqBv+xx7Te7Bsi6dUT+0cjOrfdkiyVgYVbTwQSaCN04+WefGEPCZoHSqeE
NvoVVEVLeegJrP6jf/B89EtlazfOu5UljYc/jvjYz0AjhRYu/NsNL3R6c+Yb
VMu4yHJSa+IHvC9nbQ/Mmy5nXpZEmZCfov/QXKukVfWRc4nOWVHZnIbIUX2+
M/EUYdoEJCDPL7f2CWZxihPhmClUEJET27TTRyKKodWHkx9S70iKc3iGXp3h
g4pfxihFw5y+QEoX2y++DU4LiO3kzuTxzWMimqwvU2Ti210Yy61Xkpc6B2Z+
AqOT+JiLnNJKh26HSiUSrD70ZETpJdxkbJX5szgz5ViZgY6IfbOX6fyK1H+7
x5Z4WO/VGSm16tYjPwW4Xf1CD55jnd77o78O41piiemYxDiCrkTI9qCbMOyD
Hk/xnjsRWC4WxZMcm6KWyyDZgTgfBPfaJwh3CGkcQIGA1jJRwr/lzMNg+e6V
6FWUd76WEYfLI9pIybdKsxWJVX8iT4+7i+s7MBwCQrqJ0qWTqb3eB2uTU91k
jOKWMe8BcURuBxo55ZhrC4sZFFPoCKBtufrKOtVGiUiOU3MWpWZt1KKafPaY
wMSNztWBr/c8ECjHgFMs0lAX5Q9mCVwwE5YUj5rAjahlJAkJK7u0w1wNFmTb
AnpGwEkdRGqm+GYgkSfGtbWk2E9EEGvENi056H/NzWc8Dw66z/PeIewl+H4M
0B4wDATF59FRKnsU2/Nw+U+jiud/6RJdvF2iLiy+0e5S6F95P1m3kiuHYrCi
xiMEaL6zSxXKs4SmjdozZ4uuJUsagUGKttlCGSa83O5xhne8kkdKoHs3/jgW
9uWgSAzQEYbCNhUsP4V9p9pE9Q1Xy4DcZ/DtzpaiAIBtsnC5PuR6haLaAStb
sNoalKi44HIOcvbVkAmWOwhC5JjcrNFfuUXO0Q9vCEc3Ate7HU5tXytpDrPU
vpqO1OwInKAkRH4gouqF79jb5VvZtLfxT3CnzYuDLaXjaVqooY3TA7ROfCPh
9eHciHJRUmuGGAHLZG3czrmIFA7N/vxynJQN/ESYzN2sCT1LXwSBIX0UWq/f
8o+lVuVCGj5Pm7++Eo06sZIaDpdL8MkAy48tVELqe+0ro2M+mTdNlyCN4kAT
WpXoZjtVW9SvtJjPxV+XzBTpRT4Q4Uzb9JviKp7nkLQCQYnxqGk09VNE0w5g
r3tyhHJ7jmzBglxRHc6u9fyXQppppSFVzNLDhJcpUN/uyEPE/Vf0Mb1Y1LfZ
9mZnyZIa4NU2TjhQ4dR48KEnllfk4HxjprvssFg603FW0vSNEwIhtbzoKhnR
FhRfnWdjEcQJbyDBBzwwtgcoX5+e/VefD+pgI9iJFaAMyiA9IAVX/O852lpt
5MzYKIX/Ccs2OM7Y/Osc3oEPilTtH5tLe0KHlNdAzllx8vqaac4hNSAf/ZbM
jmbzS3ZD2zQlHCQLNQ7xJK5gsMB6ACA6N+YN1R5ZlcerdduOAmOVSdAeKDjM
AUfGWBbjXkXlgj3Wcsaogzv/aHLc6v1m6Cb7ihCdgaBtpixY41K4P8vrn1kF
QwD25CTCmBavbpWYVIfUSPqSh6BrHRm8o2Yx6UaqXmJcgpqeY+adnKH8ffH4
9NnmMkvybJIzD7gUHPk/N6G2oKbH/3dgN42YslObe4NuklJ+IaD8umrq2LNw
Rm5D46/jrLPGJIP16+h4KcSp+oHujZ/WUfE3mGLx8KmehTBbNAnXX6h6I5Q5
d5jE2FGdnrzVLV34g5gttkK3kpNEGU7j8x+DPEB/H7o5Ms5Ly0caqL/JNyCC
coWU+qJQAncnA+Wj8Tsilo+JrdWulZwXpEKu1nKCKk0AjMZRFc2KQOLbHYyl
GrYBsVTaOX/Vy4ui1SxRI/GspxkkmFjcPPp99ya+WoNb9g7i262MDiiYOKHH
yVyKC29+j5YpOoPnipRpJ6MzoQzWhZDzQDvAm86wSi+fe6AUbOZUuPtPmlgo
CG562gK0l6cmikQ7cx4LNlbfy3JWm///UD27MaDBDKGDlH1tEySh8ZKggr2b
bGyWcheJO4d/ImVpSH02ZBJYdZAnnXk8Dj9lX8WgY1Qt7FhnfO5NTmfCcNkR
bLpFf7zr9gy5Oe/ZwyceaohzaFZPoM2810LbkT7K21zO4y2sXzTKqEYxyiqd
RJ/vy3ziPrZ1dNZyYgMyRBwXI++QBpxPEutgrMRg1e4/bpxPlyE8skNqsyG6
TxOuA5s3Mmujhw0xscqBvB5a7rmKMzWh7S1is0n+VH0jxWnL2mBh/yQ4iVJz
3d4KFxhD5jxV2HFXkXtdLGJvZHalEOuMN6rXLDJDl3xiZ56/1cz3kJUGBpQ/
SDkTnVSNFkm+eJqVpOzxrJyVd4+tU7UaowfGrXYy+zCfJOMGT8SaUL8jdVAl
7En3PA67+A4JH83v1mkvZ4kj+oKHu4xfp3/siRwE6Fv8Fc8e7RkYp6ZKmlsx
Nk4hNRVm9ZWAswAJsHgDIexeSE8kkTZJF1cEzjTzfQmJ0dpkL+uK6qyAntop
VDxjV/9wfMefSfiI+slUmuaEX6SiL1l0qsaX2XgRNxoYAcEYusJNBUrbG3sU
gkXy/a75MsxSNfBcN3OX4DZ1U6t3eZ1ZKr012EfHuRSO8pD7JuVk+UgqfYHm
CWyMuhv+3eDJHMpc1EIpUNtPg4cJQ7AqpIVY+/JOnACRLnXfe1jVreELqMJc
FT8x6rFtX6TBJjlaTrCmXyIr0GjOzzp5gGPIG228CYSxF5D4+6o/z9mberHc
wPb9HE5KA1FNTNek6dTTD6fNo1w8CnGUeBBSn+M8crgdtr0IJTMLL82NoMRy
i8OzK8thsDBx0ZmtczzcZr4D5kfkGOWcbid5uB7/Rrj6PGTzwsr8DmzRuo/r
annUDO01dNdk4CyWDBq0dXT6EESgxJHgwAG75bLY927Vg6ZGpSrZK76wFQUv
DgDMThuVjXzDP9m8W62oa+CWAWUcbTizRf+Kl3H1HtVolveRMToyr9AGfpZX
2laYg9qzoJAdNnzQ4ym14v+QCXHgxOLvsU3IRFMXt/AGaQFWeRgcwow1AhT9
pebj1b6pc8NuysYCkJV7tiqNY8+MGgQcE8nDn2S39EawOuYjzIOc29rZ1JZF
TPa4lGk/13vLjI7ad6nWWLNTh8QWZfHnrzyfLNnPaMwbgZGmHIjz35ldLf2+
/4YRPXoYGbY4Y3AAG4dQ7uxwr7CwjkFvoRBByOQvcN/vVcC9TgZMafSOXKoV
/IJcQGAKZkh4ecAqIDAXlsCenkIlwmUWmy9MB9arF0ZKu2lu6qBkH/XX1uuK
uUfoqnGa9XrPZn86mogeSSvi3pYN2EX7u2Q1VLkC1JQZnCuFQOECxPalRup2
M9cLSmLhGRo9zVnMz/YUvJzA2m5J5ZgSnlzr/GYI/HPtODSmMw3GXL7OkBJt
ZHZ6PPVNvr0P0BH4KUm44oAJz+JOwTg49nAEJyTaqlo4optFRrou8n4Q7PPq
7KmOSfJVBm3Ra7ml1aUiF/EadTs0mjTOk4pa+/qdaiwYfmkHH6D33wJnDcRk
pTH5x8xjcjF0LcH1LNo+OsVtos1Ra4C7CO+570rVmimMHFue1kAcCZpNVPI3
dYrFgoiU59JtOYIp9s4qzmlY8beiLlgP8PQwU7vrazfSJs5CSTWTrQIdl8VL
a4yo9wWx3O28BCUBAA7A7cdv4CkhX/T/wAQmWpyGKcm45EGk551LuxQFFHAs
L8dH4u0jCFIjHY0Ey3Q3Drhzouq/AUVRIU6NzL6QtMuIGY/augdBMfAuu7ol
O3QhzAa04j0ovXT/ZSCvhq+s2EaCQUISUg00nmIx7K+w9IAkjKxA/Rj6IZ+/
y07AAqCXUiuhjoQA7crIbD1ez6l9lm/u6id+xtSvwb8qmILZ93Tc+NJDH/TU
9Yy0INy8cqdIhat5QfjTGA0bvs64UYnI2hqSAgWPBGvTBog6TCcHbrN77iYA
/OYwYrZxTX69uQIw7LDNpjmDwCAxHZDCZncM+9rPnLi6yY3XS5EqewDLeFTh
00r0rgn5d9eV0ONScgtgFIR7qX7LpR7ESigHsbu6Hacf3Mq/J18b5iZl7vYI
Ex3+x9TfMpHxzTsbiBkVz+67fQDRhsyI5SGP6hL4ckof3ASdr2yaL6psAMm6
YZ6bzF7VOCEs8m/vk4Fw7C78DrMautJQce1tZKGFyZHSxsTcKJA08VjAef7j
xSkYqyK5s6QZMcfZ/DoibampbETsey2IK6KXOc2E5jDeN19kaimf9II8yzUL
1un/EtX8NCDBupEpl/RSCqlxJ1/Cfbf2CmDjy/36tnignciLQbkk7UwcrJ3C
/QiA+Ep19W9VoU4qbWz56sbY3VVmRzne8QI52EHHcPw+c8PY6MmcEh6guLo2
ayVCOmvXF8Dv01nx73mDD1TlQDWKCnZF65umeLbHUuS65cp4KjLxWQrdh092
P23N+l0nwtoX7wdgynGFgVHxaW9s05e9pdLH//owjAXH2JH/YKxTDmOu4Ayv
Hxzw2J8ZPSizPWsRNK1sB6EGdg5IQ/sDM8G52LKGH5hVVKDnb1FaywkzhlW4
T/s+MVRrgqLd9psPvJ86th9BPoNom0X/nXdqAeXm/uzKqiLrXQ7S/wxU3VzN
P0mTwDtZQUG3KXBkjSGnIj8QcCDikGmZ6TKQO0+Z3evWHoQ90SWElTnTkRZg
fO4OMVBSOQ1GvOECAkHT9pGcMQb2wVgqwo2zDznQoaEpPJo412O5Cu3HV4OM
G/JowE8cazzniIHV+LMT+1pMqg97hKbP8dJNB4uqSsUwEQanJWHY6pTVGc0Z
qnTHTJ8D00cb0eGFzLJ7/9ZW2L7zfMUcB0K+Xf+/TDFabbVrcv7Q+GEpcU5m
67ScS3pcJefVRvs1GNzhdXU6OOfiApztlHc2FTAt9NU7jl4gUHwP+AblCvaM
L0QWTb12QHPBjSdHMTgNvded1H09i41vWmqExU92LE673+blBlD+acHlTJQj
A/8pYwV2gTx6qYIjfdRzNlhXBbsxUYpOTi6sQ9bXS8AF7oNfYjaXf+Oitaqh
UrXQ1v52PgXiPFA2YDQyB/p7NkUcxBUxX3iD+eV8Ev1XfW44gzklr8/xnucy
4MQMeDQEyUjCq+/MI4PfeZc5wqMXNxOlwj1MdbOIlCieri9pRHJEBBg7PlGZ
+lr5b5WUVW52O9r2EBY5+PZmXasqw9Ne4PW5QdLc8jh94djGJQW8Q9UhUBR6
C/hpLLcoVxomajXjlHJhuoP1b6HGB3ndRsMuxBLK284RbykqhqsaEeamSk2I
2lB6yRa43sCoMVWrUXp/6P37XuESJuXq1/YsNFvN7ieO7GcU1gS0t180/HBS
y11J3R0vaPnv/Fyi20nTfWQUE3rUFQPP4TXeNNHBsT6hqHE87Cym9k3zt9ll
wUmAspDV+yiYJdstyW0sMq3uOFxH7NX+XJxT/Hn177spniwVPPOHkcU+GtVA
MyobxF9m3lR2WBooZL3Iq03Zh3U8UVZEyw63om3yqSi+AvHDnoUKmaTF4Vr/
RRAiKDBxTLC1BFk2cBXmqVT+/vLy14QHbqvrjVt6kBsLnaXRvGAlepwgofOR
jCH4pSLJPXoVxOugLl/ngaFiGAqvFPgo37azH3rBzRA1K3OC+Vw4KNlKGg3O
Rz6DNfsLH8hVqG/fWZk0wWbJrbSgov+HeMM8QRK5qiX1qSCtlR5GTx4Mr/to
12oYe/eOhicOJyIGrejxLLt/LkOu3zLnAnO/i3w8TzpNgGIDcSaPad1fbP5B
sVD23rEOUXx/VRNO6H4kGphUZyMXg/ykYhVOe5oRkbDf3Ud+1Z+Qe/QTh8fs
4OVdV99GAOFNaMMjn9N1jCTmfkt0jEoM8h+fM6WXIuSSghBw8Q7zRtrr6T/M
Ih9GYpg8DWtltQIYW5e4NO8/dFFBL0VCd47VDchltioXJbxhQmliHHIJdqEb
KYUo1HwZW/XJA0+eD2nKmcCHOimJWF/sqs3WW5Nkz3Zgtkyykj8OTIa7DE/4
KcXKXLlJaGJ2KVA9qcy/gLCVFNb6v/jCf9z2xTHI9jC4en+QQVpQ55ZNzcHM
2mf7Nxd/GEnxHN3qefFIxx3/u9LIYmr6AFaJfdN2WEcszukyU0cxvq57sYRd
5LULnh3W/B4TZZ2+isJKjtfRl5uyR4Of/jzdP8lk49i6SRQXJrnbaJlbcj+k
INhnoYSrt3hLfgJgLk1GauyBKclHtrBO/vYLPwlrRYXJoy+Zaum7L+KbiNwm
UPluM+S5fy/odCajGXfCDODDIwinamLcU5yqvIB0vmt3OuP0OjesCRCdfVwo
+7JewkVHh6OjHu7l27P5itc4KevxIyfCFqNbFlg7RUOecnPI0jMGS4rDa1iD
agqWrUdpzE+l3Lsiv2dTRZWrxx3PjSmqswWvY0W1QDtJ9lofJbDEeYdWwbvg
KFFGw88orUanD13C9eWAZ20pwfEghweeyG2I2v5bJnrKs856xCg+90dTXC0w
fF2BH+doII6VkIIFVJFoZYmzQBdE732DIxMtG9mg3YYH5W8HY34e5m/NESQv
T+EGUtWKY3jZm9q3Lr3jwyhtDdyAilTjlqXtCKLD1xn7ZbMBjRM7Ph+6TM+B
dU0qtANGMx7+l3a+ntycnID1irvYq2F8JylyH50EQ1ePdMk/HnuyPGJMP39h
UGwRClETHWL/TfjcxT3gDR5SOZiPiSgQ3N7PTzYjKtNCJPIMwNGFl8KiuHJX
pqehMygkw0mgJlpQ/tNxSeDrlJRKN8zbLNQwh0Zr4J5eOV+SK/I12CZ968j7
5UL+UssMwfhDxSX0oukXMVT+voJu6RNPXlkU6q/hb6GxdoBi6aO93iqofzOu
Q7KLB8mzSnPN8K0EoCsAz2HsFrGkZ77/NAqbPWrh1s1vL/+W46dt9A5Yagb5
vuhqbjAqzoMlfweEiWuYJ7EpEjwvGji97ioEvqanIT1JG0I63TRpHjCoZOhD
aaleT2gNfmgBBiODPkRy/AipFkCHH33MDzMubHdXZPJMUcBJkeacP5XbZvJG
r7q3np4FdQEuFEhwvHJrsZDqXyaUZv29eoDZxPFRSazlwdOM50O93X5W6K/I
Ujbes9n6QUu62CDKWcw2XUvzoAqWm+Y8p36oJDSz/t9r4kM/5udkYambNSK7
rNuE/DbLuuy6Vud5pBp+8O/cZ4+dee+OcMDxj8GmPnkMkD7+jsYejYw2/OWc
hSuXyzP8amzvJA66AxkacHk4EPb+k/AWUhqzINtmad1s2i1B9hiHaJSf4uhN
wAHncR2V8bOEPVlOJVQqOHghz5zv8klAhNRtaJtnhA6rAkl3gam1MGfbR0r4
9wspCbgL0saXl7QHmYEKNNEM3Ur/bXD1NWGDhGIcMyhINtePPLxifcymye4p
ej3tnErg9XKMtLagFZUbU228EKkCRHNfkD4NY2art9VwsXrcj+0N3ZTwpMgW
1s+Z0zf4+SSxqctEj6rqrDKQsQM72pilO1dklQ7Ng1vuD5uI5S+AmBD2kye9
g0AmTnsag6GBcA247AcAthlus6ALUk/6wabEjcjtDBjOKI75DDVzULN5Oa6E
usIXLnAKISlkR9m0he0BqNrnucE/sKG7La8eOJiCawm6DJZ4XuoYItnugL5l
kia2YqdHe9d/ckydqQc30y2EFBqnRZWbDKBTUvCy0R+hqnS+suYx4b0FEgG/
lH/BnJWHCeS45KuVDyPc6zYmMvfoWZEeniLHsrH1zSMwcX+kN6uuLC4eHuwZ
Nj6LSqatIzfsXh84LWmsFvBIHxJMckS1hDhB0e2NbBwvxt7tIpX1Q2XYnOAr
PSoVQQAaxKF2CFwK04ngjOBJBGpFph3Zc5eJCXLXMZD1JXJFGC5xv/Y4HxDo
yLHFMAPTlTsUGkt3Zac5t0KIHs82bId9PVN846sbg5gHkDwj78qyrPIjofxB
DS6Y72Nz3OIlWZ5A2jHPKZaK5R1LUMtD1GbloPpV+RDt0w1thP9Zsls0a9EB
omb9LbHO58ljF9NUUYBA04nZpHptSx4VsCOlDoL+bhx8Ae2NdVtBTqOriDqm
9yTk1Oy3Y7Mg+3u0BRoHwiiOwauZUMUNks/NiVpUuJYNxB4rWnmppxY83JX5
GJp1CRA+k0mpY+9k5qWtYDpAek/fs8pSOVK1jVn/x4sR1ecI9OCrgmQ9VEje
Nrr5c0Qm3E/jedDUPJ/qfjI7P8/ZHp//cRlwv1rm88Otk2EJFyTXctvgTZwK
deI7n7yKiY+Z4UiwEQzp+E7+fUb5tbHECEYYjznGgzI5GKPxli80YyKUqRW0
qzP5zlKUiSDpak5hXXfmzBLdbkzyc3yDy8nbIJldU3mN2NIOMkhJ//RMUwWk
Kwug/EBevp3kUkoJkw3D7kOz3/SjxpIJpmcCUaMrLxlhE4V2qhw8Gxt5Nt5M
QNonwRAqK4e/rL8XCYByW8G5yHFs3J6OR8RSY+wyoomI3a6NpamKtOiZQztC
v0qVpg7RxjBbQJKqamvjaMh3HJPUFocUTxnbhRIrAZqA13Y+cDiQMQFg0F3r
WRB4AZTi9HsgXAse3SIcbGW2lNnm7YhHr5E7cxGnmqD+07TcOIXxIPN9DJ5c
e39ceLTvdzUcShruzuYM4bYSJYCA1H43X7Q9/cw014uzWU5Ddp4uDKBBf6NK
rTEPztZ2ncCQ7ZKwgZW7RX83o4SjGcqREz9AQYvIFfJ8DxenEcMrfc10VbLD
LzYwTtSSQbytrfN1HI2lVQI9qhzqCmHvQzQ2yEcGmp7B6iRJQ+AfZMx2CSi5
mp0Rg9Ju6NAK1MKmSDjuO+1aBkk3fmat5dROFf2uCkRMTGsvqZQfdYUXBJlE
F6Cppyhh26TNCiCZQzfAlgLmIZ7oy1ACkInyxrheB9N/AA/LJLNzhNodFHLW
E/Jgra0DZ+vpYcpL8TwyUcCxDkRAB7kmOLttKhdD+2FNP+7zDaPbgxlPItOg
mIOUPIVt7cKJAoNjUU4r8uP4yubqm9FOlCGGGzf8+d3LCGTdgkNaGzwY84ex
Fx0VuYkFeCYPlspXz6+szb5UaSISmySovA//h/NlvBFywcdgtwYs/k7QD2uN
4NICm15pKb+tZqb4hWfjSJ4UL8AfNx6YGSQ/wpZN6HjVLXocNNtB0vDqvdJy
yCVd9DXCXKHdX67QucNCKoOTyUC4c4or9YrnXI8MIbF1h9lYDnaiiMo9Cukv
BaseXId6dV8Ctz9RDAbs7uyRgVNQz6onv/J7ciIH1OpOasnMHm6GU0aq/x1E
ksipG1srDDJtfm1a51MGGp8/zFIB0ZUouVFNDte2TxCMtS2+J5kRQdvy9N8+
uKsvhy9YWWgpYt4lL3DqwL/99/wTvgufiCUaKOEHc7khlxJf3F0mSdgozgs4
r6m3FAd4pSGwbkfvx4S/JhiP2Dl1sFYyGxc80/OoDazRmDpNvodinD0bAt5q
Z6+MO6+S8NZAMRRdW7Jkb95DMtJDTHWq8h4DlgBtIz06XgMWGy8pcdN9Cea8
m1Oe3mLpiy3SI/wBmBAJNlBiJbPETkh4SrDjolMNkrsCb4XV6HC/e9vWRWPs
Arivq06TNo3OUMgU3nuuDEMKTzfOHG1mvMO+O7a/Z2nI7Pt/AymLGD7RjOTj
jf339hJ1inB+vxy890rN9WPpB6qi39Ao75zDdSvqv39U1kZ4zzkr50WRM+CO
YjM9j+U1+BJsRl0trn9gjG1pKsHHyd++Vf6Asf3eHZ17+jFckiRJvohtrlwW
GzdqKuMm/TZPZa1HYX8OYP6h2fkZvrMJY0GnNKj8s8RVsKRgnRIvk+Z1BbyC
iA0igJWvJNSW4xyRD7T5N8Ryc47v6QPrZQlwD4OVvwRAVknhk3RDpvUVSAgC
oCBPCEEakyAwZN8P89ECNtBeXpst5Hmuyar0UQBsjQBLX/px2i334DpHzK2j
eSRfNn0g7t8ZYnYWwYl9nxp99OJNCOC7nd7T8L/UC3EE1EGKTuh+/nx+Rz3F
hwAdKenHgGWrwJA7b/UNSm5skX1toNzTxAJJPVW989UwnMcpJYNp2jKypYuG
J2sB2h85dtTNQuvuRM2rOXwK978C0q8l7Sau79FnAQE5Z1iEEaJzLJ5UVL9l
lSmuEcPKAoC7/n+JaA07+bm++G6sOvPU+ZHYushCFwnDFkhhX5bIMGrqhtVr
8/o/K/IGub/IN0ysdC6pV/zWuzVUZjJcbqmEfDxAw2F8HjIZtxGaxawC23ZF
ZFN2+s8/rTk3uBSSBJ/UJiH+vfWrrDuLmzFmw8hUby+YOX59us8H3y0zSNtY
322KvO/jer3gZKfTDlJb0T3jHF1tlNXjPUOrcBjwxAfSN/uAQ6dW4GaMaOgP
+OqXJmEjLOn400xqdwwtS0tVAdFgzIw5Kd9OrVcgJC1OB5AJvB3KjdHUPKcS
qehgRo2iRep/vezXrgaiY1gtHEcaXid3QiUWR3Dq0r9Hg4wrajq3n8UR1dH8
3YJqSYyIoFQ/7K6Ikt++vKsKKvW7JUSVKuRIL4cEveZ4yc+98PEX1VG6TQmB
8vos+tDbCp3ohgEe7aCOYidoXz3+V4NWeJmjNOl0wdW3M0gmKqQ1qvD2GeUj
s5cT7ls4NQ+xtZasKo/PMB2ZjIQ6VbRRqN4IrSSGRPcrbdpVhgxMVjSnoiWI
dNJ06yuT2KKbS16V7l6RmVCnZSR7vRq+VUv8dZwLfRfc/s1jYgHIK/Vt2//B
iYlXWZ/kFCKm3siF9P0Q0SzM2vCLC/U7rTlKiniBVt50OQdpdLrQb+qkbIjy
73z1M8PhydcSIfRsNxSD9rtO7luzJxRrLlsw7ZxvwlmWEeoFe1QBqGCLBv0d
e6vEqCivJUqrm8oCN0fz196RZGyXVjHMkKteMHj7fBrh2xES3pnUiZ6CYBFz
cjIlg84B3xmsbwVKvW7H4afx13rMKS7Y33T1bsI1GTjHiaO4hDr30jWKeASD
QBf0pBKWRq/ec9QcBgK+cAhvn+x5ICI54XrGzdwd9VHAtv3gPTQRzU3oqgUZ
ez+vNlELmcNK/jyM+uC9kPfReJfQJxeIZQXZ8YdUlQiXRyxm19eLL8W1qfRM
lNos/NQgnBmSwySl+K683MLCu/NRRmDgaZSBJSofQm0ZmCcd9aPVVB/A9tDV
zZOaj6sfBAMEAkbI8rPYSqokQzjkDvIgInDhB2AJXk6fHGSaAuvf64dSuxU7
UwAWlJAPa8kbZUfjpAy563I9D+xxQojmQMCN9PsOtxmD3RpD6L22DONvYHrX
hlWpQkmki6k623SaB1iqKZw8lPdO1ipukyqLjQZvul8Wt7Fy2snxIaOFkKBz
6jnfSeWhVxi4xBasllmr0lVbj+OLGEp5gc8uiqwWNeWeTheRUQh/cMQQk4Pe
kjY4MAhd3Jxx8ipmSVBoARcuM1pEXCGVpNoCLa5Z6nz2kV+quNwMW8qu55w9
PHtBck+Zs30/o5QseYzF8aekg7jZHhFAGZjiMrMty+4V5wK6RH/Xkeznbue/
GI2+1PhICETXrb4en4IGZLUr0otWQM98uUJuxH2oQfg8j44tUDDTZAox9cm/
ETswnA50F8oPF/6RycxbVpsdFY0KwtFGnO8bGG35O/nRJyTpWpEsi0/fWi6N
SzSQK/cCjpWlcttZcL85PVJ118eWdkBgu0AJOTln6QokCCXeNCsKqz8RElwh
vw+hUh7HiWmgXeIxsf0T0JYo3QGuO4ReTGAQWwQei/JfolrpiTS8w+dLVoOG
l8m60oXOxk7AsFwLRKFhhFyI9l9YrcJWWS7wfvTYfNyoECyFo4/paQOVIqCQ
QkfmWnt10XTWiDavuq/dRh+Rm0aW0a2R0Y4e8jSqvttOJ/AxZTHm8zgtAI4Z
oct4MeK2q0bvEN0yWAAE2wZKUXtWUyiXEWPo3GPiDhIih4rbQ57gRGGxYFzf
2ZAXWwWmn7JoBjbs+nRG08v+7MZ2gqj2Ay3JTYXVeDo4oNlTr1QhJXNCW5m9
I5SxSneppiTa0rgUA8HovmMUXLebZ7A322EXdPJ2Vc+VAe3+N0CcPVVL7L0e
ns4YTJ4UFnTw44pjXQR8kyb1cql0GYqtoPr9YqfBvE0qRrV4Zp9AgGxRzlIE
voowqFkrA41yA1+2AvFmtg5NPS4liFSbu8+PC502tRa6oFBeWxc0Bx8+gJ0K
PDZLj5RRK874VFl2le9OqD0dnjFNJbDfhAygJMFh8dTHcrF9JqTsurEkAiW3
2UJRp1xjjH9kqETT6YM9vURnIbMtaKh6no7RM/IGrmo2DI5LRLwN1mqbtQRn
RHtAaBvFgnuLD2WJirEG78uvcS0SYwMmRHh2J3JFSl6MxtRiRQBPz+kEOpJ9
NtUEIF4aPu4O/4K4Vg45Mz2B6vVmNIvIPHnt0u/tTMBJIeza92M7K7yQmngO
9KRIshsV6BjCih6eHqZa4YRN46KXcmieQATF5vCBFhzxgDAnnDEI7MdaHuSw
/UmgIhqkCAzFuYZVI7jUXy41V2hRPj0On4Ro+q20xuOSIqeOmlYKCG8CbJ5K
rEYfHzjyKJigJvorptxm7hOp+Kpg3PklJ8i1cUMKSFy4sPffZPBor1PTl+/t
oTRJzInpOQuGHkHCUUg0J8AME6+lJVrH9On4esdg9XI4a1Wm3vS9utdRVnjb
35PTJpu//Rvw4aDmZusO3FQnWDd7iKJMfefhX6IEeAXZdOFVmeujJDx8BFTE
tzu/H0UFvIT5ylBfw/spZiH3cN6UXv1vCH9X/Eq5LJk/HLJWr/aYVYJ8LoIm
DjVH1rTO+l45fMR7ekwRIgCQGnFdGTbYsyGZlLUoKqLSxob+uh1lP1UtMaTE
5eOmtT7DVTpdSweWIdSbJZEk9em4A8e6lw/JCNiQtskqQ3QDYy8hbCwdZnb4
oPTNOkzMLNX7kTL4Ex3v5LHO/4CAu1J3BcQNWwoWZIgzHgiaDJ060WdisZxJ
AlJycT83QgsIMGTBbVQSaBO0pKs+yjIyts5XsM/efvI1Jo7bZPWafJNvgGEH
7g/G3W8nA7lcbYBjh2e83J4TTIEmXhLj8hU8HX9thlgpoBnTvapjUx5m/EdI
M7CdsyNyrFHjeUg3q5lIpD9PvS3Ffn6v5ovWB8SCGaQgSW8iWw9kfQl1oBJp
JXIdLuL+LeB9HYk+x0Q01kpfAW1SdwJxWaaHzwkAJSFLGaYYhMf+nl8wPw92
kPzrHnxv73I/UU+z28OnXWylGtTnr/G8x33qHWkObtveNBb5FXa2XPaCZfzX
u8c8Rz6KmIiT+abxhZkA3v7JgCZHO+1D3fFQzhtvatzn1dVM3CT1rt5mgVr9
5U75TubVTp44HKK69LBBdlVRjLb/PY4Bk4AaYaqzBc7xX5cgXOsZKvfk8uzo
f3y3alprq2HU8G0zuT5SDXNIKSyvcj2c0aJOVJcpYmdVs1v2CNYgDTYGRKpc
OUqalZB1MUAMLibPvJJltQ2l7H7jR9n7vM8X26FV46nlLawQQV38C1WhD9hs
BAskg1mPDVHZgZ9t3uTbcb2Y+Cdlobne7N4CIaTfxmFj/YAoagFAeLe4TaAR
pwMSejmCgyYokeRn17slDf/2Tg72rdH5XEgKXve5c1YPNNoNreE0m2ik1ZzM
y7OIs7/ZTSmty1lLs6vi9Fa+WZG+ot4083FA28wlsABsz3ss1k2+tFT6ld4E
VxtrGE+LtFML4cjIQakg3rP9TI51eZyMH9vhbYmh2UTLRbzgIxWI3eRADup1
gkiDCxPnL4ZJFxM85J11/S0VJBWkDhWZOMS+Sh2pMowIEULIsBX1UK7XgVrp
MEO9yxNE9ba1YS3gcZIrNjBCC6xyp0HWE7dpIGXhWwgEfHrLI99sy0cXH1/P
8Let4hWbWKxfwNDPo3+Qr0BB+LWHRqh5iyy5WFTCXKPeveGkgMxsfYfnR/vT
KkLL0EoHAnhL0ii4BS4xvFl18fdqKqLcJveCc/DUBa+1NEsdiP0DLX1LY3i5
amNXwaswDUzUPlvRqn2j5EhnJnL+jSx+4oGfog9Ynnt+2eck72U/YrzfE29D
A3SkiJXl3ctVoJlf3em4GMm+E/ziBZsurJj6YSLIlU/ncgqs0RcA937n5hsE
rALnIbgVnXdDvYjex4enVGALRC7wU/sGLnFm6aluyi/S13kNFCIy7qa87uVU
SH0NGfVw1mj8ePjjV3Q9nn6piHi18E9hapa91v3ZiPNzK6TVZ9jrEbkaBH2+
fmw/vvfc/zWOEfetrPLkDp6Og6fs8QAW3aLSwW4A+daiPejDYfQ6VCxd7UIC
yZKotJqANpIIkcDNPUg/rHXIjXkUVvob+FPvV6suLKbTmyW7rfZCY5cfpnF9
UlDU/x0sf4wmvNZz49+SLP3apt3V8VoyZDeYv2f4rbpjUuyGIsSB+1ciCbdC
viacAbEPwDSGc5yKxwzHnrt3QndVjm64mR8DlCmkW15GAE1gzV7emPU7tBYR
lmypwoN4teArQbdcIYR4VXmSRF/SpLzFKKHV77p5gs/f0LoeQo1J7o5naX3y
6HqwbBWdL2S0rFPar5sbRN6bQZQ+JjL1KM8pmU0U7+afknjxj5P/DSxXTsjp
hpaGIM/qrXW3bvzkfmPuXD2CsAeZ+GsnbVc0QrPkOaLomg9tHKfRVMQQfgaH
420vraZaV+wKvPjyUhX1g5Ktit8XbBXlIgveKieVaISqE2dM66s0w4Szh+fU
O/BPOaZD7WHp/eZntmbRETKw2Jn/4dFsuF11wM5pCYHV4zABA93+gnMhowjN
UPZ7M+Gn+c6HBC4+Vp2na/341YpPMRLdd2TUT0Qz7VnzHDkClUonMbuS41wE
G6w2fAotoGk30O+HhwiyAJDcZag+/NpbWMm5PIeZmSxn0XpA99xgrqF7CQrn
E9x20YmxCBl7ibRiTfdbZAPWkm5kMHu9O2Iz0zv57ay5aUbsw91I57Z5vCq5
1cuT/6hNtcHdtECtxEBakF0ioXF5e1gRpF6u8xuY0DbGwcbgjnzvyYHZw6fG
ymFiUXVu6MfGIcp1h+XCO4OnL9ClOM3k7C8CU/YFu3gpd5n6k8idVm0LX/3n
qyZPLrZIqPWRwDJrs3bf0Yzf2zpzQJfQX5rb6F/bjEiBckXSx+FFUgRpPROM
nddXQnJWZcJUQKULgkkA/2DQfDHPdudpC8X0j7yIPT6KPpYtCCj1tLzAgIy7
4YHl6W6DeM5Qjc2Bi1apOY2MN9aPB2zHQdKLJEjLbEtzHlMmaQN+apx16guh
moC0rMTE10Qa1OT+WhepVenVDpPZiiDzRtS1e91rqcxubUERsaeJXZh0nXJx
lX2cVmWKSFg5a6BH3FYQCPR6pbkjrsbJ7Ky1CMQdcdnfVyr0wTkFG8itIPXA
PjZfPc6aptjiVAROdF2jK2AvRXVWjCuHf32Mnr12x+x82bV9B9PvvYsE7HRd
9Vg5xtkwGlKA8Lwls8IHMb2uoJSitm6R5hwNh8vXjPp568tD4qOExevblPnx
5ojG0ZLgzp14lsS5tMFwRSmLHa8Qe7lizFjvvh41WlggbDxIP9w3jGsNLKWj
i3hKS7ygIZbVvzzyNdF68cXzpAaOA/tDUnb0/c6/uU2uTO0dYgfrjr9FwTvt
7RJ2QlRIlod2QITsAcf568BOFTG/ClcEbeUGmVmPeAhrHMNG8PNVlb0j1gFz
A9lOjvYYzR1EWuWOkCz2/f0hCkQsJg1IN38ZsyAQAxFajRz9Vpos5suR8Qj6
UioT2oJZuxKBJ0B1BIHQ7ztzB4JDZX0PXufko8gr1I5yQ7/RN7oi425RBMQs
ww1MVdID9Qq+ovrupPgK6kXt+S8MobZN17hHNmmzyHUKGGnI72PF9A/CsD+I
bymwD0KYmaqIiSH82Mg8bkYdjPGJOq9GKkp+I89beGKI4I0dmcKSWKOl9eLT
i20E9wV9y4Jzdan/x3co+pQUxgWTXOv3z6sqAoYanqa5OJTwWSevbWMh7Sae
WTtba9WuAFFZRyqH27tKH8ou609k4yJ5krYMI+dl/NAi5R5kSMB/+DNC6zT2
8m9d6akPGj4nk9qeN+wFsQ8W0po56pfak7y9ric5Uk7RPgAcVcOPiKmUN9DM
kAWHlByififq/I8UkgJiCbF7BV+74RezLRHNxw6N0OekAESwJI3xgzr5vVS4
LLAzJmXGO50+ZQgdJMCBVFU0N7G9i8Qu+WzOacEuZQAYPQmUmgtSAy45DAR7
faCVDzrlk2gLupim7VydS0mYR6Ut0Tsmqy7GvcD1WrORTKIQNC7EPB2CxmYn
tLaBzNxWpMiwfVFzkSjKT+hJf7jp9iaHlmpKbGsb4twW6cuvxVLVBihXn4Bz
MtWdLSP+sEPYD4nm/6tVZeuAn22MzmEIejmGauyO4+NjijNuIo2hHIV0ZO4W
y+KdHHuYGv/sKEu8MBKmF0esjYkmeKFjw7wgFF7FdScWvAbESfO870WlBWAa
PUfX0KUQMFxIyPiEwTDFqwuF6b6ddLsM0jdtM4PR32aXCMNkaoYLQt1uwxf4
I/wZ+pT1R1WciXDwKIdGnQGgzQcAV7M1M2JuZBAtlAxP8ZSDjICXqakjuYgv
cXDyvmqmi07C6BA83xj9+21jbcr2ObcaRAZicagXUgbcRZ58vjXaD9iD8Q5V
OtXahKjpN9H8SrIZajBSXiuf+B/xgOkdhZBN1d7isitAPvQaesj7Mz0r6l55
WJ3YUnutw4ebwu1sm/AuZlVrY/vtCYmCRacKVi4sxifyhutcl1QbiYwmLBqW
clOpte7s6rEG1pBP+eFaaJ6nVWVRFYW6WJIZBtwYnN0J5IyGWRcQdHpG0FX9
O7XU/aGxaT/ssJmnzQ9OkaSnb7UjmnavtFJZ/YhY2yN1gaczGwzS98N+wd5s
6GakJEpwIQ5IYglWTfR+sk6esVbPcVM8OCMSl6LUgyYyyTEEHbyZr6hYEIw9
Rra7j0MeMmEpL5P72iBmMzUhLl92cT90LjntdraW3KqHzhUOc2cKf8rpuMxZ
GrEQyi/jThckG0a7Bu+1wmFb3lCM5nmM3UItfxDAA8HjCYZgmCaqO2tebR2a
84W5YPaiunv8lefqhg1J9DvCmS594juTRjhAdEU3iBFOs4Fq9YhVcK551gcd
5S2Zys4Detyu+H+5z9z+gm61zAuDQEPii+3QcTJonwyPHmt76eg7ELQ345Qp
SlgEA77aCyQwwNAf2MB7FxjGwDnSskk7NQB27zFACM0hYEddW+3DrkNQ7ewU
vlb3vJqG1+n+uV124W+n9O9eO/t3JWeubvHcrYglVu8Wpqeaw/dtG19lIxgg
/IEAmvAZVrmJQs9aEEbXS6KoGt90DWujfQ4BL256u6sydwn5Z+nIB+4OLZUJ
hbvEsgYpFigDXLf6JLKgw0R+kZ8VYVhfm+eI+4WVqGQIpEGOmBlhlkaZd+r5
ZIC8Xm7ntdeRRah0DxFNgONp7nVrB5x7wo530h7re7DSn6qO4a19NPRa47c3
JPOR4YveDQAWsAWw5LWWW0yFO8qHbUF/tLQy7/YlIoHw09TcKRwhI/PP2Ucp
C1duSRt0tw5bsOlDoiZPG+FRRa/COW9UqJ8HD5Ex4IrImwE9lHn63aq8mr74
v3il+qjgFida7QtZsXFnZUKe9rbG5FEtosss+suxe26dGao/G2BXozGT0rld
MmYgHdPuKGG04/TukjwWuO96idapLKEHc72vSI4BJZ9dO/k1rbm0DjeR0keg
NJrP6KjighscpNqSCCIROTZlUD7375onw3y+ZZorz2ok9ld8cE9OSW+HCPP4
HRRIG1+n1KTcTmtnljvz0ZOrgFe9buS3hA3f1DlXAmDscWmgds26f/47PG6W
xL74xH5DEdi91n4c2VihVs+LTe4L5b7vNvaYTWDjNUeyJMcbVltg1srJ1MTp
IXemxfOh/gslF9N8qSDdGkSq+au5mL4OhMobacncmJnRZulHmvhTm9ZEIORi
GnMFLYmj/PbrKRfAsxkWoN7aHeu8jl/UlvIz+fcil4hFYO3b+dF+JBTETUqf
TJNkybrMkjvPe4uPCdEJw3b/yUl7z3l0WsMdDgesFOkMWayQ8KJZifbrIoXT
fLsrc9O3zfPTiTR/FvzjHeRvl/vaZqk2DfGUMpQEXw+o4BxJHvLzdhDLVFqC
EBmraOhJNnvFi6pGQj7/jiOIRvLMnQxgQvkLPVeTLAGxRfpmQ2zyJAhaHn7j
QPLQemIT416nr1fwzjCMFehzn5dzqaOUhYszyXPPaIWUrYZJAxEFqszAIxmv
cHAeaiQy/byd9wrOXbPBSzQZPZ2aCOBnvN7clHEnPc1kSsPGhVpUvQO5+g6l
OCN4B45s00liivOBSAm9271aYCIknyAetva47uvv8J8nbU7ay7OszM+gF3h9
aEAtdg86497LruLzJb9i+NGqAWbt6+1fcClKHDLxnBIQ6PIdX+FgsCUNltt9
+kBoFdwNgYvy09uT9Rbio+EJTdGfB/L79sNiEg5AUWyPx7dhUI+KHboyqDr9
9vsOy99wLVJ1R6sSbcIKgJdKBeAEhP4y+IOWlRVaq12RaZIpLxdMtbPrbwpA
IGLlXjmfHO5RGo+QQs7np8uj/Cs0S+Nn0vfNqXojlcw6+DZW0o61NaDCWlNy
LVYqXs10bCVSky4AHAgua1TKQ+V+g8feWnQAgK3R18rWWfh1kSwDuycEyLVC
LzkbV7McJHA+xoTeImWdfmEI+GkzD3n6zaJWC8u/x4lY5Y044vQTXcdqYn8r
7ZyoMUOKy3VGmGsnR+VFwLVhwwdDJ8ZHzFQAOLsf0jbJ06aMlcRSVqvJE4c+
fAIMSO90zrtN2I+N8maNfEdrOBCpiNuhhadbvO/mbx4KawBACKUUvUV2iqVQ
0cJFYcB3JiL8wd3DOjUWydoKfGsPDHMSFt2OnPps3vZiD94iKIOO3idUSd+B
vaKW30Iv2TBYt0njfJnTCCCqRkKAsuUvqc4gpb+PiJIeHetQn9E0EzcNuXrd
BM7J1Dgpk0I7bRv0HhoYk4MGFPjARxLcBZD1q002Tsfy4jdgkwnl+YVvLbag
hVYx7IWyuQ6OS6jrTFpKfWY2+4hhhV6zestr2Ye9W4etDugn1tRy6l+E76C2
mgJNyZZuMbnew0XMWztjkhV8/W/SECsc25607pyJjzRxITBrdUchFoZLh5aI
LpVg/OU5iOqjpRcD1zwIn+wShfF8SpL+QhSAozO9V37ohG8hRhkn9N0reg+m
HT1XFldQU5JEjcimluFcQh2XF/jLByPRx734+5e1dfv324q7O/jCEngdDgnO
/dq/frV1VPbwiUL5wEofPcFyfMr+8CGrb5p3O2PnbpMJUqTIE36QG0RwhoUQ
NmZxB0GBg8/q4Ty/kH49Sa3h1nXiiF0k/+/L5nFC5vQC9YQ2vZy2fd4L2LKB
+femjGinJhOHsUS4sxZr9ftHCo2dBpUZK8rm4r38pb6RKaum6mR+GuxKxeCn
5KAEoSLmrZQeFSIEex2N8htXbF/dbkHEhBw/a8Jc4YamuPfXmmCmghgBzhdW
OwoP8RyJpqkl3YOONinb2UU29hsYyhArGhZTL16cY1ibIVMeIQQMh6bgTYZU
74aQqzge0xNcmuYuSlhcJocmBykITrc6B9M6yPbTmma4KLyp6l1juQdjaDnH
mBYDLgKjZ1bUsFY7DsnrDm4F+/2/cDRcCviF8YMOki5XWXWRHeX4d3ocWcWi
RTYlWSwdA+HOaY73YmtLAkQYi1Vt780+GKcDxAn75QLUeVsVU9wwmNviAlgD
wfdE1bPGEK7ApGqmTZRWZH7ZmP/znNUQ0dY0Xs9T7mx/fec7VAaC5x4Srrew
RYUsBXz/e5MbNGqHzFsp8YWpkPSE9EI8ZCyqdF5pxEP/6i37/SLdaECshl+S
egNkUMN6GLXYyWP0HS5l+0sN6PWkmdJ+gP6dEFtWzDUdVZoP93EDpLzkwJl7
d6AC/GeOf/5osO29wSzaHyxorcyalxQbl/xHWiw1Kn7Q90zLjKiapfkEWnb0
4aCWLu63Ckm+B9UkcqvtjRla8qNZW58fEWBkiFC4YzerXVjtKT0BDPgiXHsq
snVQoe5L0Irbqki/ZYHmGR7sJzVGoMzXVTPci1FZkkxaz4m7s59EtnDUaCP7
3kYOcSD7vjp18MuOFQKlePqSG9+B2zIeFgpV+mxF5quqBsoUnxvgnjWS4XIG
UgcslKa1AxbUfNcBMOH55cYJ/KztFPOYHD7/Nyx1zDAe5aerSR6nIR5fXJIx
l51TEWCFA9uu8AIpDUd+grtZUTNoK2zJUhA8U+guszC9D0NIDBs9QjEDt719
IrBgU8/Tm9ICPqHXHQXV0s2munx8qjl3JHZ+sJlzXWuVTD3JxLwMk4l+EiL+
YXFtswd1XHPd7WbPUDBcG1Ksm47TLbaqnMRcuv/GEsRzSkqxUyFJfsQCxo+i
hDQq4tkGhYnueAS8k/8lPF4hU8gALHKNZiQ5EDKcsURYxrRtgD3iED+IY7y0
KxWpyVdHtkZIqkOq9X01yoiiMNxOSOky09N1YETJNnLGYTGa/MMZsJVnJxLO
stbXzXxAxlVxUjTqIM58h3gPe0L4fe3XtLaQptRb9AVpvePM+h0jn0+2LVoY
nQWV6ZPzdmlOSGBLRtAnrG55VjlKmJomwsAoOMn7GWkdawjFJcvlbx3EdF1W
OX68e94qg/seochpj5WKM52AFeeai88pYTqnIuCudeLZ+P0qiJG3dcotPgLA
gS+UkMzOG2aKsHtKUOOVvxwwz4aOhsEReZFnjEF2CUT8JzrcuZkVh0q/0kBo
fQEnxtkzwf3ZL+00En0NN4SGfyJHlV9del3GaPr84haYz5v8NF6CFDPlzsBP
XU/19ASz6agvLjjEtvC+ZK7KsV3Kz392b+SpIFgVauH2jOLDOfx0VjEdYnMD
wwVUH3Qch9W4xsHXxO9XnAlXJHIidVeKpkY086Rg832DCZOrUBv+pQQeQHWH
1yCa11PoR9InbrEsmmOpLbv8wTvGwp05OALy2/Uu+cwka1ppSiLz+hBvAeVN
f1fc9embErt/sMMO+IQoEAireSsWB5LqLyNn2oa1F1uKQTY21lgX288CMTBe
MjDVN8w7bFLPWAIxPO5ZUTpSJDE1K81QdFZiHUoX9COzEuibcUhJkq3np6kK
IDgpHhPBFTLT6bG3Qyyu5ntC7olmz+eY4EIGi8fdGiFkqg7JUAbt7NCCjrpG
iPUw69BqD1XWw9U5BxTgQwgdvCKrv8ux2PjuLIxKnFJMy01AHYaw/gUTD3Xs
qx5t4hVuLd+TLoy9Ul42mVDzkJ5Drr18BcqQm5MSC5TN8hIu4nER0f+FE52c
cDU5azzzd871JN0GND58t3aRy2Tr3mWNU15dYiz/FilWbqxhe5k+5RizJnzW
VQnwuNTReUphwhJwr0znUYQcAqb+P9c2bSp+8ar70SWW53cZ6N2uHmHHKB/q
CTSdet87pa1NoApYfxNZHwx2TE/ZgFcLKMDP7cbcemvnQ2P/64jpJ5lsij04
VQb62/w8bPA64jgzeH35RAyk9EjaiSS/+eFV20DjK6llUqZZHBeMsg2ubdYD
Zh0LAkhAmqzhyzWRtRFJzMet5nrPXW4Fn1Zbqa7ukzeBlaJ3ZRiVgXQfEB+P
SiglZm5Q4KJTCmeLIkABeB6/sgn5KoEiNfGZ9x35iwJRYAgZXnyvNw094qZQ
rHz01u84FRFp7O93rjO6JX1wbt4PBAfO6+8+yNg/aT1CIhiqDsaKvz4ZP1d9
JUqNSbR8532bLxETaklLO5g3U3NrGcqPvuq6bcKKEhHMhtC+BDSmntEEjvwu
ioOEopKlGaJ91bS7w0+n2IQE6lYNtX+R5UVbfNjmU6sTjgBU5/F/tZAyzut1
bYwZ4tYWagE2e7u6e9/tOSyuWJyn3vD0NL86Lb2YZJpYBk//urm8+v34icXc
KC4PL6vbAamSCouhsPQrS+e3RbuZWKKbS5d3wOor+BvAPg2g014Z/YCAOiUh
Bu8+TZxmOJYLMUVqVNdaEJzOdBUlF8MaGLoou3Pl9tuCRZZNEflj2Jc4DVhm
hl3TBrjRDxAnB7rbMaL+X4bdFqt1E4hiKky+4pD9kCi641bn7iskGViiIsim
IYKZhR6mf6xgFYJeYUSxWFyXIL94v333EZff2IhvGLY4gVgceCxtI2TR/Mhy
F66mpY7m/Nux0Sw5sAwAMit4Fzn/KomekBWrxBueRced4mR0QSEKQKLt0PNS
Q45WWT3+RLxBBFEWyH+a36IJf5f+V011KgwSU9tSvbqWWrqwRTjjMO+kFMyi
CF5ptgeVbpn5ap+TJu8NQvK7P3qFra3Lt7G4Koqqpx+tJJJkNYLt4TlPGgSj
zRMyQof1cJ3/n59ss6rwDE80+9yO1ql1Y3pL++GgD/lTv9mjw8dGowkVmJdb
tcwzdXdjYkXNb/NzYFXsTyarTCrFrGMbDTzaXvpV+/9UH6/OkXjlbkkDE95E
QdUppkWzLZRD+ToNJxnmvo6PtVPRHCsjcrAZKIshFD7xlxjjSVM3yLuIKToF
gZ8ebqdcRFfIESsjvwxV6cWf1eqPajkoKgQuPxRhXH6B36wzEVHMl4nyHWUY
2l7dsOtPOMnsMhVcov0fXRaUq9icEfYobtL3A1bWgeSzywzpYNDo1G8D3dn4
Q78h6TPR8D5W6Ywg9CYNaCXInDZ4dfpvHBHq+QO/ecO8Wi3P4RkinC+ZL7qm
5Ah0AWYaKSZUQ7W3GYsqDR/g0oZ35MwmRw2nQCCqA8JhwDEwi3WShYkTsjxg
yYarDGZPZvUn25xLCX+zXGWmkuE8Kpc02AsBl38KbOpK3HTwo1xYcFYdfzRc
7hOwf1ZHbXx4E269BqObTsJhQzONbcNAcw/V6Vv0VlRQxzdT1inmcv8ja0rQ
YSTZCVLEOfP1rsFLZUqkemgpsoDdiJxwuE1P82wOnCggXW5rr3Cgy0MBFk/o
wbKUyAeH+Vo1FJxxRy3PeDflRobxImzwnjTkvMqhGSvnUsEUE/+TArypP29O
PhpmPCheBVOxS2DC1MTa7x1XKpuJ7zxB8Ygg9BkMEajXYzfU8/lGJfofdTBs
RLJBkG/y6iwEEpbvXsErwtigEkcc0hp+rmmf5SE0JgewzfU5jtvuAAT3j2Fx
E3vbVBnZy1OTh5Nz5NDEkezVjofqToQlKxg8KQ4pHY0pSr1EeKOK6ajH/ycD
azM4wber4wIDAV69NCTTh4fqV43FaxDzzdvzqL6xOywFtnupsJEi3LslN4TA
7HGj749aBiOTFWGjqliS0Ngp/z0xLGXJjkvxeSOTk71vzJs2SUtAdaXIFRu7
mtO7CYl8wLIki7OC0MMFXhNWttSNKrgCwO4t0eYbq08mydAQkHHO12SlN/tS
qWI8ZEau2n2oUDMPFB1xlOdKChqEc6IGLfGYXsoThKEktBpAPJkmeuw2JccG
Y+ugkgAmjVtPklb6XA3S29BFLIbBjcDv1U+S5Ba5omUIwvnXV5bPeV3rDLwV
86UeER5SYUHovrq9Y7z8UOSwcjUlde6yriKIDZ0kwVM6Oooqw+VOEy3ymRTQ
sT1+dkiyr3qkCOeSk690zW7lYr+Bt4dt63veIeEHy98tsZ7+5W5A8WIYUyMe
E12l67ns+lXuVIOounWbzbKa0YryM1kdKmM2JTBqtTXiGdt8QY+EX6CSnKrN
j4CmWkGOIMdd8xsDvaLfy2koIIq7rrKVa/jWh+TK0zXxcm0QOnNFdr04p34p
tdsaixBmr0fitS4J5CGr4fKfF54rstDPsDu/A1TcJSQeFTcfDbkh9c64pS7M
FBLQd28SNnxwjwMaUPyRYfs0Ct3PBqusPhGY3BtEaaMVUL973GCL5XzdqRBL
hp457sB16caSat6hBfnNLPRw2sotCmk3YJG/JjcVKCsu4r4BBSz2cTzyvSCf
3fY5Pt4+oQ0OkJzcMqIuL3xbVLvNkPSVPz27zus340/q3KntdLIMREu3w18J
sArRusARdgaD+PfieUuCElXBqClMI82Ukd6mcRGn4R4IPoyZyUS0ZwuvXjS3
1l+RkHXyRYuFOedQKwf10uNHamkT28u/xWHYIMQt7tV3f4r4tnIGl6Wa7XvN
z9uxE0Sfc214x/cBzxqET556ec0+sVxfhxCF/CmclOZdB5FIAAUdZt2eo4hP
sqIhMcIgI86UG3Vs5zAGQuMl5qL1bXMS8lnyT1R51HNzmqPwLNsUo6iDDM08
XZ1hRWwRJ4Af6AY7y4zPYJPq+5vnZlr7CIfJcHq2cx5Pk9lV/7KceW6VdMaj
ymd8bmoEKvjWFMjt75izvx94vkOlopXP4YsI/T9XF67cVzfPWozPQhlO2rEl
UR++wHj2Tqqq96WAvlKs6Lh0wKxNqp0UmKI7/NBbpuCfGjBiizIUP3CUoUSV
ZldSxk76fKNB6Co1DFS4e1uX+cwEPLcGWemzXoriRcBkmsqdTaGptVNCPVW1
sDNoRjt0g4jmdp2rFfjABZWhqa3Oc1YSXencwNh+iu20LGF/j5ffdK/RBU90
U2g5Uw2CSNGyxAkMVg9rnZnr3tevSK4FeX7qBtZwpsfnLmU7XxP9IxnKLSMd
aeqHyJFyTYQlJNATr8/Z1Avg2l7itsNMniaKdS9SBMw6XyDG3cogK2VqJzFy
xc+FWY6bjEvVaTDDu6026Q/SWPn8HSWgMEGh0ZkC7AlDIouT6CMYdnvOuK5k
Danawg1CWKw+fuZ9UIvJkqEyuvT7LJcwqnVOSXeJF2E3v3ISVGapvHq7QZEf
ZxhQJ5xPz+177Q+tvymm8OMtQZGjhFZ9ItguehoiPg7DzZBkwn2xbwQkauzt
Xf6N3Zbz+9NY5V9nmJYVrCMbsKlWHQE8g72mk37HCmyJsaweZikzzJeXxTu2
bgyBibmzySNvsKCBWNL6ukr29S7vS0dOsI2wfJQQRFMKjyn7gS5sSha/S1Zv
mR53OXvOXsm8d+7Wv0ndQp8J9moXCEkgt3w5iRJFvc8Zf1JC3+7fx1B9OVpN
1YDQEL8VeO3dlBLaLnfGVUA4JVZdCanlMBYj3/0/aMH97i7IirDUppBmh+4z
1NdD4CCsspQPOdqvgvoO/hp3NA2CVGoBv5q7aOzEnE86iwX2Yhu5oMLGZr+c
+261+nExzlZDMS2qYRFk0eJhWKVCok+cFG5Q9RttoqxBbT6yDsl3NKLfSGYe
wGINf1O1VUqlmt4WTFau2bolMiI6b5Q2et5M5ye7OMgo9yS3QKOW6/CfRa7u
MgOuw73TGW6dQ+FfukAQ5FZRDXjAy7L6WvHrsYRShodD2yiq/Jvlw1axpdNU
c+2bILojJJ8haY+53OItvfdN5sQwZ84VdqAtJvqd2h5A1+GROjVzpjdg8iBc
9az7hrg1tTq3ZLw5zNm8/eqtKWaHql3aQ5TzvauguV8bw/c0E/baOOilQoAK
0ssOiy7abRlErP+ungm4K7Zqa8N93MO5zfYqeCGcW2WKQ/ge4BbBCrFSCjNR
cnmGfmzBTZsiKvolOu7Hg3sACYpW9q5t7EsnECWZDwm9EbI+pP/oM98VJBfi
+gaHsFwWO/rP/uCQam9yi2PoBSQENbJMcX4dPAs8JMEVt1Ck4bvRfFxulD35
UilaHV6YkIZY2h0lJzP1nZPzm+L3yQlb4zBij6D2k2e4k0498Y1BImLYqsPZ
2stGgTxmnfRNX6Q/kaJIlNeTNKQou5+nav1y3MCiovY0d0xYJTQTn9oq46uB
y1P0eL7BDEEoecVW3sjKSntcUAuHc757FZoPXVqht5z2mFFipQn226P8Fw1x
qrLe+iEg8UA5tBLNtFApnaLm6Tvr5XGno8BkziNfgeotZT49rSxPzZXqoqUq
qzCllBD3HGRT5rGUXP2XhrvvyqZm739SAAy3P0gLyi3+ERPN6QAqraePS2g4
GBNG+3SGnnmDrTVDcTucX/hgxMkNoDT3q7K8xVxNTryi7bsgLZvUu9w8sach
YCYg5xoOpjQ/i+i9CPB9bu37geqIfzVG6axrd4CvAuUk+aH6wHrAah+84/sS
XypY1gc+jNA06Aqa8824V2DtqTRkLKhU5AW+LEQEFxEsa7OOqOvs29Y596u9
M5GK/JTkKXmSquu6rauI2qYZUvx1YfYWzlk68R4qVFufUVx1cA/LutedM5fo
pG1orZGTvoUlIzwv4tjJp40TjiLZrRU5/QxLB7TDBbEkkF/i3Anl1SSvyfh5
Ctxpf/JoFcXeS9T+VO/0R9JxbkwrQkYWnHUKw05qVnyoL432Df6N9pdXGEyA
D7sdLdgN5p23WcvhAuaEytE0WPTrf9Dp9EiiT61Lb3wZPMzgRNZtYrto31qO
/CHBV4/hNBNODTOO1HjnuMIKRI7YHnLypw+e18vSogd4ClZseANijXWW16oE
5/NH6L0LuI5at7SA8EuZh3q7aWOLsL5mx4YXUSI8Z9V2m7g1FiW5yNMddO44
q8mLHK9Ti5xPtdwFgGJ+tXX9YxXMFJ6c2Q+HEou4BJb6vYpWmssU5SexIoYw
k/32PcwvpjKolBm9d2kwhCFRMeJhM7v9aeEOQdqGqEoiE4MOqKiJ6pG586BJ
U6o4XWieoymTHJyKCyyAU36WMN4zVqCAPGmKZOsm1OvAV02yG5nOEu77DyAP
Cz9qzJTbb0hKWQzBEdO4FYZaIhJac8od/ngIchuRbRdnnOEKKZ1+IWGqd0QZ
w0jNil7qt/LmUe0z66TFAXtgAFpbreCHUOC54g5vLHI77qWVhABvVGXvDRax
3OM1KTIwUV/y0MDLRnvsjzncHAknSJ177D2PoXRGOI8ozw5ZlB3DU9Ahk0fB
ytX7ESCe/ZbCmFGU4V6LTK3aLlCzymLjsF1huO3p0PwJnh7EQWYkHGhMMCjS
DPOVNnmlaV91j/bPjCKyKGkDyWax1qmsaQacVVkoDxihfzV/EgivOUT+3dM2
jbjCmMs8SqOynjF38oYZVJYx4ZY0p9FpYV/M8TAZQ2t6u9qK07GTQCsJ0oop
UfNyOC/bGWdXRSCFxDwgfC5JysJ2D9Y37bRDGlvOe2EMlFsKr6SjZqedbWip
4ZbbRmBQ5lXwVcV0sfWjLBYZZLNU8bfczWbZe2sJBoiPUkpDmukCM34XMoUN
c8xFdY8e1BZRu9WvvJyl0i9ZxTCWqG0r8YXy3mVccfeUoPN2boVNJCp1qFEe
bTGgkWANahUsRfr5yoZIEHix+zniDEmx9bWZCsTfLSNLPrhb7snZEgEnfXeM
QhseJONe+vjRg0Qg/ojHlZhSdFXvzCms5txKLehs2/3Fu4uMz5i6SVix8sX+
03bvXJobGrGE0YKFXX/i418POosenWhzYu82kLpcIDt7bESrjXLLRMI3JTbC
OcDJCEelTjgTUH0QFfFBwM4zU4RHoeH3X6tEsizkdyo/L2IhNpTRMXDikHCy
VicafGpxk1gvtLmrt/CheclX++0lk004Uop72wD+gBixzSykOZ8d2U5mPOLm
G3xh+I/TP2MiA/jOzOFEyh/vir4oChbWizmRCXiYQH4zBCXyFBo1H+CvbUEn
QxQWWIvqF8a5HaRh3CNOL5Sq4WfV7t344/9PROw6Nv2xQU8fhnLHFrHhRdxa
S+7EDY6Y6SQdr6vhPc4NZBsunTxFy/Zi0AFoLm2rBrag03DNYh+Lfgu9OC3g
youhhQbFI6yeWLZZ68SbAsGkQbqapeuu4r7A/tyyasK7D2ZOaTuDHm02wJxN
ySZ+h4chRwwruZDHVCRTJQvjP2D5OjrRIVYeDIlhkj2EpBVH6uiFg5Se2+cG
VfWPHo6sjSbo7IASuqCSX33rjQD1DM5LGg/Khr39nZuRM8yPoksOXll3jTVh
B+aiYNb0sNO4yJ6NnsCdjsIEFAsd7jU7Wa9t8mJ/xBpdeK+ePRmSwyv702KV
BlSkeIhlR6x2o6MFfgwg3L/6fYpJ3RMiSpL3ZOhEG5UWDXR9usLlu0yIBEo5
vFNuKGToOqvhotdSCaCfVFtGVuBaCY1bHX12GV1NeHnVuz7yxFkA2oO+ak4t
YjlgYUPjf7fpovjkY6ar1JuwaL7di6LJRNLWrd4XJMO2l36gXkqp67nNsS/c
/VwOLetQ5ii1LFmCamKaUfCR7rXvelBklFCBo7OnoqOxqiXqi89Dw6CTODL0
k1i6p9lFbkAt3UGjXlGWtLdKNfWBDSw9qrLPPuebJyHzwT+FhUu3hjYiWvXO
n1X2BMTTOo/gy0GJcz2u4FZIYZbRgUJiMpk/AsTB1QFrS8/5+jGWhoJXf3X1
phtPJy3nvsQcaFjYCVj5TiF9tq4QI18TSaCgUryPmOJiNKibFDcHNfp4h8Ck
sRh8xbs+DsLD44ZTe9rS1/ktryvKq+935nd16GelixyDrZf9WBd3z1mriuvO
KeH1wbYu61PLBlHHDzauebj9YmshRTPLQrXkX719QjJXDo5wvoTdPXDNUQcq
VaVwW7L7QB722nVtS9jXPQp3gEI7aouWz/4293vT/0BENgogDb5E+Il4NzC+
6B4JSn34SfSUhO6LUyxb6ishJjkdeLcqWuNOeYZtV/WNe/ddn0xea437u8ag
IktLck8uyoloBZvP1/1hfQJqHhylpMwczr2bSNfgYnKrwI3qDVAhPH0YaZYU
uwA5I64f/L1NmXua5S3H4QaipwDpBjK1WdTjdzSNlvAhDihpjgjuCQcfn9FD
hzQ+k5EXOoeIS47l4CBAALZ47tUpN3T9PSS6AKx1VCFJjzgDAHvQp0SsGzYd
n0uqUdXFyLC1YjPJ562M9tXcFkaslUwnU7DxBgxXfC+ZClZ05/YEtWNmJZZK
uHBog8oVioLltqMRGt1X9iNmexHUB+C88NSYgA0K0IIxIgWGThYbYVuSHcLW
ekMjMrxhstF+kn4jZqpbLXqJ+dIKaspw9ybKp/G40jXgww4Jnr6csqMSUMvb
yfvY8LP0RmTjQTX0PE3auVgEV9a+wkgk5P2aLirpgqFhC0PiCHwb2p71FUhT
CBGQgxV7XX06OcmxBhxTiDzsAtT+4eicnh0yKnLIP58EEOY8/uiC6x8JmbVF
dxHh26Tjej9s+x1s3iU3T5c7IAnFqiFUfCB0O8KVJnHU9dLU2ZRsheVcuOYN
bj1qDFSjqdkzgFxZx0Ff+/AqZ/kR3Q4erqAio+Aq7zuFQtKwSu7H22IsS+aY
cFEJjCc88CRtT1t4CMGWcyzSQREUvBM3hhH20DOYWheVaftQAWHzIwgmPHqj
q5DgMqtHYqv2VR82b98wNCulmrKFtwUgdUB51efbXUxl/gswOuuS7hHvdl9G
C/BMqmJ8Womv5tOqBvgjBLkc8DoKxVh8pa83Q5o4OdO33658ZKKe/hj/H2qA
UB5zGEr0B1Oz/F93clgt79KZnfXrXBImma2dTdPS5oGCxOUW0YVzCp6DTTpy
rJpaaHVSG+yz28iZIerKuRMijDMSJ5vENfRalCjp64PlSCkOASKErrJneJl0
Pq85r9OZx5s3qijap0Kfy8edVtHvWKQ9FTBiMgwma3wI/Wl0hHx7ylAErkGP
MtKayxQHIpfxT6iL+ga/BqOdjMk2dlfLo6o2hEcaCCHeawZ4N+e9u0DlcFH4
f6N5bZLLQ3MVQc6R0OHsC/gfDA6Uuk2Q9VFts2QprAJwUk37VXaB5o1ECLsD
pV6t8g+P0DuLcAcflCxvKlbIs29EhEXUPo6XgMeqZA6S1dQxg2+FTLlO2Ql9
K6ij9zcUaHsg2A8nNanAdQpnRVYPSYmPE6OdyB+Q88RQZIKB5jLDD+mAvavr
qLRVn7Co2t5Xklg6WHMabTCN8b8HSPqadVHy2YfwuXnxPkzy2NHC68TKHexs
0UWe/lxfhuQZTmkjuTnpNimMiYXeHWkxVobjOo4l03r1VKgnZKmj62WzqM2N
u9b7cmvEWEuD2+hFK9Zjzyh1SnIbcoT+uwzZIhA2C+rwq6hFsRuQyGSmpSH8
hvq2lQTLNJb/b2YXgnluIXyCQ7D7WXxb602X/4sGGParjZCQYXPETDbaZFfu
BLy958CBHQElN161T2VmkTtnloc3VMUA4sQz7VVd//GAen4C9Ah/vdrTSQfm
09X8EImnCz2DqHzUds08Z2emJGC4D00Nw3nSbuGW3JTyazu6dEHcmsTOyHfQ
0LfEGRlTGGvwPTNmWLkSjFX3m7EuiQfPOHWr8rseW5CAz4A3iTMKjg56xC3i
8glw7KY3K1pXTPKLzPM/Om9u4J000MCe+oVGZitftTBlh+ZuMQoQekqz4B4q
FScjPCA3NmynEzGbl/trjYKQi3z5ZlyAdf/SBA0omXHC1B1c8I4mpCuRMl9e
Lq4rluwcGtLBtAQc3cfmObQcIOBmh1/5ZfKW0glC5ri/L9U6vd+KKAqD0l49
Zo5a1WIX5IlXKrerjla3K6k5ZjkhVGZtue/Of7qwDys3eh8vOiSE0Uhmal+j
LD2+X+eswk4+N1RU0xQapull9XefwNJUcOYJXiX1nG/zNfhLW13UEa1EZgKu
HdVuZHpSk/8uPF3llyd1u/aIuW4DdEwsC1LuKAWv/5DbE3VYk1yFdLvdEZjs
vgWkYMC4lm9KVqS2vkcvg2blY3EBzgZk83YugXFtWUqqrZ/zOuCCmbEmgixA
N2d/mR1M8MWj2v/JPVZiGSK75FFRO7+o7oOUphTgRoH878ZKmbzgHCb5c1nT
NPhK61KlCh0wrlvYWMEe1S0NqZHPrjg1L2WSJDnKFSB57nBFg/xkRBLJB95f
Dm7/OOf/XKZAKZs8wWFTqQvxvKUQT9D+aRvjE53hPuIBbRw2YRmp2xyCtlkb
jQD5knU4GUJwv1fUEd+QeajdvfuT8isnyQQhIScy9r10b4AxU+bgezDFmnz+
1WKCn9oeU5zBET1WF+TMA2nEhDtyvwHfzc3E1RW/8FnSPlCukowB7xujsbeZ
oBFg04sgCKZyC6F59G0y/7ijDqGGdqFJJl2f9tjNw7sX0bGsEZCuZn2Ncdu3
SMhTECi5XB/ztZmG3l7lQsqm6VH9pPbE65Wphwq/HfNwlEgnag/l/oQ3xbVY
kSOeCTORl+Uqd42UmDVqGBsNblmgEg+eZfOInJErrCQXKCzv5iSd7ilWU0zb
mriRNVIhFJxiCdVNx0PLOHSExJo5y3ZSfgyslXRwyLeXbK2inYnAnXWrzfwC
aEjA+oIFPQEBj/ATu4XmLS83eDs8e9Lm5PkUqE02uA3zdlu5QLedp7RppDW0
eT9EycBoF3VQFn5re+yFMxU2gOMAbeGsR9oNHr/5vJQfqrkMxkwA9B41AHyV
+7oNE9XDOhKwBIkno6O97YbsTT5O5Ynj95f+1WB/5Tk1Y+U9ZRIktRfuqrL2
tKryXa1Ttg75b3ZhoIJWWUm3Hz5Gifd3sVy2gcmqLggkeXPvaE35YoP+3xl/
HJK0sRiuTNQdR8b9H6yb1ilbzkFNhpYp7NB5BVsY0c2wwWu1i/Wwd0LNYsng
yF9HXX96Qrvs6MSES+ygK2No7QzdEUdiMsemyarpCXxnLLAKGVzFDhBunH7D
ON5AH8bOd4hc6rkldIPwKMMM3xHSvI0fXRW2ry2cxwVFd2m9ujAODB4eUAkI
Bx/prV2oJLguE1IFS5FVxOV3tqnAGfrhXcilmeMvdLK9Vgogg3EaKiK9twW7
KCVJtlZ4AlggUH3FX16aTHrw9OeWUQ8gffdtVq5FQsM8J3GgJm4klMqdXV0Y
U43sfAiTUcfSrYDvBUlmgLHQTNpzSMBTIfE1m9IlV85eLM0BRTdxJcT6DmYF
JENrA5McHjCgnpdNXlQ2srJ72Yuj1NQfa7OWespew+XcXlWCprI77EM0p4WK
RsL0i5BRmoIRA8CEmHjnBiqcZ6xv7E7cDVQgAJBkVeG9vN1zwHPYYQkGOHz3
7p2HyCn24VIQZRiRR3O2GBEfk2k6okvxNjf36kmR32eBg7HxSJcx0+P/ftsi
IQ7oGoTUJg5+fHL+C2VuZjpXk3mwF9tS2+GCsNiCOjUcm9Qq81Bl76hAjZ9U
tV5I33VisD/YugarBMynOVNgdxbhJIEJPFWTqw/68jr1F1S4NlhPXRDvoJ5m
Ue17ScYcEBU5F/qlAjqWadDSxtc9OVa65bTzxdyTcAiWg893Mr41CLtnebdp
6Wppvpgi67DPMAfbTzh5G8ieDhdETGIPtdK+Jw+xNkr15jB8/HYYy9xI/sfH
cnSjHdkgo48v+cpMKyI8RyCxRMYYarMQXE58rPIdsZgyMWyqmHdl4AEyCuxV
s3Y/AcMVV5zKMGfoLamhMbekv+FQAPx3p+NlLj+jMXXgEaXbvaGDuroJLaiY
BmUpGwPtwBp/XteuQY8UPXVtheU2Q6siHxxWoRyAi/Pbr92aDMHfoDvkHHJW
e6nHVuSR5hd1HVvWsu5ecWDyny8d97SmGaJqucE6GRk+OzsCWUbyOUXbFV9u
0n+PIItA6t4ibMHy2ZoPFqhkdn41FqG9ORD7pUJzTedIkxtpVuk+R2NbzhXy
+q2Dkti7lyb55wBc4eKar+7I51X8G8DvUbd+kYn5a63kQR1p6PHveXLYelJv
TL+jp0q1cHJi88Y0a8rNmG+TSOuGNgd83NXZfJNZFGMyJ1UVlgPnPJoPH6hU
MfDzwLs4dXiaYEaSM05T3DGjTEE38TPlld8aCyBeLAAtsOZa3xXVVuQ+knIR
+0j+8AlMZyGrE56DtOGMwepPlTssqzliHw0J6asg/+9/UGSJoQhwM8XuALs5
LUwd3vtyTkYlLcMd4O7uPiUfxxTLVuursyzNWs65bhONVWkL3ZNvbg/L7EtZ
lhCN9YzlxWdZ/7pDtFSOuMYAxtH3JIu3MU5eO4n57uApVGFhDqhR19c9YAbB
LzFDniEv6ONgzMjKgcXWJbqhUWbAp9i3JA52I5flqVJ+HU+Mx9vZ18vUSKnf
ubZpHLoDVqoHobxRvsov57I3hGd42eJjdxFYWpgVsmTW8oqIYy7nfcGqxYOG
oYtLS6CRpgP15ibgyFrLTr0ZXNoHxOU2ikLkEOOv/b+1z31dCaOwBr1s3KBP
QyeNm4jtLNYIb1XQ/GoplEjNK6MiKc/u5dJ6lguLK6EFXbf7SvA1QGUPiv2T
2Y5Fad9mriRizmeQPZCt4AuyjbOeyqfnWk08ItuQZhiUZJLJqoRjpCbg/Sde
pjX5YJnqykPpS6z684o/N8GDVUMQ75CuVlTTdvkZ23s3irWnNCVW/CvxkmZU
m+ARMOFGF53ZYS+srBnp+EejXnx0yiYAqUY3nstWjcWvfHCOw4cGQw/GQviD
N5t/d8DJFKKXr3wL0EnE2x5vjc5kcuA06Z7HBYqer4FM3/raXKa/grE6Sv2L
x3VJwH4vC4awqEH7cLYcaswAcbfuHuMb+d0eGB3RMi2ZiJp5ZKBP6ucw0/xJ
GKWYaAB/mjB4zmGy06IzvYohrHHLRFoZLBadppyiE+y79bR2tVWLyMxJ4F6n
uk2lp+A6D30eZGG1d8e7/Mp4CMj4wU1sKI6qDxs7w+uHcCF6R8DAZY0enGEI
YYDncmmqVisMuMrh+cCTyw6YZboZpcz2obhZV9lYOVJFz+V6C6NPBJtqm0q7
XvSdqHNwE19bGkafGdS5Zy1pYG+cGNWKWc4EhD+SE3y5RvvjINd8pSZDL8oe
2rD88Y0RTSu2XtkPMeEJDBorYnq+dgSYkhg7fiyDWj5UJJKKxaYoVjK1hIc0
lardRj9Sgn1FovrkXaOIj1BtysaKVEokQMZdReu9D8PrzXQ5kXJIzT3cyz9V
SnLzMSWe9HEpnXRcUwmoB6UM4kQqkj11T3ZqCIVTTyi2BNuEN1qJvJsvbzLN
12+zs9hTric76JQW4JGAh2nIOvpCYrxg89F5Chq4DqhYYF6INRJCojG5ig11
d+eDbfy6pLsQ10vIjM/cD4u49DengQD63bdGFj91Gyd92kORtNso9UBkK7O/
MQFoH9tJWVk4aREp3ajgXvLfs1HNAdm5ow3ZEg++BHT7WLryrriWYLi6E8D3
FcZmP1gQn5IAQ7Q08ivUhJ8fd7/51pNSseZQAA3t1NnUA5hR0tTNCnKYK+cl
LQrAbfeap1N5agdKrci77HJHTiStNGM458oaUGFRCf6iB+Jtd763qkiTvHnK
UcI3Lh3RZrfF3EVv5Lvai7hBvXLJn8ZnP18908c+fAVA3Q1aogLLNH2H5qOK
QOVJc/bYv0PmWx3hV3zR+HzyhpGvBAn9zmIkluqs8hxqYTduSYkKaLwAiOtS
ue3NwuMFIcgJEux1R78tOdZz54BwSunYNm3grlmOj6SqhSclAkC0TqBDDKTR
y6wfpTStU+3TO/UAW474uuunZLB7cSswG/uQKUPBSHc/ps48EhAOjs9BfMpp
kpQWLp6o18lQZuKDLbjV9U5NqjNO0/+kCClfgiwAHAdnFUjORWNxrnObT7bD
xYFyayR0FwvycaZmxbPPxI3T7Yg9fmZHY7HkhF3mLM2wD1ulGBa73/0BsMGM
3jar3nYMSYW8PB0FzYHgqApM4i/gH8vi55dFB4STKBGgd+cC4zxsi365I15o
lC4R/FmsBI7VIS4JeKaLdF7C6T5A5fBJpGEY1+sF8fOZgYPrOUBA+iC3V4Z4
PP+N3Na288zxEz2d6kmA/rYuPPLrunrP7XB3uIaN0iXoYhA7cg/racM2ECiG
qDmqpDzbnFe9cI2iAILvkgG360q0onwQpSQeimzpMUn7F3UcKgAKO+RyrPK0
liq6pHlMV4NHP5RML7p6XuT4uiaRFSavPFOWUzF79yn8eNcMmMxhyoW0rCYU
zVusByW4SuM4D9Cj2UrFyJOznF1YLWmtvY+hnbVi6GYV1v+pcBeFIAINaJAF
na01PL7kBXxQDl6Zq00650OujbbUfvrtD+tphenoYYJF0Evx4vFkbSkTzdZi
oZgrw+igSgSvqiKTGwTbbsvhCSxaG471rUCP2qFywfHmOG68ihdL5KZObD5a
2iZzrBDsHO1I7F2MdLihlWUyhIGybBqKNnev4ZpCSybhPCi1dwhnqrKWVOAe
5NXCKzEmjn6kboJ71lSMfvsC4K2he78w2NCR+/4eat3SLnfFg0e1jtACkFuT
BQHzml2V/Dnk1jvXcso859aB/F1/b1Lep2Uu9OICRQUEEY02TyfGCzNwL/nu
7aGnaQTL78RWaeKa18coJM8dO2PLfGwdqG8OeQ6FXFhKDszU7uzorNJrwZTa
BgdC1wgc6M2Faxi20DO20Z7qWpGEwEdC93O+/KK9HiVdQ8lkB5EEz+Ojlxyq
62AIvvwp1o00yS4bX/YRd2HhPNCfhc0PAEcP+yKjmN3QPnh2Yo7LOxCbrTo1
TXB3MPE7rpfEmDoG8CWZKqsOP0/pZEdGxXJBGkv/VJ9/e1EYUG8XvAK5wK5X
4WbS6bCoPNwA59yb253qQBbsunSu4zCEA4384hIYEQR5l9kFPbJRpddNedOZ
/KzXQDQVgJwqSJ8Xx5uAH39doaQM6vu9P75FRycWsVSXGB9WYvnzA2G7aa/K
IMD5fd+SOXmmxIb+i6UrKF3UGHwEBCWqjsRNd79gHhGC2sHveNTYB/xjNtfe
hqVJzF8k6rxHzc0nBuk5IhDL26xHTcQ/Dyna+zOvNM+JhapkNkLoR9zcRN2d
GYWM0D7fjpOydxx76hsxTVXf0VZWpIbt2KEcA1L+d15jFXkfcsu4WG+yowSd
iRPZUoSTxQj0H42WOF7Hw5vtFGg2/TZa9H/UAnA9Iz9g7LxfuiUI9hsacwVb
y/aTk1C8WUMFZX+c1Hjz57+xpvyuvFe5iSVicy90+gfU4ADTKe/j6ZsHpV2+
eXWFlROYfMsjeaGoWYWrzBP6qTvlvKu4kvzjnvBGncgPXX8Zwo6no+TsiG4m
11ByW3RcYp2XyMBr+dFF1Y5F4HbK7gb63O0R2XaZUpt2+NqRWlBXIumlrviN
sJBQXCxQjh4xGQtg1bi68oyqqZK5OKdfE/2ybn2lvlBPCNoStjXP/KQQ345d
zcZVg0yMWTJUvUkfobl3sPltkx68QMFWFN9OiKYGtmQOhi/rYJudfObPaeLr
X6l+NSrmDZMlYvUHr+/FIMAhbb3dulrpbGI80/S39kZc9k9ntaAjqmrmGx7J
Hho6CPfGllE9HgoYTbHrCmMEsN0RqiTBrIQtN3FZ/0CbXZmYkcEA9sFCZbPO
QZEoF7KIsRQK9vxFxfc6NywToSN2ZkksxXNb/1+oTtxbSkhKeCDU1uHeyAYz
BlBNCzu+Ocg3q/bsQUAhArODmJ1D11mXyeEvWr7oquiOawJupEVhO9y6Kamz
7ou779huEo91P0NhGCoPYrS3HKK3Rkij5ddERKiHd9qskpQqiVxxzMLWdJX2
xx76LzOLtJG3n/PJOJNvmnxQo51xgKbi8VDZNsoWUNX8Eow7YN7JAHauhl3A
xv/nmh+v5G+iepKS6x3hHitvjfQu326mk4XOizYv6So+ciUKuKfHdqYAMjxE
731CR0Voj1Km8TGh8KtKc4qN7Venw4Csm9SSj0yqaxe4+VGP6M48Z9QV0vrq
shQLftCW9ett6t3miS/TGsrioyPTqZHvFzGR4Haa5T9XNpyS2Ua5Ed28SK16
QJKjNVSgpqDdGig2Dlw26vBAZkDwuw0bGAWMsAklEQcINZ/gdQ8qR+36qHSO
ZczRZEd89Xu+9o3nBGk5FyCn9m8sB4/C4DAI84zkVcd2p8HQi4F41242ZobJ
GPZy0r/WaKwb1e1NIFX7clgaBFuCfUe03DrgXBUJIGXoas1dr5M1SWOtgMCr
x6uLoFsPa42sMZGSJam0k4LVsy9YB79T9HZkZFzD1YEj1N/cT7Qp/Jn6AE5w
fELNjQquRbEZSQKC8aBbEWZSjPHSap5HLJSrYctbIWtXGBpWe5Nb8vY9RTez
uU7xiio4QxdOolStsJ2rBaS7yzlZC612vyIrzc950vKjB6A9XLS/djbVOo1j
0KDksJbvh/oKbyLV1mEiDgv9qehKWSEC7NrC6q8i3zzsn/VB15F56r4HJ3D4
J4AQJaZfR0GJGkapW5Amhb8CAE+2hTTt0WPRcDcGmX79z7awBxcT6KIGhSbA
m7otLKDXYsL/Z7btLRCjv/bo2kzVY5u1B8+U59LIS+mZ7ot9lZ8Qg6oFNIls
ISx8sNuAJCdj4ecWfF+eLqR1Fb2clDGskljzj6cWl5wXeCZzS2XgFL1YDRjg
1tdWVCtMgttBG363kUUviede+t3hzKCg/qBfFRFW9Pp6ZLp1JMZiIK11v3lQ
HZTDA/4kCERr0MogRgBV+g02wG3RvWZW9wmSrVdJ2HSzFqoJdKpD0tZwQc1I
ZU3IR/wJZFNLvEo8zdphe/AjPMB5GScvP5SJN4rcsyQ5OlSTFjDQX6CWhjyJ
qWIPL5femv/i+DD5g2zVTDbF3B3H8y+YtujPNM847D5Ku22bbTT779os9g5D
bDcYXTpTP7Af1MC9MIfZMypiRra00F0++cr1pIy6SBiwQQgGO+/JbZhiAnqi
9wXBRYRM2Z1jvTv6ReDTrdcv715ujnoZksKG2AX61EgtFkiGciCOGltzHrqw
46hEB9dFVqz+F0JvE1j6WOslJtjkdjtD24sHYyA1vaP7BBoevLqhf8usArcu
q9Ff92zpryJSmERiRMXVgMpuwLIXNqRUO5mNYb+MIPFJVZPtHmYSGuJn0MCH
/pSr83I4LoKJR6uFz9raXT6MNsnwAwA+HleKE+B/xz2o+jKm4ryVlgxivF7R
Wx7pZkwTNc4anhA7YZGxyyqj1ZskK+GRcayei+SfHZPXOroTzyZp5f5vVZHy
vtzUGGtugdVUCcwhO87/YTm9xq/pfmucmazmGx7dncQsGD+C3OO7M2fqL3rk
w4xtcc9eMLb0AEgt5Ijn3aOfGIjX1HnUXP3v3tWLkVn8gnwCoL5iM2FjjCIX
CgdXa/JnttFCcs7btMWyXXzESY3ooS5BxIN4Dy8ybom9eQ9HNTaxCvuJUzIq
5SLaxgPvCHBVkfY4nx9fURH8D33FjNh+hDiY5leFJTbLNGLBpTtehD59qHk7
xfkXnS+99sUz44AblYWqJQdLs1xCgv3BbhC+i5oYXhtubDd0gwxr55i+huF6
JW40f0EwCpSsP9uUXdxF+5PyaL3mnA2woTydiRkyAxxufvqIEJeb8u1j7m2T
ltOKpiwmtbp8ThNqACXJzdyZBJUFuJXwJ76pj8TVDKn0hhjYymWs0KtoeC84
X23/bOmH3qH0dgFC0fXvvLY7BLuIHVwbVzZ/vZTq3HWKM49R84xejOjwVcsN
FetCro0ZSyM0X9phmT46UlTtyArSPXZAhiSkigIVQHAzuULb1RnVOtM3J6ov
t96RQwvyqbqUdP9WSH65l3r7TPZJNE/S0QQ60bZUneKJWzG0AfFXiDzjmMlQ
zdBinhkHQdeJpq2Tf49g5ytyxYgjsIBbPzThbQ29deqEtviwRJlJhCZA2Iwv
FeIy6VddpNyAE9FvaHQuBW92dEHZSTuAe7q0BOrVCVKfQ8lrp/uSg5wyRIYI
01ZPBSdr4OJpTUElQ1bqHxB9lU9BBGybabwgRJCL48qtsl3crW+5ubo09mB0
dd3KsWrz/JlbTatjxkDGXTn5ECkP0QYUDuIo7n3UOUD7enf+LgcDpGsE4T67
V+U37PBlR2p/wqLgkmWZTBq5uivqmlupWt6emFggrRKivKWPmvhXPZY4WYcl
70Wnpt0sNDLJ5o6Os+Kvuy5l6jJ3hV3zSOnbPwuUx8XaLIUtQGfuG2lliNaZ
6nGSP8nakvzIG4oCA6eJJHFAkVl51cxfizC6bJLeETlZQCfnX8aOTrN8ip/C
bhNW8SjyF9PbWCL+YmUVPeqSWH5ZGvar9DeHLWpSVmKX7vDFBi3zhTkKpbNn
+cKt09HheOgTm647GnvdjeRrcl6+rvR8mpgW6mydohnbY8pg15yl/Pvp1QLY
8j+8KPK9voIoNHtKt5kRRqOnHjAwNdYVE9aDiC2Xf891uxPe5lbCftUKBIgc
CAkkGxCEAbr6geBJfC4884eg5vZRl0Qgnq8btkTcpCZ0eS+8nR/C8ug7NrXT
2yCIr50HPrrk6TSeE6kWndDKe+d6xBZJaQUE7ozkc5p3SZz/fHv4ETfo+M/d
zpN20qYFYuFxjrpO4R/soLXyDYDVvSKkh28bJuoUu+x3AMfJUHgeAlOA8VvC
plPXRrzHkDJTshsEjcx2GKNXgcKR3HFdd3U0lLgKp/ht/MFu2oeVVDOh1+HL
uFR9du7qhBdb4ZLsENBBE9gwGIFc9rHQP3/QzOGMzTFnEI8adQqkim7R61s/
sgZ3sMIEEfLi+UFjCtq9/2w81LrNaa2nuUL8eDskZ2grmKJ2P2eKnN1wuh/y
bvBEpPoLyTowlO9GfvBTNuUWCnTpmMzSyKIf95O8Iu3FtJCm1oEzlBcWInP2
9GXdQIANGMc21N5S6btxN4w9uLlfsekyusI/WOR/anJqYh6lEjVEz8cJx1ar
CGcmsYgCxOuP8f49vFRXBApdUO0Fu234XYETwJGdylVVC+TaUhGo1XMZVJOu
Cm0rK0JzVkKJXB+O0uiloz1TpzBgcUs8F9cfAU31mJ+aSB89tArJ9oOtdorn
l0DieCIOXX16vponM4YIUzXGz6H5+eluLnZfwSIsao1PDgonCexgBcWX9Zg9
rGA3SoBn9VwoxQP3TcqxTkdAfMEMqZXwG8ZMXmPgxsRha7wbgeHB7BibsW7p
6z9gN2PjRh2POgPUhDmjhsgFrQxFerIT4uU4e1nudg808lypuTrUwMvj/mDE
jHcFPRaoLDGCvqkfBi7s90pQ+tS2pBkmNq8PrsXsx7rhlIhzKebzfjrMj3SO
H9l4RN/MMX0a1OU3X5r1VGeflj9lBKAQ5WLyYiRfcHAHXITw12eEY3COdLOd
SSIGYiuU6CT20j/BkYVdluOL8dydBqKaQo2epTZvD9t+IMF7Sch4+0YDuvc/
k/Ad+IQ4N9kJYDWBMkXOpnOE4XostDaGssjKr1d0sdcL7zLavy0sgFVKUTDx
2cqyI45C4CrSHKT8SBALQqKfhxtUVqR5hInL8xzAks5BY3UULdnmfiNy9QMH
M81EoKT0YO6UkLBC2F+hg2WsuYYAO01lxzbCECJsmCO2Wur5zd1lIblHmBbZ
4cBPGnt3qTKg7XKwJAokNdFzY9uO6mREq3cFRQF+TRK3F7kBPyo+9KFJrGy1
kIjPSt4X004Q5tFzkpmokVBsruV4hDQ0XHKtyPSYBUBfZr0UxE7A66kQFkJF
WO5rRbQzVRg8nD2071cQZeKj8F/8dkxjNnlOMAd5ZfCNUaSbNDC9HZvdaGu0
/6z5NNzDhfUmUDNl5gMGeM8TdsLejjLtDdDVodGkJ40jYB9+BO3JA3iHHKeI
ndxIsgV9LGcWBGithtos/IfxGMpDkUpXOJTQiUThx3sl5mLW4H2lcOjvDXhl
hst6wf89CfJ+i51ASqRHKbc/UiFTb8eLr5NpDI+1+cWQEXQJDwaIAMwF3AY3
aRvGhOVYAJOQ0ZDQKixK8wlcJm3FNxhMsvm8bZWL2hnOJXz4Rwrj8IvrNUyj
1eJCvLn3+f9KJzmv2ey92oS0NOK1Iq+W6MIw9w/gGFWrk0pb/7Z48UPqcoqj
uANPSMvJcjIRJfuii9CyXeAtqMw1prR2zx/TmHgS6t4gcDvqYPuskVdpXjtV
yY09XvpQ6oFu0lTpU1pqf2Yv8LyCSmwxiWRmSqO0lA64TbvJinrLi1TsnfAy
Mne2XwDvmAdYW0BMY01Ym/lY8JCCI3uOW2yZ3bJH45jtrtFDd63jpQRhrJOL
6uOK/Aia0BzJYd2sUHwFLg8QPUMNlxZDWvaMs1AHXvV376F6AhVqwZjro56E
6uotmsStWttOPXnhRFdl0PkOrOMFTB/xIXKA1x2AmvLQ4kqpCQaymwN7Zp8q
hK9B9WTjnNXPKvPGZlnGouwo5yzES5qFBDoduKkDIDbv/pqgC6jGtTcShyfq
RA3bmgY5pRkDVgXOPll23OCgQU7AigFDZnVs3SDxjcUGKMStaykRpowmFWSP
JRSh88CYhLFWZib+QZ39I/bWE5b+jfyQcErSj5qKr9CzIDu0J2IuuZaQFhTR
qMhq3FnDYc14k2XZdQwN7osIxdkAtGcidByXfKRcd4zNXRensHx+b25r8Rtk
cEqorVqL3j09HH/FFW2aDeTja4tC9XjHP9uH9osMBayF+vo08GC1mplRvqvW
otSp2tJYMbdISKA5aFuFepjrMCFheuTA6tcsod+6tzurBI57U4ia7A1itCg8
mAZ523/kB9PbZWqVlsp7+y2MKxK5yY3y7K/4RuGxr4hDWqoMsB0GZeR7kRm5
hQuzKm7BSHpPXICX8ffZKSQTgYKCruKzhMKvXDwBnsBdkVEFsozyyZYFxqMi
j9jF6MO4f/3Lle/bzx2BUvTd/pq5fIp7GoDmEzzXvZORS8hZq7HVc6mg6MT3
OZttrBDpebtYEJwY+C8z4va+007niK5u668ZnHuMeZGlxQF7YKS1VkCo5iB+
NaqAhnT7g/9tN0F7wmsGZYpJkswkSanYtyua3wLPYAVhC2PfLF7MMtuuRpn7
oFIpEvr2IeJvHqxHB5BJkjVzyra6Ctza1xjva3xU1ievSJ8dK/jxMCSdK3gM
+79ZKF9RaNHJJ63ZVno831CQwirn5XFgKBgk0g8NNb+xSx34HPzLD1/ykHwu
ABirPWBRRQZHXVAG7x9hdxVm4kJq0c1IGExOQbhtNNFLXDmhM7d0VmgSumzO
n0k5X2a9sTUzXW7bc4Hr/XVgHHEfU43Nb4BOqMgm+BMfQP3Wz5J+g+RQ8jbv
qVNol4dad2igb3j9+1TUpa+DxD8msvqdX8FYQd5XFwehMOGXyyF6kJOCFG1G
HH7G4no6r02iUgrz8fk6MrJBhK2BLyNidOfymZ3kyt+JJvqlhI3i0etuRSfe
qYgpkRRTCLIQGWV5bY+Np4/tjN8fmTA752AN96bZXTx8l9HYc21ChEMYG4Fj
K+oeRcijM59df1XwD95mVXGTl6Amj36au9ARqJnxVTz1GeSHtbzbRDoYwOfw
T6Dz1NxCSxj3GsY1tPjTXzV7s5qTCY6DfXnLLaOb4UqYZ1o/3oFAbjrwb2Zn
NaR+ct33B6+pg0ys+h2YdvW8JXNmEGSp7X7pLMUL6ilYdMgoaOz838P8zu5j
/juC82c2dnQbb9kGq/D3o3nsTY0gaSLapQAUPQ6MLZ1gGkFRAKqtH5VBIXc0
u9y0TdpFBg3BI9b93KQGXjavgqxyDL0ovejiGSClCzeOIQqOVp+GVJNi2seI
RRLqIhJcf8g4U3BdlziCcphHVmttz6pMpmio5W0jRbWbWCKF24d+fPj/qtaZ
XxYw0uE27vGv3o4qMI7CRUJcdNrDx/+axv4VQSD7lpp+MZg0LLLdULA7iIoi
4bUAeAFTzi711vjxy7vaQVhHBYvw8W8B1AT6r30Vo5UWIZVj6v+HzVkYvgKr
/8z3/fROpaAyZ146uf7gCBgQk/DoL8lY3ffP0llAzm8Ru0mdfcQu6BtRKTaz
keN+NqHpOIaoa+w5AtiBSJilGE58q0aDdfh7SYTHJrwD+Eqrq2ALvvd2eMkI
mDtPh2G7SUfAdpRO11MY+PntLWC2Kxp4zzE4G3cdbzwH0E9x7gKSaVrhPSY7
sMbPO5nl87TVYZyo59wxuHSS5DL0lxhO0xbXH/KXYDT1kFVh+v0GGDtNSAyE
/NoIYQJY8Xg8lneuXVhzu9NFIuKi9nXQmPovqaCh2u9aGqgJZ68zAsC/MVMZ
GBo9pE5P55GywSUN8QD+y7BImD1dbkLQPNghyruCMsRVJ4Bd3eEmbTwB2Vpf
5A9njq5kTLs/8wgEljByK/GvOJH4AYCzGhpyqEUWhkTVFN/WJ2GrrzkZzUxh
6qbf3bA6SVvYksLhfk+CP3IG5iv7Fta5v5n/VincbiCrsqJY8DF8eAgxqLNp
ggI/mUBJIAfffKkkxpJ3ZRN3vtW+kH4QweYLPyVskimW+feNfP6Bo2DznSlT
IuG9+VGLt0aLC6SsWbLzNQ1bQBf3Bwq12E161NF5GrQ6n+aw5OaeWt9NK4g+
cT9DO3M6ooSaEiBXRisc26mPG1t5TnN8lbifqDwHbn65qxv4pSwsgw67xsA2
cAR+vfjhv0F0P30FovuA23Gi8LV9lI4l0SgMdOs9m8B+KD9N2Ki9i0agi3I9
FXumSgMfX4pO6Si0cakFHIoChAPbFEkBJuiCs8twFxCB9e22FxvRHYAhC4Um
fQ8TCl59mQ46YHfrFUZ90Uou9ReVkFgCUM6FZcJVh22Ak5qlwcTS2+94i673
xGeHDy2Kvyas2a6nxX049ReZs9Pjy1HOqYZtH4j3rj8QebG9Tc3z40++nBtU
TZOxnZsCBxcuh5SBVNmEslKqxRNLvdQdgcwWE3xwmtROBAwnfd3sM+RcDza+
kaPtFISYC+CYVJw1Ix2Hr7h0G5uFrY0fsixnKNjGvOZN6rZwzyRV7XcJnu5M
qfqwYXv96SA2NzGLF1qHqZPk268e8IQRX4i9HHz/DEr7FzI1AyywzIXWRynO
cg7D3JZS1k1kh9KD2NnJfP6+cFHWUsyEULydXikV+qNHZHc4JGBVoQE+OUpO
rf4UMLWxpmDyioHCWUkd3yTYXH5vT9uiihWmaCDpBOlDbG9FXQt0a7Z+UvTj
kNbauMJcIw1qGY7qmh9fC4Tvm5lyZGxE37u1+k30V5MZGwF6Z9apy/q+Cobz
wLgTsZj0ggD0Mqt2Q1uMfSkqjVQcl8EOF13Z2U666nRP8kQt9B8Gy+27n18W
P3G99jpvTZBYd8YzDh9pb1WEsTDOkeovTlLCib8X6Lx87e/hf/+PvEUJn8YW
mmnwBmOhlu/jePohvt7ZpD+z8pp+K264iP0DQAook5Jnu3FtUIaQsMFdLuHk
yBbpaNVhln0i99Q0+JZI76tRQTZZREtmlUAjaIwidWNMk+jZdKg4XmLBwEDO
yvCdW8S4ucxQxua/YE0mGv4zcqvuLvJ7PvyJmwyKrlYy80nJbcEz5sHDQoaV
gYf5pTV49L1Akm4YpD/kOCn/6wxacdAdopdBM+T2VD1tmJqVG4+0YWT5/Cpp
geJw+rd1ADL6gs3rjn/HqOnqLtnym1kLXUhAneoDTR8mzuIo/LLN/pgYinMh
r0uZss+ImLlX9dPNXbpNsSixgaHpSaQr1pkZl44VzkOe2Q247sqOyG6lf/xk
kT9tVrhdZr7XpwKLOuyKKZTywf8Yj0kg4+A8L+6+GrJx314RRwtlyQkbLbyC
XYcd/d9WQZCw+NFIQAmgxdTtY7vyYTHlUu9VQwh0ZkSO92F46vwV5Y71N99R
S58DnIfea3PqkKkiWqFdZmrvNrHwjJT8648SrOUgM8jlFyg+rldFoLGB//mo
xiBvufvuKjkqGVNb1o3CaDkry3qDTgHE4S4I4f8qdVHwKwk0ZRL+GJPutyAs
LDJRUzQvRSBb5a8Ds49v5XfYqz6QekrCnyyZXjwJNME3HBUHGwbSBduc2ilh
KKPuh8PEKjgtUqOQxzY6Uwvc7rMyinYrOd/tJuWypSHQrsHfD8Vybb9Ae/vv
zN17dlya9hTh3guaGfK1Wto7nGcyzd8jc5ZGdubbJmIdyFbSP9QM5tbL9tt8
4dzxbQJMCRpnE0TTbqBOo9z1m8WzAWIT0uVSREpkgC9MOckZb5Ps27OGDLPL
dwtaEMc/ELdvI/svQozqyj2M7SlvrM83nwFPsQVHyi0CXG2wj55bkIS2ZjMB
LBCUumGKphe79dQDhGKJXUFauHezt335RvkW5Kw/WC3KuUNa0odtVvsGjj7b
fDSHcBVr1iOViwv+I7lIDUgpwxMUci7m1n4csEWFz1SPUEeL6cT1lWMem3DL
v3idS/q0oMXsjPlbTa9rEIt2xypCpoi9fK46jtH1aKr3r9mFfu1oSXyJro2s
0Gk79L8hJ9ztWRtGnR5dY5Fl1ggrI5vhtgMHt0M1p7TMzNfSORhSBlRvn5+c
sSs7TTULCJyRFE6p+tAkHvMZf5CRnBAwxWPJk3fSgmAp4zy0iPD/3dg7qj1A
jl4z+hFryVplZ9OIs2eEWPaRppPGTZEBcHa0hXqWaPDOVOiVeb3a1Dha9A7h
1UKWtx1wlIj0zl2CbXpOLdtin5nkbRbPMoxPR/IqQLT8JmYNojGORoI1fno/
78SwKaQwA5mN4RvwDuXg4QcXUjc3NRUhEDSS1vESfCWip5VfGZl4E4VQIWgF
MIuFU7/l6IqsFOU1NKTzBhGtFQJNyfxyF/WOEj46NR5xyrSzpLVcwkXYCbGZ
9ljL3OTkOFyQREzb97DEbYPccUSRRK9J1v2Vj4ibmPoLEajxonqvXSEZttWc
P1SBeD4yRbMN0DiNDuvzljhktaSu+NU70Q2bkKLtJL2MR6sP3eumgCc6wovC
GxDsVKrY5a5zRhq8mR4f/Gxw+OBIukVUSLm+5Sh6JFqhkZM/CILT8tkcsyVx
jtzBVRrzSGNTXBLZcYFzNNXr4Vqh7M1fL81Dpk/Ig8UsRU4UlG72ETkpGeFh
7caQmRIWMaLdd7xr87KyRhMn82WVSgKrBDhz4HEoINzgy++QuIC9rFUxKnaN
TIUSTAHTDS818vbA311tRkzU6Y02HsBnKxEl+ax7nLodfDA2nNa0y/qCpi7O
rqycxc5Pj/6mxnJrHvOEjdG5SPUCfzhlPJnZNdx1NcQBrq3bhdUUDCkNwKfg
zcV1YMb0m5OO0tKH3vCSHDxZwFMM0PfBRoMAoiy4nTVQ9nQ7AG9mGzeCbB/l
24j5xp8ww35jWwuUGTxvJDxjDV0JETEJCBeDhnKQCHqF8UpdPkfjRnOryTat
l99Mou9p17NsrTMqgtsprazY9dXVXlr0g/EEyHZSQckx3MmJwuXXcmhLCN+O
2Hbq7yUZVjZZbrdAqGeSLf+nJhjFI+SO9yOok+GyQAMUNhdevhizyKNn839Z
tApYvblwQDuG9AtuzB4SK7mS2bDRe02iuAU+KVYPyWxdi3cL3zjGXQ4Bc90K
u0T5qE/YdfrBUy8rOT2aU9dh6GUXGRY2hoyvELCqdp1h75tUEll7JWWIaYLq
JjbNfabId4icL3ElviqquhonANRVDZ7X2dN0REh2mAAty6exTje4Cmz1TCMM
AESXv8ZGEi/9l5XYNRKx7r7DSbqP2mr1w81iozmsvZUJjBcNPbEkj7TnSEM0
/TaDRNA/D+6JAVKJQ2RdDP/BTjaKZUEfQr4gkhsM3XwC0oQ2Zqwi5teLlEII
BgACxfBuFkwE3Aht7ynyz309RNWrXXi46AMsOLwC1LV1H3xehWN4exC2GuqZ
z1pY15L9Gw+KWBvNFcmDK/SaINCIuCjHct898IQjUceL6s3QnNKRF0S82aHs
lUjfoauHVmIeZXJPwhgJVkWIN+GHuNlU+GRjlcAbMSdSGMt8670O3lrhcFT9
ByHvBi6gmpiT4ltjzrlYIB/x6yYxCcu8JDVRz7WbKVMN/pDQ6cWIVQMOqk/3
4AuaD+cqovk4Be4xPKtC2rSD76Zwv/anWCCPzEZEFuw0J4RGOiWzpaxmP1TK
HvP+f2hkIg1s3xnNe3cMQAuDmOk5CsB6O75mMJX/NmFFw7T61ruh3hfIDzwC
5gxSAIgthcZFxp6OVrembNWvOv+OtQuTtDCn00IJX3rEeM8fDS9McJKp2f37
RWM1JqZxCcFyObOrN/mWn/SprMhJJqwuRlLljI3OswZYmB71Bfj3vDBCuGP5
7rwdlI8rAVQfsBH4QbUY5/V00lMdrNjwIyaKmTKUm+smh9QO3hkHv8rHPk8o
+4YZBO2kHUBKBtmZijf4iW08nbbNdonckOcu9m+WQYUXN456aF7DwmE3nJUm
oZNdSNzRlYHlN/Fbv8IOdBeXLeymW64BYngKGIjVlW4IkP2w9z1qMmmGUydx
XMyu5rDbTQ3OwfNI0W3PRRBIuRLxaoRMAeP3odHWDic27HcGGBWvVq1jXHXr
dVsoUAco/aJiOQj9ATXjHqp+5hRrqkE8Tcaixe2DolHPvXb3T/RExf0O5tRZ
22fSYRdtnuPWT9PcgXRRqLBX7ZTcvv8sYuJ4WX3q91+OazqH/y4wTdsD5knz
Y6YrAe8tQYxSG30Rav6w29Dgs57yL682EzUBLlcgdC+IWUo76Ceny9ZkpYjg
sXtHeGiTq5pSklo3/xkRvvLF+xtQBKERnrlm4/VFHy+BZPIlmnJa49lAqA/I
fNq4UEiG7W3MqNqE3DdJvchIwf2zfu4HrY2ulEvBlKo2aCDJDVeCyh58i2O+
wENsjGOlNfb7G8ypU5fOWQfn/PsFvpNyrltvBP/ouWZDsf/hVD8+IpCK08mm
Mob3bf32CyuZEpfdXwbHkxJ93J2YT8yCHoRD+LpN06chMvY+EGuhXZ1sUjcA
uLEcyPbgjwmwf/RE7Mg3TZowyosf2IuyRdk71ClDl+UXuemKoG15Xt8ctxXs
2ib8/JSweuaaat21MU4SdhK7aR55hWwRcXq0IJd05qESepkX/TNolTYVX3KB
WnFYeEd7pJmMAPpuXZHdv+39fv7H+GqowYKFVdhgYxp7EnvY8hcJi8cWqb9k
VLlEIWOEo1C5Iah5XRw502gLwigc8nUcN5vY84cgBUUUlrjh+XeyQU6Yez1M
axP09ZUjEEekBdA+yX29o6pn6oGNyX9D/nzzz7l/c2CbAaRnM6mNM5Vyc0Zc
exZs/POHN1iJsEAofh1+vmC4+AHwmX5cpl9tGNCvjO5ls/8Rc6kmSj6UXI9X
qk/oS8oERxvnFOVO/skq6Yx1Ueh/yV8Yhr/f5Ecm504rjNNlcuEKwxitDazc
uqHBadCxBkQejafKZae41ctxMzIVfHkxarxiJNFoCNHgjcbvOYN4LQxTFIoN
KKPgUBwBTJnwClV0rwEXQq6s02LlZzoX6GGGmHOUmn8J1GH9ft3HKjOHoHEY
pBAv1WPGAbZDqcv/xFvAa4yUVh/4OKJTqR6AI0Bda78bxWEE1AZ5MplJTleu
Ee5NYAZTZSaMe9EHshKVf2C22e2W3xMJ5gcjyfRmebu6HU9jiTg53Joa+VIK
/vBSTjboDgnE6httNXlfDpUZeCtpjbEG+TbMOdt6x2Ti+5205tjPz1by8wXt
ZNSNOsWh8KDyBE8Jr1l2s/CI9r4X+3aLYGwmFTNR4B3HbkDX9yyEtZoywBnx
5L+A0SliIb/u7kR26CBOqcb5zUXopc2CIbXnTWjZeGhsftdDMTXudSDd7qHJ
hueKcvHUkWpqbly6w9c32/AQVTe9y6je+Cg21pbfF5Sub8Ej0q99xFegbyAX
EOHTgq6pRNjEKAZqmZvStvEYqU829lQzGMbg83JrX5Zp61R0PImapNyfbPkv
YYqu/+hTzORkDQnDLyiDXGfOfsHlOxrYuWGjbEsM/6Rdf2aVf0Cjv/y3D297
cO3F3pK2Sdcl7k+x2aFizz1HDGbfRWUa74x74o1IUjJn9lHKwls6YpD3733X
DFW5MGBziuO08QwF9wjRZ4dhUx8zpQEImkM+91mE1KFPL/8/W5+nskw6rEs7
b6RZVUKMxfbplDhVuqZgUhDnM7nRAEXRW3JQukNP5xSzZKj/mFbyWOMTJ5aL
0QDBF1w90X88X54/EUww8Dk62wbERdil+8qZ69VZ+u+jvI2t1IBKfC0Sl1TD
OTyF/MM+8SCp2FWs0WF0cCNdMFK4qufRhmDR3Y/C+0VMjAq0nA7T/I7VYEcw
KoMuukQ5MvAgrEnmkEIU2q2WVlGe2+J4mpmPHqChReza2yI5Pzl94cdu+Stn
Z569i6N46csXgPD4BymI7kh4whPfPqivWwzw3Cu1mxthnscejUyvp4udxh+H
dhqwh4sZxERGkrME0RovHUJa84p4hAmUBwy+n8w7r5BKLeS5h1VwiWsBIRI1
mBo6eLbOIqErKAfwK9/pG4nwPSIZuGmi/Hc4I62/+DTPRJreVGEdxifMsgSg
w/Buq3BRByZVdKi6Iadbx8//v0oJZnZHWPKQfXNB4BooVYlZLdx3zPxDbZgG
mc3H3XGiUfWPpneY6odp+wWt38nwnZgjF5P62FZ2SjpegdFTSBljyea8xfIx
reWN9bin8CLPwVOcAFt+aUBPHKg1+pYbJ18VOfeCGiBBddyWEvo4qs29Ckm7
e+x3GUg6gr4Sa/AiydZ1N38gE7Eqb7O27461JzkxiJ/rpZhE8dkg9xPTPv4B
p9qvLmLonzidEhXyDRVHmPmFlt0EOLWphtIuweiRsanb6cllzWHwG4Z1uI85
TZjHGCfOATv55UXQ64e0TGvgwKKvs2VvevivnokAsQNCf0fZTPRJ9tdJ0mHf
64APnd1cviIQhcVFdiPrP1PpGL8h4h8VlDoc6/Zei8g26V15ArJjJbJwUwGD
QHnFDNv5XFQhqoIZ+v2zde2BNcxgmOHGBc5NSpWq2OZOLOdlRImhijK+ae3q
+qc+tZ+QMHpuMY4uavb81rrwSrWK5n27p2vtQkERlwxmRwD+fMCtnqejzClH
bEldsjFK5ljbt6AiCtUesW1/8pPZcsG7t04lhkCqme0gPzT6eqjJDAIdmdAw
28pGpKEBk1B/2NfzVH/nC+jZ0V9nKArIdf3ItGRgAFAshKQvr7cdd5dIYpNK
L0J1v54TSGNbfc33cOnTiiwzc2ExABZLSU1/w0Z/ws9OROC8+dsY1atO6n17
7zol/UOw6u16ozQ2ESSHzuZiBgB1oXPuyaOdOf73LayaAgUHhx79yYSgxdcj
CK5V/x+IHJLTUc7JhEzqmAC5gPVzKx0OMBkfG+r4LEg5tOtz4fHTolmExWO3
C4JeBvxZe0wqzsXtbrkKjtwZCiqXTNyh7VwNmHDrG6YnRlVol1R07FbWmMeG
uKVbMkIbSuQLPIQm2cHr89OHazs10l+BeHjWJixjetOtoNP4g4U6cZEs98LR
G4Zg71fBaNmZQ+ydcVGD3Oi3M//Yr4X0TMbDBOTaaMP27lj+M8t53ZjQSg9P
WMs8kz6QgMMZTTMnpbMfeDZToiGZe89/e4FQok88PPJ1aqkyhgoGp6dfe8J7
PjiuLfTz3f1eNJgoNYbdg1qWm79BBYn0UHEWvo5zi3vp0fk7801Mz3jReina
d4kvh2XQAz6B2gI3VU0biMoxbedRoqwApdKQecGgWH1q14xE40YtAyLKL7lk
5w5zFpkDYTwKploZc9R/iT/gBnJH8xoaWiEsOJIi50bCEztxelC/QRy9aVXm
VT6EceOQn79NHUBxv59mAb9BksSrtTmjQpX8hdKgcDoF15DOXrgsIaNsx7J+
2ojvfE5nXXrkrGbUBFv9z60QP6m0CA5O99PGn2+ISwKRZEQ9apAHdbpitVXL
i3G+T/3mXQSGQv1pCoxdzjzmia9Pnf/7BEw786Fwf1nxmBSNOUh0BoVrScrX
mBFI+YxSTnWbdhcPYeoQbDsDOTkC6O0xdEfCP6o8NWY8gq06VWwUNH71hrBP
ZInMnX6oRtVVXkA1x3qd8QH0/q6ngEXN9If1X0Dk02tvJn3UJQ7b2gqnxtOP
0ZdvrewI7PhYcpj8IdPMr5eYttMsmsJX9t+HohWc7inStb6uQI4Tu7wn2nCR
BjVSM9IVRvpIhKTdsyh+MdoklzyGR4YLafogXdNXnTJUR4vMBhSS1IHsCE32
vNL9QwzI7aS34tB0WambpsmSpGRaZdvM/QS0N1s/m/GYwBLoFb+6DsILoYAJ
yDgMCOamyvvg162cfEwvjM7WO2LW/3Uj9rWe8+r6kh7bbVVtgp5udhsY4nfL
PYooU00ipfoFO25UM0ln69RGuGUxxJH7+GxPtPrARV7iNMvbGGYy8Ab5fX2S
XvkYUNz0sicsO6NrAG5PMeOCaKWr0FzzffTlGK/NZrI5JA/I3aMjod5ZWX6n
3Qtsecosd11y4WxywaHjv6SB9GVJW5MMs45qwagPVFj2BSnmYtOwIlmtCMiJ
DrjN9z7gpvLn7RrxOLUe5YYUeuihwNZyjRzy/Ahw7a1/y7BjdSCh5ut2Oegu
3j8T/KncXo3tbhD7Wa2h35n/EIkh3JsQmjxE7SYUSz9MNt1GXZR9HrP4Q3na
mGu0agPTvX6gS4ihAmbEKORRCRc8MRAHhUVfnvP9IKOeMV20J+S/ZPdZ1xle
95NeWhtKPEYGU2gFV/YGcLrE6Jcae/dV2fcb47NmDwb4ZZaRtc1vQW913nXf
zk+J7cetpZCJE/+V7JWV00iLA5nZyOuGjsQkmtA+5pWhYdBJ94rudm+feVae
M4Y2L1Q7KCxxJGiVJ+GyWv+4XTFSu6UJcJvv8yf1c4cVG/Ij5gkuDnlOXqhH
TEPVkx16e/bRRAoCSlgaiB5mV8gtHgWbNB/iMFThnCdyyjPDynfMVSJkMjeo
+qkV5uUm+XGfg0OOXVZSlnUjEeClLSTceWqvAhCce+lyrwvHoubH6f4Q3m5v
S30YOuXfPs/Xrz0EwBdyHjPT4C4+8eMFEKKRRoMZsoNp+1fwhMlKld402tAF
WG60R/PyUWyLoKcR5LtaZ820lkQSzU10krNqQHSkDv97QSTgFI82MCadBbz3
ZCprHseFcNR8TbNj0lDw4tydfEqZYGn153Bqj8XxyCrOSKFOHRG32bfO3Lkz
iwXOnk9svlKvN6FqK+GYEeC1ACVrBOwacNdgb4U4YT2WUXb6EIRGloskw3Eg
sNdm/0m4nbw8x8As1gHykYV5KNoLTk7f0KrTyB3tejVax+MdQt42qt6OlSXy
yHhmo6ESU81J9MGNA+8ZAWqBrNWgY3MBLQjMpTBB655u9VuRMyYJPrI+6QNP
//AEDMXvQATza0d4ZChha8l3pspyOLlPSVwqnlpQXkywqMmUuNTvtOvkmjcd
tdsXhi6bWA+hFOZEn6FoAslU+AAlZ4wxD+zOQvdfppC6FzXOfNwZISL96WR/
8a4zw0PtjJGg8GFC1Hk4L3PeKuALUOsESmJhLqKYGjtdxA55e5uUTau3RLYY
pthnCZOJe+WjBUY1d8WdLEAjgX0FAKJaV524DCq3inGAULmsQcuBR5tjPNcC
y2dD/ybjb9tfXsO/TwdAf5Ei0wCTqusC9Xvfs+zWzHg45dNmM8t7ZDl0woKz
7dAS4kZx8THEm0H0idsd04AZTd2pqsxFiHQuo0LWLVXH/tXF1/DtO3mdpC0i
3sCwdXfFIhzUyJs02awTlN8nxWsUxho0oXRFIE6iuUOsJSHobEXlPYeeQReJ
aeemmuC3a9bJgRM24PJJidKD3KSg/hvgpEX3g4i2sQ6Eo6RQ97ICpbwGJTG/
1cZCAPp3iT94zTNFBznrkcP/knXtJL9CFanShcsPNoXbmQFbxJN/rg0RyIr7
cVa1QC/S3NSnGoZW/bBJAQzevOaF0XjpdAfhyxeyYZ1yrwwE562NEBMIjgQQ
CdvdbEL7RcMYq+WnfMNUa09D4cG85lAPjoEkSEbuVk+5k5KnYilLF1KXF/l/
Ytv8yAdawD8grPuHGqCaKg7kQh9PJlGOz4tRqp9zgvCherRVFhKan+rXVVPg
WmmRXRVXusOPSEacSRibtRiUpN0PjodB04HMteQMdsmprfg1I+ScMJsrNIyy
EXlfwSWmkBXt20v9+qGz+dekgRKWEH9AdUsrxNHinnaw3fNGSVEE3sz3UVWy
m/cabXNxqJB81uCvUGaZ3+UDteDH3B+aBRAl12yGrOSzRLmB5hiPu5EsR41M
7v4uSKNtcvu6Pf/sVt8rJlhF39OX+hyJa5ZYtXSf4zBn8AIAZVyTpJRYPF6j
pnAXAZAx5gvMR7v8BzDaduGPykQf1P+l4lrpWKZ6nA4u7A0PKT/TgX+xcZv2
9yXLEv26/N73eP94OlilpXGDk7ckJi/5qKGURT2cLeNSisaMuCtaussptRLo
r9/1eDXlzEwPkm9AAeMfKdGVhQ3geyT3wx8li0udcVogFCdPEsItzCoUgAQS
RdKyYd61NJxnwOpOSjHeMoHX5Qw9zlriazRVuW4nBFx8FF48Tw/07Mh/195g
tnraU6dDxt/Es7TAv3GD+I/bVHlqVnp6fOmsPAip+4q1RygVwg5oVOi6wrnC
9+ahF0wgdBe5IzRZ1IF8QNheWQb8RGZDg46LzkHTe0+9JTYWJh+8LFjUTYzO
pexYG2bVqrH7AaY6PCdg+j8gEhF2/alpDGOVxpNAZzh/yFK5Tlxx/wPV0yr3
0801yZytQmp0BYeh8WEdnq+ZkEwFZjlZLLCmQGge6cwEHRKFxgtChjaNENTJ
+ITU6hUdWXLTTafn1Fgjo3jaHDFCE1aCuF/1/gAMpxPpJwSHKoIoHXUwnUpb
QfRBrpA/fSKt17Ua3D14mxmwTsda1mB41oVHbdZHerVQKpfpvEmUeUkhNqRN
2P/RW5gtXTUB82k30ZXwxOu0BRdxR1GgfGJQChdPg7L2SNW33lAZt2tzMCrH
azRe0T86OwyvKXGmWEWSTs2vklEEcucKKYefRkM8xtrhPDs8OYQ+AYfBb+5u
5qB24g5r9+i0pp4IPOz5Sed4WuwRaTNZ3h6sUcTeSX2fDIEawIOqRh9NMPCB
9jhtg4WDgxjHsxjKRbwlV9diKSE9BZBBOZKf8cDEmoZg0JibYyul/IscrL3i
vLsLQbY2GfsocJuB+9QevSe1j1I9CYkKmIv8Nb58wE9L4DiJpvpq40X5rYDt
JayRjwf5kRrSp6KrMgf9i+8vwW4uzO3Cd0s/fxLw5MymcjsJXcfvZ5fiam3D
XZA24EeWq/zqCzOnGXIRjT0LFjybdC3n2KWYVij8mIwEfg+g9QGkWd1Bicbg
NIaXpKMGC6s7snBe+H1Yut1RQD2DlmWbGys1EwxB/XsRyL0Gif7vHmg7uHLL
MPpDjYA+Ni9vjykrOK1R9Unq3tJuDVrj2bHeM2ZL/e9XBsl+EFeCQbXV0yNf
axfF3PPOWQSzXF+A+lv1TMz3TNAKm/aJNUu5LFQo6OaVWPgKkCk/ZMsTnUJ8
eWzMkVfoAwImYt0h3z+vId1PHIREtc60VN7+OOTwBmwY3bfoBZJNt9CoAFCu
+nbDZCEyxbF35GhdbuJDfvyFTKSyJO6VdgdwlztkTZsufRytFWbhUYXpfc0E
N1Vox6u5sn016CK8FTtT4amkx2OHcnRSPZ12V8pkAxCFu0SBKBpZaINwLk21
gMxLBWmFacYewQB628VaznoI1d6Jycg9GLVaUxuKDYHlyeLPUDLKOc3KWxIW
h2DfhnRapvlnPgSdypdml2o551c1BN1CGveK835sLCnDmRPahUs5UjUOsJmg
ldQoPy4WWlXhHzPgvjDKPPJaQsnXKBTQXF452TBLUS5AdGtWZvbGomzW2gci
9dgHZKpMcvJSO2Tkye0FXUb9JqeIlqMqotGeN/H9KZNKUOndBwWt4m2Yjdif
ZDwJ4wTRR+XGQQXmp2JDMKptcFU4KtsgOVlaLQDOFSNfahBk3Chcy5Txh+5j
DpnMS9DJqPXl2/LE1QUPgbhSMhIQ5ighDu0jlYB6UySgGhqE4A6mkA+Bvl1d
E5BKaplK7ZhcCxBEq55bbqpgejipsY57q+bLMSStEYEV+IeYfwS51lVq3ztd
uqvcZ0TpjuJan9Juq5arVYfr+P9JFK4mYdFvnkpbMU3EQWJL4fp70euq5EQ8
quVXb3ZUQ6wXn/IKHbV4t1OKGSIFPEB2Ql4gPSzQCl+Jo1eVHyZqwi6aSl+b
xpICxE2RmiOH2+igHIcXKPGlzrVPpWf2pR/LtddwFVOj2Jcfu4qr006+vQss
DX1msBAjEC+Jb3qWjj5HOhvjhvQ9W4LlFgegln0Ie3GQItvnHo/aju/vMOiL
AdWLLGgWQ28S9HjGp7xNb4miH6M45peFf6uW3xLj2vms8GHHXa6pyXyKp/KK
DSFku6ZosKM1FiJN3WkrmvV5h52798zPvWDmBlafp/1BZeZkfach6eZ6ESI7
BqNlMr0Nd7VH9VAz2ienQWgyH2TaPMVbO8Khn3ekgLBH8CSbk8bzusZHacR4
ir72UFwJqGaRyDGpooenjo3z7n3p3CCY/7H0E9hrP9SVFM67yi17z1IYoNVn
NuIFD1Qabmep8J1lxsxjiMKOzkOcv8zs143fODqIr+bR5dbdaQCAuOHB7JCv
c2sUdORkp+5156TjDSUvgqGUpqjOfAjjrPJUtOp1WiLOtIXRb0OsKVbVwOAB
PWPKk2FsQe1NHiYiQ555FzkUNjF1/z3usBJ5ba3jHpA6wPDAQN5xrRbDNIvO
8dB+1blR4PzweqlNyNHFBQsuGXKcF3s6Tzbg2YQF59EXXqSow3vUHxUlFWmk
ojbHYXdR0u7bhYiFMZlW2RODiopU2tIU1oQXIiyNI1DdjyJI9phPHIZwAABY
8cratH9SGGlwAnc1Qxn05EYl+ggQaw54wrnKzhtwHo7VsckKh3o8OZbofepp
vc0s5+alUlRCbplhBZiJzwxTuvL6+tPbz9aD6RqL7PtYtbDBOIWigloWosD5
900ruYvN3yuwocyIdf6lIhkp9EeGXcr3KINupNHc4XLj7IIa55GFv0Ak6S6H
wVbPZQH24G0gCYSDjoLyGAFhHQUaTt9OD4VdCRXASO8W6ZkcSI+T5fvc/ebr
H+DmpFU/HzOqkhU9DUycJPqgUM+rRGr4e2azaX5ru9y+SYmIcj4yVJS0x6kF
/VZIyUa1JIxOm+qqQMOvyqBuN1GNMTJm216f/EBVwVt0az70h43x9R/0cqz/
R7EldOtvzfAuajV0S6wK/Lf1O8j+Sqxs3lepp3DyWNUtJfa5cX7BwqEw8Zf+
89YmD9oZVGj+4S5W3jnckktsUAD0RPGa3uxdo6AIf5MzQwqkpMl/niHwV+6V
Lkhicbk2CW/bht6gQFALpo6HsD1dyTWTTTth8tCeo40nLpAkxCipA2P6oxhc
hLhJo8keoXvWnI3GYlJHVJGzp+ylFWFrD9ZNMZzPzsy+iuw/X3djNyjNlZrw
FK0guYz0kBLPcT7/v/G2X+fVuF8B7Qsab5T69h+H342RxFpCKC+vYbqpfq08
OLdnSgVRmYxQ0o+z9DOrxo3F7nSlRU+qIsVu+TRFU4X3HdWXaLBMvlScEz/L
pIchSL1JO/XjOFkShWJ6/nTeJ4WsIpXicx66sFt0lc/0M9ZBkCVpyKhcfpch
VGHuwVMV9dbasBORc9/lJVJtLKg6Y2wZ7QoeI4wsAinxRQ00v5/Nh6fdccrr
5FfbNWeiyYelVsAq5CgVivJYLax8aLoPFnp0om+Ua0tHZYwMZ1Ga3vVpZsJC
WlRmcqjOk2zautnm6h9xWBGiesHwnA72H8dCOMDw50VmcGgfXIqBwgT311gR
7rhWAUAwAHp5Jy28BD00FLb4u3Ks4aAzxIqvADN9q23np+iw+ll793BHRy0a
I7aXMwJ4sRTSFmz/ud7Pys/ld2WebS3bkY9pqHm5YDmdU4QiOLkxgmhsFdFG
oErfY+tNwTI46RJUbVg4IiC0G+VZwii7qGYlHQAanBLzqEt8MCvoQ49haG6v
qbRhyZ9a+zQLJgG5yfk5FhauzHlL85hThiYLX5xiHQ3ca3md8K/NNBm2qmdy
nkkhmKdAPwsxM+5FgaOTidT7cyrqjTuehULVuKU8wUm5OBsr5TvI1MSW2K4j
IlhvUJhVjJ9H59k9WDk02j8iL4dxj2g6IlYkP4nwxKJeMeSbnm5FDuIzY37t
Kx64vEe5MlmvzH+jdeFOh/XTRPGmKMOlcyLWUx2ZZY9s0RUEzZtn7mY5cA0i
o93I4rkR7cgjLOshE2pqHJBVs5A8IW9UafRWwptMR4ETYunjd5OPuDWxsPov
dVhM56sx0kkXX/6z7N3/U6lnIH5myQHQudvsiYPkGzYZqOdBtBGraTXqUSYz
UPG/JnNiOmCE2s0cWAeppQo4xsEM3zb2BwTHTKVNqnkHKaVOG/ljw1PMa7vZ
s2SFZ5tpO2AbLSBi7LlHEgu2i8CkXsHIZLhEHtlWMts/7Ix0xSNO1IiJ6ycE
Bu8ETRB5IDxU3ZY2GbNAuyytH82ynfaetUmfqiekUzfD0MEYHqvBo+wGetmT
EEtKMSjWD/lceJ1RkG56GLj5BYsQlVgDPStRq0+1B1IsnVobWSOKHUcBgUVk
/2rIe1LM+jFVO7w+NTzIKvMA+9K5IyiktMUxjszZp1skGk7j5MnPakqLTypp
NDEBrH6+AG3DtcPqQVGbq2KSxQpDlNf4THXjUfQX+Bz0KabKzPhBCXuquQkQ
YInfC7Qmy/zGpE+sfbFWRnlskIijHezNTSTkGj/Nrjl3QEaTiz2yo8BYdXV9
i3j/uDwnqr/6j5w4mZ+yu/UQj7nhnzV/SDb8hafBmjU7E23J1xld7Jll9Owo
5tA0Fy12XLTi4rguxKVUx+nmiYnJiy067MFqe13H/wTJ9Xzgsf6iilgE29wZ
A/FL4lTj2PevaQhscrRYRbExD1TbLHv2zeSHSDbCR/V8xXUFcuCtWLBqxjQU
DoK2Mn/utIxyflkVcq6FKrBbpDGX204aYOF4qyrXef/bZ4Y/gWGxDRkusDTq
M/iHauknC96+9c/iXZ3qJZw56PWN4OEEgxngo/Me+oZxRQ12E99cNmjMhOPv
CkYOGcXOXE9bZ3NuaJOoDmP9SPccsaWVR19SgwajDQ0zXBUZT9aeWcPUxwyn
gTfyKhgvjzoeEHLnwPGGWagKdVgUPwlrfIK0xui19u0n028wYdcFUy3Jvtni
I7rH4wRpM1cHXQia+9cRyvf/9TMXISj7DSq8ksQDesYKvPAFoHuPKkCiizzd
x9Xg30oE2ey/yUvlPyIw0rpVbU0dKi1fURYWGW7rTY1TP4oWO+XNKtW4iAg/
vw/nhICzXKESDqFou4OY9EgRd6r79HBkWH3bjuZJEuh706k67l2PAQIkqXzx
6NfGetBWP4FEFMvdYQe1o2wPmV5qWgDxCoQykpGCMgblymYgnyV09TrDyjQL
9Mlh+Q5EKwvRi0ogeb5x8cXXSuicuTCkFD3jaZuaZgp9wSq34fGQEM0Gk5lR
qLNMIUTvjHczM7GAcMxfGjYLgkpS2b6WoIf+bx6JSaAHE0ClRPEO1FlC7PwF
gs8XJWawfxUNBcfbQ3zKTPu+QQV8/hcaE3/++kIxqHm4JBEMTodfG68TOzvA
QxdfW537joJBZ5rnTKylek1t7Ms4pTvwDwFjNDfNqEvD5lj4kb+wsHF6Ss2L
3nU7+k4PMbTaEvZp25RF/GqmUXBwKt4Rcw8HPaHUM3/CrqFaxiUsa9BE3OLh
/9l9vLRCX78U5iEzSLyAO9YcsgkuPMDCJSshu9bYqeBGqNhQ2F3EdFxTHI5w
Jg+HXLStMgxNpvj1gGCSExOQ4iUk7td3bBovlgcX3RZvNL93St/6y9KtM1b7
dfLmTz08kaiVdk9UEFVcGYEtqF+TGPArG3pu3R4rXRVv1ms0NfphzaqxF7S0
suEMjrLvyAZhTch2sY5VozYxt/tqXJnNBPItdr0iMe3JAuPaB2rJzdrdbn6F
i66QyxjoyExB0KuKVZFNRRkuP1Fj//RsmmvfhxABq57nM7N6xaPgVprIEZUi
gtVFqIqQGpUVo1QSFOZV28edyAD0IzOkWzC/v2l0cxeTJw/flhoaR0uHE4+D
7j5lO1nPmlXdWAsFOz9r7HdlGp40NXAObGqAcMg+B1vb69YCOjvOPaAbx2m9
U/1qhYnkeRcQHAaBagWmlal2lzzzwY2ElyJ9tMW05hHdWiogBDX4MDDudZsI
QF20FJxSQE2yH92KW9Ki/8RILpo8mh3WMB7l2zJHgtIBDtT+diCnSlwEFERQ
JnlURrCBV5uWhA54RouhbgXoW/7z8hrqxYoMSp4OnqjGPxFRHBlrxL7YNRuP
z5pljdLt3N1daGPypow4l4g8vkYPWqgaEZMFgi4DNf8WL5YE0Nu+R9Q3SKl+
iimY5VwgsPH+2lCraXQrF9urFvr4g8Qi/rt/I4z83gn+/0p97zt3x5n/xt0v
+UidUOOddWQasAjXjCRSpDYGRp9K25rx+sczAv49MtiIIt4zwHFi3piM8P3o
slJwVuCJIfWNN0ITfnY82kJtZAJdc3ZIp4ocF6ASZUHgMc2915DwXk1fMD/p
3eoctMaab9xJpAcNEWPPxPB46HKh02S9bOjzzh1WL7oOjftb4mP+AVRCVPQA
FCkrP4BoGyTN7YjucGrjdcGpYczcXU3oB61h8ur8bHSSf4e2gVIJaHCNsnmb
mSqZvy7YCM0qcxKl7/wR/cnWcyMmAVpXhV+2h3UVEs0YWKC65t1csEFtFgPs
Qef5alDiXG2kTaeerYUN6GA6gL1yp2LWB0mwOh4mb7MkDXGbrqTygXMzo7Om
8ctKEOROm43bITR9rkoRnGx/zwokKgrQPwFBFImIPIANTk+t4b4yyOx4Jn7u
snUXDDqobkE1v0D9P1O6levxm/eFp1SOSO4B3WCS7GUJQ2ddK1kpltwqBpMc
VhIUeAbKeXxoxu2vb0qnf82y0Q/QormKoEAFELJK14KPR115QKb315aEpgiW
kcmI3lvbByzXr/3DAV4naOeZsFG8U/0KpoO3p1RP6Ukgd83qyfyCY1PjlhUu
mVFQP6JzFKBDQVClH/H5451LKxl14j4jHgIR6P8HGp+i0/8AdOW5cuVefSWa
pavUFIs+1DrMdDD/hS7ID2ae1p0TM/zpAKMfrNmkHElAk0a4tdy+B2NeXyyX
im1jkykwA2VLYoz4gPro9YbDlMDa5TAE1AnTx0eWcAFn7jurwgO+qqDrOt8v
6RuBH+mY+oQNbezoPr+3TGFFlkWqru5/sxVWOzK19GaIipWrMzI/rwRh7LiO
/Wk2jzihupHrSqz3eoISPz/oWsP3VlJF5owSSIRKwQLX/S6ohcTZ1IlephRS
U836BN2MR2vorWyCtVmCxjTIQbkKg80zf+W0fGYS82jOtlbUKH33hZMxOni7
4LLTI878MQS0Cp6HlnUndRor1F5qy5D6qHnzMQHOxjmg4VC9j0Oj75CsSo4Y
qeHOoEeNGy5/D2G/byRE+nYSp+bhRsLweT2s+GqnyjTESNuEC1ieOOg/d3C0
Oaytif33jLTswn+E9GmOog4vcpuFBN6xeaa+LtH/FCHD8kO2hU8tZnvYp2cu
JfFD9Tv7wSwHWg477G65bImZzWHjBGEvtUc7F7dTJ/Z02EYGxNLpxEf9HKLw
RdxdBPXnDoWmKnjWw/S/vqpsrtmAQw+o1Vya1Alx1YFa45CKXswNrDtTbcfT
rCHkulOC4eqcEMBSa6OttuQAIOO2rHjp1j577aEjQKaBtmRNluPjAZwa6aCX
2Ru8BQBxNLpgl/zbeCiQZYM4FIoH8ZsK7EOhz4HiMV7d5FMchmpjplgUGNRL
tE7L5OX6jvqWEvAIiyFisWwBmnWfZzxsznhBGdh9cwZAbe78XfSGab5PrHyk
ISxjFCTGJa9is2lUAo8vuLax8e37wQuAD2KIKsgIKeCFyh2lPfMwuHlFWGMn
gHCtMjh0kdUwtwwM5H14HR3iIX3X5GFEkKcFdUYhb+xbnJzWJYddFf2L7FP+
Ob4RzsvY9CzY76DM/9TlCr9Yk1W6P9RGB0j51vlcvF9CYprmIhWT/o94YEW8
t8XzMo58PVW6XUgpEEK6PPR8Q062beQ0qImSpQ5Pb3xdc1S7kjWXSoj2ZLVw
iL0WeFNYPrq+KnFw1OKYD2lnBFIDAuvzjt6Tg4JiQ/NUaFfOfZ3Fn3/A6HH+
JCNqXS71CnEDfjDrVsQB6BnDi1vHRr4aTIZKOSfmWuWEWuYOIbILfnmn9zwu
OkP7JPEXEnVuK7fjunFBHlq+PRjma/4n8o+1IjzT4aEEzVVodFO/3/FPGme6
JrN4TWmj9SNB+ukU4JjICdD3F3fOKhwGmNRtPKXVRVfQ4TAIwn980Ke0wssr
6a0oLtFcjxIW3j/gBbEwYIwZEJys3DyoptSzzUTvAJqgQJVTQ6IMjvX1GlnL
S8O/3fmknC9xOk4JE4vZycCE3ichEm1Iscxr/waP4XaqeHui3pq5HGqA1YtN
XCJOin0Doe45Rt0e5PNbMPUUedto1AD7f+b7ouTIQ0bZ0I+2TQE2itiqxYVO
U+tUaQBNiwgg9dyji74u900u10STK7aN9vdd3TZg+8kGdRENhLcYJdPom781
Sb26PtkFQDtQwp2VXAnq2ljLWmwkvt0hbp/JOhEQOkfvzgZajFEGQvjkmNLw
FqH3TFqzUmATQCjpmX83hGOVnL+gqp0bcvgVWLWBShXjMgJVunXvx97v3CaU
g1wMwkKeyme8Y3AofrAL0nj2aML+MruyzqnPgN9cp+/BsFwt2kF7OwDdHcQk
N6WO0QKxiRcmLjSOt3NX2rJ2vAZAzAj7Z8locV/feSXCUUjOime9PW3hwNkc
jOC37rShWVaJfmE130fKaIGUNzol20j67PkFTKQvrnn4eAmdc3kSshALqtod
hCMaheQy2D/pEUiS+hfJb8+lTHomEW+06TCnNvB6seLn+LqmYdKpXrczrdb8
JN/6TT3eUrEwe5vylAkUV8DSPwOSQWPnGqd4i6nJ+lqAEKWEknQ+WWDEIJ3j
5fcBe3gatePgIzcbNzo4i6sr3Q6GVSKKWlnajK7/uKQmHo3KxCnbxgUbBqL7
DoDZWxhjiSej9W17tAKwVHQcE7IblqTP6g/K4PHqyktTM24Kzb5J5e2WzomH
b1uFuP+2qZIEhe3QbesJCHIkHPzX4Ne51UL6gdPFuzxGgw/v52ZoXSGn3YHm
OFaL8HE+gNNimmd9adPqSF1Fyj5nd4VK8QpM9oLnHJ4qIUSldis3ENeu3fhs
mb9yNRI7Y0NdV7KWwB+q3GTwigZ4IpgysbPSS7aUAh8d+7U4+ItsBgFi3p9V
FuDcqhc9v/HYZrbZjvojGq12zlEAagqYUkVZuOot8ZYRnraObisg+Sv9G2S3
BhqTE1RUDZDwr/Syy0sjPlJKitgPFOnUyLizyfzQpZMIz27UaONlSORrEHc/
fXWdANadLn9/1x3D1CSGJddgN3LsKcLOjvm56il77vWH/R56WQ8DFej7KH0D
nZ4kvaAs3F1zcHqu9FDT1JE2X+ofpqfLJva9buMvKfLmONs52a1jkcoY44Xy
uZvc0vuXZElxcKBMSGQMrnOadUygi0BBGiLaHjk1+/rWcgYZ4ZPdubJfUM+8
59KV8OjmffHBgUu/4aAVJhI+KuzG29bGZ9a+pquJj8wBBjDOD8nmEtYqfUVG
A0NTBg/HO9Ee9x1/NwiF+0kVJqS//VRcgXC1q0beLCCo3s/4qO258D/Z4K0F
8xbNxtEU7H1ApYb5RFq/zgHmubCcBkYfN2LfKQaBefzOeBhPgNbXgpjXiDQs
VDsvuL9K1q3lkXctYx0XwkyVNoXY6GPYB8ZV/tGpmth42pi6GsQle5orf7ak
12KPRSEWHqqXiLB2Q99DusImmsiWbkTuPQByvThmVDJbNX08/zexENVj8L52
L//WK3gNWcZ29hEN08UzSJ+UQb2iqDSpEvh5jWfMwVjqyispt5jpOcTIcTrV
en38zDrJw+Nk9eWDOEeWOZXsXNrVLD3RkpOP7HZqLE7R1MBhVYdVcqy9LQJE
y+H4ZZ2Wo7dYmYPyqKOPAC4Nq9x5ccA1UV+HJiS25lDmIOu2+zJf8aTsWqEA
ULMQhrWtgtfCwjQXHx4pEc+adHIN2zjpP0FvqUJLsC6yADVTqi45ZuaZalnN
b4uHstE1D+z/QkYsFaW/bIEzzEXhsNjdIyZPuQbuTDx9B/wXXAgbXas/cQND
WZuMEhgPDHuEQkSXheixNyPwR6ieW+2PUUnG2izZE2qRD4KR76IPbeNHKsz1
AkG4xFK0aSqwkGbIo5bEXZXif8VoRgOuhzL06wN+yx4IXIkv9ijOh8XYf3ZU
aeDqvjTpJWXCPWfh8OqEGEWBvwef6t3MGNL041l/3f3R1IVYaxC0fi1A0FCF
7FeukjT9OqABstV1/y9NDChFJAjTbY16iLwpT2Y5VBRtVwfTWoac5nAsptiB
5rdAb4OBb6aT+01iMilxTLkXZdN7ne/5/eoBoK73YjutpovSyaWY6Iz4Q+o1
luS4aXaRpZBv0bsUE/5o+v4H7VFQOsN06s5vcQsPloxwJiiz5gQllrs0VLXL
faHNUXxxVuxd88WdcNsAMDrWS+wIUAR9T0R2Th+q1G8fq+zCPKDQcrpc8KIR
v/iRgYPovQtHVVwBwJEIPhx8Nxudrp6wdQmARnrPkNvgCixq9yLCxR7OXu7S
vruDTOlVN5qyq4faB046tvVDyKvwebu7e+txJsGwY8KD3LtZ3LDIS8+Shh59
9n9FvggtsycDVnG1d+q9feB2gTDeVd5tKmYs0H2TlLGx1nx7IwaMc3JL2x00
RWWKEygodKpThiiL8KGcm1qOJw+yMHP47DJmEe+O0zANSoDt6D3Tr8ZqTSoz
EvhzYdP/Bd10zH6VqNVVF6/bEFvJ7lSZTw50l2DuQybpQYus9zeWJulYa5Wx
9wfYJf+LDqbTcVN07oa/ih+6Q5B2k2rYuZ0KNPv5I4jPIddp8vXyUly+KQms
aioqO41mBU/4v4IhZ4eGC4mKlaCmQ3GUPjW1YslLHzPoq7N6g6z/OUHZJ4a7
Nvn03q6lLflwSx3ty4FdPDrAINU/N9PTo0DcRuo/Yd8+Pl2nPUlrhmmvgG3e
Y5vRRhnhKjL6BtxUmBTr+O3HIHVbLJmm85+MpP4bSEjjUzGXF27W5TOK1I9/
oQ2RxuBW9mWcIxvbwU3VpHQTX7bn06js8ywnERXJ/VVmIHinZdWhzKqDD4TQ
q+n/QGr01B3oRr2mZ6ao5UFBP/12jFlxwet2zwnoCfIeTUi5Ur47Zi/W0zuI
vdHo927emvV8zh6dIkNIIbCsnJP73//PMTer1wbyCGGrBuj+FpCR3/J6H6d3
aRdnoHuGtOi2O5nU9bk4Z7pJTRDNtdsS1NpcXYQhXUtjW+BTqUYot0A5YoHz
Sx1pjyKNnKgi/fRxgctSl+kebkY39MZEulZIZYBxSzWrVQJWprlojrE0yMwN
AgJ5nYsWf5WjYwVxbmIpekkyPn7Rowz9enxgLR/DQbG/k8N0QaxIy5pmNQam
NJiMdA634h4EgInwswj3zKC4lx8FLcvngH0H2L5d9yJNBHxsBvxM73UlkIwH
4dUYYBMYt9VgQKKFdQKkW5xrP64JfeGeq5UNTvtpsVowTPoZep3+6PhJ2vBc
CQPGzQMH85WngFxOvGMMUgp3olxJSUb13D9SG90IPsdxjiLpY4e/zZx+gNFn
FuRfRknS1O3seiV/A3ngcyb1qmEAPUIYQoTgMWkwMDC2gnctn2KBjbEUwPQl
LZpMmPlc8XGPBgXxfny1SUlLwNLVKJQFOPvMOh5zWJpvKmJkvBDoGuwLIjT7
Wo7yq5oRTfTSBMM2YUjyGxgwtVn21/koLHshFAbJHO4irRedxuPlwvPIGEIo
K4Tbvrm+xcw/h4PARseEWcf0KTY+5BWyzLR5bxpnbLenLOrma6KHiWyUISKv
WXhZc0TATYZTqd5Hvnp3VgQSAc6sKvsGjyXDWyOSFy/Wz1d5egGbJDSzdQAe
RBT54hD9wlComrVgGFJUz3WxxcMH1XfwqqKqzkEE1xXYEZs2idQ7am6J4xcg
PQcxMWbpQRpxvt3xGrhNIav/iAlsk3pitd4iNNcM2IbQGerdsT2kKi6UkgOm
jmvX0kBtWA2pjSQyxahD6sUUcIniT3K8ok3G1iUD9MgN2AwYLx0VsJFgq/Hx
X7ie5kuIUZqAmeMTzHP2WYTSfPnKOCY4q07XZCnReKjZoXnkBrm6/20JGjaU
cTrmrjFlPmlDLUkJxuPmkhRC9UTzptd8Sot4QqCfVh5BV0IL6V8zrQ4gNVaN
E30rqBAdh6VBb5S1e2Hl/b4OOixb3WzjLrgSGXb5GK3EeSyAoWvIy22ZHQu/
uA6fFSa8PZfxXcJ/0L5Xpajig3Sgs9txInm+YDYJZ6OHXM9JvgGY4JcQ0Xv9
AWitHJ6mX7LRdH1Cj2TzJbfp57S///xDqQBepmmBjGuAtZBl4FaReUZyaT+k
j5Ik2x1yK//8XDGWWU2ZcTXlSw5SJR0YHJgQqsgDWpQ9YP4E48sScWqfYi2P
tBCi18JEU8AYFqCXE3hki+T876MDBKmqC0j89U77kZ/PWlbr5eeFHSSPoDZQ
9NPCDmC6j6vxTOxh2vIqtEdMUaPe0YXqchP5VUbEXnJF8vG40d0YKXoYr8cQ
CF/14BYeHCEBMV53oiCeZgknU7tUWgJeGZqk9CVlK4PAQQ3m4MS7XG7yncY/
JoJPuaZgIMJfTOtGA4kGMs80KF/4308eprkm+jifS1/t84n4vLZasISHS9Wd
vaWdKkG8mYpHlDeI4ks2xBQXhLNzr7tJRhmQmjW+Q0J7FL/PDU1qE+B82zFV
/EIk7r+RHyv4C5IzK/O+Fe5MdPJCp0JyPnPd9UbduYzYV4Y9ZH4wPPk5sVwh
2ZmPStN/9+yqyZF86/azQum1g1gk0Ey5Hs447jHFsWJz/5t096X/OKrdZgQN
jB996hdjUh/Ol6dGCOsUxhjn+aFGrE8YhGqneJmo+mWfCdP9fv5xc/bB3kAk
1lV4oEqtDH8dQ2Qur9RdvcHBaCuLBy16c4gamPa8I/SAsYo3JNsEBZEsj4Nq
RdjTDddz6WBIYwuAshaCAmUJvWXAIq0mZIRahqlJ2KeG2jDYTwc9hbfF+bsA
/rlUzVf1lo/GKoX1VfUxaWrM6G3szYIfjyhHREtAWTGooZ+MJIe9M4kpaiT4
iSyzST8tU6GO4z6+MWCFeWlfj5axdxj34N3ejr8I7CrhfJLd3uCvwO6AHCf5
hTRe9BVH+3F999iUnjCdVaW7cs5+7B8JHFZa1DgI3OXx37cJSFjJ9oFy0+rs
eRZJ5Zo+e8bAzAya9PXuVNZyvjpwcdcNIhyxNXATFAo/zlISiCeE+0zcZYwR
kxIJRKUgukuc/BXAYUuGCl8ZnhVALwAG3an+4522cOHb0dbu0J/eV136A7Hf
IpZ+zFGZvK16V8pCysOImWz0TIJAF1rZJ6Oy5h4ELUSuXgdR1sHSqqEV/m+f
DKTc5uXO6IWuHSFLhvJnP5ZYonAGRPKzyIbICP0MlCyRWYj8zGv1HtN9MAQS
f45TLWy4YwqCcxi+YQTAAsxUZj7RfNIkh7x0UPX0Tqlq+f+YX6XIH3/32r71
DMipiOl3Kx71mlK5wy5QAo5q6wlo4xL3RsfsgOK0pKn/IB63EGTlg/QYJbco
KA2pFey2xdgR3rSC/gLFMILDzxStumJ3YfiEBHj/zBHagaQmQMlsBx6HgXYK
slqNFsKqF7TOfms7hOLQmWapddh/lhF8Idx9p6W/WWCSRCSOckGwMNBofk6n
VEnZYn/U6d/uu6xa08KjhranEX4Q765MrMadGTLrUzSVRBoximOmKPRqh8rV
4bcVBjJfr7TqBefkEiRdcuuctdSlmmV/3VJ24lRVuXXj+EAL0mWWUBejWZLS
mHOF8deWi+2ZJ/AEip0ojFIawaxHdSJ8ziPvw3Rh4wnYaS+VrMYGEJ78DiH4
gWpMiu5mdw08YguwNMdYAmMFnNyl1CByxyf8n9xwLIHycLd6tU1Rejm2UL/R
zPRE+oOCs5naxoVm482v23JHyn6vQnfgCsvU4g19ees2qMQPshLBC7FPXkBr
SIlxrHdwipOEPLhst/dwIkPJtvzojIL8JuuIDKqrO+DYskGpe/Jrw6aPov7X
LqrsEWhRft1Ds54RI0KnMhG9sQV9mWVK5MGJ/bRuElgpOCvfhvnwgLSlebKr
7EQBXuGk/uOzkpKXeyTr40ge3knONjDqMoZXRsWQOYKqNvHVMC/aKkEDu2li
zbu4Zj9e46WrFdLP+2x2tRR1b9U+hDdkLJ8E7A0GqFZ2VExvRR3fuDV8in8D
eF0ZDNQ3o9tBx/iV00NKTUoV/WY0BLxucd+T7JZiFzzfQIBD/tOuoAcbsB/p
B7VrElc7owTClXsOtPzm81kGseepE915qa3jSOvPd850TMqEAbYQJanewqCB
BJC5e0lW3iJ36gpSP3v9IXNl7Xs5dQUb3m2IbZg7rC+qxXL53nSpm5tP8qm9
xO7s3E6fGtotgwrJ73gNoJh+Qo4iCWhwwxPTpxP01+l68aPw2J0q/uBngaJo
SogP6p8aAi1YdlTHQvTOreldk6JZu4gK1pOKD+Uu0xcBLbTe+b1Th3qdeKvt
AxDWMIvc3oCxd+gMFUIY54D3Az6bIcReJ/xj9rI3HAzBa1Bk9abUt4/W5CvE
qRgrtWvEhK/Y3lVLpQhCiXuXQglImIwPTQzmnYnYInmF9zb1tbuRKGfdkSWI
DHjOIaZFWEfy2+nJwh+YSYRakDXvUbV5M5lIU3LeXSiFMBLJXS7ELfzFf7qK
+UWQ30WfckIATv724HicrRJNwo9CpJwJP3e92Wlat1V3Yr7VU5NMrMjhNBZb
4b3Ved55vSnDq+aLzRlJWQqBL4VvVNthmN/a4c2WExoF5iloUK7YtrL721+O
LgjybTS97/JDcgPAdWLH+s7eW0SCBC7OfVdJa37KfjkkvZOOzO0rGCx68iDV
GFpW0kxRPg5Mf5hN/Gc/d8EmjDdhutgh1rVy9ssRDNVknkq52R2BtnQiXnYm
mprwrJakDYgLDvAsDDgLEJvHaRtPEAKriAs3kCZ3LI22i0lZoo7Hk5acCqDc
ZDtohkxuLmq5jmUvCk2xmQ+QoQ2kHS/M+ZifkNbPmvJjN2aDVoBfsHG0IMm/
/Pa9xIMG8CnZhP9JgFRXVLh9p2oJ933ajQaj3zFVZ60utyf3YPzPWhB2t5dE
lC/cuhLZc/o9inADPprou+30Ff+sLL5tnOMrlMnUez2zv3vQ3DjtJxuQyiQw
/wIkBF+KSCg0EhAuy5sZYLzo2lTMlvhHbrKrrtabSXD8uwueA11r0MhhIyRH
z1uRmPeXIQKIXkdvPaY++tqf+d7/W2QErBOUvOF3yzijHScNT+BiJyAIMpJY
91XaQC0EMMLLGQf8e0qFBWaOI1OqNd6u/8cCITsku88E84BU+g4FRKV5iYkl
DvgzZkx+k9pRCKE1rUTFHvcawGvW/llAqDuPLoRWeWgLtgMC0dy03+KM27dV
jjispYE8c7zJLNjof9vccrIsMem307oVMIG4rm0poN0kfW5b4aLMU+xv/5Fs
jM/dCK/H/E76SMfZoOJMxOG7Zukc88gZBEHVMM2ejdT7Hiez332HGRDkwwQs
JZEoHb80J3DEVNuSzQemXtwDXBp6xNPy66DwpcfNn1ayGoYYSNC0bOtEHq1E
2NXwTrNioflbq2tKYa2Hc8eQtYhPR01O0agJnfqPYdNiG0UGbEeqboeh8zx3
RkFqbvCZmHFTJQYJKPRbcZ9H5Olr9P2TavrFy8SipQSTKo4HXzwOlwP9c9f8
JfH5LwH0TcdiAvUVxM5ocJ55JxnBYZ9zY3tAxZsO5W+5JbeVy8BnZ4/KdESB
pyks+hDgqCp9MVWzXzkKzMaN9Y5BOpKefX0eMzYZmrXVo2kzDHS4ilVj96Vm
aFMUHygM62gwoQX07ACzFTmc/L5xJUWySHQqqMQ+8U+dwu06rRm6hiRyPGeR
7Nz/MNSfkH89z5b/5CuS+FqrOpiEZwfnMLLRyTb3VlAB/gHGiTQOV7X7OB8l
aXgMUUgTJYn0DfB82F8Ua4dsMcv1zeCyyAeiL/vBiHSTuvj6y75pC23iipbo
YfRdJvtHrLg+A5DDKxoy3fsrwiUaJxjQoYPAy5XLDf7bxXzDNbx4abLgD4sy
zLWA+gKWx0rtg4oBEcoeaGL0DaCU8E2ZlDqrf1zT+t119wCfXIdTkWneYchN
CB/ir9hg7mP+wnAATUzlf3RZ7EI+1JGiFTWrjhDO9Ky6HAuaCA+YRbZXhSMj
2+dCGrOUBef+oawFoE/ulUm1i3nbRWGmMsIemKV1qdggk+yVEZ4QkNeLtxRE
Uwfy+w/T3HmQu+xA5jrNoRvZsEYXNKLRirQS/4BCfg1C6kigtQKoLZFaMVI5
cdcaal7mvOB10aEe+1qYaZyzf1rgokXzTL4qNkw9kVBd1VLVqzQH0msCHjuC
ExaDSmaUf4g9e2nzXS6vluVd45kj60f0ofTCymHcTRdG5UC0pdoBBKJsze/Z
Qs70X1GnuDpqqrYRwoV3huwo3hmniRvFjc0EpN5zgZkFK5SZbTZMtLu8pzdi
8aEoxmMEuP5PirY4CHHCkwENGBadUQOpdgkFmjbQToo1YOvUD8/gLpv7919D
9z31nngvJ+2kVzIESdyK8DSmhTfqczjm2Iu7GYpoceqj4Lmy4QmzNwCaMhnr
ebyEM2McmvXKYwh7obBatxTqR7UbxJk8Ss+8ZnLu91baSLBiNOXxAG+bETrC
hCOTHMIa++nNsoIe/JvU7bQNC4MWJI+X9hDovwHkfB7YijK/+CZ/Z9ukVKCU
vXvY7ekWdhFOZ3XlS0erDXgRde5tYoXyjKmnkmfxtTfllSnmfEUYYtX3Jjd8
LcB8Z7k5KwxN+D5KgscfVei2Q1rodXQQC0vYzB8OO4fP7OB4MXsDNaWcQ4vV
FIMY96ZZwNNZDfOHeUQv5c5c5mPGqQIwxUAhXSkRO0Bgi0WwgT7hGX4aSFer
KsUmsb+jpxy55SsHiMmbP/IGS0yrOYqwnB3qvNnt96CSmEsN1At2nVzt53Tj
hpRkDPPARVyQJFrleSnaoL8b2+h8mikZSo2M9Ch3t3V2k3mTOyqgkHoBvYJt
lrfkWLheQIZzIosfIAmRBR7c+KHiu7YkOAqisy4HIIU+TYfvAb0XIJVzYNOZ
zKaCabpy0MP3sAEH5q+1DOvvaGQ+w/BnsPHbXxk9a+IKoXxOf0ZE0pVuaDiU
sXsqpfLxEFjsLC1OC2UxfSIOUQ3YbqMboCTEMYhdHfFkchkqKlqa2ciGsK+a
GDpWGh1Fpedl+oUiAJttaLE/yHMzzszLIsx0G9ZONy/1nbuwLsHE9m6z5618
/Fd48ow8pRZC0saL8lpbmlQ/JtS6Pe3AXVIOCjBJRLticgpWSxw6WlGYW8t2
qzOWPJdRyXy+FQ5V18MDRjCAhz+BTX3oRDClky9JAf8hxu59sNMNEmv6EWMV
8KayZQtRzyFe9UaTUavuQmw+T5mbMKJ7mYKWuP9dX4krjKkM6Q8gZbzi6SfR
DyXYM/rCq587fGL7kW7/87oVMdHUzxHOfaZq9X5L6WyebbcrRlsucRoahIRh
ucZZbGAddOl8X23f8ZHIcn/qLJxAz/zQm2ZwbkSmTkwlJvn46+SudilME5Hd
zSvB2Z2WndFs83hYZyzwwESynirUz4nkt7HZPda8cOefEZyA6i3eNi9zRKb4
3vansQXLYLwsDBe24OOfhvJBerkqmrz1QBkE57lEKdDyBKKaTStBB2zhQ+hp
tPA2BHXCp+nDWkPj4bpTJ24txLroTwnj9XxAICBdMQltkXgtuu4kUaMPXQRO
syfyjYVtnwAjpMD7FUC3RTTugqON35CMUsbTFmvdlZPCiYHwmsVyUo3J/myt
ItCM8Vq6trS5/ku/pydTU5NOd7bHdAaEiY+glwBUHxrU5YxrCb+WlRJdvH8r
bxExL1tBB1S5kVfP6Ya4QJv/nH8lDfrzygFvR7BGMq64rqH5UMnxWNi6dZ2l
bWR+fLwOezHkg+a/olFgbiCc1zViujU6BSN3hyKplw2KEkjovukbdIvdBrSF
wTl7MaxUQWvkjKdpdMHQn8yRLIX1fKjqFZGBocioo/JjLPNTPY/gbW1DGnDh
6TwPgEVD0EhjmTmmWX5KZM1wY9N5vRvorTLvcaaienVn3/+nztEUObyPDm+R
gR6OJOAORRi//KWF7MvzEp97hLalD46ZEX0EtzyPxInAlCA4hW4TMuTMxcAn
I/H4qk4Ii67efeEJtUv5dnSWlVJrgCuC4BUrv+Epl4K+aKldNOXSuoxuK9PO
hfJtMzp2rf36uH5oqN/XZA4bXJHCMuCqiV0bQn/GeeLpuQiWCZelnye6Jv2P
Es6kC3E6l9C+7YwgAoXFSHCETxivGthsAQNXVEjAz1jiGOXRnQ52mSxCy2+D
5fKGTa7m4HCRfnS64IqaYVQKiSOYtcXodoCQ2c9DvQsbjsuVg8KtXRT+ndpH
5HexHRLvZP9lGibFsh26NMFP5u+JlOTJhMvBZ1SKY6DTxi6BbD4hISyq8APj
jDYGa/wSiiXgHxRcvfYcvgWEWY2MZfwO1VJPQfAr1qtLoyGY1lkqnwU55dVl
Tr2NWK8VgRcOnlLCV4mxYe4HwKvnVWLp4oxvggdi8fygp00Y81ZME6+zNqUo
U5w0uokvxDKULuuQctnyT7IlGNQkJnyR2eSeIhFRFl7GqLQQHN8HjqGzqrKL
3+KU0ZiqP4kxMKh40JHPYNje+zH4scpQc3FCXcD/6+yefvBxamqAw36dNINe
vx4bs9JmzIfGhAEZVlPCcR5Ze4DKlqUWa1H/6cAXJFsbI+iXNkB7wD3nJf8x
dwxgho1svXDUqdYnWsip/0XkTutLk2pvYda/LNEyyohfmCbf0h78+X5OqJwK
VBdl1vBb6JM9QzxzVB81nycqnDWUhA5bSGRIc/3s5jDlf6epJT60JrXAAkyO
s6ntj9AOGV5l8PHVJz+MR0oi2uEfN+jBcdbPuLnRRF+Zcwbz8MtC87jgFfh2
wK/t4UYT9vkocn8O7Pe1hHKnFzf6Z//Nsk6Qi9tLCxDz83iUwsdNs6c0bp9+
bbMY7UKT2rI26ZY5A5PbQxeTJGPmDSmtR5FaNVpXmic697yhoj/m1X01LZuW
wTL6AfwvgPbrpQ/idTjxV9Wpo/8nJxJKU6Rqu9dkp0eGy3EK2909XYNt3Rgf
XpCwxsxeNKrsjZ4UcJV+P1XrEzrb9SXoP8LoYccdk35BgDbx9mQy/RUrG9mx
ZNvTH8ANRE/oAPmUXyC0pbjWc2tTIuBV1bDAFZN5Mw4YLHPoZkeLHXBX4eXD
4tkZ/xkuJ5s/uSQGUGllyvtAMmx4gqCy42vDPt4TvITWMxdwUGKoWXTF0GOO
Y3LdInYIL1W4BCrfQ42uwWuqK0hGwDPfSkwxT8jspBv+zR+kxR9H9c6D1hwU
mbSYUtGwHqGWg/U+CFhrxdSMXSoFdzTDb2fTc7b3XttO4snBEOzmEsDw92PC
5L027w7EvWRA/oPgQNU3+ZwJSOrhxTJeX5aHjszzRpxxQsVDIbEerQigEiv5
61VbsvHWQr62i1arucV3REdazVFbQ1bvgP+WWJC/yJHMTVkUuQg0remE3T6H
IQ33Gbojxs9fCoNq409oIOWCNFozEO9+ROiHEEyMlCTXu7vHNTS8FDKCvynU
8HsRp6LmiNVEJX/MsQPfk0GE5iuwtoXl7jX7r1XsfxnIaPhieJOi2sV9S8G3
dfLnEHgW/gMoA1eDqj4BWmv89cS7h2WndVjtp/+ynTCKk6VA07dYLmuQtblM
YWJx/wCPcLo1NL3/JrYTPPiQlnEPO181UIOF62XLkkfBGB/fDhI6qXqhS8EJ
AOolOR3Pr9L03uXvKsseLbjtYHNqsHhMalD8EfTh20qyImfYlk/RqLPGtSx4
SMfH6vfBVgNmlaqCxBxwBdoSKaFPQvblLyNtVCwCZSl4AXTSkx6edozs20B0
0XZ/ttB7OF7d5PVpzyplo9it1rIKEWkJIBFVn8KjPisLwHcsPYbICTb1lLeR
vKwc2Ac8LfFJKnC7ZU0TZB7FibatIJbi/JCcWZLMnzneGfoYB1/vhzedS2Gd
0hI8XKuQr+1DyvOcrs2K3C4tElbECeAczD8pPQH8Kgc5Wv0sdPTQFIizYAC8
UgABNbn4htqG57Pfb/2mrwFZPKydV39LO3TDTkF9kbqeyFJafbysM26I4lBg
EaMVecIcmsbXhpxB5DT7Qc8zUERr5ziARGjWUZ0hoSnAgZ0eEXUAoFQQ37kI
9Ea+1bfgbHrCgC6yd9NyDAO9gUNODnZYt0H4/vdhrKp1kl+DzimOdnLuwHqu
K6nOpmK76EjEFro/ZafAAp7k0fJjj8tsYdMxOZ5BOiPVOGeVnqRBnNWxIW/M
im4C37a1T4V4VFIM3T1evTpy+JlLRXlaWItH2AL4zVtaZYgSO0wNSc0gb7qb
saRQJlcRR1DehE7roUfvsx4oaQlzvKJdIkkSaAwRW6v4icacNteH9DDtQDo4
Hx71js7hAbgsZWrbM5vyLlgolGFJsQDccAuLG13T7W2JjSAdRH/JBQXzdKMB
j1hPfKZF1V80Zr2mlBOBA/71j+W7Os5K2gQhCtVzjAOSynDJ0NpGFr0ks4fa
L86ac6J3YxJH1oT7bVgOpNPeYfcrqtSpXAzHv5UcS1fDHaUB5PIVw2VbYhAB
LY9Qsx1LVdW6bdg3AXAFN8a1qAD2sFiFro1nDhnj+BqbhMPcIlgXUesagI0o
wleNsisbP0dUPxrF7pv2avzA9Rar0Qzr/gwhzDoJcyvZi9UsMT7qym/XxNNh
gdYtKWtZEj/EnzJhfT+ALChmXOiUx+Xh3/ZkfJksw2HZ36gFxp4NSbPM28/c
hubm1kur9l5pUg5iJYKpvCmH5SbO/Vz9z61VhA5Hd8ZFOFf1qBEFPajyO5aU
DdHEum64wS8620mDaR/LChG4U/y+EECHqWdhSNA/Ilftt7ug5QrYffwu2o3a
JKboJvx9t5/FqWm8WH7oY1iK5iwscqROL+c/hh6ajiP7k8steVqEhIbmlQ0X
9jnIBl8usIyDc4UAzrJ0Uvkk0++qSVWfQEwSsPSUYtI9cI7psdTw1azK7k3p
+qPhYd8gpNg2qOKWsTj+dlJzy2qSg/hADysk3OosuMl9XsWDInhpWKhbP1xr
EEVNpXDaaM2azN9nb49qawhIGNZ7dqEc+OdZoQziOtyMKupRcm2n5VTO82qp
+/A36ltgqfQ1hgV/fGoTCb3JQUfniTVSEZ61S/TxnNci8cL3y01xeOAwvgVP
ZPvEu7q4v3fBAV5A6CIyvOUoJvFlz0P8nXKC2WA5yjlLJiWdUQoZJimvPqG4
4piZymb6S9WEbb+sIQSLmB4EzNYEP6xCovmkP6zs/yF8aT0DoI8h45JPI12Y
vcSKTt+itTUTllOUvCyLzWugTvPsEXauvC+lT83sVImqn1lsZoPBc0FpwxaC
HeySRWaPdMYLZ7YdggQ1OJjDSyvJq+W+bdIntiRDsWeyjPT5hPfs7ieMWknV
4Ot5GHuvrTLw1JapVWVI0nDMrAgp3AD+cpEhrpnXfVSpNawIMLfYR9n0OQzG
9OZYblKbabHq/80/A4TAU2xLiXmEBSLkbsaQHVfeg3y92aPz7Hz8XpxMc8yg
w1nN7E+gN9TFiKT/tC+G6jkxBUxfajIF+h3PSAmxB/PIE2eTuHMsw9032PcR
JBlWeFP9r8V5mYG9exZirmMOxjI1w9vS9Fjc+kwcEH+iSsW4bAUU0frHkzwa
l/W74ZVApIJtAw/BJ9H2lto+35ELDHWkm5GvwxsWWIqKwTU5nJmfEPeCwng2
AmoGdPZc5wZiXB4RXy2gchkAkm8vZUvisAlIFMFs+x8JdZFIKHfTujg0uaCf
jkf9VvI7Z31wf8IAh59jsq/LGfYWZpd3YCfP5HSQ+MDeU9Kuwru8ZP0R7F5E
CKfcP+BXK9oAcY2Lxb+xBpgzKuFS6MwdH+gc3umOGlJm678HnI/SmV7ixWWQ
utYt7GEWWKIsJNbWAPP88N/1vuvFBpaQcUzER8IvRHk97+iU9bK3zHdXHL9o
s3SnfJHbqjQRxa94aYIVnU+Uhg2UH6EqgjIpkAE5Z9/qwG49qICdFVHtkw8q
6Tf7K6etYG2zeI4DYNn21r5wh3NBizM1gaUMe3wnTf9+qC8KqQuIX/PlUAwf
C84jfhGX1L1NLyVI2s4K0Zg+075jkerRMsgztYkSHjglC2vDgoFu4lw6dQyV
FWKIybqMUNNj+M03Sud/jcp650316h9Hyscarg9+DpBROosBcewaJd+VNgv0
oRlGzQOXhSkauYhCTe2UP/8jrX1GrfChkNlaXpaQa6Xulm4kxY6yF4zExcTa
hUgv2pPZ90S+WW2g7pWj4HWVrCJ0UMte2YDTRTFKAnYsXQyP4kqhmJVaCDwF
Gqhpi7hZIA39FG9/NDwpNkKKCfeQSGa+5KmP+IBIM5j4YwDVE7GR58VrDf+e
EmkqUPF/6UZu72ibDXYddVZkkjDEDM9C3gahqhN9J3XowkZHli2eR+FtYOcY
2J4ppVRtU1dEtqJ8Sdfi/6mXBpKG2W9NADmy7La1lJ6W+oPVQNyd3rsB/m60
72DoNT+xBCqZexx5SeE+Jkw8Dy6ObuJs0nM8JNc52Nm3gd41p5WFGs72etqK
jOzBy282eU0o8/lYrDUCZ/mI4/qSB9TB6uhjA3nvBeG3vs7jIdVnBn1Q3CxK
pdawZDlRhkyy72MzhSoRwrO5q+myIA+id7qkWzMC1Pe5nyB8rtSQFVnYA2g7
jO5Ek6VdBs+pcZXIkAIhzHfA07g2zzG6/dJiRdHbvNYWgDQEPm/Bp/nBnbK/
kE/E1E+jBhF517fyxf8ZqavSPXH9UxMcAdbu1kbv1aslFnKo8h5sN4PUTbYZ
tlIWeFmTTF3jSktbrezu2TXSFqpi4ckCkr27W2McD1P5jTzrzv2pZr0JWI8L
/98eo9b1yl+GZohYqeyJcC92LKLi1hgAPxfQtVy5we/zeb2wLhxaw0fWTyiS
70y+jNbnv75+y1/yyrCBkGBKpgflTh3Y511sZ78L032mEfwLQJhOCQGou0q8
11b5pAno3Mdw5K1zA1EEST24YQN9fFxMbWXHUGHqwhL237JH3HVoEm5OoVQp
CY62/5EIezrqC/EcO6lUqSw4rnIWd93GfISUWiXN9ZU0arnjd+JCptRX+mO+
/QABl1PYJiIkyE/X3BIezq/k10gC4nAAxCkvYHXJMXDPQRM3ii42ct8arIiu
UtVS9JblLkQMDQQ91M8MWnIesd/KtqjqIH/zMo2RPJFcAzR5a1uMhKHzEpde
v6SZlcB4FO/0kmhdkHfc3K06BG+F/KNP6A91gj2orsOxzV1Wu0Auu1Aj2bVf
NW9RFwZAM/bAEjxi+/vQO9woywRaiM82lsjSE2WFtyenKC8qs1YMdPhoJIXQ
7fQlRHs4Y+eHYb3T/9bgG+DvO67wqs8GIPrhYM+lcNST71DWAuJSE6fGjz/7
+K6kCT2v0mBiusLNZl2Qa40hUM9v2oekF94foZl1HiocqAmH4dw/i0ZFjcln
fC2JaSYCCnM7GKUvBi5wq9U5BktDdz6QWoZ1nRE5d6O6MCX8tFYzMt9NjTde
S8XzCMeVvPbo6c9LOwRH1JYBmgXmztKFEu/xPOM+uOOvXJlm8yv+LwInl90d
vn6JHsgLexoi+T0L/zKm+Fy+hvqGBKmliHDaIL7u5baGh+NbguA2i3ai8RiI
T+XClrXm7fvoUSalOSMVNj+Vdau4j+waieiqpRj68C8m5q7zyLj/mKBms+Tw
tufnQAg6zk8CC/pLOjE6akMrmMahwajOITi1X/P73AgCttbbJqVs6WfEZIVS
0cBmcRB5cSlMbaBL+0jdrmPpOlX+P3eDdME1qFzVcviSzxy4aeCe12CZfIMY
T9r9VspSP/ekjJCcidbN438sZiz8XBAfye00N6NgzniShqfh8lDalcFEMDws
KSzoOTI4APCKtHc4L3mYlBaPWW9/OtTdhh5eoE9wgGkRey4KMDclY0F+bvJ9
QfhdQHiFstTiFMGxvybucmWDC3ylNE+p8j48S0mqOGnOYth35fCp0tZxqQop
qYsyvYF6nQ4CJZfPZVt55UjaZyFcdEyfQ0Oarro6/p4F3VSIZ95NG+JIkOtv
6uaOta12P3Wk5VPZFvzo6Zy+aXC4Ix5a0Ao/83yM8+TIsAS9UMy/884uNNOM
5ijSWuxb3/m2jryvkUM8wixhk2aklnUvRqxBwrSy5bYv3A7bmjyVn1k88xbG
RrmwJhaBnI8C/ZAupJE1sqGYH4/DZShOebSiCo94qAg5pNdvVsvYPBeSBiWa
mWTVT4k6LVNcma3JuO8wyxSgJiEvjP0pdZsxh2C9vBYNWvSEhaHBJTXgekXJ
yP/8mMUoKURXFSFQQTr9sIorsvJs89cWn54usuVKF2J2zvCPJMh42psq4UKu
WlMjKFjjx5eVvigmFuZL+7tik9gz1sWM9lzh7FInNJvedIKhYhf2cQDkzmJl
1utMT6FgxscB238+o8nohY5Y/Lr9Us2MWZxyVomD9THjA4UnIYL30p/ynWZV
+0z8oD/3255tqKPBeKqQjFZ7kUFL5WGqnBe4FFRJtXRmjIqIZ+d9feW9/E4q
cnu5ghaptqElFyI6rTJcyKiY5CQHLJBnF/VzUz6Nf5lS22vfiDKzPknWYWJI
/gOVvD4U2atexPVRddrPAZaDCi3wSc4Vrv5WihDB96MarwSxD2JYRMyumrdc
k9m2EXV0r6X9H4YY5ELIwxA9PjPOHDR7E+7LZRvweyuN6jQZbsCQSzVfuxP1
bK59pQIU3+LsxR+2MIfo2MiT2MeYFeOuzCN8h9TMQkCfhZPZiEXf8ByKTq7H
6i4cVQ8owd8BY8IT5E2A6NYJb4LrtiTXxHlIw21ZwC02Y4hhtQDBPs23DiZ8
WXTqWny8DbB8xXAtnccverMDqO9PxrWwJxy94VlMD4OETx0u5YWClrFzt7+n
/Mp2Hv2I9NdHOZH2k7yuctrt8gAorKAeiNiwoEK8eUhBAZ1nAL7y6ANO4LeB
wV5yJiX7L64juqR4pEWWPiWlkhvEK4S5Sa+IvzHxSCMCGqN3g8ceohKL/Zkb
iS5dAmZkowwSXptn91KWDY8zUxAJC8TO0PQDMt/OZ14mJ0/4ZQ3aLAn3GKrK
AGzIaL/hSa+QVJCBgNmZFSIAyGorkY/VXaO6SkAbSA6eShzCgbenzLQVFhEs
TKqJQLWzifLVPOanDYYZs9xz6LDiu/ovRxwwPijgPt92jFLZm9CekkLTi/ic
G0Zot3M3BfyIjqppshNcQIf0IoJji1jEzxTj3jdSLvfRdNRxx5b6TSVFXpUd
r/SZ0+RZWfa0HaJZDZEMhQKBHV0fFBwmLGdnlB+h/ccrT9UgrGrUz4Xr2aBN
9zQCvz2fypnAgUD72QQu+ZpCPESNGz7tQpOKVq4j8n96EGMsMHOa/3yezPuM
o624z7yhkeFOzFpO8G3lCPdGy4xNMiKSSdjGyViQSGiBxvQ3MkTX5NMEHKy2
elwxu7LFaXwy86sMKDF11YZj/pxAF298BzRjjDz7T/O9trFZ6sm7AAADXv5C
Hz+Eig8M6Gnb+CunoJyMH/xCPUPbSYN8vsPhUgSIWxfPEt4wcoER4WOykIVN
3TOBueKnM2JC7oT+kQ5FG5xFz+g+Yot6KOFNrAYV5JE9VcnOxjsJ1u+0UyVc
9g3sDqoyntqqpfrWuUl7+FWlu7kzJmDa4tE4wbPHGBzpbZcS4vKpsbpZGn0M
27v6Wt8jIDJZAD1yKtXsJ4eSIfUm6oituXUx6DMnJDnD4u4BZ0NYdIW59jgZ
mz9U55aVqqp3+qlr9GlXRe4RGva5rIifdMZFCmHjzzMrbBu38wsqDiQSz9+c
7QNvidB8r5qd9h0SbdvjazVpxWeZXR10YhfaMHSIK7J4+7lsaYrt5VUHckrA
madyHOOUrH3XnMlHdzJTb9ALg71Devm6uWTul3m6g1HhOsvsJaT40yh16sU7
XNxnRgRsR+y10Rtl/PVIRtUhFzFPCD3qjP7X7hzS9SrMvOb1QrIBajg9vTOW
LQiFeVXL/aoBKP458GhbTpfv1Toc2Q1B3evuqpxDHd+qQl3Q+NqTYR2b1ceh
CPt9F5z5rgqot5Dog4V19AEYCjZJKD5WwQKGOATJFL7IEIurpipLeqNKOe5t
RsK7/qLnXHszkFhY4G/ndGL8f/oTnbHZ77OregU8lSiGBS/Yivkpaht/7ND8
fi1rzcIwo96zxDQvJk0N3COZV0RPAov84ZLtCxaxQWelk5WUnoA0kQq3evks
533w6wn4QX5md8COiyKcO5SIty739O3y/4/CYHIVEpS2bG9BLlJbJt+0p9qU
cWToc7cl5Dw7ct4TbSIx7mSgPI+gScn/FU4yJjaOUeJnQ6DlkexpsGEIx2qy
xyEfGNHGgsYe4EIvOyoOcg2M1tkXaYhKrXSYOV7J4zMt2tWQ6mx8rk7+zmq4
WvujXLZNg+hbVduRs8WmDH5/zMm0u9hV65EauDKXw2FJxSQ/4dfSX8deWSYM
XJ68x+af/sp1UhpoEurkXvRVYKz9pxMrAIB+GQZ7f0JMuos4+UmfAr0eWSJ6
EjBlmlykY6eiL49mxlZ9P/c+ZOA8nDoSnQIfFV3D0OmpFVLjcYzHQ6VAQDLJ
oQrZJAdgYAG8KmnOS9pnjhuJncTV2siPKD4ACHCseFyISYJzt708LnPHY9ux
FD3X6KFqh3viaojk6M0S8tiq1y6e9Tkq1mH0X0EhwL5nbrolxtuaRoAOiCer
Jn6czdz5TeJuXuMTyVK5PHuXwFv38sm0NmpYEnj91J+2OdJvUypQYobMQKpo
UHX/HzYnJxR/T91/l492AVzvdrG1yaaCJnkXTdx0DWocdWUIAIxx0wQkI+w9
QBuKT3ncVIlJ6oMPHYwZ20xX34h4h+Hk8COXD86TvhuumPBKaC/gAd4rmJcn
Two4N8lYJTCf1f1VGxYER/WDfon99WNBD5C33Bxux+MhsvSbX2vjz4wlh0TA
mZUlMPwp9zLDuKKNaMN9VJeYeE4DIkyRBUXqnyquhtfyMZald/HseMXWgkiY
CNjAfOTjellBj7KEZ3pXFJn+U1PFKoF0RtfakPrJPakeHQWube6Z1XPTdQQZ
BRb39qGSCjvDJHLuP0IyqxKt9gyO50+nQ2PTeXfTFDICIKZPpfwUkvdUH0Dl
rZS7DbjBcdsQJA8OIvevRFvchSQSbrYHtd1qs6skQ2NqCi25Zvd1JoHng5+F
94e94rvO4X/1z5ZpT5l1wp9Yx/GlIgvGjgcmEkVCdJS30Y4C1sNoBWzXTRRw
/OPclAZvkFMxfqBJgeCf00MTtVhLkEboYMdcZTACjqACTCxxjFWRdtg9eZ/o
w1axlNErkTEy1I2e7uSDWGEO9Z7Eeq6r8Q9vT9GLvZhpJVXwjqa8FmUsLTdE
cVNUNVxXlMbwuo5KfAQl9weycZXV24vctj6EhItd0ednYOs9JhVURbGBydrh
M5SBVUWgl3em96qUgOdrw9jqLj/Q6RVh/w3BJ6iS9CemOEnqemWBRO89Qs2T
/tCfRZxf/0eOl0ti2aOgaUV1dbUiAQQRMJv++bTTNx/tUUpFKX/anW4g6uWx
GbX9+fLCh7ohLB6DS8cR32iy0bfgFll3bPuHf/9sDF5tX/Rlia7aKaL0mzaX
GXr7AKnvUqQa0qdGgZPH1iYK5WLUo4kElG0/VpshTQ6Cq3RyxubodZ54M2MU
PwhYeygedAyAUTH8X05TfJEAHprFbiMvQSk3jWzzRl5l4vzaN02tf9einuDo
lIZtvA7DCd1fKq8WLMZnptAcF0wfGeKRB7k4m3xndUxES6aQ8cxiIkv6mvah
L1JKfni9PDA4z1NBrPoYr5rjCPmRAguMtpMK0MSaC9nATtijBWahUjyeWFdx
rfWFLcRXHgYR0h5FywByvKvhLaxKS3HbMU6z+e4O+35W8S01XfPuI6B9V5Ft
CkP1ag6mvzHwRfgS/55yFc+BdSn3DVy2Cz8pvZahpWaMyiCYzOvjTDChWhnz
sJnxk6GZre2gS8KGtcwr78RDz3VJk6iL0hxDF1wkTTDmGgcJiv2nx97YnbXn
Q4AlAYlSYo3gbcp4JRoYubH+MAM20CXYMx5nuHKEXT+5RSRsJdLAs1XEikVt
fAnIoZdayI3QAUIkU4Y6HvlDdue+ITtWa62Pyj77hrMRwQweHRxRsfvIIU8K
NyikP2xVe8YRaB2DPNqhGQfKO9EjPsU2eN7AnPMmi2GyiMtTdvT/0l2Tulxi
8LVTwLYgpFNPEQiWBMtj44/lV8uZi1+cQ8qt5u6MPh3kUv7ns4rFjrP3dnPK
myvYUyRitLG8OxOaUxCuSS4FhSSeWHPrXNJCKe25SzjkhY48l0WF/wY+3P5K
CzypnqQ+vk625EHt3PVbK7yjiTPhTjNmZEJbp+zB0GZUqjIa9C9r10RDkd+9
/tmo44N49Y81JI9McWaL6Qdt7uDYxzIRJaEKBt86k8JN/CkDcny6RoO0bhig
OrNjrT8l3Ktvd+AmjIqPzMYburmjl8nB41B5F5QgtBtvIzcnyomgkMijepAn
co1C4T/LKh010j0pnh3ndYRxLz0bCUqkuVvhoLoY95a9gcbZ41D42xQhqGrH
mkIBrZKNvJH8bodm4Ntjz7mtC/P5KHAIIFd7EXk8OLjGqgjgqXQGu2LMwHbV
63r3ZqBwJup1w1Cfo5Qyh9GEEK/NF5fwOXaLuv8SYaYPbeCnlKXo7SVF2VKn
dSG1puajuzkxszYAtlTcIP/ZAQ9xFz6WlcgZhQopI9mm9arAdZU94V8uRW9w
EzntEoBbURxlTKrouHPcqVZ/Imy+dVsz+pEm0jVjxXBj3ea5pgOTCwzli9ok
QryNLPc2lxOMEwXGgR7DDPzTd/1QB6Zl+MQRSrDGHEQ8/LkSDzcEbZEW8PVc
Y3NBUYN7ug8giKHyGWWGLgs2UubU1zmM46WwtAUOb/bdjVkQUBbQmEtsK8N2
aJDWfPKvFs2jjyau31bNOdsyxyQRsj4SNtjnnyxddLSGoRLYEVxrYsTdN7Sf
usVC5JQmEeIzzqF3MGHSFAksAaYpdKpaM1C/uKWnmyrTBYLRCCGLGMdzsfhf
KWpEja4nL8Pmxx8SW+AbeNys1/BCF5tcxHRR4bbNxsifPJh2vBqtr1us3fxW
Wc4BYI6vJ940vlNeK0wa4WlvbXjMUCQ8IZUtVQxDdRydmgkD7MlrvYfwT93t
xK1Z2a8W+yTvIX9dBWe8DW2Y0797swSKbT8MWedC4tE37QYvQWonh4oW2kvw
1HhTtmqHH7F7NuqxHOL4si0y+ebmF4Ckjt1ycSNixROF6+QB4jQ3KYyYcXqG
P5sLxy5T4VSUXY91sbe6d2njKEZTUetC1stSuRnY4AoiJAEws+nbHrNnNNzn
AhA8SO0ODnVVOrxuAuZTk60lcAQ3icd9FHuoWirzHOakXttxonk37Y7vS9gL
itUAYNsXaVZxQ/BWnQTTJXIgnPxu9feLPH5jTFIctxauHP9cjnLCnY/9lZHV
sWdjWNr/1wJw5mo2OAYm+oC3EDTuQbL7VRnGiRqcqHUPmrEib/qy5t30Mf9L
lQBq1ztvEF94QcZlKmGyLbcRYRIOWs9KTvRyZ5hm/De9ocRsC3TxyrmXuU0m
P99CjeFDj4M4iw331w/0uGHp+BWy+eaRSnFze8AHHjQJmoo1DWjg45fXpcz2
jclEOJIGnWEt3PZpjwRD43fxIqqsRS3l5Xt/3vhOCeEAf9e9EOyWplIlQ+vy
JbmIg4tUJFGcHlrZ7zRGUWnNY4wrjmqqaOqwFtYe/+7qahmEZ9AnGel6SZ0V
Xa7MkEkew/XkQtxxt7DOcDMkrfq4ssnkjeXi9nVdkmJ2Zvfa6pKbeDOfD+F1
AhH8S8dqaCTiSfsdJH0veONlBAZ8yMosIPTioqJtEil4qg+FUJlKXulgOsgJ
r0oM2Ssohk0JNGesyQU8ALGtqD+2N1MFmwNivMNkm80ky1gNNhRESaRna5r8
xHkK43Q1FtEf4ON8TtjzzB4g6j0I478d3Nfo0b8hkqu/p8puTiZaCSM9s7A8
ijSQ1h1n/jv3auKtBgjion56QaUH+1CYVGEDC6KJDtLTVRZyONmxmjYhb28T
E4RqR6MKWxZYS5xFeh5bzCCxjYKf+zhDs7yHL6dP822robEQrrepK18yEEgO
eNLZYytrmKg9Q7fi+D/mSvtgzkrzGRqi3YSnzHwfiM7k7jnSf2TjKQD9eL/x
8nCvyoYvtleWa9FI7NRxmCdOU/BBqio107+i5IAZBfvp65g/r64IRJAT6oUO
BwW4JYJeTfunTzVyfYJ4s8QEQ83SxMeCwfudNElevhnX+1SRAkP5JTrzsMxC
0mPtysAz17ftdAQ5SmlyJBsfL8KpoVIJOHy121mHcR3u3dI1wWS/JzORXyJM
NKzMFRuKO0hgSj8KKbYqFVWYx2VrzzQqBfMno4H45YZ0KfYTJaoHsIuV5iYm
b2lGo0bmb6EzMgMd/4sZOQRhD32l9NK0yrx8fAsi1j80MQVbLYoXgjCUgFN/
2sTfiLBbTJ/5rxAuENOjRjQoc7nOGRRkmif7gPqv0eH1Y+4iOsAj5hMvQPBb
uonnXs5M9bARFz+T5gqnrUWLE3PWBiYUtEu4u6Ksj1vIN+OGMmojPsH4SS+j
AZBZudQbMUTGeTq7S4frEarRE/BLFhKIvZIi4q47beVLcbcH+Woqay9wlmPN
Lk3G9WCX+A4kYftocrkl48EC8hJm1t6YxA3V021iVN8AS2KjLHWRbvYJSdw2
kgjHJugD0ytldZLgU4ArOFbu6wN/h64b/qVwwzk0Aa5Xc8hsZ/q32A71i7if
Dr5B9ozWzi3iIzp77d7Ewqre2owmpOYbPfLp1lfocTlPeLTQCI9/+1JyJOR8
dNYS1X/xkUgAY0AUq+XyZdorEphH/Ia3jdrvOUcILKJ5NDs7Bio0xkDVHUDX
KX6x7e2H8KhHMHX2Q7PWUB9FZcQfDlumILD7qgNIAJQYRc2lEOhZps93aHI4
9MJFDW7uGEVMYxcgVLSoABxWjjZXLcJ+alWD8lhnV1XVTbpLQDPQETLdhqn3
QGN+w+swRJGo79NN0Jv7RqlqMVITHM4gBIkzxnun9TpG6Y/gih3n52fkoZ9P
kqHOk8m3X4k0ppm2Pz7ju9P9BEuR5Oc8iz73igGwwI5oBjhzBZC+DqqxFmVm
IwV0mA38fcmF2d/dhbVUuiVh4aWTJ62JvCcerSIXpcrqK8XTFHBaO6kMMY7C
YiLDlmd5Yy7jSQDkwtD0ifTu8myaYlmma8loG5ttnhOfQhXPTDn0UXWiHHfn
3kRS7wj0bOFGDaTndMznmipRPtOJd7Raisw12iQIuN89n7epL1gIz0cbwrnT
EFibPyC+7WnQpiJ2mHMeIecNkdPjO3nU7Qw7eD10F6tqjKkKVpSVcR2P1ijL
/aNgg5N/VQf99lNYHQXNYSYVLTdljPTBFpdkw+a9+AbQ/hvUBt781gtuKKPk
KUs4UU+gS3KWNkR1z00cGKoVbYqtxCAVog+QrKvO2NN+D07cKnkCoCU4u+b6
91GWCsaD0zKTi6drFaBgLGUYcnBJf90J02AZLDRWAlSC7ps1ujk1VV3CmluB
YyBPysInSQQZUWSmJx8qNkTJOfwHVW4cQOFflX/TYy0SF4J9/CUhGFK4LXVr
l80jObVPJ07UV1uaDrIHa6u8oVTdUps/9XMWkVDOC3JHsMcyT3+Mg3BfvqO4
hToK0KyKUliNLRFihdKFGvTr3GaA6ppnE6V5CcUiI/coV3aSnrKHCtkbOdOU
EH7EI5YZXQWcNqKscNmqjuSBDZ8TgMMl2Ci7Sr7t6LQze72SJa8BDYUklFxn
Skqn+3eeCYGS3CcSV3kt05JbUx9CChI1uTlcToc3aB7ICmd7X5ju/AUY9J/o
x2UW13kfk905Zex6E/EbLTFSgldzNYVUgz9E4ebY43EwhfWCl0r9zrlPeGrV
Htz1WEi0VdC1jU84wZUowc7ipuX4LG5CWbTapBZ16hQQBB+sL7MsSoNSUv9X
bNbeFoLbhwBKUu7TyeRqKJ6PrlJHuECq9CoY1+sGSTFT+da48uKTQ/weMEQp
zX6YYkv9XUc42fFa3USdPBq63+AUW4oM7mBT9xYfDCAZgNSiTImfWmeDuLCq
DshLvoMKGqSufuEL5bhwNch/5XG0N4hD/sOLtTjiRQ/3uENivQwSYDiHsq99
bONv+9WpH9FTKuIHe/uxhA4cXilByZ8KhBGAuAPnrhxLxySx2XSSHoVfqaH7
KE6O7bi3tRSSu2qAUw8EyNhO+3VKoLXXHQJagOtc0/AfT0Itv2YqoEQUPBuU
OuNZ+lpbjp7cI1MUvzbEkJPT7yKqgvqe6Q2XYS4YV6ZLulCxc/zq2zkIF2uY
+kYDP81cF7N34KeeBwHha0jZeCyJAaCTBBXUbdYQGWAAImr8BlIT5oMFktn8
y9+6zrc6xUTQC33qFCAHO1Ot8o4kjNCLI/YydorOFTsBqgRZz/dNwyNNhil8
OuObUjQzK0RUtiqmJH442/Nor7Z3OTfaoDXaGxY0oGRWk8neR3s77rKvBGpy
tr6U6FAG7XjYDQ+wvwWXc8n0VXeFssg+iFcT1A7Cs7VtRPzRwX+zQ3yMi+oh
YWkEpv8un1tUfR0l4vDYp4HH7UxU5PVVMqMnMRrGStd0t+E4JY2YQoxKI6wl
gFni3zhewq3i9pVNeFLACinVoM24nchzIrvOdxa1VgFZY6r93nRiwDUER+UT
+gMA2JtGRN2Q+8R/vYDaM1bXXLCtUIGPDCzG1WLKFPTVksFOxwfbM9yxJ1Rp
OFeysz/1JTsndV/rQMXDcZrIK7nwV5CQ8/najIp3LEyfl8hL35PF6znq9uD9
qOB8JrKY+i4yMerTYfehWKIcFKDzakfu6rG3vUz0AjcvdP4pA4d2YzyrbFCl
p1wv0Z9WfmuYorec6gp/XxBDDOpYdcbxJxfxbXUWyHmOsbzi7Kj3xW3aufR4
yQK+aaG0a0cduDTl6lpya+AOKOm8rq7ZLEdIpsmgHRuT6L7loXQaUa7SpfkI
iLCxCcBQvgmPgHVoVeMaWPharKu6lLvmOLIZA0xRa4qVGGPw5gJP5BX9g8T8
zsbkLDJ97glIDrxx5vUjEHj7JT5Yxs/wcYgrqsgFReqJCdBXz2OFmPtmM1DB
dGiC/Jzm6Web2u9juzoSsRCyacCPAlFlxuNthsZNocKdZF+5alxAcyTyjUcz
jUmI0a9tDKf3LynRoTv5IJ1GHjvOPbaxvr1bYZOw6vUovLjoSPw2IM1bT7C7
7YYdB1Uk9ireRmEjm97lQ5w8sSnO1tIrLfs+XT52qQ6WKmu3menvkhGh5ZP9
b+yvIn3gGQYnMPWHwgvpLN0iRgr9+CiCWXjIz1a1ffwk8xiKdNo/xfZWXOJ3
r7wUqpJnQuMFyVHQ/qSRAt5b73FLfv/5ac4Nzn6RyDtVFLT0wMc2iXtquL/O
Jn3bWkNSpFFgfaEuArR7LU4051MnEClDRfvyc7DEJgR2tRmu6c5M/SIpMEPK
fwtfdIaj2jbHTLVrBMCK2DZfvhq6G8azmvg0cwpqIoNrSsbjyquHta5gjgnN
wNymh6t36tp4FKdK6bHPzgXxA4ZBnsUfHmy2I2z+B5mh+VhlLpizeJ10iRnp
7inmjVISM6Zh2/JubA9rbFDrlX3u15NGK6NIXeWjA5ivWrAF6Y5h2hZ2aLsM
ZPv+wjVTuRuH/F1RYCZg5XLleb3NX4zyZ2ErI8J0m9Jbiwq1+jPuffxxgmXr
xQMwLXYs98JEqwN/bg+CD4plSVc6pbz/NbkZ6LlCMXr8e6bmT2FR+YqDAT2e
HZj5ygKz/kVqaXRaKUvWXOKlJspp3IRWOJh1cuoSvP7Qefl7gQEKfP8/xMoV
ohr3w2hil6lO14Fav+BjuFs9IJrvAXIgmlmtMr34SjNMy5dJj1QiU3Wy7zc7
jz4Gb6YjwJiyPLisDpTZ1IDhR4Nchmy6tbGr1q7bONf5lQf2Iy7/aLam2Q7d
mmn+usiThPhFOcz+VA6wmDlG+2z/zJtci0YrQfBmGqjldAuqifLmnxNDEZs1
LGGmIbnueDYZ4hW8bLyDJJ3D7EcLZ3p8RltNNtFrf4+NTUi7qUWYjplIvD2j
7st20+4nenH1hjD+OQEC6qENFxeREEUbMM8T5hA/jzxWh9QzcvCTk7UujzvB
gIheK1UQ6wU7JIrYWKdgPtWPk+SGsCr3tlEIw4QerZkPp/j3JLVdC20W5I+8
0rItb0ERn1GdGUw3F6r4lA7BOjezu5Yyph6iMTp0skWPDltKjyLpfDvpsM6z
BQOwS0ugLFoDotxnmFqGb6w6/pY8L0AxExVEOrhWQxO29pC7pVAhBSaxYtsB
8gko9Cx2+6XDOBAPjqhuQzcCLxIT6I+5Yi2lyNZwHUDPN9dqfzfI62kK8EOJ
y8KZfYVQgvq/9RDSReHNX1HAO326pEVX/cyLmU7bLK20kZx8c/rBZJzNO1/e
PMN5vlRas93F+F7vSylhnfrC0MwdJPVzg9O6dcZPNmNJNuwzn8NjuYdjPWOm
JOPouUgoL+jlHn74JfgDi9evcf3/+hiw4gUZ0d0CrAx9/aiMpQgFvXkRUmfc
C0WX1V71Kg9cZmfWXaL5gJoh6frhVbqWIC8wzGWQ/DSZeTlb8Un1kShJjkzV
z9LpSEUW83eUTXaW2KTdLyI1LaUiXPmBaUDRyW9hL6qeWPJTAfynxFaoidoM
VGJRHSpoD9FMPEN8ORJucyMxeZEsWlkw8UpehrEEd27y0nQ0Y0uBjxu0DC5B
ezdIxpX/Qgxc+LmUbKUZ6DdEmkHY6c8Gi+GIVd+OBw3W22rKTasu3+cyggL7
9s3Yt/9SDg94nF6wO4QIRWws++4KKoRRPZzKJaFOpO994AIKS4lfDgaOK1xS
LLGx1xK+HnqCWaEE8xbLUdqUGvVp1Dvuk8+rKwuz8lpQfq3O2c3y2HoCouPR
AM6tnfRvexGCbZM4OcEj4mNAOp/ASSnAWbjJAhW3PMdfbRCXhDG1eAiu0Unb
AffFtIytQnUR0LwtM1aYXDvnSiqV4WdeHC5xhIy126Ddi3JPZQLS5XSVz+Wq
tKrZ0ehRnmk6mjtSD7emmLktbUDzVx05jDMD/xoG/s8S4A8Ms6u8x81rQxRO
tNMg7H44Vp7TGezTP+EsGqGC6Gr2R62XmWspaoF1DJ0nfVgAijsNsHW+V2KN
0KqsVaiJMofaSCTn2wKj8UeB6lSeja+gUyjdad3ctqZfZy1Z2E84s/6tfbqD
qmfro/7dgnMVpNNkkUo4CG3vZgCYo/16/kl8bCdYMC1j/qqKcpA7RmRuUD5P
OhzM1CZSkSvMLEcCzVuh0EEtRPYpvatUCBmfesHbqaZP5Qdd8jMVGAJiaOYP
W5IaI8QLNrL7+SefBWhCQYkyUVQE5fmuhkygzQDeakSW2auWWmd9N8MVxrB9
rMvq1S8z4Pskkzzw/ZKeHbNBRpMq6eLaZMRMyMdSskgtt19dMg/B73ivpCVB
tm6Whl7ybn2lgLYYy8UrBU+r65JVmGLTXIZKYFxhT8A16ZmfQ/XCPdmsvxgr
uy6DS0qimh59Hgbc4zcdUKRUkFXeUqQr7i6FSVTYp4htg3C2CRhcstfAWLgy
e10eBe3fjLCo1k4A8IFG80b5bM5MIkt6t0l5Dn6uuwY/SE/P46+B3jFs23K1
Zg7970R3q8aFDsWgRsvpSn2UGSPrCYoZnB/AuJI5q8yEFsm5mNOZkOsMT6n2
FL2zD5i5wXZ9eQsa1qTDT7B3symcUIUa185esDmMVNWgF84jBgCN7gNcu2GC
OeaiFG7qs5NlU9kNtnG/GlSYrbcYV0hutyWMdzSdAA/JX08yJuDReROYMHCE
KUQWPQz1oOdpRVXqgiWe10PJC+IrqFc7RO5P837DVQtKZSvBFhcuHFffKVkU
ZpsYMvGyZ0GaxZm4aAAFuIUrJcBz03O83D5KJLr0sXP6urJCQ7BYiYiVqfwy
uIoNbTWHmGX44USCxVUs580kz812ORTQhS7NvqYZXXGZkKalKXoYLPqs0JPH
p6Fc5axjIxbbkZH/DCUKbPeUiipR7zv3vbt+7JnUwZ35VUEN43OUr/AROux7
dyeAhToyR//X5I6800wDvDgsxGMVEBInEP3JoA1ouh182aEXOkFZOCT++HO3
Nry5F5eTWczyFF2GwSY0J1aRA83Q+CTonfrmyCz+Y3uk5IAwK0dLuws8vZXk
WIM6p06Bc3SNKfi7GUvejbPvwGCjA4hpYs5nLLyQTCgAEbpiapUD9FJfglqw
q5oNyfG7xG/uVFFSvKJpgc33EOcXepH/gMaRM491ajaxYAqubImeCvsDoRvy
w0AFSWsHQed1Katyw9clckKPNgBqVvjVHptfB1AEopHebPUE48GhJrL46aLx
sQ3Zdgnfk6LiS+k5dMmVVeEqVjMCchpJmjUtmipZn0S9ECF5APjXvWnGv/57
zPXpjyeBvlOWfe5ti9cT9v8P5H2UaqsGhGUCj8rVLmfX6hm6SBg8BfWVZXMo
VYXTWkrOdm9SDMzAc8wmviR05Cq/ppFjwut/rnqQ1LIP8wVnOupFHX0NXgRh
iHICbXmQnp7Bp3nY072WJXc0nZw319IzK89Bi+7GvSqMaSzSLfIBWz+0lTCA
FCgKqHatmFTYE6+Yf3eM/ETmIpybvQhfs+2dSuQiiUmWKPjOEg0offBejVnN
ea+17Pyo7W2tm0ydoQjtdaEOUDU5VktPyZrPYy5xrLbtieaqiAnioMZlZEEq
ovAs7T7MY302jp2/cnxBEoN84rg4qcjw8gHCT0yXMzgelw77/sdvvpCZhgoy
OwwDLK6ppgF7Z00S33uGXtRcHvfk+X/OndyYHK/mrqGhaHPD2aCjZmHWhVjW
OLLOD3yInZE7229NAuuKWZfVSerzaMtNyq77oR3AXCqUdZFszDThxH4M+Qqo
g6S8tUN9bRKJn/4sCEe+r7Ahth+dfGTrr37FZYopMGMJFeX2O8jeu6DOOwnW
dHsnFMRsieBNlYX4kUx8dsAMrmaaGDmuUromUAP+N8VPFqq64f8Uyh9eLzoF
wef3yFk77UK/7RVWM/fRdaby3Utqa+uK+8V4uypTPmNPY4+MXfh17bZqb8Wo
I9GwgiFd70+1A+KxJv73MmNlPsNprT6fsuVQY+fQZTEy8bTGqzbE1Ctd8oXt
nHHiyEPkAvmiW1rwfXo6Wo7sBvbFMoEX074vvxumx7jBFJIVctSYSQCrYgl2
ABuUqIekOB3rexJ1HO+sPnH2WegeVKeWA/pa6ZulntUd5hSKSycubA93LR4T
fz79LKqhyLxRL8TXNAYWHGYnlxIxCX0E/g/tbEFUUOsPVft7t8+WtkTsVq3s
Vxlfn8Dhf8F7hRhB6MFQ7hQ+z7/86ATLlxhbKursmYlQhatGBDSPYAG0S9EQ
wYUTpZ82P2xAm5EziPuFYngcyTizr3NtqcjwKFiKdrbGHWg+Z+aqCEWLMldA
H0KNfirEgAI6aPxCWBf0j0dX5Gjlxo1C1k6A+u8pVaA10SPNFC8u2igp8QnC
zOWvdje0xxy16YFQfOVXX7XCBfEGhCMzxeYx/U13ABsj1nISIIvm7NpVh4DI
aus5e4V3zys6Sv9BvBRbLfiqy3TqzCgw49axEqylpp7dqjuEq83nlCiUVJH1
PjX6sLVRgS4iytPS/HfIgbLxKFqD/3JE7iR7kTzF/IWu0UJpfQnGaTazwfFl
651c/dwR0hJELoDwLvwQMERPGeBwD0+grnWQfw3luWAJKtH5na4fW247DTrO
dBCRX9UtEEMzZtVVQf7m+WG0aiFvCeKHSHTuJ9qG+MM89puqNbSP+jVsR6nF
6+ctZOc+eXDf1k+OScsISvmn6+N/FdmhfDYvwzaV6fR03lrVWcZd45Hc54xt
sGYVABGHRt/LinFGYNJwnQ+lJQuoG1Ie4mnyvzPri2Vzs54cpnrEZfaVpdZT
zGoUhySkc8ZoVGre8FF+tg3Smlq+OGgAXkibkomgs5aiLaANYR+j3pPJfY2M
is32Q7KMmN2Q6Zibrgdjyx/WWB7STL2SdtnAtT1iYrPyBMx2XYkGaAsB8CJL
SWB2BAe0AUdhHa0UjKEXyLGucYHrRMIeku4dWzTY1X6xMhzgEfCtHiKDV0ek
76QYEGok9yYlbs2qag8uDkZ+aSieEVLo+40XnEIY+02/n8mZPOnHVPU4ILpr
Tb8KTPlt8JxFXjv/v7IViYzFGz9cSq7hqXLywlln62b8WoP5n1AKgM5KjAX7
9ZQCoU17sETFLehahhn9uhhoKq0o6gSsbTrYIKy4XTm+WxFv1zLaBFGQZw+Y
LwYw+MvQE9/gGK2/IEYnhy776N43YnI86QfNnvhK+5/9m3GXlldZmqco9uHH
IWHOtdU0vibW1y7z2a2X2V2HsYMAI92pjC/6Otfjg5amhZCMWlRVV10FPmNd
hQ1Q3LurfOrbF3uy5dk3wDsDhDQnNbqLcD3Xz23bUWBwbN76FJEmQCps+kTH
H/sMb/Lcsu40LDFuyjrtfqlGqCh1C58mjxdzEBWFN8RvrA9oRXmKzN+1Fp0t
KWcG2Y8gBVgZ51u/YYEADxuLv8SqKqdbp3FYjNF70BVGbdcMd5wy8YOoT+kA
sfehc9Dlzv7g/zSQhcEFWwlwCGGX2Gx9GynbgRvbsEcMwPe8Rlz7CKdnKJ4W
tXycs2QCQ4Af+wABjac7TyV2Zn87fbqARRDQqMTw5PEmjMmhvZYcUYuEgy2z
L+Ym500ZgLw62AmIjIFKax787LcMWnPGLnDn4/u90M+zYbM6ZhkRe9zuW0VI
fDF+QgubiUhGhC03e6YDR/OXst9syJ1NET4l+N/0+0eVWXjFSIxSbvB/41GU
Ym/zbVqUqyfKzfvYhpQFWFgokJRx9jstLoPKM+2u7yFkVBsoMIOIaoMr5weO
mKCCt8XC1KWA8TYf6A10WAxp6DEt3quGq3hVyvo25VaEW4Iar2uZctPCjO0t
Tap+8N2yuEEV+X3/pK7f1PHct5q5hwZ+SavpVUBbDKP4vaU+U4K2lSxXpKn1
8It+f4M2wdoLQXRY3a+YnE6QJ4wWqDYPYxpXLna+beM/+q5JI0d0K23j7H9z
M/dfNdeqocvDszeltvCg3i1tnfuVanVA1USP2efoQgLtdPvEVd6vfYi7Jip1
mfZwABat0YxzL+npNHyPXCx1gewAblWn21lkWLOCfAnQwp4Z7vSH/BTR2RI2
QrPQ9HnzdSs48+i7rLyMpTV4mlFyTQp8OuJaqSLAyWaUn6kDsAWAs41BNPQ6
Sl0nLleSJRB3ph/WYT9Aq4YETiVL6eXlYdQ+24iTGp3gsYNB7FAS1h3jytHN
v8tZhbWa0UpYgYXAKgMNgQgmIqTrmOAfO21hZGoIpGdiXcq/rKIUrKNCHryY
zP3LH5GeEA3k4PKyjowGlaVFVIz3KhNj85870yqxoM5LxFWjwgWFlqtV4y5R
KoFlccIqarHHXcYgJpWk9XkiKVPe+hs2i1PoOTmpPLn7EpbHLry0a3aNtUQg
egojINghw8G35mRNttB3AZzd0eAUh+3gGH3O1xT/hSdRKI/DqpmNEhmB5xEg
TUwq7IWMGDfAqfD49cW7dGx2qzeob6bmb7/Lr3l0uqpEWi+b9LRf6bD/RbO8
BjhjFChnc4lD5rxBCDD4T+PjfxlswEnDOMcT+4DCbFB4TbPZSSvmTfjsu3Nx
xQUYbnJgVDnz/bx67RYNZ1jffL6K2q38ZbhbrpO/JMdGr6TqbFEueK9pe5uJ
7aAtKUPoryI+0Uvsavof9I5xEXmfdZ5/tyBso2i5jqpkiiPdw9DA+QG/92Ow
Laxw/OSDN8VqXJ5exHImHR2ok1uIBGNK7TyPRBFQvCcTcmc+ATGlXJRjb5sR
EOCTrQIgx8ScMdzQHW/icJ5Ror+hteE4aO7552TXVPzcxL3Ndah4ZWLLmUKl
n7I220xCE/Rhsvp3lIhhsovum8Q2l+ZeorC4QRydoQohbZpwjWX5eiM91VJ0
GlKgzVNlrYtRyOECqpFfixw15HW+hf3vfJjaGM2T2HUlc68b6zZBP2GjszP6
42c8BP58eh1bGdjrVxW8UsIi9uNNzXh6BScEheRuR30/IeQ5u1ZcEOABYgAT
OuX/VMppakraWsaS5k4gOjlG3R+X1BNNcfKP2IKAv2Q4cvpOtlnwdSl9bLUO
xhFHeCxlzHNyhRR/pZ+ssIWvXoKS/yhyZGwMDqQfeJqUt9O2EGfNQEXSe76L
psefmwsTezV9h8oGB/xEhQu29dk97y9Jw0xui7Rdi8ogTBSGbrf1/6P4LUcO
tx4eW9v3yNQJnGGW1e/7VBMCiXwT+Z97K8F35UD8H9D2brUERzfMKQ2bj8nt
OY5A3qrNKOOFqo2mtAq3LcK64RJUwIr5d+RXKLootz4tdN89SEj3M2cJ/ufB
/0jNkg8Lee6u6XxZ3Zg6qLMGFVdJ9O3kfy24BY5Pi3A2XQRAkQ0L+13ocsXN
26xjHUIxvGQ1sG6GaWjv9+5kZopMBE5QcJ95Ep58Yd6bV+Y3il90pT6zFi3e
hm8Knd1YpZ3DXYQm0zVnoSjhKGHb2qhqTCoWhmtWTYNZ378Jg+n6ACnB2iLo
CYELAOlubhngHKsLW4/KzZRTrGzGqSpEMUwNYiTXM9RBjVcytVT3pDkCTKeF
dOTk4Kvgs1NrxHNAIObyEZ2qoJnFRDJp+RO1Tg6GzWgtBHm1AFTk9TgJCuhC
XOuAjuPER8KeMoYsdsotTVXqFe2YcxIchscQN2dISVP973BGifX1OjbhoqNp
nPr9tXYyAM0iBAMpqoWsoXsafikf9o0G8V+eAwnNSIgcj4wkyQ6kTuZr0qjl
ypfn+ToHxRQ9zGWcwck4FE1LJU4EpOMybI5QU+dLYf63ivrud6Ac3vvssfJj
ML4Ok6okiN1RjpK6JByTVYr8IbZxE3+4+T59Y6sgMo+3dJ8l3uiUYNb1O3ES
xUyK8jAuMLlF88UeliA7uF3VMpE+RzWmttDpp6VnBPHmUfWJi7KltnWfU868
bjdMH2mSjdD8hf2JVcJB6Kjr5XlnAf2gkU/WHjpwuXExDKc6UX6dabIsOQ/T
kuAA8DTMXDjp4b3Cqo2/AMi/I++tEspcRl9Frp/115q9Cu8e1unr2fEGkrSI
XqxWGDH/oHfamVdsXDjZIBmXqnwJrWA1au+396Jn9lU2ZoQvXhb87040oewn
YDm7KVFjNL6JAb+pQZStK+Pe/Cs1C4AozdxzYr+A4Cwb+87pkWt1dlnmI3r2
yjRqCtykUIxv5OaYMlTtneBAQoB+RzS/lTxdB3UKKnAle/k6uONAM6Sk9Kmj
v0JyrgjWwboXvEWQHPV8H0d3aOQ+tPP58+EqrkCEmEczEWnvs4L4GmsTBe8i
jWFC8oS0vE0j2tMHowhfcvpcPCsMZmhhrNALq5Nc0/hQkQrryyzhfe+j9o17
prDyjrvMk9H7YN3OZYhQqUvbNSMuJGVd8X9FK4RJoR8XKNQZKhWgefhXH35+
ahzmlfX8SClpuU14vdvOp7QlVo/SSI2eq0eJInlCt8nQt/TCsX4zo/OfD9HR
ImQ0jSk4VCVK3uzusUtzXc8nd5KGnKq34T2RKCODmIscZg/d+eF6ImqTfNab
RLv2s1yblwyLA78FBrMPcQrp3E2ps4WQVqWW/SS3K3X8GZDyVP+pFC5A6nc/
P9sfrk4fWP0eoFCz4REwNGjcuu4Hm36zgbmfIYsN5GQ+45l0QnHi94Gz1i2t
5wosj/SNYvjEgeJr/sijejvITRQqwWIr+tOc3YyIurls84cOhg5x/VWmU8fX
9Dk5ZwIq//8N5bVOVGo+Hz6fwyitYSTIMRn+tl8k2IA/fYHYHoBc16B9upbk
c292FKLHopmRBzxoEhPRL824gTomiAdqlY7EILbf9Z2y4Pwe1irdD9Yqrukh
QiN8LmxcFrnj/3mpk0+VxnByHtE3JgWaU1AP6lP1eZo2z4Z6qfG61pHURiHY
ZXq/20j766VHr5zD0DfRP/zXO/diPsyC5Hm8MVU3hupY1odSiuqTzl0nmKY5
Z98ejgPnX0iC71GwxF5iUGY5of3nmt9+mKheptGanAlUp78QEQ9OHLQzfgMm
BNDJhwEvi+m4C4Z+niESMYGdcsSm86LQLSoqqZPNKGSYz+W6Up/cONtT7pwD
gCCWeNzZfFZapHslCDdohmror8XEcBkZmKWuZNBGdFHCWk5+5Y0NSFFHW1Yt
95myfsrF+kYF58kpyTqluSiu+F1GV7Go+KEHXhcZCIePzn1OUpyFfiFPZYTG
xFqBRSM1Kd4dnbwN6ggJKUhfzypVV26BKiQ21QhkhuyVagenUQu2S6uUlm0b
kUEeMd7ppN1Dh1b4+SlZGV/Kp03XUePZnLtYbD+tPHcDDaihbltw36/AHZhq
lXqXPZuBzlyruFK0MhaRekVgQOi/huVqR6LTVo1FA32Yf+tL8QZYAbp6HTgY
6KklkVOdT2rfSfpNvzj9OBCnjHotJbz2UK9/4/SkQAuczUPMPIMXh9u6tNr0
dDVT09qAALgDYH/q0IKfvyvKblyVJyStLPFjRVx3g6w3ukpqETv0mQsVQ1jj
YJ2jFVjm3LK/s4i6r/UdHIKCtIhJmfyWSnXfvoiMOCIogND13NRkMjBEKquc
7YCKdBnCuGg2xHvQ1hiuSSf7jw43ezqr3y8Ra++jHcmYQWpqISNBWw89CD2L
/8vHDEfx3v7J+qbPY9AVr/qnUmY6tttFGe7Iziuj+DlB1c2oW+OWfQdt9TLf
Idzk5Y9KEFBnqMFZgAuIPFQ0VQljbcaeJKoLU0SJ6zlno5VqTLeY4HTFsNbw
66mabTz0iats7jUmcN/ymq/tDfiq4v58IW3VUE3dtkdkl2BJMn9k/aClkFD9
7AakwCKonGubS68FOdPVyzfpdmrPAf4kruJpUdAF4eLrJlZzcjS7KkRSO4Zn
jdJk7eKSwZfQxfrF2RDGEmdkb3ga9FNN8bXJ46/Ehe9BtkvePlhkpAazdlCo
u1IVyK992LCVDiAkZRMqm97E980M47g2MXnb0lm1PoNHINcsTYYv3Akabbwh
xaUhO3VHM9DiOafzWEtGudWL6yvqTsxEPWJD90VWv7gAKTTxj/JQvrXyAChO
cz2rnhoYVSJKnGzKvNIEyXokEckbetDBSSK+tXpU4CPj/uziZfWqoPAMfF4F
/ekrt1QPg91e8l8qSqYaI83YjP+anY5NtRmpA3huHmYRF6iFBqkmt0v5+ihi
uZ3B58OVBeoq4H2jgEUvgZ1PFkoT5Gi5OTOO6fZsMT+z3N9407ir+Eb0ZN1m
DsoLAkdNl1T+wRJZHJGLnnrU1Ks1v0sjeX8ks6tosCoNL6dH8tLx311VDDj+
a7Ow2EEK5w07MhJLICM+DYw72KI9zp52eFkGCYPWKB7bdnYMSMvqNw6AQMuh
iUneh7nz7jK3oMzupVKDQolDODrR1A5lRLNYwqc32xFm/HXV54i2NnFSW1Nc
HC5bmsXY3V8oOJUQ63vZzqbSACoXCdAj07epW+lJqPOyvPqc/oUNZq8xnPEi
2htJcmvvyfDdV/i7i++cL3XY0r5nvMrqrAZQXRktlqJyk+QBvp8ukk8AGTDN
FIA/1aQInuyaOd8kXB1aY0moI1cA3PpRhW7uX0dlL421RgNg+6/GiKgf1CD7
havOAlfwYJ8WDco5N2qF822DSRQAnhnRQ80TnaSfj1H7ow73fDWRatSi3QN4
67/g77aS1Iu8ua5qiRH0kZZD6MkgWYrgIBSIEWAlsYo0aR6hiG+CRo5bVzUO
8OnMNqAYZ8eEeRVwGAkWDhFVPss8UxkUv6PRDLy01Rl04I67d4bu+E7cUJ7h
9zLSK12r74IlqcYujJ3pcUzoMPD76mDPDQP6p1xXIH1Uh4T6vLIpih5euU90
wlUe0macw93y6MtaArWgUQ/YNWYNhT8MQcOXk5KEve7YKGturS++pZvA1/eb
V5pkTa6rOUTI0kYp/W1hv2iHHLlYciBBgmiXRLQJMZmQrjtCSk/9Cqmg8Slk
KrlmVdbNsubYknAqx7n87Vku9yqwPVj3m4H4XB+vWGxbnW/x8YpW/90y1PR5
gXTYVasm0mW3x1OhfUd3RgASOP6TtwmjlXGW2UPwNJIN3dS/ZqIA0+A5EsOU
picYvSukFLKS4h94mZvwa4idJgikMljYud+Q7xnqO+gDCNrPMgAdbVaN2R31
VQZIrXDoiC9LC7iu9hwlz7NvwCaqYBnACI2vyVmd9oHHqmRdTsShwJ0qX3wG
ZzCt3kvs5RTHouJM5rLYRWMaEHxKErJ3Tzkweqpm0l0AdtphJEYJ/Koas0np
WJdtudzumpDf80L6sGF6/7AkjCz0W8I04RwWLF567wVlY3zk1tx2O1HlCDUR
3j1FXfsktY+steMzNxKIAVJ1KtRvwMLwSdGE+2RSDHoYP0NvgSkFnd8NQELD
K7ZtlQD2BtRa6vj4DpIps4S42wXPywAKNQEoOUeOp/hBOsIP0MN/krnA4Swe
ZrN599xpiCk8RYBzOYkd5xqx6juMIBDRNu1gDug77gZKm2nX30HwCZhA0nWT
BOxppcROoXBcIWQ/LIeQOjAmG8NnOvnCMSF2Cr159mflFFVS+wrSwkw1AFwT
mkwWr4fN1u4z1JUO01ef2ddRN8K5y4tYKUc/T5U0N4GklsjkqSSIMHggDpvN
3d9hj88VJKlBwQosoCHaA1w75enNy67ME2LMcRxSmefidp2350KwxIx1Y4+O
Cap6XMdVKSOl9TfPZPrN5OzvuUJPVK2XHNQB1N05g73d8cuCjoU6KbkkhneO
de75vu/OZxE4tjObVZwXXGRAOZx1Xw2GjqBgT1KKrFkvw0O7Rh8ANp5DoTMO
mvi0O8bmmoxOLzYqwWxVUWzvS/9PycAcBYMs2IbPYy2A2pLhSejmZ6LpmBiE
E3O+LHExcFXu2V9bvdJx5KvnFaf5ad8BkCRQqll2ZIRYqTsrBAY0Ch6kJ2Lb
Ar5lPCt6I3Wjck7M4JvXPfnDOBchb+tFR0sq/6iu3I497IB7QqHRQnRa33eu
iIT/tv9m+5JONa42F0p80kGMWqGx8NjDsrEBSF10n9duJDmGPO3/442iokW9
ycbN3CXrStxNtftNpw9LapVuWaTeHPvPltnGNxJFTF1Jy9RTfLSoa35f7fsH
b4C68DlGwW9DI8UMv9OBf5IZ+MMtpKNrPNdyOHhe0R3CkCzHcwVIYBafYQEp
LU9pkxHmX2m92g2fjxoZPPEO7JozwkGlW0IUupOjwmXqM7OIZgZC+0FguxV/
AUkINCvUR2njV+EiBgIaSV0QTDOqRBldBimASCru1lv/mzsxA/7182JEAKkA
vhZDczztx1dUpf1T4vttyOBcXv5gCpnxkX7Gg0w7TCsKCpRa+M2pQtJk9azH
RiG0HSt7x8YYbrb0QvVmugSAZnAYyaYZGomr5daLzTzfUDrXy4CHFfbkh02L
RqrOYB0MhL9w6rPTMNDT37+CV/K7P6ZnQD7ayC+cT6JusPRN2M4pnuxCVzm4
VJK1tZffwbtfMh61KcxGRN7W3wS1i2PMEWh++HbjaceaR6J4YLkBPDOTAmcL
0VBQ80OYcTM338/OE2QDrYcORTdqjZyKpDFZGO0qWCxn96FKhYGw4aPmcRKi
eTpg1FJ7xI2OlFrnGCcSs1d2Hq4ut/vyVBZfKBjpfmVqmFhNsameNhfXN+48
tW0W4KA9JFO0lWH39ds3b4g2Ha5GCHxhG1Dsy5C7bgBq4QBX1+d1+OyzM8Aq
98mI1Ssgg8rXJwvpdFR1CD3046CTJThXo8tSkQiio1Pp3TsbEFyBMKCCBjPV
76k6/YcCSvS+jdayqlBhDtoH2p/idBmCBNWaJGY5m3GBj1SmppCRKKIu3HZ5
IT5+qEf5N9cd8lUNJg3XjUsJRT6t49ANISLUoz7LbtxjclM+ChkscnBvKXz3
TNsPOQfG8QrLBh9XiE3o3S/zGCBxteIdODP7gZ4eu/TZwHVZxz29nvriswbk
qJj97JDBUW8/f1LqS2003D39KXr0/Jg1griWkpBmye45XJ4Gi7uudjX74t03
gHNRBiLI5fcY42WSpni1RYrGSCVM/+SE8lAiAva8ElCrlv6Vth1WjIUMGgNS
cCYKYppmCRIIPqhWD8QC6fYZr7qxIq7ijLFoVp/DCZ6/IuJDv/tLiua3hfKV
bBFiNrHGEOdP3+kozlXnfqDsqEF9eO+irNl1kQcCElJUdyWCdcS63AFS/Oi/
b0aGEuJyMwvOKp2N76mCkDY3Z/cLf8uhJuDV+j2doNYZxiFEClWeGCWgSa5e
Zu7sX2J0Je+qsE1RZjj8tHEjQcfT7WcaYruWYmH/XUUxgXfCFDlMXjAPZCiT
WeNGW8iQ790t5SCfp/wLti0fmC9dovcgst1ZbzpPGIWMaVffdou9+An8gJla
qUGYkK/nL4n72F0j+NQ5tPw67nJKhVaKBxI2wJiBcGN9rleBum36kKU9ebd8
I8O7yvmV7ihGgj1phn8HJILmO6UGpuhD6AFmeoyw8EhyFlBqDKWPFIWoXP/W
WcjnPbO3FUYW758Rr0/0/DxlrRDeqAH+8ZvPl0AK7qcvSubR4pwo0kARwOTx
TeFbHSzV03RE2a9F2mq2BWTapHiSb6oAu8x4GAAsBq1/CDk4UDrBYQVGjpeS
L/qF7Fo2vBIMxpYAU0w1IGm6EGmh79Kd37OwOmyyZuPrj6Hy9Nv0XFem83Dt
M6lbmjnLXcC41rT32DYLdcbrBffjkpsKlFbI2qsH6Vp0xn4RdmSe3VI6Ze+B
fP/2rd8Jv3hBJXXVQoIiAgBH1wcbz3pSClACV3s6O9vvykgZ2WHtx2DZvWfS
LzNx6vrWxz/9RkRZlmU9y9RKW4KAkvNN5buS9PYx9N7Bta6LbxZPbsetSpte
DF4k4ZL6xcyQpNh0Txv6pi36OA2hIF/qsrXZRxeRgIxIpGqo9mshV/pPDjFa
KuHED+OJzGch+svDyKsIF1dZfyDMnQdl5pBFb2iMsQu56vIbCph6g9k6+6vg
XT3H4hLZIch14/jE0NMsJaT2DPin+MO5xbKbzkgT6ONXd3G4vWb6GnI/3X8C
2oLfz4dhgyhrffTLDiOCHzewYfIlwnqqkGRjSXT8TNJwPwdIxXGEJOEBwKie
joD6aXtMCpyiR13sgFT+/7Whxlxd6qFGauBX5KnBH7wvKrAK1+m7nlLlAKzO
jgCsa/pnGL3Wqi9ag1fMlGDkR2sKUYrYxVGx6eeLYsQzcrly7yTwiO6qECtD
2pLJizjK36yeG6wGMHo1wJevrPJpIlxkovn7oPXFiPnxZTN8FwJongkLyVwP
zki4phjYUSauyuBC5X+guay9v2PXMb6PXO31kV8D7/QmJForVCAwAv4oLUHf
HDsYkf+Y6jVir39CkNYUUONqaGCtpmuHXElAVfhIwewaWUoSewdNLBci071G
+TjwBPYRhZ66Mx1IteA5c8/ULfKFHptVG4Bd+OXpBH8AUeoISS4yN437Pk6a
FtUcBEGNVqOysNWn8k7x9CAojyMYs9nFmOfnSwrKdnYrxX0r+qryEckrvIgi
LnjOJP3zI/aawq8WzBpQslL2mx1LFVM0AYR+tdsTi6euLNtLg7iAUUcmdE4q
ZFzeXNMnz5Vd32dM4bbqenOMDx7r1irJz+Jpjo1TOtkPVWjL93j6sd6SpFLQ
6ounEiyM6lstqk5brvi16aHtFSHzYDhFf7d1JKo0e7U48QjNACrtZED60l5j
OAafzcohIqXTlXGL5ardVgWQRe0ufsVkXYmNGmdrBdfTNxyOnQHrdeao86L5
TNVnRCz5KLAT3E+aU4wh/f0pBNBXvU+BmjfozL6Cykvz3Mp24Ihbqgw+U6Xj
Mr/HS4vKaTWbBQ9jU115eolnYPTNvo0iHnoA5Ouxy41E/3qDi+tqhm00/FZ4
eaiApwBiiRusoCxdAHTnzkXqpP3/YQXFCWpcx8VD0/NVPY8NiSueKzswqTPB
0NdhFtyE4MbAvk+oYjviF2qetTiywJvHy7kaIrOYmT7nnifEGUMM0zviYMYr
3aUw+JmYr+JgqAwMf4dTLQqGnH83v4z/OLWefbWlpsiist7bgzHwWaSR+h9F
xmDaJsq1C1WHvjJ/UqlDP1jomo8Abt1tI0LL+cdybPVKNosCJoQPW5aVgoLY
gq5jdLzFpI4nwwuq534DvtfDTNZzlvM9prHBtG8LY/dPWVRbLUNka/Ybq7Lj
a9SqFS1xpqIEmeDlkmlnNuo1s7nspGJr5NgxIc4VF1FhPtRG7/zjpz+l3U9h
Bj/lPFu6ljtVZGnOCozCJW6DDMn9SaOpPRuB2/ckqyAmH6Dtdh+DUSRrZM8P
3USLOngBdXlZbFMRX/oGIqVuiuMl6mcnv+NZzf+mY8bmT8RXJYoDjJiVKxH0
XlGT0ttpbogx3ERhk8dfarLMJxDTXPrzi/cxO7M37bzK6ULQNCEAUXnul2TH
f/j810mSY065gG0v72n/AKbzSqIuMYjnCkvXynJneX6XFgN1x135SYTCHFgT
ltVeu0W2TnRFYr0MuUGB/TL16R27OA+1uxlr3tFzgjLR18R6ETyZFPu7NqP3
fWOVfeclOQtJmqkHn67MbHLhgCO+Hz+FkSm59ZTuy18/jSdFtAsSk9epeRtN
evtokDwrW3s38jt1OIGUQ7UFVxUIo+v3OVT/70LYCAJmpYSXz5s8zS91WHtP
9E9G86IfdwCECHfSGIwPNZRO35J5aSxGTxPGNfPl7K20S51wv3C+GiKQ5j5R
N4Oglo6/pZz0N1w/3q+rNSF2YCXIGNdbOKqh11/oLqDvj0JFiinTvilnDYPo
dyNsGm/K43KYunz8Vr9QDUuYGR5sZGpyd75I55LoQj+mOS4ANyutstFOHnKf
s9qOhhOHJ2aNm8XgPHnaEHwQfoFxt0ahBMGP9rys+eMwi6MHybrcgw37KwKb
+RSEwjXtBrVRlh0gIB3Eyibzh1aZ5Phu9oQvyrDIqGwe4dSiV9vgAs/aZ0R6
URP1b85DRT+Wb4sXPxCae+gN/lhHB5fbEfJNUs2biqb8k7CbdPO1NyKCqyMR
GXusTZ5yBYqTEFe85AVRLwswn9RjstotAtw4WHhTHrg1qY4CZtd7tXa/tIti
/UVep0gWfsdpzEvEFx3JzuN1aWFV83xiZWFzQb9ORlP5pjcDXz3YneRIAM5O
Gxrgq8xZN50zHsZj83fxdcuMGYSQOnIn3aKHOVkmWHS3ri04OuBopKj9ctkf
1lw9lVGeQAsqjq/wrz0vxwOb2airvb5D5pZCaL4OByrfQlvwjaAslFVPjZKJ
YzWPU/91a/Yb+PMUYAWhfTfB0pCfv+eSUHSzIHU0D1dP7cytULOZccy2jlq3
feY8Sw5O4+hCE0JQSOPiOn+TEp3kPBrcMpBAKQibFgMmO2j/oqW4BWjbVMGK
8IWKmhTLdCj2u+Q+0pNvM7dGwqIbUw4YcZ1+Vl7B9GzJk2sUzzAtk7z5184x
uBJrx1OvVMLU8fX9pv+k3Pytn4jBJrWEjAdBoM2cuXWrXViJzjZBMaGb7Gk0
RYNWkdQjARrnM44Kd/G+XupbSnjDL0h1mmSQljt+Q/V5vg8qTAsSZK9oI7p3
zDUBk453baNkxqzx5bqBrGYlNEFAHJpILcieSnwnkI2TbJuP8gxCpqXE6vwN
9O2G/eBIlB0UWNiNShVi2BkSCPVW8l2HEmGAn+qmL/x7wLVvYAyPQRoL5RKs
+qlnGs6kH6EQK2RLLHHx2Ip6JlicLY3MaLRpI25aJbacYnachviBX+0cPmkP
8x5iU4hYs9V10ebSFQNmPqrchZ2Nn37NqY5kJHJx04G/Nz6bOAt9dPOcHb3O
YTH5wJfrKzORoywpac0PQUgkYITXtL2o5WRAuZHi9A8AQZZI9PyeL/tIAjat
F3C8wXfvRbxjI42lWUNwkoz6sgTZ7QLPPQqv3pAYiZ+QCUh6wB1oLDkFLd+D
nIL06k5TeGrZaJNoSX3IqZ2LDzX9INrN5IYahsdBBDUmHa4yloZOlYRIN0hL
b+iW53UyBIWHd7O5DNKPwOn2CMTrr/9qHIAmPX87qcqF7AOVBhM4afpyyk6E
CFmwRdCXzSRRvjmb4CtArjJDG5zc4uyF0Oc4vnKZldg3cQbkmX2DLuVUtjOy
NWANtFcivJ3EdEPo2kSTGJ5Ff4k/8NL1kfW+MENnPrbBJhgi7RKb5xik+gou
CCZmJx/rJmWcnAL6iKIsHBjiUSaVjqcMgnEACX05QhOxSDl8Pk6tpuycR3KD
bs4u4M2YYWCdh9CT9oRIP+FpuW2ao2uVQh9jB0QclqbqbgkWxEyTJ28DshOP
I/9lcQui81szqivHtlXzP2WHC7FcxoTqH5MsZ6riAEUG+ivJtk+5Sm3oGhtN
XTGBkTY9rqJ6ndkHT5GHDSOnfTooGGM4QejXMmiQ9VkfX8LWI1tV24g0M+4M
mjOMnbmEJTvpjkFVz8Bz4Lr7xDdQyazg1OZtwwyMUL5dPxMaL3BezcyUI+rM
QO/lDNu5aqPb3wlXoIxrWCg8Pjba0zgfh3qhzDqVIy2aR6llONdJBlHux4He
0+Bs9rH9KMVbZ+GcnlHm7/n2GCvDduQOlRewcpsTaGUV86jenWHrT77BEq/Y
3YwgCcOiYmGoWx8EQKWbekUtLPvdYqymCTOLDCcvRyPAcjy0RJ04R5Pxn+f8
v42rT6WjHLWQTJTl3yKgIZJULspobM0xgOtW2HmdDyvvMWKZOWSQ06ZfsafK
XOFLXYfHfGnlj93xbCmEQq0JMVz1PHqMl4VRFSwvymZ2PR8cBmUHV7dzxqdj
dm/G5lXEQHFZ0qCfcDErHdr7SjjcKXawuawMTF6DFbhP7wvRsANufFM/PcXU
MkpkCxGYENXjmmUWP/YXcaqsSjKrHHwAWZC6gEf5lisrAHOhsOenn8RQ28Qg
NWoY+VUlqOdNdZOwRa5FdBv/xavFYjx/vHVQ57vmHlWO4iWfuNLGERfVT6vg
dX42RicTg4wSIPAiaKC9k6BIECII3L4xyKV+D3Np5mvuVsEnhFkTNc6ULXJh
T1KWfrEjvWEdHPhTppjkUd9wsWNxouvc8yNdZOcShNixUYWNqn/6RTIMT3o8
+eyjPyMsAVRnuLYHMjsbCKCWxZ+a+ZWzZohav3ckzi2z97InPIlh7twLxuLd
gxE4snmpA10+yd9PoHw0QcmwSarSg1l6PjQWbXAmwIt21i0zVgMv5HXKnwhX
YhSf6rJIvEb5V8IdKZohizohIHmCBm4hCdzJbOepVEHSveFvGKHtQ1V07WpF
j7kjfES6AWlnn0ARBYC9r2wTnX2W5tga/8PSryvj5MPv8E3ZeZOfx2mDznWp
2PYSw+7LkbZqHdIToFZp6UYa0tnQtax9LDJH27WYMIW6JzJ8Y94iQ/bkiLJs
M94tBqh7Bmwxj8ZS9BD0CZEFT9+OJ6IRroi+6K7110r609aR9YJ0ysyeKZlH
Y/V4X52203iZOudWhzmwYbDX5pS19zxEvXS4MvCs75QCm9hSb2E4CeJH9g04
6lp+MeMB4X16U5xcm8BgZJmH7pzgkzIi52Z/Osy5d/oi2EBuNAul4pD4Mu+r
L04Ir2QAy01Ko+z4WSWBGRqGBfaw5JTSTw/eGfplH2jpjPPNkBeWK2/G1MQz
WHMCLHFciA3RSjIs/yK8N9xvXN87y0N0UPlcRQI8pJRvePK88sVkwL3lMMJO
mmazB0h49lAota0BsvRwr95UBgMrasfXoVXumtGC5jkMTk5z0S3pXLKx8djA
eLki3F5Z9vjdxvJ1BIbP8aBXyPVHbJX5vwOnl0RjB5RPqBkrpM/g2lWN9ZYH
XsyHBExtNAEK+T+ix1dioqEje2l6/+EOVverMemshM9sYXqnRCM4E18TmGuy
QDoMuxkz3FeBwuXRhPqt2wj6pIsZNqYWH38jjcyspGBVjO3f+m4GfaMINlkU
9W7lmWlU614prX+0fSIDs5D7FKL2eskOdzsFLnjPt8W0Kfab5HYHbNmSDMKP
Isy6jxcTgYopDx/wCdLko8WqIQWo8giasJbgR9GCV7GFmvMC9NPYwmJllLT+
hpE8nR0gzd5ZoesgItK+9Il8qL180jlgUVYWWtWBDXevke1ODAwBOs+Mr9RE
jsxAFqjC+3XzdsD7LBnyZZ3SAX/sKjPPKfe6rY/d6cg3cv/2Dh/H09YI2uuZ
zfurDqdJ0z2c9vlWimEKKp36MDyA4jYGqa7kjLXnIno4c4uMn0x/YwZ6hREf
ezERmvX71LcZ8j5w/HVT/7pTbFlY1NUotdPlshxmb/hYbs39YLBF0LdrLRrR
/DRjVrGUi3pGQpca4wqVTznv3Tu2R1QWft1w/4nSh4rqF+dDbNn/jv6qaLOA
1D43K698ndw4S8Y2/tkCPdow9Vj4gDDM0meb6xPUO79vdAbe2MV/+ioXVXWL
OTUgtHpjRi8dpx0JOgFvbMpvzlmdfT3kIDwhVSJFSh4jJViyOqdsBxENZjtM
8Ge4jDs+Lvr60xHhEYm5SDSDr8I8PTvlGnBCwjsKJABydilNMV3ckqpJwXaT
x+OgGlsg6UgwhUoVuPL9z+amMglNFTX81mxzStzgMSn+7t6Qwoe2pNu2EMNU
cMxvyD8KykuJhfxJV/fw4/VQVz05760WYMkpiF0qNXVpHfna7Cg7GuB+lO4p
OVOmeAiG1Y/bbhADCHwZCjmaNp/hIHfIqbDBmVST+2fPQLarJyIYeLNCVEOa
IA2FSFU8/MWxbT9Pj4GuseZ7lD6djl7nim7mgbCxv/NrTXCls5ygcffrJFzp
GQjLwgRjJ+tK+1lLy3tTWm3MeV/G104b14cBxcBGM4F/PEryY5EJrFEOqZX2
vfEANyiYAF6f1YFv0oIhr/830l7Pg1WASoR7nNMurEi96otahwhFVSz1u0td
nbmORjm2EfbDMa/O6wACULgHODNJFaQUjtVesj0hH1A9PmiT2QkYvh+k36cU
t2LqUPv5E7E4NxBHTkC8REdewC74AnkV48ZIlN7p+UHnMPEwLp4VwTtpii5k
fTdnW1VW1Sqw6UTiMCNkGNCxS32G3HBlD2Yu/oS89Jl/7qNUQ1pL3JsYP303
2nuD2oTEJQxsM9ecgJvG/6xURTJHLuHyWx9WBI5xRSjlFPDpHF3PyTh31oUc
aFZixfM/ssZmaVN0wEdD46fpnaxMIqGKlSj1cR8BZ50co9IDr0d5bbcrM2Gg
YX5zFQiaBO8MvKT6fVVSFnlED3rOxSr+U1aijzYV+IAn1C/biUt1KcBfcDI7
1pHGM/9UBtue6yWyUp152cqggoYMmI92c/ibtgrWpZGyTbcByu/nVcyW1ebt
sVMBvxp0GncKmYcv8zFoYODtA+zLBGLeAT1Ag3rqM0eNeYrzi+Krw1wIPj8K
ZonEQimj+hPsz9/8dy4xVl7LNOzv2lfn6VznhDTJ/xJKXf3N2w+AmRAvTmM/
3HDikYQ+drzRsY8frw3J9m4HojoDaDkPVDJy8ODWOVeSxzlxEG+0TpoQtofb
Cz3PlpfGohA++i97PEZYFC40ECmtSlHohetWsLzjV2FCO7R7gJi4tgzrVzBU
zJe5C5NknsFiLIsQe0fMpVHLEg4BBDb2GB97khVNcKQ/J87L2y3KCmO68DEE
ISYziSIcOnNvzkNwBFj7YqIEHuDzHHdzcoDrR97EbA5xu8jdFeAU0PCE4gm3
VCkpABFCck+XlFZzr/2tKdlcGfXIogX8E4NCZjnvJJU2cgfrCT7mwUY5qwc6
o7hYpea7rbZsij6wXAiN7llBvcPAQCm/9KrFIZwJmCdxmUN0IDChZhALr3oy
KRZL3JXautYt9zm73SneWjUdcdtnmbM0qLAXJAHfc7vNLMVv93SQjn4kPc7t
5rCQIWIGpFuSrnZY28LHL2KFP/qZKQhUo+z0c99oIjWdxh5e/zyKyXc/Jq8c
GOGZ7jPyU1NEzvjxVPc040wvNn0k1+pUydW0YOoq/TJfIBdYmqM+CqF0cNfa
5SAIQ7wofpnCp5Ap2rdA1uwAHRxIImg94PJjRWzv3x697BSDU0AQ86C/xjW8
q5hLWxF4ZR5LSvWgHP0t9oyAAPzADxQeC9TQib6mryvA2NO/gXgsJH0qSx6t
G3rTWRT85RJrmajFJl7t2Pm35/PYbligczeiMv8S3GDB5KrJqLazkaAPUDIA
8JCD/Y0xzJGr2sBC5PThIZFYXRohyC9pMwhcU07NLW9kt7ruTN6Qh3R2a36I
6UXJGSKurM97/j9WLAnGgYD+SgJx26DcdGAVWNSFL/xDXZr45Uc107v3VAID
8C5DYFIXUN7v7yDA1cM7ZZKc0TuCibgOdCRhKCn3eozrhYGccQBqDMk6A013
Kx2SPDgJxaZVVnW4xV9N9EL9I9gf5W+51hnPdkBFEZIhWib6pu86RH6sBRr5
YZTrQSrq3fnV4kpd/VhFXfBhuhX0DOVmRx970EHzxxqdtpd6QJacJHeQ4lrn
9cnKzSVjdIwyrbAlSrE3zS8WjzEZpe2cSS/C8qK6YsqJcLIBcZh+1d9oEdpT
VFLGrsZ5sQ0dtFFAGhrIgnHCReUNaIBSeOY2qmx6S/vdZy89rQtfTWGLPnFS
2bLUyuR7wRYqeilafifYJQ8OpQa06vEWcfmyK2AZIdZcFjk2jJ66fbfEqozl
ou/ZfY0aUGC5BC13mgtAtPp16OtKfwKB3Qkqnf2DavVw5e+qmil1AQka4IQL
FeGskuVT0onmAaCY+CudtvMREMYhmNsl6/wHn1EDjVSCPg7D6QPMriS3wdyN
1h3pIJxYnon4/XK/jN9jxywU9tL4ZSn84WJsUf5BpUetJsgyOJdJQnj7Ya/7
XmiDtZ8+CMbJxWfX8egCfThrE9DyPVUyJBxJJHVLz7a8hShO5port8vZXxhI
h39r52evxPzR5HJ4qauCkpFWG5NmrGLZdWLUrlohaYFGUIalncqQuMFd7izy
unsRdO0zT5T0iCKew687NEw/ya0xpSHqD0LlJ+WAnAGDaH2MPktjmGdLlftI
rCcoQeQ8ju5janD0qCxSrR5Nl0kI/uyJ5eXw3+MxLsMebSPns3/DbBi3/+Oi
X9lycbrNruTMPR3jjx/YPeQhkaZaTehsUccIFC7ZPPjhC02HKWpxAv6ZLjUe
HjedXfyrzvLW8floklG7SUMG5i1HPjIxPzr/N9dV4PNQonlWbsLusLtxoMwb
tFVVVZUxpZqXHCSNdIm3fuiBRw9XokXfaenFx8MwJ7enian6rPrwCyr1DhsJ
gg+MK4drSnS0qtCJJfvqQMJUnc4jEvjmHGtMpz4G84q0lhVJvYvgqRuj8TBw
GewXk0rlEv4fiO5GDpxmqO5W5+w+y1CLrb8XlrxsAtlP07iE4UDLdsugCjTp
2GjVwcJ/9fjx7j0TTJvGuXOmtfDReXSZgwJo0DsFMZnfhuzKKbRwcXJV4iUa
zpwIJb7J65oFd8eGPZE5gdCMHKriUFLNBGrk21A1CI7CivwiL29oexQHhXWj
J2Q4yBv88Hg7mlxlSv7wJ5Puf/tPsjOsT/XgK3dJJjQVg9WeqljU6ouEFkGY
EIxLlDphgG0p1ivBREd9gq95ZLd7bDVnIro98IXagSmg9mhpPk11fLQV5jDr
6tjj8mDVemA4kxePu/J4AikFZSSCmub9zORBygXkACLv1dvyTRv5JqK2ejq3
UslBc2ToMy7avmcBgfY+CIBOf+CuJUbaat4u1+ysPFa3qqxWf7j7eTKCCJhs
Fg4G6tkjt62C6mzpBFV6zB4KHPwWiMmOmNOgXitRXLYvMSCyMZlSsTJZPwk2
OmORLDZuVF5rdLoUxgvs52GSPuy6gbQbgsdrSACOqO8vqLQdPxcAk88aajq7
J9IT4DQS3A/4zAbeJYYB0oPfI+V6hTIlC5Tl/KsMoqw4Sbixw3yJktO1j4CO
9+RYuGSnuC1Tze4Pe77aoqaQizrTLDMsMDErSA7fiO+h8O8bCwEcWYvLPQIc
71ERAX/XkXVeHLDOp2zzQ9dm5uRt+IhAiAkphWoi1UeOfBAy/nEr4WxgleZk
RyLhx+mAB3294ZarnPiwBzqhXmsE7q3vPjfZVfTcLsxCjTDAGU5GeWC4Ccn4
V+cIUaeG1jFWIQDQMQxvLQ35KQsMgxGPZTsnZOrNE4kpTBIFTzPhZ08XhS15
KGZaF2GKh5yTsrfT0pMXh9IZOEQawdPC45YCRLPwDISodn7y/LExlbyuOSbL
26UoBTx48wOzqvsJeIE8OGaEa8d8PN26W2t/w5uWIDVB4gI/OXc8ud1uWjGZ
jfHV/NdM6LHDcDAWBuWI5vizOP5aib2DvxM09oG2+l2fuEzX81Q390IJqAQE
SsAr+qUh+R98ankTaMWcd5i0/V62UrdRdg/SDewpEhTjxk2xurrbH1Ela6Ew
KVYQ/xjgljuXkJDk2nb/ngqA0jgr94QCZaY2GIvHpCi2LoGIw8KdSsBYp2+s
JZ/cBMqQghLNwyHHw/5mEPNmYQmLl2RHZ5e3ArC9Vg/beE3WtRpgWfVVMxbX
Z7MmceEQVXt9ovlb+sTIkQ80ArEU7uMYn/0skfVptvyfc1UcPUqxzbBN/Grm
Bv4hhJJzJH7Mu1n8J/vgewKiaImp9WP2zt0qIegSGLeXQUPFH575MHrgKGJG
tt6Wz3rjIVwRK0tsfVkCxh22uHRYUMjUyQ1RHbcbQjdjxKUbyD+ZTrnsvVlc
ylD4iaaFdu0bWSm44VEzlkMxhrLxqAgcyzo7LS6IMwPSUbeW+tdGkKnpXsMs
sXkS+IFhqUnMqmjoOMiqzk4FgCvgq7+BmF4zHmrfktavPSSQ/PEr8vi4hqZO
fpTCM+AiFW0m32+MjlFMdeSx9VFZNf8mZcRL8gC2IPBD4sCO0Mgqr6P5oksV
iByKqzSRgsjmsDS6asyuC/geIoH/6oEB5c1qAIyMFeDNn8pXUtRY5CnXH36N
L8iOIZj+jCHqxxQYgCJHkKdN/j7xQiJIWny+8GaA7BjO18mSQ+BEIjdkflx6
MIC0KCrbuSql2gT0CC3g8b1wRFFaqbaTQB77PpRR7YJHTZnTNN6NVlzHjkfw
Uqkne6fAyR3q890ksTmbvZonj0rXN6jWkcMwyKvtmFqlIlu+XNSufEMBhOp1
vqyy9nXPmHAbNR0Nk5qurBW4L/hlSjkZfOeG+gXjLyyRcdvTEvIuGrnn2EsB
KH5eNsYObzVYqMZ5NqLO3FB7iKElDXJF/EfF7Kr9J//9832uXkQTyeyvScqZ
C11RddAOf23W/oHiO4HQHz5FLWvWorClj+23rSuqAIXEx6E1fg4CVFMAKMOB
JT6UgREM8hZ4nKKv7wDHHAmlgo50kL8sksmUpLBxOaswr5fwOPKdAGlJuSS1
hGXBVgkrW4dftCGZfQvlU0MVPqrbQ+KtG8dN6STTC52Qw8eOhuiylWxl0hTj
ySWYiHu/ktMiPPGodkXSM1bQ5e6lxr1rUA5/vhTWbFgT161Pw5rs5D6hFJu+
q5v5jvjX01PJ5++0f452/IXASUTxdBJb51G3SwcK/0V4nvZ+DLsRumbQYL8M
UfG2msxjyOoTFVMLtFCzFl0t54NdYTzENtdVa4fKCMzi24uXq3JFmzATo//S
DpcyxCzJLaMsMw5tIeDn72IV1AMNnfYgBLgjchE4xVn9B1mO9qilB+GMWR3F
uB9fGnJadQSUJwnkEikGT1gwzkGaMVx9crJHcnlJZCuiYLhxbDbBTAGhF7ED
4Cfy0g34q2txhcIDDetoq8LwsM14DnNQG3wVS9wI/MDHJxml8N7cI9pOzCR/
31SBvF0HmNdRY5lPCAPExHNa2BIcOLEh6P7bP3PvpdIBvXDPghokvl7ZlHJy
Z6EzySuhBdCkHs5vL9V9h2eAEFi+VXX2aLsXhN/A3JR4KVJeKcIOuf6atVfB
BnsW6kEj7OMnv6MI0OS3g5+gj6EtMNpt+TJ0VwkYx0xyjAqK/XJL14t8mGmV
1bc+wUfG4GW3xvhv9NTuQPDmREN2Uy7F6GLEs9gzEa4vGO5GyrTX+Xn2QmH4
q5g7BTGPHBj410kHNDlirY49l2oj6c5NQUQtkmSDela2Lmy8yDC8881SZ7ET
v/J38XY16Zr3u55afdGVECyJpsZaGd6JhpTU0YtMQHgZNtES60D3j5TzElrc
j0pbHkAYM4bzREnDORL8evRwGaIZaEQFnYAvAZSuCvPPo2EDULsYggb32sHD
qxxV7DRxkuBUaHdEjjOyV1m2AI5WLABf8LGdt6IARBI0O1B10UqlIcaBInPm
1XUdbIW3H47CJ19bUivZU2vBficfwyOcB1QLApuTy4ucdvjAu3UjMhw8sIW1
Qmr1fu/I6YOxvaZGa1Ugm15rlRZQot/qbqMTzGxIEo3i/XnXgQd88THDl462
0WQVSRVvk23h0BKE21nLoEUYogov1cbM1Sfja/504D2w4AxEcVYVufVKeNvd
U+MbhBrkG0lVxsNCj1CDfghSm1mQfI3kvwZ9G9YeREQ1C4E1LIRqpj9e2SVF
Jj3QVDwmbfn4y/bGAgsV1TY+FIzUdth5pxnWj0YdPmcOMCg8dc93aARhB2TF
+F8tfCiyN1Lq90Yt+QW/0GvfB92UQ8Gxd4bC7SoeeGGW6vhonDcCjvRs7xHR
ZChWDeSbJccqbm7wQmhe/SrsN30GjGsbvG5su+swz87G3A/j+usSYHqKl8dI
VN8RkWy6VhIgiUtcbqqpU42t2Y++Rn8ruN/gxeawqaGTRtcz+WU8daWMJYLe
22POsrsBMxHAn/gAxrff074zmhPTGbtu5D2gx+4StEysSF/Vum9o9V2dOSo9
wJDT6iipOwegF7GfJqBU901JXN2/CKYDzCDgqgOo7SUKF3QMt4kUOWc2hUet
LS8PsrLdI/DyLvg3wl1/NWMQ6thaN1v0faoJi8BEqN+BtcSasR1fH946DVh4
Cc5cL1OAJq6SAeVVdNMTlU4oT3Xpzto3D/4o9ZmgsTbsHAQIjZRXefDhY4bG
sNg4LKoYMhF5jOL8dGTAbica+SgZSuwG2wEkJ18bxmDu8LNuRpV1ebvW1jaY
n/bwoNvSep8Xj1V5rBXNy+VA0eGCJdXAh9H76VHcRVzEYQM5gzlzk6vTLYmd
PDNbDJ8otWDfkOBXYI6TmZQtxgAOM+T6IzY36/RjT0jSorDUvDF7Yx78/7Gy
swD9Qbij95IzUdUq0EpLTc4alM9IoXFODFpaD9eGQWZVrWINJ4pbb4bNUU1/
jIu7/DJyqeb/f2PMUxVn3TwS55kieE9Zcrbod9RaHk/rzsiopCxcJHLbhQKR
RmMCWnL05FbCyc8nm8FgaoUGbdv3r0RezcBcWVvK1OFeKeTsMEveYFf1t0l9
B8PNmdxI9qKqBtU5ae+7hKSfSAKdtgJFNzCyf4/N3OoXDQme+siSZGSyFZMP
XOU6b8teh7eTEodvfGIDwd+alRmWMvUuwnQOBvadUu2NXRibx22J9Mi4k3yc
XTKQZNo04ABGpCwgwTgU2/RHx4xitqpjTxWthWd6YK5HlAJg/XIg8oYTw1xq
TxPYpvriZDP6PEChhxBA6UfPEQqfU+qW17WNNWbhfu5N/90+DgSy45CLbtww
Dg9dpev5XM/2dIHpuVRsmkrFWUk59tSbi1AJHM3/SPeeKV1gDXcanS8ZSfrQ
V+p2vmMIVaXFpNujQsqdKExDxC0GVPNWHhOIw06I3lIZfU36/fZH11WY84gc
OPhu5K0n5mUjLk7i/G7XU2mUmyLmUfB1Lgb3IJV9EX3Zqd349y3MoMucojSJ
boUZa7a/azMa2JAGhOVWfQ4wKJEw2GF29GgGTXoB+OM+xvv2PrA4x1lyV1ZF
u4XzL4aPWEGmctBnc1/zI0OPqZINPH6n+uEk7Dfx4dh5RzpopGMALPUSmOvb
J7cWbVmQTeOceVMhh/O7STrAVh1VuPpdnYFqnOUoitGMXjdf/K+v/XVeDsM0
J8Y8F3iZhEp1T8e4i4sJ5oyEcJB2s+CrSDCX9lZ+t4dTLDiyhGF02RaKcNF2
cjwArJegY4aj12QS8e4C/DIab3HhWPoVqPzX1Nt0mwwHV++qwkHUB+g9JrgM
VcPbMfsjthFq0pnQD372OqCXgbhg3t3A1MDIP5Q3NBwJS212VKMHnNxbb2jf
YIHs8yjnVk6pTtEGZm5p+Bv7cG4jZrsxYPIvLBgDU6J9Ft6QBGl3ZaAeaPL0
SBy9GVDK8Y+rhVxrH+VJC9KpQBS83LCjnJrcDuQGykEfZZ1A3KI5K1ukXpeY
ahooiQ0TUBTfK9cPkUBQNM7Mxo92z+ZX1qAiX55gmyrXIHM1+bK8o5ldLSwA
vYwtpuNUFv3yDoAMp0SQOjmbhNbeFUG8eQcTYEjRMOdhfgD5lJT9KmNbUc/d
00LDqdYaCbuxNqaKTSjY1xTCffJTKr/hJ6UNOXSyIA8D3nRp13PoeugwODSg
Xx5+5OTEIQzBvqdWicq0O8q2PmVv1Ue+49jnZ1qzmCp6gakDrVOF9JwUPkKY
Q5SoLyyTQWRIdGszgQWvGEOu8/sNZPbFbmp084fbQVj6B0W/u0o68tBOmWm2
+GM3FrnoFyywUKlkBgIq2Inpagl9rVuIZSLcDqFiAqAEdRt+WqngbRQhCXah
5BWhi+hbLVI9PgQdZNZoskkZpSftsq0ztfJNnyDl0ZzIZOldH8CfFb3E6IGH
mK1EeMvTZpGcrMruRx9o0MRdMgGqEhIe+DHGFj2xT6tQAB5kHy21F9ilvfyg
/CYylYwOlN1uQmG53soQKk7TfUMaM3D13VcRyJ0Kvk5T/veICnqpEgC1EKSx
b7/9ctmghlC/4aedoboTaUM/YUG8+rOoXieMTNBndRf5G8AZI6vlSXgYi/PZ
A73zW9RkZkY1yWwG4rDzfOiDUZC41MbaOeANW/yYmCFyLS8rLx3exh06MgMq
UXPgqq/PF+8fbeHLbjQVloH9koKNGFvYH4/bfgOxear36FmEEVUjqqYgSLo0
4/Up7DlipnWqkbH+y+x4oKwaqIn6KTy3449cHR5rs5GGajVlRF13KZCqqnXp
bTg5iPU52qIAEZ99wLnSm912GYTNHAhAwZEdwabT9ACMQKx2WhvD1Nmsjmci
rNmaWTIJBxGZ02XlsXwGawxRgSRjO0umhgpGmszmcMcAfol77iERKeiEuWuK
TumuEPV4+HY+Vj1VOsienQIWXbkrVD+QqbXzDjwb9SCszVg7YxIBUUmzYTEq
DRy9xnkL5XgQKvcrzlCvOTTN7EbxZSC3wmNwW5zJfDVOhgFDq8GNv55/9aV4
1j1VuLRDgktVXqB8RFHA2eoRZL76lWRR/IMEV633IIMpnMNEH3Fqfmnaj+DU
hEoEs0KesYlYcrX15Q7nEzi3jvYUUSJsIE7q4IJiH6ChitlSbttNemZ9jo/7
kVnO+mTYdtQJbNhSplTeVlyUyMi5und30RbYw4GANKo7rJU9NqS+V4cuQ4po
OTpnAWlfMkTr8fSJ49IWkw2aAiU8iPbcHCdkJFqHG0enGnVGuFdjC9/wfVFm
ii1gmIYMCf3KtNWzo6PqDTMYFFYpYy7QKAjhBUB+2La5Y4K/vC6m+JP2s3Qz
xUxmuf0XqUq3KFrE3lZ27GV8hDW1qFKsrhJ8ylc5mSSKpYXJLpYODXkiv3Z+
gUKhB7kL8IQ6DzHKrLMhqS/xo4oevWki7TVuxtXH91mbGIdPxKvNqfcVdxJr
3QjzbuE1TjxqyEM5FtevNSmNvkl+WRO2l0LbVQvxhkKY03BSyrpXyImw7Vxg
BQmCZDAnYTb/F3znaPdXqP1ZVqTNtibj+2kbZyVQWVC42XsvS6KjU2zARnDl
n86C7/hOX4mdyaBTriHJuq70hZMrkAMijDB9ORDecJ8gPmj+NVigEBugnNc6
8yuX36sbv3Vkos7EgsIxYAzf0Oa5AW/Uf/yrZhUnTIdbYUlvADT0iK/Fc4Rx
tH3HTY4dUb4NFTf+f4Ww1PLA3y0vwcldkbRCiY5OIqVG3rGLJwLiPiVbTvZL
8B+CWe6zxIc+7gAb4odGQIXMUIhZJ5EWRmNw+5E/i1+uZuEeO/ofXEZqbVGo
oXvzFGPZjZsBpkj5PituiC92q4o1Je9Au6eYGeyJyYt8f4gFVNt9aOMmV3E8
GHX3XGvvH9wpJCY74QD3IUqtM9MjofBINt1tEG3tfZsUBCQ1m2TQYq+O4Oxa
eDi0KVmcUK3SXMhw+I+hVDyO6EHcj27s0CK56M93CIuqvwLDxcRBbJxOlcht
Lm71i09K9Unky5AKtjM618556SNf8xIqylUGtFuc8qUfBMk5cnC4p59uLVMH
Nhl+tTPazDkK5rCWWhc8GckZY6EsUchG7DQmU56k3gQRqm16sKv6WJ+U3sy/
J7b0P+nweXZ5hxhdVWNMkbU3uL97B7rXWp03qa62urklZ4T3fsHcetmmBy2/
eIrlw9YgsyKOcBpPtI+M0J10SmX+P+jxo+1jHbsay7Y7Hm2OgYxn7r7bfeqs
/S1dLa6VM35W88cFbPzvZZMRO24YWW3txCfqFR2kFihQBGyEzuaI1dQ6bJeK
PbA1LE9iOXL6vPI3GbRIiMEDk5Ubmc8X0Uw/xkZq0v6KpNlz07Bg7hwDUzgS
5vUnt9sQDmJ9qe4t7J2aOtbG/EKu8oTKvD/jo8YT3Jfc+u7GzAOw0nP70bRw
znPhzAoJqTcRDbkg3JQ4qSUIhZZa6U3HnbifoVNZBRQh8vywwSUBPHxYMCnF
c9bM/38Fh/MES7cmx5BNzXn1J+C1WrHTUX2eZ5hXG+U92BSZkwR/59cU+4kZ
4afzBTzvtSn9Xz3qCDY+XV59I5f90GqpuZk6VrszZZ34TGEftikUeScwRTHr
ZFQIJmnvgZasze0Tx4UC9MOYU4KTgY/jDywTQIymW1qigSIx4bD/tsEk88b1
j3/VUpijcbnnZIyG9I1z7Pu6V7hMEAcibMK2aens3FEyUM1Z9FGgBkjwWbiR
lWVDRy5pNEv03f3FOrDnXGAakv9eDSEsdm3i7FkHJooPiGSyqvmc91AJINdA
71ycK5OGeWpOXaSP/CD4i6u+ExTruiDrzEKmoemHwfjy5HhtViHUkQtf2YCt
OM8DwzBkNuMnc1K5czQLyS9IfQnPX21Z6V1wcUqoGfB2WF9jSHv9Rbn/mP/R
pKJyFdVqCHDpvu2w9qtTcJR3flDxFb0DN8GmmaUYvdEVewcrFrIBPHQi7ljG
ajXJnaX1wlVCC4d19qPGpoViH2yzloQhe7IEYtVzg84qV1J0JGmPLcOcEPrx
JnrA1ajr+I9kPis7r+74kGbsVFtsc2MIb/SREJiaUmd5aadOINo0XAHqnRC7
Xw6+lkh04n2FNEF5MeCE3BBX4umo/TeWLF95JheQlU399BpOFAV6rM1IyKPi
0r2EcpU+G56x6Zx7gGAgpgBymdjtNDI20n3nVu+b9JMGDSWQ4NN8QuGAcY81
fXNah1WvliZOQ4kDChNKlvURyjSy1ev7Y3w4+s3h0+EvIPxYeyxKsnClPnK5
tyFeOrCtBx9pWIJD0xt7knQVTA9ETETK4OKR11yL94cSng2Ibo5jxeCjjr9T
YHGO3B43Gjaq1SktbxGUO07zvM/oFFV4Jy+IVq8YR6eOsrZD88jGBUGiQQlR
At3v4IK5AUABzuqSYqsCJHuJYX4fCXTBn/l8AmNjQOSrzXVeJJ0S8+7ZEqVt
VjAgaJO1nR13jZt6bNxvZO2XfJCZP3C3u6RI5JQu24o6l0tk/RF5qGIwHJMj
sUHwye1yMvjgAK3LGW7TVeXKESVJYSIsGXAWV0/o3d9ISO6J9BV2lA5NV8Aa
IhxlF+x6a+YaKwfbAmTFkA+6nIw6DpY+C8BX82Rvr6ISUqjaKWsYZ9/erhcD
FaHxgCeJ5F+tlMIHRPscCw4h7KvoQAd6gqMi1gVrsQI09BYC1Ydi/tHg6MqP
I++HtCm8kQQHLmJKVKu+d1RiDbEQWsV1VfBswvQ4+ifpFatF4S1LBdW3Tgqc
nUpow4MuEhUr7dYXYMHIXPVCKogXt6JktMt86eKoz5Aghe0WMAD0rhfYDlgY
tvmFGdlewyIvFLwR5kAsNoyfk/shj0HWQiKFCtuGY3B+fFMNBj9wocG/NTA9
10PzFhYRnSqjH4aeaQG+ZBen45W8wq3uY46mvgILyU70px4jtRmKr7C76ss+
CCYrBiNdHr7okaRD/fhwZKk6xT30PJBV/lnnuJOI6IMpM75Df0onOWGypSbI
HtiXSWACzCUaOBfiB5lyqoI0cXfTX/6t8p3zxZ7Io222jaAVUm7EF+wQ9P/9
1D9dIEysaFPXNOCYt7QsUC8gcjUR1UVI3jjp6bMBboMKfGc1JGy7QiaIKmqP
83aeiojH/GXulzhe6nrpPx1rrdQ5oC8oxfG9svdkXKA31vRcq6vvs7kLYebn
PYPxnNXJw0GcLdziPAjWIKhZaOx+4jZ7fPOktHuFiEj/u8tmrGUQD9OQ3QC8
jobXFYtvprjYURwyJOpHcEF7Ce16fWDnV5/ZL4rtDM1/TZkyNJN+PkhXAZDz
fwkLQhn1GG5sTc8068S6K0RuTe3gsM7uEHZKcF5++9QWi9U8b0nNJ1jBNOg8
DmHw+wmfa0BgZ2JS6Aht4FgzWjvL04yYSC6S9dVOL/NCcL7k2/oM13pHlOfl
aHDl4i9fMbUvh3dTcsSjjwnUh1Z0b4ObzY3Ua3pExM1efj0bKfmhhu6BClRL
uK8YSKeYFpqN9to/VqUbljc7yTwo2uLJfckgdcgZSRmO+LsQDy6nzEsdyg2e
QWa37phn3JgNvp9HCxtrxOdkBExmZNeG0nAnFCCH6DcoiZMoSyfKwB1qZqQ0
lpVaJgJJbD8B1KQfYk87Vj6IQSmRKkz2Ai/sut0CbQdV8YJY9JnaNStSTePv
6QkvanEi9TLCbyOoMWnRXCQiE8krx76sHXmBpmdYANKCNmb8pQ5Ubaa4Yj0Y
RKY3ka3zVYIiGgFTZfSR5Bs9dP5pJPYpUG+tLoMjROeoTZIOV+8g2T8vv7cL
byrL7VJ1EvMwHw4vuCCHC6fKxkCtV9SSdCaj0/9UfjqUU1mVFLqsiKllVdbG
bRThcE6zVPXMkf3Y2Mo9Yjk/sqIe2cC7eYxKJEBjBpRON8ELI8SsalFKHq+W
UZq2XAxwWWf5gRJf04yd+D2vyt5z74NNAb7m1TdCFR8O1QG3q7rfUhhrVjE/
iEw11anHd8OGXxim+rD+7HEvGF7UvUiqZuSqDitXOgfzi0ikD0hcpJXUsfbv
IaE0/oGMkCRU8XD4PxCLddWMNQtp6CcXSels+pwqLhfRLrTRittvC+k2KQAL
1m7+BJsQsidRMLD3dZRArYhc7Vz1yu4rsuxSY5Rie5m2Cm9Je5SFXHOV0cAO
7uqMQf8dyh+p1tRd5h4s0KFXOrJGmIR8sU5WGwNhX9exmZEvL4Knp/ncTG4k
tf3USZyR7fM9p/ZZARfDH3m4WqFvSm7EsbmomgXnxfHKe3xgwVyRioug8knu
GewSSgQRjk7gZ0uEevLLgssjHlsseO2pQeADM4ZA4beq6h4yykgkgqsnWh3O
DkK0s+hafDkQIU+vLsalInR2wG50D/YsRrZPNDqE8s9C9gIOACZu3KHusHXR
Awunr1INqvxqfr180abd1V6JI1+5TzMtTT8+9lE2fOfyAPmYz1ZhSGDsWpdq
NsXgta919LbaCDpm8grpf2vpzk8wHk/6h4eDKQt+psPsuAze/JxocuUHyfcb
HFBe8BwPgcUnm0w8Tnu57wWlQiOTSPTM0NeowaZrWJqNiQfUOZMMqWABDUXo
f3xKjgfZJRy6brRPnfwA9FqSWXVzAG1Z0Wb8QOCn5j4T/OI1Wf/cqKiow7yO
fKZrcgtE586700vQKJv963Rvnvp420cO8OXldS3PuYPj8Dez+cwjBgaZZyc6
HslhHMM+PUpilH/QCVsU1nJERQspwzJD3ppMkoAnmyapfc+E44C7whwYydke
3UEKnjFMwNJR1l6JmX5Ep1rJF6lU8XzULjuuHB8LqXBv6HCnVb2/WyR6Xdek
l49VptwIdq883/W/4HraPzCqsZWC3Q0FbxkGoIamnhm9DLBucqkgVnxZymcI
HrVvprG1kEPc3UNLYcun78RiJZ6KvRMtSPR9ocu0bRoIWJX/2w8d+ibzGvXX
yXJO+zeZVK2n82gUZxMoUs9mOFYR9D2AC+VNoSng73+XmtYGOeZpjX3Kv9qR
8q7Mt7R+/RbqerApbogLpgrQmBxPQdTKP2MMqG1XrUcTW666vJFuFuhUgmcN
KsRArRvS+cSGD9wn7gn2qjHg24TdbU64PSrmiv3y90DVAO14XmmEeywz/mqx
qk8OefU/dtD0S1OZcl3807r9AQ3rX8DdbCIEUocaoXA3vKb8l/l5r3dN1LIS
2ciMIXifnBnsdQcliF0U0rCrAiw8lDgk2HoIseTrSS1G8SGjKyftbPlY2hTD
GUeSy/DIwFlWFCIFaVf4iQSu1IWxNRDvxJJ5ZOLnNMxVan0NP+R569JI4d5H
OIMThp+I/cnCeBG2PB7A1x82EwUnZ3b6At5fvs7VXppUSRpS0dLVPSjy6pGs
MtqUo5j+3ovAdRdCi15hs5Js9eoEpovsj0oJdViMOgclEbdHlfFlvPa0cq/q
A9RStqqxxtcXndXY5wuySINSeMprSKL6khAAZRilrNWXBdxnF3BZ3ynjhD/W
qltzZTbU3u187blilBLre++/HwSzRrK3O8DVaOjEuo5rDX/IP113PdwRX/UJ
nXYkqQWhGxb1QlYSghkYZGq2wAarzmYDKdwM29aeyiuR7g1IiRyOU8ZiY3oL
LS97HtD+kSXnyJqoo4wcga0ONF/Y6JLd6y+EsIH3Cu2nbkXaEc6AB6nM1BJW
1YUHE/x2fc2rsYTNt4xoSgNAp9cqO+FNlKjHwQZsCbl5UufBxIfjjwLMuVCy
66LJhftQeZ/iXnV0uyM9J08Uxfc0emCI1yMLVJRpRwYOfSujZOwk4RRSSDwR
EuvGShuvL8V4GtoTiD7UUPIpD8Ijd+nr6vnqLpt3tWz6rgrqvYM8sAr0kB1d
vlnlRk7aT9y8oRoWzu1DEZX5DGoMX1p4qzonNPPj9ZUKeAbyEbqa6TEPa7uf
3Jovmfyf6jPcqXzI0F+tq6qYaTgGDuyXjL+DhxrEAlY6r8h2Y4H/rfXJbVuu
ZJLt5TcELQgYW1zrKnrANKfL1Nu9JNxQiEHQPAmNTG3f0marTQ2JjjCr0RNS
vnIt+UZQKFFRzoY534yTPeH3zikBeWbl3AsmG1sv5Yi2o+Kqz3YB3mymCLY2
CztI4FQ9lOUt2McETQFujZXnmoVoiYtKvXpoB4oNd5bofNbn+jqorSv996Il
KQ4auRQ9QmhS7W8gSGueztxFjhbx+YyDOkNiskwA1P4Hu0Bsuq6Z0rvNuKcK
HH+e00w4QYojfIb/mmkMn4dv6SdEVjk8NfUHUMdIF4xkaNSOLXaa7KOGREOk
oevTFeDx70IrOBHGx9cTBHiKBs2dK2YmtUXAQS2fB06w/91wSa/Igq+xC+rS
vD13mLJHeQ9QnnRAXXSonkMZ7GhzZJHubcaS75v1hvDoxM/3CU9T6l153son
lQx6QZQtwoburvjYrC5EQIxWu8dNWv2rlEZ/4NI35YmKjE6fgHSMBDkmy8ig
OGwN+Ipn6JKm0wCt/e9goJwmu+ICSLXFK71z/o9MuoLW/cYTMg0x1055QyP6
+Vl5pyudT2mryV4Cbk7eAGXgXIz+U3AjYgn9G+nRFGNTkb7Yt8InZfdKmz4A
2M86qpxOAn4CSbyb6aoZFoXo5NKZdyyYuSovRYJiewG53Cxm8k5RBVVZ8nO0
OGsUA7hndX4hmM4klJMJrdnPxw9i6Opl9qoR+bz82Q2ep2c74femDWmn2eKG
GZiIVfL4GADq0k3Uuzi3j6NGHkl0sU6oRe5g+VocsoXohhYjN+j4wLqvywFG
G22xu90M/SQEq5YNZDFunfb7XiKRp5AZ0/7x4sg/606APHSJhLk7Bo7U/N/R
DwM2Jgs8zXTNrQBsV27x5DCBWzvFfD04Z+xpgTSbHfe3PbFERmcu0H4wMi5R
V0NIDEnat2eOS09pSoZWWNcNqlWKCkSUhKScQKQ8QgrI9bIAoKB4orluntc6
btcNk+hkUYv/cz/nDDsXvSP7IjSkIrhdikp4RONuyw62eINh/x3H6YacmXEZ
NEZ9uieKylqdHha3YKf6zWLyT1xJF3kGy2sAYsueZexbW0RsBKZOJ0pYAm3F
bQ1ZlrVkVJLLqOkPq8Q71Z2XmNRqbnU+NIJ+RLAOx9+EbptHuFQoHNmxPznB
alj6PU1JeAMydAhBhEr+SVPC9nUyPUc5oG0VTWIiy9vWrkJmh90yflkYCN/q
DId4+zu3NsgHHGw981SbVSk76Z1DrvMvHxYONhwNo0vkU8bwd67xjfpxSk/g
2w098hcZ2tNN0ukcNtjXfIBSi8IAmIgKdbrhUJTnIsYUyAuVbXD2uVr8q8iX
jKfd1fcDFmJhzpCU8pA6eQeALOQpLHwdOljnDji9xc4d91QN0YD/S/FkitHd
vjK6oTTUdVED/fhR+FXOBD4Dgnu84Y5cR4nSDUnV9NjgSMlBSzz1L4SQ1wbf
vdh2hRB9sX6H1xISdmee7oZ5XyRruMRdJzJTBFXMT8FOBw0YyFfgicCgag9t
oC53QIyJZfjcWEYiQJURWHcJckE4D2+aJpH5qjbBDswScQrsHVcToEmBrM8I
s8I3TYithKOxW3lou0Fu3VdecPbu63dn/pwXXqqEO9VnVeIMd5qXGaVyOGDO
PyEiquSGWBDFtrxrfLycNpW60qCq6k80M2CuIuQFDfYR2MOk8JTQUDxpuwV2
eRyuNHpwPChM+u6XHjIY2dyIaW6wh5OfeK6DJO4J6WC9m5KhPibsKEprss+6
OhuTMXYEicVDpCla9+UqN/xSnU7KyxvASFrmo3Lf1rRgO5vUyWaV+WQ0J0UE
nwMEYPKb4LUEAczJuhSpphzrgaHLIBhFtm0+n01h1ehhZBnsuWlPm4QmsN4t
JAwdXnxwUTHc0/CiJStnS109UQrW3xhB2fXzlYnpSZL6nVhLdt7z4E9PTVb3
kp0G4edVEPwVESQNy9AI9KUMK0YF67CVPRUtf0GkdxLTScwpETGx5yqcxMeR
zcsLphJUFU8cNsMzfsuBdcBqzygJo6rK7mNMxez6e6XJW7+Y6Fba6o+QweB0
RbOGMJroHowHWPLp4+f/14ECGE7dWxk8znOLcuj8LbTcPiyl/ljgPI8if/sQ
DoKrIvV2aA0fyOMllJaAwcuywXvWIdZhQG5Ms+tfIB67Osl2CRYFqssIxO+i
qmYLmD9wKiu2K1Mkn4Ih1At1YCEynpyvfTxio6plx4KImIv04nRWUjx04ZYp
SCbzCs/C+drr0QmAK8e0oQrCwHSOcI+9nB5QrGE16lN2rGirqhtLB+LultkD
wBzuyTiTwe7JwbSz26TTtBjC9BePP33bnBLm/5GSugPS0/kEzaNe29N7iBqo
hf3OqF/gwA+BFeYmjotI3EbwbmpoXGpUTBPhs6rpWYZblkwRkuB/fB4o86kX
SIyukXRHQpnI7bRG2gvsnWlwEmF7Mbw6t1pIwxSvSeAInjHkdiiTuyyjpzoq
isDqvZIVat51Iwf8Q6ng3maVQCimsEVhGR+lMcGuVVo+KOPk43YxlfN6xw8A
kzAJqj6hvUcKyRaBm3l2LTRVzxEh7obTFTbETNsYh9igvtJHhfBW4CnUbGi0
8IU8i1zc7nLBLjchLd8npQdhnD3tExP1b8eHbIN/ceJiHbibjp9IZJ2gbuC0
CW3x2QMv7Q1cQSPu/pgYB4mYGdacKoMabKQpIh2xMnKt/VARmmsAKePfeZwg
H5kHQzzpqHiNFqApnkE15LlnVjCUDRIRR2hc7GZ1UPYwPKL9YXeqemPW6U34
4/mC+SN8ZAs1oDyZsGdbplfSHLyAJJ+ReL/mqgBvOjluhkE98m52tKVEGHEL
uIJg6hkNkpHuLTBC6SZ5pMfy/65ptJEGvBvovkcmK+qKkg5VVWYP6XNRb9af
/SgHp6gSX43wEeGqLwfzBhmVSzGBSmxEVwPwhmO4kFTOUdIDwmt1zqufWzjS
hz3MSjDF+mTw2MniDWEYrD4EFtU7NL2s32AeBv5cis4/H4Uo39p6vfvzwYKE
9C6kAVdmP5vdEuv6SDI27oU0Np+KzSGnA7giiQdQdnuCqylnl85nlOVULNyn
bmtIqn46bzhsnFucfN3b5n15hnRpLha+bm/U6SUBYAMIzfvwEZyB0Cpx4rGw
LztwtW+NBgQLrIVbtV7al/CTF00s/ojmMPNcTP1dvCHYSA8AhHv+gVW7oaru
ULOqmJp3cvvx+VvdjqaDYCuugT2Uo2WoKQrYjqGIxd4SAPucPSAvCr6yA0kO
aacWtpCRmjEMnsjTLL1++xihIwh4B1FcUWRoUX5UzHlaKJ7mBeyNZfazpFoM
iFLKTOVj4rAnahhakPr99R+b9D/wc+W9Rx1j2h1/lGSbRO8B+zQB5mMXdv1b
JWboCb5BZSfDPHyjXcotppccxMDKLy4uh8eDKKjnXsV3pFkJJMyMo935/Bli
z5LYt60WlaSM+I08oQsebZY65eb7wUIFLCMbkOkOAzgsNnZNmr4r4Qod0M5N
0WXpzM+KLS/f6a1Byf2Jbv3/p1jwQ18vcnglnjuzAz9l+zQ+Hf+zqd+ECGUC
/aq4qS1ZRmjiKQnK7o7MI+ceuatocpWWMuE5yv60qYYaQiVfl6Rj3hoJSJ7l
i6+W8lRqRhgWs/HStNq++WROsv4gzBXCloAEQ6TLnpBiyx5a3nWvaw9NRVGY
jVK2Za+IbGRtkhe0nQvw7JLr0Cy2McXXWvPsjnPU8uKVCiKX/qootGkdVwau
Nn2oNyYVhytHpEfH61QL7qzbR3PcOD9SdlFPlIJod+Nv7rVCy31Uq0O2QCGx
WcC5boCu+TgVlQGknDXT9+V08BucBoTStqGNnoolPNtz3PShrn0nRkbcETQx
KVQDUAIL6Wb6F30r50umlN7VO7XpOA4E4znLy6z21v0lDZhRKSPrMvaNxB1c
UcJv3pjEeZBM9C7mUtJ3l1WRXYo0RK9EY4TABfmj6lucuYm0QBqyTDyhNUG2
wKkVL++TqJAo8KYffm1rR+14exibKpnUMx8KEl2OgoNUgVnc1TLXWEjJkyAN
3tFjUkiiNpD5J3zMhZ+zMf183U9fJM4lsQ0eul0MlIqaQfaGPjB3H0+U+tSO
bo0pBsTfaOKquHcm8/H7V0I44QZ/0u3j8OjwjFvWTCfD2SkdK0ZRO0nMxqHY
csTNplYTM+x5ETxTtI066QinFC+kAX9MTUBIPE81fDwtsae4U02g6tTppgkt
k7Roe3EMoqc2pIgsde93si3Rd81wjXD9GFgeJA0YUrkw3oUGDHc15Laf2ydC
AU9Ga5cRN7c+M0RZMA9HNQfAHNsz4m6Dl6aU1BgccG+wsjXbf80WdHCYj0p+
3p8WCEogxk4iLIDSDID77KS6SVWRu5xG9GqnyDM6m2tvnMOswR9RGT/Ygr+U
hOA3H49c0RLuhrVv45A2mx9pr0st8ynQIUJZz7sqc0L7JRVBjiozsCx1dWDy
BX2nKBBbmx6VxqnB+/d4Yesz6kN0A9X+1zb38BQce78l/lVQi/1fz2dsuvr4
5KlZVw3+Uk5pEGeUGoCm5exKUUDQ4bMRcxIxyHyuIXSvHCY/FxjPsAr575nq
iSww1PbsJgKq5FGJU5jqASstsAwJPKjn76xfB+zMtQlxWyxTEadAMm/nrBGY
PB0BNcTmTnqYvzr9SQogkAX/NYvs5bVwmB9PsHlEE3uzkojkZqlONIvH1jxR
QBAxicQ6RwmrfYULyj6If6DSyssOk5JQosKi+011mT5zdqPfVyP14CumU6cw
gJcEujfDCWJ28teXH2FgEQi030090cX6HygHS24sCt8LAbJqtrvEit0E9di5
5dx+4KDyeBG2tzMmzVEDDntlBPw76Ds6NRcUUX7mPSpeRi0ehjhPMJ6sL6Bh
Fq5RW0UjndSDMEF6HOsRbHVdWxgICB9J+MaJY4MuTjW+hpINq5yWzPNx7RfA
AuHiOjwczXe178t94qPIj5xMc7HZq4ocdAJs0CCvs5Wu+tnEdFfS/Jah6pKp
WaBJLEqsto6qmCfYNayZNfaQK4SsCb8aU8raDEQRFrlYOBdozMBqus/AU9xk
9x8f07T8LY0HEWFCVxRgYPxAk++lJpAV0LqVcWv3simfrGpUYEn0MfNrxp6w
EvS7/i2EYx9iRJ9SyZze2+tBZeutUv7FaG1PRcZdiswAQY/VeM2orRdMJ4KN
7ApBR60lnk82YMXI75h8FSdmk3qbSmF2yoLSOGQ33ZrYRheOefu7XhDUmhNF
bwAv1UUD85iKXelMkvaYa7AIvhIXAa6S+T72f6ZKDOdxgIMsx55H3e8aTZnC
5q2jVoT6KTvRrCjsQ/bAwMyl+D20JNEcut0VCWtZOTIRNVPUvJLM1PlLM6wV
OKQspI66PbPnWwv9Y1EZiP+4BZipbEiPWsy5/oiSvLprRnkJ1+ky15t0gg2m
2osOnocODFRnJuZAbornQJ/TBefngTdeAU/FAcU1BB9ohiqLNYD+JBd/C/Wh
/2hS/Uox5QqcrtEppUmYoqNp3eQ5B9kX357UsnC0IRVeu4/UgU4b7fzSZsFd
+4t9jG3DYnsFZeGu0fvpU2pSuHCeaf7Gh7ibtUV6wbCe1jhDvC04/0w3kKrX
Sy2dkXQzpnd3HXA3Hi7Uud1scR0BcooRkWJa9a3phd62C1ISGA4g1Bg5F8+v
QZgNTKUycAkbKlBRwiBoA897qylChcmXsKh9vltuLkio/A9Etm5blKkfPg94
TJwORBtJ7l7ZysBFerO3mGULO5zK54ytI15kQ3g3LsPe0m0XZQGnP0fTBPr7
keLSVIKx1Q43V3e+SP8uMW7oAFMFZjOe/dzBfah3BDBtN1ieP7GclTGHeKmr
NJ4LxwVDSBvsUdS+SGQyud2tQ8bNXAy2aJSSi+jSMN1DNHc8dh0W3lIbWj1g
02Ecz9ICEEk/82YUQAm25HJEalSZNH0wFhRvMHVA4OSyO/2yWJnwlxOG724E
n/hIDGIfyDoY7+wEQAW059qnIqtDv7dcAgRMyR+WvVaJAK7zHwI1EJM6569R
+4Syl6a8/S6ep8h7aXfJnC+EP6pszV8guBCzx83Nj75iuRra4M9IiA0X2nU0
YjSVY9JhvsLHWBWFKds3ISJbqM8TqtoYS0nVLuQvRJnavDFJ1k5byXDQNNI3
Iy+rtXXBrPLcqdJhWF7S4cEQBq8RkHKr+hk1DWwF5GnURX3lcRxAKpPIVXMk
dM0MjXF6/+mQQdEA9sdjkGneICZ0GPH2KeX/nECqSr2nh53Re4ex5CUfPhnQ
AeDpEjJlu/ViMoT6xyrldZpuMBbAqNlCurSQJ0cSzcPTktiy1iKXFM4sR/Ho
pr9FQupVcAxbCFWZkP8aIfvHIu+hsy1aAQ85rPW5Tj5PGn491kb3Ibc+t1DT
0N8JisxPfgcH3EABIU2ReiyQmTYxYQTsAC2vGCfcshe1qdlaEqN+Mxu/uUbA
nvYaIg8l198eMxnvhLuBFUwP94VfkceDvQacKGfMxjnaCzliAKd/hCRmKjn0
pp3Nhu6vUy65YV3KmVIoncVOGzA5+BDq6fB/bs1atObSsgmUl3OTg+4YWlEa
VcsSGGOpN0MWRnYYsYrGwebD8SU7YCm30fbhZwPa9Jd8JyBvnOGYG2RWEg+f
FnOWCbaNbFDHC0fEiJei8CdOaVMLKWA5kLMsPgPBn1b1IPPP3RMAGfgE8QmT
UAzJ1p4FH0iuf5LJkhO6QQqfFhEYfu9ealOjz+tMged4++AyRMy6cBcpcA3A
3LIpCmt3a7KVNEJ6Y+0wQ49AOB3oYcXgRhgTbDY++5vYi3t998/OEA+dVQUA
WhBduOCdD76+fyS6IpPM5EsTh+vmeQjCxUXIs0RmCFZin1MBuZQ62g5oxxGg
1MlTQkDcZ7GJMf32K/OWhJwPNVxh85cP35pf7pQKwoVLhCo+vR04JTCyappt
6u0cIug3TUVlWXN4ubS9vKGQ6/VIwFea9BvfMlhxJ2CYY/q7hs7N09mpEGMN
xuBD528wNro0Hbd2Aq/uRvFSOWTXQa8OPtt0MGQYN7lOmEyrRkaxEO2HGzuX
ffD6jvH1ltuF0GJ4Fh3JPhoMftgyNv+nLVxibtTBk/7BxrQtgoBhITesiFIa
TvHnNk0JDGTVF/qade6soL3zuA8ymmDBtYfr2/GkojdPA3jfcogDOQlVvv1p
oRXInnsaOnGzS70U6QldM8vgGeft9uU2cHGOXJnokWeAoe2wPSUqKgzZu/N4
DmxPE0NUP5zycm8Ql2CtvTFmX8D6JLwnWEKEnci3zZ5clwxxPcpplQNZOQOx
+qvfdXKzXYXs/8TTFKG3D97bskWx69rK5JxAxbNMFmzy7bf5Cqrib2wAI6pv
6H15QECCqUFqLiSf0cyazX8Ki+9SbBfyCvYOb5S1A4s3CQRnaL7OG3MNwv9e
zFeIMuWKOxpB4ir12VmVPQJVSFSryejvl6KcNlZzo6SFUP2qYm/yT9UH+ZRU
JGqErHWlXpOl8M3cLb56i3riscrZre4ehYgYuwl592Qdad0JVttBnMCZ/A4D
KknO7n2OWDLRvn55grh1RykdPi0sCWDk5Dx2dG0evpmBGszF0qimusdK6xI3
nNYRlPpBeL1EHAAKin36Zyx6tVl4TltJkjT+2zRpgyoPXk+3qYfqz4Ue10E8
VkyzUM8Dro0gadPZjiepD9wtfgKzEFgEyQ6AXFpjBt3Zs0sWPe8MKdbkZOg1
qmb/thkAfjz+HzdklrgJ5wHD//99dd/KGboXTON7EZjQWgk/sdsxB18sWAzW
p18N6vGn3+7I6HjllLSnEk70CbRzvOrZvvI4TDFn3Sh6w8Ho24+hywCAaSb4
Zv4230YhJXuKFCZ36uhbIjLI1qwLC4+29iRetvEzBFZKeZjFcPPXis3b9/i7
Hjk8fd4usFAyU53hC+Pni7s0GK+AFQmGQTn+CSjrasdsubyRWM+ClFEGOclZ
zSglpy/QZ1j08//SIBvzIkFfWk96220hV1kOLuGIHiV2bm79Oojv6Mv31HYC
Bk95umkbfT3JR9TnpA9pmswkb41lJwbd2rpJ8UkksYqRfRGYB6vizzAN49Lw
otZcheZwaBsnOfwfdwJLfWwX7eW8vD5FjT7bpfTf2vMQL6FOkZB3WVK/82BC
YcoRytqQqfWyQfrdjNi7Ozo1N5sUt7RmCB8kEe97MtP1uygJLpj3x8/3CNWK
iyVtZHyPJwSBshplF5qWzIOcDULHMjbmgu1zWo9ZZcqIFts2v2m9FVyu2JOr
zzUD9IssJGqI7fNdF7rMwyrlXkYwpRdfo33dCV+iFrb9W3cbZZoc49Rdtvjo
Ggr57Xnus8WOvTVQ8Oq0/PQKmC3rJAaEYISNLLYvkL73BskrU+j1+5g87kGK
ueYqqJdeZVsB4Kg8J66U67g2Lc0XCVKoRMdwEAJSx4VtUC28L/kad2NPh+Fz
LI61Nvf02Zj4h0f1MJWmUjkXctRrJdeuu6zzIYL+ID6VuY4L9GN5u2/qGpkJ
p5kEX679XpsoItuPxcm04BoLBHThIjOfQ0HS4xd98ugi0U/Wh72RZP1jSC6T
++4Is36xRaKbmCYCDxtpSl/hJ57ezKbcsl9cwgAux7E2pZ/2DZ3jaoaxBHYH
rawIMxPqwvmyfl6Lz5t6K+RVMSwhAybfbogiivdQZ5KSnzRuc7y6tRk3gmUF
xiPi+CKjSV94zVbTeJ08HUVICxL+f6b2/l9WRVVhYVldH6J5nojN0z2YIv+S
y+IrRYEY9XB+FSzC0YS7rcbRxCrTs9H77hkTsxWhQuSgtplbkQHr19e76ctJ
d2zvxphb6tBb+cNuvtFvzal4fWQTL6gwm48sU6Ei9znNWjO4oqEuun81ffEz
USqSgS6k7QXnjvsqGkQvHxE9EeWz/EpUW1taBJ6Il7z5+pMG2yLeRpSCbHAI
m+FjZWAUzX75gQLdEn5LrG7IMU77Zkw/s5e1P+srrayCTsGX+sDyeUDl2JhI
YE32rknmPH1O9d+wI50R/Lki/3beY/QL9IqtK5/5N0kUvCErxZwicVH+y4FU
TLlJoOl+VY39jEiOxX8GoqryR2Hd0m394QdoNBIC5BgomiGbJEflFKN9AGzk
YxPFW9nkoajaWrPanGrWXmmKKc+BguNU9eToUjG0/nG9fs8y00qlgMJUctWo
4D5iZLXFVKbntSHtT1exsAQNZTlNPiVdBeCIxHEdpRyHfqa2zMdHMzVkOHcf
SKmgCgGQKaMPmMIILU0lMRqOKUkgA/2AxPseBub2RKe6oAEgxdrsRdueT4PC
93+W8z70u5gXs3hWqLThD+Eu4HhYmUQrezoN+nOGLqdBKWe0gJc8NCwxXU4e
LdwYGPfXxn+ayvmGNilZl5SWEb+v6KBZKGu6XEqKcPLdbfRcRixHjzQzWLWN
GrEukhov1Q5XVbJ7/SeXJMwnjOzJFzHbp88Du7lc2I13PdeJtEsTRimz0i+L
0wZVCpY341CzXcVqQhtMNw1wx8DSKJL0aikkLavwfo3zJIC84tCBvLg/7bOD
vC0g39i3KA4daICBvwy7pEG4wsXN36MXx7G8oBK4y81RrzAY1XqQtdcxjeDH
QG5HjnqXNsmHArGl+4QxulRvyY+Kq2Kz8TaIV0+mqIBx97waREn0HDGSKePc
cNlsGtoIcF+QAwFZ1eiF+UVj7bp03jVW5LsCcHU1ohGzcc4QIqbAvalqeERa
Te5hDkZ3MKYmeB3l8i4bqMumbsK+oQ9TmOrwlpQrKcPNuEhrELeG90hfhStf
LpSHKYjny+FclLoi6KuOtxZHIcBFNG5D4j93zdZgqoo7o2cT0iiMQMx1QXCF
sD/Nis6LrV75s71An+RvvQLcOHU4SpmL0dZuhSmptoYAto3i/+7DtDCaXZbx
zCz0ts5RBsRkfcg81EjNQ1ofb7q0ri0xv7JZHPh++wIpW4elY9u80by+E/TB
/4//gFYgHDDg3X9gxFPrMt0DUvhHpSEpj1IIQsQW0TBmWnagHSzLMR7z6chl
9uy6OFQ2FTZpNXy+amZQz8AXKIeq1NDdA2mJHyl/vKXVHHg9UqF6zNe1+M5U
a2RySeihwHVFtl06TB3CQeCSyMQyQb/gtc7CvpIULIWxH6AiVlqDX952teA6
aXL7qSiDMDZKkWI+AAFmwsDn/8GYkCQLBdNYi5vpahEFP8oHRArpMu6FdkEL
Nu3uSV9qwICvXghyTH+IWURXowgTLkHlpCQ6DVZoZA7uxrdfzh1tck21GnRB
431huDtB36aPU20tVOguJWm8GBheWb7PuAk6nOXBCKCPgyKaNq7AbrpwqwKF
KYGjVgEMWhB1xV0wAKZQfaeqlAFzAix61G836v35Dq3Br8j7MNvA1Oj9Gyjo
+oQ2DAHC/mrWq8YNRK8UcBCJGFyuJ5kzan6Xi6DxqTTgLCFi3SojPLFiHxzB
rJgLB/aeypPiN/H3h5P810CCGK5beIY8Gv62Xxr0kdBlFNtx35o03IXRt/dH
uTo32TMNrXHwCxncAB8qzfDZyNslEnyMLQKg2OCMu4GcTXHgINNjhqlDrnec
Is8YkejgVR25KSjGVYmc0z1o8y4wrYGGK3Dz7cTP52TwDxDUigHvXw1Gi4dB
kTzpiaCZ//dlRsMnZ5NGM/PtqiMZY8I7PUJmS3X/nFZpnGZC1/s1nCi36eZ/
Nkmk684nDerB8LfAT/ZXEdwGxQL5sFqqO7e8+B2Fx/8/jak4L+/B2j6Ir9DF
zXanAf6f2Udoq8wqYsTP4eRlZtWgdp5sd8H+Uh3epuffCYnRQPCYOfsHiPVu
Ct9SmaxSI8cBRwEJCICXmMNA6i3iaFxdrGPy8E00Ejn56PN+m3wO+063RXUL
tRhAY0/kgQQK2WbBBiXcrrE7I6u0cQHJZVVzsxhlfnhWs8TX13v2RcA6KrS6
zMnhltxsugxPmDZrqWoNXqfQmzdnI/Zk1d5VzvJT8QEjWfjZ/4B4oGrH/lM5
Y8P8rZOmSoLf+qWgBSHXuiN7aPdxd7jNwB3dLnb9YpFnZUPHxm8ltf8UX/qu
Eel43wtAWy3DP4lBhOOqScacQzQ38hGT+Gc5CkTiGqLh8rHnChhxoZLpAYm6
+mJ4TmoJtbXqlE6J/kvgW8HRmc4sUx+y1Y/IcvhzF2rz/XixP7fmtAvzJrvX
HfhQe/cpkaXL+Km5mO60cB1VnxnOloV4/PvlfJYnRmDfhwQ8HZgRUuEdJHAQ
H4x4Dw4YSeK9WX5Ek7qlz/fd26MkB//9vQLfbOdP6nhcr9GrLWkG7Tt/kD7A
X1XYvp9vBwTa2NTTOi59xzf4+ze/dy+0slGSTuVd7A75wbqpvafA9x/NgdsZ
Y2TSH2KJ3xMY5gDAo0vS9ubSCSKGM0SJ7fOcQ6e+ntRxvOZ9Q0xWG91TbSb1
FbQDxYR7dALq9TCU2Q5AQIDfeMeiLAhoYBc3rOaZh3ZAROL1CdZvd2qrDLrH
lr5aBl6XiBo8t8vOkOYXW5PRX3uB06ncTWxe4ktC9QYiEoNzphS/sBAjKAx6
Y/gtR3Bk9V2ZfSQFCavnzWXgQuKTJbvc7FOqzkYvNg2j9hEI52QM2xgKWHGe
Z4oMwUYjZ8dLmAZOS4ll6wNXkq1mwpIX5cz0DXqUx1Tou0HQEi/7tleT/B60
s16JOWGJUzMH7FaPVVXUagZAkTJEFluPyDPsdU1f2lEBWWGVeKv3auVAVVug
x9nYbmqmUn65IXmOHW27V0yL9i0Zhvxl0zSP02j9mMug455sSyMl02Ws/sn6
rvo/sGBKPr88X8+Fp+IjLNCyrwNF7cOFvPWnaTvzvFUIf2xGaNGWWiT6+mek
ErIgwsLV38iEndo4MZzquPJJ9VIPfIkN6XZJeS6im3TLhm08b1R0ArQvTABD
/tO42JPhNK1v1WkbHKG/WVo7X2y6fytP1rMQTCt5QzvCZwx+jswtIWL2soki
jND5FRjf6X9kFyLBMAVmkGhmX2c7P5sm1P2ntlkDQUwgEPK0KcSYB8e/LAPD
SnwDO2GEZBhMMsXi04tA7pHJHcLu70MZmWQP5eW61fQdpSgOUHfNV1JoDXD/
zgm6Es8kQF5R4eHXwtPfOA27i7B1OftFwqRO9KVpoXdhwM0qoIOdEz31JSdq
vUGmIl6oUnIftvDPl5nNnMFkwlnC6FfLqQv7j29prOw+LfboRq4MUB6V0so/
wvjrKamHVm4qpiEhAGrUy6benWATowUvZty6BhPFeniD04M6K4azOcXRxqhN
4hwCJ6Ewy9ZPoXFSARF0A7A6zj6bfYmnCdjLDy76VgKhDxuXZHYYMVL/kzGh
uDnc/lFw0cRB5jCc89rUYi/bkn27Qqyf9TqxDdJXeMcCu8TWq+SVce9B2Kz4
zi8KYxe6NstqSoNoLuPiXLu401QW1MqTM5dZMZD1SpxhNJwFdXWfHQBZQCOI
qYcgLOL26NrHoVC/oTuOlIqlSsGqCFyVjVcNwnXkXGYyLS2qQAU2oPj7F+l/
GVol7mkVDNvL5VsgKE/jaQYR+LGsUsfVlMAAJN6Hhp6mTgr1/Sxw/hXukpxl
VvB5+IetcVwF1Aj9ifIq2+5++ctatLaMM/a20smfG+t75ybsOio4rtxA8eTx
xxLd/AFpJrPGoyIFcZX+7QtZ65sb2QLBZV/Zinrqh4WcEzIL7JkRWUQ+ixcQ
b3bKCawyLz4drwqhd6QT4mbfHaK1+qz3Ka11gR/0rZ6UkurIGEk/Nyb/ZfSR
IEJoSBpc5pvwakKJmR9Sr8xsebki3Ky3uOde9Uag0i6MZZor7b/csYKmhDpF
qGCy3Hgw/o1JYfWd74wuVZxwOpxx1OMWT5O4b1168AWEwnolkvdJbB69K92h
D//8ARJOtnMQcZ1x0+s7r02/qYp2GvsccSZbNdgD6wERCW+R5/ac4qaD46Ii
Nr4VT9VP4jE5nUh1S/CLPKLAdFtyoLmchknw5Lr0xCe2BQMAKTaqceDSs0sE
7H+brhQkqK4YAiqCl7inN7f38hAKfOf2YA7qe4AL5jw5G0p3l0HdT4BPrgED
xU+X6LN5OHnXwNfTwJjpBCHkuOIAkhEX/BhRM/Gwbj1PRi6HHVCIdsjkwd7x
xmbMf7ACaDF/1K4tloredX13IaSO7brXGiLaNJx1r9sg5Koeab7ECGUwK7yQ
UTNk2FqB/0V8388ktPGrGzl537IqIQogNmdTx2bhoAHZBx0T2hiWcEVQOirL
I/KbWosqtR2XFtFdYXqsC+5ZDPbxE6L6jvEWVR7J8yJoc0TMVgUvSOJLiL5v
PRsULKvbj1YHAmWyKMh9Ab6F5PaEYnh58vOYfiSDf04m6geLl6X3vHVnzVOk
qS+hdNBQ9u3n3IXI3vNDCKKfF02ZaRlGoKWzLB7omh7RRAUK1AwvYUdodLsU
g/PfVnYAsFMoCp+BJcHPGVMMzjV90uKqPGU2oR1TgF01Aw2IjHOwYZ+4eSXh
0UHrxe1qEYusm+TlMKXKUU2VZ/bDQ98niEEr2eTBYgOPla5NZ50O9baKVQ1f
+5IYPmquKM0oe396ffAcnViybUB/ESXzC8tYPjHnsI6kUrd33LEfkpzpVZrI
gx65YmctDA8H/pEbdhBmrlKMMJRCIfWIpc8daUio3UNLNz4vOtYMFHs2XccH
9irXGsjx0Lti/LFTYCrCGtR/kIcuQRNHVqJBoV/dkajly1LzbGp2aHrgv2iZ
+uypLW2QNhcTu7L94UbI7wpQhJRK5jkhz3DMogzDLB0e8+GRRXcCYap96EX2
iGYARMSh/5pB8p264QWsbdexN8WxfL9fO8851bZEzVMxC91aKNeE5IcUsk47
pd7J51b9Mgs99ChkVTHBjUmxL1XLgwsQbzJV4P/SalV0NdLc+QJ34CiSEFjA
Bd1dL2HnY/x1Hb2zf73iqA6Gba6wM3dNiT3tcUUS1nm1V7w8ZOnJoP2yPCHX
xw6T7Iu7LM5CqiUkoejIpst4YDTqz7/SWWnNOhMLYbRCnRNGJeLE8Hy9yn57
awiqgsQHOQe2ZVgEwJdU2QDSSq27zZGKP4DLERd06Le1y1tOfHZBPfwuYOWU
/PmH2naKxXdxQy1rXxre10/TrjpUSalXLuhaTn57ihpQE5mc/EIbY3sxHvNL
hP8T5udHEYWjotVpvXQZuNNMHPhiyKQQLfu9R7xetVA1Alf/us8ZTQ1zevAH
A7MhphT2H9cmFbctAbSFOJ9fg4nj+4GsW+cDEC5K/XoI/fwb4AqQMRmtK0yo
Cq4+6tm5vGZLaBQeFuLZZcUwVVhtRTz1ez/4NTx/PT9GKEbsKgnGBWQe66Q2
IMePYgW1nZlbxxk8Kr/lwUePOa+kxx3xpuMYad9ssxcsFtwI5CYvhHbsvapE
M/1psTTlX7XqyXBlqiUWwjCs7lrBvNaJMcRS7DqhB0Gs93X8SRW7DRjW6G/w
Y4rYMkQeChSy0jP1KcKj0p8yl32tXdIbNBWiVkKBoBIn6CvWfGBcno+a4DD3
sOVtV/jW1iU/KAXMMt2H/27nXCwk68ixWeh8xjUjWqQbnBfr/wFjMJRmB0dg
gYSHKJfl4RGe9zg5q64/9Dl0n/Wdl/2wrg5wNV8ecv5UR7zqphVA/A5aumoH
9m0wo/e1ZVO2ZSF8dWl63qi2fhC1oNubL7mQVkU7PLPiK3aUK/q71UpOxrhq
CEv5dzcwf25zyN3+9rm4CugdU0GW5wN464ShbWM3aY8NjHCtrw8UvufxdlcB
2E+15M5siXipmBWYbO9dlDEI/eIV2x+XNTKZ8BBcUToRzHvWvkKRo/l7f5tR
zCiCp4o4p3b4i1Pvb/mzBykLJC2M3M4va1TQd8I4eE/TsTOFADAZdB9itwLo
MsB8n53zlkM8j61StM4Jj1LneX0LFZSEow217ynPmBh57efX/gUAPn/o6gbc
mpUOKuLZslCCs1w5b7nsgyxEbTVAThNNLZjYNqrVDlfYSs8Q/F+OGg4l6EIq
TmLz+4iSJ+bLmsOmGvIgy/4dRLja2LsgF+c1bEM1gQAqemnbPrwP6/OQ7Eu6
jEEVKOd12P4NDU6gT4gxw/XivfFmsP6RJ0i02E0LHMzVoJD1b2ht5Ynw9rct
QI0ywzwRiFaX368il37H5awhVpgq2p58csNXcCxaXtBlCHoRv2la8wzLqgwg
uGqPKXiH08lPO+KBDm4QbRMJDcWRyMf9HPB6YaSmZ/NZWAlWwn4xjO5Vp1cG
2IeqTVkDqVfybkFi2XyJhrYbgciyn0x726PHrSgbFp+vlsSdjXE9FBhVCfh/
SToDHQiRQLOjUYskxkRx23H9qZCixVBIzjE2Y0jGhuTBW6VVGFBC1yq4ZYly
iPKQijF46NYITsthAye0PZxlRyQvadoLynDBbNOeYjJR9OJL3V+ZKHD8tXsY
S5sx6PMo9QycjtCGvt1Aj07fXI+rVZHFbQVzNNNl/lJ7Ize7DmD+GwuYOh1C
VhqhNxNm2udYtIChVlc/SKcBq54HXzkLhaS3l4nvxFZU+/fhrjpYtWQX2omP
fA6BJyAP8QS/+ckiZstVERHlwnI7ReI3QLoMf7EzMrTc+ZWH2HxM8nWb5Wa6
XrhgQu1xmdZr9fpWpVWADIaT0pH4EUNbPUiylSrlTqwct2ZE0ePw71IllsnA
w8ZUvUzQKn1X4PUqQHqyKG3oc051ryE1jp3DTx9L829/qk2rTiaEEvgg+KHx
gWvJAJ+qeuy3yU7opISqWMmT3iqsR2mw/+tl/MM1sH3G+PdFcBFV47XoyZD5
vYJxM5hLsVU+jukk3NtqXAHjjsw4dDYr+HjMh0jAt4+GT73jcTFM78mVWiDU
jJtWhwTED0PHgar3d+Jb7oFvv/2ueGw72Ippvf2/9VsGTw8BiRmK96N7hW4Y
gTgtsWkjPtNlSHBaZMNMgqx6I4m1CvEr9K9ZiKTLYQAiMcxDO1Nq06kSMr6P
Tls5CWctaAdbadpom02WY0nvt63Bsi89JrHMR/5uAfVA0z8exkkc8ribPKvk
YeMw23PvXQZJszLTVHNdNw31lBDZ5DeBmGGqc5AA3lrl1nvaV4zo5RF4vhlB
3VztDb4uaqBP6Qy8GzRCoRWL94EyEAee2POCwtXIYc7lClOS3B2lmSzP/Mnx
HVPUKU525wb+a6wYdcJtVlRWMDBr7TbDX4qBeUgcqWxCxGfelkk/pQA9w0J8
o6VKNow9ySCEeYJy5OG428DSW2pYtYn9coLMHgxB6XabA27YxiJ0yxA9Vh1J
wsctaT9kQyUjE/aw4IIrEgrZ/cFt7XLPozX1w6luKMyd2cR6zTsdzDstDIa4
8piLlXQ4H66XDEwmot9IXzxCJMMZ9B2MjvutAsMaFxNQJ1HOGTuZJDGIZ7ib
/wQCuPCWZXGnw5mXSy4GDulTH8CZlEbVPyj5QF1weqzhfNfwFAvWIUm67ywd
Cyhek0sQ2X8KecyXp6fK3to4MzjlalV6wlMlOs/Su+8PqCVo1Q/AnyNEtQqw
M4o9Yna+0tiXQWZwWYu2IBLGkG31oQDO8KKCf6+lTar0DV4nPyK9/xp0agZN
eJn3p8eFEvBvMGFLVIHFWjQDjBfbrgl7K5Uh8Gz5FnIAHoZUZp4j3chZodgB
uP2PeeO748tYfQlhNA/6upwMn3+iBGGNrMJN6QOmVe8dcz5nTKIaEwt9fVVh
uHJFc+z0zsyWyMkAVdukXDCvE+QaslUUI47YOCNkWFqOf7K/EoqoRcI9Fvtv
bBUU5ggsQSDCWz8F4k989omsT/I4zvi8VfF3my8vQ3+sWTqYbg3fHuWAuP9j
BobN14aaGsAI5hXdjLKPsyQe1ZK739F8dWNvUxZOstFPEw+28JdijSQzAQWD
HoZNONJF0ioMESTUOdwaoYa/eKqYLWfrDSueY8qFaWUV5b8gIqj5E1bYbbt2
ATMG1WKW4ZMFER4Vx7DcZVabScz9ZK6Xo+1w3i11r+SxSGzbN6USsadSQhrQ
H5H2GnrLIIk83GXlZi/UhV7y3kysNSAuWuS+XN/ca1/nSto1KZTeZlfCnMhc
38cisK9Ecyxtm9HR2HSKI43/ywQEhxAhtR0Tob84xnVdVtIAWWn1kVpg41Gd
p/XW7A2aDgKw9Xmyn1VqjVJQ9KyGvb7x21LtjszoROMd6XlP7n4rApufhbpt
55LPpc/j4ADhNtRBZ2lcUf63/+7GWnfX1Dyd/54zw56a3d7Y9mfs8CyMiLsh
dPAqIPMKy0wsH1G5Far1EeNp511IiUY80qqBYEj9j4PlXaURHRaTgNs11DbK
qYd5B8Ijeqnb6XzWnKB02am58EHIZv4HaX0/HMP03HCEbQOa70GUODhak4sA
yBRZ34qVMpDhYHoAEUtN3w6+ll1P8A9JQMukh9sijLdKo4mqMfzOk5Ldelkq
PYgmN/xKK08kNkMM0oZtEuAoGvctu3eKRV8JEJmqwWZL4Lz455imLrZVpCRU
oF8N6lOoy3TM3V2wqKt77vjnri6AWPidmzBtBE05MAkEqQsqDxrUJo2cx1co
mr8LGBM/90Siz9MCOYy5o24lO2lGins0gL1HFOCXAUKvefjpuhQLeNShPlf/
4/uL8zDneWfX3XwUzmNwoBGCQVqmEEay/VV2BRK/OEqXvbMDeVuA3anAyJJf
dkPbyxbIZD1vhJDH5FptmeQbkRDM+qcQ7gRngsIK3M8bbPLN7XH/Q04urUrJ
pp+cXd/w3TFhKsArUFAG3Y28IV3gv6dHgiIcZ8JuLXdRUFrpXa1wK5ASWbDi
97v3b1Hihv/wWmkTkoeiD7xiC4lP5c7Kz6+8SizYvR8fGBZDK6cqxhjwEFvM
AxWWzg2iGkt1EpYjh+S2DA/WK2amV0liSixXrhOWO1EZguM6/E5wKf3yXeFs
Rp6mT+OfOJtka3sxINeULMTpDf7fKAg4NLnAQc4JTaqWgfc+5MwJmO5ueV6M
HMgLANWBF24wooDc6xIN/su3b240GThVDOmPtyUlEpX1XRv2hdqzi/Reba1w
4MPLwaWIuiIscyz+8TxKPX8WtqLLlAyoiioMRVLthItMCuDLvmE9eqYvgqtf
ytPf0L8XTVepQanGYAMTFeFJ9sRgtp92ldIDR8pO58zhw8q82TewLETk4hJ+
MLDVrT+0Fd5PVvlhiONHzmu8VxkTlmZEUN2+afcgocRDs7yZER3fjAYaXrpt
c9+bEPO5Dw0jYIGHzZIPo4As0CTCx+pf5KdUH+wmfPC08mSQcNGwlJLo2JZE
lJKjA/bGdaZ0QYpYT/t4I2Cn3J2ScAfkS+aDPsuvyTQL+BFm1hjLtf1MaL6H
1zv9ZVT5+OOMLb7jmYv/bgCltyrTehu1IBvA7tNqrOtPEKAx/BYxV/QhwLpU
UrG8wz+AwU1wn+G1ZqRDnsCfYZ7OCx/ZPw/JJ/xNLN6dnzwk9UBbKuhugn15
2xHMD1USWIdpBYdumNO21kdYrR3IYkRNCTPIsuSo/Gj9CDgFSQsSr2t7+6+O
3pBV8Bxmyg3Ey1d8BWfVd9F99uIthCOk8i1HLuBFjcMK6A5XCYCkCRKqzx3P
THTjMT9QnMyLYcLKlv/QC9gCfV2juiFfJNE6UaXM8PEauwes/04EVKyscac2
zfCEp1iJsiSjQxXYx3J6kn5Eb5KCuT+L4c3EWVvqXMY8BYy8gANtgcqOazFA
qT4rprOzltYP1C3ci5JqN7+GV3HhbHk5EuS+DK7K50f9V4BAEq+wV1soTDzK
CV5jj/cTLvbpzFwkibNG+H4zuf0X5btEAYCWsTfLNp70T6143C39hzX86lr6
XKDc2Zex2kJGR+SqMYcYM9D4LxgI5VqEpGcA14ut/nqMCRErg1NxtQlgLI+s
9h2vB657xV7hQgJXx6sm+hkWIQYOqyT0CseML0p15DZ5cZYcFFBaqtVqzc81
uh8fG57NWPRcKQVY6/mb8Ut/6MKgDEPFuPhWfaKeIg0DbXRMf8rOWzWdXpoy
670WtV8HA0A3XUlnLSQwDqa5WAbhp65+d5YNi350IwdnxKh8bNgB5JvhEurn
B1r6zHKgOI5u1ZRAYC8vl4Pier6V9bWvZQw0e5/rvonvdDEOrA6g8fEKgMlB
eTcmjE+YuFDweSTZ3+Swl6+Xv3zUXwLGFJ/gHnENhjD/GiznNaNS4oOu4+pD
afhLzWRlevRY6Cz+eu7PWjsZ8pIUc6MDfA4W/pvPYhQyMoLZrMguILox7PdG
+ilXGMx3P0tS4ZEntqyfC5qUMWw7qg6fJ4czWnzYcDOA1ZmQV5kGGYH4Eq5p
tlbNgmqEK8sKmLC5BpxXjy3arUau7Da7NFju5XoNZbDu7VUuPUH9y5S0fLgT
VmJwEHqRCzaDHeZFHFx2gVWg/QMTcz+qspC4h9fWjag/MQ1WX0RGeLmE/jhN
HSyCX+rTiCxw/TzcluCezej/8o4GgDdJo6E1A4sFVV7U7Sk15t3xO9SuoadE
/mr5s7tJc9JrBezV3Qs3PIGU6aJe083lKvXlgsUl1ZxwwQUpqbtcfJPHrq1f
FS8RLh/wtJBZemwKhwXz9A6a/CG4bGVFXmnt2xp6a4b1/XzZupqUzjUrMedQ
bhBDTlFpiytatgtUl7lA5MPHrHub7OISllf0rkC9CT/RhvbM6MZJbPNbT2hY
roGwyUL0durKmnXbVaXOJPkKwtGI+3Keu8Wc/fVABLFC6tFuSNC29v1UFMTS
Xiu4M7W1azz5yf1yNzpRfXnv5PILAQY82xIEEDNY4D4qEgNOArh8GXpK6HX3
1eaUryvgufmaVOh/8sIM7Uqp/Q4IjlCNWR1Sngb0Qr5Z9hM2AHog3XeMevLv
vwITlRJ7wOPDRk6ysFFu02ns76UH0fB+ni5k4B/vSF/5l6yebGLtO9/TA01i
1fuJUigHCRYteCLeykSw1CWw0w5/3o1KzFF/swVp1dcoSco/80PV4+BOk81i
KpjPv+n990OJPowF63FnIX3mvga8brJSndzA8VEwDLARmxK77oR3JCr3J53S
YMCqq93UfWqUeMMDoeidA1fSR3ePT4kXs8vu2XMk4X7ojj9qZW08bTi/E61V
f+PFcSgwboNvafO4WXbq/KmRl1RiSGBYkgCRONw+nFpaEd8RXQAZwugHYZSW
dZao2WlO5pkuoMtO3yEPHrhNOjZF4sOQsrmqllelAiyg58oII3DmF4/TyLLr
ELPwAjS5kXrsmXMc2be9k8Yz7xF+YdXl8ILeZBIjb+De7nzcBQYCwZh6s+qo
Sd6TwBE/ZJCvFs6KFndRQzL2Zqb8M5VbyQwRPyUWaNMxn6jJLAv2/SN9blp8
E4WS+ELqeKRqxwZkXjL3dfgbkVO+Mw/xOMinBOJ9TH0dsX/HASdWvK3omYtp
l2oBgyOYR7zq2LgdHt3q7QkoCvT4AkqdaByxwZQssoax7+7nlgIe15U9vNYa
4GxQKksom1yfT4A3Pd2eYC+MlIBX/ZYDYbwXe6kpVQVHhG3mFjsgWAz8rs96
le8o2uEAC+LgL2esXPnPf9+5+jSzwDALK9Y+ZTGQo/C/Xdv4Y8ExtHRnPmYl
d8gFlpktn35zl00ueX3AOl4u3qakuMJIc7Rab8tF8N9/k02MQpOe0hGB2SKE
s3XU+4lJAX7H5EAyktaYej8Xusx+RAf5ofcwB2y4BcEkdfpGjhgLhDHaQ65d
e1IPcMsMkdHq6JLH1SAHn17X29dUO1+kzXKyNdnyIIwpBETbTIrIurDSnNql
Go34Bszt0GOft/vSIdA/xazt2P/TWMUpXGRFsZGJhftNCCQ6r5vNnvCwS6/U
x507hohmp0opmLf0ZsSYGErDrKc5Ed6W67nshdrFn4Y+2PINz+hl2YKQrVcX
n5kEUqwIaK9peDdU9Nwb0DJtEog/9gmMOEiwUU4iUIXjICdl/aLc3LeC5Mga
WsKRcr22fNqZQjV2rMJygXXHFIdiuZJCKUzGRjj1CQ++OXkAqWxHmQ1WKn7t
5xpjuUX/mwXuRTd8YXp095cqsTf92dJSXLjlyfgKtVyqzoT2CzIzPCncfK7r
Xw6a9Km2rQIOstH4MjcT46valBQvbz3XC13eY3JxZZTPIz7qtw9yHzXregQe
x/XJoLu0rAHYDHIHyixan5+/tqlsKTDoCIWNZdE2EYleZ98NOzWEbLN5LktJ
kPcKgexGMdf2MQaLqOywl3Ki1YFNoB6/pEATXVWB0mFEIYs1vEyaf6aZE19+
+8LfCa/iuhrTa6ntsZcYHj1hykArwsMLEt0jyqKWzczXuR6ont6H7p3dH80w
Y6GXibdfHkZ9GbkfsyqmHeuixSFgLo06R2vJAUewAdHwigQiJSBJW/8QlWbV
cv525bgKHKeQtLqSgNnNX69cjB/hq3adXiQ5e9eM4lkZ3RzZwANoe4dav8a3
hyEgmBqtobz9FD0cMn2Sm8zZiB99y3jpGe/V2AB7XtsmPkgAaTytR3HpzYX7
DV9TvNPj7RRYgJZTB495QIA1p8sokuVnXxUmFWeTTPaS7iiO1RVKzciGmmnO
FsdNxgDdnl9NKUo9EBLN7/lmIQ+gA+Pq+RNvNilv6/r5e60oHNx1VVe90wxm
98tj5k8KWqATqqUJSuX0HV5LKu7uXRZu6KL67Q6Ls7A+9/j+MtaREKkY7FB1
JpCwovSRgatXWueWcpz7xb5OvWhFsgWzFg0N92qc1HzMtIg59nGn7AR179U6
nsMATPFyyeeeRx7NFcRnGf7sQDmtDcvfixMsFMHA0MAlrBc25++I/A+qqakm
yvbOVZP5TNcSi7cLl/xTCr9lBu7Qo4vQ2WQpl6RPhcSSeOL3Km1l4up0XIM5
5ZNfWvX8W7A59LnECB5IFhUVbfvQiP3s/bLXe6uySTPxFck9fyyad1quptQX
glTpMXy9B2iSd6yWFkMIS12jYhCkICLbMOImVx3UMRICpiHOsyWJzGa4QfW7
d/bKUcryQwktc0NEy47XudcOqSYLO1Za/yv//QTD6Ixsd3Znifp+nG5ZaAMz
4E2m2DLpFJGB7vYt8+tqEzGOMNSNnuAoi25jZSGxhCYL0G3UBfhDzcHgyZpl
uJCsMVyjbQ19hdiFmwwd3D88mY4LA7c9VGnjqW7xdqtRIvVNZlDcIZY0AtE7
AEH43on9yP2jI4je4/3a2bjmRBCVJPPqxEHa+u2aoU+v6KCoSmNiCfPu0hAW
Yxf/BjnW5ciE6w0XzMucQFhI+SE0yx/lvGWZrii0yVhyaudRjUlRCl/jyRFU
dkSrxfvcvCQJ77SF7B9Ywj0kcLo6o6V1h0QeDp7NbFexgkjcX9H7HRgYCIOZ
raHFQtlHTSsDlOt4Bpkfh0aAtABKdYqm2iVzRcpPzu6SMRLJypumxDYYU81q
RPEgv8lhJJkJa9KQEuYdmIbqVqo12/3urpiViQVdw1s8yFlYZdF1/FMWO1Ql
xVH4viAShrE3jfrc/DyqWMxGw9uhw+pHekd0mxkAcJdC7rLx0GKg/IPpyjLf
wdSAPjeYu9Jb7eGTaAWNnplgfxP+XmAQpPXpRbrcHHDh0zi9EPEpkZXm40O0
q46fmNP9J4dJTgFAtJZnY5PjLOFLQMEL+Z1C+uHD9vKWuCzPoh2fh8eHi9kw
S8HiA35kGHlEqw/HrJx7G86HQI0XSayXwmwlgQkiJAsuxGwN1mh3/mwW7g+B
q3nRlntQmqsLJtjX/nSTgrye4YHpNY3U/SsjZVEyTBjL41qNq34BmyW24ggG
N3mmgVDd7LTNLKtz82E7g8cOFKz2E/Ruwp+SgIEJmfP2e2pc4Tu4XOspZsIy
aLHx0NTBLd1vsmsbWGBOXT9zJJ9XHTbkmVIDdC8D7U5m9NOymsfwypQ/geTw
m4EyAro7AIa956rLSh75X88gfTDtZNjIZq1lRMclsnWrai+0e2MVOeS5ig88
QoRAH1ny0o+j3tEhFmn0H1gSlFZbFf1kVBRNGLjrFmo3rVvfLCOn2aVKZ4Sr
9tLl5Wh1Pm9t9wOE7unFg9SNUeHvGou1h2w8OD6//i5LCrQ+0z5OfH4IUyL4
F/Pa0zc53wwS4TP86SKSulaQK6MmElozW5S68A81tThBVrP7jLCSqmqKIqV/
ttx0/aboGRPISb8KsPtEmBDcmIabUIdHwcOkArvpjHqHvCDd4aoEW8v63t0W
vb8LbOG+VaeHI//r1EFsTiLUWuNLALYJFcgnj9IeRM/O01ZzUsKWtHNphisH
jwfZMps9ZO5idyA9WwEvnvs32o83UfiT53ohZsCd85wHTrkIUvVDM/EpKQpK
r3e2iRjH+C5zWL0O8tQi1QQJMNuJVqLwk+jgEviEWn+y2C2KVh/fhHPPl/dO
uboSa92tyrNtmKbZQO2GxjKnrfIhdOpmj6Lsd3a1XmaIo9AMo16A7VjwtAFn
I3S+1mzA568YlNbIxUOafWvgMWa9sOZBKK37YYIBzgK9F12uVmgjN/oaPuat
B1R3matG9VbA/yNeStVYy7dFZ+XuzE2Rl9K8BLTW6oDBDumoYDgao5qFPeeN
XTMhQ63zCljl91vq2K9VOB9M39RdPm6+2vyKDwqhejAca0sUaODWPOwKO5rl
kXsTDsSg/5yw+Gy1APNtAjj4hMALIYYy1faLm21ED8D+b/OtwlbJQEJcQ4lO
lnNgCpQGxQRy56Mb/TrT5SFdiQXkHMvDSM1sPXyVlcg7x7j66D1402BJgYb4
feHj4tlfBhZf+qGQWGfnEJMGIEsGXIhO438GJlF941PW8JZknEEQRdv5hLig
ViaPIzCLDw/f+X2EK6vOtL8D4SgYkEBPu8hJizx767XtkJCiKgo3DxNnTeIE
6Ee3iUmZaTv/3WBGmC2iDHRdT2qdaIfBE8FQMxZRWZhA3QyBXgEaMl4fyi8a
MoFf5BmhDjO4tMI8KBuFodfy1H081n74uPR8NrrPQzk5clN84uT9GbTqIplZ
JB91yccwQ0zQ1xb4xuvS9zUHxJGSOvbyn1mgvExQ/d23fDzl1a/ju/ONhEuE
mZViegFatLUEWH0NFQa8E5/ENL7wp8XssUR0dMdp2OHb3eN4uQoq0k4lPTGN
ZBM7ctAAls+i7C5IDMhgOQBbIi4hmXstqyQ+iEW5EJlH6t2kSJKQ6/zO3fk9
c5K7/kFxvECYz7V4braKLPhzAuEliyyjWyV0evuvPuwYEWUQ4iRZPuCZo/LR
gu1XHPOJY+NrVKyrnW4Q4PCzxF2nG+Pwo3l8N8BcBUZvyrxmXCjNwFXCc8Gm
bUdev2WSGJriK6rYkSTFjDUdMyxp4tXZw3fCRPdX0mPFE2RKOreiJ48wye0q
6zVFgStk90lBWLJaugwTcTtklrPvIOSHcDsF7A4b157UIxd+ANxvg9REJBGv
VNVij1JWXPslDkCE6c2EYge4v0HLrDuCCRBldwnFYuIrAQOeuA4J1gQcCW/k
aO2ZYFBZx9DPqj2XPcQrwwhBUAF2sB7BlS0lIgM+kIRLHeQlQN1ET5OwmL1l
ExZ3/OJNtjj9ncb3lAr2vJ/3ZyVUESD0LwM3tg7sHcop7d4nGeyAmu4aOW51
CGpoQYLUvQSYM3z9FtDuzikShj2nTTso1lMqFkhsdRHiOhkbvdybJHEgGmVV
ypTtXg5Kuf5g9bvtKDzTwHVRyMnQp/7tvC1BdUUEMATzVa+nA+/1X90jNnJV
6MMfxlPn6hxGzTKqmf9GS3P+55HHcmHhQTSCdXMuFhKTiJJKdX1JsXv5g0g/
YwblyfAYtkjjOMGan2wxuCNUAPb+ZQxT0I2ca3kEcCrFSQmVUxpWnnTANUib
vpXR+lqXcbU0iPzsigft1BJuwRjbWxKxu4/OQHNSWQ3Mqp0J5QeVoK3qoVJf
7XMkN3kMP2Dp9q36ihuOTIwNCsvZpulL+D+WEoJcnnYq/k/TwW9VzHQhr9P+
f1zxnUDWtxvJfhm4Ds1lkU48Bt1QxQIpUe7AmVt7Uj6YwMuAt6IE4bs2a9a1
D6aqYD9CrMBlmgsH0zdI4a//zQIAbr6zUqytI+IgSg0eJSIxs4lyYQGtprIc
8QeyL3Q5WiTfH2RKMJ1K2OuHkX70jX7Q0xTMoeuiT4oQM2WOIXDobEXbPB/W
7QhE84/jfJ/z6N4aVmzUn9xHpFrY8BvX34m2wo9WTrRvQkafQ7Wtrtcglr1v
2Y3DaPPMe/VPdzxG9bTEYioCkywqhanSd/HbaDjnZlG+Pd2N7qOH7TQktBMi
zY5O8LkrArQNyr13mfVV45rrD5/7ae2Hrw3KydaTQ12QIQkxfhZTpf8HFW/Z
2+9OmKxfvgmmJiZ1xua7mEgD4ZSCY2fU/3tWU75V6kX2tXBxAkGicrv9hUkK
mmu6y3XCqqHq6hLlpaZZqUfttJsh0dOIyIVdjXJEQppn25FEUruHTU/CSWqj
Vp1OIPPYTCDPZNOW7HXSwSFApDx8ErC2jmKyEJoWqZ7bsis4vauyCYkG+nmw
qQz333qzeU17H3E9oj7CILNfQzeubSFR6xKQxsReMnt2E3PnypvYnW1BbCmV
HrkDgAMscg2m76m85MSv0wPi1qFYwihdZVUBBXIKJtjfSkHh91L3kYv+eWc2
9Je0HPg+XBIeuocetPTrtocy5U6r5Kt6V1pb+8kigQCrqhXVruysCo+NEzA2
KoYujtiq1+vjW8Gg1mfM9kgLeqDpmnnvYF4U9rLwz+pjCzk5yL5WfN2htJ51
erIJ0qG4CGhkEoTnNcc8F87LNGEG8MS3eel/4EJeEd8ZX5eQEzkhZ9zNw1Fp
C7RybiQADlQdUVTepxem7qKHWUgtCW+Q2Wo5Dk4oz/dvJvJyr+DZ4xaGRDQq
IXk4L2iFEZVoZz5Im5JkqRAsfNGQCweZDVbyBtPViusVPOwGXvZmwHh3fdaR
BalP4O56gIYoSQiW8aFKCOlB5sN+CjN9BSndy054vBWb3AtkhMIqckdMP4di
ztYcGQbkfO2hR915mEJ5oeusumx8PLO/30gQupBYr6SwqU5lKzB31h1GzmtR
J6Ow2V7I12L+t+pYWW8u3FJiHf46qHyWAgY+Pn9ojLl1eGsxH0iz6nWJs965
Ja33+TSdSNDilbNo0Rh9qjmblRLTkgBcaxJ0yQP9wRioqviJRPDZsFczim1s
QZIbn7WP/9SbrO54YdqbVw3jPNOfYujiiV94HZEShisITbu+8EAJwiRACUZ/
kvZKdIfxWzX6ulAjWb2GFA0fcBndvYriLSmSGq87rrYjTa8u8PfJC/FBhihF
rI0v30IdcSj21RAJMMuYoERo6OipNZxjKUaRc9h3QoBoEPxCMDX7uBkJp1F7
EHvAMsVhijXKLJ5nzEYVLeOhK+Iz0HQJqKTmdz4wNMxNJf/WDNPUIKjg9rmj
HNWV7I4XswV99NSPdZjhtb+QjNKrk8eg/Xw0B2+kj4D8vG4BTKvcrxjWvJAz
9eaNZcQAyA48nszr9SQCtvQ7F26vgccGOqagWlYQps4dStDr1xuMxMJqo1Dg
etslCXbZ9N0xfR8SnMuC/1OdGVc6kfF8gMtnmnHAGPdx/nCVi+mOR/XSWNAX
UjUG88+GtK5hXYXW9sdVbrDoA9lqoa2NcQ1YhLtryF2rXVsEg2Ep92H4778h
90IOjMLgUFerUyISUBUd/UdsHBGLdfXtqey5rDt2jXf3eNXxY6pL6iHJByNJ
OyMNCMUvip6cJp7rVEJhDZbokF/hElD1bLbtG6lyjOkiUmhFvwZdokbo05yO
ZFdvzBixhG+TgtfGtjfMiKKfcDhnEybAnk2eRL1Q/f0Vi2V4QnFX4mQd3oqJ
rPuSbh06ZOvJoiy335ES/aCTAiaT5Ib5fcgWwik14tMaQ84WVeQuCqmXuxjA
Y9gjVYc1YOw4icJ0dsARrCdPvU5TivO/9pe/Y4D0gOTiJiINMbPjTgu09mNf
tsRhzYsmUaCJeqcVIn0dlD9vCAsqwibyyOAILEKFq8+51sDutjtpI924BlBi
g374zC7V2OadB8eoo01MLV+u2pCc/929HUjDnkY0x6vyv5T/fRyv9qow5b4A
Q/Or6jBge1eiPI2YAI+mPgNZpVqpvjRgeZ+Iyfm3Q7PQj1r8ffm5k3G5fxl3
iEI0XdaLlw1Fam+LCuzVCxVyJ326vrgiYO+UUUlXpSVYzShPu+0AsHlBIkgl
0HMrwRAzcFwZJeh+abOdjvh+MYj1v+FIKsWrH6+hWT13e07OIHo2uOJfxnSi
EDWQo615Ux3ZL5Td9dYOIJj94eR2RjvkI0RRFrrMRebhlI28APjzaGV2DGI9
81ohsUpK7HKNJHzJT++i/oTqYyugERfqx+qwjkzPdGO7ZS3UpYZSZ/vzEB4y
6vmqOKBalR9X2hVdWDVXFHSUiT/ij9eZfSGN0o9eQT+cs84sdlDTDNi8tHvL
Khifs3Mb+98gSdEhOPbSEOh2TGaNH4shiKII3CjLJQTfNqBDwSdmNjT+/VFY
hG7QRN8Su73GyY0EnMvMtd51n+U4C3IpJ2iVLnOo4xvd4u/MIyUHZbNztXrd
QyBfqrShuWi7tu7zZQUfy3oRuZsOn38Lg2v1+shGyWjCpZ19wm6fNW0Y5Rv2
Kk92OUtm8c6vKHiEg85bqaB0gmc4k8A7Rv3ChUYgUnx9yV/ZWsU/Y++kZDcq
oW11fktyNP8fb/btRn4PEWf78dM0qsHGPLqHnsbXee3Ius67R3UlhIgGqHzv
+u1mmyUrtiT1lNWhTIQ/7ks4A4gtBJ0TfLviMTFne4xVf3j0F5svaxjFtU7h
X9w6TJFwexEx8CjlshEN2eV87GHquFbBtUtGqRySOLDI5A8QjuPrjqLNKQYi
br+z2YWIfISZFEdjmA3ZprJYQRqet6uS6GJTs/jOGSc0w/YePtLzeboDzVIu
LHeEwiTlGv3jLH5bQ4bO7S88K4Kx6J8O+8EcHCUAfq1nUAHc7uL2dxKwrIE3
WMhbkVWMH2mGyswyLndOn+2eKh74G9PYoL5h5umcmVTM/jzjdX7ZzCSxDkW7
EueTIOdsqI2VVt2HodvoJUluw75GeoV0NU5k5oni+iZ205VnXDCaoiSY1XjL
pydERE5rzktbULZ57lIZmFCBrAxvGugSgRcxy60gvufIyij7oMllC0ES53oG
tasf3MJHrJAsoQ25FKo/bPkNxctKwau5wDwYNUQ5GzjWVAbwGBo3IjtP84jG
chjBo5J2UJbHAGGSEAFvVYjSoCmueKfKWHhpHCThzrVKEpUwMaoZb24WqqHR
+yyx16pXmTAeSr/2yZBAcK0fG3Fu5q264hk6pZFYc+BA4oKKwB2kqQQXp3hc
UPgalc+CF7lEqT33fJiKk6OuZzK6kTEDPtLftO+b9Ivsf8ctOTIIIUvgZkkV
HFXIlduQoFHye0KLjikllUACFWLHkp1+Y4XxkvcQzitvM+Z0uGumd0xbXq2Y
NujkdJ3bvk6bwmqelv4BcLHuuVCaiMZO1Z9th378BWteTPTrtsihDO+akweP
aKP0RwDGzm9RJ+TQddxUJMxmv9/qgjFIFChtVVCQU+DHcDeiljEj5XDCMIOV
oHHhL46xfetv/v0QkldKQTNPFEdrSLtAa9+lZBXobuqcTIuddXmyWRd6tFkM
jNIxZuS7ROHMRzTqjILHodAW305Ns4rpkug9eOWbLCWVb/fdgRzEZOFBKEiC
lZP95hGSgW9rzr/XWW5wJ23cLKvsc/DzHO+W2VgfpXxAEkYZQHUT3jaSMKGt
y27cOuVahSxWtP9IvcDj/NSw/O+5rCmDbRnxUVSo3cMDulblig0BZBvu4o8y
wJwVL1e4vj5anD7XUrkZuQvG3gtBkwrSqJ13UlwQGt64ns9S3Z4qqF27LrKR
x7y483dz5jmvy6cfLZtHxEFQ2HBq+YpdHAd+AKx/DBgE/ES7DYu+ycpK4UyX
UiCtBwL5sA4MH0J5hDxNyLfrpwTFAg8tcodh3dI/z6BlRbIfJV2qXWnuZdrS
LDR60jwozRw06X6lOuZjTlKT77zk0dBSJb6JtXL8c8XbwawACzhEJzgDS9yv
PC9T1LmKR72APVSvBZFy+2yNzM5F1uToDTpkvopbo4DzZaH0/scrlgLwf+PT
c49pRtliTfXuNY3vV59iXO3f56WQ2l5zBFc/1wa7+kUzjVqHHnGJuPr/VCaJ
yM7runF5vrhhgRox4NIxNZeMP7v3uBlUwyRqrsopTxjPGmruqRaouaA0vwo0
MrUiXMgDlwL9A4+zISr7D4OWcIY3/whXTDrhtX8QLT3ovg0JTPrcuWkw79z7
9vLUIc1qsMH9RuOMnjS1MpIrHTJ4qSgDPodIS8t5n5J/oztS6yGH2Xo2P5q8
fa95B9ufOJVGdHMnU9iw+XbWdruSwewPHnZt2BvmFz2rYGeKY8+og1M1c0bW
P+kgf6gcH2xBkd4DIudj48fgxSfyg/tkbQNSsN5Rs6/RnJwpzN8mmSs/0VQz
DQa3TPrfQsI2zVTCWgaEUv2q9rdg6CiDURDzDEVl5kWBMCy43NbfMY8hn1in
7zHWF4FmiI831U4IsWB1hwhgouLNFif5tZ8G9RnKEIqrimXQ+aIJPC5gCenU
688Z+x3jW+6BmVKl0NKQVih0Q8IMrr9lLNRs02tmz9Lf4pKHU/NH+/nmVNJG
M1iob8IHV3WWJx37am4lBuhcBOKYd3Eq/OVSWXmWVYm8f2iFhANsyvRzCjom
oy7nUbxj1GXPRcWnp61RjLfDE2XY2KxruH31DH1RDd3ANoCk1zfBp6oOJFH0
hLWRwjE6Ht6DVvN0TbPCghmGKkwZHIO0heo8cKpn6WWpXfoIE9MAk0v2kQm1
3V/9WiX7TS8/HNmayCPryHDWExg/gXVxZ9k000pGrrWiQUXDb/9xcfsbTrz5
N+tlRDA0eMncp4Y14ACcaVlB5b3tFPgi4Ys4mmlRt5z9SjWnJQVofT1WCJg/
+2a0K/tIUYp+1uwdvwPjOTOpomJOBzOowx4Cizxcw5ipu1h0PxEOYnGpZmot
KpCMj7ZBod66jUMrVh0b13DJtX7SCGbJ5J20+/QoWpRBANIJx+va3LtnWXCJ
3UU72NPUfEuUqZqF/cdp4nMZWSNe9hGhza2MJfQVXOjow0LQ6wtJBDt60RSU
DW7ZsPLx7lH0J0ef7o0isZRU/wSbLk9i0kq6NCBGLWhy3uFwSWKHXNom5ffx
aylB8gQdhUWWAOTcgioXJECyaHW55V++zdO2h31UFlMwilhADCDdKHu3TL8i
zH/qCgTn5FRAESzyeGa8kcQahx+MTnWxHlKDMo1/jOamRSM/6TX3cK5EZPwh
DdoP5y7Sd98ngIKBoje3emcKI+bdPuj+geO5hLohi5D/07Vey2IWI2mSqoEA
ppyTVARo/K0tiSGE1+fQopMjpiC0HdnVtnLsShKWGybzaoNHf1dR4ErF9SzZ
CvhYZfLEkDWULS1GIFXeUu0ZHTbcELucWxs0Rd5q+6uotZTbPJGUb3u4GT05
xzV8d7R9rRFB07jK3ia+/EJru9/tK+cviMAR1cdwzSNF00dcWEUSGTwWSinG
UFVvUDnOfrs2EVXbxzky62eXwFiVNWEc+k0VALUAwIyFwA3DOFjMjnc3xdti
m0usbVy7bKP3Fwx0yp0yG+Ddn1I0/orAgwnq7seSxNtbsoiF8ZHfLtAy57zc
+iJR5UrwdPktRxD7zMligjDictsA3fmgxhW3p0RyBJsikKVYifiC/NMJ4Vrq
soaAzL6MxGmLdv70HvuTMjHZHCfcirkMDVQitmIwu0T7oRvYmV/X323d62SM
2OlDg/vftjMld/nFe/Bkh1qUbsQ3yryfOjEe3gFe9Y6t8pQcK9Amw1TNioAE
n4q6sVF+eEYVF5yryqQZ/91TRINBbGP5j+d1Ujuq4GrOBn/IW7g4oPIBGGa7
PMxYfw9+fxAgL4KMjC/IV3aJLxOc7wk8qLtLgDqJMpCsEXygTRv9RG5/q5Xt
3b4un7Ci7xPH5gE+TjKKU+BdHFqNISBPjrqm1ROuTjwPb6xo0Gse5H0FAw+N
A3msU79N+gPWrk1gjKowj0DtBrRiiDqvNeoAVbgtkP4X5Hf/SoRk4xbfRyFK
sRsWivyQWF2rWH/5lxV9bNnlQ0xM4IAz8DZvxA9xT2fWI8lSA62AS7zu9ISr
Ok9gIOsoyDhpjtxTd5QBt6fhC2aGD2E2g6pNq2tJXp+VTJ+1dXIUS8VAUSe6
RBKyeAWmodf7hcYCrxDb/gNzrr+BCD0j5yIKrNAXd6RRG0EZ8C6k5fniiT4N
oLogOCXiJYXloBe9rn9ldavQLTRnk/5k+PqiU+dSVYXm9rodWl958lGK0QRf
IllZPtIuwYNdj7HMi0YvUZaJwYPn7b1cOe/63CJPronkE9vH57AEjLtZxiw6
DE2uBAEYO1SCqsQX88lbBRSxhPx6l9sWolxaHJGeqdNPa/18IF877DXJhetv
6KFqfpD3D9h6ItQ/ErkWUu1eFQKkbjmbaydBLFgwSSyCRkMpdYGAhkUnX11N
NpO8pmzfrXqqlpTht8irT3ab8QoUdL6Cb3KpNDC0oYd2ALb94DAaP8HqBf6i
Jhik7V9e15tqaCWAR/1ue2HDHJsl6CER8LDbSC9+oodJEfj5lzgEw5lOyNTW
neoXXsyM8jz/8kvFfFhhx7275ORx8VY74gjtm4VrSgRNH8TiB8oKoNuilhVd
8TnBdCXEBgboSdFW/bnylLy20Lh1RDX2PhMQ0mkv2rclDVjfJ2po+waONf7X
oC3hmv3UnKJB+nGOM9O2vpVelLGTRpfxR7F7CwaP3lLw4yByo6CAxNdV6atU
uy5AX/Yv6/kSrqIFyoaZ/FUNSYR2kp9x1NpLlDcueCdAdUB8YqF52i0EcMIV
rgCW3MJZo9kAiTjVy13ZmuOgdWmvl/MfrwJVJH37SjSDf88o7/+F4IDRhpgh
+HYBgtMqqNg7d6xSc+AN5Uy8kRCkX0CEBgbn1eLqWsT6tPX/FC4NqwWXVqlO
sGi/O/9yrLv2hzdh/VaGMJSJ/eWry7f6/rGchs300Iza9DWp55TsHnCiWqFG
sAyfJmvpgI1ZqiLbZBhtB0ynKeQ4tHM+rdaOORo28wIuwzsidVnhe1EYycnb
QHfiK5ZsQMauKe/XY1LheomG0bPNF5jjP0Bek5GoelmX6IzkWciAJmEyNS4x
V2EknRhcLhDjb58cFuUgv38S7PmvgyBfJwG+Y1FE/8n6+uarHeleQ+luHsp6
WHG2amrTDClm9tG0v6gzYR0Mti/N9Xkuq3q75MvQuaGZcFl9ujvzR5OgR/hH
7wMzXoCt2cIS4D/21K1p4mA0MgtYjRAUHvmLVLqbProl8trtbuA7R4WyEQap
lHqXMSQUou/yIlCj2GpCAsUR/9yo15LKNfA/Y4BW/PlI7ypgfKD9bR3Ypy0o
D4EAk7vTZGxW8Nsd3gPAY39VT9jn4vji6JPFGtw6dJjCoh9qbM8V2yQsipk3
EacP2JOQzDuOv78Hm+IvR8rqYoF7gp5sT4eF/B/QMKTN+ZHTKfgQBBTrI7sv
vWC25rg55aTsa38GZCesO8gTaXz2y4y3B75YicoT8HvT2DMff5z0Ey0bfLdX
p3zWnS/3nPAgEiYJSUcntnEe6/guUIkT6EdDVgKSsILSlP2skH4crpYJyajT
qEGhr0frEyzX9IWx3leWERE6zfbSzbaMoDxEvkLF1l+8zY3coSr2dxPZu7Kh
1h0EQot+MHUW+bIqCS4dG4LnSBVbU4jp4NsG/aDzv6EDffHqcEJdBGaABn8i
mnqOE+7Eu9UQUD59lU63HZBLJ7g2PCk5k74gTe96g2cebo5axp5yKLF53sKv
c8hgAv5QKE9HFfho0mjp1Uk4iVAWeHzbGIvawJxHIi+kGAJYFmXLBjqPpw1d
9dOZPiEhrgRvZyqDffvVHJ8CIazYy9s+/8O3+JAr05prnKGzPMN+iuH6wCAN
dq43ZH56zpqQS2qTF2bgCRpxIxbsrS7xWFGhHWS6dcJCeDT+OV8pJ+Ugramv
lcFhpbsvCL1cFrkq+vQtxW+4/NZda25f3N1f9a0OqvHgzFBkeh4TP5U9wP18
rzSethm48BZb5LT6ThZPwM6H82ZDjmt2fxHtVrVXsJaNclmrCyd+VgCoBDiD
j7cmSV2IAaosXdmQFA9drDTukpUg9fFN52IfJfOCngoExOv3U0ZrHNjDRUZO
5YW/uHnMt94/UqJsCM1B0LniXIc9X5DEjSHNf+S5o4ElO+J5hBgrR3A51Pxz
2eVAJ5ILnGE2122u46oHtzcJB/UBhA2zK+wTqPiIvd+Q1iQN3GpKnmKrbjgN
W9mlxK8P/LEOnzxf3Qfp5/u5FQVaH91HvmT+c1GdQusBvvp9lOfvPu85JfZ0
pvEOGW63EfFtslSWn9L1CM9vnlkz6AsbBo3TwSgBjzT9UT9LWQFE86Ro229T
6gzDvLMkJKcPVrg73Mj5pr6q3rZF5IoH3RyqAiJqnYRt2hukbkv24bsxmqEE
0CJ8iecpIpyvl736v2LWYdG13+1qxZarwiemDDjSpvwqkUzRzA9HW83v6iZA
gIL/PslfanpdZKqEnw2MvHJuNYpXdKQacqwM5LocGrfM+ddOURZP1YP4hIDB
x7XLTONBs7Kjz4mgT9whN/9yB7fjey3N7lraKiFOw8G0nwZg6Lh0HeKQdQfP
fi5fhoh4Ulh7CwJY0fZ46Me/NChJ5ItkrF4f3k+Q2S3RocXGnlWm8irMxUsG
CjSosjQxMVD4VG6eBrUVjquXOv8l45RHnXtSQ/ME1R6KtdPRRIUbz9O/7bH6
6VnzDTYB7gIIp+ovtluI3RLMJ4AfVIDQe4fKj/cRECQIwxf/j+d2dTs/WXnz
GB+CGYlOmRdlx3XPog+Sg5Isll6F8/+98kzMYn2/ld2IdxE4igBhbWG85RqT
UYMTokmrcy1q/BR+JL6xlVrtzRyV6tj6prmnAzfJBje2Qwf1kil0F6+/+1og
4ORBMyr3iU4F+jCYiDxOtFz3c29+ZE7Iyf79GNpAu6FwvUBHh+X5DO37wPqp
BoUYBqxvqKMc35GFi2/0lylLZNpIgBFJwELLbFEX7ZC9Xt84Aj5QiQresjyB
SSy5R0+huL8u0trQNZVycGRYyfo/pI+raSSB+MY9s2lERjxHTW4ogY4Rba6k
xKvjt14DE8HmVFP4elQg3WFuH+y0HdyHtIkavvHO3/hfVkR/84Eh1sKN+x63
j8xvcYNms1g57Q76k9nT5lcokeq3Z5RuvevNrsa+G0v1xMUUtcpRtTkB4/Oe
KT1UXjPojQcJt3ST9F4oAbf/ruSxBu8PJezFApBfb74UBk6lJQ1fqbJa7iy6
a7sbMJLLGRTszXmeAVDA+fewz59ajilo7+AJikdd6HXuuO/c7z+IAEXPDVHz
LEGU6z8YEJFWOhuQXzRbdDirUGzWyqdU9pplbMGMicCKJ42e4eQSzGY1BSaZ
W7pXYSmauOCP35se6EdxPZwc0dQ+idhguGGEAfGN07J9dVQrv6imquvRowfV
M+XgmtwEuzHiyDkUJVAOdIRQ1dbi1oWkcKt5En66u/XjXIgsDC39RUoosTA8
gc0u6IUxVoWb037UF2byxdG7bKOsYllAx7PD8h4Wya2jOL2twiC7+g/hT2ab
xIZuWaptJUeMgggO3iXpoPcoWcweQOwbbWoOkyjNInjh4KIBEbHJBtCJOzg5
BIK69uufDrU/2RrPtq9jmK6ip4F/Rp0O+xP5iqA/s8EsDqytV37byWqCh+jc
8BTr0L5xB8PYQsMuZ3JyBSGkb/r0rGerE6I91bmCVD4UOvtqx8+fSvoE4khp
Sh/atsKMOeiTuNvIhJ4H1LbZ+uf6bc8E16VpnoACgMTGdNJTaN7MzHU7zGgr
2H4XE8sxV7E96vom3TmarlgAPiqOMjOI2ekjgs+KhpZJhGc3nvOjO2MBMUSh
yaaGICr3Z8CwsAmuY1x/RAlTqI54asGVV8/Ce9TffCsWzxKXlK/qPAjyLHAV
MnZoKZT9b4ZkX9LXwVbNfetnasTfEWCWJtDGwGIBKWndYsrAmstC449ytm2B
YEXATr0OjafK8UKyza1dn8cjj6z0z9/x6oVjlIoXMFFwhg0T3b944U1LlTL1
2wa4aNzQorIiFr7w7VumCu8pzYz2wT2QJ6EuS2i6L9a3IHtwLT2n82zicpwU
s5krU6/NaWXDgCO/x5leKqktUY6Q2j6j08Y3vi3UdAiDcrwi4dNT1BUDkjHk
z4wUyKs+63+5/AiEQzZPy3BFA9MCVl/f2tEiUmyHUtREhhFHZ+1OkayEFUE7
WQDThlaUOn1kjkFPdFVn0/sH90radAh8jEiFoUuU4y2VnyQRjqdZS1XeYLVP
xUKg7hgQ1RDrGJMBo6uJBtaACyoItjRBu3Qj4SHYNjITs5+w1DNIeFL2tkbO
/KLNVvKr12V4fMmeJZ5m7/JtLvQ//g18A7SSgzAXLHMSN3r+qodPTSHNdEk9
z34LE505cvCwBQ6WuCCYlHN1wpln538g9AKos+mXQU5WYfWSUgC2wVTAYdAF
olYNq9m9hMXWvbp4MVdAL5S5NSUBHsMe+LMoJEAeWSbm3zJvcKZzhy4hrCZM
E9cqjvkoZHE9Q3rbWeNFK1w5jVgUhPBFxUbw2iSQzAS5+3xbZLJtjyJDtnhg
Qu+/lugf++kf4Qj47OnJJXVuRINl9vmTDxpON6sv++zkfP7xyaAIXtRskunf
aFuwaP6C++KbZJYBPtqBm95DEGjThmEiKhjLiiqMNhpHM/gfpxk44imdUHJW
+vKWaXAqg8ytj8c+cu5Y+yucXOkHWDob31dBw1ZPmmp9CdVMrYHYD/5JuDwq
fQaf9Uadxv9um/6Hg+G1eYjH8Ci3eB44gL2GIvmk0Ch1NAPAatqOkiAk6Knx
/qv5B2ruXstwVLchq2qvdgYrtJF0QCDFM3YMnZX6eWi7LTWMFpkQ3RHGTVEX
MiVS+ZU9nOFdSqmP33RWEeb8/x2LCpxDovlCk9kNnUVWyBF27j2rlsHTEQ/7
dWl/1MUh/RhBjVLoanfAC69Pl8ita4Bx7aZiGYc3VeOGzGsfRVvEJ3QvSkm2
ZvZd8UONRglNQMInt8fnmV/JPjfGi3PP/XhZGVsRCWa2gORsBqPk9bhWSuu3
l9657M5eICL3cGUWZ76im3hqIAa8uWZLpGZASeCwb+NXrDwVRWfslLYFDnM2
maOmzldFwG+CvheLoHoj377w2y7YsqwsKiUWjigKc97knHn8TlBjInCXMN7a
TiZZV/UWxKsRBmRsI940dKbPyKFeKdazOWSFV/oDX5vYcZVMkubHTUn3aO06
+80ZGpgBKaZW9DIV1z0EKhLPjeHHu0WEiYnd7/FVdV81vlBGxvDUlJ3dRBYi
YQsN00hyEi6qNCxvONVM4V/51UUaTnsYd6PqGWcI6VbrK3WL5fUb0oF3+qiT
OdRM/hdQVQU0tCh/wsYgLskn0qLminTXvulzjntDCK7XSG5HZ/no8Jj7KOkc
TOHeQT+ELvGcm1vZVXPIX5OR7h8992W3g3xKn9v0/WgEaRoannyWPiE1rqVN
NfoEyxttRpnBoXefF+VAWHQYrBmy4Bdi8pax137HdWJauVzC7SlWdzojyU4C
XIuUUIiRP5Kciag/2wyY3xJh2fFe1FvihpWp8rZPm04M4pyYrtugBKZafbBK
0ReDXiuqTJsFgvMCDiBkUDkmgY2klL+igDi8uQ5Qsj1ei2Cwm+GHYq2+goB/
51rLqXqRbUKGq08GNEi2BVIm0IyS/T6UJS/Ge2YsPeZMkNZjDK9i0CJgw2OF
zNZ+wXiulvbC0RT8+yjzEo9QC+MeqUNiI0Kn09NivbzCob/feikrrqxxk3ue
VpjAyfEk+P+QqOuuFKP8v5IW3j4Sw5QZJ+ODB9WgD757pA5eAPX4pHcpwdfS
aZ2tpxg/kG6XEWRUKNbDJbocsdQ7WijCeI5GA5UrN+T3eCvCWPdH2L8B6LHV
9vKVKxmK8uSeiUhoTsVFDtEJ6Ltxjl3fDvC8hXPaOXVWveBsvhhUDcoC7c2x
OLjSS5t1+rBNwfDXRglFA5H5OlLZto+kiGyeXVtYKDv3GYMpgIUZInKl999T
9xJgDmhaz7E56kbC4IUYBTx7oZLDPFVsEk3iChisS2GyLyBueVg/mcE2u8Cl
u+MiAbf7lPcXp3VlXDGk6sVl6JjHG25nW1FwcWqHArBOsxl48dqAEe1TLI4P
WhDP8fYNkv3hnn5krL/O+sEO3VZDOMgpnjIJ65RsEP8ZCW5bvIT/E53KbSBh
ecncuilff7vB8l5l6KWFvse/vmczMtEWfAadaEAdrbXpkocGSEVIc8R2eqXg
oDbjw+dDwCC87Rh2O86qP6w0WW0d0aSDKmi8mIvaW5t4ucFJUr7mqT6dZ9+J
qe+6M9+jTId5caFXjfdhQmwOcuwV+b8uFD2I8TuAYLePxBfCy9eq38RcbpCJ
/zlYlmRIGCrrzcfFtTtUFv0YOyTONT0tnhemH3WduNXGfrF8QmH1YIhTFeK9
6kBRq+jcmyQTJzFwzBvsg1URjibNC6HAg4SuEsbXLtzkTKv/A1PN5YRAezAL
TjiOBDDlUpkORIHIuJ+NVkLyX0lSXYFrBLYT42PKgZj+yl9scN/WdGnpJ0KU
SYHwyDRcez/VzYDK1di+ZNO6k/IN8LdzONADaLe1DuwYaEZyeJJkku07pLQ9
V/9nGmfM2VkB8DPTJyhzZRiloeSZBurp1Q/PQLfdNRtuTvRXWl/WSHKEdszX
ZZ7aHGxnRzdUfCVkzTkFx6mmuo9CkNeWL1FuM4V2ztqGIMRiPjPucYypJ4Nu
pQ0fzErWAhKEa1xFZ/HICTumEZipma07yhpbRDRcDHS7DoR7aDBdzTinXQ2z
hFDcn8/u83betoLf2N77hTRJe3zc9xXYjd0nMtgNKYq8AGSw083ELeRgMtHC
pQi5F/8+Pk3ikPBJnG92nletoshq1+4fpJnxmXxRQfJqERNjVumOG8mK56UL
Yay216SnjVJBMaH2vTAM3rVczXy+zIp2oNRFLdLLUZknPgh0/3sFfrV4gGHc
V4Cm/wEb6SwhCu3DXKol4ja2vYckOutb3a2uRbCHqROh4m9AK9+YrSoNfZMh
M1dXufG9a98TbZMaWlNDszKVLVwPTfIlC6ygaWNXQg1FCDXF8ItHtZzE+BDM
klXSzwP0Nsomo91Jj38BopYsmE/yudxjZpOyJc+oOJIRjcziPhnpLMQBlFFC
rFBaLRwpjek1d7IaAiDriGLDUvYU+LrzJ0LFQm2PNX5Z9qTHt2yi7kCZQHpU
vSJ6Vkl2m/4XdVUPgnGQRGCLAsKZVAMhZVaV/YVgHY6HvJAiBQbFXgjP6Q29
Yw7GxF1klmPBTzOocT1KJSIcL1f14mLWz2+zo+zV3HYy2MynnM4FFBecGOGH
kN/bUjrWAdDMP+7fwtMhN6Tisp9KHvfjTtXJZJM1yzg/id2707/doseotoV0
bMgI7r6swcKufzdmRN91I4QOpi/hg+bkcD3jcCOO8PMzkHIeOjBBGtW3q254
/pcYpzNkQ3n1/Q0/Jc8oNQOHfgQQT3/WCiuDepBzwSyPfvuc+fhfS3sCPehV
3Kr3ZZKIxjZgVw1oGYLB4BEVOBcQiG/nDcOSNoI82dRGGMq92R/y5l9RFKB7
MKDE2oFt9+nWGD6xEFze67E7C3YVM+o8pxpQATuzgN+dPS/PntFZC28Y/ucl
bKJtqR8j0L/2uGVaDOCsklidCeFZhrsTZ/PCoN5F50ekTK9wopmrZmAxJxNR
HlYAFxp0wfv0Hjqzn78mb/IstngzkppNqaw1EpfrjnwnBSPoqnK2/kzeDDdb
LY8y2IjgEpNFxC1Ckjx34/KtdZMSKHYbDPGKydqxr+jcaBIMUTy16wwWxI2s
V4aVDrrCPqiIKQpb9YmO9tpLJiuhQxPsYl1J2zZFGhdY9en7+UuRYvxL5Uxc
iq+TMnTUmLg/gIkQ8C5nfXznv5a+bjOyJQWDqAMFIyClnHQvQypqmgEn3tgX
RJsDbOvvPsD10h0Iw46YQO0sUAR6lXDbVKu98cY0rsqnAtnJsYMqq2byyBr+
3TYpMn+z+zJIkqoHixOYU1MOUub+G6dxUZmqUGF8mlH1CCAkCm4mBHgkN+mk
s1w4MI/2G2ORfjOboT6aeE6jQ0lChbju+F8lTMIEKRoiaPYfwqjGYe/JadnI
a4bFf3cpg/ydQ6OqxeM4gU8GYP4iGSWzHkCkfjiUYsdZmiGEhI8HGq/EaAOA
P+UyV3Od1iP6au2ZDPPzmjx9t3XVfFe8PMGU1Iix0OQfR5Hsn91ZT0izF7qT
1BoCHHT8FcM9R+uCal4XSVr/L2gHe1zoZUgadlB69rM7TV4W+tWDbsTLL1BQ
Z8kQgTcaktknJCqu2ujky3gE7whfkP9WNS7VXc3g2n0ip24AoJMoQgqRyJEp
PUbnBNhyxuxB6GusoLniaJKSEaE0gfUuWxcCrIPZUN8TmJ5/5h3woib3PJ2X
2mD5Fi76FZgsdVR6dgyWix3VAgBBRFlaUQN+cQ4eKl93OjxKZ4u4pATnknk3
FKhnfz7O6cZEjGalkfg4ht0iALss5kPLfZw84yME0yPhTyBCTdOtF4Oe79Eg
2tM03uBOlZh57Esf+v4NEMFcGbaTJNmlns/Yu6csF7XanfpyWiG2fJlgB61f
1HrA70Zxi254sYMmpsq3jTLBAP7DNglxK19f5Nd8W6HIsRfGoEEOVqQNPAIl
u4SPpTkVlNBzhUb9O4PHmasRjqPtfoOzPG5HZf3XZPCCqvSuExofooOTG7ap
l4Qoudfk/63ytdoV2J09DgG9TataZ7AA6VU+3nJ9D0B+FrHROlzwcEvU0g+P
8/Zyhqvs3SS1Bi8bsrUFiKplMtPdZ2iG06FH5AiDnHy7Xmf6rAAHsIadC5lj
zqmx6Oeag96pBVGgpTsykWFsKN6D67QFrTHJDRIBH34vooRUjYh/XvnH3Q7Z
GZux6pmJFR1GRshtVCKO1mlpuMnU/huESAWnXvlN492Sb2R+9XuiREDpU5rx
xxasx6soxNQYsg+KYcJurjbB6AzKZY8Tdt4loEJCBC7EjRIdqxAsuselSrb1
Vg+i33Pl4Ydn186RoMSHdYPyBn6cA235vxt4IvvjRTw0q+llQdAueRu+uJHc
YsiJG6g3rPKAnSnrRWBKO4uUdcdHZ+9v5uuEie64T2r/OC+OUu+KCrLE6DNB
Z+pWwBwLRJ7jAM+Wqk4Gs/ZeUsm5y1XyATv/jwYPPD5V2RIYO+hug3C2BAEP
GpNN3reaNsV2NBG0qA89aERmOwmmcPq9fZA9VbuQRdDgSv7/0bL+hBxZ4HoJ
rFKk9YmdTBT2ZzULGwV5zRwbFZsUT2BHoSEsFied7fDwrlf1h7YJ3PFh+4o/
SQwhyLH/+cD11mNBEFLxgJbiZSPHo7DjJV/R8FnipY/nKMxsEJU+M2iN5A0v
RRG19OityMuk/foM5fpZa0Kf355EVVPOP/WfWE0OaME8E88Ta+PY7RDVYr/W
VzT38IlVQByMxqfeQw674dRAifSGzAkToMzTVcMJgD/etKqyhZeTFlTxWl0b
/DuiMb3Y2TJe1mNv9DZKubXTgO9HtuhORMaaSKKNyKEqF8CAR5yKs6F1cyRj
5S0op1jI3XFuUOTvI8jhY2t9XaUMCG/cfZdwRZ3Iz16VpChY1T6um3YA8tNB
GK3AnF76FEI+uJh+vhIcpNty9hR12IWgNsQkqeMEYBs9NIDrRJ1o5KEy8XJy
EwLnQEodrbzh8IGoCps2QHXzwBEhChp6cqHVX73RlL776IsXQCoFWJ9qWdfc
AfHUIjC8a6CEjq1Dq6RuoDF56vIrghdLeN4EpiLgYt944J0/cSL210BBjtbl
TT0349lPFtUeG468ToLVnOnKhGnNc1pNRtFvBAL+4w9T/QE++AFYrN9a4Eas
wjG1xHbU2etYM5NaWVFW0DFpFcNpqVM4L+oONfy0lMq8IlxqQ4kj9NA/Oqia
LVyTtYfLa3rHoDPahNtU3B1keXIxtFPOqka8ypYu/JHanXPxDNRN4FypyB0T
i7hVgaQr9fWuAjeSgNc4swhaM4jrTlV4KpUUQuLXASdrsJBFei7Xl7c7MbmT
f1ZkwUn78frKYRRHWrOJHWjWVlvLDEUz/FbYC0n5EAXZC6t2nSlaXipMTMbU
KQhB/ksq6BBT53JCAmxBJHEgM1GHVyjK7gwZp9dd6KXY2ZaKBNSJjCJSCiTB
W1PlJ2OjuCAVIkLcdvLTc175pjrt9PTOUs9H2KljadR5JeJEFaLFWrEXfA33
FquKLwhlinOzZkhrESB9Gz4TnFiHVljQd2ZMCcMhC3W85RuckQtMccw43frW
eImt+k9rI6NE0bDDmrXsvgkgS83YEVW6XcxftevdF109CMtehb4a1kzw0qt7
aKqbiJ0SbaA/auJ6O4CmKvImgbLV2g5Jlf05hckdxShVuPg2sYWbOEJl3OEv
SWLYDNrssGkTdgIpmZBZLf9HdFXlSp6XUzdgCsn4dZGiKwFAIyb1Lg4suPSE
s3hktwRQlXnoGFwPKgFdxtHJdEaXvQALFaPfOneAEu3J4pgmfqjDVBswnKxp
HZIn57zzC3eJ5IEsT2SzjQ2+zNKx75ulhiEtgcnCAZgF+dyepP/B7pLOb512
SkaGfqDFySLKAPyf6JUfd/Ywh7lsOlQu28iAEb4PlPQMt8UkkBC3YEYJLvnE
UZfnzBlXvjR+UHoBE+4HQth2ep+AtTzyPu1SbAseWssSonq76HfmViZJJ1VJ
pJfZMG1bLgOG10KkUQxCzdf6UwsopypACbvqTRdQAGiY9H83G1I8XhF+R0oZ
TyHruE/g4DFemXafbHJoYW4+MECxGSkDjU0WDyGlKIXalIuMnp7psBITXYiS
Z+MXWXyGdIxNjGdvnH2pGQ40osvlbVn1BL0WjGozoPjqBwL451afQXxHU/ER
pgoIZzllcgGCA9mhbf5P2UZAAerS2GGIYKiQSz8TN3i56L2PaWI46XLGhYYo
2zkHAzktJ3XavwmuPyStvHto6GPZ3lP7xTFvAWukoR8NP61B1lMIx6/6RDsZ
tTnf0kv5QBIUN3nyQJaLdpJk3UiI1nPM1oxkY2i/TMzTrZLKxWy8P3LFyY4E
JAXMr9Db8VPgKAvmZXekq9qopD82s2xFYRpr6pIZdn+pjpzAUoKyjvaOz/G5
6TEw+VUvFZhpTeAiHamJctvePeh/Eo7di4fn1S/0MeLgCQ7KfkNpA6vTrjME
nOrPUTQBAjII6hOS7rXtEXgFnbvP7ywiKK4Tq8kvna1qWQ6mO81AlBx95K7u
vU8GzztnA7kcl9BfN1gnetyN+MD+K18h7xG8M99hcpbqrJX1UlI4stC2cuRw
2EAZgisgjDs/Xt0LBQR5H3vb4autSO8d93J7Ujlh+jXX8M9neN8llWM+sOcE
wxSsi/lg/TEFuvzSj0rA/58iU8/ZUUNYAta4hh5f/ekx2YGGdmpQmePUGu1f
VeJT6BOCYs75lQr0Z/ODQ3s1PHYsA/MjSIXpbsDm+0dQNd9sb5jQ24mMnWwA
dJF0cCCIYSsRq0C4UczrMr2pf9/ko/mWYNbLYtkotQIKmgMGfsvwTwnvnQ4p
APV1AbIZl3sppFpKM/DmcAf0kq6VSb27r5bqFz7QKbX/3+Z52ZiRPhgFoTGD
p0QqlbZiwuUeU3W0fpExUrBB88XXpaBOGGu1c3M+ZApclMwoBW0uxuWi9vyl
Va3fNEH6KZggPYJ3aYPVpq3ScdB44ZsyAnYofK2zgg9Hy1GX/8ANyfMhsJwO
q6pcOjLo3RZXpAwr52VGza9pVaEOZb9CplAzJR3kHflHuZ1hrog6poGi0oQs
XMmTtcNu/ADnv26Wii5T3Y19jY23eraDKU47b3rgX7f+EcrGUlAIS79sSxJv
ejWjAZKnDhn3x8j7ArhrHpNgqobtKPRE1JN9SA+bXqoTPZew+yQ+1FlXSe8Y
Qcxa0ORhxpiB81jNUSIidR+UFgXdo8YST2TZDtW/bFTbqSfyTSb85hpI7YmI
HUz14aYFlaUUNjjpumCyTPC06nAnV0ml+ovN9zizhMUh85GfJpp6F0PGnsSd
t1+8PLBkp39GIU9D4yrTgK5Iu6/884MQ/dt7+l5GqnONps+4OslSQBg6bUL/
GrEzpQLtURRKkXfUcuCsU1YxAdLuxdj0yhKULbVSFSTR/Im6DZw3AJZsqTnV
EEDi0vGzt2bgqOpVdj2Ajpcz9dLAEodIz0e10y4OseIelX3jELo1oTfdyIkH
cNOegwOBDpEmO8jiV5QkzRSJf8CfNAWXWbq2MiInaPSClrc/7RORiAcSlu7l
16Q9qDMQYIkXlLMeg6LIMutL74CmPRuEFStN7NsBLhY7JU4/LmFuIS5+TwAx
GIahw3hYxp8su7Me+g48y1jPVSmnDUP3kppo9EqhZJyhhrhTzObbau6IvDti
5mWA9PXI1J6GybP9I846ihAH/gmeB8emlN/QaswIgcSQ6cFiZZtbUw/OYIB8
Q37t1oSTQFwRmKcxMqEUZ+YYbSeRGloUkxTHwunIqEtx+5AmEklTNBAoRHtp
pF/k/Lg7IRG6Os9OccIx3z3p+G8UsJhSCVES9vol46P8MpWLrgmHsIlL+aoo
iQhz8o2a/4xvoNRpyTba3o32j+uMt55ZdeF0LFLU80FwmT5X5rpOPsSkUfgD
UVjW0ys7WAOqTJsLbGxhOplaz0rlnrcFfHgrahCttzsiIxMkQmTTWXfoy+nc
NHD2ODbBIubz2hqFS6x+GXKtHQnRz+gRTBZrV+WsXlrfDyNam5iRtGRczUUP
08+FRD7PH1Tdfoixs95Sw7szjNQEeySZj29VDL5jSko0ouhDa7ytr0ePyLnr
bdWfzrdaeZpHGQAaJJbWPAHhyDyZvNxohqr//SZXqrSwza0xWMADwyJfZ0HZ
OrQsF1/ZmHTRZXro95qMf+e5DYRIq1SZ0cwNGNFnhITaYDAauuV7bdGREAu+
Sybjd3/3pmD2Am+VO5KuJw9E/aZflxYCjUMscfrazyBzbJNKPPWjP31jbJ8f
CPcAJPGxtejLOO11o7VFIEr56P+ylPBQOZ3nELbn27ZZZh5q1FBdvFpsJ+Rt
8JV4lu8WWkiT5at3RYooK7pqLQdfpjKiy3c7WDdaCbLrTk08fDBuK9taNn//
2yK6K4vON9VwLQud/Z0+S/YrtNZk/xZ322bS5//A/34XFlILnFTBOGF5TwS8
VxJk5IyREYDRrM/OGGpVu4CybxySSq22R7espwGRAMNmO6ifuT11+So2DTJh
AtLszinF27DhSeQ54D0B+aV/bR6EOgTjLGpPbyDfV1IMsvUiqjW0LqAXOEWh
OY7v9M9Zm21y6doaxKQXWfe4kwZhxZie7PRrgoF52Oa1MQo6B1y3nkJMNr9u
k0juXzxXVGOnxRlQr2V0qmZsa+eyhweRG5q+L6ccLTPv0HmUD7WY2M9PhtSr
+AswB4HrS1Usoq4B3NzXeXcICE7mhleJNu5o8k3w44SQvQYuyzFZyDyvFjIu
8WUM6QzJnBIBleGWgVXNmFoH5sFQsuwQQqGEwf6SZNkPSedMzbqdqS92haQ7
iq/ETWH8hPug8LT73sxgRYckcw6IAa4Z2To2WEHdbZNky8pNPN98NFrDxIZM
Tg72cm8hJfnQt37jigeSmr8kxcsOHR4irKog04+VZK0a8TvM1SHJCn9NAHu5
acdLXKaoNoDXJtDu4RT4YaoEGYMYI95Jzj3e2/trsctZ5i+4e1WSaA2sjID4
kp1BzsMdz4622Yo/Ddmp5TMwUxTXp+rVW8Io42bB1LOvdX3AvdZ4zuxlYJAi
SHlbgT3e3h8GS3ghRTjfx1UM9yZfy0I5jm/C56+BMPSL00QpOoNUvYmTb3gH
+sm3u9/pF9r8NpYcrosVdeFTnO6Y0t19AFJs83DUMKdirAAyn0zggu9iMICk
NtsD49bylLFkROdiZTLURBReWsZg8J5ZqTCDfQjsJQZWkV26F89e5lz0mzoi
jT2x5pyMmfoso0S/n+xKqDhNHnWJRoX6kFt5+sdR0VON6P/h6H+dEG6HoQeL
PdaI53gJ3JmAzQkhFLpOiahhcAeS9yoV3ihP+blxDBrY/0QwJJpS7gJpzNvA
gHc8s1nkiTuKdVaVNLEaR8geOpWytvs7PQFINOOWFVupSYEZREYw2VnrkYc3
QRpT4QmJt5zLzAgdOGvJ40teLVxyffPeuREc/dAAR/5mIiNtOBO1CifHymPG
UuCvSn9Mh7HJsRbJ6pJrDQWtZeJ1IMONQTKyw7LWFXkLrg4TvLgereG4ndn4
xjJTcphWN/uVp2GhPySyAabgeyS9+JeoAvclvdTDRe/pzgQ4oDZS0so93/us
T8AMZM4PDp3dXIdBaIKXt0LKNFOYNEm5t6z8rRwHei3hBbmqUahjhgZkoAQj
ngvQFa9bbwqSyV+ytUxz9SgzDJxK9UN3BLlXmQGZOyN5vzEDsCptTzbF+Q2x
M9t5ZHc437l8QHeIS7G4o7AtTGxuS4PyRFoxbuj6p0b+zZRE15uBRcOtL5Ix
aEJdLuZJQb7Oe4OOLDN3JxsbQYfziJROIE4wOE/p4VRD1F6+z65A3SpWDeNp
xqv2pf4moWX6B3VG+m9g6s1H0HanlmxlgR4krbJvMPjr9E6zcmeiEwrYZoUX
b96+YulHir0J2zqU56ywGQ5HsfghQA+4L/RPlfn29ZKKNvmGKv33Xk+6DQJ8
OTkm1XUepKrQ2mczd3GhFwUiSXwMn2AyZyAHDAAGSsdgpMmJGwR6ZkOdGnqJ
xfscrVZQYaaUVAsA/sXxnJYo/g8kZXehNngzCWQui0fXhTew8414EAvfTQXG
FedGXDr3rVNtappy0NYJvF1NuiG3DeBBVyq4Du960jesWrh2yAplJq5epPoT
XUdbTRt3Lja73giZW3yj18ZrFgWry40fQap1qEF6noJkGD22kVl5YOue8uZ4
7CIZX9y1wQhwOGa7Rf1ydqRPsxAkxbBe5LwzIsIzXyGP2iQ0dui0HMHF7Cpc
hfCC1NAAHCKBjzoNHOEvHp0OkwWvo26ZK9BZy/f1BaZUhf5IuEP8S3dGlT+E
jjSrSEH1k/pjZ/GNFgUo5TzXAgvQY0+mZ94z8IcyVOy5mUemXLE0lHC2U+as
WmT3abdG4/JG17qpBczS0MrxveVPv8F8X3uXlxzpMy/n1szVQnJqz1hWmii9
1MNWAKCRMuGOBgc6CWWyFk6YtbQU0tvPjxYavqALeMMBHufmPr/wBX9ruPrN
w3tw8ic1bD0H4bNQ5GWFg8zWAysOalmz+jkGbGXdQmJ8Mb0OeI1jGnLnzJrh
mt6dRackdFVi3Lt57W1gUWlPNDikWxQi11iiKzisoWJVnk3ncWdV0FqSHjQV
msIqU7QCsLBLrHqIfbc8O6NvmdVIji788bETzal/aPqEKULxLTAGGi7KSTnt
qgBz+rPFPz7gTKYSTSyXQ8/bmLBmfSXE1pVwWsPvxLxnQciYqbVC/GDN4pYv
3j7Bt1Gc9ZsZjbjq7K7P6zhq6gjzMCePKfMyx4fLwpwz5l315Qi2WP/S9MbC
JXHkcSPZQ+sIEnCbDXC1bNFn9xCHp7/g9rmHedQPvS++9frjO+gtLbWNmuyB
SV60BGt720DDXazJntv2gf0R7bKhPQ9YOjgYc8SLRbSEnfDvpqoe/M5lhLPX
GRFM1I4Xd/8L4AzAI/Anx96kwW0t7vzdzo0u9upbWtcNWNwLqLzoddetlWXO
RSJ+yDpHWdWFfmLC7JNh/+8n6V5GO5e6OkFK+iLbdxWIuI+iMoruZKUhNddf
WWhptVR/nyE3im2Qfyya7Bewk73SNie4uvSnD4tZjkbh9ouQYMrZFWt28DLt
gH2cTy0hqvn8tWcMzNFyMkjKSuCRj1RhtT3yYObX+qdVklpZ/lu3FqKmuoAt
BVr8MK15TEBC/p7ZRrCGz5yWiLHbHwyAZqZC2uA3P9w+ZaLEH3I6mvuaSlA+
qdKqHTgiwRhS3OvYnRBtMmHUc8aLG2kc6igAiYiaN33OMO5OOg7uJ9PTWe2W
0FirdmLkh7AkH3PEuu22mjP4Roev0oByRyCRT+fTqSzGpFqxhPVf0iXrudP6
nDD1r6H7KtljwGens83LqbwNZ69M470gcANxYVN2LfCemKCpvqgrYzvn/VO2
nJJMQTH7V36b+faXxJvDS+5szCUxf/zE2A/KZkxgVPZls4A2ESG180pAtidp
84aQEGVx2qw7WB4bWEElxJ6SkNuRNbsvurR+sVJLsJeLhromRGVO6QxfAWMd
zj5H5axvXDzKmraKlJWtQJ7FCDnquGt4Mf6WJx/gpSX3QUfvLkqm7OwujmqG
UiNASaHvLcjEgdOKA+jrwovGOQDYSfcXS7DmJVRcXGz+UUQ4GXIBn8QxUHkT
cV5JiUfNfuG70kkamQofJ77I96rzY1tlb++ww3ZnC4W5tqPwRg+87xtAFMSp
4yXxN7NAfoHzxlylo3nMMpoV1hDG6aM4Gg7moBX0Ug26reBJmar6I8VpvDum
w/iUi001sGjx53s5llzUp/YqgviNgRdEjRuBD2e2Z8Yzl0v+B1ka+oW4thGs
u7XxUaqInUK81pqqx+P09YtidPlAQvB/S9WL66dAmFvhXRDpWvRV3NhADS82
tMjr1H3iKYvbAMWnv8bA6g9jLxwnhLQKPvRwScAF3z3MS9E32k1cg2g1amVw
r2T7HCR1hL5LIAMJSPGWRolXxDvP2YEgZwLYUsH6JRvn1EmpwwoYlG3+Is25
mwPjl6nbysz4EalOYggqtosTkwp/KGnMqlXNb5j6rNSkPL6bSZRs4t38Dy7R
iuBimLJg9wnDr8voH2mctygDxc6bdneRn4RP9ZIt9vGKX2MhI/1tzB9jM2Nv
zzXkQ7rxi7knUy87olScboczu1QESnRyMgdzzxCKPsZGLllf3LnMobFUNjdV
F930ngoijQql8C52wi68320J22RxJJz7qS9Wx2ReJT33JHi2a6JkpzUw0hov
6fR3hZP5qsnQ7OHlrjvkvis+7OCAgtFt8l3DFRJpdLyXDkHmEPGUpy6P3Bkg
PZgSmz1T5NoFLVhRUwwaQPO/JdMr0dQnB3TIqziBw5eDKKIV3228jwa4ByYt
dTL1lZMZN4STRtajqkxi0Fng9FZkAG+jun7FXaQ8QEpqQdA0hOLgzppRjnik
QtHt/FHAw/htfVYtlFeTugOVfD6UtrsB/No/8RDhiqfWbR867mRasFrEXtkn
6OfBMYoXhDdvJ5qv8FqrOTEtLVk++ciJJ3W2Zw+3cOCkXVay/CGjI4Bsmg2k
a5DNdZKCRa81qkLzciG45gsSMqbAL8/5mPiC2RirY9YdUNC1fv04CwlEy0ps
79XOvrZysiOJEogfQZrXmoM/4h9bsoY1G1jl+8a3eh3UwLtN8P5cVHMs7za3
dP7k78Q7cGZmLrG4d8s9RFYttXjJefo+3KZBhOKCyDOgFltMrUAi8KTmQ11r
2+UHgNvaIQTFAp3x3jaR4fsGx3py4Bks0/C85vS3bLkQEb3NFEbWKSX5Jx3h
/UxDyCFo3GvEFriIWuF8oL6wSzrm2B2qB9wyvlGaz9/WB8On3/9YjNIqqnjO
AHCPMTgdbHp23m2k3CVRE5nEmdqvIMpIqMy+F2fM6n1W4bRPTHdnIPWHfcQt
uidDYFo4fKXstdDtq7TFZPuqqcWUFCd3LybhjjMOWAXMMdCa5PiGJkn4rZG0
4UZ8uUVTxhcMCi6S6Q/UmFv6DDOXXFcJUIji8SnuVYCUcjYjwDPrYCcTgreU
W1wvPxrIZ6aaVq4PgLeU0yJjFDv/cj3GnRZzGww9OuaDGkAchwwDC4UcnXCC
NMrI1sQtY5lTkdXBVT0rnJeYGBnNTwKDV0kTn2gmWKy6LUPiAI52Zi51M1Ez
NFq3SFIoGN4ntqHbHQF485IxNz82lG7Lbn9veNW3scZhxGdhy6TxiRJqF+bF
2rZCZ01oudqB5UoN09FJ+8d8rR5u87P81SDByGk9coXcHw/g38a0KL3sjru7
TdwbOY1fmkxTXtR8H6++NmomgsokyetSTfU+dMnPX6unHtilVnrcxDT6w9g9
Q8Iz2VbhOiB1dY/MaWieYIyG1pJK5dRoErsI4W/8o/7L2icOZVdhMkOAivL9
oDkqDwcE04jYPeQg/Unyzbqm0Dg9Yb/xwNH44QEivKYYbZXHHNa5LFLwhv7N
+XKFVnikSBcvmGDod/bYRG/9w+WsO665Xwk8jndJo0UTQ3dqkxDdbOxj02S0
qDb1DDxj7CuEHf3A7CPdbyGDXTs0rHA9ONKU+mdn2qKJd9heFfpLG5+VXEI8
Rn/Z5YDxbURfom08FgVtvMXgkkZPCL0vCv9hXPWJkZjCwe48PZMj8FvBTK2X
4qj/2oSEZbD/VQSD3VchjOybvsP94L5LxZpsUSzUN4YeVuzuNN2g8RMSMw5+
4I3tCy+1X/GAjNezeD/cZa3uHITsTQMmrE8VJc7Jugt8lz7YbNy6dgCkvXGw
0w7215qF3Ecv0xvGfufKY2VtN3BR+bqgEMGH4mOK1SXTLIcpQyI0vwtazKRH
wnu4OiKeD5r7B78cSvpx/IE0VNHyclvMFM4rAMLmCCYRcq2JGyd4d3BgM5BF
6pC74RsfFLFNuau8J7tWlhjDrOBvA8HmwXUQH1pMzlybamlmyejTK3leMIcr
UuVh6bT/esaviYd4faNE1R4XE3BxuH1OMbTZdVRWXoNrom1nQVoTxHqeQKRG
A7lmryli9KWoi15wuIvwNa3oI/ymzwRlQxqmSoHCFPfozve5P8wi5tCJtUvN
iloFsQU53hEundX6F7HBtN3xmxVR69CPO4OJE+BTHEgdthILuGOcUkxtntlr
TNvZrUuhPQQOYkyCmocQHs+v/xe+WNUMY9zhh82ogbInehlOAUIHp8+YqlCf
TNQWzEYXdCqxwmiIfxpuAvTXmfPocpO9J19mfaBHyBHA7ec6b4okrhYi2Ae8
W6/4X2izwf4/QwN26GvygyqF6WTbjHGvjjPGrcfwZN9+a1teUBK2ObAidGEs
3OdSQ/rIvO91a02FEFYBUn6nUwWkuCWJ2xplrioZS4KyPXZzc2GgMb/d+Hdu
XJN5YdZKs7D7FT8h9PSHjxplxV1wQVFIE+OxTBC+W6NYZ8prOZI4pC9qsXPC
03G9o8nmVMW5Bshi1qaUToagy9W3rPTILRafDdblg3z0E+7t7jp/meVfVaKA
OQElogsGQ4qCuyQylgdHm4BgjeUoaru6SyIfL/xyYSR4jUsNdK/wnB6GjTSW
iCbR5ioMa4MTvp8+5cZF07V1h0yhtjNUkJNeslr7dhf1b2RvIBLO0z/b0YVC
cbILdga5fvpsNJH+5JQzHH6dQovGUU1MBdqfNwhMWDgiTBkHL5Pu4GowKM/n
AGkebJMMbTipitHRhyRxVwGdX6Ur5vODbBS9NMDdSBF80dhaUF1FsBlYpyth
4WaHv1QR285v2yifqbX7WyY22yNW+C8kRokqjT6L/vPGqw4+gXXl9QbYKFll
AaZE7yimLF099beTSJMFZH8QPJJB064geRGxMxTqEAOIXURUhhfqE3GyHTjJ
vrWmWOq8ZNBiT2TKgmRFxlIYW1VFrOggfEHfnUmn/fiu2nu9vT4a+KREAMfB
k+Bry7VfEumxty8GfqGs1y0b4x3LHreLSTqNJEtkKs/PXRUFgPnqAbXfVc54
HlVd1lpV6Zdc611vaQcxfCmea090f29dJ7zShok5Zx5GE2156pIwfM+r93/U
W/ep6LliXwdd6ITggJsL5ClS02AjCSsUV7wIkFU/QC0gXtYlRdBROauK36YC
i+Gg/FuKGEd/uZ5SF4h4LFogfk8l5VcCeuEyEVKPmaQOdhhvGjupL3/uv26E
EF8iuEfmaDrpFtYmBBJA1zWXaRAYfvUVVU7uanKjEAavQ+SOIFrZg7kJV9eM
Fg5ibO4iWUIY+/omfZPIlhoY2JKZ9xXrV9Mbzss3bWvFvI/r8rEkN7qJEJe1
VCDg9FyqnH8CeM1k28p9CYGNDVrunVT94KLl1xdfkBwftA6iHQ3B13SvbosW
zB3mA5nfISyzj/4wHHiiqgrGezArP4JjD6GfpEeXtqRy/8H5/alUPewyrydH
el1McGUYRho/9PdDidaT/U1dHMnOcKbN7p0aVsh2Ebxo98DzqSOOy8BjACNu
9dJVRAB9SkaLl3ZvVj+Ju0MB8dFk65DAZQexWfxx4HIncsuCwhBxFHdrXoTU
UQbO0YgtfrcC/bFkjm3/pxT7HjZXOh3NINCS856d8Gey5tpFVpGS1ZIX23y7
yG+fXLrRZA56LcjTxpGgI9e+Gp38KTJHRGLGb682jPGY/TkfhO8lpRYMEuSi
f88DH5sOG6SfckBikwdDHxyC434NKE+kb4u4qGusfK6SEBNpMznw+lTCbqDj
WqOTvvb6DUacztnXOrrAx63+Ftruu5W3UxFoaq5lSF/dUD/TR/5LK+2+rGVt
WoH0YTuLGH6aguw2JcqYfFO+BOYIU0sDcOOigiLSj0NK527W2t5TTHt0C8hy
lnra/E+h7KR2Vhj1tbBGgL6QRXTdW8+AZ38KIdyp6MwVzH+I4UUKMTMuAVAR
wvv7muTDspG/qvuPi7JXAlPBsVle7TpRdm8WXoAapIGdMvYiXVRWhW8Z92IL
IM4NEH+DzJ9fbPe5xk3Zxzyhw7Wu8m+L0SRnLN+YfhN0uEY3KhLpxQjykU1E
rXwaxb2HzsmLQ3XvwsTa4p2CCzUHtSOP5KgrJWNhfvl2qyEeyErh7W0LfIbS
CpZpijWnyXIgRbNjN2hp2csXN/sBph7y73/9Qf5JOEYHxnBSbNwyCQVpC4mq
hWT2FcT+GW793Y45tmAYfEl/z7RgrfXewamDBYDuQ6NC4PIAct+vWyOQMNgz
JtCdRkJTnHK80rrjJhwRa/enxKN3+Hlexgk4W17zh8dhBH1tPw1b8NIm8jce
+R3V16ojNwg5LsCCjhD7eLcjvVXNEPCbVTLtwz67kB30LfwH+MjnQz5jyPf0
49YDA14m/eHS8fWvH/zYJN8UW//ata9878CUGI71CWYuJS/GdgEG/l76gy9Y
AID/nTg7PnIe0px0IGrLYDb0f2jo2ZAdjj4/L/+gWxhOIfxjCOWmVZC+oTfG
Yzirck1ABQ7YqejsG5eX8MH2wuDmE1cPdYSuglcf7VEfNHigAXke32jW+647
nykTckpBsgW8axt8zWPHNCW9yg1kKApzY5+omrB6l2+7qdr1CRlzbliqn8De
B84fKCheVkFqbO9Mo9qVGo+a4J0aWO3qtuLFLsMU6XEWn55abQcwhKeTFUdl
SJRo+BhVEa9HWnAm7vg5pNu0xkeAlFtUU+aXQc02M299/v98PT/QKEsVrtdC
TbWd32226kTiVO3+7qJW/6jEJVBNUvKohmZ5XlinGSAxFb+/5GKdBuQodHma
n17PcAE5AITivoGpvUiWyRX6Mf9/euyuYyPusioPldAjahTUAvXM9VLmhCdr
QR39vks1sR1cJGkc3JRwRfIuPywXqh/z991uq1EQyiDZ0cYg2fyjguCXeMce
XiCysydMqiVN5YOlKznHJSeH0HfZLcb5adm1QUbxu4jFs+RNuaGe7JUhZ7aJ
JTjOgCkZwR5SFg7j2nMsD+77fgvXlb+lcCelQWm7onVZhD9WBPRRzEqkwiIN
PPd+T2idiW8N3SNPTDORNUAtVnNUeI1hVzF7MW1cEbiXJHkV0vzndiVeE/FA
gAW9bCAwdZbYAUqw4fEy2qarFztunVCD+qr1rTi+KNpyTrWhWBubE7sCsL9f
JBN/lSfmHiDmaCmaMzp/Iq3y17/d7AXHP4ar2XKX5wviSwkjlY9GkAtIxjYm
ML0Y6kDX16N1RsIV0Rj4nPJRBc2koCy5Fq4ZDFQOP17jK5J6qqNsRPQbdZ+e
cgoyKUonL28e0cDLZMwt3zHNuX0/CIZ6V9S1j18Y/ZH/5mFuyKscmBUIIZXB
a7FQMI1Z3ECmFeaQ37lv/ftgcGq5j388swm8FtR06VEsSKW1NRrpxVzDCbMa
EY2EPumRZGjU7oR/0yJxfWwI6GL+vnfSwN+HjmKCjWSJSFjsiazi8GJL/s4O
u2ddgnI4CZgl6AUwQC7Fru5CZsdmwspZKDG4dO7a31/7j2mCI1i0s0dAuxiT
SJXzcn+zJoY9D2FjPxOZ9Nu3ZA3GeOkHTI8ONFz2R09/mHtG1rIOYtxzN4B6
DyiZsbJ8HK02LG4faiR2xkK91z+pGRR8YO2BrpOK3Msby7Er2zoIzH9U9LEZ
T7hmrGDAd07aoJ50LAU0dGRGf6yk09UTkk/ri7ZQLAXRaA2gPJA9nii4BlDB
6XxODhYLMdldcl8TbK3oXQ2A2Uf3s3ny0lWB/SUtU0dn8Oge3zVHE8bow75x
upCc39N9GkjfYwAPn6AMRsoMtqFYylZkq2wmAHYgkZhWJwgYeE84AEjPrs5R
Hs4JFcJ/szx4EitWvnDC+OnJKnKtPYb8DDgd49kFcVeE5HAw/r3vO6OBncou
7yziPj5mjUusvWlQmyALQUSXkVloIOyOuggAxeoXrEWUXfm1NKVfp1v9KSnw
sBUSKru1npqwmxzKH8E2qEL6wNPQlApBvo4zbyu5hPluIAelsYKtCfNjnlsu
n19MQmMPvnLH2zkBatVqfKamfc84M1iCCKsuBPgklYGeUNY8WJLYqaiBZ4u0
EsYxh6n241r5z7esiiLJ7pVRR5pcs2GL7PUQwBIP9V6qaTum/dNcix3hN/Sc
OIJ6shA1w2Xp2aBmFmsBgpvKf3GH5fx91QFm3LLVkUKVTqYdzRtbXURFxWfs
0wy4d44N3Sq0Ier6RVTegfq97xM+qhwBiKR/xqxQcgg/6fS/fSfd6HqpWmW7
k403UamV3GFWxHaiuNb20LCALRz9xsDu37igwhC9N5K6djTknxSuovVJD8Df
tYuCLjwd/ivo6Yh1jMSXwCouzjcQ7JQr6geexRwgKYepMvmAQ435k58QziRL
ku9CcZztB1TLAyJABqm1vwyHDp084fnp4UE/y805j92UXp00DINR2+W7qaZP
vSjqLn4pOjdjulTBvisNBKlEERYAsmwkLRXKW9oUSzm1SuHnikqSf5q34f6l
lTnQsQ5vwZ9vBNPvsKGBs9pSIvLFzJdRzIvOAHC3mIDvWwn3Vw4NDHnoaXQD
SmuW1m0gjmjbajNGBUTRbufQ0Qw4mz/ZLauJFHv+x1t0X5KoTtd7HlPj07L7
KyrA0uBVEcmVmqc2HfW/BMwr0kvrFXWQSXYMX7vdmFubqDm+8V16FVTkC71/
hoPWDHlwM85Sz+j0u10UbYePKcbjfvGdMGmFP53n22kJYIkLepGTwso5QqWA
m6anO0Y5iZaY44cVV++vy4o7KiAMUDIyKJOmtWyuBPUvgBFfkINc3AL6o1nk
a4G9RvSaaqOUlGK6W87BGKpJlWIYkzmWNjf0UJajKs5zhxiR2zOdyRbrCQkw
V7n1dw0imSgQAprRdr9HrqGukiyOaA8Cv5MLLOyby2Fm54I3q809dnuc2A/Q
ojmmymfmXvWiPxxhNqf+6yUQrMKAFjGuSzcEBeyaydHuDKpysklklYX9wL3h
QEo0ssP5u4WCcmQRD60JJXjKiDgr7eTCV2FLLlXcRi613dvtOF5vacg8GzrY
off5M9K0ClmLkrjCRsX/kPoRIzKKoGtbJXdDwfsABZ/0fRjs++LE57jX3eQs
YeLn/ewEthLDS/L7P6zuXLFhjJhIuMDIr0fsEQbPmoWQTTBZlfNSl2J4PcJo
b0txVm01Q70noRKKesPLfW4E5U3dsPiopa3FSaSNOjNerXs+uKOFZ/v3A9ur
vugTELRdHJtwAXHtf9wFKHfQ2N5ijy59KyRrrUMAou7B/BU5GFA76I0Z4Ylf
pUAXhovBYEoH3sXFxBw1DddF8akmNh4s8CgRkKE7SdIYfOzzTnTTJQN22UHP
nk2bNp1hwqgFsk267FbR3981+HvGTVrzyjbzWiKIIct3JTjKvXpad+JHd6Vc
AWAXbzGKceslPFpKIXavs0plVX2IyBlYB7HTyZjqxoD7cArnd+O3zMNWu2zM
OP5ByCQnVBpaCKEvab7yeToXrb1fec+1teAru3FYc36RQ/9FpYRq1RuYnqqa
rt5Ezruh6R8KQ3/KWtsZCmyPVnIbTkyGyWGLOcrL1qoA3+wplcfVWgLFp1+g
qJHPjUUc2QV3AGq1ZlQllCDOPFfnUF8Oinn3RhEywsUuECApfaZmQNt4lg2P
gkEyED6MSbF4N6SurZqEQ50/4gzygV1hyK1Y0/b99lyagj4WqkujQArSccP0
CJ0Q2oSKtDcMoMqpDDDIion9dX6FO41xbMftqZjiOz2E4nMIjsJMiA0jdxEK
prgyuvYT+7Bhz7uEfMnn92JukbI77/7rexcXhc7kV7aw6qlxVJE+U2SeVYnA
8ddYmKOa4aIXo3FyGNWxG2vbZOoM108yBOteNQf2JWp4GjJTM0sNJZCcv+6V
ncMFdMtxs6SXee67N7RemiSlDWBIlrDkGn7JF5pt/4LtyAduywUKcYxW13pn
1/D1ztHBl9J3noEd6g9kdxm9U6yPVWPOW5MM6ygBZrr91CdaGHDMFW7FGn3J
Q83XGdBpBuIDT/tEhqa40CnqZnlxdRcrg1/RF5TXoF+7xESvj4NpZovS0cf4
vfh8FB1Ef2WV90Mr4IYYVae4KntATmdhIOAUnV0Z8/cjCl5pVwLaKsGwm4sN
uYI6f8slHf8gGw1X4MXPQ6p5UG6tupy1wDpj59T6yH7gEzCKq+h6dODIfE9z
HXxEAbLyy3ahulrl4Yn+Sa5av+pHrmGEa/KItmdnxZ0fMn0whdOUI3KMRb3v
TinDUmLr7krVxYFtG4Q/9P9Vg3VYje208UjOzn+bMUsqKGfocHl4LB2rjeMi
3p1IuCJI2mTe/5bJvdyuqWXxUsDxzIexOv8LyBCHni0DlnLL5E/U5a9c3tqq
xUkgqfo6OWxh4L2rKJE7LTCEvW2KQuamYSdkBQ+JkRAqdLwkvFX+crXfDYE/
W0e1yJNIKsXBphWC5kSDXLNAqlLuw1KSR2tYgT7QqdQgKg1xoCflCFpsDzhc
5/AHDyPb+lW4ELoc2V0HMaGZFRS6NAlu0bcf2jU6uvYzLKuMAEIr4MAgmN7y
trnbj+BvR7RvTpCuzcCUsCLWsZW4AS2btKFBLULXvLk5dki42YqxOYQ5HGcO
G0I05vG5HfLTWvftV5L+kZxjfewXerFzL/nu7qrpq+mlldwsb6dZDWzfYQZn
Hze6hF0/phAC4KABRskQPT23YzBxlXeJys5Yt1FV4y3TKTo7p1Ax62jLBMyp
AOLOXkK9tsmId6BaiMPGPsZHg5eDMJQGnp19QA1y5dt9Mat0MMLrggswws61
eZOe5HbFKou5+1wnvYNKql1enOEzt9Lk02dxhC5urnzRtIXgExMYhroSZYiP
Pqo2mOetYfXC0X5GrbS1J993A4qWx+ufX587dP3Dan/BF30Vc0XFOEdp+JUu
rA64a5rOVIFD98Tp5GkRf3bdjeszUUFZSequgl5o/jK+csSYVGfXGgk8QO6e
R/+UYfIYL3ymv3JEsEtuxPj1WKfOrLgUj2RlrnAO+quv3OkZz89ncC5JLJ/M
bpOSgFRlOGKq0vsBot3zKPFoVFi0aer/CtKPOblf5qtuuLHs05gAaoLawEG+
bDOwtTMa14Ra9c1jhGa1MfrhiwaUyUm52tvB+3sAQybUTT9uORyrxpGemr6Z
fVtyPw5tsTuwlnbAE5dlZraxM6StOR36S+160mUpWbpJiQNUACBbC41LP0mD
4G8ZCzSLw3vNT/aDOpyMy0witBCdDJacwECCzvX0xcBTVa1rC40o1WHSxxDG
o8/3UWys+/XGeAcgDwQad8y+MYjbk6e+CkIzyQgLHT6TrAnvqIEiaMHhy1q+
Q775rzW70vXkxGstum5C0dU3c+ciihi/mirmRryQjQhg9n9IerveyRp6KOVx
cU3lEcqjO8mEKBU5ToWvuDnWby1j0v0Iw/+bkZzwvqkBxP58eWZ+ytNwMM1S
tf2vBFHpYy4zrnF2+Wn9SwRUOcchRd7LdEkya95k+Lz4gNd9qYyOXH3JYEiY
WVwose/xPIQ/zn+uzsz6F65hOcSaB9VPp9ti4w2OhaIVFuuLXym6kJqJcFEt
ShP/WDxCjpWnTj81/4gwUe35ZvwG2/lPm7dZrh/6CxgrHrtMxR/ekBUkXJ9l
fvQqgOkn+pTckqc/uFeHjhlL0sM0xfjIN1j26cIAChzhJLXebnXLTCsCnB/N
WUITY/7MogBHaCrNpLuLmsPEjmOPz6Ff0+xqeXsYh4GsI+pe5g74AC2Prwkf
WcaQdDXZKqweyDWUE6vSsGnl6iyd460Oye0GDEP8eEHJ0Lq+Tl0ZGBP6RFDV
NkJQI4n37A6sKG+wXuwMQlQxbFeI9kjivtE1y16zJjQ3pKNZzwBX2+6sW3Tq
peAMxzP8X8vKaTp2Me2HcR+yoqs919XixHOr3+Yk4kkiGl8MGG0fN4l0DpMt
QNcEwyBdPTP8go+7WbPG1vY68NEgSvYF1nq9L+ejg5eJrVX+OQfNNHhzKyLl
d5TDDpc/VVV8X6UEJbnBYRe4BLlSNCF9fiAsvY0Wok8tt1ioOKc5VIyJbd3j
aBWkMxDyQaOKXQVIrxu/Yy2IBL/ozDxogLYZrvct9GWzdoiVTcCeA5NHD9kM
izG5OpyMMbrHCtQAAN20D19Jy3R72r5Iapg79Sj1dRJap/XaA9nIJnvkMd43
bv3jGiUSzADJVjZ8jkY/drMc2EhpTNSVDxF4TksmHBgs0T6i50Dj1ObxWi3Z
X9AcjEfsceMrljCjzpdHwxY6K6byPSidiVg5pmj9BJm0WZExX+DhuWnkH3g9
jNJGDa6VoiWZyePXmcXeQ5uqlSbPreYOJqXRtZO26qNWSuZTQNXeYctn+m+C
ZjaXKV+yBHFkGSLZQ1d8elDS3K6loCqh74Fbvv5oddY9wBWIK91g108MtgwK
EucyhQ49lI0MOueJEzRG4y0DeQx6ZYO/SVJALoyO+YJr9nOem+6eFOZQy9QQ
5VmaKVOfTk3nTIiIsdjA3VBAhq1feL79sRqBQhaDYvBY77iS92dGH7vsCt8d
5zFI+Z+0NsGDQ1yS22wD6WOXP6jtLoM6SI5adkBGq9T3njIF81Ph9AhtL+Cy
bthBQvMFOM2AsYPcOPl5f5hEhXOlYKawfOgD9NjKiE5b1kdNK55DVrvD41Cc
Bdo5kI01mvYws1+orbz/9ycQlV+M7D8ZGHYkxs0SMLbrOqKi66S+vbrfzPlL
jZbCnz3jXYP9PM1Z2RGeag7+3MDNoqvc15grL3NXm15P/DQ8PwJ4fghK5+LK
YAutgvHUsupkVjVQbdq4GnkZ3R1cJlasGqBEfZb1mcI5hrRw2gOBWFz6OELz
+ea4ztlkqD57O1z3uhmHg+JgfVT7TYxhOY/JsEEFTmMn1F/V6Q5UcyMrHWCm
RPnFg7J1NUxFkhQv2Wd7CYgZjPX3fqkBs8Zw7SXu8ssZ+0h3yNeh/oUElMCZ
/6ewMDVfXVMS50bUrAFFvZ0Hg6tdeliYjLokVyoI5SdYr/uGIgvkve2uC2cR
cWfXIt2kNT8DtXCBYPPnX7wLBzdniPmoRBg8mB/6Pj0dA5x+Y8OGEOzAUL5g
b/X7GJgUKLahXutMMBgmq8mbdtHl9MKLiD+I+p4pA1wvkBokFf7z06gwPDUs
1b873rPS6sY3IGSrCAsATnTj5WClj4SZ74fH/yiRFNGSxC9aL6YKY+M8lr9S
utp1AhZUtMLNc5JDL4t7p8s1Z6JIUwpfCyBvtn+EGtK+l88rntOK92wUhKuc
Qt2NbP/ttmLLb+Kvk4YNBa65y4+t5daMqEJCce+BxtKKf7BVYLce+bBS11sk
5LTlQCn/1Gb06igugWYN7/koJ8A785pQbhdJ3dZQpbo9cJSb4MqTxmv/kMk3
3fwKSUEV/ZAkO4Ayme2X3k+aOrv/B7RZk4GxTCjtVB4wDPuqEvXvgz1jKAfx
RKVr3BGj0Dh+1HuM5KWY/ZBwspouPgGACmoNnlSAAWAV0ppn511cZPy+KcDu
2kAusX+UUPOwDv+fIjT0PpMc5fHusURFcpLzChy9YPf4ZsqyhWeKhMUAQ/9e
EDVhO0qCq8E+C/Ji4iEvEhADWD8NRzXuVjvmyuE8Duvvm3bQX9VUH24hKbNW
VvFPYqp5Xy8bFDFeMt31LnSV5igFJ9l/K43KgNKOo487qBqzKZoQwoapKjkd
GNoiJb/7dcJk2Ib9q1DSre/hD8U39AElY8tdBFso7BzTs4oiwL971hgvhjwb
q+BN0gCxM1yt71Bn5axDjTH14IdKN1PNSEthnDulOEYIvcTgI9wGpU5kgiIc
5/ij4mVLhnl1skXv/VSl0I+/I7eS1rdKH9g76FAO667QwGzg5C/O5WB+byLp
VyqFVGVcR6G26cPpxV6BqBzd2x310SulKMqMowAciYna3Yn9oVSW+IN5VC3N
Ze8XCLwIInXfrj8L3MM8UTRpaAiJQBHn7bYf4azdhP/Bkw91H0dv+AwPp09e
BYujODSk1A3lbTzAEyyIcxQQgfWijx1e17Kjl5mDHG2c8ZeD8JC2RrkYVKxQ
8iP9P3MQhRaoVHQ4AseFRt0feAGb3ZsTzDMcC3OoBbum0//XY9t1PiP7pJ1B
48CJrQS0tvjXNpathxFDUN60VWy6ZfGeZbimriPTy66pBjM9RnQnVYN2wF3h
0xGPrXys8e8Hd9+S1W6ZOL0SDvoWlJWb6EQc8db4IFQI21mG2jGsOpIjJvzz
UXOSipSNgklV+vGN/0NVJm4VKj8TvexI7kwuD9f13T+GT0Y5QO4zVK+J015G
l8QSKFTbKO9P371rsmUr8JViF/v8eD6vWPUfYPQn9x3adCy3koBkePNDjOkg
dHxKMDsqRxcFUPTXlb3oWIM22xFyMyM8HlJtFgF558JB6LReN+pXmT/dLiMb
xH10/auJmXSfL03MXuKDn1AG1VUc9ysQoVDxfSM9NXIavnnxi/fSSA3/Ppt0
aZEVahYv1EkSYmuwPa/NZ73d1Sxrbs0rzcbyo4g2Vj4RbNRXjlyoMXPSEmiI
0OmRXUj9bvTJ31yPxO7Jm3X35atyCkRSI57WoNxFw+sBe7PHoHUB7AG+SOfN
f3ldUimwuDlUFJ4u2L6zCpOsseIC3t/9aYwErXvgf4yy4T0fIYuWrdJzLRIO
WQfnHcsXSTjG9TJ1sKRHXXd10/IGgPOPJ4cD5qmRMbaDUyR8C3x4a6vsPb0g
MeOQSuZS5b7ksqe3JNsSi390pWvQrf5wLxrEcI+UfAZWRq845F/hpLjwEYws
u73Ly1t5l2ENyZ9IZzKzil4bTgM+ElcULNRVcrvidJRWXNzYWV2n8yFZ0DEV
BSBaumOdL4aw1awEDltDQ2zot+Df1iW7k2R/X4NO0S4FXOJ2vVHCex4Qz7EN
rJs7fdWX4Su7yh2CUh32bNTkgljj6tR8L44+EjJdA9qipoxms6fN302bheUZ
u7i2GCXWMjGJSDTBRfKfdvUN0TR2Zes9WE5Pf9OajGKssRGXDCAn+1uc/MRW
2HfUW+QKnYIBKMaBzJFPRraxXB4HdWsa0hRrjqvp7rM8O1sWE5TAfuJCbQNF
ID9UwBQHnk0RE1z1+fpvMkXbBCbGxsSfIfw2GeorXYoPQYY0/1k7azhs3+2I
G7MCPbhhPum2dRVctlE158TcVQHE0D/CHrwoVvF9I+1NgeeaV0YlJdLL1FhE
Y98KY3F05fGor3SgC5JA16HtiN1w4LJih5bYkyi9AxTkRFkvIfDRFo+EOsmf
Kvu82QlxWRO//WAKK+8rlz03et3rfDfPhyD+ZmCk6vFzc0qzGVJ2NmhWINw+
ahy349gyvEQt/yb6dIBnq3il/wPE6QBJNJkWdu91rcZvw5Hi8wp6yHEELxRU
8NTYlgRchlpTifww3sLjuK+C9R9Uc9Nvud36lsoThAGFONugWqNi9yWNnH7L
xiv6hvx0Mud1kyb0WJuDRjSiqzm661UCSAegdLuwaqtoOLP2YScApdBTeFG5
/rNFRatD6gtIDOPwCOlLfoXqHLw1EBMvtYcpRfhFe2uqOjcv7/Rbp2MoAoqQ
FZtTnDDlMbAV0C0H+DNcYcZrzLr1gwjXXffqRdTM7ILoGhCG/gWbkHxifXQ8
5W9ZhA8wyeyBv+qcxjNK/ppLa+yc6GEjUxXKZ963SWO7vnqAZE23ZxbvGzjA
nF34GYEdJCq9Rfnh0NHHG4dMMk3vgrmUrdcjQwiYJg6jLHHEV8y/gqKw4OYz
uwSm/drBtvbOH/ZreYH8Rwp9fIBQIdoo8w4QXNifHc5jufMK69fIF8TmFx9z
fGL/aVdlx34QLFNRch+VEzq3i3X3wcdo/BavQ5tYWHlYGpGcAiOpw+0kIQ7Z
BzxdCCBQhxYAyCdfN3t3J/DzD+fx1iAM1A0QXmKGtvelA83WjxwwJkGeT76y
yRiWNvy+rVg9vHKZpXPYQ8GfcBF9+kMB58cjjIqMptJAF9TS5QyMo+41iAyW
OMDUHiqApBEAqKOg9pxeqTYGh/VxxlnXEI7DpjNw4qsLMICygvC92ws1tDIj
sBcwNoG5hrxjxGEXnhQr18HEoiCZSd66KcfJyT0RiMAEFxLIc8kQlul3Qti6
tetFm+tqClazjWUKBkUoPC56pC1MHqOPc3UBW8GkHqxIjursoViRKjlRDhdA
8jgH8C3xd25YICLLNRbtsWQLLm1ZQBtbKFANL8rhirfM1zkV8Hel3kenv8oU
7ab0dUiRvDYPVSa7CmIHxKuipxGCwpkNGFCyMTrosCLBYQgv4xZgWzfiOCjS
nWTsJXz+FI5UbD4l/tnDN6TQ4dX6w7bwgmJo2BpfNbwQr9VKX0BpRQ1LIsmq
DdXID7Eb/jTWix6ctCLBp8xnpLC/QrFCtWyeQnqMhhd7a1z41KMH1I9FqTpu
bpWIi/rZMsNZjDSDVZPM7hTb7qhKPWCLLSaHtxUlEFPB3u3gyjUhPPNZHgmG
jR4ehYAidZ0jvyfoQZJ5o/tRMI0GNFJtGUwkZtn+tF743k3VCi87XipM64K0
xK2k52N3ywxv7JoWamc7M4gkXV8Xl1nUIBjqeFBGTUHwWHKjDfoDCNPB6HVK
P/dn91yByUPLhkMDxZvsLwu/d6xS4pKo7BKt3+K/32KDBKsn5HDtUmGpldlL
s+pSjyANUB1/1ADt7xVKkbZnOFDrkkgneLjttCcv1klQAuxoLHDieEtygFiU
2o3bAoLvSP3lB2wbxfSC2CyW+VPYReeBMBv53Gq+W3jxtPHDNnXGkKgnPHL0
enoKQv6fwAP49YS3mD3m6EwZOhO4NbAaqf0Qpd6mgjtn6b9gCct6+XdbVLVh
F320LgEiSiK1HjK0x8XgH2lOMDaX8Z/Hu3K52mWb9E9g4Td3qG4J1IbcgSu3
QDv5+UEsGC+yt7sw1OqAPs5nsf1YboPqrcdKjy9lQm6LIdWWTuvNwUQuLlx3
uATgDsE/snVr+uBtixwVKDiRdTKX5lZvb4uxoqw2MazDtmIbKo28Dd5YuLSF
gWYwif3IPCR15XK5Q2DvNiuqx9kxuaTUfVdhC0OsR+9fGkO2iKasGt9o1S4y
Lo+/qFeZ5FNoL85JgrO0pfZZ412179UrAjcVA4WTN0sJZtdGN4lmOXzh32Zk
pr504MSk6pp3F2fY4s8TrfyVqL723RzXH5uAeA0v5ziaG4RHXJmkEbQV1Kqf
uOpRiwT0y84d6AKjrZP+tf1EhYOMqnev/9yG4AvhOMf7gUkbu8PXRliHWcR6
Niv55LJzX/c9HA8l0ACJCciKwB5sb7lQXDoNroGmEOxZU0mboQwIjzdHAg9Q
vkXjMvfQnvrzs3rRAI8nWIIQGn6oLPyb6zEIy5VynC4fu5+zkAHiWL5t81h8
Uqzw7wsNXV8B0vfbuwJtOI+NiULpT0Mq7eFp7S2Vs4pDmxG5Y3m9vIrzkjpi
90uvIaezBwMCuumPW+xpjhL2CvDtZ2fm6bZZY1SQiKwM42tEWlnI4n7Ys13x
HNPGV+1M8s3n0TWbCQQemIMOSDaUEqf6r2o/KpU5OMMNVte7opO1+DNi4yFu
sKG5XKFVYPfuQhsNe271o9h3MSHfHZoS/hAmsjDEFKb0erBV/Dd2igN6PS1/
MLUvGxelWQ5gOx9tshjZV3DtVgdGoBSNg2KG8T3zgDGkY+7092seYxJai+Bg
ARGkLYq9yQiaXVTl+wXfwAWid5r/qMUSTgwmnIer0MT5kCb2H/3RBFq/xPKf
U5qMIwov920PfYmhwqRbJv1RjvQRkwwKSzHYTzRG1M47qddfqqwitdMbCdjP
zlJFCmbEUwK444dauO1HxuQdh/kE1KRHFqn3agkpvg+H7ngeQsfWjTq/MyoP
u6aAL0md1boA2vEIzhLU49++JDQN6OTbagLMG8+tbQumPxIJ//4WyJ+NmpI2
VrEp+X9vHlrRE0L2rQlJI4QxxKhwPMqIhGgebjoP8i/7vbmeeCKWQ1L1Iz1u
mWcbrJd6l4j65Cx+u7gCHr/uwVowSUdKXYf1VQ7G/8fpMUeEpAj3tgQGc/XE
lWfDw3KNWBM9keJAvWoFtxLxTQIhJnveFYh1imSYCdLRKywObJdRdagNYlu3
QQVxq5sXIKSH9BqmCKDFeJ2z73Xyzw8VOzn4aX6hYsBNtC9UikeKVSHG2oty
4TmoN3DPHszc6lVfFySWcAL8LQqCT1EQltRmtJqHQ3PCSZOx3emVBHuTThB5
ncNaRZZM394IiEanvs2xfBN/golMcluvRfjd+S7wxmTzoC1PUVt7G8LnasEG
aRQgq+IW/u6J6+cFEzDh6PgJ5AFS5fqSmmOUz4piVzzyKDJj6MnSYnBj3s9N
+9RgOneOs1OZDP1npjV7oQBKziJgCCHbUoX4Afc+/R/C6jgc99GeiKIGo5fv
9Gkj4+1e6dW/OU3ByLiW8LoukVq+h9Za04E9bSDdgB79Y2uWMun0ZywbdEiY
c6NNclYpkjgqw9iWR7MbyLMJJRg1N547grVet9CN1igVFsf27sOgqIRbaz3p
KOF0Vj6ljEYjF5KGcwJLGhW7ZMuhR8FhDNZVZObRnWKypzILEL919v7ytDI1
sRyfjMEfJVvjeThcB2IQKhnLF1xEJnz4EeikwD0dxgFuArdGxK45MfY3V3Bx
3uTrvWoh8cFqO9ZjyxNRxRaAWCaoLAdNjjAFwv9ok4CXHYGGoFkSOVYHX/hK
U6gcQ0HAqMx+Sz3PXkfRpo7cp6quNZHftJX59fwD3zrlDa9kdkJeotCi+205
0pzAqQSY+uG0lHCr5u+W0r6yiNwoDnSfoja8lGngrobGXykRdhKXg3NrTSLN
bHRmygLIySaMtUfZ9A2JbcsuSxkbi8Kl21xwIrYo9nk47Lzo1+CuoPLJiDPZ
9DFpEvWLQxLe6LonqXbGG1JkXRZyIs2C1k61vULBvW0RSJGVpcsqtfWEb7E/
jXum0jNY4fHlQl8lHjlaoM6PTDHLRvm7T8ppnwB7PDimUWlSCY1U6LQCeCYs
my65q5VRSUg0lF1Slve/PkKpUX+xVh6IcBc1yWHhYWqEHSba/CkSF+7nWmUi
0ZEaIJbUnL2Lgr8CBSFg3iuEHmBZKpWHjy69NxtUtH5L/DsieX1XNclB2gEX
gjkcCSpbmf9mkCHCSuD+dEv5xCYcbrJLaiqG/vqf11h/myXN0k/D5Q7HeGMO
uw4Co/j+QtUWIIIlhxhA7hO0DHl8IYkdQjJwrBLw9z28uhjl8xRqWuUUcQDl
oTqERr/Y9ll7+sjvi0lCReOYWeiVw8cgr7BMP4ou8Tjb89/P40BiVDqeGkSs
LroMTCb6hUYIO2Kr6uplR5IruVbApI0jF8lrTLWZRqQnoLR6dbqY3XNEuewU
WyVBhRkKBMuKUsrScufU5Wmas7ThQ0v5wsWQ/zm3gvSvqtVRWBKTwGlG5Tdi
6XMXX8XEcgp5fVfzllK8XCtv3hAe6B5JlkawIqIPoVGvn1jlH+LKy7jUGqPd
vDnPc3rHecQJhoGg0N+Rf9qg4+22VeyjbAGfhiJ7aA+SMYPwbX/eQM1RTWur
+QYTCyjw6Q9dOWDR/3fGM6+IzufMDd2nQMr3iYNe2LV1v9QOQkaDsNzFYDg3
d/FKdQrp5eaDAB5n9/CgCW/IcLxvL1LjOU80oNg6OM0nB2Cafsz+HkSIhvy0
hMI1nOPh0gIAZo3ZF9mJfUR1nHEZHD4lf18wcVQLWPU7doaH/g/EFePUqbHC
F858nYFSkv3bfRQQjbcwiu4A484sulYQTJ3uYufVVpvFT2o5+KLBKRvmHg4Y
4oD53iQXgZEQmfndqSaTgP6V+r060/0nSh5uGzs9W5mKGytTVN41o6NZqjxX
6fWOxDl2YXSS8oLXf8s0hlEKeBDd0TD91igHvLdLi1U+zMQZfV4jaTqbcVHR
zFt6dSk1q/UGAtwglz3W4f1zjkXETy1anwL4z+h/VM7wQPzN/kdaZ1TXYM4z
Cc6jATWQJ5wNBfb5TnxyrDjUABRqF/+VIk5ylUbvO7I4uF0KWGqR14GeOuAB
v2pfvE5di+a4DDu6M7h5qdaEpELS+tYaGAntmqj5bBxHYybof/GEaoOEofed
YTcqOtYfudgfcYTcySyI4oQM9bt7rZRw7EJRtZTzRYxFOTKd40jnuECNKq+j
dDiioA2kgK9Pwq/kbfn7JtJp7/V3TSVvu07IVBIVPrcnuMVP82Ff1cjphNFF
dMYE1N71bwAxtH0Mfm7jq0lHQ1fVNkQKC3CJ0EUEuNwg4JbnpXo+57RTVrj3
/DNf6VcwHYWef90MdEE6kLgbUHkz4MkWnFEHKMLDKYCIihQ0rSKZgLYwb7JV
13kN9drOs6gH5dMsgZBZV8/B2GMw21MpeK7vlhQmgyIRiXePOAkqTamtjRFV
Lq6+29flDGarDK2/8NTlgFo3V4blDbJikfHJ/ftSg08h1e95RAkyJoom9mf0
VGmYr1K2Rd+CIhuHzZK8C7Pg6L/jHRSF9EADn4SxTRjlb9qg7VtUmHjkY0BG
VIBDyVHFrGKiZU18mclLdPVtik8zGs/5Xgo9RTvqJEwA4fx6sk4Gktcf+xcz
OgbCfXAPBhNUMQ2GXOtNK+LFUWnaxmm9GZ79Cz2fAjjYJnSs/N5el3hS+PPn
tBcwTc3kt5lIhQdejmmrnmqry+cdhS1AZ+WECFXfLu0Pe2gLrfG3LwSD1Int
u6/jQAuFAh3QmZ5vDhczRRRCyYv5sotbpQpSpjdC9C1EWG9z6m36upHruTJV
PQ0cRqlahV9URXX3afQzUMBRaa2TI+Av/KhY6h4J3t63YQbjdOWnckvWdaky
OTvXn6DG1Z4AzVepikDid5+MZvVXbIihNfcXNMbQ/JdYitnRIQX65PxhsZ8U
HOzuN7ifRnmCXwqxjiJns5Lf1ohokbV9JsR14meC2HHbm/D5pFsMPUFuEJJT
iFVmL/6B620fPvePbcEpKYCCV1FiqC9a4cfZPda0uomCrpXCSSy0pT55yxwc
wMfDjoeuoLpm6TTzrVVhg+TCE3SUaddG7f+5Cj3or3XLqxk6Z96pIIz9o649
GVKuILOsz+A14n/ngB+VjIGzUdlfDHFVoEnmMRcTX3ZZ2o5octYEd2vaTByI
vn6i86FfoaSJZN/FMeHO8lrF8Yl0FkV9AgquswiIxRVMGaO6/EHE7SbP0lyZ
6HZLBcp874Svg+lfu7eFYX4iqW+5vvZphercqdIPHsEByGf+OFU5Pf9+9Bdx
Cp4yjtUP2FIbgcWW+DG7mdwh0tHdY91UKp5Z5vX+f0dgMKI/vDrfzlDrVycz
/SJE4c2e94DnLaMBwWeiGsAVUDHYZ4spx7RMESiZV64jfToWnwpHssEJ0s3Q
Ij0asn4nO7FFep5XE1n68bYwwxooDMjv/9Wz56aoad3xA/xo5+UBpOFxrw6d
Ni8dd3ROxZZ7oBKjP8VG+jmgE3jNoyMX990mGWgD3ho6aiZZngXr9sugW+CA
wYVm1/CbzjL3UUOZYGmTp0MHFqSEquS5ye1EQrnFPn6ChJB6gSYfxOGeRGUG
RvQ9n5ai1FhA7hZNRGVkRobSWNBZQoq0aLQ2o6k18N0Gq16sT1Q8HVVWjTID
aUwgWLe32T6PS+Z73I+gwQzJF3FwRnGKtRNCYCGCXtfh0sqEWYAo0UDAIGQj
oPi51dTuaVKQ4Nly1YW+YcL3n7p8VJqAMFVzRH3REPMz67Y19t3IQgxodcgN
7P+20Zl3oSJs2NrsBRoTqX4tYk2sS7QbXv0fKdOBV9gDRithnxgVDmqOV+5H
KzwlJ8dNamnMTZdWe6VmESJHYywhruC8OPmY2Y2mslpUDemth3c9NO/uA9jI
CfENpcEga2IpRpxA1IsxHC9JJHmiTOcpH2RtvotiC1PovSAmrDGV0gKwCwy1
+qQfXWNx0zHqyA/eDbGNTm+MDh7F13eUJGQ0wsO6ef/CslLmQHhJPvIYRVNS
emUS/xJWH2ZCFQHiAFplCTvAB+GvRDT8QNF0qPj7Ord/+qzcIXdIChsqTCgd
49HsBx+Z1QQozH5jYzM0ERN8WnioyWYHrvIa32zTrsunXRKhiEGS8KCOUP79
UVdqxkLxLoD0IrQijtct+EmxNyM38SzJkK6DLWfOMJzJx9VehBIcgIjnQHx0
/gSGVBMb3Q9+5fhpXCWzuqNU6hmADuIMniw0jgfoVlXfCgwOhAIDwVyssCqS
7xteI3Bw5eCeZ9STtNlarprPfnbtsP11pzoeQu17GGoXUexOAIt98jLBVSNd
cmfzK9q6+V+s45nBGBEtDqHwupJU5FLSQt7PuLMcZz+PHlFgwx/opUWBDBEl
gvoZFcKA2gcq/seogAvB66XqPUOsByIhb53KmB63z0zfDJVroe4xIeE+hvPD
5GYiPi5YmUOuLIDTu9eSl7jU7LLw+yPYuoIN0gBXm8/vsyE6NY6PQUu9XtqZ
QTiRwFj8qXPD0lU+Kh74PdpDFGU2BvVfZ8PaDo9xnu82OcUwjSGnRYyH2YHW
6iPvc7C7MhQPgBcuPdFC3H+XOl2jIbahRK1USUKfv6t7TigYXKm6AtEY95Wf
mvp7iCuBxeTqm4NbPhl/x/EL4ZrIlOgPyOs0+G8xtsj15vLB+zAwOWeLpSKw
lt5Df8YdYu5WV8Ha2Pm6EeWcYlRhAhejMxe5pPb0L2Q/S16SC1oclI4VTXwh
MYVUXeWP4aVaWhln/b3TeS3GwYFP7O7hBbNhgWZGaB5iFZVaLRsz5VaFBi2J
lVKGJcSoSw2g2Fws9X/+mJA+65szu/43wcgwGsvbTiSoyyXEt/Sj+TuZhMJf
Q5XA+9LoSuCEBreOY+gFJcfedBbVqCHwD1V9cOsb9tmx8o3ph1DD20RsP/kn
LwVIgzlowsxqad1L5TD3B35ZDcRisdGg0vIdChiu/ysbMiBlwN+oXbRUV3xL
8VnBH4WS8oksFJGzv9cY3aatNtQ3GkPwv/pmt6MQE3caF97fFA84tYEzHHf3
TyF/e3h5FWWKbyrc6tgX/Hh6JUCaBxPJuix6f2Ngtgiwlmn+hBVUQ1NiE++t
CchshfIxyswylkMDnhxIIwjUU108j6ntegCdZaOuw57a71t+hRjWUsAT9xFQ
CJFqB9ziDP8J7zm86n0CUppqTkYwlU5C0Au4lRpIVDnOiKAq9xifHqGNGGBB
d1UhYjxyLZrV3afemhZbw7p7CT7UG6VIDElbREkuckTRlWAVND5bli6GlM8y
A0q00uB/u248hoySExzWqJ/VoG2GdQhqMPHtcm0TNdjzxEKfN1BNoVqYtZCz
iKzEBOD+aTUecWDhmeGhVgKXnz6a4r3IVE46klrvKDuUpDuwTs6aRHla+FoK
d9240EUNyzpAA7KUACKHcSGx1d801BetJRS082uIE3kRNxHEHKJzWksPstDP
ewB6P1dXcomEl2E0VyR65LrLPnCmnFZtCdL5JfUlZz8uU18XGBTAJjVs6Cql
/tjrJfQS0+qP0M7uv6YOKshOZAkiFs0yNTSoNC1iqQ/S8dkSZt4CVEnXlyu7
oM+6lbbYRjFIV/7fn0ogo0BKUi9qqQiIpD9B2M0QUnApnPDd2tgaSybVOBNf
8X+VZGlYKGbMSH+hb0salwAPsau3jKpfPunsDOgf1aA8n4/GzJg4hWj9ZKvy
GPfZhDSSjZIejCLXlazGq5l1+rQX4kI17zgHkUnxw6efwUxDLfcODCb5UJ6K
Wd7jpEP7lcdd4vfx4b6FdhXRx7Erqo6RWob82kUAN+lPYaT7TQq/FczESG8S
G9eq6wcHlohU/RI8OKFswXkhnZcEkq9X48OIqApJ7hoB/on75kT2q9cELjCS
nyshtT3ZASC3AJMGC6a4Ybj3BAaWYqHLGCBghV6naO/cpNa6U5qL+BHBSt0Y
DRhPY5ev+9RNBMr43hddtiqQ/QP9NSRYC/wJEfF3Bd6yM70m16d7MWfYyhqC
1FZI1/EEika3aWPANGjRE46J87W4eAB4tZJfXCKhB0UvwZ4k5Y/Q/BAfOj6K
im59XJXpReAbAlOQvt+PDUfx49qzjfeg4b6lWk9xwHY1/m2M2cbjJPtI8t+J
ewGAK6wM4AVB29gBMSolOoN5FXTi0HQ9yJh4c4SawNt2f6eO7day3cI8zJv/
5ielhrO1225CKsIHX/oP8o5M53bgvrIp4yvJWsHrSUY5PB7yZ5kxobIqGdPk
3sn0aGaYXjkb3Z291B6Hwq5zHdE39vnOLX0fN8VTkcYAjccShVvxVVazrmKL
a/fDOs8GA0uyiF9m8S5zlpmPbq8cTGHkyzEU2uQXPDPve9lkX/pvQwd/Bvpf
U5e9B7cTwEJn4DYJxkKRU0dekOpA8Om+e0WwwsgNSmOL++GfSNAGMQkyOEA9
UXawOyGITtHfZGOGU88yln4YChpSAFU+4G26cJX9SWSfBcDnliv6p1do/ij7
qZ9wRML9kALZwehJVeMl/lPV70imODJgAd5vWiDrgDar+jAcDbgx3PztiZdc
/jJAko442vMfegmcH4xjWEkxtXjH6gQF426mEzOv8TnvIgBCwfcE7JJhjQfJ
qiVlwe9iEu9rY/nPSWpHrmOBZl4jz30vg20QNQVcaKP6F+KlE39rmJUyFD4C
yWhny1toeZw6abDdPPPPTBUsupz/fH7IcaWSWF7QStE1epbldXp6fpx+70Va
80Er6F8B0r+SPZxYMacHkLYVDsV4MmdWf6TjwdvitovSSG3J5D6sJ+oBgZlR
4Y6I4z8h64Bih8LiONGVG4VWz+fJw2Q9Ea3D52GJJu9+gqNxVSAnAAMRTkGf
u3y71RxMfTM+cjuYQNzQDeSR3sIqnX8b7BtwzWSHeP42cmyNdDQx87zkU3Pv
NbTItZYBrzl6MIXBMR8MBeQlfdWEecKqFRsiPVZ006xzJt4UThxpBJD86Yuh
lvaznRWSxN1r5sR4K5XKc/ihDSfy3xC7sGtIB3UNb7amW/bE6ow3SgrkGjhY
HrhF1wRMWhFliHk1bPWUB8GHhaDvjDDNXVroqQC+rV/DS7KLP9QAx9B7Fyqr
k9CSVVsxBXLl18iTvhKCF8aSF3n+3j5r93Q2PkZchPgJpiR2SOpiA6xc3eKQ
N9VxaDLAmxkMmYklTP2CP5pgeXJ24hvfH3Lw61CZ3DLLsfgr3fU0zsW0CWf6
W+6aLTgGz2wA0gBGpaxTIy6E+nJlT/3wT/Qec/d7WDbSYUrbdjUYsdEEaeEe
HdxlqPniDngbUgMXZIlSUoWOPR/zAsH1IQlDmtYZ0k7Y9pZx1X4T6MItbayF
ripNYyit0Fs5LmEIqH3Qxn7tU4Z8d/56IkoPUqPHT68xi/0ydKWi7KnAhkAS
HjZrljxqHRhEejAwlvoOxRnryCuMcYUu0j8thaCbNY97fVl81yY1XuYJayfs
WkJ3H8Ttiw3aRbZAmEtxNPUW5aV7Ps/anHJpnHBzrp4wKKWPr+cDcNbmqlMO
cnGKJg3OyeZITMk05k3Hk/7sb6Bve5ZxV1qRO+jN9BIe5OQaivM1YtWi9x4X
q7mFqnkfQUfjN1yEGYLnqlVVGNFjzbBygKvVcrgJ7UC/potp40snKUZ3ybY4
TuVA1zm7FBz8C73uNVQLsQlL5ohlCO02W66LjZZRUGRNx9M39mSHvu14xMBo
HbQX1rWMNQJTSjb+p5nbbXf+h0nl7eU4F3OikjLX2kOgkiq8qGqhYEYGeq1t
8X88rv3s2J7BQw6g5niBmEQ97mmnF6XYmegjYq7OkQHgxjBMFfygg8/CNdFD
Kp499Dv1mbq0CT5MEWyjCGVq3XnV7jwjt8gzKvyJXJqMQ1fpxZawnFijx5Ne
hOS5dXelCrA6DD8j0inyHsv2eXTfZnfqxaFA7FFHbhOlJjs62ooDIs79qWvo
AfeCD8y+col5463xQClxKqEyoTgX+FyBg0XnDp9jDX1o9cIKvsh+iz40t1Kk
Lcs4Yi0Cbx/txJYhvT3pWA6cOUHGAf/7OcPQIWhHeZdNz6uU5F9Hd7wqE/Zg
46LGT1yxnAi7i412VAMnnKNvieKa+CffowvJqLhNHoRHuV0fTemIFHuFD7Lg
SBniuIymDkCtKIjTQ9+nRvj2So29xJHYdra7UXt1NASOHCLmd5s184M1l9e9
ebPs5THS1TOPBhdelzfbIF7E+VtKpnJjrRti0WcGzxYc1mUfMcWEyBJUmVAt
Chm8TRc+5AcESi7yvstv+gPdhfclzFLGNvE0+I66BCg6FWM1GE2+/YDhv6Q1
bqGyW8bWXjjc1FQFkk+BiIoVvO9rzLRUhjux71+SF/kUimgn3mIiURbO6xVu
+5GhsNBUeA+wjdX/Y6SpGQlujxzhGDldv1DGLR4vJjQuAHH9deE4W1l+xOP8
U9xjeqAYgPKtyxLrbjIYKrs+GPivtaYpkOO8MdLPWiMreelNvR5P/IAYQvEp
XJJ4MhhOwnCPiV9XHcziZRtj//FGiPBD2GcZPmhyVM+0YnnHQW5DhXhVMKxI
0dX+/uPy73EjsfwJC1yW8KsHHWe3KVLdNed/bCxVjFRfEcIr4G8gltHSwTcK
IhARUi36Wg4zkYwR2BP0mvbkTE8v+jP3NO/ET8prTdiLI4tE6jw9su6IHGWb
Y2HyiqfYpCcGjmpSgManG8FrGGtgbDqzqigABSAT1NP7pf/PJKzoU1tjltGk
rVoKYwMl/qQx6YuX3CyW8Zx8e2JEe+xnfNqCJ8D0uyyPYQGAXYpPOB/9IUxo
Ylx6FbinYTPdsfeiJSH42mXXBbkddsilvaxqdgg2XavcREIxYh6lQtngT20W
vKgzEd7ou0ywRyMlvmG1I+jHNomv4WrJyG/vAf9lt2OEHqPe1IH8Jq8lMh+k
fqtU/OqdeXn2QvB7POCbtZQvCJEZ9z9cD8m3m+dEET9sBicJChkXsGsSu1Ab
MF/0jW1dr/HhVib3eEn2Db9tJ14vaRf0jNqjyr7cbuS9WKjy/OKQlqRqv7Dd
5YvVVQ1/U2ivKk7ZCiEDZ0ucRLQ6u8gb+h4/NzJjdn7R8decEnaxRWdrwEv7
AvHWG4MWAa2Adjep7ZRKgShWBJZDErQq3QeMzbJ8OY2Y1V8ZnkmA7mhADT7F
tF5wJdjEP3AS500kenhFO+SNYQIZN256ATpUQ+DcKpVCkhdH4eTmclzhZVGp
y79vnoxqNDBX2bFafMh89/wHGdaWGvbpIuYGV9w+kwzA3XziarJXpqCC33De
EsXxbgig16N9bHlcWm2TTPBuFjUPgbWYnJ1bTYIS/l/KHgC5Nx0C//Pa7m+i
6uDWfQHYYeXJY+NsYfigxEzkYnQdeLq7QBVl4nsWgaHtNwfARQY4eSs07Lwi
CACz3OeWOIVOK4hRgtvMOVvc15PlgvDxT8vuAvgi0ndFJwGQT1RQmCNVKxBM
d+RQmCT9pnSPRd0GUrNpGLNyONPUH9A5mUSnj5z9HhoLehhx7lSM8iGLJkGO
5Cdeq2M80TELpOMvjXsBF5Fu0kImuNgRuHD7c0So5CJL9ti3EyHDEyrCb9yq
ba5jeUWV1xc/rhPlQFe3llMpuGhEh9Zozqh0goY8jeREcLf/NTKi8f6aZYZB
M/VRQNj5Mcu9wTzgJH/3Y52FsaVY9s17NWV/wAEP9Cxx26QuCsukrZ8/InZF
pqsopSlfrrjMxq1Gj7puVjhyf2eQrm3uOpbkO3Mb1j4OH+7oALyftPKd2nes
5keSZgK0YT0zTwI3VeHJI/rW/Ip76NzSfuDnUn98eDv6E4lChz3vmRB7GAKe
b6BDOm6SP7C1tr+1e06jTEMm3gyAxJjf43Hg4oTu1Y7z6k1rPJT04bdWKce+
zPxmifiWY3OJJUzSvuBPkQLN+iwC85w8bedv7BSmOpVH1UmQu1bixxNsoyBQ
wxth2zAcz9OWTGijzONoS9Z79ZgrZ7DXddj6IZDQGwwJOLG4Xtr0w2f79EUC
fWTFVBj8Y7vQXK+Sdw/spqwuG/PyCOvs1Im7KjLheHeyAnGJNaSGJ2gdB3rp
Jx53bGyL32WgiUn8+zFwhVLZiGXnUTPnSYp2tPhKUiB8AU4MF66I/F63om1O
OaVIDCwCe3x+EEdpeK8WGHEs5CC0bFCUb4m+baPB9efk3nt+HypWdKm6pGQA
XZ/QTRdb1spGXb8dWZZhzsQG6HSTy9oM1FZ+EP6BmBT0jCS1N0OcvctVcpwV
eEvAZquYqfgNJhdtrz//CNkqVJ1OyXdbkMS1VJizAVS5K1a5O5I8LozJoDfQ
YLaIhL0Q7iU1S+8cT1TDtzdt1f2c5HVczOfie6e18/trPLZ+7XKMotCES4BP
1KqFiW5844TJ7KCLpeWo/bOj8EH5ajL1SlryXdRMb6cm/lMq08zD1YAkYuf1
6tYJjbfgh5ZHVhVCwdH/hPUD2rkGj/sebr4oFCYO4AXYBxCdfjO169P9fAYq
hz+sGgpi+m9BjK/6sNnYenlCsCvaDNtV7hAUhq0+sqFycUO+G4wgqAE5FDtH
uhWZQ8dM3rnrehrj68hjP4UmdXu7VbLqThUnuHRAClBuxHjwWQqD1xckwQh1
WrYyXO5ih20O8MX4WUx1yaHAyFPUn7GDTPqv9S9pE2HxctrFay6XfVpHbH7/
atzew6+6CItfP4ZRAwPF1G80C/s+xKxhtoCSAZzHl3aqgV2BtXarL/aW3i8J
K7qlLw+wsSP3r5TNxKTXNOMMFcaGd/YPym+GngXePY8g/fltbjrSxjpCC/xI
1HXFlgSMf+vcJ9Pj/CPV3elmVXUBDOUPyLM0CGj6rab2mMbL6b/tOW2L1ZSw
Gzq6oJ8zqD07ggaXgfz9I3qJNRWz8EK8IwDUrh6WMyz3wuB6vCHMdP5IihGR
cPhz67tG5a4KlGLltJ6eFKkdTkUuxHdPxlFFxkENNdTSm7YAs/gNvOUe5U51
qwAJ7QXq7r4hVuyfrhl5Pv8cyKBOlCM5sRlCS6iBgHSSA9SbUF43eo1zQpr/
0ETX0plWmF7e6FTNOjfwnYKfik73K5TCIGvILpvPmqHM999F0A+7SbgpB3aZ
12cXgXCqBe3xPkHOpNzy8SBeM8zPcOGOqx1UGsN2tSOUQIfyOUI64Cc1Kh9e
ETjB2Y8IA5zHMg+b4X3sndn08A5K9/Fl/8g8euZ4HpEXBdEY04gYghRUxr+8
/5I8Y9VHVScRKMRFQImnNVLIS5cPWhyOre/8va2xXXvcmQjQ+Z5MjtVu3Y5t
WxNbHivLugGAM6CxJWfTK4crgu1gpFmiaAXKsC1fblGUis1lAp7+twDDUPmr
PCc7DbzZpbKNoHKEhNw4rIUdQjzrPghAZOPJj9xm0BqT/Wg8hWhepflH9Ce9
BYH1ZWPqKe9jdjyEvOO6+HpoHuqkJ4GCaVoKHLWrI1A8rE4touBAah8+w7dZ
9X5ycAdsk2Ue7+f4FamtaHvTtIUgvZjw4eZk8wK7XhfHUVnWlZFtGm+GrXIF
ylrXOS7yp9+sZu/p1ptBjtpkkIyNawWLAg+9+nPlaW6r2ih7z+3d88LuHsAX
g9W9n1mqQjdylZgXmSEGldWrArsQjOp8xmt7g1sYfY717QxCp42iQdJXqVIq
8Y5L0G3rwam39GVAslxrxuGIvbtRk9aIkEZSkmtIWXS6wmjvdbvMUzzrd6aX
/JlcQmBYU+MdZUvzS9CeI8fv2UIxeNnLmFrKePVUZy39dhkceHTHrUdGthm1
LMJG5BeWvqedy3FTUIxc0sH2T3FQrlaXW/o3cgngcO+hhZTALvywjYWvNi4B
xvqFy6UuDEJrG+aqQLW8yyDJ5iV5pVKktZucftYedw4+wPYTapHMwtVPf0PP
Gz2mloIMGrLR1dZjYRD0DUpW8uqw/Cb6xqY1CsuvtcmEWA0elVBzjYsjWgx8
0W9QA7mf6LJ3VIlQrCXYYmMquspMd0X4Kq/CtUJy880Qgc7wa3STtGK3zXGZ
aWoo3uTOlI5/aYZ71XdtDYtFyKpGofqLF4HU/G/pWcuSsO5+ms7P08KGG9eP
bpz0DHA/pzrAI8F+5F6jeOzQVGoGAmGsYbLLjJrF7a8caKNE5vzDzXyNIAfm
Kvr6axRU3OC20NewO61V4vtVukx8Ap+dp4cjxx4vO5c4gzuSaLs7QBmrwraI
g+7ChjQmeFz6Qnyxa7yyA9cd5Uk0V6HXf/m0QuQJfYU9jo75tuXyC5i0eDip
0q9USxYCQYSYVqNtv+w5rmqBTE+t/z0A/BA4ueIvcwg5PjXgqTaAZWXQvm/y
bhwrFryIZuWSY8sdG3C6ZI797IvlAeSc+u6RFAWR84Y8mCfJPkuD7JbMjRKl
8RyaJOoohiSHD2RFd8+umPPUlu0oUrKoQFDCFP/BsmnUMKkzrhuKCuu7wpum
fyGw5C461iFTQL5rkWUgL4tlPQn8ofR9FeaBsGSh8LTnJOBGgGcwt75KYeSF
8P/2tVJxuUf+IlfmcxZ4DpImg7AOj1c9t3Fqhk9GyqEsQguF0kDrtKu51/Rb
WwWu8Q9o5Tl9HJb4lXxEPAmW+Jld3HL9glgkv38ZldzuZIaUL7Xb4xg6Pfzy
lZMD0F3YTOxBf+1cLb5vU0k8xdlsXuzlBSoIoFEc+gwu6njJx3TGG8f7mFYu
G0iG9rWk0jsoeDQUMc3zac7i2Frr5F/Vx+8cFeIy2qF9jab7t2MaHTZtLScj
q7jJtRnufonCAyfaGnKv8hztvmG5gH/u4mWysOw3LNPn+lTGJAZUx70qS1Jx
ySkJfMy2CIt47/J13u35NPToWyIo2g93PBmugEo9hLQOoF4eC5KTDG7gL9wy
+CN3vNBlN+YlpAYFrh6cwRCrJilYBl4c++MhjqQxtWwN/gzq+lcFf86Seh3D
w3Op7/E+2IB4opnAX8ptkp1Lt2hxJNW4uQupuer2dXnp82VN1+irlt44Fq5C
A2/sej49xgSlozkFR9st7rw+JdXBs2VwncjUZWeW56ZZy6wnLVLiKt8FeQnO
1ihDXn2VZsTsAmQRSoVgwudb/wv/Qe6mr2JoaX1zzHHLSb+VopU7E75eM64h
5gL5ZJioEEU54aYdRaxEgBxp9JDih4+ARBU0w+5mWQM6iU5O3GEMqdUvGPy6
mUJ/Qe0aUaSXsbVCTxgYGSXyjZFrwyYWk9o1RKluCCXY3WoiNXVrOjFBjyZU
HflxdBnF0QVFxm2WVub7ZpROWlbUcpOeYWAF4pfwyM5JI8SMo5yC6T8dx9RN
8B+pSnii78OpIQKq4qlFXWghqm5p4pDbJ9OqmpmNwYazgCJZ4pim642Gdh9S
MkV0v0D0h2zA5FGrKc5H3Er4C5JLnjGqMSBYJkq7/qnymTJP56bD6aQ6503U
D18RXmB7nX4BpHZIPw3YQZEkz9XCVlUtaNxDiir+Wd1pfLgVi8pQIyaU38wE
NSx5HZ6vHA7xZclRjfWgyunEgWf2RQJG65uJBVs7gzMdoVEB9CZPwQPRFT7W
i5SPwG7FQS3m5KHR/Q2wLTfFuoss6D0noe7N//I2CncvoIJb01yoKg8TB6me
bjP7UCtA58ST2HsFUZcSN7h7QsWDoyu/tUxDCAAIfrscJ+SOvrTC7h6wiIpM
GgRTgwb5g3iyLv6jedSlt5ixzlJ69L23EHNO9tCN62DMWk+bQGY73IbNmp8r
8eGaBgaiblWFIuqo8jiAs2JS9Qe6iDjsgtNRvzVUECofKTTTUY+0pWphLNNj
Uu5omIUjB2WHJpny+rmvxyEJLgO9SABHa6kr/j3KoayJYo/FD/17qxtBXjpi
Lun4efBF5ilNtKEBg0KN4rCwZgcNR+mYcj2T+Cq1wUYQSwzd89QjSNgeDtbE
z1rPfTDgBSCNp5b+sZXcOr8LODf1WR+UKYwj9MDCBgTnl2mNziaDqmMTB1Fa
yzhcAKlF5w2VHD1F00Qpoar3EIoHyqLyMeu25mHoa/0N1cLRMbxeVkWe5Syi
UFYln74K0JMnObyEfrxazAzXUYVEryXxS/3itzl6lH4KdpxWbf8y1Z9j4jdy
hbY7wGzqumai5zQ+0K/kq/BE85liCML+Wqaaw/NJncjR0UgvakqYHruDA03Q
aQR41P7+6v5xG11R+ighI5XiWRFkbCBqP0FRtFdg1iJQihehtFSJ90RgeDwi
wfI8Nqq3rUNtzGwtyQs7gYa/3dI4/5JXbhVmyrGyvG++OEVvBmi/75ClBqAO
QAAccM+T/ylcPQF8QFTnKnPhLZYeCdbcIFm05znWgjW6ba6FCEtP3+LMPLws
WYjdsvJ5PIieLlyJwvUcLOf5Ud6+IWz7d8PJy70LsNAt4hVEg959Z0qsbzNT
aQq+GJDwSVLTd4fnVUfFSlA/rjnfOPWmDtHUCPMaT8H39zjuGrC7gHg1s2a3
zMKx3mbc81JCkVlI/TA/flmDt4DkX8utGptpNG6CDh6s1Rr6xSUNrYLDT+an
UdvqmAmpxovCRsyJwEzVhGrOBC+g+66KGpYp+YcAIr7d96sLJYx9Vtw+8HFX
I7XdygMw/8O25n8NcEqeY0gBULx5naJ/6b8c7tZ19tUxxJ6p/f8QPbKAtbAF
emAUG3n+bwq8WTYoiBwbYmobhyc36fpXb19VQdhU5t4pl1txIaXbnU6slZi5
C+K56HKxAwQg+N1YXCajJNlIQe6DJ7lMrYSN6TQ6NgTrytM2Bc5aMoZeSgdW
khRdlYfbI1NPKh1DMpaOp0GJrD3Zmz+geb7XCb7OMUFfzD7OTRM8yux8Pc2Q
Hn9M6Zudpl+QxaOWmtTfOPYiNdZY/rEzoOO/8H8x3jaPnjAUXTD8sxJkODYI
y0j5PPCstb7AE5w4KNEa6oHW0vgsd/xNBuMlKelly/SVu6Yc1UGmjOVX6nwf
Fgu9O0mef/r56/gk1N1pMhm7TSJIfh0ABoJXz6bQF7FZpqfm/vzPQumBuUM+
S3Z8Bee+Y2XrsPrZwI96yql+4nXFyAzVedDGjbjiiztUApE2tkrxXqx7UipT
Q+hOcbCZ62PTk9yZl7YW6UCGHDZgUKOcoi+DCSyoceSKr7Q3VwAvXiSBCWIw
5PCvGHlC+aKXx4KnC9kvV3+R5kjtmaYzhSjenUabItySV768aDfhRnqKvaGP
Zv9lYo2J79xnfiw0o/udtJS98DUugHsmI/xb2smWGTd8ThuJ/DPgUFCPK2d9
Ahpa/4zNZKA+qL29YUc980QE47d4zM0gRxk5H7KZBNJrx63UPzPZ+1m0sYhx
a3QVjhpSZciq55aVkzF5zNzdjbr7tPW3e0djlpzE5TjWfj7NE4rt78lU+w25
JyGbr1h0/dlJxhTE4DzvFSyPPojudpZUh1A2IusewTmsxrp/wcwvu9FGonnH
zAWh4RDYKk7ea03ZdxQ5Ps0oYgfV54STN2AymkxFhSvFRAueF7gnyg39C2K3
zJeFsSycn8VY3XiDSVMuSqrFp/PZ6MIn06czEmk0LwZfnf72Z2vdhPDaEJEC
q+Z5D5MRqHqKGhHHQTFsIwqvanY7E0yQ0dw8OBlRmAJ7C+6g2a+TSQsPEw3F
FoRwcIIpkd86EFXkOczqpqZDiLXTVCT8VpXxGAlpEW3q2bC6K2vi6l2ql4Kg
pG9EPWWoRP6byc716y/wD/V7UxxHFrCfnNShgSY80cgOG7Jf4UsmQaW5m3U2
eDaDVbUgOB7Mv15whLRA41XGfKT6Qakric0yuVp/qXoR0ikxjr8ToNDbiYhZ
FueH02v22oVXB72rpWW+h/DRCTqsA9hWBLQpksKLWp+Wa2tfbnqgJNkzHEma
9m3hIGvSf+Jis8Pr+jLuT73eG9AKuwXhAbwViIO4dzVa7vFpIvTkMm0Q0CAq
nHBtz/s1nUijG9o4euz1YIUXULRdlbu0Kn/sS3OcjjK5o0ikMP3gbqrAc72o
BffSmNAkXaPNMo073Fn/oUuxQPGMptsHNEPs5DGnQs/WTGiCbNvCLZjGRvmr
qzXYGpUmXZF+QUjIOc9r9AmoZNxSl5w1yLOlnGy+EMbrH7deugjPMkLB1JHO
tLwZ8xVJYfH96w5QdrzPLyVSte4zzzStjfrypd+uLSOXgbzsWzYVBQdqk+dH
3viUq6/VkKpr+iYjHu6kOQotmNMARa6TwhBQrTZXhdceYBJSS+5LdYiGXAZ7
1Ptj1ZlTSY/ZnW6Y/0Ou5GbkydQgY1vAnuuUjl+4Nfe0JDfihvIpU89Q/DMG
1DA4NqwJK6koNkL6kiZtuDyZtlyKJv2pMMiVUH2voyQPiVW9e2EChs3XyEUS
2T8UnMw4hKYKavHQvYmbNVu5URU4w4LcmxqUjUN49Vp3Mcbh0qmu9LIFdMwZ
AMWvjhRdoR3B3e/KT/LjE3qs16fynQgwoB04uLEXPt1I1gAxsYYNsg6k7VpN
sTvqjyOYlmYI7GStL+FZ6cjHEDXLLDhfq6KyYHb4muYzyNEaeYUpcgbXVnDI
cyboN88epz16/f8CeJwlfn80YO7OOdYl8WA5fXceZqIEOfZmstPPEvoxmz8C
bp6ewWIxtE3NWmZra59KQpgIxJdqI8i2tHXuzCgxOlFKMzkHXcTT5NmOSTFT
Wuct/jfQbwn3UxjYMuUkqmEsxi/boiyRYunh45mZ2aibwi+bBroKDyR9/x9A
tPXBwH91/WjhMKc+NZznY3FocPrY0wbYV0xRfWMnzS62lkNBJfW14BZBtJHd
+m6cRC6+lmvX2kzxmKF2pddbMhhgbwSm1CYAGI2F26rAQPxf/rK0f4cjTrNB
VHFcve6klbVh12zz+XSPqWtiirrsJ8Pa+nlHPyTFeGS16MLK/sukpxVLco4n
SszDVBT2JqNCz+544eOwlEZIK8eJxdoA2rDeWw7sogG+Zgaa+82zGChluXXR
wSrV3p5njcopJPi222chXZJK6AnQ60bgGpL4Vgvrb4SBG/jtEZLTKmKh6uq1
GNWhHBFqNsc0Cr3/sNSQECwkjIatznLkgZDPlep6d7P7a+cgTgZ9dvSHMRBg
6Xp2MSYkbHsXfbYsxLImD9TrGRkS0wHt9c5iUaxyM8w4TG+oxo+qOCmiTgas
2JYz+7dit9IgVQa+G4ruZU8ASFOeTTwSdKDG5gZJTzPnYwdtLtwKb4YE1fNj
PUkAqvRpeardGsH0NTozxcS9hOkijEaOBr4p4QsUXxxY4ZU0RqIQDu9Sdm1i
s6KJQUGn0Ywjqy6AV2cO2gL/YR2RzeEmD0cEn2V+geVNuUisurFGvhOHf7Ku
RsPFAvfFJFZt9Z7UHxOsriZtJQmQUU+yLnV2t4txlj3XhxmBqHpnjW9USXw0
nUb9IL5FEB/tMWlQFAtX9SwSTbBSASX0mx9/+Ibm2jB4ig8S1a6Sjo5UREsi
b297SsT3dSiRLzRhVr2q8NDC/cRhr1XEcZ6Ne1TouOdaFc5mNFyFQfMQI28D
BU/QmDVWXFY0tL2AHNmc+GkAhbn1Y1QpBaPodgt42ajKXT2GjrY9WJM0J9Cm
D7DaPRoNvxAv2/A7BzPVN2Bnq0pFvLQdLMAVT3naxRZw9thu5GAZM9aGzWn2
1IsTQHrsgYmW3bZAQhyG7hKPgflauqRXkR5YvS08A7VOJ2CcDLV24uSqFUxf
jNnJO9mbeZCWwBdsYJ5ZniUMzPJRgkLy6b0IiPD7O5i2sHDbRiyOIFj22IpN
lQrN9TLm4HooPFiIHXHuPIRYL6FR9Ddnj3aBvsSiuMCbw1RkRBe2PfTT3zYq
/PkcBn26b3a+PlHQsaKKy+rdEqZVrlkW+EgMzlb3/lC1DwExtYz2k6XQzSUL
Z2tf4AJAJudQAiQrugSmwJlLjky9fbkQpNQ8GhiDAnSEOg1eW6RRS4LeMlnH
J/C5ldEQ2sx4MSul75vFXU4MA2bik+jgPsONbycmPCky2PvWczVYhjLlsfmK
TbdArBNcZEqkrOFSLc1JBnSsvwjT1G6KT6jJZ0Ztl+V83e5VFwNLJI7V1GCZ
VfsZyjGL1g76KNt14AX5wdFHegG7gT6s8lpq81M76FJH5cedSFc6L0D7QM9X
DihvIVxa03GN+dwV9kMoznG0O7oSU62I0DCL80j9z1JlB5kQDz5/CeCID/DH
2kEKlfw9wvYrod5xWji8hY+xDOXucg/S0/fLik9gthbyUVXBBUADevVUCl5g
J94JG9nvp3IBTfw8yQVLUHq/7jEhaqNnfGDGjQrCrF3STmTK2qVkDdc/CBZ0
kL1NimcGYwYElYqmNVVmpc/n32aU7jZ8CrIHL2WE6l+IsHYTdLPcy438M2bh
SZnW1Cxigp1Bs3zr102qzGlnUgvQSUFIsDX8Ck+oFiBLMhSSP+xDjmx4hFwa
f90RxP2PwbLOCitpzT5BcAqPq97NyX9l+MQ3tpV3A02LbCcoxDstpkpemXmz
SrYHsHZK1u4LcVaI0thAe3gDw3zZDH/2c/mh+ZQjZHuoQVeTFSVIuwr5NNvp
NQNwiPgMEthL5+llP48+vW1owXuLPcGpJ3d2suffzmsIj2bUpoHal+Vx9f1d
a1cSEfiX0U2h+41Wa/gyDAV5YhH4bx/zjMEbJdP9IsxeCc18xEtkwHtu0DSJ
TAeaxXuUPJbnk4//hKNIA8lR2hrPVofIg+pQReHZqqCWmB/IE6tnijLSz92J
GZiEv/3Asnjt/nuKeFvBwZE1dnmwaBlNNBg7jNyTPeJjFzpUAthU7nGjB0Xj
g+iuXskeeLD9ZtFBSZ1IOf2b5cIJbdkodtgAelrbNG/mohAIOvBKkCTx2gUq
ihawJ48vhAoF2om3OGg42P7Z8aRefoFlISghF3H75cJHr1N3Xs9naP+9QA89
pTLg47ArX3NuNTyiEf38ha3pZateqtl0H9B7EU7fQLGmDkmEtkQ7gDLoDPdS
csjQtdSPqOEKOl+wPRTiEcPMwOe3V8WplOMTCXvDHbiNGVqASFTGxgCgITet
3L+OCbXhe8Gb6MsO+iLGLXlxXUXZKyZVQ/u2EtEMPP6jltdkLRvIqe26Kb6m
E6tDz2LZ00OLOdYe1bxepb3EYheC+ZaFdmRPbH17GjC0Fy9LdR3X8YSzRY19
5sA6nkF5gu5e96Do08ve618h+mRlkE/9dDydaz5yx931kbY5cGdi6dP/tJRB
JtH5BlXJWsiFP4rzcIzW1O1TuHBb83wmmaljKrygKyRTFiXdGXDifbOmABiG
CNOmGG6CwipRL8N2PSXwhYnBS8ZmzA6C33xmNBxe2bmuEHmzzzZXyVIZJuZ5
ms4VdVoek8XvNcmb7ZTDcxW0BHqxAVp5859CiYMDOVNNhRiaAfabNQaODPUl
dZ4pIPBFnXCAwTX9L8YMkHtGHyxDxeTAu64780gK9P5kxn/mB4rrnF1DXHgz
enIcNxVJUZiweEZeMixEzz6bZRuQLa4+wGwQ2Q3aPhM76VV6IlyGi8Xh59ME
KRZcHNsriwAn4WE9oDPO92htK0yO2xL4eV8FpnaUAjjNGoIueIrHJCB6o7Gl
mSOmxeqM48g+an9lsDjswOryRLKcoXwrawJanqWEnQhZBrot49JONhTjDvly
jnG9Ee/mhtEuGIidmGgVjelwnnkfq/gJ4W9AnIYN74asC/lk/Qzko1dIn6Ry
59ebvMFTgmjwASLeYKlipAwN4Zu9bykHq5UKvtjcRuuAEREY+i3qZd2uVvQs
Iw7oheoK4FUr0PdV9LIaBrGeDvdrHVBwSfCt7RomHvAP5nrWaqwwrnIbMlqB
wxRkvhi5yX7wtOQrDB4WKadMYXD5wsZmlXJCCGc06MhCFRVlbSCoiTSrm6rh
nEPE6HotIeGrX/oVCG6Nq/Y1iKHQyODJM4js/b26M+AoHvolfwEvr6Rjc2hl
93AHKFnmz6Hz+yqNez7uriKmiUn0NY2GRligpFnt1QYAOyZI7jqICqTvk1Dy
DuX0agPb9+BCm9BHOBygZiOdhQOWEO6OLQjBpnDSrWrxwVjjZjICtkmIDauv
e6csycju70lvGvaVrPZRv6d8i6pusHaYQUtvc+vgal6ycJ/w2em9ph2KTR1j
fgKFbj8ffqUccg7MtcnCzOG+VxQ91idPGYxjxsGIIdHqQozh8x6zqB312YVo
DBZZ3xF+Y6W8nypoaK0vdtIEnmmxpioLyNRxaHuCoBT1Ho8ia78JFblM9sdI
PsBuc1zSswTAbj+6sAzwCAxDvN/SmHiZninTOA9NCXphCrqHhpDcT28VRyEF
I42CK9H132a36NPVUhVBPvewtftCt6yLOBDUe/feA+BpVr3hvxi/iFqhQgya
R0ubN3q42vN6xTgernFJZKisaiVg+cGRlpgBb6Y3Oz33th0a8uKFHqbjyimT
x8Y/A0lgRrD3R99CJJ4sZuD0MQAFefTf7RooqYQUxx4BMVgGu1W5jwhDdH7E
hLsDzadxIS+SWNA3bmEE8cSZR7C+lCQYIht2jeMuKZspH1LPAG35nlO6BCPf
Wrnb447QCIfDvzh4jFJR3r3cJzqQxh4Y50u72S8JDa3ZyR0wry+jiAmYteWU
4gc6V7jlpB+osuUzMGYCk6wLAsakPB4FeoTL2/t+2D5DBMSnIYtiMETzKpKL
zlqa+XJBhL4S8Z3Qm7ejVKY94c3Nu4Lohmow0YWDvNPuWyqVCoyrr3MZ9V9Q
9dck5hJuzARfhasNONYcjVDXzdGQIfQBK+xUfukhHNSCv4yQi0bVloeRvscy
Zo4+K9BBOigfUI3ChPGLhQCeOOnpcJIeX9948EY1NsmVLObhlSZ5mowutJ63
HIudy6G87o5ZfMDxLVGsWZrpT7Q0VW/uy7rNVIT8/dUypHRmAYDSgnmRFaD7
f+Dnbu8qteGj0sBRKsW7UTehbJORwosYREZWZ0yevJHEOuZyVdfHKGmFjM1F
c613Zx7O3nxdHNFbOv/2q1+kB3ixAi/+xNzpi4dxJpy2n9F2OvmOwcCCHOOm
V/LEcRmsso3mIj8DjXumlGRO6UDRbiia44ystaF76HbwhQ3C3IiY/vfGsSRd
+AAj2NECi0HNdyPcGhejyLBj8eY63XTiaFMRo24EtB8deti8as3HKh1awbBq
P5bxWf0cnIvkeJ8GBqpYyIcRbpEXA5czvCDigqXz48MC/ET1Y9kwEqpBIWqA
4cHYvXYU+Rducmu/+PiW9F3Y+KqPc1dGMLhyVt0zP1Sp99YMVq0HziwyPlVp
UOQXzL0Ps0OGjM2sX2W7uO4DaQS1yDENXrgWwDvWVUuoA3j2X2web++cZ6Ih
5HDSwSJSOIeKSv/D3CvjGmvBUXuJ4uumNMqpPoBKkOMRzcPXzfylKcrjzCfp
A3pHt2tk9JoJEI1wvXzkRP5Ke84fFNqY+8rJxsQHsFx4MbyqSG9ujlmN7js3
7bcGetqYJM90BFbLUHf+MzC8vwxDdk/KoEW9k+4vfQYpNHB+BySfPvnEC9r3
DCGpUq9ALKJIIrzTZWOlBhfZIE2hlAs+Kfnny7nlau2CQkz8tLAR+Am+/piu
AdP4eZhSrQq0/9GMfa9OfzyO9amUXh1OGosTrv8QyCpiTy0ZoS85jQHfUAAJ
j6JUbDR/URd08jGHFk2UKZ25fJwI9fvRzt/mi43iHWjm5EgtbvjjuhcgVUX5
AR3ySyVrTFb4NJixw2D104hLYfZag0BzS/W+n1DVYkuLbqJU0OCdJWtCNarj
DbziHKTljaEBSrXHxcPA1SBG71vVnVeirxu4P8Tr7dQ2XPweGNkh4/5z8P8R
YFoqXhvCj3CVjgSG+Ia3yAnPuWqG8gr5ReBxCCPlQntddLeeh/w0X/8BQIqp
qZwQ5FWDn24s8Ku6QTdDVHGVfVpqVpVggcrAmNUI7yd6r/nN3Rd0JZyXH2nb
tTmSTLDQcAX0zR1uxAVPWw1tB/Hzx4OMIIC99rq96dywvfHLjc9RQ+32iv6I
PPK3L00g686e8Ml1MmlbL12m2KtDk+NixiW9hM7EUa+ai+6buqt+sRiG14em
FUIXOvsiso1bSvFQiezIOoqkoJU71umbeB8pkXqvq6UZkgmDVbY/+8lx2nwz
mT5FjJMTASj9JbetbtARRzUTJY5BIvV4OKUSqPwCublc7KuR9W9031mvxKtG
mscUQeeHSJh7O9/wW3Qi7hdWZfI2KsjDeadwIkv+lSq3UgntbTCMJvBrOpHe
xCzneEOVt3jWz7L0/M2L2uGV0mDagnDL4tUqd9fMbSHj4/H2+cZ1HejBTOnf
kUhwcIAiaApCRTCNJhlShfn4Hw0w5YtKhwPtkJiqJzo6SlZhnkeHVg/poh2/
vFvpXl63yNyoyYlkXtMfnoZa7fM+m5BedqKjwpZvgYbg/a5AIWHjiGhPWdoj
ZCb/EiMEAeTAwXa4xUfxmSYIxrS/8N+KekRUnQ1X6VaMZIC8fHdLHD6+rhZp
VmWW9jPtPj1ofiYYUhK+aawYsiMg3TEqBChHJZN8SWEyWXbgFHPgPE08Nghm
K1icvZbhweGC5JXP2tASelp0qha/70tUASJtCZuxynq41BEKTI8AyIlxQzw2
I9dqqz5gouXyNxGYoty820YWC1q7IoekJMA35a6cc37k2jShVHx9HxLRxlW0
TLVH7v0s7R7e/eXcauCyjyz0i59opyr+pX5PLCXV0g8/iu2oi/1rZGfwVNfz
UKjvVJTVj5g3WUs/GQM1I85saQ/jJqJrdPq+KGrrJSm/Wh4jRb1xRgfr0gWA
joQxp2O0kzyGGf6A1+sPsnd+ATUGTRES6CNy5EX9iMLPy5MmM+pypk5k2jiu
7ZjoPVpnLUVk+ijKpVlce62PHX9oKwV1Mcysw0oQkVxBUz+P1NDF0so/AM3c
zyndy0RzeR6W8t3PNxKtQlpDobMxeFOf6MKQTyrZkxsxEIeovebz4DtZfid0
EC5CdRC9h8YfHM+bnxXGm8fzbpcWy6IRuKXkE5atLwWMWz+w/lYz0XmNNeLX
WdkXyo6s/6flF+sD5nalXIDPO54ORwXdHCYcXnXnXW4q1C7UyLoBjXEqhIt1
Jmovnqquvn4KRjCQilvdI4e877pJIbTij/M3njVltmcNJiRcuUguuXY8zQ/z
jT+ilswfBmZhIGgydnlQXFy3pwC4AVuGYytP8r9C9uLmNRlSEMlclowpTiGA
qYW/YPNf2A7dtrZNzA3lbG/SFTOl523IDCbUgy9CF3hzx6h80Aj30h0uxRGR
dsrEe6wO90AnV+bZlJ59xYNThkBO+5trR0gRVTFbwsei2DdKEbBdcyB+kFP+
yOBQb1pLf1P2rL8dsyfS+EZN1d1HrODzm1tdaR3bXuvttyWCKDLh94GPuYrB
Pjuv7Ek0Pk8Tmb5IJy5XZnwu5F1K4Cll80F48cZ66eyZvV2NLOU32X7hUwYs
8RpFXnS/EuXJegGNaZVCnh9+Eh7v/6WhJXERU0KwvQLt15qKbJlSw0mx2F0C
u/W1h1n7zPOZbEF4ImbrsmtdyIdbITf/2meKzZc1h6yjGEQtlARpo41jrdK0
+LQagWVJQcdDTUEMe655gqFysG4XfqCdXqcGlGcWUFM2bHAHM9KptORwkQWX
EydBgChzAOqF4CBoX80h2z3DbQyfa8X5Kx0XO6R1f5I8GxjwTZAci3Qthqo+
qf+XSESqm6hH+m09LVFRzx3vprHoyBKc5U2x4SKe3xu0oH5AprUSKtrXTupy
bWuec+tCX3FSeeKaJCuwXQV83R9meX5W36MMTyC+Tw8eopYGJmcFWycyRPuI
ISB9Ct44Fc0upjy/B+/N3fy4HiRIyqNFJR2v5Jc195RY2+tdoNgjMcHL1shX
mjZHQJh55IWsegDE75P5/bTF/NGFE8xK8MVBg/76KO7QXO3WkIsoXum1QwFO
1u0PWXG0ZVr+IY4lPFC5gbYe8oyiXVmmv6m1oXFOt4p/mEUsF611o22JexSs
rPyw7sIvI6xu/bvaAoTmdhkmhJ4d/soBW7CEWxk16UE950bv3TiCkDFDRAyK
e7NsRY2YzvXeECTfVHFjNBmWY8FXEOulurfme7b6MXY1JFct9QrXCRZ9vbsG
yYxiEoAbI3BD3MXAtbH48+Qv5vjTfh00FwSTa8S4UdEbaO47LUvxa/1ubzXu
FIhfh/PNZ8qwq3P+7uk+x5sazIqWd4xXkUw8VPG/HhdO4EQkhMnrzmGAlyEJ
5t2QOBTTdah+oUGoRlx5OmasvDJDmUPTeD9iLSoU37Xe6fl3/1hsq6vcPvPD
/BnMJzCH696I8MvvszH/IP4NfdnNCLd627odbOJdBDuI2E9983gEYLnpfNWh
J7tcUezIqR7kkABWunV7sZOYTMHre3kRx0nUCpvmLZmRBjM00Vnpdm9I3byg
ribvbHMTuBBeEiFouLsNifwOxuv9HFl7RPXc+rJ32L0tZxm3JYh8nHPy+6BX
NC7XpXzwxOAYIN8dYc4Oq1hhmD/zmV/bORVUoBx5UagaQ4v6iCYyqc389ASK
XeL+Z4xRB6r5qPi+49jqU4ej6XBJLKutQIeLNTGr8UrYjgVapN52Hd3tF/Ws
yB2D1LtFhHYrZVJptjDffVLw5F41xzo9G252fKrdtOgo8EBKgSnhCIfIzjpQ
PHQcY/4RxRieVDkgJaZm2HHEQFkH1VTh0P0bCzdBlwGiTvE38xmFJHp6bJhG
ilHMet61DTHddgBENTj1t/EExVZBH+e+0Je1Wlsi6JKZz/bFs0kK/Cf1bLlc
SqTJriUEc/Hea4aIpoR14f5+jrpW+P7yOK0fgtSIJPwcRFv63fSQqYfnuwSw
p6tGwqAAtJrt/yiEJN2GK/X3efkAik5BUamUEUk5iB3gSkTPuhOidY5HXFZH
eRXdxwv96/crZmIdP1nSLlU1w3JsEocCujGrRvHnj85KEjJouAjQG+RIoTw8
dT2+Dn9qBFEnhZqSMAab5GNsgTJVrBrEg5lHj+z5aI9PACF9X75F5quCyoTc
w/shftif5rq8VkWQ+qEG3SHk7khiRgBm6YfiPIXBZUq8+LikgjG++MrYju+y
Ck83yzDsfi1qyGIk2l7wflpa6EFQfe6iXShCcraqQ3STZqOFq/7yCIOKL2Ou
zhVrjlIs2zn7vXciMdk0cEAfFuTiBO/SfLPjGDgL/zS48gUh3ZX1PED9C66R
k9S5AxkKJGBe+hSgp4jLeJa5kaoMstGdDPVRyYCh6esaYzCzi22GMYXgoKbG
8JLZaaRZPsC+dUaYfH36wR9kelDxETDTS1clLwD8dMH3erfJRWaAUVDD3Mmt
C5fJ6vh4uMpCgU+iU7kkI6as47zNc1/qIU+Ty+zeY70HC2ym2UyEtLsNvfKM
BWevfo2gwtiaO7yjuJCk/Gx5CV24XXnrJI8pH77JTv7ZGYfhzGLTxSR7w8Lk
I+2T+BEr9GLDXTDuOT78cQYd/r16WKGPjOfcLgNrIG7Sa6IZkXFn+B9GHC+1
NvuBD758J+NtO1T7sGNaPpkPRfBH5Wf+GA3R0KFLDEwP5UQ/00iSC9AITvU7
RagCNcOpgTfr4FpoPLzU35PzL73xtxJmJD+DmDkREzNw4KD2QdAuEpSQicrG
4R1C8AZThKmedB2OGJhFx/5WskLvjxGpC1W8IHBQu9s6GXGxGNr33M56ertY
BsCqutnBi6mj550WkZ35pypqR+HTX7Ogim43dJ7JaEUiD226tRPgWdh6z9Lp
QezMCEZoUeScEYkiqxR7enuLVdUZS7YZWrcmUezU8MvaUeR++QKRyBs/JnxO
2/HSLPrUWb/24UY36HADHQDWbwZsr+t8QMiSM7+q8t9m5J/BBV4UaTcKziSw
QQwq/Wr6tgf9vIw91qiqZm8DBQyJvojF7v3FCWufIiB3vk7XgjY1cYy+TSm4
mLeZavxra+PwIJbz3hzCywA7jOs6HEArqTwerjIxVuntO0aEdCIoNzzxaVcC
zqn8TLVy+kT/KohLPLt9kU0L1mh2Ea9iJaKFSZoK6FZtoequ0tqnwJuSA1Zk
dReOK6FouVmOZR7hXLDzbwRr653jqMDNySYHSkZ8/mDP97VX5nJHefRKpFRy
nBk48O5Y7gdgqUi8vPoUHh9Vlf1/kmKYH8W90bN/nPdBgTBFQJ3Uo37KdLQ6
cLgZJqiGjIgZmB7Mmbpss+PGcY2yy660gVsEEP1itOl1PdfuQ7UHHAOToUNv
lRc3MsET9FKfoOA/BxP2YqRYEB7JZQEwO8fn/f8DeSeudCzDjXOkG6VRWscg
JxJSMdiB24b9i1g9cItc2yLYvwyqw1NRgzMw/FkdZPENS4eQTDrq0LDbgwhz
el0E+ZnOkOU6sMX1aJVSPUf7V77zob+n9JSLm1xHVi/oZMNEnNkEqP1eTCnR
EOZCATWgtMdLrd+rho8EOTfECz/9SPhWrIklHjovnYlzCmYqO+SrkZqRWqei
5h53T2jMAwJYHiUt0s7dpY7CWT6d5PwoTsQH67Sz6R28/Cuauy4i5Q+PaAwQ
H/9RX8h0RY0PwPf4oeA/qnLNbnAtrr7cl7gb9s6m3yY3w6jeraYu9EOeyAx/
XRIZetL+7bb5AEjNdAY3fUPVUkoxADgRstqlIiupCJN/3lBUavtFM6Oiq3IA
2FHmLtJNIOW9ypqJK57ZFQ3+Vy/gH63x10aIBkFRdUTj+h28OSveG3XSDtZN
wGRswOrW5U05GfAWAwFz+01scQwxxv8TtW+lqQuVoE5btsxobSbs/nZ9d2YW
u1RI6z7u9DBIGlXUdiUeGcFZ+umNdWwz5qBZ6DROgtoF1dR1gYX2I7QH/IaO
cavkS+HZII4lXHfjAdju3vgxiLSRcwGRx+rZxLcTXTdgKY0R/DOzKhGmyjAV
4Ff1enEuWev4S9cPzLTT+FH++XeFnJthbKmoa0LBB/jzyy1uZXr5L1g4ezgS
88c/lnPMbFdX4t7nCxEyAdKQB2AHg6Ogt8qqJ/YPDpUvQaE/+Sp+qU9YEzRh
sw91eWP3DXxbNj3lyUtyklu2O++So75jIS69zv+iYDTdGkmGtz1I3WFtLJAi
3NzVY+cOZvlGNBVy5FTrQpenKUnF4Nu3Fkbc5IKA+DisW9A7SZl2Y0SW+kMQ
Ofj4RTdh/K/0qVsGdIhqHDtaT5auJFXNGRCU7bLuOoPsFcjefyrho812hRX5
99PTWzrgNHmArDIst7kRg2nMvxRhHKyKvbOyZIulhDonnrjv45JepvNKa6AF
H8Em6grv5mXl71vBnOeVwWvxCgrI2oRKbPiuRG4lpTU13uzLg+mrS1acuHM0
r5kiIfE7juES9dtZYsSZhnIBz4OMO+bO6FE6o2MugKrpdE77NbjlZyySFmMm
VFcevPF7DQvwVPmk014VIlbTizhhNssycM9enIJ9zEDW0Ljud0Q3V5iL5WmH
R39xSzAIvjJ0dncoSKycwek5mpwhsQ0SwkQ9DQqdwd8Ki5JVwnY/gEnTtH4p
pVLXQS+lhrf4oRGEDHKB1dXBtNbxmQ0fzyl3IfkplDcNMbJLjbJgWycr5L4c
gI9m3BxDsG8IlYaMn/JFeAf+pdAwBni45jNwxFCyJHaztxzJuy0mByWBFfq7
b3tw3zYRECtzmtiVJr9w0v/WGY2QKf9bgs0S+W1P+xPGaf8wLSgZsKNrOgKG
PKYN6lT5TS64ndm+O6sY91d7lj3bSiWmgSzd4Jq2kvgKpGDVf3wj1/eS5c2U
IxRNNTK5CeXTGvt52ZYllzMXwVjR/qx53jYXKLtbAKrT9GGv9stAcF+4sYcV
0QHITluuAmDI7ZwnyQFNGlKMQfsXJ533hwjEtz1PH+t0Mm9L45x/ISGvP0PT
o5IsGRe12TZE5cIxjfhosMcTLI7OxYRCUJUOSbyC+DSlHh88sS5c0Jp5A0bR
0L2AeOO7aCPjE/6WwAr5WOl6oIBD6MJdZAaaTx38WGPJ2SyrcYBHeExlmfi3
1l7dTLDQIChRrOGBlO9j6ZEo60ePlPlZrqFRL01vJGRiav6eCoSlFEdm3QAW
8BP5JyUhfuIBOKZxcSfJ9LGxLvVu2RVbMvtuOwGA2nj4E83tS0KSmcBsmk8L
gO59jmAai1cSldUT0xydcbpuyTbK+uWIoVFMi3OdA98NwhhzwaIdy9R2DWMn
tqb5k72/B1Rdu1KZ84O4pD6Cb+AYv+pgqX8IrEOrXjbnJQIEirU1390BJewv
v9wbXricroU0pCeQTA8iBHipBo/JE71+y0nbvZDI5p+WIcGFHvFpSgErvajR
KfSYJ1ORfjb7Q6lcjWGQojTGIrpVhnVpzpzQTKo7XgHb41rpoil3RIFhZBff
hZWONIlUFPK+FEHZkLT56pi5+R5kFZHjuurf2islJ16Se0FqT+zjxZqo3VsF
0CiA2rpY+kBcU6OWE/vXZGIFJNE79tuS7zJF7YoYB25UxZEKvAo6xgxdyRCZ
x+hYBRMERZkxrJrW8Sc2fu7QxORd2zQram6HXrx4MWL05oEy1sGtQGYEOvZc
/OnzbR/1oQhXRMyeVxTNBfOLyvxoWML1nlvKd4rQflLpcs1bu15onDpcu3rw
zFAt4U7IqH+kNWetNBfdVRz1I6djlHqx+uUX+fTYXexUCDDqqzVmhD9PEYGl
bUG8CVPRcqZvDWHt1JgstaIK2T6jBD5qLsInTl+R8LFT0mEkY95VJyqRblJa
rekmL84Z4ji4sHn97R9NZXZS+BKuB36/xhgVI14meEJVXoVAQA1weNXb0E2B
YNbwiNTsoBtfeZRgBrHx44BO/WlqHgMslFKOGa/HibR2z+4JqRz2cks69Yoo
UpQKSF5prDVAbwGnCoPw4bzUVtAHUzCxWgkMmDKdjwUmSV+eevfY5Ph3gOlg
w124vlEOk3pAXlMdyJG+q1xwT5P9L7MGcjUWrsTS/0icXWR3pCDiKzLaffie
c110mHEPvS3pf5hkwrLWLHDHyS6KOe0ygZRXBVTBrbF50XClN7tej51PlV7c
NGWMH2iQbraoVqbNrphXCBg4/XubKqtHfBvgHIT8ecMc/8AKtkPe8BioGGtQ
ddJFDHzP/q31XoBg5X3W8ieE5U+g5RT8dBwUmY2KMA5/H0gv5BZndqNxUYXf
wBlSEDf7fzJJ+cYi4H2hYmVOF8awQLuEl7fhqgRUCPSdicNiIuC4d9Pd8rcb
LsZcBmU5IngjFL3+cT6rZ7nEB+dwRLg4pldDLOq0o3vD2TduwYxWcc6DIjiN
EnKtI+cVd53+IoA0oDVb2QpYFYG1FAOI03j7FooWfJakpm8YKBNmY3UZah5w
V1QYGBYxNW8Ri9L21ozOs6PcQTVhKOkS8YES5gUjbpqi+uDuWqh5LThsb0KF
JMLSHR621OdmT6/j8butjVWn6Y6LAmJhFlp+QgK3VsPTV7XqV3dvtr6XrQ7F
Iiov9v7/Jz2vDqmA79RuHpQa/NVkr2WF/6g5M69tJbMoo/8I+DmMDfpCz96s
c+I3w6x1ZJzSwlTcgz8biGJAb1Zhl3yt2q9FGb2n/gREVfa2d6CD2jBCe59a
zNPbfW0FAOE2xbpfARakZ7I63crLc3IiLL1N0SLfOMJb6I7Qs+jeRByQormL
aYWPFgQ2gxNMBQTRY0UB1cBmo9sfgz9UXNLje7h7V69jhY5ONXxTREWq0OQA
CPksPgRLQoVz5t3TbhAdAKUMfMJI460FO4FkfWBMsygi/PshJYHObH5tBbP2
kudaGOAO0Yi5K5IPfyhS29Zutqe1uv7SoXxHd8hjIAUBT910G8mE4ocDp4+c
OUSKP4YnnOaGJxwIN7hqQ8XuIGGFJKNvLzdBlhXxaAXrJthPKfGOor8TJXr1
Q5umOKLKx2wAJ9dZLqqLMhmgyJe/0JFuWSLwR/7v+KFrocgNg/++nveaLf00
JNM+O5YwdtxeK++QwOL8qcTnIIzeoPJBghm72Q6+kgshkIMhaVgKRFGCWP2d
Wv9TP52tbOEi+dPQNn09/S3cHxqGvAdnEH2uXzK3JfnLr+4RRgXhM1MPLzB2
jqdy1i+b1JyyU/Rgbhkh327R2l0CLM2p22piwZWtb8sE611uGTfdh4h/GMCz
JAcbl/Urqt474miHbAWGEiuX77CLW2cfQZHYmD0a/r04P0bsdajrf7YB26YT
4WRmebEOhwQdJleGNgstwexXiqJ5q9ScCcL9SYCoWHqvFt/azLtwYbjZKrRi
hllnbo1V5QArjC2LcusBaBxLUqtenHXYb4IA6WVpTkuxTYlK9WnyNGv6AmeU
DsCKxf4pdLmWiTLnGLY95F5vca2nGlGT67cacwBmxEprg7MD3UHgbGTzuiKC
8W7aQ2nMrCH3VYbYOnrg2vTJadWxkOUpiqzyVXILAHozxie5/Z7mtT4MzZEr
R8TjzI7kgem0ve682OhuSr407KsT0xAREnm9SV5QZcHHGSccc36SUraENto1
DlMMs7IGVhe/72A1a73rkUkF8pBN6jUmBACvU37F8BMnR1gjQeJtwOthEXM5
h3+PA+012aJ5lTaXVprIyfkTwGTADkxObc2Ck7lIx2b/EqLQIXmi/oYObhEo
Fgo3el1eb3QIW4nqOmqAbfUqqUBnJ0c237Ybnmz7+P7jdV7tx2FCO006IYn+
skkSWajHzmYKHvqY2OxKz2iZfycMqIgjn3UeSFk0Y24MIj/in+Olo2EJi9gC
o1C65IiOloLGDbMjk9h1vlCcl0+kFIC7qacpsjxzksqqkM+Dm33zt4l/CqgD
e8nq/TD3lzlVTmys+A4aR8jmJAMfR0y1oI95PDzIydX9g4vyDXZ1MTekqLsc
h5zHBlIXPmrA3Ru0tFGwO8FYNdeIkGCS8h0ZYXgpeaX5/Itx69AV9ojtsYbZ
eE1USSapmfpfIt1v0zr5yo6Wg+DZLmyEI+5NboYjY1Mr2dbeybD1Spp4wl+l
3ZB8TNixUctAZu2Shsb+ARrZX28udcfz4mjUYr6NM5eVI5jvVvN/IHQUUR/Q
RiP/6t9LCW+r5Ok7h48LivwrBc7SFifQL+DhIfK5zACz+T1FF93fttUfXidy
/K7cokIxWeHbqvPaenfs/ZzjPKjEYeY+IhroYoNVOdkv/Ad4ihfNB+Aex0Xz
k1qX7UvaYSmjC1x5GLajlevOYhXA1+4CPJOE8YMBfZEXODhIq1MTSOOadLES
yAv95y50TspcJh2wn+KccO39X7THCfQ1npz/hGIFiHqmnBywTeEX4XF8ugwi
BqU8zPkUR3A6ZgOkU5vgd4XssvLd4NVuJNp5epEG0Ls1imz5sxcQ0dKpaFE7
g9beKQnzmZVdqglB/LslClLi0T2Qfx3IDnB2vqyb4VSwTIvvO4zZWznWYI0Q
5I9ngAM7T9g1DHl81MKACE8Cf8BYFcyv6O7M62kkIpFyEQOFBp47gOBc0iDa
EZhY0LDYfQO2CKqvx+raAyLdtmqPqlX7rae9GBbOkevcXwfUux6Y4v+cJ2sU
BKws0ks9laKdGdDhawlJxORMFhpFj7J6aywObmwJPUOQWCNEJkENjIWRsOgs
CZpIspacpJuw5EplrPgmUmS5tSdC2wNDmLKvnYnyKx0T+budVNscKmaP/dj1
6IgZ8RHSBZhYUCCoPcRX/8n7YE+bT37Ywh/3gbknecrXQ4KXUbtI10Xhn5Zv
sS77hwtRYAA4VmnnI8C89GRbqN3x12K4amUY6ROVuEb2q8Web6e+0vHOw3O1
1GQhrKEegKe1JLmEIBcZI1xDu3XjapZmCfDBW7eZsUIERq2REl21PW/hgplE
BoEXy4hJUa+bD3kpBsvLNk+JhwTXXQfHCn6j1v3ugqm6LWL1ixpdbVn3vbFU
Y8IFOO1MQbOpMLJUGK/sJBI3Aooz9QkykH0tYbYJJulJ0SLarm6pOSGlzZUE
XI5pjg+QEfk8OAo9qDyatO9eeh/q2ThE8KfAlbVPyyceXkykIpU2f73/WY5H
gHDbSR6drutr+LvGwt8qoJJXAOUfnWe6Mh1YPvl43DHydA+rCkVY0hWFFQs9
IqzE6xlkJGAxcU+E+rbYSK7B3QZPtnwWzTlL7Qrfgh6ajDTsfIGXsIcWXz6h
6OZSkhi2lyjAtxcsx4Com51gKxMplVc38ZR5foFGWZoEEzA8z7NLNBW4Lcnv
dzHAq7JkJ5n0KXSIhXOwh1za2DisqMFtt/tyt89DY6I2glvawaZlE0OA8Ti/
sen+5L8ov246tU7ISnj2yIA3/NP9rzUcxWNiyhrr28/IJ8UbR0DGXsir9s+6
EY5IBAsIdPt3CbCsZwm5GOkzpfK+6tr9mpnEtvYV8P/idMVAc/E9LGgen7mN
oVwR2T2IBgFytJNkkE3yaKmL3DkjAP4pOS094YQRrltu4ba8vyTdqBArcbfh
O2GLXCwckF8Q/7BmEMSSKXaMhE1TeH7AaGyle8Q1ykU/EpaEL1qKjT49HHPL
N4fYdch3aOXyv1hquQXzoSlN0+ermlo0t01GoPU7AcbX/9rQV6UwpYcdKGXZ
Li0hollOngBibGGyKJCUH31LzUU1PFFn2IJE6OYxKW5kmCwA3KmbBUo4r04e
6SlZxWlqLZjOcbofgs+NRrWuglJJ8e/Ik+gWVvyJMyByVa3LC3IlGW3pjzcd
vjG5vZJzQYdFzTm80idHILCjwQFkHI3bYSSul/Y3gJH4TWoHTg8cBSRX5FOs
dTP+zr5ZArlbKmwwsF7o09P+8iMtL9thAFq3e4qan0s5W10l14yyrEHoskSz
mkZJYJ+7vW7MSoegGJEWLaXJOWluWIBY7dhS10nq9Z/5EIMd5SqvFPiWsc/8
eKkK2AbAHk4Z6p5eS/9l+8yvnH1OZoFG3PnPd9hpnCM6N4+se0XRaJ/E+tHV
LmfiZhFlCCNr6x4XRvYZNe5sfatkJ9ytTUzggkcHAU2R4X8DgUYv+Hy37KBA
Pc7P8yfeyWlVLw5uTrY/51AShkZtMpnhjsM9NAspGiKnB3jaZ07bscs7zrHq
vktpcrwKZIZs7Nnf/VNepPjVYSJwJq/UYJ407Fpp9aNZ+W/O379igyEu2jOB
fFORCvqRIyFhLnp2as6qXf7ICcxCmiXuAB2fXKhoaXmN6XDocMJ17hgPd+Zd
cmMPZ6zjX8tbFdQgUeMtdXPsYa+8P7ixa9LeG9xfw8tYygG9W/fF0cfzARij
mPepm2WBHm1JGvV5Z+A25bZav2zEyDS6ZWwzK+ez+xDBqSRwkduu9Xe7Uct7
A/I8fpE7p+UNhHX/lijJDg+J35r517h6PyCdNPxrUymd0GcxEMBb9ddgXgoT
VJWpwpQZFdwIK6nkH4w8UtWTXfT4EcA3viodkapMWIvaDc4SrtugBW9oCUSG
Vt1A8G5v1mQ9z+b5AuwtPm4uMYkoGfJhf9i09Rgj+IQ4v/DfTxPjkgIv9g8H
6FhE5XdChZx0zE/tKeylYAB/oLRKtOEgbJxSHk4TwRS5ZTTnA+dXC9ai6Pv7
5MTXfzJ00rzntzn8PphumAk1PFMD/9vY/3QFIDn7B/QEDcXgHADqHM4oK8Iw
xFDouzJA8TNUFRgh9n6mNg0gMxw5Vrn9ejnXc+6Z5/RclVPTJBu0mAjFcknm
7fiUZey2jNVymbUvcf/Mvuxa2P1hg0hIkR4mLom7YU1VqU3ziU1Xz9UfhOvP
CiA+HoJ9ytsMs0mNqE6OWQ+ds5dHOG4xfvR1agDVXExAE4ENwtNBm0ZfnpoX
JjmpFsX7dYWC7/tu0tl3m0761Ej6pJiUuR1cyJImXmt/ecAbCx2CcvgWKG2x
rFXe9Xyt9bEp+MXh+qZNGJbaJiVUuT/q7OrgkfJx03I+a/gOm9U5XJTFPM79
PmvS2Eut0v1g5m3LKU+WoYpzk2fpl5ioVTq6RL3D9B6GYGskvjRNnTBVcaPb
fw5z2oliw9RkJGyeA2tyfTLxxV3RDy3GY/z/eabPS3SETbscjNbEjg/cMN0E
Sy9tVDhSaKt4Ylr++kkT+bzUJpWQ0w5PKsifRntRV73tlYd/w2kBGHnSDvCC
8KWrTUfcLxincMCFtI1EK2gXdSyxWK0LKWEvGo7FmeeRZlL4nbZiqdBy/D0K
urwtJtIQ6kiGbo3LYgkrMk5tPvSsd2QRapN+7lBELU2XeHyaBS3OhT5i90MP
MxhQmljfha+sdb+MnSTDAkFs8ZjSUDb9qLc+phqIgWLYN1onCb6p06AZh90b
x/MqOjxJuypc6dIdw1FH2cN7Lh5N5KLlf8hfLdUt8VjMo4fm3deVWRmKqWem
WZA0P8FiKuEe4P+/dhwnrufhQmt61K4l5M6vxIPNzff1/EYPvIrSSyj9qcUj
OnHJoV9+v+RDXlFcCKmDmLp+hs8bNw9MYSdVwQ3DSP2+PxassT1qE69RMafW
7rwb2ecZP6iIaisa0kXdjvbFEtQtzY/J/pC/z2K07RQmTuKBXhmArWuCo16L
tnIi/hFYb/GPVCjRWaXL8ZEkzp6u1Y4cUK73gsEsdE5pzdA7tBMZqUOwJsvG
sBgxCY4ojOHgDqc1q2wtl9TzEykScdQbeqC/xfRm6lPdEedJzjWfiiZZLsMB
uSCl/uHr7V2rS4fSXcmS2qwU/fllOPAC/CCemmGas/Cp6Cdy3qvBCtWQ2288
RxYyEPlzTWh+F3MStK6C4tAZ8pcRIrAa6Kz5IphS6GicgoKn0NZzhbcZy99m
OxQrlb2A8YsdHUGmfNdtiaAVPTdja5mThvyaLB1qZXVhq9HCcszs0apTVq6U
5Y4SqV82GRODrGLtZ5x/Nd4AZwM0fDe2BOX0vEmRs9eD15ae1awnKsVwcYJc
D9tsu5ZEAXxLNPbc0UvmE9JQMfcWcxyrcCvRdE4/+8+QX+mO/r2IeMpmYwEy
cRW2EJ9VJBVyfjaRZCyidTTw7UpJLD05h5CPLoYtCyKmH021v05vcaqdKebN
1TZ8XaNyCt5gMwwGcM2tP285aN+a0emQJGnY8Uj2Ovo2BUzlZ/lBdVRcQJLc
7yh+FQ//r0PLERQEbtZ7xvQ2+tnaZNQre0OPud0iOdSFrqgcT77guyO4M/mf
duNwQ6NFmn2cLo/ez2MwdfELwoD4+/RVQwf/xbiCUMsESrm5IvATUwk07rdW
x/HQcyz9X6VSfncDVpJO32AU7Up7StI2UMgVEI4E7Biy+kHZtt7K8hUGpjKv
HckcFvNK938PVUtGRpX+HjIEgk6WfKm94HV7dLPKCsvCL8b6L+rOWUs9IqBU
ZhyX/ML6qg76D/zAhm5k/9RzB4Iv+mjGhgBvoQwirQkHa7t839adocUEhp6A
B0ItJ8tLkElJLyf2zBmqQQqK6eBUUT+7rr4a6MqxQn69co7IxkozQNffn4b1
RZhOCvc7lf0sSrUTC09ChgLM2axt+NimGHgGSSZ9qwxR5qCLbhtb42nwuh2l
OGh4Xvkqycz7o6Fty6ODgWKNW12/WkQ+o+/61y21Ia0N/jn5asS+c0QnK2o/
xu+bKtlfqxJwlwxwc86DRoG8uNdcvbbfi83BP3NiKS1TnFgk5GzdtL+LtRYW
5Hu0Tqq1jW6+52lKLLYBuZ8UNnblAb5/19yfx/KCX17Hh+BATFl9fYnDahJg
zGmXkIS7/fB9enyJQymGa/kFbs8sF3lFchhcm4TLlP3BtyKMUTk5HwNvA8hv
QVTA3TmKKZH+avgkvlUzvgmGcbl83uB6XyZ2pmZyAgFi5+d398roaR9XMtqq
Ox/rTnKj3kEQMIJJKAGdH3RlJ3HRzljSrIxsZunwW9fjPdp1m26TTp2oEBdR
2VQXEd9dvt8IgDufRLdDzUtgFchroeegKLxVBsJEb98d7wI19rGV6TNH7vYk
LVCFM/Ov1I4zh8k/1nDC7IepOteUTPEdzW+Kt4VFgDSXaIF0TYnyKUXl2ZrO
CMvjEmDQa91+GldpqlOlNKdgsqOKqwdYsvtuMF0u/ZEi2+ZrUnNZHmcv5NnU
vjePnABNzEWFQkR6Kefz2Az6pqXsx7oS4TW5xXpL5aqRYNujeGBF+DY3Qt1V
CNceZh4UNNGdMGaQtc2u3d+USYk3ekoKD26bKygwiV0wx3vt1btYDX7haJsL
Ojf14yFRDXqtW6AxwnwNY/rkw+PEst1UOIUzTWqa7QqGjlOkSlJXmBirmXo8
IynekjTMUGWseC7AQDJrJhPeQp8A/KycDKOs9v8L1DzYIpbi2hhfr7VK1OF7
nNWw02nH1f/QW1UTX/RkJf0Mlq1eoBmwiseevsPoHeuEIwjntu5cxIh2LvAm
qZJ4oh0mZSUdbCgYQZbCVh9y93QlCbtJyswZz8I/psCxzjXg8QwUAyWHJ/8d
JRFuhZhVLikbGY2gM/aC541311Mns/SFpHB6tOoIKFyiioS7ubyq6JA8JmCT
1WeVXU3LljJWxIqC35fK6KZMdARs9CrmFFkRwOT/eeLRlQZCUyql3+liY2eJ
xWoV24ExRI288ZcEbsgdM4V9TQzZPaTXYaq8OctwKdlQv/UKL4RHyynvkSmv
d4jkfjbO/FHHtsuT3GMZ/e01t6pMs+t43yJCIpF3SYv74hsTdW6VRuPC5vQ7
+QIUcCmc8yevPxd26hT7DvPz/m3WEzwXVbzL3ART/dOmuQEQP4+f4lapsaIh
aJqa4nucBjK41+XwCNHmdSvSOb4dqMVRgH7BZ4QxeUVN0VK0/TJCjGLXEGBX
qLVNTzlCnmzcYNg7m93LhLcprIQkjALGxK9IT9YLlI7nsZ69qmPEcwhetlk/
I+4Uacqcu3zSLGakIBp34hiqr3YPprkbFKdi8kS1ambdB2NNzrwF5+2vONOp
vnHjedE2lNcmz627kAysJDDK84LoRNbWhX+q6CUP5RzMycXefCwcDRFsU9YU
xvLtffO91a4PLFwcQErQ2WEjsrSrgdluTozs6jnS4VCbKunylNuwCJyZ2AH+
3xRYwolBvX0aIY0zXvzQvSexGFrs1ar5znr493/bMYDrrlbZ0+4BibwRIvlO
xqzMIjoSFjDDC5J5QrCHXDpKGSZYZ+sI4XupuNxR+/jvfuLTF40oTgOMvS7M
yIyt0DbTLdMbVEou0SR4P4cJ+dPn1XZNi2whMyvNJU+jPtqpjC9QRuTxm+PJ
R4xcikJZ+DF91SOVEUBkjcmaKdiqYd1bD2cE9Gt0mRgceZ3WsEdJ5h+LRWNV
rwlUd5t0IjRQCdn5zArX61weteZsfPfl9RdFvyInXHuY/kRH+5byjEZWBNV1
r28VnzPNh78wMpclfCaSag/tuwJ/knWX5EMw88rW6BwuXs7Xpf8mYwl59uS0
kmWXKbZ+h3aQaDk2WPmZhkZ0241ZD/bNp1ajZ7XEPa/THQhHSv44llMjsniQ
4k46/Pa2SsWFjWwhEgfvKLWHd4FUqrpjJle2vzwZWlQXrR604Pfgy1aOgvCg
Eu9VxcEhaT+yqct+nBdBT3G0L3PqGL9NYqX++x2zhtpnevl977fzfn7qXuBT
SLRX6hSWIPm/EwGt8p+JWrzOIpkDaLBDWOtq1I6qnM0FIQjvpvDt4wckZCAq
Sta8XJGh0qM3EEUvp3XgctvXVVFid8BYIpwmvMUh7cQEu0tuJdVVyS71amxr
WDSvYwhVnpMmwkWi7tOhp5rC12h2R5O3/GJCPE1vmzlJLMx5mHPp/egEbeCv
RZvDgQeWw7lZ6nxDnTnu5MLlS5XkZ5oQ4mca7KJg/st4yyBQJMQ92Yv5+WCq
SVJFZ02lKZl9cATlewNm8JrPQjFBdbkIfdY50HST7BW87iDhVUDiUQa58Gyp
IR3RHooWkkDwadxAm0zjFtoZB97VBvi4RExT0d7Ug4zR4BfeVyEwslKCaQ5M
xvdPTzTUWuUfXrNrjb8n7U7uFlo1OuMo0Wi2IEszthbvH5Ye/Wf2sABQHsYE
0Io9CoumFMB1dOwqlTW9eGglxG7W9ADjeCCIhx8XjINoa+Ye20stEXpUf6m8
RGIMaM03DW3Z7vMfWjWCnYLeFGouFpJrnN0mQk1lDQTJDP+5nA9U2JTdQQ1w
KMmztfmAjtRXqHVY44byqGjNfeiIJEQoeQhOO9Fn59ymCsoV7URGBobx0pDU
ZXS1KVyU4OnlJkGh6x5uEAWzF9kJWWBFIiceh/cRJU6uA+b++9SA1/09QYVn
lOJ4yTMiIp2ik/6f9V3hO5JpeTkWsfNfctA0kwDmdO4CiHoCjo1/RQyn2VTL
8WeZgv5cpfqm2u1vSqiAHKIQIqEkVp9LcTeQQ0MiIccFH36tj/UWKSbw+Bi4
0x15gTXjy5b1Zz76O4zGjGatuXy3Ryiqwnu2AHC0GuDDlngHCl6zmacFdZTE
2ubJPHTjueXHLkh+Hu3PWSDBwb5DUZslu6qdLRGLYIvscPngMy8L8+v6vNvO
HqeONBwnjTwP2Py/xvI7rM28iJHlC9TjDRWWUVR1hvK7rEKgRIu04AAcDIzj
YIOWj+mcPmAxcS5WzFmZVAFWeBh4YaQ16EwEHaTH6pKr4wb3sa+kudkSTXLK
IqCP9GwwNd929g9V+iTLJFRbSlDQp0sdZCFiFrEqPuI0/cXuKDrtf74pvRNL
H4jqPvHmxfl71vPALUNyvJZdekMyV58NSaTDcZjY/MAYzUqZA5eDrfbPz+Gs
DfKCLcr/gW+1R6sU2U7ZZFeKDbuQRWdNQI1LSyII9rY4dIju19pmErZYmDoS
Mli06AoPq7nIHEquLgUdEoGfmay4sO/ZXTmqs34yZ6SBpcVnsnMT7SCPRGLl
wAUcCLRdX/kKei5mnkQEMQ/N+i9XE3ETAoy5NvpFdNrxnyQtsgZ75r+mndc8
i69lS4Sd8DL6p5fkkrF1Fk6NYcqRKaSt9wA2Qv82KdSSYQfFE4sExlreJLZ/
7cuIDsoZj1XDapcuTpL6dnKiu3qNtcY8JnLrfqL2ccjdEx7r5Z9neIBRMXCI
Gfa7xmPGTde04o5HvcqZbvmnBFkYfU1CYTDWkkabqWU1tl+IcdciuLRkcwKp
LZSL9zXz3jAz5H1VxsXDKb7urQ3sVTyAKw16VYLniPjGriAflyodnC7jkP1Y
L01xBY992ql4y2G2DazLQuX/DQBFFsEpdQ0Ic6p8U04ratF2z6CdJLteues/
3LbbwkE20xkJPGxRdSJRy3A6DuZHUVzfkSDgPTg9PwrvyfKBOviI5kFQn5t0
asa1zVYkNjzvTCRinPriR2DQOxTu4F1gC1n+Sef6shCdAcrCevwK/OK1hDxI
c/gGLszDQ5F9dymEOVD0um9MgIQC9u1bZsfZ1yRK2+1eY4kYnjbuvBqHYjs+
Z5s8hSw7jzIM9iag1mWmihT794aNmwjnz9WNb2CdkgBlZ7+iHralKvKLtTly
6DfsV9n21L9hx4HsPrsgEgxu8uYXzrL1+N/rP1yyuYZZj9oxRuScRRYf4Z6m
1towO6aAY6RFLNZvKhleKOtT9BGUj/CHCxQoehwJlj1t3F9qg6dbOINoRp7c
8k/sN/8C4anp40I1O98wLjWrNu1ylP3UyuubrsSQXjuzFneVM+WhF9L4iZpl
9MEn2qxhYta6GIHbTFBifl6e0mJmrrmn0KS1CLCELqes6WoBce83xwfOf+sq
DkqIzMof0NR2fwdqoyVhaAkBKfcOC9hlxn8pPpKRNM020SCGHCPRNVv1fyAz
QdpYT85BWuzRTEYv3fqrjj3vHV9jCOqWkguBb4Gs/4gfOuWvoaUp1bH4i3hh
gj/vjTVMmAqc3H+USwC4912zMlP49ICbT5GOTSUCH9XEt6hsK5JRgCezW0Ts
ecACuL+0qQL+CKR6ZA9IUIS0KeDcyPtJFlxn3ULwZWi6hp+jIfBDzgxmJCwy
x05BdcuK2cWjotTnUcZu3CXb2V5BV9LAxp+G3KryqfrT0hmoS4HSt/ujXugP
nUwV01+5+EgtRYfr3VMRDr99mX3+UgZh31EJms8dRkuuJYmjD4wkkIw9gl1a
5P0nPF9Zoxgfa/++cbKhz26dfD0f5wcJCHvMxykcqbIBwe/49DclBlMhTPaS
5IR6fvLJLPDwOX1UlVr/+v7yiyPnGc6JW1AufBU/fsgasVMzjAslx6r6WzAh
LjI3+T8yBqTDTaqvG2ZRAzYMEHMOXq/DZUH8nL4JTwaOQwph7vlRDWwGfrBm
zAOj0MnOS3OIJ50FAx/E7/LHBTfh63hNg5p499iGojeertpXsR7UUj4IK/sY
3fRvghSMKBSww5oesUe6OnnwyJw5Zk230bCivMZAB0lYlHLCENiRdq+QQ+ZA
Fpcgv+5XDFuS8DA1NtZhOlG0iyub6IS8UiPQMiJCg82qhZGgcE/CmFrgMy6F
+rKE8bPGQZeLKUKZGQOZNHgKKH3SQcOtWWbeebT4LvbPgln1PCjZ61hPj9aE
xCj9IyxacN4OaSTMAYrM97q/uvEeaXiZYe5SQTQ/bMmQTlhXLBYpMzN0Ri80
1DHDO03Z4SVpY/8GXQ20AxRo1XHd8A8fbLAYasKPvNp+3T7Uke882XQc/VgO
QdsB5MWeYQ6IH4FZ/VINDr2ubFJjwY3FWnrJgm4DVjAQZKoI0G/w50MAJmMt
8eHNZAm/PJzgTpyCVOVPDco9qR8EgfMiX5l1HG6NyBxLn2IIWnkT6r/fldHy
/wmkQS52N2qNESbAfuupvbukSJyMWpsnY8uRVBz23NQcdf2ww7G//RQvE7Ee
ZyKd9MuaIBvPgeyX9Lrf1AoEOSoK4vqzCC7sZQ/W1vHF5fo8EgOr7iXQ64X6
oNpelnPsybuMXH+hTXjiJGUHrDow6UXUIghkht8wBPcAve77jiYT/DeaJ5X5
yAj1KWQHB21koGKtk+7967diADR69lNVfywYW/bnfrrNxgfXlmpYPNn7ErxR
a+CrfIA3tHEr+6BwhMYkdkutszwLAm/G/KJpGlBR/Y4aKHsqBI1yMNjNnCmj
91zb+fUZcz5ejtSTwQq4boGwhEcDUAbdftOmGGY9JFgDe5SfdolEfyFvtEG/
ZdzH6ls460mPPZQdFSh2B9RzI7FvDqvZ6e+L9/MmieDGaqTLitFy/C+YWX+q
gJ9/vYErqm9TkTFkxCYn+jOSvca4uAD/M8LT/H5EqdE4AjIU5+SpXu02+Qzp
6L9a9aXCKF4w6syFc6Qvmo9Brbi4K0IMABhkLVQmopnhbt/C3hs6+h/4+Sf3
JWkuHV3iOWmshswAb1PgW1ZdLBpuNhPZmZJ+8RVwb47hyQGIqgsEWTSirwr+
LEMMTPeArnKWJevBrA3CHwAPV7sBEJmu6LYE8Zhwk4hyCssWjYFmAHHDmcfK
PcSuATqc8I7DaevQKafi5imkqRu/eGcHDWEVLn551L0/bYDckITRaPkHSFIu
yici3Td6IiNWQ8MdeyoMT4Kn/CqyxsqYOyeH+1R5dXCOPsngy3ARORxtkQeU
jZHYGif6zWE96gkrYPj0n/kYcuEy5WbsgCeggsbPeqcRHCiZicnIkthz+yJC
RPwrnJdGnHUpqTg6BrMusYR4r46M0sh3BGp6yIQP6X86ECXGVmn9jDNIepkr
/hXlYuC9uZqnbdwP0QyJ/VwklWRAhnDEFxYBo9Y1N8nmL2TRXRGxkgXq6yDl
sP2bfZ6iYLjOa+8pmdfVBDY+SW0skeaG4dC+g51TETa9Gj6DGDu5OpxtdBU3
3OLd7iqjlqbAjW40fVNql0h+cu81N9m7+SRwODUjp0O9WNglH9emBcrGQXHw
L9xOySQXk6d13u6o1DCRcBHsiikZtyatY78DjWcBUGV264vgN2wDzmFrMPZV
rErmfxhZqfnlfdVODcbu0ntb+sHgeIIVzbHNFp3f6HUlDGXNOmmMwq89vVWu
Yz12RokOHLN4KGEWWKrdgRd4DVXxzffTFDSF27cTU1brzAaq3uOlDdFyM0ap
hOZaZJR4p7HYXwum2iiKcmDrLmUtqKi1UwRVN3TsZy575dzcignWNpOywvLI
c8HgEId2gPR8jrund/8snHmqVlA2BzS6lP+nPhw3YyV4BKxw4QkcgKIJ/pca
XT4B/e6dP6B50mKBKhAEzaYLZsybtiwPypIeemqDdBKuFzAoYHnSbGqbItq3
lxqDC5c0f5otLSXXBdh/K9uBfCzL8t7gFIeicpTwlOvupQEIDdHPOpi4g64r
errZ3YmxEAaf/aTdL7zLdihfFlWe/HQzsGQbqhK9d/+8sg0M+wH31gNKgyAk
c3f85vp5gWvTvPGTQHx0W8t+2Tkql7jugC18E1mphlTBBbVR17mO13tEH7Sm
MKbakwUtFlFI/aD7zs83qclhCs9kwKYOT228kCD63BYl0YctsPajeTEsCJvQ
kK0bmopneKXTFOrkkcLPUU0afab1+11F83zBhuyaDzp+WLHXC7u7y/G6ChfT
b07gUw13Q5UHayCnvLUyvRvvFgi9BbTeYPIfp2agab1KPSbnaXrlJhqvUYJX
e14u+p3OTqxHBV0eCiJSCzyh6upMt49N6yfa2hKKMF5dPkRkBIJtfGI3aTA7
cL7XYl+uxyuCFDGHYPy81fUDbzl1mVw53q/pX+mtSuLhNMLfY21K8k6FjE6Q
kDL2DWfJUGpx9pK6MV39eoBrEtS5eCgBNqLXSjFRs9sx6tH6BKQt0tq8wMUP
NbVhQMX29JnTDLNZWYx0hFROtKAvubkRQbJytPjOijQavoZooXhGjEjFFK0F
MEIajBCfBd+as0Hz7SJYoQcyTNHZYnwHx/iHUGE2ts8UI7IkXTFN1B+twonM
PzBybDvxPf8tJ0dLHu2Rrwj2DsSoNUlkWiczN6a+cdsquvZXuSySgDZ2WeVn
q4Wy8gCF24M+iQJLGQ1G8Jx7vh4zUU4UO674o6d2FB+pUXFPY5mm0PCmiXZ8
Ky60mROp9S2/SUVy1h5fsOLPma2KmlXT9lVunmXTvzPENmiRlTaLiO82SFjh
IvebYWDujt2jNS9mQmLWWugd3AwXLV93b03DokEQbZo/oTNBEnZuze54RR0J
V4WSgSmoT0VM4qGCyGD7z/BhRSo+eXcP2s3uIhGduDVQwNcTG1uzy/pBlNNs
x4CPI6EPCOUIiW8KBNtJQjuY14QJAkgsiYLJEhh5OLNN9YIRAODXFBOeyJMO
NoSeFiCLNLDAwOqD0Cvtf8Hrf3wdrEXl1G21WHjqZoqp8huM5qqrp+rXYyz4
PlxopWylvDTInJa3nJLr+rh1E3t+iLlObrIfdf1cFG1R3twdcQRBxzA5TTXv
+S3VczM+i8a6W5BzMYMMCspJupZge5E667W4XQCp1OfhBTCxskGQ7pOP+Zk4
VUfv3tsUCagsIOIW5wNbgfm0jL7xjKTwewAHBive3JmEjBo8mFpXS5Q4gFyf
KOTox+xZAAHG6JjwOHe60tMTczLY1faQLCBRCcirI5/JkMLbYYozlAJNumhL
Yshoyyz6jJKH6WQBlmvnPaAxkLpxBdJe6YWAiYAOFzpAsHL+D7SzMcVzorEq
WaPkdVwP8aHOFN+RR49QqFB4CcWNCHCfxtIvfnMwajyRSifdy7Nez2CIA+Ba
t/SV5B0qpn5+lUxXIMxU0M0fJQ9EJFDIi6NNXVjE+EspmBNtAz6x0qPTOWRW
Vh+5lw9kBqLTZAQnQBkoxATDQGvJhP4RsZkuOfWR8Udisy09Z7PBEy8cXBNV
L+Q3sLde9ZzATq8hfSX6uDGnnVFmStFVrXPZ/ObV4fyrBocD/HbOUOoyLrtZ
QguZb/Ao0Sp2Zb2CQIF05Am70HGLrE4uAkrht0wM0aWN/R5uGK+Ds+/wI/Eb
++8SKn/JbwWPIP130SjiHiph9D0TFQiSffTZeKIPv/RBsQx8fBKI15OndbKo
c/wmJPEMNEYafSkKhX6R+paYXmM/wK4zsY1stEJOJcAL0sQ+dLkBEK4LpLoN
nD+T6lhA5p8vS/tIKnG2BPjn5LsnYxZnrLUqYDA45QtzCKyz7KFGcl0kbGpD
qf5dFzP4cXbnFJsZd8H80ItnR64SUrvIFnDfVYGN+HDBUhUjz8uZOdme6xu+
/19ERUGLGwcoXRvAGMaZ6P9mjtt3IRNAutqx3J0nftekz5boV5mg/bcQQKfj
U/4HKlY32JuZZ+5SqGYxu4yPqdBkoanAOHP0D7ZZgCuTVJCEdxb7iPxM7Jk6
HzSDWs8pR6clfqC8GOBSuUGuGVHGZAMmVDi5qrBeMTUu8wnKQhJDGK64WhPP
hd3n/gQKm3Y66wxEe1nHGP8yXp8Kia7Xawnezdpc5CuJkXNEe3HTnoP0ZgGM
Dw/rN0PC0GnnqvTzjdYY2lvwy+xWaURvRWtAQ3BMvlVuX4ak2NEmHc5QrcT9
75bzfu3czUoJBVhPLv76Qg/EwbC4a+Ql+TpT14PyChBT6igrlUQ1PBGfhpqA
gpwIOcWLvuIKIiiNKR4GO4On7zZ9jnvsb5maDi/kZa8sX32F0Xmb5JAhrBla
K/K562cdH8or7mSSgGrMExi6C8mTQqxvHH85iP+A8YUF4Yehe0Tgp/vh3f7G
S0ysGaXkUK58RBLZwQKokHDLFi02YWs7IAHzMDWpD1djW1tGBEd9S/VNetfZ
bCbV4YL3lEqdJRncptU3Uxu15GLYRnXcizTEKtmhhf/QmUwi0FJWTQctEMFy
5q2G4D1sCavOJtMhRrjysfgYdo6Kh6HnUW2K97GaykIT0PKpuCXngW4eQeEq
Q/qJyGLdXpRBT9aQa6Ta6G9FIeX4PeNRRuCI7k1R721EGKnyziYSEAOIySp7
gy7s+qqLCsWXR47e/0Vc0R1jNdgGFHb9gFgxZvj28VP0qtAiCptFqqW1bJOt
LRmwvkCn2lc3S0DByzJDGkxCwtgGy5dawGHGYfWWs2b78YBFgeq4KtA4EmqA
3cXqMKLVNNzF5Zvuvfu70USoaTh6xlCyMACHrJg21bHL1+Q0pQgk/rU6tYC5
XOzSbbhaKti7VCuYtbnrveHlQN9Sj9mf4JL5AfODzLoKbfV0iKwgYWVS5NTv
GC7Yir22POApycEnuxqTuLvW6fwTlaXSqj1/ejBXr7A21y7dBlJQ7G0sgrsz
ZOSUci4FLjMiYTNZVxHxod9YPSPN/8kTmp9ovHw72mzDRegwqpMXRXjsGMN0
jyxwEi8DX5r9v0LiUxpZ/KCHucgpYH9lSrBLvVntCwIS/VnYsbEUjm6YKf2J
GoLDMnLhZmq9i1c+l8VcV5N+IK868zxH3bxqNi6aR4ajfHWpej0NvFRo0Agu
N0tNgIuTGxxFajtEW1ADcWoCaTL+X8xed4/bCU9IlWcBkk5Ujr5ypTmfwODg
1TRKwJTQeJyvlzMCx5oahWql0G/fMLBPBJKQiqddKpO9h4m/2SGnklwoFUvm
kIxYUDDUG/ECAiQbqfDtlQdggjbBTY4wPBj6QFGe85a6YaXE+f7jvkygsnXV
QLiWCQdh5IC0CmAkYcch8pr1L2CxTTfPCFogthsMGKVZRaPVPh5YNj9Q6JjM
HbvvxBaCcSUVGVXuykpGSUqOR7OgI3rttSRxsukskAm0Ka02hZB9xcuNigBL
oMEL6A5DG6S1ig1xa8igVZhzBUbH7gDkA13HsGXnBdZGKBXGq2sP3yNZqW83
iuywA3nTN+z16Z8g9j5HILmuRWmEl5sherBqAGjcu9NhY99GOk+NB5RzDKNM
ex4qnIYdOpvV08yanYSbnj4xKyZTR1cK2pfRsr5xOKxNfHVZL6o9C39OUhiu
XYdeaLNjwaofNxn3YmAosobw82kW+LTspurLTY0W3Eldpbdki5WfEibN0t78
7npmPJ5z/erb33nnpy20TLMEm+PFvs/S56G2aBlOfQajAxsQJuYjIEStamHs
o4tF3d4vQk4zFua03ztYai0Td1/u3ISbhYu4R4gVCXhse25QL44DKxeQPq/4
AyRSbCeQMYPRwD3aMFQNCV4SGi3lM5ak57xQusw4+LhowMLSDgrJnDjnDJ2y
twKWXk5qutgo9MfPKrUyhIC8Tmf6k+WgbwIQvU+jF4qPA+unShDQwNXRiveG
A3L29386VSbZA5F1wSk6aw/SNDuLgUoWQDmxopDBCSBqeC+ZlYJjUgeN0eI0
k1hMbhgeCnsZ2mH6mKQv7GeJu82BfBaMIJaL2MyS+EWY8qSISH2uNOVQjNa9
cxOE1FX8NcUsEGf1/tEAPaxopX0tnzFBhCnN6zJsIL0oCqVrO82UCzVyafE4
FHUWsGIxRvJCtLZXhlnO/WMEb8aIxh5dJVERzyQGa1yvULYrWQp0ZErVVp6o
wrB+Shfbpq+DqM6gjfEDQ9Xo8/yzTkrJ3Azje8dwhwNHLxNmybbWsr/hadiS
DnIKu4g2iB7gHo8xg9Lq9Ml2pow3n+2ZPtoWg7MXok2m8aETKdgzInzCY+95
qzP+3ZNYgoEE/fs3KkCLummGiLPl/zHjM+OfsWvfmch7V6+1JGQuquEPmAS/
hW9f7j+FVy0q7ZVcik/90eqRcfXHo6E9VgXf767+OznI6RjJ2kS2LY/Rpk6/
uILrd7lfvG6AFdIDpHJe+ZlUkRA/CC/LetvtoKLFAcnye/SsG1HGSr+I1YQG
aUMbiVA81FpXjI8iwnFDCkGQkEj0jHU3rxYfPrgcwLR/ghJN+O49L3uhHy8W
BH07ChOWhVcLlGW1GQttxeM0ngD/8rj2NhTfLuVxzjBjbpGhO/Oq3FvSLKGJ
pjoHHs4OMsrmQM+A7k+MrmytRhc4/1zCoIsFr0/HcV286HDhJ+r0fVb80QoZ
2CCJKsZA4mgGE0NDigNe6l31mROkYQi0Ht6i9ELg+tlVB4kk+RkoHn4clpoB
ue2Fx/odm5OH1XeDzSX9AXnnvXNJyuEcL/v5VxL8GXLpMYolUjh/ptPR0DFM
gy0CkYTpngpLl5EdbvcF282eQ94HEpuRIBI+12RgPXqeBM92xAkC5HU1vzp7
zpMsLBerrGoAJneKEx0R3+F7OKAOscjhbIkJW0Sy+dYoxMtghqkIrsm0fqf3
/o0QLOCuR5L6J1cmAjIVyk1X/p7O0HPgnqkBjaDuRFAl+SpgvJIX2pdRLPRZ
BaLxFIDR1gCnnyqY2bvf8/A1EDhN0ENnJJVCkSIl4iO3QLvBi5yNKZFqiHZ5
sOQ6IUsTlw8c6qoqN5hrqXYBFn8uFRgSYuV23HOU1PSn/YojGCdv0eADklMh
rzSOel1oE6zW0fVH2Aa9q6Q4zWerbW0mael6PhXo38n6co5KcIrWiOPXg7a6
3qY3QUBKS95Ls0RXSICW5Jg4kgAk+nxNWL2g4aKknQC6NP7KNvGp9m1xeGgF
gx9YlOzVSTDQyi2nAXnZYCg2k2xfxH4tavl60OMsThYC25Bi3UX/aK/ex2Eg
eBuv1fCb3MSBFi6MD5kS0vds1cmxQaqKtI67oghuUy8hu/5ss3sdPkiE9zva
1/InkfvLnl1m6y66w7cw+G2fUB7tNvi4LjRkgazWFY9RkWhG/FcM3qAuJPBA
lIOXcSo8nPib1NSaz72Gsq7bQGIoOSNCNNedlZYZpKP5tjHFD8z5DTEwPG67
3MCXSGHNoT4vHKzo27XvCMkcboUNxyMe9VRZ7nu3EPUnsUHHcG9D79eBpppx
ZNRMa4WIUAtNi4TdFduYZGmDjrDvgZr1ZrHjziLU9XaZo79zO4hpSQgKrHpJ
XV5qeNRi+gmkuAagM+dpGVXKj7UhNCpYYCbKS3dOYYbeyJh0pkS0j5ISy6uw
Zg3XhCZx/y/sKyniMYEvvHMUXT142eNxTfSklil++Ya++5BlKiWokaVODFvE
YkyhW5bHL633gqxPfwrTf8IxAD+ULOGsAcAddzmuxfPsfjVAFGaT2IyRKBCs
7vjWRnybp22VFmG6wo9C+zBkYpTI6cD95WQNO85P4h5QZh2Uq73myT1erUmh
b+Mc1MToN6PXprhVrhJMX1/TVijhDNkCxcVEMCnsX5Ach3+FwBZGZ2mdNlx8
gmdnharyJ9hAtt5sEUFzcWh1vWnhgFpr+IwDA6UdwoGAQLmsrBlKThDep/FS
g2vcQehDZvjM+Or7jc1Vx/0mgUtnqSJOA9FTtObP3+XTLMaT7QEUdk9lsjFN
VtIq+bnM5leqbK6Ln/vgdwqRf81Fmei5WyTlORIQ/QRm47cb5k51FX1pB9M0
XFcFEf16Sm9BwkyOJBBppQqGDfC1hPDH+joa8hbqLCd26G+N0DKUVKJKogX8
L+rZBfOvIXHIj0tVw2tqbmbUPMq0d6xuVB6qLoIwcCpEQzaXKncHBNhRrXed
v2YRxw/7mSA0HmidZNnG9GfwTqRp+7gEGiwPZ9s9+wV3QKg7EARtCH9rnrbx
oD++KIYc2qGxeKvelZTxDJHntbjkRblIPBkhypQxXyqRqdR0NUTOw4XpYf8b
BR1x4KeBZv4R0iXQ7SySDpCCN2OKojf8fEOayB25HQTNobulzXktFunZNHEB
6GiiCtoU7cVkZ3LP6XUZV3C4V2PXGVr1PjGKH+BEGlhW6mNlYnCoWZlkxHje
9cApRaus5WODomRQPXqW9Nfey2Qj7aPakKYeOoSekrUVM945NBdImkVClU1G
Jz64Gr5pxNm61dZPCHSIwi/zV+olGlwQaDkcUUSxp2Jt7zizjhrZPYPaVCov
JPzigw8bLJhLKCbD87oDSTNKAlTT3XxuIa1kZYAUTFyf8rTvVojMWxDHBm03
aONRUPBRQTqE+qoI9fqagnqyyGfHkdILQmkJ8ALZsS2E6iKvqIOC23G8dPAh
Yu8eUA5MysdH8NgXrDLaXbGkcQNJ+oQMW7/Zy1UwdXbHzSWDEmXMaE/JpGl/
b4rX0vR8jG2mAxYeRUX8aLtTXJb+ozSTbjllX4aowpVjcITGwaiZKq/4PYIw
5ZwjVhyu3gjZqY4ketWjodL5JkLOG0F+VqxRQO8CcbEk4vWvWvbZiKlBNher
S4fgvAW4qc9TF8ECWsKs/uzloO90u0lE7wqtBEoyWYlJ7hYDZk40USmNqnf2
2UKfXwSTjtmbxlFjyZmSxYTH/YOVGxtGP2wNKKD/y+aKCn8TZCmugBqCouHI
dPx4QMs3BTJcH7qnoV8Eic7URbs+LtQlL5wFJD4rTCShoiodzrvaYZABuDHa
Fhf+dizqKGoqookWRVhLAU6hor74CjdU4G4QX9g5HJdIzbVaes9gP+dsWq/q
QN8/QGZbLnweQYAwi/SRMYia/VNpAW2J/CU7R8WSMu9XWVsLKDyjt/BwKxid
rXZf2v+D6FAoFSeJWjbgYB3rGH2DVTqXDYQzY//qHZTD+rA4WOOQ6BSCu8IU
/2ivhQyTqQhV+/7SeM4AOFBqcE2v57G+UgjJhU34OCtv8uwapJByBnw1FoEy
VDi90jEd2dirFIcxGWQKN5/rN/v+CVukVdB0TtfPrk12xSlZ9kHq+//uravE
Li0ypo0mpfw2sEtNoEuuv1B6KNs8Oa5/4EVDGqerqNieJ/jU3TbiZLaWkmyW
UIW9GJV7X74TXILTWJkIadN32/g6Vd2F/hYdwP+GiVNqOprXmF9UNfwR4byq
VtwuZeXddjt2//QZlsUBS7j8+p89k+tBCwomtpibW465HCsYjQd0HoTWXjnP
qlb5Ba+Mipbsk9txgfMJUYdwmzMx1HBDIbYns1hIojiaAUNYqubiW5fwmF7o
tojtrLJE7IcEje4mlSfWpi5fXEdqSJ8Z7CsTsUX55+3zcxbBreeYG/CuSEMK
tjVbnruzLs4MU1+K8dcj/ekxqHHmobkgFetqeb/Ox+6sz42laNv0YwmnYvE6
eIqmcphKiZpmh6u/4YTZKSVqBPU91G1Iky03MeLk3VSlGstj3zVVdxspv+Ip
KKBuCOzpu1uUAPkTWV+t4KR3xq2as/dre4OW+GJrYVtRnAzgrC4WFBdg3CiS
LuKszt2zDplxMH1px2zsfD3D+RF4bHQBXzOmf/S7oTYYwSG8x5Kz/BtXUr3I
W2330eQklJDFDMujBhDmPRDXe/q0nlF2KhfrUEGdFwYuA0ntXAi1av3QVkHg
X7zxL/6vzuGvbjBgSua/1tJdUZPN5NrzWH3XUo5o/i/Gf4Lc/79gtvyPpgWL
CxFdx/+LzWkyK48DWucURFLKH63J0QU7pxc2J2clAFyA3JHYd0Tz3XdX/83v
5+HILYoRKfii8KfqBd/KdmCOYd+0HaEDMrP14IQrb6a/NJ+jRJVZQ8tFboJh
hQqFuqMiHmWZIoJp157C9A8A7J6OjhchyB4SSZVINYPytyZqLRzr2DB9pnpc
wu6ytMdBVLaA9dd3Rp/2sTsnCw6qRbXh3lDZSwvZFNhOAz2U6Qk2bHP+WHge
bjKCbOx6cLI4DEsgUKUjonY+wmR9f2PhewpD6jtpoml1IcXbL3MHKZDZTbyM
pHKFuysN+3xfwegEKstyigVrB6jwXwNDtkJFlu+YXYo3BhEIZanLNK+7qS4a
ktaiJxfUIG2c5cttdOuNMgZnLbSrS3lK/X6tCd4Ez7WTcebuRa+SoWJNSbqV
V4B/MgzC0eTw5Ql1j7tfXR1KxF34LPUW0u8/GaQR6yZWwxCURwHO+pM7hpd9
MriExyRBTNaRjzP/SRo2J3wn9cbeCTklzUQDdoXkVaeP8LZJZvnECB5vI2PD
O60M29e/PWoZt31CtFIgpn7cnONi9K56Y8jcC/FEpPbWnooRSFZPA9ie9Uuk
z6AZfvwy+eom9Nzg0f3f4/EYvhHifEgoaCIoc0g6XNwOEx0+nHL44hGq3eKB
UarIznl7DfuJCzaoeE427L/uU2VdCTqN3O/xdikxkqma5+M+/8liT5t8L8hs
0hAxhDjrYfmeXRJY+6niUaZyRR3IL92EZOpotWMZWGpoFbkzZDQR7QB4TOVJ
g75KdpA+aIzUIL+/WcCJFv7n16HhBPYTKt5WfDiL4vZ5riHvd8tH2MJg60P0
6jqpmSwnknlssgqDWTAy7ugwwFiuvpn6ZboqKFQOjVh3kqHTzOSIFnXWZVWR
HzAMZoIIh63Srrj8kByzs0URAkjytE6o4a8EdYZQg2/6W+RHi3aBRbxt5nyC
YhBuX1eU6GJ4KVons4BP7erz2GRizae3kbsAz4ikOsraySUkvF+8BfWXBRTc
nhLBGJEOUSfGGR8OCrfEMJGusrVI4DsjjyTCjxRfRvLIn/8d7jm9FRAzV0Hq
L4FjZT4whiQBm/ifbP0j+MAWypoBZ7L8uTdGmxKcyO57WjaS0UieDDfVU+Gb
rihle734JDYJt9jfokbdZRE289LsqqqLq60r3Ps4NBiFdzWPTgnCuqLfs008
asuYy1PW2K3NCRWBRE3PdjOVhfQj/8P68SOfuEfv8syuQXTcbmX3vZtpoEBD
4Fm9aDsznLglJoBfvQe/7FKAv1lpA0QspzOAZp4OXsXn3GESC026J45ppsuM
NecNKs1NuRxeW5MfJBswK+4u82WBcJiIRYFbrJh5zjt4XadVMm56KxaHgfm0
LXUx6MHtCz0QWRd+Jldjmbd6CStQ89194Venn1qCpUMEj3dB7unQBtsmqt1U
YgBhf2+i3mpN9dbwdTWuz1AtMonzmN/7d6zn2W4XnjMWNpbSTt1px8aFxiwc
2muUF+elUuMzoCtvgInsjNrsv8CpV8JlV17ezxB766H6wT9tvo+uQpwgHHLl
2JdauMBRWvEUv8D7q1Vg8PPFJX7vHSnm4ypzB9gzpL0Q5EbPJ+fbc9JV7ejw
H+5PMkqf0eliV82q1GPTKMuAbt3203IC5vV5xNL+ge2LwVrclyAlwEkjfJmm
69Neu/oCHqA9j3vkBASJONlwZUy1ud3a24I2HDxr3iE3X7RfrXwGS4/Dz3D7
6TCIYi7t3uTYC/+/Eo4vlcdBpmiQyAGC/pzolnYFmajgvy42xXA44dBFLIRK
0oyPohi4D63jP12EnHG9fqhpMmtmh0jRkr7LNhLVdgF4GL6tADohiOkhkU1K
0vq82eKCvsRdvOrqMvASB7HgLV9DHdgsmcu0aXaxUhX7HjHXTn9isGo0yzyu
dmXYIwccAEUH/rOkbso1LWPSUMmxG4+7J5cq1oc6RZTZjIP7Bx5NmK3HtjDn
vIuABuMzzNfgMl8qeWEMQ/SMz0alWE5HwsGDZvuCUamLHSdSDAyQawrM/UFO
LrwddcAe6KSjh0FaQMRfFehmCaC0m76W0KBB7Yoynspa8Ie18w4xEs/x7aaE
DrjaCy2nciZksQiCPYLNuuHSFW7nu2AGKVAjhieQR085rRYVy5aeheEg3Rt4
eDBeIxQXKTm4mRdiJAEx8StOY1kFrnjexfcot+nAHc1+d/yw/NCBTDd/5D4c
/CP2M6yp5hQSLiFvbwwweSr93/HO6+ZsMSqrFE3/DIx+WjBviADhOAzpNv6V
pJlvHFWWhjeSQKv2NHjXk/kQHzUH3N0H7+qrjEuRBRC6/wLlpj3LQ4ByznjK
sYzXoAGGcKOLT5jEJM3IrRgY5VKhrZIiSJ9PSAhms9ZN3MckOZtmnFccs49i
bqX3ELCGxNeDsZWcJiZbf4FZplTYaD20UfOKc/VBjjXj211r9TtMVW7M02JY
tx6r+t3OcBF3qMht08e0TeUc9RJzQa1lq1dqNkufzixNI1X+FWZqv0O5zLVr
1m21jjEPQIoueb2Qa0OVnwHp3vIaNNhzMNCS22D210i0oy2hC07tJlBOhtsr
0sZ6RkVN3E6bC8+US9KAVKVIEEvnWypeiryU+9lAN6OhsuKa6APtISH8F3V1
dvb4RmuYv7leahjeQQMFMefvT26P2D/wlGm0wYTcKqwGeIo+AwVfH6SpT8bR
uWK4wyORaDd6EfWvvBPqBGrl9ksYMjBRR/ww8Xl+jyQZcdOlOE0GWiS8bCRj
TdpCwz8xJ+I2kqFZSagcMhdv+p0OnsqEM+eoTwy3YaDCI4+bE2ywPIuFrVvR
CBMzzqHqm1U0rqD6XIccfFFN6NL0KilBnn2OjzQNFy7D5fQ6ftVL4MjvTa+d
aRctRGAhr+ayF3lDbhl9UthlYb+gZYVkIwbAxthfF6ICfybnRMndErKBQQQX
s9TJpzLC8QW1zPjK27LXvjubtPeYGDBJgWw4MdB1/J3H1dP9ZG74R5xyJ/4+
y5puMbX6Zkoa8sYsY7ZPkLxUrMF9i/y5zdcN+1GeeqCPUgOSTWKfeubKG9I4
h/Aroh4CGF88uVVenmoMwXw1nf204HxltvQDvXyZoNLjwBHCQy5OdYmf6w5f
jdScwZ7oSZmdG4iBAXdvqe+YTTfBh0fviXMD1Isflmwi3fNupi04OantqQup
8bDZM2bTY7MNGstHnwPuz0GmRkD08o+EKtgau0q426JKQFeZOQIFLZvDMpB3
KJAP0iMPYYMuBneT11vGnjDIbTIHF8FO7f4Mkb7XrvF5R4oWxzEYnU6qySb4
VsI512ZF/Yc9LmiO5GbuCb8zylfd9m5kTxx3ljIgH5lH1LpzBmGgb/T3qmR4
VP8RwmxXoRBGO8fDpR5VZGzSl/l7vEpDrLDNnIo87yLL/ym7kREMzVPTXrPJ
er4rvZh0Zg9bBp/4kTqisn7xAw9ehAx1IRW/Wyb9gr3t2Uhi5XFyXNpbq9Oe
wAtflCh9j7OxUSo/zI2ARy/xJWj0kF1kdpjjooOA3QZPe3lhK03QnxylJwK3
hXeMzBo43p4b8w2ASur0gDCdmmytXp6QIdXG8/Yzm4SeZwt44/JEY1yWvwrs
ohDmQtvNhutAsL+J3FYRTsrmF7iM+rvdbcjohXDtNz+gbvy/CTmqgIWecIR9
4ABNwx6KkZGFccGexJbQZXt41LTASX8n3mlzOLCV8qVnlp2Iz25UipsxaEGo
plucrN7tMj/LvoJRALLK0+I3iX+zl0SC/znV25jty4ccletwGYFlGf849l8O
dAvmQYBnjt6NHztyoIFlTUrcU6xrO36RefnsR+R7pc4l9CUfqaR8McZOZcsU
bv46nueq54YeWFsxG5gVdRVrKphuQimBZTIiB2p9ihSzJnze5IuLDy9lWUB8
9M8d1rCKHA24xCW9Bs/7hbwWMbQYahxkkHIMD1nzMQajla9dtcS8XPkaYSCn
tVq2ld1fFnNq5ydu074bbQFmv7YF+xv1ieXRQV2Gt8k4BJ2lt/Ux/QnOG+r7
7xmOjwLaWfO+G1jahyJ4VaFIwMsv/4Sgu+aoyrvjy3r9IcxMZrO0qJOh0MaI
VxHUBtOOrrSpLvzAr+zcrYIqRlljxQoXZehNcUxz6XOlArEGal3dkCnlEtnX
MV6iyV979BJAZj8bAnuUB+b3S6CPaInhu1amVJ0u6b5yYGTIFQ7MNBCpRsRG
eS5NVN8YVkGn3/PpM0E1igUrmujQi9/anuXsemDX7exQQGgIp3wCwN7snwtc
bZXL99Y9SNSjPQHPjZW9/a9AQNbLJyvvHOnOHGGbxY5ty1uMyLf63/5aV9DO
3bUtCl8BA3K0kareuT6HvL0d5fU2Gs/6MHnc+CWXMisYzCvqYeXoIOVzJ46r
3lhAlI3ACRF9iwaZ1Imu409JIeNuQQ5b5FJ4yW/Ksh7Njr7C5E0CoyqGlsd/
7DaqIq6CDmFCiOaJRzSP1nFAZtPoaQDA/7QjIx/wtYVNjGZ1hZTJQ8vgECon
lDd/RJu2DCdkW44n+usY6zqrmeRT5uVOrmmhSVdKykOlGOhc4syB4WBrDUFO
r5wVAKO/x+F148aOm5EeMZGY9fY2CI13aWX+PmgA2euTjIdM2Bx73nkp/zBF
Iz2DiZh4cQ+RFmBRlOmLBp8R2/7ycf9G/dvCKY1nOvXYBKQB/2s7EYghz4KN
xNeVmZqX+K3Qwzoau/6gTxI3vOpJYH6pkYDvLP2RQRRqenbQSyEMlxwu1lbA
/CRL0KGCSTAf6xVq2qwwL4GdyOoUad8khw7KlgBLBSe9quQku5gJBRT/3FwC
n5CjdV8BAqqEt29v+hUHueaUWejXlxFwE2b68QA7QBT9WXS9nV87QB6/Be45
Ds0UNrj9+AsiGolr20/lTiW84i+wAgQXLA+o3zn5DblcZwpp3BrP52OD30ed
H9EgI+/I2fovUPHw00T8q5zF65Xo+iiddSg2TNnFCkSb9oYbJ0mu72sNFJdd
6Phl2FrBm9FFiuKBgGdJ18dcZq4cxh9pn3U/sHMe7HAcrlIq9BGbwRF/sbAA
2ShUXz1uw5pzHC+idD+yhWbbwCDuLWa84a+Ww3Zqtacpa78Wh/P+xeMSeC3G
eGevLzyRq+BO6sidRa8rt27qQl8NSut7NFA2hH5tZTpv+sr/BWryN+uc3IFi
nD+y0WSREgNxWRXhzA2tNsEOZO53Ezkq4yvUy0ezmDIjvVc2HKKQgmJBJcN4
LCbsQx44mgqM613u2BygkEtU0I3dAROe0BguEwTlJ1C0t0TG6FfrSQj9yKum
SDIdCOxkiBLAmeWt/06JYJ37f7AiK7fkISA29MWHY7ED8mEQZTRSQcagV22s
4b/IAjSDretz63/wvUM/W/y6H9tR15dSwnl0ntXhxskyEhVlIvCS0TF19VFL
LASA3oVo4Md1GnaQNPa7fEbVmpgQSoLevFSg1vRGRI4wHFoOLoZgUVPXxyY8
dyJ3mll77IQ4jiCbJ2fGF5L2NdRoT0z4+LxYrP09YcIU1rTz0dWuE9SZvoj0
LyG+Z/erWGOFrDhDrfxmjQFgmHdkvV3bdWd0+9QO+yRKIL3MXMxR1Zqasrlr
2+jUfpvWXUDwxUzYoAlpv2rNDHy2O1P7kBtjPgWfGK01dz9M19meD7TjmfXY
D3KIYTAPi2BFjJ+GsxqnoV+5p3TI1zehOllhaxOkpQ0uQqAHj3/L5cDQsBXf
W4DJAeCZwH8XdLkHiQSKmny4ar9e6Pg4hbtNBKuHk4/hAfD4Zbpax0M5f/1/
c6QiMp5+NZttt/Hd0sjD1PUuBr+G85kunBdTTUYWUbZs/GTZEewk7dosazp6
u3/xubXA9afMRydMuBMsx+m/l86VS3rnaITy80vXfgjYkBES/aUQluHHa6iR
cs261QwfX24pLHpxrsXyNcHM0hC2qrVlqeOK2E2XV9brm+PYrlGjS1gL0lyc
+oKdbR10XDtqjX/NNTnKGMqwBv0lJKaUEv92jhpubBTCW1vLFBiBoUiWJOlT
7Bnq0DXjFlfeRE3HfOL9lvEtKuI2yb9crXvi3bMtOOYBA3O/NgSp9USV+Ek3
MFBT1vYLI49hhdYIFeRapQhN8+uSyiN0ZJ+5ekMPWJd+K1uwMgE24tndHe96
7/DZ/H2vHIwl3/12EoGNwJdGJtrqEJ1tgf2iBVk7gn6N9ZiuX8i9vILhvkyu
G5iwziMticV6nhEuvejTXCe1bzWpQytbJg53bvwbsoSjU6VdhCRoaRl3evDM
afxtPoZqH43YgfIz0P453BshHY/O1sUsu8h2ANV5Dxhk23qtCJRZC4O7EW50
y/KzKEpgtaxczUUa359nrsINUnn+kTu+ahA97ehFeFauvKaNSQkx6I/LFp5p
xe49zmUoJJuM8RgP1PgYs8UqyKyvuc0ZfjmFrv0suF+d4ipi5FCDK26HrJq+
aJPNEo0PF7HYD0X7hYzWw4UBz3fHBavXiMcCTz6Fwr21fzEav18720gUwjPJ
q3KZGxejP71AAqsQ3a9XQs2owjpISyHY7umTnZOZJGvXZWQhX6ExWzuSte7N
dkfAjtFKvHjdYNI+E+tK9IAmfPXGLS6rNGwAs2orpgic4M7oXdFhoYmOmhgF
559tThJMDUDemfrENhYUVq2PT/k/Lc2ps4igR2xyd2ZV8gh2EgNb44rWFYZK
4+8bBSgZu1NENi7mJgPXntoF3i+mMm4eQRS5L9AflKlB98ixvDeKo6wWC92R
ysHO6poY3x+0uRgQj8x8lkuMV7W/T1rAnXlrz/0kjALYrjTCVpBR8EAheAwY
VuPt8UgpsnBn+JmZHn0340GiYly2j+bdhq1j68otAGFFOc/BDa2o+bfNLQR1
8SgR3ZErYvREGwAiU2SVE+I259IVSBDxuFnZ9WlqvAkiQ6KVldHNRupnwBBC
iywkUR+Z6He3yOVEYufzQUJVIOdaeLGId5qx11BgIZMq85gv8vitWhOrcgNI
9UdC+Ebyr+8QMdPCStUOxSbxZynzbgxL4Jo9kLiGRJAjeGmmBzii2F1XH/+I
zb/PEicJYdv4ozo4aTQPJWqyKLO5sR6pgo23K1uPhAEz7WXpI+QsRA6ff04I
zyvgl23NCuXYIq81/1PrMwL84z2hqj4xiVuwJyjpziErPg833eC0CbWVthx3
JSHammLBpUWgIPyvRXQl99c+HboD3gCq/8d6QnPlZdPRq7JEGajljA+K6FA6
RNhwbzB7KiyUossbUM6OtQHBykXdQeDBLLXmK2iQwPN5wqIPq59qZKPf8rhb
iCV77Ux6zN8jnJKtCw+68VAwFZFay1I8ERRtI54I2N22pNOXt5KSzXrFS/ly
vrOSraPeplPgLwOS2ivER9l9WE2fRCy/6wuZV4dH4SQ6atYA5qvuug4GH3oa
htUfa3otUREOaR5Qb8fkSjfmheEKzf1LhVSQMmObvIEEWDm5tjv6B3YvHcw8
Q8rlhA/BU/XvyTk0BidouvfNwn16CGfqueoG/m9Y0gWoknLXKWoAMKpfRpud
p3bvW+n0rJ3K1iLB1ckEN2LLLxGkCLzltj9rGydEob9arqn9uyBUDMyYI8KP
Ll3YumXkt7ajm04IALL0f6hjdD9L2+oFWKJXcPp6qmEl/9zmDXWJgDd4YwIk
BaBnTol1cIAj31tOHWd3Y5LBl9nQeIndHImRJR5h76VcwLP/+3aCzp8cF0uL
pd/iChrLtADMngowNBC5we+M8LXq1Mm4aM0wsFpaV8IcGeJDlBfKXhCFRbzI
CJF2RL4JztZg/Eqy1xi5NGJKqd40GjT42IZVMs/KrQvzOjDzKp1i5kaCNxvH
tyllQ+PFK432pUY9lfkSwZn5lWReuqkhXFkOpyEFbMSGiW87zJU9QQGqlC6m
QsYLDKBFgBCQ5GpTLwLtALBvF/3fAbTH6Ptaux+wimh9AMhVd3/gpARu6DEU
Xh373s0RON9a8g76Ri3ZPnMNaO7XJM+/ImTwKsA6ttZ+duLjLCU9H+xR3mib
EZmXyd/yPL7cLO9JmEi1WCY4axjttw+so+w3BEHtGyEpEwDwIiyVkWJfN9ex
WyHnyyZFoX1DehwuzB4uNajpLVkKZzcNUFKsfgcSwzAgotKzJ3rEGmeTE/rW
lS7FRSF5BcnaTgAJmvzn/3GWyhBJWKoC01KnOe5a8u2QSZONHP9Y1ET3U3LX
4eA7QSm3TJpPb3JA6TVJCPb+ct9+1wfx6Dni6FcPN6+1pCQZgOqYKkm3ghqJ
sto1OJUgp2ebpLl399lxKB0Jr6WqCWxpU5OASr4Ogj2oCGBfpqeCjMirNQKf
3W220MmHuQHs2i7RqgPo7hTdqjwHilxc0RezVK7OBOqzfJKbncyqKlp8FhNn
9kkkf5QR3sBKUEjysS1sAsXeEUre9Znmkyg4efb2/QMGlv07MPpellqEQ3Sx
noFPUug+qsqCDN9ufQ/bKc1+dN14pDlkGWOswCUdJ83w/UW7K+28uq0O0MEp
tad89vaiKsyrqffF2157bcVNTaduZPeGF1DYguiD3FbCXuDHE2DWbIPPzEOd
GTeSOmT5yk97CFKD9hyP8UFs+SrJMjV+/qimCi1XeAB9pIos40vPrIT0B5ge
CNwuGAUvDTIeyJ6v3LIcjBydCSUPzQ16KLGDzKIUquAwqPX9gdQfvslb0Zk0
XzPJ6MKtGbN1Wdv8uxpXD8/sPOH4RgGkAdXzHoejmV0iTZnCVV/F9SQdl7ms
A6ARH7ZvqUS1bDeIwep1kmmJ9aCCUd9yEIducjj+5WETm8VUyAxTkv9cpkpb
nO0ISVzr0kV/ONWGSDPMY+uHBCZS3zPktRrKApLhbLU94iJPPaWYCpsonq7f
JLjtJKopqD7a2rwa9wjfQMee8lpUDzKookAH7/XyY+Y/csizUlZjYM1+lp8o
WFP8EGyEE0G5ryURQpFE8YPNwAKlyvEHsHR2c56JmKowswIKqumyOz9YzQyV
U26JVHC85WzcI/4PRBItbDzpXx/eV57X3lC73lj+ZIo3VAgKvK3/199GdX4c
l1lAv6IZChJmlVUeRS5XnwTp17ejMj6/baeKSvLbC2gPopA//QiqwnBmqQTL
kcpHvaer1fa9LFtezazXJ8tcVOaLO9aQyIuhAyKF668n8BcKnPROZldPf1yv
cOUvS18zdnN2KlEethVaCJyu8rbLMfzVmRKi68nebLNzOVVcrxRGlvwNtsdV
Hi16oUOYcTsoFkAK1A6BV8heRktLpcxUKi4nZov2kS4bY19RLEEHRkGIw/OJ
tRNEfboI/hkreg+t4cycw+I11LlINnXm8s+2zCYtItKAz/PnF8syvKYO+EjZ
9vMp0F9QGCF/vZokIeQpPlY+Zzq20XI3jOLKJyxi9iQn9oTiW9wDc77DII9/
kBIA7x21rV9hsQYC1tyJHN3gEV+fqgKY/bSEMtyoSg2vvB/1NJOVX01ckxhY
TEaIJG3LTfzn6qgYgtJLoTKuSPee9/lEZNSdY1QSKov72ZqcYJVbWeKqBgk2
8y1SyCuUQ02G14CWuilzi0Y2MmXGoER532PQ6ktoK0x/HZiClM2DxN1ktaUs
gx6Ggr1VxhmgcB8qan2vxZKk3YuLVlUQh6heiHaShSHbdmH5BG3nRCeloQu3
khd8PDs/Uhyy3Q6Y433ZeI6h477B3nsQiSVYsGlH2SPcSnOz9wWnOa2q1s+z
gDDK2+dcc52I8+kcliMG6sTHZ0tHigLteMvdyCdGqxy2czwyM8iWJWUuxRUA
ema0jviiR4LfaRK+5YzWJNRtBfuq2iK2gVtuwXXRFX4l0nZlOmvls9EKK7Bj
ElKrd0cwNz6r7/DVECRtBBQc5ZuFmFoJd5u/HM1JYw8sVyA5h0QpIYi7iqC6
9OFLnI3DerQ6E0JbWaNP7yQ4CGVWcJJPPsSeWwmz7BJSnsCw87vcilgAH4zL
80V6yf6BfUeiPqfbU8hcEWGBu2FnmKrwBVwP/VampZ32bwD3qRA8P2JAWcLf
pj0yIdAYl68/55j5VfWxi7zDMkcOYzhGa78IxCWi4ecLXPIdcFzk/LtaCPE2
LrZljyU/VKNLSD4fOSLYE+winYp1PRaOgzB//RzsF/g7UQQE+3y5DWW8qPCI
4GObkAafXDtXkTFpqJMYQkO9JVp9xbw4dPll/arFBeXtc0oWEy9DyKxKsJtD
mMN4T1V6ZK4mKb5EWqxYFyP9fjoslUWcLLiwoLBfdvl7ZDk7sa/zJCl4/cPR
QCyGaFOD1kFr/frYO3XhtKXu8BLpKtkJjKyBAZACtzkQWPUanbFXeoe7QaqA
j+prHSsgblBAA+E/RsOQdHF//HnUbpM8PQVHtqF7/jgaxYY8rp5f/jsv3VJ+
qGqs8F5kZfKhL/wKvnB9J9ru3yvbsjGJyWWlTZMs/3v9hItUySZhR+TcHHkX
FfWPpleX1b27nIwuyhaLAEOieM6M88uLUB9TNKPEauakqmasUqZO3kYi2zw/
VGyUr36TV47fcuCzk8qNgA+vVmkG5HVNyAgnNBLSWYIRzYpHFioFRjLGd5Dm
e6UNJW1QMz3jz9myNg/Jjc0D6+Mylx/m0cIKahaEa5dvZzh8USBWFcuirHUP
a9/V/E4vuMF718eMbmRnoiRRoZAW68+K33U8rCEKxf8N8EUBOV84+OivAxHt
C47OPX1E+E0sJfoCGTBCmAsj3hDBfgrn2wslR0nEMSFyHIIaIOBTo3bJwN3N
ur1xAyBj/B35YXSGVtxG9LxsdKyRgtEZe+lxsqxV2FI7jr7BJufzxThQBjle
sfxfOu1RXbNe8wGwSl4ZR0zFFbx23BoPI8e1V1BZfkM0BYfnwomNh40ng3J3
+8uTBVaj5MzLKUiAySj2KvXWmi91mendOvwl+/rfq0G99TyH6+e9UOEJzuGn
YL/t2KCwQ0wsUtaC/bt7koTuU71/kMZUYsXSVYZWnK0eLXUz8TR62SrO8K/S
qUDM2Jdt2wtkKkRxMo1Krmb8cwBs3FlIyZOXCrOIuWRwrtDbEFBmFnqctt/1
TT75XSpY0QtoNeYvCIjR+ISLpmIzBU7R7a2oUEhkcX1fJQ/ZwiCgumaqed+y
lMyj0WxpN/vKENVZBUbWSzYZCYks+PPyTRGkgt4Ki4nAAGLSJipwhzgtJsZn
ZquL1NNsnGkW1bwRdk4i4s8BTJN+JKLwHhOlhdT+Y0omxPrdpUTV3i1P4gHK
Mw8vf1j4d7mxkxXnkiMRsg/GJlYgq5WYBO+MDv2qAYRT5QHyYfM3kuk+yVlU
NF0+q9ZHUks9hIn1hg7flSYbllpwc7j/zElsLlck97BeSPxbyhosoW4o/O5n
yM/3tZdIctd4jVbVavjZhLXOpUb+UucRUmtnEvbFRfepE/X3ulca2rSpcVln
anueDDoC2bGM2gBb8cf/7kOvRi82IyofSASovBtVFLh7G0Ya7NPHwcrQEYNb
jmwPHlVrTppuqUdgFvdFFnfozdwVNjD4vlnb0SIMextMmtGsQMl9JB6TTqtH
CpLtfaZCxU5xp+jCHUkcUb3blFfuDHjXOZZwvt5Xznvz5MygJOasOQVdht0S
vgoCJE8J0KE5qerdWrzgl453G9wh2YszhlNs53Egfr6AF7whxaJduir4VC+/
dfBwKSIpLtvKHcejYsvYW6TFCcTmTuz5xNjmaAg8huclivaH28W1UfkqIdm1
gtueqkw41mv3iMeIu0bpdIbG31L37iXBOYe/vlNBLX2jKeJgxlYMtbiEa3Qv
c9rXapVgig6PystB3FiZOwJi7rEwyzpP0z2xYOjTM+6RDyMsVIgJDneq25wj
2LgLWN4koK33bYfh+HLKldJ2mv+fvwGLhqXkq1d7DVOluEKsNFSt9BQKejCy
3PkayXnNiTGg7X/PbbAGVzoBdkMJHW2eoYyJqayAykpD9nWjDtxpkN0DHrgn
OVoZL+lrhBH4lC4mhIT77/VkodfgwVaYsNf8CdLfY88D7v04tai5nBceagdH
V0B992QjZNlS1VS86ZPajs87ibF0ia7djAB8T10cfbP+398Ugvhloo0rKG3u
A3umeBsHYWAGSWh41fVCLerGLWshLxeBA+96C9moXKoZwn5PDHOkDDrxZr/G
92ezkS4TnWKY3y/s0rMWtKYGUUj76KZbAJPOkDEEG67KU9ch6YwpLRWAT4+m
CblNWZ9cbGNLf9hm3Fka8cVFBnjnTqbw3/w8j96tcAxeKonNZjpdwXk2jQkt
smSXmNJ1SKedyf+kv/bpgTHIfO1jxsW0yfQCTj3AYjJgg3grA3AUcbMT7v7T
kdR9MV29SVP81UVUqre7ARINGr06LldUcFsuGHaKKWc38rlt3sRBrggEd0b0
DHSWn2CumaScRQDst2dSNBjsnddnZL/6Ue9i4ziIzrxXQWW38rHCIy/4HJgJ
38sPu83ZPOSr7gdWa+OYTbeHsz5a8Yco8TbXJ/LqjGp1AS76tAlJzq6tDwCD
1gPnHGRSg05lfALW7K5mdY7iLr+W0FXeo4Fj8LjOYUOfn/GNvBmatILrIAyS
MXSEuZ4RV9BT/cDOtteYecAJ6KinR2FJ3zCAr38rTCgbXOhAKVa2WRXInrOF
p99D26LSFZmQkx/tzZE+REbrqCj1Q95Khs31O0+QsS1+PtEUqx73RXaueJyI
IV6IoHwnGCPRxT5fJQcvkgJZOdFs+hs54ml/O1D4aE93ewc+UTBr4QYpemvx
8YJQYZL4nlmQ8BI5HPjkZQKCkKIpj5JbTwSyn4C9PCdxGgRYuh36nvdIfGiD
PZDmz+wZJz6/dBenUta8nskcCab18bLshyDuJuONC24Dd1JhuBVF/C41JlbR
plf69HbSGQsutsDo4m79G88EQJRESFCNwJjEkVKx2/Zjboq1RcKAHnvcMcA0
JNkwWA5yJq+WIS5Rn//Bhq5CKapikBiAJIbuLW9sORHDCzNdWrewNN1srdn6
kPYXvTomWiquybcsVLww3Kfa1vJh4joXWmAfiWWioIXRWROG6TIfVyo0Rpxa
YdV7d8x+EmBapWRQw9e91MjddqgRIUvIzcMxHUA2io4RuS8vnJBly3kno4lm
ncKoEKm4OsfL0izltdm8jVh8zmgbW/HoQoUpFGjbOZZUEaka+axc8Aq0AOBL
uUkQ8O/VtXvzCp1JEHOTZLQubOzKObofokoZybadgy+7dx7qVyyo7zFtfxN5
L7hg2Ey+j3wVMdJgsDNem2JMqDfJDAwIHF6SRDSFvwVM9udcZ1aB+NbhYZfF
hDp3nEg80EqdGwTJIxsN1f7/qj1VxKAzG+6b4xfigF8dWb/PbChSCgfgikOb
26FSQm9ivaEN6ql7c8dzy3qr9bAvEV7k2nuW+9eyBrvnEsXyncaIDxKiC3Fv
YWkSkmy4440OIkN1sXJFI5MU/ZPRbQ1yzVaZAp0UEW446AJHw3vNAHhL/JrL
L4cN4mMC29jA7GI9NQwJJD5wi4KoeXRPzgpzJ+4P0DSxTrnuVnrjd1GpKd/z
9SQj9APy3BpuT01uVqQlyAEKKrJZqit21sWsyK/oKP7a6okzAjkkpwwmdryh
+OOGLySgirljrC364lgbjCCNZ/ZPbCN3HGiVX1tSEGYTitRD+CXBuiGj2Vd5
kuoEql5kX9nUHTVI8MQmsY5dNFGsXyBKizjKiWsK6Grgnt3TLJTPJcr5rkdp
A0c2N/hWjS31J7kJ9Bn1EJ9d1RVQO8panKDGjvcSdaLrNCYBOYHuKsIvDHIl
46J4OFzXNNkS7ZY64+W7mMeZRjGiYQhkJc2CKQxm1IjuSVYQFzoj6XaX7HYE
YDMhFDOee0/nx5M/SHinA6ehyOyBabhAeaA93IIqYYo/UgUjWV9a924lYy9m
y5rxPS4fWCnKfpVqAMlsFZ6H+UBzdbRV4KiuCpBvoCmzITi/ZfdccNu6m7lj
4IrGAw5+xDniiunn9GTayEDNqt6GPq4c2jiy+2XH9cgOfSdfd/Aq44IIlaxy
4l44Q0jb6DIWGDig4zgm0EfdinRj6gX9EwlXKN9LQ0MPiX+qfTys0jiYd2ni
249Fs78TJxcmx1wi5tNcI0jjTftpws+tQ/5T3CPGhftj25o+IqZfJRil5p+b
6HvWuRhaN73Tzyy3VxLe4ihXoONab3qxfGEWV2W+vVrUonqHyrdMNTJPs2b7
m4md2Afq2AXTqu/fDSIIpviJXAZlotCcu1ztgVCM9uomXaVKvI5Yc0grIdnH
KC2jpqU7ELL/wQG3qlEwyD6O3kcBqOp+rSZGlGjOeO9tVHTiL6oguztOzk24
VMQWbVQi60hQXTrY4qs00wEEaUL2Q6dqWcs7d7NpTCuabIon+H/t8X43IpUm
iWWkxTQlVCMH0Qsmwudc+AUaU3a8S+bmQl835XRwlb0T+sSPJfzJ+rf6+yaD
2ofI9GqfZg9fn0CL0bU0hcLexbIWp/+DceL7Jh+0GjCFj/DLSnx1Vjkubzau
eofWP8G2r8cVNRH1eIV/CDFkh7is4gRrm8mM/VqDmZgeTLA6ggM1FdWJJhEJ
drSIe72xPnwmLK3qM7AFzRLOLLAHyln/AGwUIoIbCuzy6OpXJyqVV3a/JCg9
uZSymg0T4wJ7qcYUECJ63Bj0teZb2RAQmvZwSzTMjvxRdJb04qkEAS6XyI8n
jxRb6vcd9Xdw4fRuKyl1aRbjkml50ArUr7A6sVGBCAvrWkVt5xx7y9rwqztJ
LdwC/1oOtLjmWhCB96dv6XZSiCKs81IWvLhgb55sYXRZBY1qi7QayaV9s2cp
jWeTBWBAK2GZ9zx+5kazyicE2asM6+xFK22mXW+dwNI21za2GxuMxxdrDj/4
1D8mKyFBuwmOtYXP4rnWVaIsAdDPiNL9YJj/M6xoabbZb2Cv+ZeJvJLCfT1J
m1CpXrnUMMCZf2hgHUt5wejVh7xTfHQdKcBFGYF2aS0jBp5I3wRxrJOs4Q48
demsnyEJaSz71zgaxiZVYSO6gF03aGiCZ3gjpHq6x8yjtK6tkJNX3NTzXrOJ
Nhj4RAxcD5esM0xxXcSQWPWnioo4kF6fCMiMwNaqNUT7b9fsHX5xnk3P86Gz
oCtHKhTmMEZ85T1GDBT6hbH0387ooQxMnpMuU+U1GommtCXhPmJdRRX71/8s
vYKn3a7EEZBEKvzy1q242kjz3JmpwWgg88FJozQNYRW1J8c1AjGEd76ZHqFn
jYqPfLsMymbUALSeQx3N0rFbN28qjcKoDM1Hd4Bc6F9g8jzt43/80731ZAfF
87kIRP81kYOEukQSWDk3xmv7f83qIE1oy4OMXlPrj27Xu7iecZAFTNe89Izw
4SK5FCvttEx/AYKGkNuT/36XEAv7oqtsHCv8NzltqT9JdEcEmm2hulbi+fA1
TYrGBl0amNsD0lI2hhPSdmPFR9841W0A5Eb00/bF/3gAHy+a9lTzsDZUWmYO
JldRyr8MYzCFb/fRTz1kOUE3k1/eSz2nTKvpyfEl62ESN3YXHtJbZjKufXr5
Oq7/MaefJtEtQYi0n+ozUkdOdX/wBzXoDXIbA4bEiqRjsPo97D/yHEMyl1/7
UvnOrFPYvHcUFTS79GsUv7bCAmH4W/N8DOpamPa4/fAz6byYmoP2u/XDKhrj
U2j3oL9EFEfZ1Xi+12Lp7QQJXR88jL/AOs6prfEs2BGgn06utjPVV3g5pUPS
f6oIORTy0io2ayMANbfbgkK0Rkfjfn6OFZiZgsRH0uYNbYzP9QIuXylgW4Xi
nTAFZp9WLKcwJO9BONbaLLd7yEJVRkoaPiRP51EERVV0fKgDHh9w3lR0DXy7
9PvzswFr5Mo7M5nZPWYccFRUBZCAkJ93qkZHRiImdPWr/5WZOkWi/gm+/Jov
k+wHG5vm+b2CndToXEOOemsyepufmFVjYcpn0dHkXTY6w0e/MAfqeLMaQDmS
zjBGoouVaL6jI6bGsX+cKjbvtWTMsP8xp+HFuEKu73qRAYeF89QsXU/a0ASI
2hl3DoDajGDB0iHAfBlksUQAGE39fbA7P8MnwYAR47iIK6kMPP/6/WtzFiX4
0YeyPlqn8RmLMJxWPGzEXmkmsxAfub9kc5n2ECCRYgPGHaaHNVGVQZKkQMrq
QLN7wOoeB5Cc+Ht3a7VsoT5YR9kveNQxbq2xhAUYJJXvKASz/MrWKVZGlnzt
nHEvIEd4tE2czQhNyZ8CAKFkBVYsh+1L5W20jg6ldOg0ZxsHiyHnmZkLapyw
jrccvNK8XZI1jiV5N4w3z1pYVP06oYVMkD7WNHkEkN7FIADF8CR1kc5T0Uyu
J0EOdgRrf1VhtRDv4sZi/OfdJkS6CS+TreY0jjmvvmGQ4DgPZUGHCv0iRusi
aO9sdzSUTn1S8Y5+znXFVvLZ7b9FB6QFc5jPljS9/2zag3r1y+7vmGsG54mz
YqECuSxWfTg6Y6aaqrzbty4GnC6LegF18lk452++MKABBmPFbMkjf4YNdoVF
SHAeAckD9ABzqqWyRgcUb2wT04LLvFqhuqJO/Kdd7vlAAdebO8/iRRn/bxCN
aqTGhRUZMhF+QDtMNl7TeAict7LL9kv4iV75Yuhb6xZ/RYCzVgTwbW9QBwAc
nySjf2uUaiC+Z2RF2aU8eAXieoYXlFnWjov1TAuFMrHRyzOGrADtq0HSByYz
yJbQcCMTWIib7QG3PgDudmmJl3DeIx20ZY9MuwLH2UPeGxJxw7honaGNyzju
TBRl661j2XfEp74kDWTi5DxPVBb2gG3ZONkepLeT2sY0x41ow53IsVWFeMJv
Fj4EW0u4Sdzhojm/KHYHCQ869GNHc5AWa6rh1djzlVMO9By7+ZWkW1fK4Ge6
jNYWtZwLA1L/fyv5D+a/ILPXkE25XjVQWeSANKi7j+HZCmu0zl4l8jlcAaSi
sqi/EKsN0R97KR1vjTk+VvoWJXPeiAsnoxoYlX7xjLcB1MqXNREBaZRl60Kj
QVs/7Bt1NVqbcEeVEd9S+3whZwalCvfk7VExp9geyS7NPWjduJQ0hX/PBc6q
hEMAZCJIN4QqqJkc8lkwYeaYM9nKcQWVlIX8iru8zOMZYy2aR0WvnFW8L9W1
I6Ekjd++L0WQixdU9jJygdSKM7r78725oc0Y8NGlwEUXS8cV9wf2O4jtuSql
c9Nl0jEVUqWmWQgea9JOr5VQrCAqpmzKYQLMsax+g3GrdmEHn+SOyLTcZN4p
F6jMFDCfA5z3oE1R6RjThIOsKN6aIZnEJ/3pGjGigFb7rO/SiQ3U17Q8EE4f
sb6qKQGQaXGLTfIpcWoDsF3cba8wYKXtPNOqvQAc7CkjAm1gGw10e8oFTviv
UTua1pWiltGVrKR/Iv+WlXQzfIyFmpIPMlEGIuVk8TY2k3g1yegj0qmJ4Crl
G0FmbFof7/gds8ZFHyijfycKekXz66x1Na/D/XB+9IJdEBh9wyulsWUlSxGm
simQP/eD4oj+J7gVidslIWS3xX5rz5ksRW6vLDHCpqmvtrtwRl3NvCdcGju5
mfCX+8zep731zxXViiiFeQnve9u+6GY51IG3K0u5UifOd0UbNGlkMMNotW3/
GMSS0gCXdFhQGX2xRwaJHJhSjK3eNuajQI05TA6wkx2w88tb1t/634Ew6LA/
GxchgvsSP0wXMMh4WniGc34R0J2IJ7PHiagPmiexxDvAQPwIfrykSFlHFHxx
7gDGsP6Wi3jr87+wiULPJh57ZDpnamOUXtCfATPhr51+8XCnM7NPQdwFR6C3
9ikupUnlt8LAGiZjbBZk2OkwYUGBqkPHtviwCsMCAOrfl9HiKn+kVDE6ImoU
2qu1WRiP26cX+1yZ5TvEBfgM5ssQI64qyU2M3QdkIX3usAv0+uqiwSl1I9Dz
IK1fIVGCXR7geeJKPttYDhuRsBIdaqQSK0+CtTlG//KaXRRq9Jd1XY9wKYcS
BBLkX2MrWiLruHQ24S6X4aGqj8IVjNy/7xjtzbVgULCUFsmHl5QUBZekExRI
zn4G3oUlzsftE809zK9GGIf/mvv56s5zeOcu+4vzpJWPETjA0hHnO5FFY4FV
kdEc1R7tdY6NeCNMB8MHa0H2/staTxSJCXaRwXEz8TNeTzJlXcvlm9RR1/hg
XmikBeBW9oSY7gQUlxb6pUUUTUSvp018k/Q/haFpD5m0hE7tZXP4sW2Bne2K
LImewhgu/0aMRKgjVT4gSUDAcuNW/VR6uY6olr5ZgZ95YS/Uz+yBvjn899yR
tIp1llf5Do0qHlS75PrBX+aT5K4YfPq0JeMiIHJ2mm+00hc6y26lVMOR0FTh
//HkEOXOn5yYB30iOFODBBsGnS2UUob/E93MpWbf9EF7hgdtzrK41AquNnJV
iOEYP5pIaH//UHbOMKAgiP8EAqjSiMbaqPLhmEXBl18kuD83PZg4Z4VXUL7n
mC9QfJCsa3zu6KBtSAp4yXRaOROuWxZk6uT1djgfczi7JbtcD6myhiIoyXQv
QZMCkO3hjg+M7Vv/n3wD3qfAeXBzNhwjQxxVAsTF8+x4LhLtKC71lDY4a9hF
j5P48LZgeWlF2HrNN2nH/YWEt6z6zWcu7/YU01ah0JSHlwwG/gA7eTduf0XE
7vNQN3SweQ5lPp8Z7S+WK5aRwpQs/q1miJr3ZOHmKdtIRsohae3iF+Mf6YkZ
CIO8aqsHsIEJbndWa0g/++2dDm5EXPx70r5Tyqarvd13aShHzw4eJU/6wbc1
t4VSdm+N4yOYUWsJi2aC34Tbc0f9WDvaQJslABurM8qGInERc/b9IbZ/OWqH
uJnUSmNRTOPcY3T2U184OF3UwOufbuMfpEYUHPBDjdiUz3sFrgIIChmNCOGc
/OU/nwxCliN81c2a/8Dtt8Kv1EFFMioJBycjACmvRKiWORtzRkmzPjmgL2kE
4vp4CM/zZqmGi6jniQLX1ro62ylAMzUQ3lZCXFW61wgZ37T3OpcAfsztc1Mk
SAgJhnn4sQbBuIVgsAj2Y0hm7Zvrlz7yTXjunhVcpdUX8qxNIhS2FYSCYMkU
Q1H1Frh0ysqbmay88sNrJNtCs49LGiP4+5KDLHXvuMo59kgZ3OMNhlaER09r
G7yQnG6UEBz91NRlzNNDmnKyw7+/2X7jE3xC6qnDIaDwtXmHFE7NTND49Gcn
nB7HhB7DMUyDVXuSiFLw/Kokrjcv5bVJX9Oj3Y568fWpO1hAuyRiQFD3rs/+
oWHG4LgB9hp+QRzCdDirqq00HcNvmZFrbUd14x08Z3OmSX0IbjUw4RjoTsfG
VBxCrdjh0srGb9K0RHi/PtQ3NGyYjBWeD1IsHQu3PXUvF4INaSDNOjRXN+2x
snZWUepLRMk8nS53+DoqH1Dpg4bhoIWQQ3NpCSAbjH8VlkcualD8hHFXcJ00
yuO8N4a2faRxl6Y5L+HdqiCthW8ykQ+rNlDiebfbphfewdYsHgtWj2Awxdax
OU2mjwMK/OXVUIEMMIbGnqiuXnAjUsfcTruT3AqyV/2TBEg2GVL7nAI3O8eD
9HHs4HbAv+0lALFdD8+YuCmoHXCWoU8gdWjo2qJp9J84zHbJWW+tRufCRw7M
N7T1cqtVjnbY69PVmoOkoEiiLfVXfnQZXJXjYviEM7gntIRCxwtKn7uZblcR
vVmrTtQGL00Gl/O3M4YXkpxPwjR3bNkjvy455L1m007ckrMSJGPYnvmS3G0W
gc6lBTJcZzgxy8xgHl8I06WdghFSS8IxaCKAr+U8W3PSA8IOQDGIdCv0RX66
Pi/1Qtt09ghk46h40vQ1Y/DM7beQIzM1loiETLDUNjOHmL335dPB528ClZ92
G5z7xY77iNWXqlLGRsX7mR5Xmz5sCfvsnR2nRKgAr9czZ8AbkA3PWyI5Yf1q
IsovxdKFsMTAgQKc1NVM1NVf4Tir5Pf1mG2yY8JeVGEy+zMg9vVnr2hQmBnf
BXQHRzq5c1eXczoYBCPBmgOxcSgPOoADcWptyCQBJGLCcAhdXzeRGo5VF3EX
TpuwTkZJ/LWm40VRCF904QZKw3f99ScacrjSBO2ftyjxGOMdvGA6ebmHy0Z4
jxvtK5qTsIyNwTqtymEYPbg9AC5cbZDjPCXBeQ6DCksypdnddh4ys2sSRtsI
sHhRAXS6KkPtAky6rBOODJRJgwO0jYUZHjaoNsLAoSvXMrP07Q/DWj98snQz
jjCziinrPmINeG2fKSLOOwpt7e08G4f9PPrvIG9PmiIvg9mS123jYiVAUExS
6xD1sVV2KN5RToSmwOGfKPjSLp0//ZF8cgnsXjYhLmLad2qMN+CFF2d+C5fo
OwPwTyu8YTP/G4Pq1l/HzQX7xgPW7sCpcsvK8VFltmEDwR3/hv8N7KbkQ34u
aLmUWmUXKwT7y9KSfMjSeZVwlCQySC5nNP73Fuph0Lb5DbB5DJoACUauokVp
QsvPzOdkbnnY+iwjvGU0nd+c6a9Fh6rdgGnxXtAHHW14zMWjTgpIf/Dh5t6B
5cl19uuQxMut3X1bpfJBl9K1Pht7AKHzCaCEvzcolCA7tI8LZ5HbZMFer42r
bQd6bTpteLWUVCuYxGkx7nBH2K8CFFnBIWLCObKZuHNDsSW9RqcvEUYECf6e
tHK2/idj5Y1/9F5wTKDHffDzmGKny12RtYqL5R2tLy3wTvPu29JF9X/s618A
pbt7C9Y3C+WZJz6N1nuM+xJC6PcXIgI+ZZUAgjFZbao8fOCs9uSpobrQbCNe
4CHevmjOxzYmwLcTOSnent6KnGQf/5ODBn884VvipHIeJB18kjBXoWQdKzdI
mThc0rZaYU7CZcvuVSzprx+vTym/dEJbBsUPxarC3hViLaJDhvM/Y/Eh/4E5
+AvGEz0fz9DG9snkvNopV0SmGfQ47sELSOx1+57KQdKYVbcWzjQxGKT9eZvb
qpdv3Ap6k9E35+Tiqh0JSTm60qmm5i17MB+rjaE8Wa0G2ahLOuzsTqmCS9UK
dcxbH/hzmvpFydHabpI4/vRFAFxlJjsL74t8iyd2Y+B1m7JA1+4kLl5J8pZH
+V4A/45l6DaFGTF8F0My+lTHcdPsnjbtd3KOID6yLfYcHYfN60GRBIbL9U8l
9YKerqsWWTnXN6i/FB4mLsnvwVSzLpNVHbbWHfPslKrofAFvh3r6LpStmsCc
y+Ck2OZ6wqEGPPmUYb2JEtw+bQEo9RziO6XIG+yr6bQ1WiFHup3vLdJykWAR
/wXMwBGvVDb+FTVvEevb5JxW03/uxuKd1R+pTIRQ1p/Q//2m8742temdUDOg
6l7c0STNnbVFIdCvmI4wifrBVcSMrnO+22bMYY8kjemqpB0uNYi3AnwCB2mA
GM0RErxLKl3VyESi3QOzjIQFQijRnydL3+gQijeJ2SliLyni4GdHVCU88CXH
KUvDCi8t9BEaHrcW4sZN0amTqOZHpgAzKNei+9ublloELSG6cWSl65FEdFt/
gQOKiey3PTY1DL0VkbCALd9eCqnbpiK/am+cFd7uV6dm29LgHwT5MiW3NAk3
LdbHhOSBR1Om1GgBTLX3jsUnWrP4aBuag2U920VF2a+sAw0L11RD2HTykw8f
7VsEPGUtC9B0gEDH7/AawOIe8qXtUD6HMZx88yJnlFBtEaIOzZxtnM6Ta9xh
6YBG800j6d7UfK7FJ32Ju8RAo9iDjq+s2bG7h9KPF2zrec9QzUhVF3xLdixV
/jppyRvp55o9xAmZt1PL+Bcd1L9rfptPfJqIof1cOClwwhcvQmrxSUjMLkzz
QsGBGvpwpkzIK5E7/TA5lln65IRNlvUpSDMi1oSUjwrDLw+Wys2zdDgPFAmd
Fmy6bSHJw1r8xIqklwO/BgF8ftTnEhKN+EItCPYhAQeLgCV01EsPEm2gW5LP
HSU3CEHOylVh5zYjm1QDIYEVk7A3LmHiDZ/vhksZk6Tfos1+/aV6FaiK8WiF
ui9Dv8mL4NHqVaLiVJUGWIgCx8U0v0snZkIyfyIHFpcDAl4MZLWiRBZNk73r
drKsdh+C7UmiGj3MhdzyL/gf76KDC1fvSoRsyFEyz5qfC4m1ICLeKKrxrou9
GLrCLnNW2spADvnX968QWiBDqM+YlKtoq/swzbZIEtgjt2XQscJbgSVKgE7d
ir7bqUGbSwl2tL90rG1XSwuP1Xx/J9hon1mfVcy/ClStXvuU9XjhcRT97lv6
raFr/7f8Qnw2gL3I1rs+gaHaP21o98OLZB4ZuaKR559HJSLYaYlGYU8MP0O2
//+BJHLcVsAU3OqmKBS46pwJDRGENYYnSogjgJJ8oNXpEW2MElodqzo8790q
OZZgBy+eiCh0W8L2ryt9aq2zQDof+9G26d8djdBJPqE8q2YyDWN7q/w1Bwuv
lm+WcvgrVq+zzuUtBbxLmx0fHam9xJeedNinE05R09Yz3Oj4ySbf4LUffvgJ
HWEqzcHAi3noyziYIWjh00DT8w12Bq93DW5wlNSaNWeZtsB3c3Gje3+xVAWI
yeUHXjLqr1KSdXBvgnY+sG+b2ZQ4+jWWOC64VlMU6GvqcXYKKQpISnAcfl1m
SXabc+mEQUnVq/xS1GUtL/bd7UF59/7uDFs7hYWcpyHO8ygtOm8biKVs2Kw7
omHUh0n/FqHX7DATlya3LgXkX9oOfKrX77qzJwodkVsBqjRoqlwcRxzVahhN
MoHYsmu1tYpaLK5LxyTHTyEPmwDEk9oJT/upjZUS7aUn/Eg3nnAreN7o5YV2
UT1ZDCVs2ifRBbFHNt9T3QUNC4XpuiX0IgtD+Y96f8qdtVc6ZIMz/051XzE8
c/AaSmC5oOpshv1eUikSehaPLYvTPCtY2lFVknT4fIKwv6sIgXpRLhXPiMkd
BMtQlvlVULCy9IUc5n6Flh0M5bFifPdsOx63EZgQ1zD3SW/9LzggoHNCqVGo
V+Fg68uofhIAfAMlnRXtyN9bWV4fdvFc05LqCrBRnssF/2lMC8PxI8KTzyIx
md1DmQEzRF6SpuLts24OoerfEaP8/oYBc577TMuu2Pu3Nkv98eWTXTZBlS55
Dai8LAh/bAwLxn+oPUGIfCnCmZXs0avfeVKad3HmwfFsDex5YtkA/YXpXuG5
JdWyDBzFBk5SktYOCKOjgR+N/3juAqXlyegzDQ0Wjdg1YiBDziSjvuqFehnk
F0gCpVkhU9hqcAAFn4pwq6VaV7is4oJriA9oLGWul1jFXfmS5LW0cz/h3Ql8
PLGUONrxVoKEmlcLUUarjVSKMDHgrAvgXJ5RWc61k/U/2EVur8eU2S0r0h9y
JO8Fmev6MgBRs/vx4ZRv3W4S262Npsg/qw18WITTL2eccuckK5zghA6lTtjN
Ruv6fXOvwYbQRC78kP2Frq3LmLdhni3pBQOL7kgekHdh4qj+Bn8RRatc6mYJ
kHEVDDHecxdcQmrrVEKKa3gJrfdEOD+oSTIdct/hMfIk1/Kkj4K9QiQkzZPg
utacXHB3vAqWISUvegqYtboeoIS5f3cafYEk+g47V14w2xzsKB/qF/YPjkGt
cZ4wIYFXud/ujcjgyrzEvbOTujg/JamYfR9JAp/UCF/MKA/rF/Pd+Vvzw3IY
8r+Uy9kP24yLNGjEXkmJ2wsg+9+OeKv+vvGjimmSyMEGry5Ixp9E/uFmtj0B
quWAigzTQtDgdo0it3ChS+V6V4pw5olTB8y9vttDOKzbEdZGMJcRtxwmzJI1
xFMPLVlymLNs44T/wUoNNpFw7XqXhe9ft8sDqJedYVzTumWt7qXZmU46NnH6
CAFBZMQMWhRVmUhfGP5gOTrwf6IMEsFasVx9HAWhaWZy85+IrQIvNZDieOSg
V0YR0rZCrX5uep2R9LBPMkkUVH9KJcayFNjrKnIBmk/UxHEncfNoiIj8YFOP
zF9qBfFgLmyMzAfgA2xxDX+f/Xoq8NQgkRxkRLRJxlp9oBcXLT9hiy2hJiC1
ezV0OiAP9YZ1WpzvlKGo/p6XRoUrphQBkrSiGF0fO4zEzpHkRf3fr+ysJUjf
xkvgJy+4tiL4z6UucYLOR3OmepHAxI60xBc65WsuYZoCZptI2cmJXu5RfILP
uZ5DoxVF7j21zHqyTY3M01zS+KCG27LzTnEjQvhhz981wR0BxO+xm43SBGjT
L7f48JOVgVT3BDQaYOE5r1dcL+/p50UVXxVc+LIfy5VYum+qnIUBPrENw3eo
8tcoN0yg244ICsZBgFQl/GuOv172EFMQba4bkSRhr+g6q/zGbbD6zrwM9MXM
x2ma4AWCccenPn0zMioaeoSWqmm8BxklUMJZIdFEBiW9q4+8k50ouqTLy+IN
L6RZoNiPEVom5ECWn1aafAWzVaiYULI4CzoiWtz0TCk4bhTFxXBIM3CM6G5D
SRHo7y87Yynfi0CnIRrrZuzhtLCK09hBrFnQmP5t4Q/4asEJEfG0borVbc0F
F5axjjlYKlCeb0ybBIGKSXKm0V0tMv9OzDlGAWnTW7uQOqEDrY5+amFrsNi1
IYpBY71iJ7d0e4OVwqJeAC06/tyW+sGTI6B63Vtp3CwvxDNsqFV6t/JG/m0y
Xyr67CLD6BIu1UT0F7G0O2fw1CcfwG9YS2q69MbNxWtc5jFJivNJOClEFHrQ
xN5ox20XIY9/XgU8iF4D1ltzZ+nbsOblbEZK10qcuCzbvyU1/sEzheiUFlZs
W4c3GMMhctrVkuyC2Pc1MvPbp7O3i8+4fOMFe8WX9sAtU+/BhDZL+moim5sm
u8Fi4J639IQrJJDX9GqoLUkLZ/TmH0rCd28Roh6qMEhHKgQzpv5mLhEl3XBv
6pVTE02AA/EREXYPeuy0EHJfC2kWEuFzF3N5jCoM3PvyQFpRwv/xqlI0lfzg
mfMyH92XxIz/cg8/oQ3wH0+IWK62erYVWq1AZJZvMvTEahFB3xFNy1zVmved
aUcN2mXQf2LBxGiP5mX9a+hAOCvm5en5cd7VBix+j8QMQW2JugAmlxFYOe9F
EvCK9FwH63Sqj5s1kxXXIxDnsRGzIhiL09xwP4Fs0bq9T23PaPv9Y6fn9B4J
wN8582u6mdJov3UXQkkgf1KkTBpePCDlpWA6+ScMy3+JPmy336uQAgnUt6iE
ovRRJmmPYuYkDtOqiUPcak04KgQh8H138bmxP9OB26g/X9MjSseFUqktXpZi
lGsmm+TphgcCcll37daKkl/qDevFdfG2iFYWhX+VB02OLoGNR5LVrDxUXVVy
m8gn6u3QBscj2jaz0co88pAeqcJoJX7X7OD+IxTetWLTT8oxlj2CR5MSw5aQ
z5ThuVFUa7ryNbu5lV94k06/QoYCuxgjHIbo9Y0pHx2ludidoxlJNJITVZkO
sfrvLhQRzy6t7mom4CpJfF0QWDFZRd532r2/r4RXtl++/pQkBo9kvYws4olX
WhPrMIHJIgeBkDA3V/KjJw0/DuhV+6vtSLboYTEfgNxaKl6tkU4CJEL3J/0c
hSwza9j+VMGiG93Pd2NLQs63F0XgGIR7dZtPh40ZXGJihZKPJvonVphVAuzg
SGBGx81YCu4Px1LTUICIey2lfe2XvO17XpOOlg0cXOEeAHeRxKvD/RYFQf6j
xcA5pAayh0LBeSq8187NDCYs4HDfiol7CXJhSR8ZKhbFr2c754XtJy0QjSaR
O7BkmS8qJFCwCvAwbscXRlSu4EUPiXTY/O3fcnNSNc5tRMxNMVY3l2ErYLCS
JPYwNi6meqigZh8sj8PQzPfeELvGdWRmWxg6u5e6VFavV7t+BVQnSMrnrz9U
4/nl0qQJaQJL1rimC2vsHYtfsmWp7jwuru6pfykQB9KGrUBCGyghhT7268Lo
DpNQKLD4+pNMXPcD5XQ0Gb/iza/OzNuu0VOZ5wfsoWlNyTCiTx7RywjQ/1om
0Kxco0wGf0gz5ooF+AvKPhfxjhGElUK1bhyPdh7yQUBmJfwkGISEKqZG+fB4
zJiSxSlihfVtGcQT2jrwlklN/2diC78GumsdwbQuFl4wUwuqDtRP/R1QJTvT
q47myJSQo9TX8EW4kNEEp2qvuJicwYcG+xYzn5pvCIS5wrP0RUUpjO4ILK5a
yArDCDyOW7HLMK1BIqkaPWg5KWhRqh/0fUm4c+WR0GMVGCIBRoIc0Ltf+QBn
IQ7WzZD+R9HSQ4JScFxYmiEakjbS5iyk91lJ0GWeaP4rb1V+Bk71gLV4GwFX
aJtjJHrcQ+dVC2hEZPYRoZZHCpDBti95RGbHt6WBXY3cITptkVmRfKD1qBws
SNz717FwmsrBid5eAEej4yOwlFPcwefMhFoBaEVXtPZeDqAytN2aWyowZXP4
4H2OXvMp2hYMnloj0zTNsF8e8Zp6L9xUjGTb98dy9dWI0Dn1qLyibw2DvVQp
5JXb5CawPSLNKst66SPfZq/ztQAFoRSSw9PxdKFcsqWHZ1MV34SvUhETIMpu
NBl3XzLvU3245SHUVFjrtmhp+CoG5bna6usLw+EhubcyhU64tPF+ldRyVjPE
W2PyleGs2jC6vGar6AydrZWF4c8HJTekwuceUNI6Uoyi39Bat0bzawtNJut4
D4MGhmPdRSGIWbYf+lyfNYTmpPjq/ik1p+prFtrT6SRpZb6IZ0kABk7ean9M
mScOv6lofYbAQVUYgrh6rS7cIAv4A3rrPsW3+QGMXe+f/GkXKwWLIJghUjwI
zXV8jLl+uxlk1eplKBEtEZB7tGwEF33wzEvaDZ5f5CWq9q35tc+6gHR19Bls
OswEXiOiWL68/4SZwPQTbOL7RFk5VP01sQu1UQQHa5ewzAPmHwW0ya6k6Fn8
/xsUXoOhtj5sCev+Xi0ayfKwu6FgQJbruw+ttcIMTC87hOIBl+ezOErrj+kr
hDHyejz20M6rW8gKLO8ip1XkGxtNnSIClcDtHU2zck+a/RpJY/PWFujrzDiK
KvUddZoYfQv4miiZY2FNJbEYrZGnrofAAE0h68NJiZdlYxQI+n97De0Pv+ur
508ry+hP/rVc0tVntyqt9tH/P7zY7T4Gl2Rw/rTjIXCnTzq0Asonve2FQ9Bt
NkD0CJFYUKcwAJN3mbp02JK8+v3kEpHUoLAFHC//agrGzLkFgXGZtsW7iV2C
RWB0TiGPt9Uwts3iTUYk8dO9HAtQMboSRbB006CopotXeEVzcrRPox5kZRN9
yP6Na/xgymklQSCmSmbYzBxIrcHrOsSez0DcBA3KVfyhxvyuRd6de7dDT3Qz
JksVOcQAMRsborTpn6DCM/RNBtZvFf698SYpUie5YxYu0qrwLDlaPvZwJoN2
TTcqC2ySEdRD1CZK6i+XcSjeouqzyYQq5/guXOqYKB4Z/NGwbx3MPEmCfHRA
4EjAQljHcl0NEUuBAV/EqGvZNJ+HjRdTVIyjMsTNKCq2APCVRWkxz3vCgk3V
CtOkRdS6ruHkDXbenTVeg4U89qDgYMzvPjJJWVgda/ybsuAv4G0ZchpEDzI7
MI88PNz8x01qjgthAUjAxQY47FjfFAEZcydxo/yiCjlvzRUSaktA09OU6MNe
/T0pIUcyupxy19ORuKfunOdp/ZcJA+DaXsQSeFoO6XL80+R/E5qFzlCp6adz
GqH1ivmJIJ42Q6s5VliZf+QagZBqZS8ypJfnkxJB930iD5KrM1H++L4BwVkq
oWGj5pCjh/BGPMwKYFjodJPMsnZmjZ5Izl/rZK+fX7scUOUg/0uzKOgdvqFo
m1Eb6Wxedjl4Yf3B0cPc5ldgOvgZ8EfkX2JvmLLsWqhyz/8VzVNVMKwlUw7H
8gKSGfkKMeTLP1wierSYmfDE15HzS8EeIXevlwjfve6v5ttXjlYgNf146R/5
bbdORSVIPSyhUdZl+id6m1XHl+HCfQVzbUvFqk6DDtsU2QvJf+txfc8dSNu2
OULAPTkdU8TE+qmyZPrDIFhRHyHIAh23oU/dMKGS4ExEOiOIQ8x0VeWbw4n7
urTIyJ3semzylrT07P9UFLVYknUYM6/wAvEcnLy97StCHn6Sp7iWk35IWT+C
ySnH2ZOJ7XhtuAurMjeXtxl4AE++i4yB6KiWBy51zkHDq87imS/TE2kJU4fi
8RT77SHvMMF/Hw9w0Nn7ysLmjUV5lc28BWgiVfR9D+lqeNH1wrrqPeuwMrgO
QoH0WBMijv/zXpyNANctF2t9GxqG8ivkWJYJrPM/xsoWWtwkEPAhkxTUyuKL
juERol5ZYE7Khs7PWFgPF82ClUDuV7RRDlskU9RV8hfLsrUeVBKA14RYh8I/
BGoltilcXX8cLG/QK4KTTgckiqYtwdw/pCTPp8eP4NH1YWW7kJ0a5I2aT7xG
SvNhEgaKE/WePTLxaOHspfe1qokya8sDTwBqlFF7Z/IxZPtOUferq/swEacX
nDZiRVRWwjyPzbxrnb6dHL/iBWGjYj5ZYQrDqRWGgmnxlsEZMear7aT1V3e/
gAhtmh50yqR0zA2rWN0BUQvJIZKWK36wZggnVYTWSf1h0iy/UavbSVvYCoKA
TJwzmzkyI5D3d/OsNjunpAqAe904L4882qq+5QQfWOobhJ7KvIB/W7h2IBal
w08IdrRYJFF3Uoy797ZvxHaPqaiJBgXYnrQyg2K9Pmay1vKAq42znC6i3fRS
WPAm5oKL6ddw76NYmRwjhILS1J2UPID8dEPbPs2EVq/1KoHejnRF0GYhVL8y
Sko0+pyiCDkMELpYE3pFn4yJP8zVv9wHnGRYUPP9AEvBcolXyGBRF7NnN8DW
yP3ENqWci0xwEM2gOI1VyLNp8ENylbmP1PchFiQGgzd3jzYvbZqSiFI2ncfr
lxAve2RYhAhYL1jg3pPL4ibimCfLabNFOKbi9glWpS3m6I2/UsQkeHg5XAd0
7cT/Ok4P/zAPoOyTNZ4atZabYeNJIC2/aCkDfApmy2i+/qT7CT/3Rn3bC9f1
bBACua28lWDdOGaygI6jBr0pFbWL4H3RYJLJ/uue8GKgpP9BwTXl8bmTP8lm
iRJvXVjxTIS2alrj/PKbF65zMk5jN2JVc8zCb7+bz29cLqGt3OZpm3dy5G5R
iHwSJ10ODc5hkcP/XZRuDGfMaJnkdVcMNOYPN09IOgedDxeNrdzRmYG+JWMk
+jPG0ZzVDUkds3BcN++alx51rDm2K45Zrf32xeklqJw8Jn6i6l051v6HwuZe
vv3zMLAZ977jLKWaUmoZC4lDDSK4j6IhSttIh/TsXj32O/Y/fZA2FrKAmoHR
xTtLgTtQYsmMQ5uBB1P4olqnKKkIhFOsSkUr/QzwMgZoBtG/BTwZoF88iAla
NevuMVLWsyXBsjGFKX5N1hJVqH2ccLh/PqaU0+PwIbSlXYuhnkHqwMfTAHnH
CUZEDuKVnXtDVUFb3EmPE0Fbc6u40nkuIuZiTw+gMXkiCdk/Ndv48mmchAt3
c55eHoFPBXil4b6FXKEdEe7L54GbwMLZyVPBLbk1pbmN8m/WahwaV4IOc3Tz
uTyx10ijysHGm0qQSNY0YRwOF1Ni/UrELQfyE5oGLaABCM+If1VcZ4gEStuP
3XUPtKe7nklUxqAKpr7Oye09pgeDKc6XsER9feHeG/tuXsJZrGW5ZJ8x7vnY
LOyQd62abkKoyXGE8OiiwE5ijNyIjipEoqK4p5IjNGuAmS+fmvBqGor9n575
iay9n7VGt2/ucwiJPfdQg3F4c10nCadguiYgbf3+9twq0M/+CTxkjPrjFgbu
v1JeHXictE3SFju5sF+wdcosINR8Vr9eRagFRweRpbLiL2aEqk25mbXjoaFz
Z6zL+L0ObQ8uVLF8wJ/ZRjaNOjBuSzy1n0UIvCjlOneNJlhV9KTJ2SYlcL8W
/t41jY0UhBWNps+CD37N/bN8GimJHags5AgkbMwbFxaPWyw8GBvjANMBnVy9
/auRshDKNk30bbYpUUfMemvcN+UcI2ekafW9sv6ma0Vzy4crUxgKoZOzrvEY
0bvzCBoC6QVPs/jjR/lEmiGJ8LdxKz7Sdy/UZTaW7iP5Ta5EiK9J3+PQxpqn
AcnccGmaH8mg9NDZ14tEu1iUkMZbYINw6UHyvqB+X13rqiUQ/atkdIhr1sn6
woyDNeymvBki/s4MPhtEGuUP/rWkYNM3khZwAN8henOibNDP+h3Ogs++ZM07
D4A2crTSGa3bbSxfhyIMnxSzq+BvXnIeHadowREFAUCN6ccWZbPKZVz6LFPZ
AFEmjVMCtdBPuyuk3o9Ob0knVhRNbDhL6Yu//XkD0BLcOGs5PfkyuwLMpIdF
8IvPDRiih+Jbm4cBh3huntt8L6aGyKx3iRY7MPrVne63512XyZ94TB1zfKk7
cmrNkLzCl5X9Ufe0yqX/H4PY6XvEirtGxcO/ipgA8NSfXGOea/HCImWKB9kF
Q8Pz6rPHHONSVAH2IKSI0LUXQ8DL7IOU5Md19igQBRAWmIkjWrNGeTuEqEsV
q2dhuaZhkyLn6P+s4FEatvsnUVDnJ4AM1OtzkEIU5SGq3Bi3+AdXlW7CNi92
ne0gW+VcQyyKgADq6uA8DNrhyiNc9RlApWLvjsn4VFIgi67ijc3Hh3Run2+g
RoKOQMcP58FUDBWKkOgjm8kXIUBv+Hq9trqQgOvhGsGfudwMflRaGuNlZApt
yM4OdoL3QqFPBjQFjqzvnByJAYaM90OJDaxV3iVpxeEuws146oYK3w3zDYkO
9XNwaXFTCoV/mf07cKF4b80ndiUbOLoLh2yC9NCAZcdPeis06C6V748s2dwW
nGb+mbCsuofyKjEb9tNDytWOtzpqy3WJvaxhoUiqARn+Hufi+RN3XzJCmsXV
PN0MgioijXEkSkLuovOcdD2uHC77L7AkYDsh6rWfAolH19JOcSLZhBKspn2W
8GZVoSPJWsZKq7+nMwoQYkQOQkt82XaIyVL7vnEJlH7rTdmu6u29y7BEef71
L7EeLETA6saxBFIdrO6/2QA3OdinPXeXS36k/0WFrYNRTWgrLPhpqzjahH68
sOMX5phfzVeENlsU5jwEXqNb8BF1EYLoGwhUBhDjCJlxy8hTUepGRYejC+vK
VihYIjMn9+oUmgV9Ts6DRfzx1iYFUQ2j27uvVU8vS35Ie2OvgfsbDPkgnTqY
F8uTG85cH2OQ9jFamLN7882DK2P7nYtB83CCFTpOQBHVnvFuMIb5UveDk8ht
xHwvsFjZmvYQAWNIvuNosv39cfmEH62YEMCUjOEf/0gPwNdBpWZPdMhr1YCN
2ocI7UPHlny3WmeNZ7iPF2DctLQ/wvZC+1yt2fnmQXV5Rz4phD+fQTczyDyH
Ynqf8s3+8eIZpYd6FBzDrFekDKcDq1AQRXDqbkOU8yEj5TWaKtt8EeMSxmc6
fnvfplIbA0JC1W4C1TpGBwYQnE6yvMSxEX3ljWN6yBWpHE2fzAKzl5n+/A0/
Q4hx1Gbr59f85nzFyhhOEvHZHuHEO9ZOzbb11X7ElZqBZBW0mEBeukxPH+Zp
/ID/UGC/k7zD5DOzwW/jaOxEKjM9QxJaCcO4aTn3jHXXmKqN3pqpBFHsZjqP
LwQvHnBt2/xeOde/Cajqmc7ZXPzYobMMoTTr72F2sB73L8sO11Io2Ko9s+qI
PdAPPR0eySRwP8bSqs5J58YQo53ZBqUTRtR0r9W5igpSwDOQkWn8akEosAlq
sGK0PtBmlNKkUHCdMcYBnxCpfDWOpQ0rDQiBTyG/p1WjVDE46amKeJNzZCgG
0ko6SIZ/bhjDQ386ODPbR6zDY9bA238gc/U3Do40OXOD83C7ZrUIgm14kDVw
tiOVD/eQZp2fY7HiPpETZ9C592Ku4vZaJnq/vl6DwZvFwhFHkcTim3FjTbXD
GtQvc6unDKDMjYMvuBt+/MrlHUcF576qc02E9NTjng2KXZfsuCQhx37XRhFc
btBVoGTCy9fIEg/xeiFNaQF7Be8oZ6R7Uj6lCfkncGZLJyjR+zLePREpiRlX
0LLmmeCGmD0oxr9GJvzecgJUaLvZg199hwb5Ji0VtVli2k3r3YIi4Y4wau/m
Dj62+HQm0cGEduJGTIJBmSXRjuS791Mu48NkM5w1mR5cZekZxFFTSFLSrewB
dUZMAVvZ8i8o4vjph0YwLMvtsRUhXLBoPt9moTDz2lzRWuOwZxxab7gumrF8
mXSTlJ9qYJMwnrGe/UyN4A+8ZGgVWqmxxwsCe9MLRMWihOI0tAWha9fWWDSS
60WsOi/UT1dpkMBL6mOpyOh7tUBplUUfbGQ0bRAPzylr1HtItRJ1pjUeKGwH
DUhRf2FSghXW9/Q7NUfwFw2cwjTdtT3Qd5DQOgFWMYgMJZwuTRvF02si53Cb
ykKIg4OB6XJIQRl5ud+iLal4mXumqkuR/+0duA9Makg3RES75snNTLGJC6U2
TwuQeUjl0x5tqvDwfqclEg7HQysL5Vf4SzSv2aXcU/TURdePojz7NcK2wbVx
2/KjcEtfQPseI+6aapqCB6bn+FCj8FVnB9Bgi08tMMUiYZAGuhU/X2gLVXTa
5kxQW9musii6Jtq1jqs67ZrbXSWNrslfQ89C8ofroBqsl3OOAgcAcCh3aB+c
CY2TsIBADQCILuqsXG3RzlBAIxjmEhfm1R1lcduzCLeAsdnTdZS09GBF3NMj
0zfwhxFLvtKXdiS7mj/ICpaKp+/UC9AM6645glly5z4gRfcoSp9YIceqcJUh
ZH6LwoJiYSeOdkGpYyb9fmz7jahEGBvTURpcu6JXRVD1nwRA12x7eNfMn1Nl
rE80sCJOoU08GR80KzLZTymT/izOI3PL48W6XOI5eERpqU6WMDV7Q+YIWH/b
YC/nSFQjBeDYHLyD3z5p4kuRdgo1bP6aLStUmMjYsW+i5YI80E9s9cfaNVsc
aveW5JkJaHLuWxHqWNYcjupCgAjDj6RnJm+x56oYJwymDK3OCEaqJoOhpR7+
lvzaOMjbki7CnlnL767zVuq09GjYzuGEkqxOM3WdDISd/D27z8bxcDwCZayX
ziwW7171SAqgVTds8lzMMrtPaAItFbKQ256MAp1oVLxDhim9MlgIERDqf/hT
az0DuMCE4ZaRAEX+LvlIgmrKcHfL/Y0M5YNtvWPK3fRT3YSG9FZkDKAikjkl
CwwTLhGzelAKNaHDF5PbXgXnklH4rkAVGCIYwfZn42wt3ABF9vufMpTljRYn
TvgKmd1oPNFqKIcbsV1oS1nKTgBLz0aCNx17UvLYP3KEk/aLVlhcd25zH7m6
U2rPYjsh0BrzEVDrJk4+nz/dbcyU4YmgNRLn2yXFdnPjno1dHHZ4mCXxQ1en
z32377cOHM1rcVnPj1t3oFL3MkNeGQYwIZlEwm2B51neeitg6cTkAmx48nVb
u67dwY8YCOLgeMYncMzv/g0zMA+pvFpW398WbGGQY8cnOcZaD4dPI+RlpYbm
PcbuMBA7x0zCsUBRYWmmL2lVpbbigNO1wdgSs5uE9RlMCBzAtEr8wcnDyjUi
JHU7xMSf742xuQ35kesIsRVjmQeJBjTXWHp5z7s6cqAKr1YlmIdhFKAwW0L/
KGDJJm/D3L0cEG3pZWvdCMUimMiDdBEobCL+/F8L0FmFm5b/RL71BzjCMBC3
tmn2DwvJGmXYPkQ3pR7XyVp0okSpOgg/GxuXLhSYiYR4DFfLPKyxMUW/Ey8F
Sqwu+SoE8NRJIXwg4G8/R5nxpxacSrcFw5tfDgeasGgjyIHpMhv+pFdxjhKj
Sd4j6U/PndRQkTYb6L67liu5bsqLNqZFIsw3GBuujytoLCxbRAOdpZDMx4d1
M/48QxseaHv3X0fvODGHaqCml419M7mvSJNDt1w8AXB5VTUsCUeyMnmnPdoV
s0oZCzhGhP6/ewfnrmejZcYZ0vAyfoTs0Gv9NReY18CNtqZz54ugNt6oN78r
lXQR6tn9NROyKXL4/QjWMkAmDazwnPok8eXqTZylaZrayR0V1Oj8ZxVfxFFa
Q2wcyi7GzAZgeWW5X6Iin2m85txeVWSj1ME5tALNbiU3UDWwT6MethcE3UVn
K+J+lD9AE6A09J8dmnGshMgxzJcnCFNdFXKBu9EG8011cT2e72zBEbQ/RE6f
sEa7uv1h3T52KoSKjLmJJkU2faMWG2ViEC37kghoKDmA3RrnXTfxVcUEIzye
HChPqtWlriH6V6AQpedAJtaEubAgC2HthlTYa2b8Q4/R5G/jTg465OWgQkmS
bi5Nd/3J0GtL5jgFFah3ykGATqgFAEtxhfLhxJjHt6SeDjMKP1LM0CqTVwNY
fBPDshQxDZTqBCLumey4YqqkmuZiU9AJz/mft/8FjqzOjzBZw3iNj9DNDj9P
gB0rnNJ1fJgf5czGEz4Rer/IZQ2uAEvJZ9Mi8OEt6p67Px3mxF52AotAmRFT
HJt27rZvj8Ij1nfvP25TwDOhnW6cRFWyQb2ykxDoDmuq/g3qn5nXjmgGELDG
qxUkedom8DAsBL8AF9/PS+qNAhMLxv+nI+Psdq0HGy8c95Q+TAxP310HPWdt
07FAveAWi6cV9ZrkxLIk9OjNGE4WCoH4Lf92naL0Df0CiyOVeEkfN+l6w65g
0/69MviNBb1Q3OJVilzsmxXLaPMrqSCecSFDTqt/TAzLRYBfubcCAsy+CN6R
YLisk44B4pxQug2Vaxhq869yeMdaYNYW4si4LiuLu3jc+CQiimF2Gau5feIB
gqscW3iY8h+n1FHghLPs6oxqBlOeSmA6z//tdOUyury+jtamjLlJSF94Er3E
s1om4hIDl/6mF8txl0dBVIBeG4GLVrDicFEX7/pLXCBar8/Ckiz6t2kJMU8X
/C7ZPcDlP+To4/AI4xeM6uQSUzVQPWpTqpw6shH6836HnQzS8OOjpA3xjH1U
z9Fj2EwQbaGMFlFWvpcVrcGyErkBx1B24uho6Y1Wm1kcNANyrLj8CS8TDAN5
ULCaehv0cIb8EqG4N6k9bHTXzjvKXtePc2xxynKzKnepi8YAGGllTqaV5oyw
00qsEL38nm40CJLhVqATVXC7QdXLuXmchVbgHO1DJCrfWpFtoQwnECM+S0aK
ef0qGSrum+wJ9OandmYfXwVSy5hTZRbK5TaPLIr8Y1FKwtbFhNFBtAKzNIqL
RJQsns+Y3OCcQPL7sP9slu8hbM44tpkr4XiqPVRqUZNoaOhnoxczO8rA6CEy
MyMwm9DPoCsW3PH90uYdevXTv+aVodygR6g41KYGpXZKOdjEboXq+cdqGUOd
7dJhNpaUMDNv7WAf0c+dk0snIoVP8WkFTnlyZUIcEFu3sjjsZcvPUSkodboI
J1CWa3N6Cvqwpv88L8AmTlU0wgKoHNoohAdXuJ68DQ39USX0HqX5es+F2fta
FaDZ9M9/HMWVdTSH1kXwPcNZ/bzSAmiZhhXmbMPaQxVOe2qw95CtVGq4iVcX
5xpKQrXDC+XiLlfwRiKMjkfMYSgwmZYtOlveaEoExjF1Sfz8T0Lt84uxaT/s
HTLpyFzlrY4VSrRpgRWxAauZkqpxlvLmfViYe6M2atEYW4q2j1EwIV+HRuBA
B2oAXRSYVelrjBwIxtzji0ks3Q7vNINoo7eIGBtyfGD8GlRLcbEvfj5tbgd6
Q+9rmlSYGMfCTaN2GsgOVAJtuEA5JKJbDFxgu4GlD9ocTSRT9ehIpmbik29R
zir6B/LCoLwZNUeW16z65smDPfSfHknHK95Eug9OL+2c91mD+b/l6uw4UUtz
EMjUrbEXyMA/+mEJrZLP//a5RqpJOexEKeSt7lGIcyn55zoiYxj4XLPjDgJb
8XomS6A36pT0EhoO07eGvhHiak+K9WkzyocGZRvA94MqA3i58MSN8sytzsdf
+iQHSTw5uuS/iM4riz/XkA2vqjE8ML3FmJcleGprR+TCSN+uhlQ1BEaitSxL
snVhhSQKTiMQIqrkum13xr4GlppQXQ7pWtgkjOw2HkWHJgTEPe4X1iTnDKHn
q8swg5GxMr8zCXzrkJeuyVOyielqlIIFRw+XajvC0/lLqZXjo8yi3HBOBQvl
TLJllneIaRFpgTrpDFwnpy46ST/stzr1c646qXIQHC3yeZRd/4IO6LeLhalM
yVk6T9u6cTHIe0yJ0dOY6JX1xJqw/a0y4maZnCSpp7gFka6Ve+aDWFGXw/RU
SBVaMjFqz+VO9GnpUXMplLTYGm9Hp8jV/UpiZT9AD8ozvbd8Uat9OQdzsUum
FdDABiihXYsFgGBmoQ/4GZ1svSe4aG0KT0U4lcblX4cvh0NGC8LhPHbwjElU
N23Ukh3j+VI9egk4/IlvrKtC2eMl4Nk+Ok9VEZYxV7iZlUfMl9CX/VT/es+0
9cdgor7zY3fTOlp2vTi4iNiOP7EGlVc2wuua8KVxTJc3LSZ/gAkRqcEDu9Cl
0N/3EvwcEl563mS5DKfMKJjOQcEMseBO0o1Rbp3ygUmVtxtXOZH76c4eXNsX
s8NwJzClwclwjGKa4zzpXt5sC1P9fW0aPV55U0YR1n4cN9NBXtaUqJuf0zil
vOtmbGm1VK2TLP0I0WrsoImm5W8Asz5YUTrgHyByYJFE17+sbrGKXCnC5PQw
Ky5TPCeIFlGHd1SSvBPfb9OSThk40/2Va7xJFOupZVpeBoc3TDieB9KVay5u
U+Fk+PTeGjsXPJz8HqfjmHq1A7yf2lenov7FFlFA8v8+rSLLwBeFd7w0ANJ7
c59ZCYEyPv6YY89T0Zena9W4cWonuTENl3643aDe9r3TJ9JqAFSKujtxi9vO
tWvbj+CcbcphwXNBUmOLZDuuj+lhXm/kS42qpU7kM6YRdSn97wfu70HAqnYG
5J+uB29i+f/5DuQY7rfCU2iSZDLdozgyaT3KKvhcN7Ei3JDL4oPG132nG0KN
kix0NFc+z/IgcBxmP8xhI3zDDCoIcJQ0p0w7nvSUKv4cTJ+NO4rW4uHTM1q9
BsFtSn43VWHSMLn+WkPa841Eriyb1BQ+06lzzD80aZT7u32BKzt9TpSQWT2I
AvapH5A4O5exLshpJvznBltZahiPGRV5UAcgluHeEdUCwUxHD8H2k9kssKrg
blQtdfRPn53xZtHn1dssgIzxnT2bsgr6phiy06AO7wbkUGRThV1LcesW7RBu
PTAFGDEkf8Wogo8K2/ayJ5b1CAqbHmjM/jD3SZfl7yca1LI9oYckxE96+2w6
bguS4I9IG2yEfETRkX2pKbGVwJcEV7ecpJCdf9zPE2OPBd0T601PzgVq4KDc
xVyYJq/fYXR3wMUsdWhFXS6YIOmb5mNKvllPK+A5RlQzyPcY0ZyjEt+jEo/V
rd5KcOYOVn6BhGK8y8FWE3x48afZmuEJg80zbreETMxaH1fDhnV8UT+mr6Yf
tStmtZr9Mc8AOLxGpjIJcfe37e6y03UTFOnIOXmLEIWz9953RIGcJuKZGnlS
TrmXH7vWQkQAatyIlkDOgDvePT94eWieRSbtyCiZGv5XHxbTZn4yUu4uU6uL
HDO69mKK5y64/sPjKf+yWpOPdYF5M2KVb1o5UnULE16X+sfAtEEa9pnzB6we
DoS0I+CobAbqY+KSVcFr13OJZNga6n51kYAty0YqVsq3b3+Wuh/nlt42T+44
5Xvk7WWJ05ePqd7x+7wfA8lwRF5GM2yLSvNRcqW0BU6zEPCopmvYxkErKotL
srCermDEOOmXZbQIC5VUui78dMJg+3FOtakBgD2KlPNLtNcPzqRpWZ+EO/f9
xYFHtZKUDcHzHlAVGdeIZZvmRGPzn+OucsCtk44sB6C60ClwKZ80aCLibKIQ
FRRCT5KS2//+bhkCki26+9RSkiEdsrr16YtSGE3XyiM/dhgtn1S0iWkJkXqh
49NTW5DMQ+bXKdrPjGzBnp+DqKKpdaHZIEy+cVt9OBSzd8DcjW96dad4i6jR
Olb6d7C8dmqY2dL6NB2j11IkHsuyPg+vIHdsvKR4LOvmx2lwbm+KZBv2tfFQ
LuiV9KV4FQYuyYPsqA0UYBW+TME0uhDcGVqIAV+YFdyMOW9a0rGPAer+I+il
DN0TtRMqWfy5wa48S7WLvgdgCXGxXSBryp3L/d3ZlGeuEIWpmq+9ifcwfDso
O9Q38asy++56krkmGL7bmltHYebEXEPDu/wxs99unGVTTg1ojDw+5w9F0tv6
+zaVzGzE/pgbcmg8DcUIF/sdiaTx5NDM/bR+YSGgrE/EOwMKAODznArrinKx
IWi4tAOAEwJlAefq2sISiuBQHL9kpjJ0QwRhIqP9KkLqkjSQzWDdRHpuSlQS
rgqOxeljOg3IqE35ZeaQjYQXuRTjTnhD/LI0cKhBZa3eomlsw0gUCMjP+BMT
aHnSQwzqFTuqV361WLgEQZDyHbLCtmqpXxLCnwUYPTkesWmFimwgYZZZW7nK
fTdKx3SKdUugUC4mcuenBnoy028Lm/foXsXN2eVKKJJie75B21owCUUgJgsA
m3JX6aAjENPJaw2QA+mCyngWd8rgock88lvmx4bs/uZIN+/1MRGaIy4vebT+
t0CjwP7R86UUDZoZ0oJwyfqLKcaamSvPYg7pFjoBXWYLknMbxFa4Fz2UJMk+
Z4rfi4LAxVcr84HUF+N73SbNu/eTN0Tp00v+yqV47q3PFgAHc3nU/mWJUlkU
kHUhm0Yl6W7qmKi1sFs3D7AINC9PJZ0QrJMwCmZnaMa3Xnv0oIOaz5JrjFg6
R3GQ/E8yPtDrgzV4QoPk+jUQMjcrAHkRoMHLfEiq+zTjFBWklGcMs7fYtEgb
0P3MgJ33hclr2NB05bkOox2AB2oGQFGptsvVxNo/Epip8cbymFWkHJ8f2ue0
PtNV6MV2SHIpYq9qbSFmqAhh8BBitRLg5BRdL0vxfIHgUb1EzWv6gGEYNTkk
G5njsMnaBQ4GRvJyqA3z1esNKZGILMgGZzSRL2Y98WSdKWSn8ETGJWXWouUu
V+tPLxkn4S4t80W3sFujRnwC89YCcv0Nkcx0ReD7WzCAvh8A5S0WmdMdosC2
gDCWeJuqDm8iTFussOpkSjZd0z4mB6kMJczBoEXkjXWumBoXELMmVJJaaCVk
XELBQLkJZUOss/8TgDMlvZKbGm7LviuCi25M1UNW60SSjytXqmjrCHbvZYd6
glmueGN/urepl/9z+5+zkj+TmPnPd8xZSeBYTn2kUZka8Czczp3at0HYBDru
VisVPk3/a/mHYdEXn52qWuLugeBcCqEdcQ/TmvNOiMB+khHfNDuUQXSoWhuB
3eTABn8Kq11WctgQb1DQGRI0LLorO26QSk5qHh2rEfzVxjQf6oSMfOheLNSj
1YCMz93V9fkhbRk7zo9iNOKfTSy3bNFHwrEPAYV8TaX8nFqpcsEfOuId/8Bz
wIf/ebMWaDgNA+AhAo8tyITkZoeztEnbq0QqaFhaXgHYSRiUiAUBOT7Puv70
zfDKRavwuWCt37HiVdHKhMuxkULs9932tZ67VsfI/8z+ucXyhJ78cFs10bEN
QuBcpCQIqUUp+gjmg6AR+By911LWHZHfppWy6TTJRIdb96bqqsrybqZaihPP
FCdKnaCAhHUDS6eKKQWlb/N5ucPTK61DVWw3ftOlVTVlO9subhrD1+F81HT3
FVNVkfquR2Jxypo21ixX5eNRLoxbzf7e0mUIyFI1SK+mVN0AwzH7fkA7Re6J
qyIX7rdQX5pQ+D+/sklm4ng3mskqd49Qru2MTuBdihuBA2dK/rsufhAn+rNi
4wDvmW9QhtXPe9h8fK8mlREboFrvrtHBu231MIBZgjSfeoHirZz7nQtblo6N
Ug/SpoI9zY0CTxprkHYO+MAH05tlrBrrTsoz9ChSIS90xnRgZjbgOpgL5XiN
KmxsMrQ82NgNaJ5Iwze08rnu3bmb+k2zivFJ0Pf0OOivv4ADa+wxtdhyrtNW
2NCcseHBqdsAUvjnlRaYJd6XB4hWW7CMPt9W/IJ6NvfQCHb/EyQGJbn1JxKR
2job4ovcWhlLLdX27bqv341OglY7GNogE+Sb7hcUklsjYjsKtBdlF585Hjer
o7MyGWDjMlfw6ylBY2IWmQ76bNLeD6RyR0LWgQVfxGQ8iE2yAXi+9/HeZ0Y4
Hw+cEWh2jHpIuL7kF9CL5y/2shQ/3xjw0uTsHwRyjSaVjRIaFjItjLzWfTcn
2J4KxQoLkmHXE/QVslz95a6dz8QbPfd5Sgm37GRCErDuroSe9cwwSzsToGqL
R1taOvQQzcDEyCDyD7SPi2w36xLIJwM3R48Z9dpH7Iw2OilDZx1UXjoU66K0
Jg+EQZZvVLgikJY614iXsFp1VdERMVfOY8lB2xOOibR8whnqGlDM2uQVDT8i
Q5T8s3+3PWonQWYJ444BlsCzVssv0OAAX5H7Ly4xj8HiLHL/+LvEqlMJGkEH
pBm79VlEZy3Br7LLEg5v6dsOUu2NZrqtd6hyJ/pdFQfRDd73wSr5o4xHg2t7
imTmzpw3jO/6gZcA9r+HNqgJJZ1Q8F3yx6zgEHGH0WtRn31NRy2wJOU/daCp
sLQ0MsV3JyDCzdNqafd79c0LEivNJFeZ9J19F21R/yyV8yN1wbFFnLeh0McR
eqNjGM29NpzU8KX0cpodKwQPZJPP+9xMKEJuA4YTLVUj6RX5zv6cFTYeThxq
JW+3tJ7kux7lwnBlvhefOzG8MBDYvVsVsolPCPcWj3SnjYirxjcwxjXxaeZ5
dW5q6KervXqVkgBluA5WbR81WtNSKE16JKAbno89s8E6DVOQCIfL5uNhEZCL
rTILAn3PO5sIOOfZjtSYYm+u2GsND07DufvxUby9ey7i4ED4kLdx8A+IZL8c
Kujn1F1T1/K3uDBwWB731ZesryYwjHxL1JEmSVcE/O/9DZVJhPxrpNrLCdR1
SMjawQN1Dnft3+WXghPGSuu525ci2q6ckGloLtnAfVvCKE5u+EdcDeqL5vUf
ldDq6uJJ9CcXA8dHlImWEbwQq7PP2Lz0VykmCetNKbhtVa9y3f/FgcDYBxWS
N7TDUcz7GBWAYYhoHj1Ntu521mjerg54LcAbtVNzuFYrF8DBjpEl+MDNLxO1
eevwAJfLYKg1e20mX9fwsWkIxoK1B5DwvxqB/0QzKa2qVe+OE/jpkh3Pt3Pk
YAy8ztF+jLwDYoQ+xcyS3BCVESRe5YLJATeNpY8AFEVv1x90EQl3koTvZzKP
BVF7hFsTB9zqoZJXBdt05IvnLrPl42wb0ZX8z3Mom+IMqz/sRpI/S6yaxIJ7
c8HyipIsvanY0Qf+Sw6+TRtbx8mWi8AUX05si8WUGT2aoOAu6YgWoHg90hge
NU8KV4xj35J+SLBhE6+lFb54g7DCh4I1HacV8yNxxW7Ltwe//OBOzFYlufrf
ZDI7CWNtUqP9CYt5Zzqz3Ph41/lcoccPV5fIxh6If31NRe3O/Y9TS6hLytRR
EDHJmJbq/OfUmAyLAXyU0qhADnZ9Na6tu3andOFrehXebhW0RFWbEIKLyVPj
PcRUqR/z8I5xbxwE4A1rEKa3NA9YJP0ydwTLHxPwPb86c/QaWcFXwzs7MeeP
yqjVTV9b0nSVWAMrYZGMPVdcw2g0S8yksRE+gv3f5L9cWpkNP2o02z6Z2GwU
dlD07n5mKlrFUXHQXr9WjpviLdGEGwxulX7wf1CWFHFd65tbNsmeyEQmBcv3
n3foqpPUZrCxwwVBsfSsDxDqlRdbfrsUPh1L0iA1HpzrUuHtUvSf6yz9b/md
CaCMNv7tDKhWAW5WmaQETdESaRVUI0TJ8mDsx0ZIDdwiGV1TuEtWu77iwbEZ
idfRaW5Flk0a7wuA6nQ1pkn0wRpgUw/B+q8hhBcsXtacdhvK5UIh/HyeeYpv
LxBQxO8BD/+RMjjpB30u7EvTrTF3ZSwhDVUuf3xI49ytjOJVAjf/u5/tRd2M
LKq3BoFhva+0HqGgk7ULeD9U24kz/jKLYK3iFBlCbdP4PRQI+nehEckCoM+9
7IyafRgemffvLfk44+vZxB2husA9QYxDxobg2thaG4Y9J1HCUaf2JQ+kkzHR
lCpv5AAHqfGdJU35glO/3JDsnBT0n3heSee3MMWgbn9YkiHcga8doXegQUAH
j+cGP4C1Yhyz2DhMExtgrPYXSSfQ8GgjedaFiub8k/k/vBEmoDe9U/xa98GW
Y5EuLAcIKAanMcSE6TyDFckXHCu28A/sErpteZNylxmyaX+JgapZOG300GHx
VZLUmRhPiT2z6cCK1+mvfJjLta+SGKiCcLEzg5St5d6GF+Fq41tNGNVUCLLS
V0lFEv0925pylaMAL5U9G1Dxo/Neq6gXXbDDOHn/J9gMNo2E0jTmr9ci57qe
9QM+3v5Lk9xW/iXl94vZAb0GxnIVTkZSCFy5MyzNFCL0VGJNRyjGxnBHnLKX
cmaRy1XSCPg0xnDN1yuuogVx3/88c3obcViIKtJVaxUfJBXCuAdbvvFbEIcC
iGHSJLAitNVPrkM7EBAtGc9rDLUkOidLyLDA9YwUkoSSyDB4PbY6itmUFpzG
VyAK9L6Pknp4A1F5n67T3s600ysEmgoWwLlFM/+aiMKU+OwZJ6umjCg5QbZk
GDTqmQaPMUSYznsefqadTLtP4gTCV6kwSmGDFhRuMCewN0z+/wCu05myL4wv
++5IOf9i9Z2IjnX4T3VR67wt84d9wPkzhrwxKLzuVIKJEz1omPHAtQcw3SOS
GBlblrhn8bP+44EgzuY2lBXDzZdBsj8WLDsG55iIaaszVLsrZYjIzRGAUMcs
HP8IJokl4mpZhHNAvt9A8WI1A+LbC58FzaYEQFo13xFMEW9UBXI7jEXXANVX
rKzeRVeq9fmjNi/94U4W7cJDyPsPU/k24IC7irQAOcteBj3EWxrQ0eBwKnlO
pV6fhZEBXutC+pzTf16VIpPNaIlJKmoz7N6vRx8pzzLWkNzxwqd7yqWZmsDB
yIaX6gKPUH3pzI4p/qDyACcFHlp3wzfcp0wCmUGVEMyf9mLJutLtpsxwQjWW
b8DiZNZQ6ZNgh48wFKp21wXKHmLVBkBWF/o33D2BWyYUn/4mdW+rNw/jxZXR
s9zI7on3JdPVg1skE25T164awONb0xvau+Cq4+Bd9rdEta+shsXzxOsbF/oy
XSYSPXJZ/1BzmnPiFxKZ0h9pl8aTpgKuHmNfNd+4sMWCzz/UTdAlpAGN8e5Z
xTcDrpuhtT/FY7a2oiU4B4yebkDVXvu79S7H0OJHeF4/m2oDYxjWGnhuhyw/
DrIuIHYiq5PMbFh9AXlx2TBQlp2Ri3XuMa8Y08ZHuVQcyDLVXzLjWH9GcL0L
CT9QWd1EM446/Jh5v44b3J4oTS2/wKeUc1Xath0pSY7BuqtgsjMylWL5XHgq
o1Yc3XFuIfVjDw4F6+aXMIZwHfJTsfv8++HLwDbQ2ePnZ7sJmHkNJ4NldeMU
URJfHwMchwigkDgok4yg2/5hIyzhbSUxAHRcmJXbKWYANvfElrOVv53so09u
EkqqAWoaMJyN5icsjp5KmWfuAkg+lPcRytMH889q08gNIDlDYldjrMbUqVhB
SPErMLXGmySKpsVKGyjrHGGYVsfJr4baFT6CBPgs6dHeAF8waPjIJA1jBXfR
d2d+djtY7Lz8yuwdLnkTk5Wvgsm2PBwY7mUXx0NIUsQuxT4jy0hxwMyW+VYp
SD1SFDHW8EJ8Jfv/Bn3QGMMGpOYbBwczwsEqYgx1frKF++yc4Ajfq7Q8PmYm
omTxGnVEVUuBwnWNOXCJzEal+NBrCT1pexkWBfFQ6l+SffnffwcimvSFvEyF
2QEj6YPAJAwRp2OT2SL32H/0+Uz3OHT9qlzcUybPpZw8PE8KnfceShSNg6rd
1gDCch/siVztqDtdD6jF3spr68aikpP6pKPSdv3JsH4FejfiBG0xtUAs72lw
/C4hrsIwnJ7oTN4vG7k2oWisq39ipUmjEvMJB/NBUojFk4XqFZo9dxJoWf/9
HK5wKR04Rb3SAplYmpOGJPlUqoL0Oj+9MNCB4wBYUZK+W6UEJF0IAJHX7Jc4
eCU1nGySeHQ8BF/0W4wJX2wvdO97zI8K1HUm3JtGrz66sYkGvf0hIIko5obk
cEzxyPn3K+2m/Mr8yz6o4DgGY9gTyrr6XV/JQOQKHvDzZEmFHmPOstaY/SnU
G5mdoOFL5eVQNl7V3num+2uwp9LW5qdogDcGrO47I96vfVErauTGuYsFNQHu
8tUj6fZpbfK9/VkgXVC/aXKUt3OjyQ1B+F/NW6+oz3CRgDaSSnJ3+DXwc1q9
VDgqargHltTvW1148UDjxIWbBQu4ndgtWsPUfugYn9Tuzn8nCcXkHe44rLOR
MNSFmUe3Vu1nbAMCZ5mGLRHdZi808JDJez/Xmj7jxGK2CUGqP/O4I9pdce8J
FyQifugcFhzwrxLcvpxSryJLstydEPrLYZ4Gl6TT1kpsK9JXUHMZD+pbSYdW
quunoZ9r1RgnU98C5/350cMmfLhAzTMK2kzv99K1+LuGSa24ukG97rlZn9ot
wJiKDCeXginTdDpfh+ytTaAKDkUqzlLkEMLiG5qTndSAzbjPGRg1fNLDqTPp
iAGisMsjYg+XSIopPKpEJQBvzp2GEwDrJZICiALVc2WHN/mzhZLX3waD3i/J
D+fVFN15gO4VSk47HWkH90pJAgDTOb9HAAJMap7I/iq0XfwciKrwEPHvZ5G0
s4QD4JdXJpI5rvFNgvMEiAcM3dM7COqLgMusVAVhe8F4WuDxW13gwAh2UBZZ
QjWLibhclQdLmbt8ob+9JwW+s+vfOQ/j2iiAIjuJgdAIJ5moNWITbFBwdbA1
PGTRe4pKkB8vfZ5aunRtoHKllxB9Fmbvd0AGhfhEnZ4C9S6upQBrQYi1kCf3
uijP3Xh2GpQPWbGQ5LXnW0a6gTo45SOpdKEpV/2PYM/b6JKiudsXCVZyEeJd
wXcxoCidKfNzKL3SSHImBr9YHNnxp/1heRFHgnFA4dxWSUZwo/5PbZBgB3I8
I+SpONAluddy/xfpZc8gkjTPzCIqsqEOqwVl/ufEsGB2xtZGasxB5FKnAJIx
QU9H3TpwDfbaSDlCe17bUYFEL+1+0Ue7elnSSddhfZv5314nQ09iuOq9EYbz
jphawvcn67fI+QdBT1eDRgsF87FgECLUs0aVlgSDrmk+TgAhyLyL9PXp8kdG
PNgB8soeyw9arIBAybqCiqQINzW2OhEA6nVCitWZ63FBWkoYIqVGKAdQbE4W
0s8RFnaal+w/W9fA9GNKY4N6FVWAhJ3cuWuxHWtCoaa3/BfuojfABT9qnTZP
4aGyyTsYfYW/0U6Arnv3wcvxZTtThO1+SFMjL2wlJ6Ghkgn1WNHU8m6Q/aF+
iiSEI2gWhKVuSFhsOkw41jzbdCFMtDQiW1q7CFuSSEFtxlip+FGVk0YpgD4D
OyWXyd44mVWZ87Caql93VjRkOa71kbg93MDvBxIMf8G9pfPFJoEUqbQb92tB
Z2YqcelKvKCfpDj/lxaffu8eyDawq7E/K1afkILIwNmS2Q6KKTR55fhnWb5E
mBkyxRkk2ut++3REvzybrLyCp1aHgm4Fi8nMExWaaN4NsdxZzIiqrfGCPVLh
MZxOjUuqqP6iyVuNv86LjH+p8LYwo2S7miMvNYtIroSl3xhkCY2iUl+SB4eG
81laUvvdG2oq9WK7HG40+MJbJnbWORh7fkWQhLwKURd30VC/eFD3oygaDPMs
DUdksMECkowMgCIkbYdGRu51XUrrUQMWWcrk9zWL1LMOKzcEPPj99u1yFsli
SEow4syVehJzoRv/NjzfDGhkWjypIuS7FvltKkmULtVw2PGgaEYiT7tNarGX
zCI6zfcxmOgcQunfL30MNVQlnfr8pPp+CxV7duBwDBGOrv45kc5+sJsT0YTH
I1Y6RISos4SX70m8nE3dEJxS8voIXGOo2V0tcd4+ddCkOoCVGC4fNjo2xbIH
LsLO1/9eHTfBmysD8RH29BAGimYsOdLYFX6stPLR9DhDxTx1lr8CjyAUMolX
t2Rvkea7RSrUJnLAo6Sg9XBSOcoojeYm0KAZMzl1QA0er5rzbnkRyaoW8Z7O
WiCyi0n2p54KsHdLsyK0wqUZCvjaslYFD3IvJxoCuNNTUxA8GrYbJ5Gz7oen
+4dzT8KuSbUZf/zlwZWVmz7tJ9uqBKefv3M0iZnZwEgCEUqLtFMedc8673/0
AC3ZZIe5hvv2ugRpPWwKBvSIq7a1RA12A0+2v01s6aQ51jqeVLqxfMk6wJUE
OAesX4QzRhrPTQDOMESRvYRtgN30ZzvgzbnVD7LVHRpWJijHzEYGHIvx6b9A
rrnCyXi+k4ksfxt1S+iWTGOcIbTZjoh+1ci9upNtGw0Dwx/wO4AE0PwrYcQ+
9t+TQpCzmRDOMYM2Ivvj5j10/BrdShW7IHI4C4K/v7EhXOzatW+FdSla01i5
otTQhbv2W74VXMBBVl3eewVQ1pREbWzKVJDZcllniEtlud391w9O3AWoyV38
7UtrNbt8taSMZaW3+LSGPFeYdCuzxwGf+apYEBXd4UEl01N/7rRCbdPMYhAa
U241xCq+DfF/dO0atyZPy/PcAJOSRpSLRDKi+YuyxVdQgQNzl/cZlylEOITt
uDEg8oADyzfHGA62KwWHWjms7WicEfnmKj7kv6b3eB8XWNc0493CRmPPIrRE
s4BVuUUa5HLxmmhXC6JoS2dDGKh7vzvFVSpgndf//Vpyl7v9trE6YftHzzSM
AB51utnjN9SkmQ/GjXbAD1/N8xAOePjYpO0RsQWt+QbLctYXtSnlKr78jyK+
4GYqC53uxtT2iYFt4/8idzO2PEJKV29EScSa2eVPUBmuj6uzZNh9FmdDjlyL
5htiOyiBI9iUOTUnZ+AlEEAgw68T425bkhUiErNUi1UqozkFq1jmmXiwAG6S
FzgitEBm6sNtn8QOKwfOjaCylCJ/tQZ3bOux1SWJ5PliM6x3L19syYS843ja
gloZqGHs6jrxvFy16mjLWb+uGTh4ZLesjxMhlJw3qjDgbQHLJt5/BOWyefkn
tp79B2BKgn9BxdNAbTgGQu4W+JfLB7Qe0Prev0oIgbPvskOikVRWTx3mG776
3wSmkbkQXt9RU1ZvMQw7HnYQo7Z0GTa5cJ06ucJ2yYxh/lW29OC9YUkXxsCQ
eMhVhibGBAVj+k5BiPlkgpG3cqcE5gvhmMpZSw1ylOQTNGajf4R/OzhX5G/l
PzeTcdXlB2r3tblstssksrs0qKGZB7YhB4YY2Jsjm1oIWOjG13HHna7DqCJa
kbO8dNqt8IqkBib76DRa7iF/Ca6OJ5xvwY64ZaDOU9Is8H4Ny5JOQpseZE6O
6todgbfIMy/z+Y2Vo+Mw12lYUcEAzfA3U5Z4zNHXCZDTH3hAxRalPGWhUODh
teYMmIHAdhwZP8Qq6F6C9HFNiWxagaflZk8ooTd+LSqSelFw4PFMzbMPHjWb
k0H+F3BNhgQCee4Min1fAdb/fUnd6gMhKS7RE2ETPV3n4Bt3VlEsW5oJEB6f
EyjaMb/pnN1xEL5wzMK7O55QBour5AZx1ZB5diVZ630BDJbT3xT1dCTeKuYD
0JK24hoQnlvPzJHDTWX+RF2IT+bCPNWqOU2tWA/mCBXo4scQXPpOEJ1sR06K
e8X1rb7dinq5ZgnAPLRUiJtFYRkZ66c2SFvxTIP5Dp3q2fvXEFojfa4cxzyb
cGSIjufhTWH4Z2r+D1zYPV7V0LvmSXRvF+kaPgehjKI5o+M2o4HAx30LrjGF
FKeGcPTkfjvVqEENqiDvvNOOC9UEIOgQiFIE80oT2s0RB+7i6x9RyqAUk4UN
O/EoBSTueZkGT37gxXLFrXcyS6IuFLbjX/L9xr8MfGQsgUgD4DIgemvVDUQa
W/ZSEjjs5IUDufnt8Lf06UPK2oKA2wQaM83YHsNviPgdHfZbxpbrXFo6CiGa
1Q1am13uEdKY/fTIvhl8LnkmEd+OaxhUgjsiOirZ5+vuYd1a5Paj1NsQXU7n
r4snS9zTiQ+ASMoOdLm9c9ODZ6275MZ3aFb4/xhdyFhTLw3pL49zIRmylPfB
FO0gQuG0aa4u8F0wksxq0WpAiOU6wML//kvzS8/Gr7MDNjwAs/Bi41yeZixX
XW1NN7DpjmjkxfgzgUuL+m57klozp+EvNQLOtyHBH9bEzI8q9G61cCtw8Sgw
zQ5fZXlYTfbuhU7vzQ2/NN+mR5xpaFZzUtQBYZKP3oeZkGWvgzvqaMYsGpRZ
FmsWqa6mH/u/7wq7ix7ohQBFqc90dcvxykvQHG8Qu3UvaEqdY9KsrnXC1wzJ
xnrpzX9isTa8JkZ677czrVYt+pXj53NxMVqgqpL8haoqb0ty+m3uBOePJGQH
fnpgOJJ6DzKvOq/rcUPR4yDJJ/Xir8iy0Zw3gKcmKE212XPOqRGxWvFzyL94
bMVGJTEJXKiDu/gmBNOVOXlXjBfeeQiLXYw0Bz060hrP46I0LCG6YyVtW+eR
zycxqgQhFVe2OYsIcuWzeStC+0JuWtEgbY7GxtZjorauIK6ziuDnzYmm+JcO
DHy0r5MiPTnPe1xID3cvIpjMK4jaj9HUXyy6SD16X1PJotfQH77vRn0WExRA
hcyopPeEgh1VmZPxu0SOp8jvw2TRM1poVqTwdpH0bhS3dRjDvn2JdyZBAY4T
7SV2t+w1+F4dtpN8kDCaYEeewsFOC9ta5ypFDSS1ui8sPsnfiwNr6CbCTGN3
xqSBYf8Tbbr346JP3Eq82zmgWz2Zt0QoXHFsTQLtRKTpjFsrYAnisH8JIaAd
+0khXk3eResVZgwasWAxOOn92QeS4uIje9gPSiZGTALNkSuQRJlDHs4PEI45
d8vtrj26dVY8J7lZ2b8xF920U7Q5uvuWAw0lTZEkBPC7/7zNlgkEDis8iDwJ
NAvqurWlHhvLCBChjHR5kcJ4JVKVJBk5UX6XF/KX1vEMap+RT1/zIf+ZMVDP
oiOsQZkbeCRmiNT6/Nf2xDKYB1akG4g6+DOakiiZBikucUC64W3fcZRV3tpH
PGi5APG2OnD25BNMbFdE/BlGFXsX/aeQ3s0o+pYmEp/z6sV7zFdC8GQPlTRx
jq7RSFQlgmT0+VivS6aA/LZErkZuZQhp+BJ+c38kETRqglOdW9ZvFnlASxXJ
q8qhsrY1+bqFkZhkUqbdyC87ifDKGuNFenegPQ/d4ReUGyaAczappGgHpqwG
ggDhQrvAFE3MO/HOpADIFM6MrR4hOYNzFVsXxkrOYQ6bFOPHhm4yfWpV7LXs
GoI4j52Ot5DnseHJ8+eg7Pwx5OzS1xOXXhzMlF8bcBqy4BroouXqWEGSQBHW
dM3ZbnVm2zty058JJMOnOIVonfJ+/WtJ46y56xaR4LtP26ODQia5CVAhePem
4uGJ6Sps5ev4U+ePHPsEyFKgOuT4IOsz+EDG2lmsMNFST0EXACCu+7TN7cJi
cddVBJStOtQzp2QSYshgNb6l4cuKJPLRW85mOLkre79DBZk23Nud6hrQqDqw
Qq0cSFUb2ljIfpgn/M7lWFDXCWQja6BgnEfpJMXXqYzrB8bWl0VzBfT6uFwy
qNEFtIXCQYpfhpLWwyqIXS5V023QBycj+ieZorUMNVcrQ5Dyz1sXtlGaRIJF
0Nyh6isuj9QsZIgLu+/I2shpmoG7cgA1tkvAFtWlXoxdY50/6g/WRowJ6Du6
ChX/ywwkm/UwBcaevrE5MLx/gh1znw5xq6sI2E9jgwlcCz1Raoy9ZMydJvtt
pMz8mi9c150EO1GD+i3esyNg/t9iaao892juQZ5qXZqAfe/TlEbOHoedn6w+
1CyDzEUZYa+MBsBQS8Vprl6Wq0RdxzgW0Eac34EiYKiG+/8SdsSwUmsoDj+m
dqAmjUtqb8T67Vbs1CAT+QaeY3DhmP0W8G1z+w6chj8bgh710HAs/Zft00L0
kbak8nIo1Zi8ACJO5D8mByY6P1pHcemlitaSKF6W7qbN8zesyaLJg3KoyGP0
fhK/VkagzQ5JqkDdUZJtJzxzboqQ1lBNsyiSe5aOCZ+5iKpyDGcvxGOM90cc
H6qgvp/8EQVcYfyPmrTDyYRf9fIWNBMR0dFxuBMwqziXNdbTAXEWlH9M98+E
i130YYMtm+fh/ezLC0ApUeRhYHE5AQcyzthnhhp2D8yEigCH+165GQdKW+4m
Byhw3KprFFQkvZNA6snGOKdcueeac4+uB4VSHjgdYOR8/9JuILJxlYU6tlq1
52Apc+W0iTGEYw6t9evZQUMYzt4k8uTMl+Sj0JUquoBiGEXTbJRPjjoipehw
o1kOBBnrJrGJV3Eh5i8skIanHYdETnOcogifPy16W6agwyL497kLZw7nMzqV
ykrmiPrMuHwvkyesaOdzVvK75SPfGAdMZYIL1OMge2zKZhbLQyp0ir0f6FLC
9vIArm4pNBHcp4Re9aJqUBo7Y3i/Ylf594n+eyvbueAJuN/dv1Az60Mr/EVK
Zls49S+eiaFJWnGd4gg04eUGT21GuYSdGbqaxLDW28hOfzsF05GhmpEzbJB+
ebcSbqdXEc7Ra0pZbi+8at/LaGw4hivPsXuv5TGIrdQwuBD7hzEfIwheHh7G
wvwEyt9MEiaOHAeamL+TWkWneDsNTK188NWJ0Sixoo3LGzc5ihjb3v9DuuVo
dvBmEKhgvDHwcETbKyj+D0WTr1LyXUTl3/zQKxO5NucUl8zx7FlyfOJnnv88
8Mb3c6kRbyWi7Kchh/Wt9QL5MIsbfovNIQU41OeNz9xNSme6MJxOoT9Sw8cv
vB/nQBnlfX47vE3EaQt5kYTrZ3AYxpV7jbm1CFlaWCposBt/VD2d8JgamrEq
1839obPZtnM8O0TVdnfdN6r0aU/Y8g699ChicRQvkU4maFTO3d79g18AsJZA
UCPLzPyEIOjGKG7bn2LA7oN/J4GdhtlO8dB28nrNNmG6sBcXYCcvYIGaErzz
we+zCJMQ3u8EI/7qGbasaNreP2ENEjwNAY7HNjIKJHYyw1VniPjYiv03Edne
tkxvEPDd/msnvfxtz9Lo+q9iVlaj4sFgbjdeygZLGyMv8nHBNy48Y69jw/F6
/M2nMgRjRTAtO7QLRdAwbrrSkR1W2ryZsnzWGAiRwHXRJV0n7KN88bV5/ufv
kcRC/rq8FSWkhEPoyAMNGwU5NYlKQ+a4O9KKJwbYb2CDFxMNCP22bG7SMtE3
7j1dwcbyXaT+Ha4CYymhe3Yf8+3Hx0fSfPiQLug0BT3klOIh4QhDD2KSN26+
caQJm9BO4qt1q1B9w5QqOSO18o50PH8KRIyK9Tdipb+Y2XOfYjMamb4ajoym
usfrPmJxHCtd6xP7d8apVEVMwk1bpL3G4JeqYDrw1TbH2VvGaEqIqySYkwXk
CYuQFsvq284+L+uUgqvWKZPrqMgNfeCY4xoieraDAY1T+ii8CowOBc5U1KRq
CwMicfH/iTHFTdy/h//hBOoePjCAUTZtPXJws5Lxru7tnjZVqOPwDPwYWgw+
Acs8dlVsCV0Brg39u5KLnGI9HIJ2tmSzHnBeW6XtnOh129CDi+1cKnt4Ppzr
Phy7P1EUq/oSfU1T6RSVi6ke578xpwHb+C9OMeRtfB0G+1saz89N3v3Fb9UD
TOJXgsVKjOBWgURiVAgZWFmX1ndiPM8Bd7V73t9EoSAbtRPOdyn2z8gI0fmE
qLFXy8QSQsXIghTW3rDplRClz5enBcLWnWFQ7lCK8N24NAL/hjFgDKgPXZ+J
4wY6zl7FbMcXp+MyrUritp89jDVTbum5a4Y7IssJScL/iPk5CdjXlTozNZda
BW0rEpfd5sMSXEvaHYyLMIK+qMrJ+ARtj0truzQll9EW8csHURFKAcdrgmqQ
qGfpqlb3oGj5gS1SAmyXLKSELNVIACnw5lnB51ZuONGAoPCBxuc3YID26L1A
w+TvU7DFGwv6OqCaODJYF8gl2OxwrDPxJzE2zt68bdrc0HgDZQgEw3xRV4nN
IsAsrfsm8RgtA2pz9chc8DjeD6LWmJ7zzAluSVu97IMqWF2dIWG/rRzpG2IY
SeBCz8XwecyxGxodaK91CpNdKvRqhqj49oBeAygyq4h8eXZBkZiQ5oHU6Fcq
mYzDeavnVU0E/ENQrOmuTjSkSiBh/7jCCy0aJdVeJEs7OPBiCHdV+Iu3c27+
TNjve6Z0IzGwkorRjqsYnQH0qAwW/qc+QfbA0zut80lYT0Ru3jPtOLl+mG8H
94krR2LkmPIQKXGL3PPi15awiOrDWNzIpxPaJHCkHkJWTDo6OBrjA2GS70UR
pox5o5N1F/7vwfUoi8yXFGagwqHLBk+hFsQ0AqHH1MLeAP5TQdOAyjOz9cCT
RU33qfepMz/FS8j0isi7u/aIOnlcSJ47hPIoYImmZxEv96Pqpn0crv0I2MDD
daJgxj30VuOro2rofgCM7kQFRDBbnYZGWXEDw8jz5OEEEsXGVbC8J/iZG9M9
hyeWncuFjUk0G/lnrsgoHc4LjaTq4aIT2+JKi16YsdD3t5tpBY5goZMAXybR
SnGr2etaib/iYCdC99ZY5tCCbSXKJ2TSKVZcpgxk1WOmJAmL3zpsbmwgJXjk
IaXBABCk3/fuZpi9v6g4wTVJSajH6P0VEYHCUShHmnB6bVadjsroPiLoyytb
6kYgivLb/CVb++K6ibhAxrCPPMswd37OiegnOWdlMAHskkmN83/kO9tFBl7g
mvVr2lxkuP0NC0ezQQ+slkghcf2SF42lc7GoKFCLGWSGToBvU/blWPb7euEQ
eMlMd2sWVIgtbXqBtRnD1iIjgpRomdIN10gKQ8dKD1X4ZxRo5IQ4iKlv6Eqd
icehNHi1zX3QH7jXbEgP/eqLwZomyGtEPerZMgO3kqTRdo0yUigSxQORitvK
ZhImXZoYsEybDkMmIuPA+edyfSM8grE2qFAzRqnu14Vf2WhEIVOnjEfqk4q+
jo64i57iiccUjqtnPB446WpvEvH3MdyUxE2aKVjptc7cUfQItjKc9lOPFruu
1s7HCep1K8DKKAg/r6MFx83AYY+N5OboWrLvwBc2C5CARuzYFj7GMf8SWFfj
RbvDjf2QKtVjUpiJ3XI/dT3YgM8YbaiRvG76fnKrQGvclqaqHONMlbbZuB1O
OquFmu/SNNhLxENeVGnEWqh9TVh7c+Nmlco5tnvU9D28CnTBQftsKn/NIr+P
qpXxUxpTXLai0NBwzGKwbwD0I4Q0uAk8Ncg+kbi6MnJ6CrsqNDcAPyb9J7F3
sUyK7s+k5E5fKhdolw8eYJK42vCmCePb4iEcyBMAHobK3Kv9OaXwdeu5bEMm
yvIij+V2w7G7RfZMrCbR2wsiy91hpqzcaH1U7y0dMFUtEJ88PBjNacNYN4qc
tx5FEhiFLFZNoRjnMRhlC7gIXYnvq308M8DGRuojo+TQN+v1ehyxM8kDbiSg
CiYu0LqpTTslqS+TD6XZKSHH4nE1JlYla4DZqMGxvFrIjY+W3PoeRFvjpc7N
4T5AznHRxZCCqi2OrHW4L6ccud4hMuOd8HVF1Z2qGu3/EztXQX2KxWsOGReG
5WGPZO2smIJ47QTtdH2YNDW8vFvJ6Vv2Onhb/VOSbt/2/lur3EUMnDDvC2PW
nxhXaxTnWeJCc4TeYacAM8Bm9fdxIxI5DG7mXSzYdQJJVt1mXEpqgiDFiplH
5ITK3uul/i+wd3F8f8J9MRCH0S+gU/XcpDX3LYVFSzC0X7puPf8aYXvMbSSj
oFw4s5cuUVxAvLotLf2VUbZ+/Psuam+on2LpbJ2tWLzdOw7reD9HA20cN9xL
ykliC22fygs3AbV5YYLKHyKIxj0A37s4Z1ahvDXJZS/4MuoqPeRMvk095b4f
Hv9WPGprXq7piyG6wd+mpw+vcK28OdMXBD0qUoczskfM3zwQ+0kUNienv9H1
wJOUq9q9SZWEtxWX32r+hWEAtmq0FN089KOma5Yqzct/JiFb/39ujLz5FD/Z
c+emHH0BtimDX+Hg+8VJ56hweNeqCF4NnrIypldo6BLYByje6Jda4tO7LJMr
5F+vsNz0a53rR+o6/VOSNe6/zaQF5gwiKyatPbxzOFfjSZDu55wYt2qlMNA5
+KJVjJ65T4BUrJcaCodKRaB5EvfhVQYTJd4zxFhJzER35dKO1q8GJ/ZhmZzb
cXGp9yN/cMCc1i2eGKxrrcsKCVf34KacMH1zphVp+mjJ9JH4YbXQ5Y07r/A2
VJGWRuoTWxqSupFhFnsWnae/imylx/z18C8wnc5sfrRqzUp4HdpYDXoFvq67
CtAYwBHsOOkm/HXQa8oiBUFNVpXipMzUHpzFkzuEv6sD0U4IiQ8dSC1w699O
plugitTjAZeQHDvvJC4OKWs7vh5yV0+eHz8YOTL4QeLGZQW05UXG4np4Wj+m
ld6G6Al3RnR4nHs0/JpxEjD3+RUoL4FYClVo7jV3R+BlY8ZGnlXqmx90NaBv
z772yKcaB7/R8dXHseo8WHLMYRcL33iwXflpJjm2LgvmlrCKHRXSPRiglQft
zaspBDyZq3Mj0LPPlaxaAzbf2o7A5wJOp/4cer3i7merFxPsJOfWCHPEAy2P
L7FEvSAlCBk3DvrdJJdadMN2Qhao+4GJRWyEwd55qf0Mm4Xjmy+DmMnpHCr5
8Cz/tnXKKInsHRzak+hXL2VmitwxrAPXLbrAMZCBefZ3aD4QSAXZ2W3Vym+l
Dz2pg4lhd+Ks+1V/wizeUW3//ebj4dW8eJgsPuk1YbtKvVU0wfKSL4tyLT3I
rua/zPVfsARbby0hsCWkhyL++FPYzKlE6Z4TH2V9qDXBIQyd5sjtW9vsGAvv
krnkP+aJSwhxEzk/I1rHxKtRK+V6TIyjIE8cCS80Y+tEaKxge/pw0Gf9VMy2
TWIb4oUKEpzaFv7NX8TfYHBFNCmFnb8uZI9jF40mR+PoDa9QjujG73qEEif8
VaikdWsjsRgk95sMolWeB4qeK/JP0ZnNi8GtK1AUhXJmqwF5id694Cgy657b
EWiTR1MZzU1IgdrnY8F1P0Lxt01gEORMBeGNkB/TKPk2V+hOF+Zw50tyk8oy
dl7TXAudyv+CTnXjc0GQ+M+zo41S3tnoqq9qCK8+4jT07t/1sDg0gOk9fWbN
jegGVRLgaXFaLXBubqqROx0GkIy5HvOqGcoIRSiUASo3/RpxAzLGrgofQD4j
yY9ufYD78MSWY7nOI/q5P9mpwUC4ivY6+LN6Q2aiMVa0+i/m2lQy93659fHq
nauYf1L0pF5Bk4wzqMcYrSaIZmW+27yqXKUEa4tZJDSp1OBwcC8NeLbJCg5Z
wqC8TXsB2tWZiAu/zJ1GqtMPMG1Qai5EkXuBaGC3T1yu+B2x65HlN2YWCfhL
dz0xm60f+7uuyVqnGtBH4tUyy1hx5hPR1FpnA5ogdMdBJcZcok7OjOomfKIZ
JwVRGOiMuZuTs1Wgsu2cXY8ONcLk/RSSm9c8EarkuazrZzR8pQyGmMuPdyEx
UtK50epPAiPRt/8vsPFoUhILOb2ehXyQbpWeSINe9omTVqs/MroJRPoKwgMV
dBwaDm2SFypVXLMCixKDrW1fdHYJIWtRa8ozKJGEXpHoq5i4yceegMUS9Y7U
fLPZ2mcWGKhNJloHgbOfm5YsO9kVTovo34pwY7OJOM7qZom+OLcrAVjPun0+
5Bdct8q3bSrofLr9z/Ys9TSIG6gvWwTLp7N2Xi9EgIVmDy/8syx8sglWcL9X
lSVSOmog+yJlO5xB1NQNdIk3j+gQwQZc9+1D4ZG9zjWQIfFXogIvhok4dV2o
ksQ2ZpNgM8pdT1k9CnDJ9QRrtJas/HOHOs7SgPstnPRNxwgFb7+ILWCc5wsM
vwS3igYPHXB8krW5+UbXyV2PM9HtHrzH+MTur2/haCxGXTwfO/lCooMqh0tM
wW/ancnE98qs0/DuC9dnQOr4I1ITsv2M1+MJG1+ZyX/P4ycF0hPp5JxMH1Di
5yxEoCVH95mzn636HUDxGObyIX46un6R8kSAf5y00h1waf98p0OzAlEU0jvJ
mnR94HBcEb346E2ck+eB5YjgoqIWv1Eur/RCJr4UjKGIdKyi2iMiNYX1wgMd
kE9H/PNAOUuXuj7d7NAVNErXh/A4kW18g7GseIvpVdmoKXOECFr6mIp2YWEQ
bteBdKUIKB1SGLlKgbsOJ96xTz47t7yQNEFKjFNQJw0QQT6LoqZjEk5WE1mh
jTrBTmvd0bYiDiz28IL86jbxwNiXiBIVWJi5JMP4XJFFtEwuPd+zYkzsnMzw
wfXxvXW7UJk2RAnmJhRQVFSUpWa3TVs5Ps+81U0kKmRtTY+02PdVr/u5Rbk+
oheaA9lCe6QBcdWGlm94GCDGJ4FKpXT0i8YStl55AZkMSlKS/hk4UF/oWCsz
Ylc/cWPs6erZ4deWWDQ3XvMBLpJYXUgsv397LYFNDNYu12jE5pC31+klo+He
SO68o+22Sjk7pGcWlIZ6BsugFBDupKb/gIQc6jnojv8MVETXfB9VvIlE7rNY
elh3nX+D78KqPpD3djBXcXiHj+UGd/QeZQJ6IC3pvljznkKEH165AnUpOUBB
bk45ZQVKA6pagw83wz702frR7r3hFlgiwmm/c2JXghVD51ekOEqi8hjvKn8q
WxtkCkiNRz5soyVsdd3qxoCkpBK1s/8YGcyW8YmF1C3qUphSju+g1faWTuuc
4EwDudiM8vr8AyPrg9vvKRqJ65Xbj5+qc/nn+29Do9ngbvuay67sEDyyj9Hj
OiOePif3WY8TWttMbLmapWLOJ3xOtvVYGPV87aSI6eVR1+X3bWO+ZQ0EfZHz
QjCd+aNGTQC5Gmn8mDR8sYjkj/oxC7rEPs7vhxyR6v2A4YRrNbl6cfbm33WD
lUvlDOVJ/yPSe/ObdsDxQFt69enAdircyMvnWrpyNs6iU2pyEawoJmDQ4zN1
WyZQn4JwPwf7ey+iJVd7txfqhEmbczKMfl4nk++v4+zQBrJjQcidL+ceTmqG
l+i0bgdoj84oAyrzRWewr6iapt9QYyD5g2Rhlsh0DNH23FUVfPeQTuotFfzR
Sqk41JkPU76GyazTPPMxg3KKEVo3VHl0K0C1YcY/k2fEkoTnBLinx/bZM5RD
njRw4im9niSJEB9chfA2F/k92KgnOAAvm3BSPaj7GARoLmTpuh0g6ptoN0uO
K51gNcOJyLLCqaZdbfXVk4Qq8L3qMTMJIqFFtSkgvNRa3RzsYufwVJe+9KcF
Dfu3RLEB6MeJ7KJFy3V+oxRWBMIBBah0wiztfEHBtnbTrrnEPVmwrQvb7ALn
NmB1SpnWC/vjywQa/9NbIMeqLvvu/h76dShHl5YZ9yE4WQv+KyDphOocD9PC
JLr9UmNCmqC+r0ithauyLzmqfzBIZ+CFONFOBIFlmQ5rca/dTBmT5qYs2iwV
HDUpGVmr1ohQCKWvP32HLuv+Fd9LXw0cXRQe4roKD/Cpds7Em/NzLH/wvZ58
m/9/x9jA1Rx4nm29105zNkNrDD8QwYYbHs78Bsefjzfz5llL5LFIHkt/84yB
ibJl+kbaeJrIbY1yFv/o6asnGUpHKd39ZhK4ElcTib59WpWfdtOGbv3diWRl
82w34aT3BFY1eV9sKw1ruVd/I29XC81Xt2Wo+lHUduAbF7jLsQu1exGhywXP
DtfMeDiZMosB+XUGJBHwnMp6A2bU/hKujrD7HzBAU+bD4eJI9YaZOO+Xnwli
EtspRizy2KPcWXCl51+lHr5FVSZjB3DyI8+lKEwq2o8wmGRNpPGw+4X5rUJr
8+T8ftgsHqhOKwibG8unWfoZsePplNlCSUzdiaxZ6Qkhnm4EDZN2awtm8CIO
+rObivctVu1eF1Ga6/7cxp3c6PcHEk0tTpnpJ/2RTusosWILANRBG9TsQJvd
Yyt88YU/59K8NE9sqaiUKZ0VqRArtRvO0Jtn4zeMo9UyI/Yf9yBovo3GYhqe
Cbqe0CDel7Yd5ioCKlWxJfhod8B3HyeS/1L0dDit2d0e4Q+rRHp+4oai+ptf
GAEiAJL5K4aj2zjuFJlYPkoCJkfo2PJvJYqny8jHs8ACzSkNa5eX7g0W+40Y
IiS8/0Cl4JHHbMy/RslKDIlPvVtiyVWfXpr7uba41lQO/iiBZSEGci72EnUj
f/DH2VlNN6Cjz/LlCdV9O5/11SpHStV1mc3NXTlVSEL/NL2tM5xRIL6Sd1RP
E3pbZnVpmMUsRpAgfYOWNup+2D7tD6WQPaehDy7GdpQSFA9qsP0VGNjRfeng
xr8riN6f6t3UqtoiKYfp/TZkPepQhJyq9FmJf0DTyraETmG3Frit0PjwnFYd
hog7M37HVG+bwsLrSNmQTDpObSsElyQOceEM6FGHYdTUDL/Bl93zGLE1nl7k
Qm9SN2N+iX0NIGJ4q4op4sNbDb1TBQ9WxjiGY+xxxWBrjgiKecNxfSAmc2pm
Rn6p1Ao3CnOA3rzr1lmxy10PA2SjNq9hFARH1I2mMgJJKe8n9b4Up78eRUcC
TG8kt1qXt10mHZfmNdnDg4rOLuJIsPnyOoNl7F+M3t96kU8aPjT3gUtPu81l
lP1y8kM1fM3o8CVvUj4COPJI/nJ0qJqF3LttWX9jq0IUgUXe2AC8k2DC/PwA
ped3naw3FyILuk7Nn7aKodnfaQZk0R6hS4V/4MnYZJ/2NYrjayflbEa4Rj8e
ccttXxPb1Zv8IQx9a29mvJOa0hfLtWIMeCXgmi3Fh7feobF8/R2e3xMYzqsr
7CSXHoa4VdLnZ19LqUg9Ag5MytyfUoSGwHqh5m2XmdT6/xsqPzMhugVBoPz3
QlfgbmrZPvMIJMVdnOZHfYZ8j34vW9WFy43VXl6uF+0i5uWlCk2X5LLcFJkk
n+l1N76P1gchyZ7lWxYXbhzHNNS3jF0/yQWk/Wtd8YSXR+/CeQMf9AYsBCOl
HEsIb3giuKSjiBaLxIvjh3Wot4wj8j6cjxLs6vyRMilOu93a0XJlFN4j2xkZ
swNHr9r3YBeJ4JscGh8Qzjss1/Ju6aPR2k60kYFIxvRH/9KpkU19iz95x54h
+iah2gPYnMr0HtnW5Oz8C/mJrZ/Sejp/Nqm0kQMP5RrZe55aJh5+NDAxVJP/
W5h1DYuiUdlGvD7PpbD/YcQYNVts1l2Jvv34t4KxT/YofMOCIDuf8SvwQTLG
azFlgb8gLD/3zoJzu9rkFOBZ240HzRO4BN3QM6Q47EeAJhFEY4JBAl0InNFz
Stlbl/KHGUdoWZS/FfuPSDCSrNNj4lI5qaS9oTe9Nl3wn64IuC/8md+w135x
7/SySJENxxn0tccpsqoKL4Bs8tQdpsy/w2L+NIMq3S2kl3UJpXkDgtYQ6wGO
5nQmYYFDEULaGT9DqHVl68m7OxGWr9wLlCu0jpDOGLsaRDNcsjhWQYH4nEDT
H6g6mCLnvG5rH1Eq6Ny2K2k9F3fAWwPjQmPoo6j7u/+HqrHWjTAHyuqQcM/M
VaeDojNV2NSNjQJOFWVyrRVBGyjGjmP1tUmD/AIhDiffH6t3fCWGCIeveYQo
VROXRcgId1tgfopdXAPtaKxC6BlRKSXY2UHKHjyrywJ1ZhN8YPKxne+SZcaK
4xS39HExUz0GTlKZTjkPVpSfkXL8XhssyQCBCvGWn89u/wtV8BjmEvH1GUYM
suhxYncx+mUcUwtVZtspUyW9/Xj31aQl6sMczo7DCTELcfANV+uQ3sC6+xwt
RnO+PXfeVm5reVnHBDWglHdLkEQninbjkFp23hP/Pb61UwakFqZRvbPX/sMx
J/Vsq7wxb3xKbC7MYzjEwGCGDJTOINXThuJZnaW3S652GNni7gMirEmKMTZp
1CibbjV/roabUD8Re6ooROKk1FjWmRNxMGe+/zvZynbbyUye2VbArpnmcWLX
A6kPL6d1bwGb1qPoQwklElVwjqlpuWSP+CL29N3x/AIzxyCrcGiPwYE6cQYQ
IxquosMRFXv0HqtyXEEu6bPb4T4zMqAZYC7v3Ue18o4Mhy7UmiPysouLlrDk
D8JqwENNRwEgFLwAu9OWYXKKmHnSa+SZYBpFQLofjdq3pmFXkZn/LplsTlO8
7HxyIurCbwNQMdjQUQX4Ma6xCNXTayG6HJxTgZWulr1Qf+lw8JTbpX8xfj4t
0C+pJFIz5HFczoFOWznbWwAzudPtxKdout637pl27Mv9YUq0IpVnU/QXlt/7
x237s+ekdirEcDo24rHPsz6IwlIL3D5cr129cjKg/IiUcpJUbbQxN+A6MGZG
AolFJ4OFyyRkoe1BkuFA0xn0QCwknSczlIev3mcAUzXuCTlxCwJEf1V5sSFJ
0nqU3ODCBaJcxJHk5q0ejJd1OsJtJfhez3/h/ILKsukGtMXcSvaRBMCNCTPl
emqfQeQx2ERneB6CVX6l4SQ71W8ZHkHx2DJZHVWTlsJu02WuKNB2S+hNYcVm
hYqnsIO/qdomgX4uhFTaG4CTmMq0LmYdbfz1xsX30bVk5nhXNHzADoevSVL/
Jp4KEdNJm9vMvstnAksM4lMgVRkXCemt2wgX9cWlM2c/i3jXPr9RUW+lmDWT
Y3rqnlrTGMnVU8aTVVO3jlojVa0FRDv9OKiWegJJ0Xes66WGFlxWYiJrbQDC
kaTuWM4TIfWLxT5nnSaPIdjax0righa3x7Rx3I6L0SOv0J6wigsnYdVhC6iP
3Xz2MPBONj/eXHp9w5fD7tVF902qHNhcAc7juCgMa4b5rXhC6LQlQLzenZAb
VXNs5y5Oyf9isrtMcTp48dQ94cPAZTi/sw+RXCisrjkvRe9+/C9sGo63XERt
WHqhNbBXXAX/k5iWjbYsJalgL+4ftmfTZLe+dh0X8MUbKUNmF1tqAx+uMPmq
XZo73S5R2iCRO4ENUXZbSah+YwGXc3dJULk5RNee9FPdtOswrvtT7kie78mH
KUmLqYYfjHZMuKX4DloGsy+33oNcsY990PaVYMeAgR7OsVMNdrMYQseDKF3M
RJ+etmt1hONcrYN7oImtA+fKnpiJEA9bRV4RPZtI0emKIrhfaBtWVhDqRUZ/
Re3ZrAxDg7pXaUq5cIvFGpAsj4P/b59HY2Ylih50U+fQBn9QzwGJG+dahbTn
4c/A+75O+VkFmhr0rON9Gnfg3FodkVp7OA/sWMhBGDB2LHM8G8EAjNJZ3lGH
Fd2QWQmE/Vxuwj+uCUZU+NDYbBNRRnXaKLzHDrVoFimU4NF20F8tFvLSooW1
zU+1j2Ql0eh8DV/0Lc7bifi87lGND/w/z4RUUgeMZz6oF3ad1+N+H8nJaDkd
zhRkAX6TvFwgZn9CjqeqhQ46Bi8HZ0kpMd/qRZo6fi2aaOcPuHriMJIQMx1p
xLj7vQWe3pHgFVurzY0OHnUvJwel4snSPAXkbTd2ug8jy2rDD/RmmIUfTGON
w+FKnrNTXOT9wffO1HNbJ5EIr5iTdtVWq58dT0Iz0U48N1vw5JtI5W35F0vU
Ek1bHE4ORD8V5meqgKpMEBvlkA6Nx4CR+i2oAqxK68lvByUllWwiRHlLAeMd
YBdkogYWcc1dhkB8vZUlJIBz9XYvDiZVi+d0xToujzoCt+2o09Aos16Q5y6V
Y2gYILwDSxuMZoWQxWjgsi6oloFR5jgQgtrqX2nXL8Bj40ETTwqLAQLq9MCL
adWA9ScAlDTNUXdRjPEZo/0T5Tozh/sMjbwuw+bzHES8K7W04tns3kIftZxP
AZ171R5RisG+DIRv8YFr3eT7m03+VnJdlHIwfhzxn3eJ125U41sws2QfdkmR
KuBzqMjpAE2zlAoHZI4EtP9qL/i6tS6+p+aKQbwNzBzlz5TiILA+aeYCElTl
8pRdo6HdMlEv3J3ErYJ1ied5pdtNISy/x1jpjxtOHeERDtM/+gFPjQoEZBKu
q8LWl74wpA7d6uuPi3Noitl1EU5dhI9bcigJHwVkfKXOr0qkJZy2LBzZH9x7
6+Cao8SgmmHKXO1Z4gvvUnLZPkSp/XqISvZirb89s5ZEI8x63BuwAJ/eopE2
gaX1x/r7hoIGrOLUv2KOvDOfE093hwE60XSUsdwE7NVthoBis6y4p45snHu1
Rqr/AkOoLn5QmWxPp3vEvr79KOBmFNhWyPsLjMpvkQLFEQJuvYpEH3HYiLCu
UwvosC+MpL3VjoeVFLCWTpRtugdDHXX54t1v1QZG/Mnr7wzWA12V2Mf96E61
hjcRZMlMdK49qxqFvKOpKQaEVrgkb9PXhUh+4ice1FeL9fksZqaMB3/Kyuwg
sZUAepuhTUXulW+8w47LOMUEWEKVz5o7UfHZQ1fLKaz3q12riewDzHIffyOn
Q5kpcNUAAzsS0GC1qjyTv4nv9MvstXpoOZhl/uUEyWtW5iVPyPWIJ6hoHWpH
PMWMwOi4Za5BLTw2dcTgRp8kupQFaNoAgcuvhZC/JKaa2rJImb8FQG5HJp8R
HA4TFAwci/FfIKFAl2T29pn/TMeJU/hCIFpP0zuYc5eO+0P4ZmGAOJT/izB6
rbVuyB0ThCeyDIPm90vJ6/nquxsb4cpTvUxbh6S52wqDFL9+DokZmDnFRd2G
Dugc3H1vk1UEMdfmzy976wcSO8eMPYUa0BpIpz+TbPTzH8Y4bdwHlw4L0z93
VGlgm5rwntZ+u5Qjt4+0ZdiiXhwPjyGSKJ9Qe/oogl3YXXFML6ej8nCbdw0M
yIek9/6UEXZfZ4YbowlDmTSDvKnwdmiEvWZ99J4xCzr54jyy81IcX9V6aRm5
RDc9VxwkMRmTNLNtHqqhu4h8nqr63C9j5udL3xwNOhoXBLiGgkvm97hWSwgE
WY5Y6IBBaPstUgxfF3s9fD2lxesY3IiD5fVIdBTEVTqmnxgdWKAK2H6E8K4n
9aWWKF3bBxD+IP6HVPLcfcAB5bJeB4uKJQLMv7kBwiA7y1AHQfabAHIsinpR
LuxV/pRe+CSw6D7hNlvpvYIot81GP6FzZJJE3xURrreJCprsP42DrqoINtkh
hpFyMa9dq3xfsYwy5o7FA/IpglfEu+NblL+XI0M1E2YFEUHUDWKDPOGaBhvk
CCrNYCHuTYUgHRx3sUNpdkH85Bt31g3F8i9Z/zMhrPsDwWZksLgBuQa4XHNq
T4K4+1tWFSPMX2SuJJYGQeM1QHGmvq4z7K2zXDnazOKRFGn2I7U6wyAtrTsR
jDoeHvBIISlq+2i0Daxgkbhqw7skpd8QmGPCivRXlZjXCyPa2EScqx7KW+U4
nsjFoapSt8zWeeNvwxVlAwVR6171TKK2OfpMZ1c0a/2uTl/xXZW6AuYXVZXp
fRJdRgJK5I43nmI9CEOznMGQLvCUlo78yfXvabisp96IShITtZBjtBZGoI30
Nn1gmamDAVG4MzurVwhGnvLouuaesjaB6XEOxFGhMUy5Br8izRl+nXyx9NxR
e5UMm4eZu73aml7SG971ecdMsXBjX8c7Si2lxtPuwyAXtF+uo2mn+vs7W8bj
sDhC4jYtWcKqpSiJhA1uwFQytIHPSOsxA9SYrOjSEMkT/QNUCTj7g+OAWMUe
7gCCB/jbGYvrL15nZlPVO+aVQxse8dC5fLEklCF4WUZuIKvjZdcdQEE5h07V
f2Qqkl5EE1yz7QNbmTJOoDo/zSBsgnNtZ/3X/BgsPpWscrTx7zvpMS8lAHVN
JuDgtOBfx4xfmdBy8parwF1muruLwf/mV2DvigHHcZMTU9eCX5YJehb86CAS
wjeI6OBCZ2sC//Eq8eM0TS2/XlHIUP5DlJ67pXgOV7q1jypaf6kw5OzDQCtF
zwm2rInY0wO0pwzoKbNi4qWeLOXeW7tQZsJVZtd1DaMB4ZW+AOk+eTCoviZw
jv8sGtzv4yjA6sQST7pg4RHzP6va8kCUyl/fLYR7D2soNDBG4C3faq/4H0lS
/Vc4k8RM7o8kQQHAvtMqQTnEKwVrifOtOWlBbABQvzB5pLC5J5LPUfYMlrEU
MMcmva4LwPJXneYpsMW+TizExdCIAXTfm042Ex+2qP7KeGTvw4e+3QbJgxbG
miTRMLwrNxqvSPW5gxwbgc+pV020IlG1WwTJ1iPYcXR4fIhTf4HjJujrmucd
Wq55FSMmYCkJsLCgxJs2EhKQBe0Tpj23y3PZKI8SRA50GjEvLpqoIRBLO4LI
084VrgVTUuAMMF+SazqNzZyrDKgzQX8AaxccizwGhVk/3xSjA84W/biBmqIY
oHT3doYblS/3pyPt9Ou4B8lqdOSnu/p0ppNiQsNHPi142L09oKWDFzdiQDfS
WVm2iI4qcYPf+1gXnjtmf7/EOw3mcnIR/A7fYoUv77bUTEHIzmgOHW7n1lAD
3/ogsC+sfOZmmGI2Uuc0fBjoZS33ZpuwiNUA9Q2S712HsADf4nVZqR/wJabW
hYhNI7hAyn0AIZNIpkSbmktwpZn9VUq5+MPwM8UX9FUJJzXP22urW66V0Hxj
MuXvDxdRUzFzAmrqZbc0UyaPRJdRR5LkUMSH05QIjcylktfFhV+0u05YXnoy
G7pspRluk6+eTl7J390AFDaiskNgipSG/lnYZ73UrxeI2UOG9AxiaIlqwtAu
+wUh6Q33088tAsoprzemIxoVDvj4LJUHEYMUmLIMa3ddfnoFV/0x4SFJuExZ
2tHRB04N1yOuWQiOz39lsPUja88Wcnz9nlnusUsvVazTavQfiAAK175usauQ
XNFJAUSh3VXGPieeSUJiVzsrqzjLoVf/f/RmPa/CfVLq22iwN94eT9UapVdH
T4XWCiq5i21SnQ8cPGUzr44uwVYxLTXUi1QjTgT1+Kct46abvrRR8cc1xlHO
EjaAcSV9F/azppW1yACHtHyKqC8d4PzavuYDwSQ/eH0N+J6ySYi7xZVvqP/r
lr1x0Luqi8QQcZ918R9zGdqF9KWPg7MuCQv+CObFjtAqa0rbnHgZLpjY8XeL
Mxc/rU25zUiqG6j3VELN3RBo1e9bksoPqbJAMuLdWN1fwVkCcV1rsNBnrx1H
wLnv0ZZAIIH8weBxlEJMDGi+b2HQvPwee9mI2FFbiVzzpi2GTWq6OdGuI7V0
23WTZeIn3KxUPuHHJkMgo7Plvq0GuspXcAevtUoRJPtziiBxfBcVQinW8fph
plDRoTMVaSLWyd3nDqO83zmGPAKWgaJvbnONgBzM1fIpZ3Fou+gh0l+l/8bu
f90P8h2n8KsViWZZI5dLVzL1jrfxx6XrUTCV+WUc3vaFyIL4WCcF27K4H24q
sqMbfDty8Q7849Pg6qhRcN7NrWv4oyMKCLlmVLc3cvDCufOfmmj3wLIc5m+J
7Pxzi6XHfKxSWm3iftJ6+yoX2VrA93Kfnz+Jx6RXTQgK6M6W3VSRSHPm+XNb
KnKLkPz1rBlCPDOxpgf3gQK1sLFdMJCfjdfUEcovuOyloYLshVgfMfhBYOwM
CFnlXrh/CXsiO7aU75Zji35M4Cnr3/xLlANWj7qn0AtjDcW+GtJNQ74Q1xkx
nY+ybIXcpP9WTALB153z0jvLtzpXv/OpjYVHwXM41XMS8zTshQQr9yUQRQNd
5zo+17gf+kx4h/i5aP/pBdixAAYmeQeV3SCwtISlmT0Ftfb1CBja9XeTVSP6
DUQBijxiEII96R1zI4b8k07w0qdQHY1g9RMcWxVpdtSwmUNH64JNshBhuLcx
my83dezxyvVJnv2PrCZt/qW4GYQkWA6Y6GEV1NjcvW/EBQt+6+oQLzpBqrAA
LJcfvoND1tn5CBWf5fbo9Qp7pTwiBd22EScg1SuZi7p9mY6Q6bZtCFz800W9
9kZZb652nPvgmk5/mlcvZZFGKPqDcfchot93WXXL0q4qBciQGwWEsI37xYdn
mmIlcdUG5Mbdlej6YCZeucJLtBCoOdDRs/K5phcZd93aZIQsDoMPbpj/GvzT
yvFaGMePP/tFOECMv4wDAj8NoC6LLvpZoWZtWGddGCuQnwCsLcHizLXncU/t
60JNl6Q1Iq+8+tB2qLWk/dJ8lIDd2LqW/iDvH+2hWi/CC2pPFqrwNzNhRl6A
hiknCJtFysgIsUQpCgX+8stIPt5/DnctnORKJy11giklOtBM60lFEu/yWQkj
M2M+XA8f/Vd4WGEawsgdaA97lGbwqOI62n0VHy88MYOVnUOGj5eynjC9a8HS
FQZWWowMje0fqZxrN6COUf/dN1D3OfKyV702AM/8WmxBzKeiazrW1Z0OP+qh
ATFYA05EvJX8z0KxHH8MUaG4nyp4xqARJyt5CTO7xg4v33ulFJZoY1DEHgVX
rSCs6cjCIZCjSWGMCI5+VWAeH9k8VIKESMRxJdKLO4uVR28CIPyhfQR3bmd+
4O2Wj2gRtM8bm/DRYr4nB51KhUsho0yEF4jQfccx2Jivp0uI3MOz3UIdAX/d
C+5bxXBs15cwBq5HP449ztCagqWGYh/iQk7uOivlhlu6j9xNm3VWp5ki1d9t
KAMkvHF44egVeb17/0L0pwqLJhzLYb+7rCmvNn0oxPxa1cYPIzii3OCPzrJY
KIAPSPDbestKoT6x/haiWAfWL5HylNTV1JZaJFtCD93mjZWS9DsrZECH1iZz
JpX0xpEO6dvOxFPqA5ghzmc3KfPet5pOE9O7v2W8CX9CN3HZej7IvcXhSFv6
5Kv+5w27QJnW4/NM5+CVy815l6lfebcap6I+o7mIPMYAQsDv6ch2LZSQGI51
pSmimPuAvjlAEcx/+Z6K2530O22ovBpO7H83X9V8MwVTGHSHcGn50HxviuWL
q7okEbXmjrlWY4la3SsTAzyQH465aZnurD9sphTjOq04RVADu9S9JPXCI/9B
LGlxBwbelcGtKWKbxVDYmNwujUbssyNWvvjGAWtqplyKeJ6GqKyz6c6jo/hI
TjZXT5rExuzPBICRpCjSWiBdEMIeeBWpfmiji2q17NkpTSUUk+aWKNaGqcqO
dMqXoT1eMGyOdcWmWLnVbRhEmoDeao2i4+fUc0Jlqkrkj/Mz+XYxAKXGG6Ow
cWVPfxPPyvTBgYDVNImK4JjypD29lP16/tPc56C+hNiYmFcrPQ6w5duiw2yi
YlugWk0e4auUQkA571etUzppY+yF3Ar+/gJUxZNIgomlGZbYImxDvUzvxNEp
U73wVZWEs8+KxQt7raas5eZ1C4McuJ+sZa2SM8/st5L/V9MS+HFuOVLsiDQZ
PyIjvyzINOt88xJUty239y3I3ub522+GMufA22gziPOdIJmT+e0YpwCMFRiz
YNRnW3FH/Aiuwl8WvpC/vPC6AdMqXAxf0+zgWysVfMR+A/+N1z/edWC6mz+b
Jpig7ngQ0AXP5Qd3FLMW79517TQtodt3ACWNZD5jnQNSY5GO9InrsK9fyy9J
eShNJ2gk2Z+KaqZIn/1jddEED52bV+eahD+YvUcyEeNXWj70Jsw2/UimRTrg
bKmqEJ+EpKb+UO6e5QbmOFaQ7yJzO0y4WyhFA/fe5YYhrcmrRtJKnDpPddhF
YASF2EgTB+rtekSA3SLoTWGhsr6oMCwS0b/9L/recSgt3tahtJSYG9z3NqaH
QeHe4Yd+Mh52hDRpNxIqTdeoEcTTZs5CB2BST/ViYVZY5EoR6x7eAR8KqXh5
xymFXAbSfPkQidIV3VaSm5e3iazeOQgu29ADd4Ze5ZluRj0JFJ4FnoVoR0M4
5jVHWUInvXDohZG4JetYPYtNI3gjdjCKXUVN7ay8+TPSp+JgRIyLyhH3miAJ
WhBvz88zzPv7ijN7mdZFZl9lW6gYYmbw449kh7AWvE5KMJxBi1Qrw9lmnA3F
OaV1eRZm7pQj1Ym6BhdYGr0PURxA00pLhnxI9KlOp/myS2GqWuFGx5nFI+Y7
McsLRG+klijCuVPv5iRALp7+9svJfmoWhFPqW2svBUPhvJhZ/d4Vx5L2l9aD
/8oK5saX3sUKb5u5ItPyl9RBkozI5zVCJuBQG8U+zNKdKJ+G/NaVduEP9Y/3
iJHabsSXCqMRirBWTGU+7h4Q1nXcz271ZPY2dM+MMQoVwlJ5iNOWfLb1TaQp
RM7zt1HEkyO2ZBkLBLQUwxirYaIp0qUm3h2uiF6qUkjSmdufsuq2BlllCWbs
i+xqz4xFD70MPBz1HD6SIMpTPkNUpmfsiAvGX/MS2gjPtTaJpPTf1HBlZQYD
lN8ZxjI+tHTE3pbguGSvDelmun5toQwLdwTLdarpivjhV3iXKv7YYAjivbdy
UXBmICsmykjqxJ7l0XT0KQg05n4prONTGffJ5i/TaKRBROjWNllEiDq1pchb
vMq/xAQW8UX+8rcH50b2CeeoiD1Qgx9iwFqqpi+UkEcSVj8LBkh6Z1FExALb
NEKxezooQTUiKFuh1Z/aZBDl/Rx6JcocMp9VC1DDy6Bd9ozQxfBfnm+pYCNG
Kw+3PQEYglTXPa5YQ+mou7/l9wLfFYdEWmPZhKFWsYnhQ6Nz31TfPuJxWiuA
oIjtVH85Z67xwkJL5DuFXIF38ata4UHtKCU22TzKs1bMv5k2qdTXOfb+6c2y
vtwRx1SiD6sjRgtI7AfoxMbyCvwuG6vD+g0vdF16YpagjHZuphw/EobhwxW6
fvx8joY3vEZ4cK8t37ap+4dot5CPXWVi4q2Y1uXnIMKV74BpMpNMFcjHvlNt
aih5JJCBymHuHbOG2644c3AbXaN073sMTfBjFXnvU3Q2fU3cGpQITifWxLAK
ukywevED6Vwnb9BCUjfRqZX8UMmfa8N6E/3z1/smo/284o8wdah3k3OOaHDZ
ZgId+EypQ/pX2DrJdRZ5KzmKLDk6ON98ucUvueYNMRzzm44srr4bNjM9UrNU
zdEMTjZGi4u0Wrv/aUAm/qi36+Sk8Qb95lZjqlQyErtXp5EroUKpGS1MEgVr
gzr9e53CEW2WLhbNkXJMjBcqEfclmJb+GQdVXwlcZ6YNky/7Fga/PmLLek8y
Cju5IdOjzahk0sRAEqMxkpWl1IalYcf3YCuQmaSAdmL50k/oxpO0RLNye2Pe
a1dcA4wIY5xoMTKEhu92a1Sh79/1txSEWUFqJLBuso8f3Oi/gZkOCyNoTbKP
heTZ14hLDj5ovJwWBWWAFvl47Lr5o58Wcy8KDBCYYF6XxlsvtZ034n4n7bcA
A0iRDf7W2JrhtICa5qKJfCDIH6WYqYuwF1g+0v+iEAPqWQiiWmb3yPCEwM+0
Ja5k8JIKmUVHj+DTYDuT0WvRnjXuf8bEplR3ooWD9XJouxr56NQa0DxbG9t1
x1nH3N+aORVCB7Ei5B5lKik12QcwBBP/VV2c+GZBYw95qgCuOFifYX0ThXzY
mZZdhj4Ui2S4egCrhPLQH8S06r0RbPq5512O+lIIWTtRhxfoxSbrql3H0FLz
foCtF8v2bIZBokg2Taz5H8bCbp5PwzC87WCyHNIxZmyu+MfhbWbopiXpyzsL
WRh5+qjkHX8OPRk5z/nJd0P7JnDoMPrxh1Nnv3J6vK9BFPuY+j706Vsoejvn
yHltEiwV4qsKkYnd+SJ3RTKWVfkO8yyfmvvyJWIgmIHbjEi+F0FXAV0Hwq7C
WI2wEvCVR58Fjt240zImi/k8mDbdeyApbS3eqyELUUjqU0yisHMrp5MNTmek
bAWL+Ysj1AbN76B+Hwu4y40vNI/O/hE4Ln0XxtiOb1t6/thkZQLRc4gwcUh0
RsguMNSv4IZRr1H961HAT6d9EyPQHuwe4ni3YQG20GvCtTPg3CVop8fzrFI9
xIZK2vFyV+NqlaTQJ0SJC2sAZElLeSIXrJpgX2o3RuulV5zcIx203eLY/g+b
sdC7vvR+WtrD7IktGkI/M0k+xnwFP6L1Phcmp93vpa+aQJjNaJcyyziA7tC3
KDAfbN0GXQTNHlE2EKKhIv6foO0lQl7SLOs6mes6b5Id4Spt7/ZyW388ngjI
CSP8nb8Syq85K4Xm9FJHvKo6jfcbeBOnsVrm2C3yhvdNzPjWj48/ktUXhkoS
iY5LlWTc3Ba3X41rPHc8Tb0OCcR97y5iJ9aLw4h9mhvhGlb3JHOGSdtP2hqe
Jg6lmW3xhnX1Wv5RJMEg7f3RwhA4luMGjoWHWA9z7NA7Kve+rjRIjUVZeohl
H8CFIE315WavimLu+X5M4kis84b+1kxjjpRXJAD5O+7MceSNEvvPcKIE+v4E
8bJA+sA2jp+plBpa8sUbdtXlb8DNYJ8pyb9ovcRdgXucjfgi7nGd8CS7eDJw
gS3BCBExAYU5gG/wsftuSK4zQXYHdpP/fi6KF2afzfhRHrftk7ea1OZDvr8H
EaEmmN1oO0ZXBXQJsdfCfLhNDbAwHXI+fbFuTq/R5r4eU0v01mtjkqa5YpTX
VpBKITySrzE7/Qx1E3tFCJoSeEp6GppCh1R6VSLRhxc0jU8ngA5rEJmvRwHs
tMW4JRiPrCNRnLJeT3WbIehzk7TcX8Dbe1mv1HIPjRU9PdOPMPrkUsEcmi2i
4fknGuBvK6Kmmo8vfipZHCd/3WaWNhSaqPUioKzRIggEn4iBLOzWmw3q4HKi
3z/kSvT4edl4RUZ/NClwm31RAUywmrGpUPN7Ce2Sv9DPDgJwLLJWILxu3v0o
YKsFM2ZAW/HzkUlZXdJhq+eGC9QGFI2SqyaOldAUF9ZhmvghTYtLvPLXuLpU
w6BBtIpjH+I1Knu27rAVkJ7Z3giPhFhDJIZo3gxEi8ZQF226kXgnmJA6NLl2
lzPgeB4gCClcdLZPyS8UlQwTM5SnjhTfFv6FUNPJ4iFP+z1FPneqTgUJOpSE
aOgCcXdXyW71VuLukEeyjKoe4r+lEa9tQayHRzNVMJalmvw43k3Hdf+VUjwH
WsMw7ymZHWZmS1TkRj0M59nnEc/kOZDj1Gk5WQ3hLhlAUFkmXCJRrb9XCjkf
mIDysvteTcuwcW10dO6iADeAmyaofKJJd5R4OT4+D1P9rimi38ecEBE2sg3P
wtD29grnpCLUcdCbeRY28WfxbPQQ4C0kOFWFXepv/IRGmrHiBjP9nU4DnN4F
fhkB8lWDfvjtmFIE/D09VAR02DwXdLpQ+hY/0dK9FzVfCn15QKkPF3vrRe9A
WFqB3Z1sN0SqbLXqWW1nMiER9nDuPp6euuYmbnMqTXkhsg4EcNQF00Lrc+yM
KkTn+2Pdc8rsspQmi2X31nTx9FGbE2qLgiA6Ak9kOO/mld9hILwbuSeTZ27L
uU7wwHSZpq1XdhihH6tdZK+LANmu491BzmJuVmfrAXq5z6iHYHfTga4anuC3
LwqymUh6D1OQO8cEsrEinPtepEEqWGbzn9llXA+zBcTlfvTUPE6VxjTbw0nt
sWjJn7M03cNyDL1reoWaovYHYJRqxFn0EwOvKQME8btSCWmKHK/Xf21TUU7A
m20dvANJYPAzDDpnZs/a3eX+NIca1099E9H+2Ntk25CjOmoYTSM8uXo05m5z
xbCF1KUVvdVc70rO9NbNQNGBGha9Vs7BYGGajytjav08hnGEl0Xb8lFON3Yd
vNrc6KnocZndXglvNECNn2KjLfTz905d8Ra0prU593i3m/+GxHOQXkT+x+Hm
IGrIIy97k8kNb227yG+4J9mVgrZouqqBP/luW07FvuxRdgHO6EaOTiM1a936
d7xgiv4uN11l7LWKhEUkTePVxA2DMD3N6ViQZSFqvbJJXqpeM+XiqFvfrjrE
o3bQERNHy1LyR6jm1YBJUpuldEkH/jYsXSVhZOQ7yXiUMFaXXD77b2kwSafd
GWcgiaPLc+uF0lpYzRvzcK+tI6j+mr0qldQMC7xXgzSrAEi0gatmJW7IolCt
4aNFylKfUOv2hq0YBfUXUZnLC0IPcBn1FR0DEyBJhfayvB12Wuauih3mwCai
+I9Us54UcyJtmE1nRio1M3ExrXFdbOQHf+t9k3iESva30nARBHDdT3UQNg3L
O00ti8qI36ujeH82LFct1oVrJBabTL+GUW0i8h+F6ZWX5MMxZRS5vAemytfD
BlKUit4ijauXu6FMBANfUTKMLZo0Bx5htJdzfitjzw9iI7Ca7vM4cJTdd7iG
OpERku8KMNLlr0R26Jj0WD4+E1YQfknDdIWwOy+dTCsdYxtoa6iw4KggaDgr
+QpIaCFkPlch/IgA2dkWdKWRklr2TJvwkpwWD68sAP6Ratx+qtiZYEbB0xf8
N3NBHrNFBUjW/A/zB+aoDWR+lA5vnulDrbFPNbvT47Y06Jurr2aBSam7YUvR
xDsnslOmbT9ykI/Dd270epSPgOvYslRqHl+meiyfRGcxXNYoltGmKBwuB0AC
kvTKpEmPfaGaleREir8wRGbc0HQAVCxsv3nddPgf35raa2MsCNHYxm7d9pWV
t+OgYjxDxm5g6MVRMV60x7+TSox2IO8ZL8ts3k7NDS8oz+FvU2/RGj7DHvYi
8sUkyiBOdmrPHkxnYcNQPHvDJGpGHuc6+h5UcLEXU4sPu8ObCqSKVur4Qqef
BHuh8C13ztMuBBxFb1Bt7YeTDEWfoMF+9tiBHxw39d9fBF6bCibd5XWyKqAK
qjFu9dIS9pYqFuWzpydJlXhweZ9bj3Eis2xil1+nsEdrjA501urKb5OoSQSd
Y5rpGAX8iZ9EfxseEAkvdkGi+G3NsyfG0MjDks8+yRoicCg9Bt5UbnVxN/rj
9OaPANncH1pPzzadwyQ9jXTLWCFpcvG44x5DOXCITJcpBUQUV0zrkwWBV9Kc
A9gwYT9+CoWMGfajiKSCWt6U7GSPcqEiAH8mlB1qDtcz5lqsE7sAhvnQ61kV
O5FTB9KlOGZeToQOwJA0r6pMJc4PNKbo9+H7GO+3TaIJmHAbBFtNRFjyvfSj
AmAJD/BMlH0bMZDyFoQoHojMZRFO6RNhhe2y4a7Cv+G8/LJwPfWJkbcOMJyE
Yj1HJ7jCz+1eD9APu/YxhCtMpCpv54UI6Ox65hoVThDcPslTQ5PipR20cclY
X747zRhEhpTxM6DKZLSkDxJXx2//BOQzTekR50m/3SbgHY/ABedB6O4Ldu6a
qcyUmNPhp4W+ZB4wk/Iup1dTqUM5lL6/9fGkr8OXJ+a7XTTW9ZD2VqOIQ8ra
7dUMs9WiP/8GUTPtmZ3SSqB4fxklSdkl2hznxfj4XjMIWmNBI1yqAwXSh+JA
kAJAImC7aIyJJ4jXbZCatGPBxEZO13jY1A8NrXc1Gr7uSr9+LO6e5/X2R9gk
4iwW5UWr+dbFzh4jYZJfOBjNW8vg5KAOf+Rm+HrA6QqdxvEYZVT3GopLXU9r
VtbjUU8laWxQKHx3927hq1AF3GCB/1LrK5nj0F5s0iPdHnA2yRbRUiPxNYdq
StUDEqnRvUQIrLOVcc8Di6i2kjUPgmhM8CURAyUFe9IIqJgBMHekz8CgJwJx
fTvjDhDRbdT5etEspZFS4xuso+VtEGGwXsiS6s5hEDUDXbme5FDEgidNMOOP
DUnHkp7s6b7ig3B0GPq4l7e3KUoRBv7p5lUAk+pQEnAUVP7NBMkd73iarvIi
M3c2VvxkftiLj07cMDOGpfswbnCBSgcG6K/9zTBc1hUjPG2mkJdCZiOcarI1
opnhAw798I/kULyuyZulpEpHoYN7Vt4N/KlAmoUB9VmTTbHH1mvJg1ulhRiw
vZYcjyGLGHEfcEAAClLT674GXfRTEdKF/mXJAfBefnu42q1ZvnyPBdsd96gb
GqQ/jFOcbTl5Ba9aQL/zcd3rcIYboMUjNypNWTos0kR0EyMc0O9yL7uyFTit
JInuHwAzI7BcGXXw4VHi2WYgBdzr+lAauYFFyJQb3sMc5NlHFMKrqMi84QkL
N0tOY+IIjPfMiEuPbIi3FfAvKromFAh8NX7+bMVFymnnWPPAlv0C/Upx0+hv
JT95dHQRF2cxywDrAxDQwAElpr0uK4pQWt8b0xfSkEqmFxmNZOM4nuYIkdNR
ECyBe4RjZjDIxXdeeu2shPDp4zSqUalh3ZdIhAoGTesOK9gLfIn6H4VvwbRt
UbalG17hmpZr7l4z5fgpnrNIAoQE/OpmVg4maNq5n7vc1rGgVW/+v6hGBYHv
pNbTlzfuZBzQKLya+4rVnq6oZ4HQu9YRPqDwH75r518OieDWxWD4WtLd38bF
XZMXcD0MRcM4MSy2RO+6QptaLCAFHY3ElzCGQ/Wer88Bp5Y64UaSsgSJxs6D
1+eu6I/pSnm8goKz6juHYpoRwzVBDj+M3oOOQrUoUgXXK4LWZG0gi4+Mk12v
uWh+G6athrY57tod88OFaLEQBRgx1P8+iNLASB+P8l5W2wDhNvk3YAScstNO
vHgvEd3laRrScXyl8u8lJLshoDWGktCPQuULB+h7BtuIC22F6hPvI/d1Y0QB
xQpKRPkB/9N9J000YRm7dvMLp2H4bRR/A6bVMBxwEh+1e42OUE3nq2tQemV3
tCje64RHyDVRWhkOLaJsjTACQbRmm3jY+wGZ6r27dzp6NwQ9DYy6P4SG75sp
G8NFPXk7xkXaoO/wHmPFhwUXMxSM/dUQA26Yj+aUBxm9v1tDGvqZ0E0FxqTg
cD1L2iqFLwjquTr2Wt6L45FrAGuHWmQ7dQ9NlN5qoIOD/yvaAxIGD6eRBavL
GXplcHgUG7pEY8/FLgPCdSsvp6ZbHnvQvIADdSJOlUQsd4tKnXZhXYDdpMdn
dgUCg/FALB+il7Wf3r+ZWGqoyj+WF2bkQMp/OinbugpUgJdyq2I/VwcWOivR
FnQyvURq1re6uSjXMYhwligjXbFGpLCsUdf0FzA0q/gO4f5v26NOeWvfa8RG
NsK04USc6agnbBA0HjqCn4SEpwYY5ThKhxSYLjIvX0wr0B944KSDHWoByZ07
Bjq8xdGB071thii6q8UIz32tu7r9wxUe2yBP275NnZ0IDpH/BSdrM67IpMNB
B/Q/3W/8M4a0raC1/QC6VL7YtcEsa+TNqGuUUTFRQV1hu9ZxfN71zd35d9aF
oR621eAxkreWPh+w8g1dtUwkivhHLDO8SckgZrYJB0dew2Gvr4YBnEiIDDcW
ve9t8CSXtcaAGI5FtfPVipx8Fs0ow0EtqRryDBzeQVIaSsI1Vm9t6mMf+wll
BvPG50QO4oRwRyvMJeBQe3dxrkEFKLofAKjmyha5E2Ge2fjuhHHSnqBnu2d4
yhc+xnkc6jryZrh6RS37VcnxrkhdNOYSAjDJ5uE9iUhhvgDEySmUG2gIB6XO
q8QA+M3VSh/oIwkseNIBE3XQHAAWjKE9uUvjIcHx/EjYTY5M+4nYZtSvZ3Uj
LePsnjHsCrbeHggi7w8FpgpDUmy0TxNChQqdLEUpO6pQAeBTpYy8OyAV1Z0g
0VTK/Ndysqn77565IM7My0kKie85r/gsZBdp6XDp8f+2poTO4D92QVh8ZCu/
YaqWSF7rHknBlQm3FDJ8lsc8sjKoJkyB+GBisxJ2LvLkqZ77d02g8UUGRn5j
taYM3AT7BiJ0y67peVs1FUAzS2IvhuIjEy8tudWvUv0KLHupUn8Cy2C1C3Qf
d7oqyIttvl7L6IrB9FPCpVVzV0kk/BEkEQva25wpcz9O/mVS7YFG5eiHlw8O
DSShvFNI2VwGIsQFSdBR6xnhgvX2VyCGzZNcocQW2m7bX7lhllOSm538nIqN
bOdi83xxnZ1a4265JnWS5NSyHqja7gJCYnBTmYPMqb2ouMj1AF+n4yKwuaxH
AvoioVmaHf6a3aEkxsa85aCdWfSngA5rDySJWkhjrrP3/evykJEBG2r8/MnJ
lckiFUnt3Gd4k0Xkjvw0isojZe48lXQkGDNUR3YuzgSE0dKBz0LvdAwTh7BR
17eslreO7CzKz0xkWLzPhMoOQm2QHC9mhhewhCt+fCzhUKxGYZnC48fcpv7b
uVnhYPl/zvF5yV7vQhAx6QiyFNluDhCjPjjfS1rerkhGq7JOvqtgGSu8tmjQ
RX4aYCrL9NtdLUa/9pr13LhXPRigSo16DoQWICfVPAT0HP/7o9zF+JkMHuNg
IJoCwob73dBP+1Csb4OifghKsBsUIzaIfuwcOBLtyfWXaARiY+ezaRscyJcb
8iGBY3hmWQueFRYL5wUHkVNzAWwXKTskw1CtC6EXgubDdKRLTIEqhGKZ0Ypi
QNlS2dfir0KmQJ+Qo2l5Rv5I5VeiHrYijt1ByAEH7rUwJPq2+Jy9afZxIeiG
R5qDnHyL6kJqmvRyVVs01y/So6aMnCmPtWq5wHW4P0LLbsGvWwNn28kbiuxZ
6UE+p0mhVzUyV5OxANUirezxfB/yqTA274oYDYGFk0ku6nW8bsrIsexdyTOM
qis2sIS/r2NhK1KlXY1CbKd9iVZq8mtYvJx1PxRhMETdkkcG0lHtTP2PMKP1
Og3xlz8Wq6ah/llCjTbu1B2YxWM1jOfLqG0pUEndIrSx66uiWrL6UVw1mYTy
EbQLssTif8jWVzNvyZognjOQI4HByhBBIH61KSWeL4oUE9ksIsgGKWIM2ZEM
hPVaBGSm+i0kxAaC76ZdkAD2nnFeXZzb4gaQ1iC62ox6LjOxs6njhMD7SiXb
ddG6hv/KtU25fLLDu6g6NEqqeZq4EGTWoC9pK/PUH6g4YW2CJWS54pQ3Eo6u
+OgH8Hc5TkHT7UFwZxJMEw1iQ35eGyfoxAayrmfQCnwT03XNGeqG8euRkiDF
e3y1RFxDZHu+UZqHLGeif9eWuP9rlFQvk297o8nnF3dBoa2ZC2YVqDcAEYwc
kscmie0LjUMoJiZ862NqXoepFlZ9ZsAcMl1HbRQUPYxtFHzYLDSAboqtoXkV
g2gMmU3t6By6gjDLlJhdtLoL6D/RlLWBCTilu05e0WOaQqU3IflkrZ3pGZhD
RM8S3n6+3JVKkQRfRM2fvKj7UKLuLVh3QD3B/UGNgsdqn5qBBbHBHKHlTTHb
DPwAWiOECOe22gCcjC/DOP1x3UPHKg98+3oKsNpPB4be8f75bSfJ9IBuI6TC
ZK27GP0kivO6+4FRnU38lCfGpqy5stlMak26YxM5unjFDMYguoq3Ysix5wig
8JpAimE+TjrecuVpkvx9jgO5g/iAwZkG3vRNDpOEHRBMhbTkLnxLqDEstPNa
Qi0WmQ5/rEb/PUwHYKinZWEuE3wzuJcVEuTatilepX9FxddEhFqVExGZrx0B
i9Lal5xRk833c3mVD76iWCSMHsedJieiDra1NUh8OdcgdKMsL5UyOJkm+wNV
0XQNNjlMGPtyWqV5I81+NqSXU3FOY66cbCOUgktrUeoHYGM4NiEylpnNEcT8
H/4Kt9Yqt5/AoM/06z1DX2R6iCH8ln8PXm0H5MCI0g8ik3YF+AwSoSKpIxOq
rWybGTtY1Ue7tnecSFaShLgDKG+kurG7+9WXIy9Tn50pukZz9BBL7XLUd9PW
SdCA4JAi+Hi3VYjWYUNR7o5hvDKClLMZxCSuLxz1nlKhJJcs0mtQZzKk6qvI
h/dswGVVl2mA5JCrJCp2Vz3/dDKbdEx5Zyj/qjOND8+OOMTCK0n6wQIlLjvm
PURCLOx6UZ9IpR6jSx3/EhFrVEcy+Lz6cgKgEeOOrFCHqLsqyxPNa1wD8MYA
3NNdMYgZ5/iZuya/DFFodwHJ6Lo1fAZFum8ZNKTBwd0B1cKjUzKCdmhyJGvx
TZtY8yvxaJ8DV1ITyt60nzbsFXujdiZJ78OIwbPP6PetbUhVA2gpUMfoTJs8
Qebb3b147CaEIE7xVF8fPOuzqnIND3ZfrltJYAUCbr8YQZOfUE7TuYhQ0ZRL
szr8O+x+mfLFwFimRs0z+upPf8UyCGUgkoeECw9LnjX2sqfQ9DumomumirNH
IcxiklGCt9clGkt4D0cskXahYnSdemAMIUVwm/g8Lc68b8p2OveXx1Pk7gw+
q0ydrJerhYNlofYmZXBmq4Pav+ovcoBTTbmirgIXRtk5+bznftHy+ojHH/1A
VDN/XpyT1+uGrdrrdCcWM6AE1cplCI+zkAyvEDHbCnNbH2iP7f8u5hUEoMWv
UvXxNW06QBaE3e3KFepppX2JV67fgydwFOtM4sQGX5s1ckYKCPpPGgrjatuF
koGvcRKvuPm31MokhAjnOaEciGuF/fGZXN6Vw/acDjXZ4daqVRbBEaJ5CTKf
oJcqeD/mVkwixXD7DBscoEQZa8YZ9wMfy14JA0nF6qGJjFokUy/JDPy0pq4m
RD9Od6tFBHLHgS8qiIwWktdRmLLjlEKBErLvTcAE2aL0qQMpL3MgYsoVSYKA
XIik+GOVCJWP6BhZTRuW5cs9FFMjRhVfhXVvqAYrkvgiys0+ltIryV6FRrrb
zZd/JVC8aIWJL+ohjP0SYPvbmqRq7urgt9jZvnj2XTsqvL7/avkNW+qm2v6/
IKKWH8uSTTEMPz0tzILaORCS8gWLogLp14dLjKIBm//e+zpgPLOX592lUPQM
bm9fsvkSC4sHvkQf9VYi1MamRQUtatb+DnHIHPGBwb7iILQL2rw5LEMmjqIW
Eq+COd3CGBXWi3iD/1F8d04ND8Ej9jqkL0yu+OT/VkOgBKAvLFrPfXG9rBmV
5AiEqee7oVYELk6Q9K8zWW+d8TG2a1yZpnYbv5CujkxKUUqCG0BufqYCd/zf
MfmUfZB4zzb5lhK70XS9IdLmSHy/UrXx33gZaXf+9qRjieqvoSMqy7j7YF21
s29sIkdk/9Yk8tk1N2z7uAyZsqKN9bt1glpgIjjcGFbnFHK7ARPRoJZE+LBd
Ju6PNqRSFTeZyZTUMq9FMV3yZSlr8SEbkOveNyPm9gJFHK6EG1mIBrHEvskf
I5HIgmQb9K2Gdg4fIHcxKKYGdy3JS8menDRsbP+WJKLGhAeckmyoHakvnJY5
2MUJApJUIdjCHY+p0Hlq/t0X5K8fhsPlqXL7vyH6/7IF5Lxj2Tj4BwLXXIQ7
dU8djuVfACmz/L/F7MjJtLlgdTSSwXlCJgKPju4Uyr4IgM7mpTflnc29jZe8
enq55HkKtp9uZsyFFtly0ddmA4qymoA3JUnvoz3na0W5lnegTssg/V89B1gH
6M+wUtjm/uE5QjEDa7haf41lWyc0utWIuXFuQQOfh6gatpMoiHxxKkeyV+y5
ptcY62raY6vSJtAWBlCzK20+gpA8fuj9JsRN1K364i/Oip5FtkHfl238uvre
W6zXkO3Aems/tJVmLxHlTfXpIOjGPWW+SFeid/evOwt/T4ThYcf+lpOQqC98
OD6JiGc0rJgqTlW8Nx7nmFdsNXFLxfUjSQmOTPxKbHtVHL4uC6vAUlWusNk6
M2CakDOXUlXynRG9OhYjx/wA8Hb1Yy/WpKo5tZtVg1cG5auPtpQgkRVpNkPU
LHUhopw66dNbWumwg2EgUhMRJL/I/mbTzV+rsmtk4zW7wnRycxv3C0A8srJu
CFlZ2I3nYuI5DE7SQmUx+b6RKaRf+jnnyxpbq7QptmPnmyuM89SdhEJyzASO
2xPNW1HvcbqWSENpq56JBevHvLh4O1TgcOihECv/2McUNmJsKvgXWfCkhy1m
O8h8ned96sxN4qV6MByOIKkv3jF+6y84wLyEgYpfdBVcXXh3FlZR7r+QX/iY
d8Nf56qU5Ik9t8RrqMKw3znK3xOVyQavSN5kTSX6Hbt9Ha5pcetM5zC/GP5L
/248ylkmKDmNlVezQjO+ic7ZNgdQXsSRrelo810Z+/BicimSLj5TkkXIaRtf
ioWoTPk0s+qfj2nn8n5798cnU/AezO9YsKz4f6YB3wvPXmtaZ0ZxgCpOlYQz
Spz1n0UBm7K8fOmfb/tY9iSGlqb3ui2WIPWq9h34dQcEzGfWG7JArSxRHQYW
ohDXpAGK3DcqVKHTTSPZOWcvkG9su7dLcW8e07ZbHxVZKFb60HPsAaCgAtet
TzL4K6Mz3aHwLX6KsUgWqUPgbABQ1QpqJ9/LRvY2LmA0RuJ7tHf0ao9YRhci
RYuCJXnxqJXhP83zqx9gUytnwlbJPU6lUxh5QgnhLpv9vKp0qYyex+Dm7dPx
BRAlFv/AkjCzb6zKndfE6sxFmHdP4dGt7P78v27me4kfmra08lWX7AhNsxIG
XXZInOk3oOnuLbtgjUR0t09eYJa9LnRSlNpcTXxn2iJzQ45HUx04vtwYSSff
4Pzs1p5aQrKgGLtq/88tco6UQ2v24d7f8jwVCK3JePjstJ4Ds+7JxVTqwJQ1
B56vT6UWY9GdtDnDkkezxp4UGwhfojJYblGT77upNmvPyoiYyo6h1hatOmov
dvRmYo0/Yw4I/KZ2DL1XYEoVgu5kxROzhUir4wUYcEJEkCSe54E6qREknfmJ
4rGcQLZhnvHt2qwJ71bGxAiS2AbznRqctjS7rEh/xS4G/bP6nNmuHUFSopK0
jrB41sUvnddU5YdgIqq0WeJW4U3uo7+g0eNTZqhOttuNug/yxvK7y2PSMxvl
p5LJbsGksU8JkRlNBBe+T8nousrdhTKo23rThvGGYvffq0rF9VGAx+TViKAY
BbFuH9bDrUsGLSofYb/p49PT8+mjXN3zminaYb/B+lAwxie57ApTxXxDTOpz
0ua4pa+tMQPNPMIJLquO6Sg9ykzttgZQCcMiWt89ZogRNUpZkRuBGtYbAgbs
jnpnNC+kdYROK5fHfzXuY7NeGwpW4NwLXCqOU1KxWEtHhDJY7h3IiisOxqp4
M1LzXJ0oEdfD2htkBmJFVAWJTPaWWPB0P9ZShWgNHITntGamznf0/ghWFix+
AB5x2gR406l+p5pmnIHAbzDO+jfzgSCHlILtIXl20CBNCeMRcy/ZSxuNMVdx
V/kdhU070ynIMQpmfgBAovCxBy6L+EGcKzGZFj+ms0d9LTCiyLyr5yRH2lZv
hhY1Dx3JtXebmSXxi5lkQeMuLkNEsoOS66Nx8U+lHsk0pSBRbwtYZN2ZIedg
Thc2GmZ0DoloELlOqEQbBUWfrqErIzOpc4Zo2eK3lZru5TICREP+i5dtX35B
b/y61FzkClYK6D0C4pXu+hDnVSqI/Y7eYn0lA1hvWzibubLxPzQcuTdeAhEd
OtLMv3o68Q1rDGjqOld4xqUiFlBhd4LgYFdAq3DcgVLnT4HkwkKhsvKk8QbY
UPiPO8PqFyM33yKiQdSLhp63KvF0CGBGVPsNF3IucxywAeS/ga/xgwPHp6QA
Q+0206ojgyLBgx+/JWN0vHmi8PIZdLuYEaFstvEo/0XPNmDvSaSuBPMII03l
tJLxuxDb9tq/3WondnyoPiM8jzW8kOmvIEKvITy6IhihVHRp4XUSR/oSlUyb
SqKeTmIe07z3qTR9nf3wPd96ZNCQl48MGBsTbupTYv29kOra93gANfM6E2dE
4KWAysfUdNwyBebkVgTmXMhAZdvmvHgsbulvwYQw8kjrb67DO6Mzh+lQ9ehC
SAIkDJW1k8vikiaqo47ICf+CFG1/qRvajyiTg0xoIDon/wHePdiOH12h1Y94
B2B2auV4mto2SYWty9DJ34AQrXpLf7K8BlizLl9sYs49oQAaD8V+oATWxFn4
K8sw0C4E4LphJ6AvZ3Tf/hhOwS646sdMV32NxCM4LcE3FA5iRhbjb7ZtDEhz
T2LFA7Cv3u+WO0W9BeqImRxmD34JPw5XVSOdB1wT6mhSIzmckMsjomO1pO2M
Kg0miBQyVWGbCazroh3z9pw7B8OY9k+VUg4+bQZsEXJVbj88oYpxWAoHdsE6
88UAx/MeRei4D9R/DFhafOhDU0CihYAc7+tUTCcxfk9Oh/PO+5skmz5p1oLP
4RE3iBC/5H1fMtRBwW9+JxKvcvYmQTDGg7w2Ysg6a6I0oQain5RHk2l5NGCV
8J/jAelAGnj0zYdXfSna2nmT/N8Q7Z5caUIxcvzNhr+3nPOe16ovuC+ggw9i
iwCnhue4DR+b2zJmRfssLb1y65+hbL3cBmNroc2sPNuB0bC/d/2fzt9c5KAQ
HyVEexO6oT8/kCzIXKaa3+ZDWStGxrUdfsZ12Cr4j1e++e6QZFhB3Smlad6Z
/WaH/dOxDqLxwoaHV8W7Eall/LAaFv/e0b/IBDueB3YjGzcAQb8I9q/i8bo/
5qoTjiPjf/9WHV+ML56V/SUkqNvcoUeIWfZyoQDzJAtur0riraHwUabBRzmO
0X5CkvxRhba1X6nle3X8Ntc3Zp2nLNKUW04ClipefI6JjxMCX0K8asSeQQih
upqCSfjQDB2iwNSIcfb8lUSGiBoQdRHliukCxd1TkQfRONUZMkdQOdYAsEdN
m31XlR9taQsEtcd3GhstHAr5PEHZKEc4vTpPHNPINaiWHhBWASrdYnxqdzIq
xhJNYD15d0vkMGaK47cnM2GVuhFjdqy48jvTdb/oE7i3xqUGYEy9e+lkbn1P
zoEpnGQ2ADMMuoyQ6+8noBAvpe0xEcZxvCL7+gxuXlOnW0Q9s99B26k3Bung
CLR8NIOjILM2M3Ls0pc5jue9oV8fbsLJ898d2eOa62gtUOYZ5/FPhh10QzNU
EQxvj/ax2E2C37mI7qiseQqLGk4PtZc58CM4UkeP5Rc5LDJgNLTsJoDJ3zTk
67OeyV4RLTwCKzVUcscvuJmyGjArS3op+aXcw8MwT8c3N6sualNZ6g4BdZbz
1OKWdt71uZ8ua2VlVeZn9X6KHDSbtGrfyt+I/ZtMsBJ+d1tLVDuXR1rvO3Mk
KOKGtOTlxYQ9dFfGlvASljsZhV9woPko2LbmzTlDtKX2Z1jiJ63XVeBY5GvI
3HdtEI3Gw7OnfeXZPSeAziNh0i00eS2GSsDAmaZSgr7ZuwO7D7gc8CU/Rka6
Kpd1XMziKszdzoAmeGTWOR2OaMm/4ZppOWF6JRqc7S/ADwPWnsCCP3i5xGzL
/6HPHEaeDWcIXh3INOckmqiCQw99Vky+iEt1+07FzkcyqJqxJf+JyPE/Lg6C
gzl0M72aZTFA/kxwI/lyspW1DZnbox2ZzlC4Q0MlXHwPOxy2zlMptCeei8mR
ED5lqzfHvqG6X7blb5TjBfESvWlW+qf6LCaRwZ+ebhq169STNAq0lbPkm5mN
RJjBW57TvI1RmLBuvq1b8+sJUbii3ReXhBSQYxsBDcSavdg9gSsEnYWej+XM
8tvAXplf8WmIEkIMWOs/0b+noI8w844KwU5MMrx9pKU+rjZO/RnyczdlnrGr
E7rI8JyZICziWNarGub/pgS9bavbOpEWlshfXuw/W0CyqyTFve9vD1BxG6cU
slpXB/RBmx5NRwpucl4mdQFKxfpUTbyppmhLCXu6wGjeD75BoFw+ZNNJQJMl
hfu1SyuBx0jfsiBNXi/xkmwv2Own02FrvOhARekYooEC1uIFGcufUGBtEAGB
rHAMBsdwhIw0QzgHf/gdX2MZ4myg3ICDx02cIytJdGNfZM/sKcu0SUvZU1sL
pjo8Ga0Jwvou56Lv9PtgezmwHEPwYnv/7fgxaaRyJYbJIRpQWWOhIOZR1qjv
IFnlqi4q4OIdJanaaQFdNWDI+XF5DoKldk+jnDYFhg76Lz3ps84M1Kvg4Vce
0PIYxo2WfvCDNN4mAUcyxWGZJJ5K1HAtFLFJdHjzmL6YjlviH5VPoGpezp0+
5uLp3OEb02MGnQC2ESX1q3d3/Epw9xOlYcueE3EUKMVz4IlXjBzzJAJW6K5M
4igUt7f5DHPPj8xh4KYyWOw/gKCEdq4zuFZWWC85sikIldCogrQwsAxTvaTM
KlluF8tONdfaR21XD6IcHaa3Kou9jrJS8+frupTcaoulo/m+9rlWilyAd3da
cJhR3n65SWsm0WRe3jGHfVkXzrcoYwwwAsgUkvfAlNBT1rshcNqlKNnH/yo4
nRlKyx342oVsRtRVqRxgBlOgMlygdiszcNcasrZjsDjJFrml6Lhz3kN+mlSD
iDZubgU3wx+W55+ADZ7ithUkuNzbiOnMVdNwY0O7J+71NEw/CG26cg4XBkAp
g5b21OipkOLlz6Kud1A8tLN0ilOgZO/DbZtsHuF6VsS1CsM0Q7XW/Sv0UJew
ko2azUwxPNcNLMqWp+7imk7qxgSxxDQVx1SPD+oueq1mlbD/ULufWe0NYLw+
qSlDA8dGpVAWGIXtGeDpnCDJMz5TTbG4Ys7YmK6pBE8iUNI/RkS3ruZPCeEF
KjFHQEamphBEjLa1b/XWWEv+ueZG4vpyetozvOmYJPslCqTL/TU6a5POTwsK
CyrvUVP4h0GncdowmdmhFEH2BfxKfCIUdLfWL6BiQiP9Qvr4S2froYgrmk4w
d8vzWBAHLbh4QpCM8cpA2RpBcrlcjMxFaycxo9/Vp0cHrD0Y7TE153kvbqPb
efRjGV5ZteUiChpseiiXHC9PNcuhZgCsu9nV8l/GqRTJUKeP0ghtiaWiDOam
0Nut9Ww+ll6uohxc9QcbvY79IeIp3K15bD+QuJRLSUrIcv4pUH9PegZEmgsg
KxqtT0SMKwneAgaasu7rGt56a4fpTunIGBWrc1OB2Md5QVmYP5WGdbjwuF3v
8iNF9DfL9cjDMq+WSKTn3bolgBMjlGGdxPE3elm8YkRaW7DMGR2gc3MIksI8
kJtIOx9OeWZNxWUfXMXX+GP7Q9UpW3HrYYTi7iGb8hzHuRHk6fH8GVwSzzU6
zzhqYX2Ffs654sOTQo6LiLdByERa/JUfSQ0gFWxh7VggroAOs6nX5g4cYaBM
VgUTgg1PdlBRccUUK7W280DDUsLtlSzR8H2ussjd68lIcj4ug/kg02RpWtcY
UDHA8TD1i/qnpkNCFFcM0Kj+tGk7YriTFvpavMsAdFAya8uBVyJdTzy4Qlvo
nh3ojUPImyewaW5BKJR3ghtcsSUjLcP1DmTqQEvA/zD1gRBT553UiF7Co8d0
8n9X2ma9WiVcWpa/vDY1b45PetIdjHlgtSNjBzALAVbBFcCXHQY0G1OEf3zj
fGzm9Nu03wxuyF6q3gOgrA4WZAbT6eCh0vF3V35MTHMK0hY2699+L0PJ1ApZ
JOwGwpvqQwCn72LQnbzg6rSwGlpXFuDeNJ7YkIZ3FOpLJvxU8bRcSe4Ilt+G
VO/XNSOL8I97026Voj5zsA4Qi98e96DQq4Wjv+/vpugnP1dRkCgd3Vt8RDhm
fF+EreBHRsRsNhi8b5ti8j4zHz7wUzJ66nGqGYqMbK8CfdLBzluDNSoPYEST
QtURrzONAZB8sQ5Oc3e9y2d8AbdJqwCda9uxsVhrt8LJzkES7J1HviibY2vC
GLqGUjbQOM4oXnx3S2G0MY5yxlPo1Umi9J30aLdeSmKBVvbVtIN1BVL5Sb2P
cfR51GtFYE+oOk/nWGfYmv+u1+fOaNUh5eneJPD5hYa3/SQkKBl/v1flXfZz
ei4f2inNuQIYZFd4dZefzZ98+ABRMsD40yYLJBd11z7FB/ap1l3ZPX9ewvCN
Zeh35R9gBkyu7SSg8Y5ftiUiuhB8notc5MznYizREfNyB+9ickq8WL8FwABR
LzhRt/r0Z/7MVaJoucaiglp+sKMVE2a/o+k9i8mprMqoJCeqKnH95au2XMel
fn09w/UUNjZvkyee9xeYaxTUXWreLeU4eSOuQdNiA2Oy9TtpQMcY5E4kPxRq
HPzUAFj2YpxUbgSZ4frlx6ofrC2eVt6H4h8o5KfuoU4O3a8xASN7F17DUNO/
Z1seL4vigv67Mt2MtawgaLjvFfcBejAx1n6vWAEMsl9CHYm2vvhYjJRpjf+L
qK1LgLIztCAejO+Bc1ScHkt1LoykWP1SksZB0fdP89E5nQADX9OQiW8zQhEF
A/lg0NdRTslMu+IrHiL9hk6qkPO818Du41gOIk+PZsFQv+aXEX1UBGwZP8Hc
ACRdgnW3vHNmc1cGt2QECI5T9PX5md6wNEfF34vuUIGzWToQ/PsUYY6p2pC/
1aXGatEk+SReQrzNtZevje4vh/KNIiBorDYioxAdFxDcnLkeMSLG24+CLVoY
iz3AqmJTYBwwBAu4op5mYYl5I9sN+xICbCGR1bOcWTuizwXBPu6OhPBiM4ss
CthjoA6s2Psq7CWUDz/Japb74/Q6QDNwdd3Aiv3NFpwZBwcAyqQdDRhffbmX
9wq4XAj6zcb34biQy3ER0PSiWbG1XKW4BTn7T9BuqKaTMkwFEdSH1guj7L3m
9Q4Man2OWV4OaQ7SZbfjPNF3rh/eYGwDAhz+iQlURAppmjK9Iy3JVYldtH/Z
Rur4mFd9Jy4LIKvriOwcZOHxH3tXTI3ljtVeaCBQrNKsIlR8fBEF6l5xJQJm
CZSVWvUtWTS5eesXonSE2RTgc5ajOTtcV9QYAuPDgKyoVh3xt+rj7QQcgVjZ
DOf9Am8hpH4A0+WT48v3JgVWJK1cUL+tdNZm5/JO71bwQpv7/nPjsF3e1E18
JSol8aOCmW4EUSE6GNIWj5yZXSCA+2ZjeMSOdAdxbFFDA27D/SGuqMKMLZHQ
7aFZEJbZ6ufEg3B+ZxSomJ5vf1cHPEZR7oHieKdHCFkzOZdmqqTU0fGObU74
G70CyVT7MjWcXLbe8+cwKJo9dUEEpq3KianA1UtKRlwJrbIsmH41eNnh9GrO
ALngJef6lh8pTOaYTI7BwXR+5MBYQgOk1RDxjuZpsfwAVM8Yt11MUUiMFays
oPJSa8sJQ14lC6kDkqQ68ihVufV01wcabUAmIvDjve4DQcXJvYdBWAlQB0NR
3JzrbDoSc/WhIoAH2BPGRsX+QzRJfkloL0rZCXr8XTYRgxPFDAPliUHaLSmo
yi3Tf+ASeCqT9If+RQQZvT7FTBEHP1PG/eCJqx8rxSZsa2q5iCvDwAPLthup
8CtWo6wYkkMXH1VSuse3nm6ck3VVGY5r3gOyaA+cZpMccWf8p50pNsRNh0A1
msYYo0q9k1yhDp4TQU4BXD77JTxehkUQIyA+jbkcr+ufJBCeR59q7hd7wqFw
5146omNYBSfI8MFRAi69PRp4d9OP/d7j+FzVgs2n/m7o455mEO+aAznBAynJ
ztnmz0n+OlFDxDhYWmdTOtknJGgMV2kRFdmWjugVoPd9qQl+Y5uxmBXioWtK
d9QgP72okNnd/yZzYrzqOz4GHfRnUoy6iYC+SyY0R/fqbqVKUY7xK8nP1S3r
kZayK2H/Z8s/Zt/qlvSjaBTlt0FmVRLUwpnOh9pF05M/HBC05HJH0ojRS6Or
gTZrIgRLyQtMEsVvj6qBaCQvJlbWXpMlczTmto8nQtPfTm2f1JitDnhNXnEj
ElqeiZPQtiYA+o9dP3sNI98xCxL/AFkXgYO/y1FPRSh9/n8Db2mr+t+CDsWI
MiKlaC47viqx0KE4q+lEQAaNkE0cvvsElWy9KKK/mGB5Viz7+eZZM9CXF7Y7
/Xiy0o+yndaVwzr0wdR9u/e7BLLq4b7J91ZsC4qw+Ru5NbF9PgopE15nc62P
0vdI7SeluH8ocDwbdrOvQy61kQkpYhvyI5MqOMDvQN0I5N96XPBCPYDMkKU2
uOUQZ8BHP0CzsAGv5p1ougNakmpmS4Fh3wgoBS1GvRSn3YvYCqaD9jo/8GtE
uH1ka2BMclRM+XF3YjWR1w5yfEg+m8ixABnlucP60sz5N+GBPv6N8Zut1UTK
+QsbNL+5f7iYGvv0PK4kzYljbuLOGeffZ1CeyrxxkwpBmLMmEkkEMU/9fXEV
bZpUNEbw+e+lh9R1trUsPeJrjuikBBMZ0XJCCisQYaF48N7MYvC19BhNnRCN
8Nc9ELxxjM1pcHQIgpCHSd+3aDskmp6uY4V7E4sQR65HEZ0t+IeWhhIp8UbI
ZQ00mPdyXU7tDoLqGuyYr9yGWg4WWRRXfsPhUOC/ukSbRy1CSxI+FiGUoDe2
ERe7AjuovFqGwBx58uZCmYtx9Y/Ul0TbkGV5SAdfq0j8EsKCWn4K6r+Sg32J
PmGB2BBftAO9vzCYjF4Nr/a+H8KGwebHZFlvPwCf+M1Qc6ixl0UfXyrPO2WI
DzRx6maiYm+JrE6ImC2BweIkfk6lGluofNqlMxJ+dohF2pdMveeEnHdcwvX9
NPYiNC94srFURWs0KnKwy1JReIzQYSpf76UqEeaDrj5nG6hOkmesyd4qVuTD
uar/ZAryelDqmsggNj805AHx07HPqiYGpZ1LNAHSddq0oOvoyNj3cpDYBnMw
FwMwfHcJW1WLIDMp/C8Rl+ZAMFnCFkRo4a5RWrYoA3N0hCGlYxsnEheFKmhv
hjf0+S8e7/kYkR7hpImQcwA2dVOdYje7a95+cTVtBkzlYUef5fhdapYWFIjT
vWvt3sh9fZC1ySMorL/y4yK7CaBK6OQ3aMLPxC5ZKq8E7uLVPRtdl4tqp/jh
aR56QwpprQM/AGztaK7RJLKqKd0njqxgr7kllNCMRP1fNlZHbWzLj24SnFPM
6Ilbbiq723VJlOfsjHpMp2MSds8sgmy/RjXAGeSJARICCPPJiiJm+7PKe69D
CDL8cQPxkXmMkvVKVZyBWJ4ffyLrrtj1/Gnb7COjNdaVCyaAFd4wmCMdzeXa
fcGr8hD7XPghS+K9Rv9jAkopJbrhuEiUhZxqSBCQLUxZY17shoYQys2+v2ch
oCeHPBmy++eugCI0YAUj4CLBgEXcu6KJGBXUQPfdwUUFHlNTxDa4EUBRoHBy
KgzD/RODxBW2ZIPvib+1AxMNkZIBOgH48rjsWgd9KG2Dynxr1ORr+wKXyAdk
4n3kzyII2vEIKPWy61SX9Ny6uLdim4+5iMNAanU/m+a3Ccco5Ov1/8WC0X6r
2s0kYMrqfBdKVGABpmoj0ErePTifbeiaj+YgYuNNLAF0imJgfhcJTfmCRGDH
wU90HUg7Vz4jgE7DzTBpZv8x68DIM6U58A7+9V8u6H/RNiHbJAnhFnaxUFiI
T1r32jvu6xohNHs7d/QgjXThfZXFJoSfOQBDBygLaHlHXexwe6dmYF/U3PcL
25oU5lhJQRTAHqqpchtdtZNgpznNImRpL8MVzXNC6AV6MtB09IT4VJql9i+L
mGljWrN3A1N2P/65lV7Wtz5ujG86qoDMlRZXVAhQ8OkefXRHNg15RwpTmHxb
ZHdQzPbQpBY6UVHOB1SOWPECoRem6ZrOsZM5LpvqDxEEdXK64oqH1OzaY9Gb
n9U0VPvq5Uu8sm312mVYOfkJaro3ERUh0NKT7PMPjrkQih0s2oDlKOJ7xQou
MWNgYATSZmggFCmNMdqG7dGqmQ6a2RzYPGCi9tu0vJutGyosFop13d2gFnWo
XNBQvrrJYcxJjQzWGJzBxYz+F5Bv3VzW3sUiHlB6KVJHM1PAfkyDIaEGaSCK
so+lfHwDXQULO/YxYVattLuzfkJsXdF+rcWcevHHq3Ag0+12dZcQVYKqL20d
LmePdiBojz8AVHJ/I9mE0UfrG6NGDQx59Mj/xnNW5Pd8EQ8wbXw1kTjys/c3
Pd26iL18dPbAI0FKw0En3pLRNniV4KFcYT6YP34WMaNseob4lbfnyXYiDfQh
vS4dmWY7hREe1HlfNufszeFDhvQpmXPTekNEBQAjgT8OGbXct5QNpUiNdulw
31xOIfa+Tu1nV/z46XD+R/CHcMxneVkiAW7THTWp/hlNweZTZA+9hEvf8ls4
j0cdnAgmA4xz9gEBqqM4KNKkjGVD+1vz6JcY9FN9TWV9IitVwuWDMq6n00eD
FVds09aT4zFPT6B+/I0MkVhQ2HAizTYTfNGOJ2KGtS2Qk8xxr+xDuVS/PU2S
2hQ+Ry/AsJSPv2bIELxUVAT8xXTJjwvww74h27o633AFwB+oGV3WDIDgB6SK
WxnH8vgaO5HIv1EK3QgJKvemDiJ2mNd/vH06dDxYIZGufei0bUpQWliPpIlT
EjYXZAbRqksvzEv8vBv5jpVw/ad70YzzrgW/dDPMGMRX9Q3qcI9nugsvZO7c
OQWUiFGDXqe1W4OlzWs5G6lOzwd++Lb3jXTPJybkTuvv/iNxZyc5VVb9ScXR
oNDS6uYhGaS7EmF2dFN3zIZPLhP1b+83lnkfhkQ+4IxfFzE4u4cKWiu7gfju
x64HoSwVjm8X18GjrGLJLuCCb6san2ipI+puB2Vfpdhqu2MpiaV13iPfvwUo
Cj0b/sSp2s7xpNj70OATySESi6gv0ow2o+YcnQLB7ytV9dx3lFKmoZpFfbKx
nYf4+MfuLXF41laxKh2vtQACL7+AzJsCsDoPJo9cKwrCqkvK18GpHuDpmbhR
KfTfIGmTXPMFnd4ABfbbH6yJIvAyBZ2JIF3ws0VRhXnVpmWeGvNpuSdqMYXs
A88Qp6ibC0ajgRj06XsItMuJ5FCj70m+bNlzJluuujrXlY9pVtoqoOyXsOgQ
WGZWXQ4tHrvLhQ7oHbGwt+OIypOz6+S0/QZIHrbJ93WLFLrQc1GsvAaTW+Mj
CniPt1rg3ajD1BbPBYPcu5wQCBiZe4XfYOYKL/uqVr7Q5BmyKkxiVlDLAJx/
OP6E2OXvHDgCDiDBlaXNyO5Nnw27at5Y2tN53fC316GoWxZNEmwXpA1c0gEH
j9k4YrY52KUgmDx+LZR7Gzt536JpkfiYifDq92D3qSXt8UVJccixPH8SQb0x
kmo5UIKhGl5XbztjibM/syff4zKCbYy5daR+ooboYJiUFhNdvZedYarNwTzz
PFdj94AMPswjh34NFj0YdFEZlRXFJmfZLE6iMTSGN9CdFs8b7KfM6YICMedg
jamBfpIsN74J8r3g+KPQtWrS54G7XYrRprJmUqPFXaXtaMYOG8vYiBjt6l2x
b6NWV8upYKgXB9Ttg01lqXRMzdQcHe8FHKe3+5xSdFV4mF0F1LJxU85QPVPd
YG6/9FSDF1I5gj4cLDkT7AUJufwDutLSGyLa7av0EQbb0YbQbYYZm0ni/KQu
t3w+raVBdkUvKYmVaaGpzCXkXimpRrM1jgONVSDa4pB0VW0c7G4MBfJ4dLGi
i+TNVkAopTRtLXH5fJtZ6ZjHyFLNUGpQloNLsjOF78A+llkfUestioMhh0J6
375DNDrTBaU3+SdViu/bAYU3uHNTJhzZ3DNsF8nT60y5SacuI+buDE14E/PY
9QK4ceIpSxfxmIOMqyDbbzGoVcat4W/oiW1aMq5Vi6YcCNy/ndhDI6IdkZQM
tCqrIsoF4fbPlEfvbA//vFBydbR07D/1YrQcOI3mCbVdgWVpd/tYxPo4Mntz
fmpyKOK8FcENqSzL+fy2aBjNKnVH+4DmzkPtniPdzclXi7XwDOesBpaQS0Yb
PyZ8JiqL4DR8iVW31TUwIK3Oz1CE/Rnqg6qTb9gBIKBz30acFX2kpZGmn5LV
pi4yotry8qfO3PK9ii5sKO8HWKK5vOunExJtVRijn6EV7PmFpE7NV9f1YmKZ
LfAC081s+3JQf/9JhSs0CQ+SjccMy4AIBgHpZOnN1v/WszBJxVbMkyZrMucJ
HXVB8Dr/oMKCnwjfgo7U2LMEwj8NbJ/n4jx+Fn1tFKxYeBjqrjKXDD0NPv+w
grBgYp0psJIg+oUbUatVOcEtW9KZy5LVlDA6+l5GR0/VGTmIuomxroYQWnp9
fdtMmGGvQzP/MpspoVJEsuVAb+KcxhdKX7aQU+6Yn3GQUY0N2LmYSX5rSjra
1U1Ie3yS3KX1y8LpwYCtUqCuAhwJoea4EkC4TNaMKl0Vps+CW+v5WqCgPx9B
TfNl2Af44i+ytod+UbGUmf54ALIYdCwZfjxDdM/1Wg8hGxfR5JkkBhjiFZRN
Q+1+F/0HOKk6raWy2MRaghMGvip8UpUKO6acU7nGcE3kiZIwF6EeV2hEVF4a
4Vev++B7rx5XSFrqgu2IKypniofThSx1V/dBH0RwBeqFliJcv3MzuJhQRMhT
ow3O65qMWUok5ROr7xeL4YqHN/ZcQoPXTsNqwMRH8Ja26ZwPMgfkzAsFDu9L
jqcqrd3CFjFKS6NRi6aYfk9485nPhoqJH2BWeul5p1xIc55zgNXrT07bLsN/
Pz+TIdaakZCzTN+1EO0z1XlAu9sJa0FDGRxm4yjMnNm/14l2rcNvH5i24YzJ
NKbnTq321ZTepUTCPtl2I7AzFB9TLuoeRnhB33mP1r9Jj1RowBS/SPJaYJ8X
OVk347qUwNmhn+ksh/IUzEGR1iCp2zbybbLyodXFbiW2M/Eewy6UpsTczTD8
DP5aQ72PKoJpV4oQn4HAJAj62w+7jphpjBxD++jKIENashzNVSwBuazCrNAJ
wIioAG1FsZfHxYsKtyFjN51FGScFQrkunEk11TexVLb8EskxoY0w5VudIRMq
nWM6Y5DySN9nfx/HZ7FGDOfWtLREtRin8eL0MOZdj1jMFgzsF0ggQfDG8oTQ
o/RYc8I7aQ+roIUt+c/BByqQypLatxLgpipjRQz45RHrXb5BbgejRZlH9UAx
S4P6CbyIw/laANeskc8za8FAXITP0qCdJnPdgK+AdIxGaDpLg0g0E+KqoGxd
vhxQbXbHMQKt40ZZpGGO78cVXknpdmVbP4U6Wl1eRP/buQU+72FXHnAiC7Hu
S+QIxIBI7/FZ8IOp2n/UAtJpaW/ZS9dcRikYWHTggeofKGyAPMf3/UijCCo8
R6SzIC/lP37l2qARMqcYUP0GhZne7npcDs13P5UmXOIuS0XwXom1Yd58Hm6z
buTHbIBDJQBtP+soRxSR8W5/pCWDWcUcrXg8ekiEjENLlxVt7L+KGNjImDeV
vvBzx8J5Y4ln9YPNE0pokaUjtKxHKdqtlObuHwgFxDAr5NPZT6Zzf2asZawi
3IWEFELfg9hhPaWYGsTdKNxMY/c6U/+ZNrHVUCOLRg9RTcSzD43a3n4P2Z4H
uVn2nq3tcZh/Tejj1SmH5v4IaXbl9Vt8Q9WzAz7lnZjP9Wa68+7eci6zhHae
wJgy4QtM9L8rj4Zn3G1NbPFOawrrPieEAG2cI+Fljp2OExXeAos39uQq54/Q
bYn44T8TsiLjk37gDcj790aMZJ1H2BxiKdWqFUcDoYU+0yCTQc3jDZOmW1Rf
smCU2iaSEhNX1+NWLP4/90CdbBV/qydGiQ3r6MLDetrNRty+rgQqgkIp+L+I
TUvUpOlH7kDKBWmfYV6O/+k2TAAKaNvzFouZma/tJlX6qhBUC7wJSvZ8ReGO
7SJOeW63WH54Pf5W+UYPB29DSoHRkaPhcmiqoNQADIJb3HAjEywf6lI/8VL2
1mgMq5B7hTsuo05oRGSiAr5XqqhiTj75m9Apflbfy1HT6rfjufx0zZYPrQt7
LPJNz+SM1VpiMB5YzjUMMwp1PfaynTjRID/ihhYfU3IlkTVs31cukuMW/7uN
TmrY+RdhDfzFbX0VF4obJZuZWZZGmrPWj0LMGgxFuSFdtNmOh+cq+o1ftFMA
BKqNDVi3cibOOebmv1jj9dofBOYuRN/kgeJnqs3uUcUii+Wnj3JJKUBgdK4X
cT1D7blTOZJptwLcLq8Aim5A877LcGk5LWHBkaoWx7UJxIFrBGJVzMjQJfZx
VlNNnLBVHxvOPDL2Uu3J7lvdsUYHE/whobj2u3dv4aA3NHbxZBZ/+hq7mzUj
Xipvk61BukooX2Zd/5Hdi0r4p014vOFCXKHTXl5bwtdxRgu9fB8ILOgx9Trf
/gJF/GL3PxT6nXPxvYBciItXS1H4rbt97Q3GHbxYcL0AiLwGTAQCS1xRTFUp
pOZyaBkSSxbS2HaUI0OtPSM0NR1IUHKp83/Sm590rYOGBX9IiGLV5fonCNhx
1GGkqt6+yH8IfsCG0uw9AxB2dEjQtCe4Iuf1VU+WYmTUP7rpBTcFSeQa6s4S
SWRzpfwv7tPp9ma3CUwTvDnAIspt1DO2BUtEjmpgAEsPoBrJPnZ4aqnaGMXy
+BY5fTbKFo/swJc0krobj7GPl/WddyGtQTo3WC4FWpm+jy9k64fsQgXoi0hf
hiNgWgfH995shw5ULK5R/lGCqD6P0zlLQoL7SXhoZVdBslDG2ebnoxyj6mKB
wGRy7bsEAYw/v8U5toc/EBd9tzdxvtKvsz4icWiooBORre25GjMaTilgkj6O
0i3F5nlHUxn/qG6lm4e5Y8nJTQEZ2jc4YdMkU2ODikqS/zwG4JAejCWZhrUF
9rOor1hz1MTH0TfsUYqzGniWeSqcDmlfzJsbCh6LLeP8YxmkeGe1SfFu5reg
qoHQIGwqbdrDpN71ZuI++WnjxMyt5TpQUrPmu3rmsUnKiL3pnIBEiN6Z/wqh
58Iqei5j52/Ce4Mh+Js9+fS8MMkB0/E4ayLeUF6am360d1keyOqgeipCVyJ/
q1I4zD+xRmqqwrj4xiJqYQFPx1YGdoPw7lfdLS8TQXAXRVcjOygQ3XbCKkW4
VAtQoC/t1mc2Vp5RQWigzbvRRTNGY0REKv9D/+R/VUiiebiR7RzyiVGxinnA
QrH2icgsZ3yFT2m1v+LYsHR9+nCl7iiruFNAbJzLM9CQSo/pC3kOLNLn2wux
3+I7/+Ol7OQSJ+JWYPw7oAA+Uq/dc2FMz/UfWVESxnVwRXYrbAPW363yTSnj
EZ7WwdDS4gHnw6O2iCBJqoHcCLbSFZ71/yAOi/Qw4aFu6Z05vElqY5/gpX+e
bHQRVTBK1roxOztub/aefJqRmopFNBTd3+OA5MzEfnXZTstDUfa7/wtqXCbw
XkFQgy622d12+XX1xcuCQ0jOdiKqNHaJ4cHH9Sjok221evxoPvmr1KhYrc9f
ftLuLBcuu0ms4TkctsVG7mR0JPUq76/GwkvKC/R90AXL3iZyHwn2GhLeQ574
1qlWSn9fNl6bTPNfGdW6nWK8U1HW7QH0Px37Sarp3AqCR/+lnk1bh+H5guf5
5DLI37Ft4ixhmLyLVQBfBDW37erAcFsdmgeKqqVnZg6fZ6ZGEAySgY+l0Xti
/5OXio5jjgzNlCbukAsq79saMHVv4ncgAJjzrQco0E+ky0iP85piBAsvBw9B
nTHDXaTUmHjwdyzHf0NVIWFdkNtILHj7qzVl3hTXLc31RciBtdGXu7Jao4tc
06x8j9GmSxXdtQ4XBGoI6YW1mpdSFjr93zp8FvgL4XQd1Zw2LG86KFrgjC5u
4ZeROFPDRx7K+j7yb07WQw1bRmAaQHyJBEcY56H0dWjlIJvM1NLB2nBmMm7L
qC+YgEgfXHpPBeVmlaZIqFsS3c+X9livVhigvS6e2Kzdaxm9cTLbfdxB8Wnr
Z6bj4VkMGsa2DWO0eHffvwsf3vx7sQ/tm1e8gykfa4Q+rpCiJzuLZ0jHDI/7
33U+KHNeBt5TjlAQ0YrV+35xhPP1VfH3huhYCoi6dRtmN3hQGEe0KtiL12iz
m5xs8Od9AVQha8/nrVy4tP9zNlNvjrwZBy+DnLLHDLQleOTD+uWFAkaHvkz3
M0/tGl05F3ltEBxLpixrWQdFOTs8irfuMLjp80bJZx7b+uh6aGTKuUdhC+oC
ADJ7VENzbDAf43AX1KtBOI2YEIWRKnF0RzLF9kGVwJ4L7rDCngn9JTJ7DFjM
z4ovrUV+LvMV+3uXf13IuXSRr1qlR3qTLk6tOhDXIFEdI9sri5pZpvi3qbM2
8JK4/XLqh4156De7EBdfzCZBPjJ7o0emRmtcsH05VQQ2KLtvK+/r+9PSPK6f
s0+SFizwH+qnACbeBKGh/CIc00c8rgJxaLoM6X0nIbIq2DMuaqb0cboX4AK0
Ao6esvCYF55V2KT1CudSKGK8J3pz8zUMhCBbLTbx0GpIIANwq4ytqA5lj1+M
BSocc6TcS1v7JojgIj8l9tPTldTHXHa8GXUkGqCDBGHdCuO95bAJy6hmhsCz
SsbAoi0LfVqMBZmQch3dJBXHcT+Nbs89GAXRNy8aOzzNZ4Dn0IC/7riCS2v2
KEbM5/LNREf8SIcBe4R65huYxOGf+/e9Y2XafXdCvm5ngzXMB17/IKV2LG4W
ZGkCsDtzm7aaqrJkdVqztPn33XI05NcfkQ0iUqZ+VDa1vxfNFPg2PaJ5+B2g
8RC/EpeZBb+7ayoBZZNBq8I1Vcengthn+3VVl6rp8fpm2OX085zDSuVcUPlx
/fm7NvZKpfitK2ivuXxc47MQbONZhtcl/C4eY+dtb9/EdUI5w3VWGhvnn51z
MZULoDqjCXktpYK+7Tlw6VkVJAk4eCzLt30VaBS9sUGT3FMPVzBvd4sC3xWz
CLCmbNcsmdc0gj4ZmSPpV2wBi+E8fI4zkoYjk9zqnDlIivJ8I0Fux/XV83cz
MRR2PVa8IEAIfoJgbE4XC939955cDOADCMY6WGMwo1fTeGOXO45ShZDbQpGs
n4yKpppFIiiGFTar7HGkxf9LjL9arUnTnaAAHZC+/MeqxUgUEx5H2lOgyiM0
VxxMnSi+d6YtYaWIkLPGAw9NIvXjVVE0/POgoPt78UsLAQnzdX05xrJePEd4
ePqKGpyEePvhpBRAihU7u5NsembWRKvX9GikmFWeFmHBkiRjWzgK1HKGVvJc
rsRgBDBymK4CMhYuQpPlNnE2RjpnH6MugkMHd0BZGWyPXf5dXBc/U8JSCzKM
FTRX/tmXzGjgELIzesImg11usQGthfX3qwcKvoRbjMZebeVnZH/M3IfIuDmJ
E7WFjjQ/t2ajKwNWnfJmMsUwySRM+j3s1ZPMTByk/GSt+jMeZUgwyisIu0O4
myVf80CVBP5DJNNOi7fBsFOXHbGWf6oDCuDKjgWOGKPXBkN2FDBp5AEW0nWR
B4KgBd8ks8cwpZargPWQzCwpsE/vDw5Q5CtNeZbx418wEUrEhZuapkvnVbKj
KJw9LcfHxKnNm2EJ/cwD5tdQxKYF2hQ9MTdbzVucOsgDxR79uDSYfXt1aydV
AKP18DTrDtZkaqbw7m17spt/TK8LOLD//QeyNRst7fiDSI73rU7so88VNoMj
sRgtk8Os+JHkFUlqMX+e+h26tH1fj5amuXeAAfJiM2girb8+sKLqqLxNzCJP
se+8taLuIh4rForPzcZD9ee7eXqjCb8mavJoWqK7A5HSWkr+L0DeoEKhGB0b
2TIfkgJRzWs29V3Uez1hLmteFfUtANZF6Y+GsKSPEVEwrBnjkxx9MTZ/AmEJ
4xdB97ltQuR+hwtf3yj83enSz2KhEJfVe29eKZIe6mneOX/ULxHUK2//QkQb
WuoXWi6Ek5OqFnLbTWWgK9ljmqZbjnw9d/m4SzPRq96GoIWBC9PjT2Vp8gb4
BkzS5Wn+/rY1JBqHl/NMDuh8dcjD+XudY6J8dhd/sj0jfS6ZCcQRMQTCm7OY
ZamJd975fIqzl0A3ZKVCDzQzVyZiR5jobPX9rz1Odbbh/eaqrGvpoP5GYB5b
S7q5VD0VJ6flNHDY94MpBNZU9NDIa9FC/zFv4lrSPKmcwRJQ4ZxHiikf80xv
nfF+4vPO1/IT7DlqROuoo/fR+mKlWHXAl+D7FtFN8ek47lMO1GygjiX6e1To
buaYP/HixQf/FWep5GmrgByZH4c/Wngr8iOMUs/LXEw9iBvHVlbsHkToXt5a
TMPlL2VjqLzqyZuSSlIBzgqYfbhPYhiLrGd+s8ynaoOGRSUg1l5bc8VVHWIp
sFmy57owt8lCe8XrH8/vTJcQ9D8kyx5wht5YREVLfdrwJYFpqSyqp/11cyqu
oL8XxJzL6Z10nkddpdAgoLQyMPmb6mdOPHjUpR336OOsGyozKEGnWKgURBXD
7jj92jOU0ERNn53aVKP4LmmAxJEvVBsjMb6HY5Ic3er9FxJxiigwNiS8Uqz+
mHY8xQ9y1h1ktGmmg6zgPC2j0GbFV3VnQQhtPF06qBYsvD8Dt+DXzJ0g48db
QRj/1ZdTaDHv+6erRt/wFZb2cihbGOf8vCS6SBGNHWQbf9QuyJCNqTI0ELTM
gaOqZy29svGTciL/LZaH/dFs4ZVOSVnGIupQ/rPZ6qdi/w+w8kfPQLjv3Uy6
96j+B/lWImYXwaJSu+MK7Zais6mAKSRrHIQpuU6mSjWmG/hmjnJEy9yN/9ww
3+aQ2ddqtb0+pIEOq4U68CghvsgUBKpO4AKZHrLIm9nNhhWwSrOPvMj7iQF8
wSdz9tyslK9ydPv4GHvVGYOE4LC7rz+WeZ4X4fu/eaUET96zXp9m4XLw5FYs
U8rJQ7B/IPUiJXsxKYrBde/DvR3zNBL7OvlNPDYXLGXirUmnLJ9MfanRQhQW
quKMoKBKqZcYBvVB4SkwkJLklDPuVONxGA/esOluLP3IhpNDubt2AyKc7oX9
78A3Lt608TSFRcHf8A1PDhm+6kpC/8KGoM6wy1t1veXssuEhhkOZyNL1WzdA
jPUXuNz/Jh7I6mtbqMdTqhTZouxuu3wVuZ33TIpl2D2huTPOWDXJhEwgYdKe
VGJd1thuunHgmUhZt/x1YEsriqjsGQTzOjPZmtHpNa4WtecrMiGXnkNXyQiV
/zlAgxoCo1G3ApS9D77YxLU1g9//jmgKJhBz/Qlr0iaHquXPGHFx6LcNn71U
ytzf130TvRHRB0g73DZqizUcMr2JhvJyOknmi4g7PZ6u3AQUSr4GOAKNBlXt
j+fg1WOs1cawfdF8sDkBnmGwUHOEe1nS41RZJC1TSzgAj6Z1hGABMiWjWQYw
kYuOOh42dZzowYAaaNtebNQqTkhrVBtqRvrfk2n32HNEtL6u7Vz9fH52UB7x
NwYY1KDzTmI7TiENQ4rA1jud5LPoO/QPNOJbuEZKp8KVGt8uVaghHb32j4uJ
d77TC1427mhOlSGX4VEpzZY85P0K5WzBolRQ6c/XKYPbx4DinQUt30CSRdf0
DFjZWA5pnlRQ7Y5WPHRrpf4ZFPibqnuivyAqHhCmeo5ClTZ/yy1HCeEwXpWY
+/4UQmwLiUgv91UEJJATv87Ymgb+UttZM/nFTwasL4jN1Wh9EsaM722vGaIF
Nz0t9hKcMyZfR4N3at8N4FITelZvCIqH2QEaJ0SSAP9tFPK6NJ2/M+4c7yS7
em6rIbBKFcB1Kg0cARnbkMg01lAPO1RSixAQD9yq747+vFgrwWJXlS0oKHXY
NgF8dbHYkTjlzrKg6BXR24xYOg59IVarkBjwT7pUjwOeiW3ExyFJz9INA3uh
KTTltKI1xi36ay5MF90rp+whNpLTg+W1OFg0E5pQIQWl8zBcQU42e6ks/GXf
8FQCXOfU5yzDfpSXvnBilWTZEq41fu8xVY4TFk3SvtgZwsc4m98lPSLrr27L
54orcWxnVTh/Fs8VycIavxESk/ZFkrH50elx+wg55jDK+YeNmRlXdaL4D5Vn
kibtrtBd9/ax4aNvrlYoY4yhN9X+SGpw4yWBuq0vaUnP9Ll1hK22TNk3H77/
AC1a0DvzwHDjOJJbFAsSahlA3h0h6nqlsXM6kCp0spvxwE7/AcW+pZF/QKhE
+i0A5bqABChbfLherBa417yorz0mMF257fQavxar9b3anplVmjKSUi+zNkOb
ZGoO440g7r+gDzCX+D2ycIrJTtn7Ftu+rd28jIA6PQzg7nnhP8oSqInNOlDS
d7xrMvTvCOdfuxb6ow0OTYMfP3QP6kQFCHbKgXKeaiMlmPazai+N/QqQHK52
Cu/6bqQ1wZ2nexePA8zHmYWJM+fKKdWyyKU2FG7mS+kOaBSMIOIpft9zG6Ce
tfrvyu9B7LtOUr0rjvGUT0MTOK82VsU2iMQIoK+Yv1T+O/akzacIDO6OTvna
T3iuRDWho22hC4Gyk6Qb7x5kR+IV3eEgyi8CmWMSxbeCFpx0JM8+TP6NH1g2
u0CNPmUjXpg+qrR9sEAupyV5plSawoTDbNiHN69p3eCJFRWae7TQbfzLwMn/
rGkiJ1NbMYOkGJKfw4HKCQmyQwjFZoiknvwfnajUZODm0vHD5vwxy/uukk84
vzUs5cM3lzITuwwLogpBOVzqULdUAFM4u8ispCx35fBXWtquevCk/eU0mlXU
UVQIf54Bv8Uf++WLJsGJ3OM25rSLw7MHbY5rvOk6JD8OUFJQ1HLDdkaZaepr
H1MTEFJYki3Jm8IvPgeq3ZMAAaT5lZn2G+uqrG12Xuu/NEc7FhedhQPQnwtd
WyRMOeUU6ywpOvn5SqqNXk/GQYvhxF7bpYsWbxxgCUhT5/pPDLzXYjcpJpDQ
S7sY7A1ySPIdngeeuOTDk2E3dduAo9SdW0bPT5m9CbuUtAxF4F99++DbbIzP
rhqsvYc7XxJlttUjPzSV5sOZW+VqFQNve7yLSnp6fSm5M9PUip7RmdcBgMTg
oyV1nOjGWWpVNrmYXJMvUSprYIVqL338kPpi9QdtMmVzH4Qpw0IRJXtWzqaK
omHkDwQpyYqGk4FaBFcwJeBAITReTeQwabD0CEt30hWkvl5NVmxY9u3un7zp
Z8fLDGJiLYeYJs7ediFSuYWHwh2EdjmGkkXEEsdAvB9W0+kF49NQoITnxm4p
Fh7OJIRiq6qlyEXDYEsk2/29zwCW7qTVnwj/bRt82kSg9EK8CGJQDE05pzlu
MKsDNHBkDMtmtbbUiQGcIZKVJZ5CHEq/SO1XT8ZAd5Gg50Z9mYhi/Ip8zXwP
BarEr/fKEu7k02Gt8HLgwiUgt7GSPEGexw8lqFtpIPlNkwKtXx+IURFziRPR
msS7pTaKAw5WUQbbDl+5XtoYFeCVtsOCG07/el8fOFv8tL6xc7TDwNQItAce
KHYGdDtI++j9OHHXs89qFcptWA9YV48Dxm9vHmDF7XLKGA2D/gxIsJpM+1D/
QPC5CAbDtf435Lir/f3BIDzfvsuZ0LUyMQ+Y4AlhZPNKgXtxj5rapNdGgnjJ
GYNveSZgcvMvuBbpU6Yf/pkCENZ4zrVu0Pvl2t5LxJYM7B1PhjkbjaB4ubfn
G3DfQxUYBEP0oOrE0vN+pUMG7xKt8VIFsILySvX62mUzrfnTW/JpMENb/SvS
IexFgKtymgpnc3haOwHoWKv2KyEK7yERdIr3p9Je3k3pRGg8VUXkrMzx2C7g
8+ko49SduFn+7GOgPBgP3SXyUSIkg00Q0q7N9MJMpL3MKVmtVmJ9JFZ3mpdN
cR9kwfvEDutkRAyVCIFPCLoeghR1oMnU1uemRDWsTCkpk+g3sxz8KeyLFKWJ
pWvxeT39xl3x1/T/t4BlAPnLQMIzXi/qaI2UtWZUIClStSsDUnlH9H58Vg8z
j/NRTgF3k0iHWmZB7ZkWCCBuoZQHO03dBOhhsmS5503YYOjTuHBf1N76I5CP
FFGNCFyj14o9JvteKVRKClwcbx3s4AxMMbkjzqr1hpfe4u+K5IXrO3tdEWBS
J2cqIHJ85rZ9kOEqnOVeqcqx2U35Dr9cPlE9Q5VuGc/lEgWATmJjj4Knk6wT
jePXkQWhjBY5eY1QmoM36Naw7BNUts2GCYetF4isfeNsc+9Go327YUvwxZ0c
Bi05WjLGvlFrN3HAc543/Ma9xTcph+A7K5i6RVFor5ByQ3/ObNvf8A/dTuk2
MFVtYglKcTfuFxJ/S1vm2+4XtvHHi8WtQozFZNWg6Dxw08KIwVcy7hKgdleT
XeqWL83+J/NZor4sJz4642BvvLcQzfnSxamAvI0qAOB/aSNlxm3qv3EdNmaJ
NzRZ5tG8tyIrhM+rAHcgNy5G85Tn+9oijpSlr6immyrBM3wY4kLL94QyYKPE
4fNxPPQ/uWBUc2U9rHhCDHnOIMN9WHQg0ueVLXRooYsMkrUHGoucB5Jlfu1J
sPfhOTjz/HbaBRuvCABThQ0yN3M4MqEI/MpJ/QPOMDCBij7J4C0Y0eAtOb7R
pio68eiAge/etgDQewoI/SeUb5Sa7eOn3q+CqYp3P2b1xp3BnJg3BGuehI+6
fQwFOCqfxqJhFoJl8P1hO1mM+s1zxApiCdC9wsYv5S1uemXfI6MuQS5Cyzho
Gu9qf6b3VZ0wnrazbIv9PApt58KoXs2OjaWm9D7jdc/Xm463oGqnrB8B2g0y
Xd4qrhAeH4A76EZgEyn0AR0CFHEhQEJYTcaUpUViLzEFHbcP2H9+Mc33HLJx
p+AH8TIhcuL5GtJIg0mH4STA88IFKCjLQqxLIxJAq8hizuFrB9AxScIdB8tp
oiQZ8h31foMRJgqIwKgtelHRK1fG+QII8kgbi+GTz3bTbb0nvGT6oLnYg+W3
CndmEGpEOj3WlnW+0GS2LLEp3OE/Q7kzzlEWclavSDjWvf7mijtm9XH45Luo
TeplEn/dRsfloogHbpijIpNbtjxJyh5hEbV+/Uw2RALwIaIME9hVPxiRT8yj
eVbT7gGnLRcve/mVLUyu+gfIsTe9GbIetiZLbyeLYsDZTlAOkKM9+ynvMq4Z
j+D3gAvXxEVYyEZlVEizHWpDnTsXF/0+Z+nuTSubzgt9Jramr55rff8Na/3o
OFCh/phyW3SKdwSMcGhiNzW3UFyytRvtbmmfAnURk0o04o7yIXRclIxG7oJx
abj+3bgcoQWHN2PR8Z/4XX6W104CFqqbLabexudqi9GFaL7vVmbQZGTNsdgo
G2Gvu/btgqvQ7ZMd7pVqpBbT+r+2gJuX7tV16DBojkJzZlHXLknYXn+PcXbz
mNNvfj16TWiaE0B7GYwhB56fZLON9/ALlUUsaZW02Bp5MWF+Ij25GoqGFjhJ
01Apg7c9zPAImWR6+B9aWaMe/97MzOAQCPiRu9IdRXNpxHs2VVR8h9nly2FU
AD4WzMECGWyl20JZUa6lck+UNQHb4mJqWBUODtqb1rXGBOhwSm6nZkHVRLK5
7DmBrg//kGQ/SrNM2PoIEYndVtI2imbknv3DxGspQgn6O9IF1BIYNkMs/kRi
/M26uM1hbuPt/U8TwtQ08ixZ7UipDjaTCxOGJK0U0IljQ5TEpLFz8nV4H7fd
mlcw2oOTxyluAf8wH7ypdvRreWUhIiMMDbjQ86+lKc5WIEkQc7dirJLfNtvg
FcXDlF3mAr+GJMoPwBWMDjum3wAoz+etsfL6CHNyDNTfIWk87d8lUaWAQ0LJ
CMk2z3TOEHwZj9T5Qfm/FNw8lxvZXw569YFYrwyae6UM++5M08t6hKpjZSUA
X9h+SeRK4wD3RhiQxGqy9pYQsgqkpG8BHFBJsY+PgrkiO77GmNt3xnVX5ATq
p8RzfNiM/dTE+GknwhppxPaXuaawQV+HAY4ZFBm1aDZkqeuSxn5L9K3UhRmv
76E2DHWYg4Z5pimrpby0QtzPmllzQgFX9xxyjz5fKQclcT6/YQjA/siHGQr8
afx/sIatH9ti4oBJbV80kvz6gdo5F/O9ejhkA4zkyCCFmBkc0uJRvdve6MZP
k41rCs4WRjoO16YhPbT9cIBO3RBYOuSG/iaAri3OSB/o88ABC+adW5Z7p1ud
7oAul7KId1rYbFT/30MYEAiSluY6P06lSzMOGlQzkWHApG9WfgOH07Nwt7xy
zDJyIJDKx/tAG1L5FzA7K+DJ+IBdpq/ksWS/nlOXChzomZZk57ziBOvYsTIR
aq5BgVyD2jRtVeEzctLTv+9+ykipuKqryKyIA5fQNq6tyc8N/5XhO0E1PCSl
V1nee7tpt3LdKyawPXaDv9t0y06Dxq0/xhEIF6AgJyHnzukGcLtASe3w34tO
6Mg7HWjVCLnF8t6n8Wi3iVPCR8bsaaa3NXivZ7eb9G2XjvcaHc+ybFQr819Y
Ri4WyB87v2MG0imJjrRQs2tMmR769t/EozYxl7WtNeN29d7gN+EwIqRyQSts
VH5JbRizIJsusm/mA/pcSN+lbC/iSdLjOpmszcP/Qc+fByQ3cRj08q7Tgzw7
jr9JLqzHZdnacjYThspBP4YQ7qAbgBHzwgCneQAhS+FxeHhUhymSJHsm99/y
1TNnu7hMP4G0//Jb3YBaFKy1QHQ701HjXvUaKN5M848XsNN6+k5fE9R/w0TO
oecQHlcrfMO1enl3p+ejl1xlUWHCRYCZwGFdvFkqY8lZkZwwZBm/IX6n/sOz
yWXwRjx4+9gMTPmrsH/7FncCO3sokOfNElvN4gLagCpOsCe2smII2CIKbPh3
ANGFDmhZlWILTuzjxqf+cNgVVb0hyZC8hbuMzd/brcRsaDtbjx7nMAbXvyzh
Pg29Oqd02lrj+pzZqs4zN6sEVqRYJ8p6SrT4932L1wgc0VOq8U+fHuAoS8cN
Vrc8YJuBn5BvLH6ZZuM/aSfJi/IsGQtp1eQOEZMY+XgL6oOV4BdtEhbvZ+V7
voe1BJc2sQG5nIq1eooXDayrzvPp9lrEyS3gC2hfkJ8Ey8FG0kuCGrMw2w8I
RNAgN/2JQYYqhtDgwiPp7PSjb5z3AlMVffhP0LI+RG9ajsyeIXEXzDuzYD22
DR4Toqmd32QWyD91slX7aOa86wO3LVnxlzwOxOxbs7up+h9+WGfnMPzMNsQR
PU6i3ZCAYd0oph+p9ECAfUjckVzTPhim5u7607A9VKIG78c+StX5RWDOOIJs
5kjcQ73RMmylNAdxVjNvJEUxm3os6ADC+UwYPYITGyRu8v8GOmAi1021axss
TSmS9i4aR8sbBxVLNS/dxMzCMunBRhXuXb4DE9DbaMjiKX3JbfLddWotKF4n
4LsfETAS8CRwE0Sucrogpibcvjfgy4Z5/V/vACgohz6Aul9/p6T6DYMot0Il
CAQR+IfxNAKtzBkcLK+mbePzEnM08I16+0J9MotBMaNW/T7Ip69N0LzLibkg
yofMJMAA1t2Ha6KV8mH8/EWHiy7PeEiz7j8IIxGpmuwnGBZPqBh8D52B/C11
ktXN18mXC83qPpXfUZWIter1VygEjkdFRqakyFcpirCsW1zjIRByZ863DzTA
3dXQFZRg/n3IgRo5gQNcNKGEp5BG/DmOAgio6UGRxl9C3SJ/UgPm4tsMQPku
xYt1JBCWpYvzE2ZmZpf749R7C/lIl7V4fAX3KDkJpG2rMwzdQ+Xi7Ovwh55j
0I4rE3I0GkijpWnPBBu9L4JcWKD/dolTuJPMdv4qwIJgYbXR1wwQ71m5uYqw
qgZhkAuQt17xUgUwV75MF4CafYo5F8D1ICRcHLXfmrTHdtXtCe2OoRo8wmZn
cDmNNsJpHY+sh4FP4RQPv9uOLWhAJhVybIZFQjkNJwoIe44/RL0fTbzp+RTX
rI/8iaMbrq8ws6qGfaDUd5wbcmtAngipUPfSY+WIoz3IvDV5HJqpb5mGH/Hk
/llyr0bI8Uvle06Cradd4ScJPQhcFO/8sj3UkyoD599RxhAfN3udHEoC/pFy
5rbYmnsTtptBD5bCiIPN7EEWpUpgeiFVFeZsSwpjKs+cDRJvqHRDnUSiz/of
Fo0d9xMlmF5CkHCbcLUM6e762eXy3KQYi6PHmNjzapsglCnwfJgh7hKnfSqE
4c0yTfMqXN9i6XEPucC+8IQJLoAv9BunM3Lh5JBO4O7HAie83IA9ADH7eTL0
Dvk9LuaN1aK2IJIrEOOZAG2hPaHBu7iDw9cW6QhG1zdlnHrpCebsVBgl9jx+
YJYcECqtB59I40KxysBcuQIklmd/PcHXcuyBPRC7gOYKFU4Aq+2c6JzIKSUT
964mpdGoIb655CNBm5LJ9W0stASxISwF/NDxjLIAkepYCwEIe94CYUS0HTr5
GVSOp+YtF31XnAAY9yh5zB4N8r78dDSpIh2wOG9el2i7kybVM/3a6hh8mGeY
IgXXHCmNnHx+PhigyFOA2jx7egqoklTUDEXHSTMs3ibf4Ci3FQyKigGLPV/C
mvvIrk2IBtwAkDk8Y19Ca/QttltGtaGtdekTt/MsUM4xB9Q8bBumxsOf5tJO
+de81aKMinazwt+ApIDKyMseQcHXciP1K72uOCMhkXc50MKaX6YZf0HGLdp4
nIx77KAXEOqLtb0ywh18Oi+P8v0FwQjOSB5qqGLbXmK4lP6gCZ7N/N4/e0Lq
qYixKEVFFeT1iz/dGUcOpwUEVI84MP8n7Mkoqd3CJRaseKtFj0W+KhGND5uv
r2ZQva0STGcjm9cxVQfrcvlGc8laMWd6mNlHBEJhlEa+SAVinJ8xq3I9Hmka
EhaSV3A3jzptLPsHpqFIRogcIQBz2vx8GdFlgz1miumVEjhxN3pquNi9IxLH
5thK6TU2DdrA9biDAcB6tQP0g2r1zzzD+llqVyI29oTYSoHPpafiBwlWr5yg
qbxYjMJRPEopRVDsnLsoJJRQSH7cb1nIowF+DFKUnopeNktR4il+33Y2D8jv
Z4JgOli9brTv23yieYqf9lIddV/S6/WfwI1W/2Nkumlkgd0Ul99ppeDFlaVn
llkKSbhTXkvGxik2Y+a7Z6zxkplGx/JPcjhp78aonIHCjt/CSUyHpixW1yFR
xo4r5N0/CfAewiPp6n2b+4F3Ys+XCl9vRvcPPaR9Sbob44Hhi4jXHA62NXmu
wcFAvG4x3jnZMYMLjKt2jRwd3QQ7wqPQCXdI1LHu1aEf0F4rXIn2a0wMHIBJ
oNp3A5THpiB2j1IMoY0KS/zw+HpXNEXMThLd9ram9O/h7Fx6yt6Js8g6Tpn7
DJgbpOz15i0hiZn5R3RyCQACD26+EqHLfSuKpMo7BpGem44ST11KL3Tdf6Qu
okiiS9fh43pgfVqCvjcWglb0ZLU4CwxElXTLpa4XTCNXEtC3O/62Zq14ftmY
TEoRJow+OdlxqLcpAkYuS1BgHtf5u6clOCQxMPAvWJtGZuGJIK9ANnnl7Lyx
OYn0rnRl0+TdwOW8CzEuZapOnFvNz/CWrbMcGwxAkgAIRhbiGh0Bktdx2nBA
WVvB5FBQJXY5lCm/Tr1LohDnpMfafoQLRcd3V3WdFdklVTv1YXALUSmh4D+0
d0zzIlikBXw5UFv1spmj0Tpwfn5rE3sAf0EmvGHUfNns7wyAnkyJ2UPbH4FG
I4pU2zA7nonxfIghM+A4V1bhl9T7Km/VTsJ4LQkQYhYPkje+edTCv60CeLwq
LjPGJBC47S82Zkl/x2WLZMP1OTP4OHAsfDp8848k0gX2F3WeO6npLGCGD5+4
XJRPfd7XEoeyOlCwuIvELIOZQbTUpru3+6oDKHomR03mmEj809zgXP+ZJSdy
MKJRb235fOQ05wlfv5HU7dny+5jWs8fTCuDwlGdBlRNqqxjAb7SeLP+UChr8
ehcXh0z+HbCvwV5GP+fJd36hQsHbnDbh0C0EEIzmpalkoDhx1bccMVIcVgWQ
9iMfqd3KcNEqRAfhHTQuu/4ZdBMURlocWerJ2457/rY97yF+Tpw+xK2Pc8nd
Ir+L3MBPjdOQcvNPrw31a8I3Rfti4yXCp5RhoTmv2QnRGYb7fsQQtoNFIKXd
PEfH5b4qX7QRvp66s6yAVbgb/BpCmwfdYk5Ssz7fqddDXIQ15SRIn1bsHvJx
y+kOlZRq6khLdJ8mvs9q4mF1nWi1KJheLteoPeBUpMKk3fIa3ksURGO1yFFg
0AanznliJ00fLBDikMSFkKx0vncKUsOqluBYkoUt0QUGHYnFDv1/pykUhIg9
SIO2XoViUzbiuVB/CAsOTTbzd8CeRJBVqVwof1iB5/zU/QcHTwsVazGw6YPT
bYKSX6OwYVvNXQAAczZGrSTiyKdtr1c/pPLOVGRHQzCS9Nj3C00FDnc9AbOv
XAFW6T/NMzJcaGl4hZTTotpQpZyELXJVe2hHItTevxjwY9rPUu924HswsGaJ
6KkeAvzK/yDfL4ZiCueSCuMlAVzP+AssUk+iA4hM2xxdlVqLTI1XnCZCu3yI
9WX1YAbHlLDaU0ck4PB/temrpmop/tPZ2ioNpP4AxaAGssKKyBVXH0uS9CPm
38be8jWb3N4Nbjr6o6HGRdDK0AnWQFdG/19Ko0MBzV+L0v07D6Wguhh1fHAD
59gBnZ9CXOwn9UjRUkzK+jHsDcViJjBhokvKm+aDCpTauPjb0IO+ZqZyGYGy
5uoUn7VIbI3nLQbNw5TTAqLiTFgWALmNZjkS37dQSy5jqGm41A8X9gnGfGq7
UflUiOUbv4gl02xcAo/VEqu5duneM+EWwlc3Zd7rVjfKD98Za7TeID76QwEu
NGUedjufx0U+uHdLeGDYXsuNJ7lNmRYPOYYoUmnP9SogpsfTgIEjSYOmAuF1
SjTjgBc2HXlqw4C2qIsaWAQYSSi/IxXQOXXJEn7wEeDx9DBZtNa9/aRzKxpY
0h37dV7E38J57MXWbo5wHlgrXVZBleRxX+qdsw+9LgsvOgHHcXaWoSnmsTo/
31Pl8MFuhGjWmfqJPoAlgFL6jaTWPa1PMIOdDMiyH950BDTZk6vRaPscfKXz
/lTiyIUxw/K8P3NDbUKHbZtTbwHx/mjIMUh43ASVr4x+fvvCXGJTlWggwgoD
bp06HEkv0x2ojrZzkZL06L/MunyscjQiDn8QpkQrgJbVEQJ/U44TzW/6rz79
VWkkryvSjopOAxQQ5QE30F3mShPec9tpBxtNWlP0KHpQIybYMDoNJEASAd29
XK8A9LEP/OJ0/BsyrgIcTqhxxV6eYDjVeaoOCwLV89L66bWCpYcoMM31r/7f
xQxetLmRE0XhfUwGpOaY7I5vVhs5F2SJ2/BMA5vLZdDF3iwbv57PTli5WYMr
J+9DoRjb14NhI0M1tQKANbP0ULOxtnlHn+1vlMP4iEOiHLGDyKgTCI+ZhQHe
eotSn2YqlFHmC/rjH5bjxya32aQlejLmBuSH1VFfO08Y/sJqtv+1dTMyMhFS
FgjOhUq7mG65nzGo7xkEsVcvMxPpmf7SPejM1v9t5Zl1ZWAoKX9datM3Dpif
lNdZ98+m35+xnFnz6JkknLAcY9tGjow2q3iWq/Pv7szG5lsJ7Vy9tnWcjfio
LcspHV/VVpkowX1oRZzqJJMXxiV6EXNCVNr1jphinkPAbyMsps6rx5q+r1cn
PGO3riQvKEGDl5lHc8xB4F7lzu5QQsIfz2TV5Ti3g4ZR2MNNW+vFdtmYfSSF
1KtOG6+dHcSEVJDmspl5bOMnh5q+evZmoumYKAB2VNMChu3zeU+ScaZbapHR
/wqzfGMgbj+k4iqY7xbWUq1bLclSl7oOHz5QRVC4hK4EJlxUKcKFqjDKTrIU
rG5wxO4NZhHjtQsk9fBsNvz26eRP+zYbfagWZANyPOXnfQP7CeBj183Oq+qB
bImGqpdg6ox7RV2q4ZtVjAKaF52vyl8csno4xxfOvmqrRFaSAkY+S6479Xc1
qp8PrqZ8E6pLxQ2dUfEH2ZehUyj3VknWq5FgqNwdfc4Cs3W/NbusYMIrEHI1
EEF7RWx6SP5cN3ZhTOBou39O/AkbIWs2FPMrMF6jfC5I5nSq/IolhqZb0BDL
NEsVFcc9TozVcB4yE56mA4eP4rEZyER4T0bkauFtqXIPr6bhANHT/BNPHLJz
MqM0O1Ccr901+fXdjt5TJRozy/Bn3us5kySXKNwJ+KN1Olt1HYqFyzsFuqY/
5pu0NCz5D+qIlz/4gAQ1AsSJ+hVBSQ7XkXfBWsrnsHDzlgK0OvrQrxF2e76i
1jBTTYCzq2Z/afwabNBIPDgvyxiyrpYVsB2xqSDOCAbgCO2vNV+PW6ZCCUYm
E0lQxNICC5SK+4a7dnA81DglrPDYr3g3ueQm+r4b8OHXPLPTFBYzbWFSxZcM
ZQ9aIs/aHXJye2V2XrkyUnoNfLJvKQcE20r06RXkLuCbt/Mhfi0T/XmIVqYh
Lq2A2AtWkNfQMXqQVEN6syZUusU4lggwE3PHOJhWSAhydojPDQGY+U/DJDHB
VOXf/yYFJ4/70X2fldmCeY0K4PMtdJ6daBVfBfDQ0wd9ruf8qiNTLAk9m9S8
JLXb19BHgEDaYBYXJHen59j7MWyb6TVYUP8jcW62tHcalspbYADKPo8pCTNk
s6EBkg8YWufD/O7ULfIM0R9XUW7hFKVwyoQ2dHoEZ3/eTgR21aManP188g4/
JunldUpOpq5oEHLgOdipTgW1lG4aR59DbQJP/h+DD/r0H+VsdxUrJEwySm0o
y0F7HDV6m+XNY+2bOovB+n/EYZ49EFExIA41xc8YlTHFrClIsfFtCknLJeF3
j7yTFW0HRSC/0gcMeu3B+ksTkqXbB33oC9EcCkL6MgqsYzFRDY9aTfx5sQe1
5RTsCO9nL0ZDE+JZxlVbK4ts68lQ/boeRoM9xxcZlEQjiP1c4Gpi5yOLt14X
4cjjVMAFxaZtNgBw8ozx2vxArzGA6C7L1mDgsC4QYBEbSbS6Nzz+kPMup45N
KkD7UrwbnmRUJ5tk5dn+vfFJgu3vvVnwPY3zaq2Nu+kZ7xXQLLm5LvvpDwym
zWfrwCEPkROtVG6TAwQR1i0g1LFA22tSnLFlPxIqR9CIMw0YHQgpCMTaSA8A
seKhs/XrKmwK5v02xO4Wt7QTXDMqMMS7Iov+X8KMWkYU17Bt+eIcgDXMIVh7
i//xGPevRVNiXKJ1IZRv3t+yEgCImnwXt8loce5ufkKz9qSVQGMtfDP9Hze8
qbam9A092hIl3cx0i7LAOvs19zD5qLMnlGElKXkivyFaYVgTXKWRhG+vJUrT
Vja4mYPEaCjptxbd/xYwOrd4It0a25G9A+bJNTw0tAiGJtU6QVwpjNqszWut
MAmQN+U0nuN42SPtSMgN3X9yBNInOTqtevxe5qlUMoSIX9WRKhDy1dWMd6Sd
D5+bKPUSb8qMumwLTzG/ezVf7IqC4jhyN7zP4gBoGt1I/BpSJhEW9xAL4RFf
O9vauaQeFkwncfHme3aDCTKGxdbUfyt7OSmQVuTghNuuJWC8qB/CXLpEw7Xe
4j+sJWTQJDBIBoKgMiPG0e2T+SAax27nWMMy1Ojf55Bl3ySP3gXPWmJHfp8s
8calmHnn6ReyEp5RVlRgywOcgasRYepcygJY8GaDwZX9WJ5IPHE+mA7tr5RX
h2qR03erJ2pLmYUr6C8fb3B8DDhFrMUTOahnJqX4BSf+d6r4wVkjk2rgeA88
llWFscAhyGWQY99BNBzha3DErgOMA9LHmUDQ+LrZ7txuUnUdR8XTpX4A3hhl
Bo4olTP16YsfrsFc2B0/wz08IB9t51faPqmmSoXp3tszDzHu2qhDk+GpSxiV
IXH6Rz/nnqc3MO1nA2EJ5aQKgQdyS5OISgJgRq6kxyVS2zKVURU7ULr+EN+J
zVyMJOFmUtD5pljP75Guj3oFXpezOHn/rFsGrsV0HcsKCIDZzxS9Qu7/h92q
VH1hAbi58gKzoG6Iv67ZINMIgEhBVwYpJSdsvieLK9NV1itYRZ5+MOEPPm3K
qFdHLHEkXAJNTp7QPi2heP0R/vo79gwRQVTeGnfmXbIjGKUtUONTpRvYYUNX
a7Rcv9/0trmqtuFa35pe7+WI9heVgnpiCPQ7LBzloirCuoR1KulguyKSdHTL
NnY8zmGe+fVdB5ztJ0+nQmWYOIptMJTgTqD1Jaz/RnCm6M0uxiG/1JL7XJi9
yNVomVl5bfPvQAbw5MRTC8Hn15UR8ntsghL4OrJolN0qeHxkZJULhRiIq2u/
9W8Cw/4+sDEXx+dCgsp+/H9rx/i7Aa0Iajwt1pLevAsTuulnvyucnkcb2KV/
Tx6TQx/3yh/NWfg9qykKhR922jNFGqqjcIkqKiAmlg+g9vQXRSC0Fh78rRJ1
zN27LaoXQbBXs0m8DmvzvDskrxwEitQMvBYLj7xIxMn9YdJUCQ1ReU6gv2H6
IcEaU1wHMVt5TTQ1U4QMlwB0ZPIHdjcIr+4TsPGTS8U8MC05J7JILs1DIEgc
m52b/z5PjCmBdRFMsL3TWsMhOPr7xQ04g5LMuyh0/8KzNkhg9SeZgMf7DX4U
n+b6f5V15shRSkdGsXx799cQ8QbiSw2m86VdDIr+bvBR/9aF+ZwYdSZM59io
jJ7w9Hoy4OfJp9RSCcBXL23bMb+OiFuWm3Ybsn+H9+JjkRX7m2fkAPHYoQjc
yYyNlQdqEBbyIJmQDjDSfLe8D+ttEIn9gKsu8/JmcXvMGquQ8yyudgvsmFEt
0kEE9aHF3R/iWF28p2SIaZGdolF5MTHxvZRbTjSMlimxEyGZdqFEEIJ64fu9
9sPM/inrj2lB8R0Tu8L2Dq6NYlOvbAPuHyi/4pB81+wbDD8+FbHVrmo25anG
hYTFo2hNuw2TchwYSkBXHktkAwcEQykDHWhyRohgbwN/wMOdJgB9+AUhXIax
kGedURaD4kkZPY4GdZQrsPi6XCp3DR2/jLW5Ng5pOiXO6DxLNgQzINHLACnS
PYS9KbhhezWi/UEiomLZHULTpvGpMF8ese8C6RG1SCd/x57bS+0v/lXBrit+
1opjisKgSJWcQ+ipq9gRC3yONJN4Rs0MJetJcZN2AYyUl+tO8T4xRc4m6nct
XsfWYWcUVxFsE+V88Stz0BPnxkBjugrW0KTFxOC6eXHHoB5BDxprZje3o14K
nwK5QSa6ZLa/QV5N3uGdicM0YQkstYoQeMUTIUdl8NN9nhP5vtleH0Ym+AnQ
TZ0m0iWvFRd/nwHJmumJsBy6nGVUD91+F48nQvKQeVb9bCae1Oa/XGPT281U
Vp0d0TIRoYaUsG43V8Yvz6qjbwAdHNI4rH5DjHVeJbWnpof3klpyn2nJckAF
8YQPgsBkwxyokEnWj4o96Xny/p5NRpzjm9Z+5UBzOScc+4+Ay4GDAKuHFb11
M795ubyDtL265hf4v6slJqX+Pz0hUhQZNC3DKBJs6FnyuHpVE8zzS5QjrZuy
4l1ZFGmVqSAJi+hn1PkLuepUrzdptGnwr9cigYhw/Q/T+xlLzUlUfLqWIrH9
9TMiS6Gz4j1GwVOcAqaiVAtzCep98ShhVMKjpXB6pAdJTHyasdF/FsKTnOPe
GxOFafeu8T66yHX4dAowwllzsyU1hodIg31wBc78jzgWO4xJBH8UmOaklcpT
K+K3QLKtQ+InobCCSD285zAkk21LjycBbqnFZdskMVwV/NKzl0FQKBT52281
rNOpbPHRp6v+RI6R/EimrmCo3qGkHx63Y3IbDZdQ7vc90rTeuW5eBOIY8qkG
C9sW8jvYqDp6IfNCWR8m2nMHGXB2hKW12bmg+aBEtsIs/TJTtiliFH2q/g7Q
a00zVnG+xifO9lVTrAQ7kcFWsf1TPeh3A8tdBxmpuXvjQ6AsLezfr4rUrIu5
ogHHz8TDEComHyfAM1TVIN83/G4yhdxNKM9yqyAKsRclEmIZPImyidT+66YN
+hfUEO8GYnU2EgMK6AMKuR8y2geIa2xCEVBBWidHUaPjpWHg3cBtdzXzF3EF
Fvbk+ez4mocfWwxZTSZg2aMZHY+rlxlf8ZX/OPBqlf753FByu068Aaeanl0P
Hu/Ge34/0+vvwXuxlvBORccSYL/y5A8C+AlklN6zszre8IVWRDFfQUTXuMl6
+TaYIEzDj6CF19Ssxfdn6p2lcMqg1sKPJzDrjweGsGG2EMMmaR993i1riwO9
CcjD99kUOV8YkYNY3KDe0sH1ZV+Kz6/EZ5X8WDQe1jWwCAXLz6EMzyxg2qUA
hRiGwtaiCQsjIvb7+umjFdaWKqo+anrmtwqOcomy1clLQPx92vDejPWTIk+1
oDx5iVBiTePD/i387+JLddGEN02d6odqToWd+MOqqhY6EtgwTzwKLKgszbz3
GxPq0EpB+9JlOxX859wZcIDyG6Z+ebPtvq4ZYP+UC0lXTRLQs5rCfbH7z3od
LG5H0rx5L7cBiBRhm/gzjuqUqNLjxkr5X24ZIXi6o/cFAbzci/8WVurNQgQZ
vdrUMiqKitHYeH5LDX7k4AoqXScQRMVXvrf7/6XC0Gr7JTyeadS1TfmB1km1
Y87EBzOgU2rf7CoIZvbIaRXyMv6joZUwUD9v7eW8cJr1XkDg3SjSzp0KGLFa
m/sZszGCmyMibVCSnekGSDZAjXfuZ3DQS63n+w1ivYGfN9RcWahBtgR2xXeB
qzS9kwsYvIjwWtArXcakLkBnZnNMoLiRAPUH5uT5epxypC9onIrqxdKELWVG
2zqg2AzETllQVnh2xtCaMYPrrLHGJDSg39oCLNfRBTmOCfrNtml9w1jUd4Nf
veIp14B0Rlbp10GsflnDJ5P2BD1ExIeaWnvop9Wqb7Z+BPgZcypGYfiVnafS
8qx9MR1DgvKpWp7tnRlUoRXTRKVjbQhLGLS3ZDIaUj1iUxyV6eZ7C4sEoKxX
6FOJwPCRv8oECe8hEF5SUK2GnAmmhUin+xUlWciBXvekjVP+/KOj0fl6T6Ra
U4ryV/ZwjhPsQQx/OSHGmeSZI8oGdOjnvVzWhU3LOGDSb+l5XKK8sob9yBBU
wwd4avlvCoAcsYCS1PIep2EHddNbZ/64hHUW8xg6Pa+o1G1GTbSCohDO2iix
HjrhfEB7jiqUfZDcPV73hexwHBsF8P+iC8ClPD7dlCM6Gx998CQV/4yrQ7zR
LzfoNRc4TSl4Oe8xcf+JWoC3Y6SKn4MGpUCHdNWJH5M+sMNTM0IJqfYQVN/n
V5Z+dNBJW6YcSVBQ0lIHbBnY6rS03HQG1VaPv7jlWz1Du0XiotgqGH23xVcY
PaPg85LpJObGm3M64rop+zswXOLWvGN1U3qaU7lWnXhOqNfvU8uMzriOMakM
oM7GiVfYmwtYn/SesS5/A/M56WrZOXnfh8j/F8ARiWsw25btLohp/tPrmuMu
Krh++4Mz3RUobh5yM2mBWHQlu/D72EJenSRxDzqzgEWzIuLhqvzCOfuHZDvH
yeQlqk7yCbJkTyBMqNXoIkJEW4F86V0HVTIHDKl8HllMKHQe5BhtIcvDCMoL
Bx+pwRCwDseHVCnisguQwZnbTOJx9qIS698lh6pUbf99L+6mJY8wiQOIdSFK
Fhf7IgqBquj5afQtGnTrYrNMURKOEfGEbg3btNwRW7k/ifG+Ml7Q7kfxe944
DRXMNtTMesdHJGsdXDjWAvBuF8toOxIqYXTo8YsrV6shjn95Rtbb6pF4qcDN
WJ/coKq0xdQcY1FXVGWTN2QxVBaPgixadHPmBPfk0Wozxzn/NJgiz/sKeHZL
1YYs606jJyPjXzRKAUENiQ0m+nfhhOXHDXi9323Ek1hsKzk6OwOqCf+uXZe4
fQTrrQSw38wn2mqueNaH3Y/r7dLZdfR6nvjaYjTpgomXPvPv3cxefzDKElWB
VqtEVwVcsf5kLvBCdVYPFUgvQqXUUioK5w9M5FUlcSitoISFFHSipIaKwM4u
OtEA0KWYpBfumcACNgC4jq/oLuiV1JtwDPD6rlVeIjOD6dZ862FXRjUhvw1a
ZgGIfmIhJGEcAkvMtERz//8qhFkuC1Qxv27N9/f9nEYopHNygmR1ENpKXxxA
lXuTiisUjy5M/lruRZmz0t7CQ2f4moHYbqhChXA3F5c+ThFyC6ciqureEHYF
tm52yuJz+rbzNJW1mihiftRsvH7GAwBOhZKwNNw1PMNF6VRMxlS18yl+qxfU
Jfh3dvSEYznDENbZdbP8KROMvbwHYh+ZS/FWz1CJm8n6+rZ8WeFAoDxZ+KDW
ZumDryeKIyuJfVdDOJAO8k+i1pMP/xt3Az3nurkdWTNWwk1fqRdi+2qaVaJk
66dqhSDDOh2HG6ME8OGnToQUckk8aiAi/1UFEofiQb+dKO6c6Gzp+gKjfvTa
8CEglcKBzCgyIjtT8yAA1Vjqm7/QMg85LqaI47Buvg/T6qv5Y1JHPplqhyo2
8KhE6DUhnu0SBjCFNLsfxCRkdHWsVW/LyituJLn6vmf4KrP0rxDQ1+FiS76m
2cB3NjR9+FFz5DazUEF7dqRJ5RIwhIfgAN5Pd7SRCaUo/7KZBihI4YsdwYvd
7o6Sx9XTiQB8HLqB+uI2pqq1CzBj2GupQmQa2xmbkKwzGxvbMXHcmJjcuzQZ
uqahZSmTpjqv4E/GHCRQMiTVTgmb2WaTfzyoN8rYABRvyP2f2KdM7wk175S0
0YWnVty8qvF4pu8oM/VyGaMyFJIxNgTIdrKBx2co15B0f9LWvS5UbdaZsfm4
Kgkd1J1BT1SKx2uqC9Pb650W5U54nP2Dm01GjctkG2bb8MYGaqBVt2OA7p/d
yVTkt1sulvlU5zUtw+3o1arpGThytTmUyxiWKRUcvDyDij7kWeKbR4rrCl0d
pjfpah42uFnoCMqaRljYJlrEgwlyK3tjSjwJqTH+mR033e9YBveab5wxdCPA
SbccVuouSwVebnWv5YO1+KO3/ZvoROce2+pY2/mmdDqlJ/wFFJm1TKaC204z
G+t1kOjdPXg2Jf+DZJjWKHuAjAYx8YuPE7AGbVidi5ZU0ufBU4+ry4nn98X+
3bgV13wzdGAADMpdhnjbbEy8cVcWMqWzN9ZHZt7D+LFWnltHq5cLBPKSjSTs
Nn9tnoYYgdiL6pjDNO8p+dg6HDmrV1r+VkJX3Wj3lDnE4F6O7X5xNOL15t3b
8V72HxAL9cjCVwQh+WLRX8V9N4qWobLbPR2etWGdhumkhhaXaRLxunfaVRu/
BenJPDXxbRUtfApwLLfLRY2ikp4NIOGW8luYNdtOyFEVsSoT9ySm1+2rBdNl
aDFWiISbU2jQN6PnoCtRoJiBg5FeWkBl6BF0M5aktzbQDduZ0oTilOArSank
d7w6OUHbyiMiTGqoutkeISzckRbpRwRiakA9FcxzNAvqo3yh9MOFpNrNRCkt
mcPYpM8jh3kET56MWblOvK2mWZFzst2Tqs0YVQq47R0exmb/PGxgb0imNzmG
0nZ0tMK7aliDZZC3/seEOVbiT3EIGpBDA3mZrfya2tMwtwDGfJ+isp0Yg9QC
RHTcJDD1m5/N6U2QimwQhwEXkkLFI2InF/USfksw/suEPC/j4IxxfpAckx5F
S74NF0rxSZ34uLPhpN5s0g6BQ9laNOCewsnqLeFqJg7yIWwD1guBQwWGnss/
lRBip/ixNRrQrzLfO+IWNELfuOduNjDbnoCpq0ky3nsEekVKtli23Wdpj8qn
TR7CH1Y64abLU2ls9apogjzs2RN5aPoNqk3dE4hvsDUvZzo4uhQJBAg1Z7+s
GNKIiaJ9RwnuModT1rNoZzoR2tJZqu/O1Sy4lIUYPagTkWhO4fC7JMC79KCp
LlhiZ6e+u4sWa3ZhB/qWYizRod8vzXIpGtrNll/FFDwbjKoieQjjH2xopEYW
pqET5agUEQY/U5Vb9p58pxoIZj9ZiCLmyHh4HsAxebsLChMYL+WnmMjQB811
EbxTIBEvwU6eGr8WAcI+63wkQl4AfIPKruZ+x27UI01oUt/mZTyrd3CRrIKP
NJBky/7Fy+FOUao62RlPRmAqtu6mP5sc1ojph8k54vW2vZ1yPXv5CNhWYwtN
sVOgVIvAIe6UUko6vWl9zNmceuO3WvlRc+gHxIx6w17Nq4E2/rLuhugK/mVK
An6V/SPZ1faDtXor2uTq8Uxxjdqhz/AWRXX3fP2yr0FyWRHMynIAPNA643o4
XqzKY+p+AcaiVGUEsGwIEIKCYrTE5s0IQlKA2TQx5TV46OEs6qJQa81UDpCF
bvn+F/ueUAFoaoOaIDSMNUsyI4Hbb5DRd3gPTVfb/EbNu57ZoERJ/Xb45ltC
VfrvDnrRz05qRgEfAN9ak2fNml6QK7fe6owiytrY7JhyeDFzrC5/YP+5DpKL
Q0aA4WnjGhXlJHtNSAJ5RV99c68yXICA2JXxuXhpqcl+i5oDqF4eH3nah+jy
V3l68cdYoTCkxDLLflkeIMI8LFqsN6ZT+HfY7MBUsaNsJAEgDt+6h7gY8jBU
JTOkwTvfOPvn2pOB9TpaKCeJdyDyDyW2smaHMMh9LOWVyXLr9/+Xk2lmKRlU
q9Ja+ZQan2QKc++Fj2A6kQ1/pe10dq/RFl9oluLEjENrbomGCAMiskkmfsQM
m+/2i8yOl8VEScoflTuyaLVxfLRBJLKFouIRgq8nTa+FDwLZR8ObduFOZ1da
+fnnR1626XvPvSnL6yHHsB7ZD2TOmag24gM0iU6Lsd4EPGKaxgcBZ9RsD6M0
fmD2LwwORCYUIOW7ot4NF8IZm80wpxTW1dOROsPLril+Ys5fBRre3S/zCk6m
TrXg6cS9MMs3VQc0cxi0df3MuDooNgp7U2Ci+er2cW4K270D5nUT8GOsmjVM
fi5k1s7wfhW8aLZhG8iY4xyCwf/n3+HSvwzclnxM1iWTdGcMIOj89tq5cn2Z
VWTh++yM8oVuzVbqtYv6I9A/XSGVHJJi63KZ/qR3/rEPtBDwNF8iMDtfeYb+
4UB91oL3UfvA6lBRX4eFgj1Ap16Mf6yJi1nBcs/qIt22Zf1GS6VlwIL7uXfA
+koEH4ZplMZ7F8aI3ml3jqTgOwQUl21aIe+tfwf89+ssQnspCV14K+0WUgz3
W4uqBV+Sd4RTnyuu/cqskJHratmlZQ2sje8IcX3NJeIMZ66PDhQO6+Tip0Qw
HCdD0lllH3h80exNh9MyV7NPcJ9REK6OKl2RN/AmumvTsoTI64F4OW1myU/o
8v8SvU70PJcAudgbIKeCs1E11QOluhwlgKVabIn6yJSWrztWvIpPndFsvyXd
YB0NFw2FZr8BPxhFPTD3QuxwT0yf7YFQg7aBsTTDryQoJDrj7MgpAMRdU5cQ
hUo/Wg7qRstcH+Oil9ovSVwvDJj8J/e8wx4Ow0ZP+gyZtEu0SVgY9V7H/b2B
eSQJfrqJttMm17vkWzApt7D8GVN2eGEcpkZFNaSFxi1M2O5aZ1R+1aG4jLvj
WzjFzSBggE5xnVO04jLta9HO+YGY6GRHksO4DoUCZCitlJVX/1huRoGBqwGZ
YgVcd0H/UoJd6P6Lw/w9ESJd40ZFjCgFu/g/OCpq/SlsK5nZ8Ti8c3AoPtAz
5waq1miQ7Y7KF/fAzV+j1VEs85uhHT1cvlK5e5DLSmTJp5qOQ4Eo8amBX4lc
l7UoQALtDFqXbvlcbXB3gIt15N6UM0NOImVqnWALt2SmsrHogxx1hao99U6j
YFxIj2gUpHsl4h1llSbNU/MxqenjRycodHigL9OlxFHtoVk6dR1tH3ewtRmX
DaInyqlk+RbST0kW3j+BVJM+ElspXTlPpwTE9wP59HIp9drxD3nhZJZ2Ke8J
u9OouHL+iaUQzLWAGxkktu/MXIad95mywOiMIi3Gux+2T3K+sJUPEefMZdGC
Q9ohBqwtdMwjJr1zfZgNmTydJvjECzjLuEgKu0fHPFjCk203OX5mxdDk3ivc
HkxJBWoytQ1+fr6UB/sM/iCKw3ejJ3JzbWOuFLjyHyKFJUQhR/ICFW63aMl6
QJAgBbRSh7ug+xKucg3o7hIO5ftNWxSo+W5hdeiM6UTbglnjglTELU/htrPp
wz8Vs6uHTRh6mHPgYt1Ffj5vLu7SEIP3FPx0c5y3Js06LpKsAw1xepie7fFr
IJlepIw507RdWQNVa3UiQvQfpwEXHjVkidxSfV//50WcdX4f1sxlTlXtkiiQ
xwzaw81OwrOPB8g1lpBMOP34TDuJipDbSBi2ixDt3i5VuRL+KwdVjhLS8aSr
ifAhUgY7O58cosGDRW36YeD510zYKKtdw+nSIQ0Nl2+kiTvCv89X7taswVJl
4Ky9zn/Be8AOKQ2NhT96S9BLYJvT//5c3fKrjEuhk2aspj9Ex2ObBrZYBaU7
A6nEKh5Hxx16H+QapeXSdkSEgTi8edj9g47oe82K7Q9DUe4ejKlElOyGXfgK
lx+HDvsSDABXRM4K8uB9vmuTb/wYowE3DKRlMmQ53U5tj90yHmdWGocQOJrG
g96v761TPAL6eoFMcLlFVonZlcUTxU4rxzgoD5WJy7hrqm1450sdaZ3a7LYP
VyfXmdxXoSWe2IgUMPtM/J5H4PSSuRgvSsUY/BF9HRYhs4Yra0Jjoqe3lBGX
wY9c9JpKEhZVOOlEZz/xu7CkSjvFMcnib/igC/qKZzJWCGA69dw1YrUxcCaD
Fjfq74ZsRVB4JyGyV428xMRKeA8Jg9EcHlb3ZRZSY17HBFws3S4Tr9bsLcIO
5Tbyusf5xckkmXL4DcKkK9T5GzCCMmBHWap76xGRgvuvZx2bE8ShCmZylpwG
bh6wVqc9Jm+aiKONa3D2YoFah8lxKqNxLxkCcbWJRto2TFM+9lQe4Hw+iE2i
wwdAo6aEJjJPfmtKw+s9Piuv6by3mMbz+bpmz443xWZQcwf7HRqlMUzpPptA
Dy4WXN2apyOnnVIqVlro1FXFU3lpURWTGy1nv+ffuLarMEcHQjgVVcfR0Ta1
KgfZjRKhaDG0egxFLPCIHK8eM3E+ULBk/+naf7B67N9MNTiNGhOPBkn+rZeF
OckWio9QVJD5/Stgv+IrkNhXOPPWGQ8oi4YnWQxsZNbq0039YSgUl2H+ZGcg
PbOwaLwgmUej0UJYeQUPmINnzEUZ3x2YDSD/X1wBvAIyJp601iYe+Aoajjdi
z3QiX4w/sSD3CDfmjDtsiT0hRa+pYb3o4SejWoBjwmO8EcWyP0ObugGGjjZV
n9wAMlvvpiCuHScuHPjuUIZKbvuFjbJq7nqJ135Z3cOCnOwIBNHx99ogv4Rp
i8XAeEDwQxRbXtljm62/fGxiWN6gUtkg99y2c1jayxkGBVn8NhMn8rIZ9cyT
vs3aExB0OyvyQBNUvWw5QsEyOreqFXYJi35k6aBGpwRJxqQM1vpU3iEJfP8M
Hl26hEkkKWkYj1lb8G+Af6uCgq7vdvjPsIKzTxM8AWdWq3D8Tf4D86W8xHBa
7slt5NNpzjTOO80kiPFlXeBVCQmHIRUzqk8ucRDwmIYnkuC+5RWOYYwOAZav
VcMZ/1mzKvCT2FiL8qjLIlLQg3+Qt4msunXRh/7EraWlyu34zo9XpkHX+g1h
FKrT0E5MAkm5ggyGW3bpGwAa1H/MyqXnTuBgjveoAjCv3Z8zyulQEXvrfweQ
ZzkiIMhJn1oO4USqrYAocYbHHb+Sh+OSklvxnysiBTM6QE6L8LrwhAoGqPBG
UWCcpJxFFfFKEqXK8AxFPGLIdgBL+CAOjlEga/EYPlf4Rz81jA9I3IyeXIML
/vKqG9wh483i7MrlMIk8rN+fJX/zJe/eVolgQBh2HUPFkW7iI1/ChaW5n0sK
9VFD/23xvaKiEHf7IzcOFmB5IOVbBKAC6c5Bm9FYQazBc/j/EdbTwNI5xeQN
xowhUwzwR0pKeTOjuQL7nze3gyXbfjuJ1qYZYqWnrrn1paZlleCr2S/iYy8S
/7dHnCnF0TVuL8cA16s/asTWAmWbopjzcIswvNDoz8Kn4e6pNzEl6maQs7tn
78A54a8hFEz3vK6hjvx7qeXy8r8gIgXpM5tIilsem00AWWipcYhJjA64HWQC
yVrtkGP7v1aPcbHqJw+LuI4ItgKkAny0IO61PGJCN3cF/YDK/BbQ3QmGgPQ9
uVNcVN8iURkbPU5vIssazlEdLNN8u1Ik45y+moIWpCQBG4R7CCceQq9HStSH
SKCjYsrRpjHpDZwQOz9E7fPGGgu4jSNnQmiYNvevwDjq+QVC//KM5HRPJlU8
4/SM4kqfiygDWT2q8OU4+eeVqmzGrANIIFM6JY3PdSFSo7E845ns4tTJmkE5
fHAaUNd/hrhYtfj478bfgOZYR3KCtqBGTocugAD6v64vNAaH8ie5XJhMLj3D
9U2DNlt2D/efqoboNyoHHQFhhm+z8+8Zp7ZQzB/ZEFcRs8BnbxJF1tqb1Rd6
h7RoPp+nc4jsDq/1BvfXI4dZ+ToSs+ltf3VkDzTCMvIuTd9LsMoQ7zz7NfaT
cnnvk8BTIJQ8lMw0vw+jXNH4cjJ6sX7Hf/DJ3pkxfiyX1RW0QAo/ugs1MbxC
QqPluu4s6jH/ryn8swQB7gkx8oPqcoNQR8WhYjclzz0Ag2csAUOZmzdWTEdU
MlQgfbGvVMTNAph/Khurasn1xkAGPIYqsUOXRKBMFi6aF2aYIkDzSHLeQAKo
swDDcK9UCVJ+k6WXUVtI5tof0B///i+ldSTcqjh5PHFtohNXvzMTxfwSu6dR
CXC5yeEEkvUVfrXhJ97ZqsiXmU6zVNzKsKqajrLG4vBDYXcy0OldfveANJUU
eToowLEM2dUoFDLkYm6fxNANSaP7aYIaegTnjI5aJpg4yxScgUEGrTPNZhpX
v86JpNpEhRC8CmMYf9UIVPiHedeCNlGfk7ttYBjxKgnft7JzCFOXvKishZVE
Pp7Ltt/l1+DoyqRQMBeuMUbOJkQNasgRv6MGwtVnYeExco/KubflfYpLhbub
nS/V9v5SRn4+cQtt1MRZN/TCccHLHLWQOMZxt6fBKU6rdgoKLukNbbegHhJ3
KRyxqXYKNRxdUqctpF9rB09Rz1gzuvdcGWQAfu1SF7iPVyru872s0EYlV4t5
vnsMwmLkn2B05uvUqqt56Qj57f8Z8WQg6sv0DQUOuFsk6cX4w48Esy3/8VEV
3NkRLSWpjx6/CclyYOg8JWgSy6BhOUMUmfvMZcyHnAD50Uydbq48Ns1Yig5V
aJCrIQz8wj0YcZHS9HinkGOnTDlZDMUsSE9/ZoALy+bIUlz1oBQIRUGpHM2L
KNURsls8QMj6GZABMThkKDZY9+Rj+OkIRfQ83tRNTN/fJ8Fkx7iUYpfWdKt6
dASHo8kVaiMnrIbV8BSG+lTrYoxVQ9TGkTFHd+hXW9bzoTeIIDUGEOP4BSKF
MY/Amz77f5ZcGJVL+PMU9mtU2tmUVoyqHFMmnVms4P84EKjMvL6uUe4Mij1r
cZ+o/ATfiWpNCe/fXLlMjihmbCYcdzKbBnvoGEjTSFU/DgOxTbHoEHk865GI
gH3ySHYVj10zwjQGqsgH2UQgnaXV2Xi5VctTka5H7rtPy0tKSJLFpCXC6qwj
XL7NToa+Fc/m7IMKo7n2pyscfU6Tj25ADcrBYkT5LwWH/DiA43+9Puybh5or
YiAtqZnMoxE/7nzUXh8HPWKF6G0SxHRQyvbXZcxI9r5yCw4qkSQCzZMu1LHN
wzj2fy+CZLbga+9OcmE2mRv4OCY47dOeINE9Hbc7taENi9TROkHA1sySJTgM
TPc9ccjsjYdNOP1MRhg9KyE50Gm0NYK1WRl0DGtpGm6r4yHEBSh3krsMTIF4
VQuqNlJAZGp9lz5i3uACjvLSKdSIg9qpgomEoBEwglUfZHDUVXFk2URIHiR4
+nylD7KAngIFa5SWcQva1++vc0byso1E4TraBKnEoxbkEeBIRxVlBXpozeXj
XpY3GoUzetsYobzk8I1HXsUySTZwZX4OPa0j/F9ev6NWymuSU1GOAJxBovht
FMdmY6R06DwvpvGqd3LRCZVEAKqUSG/tLfZ+/BlN0cNR6M+oZnu/oEQeO3ls
fRhyQbohmQNPgGLofzpQnuHpLtCyp+KHF6/OiRb49kDYMYzZ4YUq9k+rZCIX
rsk1CRAWDxWBLNy2JbSGg6Kji/97y2a7qcaCbsoilSlW/ASGqZPOvbMrvXkq
j1SKPev/N/SyrBmbuSV6HJQfZeVL5zHuS4LrGgPk1J7oHyqvFv7n6jY+quar
iD9fJ/RlCwAg3RCG9I+OK5uzGEiysrzLWr0pHf856FuCJzlgK1pqXqOCmMVm
jrU4Z+V5fjA/RZ3CWz2oSZ/qxcepTGY3dlr2LxPIpoU6BN9QCxf6GuQV9zn9
H+BAvI4UletAFiC/KqzNCAF2EY/z9eVpfLaC2qqRa/tGq+SHy/iJchDuItSM
fuLvbneLeQ48066xEK3i4ZhrYrWzKa2bYyUrJV1/+e8+Ly2Idp9zfzq6tps3
aacPTXaSprbcPbvtwWXPLcpwcgvkm9Oz8+eTLndNkC9ADu0rot5ZMB0bF8WI
vn39B4OecjwRrBbZv1AobgflSA7Udrr3Z798oacg7iZ82vqrmIH9N8zT+eaN
1+Hv2h1VpqG8Bz3kC58mc+kxyJOuVn1FQluJ4J91MtPutiBmjUWmqbdimxfe
D9BNk8F8xpsYSOwrPfRgpWlLYALlPLW1Zk/QeAP/kSZZcBpiM4AfIEmuDoGN
oYX6fmNlOKWIodTMUa2bvH8z3D7AXPkiC1O7gcJ2ldwuou9PUzdSIGIuUY+7
ZnWcjIR/Xe+P59Bm9BevWhospU8ghCvDMthHm5MMQuMho4i8LAfGNQr9DmsB
QH5Xhm8K+nZzjDLo9AfcF92sSZ6MSU8e/EDmkgmbtCBX5ojmUeolkjkRcxHv
OomuWHVYEZXg/g4/+IsNYV2pwfF3esY52xfc6SXqf/DDnal5EqFeBgc8zCLJ
MiRMU/Oqkk0NCVlWwpSfkmCuDrUkOY6vVWnyiUuVEqaNHuIXY85gScH4a0kL
sV/Xfh/sspPWonVlwBEYDB3Om0KvqocRefcaruj2ypLmb2V6fKYUoTKeiKM4
XZQIRzjIUNIGZ/Yma6/xXPGfRgY3eFjfeFPYpXcvASmOBtS57fuVl4LSxeZ9
wx4Vk+DY/yHNE97usNA7b5OQwFznJe8UC+zalRtjU7ZzTGBLUP1bc/bdc6fC
N2/V6NgFDQ2wWUAqh4Ek7N92beRdIZIzvaagY6b4d6So8XUjrOUhIZyNO8JY
dDc7V+i1oEvujiQXvXVwxn5RvnjSbPhm3hF9/EUav9VuC16BrZwnscNALOTs
xrK+P8yGWpsnfNFKs+5xSh1o10v/dqdAe+YF9tLRoRDqkzCAGcJYalIzOOgl
9sZyLirXRvoY7ljVaI3NsYUBOW8ITLp5vItYMWVWD+R8iRN30ChZcGw0RXrs
2dYiBix15cAmR1096NtPXcsguFe3TsOkLShvYlT88tghfZMyvSGQpTsd5/KI
7Gk1kgotbiPDNp+w3Mk1XysFBzkZtaQrwnwJ2HMU+SPqY8IsbymL0zSBAeEv
S7FD+8ndPAmdE67zxZgBtM/rBu9lTLn6rN7u85fpRG+VufP6QfqE1o2s/F2+
MGoeJLE7vj79eag8HD4H6XL3X9V4Cw6TNNC7aim09gxxVariUORJSY+gExm6
IHIcqr3u/uirwzzZoQsClSSiVLi4KZsYask5jGAxiRM1trFXndppRggRQSTW
tl63vrSw3/yLAhg+YWBsOa9ozmMWE3F0iym9Faci+ZCptluz4dYjHQsKs/Mc
RfHhII3y1F4Mf8ijJ3Uht1aPeSh8JNK89xW11G6xhAZfbZ1xURimcjiP+bFH
spPq5KSOvIJ3JQDpRpgUYAAe6QIuDuV7V2bQerGULxI3lOVV96xqaGm0dex/
THdC1Dh1mdeet509QTSZA0PYJRR2Tgo/BXCXpQ6iQyn2PtTX8uRM8Hh+JeFI
9cwJzHzqkbLwNr2wZTPOaekOC51CY4TYdId68S5hQg82CuQ0IG+Afc2dKMvh
jfbtKkkAhnqTMLkN/NhUDsjifWEP41JW/cW95aCymQqjgcBupbNAl5WVycjL
HgmHEMq+lMWVrsHesM8jERviCiy9wiQntr1/985BBowS4JB6SkNcs3vwlKQ/
M67UWSDKYQ1FtS6nYw2M0zLJqN282Ygr27capUpFPn1evUYByMs2dMtJZ2H2
4b0UiRzfoowE4AZ0PpF3tc9oY4HxixBl6l2T+CbK4TOrLHA/6R3YlFZEmsrA
YPQFpz4ApD36lrM8a44DCVv3NKz/jt9f2YE0YRuFMc4EUoOXUoaWSlJ86fpk
zdZ1tNqikRX/DCtyQXApkwsRsBD8XIbP8Dz2AApPfueNDOGnaI9NA0Wq+EqV
ULoDV+W92PIfvgYhIy1ElUrvgd53hrEIcjEi7LbgLiQ+p52/mwBP0OzhBk7p
hiWJYyO5LYB6IVZohEbLFhh1rQcWbgF1tO9AGTlHZg1el8qulRAxYeC4tyKa
ULZGNhZfAcoemc6M6cOtK9r8j+LUgnpkmATvUvywzBXYOilO13IUXYeq4O/e
JZO0aqKaz+tp9WLSXN18u2chinni/gqijrjUuWQMCE05x0WTcsKUZAJbDoGb
YNCcsz/nkz3bwfEUMNrMa9DJEOulYDCW+eDIZtj/5yl1syM+4i4HV7179SUD
7/LbGat0ZI5xVigpqCFRxFS+VNIOsJ6TpqPdto6hRkW1QZruTODqUPciTcbZ
f0EigJ0uQIVT0jYEKNfusx6P5p4de86vaHg9GhyAvU7WjLtPJFOvVECk3OQW
LfdU0paQDJ0Pt378QlCcpfKpyi3L/+cFXHnOhWQo8PjVfPgkV6kMTLU/CjP9
iBcQauJ8HsBLP+2fltkH1eh4szVu8aN5xNiDGwziCzdFizicz0Q9tOfdlfSE
t+VIWmc/prVtOVj6ACrTfW+2HBUPbORydNb5sWZM/veJXj/AynZ4jVQGlk7w
ZJp0F2Cwyt9RIsu7s2dBYxJHlbE9r2Rl7uRqsQoTY0CEfrPh/CdL1wsgNWuP
JtVoAJ28xj4N1Z9fXu/KXu5nbmWadCweDKvub5drKfFWBR1LzDIAwgQMzQoj
EC1hWinHvNr+VgOu8hbZP6HRoDQGytUAt9DZs0LHUWJBMzhAhpy85ns5A0Wz
AZNe8ji8vUp8ghkv66yirCSgOPciLlVSPcjxvWWOvv2Yr4TzIBOPdZDqrpLp
hmav1yMPZB8fPYsug6W5nJ9rcEV+gaCG86y5gMarGiBhLGhjasrCUBzmacP/
Wm1lIflTgMP/fuvh+FhAOfb88DvhgdCF/cNpMbt9aTGKcmDPrAdrKKCyGkFE
wY6PYX6VE5tU10jFV7nrcuvDJ2twh3pZDPSDtIezbUoooQIcSI2GgytYFnMc
F2KfiIWHY/+v//veKfK8aRCTOtyOIxh3G66OE7E45eINuqVEkKpWNxSrhJxj
p81qjmiHF30+mKNS0pjAKySUGU+6MWV1lIUrOdpE+qgVUQULbT7tiBs4Hhn2
VqPQ5Y5S3Hz1tYi/LIz8LECVR6HZ7eoO+LHyALeCsZdohHCTYWHj2q0gQKLK
BDyl1XNcnGq+Z4k2lwOrUVZykUGv4aeKVrh2RLrQzxNyfH0pTf1E/DUszUhb
8KBUsP96NO0duJACpzC8fYeNPNSnhFuUF/JK/k5utTgSCkdJ0woFoiDbbqK+
mm8Xm0opj7cqra/7Wb1KAymdyvPlBDHf4kq2qqFVYz6YzXFvg+L+z3ADtdWh
zvNvTmT9+YmNQs7/rGtdwDuNEZky3ehDqUDMbiCqGm5AWFGUkv2n/aP10wzz
bVeuGtysL5dBZRExHKhGJKd2slq/d8eHAaRgAz2UyDycxgiHJ8PAXGmoJc86
POR7nDLSjBHU94JZzRMFczhmOCBP2TYuMovi0d0b0ml253s8mFNgTYso8+/9
xzxBmMuA7zOhzP42Azv7ZT8RFI1d+BDGxIiV/O51JNmCZu/ssdR1bE9LLKua
uDF3pdivo+kRXmPtVrmwZ+MrmbpZQPDSruTqzRZEW+JFXXfuNZ6QRKnT6+F2
zzitQQvfjpUtyPmk3RbHArD2BGvOwxT+RINMZsGGw3tkfN/K76I3ec6DegJ3
ILUw0IAqNeENixmwpS+uueo/gr0PJlMqxGDRsY5NElTH2n/0F3c57Hs3Kxi+
4XTkK0J3Gm8kTp0MHdQY9eNxhapfGRXoHRP70/JbEypFQyX3yRlWwN7cGb7m
EXzBpuk+rF0Cerc5cSIc15YJCVgxNeiNqZnRk979FB8Dg9yZQEcNbJk8edt3
ZEgVHNGRB0cKaDs5ulsgevTWx5tdgfpe4AQObXvikbQvOBIqs3Up1t35jznO
tlYgc8TDcH5rS/A/M4nj4xGj1wal98Lq5wFYMcwDFoQlbzCvknkroxb5PogM
t39kUbr96I+k7hMII1GmQyUHUshwjY+jWjs157+ZvKRYUhmfI9KY82j75/F4
uCZKwVgQEldN6F6tKebDXbAYMG74qbGHLKiKS4VMS5S4F8FqKzOX41vfm5qR
HP4aVvEj1yVVlvBwrXy82zDY6azEObOsiHNAGgH9x7yZKNUgYVCoua9dtUgq
v+KIQ2Ek5EXp/SO0JZsx6+SiqQqh49S5X3+H3QKMjjS24mmod8AUMpfPxpO8
rJ50codbZiVWsxHAY7KkKo97Tc1Mv3YgtyokIpjV8FQ0Su6iUMLuDVq1X9kb
EIFfzSiFGH5nnSYM4lvOSKsOlm4I6fQ7q1ISU4IOuV0DT4Xch2K17Sdckbj3
1btJq8efQMLL9macYdcpdVWWxtMdI0hrxXVuXY4G0gJj+Qk6/qlkKQ7cGMs6
KjNdP+/Udr8Cp2wWHOEA03TE4CbKqsC1xdiho2PMdqeu9RYJv0uuphvqDb9K
f1ZoXkIx9vaELK5TA0hr/i90KCy2+lQgrHLZZsNrFVUDeOZuX049SiNZKbZO
MBYBm/3UyeWqLtGg6oSOU5gSPhY//MYs8ErgcqyY1Y2L9EYl3WadRvIiQ7vb
jZtfVeduxS9kehCnrm+jFE/eerz3bNQ3iN8+H6B38TTJtDL0hUgKkNvlFseH
9RVmf/KoF2wDneh3TZHJeakbV8ltLh3PSXyMy0OJ4N+/VPsZfAmR8rLSS6gu
Rqk+tGBKblflYa0v15HuYHhF/mEsnyJEPXLtViVieRB3WpofNvljXFqvjEex
FavyJdJJ68u8i+3bEhfCYvnx+1wqdcMBOBLaTnMk9EyCJs/tBUDnl9l2aHF2
jtYa8Mp9v7xcoginVthFPe4svL1EozRTGxfDqi0sjqGOPfnwFalJNO/aX3DC
imb6IcJlvyIKADfzVf7gKK4IQT3qahlsUl1FogrZWn9uhpMwPTTu1CFosmOd
8RjAMHTEl5iPBDpy/e9zyKwJm7DiMQRcvIOWjxeGxRxuSa8okkUlVndDQH1H
SBU3NxCJxCmrzx5y+BgV7QBNLA359ghdyCXTjMn5TYUlLRtZEksH4wZSoCcv
iGsRtzgNzY8NidP4QmQRI3ITMv4bYeRVBvGmSTGBLLM+s9p6JcaZ08mCZxmG
1yS1rKpkPzpCRckHG34JeGoMPk8tpT5O8G8Jkk7bhig1WVI7D6fwburOyii1
awOeHhLMVa+AJ2BV65RJsyH1i0DdvNexiV5IL5g/pZVzp7D0s2AbMx9BQBOe
iJ//mvB/ynLHMv6JcVl7qgKrvX43jK/yCo8O4xs8zRMQ2PfkVXqGnwqwOajF
hWl/gPdwkBQGmcs6mQHwECq4xZixIJNILnNUs6nHotjaDyjr7zgGTU5GSHcf
U8ND1GpeCXFhnWBJQY2o6nPXr8g083/r9L/td3/FLkfKwSMX35blB5MHWBJZ
t1Tmt6KOTTIJ8ltC80EIcJMRv8prC8mxgoj1iULzqCSS4oQu+gpfneHBCJc1
zdOZRWp6kHnJF4CZxFcXV/ZLoLSwUB/8Se3EMAWOdrEt3T4d8nppF/gkewsE
yVlLePKLXRK7quLf7yMF89E9ql+yUXbEJHmQi93nTbah1+dGyowYb4qWFjkG
XhZ536MQcS424Uf3K+O/seyYEAV/OanOd72hQgU4V9kCf+5X83CHPiFq5vzx
lFgqKkalEEetjYlJOC+v5AqIv26q/M0u47tnxjFEd6xgB844o206VDaeLW95
6cmJ0BUvQEl9tT9FwUWFu/vACtbdXk+CHJeeLn51rHNYmpUMcxCQ00+IAZjG
RwryXl270IgODARvh65yu6lgnvlH7m4yXpu308LXsrsqAfPpWTPptWpx+YMC
No9HF42yaS8JsY1va62htpeQUbMn3qOOVqfDpVOkbKX3AA7dCHGESk4q2zTX
d3TTZtRgZem9O4E4dvldJUcN8WkRICn+bUqVy7RtY3u/BDiBMUoEfKDqWDq1
LSU/+VjuV68IQu0+aY/6pqubbFBe+/VjunHWs8nZKvUuP88WvKpPmEgCE+x6
ryFj9oNjbu/JqN+orGmYOJ6Ffi/QqIKfzFY5RbSq6Qk4yeOokVZyHDcfuEJs
UvavodTCKOc8JM8Fo7DaYLOLV2Qzw4qgBKXfX5K7sPdejic4FAblWjXqqCXX
IAG1SFaFg66n+wiXtbS+vy+fXv8dlDjdK81zs0mgwRmj63joM90teFo9jFDz
PmPm1c/PRkbR+Jkqn/sm6kK/TzeaK+9+XypCQRPQf0IYiD38sVy5tH/H/w+U
jGo5rr55Vh0anIseDKmQXj/mrGVR3hIIJBx1qJlv/3FRItC+J0nDR2z+irQE
TvqYEVfNSQBHRVXLN7m3baS5lj/FTvBbRWL7b9lgPRoIPCYpHZD664mqoRMI
Co8uwHgNwPyQPuYoQubI73R8khYDb3H+8bgOx1ehGq6VW1PU+D19obv0n/lh
ZfdhO1ppggUYdXYeW9y08o1VrbkQShdHHDmb6OuXfMvwQ8B+Joh9ByJLKcI6
ev8HrzGHIIhkPPDpGomiSGgpwedGo+pbb8SXQe+I9w+XVwF+OQ22oKRuLmM4
BgEcDiN6+uMm1Fv+Jkt+qH2Ih8bRA4tLyRqucvl4zz9A/pOO6ZgPwpXZ9WyQ
1St/p7SivxcazwEHuKXOBbeR5RN+2pEYyD+5VnkoVajeyurjYICtCtgmTetN
tQChhxj7ykVk7QiSwNz2pb8c4P1Vesh+HD/wvo9jXjza+VXDbACVYuQuPy4Q
Q/pgPJ801IEpsJ8aIlpRf7jwMbr7AAlDJ5cXYZuPcOLsGjqrtkhilbZgpkez
RAxzt8pUj4EUwVYluZPHf5dvE0Dz6u0ZvOCQQ0w4CM8s75X1Z4R2s4cM78Fa
Ai7YONuXX+e0rTmaBUzhdV/1Z/oiffnCMM9ZcPDq3r4r+6GQng752GETF+WS
+Dz96t5S8chCDmRAbNfRtDiUXFpDrvdHNCNzqbq3W8ANiEc0tbGMJ/cLFtJo
/QYlJ2eRWMGuWfE3LQvJRBwTifMTmhJKNNuiIkrkYxpIT1sUNJdFIsTcLb0s
AZNlgZpPAO65OMbEyGgXhj0OgLUJ9Axtmb4o8CncpNcbOIEctJirvYLHue0a
9bPm4ieDe+Dvlco0FzfIVcws5rLyhiFQgCPvWLPvzwoleEyNZROSptQm9IR7
5iGlKkNuTUPhGail9L8FUWqgsEZmcCklmebdCbnAGNvCm1Dcj53rv3zeQGtB
JwY5jgYesx6PMPyYawSZxsg90pydaOjV1yY+r1HKGPwCV5BXL1IELT+KrAB3
Xkc5jmB2Htq4dFFElJQm+OjQt5Y6wTjDe2TycoEohpvckEHe7144IiyWZhyA
lQNmWN6AXXrJAtBQ1eBTqOV6XDIlM4PIWFmJBRQV4/oCZSzrGZEcZi9ZOofB
pWIJNgHwFqUD4fCvzER7nzwNRA5Y9YtwyvaZL4kDBj7rDKNUlvPaZTwRRdj6
HaELRQ62thsyLfnTNQdPg/zdpMUdjOxycuTOrd/CAeY0Jk/Uf1ZvHVlzsIBs
Pi8d81Rq1O2ivGuSHTvtq8tyRdXaUHVHQdgRR0nvmRE1f6qY8iOrI6kOE1c+
0Z539nUsnZZBF6Sle+Ktw2NDBJ3fOo8BaXvWxSgeJjbzNf1TeX2LuEFb6si/
R+FGRTa/ceXM4X+HGUIjOteF9d0gogSF74KjCXHlcscdwX/1LB8bEMhxS9B7
pfMUe7u244lsErL6ePUUWQF79cREVXVmsYraHW34FcEvVdk4b2eMpYNVDPuf
rRtoI8aZkU9tuQ8kVvDsR54oQZysCG0HRbZ3Mf+TOkIWyoVwKi3Qqihr2zzh
IuKGxKWvG/92or91pdGmtnZjusQj4bsRvwmR6qWJJgKCTzYwP7VsZ9y60YuV
v3rZaZfw5CoBO1TGiX1cOJ062N9FAI1cDwrlW3RombNvMoezjvSckmPRn44K
sOpa3lSQAcZ858YFdcZsb2XksEzCPci6t1gtMYg4KviDHIxmzqrbbCRbn9Dn
9ceRloWKyKwbXuSNRxjWTYlsN7Zfu9Wy/LxNzwmg2ZZbfgwE02ql2/Y0N0c9
CYTbPGfu5DsMQbx56X/c/R+syl9d7DyKpby6CP3l5uQ7TBjYRjlHmg/I6EBf
a41httQ3pF9ZDj31e3YJF2OpvcKiWqeAMY1Pfr9tN0S4X3lh3uv8rqcu0+7z
Cq4zuINeVvqKIM//DtqJmOgsTZnAMnGkLMHZEo+nYQZXhBOrupCQaxLEEOqZ
xjImAZUBsko86UQcxo8w6SRCSN9DUimx4psOXDuH1CkhgdhDFQVoQSzAefvG
/m2h0Q6k8Opy1gPNzLj5qJbYzgcxQP2DVLXFUT280gLVTI/ljtOjG20nD3OX
ZlrK9CROick3AaOtQYwK96lW3VGiFeY9XE52Uoo7fmhYuQtO9NF/hK8p7m/l
4U7+KSVsDjxdt9mJbMO05r5Pu59mPK3GblzI1GHgsf+AnBnTRoB1cgiRTXjb
XkB+/i/tbJH4ROrwxR3T7+zWqMTjCoQuwZZbh+AgyXVYFAllkYtMbhfOQJrp
OvIIPLcexxzjUwkBBAOcrqdnxYRHnTFmjywRs3vf3qLhHp1Krn60gyC1R6IW
nltdBl9tavq9b44EY04JevKHo/jpLjGrh6fKRGaZ4dLB5aw46Fs3r9KnPEeB
HFZD+isdtY8o2k2xKoS8OguGk2N02GwpdXN8zO/bgH8QAARnGTqS/wF5RP5N
Z/g7P+3aVhsEvmvoBMousPq2r2R9cnjQStaET3RncPD/BaVUtHe7WaNpfjzL
y1E1M4k8/e3btUPdI4BfaGdYQa1FFZ1c1GV5r11LznRLpjmagfc0r6ZC1tLV
ElbELkqyxvqBjT43zYxbaHJa64CyFQbvB0OaS2V1UhQDsVt8NHdvuYd7QUnH
5BrQizeSeuJGbj2YRikMCxie1cdzrjKknMmFq6CjVXcTWB1oI7dqC9cwL426
v2GBzV9eyOBpoX4yTUflzqxAuT21LW91IPoRvjP0afeE/Ku2yc1oxdGMa7SV
vz6yA5bv6+2MegaEvtr3wP3ljLeS5Umk20HHhbJl+zZKrCjWvg0sdF6roV2H
nCKuKWnvQV9kIpslYF3RKaqoMiWEim9k3shomIhyLlJNwg9OoOyX/oCkNR1d
8SiNmhyUKNwfmD2lC4Cg0hA55COYrcEIh0MMPwIMeHmdvfClRJQyvyhaDoWY
/OSO0C22UMbl5ZoNNQXhg1TqVtOI8lp76bSnPxt0ziwmpF+kGpmDNRkRhZ2t
7oyNWtN9+vPWoU/Ivt5PgI/xf2gIcm2Yl/D5RVOTtLpRyV+0eGbhuBYPs+My
7Igw2blyZ414FoDl1zpj/N5Dme3W74mI+DcJIsRpLDMCwgwYIXw986xNsrwY
wqbjVlTuQXF3z/OpAx0eAN9DuZSBMUVcxY8wiWqrEBlTnktai24GeguOTy/x
n9PKAFGBfPGyVB0UhDhb6fDVFWL0JKo+SDi/fsNULgX1DEyi2yhlMxnC6UKV
n/xhX07gF1OuWeKyu9zvQlDzXyNyqYfGJGcsi8ThfjK0NFrvoZiqpDk7Iu2u
sGvy9P3lP40fsqrrRfDLv9V8F5qIiTOTWka2UFYeNZyexW3c5OHw2gLW+Yez
SERPstL8MzWQuYZoGt8dV/coCPExW6D3WL/VE1Yb9eA6788oYEmIJBm3XPdj
n/I0Wec9VAOte3GYjA62XBUcMNqV5AO4K+mWL/7uoltdAmrF1EclqBY3sZyc
WoDaQz/FW6zChe7KqWT6W2yq2IQH7WkGQy6qHYOgS7YJMbkzTUqBBtmSloNP
xQibSmq2okaXiKY3BNfMXULddhS6875xLiZRlCMP03kq6Ndm/twQGyJS0g8w
+VHguSoi9AUl2yoFPOaR9+kmMs8jH7IVAjckEr4xiw2+AYVbYQCzynzBP+xl
3W6h8IdVGqXLYnMghleEqnt8anQ0zYPBUdKT+GcvmfFx62iy2osxhvPnqe9b
V9Kc986wlmhWDXpfroLiHZbb3dVdsEaztX+W+RYXRd6A17b9dV5IvOYJ0XPv
tEF66dBHszmUrMBhmmHwxBxE+Jst+6ipdPWaXAf5Sx2afqSrkHynp5cGk6is
Mnz/MeYYFYQ9uy+prvOmrWgVtpFL94YE+8Cyi6XPl751hmIlctBFM4UmFhWH
CvZtPa+ZTn1XpasEV5X2bJzfAuwAmhPUc2o0WXU04Mfko8jskipcA7rYYqM2
m4q8WkjM8KkOvAYTEhQsrYOfu8lJjgx7oPVweMMy3krHNda+9QLBZ0XiSD1z
iIvFT/9B+2wfqBZQehquiM4qyTOBfLyT//xCUGNNGVXuyQgNRGIfcp0FfbSl
tlqli51o0Ga2WYAQ+i8hew7guEIMkVpLyuewDQVb4R16+DynLu1EqEySgXDW
stfNVLRWkdgdIhA0fKLmPSUI75IDB77YwW4JWMQ1/rIXubUkJwx2hUvx8294
m3m7GGobzThVwnbo7hZt2EJba5ZA5vQkzMghnAK/alDM2N/JIFGu3K50OiVH
puhMC6VwDbGJ03vDsDUFf0kQmemv85kBkw56ge0VguvdWBrXjnkT7rCxqlHX
P2r8kYD6faPyXeAf9wYUji/V03plMmSvuE3MxkroUyv1zt5OLTprCQk4phGJ
u2g2oATj31hdQx6Jt6yFrtuF7z9/06O8JVAsteBULXO/RS3NjTv6mcBMews6
izOsQXSgXJ2M91TrhjdhNGGlsZxsXvExXX95XMsNfhN015JDeKIDfBZQqy/N
tJzplP+0wJckmcZD8uUVzCSUox27fL0wuN1QIvh1rJ7eFX/JgZwkyhv5Lgj+
6owH8lR5U5BzR38+dqebWCtkOP/C/tjZ0Pd6znXDfubmIpMHh76RluadFe5d
75/0y7OS4Hzt93vu/opeWepfOwnz5uormOzB8dRZamaCX58iuILz3o7IWxxR
TLX0B6vuQF0yq8arwAd6RxX+v4Auuv0Ag2RnIgIfBrMliVunqX5zWCyaYGwf
0M8IDKyhddRt0kJMLuhCk2D66K6QevLRlZ+VP7xZAVX9YK4BGn/ANoZAI2FE
ckTcgbQmjRt/N6xEMjyu6KbPo0O7XUsVUlYxed/kCsSnUccEU51waGiMLI5B
7DvwnB+YOxf8hNLE7wJuGEg7HweFyJJZ9asG0G8w8+ICWbF2H6TQYwKcJX8j
HlTVCPH5cHsOOCijovzAVwsqXYoP9u7QlgfLvKTul0E9M1h8WWYEEq6rcL+c
iJ1taMP7A3H4uaQLfQQrXRdzT2CtXorzjTfcE8ue337nnuPvRVzoZ9JyepdP
Zl5nbOyI26ccoBoUdTgrcBO0En0xxoLqdXQ5IkQjZq5xnZZb1zybKZqL0PTm
omzw28gLh1uVBjmfJgiB94eDBphS24Wk3ajFOmM5tI4EiZmRx7zQfi4JZn//
5Q+ZUXfBFZhcmevOkMBopPyNG7hlH8m8FDNBXCcoV19eitsj5UEDBYXwUXBz
1/mflNKZLT/JICR/FD5cZgLMhLTr7WcBfYz3rEGw6wxey7YP6KJyRXXXSEa2
ipJvNOiKlqLSqyEeLqfVQD6hPL6URHl0hsMBJYWHmWoyWpHUuvnpS7Guif5j
64b/9mpaosOEM9lXyqBm822TFPnydSCERszI0P4FxQ+9gpNIoJuWmg8mZ3AI
4Phblkbi3DYnO8+bQ9yW3QJIdG1Ko0KRMPH2E1wuvWA8m4zc3vWrJI6/qd4I
kn5EDIDmogoEge1Hi9OyHu6ndx9RxOmZCKgGIaOpwh8yJTWzbNdKzWskxqKd
La+2tVpjhIwDDOn6MUwP5TFejJ5B26jq5gMhQcTMFKFthDMKK6VXNNZGn3k1
6VclT8J4dLBUC3D+NgWsQJHAghYQPUBJHVBxPO7wRzsGFSR7yHjDcnBcvq6E
i3B+CChdZadNDoPzelB6xWKH4RirU58JrbS/BsL8NE3YKiU16+qb71saJ/74
i/U/K+unE2okkgkrmzqVbhpakD1a1RUPGF62mUMr/guFK2XQiSXrk/2DNpup
wIW1UbUq3mttcnxhgz8fB35DIoKBM8sz85VunvhNDyP8RbKk6sVM4fUGlxdg
UvRJZWGpblwpSNkLWjO03PtkeUo7VSvxLLWpEvIKGqTcc33DoJ+w7y5tXPxZ
g0pcgvN4XIgkXE2OFbjc0SFuRkRD1MQVN9rafhc4vSLPq4a5Wz4KAit3WvuA
CqV6hJ5WN9FMhDWI9P0EMpXxior5bkKGKX7RZQfdNvH8+QQ0hRPOGDbhTL8F
+dYsqXmcAji4DJIiI0iIF5kolZOuLnsIwT5Yxtxvk9oco1tX4HdCztUR0RsX
k8JfvjR0/v5uzUd1jkgvCjxQ2H1bku0mZa4QO0HxuePYbo0VjOfhkO53hU+s
j6fW2XGe7qXVPnBLgZiR01q/pdqpwEXkkb1zv6CMzmJGJEjL2fQGyEohEnPq
fY+Qen5IcsER4Mz2hh+Mt4Ypm00CpB4Xbjbq1YVHvBrcTGhQxQ1Xeldr39uA
Fe+HOm9/gUmaMPtcvcAH6+4m9zDQqEMASC1Sd55eMmU/9ER9tsPc+Ae1ChSt
JNZsdN619N5n/WSPwPlrUINsrcf2rFksh3bL6BXR3Ryy2FBSt2CXoDQTHbe4
vWeM05QxsQK+Y6xZULs3yeVDw20BgB0f+Y8VHcCenEggF6cRp/oHxUnKnBNH
GeZp7MtOfpPzK9FN+iPQAENxDOrK1xY4Karftd6/iDKn7FM+scI+UNewoZbW
JTMPTGAaTmBANkUHfenPqhYRHAmYzUlzNdt+adLQVDb6okoL2zyDKdFOTlH0
b9SEk+6qG/wE9zoEBc9Suoi3QbZCoMZbRaWfH8A3KttoWB2F8VrisAaKIN5u
ggooeu5U6YXpHg3lUIskpBPWfqeH5uMvOtet48YNHYOsWO4ca/OIyMIisRao
ViD5Pm9dPVLA1FYimV4rqsbuCWItkB8tS4FqPahU5U4CVVDyUqCssxk/FDNh
N/0DlCkxktZr9FTpjGPfcAAZ3LFQPHnJmbbDmaOLY9fkEscYTeASMnDRS0NS
5XeRh7vZkLMPaqC5rv7M/MIiMgWwgM8JALe8Q0peFE8VgVzUIEN2CKROx09x
dwFHfymfHyNuLjV74dLlYfmzhWgNp77w+MjLB6ncO5VLICzCgFXsuH2pfsaZ
NykNCqi1zmSKLhPjXWwwNZ20yFfSX42Srh9Ie2sFOXLaAaw9Jv76Wn7dcZUZ
H/eHtL2aDbVwnzWfKmWeEvKps1TtkLOgildKJqQwaXugef59lZqOlaOPrzqv
BIzPBUNfBKRoYefQyb7dtGMRQ94TT43z/VqT39wO2aev8xjbzMNJuc2zhl0/
D4dI/K6JgNe8mAB5wVmRreJOYyMRZPt5zrJ+Bakaog+yQS5al8UDw0daAk0j
PzZ8IRMZDnJ2H6l3eSLN/PR28F4clce4grpo0gFi8iX1RtKDIpn+1aI38qkU
FUXz6J6T5iFZns4vtnldEretgl3ngKdgiDxQv+UxPkSV8ihdyz9co+cQBjya
bo88ZjP3IAStPV6SSbaRmTIuD1ezvukcmtgAZW9hDyvB3llp4WlA6UnBXB0p
gl4LOwD2UOHHkrgXWSH8GTJxJQrBGW6EZPryegxfoBs81gaSyHMyvimzCRkJ
PcEpKCfKGIQwakxtam2PGcqZevXoLCOzRYAB0r0qPszWLvreDjdE1ocpvabY
yhbdf/iH97Tfwa/JJgme4TkDpWNxlBug8gWJ6voagSNhX8vtwOqx59nzKo4v
duuv7pASIBjiXeXBV1/jskTSTZUfP5o4jLQOwYdNCy0fboDMiqlTmlgOBY5A
YrSwPz7rGcnRNCKbsQ6DLF8rYs+gUF4w2qCkqq//+PlhGqxnZGW+TUEtlslU
PnbJzWm4bIW6cUw8pUflKmCmYepuL8jwh1kSPpGKq2sVdXZaG8kO/ZCDaqDw
o37A2G3NSZ+XwIoCJYN+jL07j9LT01Id0mNrLiOqfBSlc1ynTIzMqC78z+wK
6TM4CVPIaj6wgEpY3Mv/NzzjDFHYk1ymGgd8VjExJbzmYvMNUCmLEQTHMnUn
K5WgQyQkY+HsYJ/qwf8s8loxNPmFQcB58mbAoDscw5qeTMiQBBNLZvs2y8NA
2CMJru8YXvBiRWdSi7QIJN4uhYbTw6yA2RNScY+5nRDKbiBlBwJp3b1dNNwX
cCGOSWUr7CB3nLIQPcTQAHZA3zwRER10zv4Nph7Kup0Oeaz9gRPx27JVx12J
9SJoYWIaJ7hUY0grZEVWd5t/0qQOomUdF31tHaHZFLUV7HibTLrS94xUSsvC
0NYj/f/Q8q2ed446fh/PPvxg9V5OncdHe8q0HTqPLKYgLQ4vxqtaAh1l2iGk
ks3RMWgCRNzqWMqSTF4klHkCAtFoTiS/9GmXJ9YDUB9WydFIXy3qzF93FB28
Lyo9d/VTQAJrKVSFV4rCSbfb9XT/oSSjI07Tmw3V6BeJNXNIj8EmU9QKPwug
oAjrdxv9cVH6c5xlzf7GvNF0uIvpncGjzE6nT7SF8mXFya1KV8aGxb38I7at
Y5skuR7R8eKVJ1ppJYFfV/e/cxMlrIk7E1yQOSrD48JquVhRfH+O2fkmP1vY
SujpYJpdIGrd8iw9wh7QS1hPVcu8Fvj1Irp7rt4mW0PPIFLV2f2yp3Wpsxx0
HH3XPOlzQBa2NRo6/BYclfwm3d5zCGJ0y2/0CLLR2zgFeHMyDH82WfwoA/LM
J5ViUWdpA9BOaAz1SeLQVPXryiYTR8JsmL3C8ycob7HfocG4/V49+HBcGfT0
YE89UKzBfGZg3H62s7R++976UkAfAkl5H92sshk73lE7WlJ8mcEvs6G4nlIC
AjFZnF1YYh2di9jhlUo85j43mz9gzS6ClreZQb9FNt1Po4U7xGpF+oTIN5gF
g5HDo5gGebga/qCrcVlFLv2HYoLCvpIHt7Rb1V+f3eaUodGH+J1GWSI4oY49
5ZcKq7/Z0wL2WiQ3yt0kBBZL++wbj6jwWgdTHGqvH0Tybv/hA1z7rqirgE2Z
oG0F/XakrNtm7gemJQODeIsE1Bfg9pUtzglCrD010pJSYPFfmP2R7CmCUCRY
9G2WLrRATXgu6654ps+bo0fkVtui+A942oujBXJjerGHATM7Uzbwc1pcOLtb
zSPUnZ+P03cVSvAFQ0q3+llVAuhwy0Zb5oi3ZSwQtpauYU+bR5+d4EYkXVNs
kzz1VL8U4hHz0fNnGwB2txam9Vjw8OFYrs11gCBMc2AAF4o5Vz9qCFvpfDjR
TYj55nlqIngIumyeHPuWKrO44JXEuWYd3o+Ny8sqEkj01XfF8K51GCSiGYeF
NHo8huH1jOjF6KtFabXezaE3KOySFx7VI2xTmCAyHuZzLsoKMHYvcywZytd2
FSmQF7CkTM4/Qzd+W6r7mzN5ah1ma730yh2hsvzFG2DQpzu+1XKQV5SV6TuU
CjSsX1Yus5LV2DiyNyPOpy/n2NLTRobCJRAs5k6GAaOosfmvmA4vMyqJqOk0
l8najH03ROk6whuvjTwVCKFwOzvJr+gJ3BFH/h5F0v7eSahWakg9RlekeE7V
C1ytiOz/QVZlXeXv2wnkSQSvJ+N4DAl6n2zUOu2+9OyNLpUGZhsmSNrQfKh9
cNR+oyH+bu/85P7ApAahZR/M5XPdFo/B4TgEL8ne3JKttpRfCbvETR8kS7X3
zRXQ1WUxw+N6My6cs7MswvkH3SQ1f2fVyVxcTxg3kqOy5NtgM4MBr7jA3mA2
mUl36skc7AScRrnfYsxeHO4aAPNdQ95HUhJOPCqeSymYd0an8ApIxrqwI7Vz
moBOVrVJ8Y3PDR/B5ZTUP2M9wcDUX2y2La/w1IpU4xN2o/bulGMkpHlXdJuC
fBbME/eG30DIfEUvw80NglW40nacoQq4i11R8oGe/RCq8k/vIyMjt75w0YLL
V4ZEq0Oyguh9/8qixLn8AhEuaqlrX+XK/ZdTS7/beoflZCZnMtC3v4YZLlei
xERwY1Uph05czEYu+9HZ1T7aFvNKZUQfudK4hPBGa2YRNKzJKsJPrvcEVbAU
yjy45wLRFPkHTzyzi9pLPrULl8F4eDXWdYi3aHx6zmzpmFamK7U917uK0JpS
GYKAp/cw8+2Lko5cq3tLnTpsfKbeOiXKrafl26DUY49/JLbOq+aRPCdo8sat
fJhk9OO8XiY6fHu0YFxI1V5raIC0OYTk7RCFFQfRNEGs7xkMNua6wu8TuwCV
seT3EizF/fz7LLcpGYeDGpNhmEeAfTSgsEnvZf+ne17Lx+ExCguUnvY4I7WV
Jeq/RXTw9tmgjndtlYDKGAUjoFNAaTznOEnLvGMBfFOSpEccmCQfPgokZ4E4
LGJMx2UI8Q80h3IeHt9qFmbK4E3d1enl010meQXk26Ke5Rq5YgNgwS/9B0i9
RHXdwOovNmgnN5olwG/GptW8q64McTCMeVl28Qx36UakNZc0MnB41pt0WCSW
SJtbSZhFqvR8uvHAcFwfoX+NB12X+7/urfVx0nZHmzXfpy0zQtY5ubEA2aeP
IDmLmzjkbFaPsxLpFk1ZqA4CRJ7ko1bSsCHymYSeImb2nXN1aTxoT6SjKX9I
dt+xrCje4esbp7pVgUn+zukYpdU8AYsZ+lIQuZWiyEPr/hQED+9HApCL7kxs
399CJ2Vgz1kRyToE8NXG3K6aausuRKv/fS24YrFwARor3eHjESjFuUwy02x6
ZDd4QOZneR0JOWimx38Zd5/5Wh8VHNzAYatWLC9wI2zAzqverUMRfnAhXkz7
6nMyXdtHKhDetK7iP9XffYPsJHFFlYchkWtZMW2aLIxKCr/YqVW1UwBy6aAs
ob91wlQ56/jXj7MJLEcvGP+17RV9gVxFJASOv6wr+ZkEHQ8jEREsJm30p+0V
OsxLmKthemtYYv08nOc/FF6qcm/4khizGpAkZpWKqZk6fTIUlDxIbUS+LZPE
txsY4mIBuX5EoZCPjYOU0FV2ggdttp1uLGzhhNIl6AvpWKDQPc8uJ/17F7lK
Vf7aQw8x8WbC7g/vrDbkyhs36qR16WqbIO0lPzpR37XSe5YAfw2E4k6pAsmD
+eTFuciLs6Qk+5AwAlXesErQB68zQ0XYB00nhIsUkRIF6ipI2otnkC0GIKfU
aJyCAhOZzpHThqWeemx+p+wskBsspVWd86FjyK9hdAIhh2ENd5TTrm1cQOaP
B/b0H7FdQYCaHszDvDq4tmGtdJAFb+RwYzS+3trbWu5Q/x0VuHv4X7hiRklL
aPAq1tTvB0a1IUumiKh1SSBIrguaiqUFwkhtKEc0jX3ltfX4yZRpSejKyLLu
KKsl2kBZoUcpofXmM63jJo+9ceJlyXB/vv1NBAabn+2iE3Oxkv8XJ9ZXkGbO
3AHG/Sv1GH4a5z1v7kvYTahAhVDPKC5RkfDB97EoDjGci7rKWjnuEQOn+Jx/
OcV+RhH3M0BVjZh1PqGAn7Mncc2e2ezp2W+TakWEpBOa/XjcoiZQnQdLm+DS
3m6xIhsrPnWhlN9JiAmxslJcne4kjctcGUac5AIpA/tga0Su0rNj3aqNoPkq
WmrR49/YZ/jYOtNwAXgBT2KV4/eKYyC/WjtFGEKbbuAJmIsk+TYN+Mk9xOpq
ypOzYKycVRgWGpQ3tdmotz077Fzh5JtMI2xtCVjV0SqrZ5yGyk5K/E6URJTh
V1EACYDQGaO1C8me7OaICfzDou2XWDH12pUhv+uuMCte9wfLLtfQ6bVlhOnG
U6okm2P2GUsgqHeg5TZIbyPZzA16Fr//Ysru5ZredV6MZ77LpusZnpTYeTeI
NbgcW6fzfQ7icG3P1+Kh1J8gvPzkkfxleH3wKFhkTR5Huu3JL+8SR3pU5gUL
792lMH7QfJYcSEU6YANNl3nOriYw1TCzUuty+N+GDMBsTYXfKMP/4cXNrswQ
0/JTm7lHQQNbwV1BRxFhiK9U/J+O7+C1E8vLtt2syrQRSq/krxpw4ZtKstt4
11XtNcBrRaExiB7nhBjscrMLuOwQ+jS2dO70ONrwYX5T54/hIE9Z8jKC2v5R
CyAw4IMvorgrS1ChGvf/yj5as6oE0elhSJ7531KhJHBhBckjC5WN01I9YaHK
wfVpaLN9LYDyhj5FyjAb1sCi3lArWb3wjMaiSUliXWwfsxHBklN6vUeDRbiH
ZHuS9dhLbgVvcZIZBc4Yb+dModI2Mmmt9BRnUs5dg0j0H4KnlbtzvEBbclnM
lyNBBn8zLSPeIr5anyuL802YGu8dX7EJrmh70Jy+87liS/KnCUNcgedXpWGX
D6C1zi8uyXVpAxi9YmHsTRr7A6PvurlPTtwL2mlz8hZbdUwQOcD2DIsYSoyV
W4h6s3NUeUy/qQ8jU0kUOx0dNjFN+B1+6MPfxv0sfcjwWR1SegwUdSUu6Zhl
+32lr401MtARuoZwZxwDm6s+uDHdbVYJIRlXHCuDbDzspnHkZ+pgsVCWq5ri
PrVAVnGLnO34gNRQ6laFloAyanhTtBizovBX5Rf1L/tLNfMARgypPQQe1UAG
4Do9EC2Xe0a/iTAXJWRE8W8EzPmf1bLkYf6y6LTiuYcbdQa2c3m1M8EzGq4L
TnGG0Kz5Z3dR4At2oxC8TWbCY8MXmXZEbvncuPp7FgXghGCWDA1yU1Uh2FRk
2NYqGY/+fFrlo8iQ6Cm0ROsQ7Bcm+AzaOIEpKxprsCfv2uaBRWdWe1PxY3ut
qvea4QpNr3ZKFJ+bo6hWfTXsNFeBunMfxf9psI1AsRhf54mXmPO6w59FGCAU
t2c911vM/NUigdgSqEWlWff1cyyXmtRnz4FcbTETg2jawJMlXG56oYzCFQ/p
77A+QtwhrmKH37hdPajbOAVAvQFNJoHFsxbS9m4HFJODNcu89i5jSVyrhaEl
0sGS0iogPZKKcr1vadm7noOAHpyPy4wBbfmhlr/TfLawK9RCLodTZguab+xg
0Lim4gOvHJYQBiXJOOAx7eiV9yvSdmQsRJa0iIt4vIVBk7yl6/JxkBmiVGnH
+VCib6ampwg+Q0mUJpW3cBBF7znCzAU48giOph5elsNUfVS657VHiMWWLcJ5
9JVwEBQ6xsyR8ZXf7cjio0WSUC9vcQsIz1K26f4kW0Y6LGYlS3Odat+zgfRY
MmsYeKM8ympd9Z1Lzm+FUUttG/svESDeVqnkiojQzvFM8RvQecsbHGdafKKk
lQpzHNQWlipr0ZXX6CciU6yZPPUPr2bDhj8Ec8l3VAGmV+7rBRgEhyx+q9qv
Z3Fv9UzqaZgDoDJmyQHnwD+SDxurwbnQ+ZSfPTCVgBzzTTle3D+KOg+F5kRi
xzo2QHbmIlbYQVrSvkgkytPuMPbSL+P2xZfYhQjFc8MuhwsFyMZsxBXD9KNf
x5Aoi2rsIh7EUUyZ6wLvv9Bph+vmQi/pSr9EBU/7lbVdqlpaWO4VigFe3g+Q
a4iW5j4us4qMExIRkL0YhH4AZplS8KT/ZOH3kX1l03H7CZjzOpz2iBmV+Wi8
20u2rSPx7IvMt7SmVQIfMPYoXilroPR5ZiXEZwMy6T7z/Hc6dq3lbuR5xL3o
jU3KOko4/HN6VdsVi3KGJyUvXjahqL4gnAD2CRs0hiZ/wtd045QJhls9sA3Y
p1/SSEDbKsMBggPHVXTIt2n+6g/UsuQSi5sL7EJcjj9p9GCeJ3tIIzlzMa8C
pVjqHdZVpRh8wi/Ko6D8F59VhNfh8lAp2zVyxywtY2CLPuBgBZFShjddwZfh
y5xVe7HStD9Rntw+I6XHqvdFSCdVcrbkogqBcrI6Gze1ECNanV8F5l2fj2dc
eU7zFn1EME3rdmJ3VHK8UF6ZyLYkDecFQNG7FgS5FkSWu63fAa0Glp4RWgsm
lFtPi5oYowrhLWP+GBEA+qjr4F4tFEgSoeNlVWKs4XV89i/qIa4l5Ydufiwn
UGK1NgHpyxfsxDmkmUvmdQc7YvG/6XxIgV+gHKSITwd/8FyJ0dMAuyFRu7R1
ZT9Yocq4HEKay199rQYxH96kskkSF6psv1WmQcgZPr7eta8UFnVTNFiGPhj6
soXFuN81eOb7F5QqA2wEUec8kGwDm6/6faQwxwRQL5y5Qn2MPXRpveXd76TE
kMxV4tWbZSzhVdDFqcZR85nv7gWzcPVk76D/C9XJqdeHQPpu/VkGcXAU2TzE
GH7/Fo6WunfoF4quaL9aEIibZTI99OROah7wGGo4ojErXjIHMXZ4W90PT9Gy
0fZilfni9z34XlcF46swfyK0PozcYQYyUANdW/BZ9DGGXPIzOTuXHg8iUwqX
7q51Oi5kT5AT9IR/jvuMyNIBdya3gcc4c2n1IqS+i+X1h5esfOsu/LMMw8lT
nKEmq3Z7cxmatXLRxWAxuOK4UsyA7pF1uJM6GxUMUr4DemLzFygfti/WAPU9
5HiU9UsYqonOSDBsoVjh427DiUGXlt6ivUvHhKAbKfW+xb7Lopa0+cMqTQrc
8ViURla2SyDShK36mGlqxj8m7dDvz32gEnCTXFNZ3QJH2b06oFrxEiQdAYKj
ILkWULSF63xfJwkYgdMZpV3GoqViaoQdOCS4dcIKAOPb4ZGhcZ608HKxnW5c
xr9oveNkR2fhaEptsPnBfSgOeymGJfq5syTvsIHfYQFIRRaZOoupMIiHXY1D
kcr9qa1gbZ1y3qHpl/YHM9th83tZSALSVnmIPxmI9JULI//diSq+3zrPiDsc
gI5v3IDHO+TAVyLIFqU9htLB5MO5k4bmck+Wiw+rFFg+rIY+wgJ17fIsyj39
VS82sZZujO1/c+GqrXJwi7hZhkdrjvzDaiYh4G9y1N95GIjD66R3mT7owu64
4n/mbsBnrl7OBIwA802w4uxmCUDiETkd9i3O1S+taDZOBvRSt/lRtCXfQarY
pY1zDFk7SJgvU9gnjAVlttaLwvxGdX0ZGpYYj6JexYiMWkgp00zOHw3w0jFA
5OHc+iGiEGldw2qCE4eKLeihY4drUFgqr/Y5VuJhORiKKiYeOMj7slJmIJWK
dcsq3T0Xd0/3XZ9hdgsHkFn15uX1iOn/Zdlq9J8XPY3xO45y7iFSBXZ0AZ6u
Kky3IkoMBQSMkvPsjpXa6xGPZwOXUqEsMZvpBzn8P9dV8xa7Tsq11PXeiMSI
u5z3MDUukNueS6juy5r/oiFAWLcq+944Vv00CKbweaY5pOPzNODVJDCILY5X
J95wrwJ7RpjmmBZtcw28+aNX6ZBwS1QeSCcT2H8BahQr0XkJkhvfbiOQf+UU
/vOdReIahqTOF6Srf9nxSvv/BaOePqijWZ0t0vmoGInrUdJIF0GGjumShFvd
eXPvUJXLvsOsKIH3rW5hvI+NsTAh0MPE7egjmcZZSD8OB5cNdDdkZRdRw1PW
f0VMjmuc3MebxxnEhvsBqKqOOUOGhniKBVHHSeok6rapsWZsEqggD+xB4JU1
AAyVa72LbpTrkB0EzCRaYLgvP2KUtRFGAHQCqDUlzRbb8b6UiKZdrDKTE1Z+
Sl6JBknNSwhe/DwkRRPTUPdl+TG46mPB40PWjkHzZNwRSGINY/jkWikDILrJ
AkNIcVmRlJqxp9/kdWcKl8RvZTh/0lcXpdpjRakKaonAhIcw7k4rdxQbvxVL
l9hT5t4IE1pRb/0DiWIHeK0pRqJPfTyPKLVoCnfOZY1dvC1YxmY4Bmafs4sB
wZLqxLD8j+LEIDSuVTSLcP1g+a96WmxjNrrjpwmACPLoKLbmk8pcBj79tFAN
7ApcDGgrXH7xdHJjkDOjg1v6XpgablwPqAC0WpZh5Vb6/ww2m5lY28k4zv2O
53wCNpoHyV+DN0hzUXYsAHzw/MmGDnOLWDRUac0QCK9pMfBlhO09gyaAOyKI
q0hG8kzswcU5UzlfYgbZ814+EAMdeifXhla1gJiUvuFB2FltLvu9yqeNqswQ
YHW/wn+RIGbTC86IboDfatw/jM60uhUIYnvi3qPPTQYDyoMoZ21jsDbxBXtO
dpLZWTeas4tRRjUnAK5UFOZkSs7mRPg2S5QzyLAD7U+GbJzSOCKWCtvCdg2r
PZ3s9QpFxoXwXDrN1NJgJtn+A/HkSK9uANnuReiQzYt4MZ51yQgmISogAXnX
wIK78ItaBgvr3/j7cCX78QW3AqzniSGG250Xqe4cdPEbliYMfVwsHI67n07Y
PFO+qnQ4ERd6/UfRM3wMDklcomr9UKSckZ6cum/D/2swWSQGtLFBb1RvyKIA
YQ1uBMBl+DQm9YpbfHO08gtOY37Hf0HYFRfV/pEilHfMSLlpMi557m0i2bAQ
UObTsHeg2WHCtwG0SklT5djWYNDFIDXSpvSd/TakqiXWBHKfFzq1hywOyQMx
sOCWScv33z7EhETY1gPwCI1Ve72jOdUzDm6GBn4u8F3g7jel7RD4gIzi2sVm
ipdb2EWwivOGs1Gypji368O6nDgQPlG5mWIdDkhNFisGbO3jlnD60Wj3rBOX
LsX+J7vXGSF2MiTWH6bgyETIkJAY0ha/B2xSCE4V5zGLcuTygJYiwOSd7FhI
cgdJk3cFtI/rIF3G9zgse5iV2xZIC+0JBVo2Gb/EIT+MDHwmDwGzeD/0un7X
NagbKT6K4VcBNQJo+yYw7N86DC1Fa4CBEOC32u5kFehzMEkyXMK5rQJxfYpb
yBVoE0QPtrXpYeha7DhU04KKMP6E6AeV2cSJK12kYyXZIG0QcGNkgb13l3Bg
6yFv/O0Qiti+bHmk7Yh575nUcNolCAEbpWZa29jy8KpoBWN2iUmKLNDTopLR
VJqI6Kyau6by7gublILMmliyb1rFIkGZcUMYeKbXvUTH4QYQgbug0AzqlRnt
io/+bnj3w4OIjpaLzrhtRpWBRztXQZyH8WT5crjLeikdF1aqrpL05BahrQlf
KiTyXXXuOhqrj6OMcAt70W2JpEGiRpkRYb/n0Qe7llPhFCkSCoyB6U1t4cFP
e+W8j4KQDtqNVj72M52fZq0eYLJJ8LFtinxzSM5ofRod2Xvf+Bw7nkTaU5Fx
8hC4F0WM4OoHzdOh3OI41s9e4Em6RQH0r2Mbs3ATfqnhtaVSr6j6QaFm+3xA
O8WV0D8s5RAqLP2AstNF7yjvXB1Sp5LEiRq2owlTn8h5bNnQelBItEin9f4m
A7F6tq0IQJ3P0e01fRNfTrlEyZ8/iqc/+7E0HuyQwIihMMt1FHCT0FJF+ozH
lHH5Hpfw66/IV1YWLJWZE7Cq3M10p8S6pifEhTrws+zQ03CrMF/U6hOyeJ68
cDucuT5cKXO7o94Z5d+x0yMe9CF2It7rgeMa5CVLVzgTWWc9sSbbM8nI/5ks
aLYAqA2RQoUqspvaDsCBVEjSwd+coAC3WknX08rxJ66Tjq65CMnl5S7j22/W
198SlgDf6KOWOwlHmT3dgBpW6UCaHpiGGoT+FoXTSZ8cWwd6+bR/fXDCF/71
Btgo6Zx2gCtd5TVTN6+UBpgQwAzYbbhdcU0FvEvjHpSV8fM7nz/60YEFCVG0
LRy36OKH1mGmXSF8ypysQEgjXfR06lyiEnadlDkz9g1IrLcUYr8I9qFeBdTj
m1ff+Wg9EH2oENTn6tkRegHVm576yoz+6sZH++e4I0+wnCH62w3NJwo1DjHX
WSO4u6uNSZlNHdXW2OvBEHJ+O+CUIX+rUbHbgHSOI9HURhbKKzPyxCFBoHvI
erUDrqyu88TlfQAey+WvkQcEZV+2elO+Mg2rGA+3bjIK4yFWDEO2J/CuXXkT
EsJZNaycbmBzcc54RZQiSIh1KCBreOjgm3hcYtJ7Lv0xL9rHHN5nQc/bTScQ
99EmrAWOFOBUhjQbLZPW5mko0MumkSI0ndSidt4MrLHGnABB2neqsbEF9VOH
hQ4ss4TggrP7iZvaWkt6UuD+pc8LCLcg1KDLMeD0yYfqjuaiTPRx6CUKW1BG
BwUhvOY7K7O5EBjQjtZh8Uvf2gzmKAXx6wv5B81m3ybkGFJUovQ4oTX5BXkr
8H9BBVzsDdTHuztbythn0wxDzhzVL7ItrjzWSvMMTiHvO4OEJmj6r6moaLlT
RwvoBP0tq7+aas7+EL3rHdiq4xZTLGwDOPQqZpOQ8mZxBgbQBb9JD8mHyzgV
ZEWMfqAcARG+GDeBO+TRswjkQqPHYsfczqYX83SNN1tBd8j3jCma4/iSjIYz
qVevAA1dxVQbEzDCk0oi26Hc8umxWq+me8WRrdxcJ1hhhX8eIEHbiQ4nXGnB
L3Wr8V2kfqzfi7zCv6GShZX73pQ3zTLWJvgjyWbNLCiKa+60PsyTQq/H9koj
Qj40MxCtSSyupo9tsbxsO5ix20oDBSTIcFy7YCCXZiscGXX7XItRuE7AKtQ3
E/3liXwI292yNpit46y7iafgZ7WsGgHn+XSG15Gdfu61Dt0sm36tpy5dVSLC
4kOanCRrdYNZuGoBVcvKxueSkkWDPJ9+f7bW5vZqDjlHuLVK2F7VegyPYqEL
QKk6RRLT3CcjIdzM9Yzj0wdxhdnH9SD3658yaZBHl2U0M7hZSM1jjZDB7c2y
5jO9N1JuEjsLamovCeGF2ZI8Pwo8GY9h4mY73hTAIrc4Zbm+Rv3bRRJkaBZb
1yMs1bRP7PG4ByLYDgOHBu9u293ZRetAuu6cb7sggpR5cxsx520TqSQJ7apH
VwrlhsWsgPYqI/DpISwtUjAEfxxUkA3shU21Ml908j5USEhnjJEbcQLytIV/
jmf2b9fyn92H0FGBoovsKnqP2SqPdTTRU31B74kBYqWY7sabPnVzVHNAVs8O
w5Cv+/n0t3h8MNeQl9P71GyuCOySgmc2dcwFFAGavPH+ZiOMceM/xRotg+nl
iKONQ7UlCzq8+QLbRVaMiLN9SlZuxDLIuqS4RxHqg7EfwcNnDDACLRuMJBlp
zUM4zgMiSdeb8Zoa98ltOp8iGt3uwCrU+Ts/1kB8VPj7JtcqdCwxnJxV7okg
HgZhZ8mGBoCcMNGriXvBAMEpLkuhtsLKMj0IOviTIhZqvWfPSCY9/esRAWfs
7ztiKysGlsHvWs9TUtoXbvn9HP86pxFkF30iSOnpiUNWjZeoPK9OhQ6b/as3
ryiPqCdPTGOuv5tW73m78zwbiANFa4N0LiMDQolHe1GSyeJJSUqoLCqGJvkt
R0G9fSn9ckE3+MXsIhuJwNn7c9Wy1P/NQCMAOwUIAaI7wc1H58p5gv7/9svP
qycjUwVOlXIh33LAYUasvAsNJmwyKhpOUIMtGkntRObKBmLp6XbYq8GwpRDU
Q5t0Ip2a5sClHRVimkgvfgyBQzybJk+usi6dwMhLiV+FKqg3K7PqzvUTw6CZ
2JRC7H/yIqudOkEfrA9teKi3LeOBPMMQf1FKBBoPB5/RBsQdV/eV6+1ab2nM
2fDGNm8olV1Q0RBWFJoAnLXxRRLUf/Z434Bmsi69wikyGM2w4vFZOOm7qRk/
9Df+9yi5wg9fKxfEL/fY4odgnI/9lSFpFTrVVwjnURIDG4VD6y23BP8HYJwf
94kaAgSXIcohF5NSdFaOWMV4OYGL9v3p0j6lBMdjv3jNtT19DKxR2qhF7BxU
KnGqkTXuSkQQmrPhms14cq1uH3r7NaGEDEKWsNTNsV7jUfeEEwhm913jLfpP
d4Eb1YLPRi6WkPV9/FUOZAEnnxWT1IPhvMTbJTJolBhR7lO03uXS4pghT8M+
YdgOCU/6CnIAZSo/VFJxUBGgK6vIiKn9wnGCXhDXOfPFYace5nhd1Tn6ZAKt
dkslf79hEE2lPK7Lut24ikTRYvbHu7pq8TjozxuiOH8eeXZlUzl6cAkQetAt
cxm2SGKcG56aMBqnEKsOs2cRh3I8pb3zm9BM78vUU80tjLusB4Lkyuf8SuAg
DjNo47l2uXr/iS0twwdkS7QFghAH3Nk+nw/0GkiDZQ3l3Rbu/By0mKvs8EEc
0w6jZyNkgCWU6xmpcdCwd99Subyz5zI9iADQsAFfnxt8QIcteg0ALbHhC2kK
TpFlaOXJBPAvGfZ9pdlQbupcF1+vQNgMNFe5O5jtTWQruYdmacCWSj4Jwmtl
CXSWNrJvio4dbZPbN2B7w6HOOCBs05EfbJL+XI15TxCUT5No+sAXfyijjg2v
4zMxvx9HKUifcJUq3PKBUTawB5bpT4uhkUM9nbnclh343nU9XnizJGqXz6rQ
ybuwEVaFhUYmMs3QfkwpaAz2849JEOX5Kk6nTksdm8qeeDJ2rPHzSSTaDT+1
KhPvT6edJ+bSSyeqGjVSGhT7n0HeiJMHIJdvWpw0cdmejM9wCEYphi4emH/f
q0jG3Zhv9IsY0LazTgrSltuYh5MBkgwvnFzP9pdkdZdEIRiSuTHak6Zm8bS+
bxnTQ+Lcl3zVxRf2SyneZCvwdI/i77cDvouWOIlEKXxgbzd+706xijDNn3wd
957Ty5TsUpwDKesYFnipiANkbijjBDpHVE7s6qgz75y6jMpOdDr9HAh2ftzB
/eaEX1C/22sD0YzoV5WQ6OndqrdlyZOqiJ0whRL1iq/21kKjOK5w6Pmmc0s/
W4Z0qP4dI/1s/fQ1d3StnVkQj5xNPsqJxHXDVUOFQSi6pobtTB52xsrfcRaH
XQOlutt5toM14GCj5d8m7HIkmjX2MfpHawb5m7aGbQgWUFp8tSPGt4ZCtkT+
OziGOj1CO3b/qPgMLQmvakN6eY08RsJWeJ6y0em4l86T639e7UxsacDrU+Pz
OkxhXPQQm3F6NdYOUbnccM/JV/Nf4rXco+d3KltPpeX25YtYoVFRlHXheYXK
XnqZ6iIIKMXca91qNFfMqnChuNRFPbaSko5SnAKKLk030c4yBdCGvRXumY0Y
iHmXrFu2+Kqxn74e5cn9zXorH9xkx8rcDrr+2GnJI7SVizp2UtDPbnEDpgmC
zPfzzwers/RKUggPLv2X9uJT8PQfvzMib/zY3qOX0LIJ44sk3S+MVdtxNsYQ
8qmDASZJCQoansSob2TAwuC3q8or+TJJWE8W5Y7YacfrmiXkYjoWnmfh+xkT
xhwFTzuesf9klto67ZNDJNO3YRRb9oDryABjgd8OSHY0l1Lgu8HG6GFz3hEd
uwZLlGfkM9k/cZeCGB159xiqQ1RT+w9qwMFbAtB4xfEWVV6lq0RAl2kcNTvA
E6mYHHnvrem9YxaCcPnKZyneJ9IRbSEnszGSSK9UivEPZxKFiLkdFIV1eDTz
OXYekpFADi/pu9UHDFYE0UZYoRgmqPN0JUgZ73FVH1RkjoyDV0LJsUNUwyqi
cUKtUfUqfyNXy0cKdBF+zy7aLWWF0UPwn3dH9GWvWivZ9mcME4MSMbsidHwM
Y34ddcT4uLpW5nhpvdoLEJ16/qdDEfqkZy3foOrQps8P1DOHxg/coScAMZRp
mfjYemL6KDo95l7kp4oY+CwVZ94rjCMeu9c6i/CSR0oIKgNeLOf/ghBUsfG4
dsWOgTIZktN3roDR/+vKurR+VKUQ9atJqtq3OQLtKsA5h1fQFoCN1/rUdA1Q
8S8eL4RXE/rbA6N170eCXXvw78+5ZemW3NDI9le9H4jaH96S5JX2S1kK3a1K
OlxfwmTXJxR1HSTPPS4Imbnij29UvYiGs8lUwA5kV5O1E7dEP7+2n1H63etp
DWEbsvk5TvdsUYAgPIsFILaNzTFu4lEbmv3b8qnW67Gb28dcgQOcSvA5TeZs
A2Tn/wTKcwLinAZInH/oXKjjW0gpP1zh59QBvf5zm8zILnKeU20fyG3t3nl5
7Fa8Tup0CdoiVRaj2t/oTam+t9T5KRdn/yIrbYNPExzesPCdtOB6grPAj4+j
9MYOTjoSb+1+oNfBRjjDbLcKHyAjGO6wTU05WO1os9zQvWFUVQ8GNIG2SQ3m
qM0LAL6svcm08/bbNaKdVv5VH6VNJmJdNaBR5GC0VBMofvn+4Ik7ZcwRI6fk
LbVCw+PU586vm+fKKi6erav5xdi034ifDhj8q1WvsflYDifTgwpQLPoYN11P
1znlHClJJHbiHNV7vxgMklwYlnNsDg9LsKjDZfJpDhh+GpjW2WftbPOJEn/v
5FBSIW1rn/Fyf753j0Axbp6SJR7v8TxSAw8oWoJA6iRzG6hq25c3kj/FBcxg
Cy0ZLVZXE/WAzVnJpCBzyvp6gjbACIO+oZNZx1txnxUtz3WGfRkwnoOHIRET
+hB6NB8FrRNqR8tHhAN55Xr84QHen5EIqUn2/KqVNQanZnL3xaTDS8vnfKgn
WLHtZatwxmfCp/Dif1rciqici1lNvk6zddwnoc2CyN6BrHlwgQl+eULhHrR2
JCPiyVCjidiSD0OHYCdof4vKMCLyUDo83F0oNrDrRhQ3438hnYcUu9D7xomi
kZMeJ9fp6ZqILghxQTHsMryJXazPlpR+/W+QvsvZKqLDAnEOapcY49ZOYff3
aDBfh6x2KHecriTzvT+Jw31XcupZQAWouSyVPG+Pq/uoxUtfnEkWfiL4loV1
SGnCNxXlnI/Sk+96Ux0ZQeA9yQ2lbNweePkpOV2WPEL/oi4a/ZW7WCj1hUMs
4ghw6UQln1oNqZz6JcGloZKuFddpQjA9KA+Y+qZFuE1SryGL7tob8qorRXUS
l9P5yuxDQMYdZMaDL0fkIcBPoYqf6BB+xiyiEeriE1WI0zcW+yXW6xdv95gl
jvEU8jjW/EJxtp1+2ecR8B8Y6zo2lPhRrYaqvcNtUCZOvE2nD3MCLOAiaX++
w7Df/ngBzB8gF1+/asMEgv/4j8f/nDzrHP7uJ2BMAJQC7X5D2gUkcnXZEfNe
970l46ZXLg3cZ95x0j/5L0CX5/+dFI5YxqfRZBP1Ka0fHLA0C/MdXZA6nY3d
hJEH5/VZoU/KH3mKT44n1ioiz7zC+AYZtnnxg538SHfZHGyVpsPIMCCiVbb/
jLJHY+kECPaLkvpZSJz9O6hmopb3gSSiHISsa9ZbFe5lbDDT765KJGUZgyCh
nOvcXS0I/JtLjO79H93IqkqSwdTbTg0shmsmHdQh7J8MW4DfGh6z9nSBsHGR
/jZ+FTEtFTlLMnHnbuJAj+xaX0u6WWTbVZKdzVfCbfVbVkuTWX50+ucuGOyL
L5LfaxekA/6Qw5dUtrxJr2UvhJR+aMhskg22fJQhWrbXcJPdnXB6bcgTRYUg
B/oq6VIZFFvk2Ugyfid1C761XuSoiW4xn0F7M343OLrimkF0oSURm5rAyzGr
Jiv1NpYL1q6BVGWeWzLsH+YtjZ8KGEWFE2Id846qaxwVFQu00/HoJbQJ3Ny0
a+zi/2/RJzScwSpMU5+gai3ohadkTRjvTahYNDwjwLyzNnBXMr8EG0Z1YAn4
nTWq88sx+vNfhqtS+gBLnxxj0blH3J8t+VKpWwdi2BKwy4AJKAsFmObEdAea
b07jxWctzK9EI4g7GJU42k4Tmfly7z+RPaIyuL49rX7que4yT2nhB9zv/eXQ
HrRZRl2QffjqCaraWswt8zQpXL9G++ZRBr3I7gC4IOsU3Krl+EGyZABLe3zH
etYyugZN8wyEqxcxin1y5icpd7zOPQ7gfHJMvAwzpcanG92ofwl9tGSjImSi
56D7m6ZtgQ/zfYp0ali+xcNJPu5solSuhakJ/Y3ZjwOoyjYGvchbZbBB41Fz
5FrPhKd0XDI6RnsO1spsVG2go7Zy2RsD8v+sj7s9uu/OcYD5yQ99nBKdLcho
oPukRf3VsdQAWO1DrJseKlFeO2UhEIGm18JFXcHI1Xr+2sZ60UDHXQ14wCJK
oCPoiTlukOoe9GWaevqRb9FAMonN/zRDhXbcyQJKoLV/jXNvvNSev4pY31pf
T6cFj8+iwm4KYoXzgj0A+pw+Jg4BwoVFgK2XapxRcuoJj8N0m9PYKXx+7jnC
ldK8dZ8bzhLPe168uOzownssV8cnuAoiQTUFS1x7JAKgH1iTaiQxnKK/vofD
k6pi2LdDNIpi7G6jtO2prPmrhkuBY/E0nvZune62u+prRhnZMxJ0AghdrwUw
M/s5so4O+gPZIoY4joWpPOFbtW8J0Xnuy4crrAtF7zwA+5ACphllqESQKy+a
xCKkfPLyEGtsS3MxaQxNMEJ7GcKF2A/kxil9bAX4fIUTv9SHD8Ge7mjxnDyw
c2cp+a2GjwOcqhrtk+IyumqUqsP0JVcXPwGD0E7cuBg3Et2wTUHvfoaLWerl
j/sb2KednbCWN9jSbthp3D99JGZtfDOynLPptCtQVe+GTRkhS8a7FzZBsABP
jXN7VReC03gkmuqjpDAxoHC0BVBa7V9J/7/ix4X0zi18+WX0OXIAJJXb1kl1
/pVBaeK1W49SwgFbDltd0SfL46oxXCPIDQX2OkukauRxqQN1gjce9+L8MPKe
KaLEsUf7v8UkuN12jAFlm2Irem9/5/3Z5Q88Pg9ao4b4BPfwaUftaUK7+/tr
mkqSEqOInvoDS2FWnra19X6KHfMJa4a834954K3qYBgBamN6zFL/aOTSuhTq
47q8cOlCGykY+RCUqrX4KFl5wHBkqdTOAD4Yc5WHNpoXgRk/hO23B2Lf10/+
fJsmkOnPWL/pwcahcXCQ7PsVjXhvVuDn18NzD6KHS6YoPyBhI0XHx8C0bGou
L4KV99YzMFkfxZcSit6onuQLHGVJhWJBxNIJgVarherrjS9Tz8ubFRG4kUfq
9K4IeUqTd+HpVueEAcKeXA2bIpBf3wVBhQSbhDZjj3WG7DvanltK4ZQTyAm+
XRQMzNEMxTR+4lWOJm0LGpoQpitBpNiyJ22v1JX+0+6R8o3hp5ilK6qGz4/b
/MMMCh1eCgUmCUcMkP6ER2poTXGVz+KGdwd4RE5OSOlvCFU/26U5l5WBTrzh
buLwzeswx4D2FoTqxFakiL8cSeBvSOHXYSDIyakDwhowIeYqTvCYp9/Yz+4l
xdO/eZXwl5YO50tVVbGsm8QOGxH9iYcuiDqlaMjutTkNlpNAHEqeeW14xSKu
1NFemp80epBPcinhQE5uiIHVTqLrJ8S2UDvnLFSAQ4XBcR2fsQYbnAZH3Vwt
KfVFwj9+IjxZ3MvXAAWA0GF6fNtgAGUjm79t6654VCm+L9pGmp+Bb84Bh1kY
QH3IaC24GPioeDXHu+MQxqX8nuGh4OQgDY0QBuwDKDoVzk/bonumyKs5c+oI
uk36aghnwp0z08TA/R81BsbhcUxkcoyH8dgh+CowjVTOL2AL11PQiOC2zIER
eMLjugS5kidBwb802jyooOF+WsSBT+Vm4w1TdT91Un/1dCqYroodK+xebpso
isorbLlRtIB7tvbviJEv25Co4HnMFnNSMTfG9DrEbT5hD6Wm5NLa7reXd0tb
Y3BGsoaobwp2P7ehWgo6XXny6fHOrnFWFzjar7uXuqq38rIT6+qTVgKF0igp
EoQB3m9XZ/He0CftaFaygaDqDH35yshpJnInGHbyPNeMAAQnGoA7ZflGDDfD
CPcHFF+pT5om5jWdmLrqPC2S9eCuthh0mDFwuAXI28orT0r+NsaVvtDPnU/o
d4WvVzlKNohEXtMDG9Wms/R27aZHea2zmD/2nNXKgKHpnrgpZBilYFviUa9D
JEZJU8ac2n8DgDFVtHz1y8Oz+TXkSxStEdNQWjcvfUs0cUpuipnRIXqnemqC
Lh9eyB8sQIkYDl62Sxoi5BghMadT9HAGrYamlKHvP1cDOz7iFTuIZ3Gp6seN
0YN8Y4Bk9P/COwQdZF8e+nCcTtH+pgzIz+A1UgT7a+kM+90cga1aYgI2/1wu
ZvRNMW4C3WuUxcn5eVEuNouDMJYZ6mRC7IDe6gxQMFdBLrr2ZmRgFkQl1Alx
9hxcimzFjUZSnhX9WvR9QsCKW3GTZoiehAMyXwjASX8QvpltQtE4pBfQCqlc
FY5NDml3PBu5g2Cse4781BryvPehBeGgZPByyTzDB768emW+eYencrBErlxn
BdZUZa0czuqWcFqmSLB5i3tYqL9d3fFK88Rf6ZEKUVcqVya16oYaDx804Bht
UmwQb8ovDqH/nzRK75QKBLWGYwWVSFFOYgbSOKaQOJHca4j+aL1o4w851TEV
Dp0KqdUepbnT4NOXbfKFFywZ5HEAg7SenFnIyfnKz+BTz24dWa0voEPKuf0s
29lA+j5L3xpDAns4K/f8ql1Be5tisuWZRFBK6/+TFmIzZCZYLUcH8W9XYkGe
c6sAWblQmnwK2siXkWsIweU47r4VmgH4nipyw6t5mxEn+VE9WH6JCZgtDe0l
O3xRCdpK9wqLAYGFRyKZijBNujljqtW3oUy5pfgZyJ64fRtvhG29hFwkenL8
3l0fVqzRCasnl1HO/uBOcU6obnqDxCpd1IaLCHo+PFDjHEeDrex6Gtvu17dh
abQ5jDCaXz0YuKJFD83GxDmuY8bmRbG3mHmmPXPIF9gmW54S8c1B7joDv5x4
ok0Iy9wwwkqWRIz+jzIghChYh+Hp+V4R9eo+/Z8Tb0nwqV6CbLIp8DTUgwR1
pfdPJDcc6GqNgWnWTdoHYl31kZ12HSdoMam7qpZbmDOIXRgD5wabXSgt18jv
OGuaWY36wOMrZSQ0ucfLN/X3JQx2PNTI2VWo+pqRW9eu0mzrJgEdA8+Z2eQf
B0UHwH1pjaOgpPdwLECUUnEE4uURC+VU32UMEjLOeRttozryv4Llb5KpD6yn
GzNbwSSxWi5yp6WlzQsRjvQR01mw2NB25eEIBeaJygBvAQFYsPQ4Woc7Ipue
IawMwX1dmVt4Z8dlz76QUyu+Uq1lZghQyrF3CAnHtCEzN7YljaK+Ntno/YYE
TZ0XbRy6RUnSniZZbFUtyS+R/V1v6gqkaBKqY31zLCxainJx1nQe9/frtYrd
fjFOJ4kDH2GByzP6PshXvjp731Ofjhzq3GUo/aC8wQ+YU22kAoKkIT7Wcf9c
233+k+mZ3uN2hqlCIR9y56zBvIkGa5gs/rFwAkPBnLuclBr0CIaLsHzkxcyr
Da6lpq0eWDBgY7LtxYiZZoMwl3T+HLff25UeotafOBxKuhieu96y5jHxzPab
f6uQDKkbnl6EODuhAenMgXk2UTSIuez6UhyjuzbKGbCjbYq0DBvfXAxSSVnD
t+2Xw20s/ICHK0rj7ba6k4q45P2Gqauvh1R1qwunan2pGcMs64PcADGLnt/y
1bj1aS6UgoFlp6y1kl5Emw1O7i9w1e5sXEA/TUfdA37ig09y4y5jNF87ELUW
Xv1ZDg/9XqcGWQpltacSZ/ACtRWFbqWekK2pGpu9mRAC2Fgh8qOqKo55h3dl
6nRstWqAxZqiAUQ5Nv4BPp412cprakhY4vSymHfNcvlK91NAyUCdYMuf1w3s
vMnecUXDUn31YZc74k+0ijNnT5AdRGoqad2/VodBAEmbyHm3tpwfMFSICG3v
YfRnlPZSjWFerwL6Fwf2XVb14xINpwmGisE+uqaY1ORdQizOskVaRzAPSC8a
SlhTiVGjB9BxHnTxogvRbg1bv0Jor3HE/P4X7K9QSjsmiqHhMnH4QSuOUNHz
7uU5MyS++TUZc7yvRUFVuxb8Hs8bcRXaYpx4rLWkQIr+d4+R8o+lny+q8RrG
BGU7eOfKt6hIBnKReJYnsDOsqcuPsQ3B4fGTGnGQryV4DZm+M0n5jZO3rDYG
KHgsBZsnd68dtRQyXfQFK1kP01m6sk3Ms/ZN95klCK1szBDLvfrwoe2KTo4d
kSNfZP2VKQxYTvxF8o9h8/Wj6fr6neZ/00F6E0TCrYUFO9dSVysK66dNzlqh
8AtKhAbkiUy7e2F1d7ZumQXykNhks+A/PJQkj6TmjVziFvD959dYahq0lua1
Gg4J++otY0EmWhOVhI6V1sYYVT5t/x6rBF3qwkROazK35NPhieLNT70ycvAR
mIA4Q90JCXptatMAQkxHf49jen53mv6rR7Rh/4xR6R7SFxztlEYPvdW/YeRt
WPD3q3nDQ2DC6EEPP5FmeIBZAutx49nsWZgS5wp4O9++kkGaHv1NzOj1Xr82
rKbykQB7OnjVykviw1VbvaLWUPWYdZGdIRxu9smnzeKmXbt4YjyOCCrzFfcH
Bl27aS6FgoXYULRysWSC1zK5CPjvRtAfD6peEAne8usaavFxL2lC8I0/M/Pd
WohNs5oUzUaABs6Ph2AmTwzaXhXVdwjhY7qFP1B1LKpCE6g5S7XVg3vBrWJZ
ksctcVxeGJvjcZhWmW4oWzGMug7E+vsgsBrfwntIzWRFUl5ob0apY1YIver7
PMNgxaf5DIrrUomi47UrqU0KOtV5U+a0jUx3zOG9n6LMmDeCP2/t7Trw1YWH
O9DwSbqM+sP6H67F8zGYvWK09FFuZg5EliI4+miqWxVw6TzjyYr+eBgAqgPD
CWCDaYtwU6drVo8DsvYKr4Mz5aunhXVL5NK4mzGQZ7zMnGoAoFVKul/zNfS3
wP/vO7FavVpMbSJeroovpcgTY1/NuG+t35H1qVgIyGJDNYgq+zigMQCr6iBW
vqNCqFwjz8dqTpaCaxFTFF2tVX6uSzU759unQudRv+3jb5ORBYHqjUE6nTVm
kQINk/61pX4xphSvIej2WhwfwuVjk3WFTzEr5pTTbWdHpunq41uS4qOs3DWM
2aaIHdmq1ZWkE3RdgxpbyVITuZufKzZBCn+XEnz5U1o8JNU2jf1ajdlLH5M6
zX5Trt1P3kCc5viAME9Kk+/ez9EHhaskGXj8JJ3UwHs91MPiYiA6vmv2lAI6
f9HaXNyXsq3KxAja8z3PeyXpQ9aaGRpUsZtCD1j1nU8VIiwkafpsjkkfsXOp
wVGnapUXCBZHyI70B0fnKUzi39WKaW6yNQ4t9PzSB3m0ihmHHWL8LHh4E8qe
ZjJ2r400Lws5bu3jlu0esH/134sX3OkeGpe0lrel4oejqOvTTrCVmCQZZN0y
+8WR9l01LWb8zyzN17xpnopX0PlpvjwZ1GVZP5FNZF84JNj6aNQ6Pzhzh0eQ
zUPq/DXAXnSYZ0ejvTO9BoOghzbZMyaNCWlCcbq0NMfYfnOorEtXD7dYj80C
xMVB2g6DGMS2Mf/3AYmr8xn9K8LOivSsMmieBb7T4M56ixUWLpcPxv1bBzUA
xfegY8egUhmf9mmpPQ87Qx9jCMJV9IJnm0ADWkqaYsP7ZpYwHk8jCH5/Rgxq
sqDIKL2LvClXccnUXZ7949IDOM+xBJtKEuJLdAPtrFtUo4hT02+uoLal/zhY
XQ1vONarloMyhN/pnAo41+Ism1igKjQ4z3hl4+mUw3Xx1mVWJ/HAI+TDjs1T
eOrnNKzUBgxUIHewrivtJRvns1W52Igf2u7CM+rMVD9itu5AhBBPfF8nN7xe
MFimb52fPY8fcGVSnSz8hIphCsTexWPnZtFEMKbVCRwJsFNusVEYU0tzjBFD
dRwF8AE1T3N+BOK69JGOzQuLyUQWIQWauoQYFyQrd91bg8LvWyPSxGW1iufz
Jn5V92PDaoeelBXqyDRjNBwDV6ivowtbeZ6oovwZ1kHePHPyQYzwG1XRlppa
lSFcra6q/tp54IAv8gnCNcrMbkQtSvvvSVPUCIwACSW8ckxjxhsUFwB6euM6
tM4obCo8Oe7a8ItSgFXBBYof07bc5o/pOdIUAhGTpA9eBfDLNmpUeLfwOkYk
VphxnRxPzt5wT0DF1ULJfOnBsLqQBvs5SoDM8mgYuvzYMQ3YfSHkYcZ8mEwL
Ew6KLl3uLowiJWaLJnHOchxVBUTEZltYNoIRkmVw4PxVgHwc0kNNmAYx8oYR
sCdpHdjtbmyW6kOUzO1sZPCV/rFc5qbuSw08pDbGMhOBDYOBNV7K6Fyuh52x
Zv6FawPSFLTG17glZWTmJVkkk5nL/p6Apc9EnWBRE3C70N5/ief7kWqwQW4J
SxcGt3us+2uad4rxv879McjdgKWxL17juIdkpzA/+gxnfFYgp28pD0xgWiJx
dmQi854fC0uGAAj2rj8nd0kQsdz/udQwDiXR1e1KMIkNaOdWPggiSaMiyecy
cZqTfe/+bkHcBIA5PzVP2SNaQN4ufvnUl2dCxHQKxwLcr1DizI2VfrV+vZXK
n9Zko+F/nJloNfYlmrQkX+GU2wcHPFvkMXNejZDyWJtEoQdlRLYLGyt3fdPZ
qLhHBxPc7AnjVXMsvgpQLexnzTgH3j7LWI5Kuz6q72aQerQb+MTf307f2zUu
xhFk0+Y3DfaWnOvkmotuSdSjs1jV7EFASyRdIs2DXgQATky8dA/JEpoY5GcD
Yri3N3WD2ZjAvXRL+W3d1glabAQr5n2Uz7EWOfJtJClcwQd1yMOQ86VysKdj
r+iHTGG10XOMlB7WDr2SWLF7UC+JLcmmAKmkcDYWQfwGDk1RORrhwNn0HVmB
vwWf9b1GrgoHpaYL0DoJ8DBWikyxuxs44FRGxp83awQQNWx60Q74CuIw9Cm/
LN8JObdG35d9xe3tez4s5wd1OMutz/HMPv5m1aiBn0SEFUNA4GJGkYHkOmSX
rKCVqs8iePn3LCu/HxkVDDNj4s7p1m9Ps7Ub/9obIdSCHc8RGQ/6kc6rRdbA
ivLD4hzW+OETvQnpJ1fT2pT9ONrgG6VUAtM0gkRSjuGbWhe7a/0fXPvCzjPX
CGebRznNnNWKnlknkbWWucVM2Eg4pX6lSOykFqys5chLeTKVsn0M7Mf9eeNp
4hiyE7wTI0qpxEtPEtnmZ65MbSArIzJjZg4McNw3QAcpr/J/nFZJQ6cA6KnK
2Pq3WTcQaj7JQzwpc56/ftipVNLtPNxB6ovjJmFdjaLiZjQmSPAeRFEAev3C
vnQsuvO+CdT4FmebzCc12zAXwaiUIeKyUoHtA5xHC2m8ZUymQJSul2JbGuL8
szKfC0JbvsRN0Gsf5bm2kzGGYBmX9w9cf5dmmMWTgHa3txxhpoR3CMXeqclQ
KnS5wQtV3aPe1vgChWxYDaJGyg70a0Np+K8D+d5AB80/gVUTE7gNc4iFDMHt
tX5m7vxw47DxEQyXTFgZ/ujDl/sEwSkpUdyyb9auyPjnvAjLyahkg7jml9yB
Wt9cD5piSXOXVuPGXG9yF/GB9m7Io/JkMN3S8iNE89KSC/CDK96EAh2Id5zO
bn584y0YTNJfRhZ8Lc1gQZ5aHbIV3E2sR/rvo/dcZDCFH+Tx2xi+aLv6J8tJ
L3p/O4fyE6SJIOaSpVFCsK4xr4vOj7mP9hw+cG1E+l8RW7S+QDODLFdT27JG
oMp+q2QwkZykNK4cXSd05QzeskwKV5nLJxjpxEhQZEGMEcqyTiD0Sv8sBNnA
jTTn4G5Ee7cxV2h/7FPJA5N6Frk+8zJwDvF9tpl50e0Sc4VqiVv87F4XORTX
/ozjkf/fl7rECP9wVbWXqQZeI4/ilifmlqCUeIdOiYcIYstjAGnTmFVL50ba
4qsghrb1oG6E04LPktPgDdcjgaKvH6RkspCQ+Ckieo7DNGDv/dyB+sg/6Pd2
oN/uopEnYNlURBiwnzrY6/gAidZq3WlPdrvtzPijyW0f60kObg820oRDdINp
0CAj9aO3ZrlkzkL51+Yj85kokfDMQ24LckrsYN9abIgm5eiiI+9ThVB2OAs4
uMaYkXVRMOsXiokdzykH2cPnMLmCiUFgs/Ks1iwwnHXoxxUqBU77v6yTjHd+
eI8zNmQQYm9dDQW2zi+tlBphz5uHyGhRVAh810kFZk/i2IuUvrowU3MdbOcY
lN+EHZHorSPjGMcv5VlmGa2thrndlK42Ef6WQdtHJC87IU1eD1v9LOGNYZut
RFYGdly7iVnq1naXvI4yZJukjZOTnfIoLOs2ziMlv2LcNvCNiInkzuzDKDGB
qMNKtAVC/Z+gfP1DeXNucMG53bnIxcKsgwFuhtYcgvLp89JdtLx5e1ca7J+W
Wtoa1JRmAlJkh0UVBGIvyNO5LVdzF9LuKJ/H8QyfJYp9TLDWdRk+7kQmorVy
zf19NQKs9glTfJLbp+bHBRSWi2HevA5s3TTC9mrV5CGGuYxnUobnFYrdo7ts
+7+70lVa2UrGH06lWJsFqJ/sv+1dpXHRat7RV02pSefJZyMSC092jYnqUwa4
DNzhUrD7sPoEGJ/iFbWgZoYO9DzWBFUiFbaFAj9sB700UrluIwARxTnUPFkw
skQi4U0dx0TH2PNqipIwGkkx3DFGyTHfhy2BPlpG6fHFIQl87JilCPNqYmn2
X7c9NGy9TOdMZwD7y3XVbQbW2lG9boSB3AHiMtFwGWKjC0EQBD0ZvCGX6M9G
z/Ou2E6e2ufSe6lc+JYlhF4/CPPdJVath23SamVmJASoMcZlB/44/BkEjXq7
G/p1WJljxzIo5/ujUBdof6RujE4o5dCtaK6B2AmOsCtoXNCSrJ+1R23CN9m/
KgOUdcExI59bp1I563/VCtbIqJfI6y3RKylPqVJ3tFsOgCiyCpQUgkyCsPZ5
RDjOmIIKYBbz5i9hj4rNAsXYtGyYxvAFx8TEo4oocWgpUBrEQIjDGk8EhFs4
7xwfSY6GP8Ky5Q5tOjQFpbrCoTg5C13qGPYMcl10w+SnKpKmg1C9pXK0Dmj1
jKhAch/d4XBqy5erCWU5aWEy4DetAevnYFROy9nbPP/ITRO6+zTF0qR7WTr/
Grnza+3F4i3llVrz6AbeS4C47sFl7mdiofjh3ZxYbclVn6VIxpLF+unReFFE
KoRj5z8xfQsWFPyALAe60tWsdggMjGbN0ssmlkHsAfVKTQtwPkOXn2EWik/c
hvRAV6oRiV/H5GHIfVu4d2ygfqo0OTxwG75qYfj6OG16HMxRAQlQPWCAfkE2
Ks+yYFXuEWI97CKY2d9tSvQVGICreo1/PVO/zikKCyKVhJNl+AQiwdqJmwj1
6lc6k7BBPHlGeFM9jG7nHFJn9MoRZDi6qQ4ayxq7x1Rb3Mo/L4w15LNdlkMb
jxrUAkIBevKXiSSqO0U4tKv8aYATfLNPpQCQtJ/ujHTKP2/FAhwJkFPHmoAj
rVvQMVXyTh6xin/vEac0Or88L3qzQtbWQ+XTN8gxdXLTXOFQ5cq7Kq4lxL36
jBsE5I2VyqL5BDT3HOvNI+gd9h553Y+jhENg6QSkmdkxtc0pvHTujVIbotoD
621pdVBxBYOew7jcEFQBVLW9kaW8xTplq2A214fa96aUYgpT8FvYVfN9O3zU
ceFBFsYlhl1dlCbS3ia0cjmE48ZcKDb8Syuz2rQ8uI+eAwkOo1qVVo3yAevY
LmcLRuKBDYZ1Jgrcy762HML8QkIO3gOzFug7yXLvMvMIx/oOAqhyI40+K3VH
Y1PzSXcR9exih/QWLIuGCaPFcJ6lm8uzGRuxH+0FnGWhJzA0NY99Chh3sjXt
7yTfJ8Tiy5aV+21geIa8zamY2GIhlSMU/47cMBXtFuiFYMt/U0rCeZJEkExf
gvYsSDsA8eIq9hROIOrtGRDJ/d8SHaGcwO2COC0rGqjGhVk0Z7KyXWolc9d9
r4WVfn2HaUtat+tf7TPubnsB2qb/k+/X7JLLHgX60DWddPwHH5sfK2AmHqyE
AD8Fz8KWhKssEj+UsrglPFnD0Ys9acDFgDEj60jE4V65bDCS3uQ5ruN4GioT
Gc3EZN1EMSCabNs7iZ4FIlcW7cVvnXst2FIztNVxyI8UQr1DEh8JlmKhGsQa
szhlGtadaOlzp3efoO7T0TuSHspsx10w/M7d5/nAUHmGIW97DRuL4OhmzJjQ
vm0Z3cmSdxIwsOsZCm3jH4RtSlOIuhvfm3kX8j4ZbHf1gmJD5KHNvj1tiesV
pjkC+jklyRd4Rjaqj8bHs+XokwUdZTPuA1toPJYGf7RWEA/ZpF82UmrMQkaA
gWJhXbmuZJSu0S8tEyFOMYR0any6F7SNGhzBpUuntOkNCYlX6QLvmwrVmfbh
Bg+WLNymFVuGtgAzj0E09ZeCHlKu4Zvk8NbqoT2I7W8c0C7TCack5EuJ3D7K
0hnNLM5wDms+jhVwmLR5/oiEpU9Y3UJsgivyOg3v1HfOX9krw/qul5wRHHWZ
KrlQok6hhboMlg8UHFAO24GAXQIdsM6BIRCuEsQpJun3RjeBJ14ueBBvmqAU
6QV706Q3nFvwDMDSeY0ss9pF7I/Iv6zXDgGCXI4B1w19AwNvQR5RCAhH66ht
2S3GY6KPMS+Lj23N7Levsamqu3KCm76EqnzpNrEL+TxiJvuOD29LEQRZR+kc
BhBozKQPrGsUNRhJDyH+31Pz/Rgy77A35UwK2J1NucDpVMh0YukQnOAJ8JDm
37eFZV8lvpe/2Pbzx8I0KfJN5jETrA06YFv8Z7mhgXl5bHStNF5V4vPXB/4r
oBZsMow1Ov4z37FLk/btMQ3Yr+9DJIkQrmegfjEtv2Lp2ViyHWfkzImv3btc
DIz5Kh7513+7CvtXU07Ko+Iklac1suSYEBf8nC81FTOY8oTrExvaw1Ya812/
iMohY6hUwuPiuPSeX6LSj3r4OaVrTR/h65eFJJcWKlQMGn0zRCOSRajAThIH
eUIytIIekuyG6+sLof3XCJxNYq+0sKW21cbUIhqRi/ON14Ftt3vFCzsYusZf
jYr31SUsmNUrFQK4fvnt/zFIA9ZbIxrT9O98srwPr0YK4RZtJx8YZswPy7FL
s37qW1cxKDUib93TMeBHwHOgbZaK0iO3oVjc4azTtWutlf9Trd1yhdhHmBzU
4EvlwSwkWBhZ6NqbJeEGQtMkTUjgBJ5CbFiUEtkADvkHXYevrSwXVe3J/95V
mpJDnSiTG/cY9vwxUBqMR+wEnUV1oKyB3aA71yQrv/GDFemCuQQgE1Tqo6jf
fVN3/Fyvxsgr/Z9ri64StHlQb33znBRVnxoz7mlEfCef/8Yk/zjU/i3pzZUP
BnnUDeGTinzKdxUhhtSf2mkuf/n/fYGk+fCg24FJV6ajxmn1TkKIqpZTIQ12
FhFe94Fh14xAeNzy65Nan4LmuQTc4JQ6PJNX4P3dAMnhbmZh3pB53dla/F5r
aydkLEzBSjExYaENozyCgoCXjqY/qlgZPuq3iNezK12jpwqEbfv062GdXmBN
grMzpybdVo5gCAwpERt+SBaeDuhkNaf9YElAZkUYwK0117ffr8Vs4ABwHebT
udCMmaSLK5f6NdeUc8J3Wvq55LhQBS1kNnXQjgKXQ7pCy9QaOSKD/R3s+s2b
zDhQdojnA9XSFAX0eca/e0zWwmKS2T09gGT9HDtpPgs10uiI7W9SFemO29KI
ZOBcWn31+R3STa1bxJl0N4mYC3N5NxPWAPTQGVENkCyFH74NCOYwgcE+s6Px
zx/ol8Yj6MEfqQAVbdgIGSmjxKC9mhmvVrtG0W/TXU8m62aGd9h9dzk3q9LG
ds8iGSVwAi2nyf+ER/PQCu4OYaLrkoyXqTK65goDRr3GH74Nyr3/gi+O5V10
/d2g+Diyy8XPmvCrkHqHF6czDarD9lHbaVYOdk3MqYr6bT7HN/7FaF2vFoTY
uR1qJVDnejsPzBtXQXpTcZg/Ice8pm2VfXHTUzGdJ0l1rPbmP6SQ1DTvkPBv
g1mLttAG9eczVCOInsMF6i4XTchh3TDpbVfNBwhsHGDBexVmCgdVc8dDf2JW
c7fp3aCkVz64xzD7IEFeEPbxm3BGaJRy7mV3hRK5jY9969ytC3V2OhZd1dKz
+s6JtOuWG+jp3HUvENHvQZPR4CZ8tqgTXxRf8tH2g5VNzVWnqvOMawM/FpsA
x+NAfuW3PkXvEIXLaBO/YOO8l81iDGJTuGWm9fGSrfcLuXy37rGEeWuTb9RN
oWuggyThkbf8Djt7fXCL/xrXWmlXs5q1IW81FmCdsn53TcNntUK/ageuSQlz
+qMa8uVBKNCHiP4J8T8CCpVnxSxVu5WNMjTXCgZT1y1pFIGkgzKGwpI99rkJ
kzFaFfAor3hXLFriuxaxJPwgN+TNDaGem7eA8E5/JDJePnVzRpHi0oj4jW+2
hO0jyviVmX+TfgwtVALfzXfWlfxyDzCbiXohhJHkInEVuUO7YJPsY+FH9uMj
PFw8KXV0k/otQoHnLXaqsPSMulv1TLv9fE+SSaRlpodYB/+SpbAmFPwXUOrY
QQAU4yi4pKPhxDAtTYQ8l8KePXaeYrIKsXsPbjs+VWapTfKKaGHocVFuBx19
1s+8TM+mM0/vShyzM8X4hU+VDyxwNP5Y5T7l0wLPs6Uf1knjJlio9DuWCRjI
HIuaNKxVlMjXi8ii9TaI2PXwZJptOkvAMlBZILiERU7lrj1qIuvvEyNXuG/0
y1DWaDimnKIFNWPDk6fMj3jrgUT+NvCIsaGrFrGT6B/pWuZlEgXl/rKwkk80
dgFOpulqxwae/usYsZkpuW/7I1xVcTVfWwx3Us2AcPBxcBK79cYnsU2oy/U8
82awH335SQW8VQFUm2is6bCiY14JvpsgL78Ac7ZXIe7E4qqUDa8N/3PndP7V
4DAZhQeZ+5Zb8y888M8Z50/mT8GFul6NCJb0wL26b37Fb2edJ+tCuByzpEX5
87tYlHUSNMMrKx55HPesgoIGPWZOSX6lU6E0/PK8CuFeddLZFTs6mZSMWJUx
TCUjUe7oSK5i4XVNkQsYojSz452jNLkO9020WbwKNEpkMFL/rVjevC4JF+FZ
75ElrfqdNL89X+S2MHEGxgQYZk+KkRXbmaT69PWvF6Op6mNi/nwrw1rHH8BO
6WcjiNCKBn/JrC5nsaJ9NuxLSIh+qbXwaMHxOdLRyG15v2q76ZvnExZ47xbD
YoZc+vMKQRMXQ2Myu3n7I44ulnnsE4RHwz4BT0EPk7oQaPvI9AykqG7SnqSw
plzDf3PwVtvk+zwqp/EqVLePj2pxAJi23DHm9leTpOfc52c5FlXquQ9PUIon
rVvR1QJbqcTTfEOL0yiF5PcJn2MbfX2+jTtfSbm7zrUgHh4OLFaUrhZDe5bK
Wh2eykwdV3ANy6DZdtdhln5Ca2ozjAQ9tQdRwYzRbyh3UlMThWeI53dDZm/q
n+R+aNzbbgbnVx2VmAtE1w5A3k8wL83BqP2ZmrFfnYbo9FG43LGG2Aw/3Xt9
2Zr1VHOW3vVpdgUuoI6uAWkIp8CuQZg8lWmHPwzbbOWamC/Qw7p7eM/XM0m3
yHvj+YZnYivAXFlu7qL+teE+zhTRF0WAALqb75Fd9VWLStyRnqm5mLYxKVMP
pWR2baliGhr7ywrTL2zCEBjJhKAVPU0Kie4s1ehqJOGi8mKp4zfe2KpdVlWH
X1q3AS9OsBQ6jWS3nUcZiidbUGsqPTRC5XVWAA5QDd8ApwPRbKhYyBP6crwo
2a/nQbD6UuTohnGgQXkDDO6koTFwUnal6VH/sLos924tb+gILuhiY+sPxuQp
dwW/l9GYOUL+dQXlqHpL97IpPxS79s9/kzbhPQnjLdNGQldBtt5zcSVZ12xS
KxFvtpMKG62xNVoSKdjzp/oIqc0gIy/nfemi9zaee1FPXOVTWG1IbcEVKu3f
4E7qDm8KZXNOWxaE+KNaf7CWN7Hp4ZPjRmDaMz4OLrgH/WEko4wvZWjFIl9I
xr5efoxrWEgwXmky9najeyyICW/c4VVmW+MG0SEIsg41rLl0EC9ddbvBsnY0
I9T+pgbTuRsKlZqEKhDFQ5XYUpEO/hI4zvtpPeJZrQbSdFyCYd8ZPlxU7+hw
7zN68fOWMsreib7UFMdmwGiPtJlBC/K5YDGQKrv5Qc43Hvf3Hpi2xHd2ONLT
3uIFoHxfy2/dhVynovEyP7vpoyXXJyaGBVtDSKq+kP6orcPiJ++o5KUYfi6i
vVl0pXGhggjXYOZCFqkV3ie6PdLSSfPdKiuUmH7aqLh6GCNdRSlOdLtc750S
BpCM2g9CSQsdZnKe6e6mXsZacusNd8mmB/t6h6qbYD3dshnxgCEpqj0MKbLU
3I8+zSRs/lOsdboxZCx8QR9iFLfq93A0fCj9Cr8sXPP6+vPflBvCu4jpmV12
fZvYDq8vrjLsac7RAb9qKSE+zADthvo6EURYoLr59nnPJ3lZRd1KcSAG8q4T
oBMhcLdf7B1kLYimX4swXuuUIJSymMq8LP88py224qKWRiZfBgsMKqi+x7S+
zGyeYNbCGWMBjmte9te8JsNHc81eBCorj1VoDwa5IEmACjh/WKXygUzeRLoL
ugDRwqg/hCIU4HhdS3w0Jk66gx3sdGg2EVNUIWELpIVpHWcF3NJrlEWXP+ms
MuuSbIITdeV65YpDDueq4o1C9nKOnzkG5ekRBKPmrjZ/xVt14hH+OFd/ois5
ur18lGGvwXNdKwzKEz1n/h7d/aOfomMS/TC0KDHaunin+osdLC90b2zZ7kS5
AY5qNfLvNksy11CDzVt6JcYES+IHROAhXHr5Al/1r+X4mkTtomJ9KTDLsvEu
i8gjZ4LB4zCpCc+Sn8ddyT+7YIxysycqGil7B4uiUGI0RAJ5J+nI6WgpXmgv
3oAuxITzxB+2yAPDzDYJSffRX5p4N7vA4QOYtXTglrVC9MENJhInRtqQ8WM7
2YAn+fzsItIuYEmRYx+xICSeg3sKA7TXxjx5kV5+1b+WR4AB6EQmyNWpN5Y1
gbIu4hFUEknIrUvzLI3BQDC+PNdf1VdOtFYaLJdc2Gs744C7C3jn/urjVBDG
W1K2oLgrk7S9+UdexEc79YbCdQZltjzTuxsjR5w3aa8YtQqevV/fpGelAKAT
GwG/dKvp8vTi4sfQR55XOzgvYtU5A1qT9f1RZ8vV/0ydZyyPCprbA4llFs0s
wyOyy/oUM6CH8KolavirGXqTQ+BF9RF2w6Q6J1q95EQgMdJwG758zS8BtGdU
oRfY3Gthsh8WaqVWJXR69+MifHRZI5WZoSYq6sv+MZyLX8kzhljXhVKbGKjG
ZhFdN2kzhokNWoIszWu7nur7xw77re1ScX/YVMATuY5KL7BjENztUGIbx6n/
sEycQ4KnSFAAPJqyswTewwIkUpj5tH7PrZHuToNoYEX4FKomh9uqUl28Ts6/
VUF6eHeB6Xj+TkPIps0BA3SyObIY+FIT1bomY7TaW5rCsFJZzL5F33udfqm1
p+6O0+S26Sxwidh19gRW1q3Ob1uW05gVSTVidpqDlaDA2xv0gpsVRmsnrLuE
1rZVQuoEEAr1eeplSw7W3/O32sB8vHBWJtgSF4ZImncxxCPEaiZcdS9bUUss
W8QANZ/AdJ9cMclXmGtET0Rk8biVb5G1yz8t+8Ljqm4YrjHW6N/yA6PGIAfI
e55TuiZ4czEiYaLILDh4puBUONuxVEMu3oq7pfdSemxhd91KkugZ49Ggy/NF
JWY9WJBr5zOISX+eiysBw/MNZxTV/rtMGBN+oHRrIBrj6kXoEcYh4GqgqiuQ
g2m++EB5kdUqnKYEdhi1+BnyxHiE9WZlw0B4IJa/OZTcGixcjmdS3SAtir+a
iQIjOsrzPbW0d+1CYCUHfpSFzpYhJUQOlqZHc08W+iBpTlFgqojJYF+JD8p4
dPIea26VGsJkYsxUTi1xM45fidI98THnjIVWMv2cMwSYl41A1U5imv7fa5KB
+rZZuCotGccHx0Ra8i5T6xQUZbWUNz/rLPi6zAKvmqzme41u9VkRTw/wXtYh
0HDUxphBL9sEHt91xw42fMVGhANUOqneqAvkrpAPfNp/tfeFxyxpouDBofXD
GmYX5VUDGWDprIbDE0UlosAFWw55xFHqE2JCJqFDS5AmiHHTn7d60EB8HXmr
9jJ3G+ypRlAIpmSysFqQwTHP3UOjhWj0hNYFZR15I+CzmaLwVoe4wODrCHQu
QInS93NopR5r7d/WnSdis3LysBiR4nCFynxOE2P5OD+4BQzQIu6as96ToYIp
DzF0rJkZVeTKOIsliqRSNYqAIkwnPI5uxNZLwSvSE0Xo8UYjSsCTWjQ74mGM
Ya4Cjz+YhOv6Emj6ZnHf/fdUBwKf5wHSF2cEc+j6PW2xpm1x7qIE/pfMoCNz
im/MV56i64hqrT/rzwEUz5OkwEGbeeulSZ2rFD9d9n65ZKVMQlJ+wayFeNPw
hM4wrezF3izsp8z7xeBTwvnmyvZ9o0JRrw/IwHbh2IKt2P/ykMSdkXWuqNFZ
RhKVn9mA6SZTbTx4kmHuJOvXIRIPLcDpe7CWyjo2VS780HN6LBvEmND8GXJC
sgbe4uL2w0Afr5bnxiBlOP6tg8027xGi7gN/qmosYyQvIepKakDs+Xp32kSd
eJ9hETsbAwbodRlMQWwkBgidiJpWLQ3jYYtJHF+n5ZZLOVWzs8w8sga/p1vx
fVP/sABPqbK1IEmxSw7ecaE38JPqV+T+Sd+VwOCIgojgkqTzKuR7T6qH1VKR
VvDblnQs5Nm7tm7ntgre+doV4rnR/f9zzA8NJVws2Z/3PbeWBuPTYUArv2Cy
/pvxlPRG9Mvpo/DI98xgPYECNRJulfEgSDlffk5fRsufogA8QRiyPlxIe/H9
LdW/a2mEKXnxflnjlXntb7lrTPPeUUi557UDmH3FkwKQd2p6PagNhSNgbQML
bRSw7zg0emsqVCLQjZKdH9CdQ59wS4im/H8iqKx2BwJaOWmHL9d5HC7r+aRB
HRWOUhL0MCHjeldlIVOY+bn30/E0r7gRP+Z9xLywxNTdsIOX9FuKLrGVNnuz
96E1bz7rkY7ol1OPokRtHyLB4LrymT9EL94jVoIvK0sXkJTNQ7GUDO2gZYAE
3XHZNdYTCj0izchBjEYSbs75utheRqtyQ2Yx4CFqyQPM0f4KiaAes2MVavRd
p3yf3U5SN2pY2O9EXdzg3Le+OgkwVGdQ/j3K67qeMlol4rro2FpXwP3JS8jD
jKFV37prsu36FtP0zEmcyvTsIH3DgrzJum+1NVTad4F0qw1k400IAKaAyAJo
frTT7dpHqYxISAB9mNX2xs4GvcAOyA1qoFjGX6XDI5ydiHUCoFi8TLDTqS1F
Zwytp4jdeR458793ZhYQuDdLe9p286eHnkdDGOEh/Y32yR/YS4eoXZad5blk
V1PHUSy4JkomFZYfb89khzAE0Kt9TanmC+lEKKXXaIgTbbqcqTqCCN6cexDy
Fzf6MqXufyC5F7awPp61Pvq7Izd7CouC7c+7+58mIAfiNdJgfHZ8OEha57jc
Tj5XUWA5yIZF126VSxBITOAcoELzpIoxaHceQUPJAsmvjANXw7gcTsYjPxV1
pTH9gQVizKJSCNdqIlk/de9W7htToXvzwgy5AovOUBrUnY3uV7ebUTXTG6m0
kbjqfIJvC+ufeZ6wQpyqDYPCReMpekYFzik4enjDgFGZJg/gbXnLkrVBZViA
HDNHcLLgcJ5C+dZDXc0ZeWjwwtnpEZLXs7WXJCK05Xm0GFq4PJ1w2SBGyy5M
40HyU8PDOh5AUAh9UhNNQSXDHNUUo3ox0fuKgFyd665L5LXDKBOGKmaKjF3d
eEfmMAmw+q6Use+ACdQDeunS9Sp/seMr2bq3OuScjbK8KSr65n9Yb1LdJy7x
iu3gsTg56R7/jIjFqBTExJX8DmHV6YdQX0SWVgpEYcQJpKwdFl0JZR+HZN1b
WyjNhRjND+jpFt//FopBrM0wKbOYiCbHaN80ke2oqbWATJuzved/1wzBOxG8
8IuONEihYGSSPbxCbr7e/4LpExyFBwekPixJJ73wPOqzFrrwQRCqvYyIM8hx
8ghNPm2R5Hho5/PXNr9CzQGjpd+xbn4Gy2iKVMhScqLBztvkJX6ARwhiaNSB
tXeTFx/OVyRWzM5VKXjcKtFK5/2Pn3XL2EdvSi42dSjZjm2bLpostiSrgzDz
QPjJ96uIbgkbn6wGNQ31X+ZbXdAl67b0ZD3cBYBkraNTMMFTctulEKbPMkJq
4PA28eWCYG/unkFzB/idWqVgody/iiruihRrCNE+DkzbVcesS41h70wNn4K5
Usc0xck1VfaS8eAqtwhdDeXo4BHCL7QkYD9cv11DcG6OxvJqTeeQI8ggxroc
hOeefjO915zDvOmXwrO1Yc1yptlB5TJ1/QmDCAAi84/BLbk6As8LWj+o44Ft
xFzSPDp+dZljKAQ0+om4czdYp3OlRWyHs08M07SavmNwILoEtkIyC2z1byWc
id3ponOv1h9xnkfD5cF2Qv8eeHLf8N7Pq+MIEJYlz1WWmuelRA6KuEalywFX
1AcXM/aXRCrG8fhRvLmJ4QXhiQRxgjlruJ1kus7QpDy8I0dPf+dFOJTKXEv5
KXVbeH/+KebHPpAsl5xUJGVOb8FdPpvkss4aWHzRHATr8JwHseIF5npeKwT+
c3hQ3t715Lf/cnGU0QdAEj7BxRgkEqUuYbCwLhv99Vp0UDXi2jCtYHatImER
xZoCNi6MpTVKit9p2IpE5C+dy7BkDcw8zVhVrmswM3zIo+tH+ynFqDqII113
5p5L+20L2UvClQJBEG5iTekjtedWGf8W5jbuvIfyxu6bq6QZz43bcU8JGJ/S
vFmeTd/d28wVZbujWQRB6uke3cOfk/4APG+cAbkZ6EDz6zI8pHphrIqb0LxM
pahQ5WrNfaMIQIehETEQM+N8hLnVTdLTWcRZl8Nm1T1y1nHpDfN5w/N1sdYP
NqiTe6Ylpd5OwrWo+skwxH1RDnR6VU/lWAMgighfoAYTcd60skn19wNAeagI
qehm6eOM7usYsGbLKtzYMfdwxkNZN4LTg1wKMiADQP+1SG5RkvpE7LfGxknn
lvf6L0iu4vzKbI+Z9z2/i5ukFJ7b/Ofm0G3rFXTYfCh47l01mpAgUwy70V6H
E5a/xeSybDNTzIrboQLOZAqxTofC7WUhV+ljP8jz/ckL5XWj8vb6RYqm89lE
TTBxKePuClyidZf5+XCxMXUXjk/eogBIvxFYSLmNOiy7xVkz6MVsqu+vnCS0
s+KU12yJjJC//A4PPDA/+71OaGW8NuLBTayNisweMhSMcW7ihFAPaPkHRkqJ
GnBUvnYDf3zQylzKcUGUn1ByB+DCX8JfsInZj7ElsWlJun1B5cmI27YZwocU
tqiOqecvWRNyZeA+EuNZ5LsFEKXikgr7i3lOe2mDWNnkSHI05Ta/PJ4wt1ok
7xwDWcvyRLOYW1Vlj76TT+TyMXV4c1iaPh+YJFDV4VXdISAegQxzu4vaauXK
28p1HTdV9krezQLJli6HkBodFfDuch7vbEEzdur+9sGFAtZpdE0MEsVmYTmE
wn79OZbs+c8DB9aNKNWaHhCB+RgSygAbfJVsZiYGd1r8Y/Rw+xdwCiVwRcSA
dy1Y5iIisNA3ihFw7Xip0PXKtxJGPlIb3CXSGxaHmmiPNusRQiLkZAAHqvaZ
nl88DvVDBz6NWld2oyN7Kpv/72BibNvJcdpoAoJB4DZvgE+6anbOq586Ep7E
PGB7xQFzwz3WNxaNfughWrZ8YP5SOa/Uhy5rlmGSaUCaJHCJ6XrfxaVR/GPp
B6MUto8fHJlAAV65nIhes+BYOuk/3/JCowq75cL6z6RYcrkbxlgDJDsaNe4W
D1fKlRmTNJmFUv70rmAUahvJeXIjBQoJo9iDuHg4bp7rs3x5xcMuttMRgc5q
RDRAtkvIULzL2pxQICe5JngluDFbjvXvO4acA1ldIfr6EY87fR8dyN/uoZEc
skst8/Mv8XxM6XVUrJ5kuQCY92f7YNMCIUglOrOZsdRkaYn/o+gf36myse0Y
Sjd6dQptops8cGJnqFwO0oZ2fIToBI/rj5hulo9AaFQRhMaXUcmtGt79Jokd
Ph9OfYcoR/VtEaTqxH572THT07Jgw5oqKviVKSTMjvReirvOGtmx3gBzodvj
517D6rWUs3cAlXBvXmtcGkM8UTZTgqKPdR1n+1e3S4rGIfvF2ABM/BZSYHrW
dut9FOh2NlF/rhgphnSkDSQWwEvT7vmRQhUdegZynenBW/wtU+cJ/XIQHyDL
t2aOidtOQRTuPscawVyvyUl1E/EA/J9ozQqnJWyiXLp3ftV3l/A7MI1HH16A
My5ImBjHoikTXGlQnXvhrKRXyqzZ3gRsh1n3+WDr3md3lQj35VndyyhQbbdQ
ehc/Hn658HNl+ulM6MWDxiwWJnuFr9pckBpjfp3Qq0THZVIGS4B7ZsEkOEPG
CqfJgrQZr38WrTjKsQkSzHxzZM1FnGwxgcACPXw8+8WvRD8Ec3q4ktCVzOKw
RSTonlH3ha/gtZD7JZ3BDMQFC6/nY2kKx2wH1mV/PeAMbBTi9NsZ6dTLAZrJ
UDNWpbRBY+N3xgtZ1m5dencemvyXa3PdB9SiJVigjUzsFLiN9+AfSjUb8UAc
P40FWb3KjtqM99XlDqpoaRSNmqroI5eZTnScMxhcWvv6xQvK9QaQBB+tFFZL
1mYDGn3nDydUoxMus76tzmPX92sZf3eWhXvtVnYnOD/RlQ9tydRWZ0Tvvcdu
AlO8uMZdiLq7xAj5bx++CrvH0gUGqbIcr7Z/2oVHztbm/MJy9z9YjB1HXoex
y0Kn6XIHh/VaiFo1Z9D/r0oL2ydzyD/nZgUAlSnlB79C5g6fK1r4wlKp07DP
rKCny/FbPDkFKPDkDluJrb3Jg1x+v2/6MVtPMeuCYdvs1Wi9eiTU33VL9SUN
4rztOBjm38NJnZqFn+Jr0OLCSOwoA8MpF5XxEyfOYNyk1b+vbRhhRI1nwyaD
k+Pa62IB69obCz/6Wu6hlbsMCNC6L+ZjOoTGj1Rju3ljpgb4NEl/rJ+eHnwa
PIijC+yuyx2pwwHqvt+be26WQNGcodggBH9l0j6eHfUph3ivVb+095zK9od/
BTTNHpgz7xRjDa63p+Jx1kY9ndiobHBuEHFO4Qnotezo21Y2JbTBtDhn4JGI
s2CHLNeccxCrE9DG/UG88PwysP7nk52HY52kr4j+t9xF52zQlwGlKuUtr5bs
BfwKPtqt0zXNP18jHlHycm5qb4HnW4UnVcigBY2nJejGsacmrikwIEiTw7Oo
Unm4IYRH3lN1xceBZM3Zc55CL5qBrqqDmEqbWSciDsV4WrFVrbKgxgFFbAkp
n0LW48WmXvci7aksKoJwPnqhJyiAS6W6J84fOvmP/Nwz052dOhEOEC5w37Fk
HCTzzhC2JNv+y33FlX9YttHuIWD8KRgbpqkFKl64dWMK8qJITB6QvtSU/Txp
jbq99yjJn9RWmnfjWZs7qeYdTT3XPicooz6Fy7HjTMS1k7ntkHp9m6eDWqQd
XBeD6quRMKFTIIm9Nk3gIJRmxUjvtQ8xxreLnfZlzUwyPNOjkp0j4cfEqqN8
dZ/TMkTXgwQ1xL07mZ98C2H6SqNEM8E/c2v75u+/h0iCrFCQjj4nyJdzIheY
BKqdkc9seEeIcu3woFCLadtQdeHFLgIFvemv3RqSaYt40aDesPwDc8YsWtg5
cSkWuKEmz76vGE0ZgZzkoD4QutgJetgXnSPLPZ7qAd8fVQbxLkrZIh2pZP2i
9OW4MckXoj03tOr28bleMfKyS2jdLawz+eRFuXCIuXnN9zLp1I8uab5r2oXb
SNSYKgaKVU1ISi/qNIAq0CYlg1q1qHOr12r8BcFrg337o+nJeldqvzlgv8qT
6bhSYp4gOC+xXABrm6AwvI5HRYa2IdCKKnlnFBqPljYLmT2zQSwsLiZlg91D
iiKHWT/54fXheip2shqbQDMxdgTh/trIVLa1FVfc6m4hQ+XKEm3TBOCr8suk
XuQVNq0PhWCum5x7NPyDEs8FTJjtaH5Yxnvj3FBc8WqyZxNN9VBUpQvEqySL
5fYzUJ4WaF8VDePfxjcUttmKZb2hcIEoMnxgFiWPKPn+2oUvbAX1jiCk94JJ
jYYt4YKJ5XWHbRv95w6f1GdJqSLjdcctU4lX9M8Yri1qmB13vW4t3SQmHdX7
WglPRSuWJeYIS6/NnpX/FeRaAzlCXyF9W6l/Bns7geI4+uoZXFuwW9zHfm5O
M6x0pfaUIl+5mBUY6LU6gYd80FLvrz6e9tgMtjXzQhaxCjFLBAk5/3gFg4sk
ijRY5XLHpcBtY+rYglmKeN9y+W8QgqsIqZa+cLu1ndtUfXBTkAV6ZH9aMM9L
ek/vPvqDOIJxP8z+csSFbLYh1qp+h5BAHpK/9s6GLJ7pSd1rao1sSCAxz1CD
wIyowJqyaOEoBa+An4h4hjnyok93jEGs9JFOxjAdHMK/QG8WkrMc0FA94Drt
5LWSuSUncOqfwKCWX5GYukmmDQPLCAG0RGQgHjBfFMgmHDidVhmyCcmg19ei
WV5d0pOG4Y+NfMUJlz6G20yTRUtcA2tDOOtB9dAc4dYm+Jp/Yw6HhsrVCfG3
WgbzjSWwu7XYLP9skDa/LAKmg+yhxqObE9mZFCqO/zDTY4iLqGiYQmIKPBZj
pmdDb+ReugVnoBiWanfTEZ0hu/DcXz5r36d+yPIYwvv0POWmgCCmDNED9zoS
+hzlxZOVFHr2FwKDP/4XS9eUVkAqOcResxCk6dnsWsyVVcB64lJSvD6dj8+m
nTdMvd4+25WNpO+fEFV1IE/FjV5VGZKds74jXB7qwS4BPncQZvtntWn7TgsK
xvpJtNs3qrn3khdNg6/lBtFnvoj4/24Hjt5mYaTsK90ncvOUlz1glxABQ2gT
xq6MBbu16kZYPHZ3CDZ46py3CqsogRvhr8D17pu0lV7WAd3gCQJ2XW+24ojD
VDVs0qlE/3WA9CfXKWYe1baRgecd8UeBVfGaOaNHi+uw0UUdhZd/mvmCR43D
kKlFfBWhXev3igxZbwyAY6U2aEUQcJg2ppYAndtj6kDr0mgwWbkdIimGNue6
U/Dj0avyWRxXbkXdAZkCkQWJr9oJSA7VRs3bts96hva8/PxSi3iwm5uDKAm0
rr3vn6PDL6Yg6u7W+OQisSNtV031NLvYcjoJD5gbw53U/non9eTU+bZIxLgq
+oRgA682yOfk+A0WFrXYVNx9224mmPC2YkyZRHteKcpJwwWAN4KacDNyN2QK
8x311p1maWGOqhF8oInxlBkMEuBbn3rJKIOZjtr8YJr/bK2xjwKom5IJr74Y
8lZZPohdqc3zB5IzVGad8h9Y9mPmkgJhANJxlMuI9aR0RqKbgp0kQD5+El2+
XKBznXsxJ3XVKB37ImuFmPh9fTSHmCUen5Fyyz5MEmRXTjR4rqzqBQuI0lx6
m8v1QveHNNZb+8bml6rYd7IQiab9w0KJnMD9a9ryXWUkYS85664FZFnz0PiI
OXi42VqH14IQuPlv5kBG2ojYfABnptpSvNPoobb2Tn0iERgfeTicvycvIFh1
Ml8YAjFzKSadwhEEnwOOV3r94BKZj/AcZTgHsvzUmNRZulPo2AxtiP9ozIfX
5+LspDo4gapUxTGsIuD1en50ntqC4wJCCKtxOJ7wy3BWRPxfAHkuN8HwUMlF
C2T5wdMCYpXZaP20cGt4rv9g4NaZDydfUEhHNuH9UtIfzTrhvqFtwqh2Gdm3
o7qGJJIc5pWy8AlKQcUY8gZX9Q7q2hww0fI1nXNpLk0oKz3soqH4MmLn6MFL
0Y28PADiDXFeSUPPlSh4RuP0jcBeZKdy4Tn5FeCkZdmk1awltP/DlgwUW3kD
+qUmUlGOQoBznQMylh25r1RQx3VWO57o8syQ3rYPu9O36v5dwU0BFNk1OKG+
APrZb6HH7ePY9h+O3XqzULHFvOEyGdUf7O9PrSKW+OtpCMahijOsLP8+3KGI
kzarbNCG3AL0/qM2Z/CMdKGZane2T3onS5Oau5hHVx/mP9Bm2gEl+HBF5+UV
r+j7VQyCTMaSpGix5wTOvQ60MwVLhCyRpE05WmM72e6A/12e4GHG6Ke4OiGd
KeVjWht8eluk7umTY9sND+Bgt+xE77TixpPM/ExzxVadBWSQmue7TSXpJJ1E
Ovd6Z8bmhsn1wpdNV/GvT7Hq4JAA0n82ZR7ceehbheiKPgoxoYE0GeFp+Z13
cs8CzX43FnLLGk4N+5aJpRkxbwADH/LuNCQmANu9+g9mSH7QzCCOJntPFlNp
k338gT8dcdYuM6gpaGzF85ejZ9gHv949GAhjJRaD5Ltd7ZtjzIBnrzu+IQfs
5Zc30p+istGZx4RvpvKHLefOgAuPFL3gkBiaubhlCle+oXmwG/hztfGxXpKn
kyjcw+SQjtNu+Kwu//XctfPXkZ6iO6GADVLEsfzmEZAG+YoBRUsQJdPs8/SX
jsp1oGU8yZ4FMcWrA45ycR3RJE1v7xUrQb2Uzd0B7G2jyAIWSZNXy/QGrWPF
rj5eNHJoLW6rb0QSVeZtEqXzMtAb3Esr/0izMYpwE1ex+QLifO28f9Vyt1Q7
HYUtX3AdXF1XzgzS/lRzg3tAlTp/H7Eo7SZa4R+Q18aFaYrFSB0Ww/ZjEOYq
/txlngZTUoGCtcJudlKIPLhC/zDbkfYE3M1QAxRkPsTRjH8Y0bibF3HkRJi0
EzVmz5J1ZmXwZNTZGErvJSgEU7vNO7Oid+MiGOrWrcJwXD1hvqt8X7k+e1wW
TlWx1L/Ql6N6z0DlB9VhH/9u6fyWuqmQUinB1rbVGfP5ymv7dSN1EQKDLpMJ
h5tPqQmT60rvh6Y439YeTi9dn/bhCsk73ye4YR2QanN7M/0VMVOWhuQqj+iU
G5D39CY4wdYabPnIMhjsJTcbBxFaa0DQq0rvTnFXZIDmlAO5y386IzAEK8ie
+kW24SMcwvVPN3LV5+kkuyIImM3omNsVtYJe3WaH4NErRUNUESGIWcihA2Sm
dla/BVLtKff9urE9IisyQxFg1K6u80XXEOTFGqCvZbTkCyw/Cw4W1R8HaqkW
cgzf7py0hIzF6n0s/LSRvgN1ECBLxVkFxuYs7sb9S0rLNSZmFJG3xFc3A23+
wCnZxoTT6I9wA/0vA1jnmECCZwkppsqJIU6APGvIWHWD9tU7vCEmqc//VOwm
d6YENbL/JBF1wq9lx8UXffAXUx+IPeJr/VpuhWRLAmL1f4V/z/mU5Io0NTLv
cmn02IOHDY9eMt/otjGA887D325vuHmH0uQicCP79oUihJ8xSys9iiY1xhW4
lZG/Wp20WI/ku9XjtyuAzkPOdkaOHAqWyiJ4obuVnP+jzkIyqJUDq0Is8yRs
KIa8pgRLxq+/P4Ot93lfTbY9ItnE9ygmgp6hr7QyAiFjyE2UQAQjadmnlSom
ntLmuXD/vlpD5SBncclBgGYOTR3HN9SetN22vz0flfhL4NPtS5nr+B0Vc9jB
+i8itV+au9leeuB+2PXjq/ZgyJ/wBuazcAz2zwir1ayNHy9qMQtYdTC5xnoh
18Vw7y0ojXt3lZbpnaYjXTTcZezLgoMmfgvqrl0FmJrCjitiNDMppq+5WIhl
HoVhe6YEIu/cYyyQeMTEk6qwLu0mS2yUF7yvV30G9w1e/rrGFt3IgTknZHA3
VnDMj40v2Q/ZnX3p+vCW1NBE5mn1S4rxFMg/3Iybq6H2R4MLz/wbAmzmN3ZC
7D00eM9qJGt74BBnyNwcpyusEgm4CJ8RD0nFKmGIA+TbsDWu65tyt3G7df5S
vsdI0H+2iMNSH0/Ou0KiPnSbCMYYwctLO5YTmj5vfc85w7WfKtJyt6yZdk8Z
FTonhAbEjIFc/isi30Uuro/Z31A70xhD9nFuB2fIVjVvH53YjUoAXL6lhDji
vMotx3Hw/LKnY3rOKQ1DGmmkQI45CiH/YHQ2xBkvJsepMUQxTw7TQkGSA5rM
occoBCVEvhtRgvXG9HNlfQ/Fn+qmZ2pI76zBSobd3TNuVJXQ1GSxRSsjp9N+
kCa0SHaT77u+Fiaa0zF0b53nDekJd1ZcpmhazbnZa1i1t4lTatkUDHrKPjfT
MFeqQf8unWKAoW6puvuOaItjkpSgsnIMC5pvSyR7tYHMMKHjWYEpH8bLFdSQ
IhU9xdMs+7F96LiSwsNBtMHVW8a2HJzt45xEF/6J2VcN0/vfnREnDwiJvBxf
d6lhNTheR8m/wzPNIUAB/xHLIhiowGIaMZr3iBlUZY88EheMGzQ4L0qy0Qro
hTLgiTnI9ecx9gQASCYUiem0foa31N+AFW/5xtNX6NrIojRUxIPvwWwvHLOU
96H21/tc9JSqHbjfLHNUJQc/e8N+7whKLN7zccx+H8bRoG79MI75L9nl8GGt
H0rMtQBMVVcXlFhsYWiuBZV6Scj19cpfvOhR/eMyyhO2xS523TR8TmJmrIEl
T0umFOOyVloS2sfRUJHApXJ1YvHQpvAv20fwBqL0mV3Y73F+QtkEcKDfeJ4W
vU2yFkNemiX0ZjitspT/2oh/Z5IgVvNzdncTO0ywkpJQAfhko1/f/v09auDg
g6zvhVrPwZVOF42lFvQ3kvHuK1CBhGoI5t3j5lD3qcclXIINtdhSxQNe5QvB
fkPNmnc737Tx4stS527E9EpO5BKVSrLBqXbamUCEE0hIMHcpxlSHSB+kGQRE
9l0Zld5yxYvnpi6WsRaDF7oU5erDaV6DcVUOKkIHaRGtpTI64OxxVcpn9jJH
cmB0smbMiEZDFp7FIZ8Y8mcId7gAUTOE+azf0Hx+ty8kFjudKckFxs/hH6n0
tKyyy7klDdNdJX23LXewLtTrgJ8RN6JnMxSlNUd9LirRjnveMMExXDm3cuZC
f6Fj3G/+QoSbRFZd34SU4DUz6lE5Wunou66v2+fzgktaWsMmdtmxyt8mMDoT
gy6gLi2oCEdbm/ZRmWQ6wvjx5pwGc+My3r+fdPYFqEY+CNx+2WohvA1iplOL
t8e96VWmdPRMJIl71mRviPlR3A/wn1qAtacr1xvh1npzcbVl1TT8FTsgDktK
cAEYOoaF+pjbodxbqr4PeR02Y2Httz5v9nz4Y3LsPC/FINiCUWKiMaHvN6zu
zGkz2Z9p8FA25HVUulbwRH2cYVu/mTyoFkJcTT3Zfnb76MpoxyD/ctSh2I8p
Si16gINvwqdAnqoRj6mGj6IfJJFsxsb5vo41h08UO5eXxvHfvl+BocizLIEX
3OwpWAOwxJHk8fRaFj1VzbtR+5CUQ4uRi9Mlv0be9UT6u8fSlHT01j2iHGhH
runSyjJ2Lmez5VMHq0QeZGMP5hLwgMm01V7WNv8YbxnZGRgyDdYs0NZ/En5L
CqWRSqe6HFBHtlRm1Oz+yoe1TWJKg2dWMY6pMyjQHwqkGS/cOvMmgoJogSHK
kClZYMql4Yqc3hZA9asy4OuP4/cPMdOTk23p8SeE75vIJCH1L8GU8o3JvVE/
3Yl/llC+aOWxmBmlh+ZbSKKKWNniOjirn3LS+jm2OFjzV27BtgHiCq3YfKdO
l6VoPGT1j1SHD1UIrfMLBeQdD1DnQGuNg8n7UffBA6zunmqQkI0cLFtxm/JJ
7jV/ikuhy2BWxzgDHDK3JIqu5mZFLe3qxUAzTE8F7f37jCw41/CkqR32JB+Y
kSuObj4kumXbCvFyccv6HPbVJx5w704DvmZV6Cn2pcqKMXB42WVc2diVhZNi
XHBOtj5GGH3TRSZ8Hk3Bk8Jfh40/FI/lnmcngQlVU0QRIkZ4+q+nzIN7Z60B
ESM1ohxelu2YWDZ1+CtMZF3clEXrjnbD0PUQfUn1/gX4VsY1mv4njstIejdM
wUjxxA2Fg1+ihbsY//prHlUx5ULqzRVZ1CR5W8ToLCvmrtOP/73TTVLuholE
nVwxLxyYktoqrzZpEEHXdvMBOEfvMEm6R158ZAwUcwbuHaVgZ0o7NarJrfra
MQbNHR8iUGHtoPUA+t/oLWdzNAQFyvLBH6EGQl+JCMJTkXZ95usX1zYdV1Q2
vliGwXZGZJfDeRqYFZXFjRDyh6aUrQXwKcoJydiAkPZyBSbMj+TL6FrxP+w1
52CEwd1GnBZWGAZIpCZnYC7Lo0fivDYQuDzZHvUKBZvMzRj2fKI0eLZ3deAR
1zR5YSWGFUyhQH2ino8l8O04py/Ab+fhXlp8HifOTDq3BctoBMzIuZvYIROu
duQngaKE71VIZKZEnJ1ZaGV2P55JDnRdW5OJ1+OaMBRiHFKF2YLKHALF7cpH
OJz4EhLXaYylbNhn7pJSF1nQC2PzOUgOx/s5HHYUVQ+witMYSiNpwtrE1Acy
xSX/YFtwWww3mrhRZPwq7oBpkUgomT533Oqfz25KY6WohcrJ597FQuLdJo38
nc0plaL75eQwaDsgr7eI+wK68xYMoL+StiMKirkgg2Wf55gI16qmHcjYu7cT
Zq3ALf5P2MM5rNcbhShOHrT8DWd4HQOoYeS5f2ZZNUltiATxeVT2dmJ5apEm
wYC77rfNEgkaWPdycBohxpUY8LiJ1xdh64S1DTJuYFAoAeTNW7giN4gZyxzE
L1mn1EOqivdFV7Uk0PIUkRtQkKIcJZBdRBZZUi52JeiSfVaeqz+tlXJbnMAs
2sDHK9danaHnt1Gg5NxCvDaPWE6ZQkd6veNhK7t9KfbBAew3HRVtoqVcwtdx
mPBjENcryPxlgTSyYPlOkcMJKhiXgGzC3i+m/FPt+LOL51i6hy+fchABD4ui
2CSCYGpFXOAYZhT7QKp8qim1kmKL1mUkLMkr99RIG33rMxAemBcvjPcsBg/N
V7uTFjSE3ckUTQ3oKI/gStOomMKtVUo0fJiueDAqJdvs5PaEKiNoTugwSpyb
TsAb0oDi8mhBn3N3yePQFDy7vm+wPvUd9Xooz6jonJXauS5V9HMc3lW0R0SY
Vqq+kBP+jpeRfWzpNY4IPZ5GpXJ/4mrOQc7cV75ix+/V6uCM0MZ+43nrzRha
Dce9rpyvmOElQonJ+uKcFJPVe5C24b4MVLHs8tQzTnmFGFB/2+sYj0eh9pfU
X0y1NFi5McK+Mdc4cIcr6iTt2VHy18vENqfBJWwBqoIpHufvuf6W4ogvkog1
2eJWovnsslvTwwlbcZJ3Fmx5BTTCLi+ZuYlDBVXaVvEJtCNLSjcoC1ZXZcRi
rsFeqGKx7VxI5641izZR5iQUP0Lx0TnbAVbX3yMAnaySBlau7kfn6HJZHNh7
sO0x/JfdKRjU0gbTA1MyGM2tEhOfLcS2FuAc/HWWsgTV8ogfqHWMSvnNsJjy
1slhZpRKPFZIn2cXV77irUNN5MNr356XervSzy6385aFKOihdEQX8iAogQYG
Nc9Z/67VseVkwQYL/6EeEi8errTsmwdLTLiREysMfcDJRE94yEfPq/u0yaF7
LrYzoTaWxvO8hW+oJwuqcBujLWTE/bOrJ18ROREmmHorUYNSsUnTkM0gMBoa
9ae8RDNlkVj8OuMdWjAxctB3GECSOVnuCiTYMF8nx5Nij2n8p18PCl/K8g6B
EgWCTq8AMb9VnkaPdxweo+niQN1F15c4fDZvjRu2+bIUiA6AkjTtXp8EWSlK
dwdJmS3ab95PSh/Hw9/CWj/ksMkxIMoBZPLIQKEJrJbAn1orOkwFbAGDkxMs
MKLWn/VJ4gn87z8ym4tWb2xDZ1e/J4aHccC4PZLiZpzAAaIYDmwxMD+QFyCE
VgrpijbNBEGEAmLrBSFODoWpoRtCUJlXKKcUgqF5ObEL5gJaoDkjz3CcyoIs
vG3Jl1tWyserHy03XlFoSVryysYpdXJJUzPxMuzjtAw/Myliu77QjvTi2BoY
9V0jJHQowY9cUzSScl3WszNKjGu4kgEg07MAy4wAZZRMFE5vwV8nbQXAkoBy
VvqdchxVVL0Qwx7q568juIlcDvOHmgTBVNFuSI+A8nH0i/mJxLfs97xR1m/y
Lie+U2lVp+MC4fePAStD19tNAV8qKTCn/5O+aX5aUjIZBFhwYWi5AipXLRwO
vaRzETIvpgCufo5uId4zxRxXn3T4FrW11D/2vg22aIG4US4xFxKhNpPvgnaX
0gOu+cxPReQG///1uvXtk2sZub+pgLub7dB02nSSXcZnDc1S6lYkCG6hgKmK
Ori+LNNbBSybsKFFqUuLQHvs3a+8Q+x9wl8iwhe7Mji276BsHewrfEGHW8L8
kugPyK1wLd7Q/9OfSNpBsKffB5WVQwneTeQdg2OuITD0Z84c94BSwR6eXmna
j8ktqQkPPOnNG9KdMsWoZnWAnbsFxC2XlNa7lD+uQwmR6d8wtH56EecmbRw4
hgWl4sRFpUt8y34YWWrC1vCuTSfbrgOv1mvRX5dn/r+Wx0j2XGMoyYPos51e
LCN6bxDwcmS+W9IIaOJjcM0UT7MtudYRmoLZwYWCd0MVkX6D6SRD/dbf56Dc
q7jaYB8o0EkJawBmmSwPf060DsW+VnpwWmS7X0/RvveYuSvbAnQePx7yd5i+
TwcsNl5+iWwx3zshM2xZqB1tAJjdM50eefgakmtEoVr0HlIJniO9S5raSZkJ
CT9tNxOHF/AcEtbqPFdasaJWdgpxJwpz9y7SpsqKVPfeJqO7lOP3ndy34Nzw
ON4HQ+xJ4OPEVqlCP826ED2T+qMO6bbw46frFRMQ59nrsoCjEAbVTkMsZtbX
5kFM2dDD7eSmZUOyz0toZpNwAGt3SDMleDyG+pHkvAsVVhLAO7aDNL3XyjaY
RhKQa7fbJ7s2D/HKicozKLnT9cUpvI4iwzMJUOwxFCZRZFKvvhs2Gi3sSoh5
1WVOSXHgl3CJkJExuenwyiv0HizYE/6KsrVRaXdInlGLCn+oxhq9hxehAboJ
EMzn2MSqAth11LdFd+yzXCHW6dmq4td0c81ajEsQof+6jgvntCGMss27moS5
EhQzsh1huKWH3SMY76sfASl9L8Tzz0et4/yg8L8V2MQGU/eHNggFlahzwkw/
ASFFLbZuN1/FTxBQmjT8f9Y5ziNG4i0m7HHPC2MxctYCSzF0oYBwUvfmAKcF
xgyH7tHK1nKjCcrvqFxh0d0fJ4UF49FmuXHSOoqfIpwAOwfke4ZZswkCi4u5
l3avcdLCC6Zw7zxzDMzSB6aGx6t6YGV8PH7YhJ2SQss+t0fOaTAWAEHM8U3p
GtV6/Bjjm3HdQFp7u18CiHfQHBtaN3hCgu2UaVgbhBJdRCV9LSjFJod2y8ym
dam0ciqEJYZlORs+jve4rMP8u2ZRmXIHUZ3a5K0vEWq/O2wCMf/Y73patjqX
XuRgKG4hlAXm7BuMAWYIOYTyqHhTJdzO8p7JwdIpqwj1DaCCqKiwdUDYEJm2
V2iR609xt+hpKGKVp6wssDBtDBA4BoJFengeYya2+aGOhqo6yJFKvXUnin76
q1waWrqdVNrgWpgf2tbyobkur4sosJeG9GcUJAjgHa0/PCPN1Dfq9lV9ZPdb
ss8VvVoCRIyRIGeTbe2MTf6N9P2AOfrmgmJMHP5nyd9ljEvlRKvSL5oICPCG
SDpu4Gm3RHr+lc48AkEApepO2/78cjOpQqN0KtUtTDghiKDMvbnKAseN09XF
Calx8jg234XeoeZe12sd625jRDvFDd9VRDKa6myvOCLDYlzLYF9TCRTpncWQ
05myZIZeQTTdwN1UsVrrxzlCwtBZl/bN3cU6o2rmYqNPE2oKLh5x6Ztdeeek
DUixKRUjQ2h+3XpdADn7vVoxUuiObMYLYMlOJHaZl+8mxyq1jUSWfrBfOpuW
BTNn+fnuEzI8GZEWprmPERipMlms1OuYVS1J7HafdS3rq07kQIIKRW65omeB
EIK3Q/IFtFzJ0n0vLnvstpHDDU16ClKiBU49mj1ar28Z9qy78Rpkt9dA49qt
2MF8CTYJq0p8R9BvON3hBTypejOtGOVzTDRezlu4gv9e2/eVw8ObA4xcOgVD
xEv0jV83ZqlVrulKUsMI6bswz5wTRr6ZVTE50YlNhaf1Hv9dDkDNZaSD5tnj
QqWOm2l8d5dhVo1AodvHADrF/EeLCYYR8aMWqFGOLJONO7tZMmBR5i7IokPv
lyRcwFZ9QsGBU41KMqrJ1GWp1C5LeYuD5U7JM/ZlF+MR4K1Ajp8S+bM+v7Ek
PR0GkB86cy6w+R9Sv5VoFjs60yh67ytxzdmUsjjp2ElX/E8vCEAQlpil+Ex/
DvU7OVkRcaG2azJaIPM417W0toAZn3A592iH8D0NM2Jl26yMYNEsaD4/jJRy
ciaBZX1f4Y6rKEjef0T6RY5k2HokZyaGSdoKufGqltaFgcFbRF97KvK6MNRy
qKE6PtRUhmn2AQ5YXwnRG/A5FdQag03shCXTnM8YGZu8ERFbxx6OCL8lX3UV
XzLhUvQgg5vHIKf19o+z9nfW4wrZLy661EzTlSSa7S99O/FI7UfP1MhOg/jo
EkvoXktz5XQYDdk/rRO5i2DiGCyBWl1Pgi20650F85GZIGD/Ykynn9OEV9Ef
03pImjKUHLjSp5o/V9cBouryUJidh2XatWbTpiLWCE44duKt2jCfcgfSJbox
KdvDHXcg81qz3Ijw5UXLVxGCAc1Ts5YmcxVPvhap77vohPR726njEacDRwOW
6F6OeApTtOEnRv7e0XYfa/hwTQ65/KWi2m0xUtonq1wm+25/5M3jYPSjcriV
CdHyb9S29isA0pbrm4VLhSNTxuro0OPtcUaSCor+cpRgbax9K4ykrkWdPQNp
bF5hm9MymfMSOxvmzimItY9v+NmZgRO6p9JDQaxQ4FgYIsQWN8Rvj8J31ZHi
n5v1y+TEnQpYciBvp/6RS2WUjUgCAdkszBw6lStyITGJns1AEGvhoYFd3GcX
bL/i1eKZVGMNnt9vQNYwjfhs+ZNmAIUcoK+enJpvssyYtYxyuJ2Et7Qr820R
xRg+AA8y99iLbwgMV/JAS+9lmacQtdZEcnOKbPbWQAZI9JHIsqGq9U/kvJ5T
xKmKq7KtkKJsaJRGON5UcPTsZ3XfQo+6BtEYOebWdYkzu18kbe1g92WiSCc4
q/qkouJCvate+6QsxAMG2o1qol1RgSlb23Dz0fdC1jtzjw0DGOrByGHhNmgN
wWyxFyUqclRFyIAOu/yNabQQOOj7yrIz7xRQVV2/CpGFkpAw8hMbp3FjIr/j
M3r7le3Kk169WzkAIkMJAHe3G1s422KnqbphS2wUn3iNIo5PSfZ88S/iCEpC
+BHc0cr04iqJtumVFM4lUbT1C54wImzTMUrhrie+O6ArACpbJtvBWptSprVL
GOKZIoOHO6WaOPYGAMX3eegPII2vmAXBWPpnt1OJSRnFKcroaazoNltoNlbw
3Njrhb/t7iBNhPKLYXRVwe8/ojGlOYjbzus0ajAzYWknzfGfNAWb7401RtWK
aMfUo/HQs72v/hTkKk+vGq31IE9Tj7KHgh2DVCMixJKTRdnPRD1RcddL4oMP
en6Ire9ONGic6wmY1UuKfp4aaT6HpClcivbkTsADTP8yRItZTrVO19JMxvEy
eZamzZgJfbCbVo6fWAD92S2UMx+9ASQ7xOlFkVaYwDrQkUuqWnTA2Ehuke3t
JvmZSrgqYCg1mhdTlajxobwViTUD2ibEVc0mO2Az+LXDVIWH12MV6RHSNdnQ
jikgTrVjkmW9QTETZk8CExAUIXQGPcanL8bbPiDBcMOA4xsce63+4YT2avDe
YhIMl/9D5FAyQ36REkruL1mCXnf3zBqrhU4sZWGKabqZJEQJ8i+Uz4jImkfO
MJkqL1UEwW3iVWXRaxI8ph1oKY3X1V35yEjMwLWTzv9rsmbeez1gv/rX7N1b
fXyO1r4TkdrJgqcqrXHJpwtl64OZQj2iVgda/Yer86Gnbi8pWjBz6a5IhMaU
O0mJ6pYvRsfhFsYBav/lHa3iHH0yIwjWhzZ8tsRa9eJZFwLElhHBQmTQK59e
Jb5I+e6FMoNAYxU7rXBjQBYNKD1TcS8q16pzE+lAjT1jWxvnY2zazRtMeAI3
dNmlrCWpzdyoPjGqc4M08S5o+mYOVOfbu4Ie7Z0uPo5bEV8zsTM4wPQolQHz
pch9T5WRc3tZ4AO946jALiv4r3rFIIhk7l1emPxSdR5UcmAeflb8qjg9kMLA
VMODraD5+dncua4q8NSK8dvyW5gkkHQVdxwWU72T//wWwDaf4JZgC7ukmwTF
3T9tC5oScwCATnHCx4nLNyXmtBDXF7X0HIQEO8PuM4GcO39GvQpUP/kwfxjm
2fNdZequVriDFV91+IOEYu0rVWEPRM3sEr9bG3bNc7vkpMYstajbrx4DGMbd
CBIIPG/XcI/3TPeYrmOsgZDQR+3pueRF2jLUYhheMLpwq4P345D8egu2SBdV
Wx1mW5KJUDDgK+78RjVdMoSrQKqTw2ob30uBdyoq3KgszzlcCgyJ8Z6Tqus5
IvWkUmYSrUeAOjbhWlROyQs4K3iF1xqF9BKdGf9fnS/KdRCNho0lk2pMw4j4
AY7V76h1ULoESpGSY7UC8YtUyX011ehcoh6NDSB1/h31f79h9qKhWRpE6tDa
+afrOWrpUeqFZM4MypKQlugKkkpSjE9YPXw9iJuapjAYwV84hOMBk/vvwlGU
WIl9Mw/FAnMCWPcOUL0j5GE20BaLkz+UWeIa2ZYdVAktv7YcchI2pIDL1skL
W9PLDSsbn9Z9TrRmU1BQBLuDY60JD4uAb8ld5z3dqYo/YhBEc+BW9CXyVRZQ
E9vN5S6tdiWYsFDKS2jTETt9zXf/LLCqM4UyTKtlKuP/Rjdn4wdywGn9rWo2
1hpknZJyVYdvfjmr2TYK/JUi/rReyMElR73yuCGqwhlgeMAw05pjIcG2CgZ7
j5BAcHPHj4pIWgOsH1xBVfdaxB/Z7zwf2xNATk8SGQqaznTh9HCI3nwnBMma
Few/L8CoH8Qp1gLNDxzlBnLqnWqfehmlDBz7n4mUTQYXh4wi3GNijwSI7cgA
V8whKxwKMTQK03FD2J0wZG2FLZjv5Dkn81arUX2/a+Qb/nHpQCrnqct9Xb7o
JY95j25VURXFlFBLSvR+UGT/hZ6Ot8K8zvKDSA1Zp6HRRhtr08BQ9GXGtWzI
48MkkI3UJ7yNtl+cG9pc870oabKaAEroDp+XXvTblX48fUVl/pKoDXszCQyW
Gj1eu2X4/aIeP8J6QJIk+ELJ1jJ56XPF0iJvTPs6bej42/d6obVY5aozD7zy
Ima1JnPBgTNwx1nJ0jB6feIPeXdp+V4STt40SOktBEerwxlgqVCWCZXXaAr0
QFsY8H4O0VUUGO49JgKzNd6ds1UZruiOES+42SgqqIMFLvDWXv4p95RD7nZw
QQBixAzQZPG3mSDN/bSrXxA02Or2SMv+9Uasfe4691H11SZ2oO6OmKfzAyJg
FlnO4H57sMHTP5q4u+4QhpMbSKsnEwkThT0fvV0togGEhKCiYF4dtOYYx7Jb
257lFw4UeEWFDCO9J5+sCL6CwT/4H8iYaVcyfHCcuLiK19DIipEsRW8wEBbP
5Kx4d5+RGxJa2u4Hmr6KbvjcLufwWfCwHQEwboPGz5ByorrOAWmjDWsSoNVZ
FGDAQgw93CAX1OaKHaod+5Ld2wEZJNuCw8jdEP5IYUnjyyrYC5qFjbM0N6Bw
xmJsIj6TcWP5S8iPPSwXryZ1fS07zd3RZGzlVWobP1havsAyqY/TSC6cs0HG
dV12NyvBxg54pk5VoJSSdjv8G9VQqRtM7lvbft1XS5KOHzs6LrmY/QheH/rd
DtlSWPa8Ac+JIJgYrmFf7dKDStXUQI6GXUUjohjiuKBCSIS0qeSTggiLclbc
4QcYzc1RapwKbUXIR+7j1Ba2ZekQSMPlnqQ7kkSHAKq/jpmXFuqVQjSlY/hl
DuVNYJXvBTrXG9mhQH2TM7kYF+ghF0EYbuBYvkNEfTYI4PZzTFmFvYw0bYKn
EG7wmg8rEJ4SlRZLJaBeyk3+5mNjmI7vcJ2urjnLn/rbP8Wi+LiEXYvZ2jDs
U38q4TPYcnjnLRXZNOzM9i5W2eKfUecXeUZQn1zpE32fYC93/fDdVrprdOwd
zq+yxdS34AdKRWzuULQlbmDUMLNql46riz+XRyz5Auguo1ZszwpUub4mGIg3
kb8YAB9Z/1xGhe6ZfRlIKtDd13oyBBmDey4jhkXjcNn3CuBGm9JAjWvAE5cA
e95CdIWLhdLaFNu2cG+RVdPZPXqoPqGfb26s1W48pTkwNLuqbagARZPw60TA
F9IzXoZrb1lUv/dVdmdLywZWaAfuyJlQh6gPmtUAH+qNM1lU6Den4iBGL2y0
ys5+Qp6aGPUMcJw6E6hvRQcy4EtNkdO08Zfiu/t/PfOEegLCE4HR7UKCHgoc
WYDdFVZz30sLAOIoOkVMSBKO2ruDzRHeHd9GPojsAo+pEOT1B3C9v5TSqtFS
zCiJVCoVP+5r4f3wgLLYVyHEAJ9UkpXc8ZlDwBZ0lWRdII712n9rLMb9sPfx
SzrEExgnCPeap6imgj9xq/f2I1Kx0OROdQ3wx4VxSu7rlRPNoXdH900fy5Qe
Hp4RcUEC99Qka0ETtRvdY6h/HQrSMBhwF8IWcDOzLiyjsSn88qayNhas9rxI
n3UTTrtxZy4EeJsq/O93iNNNwhcUTI89uNqPk8a9WBpi1fIh8G27WZ53dKbB
aDVl9Bn44qGPOlVQJwgKBbXOJ7xpF/cynLQ/y+Us1XYPhiePMVNiUgpkYSL4
JPCFG5JkguGlxXJYsv+gZfRl7/xrAdBDRrjtMVgDhw2Fv77FRMQv1fXkSUIz
GXAslQtIOzBj9YOXPkU3KEGRHDYX361Ihgk8/BuBxFcsq5HCrqi3mOE6OaHG
V6wLIf5F90GXzybbQEclBozJ0xmI2pD9eucv/b85A8f9OtPBjhRY1AkbKHp5
1b6X0Qr4YSkudCmHBRIMMEqj0zgmszy/CjPBu06xWzNLxGkkd9hX4OcPO3nr
u6pguyXOTe62UX/SxpopGXkPuSRNZAs7lK1eCxQPkWmkZyemY1uXNgyxDOiX
+5Er1shI4+Ia6t8VwkiXvlyySOrsp3sQMIE0cLE/aAItq5yhxT0Gj1NHJyTj
gaPdSA0+TDYcpepzmnHjiIEy1GI/Ovu1TZNsem772NV7zXVqcIaLf+UJbowZ
ZZ0bncS0CudrI1W727P5tZ5zS58LYSCi8wwFy8gqsPyRDcQHBuygYBu1pJan
dttXNJs5/DqnNJtmV2KXWMbt8aZjSyz9BpgavjU2enuZ7/6raUeExkkTg/HV
Vhw9FUChClJA1xVxuK1bY0jQ6q2vLwK7zprltB5NgrQteLy6huk6x0OuZmqf
N1uQ11IyLpJSeeF51VDPNRo1tQOS8UH+pFWwedF3AUxeHqFwMiSVi0Cc7z/C
flmW1qSEnBTiixXSIz2t+wOk85nz7xAWtWYLjNuYfmzM1rxwoRAo8gxiaxrG
wwKouKNJTPTlhbOgMfbk9RcLptvpjZEhrcFzmPgOAev1V/KbEKNEaZaktYKz
XUBsUPgt9vBgK2+XB1zaGg0svhFUoKImcYCpdkcFVEKEOfrBeg27j2UaIv/u
L/skdMiqkWC2yCaEWub+xY38bc5DrqWELCk11rsWV+URq9OiEcmnQNrsX5R4
CqxHt6VmiVr5oOjr4luUAMR2abImmF0T8f6sLuyoFq/2Jgn4nBXjcaABiGbN
rFpstvoZzz4iN9T9qKd8ngWygoXnC3Z3VM2dZ+v9wDu3CFp8Kd8wTbqOWFmT
3cF2gjp30foQLXFUnseZD//NaxPptdHLYXp+Z4uSkJcJAfmf88IU1+cP3jFV
/+IuNJfmBxly5/t3AgMaQyDTGdX8LsTyUGNjdo6Q3u0rWEoNrR5WCNXQSnhW
ey3Te5KstcAO2molbZ/cs7jbxHOTaA/vaEMAk40GU6R7UtGdpjCHFjvsfWRv
osYbbdl35nezUX7Odog84VdcTw2pXUADNq/chtz//qCyQ9FnXcjPuY87RC6A
MmbYiyN3ZI7chc/QzguY3dkkpn3f9azf472RigJyCsNYFn7SR2A9eIdhijPA
djLLl1wU/2BVWycw21ZfQNMM/nEGIRSxSbuIfk5pnyyM5sndbMpkmoQ3UncP
vAgxFsdWFibMWIwtyupZE9ekqswht1RVkPfndxkykUhaSLB2zD46bmDU8YnJ
ykWydNLOj4t6YF8yZTubrPm1ZVGMBSJ48JJRs6JV9ob5BC+LfAbR95+2+tho
kOB95dyhMZH0tyVrbH/f2mihjig+7pwphCmXowBVSxYGYuDNg3wXwPBaqsJW
yp+rqoEgWwCbjsOd1ymPdpI7LIID2b2F0Ciu2lk2vH0ZdJOrZgBJB2j+ZVEW
enW9jDJJK92yWGW0/v3uDHg9HArj5l6ZDs5QIbcKPslpEK7yh4DEBVDwp40E
OsC5yuoAIr/gs6H6oO/k3/vuWQtgsG0mICwtzpye/lAhCsjjAWXq5i6O3/xr
3qUfmEQzZOyYkjLW30e61mE7vs06sWpn6J9Dmv5KkzjWmCX7R+LP3KJPW09i
tjGGrTYs+0DRntOxGLSGkmtsbQex2+DN0HiZ6u0FALtqgrXFIf4VJvd2Kjaw
8K8aI0n3n0vILZMI37Qje5DU+c2e1cEu7Rpp6zemBBzAmxBDrQwbmSE+hQnv
1/pOme2ic+LhbpSgoXi3acO+liCe973StZUQm+LSfaW3VQjTpwNL0sX6LLeW
mx4lKz7bFP15q8Y1LwhlIJFtTJn7ng/cs78jj8o+i/Tvszm5+8TEx86d/47f
0IObPakzSG+X3jaKEXAmYaWa+oWEVmVUhrucZn/kriyNux9A5+CTK6sEkuZ4
59ljxdxdwFv/ysRnkl/mNhgzm2XA4noDgCxMQUeIEzbdGWmPmfVtfW+Q9quN
fmBmPw7Fvu/NL17rdLQOnLPnlhZ9Yi8UNk0VDbzOuUMpOFNwfW8UnEZ1nIy4
M8fqrsl/VT0uLbVlAxS1PbdQAh3QjC7/ot4ru4AweLseZnqPtSluaeKP/ZDi
qE7eBliTeTjyYNro0DuBTMBAjjH28K/T+g0k8tueXodTYLfdE76mpQq9CSXS
NXwiddReS2Ukz9EkTirh8nH0gUuXGzKPpdPgV/EFw+7ASFYg8F6K08dDB2Gp
VAK2YsaRh1wNKeiznj9ZN9/4tOUlueCYxXAdCYz2tZn+bGZWXKG84oQORnuW
aJwla+4L20E7rFiGPGM13W8DF6y1x+BOSpS55fCF93sxlv6nzezvcSr9KgZZ
M+ArQj7Y8gWVX9+f7uLyqvMMn6NHFzgCMzGnzMm0oxAT9hsPyL/16h6jVA1v
leBYnBbzvdEWzTI9JxFzTx6N6OVoy02yKUIvXB0p4po00+pMyPUl424eZpUy
Asrxf7p8ObjAXhir+/1KHSPdlXz4YhSMDqXrnjgSU5dqQJBtia4ioh5mI8cE
aBMJ00V3K5ldlO2W6AiEFkeHDXZIHO8DS9Cn5iDSHyGUelfpLsDedNk256F9
6wm8lsHP3Y62GqzJuUeq4fS/AtD+JMIzRQZVJPq8iIJgLk/FJQ3cprnEnxFq
Ca1iBQ3aQBmexoFnXqCujn5TrkqqkhcodThWmeSA8T7ltchoC4Iod9Bp9Hd7
bwgX7cuwMajieOo7M3v9ycmETm5XmFsYoj/2Ah+gDClwNbWtMqR71Im7fCg5
oTWTpoW92s6Jht44/2EClrSLN604xk2ML5R45g5hVAZ5E+ptb0Hn6O//N7aF
gqgsg/5GNFeMK/5b6Xg6nTgyAYWUsNlm0ce7RkHkdrgMRszgHqj5RHeiz5cb
x6sziWF423GNlG69CPiQbeNcSY/uMiPAC2i+TTS7Lq7kd1NIPBmAvwI15D9x
XWnFV3byH5lpDMWkB0ToC/bdwZiYfclXRNzQNQhaSTH/xTX+CcaLjC9Xqv+l
5yeunPPt8zrhQxaQVWrVa8Cq0SpdVr0OCmsqUpp/bTk00t4C3q7hRz9Sh+qr
gUngszZsnLH1hxcDhf6GEehPtaI57q9KRPpkUE3+odEIUYyzay/w+pw7zdte
Ap3XE/A2DfRs9j9ZQ8n/DS/0na7caek8Fhr9Y5rCF7sfnV4sccRYzNFXcpfF
9Ah5FunLOGsP1ogCBFypdv+J5wW4qIz71NDUp9kMMxjz0vlAkiUgS4FGSktM
nHF7tzWd7IP3/D+mFlggQ2BQRWRBaml1kFOUIzNO9eSW7z1TAcuWV8E1eadv
WjMBGHoIoOKhWBPoelmPlLIvqjyyz2jQvARIr/Q5hpSoTCr+HNSebczmwHuV
pR8MzWLKOIC6MhkK2JPjQhKqz7Q91uw6otf9DQyrA2bC6P4h9fGcOTIHQDEC
6sgmT3FJyTIUiQwtT+xV7dlEt9PuFHwUQkqo1Tx0o4s8rJZG0jp0FdmK+3Zq
/MMhHsdGgN+AlP9EDhQuF5Y3MbTinik0owQwFC/x1y4CTEDdGPGz3cROgJko
RHcZ3X4YqSrqHpo13253k/eYjoZBxZKNP9ZTh7/2VV5sy1/YBOgU5ELt1VxI
C4/Hjg6wkwt58hTI6NQXz93E8fqGjf3PFZH2OIAd52nHVkzI8xgMIvmg3/QA
nmxHM8kosv5/FYgzFQPxRRgA9NJrj8hzG71vLl2n3ohVdl7RFjmEF35udrwr
GnOZdDEfJcuCow74m9vfsZUQNXRjFFA1HJd9/g/xx23viOXVX3UjDAUKxWXi
t180Tlkrm3Yw+3agI3iG9SzM2j+9CHPp3tRR5kwac6+xkIWnaNxedLMOcl+B
ERRAvPqdlJBORN1C3GYfb7vPTSNlBDUqGUW3CJGggiRU8+dMQxtPIVaDTNVU
/iMzrTJWKdN+lSC7vD2/V6dQOA5t0CsnpFYMxILfP5DhoOAzFgB6YKGheCSz
jPETIWgTeyBe1HsFlJrVWEqEqhozibE/v+Jl+5ci2jy8LaQiqM0Fa5WCDrIz
uy5MTOqLuLgUniHCLHO358ubTgJ1xOo6T7jNlIc6hh1xCYypAiJ+fDt+4iNb
jGM+qrMlk5iUbPE6pN/92t/jMtO8Gbfsa7nKp8RKfM3VCwHYvtnYKV+P1VOu
E0J2V3yfpUyIsh+uSwXjLWgaMU99XP8mvgW8ixKUNIXhRqZzW7AP0rSKw7km
S2A8YAdAs3Ew8/orMURNBdjf1UtF116qL7A1dkI2dxf40MlLUNnY/gA1/p0+
f2d+K+7WPVB51Y40a2+ApB3IARTRns9ZLKlaCUJTl4g0VKY9ff18pIcuA2j8
s7g+5zZDBWriRMBjU0hF7nMdRg4esdUqry7XADLBV3ujAWektqpjZxNDbtRc
JEIcBFPLHHP0XjUJLXQ3CIt2L/VRn8y/3jkgL/r7Y43WFOspHRJlKUQr33O/
m37+IpX8YhBZum46vB2vrdLZVOo6tCSuQqBBeuW1NAUf9XX3B7JfvGuoFkFE
pV0hRHJq+BM6PkYmEiuA23/P68XEQFOquVuR3FsA9LPCQrI5yGVwh2IiU/cP
HCJd5TCqGEu00u/pLRaZIU9oveb4KdmED0/034Q4/tegJI5b/6G/TBaoYIwx
YvafVklFMF0+gqNGcrCUy0RbQBUdH+NEZFG87S6JpKHTpPZL2a0UvEMwVzbt
MOCfXbN4tuQcRlWNVu1/mhqT6Gk412qYypQBb+t5ZKbmlVX3yO12SL4JhOsH
Wzk8NYnNMZGSMdbMWXB+/TtI6YnrEY0BW7U4cvq/EagkGuf+Ak4hQTpRLmY0
o629/uUYJpwIruNeBNLDEpyOKoT6bpH6UDCwX7hADyXxtwUSXxyvgwLHFWlF
lipQUIarE7DyXK+UFrAYlvtywA4ZpVOh0bSreG0CnEAnSCQ/TqzSJVHpI51a
HVBDIxbSp0lkfTeq6gtjNv1ONcE6r3/pgVx5LuZYNIwqUgRAyFoLzYGd9wAU
uFY7WpGzhcvDVep2lXix42I16hMw6NGRKifzzcwXdY+xLyStsbJd1cMpcHq3
stJvJT3BpFQHEatvNCIsNp0VDBiS2efjXi527mHg5Mv7u+wsFLNqQrTepZlD
pqbeq5o5Z9xIaH+mcxRSh5/NYcY2qP1709L7s6585T4bzFL8XVBJ2JfuMUlT
u0/P1X8Xvt99OCmn9fAhxKF/r7xTJKS/VgRo9fjmWXg+ajfact2SFPFIlNhe
1dQYTJr1l1QpqAmhB/U3izSi0FwSPZzTz8kHLFM8lTGCYIItpp+j2HthxcMO
Q3imhLMX0lKtQyFi2ZoyJ3dwL2F7egqZhZpKe54IwmpwMZzu+ird9gD+/mQb
9UeFoduj7ePRByo6VtOU6RJNTkCeP3zDDjxkLsyo45rQSwUHUVp1djwiGX0y
4LYRSlwscJIGUWLQ5kDfgXdn4LGHSHILCNHtIzh7O2q5+KS0FVKLUnFcBOmT
17P1G0BUQnCA71zQ3SziMxw/KPO88sbCJTsDfb0Bq1KmgfiIH7t1ioramxBk
jskA8hD3NkaDeEQKmU7T/qHcQOp4tgcZ2tR2+47HDS50DqdIQsA2A8YIGpfK
xrPCB6HbzrS2pXGSGBRlWlQ5G4UL0qXXZh+F4qKrF6d3aSvhA2t0crQ5ry9m
31/bTFcUMpYwwfOzMfYLaCGPjp/z2Qw4LjqmSDuL/eNAz2aGvy7/+oUUBpOr
QP7mM+Aw+HpSGmt4voWSVcFUcxAYm7INMkT23vMRloCw5To3/qAPMPBmsw3O
wWn9Xe1+3H5N/oL7Eb4iihlFvUNHQmKvY8m1cafKJdCTBU2ngIz4olSok+qd
xttvnS1Bl0DtbqICPsydxQ0o7c0AGfnEf+WU1znc8T1nm1thBe9+L8XSw/a/
QrjRhpKUdyxz11xV0JF2fX2+R/a7W9suS1WijqLdIFGVKM42D6KtxzFscwZh
jkxVdY0rVKrKqM58UGEe7fHe2j7LISGbfsMJXk2UXZhm2GYByj8d+Ay+qBGk
0dACUECzWqVT+WWhRpkp7ns6gaVgXqi36BqnqujL2cNnfgReIPOfURDCgLld
9KiXejIX21BCaDmGi/tf/iyyjs5IHy3SlPwvQyPcU91pVTGdMJYIu5tLy6dM
2bTKR1VNmbdLS1xDzgtLVuBovaoBs9W69/aOiLkpOfX/9lgyKd/C8pZJgS5p
onT1h/pltDUEnPE0WRhnErppmDLuyXMPMxZGpESOIivtnCxzB+xpPIwxb8Pg
4paonS1952I6sgoglKwYBaJm9EADEJx0n6o328yLM5m7mTZ54UmdrLHdMvj3
PY+RvqOXHgZZIYBctxgwWcQ8pwrNxhgjywTQ5yfwmshw2PVcyFLsj9zZ4d9w
oRCeivcycHZ9qSVkto8/qdArBk0AKNlp6I8e+b8I1xwCXpEm3sDjpMFBC9uL
/rLUwiezbPmyxm0gqoQ7JT5AzyBIjjm/5KgXGq6H4RmEDtdM1uEVetAPAK6v
76y5nlloZ55+pKmmI3ldZL3tXnxWx5SqPfLaET+jaKJx6aXAs7uvYja1OTmT
blNFZruGkctrH6D9/BQpn9S58H25iiuaenzWPTksbXlB9SI9IGTm4JlxSX5r
td0/sfYMPXP380qPDQ2rLXm4VejHl9fzAtw5if2oQoRw3rHtcBjgObBYFgyt
I/kntE3cgNOqJJa3J/lr/yddZIoswUR2fKuKX6KUf0MELb6tvmxeD5IQUQGu
zsXt5QG98d8BmsTtlAfoBJraoWyc3unFNrDkamAchbJcJy/HEsBQQ+EnC4ZP
0HEnGOT2865Ucc07X7iEc8T3i6XU/5BBLINdf6QRxsh0PaiVlwneqSCojGHV
vemo5YX7DA4W8Uq86HG0gW25oGCt3gfiNmCnguQTIA790s7UB+RK8wW/gLhf
pnZ3bN8SRgm0zzqudTzQfMivrgZHyL7t0b7UWfYVBGwSNGKb/IM0oVaYPYru
ACgpGXrGZSYYoeFoVMjgFPZUGNU4uWP+s+1/iNmtVWb3WzkxDgQco/ktrfEy
vF7zkWYGPju1LX1qIwVGg925o8Gfn9w4EJWrLGT5zTpJ1wpx52Nh2G4o5ZzL
f676aOzQgmKn3FHSumpg9aVUb1lacyA+BZ2F9E0l9VQ99evxc3+wXgiybTDt
dM979oDTpsSQzJURo5K0rkd1C9apEsA4Rg0jFwWH8YEuBrrGM2GZ6/fKvL+J
+H79mGOaM6h57rnMEJxk2FxjeMjGttSMQCdKvgfC91ILn1nk/u05eRad/swF
rgHMUxBTlULKdYfdj27zX1wees1wui67z4CQz5X768GbIcCXXBBx+lEHJTAZ
NrbnySX64uNK3gWRIi7xDgLLAQuPdxyZ3IDYZ6h29CrPb92sDNh+f8Wim9XG
x9NA6JCTP++7gA+RAI7EEqs4XBQcV/3bwCQhRC+mC4HJCL3Nk+xJQwIFIu7L
CSx65UbsFUgZtIUuEQOAN7gKB1HWgvgnSGlRrazlWkRlvteMNBwQsqh244RC
5lMvOSoVYfXS7GihVfqv/Yuv60qQEZq41QazPFjkPwmij+NUDd2hyJbPMmXV
ZvEmYqeivLB4GDfuyCIq+SFnnDksnZ0lH2YR0n6SuECulkgkbfdwn/9cwkWr
jOlCB0UY4L7a0GbbMyqbejfablBBRPo8PwWuSi8XXAnBXoyx8/ifkjDsCLHC
Tc9nF16NaFbL/BdONxqbtVQV+sOs9h2UOnBVzOx771lBiqISjWY8r6sVoCGM
9sYHxzraRYPOng5HBQioptcd46LoG4hBBLDmsYKCVnswHZSAqYcEYi32nVHR
wgMavflbfILBdUls5RXHoopCVPLuHIqxR9ZAcDopGsX28LFjlSn9rXRgJItg
tEU+mGvgUIgfuc6pVtvl63Whrariai38Izc7cJOV4plWPUs3lXURM2HNklcz
miATKdH/j3tZy6Eb05k8qgVwEOD/9YX9b2Xtu6Jb/pVhNEqULyeU3UxanwBD
ffd3I2HGaByKei0p/I/ep02dlswq4ZE1/n1ToxcQvB+9DuwKNJPoXyqAzY47
oTTdmxXQ2RjB/gr/t+y6PGzJ0FCAXYvrE2Tw75NvTukLxjR9pW0xLM0Ym5SC
UR0PyfMfPokc2kkvQQ7SmaBqNXNQzjOf8jeztHXtFUi+P3SQZy+IiFenEByY
gAm2vR+LRLJP/uizxvq6PsrC9ws38JeYFELrQp2BJ9KYdP84QkWob4UPpqdw
R8NZ/cLbd++oQ9k5Jrvkg43roGw7DyKmzHDh3AkOAzGwniDoS1N0G/PbmFDz
DrbmzFJcUT2a/fSp5xIU7S6GjnjkwcqzzLlC9p78ryBc4RStz8WQDpMQZqQp
7SY0QBlfBIG/b6Zs8ie/2bzIK76RuskLULCikfeYdWoZD8DIHY0e17YBDfMW
vTtC9vRK3DliEB2luVI+KNYpMnGSAd01Q7uxZjj5RWrO9qvWq+f8oAd0OCDK
A5LVG3RL+oSZusxnrhPoLl6m0ZUSOOijgzgjXL0PgXjgMhwebQLu3+9niGFY
8rQad452Iy7aEZhN5WNlzimxhYjz//ocAp8sRnuGEhX6LIHZd/Blohpg73kE
5fTrOnEw8RD5wHtgMR4ILgat1h0rtr8d7UpeGREDDzXBH0Nouwjn8Lw5YimJ
rEbrbr8sMG7QS4nBDot0/XmiV3gwoZ3ZLSgnsUEU6c4HMw7zHjMRptcNST8a
Y68HAD/E6xaqrhdDxXhmQ/hyRpQorj98pwaQlyXiYcI67+ybcfwvDd7OeL69
1Ty7tbnDVCIJYgCfLhqCxL9uloIFS+BJX6Yr1A6SxkS6NImgcmwOuvfHzB2m
87XSXfyNShSZDR0eUiqUg5fC92G19z5PbSkLkBZSwqHe5wiV1pkMt2YkUCPg
rHs3xuu15t4eaoaovjzk8LHh7ql/zFg8h5LOU7utI7fLF8wgqlp/1caKWQC1
79p7CmQ4xfFb8moRjiJQThUaum7BFriW2WxEXDosgPEkVRIN2+2d3H+Q21nn
7ldSyfSfsJ0XzsSV0XdJQEIg9K7o/Nm1BHFWxHcGAIylivRcqKcQo7SFVtT9
/oKC6hgWNOb/Pj2t9S/j/b8qgIQu76mMUixoYUTAHDgIikgmeckelwFl6F0l
m32w04NLiN9qOYg91/gtL3URwYMtsznICNa06hMl6jD9tJ/mScTV4U5jYa+2
hJnmnZKCDRHcTKbZPZ2bhTjhpbwYSPKLdwLnSZcrNx1UPzWvf8k3is0QvSPf
ZXQcDMQpHI8f4tYxAButaopJsLEQF6jnS6J1djxR6EIi9eLzjbDVK1Kt9rDz
8eEsmxRn7ICBwnUV03Rt4v1jH7ZdM44DS98YMtGfxVW6LxZ5hNYuCZ7+mpx3
ggwoJqRLXy4UyYdXVTtTwrViKwUVpyVjqO+qWAnCMeyEmSOyKNT14fDHEmr2
K3aHeFnXkFt+22G/H6+CX3Q4yYF9oV5T0gD1x+iINSbYY4sF45zP1aORVyqS
GI9lrfgqr56ixj2x4uUdYWwIQsRUQiCysxJ+yOzTgrCSSA24MjXCv0jBN4vk
vfCqA1C5xX5WqX0bV+vgb8w5Izl0NtweQI5cJvsSvLtuTvCsrAsM0geE7yf1
5751633px6L/F+V9tE9NCP9lavLHok4oXa/e8jC30iT/TqT97u/1lOG/z38A
aE8CHyMq1igaIKMTGAfs54lYEDY2ZGie17sCvAwjtq82hxpea3hdJHZW61A2
UlirdTSfIb7PYyme0cbCMvJA+G4EyZdKhyEUm6iLUBZolgDHNwcYKCNvExJl
7QU2k7Ttn/cWt9WHlhDhzEkeuEi5IQ2VoKAqOqc7la1/Up8BBHPmtxQY5Z2F
yvAF89qGqCTHLEIydGao9G19SKfqNvaAgCUBKuJq98Tcu/3rja9zUux/iZDt
7dP0KlFWRTPrXFlh3g0+yuhUpi8iEsqXxLlQ/+PIzWIcbABbTvH5Ud70fxPS
JlB2i0VobV2Vn42GxLgaKvxLEuiwJj5XNEEbjbSX5W+QRQCV/DKkbaZcjOOS
LUgIbFZrLBdEGYNfu/6qFfzSPhBeIdrhlb9rif8IWmiBHnQD//pgB8UlUdrm
zz5nJJam9/hGmReK7EXbqByHxAVrW1yGcR1qMBJDmxceEnHIaEcdTBQX79ZB
Jo+bxusE3NUOJRqzKSRqU47Z025T7hvvN107ocGLCaf8VEL+L1NX4U3kbpw5
xYAYR6/sAFJH6Do6syl32OB3nRP6Q3mk/oeDq4KcidTp49XF8jBjrCaJsl7i
Yiv+Vavxdcu2MSViDYAYc65Xe6o3QxY3dDH+zqLtmjZyu6CKfSuAqFDDx14H
aNuzsvqLvj8uJq3GnXeoxgqOtyRQCyoC1uqXofMKdxqnZWfj+VAv+fMu+2Oe
0s+wSeNI52H63g6Du5Lh+Ns7IfwfofX/FNsMycfjN4P8+lNZyMo5eCbSl02X
soKrhItPT8HDHzpaCxnbL2dAdzU+56Qj9i+YHRSe+Rbp2vRKimaBpfTnuJFY
z5S/0I2fznQkG2WW22dXD2F5mjgHmoga4UWXctm2jeX0a0zMSVkk7IepHTjx
wK1NHWPl+P/TS5gUW7dsX46X+Rbg42lwJ5kUEEmuQ1X7TbkWetY15Tv+9EgD
1Mgmgm0XmnkH3EX8IcLVO0sA7yLyc1SKwBtXM5x0aO2Kw1w3vwQK7eLJnFan
6P3/+AbHlspdVgUSqgTZjlv898VJU050bxViw2V8vktG5qJT3AD+3RQt9Utw
uYeeDytEee7m8fNKL3GnqKxKOmX01WDkZMLukMJyAr0ktlX3t9RIO29C3dAi
vCmKDzx08VoVBVIjKhsJuW1hqWppoS49jYx1EJ37Fo6N5M7m9DktnfpnV9P5
XqlD/J1NysBqSqvkniKAh7hZx0U6t3alPgTdsnVYeiPy49pwz3ehhFnomQtV
J8BaNfNNnxKlyt6bKuHK/pCt6ufKS+LLTknfneePyi/kV5e8j1VdWiuwyvhf
XntwhnD+yMg1Qh/YN8xDEE7tmUSM0meJRn7B+Jyy/SOCsLJ2J1JLmLhbRztC
/g6XIB4/8ATHZPKAFU0VN5n/a3aG78kp/ZETg1V8jaOSOEvXYlruOIV8Dnw4
gegZmSMCxJcq7PyT/FCgywMPJUydkcUDoiRWQJwO1TCuRyAB0J4SZs3GwnWO
+8vjsIxaV8SPypQRROx/hO0I/pZPBcVfwinIHGV3DYhWERQmNRJUBykxzBqx
HWpRA/nyi1GnDvBKjling2rMn5tShROp+T80aY2YM32AAI6O4iE7/MONjEZh
bsl8aN/k46JJKxFQG5HGLNv0SOg2mgb0LMZC1nMiQ/PN5iIjzXQaACJH1x5y
oF/JF+de1Oa8OvB9rFT+8uG3MRa8gIJMXS0ykZd8obPeDKKEfT3CvBf8cXvU
lAAKwR9V9xFcXWHQK/OjcRlL+mKVLHfO6wQnC1y0vcKAXkobcw+GMkIuOUS2
F+WZXbvs0wixvBYt7QYi9XCyAyTM3IOGLPAmXx0KeZd/cXuFXHwTmaqlQnA3
/IPN8QNApTUKGygYMYAuk0xuOwy2NSlQ94Qm+cFl+FOcP45srAa0gO+s76Zd
l+VNtMyHr/lqtEE0jySodO8MLUKIRmuul4gL3V/8Ed3KNDxxQlc6cn6Lmtvs
ENJUhv7rU8sIxIzUKjo0MRTdTaJa7RpXsMbf5Ri/3K2ZGxJceXEo2bAOxDsG
7yVfY7JyNEWRGlvkWlk71Q0TL01DaWHIaF8kdHeZc/xJC7d6I5qPQ2C73Xue
ddQDlsENP008VaACNsL0jKBqxeG1cn2gwIZ7Tf/hgbFxFPa6wbBc7K/rhXPY
FlpCGjhKoGYd1gZh5pMx+fmKnzh293kVquTSzlODK4t9mIBJC124ykx0dVxH
ELPEL2MPHvQqdRrNiYZB5dSN0TKLW1XSSfALra9cMXwASf5joTBPENIAPfGi
ZCxDl4cPHzfu2M/fX0OEOsq+yAbCggptfWunfJ9vyNi5VyydrwUF+h1GCIrW
foFlde3ISyq2BSShwMmdX22NASc/Sa4FlrUcWuPsxW2jurnOghjhWLYr2KVx
NPDdKGx7N4WXJbqnBHiGtoPCnnFv5FFaPVsIGUeLrJpb1hzEtBmG0WYriwQR
nLq2DxslFJntaCtzSsC3v1NmAaOQN3d/ejN0hMlXnPyXMtppnWk69bLfLP2K
iNAKy5OyTWGNgaTkBcb4L2FhWiwQrBwAj1eVR3eVO+WJ2SaR+ICou/2Rd2v3
pxlIZTjxDqMAmtiPczqqYJQWxikujm3fgT01UEBiLhBUh37ScS3Pjqc/jfym
J+z+GbjdHWPbnRhXvAfVl3oGxkroNQC0mqoibxzeTO3SAkg57Vv6fUTbg7fB
J6ZGHPwHvWUhNUykWYMBnB+tkT2rMAgzHqG3OJIsUdcM4wb3WP7yEyN3egeV
WcLOkxNam1wAuVo6H+eQ4ryQr0dXcV7rTqiGNfl8ZP9OAbQXJLxRetF51aN2
BhZx3MUnYQm+hLygJIZTdEt08njjiE4kh62lzv/fhommpwBawKVGb3apPNoP
vuOA41MPFhBMgq//MH7Q3k5lPkNHf9hzI1gxAIH4YP6+34Mtt6Bp7iJGKE2n
6WQ0Bm99jRtnvyBH1v1VR5dAJ5OXFSp271yq6WQrLEMDiCbfV2l8eS2hPMfA
eBeMNX1KXsraNALcvjfqAW2agKBbanZ+7KYoClPw8E6cTlEeExLpY3QK7E8O
fxuKyWSg2VAZTCkw3PlUf+ht91G3/6bR/QlX6Q4TFjv7GXyZys1cO5T7WHKm
U9KzJHqp1ZAF5ZG9S7cOK1bApXDA0rRx0P5GGWkR9UHZ+tQgJsfYjXji0Jsz
G09TVjmZWzeA3zVg7X6pbuov9bMET/06lO0OPs9UYehoy/YL98exYybhFz98
PCNHSKL8htA5zgD9sAeVMw/N14JooHYEU1mpMCPJ+IVBbGBWEIPkI0V24fZa
ywRFXcac1D7qGiyskEiw2y32PtC1WStygjauPptiSwGN8jPwldfsyRhVj/bI
sSjCAZyVc+0ByrICqx6+we8fu2Zy0Z0g/zQ/yJjwnH4YPiUADBrkPU04H+Vz
6Wps8U8TJGJKdZa/DLAXl/CLJIVfgsoNGA07NdKgxBZ/uF4SYNtO9bi3jD+J
rdWdlbR4Nu50HefalHNfGA0qXn4PTmrWfek8HLBw+9nysY2z4mMFcsAY1OPX
efrbyfOLzo4GtsN8D8xQXDQPnUSIv+44+cqkWsGNEVe/WH2SAmdKLWrXfRy0
+PRvxgxPrtRs5rDBGjRbP7d1+aiNR7blfSG+GTon9e6U81RHovKVrjhmHqDA
4sW7AIZScsJG+L8DBZ86dMyU9n0F87gjZbdJ9lPkXB1Gryt81up+dzkKkzUt
b+CIcsYOkhB6VGkmg1YQb1D916nKn5AOVnAvZKL/SSZJhJSp7ctD4Y9QxQdR
82U9GQa/emzgQVBglOGKbF2p2dRfCJg/DN+1VMcZ15qVYgXo5RUCYE+rv5de
MFQbEJt/SlXK0f/n6G75cB8iUZoQOh6sp5JSAx+SVzrOtTHiWb0LBVqFbeyx
d7zCudyokgkU9wYGVCJ6zaE1/CZ5PYDp8ERFKj5AN7FH+/de8HojJ3nS2CNJ
PhXIg44OmNaYkNc4fUft7zIKL3TSvYQJiKOoO/j7iETZ5J5JA1HqdDaFkEtu
K+HNmeCGpBrntqvlFWtxyqAFNpe1n7XltnuG9dUrTRMW9G3pHPQGYz3DRRhi
oqFm4w1j0NerE8+dj+qWkbIUDf3MBWey45voSQ/7e2QaFPuX50zrxOAnGvXj
ne9srFpEFoKKvfBlPFltwS9qqlj7fMQNV7vJCTY4RVo5l8uvVL2Tnn3fqJDy
XzzXZTf7TI4bdkVgxBIBYjtA6SFzFDulLjBVGYOV72bTbmskLNLJ9uOJ/2sP
zgFygwt4r20zeHL7quOVLv/j8k63d8v03+IO3Mg6ZI3hjC3B8Wlo3Yqh3KEG
VONdYXqC977mTrSDUfvFGu3uwtYFb75l4N2JyAaNcqJsXV9OPLbuIKmT+6am
YJaHy9vSdTZRShRxYD7qxEcDJ9PQI6j1A1voKVAwhNjCOBnlR7p/R7VrLGwd
4ca2w0EpboanfaurFY7mvp84Sey6V+mJLeWGW3uWrvvVRjZNbYdYxW/hQjFi
I2t6+o5CuJRS44uYNHhFsLJ6TJpdU01jpIR+XVKY9Mm/QKnJmIDNHYqPUjW1
JFw3Ryt+RQtKU/+iXn3wePcFYGyj3djlJWzhfw7xFoeRldPsiVuYSIpI2i1C
hyn+OBk+XlU4jg/uqmgXcTYSephAHTk9JIa52awXl4KlJovERyHY7RSCMtSC
T39roWSHfkEtvWAM5B5UsB/0V5cx2ONWiZRGMbPrbbj6nT+QVM7wBxo8qmP7
6mXFpe0rqNvxBGOA2jmHoKRbT2rnNgkRmqMmKfF3cqe22S1ftpvvIdyTlbmN
5piKFcvQ0xtMTbNqCRQ7uVBrxGrTNDT7kMBFFuHIx2616uVyXTi/MHXL0Fdw
OB/k9/HwCvroUtC3F+QZ3+LxsjD9MS7HTN6RUc+6XAYipK2M5IJHUnjTTGhz
ZLd5nrr4XN3JSj5nrIkaU3iuarK5MnvsplmJCzqogIazMH7fkfy8Wp55aOvc
kYH+a70uPp2bXGGJh86CcBziWVtB1KLAfwSTbubbw9gYMiewy47eJRoEqCB+
INYVfQ4CmpoJnlUv7bk63ky1Lh2ipiqPCWiFRwA0rl6lERiDd++1+zH+MfoD
wTEEyI3XJ1WTem+7UXEHk9XEzjt9LDLmMB6YITMNjFuWwUZeyNm2peT0rBqb
21K90zxspg5/ffYeqchzmwzfPyF+eP+YOrRvQIopEEZC4oxRNPqwYwPKwHx/
k6R5g3bknUlIULlx/oYO53d3nwLA8H9wEVFsTReYPKEAZy+2Iq2keDL77Hin
xuJJHmn55r99i4n7i+64Z3XII+6pFdG8kwMzZrLaBQJ+skczJMy9iRGraD7b
vwqAuUSbMRLkSgr6DurzLh6AquDlGTTtp3TAo435FlmQvcShsg/NnhAQqnpx
oiDaY8QB+XCXkrjIcAFDSyPHQvlKM/cKuyXC5JcIalxhK82J325FInpsc2NZ
sIwGX7XyLzk/wH/wV4HNRuwkRTznWpgDa7xABfxo4H086LkMWA6tg/K2dHkY
zDe/oQPHexjo+djnmmH6FX3WKGs0NFHV3MvOvV10juOXxdLLziDabojOL9G7
PDY0KUgRIhzNLJOS9HMjXATW84y8X06ZoZ1EGhCdt68qEshtJFUcWQJtFqb/
D/LdsNfPo4Wy5U1ipc+O6Ae2jXTZkokuTTDC8QCvpxqJNWdXSHohf4m8iIGf
8h5OOQYTjzqI/70UveTjjvrNZl99fwxd+AkCGWXRDpGNCG5r3WZTi55keMIT
hZ10EBI++e4zBtVX9MQTjR2VRda7BEqaN8S3wJO61KLcD3Nr7enWsbzlPoqT
liwN6b1zfCLrt8MaQfu7XHwd2C/ju8BrQpCy3EmvDQtKvlGckmvS+W/5/wli
TCkkcesYzyUXoVm5mwdaec0VY2CiHqKSORRbk2p/CYpm1nQJN9iwG6lDko9B
o3CevR2u0Ayb3c56+IycfxP0iUgqWR25aovWe3mGiqkHxn0oeZLcq9O1bBtE
4sGXCKFhGXU3TpAeBR4FKs+clOdzPniI/DckE40hcVWajQTc1TqmNj4ZiBuy
5ySwZk5m1Hbb2jUOggJ/so2DrDR//tFgmNDfy25q5HjX3bxaZ5/X1i48xKF/
nJZ88dlSaHruO8+4r6KXIuAuWJQXRJiqC2LhjjJjJVqj0hbNG9IAd2vXc+dQ
hmjU9DuE3mwSicR4XTTT3PYYydD1l3l8XibO+y5S6eG1ZjUekOPnaaXYk4oJ
VQxyrKJdYzvIkdR7YNxByg5xFdSYculz9ebEWsHFOoMIwf9GGnKx3C1QsE8Y
r+9gbaWiBW4kTVpkm8f0qKuBrMKCs4rcM4hLJefmaDygeaTrhJrUs2+r6wlt
+0LzBP1/Wq2kRQBp23j/bwRkIKKgcSlCgOM6QtxZVagAFKqoQlknwmzWrA08
z5+0HjXDRUtbRDOiNTgtW/G499dpSr/uItD0I8IGsvw7XBKbPJ2kSxgcadvX
bGHPWGmvSFNBdBEt+nQsL7wpxqLpTBt1nlnJxuQhGdPGgenx4zvl2bptgUCt
T8w+R7J1oPZBtaRhqEHwKjjWF9hGwa4FUEBvtzHEJOAV4wu2hIYgFZ5sFU8S
PicB69kXPFQHkGAg8w75iM+JQ1aQXykWbKlovhheOUL97QjxDf0Tc2XGGV9Z
hcL/RIuKT19o47U935XTEfPyonlx/uAsd8B+fZWR1Fk3OhyeejIrc9aFQrkb
anA0EXgfhCulqGF+KJoGpJVhdUtx9zInmb9Xevo16F3Sc58JiEof7JfgfsKy
e/W/gWKE6pzYAp08hUjMzpHA968D2eceEtigoYcxtokSKLJ54JWeQUTGnzPW
Zq9UeIoZ+BxiB5oX+s0Z1OCw/W6JJ6iimOMgW9ZQCcYUREC/BZUAfjmOyOrr
Nqq4y3kIRgskxAKQKFg87aBBCrglTsbDsbS0BsL3IfmctsaioJoMAocWt0oS
P7s8h0PkrdWol85LDqtj1XGFULXqkCAGw/iZpJ23Bgp9RbiAyQJECPaHeCXS
uQJzi1Q+AuiR6/m8IvpznbZbb10jgEzMdWRfWVlG+Ua+7yqZarHbWPW5RFxW
WfvTn4treyqUl3II2/YSSUPGx9cPYWHAzrU5HDknxjeL4Ho1HuggSdVPcmQv
EzKqZw3tnMZRBkxyIM0LKHtokIEF2umP4LW58Ccftg5QEVlsGomxm/Ju47r/
memfnInAbIpczeEGggYY9sHtKn2YsdfW0NV+g3F3IBN9fQoxKFxjjUDoylAH
y9om0zFY0HM4gUaJCSVKhUGpvJXkgLhuBUwvjJ2DH+Kz87avgNpqZxN8lUOO
z8O1k0ibnm8iVZCLUUXBZj5BZ4oOx1QQ4/Gkb6WyiDZmcQ/F3jhSP28ojyug
EEqfOfaYroi2gFx6uCIcsRUcUA7yTNu5MLVLzVnOTMjblqJPuCGW1K4mMckB
Kjz9SyA9G0weVcH4kBGZAS4hSIq+aypoeNlAcfaUMWabB46L5YVDVYJ+wahY
KD8n6dVtJwaAHdUEY/04aKKxW7ZDw0w+5zfBLPeIOAXIyJ/6lyOM1BPXv3oj
jjMnpXTnzTDGhSELB93kyCIfkXVObpnwKKqU450OJUSkCCKNJuCKtBT1OhzP
wQr/vSJiU4VM0uwPpqCu6ho800UMaBf8nMjKD8tZX+OB8GGbRRiHb+slGUD6
Jlp+qT7Xmi8asZHK6k7rwOuMQED54lFKqbw62GGZllQN3m0VcEXPRxnGO/GK
ehA8bnteiwRP1Of2iVbDYwH8yMpAbyIRmgOqxZ7O2sepjaJfvFkIHxW27dTI
9Bja32vIfVXg/IsK357PaRlrsafVbkeKo5JX+NM0WeQzHEwn8+lb6OxwmLuH
AH0PLvm1mf2koq97lVXWvB0bFe2b8twSRI1N2x5Ahcrfy1b+95rP0a4Zzctx
79V9aq4Bg1FlQJOLux5e87OmBFoRq6sUnimiHE59/xZTznAGI3WEPYvkIsyc
AxScOdpt0G4xdHioDeYHnZD7aZtQedOGyjkFETHwDpA0xOrs8wWFAmImINla
X5IU2SStfp7DKzYhohEOCtnBvB+ndHew0QpCPhJyuJyH5TcZSIMXxlXL9RnC
Ih5GNHkmo/b2sZL/aodMH52MNumelJm+ELMbB6bgRID+nnASUkI6OnBQf8LC
eGBtSzBfOJw2sX04K5DxiINve6VmvK6nMqaYMbnAgupRpw6TeLdEe3QzwIP6
F552uKRTU0Rz+/IGUcK7/SslfkkDeQzZPjJn93eWWmayxIihR2edNgd+5URt
KKPEWCxQ7M0v6mu8SSiEsmL2OYwvUEZF2LVnKeR6Xa6TmpK1joPStvleAUr/
23qfn7E7iKw760PRn+BCDqwG82B4DdTOXe3xDYG163W7QLrAvdiK3AEs9xbe
IaOj9g13IzaDLgrL/Dxu8PvEDjtLw5rGWj4IMmfJFN0pCD9Z8sM3MSalMleF
AE8idNc1o2pBIlGELNxFlQakQ5p8BTEcy/0F3NDmFJbHeqjsCELl2n/7o7o8
Y8N4HeN7vSCssRlCVmeVLCibn7t03OWfNxgCQeUj6VC0mLcirENbyutBJUol
/pAOjTyo147Gy4tfBmzhncsYO5yw8E/utjjTtIQv//MaUCrB0IlTJc/ZzTfG
9w8FkS25hy9SeajjJTHbFip9ZIX9liJJl4JzYKYV4oHWqCnqPQ2UZq2B9f5n
YSnMQsF6CjNC0h314gKSekwkhedtgram5+4r0MekSxLtmXgMLvViAqr3veFp
cUSlcpkfPWWB6OSVrJwjPZ31QcigsygzPJSeD/+0DHwYDMJHigpW8d//60Ds
49JNqj50AbnUTOh0N9ORNvflKwOFSyBjPPMHxzosOy2l5QPFJJFMeuHzPk/+
87wDyd8eJ3iOmslOtTG9bM0uMjQLGMaq09e1/0FaFUSzKgYRTe1fGybAEcOi
bK3YYAVF0RnaT4sj5H+I7D6ZYX/LCjTizIAemojb8J/BMggyhVqK/PKoJKCc
naM0cTzFdyrsZ1GC83/XY1ec7RgCq1nSFnOqiw9ESVvIkAC7dDUV+ALILMIZ
iSjwlOkBgdL+vuJnquWlIwvMGPqFcBIGXWnhf3Gc5m2/ahfZaiOUqtrvp2zH
kJ5qUn7Xae5/7ALwc97J+WPWE712LVpn/d5SjGPaKE5ECoazUvKIYU63BH8i
cfx2y6vWQh0CwcMT66OUlPMSouMsDWKq1LzWGWVxGSgkMA20LUFumuSB5QK6
qciFVCWlIKnj6vpI3QER6UNjHHer5WVLYEtfC/NOi1RZVXtZ9HbQwcRTc7Ag
j3xTdeXT9FUHwsRCDvlq6h3ygm2us7xgAbbC0GsZLY+YiUC9aDBAD5jYi6+W
Aidrgb5EDqSPgTHl6l3Ps/BgvkVlinDc41QhLXHbbfimmuIy5Gu0T1DucUbd
fvKT8/1+iJNcUpsInVBuLkhwK4UGDiPLDJYMGEaZp5rrH7OpDuA30LLArLrx
ikxD6McPloEUI0DPNGwE0VehxjXX37IiDeqVj2QBM7csFyuWhZvRB5QtCNO8
eBTNk8ABS+57/MUEJeUKv+3mQkAvUuTq+T49rpdg78NwjrBaqHyr7A+wYFkR
TlSVvSi8+rJqRtHfoVVDFPCqVpSh6ULviDJQKg2k6Y4SecRE9bnTr08sef7/
AOdjUXTZ6/2DWPTL6WacXbrIDdLVldSj8C9bpwpiVS0Fe+9vVKTKpOBdEPao
NHhG3EroWHBfzk3ax7yGdTQvZxSkHvEegOOlYqBq996weKFAeMLEmEertFyv
VQdqB08jcjXl42MeJTphr4Pdh5/8/YK6MI5blnhW5i7e2jaLaJD+MzStWUsz
cWpO0ZEqiOiJEdV9uFyg8AslPlAjWf9vgBYRC48/PvLx6U99g/X3zU2oWq2M
c/XaXZFEMESac+lC96bpxWBU6Tp5iOSMZ5bIpkekYtl5S9NlHRYA2wOgrPGh
Zu147hXIENVzeKZHbdwom4CRKtG8HiZaaJXPssKTmG0bdJCdFF1oeg8clWjr
g4X2PmAN+jgtR8xCmx5SgAyC6iec+uUno0sfL08H7bh42FKFtVYZs+01xsaD
OzpMFikFAvpm0K3060ImOue10zhQEeDIjlvS5Rtw8+HsIS9puclHEOENcyGT
xrzb0jq2RaHcUtaDZH0W5Hod1INB3o3FmzNTmrLYFa8UYvn7/KcZCeG2L69A
U+tTFAQ43MDSk+gwopd1qOG3dcrm/hC1VKGFm5KJj2b8Qor1goR8tSDcxi93
mt1MwRTaxMbm2qIZVtggGfB1FSMg1ZmfXjP0iggvVweM3tZ3CvJZrBHSHVSt
s39PBd3kTKMl/3kMUJiOdrwQDbhpnEu40jfa4BDGThm6lz34v4tWissPePFH
N4f/69Gym193UPHewi5KfAIRWtPjgpbld63ymr00QMDRqcyMd3OgAw8zGnIf
ho6fGpKUayI5tY78VFhOtCCaC7+LoQ6+3PNPv6qC83C3sFgUBLAnT9QTRTxl
tXm0cOGetIqBoxivvWmrZA2XDVsVOYCjdx1BZyG0KjRgnN93tiNbdoJEmG0C
Wp7+iW5WUfwBRQ83xeXwhgfddJti/9DKlMl00ZcysdIQbKUJEcr5YENmmTPM
47D42JSqD2+3JYXodTPwfH8CHave8e+n/rfeSx1fnb9vCRY4Vpc+tB4ZDc3d
D75iSDPGqHQU7DQ9VsUGraA5a8TMTzTltwRqlQI9R5PjJjYc6Ft2PHKFwf5b
x4gNViSbnQyDJBDS/aUCTavrO0Ss+AoEiDRJciAn9Ssg+ijEXYONkLTmIj/C
jyqyLtbffOLXZ9sJtShutGE1kCI609k0I2/G9vyAZaB8nv6Zm7l3g64yE0I6
QiHhh4ogAh92B0eZ7VSNCK6ndA63jsC7ywdnHidgvWBxvNdKqmtmc4xnE1hi
BAAH38inoots1uKXRBmKUtStyOW++71/usaKOla+trwn0I7z87d1jCtSeTYg
OhNV7GOmVHRTkhCTezSCivXARqAABnn9rEJ/fKN/GT5t3WBFWp0SYpGs03GQ
Tr6iy+8ZlQAUzw7HkQjp77jn63aL0zMMLAhSVgnCwtiVh7e2pSgknyeYfsO6
l11urx3g22/NU94dPNmy1HNH/FdADPGsN+dHa4Xbh2XHzjQNkebnmUtzJQN9
iykXTFsTWjBkyNAercX/6tZrBa7acehucR3aKkM+U6RxbOV50pTxz+rwvS7L
UzOyE01go3TSYPAwElfiKfFS6DQATTx1Cwdm/sHeONKpZU3XMTSyQrG/AhI+
VrNlV96QhraCQffG7xaLGybmPb7KXd/3LYEKZG6jbB05I+llsZhHGmObKUCD
JJ2A7+9ynTN0fR8CjoevC43hyMpmuxofbGxVkF9ZpIgFynVO9hTJSjRt6XFs
xdDDPcr/rJhEXywHh55YLmkGC/GU+0uW/0At+Nb+qGn8e2s6EU1XBsEZDA0d
DV+AUoTUIn0tUjLAl+PTuDzTXgPySuQXYBRcsphIJf4UPALYhD7DdbAFXMfn
H0BKxD74YG+zi3SsrK5xjnDGViRo16LHEX/VojJedW9Q7d2QIsitKddkcPcb
XXKBVHWIog59LxwuIVAf1Clf2J19eiIS9YypgmM+x2OpzOfq1W2wblswmzAX
0Lu4S9O8x/r8+IxNYDThzJFfF/iSy60F/a9uuYOn2xVMkkPU8xxOCpmrdRL4
RIiWLfoNPhdwBEGgH6O+M6G4ucJWL4mSnHsIyiJ5BBd2UTsNaPSoPRjHurpa
CXjVujww9xTfk0gid1UX7Ourj7eaNBluiH9H3z7uDrEnT2qN4OGooXt1FwyQ
/PUgftnqhD2Aunoc01HXoQ7F22bABkkAvCPJ8disRc205BVVlfFIX1alqFuq
UBkeU8LFnTTgirDZmQNiNPyojdSv2urhQf+DZF+/b0hoxwbGd2/uVsx6mQEU
03dfzaL3YYsetTp8FydXXY6U8uqL1m3HyRkqMfLnq4dmkuk5S+28rPIckir2
3NVBEUnm+Pw/FKCqB+JXqnqe1TJ8gKJAIfK4O150wZG/3Dnn9UIaMihZVtmr
lWUnXb0CVIQo7CHS269clYyB2rZEXv5WO9HH2DtTbAcTcSjGuM/Sk6EhNshq
RHh+STg7U/a5DttMQxfd4ufsYmxzSSbTjzm2EffAcmEYXXJHHDiNVeZRepQt
4+ZAQo78qAO+ICJZqhUiqdi8ztElcD5SM9meeaNC1VsRBCr/LEcD2iudTy6M
NawKdSJNnO4wSYvktNEIC+Hx8Jeix6Ehk5Gtpxt/wmE8fX6LUra5t4WG2xY6
ruJR63MwkSCYQpCgGxRM9i5vtkymexzAvqHQT2XCZCD+u77Uw6xOJdVVJ9mw
T234gDfKFFM2YJybHHLh0li40LvBc8Biy8OHp5AqGUK6iSgiJDuafFN8YEjH
R8XROzI6TJaLz3LzqrZUlasItkAZtL8/Jew3OvlzlAFWyv9Q+H4DsnKMRtZa
MU+XKxf22J4t/xLA03wgU68eBEDx5bbidYXN78rgXUfd282mPsXorzAsP2z7
1o/EqexOZ2td4rGEAmH3/u8uuiKqG6vzijFrzvhlRw5kYnTjoa+wO3H8r+F2
tJl4O3m+v15/1Ys182kqQxqiGUObLmm91AgNP/zIQa3Tbvy5KW3yenaVzED+
r3bMleh/Pmzl0YKP4qlbhkGjSoCwSJO55VsHOXhKiWMYxy9kKIzP/0GpzpIN
KmBL6jJkQ3xR7xKSxe4+eUYf+YtzDzy7GFlFPxYhFC7KbFlIM7QdsrA4fiC+
adzP9r0mJwGLVYwQoIUVoTafQnyPjramo+1JflfINXL6I1N8EHoJr776iGmx
yBO9cqZBIH4GFiu2CA2AgDKo5JJ6G+FInoGvFxaR2rZm+iGc0u+KajPprRof
XZTrdTysOisomKMswFR2QqZ39pUYyJAlzOaVmKo95v9KMs5NnfG4HDmRmH/T
eoWnaBiKnGJLyX06OdZZ3da/aZ2vL1QXeaRMMmPIK3mjabZl0YGpbJ5qqHrW
hr4cnOJ+L5k+wK7YRzKJ3dapCVVDF34qQm1lZarByGhbLAGazhqs3xCja0qR
+tW+HYLjEUBw4WFWQQUBdK3nRmuBmMPbdhxBlQzU4J/TGgYd1bkbXCAR91jr
i/zeFc7shciwdlIppq15d8EIXaYqGR5F0T6wcZvI4Ysd25hC8UH1XE8p58L0
JDR3ZU03g148itZnAzPQ4UsHmrx0n1ArTDD+3L6Sm0aA0F655iGT8a5gFUbm
gi5MMvJUE5uManpgfAL49+Y0hxuIAKgfehZ3ftL7aPUytfvNSOrETXhRxM40
GBB5DAjFPdA8PIWkyagx9kLawQWC0L5aVVRmX54f54vM4L0dSqxCRAgy5ymt
C+3l6f16uSBpU84Z7g20zGQdYRsLfok1/tJBqkCOCYCAeW9UPIBMb7+DVWPG
xH+ZuzpEugN0YrhI0aFtbCYNslmE9QiUDKlBhp1Vx4knFI+rHjXKSxIha6rn
M3hyAWBK7LL4cEJwXSE3VXImQvTi1o1/7IUCoQtEcOEKTFSGX/NxGTgiyQOn
HWOfFmDAgyFu9WrAl4Zu9ZBrF1qKOA8HaUla+DrFrJUrFCuPHo0d5Q0ZOc3r
QKsBG7Mtj4hDdgjEuGGC1mmxprHgMpeq1GSTL0PX/NMH+r5gtjiKjt9aAUJC
zKPMXBdxDs2iLK8gAIH+3VldUZ7wveG/uXINRZvDPqbwhxmNqSwSyNvAI0Qx
YJL8ZszCDEjOhbwCw1OzD9ZTGUZ0NdIyGVZ36qSv2l3J2kGmn8u8nBfEKz8c
T52qqHcrrpO3mr1HbP1p3FzaJz2hHCXoMS7N8xX09/8xSBkwObsw46AkgqTd
xi2vgscHaDgAqx8U1fzjMZagaygBlwjo6lpCyTcNrD5pT+6/gKuQbrwZYhvo
W/EEnEdCFCDNjS5cKPn8qiq2tro8BVfasKt15c0jUNFE/zlZymN307I8l54n
Dd9xe0y5IjN4MFA1XqZY+uH4hz0r292N4vD1KZxETzAXgX3ywHQ4sQckqA+7
nxpcsJNBxBQJAjlqJ6SkIA4HjeWEUMtnvW3pO68cZXcC+uDK7j3d9bPw7BwH
kq8KMZ0cEFPSm5c9cwvC3PM70boEipSlvkthDIBEsQA/2piH16KY6UPrC+DE
XcyHN4o56sWIcECvIUWDMaWFkedcaUkymTIJTWMD5gF1TebtiVIss2GH61Hk
KCzZRCg3zWpF5JhnetErim3zXtlmVzLCPSz3XoUlD0iNAvHy7r/w5QFAa68i
L9jz9tMe6sAptq8SeYzvLxcaCB1QP+SPhic9qrmG3/pngqsf0vFcXgu35sq8
iwRF28bOIR7DuW+dChUPIRQMazbLlLaETdLUg6gq2KpYFaxPPt+Af+Zx5vy+
6vHcIVyNqhuAkRhj0l/UBIVOldg0miK5DhDxFnz/rzL145OAGQOyuy/1ygoi
Yh3KMiG5T041078yEGA9l5H/fnRbGc9c/kjOujpDWhMMhNoa/OxMhQkY1d46
UGQbg15j1zVckCh5qDRGEWtAR1ha2NBanGAiqHMQBri1K0o74vpLTxIXK3GS
pKpmFQvs5TijGVxBSo2gZjldJufq7wtIW4y4hTrLe4SZNSZylHVsHlmHwEHX
e1G2W9fxN9YlftiKpczXZ6G4Vw6AIXVsEMWatLfxIvS70SBdC0ybeKiuLeN6
3vsL+iO3FixVYrEABoaEZXq6VWHR1BWDBz48ehu8TlyQlKnOZa86lHToHxPk
iYg/u7nhkO9AoiCfzhX0wmCm7PcC9cAhpPXjuRypbUMjIsVwlpSEUpj0iJCK
oRp75sYvAvBxJCk1oIzlr1Pl6a5HKSL8KSj5NlStpKmw5J0pFNuEdI0eveoU
VMf+cE4PKOKels7iMIJoAK82UJHAjX16QPt/pHwyiskEHaQUmaPOnSQZEKfh
esMGIpFkYwZN+0Q4qMDeXoMyrtgf31iEqZzwxcsxLaQGvQFF98B24KP4lxEe
BIeynt2WnHPSXigRCqenjFY/Ar1A14unJbk7GIqf7JGt060MbznCXM2olEW1
f7GZUgrdGw0SJ8AeIfwdzc3MG+jABAtjSxFEHW3PwHOmrIHWtamy180s7SP3
0NgUVcNQgGSZZj3htct0Yqljz5ouFcWI/vepvuCGvdnHaQSuZMrQp7mzMphJ
Go3PH7bI7HeHYhxOGDCMcwozJ1jKz9R5qjm6fF2rLwTj3ONLflIYKtFDsGMP
QDJkB5X7iShkJQ67GwsTdyLMo0sINcBWUSLZpAEWSVKsmr3Fp3ijVxhjwXfM
mnyR6HxiOwiI3f3/ENBYeuP8OLl1EXJzowbIP/OvQmu0kvImTMBLE0c37qrf
Jr5eoeGCPtmpmGzgbspBLD2NF1+HPUpDYCR5bS+NZ4BuKFvt6L03l9UvgNcA
9Ev1FILp0xiLcIhdp2j73wUILN34Lbrjn3ca/iPUK54EeZbpOJ7t6xT0pplk
Xs0yphYM6R61tEnh7nkT8ya7F6G+pxuJhmvfuJ5ofuAzfb3/kP4z4QBY1Wdq
IOK+273GVUBvRO3i1y+8IsiQxA6qacgr513PHjpfpeRS6NBkjQvYNQsZbaSI
hBVM8WxjWsbutnUuBtnWVN5tBIbNh3RReTeMeIhdtB4Uw4znB9QulqKM9Q2y
4TKDvnDTXzBSJ61MQZRl+/DlHSmhDks0o3Qnp53xCSx7eT9RpaHUhiGfEk2I
mOQdspvT8LMNQM3dgrXLDnXeI7bp5IOZtmoMcIB7AOAoaBHRhjpHNhs7qOBN
pe5WU1Lh5MB0fFUQxJ1/9odmmiwXQ9Fc6H1CrLeDVEq9mlQlzUKpD/SWqMnK
oHPGWcTCzgrY4OLDJJPLQ8xXMvOVSu1tl/hHPXKXpMKdB22HoU1qVx6Eo8Wq
D8gdCY3DT6/p9lfRBGcQY029iGyfMean+wLeskK07aAQfHbIKmAWUmlRopSj
ldumHF9BMNpUGUSDVsDP9bnd7fCinxOhsHR2G1/z5FbelJIzhe31xYh8ErJ5
hzD7TS/cBcPaKhtxneAWx7YwKK7ZKIy7VqNqMFL2phreRMJ1063GOhYdbDYT
iGtZBxFOuZPNP+2m0EFtCAKgd8P4SsvlRzpMm63/+ywbL7ucdJSV9iHVakKf
FI3dIGDUkgJpArZ+wd/Btlm4824vqHPfjB9YeshvML4+fT4Yqv0mQmW2vUYc
SJlNkAPrVlhFV8z4+OLQq3shVTEVJVhs3Sg5fZMt0vfS36UOjdSAlaoEZChw
a4d7Vyl31TP/9GNcM0yj94xpZm4bSzPN/vappGDK3BscQCho+4p+e1vG8uLl
KQF1AnfAIJH4OfiF8snmHmpyNaEVEwhHxSHZ54xGtlBWafUJYhbteIIdKyyq
AIRC9kaalSECKPiiu5UYzgFCARWjPpI93//IJbp3nfKxpQVIVs+y+vAWjL49
49py+TuQ+na5Mi0NAHrBkou0RJSlkK4QiROJ/ZZ7Pcjhi+ZGL9enZzzuvcfU
yJkZPXak12k4AV5Sw3PjSP8gK+DTLUZCvAkrUq1nGRDjHuWW22SseL/oZ8Jv
2UogsP4k7IFjbkYq5R2OvasRslc0YvkE9o4TMItS9tcWc1Wwo6UVeLCJlGv/
I3f3rvNWcX3/3RGbAMlU9HjiPmXiy9CVruFTeNbUzA0D5VzlQFbmtMk/K+17
wW0AID4VpSRXCZOpfCNMppRAa4qj30IkqyCEdDxjqYA8OUQBbnZ7a+maLVlx
xjmYznihxeHLC2mBEhmbkjNEnRy7/Q3WU1oeuNoS8U/y+bid3vbG/281Vn/M
vvmryhCfVXcUOOImmAKQvNnMy1ogq/n4QVBD2udJwkA0uPI1ihFz4q57w52R
OqVE7H5bZgi9xiM0kEhX2Qkrg8zvvLap1iJolArhWwyAhVkOINJnq7w4IACU
saY19RgUHpR2uHNwN39QWf8ez49Sfx5VzIUENWrp+pMWVLDe/U9wfCJCWEsY
iQeivURQf27eOOORAqeTz6JEvV9A6peP3T1vka4awnh6xRgKzk/yUWDMEdxe
/eQgHUWCmVMdgd3vQTNPLuZuRs6PYNEsbRbEY1IYoNcd4cQWuIj782teedtv
iJfot0dwblv1kydYBM0Rf9V1ZLQ16hnOtgNv2x81i8vuHQeKa3TkqrfYqQv/
hvM1yowprVxI60nCiaH4fS+GhoEHilZJKjehuZ59Nq0m+yEl9ugeTMGPlvik
2wZ3sccmdblrF1do2PSx8IO2QnUBGYF9V5Oyz78T7ROsUa6Lpt3LvbsyyAkl
7PbGGFxlzk+/m/8QAsbSfVk+RMvRNWFXt4A5GLsbg7TpNjePZv1Ueexi56WJ
HT2Cm3+0LiZRAO3Xa6Rv972XReBuIHbx8t7bv9+Hr1mhnGyOMT6T1BYjOS7c
p6RDqZx3ivK42YxMynFbPhsT9CEO9TNVPL93Yi7Unqq4TRP7AbI1T5UKBsQq
vp6KNylT57qj88tZVUpwsvmZPcD5dBsRLhcqLv/8q1cpXVLT1+9nP3DJ8lqO
QHwqAQJkhw22PnnMtR3X2LeYqN5NbTfFwGLh0jrPQzNXhfR3axq7ha2cu11t
wMn/CBCRKwLCyLdqdZMq6nNzS4iXBRyzSdPkxcJm8Je/41l4K3aA4ZbLC6Ee
tx3twyW7cH6zLy0iThdMF58tgDh5ns7cp6TzQkz9++OhgEB1oi4MMgd7KIaK
wThP1buesTCy4/PcMWmbGzgnEUGYbND4on9L3eyyAtYkijU2ITULZ9rBxBre
I0yn9ybUkqLFSuztKqQP/Jn/Du5kjxWGonHf392ztuJlVyoa2AGMLBRKvJok
crKj2EfdePk+kLUWg6qzVS0YwQVKjjithL34zMPthpJUmKI09WueaJjJUmaq
5Hs0mc36PebhzT+e0PNBkZxeX5oSyflEmZ0IASreVpHt2lckltvMikxXhNfl
11Ch+0Ymjr+1Sf9fW10dGuIPuVPbrrZwYJTFjK8Qfp9S9ghrR6442ip8L6S6
1IntI/gBfIa3nUx7A5P8/mnI1tMOynaU9oN6FDMwBJ/1NoMaH6kDbcKT9+ug
jhbnAGuqj/wkUecwcevpWNFrv9JxJlW9KZsoIl/Fa/jNrpddVC3n07wHR7SA
CcMvOAH4Frv7XdZMYFqYwV1fsyW5H7iDJ83aFk8y9YFz9HUdhLtY0rVkO+vR
XkMKYFwH2UlgZ+JQLQ6Z16Cj8tnLA9Za/m0D2VQ1ytWOJDYweqp15UDFcTTb
dkTbfhUe1G5PTDq4LifuM5ywaLJOADD20gFhmg1+atmn7x5yaM9h0ZcCPqpH
dk69qKnKO7RKd5LW7kPQfoR9mYs8gWr1cMPZO1SEHioDhApBqE/KwTRQmq3a
s91XKeE62b1V7YTO+lVNhLUiHmlrY5DNplvECnX6GrkKtwL7Ht3R6cl5QjBD
N4qS1OI8nH2m1P3N4UFAQNbL17EiUFYlTF8JHM6U+BwM4ybGlhhKEK3/CSvL
m6dkkamH/hOV9m8NfFn23da9P/PhIJdY6/hYl3m2xtDmOz91XusDQ0r8Yw0O
4QBVZHKyrbyzF2D3p2ONLeIUCST8ByEcQLhoFrbjVHlnPbmexc+n9HUePNim
x6k36u8KDo6auqhmZKwpVfDiIWvZYehwTSQTIO33cBggSLuhgHs8fs2F9Waw
30+YLZM6aVCWr+PzQs4K6FfoPiHtnGY2TFdOn+xFaj34ZBI+XRvjihDR6RQm
pbo95XCwdmCxP3tIxjQ/nOmdPmZNDKXURgIaXGL6SI9fnItFq6IL8TdAL7Uv
sKhwLPQF8BdstuQu6Yaa2qLKasYmbGrF/8zpYE6M8HDiZOzZem1ypX6PBNcm
N/dVI43z9zJKYiq9XOHXb/UYYfpIDbSfGf/h6RbM34l9FWkq7Wt/idfgnq6L
hjT5vdGHQIY6iJc1RXjauNwmqEWlNLCW9bW2uVbCJELr0o6n69iOjiH8kV+A
ECl3U3nUCdsNSxVjE78Au6jEUX3cRcnTCiNkGgA/6X/p2LYpYLFeRI0ybK8z
qX2FWjsbRsCrvHZ0PiZWXtPo6404Err7X8bLUceNb9Jn6FzxPk1Y3F7zAOAP
81M5C3uWduN/HzBx5k3BKcc88rxY9XNA6hFLhsPxGCm6zFZALDCq9m3L6cij
YeMKREdC2SynROSOLT4raP5MgoWsm9dt3IGz0WrkhelwPzieHeUbhEV5755U
+X3Mq81bDa9YIX1E6NHF4I9XsijdKULhgAOHUDarx/RdZp6RKWV3aaFLjGQx
f4kGo3y87+Ny5Uu7yO0nMuZR//7hY6XUBCWs82nKQMDKeyVcj+RX2c/vYwgk
oQd719N02hK8aBbnYZS5ZEz//wkMEnzJmjDO/JsAZ7lyCZAy31axu5R1ws4s
KJUyAsydZIDrZ3Rd6k7bvbfzjQnbh/2Sh5OFH9Xqn6jStGsKzfJFq9HNaonf
sQreMAdIJaQ88mTSPLuv88g18DazxpCPsshkueuP5Nx8jtmWNyqQP8YPnCOu
92/n05uQpUybwc4c6DcgI/KMf/AH073+p9xgvk0++MfAUqrvW0ZR7fyS5R1q
wQXNItVHq7u1xHnA1VGW0OVafC/7YZC+9LlFXzyWJUMXPUb1oGO3qwmpd6Ae
si69yCqnhFUBYmjusx4TvESSW8MNgRX2r6M4ewdcwe50EvRAZBIxCqS/uHrv
HoWeBfNMLysWc6YSPs9Pal568uzU+3QrlZtiOWyN6PdfGr/Tn6gVKF0rYQY3
B5NINoIDRrV6ILECr2xKE8u92K6VUhj+7jIPk3xiswTTyXACZkZ1HC2JaBe8
jH0xnW7Rx5wnahFmBUUvVuf8q7OOtK1Lhrh+h9hR7xpR2HNFQxpgjwRkWi1Q
9qW9n2oodFOjiYKe0NjulFMeWG8GgyGx63pLr1vEuAf2MgNEO6F6P4kHFRhk
9iwZdjAn++f1/n+o3rjWChQjNl6y2FAz8YR7jU2U61j8bEjByVwK8WT1zwk3
L1ZqwDSRiZKxlrz6yavOcuPHTrpx6Vq7cf8Mylw/QECerZ0kjm18f1/i57tc
ljiLf5LhjK8jmrgdQlpRTG7ImcQdpt3iVH5o4jZJLvYZhanWmzq4XEZNedGF
IYKawcYNu51QHiZgVtOf2t12FsS1sJwDOW62eOpzv2NlOkOPRMYehL0WrNim
CXkbSq5tEn8jqVdpNdVc8xeS/EAEnczADzi4YH1mjKd/BkoAwynzrPJfiw43
HX36/jr57B3I2jYOwVV9cMIiJy4CGVbRWKHcOLYxBmEbgJya0pLnRxws6NRb
AqKrWQ7aH28hoHAp9mIMfqljA2ldwBPcqpfQtdZbll1AEpF37bbuMGzaziTy
HIJK5D7sEHWH2nIczvQyc7L8W7hSZQc9J2x2anIDQBI4vP8uXqPkcAPlY79E
7OC9QGi8/yXdA/ZPn4bep8/bngs9WFVS0I7G1+sJBJAgbOUoQJvks+2Dir/3
/InOQP8p+nHMtTWAozIswyewSsgBAwDJc8FANxmuiYcD/0quEbDqiNmYW3I3
LEkgTIjouNTHkMMD7j0MIUAvizkquvLDXoaDfnLAoMJRZDBqKhy50G0qsQz0
7NnvYvzLY8dMBgHeviTQW2ENCH2qbfRwm61pmmSre1fG3e0GsTjSUi17qZny
YCdXmhKz69EsvJCm3+8THj6rCpX3dEJDsEn3xI0DKLm5iFI18ReVAlt+ms/X
REjTFUAz8eKk8+4mIqz5Qy1Jcil41lSt+3j2Pmu82WrEewfNNfm5kiE5ONLO
VlqOEhphNBicSF4xnuacp1L6pqjVAhFlxsNc6K47k2yBcfDog9QQb2pnx2Nv
cfx+U74QG5WYrNgb0TwlvIWL/LADNmLbylqwOC0Pu2agB33vxqsEou3LV8SB
fdd5+YNemQT21CDpc1c7PRa2ELV470wz6YPpwGO05/0JeueaMbV8b5yVJpRL
5UpjUS90MjvUH++PA32meG66+BcZYPUut7iFyXMyd3Ks5RREU2NBsizjZ2rz
bXIN7KfN0RS3GsJ/aKYz5Cc19gdnERqdrzWznwkOXqNSqK6PaQnXM8zO4hfE
HlwN8MDj2QjnH+5w3LCUlKEDKb6q4U+Y6X0Qeh3HFa0GltNGRSPqURno8TXa
01zhOGZoCcp9MMrPA2bx1ZLUZNL0jHI9ey608uTs7sV7o/rVBv9tDmew/maO
a8VNPuLwJKh+w3eC36aCrpR+2r6nV+NTpArRsESiY4iv1x56OZwP/g+efAJM
32iDyqzE3/31tv1WZ+dy6R0XtiJO3icNfcVZTm5dygqzoEUZCn23IsYGEqqR
WsNanY324y17Wl/Kt+nHuXBtunwxGv9YdLRMTNokQfFFUv90LIOafY1ENXRL
pFJGq1JmvQtgtjpHKt8c3tNr3XcdPu/rj/IwGgH5cUDoMyl8Aln1AReEEFob
0tTTZkTT6pXzSECRqZTneQ8JbCG4HD1mgE7+Z6jklKlN6NHZ3mGivEunoAoO
YwOYRnLMZLXDcaX7EGdzk8F2Vkm6G0h/kgm0tE24BhFDdB8zvxchjjhGN2Q4
ZTkTG2lnWFe3zIBMnGNEsH7x38M99ek3TWMh6xJ7hRc6vTk5dvfh7AAQrtlz
lsPeUv/UD/Ne86SO2ur1zbqQe6PDKqobPGlUFuh4QXDuS/Fo486ehZm9pzZw
hD2/m/hrJXjGktAssNby3TyHq/BR+J2OcyXyDH+GZJSRiDbhcCvYR6ZF+3C9
kOXUoM2n8ffKqNugNQ2pwPXyZbTQ953FIK/WFJpZQvpwvVSsRQu8ZzS9LsuP
STQXLNIGEJ98M+d6noB5PM5YPle6fx8IGCymKCQHWSzwSf+GmgspRGOKugYz
pFT/VWTrDFnaLY1F8dHPFdnkELG60YeIQED+UH+AsDxoYtw9bAIfmFcZGzhp
lluvu7YhnMjPipHXbTnms0VFdgX280EXOiZZoizhKsA3icP5DJVjbIzhqWal
6y7fCLF/L8FzF/E5S70MWwgW0BThQfWlLJcm0SFcMDJPtQhqc4xewnbnoAHW
xmuNfjBZzcn9ct2jgARyTtoAVTvMkhk4RspSKokQ8uW0cW4U8isXjp2Nl4Tm
/kHQCJMwWCnWhSKxlQ9ZaqrU9tNDGqE+4HWyUBs1fp7vMlU59G6AcuE0sEBg
K/2RRMZf3Rx8wJuD86fbT6+/+0evZAbWvVx9lTUhX+LXyYUPIKc1r2m5M0bw
5TkkmHGdAHTgs087ox7rASjcK/saBp6+0NbdE961fKrQNtROcV36Yyh89lN6
2REZu4Rk1i+jPD6plYSKHxyVIr+bMcFrQr4jKonw6wP3TNzCyzuBLa5ZjBTM
5fpqxJQJ5bPJw7UAC7sLr61XAfVItczHBAuSvwlHTcLZ4gYVyGHZvue90lbA
oVByXR8dKnmkgTbBNr3RytjUF1Q7fPOeOfFR0XPYfEciEux3tpO2BhcsrzR1
OVBCrz2byyfszqdfW4FzR8bjBvtA+hu0xgBWqXaOMiFbdWkNOtaaFJuDG1N/
ElLg4HpoabK8g2sRC1y5HjoFzXh5jXw/RjH0eXlpLcV+ZuiT1mKRFp91GRGR
WSZ2vJxSRWd0HXvGewSk9jyS/Z4PNa09VZt3h6OzU52yzrSkeldIUz2wm8tV
36+chyrbqgqBp4ED0ky3qtnuNvW6gHpmwMPbsLXOj+dFiGdcrRC2IJgkP2tW
6LYfU0glcU8TUQqAvjzckUf4pWT04cb0772Kl0VVZItznqqmSBtOLIKTr9En
Snzil4gLDFeCqYyHPSKhqHtZcE4hACbvUW/82wPIqnFpmjpkS1GFE6qPF1Tv
EPs9VWrp2BI7sq29C/UUlugoNo5Kj0MVDTyMDRK49+I4QDZzfnRys5VLGVke
SlGaRfXTsX7NKk+yrExp0FLYmFafvU24eTTLBmuwz8Y+5kO+YlLbceVpv9/A
jGyTPjFzTuoD4sMiEB/WiVDynafB2fgzN/h4GxHDbrBdT5fbPAkmDRvQQR+S
y/ADOl3LL99tAvgNrWekTmEmbYqXkjco0BojnXssiH4Iu3l9QlhFsm4KuM0B
whbDP32jazbyh4h3SIsttZf8F0kDkyuyk0u4X+qk06A++DLIOKOuvJKV8fv4
KXtiWHkZc/c1Oonw4+XrF9sGlTFxzfF9NEQcDf0ukZH42Oj+MX/3S7/KJDEF
TGNkahHWJkVNd2Zx9+lqJ7rxB7P+taue7EaI1boUkmtaO0i0WaKLdoqup3i6
GyYek/DBGpB0J3KrcJ7TBH8IFXUuO28IEkzd/9bgCa0ke0u58erNAvsWvjFY
fDg8ZakZl/N9Og/BGlmJ1YW0Fq0+kVXKeiGX8sWZ37Dz7uLvalwAehlAXswJ
rxAVN+rhOzMGj/B4MagMi2yBFPKT6YksaDTAT/n4wqbpaP+AMQoidJzyPiqC
decAP6bqQRYUfV517UETEu8l/WkqyudOEp+r5LuXyji0dJQF753i6dNGtOAP
k985y4+PZiQq96NEfVhd0GiRHh2huFzjWvqHKBG7RZsYOOq4yRIsGTMZs5Xz
qdCR5/z460j8p3Mz6ktSYlhWhv1Viady44UVSzTNHcSsLMCogiQGsJMlllb0
SLGAMB6a1Z3Suc5ORcq/eUVsAaHM5WlumI8UzEoP0X4sRNBnu6oxuo5s5FSD
QQuYdV93vSByinp3T7f/09UGUPUy+Dk2ZRF9f1LWCDPW/4rdIn0frxBzckY6
6xjkVt8BYxWmiXnvKhMyYqPFGKhqvtmst/m1gfl/mRFWYDXB5iOiG8um0sON
aPWIFmJm/+CoOqrBeKPOZ27U2oQ3t/vivQQbtk1Sd+muox3qGqDJbz7Rvoxw
+3A60i4CWfeg/muDVF5c6kw/qqBAw7AfZONzy3J+DO8kzck2hYXE2+qV9HUF
IFY3xhVFR9k3mtfHX8ZNlN5NiQEQGmAJEjjvF+HYvHums7HgZqLyzcJ6uw+l
iQrdTJTaTtttuHhlVZF303jnz6yXj/4vrl3hp7Vzki+aXq9o1iVixukb4Fgm
cBUuUbAaptBaF9VsEfSUVL3Tr4+gKVugBuFdjfD9E/8nFuntifvs2AsFixvG
iFJigwkmGEsV6BDisaRFUltJw50Ilg76Mdtj9/5vV2JdcPpjOPq5yEVzUXLD
XAv2dyw9FuRkMGJk9MTk0XJH6dEyz1KRYTNM69qSaVWwEPemoJi30rtzhN4Q
SGJjX/Nd2vixOE6qaGiHLzyaigMmromHWcxElKsxwL5rJ1awVoFQvN7Jmc/+
JgO0UqkQs371bqywMSPunCJFCi412sPHDQLUe8qcormicWZtvFbE7FYE9CLM
EM7KSV5F8xOLKLHCovE6fnbYkFScbOx/7KQZjzExFRM+Qtq7r9qaHDFUSHOX
g/zhmdBOLLysVhaUrZk6k54sHl4QemAlsrN1jtYxdY2DiHCWEp5klMY0GTly
ISTQduh2uTH3UDxIkJkB6Gt0icNeyJ75898P7jo1XRDslgJFYUCmoIcKofvn
DnQM7MUc7GINrjsaNnbg0mmTC5Kv2AiMMCpk49X7oKX2SNTUGQ1DnPoIpHNw
Z5Fj1aslCr5s5xVTWCJ+sGL5+5HTmqIKXtdB2J3Q6Z6ZA5itBnhkjw8xFhg9
VC+U/iOZo2VYTTYqMyfceRJwhoJpmtoyVYh1AJDJn4hsgYBFq7f+8de6RA1t
nd5N2Fh+81uX0jzaUMS4xHVp1VuX09q5gAa7+3w+RHb1XJ/YHo+1Dk0G7weo
+wE64WURSscyrzV58/50nV8jfRrjh5utlzxZcxUEr2l9wVNphAsa57/ZQchp
Id7PXtSVelWOAI84DrOh/ACtk62Cv6Rip/THcUTTuJE9UABni8kqtgHiLxJD
Xj3p1JESuDBBagHlRvWn+Z0LQl0taWwazbRzK4Fn+9PY+oCL2NfVGQOepQKv
JJDFmiODmU9vcu+RzE8HaKn/77I4e8q7W62BccqQx2MW9JZg8f/7ALA/uVPt
YBd4ViMMjm0w3e6V3pQ3udehGOO7eh2D+KnYAqWwiUFWrbF3puQ9qNXP5TPO
t/HqYM+ntFkhl5rXXV65f0rdHajSmtTrCS5EGUGjEX+I+Y6JvOuIZQGszwge
2pNLW37IxGDPKZ0m/eksRXkeTYHyOCqakXPy9cl0soHCNy7ekkh4m+m1EIy9
o8INTTaYufr5f2lauYGX+meFSQBMhAzFmJyPgy+rmiar5ZagL/WMJWeZX9RM
5+WWmIfcj2X2YCOTxW3ii3Bwtj4vFue1WNfH0YF7YVpyYRQ/9CtmoTZHDIAa
SouiXMRcztFH4QhL5WCotnNT1p5FEeUJlT6EPzFHNmvET8D52quCgydDGaXB
PanFBngyyfWotjMUhjlIN+ZW4KRhU/A9eAU8u/GcgmYWsyZPUVCQOvyX6KvW
yyrsrk1oLn3BvNqIgL1n2CR5G3OXITssqsngaOccD+STbdFl6WN6m2TlKO2z
rEIQAd8Qz/Q/hpWkPnu3iC5cSKsitKO6Iu8+Xzkw7M0YeAdIj+e2opcllBsA
BwGHXimsXDXNzY70mfygf+BdjqJHj7AaQN97F0JIV7jEbpyfRSC961O99wN5
8LeJwKDfZOOBRPYeAIES35zp6xa/uk7DVEeGVaMcMza9K5ENyhafF/6lf0Ga
fOgru52u8zr0XMkcVVJT2f3WU0G3qNhpzUT+jDPLp2fvvv8NtIgrUEmTsw2l
MW9BEh/HVoUubmDPDEBo8MYK4ExmK5zHxOy3XJqls2lxeFigZrUx7IVoiCLo
1LZv6PcOObkIm/NIFM3ASyM77itHn2KefqUso43o4U5E1XchPJdRw/H+gI3u
Tz1G7ysa1SUqzPzGMuYjhzkfBgBSd7uhiaCWzxG+snCfCGtMqueDXIbfcJVU
iPWl0TI/V/41+JsPKPKZ5arS7dany64WA6dboPBHq1tEra6BoogXKC+92LD2
ZQPBAn45gLuhkSna8uC867FyN4HNJ32B+o2F7SdS4rbayu2RlKPGnWLVfaoW
Sq0jqHEzwwm/AHUfwFEKo4NC69AReXZqud+KxJcUmdGP0R+7uDAN7iEePk/E
zAF/gYoPyYPSMwSm7W8BaJ0C4fK16cYgp79DVdCESnTpmhJgHCVVpiGpeOe9
dysoZeT2A/fIAcMo3Hr8MEX2aF70+iFQX28Cyn4/+gj3QCCck0nfBdoEPv4t
QAgYEfnPFrKqX8RAF/ZzibnA0SaXRKlPtt02DaIB1WieJjqhLT/4mvxQ3kX0
ulzS94jwC8pRBzcLYixCI1S9nIJwf2DHnRimC1HCjKVoTJp62ZRPfw4b/rvK
NkPmvMr9x+pyih/ZUeMF4ZFouzPahfpfzTwnfA/uZsQXix9oXa9VLtCEjwWd
byssYDUtFkvGEB8qdLEySQPRkuZe+kHDauutrFVHPlv59+1dnkNCzRnSct4B
geBvJMGutc7xcJ70Unfybkh2czz5+NKyV5WSBMa0QQ3DAFfnS+bRchdvpTD0
eFU6JGRSjnLLuO+JF4CaBw0DM7ouI+SByitEPHvuStvhHTAp6EHv1Mf+Yeat
yTT81FJhM46KLYmL4aqxuV9UHbrUEE3nTeb50PF2zLcLnoXnWtylf2mR5e9/
Jsx/E374lLz/xE1sxMgI7SI/EXZp7j1JTm4QHpC/31uGtukAhwVbAawaoT46
hO7Fh/qw1su7kkkYxR9ELXep41+swwNkn8Q1dTPimFt029iywk2+9TvUO2wy
xjOLfyuK3nyn1gRFR0K5z3R2bM4G/X+yq1vx6Str1vEjxmfUKD8CBoj+cUR9
AWx47TuzJVR8dNz/JqnvP2+Qas9qlCbcRVdW8DqIz/d8e7QYrwl799tx6N9N
YFZ/5amiS8rbTNVobzAj0KmBpx1vEpfLUfk/rlSQgSgyX0JyItHwfotDFaYA
WPRyFDHfuqtur+syejBIf1Fs6Z7XxV0Wqsd2ACfnLD8kAylQbiAIOUrxxc7Q
YtK7nrUfqx/7uDyC7yh8f2rPJDOxBKSFNmbxy8gNw3ZbSSXNGTrLdwOTQhFu
X+bAMN6hI1DpLrLd0WxkKLLrInxwM6E2Ayt/7uSBGgerUoz1/u7ubg2o9gSK
xDcYQXkGh9A4dICPoTdn0Cpo8ngSlOVjPEMg/Ao80mc/xPyWeAdum9vJgjGU
Kg4lFiMaBRRvFwkLadtJSjjJyj4R1bcyvJLk5lZ8CC30xU9M3hNTM1H/m3Nj
aG5PElmel7EB/1ans52CdeHblTAQJfgOUIvxLtIFwBA09q9VQ+1CQ0WJ9qeS
6pC0335rlru907ef67eilMLpw4u0KOpnAyNRtdcjmtIMbW7GSOHomWzQc6xJ
HkrfL6Cw5McG3YIZF6TaieDpQ4/ZRLif4mlqKn3YXhwcW5mUFFjd/9RYGWF/
U+dpoSr91yDk6/EwnNDb2xfb1p3ho6m81/uSjQfACj703lU5Co2WnLeSCBH4
m6hGFKykgf/o6i3crVr0sGjSLqdlpVddD8cHH83uxQfPpHEoHveA9WyqbW1J
n6CBru1Q9vUa/fNEro2XlRrQ0LN/DBmMwyiD4Jy107kGQPrPf7VCzfp/RiHa
4kbihlIfMFxEEpACDg8LhT6qw/yqxLyTb/qoXCsuu66e/KMhwyQpMuETo6m4
p3s4gpb4r/bdw+qrddh8mDL8URJSMDb83KK+oL1N24+c9qvZIe+6E+rpMOo/
fVujDg+/GvmS9qW2T3ps3tCGMipAch0jIxD9pyE+pDLrSGjfpajo6c3IH3PX
L+SwkDkU+9vSgnWBxOBkisORbFHqgmMeGda5h43hti/aBm7IbrkYlndmrqsT
L/dWOOsLH2Q3ucQbdPP7pgJ5EQxd7OMHr2zJndXxsHCLE5HVi9mZDttaU2Mc
d7hdpbtj1v9B1GnftnanF1/MQmzbfJBywHjXUwz7rktNpqn/N+gFDTDQjrLz
buwlJaxocyl8QPsMRlphHzwlRO3sPavEgL30sMQuuZDj4IXZPsV1CCHVXlXH
CaRZaD4iaWn1s34dGxy6nTmwQQ5TykYkRiHRIym8z4WH6y4A1Ys41uyzlM2o
0JrulKslTP2OZa0NGSVDBj4FCADJElE4ice/B18z+hvfyNsJ9fbTt1cXoSSv
uSxmUdhOI6n2onYPvryEKG3nft+KBO7o+am1oZ6miNiTYY1C7kbWFuxXWM9o
Vy6jtyIvpbMZDH/wc2n4AL5ZgeJ+aAbBSWTHQuN9FLSmt6t8oa+dpbuQqNQD
SLeZH4b6/V1+BaEqJBI7FZP+i4gCyqAHEb+n36BMFGFByTsbdUykfZAe75Pa
e1ZNAMRU2ovIzPwOHICfXShyNf6N0salni0OHhTqfoxHRPpdT3Y4WZRI68Us
2PXsxOt2wDfbZ4HlEdpSooCBszK/ubsXGVyj84nKeCSUJ975BK1X1zuwx571
vyuPEzgapgBw0PU17p+Rz38FxhFWedf5lP85d2zU65mUG5ymtrF8/wiwE9up
LsPh4qCIfNG7qaUUuMJrmdNIP7EhNmTmZ3Q8lPVgdRl/ae97j9ae7WVgmAYc
86Sr3S+ualBvtNTegCXlG+Shhm8IDApfNcK+Q8ItgNxfV3EyOjQRf+etgk/d
Hzhuxs7nYx2Ha1AggY6PLZ2BgF140M9YweDfyHAWwNehqB+j73UjNh3uWB9Z
PELuUI2t94WaKOy81XVQ3obz79yrDCgCHQEb8LTqR1iyop7lHqvdXz7wGk2+
55D867V+X39YAQqlxXS7Zl5IvYC61ixX557ZarlnPLsQqhsInM9+dywGMmhU
D5HXPw6DeqHphwHWZZUv6ym8DS9ZylmJAdzhh7NqCp/uYlCSm3rtptWsBU/O
jLMc6kOTpJN5YTgGv9HalTs/Q8PJaNhoVnPFGrktShTyAweI6l7zkKBBvYf6
YGJEjfbg07iL7yTd+uGJKKh7aapVoI/hl/2kJcsG2bxZU+FkpcUPkavb/P2/
Ln3nupR1NkEgVuYffVrZkot6pj1Kd69T1EDCFxUllV2Lp5E/IqG1VPw7L8vO
IyB11A3Et5uq/jtVHulDGqQtSqAi5lVC/Jmljkt3dayAFZ6rl/vH+OuWAnBN
ti2YJbOB4qxKA+2o/OfzkUN3zXmFClu13PKZLzf0OQmsYocF7UH7Wpnc/vMc
uKNu72YFy6EoSkItr1vvKxWmdlkoeBk/hINf4p6IB1YUGVta0ak/txdZnaLE
B4s/iTMJiVZT7WESHfMR3h6rnvXVUz0E8AlEzv13ojFUnw07/8mtJThFcpEc
a67OZ0jvmnmzsuHIRNo8/GRdlKNEErgpz4zYOEuRIULweukOaH6GPOIZK8mi
wcKMCkFPKU1ClPW1siW7py8yug42wd9et0LmuqJQkjPj5mmWbsDe0u3ydyV0
+5cmHOXxV5zKixj78cuK/RjoVDkIIAh8QDAuTr0hF6CH6hnE/ibWBdSm9QqQ
mjqftgTI0PVkQZ+oxU8YejAPHajIdIVtJHr0kwutLwOsovK+u0r08SkgavVD
baDZ328L0CaUsNuIKRSs0DqWVikTRHjyCSG7guSTdwR2oQj3vxBU57vdK9ad
HgulO1bp42fUjJVWuVFVIgYz9FLHPjtu8nLdEC6ZVpNxfD1/xgy6THfHKysQ
QW0SJdwusWQ2gO6ZXsKAr8HxQYOj7pkWVGM9lbZGdo+l8Ue05z5PRsM6cemE
28YnxLTA2zJPBqL6nmTCiS9RviybVKyPvfvFIDjLPsYILmmTt34/y9GIewDE
dRslu6aMWirHjY+CzegemrjyajafBLvKbkEO2mw3A8+hIFcrNO27riJxXJVS
+Urg2jHJzwHyMoerVKXXSRopZ14iH/tbSn0PC6z3+rYKKO26M7JDiX0q7Z0m
3YsyvRtzjkY4fhT9YdFjtRXnel3WShI+3hEF2gBWvUngskE6s9EYrkW2L0SU
QVRF5VI86DAliSl1V12o1ZXXBgkkf5Nx93ko2pVb4P//pzDcTENakzNVIqMy
dCv4a2sANjHSnBFW7TKBvEQNxdSvJr0bRgVAKsH+yk4KWeq719RHopDfAB2u
S1Kbj3lDVwbLbEnMJIi2EyaeDKbitJ55cX1yXp5yLIx0e9o4vU4wjkyB1gdX
llw+u5U5KZeh5795iLyjh67seFqcsFE+gbEKLrrzyKfllmwbNcajHTHqhK9a
VQ0Mnjd7W6rV0K2e7jaD51O/oZDK9z4PyC0+nxCQLf8dwYMT2IqinoN2TG/Y
OASQs4Cx/q4ot70c4R9VNtV2Ew2KOolXPb5mng7eocietQNV/nJmgOe/TKKR
MAVzoTdBfJsLbfCaURvPEqoAV84cr4wPfMHJZQMwhBLLS1S+zAu3PZowgutW
RJP1WXhKu8aHZKuhbsKUU2b9XD3TwwidfiZDWHWnyV/tMz70Gmu8YbUbwoBF
KtbeckWSaTFk0pdJLHYLDGZfuoOyO8Iv+DJplNinO6vNPU947wl+U4cvn96o
xwLPwUgJuOHugtd0Pv4Ud1RiaIrar4JHBUQZ36PnYiPb4ZgbLjXvILAG+K7r
SjRHIXm0VYkawaPhsoyC/rX5heaEP5mo0udMtVRoL3p3SWS1HSBj5/f1jgkJ
9G/qUe38DTkcM81ZHNtJ9csji1EwsoON+PBQdghGbMTfk0Yd4nIL6BOnVOGd
Tm8jh5O9CiStIrRqxwK0U2RV27FS4l7Olcp5Pmw6F+IW+rsOI2x//pQZZAqm
P+8T2266CN2lvEvdTaeVA6xg+WGWScTJOOtx/D8T/7ex4tPeNPXOmyT+J/vI
WBe77Fv4CfVsX2kjZrAr+OhP7Oz7ZylPYrQHBq9gy5W8xANAMiEtu/R6oN62
a2skuGlfKfbCELVupmJsleDOqS5919CIEhiXtdB5Ka/K2655c3ieGup6Npnj
YYdan5WsoWDQ6Xn9XQl7v7lGnsdKw7jzTbrwfg8mkGXzw5jsBkOSRxwZPKiS
e0XRI4xNK2vup4eXTmwmhzQnERyhuS2yVSDmE1BRHSdmFYzBGAPN/rcPatnR
aJGl4uxwfBG4N7wVm+p1l/WXJM2ECx3D/9CO/e6RJkRE/kQP7dtYF0ZhK7Ob
9mS5othYx0oM+wp5lCL1NkeqRoikRzoTzb8olpLFm9q1sm5KfJGe8VAV2fq3
//ZxD02TZgKXCwEWX/vTmIomNg9AGDw3/ARuVhaTlG6X9S/K9YhM8vGv3zO9
GeUrUEbnbueyGG9w64eemKiAAWnJomt57uUtgBy/+56u5yrf6Qx2qFAJsh3A
CMlx0ptZhJF4s59pS1eNYwxvEwaEnWuNjHh+3TL544EyPDp8uiOlfNKxkMUs
9cIomNeNdU2S84JLPnmIsw1UTVXJ8tO0Gtpwa+Y6r47SE0aHmDAi6DjL31Gr
3j5JvMSDpNtJaKLoJWtGakefz94XkzsJqX7dn/3EA3MW1xLDbj4Ujo1fFHF9
AG9wCOCUvvdtmjCwLfFxOUPXawMq2YdIVYsKiU9VSa4HMnfUbGmItN9ys4pK
bM1ZX8fJ+nz/B8YcGvPhVHVUhFfS3xpuSk0+vQERczv39+rl4mZvHqlLm2i0
a8GgDjAKMfrKN1olLTQULFvVwrJi9un+vEOW8qmnQzoVC3+EmVg6bjyqhiWU
7qCI8GSlBqJ+WhY0R4aD2cmsXpk7e3P29qNmWITCeXVoqVjeRFRuEOp76zQi
vglxdCnQi/ppscUZJZDb3rqKGheEUFcrDU7A4mtW9MwbTOkmgvZchX0Flvw5
MosBAX2iu2UKn02xIT0hc9ZCpFfPbF/gV3BSGRQZtzkC8UDfaObGY0b1EyzD
3GYEzKMKdqwCJDw63bJEL2Ikf9wv2S7tEFm2eHfjsMoNKuxF6ckwW/ry9bGn
hrG1WlPjPx7LERHOwbYHI0nvIR35GciPAEMUm7IR50k7PRQxME7NMVoDSABd
0CBDzDqqe5fwygSzAD7SIkFTxf+uQZ5UL3IhCcIdAAuNkNpHoHJlIcR5f6sg
6vADv0NI7K3WnoxDx8SO5ORi6P116C89dl1TPMxdqY3/5mik9TEN5TvOt9IF
8rWV9OqyUXZon48VguFz2D3qYdxOQuMOIcfBjYnMC6d+SLPYv8uUQ3OKmKTT
RnTar3zfpA441tfncXo+ZF5Wu9F519RBkXC26/gmtxkP8Z5+ff7jkL00LKQ5
elKw8BN4MKZsdRiPBS2w+37KP82Fx36fXHCr921SEp7kru+aHXGZoynwqcH2
OaarMu6K2RrKYqD/4oi+u/wobr/eUiOpF8kEAW/RgC3QUZLlGZ8HcRbaVCKH
Dfb2PXdRpnUSFF/suthvBmDIxe4vzpx2RvVXRB+T1sIbfb86qS0STV68tHaI
AdI4kIlBfPnQ0C7fLviMtRPiNqS295FtCEr9pEhpEVYLa5TIFzg/WH17zS/Y
ykzP6gCP/jN+cajAYMv2Lfo+QobMqKwexNLYc86+Pcj6YtbGIPpK32bvvVNu
xN6LDBfrtsIQkvdaxsa2nVh/gNTMk+ykcHoVNmiCo+SfH8GGiPmChsXKuCg0
ZKkWP7ZfAuxfEm4j0O1FTAPI5JNm0hBBlPjVBR0sB6A8onM0GQWV7M5vs+so
YQPewTFDMF3EAYt8KCnrQf0z4qkTbrz5XHGAXk3ppakZNeDiRDppY+8yqQfY
uLxuKQO8V4EwrRtZFzqtBJnkQ4OvR0RexLNF5gcUu6CdqUGWXbwpnibG7fZ/
opxRkPuNRaOWespxgioZQWgB8tHprdNbVxFDh1F6Qv7Q5VQqhJCWxk8YYS9z
JYcRKwvlSoAdMo2BZDw2fP7dnfqfIuSrhGK7IdMH5xUOy1wTRFLFTnqzvJ/Q
X68unXtjJhy43ggR643JBaFK8fjxou3txr+SJHiAcPAZ/ZZzSz3hckUAcd4m
qWu90/eVPQUOI0Q1IBMkwGLhu96moSQR2+ILwW7IhSCPGfhtTR4UvxZMOR1I
QMarNCsLbw5S2oPg92d9QHwT7iYenKUYeANtwdHMsz0zlR+Vrwb0uZolVcjQ
WwuBn+kPhiTY3jLQOQIjGYiz5i+9RR187YnauYahviR83ac5gWLoaZ2ndvg2
+kF4uBEYk8lqEkrPuCiqzuqfQT5zx1IyjUYkDPpXbjnOkqKaoa9la2IeRAaE
MU8Gq/tnzm/gK+k7JcSMp9wPXy3E8GR8fKG5ZVaImEalOfgphLfsBfiG5CNz
CStn8BewfTS3pdv0Z8e4pBgqh5MXmtdLyVnyRHgccGbIEbXVz87PWxfeBlsl
5OSqXWL7X1zL84EBJVwzHH0kSpQ/3RDdmdxRl4y2rd9PXubvrzlqsc5rZQq2
FH9r5bBCGy5ao8WBAZrvnbM96ss5P3lDt/fUJKU++iqcpRYdnfuQWKQI9GQ1
48fe1FTXphHAPnz7z93kln4a1XVr1kNPjfyE0MzDbscxBWl0z7K2YWavxTqT
AZm7i2ZKEPfJ1ARUjEL8hdcBb9DaXmM7hMMaUmvu3EcOuIHeSOdDPAO17MjU
ZzSyvR82lAUENN6u8GTsH3uuZurAzmnX6IkO4uSLT7dwbwVGAwBZ09AALw/+
0Hf0hXMUXymNO5esJuynHsjpZ9TmdBsfMde2o7nzKjOpvDhju6gTmgAjK8SR
ORXUiYHfv1RoYdS7Usdndvedcy9w5yNr+tMszQbgrn3z7ksni/MEBfAvEdve
gHhi/WR7UgnPIQtmaR3Nu5/6JTkeYmP8Fsg3pZgL/yak3+9DvUg870OLlJS3
RKmg6UPUdpl5wipqzMCkwB58HCF2xuC9rHFuX+FRMF1uR/BAuiYeQQLvtSKV
QdXSa065cUBrA5TeVSrhNds/UJz7D5toxr4EguPMk5ANGslWfRdZdNymkC2a
4WoNFOiYZc6U2itlZsOlw5bIwEFrMdr621DgLf5tmlu+fo0hJbQW0oeqgLUy
Q4XZ8Rjq8ceYaUz7x6p/HWaSryS02VKnfGfL9XNu8Q2+L7nNOfcCIrGAr8Ys
8SOLq3GO5nWkANqn0XaziuI2XgssM+O2l1BzVqM5tsqC/r6oQRevk2lxn46h
uxr9CUGVgzkMtkmmAOe4g4zVQ+x/R17rkWmsffNAdWTefoC+DyVlCuZEtdVi
bq0yiy+5YwlMQ8T3ytN86QqVwl2I4t+nbGsrZ8IdAl0qeNfK7tdHlqJ0KpGe
abZzmqKO3nTDsrSpuE/SlcpX4whNqwsLvUfaIODJQL7z/pwPrsfWrljAwkAr
c704eMs75bs57daPGcs/nUO9BJ2mOCHMa+jsQY0oPY4zdqnOndeEmdjwDcDR
wYTY9uB06J8+3VHMFEDvg7xTU+WSkEzs8p0B79wgpuWgAc3cvCcChPh5Cwfk
BjANTr0KeUplX0XWSETOg9C4zU4jw8jGGLBmADIUNn8O7INhyBOJYKBQ0ZaW
AhNEue7K4Wcki3lrckCvZXgRK+MZr27WbW7jcd3hYshDbXTLXYuANARvv1f4
i9BPyVL93JIHChyOc0TWuxypmiNyT3IfVtyByTkuuqLirfoBuamdN0TOTps8
/nBT3SZHkQmuh+RSG37co1bW/JhEFFYh3Il7jHvf7lMWGVebR7D0x2MdG+lT
L0fpXYPF2nI6/GLAsUteFNsix2/ZJgV+dR8f+VOGIlFv2odLXVp20giOmZXJ
ExCQqpwHS2YPMY28ObX5u9vn4Ua2H5qxkGkbXjxqVbNbT+SLpB5IKYBDkcnM
xU4c8bGHrrieJEiMSYOtcfz3/3A2qPz2BElZjTjkE8yQTztu/A8tQhktm2R4
spu6h9+HjM9IijMwZUpXUQnaulChI2sJKv3ql5/FJTiq3r+pG3txidEzoiuB
fRvG9DPi/SR1eyBf4W+GCy+xYMfu0279K4Jh5NTovuwu0/FPbgpACog8Ay2F
bgFymV95yQAuc5J+g/Yrt3nAPqAzKyAyM2830l+pV3NvRkAlPGK4AVbmsy3B
WShEgZ1oyaElPyvyK6oKhoFTc0gshx7YvKSETe9cYpMsnG3aXZOgqnZ9wny3
SyDKXulQAqfmlOuipn+47xF/UeQpTVZNcJGzJ2SHp/Q8FwgjZv/2GlrqkjND
1bgS3O4QryrzX1EZ5tTrTD+JLPAVl0fG7WpthEb9b6UIW8ygPw8IUa0Iv5kI
BRHg/6oNXpX4o2yySsI3AOl2/7QqyTfsRRQJp4BUPPHDGn+p9+yd9CE1P9Hd
G2ytu0R+junw9XbMywI3/VsA2B5XqCERYwO2We+7Co5gJ+uvS1myFuDlA6tq
6RPjvWxtsqKql94Cp5eNnW8AGletfrAlgkN54Slnqhi9J+l5PdMI266cvBmj
zGyAWTZ/ZtT8d7XXaSaXzlEQwKZFcKB9z09zqD8rsk9ANSJmGdm5TfXLat88
kcYMzqMRO2pZdVna0YxRUS6bak0p7bIUGvX0vWtOWkxhQphk9byUVKG6i1z2
0vH2YrNmn/3pNFwOIElUeeSOZN84snybD1bDgijPh0/IiPFPjTlANZ8HPi9p
juRudQMGDZpYQHsUhgFcaf4NUgdML7ow+BAmy65d/+5Q82aCwB7roqXzi1P4
fWYPJiKeRmRKU+l6/2OcTkv7tPJyM0LW7Cv8/605Cibu8lXsj68QcB4hmPrG
S/gwbSZjXGWpXOz9Y2fY6rDnCCeHAMWlZG+bcrg03DuAvNR9kCMovvJ9WqO+
Pa4W+hLiEcXoaJKQxn2a3q5o2b3B6JKmtNbPapOCrvMZakR1/8SbmwbvyfID
rMZvnOa52/RLsIXZu5o/iG5oMCQoWAPueohYDsBjXoPqKAkQMeENCZWNJpoS
BC/3wF+cfbzhU6XccyWhAjIZADzeg46kwH2IZEern7MHMQQvvl00iNsYC7uC
/gpjYKIupOpFvE3EV5Qxxaa/Upupy4lNWMSGfgx6yKzm38LsiqHkH5pPChvt
jN3h2LRdSN6TUl7DCRJsKurJbdfiWaGA/hmzdhQadZ+M8yfUGytgTx75jVWU
3B+NPWtXuXRQhySr/bbG6cph+qu2hcMsGakJdVeq454n5rDNbJQYqLW48FOK
tDmzvGTWoGlohP6mWuBKVVmUQMCrEQNtqre2dtv6I8C2QASF6IkhIfq4Dl/O
KQVW7hvFXdDmE5pCqTTaXyfJ82eSppIHpWIuHVNTZyyMKBSgxO//WKdYVpo8
lDHsWjWcb7m3DC00hCih6b4vzBBCWOBS34FUQ67WC7apCEzM+C21vf8IUTN9
MIRuvxMbjD8g6qXRz5hGWfwS05VPqRkEPOh6OgW5Lu7OJv+apFm09P/3MQeV
7a1XiJ9T1xDbQV/GC2L+XfgGjgqsdqUIv9TrLZDTnP8Zt6cS4n9W6evckt9O
X5GrEE0h0fBUVEjftmvwc6I/cUJB1JKTCC6EGRM0WRMlRWBRSndsioRS4oTd
U0rwM8T9Mk0j7Fwj7gySSEqCm1/Rrara5SAJCyoX+IKUbl953t6W6XWZm3jk
opBUB2h2U9K/cX1LKh1BuUOP0LGPUWuniLDxza2DzWRS/wyU0qDjwdhBMYF4
44z9/N6eMbL85ae9FRuFjBnAOL6mv2jweyUmbQHduoUjvHHnj8x+3H5SwZ85
iYu/aIjB6JBPPFgiWwAOgNg4/NPQ2qH6R8k7GEhPB9+mrMhK5SYCeXmiB97N
7+wJPOPLP3sr9CbIklVDHNtwrqUhtawvDiAQAWuHNHsBIqkYk3pFYxg2yREb
IF4TFoChanwWc/Gdl0ZgaRglxpo6Kt5Bzx2ovefpMyJF1gEPB8viQwzTllrR
079yDoXE4/SGW5hkTRBngCX778FLPSirEuem/5ffPsxjy3ZPsEBmNtqqnU9y
F1zq5jh1TKA1PoTOvtM2I/P3B8ihJzvLwBp8qyd8lQkmfNLJt+OUTKVS1ZX4
TBkrU0lLzokZM4pDeOoaru6zfJgSBRPhMiMgZHY1c2/FYixUydXlmWsclIee
A3eG2L3xEhY/41bWvAvywhY0OYW7bv9ZH1TyF6qXS/gwl6YfqLEMK4r0+Enl
nm6cTkXpMxViDO/jfee6TAasrAWJh7/38cwiEfmJ2qKt1D61TcSPRvhhgncQ
dSngpGUQ6wLlImcb5cJUDAhJtqNFBQBhnEdTTP5DSenI4kT8dBZZ3YeuMcNJ
BWriE2jDu9XJ7/HEZcw27m1azSb5l1oePqAKnaxF23HCOJoKBKd61v9Apl/0
zpHXMmXQOsBx2iVNLCGTrOjWr4rF4+QXfdRv03vU0G747H2h2o3Eio5CMURZ
ho//+tVp5nA66JMyBgYN4DaGSA6Rud9kzAxhNkJBTbm+GHVldAVbea0OBppz
mDs5q8DW/MfPGY8Kt9tqktkGe5R8nZOQuw3iNxmwypKvLjtMCMpbnMaXrhgk
JaC61bGnFYlk4mVWaQUm0mDBmKL5QXmYI4NJmZZkpfuN03YgLljf/Nk9bHav
4XFcbNzAoKSelA0SKiHzoGMT1J0EeOqagrwC/L3Ab+lEGX+3JY/jA1DaGQib
PkSJIq7R7z/vjWcPuR9Nmw/BAMc/H0qs09dY64tOtrVYtcZwkjsrI9rl8h1O
v2bhiYJO+44AvU0rksw8IGMiVmTbIq+xtYGGEh4T901OaGawjTfKRDc2cWQ4
B6zn8/4WpNGe0TVZ6VgP7SM9szyF9/pZVyXvwyu/zghvRcrxLP02DaN5KcMj
8Rhn9yg/6oAOEvI5fvypTzuDtLf3G1uiY4TXMiMGRW/xCNne/HggumdGG0MY
0mk5RwNq+O6y4A5XXiY0KoDvW+B7OQ4Z/Et3Z2bnxlCErphYNbC4buty83qB
68Z6GeVz3ny72R3+w4nCJ6HBQkCwtT+lJFsYZU8dsbOi8kcfy218SGRT2TQk
Ka0ApFv8SY7oFHgbCYSvKB3oMasLqycqwAWf8YFt18Arb2ArqTA1fq+aVI3c
nRVHBNYVMTnoVQuTAEj1eWPrG+owuIXI7OfFNuq12RBWO8wLs2XoyeY0JIkF
54g/ufE35lLfhiu491Y+UKQIpjo1j/NITjQZBTDHcp54gSIoqOevjWaFqm27
3mEtqV0xPRziuHy2M8ApFF2bNn/uMmnI0v4Ai8QSqpMCqbaqLRJv3FeqYRrW
1NPFowEPXbrRxrJ/lVvVJFeJHw7MXhwhYoK8rVvZwu2swf3WkuIDD4umvZhz
6/hmEnByL3z6J0o+kc5Vm/mLeltNky0oqKb8Dl0cz7Qsde5hl/NmZ+TtwQMM
x18FaQloXgKe90TiiAMyXzQazPyaFHZg6jMxYeakRknfRSX/VztUrHCCgJQN
viL8cu99pLEpfxJhi03SliGa1b+vqrpU/FcDhiP5/pKTG29fFyZl8a56uius
UMIsDex0Qtitvuh5P8DwXo95hazQnFto745Znvw1nc8yyNv6KBCLkTY4M6Tv
0FA8tw0Xz2DWa3qMK4X2WgowkKUPR7L/CMG0j9K32HCLOGweSWim6Dc4i3S5
5KuTDClKBs3E2MrimJ3cUAUgO9yMoOByu5XPhajduOr28TPoumyCuq/TSzLp
0ZZCmNCkG9RogXvKZbQrEZnjhAHCE313hBY6418UHwDgkSqGTeot6Mkto1VL
YosSvsumtQ5zc8XJdsiRowuAHuq8coAkVZJ1vRKc65aILHFXantXoANOlCL2
zkzT9UtzeG+nCXCihU1A04iKtNig2I3RzjK/OtSqinlihRemKRs2QHXLprfx
WQ3DuhtC9o8F9NYT1BAjPe8p5ObzDuGbmLHWL2g83QIf0xKIvaP8kqdE2fX4
2R8eEdvQEKheHIUjT9lr+QIgBhveADxJzGMSX5lSiBcL/hHKLQpVW4PxcqxJ
l8Uo5xcO0+VKvYMMh1ETY7BBBPglRviz4FNPCxfxkkrSn4mPnaddhjKo9EYs
/Jr5yyT05wIsO0SGBn7YcM7Y3M/EHCscc5y5U8IiabEmfXkTrolI5QeXoOaY
Aq7/VgMWI1W2ptBivQRYp2eKL0jpQD7y5OUR+ZjNKCkw/PrOiQAJUglTwQdS
V6htogJklHKhmY4cTOCSIhfzcFW+/wkiDa3eNBULPCfpwzReWIu44uHUZBo6
rNcmWNzqFax/NKptalJg/NSnDA1wqsWmSiMw84+ozfJeqVG3bO1YS/GbDlid
7BpykleX0ceOiXgf8lY9kWkoNCfh5juHyR2HbOuuXrQhhpWzPs7vzJ2fAbVe
2HYf8fotCYl6B9YLJYJ5sRG444Cwj2aZky42+7n5G6WyiMsay4g1R+cpRSLF
BtyuhbAmEKu0e/sKNOdjaUzlzQs82KW+krpPPbb0iBJqzCOE6CG4qwDt7T2Z
51GvK2DUQ5mg6okLHmuonh9riG+ukqAP6s0kMiAd/EIQs8vj7JivzL8H28sS
177MrX2SdwKrOahYmo0IIvUY8k+02xTUbMRzqpGLewA5MpRYAdHqnoRUydH7
O3Uc1ehZANqq2/Hw1EgX8lTBkxEHyW/MyAsbUJAFVilDHiJE6dOyHnoI8ote
a3xlhBLrZORp6G++imSPUtlw1owNF3IASXD2uAyV5hT8yBX2o6phUa1Ku0A+
1XsHpGUWgQSd5oxZQPjRd6ZGfVczP2AooWmMq0Wv52X9cbbOEXPzfNyxAZED
cjy4cGkqgPwX982Dx+2djuuIQyq21HzBJwdC+kaj2KmKAIH4YX+5YsuCLzSg
Xx2lNbw5AeDYEYoRduxybBTIEOz7FuObH+WnayiDYFDFRPZvg2Gw3gmrO5gC
ZEU0BaHoPl0rWNiI90UGWJ5sxFrDGpbfqgLcCtNeWbiJkji4CPti+WftkU7c
OdnFVcwSxjCKID6s58w3Wi59K0TGst0l9wIhmuB+j/Zn3MRdsABQwI9ef/TG
DdrZTQe8ojXtmCyK/rBwlZZIZWhNFezilpEHdx3Yp4becIpdgWb3w9R0gFGT
/XVS2BBhBkvrf5WbvXjtKwr7s6Vj6J3jl4oKDpN3fKQFh1YvfRhlxlVwrYoa
l7hDT5kKGAd/NYelb802I6UJDUTy0RxiUFyvJofLRCAhHcoibi4hDRrZgakr
N47mLueS5luI9Gss+WQUQ+m/5DKsCxxbO0NkfrFTyj4h+okzUJSf+iJiPwuT
/MDIkcPMx6fFMu+83T/21xlaiRBnZ33ajCoqfWEQLAP+eUKxw5rTgz2vZ6i4
5kDN5DVAqcUBLo9qNwoIibTo5B02DWTLH+FvUkDrPLlPXxOcc8JQL6IP7Jte
ab5CQ2NpZJxBezu9jzQ8RxQSpQOXHttccEx078ypXbnr4SkHVdFVbzKcYPjE
s799X7/Ft6Q5bFD066NaOZROIWrBSiJcFyvA3k61Lf2GZ2DTixw+ISAze6zj
VFkDucCeQWWpzcFNE0AnnQMZYRjJtzYNDILXCWC9cL/k2g2IZj77o8aRXxtG
2j1Dv5XbgwpTmmsDF5Fk0ERGXpRvi63AmcwneDWXtPVtAuFi2QKi9ep8+NKT
Now/2nY5aQXwiFTukXegvwjDgGxCcY4zB69k9TNaSMeocHBLj3v5pi33kHGI
fdXh8XpRW5mxv/Fwefm8D1xwRhISfa/tXZVGYS1nvdum0lZGYLaXMXYFQYR/
RT0e/4kv3TPGQ/nFT7G0PQCaNill5+iojpApMvh/mpFKzwPHMEVeKbqy7ih4
2kv+zEadP/C1lCKwwGRwPxsG/xw7sSL/IMv0lNLj6KDKAW/3V2BQHIC6CAdo
BO282Tf99pqH4DGJt6zUUtzYMm3rHUNzvkjbP3CVCJFzFcl9FxcsLifqc10f
exyozmfd7ObB1lmygQ69gl76HZED6rdCR63jYHvw+hmNWM7ouijCS5GIob+T
uQWIR9YA0nVVY3ponQ8ZVxYjEclju9vDLN1xI1YxzjJHtis562SMmvcDwwCC
KQcehEYaQTTiTdMWcoG9uXct6g69CDzBF7JaiBL0Sij6ZHbh2+IEggWz58Te
2TiyazdplR+AHt5rnOhXNvykpYpEWI4nieibm/cArCh0440G3dbus81hGvUR
/G7PK4sP7U0AZcHM23ExK9QXADyoQJ+stbuKPsI65V9pkoeQbEb/iqnhMN1p
LbFajYD+af1v7O2X+Zk+y96cMNivS1dLU88QZBCOLbOfLznBSupMkdY33+8d
Tm6PybyrymnfpTj4pkS6X7QjNaZB0mQ8j8Mf/5eimMInt9s7oBnBS4HrkCbz
fk/CBSA9pPr0R7Qvm6bhNkGMOZRy3gGYS43FlwTRCeBCk1ow1D/YIsNLX+OJ
7+IUQdYmsN3UzSTuLU5PfajShu8N66NQ/a/M/VO3FLl7DB3+EDTJSqxn/gM+
kj77xI2VOASNEkqIeuwERRWzxWg6JeG+4pRsXyCxzOE6Wo5NRXcywSqJxHJi
WGgH7hSBDuVIHVAKOicA2LxIahulCCDN+dt0dvzDqqH9N7Oq1ly1QTjtfv+p
DV7qupfgnndUo/TpXP6pk9Y+BZWJIfL4Q+uPSAc9P6EMuqCtLxc2yVM1OyxA
0y2PeJeXPdmNnBdmSfOxBPXDLopQIHs+mHYgjsqBPKD9znymVZtkpRND4P5e
S3+B8Wex86fxiMSUOV0FrIZjvxn7YTpBYEVpX31ijSxLJPw4O1pUvTsiOBuY
yBklzZjBhPAvxeCFykfyC0yfGbM37TuJK7vOBIntqwv/eBH6DeZ7KWByIJHi
g/eRjzPygBn746vhEXhuXdPgHYn/y8O3wLW9maO9HNKB5wtqGejaxFhv8qUS
PMoOs4hM34B0196UTTdNEoF7qctEWHp3oX7zvso5M+6rMIr40xWRrCM7LDyZ
QnBboY90Oi49hJC9pPtdZCFENb9SA8xyd8P+IMlrtoBHQzV/Vuod9jjP9axT
Jt67v7jpKRUQqkNZ+AxF7hDmBDnRxNQoUzhP3medUeDglTRoL3y9aUUfktkq
eEaYT1pHHf9NExAtdW0a/dPXoxDrS1ZeIqGzL7Gf2Z4OqTeEJ8pjHybntfru
XSHtY1t3C018AHY3Ir8bjOx/cYK51LYhq2KvtIJ3yCwJunuwX+b0d1Ka7Oyl
VF6N+a26Pr0NQqOYBtBNYUFZkP5m2pz6H3Uvi04DfX1iop1khfUB2gbz+2fX
PbhVDPEsB/ScDgbm4kY+/SJI9BYiUei+QxXipeC1Vy89++3uSjmZQBtsucUr
wgAkEdxqNphay6QwFxscEo04YLZ/RYpiK9FtidRYhoxyqpPneom3l4Y+LgLo
HwMW0xk+k/DbFjOFKXvleCC9QoIXm3mFlr66nSsA9GtLoMwGVQXXVdwXWYEO
s04ZiKhhKyJGnggSRQZMH6504gmRPbQMhVX+Fjpj6oQBzEb2keSWJ8maWID1
2uBaFjqJIxfONIWMTyeJf7PYh1hJfKwPfuu1kXFaaNb7Ed21hkWOSyskA2Yy
dKwQy/2L55G601e7fBhS1m91U9AUm6YfFcbb+yAhWMEV1y5wTLf1yobAm5UT
OfzLCgktvh6qZ15pDr/osZt+0F3VwTBwrFLNF4x7uTATzTdVdiwxLaHVtOQm
8Gq6gFh2OgBeDiYpXDoMw7tGtwV1kC8WoXb1vgMH8cNOk/uII/kyhTTELBNK
pR0lRaaNLJxRIlqTEndFyIY/HIWUqy6W5oxdFC5NereXbjN3hXBUX8FndJr1
qTcWm1n7uOhWILSFKvWCn95Y0V4algDaS/wPMSvWjmiXpJHZApjOBfIJDp66
tP9TAuIdWzyaXo/GWFK/s/Pem17lCQVZ3CHtEtXGw3ja4jwI+Im2e+AN6t8B
tnzzJEaHWJ5Ql9Tw2ZIMEJJKrQIOH5SBYJmUDyZW4n57Lx9qXi4c56l0m/9J
i8wTMWd3LjSGfXaoxaCP82cccGw3nM9IgJIxRXaYUYPliSpN4CNoF6LgVD6t
/kwXGTdbl3RxaLt9oR9yfSaOzBVHGT5rndotxu4ju9J/BsNJVOT1goZNTsYv
iEYKoPUIx1MkutDWy+EX+3tEh8E1EXQCJz4DQezPxGnGwCNk4heWT7eFuqcT
ciaAUs8z8/mgg+nBVTwxLwM8gT+A+NZZjnhxaIbgDklCC3ARaIKlo/8sOhau
6Hxb91ymX4mTHN+E63GyPmTe/6u28Nt2icyNDiWWCIdH8m3jzRdhM9Ulbh5h
zNs9P4DqL90Mt2X6CFk1MRWBhzHlC9iM/dFj89o4wDW+HYRJ0RWfVNw2GHWf
q3Lsfan49j3S6iQ89C/037l7QuLb9gclrKD7f5MaNjER8ZenjAGiNEoWHtmf
8W0vlZgmtxNBwXciINwzHo8UyKZG4qUdLRatB5HXzrU6uF/p98KBcOTllHpi
WOXXE3wwGymqcqcsSrKOmXhaGa+M/0itXoi7wTHLdpGJiM2ocUIA4stbCuWN
y2AvsbfwjMlf5vw2rcK+ayhMw1cBdg4JoHEOTduxTYslTFeuTNE+8rWK/36k
/R8869Tw36Pgcto0mdb0hwJrgVagTeDPewg1pYk82PmYkJqqoK9RdG+6Vw3J
tt0yp8XgADe/Bqa6dMLA9C6ePFqkEyIxpr4R3TaDohHThgSK9OoUu7dIUHr1
uNI2ClTcl9fyv4ZscAUVSQYfKfNQYSnr9pot7d7vlzDk9xV7wgTYb2GQjdlg
/N4dqgPp8IzHMV4xnr6Q645nHRyuo+hqI2RMuLLEyHMd+w/Xsf5Sn/BnQ6dw
CUKu1+ruOpJEC7AUnjqEauydrJDqaEAMecDNnqYjsj09P3B1ipK2MgpNQ+ZG
xjZpJyfZXUBkQC0D0xMCNMmeTLRSTdwU0IqoUQ0109izbdWx3cT/6XbmM8pf
y0pOBrp53MIyW7Aj5quzeay1vtWYW5KLr+HIC9cApEVu5QKCOIYe8ANUCq88
aKwq2cCraKuJIar7vaX9DSicORBE6mpBlJaU0uu5PFYryAaYdgag7cn1a+6I
KxFWh7nWT6VA4kmoXWuXn5qj4YOvdlMAJBFebsnKvHeaReyUrFOOMnzLANgu
xa+Z3cv7BQZIlPbYzX/8K4TIB4XgExf6SVl5TvNSXzeXMaeP5DpUp5enXG/3
rt0+zRpSxO0qyjygAwUYT+Xa+TlDBD88iAZvEWjEpmK4NrkGwHnulWcfIxzt
1tOkJvuFYmyeZ55QFzfbSRfOnMJokx0iXnb5Gm2HfArLH+l+YXimeTs+h0Wx
Bor6mSaflSMg4ojaizz8FcuvzcVDIdkU2l7+oOxLWTI5pADZeBQseX5/mQhc
GC6PyVpW5LIkRlJaHNIlKaS9Zs4o1rc0vNDiLj72EpoNOKKfXoQVZe2vmhxg
8asoaIy3yy5YW/1nFgg5Se4ahnRcuNsmiBuNE6OxL2kIEfOOLUSXEiz5ZhB2
FD5bG88BJHGT6SiEQPikHhSstbZ80Xc/Pt9Tl1XU3BWbUzVvNz2mzFiXgK+o
/yiZcTJRhinv4CT2Py2CrG6c/v0REzJxy9GI896714fLBJpg7MsBEhVeZ375
ZaB/pPvBuu7kTf9mWG2bsihr36Do6VB8fMby+0ZaicMQz0EpJTMhOl+v6Zox
pQ8cml5g6igVo78B7J7++u5EWfWvxeWG8q29jW6Ao0C+HEjN6GMNetvUFNMH
J3n8sL6nHLIyQuqWDGLcRTtU9M+/Jro9R3yUN3N3FcLTtEGlysLXx3Qie5v/
OkgwWk8yhcjQqHaAxrN+ge0Iz0xZiZWIwpANpMIdwwxPuwNao4kl4Mgq3WpI
IsfC+l1zmAz2wqPJN5mnhPuw1Q58ePMT9HzlJS1N9aR1xe7dqjrU/ERpkWGy
OFnHpRbmu6hnTL564pfg8beXRkHXFeRX0sgMNad5tCdLGdQgSCxzDpJN0osQ
PcceS+tSbVkB+YYaMD6kEdBmSjKxI/Ap2LzUgdwbZfSLXCzsmziPe0yfq/2i
mTqrJpt4HTDTGC9HaYApLfhz7T7UKrEnpC1EkWnwj/rlpRfY0PV3bZZcU5dW
D2aT+kLt48mXK1Qfs4XS0YkBzuR05l6UEC3Ii65Wn5/BGe4mhF7csKQKvczh
pNO9K1hDUSV8RI60fxDj8Po+W+9i4XXc3MT+dwmBcMkDKgsgfYMkZKDUVYSr
iGU7DDNdDcflwjwFxDulxQc/PgLPlEIuhXCVch/UkSzWfmgdT/w0F124Lcgu
QmTTncjl/qcOBAayhZuEcZo8pTk8DXAoXlhlZNN+iT4JsYCHzmZxNTmUs3UL
imw92dOXCgrpJYRZCq4VkBRTupzMOvA3RSHAeUAR8Phc+MPj+f+8XqbkbJyy
k5y8QVfh+PoLql0gZtqS1/rKmT+/82mudHIZichGAxaXVUnTxSEovs2lnB71
CElL2gyYjPSDL99UZ7W5KGMoh8nQmBQZ9oEZk80dGzVVGAUglXIgJsAYuzBU
nnNVBHccSJhaLUzyeUF6FW74EJ8BJPcmUu6J1tbdb1AmYn0gbFAj2MKX1lBt
/TIUsFK9L+jM/FE5p3qov+JYwAap4xTGynml5KSsVSscbmcgPblSQuhX9tMS
ORaaSgR4A2Kkeh1cI122zEP/nbTzpcuSaN4h7RDjjxnapf42gPQjwHi5R+C6
lPa4l8iCHCaPUK2Hv7N7Pj7rfnzlJ8ZDpzI+r51p+uAkkhEqIWe+yX3m/461
6WKuher9xXzZAYfdvtj7xdhVUPr3XWgW8E53MgWd++ftTZV1EHrYPiOF3Ure
ZwDyclRKoNoNgKxuplTYVRC/bn6pObqI3u76DZ0J72U1vZAyeWRixLoOZ8Mf
4STmqVrVfcprj2uuBX37lpZL6Q0BX4Y9DSyEwe+LRJICMbMfn9nrWkFqm4LY
fQyva7mf4b84c3fqDsPlbfc/loysjtuOrDppERwk6fBSOmxZJz/qLqPJJ+Dq
jZWhl/+jvh4xu1Jz1J0nb5ieF/4b0AXnUsm6KlGiTTqC/+gmIbHI+MW0P7e/
yQiwt5CwSxPRmMe60fSi6wOsW4YSoEXSZ3ZQ5uLIgRb+jRGbvKaTm5396TNa
rotnKQH2zQXbjZJga2JDNff++wnLc/7JsF8Fs9f85WTMMTF92tyUlLNgs2kK
94Fp3qU68U/AXB9k0ctyHyMbb7ZjU4ta2boQ64Teh6bSf2ES6evsAnTb3UPc
npV9mMOk046JOVuMP6zC6xN8jh1v0Gq5De0YN0WL69brJWPx1N6Wy469RmsA
4TMgoND6EolOn4yK0Z0GgMY1s1dnzMXhn7HRGXWtHyCv9WEYzw4fSGlWXupf
/5bMUUb32x2t6f7IoT1WP+YF3lx8t1RAj47V89wvwnpzVuuJjaL2NnmU7D+j
gKDNs3y+mFejTLrtf6pMgzfWSAbio3zRk0+2/npLA82rvBAla5FaqXMfz/E1
pE7DUI7JHZ5C0uBhMwNMvJFNSZ62Y34qRCjP2QNUIhkqhdT/4kM02mIvKlhS
VDk5CslNaJUXtlZHgwkzfzYL8T7QFXyGWRv5159XLpLFsHELinwPO0NAYun6
JFdH3tjPJ7FfH5KsebL6X3Dsx1oRJjR6zqYOOJV0MhHqYh1lSbn4yylc19fY
ufCvlHZvhKXOgB6Huus9Y2Vw1b90aTDAuKT0QHiY0LEQbTHBRBjoK8kGLrPK
H/E9B5DmFplsx0RH8W2+2RRcONPtcbi1DJAqpZp7aE+YEavg8U2nTzC9LLDH
ol2nJrVq31WuUS4RJiW2ySe6U9pzY/SgsTBok3awsIlYfKZ3ZcynxxHKpDkz
Dl9lpThPfiHWQM+foaPYc8ELueJJ5z7Sp20E1TKaBKNHivmkiHWeKeMHD9lk
PEIhb03OXeREqeF1nHzqCKoa+lBdeNa7sa/rlVKeM8qVnN176SUzvPQu8DoC
bAFiIeWzW3AGItkkeb/FRVAUgCQrwZkvJTZVajMjUuM08eFydXtQvcFPk94i
0+4hfmet7Y0QEV8sAC+FAJ/l5CfrqOSP7fXO8gqz6GbfeEWBzRYDIdtFLBEA
TmSfUS87/a4fh5ZCH3Jn/RBx4/c78v8YEFL3VVdKeupxuKfyNmntK8TlpHtE
GTcKSa2no3PrO7rm7SgeOouCKUVZQQqqHQn5nAH2ztCiELND1A1JXUhZIipu
j8OjY8j3MKSuDa/jGGLtL1hkcOZhrNei8pxEDqpzYK15y2JzPx1zMJEmGA6+
z1Jz1ZS/ZqNhQy38kwJ1mUMESuU0N+cl2W3jcHExUlkR8xbIVfmRqTkLJvLN
IUSV3lSY64oUA0bAdoT0BkKTLZlbiqAfXHty2pK46pzjbOcASGJ8ZZefndgB
8REmP75S6kLDqn6C33A3l4BSD7sJDT6sosaE8zmb8IZU8UMACjPDZm2XQoGs
cFZ6Mk8xEMZQ5WpYSGmvazJHU2Lzdbcf4Cbpe7mM5D68AKsgI162rsd7RbbB
WhFNBeyj9GTF8sEkm8oQpPZnXWtiVmsnA03XsogVcv+31qxUx13Nts6KG+K4
Kxzj2yzG0DbTPochf8Ql3TS+lA1CtpQM1xBVfz1KIl5exa6eXsTQsKpJ3xR1
iL8rI+MRrUk/JLqI2mtlAltBYBGNG79tExw9VrXaDyaU/9LCPS3zG8ARDvnC
JfrGqHEQEqWkDTRxa6H7F/daXq/z2Yrn6n8GPdhod3fbihtW4JqU+MV64nYS
7bVB8P03tGUqSUNAUkR2SstB2FwezvrWhN1ZQXShDceEaikw6nQ7V+sFKh+a
zf4es1uDhucEGBn3vUqktp2jdYRxJPSJ3dzE0Yn1b0VMUh/vLyZ4nHljItgk
rzLFMWFyJPIJhUHzTgmUNgZDn0eI8fpkvbv78O7m9vGLEkWKixo0u2zlgAaL
29vlD44owil0+3tskt5kWfGnB5Se0MvZX3leHZ56Rp0i/0ZJ48MZtgQxHD+J
PJwajoIj/0VV6vhTrFI2klaIM5P2cfWZ18dwLkU52PNk+QRtSajadIyZEW2c
JwGAFUPgafljcKQ/kKLe8eR9kTm6KzC9uWJUnjMEjxDruWZ81XNmrPZ0x0Lz
G55D9+XLxepy3b2OXUKMWwCr634nKgPoeejPAmbgyz/kQUUK/V1HoHvJR31p
qn2s16c1dcG/4zFzGoZEl0CDC3nZbPxHjRsjyivHS8TD3UhUPBVBgJoUm5d6
H50F8QvGiQsYKO7jnGgt9V4IB4dOdXlbqNmf1e0ZsJs8B7clAvetbJeK3oQ/
uRzyaP1yEFtUG4WcyO6dL3vSGNzMU6gc6cwmsxZ7baOEBZxNokhTFwaaqhX9
Usyt0E1w+inEL+Jp5rSSoFbnvqQKJmKPxPAl160r2yAuK7GoW70kaAKAZA4C
kuo9wIXDrVMz0wOZ+yDGxLi7/6s0S3Vr9RkRFhLj8Ajm3Oyx/G9ZCIsSuB+4
liQEuMfOSXRteSnxGh3dn2Gq6B1zowR1aGjSDWcAggPWl2+OZliTrOg2h/4h
YoJsML1vy/Xkd+wFrrAXNY9k1V3ok6RWo/0bQRZy+2gTGpGOYJZ9IbSPECjE
Slhp90McFlRTsgcR47NPK1jUF8ZmH8paCZKMCWJJxKYBN4Knw1x3wbZx9Kf5
KPFMM3NZFstd56qCMJMl5Jdjbazdo1RyHLEEdCnvBs5io8ybc4gIvu3+p06C
zzKg/A7qQW2LtnFMrIR1SbtF2DGkFGrgGE8xKQrYw8HHel+EMcZwf9mdGAkm
F7ZVJTD2HjLKUamE7rr+8NhAMAoy8HML0FvPGROVbHD7kz1NHNIfRMmw9xDQ
6WThMNsJvf12TpW0hLKi+xhaXDLzi+1+lgOUMT2sOHPCUXgbR5Phiw9Gk2JA
MLXKp7VmxJwEtNp5LpFewF5Vwygj9qK53So3dd0HEJS3IkQWTcnuTJzGgbYc
tuFBvk4zp8pzkaoMrBKGZT/yZ+mpWB9v+tMBt3eZvJWwGwsd1iviy20xmxtH
7zJiKzdHgHif6aRDyB2Xk2AcFsahS+JKQg7kHNZ3byA+eaXcK4JBgD5+VPIm
RdZDzorNvGJy7KmVwlmmhtqGUM2JGu9UocVuZCLgc+8wwBKvQYUKg9wZSdVE
F4J8OPxi4hlsy2lJ5RauNEumTTJuXOi6U76Nomz6kgu6NULGcBvdJSm94OIT
I4BLL2UASWECkUGc4vF6CHZPpYjeS8coQt3HtvAE/z3naClgBRsnlHhOeHGf
NYpTkyLbdSBQhlNdhzot0I+Gr5ytzmtcW+cecz9eHFrx91a+rhO/r5vv3Gfr
1SDwiXxp/y99g7cjmgI2o8cXjdTqxNhdrhHmEPG18yEv0L+Y9oVCH5ctjJMp
2hc++3v2P8eYEV26kqFTfqUEbiAZgUeCMcsEGtmrwoj3lZ3dTkwwSK/ed9bZ
t8NqVSndVbZoMtUrGpBcnPnI95orMwmH5XiBOJcjtVzeF/L/1OsGQe8bofTW
Ru4gBe+FiHWjsyirnxsYU6h2XN5Ej7cgN3b1A2YbRT96qw54eRUQ/K/LofE2
ZecmFSaCTwHtC94/qKagSXv0TfY9Ac6q2BlZoeNo5rzpREq2tUgHEratAT/a
Y920qgb7Hwfv0xSTlaL6XeX6qJndEpIwcY/xz3eLJj3BsFieE/bO7r3zjVj5
T6duHqbKes4ymPIFD4z/mOMVRF9pEOoPJiIdUBm/NBEOvW/9owdZpBGlb/cZ
S128Fsq8VzV7/1ANW4M4IIxRBRCSMK6DdWyGrNytupu0TWDOd7vlWfFuY/rm
3Da1boXNvRd+5TzHSEG50dJ2SfTO5vViwzfGb1PB1WAeriIhVm59A++WqFuE
XLJuNuiPZ1H+34NJ5LKGYghKgkknSU8RMc1MUzYW8UEWw+2PbNyIT1MYm9GZ
pIuryOHvYjnvS2dXYE74601v1DQCOmJVLAyqCt502xJHY5GWSZ1BQJE5qXop
CC9hOgZeGPUVSIs8WOrgG4i4j/YJTgH+8xwpp5s4LeykyuNKdBbe/fSDORII
iJBK36EOYZr8VpLrMX4jFKGi62gBq22ndJync+cgqzQvWfCY8Pg6MEXxeNwR
ZhVyeDiH62av6yJ0/zRwj1Thlx/nigoaYQ+hot7xUld/eBcwhgCRQAETuAK/
XyeUnNtBnumP9ODm21wnCsMnPgF+fxeuPTpmfPwZQf0Tz4MQKFQSXTD0z0Sn
nuQSR9fivEeEDEhvIsu5Ik9c6ZhMVV77681Y/JL5YWKXPJXfraPi3Qq4xvsM
FDsvEpMCKuOuFjN8e0OoRh0TPOKjFMqHHTpR/j0stlxILx6cjKTrY487BJql
DQoUmvZEWAc3NTH6UZJK60W6te1/Iq2qg8+44INb/4wkXeDGyRs0imam0SAt
NjlIkxzcBVvTyoosUox1mDgDYOz1EcqFqUWEtIF3dJ5IIOLEUBpjLlVaw+Nu
D2Iy6XUWjfq1RwPY+0BKMXgiTrEZqKdf4FMtEQJpbWTTXrFQXQV/JRRDZwXX
2qgb6JpTcThpSkvZ0am2T7S8OESnXLky8F1sSjxINWxZPvzJNWSLHu1v0LVg
d4XD4x/AQMClzlPELkLDB2g0me40BD8BJ8mRwzzWRnDWNv8mJcYh4mNRYFFZ
2zldZ6EEpULpm3QAP58xFvIpsYv5QiqziMOCMDEnETTadoaXRFmQl+D5lEZX
ZYViM2sqYVbXA0/gdNKl6xkqngexpPRlgs2YKQObWk3saRGEOAOlLGxqHrGm
1ABOzOh1zKV7j32LOwyox0Gy8C93686Lt/kPx9ET9GjWYStAy5jak2tn3EHP
J0+5WkV/W3nQOjJxkM7DlTJQOvk+sa6BfiYWLLp+tc5esSr59NacsKNcFj8d
ABycVr0NnEd/eyRl14Ac9RwHhx8kxLfE5ZrplHNjiwmixeyP2G1uitDKGY2C
DipzNpbz71NuSfCDQCzYEXMIjV++wjSdRUkxsLEcerZ2FYqLEFEGHYfijZts
+Pl2Xx74EzykXxiZEwqw099PKlTnMDjGfgfngME24y/lIJo8/0FlhYwmyn99
En23KcoWhhFJlOLUk/64iZ9ChDj/xEKFK30bxSntnikgUdH37UICMMu2neWF
qQpgQkeKSth65r+sRFyZ3kNwZJoT4SXSeNYLFvv3pVCU8sLc4rvK9AX0YsF3
2GgouBvgZb4LIFc0EmgDH4t5FPGF/l8vHsWiJwUb9gnPB9qTUp83j6Vfb4g+
mBEUIFbplFb6DSsyz9fDci6P8now2hFYQHgkh2nvu/CGkomxQkaqxnf8beoD
Wx44kXxPmeSUrzngvXSFJswo2pvHa+sNnveE6TpfujAT8TgtV0HiYqVBT1/2
nnw13ARCxs0wbqIdNM7BIRy5JUgc0r5JBKrzIBvpKzpiykQxw7XV7W0asvLr
glYTctCphYSmJJx5YIYOarSSJmVdMdDZPcFGP7yOR7MyHFOVdWa61hmKQU1V
N3YTTsR4fLy11X99hVGi/duKj6V4INQcX0i5kSj+THEA1/tqBME0ad49PMtX
WZs8t+Z+H0QhZlYm89H0QYt9XvO4dgy3udDRK+/7nxh79/JVhKfKhJOlvsAY
ovgGzs5bIZVXgWSSuD30XmUjqrbCGjlVtEy5Uhp26nTOxCh/IHGyY36N7o5P
TOQn6QAIuz9mGHmxpA0LjLmm1xQlDsrOKgeZDZ3CzIFJ06tDHPU8KVdkNOQp
pzo9jWGiCH8kh2GovGTQGLQYD+HcyUIr5+otBa5jO2ipD+5yPYXedsPFB1Ht
NoeW9fhCiMx+Q/8SsmQ47VffOmi+q1GAyp3Z/PNhXFq3h5xlXNv+dCzteWFe
BVCxzsEctaaATdMmH9hZJS1mMJA+mAG1ueImDE77YrnxOCUZdmYP6bCZRV89
JSk1U98oiDNjyWfg2m7lJQc6fp9PRsAavo+xWw5zywBLayz6+eZjTL3F5d7/
hFpAm5GUSk1+7Fk30DkspygmUTIdk2k0o6Q79b+fDMCKAo4ynCy/uS4Umix6
Aq3ndJvVcSpJcm7DCDpL8KGQoDtcW1yREFvt205gu+JlDu/LTHzbNa5dluCo
yYX2gh76K33JfDENreEngdxGllKIGvmcCBZBSt6I2s3TkaUcjpnwkK6YTRp2
a3BlxRDJdsYZcHHa0WsjM6GwbdoAlh0oJV5WgUlGkv8cnhByrTMQWiOK1rjT
0yS6L2rKBByVitAIQ+yE7MDn6Xu7pNC5J156nSemeG0ZHZ8a2SHCd3Ucdr5G
sTnNCrpxvtYV3q5wxSnDwjd/mCpQnR71ih/Kr5LlPrMoGZMX6flk/keRCx8I
lcMEhSiodNKF/Br0/mh1eHs5S5k+ADlhuxZcfgr4Ttbfj+fio7fmAWWFgBK0
qdYbaeSp6Mz685pC2qFy7893rPaGz1VgVFnrPiGG3eMbhgDinbPCksGhKWcp
phunST92QiBewc4eCeNBRJldijMombWxZrNK8cPLPt8Tay+eMRKCGaOQUHqV
Re37AzqFvE9+eumlvMpZSdlWQ6z4TY3j5gLRRce8LMlTmqjPcLTHqUR97+X+
s3Wr35LexQE3A+sxMlAF/OAgJCLDeu7Gm5aviK1FUcn9PHQ0t68LU7kCszx/
mp+N6uo+iyajOokt7z3BspHDU4xEfZ7hhmAhHkbp5eDMUVlzQz/66cOVBVaH
Iq90pWDzIPzxu1g3ZuNc48/dygNIOyedufU1KPLq8yg5jNS1+dPnS1zuH+0z
Xm96FoHyvP1JDeNTMy3LXrRnQW6G9XuJM0d31P89bHeiHrhiiuywp8qxDgtr
6xblx8DzBSkihFLBqsQsj3XIhVBaQFtkdUBG+JFJt+//NFJwKxlxutj9Xig/
l2oE4IULjRgMAq3ge1/u/JgxCsA/W8tEb15lWg85996ZqG19bAJ8c3fRT8ys
btllDjkRmxx5QLbIOkauIBsLt3nIfHUwT4r/px0pZJ99zJj/FwG9DEzVQ0f3
k9qDA6NVtxpOwzZ03r0otupfBrynoAQDga8BCtbFz2jbDRBIGe1m4Os8oo7Q
ia+LGx6dNvw60h4Td5u141j1pZkOXW6jer5V2LRodvCXpFYsDRYvwwCd20b3
9oDla5KXUNX1L+gC7gtF6T/iyznsVlsW0l3wnK+btT+67mgzIZfWdvE8g7tl
LHcxqt2lXE2X7hJY/+tz3i/6An+qUsxGuE+eFP44cGA8zecVyAuwFpVdgBua
m4x4SmNC7mM6wR0ErifqBwcoua2BkxjS+mtoZs3LhhkZxwzNc/r9G6c/JLHO
1OrGVGecuVKWlLtlr3rhwesI0Wv2p7957HDOwOQFjPZho7DQ2JVl+ZNOb7GO
K+mAeVIeKE+0oBo19Ptjav7NigAJF6pgtnNMMEUGlrnn1nKs1MoCN7OVY1uY
eUpVOfjR/z39ae2tdSOSEnLHNyoZl9sxf8Ru6McvwqgFPBi60zqvIso9nrIF
mprIZw/oTk0lME7FCa2NkgHpqlX7jXMjPeceFJpYn41YvaMW1DAxgnbjpfXY
3h1wFo/lThh0QlC32anM/W+MFojQb//FdYuX1Xep2VJz/YC9//aHxqWjWtr4
EUxDmskx+UOt6ubauIW95L9bx9w4MjEUB6uqH3K75yRtXxceea4EZHeMZiKn
p7eNihyfj17shJlcrxYDcJvN2nkhuRjPeKJSla+vmTSZjk0/9O0N84EBHLWv
/CRdWV0vPGp/vG6rK4PkSLHdRYT615/sx/8p40zZMQpvnPnvdy4OaWod3aJT
TwfZzLIfjDproD+pqncMFDq2HdZfh9ZtsW6Fjb+rPn0ZxpK9+T2ZA8WqtvQU
HgFGgBt3mNePjWx03YITQCPgWrPvZPMf48UXToU4ZhG+8t2fctMaVRM1iLbS
UtMD1op5/A6mLc/uftRBCuSgkTyKOdoJfKyRe07LoLzN5RxJVC36z43+BdYt
Jv1hCgIZolcU0Qf2+1PwMpPFVZf0v0SyzIgscsZ3tWLAQP6pEyQMhGDI35hS
mJ+WLXFzwctDGARNZiticRjH8Ta+hlGNxmGNC/l8u/tST/8sxe3wD1QLfT0Y
XjNfI5MWZhW4oj9qa73XEhgY16tdov4VILIQIvaqbU9q4m/pGVmasIEeSOyE
BhtYqa+m5aYUjBaTemFTpcqycU/Hfs7/C9HKmpQZOMRzton+TFrZzTWpkSBP
fAUchnBsLGo01ZesdQ6ti5aOuw0KJ8EGnQoq58j+IhPFgjuFq750nUjYq8ku
TOA2oCN0jr9QMmVaZY8bAMUPZkq/t3tL8BI1h92VN5QKR14yGhFo4oDD3yTs
LSHp7ZkvS+/7eF5+tLv6VZAwhEJ5MAkj0404eXgGcAz4Ce0T5YnH+DCESfdy
GPGKaui9jF9/AXOrgahjBVA7aadFZW7e1dVko+WDjX5ipCRyafzXzUIwM9uS
uBabXZb4vZ1nNbW1q8u49vu4MFgHzftE7SKYRnSUF7pIrAb6mIblkeWhhphi
bwcKveOLLC/qe7UjyqhLSg3ux1PJkBYcUnGp8+RSgI6ZrWayXm1LFoLbrBLa
M7ExUejUqzNeiNJtqhiWHNM4WFE02SY1lBri/B09H3J8Fpj+EwoAd4EV1sYp
EG8XeoeTg3kXXGsV3DoiTc644tzJo8i1FZ7QKS3SvN4C7yLuYWuDyqC5ZhPq
m3vOEQrb6avEatB6TH27nzorTWBy7Q4nxR0+OfQGTwQkPd1/5krvBwKeDIyv
0pNtPKM4O/n+oUOB7uqP4XYp7Qi4mKnDmeVu/q3huSQB0Gllvh2cwfzZ/q84
ltUy46GTzNnSRXT0s7yjo0t2wl5y9VjaE6sLS6gR9fb0QNsYKsiO4p0ORtVs
4/Mx7mKXu+dnSdEpfhDDPJO9KP8akXTPSolGveH0QGOKcxGiIQkJ1j+zRWON
mkqG5FzFV5sThXPsZLqPwIkAYYXrzKHkgmGzp5pYgHYPZDj64V6AgNZfOYrj
Ct8KjDPLqW6kIKEu+z1crbt2oAl8iOXNFAuHNt83ljSSsN7LogYe4Kla9fE8
hpE0s+wdsPmwzZ80LaTk9K62Kk7l72fymGphedlH5gIlOjJuUm4Wc1oJ3gRm
kgbWG4921mKN/o5GCbeLwwcYzMHh+lZXNYWdxQ02jOMicV8SDRY1ViAzqbeB
I1pRpq0zn+v2KruEQpxkh6U5TauMYPCt6ZR7B4840VE9WTMdsE4ENrMxiQO1
ogcyPcOQpbQy76GbqrOG59awA/YP7TauEI8CNKkEF3YSzePfByoXlX6bMFa1
qG1ZMAgua9y5oqfQIdS0JOjn2FEkrbJUy5hvusiil6bqeltrytUC2QB2MII5
e2+dwv+9QwZ2vLZgZjDrrDgy3TvbF3eaRIP3uIJKGM9hlne3Ov6A0ynNfjWt
kUnx+ierEqh8sq2ehI2huAM44vlqQG7FZG1b6P2NuXUPs+nPxoUxnWLHHGEo
uFTpZNhwTgVzOvVxMu7T3/ke/wIK0vMzDvt7zWM5NDyPbTr5RDOnDYQgtXPz
gd/qwNdkCC0iO+ajUVGoyo4W954BRVaFIC0A9TWX+ppAXRLXu0Nvn8Z5ZGOr
sGTzqKzjsGa6xeQYmX6i6p2JSxpjHiSuyEZvma+CZLT7/P9U9IPdkP2fzFkY
0VhDQmmNZmTfXVhbdwdFjLnN3iIl3BMK/u15xEMMMyY774JKELj53cNweXAg
XjQxJqLoG0+ZbZ+AC88X/XybS6JJu7SyUgdqkyS28Jxfu7nm9DP3dtN+9LBR
zrEnRpSmgPTbfirrdrGIZWNXPRgc6nY+0TNebndQiSUmexlQRuzCNceHxiDw
ZVX83MRVY6Rl5vOk9w3T2/w0gQlwWTQ+f/PBU/Hn/gLPfPfGO5SZvVsslYZT
xCPpr+ITQ5gjoi/tCYJLbt9s1HokAVSujK29q5sWpnP64noCn+Oykw3/PmWZ
stl0QPZSkAaMfOay/gv1FQ5qwKNIZSCiPiHgYNQqD9VucZrUkXu0BfnSX/nM
+zpA64S+XFB9ZngsbHSAVf2KsN3ChIEXt8nDNo3syWFvH1MCgiLMnOc8YgEg
7WLpEtcTnVODv2dLmazKxIFefWqNx5iuJSzxVVj6gFgdAC+atSRWrTWRTcdj
emoKtJ8XU+Dvg4uabc4n9YqNnqsURgsjdrV8lpePA3HZPRO67tn4OLtCHn1n
OcTyFN9PLypUW5BoEPli6WNWc+AKF/28JdOfBovkCsViMqEVUAj3Gw1lpBI/
O9jQ38Om1loIpGYfiuYoHaa7tGnd2YYtvO2q/+rA/a05X2WMIg8ud7+Fqtvx
ldVA4cv6z23y79odEporuo4hKgLFEqaeyNC/ndfs0UGXMmGPd9YuL9QNCJbY
MLcc1lIZrHiP3YVnEPJeZo+XOR6yd7nm9wnADhFLruhAOIDpRh6WnS0CysP0
7ps6ws6M4Tt9U0iq7/wMX5T3nFmp0qcg8Kk07VnfcmEQ88abqXCS+bRHhZz5
pZ0Y63Jdo3yfHt1+1KxzxiVN8R/EhJQWQtSu0uojI4MkEAXigOnqXKdav2dz
5qQCmGFM20jRxUMjg2P9WccOAbFiNHUs2b2sUZJi4UUqAp3XoRqJreh8rFhS
h8PKG3QN2yQ/CzhEvZPgsT+XsBBRBDxrWHYUvFg6ge7Fu8zO+Xna9jwwpeNU
9Z3NacCn2yCoE8UGHePwO3kLb/X5wfuOPrKdlFy/Iehp+jdE0doIDL2XSaNy
Us5RJf+Fzqt4pQ+B4eQ1rt306K7SKCBpk/YlhPhEvXDFunfdWhjjVHB9BYsi
i2JzpILB8FglhqyGLf6e6BwQPbV/N1DNV/hgrirytpTMYNqVxQGl7cPC5aW/
qJfyI5+xHNI2SdHHEhNy/DiGikg03JXhDNOv3lYc8gpuRD1874Cs5Jabut8s
S7rN5TzzuwGw0rC7Q7k9xm4kTLQRGqR9lXKAFqWuYN0B86zBSqzTpDLbInL0
vR+h8utuHL8jan/cYpCqrMoi06fI1XKAVqdUdoMjl/AKAj20L2NjMmIWJup2
uOIh7wNGQbEpYM1eor6DerD/LGFQTdbJB3NOahOCE9g2TQqJZq3EmKhhBVxP
cLFgv6BULTlhktOxUe59e8bvRMPj/s5mo9cnelwEbplGdnO9XfanrUVAezwQ
J9NMDNUI+nd/YAVVzSHzMkeqSCmLngNtQ30+KOO4xIEV6lHvtKpRljsG+Exn
+Jf4BFSytIVfyEauUYuYCe/c9HSrE0H+pdgyakRtsmpm/0vSv0bO5MsuoUoT
CDHxIwVaOCny+Ny0Pk6qC3WvUXwXKc1z3G+6mdJjbMagyyTjiUoCfp7j16pV
XaXiKJm0XuQrTv/CPCCF5zMXWuzP/x9+lICkzocidzNty5nmyRghKISSeVPi
IGYqr1TRWLhMQl99u1sDobLJs+yfwkm7TKFmQbTjce/+GAB/49bGl4Sj+K+R
VC22nSTKcJgZOT3ALK4sKkGFpkiU0Dn7ZzVr7U1Y5tyI2NAAtujWVx9XIaBW
7XpC9mLYaKUvRgDfSFqL0XccvAiDRE2nzcsB/r9yr8LgZxX/ulXQlmCOWhji
NCiuE6jRuAsZZU9nbl39J1/vZeHu3s8kYtQkro+UxnU5Uuy7o0jop3BGtz1A
hv3XVI8uv00d1bWy84QBAqw9uYBSx+6wt3Qo6g6jp4VHSLmMwy9lmyHAlfIq
D2Itf5PZt3AVZOhxQaoDluFmgsRqfj8FcghL7466ARqyvh3caxzQftUEt5Pj
d44q4MEyWc8lPIWQOO3eqE3co8/w0cKkfI9PFSJaUUSA/R1B/uy4zGpss6zL
3Yln/rCrzUbS2w8kEa2cm9FeMMEorkAFBECuhH5N3uTjTyDLc4u8w8/9KE5J
1ijdKFrv4mjenqDToCxgLtt2bwrNO2jWnBvLU4bR060RqpM0O+irgqTC2ItO
4fGivs4dYbYxQWgBpxWmUX2NFDbuhL6xLCJFU3IT9hmCLr/nSgyK/ziqvm7E
qHNSEvFOuSm/xgHuI6BUX1RZlH7+Oz3fT+3v/xnYIsDkn8OvYEYjQbyqly0L
EPvPEtGClaNiAhygS1lvLT3UftOQAX1e8ODH3tCoXUwoj9N2QoccWSzK7ZX1
QfBaZ3R9ngVdQTzhkyI2S0Yna2yDvZ6JLHkALNN+xquPo1ib23uttGt+SXHW
rejqvozupsOXvuhA5Di+FQQqIIiFNlVJE/r4tpkUJOGB1TfJ0fQIn0GjWSl1
4oayLtsr8FD6gxMe0w4agDCDHUmHbYOpIMykRa5O46JIuzF35vc6GOc/3JLR
aRwvLdZnyHVgCMfhmSt//76k4NlyBAUTM9vb2JuElKhNb/WjpAU8JEJ9j8jW
Uf3fhu9nQnzIShDP8/r35yR4QLdAHbeUvGVyj+7Fe58gAVUBx0F697lI/+nu
lOrBh7LdtsQI6ZgGX0NYdara/1NNZOmjI5rrkfCQDGlljZvPoiPil3DP9fRN
Nmbx5am/uQ59GQgPdGucgbq1Co+XURxFHGIwhF5wU+Sm0ROtGa3DYpSMHfu6
2PSkike503k9BqGGQ87ZhhH3xbK6KcaURtvdp+vsEO0JXUJqf9ktLk33QrVW
lu7ZgUMqkYuRbS4Wc+3SdCKIZWojUESH88K6Q0LAg5jJ0MYVSR4L5KyVI4Et
4ckSquD5Oa537munNRFfS4z7G2JKlrgZ0hFZsVOqqqmiF1PgiaKw7gNH5KuY
Khhy5K1h/nGKEzX71O0y36E2VaZpqpL3+RtsaxfRkhwSfzbbOsIKxx7al4c4
mWAZcujlRDB3h/wn5j+KlP1fMAQW4zcX2B14GwpeugBJaQL0c9OmU4l9ByqY
tyqin4QXtcNdmUgzwkO1ePOlZfv3BJsE/ynmjfD4c9xiJ7cAT7XhJ5+e5BkR
nUKQwV2qGftJb/FqBSJO3QHYEX4bNOg6EJj+Ve9Bp/BLnR5YR1qm1VcpNc0+
0djQdH7HZJwsXd7Z53lY8O1r+ShbuirGF1s/ZVWgOWEmagvrPfn3sueAfP3Q
h0SQw7WDMC+7jBRstWHWKTaZ24drHhLXIFM/5Lv12eFLmDw6rPTHCw28CO92
s9FcQW2QjzTeeAxBkhGWNeEX1gmmv62JO8fSrpN45N2FIyPfR7PzM8pYrutw
lqq2PvpSmXAZAXjMty4fqd+GiB3NmAth6kUgB4ceygRHIP7jvG3K018eIARk
4VcnvsIk3FZrkqA72qFXsV/gV3duY3qy0t1GsE2w3nddQ9JT3uyV+db0Mijz
4HH/apye34fgW3RENiXH3+cJOnRofy/lIySTqcz/7q6rpbaE6i2rzXrS6kQJ
LOy4PnXA1dLDxX25uv0Twzuagt5FjQebOMxbP3oVd3Y0WabUhxTFUb6yUCUy
Qt4oH8cAprw6E/jisxqo829YlnXWDpiYQDjshOZmvLr49F3bM5wrevanUIqp
woTrgbgjYqQsQBCfbkmR1CrG2QcJAAcrtuR8Tu7QL/kYms1201rX65rIBKDp
aBlRX/J+GklLuETjAe0Ga/3CN/cs8se4dPZR/4mQCe7hy2uvH5FGi3jijjLC
cB15XMgwzTmZ4aqCDC21ckKal1LqThm9F5nvTkQ1pxIJWLnnFotj5LFmh/l5
Oijm0XS8oLoUW3qVkg9O5sGAEyU3rVgKf7fnTH1noUjdEY8TDBgQlTPICEaf
N7PcmpF7cv3Vwnw5a9sRNN3L3BdY0sjv0yM0w4eZayGrKg1I1tZhlFyAiOqv
rIN9y5Fqx31Z7fxLeig6OPjTqpHo7ROtKvtBMRWxh3oh/2v+R/3KxCZGSdiP
aG58cCC0X5qxnqPQMnscmINEjwgcu/V+uyDMQbwZmBUnqlhn7TOruqC0QiVz
BT1wVrRKOOOASojkCyFV0AUhgVITe8NLCdGSqlnNmHAQYcoomYAllZUelIpb
XMHcajqhMVdtOMKCh7SDkzNn3jiYtqf5nj47V0Ee97g6IPmKTEk4oK0/dxfr
unIeZOyO/l9GThfEKQTBNkHXTkjCTvUtL7nnYCLexnu8Pgt81oipYdGByjb7
TTJ+zjGem3jxUMPPP1da41ExAwt8pQG88ObGi9Bbiofjwvh/5LvuH/G4g2ts
Roz0qxrTM69gEcHEsQcOFLNtwqXotvFKAGPA+P0/cttTMaz4nJPHDy+cZTrz
nQ5CCVm1Y1tSUgyBjwOgn0CdSRc7YWfjA2bihHIRfx9qjD+SLdfKhEpoLt46
YPoFuDC1j1xaIOraprbgXdzwltFLr3T+FrDGb3A2sDL2EY6z/shCy9+9kpnh
G+Aq3ALAwWUFpWCKhuSol/m4pZahIIMHqQJTr9ORkGh9OM7wZDY0h8U/w3F4
NLpE6f3FoK4aVrCWQFwHNxyS00nnREqX7laLVJmRYY5ggrS4H4N65Wv5zRSM
gPACwPn5PO7oSgBP+e2mODCzoazh3tmoki4yLPnzZ+8iPoUbW7NLFpLmlRsY
oG+r0dhJoesEPFVkF0p5+kDC9P+mBAcdMohOj+MIBk52u+dppFdQyC0hf9fM
HDhK6ZKQxbs9sDWjui91QHh5CGU+B4E0wbRrYs2Y/O8vEtsTfjZ75tYL4Lzc
1CTw07YyDU/TjdLYVu3MWoDWtUCztbZgcOpZgUkvqtUOhf75lyc9bxTO3jXF
PL0iHgmjkazAjtABgmOEZmGCDSQFij7dk52FsQV6WHM7gGbbtSaEeDLFDRYQ
pnrFPf4LllaSM9sijZMuOAAegKJt48Zrr15BVLFd/lIA1qq4ZirbcNc7WCv2
XU8EaxaUuSvz82dRnJDqM1tKNkvWyFPpNc8YGvH7ksJbxH9hnxQdhKdgrAQi
3ppfhX21B5h2tYOApvqDpxfOcUzMUSwcE7k5Wb7ZOhqup1o/2D+KTebMeEDp
VAqDkqhN268zjxmDFHO5bInqgQLuT0QeU1RS6xNjueDpm4Ca588mPWBsuMMc
P4MmzIqISUg/oK5D643uORY0K6ZmNHIzZz8kHt5oIfouXVP9PtR1xmGqTHuz
v0zrsks2QMfHpOjIxqRtftWZDBChdc/1IBwHc5OvYpeRgjkUH38XkZ6dvTRe
SOmR/5Ii2VT+L3iIL/RPtA/aRTBSzyDLzwL5ZXDCCs72rcSlGkEUx5cdGZX8
UDCjOaJlqRFBw2Sa5JmbD530Zrgp8M+DJLED+08OVtFEWrwftlbNeMflIMae
pUPtr1iF0TGY/bf62i3fGHMoyBbgXl1j5w25+FHxoqs5zjKpI9GzksdXOmgC
gkK4WN/hgcImF4ZVhTy2W2u5nv0HBPtgS3MmQz1sR2nOSPqz2d6mKdIR1ppN
cj+vSm0kpb8ftjtJDvLxMNOzbEobWgFKygNusXlBITJOfebQfPRWIB5y8UNM
5rZrx3nYF040EPMZAMh9rz2gFmlx7s0xBdrDK57Won8goiJgUUUUWOzlmCok
orIodP8TcX8K7M3dYPmOY5mZ4pefPV74xzhH9qpcQBQh+IEOLJ+jU60XRipW
BuX3+hqwFVEdmp3BMBNssE/AqwARnlE18V6Okk+1QIgavv3zxbMbANpKJuHa
acuzoVdpyr3nNtJkiaJFs7j84/NgAqDf0N+rc1+czu6yDzXPCV5D7wK3FuCF
8yMUKiv99nHpzNuUI4iNl9HEGZ3HuAO3aIzF9fWobe0a8pnPGad6Uga0ySNV
m9/kmAOYMcYioEEM34NCfK6rR+L1a1De/4A4yekwhUP99RCsTfttjRIb77Ht
BWf7ZvL4t8og48uABcdcD0dzvkd60L47RljBUMjs07weQnBp0wzotUMmDZJQ
vZi8gLltaV71lqt3qO5bwU7nPiEGUGvj70RXfgDqwwbBCzHnNkU4+Rz5lzuO
7Sl0hxVEad/p13f5p4CbkGt2OBKfRuS1Ns5y2NdLP0/MJASaMdHK7VuwoDbk
KxkyB6nnKQ5pBaHFE9Z4SNIQYIBRxIi+DIpZdSrlX2Uv9ap0S7xVhTon5Tkq
jr5UVu9TzmRb0rMKgT6SAddBP/V3+8yd1Bsf1RV+8Va3P9xsXAM8WqYAo/S4
yDBlLlN4qTdaya1Qm8/4ZMEc5n43wIwm4+ftBhMWZN0zWtwV5lUxc3nFZHv3
k4o2DyyG9avA446D/DckRe3OJXb19lqH6HmUN3MD0Ch3OxmRbZ9OUhJe/tBq
nw3Ry7SD7fmPE3XRYvLqVeJUPen5eqPeh79i+Iqi/KY1o+PJhdrT6JJEj6C7
mVSXxg9Iuiabep3zWw6jc7IO0S7hXK5l7ktsABDU5WhN/5+AAifxRFfXdjfq
QxFnAcJ8KYyQYI6Clb+5HEzH9Z5JbQdgqV6jGQnqQsJaObEhx8zxndp0at+5
NkgNtRtNKLVizcgqrjvUchktccuOjxSQedbDF7PCvacK26BGxiiBtNzT8ftN
yWhvxPFNFS4oXWxfZ8zeHSBVA1ftzgEbYSIIi485EQB37xADQsj7L/WOCZmZ
Uo/N+rlHjbRI5IW0diGdxeii3buPlvpmhjiQs90IvCp3X8yGto/Ioxr3i+vT
bcmpaPvIGZ+cqiegHDpd43ysLz0K/mT2+MO2C5A94ElEblspbj/eI6eb9bdU
zFmT6+9ozLxCm1onnVcK1hhrBbgtRyk1rl9Fi3EwFVn+J1l5VGdry+7kjmQK
IhNMyrGF8Cv6n5AgjtaMErtcr9NLxtyQflRfKJl6eexJLcdKTa1YDNaBaGC5
JIPWhnrNHZp1xgF9vAWeKs3+yfD2DPPhsfSVKlscjDsb+Dc+In479FkE9nfh
rYyaQngeWQx5tvdYSMhUhY1cfIhemCt3a9NGNTtHIGMLfs8cjvie0VssH+Ny
w6j1MyVlw9qMQW6aLUczczcEg9XNWci74LdDkEzwVVaLT7cwC9fI1NUk+//J
2Avk4ARjBecoP08XENsHsHopRigUQotnxETmopwTsaF7TxXJLg+4cy2msBsi
s6PZwdWAibCVCxpukagywZsbYTO+W4Y41qO+ria0ZwnOOlnwz72NJwj9cX9v
duJJtnsWkSJ/8sLxfOBEuYX4HsufEUwPlr2HNMdoglAI3zzQyQPj7k20nAKD
NsILntUxsDuk6LdknAhVGJ7mS1dIheu1eNEqV5p7eKXgZPwpHIPrRB4jViKd
PxOoNFCC1hNULPaouDYO/g33vSqKpGOD1z+bgyydA/DJVi2ernzCzk5x4cNb
0cV9zOriViFX4UDHd86pysBSG8eSZb2SbiHRwXuE+UlL0rvaBk4Y+tSCimz6
fZ9AlozZ0PeDWzhq9Yc08Ca4b4sGkL6pq2EzY9PuWTwSqQoMK/23LP4WL5e2
KizFpCQoKgkU/bsBLDq/5KrDg8N+WGuOd11k+0XoX06Prx6cirFfTTxW2v+1
0D5hpNr5rRVTROKt7cl9fvUUV2QOOmdseUIggE9mp2t/4UA/ORvuF/WwRrst
xfQ4FoXcWLhtHm2L2xtiZHiuSchk+hsSA0A9fuVxTthORvrnyfgnkCB7mNTc
gWWPMSqpeKjdE1P1FTen6RxzXqcSL9LWYBJqpTiuHs7L0RNVlpmsuUbiKmsF
kpz/Cn4JlRU8T54ASXyIouCDj2cWrjv04uAgQg0J7g+D96AXn5BOAL8ddlvr
qEb/YUdX5gNQ4ggtRa+IYZ5dECJF77kw/9hcZKkGD6jyhNvCOGnAcwkcjlSm
wD6eydPUMPcLVxbod7DQkDRAvE2EfT4eIbH6kteEca4wz3+X/x3R5GB0fzCu
Gp8YoQ9dZLFq9EJu41UmkOY41HYJeIljFlLiQ+6OZktID7Fwg7qRrNqJkItM
dis3iSgm45eI1zZf/lEss0x9FFTnV935sZ8x6vIbVjCtmpqzDpEZkK73uxVr
OmbMbMVg7XA5n/IRPMV1fTZRWRVq0w3IivaFVbeNCLvROHpXS3DM76FgtqFH
3t4CCuzivF6u/RZ2fApQL6kY8QPfE8fx8jx9do+5BCwvA6NH2k/Gpo3zS+Un
aqXEDoHC2Pe2nJoa7txSdhlQXuWq7lxk5BR/WsQXJcnBH7DenqSOLMIFLO06
PPwG2HkfGtOAAsgWTALE/TBIO1+DoID4RYPhBU/TFUWQnOqGHO5w0SJ+Xdht
U+j+TcyJibM8nDCz+6riYIVljlrbl2L98jUaQnPx81g44GBpYQypQFHD8wvw
XLoVyUCWfzqakoSE/04bnpTe0+sTntH/HNA6msOXEryaRYYIlsQUwUelefDV
iuK8SGepwjt6n+wO8HJnbK6Ek/ruZmuHT+cwx1+OvSVeAHoT8GPcSMaoGrqx
MTnseHSbnkRuZSH/d0AifLENLMnf//GNzkZ3pOUt53b+cKT+919uK3t+BZCs
5Wc1qNOerKh+bQpG0KA9DglljQNg2W064X/T1uXnH73dc2LIcOTLnijHcz/D
eZSSrXHnOaUDdZLDb2lfnt+AZai4a8k3oN2n0TjVJHQvXMY3vAajlvrLxPAn
05or2ItP17B0QZuFYQI1tRr4Fx6HYefYAE2BZ68WlO+6rPzWZCbEsLLfvAKj
hL9jlgGxyuUc/ORPi5quzu0WcRDTNklik4FCVY03wlSmaZONSyo8l9fGmAUD
Eui8vztiT2R8nvG+UIwwb+whNACMBAW3iHp7rsF936C+XzvIheGnNP1SyhNC
236ay8e0aUgr8BEUBEDVM90utAEDp/p6D54GFCcxDTZ2rxaQFOOsvRZWh0FG
dQf5mbyPpTLeSC6UJnsEErXQvKtGxAORHazDWvLUqjov2TCGilE98igGtXaj
kMBM6Igvt3+QmE4PpxUv9nrQfjghFfScysSv4rOXKvX3y6cLQUo5+bzQPoGa
8dBcIFMfyHrDHLmfpMSumAhEkGTSqg1HS96dc5f5GbHAKIyzC21bVtGKxXtQ
vkLsCNCx9Lk7g6zSmyJRUEh43JDjRPpR7/0fRXSqxxEK6ukVQOOUNXvm/Xlp
HqzAXlHPspOs6DPLTlQ42lJlc7kq7hQKbj3Az9RaPzrDhyUgqnA3QDXa+Vdp
26JiiZUZtwFObrWcP3/JYlM17PSzt2k4asTeIpmkLR3p6KT2NOUE0Bj+1frQ
BZNLXwu6IWG/XPL85WSn9uQqG0dHCpIPjNXCARkVbRP2kgWAqkdtglGJJ328
2nb0gdmeWCVSRZSeZzJVv8A4bgUIw4ayV56hpKjMrPxCmH30v1iOt5HB6xfs
tGCwSd1q8Trg+spfYnDsJ2BH30tBDMERrjVo0/XckysM3rObN+NHIhKgCk8M
ACTvWJmaWrLVmDO4w9jk36n86XJ2fer0kT+s1mqDkVsN0rozHcg9ArPtDs90
pz6KJPxSehO2JjpZ5+1nr2ildxFemL6slBRxHZllHUbw7oCUh6rM3RqmO+Td
GIVbW9nspAndWA8+AgdBEex4GxhxH8keI3Fqtv6ndviQhM3gLgAT3rObD9rn
bFO2/YXF+ZH4dy0cNcVqR59d0JgqY4zlQiLHEVu4+rhlm3KcESoMgoZiE0yW
bdopAgbjzu4x7qLAbV+Alz7cjrwOvY/jXMDJkbczj4iHWnyZ/c7VxBrOZEQc
MaIJE8UBm3H0X+hye3REeHvELsIXsbVQdhK9UBIcMhRR2jlxCIVSo9xBs+2y
aPrKCGpBk/y2qpSe4npcNRxpBiHv0CsXNXnRk0lrOpyk9OPh8mDruJvIZV7k
IxWDDArCwQSNA7NRkkED4QtyikdMT3cFmh/phBaDd0vxSU4rTXd4EASABRjp
S4ux8t728cJQUJqeF5LYYWjbnwVLYSTZemuVGaIbxccEdUu5rMbcN6kyR+7/
K0qDUchXM99rSnxa+i3iiKgdE+/N5U5PocnvKLrWO7V205U6UwyOgZnCx7g5
wG+3LYSSQ9KXIast8Wx4dzsv4QmaAWKOnd63TAKoxnKg/gOtosBH0VWU28VZ
z0LJ6nqBAKAHUrm0gf57diWXFHBFXlDdWvJffYqBLd296r5t2Hrh+1gee9zq
4WVpdCbRwu9Eb/VZtoCoKoHRUPofxBTzAJHREK0doIZqpVmwm2xfby+p1/TD
Zli02zs3wCoHtDT9sS6dxDJMVltbCj2Sx6gIkJyfjc+CWE3MAzgG1qh5xZjl
GcUkJvGbP4Hodo29avdsM4c1EXj3VN9d0CBZ6s8UhmuJIyrCQaCJwbyTCOPg
LQKYsLGkJOTpFf+8HM3u5wkYVYFZtCM+cnMHKYWn3E+JIuJg6rPYsTknVL3E
785Y11FQNuN2IUzxwTvAB5XbQnqEUJSYiiyDTlR3avkDn2uXFumD7yE3S5AK
Wj3bxopiIqE79eOBTu3fpNJJEUCEchMJzOK4amKfIJX6eYxJFZVrKtMeoDiu
vJF78Zlu8TvuEKmbNZLzcwcwiRoZeoJeNBs5BpVE5UK0QytNRRgCTxzxl8MG
0vvEArWQIObylTWkGxjy5YNrVvZ3IHxBScmbXV6Lsmr9gaGw9NRSz1aruuim
a82tdzIB5R8dayxlBGfSKN2yl+IXE2I+qWdyPrgtvYtpHJpqBj3hsg4ly5Y/
IxtqkffLRdxTB/5b3J23dWrKuwy7q6wmMLipP64EOP7TyrOoVIQzpx2nbmSe
+pvJeZuQ4ZyE6naD7EUUtTkqXLoZok2/bQM4WxgFzxJKsu3Fg1/A2Tyh/U5O
LYidl6towVabRKAmgNVUs3o0V5TWsNyvXG9tZTiuKVh2x8kAeEZ6qfIWmIh3
wj6FdsW9Xd3H3o+hJXFpBVjTsUj+CTNVHEP2EkH5Ur18zyZ50UABtxBMlROf
RkL0KNAAlga7nHiSEPyyP4frha2/OBG50D/MWWyZnLe+byeiM+A5swITGr85
yaz0Ol+j9UKSstmP8zf6NBHxRL0fQK3IpEu4z7N16Y3voY8z7YH2NyIEp6JI
XXRgwdtNPUQPjvK59+V3u1BMwmyilPMSTK3+fLJi0yrCncuy0fIMBrC8eewP
ppeKAw0skNwHEz5WOfrbISOSKMi7h+KTVNKyCKPifnfVpSo6V5dmvMtejWVJ
u3SHPBCVJz9V4Kw9QV1vjTejDhgDiNb/SdfQeq4Y+cMeftltNE+iBsCXxQ1p
PgiWVI5XbQgGdM5pahlg+gAxOC8Uk3BU97Tk1BGSIwNb+vOBQLu3tetYEXDa
BobqCzaUpQOxr4FxjWFNSuYPpwQqwaj20zltJVqX9urCx0oCR/2bFnSc1nLV
IOveWSea4ohRxByVAejyRbU3BMIxFp3iDR77vooEXtbfEJp84jlA9VM7FdwX
rDZ2NINof5V3XhA8omNUaB8WrwNh4tZVM74oJ8S/Mq6rN/NcVOvOVqHQCOeA
zet67vHA5aRG5s7Iw4qC+bP1a7J2WpbHWmUCdhS0AhDG1IJw0rpsOknLaG/L
ZEJ5iZucCN/SO9McRiDJBNaPEpWhRSsx7s26yC6UzVcZerAjh61fFZiEUqjv
4dO+tW17zfRzNKaqoVWSAHuueYBPEmWu6bOznyh8TEElEq3XTTdcwWwvPPj2
KfuRFj7yJpYI5Z7vIdOM0UF3jnbbtSYcADlxYxuVfpyFiIPw9/CiXN7KFvWI
Tx3rGwrPOP9Iv8L7hOH5QxPk3jH1cRgjFYhT3NwvIx2NjDPqGHX7gI+NIN/s
ThwF3DcBlwU+6nft+KMGTl97ENoX5ViwBfmkiHct08OIGqYj5f0n7h4cxxfl
5j0HIj0o3AEjI71mykyWqCQV8jeqO13vOFcDRgjOPCupUgMw5dRE6ge46ZGK
IALo0qhXaxS0l3FM1BYEUdl8sn+dG+G/2GYBTr8R6CbGJo10y9TjGmbueaR2
BNH7I7bQL2o7UrKW4odombuS6zk75qqsrw7c95xK+pDaCq/EZZ/hdOo1g/BY
W1tWJZ2VvPSPy/f4T9FQO9T30Xc1LqYWERU+08YSuZsOOVLWEplF5X1ZK13w
qulzW7tnaNuFhxp1NMGd3bg5qqVDLhymgHjzM8xFiN4Z8w6+GBZQGmWRy89Q
2cClKWm4Njp+kbEUxneHV3BFK7gQCYvD7pDjpW0cftoTUHWdctFn1UQqKWlq
EvFc8Dx4meITaPJ6twHcY1kHVb/tamdCBBKSPmRkhXbGSce0XdYYzmt/W9+D
+Op/ns8jM7flvFJtXuDOo8zU9z0/I789lVjSFqdj6RYOx+ybpuck7hcFxAqM
7aSHfOpE4jF1YPa+rbvuaOIQpPX5izZpfYYtjr9yL1Bc8riii+LqrnIrHCsr
nOXIq7CZCoMtsniUyHSUwdVIanjsfYAZKGd/dDOoHTFKLys99L9fG4BQz4Ld
jYm/n55R8Ym43LpaPfJqW+ii1RCVdaWoqinyLKPR7j6I9Wbx3SGFKpHBsKf2
snTicW9QAtM3kjUrFG+f6ctpH5EIW6Bhy7N6WE8zOpfpoDCdGJ6FgVXmMu9d
bkGvXNXGSUSuVo+XJi8qQKqhbRi3p0ewgSCF+rWgjJ1SR1SjldLZE1o0tYh4
84LZCGg5VGSeWDpcjDtJ9aQVxoCbQbM7xfnHWFibmkhRb0rEeJSI+7Z6vP5R
NRY5yE+lhxBwaTGGhYzM7/+IUrf3xkM8QRNfaHDZiNe0kbifdr4iJclXp0ge
3snl1ALLkPpiHoPA2y/qeE/6B9B5eQdb1di7bq9TT0mih0725bu37md1TwZV
9e3+UHfgpet96LVji/5DGuKgb57sZHIj3uu9yaY7/ZIYxP4Tu+LjntAGhcKL
td7IYuP6p+Wl/F07u7KmwhxkksyJgj/jDoJ5QlkFBA8k/n0xQijQy4HShbYk
Eq1P0Q3ZObM+eIGOzOxfbLqzgBdWlxdb5WRpy2tavyDTYl3KPyii2Y0mQYGz
VK6rPBKOD26UC3smjeAXB3vz5kgPLx2QGmVOT2FH6UoHjtc7mxqeAGg3OvJh
ob4A5xoPR+G1uw1ChVXDuCaxtdyWch77qGa+bmIo2yQbhF1UDiRYLfU2OiZC
40cdLIxHWtVsgrENzL2XUTpiO+oqPNAv487D8V6EBrtv27q07AR8Ve7l/75Y
+D4J4o6YOvvoXRPmYdz2Sq0JN1Kn6Fvdy7rKNpXP/2Y+2KZZSMHCUzTXP+xi
/Fgoa5a15C5DiyLUgMeS/daArgJC321AMI7wxIAki1xkqxlQd2xXlREXX+Zr
yApckFc/h73wieuuDWxf2w4VvWe5euZtDtKcNFlaT8rsQ/NoO/Q915uE1b+V
c+YrCDxQgkkVCwEx50eKCOkaejcLY9jM785DwpXSrHUkWQg5Ndn6ASKyp4U6
1vgLDqcASWPdMaumO9+gKlvYyt1RPHid82cRR3aymD5kmkOlCOByeqtmCh+G
15MRyB+RPRJkt73X2P6MflEP8O5pMWc5g7iHeubl5jmlLOG0QXRCs5axbt+j
oFomhlzLgHwRgHkL3/4y0j0XP0/LFOrxNh/SldZ6OxEnjxKP3cCkDL5026eW
rWmwgrZ2/K1HgeoOb50edRv7uRhaJsYfl5KZs7XHijKysZxZruS9hzoZY2TK
KTm8Fq66Zwrx8Xe8sRel0y9XacuUBYp5ujQKfR9M/jxUl82h4ZfUaLqgjLud
aiIeTFTgWOImQ9JuCOtv1oMTcQZ5F35Bf4YvkenFnkxuFbQUCWG7vLsGCmsF
FGsH1F4oaJV5SvQ/qiy3Y88VJvV+199dBV/0/ZE+BORgU5Hj1lBkPcleLBGZ
JBTg4NguvErYCmyEOACijRuv582NJ2Dk6797oQoHiwr1ofWiIZquwusEXY1e
5JSmanu62/W3NfdmTNNVn4tpTGJKcu77veBP23jnn7OJCAdfheHRLxADh6Zl
BDfjQ+l/VV9jiZ/5rbKobk1bCcAPbHajeEZPoDBx92EMUJdbxQblb9DHbFXd
M1Bble0IU9ZvzWh7pXFu+wrJJlb9zdgkQkcocoQ+aZ7SgoKwhy5AZNsoYQIe
OKDa1UOIXjwxjpGvjzv/kiU0Xe/yf3H/+8++PpkHlXbPhgzEynV+rnqGEF5v
wgyE5lj0JhE5JN5Is2Tan1SA/0awtZW4WJMkp1ZtmIzU/9TBumYnc5grSQCH
JdRoLLh4P/QyLILCA3JdowCyDxazixYONLDQzk4Er1hWolDHW6QSEde/lj6G
hRbcgMnApBorv7Z9m54bUH5sLH2LdeMY5nuGNYMrv2iRABm82B1l4AE0gi0P
75Qj0d+5lqNuJri/zKMPM8ChbGk5SUWWUr7Auu9AyfHCUEtUi+Gm4s8GN2Pe
s2NCdOJKZS/UbnGS3yrFKdrVDTsaVzgdMfP4L2BSurhcHOOAnkLqWvhPqGP9
ho4H/ZdpdHgKy0Byr/c9WRFn9NjgefQ3YYAXzM91N1UPkBTwNtgp8YkWmWOd
wT1678spb+pNbnGANl3Sahl5GirsFAZ63zcuqd60tIxbFodG7ST8UqldDnZN
MtBZX4I14vhmckrayvtoxT9kD0msUriKRAj/MPLpTexxs8jYg7UABpZjA1k3
DHEmC9qo6aW+EAWEDXK5sH4m+rVcsz0LjKhPyDAaIn3A8kgUI0tE7DEyo9YI
XILe9kcPZ//dOAZu+FEQjKKp6+hjo0GwZGJ0wzuaP2aOdcAc2pc+ZapV0API
kRp2qObL+D2aTl92pCcoXNSIPU/xekV7jK7aS1VSgsjc2TNggOSL6eTgpQE/
zroSdgzy1S3KePedYaOijAJmKOoCcCoze8+kPpa/eJh2iLfZh4ssQ8/ipb2x
FoMXMvmBlBAIZnJOifBGd57sVSa7FMYG6jTbonNYwvoBPV1QpLcP5Q9GsG50
uEPm+Y3Q/kX83A+ZjBh0mwQ2SKD1EokptdCS81LQU1rnzf21ihPjMuN6x45w
61VdstxMoTgihS4bt6d2R6kvmUnAkPkzOf9Em3t8fTWbIbPiSFzlfvxDZNeL
tP0IQBZjyG57VkpnroDvMbVVmCrt7dhyB4EVjIYitra2sDI4ulXZQLFlqhIk
rZndNMjNKBvR4hTPKW7kPKcSq/CLIL20GY7VuCFDhr250ezjJNOgyxIOFQ1X
k94doL7GC9gYb0KYAPhZnnidsGVtadAX3DuPDRY68LOYDbEmJaDq/Ukbypn0
k0GVYWymMQD3w0S08DKC5buvEdGxobpeG/6fiHTuYNb1Rk7oHsSEpLeJH3RN
1nJdPVphz8fm93+42vNRi4X1G4du8+0en3Wcbnri7cWFk0svuh9lwG/qeNdd
Uf2/60VUSXUBSyRKJPRTQEG9LwwGpYZDEBfsALiMbD/JFsudhkIP7AS20oB5
LmoQkPc3BgXaIZtPjP/GL0Ahyf5oihbC4fvKaN1FwdDQQS3PUaQYJxZY9xxT
xr8Uafff2U7E/T0Usz4VbpP38OfLnU7LSWkLQgqJEUaDc2jJaODZBTaRtBs2
x8ILCNtRGGBSr60SSD2lhvp+AKTSVOjg7N0MPjhgKouH1r71zUCD+57Y/KCw
XFN/tR8t4vganDbt57KkS4sKbtRckhYXc2WY8rl/+iwiJ2lbvPJF2AoHecrP
aSeMNBt46PvdIQNbJ6D7s12I4OQd3lvZjA+klD+3lf/s7pIt1Ow/I0BCI3sE
i6l0tqe+iluZhkPcfTYrpHfnw9ywKCQ+Wfcpn6LytpbjUi4G47UjQxZ9yuyl
eymgTPQhGQklgjrQ6hIc+lJYRjqEWnK3GCtMqb5G8oMu5IKC5zUjO+6gdis8
L56+ov2Y1BFkaO6iMeNraP+I1r3WvjeIXAO1EyFUFauBfGGkk28lhiPA8Gh8
KuLL4XaQgOd4MAY5DQm8i/XeBbiUsjJo6f2XE1e11Lqe2n4qS5CBIm9q7jX8
IJZIZ75WTJ9JayMOmc1K1sp9JwvtNYwwWkcTDgKp27jCmD9ZXJM+sK4i4eft
8DT53yKotoiUCI55sREq5VGM5xK78J9u4zwu+hnVcOhIOvFkhbSe2ru3CGxi
qT/iDJe/1ZJyINB8xjqc1wa/BhgUlnxr1umGQCL8JURBWQh/Dt5ertdAwxai
eBkRZwZs2cca62Ut3SXfOgjTosM2uQNmmUQBjG+bBX5/GMXwlzDu06EnaBPH
eMwNghm7Fm33uhl0gEXR9tDfPuFdxA5C3pNfgsQoCbzjYrEvBwy4q5gJpz97
B6mA6jNiSfg7/dcRQatdkLl3D9RjcI4e5W1zuHP62AVcEBEv/HEWXloipjH5
2hzoGqw3WA9TpFjKmokICrQxF2yF5eOo+/zD26knO/h6n+46gvhdSfy65ORu
tOt7yeKrYsZgzNAGrSOJXX6A5AFReKaZSPCLD15Tm4bC3a8e2hIppzxvi3wu
YeusqcwaT1+CH7mdH5DycvqzhsR3zU4bCI7DJWBzsRgaf9fFMN570FFredg2
J0Tee3jY5wReU8RHitnjBKAsL21FUS2mq8uECnfp6Qvio5Sk0KHkffK47n00
m/oZXese/4OG/WbdJ/JIpSu/+rmXttLDzn5U0soA5vlOIaROFiU+MlmHHygT
/K5+m7TsqaeW6SfsbJ/2yYeBFSpQV3YMdMc4LFuUhmN6mHWvu+g4A5cCS9WJ
FX+8tuahWlaZNBoJ3fpVGxJzjOaNU9Z65Wt85azdR6GfvYZd2YXQ30uQBIaz
zn5CoJApCTW6xRv4uuJ8INwsH61rDjjy+OraikE2oUw54xCvGS3aEc479Khh
3EPY7h5kcyuBctciv/Cuatgg7Z411nEKATLFXPNH0UfbhN3rSYC7AvgwnAu9
4wj5TXlQSHnf8t4TCQ128rHyWmfy2s82vsvQvKyWiIrBHuQ8kAHO84yJfLQO
tY3VQCH7ZjI3r7CigMuorD07jyKqRWb5D+fLig7N/oWtarxj6mCCfqb59IyQ
Dcg1BgcCD4TC6CA9mrciXnZb34PkI19BS1aIZILR8K0AqYaanacMTlIiR5Sz
MfZeleg0oGP1OgHm71Yn/y8tVD01BbT/1fFLTZWqTz6s46AIjsp6Zh/CyiJU
D+jU4SRkRlRbpMLL45DInnAVcIRW/xvKHhcu4MAMuManLr0l3jj+J7fzYRI9
sEnioh4TDNyEkkKk3mPQeowPXGenLWNTPKrcXMHwvnYuh2VKCEu1GzUZiLIz
boj1XUz4r/T08v+Ke062St2vRx5sZYeZbMDr9lWXOwESTpMIi2VW00dOrox4
3o0IZQUUgjqccyMnZXFfmLJbjFh/4vTiJ3xj1UwbPVtOG0s3jwf95zg0U+1J
W+lHM0KJqIxBUYpnq9JDfl+WhJsXWysJVUhY7jdE8cPqCdY4pyIRhimxPVCF
BvaHp40b1mTIVjVMlVhfABdpG2N8uHSNTCS5JZ6cwrvAgmlKTie21EXZFVGV
CXD7Sdo+Tnn544rcTv6yXjmufOjPeAJJ+Re1NUVkfjcfh+cAOXnEQC8MT/bb
cCB2Fu+4enXr7zWY3PHSVf/SoFtaibqXKhMw5VgQIy9h5afx1QjErZ9C/dJz
0DQJdp7mrh+B3woVhbj4m7a9bEgh2wepBIpwHfDBF52nEkI1HOXVsCf75iWC
q6qxzPIWcLuTNVC+muqAe3n37twr5aOujJXxwU0JssNsyIglESbbMmAU+tmt
zuet6YaoskrolDoX56jVH658fr565FC4ua5UzIu/t4TjUg+SA4QBUL1ikAjm
2O3UKA1moDzLqr7Z6JDvV4x2Sq61xEpn0zwyoESkyQxsm2Kniq7aocx3VowN
doVj5wJcm0fM+ygRaWxnslwU808f0cXCHSHZFsMfszRkXKHqOKFy/ZzNp65h
CvRP+qFwZiRP4rl5SJNdp2rutct+oxWEBFJD5I47qAa2LNSheSPHpvnnGEHC
d91IoFyIS1ApWmdnUZRZS++b3Shhxb5yWnlwu6bvcxKFRKF4d8hSQKCXrGpa
fhpobMc7NW2Afh94HxO2X4lqT7K70KV/emuYJKbHjDlNacn2LQ0hnGHBgGcj
cmCGE812jjsBAFAJF6x3eXylntkVbYU3RuEj5cawsLyBldOp2AmRfCICEE6c
VO74mRA5R6/2GYb250v79XV/cUqNYvpm29fOYzOXVlevO+eDWsuGvlwNiD5H
GgoMUzM45Pl3Uuy7qGlyfQlMVOxUPjvjeFNfURVvybHoZ0qojmnNtPypLRTX
9zvWq9kdlpvJnpbiCEhKdAom5VUqNPLfapyMRJIdnSnpIlo5WLuF86RdEJOO
YHUwJ70IO9xdN13aVRSaCeunE/uCQm7gsbricYybMq8VV9ff7xLV6UUyGcb1
xftgoW8faVlA+AUTGFEchLlhzHsBGfM3w3GXXCfEcLE1Ns1CWY8amVsxIyuB
e3ah37mDNOjTZJF7T5Q2nlA8ZDvVnyupuNB+0eqXwE+5oCwhtEcTLexRU7jF
m7MmcDtKPLRyEpBJ82F8qtahe/BxXpScJ9b/Z+GwGZVX0LuVRbW2EFjI/UI9
xSb7o1kf4aQ4bAQD+5TkAL53FEbk9Kg8ZMOX0QeWc6UemHVO8Wuuy/G6eLdu
oK2yuc6WA3iJvKDKOWxK40moNP2ZhBepVA5DZhLYURTs3TfZBdGTkQBgrenQ
ecWC0udL0jVEoJaV+RLVR6Uth/SGOSliEW5x40FMfPhIJql3+44RT7qh0L8b
CsVM2UKiCiPnKe+IeVn3Anv+FvRypzTcIaLZSnllPfSEuv17RSc6hfibD+aM
Jt+aQdwI5YLGdHFVf5bbRRpCMu6SqsM707qgLK6t3jaq62nbATyj9lR8v/6c
ef6i21fRH6fjyXV/uOSyWORtq9xlHiCBCNn4/FdICv5FcMtOC82ZzWTmHfUX
RRYUR9OiN5hvLRvaC6t+S2VaoZtY894WfbT58ox7eXfYpCkzpZ7lSOsxg7Ld
oT2VB8F4Gb8wh6MPiGlDh3HLxzg1Ykn4ZdIT39Yz2n5DF2osbLlz2eyWJi/U
jr3Upi/87sQN8UcY1wzuu++jX+MTNf50wCI364LyM5su4LQUSATuGS0sV3RB
M1ofddByAl7+IvnRBw50EmR+khyX8ntOVGL6OKcawbk5VlRtfWZGUCgSnAO4
apZLTR8hTROB2AQezBt10IiLSBeKm6xbVpVu08aXP3KbFdrls8niLAH0AO8/
eqfg/FwgjlL7MxlnKnMwaHByqwdFqRM/CXrKXVk1xY/2PvGlRbsz9shpxmem
VGpl5Gn2cyWNyv0OkfDYUwN1/JkaSFQTKJN4xc2jxhck2vq+6w1MQRaf9+wT
xs0jjITdI5QOrFG2sIc7vi9llR5qzABzRTIdHOKMUG3NBqvZCMHFGqwcqST2
roZoUAZC77DPtS7aQHdG2KyeDSAirzFw1hRGUzgmG9F+9xZ8Su+qmbgEqRyK
qjGsLu5IVaN8rZZIpFd3lv+0thyjFrurDXpjAv6tHamfd6lv5A/FQKkRQDD2
D/tUE4bep2ZmgMZsK+wn0p9OL5skZHb3I13ryPNeJUzz676G2tsznSA089Cz
jMafIGMNTFi6ueqomlsApxEuqQ7t7jO+GWjXeugmL1ldI9b0vlYgkTlia//Q
Ba18x/h484d/rTci/xRhd823G/c7Hu/HJoYtp6GjW7HPiSEzABmw/5CbiQ14
uYGoV7z+Jh7DqTmNNKf/rw/V+FU0Lu1/WJR9oLdVhBQ48taxarstt6iXA5ed
aSPeai9RmQn537kw/LKrHNH5hgOmm2jKAG7Uvrf2wM4wDPAQraA7kCNAL3NA
E5vMfAgmNLB7lb4rFcFY6bfnhztdFIwqwcrFe4yfZ8y/grwNKX49mR6L/b0q
GOpZEidL84W7fovj5aJqt/eCatuFjj7ToJJifvNkuYHTvhgYXUzSAil6h0H3
5G6lRnxbvxfndEICqkG9RPfpHmZ82TPWdsXWv0i8P9BMCOKbBZRDIsCNqhke
xtFIVS74u6GywJD2+23ReKTS4jNpGZvNmQNr6u9SyimM7dKpeTB5ltuzlHy3
HEVuNHp45BzLAql+cBwPcWaHN3coc9wgDdy/4aGpfxMMs4B+eCyme5vPN0wf
BAhvsPi2IJU2Cssx3I80PPYfIw1kJ80233DFTF5TJBiMEO/auIJVdyn4nm3w
myIsSqw4ubm77+VrnRLJo+P1dBxOBYKTKlfWGCmgSAg8bLwmlGNIZH9I4pUN
dt+rEuD8mjAOhIk2l1KUXTEBwHyOA0qUplWTdODMJDU3pwR0NTWwgghvaqBV
WYOmTtgJCL29FP+laG2MWCuGiDpShvhPTjOiBa0mc+LCByj23LTH8sg50T4U
ODaGkwLByK4xJcrBnBd+32qF7O8LsXYrgD0IoGYmONtxfzojCf7QjOrSlbvH
12RkdGTpi6Ah8vJ8/TEb1s4wUscti+k5DTAcUz9OH3FTBKOVlM14YTIy0OOt
VU5KJioIOHeDF1+HLU19i+fZ8hmaMqzUFVuccHNeKFJjdhjMDfBDCZRX9dX/
yrYKzcLP+911U706BKQxdaDTO/VMa1p+E30CeAWaTRnbnRSl4eNED8RDO42m
FXfOrGRSREP2vFS9u+8AGNFIVHx8eT3gfnVyfWIQeC13OgpoEvVzskSIkcpC
A0VpyslVqq1ApdF1nIle1VvjOWOzUmAyovT2ZPoU7U8cl1Wiul1cboSLWqeR
3FbsjMVV0TuIds+d+IZpIDblbX25vijh1bVvVpXn9WyB4wzWN/C4S9k4lAsW
Jx2XdQvWBWp9BqF4dtsWVDbqEqIGFLkKObJADRZI7vawqYc7YGZNnFZLpE9O
DoG04JPNrghdUWTwbrjKtHgzEhZzZtU2OyVjVAHAvQC/ww40T9eJKBxj/E4I
o/RRPmL4xip22v0I73Fv0IpMGqvk35vA3oS8XEdhI/dY/ukQVqu45d7bbB69
UZBwyu6qGv2r9oatKQ/qbNFlNcDi3PiTRjaOKsxTDqJ1qpYVGmPCodbVJyOd
xXIzosEcWE6SJob4I14KzNmXHKmLA2UgLqnazJIRoH990TxqZJHlUK/fjI1L
ZbaK1850VrWK1dK3BOAK7gQ982jdB1HgLW8++ggjokCdkJMrICUqwIUMXmgI
cT32ojk6gyDqsqMV1km0r96TRTFuxGr6ktE4LeSi6dBSK/xwz93rpDg6k5zO
94BIF4eBUFyuhpfq9N1Lfd9TQ2XFn6IXp1qX6VvzzwtPemJoFSg7Q8VAQrE8
Pv4dNXj+712NOwbJa5DNU1DKXmUzJNh0zNB83R/fYahNxMo5pyEstYLbiI8t
FcpJjNEEQIEOYvD3OKz3EMznhvsBlAGJRoc6eWdLXPf6pt4lCs9H61TDMxgy
7qu76SAOSEWM5rCK0Z9nEje3Mqvt/6pFqs1DzHpTH556NpqiLOdJs2vDsGiP
eMxyh9HkYbh6c1Z/sIIhLiyOi0m3s9o1ib7EOiJu0X8sJLnLu5yEmZn9FMBx
vhbKi9T18BkRGykjaQuYV4u9LcCzRXNx3XufLMZJjZbgRQdEG/anigFn4mFe
4KjlY2stZ8aDN2sOJLYqogX11FppzA+ak65sOCYdFuBImjZa3bXphJh9tLoa
rxCi+mv+lFMNJIQTcRSPW9LEna3t8E64SW3wnrg/PJLAAabIrW1/S3MRp9mv
bJhz1TgmkAwfnDhY9RTJBY0ybggdcg+xiB3OmwNUtfrohnsqkoELQqiIko4k
xkyxXbS0qH6CvO/nRiDlbqJrC8PvFnYQzeHjUW28gYiHLzqfJMXd9bQiM0Du
uxc+d5M0+t2LYoOpYq8vrjObkAFfeWeIu58aTI0bNtkslLAVnCImtYzkCHUF
sQdnVVov6MEMpYN4cuEfp1lyq31bCPaGLub+xGBIYha4c6T8FSBUy1NDiLo2
vv4Cwvn84v1Pgx1NdVFIl/Ay3AdDpGMhIpuMbPOKqarbWiVHs4kJE6pG7j8s
nl/IaSqAyYVbjFJGH9+FxHgORzw1xUoxUQKPtx6Fkh1VRtySPMDUOxc9593/
GAjgh3+v1rCuIDIvjpSo9CA2esw52H+zkZL6GXpr6teH4HQo0tbIUA7Lfdzn
g7TWdU8pWrg027xzCMPhqbGd4sLeP/7bpgPQaesspj4hoeuYZ7ylw1jeoHhD
4o1t45KSRHkr+FacIZtImX7DRbi/za3XvI5p62d4zXoH68aDLgbqZh5IJohg
BA1iczxVi1Wq+2aqEt61ByerT2f+HFqXUeSEFIHp2Q1/TYQbk9R64oCwSP/s
KXUNa/MUXV8sKKb5G7AiTvWhBjlBvVbK1Kc0EW3759NATewKbOw7fCyk01AU
wgxdsye2MOpsXMk52rgDHHrSZapw1DmM5kDbvQw5qVcYLjld1VmqiQZztezW
YthA2xYqpFZwipnDK5oAhx2ipjgX985PWp0qtzLpxcgLFK7/7q9QQMF5YCGc
0EtCNvooO6Rp+afFuZSYdnpOGwCuN6qKuvgFIT3suXOd9SCzBqMKQxy6Bljr
VQVgQuyc8Ugeq+SY2CdOzY04zF/eiu7xWz9RGhJ+ogLrNv+qpqvfPPZ1sdB/
p46P+moK5vg6bk8g6EOIleobdOATK0+OoyZUI1Sr1ROtxjBKF7X21pD49vV4
MPvXaEmssIzb/CzIPbXSzRo4hXDeLLMyxJq5vWQYEKIdfM2L7OoUnPWB4Oqc
Scm/BQfHGaVoDfbv+v1NBxx2RQ25j5yfUzDfI4AEEPjeCR8BVgJltCqRXAbx
Q/84qqXuia/rkC2ma8IZja57muOao64PFEz8POpoFe48omNSK0CxeC0gTIwr
yjcR9gRnX5LSr2I/VLYlNciXu6SitRjBp4nQW13TyPUwF5PZlst752WPMXlE
cPUdRcpxX/nqhnEUS6K5IS+dAQwHnj7a0HyjIPNGjIMknYgKSUpmmZKSfI3Y
6qFsIm3KZEkdbNT1m5DY+RlMLnZm5dCksTLDOhYxCdtV7SBJhAgIyTYHqLn7
2DGt4o2HC5Y/iTIttrpk28T2zMZNaby27j4/PqZ58SuH3YO697ZdfMDIVWuu
7CxwlHrydKTDMk+jCWbS+RIyPPhgTM5ANIpCfO8F4svDWGEI9/eRZUBUXYhL
L4RyxlRcKFEEh0Gwg5WEYMQdG1eMB9M1iKqbKo0GpbUBiedWb7dDTeRQyH0u
v93FlegdTJ5jvJElOwPiLZBjB/Gi+7XsoX9lWUt/LfSk2cv4oz4YCcXtDOH2
LJ9CTHwiO9soXMU8jdgNLIfcsih0SkUbLVUjJsEeVi17pV8EHITN05MiGqyt
tosTj8nraOrGyqcEImV24w8eeh2arQa4ymrRQNhNZE6eCDc+HgJItrGud7eU
es32NUXlsrpRV8TyGfK80ulbp/OuGnIVu7a9N54X691UQWGOUciGIxC2Sqpo
cK0UfVP+IhLc3H3xoMsb4af5i/NDg/rA6wGsrBw0xgABjD/S0qM5athFPGnC
HAgBzgK9/WQuNhemy6mlWEXH4+8zZLQX50fOKdFRDE++Epk9rJ3RX5ZRrDE4
j75tXh2onFlaH5KD0qFYqBKPs6LhqV+RigEEzWsSaOGSMP/9Kel4nPDtqdSW
h9admteAZ+LIl0k6PHnY+Gu+DtrT/3c5F0+vlJiLb530br4H5Ye3pVN6DBhv
19q8AX5sbZzMGMYyqJ5yozUC/VDUT39G0mYJBbLPGthZIIPe+BVtbwmdCvgr
rMs77Btw0b1XiwG4JCpQPoS+DgMYxhFGf610qWtL7H4Sq/I+90Np8Drwef6n
gX34QunokIjCDhSj88Q7BVQuuJmiKrdVh8y0HvwuC/ekGPJJPEo+NlXUcuOK
UFsF/mZCGQXqfpf2ozhYXF4ctE6cYc2NayPvPVit9OclN1GfLUYfKSFU/FIg
mYVQAR0aGN5rQBfs36JUn0ECgl4q1MX3rRoO1vmCgDoFfa5PhgHqw7CZmcPl
CWbjwhsJ1WWKnJtIiKRZQwqef81Id6N8l3Rfq1mq2PkbKo6TOZNUT/0fFoRP
Qz/0jN3UWYnerSeoaG4WefJ17ji5fNkWpL0fM/ManpVKZPddiOvcnqw4MD42
+venweALlJjTQBlsTkEYG4UO0u9hCdcEVrbnEvVCNvBeblvxxuHU4ATWh+eF
d+2QJZ1HP4mRd+PULxfBRBu3aUvr753010LpT53baKPHrtAOgHqOaOKwXh+b
cOfIcPdZamiJwzpkhnqRmhfwKJqjpi4OuylZoXmCMk0b54sAuV2eYy30W8FB
tk8YxHE9G8u4u+g8VsE2mPeVqu8d+cjodFVSW1cLMoLZcAVsTQVwgb8O5dvM
q/BEXaeXcrI1Mt0+IEnsjNlBGdtWnGNUbK0HphMb1C9mgZrQNOPNY/rhf8zj
Kp7bbx+CWM1kK11QjNdGq2W/iLknJgxluJCsGPO/2BL6CWjHomSCd5gdozmp
eY6GxrdUR2nPSkXjXevSgJpr7os2rV3QoEl2R4teaZFD0e6Mww2qWERnIsfQ
BTPa4WRagefWnTRvP5GtvFxpeIqcFhToloGC0weYTsXRbXsYvyfNpeJWV/Em
rfUvdKIvJdRUNtrOJULaSUvKy5D0vuNMx0Tgf0YyPlFH9dJRmLqJV6rvN7yB
Bqu+4aLLWNHNoQKp8w9OtTreTSXlwBBe5WdzFwl9RG2im4cmssOQd8sI5iL2
TQr1mgbjbiKZBLgFt3auUKfazdSGt2my5XXEvnFTNBSSztvAmr35/scTDpEH
BHmljCOqnzFForcsQ4Fo0RKzRsLlq/VYiNZvNGmJCvgePFjsnIm53cE/gxCu
OtsXvPnwoEYIQc+XVgPIeM222uubGyWBvdTd8wAlxelUd0dYs1OjJIAbR2ZP
N3UWaHWZv5lY20mMwjjPPaxnHgCPEB6a+/I4z++Su6DIei2ioWahj2W4DwSA
NSXIrcOXz5y4WRVtC3Ab9ryDw38dV9+dKG2hhe+O/wzXYu6aLs1yywNOjEkh
ZZEmQzdqRqmNHYUtX3TSab8uzlli9efMsStJEW7Mi1nICHlYc8sQDKAnwaAR
pNQlupDSw/wRdsPIDLXrPufWEuB0b8bSBy5GjRLOYX6RlPrzlnVaLEXzSK3J
uYp5Sk6lmP/nC2fCect3xy3xkwHZ2sN5OBXeUJYb0/tUGnCSvD347afxBWAb
WKX2zLuNpJR7koorAqYeaW32hM31C7hJH7miAQqaT+/FHDg7YNwYnSvfScZn
CkFS09Pl/XeSxIcJRpolt1hlahxw7ChM1GrisuwRcS6iqF8avB3lpvbkMHV7
BHNtsQa7c8BN8HwMvRQ+zob5KPeVdSkLf7Wnunlk9vbQ6Q9vM129W8ohI193
6mujldvKEQoAg3W86mJNpkGpkWc4F+ezcJW15FybCGi7hqFTY/q8Lw5qfaep
+/2nt2zxt/wmNzOGOUOSPLloHXtpZ67MMdVrcJzovE2naxm6jGlTMnwuAGz+
zsuweb8QU4unL48mCwbiJEHn9lNzRwEhjnprsCQpUlCqnnaNc4ILYeJGs/03
/wGHxFZX1U6fD7++Ywj/arqyuuG7nDHbf7VEg81slgaMnrKHvSeeWC53103E
aCOjLRWEd7imQ2vjDkb6zBJJBCgX3GzkB9gzJWfJzEicuJYZPwOY6tCSE1jf
zbshCFxrtOXTT6mWgLuTDeV0xmrQHwPzOFgRqKVI8miIFav+nvu9jMKgN+tF
AWbHqpTBlXlTIeFfgMXopGmwJuSFG7nhTugg3t/K9jxsteh4m8iOMa/zfuuN
3u+H6XKDiOavPZYB9oH8TQNjq99ciLtfNzr+5SUe7aV1tgDWWSOTEhu1sltb
x9LWUgRZp9LJEiwL/ZjS2FRljYg5TgKKETikX+8HNfnXpckQazu0dVLFeuo1
oSol9IeCPCYI/zoPn/xo0ip+q1FS9k1Qgeqzed1MEBSFEJQjoA1R49wQAL2E
Ofstik4bSDr/Opx2lTFbrDPHuLOcPBCYMRvfK2JLCPfeTXGfzVzqp7HN+pte
Y+gQW8j+6PZJXWSQWfqgBchxtJ94S0vsoHm7uF8GohBOGoF894cwr9XNq8VO
VJrCI9P3496OMwXazC450mbiwPhrfBnk9BglXKmOF2yR1q8+3+vC9RXmYOix
OiGbcHaBoPCeg0XhKwDpovhKnOvj/szz6WzeNtEPYxp7i2LPgp7HSOxLuVgo
VAJwp03gpX41iSv2q1613y+OSS9prmx0jnsUV6IYB8Z39akYyOAQRfxdaJt1
yD5ewivI7eNXq27lwLmfljU70nOe8vore9USb8UrbAC6xXwVOrJRf1XPpMzy
KrMz2Cs2io436aDW/PEtsyeqyAxmJwFd+kshAAvhXxtWxcWtN0n1YTARfO3d
HncPtCazdE5Arz+22C7CBRVe/dwZJScOv1FnX8k9qFRptNfDIWBDoW21mh8d
W4z559DIsr9kTg6tLwcgoVUSWjwdK29VFlEPPB7evsoLQk8DALDITqg51Lj5
Ix5gUVTQDUM+PBhS01JT+BPNxgOHaa4UEtdDcWVquNbYzQ0NCa7f8zXv59X0
mAi61D/7I0N+8da98GQ/MhMZTFswsVA2bGXe8LWKh5o5c1zXalsRDdY7ky/x
IckUrcEEpIf8ejcCxGmJ/12tCWleKCkLSgLIq/tA6Tw0k43kLlqut7CldrQU
WPfQYA4utn/if3lcq/IOWbk7E5hxxXsCWlqlmhxgBjMIaYVmaV2AgaM7Lj7F
pVjngKxlJAiCupVZmimSgJTWAXfagTaZHDjvL1Snw/ofTpjx6YZyFikD+TTw
uIqLpXZaz7yNDUEop3mhwAOQDFvaPK+y3ZNmRlt3oYkFAuVoq/t6FIVBpKfB
H791QR2t7yRvsLftVs/QvJ8mypt8Tsz3tHb12msZg5nXlTekLOFadV3EImJ9
F4gaMa0y/MUZ6gNQlWJwX+LAG3Z452NqMO3q4VsY3n4TckuaxOqMfAhTEehI
L2zMdnDD1YeHWvEwWS42TVFao+lnf3H1KoTBo6uOPOIwbrHA7ir7SjBLt/ZM
zH44QwtqUvLcMj7uuhBhP5AeGYqjsV+1Zg71yb6F4BNfB63bWx1ff5DlZohb
aobKwgzTBNmOVbcrz0rckvNiZc9fissQiDQN2ZFBdm+J6LhWm+pirvR5ORE6
hPCEeTcuIbSs2F3gJFVAH619KWX8EbLfUJaSVg2J7v/bVmMtal2DR0SQpWeZ
HkrsybMnZqWfToCfbxAoxRgnQsw7m3pjsxk4X5Scnl6IZWlIEZ/Y1YU6ZZJO
NiyKTcrVOa6ptfxse1byZrdI0ietit+sgB95EthKjz2op5XLiWfIlv0MKMd1
YoqjkvlWqd/RdFsbQ47fsFnvRIiYnfUzoj0s4crITCy3NYwYKu/imcwebO41
f8P8iInCc6CuXx+MmAXwJ+16bDtJ6tzcsGKPVenZZ9895Q3ituQsNONIV5di
26XFucPrew7fiuN1OdHhQcdvA5l0f3J54002wOXMCPro0s+ExVv27s/pYTC9
kVRA/KUFIl/STXfIWoa7krzXnRocS5Btm/NOcsz/mA/TBqRlx1nYxJXg1gwL
p6zq4uZpJ3DldJMEOW7ut7uxs/MZ9onBXLoYG1BlhkpqNYi/3FBk38Yp3uBL
nFOfEqmVcAhRvn6WRXDl40Mh1JaKbS7A3INDVOYmDLkLhOcCD99/y+BtKWjz
dqYOKYJ+g3rwKkgAIGBdEOXeIcdJxt7vj0kx1Nb+1uz7lJyi/AgsiRpQuTrE
BbK2jRsXWDF3Wq+sijANiEt8xJQFxf5DGx+4SU5zbQo/WJ8jMmyfg2It9EFs
Gw8A30ViKmcIOeti1oK7ronTN19hddr15T4Rk0WtDdQr67+n8rxpIvk8fOqA
HFFRjyz2vss050lq7AFr45ZdZ3scESyvd5ZnVQxYe6BOEt53dK7ZEuJOj6mN
o5e5vBt1TG2qdoXR2SZVNMq7C6ONZDslTCAui0walSpvu93qZGlnkuqFmRff
wkwXOTGd3jWoVMJ1cFZ8Hfpey9vXDCDVdQJE3FMas6n7ZJAuFmW3yflw2MSX
rEfguc4JCbLlj3V/QVtK/VhLpQa1451s9EOR68Sf8HoJa3YnDiGGpBKcsIiK
AL2YcrHUO8dHxo12bB08s6iey7z1H+EOfKS+LQd5vMxDknz8XyhNZvK5n81F
CAn4M2d0Y+AHX+bv03vJW6nDOg1nLiBpdeJagPFe4CnGK7f2/OhHxJGlNaMd
n6v9Wy9DkIoWQMCPFL+px5Lv1hMw88ip8E8xmSeDRmCAv8yVXRr2U7KuZcMr
FxqH9wX+5yRJGpmaXMwYoVcnhxcollV+1mCOwEsy+uS2bv7z3T5+9R2UiUpr
iKC9Oo4awjqXhDXDEFy9NZGP+iOz/VY8Eq0fUf+Rx0NUchKKRMtWCPB1M38e
wNp2NhzUlp58OZ1HsGQTjBOYZee3QHyOUbJG2Vc9hu9uY9sjfUjCMF+kAI7I
EvABlL+jM0QMbdgJpuS2RYy3Ik3ZDaMmyBtpK9dtsjFB570NV1/fHXFa5SBo
5LkSXSxOXhTFnr6nYcE9F+A3FJlD6nlqb6U1F+1HZ8GXHBCgzKd5uSWFrU4m
SWmlKByp+M+RC63Z3r7/6p1ICUnUeYbHKzBZ5Xlk6F3Ine2vQiGAtUobkjNR
6iUYHmCYMHz/KfKLr6T3g3XgwXAou+Tqtc04hfhEcKb+tykePAUt9dC/lZNi
TELXXK8npKJVE5GGyWXSO+MIvVsxhnyUI/iZzogFsszl1HEPeLoZ+oJUq3Lf
rIb5QYahVw6tu+bvvqCRNfYOP4Kqokf5stXIFA+L78vYLNsr6KAl9KmGjYki
9pQh0MfarrDjPDdFRjNwl7b+glYfT5MFZfXf6MhPZ1sqVuvOtTlaGrdzzMlW
5KrlNkwI+jEbAuPei9+Law03c12OgcEOYw+sxU0oXd9NJmCWJdTztGI2V+05
1wZDoicVbTmyRTXsBPhJViJBc86iXy5E2ghO+vyqrBznp0fXD936STky3zQP
qcJm8jfauqxpXP1NdLqF5QXYg5d9PAhFH+qIpX56SB2Iq3odT+C7hDah3yKs
ZBWJvZJk+oXlWFqHm3Ruh5/rYcXxnTfuLtbCWYoUxtKPlSA+ZbRYyTsgGtub
MZECdDOyp313RhExSM5XccwAD725lYiVgIi39JBr/KOzqJC/zvfUxxeoLvhE
IImznacXno/vcEqazY6o8p9tMu4gjABSDrGHyXa2ObtOpDrifYwFl2LyOdLY
Hjvddpy0s/r2c5DE89/BRkvEr3EC0UV3g4z4+tatkt/VYa6Bz2zdodgT6KmI
POlYrg/oIHzxlD/TfHGDn3fjrBbVZ8iH0xKpLP6PPwqVfth431ytqMylku+6
3u9OcH4BBrAe91anOPEm/tH6ykZJsc8sVjACO700yCW6QKswH7Ui4IKUoBTc
x5RzS8vwDga2uNqlSvpIwPoiPjUjLctr70MrJe7YBinFMSKU22MrwTYWPMIt
1psSZJHaS+TpF8OcHDB8eZM4Ct1vEBNLjz0hsORsatJiubArQuJq265kM3RX
K7gxvM/Ffqr8n10nlsPuILYYFiteoD6mW/nR6DaYloIne6qe+BXkc6ARG8gX
xPpjj7bKXQ8XPVxXltSFthiVANB9B1J/BoM2x0PfmHoaLtvC0pGoZ2Cxo/CH
1UtcL+oVrmaUEDENoOEH6oEhgy2c4z2dz9MgUPR02AxK7YNMCUy7WIW0Lee/
9waGm4qAnY/hm40vMs+aNP+LpxtQF6+zFcGuMxSGjQ8XKSuY14QltNMzXodc
NsnUiu0ISxi/IwxUu1vEbwACfaPmTNLs3GCyfuhy6RXTzzZRX+RBZdTMvEiB
1IUk/hQxQtiXci/t+JRss7EX05wxl+2pGpjR0vYpDP+qMhQ56dagF/2bhE9d
x+jRX3xrdAYZ1GRaGza60yDPy4QDzKXbDpBroIs38QuH00Jy4mm6kuCCa2iD
RiHCy0b2pogkTrhlcLAFhGV2WMTLQRoQCRYrllBHCYI0ds2PYuzcC6OU3neF
+4VBl8IYG8izHyVzceCaK9Wqj9Gyt64RUZFvb2VSr5MRvILK9m6TXOwhH2p6
/E7Xvx1jGzKuE07TCwHHgb3zwTjFOBLzegKSedlF+CpAK8l6xzI0AnLALYGx
VDYNYGvjVscTWZCj2CNQBnUHZO/IW7loSZYKfHKT5pjogYaxpAZwwbTIlBIa
5e/gJ3EPBAPuPk5c04OfOFMsUbQro7xTX1s0+OK1xjzozmmt+I+AVcIAXRez
gyw/+TfMOZIb+GCBiU3GVTFeLJdnYMyzBbv02zKD5DPAmsJ1ebirj5ewGJdh
jIynZ8IC0SzxlOnR7DpN41MgNlEk2CNyLEyNH//LynuHCSI7fUsymszYcstM
017aVZbuuKD2UouPahAb5S6dz4HpY/TnbcKNIiUlpcHzdSPKKt6z1VeGPY7/
G+nP1aN0P5ZTexdumiYTkkTz0bUTv+nr7Rxuww+gd1jGa63nDujVgtund4Rl
5Kc1GE5THTlT6I0J3p2vYT8hLJ3cteW/u7RxDLp3FAXRNtBg/7qGss3Q5KrV
iuqF4QC0LfeAF3lsKWkL2DlQZyAR05Qw4WRtjwetJZCpinDkcb39rkgeEyu2
mXz+NCug2KA5rUY3GXNxmuDi2fbR2U4ju56cIt4F61fdxZwk17wWGbAcYCrI
UnN8vRKQ/nezpPEfkfelnIityGdKmV8cSfaKWHsFO+LXClMp+7b6onKAK8uW
+2h4W7Rlh+36/qclgMnug/o3DuhqNGOfFfO5vCwLwoLFPrcyLuQMFKNLUwhZ
zMQk1gQi35CBgvUI9MocHHTfGKpI4M8EoInMYUuaGwnSE6OEx6lO2Bj6gQR8
qNxIelUY2HbvC2Jsy809/6r9eoLYdj69lylqymuBTXNOFG6zRulZGCMJxgha
UrFGFQ5R/9VHJS+Z+WHTspLm0LlzaUEa+imsPLibX+OyXFlTsNPKdEsehF53
oRloow4qd5JVujZby+j949pFngWGwY2aRwC5x3xfRvg6tzxv9o+WyZRFSo6L
cQVHFFdDFvl8mGB5vG9uRmWsCk/kL1tz1wsw1X2Zst2J3+ITjsXIO9Cm7kuO
1ONTvj3nNaeozlysumZYH+IsIhYuavya4+T6AOoo9kBsdi4lKIiDuYBqv89y
Tv8VBLXfan56PG8VWb80gWWCASt7GpBXKyhplTvBK4ld5Pnf9zwW8CraPHRW
HjKx+sADcRD4uQHNxzqVgZek3xu2KPriyr172yYuYf95uOjkoy0VbFfNTTI+
Y1yR7Msf18fbnc4I+0kWG4KFXpADSxOtQ2YPQWSR5h8CEwg0V7WrQN/fYkzH
OvKupobqJMHdbBfUrd7tIF90NGtGyS2ME0Fuoh8bFmCO2MuynFKIhsAEnmrm
dYthz5C+woU6xi2br+UekmMzuUcG57EQXBvzJUoJHYmh3CbT5ZZK2OFsZiSL
LBIwDSRbHtNiSxvwZWZmwJgOWvlDIlM93rl1bc9bYB34uAlL9MicVr+F8iMm
ZG+rjU5GY3WHy6z7eTq1sois4LjpfaArbmrxPhYcH8YyQPp7MHD7aUNzum++
GNRSxwNH2pGto191fuAfPEI6M4lpEjf5r9iFHOfPK/Mseyc+Fs0k8hwo/RHt
aPBu6pkVjBHFpJgvcqQKYnEJ/cioitZvP+1A4DwdyTd4/DNgkLq2tDE6QPY1
NKyFoQHaUhSnYYBYhBM9uZj2RDZk3Wvhy4pes2KRpKICiDbnb7rjnlnXanzZ
5vX4hVY6ICqzdesIl2lh2ZNkYfYSF+PmI+UdSm7WkpfcLcaYHvSK9fKxkyIX
DF7KJiNwU07nnM9yi+w+LHV+buTNdfEJT8VYbxoGKTs5N4C3df0J6JuCD3Mk
/f7KfQCd+GPJq0ZhWNQS6X7zaI+XMiKv7dJtp2CvZi7uVbJgrxqRvb0u8M7J
CgXU/P2LOLLtOOmj1qwHKTsKEtkAGGGkWaQ3exSzWiP118WYd2fuboOF0vY9
8SIUdtkqEF1M6SJOv7hCEyHtgy4WS3Ypw0NCLwOGAgWMXRYez98o0Ecv2LJ1
43x9/QpTP4ANsoSLFQVCJvewxG+h0WMv/xOaxGYWipo2DskKq4rOWxWvxuLy
o6UStKc9OlHD8m7SnH9+LBrXJtV2m6Raa3FRos66Ftu148LLoEKU/1G1pN1c
Oqf5oPrzwpMJjwq/VpTMlZIqP3XswHhqacxgLYaeLSX9oqA9ePj7hDwzqHx9
115RMaw6SNAYZ/p4YpQ71VMMhL83OGR3Qfym43boyc6BF1Ub75jrt4q3Ij+V
r/YiZi9VR+73U7wsFFH9HY5IOIs5z+rG3c3DPeTJ0e9ab661mC657xt9YRAN
7B6m2f3k2wT+MviJ/AI+jvrE+mNo1/lTqmyIL8w1ZWPUyI8yFsXSpmDynUZy
BqaMbrhWmE/5OabokFRCh7zJqR3abOmuBXED/Oa8dSWsQWtLAjgjxbELxA/A
qNoKX+L/UcrOjYJOq8LxLHWf1Ksadb6w1QaBdfi7FOsxNNIh1t0yeCQJsyYp
W39Y/fE4/Um0BDoE9r7pVL70qldAZdmBVMOL5Vk0ZWOtJrk1Y4mHMJvfSF55
viO72kAwXlK6tTsYOehwzj6RsiOVxzuVv2WxI6r6TPKpQutedbMxaXqisFGu
l9UCb7YaPgB+dwLxi9PYe9yvWyPtYZ0WafnOaJJKdOvqrxuHABnu7n8tWKy5
G9YUHx0acQ0pKKf/5CEC2rgYW3Qt8/gwW1sNxhsX47fD4fwgoXhq/TdUvzzY
9rCnSWz1rgFU5RZfOVvyTrU/UzO8rh2qR3Y+PxkWee8hNBMQFoexrC/dr/Xy
UWOEuAtrB81MckqCA7S1/qm7/QeTo2U8oYy4o/aKQfXLOPfwqsmvMvAXUA5d
OPvpx5Cmpzv5AY6CK+zFGKBMzZJ94grPobOIQ7uSPZvGlEfOR415iWsiY58/
WnaFXkR17ZZh1sjUWBAaeE+Y6r7VEVXQta955FIoMDjjyyIL801oIVcbhCVe
WUv3I+v0OfFsrS57oX3RfCEgw+WYS4nuAEyXcySgQK6PPEEQku8FMcAeLKQ+
9p4ww1ma0DbY5slpCe0i3W1VT3Ry+NyXuc+c65DFvLFEaX9nAKdWhQzu4+50
JIkWfZvBxIM6jOogSIWNXH/OTmZQPsiKIsEzqpTcsG634gZ8GnJSD8+/o3zm
aCWwC9akpNTRobxM0LaFiChXMJmxemNY6gAgEI4DbkdHyu+aa1vJdxM0EgGp
TV3Ul1s8vUx5lAubCCiZrKLACQ9UjKh/B2sdk90bm6gzWYQM8DH/kFYPFkrS
f3HunVcRYAkm+zDaL+E2w26GKe0it7VV3BIpQd4yoB7RoUkcATTC66gCpmbe
Lu1khNUYHGgop3v3AjjbYM1QO8V2YhaqZpxaGeUIaAobJZbSfhFr0wjkbBT9
X+lOkPkYvK7ocJef4jPuafsxnI7WqNYpT52qf4Q+VAzp1QwqR33tJ6aI99P0
quezW8XydMKMZeqHpY5uuKZjEEHUvUiayRbw81+B4+GGup5zzuPCwrAJD67j
EMjmVGUnN7RuCtV13Dai0yU7jhzHXJ13bwmTsSsnCzyzbZuH5jhZNCmd1lwF
IbVrG2JsKnWj6MsojYSVVNIBulpFOAiE4buEvi7LgPNnubq793IXnWHqOWmB
hJL0SKx+ID7J8J7d34rk86Zz2/xIHWVlMZPs59rZ/XtwrhxeF/Hps4Or8Sqk
Lk7wiv1Y8UWbyuh39UMTRMoLiCXZ4lhP9F3Ss5cgcXnVzMH0BYv5oVyxrzOg
/Deivr8f/tsrOP+9OC84iWSgsHBBKxwQ8LWVB0icquka2pUQqf0ImMSKW0J7
jbpRhfBPpJUBKXQWwwUP4OW9seRlipMRly5LajnYXLYe0fw2reU58NKwKOZA
XSJtDVu+tWr8nD+7cinaXHNirWbcitGFSVOoC6sPeufXprlihsiIicXvfl16
VPRh5A41MLKHHyu7wbf3nIjGudi/36UlCPchtxuVEQDZcYd8FbyKm/LhoU8y
al5KeIiBH7TsnycD6c/TpQ3zA8TTzXLaHR/kYLoqydT0cWOphC/dBml1qDnJ
wOeLKjT6ZHT4Ls4jaDK3GLHnsgm990MmVCd0AGB/QyFfeBBCiPEAD2kTGR7Y
5VzvO137df9ke5yU7W+Jz/j+XwgO71XpRGAoEDyTx7YOpZwLMaiBQCTDEEGs
o5RVzMyiJtuSkN4ccEdtM66QCJXG+OKIYd+z+EYHqTsFJXR1eNTr5Ss/G9G4
TXIynJbKhtDO2N2Hs//nZdFB62Wx+phJd9KoLnZ73JShghT/FXlafpMqwP33
NmDIFcKXvtcfultAjuEMxCEA7WMtCSAbqXWvbwFAi3Z3kBtVsO/EpX91Sau+
FQRARVvx1yN6BMFZJqT+y3rC7JBK2JfTV10bN30OtB0PRlsdoB5qkaGAVm1y
RXhi1gGqcoPdY4GJOumarJ6sdQ3/dqynJqhqOJhrETS9hOA9YntGGmLt5oWJ
xlv6oJdDEsiVLNnK9aUq60IMEfjsgROp8++OZFoWlJ6anAaWNL8sTdOtZ5AY
0zDYQJUd0iJv43y7PSzKp4yiiZEDOd9T1VhKPbNEQ+Cy6zuYiHwJuYGlH54N
Gt1SxfPJ4YEOdl2yRWlNlgrfopMete/B+Mi2jgw2Jw5xSGAuDZfybWAS09UC
Y+QN/YP3tRhOcu7tg+8YrjY8AEyTdl1cz3LmBrMeuSrveHfebSxnzCT85uad
TRCkp5isyp/FHxZCl53XWBGnudZ1W5UQNZmODJTzSYNELPr6apFzuDMoL5qf
Ts1ElCjnMiKKt6kjhAuK/TwJIA6x4O7G6v/BVDSbnTayIpaDrYQgRkiqLRxi
79umGOGveKcZwevJlSTZzYzN3ku74iQrZ4EGVCz/P2nEdC/tDVnsqN9JrmUG
pNxtbMgJl/pPN18C7qnlzrYvN5vD3JSoVrQEqON2GP003Oco45COhVXMvFsA
gOMUGgLt+B+EXf9r57wE2V8Ne2tY6Bm6TRc3D+olUXNAabMKyss+Qm04v1Yh
Pm9vnjMPeVR/tZ1EnX/GFUF+5hw8F/uBRudTwRxz6UWbs4Ke9E4bwlHEZVOb
+BFXFDPtVUi23umsnjCLpEnNJOZTmzHmz3QE31WfQAIYgoJQEWwu5HGlVcqa
1uvyWjbJ+yVoMLOUOApZxcz0CVTq2h1ODUPI8tB/o+zidWhEHkphnHua8tZ3
QfBaQD0xKQF2xGrJ5UKRzlLalgIe5SDCjcdovN4Upg7TWP6PABgMmDq5ZTQr
c1Bfw8zQWQNwrUL2ZYY3HNvUzhHsgW8b0C8Wh4X1FL4AOGERevDeFQkLE7Sn
i+6Sn2BqjLzXtyqKE94G9UfAWHpnLTE1O4suH/9w59FCwXcXSn+3O7AV9pjQ
8y64pz80fpPQoYLPxC/ZdIlIRCCyi9Hgr2pGQ7yZnFVnWYza75vUSxm9Rkuc
jSqS6RxhxVfOUneC4D0oDhsbYK3V2UTL5H5nmfRRk2/lNoVTnb3G0wqPxzda
aT7HvE8oJXGoJ1v1XO89DFixBT6bUsovTUg1gY8+MsuLrD6db56QHkNm372T
y9RxPGsHtdQiwXsM52lNCMDlRnMMfd9mf1W9zYZRSFxq4YTw6aCT+GxYeUJp
9FHvKrjisPDPmALD9WCs4yutf6MJcVNi2+iIdssF1kLKZFMSNszcai3Dmwq7
z5i1akpS8tgbDDgv81XdKAFD67TlUTiQDQ5zPADEjf8ZHoPopnEAzgWtG1Hw
mJLtuxy+eB+dlJHZ8mWL7JNI4dUxVVSWLYPGhMI+qLveOZbxX94zno61Suem
m3JiFPDxYLpsZGmLcVRsaKD+obaHgy8+aKWtV60HYtIewDCRRhu+WGxKNNhi
cndj6q5dQaVJD6mciXVEwXfmjY3YcGHKXoqhOe3L7X3yqMPfM31Xj5JcNSTG
SNGRXPvZFPBoQXg8D827S3JSzBSpJNBF/7btgrklv8rSkDGdiKvtrfV2M3to
6nQN0Ge6+Prsehr5a2oldwOpo3Ma6wXkmcSGhN3nV+54CqP0LHM5214e2GHZ
YKMyJ1pQz7E9gbMysxSUbQCLegvK8PSJsrG9ejZcOp8dn4J9X4x1rjfYMCbx
ttyrgNTilKRcHTsolW4LZXWqdBpzYN2W+HM3WWsWddDBBORdzD7mgd6VkGCn
gHYzFvXeWtke3U6sed5+yQXYrng3EL2Id9TxNOmzmcyvaDOxaCDgYEwjrHCE
wJADirdbmF774o6WeGVByO7Hw11GipMnh0QJOhX4tmitcSazZGNmxO4NvyUR
Jo0N1W/141t10z9JvOtXkUKII3VE6DsTz2OzxqJatoA8ajZhDP20HBMLnlTi
Pz44Jmtxw9zBHN/x8vC8m8zGzWGEz2vFEqeYS0z++OHMxkYoTMstNh+MGC4/
K9mQL9Kgyo2iuoXOcPciVFPL6rM6hDJpJ5hWarX7w+38xvdT2iN5e31bXiqA
LS7phHRtyY2glmXnoqDPwLO8Pe/UTzYmfurLbFzTjgJVQy9bOFxWx/HWS+VA
tONMsNWkvzDSgwBPv1ppU5kg1XXR8iul+NGng8WtOmRdE6MxT7L77VEzofpr
Oj/OXvPR+WNQnFAsOso4qEkndtnuOzXGYJAuGBQKFYqrrYEUfSscpY3UHpBH
GT8IOxS/TNC4gGvuZUehh5BrBP7nt9VahuLj9wuVzuGB81MJbXO+JjABpE4X
GNCa/eypge2AzWbAmbAtxbfuM9/QdfryM7tEhOlqPZUDTbTjBIAvX5lpLATi
UrxdB76FiKEj/HT8daV3dAn06ypGIv77Xj/kmnPsNZb2ZsWxEssIyP9D7Amv
IJMyPlSAzFsxo0emxH0QhVaXeV2z4MMWvjAyhoLqMx13b1PGpUCKMptQ7awO
0CMHXqPrNI8QG6Nmcc8fAMRrikPkDpYtZk3fv9gUeXTFxB/1vRMjBCYGyunp
1tXsdyNdbQ5i4qV/oO1NLdsMQVM7z7MRFL4cE1OTR+MfXPUy6XZzXKeliaUR
386OgpV4T7yeWjCoMl1OfzlLnP0USl4grkGH1GAU1ml9+wF34kwo98Ri+4eA
A/PZPMtJRKxy3CJY2cf3+gfEgXOZcVkg9lHYVIlboSR3O1EaLoDwBq2GxlDA
gzlk4GvbX9APTz0iDncDu9qbokQDeiIZick20BykVAJ1+g46qqflyMTTWGHL
6O3z+MZSGrc+9EzfYFd3H+FCyZ8iexsKIZgQSxg/kGVAjCQYi77xAuLhUlAn
YFKVwhkRZb4ND8PTQuQwFbsUbmCHP+e7kiLac0e6hZseJBL9RPweMN1EFIVu
wn8TnIkDqLx/Hgrujz1EOJ0jPfUM9J/SFlTnIwsRZY6z5k2xdiiVOaMMn9gS
V4dy7UVI2SH1x7GsfkmAbzq34dF7VbX1v/1b3Jchp2NF0ISF47H7kpWjtraV
XP+BXgmWb3kClnGCdSoq8Yq5jh1Lb01zBgqJCXskiFr3dCigbQVTLG5Nsc92
EGowYjvW/CoEM1gn6+VXURYkQuXYrlRB29DyU+Up7OjCePG6YLlFwhLbgQTs
HMKpdGfKNnIdJUa/rBPNOKSmuweFoYOJzA7C52qpVLrfqnsJabW6I4YBgFCP
Iw8+QjCGgY+DgR+0leS/cxdXNTLCu5xUMY9bi9G/tmJ7cdlWc3SLdGYNuCz2
ZPkc1RW+A/bbGvI3M0KFUliDo1H51uoQZao6Cd8HrIsMMZO2tCUPXLjJCR53
XkwdcAay8ZA+8dlv8SU1dNO7kJQEYOAtFyMbNNJUd8xZcN5pq404lHt2PZbm
zjV5sLaI/SPi47zVbhhSwrghUON3bICf85Jirk/Ls8kWsfxfsoOaEs67G9Fo
uIUm/YNMWr2xrlVJyYgKrsUZoC3/ohlzN2p7dm8gJEvZ6rEPYWLg3+Nsdp+F
ajPrS2Hf965rQLlsQOQIgfV/sNaBt789KQoWg/uhGRr0TSGLMfZSQsI1/xC3
QO66TI82GodzL3wzy3/piM3o90pYQLt5zsPUho2qIEcYlW7t6msC4dlec5Vp
eu8xfWZZoqMISMOtBybo9HCfxb122BIGY1wt41Ipa49sJrTG9u49TBqMcyTH
vE9+ZAuAofLM8Ojuy9b+FbA483Ds19fJIUkcECjAntJ3scNQUd2o9X5nTKaf
MrRYuY423SQ01N+XOuCpeqTfS1FBc4oKr0zZYzvuOJgDQOIp6AVf+PshzoqM
BEzFvDt6hh1LGJC7Ih0Qq0iVDzSPeNjA45ZUTXd2t2+1e919j2JcswFPqXr8
b8cwgSGtG34ZLu9lYEeUA0YXvgGwLtmaQqURuZtHEM0Fvm1Tq+vHAllVJx9X
lfj3WlZIoTj810DdOfbpa/tfr/s7oAM7GGye0LC7VqnoJHbrQ36/Ly+ZpQtC
gc3Ws44uNdQnxsfg5h8P+sOE/PnIR7wzOOcBf4zLLqwDnkHF/jZ1vz3tsOLR
BfKRdBZqbLzeSH+SbGG9yzhv/IIV/uDxCe9VrFNECsGtGHrgriz9Rlz9YguE
pQuTTAFxxR1OqAQ5W73U/3Rv3yRg3Ffnqgbi4sG2FL0DvghlDxbH6UL6M+4l
TFjG/zMlLNovUKveMIUpXONtFSpm5DNfBpO1jRnamD54I9M6M8NMiiap/QwQ
BWxuZVX6vgujCvB0VzJAdAp4DNy2UpT0L+5H6sTCrGxNG6bfrcQkPPzp59Zx
fHSaTyy6tptvZflZ4U3TYokE69BbeZfv4ucQO1nHu7GBj45n9o1unWD/PzGR
0GxlSpzTnG0e6hJVpX64MQEpuFUjJ5nzw+Hs3tw0fdt3zEBd2gMb0a3rk/lY
Cb9yDXOhLz7eq3SN+oh/LeDxq8DXzj1d3IhB3Ngw1+Dr9tnOAMWpkuS2CMAl
CwXe1yiB4yw2dLNgfuY+zd5BIjLmaDeFj2xsRwkb8Ri226tWqgzBoaTLDgrw
ScDMtdwIVtZ4RwOJR7iSpi95nMdK7ZRPjNaRJP6kzUv5sU6oxb+M93lQW001
FVM87aSdoehJzYpjsWzNhGwtkX9jDqCF4sl9P3xZLr3DNOkHGvXtWX6oceRJ
xP8vfTn67PU33loFwSK3WpL47cNgPdHZoAdlzo4CSFt23MHJNIXAm+/wOVPz
VIguYWAsmb+Lkcls4PNJvNguX+jnytB5GWAO/V17j2NPkvNPuE1b0Jj8e9wP
L2O75irHz+g76gfj9Wngb8HQZhxAJq/o2FhIwICQDrrUAhh7g/ETdEn5b1GD
m5L8bNXbIlxI81JD2THN04V0mvsjD2uQQu2SWtva82mrWWWysHl+QtR2u1wK
nftxlJfd/QTq9Vv73fK0UVm2RGJXcBnP/J4v8WRpUJ65fBMej7ORfsJMiHUT
icPBfmQ747vVNRZ/KzzSv0wpYlyHeWUkf3ZJ6AR+bV6DmN7y/9lc0e1Nj2tb
IDvPgfMAcHJvshqaJaX+b497M0GdghhJMVFL4tEte0xuO0sopSc5al3A8UoM
v2t6QkZ6PQVY4NMJX7Vv2LpFR/rqqHBEjRyB/pPeDbCC1n9oYEpb8nP/1oSX
tAaZ9/zoLrCtWIG+2IueJ0C06KviOx2p51i/Oz6Q8C2X2C+7vRwTKjJKygMA
k9N9/9quQLE8B0Q4DD336yuoBR+lWpB+SaJbg/4wZ4VBsW9yha8VxdM7v0YQ
NFvW1RgOdg3/4Z3SRea0yVD4myyFiX7ei5YS09TbEMA9j2uW2+ZHRaNdDxDE
GkT50t8qlf/XzMdhd9DAot+F1dlRDALCvNZPF4FgF4gLAH8GO6DzGKA0Ay6x
bew/9ipNzULvkJ0RBgLFfQN2zQDavTm8Rb2fkPVJh6UC1+7mpivvfZDUk0cr
uCJHcF0we51C/ZNA40mQ5jc+GqmMJmNBKIcRiI3nEA7NqMRAR1YrHuQUXoF4
i/v2NVg1bN3KXKx+Ygb6KV6MZWB065B2WotLV9Dg5rxLgaJ4e1AJjc4meYfp
FkYgiA3jmWawpuyaJb0sC7oHnYcY8DrwpcXcmvW+8jJkFj1hhxLfEuOSszY2
6GwEdGkNFzlOKNooarDrxT5cksnnaH5nXx9mPq6rJSpq6YEH/M8zz9Afuwaa
GMqZ4JMuKzjE34qvtHHUstvUiEu1DmtKFiwCooOA3FJ0FWz3hpHihTRy+Qz/
pCXuoctAkz0KpPl3zyyOBqiiycKHqwJxMYqdANWJ6bynwq16OjSZCa2n64d1
+oVYKX4sbFeS2EVE8G38uQgcpBqQ5nf84GB0Za0xFL285zq2shEOSmxfGL2V
UWDZBwygwFwcq5/mCt0IFjCjoRdJMwcb25DP558N/vjRUMmvqdfYdO5HyibE
T75hqdIA7ulM+m6hkBFZrkIZ5dfaH2jJjZ0kFENswJpVUpSJ1NxnA/zu0O67
CtXoW6pyXfNQv06jiWVUNeoHQygp+kNqCljl8JaZWK3mcBO4RMm+PJYIzBY7
DFFcWgwjYJwV+OuQDHXcuAc0lIojePcPDb3RnDEVgzhAyBgl26dCOWypuSRN
SE+ustgQ6HuYDdreqiSlAo54NcDN4bbyQYqlKjO5EIr97EdrXhbhJQORmaKq
7+ORZehdaG8sTfgyaV3BeAeGHSXKz+A96VzvLuHWhN8/n3RnDSBX76mnpZkZ
y1GGj34qbu1E/Q0I+J+nqnJ3gQ4oNm+2gLFPUbwSh9zFmECYXpAhmDhHa9AY
z2LNf6ydjJJmLct94bhqCvv53Sl25HbFv0VspZx14q5CmumY3NtFrSrbuYxt
1uj2mSHPRZZyM5jPk8BD2vb0G5LtUXPo9Bq/TjeRaxHQrasW9FqsvU6Wzfzs
Aw/U6kTrWP+dWShbxVLrXdtDLcBZBPkzu5VCAiodkeRzBvLOAdm0I0rgfOyQ
O8wu3bLNMXQtsQwjQpjjddQ24yLbafsvxMWmx+wZ5JPr3A8ZsemsFfcRyJUb
+tXWO7X7pND65CxuFghjdxLaihCmkyJB7BLz1o+ohw56tw+mOtwSKKiV5QVr
pY286uc34r30hOO8cGyA1qPUlAKbs3uN2MN5QmrzvzBRiyU554udeuC4garl
p+/7UdLr98El1wocQ+xeUnZ1X+lxhez5jTOQNUvsnVsg/jeppR9f2ZBEb8bM
di6nUKlQdWJBbuo4M6muwPctKarXdWx4irbqCk0zDYaPV/OgDsqGKkdnMx0T
xYUtSB1r+qDG0FSBbO+cuGXLnf1uYLu3Wa7mOSB5L3EO30lE2XckpKWqJuDJ
LSsE+RmGW2Op5OZsWj7ouUE/fPX2lVrUJevYKhXgpdhnwyP/l1n5Jhwb05Lw
iNN7jBbpwqdAhOFyGDCNUqQK3MVF0wolOXoel6PyeQKHSoCtZw8A7+drzYl5
AK4/yy/pgUPdIk3vTxQRwX5XypdW4BfudgEe8+fcpv+vR1IpYLARSrpgijll
ao72bW1q8sN0cgDr1RzfsO4vCGP+j6aJ5AEq98v5LtDIVz4e8trUuBCakcNK
7PNItLBxNXr7nicbMSzzrsZSkCG/+ZoXZlPUTqmBlVAerq9EQ/UGV2sAOV9W
ieqqtHbrwenNDxylcjBokaJDjijd4p+8J9guXGLkwKZ5AYTzcMgOary7WYJF
f7fwnufRPI6G6GhCtxYfZJODnVJgXZ1U4t3o7nmReFloN8nZYr0wAO19DVYZ
HlzrbFfv4CVsEW2di9Ddrzeg6MkSTskgJPspDAoegMafzZMbyWw5+GVVd+50
jgfILfsEq/90MGXCTWmHZMb0FJE9X3dZK6bNCJSPgs3Ms88OA60E0alBX5Qu
uLokbAx0E7xb9v6hbhmdvTZQ2wyP+AATKHm82iznARSzolBioSFmXQY0leoK
6XOGVH1JZkq97jGk1EZP/IL6id2FpaiFFqpmSSHyoLLksL2NVRk7JLI6+7Tm
g0bAAlIqqWSNxEBflX2PdV0cCjWymjwuYZmyRutYZ6sAytF0sLAwUZYtYtLc
rFmG4ACnVd4bMTEJwjhVPkbDHASgos3I3Cz8lAkPDLNhB1etBkQ1AusDSYbd
TgLDEGinEBTl78VJXUcGPD8VmlodUqxdjNNZMkXVQ6fHe6REVtkCXHFXzHm+
+E00h+viFvYNz5vYce/hJawcZ0OU+F09isK77bw221rBnFx30krDmTOF7r/D
uCYmzcxLlhRfUzGZMiPD4R1KYt9erSE/MbRA5AHrm2/aBwjSBCeWo5Wd0KhF
zTV30kauzpg+5wGNcXLZ9sg2ZU+DgKV79sKYWFm9Nm70RbOIcbYwe0ox1UMj
/9b/VDLdHB3kPZ8uO0MYRjh3vgAg9UXfMGLCl0fVkFdxRLQPpjoTz/WIKIdo
mGuQ4LdWEEEJjB3Ve4P4mbsBwFgtPZFwqFHaX41ItY5b/AKjjqAizfubEO71
TSTJtnv8zM3A8qCiGajdHp7W+zs5AYvpYzuXVnV+4QfiKxuEdL1CdecQK71H
p6XymNehc6HVjk7mWaXcUFkAsfG5r+VkG9ym1t5AeBr2NuUg+VToCR7O1rWG
7Ur5VYtDcWQbJ0oqKW+BU2gKSfYWGLY8iLgyVfFzcXz7qtchurQFP1EAe44v
H28bEmbsxhefZHw1zvmUc5RwRI1/Qyu7Img64Obo0uZhOXvcFnVgDAvKPJP5
iZauK8fbY1Pm66YJhq0knBJDSSiyBWDCTjpVXm4vR8l5UCd3AjPjW3FgpGUv
Su2QPOyUbL6IRCnjG+yHBF617NcZaWu4rwpKk4oheo+7ff2Qlsyok9tsNysK
lG/dGvys0+2ASa7cKoJfB3pFdneF+PjoRle1JTl+8Lp+wms2VehUczj/YUmk
wmDLabWLqXjN50nP3ASgVjJUTw+/n6T/oEYre4PfKyEj1VOSCwkFobB+2kCI
u4l7LVq2CI5TzZzArcH/55OjhueIgx2fgPKVKpdgC1+LTTayXZ89GGLtfIlN
H8wYo14DbIV9t2Ohn3cjjLXEPaOQwmupL+HnPHsMX4fjnwkIfKHCxVcJe8MS
j/gXRVzQVW5Fxv9Uj4ArLDzHpv/2C3myweJFYkkbnIVkHVAoJd8WlSy+p0TT
4klhKJf8JJE4wXkAqQcfkIe9VGOheWL+MQ0ub70q+CXKiXjlxx1F9twAbf7K
wDyOlnkmd8CrgKIj77affZluvO1huab19fTKJrddcUXokAnzVuXixwXqgGpT
gew4+TFeQZId6BxbCSf3FxR5eWg7/6UzdLJJyGESL3VMS9y71vWqentiqSal
Mc0cyF5ArOlbrJVD1U27Mbme8Tfs5RepO/6F1GfgYT7NjI90x2hJ68TuWPNl
QQobWENlk7zp6sD313b3nwl6x+yPRIFRFUyusLZ54NEnyvLWXOR6aIDgzkOo
B63HMFYUCRpgR/dinAAYihStP477N/6+QkzBGaXI7X18//eo/DLrGJjZuCt+
ao9i0d4xWDlo+J7Y0NRN/Ur3rR+jBXol7EoQuMQcqNH6i/vYydw+TYWaYlrG
SbFZX464DDqzfyk98wxYyIC0kflyRocMW1n4KqjfpklYVdgIF2/OVidKJz7w
+Wpu7t071mmMjHOnqZ839kIYa73Cr3J5Tn3qHj4jFmJvOkePU6TTQIj2sg8L
4wG+M6DfTtSaTEIbYJ79jPpe+xLtZ5z+F77sWmFNCH/tbOa9IFeoLSuMHx+4
XkD9cx2+myLX+9Eb2r9qfKfw5vzbmNvdmkkv7/TnPg3NsSIPK9B3fLe9UVFm
uq9zJY78j/4hkmREo1m2HtnACZkmjcmU8n/kSA5S8dz1WE6i/EiuAnCvm8vQ
sBIrQibdrKJppMgYn8FkWZp/ldRZNG4CHSE1WI9YDBd/VWTDiCs3thYlw87n
7paqBoxVIbWa32nhEiYxTa7kXJp/nNtqWzSHuM/NAbG2QIGiVBylKH8fRF8u
7vf8d8pfMcNhJmiEL5XdNo0mWzpnDvVWxkubnCNYWdIaODp8TAsXvRqtQxie
ULEQjJ+DWUdVm4kPeRguja9WNDRk8VELaUOvqmaZm0LW8yp+0nM7K5OhYUsV
LnL3GpRhgDXG70FKCy/ZefwJ2+4+nqb+qRzTA5a/jD1rjxLl00BeHBMe1xcP
DkFCM15c+2g1kRgp1XpgeyUye+SqGuVElG6iRZUXJszZneSF6AWO/WTmNNPW
mdO0HVOTH+BBgGwRa4zfPtyXPqRmDX+8/ydyETZmHMpmFrObmj8/0Eg0J/+P
ItkZwyvcr6jrc22oE1GDfTXEWvAkZfRXyR2T/tDGxVJaHMKdR9qJL8WhCsw+
UMSqb10Uy2aqKzrrzVK6Fn4nmZJVb8PtHE1NaywNGU/hzCOO+nW1GAPsAEEn
cKqQjkM/E7bKqqwDyl8IVXSgA8hvzpNK7qXSErKtS+ho6BwAAodGEnSnfXNB
oTWlSaOsw1k9dqRmwNxODuR15jRmy7QGalGjfcnFepnokY9G70yo87avpkGh
j+9vfKa0zeeHxCsjgLuwobvgMKzSUD/3WXap5AKOQ2ZXr8nFjWLKVj/ebuuN
KporpNGswcVG7Ofm0OVmc/kVeiFJPKVYdcY4RKQJuI8EcRnjrT++AS2cvA/P
pbpCoxc8vBqOh2xDhhByuKHhKE1LKwVk+ym8NGeISQPvlS5CU4uMzFoa5FWL
c7f9x1hiq6JpTFa+3GHCjG2RVcW89UAU0Sq6Ej0YOhx6CSVCA5dxH63I1fd0
+zOuKuG8Ijrx/hnyiLO64brILapYR80sQN1ENKBfLooo47361LJyBAZZeYmO
pioGjzalNWR4LrK4VdAtmNucwDYOGoBy8iEbKNmPLJtA5y+ZXMCBD3UVlCU+
g5przqa4cjDDmiawZhDzeEV8WgWLr9RpHjTTg+/g1BqSQa7I/ipPzVsfPVMc
knYthk+F9PX+ojXxs7gArWwTT0zzl0hNg8GragJGaDEQyot8R+AHRfxHFrEd
uRWTJmlUqke5+jIk8ALKTeVR/TZdlzW0SuIfAwuWYxLR2HA6z3XCcqGZZyNv
mNalrneiVTIGcQn+ntv9jhGgoEs2eFA9Jk8uryR4rT8ScWtPtuilqdb/U+Af
Kda94BHWSiUSt4sj6g7XHwfZXVtXwsuelGyF1KKjLRYeAS9JdrmU/ahQmbsA
KApz96TIbHYU2CZcHLcUIBGhia5jhdt/TpzSoSC3fwVc/qYOo2mVCQu7uBC6
zy+mEMHyyBOSqROlDbNQngjHlWrWnFod5f5E3HY7MvAhW4sw67zhYes3MnAf
l9+4o5y5JeFK+C4tSD0N6FpuEtyV6hve3QUjDG5jxFgM++jEdPdBX/J08FZS
3txsgz07je7V2Q6Jfx0VgfHk/GTO/ytnWDJHLcbBPHYA1qDjGSAAshIc50JY
8Nps2y1ehhZ5tXm3Ey64trqNXIkab2TV04W1uFukdzYhOzz3xseghF30GdqX
VlYkINcwNz58oa0C8UE8q1pkpOOzUY+XxY7j4dvPc4B3KzfbVK2YfkY+qH/w
mTMjA1bAeBkey/Xj2Dg4hcE7iEhamEyEdM/p2RDCyeCJOEb+A3eOs4WKHsf/
cdVkPNcaBEKEusN4hzdKuLQXfkK86KJuxd8UnSmZOkrdh01SHjXc1h/CM6Eo
sLjAu01NLX6ceTDApZ0wf4+w9lFHfZbX/Ei5bIXRNXqEqGuWjg6fD1U2dPb8
rbsT5jkkOcrfDWgYQ68EIviPcC1JqjRxsz8X8i9plN/9EJxkcHKE6XAJULqg
6We6b8WTP46s9lVk/Dz9+Fy8jv1+lV88d5NVfk/AmqMPkcW2cImocsfjoIsU
hlC8vvr0jc4p1y8TmnR5vBczZEd6Gbg6qvllIRAUIVLTaprHkRpPwWILDAy5
+D6CKW5XlVxKW8TK0qLw9R8QmGVLjptlo8EaMXp2qmkEx+DQxVR+c4ypXthl
uOhXDNoMLXq1sYr0zGggzepA44UJWFQqmmPqq0km0+YUbOFef1QVwtVHiKfX
pK12db4Eqh4ktn6B1jC6jagkkn3mZKdzwTIKJyrUmJruxwSyITZ+yLMPeam1
SkVZnrovwQcrTAI1UTxPks8aH/4w3kNBk5N9PoO+Pn1rdiQfhfxYzqhIkfSh
Ftv5VCcNG642vD+h5RRCKDJ9lUCB5gF6XdW5dkkIgnaKB5Q9VEsiO3LfvJZg
i8AxKQXRSUOXNsR2qgPPq3p8kPvvcLy/PaoLVz4GbKXlFooQHvGF2iCemZeJ
sNE3FVA11L0rItNpE6exrBhcHn62R3zxcMiSymuO+YCmMOw+4Ih+QooYDuKF
4A/u0K/x1bnH0n+kTux47MM78F7gGs5SxN7TKy2nmI8dL+tzK7BL9RcYhRLO
j+yV/6S1iWMVbtk7coB2rt6aUi8+QFxifCP4kz3Piw1A+4PxKQz8fyG4rFEU
Z0BOA6rAWyX0a5vG9O7h9el3Cyl+X7pI1JdfJXw6j9LO5Oy2Y5O4Qae1nVNR
KNMxEKsbis5vz98LKQMEDWbkKNyh57utuEpnEOKRi1nBCmqSjs79/XltfzdZ
3owLEQ527CrgOpPbSjeR7ou7UgR1Dwtv1oXh44KQ7E3qhrUvlQ2PxyYlenNv
/3ZdTsNa4kh0uV4+IJfvYCLNcBGSSCEgsbwI0zlwaSkTGGLS9I6b7beqy/2j
V8cEJuj0I2rrolo8dlbUYnRHgsWH4tLiiWLdgvxNpgjaNQJt3u9EpB3q8jqM
hh5qadgP6iHcC2Fa1YrvgGmzIrWsS/xg9P2jsGGhmq5BfrvGh+UQYCmJ9Od2
4tzx9vf6HsF5mgtZjugS3TGceM+7cauA1oSGNjzRaWsCFxJqMltyDKP1Dmiq
ZAhS/EfszhRY+RddFMK/Br8ACWeuwl9njtMy/Ss2lVtpE9/zyMv4NjJzyM9a
upzvW3xTaVrcmTnubScd6qfvFkmsDhF8tWYyNrgQX8lu1kioWbj+yhXie4i8
4n5Gno3Ol69nwyTu+9yqAqpcp3Lj0C8OnKoTxnTRlEEmzv9+/sqkpjaOprzZ
ZZ8hcxnBKXVC7zColQUqTcSvDpaGTqefxGAE5EqLXPNtOUITzdJ7162NUAJA
ccfSCrEt4btsG1EApZfcYBBK5HTB142SuaivsAq22XPTaKZr/IbRVV+urTAS
rnGG819lefkMAUcm3hr1N+QEHeMOt/ZLi3peRauIC0+rWpANlOHa5b4HsGwJ
ukJiDwi0V6mu22pbWtVn6KjFplvUba+zOg00NmPuwWn3lNDUBnakcK5IPwqO
/CgM/MXBmVh0t2LmumnpUpoOnXBY2kb7Q0dMOxy0EH6wmLiiGe4Vp/6aUciD
ZUKUDyrZkDwQ7+SUOmcSy8FPMf6ZVWsaYH3a+FMHge+k2InDhwfQL6uN2CUo
HiK96iTD9YL3PkdW8crJsQBIYTs9SRDRAZNffC8hZcn6YQf5+pIlOBbA9r4M
CbzyOVAGS6koOasbZmzYXHoUG2tiA7UTOckprJAkw2HCshWd3iFBFtAieNyk
VtF/kNqgnKm2h9B3INYiadZ9iFX2vJF1Ue37wzsAdyVgWycNuyFB93lHFFJa
tD1+I6X9wlRKkLTGz9cEfA5FqC0hdSBr7udAy3T3zyu5fxP7gPI1zxiibRr5
A2L1e2Q8Kp+nDotpxrngoQcaYG0HRAN5GwEUhtdvo1bjMVh6ilIEJzPcIb5h
0DMvY4I0BAAbXooudThamm7z0EOwVS9bfEY06G5dfw+r3Es3a/STPADI+zIL
AHzFegSXYaGrVlRT8LXNwDFmvI98hmZdrVpalfDXpjdR38iQQhLc6Bin0n/6
anoGYfdSrl6pnskuLi3shoT9EI829niqfs5pd5a2Rv87Pb6bhBm65uK2YKBM
slxcL9t6ugORAuXLU0BSFuZXmj/z/xpJJrVF3omaZeX0D7l12AJdyD62dKNH
xJJS4NVVFGssXkHkVp7zWPLsxoaqg7NHtmZXhrYUeItJHWz8O9sRNXESfLKV
6BwNXyW1nnujJbA7m6xSCaVhqLnF7faNYdV6KlMC+145uxzqBexFM5bZAocW
mA+JuIcSGi7ODhI99noUvu0OKEpDwq1ESZUHi4XTNoevBRfAZvuzmo3+xyoL
EyAo3TxOtxZ4whG3cZbwHSN7w+s+qgGGohA/aVzN7sEdoNU5PdzUjccO8c8w
2iFxQOZO7OCQoXDJTvAQIMijycSKEVncuWIBf+SgUOA9X9HawJZYy38jB+yZ
Ar456w7EkSX7F6oBWTOWgyoEjE7zDl2c3PXFgXSwogNkZMjaaRHa4we55VDd
Zmupn1/snLi/tDBZAzBp35EpUiATk0m9KQv/ewzU0C65LIsPz4N/MqMLJZCS
u6V+mO1rvm0YOJ7A+p6ypqJ67GdlSHg6eKHQ+yp60ZXm9j9bYjpOuU2LHY1W
pkOuCkj+EFcvwnY5HGTE/S03ommVEBkO4p1wlCUa3WgekhyDn8pYE/xKgdfv
wMepaTqvo0VLPYH4/HDMViUBiAgKzmUQPSTsvkdStLYkkoyLGT0BMWpOAB/d
ZIcgjPCOAvajjK9MCrWXOaZW8AfHbXYGDI8eTxJAMCNcMIkJeSFciASBbmnm
SmjkyB7+nG1zVt87szxHwdz0a+InQKW7X57Wblfs4o+QPwb4U6qLJbC88Dca
AqxF0yvCXPpB1eEUsw2XXFoDIg3wf1t8eIf/UIb9fAeuEzcu3GhccJz8iQjt
NZWhKLE2JvAsff3xJBr4YXBezJOzM38AVwy6xyvXeNI2U3f6xaTYt/pdS5bw
uF3GuaIpm18qpgdExJ/2GGyeav19aNocv9+2Ri0Fgr3FqslHvkBCaqz7HENH
hWKSgqhVChhrA3fzFG7lWhVpRpuW/kGer+Bb2hhPO9DkGgU/61krk6Ae47RZ
JTdiEjFmeD/wNd4crpQzi7jOrXYxc8DdHnGB2F9+q3oAPNoI3FfV7Xg57v6e
6SlnHmFgM4SuJ/NkQe8qFuY0MnT1m1NPwkyMd8bouvw8ctfaCV5/MZa7ETXP
O8k9Tbw+KF46jdpcwwuXIm7BxFPzBwRREX/shjHXhMa7seNnasuDI2fZ3lwN
ECIQPOnvkaYINNwfbj8vy8rVXBSAcVPkwsKF6UMlm7t5GzukcF0/TFy8mJnd
xdb6v4Y5eRYiWXW46v8GPrvq9vZUvepLpRBcwlkmrj2DiIXQXu79inLvIOgN
5fHOiH3+Mz4eCr2OC0RvcLRZ8L/K5KNMuJwSUo0fcoXRvn6sDdU6ag4ugcyA
dtrjGJSvxQpq9BTBln2YWPjl2IkkCfpm52TRUUG0Q+h7GiE8gdGuLYDupzrN
Nn7iJqfWgUWWPo3xQzgte6ZeJpRHdCsRHVY5s9UvixEVBb+/WyVoLWdgEAGt
wQIYgmIT2DtVjULYDOdHhWw+9Swdzqm35hIVL15F0TGedX1w3dhCeoGTJxKI
KIIsVySmwcvPd0hvcp/Ycjs3zBekezTALyNhYXhsY2Aeain+z3VGurtMQIuD
fXdPk98s6ueq5VvZwaj/Vt4kxokIwnhAdifxi6QxX60xhrztEUG/+DY7bLUw
tIeDq0UtT1pVz2+tVMpBHiNALPfGgiSp5LBYUKrNbUGvucVloRBUryPe1o6M
fbZqYyqIXzyV1z/YX0v8++YyD512nPvWb3nlgagdV6xc9BYRkSFpFUyMJSNj
Ips20pqP4z43cPxfVpRZZRfZDRQLlXtZuGx+kPxp5ZqQW77feS5J5f5A2gHI
zaHMRb+q/Lti+noieme5rPCwTJamSUFzU0nJbxMG9Ehow5bOC1dV7RgsKNvq
lQtdGymJsHyrslgxYu2ulhFhvfJDnoOC8J1YeYphsWBhhZUuWwInHogMzwxf
R1KwPTM7+s4bL/Ol6EevwHykZ7IeCTqDqtqYpDNbSVfn3SDKXfnjiksqxcRC
i+8sA/clPDIVKX5Y8a2WR4ormQdNeE0gylN3KMcy6Ypb+wa7CGf9JlD6/1wd
CvPa+3rP9T0bXoTHUPZHB03UgUIq3I287GmZrkrgHyyh3NVKzn0CFXqSvCIO
u9LVNHGvz1JRmN4y2VwbCtAGmd+5rmBTkN9Ixj1+hoaVaUVqE8D3kF9dXPBh
DJCfh5RZNv9K/6Tz4Ha1yWsuTNcHrM/oCiZnVcDESe2By8ZHSHxp26vimatR
8lsEt7WUWT9Kc0cq9JzOCGpDeqz84Be0f38d1Z9MhucV/GDGeocB6Fwmw+Gl
+9T7y80xnz9M85mwXHw1ULL/F3ZN4yB1DEXjaCjEAhiy136aeq2xImoFxnh+
YElQ2QuWzbtCilOmknZ6WnxyM1ClCvCxxIc1dllxhmNFaNjNsK9BMry2huzu
13NgPcrdMmEXA1mQ09yh8j4A2Lj/ANFagIOAWJ7XdH6Pd0bEvM05zSvctf1J
8myj1uu/cythW7MKJRVcuu9sgBEvTSYyMrZTw6kMAK/wQr/dqm9Ucq8sX5b+
YY0Hrie2Z1xxq/1uWjsJX+KQs7dOU+QBut4UHfkDg7UjeVT5WpvXAn16T/9W
p4Iy2PUs4c6x2258lF2dRJY0OOnh4qKwEmubFiVnA9F460Y1NZw2gqXDmnNp
N3nvf4W2ntiF8IJAT55jJ5oFynbRnr/RWSzAEfgwitKd2mSamZzlzpolwQEg
crHYa8KgMBPf7zDFljPJ4JEGYaRUMoWeJ36LGhXs0FJbx3Brp7BaJwDkg3Wq
s66IXpjcnp9kYhKRa5q6spc/HQZdn9uqnjYaPVqdIzIMhjqyeHlZRz+GjWz/
wUjS8wvI/4mNSd8FilJljNsaz9P7FZumpuICQ9LlfiZ1cmU4t+lK6j7JBqUL
RD1aAPmC7wrydOHrKu5K+7byMWZeg5+RC7bOj64wAkJSI4q1uE41Ff89ISnz
Slm7ikZ8rq/r7ASSQ/eSs42ETNtaDK6E1Vmp81e0lbyAV33LClE2YOoMMH5+
6mz95hYMc5S/eM6HIcSNQtRPDQvynGwpG5Cbv09MEGg7qzxfYQqUwvN6OVzH
b8JODeQpMXrmuF/kEVMwj5G3IZ4uz3E+AeZHpNadgmdAiZE+9rtZmjktSIp+
drYGXWTZ29GSETOOdIZl88xF/uX2HZ2VA6BKveWK50tDJCqU2ymujoagYisC
60CjyaAnil2OyDVQOMEraU6XIvXnTSWUbwQW77vhyOTcAPOjWqJFVjuCZzZO
lRQmNlR0PxygB5jGopUQfi0HUXBU0P4bNSab2dzgfai8cLwkgm/6J9KGIJmk
P+eqr5cJzi4piVuI7A3LSTxdZzEnh7RES1kcn6MbgDL+3YQScRou4sR6hvV5
4Ouc4TwVT5Zvcv5HISa2DuTeS/lUbKmcntX1lb/QaR7crIsJotq7itKhUpTz
iYunjW/zL5WSn33kkCiErSf6ZKkSbeNdEipfwnRzcDf8hf2Bw35IH4GEwvga
8pRWnIpYeIzncjv2Befh27LTM1EMXQSaPBtWIYZjegCCki3z6OTr0qtlS1hz
nqr3st50CQzKoNfbaj1nonIANQVXcymeS0KpVRJLOMN2hY5y+KlN+Kb7QW95
Ak2FWc0dv81O35erwOEvnjYCWKc2Uk1+vMhatUM2VmrZFvWYb8CqAxORPpl/
HMQEm/MgeZV6Nu6y7UKLkLyeU5RSuLfh/jaa0oGFQECj9RCTPa/UWLG1kPrf
1e2LClKqtV6yfGP0wEKPCHRy3C85h1lpizI/eu4+4vIoKUWlWpxqT8EfpJ9I
15xBoV0m7a6K1N2CAJittLmQaVrmvXeCbYKyP9U5QsXKvaaizilIpb04l9yw
eld9atkOJvda2p/gmdCNrgqLYWsyAcAipDcRxT+iz6D1b43WZgn88Mr52a8v
qkgShe+b7z/Xudt4BfSsDhQNlKf+hVAPSwdD7GtFv8ScDHoGxpOim76zTaIY
qMgNUcWsUWTwIGh83WRgzwylX8doDHK6rptK/sTa9Lne0O5SD1w1BacXu32R
TnTCfEa6a9TAm3sRrwykrqHYyjSsWTiMs70+8iHk33pbueyGCjLsO4RkmTD+
mgSYtKAghVsKUSC+5QjrWHXkG9eTL52VaFchkqljtMOzUAsDCDsgtH9+bN4D
mepwcv8BTTFebO7iumhbMGyaIvM2rIvTB5dC9e3h4UvioOLS2zkZRY/X1bbM
OLQZq9b0aFuvAOHaZdrWxaMW9lBJFamGlY8MMgV/FLNo2O8cWAxG/xTrTB4l
/jiDyviP57LrFzdXtGrKnZK93wZr8CZdgN8xcGX5/1Gz1FC4jzBc0F4dRPOU
IiVLRUYrWIAFGog9fCu9fz2lhZOMGRsjbONDU8DLu+a/mOl04pIXfeE3Wip6
FMhNnyJV9ycZiS75R55Sn0KdeRpDllEPpiGhDCl0HlF74odJeCVKGMMfkRvy
BeaWn4f39/7NgGZs4OSetTnSjJzHysJLWUmfXQ/Dc+/l/ROKVBmmIbnl9jSR
Dt1UnXzfE4OULUPi/Qz6EQ+N7SpPs0FP806DcpcAQPw6FnfJ21gQDK3FXVai
6OKYuSNA7dJ9LtopTLkZoaV1KoAnBp4qi+tXHfNAr/EZQ6qF+GJfzQJRtw4e
T/dQrrE4T0Vd1IEWW0e9wfJeywFAUHsAEjyc4XZUgRyqJ5z6br2o7bJOsra1
Q041ms7fUxsYRbxrPqf4Vihv/SNd+LZMd8h0PZvAsPD5NbPGlXzoIJ8MlkqI
qgpewbHRUj/xvrAFvLu6YV0/5FyThV+dYOhLrkXzJ3N95jgFUegmPEbld+m1
+FdyLF9UVyL3nu/R++ojN/k9uLxKZ7+DaMx+YkvCB9tJL7ABHUw4f/5b3B7c
llsWhjf5Cx+G0O9oxGOSLIVSYMQy7y+MXTrf+eCYMcGtqp4FCc20ZKjROnuX
G60Lw4OhSWBwsxn3VhRxoPgYu+PZ6Rf6AkzQKvSkpfutWlXmVlY7xSrzlLhG
AjA0yVSrt044DSsvdksWqLnayLbXRP0+uhN3QutNIfY4mJo5I+ZyhzlVK5wP
KOXgFVJS685EzXzY3LIGcw6UAXk1vTO9RrG33QZXky2U/x4h6nPm9sHB7fyr
ApD2dJQj+BUxjPyREtYS2EQb9MK9wIMr6Hmgqm0n6gpCb9jDx29EUZJTaA4L
Y6eKCs+EDxqMfeFtWmp4DLwg8fV5bj0QTgBJ4/r2/dqL+cL83LdiRTNG2DX+
goK5rwNh4zvM0ZjIHO3qKXrl/ZwDpXg3sEAbFSQgcaFCGQ0BMGE46KYwMMQc
WIahq5BTbZ1JA51pw//Zq0sFqJxA0VbxF8F93YZ+Wx8vMSPr9QKZ50g71b/V
5T07vDv3ds8+JiG5c1lNBGyc0vlTes7OouUcMBZo5w3q7Gf1Vm4B30fgkIAa
vHfeYAsUYsVu1imCnB8WNO3mRZueHVO3qB7LgG4okSAVvUuFKGHF7EgEf0Zy
J743UL4up+WQN9IN7sPaAugZd6KGtbIIrihdd4RciswE4HfhDOzlqLM/QstX
DlSv9X+s5r8OmdJXe7FfKTpZANM9Na+Idziu6vntuYH6mtkVhjmGyK98gu82
kP/F/52LlMmzPPp2nS9jh4RUV0nCjIOeMcRkHeHcKeBSlMMB/eF6zD7qsL0R
9FS4dPXABcmInjHXwTlpt9050CwvDXdgC54uhTdy7+zrc9NMdJTCJBlfuG3+
/d11CSHRXk+cYvoiQT0u+sXW+9AMQ7R/t6lqCreUvIs8+kBbWVEyihDBLCRV
CN/QD4/RCd1b4Zo9svL9ScGfOsxSNhOpBbU114aS2Fxd2S+Y0ONfyEzunZ1D
KbrXavQ7QyCC89yp26q4/l4VYBWsMBdRtpAOh7OCbcOCIZIl8FmJbkuIhNvF
18VqLvv0nwIIsFVbWC2mlu8rrm/HqwdMShHni3MImgivjHf2HBSggNqBvE1a
kGz99mwbryro4JhIEBKwi5msrI50asW7Hklt8en85oGjUKT9Weutwx3u6bLd
wUpp1/g0LIAjYwau0RRSF6acySTlXS+ectYn6wMG5Qa5c+GciU5iNaRgRON+
Hc7eJzO2g2Vgncy7D681ZOeR1AlXIzHvZ6AQgvM2WGEzS4gyH+iPvHH9cF/3
KJokGR1xYgBObKK34aEgI63sLmdMi8mCb5iW+K6i6wZtZ8aXLngmi1gfNaCv
9glJ87HbEf57dJWWPk4R7aZUGdbeiKlrP+2JEJVjE68qTHJZtIcEXk1Uxy7a
6Dk90lPIyzHRN9E33VSAy6qomNQXhx374SImGBZUwxyutHz2XBSoMxzZ2JRC
SbPLCR1Q+F5WFatEfziSK31v4zPXs3qrU5Qu1VgLflWZRPgVI9EUpR4WEaaX
lsOVnyP4TW/iCqK/iY0tfZrTo00OFu08CI1RqfF9Q8P8VYXhzxW6l24xXCBA
mZu7fXMnpvCeUCd8mMwzID3p0K9t+SB5MtMr12+jg8S8q6zXf6Y/P71xWWpl
EsbmN54Hfdm8pcuvT1aB6Xq9ht9zzottdb9a8Yv+2VKbnrhw9kzpqh3UCgjP
budF1aW1c0mz/9EcXtSDHZ4LL6sPFj5IPwWE/variAxNAsfEkRzxXa0vWkMR
DShEZ+/6lWxW8egldd6K6C0j44veRWd3+mXx3rkxTkdkmPp5ja//1F1o6i1J
Qu3xTzvm/zBnzBV3oVXF8Q8u3xXAFRpMfUTsE8EyHNBNEqdoBK03SlhttZXt
oV6NCoa/xuFR/p6B74bnx+gtLOHgIKmT3JdKarll4WJiSBHkln1TRkCqxaom
Pp47d//ydIVSOD60kDEyplfRIwi6TVardTnCBJTEioC7VPiDqiqhr/e2QXHP
BQzBJzTdAJUyx2MejzbtghAc3QwyxRt1ApN/4OXmvKdm2xN7GxyIcm9YvDdb
UsLFWVcXtQk4lo5MXvwb+PiApDidw6lRhOV5SpeKrQmr/Kuv48C8fG6a51yw
YGTYB3eZkPPTNd6zd1bM2BZgEaMwgeINQHXgrzc2OgURCCe4W2LEz4MwQ9HH
k5RcoZkQjlfgQfxuTSJJMgfzZ871VHRwl5JAKAU+EGKNS7N2lwaM3wXjV5hJ
pBYvM8eiW57xDGZsbRbKwJky77w4pNZqADqqfkuntN0UzyOXUNwwiQHDw5Z5
L0zJ3gzZTF7zaiBaR1+PP2T3zdmfRHntc1eeVb8GMDwR3h49GHK/NfnpBvJX
h92JWZ1bH2AobGuDPRPxt2mHgRG6N/NcaoxHbpe0RU0qaavFo+w+Ze1fdqpT
Vb1xSAWZIfRRxOGQYugAPVHtjCsMKmfoez3S4PVoWxWxIGAbvFtSBX6aSQZb
bZW4NxOgc1WQfTZN20R+sCXkYud2OXLboL6h8A72gm7wErTMPzKg8mrna9nM
YvbXgrNJJBTBjx/YRPejTfY29KxCBIMgarhaeF/dPWq9aHX63maWUP2/ca8F
4fdEyDolRcCo7oLXCOZada4fEPCfuFb3qViojdmYpYmrhrW+i14wG15liAVx
tQ1nH9H5j/94dXRWwjJw2a5XgeC50Q7msm9JaykgrE8P0EMRQwV1xM/WwCqR
KzfQqv8iOGCVxvlNXilnm7HI2mrsaaEJMQAOSg/UZDdd+2pA4cqDgpk3FKmv
hAXzutAaLWruCji6nEnyJvV5Yeay9p89VlsZAA/Q+XmAh/euEK+8Cs/44A8p
UWqP3ukcOUzpLrOu5NvREFKGu+DlPTuKX4WBmLFCPv1fSko+JXz74sy2QBRX
JlThZxzodcSWwkb0wnydAebKrWXS6nihSMuhp9VG49KUM33OeL1M1whT5+Yc
99DraCpkp6FgizXPFZZj+h9AsS9DCpUa9WSt7JxpSF6r6LP8bvqZjR6WlsNb
B/U6KhHhMjK2yV9uE/VS5LhGDpkcWZjzrmxiTFHgfEj2/DX60PRx5qe9kIuJ
/sRR/SrvDfwSZmBvwjjC630tYl5WqHrenf3OPg1Yfe+4P1a1Z5KyT5S3Taio
wH/6PKg7foMy/mr1tZ88ig1mDbausi5RRkhsebT3M6ynoh4UwpVr2SgQPZEr
LLJ76Aw+gtUa73IcBX+O8RqLdpEYy0QQ828JN568XiBVHXboXXebDLxhITvU
OtEzUjzh7l+Chbl2eVKvSbD06oJeKhFEswxcEocmbmxqkma2HMzbSwLXa0t0
mtDxHICf4GpSun2IaQQT7RbEsB7DeWNuY9AJfqRFwWO8LOkfeuntxNn84wcn
l8CkPBf3Z7oPvjaaLIEX2Tmag3HrVsKo0MxkJ66UhWNTZ9MYl7sUsnVoXjr7
wxS/0vLHxWpkhHHTXUqKIlzvnJjRKAspOFA3Z+g83eS7EE/v0P6/6h2syk2T
nyRGhUykbTwuAg5OBfT9f1q+J3aSFkI48B40DCiAl8bWOEDq1w4AoG1tgdN/
FtiRyejBWIb4rCHT1IZpyqLVZQ+65BPVQyJoWqcPVOuoV33t78c5n0jHtagx
E74kyylS9lVlqgEWnME8gTNq3RpCF9ceOofqCd17ImyjiD6svChcs1fusvw4
T6rTyg76l1Ywq+uE7NdOhu73bcM/t0aUupY1wFQk88MS5gU2MFuLxZWlROCY
UPJwXvdcmnrd0EFPGaxIOfXwt1qeDI93YnYWbpmChVHk/wJID+2XQ5xJ69tZ
iJneHCnqHIRvDdhqY0rNokaFx4m4GA/S79q8SINNdstrXBCHw8uwLInXFLOo
+IEFT3rcsjw9Z9m9cClEnQF+LOHRR/xS4lAU5jGxNKAK1dB7nrLBmHJEoFAz
i9D+wwKqcuMXB9XTmNszVigyZ9rsGNvYyAGplLB0mQtS3AIT0RPn2SuablyL
ij/4NtKwoIhwo2Bd+7jN1h2cqWtkxDiNgYyePkcAZ6mdh6S/DJ4D0DASe6Nw
pOhUWwJ2aURTFzdRXl2ZfbaLTj2sRKqB2laJ8cdLiMbNgHgmF06L0y6TmeO1
bg9n48qKzS5ZQvUFaMCf05iXzt7mDfCQ8/qjBRYHNCFTvGBXEZjGwADKc5Ld
7+2tIcua4O9e3CHUEoyxEbaxiDhJM+p6l7ZM4C48i9Oo2HK0locPTY4uy+sc
TbBjQEzyudkm60IVCFgeJtw1nlcFCmPiBWR++kpN0ZIalmHdEy0vc7MvMWd/
7QBpt9i+QI0EVSd0+LNaBaJx3/Pt1vBFvgy91LHALqmdRWIQdk79qYIRJ1R5
w29WT/DrL5jWCxauuZvo1saqObrdXYHvba8wc4kozymw0txR8LHbfUL/swMS
TsSe8Xx8MyvFS4W3LQQQ3/CKeEb3Dr0X4xt2ryCRNjSiL96QU550Jd4ZjhFI
JrXqK+QBjyq3u7+KHlZauMuc6Q3hZ77cm7V+WfYdq1mDQU8QxTpkVwwP3qlh
406FFHllGyyQm2Q8wVEH8mFCAVz5F7fFjsV8wc6UP8sibbVlqSqxnPoQdIkn
pAlS0HiRe2sTkcxs6XLdn2tyfPERvPMc8PRU2XnIIFoC85pyW72O4VBCf7vB
2CswUVO+51SChbOrLMPCdHEIVCLOhFdLddAQqpOovZjpVC7jSCmdovRfMMvh
lqZv1nmbnaTcEklM1wbfGSFyvISTD4+am8IKWpqOHrSCiTS0ByqTZTyUMO5D
Ch0ugHVilxy6eG4ESjM+ORbSBxCtrSfWiDlH5ICaYr5K5jaZX8+vWEqwodbC
wRMIfcYW4nHts54G5RW3NpODTpEUk9osaA4jlWqUhNMoihVgV1qaE+5XWcgz
Lo2hXyj4d5fUfaWtCwWQQ0AmLqrGdBN+NOyOSjvGL2f3vH66pe3qvs4AD4HB
55KhP6R5ycag3gZSnTfU7UR+D23qQTBmJThHIj40ysETaqtsPLctrmkrajq2
7nRTkmmPyxCKbPO0hWO/kmbERKld5+2uJ9bs0l3AiLBEu6Jb3kU9RA+Lyf8h
jbLGiRZvY8tmj3EL0m9xvOrxY8tBwt2D7OMvCDBhT5XKZAMqpvxI/rYnwTyO
REhz3Q8YeZqKUxhBLGefLV1k7tyMxXwMt5EdF+yhPIr6rV19Tkl1zYGdrS7s
l02UYNFUrhFLPQDAtAxMNS7U2GBlILCCzClHxfCZCRbNG8OsYq9b9dObIshg
42srLTJL6cPFmUVCLFYDx50rziN8PWwN5VSdkSDCdrqqVSPDXHpg1HKSFnsa
DTKdip993iGWtOMHyKlNZmDPA98SJ1IVZMstaAwYWKfc16RpIO1gHfB7Wdaj
idHvojhwPlsNdQXwRE2A60IpfJFMocWYA7TQLQpjrUpG2suyGFFm7rdejSM5
R55EdiCHWsqLGsewNWzWFWpa3wc+uxCHU70KI8InSEpRBz9V70XddI3uXIOV
/gSVrRSZreeoqc2CDOGfG6FGQMtCoV2zh4a0LZWW9QkT70BFw0qrK+lX0L1z
DkNd4kr0Bn2a9MJIbnHQJt63hCpM9rapCmU+T87SZ/o+ryIQva/7gpOUAnP/
ivIFrwZOtPppASAEGj8DwcPNR6I8h/8lV0g01DtySzk6ptxD0IIlgG87d0bZ
iq6ZpcRv/VRS2XlSTGPfLAuT7IMIbscxx0gk3nHCYGUjq1TApAaxiOcmSaZw
9pVa9q8pKVO/ofkTtGHOCeQ21cYhyNVcMKtOgihTQM3m1t2Kt7jxUVFP5j/l
YTOOpZyars3EATuXsNOrHE0KSwrDUl5E22NQdx6t2T/mh2GxBpFPbgNGxnTX
NDXYITci/coxsZaMKAPdy2paVmNXoGjO+aWLxk4S9Bo6fod2uLXi8eCDgL0J
Ttv+huzdbxPE26nsS+ekaWnKlIEoVMU79MuqB+2aXH3fHO8ehP1tyDtEanYS
Q1tb5MHpTFb9lRa3BrAUKlnEUwZvlnfE2bRVo/O4CYGJvSFzod83BkJ+arMq
gUQ3HesGRCAofpT+S2salJHazGy8Hf2/2Q6GTYDzfikGto5uiMw8J/EnRvKD
DOiFgBMQd/5zb4uwnVoTzIaRQ/HSDRr5KZkYeOhlAtYkcxe7O1UniUgWl3Y3
U2csQOpzbT4yYtdtuutbliiseXrgq71fQoKBIQQ4vOYFxnb8yl9xFXd508RM
ZDyY+99Ae3Whyea3MXIDWrf/7JUDLjA6efXxWJ6yVkFFuAqZgQMq6HwQBBlf
yNelsMFhTMPlzg6F70NSuwxC+w1bWKeGx91/x2pn6op+Q2QnQcj2OWcVZjYY
LE1PBKo+GDDywsNBs8pVCuCE6+Kr9KK7c7uaUtMcabH1yxJxz0FFBFxGNA3r
KyC/W6lGmWGb59QeoerBF3O/nUoi5DM8nVpwsJ/XCu6YX9kHqOzCNnyB07y+
R+Ig9tghgh4X1zIMAjal+g0603nhbjF6noxLeGyuhtyOlbRvTYbYSQAFoe2X
Jvg9Obsi+nXgmxB1dfZXx6zN3PATG6e9vxsN0untrJdkKO6QvohUANcOEA8h
TRV7/4vOU0I955vWHHvThJEpzbAQOprQ7j2pEThUpnysvpwHRlaCtq36/zDa
xe01gN4iYXUUp/BIIeAnluGJp7Kz6kDEKmsoMAnj/CFN7Sk54JAciN7VMr01
z2nPo3KJHFF4+ij1QQw1/XMy6eKtRiOuCtJ02QTpqf9X3QwTSE3QmqAWV8pS
ZqOuIamOpkWWPJho0OlxFDd8MLkvRB/FMx90C+UftFeIsylXCMWGGfZ5WGfq
ZvD0sC+tldbc4oxvHqRED52sHxJn9hsoXt7V0XDXUq7dsDFy4yzsOMSvq3sc
Qp602IQhx5yWbLR7dGIeT4V3343UGEChopOiFJ1deu2fZMULzizuIK9uiZXR
ASGt2PTbwAofUNXbR5tHPNwbF5FWXCHI2vhtVUmfPTJgvTlax5XzjY8s7F54
VhSsNHmoBZujxg1hP8HDU/ZcSFXx1C0ukdwZql0z7FhlupPvvVHC7wMp9y8d
z3SuIZbRVej/Bj4IjOCNKEdTA4AJ5zJkDhyna0x0EOoUCzlLM9bSLK9IalHs
J/WlVKlFyHQmwdz7IAtedaGqvroLOJo+AoAvMGgAIGPGo7YW49m2W/JRxiXu
ipH8pYXey19VZ2WdUyytl4oKLzwROzI7Bb3PUt+AH9S5XgUnNHvYlDXzr18Z
nVVvICMJ68ex960uNGC/qhBQBLdU5pU+93h1Iwy26FuAG5e0FNtltdzfBuM/
+IB9mOafqr1GWtwjXj0F2eJMkoZZ/OxbyApyCp7HhIIf9Fl8jigsfU2zQMvg
Bx8oDiXu4T/2p/PG20skFES7HoSLxY5IGgwIOaZ8FAxYBr48Y/Styv3pnNt7
8+Sel64goMP/slryUfJOw6//x786JRrl1ZUQo22yuZsS4tMvFR0OXRQPK+zf
jro7Po/u4VdR+3eiyAnkQOzJbVurasIzoVY7YcFuZhJgKRzEkAR2nkBqIUNW
YuydE7En7/7hHMAPzr7JpKEn8AqA7HPegB+i0P2T8aeXBKbf8+siUuPu+clU
Po4dJKC8Vz7I9K+w8QCIlfxzJ4sbSXUh4OXCRfnpQSaRwDSrzOBCEtWPENOT
poaUE55Wdy0QoQE6X07Bs0yCqR2+i32FLh9YbaQglo2ez8kP73u8vQj66BXk
uekl/65vITe87AFm3A//amtN1qVia154vy7/y8wOpwXgNLJ81Mr3DFyG41Zn
FBr4R6uvSmwg5kUoBUfA6BRPdooeW8L3EaCb8ArZBwoqojCNdFzb7fDK8a8/
H66lqvgCLQg8JcdZRCWG3rz2THuGlCi1repLR2ztEyrXwGaemHs6i6kCFLLq
5asLphT416Rc4eF4RitA49ZViNf4zw7D5OPuXSm9B37/yzacC8vYVAj/bGff
de3LjY7yXNcX+3cN9LxSBcUPW7tmbMuaog2J5sHXe/Ox1WNzXt/xKwe3XxMK
rwd+7ckR2UmrlB6Cg7fwMVOqWI5sDD2nyIOCS2xmOW4w3viERwutb7zfsHpd
kNlAwkA8RtnFks5aTo6yyDnRcngz7Wek7u4RBRYWS5qUoA0FTPOWpcWn1gC3
Ze/TQ7Oy+RPrNmmCWMFuTACRoNtcWJvxsy12zCEFpiNH8fVOedqohtPfpReL
cs1lPclClWqn+gA4Y+HeFk6arcKnktrJrskaxHQlJ84J7HPsD0gxoVKXujPS
wcPFvGl8Lmof0+pXINA7pdAkwmRkl7AY3Iey0S5zGRWzY1ql8ozprnsO672C
JfatMQf2hFurUs/8PLGU3orMVt35BgTl4SwNDnNrWL99iKME4Zm9tDEWcDQa
6V0D/C84sQCTVvCwgONNIlf0BcMv1u9H/Dr02Iez4JWNw9QP4IacO5dB10NA
bTWA1wtdTnlkWlhr2hp0R679Prn8NdOylLJ1yQCWI5BLefd2F4wLYB44+4Is
uhM65hwwk5heOjKUMgZ1Y//VPoP5ot+hQall4oqV1PgsDWekri4uB8LlAfMT
eO5ysG9G+TYWC4QPEXKcQuoqaMdwdBeNC9TXLHhS5hkBjv0dnS/QaFmC4oqd
u5GYXpuZlJDS9zoewDxquRroJpXoATJn5bH+dXY47QU8e/r0VUOkm94cPV13
4SQ/pZUqeBjFM39AEfSDju9sv8cITVjfj4JCUSnQtgLqMikFYTu3OGpABiXk
KknHE7vWrBJfHI5kflIgW/ma+qgvt8phc3aLBmfvNUhKh+FKSYd/Ic23yeSa
527HI+XWqCrathmJI81vakABIpqhDr9K/EtVYwyttCjgYsxJto/HMUTdH76D
h3CcVlrhIo3r1r1G3y4CKeqdkAQsawmmGZ9EHiPser2eWUQNfIT48g1N+WZZ
xWqwR/Re4E4B+Q4xBsZcxGIBILHa1XWtdzDwPenAb9d+8BezpYSuZwedD6U2
itLfiQ70jvPI5wUm9OXoeELBd1Dpig5lbV9hb4USjHMlHr5hwgTxZm7Wxpp5
EaqORZ5szQuBF0H0c6GYMQzWVgiI1asH1CED/D9Dvv9hEjESsawkPGcGkmOk
P+fVTkp1lCuLFn7glmAu71MnXBz5zPfwUpfAhRMGy80WIyOecGqRuJUPq9+Y
gZ72jySE4Oxy69OSVOnDtWLTh6qlPG4FlePLVfbCRiPnwJhHDwYN4Gvwcu4i
Zi73GmGRJG5/3ASReq9wvLIgYp0alIL1UTOzLTvakPLwNFqOuCiM53FO0hQv
4pSLc+WglprBTWwcaKAoPRFiETW7WsRi6+TruSQ3bfUQ8tnv2N6IbZJA4jIy
vTKzE9mdoDbaCg1yZCrXrwDYdlbVz3NYAQebimqsmQt/tb+Rx20P53sTwoeh
bHWt0Fac3aapQQj0fwtcwZvH96yi59Ale1TjpWNGS9cl22U7kuKFPzEAX7EP
brjGzMIe6KrbG8bf/LX1sjq7aHejpLEJodC09PGnnwfmxVx2lDpQE3T7aMqF
fNzfTCk5EBpUwBsKYdk1iBfAb/sbKepNLWsGhRbALRcmF9EMWqRHtwaZgT+5
Nvx6k9LemQd5TrxsnUZqGsUHHQbZX12Y6kkQmKuOB/Tl0DhrOTDKPvaGvA5H
OX+eX5eX3e4D0xiPwes8zJtbkynrdbOL0/E3WYaESPfKTWwW5b0P17hXV2Zu
3cxsC4WPXGzmvOEXPbajfDQT4wBzkb/jc5qqPvsTap4Cwku2F3WpY2ahrEO4
+ZnAbb6eLGmTgipVxn/54yuremzgQCLV3mEtDts6tE2gvdV5/8v4l8N/5SS+
2KIscG+dUlSbZ+EEA4GHfvd8xBR+pxd5VbJUSDw6oo4lkn9biyt+ffU/CNe9
1NLPHyNQZ8EIY6/RsHLfYuH9kOdOqLCqes0SQ1oDMwTXU0w4vctyLGtEgSI1
/2GGM7/IvXP0d6dX8CpV+wa/KhrWJBS/J7c2FBarjNtyPjTxr01FxHnD22TP
qDKYTiczp9qWvcBHOTy0nC97nSJvloSlA6/JO1LNvKI9wUumqYVLRf/L4Ef0
T+1XtKBNpJNhMoe3CDPO9vuJqACRv/dN7ZjLrtl1JsXUlVAJv2DGay1QVaGI
DFdi6RuY8UFadA+x/gtHO5sgPtkE6I7tlSnHb9sclP8gI+W8IbKMKxsMyoPo
IdUJy4Re9BukNyjbnL7Qn/1Jt0KPF8qoeEGMVNDo4Cn0KRBqFfrglS8abBxW
UlOZvcd2+yuwLXMuu/3FVXSp/AedGQFDm9AXnOh2N/BqqZgZ42h4l2uQS22h
m3DFUUQOTV5KwW3uI3bN+3vG9k+Jl9vXMb6ri1VJ3qdev2EdPWy3p8kP/wF1
tYgXeKHN7tm/BxnosB7fRt/lRrdJaZF+E8ygxg3jeI+OFfPf+S85iqlBneo2
XaOrn25H+GhhsCMSIj9GiCv2arLNr7l4fWY/cM/bz0lqbM/DIiPROU8IRSAh
y5qtlgyCJaQ6WQTey3qEXnRuhZ5KRcCgv51G9n0X7Ww6xxsrEArX4uu+qI9Y
LT2DFGg2YHn1bvHb1HvVLLqIiyumEN6fi8x2zFee5Y2pW2oXZa+fkuRyNpFm
f+8tnRflSGdoKZ7W8aRzbkTflclcK8QfR+fZbpsk1k4cFXYIRVN4vsVk0VnH
e4WpFvO6E8ak9vcAVgwmx70AQr7eWREBoC7vQVm2wJCr1PCdh+MLhkZFj1Fo
PsJPvuOZmt7oieLBV5ZzI1Axjp1sf6OG+r4XXHy1My98fhQHJNzy8gArLWVy
RaVXbiKdiHUVqS8FaesPp2wXSh362Cvdls3z5CK8ZtnIePkSlV+5ki9cwsBY
1xzIAqi5h40bliD4isUHPIEPWm6Hal4CvgE7bWytoYSxCX9MAbJ73J6dxXaC
aCmPXF8YYhOTa69Rm+efCu8lqs5DhykhHwTtYUs36N7Da1CBDUq4cg3pFlvV
pV6rYJxP6YtelMamfwnyLikWXYVHZmQD0TvWSM4b1RJIgvFo5EtW7SNB3jrA
8/G2Ezxt191oWCj+bzFNI2699xf0RNJtLWOwDMPygU3iXWmb4jjihwGcSpo5
cT1m6LrISPkuwUJym5xYJJ4b64jTWqDkliWz2SPRM2uugTuWv7sPOInbhTy1
e7wze6O4aFsziBDrxyKilNa9HLgwN5DCjDD6rcybw3Q4kKZ52MVeARPC4+75
QfTicqI4Xo7O2dxC68va6PrZvXus6Dea0v68fhL4ualKpzPljdPtrRMD3Far
tVMnTz1JXxRE5XrY2mByXzMi44YCUpU9Uc4q/T+viIP21aZfVXM0E8pl99Hq
GfLUA2g4dp0dVqu6JN29ci9G/ifkzmbjbBQs8MdgrxjVKiiSa88s3mV0PpYc
6CBttsxT4h4yjTYbZwXKQwDlo4VsYqgNiImtU5y6yQzVT4bHvMwOTAH0XPyN
wBVh1nBxfEe6LMQ9+gXB/G/g+rcoJjzgbkjMNDw6eshERtm4plp6A6sf6/a7
kVrbmkMIfieym2kyfJyPjlcy3HWlSfyXUEthQxJ5nyMspTwiuP1ZKt/Of4pN
AXGb7ezZI/bEQoK/1d6qnsDod4tJRUGyqtihECpFioHDcu9H9Z6IaMznrSL4
UH5heN7mmeug74waMSi1aDwIcKYr5k0WKEQ0hmUf/f913je9fu9+O+aYd3B/
KE0VQDGo9Lci4dGu0YJY0Y80qWkPnAyly/x0SNaJE8ux3REztgKWNvMceFoh
816jGYYLpG4jzu6+ix66VUZEeBIc9uaiq9Abfet3wgwAbXF5QPaU3DOkZwOt
cLd33Wu00RwCgCc/0ZJao6CdtgeyItHhIM9/aN6j6RwzXbmSTK4lJ3qKMdE2
O2yNLOyd4xQ6B6aAfnyAg9KSyVpEvxZi9LM+jz7NjEeUo4RaXua7MDqhbSFZ
fg9BNGKmFLtdJIiajqq9eZ6f90XnkMsr5zeXEiD0YxQxa8kYATIZpw3COUFz
/WLEbxprNNUuZ73iqBeFux9G5fqyTSTSnCTRQvRSvWcxTAg8IpulLToJKGf5
q7FjG0vQ+zz4xcOadGsSM7XLqR4USfkBEss3zqBZ7iNvJIkyn71e9T0PkL2F
ZZHDgaDlAe9BJ8gKwdKcha2L1MtnrxejzEykTI8o9pb4I1LMkngyyROl0/mD
Dm3ooUB7gudahorzGcmeKG2yPP2WyAlBjM5GEt5z8n3w16PAAYirnjUwh+vr
uFAUM3hscb+iVpaSORmotMuP+s+uIQsK6nbF9QJrIfLxEnUVsF3TEI6ly3RJ
3TFgrTp65Krdt4aRNu9aZFWSEP908EJ/7EZokFoByFLeXYVu9fmNaouXO3Xv
AZxLBYZLJOeCGeGNk51ZoTI5oXF30D45pBW2Hg2XaKSQvnfnW5QFwzp+Rllr
L9ocsUuXapn9dz7B4z1xUBAH/kZdbXZMO6Ps+GBiS4v0rjmep9xC9+8pA2DQ
/wiF3aXFGoT0LKIycfSGcQDTgZp47YW509JYS/QVeYMlmJPNdzNE0GHgMxxy
pjymwd93+djT572uVQoeh0GfzuUHBQLDOEEUux0T7js9Z/mKBr91Aqpx3YUz
vp9y1djn+D1L6w35IuJknOb4Gjkt8uqWpNMca6LCZZVFfh0F19uqj8Fd7g3m
foBk1LazkSy07y3dZegVH0miHfB9PTNSu0eYSJDoE1nkdEg1zRaQQV2p3/u/
mWzoYqN3X7eTwITM9H4U0nMvAg/IBXmaSoAFaovqr5VKKqwzelpKuyE4apSD
DDIeTPBM2fzKr5TK9B0EYnqPXmWQo5bsn3VkNnWauAqtiqAZXbJzQUjRCcHC
jp7g8jN8HBMdZpn2PPP5YWPkAk0iR4MwgIdgbz+Bt8kAfqPeSp9Hp4ZCt//r
oPrA2RxwXAmp2HMohELqG5EOoK9IS1YcIwZmI7jZKnsfOypNRKAIjxq/MoAm
upMtIBersdiSnTfTafAl/bZZWJxF+y68Z9kb/NNYnhj6zuIBq6Za7dwnOT+2
8yfF4iQuur0ymdY7Qi5IN8RfOh4l6UTDdvhtHVuYuJq6d3Um1G1J0g3qPpSd
2FjTkomTdZe9PyKhiiaTJfZ715b5pW9+x/WjCBFV3XoL9OrcuUsInvGgqtiU
+XWnKCIt9K+gmBlZibJBehG7yPuqC+/JwPXtwXFwyRfXlJM6NuktW6vAI3RF
FTrXZSE6m+tgvFkurbIHqxG6368IXmozLYVm4mCzwI1SFUUuia8ccxcaZjx2
lQQ+O91uzaEsjI8lQRjE/uYiJx+oefq5jg3xJNz2vfRd730nibjaeU5f1jtn
AjE+av1E12X5SB0Y1qhFVE1bUA+K4KcjeEYBMBQTqfDdiKHzBLqAXir7o7YS
PJ/CcMTOppslnzIK0zieiPazwxL+adGl8Mxq73IoQ/1qamUBVrtVyhfWPFzE
SJcTV5redRIJraKy4/0Vj7ELS2CUcX4ikb000CFNCjuOptPhBju+0ZMqA0hD
SZcdMbtfDk5Y1vsMDYRYZn2MvDfviiTylNgI6J+MZA1cShvLkwQgA3KV8xDo
pq4ubvcN8nX86Sd4j0XQSyM8YMDnQ1fOHCdvXYKu1fmdPsYCJ3LtBC5dYp/Y
88JdyelaMxzEGIXNySHa9Lb8Kun1AjJcNRIoMhVvAbk0HoS2cpgDjHaUsy9Z
sN+oU5X/wE6+Uty0V9FyG9XhasYGcRjdODZ/BxvZqXxa7gi+i13qoDTB/vpE
eJCuQQIm8NhPbRjqi+uiX4vtLkpyxne6VJR+0EKgsCNKwwlJJCYjNW37ROTm
ZJs6bzZk2ADMAPw8PZuj2gl2kOM8t8akt3GakyXXdJjwGEFuu0hIURO79aBC
NZV3vBXB0J3WN8UQ6rEd7WVNr9fWOhLvWqETXHcO6f7RT2WAvByNd4DEah96
UHnzVmMy/KS0+HKJJTDUHPe4tsvnBBIcf5R3cVUvg2XW1bsfUjoYE66D+F29
YO+BkQ9fqiZ5ltkf4olVCYP1csro3duDbvhrlaCrQ92PM+Tut7PvVwKGc/n8
qUUHA6ksDyErx83LpEK0aRzw3CR/SoAwv4Xulbi5vyMtbaSrN3brZXsgol9d
9Vt7iQuoaSI1vAw0oKSlrCcQ1/uO3V7EV40pzQ/QymiutzKyEzBZYT5itpfi
J1ArYienK9oHGyQmSHtC3N8C71uACtVqZ6FjXvhkg2mA37Vil23Sjn1QqW+P
OO/ktcw7bccVZ23QGLHZKgQ2SsuTEFz58nJLBLZfeuKn+9ofxp16b91yU64I
7U2KE2jl/VNxDcIBOFGycGo0bS/kv2G+AR5lWgg4xoZMCuDEat5kys5lQsda
N4oCGzaFGiwRzqIRY5f3sflX8EjlG5aFuOWgNAgLatk3MdZqmks8JPgtnNJE
3e9HB6rTQkh0enXijt+ArRNOOycrSJUDDtw37PSlTgQMBEw8xLWot+8080mV
tcQrxrTUBBspVIyxLB7jI8jg7teTeXvYD4kQ/A8FCx3eRaKJg78Zkkxa/CmI
WZ9Aa27n1RwLoaVcnESfzFcbxRmGKCddigVFsq71J2RUqkbC4erzX8utpZA7
S2/EIac86KFDGVSwbvhfId8JlJPAwUDr/DA6b7yxPAI+kuIKg5YYNqUpW9rZ
yxFfhWueAf4AULfJkekx01PIn/Ny6f3x7pxOLLqVl8OQgymXc15zJGPktZhp
pEqaGZqhTyE41uUSFdAeZ+f8FWNGpiyal/i57xYm3vdxaEtEi5SHqxW9e6w+
Jb38rSjKO8m9CrqucbcOfdTtxhPqj/DOdowW8JFOS8pi39bXw1xk0WS12yua
vix3LdYRxwORyYJmflmsCIPixUNOlffvNGl1zPh8WaYGHSGKHFdGPyDzvpkf
PExuYmTNQnk7kagzK0/JCOGVTRrIg7D9fg79f6vW9sgKYbaIDtX+3g6TrGSr
UvYAUvP5srGmz7/RAGFNCcEmCdwj55fsBt1ykjjVhPYwrh0wvVqvPzYAqQnz
PPoodeXlDQv+pZTxniBxzCXST4DEf+CnEZOBCrRuCdeQYdZkIVrBFeMvBFzh
khu0Rphavhs8uYbS6JUxwtjsnjF36+kCUDagWbT6e4TbSm3lwQoZQAXRsSZs
vVbRz71a3P3PSlMTOCVoeEwo+vePW8inRQ2KgKK5bCa0RlI8KPu7vkZLlwzb
1HgL8qOwrFnpZQIL20YtYWqGBsoX3DAAFcwi4st5LWKOMxYKZs6qkS6bOVQ8
l+Y0ciJfnch6NcHmhEs1M4/+yctB0NDa/e+rTffi7S0XtyD1zcqOkfo6nVTX
FGss5QzqMlN6TKpHTQpCaT5ew6T2UMpy7vosSajDegSc/QfKblCky/zUto35
PYhGsjAoS/iyDY57wYcgMaM3+gMEXlF8A6GBDe8EfNYxddF8J494td2gi+t3
bcHy+/HZupAOrLztY6/KnXmy0v0u37KBfsKzPD86S36AJ9f3nhePdknsFn12
wQsk+0aNtMq0fDeOokuLgxSWKLZt3f88uWHXHdlmxxZHj1gSYnD1TiDujlPj
DOlLZSMKWmsKtvlmRswlLYi17xEshDqWJwOEP72qzvKHqa+OFc4dtLnvu2mC
zVP0XCBlJdlthQ/VNSD86gtC/n29fGX2D3eE22JFumsx71Hfe2A1kIIEtvFE
GeqnIXDrwF5V6npdo+jDjJB/EntUGc9Z/bw0QJexPjIoCo1OiZEywg5811J5
igqryvaXVYI14P/lZMPjy+I8S3dRGMB7uDFmHawGJJMNn6wf7O/SU1ALBF2M
MXyGQ290eD1S8nBxhZhaJiaH+FTLieDaC/sgObqXSB38C0RfuWuSEZZmyNDh
opZHkBt0EApkGzjO9V8PxiOanh9ext1M3V3KF1fSSN5zOuNLR1InwiivTtDA
TXa2hoOF09XQwNmpT6O3n1cm1lTdAhKqrVt5LkPQYmjsDb8etmcZiaChDkmb
bIqTK7pxhTRLP8nMxD2Cbmvf9Sc0D24B485M9kYi5SnKsfve4MSzavFLSkC2
De2mj8BQ88vwq8CKYVXW27eFhUKCplI5qKhgvZ7Dl1Au7fxr287s9iakYjVg
jGyoHrd1iiUpCMPykvTjr7v7ENWBw26C2MY/j2y3OZjWSVtMy+xm2n94QvoU
cglIwS8izzA/UyqzB4VqjJLGhbYU8nf2eIjDlXy+V6mjP5sU+0qSLWELmcHd
y+gABgqw+ZJPGLyxNxS5J/qwkmD7XvbLokd6LtDc2O+HGI69SzxwNnQtX9VH
tWoxxI1gUo9OeDAXaxCnkVIgLLFzfaBmC9lYDD1YYSAg/IVCHG/MX0/m5V9C
hq6i08rrzh5Sczdkg8+tfJnt8PCYGHwnyuROlJCDSDinH1T6snyZWfjxs88M
Mk80hIRYoANUcIj2JMdgzLQJTBJCzDtYgQQun6u7OXnjbNqc/bqNxdQjaKwm
xJXzYao8/RNOYFTfOMtdCelIm3GWLqGL/EXQjGxWtVAJaFnkFMsyF5ilVYmK
Ewt0HN1TthVVv6VTFKH0lR0yfnkYuqy9Sp7rSAw8L7THx2ps/mgti2tuYm9V
5NqDo/2MqkDdwESN+MBxpX7T4TnxvZLqL/uVLLNX4M8WEJGcm52tNfBhnvnm
JSSZLitmGTRzBn3VDZCbAgmb536igvXfsdoW13GouDSztHDHWB2sFAOcjlIZ
fOi3+ZUIqIrtDujpR4Fp8wKCnAHkGwJP845U0RROIrUI9wiwR7NQPl+VEyxK
oN1A8HNbArz+XMBQuthoKjAf/RoSrygmr9Q4iCSYGtvXavJxfkFbRvYNJIG2
iiOZlyRIgoXcuXD2zZ66CBwa1ekqEfjaHHLYHm1Zvgbo7UKuEcgz58xPv+39
MxFcUIwtZFBcfWMqE1j6eyBHXwmEsDOKn1cSqx5VX/qBSf9/6qHdBbWZcbWJ
mNEObuntGjcXa9f5UliicDhmo1pYPgUFnP2ibFmRZMl+xJq8dGl80Q+UmcFA
ytwqsrkLtnHj6DuGDyf/XfErm0R2gBvKPCAVcdUrM6iFp/eqAw90OxH7OYoz
HOl+Q+6RmJOzDMQkcHYkfR4LrhVFdnfYKyA9HFHRx/IYrhPkVAlZmHPQztJJ
3769qQnQFYgp5c/oWMY+s88PSu1U9/Wak5BZLEPxp5pyob8HMXD5s5RK/As7
WNyt/21IzUKo39gLxTWu7nYgHpbMOeY124pZxgLYVpRnhkco7KasBh3tVynr
Lm063pV2t1NpsudbwH5tji6ETNTdTIkRVbz+iSQ6vsa9eDHcT/hvOC8rocop
yFSjX8PnY/5nW5GXk+fCu6nJtZM1OFGDsQ8/FYVqXZO2iGdRSMTiGF5bg9IA
vs+orJJGpLWAstyr3G77OcbCqrFXCoA/jIg53GqkMnpaxdvwLVWdO6ivgbHW
bt8BTPOMzW8BHjWEZ/PtDsZ1ys70jR4bJ0lG4/uBHspcBm1pZmI3iRLQFACr
+QTTGeQAvpFMp8zH4vx7jjVfcg9F31LFPHdaoCiEhyemQiKP3Rpud6EaTPK9
nU0x7+q8egZCnfX72uB+kgvk8xgZ4geMVzGTfBMTNu+dMotUsO//CpTZWMnx
C5amT6yrlvcbV5M4F6dzImuqpeS18dSQMnj3QLlFxGVc3br2JABfLX1dTL0q
dN9difclBazB6IEhGOLtvLMhDZnBwKMXu4jY1zNA0/JVWJlXKQAhAEBQDwJ5
IrR+LCReY0pOLhObTY8VCyflIMzrj7tX30i+CQQAn+Lohktr2UJFjdDToz1L
MWTUx6DPQJr/joKy6PGFHnKLAXzxlkNT7QGOxXD7y7fWX9Ku7zT8g/y+nzTT
6T//WaNAWOV28OXSKAVeMYeWmYw8p5ji0BWamSCQ6LqY+HQhGCZrGcbRLAKK
hfWue86e62PRnmSRevyyUZygvLhskNDA8EyDkhcKGJ2lQFpFSTBcu3CDoiqP
KDiv/qkdVerRp+WzQxswCSYwHIGPocfLauKP9wS4BOmOtS7si+ma91PtjYuz
sd86MF05CAdHImUJWaMxQSuvkKKws8LX8MzbP+qJCP0qQ4pF5+NeDkZFhFW1
ULqx5zG3DypQlyaK9+Lp0X0vj2leKV59gy6CegwJLgQ1mkmVTn4s95kmMDx1
ekO3FVChkrA1X5Gv74q1UQ03gZ6/bzx5vP9/T6Gm60ZvaHZEh7RtE1V4EaDW
A+3s66WYoMGAnWiTNltv2V40+5fmMN4Vr/fO0XZRgNAcIViKkZwMrfGJ240J
a3ZFSMkyvD+eqwc6fDLNrKeRZZnjsfKKG1dYA33E0SjGuELJBtA3qytlw8ot
a66Su5eH0LlPkAuNTeqRrhpuGpwnIuGJNS0cPQIPwiRlfjKJRsT9uIa7zbJ3
XoChTWjckEYgb+H1zFySIIbzFF5kvG5TwiQn3GqSgJNdVz/cTi9/xtpUnYYf
mldysatyK+JljiOi/zJgSniakI6uP1Q4TXXSB/dt5wSMTkKQNOWg7fNs56G3
a25bOWyHxwjyrBnTnyz9qj6EzPeyzc89wKilBsHb3Kx2kmrRz54ZxkCnCWDA
xDeb0kVJrY6RwbctyJ+2bJNat/pHiXQcZPHtWdUgGW7cQnM3Kev/PWZqAMvB
p3fE3m5l2eI8PrLRHVRoW9u6PMmKzja0ujE9SvZPtLuCVZtKxuHDPzmInkK6
XLUxPz/nMfFpFzDAsb7ZACCADmrsL5BuhevMnTM+lfLIOdx4T7qYjNKOJZJB
F36FAyxoCAb7Jeh/NRLH9Is8ercQfwZLlavnglPzzb7WUjSuHGrImHhrNiJn
kCi2o8akfMuSZzhZWt6YuoBmP8GAK54i4T5hSMDggK2++cEP4SXoZ6juHO/D
XfmptWFod/5LQGLTfP1he5ZnflNGmQZ3fM3IEiW53Khr0z8FWCKZBE0/fFsX
Og/JOVMf+OZQsw6fyMXmem3cayvN0OVkQ/krxym+IQ7m1GQs6IV3nLmtVf7w
wyfKXiyCc/ghyf86jhi2TBrOQnb/jbcnYM4PSA4h33XwMaxGS4ZaR08ZRiMV
1cwoRNkFZQq56LLe7atI3uX1iG0hF7PjkDNGmjGy7wT/FfmgY9UwFqHAiEwb
lac7l9bPq3EajjSGp/PD5v4ZMeVNJh2J26mDZdhcRP5XPsfKOuEDezxDGOAV
HkgSJP7N6I24FKrrH6TE0GX4v1nmZUQVPoLwSWL2Aje61eOJLXM5ijdDQ5ul
n96EGiKE1JXXExmpE4F5uBDe/kru4ZK5RfJBQ//eMmTJJDr7lTx3bLPsKl8J
wgSaMp4gb1e0b1kEw+RYEyl1wBPTnTVruxEhVmZgPqXiZY2yh6nA3UMFL5GW
TBXeCAWF06fSpgNRNjY4DyYffYc3qWE1shvVcazqS7KxnrETJuzyKFzGh/Ra
vojFa5r6I4PlSNn9fSUoTlH6lx6xsakTj91AkaZrwOY6NhXAKTDNtJRhGi4y
nmSJgQzoP6R0JJ7GZUzuwXtV6MIJzgS5mo+i0R49qwS+XS1/IkP0C5w+QrJw
j0zyTrWXOKFwCEIHtioGdtpbLtdBMSpvuKYiB/ZJWJgrd0vnGw7ACfd/Cgts
kiU00k+htxphBvscKmYb3l190gnEsNRa5olk41M9ovp88tFQmvMbuGTzL6C3
Uug3xIp7tLPArcndICLyrZcPYfU0Vnww3aM3KwV12uSI8Pyakn3xWUR5FHMR
ILT+uqm9CRXVtWIlYekwy2MU1zCvsBuj0STIK4yNeTbnaBC2keOxWm7PB6av
82EEYgr9SNnOKTwxY7r8McUpJjgy6zLaxbJ74ffcLy/+KM1ZbUv5evpshnA2
wOosGrEmXPuzvn5sYQNg5YXkRue8bNzmwu6LDkRutgYPXj7cnaGlpuLXacSg
pf7qon3Ns5MBuWkfJMMA2ytNmbp+DFv7gPHADYJdC6ng6e7NpdMOgDQXZA2t
271UinPWycPYSUtxCCx9KyAnq47AQ8E5DezxkpYpPvgtLfZqjViTQwzePQ/s
tdiilbW0LfUhLSYyX2X9fDYyzeAuPCBwkWoG5w/tzATq+xf8OxwiZKb/AWvI
uYo4C0pg377PWyFGAT7df9r/ZKJytmsfcs1gzxRnf40qdPqLLVvOBiRw7NbX
namKi4faILhBEf4eSyXmHN67ylN9NBXprsvKiq4aeVCeqs53NVQcqIhBdFV6
qBnhVYZXwjng2vJrYP1YhdxsK3YAjutEWQIuQBTHgKTpsnWXMEecAwzJmqUO
Jh3VHGrO4SWOc8+NDEY4Mh9b28rCUP3XeEfELBl3SGCAw1mK6ntUK/bP4QPH
EXBelR5lRkXvT3afC6WjHumOJh+wbQFm9wNUJT1ZpoleKd1nDAmxtJXCOaAP
bGZ8Z9YPqAnT+cQ/DgB5ZgsgO9Tgzyk0DGnU3PJqN2GA3NRqyohlCuOtGQ7y
jp51lNEwjIhaFIeu6Ke+Ii16lG098M2fW1jM/l63dBkS1vCypEOZ9Vqudwb5
CscRZImJ/72aRdjZH6THh98OGRmr/5X6t5JoqX7SolDqMAtGW5AIXKqJhOhD
aISR+pTx8X2p74f3q/ShuHaB9nVNdExHHIQNS9UHclwZheyJJ++/UZCx8nGE
EPtDU/bS9B6kjr6FBVKW/GntzBo4v2HGi6TSjrTEk812SbpYzw0mfW59lCNZ
ZjQl4lkenEDbdwWibtXR5Bp+hSY0shWnFkiqNvggztTsRRpojxMDFjbJWuiP
ND9N5/KjVrAFCleTQy5hTRDHl7olbb8456n/yefLz26uwNpGjhpSl//IwxLB
xkbjQuv/Aga5hsLGvqgvByjeQ5wTUKhlPRjUevUDigUKFcQyEu83TbMDN3nE
HrSTaIQw7cG1f9WxSseGXbHVO/RbnV83ACcy3D41kn/gLDU2AjcqmHHTNEIc
R+CY/9K/P2dCnuP0k633dsnfzy0yvA39sJhHbWYmqlYA4S904J28G3JI4KaF
xlC+ezrcRBPquCZafNLQUsmguQ60tXx7FPZ8txTucZ3kKF9VOFIyDW1sRbiS
Sreq9DbcXSuVQRihOpg5a+CNP5NZ5mK4jO6Ki8CYhVFDuM3wHNMYSMZclLxU
+0LE4n4NnrsG4ddEqm3BIeS83RZUGZjB1anHRboYcHuwduZxXy8PPYYDS6Kd
6R96sU4suqC5kcOLITJukbWetEipY69yv79gUZl5OPkLCZNp5BnAW2rAdlC1
UhK2Wrqm7NQEVY3y0CChv5PSpZWd23OjNrKCh9QNjqFICSrOjlVtpBDzqvlY
eAVOxLtgUARSFD09pZlBoepL4FuomwInIJbmU/52cuFAG9f6SYvGFSX2mJ+z
q4SqQQ6jCUN6L3WoSr4xaTBeNAVSO1yPwmdx7UTZIekensshqT50EFAOAaM4
X3rCGwZgGhJFheefKnHzlgqEYn4eNX1SJhBkTI1pyiVZbDlvdDwos3vlijH6
GyDD2i8p8i280FKsQER4v9Zo/H2i32KU5G48EXzFzVslDOxC0awY72A9AsJH
hEqmXYGJ2H/Va2M2HfPYzHtxgxWZoAeQ9zcKUSa2xbRA79vLTLT2g2gazHai
8QGlNzFOhazcFCRA263AriIA0ubDMZQJm06DthGMsYsmeP/XaVtU5OxFsTrw
TD5m58AW87MGG5Jj03jjLuO3RoC95kK6dR9cbawTfSa0cDpW6ALRWkPHduqO
jE7ch3uQ30qN8ipdvIz+qJD39XufjyZGfagybbzFo8kh1+T+XT0vnhbILlZO
eoAi3eNdR9Hwu1syM9BOerJ+vsQxNHfweYJva3rtIvp5siGFplmf3GyMOXmk
63rmn2RwRrQEWr0wNF7230cunP4BgCAAWiWNC6SsIGTu+MT2EtDskXuKw1/M
7vnBzuKb2gB0d0hLX6bI1Ui6gfE7u1vNw/9Piq90ob1mCjeFW1uxenyuADUl
4tXmoi3fNBygrBPqEpidxj6YBlqbshutzumBYgyUOkvv3w1WmqQl5/QHKbg0
PYfclpv+g1yK/kapxsxwFrp/ROM2CcYFT/GBssBfzw0bH42Nz9yQfqIJFeae
hhM5UV0wv8riXTa9wlGk+4+y/vyH7KxhWGIJx/q8YqlhWXUPudLCu28eX/Uu
MONPEK1GOwJ06e15uUjX2H0yDqj2naCCKQsrT659CbBzKmHcmrtt805y930u
oYUcfeXWbQHO2yPWolx51X7wR0lhDOA7+tkqZL19y6CP9xBuiSK5xDZUR+/T
Nvsr0TW2n/sFeG6U3k75PEAwuaLuDonorbXcnRTuOHl36fmvz+zxwtev4RGN
uUr+DosQgW27dOIsxvJN/PCnple0mxBrai9ViFq6Mjrk+MhdGsx2qsk4eGRl
rjoKeAXc1rVIhqIqpQDW67jcMdHvns/MginDB0pTQy8n6bD1VluS0g56+YjO
QamRZS3kn17zOYyReqhOvCsnxik18yn9c74t+f1ijA6Zncl9I844i8tEBXQC
q9VPnngz1a8FR20P9ejpn4byJ8PI+xo6mZ7IT+kpUKmayR+AMVerQEXBKuzJ
Lwj7o/cIw458xEDMAb35JhDkuOP/dENvaNq7dy7MjrB8CLjqTPb6t4bnHOT2
Zfziv+5vkuOzDkAhITkIN4S8TdoIkMLyW+kSLuJjFa5NqcN9eBmAGb/6AMKF
X1UtOhj7nqv0PTs2z3lKirCfTVDPWkoopkao3IUFlOEKOrcm0C7XxWX1jw1l
lw6i5NY6rXEPN8W6QE9IILMywqbjx/3XIAo+orI+hy3xkfM1GDHnMclWmO1Y
ZxotiNQMPbDp7cBaQQmXeD2GpUcjy7IU4mKqQD/GVwUlrvntF64z8u6+rSf1
yObYFnhDd6o9ZyUqjog9YY2hBUzKLUgbDISEpeHh355iSqzlRWRLGUINYYVF
AkWWkZd0AYaJ1qYUYVt+a3QsxwjmSRGJVyV6rBYa/Qp38lQvB2qqr3ukggXh
M6g2laJx1FY1h88EMDW+rr69w3ii+hUAjUOyOi8mhdgygVU3XJ196pj2vLMU
ykMkFvG0lZ52oRxa6JXMk0w2NdAjyMYw8BT7vKWhs49pyktL5tRneZvh+Hzy
6KJ4aS4Pz5dVSDqhHZR5jxa1jjt9B3/oUtjIiRR6c8kUPdlwNXgqEeltYxnB
5MqXdEVMUuHt8eoa6GPPB0tAR+81riWAabPiXcE1L2/4X9eOS0C1NJMDNGwz
59FvJlzbRwunmrlseqO8IrhewMDqmGSuL1xnVxL7MzCcUjPiI/XSR+W3n2b+
f9vTK7Q39lReXBncIn2/EGkwMFLC3jnN1AZmvClPn8FJIaFO7248j2TAO3tC
9mTgHCmkf+vvmEtGm5G9eGufqQualmKbZEJVt5GfsbkZPoASj6ozTE8y7SrV
c+6uBAb7Ouo/WZ/JKuBEXdc9xWdR1//rVqFXQy7KVLET+9GD7mDTHMyzLQZC
EiEWh8FCAlC0/riU5Sbr3r6tZqXWCG0/66ua1kci18sIrB11IdbR7/GPETOl
+oPC+4VBQgX+8yQ2MXioBG/JLcREwHGH3hORUpnGB88Wmdm2c8HAfhyOtY/T
v9heRZflhPmhg8todnLzAf0ynPw0gNqTMN9eVWfLygBKGVxoeFkUmXdeeRRc
px0ACZmo9lJKWRnnOqc4lSSGL8L53Dhu5tK5PdQg0IsbK7/1vkfs6DlNvLix
AUdMDVMYgiZF9p4JUXplZM5U3UPr71zk9eSrJuUulCtCZ7t7h68NYnV5T9OR
9aAQfOfRey/byvoy160mmAS31h8NPxl+amxPaon8W8ceIiHWalPPAcyayld0
NA9hmES4Bu2NNno+ih0fc03YPGLIuk1o0MakLu181MxPh21p9RmajwqT1qWE
Xf/jEimGNYSyxOAsAOh1lfLnOSTu62ghEipDjwAMmEj4hldLvDfP7ZdLdi/y
7RawRSGOOe6cDHJMmw79jqM6pQ0QMrqgKzXqzFEYluX8dJQO7PeR3UtE4/0J
cU9QfHu+8L7FOksAfFL6HShJ6uxSGeo+hKrSdkGDMW4tMYHmzSQAcQwvJj/Z
I0a2E/kne1PaJHzK7zY36zkx72M1klDXlpk67TMZ/Rmo3VGMWU54vZKmCpMx
l232kOZGhBAqo7FukMnftURpeu7OK/D5Wol6G4kawUxsbvq45k8vu/wgPYbh
uFqdZdcEzeFK2SwGW/dQg4Xi4BscO9gWoiJ/KCScwziMSy2hbbUGSAuhXlGG
npp87ld67Uf3lyDNWSz1aZWbvW7oA6ni1hSJHs2aUP9aq8jxdipjiGlt3my8
n90AlvEIoZXXbRQZW/Q3szjo6xQwLHJl8E3pb1uZd58bbmsFjrGwKSYRChbm
9QFQGKhiH3/AGUSI1BRub65sI6snyXQjGheVsLnJMsoXBingj9YOc0sz31iB
Zx/dV9TGoA9h9HTGYiYY0zGM4EVNdqETlWjovf8hetlqXCkiH7W7AzisLgD2
/QQ+F3xPG8uWcQRdnAIPCPZXMGWHcYr9Pw+X36PMiD2L5FqjTOroxPraLkdh
KNWgTJNX/+i7jkITRqwGLt1fuoPxg8cwS+rGFnasHOdYKn37M5qVNxiWsBlm
KB1hpKinhdI3ZNJqfBZjrOSatubUcA+PIO5bacUr7l1sUA7codxiWcmxAh0i
ww0kh+LZB+1JYCBKx0MkrgaRxL56xZQBfTupdfk6vI9CZahOG3FIb6T7xvVG
ovX6uAmDWxPh8TUzdOZqFl/cx8nCIDiGDT+Shuj4wee1EoNaoTck9EtKZPop
ugxyf2sSEUugTPmB/+Q9whCfow54ATH0Ym2FnkAhjEfvcbPkt06Nm2oFMnm0
pZuZeA8GHRPz5sDVbJ9cCqjwef8KyKqqMaecC9VWtTsHsRpLuv7Q9f5GdHwL
PDlgPRMgpeWBydkVy1wqRGGB8av78VT34PgnZIOZx+3hD5LzaMw0f0WU3JC/
6QeIL5Ur/jwTJjwsKe08GPw3rhs00mwxKRTzTk5xdsyAtM4u6EWW2t+SPm1t
Nxr9XqnxqLe2+uMkrfFScjAQC12P/L47wdtYGqC54oqvbG4WHPckFGOFQDZv
M2H88tEORyDAmw1h3ubmIRVdgLUbxbBslyBrgkC1qIU2RSLRibnHIqxmR4co
m99ODMuW0sRnpP7Qnv+7YJCBb/z82qBawZyXcWWZmSDFUFYStdUpWHSGyjt+
qTm7XWfV51CwuSv1xEekJ6PMoMetXRQJj+9YUeu6qX3mFy9BWO8w1ObodDzG
nluCy49ij2d4qNHyMiYhmYV+u6sPXqVKpdy67L3yotH9610eS561ef2i94uh
1/Y4bb0k6uffF3238kyZv7xabef+lxwdmxrj3S1n/UV7HVXSN+yJhUuQOlSc
TEzzN1+CtohEAp2EIOrqhtX7WMS0BabQZ29Qj/oKMZ2y5Aa/iTfi453foilj
peh99eIxCGgai9eHCS6Eafz708czLBg7XcmUwpM/gKyJd4W304OyNaTEqqTi
2htXDhZX7Hai3KifHo1ZEvAidOt2Q4vBqEcyPQMMTmvNjDcjushufOB6oAOA
4IWKDROJ/rGnbexyk68cZr0BYJq1o0Rv2emfb19FANU829+iwAb4Ebjiy/Bo
hGEvVXR3kKpoipb3sU+d6ukhE6dJY9UhgKucbBSvszD542qGrw/JnFf0zwCl
Pem4Wnf2dDUioEFsyJxIxaqinSWLgIwgbnI0h4kNMMysZ7OH5tdEXY3M6R9H
axQRusLEZ67THyBxf53Db+Ht010/CuOA7IUmbUmXC7SoTO0sAVzUH6eTM/0p
WtY9nTwMZiptQJDMkemTHsrwl6+wk6Ts5ubvBscuawj+q2p4EpVEqqveLazy
yxvgI9gi5COxDohz7lIDJJDU/14ylaal7fT8Rs0bL2yxlmHyla97M3+17TZt
qHDFqz5L7NSlTNSg84LjMQ07xby2qnGXlYpjM9F95El89Zz0RQnC9jBlUoK7
4wMCyvflmbuOM/OwYEIzKJykn2OcZI0wo+on4V/ajOnYbcKwiCM6FZc7/VlP
aqxr+D8fiJ9jZ+B3sjazVnIiy10yVjXfvhVtlKCM3U9V8INcbhYnRjHcOdwl
CM7GrHetXemygVgm8ZZwHjBr/xpsDExkQlyquVPY++EkyyfgFWVhwhlinvCB
zv8KosaVAled6XdjjJvDwflxlbCmLqCxTuTcpUAeWB8l7H0fLGUBKADd8PEn
uu+td96EYqPGsP5sMGlnR+4tdRhqRPYnlon2ZFtv4aUu355E6hGqIEp65M73
/ey/gEYTR+lSnKiDuEUlnq2CmSYvJOqOrT1pUN+ahD4z3YpeWrqKI7AaaPQ5
haMa9SkcFEpcqSUEnlkkMF8hCjhfXr+X99lS947XHWsjCV0nNptTpnwz5g6T
vGBhOFUGK+ON55/0Gi9DwLMwfGnAydQa4KI8tCF/BWi+m2OVf4ouQe0DIrvu
jflXQPnB6o2lkpGL6lZdy7rRjZ8Sq4zyKOQEvJ8OrpV0wSjSz3rCWPEtL3hi
qMJpTmvmpSYWYeNMiOWTySs/+BliMDqTw2/ISlgSZVRIHUYh+Y66VP7l8buD
UG02x+rO8vR7KRa64evLCNwh5fcgikuFPAysVSs8hpFEnfvI5BzQDpD9QGPq
Btvb8Sis0BwWq6qESfmUj2Jiod5SzantlVQKbpYE8Fclwe75/cSTzcfZwHDr
6MgpLGfm9ELjkxpGItwsc3lQ+tmKQZ41rg78Y+5mBOsPxzLTnzfpJWarZ2Y4
Xfju/J0i4XkMvnqoX0j7vX2NUG3OvmsCk3sS6DIAJpqFSnRVVSrRKRktLoz+
uNicgpzzcLYxNVC0CDSo6F/iT0f/zdzc4Y2tCdl2HrXadp5W5P2J7CPf0ruQ
9mPHkhaZNS+XJ5lfThsaQ77buetOI/IVEmYfFdkJ8L96BORgh4lscxS+6l3R
Sz8DHQI9d/Ozb4Ewu/37ycCu4IHCbntLrgBgKxNmhyR6WTJcRTAq7AaqBU6A
ODz2OWlXFffZgq4k5VWb0LTb31wlsOJ1DWwmX8JnGjztMeIYUPVT7M/9jo0D
kYKYz6RzgaN19h6S7GpDSdOcA1YghkQtHbmT2FIbkBB+aY2H4HC7LxG3f0Af
dtaZh5cg3f8VvdRNRRkI5De0sr7CX8X127WDfq9KA+aiQD6ZGca2e36TZA/3
SMaWeYe8UfOOFvCAVzbOhvao0qKBC6N2UAgn2Pk+tZfIThs/9sP3a5CrFBFK
wa3mTNYHCeowylLjQ9+4nazvAgI04k3E/OclDC0XTK54Lhtzd1kydjLePcvj
EVl9IdotfY2dTSVow+jZ7vPivKETHya0rx3g5ltRXRcVKtoRJL8Xcyy2Wmh1
rG+nNudKt5AoOhdpJdP6Aof166B0z3yveUI6Vc2sqbN5nH/4vllC+V/yXXl+
br1rQUcX7sNxJjvpLTx4Jq6T9azGW7mqEcHXh/PYCusLJyWBnQ6M2Wh4EpQH
bWMQS85H8QLncI763FSILTAvV0KmB7vY4p4wv2sPSTLP4lT2K90b3JqiA2mR
MBUsBgchvL55z90On96mqA4SOaOXERFnj5TutF7ppG4qp/idAcbhTc4gQwXT
LL99c7ZG4LRK4rAo24yP3BCuD5y+fDTRCTzq6eBSPQhkZoLtwAFJNMPcZuNb
CmmeEjNSib5pJ06pq6AyLUvLFT/FxFtHvt+YTzbD25XMNBL57irbxBlE2dCw
EFtEFgyyqHiS1YBK1om4cpIOB4mDyqiBr2Z/nfwZgD0c+mkWCZ6TUqghKeOk
tlzH86AtRJxQgSJyaaBDwYi99BRTUwbZCCMkgkmN8Gygf0QPoWpmBllFyMF2
rCOjY/X1aEyFjy27q1e0DbmWORCEw9kt/coFmFJ/h2C+vAJ8pzSbk8rnPdKx
G5KBoeqwGagAp558Jwa2nrY798iCKfmtYjssM7rw+lzzaPgX4owoOA4ADt53
d8rlB88zX3n0J8GwVWEjksZbzb4Uz78MH98Bzoc2aUfxxDpsVZ1UW5K0GP+U
aPWuwyx0mlGBhdjpaaD1wjbZn63XI9smIKrSCISaDSnaxa7JU76CW3xPcCJW
nM46uzWIgLfDnLXBZFvSxfdqRS+9UZEx29JRlnJO44LmOf6gVv/HwyRxUQd+
GRV1mKgxIdUXzzrxs8qr9+aPKUAa1E6Y25r6nt9yd+r4cMrrCOG/5DW1mr6M
n5Mdsl+bY0HcEbuTYBuP3jMX2Fi+UabSvZk2BOU9isF8mGmFTrsck0M1/gWK
WyaRSO02kFE71ta0Rv42QcUrHU32ehRaX/4oxljKwibVH30ESFOXBsRR+zBX
DW1Qi/L/0PCF1ZDkr5ES6iTzBsJg6PnLTIwE9p0Ejqu4dMK1Cv6LWgpNx8Sm
RtVILODq6hETn6xmv90dfyOwiYOxFcVyPzWbPHLWLm2BnknTh/Y+6doXNOsi
PAHD0tEFy10Ib/stLXOYiL2oVUfkQd9OYpiObnA5uF3gyAdxzhpVPPqjqGiw
oOEAy41+DluEgs3R5gb8dPMLPdRcT1O/0774iKT5GCP577aZMQmy1ZaKZFNx
jbFz2k2ZyzXatWoL0Evgx+Es10TL4eGBHG2bd9Ah1h3SmQ2CwDkzM/6IWHRP
+x+yilHEHJpZI7SkduAixfiQYJy0K7L01cL1RWzO4nVdQe7+EwD7YNcV+xIN
cJq3X/DSfx5p16BGItQg7ejHiZEJRYPY4zvX4vHm2EqxMigqvOInuKYHFFxw
25NHrTl8ek9zYv+z7LqB2Ue+1WiKgbVZ2s/Uuo81J4K2878x+7S/6BjVIPHT
gRJs5bSirFeFeMbtBefd1MvKtHLvh+DO3DbtKGbSie6+egEJfgcElYHdyLS2
XWedV5PCsegwSEj0jV+3T3kAYyBRtKMskvQOBfhNaPEnTwAsagxTqwIi+YAg
SOViWVnvM97KgdVTRVSxeLIi1v6ij5vZWe9xiLl6Iq5mSyQHAz7n4r0pkjjG
8wrZ+gm/6LVMN7XpEhXREGLT9N9MdH0vAAaWAQfhvd76zcNhNIVvZD6wIhg9
fLlwt33v1FR9Ddn/bkUoCqItrvUbfFfKuXEE09dcJ2s39VpZ+3ZRHz4EfYCb
OwYq6xGb4GiLarhjxMxsgV+NROD/k5imZGIA3cYzvcjoj2kFf4w12t4cmTpu
CLLDsz9hwLrH2veb1sa18Kd5PT93yvNlTHOfpJQBTREWB+1o/idOxPju7qEW
zmbQONq2WEHNhn1Fq3qm+T3hstFxiqTKMmkgtCi1gSPxUniPNpRlNQbUIwXT
iAvkj8rCRxyIdzR1EnQYYleCs8jpBJOSFRjsTyKHpsW5aCQgEdILiF7JHaAP
SS74QHKEGB3HHT8zKyTczJqu+93qh3TQP4htrdskWpiJCPorpMySr3qFiEai
1uScZDZFiaUjdHJ+xpDCwc/fAdqteveNDaiV+6iafygpfaA9+on/kaDf2Grr
mZd9GV6KpHCken2j77qKUzYvhXFoxR2uF6np6GumZ9KojNJALWCb2KP4h4ad
x/zl2eEn9impcXV5RQlCD1jGQb8jZU7zSMaW0gPre4TYCOIH+aWsjCJKYQAO
Dh/FUwOZ/0vilydkQIxsxQ5ILamrOzHo4vjSMUqQkDGGl7+0SO0IA1A23QVj
5wkq/ojj0SyNTs87P6GXE/0JkVOTbdrwiMCo0FRh4JucEbfWWNDEGcnAqdCC
O+NSdmT1QTGEuhdFtRyJz6dDHWKkM1LsSPA7KPNkJG2aTHJTeDXUtZlahcEv
nPOmybCr2qDm3Whppevoq2yz9ZUIUqJLM7E9KMnQBJ4QY7QospQ0yrO16phG
xGK4d/gUsKQY4/A6frPLN/iCWee0I084W9FRQeQC3NHLyMgTdlvJIvN73+on
eV1cf+lV6vfWf6E40Ui8MH4iaoCF48QscHTMZ/pBrqxCxcKiKG6oZ+JqsOev
UOwzmOqg8QjOxZ9FcMcNvu/uqqAR/Pw1XyYZB7OsA5JbzdM6xK2qN2l2e82F
l18VsPLlG3ULgUzNAeyU3NqdOjFcbeelR88RXQF7YIHkRF77tjTdXAjuvu/C
qWFGam19BkaiwH1zcSZlmuStctViSM5AVygM5XQTPB3X3yaOyBUFDdXEc7SA
uTqBh74GUZCAxyPi3gM7lWsPWqQa/pu9OnRvkSuSl6GSC0ghcQl2ossUed4/
xeQ1lDU3E29sddUSZO13GmyYFv8A56S0zDgnIRtuBumzbhf7rgIUgTw17xYa
E6jSzsZxoQ+TsEHwmC/n0Tio2p18wlfAzbRd1mNTN/Zm8bNZRKz0GFRRDCrR
JtqQmNAEWX7+UsJdAO4nyM5dAnD9bghK3Lzq5LpLEfH366RfU1Kyw9lU2PjH
KPT44n+uQ3GxFJwsbG8Kj4QbrK1LS4Yio0g2+27yzPLwUxuiDwdBdZzSVRmi
NiqptO7byNnqVmW4vTLcG8sLSB5JrdiXaR0CYSp1LN6uz4PArMlSlYRN63hV
7ZxYQVnd6D8flDKTvU4D9gf4jybTRdUjdM3Oka2VhqC3e6bD/rgKgpxaPmmf
oOLhgvHETBOhox6Ozu6441WmbxtM9Pxi65drsU5J8H6UdWoM4uITXUSp7DRh
17KRhmYye8xAiil3UsIXShlewDt2fHbdgvyzU6LfXGZ075akMWWpOI8o9wDf
HuTrf0SL/MM8JocMlohXwwIDflVKKu3FsAXG5VRMtKuRbHz/P48HUXjoWRpv
tX7urCob8PdVp9qxHnjCZmQO3y/8MpDjzJ1BMk+8jSVcX1ZhnYqa28EUCPT6
/w1LESn02eryTtJ+jzV8Sz0S4LOa0mrlsp05ZhiyP/7W7hugE/cmwxqwjmdX
lMa7O91sVvpbH0c3apE1E3Wn/pB7TeDtyAiXjME39MadJzv6LGALYtwCgpoZ
Xjc5HoctwTi5JDkmvRER/urX7JfIm84mVlQxCwd+nt5MHGwzhP/PBBRV1M99
OISGnJJCkjP3NW9WouKiyu/sSvlYJM6jp5BfctGU0GBEcpvSaiRf8sbDXt1Y
ZnUjQyMQOChuke+5ubQf+MI4zy0ia/2y2kOiKZ639dWNr4nYkKSFbpfKxZzL
o0GPezy1rDyqEZ8R+1mx/Jp530uZW5BDrnOyNpmwxK5dy2QL5d36FnC/R1GK
NEh2sypHxcdRiB9aHA+qMATNkLEWcW2a+3E4GvlVBJ1Aq/0+YIOrmnVPojZD
4hqDCrrsxtuOM0qO/0/uZne9FyIHAHMfMmmYD7ng/ZnYv9Q4LdQcSKzEutsV
BJYAYSOST7G+YMZqY2bmw8+vUEIYCAkrDHkEhuSULSJ5KqppJPZ00Bmu6051
osUXXQRTMWYsplliOEjN/jfOB9PrEat2Hbc/EILTRhsHO+f7iEARq5NyHIJc
FJZzR/DYdwBiMa9Kb36H3VhvNByXAcgJDvznx8Er1U7VNeVWzp/XaQJF/CrC
4zTUFwHXRPT4P+q/cHCWnLXniCmRBGESxoUOG9UBjnsMAK3X6vk4c+KEJbPB
Kav3VqQVGf38K7wSF8yXQn4cWXxqqyQiyI2Pfu1YROzqGIxqATxv/tcL3SlM
0wX8Sx9PfMKfw0v2jY7Eh2CQYYQjL+O2dGbrEa+wvaPm8xslHOlcU5ixT1Hn
/rN17dV5rLHl3sN6Y3/MdJZwh9NorJaJgPiBT5XhLBwq6yI+JyUaWczukFxW
kXHyO/4OZI+LUdHvJ0pxYNPgK1GHo+SnN9XxooUEQ2k3Q4rz94+xlp92hYf7
s25aiN88Vn7flgP36a0T62W9ynLN3AmZTTTygsogC9wPB8gwD4/NovXAsrDP
82vNBwWqg2rh8TRlMu40vFKYJdOilRC5EcIipz846zPbVoPOmkFW1h1WlyyY
ePagJX5iNtHeuaWDUVav5PvLrwmjKJmUIKP02mQwcuPBHOTVwXG9kfC3oQv/
KgDhgZcuMQCfjTeD0ks9AxxytT6ifpeXVQKD0uTsbV5CQ/Fd7s0r2RmZxIrU
pfwCa8OrAqRqwpCGuw2tloQfLrS58/HNUw8I0M1slYUvbMzVGWinW6OSFLpd
qBa8OdhfDspUBXVXscznMAAH3mAgHHjozswbapn3hq36cjnS+UtMMXE2JYBl
Y4JsMZ+mkxlLSNJZwV0egvyp1nW7ikGYOO44UXGVWtfftwvZ+ggsAH6XvGU/
kBYpHkr9w/4SL4kdo57wGqtG7WVW9gpIv88vJEANeClVeBl36dKHt8cytnut
O2PB6ZjAiTNY8Uj+hzAAshGqaMNthTZrRMWvy5dRW7lnaqhjzA5XQYGVEtst
WtZUO+MtBQeuLX6HlQ1yGe5O6Sv2r/w63Qa5joP3GYJ40P3sOPCq8UhxvWTq
hac44UJ09boGaLi/wflxyRSfxpfzLl9n7pBQKsA1XhV/ceuYDMrCymbBfeHH
6mgzN22dwS6Yp7/+MVoLnsTOLtQkqOnPlqdvZ8sajDcd9MjYrid6qfbCUNPF
nuEfk5oN9vlRW3qsytSWCwTgmJS6O7E00K4cOCccX4q13D0sxU83CtpZQQT0
pCNxGdq1Sb2ZMw+IiHGx16NEOE+jEJjJhOV0dhSAMnskfsTk+APizSoeIJuB
1lXl7GGButlfJM22vSH3Ym915g3D+BoltccNqVOaEg0pJvBbc1HZa9FnsyW6
AFr85XAsCpvBTjb9okiy1u22rrcXEJA8VpPAlG0HRKa6/nWlTPHEwqHNW89F
GKKs3ADWRHmnCmY281eG/W8l07vaU7XNKRczRAHq1JjMVq5RBTzi+JMNIVM2
bwmFZRr7o+w/UBK+3CtmEvItfz1eLORnRKrM5h8skmTpqhkCeNQtb4cEcRuf
VpT5M1c7wwMYeDXE1WTBnnYSOfjqVcmpkqY4PtiJ6+I3F7zKYkNXuCzS4Nj3
zVoQ6np/Wr7CNZhcmjxtcmEfodvDL0dv1RXqvMsc+Q1St4mUS6ZWzpBts4w6
vYT8HLDRT4Q/0aojQiBalpCttMlCE9bgA9wyVvHSx880ejL3vBTHACpY9FBS
eVJz+uYHAedbA5yLCmy7JjNm0Gc4mxpO6OlWMcc6hfVlAUd8BuZtG8XFC3UX
PTHPgUJzWayTjy/1/EBScBaflaGe/Cneney5mxS6q49//Xr2hPPqB06eDlLg
z5lt26abuAA7dFZfZRXsK3cmiMJv01zWZ5f6xhPPsCV7/JjBMdkgQYvpHLh4
Vu7O9/+LN/9Q/fhENMekZKvtq/4Tcm879poMiGZ6d8ftMPsdDtMdGggnk9Xk
XzXfiMmEvF+q8OqhFcv6bE+JQYiohv29mMk317KX3HlayAg6eWZHrfb9kee1
5+YHdkcoakRLwkuKIAZkiGNqPadusMoTAphMsp1I1SgEj25rqK8lfeeQtcPB
iMN06fBScSGLvlL654EykRFPVhBJydKfQb3xzx3rgiRhbns+i11PAHIS2fwI
utyghvIt8WmVX+HJQV8riksPZrngkoY+ZAGoAqeoxIiek47P3krg0+d3FU+y
vS1E11LoMtSvEGlB0RiINyc5leVLRPYrREE0A472F1DCwajULtTlLIlcV5NH
FWjMsMFSxIQW9JzJqCM3EDQ6/sKQHunL3nkdBoQZBg4eKyXqwCNZvZV+wp1C
oJ6xNxUNiWox6Ss6RgNOO7WBv/U+tyzSh8YawUYVSzQt0jzVRbV/q0+COAgR
XIEFRq1kZh54nL/JiTVZyX1y1I7pNNYn5lpJEtXB7d+E8WC2yWtHz2Nu2rOi
1aVF92dVw9uywiAPayyEhPO32uWx6Y+Vzr22YYbEFvU9SENd7HpUC4Uw/ekT
Ffqb3ahZq2hqUgStmOv/R93mPifj+2gN0VwLBthXoGDQyifd+YdvTlOWVw4q
lfNKj/mRLhW7ANZScMKScurdC6PH1FBK8nKEhSznEUDXRgMlj4GlXptM2DHp
2iK9QzE2KYvfyLngEn7ce5/EeLV1ReNKFqfgkHIZMg6wtvlIwqEgEq2xXAJr
m2sjSdjmABlHMEcw7UfT4sAX/+iy71sFZ716rNydQQZsfC+qgeYsdf7c0UEb
uipJBDny/KwS0LmWZryML84QugAjQLzecEH3Tg5LEVCj2jfkyXAMkbdEnNrr
QjT2f3eHEX99ILJUybO3AgFmC1kDjm9ZsqULbx6DRfTrlAsWAW2JGEby8els
QUYdsiDBVA16BS9N3y9BKeBYbxyYhm/heQak6wDNTErAFZfKvS2a+Ag86W+9
tluTfCcC6lGVa/vShVPaCmy9QwLPJfX4vru/PsZ2ODxCm4kt7HfPEDLmInw6
tZOiUXmV7cXW3k7ZlP7/y43+0h6QhjOMI8X+YzaZpVkihHo1lkDKorPiWMhS
9Hoqck22UlY48Ogdt9zRRTiCpfkzMutoMRqwJNmuxZsynEiUiBG6U5pOp4Wj
0OP9dYxiqC6uLa3xtulAfY6XT2baFFQTLTVfl1Vl69hi0YYUzpgS9riqXMPo
CeIES2agkHRmpbwAge5UOrpODvejrAwfl30eoIz03kka9pROr9GGx3nsEwh2
WylbXrTjSh3cfOibAP7/SgjaHEG9duxYgC9omRiR8bcRsD26ol28JSNLzpqV
TULLitCeT0EX/9B0aSfingz8Q7vuo23E3MkilSMHUiQJlZrPE1laBD3cVUOc
IUVfTQYlk1tLMr3YjYRHHVQsrO4dCPCe6f26s8/olWpgoLiNhmFxfxPs6Dlf
8iOjATWBe1nUTs3QVR3+hC0cFmN9mjUtR+APcwvBBUxzQmT3P3pSFrvASN3l
+NNC+93JrMFVx9mfINY5v1wGHnR2SUtWLCIaAS/dp7Sn70o/tA6HwpuS75Kf
Sp/Sfl8lH3AuJ46xPKEtUBJbbEuiiaYLsrIiLsy1CH+W8rbp9DxPf4j0esjJ
neKIyVcQ4rs34J70TToa5AHDO6U3XGDRV+EPk971ArCIi7bzfcZsYePDBH07
z2eij0s8YpTB2vddIYFn/gTxq/HIlK/eO34ozaHD2h5RYC3jK2svvVcnDLJI
VX3unP1LR/jNzUcfhn9XaOMXwNq0mf9bfHnp1H71ARpj+BLiK4GXxJypkKFi
L8Dk+AyLQ0FORAOxFG9ZOqERAalI1K4B3wW8mPGaKGJ3xvnPQi/Yo10OR0YT
i1Vxo23QmP5n8WCGzgnSB3NgIeo+O7c2TEA56Tz/RtLRygyWHxt/K+jEPIcG
42QWL4YMyQTP77yjw4f3JfgNShizs84oPezOLZc7rUFs7PfnGtwtT2CIlBbm
wNFUc/Brg8uFvpRFfAp87DfshlvGZVXGBLH7synyyWX/3+CruzokZ18FmIRF
dxE+got6Hek9idjQpJoR8DG3ZMqUmAVrQh5tw1Xh4ubACnpH7nOLwGKepqdi
eQxEyHtzviPh3CeSSzbvBOeom29dDZbrlzaEJyBkycJaFg6+w7Lb02iMSu7o
qFV/tBZDWb43M7kqYqlA8XrG78kRSLJnvl9nQxVyUjn3V0pB+haq4MYMze7O
oodP/XdnnvlyUy96vgsuovztcnvuZr884XjthgeCfdr1nFL49E7MCkpFblg7
dibLjONh23z0iXNngiw1XmIRVILbAYBNYz/+7FoMmzGxkmh6ya+TZAQfZSO0
6TL/8n+pkGdmYzUAHAmhCqDQeEWHxj7Hmv+l3cciAmhHiWHnGoGvigWtdKIq
36JxjIkXaaVt18hUUvmuAPg5dqletxKTvBiNTOAjBYcns5Hrf0798gjbp7vZ
7/vclOVcP1xBQItSfiSJlTc3mIMv8OcZsS9deryH/39ZDunh1WJ0vGHwu7qd
n2SskPr7NgkkpYzrYGQtkCLzgJLkpiEP35v/YgzUOsMdAfs8tMP6KSVvAGwC
GbWAaA2qkNiRNAe3RM/Vs+gIwS/Lqzh22xLENsvPkAW3yNy07YsD0lINCOMV
iWn6Ah8xkY6WvwF7LohfBtMlKwOzynG/M1ZDD+PhfPbZg7Jqylkx7io2BoCU
CzjOZH6s59MHvVHGY4sHT3srT/UNpOU5b+hnhxiVrYuWb35LXKadhQj2nMFe
6VRdaWBET6djEwr3H8NiHafGXvPa1ir87loE8/YiXlgOlaYMRo+8vAuh7cF4
u2f8030DSk3vxKT4AJn9/89CFTrYT+2M9j+kCOAAXWaeR+TrHigyHVh0SUXz
xNX0xSNfIl+uazky+R78gm4UQgDf7wTsKD3q+selxyvotUcsRna4cv4s7Uol
1we1CFqCT5zXy5m/Pk08F26+JfwlBwWbImuoxneWpVzoQbhSfwGnZNbmYo1U
bKpIwfrZRFzyiwEI94q0vwYqdmI4/p06yYwu5zH2IBcqexR2LT7/wLId67WN
E/TR3fza7/JxcDLv1BYAUbTcwdqo2OYetBZp2GAEYmgaXG1fGLrRtXvxhDG4
9R+uFdnPIm1DyTIz1jL4QocZR4DjurcMy1NiZWxr8MEQLWpO6Xc3mEhA5i6c
636ETUoZ7iEfuE5MsojXnNkNwpoId1A4ny7GC1STmsEuT8aXGkQQtJi/Pl97
vGRSuQp4gtIQKN4QfQc+5SBohCA042TZPbRcNMi1JZW967ldF+a0SiH1mnBU
7wj0AIpHoxb7BPXCADDOm1I8vW1AaFrWHj383qFbQc0xkXllHiC3U7bq/Y7F
X7sAMU0n8tKZG0BPNWR+7DAHEG0hPVhsULjis6Vfxd39/HgsMegqtQ/+ndLe
4x5dxzDaQMwtGB87TZhe2EqyvKY1WNa+eyBJ13EF9CrdlbMVdbwHV2vtAslG
Uamrr625gtFnsuZuDU5KK2ITwY5iff88CiW4DbHCeP8fAk9+QHIigaXinQyI
K06epf7Krw4x5AtY/6Z/KaxLaHK/GlEBkArTU99U/tnj/f+l8wgTtJGQJVWd
G3FB/M3EgAsmZ/0aMZeCPgXHu7wVl+mCc2CyLpAxifAhdrwLx9EUYoYTaj4o
8u1WRo7gopNn8b8IRpWVAsIdOM3bb4HgNRO+A2ohkEkmHeWnmYJoRRzqYdih
bppysJCqMr7PgXE1f58lhr/sNSCp0YYScQp7QxPittWldb6/NHGdbj97oA8s
fLWNIQK4++nwdZlMgpnA1PHXu0mGBdJ4cKKqX2envc+Q9CmzviROARYdWk1e
71mIcnhrCEht79EKNhISuhUFSpRYweGaiquJ3nawKD/z/DPCXBbGsfh9bJTB
D+PSV02QaYKwGfMuO8HFQ4efWSA82wsvQ7Xd4qCVM2ShZ5Bzacb7m7YXQEXh
3Jcog7mJoysXx2xP+7SfTKKsjjR8M9gBVv/o3CZkBykx0UXG8qcahLZKjuxO
5eMYd8QY0/tCEqV7YItvLfuMz+S8SaGJirDB2IKusMqvcUyIAp2GLoUS5Lmr
lCaOhC7tG13FrC2LrCxREOXM4j03BnOM102EntTEugJvsIk1jt2icc7bQPSc
/U1Fp5qbNabj2/DCuaB1qUVWYWskWUATWnzRuFGzgP9Nq7cLh9O098xGvGTs
NCL4KFpqnXBFHG7V0UBSf6ofb2ZGDW2MIKQJC6MXv/5JKOFymzklGKN9UuOl
AM0gnwDQWmkFzswKL0dpaknn/bySBgtIigrLFdpmEaYmQ0pyNVE4FD+q3gO9
jlM8nrwrTAkyldfaqb0ViukyaL8GR9qi/uR+AkDx4J5SdaeChP4Li7oY3qeV
lTUa576AEVKNH0w3SOPxq1YeW81kexW4AIPRZRdV3x/YIg3roB6hKE/N2qP/
HbMHTVoTs2j51abaFqiX+g5tTeACgQm881WqFEkzlgYVQQdT/Qxh45EMwjk+
yyqoU4aRbZ4WZxpSAUdgnDGCn7PDDeE6aSVi0gIMmJhNnjPIrKoVHMCi+ssr
DNGuzwQ0C+Rp2rxZyx8FWvrA1oXRoXzwLGqMttGizU7Tsbuepgnwlv7pKRaA
TF9UwRYfW15t2ZQHoJSDWdjHMBEhANbQdvDSPdkXsUi3QqAQ3Z0YdzmOGSLx
JNPPndlBnbS0GZ6RM+PV5gxLRq1WfQUVLU38B1LCjS8I8LEC1lEpADsH8uc4
JXdI9niPdcJRqOfeL/ueHHwBijQvBgZvIRuGSje7jaT4g6lw79rRP9O28rdT
eK7OwNSwM8bOebFmHJFRyzBqMiiNiJ9wXH5fBuPQ88DNad6hmXbUlD3EmGS+
Q6fbm2nOQQR87yXGKVlR3A+jdKAHVr+zwO7hCnU8d2HCjt/AVSGOu/5FCYFk
nKdP8JDllCSBn9uwxHEpUTVVvV5WBPiY2T8I+7K1sGERICAtQZ8nFr8NQDXM
7wgTNDUakElPxy75HvIs6cTLYkVuC7vb9/Rq44yLUS9TeUklRO41L33ckKBX
IR5jgnHb0h0ZjQ3pe+hmaB1woIIeSqNLH5hMMF63Xab4kXfqoyiX+foG8RzG
DkU8ZQzJ950cx4NoJfa1kSW/iv7hHx+O0erarkasvCeYbhNUdtTjTb+k9wPS
6HLz6Po9GC2LIkAYFtrKgnzwcE6g1KGQwnGJuDhmSYfsY8pQLLNxFsVVE0yw
9H0Ecmzdj2kvV3U+hl96dDLSou029KZe2VU6nY6hi6vMMtiq82PXCvlDSopx
hYrILtR8Vui7OLBGMDchLSpMxG804Ma2ekBkxnvx8EimNbILzpBTr23rYUqn
OMN5qowdRFgGwVc4pgoA5+ZO/Sm+k+ttgM3nS/OADX9BypC1Nhka3vyZZyQx
I4lfKAbxaEsWslBlbdYdmU8lzKZa+eP0FJfHw2oSlpJErRid7HCTMFiLSXzo
Fdw3btcD99x4URcta/jzAG/U7AgpaMUm2MzklYq71AhngYFeE/hGJXDvDn0t
6sOwnUZPhZh1ZKpuU2Or/mOiPXCmBxpIW3pUOX4axDpE8iCPqhcp2/W+7l64
uNFKoTBO5zzasK+hda6OAzNytxs4BrGrK4pj3rhySomiy8Cg7RXYGG2r0pGm
FncjF03WKl+bXXr8+35hrW6IUPmXDi39V+hYFiJ+enwlH7XHCYyT/hkoLW1t
A/SeRRuexHO97Ac/dDh8a7C/nlYp9fX6IrrFH0hciVRDGZWmjRU8Hg39qnbQ
OeAL+Lpq43iZDeMBiG1zJVFgbesK1D2/fNX+5NXmMb974JkTs3Y8IHZ/M9cA
LWhOYa81rK5nneJtzBZdpt+j9R8Jbxb80qRwZ6WGk/tjpZH0Ng+eL0cwdu3m
S22KT2ppB/W1wvp52ZD5oT3Pv7ZQcYfjvLK6LN/kH9Hv/tA1OBdpMhLuNLnF
o4GdDxu5EDHR4R4y7LQo5KkJIbUokwk7of90SYZgdBKDw/5mpy+ZXTSpvVT0
RPvZtvRvzXVqOd3XqY/viJHaxxWxHIDvpac7sOcfrtjNorXBjcl5viooc67H
S3JNsu0b2BzQbDjJ5h1vQ22qKRWK64FOhJJ1A9AV46jjcWBmoWvwGPNcro/U
JgJ4hEG0zg5f+fTNaIW644cXn23CRXQLMmLiArZemgibK9g6AGr3PqD+Knjy
6H/9yVsw3LnJRDxlgZtGlltpJoRwXQyz2ClSbhzueUYCseb2y/m1rthT513E
kOPA904xG9xHSolCtoVDDiAeeoChu+tnO00prhajB0bO8EIgr9Tblf2VD3n2
JfZZC/7dX7rH4AxY6zfYtaJub4Af5D/cAMSfWZX86hvYpXIikLpVoaulYojo
ndFmxajZBMCr62Ouom60ybmebLU0w+G6lFS59kUq/lJazuPeRZwxqQeKB49s
3Q0247WAjGR3tIFSazSzt45dDRthGXdZ9in4B96DsOZvqDAqB8beP1xVX+xe
EaoFccRB03Ja2+zavrVFnp9qVDpmfpRjl9lmUKlEk92ZzAtFzdccs5rAtlvr
IBK/GG7yHHeGZS0k9BX16ZVK7uOwIXq05uCfsROsCZdZdguJeNLX4bDaduej
2Pc4Hi8pIbf1Z1wSTaZEKQZdb9jNNe8x2lUgH9r4JU1hr0XnsB2ioMXnlNVF
6dmkrwGQPKBDFabNfXZ33Z6ftMnsoPrh4IwA7ejmyRLOHgg+0c+wCUvnFFnG
5JFBTjHaJpImD6KPff4DNig0AcdNwAEwQXYTWRNw/lCCYZofLBRd5q6QLOAc
R9WYvYf8vGJUFiI2BUiWknMFaVqqMIexmpJGfpjw6ogiIwYg2k/cvN46LFeC
5qz/vXz4bgfAbPlhpnqwXk4G/l+pPzKUtWsgD5jyeeBQfmo/fQYJVVChpowx
nMkypYSNFoQqwGm+FidvheOBKxi072BlOhHfcrCPpGyjd0d00tSq+ITVBdl1
4sQLY4oWFytx9XCH6X7tmZAR+pYPD+CW6sY+mJsdbbC3c8vg1ZlE8FMyWDru
Sp+HYxKJzL4AEulr1499i2oGZt7RQAJ7d6VhglakY40CB4yPSFy317eFkisY
amLy2maBgj+UHq34EwVK5RTdyJUeNHpw71508anNcOZfL82VuO7rVi+MNx01
bO34UTL4Wo6pbVEjQmEnq9g0yfWItpKUQG95FR+Os9XaiZEjs5rTdXHBYWio
/VZ+d75wMT5g3ylvfw55yAWD7MV0B5AomNecbJuEx+zqmZZVdo62smBUyfuI
/GFLCOYP9TGSrOPgwcAdpNyv2Y3tQJhnPBHW/OMYjJim56MVKJQFoxaldXHG
78UBTMdB5uxWC3x+beJt397lfq2tGPHw3B1s6uCOzm6UlzPQJkTQGznl0ndg
dc+IljFl9qPg7cKb7D5cbu9n1apQou3V5+bXcoXtIG69zFzjJy8EqF7boEKA
DD+rCoiS231h5+R4kv0bscC4BfAd5345DpbXPj9sfj+yslq7sp7ezYDq7psN
eOCbc1y1kmFIFJqcasLjj8jSfD/+VVmm1FwzxW6cQk4vfS03qJq08kiIyF0j
SDPOtiKcI5PMTwXLTquP3H2A34YYIU9tE2y4mgguwwo9Wo5NJ3y6WA3v8qIY
2NPxPSjlc6Zvy8sMOvwqyTTjVxfNV2eWuowriDzOTLBsMfjCwdcGjZiMKGER
WE2xeiDdjL8AM1UzthfDlVR/t/14F7PtPw36X6dTK8ypmmL6D6lIaR+qLe46
j6V5NPf/beQyX5UnkygUwv4c4v2kRkj2d+EH/BNUqj3EjI0snmZTTqDzh10N
4BRmReBZUAmGVpyGXbildqaE/H514FeflKHZ95r8ZsK2FqJATkbgLtWJHb1B
uxdW23+E1RY8/vSlKCIEDnjKU7oY+ood5DJkR4c11fHAi5Xmy/puTMgr6s6O
siownbHYCGzzBf6d61Y74NPHULw2NxMEO/biGeBx7xSwcixfmD7ny0qVSnU5
lndK7748pfTYAasEYiR8EV5RG+L3O8YKRt/Pjf8x4k72EFHdOyIZT1kN664z
zm+vI5kxoWEPPwVqoCnI0hSaQb+sM+ICnK7nd9Py0+DVav7LDZ5Sz9wDZwE1
zPzRbUsiVcXKI0/7S5UIjkVLZzIJ3veuh/HfoaisbR4UFqpgIPRQhlverypV
db3sjjCk4KiVMFBXDxUnqE/eG7lz6cUS8gzSxT1EC8k0CDACEOJdOWn/GVKp
r0OGDgNX2tNO0euYV5bH/KDHvQxBKTLW1SMFVPIRJwfyzrSW/7vW2hEkVvmq
ySOj8VXpIHIBJVqxlXsVU1VyE7suzbECzigj5l4o9hAeUeypp/FKFp3JhLQD
3mD+i8DZb4SobgE6wdu9T12pwFOPOoY59JmdcqfpsdrVkIlwkQ8KSc311Ky0
nn8pxsFWy3uwoe9mVXoWXsJsUSLUgygyJNnYh9JIQLxrTHTj/SeTtYPdu9Nb
kI3wzAZqhMHnZ+HF+ItK2nCXNEdx7ag3kh6hTtkgr9bYxlUQXzGBxp8o+jJl
/DoKEWgZDbS2Kk5yNtQQlKFikKFiKGSHQf8l/GjDyS+X7rtWSsWU7rn/zJgJ
Qy60POZwadzQJtNRGWrxp2zrgsGFMlMRJJgL4KGePY0qjCbxnEs1FyLsO/pk
vAErLyLzZqqHoKU/5/2f7/cw/dIZvj9YGkarQXOmrJH5ZyC0UhVX/JZQgEx5
cuDAm2q9RqSUpY6xYJxzcoHj7rLF7JFHivedm7bADlRs/5BhywlKSQeSLKLm
BCLn/d79iI/BUq2abIynr/qK9LV/YEatBsY+Wy2r3J1IucYL9m7hLigG7XOU
t49I2iXv7H8MllR02PdRPK6Tu4vwwMdUJQJyRhss3OniPAhjd9X6T1PhJcBY
Je5PBvL6N804zUQ956XcbIlRtpjJLI2QO7nU2LrYmuKSihJv/3hF0G7DMg+g
eMV2O39VKsE+Y8kqjV+eOgKBMvNLbH5HaqMTm9uBBsfJF5OcvQHHRh84bnY/
RlN9w1dDMzGap9oNbCurOrtIPnTlTjHRYr1KAdfhNtIb65TBIZzyUiVktn4W
rbqHimDaHMgI9kStlV1kgEIXLaoSRGdrm1ACPSTYNPXsJ2b1HX5ryowVy578
yvev/M/sNnB2bvAdp+WehYIVdAYg8uRM2vCSaBVf6QhM1IL/y4inAbQUj4Xb
fAac9SpwgKrnCDsDpsfdqwMgYzthvgDoJJjTBEb2nSKXOh7MKJLH5I1pQoz/
Go20FAyW0gaqhRaLGUWxCc8ray2vgJzHLQS/Pioog+sPFoXY1LpTCSmK1pKJ
szvv5v+xwuxOgPTbd/OnZVwo1wn5G9U5fBnZ6IzG5aI9+GWcRKfHmEQBuDyK
0oIEyNDFI7WPKWdFEQTVtzuRZ7GBffQ2bH1VntlKhN5dZTrrVa9uKvjAwLBi
f0Ju8dM4RogpjRYZHCs4fLwkZt5w6YmLA570H4PuvfEBKyW5ELaM5Vsh5+0I
H03+HP4ak3g8hBzsCxKxhtkj3g7dwalQexLPJTkxQGQS0OJFFUnW3xepjgIt
IxT+ZKcTKSWj8/CKTq5TMZb/CTQo1SG2KUhidrF2Hetp2hrSSZF491FPkGm+
dsqN/beyVobYudYFdKDeppg0GqlRGFxQ9vz5bqhF8U2oxf53EFTAMovftR8k
BzKkimp+ZIBUFUYj9jvMFNbE13oA0lXoNkUIaqmBs9FeCsBDYBX72mFml01U
wAXZY7Tbi3V+b+rFOYRcWFxikZgzKJCLRnbnXxFmbWhPp4kJs4WjmyQBNmAS
Zt9yjRkpoMc+hVeq6y8EHrtPUBePP7jVe30+HUie9mEpx6apuQZdXuFi7N4b
2zJdrJrugcnU6JbrECPtKIPuhRyYR6/kitjtUcJxUfzY2+2OsG5WIVkZDkqx
Io1JEJjntDJnbDBwFsd9xpyE7+wLA/62JFEqzLFvRXCqwBjn2xp3kdN4MvhS
QDRGnvwKvuhFgT7SBP5C6BfhUptQi/+VuRcM9GOGxnl3DU/i7D9hc1uUmHWb
3MAHrvsEcZP7I1qdRwJFLkOc0k25CbgEK7LLTGuy6dDNOYVhTcsURXzbKFm6
drUfCpdG/phGcpJxgRJqtwepE3Mt0i13p6olhF8p4secOafRW5UBg4FX1Frc
abNEKgPhQJNIW/mGgw6xpUY88aQmfR6fIcindyoOg2IUBcwu4vxwo3xnzOBt
AgC43qrU+BeTgOp3I736M6FvgiXp+QN8HlPvsSLAOPfFbWskLgnnJmlu9/If
KmfOWTdYkLg8eyG8uqRQ2dqlVII0zRlkbQuZ8PjRpP4QO7zr349WY3z1gr5B
aL6mTZCNwt6ZnqVZ/uF50/GF3Zz3+SRZ8hlU6fR+IkyKgclXRB+A6qShRVHm
no6WBmQ8i76/wsFpisrA3llOa7GAA9drbSZbht7fFGojWjQom6g6E8z0ZZjq
W9ywOoeUyHAp6mogzfCQAqIBkVAV41kNzCRR8nz9jbkItBavIY4ZZ1+tc9ts
Zh6BW/9aRyyFPd40I7ZB4MBXW09KEyoQLx3jCs2lweQwvLuLj+eeQnbWk/C4
Q2e/05c3fR6gY8953leBogAktLhhKS4PKreQz/y1Xt9cvnFLC+QzmWXm8Eqd
vivg4s1FQB3ddr2uUCs0j1SOWyUlOJhEYNieE4RJoW7msyUz+Zugv3ayfh50
Sihdm93/4aAM/5YTzksAf914qmh7g/aSZK681TrfTUbOxRkwQjTBTxSV8eZ6
uyKd9ujtLNoufWjfWg4B85zqVAmbbK4zQWxHPmpe2L4UoPSmLywj9lQ6mWwd
1ooJg6JcnJUWPwvIuHZXnskqnBA+HEVfSbkFyp/wHZMXmZd3EAsRAdd2kwG1
bq+BuiLCe0+/AOZ6hS5fhMviRTjPEZ+NAsTdTiq/dpi3IUB37EXoyT+ex8Oq
jQ2mfHFRdWlefjUBehxOeY55RyYypfhBOYEZoaW4rqQdNeCo6gJpa7hnBpRI
sbzieNLfII3+S/CsKVGBbYFwQ02r9h5siB3iLODq5ffgxJn6vpd3QjLV7Iv8
n1K5ffPwDF9p/br6sFGV80hlhYE0+Ad4wScU681EJWHw/bi3z0Gm2+P4Z5yd
Q8W6exYTUTScf65jRRVZHUnAGrGy9zmkMaVPYl9RwARqiNhEHyAsOVA2vgpr
zuSGa5yGOlyrIBzEKebYykDFNuEsS9/I4/mt9mVEM/IOOLyCXKYu08Rym4BS
YpDcn6Ph5wpL8+P8BenYDguelKgFOQDp+DfEDklKPp795vxpK2+8Wy8rFRDj
WFPzv1j7d1kHw1wCM7tJY5KzdpsXZQleYGPHUrG/MQDJj4dvZMRVIyAQE/+O
dswUe/T5JatQPNIl/VP8gfItaYLkk/tDIKaef7S5O9TtQ5Vx8K1czYmHCUZy
TOjjFYw4uPWGX1CKRDPKXS0dAdWWhyky2Iw9ttbf+rSRz3xAKH2Jb5JYvyP5
SR7cwU7BHqzYlJl9nvEXY5Nv2VLb2tM4SDHrQZbr/Ctz2Cil2SHwhAhQV9WF
DtgQa+dC7ZUnV18cXltIyWrsqy3wfeAp7Cwmri9uOrst1H9uArorvox6bzUT
7PpR8GcWX/tfkKN9Fo3Unfkyy4upCULZNWc1Rs1FEmpbAa9cBwfThyTfQk+O
OKDGkqR9PcdWiRxo+Wh5/6YX6NucSNE0TtKCBpd6yNhkzrxmt496vad8Ep7n
MXMSQz8wbmuNrH6CSMCmMoRARor0ygVZ3EQYyye7D3ghlerOKGg5xhj4Mcrf
8LhVuwdWsmxkQxc4Dl8PrIseoH/zM2D/uDzlxEBzwlp8c3srP/DHdYELafSL
CBu+7yZeaBGrJp7jlcwH0FHnlmK5/7gP5r4onpbqunlrqGis18/ePJIwqqno
itHYWSXjng+muG/Js9kdvWhNzZjc7ArJ0h6U9drXMA5OX6XbR5zn9yMeLUHM
Upb/MEZUsVgUcwg9OtXndZDJ6L+whkdOPYq+gqmNqtIzOADkRpA6nwzuDbqH
+or4DgfyF4yAPS2NDMBibQ1EgpnSIhhQvcVy+IJomXWjoZdW90lC7PM+2r8i
c8KhDvp0OQrwgIzNZEdguT1AkhuMIG1ScrOFFeYmdQq1vbym8Z7nCG2Nhava
HyCAgFvDt7KPhWwAZwj+a7oOFpjm9p4iFO5lTkAZWnzz8pDtZOXN15T/5f0t
wAvV1iHuaUwdM00POPz1J7ji6Yk6u7snYqkX9Nt7Twu2dbzAltDeomCKO1hz
u7k1qhjGJuZcphDJ5VCmpCYMbnWdP6qqvXoiKArkEc2ze895ozGrgnOKMEus
iLbm9Xq84J+lEbBy077GwhgmDAxg3qzyhLPPKn251mEj7zN6hgDLHsTjvl+D
ZH4gS8uvDNvDam3H6Cph3EznqhSz5/4WrGWY1HDH3xbxMXhinDp/lQ10mAwv
EhmyvIGLIngsHvw26peXHzG8wP9MlTSFvbErICI9M7kN3Hnd/k9hnLajbtJI
DuPRCye2lwl+VxYNuxeB5C9Mlo3idwTsQzXGEwIsQSuO0CbahWMPaWwyQpOB
qbK0ihyEw7gua3PIOXjZq/u3D40IYElbW3emwNpK9XDF9T7YMAzNJd7j7Btg
TkASzW8VOaistfepH6duOBW/BbUtzh3/ylt8N6IaKbLmPXJHznEQRGMlpNnX
hwBbJLcFg6L5W0USLRb1ljt0I5j2BDImvKHKU1HRVfjiOzFUQS+C0O5cNhy7
gxkNQ4rnDCM/TtdiJi0gpTdh8xubeeDTMV3uA8C1SUCkDJ0Dc3pKkGA54HTE
5QtfPR8OKET7tfrQAqfKK5AJOAWu8AcZB1zlSw+rsGyJVAEx2MnprnNflig9
RPI1HNbPDgYezuYaYVo+Wh/lgeE7aYsiYLi6287dibuvVUlZAcEWvcIjfPtV
1OVRJuFYvnfP1oQQR4YaN937f0m1voIc5HMRVkxS/WRzelBDvS5Fg3vUVtwF
nmIKSuz9l/Cg/vxLl2lkAGLjvMdCaIiGoXfKkeaV/r4IzRD/+tZB0WMXKGB6
hAF1qjszbSuYXKVab8YGfQG50aE7adqw1MBTkqAG7qxiNFmoEdhT5T+83FiR
cHznLHpQ+KuCKqSOkeSzPb82NostB5QuQxmKe6Zlvq0ssj//kThgluFk7iI+
eBap1RAYwplZUpJWgY4AfR6gHZwSHjnXO0rMLZnadwklKmttnxdX9YIv6Ght
nvea/FSY297BcevlN/7YFWgBpUTWwlN9reynHN7aEJt9nrLLvgJ12xdoE5Rr
wKJJSu6E1KrplFqhAnPYBZWdl7jPZC32ZkF08KaTe0DuIGt9wE6NdQxD7YXf
uOgU6hmapRZzQVlbAUJ6E+LUTN7X/EzlIeaYuTGs2kWlYxrtKuF860qXDQcr
Fg+KmX3lOYlhSWaKt0FcgvoxMjW3ZYXNIdL+JtuMokSQR8XD2cmmg4BkYEyf
ryLWWTg8eON2QoYSJ1XTW5qeqAXoieWXmRvBrvxgZLMZNx6KfF9P6F3EvTj5
DWyj2kf5pU33DM20Ls5IPws55O8xO7rZBOevbdGEmWptYD8RfrHz16JC08ju
3SdBFO5OAffq+1RZHLtqMGV5hl3380ZV9rWS0PmbwHeF6XiUIWeUzFbM8byL
sz3O8aqXoIeOHRJjcey/bJmXhRE5FtXlhXiFwuHq6OxImvbODEKz51Gjulqi
dlNvJsUMixA08mwSRjWm9Qm0y0vI6DfN+puaNRfkFrZHtD1xN8ZlRqobxyYs
C5+JtDrNT1o3OTMY09oh2RV48730m9TSXrZPL9EKiHf2N/CJjZ6lYYBtFjQI
EPQmr4IS/WV1HDl1IcMwXAzC+DP27Hgrw8GY5D6LJTVql0umpF3n1+tAISyr
g1eBrr66eDDhu2W667cMDQHxZbwI+Hh6IFYHPmqS9EfpBVbNBTEGeky76GTV
OEp7XTJ9VX4Ykip1BgjF1orxSVOG7Xk4MUH9v5Qc1Gp1HssGWZTa8KQW9896
gwygt4b2VMB5jP8uZOI9nNv+DG82R9yOYN5kdk+GSDQHfU7j9b8P8HrzU2Xq
iV9AKy63P//X7k5miOlm6IO6kbsbvACuqH/rNkV0FtR5WvLcaHHmfgZP6hue
ay0l5mzlgcgKgjAUC//uEizNtTljItGM0xGWrfEkg7JH3FauYN4slW0C+IMY
EB5WgOZeJzx4/vV7arK/VHIFTeGuy5I+5yIMIXApnAGoo6qpSUnIIZyYrOu8
F7IH8xgWtwok674qtfjjkHTTmFS3qibqFVJf9OqWp0ucwQJC5MmtpSiKz5/8
cJ72H08uzkf/I02TgRqI4wFA7FMie+kgMuJtGYuhR5Or1ww5OJ3fA8oqqV5/
1JZFJ1MRw6WlYiw2rZLESkwP9KnDzOwWRisTiKkMNZZkAUiVZsD5s8/BrjWH
eAl7zfDYxZP7bZKXWmBx8aKiHUifs3uDHCXvJO0Rpgyydlnd8YpNiZpxfgqX
R77XCcDALe5N7sLcgZh7HLK4jPleo3lg+cQBsIgkRdmqykQ1ifO8+GHJNZ3+
Uhp1ZsJ3sMvBxpRSZKW7PiPswg7C+q1XYac2RNptmyrFhWwUd6JoOfwZoREN
xb0+rRTfkYfhOgialYnkpMtK6NwKIDkaXeQQLz8VEAHJ4/lFNGNdPP8zhJ8B
09NR5aigjIhhyVY6BDuV0p4S9HBd/7k4/GqwPff08BT1YvVT2oLysUWAseKU
KEquo4n4TF4aHe/5HmSPbfoD22yNIc0h8sE961lMl8w1U38Cg57yZG8ws9RF
3W1KEXJxtb128oTESCUhLCTkWfaIrj/PpsgsdKou+QrsJvIxf6G59otJ//4Z
83udZsEgJ7S8U7GaP6udC6/jZ5/vJIoMfGA1bjy226VCraq5H1DTL6LOYCQL
QGq/bapKeeDzQ3TAH0Chf6s8cTKd+yu9Md/TR9FfRYFq3zEkMY7ov2zRAHc0
wxxvo37U9jY3lnayaogqcgLDg0/aspmF3PDrOYe5qycSjutNBcabkX4Zf4eI
z53g/I1iWe4oJAXPYQf+OTLRr/d269oqaRvCntoSnJuwmKG6aq9Kbi11Zla0
n66v85aqH2//Nsjdr/TOSCV9zJjN3qdTlHT96uexaZOPsKTorZPAuoz/+mqy
nZgdruqsgVjUdTktjYCM0jU8R6tubkCrpd/2u5VqQW1irSplhXH4O/N2nxxP
Px2cGpm+RIxQOrmS7yYm84Hlf/sBh2J9mvKEOPmiNXvx+/mbQof/qqY59ctX
tccwNSqyJ2OoT9UdZq2DWmAxwG8bxHXYp16LrRb/jjn17eGeYEP2AkKuntHA
RA/A93t0gYw//jN2rhNbiNrDaxZ0/ulNLgC/H6W/xNADc9FGt9XZhdYCfTvX
6I1zr44s8Q9VegLxzEuGkQxLyUMEYUu6h0X5DBAKMeuD3F7+jkSWk6qwCKMa
m3HwymFGgF1+qY4E0JT44VUhsY7y5ITOs75Lx+RQblL4H/7ta4/X6XfHmxD1
wAFjc1vvB5WlpTf2ehEAvGKhNu7ebC61sYsY41hkJWn3LdjW+pzEty8u/0am
jPsE+wC3GjxcuhZP2+nfFa4UzpBwl8PjBvv08memPsn3qCMtXQOKnIe8EzIx
obz+YZKgcdQ1mPIBtAeITDqpqYQvZq+H5DYRkg4DHifn+su5JZTJG/x8R17v
awgIAsNNUDWF7BKZJkPbquuWyOKW9tko43Qkv8YH/HIkDs0rLZrYLRf3lca6
9PNkdnqcxjBvo9ItA/LWwv+Vb7swht0/pwDkpWLkzwaWHwzB4jdVI/o4sLlo
zeXp9hw4T+WueIWbQXQOqG+okW+2U8NzsLVS5jkwiLVEwKOOqe5+LwWfj5Ud
wL8zpNlHcinTiv0cdxBuCFyk7dc5SebYMB+4Lkq4er2Gfta656czVw9oASRq
/21S9G9PePws8XRl9A4hPzVExd5ZAlAvLqsoSilJI3epikuinAk2pfhfsKDx
UmHebpxVz2oAtPv6l5fweSqDZiEoLmNaxb2tCIWnE9AYzlyAmw6PIDbD0/8m
8nQmtP06Nwwstg2uT14qiI/oKbJGQl/S0nh8RLrKmWUnaXIMWIPGbZzvwhvA
8kntj/QSjYMKyUbgwKmRykMIiocsiyTG2wza5nRMf/4+SvtIgVBgQ6jtJ74Y
f2eTlfBcL8gOHeowzYGQExH5eDYO2E8kJnuQHKcFQf4bvvgPV4Is/c7vL5QW
KPJ0gDnlgUe9Q155COX/+7ExcYOxAEq8CQ1URm8O5ZUBvRB+/VQdTIMI3ELi
q8VlaFp2Tck1JFISzrOjCQnJzgb/jFPFsmR3IQsBwRqGmwVjftg+9ZFIYTAe
xX2W5fnBtGYPCMErmD4k3FzrFllB65cI5htYuURvSFFdDhV21Hc4Xbd9H37S
DZDi5pDLJR+AhfmuJv3gFGfJulEIyT21j4LRs5eyE8rBr71re32ZZB8lO1tP
AaeLIDm560nRiFydpdMiTED2SSRU/2ltKAZIPZuOJWMIWiRFlzH6Ws025Xm+
YuEr5pSvAcFZ/EBFAuCAdjUFQ34fPnXs+Jj3867MSM/q+zovu/MlLMpOZGmw
RHOzjsoFUUY9djm9Qr8fZaUlmfxEFiSBfGgOJhUP+AwgDa4p6S9dTbHmu9YF
O5pAcuYO0xVkeQZUV3l42y75u3ldZS/05R6+xo0ixFYrZhLX+DkCucGEcUlY
wY4bV0P2L+YcY+Og2jD5ZjQVanzLkc65NksfM2cW3CEEkNMJ2DY+OaeR7zlC
/8PFyk+r6/P/t75lSjwc6Qf3V2JsbSaE73C8QuuMWJbmABMWlE8qZV2D2Gvt
y/1riwW0+OEUMVq70fktpFlb7schcD8UX6oqxP9p4mtozcLrE0987r2H3TPD
oug1rWGlTqDbb0wRPGAFeC5jzo3cN2eGYatkHNM3FPE+hDu+OxAF/I/WH1TJ
Poi852q38GLff14ud4whMnzf7KH8pXRdDmKGgRqw88qFesCyiFSw59gIKwyU
042DATJ6pksv1SnZ3tOMUu8airyJ0WcRFwbRT0sahmY+3NPt7cjlXeY51yC/
5pfpLb8RD7CJ1A8fDTe560AW6og9+Yl7z3mJ2xklvStU08Xk0liATt9UVa93
H5ri/ipEel+SwZ4fllnCC4FkP2wiW8I1EMN01XiVmdX/6yq8WFY8Dp2DGYKy
K9sK9sYbrI8Cv8sODPvdnUJQmEjVC51/Tcnu2h/txfU3Swtn9+x9aQwJav/Q
EKyC0Yx2fRYm+YeXlhLvxA1/Eov1bem2f9YZVnVfqyOALvOG2PW2BxhNgEp4
Z0wauqFBzJ0kCRoOIZlWJu6DTxgZqrLoAMmq+Vev2RxjlAIXDcBFBfDgQ92l
9GUVEE1wnJYWZbONJdNJl+LwMV43lIvgh7AaMWi0nzvvW+/07kVO+9t7p+qJ
D8B1xkry5aCs+8hXGoIo+tMq60hh4FWeFQ0GKsIOowGbqS/O+/vMrAAgxfE0
tsD67dM0uFDB1WciUNaTJtKueH3XxsZ9xDPPq0iaAZg476h3eJHOJCtwl/wj
AvkhjpBjMsOf+Uw9sKi0MPjGlyb+S2GYsQTtOE/T5Rr2YcWp89CtJSPm/W+T
JuGHVQl89iazmev0FqN26uakAvCP7ngA8MCKQMV3zRTWthASGq5Aj6gw9fMw
H84OfeiizqqjcmjA4Tjt23YPx/ci2vTjRMrQNt4eYRTQuc1L6WEo/wggGhhu
Ips85vL0tCZtCVAUV9Jh0jWayHdDFVzRIKrLcD/VJyDUSKN1ZcElLvtAPDEH
tY+He518JRhcQhYdDGB0BYqSWnVRrbvcE30TZKNGJo2X9OOkV6UqteKX1m0p
RtrmWewL1Kg7GDsbelV+atsJB1WJ7DAAadfdQqRiQa8NEpoikPI7qUcxGM6D
FyROpD68/1tSnpb67kfbdRAggmVMXM/U0WARgYo7KN/UMLEnJFq9/voG511k
bbiufZw8e9QBKoTpJ8mtdFdhoiSRuS8/Ou2u+9sek+WhSFC5P8xxaFQrjSla
fSxY3t4e1E9R1SyP6tSP30Va7Fx1JcQxNuXt1f3bKBSdkJLx/TgnlD4Riprv
8gxZ28/x5sg3rycuRFrpVckoOKjO96XNtkGMHVdReY8jTFRx328kl2RbS96K
Ihp7R/wRn6sTCZXQypEArGYN9ykcC8aWVx4sEa0Yo+LIXC80fYfz84Suq7Ni
4oMC6uk4s3pFprXsbJGToDcfeTiLGJaoLBufmOpgjWhJVSUnWd2O7icoCXZe
03lz/dEUtrZ9A4rWlaD9akS+AEbIWJGJrQT64bpEO5FCjqvXjICFFQNIE6fV
rcoKj3hbuiqFt777cMNQNDNdu/l4KL8j2d5+mkqfnuNwfH8cpk5F7G7SxfI7
LqTeESqWmr4ukj484oWhNTmmguSilhVATvbG5TGEsHjiE5BJ2CQ/EYxvvj05
8FcgzHffvna1w4iNvF2nFXKL8argwXAfc673wFRPvfD0yHZyHosNhH7yAcQA
9cLF6vV9j3BrTtOVdKezb5Omuq1XAzIzFMZuxGk9/xLChP+fZl1ptUvtEGYD
hutXfFPeW+25wEitV85iUkGvg7v12d3VaK/esqZm4E9c1jQfHo5FVLT0buVY
kmg9A3HmjDAUKFCM6fhcfUjwfOuvTI6dVbHVNgu3V98o/GkeTSipdcHTqgm9
50R9gS2Lj37u6NRAKYSolfM3WjGTZKl+NDlI2ri3R+AMVHtW1T5GPuv5qsjk
ACS39wRGtvlNuoeTQlgT01taF6+ln6q9e0n27f0Zp3I0Xolb8pHm0v6Cd3+r
V5z0aJru/oBmqj92SLBOyBzL1EySu9lUZwvEGOf9HL+iA4Ia+pi6/46E+xZa
bqgFjotApWjbY6OB0vtsmNXebzfl1591vmyWdu5M6qaGM9s1t6Qjp6NeGCF1
ROdpRC5Nz7kQj6l2rI+5qQAYaUMXN4a/V/eY35WWmqYS8RMVFrXpmahcShFw
2yjBBFMsDfmPE2U1uNGNzI/vs/l78NJIFeBHtXK5LfCAwF532Nt3NBV3SJO+
6gobpD7X5/hPpqwI8UPgt4CRz8wTNyakJKmMhfuFm0s19683yvbajdyOVhSW
jPzZRJYGnYT2jATayikwGLa+lFFBmbRxpvlstmRPQRerpUa4/E57lRT8DX8z
NIkWdxAHRIDt5qVhdO8BjQEDLAzi1OO6kwJYPFGOK4uczMbn6SmnDMYtVu5R
1It50wmwPwTnuKko6dNs7MOdny2c/IDCfv5HLGB/xmsw9lhu9UQqoGRIzYlI
ceHii1LpUivwblCPT2Iyl8fJTMh6v7ntHx/nohGRQwse/XgHmn715MEkTzs1
ux38A71reg94y9Va6txC5bc/C1TiWOnC4fB2KI+dBYZPZJyGsVFeNtFDYq97
3Cnb9JldOOPtBRN0tRLv7FE3MNrdr5sMpnE45lmjKnmYtcVgNOJ6fPERpsM0
r7T5zU16B12wn++KZ3gqfWUGQTkipi4JzBJ2jKRouqpMPjW90Bce4A0DBSOy
5V3KhsNZIUKpea7JRU9mYriZjmIJXT9D5kLDvMSk+C5G1qOWWP5y+Gj9eWrv
nvCKPD/YJUjuu9DCB5Nw927QbjYIHCzTmvWoFk2B7Jv56gkfhs+dkoVTR7pB
9GHebB5KYPXXGwZnbe9VQ+TBgqkcdWd9mKUPydcl/jHeTqBN0jckDG12j9lD
wh/VIHsL7Q8we/Bqvy5gpztZ3WnIwWFa0Ha2XRVZnhNbWp7mKOrKNS5Zf6Z1
TnY5jcGtI1x0yHnOA6v1hy1eRATnmUTvyngnFGirZ4yWSbbao3A2IbSWLPxe
nC/kr10Hz1oPPuV4qz6xiZ9hQnX6EbVeM6Cwfw2ITichzrQ09aH1AGsG8bea
BPDqpi9031T9/8wgUPL3IoddAXRQZhXPf7XtSxo5AZjRmXm8SSvt2fDNx4nz
WsnJFKgBXwgvvUsghqB7xSIvNkap2xRj96A4xcSerCYqb+tTCmKxZPgFhFH3
JsdQLTyI2GDLSxoiKwQ49DRpUK7LGH5f6oW5d4Zl5uD4xlWMjqj/n/RQPSOu
RvZ5XeufLGPW8G8UyADZb7wrGnmP2T1qfI6QdwKhrf/5S03QAPiy663WTd1V
D4Dtzq7BDlNdKN5P8KXCSc5LMzcl8aIMXo1U7N1ormiyxGhOahUf7HuiqO1d
1loJaenhZR9EZ+8y4lypTooj6ZsrhZYceaG1NBddYl0fS6KpN7CVNGxjXjf9
jgwqqf3npNE7BndKlQ5P+Bb+Yu5y+QV/e6UxHNWpsZiJwGERLQrMT/BLLeOx
LzEX5+OlTauHH1nyhyP1vyUoGrioN4lVgdXFmYe5tYZBJvY4U+7n0LyoQC1e
vHzOgFf6fBK0HH/GeUL/KFQ9r8f3CDl6+SiDmNfVUpnSVxaeOde6hw+4crSo
lu6bjz0tPQYhj9Y2ElR6ho0PQ7Vii0RN7S0M6NnnI0ySgzw/xDj6snbtigbE
WBjDvzvwvEliT/lPCr89rpCi34LQUBYv6jg7Crnj7bCrIiTTEu7YVg3Ey6Fh
72Lq6F23U2BAt1VtCFJSLk6R6Mj+Hx5k9ujWttFzljrtw6CfrXlCXRkY+zBi
Mre6khA+7gmWtvXCK581i85XwQ9JdO5YmE7G7s7b+Icypry5oN48wjXlqQ52
Se1kb1KYKCJjBV1pLaBKFUg+Vt64A0Rr6W53MaZMyY+xYckVmf8xzK39usPt
ciO1UwtkpAJ04TFtfkTqQoOkWCAVZ5BuoJIyaRh4brsRk8fsoKnOc3U1o8X3
UZbQM4XAQtaYojRDMOTV3p2SesORNGQ6257sNppK8ZpdcfyXIdLe+r15yaOz
0BqwfDcdnJ5OytTHXUcwGR1QQLw0KVH5Ck+HLTwUxaKkTLH/I7xzyy9uQR32
TH2zg10g8XTdIwjw573D5Gn1D71/RU+Ztfgvdz35E3X7wvEnHwvZF8W7iLok
Wd/lIH7Ag+h8OPgo8qyTOeKxp/jqmBnkcBoJ586u4Mi7pkey173cDdsZzJKF
+yI1N6gNYUgo/rKBx8KtMK5dODCFFB3HBDyJQAMEAd54eSfult9pnP5uardO
9qL3j34q/iK/C41PQuv6I6tQres4IpZ5eUCxEXY8zFrj2fNIc79FEgk5O+0O
+d1GVwSi8a5k10a9T53F5jEuFZVt0NtEmEqYlONgMkCXAOx0zSy4PCJ4OZq+
Q+2hytoxWmAXT5IYF8d3ULx0HSzOqYYM1nHVJHetozLs0/kxSDEFoIIQzHyz
474s5ClbSYvr//mN+eBx6k8Rgw1xuhAVDroWxdgi6dnb5DzVDtjmHLQJt/6f
xDzt+KaG6CsyfQ1QnR+OcbSezxgAb85OGmp6EwCeuj+UVlqqDDw7Tn1BXjyA
2NzPF4G+lMXLYlSINFgt2ASoTeIYeWVGr+/hxUkmRu7o3kr29cYy5/gPoZ1j
d7FCJj7Fn7y44JTXx3Tjxlmr9kT0t95rLem+XvYjzeAfjBuZOibBqOHhpq1E
nZyYlmxIPv7quWjL9sP4iYNKEW4Om6jItMUjINCZTrtZnyO+ylznXoVkbYEk
Cx7Yao6P6SFKt+XKQ3bjgUkmkDQkTpRKHWnD6+z5zfhDRRT9ysQLxhCg+ka4
5roIidp0C1F0UwHeH2INpZJtSceJbFjv2a3/r06Ls8ep/hEvHMTFngCsU/7S
SYGOe+vO4hs3DXjz3YtFaTd+VqRnxoviV2YcOhC2QKoygxhmzLzWAYjpsr2S
uhm1U70GPip8dUidXKlclz5MA1F0kgwtYPtEjgf9FcSnmo0TffQNDasT3WnX
/Z99bcLe1ZbZlzoEGFyVaQbmEibKzLbIVDkyaKJqE7w1wjIXBwkQKndGlaWh
ej+z0jSfAGabZ2dl/drGlPuqZdOO087KheDfKt7PJQ7fXfRExFyaRByEZ4H9
9p+i2sc71ll9ntCCm1sNjPvpMgkNJALwsAigS5ZxqCMZ+u7U7IdSyrB/ONNw
HbHvjA3SCrMyYctzMhYrwJpsXf1eFCGB7kQpYZzWlUeOiLqr3mgBC8r4bWZV
rx5cX7x3GykxJk/ehTsp5cPx+Htv0Cw0kLV7nhMVY0OXJqg7OnDNsHJ9ri3M
KT//JXK2ugDkbd9B06aQGfWGJl3u6Vh8UsOZX+0vDFaZQKCLgn1FB1ybbKQi
ghI7Oxv2B9jUL5Q/qPQK/fsoMIUBgqWgSXRXV8y6K4C1C41FhxQc/tHvZbJV
w1a7tOp+pQGKq6f1vArSBtk3D5W68YOJWfz962ka9PZtzzjulM9/up7NmpGz
uQzLfpT4DKEGAkiRTltWjHXni4xazMJdfHYJAUuzr/W8cl2AKz+Bwag6RcjQ
Jl0pKwm7ibLZI86diYbxixFYkz8ISjZN4nOVpXxVGvf0qjE8Nqb3joJX+InU
0ZOIy3wXI96+yTOJUAXffyC1RABHEbfeNsHDvqSnWpR2e4nrCRKBaM6DESFN
VZ7sWQ/zSm+59zoN2lyzYilZmCYwTs3o9WUujTCUlvulqS4ECiD7pgE3IjXM
5jBXoXCYZJtMwzE9nkYOs1oS+4YOYMdSk1AoBZrLKJjGkEM8lozHEhEBrkFY
riprgxQv02Hsmfu+EfGhqMFwsQYzxRSu+PEsQv8ZJ1l6KOtxrb4/LUSm7ZXa
ScI5hr8j1M6a1A0MiZplJ7vELamtSm1AL19unAUWb3sZBw7I/m/dIh6Y9B23
/zB77qJ0K5RD+e7VpsUUr+z4oQTDwIUIqP+ZY3RaAbCRdj5rUHWXRI/oyjc7
eGhV01nwkwsrM4XJH9/5M1GWJuhIiSFAWrGpHWzqCIxatEV9MBQhCw4abKD/
kQjXqQHekAtGNdpJPRTgnCZUWD+anpnjteUQ91cuLWBL05g1Ut4DxR2CbMUn
C8mJy2oubBjsYR9Y2f/vHXqUnIHM8pxWNR1XuB+wp13nYINpRh37i0laCxNs
xGKyKSF3hjw+Gw/zFB95/EexMEc6cBsE1MsXEWq9ZNhdnJqZncGR5mruRvtw
KtNYidz3Sn4KViA0WHAA4Xh6bj/9UeTK9V3OK4nK/LzppUiJl41u3nr5yAAj
i0BYHw0m49+xyqzeuO8rkVDnKNVKWBdl4agjJ+kC/kdyfT8C91jZ3Kr/f86X
aE4UZzbsfd3EQebY5G19nq9xCR8G0uWpA/TPIgOMB7TRSk8PEvCwAcCeo0WV
zY2QvaKcfCjzPcenFFlisuL4xTSXotWeGdS2Hh9Ws2ArhrfWAkRhTJQG+SSR
90t0IT2Z9N/VkJ4IJtq9Y3TSRtlDDsKKWWBMjbpUEePliGQjuC9hLpBzyW5E
1TMoL3AjvyA67KwVPDwtUSmzBXms3qwzSZN7/gWuBw7sphFKr4Bvl3yv75lM
GsjuEz/v3yKfgHRUQdQo2lFiHU9e8smUVgWTsqQtkDoIkqmdBNOPfUVUAxc2
5gu6+iAgSEo83hm5BwSmbAg1fLArn7rb2i6SM7Rk1piCc0GQA/UdIUyFqPJ2
Fjn25tFHWWSAi2KIAL4OX5glXDPFiXd4+Z+NnGu56kbfywc9wSrWEMuIrNmN
EckXtlfUW1f0HsnAdY8hkOKNsY/12m3/5eJ2dRD+HqppWQUon26mJ6zEEdT+
DLKA+8PN6MJQ0pllIgyG0fOwEYe8UtFJL9X54ixOMqXI16kO+1x13W44rfxu
q6w1CKcEDEE6pKCrhlILoSsBVblRTOfu6ktvrAQiVofG6e3c2J2QIWWRm4EC
QZ+rAn693FxeNzeEOa1HeYwsNfIh6f7MFDDgk1xIPTP/MemDjwKPwmyrR2pr
tBtOJ+MmoiIY5n1qDkDASNo9fGxqUeHsBtadqI4wPj4Hz/tzSPzDJC3zNqbD
89AsHy2GHUbG9Sg3KZYuOdnbH/DXH63YUdrfGN2YPg9RZBVhYRulmpIAbRCm
yrQMwUrNHBW27HW3gu9SCfLmt1yk2TS9Upw9eZrsI/VGtzt8blUYMzf+UYxO
GRIMFR96GktaoDOp2ywu+EYAynkVw5b76uK0kgP6Jy1AHVTZLv8OhHwpRpNA
3fFMUxuS1uA54vNm6uHdgwMWXpTd7gpKgeYwge11hUddBHG4w8IzRRB39QyO
eBsbv2hm7fQ6HYoO0WW14nFjooEccuxIU3kFxyDW0Zp8oB5pzCPGQuliPmpa
HmuzYDYD4CqQKgdDB0f81p0qIEGht4P7t+NxyWoOW8oO1g0XjHrZgpEWsY4M
JGRk3cVtzU0N/dWlDuypEXC9hqGVDBmSLr4zBpaToewan/h+bXS9NNi+31bZ
nzeOnqmiF8Lp/LeNba3yfLV6iCKFjLpxOywg4UV65QEu+ECfwXTdDfAZOeC4
hmKQ1fV5QMrmzxe/Yh5vnGfV5/e52L6iRr/PF+43dhsBTm7uo9JN+yqJ5qHY
Lfy0XfYkl7/8fCbSsUePgeCHoQ/ml/sU2vQzXL0SS1VFKrF3s4Mu7H/KCLCj
LQ8XAfzY9E96FZkwTCFDiiIcMMB56/2TnmRnCkbhgc7tSSoHZAntGYFFyamO
4dVZ4ZyOyXZXUEIoZiOnCMb9KSk0EoD7TzC5+AgQxJGCriHz0YoYGwOjOMUO
jprFHKx1HcSQTvxyaOfKf+HguOU/N0iKPt3OKXBrO9wHDjHK/QQ5D00JwwgT
++0h3XIJb0qbXbxHAubjRdIZl0UR6OM0h2TfGQnw0vVifBrVQTvFjjhajt+r
A/9HX1MGV+XcHBWzBxzAeYRVdnYkgDzG3RRyY8JCpAHfndjjV1oO1NbFn8Bu
fYVF6AmkOUHQVW6OdlWqpuYZDgh3qs9xTr60IiA83rb3XqAhnAMgkrGMHKQ1
UnEWxZPphdl4cpFW3yNosnT/Cd/VkEcPkHWUmvT1rp1DjSGSmd1vl4klS+Zi
Go68DtoddlWYDH9B1rj8HiWwJUFfkBy7fi8q826hTMd/mPNTvIYzu33eIxhA
k5Fri+I4JgEVSnwXzh6jbH5uwjYH45qtfJfbQd9ChphugrcR8XQ2bP7jBtHj
h1H+28B3ICSkMfMasooMYlyC7mrKLGrFRMRBajpegHRqHjFT8X28pcgSadmh
YmNGUcnkMi8iIYjhMb5xQCAfd+TAWmuXZ7/8SRplwmpkM78CYvqcuhC61Zcq
+AN5dXFXBPNExVxze43yjqdb54PTtNb1Medve8zdRzmEk7KGGy28fHU/0139
DukQzCRZ+9E3+L+nLIdAuC56TAWQTi7vqqsRZ+LM+gkfjD5silekTBIumKKr
C6BAtaN53MykN5u9L2lqbska4BvPK8LQj8cK9NboBHFl8Fpg5z5ar6vxDy1v
JdUsZ/FZZa1vrFX/PxIj2uZIQ8RrNePkA2ywjcwXfWk1UIOymQXfq4DpuoSF
JTW8b7YeaC6QJdGM/bz3K5/mTyaVlQ6V+XvPsjSlIJqr+5Yizjw1M93LzpGF
AqDYIwHnWxAvMruceHpbt9UAvE+CqmVLkeW6aXc6vrcsFV5bozNzVSSW7DzT
ZpX7oCnbLjHAYiTAOFtAMNrM+7HjRA5VWkY+qaxcadXzriuHp23RgSkDnm/b
D4ihwgRc3z1+CuEx/DwX/s2LpHj1r01UI1NvVIfZ/9xwYu3evvxwOoSr+817
Ok8oMqxs6by7bLUDsGm9QkLgeMwe5y4m/oSBLE2dsKNPZDWCkYSqy/JETbwk
9Tbs8L6djm+8pcExRGD9ukIsIB1K35NkOnLgJ9RFtwpIzhIkIzO77XAKNfoz
8IT4m77+L0UzW0Zo7tSPB1UnRy128uCQS82QPm7pOPdjXS3/TGR6hWKGbEMb
hQtOA/v/uDU7ygRLT0UgNYdM7ioVCzao9tY70lkoYQECFg0Mfpd69+dbqzHg
126ArCI+flZekp9vgJDJq8jZ+zkE8Ay238m4+1oCfrgeSsp29G7rgmd4ctCF
EoVH5e7mtei8+0Pp2eJMBhwzoSxlHzsbGgjMiZBc1ijeZRGgwSK1TE3hlp3y
3U80aMjpM3gqupnVvbs695/WKaJT1a8ZVE7CEvwtArJ2ddymRDLjZtgG/Puc
7bbDzgQgA8iAlY+4nKBxkkn8g/68wRaZMELQEe7aEFEQ+LBxrjK4+R9UT3rF
1X0k2EsoTNS0X0Ta825NHYvKbj0fXEqfv3/Wmiz5gvuSh98yGrtetNZyeSMH
klhfWYTe+tVfRxpsE+z3Soq6HWxTIbQC4JqMJa/onRfVMvyaZRAV9ZWdlwGi
dmCftcJCm0Ofeme1SqA7qbJd0kfYyt2UUceOjgvKQv+c+3XFfED6dcaYeLf1
ZRJh+MUs0m6z/Ih7LgdYrKLR9R6Xnp9Nul//Axg4W2r6BMLWTSGpSH0CtDQX
N1VS6l5Ravqw52ipqJFT2nzTCbnAz298LZMG60nUs0jIyiilH6lVWgm1QEcV
uCWJ7md/xDEsZdn4UoUNoDsdSN9HQZGU61p07IHvLjWeVil/MJCRnJHrl1Nv
2dHjMQTrM4IYOUVkUoYCSDSDj5uykmHF12pOTGc+IbGmuYRKDnL03sqDvqVm
5Mq2K3ojN8fkHXYmDBhe2jV53l3FkbudY6JR2ppD2zWr+LW0HW66/6WMxeFQ
yvtYYQxM8xgHiZeFjQrp+UwYWCbN7+kNbil1z6bapiFRAjZs6nEqn+lZkOSs
JnceHJMuwrMYJoW5u9F2MX74cizNFEanpEUHvxQerhr6sfIiKnAYAeXyX/cf
ZmE98ToHEfgDKqn7lMuj+bOXogitZPwCglVTUXHwapss5GY+P3satLJTxogM
JwEB5Bhi9ANhRplqxrRYjQzzsoajab71UJHKxoBDVIj8BnutxJXDQzXst5F+
SwJv6qGQ2ydY9fXvxsxVZgWoj0Cr9osRpg+wHaxkqeZBD0bfdJQ6mIjjV4Fq
4PqKjna1zQK5Slv8tQwHU5inlMF0UmRRLeQMV0zlmdM2YH4QarmgczRRbaMd
uEfWaGDbZv1o1pSECiC2BFRZO5irttAUfdkFc9LdBotUHF/kBZXac1c+TmDi
rYybabTheMy7iblH8fvJ97fu0D8D55hYu/4YSY8Sh49PLS6mRq65pSfwOlbC
IxxjLXR09AK39xjMuXTPlm9qD7m6R0uDt7ck5k+P3o7brpiip43VjNp8ebG6
MEGu+/3VYGyj+NzMZ1Qv5uXCJz4nPiHhx9E24ieXmXkWmOav69710TVbYLPK
T0OtcSY8ASC6pnzsHeN/uiGsDc3b0quvjlfDTkEJ/1uP76PJk6a4eOgbPGpz
aypHNkMVV7A3pWh9at2wNeWszsCa27kyQHhE18jWzZ/q6Wnfl+3UWXwafcno
dQ6BHe0+ktb4fkr2zB4+Fmaw6ZBQHwK1oXa+9dF6KFyCZGQKi6w8FkG2DKet
wGy7S3/NT4OzWsOBPcezLcC1Fv83RcEPcVDcPPJISlypLLmXF6QIx26kqYI5
rF+OUSFtUfbZD611xW4CHnbUwIxfeoJlPl4TcUVHz/6ovjY+m3UV30EjCgNM
haISA72hWlkXUZ3tu0lo9XxCtY0cK1K5UDvl8uwIWGh5dFWeLgvigKlKM+9x
GvZktWW9Wp6xSTVNHxQxWkStE5tFrAKg3pCh/fQMTc1Z/0CzdQC1icWxWFBF
Gtzas0eoILKTv/KigA3s20v93LISw5YiLsnLjU5M4QhfWV3lz9gmRFxP/Xdh
k14jov8bHnz1eav9Gb08INpWPyQiiKfsaaE4IH+2QNbKSCXIlSxcqm8ji+qO
0uD8btPYhBu9GO1jNHeVmzsw9T9ScWXEaF62cpN/fVFCLSVVFEp3twYzBr1S
gTRXafMsVYJfcNQ9XRvH83Kv/sGYx122IKs/5ktcBSvrsZN3qc5sja8ms6Jz
ih7YlGE6ygVClVrmAgc5cJgubihUC6M5e70QDXjFe/37IMTiSceny1dyfKD7
v8do9aGW+rVv2BiSAJN/P2e0TeoPJ66t+oi0rjJRhFONh9lkkQWeXy8bt6cM
Bmf15dw7Ybm3ZNcASgZilnr8w+4xSDwoYK+fH0DqUAAZhbtXkklgVp1FrBwP
he0I7YG/JAOuyXyHovHxuo4PDqK+ZHRlpYNNjFRrQZx+dHr2/THqYRlPLxLG
wBuAcEWU6F0sOTb9tkfOSotFljUhoaKs+j8t1ruXb/7ot5nrD9pPsaQec3Gk
Q53kBkzidXgY/sDUsTiMDS+rzT+34y8qRRNvMBzlONisAyAypK+Fn8PR7vjV
W/7guYWu1DW9hlmK681lGrT3zddNc5aCvWpWSrJQulMmEHtbCzqKDaEnuVy3
W7psBMAhTm29PrAzDT0VW1j9BqdK5T2J8xs42lX/bCwWyt/k0RQbXuTTwxjY
77jkDQRveGn48iyRv1B0/zTNxggvZj//O3DAPD0/7a5287lsB14jhviBlXLI
63e8W9ckZA5oYQKxCg98SCiWAyE7V3MIFzCCKFbzg2EAMT2P1sMdxh3uB/7x
/bLdCz26W8n+AGzMf4SXyNmJbvtHLrYjbXUc2+cy5rkie2HvhluYqg0zjsbo
73JE+lVwOGo/E24WYq5xzEfG1ihHG6smqKGElITEK74SpZlGs23BdxsUxpEe
fU30OsmlWKDCQXYyhpHtHZgU4vkvnFV2YNzIfGbJ4g6YLJlLJt1epbGUZKEo
B73IPPtuRqLrpu6NJcB0DUV/uQ0ztJrsROaumEt1GJKgzXcVBmtp6aJpxbDf
JQ6W+HPbAA7RFqVYWUZPkJXPmgElgbC6q9uWg1bviweee/o2TSNrJVwb/Ruv
kTXOUz9YbGI1irddRMMB/NXFo98fva/rFVwJXK+hCTpoJ2QEC4QbjWGlBhKT
71WNTJ/IFMSsygFFUBaSOODPCKSL4JGBfvdp43uKlzTxSXaugNKqtviAN8p3
OB7q6b6DqZb2R1xTnPxZyz+ib+5gX+w1mWlxgjxOzcgB1MKXB1Eh5brCjvAx
4bPU0Rwz+jnPNFqC6ZQs/BIv5q1x/6LCh/hO1HEmEu34dXEjkk6ogJI+yO5Z
jcU5X1LP3WwuyxTxf2CsShzGc9Cd62GdAq3hDVbc0kOwQrLcF1vVnVfk+Ah0
iQY/DpUgtLnClQ0V9qyRb4V57grobP//LEwVjfaLkoM6z4SNuLWtDnBzzKoc
fMLtS/dUjJdz5JYEnCfW5Z5iBYWP1+gSeLDy83f0D8DIoSZj40rAvhq/XgiN
xJoFGk4km2TIMGfVJy/8q2EUBWEDcOiV7g3STIVmM+MBhbQJIYbgkxKs2SqU
m4VBzZveoTZG/2vJhI1RfE4K2Tw+ri3/FzUmsEajjnvlfTqMfHPIXhKQDfNA
+p8Naipbl8BSXynuvFLr0z+TwydXJkahm1oooAHiuU6vOSA3hQnrboaBFeiM
CbKmdik3SkvrrVumMwfFf5SagEZQN/QFWtyI5E6rp85rWBIaO6yJ5beQKIXg
AOYhNW2E89xVNaghYcZ/csTvv5kElMeZZnozXs8TGshfOkeLzxMcfA/pxV/Y
KDwc7HwTbE1v2kLimEvcIRr46nXdt5ti0TB29o26wF5NuoMbSWCbIPm0z8bB
d2p3BmHAwPRLr4eiaaINBlklatqMclQrvLlMV93H0bw3chYmGp73ARwV8xVZ
momDZ6r9lXRxSO8LwSEkCEpUqcE74/J1BkXJGWNOZ/CVPgcQTP3U6TQVhyBU
07tUKrWe0T4Ibmy/H1aIwjJAm+s3MC+iRpGl871oXZLVP8DLMyqfpPdLOpO8
MVkjFFy2OYpoduLerzkBCw3xVPrXvhFz1N+BPRrMSMExyH99sQ3y/Cva68Hb
3PRCCAtKUVgrZKfRgs+xM9lQEYyaJwXu/pXBOCSgMp3TJSyjMSM3R4kDkdT3
hzRl2qVYJi/owCeEgOOs4rUrVSp9UdclHq5Pi9aucBqp2JvEdgrofxIxrObL
TJda9eoVSpAQxN+EzDIEjXgXpF9tKDGdQDgq7nVoPOuxBjriwoYKg/2MxMEU
X8/EkM+DKwow9wXIYFf2pYrlnri5bpjHIZOJtERJZMzqVehmG9vTweNBE8Ie
qJXV4G9YnXdj4nAIJH9CuvWIZKIyHjNtKFnIFZT9CDDqkJSXwhe2vRQF38Py
l/WU8eDJcUJaUHpFDhpqaisEc0sBAv2YKQGkcl3H3qlW6u7RgVf9717LiriF
axJN3GZwAi/Um3Kwoab3n5NVmlHiatYZNFKwwZwjM16HXEnmqrFSVTxgAPqZ
QhbcfEyCwH6L3PLP2vx9bazQXBju9+6iSra6zUCPuhJ+2VwHaRWmoS9zk1dk
vgX5e6IA9Hk5D/GYkdoGigr2zqvvgMGwxw2amYXD1UIdebMHbhcK5YLk8I/G
Q96CFOstnSzHQO3Dtg36/vY2PW75eMi2lGpCBUsxngfWQf56OfukQuM0tNCd
oSxBpakjscR6MX6XNoz0UTcD0BSX1m53iVlOgZj51MnHSN8nGJm38Sd0zPtp
1vpHXkJiGI9fXyW8ijxYqR4hvcZ3/cdgmUn/+sljPc8OY2r7KK49/KAmUYSm
BXt301j6YU0OshKs4YBlL1u2BkgoEQFCRmpZGfULUqQdcYCPG3lwGbcGAqf5
C5WT7e0VZkBEOXHVd3VgY1+BJKynDg0CuBJzxuzlKaLisNaAOkK/GEV1Pz3x
IOtjwBUh63tKUfxn9VJARcov6t5BVaXe/tckmWuATcVDdWmBWcAIUKrPESL0
UKsdcC+rkJoTcE1MStskyXqVp/jsUn/DWDppXONU8fa0ghKWoljTtY/wxYMf
ewE1JenjpAi47K1nVDXhAXPxZ72AnAVuIeOsomS3fAJOGDnoZq4Y0+vgaztB
3J/NJih7/aE94MnUejKeGlfdxSBfFeb4Nv9mxROfB8VuK2hFGZS7W9D514tE
iyM/uKy/Rw8CSFBAig7Gtni1zWO8W+MVsGkdWwhtvJFUqnV4cBOBrqyxyNgD
h+lW/lun8SFIDtgqSaauq8Ty21uFtuT3wOVsvtqu7hyKRg2KiNZiOZpEYGJZ
XSGGu3Xn3IYrk64tLopri4ntqysU1q8M754eQQ3jEoBUjFXROfxfUIc/2+rn
PqsnV2dbWRKy0DicqlAeER3CJ7x393rx8y/yPdvzTfKRNR1PAI198U12PeHW
I2wgyS2YSVq2wyEG6m6PlFnCI4rLMGHZ5InbNKdRYQdVAndgUvoD9Uy2giyW
BRIibSfXfvLp8ngRImAZholAshQcqGoxj/dn+KgWCH3UQCg7peJzLqEY2Qs+
x8GXFuBo/fmiSItsblVDxW78tjFtZkIPNxpASoLNNF55Fmd+h5HiJ0wWgmbz
2dRGcfW93P4ejtA7lMxVy+hadW8iE172yH+RJOFJoJqXPQu1cSIpg6NJmJyz
QQeLylEPg6GLSja+egMQx8WkedFy8WOn2TYpln1xPWpXPQgjbh25w61noybW
SZxKKSPJqeeVKTym2+xsVXd6hQLqT6S4mqzfmoDw4ZBqlSbAy5Zif2g9g5oK
AUsVFKDhKaUcpIJhsjJfddLeEp7YN0ew49nUvmHZ8Wl7si2PBXUIOCdlNyt6
IgHq82FyISdjJhuNOxx6cwzEeZIuSRmufkL2jarKePzrybMUdqg1KnbdvnVG
M2+eCBUmgUG5AWHx6Goc2LzvhOkpCn9cJX92HjttTWExkSmDo7lR1mZ+izjz
TBcpV6QVEdjxOHKeBqSrMb8wzKsZQogaC9tps5SRJr0Xpxj7jeO9AGp2GBUD
UATx33ooQclCixcVl9uyINmSM6IJYcHtaNun9Ew7i8pLu4glwhSP2Y/nFWu7
zXTbkeDmrxEMaSTiqYjg2BmDWEWIs5xWd5CQTjVxcyV4yQDBTb46uaUzrMjI
HrNg8VTifC/8pFcVbE8ZNmm29PDfGyCAJhdRAxzzXgnymHaUIsiLDkPHj0V1
8vzwywUbKOiEL/SSL0YPSxLxkRPbPPI2++doQAT0Ol5u8Bj/hz5fNPwCOVJN
3OfqqL0Eoq1ev3FtU3xpdX46laUNTUCe0kKxhQM81/5ba+O5ythJ04ZgUIRb
SgYTaVR960F3w3oQtzHHGVtz32QkeYz8abiXxhTpmczP2VmS8BP3KQQR4OHU
YsvcyOfdMhIvPG9u5DYNFDtom3YMIXEjM+rrRWH1H49BUGVwzjTA+Vbx60Fd
+ssFdkoZ1yb5A+NEAKbM9AMuhp2HgD6zFsHOEJKLEayeeFZtxpgTr+WlxjC1
C3MAjLuhSWCZW6g+OvQaiRH6y3L7vId0KsSmszaXLnSJ5wWQuZBFnM7D4Cjr
GkLDPmwYBgCE9wj7ZRHbp57qlsFXEVmaxBZdH+pgqy1qYAcirP7gZPcsMP7A
xRdVgrWkomUNBhEcWnGX0PRq+/SsOEU+7Pvy9rykZwi8rxWDUG5CtLDto4cT
F2QfH5W8cNeKnOxZmWwOSfpXb++GHA153+JyJ0tSjW8pckWCA1Tm7sXqxgz2
/d7FiaApnf8SHSxlTiV7uSAMty+tK2v0QUnNkZao5iVTuQhKItg7WRxdva03
Ag23twrp8ppyyDKkYN9lJd6TwKIjUa3CwkEJRHbtg8LkMpmjI8Iey6qpWzOz
hf2OuEWyZLmUdtNRrTCkzLQ7dUAD2oPUXYyX9SBzelYjM1Kn2icCOsviOR/y
HlsgRS38SOREaVE1NzAMOz2lWEbYrL6L8A9Oaeql+ne9/IbdINzW02WnH6Lx
4APoJDiIcDYoe+uPBKcaAWNJrQrLXt0ET35+JUQx1CeskTCW3ZVGXnsdfNte
XR+dN4p2xIjwJMbIl6V5IrYcb2nbCCFs5+VUfw1XPvuGd8/S6EWfAit1odCU
f7Rc3vYqsGkz5DbynMTPnTlazigc2HhFkVx/RR6rW1K5KFl2qNrQDD8NG+vM
okk/uibbutVy7+m8E1ZV9fFAOsLksSOdgivpy/bYqd/FKQcTLUHNRLlDjPRM
s6SzGSpS6kF2AFyAVyhyvtK8yMV42PPCiY7bhEUvAnWfwbpjeahYoYzQlywL
Q86gUTGBVXMbvpyoTup869obMZGo78X+HyoylmYmGbH4K171WcFqF4DDfJaz
VnHEYEdYWftPqrkE3t4gmW1Tt1ZSefU0/PLHatH1Zgh962bzbBUFGa7lUIk8
wT1sJHDsn9vzPWsWIvXX5MtSAySSUZVwRD2WZ7jeDuz2aTOlWlYG5x+3u4CZ
x8cA8I63racLmQnfEOXk8cqdNK3Xz2CrLmtaekqEZ0G0u8sbylLYWOwM3cd+
gHhxbFFyoXZqg4ZKyrh4mLuHXoM56D/k4l0hRTYe1lJiqbNezOLAgTHqrO+u
6ZQTVdTF+pmfvXw8V7WoNzJ1R+8E2pk3xebsRWsDaXskwIeEpXhoM795Ogb9
Ik/Fx3AtXj1m02fGUbfccTZc/BH9QWSXmS1kNaXCW2hia/4D84KGZ1diwjeP
V1Ur7jAz/0TrrSBJlQwucrwlqAyiSnQ4RfUOhIMLIulrvM87tPR/b5wBU2+G
00LQXkpyoSbo+dw0dXwklP3e5I+xZ+xaste2hjLmlPuGmTl0F8A29n2HxfXv
eIuwJAAs5IkVRQnALH427ogUWQZLSDEFV44rJaFZor+JNilCKN3Xug0re2hz
SmKD6qkkFVyiQkm87zrMtgRIGBoXGuo3SZC5x2x+eTzBJVFRTtg5CHlNSLTA
xxCQhynz5FOMfwoq3nnKE/aeqNQjMd6GEQ5z6K8q/MIUGS3EZPOaDnCb2EPO
rBHVnnSGW9dwOo2uKAFHxyiCCevC6RzrOLR1zA8c9U5iMrSZgESMC3D6ob89
RGwcSVSM9/nzGYl6Z2veFliOx2Qi7FLyDt1KfL2GLqmO3ilo8LvfhkaK0Msz
SSzR6oKG2YCYlANGKeqFfx1VrR2t0n7jTLo3waj3Jex1O/sL6sVa782+vPP3
dldVzbolGtzvAqcOZJP+1miH7eGqTIGBKhoJ7kBIUg/ssf6NWhTNwgJ/LjV7
XnGrty00JV1WT29NY9GHWxaJEMUBcJMv2gHjDYclg6ttKOLWXwF+XD3e0+a6
3EoJl74e39n5NdZMKsRbzfiFWjIH7zdKKN9EmHmu9EHQ6Yl5f830Ipf+ZTir
0P/3ONoNHI/Ta+2uxd5hStz5b93Gs8segDshKC8N9/Go40OThIafIWoSRmq+
g6pikICbe8DUL6PRsn+0+o3CRvams6szlxjnszDrzOJrUTE7yznwcHtX2ez1
7hpSyw+E/+8hHK18zc5fdoRJenb19NRy9HpopKQOwWVs3X5TOOzbcHPzU4wO
1U9UClrBBdrn7P+vJXO3JwS7SWUyVgOg++sR2064ppJ6FnsQdsoId9gXVnP/
/BooQjwFddobO4hM1L2Ze+BhATZvQV2pGej88iSyjHOMRtGMm/26BFzK1XYp
PSyvNxdPjEucPXErsQolElKcXj0AHWFtumzI03nMY1foj9194Ecjr8bKtwMv
0jp+S7RrrloyBdK8FT7oBw6KzZP9o1PHtRcaHSGwGqtC+ar00Rwd8zvJsN7Y
XvvHDKBj+nsnch8Yp7lSETwL6//rDajgXF2xZQS/8thbwx2ockfef9lEqdV5
iuhyjYvYxWRyBicgt3Dnyvd+m67TRw0SH1weaJgmqJiZxXRt28sTv+7Wz+Bo
8gbAsPwmaB6B43VXTz6rXk4BjHFROJr56pm3FxXye57hZPlKc6s+R4cNIphL
90Z8WdLif6gwHLkNzZfcutLJNDDsdRoaqMTuW2QQvjXOqyQ+gpdqrh9lzolh
uRD0A9X7pcyqKcDOpE0TBltPS6AW1l9PCLzQz/seALrjyQqN0o1quHUeNmPh
Wa41NxYXkA4EUVa8ecRc1ne/71WMk+ofIum7oKAT2J8WgiSOV2lDoRjb+c6q
B076oQYjCH1Hyr3a0jCAQ4y+2UW3ALGytpC2Xo5pyoXBRtyOoyGPxUfLrtOr
PMKvsbMXf+Qx27SvoTNxB5fKc3DzQIr+1JuRrcBNzPQq514UPm0a4u8W1s1f
9n7D9bC8ycxt2VXjuF1fGIW0PF6rz/5KRBwIG8VOW8JhTnARm1RMHPD4cXeW
+pO2pJ3cLAMOndszK/0SeVE4W8ilEX3+sUoQ3F5joitC2O2AO18Ng7dyC2mC
P2rsSslvobjaewwIxD6QQ3HxNBQtb+QITnOYDzeeQX9wef8+buTmFlueSKtJ
ilb+EQMlpTeYUCyyDyHG5ThpUGf7kLA/ivdmeUGaHD4vw4XMa5PhITm0SmGP
ZLv4wM2GH1MxjSwUwednfiV0qvjkKWenNlnD8zBYvwqhNGC7B7jC2JggAXsz
jE+aJnW/sWlvyjq65SOrLZfs7D/NElDbEJsalc4vNjdKPBs/wNHqNgWIJepQ
STllCgHoF4gWMWt6sQGOH1SEnhSEYHoO0oumjahlQ5tPCsbLb+f614m4xSli
eUqu0fLfZ3bpvmYg9RBZC43xEW6lJMrZNFRpo2ZwYzl892+f+SKEUttLjADa
Z6c+4DnnDuXEMt4LW8sAuWt7cokOomBGPsyyff0kOWcRW00SEQufEtrbhpGr
FQFj2zWZFJiWgnsgVm1pzDB6t2nSLmHxJqrAo9iDBHwAfzron3hVaHJm7pB+
It/FYHZBzTtx+5fmHMV0fjS0SPRTX2SUr95saKM0WrW9Kr9BYH80sr/L4i34
lEaU6bt1yo6asjy5e4GQxP1zseFNc6AmntOeFM8+uADC12S1LHtzd3/NyEZ0
QyhQHt/po4fDXbijbT8dI8+GjhPlxG8pbimy4CZnD1LSU1XQfO/ndRPHI6jJ
lqJb4VeWBQoOzXXrSoTictGqHs/ZE53gFenPu1cRthgjU8a5Af40Cdo2NnfP
uwW0Co2+HR0mWUba80ZI60e4sW3SNGCHXoEMpZWmHtLw4G9t9dhbgd6KOZYZ
K3gBadvFGUU+lH7xVFIE09U5Ep9OfBSE8wrKL88zhg3tYpINXmz0yM8iiYLR
dZydjqsQd7Xp+s9B+0l4RijHlI2ud6idXlaaPXUzNHs9RqsnHS65hY2PIIwu
piKqrJy+uwdggooFOAfjfU1DeM6hmxNN3tis7iud+HbzcdwFQnu3YVZ9XNgt
E5GxeSP9FTmKp/l446CyzB8TiQYnqQVDqKZM/n0tLjIu1/tFHojpQavWNpJQ
MQhEr1X3Ifq/qq8mLdKDq+4HRAnr5g3fiCYUJqIRFBqluhLjhLlty41uGyYS
/yTEnQs9Y+RRqCaOuEQdFlc40qTxtl2j2gl3ONKot5ZX7ZEr+IkclN3Cvljr
nW/CEdv6GT5I9j3zL7ITLacWawwKfwiiKPLBWlB6yFglr5jNgGMYBh1BSe5O
74bLZXZHUeEqLKmqcBeffWNDxs0BmWK2kV7X/1VYamlNlo1/WwwlvmfKdqcx
5ZmBNY0xzde/BT20gyje3drJEsfofyvVKPoe8n7y0fAWjDbVoZAZp/mkw3rg
mhxWASyBJlf7ZQwGDjEJDR/AcfL420o/N3pzJK++329y0sZ+uIGZk7r9mZzD
hMJ8b2ChettodtvszR32sHDM3U9qcZFBmT1sfxCdGSgex+DS8IHZBt9JAig/
2gV1RfOnEqrVONEJmtyEgSCBMd+/69/1FAJuIv+UUyTjUh9JVuyYsD1mCj9E
Qc+mB0gdMvvccIiBep/UOE6f8+H6PMLx1fKBcyJtAetamXypaXpXK6wXPsc0
A1hE6ONDcc3wgO+eAptTIxpvqJhraX1WcBSlbOlhpUAD6COVioRSl4AG4cLZ
ZuyKzq2+Oq2lME6cYu4XTAbcuCJlCwFtlB9DqLadMLx8CzYi1dR0Cgqw9NAR
Zn0W0/tWQIBblrLKNseRRnjxeZIdNF1NoQIdqW8gh1C6P+I3UsZ1vhUYdK8Q
Kcmwr4WzfavlseSKKVh47iglzqaoYO8VophXISHyRVh8tmMn74S0dEsRxiIA
5KzwlzmAmA0+ICzhT+SM41lKgxDO3FiHgEaF3TdtRcNCVaPOHpvj8AadPpER
i8OWarubWOZRappW7tHuBWZvzNkDW0zZjuL4mdtkP/KfTnQhNE6oGPgFgsmk
4hI5OEQFZlLfAx7e1xFZp5oesFEpdctS+IRLLnj8GDxQRXB9wBh92EZbfe23
RciTfze+tRk44PJua5n/JAVxEpKuWMlNbVzoZloxg8Sb3lqsTDfOXmapvoxL
5rLG7Vtxq1v+RMgsiIaU1Jazi2r16rrj/45gOstXl0VamGCgoasUSwMX/Whx
uysl+HZwZ2X4XCZqztne94rBnrf0FuSbVEQqNOjzQ400+z+Y9rHMOOeJfsLL
mGjz6gYkrbRN/vSa72uWAWmb+ysEJLrh78RWxzbof9GPuXQGq53EfDVYQGpj
A80QPUIJ2qp311uYcosR7g5Rk3g6wR2qK4j9dd/lIto3Kwn/pZR9kr1aJ+kG
mdYjRvemWSUSMJF4utBIWq8u54i7NzfYp7E7RdSr+VO1tXkjzSqcdEU/ctpb
c+hgbD8RK0vR6ORNjFAxgMf9Mw3Q8M2yzZs+CpnM1iRV7n2897zWSorad5QA
06Pdw2UD0XiC+LvwILbgaQ0FkppOJYZJ6/0OYB6nyGhoXoeLVdDgd0+EDkGB
BbU5zCLxo/vx+5ePxo4JhpppuROwc1rDFHai1LHwt5dME4DCRErGIvdFEpVD
AoO/+RsPAJnd+87S6wL7U9LxWEQWG2wHPJ6iFHRnodO67t/7CWKJtyEyErP+
8FKz6CIkj8Qh0xXMIx+tTL62E3f/s1lJlGDR4s1CXbW7xS4w8yEZuQAHMyaf
ZsEG5rzldDi9t1J0x2I6sZs3mcMy/NdqO5Be/yOBM9lvJ24Z9xsbqNWyKVNz
IGT3+gzGnjgAYmM0/U0eEdiE9QK4THZLIwYcJXKwHsCip53BRcVbZEqTPdIj
wb7QqoZiEnlOrB4OlKefFJdabc2nuhKq/oDLPxG/uTwQa+1Ntg9fqX6au4MX
seX7d3+SihV6iYZbhAH/hQp5XpxOChZ4aCUXArS0VnapTpB8jbMW1YXz3ne3
3Ftn53ZlgskeZ2JtcW3qoO7MFn0K0RSH1BiV16o1L1yBkPN+iONNI57LDdBv
Um8jWYxRIswijhWsSrgzEMgc3UnQsIzySxVWKePTE5xcSJfT/qsAY6OXCd5C
jVL/4Y43qE6qMuLNfslKP7Nwg+dJ5Zg5DVK1+fAh+RbzHN61S+dXPVH30W5y
HV4xpXkKwBsKk11R3rryRm2VQbtr3Km17Dh7gKCSJiiwhMdgdKW5oMCqWv/0
hS3LxfxvIgHx/1LC7KHKG/cOexaZUYdSQGvmT37vci2X30V2LKQmmNH4W00h
7yivbwq4Z7J58dRWISvm9m9lWiR760+eMsnSj0JybuPl3pM+OgXexDzDb4pm
34vi6EL3rF0Zez1SC4k8BFZ2bgxXARrGVRC2OdlISDmMv55lSwu1bGiwuItP
wDuwnrdKrLVJELQRxpJJNWVf72oCNSud7xNjeJiG7bCZvKsc4qODGDw6v0zE
SQaUlJIOL3QmkTAleQeVYdWsfGKYhkEwn9ZjbombYHA4Cm/gYZt9poyPmBVj
VRYzqVi0YzG7fjHtnV43ABujHWUK7+1SHtxHXQG4oac1hCdwmuxs5nHznEar
oVWIPLlcRMYavG4aY5ZkIHEBfHqxD3+8vCVTwODhNOAZRZJOAyuOswiFJvHY
6IadkkSnfUeuTCdhiHDhjXgmoX4BG7ny4L9VykBoEfh/pKAOPnBIcrFmZtaS
Jd7ZiXtDvqLxYUvFHTDKSLGCE/25rX14Limcf1NiHJsPqDbdIpHd++SKgy45
bRlJmCQWCAlx0Q+L7r5tGmDBgvuLSjJFacu74njAOO8LO0C+Df1vmN8HQ8RK
RsPphqtMfGw3I5eOyNveM41kT/1UBbswl/jwRVAAFYk0XJ0lrSf3OpI6uk0t
Xp5Qw+KlrgOKfXZmlaMtI548hDG8eU/eZ/MITmF+pUVk3Ptjj4/Rq0HjvOMt
1E5wmIraQXCbEOPf2jKZgEIa4BySOQgOsoVukOen85LPU+tvpFNEUkGId66V
MwGnoMTynqBKKAW2A2PvWv+cD/EZ5XWjQgSZi5nWD4tXwpkB69ShxfQM5DGB
OMUtWAQ2L1QAnO1HTjYFQBOxNDtcJV/vajVZN6fZuXqNl76Ay9xYUaBcsR+Q
vhuFDU8fV9rsrliOvXH7zwWu6iDE2P0Scda/8e6pdm7V6l8EVwxL5GY0r8o8
noTXbUD4qJNJVJnFhnuSGkIrLcSaoZcJskIeH4esNSCkv6EOYiZPftLXrtik
bYYB1e316l7EfmmMOflvnkmmVMDNo25yFkZ0oRoyJH3F0a7+p8T42DYncI1S
ejrIBUfubXgUTv3sjFGjwPvVI3llIWO05GLGf6rqSnW4heNxrGybppNvHAsr
2ctTi4Hn6oxabqL/dmqfxCM+e4Wpt+2EOVP3QXo5f/beezUjCKq/mxPbZbVT
ldAijrfBWIa4SGDogETrDc/EDRKNLI/g33LYMRaXfcjJ/fzgQq0aiEUr/Yif
C7xHj+WcLaV1eU9htoW0KXTeEXut/kZyVt8PWJPtYEhL/Snv2y+F4K9IWzIg
vyZ1Ox1Puiz87Cd+alX4kGm0ZTKWN1K4+hGN6rPaSzeQvu8XojYn+VreMbF/
+vxhRMHHo8b+prHYlF0+zqmbtZhdmW64tuJpYrqZlg4QWgH+2E1ukDSFZnJ/
89L8XnUmRHhvkU8Ed2yyl50zq0jYVDp6AabAV32M+YcM9ym1RKARR4NJupQa
6Owljfhy5Unbdm8e8lEOrplrfrfRcRu4IaaNQYrVHF+QiZUp6CgW9WhYAWvB
vl4gHvRWd0uaizawACZrNFrFU+/fE8CSOW4Yy1ZE1XXNf6rJnU577EsxRqRV
DPG8arLJy8PbkYCf9zy128oAjXMZScmn8Q7dZem0JAtednEhhgDhuhjDvRvc
gO0QwadGdz2+LkQex8yCkGBoNLboyJXiYkndkvrb9wM+ukDqv40gbW65psXW
c3C4ly90ZXmSmwRTIfT9S8D7oTyRWGmqXpA44t+OE1yZo/MknI8ERvbHKafs
BFmKHXVyfx31bEsQWApfRtk+wAUrKuvB4yqyBpUOGZ/Q772zpjc9rz1ediLP
LQPi4y9veUw8AHAXG5HUK8StFTMhmXuznTVLFLtdvZSyXCm4IVgXRbb6/1C3
85BpyReAcQtY+J50HkEK5dA23TWIgi7yQGKS8jWnJjClFwWHqrNM2c8U3CrV
pxH/3zOxNTCj19yb/RamQ9X6fnmlsD76qR5bJnWEQM7ilOi5JmqBQdArkI3p
XULkPWdmeUUjzJvPi5Ntn2LZS60X+gUSkNjALoFgGj3pwVW0vX/vxdr5slLD
t/jY45cRcIee1dYfoSVtVbm4xKdnCpV/1IP21SkAXLSUYdp/AP71Xguoyyx4
eSVTXdhcSIog6xQzpN2lgw9C22opbb5EmpZT0cwkdvf6Ui+0wAkaHC5QW+73
5IfOzAG8ig1dmbbTn1YNLamHL5yY9fQ+T0c/SSCY9T6WoWBZKRdcLwRrIXu/
20iQlvM1DbGEXEYo56dPzaZ3z3rGt6ETiJjWZ6qquCaOm4ADAt54yF/ekJQC
ENlzKEE01z9N5wgiWvd7e2zCOku5iqrhuTeauy97ON0n395GSOlVzSbPJGdY
sOiuMk46mO1fzkTDacBhh9Z6bMoyQ5wAbD4YVDacONSyeu1RJG5l4hzZH89Y
oi2lLy3noQ1Owas30fLut0MjhIE0t9+NBfGTjpA1AGRceM4qJN5o19z8iXcY
pWf6b2Z5R5ByFom4CO97N4aSZQ3iRRX+Y/9jYApeKaIn3v4v7jO2KC6qGX/H
uns7eE6qSOQTcy1zOXWf2lgW5R63XU8mXdD+Ne+nBpvTqHemMiuDooyle80K
eKFdRN2m33+O8KSJL3uc6MUMgx1ioHB2aaI3blJmAz/tku2LOhlmmwdEyhaz
iJDdmZzA8mPAN90ccf4xGQLtb7gvPMmzeRD6QpJLOV3HtK7+ClMbbPo6CtKI
DCr0c8M8vaShjMIuTVew05xbVk1y83a8DljJJ1VNXX169UJwS6twXq53aIEY
q/uRN2Uau3XmK8JaxX5e7T2PDgzahsaelYTEnicCnVlWJlA8fpsKr9vbBWb2
NFS1bJYM0Etz54gV63f5iXOtB35FvzauiyE8DiPKQDuG4m51e4aVtswECXc5
9F5l9YS/jfVmLmH7WP8N/IZgnAaRlyKHyvKB0S1Bs8sfVcfNhVRJrX+1A7yM
jWPX1l46I72DLENQtO4+4IRp89Z1YxI/Qw3EhitHwaH/uTPGM9mpbVapYqpO
K4bBdZOGNvZpuddNyMrdelTl7a5ko9j4Ve2bnMuw3ROXDgik7VQiHYc7CNlI
HTSoOxYQQqe3R/6kNSltXx0z4U6UQMxW79dylNqJAsWvFNt+/WqRwAy/oN9u
JXdmZ7uav+jY2HfkiGbXA3Bkg8/uftneZhguig5SmsgXIL4slgQZgyYcSGz9
kYg2OQYWCL8CYjQ47q0K18OG4CtMkMBCc8ZizMNT3VVbYwIe04AtzdM81nQj
lAjA/hrpSoVzXFMUijETdM+HGtOBjfTHxLyHHbTCLtsCiS5E6wwFe6ZRpGq6
7YkZbeQ2V/Hqd/XUBJARBPZ+O6dGhw0kO/cgpbesniuBl/T40VM3OtJC4vHh
5gHRQDFBBbJCH93Pe54qJT9F85kwOasQpCAadAhlOeynLBSqBZLZxDKX7PNG
bCB2Tjeehiz0COga5B5flxCjO2rQKxhJvt74gL3JOvV8k+qxFchxn6yJ7/uV
IHXS+CdYB0N1nodWHJRpQyQhVCMBLL8QLhVKl1CmD8fuY6EG2CKVSCV0/Ml5
OPpv/iCGLlu1Vwv+D1JC3mYz89dCfVJuMX13H8XbXmoiRoQf8KrNsiT6Ra0a
1IFeL+AfMQhcNoM0/PxAGVygrQ8NpDjV1QgwrI05A3TCX6H/bjG3Kjo/qfuM
rqgmU/c62hHGmMeCmqReSUXScRw7/TR1zOisR4X1Zn7LAmmPoAH2SMC+J+Si
Wz1mE4QfYJ/kXjdYBp3QtrTvtqPfQi1jDY5s7WztjlwLOWgO8TsTE3pdUFa8
KRHaAN7ZYVsWR6qHKt1swGg8M5XAyKcy5L66MwHtuY4rxm+axpPhzDp8ceMi
eB9lGmu9IG4DAGcnIqlrblaV8f9o01ysQWnn9Pe0O/7iU9YxyS17xF7ek5/E
/tCil+LA+4o7sIl3lhVwkuwEkiDZA/LoiUGwsZbWYBRGjjaUz7JuCOBiPtb0
TdwYH73uPS+4p2RNhI4NpUQZwz4XYyFckWYxIiNLQxAnxDsUVIcYL51C6BPC
0PB42o49/ETu0RcnqZjBf3GoVXmhhRehFO1+2SWGolmdCcn1B4d3u1fhxwvs
aOIcclkdOpzoYaR8CL6u6SqoOP9kBLDrLdh8Cm+TIH5bzQ/TIII69f8IN9g+
0QkKsR9A/yT5ebRjKp6XzclbsfqGCcY9sprMg0ZOjwC9BYQOjzOH/jx5kqMM
/Pa8Y/1sNfhRpPi1YN1t3rwe8YoSQ0BKJxQr7BRjI659JGyhDzCjVXC+navB
WmikOPlDVImtQw1pl9wYXQbPmGnkrHAAZNsJWRifURIwIv2Jw2a68gGBQjGy
OSZzti+BPTg1iPkOtcnDPvPmafbNum6j6uLjPNyhxkos2F2p1oJ7MQc+/Vvt
UeQ0l4lxg6y2L8Bq9zwO2hqQcXj/yFLxNkWg0QS4IwZSTWiI4gfwOKxujh5k
GvuNACrzabu4CcF7oqwfWslnFnmAKh+XBa4cW0MnQQSpab6dN30/iylO9Ahq
54jYzohXZBP24pWvqGVGXGpIOfYkO22LrlgavHnXD8mEDZw6X6lgPf+VeKLW
GPy2vxo4g/nODYDDAXPkEMEPYUzH7uRLBG9Lqx5M4yzopB46l2gxAPskSvg/
R5HRtGk78Mn4KDONpNPyUrw+KCN6/weCONYdsbNpVrvBYadriIosEt2Fkirk
QSoMPTA9zfQWV4M4W/6zPrFo2aAJ3hF7WGqXSuSFGrH8mLdXcZGD4xq5fQ9z
redBmofcyGTKOFVpVbcp0jnmWHlGc6xqCbNyhIWW4ar1CV1PKVjsLJe46ddR
ZLEVEOYS1z2PzFDSw2F8OPgkOEaO4ncwqnnqovxMJP+vOSeZ1jvrEagsNdNb
Z2xIPfuUyIAkUKBTpcAtQ92AvuucDpx0PZlQ+o6KB59SY5rJs7v8tHrUKL5U
QhjvDyI/ABWvT2FQAe8Svx+0B5+8YLzd4i+FaMwsKvyjPN97JRbX68EHQwpZ
eovR2uneL8uu6wWNlUJxSMxgQEOAFo3w3vXrcMa5/SGTJp78Ksasqzrdd7Sk
yOFHdyn7KbbsKdHLx5mYfVhHzbRLqMistUOUL4J7JVJQMbAatp/1H9kTkEDF
z6hbpqWR0uTFKov+T6kmAvRVgdmNs/3qLSCuTUWsexEDuSTQ550S+u8YTQyM
2maQUVo7rVUKgc76stz7Kc6CEQPbfBSAy+FG8AxVPFC0sb31LQm2cgZs+0Qm
dAqriEAAYbIaUqZ65m5H1wBNrDVXEVETUTUdn5XQV+C47jAmFh48ZlSl+TKM
elRuFFJvgnlcIV+z2zPilppAHPbA/ikmK6NX+XlyAxa6U4QN8TP20s0dR3Md
KNMVjgkOXdpeoEIw7zyz0b8uZSli7x4MGEI37b6lLHvlMDgOg7YOgUsHSAhU
s6g32Bdbcmv5DZvGSPhu+kj/NX/jiajWqu9HVxl7Tbks6f1u5UmhNxoJcTwR
dsZtBnnj67OTZ7kmWiQGq0guH2yPc56WlDP52db2l73DVna/ESwodPjAhtA6
XrIxsOJZVPG49RE5aZqV6l5RP2LyHsx2sv9LaA3sBVkhuggEaTbQp8noKDVK
pBjn5fd5pM8pKEwdr2NA9S9W705oG7M8p8Zs6pBPVSuPRqU3/iCllxJIkI4w
n1fSzw1rE+g/OPF0G/9uB64woVOKXVd++hwbhbIqzfkGbqjKEM4pVdcQGhvS
fzd+D52UctOQoOlDtX+yZ2leGNYhZNkKoBn2PyFFcRjwpYRDG3jRgdjcl5W4
3PwRDYZHZRuw2gGi8PvrzojOAv/GE+as2nEpaXvGh2Wndmbeek1pvA8Eadk9
6KWEi4sjnZo20ey/Wa8Uh7+fek6abWaDy16eQ/JpNSQPtZ9xgsbAtVvc7y87
f50xN075kBZ8HN0MN8FOkxuUaruU9wJCZTBXDNv6kyHchLM9lmurKIuhQ74y
mIU/rF84s5EhdD8vtZC7RcWR9T9A4J7NZkbkggEkkh1oi27KbWULxz1ocgNS
aaRK7JH+183Y9Qj1M0dogXydCfxmNIOuBDG1gNSww59v5/Ez386DO0g2RRSf
gOfTdFn2HC1ZsJlZHHQ6gsGpZpkFxW7qP2ZE6V7eKB6/YUrGkrMX8co6Ek7j
R/u54oe27tBUWaAvoCB0I9JzutWY7ACJVKD22T51xCjY297xhoWcqzdIRlMV
vq7uEjB/dHyBGuvZVp6QyX+8OYbRv5icRh1IZRso6LCnGRdqciQFTsDdvr7p
bhMh/+RLgDrUyLzblPPTPkjVqP81uaEIA4CltiJsvBCYWFviSiMcIHJXCcDK
vGRRuPrUFFaP0Hn7A0+sl4JsCBvs3663cfTh3HZ3bDDiVCH1NEo0fQznUFG4
MICBUMsym2Yv7SLgbHKZeiD/AvxPjvJ+KohN0fLvPeQjrlp7HNb5Zo6uYtNw
OOhOo4IU6D8+6YhPp1/grzkaxLEwYLEIysbpKFaExqZQXNec/Gg9HMVuKHVI
/Id8oUN5MN+BhYyGhy8OS4qmNtbaOC9zzSDLpbi86Lx2MD249hpT8WvfGxsQ
OeoPzlhPE9e8N9v2Pi426jhVUvd6tRanbL15LpsH96GNMe70KiuKKWdYkr8A
1OIqm6Q1dXld8tfXAGv4iK2mYJU2F0CMaFo6EvO38+99TOtDhp80M7PNlwBH
RYRC+fwfTvM02dz/+MH78MGb9rlM1OK5M8JOLkcqPrdZ58ujo4DafgOZbp2n
qWSwyvqsi+G+RU+ywJheJEUSp1sZT+Ck/CbOqWAH9JciuwQtFcWNPcYoYf2U
8Ufw3OhBhVo6fJ6S422HYl8NVljLbF+3t47XwLDwf5vykAYWuy3X10xUVnDB
tMHgMuhaAUQla90nFxN1lQlUXfAlJjiWaPQZL3vQszmQ+A8wKR2AcB39Xu0w
eWVuYCwdLzfMVVPsJYHzFOh3rmTP/O9UFUfh21DdV0CwrkPDBKM9JQaYwvBA
NCx/s3xZRoCSEirn/nfM9bdr8EVm5uvAJNbRVsc9UVKifnaoXnWYtPUFcto5
VEvMhV+C855vXYuk7Q9Q3FuEDz0NfnmvISn1ywVGTABLBOQKpwvqh5ogtXup
Zx7yTeLCo7x0Py/qSVwTbBRdbA0qCPQ9iXj80aIHrWJhIzwKrNiv8RwELhMu
1RqOUKY/yd1US0oWPQjsHaGNKxJRgmkQjOGYT7/HnEYviPJ38BwZPzuUE2v2
IVKitRAB/omdy0Fq/s26gIzTh1upr1Xilw5oXuq5I4aer7BocoGZlgg1MOdR
5pl+Uo36wWgBe4RYuToG4vJ0ROSAD6hs9cIAE9cipfclmGbsR2eLwlbo7wmV
U4rttmO7jkG+73tBKBA8C0g3Lk5a0+DwYPdK7sKtjokS9Bz+Pi8KzIQRlZC/
qLhEiHeogwlZtV1vMDvelV6xDL4bxMe4/Q8S757I/wNiZXgTvtMHZVx/PG4g
XIWgfiv0hiZTA4EkIkxiUCuWJBpyRcrA7j8e5bRa+a3TT796HZaxyvQmTFaB
oHfV171hQmfuG1xFSW0II9W+cgKYaOBrlswspVRMxXhJm26ubiIV0auZasq4
z1Hcta5U4Qi9FjvrOZkT+jqZx7AyIh0rSjZgSIL8qUasHn1EhEmDZ8NJFyJP
u5wQwEeVQptTncLyLNGfK++0c4i0qm+UxKpR8oN9yAyhsOgmQXYlNkg5E5YT
y14MHm8Ac0YhOuJtP9Aux12/Cek15QrJbQmOWM6/Hj1WvLG5VCJSlT36kcBo
TGtfa2erEKFBD03dMIVnEK8jH+8gjFJ8UkBPeq+3kL15BH+4Ir56mmgDUXRC
kan90Zf8HZ1jUklcT37UKd7B6ViucA9+23diQ5lbTIlJgxOf8fI4zYbhNUGf
1/mmarFGnPYHblHpmwRmMH2ZGwTcLTZr5Ln/pHtwffaljD5WCptKCPcqOUse
QbL0913WT8DGWDWyzxFOL3HzQ/TLvCnQI+h++Bru6kUBxOqyKQ9SQvg3t0KQ
ebFFkX/I+lR/Sq5gnDW0Y8pD1KRosG+ACSvI0GT+/FwAYGS9R6f45ehddk8p
pgQc7e2zmPOIWXqEGeZ2wJRnywmHQLf7/Jwc+q1GoKOpDgojrFJk0CLw17iy
X4nvyoLY4J0DFIWaaBCx2ISR9LdaxUlfGNW3HyK7PL11jpBasmoNc9LrVMzk
qGJQyy2ilWXMhL9gg7R9c/+VFaJvb0Tca6BIc6m3/TkGe52FnAqbRiD+kBmf
+/pSSKtQJyyZwzOdScPLTB/mjcyhKh10Sbv7sBfDts9k28eum168EqZbsZNI
M+P41THD/jlIZ5aMuN7mocPTmX3uohiU+kUuQiK2nAOtLkNzggmVuwGl6UGz
92zQVxUvNLUw9NHaadHZ6VqQ6cUlfpvB5gyw8FXiH1QrxdRNBZckZdzOD0HH
l9m1+CN+/9JHbGKfm8nwELXBZ58LRPkN2sHqT1UIi9/yF35+C9zXGpFOyHcx
DWhEY4G+hvS+qTXJXXKfCakjolQZ/YDz8L1hyu9bfRk8AObmD09HpkRUjDj5
ZaxmI4jOk9NGbUinIhgX/Z0mPxUzWvOpeERc5Fx/ZIURixZX99ISyfHhzBY8
TGD2DG+l1+kdDIdwW8wi3DKtI7mEaSacaI5H62AA41VC8t1SwBnJJE9KJzRT
m2ETS5w1W3kcmsgaeJb0kMhodIpVscdIhNWkqy2mYa5GkZZeTDALgAibgIiQ
BZUNdAuDTrQfKReZKyrRZ/EDHf0S84r0fFhNIOVFpWYuJlffc83Etwz/NtLf
bsDvWhEHhLhY/eZ6EPYwfsYXWabsYJWflsiIa4xm+42znrG3sLDLlcgisizv
I7h0B8I4F/MnnWhtF6gjl0RKGGx0AM/fS6CZEZGA67EXe/T4i47/jnAaHwUF
KpK7mwmjMhV0hQxR1evkshbQ+aZM1iBIbQ/9MLelX34Ii+jrnJMtY8Ys9nOj
ofrvQWaTp1R5jLcuHwH5GViyanP22Rjn9beZ+em9ZIO6uSvXoCSgU+i3Szvs
dGBxRZzNc/QhGpBQzfaQkAW/j1DjDZb49Z7IjCYhzOBTdTVewytV6DXb+7Rs
b/roRiL9SZUZT4fx8hhyXxmmL6qk0h2o6BM0/ikobc68FKOtMZrkXeeONz0l
GztkAx5nH6gbT9Y50Ldw5JsSDAzlcV22o2eRdtv4P2K2HmDI4301VMg9+wOy
0tt6C/Falh2tt4f8yVUtsyrzu21V6nmya4RpFnwnSL4LyCXS/IUF0Xgpo8GG
i/CPL2uJ/Gm3X4aYWcFk/DfSoXrvyyTYwdVvHhxxeaVmEN3s2OlnRY2H0pMu
G9OHL/AvJ2DVSIsnsmOYy/HI3emLHghhxMhHQQZzfFwa8KUfdINOoaTAKJd5
9qeLgUffFWEXd7aHkjZUUgE5RhrszhKUzo1+ufvNxA/cR9ZAy38D7ncQMB4A
/kWay8jfItWdsO1rSuZ+Yd7q58SW0c9V+cnGc4KdEZvL0Hf9Xj0QPZ9SZdbB
1cLfcP2/cwXfXUOwwMwpOFllBWjiuJ7IfWZzkdKlhtPrTHyOB2yGp5iS6yma
PGCO+k+WcmCu63/TGxw/QEaA6xdUc38/IcDc8zon2tphHuCdjAoro7GRNbaJ
+eoovuVcmZOsURzUaezkpidGveWXYeOt1rkwFFmLrzCKl3wrByAFbr9HQvAi
ion2Hd1649BdELclhZvF4lh/7OezdJlb+59v6bR6PSziP2jcCYW8rf51dDFN
oAPU5zDTLLB/z5ZeWHjDUDUQHowrVYyx8tEQ/SERFa7Nb+pUBEsJjAiKdguB
GLWqZAbYECNoBBJWkIVqrDEVAAJ5L4/PD1h3FOgCKx97O9ddSWOfcES6ItVI
UQE+Tby2CidrGfrUP21aOZYAIb05djjcyoQpp3BBi8Yx9jrP9R4StsmX4DjR
YB/2mFhIzKd12fz5XWyM4g6ZDqDe0dvj4WLSCclgpdyGsBC89+zwdQDMFk22
6E79+iqvWVZ5bgMuvz4nfCIDlIvqB21vCPbbaUbQyOgNXNCLN+Ddym1+DeDQ
f4+uYLKsdVpBaH8ZAX+jUYm85x3oKCtQqMIw422Fd+S2yorBXlhzuGlC3P5H
u2Z5hcBSn5bq0cuBjzc1kH8tL1zlJBvn3+Wak32zWwAjPBtHmGcDyY9ZTTs1
3Cjy1GkbDkLpaGR5ufq9+UIf0qc5A/J3BmaFDZral2Ve/OPNG06E0MjoCI+t
8PG90U7hyPVmGzxsSAhHUKgOgNExksWLIpGImW++gMrMN4+X49BvTLT3/e/g
TgJ/yimlVaSjEKa3vgilLx6t1JLD+kmz7dZLLIKKCEEdo4MRui/AeY6b7nFP
XTfaWZc2tn3nIBXqvCUdWMHRrLNvVuw8yo02/CLR1BoHS2rJBNTfqAB+WpvP
zaLGfGYIsyJbr9PmzOKOE4v3nEE1HTi8iOOLhAlzIg5TZ3a6P4EJLItwZxDv
QNEo14wcSSRV5JNL/64T4RAi4OFjhCu0K0MaM0R08V+eyo5OEE5eoBYqHPpb
kHNzShw42K/WlWt7DPQ8WgEIdblwQuQSlFX1qg5DresewQ6DlFXH8bCq/Iph
6RBqiJfqHWCZDOgIitVEDtPHUaMCbeavgiJz8squ0Wj6h6kENJDREEQ7OiJ/
mKoQ2PGoWcqs4o7qABXkbch1/pw8xtq6bz5ft9hQxl8cQgF/0PXE4XuV6u7K
tSkCdQrNVvBWj11LJIl3TW6y+lwXgebdgth3EVJ3Qrai8SikSMKqg/q6QCEr
RggjWlHeTGr7k2Nwn9Sg2OeuNVoAVt5CXXp1fQQbF50xXW688HU2ZyqYMfNZ
0YDLI3t9xL5moyEM+FM1EPVKfhbitjL4zHt/L2VcyhpwIdWLiy8UFPBcD4U+
M9MR39AEl/jvgT2BEsvHVARvsxg0wmynb5iTiOxb4bhUjZffyczoP+uc735+
j3oXrZAfajg6d2ZOBPir3a5OnlEUybp6SBq/fN5Ba3tAPkaYEJmZC/5rQE0j
J/oIetna00H2cRyyAgAMv0PrFV7DVmXKqXHoCiZNZyjXuW6DXKKgZbR7MiBj
gkct2o5gJ2mn3BkX2Fy6pPEqCoeMcihYmJa/7bUnZ/6T2T+ofl0rZTBbF3j/
Szk45nWU64FEg8Z3rOX1ARRq8eNPPL5QCw1/iJnh/LgSA+AG/suOTOmoUbDe
UechowEJpx79m1PQJM5Tvm0tOxVN6zgAxSXcz+ZNCCB0rqW0egHatNY53x+1
8ibhcAVi3Jsj8K2C5xmepKcuXjBVeu0j8oQTpiqVeiFfHoaxPdDybWFMA81H
mgzT0bEETgQ4WRvB2PznIylu/qG+kRwr+t33WXj1SzaZgVXQvYjoKEpy8aU4
SHBQh1G3wcM+dP+6m0fIj3oyNANaWQD4Nvm5O7A5cmDWGLLMGGrSl7TCDe5T
ain5tMv7vFiRf+rH4i/OycnV47sUHj3pd+fEUwG/4NNANn3u6wRaLK5N2OLs
SnPGaCk7lnMk9LqT6p39fAbCpqeSWpWYKmly8ZJI6TVtlWjaI8cNcRvjqKgs
w3qRQZsWIfWcW8Oyl5tvVsu1ddHXJAuBwkEM+w3HzJRFL6k+0qYlVW4c+mDD
N6+sST1mNGmJh5vLSeb6uQr8fc32lmgXTYY/yPsGhoUOJqAv+2T2JtkrTK3D
yrytttbCR4XiJDr6FsDXT3Xjft1iqEX6tZa80p/s5pOVK8YyQSSpu9id2JWw
rkkgtn4lV8kowvZ20PsrgQ16xaKdt4oGXmNXyJSKbjHMshEsPYw8s3D03YOU
QROPZIksxtVNQ7D5D1A0FIzheexUOkoa6dDTqERnOKrXNAgaXmeyn27o24aK
OGxnUU1o4fSk9BzZVhCOwBLaJ9A6xZUk7U5Qfy8N7tfd0mocFqRddhcS9Y1l
d+rsYaY0K7NcZ66mqAu9OdUroEN+Z3nXyVX2Eed1RfHvmrGqrTiESm7uAtHn
QH5gRtorS4G+4i+z6KmbiedOgjs50cHNmdrmi0y343E1NJeGniSOfECVSjiJ
fRWPdTA30xfwk5QKM4fg5QUI7zz/xhq9nzAsQdBJ8m+7HfbkAlECeDZCzhMJ
evlx8gEZrF5uH1itgT3bo7GcPs12celCfOTYZO3vvdijkWwFulFBpkkkIvhr
i19v8Omd1M34Aa1Vj+scFJznHTOECglGU4CqkorByH4JVsDsCNKR5iHpH+FQ
CFranZ4iK4d9qm/4WygGPfMAzAOknKVwN8d+r6NmARw/xsQ8GeYeM+uKTQyv
i+kWEufhk35QG1iyRtijcp3/uP4+s0ZzVH3U/Nk3PEBZYiPD92h7km9CQmpD
yo5kFCiguPRBCYNI3QmvzSHIzyp7WcnBbGbXP29mofWuPSv1XLCZYHC/2+MV
Vz/PVTCbCitOBQhlJgQ8iNt7by3E3ozF3msXVS9p1I8gkiaGPWf1l01KH3jS
nO7v6okj9UTcASlaRBleOMBiUijmH1JnzWlNSCzE61bT80GMawknHnaVjQFj
Ta3bY6s9D8YwoubWmfnxQDIO8G7bi8bwRjLxaqhayLe6YxfVZGZg17Eg2Zqs
OdLVKPfYRvEPXPgJ9lBzMjPhiSvRXQPlx8RR3b/7qg3ZPvN5mzf/hkcwnNLp
VY1vVkwEOGHFUZjwUzXSPmyVhv7EOPDFDBq54pjDZLpWivuooQKO1dWg9VtA
ZLlY8F6KpjyDQxMlZ2nJx0e6948RgKOM2yAB0TI0/d244ZXslsDKpd7u5xeW
HlGpd6I6Zhj3yupvF/BXGMOH3Zln77gd5P3OLM8ejo9Aj4adsfu1tDMwUGQx
YmQ2IqROAlHfdkdmHd3pt6iTqykD7XhZhaONIV0tFpxIqlPxPIoq95klFyFC
7TTjg0UuU/p7dMsGylNOd/nrPHkxsNs1d+dvncAGfEpVEjkORPd9WB9qZrgn
UdzOBgzozZrL4fEIpHar01h/j6glcDZwDfVUJQy5qrdnB8e0Es6sobIeZAwg
REDKkSR857yCNQb52PXsAWr8LYn2LqN8yfm0hsOTiGKnxEwHZcNZQmHsfrwn
GG/JjEfq4EAuPwW/OOw8rJRp0a8S34Om5Vui8fRrHZTpNVE1lAPf3WkIm3rE
62t0r4ciJcIoe66ADYmMs/I72gZa+k4GBJW2iitRs04zE2OkMpdgUDg36Q+J
HTbXfi+L01oe2pbB/p1oLB98IgD5zl3AiiMm/Ku1aAD3x3rp0YG18glhgCzk
+F6rIqDL52X5+dzGMNXfv5hTjbIM11XQsfh/BZ34UDo1oIfzuyx1YgI8+Tdy
yiFwPit1IUq/ov+/b8nBn6jUfFFM0+4UNQ1hfKbTLx+/mAUkKtLKxZI+6fqQ
v4mIQh5uv5178KpIO37tY4Gr0mwR8vNj9jxwhrwhhxCaMHlgjaCqc/g6Kctl
8F5lOhuHBRI0DtIliq2c5jLKi7mYKK7OEsG4P8T1sVYbDpIcTAMPObrGkFma
RmMWYaZ3vX5eqACa37DqG5j8Nrl98cGMYxK3yvpnp6VSpv5lCmt4Y33EO7em
VjakHRiUAm6F5mI/px9uhHPIrWOavUTa7iIRfpxjHbRqeNYoOU0CICkdCdTU
xaswfJYd9rd4cTv2kbW03qxrZM9vlpFTdcs/MO6KWILT43ojrJWiBf3A2T/z
HrRyQiOBEmY9mz93BLZ5/uLfGj8lz05finZ2TA5OW+tcjWHFrCpPx3xS26Sr
Ijh8YKphwUWxKQQ9zIo46bt6C17BQjL1+bZNnqIn6WQXZHmEVlm3qIcucUBF
S/RMsCC/v3c2FECxhrlL4GULOpnBj0qo2dJudkTe8Cus0wRU2tAqqJC/eQSN
C24yrov7qg2nBbTaqTgnEN/Dcx9CtAIJVm9bIKsnIiUkDsqLwRcjGOL8Q+OG
5Ze6lTiSv6eFOIheD24IvoHUVYQQFQznYvNv9bpXn96yzlx7ZfNVABSuiUNW
eyQdY1jWeExzB4diEMM8Gkh+6PPejA9LLvpzRpNa6wTY7Urb1D9vAkUHb5vI
MjdjGLEjJrI8nMaANDXwTqSK0Y+eaO1Z4EyM+Wl47EzZmv+ZQIlWwu9mvoax
xh5sd1jak+khgeKAYN1JE2x70Au7dv9GYX1uB2d2b4YC/T/BYYZxFUTFvBfJ
50Kf02obID60gwVEX2R0jyd7XBd45a04yA+wU1ozk2H7E4A7S3ZCsEpIphEu
jFr6Qq5I5KKi8NXsxVxzWJXTa1t5yxR2aWlonQDlUODi6tZTW3A1WF6QVPgj
9vkw5HaSh0Rd2FxzaQuOPZ+MgiZxgeUat4QxtPTEBEynfrHeEpXG561RRJ8V
anzPE1Efhw5uGwp1iOclnEpwgYkN4t8adU8fO0ECviOrFFfp7TyTVH3Ap6qn
VPa6EQXbj6VAcFXXcZE1aqDeBsLR3M+KsNHZkRnCu7Ae9mi2ce+Jk9QNc9ek
guMKehDpbCW+cHkGdJN4XIr/syIODV6XriRZpwaxjPTK+vSmTNHRtZ/FlKP/
F1ilSfCX9AG6FgxWMLwzuZQYgMnU784YvbumAe4IqR7/fVT4DEnYwXkX/Z4K
HB7qtGM6ELW7qEEjTF92TPaIg87QDNhLRyC15QQy+MkZEbQprN2GCIh0xj6y
V3E0vVHcEMhmAHnk87LeI+yeF6ECDhRGUvXrwVSyxrQI5o1arkuyWyBcmKAx
ppT258XN/IipA9xoGn/Fc1YS0n5nzA9bZxi5vN6U9SisD+xnM77byiquSrfY
j3Cayl2pDfWiu40zxnTH+RMwBGiPWPtjOSNyfVv+W6lUr19yhXdK1xBZ9QsL
HWkMIyl7yJSnhnfvgjP35jhFdXLQ3JxOr26f7aP0qcgZhWtkkuvAeSICW1HB
gUWJ4P1Zf6lnTLsV5dMTEKlZsswSayTXr27mRIDzxECENzOanVRj9guODJbj
FE1EyeNeviQ8xo/uMFX5DHCKFcWuGNkFElnHMKiJ6jBUSliXarLyPYIZgY9/
GYMoa8pF0moQRoAWtygVAA6gX58D/GpTVlmGM0pJsNgnyCaVI0eZifW6GsrJ
73LzUhtEmBey1RVgAT0W5J8yw9VLj63p+6VlV+VXAYnWguyUBbLFM8flU6Zy
zZDwvAONiEUcbkct2+4Z5tmt5nhxA2oSJEqcNNWpGJ1AK1AVGEjcwvjB16XA
mk0xs6G8SVr/gY451gmj/AtfHz/O6ynOOZfiIToTVENVVFdwHEiK5m9C2Pk1
df2A5yPslGwdHHnRxi4Sl6EYPSeVdOYZC2/q/4ncgj4z4Pgxsx2W1nbqRkyj
EdMVN3yGN8T4s+SzmgsjWjC4Ko97Jzt4f6aKLV4wFiQdz9u43so6ac4FMcBE
ERmjnIBPcUs7fMZCEXkXJLUzSMUKTDT1id75oJlBp3uIoGCFOir3kY3b8oRh
XwW91Izy6sANK3gNF1SCLKXnf0xVLn9iTnHkykkSpyDMprP5ctIHoobjyZTY
LqQI4Z/WCKHzsc0NJeYqgP57Ul26U80H5ymw00FXKKQRvLKyai5yaytOQ0LR
QQiJfcGWzaSakQD72NIrLWBUcfGJlHn8WVjbVeTtklQJDbpvyQUHgcHKllO3
rgx/NTeIf4Supdv+aLYHWNjkqibiFB+OaVk07XIK5vBD0h2BGQh6ZSp6Ynx0
+vZ1XS0Ev+sSld+/pTEvo88DVPb5wsvcJCTnW5sbPJOfjYTg2vbljCKzrLbd
aSdWZjHqcrqSRBKQpnG/6xVcC10V3zJSW24G8oJIxA49EvNpuq6g5pmZJG49
9UsNPF31H6CjGCiICBT33QakSaqWN566AJHYExt3nok8iqoLIZxhnslGzAo+
F0X7goWt1+2QOdhVl4OoPvTP+QWWRuXeNEodGxK5eS4CJlkxsfAmWJFLpynR
pE63aXA+dCkPVPG9W8z86lb58hcrFEYAv6AfvTVII+231i08EnkcEAgt5pz2
14pjtpWIYcGHmdDScfIGHlBN0KnNLWN4LoPleFuaGhutp5S7WMvBEJFCiH5X
c5IbdhSxPbeuPCA2K63gmozxOtUq54saJHwuQp1mioz2cg2LsjXnnut2NWoT
5i4rqofOIKkW7B8zRE0C0y/FuyWhgTN9CzVMZFyBX64qrrmEMkaqvX8QKxNX
aG4uLaj+qzCCpfMNjP54MCSftPJCelg4egKPGJ/sq8pIfnHIReGse/JAMWXG
IfSywAXwxopAP+6xJqBzi56yHWe9QKuQpnguf5+5JJhKc6X2Zo0XaiIEPbvE
qlOxCJPoVDVKexoIJGiQ+hrrRn7PHvgY4/8amXSJP7p5d6fVXP3vHWzFv8Rt
dzcF3FqE/WbYy3wIVcYkjSLolgfZaEPT1PxhzU9UBJOOUiDq+gp6ZrcRUbJR
hM6xDjT0qXQThFFMm/MLJUaFbZGwap6HrShFy+tA3pVB0ftW8Vd2Xf7DS4bf
YG5H5IdTzXt+WbimbKvMexZ0y1lAf6n1xR0wr5tyOWKahwNurTSEMQ6Xiz8j
QMKfhxVDX/Rfn4rr9XS9L/gx7I1t1mHDierXTLXwfGocY78cE4AK/NiPORNX
bmLz9g6flsaB3qCNLt8DgYDrPNoICltVO7BTfwiegFrAkL8ydvq8DjB2pGKO
9HG3IcTYIbwWHYROmCwgGyWdiE3EqoebAxduxmQC1huWC5KKSDKijy60V4SW
7CbKRWIw8eGuJCG5qv4l7tCMx8XzRzUtpHozPns+xP4U7R2bX0ixYVGT+XJP
WR0jP0o7UW7h8Qodg/REZUFvwUIoRkuh41EPTs0fEvzhdYAKWxbGKbS9eGHY
faFOqABJVsMQjfsWdnzYaWrxWusc39fuVTfSaRAFz1JqeKPAGXfkz0yupU0N
eKkbPNrFPRyIKZbw0ehrli6cBJHEwq5LZ1TPlIG9M3AwDT4lUqqDaCjGVHwa
eRdswmHkQJW8ev0FkoLeNGIrJS4xh4FTFHiXWdRqhPnrYnUzBx3kXigHKBHE
6kdJuGfnRXV2v6mkBNETyxun+vaZsp1Wi7aqrcRp6Qvs5Nm5jGKnqck4Y9Au
PAjv38wDIjg5WHKzGwaamKINgrSytoQcQjeFN8RODqCZWnW2rl2y6ySQreJm
TgC23+03Cdi4cRB8Ascl3Du+hKqSGjmuI4DXcsAeYysnY9/0YaeMvl7yd/zs
iQOrgnqNI7Ffs6LoIEfZY15dkcJgtvTrNqLN65U6eEPlxmwF89VLCYNrp15R
QJhEVzgvKov9tqJoZmQdn3FUPzjj9zVg5uuS29rSuGUQrbfAS3Fb4Uygwb2b
X7UmQWM2Gy0/1zv+2LUit4mMPGVH8KrFEue8PH5eWs7eGnvUyQgPniExTDXw
orqPcLIEwvojZ/6xfon0W0th3ldzXx+JbxYisanPIeYVcKPze6VQqV7rlPCH
llj7D5aWIxL922vI9TOA/GEEx4LXRaStL2uDSGTb8WhpjAqQE2+h2c/f5q56
7TOng+gs2qKZVcGU2c+zsonjE0jO7fkDSNfXteJ9ovGTLW/sB1e6broTMTKs
1XWaoWuzaicVxWxWfqcLAXOWKsRlyTiocux8YKMdVie1zSSTPxz2UG1rRGhn
Ej5I2NjR4mk9IsGmu9BphcfsV7k4eIYN+gcdJgf79eZr76x3LeJynKijzVkW
M9rLsqiu96cnw+tNWVEYA+VynGIqc4e7OPzOPAsi7utKPKtYoWo0nal2Z8c5
usdWucppuFH0E3gmIRxAWaxQhLIbGSvUMEwkJTAyF+58wqFNWLAtdxsxI7cT
W9N3pT0u8iH9RWfas5S3B7dNml3zVOClnxZn/v4UNSY18wnBa3/pz3dMvG93
zKvAE054IBpIZfpmro+O/lcZ6kAIF0zCV0QbkTgltxdd07kkj3L4MfK35gM6
M6ocLrvcJH22EZXQijYtTmTyubGLbm0Wy5EYzqE1TgucnkfYafbstzIdglK8
xWxVBFTgo+f4KyScHVG53ugXKvQb+pXWddPtaWSPoDUNLxv375QYqmI2fQUV
u3/72aU0ACno6U/BkDcaXUUhlG2tlufaHVISMxtCsCdR1Of0ZGna7oE0JKkS
jUGT3jpAyz/vT9/yyhk7uGwqibkkSVwWpRubKYxzRk/Hbl+weDnLnhiH4CVo
8b3rmGGgmN76Zm/13uAZqdMSP3AwNBtGJeOlXyFR0KCFS45Iwf1mjhOKtOyn
YNQiSpecFamjQplqMMENoMbwoytsxhMyuqT6np0krxKHrvqWC8MtlE4S8tiv
Lyl0ntUL8xfcAW7/GiY7R1G1KpIhNekglb+ZF80HNE+0/GzIFtiuey+1UWEO
PomNdpjr8DWhJtf8iBfxvFp6Y4e2S3Q7BoHlNLeaJaFSH9dfybWUfC/KUpdR
8AmWx5MjMcHpCnvMKjF0qpjkKa1WE1w8iDUSy8KDnVCbAMSw/2Am2IwY6bYA
afeU0MFgzTFRWUOn0jJr9unFG/jM1ukGOcHwqnQ/qwuN+1l+LbzOEgzfyPR2
ujuWNY7qq5X6gIiawps5KN+hJijcSlYG20vzBnjnzXQDI3yvoGqzZkQS0Tgx
0lzKtSCI4C6DCVaWk3UDTOnU4hKXlqlPXY23He9ua3GqPRAww/aea9+BK76f
j+S5yhIe+pqQ3O1ev/M3pDmX/lPf/IwW5jzX9d8Lz+7I8M4Rd/Rg3Js52VsR
JDdV9KQ+TMnVZtbIr+OmSg6yMBz5oq56qNslfyf2d2KF1xJTXu02O4eSUiK2
R3sGigvftINk5XVVD/miLITwnRbbrGz9vFdBPgSEm/0JJ+9zDNdwMc+fcd4+
eyL5qBReTs2IlqpGR6obTAM3sHxm+eDn2BrisFCNLByOfzzYqrgA+8ReTVFh
7eTa+oD7GFl+9VvINpikEE6xKex20FYeY4AasuCQ23Qu/zWPPM+fBTt5GGHm
0mBhgNwSMdzcgpS/VPR0ByZC9SdXbQuB/1ZgVwBoCJXowUQI9qP+bGL+9yfk
dHz37tGqgxkkZz2NlHgW60gysgfag/I0tjmeMm6W+RkxQB2ekz1MKFIm0ZRc
7EiE8KGB5sURPf8DwvAEq9OivrAWjz9AEAfj6eYAS+UBmuqK2tGCYIT/9Zk5
gBQrJOnHfCACND0ulnws6PtS2zaC+pXr/LGrypdk/TmzMezO61dj/PAFPqc6
e54c8PKb0tS8pNiT+tReS0aefJ0TlBFp1YvIQSeWcmKJ6uAjy3FMMPkqObvt
3dAN5+ikcr60U8L2ajeNdIpjwiEIZX9C8nW7zwKjCts5aDH4q25tPYgthmsV
bDCGdWRV8d0RhRuQoVFFQl6NRcS9z2t4VMYmO56zF47boDulEbpHS8n33Bky
LUeROt5t7k1b+hXA9VoPv5FkCXeq9uk3mLNfxkY2IVJCV0UAaENB7o0AqfQu
Uefk+w7xx3bwHJ9pvV6+PedsqJy5SPOocfEWyzW1/UsispF9PEO/dI5IXGc9
M+bpT5ZMJ7TaI92cSzHgFGyBAB55dLwTlkB8E+fVNQg/XR+kTHd/ohsBhkrI
TRq4BmkX4/XoAm9rNgHwGoBaZEyVqUkSfkM3bEotd5upZJVlIacIuO2VavqF
pL6xYfd45X9YTsn3zihF2WQWdIgU42KvXZnnht9D1Q90NREINAKKOuLiqqRt
Epdu/wYOeipegjgo5hc4BvpcliDq6lEIlx99thnsFZ33UP1ld58yGl6shhH2
zBehion+KItjOByCCb+cbEkoybpAZ7+580TrKb3TVQIuKMMITcfCjmLiQC5X
oyk7I9M+KQflw5PUPdwMi23ne/Gjpvd/Nd5rYAEKwj96O/npXiv0X9W3PY2Q
1hnSqAVjwHt3oArGX41CrT8tcy9Ug/+7x9a/Nf4YCABP+gDDF1MEldkDNBPb
XCUs/JKrlJ42NYyVUYyKIXTxgVDB6sDT3wyPjqA2zKtxS9D1XngrXYu1VIcq
83EJCk3wAqM538vzmgxAGgltFNDB6kSdmlreznrOJjaPurXriJ4QeAIaHbUZ
vfX05hIOZ7WenCF1XoZgNuzjOIVgjVvEcQLK79TgTYKxASLmO1rrOLHBk+3p
RriNEJf2ViEUJlKBnbhxUTYlA4mPaHh1kkfP5HOQSFss82gbwXGRfUXGS1gy
+NWXSm4KbBTDm12VHrKmYO8jBTzpn2ZA3+mpEy96XdVKVrx+I/XRj/qmuLFI
fnU8H+fiKoeKvGctGnx60PPzqLbgU+5aatxYDGDDuH66GPo4KyNiOE0JLp3c
Hz1expueQVwcsbbh3WUVu8dXJs1Ilh1tp3oWpVd+hXWySiNbxNud+4CAnQRS
VjDlJMicQ5hfLRNsNRFVVX3tz8nT6XZiMZFm1tZh74lSMu3tuS7racnnYudK
/R/0GyysvPxYgFVqZ2I2hyehI0w/I3itVgu/eHwaAAdQ5gavLVDuldDsvr9v
k/5DiPrwI7zpN0WfPCPMfKF5LhlRyXs+aRV+nccNVVwg/lR4oKrHBLaWc/6O
gJYf56ZzYD2AB8gbY356G7MEidxfE9rFWyKCFDMh8BK8pvY5ZqL2020YNT6e
Xsu/I485PO0oSFUzLm2DCeS42kbWfkGSGj2Z6cLjDQrgFnUv2uwS6lOP0MXw
Qd34mkYzX6zO5+OW1Fc6wBS7GXspyEV0udT+neQRGzwGZR23I+x1UEfBVpGM
kAkq7p+hpYShUNRSSblAMACwJmXIhI9zrPJRMNpm6vC3QSDSN6pZ/Ylbhb7u
iF6LqJX37H5wM7YdmumTzdXDIGWmk/Uf2UQswhREtmIV4hH3poJwmAJ43qRR
nygZiHK6POh41SBNiZ0RAz4jYAEbFMGFGUTLJlCBCIsp9QA+YJrMUq0QNiuT
U/jNzbztMaDGY/yjH/3j5HYzVVaMA7OGUqEpXgrXFzgZX2JLEEMgt+uo+m5m
sBEMbRhrlyYlV07G+UHJVHLp+YukmWfv+fiP4mdKq1tsT3Ryg0+f9dlc7JYS
dYmlqmwmiK15fRUoKqmGUZODP90dJCmjG3+JIPi5RRqSK9Z2t6VtN9D/12hS
bGZ3JprujZNyIlNbM3lVTNjtq+K9GzQrs4W/3OL/Xjg1/ikVUvkBO96MBzzK
rc0ubg/f0gLW2HVbUZf9YuU6nB/UrbF6NkJapbepsApCfX7i7o7apX6cjzKm
/cofowvkvvi/J9VW9tVRXAvm83A2DzWUf346Z9mg/UzHqD/JUQb9SJOLEWcT
O0SqQwLJmVk4DK+E1MIsG8WcktptntPzUkMLRopu9D/RuAefshkuj/dx9qM8
V4KMACviVqr3dJJCMiicmmyamrZmmY95lXIFit5Abk4cFvMB7NICFN2umMp0
b8HIRtvua1oGLJ+dXK3VPrVjAb0mxgQq/p98Ra/Udf4hFQDSt9/5j+yrvCnl
3XMzL/BFs8w55Fral957koITIe0Col3NZ0W2pAS9yLK3kVA1I5Wj3MQRX3Rh
qGtqzilsLVAwogGVFf7PDZHQ/Zkk0waeaNfYGiN8T/JFtdzfz71zUspoMpB2
DZblB9qQ0zylyMMuuvz1RGod+hRIyJfCiy7yXbFz38T7cAp2nikl7/CXAzAp
lZIMNECYO5FLE2nFEbPoGgA3Ks5AvZbz4FjdDCNe2jmr9Y+XddKJWYTOHkZm
ko6KvX4aQxNGalWbIdd4hoTu/VeSty+xV18rU0+btycLXJ7+ALCVWVvHd9Wi
0SBXaqet4gk36qhBU10f2CbtnKspSqT1ukQT/lMx5iemHeVaXAlmxrrtP1XI
PHdMhzLxECR/zoNcMB4MnOCtiIUoh0j5wP00QcpDXW6Qgt9IpzleBj2V70H1
wOul8+j2hBiKg09+hQZtnZiWvc+stPMH3McmoxS6149AmjTbE/S1JJqZvDDD
gx2Opil1jiJaTc3ngzzk4kSpt2HMe/gE8SphH8OtYlr8u5A6cUiZf2nupaRt
e1MwD05lfrNhRx+GgysBCzBy7Vn3CW9H6Rum4Y5fOXxFy8Hx0a7dZgvS7vRF
g6E8aEFoXdgZJgeiMPTyoP6Vh1Yh9dY1jNVUyuq2k9bqmMmjNkeC7U5Pp2XF
ZU8G27/T1+8dywyH/76k9v6jON8yH3qZ+czURYbLJ55r3S/k4aqs+XRwfzNV
a/NwH7PWCOloqe1rE7+NV8FBGlblMA5BhuOTbTpf011LkYY07/PKtw5aPeUA
NOVRgcxede7KsdMffoLdL4RvAVmSQ1e4EVlwjsQfy3kI68GZOcZTMbbAPYak
YMFg/59bK8Znqad9h6CSNXjuhcfr2YZNzKjPYZ5JBB6G3UAcGb7m1YKvo3So
n5DjpFO1uw6u6cc9uSDHpI3P8u0rRdSPg2b8ePVTKN3po19mCw8j/rc1g8Bu
tHlJy0ux+FtfKTY4VPOFWDAUkMBwQ/ILzJR8tUbmIvUvKTMahhHVITn1uIzk
wivNTKBp57HKQs1QvCNKbcd6gJRfi/HUxyXtdbBXLu/YxNPaYeizUoScR/Bn
QuGDp1j8vLa9oU7Z6EswhUqKIxkgLhAz9+orR63abAhgYUIlSpa/SEoLLK3z
MUwEEntx0Jm3HvS+d3fSctQfes8Z/vH9Xd74VqtKD6CXCSNql38oJDpY4gvj
X3kaXcDsQoFL6jYJYA5YweThVTCTB+3J0FPLNNXSROwc2JTYdlkFX/J5fkKF
3VMZIUsgaYoKu/zPzegRGecOfS8kKfYYI2trQJIyoMVUhkK7Ejwh9QayUdAB
yo7Ffb9gZVr1e3+8os9azRRAHAbTehhejnRbNSiBZhT1y6qpQQ/qqpYSrwnT
ipK4MEdaNyuFjjQiKkE1o3GSQ4CjO/2K4eh4idav+eeHi83ZyfPeW1asgS0Y
7UKKc7vmW+84tYhaO+n7IorG4L7RSMe686O/6vUlNF+T0eQCakucQdrz/v0+
NdKP1lsr9HDBsMs8CFjOa7Z0kZJYl9+zBuSz126d98d9J1KTjhTtB+cRxMMj
RLMhDdf2FP2D/o9fl0MEKyJStGH9jkQC2ks4EaG3J0tQL8cUUHVenSab1V8T
+Kh6rbFq9wwI/RBYSCK61AjS7kASfqtGdnaU8PM6oMVE/WufIj7+dplNm0NY
22UinmqzpMFI6TYHrqQ+UufPygYg1TKklMrrm5zIjAdNBIUksLHf2Mf4UCvo
Dg5rDuirOg+c54BrJJ6ixtgFB88ESnGszqCgufOSB9aZ8J8wnlz15bHMngVD
8yN6P5urC5OUFSxvyRbUkoUJ9FpCAZ8xU69l8Ya9uqIo01W28miHrIfrtZDc
sL/1nG/RaSr60M7Aqgkpfjpb7MmWuc6uw636qUDy5yxYhC/4PljfIjTpjI1O
5Vn+GtKRafAGWVDvOIkOzEd6lNcZ6D0eYi+IWOmZmPhD8sSo8kWwy5ARj8ui
zkpnJW2rkF0XNz0puKAzD1bSHqxDX9HBM4qNhD5qdKjj52s3R5F0doFVWOoa
Hbx9qYYaePCja3U+EYjJIlFYjXMmoQSj5jZOefGOSw3MWyLKh7YrgG/4u363
IMBKNzWpAlD2K7FzRET/argn6M/+wjzfUkjhxLEN6tmzYkqqceQoW00G1ONf
j42dtEDPA5YAR1KYsdTzdem+H+msWECxR2EF14XxiOhkl7PJGk8w2/m8z3k7
Uzl5bD27KHLv5oM7gOelL22RdF2UQ/4JlE0umASQQkifln7aTDcwgc7oQ0Ra
AYpbCBekFueIY8kW0y4DmuKSERMjk4udZT3JFKw8v51EgZnOBRBW4w4YwUaM
XOkTXO7mnAoL+xxSVDn0C2uXCISEj46xgim4Vrd475+thODZQYqF1xQNet/S
o4GBbvRYmKn9mtoxqGM1fA3JnRHrbb28vu5M9rqXd9W56DT1IRNhtDUhHKGL
ReuCUvgEN6HvoFPvvqPACLN2stDx44mqcps5SKxBJN4xGy81KzQw7zcKWSi2
uYeG16j6nFWIMtmNzLmH/3KOqdYu1n09y/HdZkyjfJfFP0SZn6FgTxrJikyc
eLR0Fp8AOFiusAaiKgwzYwJFdAOOKIUuzLJKa/XKjQHqcSL6ZOQKxFh8Pudx
sr1WTS9r/+1dvzEIhH3prWWtx57MnUQIcuLM+ax0Xr9WNbBzdZatHYLtsxbW
CCP3mPtxUyCQ3dDmomDsx/YG0vgMjYNKRvWPYC615iWNfxZ/DyBm5tx1GKVJ
FR3B/l7Z+3J2/KX308lMnf6YVeZfshaVsuwcb965c1n95UjaUdBq/n1X1r8A
sg8TnQFzdLkqA6y3eRkFUXBwtkiGdm0m2Vapsf7rzi7SoscfGpNGpSTebhmT
zdgV5luicpkoPQhh7uyAuJv93HsMANe+HR7lIyQuwR9ynqYVZFn6uBomALXn
B/6mHTYgXHGH+ddY8IYv/UXaPY+sgop7GTVzh+gGxc7n4UbkD35ga/fNG5dx
7TJeZo1OrxesUAyGNVUQnJMioe3gIjE0hZqr4CzH07TeQGH95MQ1FsSLmh3P
31kKevFgEF6d8oiqUNzjz/YC+jM+Mh/tP8zRuLptlixN+ufyEtMeDbW06HGZ
sQ8YfCxePMz725MIiL0Hp0BpgQw1kAYaj4O5XUDcAi7A9ag1l40QXkJ5UlWC
soeL7ofemYEpj77prrjm/Y9KzRRqSP77tUZj5jxNLgqud6sr3tFxUuY4jIOV
IN3hAEbcgZ1wmYj9/bXdFuQUmNPUYU9EwJaLb/wdQXabBG06A56+vbrVjbSX
w9TUVXXoWU5GEwUEI55GxmLt90kx5lErzWi6UBZ/nOZgdxIuF6F/s/B29wiE
VxA7wceEtuzrxS+m7fDrAwpsJTr3FLjCrS3gy+JVpHHaXPLVY35/+JDHT05L
oY6nlFEayVlw3jjyv0MAtZjfuTiqpOiyKiZfYDyQRZYeiiDEutqs0G9Q7fW6
zse4jMwNZKNPHHnnr9fpHHG+4mjLNcqiZmMXgytgZ3CKBLMUF9v1Es0Jy0VR
YjjPrmGatFXOuZp0qP7T8fGs1x0eJk8EuqmHMBQh2nXEXoWl6jU625oHHoAd
qy+TiTUCzOzvMSacgfz5eKdo7siuaL5heixlObx3BLthBBHWg3ivAFqGheHz
ryIimt2F5HctbD/XRN/HxfCModvUjFGsIlVtquKNwuglZVxRv5mSgpTc4+lZ
u+TkL34tZ32l9SMRJY12PlzmFXsdHiuCmsdYGVJn9tzja8TaQK+KC90A3rcG
ElayLDZQmTr+hrH+jb5GnlqUbLNspdMLFgEhuy6GmYjvUe0GSpLrKDYc62o7
g3Dyj4fEvoIguIHO3y1zE38l3iz/4dDMoeBC5Yk+c8E4S+b6x3pIkHz4l8UF
aaY/qt5ko/to9mHyt6TmxE4v28t7mlycksKolt2R8fisoEwZPqMw8Nd6t3Fr
DL7gT8kA62t/+fIFXec61VApJR6yGPkFZ1F2eFCBVynOUNye16LLRq8X2XqT
SXxwXh3JDXkPp1El+aZ+d2MAPu+CvsI9t2twJQsmzNmNOyNhbN/pBoOD9AMw
nSsBin/5ItSG4gxW1jZXTgKm2BxnXVPsXoo4f7nhwhMk6JWlvRf0jm1SC71N
2tPQ//C9XhO9hwDXSVnMCtcvJeTF1oOA2HMRliXV9fucmiytm3NsOSoa+ukt
dLiIZ9BxIW0zkExF5CLpbCwrNWB1JZs4noVG4VwD4a5nDfxoVGDpXktYCAZb
TLJeWh4v4jpCoQTsPoo9kdpcIjBD1ZkEL/Mr6hODNeNXTl71+OFdEr8hqa5O
dfwA8h5O0dZjqhBUi4O0JMI9QHVpm10N8eU8+tvyO1hqIY7K+C5mamhNeFZj
lImRPKpNw3CQUMoefq4RmhLK+sv5hgxxjDhLifupsildzEHDBoicx7qfcgWi
EbWq8/CMg8xY7mV3thSDglxC1tAoGP93IiKJaC5QhfKEbVWTu8raJXz2k0HJ
pAoRxG017/1iWnADA1gKXjqlZYiJ5B4VE9JGMVh3P7zXKFnF6Q1VZhuFrGHo
vXhDqzNVfb2ARDID6wU8+VX6BwKMuOSMG5T6ONDuIsE9RHUAVgIhwA//MFrD
dj5Nme7gzdp7t00Lqs4JsN41lwrXgVEh2QgZvHVxp+FDfYMcSeT0dAm9fCI8
DTuboUaFO4ZP9PvOVKrQuqgk9WyJvWpawosCzcLown41crrpHGorlbrPcPPW
M/4vc0Fp68t1BDulHlBPvpJ5X5AA29q1s8dp75DfHJAKj7ZaVi1eVF9dxZRF
KX+JB33HU9G4TK4eJL/IZC5KScByVWVeDPNPvuNCini08sQHGxb0tGAEZfi5
cvfM+nV2yuCLcwAwNzWXw6VZwVgk13JMIz+prjpAOFgC/inJ2sNIoABjXRmV
oivw8Q4jV4FfSyD6mr6PZ5sku/bYGeZosyNvNjjXGW4FO9RZ6mEI7GNMLp6G
IRHByk0XdF6QnW9vzDGkilf3RuJgbnoS9dfrb//6YRuMMjfLufNtV+5Ng9RC
dgMX5o24AOdDoXYEU/K004glFH00oXJn6jSoiTLfdyTusQiTjBIyd3Mzjwza
xYFodRsYO0ln4GT8UUyfDN4AmOWGACX/lyK/OKV90xjUDI3X2yPackKWAbev
g26fXGW4FWVL0ar9njHSHAotzULBqpSMmsuy82t+3ylU5PnWc2IZPP785FPd
+bY1BRQn9p5T1Yfzi5osXP/OxY8QmprpmQ74QmqG2vrtZaBL5FBdWd4T74f8
HfdwB778+bR81KfpIrYCopbsin5sHh2nHclZ43LFQQwHrfhPJ3SWgPaqEqeQ
VWnJcZc56OGhklaGgSg5gHxbI5D8ch+BMo6JgvIfaBQHf/g/LT3UpFTQHIS9
rVqctyfX3OPB0GlKxLwNzJoOIDArtCfKAmk5P0Rg7fipWfjlkgf0etUuwP80
HnfSxtwNxSnI/rcfk8Ebrgf4ldStjJqAeH7jjk02vcDG4cggh79+lM6d2cgN
KhV6n6ABYydEVyjXGgKqqjQiPHBi3P6CWsNzneS+VvcXVpBBmMdlz87Rg/5G
Yuwu4VqYNU+v75P2j16X5DjqC2Cg/gmma94sKPd2X7x/UhPV0k2H4ioH2pCI
ufEFVFLuSkZVmfEpV3nvEsQFeiU4sXLIQLci2e8YLRqHNvcaY4ICV+e2Op0r
rO7YhSXMQDBcg2KDwSbSWxdv24ua9OZ2g/bbUcXSYIax4wHkZQqCb9vrJToS
Qhy3EPvxk7cYE8y62vIL8rAnA9FrH6v8FbP9xq6+wxiNZtdJVudGGe57y9u2
kboyB0FwIusjyZxFsaxSkQva9CnWs/tlJcuzhbiVGqd73s0oNK5HJmX7zLqK
L7NqIkemboETBq31WiDr4rbDlAJHv1lmxEITTQZf3RbfoY5XNv6GtrU6FMQ3
by9ZIfCYKzqHLHJGeubFaC+kFu7GEf7TLDcZGvVfq9KBcimfH/47+Tdl+NqO
xDcBn+7dZiJ0fowyT6XOSEOgOUEUeWZlZLo0WlkihWvprLfz3lQDkEuPBeg+
/CV4fykkXoCg12v+y0Tvispzk2SouYhRt5/gCoduTzGeYVL6ckbvDWeCtfzd
Tyt+6ERVD2EveAqYTdkpXKnSurvIpfxMO7DTohfC4BYw3Pfg46q0bVa+f3mZ
8gozy2uaqY8aT0Pxuqqixb1B+2WUky12N69a3W+xwQBYcp17KFAhL4T2Hm3C
qy8NnMp8PIQl56rVansA/pK18tnpNvWsE3Zibnu/dIHbw89E4QLN7yep9Xij
CZSloXmfNeQ/UhWlG7QHAywsipW1gQjbrtS9lU6uVF8YOg1deEwjW8aVFuuW
S2M7LXyo1wHBcyrAGFenkXaLUUYBLz5ghLgYzeZ7ELmWWUch8PhSz2cLKpxT
dCMPyWVHblf/TV7fTIUfU8WZUjTzTDnXRUZ7Js+VecaJsAApbsJH4O5xpylO
z/wjoRo6kJQIkQM2QA4N08iS1G5RJe4Y8h+J52BOHYvte3Ld9N3urifGRMys
AEc3vxwhWisGJpMv855ywZM3Yw+3T1/ZvgOM2dsw2fnoeLMe66gg0SpIuh0J
vcmUre8I5mQlHVre7vQyYdtER2etHQX1QQGFA38FcZ3VsQ6L0yKiMniklXrx
2uT9BC69q3Kyl9y2sJQSD0l0JXfrImBm2HoNf981JfhbEu2nCdHf6f36M+aa
HZN9fVjAyoUrNQbljmkG8hHIzp6xqCFk+Ji+xVPGr3ZTu0q261S3VFW/U+Pp
hJ8/k90UCRLRfWp30X5VOZHm7rbOIlyN9A6o0oN4K2fd0nX9fLPSYnjhlRdY
2fblT+/suoox9Vnay/7Pa0CES5Eth2r2KNn6/0eYHNN2d/0PsW/pJVUtZqFY
drX/yjJ2W+hJ/vR0Ic4pmXCWYtnZmIIrscCIqHcBGwTGA623Ip/CUXqMCxxq
si/NJhSk7sW+QgLy+SPT3r1r2Ga4KCSvzEOgbhrUvKNj6JcPem4ff171oHbG
7Bj3g297/O6vEtHmrC0uImolC48hDRCLKz7/PH/LsIgL7wneofENZpzsdQqU
9WETQSul+CmqFQgA2jqeF1YUBwN124/UYcLtSTDh6vWVKHlwBy0Lfc4ol/tB
5dvRhNU3Mctxvw3pVxb2nNVBQ6HqTpCzmR0tJoQOHC5nLspF4tg+rpcDw5Zy
3Gc2BbtKNanhM/tjF0XIJfDkQVtD7XOn/I4gIzuPZPjP0jRowLvREFhuCtj7
MqLERfHkPeLd7Ehc4lPJui5n45OOgvy96fmoKwQBuPddOPXEvUIRdarQ8I9u
DoIV6PKjMFySuGJhgXDZ/fufZLxkCZHC4fNBuU5cuOWEKkzoaggCgeAGdNr3
pmY+V+76u6f5TetmSbUQ4NMGpkFBIzWj81s/FT03mdxaKVVBALKxg/1QluNf
h/gNK5p9eCO2xZOpqwZ4Dwyfn+i1z/zOrUiKFj/lO+wfS8UumeV8cU6FU2cC
nXN03nNhpVAJSRT4Cg8Dl8z1/GbcGJQsn0KJD+pmq6jzN8qKjh3FADsyCFmW
8+bEPlbFC08CNRSDIIwVsMz3HwLKyX/maDiX1C4CKc8CvVPvGU+xhNELy+25
QtLbsJoDNqAi1YHhUlh2r4JqPLrFVi8ecffoKmu1W+ooDn38G7lTumKhFJ22
rohcqt5qVrFXUf67b7mbc9hXDdOvuztQdTX53O89n0wwI+irV2jGsubpU0rY
JqDTscoTOGyxokG4OyPgl7VxTP/srUrZIz1EfBva8JyiQSaDPBRG3LxPo9DQ
QRYUduxV8neQ/JnhNPid0kPumbu0H6qX3voV1jtsQo7H2vP6AWDKbDG977c9
4kTsrOj9KOCLPezSQfixc4fd9WQpIH507cRqmTiiqmTEYMohIiY1TaQ/YhBo
wgncUcAG/YyODlaHOdh9c04H7UGV6Q1pdtKRa8oDTNmynGf8heNHA2SL24sp
1AWdcmy37SY6nCa4Q6g+ct1zSVSanqrCgvV2B/CNHbdvmVxMOjW4BDJ5m1sW
prUfyWJRmp6C1JbbxDh2cBrUHCjVl0zvHrqEjE6XkQotDCjTNWbcXvhNvcTz
fbQJ1DzR6KMOlclGrm51Hpu24E9CuIZ7EOqp8tWcNbAe7TaWEjpEpskn8WFa
4Cgt9mH1zzNMUDBv0KKAx68+Umz0P468WJD9P6+I28KwMkfYhfMpiw+MahW2
ts4eeIU2QRBjFNFWyEhh0Y1zw/6SlUf1jceSsJjgJ4wXcj6Ju3TUi9ucDyYh
cJe4UCRA/eMYPyDwOhuI51XsmYwiYa/uS/NSo176DLxKN3knsoaZOOSgBmxT
HvLv0atRtPX5XRbmDHhE7CVTgyDMicYZhy2h0QQz0hDD4FUIXbsLDDwbIUvl
BChqA3aNMrURU7JWqGHwdpMeZ682Cp2hmkkIkgbeYy2qxa5RqcajthSNarhS
1aMZByl1IikAVHDjvujZJI+8jEftKEj4PfPlZy4VBpZXRD77ZMs4pPsYlfmN
OK8aSmVnqRdOELRC/Kjfzd2YZszHZURsvwS8uSmVNHmP1SMOvrPpiHUY4Vku
V7up1YORk2oIsbA5r986IozJIL6x89N/NkNCyzd8dymBwZuq0kUMiF01LZ4i
ZGPYMPGiPM4MiOK6K3cOVWCOHUtGsMrCikYESKJqFEbpFetw9KE2Zba5g70L
jLV1f4EvOXRXNTZqlyChl4d8SnBbzD1sYzDg48pzyts7BybVdh328+52mOOO
M9oXHSl/cuK3L9D51UCX/YHCLXpJxeTZaLasaDiumZCtrBnWRRwKwb9RYRbs
Bv/NKz0tFTXQENqIqHBl/CTDMnKYBXpqgAOaSO9tkLjcXvrbTcR73Y+dROW6
EgaPVTOuymQyIN1hmmaflD2mx3hah5Xa+s2j/l+opBFsNE/heNpKQdT/UDcI
swuwHUYRMWj9j7IEVbPwHb+DyLyyDVU3/s9jMQ85bizwRTf5FDxGyWHG0r+I
a4RmBOgP/GiQJH/ha9+fjM7/H2bQ/5i5sxrpXwKuUK8ck23ihSA65+Ma+ql9
CrE4MJKclr/d07t5Hx9qSLrygtp73151KsU1OE3EESwlZq4Q3YySdz8dOyXv
vLNsx8cOnEvoeOG9P6GJ1msmfHRZ478cEbgs8zmBJ3V594LSW+Vpi5WI8WDc
ZjSV1feVbPVsKfcjV7drUDEG4x0XIu/wPL0UCcpFu5rW/QuWqRqgAZmEmIbb
bB1CV00m9JsWIMuy77wcwQH7FmCfcG0lxN3VfLsXvQT0D615CA1mpV811QUY
5UEn6kngsjNnqg3fyvY+FaQpPKTMzFW+BX1lsUVWkbRR5fDT/a4pzI/ZvHBL
qcKDYGo6P+B/l3dEov+/uWIFwE9wu6r+nvPUpLwWGt8jZsJCNymLEEPFYHAt
0l9ZgEXycjRaOEJB0TPuV43fsZFqwsS+/unKTnly8RDk2EQp58+ACqhqvgMt
xjtdL3j5Wu7PRx+ofQY5TydCdaJaar5bf9pmOUP5WR4EInRmnOEiZhdYOUUb
mARrWV9Szbcr9iZHqPGKZWiZAA6UxNzpbJ70T8J5Uii5vLhTcxaWherv/zjv
A1dj2EgGsUXUt9lC0tbEgL++JxfuuNpsMIGrCB4BhTcRiX7eW51A7MK67oCu
Jd6WpAqeRgSa6nn7Abj+h2K9qECu6Ux3yv7yloAm2I1dRvIANKfy7FmkdHTd
gDWgb54viWl3zCDb6iHCMV7nrnv5v/CB4jSp+ur91fFXXgZ6VMxAaGuNZQpy
A8uWrZOZgZVybgqDg2PBWI+pQr6XzVX7wflAK3JSx17mcEGQq+Mjs9PJ8qCF
uQtkl7GO15SpZyZR0wSCcCZHqLAhA7kgImahSokoKsGmSxiuEXuMxwFJtXwi
qWBVhV0U5F908zntvf/ZwOtBhmGSuLD0WUh2FCHPvLW18GENes4ZLxsOxZq/
deVNQxiEgJ+grsw/ud4FPB3fz5xFWVcuN7SYZEuSHvzWGYEyuEdDVsxy/VGC
roK5JSTna059G/yKhSurPlSV8m/+q8NI1LbiA0WaS9fBTbeVTMN1f0/rUi0y
CCSPmAfQHYMULsPEtcWLP7hdxvlyU2nNJpz6FXl86NM+Nh3HirVO6A3USmlW
6R9gPLHCd8E4t2yRqulQIBts1T4jmnMfpQqI25Gb+sT0Qq8NMADvAyS5mfta
utCBg03WfWUenFAD6YwNweimmrSDmVLk+0YrHh4Uv8v1jEqaphFGaeTSXUcL
rFUZtbKevQaTU96bcchhNaYeEX2GcviEwWk8d7ZwM91Oems4EF66q4URinTB
ut1aphkVCsLmPu5E579AaHO5B3hKWdJcEn0NMgSFXIUBOKRtHoNwoh8a/CvX
3yoiAy4cPviXZOZGNfCeN6b9dx7NAYeTzFFADNLSVavMHXXf912yXJObDHgv
VI25e9PTzMwmYZCzlG+6slwB/Iaxzs4dsVn8peD5uvOBfzRqSEJPDY7ef7os
7sxpPV6JY8ucZZhoE95+s86u6O+glcg7DM9TOLofKih2fxlteyGMFyekrKJ/
5VVYmpq5YnbruzGZRLD7an7M5ny5Avx3Mu4d7I4nThY2NJLgB0k7AgDfBl1W
er5gqWvrlEwZGgEB0o3/Bqxo9Gwpu93WDbJ0JcUqCIlZNuopKtrmYKYjj5mr
vD5p6GOcOOqH3RSIHdGTfiRUCFBJ+yXws2p8gPaaNCcfSuuGpS9bPSvEt6r5
jvljoR1r/qJXZbyd8SDXStDR2UiMxIg6qGXAXzn0r1uaBuL9Z85eyLPCtI8x
Tf4qZ/o/4Ml7DTUGen+l+bhq2OCbNX/gn8s80H4OhLj6hFiTD9d+9zYJpRpX
lkFPBRx7Js1zpg6jU38tlS7uyt9rgGwAd3HXJEbPx6XL9Mpamw0CCxKVvecQ
j7mMhenuvUZJ+MT2PimBEUtaDcr2iOVZrI+vn/WpZvS3XelSE1S41ngX0xrs
fxT99z6y8bStqmxodc9TQszczAbmp1lsZo347MTpM7+xOl4mPdkULUTVQJm4
qSE0bB0YYdqvuKrQlxlQtnQZe09c+0Q97fE/J050EsX2j2bGjW6g0kuD5em1
xjlDudwnOy5/TSko8eilkosolCN+tlCATmi3t+UcDa5ClV3aN2SLyg47bbl4
DN/UaEyNsrJkoZntxW7AyOnV2WeTZBPSOnDfaNNn19/bWX7dohH33aCDkV1+
n6GdG+b6mfA2UPvx6vooekM/ZNLD8QyMmt5qzk9uljdVH2LUpRK055xvyT5w
rBBQwO8SckB0rC372L6yHwauu+NeIJ8vf4gpNXTjUV2JGcUjgYvFCvARh+Zo
TOlF6G0ivityEatSni0ew2qvSN+LkQ2/B3/rDGbe32sbKuHvOFmqSHU23o6d
8Huj3rHTlkdHLkv5WeRhpTHQ2w7Kp1OXLqssXSwyUp5eFckn3lCM0euettIm
7RQO78tnjOuJVk6kB1OdYbLM2eNtOShsCiXhguKRjrC1D0qrUW/ldv0z5I4W
ucRksqgggFY07iOdVbTE5FU1SutFYMM3PtaFQ/VWAexfC5rnI2BxZZvDS+s7
S+fRa7/JxlQMaU9HbMi/mrqCKSsSEFmWrtj0cx/lEmvueJhKs2s86h8iYwde
0J355cQT85Mzky98yaOkQfLDPbCpqJKrUqiOF1fMM0Lve598UkTM3mfMQWp9
BtYBNBV5GtFqDu19GPz1xW0Y1bAMvqqEwKTsF5dhkfDH/yT2MbkLticQUkDZ
H7jP3PwBYpWkYZTt8CW2x+pZpxfNngMY42Nz91tgAsVbHdZ5QI99Dt1hbSsa
LXGETl2cv+jDRihynMrqIx8bQgSym6VXPP0RIzfkjHDNfHB0a39lhR1cNc5T
uKukpcKndHIoojamtmDvrQPqdVt9jM82xZ7qEhyk/qOQdkBroepLyRdL1O8Y
S/jupKGWy/FrhK28Bxsfw9CrQ0G1hA6YX3UdOakK/JOZ/vKW1nNnE0s93N8T
VBxWtzT3yK3fAgYcTh2Mwqw/7Y3bcjVTXtPDSr7Af6IfoTI/DyDwo+75OxMe
MqtxeMTIsPAnvNLcjP2ZjmYCY1oIJcZFVGZi9t9+G8S+aCiXHcNhW2u2nUie
M84Oa1I6e4Y1smFXTDLjqnfWZIlXBttK+0cs79YsHSb61Ml4KF0z/oxiO/Od
+bgzxhmUfAArO2RumOAB+5Hh616XFbuYXu9/HMvB4YSCCy/UEJ7CBelHTus6
/fdagVAxXtfOnwFGDdMFwnLvWw6gw51VCvCvmKQJXpBefPPZ/spxsYo9OxR3
8HS+PJoC/zrw2DYp0HCa8MK5xhDuPjAm/xpjgqclKPfv7JgDUJ+gM3gHDRzD
KIrUOChm2oEPryH+giT1daeNcPyU0HEKiuJd0HcxLqPTTxFAD1hEEjLhTG15
b2h1cx3x67qFuBcb2cp+L29pTTBKQlull9810lfD0eSIuMyAG3GEoR9fhL7h
F5L34PhtQqF1dlNLkxEZxlbBGaTTHvVBAUTdk0lXVTr09jpCOJycCW8wirzc
3cI5LBwN6OMPcz3mJmfculdWinB1sJhYInVi0BWxWbDrvfo0HGrIO2BRktw0
2FxljD7WQYDYUeW5BNfigymnruNKE3FJsJXfEaxDqligMElNsxJrkQ8QWnKb
aWelUvU6bV/KNCbIkdr163kLKC5ekmQOW5EkoTBhrInmAZTIFbdgHa2o+2nD
Xd19smY4zz5gloUWqsv11KrQNWswdDSmurGJG7R0afWTPMmzs9aILH2XV+17
EFp8CDYMMWEtHZL20Dv+z+tzf2HrHCFMQUXbNUKpy3XSnqlMYg7i+RlZRcFB
j2BDbEionKYqQ2y2PMple5A2VRorA6GtSCEVHPc5+zs3uuYWnxjfSbkPv36t
qoTGqC0LmktQLy5FAApBhV7Ze+u1D1OfDciCthXpbe6VII/r5zNeZF4AThNP
xjD1Jl5OEYCt3uDewuKsSiOVp0YUAWk/fuGgew5bMr80TmGskVaqU7otGGOD
FWzgiQiS8uLge7gDUP67P1Z7NPh9iiTwKoJbtrFkDH9HFOboUTpkKolImWMV
I4VXR0X79+21YN7PVIFgmYsjWW4aPsnIEjmH0lf73gMMAqzIsfViWsfszwzQ
8FagZr4r2C9JRUjYI9J+D4NNwzDp+7PQ4pOR4q6jD+5Dq7hlVLfnGXJtfgRd
3/M9Q/kELzCHuLwzOyHLQBR8y1WXX35kCX2USFVv5p8HIzSVZwYZqemIoKtA
9KmkrxJtIFKan0f+U+fVseokNWBRw9tkFJvg6olviNUW2SygCqniC8ZI00VN
o+QULOyAPzrQGt660NQgEHnklKckwtz79CJZAZzR+7tfb+ap/PiB5I7Mwroe
QjgI3N7N/X6bs7tBL7CHzK1gokzEjkVK1sEstnckSnUPzZeVx5Lm6bVgBcS6
62RMtxufrJovL6KwutZhlEKEmBpoVOthlYYSaKhfvollp4HCVSUeP18W6mee
UBHCQtiwuZN457yWehhHrCeZNqY7xQLo2NE+dZLJUnNRv6YqqcwC9KcO05Ip
C0ZAyNpx2+Jh+Bz2ZVGmS35gGrTY9X7W7ws6QPINqNWHj12viksvGv/1lr0a
gFwiL9iqWiOOniMPMahwG4syBSs4ggKLDsjC5MyWqAcMkGUKxjFG5uHJK4Eo
SHt9CyhEIrI1/D12IqrVifmUO/0GvealkbQZVT4Us1n09p/2wawWIOhvgE8S
mUPbz6ARL4ia0GXpXf152WaXsMasvmWu7d9VTR95gm4c3Cl5NEAKrVqzjopJ
Lwyr3m7wO/7qSXWzOAxPtWT93hRV1FYRhJ3vyskikjV8RRb4bb9YW14dx9I0
R+nQB0Hl1S3sUT2teNneoCLH349/IiOLp4w8AKcL/UpOf6xl5r4dzT+EmAj5
ercCp9Shx7b/iXdSz7uTz74qRykAduysZpqzRJB8GS7O3AElzFd92DqqIG+p
42Ch5XcTecSAr8/KEhVVYhRJenGabFi2DedGGKk0qgRhjyJlEasiekU0xazZ
nIAb9x5K7WZeK4/BcZ4lZ9yeEDqXdj9uZwEPDCRe4/JfNDOQhuFsOczy4IqU
UME1ulIw3TQAD2hvkEqk9fvatL8FglaO8YP86S7f5wm3SS8b4yvM/4rGqevL
+l8b+QShq8HOtN2TtQ+cTMzyEYrZV1xBc2FzUNFrXm6kZJ9zxhOqS0yGya4U
HI6QhfU/TsiIEuwZQH7qQ+bQLwM90XY34/wpbzrJewT+Z8RZo4hle4YjUzg4
pbh7Psm940BVTVAfoL8z9hDd3VGQCf8h3M1ZP3mjYSo6S6btXkM1mNGqwwio
LoZUTlJoBTgUlEDBC25zNatK2b4dZJbKNFK6ZTp4ZHVy/dVXhQtltAPv0pnV
RWL5VBOBgJu/L1KMwpE2XAZd8HXXvpWSNwGu7tBm2WBJwbMENYJxsRavy9fm
uDXWKZEzpymSzJZvFdqcrfnuxlclvFZeZL3UNf7KNyI8cfMs/xjXs3Z0MJrB
PfXTCDck5791yx1YZZ5xCYBExJFXg1NZ0rvOck8Q5e7n8yGsMIM/qxEUQdZY
ayI/ARmU2i4T2CGjVoq5hx83oQRtIR3RFmA8H+eek7wgXj/BM+8BXqhU1ha1
fsrdv+Yq0owBhY5E3wmaGccQULmFv8mAwkNVgJET0KT0F7/cfeXAUyMHftEx
M8AuwTDJ2BmT33b/58YD+6v+qQ+hCAfS47D3yG8QzxA6EqQv9psZdlLs7aw0
gZ1n9Je00d5FTKd1HAcuEVUfaM+AXNu9he5ghV8EE57XV5MnmMTWzSafu3xE
cdohHgNNLjKd6Wd6x4q3OGXQx4nDQkRd50+0LkfjtM+tVZSMccJgpCct9mQQ
WvzbqDy+pidjMvd6fYXjuYmlgufwa5Y654CR19PKrKYosC3VzOexVnskV4ZF
aQkjN3XkjXv37ZC2k+CJC2T/092Nn8rs0s6iItfytriT6S93Tr/P+nwqc7U4
x6xo5xwc3vJDAHoRHnmWGy2j+g/keAyZQIPemlF1qpn/LCIP7WQkRaQKy3fZ
dX5yrAPRO/5slIRvPwR0bjN9UVFopA4mk6su5aFmLt4DUoOqtBx3Frp6raCc
u4chONo7nqEY/VnGgoexfL0aUH2KmScYkaRK7/rDI81ek8B6Lxwz7r5kX9Tr
48cNr4twHqCHu2irCciJXDLXxFAimapZ5wInkZ15Q2mVuqUTqarXvnfkBYq2
Dbv2q/JxvKpFMVnJiwHGwr2XfCoLGcy/LJEhuiVvSZWWoIi1ae9MN2IpmtFb
HEksNQRJ9iOLflPoiP+Q+Mt/BayoFdJIfG6LpUcmWj+UC5n9tapQilc50cUm
PzayMkpJeyMQw25eqvKeyQzUqdQK+MLAkqDURnaZvDSuIBchtSsZSWL3Jgu7
d/Izk/aIvidbnCkDxvq51XGk2soYxh5CwnSiz7yK16rZvyL/OSDxr5GSxKZ+
iqqsMSWIYSjIhh+9q/6T0Nktau+Zocy0YH0xpuTwLSXVGT9siD+l7lyxdnph
jDk1MjQD8ouRppvhxZvcTCIiiEZ2ONDlBkTkkGKNdWU0BTf51cdmjBP3Umd7
6znxOsu3hjR1IKFoXMRZ39GDxax8LeRe8NVXOS7KYiIQrPqp5rdmICNUP6IF
9YHPG6u8/VIu+CbxyAgp4RmxRR8mh13DUGM9RkAsKGLpD6yyyiMFe+vcjEU4
E6Ve/iGKU93xcCBiKA1hSd3vF0HvGpWuR4vByebryuBIcrpmLf7i2Uj8eUrB
SlgD8d2zcjNvNmEuh0Cv5r5r+MzhOs372290MACqKMuRp/30SVno/yO7x1NH
b+30jOYGgv1tVxpD6Phn+0qevtafNP2dYvacc1Yshw2OdqkD+FaDoMgSD2P/
N6DKeEoznxnb7nVGTqCrHVXg1fD/JaAqLLU1eaNbs+MoxIzdd1IoujuQ8oyf
8qzYaYLBPfLVGX/loGYq4KsSXpZUJsIbnWRCtrUrpO3fWmhEbExwUppar8mw
q2jne2qoiPzdd5cU34nNMsbOWyX2mTNZYlkC5gZ/GBs+bVXIkwzQkUct6eS2
fnLZoxvJ2r3KufUMFAvxqwLwE4qINvNOAeUAxcmTwFZsftLydpYxvibkSWEJ
B8MbYLKP5HMn8l+PQEVv62Nb6MH+jdajLTUxtu0NRu8RCsA38ONB4bYyIofY
4z87V0Kqzv7Ax7eOyW6neiFYeWaMXKIibAkSylOEWpcIG8DuCv6ZHxlNKqdY
8XMTo4YllCA0aLhH6PwPhG5Ey3HnhUzajewaZT6U8xyd8SacZmjKU1ighmnP
YeKzDZWrtZ2iO78zoQcZOxw6nDLePHjryCpDK7C6XJ+dLpCyY6W0ysjLY4qK
RVhAGP4jtr0WgEysJ53w3n0aAB94JHnYtuyiNdJKWffh68IiUh2lMPyrl6WL
FvouXUdsn1unN2eodmEsDAzs9XXFbSfImmGe3Hr0+dtNfcBjRw1QjBO3jwt7
L/tdw5NfJI8yKWgbuvrmFw7pKxQ2h/M9175hxFgefiCNhtceX9stNCVza1wO
3bNj2ETk5ngbCKAccTgrbZgl3WlHxoQTXNfinBPECuR9D5Y8vApWYSqep7WA
GaIHUdc+U3K8sQznSKvNsXhVrGL9TZVt8kEq9yyuNJEM4ipw0UIhZVLwil3P
Zkm0d6Cict/AhWFwa7555d+GoqCkwKL+tSEC/NW5vY6A5ducC7eGpMK/blEA
UVaJ4f/UhpfMElA3XbHGSmy46d6YW409fSP7zQmwypNrhKsSrBTuEf37PRi0
BVYjWQYYbDddeJmn92Bg2ErRp0JHHJn7QNVE9rpUxzZTffqWM/Yklvi1JVZW
6U4avVuvphhE2TrIkZfYdvWwsC4vbQFe5nh6Lbn7Iwvw1D4IJxVfbeXPEly7
i94TXS06C4rdMi1hU9s7zYZ6gdIHXmyhPuwnHouAc5l+r7HNTpOSTPhvS3/c
Cj52G54Izr40tNVj8GPgIAsS761gnvMwbPP+mRU+W+Yf2m51b6LFZ2VqlOff
V2n6knbXOalPkEOqR1qEotiYwbwmQC2fUvnB5f+rIra3O+rYwB7RRvHCp3qz
jI79QX6rDzrzunxaC+Z/dvx10Z1uPB8qXFTk5t3owhyjM4LBBYAHKSWSJ/su
v7iGgdSY+xbuxUJmr8ZOIehpYFjPbs8XKx2dseBw/Wd4JLRlXKXaCgAygQRZ
vL5MsCGXzaifll9iVcczXq3CtfJgQ6WfV/RQkGZmkr5q/o2ae+d4OjBDDQCa
Ocd4K2DhA2esXwSwQh5sza18P96fiLayrVmJYYPcLflSQkHsEK5eIYLd23Xb
aG5j9BhPbefV7EcwSccnwymOMNX5IVXc3eyWiM2+/0yHJdLopwUoau8RWum0
LlAf5LaouejtezYwWbbwCiSVlc4Bc7FEV2rYzBr3rgRSsHRrxeFv+mwmMi7m
gPQ1kbw6DHjQt1LCN9Ui47hKwO4AIPcK2kWvLwCgkCnYyxfA79O3TEYpx6j1
z9Ulfaq3zax+nYr43u2XjpjgKovhqpEhlc7+SJ5+IkExjtAfkPJcjoBZNGzr
sqk6W6pQWyuCj8fEdFGELfytb6UZtu1wdTs5Jtlmxf+O2g5iTXKBbgVFWGRs
sQgTlOS34TZG6U7nTDFKODlnwQMu+qKYwSEE0x4V0oeF99KCpYopuUjWYyms
l73nAXqUoDfCBwLlxDaNdr6KaRncN0HY70pEkEn0m7yUtFtvvwj8wsSP/D7C
yH0sD/tZttNTIiMuhy9eBwX1JISktngeu9YrX9nJ20qaPbrbNIVt9qkQHiaV
4Xkx5AfDd6FLAK8P9pvJXfRYz1JHk6nUgthnkeEMce+t07QLlXXacgwIliCf
228Ntkka4cTYDtGxbFHah3tFf3pDlN1QwjX/6NsxIoFRsYa0cAB9zPWfC6xo
bPHkWoTsy6aMjgAhQ9xea+/tcoYAOjlvLpPIccHUDIOkU+KHvzn1ZvkKEsU/
b4HTp0AIlawO5SGM7BY+FVAcvkeg8zU1bS2tNT/eiXsIeWdkE+wxHVUty8ge
vPBhb/4dWzfJmCVE6mZYtmyit4aFxy9WeqftXiht/6LXw+402hXFTwX+yHNy
gtMviwFOPAzrp+oK3STE5tYFSebtuRDnSNzOCwn1ghB1r+kSkyIRtb5nUSVg
mG6TK3a9KWJbd4aBSGZO6g0sJJZURwEnlhhrIx4mROAo1PGDScGFM3SKHh/c
unWj5+pRH7CqDZ1Q3B+cRnb/yZbxcYs/QM+RdIAVoMwPgmVfmNRDkychSoo1
iS7HKiKzb05SgCq2EphLMJxYbaSz+Vr4ApCHuQtb9uCYMt+LNv4lA57LOfwI
PEpHECIYnzAwhp2qj4NCfmO8MyACT1lCRYK7k2gOfaS0Ctb6HZMglNn+qZKB
kfWVTWWoZhsAL2h7BWEUznSjbSW9HC5DhXiSpX22QAg3si/MUJFAalmseb3l
fH0cgXaYMWk/5tUevoLhPoMEXf7RjOdWBSWdbopSYuhsmmjQUngJiMGrCSxd
N6wCLGgJcK7iSE7wjSLU3Alud7F10fnOKfgrwgm1gOAiJCULLfF+tKbs+PeZ
eWVdtRdF+aEENQhgsoMY8VokdGyLRwlzXxca8I8UBIQ/kYbpynqCzwFqGcZc
9/S12l2mIhUcxln+k15jT3CusMTsaLJptrf2c4ut7U6F1/vYLtzV70l+/U7X
jBzVp3WRKtmazOCKsHs550o2f1ERoBoqUK8Rs2Y4vSWiGKh/hrLwMjyb5J0c
iflUh2YPkEIynbeu+x8ESsutYHF90dcaiqJi0R9Rgqyr7VGcK/xCelCwyk6X
ORN/zPGxqpe+uGW4Yf3T4iuAY5fuGR4LbuSEzv4HP8HCom2LYXz6fK/iuXmJ
5PnVLicxWgopj+CI161x7clYQyHRce3cL27ZVezfXrNvDIv/SJEPWa0Wdu94
JQ25fRrLARku8yvVyZvQnrN2fxMAvY7iyUEfWX4BFD0gx0mG34O44LrOwHwR
DS3XBDP7DC7mOAHCYIYEdwS5GkfnAiTeeyDE3tYuNr/zPY/dt5V/VUSKEZiK
NL6cKfHlZ1lejreeN38WUEhm1ezgG5JuDliWiZPbiuTLiYoMj8ktwn7O0ayV
XQJmGUVLSddU12QHh0yUF7+EuUAY4fIK6CeMS7e9wYs//5l3XDA8gBbJVPcZ
pzksLrd5apBkFTlKVFg4CHXbGmQBTT5AvL3zEoQke1uQZlf2wgaWQlL22sfk
niLKnqQBrePzSeoatZMqNBHqzVOvKh0N5QJV1smZC5m5pYR5nMsReYmNMVh7
xkf+w7HcRGErMwvGP8TPmpvFbcoHzKvXXx/5YhmzYIVYYKWxHTUA6LBUY83d
g6XzOadYQlbAZP8SfSnWPy2Ksi+FwFdQP1opK/W3A6VATIzPBDUjCAFAwEee
dRBAd2MszvHzj3PVpufg4cDgNsBx4VfyMUUJgYQ82UmL+RlBqC88rlVUuZmf
c8rOMfjHLJCWjV8CcJaHQQwE0L+9BwRsMn135KPNQcg8WthZpRHpv96Slg0I
fwhg1m2tnDyDd8iAxhLhXk4CnlrKXmh28VpQrDykVz/tdfbxtEJ/O8HnxKIZ
JxBibW5c7SCZZtI3Z1KKpN/F9rp0htvAbZrC5R3am7A4cdLxGOw5BsczHU1k
fURaeiry5yZHwEUjogfALkq2ynZDaQ334Gl9JAokjgKjx9McvXyY9rWhQUSQ
fGW3qijGxmPtb24sDIa1hH2cjzrNFpvjBQ6p/pwHvavk9CSnsVIlCqLWSpDc
Nxs7TIJl0x9hUI5ZsJCBsNdll0D0GjawoGO22pWD1DJ/aeYIh94aZsStJMDp
GGQISCs4RHE6zifB9wB/W6A8QDprpuxrzVrYy+d84N6W/1F+450PXiN+vKFY
O4E17LZqyqBt2i6/1YTx3qxPfjrWuHwaH+MQrPzD9cypiA/FWsCKed69VrNI
Gnp2mUey+eJojNYb6kE3nM8S4SWJjL3DtDvNuzgyUHqns+Bo7mnISW7DsisG
2gOccaYCaAG7TNP3a6ZKKw6qGkv+AiVnsD4ONkn0uT53nOUJD7Lr3cQKTGjn
M62J2Yhxl8TTGZ0k8zNtxIxco1XfF8fut7swQJizMxXEy3S34q/hGzxjUZrZ
LzFQGVKLtOfdkJVlQoIuseU1R0QK2Kir4ICr80ga85y4vIgOk+6TwvAtu7pK
XNkZzzYqJ0tPpZhVqk9VzfiG/Xzg4rkzL2su2rhQIhMI29HQVb3ji2fOdJ7R
CJiXkkYePiSxlqKqMdZDJ/t0ZeZfBvWZCuSMyGtah0deAxV39zAUa0KrfiOx
Easy5OSVErzLRPy0nVRCyAKkWd2/Qr4ymJZeh01n3H3zdKCjzyS0NCg/tZD1
jZDNNPc7u7LlX1KesukMG0dpWpYfcfjZPGRF2gKXLg81pwrAeqG11zWQUCVp
8gB2coj7qf/Dq6xGd3Wfb0xA5OXhDnuvDtY7ca2qL0e/epmEZtwOkFNmmAIO
P34RWpuF5lXlxHDkTJRewli3zuNs+n+XERSsDwhJWX0INGbTtnQo5vfMlUqR
IdzMTrVNFr+Dor+7Bf8Ukp+iVOPam6GzwDyNIli+x1wPXTCcA3GPwIkO2X+C
0Vd48Zx3HtcfBamgcsgIyYrgG9TeR9IVUrasZTVNG+Ytz4dq2CT83XVpRHPe
PhVVt8AronEGUwHEPE4MHSBefYvz6xopFWwufRlnl1Fbm1OeYIeGZVsKr/Oa
rMBTnNM8vIAmBD32p0Gv+BGHlVJLrPDIiKN0jP/w2xN7dBG10Mccd70U2RYp
R/271OhxZ02xzklbsV6MqRh9VwtNo/kHc4sYjIan1rxRL8nj4AoBiHOAguO+
HeM/yXs+etErxAT3pLu++kPhwRbRNSQF9o2JQ6+qb9Y2oE5OsiCxasQP3cIr
WmDXl3ZP10iK4G3BVt9E6xKM1mxdqYresRHrO9D+0NANhPXd6tO4vJSEk/yg
PPrHUbqLb1ZmsQ3JATVk7x/iF1yeeUvR+BLJecC0oF30mMvIEg9Yeyhj1uvS
A+5jNxSS4154i7F+yn48r0tMELjuYDp+2PNoU4rctJT+aRtDfca+dQpKZZ2h
yL4ddq2gOrqHiM8ktPu00aLkhsbA/if0lAXFPAywQM4ixmSzy8Gi8CiCRSWK
asoo9J4TreBx3P8E7gyGjz41RylqcjbPJ1wqLw+PGTgyd2TK5w/MIX/TnpHV
P+hdPxRJptEDYf9O120T0DJXXzbsBInOV5PSNHcNDUsROq6fquSow+/+5djh
4fm0Nq4k4PBrqwO/cnlgwowOVSCW51OHsSG/qn47WRFL0J7BVrFBwbESodIA
0IgY/N9ZSNTJmAifQJxv9HSXliquh5p/ItEz4HYfuEmp/WHN/oZpse/yRPDE
WnHeyY6zUPsxf2Xm7sLYWB8CxhTpOdookptq+lbO8t2beAMXU2Qnk5OUnYwv
nSfMc1OOlZdfwH5jPc8aB2ckZJYzoPDgAanVeNSO5nYTLdnL/f0gD3POf3bK
YD2cFebEUb1Ws2UJezibEDcj2c9rB/e/LKdxI9co0Pn5yFxSXEQeLH9cjDYR
wT8Ffs/N+c241EuUQ5ROZjAAW3wkOC0Y7i3rrvFPbEW70Tloh2z7Xrj4yGLX
8rQLx5HM5K5vDC90bq7mOpVJlL+UqUkUEt+p2gukztmFGno3l+7BxrnaTZTj
w0gWv45FQjzDusEbd4Gcff9DFeYsm/4IalwMMC1ZtaGtsi7lVabOpwWZG0uV
QmnRD1+hRvI0pxfE9AOS6WKfIo9hB3T0bqYZGTMw6dIjwMBOw07n1P1R9dNQ
L6zIVZnjiZY572K4RVb532zzz8Eqcil3EqQt6CAlwBYyi3N1Weeu4bCbB/tV
5AbTjvIhzaVWmoXtJ2wMalBvBbZhELVsbu77ZTFo/O7nwGQF0PNVVFoH6Fl4
Qr9y6k4V51IVd0KF23muQhwAEIM3pEEvI533Tcs1GrQNagqi/QEytun5WHlq
yFKL+Vajvw/vbX6oeZVQ91XDQLkJPrKVlVn1uSXMSeyXYe4P0T7R6S2Gk+Cu
OR67RRbkD9lDA5jzhO+HrzC9vSfybRQRHiJv0RmqQBxSdDE0PqguhIEqA2gX
LIdjgc4VDHfe6YtsJ0NuaIlcm3nJeWQ55Sja5kSEdCOG7I4hpokqhbdK4694
5ZyNE2kMn3LCEd1hGJbVPlopiNgPP+vL9q7W+Hq9fQJql4eUN5IfgGLXIWiQ
BlEWcCcYRgEMjJ2VftPUwsJyntWKQ0H/4BYJ/8k/2cLo/5oPdMzn0gF0llEe
qMcQQ7vC9IWbIWfl+tQ20yMqLAXsxtneljej3fEbEXvbzJmQbwt16Fa854wI
l5Xf0aBWi8u67J5t8LVzhdoMGejZNXPo5Aki+Mq+ODf7KdOnR5Hd7mxsMe6F
U7BjqvI9pEb1NjpJ65dbpCpH6Uj7YjfeFar9BrAsTIq52i82bT9m7F+NVmd5
0jPeE5NgDigrWi30YhhoiTkJBTTc+Pf3eq3l7nEthGj98qUFdm8Uru0yHNOE
/3Ml3htNBNpCJr4HGeJd8YprNGADPdSdfJ33bA6vBVvZcYhb0JxH4M72ViVY
mOemqJbEfSY50YUEe0j4TIldFROM73e5xqmQ5MiyQb77SwTxK9+ZQenwxLMW
n0qQMx/dduHF+ZWiKYWBJLAvIzb/6NidDsWKN9sd1wZbaYr6Mqu9bWX8xUlo
AIqnfJljK8KzNEM/LnsKEGxFBXrpeziAmLiU+aG6LHCNCV2UBMI6VXYlKHim
eD+DpbYxVdIdOx6U8uJ/KBAMqZT5ZQ1G/9dJoADTw0lnNflXgLsB8twJTMat
GjCEu4s0CpB8C0IXwYul7pcE2nc41ig5naHGbcDaSSZ9fzM29ix9TkAFli9S
viexErp+TKELn7XU27UrxnbjKN9BlB9xP8mLmkToJZmckHxhLc6Eou8hmXBC
kSKgCxgrp6txIoLXWjJFzKo8lH6skUsditNWzCQQujuUJPGMRYB7MKFhgYjN
VCsnYesZt5+sJNmWlvCJdkWzHIu8LuMnI/XNyUWEux5l+MYe38cBerLF9Tb3
pESY9Mw/5zAz0YBTaVbIeK+9kVtH9jRpZ3uE+Jv3OQy0m5fHqXQm9p9W18fh
FW5XptYGKbMDHY2f1+fVVL6io0l4w3ggLxqJ5UzV4B1NFcs95kq8SHEgxA2G
a7o7DHc+7PSYEky48iuaTExv4tSpY0PdIrkx0YE6aXs+pw1G0JurmS8V8v0e
hawLa/EhPYJqvJe4og0/yrd2EIpNVXtjpRedpz2EaHaAeoJC0DRy7t5r4NEG
JknyhdhsPgWK4bySmaCW1ipTokFjqOf9FM8nlDp0NpygD2mh6YaTGBSwwqw7
/nS7vHuFjIZsnjNosZfT9Cb8b5PCRM/j+VAYu3+XdIepAjOUlXfsYDqShJSs
7bvoR6yXbBWv0bA17F4ZfmvzabbWigno0IBfeO/icI15wSnjCVkchdp+n/Ib
ftxmhMtD4KoPagul6X76ErHIPsPTMCyYIRejQFgLp18T2Vau9N/nyL/AgAY8
OrfTgBC/lJ/+c3MZX30ENHhDijId8TQOMKN1ybUAmjShZevYxcytRo9MDwaW
WZAYY58hPXhKknvaUMQ3JSbX/99pP/VdtCtZjRIbaAGY0DQYiOAeIWv370CP
+kn3ZQhrPKRJButvldtDT1i5ix/B7rdCOVL8wnkemhH7tuUwBkEfDV7ivv3p
/iNNs9y/6y4pLGLFks41Ul+JHsZ4rensg6F8tsTzN1kOeVL2JgM++ACDlwoH
oW+Mv19sjiHy9jHOCsS77MZfHDEkhPuNocxzcmeWNNuy//WwzhvdXiET1kJU
eCLRnePaKHuyYnK8X9TPf7R6uP8D4s1JJy1fQwPUiA/BH4AGj+2i2Uk1u1dh
rTvFn2QI5OCQZJm8fLTwc2sfNIOLcFFAF0wFR4V1+GgGFtGWwenSpK5TmJIs
iX3rgYEJ8ydoYWu9UoCA7Il6HsE9cv5nDPjDjZCiE4MqiFCq4Abcxu5EZaBx
dTA9CmCERXPfOL0uQh29EzNa66b5Ey6LOJuhfEVCzOpqWWHJz+Vh08nuW3h1
MbnBc2mYqgsMtQCv82R9cf1xoXwp//UAx65ULTFr8xU8BU1Geyqrf9/Q+l3h
vdwCVkEFfiLG1ydOM7xZftdT8uSRi++Y5pfvvbjFBAXAwjCDoN9jQyudUR3l
q0IxMbQIYNtxRqibGKPVkTu5eUpRkU7A5lvTFCH4yDBC77svOVTE9+NnLytn
t29botCjmAcH5s18uVJpD3YZLBvJwz2v4sVWl+w6sWO5rqb4mKzUNq2iGjtI
HVkx6OcKff3SbyWB5Zy8jfOxqANUjFdGzRIqMuK3mTyMATsEbN0+heTvLVrs
nsUBMLhzXvXV6SQPeNZqLFFobxqAYCO9kCcQjF2UgFNz0M0bYn1OdXYvWjj5
SBhZhne9YUpBckmLL20Aye7pTaxN161ILDQQFDfFXzWJ7KWEpIxIKHOSy7Tq
Vvw18w/HVoU00esfEjZzDwzhFsQpnoq/mZRj4sE7HjCsPeWOR8AucPjHmtMf
0ivYbGOTdyHTDI3s/xSAkpgiwcBYPmUy2JxAD/BoEJ3DjcTeyhJeRyeTusv2
x7tw0Sd0CEddftzGDaZvkuuSrL24kWz3ZUhaI7H3Ro9DgTzawJihweFFQrb6
5Q7JmkplKKUeN+vjNiL6Mn3wFARmTDOkXKqMbR3aanS1LZwxD+Ih9vL78uOc
/40FSWMdLzoAe4Beq+9MUsi5HlB5I6T6YPYK+dlcem4OHXWMY5u5XzuTuzS7
yp+HtPGSbGckzXmeuVESV/RxzDdpeofOBmJUsUHGkZllnH1OYJg/slJHuVI5
Aa3Kiak+GVdFJiuu3zqFM6aw+ZLh5XHvko88lxB+EUO5e/22TgW5qLJiqcya
iueNFhKJvV/osODQ/NLllOrp5nM/H61WHP/GsYw9D2kxnm1Q69ipAnT5nk4k
brQcj7FOY95TBKy3MnV4qSrY2BRDyP3ph+pb0RVYJhO4j4oPvGfZVy05ioRN
t1UWH18EeA46n0tlkXgmhtNj8YbVorgaHhYbd+5vnXLctpzTqfZpvrIrEJqd
1i7OzLi/VeixLP/rsgu5yKaheEjZnvH+WocFzU7r1WndrFMgBq5KtymllE/b
KI/c2BO29Xw12hz2IIuzuLc3Xv+WJF3FijE7ivUOVkEKC5aOFFgqkYyRr1r1
v8kbeH0oXIni/a8SxqbmdOkWgtssLGcvO/hYikVL6C4jtLvt44D+NRJooxKm
Ab/nIZHZdDERlr42MgoZhm5ZTCsF+1XWcq0ZBvkdKVqUd7jmvAhwvfvP6sjC
pl+DsMyFgVNAK32mmr3fjvLb+47tg/ooewwBB8fvd3uW3CdSPWoej8/9l7hP
sr3RjdvtJIudHyqZ4RoEYtk+8nG+C4iJ5LfDco/74gX8uOSScePKcDngPHYK
xOT6s+NTH/een4zXFFlrT0PAGq+5ZWXVMTeAApuGKx+nbmUNcVRPqknTkOSN
pVPqUOmdurJ2n9qp53RLOkonp3Hl4DB4pIv/boRscYOxh+OcjIKhuXe0N7kU
1mBGdVFzj1vdp8Ms+Z10gdPAjkL12/F2MirQqJzYJ179gn0oQbXGQDF8HfkQ
EiGghcJCLjw2FeChwo7me0m9lWS2AY1Xx1yFA4xouwyRg/21tSH0coY9ulTO
paLmQWcwd2EfmD1bFS4Wx0OuRNQ64sVy35Mae20SqpYWgAeYRMwhZNJGK4pk
D+ov67fIDoPfFomZevUsfS62Yg9zDcvDSif+XM0sxxXLjzP+CuuZ8oTEOQeL
FEi9B8b04DVU9gqL6XTqg2Xyz6IsOvLlQ5vrVXIRw+d8qrmprfsD7Vz/kx1+
r6vims/r0QXTTNF/XHru5n7H/YZSbhuEMPvACLkTgjICppFg+fbE1AXRwaBH
7dERhZoG/K41sKuWxzgTBUFA9+2Ww/1vm1OZoXKUKLDLXwHKxSWN45LC+yrp
52vEc7fIX+AWSKTkKpsieP5zbuTsRuAozQsCxYZZeRgjhHe6WKfwz0p3UZcT
rr7li2oMYy6o0kymGsrAAIZau/q9j/XgS3u5p17Zcu5Qugi2L8JYKQYHs/xi
Njj/pLQYcW9BZVpwN0JwrFRXwP++04q6bAdFgbDe3WE3FuIbECWRp/qEhAMh
HePAEgwRoS9kmbOzoO71h1SdyRARVT+W7Nzrd/XnCeGCN77HURpAEFE6dN+l
4LgOZzocvXwGAgMW7PpIErb/dNUqVrOEJRLOj/otlIMZ/yBodi/rQud2mmRf
LmBJa0w+P1osiBL/bnks4rXmc2eTR82UZodmj8jcrDxkyxpAP+EHpBgAnIv8
qI+4aHABds1OAQtvCVoiX5lA4rIIwODvs4/bQAsgU39cPNSYFijlaOVMw1a+
a199fN8yZqtGkslaAGR57Sb8crMvxZPKzKslQSeAL2B5Ug29yVstLoiU9g6C
91Un0yl7A15TF2qPJEC3rrB32NwxphA6BOEHKASxy8ZAu1f63tIuXQ4iJUks
Fb2qvYLYFZVYqC7jsw2DZ20/okaAZgxYpiCNnEMjYfKF037WFXVswGYpJqSw
fyCYMRosohBDI4jxFCij0NDz1ow/K4JL1IWZPX7oHogs+QADzsNJXYucdmTs
iuIEvgLe3msmDlq+CtAjq+Xr0XISy1i9F8sXR9JZgdbwR5vqaBFTUu2mMr59
kt2SfaH5RPclxPxMs36l7TDXYKMATJNvGvPB+DZu5lGCMfgqb84sk81Xs8DY
ZpZ39x8cMhPLyRUBOu+5eJQsJ6q/yHGr0puIgDydvgGzrTMMe/LWFc2GgDSQ
Bu4TL1tnmiQNLyoQuxmDeUDzZGztLbAMaDnYRKMAjFYi0E6rAhMNGcoHmf4z
/9axws/X5CuiznPKeHZxNTTcf/eV2nLqplrozsyG5pujFOONGGAxJXR/Xqk/
n8MTgXbjY+oNUWFMs2YCsRn0WLvJFOrueMneWa/QFu76X9S2xH53S2Fqzdhf
t7lF+xl8MKuN+IPGfc6AQJ0L3uXe33Cd+wPgqC+e4xDqwXZY+uvOAAhvtfjJ
zQUXoPl8iK4Tt/wikZWoVLfcLRI8lxvssjMWrCgHnxsBgyzXEy1zPNeAGxMu
8wf6eHjQLngFxoRRF8vdVBWk9fpSR48oZiNVF6Kcqw8CnnnIGsSBEJ+lGYeA
lXSqciUdDvQhYhFHwCzZT6pGGk46xgAlBIrg+43+E0fFIGyE7mGvnZOSkrXX
BCVsYq8h2ExGqm2y1VMou68iMKfeTj0X3ikpvlQ7go5SATKRCHIFP05FUJGn
fj6C1ypjaSmxH1brJsxHID2SBVM+e/39F6bAfpe76ROss5B4ZVd11FrCGFPY
fVEkU40R351AtkMwcVH1P8KqI2eJIvCoWgbv25+4wnaFG8HMnUmTQ5a1N4r4
if4U9DfRJvO0AQ4OrnI42upY7VOMRHsqQBQNZ5GwrlWOxGv7/en/68vLFxbY
sb2cOwQfTDkYUJH122yN9aOPDaUvApLAy/Kw6FkE9qrmNI9KG/dPUfSXoA/l
cgqIJLRIYtDb6e1cXtyFMToEvdF83XQ2sNCDfroFsI1YGz9Hcc/nCCBBMkLn
uc3XrMzg/wshcboezCTns6c1MfuE+6mHPpjj+YkX+YKnI/aI5uFTZpcDals7
enCX98+mw70oFe+Z9brdUTZ/FeorRP8zvFC1xN82GGVG4WR3VA0TZAp90kWT
elVZN2jn2wiT3WT3/UOp758A4nLqyVrHHWT6asbZaPXFOKLjX57twDvd7AiQ
6Rxl0/6grC3TdBC/JpUd1S3jvSJOvaaOZYn0/dFrEIVqZ9DZtqAOpOBSn1Ip
6utO97ZNHa4ugROyTlVcqb/IMBBkq0jSAR2D/DykRvenBG4NH0ttascyXug4
+sIdoGtArY1BOitCFk5nWiB+/Z8TFiekn9enzWgdSCvebrP5WRNv85ayVipa
lJalDk5A9mMSJRNdetcO92mmghbFP5WUC9Pyv8ngGyX6iOZbj8bwFU8hEea1
39lwMhckUh4HpM1NajFtptmYNZn06Ydv2WA7kurmKiYEKhWmDzo2cVGV/AQU
4lhQo57Cbvpu7TaD+pHt8O6eA9AYrleDmqgN7K3dwFpz56bnnUWYCcBcUuqA
vbuEODguMWKiHuLnea4h/3eIsv2BIjdqIXbiJd3cyKoGZGGZ0t4Rk/seQ9Bg
BXpoh3k6frZbBRqcc8CKf6w9IRJ7+z/qD3O5M1sPm56S6oevkujHWl2kWHde
1W0uvy/HSr2Mg6EgDnFxXDGMwxIyJzFS/j3gjWDoObPlAy50uQPZjG1WG1Ao
t9zuVN91rKzCwZylKawCemooCjbRfIiWxKplTbpKXOeH86O2mb8ylNbKPghb
V0wBjFozX7bCwx1TzLXSHLKY6EFEeZabKcapauqAMJEPxN76kNJHQMrznDYV
BIhXV/j5dbvOI14lJhlY3CjY1gSgtpBj8Rm9P4+WB+8sSvF9TRqfj5aXYxnL
odvBaMvTXcbI8buhwhSlWX3/7OGMvITSqA2FFGT0iodCiipdZnQ/58qa4Mtw
TiwkwxRfeJAwnImVClVTfP+W1nUSUDlf+DixQgkFL0tqSHUBw6lE5EkW5vgg
dx8m2gk1DhwPC6fcECQNk3sFSACrj0VVNWSp0yYNSWOzVhQPCL3A/Z5JTJrH
DG0RB9L0ycM7wGqHU5dwrSjsXPmx6t51eDomAdYHVjZqKU7v+MGk3qkn8rp9
HraHj9PUWllXZ/cHcbO5hJED0DeD60iaDHiedyzT+e6ZERLR7Eqst6AmdN87
BsBOlP/5ss3/X9Fq9MWuTt3Qm+gmHPSu3VoYyRj6TqeEMcC6mPvrtV2Gg5gc
ghqTl/IfB0ANG7uFxALI3fbXq4Fw7S0PVb8VPI71rMrE/IUIOiSH8woJL/CM
RYb6eJleJHKoCMfawOI3oWQ8yD/ULcabe6RUwx20zuoUtH/YAm5fCPMBjL78
5aGKcEldz3wD+c0UWkNjm4Fg5hxviQKyKOvLTEZ6s1ONm6CylFweEjxXdOEN
6/E8H6C0r+347PUiDvMfL+jUcFN/9YBy2MCYfCB970VG8aHv/J+43m33pvAY
oZ1ESJia4WdZcy/lXAAGRHTZT9htQ2HiXwSCfe/i6yIUVA2iijyLSCP6MReT
zEMvKvK45rPr5mizCxNDQ/QXqzMA5C8bgCE2Pidw+qjpbQRfJJ31oownI5Ok
A0WbNq0xm8nPSHr/kAjADcghPbCDRTtldyaDVL6/jcGIcoeKtGJg8SwgB0TJ
DDEFcuNML9Tk9Pu1Tj9OE6Bei6dLWJakNTyeDB68ZS5rXIZCt0cDvaem2zat
UpM8spOIyViQdGMfEObgrfl3DQkMbqRnUeP3myWMfqnsC6jLxVbcKpD4dpDA
WS6+QY4H2nK7mOG7tnAzoGeK3xAikV9Z4egrIvi17uCnJXGcE9kuQKjVlGvp
8DkSQJGY9dwZriRilNQZtUErTS087ujPJS8bi8xiSEW+j9ucjXH4qZO+VRCT
soQDBwX4iZ2BVrPInGtjafMiLxeUQs9N+yuM8e48uN0sA9Tz1xviRpxS2/Hn
JBwWw4++pluNdsCNEO8R82g+0jnuCpCCsq1n2JAVdPzQM0vMAGYXY3nX0iSO
OvIVK+YJKu7xlNgJ/DU+M20FAjKAku4k8JzZKsCH57/JvnHGjjHuKYG4bg8I
/fX5dw5NU2IvqOGrhmny4ulFyNEnPge3mJQz+4ep55U3+HVw3kgmZ+5MJ/j4
NT1nPp3KWJaCx47Hr+z9dZcBijDy1kNl1vaqEX/ZA11lYmwOdmLRzfy5Zz82
J2MHYQSf8KRriqlGwTBcNoCGNWG21O3M3QvBayrLtuTE1DYnvfvYgkxAMCQS
sStGBmYYoT161jSCgf4jkkVeQ72VBtXZP1NWP7WnHHR2HcKcRuKXXEuaV0vy
v+fsZvlJDBxhBc6V67MegHe6EkRCzzWAv01brIdwTzK6mFV4hWuldGDiWa1u
ru1sd9+KPY4SdQMImWxH0PR+at4egR/oqFdbJIPEjhKD6u+5abeqjAsrkpnU
jE8JWMiAmlO6ixzILLrG75A55vnH1UYQcvuPfaMsADuOa2f2+PO03sDLN48T
yXLDvJ3hiOhSszDQnCOU+YcMsESVTaQrrVx07Eqb0s0g5Pvj7+72ki/DMti1
vW7ukS6IoNoJdfR5Kerdey9SdsODAS5Wrsr+J2I7auFcEor/JJCFxDQdvuV/
Ja3O4EG24A/T6+RjA0qJImcKfGGo66lKVEiO9tcIchKsGkFwNucewpAbFYxM
1Yg7UUZufrHTVWd0EnzMWYqSg6UIc29pbTLdDAfSsz9l6GU13QrQyUUWShmj
DVPa1H4yyi4oRvPKBP4OreEEVumhWjdi3AKdN+Z2RmeOZHloEAEJrN7MKluO
yVtZPrGyLECiZPjpIVn+9Xa/KSUpJKdA09+b/PXwRP/wVZ158XJJSB3ZtCRX
E5IZwX0yTN7DxuOO1QHB7mqmlbVF1hSd6uTI+LrHHttuyP8JAvesESt/OHpV
3ZWGv0euQCpZlo9T01SBITGZAEzD36od2vl8R+BvgI6kd12fYK091rC1JLb0
wPQB/lf0JUVQ8nnXgyWd1HkWV7FKzutZDkRLbdhdxgBnhblsK2x463aCa+Wh
Uevf9uUDWeqbX+9mR3/++sLpXAGeMZQ9rEMJEAbH2sjKNOmRAktD9Hz7H3Wn
A7pN4X+OubkeEBA6+VWNgINwJEHqiU4OCjDdEEjZeXu2otGvYVTqrlU0S7MP
/dToGEbmHWnvy0ef6rY8GCTDhqOC48u1p4H254SflJVcy+9WzhrzCXseFmUj
L/o593gWYvCw1BuVAmHmORck+oE8wxkwbli96ndEg+6nYT5ieeINh9quKlnj
aEDMJsTl2qf7Gm4MGcBW4y/oR+pcW51G6OJ15hhkIANuYL58k9LWA0yjOORn
uGapnrRjwRapiw0z1q3XeUhkwo12SbuY1BoK+iepe8SVbka3lwgqGe7lzsFG
16REcDE0FXVjY048BWbbLea+8riK0rRtJ8ov8se2Qt8Pw7p7lsdOMhNceygb
4JxKx96dm4lBx7uW1jYyOmQlJgCVv5d63RIgkihp6Y6HqVimGRRz4vtubz9o
EcTAj+4SlNYKGCyBpEWQkuOBNbrN//A2GL6qTQXR+WdlG2mGOdr0BRsY5u/2
x0i81P5UMu6gPH45av8EeSn7LqjpOmrXtKmkqocRIkbytiHiFYxyfTD3B7I7
thf5pUe2ckw6Y9iHwZ8LlTCQPnbgsBRNx/BfX5uxLQ+30x7rwQ7mtJYjx9F9
yGoxaWeWZ66Ht7012LkYpAH76D5ioJq+J3xx3H6xdOeNd916qm3QwyNa/xAB
OFKBL3vBTn30mn5YKWliuj3XlMeQS0+kXRyhrOCy8iO4ldKPfmmTizLOmy6v
a5Rc9KvjSxbTYqntksc++T/aTRxmR8E/9RxLSFCGCJF0GMKKlBQn81fiM/12
6UKHy55lW1HlaY3/bio+4hiB+gSMgq2JgNtijRkEjSP8pewv39N2TpmfKoyI
uq9GBhpdVX8H/YhJvqDbfpLnb3XfTQrHNyfdqWdMU7uFAmQQsuzsqDx2Ra6u
Tf/M2JT1lQvqvkKvrm8k3xLQck/g5VMdmlqPyFCQHGnCP5DE4CAeI5PSv999
zFgHA+mvSDia0Ucrpj/E7pSw7mpKtqg5ew2yJq8u4+2z+uAH6BhMK03mdmF2
KcfxATKB959VQbHUljuhbqy2Z99Dh6NmQqRL2qvoAVIiuSTM/gYllJ37v73k
9VZkMspNHl1L76J3lasJ4ifBFm4v/tXGxhjk5cgVy/iJ6OAsazZ59Th3XD54
le/j82KB+Yh81f+HbJ7TjweSm2kJKoHpQI+whOWQZAKxSc4MxpqMwZKx/h9u
KS5t69AHt/usvW4C8Q7jntazMXIFVUs8PnvTeP1KXc5ZtG2uoHhzCYhz9QnU
+KQBiXdCIQmCBniA0/4FRYhRGo/kX8e5Ti27LI/iT1EH3IJOIftI42Eg7sG7
CIRAF939BSeos8hX8Y5pEOa73Y37zIdYlvnwSAtnlAZSumIrUso6hX/3Ng09
7s+XJUbCDeqBOjVODpKo6mXSvpz9s+/PjUYq2a0/cVNu0Z/3APkGvuikhaAQ
kwsoueTwnie7+NTEz0qkpuEu8/ll+4oZEMiRnNfIgeP3aDv9XoVqN9xo+L1H
kOV8WraLa5xRlLU0hM1IHkbgnyJ8c+RcKKJDStKut44OQLkTk/DoYdVsM1LL
nhbotUs9n9S6nf98gvhXP4IJ63WMod65rs7+g11s9ouj26XQ6hQQeNQLqMdC
0kZ3HAOqAhF0VSYU8FYfLdyamOgClmm+AD41oq/ElgVeZJKJ2L0WxgNixM0i
LMsaShVKi4bI1CALpwPDS8ADdTDzSsENKNGS51ZSK1FWMzS1u6cfugGtUbwX
H4/03vxA81Gan9/j1UtM/RNJ0kCgL+iyvCUiGRlrJl1WOkZcT+ruo+G0Y8ZE
n7b3G5cOMuXyi8NLAkVf1p3sWNQ4ky6fseYXVD25TXm20uDASf06a422vOr5
6lGeExFPqA6EHOw5Bbx2n+jWoPIE+v+Fju/FfuzhUa7x5GZ1nAdwkHUOOJXT
YBeymfW3WoWsyGidaeivFidxWv4BJw7pX3kFDiAz2WRrIXy0h1+b2jotjyhO
TSL7U/1LhVIsY3VS+jf84xmO6h0TM4CfbGK/tFeGVObtKdx6nqatJM75QPxg
6WKnOLvT23sex20mVUqTHY/Bd1FPPjQJ7pCpfUAdMNqM+wbAOVtxzZ7L6Rtn
ySB+8qkHrufTkMr9fksZSMdxQdEoySBfgB3PzN362xUjenp4rKKjs7ML604g
nv+PL9p6QUn5YLqpjLAlIrnxxlv92ziYZfZCMnycoUFbRcVa0/UM9qYZ5l/b
+a/BCqustonkQ7DRLg7XkntREvSUVKGEPJmj4a7ruRwN/wH96LaMGqYd+m1h
36+hn6KG8gxbXOdR6GUTwXcmtJ4d5x3WhvmgehIhP78hPU02OCfYGegYOVw2
M74xq0TnV7NkXGRRFtlRUlJG7U7C7woJEmQSdXMhNRt5x/sk1bbHB+Bw7bmD
t12+NqN4F0WiJwRD00j14BQUV1YDm8s4VvE1w6o+PwmJ8GsTOhbNVIgtu08O
3N0c4sp5VjcVBy5zJRJ8qatfS5B+xILYgL6UZC7g47EQT4lZLJustVSTDAjm
EDDwn/u2ORaS96NN8r/UBF3e4gs0VTOY4xJxZY3CqUlJD3+X7IHqR6x3cnhd
dmvWd00A2wvWWEVWLFWa11lVatBJcxaGvDBD8r0kyXMeSHy9L7vkEU+dBlxL
C/Cyr6MbTu3FpQfwq8UIe2cVU3Bzk5hYDssn+MiUthSDmD6/qhsu0ZujPL/H
P4YzGslOhHb39Aj1uNrNefqxcSrCqVq0A2+nEvGtSf7I1zI30SxSruMjnZHn
GU/dwOF+iDAqfSrW61PlCKicAvOMA/ZWA6FzQuiemEcWG4OlwTyPEmtXV+VM
Z6pFwhtclDgZYCvtE38ESe1QBVlQpi0xjdVniyw9saDEgWE4NbqpihRjmzNf
cm+2XH4yEXK0YSmdOc2Px7s6+YOE9qRvfwVbxAnmTk8wYAmZyAiSv6xm+t1/
rZN329P0kmrJ020de2MWeqjimgNPnZiF0/7dgteam7Pd+MKbNwFv8d8ZwRCs
tK1tauUjowYKvO0rSkPJR2Pb246RyINyJ6VOtLtqoG6i1exRNIv584ggU3cF
iXVrBRA0OuAiada+JzDn75vc+2klgK1f2cw9E6Z6u0xg2OyqD9+dZlq06Ykx
CJ30Gq4XSln+Dr22nShFM8JZIO0q7Uu3+PwgYn4F6AkcIjSO6SQ0JrrdiHZi
WORpF5F6vlzkcLyrN2WEzSPrm1QB9xA0vd6JQCCEvjf4zRAK2V6W070v/LCU
+UtQ2HuVFwFLIJSHXhSGaUeBpM6Em/ETxxak8byDa8yrGPEQIMpoWeLEJWYv
ejc1EyE5xVby8Pck4t9ik80zAfMyK4+NscQje3zIwEBAaVfIxC4aaGnJ84JY
6gUvEWBI8YWpdoBx7/IhLNwoaSmM+SPJsmBlun4bf1LzBSPWTIy+V9ASCjoY
ZU1eSG5WDfQzAwoe0DZouN+kue+ZgpHtZ9Ih8T1ZMvIBBJymAfa/Sy7o040s
5p10UkQJ+OeW7QoAiVQ8LxnRfgYmjtxNVKl+PdW+J1MVNKcxDfxqx0jWP9Xy
qR6B3vVUVHjszQfq+9Usnq8jZ7v2l/0ntAWaWqIVp8nHSJFdeOsUAsQXIK2X
NSg2gEJjzrDdFISB/wLINcDIga9Rc4keLW+BubGmqOUdS5p5xNlRgTMhAYdh
ospGfCTOi8/zh8U+D71dq/fNRVGYIdUFBvQ5aagN9Jf4cVutmTClEdON9Bko
76avan/aAqFTHHeQTbY4uQ0xss8SPTpEDtUK0XYp1vBo+Trmin33XlnorWLQ
m2xu2QEeh/f6umVAFu+l4N+BPq33BsrAUg/LeRYPzRYD2iuo2WXm/i3sfBNi
XDFqdF2QirNvdT7tyfCWRst7pYR8gL21Bfpu2SEg+OrMhkdCdnlAt8rnV3t2
lWZYzwAElQD6ttlX8upHWcYN+cOB09Nrl2IGDhawzHAAG8R7Xxe0lZ+4WdNT
8gSuj/UdOyiRiwfOJkBTwqTFJLdUiznnhnJSd+0pUuxTEETUoEQyj11xZrf9
xvQaW/lS3gcRJQGiYMWL18tf1S8NX2TaEtoFsaS8CYQRmZ5uGK0eJXi7MERW
wG1CGEmmMWmiP/Gzu1GK1B468RBzUafOHvlTsdEu1WEdQGAzoAdDR8jtS1JV
spOsDO0TvwBn15DulJZNT1Z1ofEOtLI7sYrqgHpeMuA9XkZ32CFMU2Tsv7dA
QczWuLoeD/75du6e9Q7VVYIcUcdUywijYS56HIgtUgYJsGq6O5oybKZC2huR
ofrJpNG0UWmksPhkn/8nAzG0Aa1ctT3scUARCvSXwJrc1s0yFeMO41Yi1mPA
odhzHemZF4hEiSuue6swKQP4glfVUJWCWDornnAM0mfvSJxVb2uEz6YRgmyU
L9GFKfOKiOxoI7V18Ji6RnW9eLGU9qGKAITjcugZTxhoPrrMPAE9xItZedtr
RY4WebkwSFLPsOez/QxRebkrqd7zNqSZ3wEQQijoG/fJE7E74SUEOF2VFg7t
7Gq1cERE41/UAoeOVPsjilPlu6FQ0jQzZuEccSyPjgw5mCMmnQkJymWaMHrD
6sEx4xvj+96KLhNqyfxzs7bPDwcZflcg5Hie9kZtdAaF4YZOYSvVN/EfDx+Z
GBzQnrh8SVtA0NggJt+A0+oA+HzJ+mpf/qYJqGNX933BYE4eBZpmw90XQbXN
A17GyQWaFZTGwxxktz09+AFR1SgxGYFQTMpA6LNZBgWZHEIaPAP0k5Mmxqv8
MO9Q6mim4dorpACQsC/g8pX/d7OQNE+oaIA0EkO1nkT6pqLXCRNUN+Sb9wOY
zkZ86hrvrsJUBbwTnKr+dT/giPx63W94CL0FFg8Nqnddtn+/7MqhlxlswBCW
JT1d5eJbeBw7QnzYeTnIiTlf3FwSoBB+K8Kt71QJyko1YAXhNIN/JLxIt5pa
cckK5vdVkdiE07oCp/RXj+jpsP7UKyCJgvZcda4DTApniqB/h/9T7meZ1AkM
vlnSQd59z/155NCgczlmNIk6SIjz1SU7yQ94OhbhgmlSmuTFKdYKRFC0cuaG
OzL17K5JXYbv+toU9W0MHRxwcwxvhSbwHZVSHa+OuSoc4m1oOVFjFnvSk+aI
luU5Abmaqqt4Ib0VWxNjPZYKNOklrPhDHduI/UzTH3B97WpL+d+a0WLjodB9
oSVBWtBQJOMVT9rRs8SSuxpVOfO1HrvC/vLd82PJrxEN6uXpA2RGU/sOCO/N
JY8HdAwnxcf5IKaLfEUznro97W2ixVXPIV01xOxnlojb3D/DJ2hDAJc/jlxW
B8+JWI5TKzFiswcM8jmDmLJBLlvcWmRBhTm4x25MGiVDRFCICqjbvq4IFjPk
dXbMaoGdjZSVqgppo0yUF8nYVsrUJ7dd50y+UuVpUMJfzsXphey21kKqZJuV
00Q1DvLB7swESdrqtEsJeZY5nIQ4pm8ru6vzEgmDA/gHnYVA02I0QUwcIj9A
xwrTnAzYPhpa4wXcoTtENLDW/jdYCPC77nQAhKJacISkn+xF8N9+4uE/5AAS
Gt+Ad5dxouKjlKuhQLEoSf+0mjz+pTDFCr6a2Uxi9oObVt3ZVuGNyQQ3xUJv
8pVseFyZDny82CEqh1mC3t9k7Zc7yt8FpYNuqO791ZTNTiSEi8IXzSpOkkYY
OiS+NcZgYG2PstYYWL/aimOnAPfLIdLyLki/V0mG3oRYDjSqSgC3o4k8lSTP
jinSfiMxOEL4BOeKBTXn5ne+rUupZsUpfmq9JT7d3UWxj9l6y8CfTFk0SY/m
bJ/jzscs4pKobIQIDubEZlxsrI1aRQJKUQ4spOSt0sKQj6c777E/OMTUOvk9
K+sZA0eroCpHGqV4V8TfEU69NskaY0/cEdytQUcb9dor2NN9YHSZofvwV/gw
arVXVlmoNN1BSjwYgWhh7HZp6wDZIWVB7cpzybFfPmLd/Jsfi9NGzL9H0NO9
fblenOepLwsDi3qKZTg3NZ7dlM7uVBo1XyEqn3pAcsshiG9vtJwZy4HDzfqW
ukzcByUNoCQrfRBh6ccPDuV1tIzOp+FmVsnbxfzKo1gMmUKTNGb64nnmN8YQ
84VnRfdNZIoAbOTrQYYSe5Kj7hxyHwhCsgX8EGaad8m7FSMSCchNKYarJ7DR
nXp7tTagokZDROrA0V0mrkeuJ/3nBjBo0ahoiQ0lMGIpg2sEaTgHnvUiVk23
kb9808vBvgx4Sl3FdVTOCLNez0sDjb0HPngXZv/bFMohUvB5GCBKN0crYmF1
MV9RdJFyukSm6oSoD22nOo1FlqF0gLFQjaijd27E9jA3onHWgdJceh4D225n
GzIJuKFVJeh8nie2bRPBB9lXTyea/ykmZNpDUBN7yjD3nLbnIwUm8umj8ZQ6
B5Lm9n06cCxmObnLWngoe9c51iIUdEL1hNRd1PgLcU3bgl30O2fG3MouWcxT
vhzks8dqrCLX74eau8MdhijZ9BphS53LhJS523MGgLq9RbtSvreHCtJGi/vj
IlxBpJmzHZdVAhutLBzuMPDE1o7AwQGo5vCaBvMQKmEpRe1qE9VvQkWDvyUH
FNuDJncixfFC7DYJfi+lvcCfYDQoTMM3/0tHj2HeVjWEdzh3sWDxF788NLIR
8qAWOFYg59Tg+3d/KY9M0BoeUSDTIyBGEAKIW3NV6h9TM/8J9ZyhK5rF3xP4
MxoqCW6Fqkwy7Db9G3Zz/EFzwesyGZ+2bnyqJdylPw1mQyNDW33t87wWBvLZ
7JK58vVzgWWDlsJ1MPyYjEru2ra41vfCGO3YUsnMg1P7ZmxvDa3cgmqyHjFF
SKoh/VAA7YYB8wY5BQYsZ2rbfAxYWkpFKdOm5QmZebQTquFgJ8TpbcenS1ny
KnfjF3hinjNUuy88G/6iGqZHiDUI3LVlqFphgZ5VMRMPgt76dBBo2fuGiQQF
GLhfK+4WQarJ1Ip5Q8f9e+vmiUelXPthUmEndV2QxMi7SccSnLh4syHXVDaD
fA3CoWjDYHL3kAjExR9b79D7m7ClEfyKab3NV0ozuSaC0232tFQqk5ZUUgU/
uKyHqCM1hjlhLzpjyo9SQ6Cnsl1XZgM/VYeIcVbWTL1HH0CdHIFXM4FtaW8J
YRbpYfJylmra5pkxrZVmnNGlLrw9fFo6d2sM3brBiudfntu7EaFOWchuCOab
gDckBqW7By8Vy88inYOngibLsM5Thll6HFZ7kqMlkPivDucFsBVH6XRtRqeG
7e6dJkKsPt6AjS8CL10bEJCV7X/cSdFimbiRi6xlIt4nl+PIvXXg97C4L1ki
48SG+hufk4vqLS/geuuXzK9QKJgs66GiqskNw2o5C/MkjtkRV6NQJCcDetNl
uhYAvwZzTpMQNIk8xhWqTdKCjt/RdCzW4zayRENPmX/qNe2qzJ0i5IHDrl1I
0b3yhelqwFrV9IgCRv19mQS4IGH7KyvxopnJQhCvg3RDaptg3hZyHzwGKq8w
Yq3KRVpJY9cKG1+stBQnFQJcOvoDJpe0bXY7kY5lJJzwcXO1IC09Vk31BqBU
z8S/OJ0dYhIzaoTMbJDTYd7eMN0cNlhOX1pkYuVAWwF7neIqi+AMBOpge7en
4zOQbePvHYUoEVSCj9ri3L6pz5dkYuiVYyoCIuw3a1KnIBLB5kvgaWk28tkY
eACJLlvPRGiOrQl/PFRlycaDmhBmHRGAUy0O1l6nSfXjqqMwAleeh11Hg7y1
j0QzFgS2+SdfbQaqgBzdO9MNRjktVXmrUMoJ1Ns6ganfwxK9HeorzJi/ugfi
bWlNbr12h9isBTCZK+3e34/9Jkt2wuRMRlRqj0qNLIdunjiqf+u3G30nKfjm
Ma/0PhyRcnXsr8cRGIrXkE+ukLzWzzpWt+exi1ohYdLKRc7d6tzI0sphDEhO
A390FeTqm+IbRYCGzn6iJ7LD/6aOsljyEt1zmEWAuFDoklFRxVsBfeipb2cd
sycYHcdaxCywCSTPnIESZ2yT1pr/GegHpTipZZhlUM0Hkd5rD0XZf+SIC8NU
yLbmxOWWLqL9HJLiDp7Ms9mYaHIaf8h57pCZfHPS3SK4e/owzA/lTOnwm8xy
7W29AFSBZBLzjG0xVcbQiLXs6A1yRMuvZQjS27Qex/l61uZMifsIxabHHDWO
mODjB/Vua0lH4qPIJCDBhq8nK92eBRIIseryAYosoQ5awTZZNmkp8ncF+LkA
2f/PP+K22bdDOZOYwaiHXd+LUyWPZMWVDUfB++X4Y/Iepjv0uaJXGGud5j6d
ehFuAHG98LTb5r4J9SJVl5sESQFhpBgR0HIv43SbOHd3RTkQ0RHjX+5Sii57
FSnBkL8AhluDzYBTPfxc0RXlUTFpbjwenDjyNq+Dm//5OaJuKpT6aaCepHLS
6gMDCPmFDz7PLkrY/zExti+yPf33mPdI6wjQylgE0NHEDnFwFgMStREzvjJ6
NBmZvPjZYPIBwytf0dl7i3t2wOW2EaXPPqq7SXiOgX8C0f6Yx95EN5oz7QLf
zN4EHGbffvnFLP8w83+07iDo0FXm9cyldh0u7YgCD1qLef67EWiExanPwmB6
exT0HCuY2b5hxEjrX0J20ZkjfXXDnQ8uteIkH9EsKDvggRsz6rKCprGrcB+0
bbol6kXF0L0h5qHB++IIU/ounZD412WjpoaOHTw1XgWnIFNI5U1Rx7Bt5XaU
1lBiQCbOn4G4gSnvg9Hzi5L167teDC78fncWQ2QrB3HR4QldXRaihiQap4dC
3l+0hshy5WTx3a5UZgMzoL+rByKdiq3VQRdEG/+L53Pjh1JoCJ3G4aVgyyig
/vhlGB+DD95tLcQMppZVPZNXd2cuqqPCZlH9AmetJFeY68RxFRq6D8mORQLj
0GQiRoR9MjCWaIbRkaGFTwKhSV78vFK6AgLbZDzmBXl7PEYuzxgK22lLBq+E
kjqoImDgQMSxDSKKUTd6UVu9Ny08IrvBQweSK27SWWxA65MIEBp65s3HNFHQ
EexoSwYXlOct5x/LoCj04E0t149M3wrlfBRorS3Tmwe7ZzdaQAVet9VDZZqT
n4YiTMrJpuUuU7gl7CmuFfDQyO+hADJvTWJk8numB6QDckwjjR+5oGrO2dAu
T64l+YyW6n2K2eQuUM2lSlTBjaRTdAgqKK/bEN3mWBV3+wbU8C4BlSMZIBV1
DucYjMR5LwQM9sLKaMyfIRNbXf8xZlhQgFw0m1YeAoXqZ4e2DTNVx13oPjFy
6XUFc+jdR8SAIkylXa1JIcJAvo+yjSl+/5zFaBzSsYBOpeHqnBqjpkmNwFCH
PrkWtGSb8AzhH5lmWAr+OBP4zoVFFZo/KVnMSYI7cKJtFt/+M6m0/02BNnky
oSgdh+qbzlKPDekw4IFXflT+kl9cxxXxdigm2NnzVDlCx/Ic3HQaHhQ8d7tR
jSFDm8HJiGsGRmp0wWQaSEw05J/RVdbLvIpraJP/3ZffER1PZCoKbVdyC5Wy
Z8VCaiFBqW9SwEhwnTHukaMqEYfQ4erB+ZVE5TfC+vXnlqTHMsZklx5YluBO
WfqDNRVzZwx2UWxMs7uqdRNN4Ucprw7+9jJvFgYSgZZDKiBK90wfzogpn1Jr
b91IQZmUTm3yUoHh+Jx3cT8T2CgP+EhlWsvNfIe+Y/aGD7S10mLfsPSUb/el
ckr3OUbKMCEOAgZdboPrmTrZe2urykVAa3fbkNy2jnoeDECN00Ibcn7Qrq3t
cR+LsXGCgH5g989QBICIKSR//DhCvHNoc53Z3igTnF3x6MiKz5buNtlYfByP
EkWWbQnU1xZV+NeB5opu2BAjuU30ZmVctHPG0A3h9CoIe79NU+/JppTlVEzT
+CykHwTTiRD4nQb5MhubrMEvAz/fYOigpZ5LpzUbndkSXgIBKIQVNDAJp3lG
/+AmOrYW780wyPrtd+bxwStOwmOj1vg93jn7hqdcYpjqr7ItfQ8E8Vo1FhB0
vFPe9DObOFbmeUlw6CkIq+RcCprhJSK/UZ+X7bzQbj7xbL2ThOUdBQYLOZiT
iuPqDgsphZKfGbzZ9jPECGLnWTRGVkb7KYgE8QBbG+oSRgI/Ly4MjQgtSvBp
9DwGaDYAfzr8cXhi+q0WuLfEYzOAMuMUnXxhohZR/7fixAUn/aHjhzn1HwVz
LoJ6asqBcB7L8cutgWuG9aEotKxmLbdWgMTtSy+mqDsREjlsf60M57rlVVmx
QyJGDvcpxWcHI816tZ12v1vCNJClQyv50KON57v0OH3aKIBRmmhA5BoPtGag
BJl4DHpYOy9I/jBdjoCLJZGwQ/3MYfzzntwzY/wa3Wpisulrtx08mUhzNPzO
Nk0FfmGULyuZp3PiwCyqZIIYttfqUw7NUWM3ImElIM2BuXodCK17l4QlruM2
Trt9u7F7+OwAyx3Lx8wxJ5FtPjIpFnG4yplbjiOVFtp/6TM/Zy/mqMC/Uvtk
Z5Po5jVk10J8gvPCsP/QXJzVIud2w6rPwYXcYKOplZJYcIPL6/LrFcQCLAbo
WmwxtzUQJv675fra6/5h5sQ4It+a/7F7iQrWtbolUPfFVokfjdyAqV2VOUaJ
lZdR91JZYKi66OAsyEpH9dMzP9AtQVMUthzduBnhAP/evV+xOuo4nlvt02uH
CDzjQQdoKGPrqF+FSUGtdvt8WuGGrkE/xptBg4KgZRzQ+AdjXM/HO7gxMMBw
cZjZvPit57LgkKJYomKpPg/WcwkeKk8oh5zwy9+y7yy14QIK33dfKReg6ZUn
th/f5n9LuLzzvO5WCj4LxNB03iJWOeJq6BQ5hPXGXX63jFgrZ7NejDs9KdtV
EAlRl9mZw65ZkYaDayeMdmG9HjTuvV3XWslzygOPHmfaueG47Iq5aFv39Ikh
3IGPnB/oD36F5JbVJknjwpzhVX4tMeDattiwEaYrmhv1PwecrY9mzpUt3iDP
ScBRWepR44qjT1fEeykUdj6vMQjFzdt9/4xsQ3uPQWtodBiFmyNYlRZJPIHW
gHhgviwCnOihhHSOW5ic4NNeT68MZtYN0zHzydJC6q/WfJgGtTlAjCfui0UB
j4QyFrURQIRDYzyKcVBdY8k7+lHKqEFDHriqZsEzXwK5NqDUeZVigtPP/k++
EJSsQCEl4S/Qbt1fBf5NU1WTKnfBWJNz2BBbsAApMcWUPs8uBjJOh9ArxttV
u0adJ0CTtqVx1H1dDO0RjBQ89nO3tj3wTiGliFzgNITJjtAwFBo04EAg9kiG
FK79MKX3jnJIkWJ4exe4svaX70wxo1Hu9glvGq70y7momyOkjUOBC8yDHK9z
YmBkZ39tza5v1KitSwRsj4XzYXbet9/5H6kLZ+/Nh1clZWk0GGPxiU2D9xsM
3vGrfhs2icgbZZC9KeJpUoCl9UsdZDi3BFBqDXpCEENqy2jIlTDeUd0U7rue
qF/T7NJpwr5SCuPG/A9jmNzDBZN2naBEPicchKn+fwViyPl7oCSeHDe0cpwT
1VNwwazZkbM5GJraUBv15eXyxyJzjqDf45D4/GtMlVvuS5XcA7blTAyk2m1L
Sq88E301wJ4RpLjDcUUOzgVorwNCPBJ43gzJ7SwwBasy2msW+7XxJIUaDT8f
w+bUUwtuMwanWC56kjhyQXPiSgDIYWk39jPgEDfmikXou1MM7UFn4eqr9N6j
NMBuIZ8v+FxYqrd0KHuDkWqjt5o6B72kcAW/+QeFuFPVgMuTlMAroX+O8cIv
JEL28OnDt6S09oI3muB22p6Kcq0RPp8edkorNxyLlfj/qwh6oJdL0ierRNyI
iyzTM9GtXKFLWe+7k+wLiLzc7swmgS/wXbUCXaeiAgVNTNfc0pmUv3EmvmrT
R26gEABB4NmgrPUFQtIzvgwkHL51bSH9BDjYnnFV179K+acBRhpnzXg5Ahts
HKEHC14rqV+lPK7wERxA/fz4U+c+IOHlY5v3xrrOpp7/Bk8U6/c2YjBQorOv
GnbOa9d8mmJ8aEQPNit65SNvQNWC2oiBMga3O4va7LwFZDDv471DuSo58UqN
13TLxX7hLMzcnrkeZ5bh4Rvp8RDzGStkKs/INS6/7kl3FRePSpUthI2PZEWy
nEfjxu/lcFAn+xPvBxEuhOgqkSmbe1s/Jm3kIAYe1FfNPZxxUzu3+DNeOXjr
4rKxV0a6PIBkiaOvAK5LNjg13WbRJGRRvzXDsHVeVj+hqJdNBbh7jfvRrFhA
zQTDVreZJjgQm0tKvWBJMQaeCE75zSbRe0pdXxOeBOXPJ07S7d9jBgInwx0R
uFXZ6Cf5ZxZYV1T16lk+xRdQGrTUKWQxIHm4fyJGCobHXicCAQHEHOizO2L7
3ARgM8k5p9Te/wCpCpxhCXYbXFd265aqdlUF6GvSD5Vt6ZWVF3/fcSvVIYhz
V/O6KSMmWY5mGTx0EQORRH/zpXPPuWKgceH1SQHlb7Wu4pmuut6a3hbUPRED
aKeH2gtX/6f0lkWjJvimhI6AiKahEgYXL9FmV4a5x8v+KWge39nl1yAmCRvG
5SgHg4xHUZz8dua22SAjg2c638Y3dKkcmAvVwn9oEFTf/S0qs8jfZ2nbYXAi
0qBa1705Nc8EPnhQS6+UQHbWtzWnLciS1Ef+V5Rq4wvYBc91t6nJ3XWt2GaD
CKzrHRkU5sZNwMznO1ZD1Ien0VLRKFPy+4keKmzR5fU4pLVwY9hTrnthXgLR
61PudcjO7CdUxDr8EQC1v7b0CKuanEFGd0ynEOZ+u6rYNgkeOuOjdYjRnrXf
/JxIRwcBw3uU7HfSwJuGCpLS5vzG3RF4eewIHRPWYv9UK2ZnTx4I3b/Dzqjt
2Oo374Bqa80probBpdbyQORORZAmIzwvNpulZaNwGBiSSINreN/vbWm1edgH
jht2i8uv/qEj7K5bRr7ZcV3EVKzx3JAIiMdtZb8Akd9J1AvVY3FtdkBR9iQh
eg0jRLydHD2IuDswfCWDFR614nj9pKBCiRAJOb04J313yzi9hKeh/M+PQ8FG
ZOHPT7TQNPIZRKTGX2ukJxyfAUJR9mVT5qH6BSV1p/PwhPy2824Fe7anCY5Z
iBrJq05DiL4qDOJJfyRvUfpZkPEePvmoEwNhYoxI6oa4FjAq+m/AHnkhFumF
EbV7VbnwUbNaJ8IFcIP8uZqoN9Tpe7NImDNEgSovHWBeAw0tSwq/NOWcVwvI
cGANuqI/N4yoWDIsxzRFFy5LzkQxJw6JkEuCJYNmqepsRvCvFjnnCYrogNAB
c1Vabq0nnvKxq9WlynQ8qgvAouq8WAI47LzFXIf7EYUt+YEVHvvct81ajXb+
bsv2y2w9/JuKo+wszFLcTP6L4iek7iNpCJaHIAWqRrQovge07JDtLQ6vbdxA
V2Pjo33Zp3reAVApqpNMHcGAqeWmS/bgZHqTewJ/z6VkMbKR0mIbMsevgXrd
W9m9jPC38/j5ByHYBUyLSJRMTEdBUaxm4HF/g4+6y6wvCaWtg4PcMgv6RuZ2
7vpSSMPSYSUSpiYvS04gyR4RbFLF+/2S/XFzwWCiLHAhJA7soCZM++MEM4vR
g8jY37NUPn6tqQ7kIpTiL6djb4c1xnw62v6wAkBn4rhNhCAQpQFoRjI/8q6I
x5BAEk1Fq/yc3yIVDebLgPhVpXObNuskSS84QA5jtTnpnvDKkEtQDdRHk0Fo
NCH2kb6pF9ssl5s6IHBsIBCG+UEn7ycT5E0Ex8snDLISKr9Ik2paReTz0wUU
6dUuzK6WxhPbP8CwLvCS7CXrGuufNUtKC4fWgJJ6SPp9iADHcyPaRBXTR0DC
dk5Ho+e4OZF6FGTmunkKTB/9yw3Pw87LV5+O9fYcoP7uCp0i76tdB3cBIIfW
TxYA3u5xSBZX7e16o+AHtDDh3JE4MujVpDkfcww8xFQp+ChCflt3b0IjdRFh
+JTj8p9c3Yc0qwoE8jDLmV9kw8J9L0RVHrKcQksh6EQqtlwazphq0DQYG4tX
71GhkQLm+Zw2yy+PQ7JEcD2A9MDRyMhPmXwppm+NKmFReJg21Tqp09mTemcC
5JlW4F4aF1GamodyF7X8uqTolR1QP/nonmZRRblHjSXgspWzXYRtZHJHVUZX
BWN2euYwiLmgyFXdKAXTr0LxbsrsydDf9L0w25KA1NHDzrLCb++3sKD7IvrQ
WfzCEaT6RnkoeGfoIwvDg1k6EEWt9oMttol7DY2XuF9wT9/DFrSqaA9nvCPh
fsXf0cDi7v2x/kZ+fYYW75FGbd5ZrwHDYeX2hXQlYBiBnbKIcAvQP86Oc90N
t6srDCxtvtHhWd9sABqHt/7ZibXaIaj54UuAtc2KR5PDVw5LvwTXT4GnqJej
NF3FFBTCTffEmAWnLf46ifLRWQ0N4hPSiZJRDD+3j9TDhHO0C1dZaW0tqx/B
NteUeKTd+YARo33HGbk95VauioaCX9+VuynqQ1JprP7BY/Ets6P+ScEk18IU
g7NhVni6Ac5YliLrLlV72xrdl+KtI6VTjfKgz44HHZPazfEiqTRrEQ+gDJ5o
G3S04bnFFFclAMv2lmkBZROfpSM9gfrKosxR1LCAaoG4KxG9/0X7KmbNeQbE
SuypqMvgIiyha5ja6oyNWIEFLs41Ama6wkDxMQqLkk5Nd5o7zEzAy6DRVvWC
HXxejbmGUdGTDhhOFz+UuE8ePMt+vKhJ8ZqaMGwjNWbwiCv0XC1IJ9Vhmn8x
CFqWKMJNarxijc4CmW9Glb9RGfHpBPVEN+mUYEKF/5MXJ3fCwT8yz2PDBxdE
ek1hsJEKkkqhFBdrcaz6FHxMgm3RMjT8cEOmXQBQrbOrOsiQE3Ms2zmwM+bV
3SITaq6tBKt213lnIIJybTP9MKnEne+8vJypziggFFfb6XvHa23eLMJMsqO6
6cvc9Dk95/Dt77PIZIFvpF72KPPr4N/yjW6G0GL8LrNEsongOpxRyvuoeT6t
DtrkXd23plzC8HLGyUKNotlKz/dQu7CUc61VpXTFEW1IbRq7uzisvzAZit0D
KaF7Tsga0AeGFEmXrmRBhS7BHWitVR6LPbbZ0fS87GbuywOPs351OOHHcZEa
Z5fAOOf1HR+gm3FOY1FwAKC6dpxvqvEwo2pXksvVGzm+lpMFCyhHTVq12vRg
UQjNUzvXV05h/WO4atLs8XvyYdtzGmsi8OQqkdXaW6AjQiQ+oY8dXrBPLwrE
anV9P3+z0mEhV4e4L80lrNuMo4AboEjBzZjD59R8jAUbYGgcr7VWWYvpZ2BM
Dj2UjiSGKa7FEuTF7JBKpUOoeqEtof+OYwUWgzDfhN76g/lP0rfNa7iYlCM2
DU7q/an7E7Sj3Dto+cmtlSPxcBSq0UCQC2IYqdu1kzde/lyu84cRD0U4LK5s
u6vEt8HMdAXxTrBQDGjgxvaJeHsJR0bfJbEMu3lb0/rzReuzwZwJKpF6FH+N
poAlhZIbrgfMGwbXLO/QIcKkYKGmJMv2yo6/bYo97vUa1dymBJjCUSHUYIga
s+hioIWNB9mMpuPkEFJ52YrC1jdMl7dIbbX4dF6taxCTm9u/+5gzrm+JRBgw
r2rFbEP8/gGVIqZMBf+jsrkUU0pVxtZKXZriYllLe5cmmPcly4OPxxjiekCg
5nc67UOk1Gs9Yt/Ef1S7PXg8W58rBAXKfx2uvGkx8MflFs7enazgUqIKkYHH
FKvvh2B14yaLqB6Yvht+LI/9gLp85H5hpqrUBvscflkcMsEvDoCDvVns2c2Y
UmN+9F4Snwai0vEQndw4jZGxti5drUT/nM4NxHbovMgBFF9vGKWO+N/kjY7k
NakFtQsTjQNQyRDUIhZnY+mm7U775p4/JmYf+MK6ewQRskI5Qz0A3ty6XoT4
DysyRiJDaNRcd2DySXAMabRkufZNJlM1udULsZcHIvQt6JmwqN4bL54DAKeu
z1JoF2ou6QGnBoDPmPGaOkZqmdmj8GXbkUtSS5HRIx8tBo00RC+FwF6CoNcB
w9eAtT7d89h+UHUqROkKToVemWAzwTm71m2md/89a3vGyBhAf1vU4duuUOri
e6BBPgeUPX2LZ8gHL2ntSAJQfJM8/+5yQ+oGzxPaxTYrtMKCzIsgGDSUncPu
u/uj8PwpKlgfaPHLUjHkS+xn+fcnnDyKEe1FI/Ey5TT7doLrsvr0+bf+kAPD
/PJ5UlLpfmFtna3KtMUveJOlXqEUu9TdE3Y/1lPeYVMRM184/P0tZmyp/61k
akeBNAr2S8GTNkfuJ2fmi1COWkOhk4E5/ziXYSNXkh7mhHrgjlz5984FWyCt
UlRghNSVyjd40B/bnQrBbmMB7jcgvk1l24F4B2u8PBpaOpmTp97L4M170zbI
nuQaO3KcNrM86mVd9W77HiuncwDup1v0JAIDnKcTtFyq8g+BH8jCkrv7cRVr
FwzP53pioqjDkkY0EP1/p8pj+cfwMgdyVQ04A9IG0Ho8PxGGvs/Qvngp3/9F
yN28Hc8xD/ncNaAzMhuK5MN4y/VPxuzIMXJ7YHAuML0ILZNS6zZjlVWXYzLV
v8rxVICXSpuIRvv8bEDbQ20NItQZffN/UGmo6E8ZCk+bTySfjIx4HJxrfJpS
ikUxtPu/8k/zADodHfx72GIqttc5l1IGJiUkjModuOJiTDZeIXrier4typ+E
u5Gwg6sOlrhuzSWxaUGMjuPkAdTu++XyKg7aCx8XuAs3P9GrQf2q8wtpW/FF
RrKzYqg8H1FEG078Dn2Mh/+WeDi7vOS0kHOWTv+cbLbR3xy4umOWheBx1xtM
RksImHopO1vm/moSDjSvv9HDgVtoYaO1rIiz/Oa/cNuDGTVOlRAlo8GdFLYD
Rgurzb9TejrfBX0Mzn62wiDbp92652mXpNtsF3cIqTiyIM1802SAPNE11pd7
JsNypH9Zux9Eehn6Fq+S46/0RE6BPj66pCRAWocHJ7s8NANILvfMTl3cprU4
CwxwSsXbx9IB9dmkHLYdYxOHt0R3sIlm3XoVZEzB7VwKQXpRjCyqLUagUGq/
r5Xi4otNjsCIZLXISrQ4XAEaXB7kzP3ajvJCLqrexyUfMJihWL75PaBO+3/d
ce2HzxGJc2dBj3mkTflRDW/swcHsF3AnFCDTyCsq78tjnWv6TRKLhQZl7qXs
JY+UB3LxCK0SRK8gANzmPbFeTNdg6W3fAZmtJjND3CYHNJnWcZjWGQxL7UXy
ho6JFGyjMzjXFls3JzrPfRrq1H5CDMgtFn2XkG4TFicz4jvM9cT61pNjrFpG
w6yuMkNQRqB1pmFBi2pNafZVjfzUE6ghLcaCETy9wio6Cv4hS5rOiLMPrz7Z
G7YEpzcfDaGCmREsj3NHhMyQwjnm38y7QG2dWk5gpCb4ojoaBWVk/R/ZwUy2
LBbka2459X7Abuhl8X8vQECLIszBJukxnjSJY5DKgof8yuzUXIx097YuO60j
Fo13MaQCpuc8rqA5hpgePB+VQb7XH6J8MFeiuGKngFFSxD6tzngyJqhODP29
vxn7kivbT+emxCYlbtTclO6yCklMhyxYohq2H0Mqa7dJykE9zOhoeJgEQC5b
LvNVqyGHizXRVloC9g69mWB9kOgjSCEi44xBj84ZvGUqkTbS2OohgkR6SXEA
nYo+lEMcbM9BA18fE41Xx1WYsq+AgmwNMbwQ1ktyQlT7ZNX4ovR5Kls4H6vl
KB3zqxePaUkPo3+E3xDSwWfDuZhODBGh1dx+585sFLNrBQlNG5xvcFylFfVp
02KEXPjgjDwaXH6xeSeEO5VjsjFcCUeOTSO7fsyIzddn6wdY1zLd66qX1T9W
QX4xvzz4dKO8kXlHZ1Lf3xIyrPBrqGIUiChPbkQ5PLo4JESgMcrNI2FgmrOJ
Tb2hn/qeo2AvLbtPR8/TePs+WeKqYIUVYadA+dCU4TxZazv5DXhfJdVgcaR6
LLT1ViIxwRxaIF93quTdR5icQ0MhXL4R8/VogVBtbeV/MJVgxFP8d6+N9M+n
LRnlKaksb4ghiC8YlOTuC9Y6s3lyIEjCiQcArjRDWxpqIJO2VOq0l6zXSZCl
rn3QBxX2WzMdlsiKP5ViS5IBgl2Gjcz7LTRR2Cb8uFbhT9N0Ztfy+yjXSVC7
Qhgqy22K4rn2iwmTTwRBOSP40hNQOhFPYR79rF5ZNHUP30poFBE9y163d6Ns
qfaYJcG/8vVithRhZsCsgohdvPrv3Q/zFWgExwawqP0YsrpPR72fQZSmpOsE
jcPMj4B4bl+fOSqOo8zK6F2+3REVq/1CvVBDtLkp//3eOP9y+s3APImljDux
yySmE6Qvd32cq57xzf4B9ltns8QTCogmmI5So/lqRceJjxo8fcSH08JHgTah
sRZO1DO4nhkv12MLHgAHtJ5ywceXI1rbMwU6shxYtl0+9/aBlgkLPVwY+ev/
MsLI9dH9wHhqHvGuwAgE2Jn2lX/W7EKcBhB+YaIa+seaAfPZQlzdM+9zO8j6
4dfR3jT9QuabXLG8oIVoCi8yqPlW0QTQRj6jKOKEHbK1Rc3Pr4HyfQ4EmIxA
oALyP97RbXicS+W9YTYNrQEZObntmT1uBy0clvVCchtSTIs268FCM7WlVW6i
MH7ajfP9sy2Kw3GjL0O98m8t0MB728RKKvM+7dWuWCGg5wC2khPutD3sdiju
rxrV4su5IiuJB4zo3567VpLgl/gp58bzZfTiJKMYyB8oZbvogjFZIu1Qu8T9
himtV+Ci/mrglxgi/b7H1gRxV0SqhFphujq5jwmFVkivf/85Zq0KLg/Hresg
KiT+PKi+gwv75ibUSafPlKNRIFnqEv07EHyCNwoYFbRasxDdi3HbrVOUhCNs
tE/U8LYx4ncKTodq0DYIyj6Y6HX6BGhj38fnqiL54ICfez4zZilxW17PuD4I
WRI/nxLFw247202uJrx2U9UJMzkjn3oOJCC1c6GG5SW+cIL5FKQCM4AZo5UV
KRZ7PeuDhCwCYHUBbsDq15r3cAGJ2jP+uR70uRU1iyfTrYlax1EnoW6vW+W9
fdgxoKwRoYF0Oze1Ba/2FS2Guej9ivjfIVteqtjgPKPHj7yUBVy4bWkGBqtT
PAkWUZlfwA7RsBg6ApeqDUffR+2DT/UiZFN23/xzUrE1HwH2CNiwnmlnjVOn
V+ToX7xRIdNjatjlMgm7ifYmrCAgF6hUiPQTR4j8WEL3XJMwkoQv+fX7aEPA
mMgKk5x5PGtwMBc2spUBU2jThbf4FqVN8s3nIpvy8w8KiYDNpYd1+B+yL4aQ
macstWhZOBIJzhHpSjKVvv3SJysfmGC3DhEupvyqb5azZ4Wp1oDMmtOfgKFf
Wfq24yoeiiKW9E52gKyifY2l6pLa2DYAexSJj/RPUviUicwR0xctQ7SB2rQ/
4R/8v0q88BIFytzbpdN2qLTfRpxX72Kqvw9MMI51QVTcuJPw4t0lRZcB9EWI
Oz6wiLnctEad+GAiHV2Egvpd0TEmIw0m7qePvZ4DHj8IM2DtkmRrSTgsBCIH
oZJ/kQV0svwMsBExKc3OiT+zSDE4j1Mywqj2zFlhwLLjCEz6OQW3CH6bRe4a
kWYJ98y6qZvD9hQTcPQLr2YgzDxt5CQRVNfmjPSKBkTPb1qL+xuuEz9h1xtI
FKbZk1eYe2WN5xzC8KmJu/O2BMt4DbzQWC3WfRduXJX0yejXseYvzfsXmlM+
ldTTlI9gw6ilnnC2yuImRZBejbbhzI+vd1Uvz91nm5d9b982Jtxn/gPGPepD
cgKgRHCmMpgA6hFWM1q1VvQxZj1SKJHZere6192q7VWe1oRZ4QOAQ/4JhrVl
1CXPj1xvLAEceZyhOWSZ3oL7+4BEXFUjlQtKmf6dq6KeET/+lDIOrjCxY7vV
BV/dY12tx204ufsCGGxZf+tyBYlsOhy+dqmraMxBlaBnjRLv3Qom8toebBhB
LxpNV+4T5fdIIOz5TutgvqTVBzWF9ffih+pFznUCQEhWM5bULqnkXhfYzDdG
hOj2EONREWLiiYD5S1ezbcx5JYtUiDorBs1SV4LOYi+CceXBOBhEmuOJtU05
aMaLk2VTj9M3LgV3kU6zRAuspU/0x+I6WSwXq+S3U7wkVu1QTG83JISfMiU9
hOZmT13zWjFXimwQkZZNTxago6xNFv7jUbDjeCWAQTYczaIZS0vil8Zv8QC/
xKBJ7cnfYZwKxEBPLJW08KJMWkbnixDHpMdfwpJbl4ESbTPQAOyLLOCoXfnD
vAjFUUdE7yPgX0kHHNuasMpdGNuP1XCMwgnMfU2I3rslJTUA8lM/pa8hp1l5
nw1lyZlaVJKlyRdayAp+qnyRSWNpLTgX24Pu9a/CJHpbzvAdH9bw6z+jRhZu
v395U00TNnHdlm2KkDGCHMJrzJ04KblEhuoXllyS2q4Z4NGjKeggX5N7b1U9
AM3c2a9Crb7FQGRM95PvdOUFN57uifjNVjga7hHETebIdR3owLy6oHkedmyF
bZ6fMpapGd14BzlrBEE5K1NAA4711I3Cf2YU4toqasrOf8Tu+d6ZZUoLllkS
wpLi8AMUpVY6zekmK2GRlj6GVcfOdzJ3xU04ZsrSLlGB8/YjOCIit9I09jfS
rxVLkQwUkw1leJYr4z5Asse1aC1+vGERO/89O0ZbcgWZ5MFlj+SyfD9xiI0r
uTRP2eMhoNfW9Pq38/FJsjCMDdmahTG39WHwJQRTg6anUEcpUIcv4Ddt7Mbb
z/LKKAr6iwGkubOls76u/xcOo6rQv+2u7C/r12LBf9jClrBYs3bZWU1UWCVm
JaRsk9uy+9rTBJnA3PUALuYfbu4B9HT7c/keHFEjkc5HrKx57ZYeGXzvS7qm
uvJSsiWDhCa/I+mxFJbf+P56Y1WAakzYOwP7dfXt+kuqrrPz6TAF2SvblTnj
zaZ4G0Fdb6SEAC1ctvssBN3PzDMmZ15bAyTXf57fymewZLj8LyFVaFbOBL/f
wy3EykkhAPuF7wzk8ex9Dcu2uqRAdVQL12UDNAAsFL0z1LrPdlRj0tC0TVJ8
I9sfIeuph+q0CUUtrVwbLNoPw5WvYpK7iNzlxr04pTrOrt/d6ilMH7camMTq
qEzJU3mxjh+a5xnUSjeAHl4FKvXBulaIfglRB10SHOoAqR223Ppwq9c80v35
CD2xCPA8qsEoylxjPwUi61hHL0WWQXlws7vncw5JF9o+Gyl/+n0VMcP9gy8S
xPdubkd42KsX1fQpF/8RhZlXf6a36fWr8DoSEKKfEMNH0xpvl9bSIBRIyVJ6
MUg/mqp4ieEaCW+6UTOnLeER1GLslSUAH1kn6ycfjhIhkzIVZGQNHLOxK3gd
QOjIYd/NDCsy/PQBmw6tATs1T5Nfb8+ZYCKVKmW+G51DX8U39CdNra2DWSkK
myb3SgjE5+dZSkKzVCwfjDdZ8ekdczqx6wvimS1653PvVBEwSuL++stg4xqB
G1XDuiF3yQitA3uj1EDqEIljmzDDYQJuSyiNmbv3zHaylEHwQt0zQe3iBK5E
BgBJPbHhY0j6q+XxsDwdUyj1ON0rG4/GL7S7sJSgYoASfhUhQzlnKmIn40Td
qQH80pRVmVHqvq0MaVx+xUYkEVgsrW2zxU0Jr2zVqHtcLMjOXsulfwZ5rxoH
kHiCis3h/VHFEeN5FADPKN5GJdqsEl3cAbd5zmkrerSGAzyFCnWEcNg0WfpC
CJICWXeGj2EF53TvjSnvYPPpiyLqSPGuxyaRNteoJgmdEcXoydZblUCcHYWI
YXUSlfYeQnQf78Sj1wpsvsopjkuw0K8HUbCFnQOpj1T2dKUkMwC6hsXfygQC
gKY5st7LDnBTBzUbOqrWa6Y8bDOffx3Qbg0kw+2U0F37ficZXK+Dzyos8mC9
r4rqL5KfoXXXeEFvhxtvzRfYZoYi0FyD8XPfecEQVuCXkshAVaxIh2w7/J1n
g7HO9QggzQ3Ef6f5F6YPyj/Isq+QCMycrduDebeIsnDElX64hvbutib6ChwQ
nFqWBKr8kqkqvQ4ru+aZPT4yOe5BofEyAjdjMz/KIXMT51rkK0ZXJzmHqn6s
nTEgns/CT27zPWCCG83QDFtVUeDiECHj00e1HsPRrHEGOL7Owgnfe52bKGpt
27WLsjcom0ylcBe8CJ/eH26d35KxSNzKjFcUNJj+IIe8R2Dzl76Slu0tJq0s
Ubb/o/gi8egTv36ZHt3ptXBttsL6boVKrrwXw0ZnHvb4CCr7bt2VxVLVYMAs
ldWCUfUUq0uTUMuqOGa4/bB7/eeo1UhcTjNBPUaQIlA7XYl6X7ILE9I8bjTk
XAx9G9Nch/Yo9b28DOZGrmCKMTpFN9vyPVXyAR3FpfYOKF3rablwPonTZdnd
EOWKQO3r8MtSHEwW06kZl9leH23e5We6TPuOi0ncolPUAs5j0vvGA7lhWIYU
WTtTcIVo2S78zX1z8K0xDgtCJeB8hhJi6fo5b6wAzCpALjeStg9E1n4npbzg
aSfi7VG9fhHj25phBbYcWmh8Gkjy7UXijFRUS0QPyR1AKNTew6mae1u/l4Dl
uJ1SIGH9HJ1oL7oqLTpZ5hLWFhaJtyvwHGiwFpkTN48JuesNW+hrtsQOPVHj
+uzUSjCkhWynSHzbtW05PF1PITGAHMp2hBxSizVMprMJJT0yF6hEHG3dTME0
5T62em7ZWvN8F53BLGhoaOXDBZB2W7wCVzUu+Tmsm9iIWS9sJkPC5TRAVoKH
pu7TJmwDSAD17nSnzMxik+e+LAzkJhW0uQmLvBkXQtMznFPL3assVpz2hAn4
ulT0Unpm+ZnxIQ8ZTkDImkUrdvClVzA9CaeTyCpFN1+pkCjVOlyGH0ICXhdF
867lqlwcax5NTHK903+oLDrHN4hHNaF28U4uAwa+oHyPzAtIfkLb4+g9Rtz2
ts1wfpoKPNGI6PEVfg6D/Oq7FElxvhRMcf9ThGGt3lQ64meOnP2Sk/VOo/r8
TonXsGXb3h4McjyYgOzF/pva5k+zRErdoT+Tq+R6deF3nEHwyhw0idMMdOwh
u5t+Fp6tALbHTiYkhcii1XIbywpeD/pw3RT/jBDEfu0w0WoaMxUyYQFOQfb3
CVcmsvhGusZ7Cj/3qtndntegr6bZgu8eDh1KgyKq8+eSGD/v5sZKK6moulMc
WIisnNJ4+HFWcS3u6EU1ZGpf+QuKDZ22zw3p5gUvgJnN1sASuebCw8p9vYtB
YRcZknvKZy5XwNEw5StuGqCdl26VqCZdsAF+RvnVFFXAYiQU9i7MX3Q3BjNO
wNSu3pG2hrV4m8rvFOqGYsoden8PZUk2D4mBDciv/8o6oA6iSRkaYfuva6NX
YHhM6qIypYRjFuc0bTU1aJh4gZdH4i1huMkIb1v96XdQpLEBqly5X/cyNRUh
+N6k3m8dDNUilszhjxoZNs/0jG0cOM6W996eyWfsTvw33VEe6mxVSYluR4SJ
qGU3FUAWPQDBv7KuflASB+gEL88S0UC48mscd9fREbYRlWwenOv88BNPGUF0
hqaaJU/CScAXa/6ONZ8NmhSVK9r3HBjyUbTrZ5futMc1cieE143tYbW0taM9
0OgekhlyM4jNqRNwritES1jisVk11Mkelht5C3qkU3BXpVYhJLyDs0ML5WtO
85sLWKO6TwU68xvmOprfQVX7SP8/+xumyszKiBjB6oAnZBIPxBs2iBxk+Isp
8XwoSulY7/pYqITeGBGoad6Z9OLspMLevvWBG5pPmnBK+N3AposZArbw/sVC
xtaFeObVtShVz50BGpALylXdwuM6fNO8rxPliRShwNHKWOsYczx9C+FFc3wN
cP5NejyzYJLbvvOZzyzkd8++7J8oykWL84SYihzKZSCP4mzXXqXhKKw65Mqy
WPNtnYPm5pQ/RU3LwQqaOPLpY4aq4Jss+CkDb6WMqb4fQ18otYATUnLU0Pw1
umFvURLU7y0hhogqfjTiF52WQObBNvYXczSJ8cn08ErMjrAs/WxlGda/DkCt
EmATv2vhJ5Ghp8LRpbldlf/aUvCwzcqctlpI9Xcg/uSpi4OBJEGlAWW9xfRF
efKw0W7oDBPKn7KQyEPlh1C0I66Wt43f+LSKBBBSqJ1tYdFD1owKV7xGMRb+
Gn3YbwPTkzO4PyYQzEGS1TNQbanKqm+LA2XxJXoNwowf/dBckSxRe+udliZ4
wrtiriNcKkYpLW48rPgGOND2ngIrld79tq5w7I2H5NZNgtc7OdSx5Boku87Z
AnuLN/+9VRsZ8gdJ+j7PdxgsTu2qC1CHlzyUDGjY8w8xILdz8S5RtrSBQxGp
KhxPDQ32VLQNLc9QQLRTHqdY5ErmfRz3W5pBsh8r/wasGICeyCjHo+iRle1k
xbHFa/+ZJQNtIkRyMiGyKAKDsxfON6CENCZdpUPsVixX/XfqiCv8g2LhVBji
FC3Nz0UjjohdSwbmdmMMKHXfH2pE/E8JNWyckeD3IzpmRf67aeV9r/7L8Cw4
KYRxhyphiw49su6BsvkH7o6h4Kf2pcVwc0K/QBfLOlAVpwrIgVcAs1DYYD9+
l2/v3WuTpYXw1nsRsAm5z9ueygXUEnh1zglW6FkJD90Mg7d22YLjK407DASf
6XWwxh00rng7Zc+uNQihhnrA/BBavX1S9ICGHRM8nZx2aU++1gydoMyFvvid
+Am11kP3hGHkiOYA+4yjieeWeAImnX4Po4DgW+ghPmjm/msIt7g6qX0m0tE2
fw/6ykjUDMqXqFjsdZdNyqxkaHLtd3K6g89+pmLmc072Zz0JqWnv5tGkQLGX
TCHCKmo1SX+m1uGhu9CPf9eev/mTGIkjY2OhF3PWS8iO031hceq1OtNAsHcu
p3tMLyAv93/6FlWjWJv+B490vhYIkL7LGX+q71Ue53qMsc3WVfHzjbd4cZea
G2Y0RqdmumWnDgaCPCNX+c55rd4s788sSCR1t+lvxTZqiWgJxPzyDAimq/H4
NKUP28R/SBL2mZpBNqyoclgqCci28molQ2ON8tFL6Pig/l1fT2EshFKBusEO
urH7MYo3yKlqjXSji7Dz0cYHBOb0BhISbAyJVRcuLMJXCpCn5CLg5ubdSH3x
Th4kqKhxd0lfaoQwnQY/XbfbrkGcJJbNm8ZO390LE3OyA1pNgLFwxY+T2xlh
4/vYU6aAik0etXptahAI1Zcr8ae0ZgYr4dD4LjFieSqa19UOWRa7ofCscWnQ
hddPWTHG0OdrhMu909k5qIS36RimBVx1H6WdczFZOPnvVMLcDellwjVLHPtu
rh/e2QTeH9QaPQIMi/CFriGdOQSmTrKUZDglxHDshL0c7/U/P9vN2sMDOFwQ
j+U/vMSNgAgFvMzcG56YEfusoKWL8eawx8ySf15s3351vwK0m/5y32gJv2GW
dwqXwSp1z/F7TZO08kxgdrT+By5HuQ6BW02DGOETiTE4yI2ukkAO+zajKSEL
1zqYF/nlxoOvLo35+VU6/Qht/PtrtXRW3HUQVkVLYMdIgGcmu2vneLYTU23S
Y4/DnqFVM1+97m7jmHsm4ejWo2Hsn21RQhUd+cu59Yub1qDvRgOvKnWv1P8H
7taq7lU/H9uhaDh9/GPm4EVFrjxDqnYdJMiXlJ3EageuoB8iykVApsvfPCBl
itSaA/9KRvOqEw6y/tiaD7NL2Gd8l58FKVb+vwCzJdP0wmWiaQdgI7emY4Z+
bZzQzjbA6mNiNF6fr0shWg7Y6bOA+pGUcjDE3fZcFifAsht5zP4UjuFHL0Wd
ynxN8IBRRHSViJg8qYboPahEyyW/ntHALz1ic4IuER5pBoA+ozJIoQqCgREX
zYy6FaF/dLmP4fIjkfaja+Jo5uUc31A+o3QyK0DD/Nf8D13CsMKimMeHwgRk
20gUxU5+agaholvDwURmNy96ytMpC+XruAOutVsHwbRi+2aLv/1T//seWclV
0cqTxOH39KhnCzu8rOfw8v35qS1dVRXMvXv08tfTR5ZGsrM5179lBTeX7Jbh
z0LkQeRSiQSo49eZwLLCtqQHqB4l0s4AC8d34wHmLdfhCQxZDNFAOdQmCByY
kMYez1kWDbNw1P8zrOSmC8pxCnrLUT2Mi8b7GPknnuKpXpSrAgSdfUlIdJk4
E3wUt+9h0zeJBKg+cqxoP6OmO6PFlA28yyVsdFTpLznmr/XGe5kJo0OVwcUv
lbKrhRArjHeImG7b98AzrZeWftP2Lb02UVtlUSxqEUSCN3fFONmGm7pFgSms
fW7gDiN+0Gtxbe+nhWRCgU2+m7ovfCXC/KqOdBZwZ+4cvqApXdxYTQeZI1J2
caeKszFDV+XULRr3B+5v46OYtIwJK7RFw+L2Mu/vWRaykvDmL3rGuB74wE7z
GDQ5fatH0APLRS3ciRtFT9SI/Jr4Pl/34QXGb25t0nLvN+N5stB2gnrsHXOC
YfyWzeVqRNvrd4oCTzHkSbAChYZ8LIbXre6CMs9HIVpeSKyt/rX2XtdHZ5Sw
1lO46jwMXHy6ghcwuNZ8QSFQkpMkQC4NnL09LraC+R1cDOMlryj0SBDp+ucP
vKTKFqNXjhgNxMDBD4N5IjofosccCtYnLCwbwYxTyyS2Q4LOn+Y+8or7aE4X
pZpRNPKZtEPpaOAquzY/Te3FsfxhwKzi/LOFJ/T86G0zcSoTP1hUah/qq/qL
4ZrQcNd6am2RjdAT/EndhJeRKHA7/18/5o8kv3Rvp9BpGFgegeruXIPU0rcR
0XmwdeM+p2N2a0jmDg7yglSDtink3Rv577wcwqidlS3keuCylnRzTuO3ITJ2
cipRI6i5j5XmSk+PiRjDV1g9nPXn6Io0N6DCCPqAKVPWw8IwftmQLvmHaDjW
g6STkqHIrEBC+rctuoeWYsCVf1ZZbsD1SrQfFXPfvthn6B7twy1Jcpb/vMJh
jpcMlFvoq3gvMieE3woBLAGQFfhTZf3QixiM/9o+QyscQD4Gr1+yrMVGzFg4
XrI7SFsrsnQ+r553hLfhDqBV2M/vCuN84CuG9+rCQiGekCHwbkt8CXw8RB2H
HgOGRWI1Gy/HzY8tWdnUCrYPI+CclxJ3O1mMXiQpjcMUlIO/6z8p2QFSzR8V
RwRyTkXXskQyuXoWIQZBPUyD2tv8p5TKKso5n4zDI5+aTW9k+mJXQRx4K37y
uvv1zn7hW8RSvJmwKRVxbbjn1/6pP6Hz+xhWGjRjj6hYnm50ooA1KUZ/xfZY
ntjS3D90lbddJ8CvN8v2lJeOs3la0a2xHwE5iDU+SvdDLhCWktUrI4kL6qvD
HHgpnCHkmojL12Dy8L6IHGrW2eGsN/gx5fgVk73mcAuuBN7a5vOFcoRUjB5X
7Bcz3EnLRncVfMWzYvXMN8y6o+VheGN3/mw5wmsclIEAMPmmic5NpwvW+QcG
zteFyTdh+mQP1D82erSksdz6qSmfo1pPEMBs1a1o8WWZduKbzIPa8Nym7689
SiSDZFF0Pp+thps5XrgXHoAz2JFDyU8Xka4EyrCXgh/a35boEiEg5kZkv0qe
JGWP3YsBE0ttOB904qfW4br7lv/MKs7hy/cMe5PmPCzwnexRXyGBu5mPRNnH
oHu8j1ek3UqsNANKGEuDE9vwVAnLep1+FBv+Hp5Ahc7apJFqYLD2+ehjLVPu
lzp9CMaYFinbwwQzfe4maH7f7C3CmMLMu8dWZbtccvUF4M6qKpsQ1bNa5WQR
qCGQ3T8ZHxant5QR8XHkt86KUyPNPeXCGIQuTesfcCTSLUylrqW3aheGfxKq
rs0/xfp4Zxl6KfrZBfXwg+8Zt7FPwwNKqDYxoCqm4xAu5CYrs4SCFKzQp8/g
8ia4NxQn2NVnQQBiulj6M8jba++Wpn1oZOBOra3YaALu2JYwXvcDwYfHFU+l
CHibgGSYrGzxqDkBo76Qiy1V3xcvxb4nE1anRHw/tUldIH0RI3wGs+Lb4xG1
DhqbKB6kpl4TYme7ehYDcpC2FrhzstvUM7ne2vWhh2cwwOvMCTqkDCNHcpy8
l1ry5oRYr97cBZW0UFFqW7jWJ+OLaSr0+WCFGT9HKnoU6RXizbDW1mfYozbV
VhlhKK0nhA/Cb8q/rBVI2xiM4Fq08WHwDye4Yr5cLbH/CZ2qoPN0IeqpA2Yx
h6JI4/A8bPmBOigqnTeMtnzxFZ5omczHpwUL4ZFdiX4y+7rVywvvpLpvtu1x
Mi38PDgPu1v+AknjOqaWAIRyG8xrgAOd+LP8n8dpV7oqoBwlinUwLXUA/6Ox
hIt6o0CAnkTjgF8jpjdJ4YravGah2aSSVXTRAIAWH2hHoCqdOeqdzuv8DeGa
dK4sVtRgt9RGmvrIFJJkZizVbIPV0lywGS0JgXE5bNuguGQ8pNHDP9U2c1Yq
RyJnp5h5JSXIc0Fa/PqQMu10Wj8UUk9nc4Kve2Fsf12M/0r0cykde9PMPI2+
DVryk5rQlp+8kH0UB5u2LFmdcCiBoXinUpk3CQzG5iKOsPD8JvWzS7//7O2I
i6e6Ku4f1N3oKMWNajz7A//o+EYY3nDFz5cuMBCsYbxfVE1mQ6LK09RkBiSw
BU475BPQeh/XG6sp0O9TxPhQHoL2mAeAGO+6h5q+lV8k872wQpr9o8aCl9/h
o8+znduRpabcZciIVoY0YW0T2KK5LklRiHTthF1dq3pjtZFZnZ5KO8T3sfG5
w7LUnerCYHB37grUb8hWhkgXxS5ouU3mjJj+U/dDMO3oUtSX5pr7cMMiSxf0
xKFiUY2X7To3wxpeCDpwqkf8rjmYeVAmPMxDtgSo8Vo8FYl5XFiTKIXsbbQR
EwyFU27eqaV9toEmSqrEZJu9Xl2l/8P6xl2Xvh4HCFhAibmZX26xl1vpzJyC
2w1yDoSNYsLC37R85lU+/TxfpM39nAp88c9yjVUvDlBbiqXlIsjGHxNU6Viq
LyAaVFt66a5YukBqQvw+XutZlyzuV5I02f0jdXLT6Da4EzxxElkV2hfUGLv3
mjzIYgEFg+I0YQ+IdKcmTxuM3wBtkH+QkuG0LsKxBp7Y/F2gM2/xKiYpiOYx
jiRIjU5H9cDmuklJ1kt8JsGjQs6D8rkTc75YhbxrKUeE96nNptv8Kacl1/f0
QFOvWJCabQx+13DeBfa+zXXxjeJKEwRcyf2vJnil46uWVkUpbPFeJLIa7nvA
kjozlWonTGqwjcNffQkCU8vQGJop71Kpe5Tq6Pr6PHl7qyvwgSJ/ODcotX/7
ZZ3xw4cyXNuOOBuQtgG8JFM6g8L/ljN4DUM54eSIk7BLWDkai0wW3nlr5ciE
y3DQXXAwRypXXr+G+nsqaEAM/W4ULw7Reb5CViOiTZwyDr0BE/2oJfzhCmCr
mOpkdeHnp6m83/vv23I1PcX18zKUSzN7iltbjDZDGA7dtjKOM+hIRZUHqDIT
XGzXSGMYcdqZSRUOiDm3Ev/Bn6zegd5Uf+eM9Vio0plk6q2i4pM1EgRkF1GX
D5UTkj7zgDbxtGXdzYg4Nqd+jz80b4QxKycqYPk1+mJxu6KNPRbkuSz8mZVA
H1PBAx42v/6S6vSKiiZkeSkDWZn/tp6cz85RY0KlZptuUVGshbNwQVLOW/1m
m/KWvb/M1pqMKfy1XeNIKrnv2/6pR+C2wk4ozCgbCM/fq255PxB0/+7vK1tw
T6+w9vex8LYxh6B/y0l7vmaLfFD+QXdzX678DCseZ+GQzuLe+aJhD7ZKtlwQ
hvJn30Sd1Fr2igoGU6IOdu7Kny7RTnhcFhorlldYlzmaXBySiE3i4wBt4tyt
fSwGR5YIXKB+T0FpfgPNnuCsPfA1ClrybLyiXJr3nuQJc2kuz+2pg6Nc/+im
Jr8PapmgjsWbaiXthS9K1O1GyDiVUNFPss7L+c9qmzUatbYaJWU/7YOas2T/
rQJZGgNb5xuppfKCCHGtcGzRxNU+v2r7kqt00vf6RuRKmNL2dot9vGTkiNWi
Wl9gWRLE57YJ0Z7WLNRQ129Jnnh381SSBSixhN3awifoSluYY5OEjMbLwvnt
HXa2Af4SyK6KK4D4R8ARqaVA5FzC3hzLD4tvt94/ZLuQyv9I1/NTtJYqF/iS
wUXmQxgwAjD1ploQfaej8acFv/MBP1B09pRgC0VzfY0xPGFDB71cqY9ySHi5
M/F7tf1YlMBrqbQsT5/a+vRdVXHUBn0r4zt7LgwvdyX891CiMoiwW5+L1dmX
sQRmKkHMChM+kwkWKIs9Z1MiO3tyjaQbVfvPJmPAjN5gIx303hlqIZn9AC1K
I9GQF/Ltk/NTkFleppvtBylJlmOKacnAySBgBFB3OE0aVgqi6hUS+zqmI0Kp
3Va6QhB1iEctuCQhtgPs4nb+n91h5Tj5yACyfqNz6c+e9w4i1RqCEMyaMbOx
fFo583v9UblaNK3vmWHjsO6RkCxgAcd2D2kunwYYFY43BJ/B2exK8tQnHuX0
PMEe+DB2ROdwnKeLpaLVxjUs8ZUG4a4hbJCqQ5JKG53iCK+jobWIkZIWrzoG
wZ+0YPRnTxragraa8dSARQHZG1CjJMdBa/JNJdSMUX5oaL2LnFLc09dhNJQk
1g/sUa6mjS8I6DAB4MNA1Ou/Mx30bvM8ah99iNizyOYhaowFGGbPP1tkW7fN
fxZXsbNyrumNPJ//P8Nr4TYDyR2CrAL2IqOgzXMdqis9R8EC5G4t91MkzELH
j8iV3O1dFPb9FYD7Jrsnlv8v7kM5RiKupCywq+rRD5Tz6aS8wKvqW5XpK29V
+K0KSM/Lqu/hdStVE9yMPyL7FV2hNyXhTwd34wo/n7BTlzmEP7PzE4FYYhP1
Nd7JZgrX3B9rr3TCng1D0cwexTyl9HUmpG0dO97ejjoTZPXuJcbA7A+aKpHl
l9tP0x1LzTz2UwoggLZooS+6Jgj4YoglgLPLbv4YbjqLXNVe4ACmMHyr57uI
2wD9KpGqmdd25+JqrJJzrfL9ccuy0/JaQYaIcvA29FtoMMtaFPGJ00+lEKnO
6QFpi8LxrLprgy9Mty0em3LiM/wnhZ19f9eCMNqI8y1obU1NGW6X/aihSkf1
SQRTn2goY7P5P2zKDTv2QqzzW+ScEOcOmIHbiuMJ2CCvBH3S8BP7ZwjZvQG1
vBP0IYuXVquqk01+F1GXpfoKu3jb3kOyrRet6l9VRrS0vcfhque5vZQ+XC9T
5L0pGAl/sqyOuKu0jNshasA+/npSWhAFc2XUsQcdRZxZIqhwNph6vr4XT7zF
lDWcRkGjwj3K8AvRS7vNtg3/8KN3cJIeZOoCk0gmw03WvQIKIRfncgR0VQDL
ikzea9DEsF1Pzhypntf3DMwEmHQ03KtZxar3203ZsQytw5dzGGziPIh5KuNx
zLxO2FHTJHvF7/zLl4G2yUoj270xhqapz+JCUmphi2RrckQPWCvmpO9KdnPE
FrRBr5h6LzHOT9svmPjXgITfR2Es0OwFa0h5NH+Fprcr0lD4CZcb3d4k4IL3
Aa9f2UqGzgcF/bIi/qSRC7NtfYsJqF5Q+c4FNlx7JOQmoO+aNyPKerlakIoQ
JRjXAO4mGdcAwFhA3eM20ENbJDEAv/UmEIlLzkz1qhjMsiJeBaO8oo8J1cQx
knjNtx8qVTF1gijm4Zfuoh+WYA72WuT9dGfgj6ZVdTfna4bcxQ6wDcz5WwwM
AKubsGJ6FG5cSEc2MkeyxPAF8AnC4ZR5+IATC+3q35RYKBIdTAWkHLHVqL1F
ZqwFHob6PYvTlOCfhlvEHS6mynbVeaFjv4or8oNAq5tbxCxv7j2tGzrz9EiI
9e4ZVdzAdN8xPnwS15OYVTLS4ubSBbwLQUpsgK0ODL9S5E3qYZ0Ix4rUvLjs
YZgTQ+SmzmLSj9Ap5ou96j9AFCmViMvGHOQyp5U4Si2RHdc2XnEdI2AWCHnb
LNE0pXL2FFZRFMarETRnEPcNWO+xatlT+sqsag2L7JQ4GMg2FCAGH6mF1RhP
zYbyRKgx5XzYR3jDd1aC0utNULiupqO1xDKL4aMTiM4LYUGw2koJpmwCgdl5
pSbZQ+OLFE5VvHDhocZNyTHjhRT4T7FBq1SZ+0QkU4fzb8ybG2I90V3sHPia
Xci1BOnT7GQXhKVAnbnmKoAekcgl+v46v5IwhMwTa3em2Y+SoaO2Ok5bUCfW
gxAo3Mkm4LIS1NVGltwlyPsCeVv1SRG0h7SCzEdArN/K7mY5J4EclYSC2CwP
VFD5tp/d205dk+dMVUUrb2p1qYctDvpasi8ssDR+QbaegDfrGEPILUyMNZlS
94UjTuYMf513RW4W0gOItjWz3uhbAvzGl+hydxUxSFa/GFSGf2337bkCkbFd
JfGLdB2+E8Mc7LlkjlUtL1mSa/GWeMOyYmVfv7gdcxU6e7YCYhKARzHuW8zE
epsaeOF6nm1amK/pM3tR7SBYoldsPgcpgdE4b74aX/HSx9lDeyqMJ14QfFDX
Sso2PE4T2rpy938mw4v6aX1sPqLsOm7L6dVu1aBBOCKWt59R4f93wj3toOja
0ysLciPSc27YEb/A3C3GoxHOzcgdvoA70yunLbgnnW2NmMHDrJ2SErwj+lNn
DSl2O9F+8NFSVlgjAQxurWWMHIVVA4rO1BwDeYtKNEyu2y+X6vGO+R83xDRT
cc8LKAF+ERtuVeumd/8gaC+gMiXO7o4ivNZURc7AKnHnKaHzyNO9udam+slb
TkYBGwE3FRen8USvsBOOsCRM+91MrCHZTf4pjNLMaOPSKP/vfzBMzGv0D0ql
OZilXnV6AB9ZSsN2AyAQDLdBgpY7sQ9a92+UT5OonxZ/Nc1uv6zd6pCaXbIg
OK5fBcERxkRWDNgDpIet6LelrThC4b+Btn3dMCkWJ36hUYDrnezHXZDKL0gE
w1i0IcujVREkVn+SofHMc4hZQ/e6LKglNTVGaQk7Uuc+fdQozl8zhZRcp0fr
JO2xuiKD2hEomqGrgPzdh79OqFMtcUcnwrvyG2XnI+XuxMmL/UApuIi78X0r
7kiDP0LGwfJsuN2oiUjr7FThVQrocH2o66bYtFU0+MrDV59wmteBAGDkFeBe
RGjf/60gIh5WaLsDxmoUtMFjV7wqy+Qk9vEZXhfGgBg7i0ysx3BqIxW6djzI
GoBhZmYgLuW9iu1RyKTooN+6XMIUdrIT/ekolyh29uG9uVV8NNjSoC/EoKlo
3dGSXe74F+ioKAGK/+90Cf1lle0ij65uQF41UvaZ26MmTd/4noaHJMxERv5q
eaUr7CLzCAR7blgEtA5q4mM+pAJIonWZSSkG8fRK2hCF3kCux7yOPbJDyDEG
E0QflQloXltxBvIyG95DQ67PkN8/MPa4mSw35SCgHH2egfHWCsOzfK1JNLC2
ZTYKnybgoAMeeYW8udVrO6DT+fB1wxQlfnHr6/S4oJvR41EQd+4m6uKKx84x
zQ/pqCCOOuEYZiku1HwB/QdFlKdoNY/QAeZSWE+6eP5p4mnLyPiNNSrouJkz
hcUfBtKdld+yiVK32z/PiPR5Z72rSXBwY9mbGv80hUk50xjjwzyRtHKdeEfb
1H6p08Dana/gjqCZxunqipDCHLInELFQL7+K4DM5qjUurHWNwo1DYkr/0Buf
li8jWftPnMbmrf2exnSwGV+3XWeXncTiwbwz9tvyzbnOIioDaUgdthYmaSNd
wCelzOJsygWPrfo2kI0P9693FCz7MR8Jn9lWaRo7CQo7tgdE39E0aI11vojQ
S0NczDh7uK98NmnZY3Y6SsUNh+tNDmXTQh6kvanEFDrWqkSlb6oacQqxeoL+
DFiuu7WFmooSSYLW3Q+jmtcjEENG3pE1b1pDv0YhoMn/m2iOfarmTWTy1s9z
aoH4NDH5arY3f/y1S0vgybw54qKp5BM1Lz56//JJdLGCBrQiDMX3zmNqbgOL
FwySMGCUQLO567/wEbwztzDw93hLXAeCteH4kKYCaPCVN1o6wXC/ks+NqiRM
ZODbd7NnhA0dHGEPNQLjCWCSNeG5a395Pmzpu6YdSb06odRAwcfkY9PTL+y+
ZuR3W9ANbWcJk4LdxLOBD9NFKvwNwTC8R76reYNlo67E9KvVkEM3NSYrg4vI
oYOZe0Vc1mSi1/7Klb4yMakJx/t/QL+bjzBfnryDMHmjGeclIbPlJQbzQj6T
32jmdaGof94HaysOOa12LZQQ+OI5OUjBl4wtfEfL6OgkCZgNKBHx6K2Ktdmq
Yrt+qEiGk/VeCrFJ8wZsCH+1FstIQhpuyPA1Ibq5/L3j/qkXTLSd28BpsgAV
iKoDLZ8NS0mo6lEk41V7yHtp/3Q3y25O+zv9/ihjqfqvAEOYFDFCxglYATl6
43nQ3diwfaellcfK8Bj2mO7E2R7Ohs6Aym+6vIFo7PdEjud1NCCu/HEkHn09
NklSFDYRcYJ9IyX+V7pJrUY1dORIHRce+GkStFSE4OY0/WX+G9thfPvwQPBZ
ZS96xmKhmQ8YSBSQc7lu5/VuuL1Q6z4jzx2abi43MTEP+CcHVt/FhOVjVpGN
FoEsU6hvTp+26SB8/SWUJFA3CjL79kl5UmB9FVMBWcQmSnCrz8zN20TWINCR
Sxt19ZOmbkYunUIc1Gt8chQ2HHILMgJCWy66yWsm3VOT76ZOkJZ0TXCydQFl
Y3KubMByc7DETt5K5rEVBMbBGUjL9c7sS0ttlmwVHV+cXKTSI6RgZDiGBAD6
zqosqAGbcNUqUguiMKNxFhzSqf9zXbhk6aX3o8+tqKqvqDASRvsJtLXiAhpQ
Fd3hcIBY66qmBdCCJuNJECpV3zZaQCRltCAf2HFC2yJkvVt6cpaa+6WPsqgd
/S5zaIiCQSO/NVKJyj4zU9eBpXCioy4h4f9BNQml39NtoAp1WZvowuiibx18
4DAj/XX95BKt6Xv33hxK5AFQ/cZI0MMGFNnmiW/VQKsHRr8NkCFEs69nIiDW
FpG0SDkhAcdO6CDYzs/IAwIjMVQ5sJpwQ+bWJoS0FjdWV8AxSeJ8yBiu9P0O
EC4UOSO3pfwGtyd8JOhzc9JtOlsIdxZuvn7YRJGytrFzV1jKVkI72ulhud9C
NHT2p76OK3H87q4hhaieYRaPgzf97Ol11xg2zFAK0i5ij/CAdK4dx1TvZUaa
m3rvyWnqG/mmDFqOgHy7FSuboiGF2PXuQhAICzIb53z7pvK28ObMAdCt/LLE
TjUwmx1TMisyzEoq6kl7WC/NYtrYl/Wk3nfT0SwQsevzVSYNHDjjLNI6ZWIa
ap4LDbr+yEd8yWi6WerceXhRE/NO1+p0JczWVDDQzjxjOqUALskhqLieFkAO
pZG0oSMQNbIvZT3lh2sVIyUYTIgSxO7GUOhioz3LZnFqhdjdTe5k9x1RWnRP
legywg+ucY3XOCDmew6TMIkN4F6g/0yqL6yxlboLxRiZbBfmpEr2dzlm3DWh
wrjzQvqhxF6WoeZy303BGPzrFIDqD4XV7yUd4TKsd1nTw4h50msZSYWrhpF9
XhRl7OcJyCWTPMocZLG8f13CV4hK/U6YBqx76FlrJsfAN3aTro2714VtmLXj
tpNz12JX3URvxkZhcDul+T2T8KPQsbtseJAXWNu2LAlDbXs/4nbDlwYkBnWc
d7ZtMRw0uWVSYIb/UCaBrFf+xOsQGcJNvg5U6GXrtT0z2NKKeH/PSHBhCFJq
xJL01n6nc1QTzP2dU98uWBACpLB/RhUc03i/vqvREeIlS5CLvDOcC3hRqqK1
YPpOqHrQaW9IV+KnFP5llANMjXJt5na5XMnKmfJZAowcuvgS8HaojWv/+Rzg
xnYw4Trchf79CF2qzjJuP21cZEJ/aItSDohAWf7P1cesMUP6dyy4rWS2Z/3x
5Rpyh/MQloQ3I6Xjnv+he17lhwtIE9qmaEMmrtDPdIl9pDqiJWE0y36XDPZx
oq+yhLkJv26QjjbdR2METia15ENxNn8ml/EwPjAQiqGoOW0pnLQWxssxvRTi
tClMwlyAx6PtK7eBWo5Z9XTKl8zV0S1t5VfkIK3IxvjPYoAxXsnQgavjbA91
McsoMaPptGVAdDtDxMo2pMFL8HWONDFyv2fHz6nNa0cUiIDyBsTq3cfVytQp
JjKgzSfenGJ9yjYuhDktbLl4uThzc3r6+Z+Bbyv9ib/FefAFqoTxdnesa0CB
o8d6gKCLW15jGZoIB6kDx5XHroT//zwLibJ0HzydfEq6vuHq46tZkRRuq60o
CvxM99B/pmYBoa7MimYXX/EFBcVt6l7VGpTTiueUU42PlmSce+eKTRQwYRV4
2+YM87fqtqK+00cMSwPekNUvbm+6P8D6G0uw/MsFSA2BIXyi6WEADtBT3prT
8Iq/Ubalh2gJs8rZAg/K4LVo9hMsm/gaZmYzhpRm0tsnor4RKNWZzQmYR0ex
ugV+Dneaogpr1MW2jDdepmhByeKzDGCC3L6Q2ZWXNhsGJEnYoNGyGNHKwk5e
5qrZuRNLZmOnr2JqBBbq3rpqESo1LJjHl5fHrZ/VgSbMJTlGQ+mv5BWYKWtX
UAPG+dGfbjDVNXGKQ+CMl9AiBf+Cg0fRspXeBl+6PSI6Kt17YlWRmtGPxqUI
ZgB5uwzUawRlOllR6rcdDQzZ2HFMx7/OnmvcprT29kzojI4UNRvRKsHA/D1f
wKjhffQyOM80ugsTblI4Krhq/BpsNcJwpwR+9FYIufXcyZSLxELXpi23HgE6
0tP0n24TFvdPi2AU9c1HGAihq5EDFdT/ZcebNl4v81LKBxmONUAPQGGK8orF
hwMCRqeItSwnTjxV2htGB95kK0Wnb90KnFIplQEdQMSNS7OgX/gWi4BDTgfU
ltAWLc6Gi/wnRim9QH1/kF86K7x0w6JcUnZorAtRPV56yztu5ODgIxs4vIz/
B2EBiL7/nUXzZFtEIbdOspnfkVTjfzGtLesw5BGNb7itis0mhlopSNHlUbD5
T7caRKBFfCEJZPqh4eAKORhcMLdOyM03IunyHsNW7T6v52xzMPO0etheZl47
ZHtYduT8Ifx4LxkDKASndtI/TwtbBlOsc+JUKPb+4D4HX+aToM55kKVKdfpe
eIZI/m75pLXfpKCdpJCHqn1fg1sO93HA3lyCf2EQOYMX8cmWuPOZq9O93IFw
+150B+t0EmrQWYehaTTvL5CpXtSsVMc87GLOG92r2BCJR1oP6YaATWOvAZ9T
Ej7y+MP2uGg1Z9SkvVD7/zgLf4n1Yu7QmqHZ/WoGBb/HXvRpXMWs2XNRu1ju
eMO0At9w3qG9lqBLdpx/VwYl05axCNbtq6bvp2aPma7oTPk3EJkL6wRGZyjx
bOd/kCfyGIWYLsADhO7oFe7mxUFlSTR0/8cDV6/ZAOU1MQ8oJff674DpI0O+
APBxJbwlE1Gn4t8i+D5F1ABTVd9/1/EH+sGi7FSj8CaMNlC76iW/6XA4e14w
SNNfhn1hXjr4mLvDmx4WUAsP4i7fR2tgNsqdjm0tSSOXmONH0dBkzu1OvQVW
STQaGAXgLJFaXwmccfSP2lbuOAlQ+mhEZTEpoGD83vS4KlMm/zK5p8EWNj1F
ei5Bg7ZCzV6vwIqp4Lmg/6vRc/Jkcn4OzgjLpHweT2IlKIyMJsKZ3zzF0z7o
gI8aW/YBvNkoumLzoLS1R6kMWtybM8E9Pbmb5ALf4s6TyI4nCob5Rv5wkRQ7
38mSTtxcqeWVCp2FH1qYEFq0itjNi+vh3Du7eAoShIt1gm/aTMnp3owMBhQu
h4F8ViM/i5UZa+ER7PknOVYIJuGep1ze3JHUFsn4YbEl++13VIa2bjD54Pxy
oQfCOe17hIjbel9RqLujAzxlCl5OjqVjpbE4aY51Tue6WSKFkr8WqXM5DuCL
h7kxXTcEwUlhRYLU2ApR3Z5uI1rPhPMO0IhkZoAZ4t1O+H/O6DN+kKHcbS0Q
0yE+kbJYECeti6bJdGO6+USvYJbvZMj/og0j8C6/0FLULTELoNVhJkN5eSuY
Bw9PscTaLy7zEHjBSSLRSgDMsjR365dvE4l1D5GNOD7sVDrS3+iyNAJDgKQ2
2C1D8JIHj/pdUFejdSJ+2Uzi7Ciw63GkPtuyqRVdR1XjvA/k/RAkhMPSjxrM
RKTLrnU5hRQ7aVV5Q44boehEvXKqCCyxmSXFx3ru+MzXRU1jfBfU7NJPgkon
xcTtnwM/XlXQ3pUo14m09j7+G43OLr281ZlPAVi80+Br+Kf/CywjL2kXC3zH
mqJ4QYr3lcr0gISaL7VOuPkzXQAozCjOmb6o0qOaJbFX72RSElHluONGMCIY
+2T+CQvVqQegOtk7CAN7f9UcHG36dw9rw6mw+0fHIjeGRcBLXn/Egd1G3ynY
mZ0CDLzU6D8BYmsUtOelPBRfKcClfSFq6Lcdd6UNia0rh7JMRsZhL6K0Ts3B
Ym7vISiBiEi9tzoCLeShYINWcY3LDWi8pWQnQIUXbypEkXodhTRKSuvW4R3C
jipCdM2cgL7I7zByinPlFfCNw9njCuStbuYNnR2G27vX9pUkdv+GYskkIm+8
9BLZScWu123sYbLson/q4DnRaoGw/+v7fHGqJOeo2qgUK5jZKPq2uinzAPud
Y2jblZ/5a3wU6fVNW5H1/z4z/n0YeXRW1pLX2xt+dr961LKhwopi+GxqhghY
p4P0XFcctcSxf8lA0Cev2GluBpGKlDp4WtJuN3cIFB8m9xQ9Ntap4S0SpNdy
7jtnNKJ8TnYDBudw6MQ2b+MuHOWRoes8TMCCKDC/jgeZHdFtUW1Crl6xahUB
6lOZ69q17bQ7GzZVVTmBIjkhTUnmKKUhhxUmKYZd2cpwtnPIppSZddpXu/E4
FbEhJzmpHljEX71BLW5D6dbFhtOnwacm/Q0b6/0TgtbDLgKr5/Ek7M3guml6
Ei2Y56i90AAoFeN/fWMMKE/yZOIU49FTXtJLoN8uShCoPw8P52jPz5fpzaxS
eZNicgtozq9MsGOoqAfEOaJzPAcUxJQYuJMIibth6Gqzo83T4vmZQ9KU82VV
T4Z5NtsENg3SgTo5K+ZRY2+K8VKe6vwuwzfB9nF7ozoQD1/7z2siZVBaN0pk
oe8wxsTov3VbDj97S8A2VwZyasU9TtPdnWKeHTTgBdNkYzMm1fM5aUf7mKS+
ZVcDCvPpTnyZw/XskvDu8VohKP/NfTnS16PRP/irndoxT9BJq/XvCsprDklv
sNuDqpF2nV+g6hsVTC9g0LHOAbwt/xuCPeWEXz+L/FVAl9hQsl+xvZK0R2FT
jR204O/yOo7lN8aKiTxG5BTojzMc7+dRXCbXX34atNFmB33kC1PRn0ptwMq3
T6mBnH0BEXQ9FR+0zwChNIcfAAOYKa0Y+kdbSfqfTafnYl3a3uvE3oJzxMGI
eRO0ytA25gCAPuu5uUdCT6Q4ahi9miuQtx9MR/zUF3k17vh53wiPyt2AiLDb
20+llEkjsRoMH8A2x5XLAU8V2TU+8E5HLfiUdxPUS7+3/2l6G/87jj2Yf1nx
bvznKcw5z4RmQTKnfHJNJPHB5ch+9N4IdtpV4wxARv3Ohlfnej2ImQtz+jw6
J/jBLpxRW+MoUT6Ywn7AmUQvQ27Y36VXD/rBW7EwKJvpmRNyH7c5AwLCHIOg
aIUMdg1gQ5xqV/uXtw892eOBmaFBxLFNHkzyY7+ub/oNWT/gnxzC537aQr5m
wOrcg2KQNbgiwZZlg0aSxZt73pTUxUlOoDiRmePUqtVwwPpfQL6UWTBwwmSR
5SbsqCvf64AsoRHm1nfLVQ2nnDh3xQn39AU8eKVRL1YlqxrY8ugYwpyImUqn
pQLi5Jsne3PW5CqLuOMhXupL6OYLMeyHm/Ipt1lug9TSA67GbnE11tV90OQS
IdZ7mhmqZhJKG7dwRcNQJZiY+usblwLHLSHmU7fWZWdv9cppZGu9IIiQ4mbC
A/56Cx3X3jnfKY4NU37Q6c3enfbRQRy7vEpkHCHT4xvZXjWSfMZLPyiElkps
m7o3bzWQBjBZX0ICJ7LIoIAN0X+8nwQH1cEeEgSgSSTjZlYTvJayMlCZfv2v
H7TW/+RFKoCcFCwiok6ro9hZnczxBB3O10gw2AU6CPgYXpGPzbCtBVt3obBI
VIoa7vkPSrGp8bPTg+GjlO550X4EXdlDAJtIipbUEAS4eKXB+7AUfLanUoi/
U78qCzLLvs144QHdScoW9rFBAYHGEeVztOR87nNAtIWNt7mwz817oVeEFniV
AohKRkGtc1A4eTC2fwyt7k7QwwwHtJQntzyrqKJBJhccPvbaHC0Etst0FF+Y
SZIIauJsD9m30XioTWqCb+fNIz8+9JBIAHMh6dvq0yLKj5wSAg5w+VvomZvF
5GswIpVM5goYo883fr8qniLCw4QwKgG7MU+u0nybaoOS2+wWZXFVfVVGNh+V
KPPXh1BgdKh28DGVwZ04X2Nm0FtSizbW0rlN4QbiKF8fpe0HS9j8gt6pXaip
IDhj2RlJszw3z3YI/WBakRClhzc17e0I1dzLYVBG3AT4u9cTrQTxIT2ftqpv
FXA04enAh0UxPvSAtr6jsozk4sw8s1+VtzfRkuEQ0Dl/EFXEYaOUVg0y61zy
+zan4AVFt/JxHxRnnd0NMYTelPciHlCitdG/hQZgDmLVlnSAUlKXrfKRYWfZ
g0PfVrKe5GQvOk4n/ba30uXIhCIQTKFthgH62QM9GRklkyuv77i4ItKIO4Wg
mXs9w6xv1j9M19ENw7PzkqsBdoAFwLqG48m7GSDL1tonAzuOLmSblFKOowKd
aLWMvDKclEbiQA+3iVi5nYH6orgtC6ghgrk1Ll3H4+HvkH3lec5XRz9p2nrb
Xl//bw+ZE6rgl5UnQyvYpEUUAS6aQt27kZ2o3pyDzAlxwlaQyD1sbejnwPB4
GCOOJjG/c/DLawGDUOx9nEMd5ewmdDA/cwW3vR/wD011qSQ0xYb0m2H/ovCE
C33F4gZBR1q0fabBu6Rp8su8a6VMZRPcDhkz7CvsQTckaTLgL+S6q/2+rPBT
zgpCJiJATrdGdDiMyuTE3IaSHFzGRDqNAiePlVJWvZcnoWftmLkXYZn3hA+b
8aEmHa+4lZoQRUiHvs47R6xmfvRNORjuAhAo1X2iAW2KvtFBMPheE2izmeba
xDF59EzTmDJhjF9PEWhZqyFX466w4Pdm1oLfpsmdIb/YrcJOzOEdWcTOZLw/
RknQVrWR5jVdtZ8nr4owhwKlv3iYJ2EFSFExfCzAVjlGqRQAwT7haJqTfVVx
mJ16aF9/q9EZjqeeScyr3xEB9NuXvck5A7vgNKNWZlTVzXxFNmS2JtkYqtku
4t592mOMMMA5HSSDIJMjYYWLzWv5hOk6qfgvraOqdNcv/bSPBtcE7bQr0/Bj
2aLkEL9qwcQpxESpksstWBQDqseRbgfRKmZ66HbTKDuVb9cGekw2OeCVnpp/
iqxOEyy2MwS8ImL3kJiTMYu2tNk394/CgixhTf/KG0LviLLCRdWBCvJX0JU6
BLjqxpwIdnqK1ZFrxrGFgYSpFN2Aoplz2/Ez/teyuxhcWU4AlItSJ208tDkb
CO4W7JIGtvOiveDY8gEXimG6MKu1g4hrFOq7tafjNQ4CNCMUtmssJoex2Qt3
9G9xrsaiRQo44CFqzF0OQgg1ojkVAJzr8r6Ws4JgmqfiQ9XEZgEDqKJFYBD1
f8zpOd1fkoQKCjAvKTaet6pICikD8nhuHwfN3bknnyrhD+sfpn2e2nRe+ez6
lZYPe9x44XAJEjpBOh88L/uhnaxaTq2XEgM6ainxRlT8isEodGSUSCGmieLK
mSOjEHVN9+PaEvNmpNvhamx8SVt+ssBLdCGW/dWkjOSLMaKdNQtk52G8L/MX
dO520EScgdr1pzClnfUNCEVe79XcHjYqS9ima9RCgZ+QS6RLWDBp8kxPMLNS
kgJ5m3Df0zDV71H4K2PTn2FWYRilTISyE1HOOamn2qmNdHOo5MFfhcXqnYte
9zbWmPWri7vWboleUaAAi+uZRCbcJLYksp23CzpNEVqtw8bSYN/G6O5L0Q4K
MUTsdqM2ymmTiMJirUmTleb6G5nf+xx5OT8vweT0TU8QzCOrgkVd65SHXm49
pSZ2D0GfNuMSCfmxD4w6EbO/2naH5epzVWJRLRPdC6tqVhJV7jhOG9++pgX9
rZW6RdFPwQRpJxaLsUTWGwXiLsJmVyhZlXT21p2wLUY5uqnrkoyU13Av+Rc5
46g/XM7PFckIgH8kS/yVMfuwW9rmG49hXKvmXgzIuWHcoLQimv23hLH7VMHe
hoMHm9d9jiL9QLG2CwF5tXKya6BnZgvUw5V9U/P277a08jFFFPKuu1JszdpV
W2+YP8sZgkcpx41SMTGGrIfJcGE9bJhzd/KxLl9hVpTNtC1CQ7MKYduM9J6D
3rRraN8BZ2/3lT8d9Ds66kFhgI96EWO0uPLnXOXQBvDE4eOyS6hBWeTL4BK2
CmfMoJRgFx38/cN7sMIdvlzhKLcGMd2sB6CyWfELzHvPK2wOuK1O4Bkvilz6
JVQMUs/OI+1zv2Z4qn40YmBy6xiLpRETR2brGwaEZBDeONywrTgbUW3bSDnw
/l2e8qhxW/xccBJAuGy2GThx3d47A2hhBSGijhKpUIgc2i/zaJmHBS6iHwQR
9lHEI35C6Y6x7olS4pwZLvM9TYhWUr7L8PFrLXqMJ6fAwU+brT76zjP4rO8o
87VIeyDLPzL/BPlD7AYTMizo9d/GCDdcKoyslmNW1vmYjEto1uBMCnfaszy5
EFiL1kjmFKBnoXEmEZezZHpHDciVF3vTVHv5LHycrRFz9U26n8/nYVKTRhrS
6R2h8zjsK6Ckbk8BSZuL+o8KcaPuB1q6QRKuVAFvqUgatoI3DvV3fGARubhP
B3stgFeMMNxCqURzvfvEnTEVqRp8Y/j9ug1nV8QPE0mfjsAxZvBOPI0fkQxB
1+cBlzNwSehqH9weTSrAgj5fRqlKM8NxNancFaLkKYCKYLpOcuePElfvXpiF
8XCB+dvHR+96Hbr4zgAAG7eOoxd5H5hljKrnjn0afwr0bLFs1qYUEPUgaV50
18tCCV4OnF2TAX+UBc87e9MwDG+kpL49f4zxQtNrAwsu0chcbCzt+IZuqOPs
+L59PEIxg2nqNzsESiXWvP5Co90/cOFrpsR1M3ZXFFUpKVdXbKAi9UkTI30R
hxg0DcLWAPGFUqarSHyD5JBOn4uAMyPN4yHRP7ZkIaP3XBnWggA8Eajb30eg
crKtmFDRV84oCx7jfsT3M4JxxgdJo/wUO3PmIDD+snZqtDFYXsH0eIoOrCKw
721Wrk7IkpPd/ACzuxQ8s7kzpNQKbz/9cdS0qosyqSahTRG4W7+cmO5fRdMb
Sk1llHqmEWmm83nk7INyELX43pV76sCVi7IG32iulnSk7zwcM7VHpE/oYtgj
5mmgS1AG1l3NDpkDjqweVXvOclpxFPMEEfgiPRG6ox4QOw3itSD8mIuO3BGp
FVwRLGCo16S4qM9pWCmh990wiEHhcgLKjQcZA5U/7HRIZEbT7FkP5TE6femJ
VZyoCwwGzpsQM6mbx2mF8TkfdqDkx5yai+2PUT9rJM/ARtVHKwdLlfteEEEx
0Loie9f2DuminToQdOy7fLVAXbaaZMoOAGW5f5yV8AF0l7N7jEXqNPGcCTnU
hlZsimKQkS2HWV3CBZ3/76g44IWxQb9RL0lE48d7cDWwVtJlhbSVHEZyVumA
bHAZPSnX7Q/vWPusLIZf22Dn7lFuYE8uONrMy2MR+XFg+ezPxOSWc1FmoohL
Kx983p8vD1Oarize9s2dNz2Tl5vLUJbhmg9miBsXoIZDGI71S6xD4LqZpHdo
3VY6jIkIecI82pzlXcmhA9fMe+NtlWTnAPOecFELWIMUrxG3QYuDiTFSP6VF
Tf8WsK2yEfuZLgRjpJmjKfqWYtmqH8l2aEzlG4k6mCbSCa/Z1pSlraetchyR
yPCU3Zf9xbPXP2vPhI5T6yeKgTGESz1v+r88pbx8OotewHAmXNOHe8SrDYu+
9kYhisH2r8c4Jtet7YvoWRToA5xD1VPiK47emydtZVDxapD76/CENbTxWIpD
KgxqgPD5wpZLT4ZsdB67yS/x1o+pZNH9YamQHjMPQpfqtc/HzvY7+A/kD9t4
UBRJKeggoITjxpnz3WPrbRKnyUco5tG4mRTYXe2hz8ODzVs8zhMuW6+BUUfh
UsqsIREFCfTImSSh9ub6RbOuuSu50oT0xg9eUEPHzIj6o9TTw8buyWDPphUJ
7rHw28DODEf85QL00cxCrGpLsdOsbmOh4qBpafBcSwyXfbBRwwEx3v93B2dK
YAeS1zU0Ah35/uTCHKq7zz3+B7MeZfOtGZkwXSPZFGHmQ13YldJ4iRrKygij
H3XIwtiszzYnhMKRBIWQejVmDbObZC9CgSMnU7DoJGP7EG7a1mhgzeFKNGn1
KdZdGoRjapTfsmToFZQqxyI/ZzVJSua9SdsgY2LCHi4UqZ/b3dU8Y/zr0fN3
U1ygu7Li+lW8Pw9KfvcBG0p5SKDBrGUNIt4zTEggdQkhtb3s4+sXQ4Sa3OQK
DkbBS7eUCBdC16kn7JJo6hy5p4FN7Wt095hk4IGSC4H9nEX7waxsaGqWBL6b
oI5EAI75AOLyAzP2URSm87eJkKgrx1B90meocl9HcApWYPMI0Oxj3Ld6EB5U
JprxlOUxAt3sm/c3eZ1xKxJg30QfnOFx2SykCD6Qocoa/k5MJJ8g2M4JlWlx
VWjOUUAU+Xvd2PMXUhwJRz+TunjM7wIawEdeVCvR34HCfotZrr5k4pxYYumw
rxx74Nq9niFFilMC1A1Mvnpt9afcUrhPe2x0xBEOeBvRG+pcFpxWWlj06QZj
k7MGAmPzNuBSaBIXOM3zYqVAzIp2F3sIdfQGlrLF4GGKG7hQ4fz7gVKg6oCL
7nL2EI1DKqu0WMx2KLdMNHKktp2C3fT+VIfjhnE8cRKsTw7VmjFi3sLxkqqc
nkI2h3fCtkO53+vUWGwpe6maBkSFc6fhDJ7Ay3B1iF5Iges3dvTkQLJ+CMki
2d7w9kFqrl2v6t4HbTG/sfSfFILcEPZgxcKFFmAATrjUuumiIrkjQelbysMK
zy37oOjg/IYO6OShsdX1G9/Bcu6A5E3wTxXtCyao8u/3QZ1Ws6Fg/iBUnyyG
dvcPuuwdAD699aSQbqA76u8/jpOf0RrlESt3sRn4+9k47ljfTpwEOxB7fzM+
ogTz7Awx+2xyBzetv/JcXiY4+S9VjVbfbJ2mE58b8PhXauPzUrJ39H395Ww6
j0MqWbsKRoav4IN8/ssLT0GSnc4IvioCiBLeKpZVT1VtB5/m6xCJ7oTW3Rmq
zEwLUNgGw5u2DHe3RxAl/Xawi1jzxGo32fAGKZX9oTlZ6h4tUJMivgCXX+pB
C/OgGMOekCTGsKy9ojorq2ZEaqCH6sPyWswiPLYglWnEyXhGwyRnzbn+3vhp
oNkFltxKiKwQLUbxVXLQOSMJChTzz1hOTysCq6sUGrKiVUjmAO7fjSCnQ7Q+
cdjwfHkb/+GqvikNOBmCCIj3GueIX5DWjio6lBVrepFpXEKncWk5cpFInh5i
KeTkgIlbfmoIQku7/BhTlk4DyMlBSm2BhqVvCy2TYogCwTB/vEVrIqPSy/dp
O0xm0tmV9ZHc/CVWv4xdE7Je/l89CHPZb49zeDL+t0V0vkyeLYwLzB/kbZxT
pzboFuVmElLPqb+E9JWVTxeM5jL/YUReyNL/uZ0E/PhxRc3FSby0TkWJCEj9
mdfE2NLN0a7q3vAWSE3mdunetbwrr1/QGHsoknkEsyeCKO1bJ7QRmRcawijg
0V2pDsFxbNYwFoo7CLk8meYFqC32oUyAxEm/dF9Cz0alsJWg2a8hpy0MhhpT
0SVPMo9AQj9OxadwsuyinKt72Mg8GBpBMHoUY8rArtuBspuvjrAq5OZFHYRt
ZTdrqxWfShYoVcoG/6BC+Z8ErkwRVG31CsOPIf7ngyjLcf29n0NwSgQlTHhJ
c3/25YBSadhrNY9hMAFqy0q1ZdKWeV/xooOtNAc2X+GtLRJZpgWkSV5D+WR1
Lc1Rr7naPGiX5MNux5BFUGymL4t1fr7l98b5dEFly+Z4eEGv0zXJoL/C2tN5
ORIhMpD5GlfFkmjYqD/iYElTBowoRs+Gx09+yccQ5JrvmzJIPAc4+/Rl8plK
/Q91BtIvkgGs2wNj3MuRIr04AQcspCqRkaeldCErRdpy1GogmSW95Kgny+hL
eJUZ7xSjzk+Sn2apJm1LKi/TUAE4hvgEHNSldV61+0sSoasjldPIXdU7CvDO
wppB0mwdNM7ra3/24tQJ2h0sYhk2j/mMtLBlVAMh5lp5q5B8I6vWRzsVpJqr
/gd25E24WHJ+P9zOehXkmBqC6gNEoNvBv0GQNGVdNXyb2VNTNnz9gEXW4HwV
BR1VhnRbrtBBpu+O/E9vNB05RtXSsIYkMvUm0ad/8K6SGEDNTP89WoDvp/le
MPBvoYNx5RnTDTCWXgNq9IcJoyRnNNtDEmjUbmLDY8SocpUYSOsM1fRoJFAK
i7gsVA0tfUbWfCIIMY0mSU5papn3/cZgtStEgce1P91zJh6ofr2u539PP6US
3XK5QfgPY9KrU2MMUfv4N0fZfPPje393E9Wb3QXzMCxSN8zXPHQ7GmUArJl9
CdghjBNcVrj2CszpQKCWI817mp8t3AUHruR/5qAqGrhTKFY3bB3DXww26uoQ
7QBQ9P1w0Dxc+Ak35Cs8oPfCqR7IJ5J2joKMPn3kQePj8zeUSE2g9NgTmfSR
KW9DR23pLuGqCFziZrrtayZIK6X0hcrHDxwfwJXefJVuv79jyKGqpx8ogCvB
CrV5ZCAYufg5etfqrHEe3WotOTUAcg+o92pX1rtDfTEfneQSy294CuYnOzqW
JZ88n7TxTaYU2u0sm+gxe5GaZD5SLcMBNfX0hgl9xDaFpkCSv7oKFiD12MAd
OxrT4BxuRtN/EJ7hJRXN/jBLRQl1XU+P+toy11qt5L1u1/mQatJEdLxaadMK
5dIo813yXITbMNHDL2Nwb9/mnIy6kmSRxh7b7AFV9KwdfxxWrDCH7CWOFEEn
yjOmVnbUZk8Q7gdfkUDyAOfyn1nwtYxeUiGRFrRoi+/9OdRkIOrfUka4rpqi
BVUK0F5V8TH8fTULKPDuqg1RcxpGd+rugUP7lGZCeN9TqbV2jXjpEgwzUACZ
dQYstSdP3y7jp6HF9KP9j2IgWfiVMFyEP9gIaDepsm0/A6xJ0qdyBZX56jKd
8GI9OQ6B3UQyn+wbE457oP2a47vGyJhveEC7tiWgWoMcbtfAggJbCIRy9dfD
gedzJFrcxalrduq6f//8ONO48rjr8mwMMOCW2jURsHwvLePEe95wBbeXB2Ci
JJ01UNj1XRP8BD9aLo8OnKMG0n1vrWH2zQsWUlkktSI1regCKNijV05iaG5r
JJTrFLzQ69WJDVCNnL9aMA30txAnmL3ih0PtD+GQoUwbK6tVDqrXmXQtTOYE
yo/AyZL6Gkfnrj0HE97u+tgX3Ld52kf4+JXaaAQW5uJ/4hlh754Z8JAlPn+o
wUBjN6vQAZbn7Ayxr8kRaXnK0ZtXYSgU5sl4fNHHu9zbOAc4W0ES/xaO9vlY
c0kE4EPV3GGmyVIEPMaswFteQ0sfpTrBbMCNJHJBARR8iikgVUASWpBT673l
aN2c3sQ8vIhjD3GMw313Qi1tQfJscI07F8lBayycucC3DPfVtGoNDAxu4Pfk
Ty65ijyrB89B1Xb7P4h0WYI03HY9GwXmksOvoHetBXfuVb6kkrNhhROaEF4i
jxe6H2jOmWDR7UJ+QH0Pear/EqAzw8qrGTJCYq7o5xe9X5+O0+Ds1HYObzLK
FhuWqrKqtomjtTYH0hh6EKQn9yODOqN8GrEqHfpgb/I90eHyuU1DUQzfrBZ3
j8Pxou9uWcd+PmLAzNGgbII1J6fIxKpnSYu7kzUxuTD+I/XLVzh9Df8lGavU
MojUQFuRMIuEetEdYbUyvPA2CG1r6W57yOAuEHwp5NA8rXhvix0wArLg+rua
4CNdMJwz0y/STUv2BR4+l9hGE91NAeXYzYMp6ptu1vpG4lCiJV/g+SVFrb8z
DYAGSghs5xAGdyUDsIqGuG6msG0/CpMG+6xTLhGFqOw6Qucxp9F3FDsXxSOW
bszEBwTO86R0bSZpi/4UInQ97Pqa9OwSC0t/4/wVv4OX4YkVDLKCOYJwXV6D
VpD4uZ3vuVMisSWaH0+/Le9KF971Ykzx2kYG/ffzhoV0rWT/8uf7i3R6+5Au
8Nh9khd6Toh9czN8fiQIvSJOX2vlBDotLJXDTN221LV+8aX7HtLPAuzobMT2
DfPeD/Dihhk4quJvGJYvFOTZllEfvKkGMHwb2a/TrbhqBPVguIgJrtz8rkDD
ZOztYWZuOmD/IrjxADmOpzk8PfYQsv5fpi5U2aS34xTDONfMVzckYjcE0dnS
91QAyPyfqaYBxjRhuP2zPWgXlS6/WxyMG93bqfMd9yK9AG3Z1B3jfS3z9ow6
bwnrYilzorWQBZiYcBPbtIJuBA57A8we4hfWcbIq3iZgbmcSxKFDkqogSRin
5lkZKV/cbcbrk3g3SSypIexPMfBaluXGmS/0oFWxOIZdkfsgx7TDajw6UC30
Em1PeysjKhyVYP3TtSx/t/fCd2iiho5wB76653+LNy6xuMOV+0dSEB3LIFXt
C2ZQQeB1VeO2fBdNtQD2co1X36PcTky+wpN4vxczqFbKxb90TIRHRVhgAi90
OTj6YcAaPdZv8GidFJ/HyEQ7cVxMg+f6LrHIKHzME0Uhafc7VpqURqjrlUEI
5PzDaUu3/Fz5qZkVPbYiNWKnTSRsuFEfChFKssCrOmAiBowvvelO/pFnYPLa
klHfdkn0sjIbFcpTqNhiE1FejkFTLDH9H5bZ8GnAYeZpDEUorgz2WUkPaUb7
avEfTJMtCSuaKm+fRxfvlOn4twLYED84qnv+Y0XKiB1m0eQI0tRL51pfszsA
/8nrFshfPYZl2nByGod9K5cT6WYTTj147+Ay7zIfVj9XXv5zKgpAHLDepg9K
LOihDC88UlNBcWfVRy5Cqr80x610erWNHn1R9hlIMk3z5WQY9/LmKU/hDGst
bq26SwJweyJYEjtBewsomTjqY6DDnYrFm8sQseAMOt6tpiK7iQazA/IDcSBy
xB3ZhkEWKO2WiiHQZkS8zZfSUR0TmGchVSd9B5OtLH70qgX+EQQ0pvtLdcvR
djiYnLQ1W87yz7rYseXUtCw474tGt3+Se79QPr/VlbbIvvZuIA+z0ynIwyaW
MPaKAW+5m7XrGMAfTOFtY10I/sX/S1UdPgZDZqa8wyF0eD2vqkfT/tYjnP7L
Q5qa9+bQSmZ6H7dcLsztN7wlGnzGJ5XeJfF80hs54VSXFLjP0exCplz0dmm7
AHH++C9uOfKmvayfzo1SivkNkfJfftR0nY0YTk5HGISeI5LHmqiKeOtQ4qhi
lpLDWwEUGb79lU5oPO5UdWBYFP7dTZx10bkAhBV01Jh1xvgUTT3/eA9NyupN
parDcaK7L6gm87Ja0ZJrfykScoeA2udi+674H+RDTTk5iNQ8KYwvjsZ96RUw
yV2O6N4uRsrS7F/X1aNtMkZa1cBGWNq2dH0vpxl06vSwZ5Ohh+9JW9/6HpxW
FSozZv7084tbgWgFSwv4/3MtitKpqxaTVNrJ1LOao9ob6ejzG+Jbt0HNWeuB
fXCKtihZbMDL2AkK/DZRNg5Eb7qYVmZguZ0FXsqhVvzLLfxkATBG4dRrIMt1
Bm4ySa8oKbJUZIpyHuaFnXGevGG+sadwiGDk8cdqbbCE0fzdiQ6RjmpwCyxm
11mn5Ti/vaNAIe4wvUE88ksZeJs3bUsy9GFYJDqpUqMH6apPHYqx4coMCHz0
ssOW2HKqgvAoKwNb3pUxxRbhtNNq56TDwQhmOc6wsPZsJpelCJ87XgoZK8Tl
vAqz6oGd02Ogw7FFeZ6YmAc4La8ihe26/2uIsrrX0ti6n2NoNPOIdtylfpF8
RCfWIkO2xw+UrGYu8Q30bWnMqV2gjZCtG5rU6ab08lSKoRuk/v0rKwyEkY69
GuEgIrMh9RGnKU+lxhUzDyzRLXoQAzwc+V4VmOc1k9Tiy5ikGXNMV26+dEPv
5CM0P04WbFCTvfGeFoEnhKSIJ+pUUKH6jVcmoWoU00c99YvsWdFLn2RVNAIZ
k1JCOKVFnNXall7Dx5jtrGCIfPBTx69MMgrAa1iJko6QSdLIwDfk/Ja5j1un
I69H+9fw6ffIJVr0LmvODYRlwbbfd+wuszXInm3LVnqypjiqdQ3kl4poXRsM
ORvtkxu0xfrWd3czc2g+Phg7P6LtKlXwLh4WaxDQRKAnVXZhy4sQBsVnegFd
Z7BJvF3tJj+BhFUKhMEIer34cn91PYOB6Zf47Dx8W/YznZTKQFIPObbg8Qgy
/bZR7GQuYt3JZU0kz5oMfSDEoSuHaSN9vkSaOpKplt4Ng0JrWGMjsYZ41Jzr
tkv91z4cactEo+XkKiYNzx3mCqgmACG7slTkun46odbR8NAzeoexrWeFZ6TI
gnPv58cACc+wmP9KXo+QyHzmQL8KyS7+EzGtDlQzyZtwvtFQsxlUrc/Y/9hY
Hi/7PC+693SrJbj5CmV6N8h12F4p5o9iuQ0h/Hm0KJ5idFLT3h/atHigBVOX
sZaIxB08YnIQxem2NnODwg4buRcKbkD+M1skwCqh/+0rAHPdy9g4Rp3VTIvz
kpxvAFRoKkFEUNEKqryg2PRJdY9o80tk4m/XyYtgYattKw37PX4wSrcsmvQr
sKbAED2VUyojS96O10d0iOafxND7zrvhhSGYb8nrNth9UrlXokEYzA4VgYwQ
YhzNPcUsKU30k69Ci/HFh0WZJ/xREXz1rvqgyvww5wscwa6nVz7m+N3PKItG
1EA/CzyfItpSJ5lrW9zo7Q2f1XlgdxUnn8az02FRuJOyYWZyQBM0RYxNh/pz
Pyn/QXSY9r4kL5T071BImbfMQCPwb7laJPmHcvAGdsiLqTyXTRvqPTICUguc
QFRTPVch0y1J7feAREtmci2IFD34H6PWDyncgHKwd8FMwmkmm4tJigAOqYIS
+goofuf9sAiJi3Be3Rx1Kxe0wYRzF9l8bdvcfsB7SAs7Pt5AG7zLnYpOpk5/
7zo4DUYtnynW/5PpG+K/toggoYkXlzyCTQ/hWYlzIzVY3vccHlTqqkGmMa0l
qr+YMG1CNqsIQcNpO6XAleRPfUgwUO6qMRCNk3TpX7ktiAlxhPCUzuVQaD7j
a0kaxAA9RG+vQ1fSgKMMJ60C/qDy11iEWBanx00NrwAHhH/MOSe+VpxAdk4z
S1RJrp9cbzMSVKoZ/Ap4rdl1dfLaN7r5W5blyN/oijybqJ/hrQp7MuwRF+Do
97j8q+cHZlfnL1dwgwNOiX//oBBN+OhZVD/2U78VHilXNRnKxnzs6Md1pmzZ
FphRkHnTBUOITviDKgcH0bNzojz4JXVBuTcItqIt1n6Lbiy+ySolNetTiGlA
slK+f6J1nSaeueJn4+86X+wyqdHCIL2/UdYrEZQqb+6b/Dqbhcc9QU0Z4Kqd
0ajzBeEyO1ZSiwdLVeHbeNChp9xlSVI5U3FgMc18ydxsUs2VqgSReAhPu3R8
FyzwcoM2nWUuSeb/wzDw7gLNLhbfHTeiLd5U67HLqyfHUU7NIPeSVZDuGWHt
u15iDxA4iVjkWiCDGwdoTTxi6ONHw/kwBxADpR3540utERCSFZNET/3k8R/+
4Iy6HP0VskR5qSLjaR/bIYvG1PeeJV7KYX/6n7+AJ2J2J3ZXxClC9MbOCHPS
N3rsitJDPqpNcrxFb5VeczuLXPCNxfHk4D/+9gcaaIHUA2QMArbla7+ZXv7T
LYyOb5qbgjTaOl1zsIWJKMoyEqq2c1CoWpFiAVe9bw6RKBkYqVn5JLmahk6J
qNCXgZCP5M5LXTt3XhVvQHL7JQfEZEFBKtLe0X374K7uZCXcjtpvubQ/V+Ny
q+KXWvc7I/1KhE2d7y6RE1JPSrk0t89jvGho8R8QrfH5HP/a5Aeht2PKMABc
uQjWt6SCyp3/n7rnfj0kq0I2LQv7/PKDs/yy9f95ikrQenS/kiGUueiT0DW4
vU9XQOSwfK+KtDIcwBs60r+BP4fwclftVuedH+vEty7rcwaxzEZCsY39zNnY
KWagUB/PAqxQGSavpjtmnXTy+FUJmiT0nPY14qzcIT8yskVVX8AxMu85z2tw
AG2+OjfFsJvDJWVydLM3PtGStW/pudGwJujJxOUvGnfRukjoPqElVoaaMykB
7nynnetyWggbTZIRLWC+c8f0nQkchJaAvWg9wWtuOS/BIV1LmK+QqHsHhegS
2H4IbMIi3pAZwquwbyISxzalNshNGeIknwGy9ZknMq7SyYoQQrPSWrkbGwOE
NCjoJXpf4d509hnkmOx7uiAIFc1dhHRTcTYBJ78e8okM9fKcd65Cw448aw84
+3fypnfVypUBi7rzPWqNtttUVE1X2e5r/QReGSbORWCEr5wpCno2i47mMA9U
t1hWNx4DupP2/KTNx7sUVgH0pEaIL1W0a7v1Hh4rYAir2HaO+Of5P7YP/iZK
azyTsOhOVZILdPrk6lKtmrUxwH+osJi5zyNewerPoKrNAhBo9Pi+MuE+eEHj
t9gVbTR/9ejuWPT2R1FtxjHloKpULfDTqG0a7+wPvG9SgsAYU0ZU/OK8ILQ4
EG1s5LxV+wB9VLEqfkiEOUUUtngNZ53znj+uUtMSLdQH6N6Mubd4JBnBBrW6
o+I6IAnrGXZ/pvGIfnJdGZSUKwTqgDkaTZK7L04PgslzPzPKsOMiIwr0ms2i
meGGAkau8syFXkpnTJHFyIMtbBJdDP5cNupzfu9+jVLY/IItXZQw1dmtt0Ux
OcEdR8ht50tixy3KPfbQedCrje2/fUbXGjpuFmKjlVNku2nCmPwVIR+iR7yY
acsbvBRRSX+qdbgHSWe/DDVVeu/v4SV5krzp9nLKZ7dXAFN2FQSh1WPyxbP6
RzQJuuVeU3KhTCYfRE3B+8bjmzToPm8jtDMPwJkuBka237f19yAGuxkm/5CH
ioJBnSdWJ9Yg8C//2J5F1ODsuCo5jJnLjDXJGWiWLDYp7y3p0+R+/0KIge4J
X7kIrqx3bY8eRQHmyLZwpkUirtjw5VSFxEpp8gW54zB0dXRAQYrXXb62Znev
lNBOQnM9Do4Nugp/B40IDf0TviIql/76CSt7/p8hm7Anm8/DtM0R9MQV4ZB7
k5srjs9wvAQSEgRSQ2kxdVLCh1CvOKrgR+xbd5ugB9SWTL2UJxbrD20xyEaB
sQcIyXtcIStzroHRfBGdjKKFuU41v1fd3EwdhKwK9dIcE89yM7VH4WJiqcxa
wN9+HMeiZDPOH5YQBmfXkVksT+JgUFgRXtzIFUgzGDu75cbaKRGlqqjEhLzS
t35tUNQfpcCJSUD27BSTT246wMyyEZ6icZGOJNioW3d9Y0g2BtRnLFSoifMQ
gMsx+0rrOmIQaSKvtS+TJ+4MmGVIGBnO3QzvdvU/8FhELCdSpE0PeFJeKKtZ
GL0rtcvX6myXgBmnGdvmb8D7L/9243T/IKUCkXnsIoKjgvWCEf8rb8zvj3hV
CJxmvQ5Neh17EQlZaDI2gaan5Cr5LnJbSlzEeyMcgM6RhsEk3DJ2B7Z6eK91
CtxrdU2Nb/O2V90JnocMlte9YyqWV0ZnYVB4E+OWH+Wwx0B6N5fBGkHk5CUl
oX/uK03ly8NXMzKHI2aL+9j5voaLmdL/cBPTPrPTWrv1Pn/O0me55AaytxGL
mrZsA3jIiwShOaktz6v40PMa2EHFF2INQ1xOnKBEe2CqcjSbpOC0mj50UdGR
maX3hWf/TfFhI/WYwyqJlt9wE+czqja+Cov0jN6hTuccQoXXX3Uo9l0OQCk0
2AzCiVH0FKfe6KEmyOXOQFm/zR4QkaInYGn+um6bKgtwD1kcAvSCd3vCMULa
ckYJNf27qycSaH9Rc10b3GIXSxSgQSNb8fNYCJ5sKf8POBhL+QcGXCYYn1r/
A5QvbaxPv3YdcjwyOH2Cn4KPio/0ZZMMEu01ZhIVXmdmLd6mtPLdCFhxwp/0
9AHZmMasRS9p6VcckMYJb7J1TZN6ZJILSP3peHMuuCz8toAomYqUnpJflsg9
gtj7xV+RJgwBEJi9fM6zadAXHd6ZG1o0igodvxNfJWhifKhBeibZkNKkScVg
o/lyBzU2+/7kmqiBiKEdDqzbNJMkiYUPiH/ZnhEHVl7vz7PVXIZvrFU7niQE
MbM7tegAFGtHB8j39Xr2VeInGu0ieKLDJnYOLl7bnZfqU2pIth1MKsNk2Olg
3jhBb3AP7uNdhvyrJv0h58Ki3COyE+PSLGe+tn1IDvisRiRdCRoVARDuo0z/
5qW18uUv6Y4sMviignnLFWjOshp9Fm+2PZX2ZZdqSJOViR5LcyduYX8/bFbV
KfW5hOYmRMkuR38mZColDrvpO/xD3sReJLtoyfSAWpq98VY0M5ZdBUS7ZYG+
StTEHnVneigMIVMAxkimkMLEUA/fEgxr3zhelvQpYcOoJ9LV1hrzq+1o+LLM
ASzuR3BuYTX/UOkQ+Wz7lozgShAtGNUatdZbYfAXZPYSYcW6PuBYfO3JRA5k
j47diX42cWw2tC1dhhivKAJYD17oT1UNUeQ8smx3bb1Kevx2ovwQWeJ6pN32
2BWHNXXE6aQkkiG0SyHt/djgqECXWohGMvMY030uus31x7up6KV+ftOmODo8
cgc/adDDa0KzLIr8/zb76ICU96xecNosBvnp2EfPvh0+gc9Y+jLwmuPZY9WS
cfp0FmqgF8q+7uQ0pDtJVAYpWzf/47TvIjXZkIHgWe7mMPPn8TS5BCb2p5jm
UONwOzeK9VaY8oarBnGzkNOwMxt3qStTGKCLaJbQRqHRr4dkEaW6ikSuEOIn
feDUWSAe+0WwxIp3/OhmRseJKSxDFOAHIoZlyXuF9vM6rLjXpspxPdf1keTO
4LRPqNCT3V4+Lku5fUOup76mCtWyBjvUi47Xy0YP3wF8NjZji56UT0lu0LwG
uWtc4JBGHpzYrB5uDPG6fG5I/TeOOag6iUCOjeR5/zktlK8U2rDQPFgYZxQh
uYVn20K89TmBAxLvh3bAKbPiTlR0r5E+OLrlsPAHkELrV1D4Gzw1Hd0ouYyI
OI1Qo/hdgnj8xBaiYxlQELWafFO18XBpYvBXuEjxHMxxh2xE75LCwxYmi9FJ
pc/8r27OZmiElOn01gMMyDrMAjofWGy0vPZctOH/zMfQglM50Vv+aj0hpioV
H65AZKZiH/Vp0FywXIrNJ0MsxnMXcfQkfJkwbnezgrSHR+7CAZXqdyZ6YzJ+
X6eZtRJzc7XWcQxRFiFNz5Huxw+2UIS5WKUWacxPdgfDpTuvzVvkjb9C0lZl
K+OlAn/V44A4zJ1iVJh4K7XxhZrQVqKhkjTXUw6BTpBUC8Nihnecv6ZiaaHp
jN+UDpIdyybmAQgPBgUf/gncWYZyyBl1DlellsC3GRLXFZypIuPEfeslXqak
fbf2Wec1dlKu6ulCxZFcag4ngH0xL+hw2JtCQBsUU7b2SnTU/qtg25CA7nTO
k+jHIkMhJNZNWSVIBkkD9GWXvR/mDbt3ipDS6OEsEPgMny5Qb8wt9x8qC9Ak
Kr7O0bG4jRTsvjF980/WnWJCEoN90/5sDIy6VNyaU+hPqsdVHfy6Gzhrs5W5
kL8R9bqf03mV2R8s8//G6bSAjZTOL8Hj5HyqNAopMVo7fU6Q2ljNCuCKRGEA
LU9bqF1rp2xBh8m5iwAsDWdt77jIsJVeq9YEDhbRK4ABI5R9sixYxk4KpVe6
QPMuODSecAEzfIuoBwMUimO1aUKcq+3CnejGk8uGXTXrcS7GZJQwY+cJpedh
H/jpgqHvEwQ0oSQK71vFcj5/QoCw8XIjvT18hTSQaHqZbH0iyuDI6SyHPYh5
LVIZ+bCTGgbFMN0/lCXvGUghU+R5U8ihwA+7H+9EpYfYhQmrCns+uYTx6jLB
IgP8ZpKHAcveQLb5Ex7ZbkEDNmNtMpOi/D0zD5K5Lq64SglZHVYtMsGFSIaP
Vi7cNj73sA5yW62zNC+V20fwrpGLUHj6Y5TCcQrL+m392kqSkuGXf3vWEzT5
EMvxZMAOWt4s/eNeOAZ6X6zUxFlh8Qt2S6yF89AvqMSUpC9GEoJaWpSeFPrq
UwLNvcZ+VWKiMkGm7FpX6ejqDcqbJobZA7CacC6c8bUUQ62WdKey6Btc/fSV
mueAy7TB/Bjwx7dq4PKpGnmFUwLEIb2LjiC/WJsG710Nr/9w9e1e4sFiYA9R
nLPsKXcw7+BeqRA0I5E/z9/xukfPn44kRtb095hnIxguKHm1bOfxnbtZ+L0i
0zKOJlePfnokm52Wz4MknGDEykHalk7anYjnP0H9ebLdfO24bWFc55n3yw2X
G/q8EFM0lYBN1dcADH/T+N2w2Wv4IoTgJ2lAipDoc3IRy2ohPOwZeVYGTd7V
9ez5lQcCWgpEgvW5biifv+qcWKkyVpqppxHDCK1BOt6F9JeDfgdeIid1bdDu
3W6YDhS231N3EnSWbHt81HbswKbXuxQGxHjGfnJlVra/jICwj0Nec8aphclz
FDG5d0opDGTw2Yj7qb/lfTYBniZHt8kpmrF9ZmXtaf1CvTdh61dH2xpta0tq
04ea+29HfZ5d0eJZ0NNr51FEb4Q0MHkTJ90dt6qTiMgjCOwERDTJm6YnIpln
AHkqh7RLm0YC7zFsIpA0DPXrLutFkajDhC9IcWo6sEuy56EdXGYEAuxaHa6K
bv/cdZ1hN9hrGuPhEKC3U3GJnckSnsCyinSSdWoB4iiVWjTdmdWYjoZ9wdTa
dZfSj7j+sp2HpzsxUebkYf2J7PSEGH+u7n2fp+MuyD7gi0CQTkGfKG0cJerZ
xZ1GE4lV6x/ZvJga7ScCW8u8OxZhb3guWt3okOUjgXKMmZDaphunVNh3p0ZH
ycelqhqX+cgiF95XnmXVv9U8Y/91d9nd9AqrRzEKU2Xm9jFzNsBHMR6s9qKO
WEzjRu6VpWX3q06POKBOrSmRRHiQ/9+R9KWv2lIS5vuW8nP6kBSgOQQ3XhpR
6Rez5F6j0ACtE2sGXZhPCpS2OKWm2cQMhgWThMHW6278sFh6HH44uhiBHN1g
/qiwA6erUogJwNrX6re/fAObdlFaykrybfy1Dr3IFI6rLmpuT76hxiIbisRY
+N11XkcAXeJKVGxbav89uaSz3E5+Ck3GRbZEf59psgYUznlytGH1PbqNR3yL
ScRXr8Crwxvb7eWZXYOpA2GRUAmP1M99CzLL68f8LUNhPu3j0Wzpm06fl/n9
7//ZDEoNRr/8X7nKc1jF25/ijEqvGazxJjGrUtDGoGXoRTjRy7pmhGNXM0rK
9foXbQaPGNssu3Ua4Hv7cv5eGLQnW6meBW5LFGlWlEueeXzQEB7yATpe2y2B
iLQK2JsAZc6LfCqLTYJVpdKldkNqnHXIO1SkEr8iCIRe8exsG5O9QyS6DHst
e0V/25urtlLR4/NkMqB00ngaBZc77Woz2eKzgd6U4DGwOkB+8IdSbTl54tYZ
fGxX6r4v+sY/6JLY8FdYHXwBT53OlQuw+fC7DAi2LBud0RZ6X4H5ETBp5sSy
BYi9qF3SZY90yvAypwhY3bIcJXGgOZlFhT6oYNX9EQU2bMMN7cjeUhQSQag5
F88xV+Hsoivvigjddb2zUBZ1n4U9AliHe7iB2kZH9gDdU6/fMoZBcdhz+8OC
QVxSelEltFkjOE9ttOaiKz+nn1X0KPE2TVse2dTBU8sO86TbU5YHjqmnmd4j
lNdtxBWwr+/qU2rKURWxcd9TNaFPIOgyFkasPDBiF4LhEp9+6j66E2okiENH
HGtQfQH62DbQ27xaC2s9LlDjdy+NznI/FQv7jCYZLpwGjfyDBGgG42l8Nro6
wWmMfkdidFOLLgNuVBt9drkeZnCmp0mQQfuEtitB5vuWWxRaApN1pObr6jjK
OpcYcADvTjWbcI/dRKEVUIal6QZzeOESvCvssIGeuCeWwXDhvZNFxEpbfYtv
ojPi+VoWxbqJ05Y40PTDFuUiuGtmCcyphILvfrQLAClRmBHgso/FAKmDX5sw
hOyGLDRoEr4vwgV3ND9BxzBQVQefoVhIC0krTUsF7/d+OT3Y4ZulI40bjLij
DbKFs8CKQAhhllTsxI9A+ltd4nnxIjMsf+JjNh9/R4E1QsnL9YMpgqZIWbUT
r5QCByWnjN0CQijJSapvFHuhRfuKmo69MgQbw/cPP54IOKvSpm9d9zD6WaY+
aG4Xks+c9MIoVHmw6aMriIRxYZ/LX3Y52LMQFiF4Ir8cRvejrLNlzsbaV3xc
BFd8f6uBiH0mhMT0PYCIy6F2McRZejCCGnV9uBO0BO3sd7iuEcZtk8ItAvDx
OZGNgjdiC31qefaMxaD2lqABJ8EITQr8k3SYlJOLUbbfAx8Ri3P6Qt07WT7f
MmWmExdTlf6DLrBLg6muLb4Q9erVBQeBHYffstAOw5Muzo/fc76GHPUP/pyJ
hdZGmTt0vtc7hz8KGt4E9qn8gO2/3oxjRiQ+9m5Wk6WbZH9ZIaubbiahlAUo
4nYWr7BXdXTalETS//FMn82FMeFtfNN3N8BRhztMNcCF9ybWRbX2dwLw5A1R
bL0UPD9H0F1/Q35mhYACAVVOVhdnA6UF3ey/4Z44n1YGim+X777AkzcgWVru
R4OIVpv0t1GiizfLmSy8Ej6aj3BvVB6X32D2GePHwsmPGZ/WkB7HicqG84Uo
E3VPjWSvBxOTFMjk/znHVIh+cHKEy91RJ7otpDYLuHlgr8+DqXh7G3784U86
1m6JMl3jnnUcmyfWqG+LdMp/rgbR/X2J1HsTF5bL94ZEHQGvuIzb94gCUl2p
vjlPXjrRdSAeQX8vhwFXrjzlmYOMHbx5QIx8qHLka2N/6+K1eyMaL4n3iuRN
hQXJ+fhU12peEgDhrNAcufgJbgvWEETlwZu5JRZdqowuFP/n1A5YnsSAtj3g
8tlK7ywEj3vBa8LMNYfWiHLdbnmuY9Rh5pTK/aC9PaeEljh9YtJl/u/xvulk
OPlghyBo2qpdcS5R+XxrLv7igF1kABL8i+CYmOByHvzoapVbFFXGOZPC4rF6
CWgxDmhzQkfvFDCMfp3YaaZ1h7B2ddg5Phu54XTKOiLxH7eZ3kk4DTiCyW/K
n0bOrGccRliAX5JTi2K2tcAM5Cf9WCCgJC2KB674efnn3AxMyFsiZXmcNtZx
ChjvtBPFLZm27h8XEv6j45CJQof7jhcsS64BDRtjfJ3k7xF/RnJIH29htOgK
hhV+GB5l2IkpwOYWSD+83DYtTquFEzE+4ahsw6mpp8+h4Ege01o1nR7Mmcts
w6vF17stVd4ry9z2j2Ffc2O0k8UYFrKxIMO86ctMpScb9N2Aq9QqTihn6U+7
n3wCr9JP6bm8WkoyUn2YE17RWRwUtxYpe5KxVDbk/WPFy662mOnykb70/6Su
1dp5vXuMN7ULfUIVkPiVhvyDaHvGb1PuXN4I+aeFSw90EAERIMUIpFI3h9tE
PXJ4gteoQcAsN1dLwI90z/1gLNTUD/wL752lexwD5VaeiXnixpn/KgVSD7sa
D12i21o1UkmKp6UNyjqqysZ/8vlB1KrQE3H95OdIPfttOKt4KSr1xVrvx17c
CM3bynYU1vZ+tug9kMJHwKRCKK26YlDRnhEaoVX4FVZsKh2vBcwVdAq4HHfo
YnLTUriGCKwZisyrAcOkXBpxhIMSoTEmCoqL1cYnq3XT2AeVlj+2MtUmCiAL
ylXZ07JQRfzjQ3Ra45Z8YWIYvyvGq+v0QUfAvwUiX3nzJdcPgO7IyAGD91uo
22Lrb56EHhfkkNIytfxlBIeAJhC2ZNsKJgug8EYTxuosMw9SotGlzcqtjguS
8331phdViBTa3st1r4Q7II5DkKI5Ae3aHwcB0vFQELyZFEmz6Ul2JIBUKX5r
hfP/F3jrn+p/DEtxAhsKPEqlpAOawzqffjI0KOptc6AD5rxOZuKiKFJyccDX
AMmhcVQEXI0q3KJDtw9p9HJURzjq6BmeYJlEa7XNY5+4mhNdZoH9F59+zg/b
fPH0QyWh9AwMNEZRyHCSOubJqKYGHwOehxzI97/p+hS9sT927d7CMmBvOySd
ucPBfN3QL5tnslN/UywLkU5EqR+PUdiTAvevRjS7ujqL3khsK1/m+3hTmgTP
1CA0Nm/DgKwaAdZe2Dxhbkn38bklfRbzH64uVGqKEu5WQa1pkTu7DlcP3ykk
S2mhrl+KkpEaZPxp/7ehN58v1osq0u+SYfsRp17BOGPdIFOOKx88S3jW7fu4
GedXXV2zanDjl3WP8yBWkqAP4E17n3imuAxatVYS929Z07Yns/VHchE4+QT4
IQ+yD42Ct8pZHFvdrM5Jy7xNhoab45cKRHmPNPfY3a7InOfRu/xK9is0O8lB
BpGi3f9XHh7/XAlgxTA3xtR4hc/so+OIjxfohnwOkdg6niTBwm4/ccKGMA2E
aeWYOObZgLJi63y80+K8Vm8bxdYJhmGiprzSaX5x0zhN2cUjlnJTDA5ASQh+
6PqiUIwSGjYODhMnuY9U+Unf0sUXfiLSkAAaTBmPr/3T7e8CkFYLCbITlHlZ
bm+DSGQ5svQC+8I7+4Rmu45zWlncnfwnkpp0hC7Q4FyQn63adTRrTvKxiH/E
5eemjDMvyZBdZcIW0O7DDriWjqiNUm9E9tgLykrCB+kot99kR1wTFvqj4vBT
P2hEmHMSAFleKvbqrVUEaDoTnSCbcincxd/mdZWNrUnMDi7Waes6foROyjHF
gzie8yJaxbzKOK4u5UNLNl6+IFKbYZxC714O4E6j4vOyEPiDiYU8DlOAaiIK
jsjDUUStbD5ZbcFblWcFwJ/AhD9lI/JQRXJybdeTy5Neb2iZ4TS/edlT7Rnf
LVX4CrKw4YY7IigPk9Zxy0uaUw2Vh7C6SD7bynzHQ0j2qpq7br/5V7phPtr9
5uUjDVZ6SWEMsbR7qHRMOd8YH5nBRAqpDLX7ZDqHntGVp6B09QdfmNqf5Cjz
/3r84AaT+U+rP/OnALChvwtjH6wQ9Dc9OVLBlj7tk0IS3PsQ1bbVylA61c5l
GsY5u3FsrysEtBkmtcnJD6lqGGRml80+e2sqkQfr+wdN4lTWEhWbwrS/vQcr
SQESr8PJ9SbtaC4Om96cDpt+pp/qtmbfnzEunw+g+n/s3OIbFE65uC86cSLh
vi2UUs8/7CO+ZWatZmhTuVdV3hbcO/ogAK6LRc225HfeSni9EJSny+UncWVi
VUvYF+o42L5cbVrQiigsyY4XY2KYPe52VHi164NXIH7+knR+CQMUj6I0x19Y
kzoUJt+yHPx/mRiwshBhfTfWEGiODScZ0PzoYu9zraq4xC5gQkEV8Ysgbg9I
8wuBgsRJWl+fn0bnmS/vT08u9qTmypPJ2ke3std/QqWvtZug1M6N/LtZuwRu
EcUihElEqqg0Ksh0A2GFlg68neGfHeiUdnMmwGG5qx58Iq/RS/7UpoPcoNrz
OwVCpt53iKmf9gY3lSl7Z0xf8mwvqhjtby5uQ9JcUfz4PQ+7BH6yNj8hcF9B
0j2+N3MuKuHefVn/66SDYvIlG4nRsLqoTZONZS2VHT9YcUNc3YhbSxdzaO2o
E0wu9KhiweohvVV5sU1PVKy3fVeQrAhRgYtnpgg6byvj/HLt8J7LIo1h+MLt
DJAebeHpWwYGYGI5diWRkfhkmrNF7A7kdyjKJXHAfb75K8TjIlwgqQM5DJAP
UyvcoSGmtjCvmIx1bBJ+GLQc5IQlUR0ktOa15+s/a77HibZVtfxeQY6y41VS
aKqGZQi+RvXxxtpkvTayxMUBIrGYJl2bGJ0zTKjmjKOdDNpKq8MDuTQESkDb
cPbAmojgD/XAj3InNtvEvd6aPsT5oz0pUTlDrQ+EwNJDY7Pw2PyIOfuFwbZf
zwCyzw4on9AR4eSz4BHr3pKp/zxU9DEBLEs4qg7NqWrWdT7J2CinPWFOjlIc
upNsqxx3SMAD1BLM62a8pEp8aRzpm8/6W55PfjT0s7FjvHsm4VVlqA4Shkzg
T5qbPBmJTiubuF78bHHiS7Q2ZK5pMKLXGo3a/oWq4RfFASYAbZ6xMQ9tspvL
DV0BIGkOoX6LG9CDbbMvJQ6Ci/tQESez+U1eNlwR2be68SSjoPOtihzweXiL
tZSRQEJKntLIYdDRqzk0Rg6OfP/VlPcCiZj+oo8JH3b6/iHmtUWAJG89joBP
ilpJbX2IYTyEyPzqUd2iMN3lU517S9p87qqqDEbGKjfMwWTmlOxdKchLgaIT
A5xsngCGB7wehOGDV9groMZyJHEXdK9zZLWvIhGB1CEB0kMmBPSYFv8HVPN1
VWHUPTwuWTRNFVifMmWe04xHfeE9XUzinCp7blqyvSXhG+M4nRL7TnxCr0w6
QuBfFkSL/ze5FZMX0Dfxnhf0JpOpgiXw7zRZut09oZqLNb6VYjUCTts8qazv
M0Sm9Vmuse4Ak7nnS2n1gfKFJTe9az1rQd7EtQz2000UGNSxnJv+BcmEvgqJ
DYFw2OS6u/6ODsTIlgtxXkttFMKK4X58HtEpg+WFhjI1xfjV1YG2Qz09cA1x
DMmju71VbLn1pQC30cqx0FEGTmJ+sV21ozCbxLMzKG5rQed66ziqcYraK0tG
lk1qpqETe3K3BAU7eTzwGr36xvbdrMeIBrVMwlpsJLk7ZVT3TApsLGB/NTF8
I22GY1hFSRp36qoXGU/2Xy9/9ddoSyPb+TYBBqkZy/KsYWn2ZfEsHdaAYIdB
t5nLDktxiwtSn3lsvJaLmw7sQrIGwXnR4dSbdEBG2bW+dL+BiETLDvKlbidc
K/9qqyPsBDqv90Oa/q2JcFBT8yArlXXOF7gANKSMoiMBH1pcmexqasPlFqKQ
lgSbeH/s3YD1nPkDiX676UZT87obSaFKcJCiMllxYx9ksOqE6a9wKho4ujZQ
tHOW8EqmCsZG8i7onLt1HvgIzABC4cLLIbQNToLcMBGx6Gr5IilKuUlgP8ug
N+NtYI5jXBeggWKoG9engAUJdcUiQ/veAk3/KoaTll1qbTkvdYmRj43+rKQA
Wl/Tcul3tEuvMwmxbEvS10VhrhAaEhYoAYRLJO3fgXKC94yJ2KAaegVztm5Z
99JxhfalTgkUQ2YxODulVszh1OQLzXP4rbdeYobyuGqhzEpt3rO556pLuN+g
Ur5QreW3jSKTQoU1xUTrOfbqmb8eSfQjeKQltsbWl35VGxBKkRUAHsEl+dy6
2iPCsNP6y4RjbSN5KovdNtY+KXI82yqSFNaMskwJVC340ijzUq4pKVNOswQ1
XTWZY+mkyO170J3h+HykzznkP2HaDvpq8bAmGNUqhwDQH5vi40h5WiJwlj92
+isLkslQ9geqaW0Nlot5pf9ki0eNnwQNzO5mlqN2a0rX1Hn+t+yijkFDP1CD
ewlnh6wMwZNpwFW9UYmFMN/OOKmQ/WB9VnwJGFSJKiBgmrE9WN6W58Y31h7l
F22nukKBb+8xWYoGwRmNp/XtdTQeaZVUr0oYxbF13RDtrhP5HCJ39htSJIXS
3D9ftWEbRsyHoAouWMldhDZ206jbp/A2Rehvf2ulexXwIAIMfwK8NipOfR+v
T9amc8lJH9zYAwoEXgq2k/nm8eKCEL1FTkmfxLQNB+cuZJlZ1Q07BRIpI0wX
ERnntkVUOqWqtt19i8Sy/DDbS8YAS/O1HojJe27FS2OwX/qGiFubAfaDPjeV
z9RRgUDPcu1Ju7ooWEg/lM/C+Oy4K0f5BtJFJuu0KU/waNTsAcRSlNt4G+ui
G/d+b8iFLJaXci/5zgcsnb+jboHr83PVRlJ1giF0/gFVX6Vog6/h63UvX/uy
01wy3IfmtUa0mcIW5CH5I2sJNvNnMe+vr4pNeu1Dv+Pjppx5YhMDrjazvOhm
kHIqy/Mr5WrbYGDRZzU22MbhximQ1kNWlOAjTw7Gov4PF4/GKCslKUbw3yev
+CC09/GN6xoGnZV/lZaMlusNdjov9aGsrFny0T9QqA8Jpf/1NlHZjG8Ksl8h
aO9dTYHqxdRjKOex3wzi8TTj//etv/VE8tiqgMzxBP+sSfa09lNL2c56frK8
XLDVkckIGlhbH7M1LrYG/rNEndNKmq94IO6Cqi7HNFbywAdkyPW+DjuyXOer
p+RYwdhT7GxSQ8rDgTAt6iLcRM+ESwK7ASkT7yIRp431n9jUtYlxAtG285IL
T7xxOW5ePFW4boqMl8cVQvU5E7ipbUhvUVX5wbhU7+XHuy8YWt80sSvjKpUd
YDWqbKSCI8cNQ5KAinLBUtG375rLsU9zs4WspxEJte1LR1cuD6CcAMVwTbi/
Xydn3dDGCzmYho90t4Xogtn7Fgz55s968BQGZNigPNYes4VjE7Mq771kIU8x
crX3QNxyKSrgF0ojOjT/6D8JGp+EV1wk/b/bWR3N+G0BP8d5sE/S52DblbVn
uvW2rxmlVrWHjtzeyG9afmSRPHNimZcAJzNArTxRsQOw9C2JZ0r1RZfRwfH6
Jorfj4JyE2ALOeStl58Kij/vngG1lnISZrd4kSgh2nZcGOGkgO5tJCMwb135
+se4nOhK2Os3YFWkOYdFbOKzi0rsJiqKg2gvgQCxUSp+USGACRFp7fUd87QS
NfsUUJ35WXj8oLsS7Cm4qecTrOL0Sk0JMgKh6ox9k3IcijJwmIr2+YSGUblF
u+EZieGZQ8jiiDz73vH3fEhqBpTW4TI3pTGUn4qCFY2jzaxSZI5S69zd6U6U
Ooy+z9wQomWmLx3N247QxXDIL/BspcqU9B3vQnrleVwfmrWpUMAJajYr0L0Z
dyn8Ehazejwn9isyDX5Rd8DP5MbUTg//USV0u/8ohxbwouvtR2pYqiDavlb5
ZL4qA6jh93A5P5joHZpibqKrVSyi0hNym/Oh8JZ3Svpbmb/+jOTnm2yj3AFE
G8mTd35k2y6/h+yDhI157xEjufieYLONym1b8OYoAgH7C1G8Hyd7dDQgb0/V
1jjm8Pmd1vdUBrWslF7m6gMAi33EnkSS1xuzPpWJKfg9Bs8HELxpHr19u4ME
AcnTRFwW2oJYFCZJ4bx7Sn58gIUs6ZDjURz/fRe4pAUgAzfgReA4nHSTB/do
NyKMjedYI1Il2gxkdGTcbJ1zWeAiMcq5TRw4OQDFbtH8bK+UR1kIVS2lPDf2
Rek/HBt2zhg4uI9OaYFKoaG9COVySjdjwz8xx5DhYnlv7oopGaS/3KKITywE
D7D3ddUd6Hx2E11MVR/GKDm2q1WDW6TC76tTWv5DdQ0183MLpDtqr1ftjJr5
44iiqZvNaVL5GQJiFEFBOLiwiarda6ruV77ZDD50enOxw2VIw0KGfcTC7Lob
2NGCzsL1xSH3lKZv6nSnshzoM2M3Dmky+vbKY9mf7qZgiEZAO+WdIs2FLfv6
GfQTw7hZxgMCt1iETLkLde+WGNT7q6rNJYzSYzwpxjMhMnjqSkoT/WlIIAmo
7uRQSdN9ZDrY0zE9gCmZmpgpnlJJiTaC5SZcE7qvXmcN1wMRuKE5Fapjie3N
8vEt9UAxiLjSmS5y+7eH0CFowMy5xgvMzw2M8H2zLHimnpFSXFyVx4ZjSUlf
n9QkAqIq0+usvPsbo/PsrNP6axB0PqVwAe8pgesHcw2YGePBWmiT7QujgwXd
VdinoF87Z52ZKcfRi5K5FaDe5tlFK5lCSvXUJedQQauEPEAkI7cV0/I7BkOA
ejbEreOOeTS5o10TteFhd0olng+JyInDnaFrj35gTX3Blplm8wRZQr2Ze/sH
NkyasvktWAka+KofS/zZrC1aQM8bRKUs75ANTcbhIlQdIS59nXVvoZklBuwI
dXIu/ekxnM17xX2K25EE24nVKdYVfs65RwxJa0EYP2Zhw7KxWgPMbUf9JyNv
vD6xU7AEnQcKpH1SXf8Pppzwn6/dqIdi5IDvGdDnVemnKWXUx3lhkyAyQbx6
CxWXTBue8f8W2sILJLaT7l+AfI8qQIZM09fH5oPitxBxgEMYuojvjOzz3lMt
cl4XvzORmN3NMvTSVSfF3LD8IDspglyE+uNN07Cebhl0fVWPx3mSwxSczvVC
Ry4cVkf30IIq81A/ztLkpOK6G6kq7FXTbXi7N+sLW3OqcU/r9D2s0AiN+Cm2
ltky28jOQf6l65i7a7FElcMFskzmvMWLGb0G5giSA9+VkfnAldoItf4pz4+E
9KfkjVTjqk0gPK7EAthzbIYreVtquYFTyECvJ7AYX1WkhYTZwYgq4hglIKb6
9NdVe6TJX/FunEkXrc5WXh3XwYY73MdJNBpEfj341WH9LbI+Er7OwtLuaL9n
dKy+g4N+H0g9G4GKXl6pzFQyUNnp9k5TvNUqkzkZS12CC7sPZsKjrc2DQUxc
LCNxEQsHhghoE8bb6Oh12GTDV2ewCawztyCH4Qjedbx2jHInDtgxKAgxSJjE
HiDn0y0GTac4djsM2G6EvtCUQADU39VUHetpKPChqB2DYyDqBeGUx0Pc1oKK
RH9PgV4DfxJJzpxz7a8hquKaLlmZo/AQMA9BRuRrP9R613VoMbl5PUOsIUsf
4GRJzRb6KlpMAA3DZ9dkQyKNiE8Ck8Qr0wnTOFyRP0wLp9xJpbjxtOyQ4FpK
3k4P90oCdySVwvpzWNjJhPEpbgZ7GEx+wSOn09rh+xaNK8AZz3FUkM/uOS4X
VSpGDIYSA2XVtyjP+K7+kFA1UUyIFRxkfPE/da5xT7qQbuxB8rH7gWJll/lh
BWhZqy9wkwBGcW0/CMj5oUXNywNjn4P7m03hxcp6A6mLP0SHwaQPJwb05ZSw
/uvC7nMrzU7BuQqz62To9c4ZM8s6H+qWvV1rnzdnTnMctonefJcuw40iOHVm
ee6GUSiaBZXUzXq4/EJWDefSqaON9QL2viSxncYzUzEgqUGTYcC4SpVgAanX
E8/TXp2YZukY0chRIvuNrY9H/yINCTW3rj1wTytEXNJoU0zf7EEZEnM6KhBv
KZ1erSjmPxeXvojEZFAq15K4Qrn47ZLtDtFsmYtwp6LiHn8obSn4HYG8trlo
qVMEvusNlF+rZFI7KOUB/ukeE8QdvMQiLbojcF76EQCpbBEyrx0poSv8Kx/a
j/mzcDCXPq3MyxhMO/8hsgwMP0mV9F7ehF/Ul5XAny3bGXmcU0lRXphMtTVq
g+nKTTpoX+dXUpUrGHM2J+S6Y2NNelxwEZje6yFFclIw08skMFFEG+DOK+7b
7W/hrt3WKUzGNKJaG3vvJMli8DJHGut4CTsFj6WsZNrwYHRxAvb6krH3ncGq
PDbm7xBSbrnMVdqrkm+WA8cVU+9ENXqGJGt4Sl6ePJv48ycCGYS6K0K8MNla
eZzKrVBOFcphH/q4wFQJep7vjjbu4w5W9O2GV0IhstEAbjYL5dolMI4QRFgS
/0T8exC44sZLq/poPtPYodTofv80BS0dfz8o+G0aIMG6bMDJTRdkMlmsXaUB
4yQMxdCHWG2kF9KMpdA9e8uMgjBrsjO7cpEEU/yym8163tYd8/KOAC7T/CK4
z3hPdyPM+66tywkSEBuK1vYChkba9wrj9nAgzXE2VNga+5EsHFbzfzTxtv/t
mBiWj0YHQsqwIyeL0bBAY1N607eKM8m7kfi5h4KyOZ2U598PDQc06dSBHp4t
FnMwP9fSnuhYFL6aroC9kg2Q3slOJmZwNV2neUxfKYaDw6GLA/hSduSjAe2n
0jP8kWEdMpivOn42MXyOm9C/y/A2c23R3fKJyvQdAKUBFtnzEiLguBdse5O5
6sL/XMonErEHDNEQQuVrjZBjkd7ykkgxL5ysA68GrxGzTaiCFk6Ef6OMq+Dk
CPZjnt9PCmFTTCNG+Mov3FPWbzsjAmdt4mDnkl2GZKiT443f9XTBXrF+Vr0v
1IBaP2wzafX8zObnBIYZoEEY05eQyE24qg58kA/TqrTf4/lxLKko8c0yhCBb
5IQhs0MpR2b/ZxQQ5RmDfb6vCegEhE71Ky6jNuJT55rZTXOd3+PyBW6kIXa1
fPvEKIUxQJcyzlRJA9A98ElT4o00rkjXBft0Hmfo4d4Iae0WFk//Tu9i6QQI
/Iifpt8JHvNnSFD/loTIxJfk8yfn7x3EZYX5KySoQd13kbg1pcPeoSwQks6/
NN3uFZHRuS+HRh9glRRd9UhRIkDYXwb6FqiU7BSyK3GkpcqE/8jNnvvO84mh
KYRzCocEmGxmWs2pYf/PNYC+BRC5owYJRAEUzsFKRZCtKAEMp40TRXMq/VOh
+ViwlwrVxLbdLToZ5zhVx3sk0uCTb9k72WM4mKW9y5yIwl2sSy0e15OZqIgA
moXjovAmyq2Ee4cF0rz5Fz1+1haoJX1IzTgSVpqrd7FT00Np9BfNNfVhRVzl
+43HZxDUQ0ElTpOIhgHB2A3EvofXddiEAgJf/zMZPoJ47V7Ouz5UA20y43nb
34ccK0ab+pJdqUnVv5mLD++3M7Myzs6WqKzJ3GdFDJ1X2tV6X8FLXpn0iwAO
qElmi0IiKbHTu/MXiNkW9DJcRAXd96KqAj6Kc71VrkOwwRc9WnwkyycUxBGc
7Uc6np5EOCfygqWps6oO9jSFqTL6qgpCbIEv9WZ9YZwuj3xbInOon3zlu28H
qXY2qS4hjDWeqQqsArd2HX60JlSFP/06QGpORGR9hZvIquWD1Dy0tgbUrypq
ckHSgUSt6TiKV5rXEbU1bdvsragzclewDT1WqQEJj6WC6GHnfWkpbL8nr5iG
jUBtfuQ1xmrCMSDQcgLbL+VUoSwL34C2oEfzvyZXkenO4FfV35klujPmw7Wx
7NJRkt8VGj1BB8FJmTRU39Uj7C/Xbq0tafgoWqYSLYTwBqSwyK7k18ArIlBG
24z7Vp/QFKoTcf5SzDugBx36hFRRo+4lr40j11RHeTcsT4qanxKqfyYg2em4
B7rgEwMprRrZmAJCklTYAcpITuazBqSXJGzGH3vzy7jGk01DHKNzIwueRNnt
WmPdSMyx4iZ4OkMxREYJtG71LWiffWiIGPHvmK7aoCEY4SZe4fF74t7ohiKX
7FP2ysny72m2mCwKZB5AWkIssQtTGNz6LPIiGF9kC0rlqrw0J67ouEtOEQFE
uH5OWmRR88KdjLTjk8jG2c7QjyCNxkyQs0143lnTrCsYPr8Hga5GvE6pR8c5
fakS9MSyzmgeoBWnv7ucqSb95co2H5IYGfCPTEC4RrEzB4O4VfJ6se/h6uIC
p7HR7BueF1x4iqrAu2Rp4P/4nDwQPKI4KVZTVIcqwQ8cgmuTL+LHY/rtirj3
14uyAl3o2quOaH82bhHFDKoA0rd5Xnlo/qcQcgeqq3yW3UaqnMPCDFGmQg6u
P7O9j70tDkUiWBY6pj90T1965LoII9T74BAnZ2AzRxpIeqsP6QdCIcFDJ0vr
5+YeCnB4eF9fd10cjtWA3hLd2Rcug2leQinGM8JRf443/lGA7Wa2y/8nEJ6j
0+yGWHWE6erm+vmo3LrH8ygMDCvOgXwKSgZ/ipZFMF3Tow51dcMhzD8vSKpb
XZgHUbGa4P7bbUDEfgzPSUGhC1lpMeyJt6wEHACVxSD/Uiu71F1TF+yY8/vU
0vkICd7xAnNxWyfNWyH/m2ozVoKziaVuSuI1XtNRlISnyNxPhfv1Gdt8uRQa
N6+48KYJi/8TXfDUHvsvOcyavOjImgaKNeOBql8BQBr7WqKzPTgL2U1mB0BR
f5LfdNQCghiHqPK2lmBV9dsn4rYT8imDA0XXMZxY3rCSJcNOjmdQ746HTmOY
SeaspFkzigT6OcSqdo2rstqJgWwvv/wcKhZt60Q2d9/CymaQmqJ6mGdhp3UB
CwCfPhbYwjBB1OfVx4YDLpKOix5sbMBRR+FD5w11deXn4URUcB2pI8o1SnFs
/PUY26AQYA8aBCbqUsSGBBvOZQy2ELgZ2J6l4GLrLHlVcMShIKqBPzM2t8cs
feQh71uG9lQfiY2yC8pzS9stmdYGDY+zixYS3znuxVkJ1bvX5LM4Ctj+CdTZ
URKw9YjPKjqN6HGIFnzszgeXp8gzZhRGIi0Y/pekpaqqn0Lw1rsqUeOQh91m
vkiLlj7wz67d4WI6Pkuqe/e5yxhDoU5BwoHabYUGyheHBHogJZUM9htRBTou
fJH5skWRqhDbbxcA0SLtNb8UJPML2Qng548+n7foWfkCzkq3gCSHaPOD2r17
zdgctrCQTS/EIwYx0sH4ZY7px0ZaYk1F/AIqaizC5XIK/IqAUFvVZf5LDyUY
ObjDZ7oFw1IiI1kszpFTcz99cY1YtaKpko3FTLrvELsx1Qjsbsk8U/0m4dPQ
GMjjNm8dpi6BiU4pQ8WGXF3RKxK/JoKoDGdENnJSMaV3PCd4px/F/mm+KVlV
uE9ou4JOtgjvy7pQ67Ae84tGlxO/36LVnb/qPncmtodl4hGz6caP+3mbEZQi
SlGgZLOOPUs+guSwUu+InGfx8uylJydFlCakSeBoBk46yfRunnSp7+4gcfX4
WAC+XixCZaMni9djJuPzFAkCYz3lD2ViCtRBYJEacyIC6a9oM33qfE++sJS0
cTY1cZLfh/fbCxlj3ZoNaUjW8XIxIkfYXUobnIeE824+IJTEMJYMXP+OLJ3C
ouboDufk349e7qRsM8ogtSwXTqs8sAVe5itK2ONcEFsGJdzJB4wGPly7pk3p
Cq9H6Qj50E6PpCSS2c6mwgyyCgBJva7WT+NRkHgjo6ZV+4sf3vlexkhtdxQ5
nXTg1heP+AxrLXdcXUV0udvLklFROHQPB/jN41qIzFvgYk+kPcKOOOCYg6K1
5TRdsZTX10nWV524XEQuWQF72RLoBuyhxYGL/IpV1eoZf/kjwWcyppsUSrNL
GrOtKONf5BkaSUo9B0r2rckODICFkCK35cK8pFbXD+TWdinrI4vs6jSC6WRn
E4QBSwTq9IH7C9+CwPcVzPJhhrXJEuPHSUBQU6faTIThtK6BSMFeJ+Hxe3qM
xAxLnznZBKvXZFOx0WPOXZTarpFFfo4y51vhsX7LrcTl0CUUocfMZYOns27z
obAhwCNu6kCzOvlASA4bzB2OvEViJLvVDXOJVLelFh5wbk2O4whRsMJe7xXH
7Ou2MTsVOgABgK8HzIs4vDtHcQPKRP+DXzjsVOU9AUr1WbBkqSmkHvNrxaKH
aLsArUUZK2Dqo8RKyBfyW+VsoUUrcoXNWN+xnoJtUxqUv9YTNMM130W8tU5M
RzEGi5Tp5SweTiqzE2BcZpz0xrBckZxcGHEk+ld3Enu6mF6T1YZZK+wABW8P
jPHhhZO/xUCwwtLBNWsZP2UbaU5l1aNdsOlv9DnkBcO6GSQ7t1hWVshpHxQV
VLw18CeRfUjsnxbYbo+O/REFAjtzJR9L3RzoWDuOBIgt/oY7TRp9ReEkV8Ii
4Q4DtylVzQBpUdi3BzmLpFGYjKnhuyloefO2NPRX+CvP5X1DftjBKDtMTn6P
EwvK3tvSXHCnfyeD7V7BMXTt3tg2DcvzrP1IBqQbCsLcvvdgmlxfxgDIESqA
qomgWZED0YkOeykVu4N3o0Nk8puLpZ+ev0qWq1jgqfskBTdMMQRycnTBNemH
xlDsovNxjX6xGwXsob2VEbpl+t8JbFGxDaNtAgz5s8/nlkA+S4x0rzfh3E4H
9L5oTnwUPa422B2PDstkxJ/02Gmhf9AfTe+r3j8oKd2oKEWApfGietrL8YNP
iOMS8GCMuCPMoSYz6sZcNv8F0uxWd1a5mTL5M8vs10ZQ6NAIsrlClsg1qLr+
jOgtE7a9WT5EWcjX6rYiATVtRbcmWmBIFJTH2JmvxiUquPBGyoc1Cg1S6oJz
eYjc4RZirH5+KwByIotD0iEvde1d8Lq5RPRHWKgfGfhKMnqHXuV3+NbACujd
XRLgIro96KEPUXe9sNV4DZQCQMJtj/AI+h7QD1dF92QeUQ1FJbJgeRMPgRRG
2++EVKtvvBSB1UJhNzR73qUG4zNbMvMOiMC2BZe928B5RmSzxZb1cOlZOEPx
/i3e1lhJMqkUjZM565fUqnHL5KkwWbQtJTOj9attUPpUsexbB5GsyWES48Dt
EX4RT37bhWdUqEpbyUZ1+b9yzl1IlLPj9z2pEcgm3ZCV9KQ0mVbxjIuRD/j6
52yoT8fxMsIMdWNflpYvdaVLA6fnkghbckelYbd77XVmdKYp9ErE4Gz5ElCH
q4u93yEiES57f5Qy3Yji1Q9mHdyOf+bsYxdwrj9Y6e1xtwa4OBxjMsfYcm8T
5J8I8/GG3dkzgXr/PqOofHiK8wEOkq1YkS68xlhBm2KPc1wwTd2TLY9QZ5iY
r+XBIW4/4oyv5KTFnW+0Hp3uVN6qMS/0VC6HcT3jyCKoWfvJG6H+v2zx0ep/
8aCVg54Xr+iL1xssWxDDV7iE/1RdJW/NXO8B3UxXVdhpVZumnDsm7m5+IZlU
8R2dMf2M8Cru2QD9azeiRus579/lg4R9xMu9LfPD/LRDwo2mdMY7tvHi/JBb
hxr369t8xnbH/OVa0zAIv3Xfiw9fTDwWAcmayNWHKGebsCU2v3YwL8oTrFfj
f8gkbxky99WGkLfi3ULze2ZgPK8EWPJ8Iw7FkQudeTKmbaVgSrjdhZpJ+wQP
5zqKKLLnLHv8az3giviA/WrEw4Zz5XXlpU/CVrkkCob5AfieaLBmiz4trc+j
DDO4UJF+Q8isl30ZavgMijyENtJMoJDDxmrNZDtDYFmfqQxVkro8GyeP+28/
OF76jJRnMlob1Sw6BsJdPR2LWiag1oGi6COzYcJ4Fs2p2BPOXhvNtABHb3EM
IXZFJTXNjIdNS//TR40OaLWmmwEYv0N+JtleJSOnHnugkSutsV4LgHuYpqr8
G8t9iXQVRepBKAK+hHtxXuxpaYeLhrIezJSUoCkJ8V5EY0NTxXS3wVk+tU8L
/Tx9rhGD5FcB/QLJ6nM5jJQn4fkLg/sWVpjgGoCAkSOcpy7h7nu3in9UqXGl
9rnaxRouSFgM9Io7fIc2eOsxz//X9TcC71GdVx874Q5rZzFbpTZdO6Ko5GjG
8DQXq2u3imvqeEp5llY5anX2xXlqNFTjtHW9z8wLMjDFQNhMnFX80LwqSDh3
KLxRBZOk89IKS4tx4uzX9wvYcsJySsQmfagSb5L2xLfTgWaR16kvKLNpJySb
sJmuJKl3EVRs+WBRiIYrFpgPtYmJA9gUjwZ4dlLhg5J+drvuYlr0STg4MzkL
cHjF6CUoNgy09AW+Q7Hz8RtcV59oqtnVZDaeU8jDrIfNS3+up7dH18GOQrnw
ThSCYhC+N/gRA7FYPudUH1Yk40FHI3Q0xbcTuYJ8uIwmymC5b1ER6mLD9DaI
3bDDyXR9fqXAr+BiULgf9MChOcQoUN9SiZjHx0ASPhv6ejIXNHSq/ulR8GSv
/fiVagVMDKgiycDXexYrAS6v72SjC5B+8c9ZJAvRdRsKNWd3eVVpx1X2qAoh
uP07emzLB0CTlYQ1eN86O0IJxIs7DXNNfXAzet9lqI+Uj2wFc+xoK3Nv9Mus
mwtC1aw+6lcvoBN1OeyO99EmKxqAvQ074jnO2Djp5S7FgpGqJCHmghQLxXpK
5T25R1884F8EC0/UPUFOvstJJFAQX4aDPiUJiRQJQjHbJsZBK/wjhfnSDu6C
HBVtVU1j9+a/qAf+HHDIb0HEjSk/F35iTKZ1y2Doe8wcIggI4mNmAkpfbRiq
c6dCFcWKRcxRG5UWDgEHurtghum3L7woTzofPaEOc8woo4Dnsq1BH83r97bT
if0WP0pm01aK2go41MkpynB0hT3wgJf1a7pSeNPFW/QqTUYvviYiXrolSg9u
N3tLALst/jUD7h8r+mpSFrC+1FJDo4qgIbBRG2RcQggJze6WJr+FewVMCIh0
5qaOV1dYpbASImcVcPqnJ8LVXfZuaazSaQBKabKgqr2CsI4gjC2Pj5FrTzj0
YWlvJezayjC60sCqzydbHYD2K2xOlXVR7LPFTH4OcxSrTAALlN0DCrfYtNfI
ZyPeeOEInDwycEGFaf11xjfIx0uEXU4yvIK2x2Wfwtn02n4tzaycH2JSeTwU
aD4lfa6+3mmbwkMFnxLdDA81Ri7YnMPmRIH5Y+L6+BGrtMeN+n2oD5u4tWfQ
gVfTvdw3zcrG3emNxRqM2cm24311OrjpEDkq/foXP9wnrOnQ5yKN9LGcjEbF
hXJW1WG+7k8OK0D36WuC8B8CcA753+/ewmp2JJBK4Kg+EvhPCk/jx2QmVRoy
wZQ6dG2Ew7iDh7OsQIqDlyp5lra+f0az15rweeUiEB3byNTOmnv/HUZXl3MG
Le+E/6gZBFfUmVsT3xioL/Z0u0a025wWf+zZ5twjq8xBw3W+fDtMWOw8j8rs
8UGBjfUV5bV/168rLr4NoxqBgfMh2b8Y4RkPTCQ8pQuv+un59S+qbQSWKpXX
VqgDCdF+gr7BS5kn2bUpOdQnpmhUdryVHVGe44OsuZxW3zUfLnot+DQBveWb
C48XOT4EP3f/t/PJ7BJY1aovxqvAJW8Z1jvhxVNMXQ/JuUJT0DvaJYmS7bS0
C81AstxdtnelSyXKW+A2V/QefDfNKzUFN//aZzS9fv+wnllQCwNTXgpAWgmH
A2KP7akwG1FF9Yh7u0CosnG9Yb2Jrce8bueWdI480wVR6gPyoKVrV+v+SIiv
iwuVuIcAcZWPrXlEzPY+5SYgLbdwaTzIKt/eB7fAak2NWr07GFOAs9y7SJZK
Pfm9Oh16jJ6PeCX+xRdqgxj4FKv+x/wX1M0T3KKlEmPkTzcbXQY7UcvqoIN9
bfWawBDP6axTeUh72zfmED2GvDhPax+umQEdBaZhJgUt/2wGn+Bg5mzGTkvi
HVMIXpTwbwx2u7hjrqcVXhMn1FLdkUbPIK4gIMTPi620pg1/WP0l5RzXEits
K5lLEwSgVJTefidrdAh2PYwXgSpp3A0c4JkC0ZHk8OjOWFoagXVqmqRmXn1z
g+CHhVsYJB1Bp+fkwaYeCRAIgaIwTNXc75btaQwX+ZOEDTSGzFPazl80PHWm
n5tnZKvJ5NBbGljrXphVOcC34nhG3xKpDaY8BfZ1pxQYB7bPcH8B+jSeZwhm
0BoFFM4yJ93JyPhILEPK0MQ/2r9fDucIxJon/hAR8qVx1BxbXTBXWINoXp12
oeVSrooHmPds07+JsAdqd/B/ZphlZBr2eRpNJpEsQFolFMTvU2NU+R3jbmIu
apZWexRM0atK7dp5DDbrA019UOEh7szK4g4c1k+qOc2SoSfh37OOpyhYdP5C
z075DoTbIgr3+e/B19HOxmuU+2Kivz62CgEpOB6NuEIMB05noRw9GxjZPa1c
HOk3d7+kFdUjDmPO7o4eZEoXJaIfBVFaGlRgs9O2msWEjX3zQrXCTzMEyMkq
hr/Bg41cAFKZG0T3KaLvEx4Tyrl5hxmKCnsH7HDlzlZrN6a8ld059Vh8L5yK
UFJN52eq2nkX3Fz/4lToHLvAr5GMp9SEG7fRWspGAxJkf1UgTgtDD6ilUUNt
nEXYyrQTcqbeSPqmmE2PxOgA1HbqM5qdujgnol4TNR4RZx7IIfHGnv/JDgTM
GxxDVslbwZt+K1YyWKb2KjPpJRyfYSjnfA2hATFKgMa8IN3DIvr1SQ9+ykp4
oeAjv0VmhNpTV+548SFvLLKkCM/EJghANKW5UVu+puhW+nK7nLlfybxn6z5L
vzaPpQ1aDrCsaftByB+KymVRy2bT4e3vGnFkG41CaBHE5W35LHkf1gxBge2l
E2SjBlY/EOi2lJIqCXvCExbZTJZQIEgfQpvl5KydEPgc6HBolHgqI+kzv6fY
+dxJKdtl282nnpJ3zOWhk6hXrLFPvwiOTUiNTnKJ28I3KcOoPbgtP7aE5L1O
nkzLPM0Rqr6ziXKIsvp52c5ohba/yj8nJ4toKTcoF2O7XINqIlEoYsQwdg2V
L7NVnHdybN6fNL2U0fU//yZP240PT1y1dw0NxihuSQmOJLSFZplYEcoAHK53
DnKy7CxlMSDSbfr7KzucokeUqiMx3zEWqlH4OaGnTATFSRl5Uwf96ifu3y4p
9us9O5566N8J/LACfnzSLo1GEdJFz5OEm0NEBgx5oZH/j9NIgE6ck/Nb8ekV
lbyKDkbIgbQ238UYf6/9dwnfvgtrNldtCKp2kvNrNuZvtHTmSrpvanZWc7EC
RPY1zmPskogmPMr4AbKte+4zj6SbH2ePSq2k+y0s6tJGw2HSlGrXOdtI17P7
PW3zSXa4/LOyiMHDdTI8eScpn4CtzrwUB/R791pw1PeUyptCaPkeCym8w1k3
kHMWbd8j+bIE9diseIQXoe/Y/VDnB+35YCytTBqXyN8mffro1o+iszhvD3MY
3KUTkeRf9eda5TTguIS8MQfwAYt1p0urn5TnpmtzTTAGA1vgPL0aIvkztwhb
nnBn9zSOnaaruEoQPRd3tfjOU5oYZ4d6AFE5Zjyyq6IeKgACms21yDmA/9xo
cMtuub/EYqyAenN7UESwz/TwFXucmiZKAhtTgB4Rj7fpChyRG9AdbkPgvH+1
178i4mNMMl5HLkyRGTEFEjlC9NXIlKv2ubEKmloljNcYx0+wuKZlSIIISn1K
aguquiAn+htkCiBz9xlWUdJv81CKOfO0yczS7SuZNd2+ziUdFoDTFDj6P2Kz
ZSdO7SdQl1RoRpY36f/DitjIh3uuNXDuedftNDgaTdOxSGWGtG4i8Vzl+Tyk
SWyTLptJrQluQ1UtL2YO3oDa+TaRMdnZCTSD9TTLIgjAe4sgXs4hR9/plm3d
i+ZEMUSzHUOJKC4T3efkk+3qP/6AkJje6DK0KUxfVzVqn7sPNU9D2ZFtYH/M
6D2FIAJzxlFF/4joGW15gcDniiQkFYD1cdIn23iQUHSe6fTZWoaXGQK8jaZZ
q4IJyt4eXzqL5uJQUHArmRQS3Cv4rUIyO3FsQTSxoVe6BGLL1r4JrIe4PLS7
0fK8BSihzv0suFJOQW+zMk920u+xWkTkf66oFvQeajH9dMJ+EClkOm8xxZf5
9opgcVN/gdW0P2+73/VO++VyBwVZCFq5EBNd1gVKK3tTARC5CTBNY6aXPdFQ
icejJ6zZJjjLmHcJEPKOsp3Q69mQK0oha0FHtkXbrQBVC4a0KTi+gCVZpEql
W2nxeSr4Bk+wtXGSgPTVTbMJRkoVviUz1hTvQ4VwB/ZqS7atzd+Sk03aWx6O
1DaNIY1tmaQmfN16QUk4BHi4kUHybSm52VloaeIuBvlcWSJCB5aqJ0QkulcE
Z9f1zH1p+fZRHQ7sDW6IdJ7Jqycq7Q5Oe7jvNGL3SYiRa6b/NhmsILCgBVAi
xRs7Da4A8k/T/0qRUxsCOYdWMg4RPK8eudU2wxLPLxVnn9RCZUYCh8e+Yqp3
PFbeEfNzdfi0/w0N5IyjKCgnOeiL3+PWBjhDBXyYyaYl8yFESrm68DXNRrJe
bJdIop8yHs8K9blHGxZn8szKoFtBSEhCodd2KVEo/1/XHpCGEAam/cLUCLv0
ZcM7BMcxRjXsFyOyuyO9xopwLWf4DF4hPsFPALOIM4GObNUxirNR5YT2tTSq
ojJ7Aj/305ZOX+flblbgj9oOR6j4V4GTfJ4JCzuIyK3MsBGzDkiRXDeDtSKT
pWdT6YzdV3Up2TuzNzhyQm/ixu6EpTjoKq2dQfYcZRg8IH5XY8r6kFKeNV44
VMbjAzGSN/LUC228VHmEPgOPtVkhU2JIZ1kndrNviHO2OeZpmPh6Xwh8/+7d
F8r0vt97khjQ/M6dBBO2/z9wvcfG4khyzl9u7dPOkZy4Lx/7PWx6CVo7/Ow3
RbrzTO2agAFn7U+PRFYHQeR+pvjBkhFJWQ+zrNlip/7tw4Z2+2ElAOxXkHAI
TigRNUK3Fliq+1XLsdfJ4kihKGdDz6xvc95txxuQbtcDlNqy3eLjsHSy37b9
BJO0Y8+Y6SsoOfHiOfiAKJDM1Sdb5icaZJbci/8GvADBtc4J8e0whoB4zDAH
6VwqQK5HaamBY0lj0Fgi28vb0r+WXheRHkGcQe0Ar7BXtHGX07iHF44WYfo3
zo+u95bUFMt4uuT+1LyUChb5XUBgNLb3TcpZV9gi+YUJO0OdTw6NbfmsyeET
L4eF/phDk25KO1jBybdhlQZDyVKsgUXRl1PlXeAUXp/RPfIe3q32lBEIi7nf
Y04KlEWb1/bwlAGYDB9LT6WpfBdJ5CDpXLPNkJofhbKxR9RMc6VVTIEe9x8a
teALIaNLgusZEm8gfVYbTU01/d6sLZC3EbABNwd/3v7PvEyMnsZ4/IDZXH4Q
EGvDqlxwLUrYKkDQ/TL7xwer+ey59vBWOk0/kANmoQWSOUAJeAWGOlRXhJP+
sRIu0doAfqJmQDgknnCEDBByKDFgVKungoitS0VxqqxAkwTwrYmpKDKgIzZ1
elzoyc699MeoZpJBKInY7qNl4Kip698D7/1QO1MdNZBm8x0YV3nK1JULlYce
wryvC3fv8+Z3cIw6Q17ubXYIK2pzNKrbiQiZDEj1Lo4JceVvYO9POnrD/F7/
jK/VJ8sovylEyGipzjkrsW2Jhf4gcTfkTXZdFF7S00/Xmz1ZK9rh3imcoQ5T
QxXeex/lLne0GINAoRo0cCl6xAlfCY3kW5SMXzmsCz81iR7tIjYVldWsV+d+
QbBDehNv5p3YmiST/3SyCtPd/GdC1tyVx92pzKemKFNw51wUHqxyof22Gjth
IoKsU7wIblFt4aTVz39PXQ3qWNx3h9i4RlJgjgP4jylC35b6bmJpbuLFEBjm
ZgVnmyVfBdjl1ErobctOSl10P85PeuWkVQBEtT8YSEjDE+HU34X0TaYO3L4W
fOnIgBbGxucbZHOnucPlPxm0HfaHJX30GksEcCBO8fd9IjmWhQFq4eER9JVo
V5pmsb8DpBFwz/8CcjO5YLfY3ohamQdgcMTi3FbcKKIR4NJpN1Z6Noly54L4
XPp4Q/dMPZqD2wmpEvMcve91yGL9ckrscE9VswHLc658y04mPrvgN405IzxD
7iRSuOHdWDBpvFokbX0zM0OWOxMuiucc6gz77y5A5RmSU66/KVf0ZJkDzj15
bMi3Fnj2Fw5Eggwec+/0fT4p3oyRkNem73t9Je7hWn5QNTyiThmWKf/Sl5Fg
raXtdNx3NZC8ueppbDPWpm43qVnJUubfz8LH706n+V49DTA6QYuEqI1Rbrq2
me6auikCdUm1gg2fWpcHP5aq4VZxkStwDCJvKoAqens8ngyYoI6ASknx4SIe
48r+FjSePczsCk6eTEw1Dlz4tlHsbQ48Klte/cmekJNq3HT9vf/bPmI/2zGF
djeWVQe5OhWnfukbum44IRnoiSxQdaW/O4Cdw+o14WLLPNQJFjFA62Hu3lW8
RfskB0344bgZkmGdKfxf+OZrzLSMHctdRYJbYU72KBA/1/ZtoBboWgryTNfL
NkLhQpt9joeTFBd6RMeOqSK5D/DvS1WZRc25qSAQZuW1RiKfiRS1xSYWswjb
Yhw804t/rLfVjeStjaap8TXgSxZjiHG8klLhlxcczIIi7AZmMulumLiNRcz+
kk6PB6FAEOs+4O7O54m6/1ONZ7CRpAnonByNcoEdXYi2fMqoo1JgT/e/gEH6
CeAWKNr0ZAUOyJtS2Do0fzYwR/X90sOT1Zmxz9Mn3VWcuY8LfTokG6PB5I6x
CDzBcfi1a+4ASdfS8tWRgn2f0NBirUAp/e+RHUIYAza+epTpCGLP0/4uVXZA
bkrSxqySDfcjcTfgOkNwLjhR6mOtG3ceRUYLaXFaS+EjvYgqxq2DhDgeqtIF
r4IvSe97qDVbrd5grYdA9D5PPaTJfCprPH97HZHT/UiMjc0IByjDQTSBgZRu
7ad7t5zJaKG0xt3s/l62PnC5/ZyhvMiqpsQyWHmY/pMfP3PPTnkP4Coa3gaf
oYhY5ZljfdOsNSymisswPtWWgfgxs4Q95AuzhMI4oilaEPY49Ivlffc1stKU
FQ4XZZL4W/RAzKxC2grDhc+rcpC91oMsRzTp8LD7/Gx5iaXK6PofbneMAMjV
znLWIlQQS5ldubpUY9YXTLdGY+QmY8Nh3OEU8xkqA8yJTwMvBPqc9i7W1H89
k6FY31LngRguopMtEHesRwhe5kLu5viroKqs/AwwRv+wTvU6ekVdKyVbvJAP
SUl/VbT6I5WwH3Kf6YGZO0JXTPpLjNMVHv/rCwC+XprYCEvLbGBZu9NMOHnq
yL0Z32xVvXUJuD7B8V8lP247SD0fWylfP0IL54/J4u4nY867TtRXRfNIx+1e
0Nflpo/8Xjdy6RsMNFQ3DlqPj8GquRWzwPrw80udIdVjQc+iE94eik5JOYkD
pqDqimx6nK0dztCWomvZooPfgVB+NuBON9qxlea7GeyVATKMa8Ka5yzagdPC
o2e1UZfljLD7N5MvOlp+paz8ON2Rh5RrbzFuxEz24dmHkIu+i+y2yq4zyDvH
FH7pdw2rXrkXBSqYm+LTrE5FPneQwe1mpHinm6W0JLgrn5I23ECMe5RR0Gm2
ga554qko3Y9dpiN4W2CP3o03e1XfrINTIyQmCCwdw2AJwFygThfKTdgJicLX
pvAhyhNQ1WMI72P3d4QCopZ5BCU2I30YTuYWAuYgPhGygrWqKXdKF4w5sp+I
H99kz9O1JAjkqmcBt5RzHoiXbcW/Gnv9EjfCjmLZnpmkhj0X19AA/vtwxXfl
J90D2zVli0k6bSDrl4OYu2F6l9vnmIYBcMVt8wflqieqSSmp7KtIUX5cYPfV
yzKEk6cN+GHWqxZm0vhlEW+L0a1I+jWjje6RklGfnKhnviL9B9+sYbDeN/NM
BqoabbaXHhiIJoMv4g1hA/rEnuHvQTC2RarKzrecakzfoMAcvveQH08JCwYp
j0WPX9L2U2v640gkiPzx1cGeJMTyK6aczuhnNuttYuG0KVsyIM4c37VnSw0Y
q7yMoE9X1RI7Fx9uHFqN5QJWPjTKxS9bY/UXc15GA76KehYnkt16oWgP6Tbb
3+khAkhlMu6fVWczTn50yx7wWvR2ksxZIzHjeA23pOwnT+zj7M2nK2gkWIgA
KCyfTeoUTjwELgR6J6ws+4CMtAudP93coDXT1Rb4dMnlOnb6IhHb5kRzIy5x
e59BuOKndR9kKAbzf03B7hdGV9oFq5U5KzK6uS4ip/1Mng9bwHTpVqT7WHKh
n4CNmlVOt1S7GePJrr3dww7ut24pB8v9ECnKf5IPeRhBy1v0i4KDaqKYuzpj
1SmAO65N4GbnL9/EeSxFAF/+YZ3R2WrG+ypEfUEHnq2dCRknDhYd11C6HSxk
JzIMs1ILeaYcIof72rGanKKIvE7lti1+u/L+VevxvaAz+p5ka4fMK5eHEvoH
kY9HgG30pxy0oZtggJKvwjL8iOsDbPjCg0KWKFetgy+okmFmDwriOs75dBpY
5X8qkm226OJCraSp6r6xgMEIq5EFGTCd3OUFnalxdVxHKVvA09dozH0lTLhy
gFKx3xLyuXGMqlAjfFgw6eYWHMDXsE2bQHLHREaEFzQd7vnf0yicrhREXx+8
nJfcR80BOmYuL18U1iK3Un55I9wFgbhZFfCGJD/CoV86oBMxDBhyLR8qrFdu
5TQIpIvoHbxN0rftBbaUl/+c0JInSy/bT3MxKEwy3vk9DP5nukmZEz5q92QK
knRc105g+EpZ8pdxYWNXijvIZP4C645aNSzr3wmL9+unBEbfc4nfALXiP7a4
WAz9cwnNL3gsxTBV5OmFnJ57dOlMvWAMNu4ex+wVpF9O5aA7vXIiCeGNxn7N
joT4Gk7TY5mRvBrVU8geCTyYuE22kHnlGsxkn0cq9aReTYhXeXDDeCKPWtax
L29CplsfnknkxgJwwSy5XD6QbDvVqa1/epNEW9ZaZVBd8/Lgb/G7yoqFuswP
s54ChW5jePRqTsAL9JfmLcTbyJbuqTHUAkDrEliXBybj96l8YNndI7EqCd6R
rFVwqrcb0hIaXsQfzNx0Djgt371scD8j0UvAfclSgnTNOTL7EjUEdFgmx1C7
UGR1QvqA2G+t0RFJNa4LvLZ0jbGawnVnXgzY+Pjh+vwysLVEUVnc2ALR3E5b
EkMRJyu9q7lTnmFo+YcyCtCqL3b75DOxwKDBxd6HikTdlWFUSQLDictzRM/F
ztRPBW6XS4F+JjAl2ylJtuoeumO1FYRguLW3CkDOU5OnmNulRG/32Vtgy72a
VU39pJyCzCDAYYyc2ZjmS3eGsvR/K4XMAh9hLN7CJLH6Z0XjfJ0Qv+NgdArn
83+beOJrZ27Gpkam4N1wLCPXfpxIFVeiRoaPYDoNE/B6JDU3lZUpqPiseG0e
3SE8i9v7TlJuODX0iybJkRD3lQ+F0WMoHTpdsTHnEeI90vh+LnjumD2nGjV0
SMkAabbuw5LL/KWkm0zL9bCFhlvtWRvbs60yovIiGmYMULSsDfIj3MliZHzM
fUadVky3lFIL8KxsUVbo+HhesuZ6BKNWoEaY4Cmd7OuW6C1zksRQ7hJUzBEd
3lI+BXvBhrs9ZpYwQj4Aep6NeZFC05C2T6H7X8NUCf+X2f9yhpk6VTzIyKMv
5bys9sa9CYyzTm6Y7p6+/MjY2qc0zG3tN/dFug177R8M/P3RQ3Mq+zTDvxRX
MzT5Tj5mmG6vxMTjohO8b5+yRXepYMcnH0oBVyhsMfqawSUbM1e/ne7W+V3Y
tQHzk/AoHuPykmVAxM+32OWjRR4OBzMy/+nvtpPMF7rzkuIWVPpvUlBHJaar
wlVEzp/FqC5FfO3oy7NsfRBXxoomBBfkOMyVHo83spcdM3QV0zDvyXdD66Oz
FWiNrMOBFuDiBvxeq3IQxPWRgGTMApzNX1dcZF8mzFQJ3EboqJ0tjwEqeg5R
l5qj76k7/fnwM5D03pC4FOwG2IAkWpiYzxdvTcLdy4RPpL7K2bGXwPvB+5ds
+v6PCuMct8MYf3Xeq6WhAI22LG+K/uhOOydZ4Ea55pxSBmdmysxvWmF/SDW9
DWSvlJnocxlRLNfrujqENyfwX60HXVj8UIKylsPRYt5fUSGZ07He5Z/vKH3E
R628Ffh10FO/gz7pTBHoNcbdA4GOkXaHxNElosdGpMWwk/DyGoSE3v8Zq7KR
EY7B83pIIPsewAp7o+90cT+n8vJ+N20c11nCYLRHfoo3wmt0eo1U2kSx4/JH
7K88fo9hjzQIpZyDm4/Gbhgcbq26HkDCrp7ictrzNwXAV9BIhX1sK3Jd8yui
s0s6P/Y+SUTAPWynzcEXb/qC6LobA2lsnESbL6Fu2EkcfmGTayr/tIs758GZ
AEBSFsJBB0itgWC0TDOpffvHahESl/paiAwKdVWQVAm4qNP1nohpNVbQkFGX
rwno8uZfpj6bwWfcICFz/kHYOEvB2i6uePhKCkZR8ACxzy6RyXz0iLIHRUKl
TY2C4/g8UNe7JVTHpkjhd4Mktbh8Fj7Ih7+ht/bFuCi3JfdqnLQbVz/rcLgV
LmMUoCht5cflrQqn5uizehDibC5rlsXtnNwBpirmFnEVHfE3zq3wDhnv3hCQ
nsGPjdF6o8di7NtYQF0PaxKtwtzyvRBimTJhSOzSO1RMAGPQo3L5xkeelao+
VbBiTYQyioNg73viOIqwjXihRgkMPKgHWaVlaXPViCKSDDL0jjpEcjvVTH8+
JwQ8q6+HKmfVf76lBCVUW5mOB3Q8JMAPsmisoqx76msVh4pc37+oCRyYcwIv
2xUeEC8jLwLLr7FYgheCWitwqZg/XmuIWHuj4lFPxS+cV1PzL7ApsOGw9p+r
G0Fnn5/ncNa016c0/cXJ+4TeAICO1DyIVWHnWz8dXvTSMJ+nB6rHc6EuBu7N
MonNZVMdQ5fTRdYJjWownWSIZT7z9N9ZNlwxkEjY3cX9aW/GoIABjjTh0fNj
2Kpqk0iT4RDYDrwD917axc2qUcIf/PdYsulKSsH8F0bDgikeNHAN+fmwK47w
n376geCPyKobUfunsgLGt7MG4RbMSDjx1y07GpXTcmZ59jSXyYIHRRhBo/Sv
+WfneACxtLhIA1uJck6rtaEwLh++sFEXy106wLDBfGw5L90/Kao1CAoGdSX6
QQaE7yhd1piJ9JMIgaJvF4BSDma2nmEwoxbFgQK+NQoh8aEc5hx4q+uLmJFC
5muW9MuifFduSwBJFFyN9Q5KWau1Wnn5MYyNsU3Vt00KuLVTakz6BHSAK+uJ
UookVPm+4O75LSzzB62iWBntI8k/QQ6wuw0E0qGXtNokYxCfhGf85E9epWwB
YPko7AX5GNFnRxrMha3SDoS3j5UNMtJ9LmEh2Q52MabR6aVaA1Rzw+O8nd9m
wiZX+9OdSaHhNWlfXB5kS5M3hLJEV/2Y6Vv1FVdK9D3iTuM2nX2ni03bNXS9
86D4PAkOPbTwVwL2pOk9fACboweoyU+JV6TdaOKoRdZZiG1omZQqtpBRl9u+
V4uc46WRCawLnSOCIEsy7dHxltyPg6d8wLy+Ytnoe0GlXnV12ued+hSRSxby
17waqNd6u+f3fBt2Fft5E4mfEAd5cIVJ7Y0N5x0CDqw9sagTUzP0/3EHlGlW
i3S4oDo6OodZMI1UOaH7fAAAEReIHe/NYXOo8x1hvMIHvmENRubN192sP1kY
VdQrmaX7dt/rVaXv3VE4QpJ2exW58kCQZZOMpFUdDeC5i/9oxPpQf6htANX8
OI+enP3jF2AC96zlM2oRBcoq1VuHzLauGsvYW8niqWS+1mKNasJ4jlltq7xC
xgID09ow89SIU7NdJ7WpOxNZRdcXCIPpiPdlWwp+tyOGi0RbgB2NbOh8lCK3
+XiVYg4uDVXgXFMCoiwCVc/shSzKpZJ3kk61Fq+hzOblXqnI8ZZ1tdJN/grG
MRwKKvTkcyS5bqveXqVnKykDFoEVm18eo/PPi4o+LSLsz+JuKunIS7ToMamr
gDUnwQOjjf5sgOMHcGj0XknTmVWt7Bbi6TAVap41Fgy/GDve8AgLGqUTXlrF
XMDT1aVDgNqN+qdUP87wx6IE7sUvlpsBPA1EhSEf1joXszeiZ9x//3xVPQTJ
iYu9wlRvOVpQNPIOB/ZY5DKysy99Oq7TwW2CLzPr5xVJOUkkG+7/G2E49Rr5
e5lBrkWcW+J2mGowKB6SS7u5Mu+oCrburX0AMCoxyOqG6VlX+ctnhodNCrhc
Pul6CJd1yi+lY/4oMYf3Nmzvp/fYmrnn0QtYAYNazZjdr6MjagBO4tlKSGwi
l/DNUjtZiDq8cspW+78MSkdkKC+qE7LwxWToTJasIL3kXv1hoTLjilW424xk
Ce+azdRavnZSL5x3/OFuOpHuF23cnL7HHaP8BvKX0VhAajGgPIvJC8+fWhRo
KCgXrJ7jCej6km2lYy5p164H7uUp/03Og5OJnyUPw4cUZOlM9/Pq+05CzDFw
xtFa7L1Qaz7AL9sNBF0hWXr51Zm8i7DKsc6u2/WkNkFXHovKXj72bkTTY0rH
hIpWA8ZSwRURYMCXgM5aaJlW8RZegRIcgi3QRhwuXNQ9PCByeZcZXv8VjbZb
I8t16FWT/lje6ed2pThnrxhzbeR4YiWsYH3D+11hefCSQt8Z/hIvOmLdLmce
/BK+I79lk1iNCa9P8zVpBuUxPeIS9kRjt2matLiSINYCDYx/MHaa9zWJ194o
ZAQvz5pY+Ga5rKnt/YPjsmDdcela26rU9k9BGHdD9PbKbr/NOzvSp0/TJ8/w
wBLCnluCKp8KVCTyb9Kcg41DfFA96iXY9UeKRy8Z1kjLT26O7wXUS7FJZ63f
mlilH8//InknvIJBviyF1xsPfC0yNtdcxcVBTWrZhb1sZo7DZYK/fTSTKjMu
r4hYboyz+aOPR8zY432bGALqIC+FrH/mX+7sDQNi5O/MXzt3S2p7THVQOGSg
Og3keZWKyPFCIG2LqcbHVGsUEt56l5DKj7BG+bzo369wWRRqQqGHhkQrAkih
JaM+WFG60kgD+y7bucfVRWp2lRBmLen0Oji1u56X9ymDuG8aSe9x5Ptpwacv
3GtpXknbTvU+kFrXnyLsggBG9/Pye5U3NBQBcntATcDbpo0HiiRdTWILvIAL
+DxCsPuAI16ji5p2f/qiY+eXw8dwIGtCGp7Kw0cw0nS98XgU7Sy9A2Nnx/hi
VQKa5U1ENnCBgjHbF+up/kl4hGADikuzl6JeNd2yLWNzspDrRB8VnMmdRCVz
dFClDD9yYTixTTZEYE+Hkmk9M+U1vtxutmONLO2QwNVdlTJVyxMHQdkTFPPx
35mA+dkXkqNXS7aiMnGqw+nXZzV3sPbYKokb8lkCB4XuZemnstHKsz/9ztlk
aUFJWGkyDgPVG1mDuCBm/or2WZfQAortO1SFuh+L7bVcXSIp/CzzyhS6GMrY
X6NwALNrAQITsjJCPPSVsfEBhTZLSgJguvBV/cRd/Vb1dR2Yw/vLRXxdiVoy
QITJfT/9FHzB+XbCUNVOhXelFFrv758IXmJZfCiGWJ05THXGD89K3YtakYry
fw4Y+RQqN0XaRBdg9pQlMuwGEZ7FUlU8PXqOkajBC4D0tcIK08ihCFOy0+XS
5VbodRlgDE303FLKp30PMImruN31KUiNFMQ8jU5ESwqWO/h9Omia40fyGpBH
msFQXmS6JBXJqRPhb1ubNtKEd8z6Ype4ys03j6LfQ5FcT4jq12uX2gcwp6hK
NnGh+lli9Z62pfgJaYz+UmPBfT/4+kI+lLQ6pgd4KNbe/AA0D5GvH6PmQd7P
3OeqjOmdHKNTd8MZqCb3aXDqWFyZDTo/wBc9e8DoL/pMXTG7bSrREcq0czzv
LkZqf0A7zAfd2FggYehjJbEVv+melnKmzSgkbhxDQyMXByt1WnbaFE3sUypy
0bke5IyU0lnA9uxaemasFvgKWXyzpFFB0FvyMEZInD8PWGm8sJuopvwmyFI0
Pmr27PwYUuBReu/Q+fW4KoP85+nVrkqTLpvev+xzm5sr5olPhAKKjfH/kLNp
/hUiKn82hZsXW5YwRIIHZC2YfVL4hFh7WYuwOEGiOTGxJ/u8s8aByzuyUMdo
/w10rHrt7HGZmSeX2y8mgRzObjOMibWIYP4VxPLzxDkYWJlXDtxfF69NPbdQ
M2rNHGTMEK4QlsLAcqVzpO/w808GCLDii6CVtkUv5hf3EvGp0uotfsXYkVHh
Nh6klMUgnUg3QS+8RfHijyizQhlos3OK+C0M6YrB4vkKRPKZ3f1KTzE3FRGI
2sJNMho7nP//i+BYE9YufjuJnOKDIi1CdFFc8uGnDlc4hhub0DEj3GKR9+2/
fEnYrM3j6fWAkQ/mmUfczZ6DWdFPn27ky1kDV5RBb1UC/LMeAZneR1wtwKWS
AO93iuH9wLK5tPX27LB8lepe7AhDs8Rzh1K/C3HT/T0zGUB6O/tikJdBd7D3
ZNUHnSeofbs6tkeUAyA4NYzIDwVEKM7wOOwM6S4bBNWjsCMaNiJeub4L8+Rg
UK4doeSs4XAyqRWewQb8HZSyDjKP3rNsseSkXPHBA+EXGc4+j7rIVtdgSJ/O
aFAhsweQwYROKFMx3obPNMSFoY4GyTuFIAOuFnZUknNRvJd0DUpGe0aqib6Q
GQNEzrpuNmgbLCO3WR2bALRX7CbNqv99U6CRsFL3rGIaZJ9Bpr073SykWebX
DPylz5KY92Ym7JVGVgwOjk4L6sU/5+2IRYklYv/WuTyfi4Erg8JEq53vIpC/
Y9MiFnQeLER8I7g3Zkk/vp1l+Z10bS71ITopVu6Vt9MfIW2+ax6Td4iGJ9sY
BSImTZ9G2fraUAc64Xi8mvRaxY4Nl39DR2oX3oGcyig+WAdhvUVmcOkXnLzn
yJEJVOuwFm2G1AfEVnjs0D+rDaaIQS/H/OwRYToAn1SNAhwSyMZjTyyKfP3h
tJdQ+dblAyp8hInDCjSrJdDpIBanw+xAS8KAFkqZWLsa5aCfdhBmzAjPJybx
xkJcCP76wVkQlbwTPgh8zxyVS7+ghAncZ0A8152jZdzvhDWviJuY9LJF85NO
qCiM/ONap3P6/15Z6rGnQiOw8DNPw4RZ2DnDtb2qSX4uyhiyc82mmfGvgisi
c8H7GAFogIAWpMLPUEDZ80P1/r4vXAmmYh+nnNkBzGy3JN7UKVmg+2zC8bAH
vnQ4iE3zNp51uNa926L9VGDRjqNUJONKFckhJplivkS7NMkDNSJaJ3Wv1hcH
rDjhgWW5Mt2VJe8QbOABE48r4UsA0z5ht352WhZNhBnRimZhCl0dH/cu2eCk
RxiW9y4qhjbs5rGEF3VUAgpunA5uSzllA78X6ZpLpLaxj9cDtmkGgJcTB7gI
hiEt3oE3CdMLqJeHgsn98f5v9IrVbgNAzbZjtHMV0bilB/RyHb+K5DSUj2AQ
jcyGxkKW3598Oa22fEBaltzO+ID423/mvVgO1OVo2y6AUOzbP2oUkjWgj6bH
vZBtTzmF4Wpwq7/OwZ0enW2bSyaNcbOVJKtzxwqI0Q8Vc/lA3PwgvpFR/Q8s
jyUkOlKPG3OCagASjHHgeOTi95Jp0+rSuzAew0XnXHxzTZqjr2FSAKMi+3r8
HNvV6CS+4DZvbhAIdJ3877wHpU870e8ng2yXXQan93FpMit2fhVKLnb4KPhe
bMitJX1YOq4WfLG/fsnte8XyZPJHpDyPhKiA8j5Z5XDqqT9RnJLmeg0fyCfY
atfJGHEdxq+G0tD4/XhMQRJ4GSbnmqiHUbBeNBreoRB12tUDAudeLjCoj6WE
ODis+IcpImgos49PRQ5vVDXS3tBJs6+LEfx93M1F7MYThQoh7qrjIhBGClIh
al5vZD6JyVpHjZ0hM8Iod65MCiKj7lIqbSugKVxnGu9dPcxAL0n9LlAIJdoU
KHdNeH1FZ3tB45hN6REqRz5QX8xFrVL0zjiJXG6yTSA+jPKvGSnlUAovvmb1
2KFNcBNMJk6wtOPOFeuAaoIr0wXzVrSFz2Q2Q/ZZaIzaa/PNzLsmNfOP2cUs
C5LrE4btxiooMzNy93J7l4iHL0rmWJF9XA4ArG7iKDfECyuEFgL7nZY23T8f
DKxqwK6j4DdpxJEG3IwGKBtJ7MqITG99VX81gbqT+M7SuTWEG+EDG005xZMX
/NOlWDuvFiRtDT+q0NdoW5Q5+jQUKu8NPn3HdqBBq+swlNAU4DxxJxOu1u9u
IztfR+nuGD48OEARVAygS+evWK6u0aDssoC6jIkBw6aZO/ZXZ586nvZyBJjx
6KvtlZHMzW81pTtbxjtBU3cvocFqeyp6woZSigCZvfd02PzRFZaCPiHL2L79
FrxElDvmIuC7LXKXDZLHXPrRPUZ5FO5eBU9oYlA7Y8eLtGv0zqlhbCLnAh5p
qJWhvpXE8cM/7BqIwQAAL87QMXx3+KtOJDqRfsCrO0poxRfLbAt4d8WviHXk
mrxszJPCD2hTa4uxF+vk0weP6rzQoHiV3KHi8u3dpB3qThR6JLbvEz9pQ3ob
RvCxLFY5ANTUDdXKtAnPrsCsMNMG/oAkkWWJS+DE6UknaL8BJPMF0IKVCUgF
lcVnUQRfx2cW/s8+1qCNi4KT+n9RWkY23K/J5+9wzpsR4bp0DY/5Qoeqdusy
spqVjR+ZWyxI50deRVo7RuhrSyTZf15ndnfFAFa541/08COmRKCbsR4e7uqA
ChK2rAjz5CvdQB7PdDOViXjOOzNHwd2PgBo+epceXDlQAKMSmvwewMOGkb5D
EBpDkjbzMsVLfE8+nF9iXjoBxCHIIsnm44xh7AkY6ve4brUAcpDOgeSclO36
RsQ8Wzp9I1GoCxYxAXAXVSVpB9S51rzpUYX/IlloQLsb+UEX4PdtUcmj6Ixa
DtZ+YZa5R92/zEWjtsJPcA2U4mlhPrOveUNLoXFusRgpqxoXwiLq6t28HkGp
G+QVjU2xmlQKQ/DejwKW9cP7q8pICj2Ntc075t+nYQNb9PntOQf1rbQtIsAe
tA421GNm0wMWFtuX4VAGBUf9F1yOeJtXuFhZ4fVJTZfNpvdF29jyYQLr+ufI
Apas64sh8IxTn7NIzWkA5W/sDHBb+YP+IXAl1DSRBC5KTRFoFNE02mVoN4xu
j3Eql73ZgOZ/gkAFqYGvUeX1DnPI6lmeMIbNM1ghKn0nsUURklTEzwn8Posu
/8eiLDjdbEDoEOGSXVuYbosQYsMUwd8Bwe+4PbhmHX+sEg32jGCtCTb8OSwH
liw4Qi2o2W/K38sEtXB54LFJqQMlebcpp++ioucANF11wcr/fv0ug0R0+Kv8
FHqSDxaPnd4uCxLXaJIhZVM9o/WgyP+xbLmHa8wqsX36Q63/tJaO7J+wgGVf
BnpjSLpxC7DbsRqaosU535d/t4fpuCDcuvhdMtqFOdnUox8KA2hSq3BqPBwk
GTD7wx/XGKz8cKwIjw3iV6g1wxMKEYN6v9c6Am5xQDhZK7/ZH3bB4mJiXP5N
X83OmG6qviRIn+d6RrzkwDSgWbF+nk++rNQLOS5MZ9ps8mpa0TFuCrF8VJBG
kBlVIxDwrQ67w3cyQDLwkuJkCFsatQqqvt+PJVU09BJQS7u1LkPRWnGrq0OH
HvEUQiw7HRZvr/zGT7fr+aLi8odd70viET7bL8S6fOpIenur3oLcgHNsjIL5
CBBt5opfD8M1rY32RpsFb92j90VUwC/cner/2tXR3LYEGRNlmqIhBNx0KGsu
Hz++FAmDCT9TFZSKcz18DogBMPzN/bcA51CZ5fTyfrz1SZWA9NSnvHr7UOiz
5wIJ31DXB5VCoEhxgOqIEMZyqOZ2RXYPWnJh9+nv1Tpy/RpYlos1eMckgMHO
R/UiwEzBNcYj8xKl2GhXUXHzEyajD8Q87lf+WTmmwxuOKcdcHr65PRbft286
NYucnvu7S3B/AOph1vVlmnmlhLb0XgBI6DMt99v5TbGS3rFZmaHEhXv3xXlH
SGUQ8VFO1MMXrMYgCoLGqoc6nHRkvzyh9zpciCiwWJSTHtopbFDMtz+2Hpl7
gM82PYhZSjOUrSn0YCnpcFQRWmxCa3Zy0KNbNZtn1sYzs952fPnxwt6kk60d
wReabv15C1kXddYdYHbmtpnKGavhBfKPwF/g28WL5ETw+oIZPk0T0iwmzLYe
y08DV2BP8Zl0XgtdrLGYA3wLySgtaFSpEX+Jq2kJI1YULEkZxQJvATOhx//c
KiwpUZoHBz6aWNL2EsMua0k6JJ4ZX2+sJ/F5/k5T3yKGGmFToc9VUrxJsfmK
LAoLkHfCA0+G9I+TvyCKZLETJ4KzfqccUbXEOdVDMPaQwOmOPpFk9pJt9Yko
/crG/7W0XVjUgetIQk0VlKpjHVSRKC79OwjxIwqaoi2h/gLMqZ9MQUOUUhql
JnqrQCueVRwWdEwLfxCx5/NJPEi05mI722nOOnGqxxomHcRaoL4cyq2T4Q7a
w4Dwu2UVFRRXj0lWQIAAVQnK43JPRHuAGdJGVnHRnMqMqdn69zP9wL2rlrRi
0bXN+//5OpGbjOPI9p5/8pl91GtZJcItc8EAHyX9qwsKO2SJ1SPG/gsX73o2
ICpIgkecEpUiwo0c6x4xfVUAOESo2b6qEh2WiHFIIR5/GfOgRmaDKgNWGyhB
xjW27Eck0P2yl6Ol+NLYUB/n+9PdccA28EKtxmWo1DCgq7Ng3yowcRgHfGKw
e3O31+lHBcmcoo2q5LhTb3BjUyRUwjScWts6dvK49nJtlN9lEGOLP4f2A0dX
lZ0sQjWtZTsKVarvGa8zLJ1mcMcWpE1368BOP98JthHIQ9Uv2ziZTvxsY6WF
qW3nN5kIoA3R/e91p3uA1t86QmibXRp7Kroa1un0TSDljIHOSFScdESGFUEW
A84oSEu6U7lPsFm2g5gHuBEhuu1oNThR1Mqm3HaUltxqJWOQCwK97WlOT/Y4
z8PEno+mU6UQfK3Xxs0i+TuyenGlbS7NT6NhH0D2xbuR87NgnR9r+qvQYMgq
gU0BZUHo4WNd3rWthc9Cn4lLaUb88XsRrTPweOv+IqexvGIHW65AU3/ZFlU4
IEq1YXTZMntqnslavakqlYDx3rgZeQhThD5IXXxI9IU22DsTMovHpiPb3Z+4
OP2Wz8tXFVfc6pHh4FMcSjUE4UaD/ih0jDm0rxLrSkpANAFH97NhUzCDZkOY
n2GorUmvvHfMG2Zr3eXPzxMhr2/0D1B1mMQPEw/vkeUUobUtg7qQ4ZIg1r1R
B0+WVAvC13UPE/P+QaDSyGqchtDeVTKBvcnGZkZCB/mDUsxVC4fDOFspwrEU
PKAvNSkLAV5jllegZ9WwaV6C+BeZ0QqS0GNLbYfVaDdeLWOTTWIdtTgQhsxu
1cdZ181iSlST8jskXXJKfU852GFpaOtObgq9rXnHLfrYmWMkW0bDyYFuAFY1
+ILhMYPtpuCG55jTdSzVvB5vOEB6nEQBZ3KuXA7CKph1Ee9qVooLOM5zfnSY
QAr1tBXnVa1KTt3EXBjW8ffyPOtE6eXh5Vt+hgDxde5R0ei+hqSOiToRykcF
W4JD4pmbaLgGiXBuTRw4FLURbiOs148iNnBwoBdIxN4prD1Z0F3BWGJ7MJ+C
rlhY81o6btDgrGR0rPQSdJc0B0FEgRdWtskuBaYDplVkVdvoxsnpKp5RKq95
AbsOx2KcLh2lLNX0JA4xQRPgNIUev7oTnZ35YksFvBqRINHfH9flOjDkCcPd
WXiWOwXoJZjHrG0OMbyY0Y1ewonF7PGm4v4zTweimnBPZfrseen3D7uqSmiH
GD2+qBaCASZ4rVNZo8b+clsSmZGa/rIQLiA0Ni8HWfQLTJ8uXcnFtioP5Foo
sonv3vocPmqbTL5gLaI3YGY7KtGr2NMkPV+c+lAIlJ69Q4DVmVq8hk8mtQYb
rIopG0SPjS7u5f3GsKc2Hv8CLY4xrKphL8XSkRDHxxPSSBqYbCVyAmddDQ2F
nvgrnILzEEu2t8BtdmGWRkliadn8h8VlMBj7kcVy7Ez0i2oGYxPNsmFdsX+a
bGsdFvmqJsSkk7bVpTvOb1fwVsI4gVFPW2sNdk4V0jPtAOy0b6OkJSSSxXPV
YMs+7cASRLz4tLbLqbGsvWShL+DIPxWlx4M8+O5sHlcYil9xEBKq7e9AQXpM
FchhnQEjPb4yOKRELTQglneEBuh9oQmm12sJFrhM7JK92R9lrSKyFpf3AH8B
/lHVPa3klvnwC2P/eJ3L1u+zLS3wxS0Lu6VoaexbymFZEivTT4D3C9SHexFn
iwnFFYKx+GTgN1W5ACyBgUy8mo0Ovhcw5jljgAu03IWMj/Gg4Za1fgHGDXpi
3Z+kf4DbtofEDQMv0GmhkOZnX9jo6cWGGvP/+95cBD4X8ehc9xQAV+kabljD
gKoMCpGAZtCHBROEtSaXVs8JttH8x77EkrNCbFFU2yJ+nu6M93stbDw1hfLy
ipKHtijBugjfv5BzPY1ggOjNphaxEWgBEsMv+PzEvlMi3j9mKMYM53NNgpGx
Swrbrf6Nk9jvPUg70Hwv9xyH/On2a4mZ28+9NvsUSdVOvF0MedCVlPKstvDw
12udfZQsZE1rIpGTTJkPfboRtXJFeb8FekhdRDFM7vRsq2C8LJHpUDElJYga
wpnqRQ1DWjSgGObp80bzvIZIpAfWi5ZlQJ9/9pzNgb4x9vF7UVTCvquDF5/6
X250EuD1H1dLq2LucwmdC6S4mQ3bHLBbjbvHJTHaalbaQkOJcJJnyxEScVIL
fbxDDAVqwPd1GfloqgRq2rpBlOc/8mHvMzgWbatGha6HS0pgotdA78Kf5+Lc
Xbo0LvLQAqkLNog/Uzx4qk9jpc2yLIvFgUB3KjHUXIxyy9U9s+LEF+3gzKNW
hDptHeynQEDtlCtKxJCP+FU4bDmoZPo7sKI5sz5HuRHOlZV046+SHSLLeCII
kdIP0LX/llRha+cQ9srb7gIe5ZC07gKscXEvNTzH601yaX/hQGcHUdqvoJhJ
a6Wgz9BxnfewpOQGFqhUIcuibTLid/8iJGlIRBbvrnR0/EZTZQ4xmDM7G8CW
k+YrFzgdrxMyz57rZ2LK5fntkvphWWcgDJYylFFFG2mAiXA1Gf5Sv780ea9S
WDsjg3/kTxZx5Db2kyxDBkwzzvdE7589+ewTNxJMF2TapZr3i2istHRCaYj+
Er0j4Rp0m0SjXm27xBOkVAmtCsQQLDFnjQ0nkxlED6THxMexwMpu7VHuqjOj
pKPakuigOXTWtaZTWybPY+AL0MGCNqUtEOyuCd5yNPPNJm/XJaxQ+zoFY3JH
qjl3xmquX4hPflnYgcAxBxiZvv06T0sCTyRe3j8aRsLahM4HD2EC+aBPjJJr
F43ga8NwH/cRT6NLMz5n5T9FgERrCrAa+uVszqCJtCAE9qiBwxncigb7G8nN
4zv8dikYdkdWlyj+2VaosF6FhC0ZnFhPEILnyoSdrMJ8qPUf2FglGqk77Q1K
bJ1c5DJzIcMlTvru4jvwxU1DE7euIY15bS99n1EgS9KanJmJ3gQbO/81EHI3
EiUdV7I+OjgVKgcSJICvpKQ+JnJAB4vLRozgd1ILeR2tba5oN792MyGfpods
GPP7mc6OOsKHNyFsg+dazoipde2ENJ8yYG7WaMDxCzdyURKy+i+1kpG6AGZG
KZphScsD2vVRaAF5DZdDafms4Upn3fs03BdU0CfzzHk8FBjTdvKMCI3/YvF9
3TwSP3zt01Cte0QCBvolC9we1QJYU2nEV/xU1Hb+KY1IsZrfqXKhhUx+fhiZ
tz2cy/5UT+9GVIsLCndwSevUub+B/e+6nPALJsPo7ombOAU1tyZnUSIsldQv
STnZC8w8hBGcnzGJYH4ut5mK1Odz8leHC5pQlo1YvQDG51TFSjUid5iJhNis
jryaK7PmSDEyO0ty+EsAessiJrLfHvK6v/LBajR9Dghx/dbBi4wOr/q48BOL
BJLu4Hc5g+UdqphBNMfPuYw4mIFi5pceNwqkrFV+dw0BKNZVGvUnXUZqox5R
ux9JN2YoUQl/tlNwg/2B+8Ot1mo8l5K2LeDZoJFRq7zcREdllHawNvcLg6za
x6kn50EVwjW9oWb4h7Nq4VEKeiNq4h81Rr2bq3d6I83PXxivXGn/q0ayY+UN
u0K/dHMetqCs0VobRkQvW+78/aIOCq+9knfRjAfZ8xroyjLrt844Pntph9dl
TyMo9LyWQ8HCwB/MG17IF3SM17hcQdffZs2QOhrykpndwQf14p+d3ly8SN3U
Ysmb1xKoQfC3okD71gyWi56NCx+Pr/iG4vMkPS7YnHefEYczxjKNeY5RaiQX
ThblVOu3PHs+3X4OClGwEwkcrf+oT49dAV4x7hGySCsQjV5IlOXvI51NsYQE
vHTDvY9HvYd1mJ2E5TWPKDO6AjfEwyxYHY30Ti45afgP0uw0Ga5rObVHlJnS
9whkgQohTXaKez5XzEM3+dFlTZ9Iyzu/W63Pi1yLQI9IgOCuiFjsKID17y6T
THFncLuNCe3rimFyR+dKHtgPFIhcxeKdqewuJRgeN2G9yoTWdBZtSHrfZ97g
xMGXD4qLmi78SVLv+tAO56aAYQysmUEkNdY8UFK+C4a3KCrZFdMShrkXnk7G
z33HQj82NeWIC7vcuDjwALwo1LO7vNfVIhOQHBS72VCHQaTZdUG3deAT5W03
UCdQGtH35L5yaBzcBkxBIE05pU9LXEe46PsAv2da5AH8PZFgedDbZ6GxS1O/
jXgLRuG8oA7uCIrwD+Bs3KnDAW995P4M6dkRYhPjdmUpLDzqA5wUKgTingCa
ZebLEamlqsrHqWvwEJbfD89J63xlALTVMbDGbD3XOam/QbW9B5HWhvUE2BOT
MMI9/zPjVl0JghgYBYKE/XviRll7RrXS21lzbvzKTfl7WxDjX1UrBJofAwYd
BP3ZaXEtc3La5B6H3mzWTTS0csnTC2QhRjJ9AlPr3zNtaiyB4L1l+wFyT8ov
whv+TXYhRkmG6S8smy/kEsF0IudDYws4D/6T88fpwa5Dvn6/ag8ENlRY/y8x
MtWCpN45g7q7trBAMesQ+e0NVa7f00RPL5QW52LmBA2N2sO8mSCLPohuDEJT
sY6luYaLfc9fuSYUqaCTqlTO9EQE/gKFdL6LRwUn49AGT/hb74XAipgbyyTf
7wVfk8Ki7vKKhXYjuBpPhybEvfL9aiE3DULqbiqnEJR+pAhuo2rCOj9y7tW8
ExM/wuUGDWExpKQ81UNn4ibO0WfYCHFaGmVkoy010GLmVoKQeO6moMcz/f/g
YhjwNSMc1/1Hzubdqps8lYFyy1zbeHEQ4s6mCZKtI6nSaESZ0B5CIuKsx5JG
YsMzipMsN0NkebKp64Bse8+H+oWK2U6YMNbheFKwUwdT0u8ObloqgCl4mATA
97ai1iS8x7EQzLnmL1JVF50TmEblZ4ab6l8hZ2BJqKLceBi7zr7y15J5uIA8
EfSCKyp3ZmeG194/5wMZJmfUondDg/+X5FbhP/BXkpyOnAgUmPl+6lFmaA70
2llym/5NmZv4fVveKabfBKUdr1KkrL1K58eqJ5kkjv+e08H8LmMmyAm7QrJo
2KG5UvHG5if/UVRL7E2A/p5dd/Ry8tjyYKpNMnpi+Tkcc56tYzPCdcyOO1x/
+DMHsWgNaMf/5O0Rx6/D8e14ik/KDifJPuGYfbqixTLzazAiEr31SPfkwUuQ
T+e6X8lvIaA4mX/7XNpjbqHOihIUUB9wOJC9DpAvq0NS0z2IGyv7ise4XSyn
vQvjPlQVZ9ufw43e0IaacfQW55SNomgu+s7e2+twrByS6TspSPCg/lwJJFCt
wrlgxXkw5nd+BAEoxGSLeMs37W2J+2IMvxwARUdozIsCNeJf1oQdMXCImZNO
ggmJtDO0L9wjX/Jsr8G2HTKgiQ9390jxJ3k+hnymM7IjIZYZ4WHnEAyMEY2/
93mEO78714cigi33kjEBEmWTgNoYXyHZlayox0vEupPLdXlXtWkeUPwHjHC6
d3RZxVVtcMPaxxKwbvbEWeRJYRbl8NxA7rXDo9lMR63deNNsOXn/DDL5YsIa
lkT3gh5MoSe3KXkwe8eaK/f7dI1QTj/hjpqAwpgb6rO1JIcHkBBqbK1z46b0
JLJZW7jUm3RphrADCnyd6I2mfEX1GduqyQ++bWv6/UmZEPySuOd7b34E1ows
N/GVI24Akm93M6RqX7bVCdoQ+TXu96OslbQ8J7aSEFASQE61jbaFo17soScS
7f6FKW2BwqYIXB7bbiYJ+X3oXByIqwQILSOLOygOOe6J8ZKk4Nypq2Ko4fJk
uxJ7w8lMDYqTEmSmVQUfL8BF9HsXfkc6tmlgv6UzmSNSpKtZmRSNPeNduaVn
hlU8pTp80vb5l9pE17K0x7InglHRwCHK4dtTVSN2QU7Niu3+4TmGOwyiRxIb
FA83Gb1k/uv/tF0v/SCWt9dv00olq/4fxZQ3NmhEK1RcSFVJtQ1dAfZvDDQp
RRbquvCCaOExaMI5T1MdxA8uHJxKv/MWti/+3FB8jUb446wJPBcvM2IiD85O
eIzZbcb/Gx3MeFJWn0oAReMX0brOXdOaot+u/nm4nq64nA95dhnJ5jzqzMHJ
cEHM2GgJrWF6uONw5uO+jIBCRCKCTtMqnjytiSDAjJEbg+ivpeHnYO7RL3lZ
oG0gtubDO/JrNpMAIydIUSgELYQsSkWSSR/nNMo/flG1c6fnJcJdCyVeKOHf
T8sXBTeVB+8anFOmByVv7Fb6O2ChyEu+YXYDEITdzF+eeSsWEwbo8HA6EPaW
+P+PpdYYEZHxhy9SwMBNLce+1bKdxupeoBF5vGkJCRBKYp4uKWWoIeIowlOV
6S3ld54+uLNPclRcXNKd+8XePL6qUgPCY605cFwSjKMUfBR6Me08PNzYjsMt
17KOhOhlyUGhSa5LNNvnKxYHC8q3rrnnUCTqAP/RUId9aMeqjdTMHlXUkkVV
yqrtAGzfnDoZMdTE0tpp3I0MUVm/pJTWZbZAZfgb75QEl8ZYCLZFbgpaFjNM
N2OpE7v79fJG1FgyWJ48R1ziA/ZoYehyYb80kdursAhOUbqAd7Wn98Nr1peR
q22YTPLCq3NU3UfWupLsVQqV4LnIwGhBqPNWydoi9MP7qMck4xaIA8SAs0yL
Zb5ddgU2Pq7rGRYFXgqWSGRvO698xIjIH8JoVMwDSSaRHg7OSL+Yu1L6tayq
yunMaGy+4CRLp8ZLv4z1HEPAd9KVXNuY8/vm5ov3yorZ5+vw0udvRGVhDh+l
QptC1lW8dWEYZq7VBclUcp4vFOi1dQ/3PVggN22yxmkIFRQtUZorq0y/hrLH
gYT6kE9eWNzOUrh6Hf1wkWrbGZM030OnFGT88XWjQQUK72XiT9q2eKVNKZ7I
144bdOV/V0rfmJoo66Ualbsd97eEjdBaWzTk09rDTjbA8zH7xJpziII9x0Q4
T5Dp0gQ67OvUxJGe8m530W3Eh9nOwEE2LCVSIPbDXESFvKQy1uRTdjZqnqBV
RaFBa9dNEmCQvsnQsRlvFCiJbHZUasgL0vSEFM65a/jKW4RTEvi5z0qQn+4c
QY1VYZrtpDrsccUFxm928omUBvOUr4fhgj9XaK/M1yk/o1eK49bxzgRTuNIT
LEvTb7t7TDXMq20sHk3MRvTrw3AwQ1ETjuhCaQqHj1jN7v2EVf2SECYeemul
0B/7hmGtrZQpQlamproRLxAROeGMkvCYC1Ellqx1AlNv8WqVrfI5ER1YpxQc
1PdkyGNpCVMyCcFdOqc4mLp3cAyu+SbgJLT7sOUhIduzbeDPs1kucD41J/Oe
iIvbZeDj5D/macCEWx9NIHyKROlQxlnyyRj0D2UgZ4YHPugUuRSHIEnyJng0
oO4aJdWJP2cJOwJW7yiLUDmLoyl43tns/AlckEND82OEytO5rDZMliuLtm0F
kl6Uv6WNp2egxU+MBSCyirBg/6MOujNEPiu/Brn7LzKlNbHnhfQ4vvH4fty8
tPQqrIJYtt27CZfClZOjezsQw79bRuH+rxXRb2D5QsLFWgLPGPZhitYKq5v8
00bGLdQ8sWvkd9dH7KnE9fQDaUeW6GGsLPCGtI5jSJD4lBpnD4urI4yRShTb
vf0EPC31QUUL8yvMgTR/VR8vIkvomztFr3s/RGVBAOP+A8di/3lVrkSRxrVa
Bk8vXLW/VZAMPdsOcZl2B7Ryls37/fgiGAupzfWjvxPjcCB4Gq8pJXwMC5JD
2kj2LgZmpCo2F+4ftJxj54xkme2xxiD1DSZ6YvHfToalSYFm86DAblcNZEfJ
71aNdgpzma/MtnDav4X+szJHDlYaQJe6XuNb01WnFS1oJfJ0bYMl09p3tSA8
bD7bAth1wlhNCqii+74mxpUgJgXJOz9ue6YTu015zPtlVkhqFFeMbg1787J4
CqAEuIbsd2NKXCj4A5MPtPNLwqNKoNOx7A3QZUvJTeul5qSGPDFZJ2ohFKBS
3rv3/iMl9RUQVYgpUyoyvO3J//QXZf7CPux4rDccz9nfDM+TTHm/uhmyEjPg
XCvWIr3RbwvUS+1lkKZjwtWf36LUgKAuzel951baPeHaY7JO+mZZPcicbC8x
gPUX8koGA2yq8Swbl1zkW837wpwwXL9nN9+yhrG1I1US9qPGjuaijct7Rezn
FViJ3B+AHSspO/Zot1s0WE+vOGfEJDGx5TX537lEKjiIwcv2AmMtQFiMJbmj
b3tg6bP2jU12JcAgF96ot/taEJjNeraAJkBN7iA6g0Rx1U+zOt9WGrswMa28
nWDjrjfr02bfFz+18u/+hTw6BoshklBr33SuFAfXO4isHSjX0xeOitVird2D
ZZGeOpODca9WAiTy77+5Lng2w0iKnb1aDJ0ULUBk5lURfOgD+2F0L6YCAnE8
dPi6Snx84kLWa/irmRXbjow/kjgokp22k1vAGfpNI7TiE8JU9QE5GY9Re5X8
O3YTAJdxGMKeNujUh0I80ebKgr+7kgWWhXDt6V0VUs/nKA74UJgu0Ga/cfcN
qfAezSs0+LT+7BiZaZE1RxJZU8Y+gq43SF5GqaaQ0yTu6ihnC5g7EkFndMl6
/2rVlWsUuNoCadn86fKyrVZbw3sblzXEtn6XJJUucn0A/WxS38HpSQj1ZcwX
zYBJC3/rkaYYaLwgIHZehHDdpLl1nrbDxkZXC/+L7BzpbkQZ/CtxD7lhsnNJ
rApIHk9WOEiVJZKXeQQ2enuc1MsczcrqWlAYV1LpoiMrxkzw6CdGW4N2OcSA
q0QZHRNRfc9bgJ9Kwae2Z7x088w6DbXD4icYiWNJB8qr7THZXjM2T4MLXO/i
PgFfxhmmRh9HWYdm3hAIEETvKhp4wZA0AnjUYyBTt5g2IOSraJUJ74ydtiRD
SBYEMywiteTwB2ZgpNQoSO5qq9w5muISevKP6CYvG/a+hWjDEVlrOUrEhpHW
h9XR9rC6vt0duQIr8LoilMZqK39IIZ3zFTNLtm8ne8oHRdrXxGqcLz7HdeW8
5sMw4YgKVdxABNyewZKC3hxU9kbnbALyvduYG95A17t/552G+Yk8GS7V/5h+
vi8VMYxIqbhrwssjdnqYaDMPu2AYyv5NGlex8WoKK2AiJWOtUKlmVihCc4RA
6/Fv0DOY6Q2aox0okDTMGL47LMzg+hC+UM9o3qtppXyVDM3FdmbN/vOe90/s
4sOBjz/S0+ugs213C6T/DgVfNnBTMB6yR8uF85E9knfUeOqBjmKU5WRnoFd1
SXYkfWu1iOTKXWw3zqeWgQlvAZY9Ev3x4GbB4VaiLevT+LfAJJLIDBobcQX+
LQHObyCeUuYaArDjCrCfuB53jW07UYE8ntuDHHRmNUHb9qPxvjFiAhi0bWm9
5Y0F0tuahmYenalH49JtpR1h27eWigT8xaqhLlG9X6hPkEEUDv/9Jv+kulOK
973QZLrph7vOd/r7o1MtTfhNsaILfWgcwZqJTXq9eTzVDEGJn8eZwOhEorxR
uKMpPlyMs8WRzv2Qy8Xty+Ewkvr4wwkyP5lj+E5xFz9EVg1x/iplseu8YPUx
P27AcOjDdD3NS3PmLWmPvXscCtIw0hWeTa+9OICoMBxMsuHEAH4kzNEMBQrQ
mSqWiAclPi4dw7RtUXo3goJi1EyoyGCOJLvfiWCJNZ6x2OA8pT+VOuz1HHp5
YWBvM419fV34tc7rW1e6bgDbXsl5uhTmWwAeGRCnTyFJxT+SszWHdMNrVoEH
8mgHNT1zRDyQCcYpvThuj1zazL+lUVGHdRcZnrWFUn5GhA6itPdSQ9QEcNKT
cgVRw9+71D9pafTVep1NPvsoV8L/AyJjV0ck44j45Oku4plwUs8zV+abenrH
TkEKIpA5Fc9neDnBTz6I8teAxgBW9lEUnmiShj39NcxN83VDpgIT373oyCTC
wPF4wTYgdCM6+mjl/oGlNkV6ubjMLyvu2bZYSN01jJhCVu359Tl4P67H/7Vu
cvHldOTSTaUqYEe/gRIOsM9XMWf8SKve+vTGhNCt+CDDdJTe8q5HAkzI4ujM
jkjzWaO7imfB1kRVyTURmQEzCVfd1bueGkbc50Kxilmp4BLXIwrKbMKBU0LX
9o4mTp2QYX54A2GgyZWpwLeG8k+o1loDshCWfX6X2u+LHhRz+HYsDQGsscjq
8Q11RPan+2xSvCX5oK+VEFvowG8aFTdfmX1/U+aFYH479KrsxqLW/RXzR9YR
lAB/Xe6mPcfit350Zov95HaCA1jku4JT12XXIP79Yxze9a7MMX4Y5k1Fga6O
SZA8/7JyiWUo2BcDt/hucx1CQMu/rsbbP0WJKraU2s1QBeU6ltqbuLEQtZsI
fxAn5UMYc1kTTMu4AqXt6GfHLUNKhXD6IXo+nj2icXAOvU23XU/nvSSmDazO
ZPLJyPVHN3Qbr049yJ9OCT5J8G9tbFHnAp8i0XF0dYrq4+v0fkPNO0LNojBy
rHkbx9PS/JHdWng2oeiZkmOKuF6lTsUdfIMAXSf0hGqRn9Jmb8eBYhyqf0GW
JzJXENOsg3BMKgC6HwHJfms15RDLLrKuHUtSBdsSURBLNJDOMxIOIkcAtODI
zdcoWthBoJwnDWawkmmj6lD/iuuPct7GtzNmvSR3XB1ebbpj+nX3bPLWD4fN
10HXj8KMQGfNWGDPbzOGU9w4S3M3kGBGwk/fFc7wdjAwvOkdw7d159pnKbAe
tZzMq2H0c/KSgGTKfK0mArOJ9rRiX27XeSM4fALcJxTq6WC8C772EcfW/6N0
5NW8vlQ/yIPsf+hquju2SWCvIQ85/3GHJvJFh69+u6uFu3fTwxZZ55DYP65c
Y+aPWXg0UVKCVcD2bU6UkQxeOBM1fJ/Y2JFwOYnp9i+xVdtc9TPhKCN3iu2l
IsI6T0NadLK5IyzgNjcMWY25gCDuoPAaiMyt2JbofFVumn8Db/zh/SR5hPii
RsatGSn7OYJ7daOLlDiXaMB2eT1tDO9YR4jx7e4jp+Yo1uhdAH6CNUzr2abl
VTfZjD4N5pz8vLQ76YvHee51NatkYF1Hdbg0gjmMeCSVM4yb8JCy58EQAKbz
XW62bUQbLexdNPFeG8+ckGtXhBfGgtgbOr2THFhi2U+QQKYVz8rHxUFM9JrA
UGF+vhQaapgL0lLX046FkVXdeVNW+pknbAEtZhYeiX2IfGepcofuYpOFxwLq
uwOXVGwwPj+M1TCIBhI0BW+GugZKyELryPnb/sPhJ0RXiDXaHUCr17PaR2Hk
DQcfoZYPEhrSDbC7GapisoXSClwSE3gRQPeMpCSdhwySkd02+Tx8Fkq7COi6
3CsbupBeZL+mXYsnejXt+1Jv6z+5IlmVV45iZhgVkbW9ZRsyOCU0GnUz57SL
/b/bfiayn7awxoA/uT9NhTf2n0h1ABt7UxjXfkEhNJOEmefSCiqFtAKFxNbM
R3YGKu57R39tygi6rrf55/BhLgq4gcsQVnJDKJdwYtJ8JBKh/BdsZhRIbva6
bJlcRajWqa71CWDC/4ESPY6xUSwu8IdLya6UytJWO43nTlTeZ1B0WxDNLC5y
YoWtSf9R4qIm4LN+gaWjAi3czS2kniZJBeGiZYb7JgJILlKDMBXcxHcOEGwM
sKwdzoeMzKFqibGQo4YBS8CKNUU3NSbo1vK0PU/zj1uuQ7OIlrWMDwaj2dyy
X4x67k5TYvhy6YP/pbu2+4nf7u0bnfimm/xupaF8scHSBKbwck4MYwhV4clE
7na8vHPiBp18/qKb0anniEStl//ot/J26Z5HdnUci3lMmyKfoue3L3/IYr0p
0YxyZ188mVA9XxBr8gJm1TqPsSJ6YnzkIioKH9yvqU1CrZvCdkS5t3k1UZVM
Dn6JxnMndzQzImxzPX+XkKWTmsIc3g1nxupVmVB6LzYcdcVuwJGyZoG8/mDM
AlWip7afuIXu7RYsb25vfeQiewmLSgztYUV5/M9MsE3LfDMFWPksKUmhnsA0
gOBxJYTXVOQ7jqekeIuUWOnmtoQfaRmXi7I1o52qwlmDAQzUSzNICNotPhCw
n/Vw7o9b0wvOzNZ8/esLM7W734ZQoJy2nkmqNEgYKPVt2AXVdHMIxW6u/rEd
vnwel3LLzyNghU6MqI2gF5LXrBZcphN3FYHXZKl2JntKNzaKzoKt97exhEdv
aAq+924jLToxIIw7rwqYl60bWDwa/+eQtWXEmPixK/NMDD5Kj09+i5mRil8b
BXhY09A4VO8FMiQCTe99Lofu0yzmtsbBMFnMasi89B1Prt+egHkHZRPLunWI
Y2j03LtXdQ5o3LTNip7wVI0rAgEsh8blooPSaF+Hg0mRFGGErqXHMiCY6YZJ
ZPpHNrWRSUI7AK2HFczlhq27PTi/aIl05eqlvBHuuE7gwasxxdKXCgXFPds4
d+P5v2yk73NZH555t46wV+UczOvOyAbF9KIQx3zqaYihpP8VhmIGSyVRVlLk
y2rK50zpyPGjQ7njOrxXLsoiMMl/RQz69VGG+zHGAbcG10ZdqdnXrl8nw3jg
lr1nImHbUH8dHVMLPN4YjEIl/Cf2tQsNz/BOP39toAPkwb0Ygp+AfzYA563E
jwuUYZ1/pFibMnlt1uMpyM36lxE1LpdKIxuOSzaF9kIgIXLWxTOiQB1vQj0M
gmnA0Z9XabYABTXvOXqvcPAKOP1jRhfSy6g6jriYaRsZXPDd2xfS8htjBp5b
Sgq1IXNs/VnolRS/O1bBW0/ciPG9jTWQLWuSE/wODlFukqfocigKGyhuAoAT
EAjG9ZwtV+JdfoCwkUIUY/F26VYTzybyTWaIQd/iLsXb5XnASM2zH3rRNR7p
4dRvUVh0fU1ORShFz1Qdqs6pAxjUq9bVq7NrhM6wtcrVeKoJ2ENbFUfB+M7R
pR/h7WnloqdlxwR/jUw+wxA/NVBc0ZWqwT2Z08+FsMQSQ5NT7SFAefwG4BPO
iJUbvnEfVtl0f8D9+MUhza0St5z1kLi9cBM+b2HN4wxuNtCmKo5omOBjt0q9
tqN6KiEA9Tt+e0VZ3hiXBT+4ofvV8YH6wIIlyzl6X0QjnvAtLb5e8is28Qd4
1FboZ7YcoCy+fMB1oN71szR1F6Z5u/GR6BfAg4cdQ4tarMNkk7+u43bNZHuK
+0uTfL5MQF218x+fL/+e2zinpUq6TpiDEbO9M5ZdbA7vjELxrHoKYNnvB58r
WeNsIVglKiSox+bWFELA48GHq4HrA6OhjXrThiJ18+AOfKt/a+63TDgjEsk0
C+yEZczCjvbeyravb6tVprV6TXptDsR1rJQR0XC8zAvDlsh78i127FO22ZuE
CStt+a5/MbIZ/fGzUL1o/PyLyK07ldNmwmiBsec4L+mtlOSiOL4O/O8ndYW6
fWWmebIP6mk3n7i7n/flq5ilWw/YUtD22zzBLsXXcIf7GIc93IxR5vtLqe7n
tNUPqoQalLLml4RRwV+mNTZxb++CYQKUfysSL5lXR5iHlEUIe4U6hokJJTTD
UX51Lax4H1RW1dY1s5F7FprbAmd5YHXd3dDCj3JFxFFC81mvV78CIhihVMQl
rCirdfO93Ba5qLfMYjCODUWruvAkr66ER6/lv7+yL5CiekFHJO+kbXxtCPda
IOYWf/kgfLa4IEWQZuqjEhwi3sZ8JGkucFHnXSGxE95jEIG45sc82VzWVIjj
V0DcDS3oKXfUVirKBJV1g8lBjIJEvUl1SLVFtIf3tOCF1iiJcVKbHaNt8pGp
C5NiEnI0LmCCZ9i1heJclaEAqm/BYhnOIsqc0sq3rJB+H5DMSOuIEbW1mgKL
OUoXnwl7/ujyPhRjGwY464HxEKpapp2xAj41KX0pcF8N1SLrCb5Hu/ewSHSC
jDGP+gYC67tUQ40aheaLTlhYMsJSG3bYcyb1WOMePFKKpW/YRlaL4QcbMbtO
SkTGwLYSELeUltfI+EBw/vbQad9Lia2bWtHSd74JBcQBCccl3rTUXHJi7CEN
2xdJ2m2+ejYcDcG0av3FQzvR3dWTW0nL8Hhqyda/qo3O+7gtJhn4rMFpkFsq
JHbE2eZtX3ShbbNcfqRN6AJ5dPU7K8maFTUU+KTffudIMa2atN4qRCRCeTTf
R6gcOK1QEmI7RI/j9IMVsQ0xMe1AdiwY+doVw6d/JBafXDeLwLbqv+xofqfz
NB0U46xZfgFMMOY1Dh04iCbFzfb8XXgsV3e1MUVmlMbJB8muWtA/8m3d7sOg
xbEcoWRYTf4vW+zZv5gNGh/zAAVqF5+Lp+Z+RVfs8Ypi0Uk+JOhdmfiqTnGq
haKqklGTopmmfwqT5lnvBPpjt68IMukZLXLbaDvZEp2h8wFkTvI32uSFa9Ys
PghiAevV396N829M7WNB28eRC/GFERhoImt7ebU6r0+Tl5QZ3uMyX9fR5Vyc
akiXYzamQbplq2nz2EGFbBr8GwdPMAZHvma32hhEaW8eoZn9b9/bpsONwr+g
OTrDGOgPGufMluv3ie0SW0QYOiclYp0y6rMkmpbLum4ZsIspu81nB7IwRkC1
Vo/ERnk2zxJKKw2wihPZj7KfpZu3ghJRmmCZdFPBGq8FdY7+4gYqTyKun4DD
d1lmTDlIzwiwj8zoqxY7z/6jOAqLKyRvFYaA7PA7PY77O++UxwygKbKxZLN1
TsEQJ+30dcjVuyL7wr+n8poEwCObGEorKjLeor7sgwBlZZOMXMTBkyMVCWDd
nXRoEpWkSGSS04Fbmm0d6QfoDhX3g2jOBANI+w+FpnVDpoGlTEBE/+eqBt0c
AojQQaPHVH93CI94Jh02I69rbVVB7sqTgzQxaltxg8iWCDaL0ko+/i7AkjHF
6j9vGEsB6Qus2I9tkmxZ1xOOWuXnhey1Dobl2/KZ/7l9ZRFq8B0TxtAmsUh4
RLwWQ64A+IDrvom2tFBizDFuAPAbnhVVb+Tsy7rOGtN36amOZYstwNWI8ks2
KyZp+MlQvz1LtkuX4vXSEqatwLvXhSqOrsJyGGIvrx+l3uhB8/ODaD4OeOjs
2gn15KG0tDerpAuiSgKyH3ghh001w1oxYxD267vdTKKg97xxJOmRCkBTPHKJ
9yrfBk0PEhro7eDxyd8GlDguXuz+ygfVYgFq+VUvfH0DGFg08EG7u/MTBKXJ
JagVnwXIJ6VLVUbL0HNsJPdCKpamOu0e9xEP1aWc6NdKIfrFzm60pojt76YZ
jK5njdtkpZ/QOF+wb8roy7DEM7xUYD4GPVGbvARQ+01r3t3KP4JB9QppmEMm
H/uDLUGxjjcsfEvEbVySGdA4k45Te75RZrcp1ELvXJnNfDWQno3FDA5qwNxY
BqhcimvIewCKoQWClMSfo3ogyndbQeq3R6ulC2U0FiDmcTgQhDrd5Es+Bc41
32g2JJs/vwsFQ5YspO5bJ0O4ch/AAHtgnTXzQqofNONDgE4+C5A37V6S6TnJ
cOLnM8VnEldUFaTJUyzWagVVEdo4V4G/rFK9psKqkuKOlgp+HW9/WBM8n0my
I55NQUMZVXvOlcYt4qlSX2OjL1lLZuCT/3wpPm5dtxV1cA66JgIrLN6ZJLRI
l4F2mWmOmRTrtwRTYNzKeDN+YtlkJ8WqQTIuplyZcJlvovdWjiox5G/gXQdu
2WTM5Al4PAcB/ryLGqkA4OSeDDTi7T1gJHw/Z9CSqx8dygimQpQRkwtxi1Eu
LOrt8+TQdgO0arID2ChXvgu9gqBxqnjalAsotI94Ke+Vf73VFNhqBnFvssQl
u9bRoZ2ochq2VEDa6xdXP/2SfHCWQ3kVBUjUGITCIqv/hw/o0v0WJytoqx2P
HhkP4QuXYri96vFBVi7BLozxb/KgkFRMheDB7R5Ge8AaWN47fBmfbw4kZfbf
YT3OG4zOUjqsd3tP/AaLLCznjEyrgALEu72e5WVYhZQCjgzYx0ZnvNd5OCE9
h/1LJxnMVGG+ceM+1wYMmAfaFvT9FcZGf5HL3xEUr7/OhFev1e2ThY2gxUND
aNUQC9ybHYZPLULZp3tInpWE2GvbnIN7nmcA3ZQVfCFwt7yRfCVpYLKwx9r3
qFEgwBAPE7X2Sd4PxAtqmWfndNPeFWzGezxEbAQA7PdiB7vV7ysx9/jyNctS
TbFtf3r3e/KWPsBI/3a5FJpODOhQ2wCg7vKtoT+fqYZKmXwYwgKI+/94KMpP
4MRjVEHryUEOSoIRPnHQjQdv77bxkMw0yA4vbYlW4iSLRXl5fMWyWwoeIkSC
Eh4rB5jUdinNvD2X1zNpJywt4nJtL86S7L3Vqitr2rOxqs1kyodovRHsrpnR
Afun+M4Qg+85pHeE4bqb55Us73PC59uPj/SRIvUB4tYhFSztSoT6a/g6NpoH
otm6/d5Euh3MK/UKO8FTE0SGlG7AHuPAALbyIoYQNbmCETPQK4vV/o9g+DBw
MMDNZNl0XpIQH7JnctOUqEED6h1rGfCR0TFrGgzQs/7nw9TXaMpaJPDQ0NGl
3PxcAu5CLhr9DluRmCuGzl4Tff237FU4Lam0j9ySBRaHnjLez3MFvKkmJJeZ
+aikiSxjI5uiyp3rbBzntoIc6DW129/QvSGFFXbqo3wS8PKBH6Ru7LPemNb/
2j/2n4hOCPyoSnpH3YGFWAnpF6JQG0xMAyUBEqAccgUhUZldO7uQ4uh+K2wy
B6J0+5ES6OJMV0qUTAnnFOfi+8WPSIr+bX8m4JUMLTyS76AKI3XsMFvA35r4
cW0YhpWkQwC7YuLkJZO9vTQDEb+xySLXk9BcB9KsDMGC9h0cmBk0O6PXO81L
whp7zX5HdkBANxe/uG35tNFHpMeHaYSqwUv7D4lB7FtaOFUM/G+zU8OMMdWH
Vj7hdj9DR5/RhMffurAM+dDaxiMMYSQ9SeLMoXc8rDy3ofAKc+jq2bRQLfh5
SeVIvof4EYFUCmGp0UCrGx3bRtM1b1iltTESEfOAnwNZ2LsST78hNJaewalB
430rRmCoe2XrKW+0orPz8Hho1gdr+p6o1IUydT55pyVO9Mg8w6G426fH9fr5
WPC0W683/QdGy51KE7s2QIsO+9ZiR2+W2iN0LVCfPNwa3YffaqFkh/UezHWD
QEokGJ82GLJybURyAjEnSocNelhjnWup+DFh9RP7vaFG14azAwyoFfa5aKrH
MHtzDvtJafCahbRcBZ5UXOLDo3kwUlZTz5mp1AkQY0CtC8uinMsJxJ1cDoIE
Qly+o48VAukBzSJegEhUoFltkHKooxP7w3FDAk05+SbH9rPYvOh1Oy46nklZ
PQKIOKG0kuaZx/sgZFTYAFgF1h3KkiBciGiCqFT1QYLUQFvPUCHI5gEvXJ08
nMZK8111T4ArBCrTy+QRMr1NBRVllHlUrZwTlIRD1/a3t91NcO58sTDnrEP1
uOPCAtoad8dy33z1yAb2QxwpNGjvETw1f+7oYShsBNO/d4LMbjdfAVKbMw3/
GvB+oMzdsTuBkIzTQk4sRPAr/zL9w3Q5R/MhjH78uzpIRensXCegk/9ihxFz
artspJh8Aau6C0LCkhxj+u15FNIETTo5cgsLDuti6ayOCwqq8EM0OqcwLJ4q
B+7+Qw9+j9ubMpuKdMi9KMyNAj7Xohq7I8a5cYbny6w9PFcOsDbrMosx7emN
TyFZAHalAU/QQlM7PdkJ+DRKfk2uMHRbaQy2efgWB8CGsoJd1m24tXCKZbWM
rB9nZinhf+i4IyqLMNQk0d5DFFqkH5aR6rbzquRTGIXLARcR0euj/O+Z/lcJ
Ah+AFlm7mS8zIwB2hKvVuHht40YAj7Wnv6dMSqWylbCs60w9bdrNmvcpRNHp
EjRfE22izb/UgXNy5hzzHywJIexiAM++4MPWlHIJVyciA3ufKwvxZ0hJA5Dp
8A8XDHJI1D0NQGPMcXlagflFV4Tdqz9rf4x0dnNL4rqxmJemL0hTeafaMGC3
4A4DJ0MwUOjcMb7rGFA6GgIjRuZFWMX2f+iowHJc5Plj0Ssa8SqxcOFdNrxc
+BLl5gd7SrqLxenuD7nE2f3mDwqAP5ZJGyCBFheGiSbnjYQXDvUA9tNAeQ7F
+AgezziGnUbdwQDUZNDFhagAysjwxa9aBOOin0IVziKYgsb2Cn10MNkrcNdy
sqAA39LjJ8FKxcV/l0EN1s/BJYO8SaJt5JTNaPn7QxjaB2Bat5aN1pGLPf1d
vX0hE2WZbTqhOKrHRHiJ5K5fHNKkatHe+jFMWbp90Ha3k8mdM8jjm+lwthMp
1JTaxdqYj1lITw3JPqBzxLDpNkb53cjMPOYVWy/Em1VR7HYABlnXSaCgT73X
1sOqvP5RU/n/zyjC5AEvYxGfVPk/NZ0ESfd+wYpokMi8sK5/oTNw3AQGFEQA
rU6y+yR6iUGAK95hVyXjLWwTIvl11faj/+vfbskWhBE1fVDTUiROs6DEk7oT
9VceJR3e8V1E6Xvq3VF5UDzqhlgHPiDuC4V5MbKMT2rm9O9j9Ua8XodXaUUc
hvucfY7ooC3tR1phcG1QILf6MSmDoNFRuCt5bd6bYiL5fV/pL9vz0UjPF4Vq
MgVuQOyEwe0Mzi3ryipJqznWsuxCpFc4C391o0L6lOMQ6ktsNAzRE3qNHDZM
BAbABAJuL2QDUig22RwteTX7PvJb3FuQfRy5TGAiMu+jIirCzxuVeav13lrW
nzt37f9ishOQioMYZDy8P8RagC+PSwlwiHEVul4qGhSrUfQcCoO2h3BKKMf3
PtWvApGxaiRK5VyXBWPShpWGMuMUmYrZVnwbxrPemGF7HKD6W30nS516HLLN
hOVLZSN/3RW9FQPtetFb00tXIo0lifRlEMAMoW52m5no9+1By9wpXpFfiT0Q
S5DVQl8CRUBHD/WB1cEUDKoxY7kFNsUbPhSvHDaVoRebDv40v39JJwt/M/OF
72mhkTNqKgyAZvtqBX8ZgWNDaj8z/vA8qk1jXcczOI+65i1AHU9iQT02hRdw
xf//jzMNpl08rLBiihGxYXV6sAdjJ2Dp8zffc15EWAvB8o9/QPSc9p8sMhFv
xzO9EuqE7A+a3nlwtVX3Bz11W9NLYpOQLmH4kfhOVZAAB7v4ZIXxTjgcywCb
HPbrk2PlXolsLsfKDLMS75YDKW9wd0XdcvSfEOdyZ2FgOXOhrariWD8yoQg6
Nu8yMrEc/seHMsVtYazAUDTHRitibzht9kxUinF8tBbY3E9iBGD2ahLmflJd
U0o/YKNZ45MxqKF6flH7Qx1jlgvvcDh9Gf2pkzDKZNaqaM2fjZLsVwZ7JPzM
FQ5cBJ8XnX/BJ2PMTKUlREzzp5PU0GdP3xTPxaU5rgMthVGmlfkCj3w+7UJq
e7IxdORORHy/mxIlTEZZr76KfujZYLgn9VHkvHddkakEszRMAB8/HcXbXJ1p
ZCseDzHybGuc+uJZDDI1wbOeF5Bp0msnxVLjf6z/5ZKPRCCbVf955METyY2J
U0KmErVeHf8wZLmMQrptIxNZeSwB61Q2BI3tsYbYWBOCR4v6khohpfj/kP9/
CaMQKv3O6kEvpvKcT1cChMWMrcMdFAfN7B9ga/+Zj0Byhe/1lRM6viaBs4y+
xigTbGRB8ukp+xIHjT+McqFMpQZePPmZyiKZDzylck65jcdNyzCsL7Kamofp
HvkhWRPqxWqL5dJ43FizUNTeJgOjXjbTRpMOUKGol+jTuGt9H0xbhmEOnC3t
iAU02De7fzRYNZrnmgl0v5wwkwziovsb4+MhuqT+ofBfyGyS7ZYftTfBIvjz
zGmVmzWc8V6juLyJ9EdhHcGa1xJucosL4x7ITLB69t7+h0mJvn6TLs5aQd/t
IMSwonyEZQ+x7FmmaY4i6yx15vukvQ2OzRGKs4ezLBl9l62RIoFRbne/7Cou
H3TWl6+uxDE0krYT7RpDfT7shPc6sr6lYOXk6dUw4XxZyv4yyT4DEZoJg7GO
jWo21KkbQvi21P8KmrNtO4EauUHzbkk4OrHMsGfPncdOe37ucNuS01BxU/H/
tbV5bC8RF0z3Nu11SkG5dhWYdkk+sqdKqvRYZUDhawEUnBbGuUw6alUnBdVk
nX0vzmBnp/uTpK5xl8kBJ00LsIu07UXnhhzBCJYoRROq+H5+b9s6/J1lWyyn
f+f2/BMjsNL5Ktpf0mJIt0AOW5r65AAHivT5UkrpjvSNwefblodDAK8Z8i3F
v7u1K5FzD7p4D11aOMEfbu7NbvpnWvX66xZuJ7WYgArZ3bI6et0WJkJEKd8Q
f+6u4dvUi6Ib7lXcKQi5B4ZEycEvrZx2UNxgQ4kVn1IYEX5kwRyUZb75leYL
AHRb1YLNHfH0XpYJ8yewGO2CPhTvTWUU2xrj5BDUVcqvxoBQjOHlKPNpVMEa
cEiAqxyEc+NSqGR2AT0D0hr/cjcEEM6qANchR7pH9LSku32ISEUo6cLyiu3P
ymDyRdbU22tmEsAygNU9U5If2Z1RBJkz/VP7yOW2QLyxe3uvlQHsVr8rk7fm
ZfSPJ2x5+LSeDxaNd+uLE0r0YniPj7wUIA37uZv6M7c0XtOGYcJKPDBrVNIg
SvnT9j+Au30zxqt6tQAjPgCbDCvwn6LAdkLz3vbmkPsr6AesLCDKHvNN0f9l
NBpkL/3X0FXFRotkY3CbcaDDoVQL2W952tBoWXefcISgQvue/EshO/G7YeWJ
1YEQfx7IaKkwVD52dzl1SKrYie+c8dvMZoBNZJ2OVlwhpZR0rt2SSoS61KA7
B5PlOfTJ4T6RSYZOxQMdhWZXlQhS2L/nzCbtwchBUp7loH/tFUp+YuZQ+7dD
JfXuMzh+Eg61YdiDnTtu8SpmMGx0fG3+SNrtH9sjdYDm7Z918zgy0lyr4Oox
moot23401hneBe1OWjv9WtEOFzf3KEbX0T9LKcXx8TrQTu8kf9DFfmMpBoqS
nZN2cMTArMpjeomy3NnqQuj+hrVDS+kSk6tWwsbEyTWZ24OJYnHp+NE5EUNy
0SRghr0GvaS/JrF4zFBZ7wNk4ozdT9pvIv4skhBbdeSpD4AH89t4NUxTaN16
BbdDEKdAqhALUfOs8r3cX2aJRahFVkdFbOYOAwIu3hZ+TF1gO3B67JqoI4Xh
BYaJ60vQXHJioF4yTvnwu9csYXyA7Ul+DHGwoulilCq4bg8slJnO/+/yveeu
GY1WoZXniIqFt46wCfKZJmpK5fMSY6Y0cjtb759EI6oXZ/6jyI7GTFtL2VF6
VNwnvjbJ3mC/yAacnWJaRSBL2hSzH/mc1NIF3GYrGvEQIDlAtgVBC9HlduNn
JYXsoeQD60HhXddDgrbNpLLs+Jy1Rz8XMnWtJpCf7UCSv+b9+rtU+zldhvW7
13boE7dmbYKME4KEM0qz11Pr+tm34hNEI+dNcgRTD4jzd+yFn4Wbr7aY/q0Y
LJzwTCavZmZvtTApOm6R+xBKrI5/xBJiKx2ZK+HWVDWMQ8Lh5+4UbMkS/HtV
1Tg6qE9kWVA97d1AdhkxzGayeinrkVX1loFtEHr6pZjEudKX+FKcJ+F0BUxI
fAZPhcRwMobIuCIT24EVQYMiXYX5yLYBthji1VYZHwltwSMqp9fPCdJPfVcE
WZm/CkL0/QuLHuX2xThOv9U2aeZ3GVhR6EFsOoHKQ6n/cTdQyrX0VtTz0OZ4
eL7LD53zn9Ao+MU81bkWv/8SWBjr2zcqR5EipX1QxULSacGjmtzY47IEXRIT
3mDX8ATqSTYNNrRrPxp6f5w/LoGcIHTM4ON/b1Qd9uWHjMEX2VXk2CdclLnW
HhHUKH5dxxeSAQJ/xHyCRNjFpcemggQ21bWuuhYPCgvxU+krxGM9h8bLv/qJ
WCxcr/79vOt9YqFy2oyd5INLs++CpNzcbYgIXQ7x955hqp3JC5WSbM3lYte2
5l9gYOEW2rFmLUTpFoeQI3FMKcDokJnu40hRr/GiXA3A9+xbJFvRaOtjm4wi
Kx0crrSMRqnzt03bp4a5hGvtXRfEAs9C+y+dFxaiTySSs+Gy3Llw17Ib32/O
v1f2pq8y/JX0cJWIZYcWeu4ImLiQOeQ5sk6opYI9hMUgYLZ8a9IcZCsuYP/j
weUwDmGvLzTo41SQmagYR/sr/gc81RC0xQgLdgIcP1BzjDaQk2GKxFfp1E6P
VUXEIntzKnyMZl+WGFb/tl8m4Wj5lKOm0uoI/OFADXnKGq8/eqKIYtAcqSp0
Xy//2K1ZBGEMF3NfNQx1DljuCTZNnSViI9VKouo/mbJkiQLmAnzpRLlU+i6m
ORm6AlK9s3Lrjc2YWUYvsJOxlaTx//rOWCWhMrNygx2Chex/jxD875tlBSxA
x1z0PjpwLGxGJ9Z0IiW10ZJ64fK2J2RjpST6O9/Tlkh2aDBS5zNW0MYMHfLw
hoCR4dx8bc1ZbcTMQT/6Ae4GOLKmkZUVT/xuYD6GU1dCFzGpsPOheJoTSNlj
hCPdffqzwWq2fCXt65aelFV1syIb0xZEKct4iY9VJ4paxUN6FgmHq5DTF8XD
IkoSNuB3PceZIQN941Vk5MBkql5nBvVtNRY9+1bIE5RkV70N6ntBR1g8lUB1
O3CEp90KSNO0DdyUVWgHPuwUiOWGlfNgI/cTtXg9P0G3NNLr87wLgYyfNMGj
I7jMVDIX/j4IQDcY0sxepW+wwqedxgNtcuON14iKk4TMLoONRyqV4Gmg/dPc
WItR/oL2a1R2SHVgGIsb7OgmkvFXgVinF0xtUTI/kMytgzRZ6OTZQTnRiwxf
x1Qf0QLbBXRLSSHoyIvEZboeA1Fmyz2wS35zC3wmgCr6fNX4GnS/off2Vp+W
HsGB6hREaQpXfJaT4hYaqbX0J8qhV++dtvE8luNQZetL7hekMVYeo/GAPmg8
Ok4QtJf6vRQwLuiAPhUYEEMx4Wf8stnY/ffnVisd+vsIrxImMmiHedc9CdwI
fONl/thIJ2tt0Gf7DqYBR0W9wnPEURefF09Zoe28odMj7VMIAbRW/UueAY6k
BIsL/vIcw9ekGlzR04bIbc0rNN2D9SkHjNe5q7VGQTwCyvPgxqfJywAqfMGs
uS11BtXRSO7iWrOUyBcLCMJoRJLbK4QL68i0FNZWcOkTnWGq7Vg6SmZFzi7/
xxXt7jps+zP44oTQWQFGAWfZbfVXoM2gDk/si2TkeeHuBEsMAQtnfJcmdfI1
jMGyft8fwHUc5jy4llS43nhA0lEsvPklmizER6pMCRjW71HoUUq17DKf/hMu
8+TUO7inA5xp0OTR/rxOotrbzzApPt8KvvgnAYKTTYrgfUqIZYrLpIM1/SOW
zwTs3rvY4BMsDDodUkdMebGWYiVSml8KKH/QwMSZNdxClTG+Ma+l+jke0K/o
D2GorYWldJzCnriInWY0ihdIdA9/CRgVcRutGie4zXZjTdOTjj+PXHyV8ePX
siRX2UZ5OtafWOIN3Tj7mLQGIcuxpDs7sse2Gv7jWLFxHzUweRsTtVLFM2sZ
3An+LwmkdHal5Mdk8R7yX6gtT5tloF38BUryTSFQ/7L0SE655RCMZR0PkFGa
sFmv1z7Cl4DOhx6iW5jtnHCEV+NPVLCFmkoKc0M0i5zeJy55MKJb8T2nyMOr
2xsaPn3i4kvuUnb9ezNjpT4g+mU1m0sSjP4fBhuKiXUQUXg6l4LfCajUDavU
uKFj0XZbdiwsrDR5PJlySI/xoiqeXlJAwyXtGOJDJTWEoTuiAd0ZTJfs+vO4
n3oeUf9m55GdqRZ6iIA9LpwX9Gt3rfnptz/legCJvHf9oFRqyDYSDLm5AQZ2
AY0AME/QHTkPh7qXvbqDrdI3ml6leHtrZ2/a/ZJJ0ReIVVnN2YA8EQCTbSPr
xjeXX7hLVbOAmY1xBTUj0l1APlxZASsKQE7FSFA340gvzqOo4ngnTtMajG+4
P78JVbiK2Nn6GMAPVCihjW7v2tqzLNhlUM/O10u55FBFsdZW8qzSXzfQ7j9J
T+2UXErhTMr6RIsHrB4dwB7babXGZaCJ8JvG+xCnpfOLeg6kBjqSVP3Ow+aA
frsP9U+wbxbUBO7raryKvPb7tEgq04DheWhK1/hswGa8+416sAAx+zP5wNS0
x3crAiEqr3tfAzUew/G9qvmJb7lsqShpbnB8ZCS+jHJUcp1cWR6IS1KhqHlW
EFcxeuCdrhqU+hrITdSHAhKFFKOgn2+nbGKNU9kqmvB6j4M0mbcdA1+9MTmp
eXihVpEGhvdpytbEa9shVwK1C6WsoX+7Qt+2OS4++074Z0deYGnvRlvr8oOK
cCyWz7KmPXvWKgY4AR+yGF6cZr8swLYwpCL98eYnzZegL98w5AclxVoKMHjj
5orknNq9pzcyt4AvUM0vYvGjDUKTN8bs62Tolbtwvj1uN/dmtFc8Od9l4U2t
7XBGIeCNIkkKPBkm9tTunPEZ+ngGVhjfQcK3DbuBzL8z9p+wjx/D3YDPglCc
0OTT423PBobfmGlrzi1yv7av6Ir1JmRH7OG8ocxO/u0yJGT9+5QR8X3/YUJo
E3vFcBE/ClaJsk4K6XUEr58igvCywaW6Rc4Fwi2wA5bsIjb1OM8XClsT9Yzr
fe2JJ4ydmLzSyItFfqxSQlQ11o28Q1hfby0NyJvQYMlMaQmKisRx84ufAHcO
T3mLuOXCEgsEc8/bl15QljYZM++PL42uRI1yh8D5OgPCowN6VRMVNHjPyM35
AiEm7rLMrQtJjSzy0asTxT1qgGwzwNxtpIrCW9zH0oCbSVt/z+p/IFZVLf9k
aGnpkyB5Xqkjy0t0VAKh7HVQBty2jrkaOPbleJu3R1gOcu6a8vpRLNc75/rR
SiJSC98odcHgGZcQxWLhacnGAxKs26EnKF5mPVcZFOcTPBIucbH2X1ryCsYN
lLYvPksFnybRNAEjJvRZZpGsNQIWEPZLDENK1d9Suw4CGBfo0WdzSqvEKDG4
oNsB1gCRUzStLY/TNovg8HGkUzdgQ7whQiJD24ozOjxw5oBS8AjUIEKV/uM7
J7VXks+sPBUFv2KjdlilxIiwiGAeH8XbW0v0ByD8SJ35RH3e5p2C2n2h8LCm
rCLt1ixTNPJ4S3jWOUXi8Rr0U3OLSHJltJGAogeksthgQJOby6JGzN3MFXH8
u1NhfUWoXpkLfgzxW9WD7JIwrq3J9IrqZ9vbryAaxcovZns5l0ArIXvuFoU0
qEKTbAxjGUAkrpeQPfZOoq5VoSBD6aEmtxzhsg2K2nbTXO6/Fbmq5uFWZEVl
HPuSVV0qawHFfE+EtFpDNMOjQgzA39HgeCvAmZmHeCOWUJlNhLOviqJfb1d7
QF8R7I++A6lGA0Hz95FsFK4c3Jh0MgZtKlRoZoQZzGh4yk3f90FoLp7fMb2r
GO2WbnxuLaqUfBTeC/Wg6O3QQhMftwSWVdqklSSUxMXlyunUswcvklSEE10s
PqB327c/Ge3FhHT7HgbFH703XR9MdqNHIc8m6ooeABuRP24hDHmxrdxDcUER
7KIbpaGdSmAVsrQ4v/bSpKlmldnLSL4YZm6KFNDxP69/mMWHIaxVfCJYYpJ6
QfjuyfJrrNQBWlp8AntBxaFoCPz4y8zH+YJ3ZcVZeXlGYcUSOudBgUY5MFmE
6a3AZEZWuSRzvxIalssn71IjyH2XjUMXjNc0JSfUDxB+ZNGyTT0YdeN1NmPw
lZpazPQktCjwk6FrNYN8DuFVEx+czCdt0IKX/WDXK2tADL/R6yGECZwkd8xV
1WgdjFDLoTYNRl/Us4XZlA2Sr8jhmV5FYY5/Zgc4D4BOmVC1AT3jf7jSVcMG
DwW3ZiqyLbfHRacQBbyPP696/CpOTNwoSTtw8leVGN1A0PKgkTokH8s0DuQj
ywFuNYgmYBiEcTATeiNI67O2FKPqaMBb6q/6/xNO7+NivB1WDKvf5EjTKHDp
P0I8QfJY07Jt2ojbP5vmS2zE/erUByyYAtS1FBeg+gFnWCphRq7O7zyi3GCP
Q1ukSlYYS381/jF3dZriLKwKdnQF6ZBODPmb59xGolQT5AUX3eykeJbk/Yro
M8pmUeFkCuXNmIRpOwAEN9EH40+DZ7f8WwW1S4OQnlB6AubU59KpkYqmV/v6
0qA4OVAt+Y9ZiQe9V33P5ePcsAaD12lxIj1bw81GrFpwxnfXSfa0IYehNmu7
OLHgb769ZPaEjQsiI4mMEnmDsYHeQ/TbjYLpvmwWo2oKKVmxxaXq/auIfxfI
xTd15eZ2kO2jaOCthmdNQuJolUYLAO2vlpAUL/Qg38Q2497USGskvmlIqT8c
jXw5Dx+/pahfj8klpEH9O8t1ql+3whcxn1sCgbvjIGTuSt/3Uh5ruhVEuiol
JB8SG6JR+eORzA2Ipn8JkzmLhMFJIsYrSk0kNr15KMccBfdB+zifnzZQrPV7
x1hDbs81MKlrpjKALOUioI0Sjqrnn1CJ98VQW9n1/znmmhQ0R8XLYAz2fu3b
WiODoGtSeKhDkBPfPrw67FGv3G2l8qa7i81n2xbO5aTdaOrrkSJ+VrWMxup/
uFc1YPkZXWdfrrZba78P9DhGtGyydrrk0yoLj3w4PM4E6PoVsRdhkfPduWiA
7eFQpntLSr4eOnIFXLXNyYS7DzyAKThJjc/6UKZCAwG4n+OOb9zUohBFJXGV
5MRNxJAp7SdbdVkKOuqgcxavyzw1C0PHL9FblMCI8IieqQv5PXsrHrAygGdi
0AvNj+bvXaYx6GfcwPP6CqeOppu7mydWyK44+oN/iaLFwuETO8ANs7sjnnoN
gaHDS4kq7FpgxtPHAu+IyVXyf3qxM0HOQI77lLktoLuj3LZ9as7okalHdbi+
kP3J/nFJOa0C0F+ewLMOmLyyZsnoCeGLGPvzYCAtbVb6AU72ehzPpwsgh0PD
eG2uQD4WmvwJ2ZEGxxFEnfTWuZbk820a27SltMDdAchGOnaRsqtqZKvMcjDV
qXzC1L9FptAdcJQo0IYuu+3Efi484U3a8sAwvkPUoc8cbEOL8FmiWFyQyi32
A7zdn4XziJDaThkhVkRbZ9HFsupLNJf8v1c+RWSOa4HQWgmoHIBUI0/8a9AA
mbrMnTgKZlftuu/lq4mDeKvJCU8KponofXz2Um4DRp+QqMlznzgy8Pg//uLt
QG29OROm5lXpohX6TH+W6s1nY9ELJsWS3buLf5L8imI+5CzyL1pTb8iLL8qI
6E+A61TMf3feWxkHGmku+4UqMxjKJlZjLMVdg7mtLFO0u7vY2pctS2I0vAV7
iEeCWh6mA5SRvrd74qef/QGiB25wEH2aYbt0/F+/593t/Cw0gKDzEnGVPcq7
W/RLtwUg20SKhRSQhfNgzgi2UhNf14zBHq2jcVZOe9TlaRZ3xYGuGHUh4gq3
umfEGra2jvql//cK6pjKd5x4eP0W4vC4vQahALTn4DfHw8sBsi+Q2U0lMVI2
xuxY/jH2+X+HaqfBZr2FDrQ2Pngr3fjaNmGe3/tD7mYBCNUL8wCwIRS1dLLl
/O/6msuyicMQS1O355TLmD8HHmSPOJ1jg77ljxMelKNZvzj5/zrIZps8NEYB
aclwEhLjTjDeTmzrFZNBu6+c1TVX28g5R4oAbWbOviDLcRCwX8E8B+uUZdKi
7ODjyNA1XlmbgZx6SZyzOQr8aPbr1tQRsewCtOrguuRfI9x9o390jyD6UUBC
EIb0phEZ9MjWh+f3m1qtHsLE/ppatEA9TfXPDdZC96OVY/x7J032sYD2eCiD
F8tHzPKUdJmn7vO5BEohQg8ErlJ3fTp3uPUOUnZmYaV85zFW5wPWbe4/1z74
T/dBNymac8y0JxfrAoexn5p9Z74Dmv0V2ZMQ+XUEfdVIUOvmf0S86465qjhy
omvi7awdMg7Iha61MSESZDMIeHOcqm7exMDhMi1JMVxW8v9MP3RJBfSdeCBo
/0tppDEXP6YjzdpHaSqe4Z1xqy7eyRyFcgXCG1ZhKlmSQ6LYFeCGrG9+DN1V
7c5O+ZmcnAn/cY1ybREjJYboCslsOGgfVlDK7Fmbm0f1xXyyHRDe3bGtVcgu
2l3v+TgkTJh+maRDHeMMYiNSviM95Hlj3lJtVvIqPZhuntp0zE984W3MMocS
QWJLUjDKcb8Pr86xhuyoSJcePP25bKrUeWysvlVU5Mg5WA5hdX7YubhGrnvH
qavVkjG52ic6SqhFZVUqFYSU+IdEUQtKJz5LX+WySYoGmJLpfudmBDZgbRIf
hWSFso+brKD0PeLVXzN8wN2PCXll8y4zkpBZmPFZ+LkF9LHZfFYTSUrXtPyj
HnSmKCdkyfdGzmSxI5kKPgGimh/71eQgGpB14qeuSA3cjQJF+3EWc/25A19C
rEfNZ6SuSeB+NsE8uAbSiSlWVeOwYs8xGze9wWs5kz8trI2QD+KV6x5wAZVB
9N6KVOB58TmT7Iomd4u0h3OMIWGV1z8M7Zw7ezAQw9Dlk87BSZc1pkJIttCq
A9B8bucvJ6FIOhN3fKIK0w/DlojLbJXmtG2SHjoX7eP68WHDFCXMAFeEQK8p
KlP0OgR3NC1+0kwNRhp5puXfIXCPmWE5PRuHtFOoE/BRKPPBE4mRs3Sy9m6k
N4FBjP1X5VQ+36ubf3RXN+fpij4iIIb7gTNXIdDt2cHz91hEO0cKq2GCbWVz
39VvjnjpD27Nu6cyILs6nrKp5I9ZMyigNYHtahmiXFo6VKAg5cFAR8u41V6s
SRY0YbfHwlxyPAJFZs6bFkdsdElouASF+S2cP9qtLiRiaPcHQyiWsSrHdS3O
spPbVqhSN97G8GuIApQISO1BV0z8593jk3lTqhoFHRznYIkEqUazTqZKWUrk
X9DSNyJYZSGVTL68YUnE72D94jrJNg4c2HNktXEXIWEeY0+AR1JmSty9+0oZ
UtK+2smf0oQnlu/X7994Lz2pIFlmWeo3KI+5v60zqhOaL+CtcQZrsxM0RX4B
qJomZpeiwK1dYgpa/jDIVvZAUqx3ATwee8V3k9Hc7Ag8+oFmxPgOfsyo7ueU
1pqUrkZTP4pXTdAFFB0Ro64EoUt3TMNLIHVgeJf0s12fYkXwPSPY5MspPAxy
/RnVT9Q6IpsFdytbFwHU24w5tH0hL8yIWylxNXT+Azt734PHCnbMkUCmWIj7
9Q4xn4z16x2/+mCFpi0eAE4bHVyRB+3JXiJi537E7pfQQ6PQhwNKbYScW957
7Y3DEw6rnuono1SLeMt0woaFdL+TRaOFlbUFFATUgUhkUs4gz/IYlFzSzqaD
kMPaJbRJLZbrxqY2UG6bhaJodBSj6wG4agBr87U3rV+0UvbiC9aIWe7qSAPA
RNkMOaUwcs+kPq7fAlXna1xgaZm2z6ghiIOr5YH3MZqDRTnMtVLSq9IA+o4m
r/v2LzDwSkeCtGMn6h7xJ+kJdowLuH+EjIMUTmVAv2dOh+cLNoQ0R8AzKdul
lG52e1xaz72WwYhBMw9xolDEAT2LDEn05kSiK/XC75XBWJYKW3xCqHjGPLW1
8rG6bOO9l3GhqpkhpyffKx7qvSnWOKapo5xfzSOLJsfXNJKCdofrstyw9YpI
vQsso+WQfAjmF0wKaOUOcs3Lkh22WZ+T3v4hh74GCf8uQvJ/syoFtaYA34wa
nD/v+iwOA/V3nBiMfAAdJCD3EnXrAbUQyEdcoWb7pP5HWUEwHGcoCAqP62k3
pYlcPHgCD1+Up24fKjEHeIYKJBlf6J2YdrQRXYvDHpIGIugu+nUwovZFFMlo
riIPfoUFiL4UWr7fiAfAKxru92RiP5HrCwIxq5PZoyAxPR8AdJye4lunATz/
dmdZD4lBkqc0w35hGiGeDpIY9kLQyUAI4xDqJws0ZRpH/iVKN2+ec1mObsGM
T0AGiofIU5D/l11eqx2fxlxWeOsiIOgsr1WhmHUTCq07QgvlsUxwnL9QRYja
54hNdjuY8tRXSD+EG4Pnngjw0DcHWr6UMzwQ0GWPHHxvbP79ZVtwbY8FiV1t
3TrbVz1kd7xHETMEYBQ/mU8qjyIE4EOQ/RvGrQyNc7CREzFeWr6fIYiWPup0
y3Xh8T9gwFyeL0aeZcxpLT/Y2f9it4wgwOdPQBWrzJAgoHxoFjStDZnLcL7j
5T4ANnXLcGu6ajG0WxZE/n2zWI4w2/H4sCW9DBavlz1AXjdXsqF4SmdB71RG
lDKxc34UEpJcJLOVuxCsaRzCDhEzXmAqw26+vpSpPaKvgbvb5rSG8HniJXGj
0WGz1FxCYXaSFouupyIJkptOAcaWz5YwCcEb99NUyjsDvmhskUmoiQ0GCTZO
f/dywpx84dN5GaMFbg8ffIt8poAo3CjR5v8t6L9ah9YHP5or6dZT+2wCdXvx
8U68ZnCt26I4Qncnr3JOYKSLUOILZrUoQ64fWCSqzy/GFG22bTsPwLnOPEXL
bekIjVzxWtpwT60Sedd1C4YlDcUcb6K+9+BCXK+1DgO+XQL9h+nP2ewAig4G
D7tEtOjV0tMSnHUV4MOwDnBp2ke/UGGZK2nD0AKZ0/AswvKwkKd6lWUXUiKy
pv5ObxE3ZoTkA+1KkiZqbACauskWGoWIiLXLDzVBGjw9L6mOdaoR8VuaN0ZN
I4TSDXGgb6/EwaP3ofTkx6WW9aMjloYqSWiJJ+CnFJLd2SHsuwiQBIFTfMWn
V+MjMGD80T2JIRux9ncO+oA5PoWtN1mhb5LPnnV2eZ6GE+0b15QPtvGfbijC
ohoiIShxZmgho8ChlcA+2dcnB+jv8VVjQE5dSszMl++AE4XKlpLCRod6K5iu
D9X6ovpoXQYBDL25i9rIX4+onbwXrjS0Ys/j8ysL2aNiZtqUuLbwK2w79SlO
0pWMhS+2Bciyz2Tv6kF8ieY6F9hagQ587pyd8ae3wCGogUahwyoYVKwLtTU+
MdnSplDz57ATS9BlVjJtol3Vq1howfqkrbDFIhLrmW/bj9G8qg5JjQZ+/nht
BA6yCPoTO2R4t7eCbu0vQKaQNFAWyVuM3Ijul7eNqLiKJUCWlX1vrjumYaKi
yA/HdysMd+W20Lc0Q+99mVMSjPRG795QJCp35XZXv+y0iDmhWcomMLkEyyi/
MLLI+moG7upDYnijh4D8eAfF4y6merGdG1Pasl9bbGwVkV7uGfSoJeXttYur
otFaEPTf4cys7YYPfLrAx0crmG4iDfLFUz5x/czVwRKcWEEwiPOpFDYQTFNN
9gegvolbDXzUKdoqM9UXjLJQu7r2VgIu9qWV0PCYt88xXCVoQQlfBI6PABY+
o0/b3FO7ZjaTQICYClUberFzYfablhV3Eb8va1XB0Zx2XJmuzeUJKlo2/deS
D6P68OadLzcz2WKuD4DWRrdZxFvTBN42CBFVYUOJdjL6Rl1j+w4gq/bHAmFU
auwYf9xHHb1PGcfdFhFw9uWisZlQFiVrrJeojlIn9J8eJ/qxX8SeBWXNkUr7
hIakA5HN6hIcrHumzfYWU7PPIcEwrVlOLWIH9CGz207L9I8Yg/dLQZLFOzWE
ny1bO9mdmChBT1kt8bizNZL0gGcpbDmTtxUEUMRNFUbY1TNGjdNL4KKYlmP6
xqrYyGmOHzrqgGoWoI1I1KHIvNF5pxnn5U4o36c2vEy0+8YVxccNatBil2vb
r9+ZpMu8oVgd6cWJjzqdKUaFCfbQr6cavuQmw7pmRENkA2mr4AhlaAYRsp4H
fnLzvkdQ73VnuHrNXkzzj/u88QMRd6QpBnnPaaZ5yXyr1QmwS9CWfuxz3pTL
gw0T6DJ0ND/lODc1U4fSc8fmsnDsgz2uRYtwVb9slzTwY3jwny+md6YqY5qK
GErLuYZ14CwNAqeKriiTTy13ZdwuE3lbtSJ+KOiWidm6ruNGnOdlqe+eQH35
6P3o1Tw6oBxEIIRrfPl+Yp0hMPXKQgJ5B77fr/atRSyo+8Q+ulBrO1+NS5rD
wAZiVxnj456T/lP/KB2h4IGi9PoQ3PaCREAX7XPUDQFg+Vt35vB6qyyW9TW+
CJ0C1PlKDRLLkxt2xC/SSEU4yBBuDm2kBTeALxBDJNvkp5yNXKcx/hT473xf
av8lhikDk1s1K8X7bvqs1EaXC3RJCYKet/OUshRQWjJag2KenRbtMn84U9Ws
1n+oL05ynS18AnSDfLEiWhG9j22R1dqQtp0CU6vZ7nfb1+p3D/yg+dNQEPeL
UP/CwdQQSkX4Jd7GNzlg8ZIy2vH90pXl281ma/kJpQlUG/hYd5kKOBrCFT6U
nVx+R1i6F7gjZ6K/VxR/hMMACC8boLpWzoVcK/LDjP1csTerJLZmSS7jyPm1
dSzP8vSP6qe/L7JWozDoUZeIWRSGvvoOPSEL1BO8T7tbVsojjnfFAX0jPItu
YbEbc21rYVUukDtn551qy0K27cUbjoudvEo8M/Dmdp9pxhYUahuaOFq/sWd3
QhquXLZV8t9DPxEaZFf+sVQdiQYRdrdWS6aGw/2VjRLBCz2jCY6kY/AaNvNT
QuFJC/4Sa04abaz6yXad2Xu38NT6NztQuxXQ0sarFr8F0X39UZduOWKquEkb
SvZg7V0Y0FTLQJ1CfJfint7Pxd6K4t6U5LWnR2cy5ZtCCFQJiA5e2ZBRVeug
jqsJxgc6KhYPdCcRle0gOJ+vl9CwOabnFIxwUWBxWiq8yixfw1B3mCTfZPSQ
2mEdEDbpAdCmSQtrsQudnnfZdV2PzVB+sDrbdW6OKjJt6ng/gBthUDuEBXkN
sryYfyO7hWebNryB0+/FS22/XkHfFXAdbmtJpFZfbO1Fovxw3jbqolPHbeJQ
OXnKCn0L/Bz/VasDr6TcxajB23f+CqdbdMt750ILJXT7xCaIMeIUUpAhLx0X
/kdQ9Lo6CmvUZgJT3l/ao/KHJrvgiyQpt8U+CZ7B5c4zCS09Fj8/nHMIdxcI
FOHuJZdREWC65D0mKUKPvNa8Q3EBYNMG8tMKt/3jCu48qfUe2FQPSJPHJnW2
z1T+7TkRHOZGrG2L/tbf1g0MkPRU3tIbazxZIoO0DoMjlLPj1KtQAcaGUrBl
vTEyx/QGQvF+a3OUc1KepMy72xfNa5veM05yFrQQz+Z/k/g+/pWaK0egcQ63
WnVgkmHwvbM/156lUqgPlbv7LdEYOTidszeLlSLonDqXurfO5Zkesq1GCNHX
2v1E3vy81/Vt4cheXmEu8XfDpnfVdqkiVKSdgYuS3KPnifidpN+GtgIeYjd7
LMRIYyNCMAG2BzevJuO6SBl9Z/VS6qsIVivGguURj8S9XeM/V7yOLBQTyakE
gLJCAil1IyrKa2ES8Ln/jamytV3m/ZNVAIGS5MLr9mTGFS/OQyE9PlbedWoV
CUenmICuGt/A2hCxtKuqpoB7+gJ4eA9gk0vXxlhJm2d5l+Ff/g8S8zEE/na5
rTO8YRR8vvryLHKyKVpA1rTfb5nTN1dmmNYRo9YCQghOhoSatqcp3DFMtfIN
BMcFDWn5HQXPx7tcC4uIMRX5UtyGNM49+zIh6NRYJaVzdxD57pviVSqHLRl6
0LsQYK+L/m7T2fXUnjaATWYqmwn9MX4XaPMZX4c+NKEEdIaCQygX5C9gbBo+
UYsBok2F2+pqRPQX9giUVTl2cmQBB7pUXa+wPaocXHzcVgQ8rhtXRUEyDr+5
z6eGgSu6Z84vO1GPaqa2mDC3zpzv26RIQFZwVLgjTo6qCNjuKJNdFuQ4UR0B
Lye1kD4OaBQJsNI+KzMHEIXcHP9zxZ8HHuJO/kS1of0p345WoYGQnki70l0S
CevO1kj5h4T+a4MYmIP5gmDstKHQhrqV8e/IIZ7zkn8nn+e1F8wL8zbo7fTj
l8zWMOddpxtR2+afmw3IH5n1/EAhr1W/uvgidatA7zTvGSRtb74xJ4iXppzi
FPUPov4jJ1FsNzRcTRSVu+4S+ndEb9nhpRjDW1YPg62hy2yauw0+OjQx9AqY
9XXFrFWRrWx80TrhW0eLfM8MXJhDfxz/QtJurFPVUlpJ6WHtlUni60s6hBHn
PRmfOa34OsThk4H1hMRJL2tsiAVTXluV1IwZJj6G0rkGEA23I//NTJ07CoHH
Xvmhh9bUWju+q09HK1S/aQejKJBaRmLJrchuwvrpqMXDuuDhKXuHSjU32r+/
Qu2yEwsOljcNbsvf81iy4an0HynM+wOCBZJpRRlhv0v+4a+EaglMCza7EopQ
qIibcErTYCktp+0vOGR5VXFzZrTN11f9W8shi4JrHDh8voHlQt1aD4/yNPpS
e7VEHSFK5EPifydj+LuzCk9CJlGDR1d+K99zWpNoXoKcDIVFnFGdrv09Mv+S
ov+Oc39ViCCjEDB/FBbZD8ztMJuI0lUHUHJklzlg2sOlKKp0mpWAR2CGmRI1
pAjxNRZVTPOWsGVZTCw6AxC8fBcWcgKzeSYTi8uD4EnPU3VWcrnDD06ASFcu
B8p/oLoZqFIH5G0C9ZfwMOPtVrQur+Cr76JeVcASERQ8zZajQWjC/k+zFfyp
PrE21Q6rNTZ0tCAjZwyMvRSqFrAwDzWsLH8MfI4Hz1I4B4yQZwttYfHpS9JV
WyWp7863kqOINCe++G3H2BURpCjpIeM3e6eebpxM6iDV7NHUO1Pc6aCuFzW/
ia8q8MHK/LfuYIFS2bF3/s7owWgYr2ivKeTMFwRhkYbN9pMIuN3Z29cExdYB
qS/EGO2dMj0HNedLet/nurnHAkBkGHqnSeQ4hGlexV6O3bc41Bxpx2Fl9ftQ
kWMquSk/YDL+6Jy246Ymu9qXqNtDjXzWwla/qEUmyPdtBBYfwCvqiWbUNw5B
4Zlu3pRk9uGHmV7yy5CWj/WkVbNdV032BNy1Zq3sNKUBc3B9/7gRwYA0IDKl
acwJ+yh+ykwXu1wvOO/mgs7dWsuFnaJax2vCEqDZt5RAqMKCW224sZFPO1+n
afl1HA0jrImC149NctWXD2bo9wwAvVGkG2Y1JR8olOTCr5baXwaeBZmOtAqG
HlK888V2y45ZC9yAhAFmwVBhrXBsfLCwx2g7RMq0EX3+RfAF4hmh5mW/P0EI
JQiIbcZRkYl5kbgZ+Q5I+Ai1rYDsSJw5gWe1HZteQDWXBbhNnjo43a73X0JV
ktj1B7075dnJwaho5eJnBE921Tzifuml2ptDOjL0ooZMQU++kJWhJAQw75WN
/3OiSe+DA1mFmSUGcv86Rp9nhbw+U0FTFtif/UcHs0LHHSCuohviH02PehqI
VJSlHIbcNJIcKNjgGEXvXPUCr1sGfsJB1NYXRP5Ms0N6tAOcudziax395bvI
paODiIFI9qbYXFMm6osYhU7EFfizp1yvhz3wjVjg+9oVdDT7t+L5tJeTbILc
3RcwtE5FdmmjtaFiuer/N77o3hLBR3+MIj1rIuDRF4F2TdzZnAAVOEtb6jqI
0YC0C99JWYa3lRwkIAyhkPQlTSRdkWtqVS/RMX+daVRNCh7FsrEwNnT7StPr
NgB9dN5T8XiXbzeLSLN5+1PlXV7sqQKv59SmtFqS3oHISKZX2kgMWmiymy70
tqmCFrjQq65NiQkiw/lYM1etg9wyirwJGmXDgkZF7NK/gs1UPFYH8KmE9anP
KubGmxsW/Sosn8eyt24JAi1cS3mYvfb378xZCUXuTfODzO/6sdo/lM5qNGiT
5veRoLMWt3ISm7JJBqqpD66Gqz1QB2uu+KW7abgkwEd5bebNzkbJ4Z8c6EIf
VnHm3i10be4BUPSgMnKspoEu8a58qF1+0E7mxmDXAf7ZRX7CMS7VbHTJ/k6q
5hDlDYsnWhiSGWI19eeR7LW1LGIxGNxlkteqJCad89QpxzSF9caRmaPwCSWR
uxmddDxvRNkDt4UiHsqZ4V/TtjhYMTlrbs9D8Xnyd0x8PKjpV5FahFSQQJ3f
PAuG7K7tdlKLU3ACGXp4ERvlgD8ijnsY8AEcg8cVd1u4fXz3o8UpQ+7kotJc
D023/jg/sdiuw81nAZRqd6ScC13Sy1u7f5ul29z/YvE5CvU80L6MGL6JuF3M
R1G6D+BKSCWh+a6vKbGCtzu5yz+FziEk+q070iWCq9kOtRVeHADFrGIq5B6r
ozBDeqHQ7inz4SDNVsnpv6YynJ4Cn5Cbb3FTcvThj3beSjX0M21a2Ner7jLa
8Mt41fPhjAFXqm+3DwAy8CDMjWFhi8Pq3UIOrUoCfYyKuzH9vS6kWDKaJJrW
tFMFwG/sNnJh3GPI7mjwI3Dyw8r4s6fBCDzjW6fuKNT4VVgFXuUC0376Icxi
nNY3FI+0Nb6k5CZ0AMtmk6BjY/vbwprTYtWqaN/7FJ4m7Ch8yf3hVJE2XCY/
/DF8Wbv+850S9Fmn+WIns4qEEla+JBK0YVY2dZPs6HDhHWx9U2zN+CmFy1nj
Tn2z9ZlWOnA20GHiI+QvGbTk2EWqYObV1X+EqyVdi8oknHjTYeyCU5sgnXy4
0fbmm7kx2PQU7pAE9IlTFy0LiQIrIlMnBgHSaQts7HWyxCaaUmJO3rYZr8Ji
QZywODkxHOAwxWqUQz04AU47Dz8zf27O0gcGnfs7FAQWJ/XffHAPwC1dRw/n
ejxAnP/vihqFBLkoegU89vsottdozxJVjezizJUMGnOCQg8iiSTSbBHa9dYY
J2i2cuGqh//egk/bSAPt/HAWwr4W8X4IWg5jUr5FaHP/B93sqpR4WXxfPivX
IfE3Y0lAr1oT5K47rxJhcL3G+G8q2xSxdJkLajVmwtn5BF1snYTpPwnOExg/
9V3uskB0zb1clRwgglLx/bCVcuwpVjZv8XZRS/sKRM0S/Q6CumE4J4SgDLUs
7SPcQhD0xBjY8HcevQC76kmcI4rZaQX85w3T0qBmro4C9mxu4EYAKPaPxscm
kVP7fj9oHlUtfmoefgYW+NmZLL59iSziyV7QA0CeOg+yh6TH+eAr2QARygrM
YVOmBmnh3cp/wSTaGdXN6OFy9P8jSI85xYQ+gIp1aT75bmIAe5iRZIQMKpdO
XF0M9sgTrp5GStvTqInL4dmsFSIEdU/6ZTocK8Q40Kkwld7qPaIn3NA2kiP1
D4QNvKq5sOxAVKwQLXwfUBZDDDwe8X6kWzWbeBPGei04bSsXZrqza0jMuGFy
4Gy0pD1HaCKi1j58RbMzJF0c9hJIpoGTj0+hVSWb5NZHyWHdNve6b13fVbh4
thFPjRDDcsEbEA7/S058rhftRLmqo6zNqOPKFHih63+BPwMYM/uwQgYYa57x
RFqv9kkoH8QYK9n8JIUv5xaeGEcpvG5n20EYz2CS/Q7o4nOBTR7yw9o0bYTU
HXzO3TEpozhI+kNCCBVfE9PgdZSNSOR3GWd4AffiNe8229tDJc/jSULs0x/o
wD4KAB6MyNMwB9Gr+GuELbi4HgAAylrzpWtx9RadPo+Do4C8WT9CeYYxPR5l
huFwSKF+E20lx8KUUEDHvqTw2H66MTBW8+tCx32XAOAWzRNHf+FTBMI8BQ6Y
rNfKcvfe9StE2m4WN0tS32BGqaF/ujdTTMtWUN1ljpeAeLZyJsLcQuTsFhPy
aZzcBIMExv4XHyUrDq12zH8HLtccRzpt5CLfrAcUPnpscLr/TCmj1G+YjxeV
wv9oR58omCv0rlV9vtdC6vOrBXUtnc9YXkjjqRFN+t2OGAV+OdIxl3A058a9
jJpGsg7o8ZVoSAcDVXn/OByPBlZq0O1xeyXIFeeeng+FCG3aTBk07TwGLpzh
RHdZ9ptd415y1MSbTVpKSSxMRFDZIAdddRjSVI5QawGmO6Y6oKDGgSPy9iIE
kprD3MFmBClPsyYWfv4/asnJUab5axFsLtixQH8wRS/HfI1SqkvdG+CHZJ82
AtLFbN3J16KMnDQK1mh84L316eAsOsSMOPOoFr+yz/0+37HoW38w7COSxT4W
cgkwpvc98lNn/83NqUFau+o5oWzAnwsat4/01TUoEAlUdWWqI5DViLL5jpL6
u+o0wSQ1OBiepX2TW9i4Xie+dI86Y/nQhuo5dk63v/4ukfJAn7/BOuY7pT/t
vpJuBZ7aVZRDfgFpp4aTsWXz9I1aUqcBRa7edkq+p33eUnk+Y3ZiB0WA8ksG
YIVx2p+g/0ZADKr7sy3nh9EDnO4MhV7ljUDy4VAErd3kCNyE8y5+6yehtziw
V+2PxYfFQAwy0A17beS4CH9G02ReL1DWmIk0DlNo5DbjrNrbVbMtB49oMl7O
ymhsGGqGcr9oZz40i4DTDIvWOr8zTnuVZ0+9COCDZJdeocW7QsdXVLjZ/ng2
SJl+1NsOL8OPxgt7aBWU+u95wTdmG/KkLqf9/JInRxcunviVXDi1NZJ9by9q
OJ4R86CKomoNhMqEQt/BRYm5krvvYXbY5dPVcLhFoRCVBSFverjXWXbWkrmx
kOqM9Ed1Qj5uRU7QhISRt3RCeNZAQKntMfh64xcoEUDSotc9PVS1qOSN4+Y6
Yeq7cJhradkR65HU3/dTNYYixTHC57nFh3hxcI2sy91JA4I8e1kYNfVMdQTA
fTRqootE3zbHAt/sQTplTARmm7/CXMDjuC5hh5d1kj/22/Mw+lDcISyqSg44
eX3I8MexwpZjp9sWLU3kWBNe5G10Pm6x1Q1ABcTVJ7t+Esci5HZ54gyjDea5
ehKwAlfNbRyQxXcdrLDg9oq9qAGSKkPxkGR1yQWvCVI9bZQQLTJFfpNAQwI0
h4G8DXnNVEK9HcAWMhxloCD9GnajfEOZz/betwfUJ3zVyTOpFPcMALOBs6bE
f0150lqskyE3IrZ8ZXYubP5aisEEmQQ2dvttk8Uv2bq+4AgJNXINf9QF1R/X
gj8fyOgttZ3ceJlDsghMvM4qyetxW8imwV1DBjfYWTnO6vajYhepJuHkG+Gf
9WQe/+/5G7AeG21U2XCiLtil5sH5WT+xqPvb0oSqFCVQxTk0Su8kyBzld4ot
WVdQQ+o8arluynNmG8nDJzoM8nwn+9/xl5lNXBRAFU1aOyuLqStqNW74QaAS
hLepBhFv7p/+nR25hYYDTYfSCRuLYOdke8n6ZNUmDYftytRRR1EnG6qLEiLA
+9AqHstNZbzSbcFfbaPYe6fKXLDpiXjDeRV2nNnbsRuhm0LEtEGGRdMqe9Kq
83o8mlPslGaZIkbsxWkRSjJdTZQU/7/gCp0591inHZDi57Dv799R4Uu/dXZh
6oDPePvapJHFC0U8g+Q5SvqDATLtOvkU/YQI0wjEUsNJAwKV3NAc4T8Hcb8Y
NDVBhDAY5rbpeng1OCvUGanB6UMwoeLskM2DT7OJ2BXuBTD0+1dL0gzoqD3Q
qUMZej4EdADnfT2fWHPj40WxUkg+y9v1lfanMXEy5FdURv8wA6cRfywZSeNz
IkokldFzAuH4CssDzlWLZ5RCwQsFC8PR3zqJ+i4+Cx7shpECaaSUUygmjsqB
mJOQ1FpBNqkxYr5CJDH81CCqhNOWCdi1eHvxYDTmpszib+Ph5qVpkCYtkOA5
Y+Hw6SvRgNr7teUH9ObIatpUeRt6FqUAvcvL+6HE9No5B6emHsjLG8oPDOV4
R74t7VfRrftBlThO5IV41vefgJuklH4OlWvw5JNwuX24dbRXVMznOaOCq7GO
AiSRwMlQhJc4A1+EGGunEKqQNe2aWdi5C94CgK0Xb2raKSAIJZoT1CqUnIZu
e+WqOZqUxlAMx6lKmiq/PbHNKJHzR8lInuP2iaNYtR1/hE8wS/oJPKIoipZg
ZVEQQ3mI7UdvmwVjt8KSZp+e8zOmCz0gE5O1QANdzz0aVqAIbA6N6H9RsXgR
y4vyiSqHVnJymSTX6UG1x3XgCkoH4soFIrJxFYnWUkb8M00Xc3rtswnQrUN9
T5ykUS8stsYAhm46J6dIUpKs9bpUX144CvuEaV2OqU08ZEDmzhD1vtnXdeqT
aeJfQxumuAWbIq95kTqWV9cQcbP+4NOm4YJgNFNocsRY4RnZYgYCEIevIfwE
+W/7tIfdwnJLl0wCiXUepzx20ZoWUB+RNKPNRzT6DwefKNvpCjqKodWCzr1N
Yo3nb6/NkgB4srWevJRMXlMYcfGe+HvjPIp/aKnopBboUyL70OUGV6Glw34z
LPkMN9S+YiyXHM863Gd7/lKgqMw8uyoagoypvZnkeff+Uoid34oe/VB+tbch
t9WntolOedaUt72Hpzaoq/ZtvIJCpzcsCjRhaV/R9gVDj492tkYk7ofUEAY0
wmp0yVYCylyurwtO8tb66ruzfMPQ2I5IdzCO/4ed9JsDXsrUPK+bMVHFLrhQ
pWVJrsFQWSbbsDywT1gK0Yo6pAZRtheI6e8mN+ESEeLznZGRs/R0XBsgRc7w
/115njHZvlCEcBUTx8aRW12Enz1uj6a+EkvGtRXZwbNV493H0R1JiOuajpYj
pW0qKCG2NLItLT+1tyGfXRaGs5S897GBiZesKooNmFot3fh4Lq745ctmlVgy
bZMjza7ReBX5q27qgfEhzcmdPFaCfUK5moXaBmjumP3q3OaFIM7IWQwfndmr
kaclOgA2Y/8a3SAo+j1zKV0tW4tRBRnZixakBGyr3zxdiB1X5YZdLVSKo3A+
Zy6MJjgOwu8F+nZqB/v0AEJKqa+txEMptvxbLqID35weEDY5We5XLR/OpuNb
GixhEtH6mnZADSjHZPSCdCQ46Y7M/TXS8EsExEQ4H3QcYEXsVcoZ4Ajj7fh4
g/xrs5QQhcUJN6viGgX0c7Lr9uQQIuFiL4rPW/hXPhC8NFHDJ+nUA7imuxw+
tAyPWfwpNDXFxDbs2pqkqCJtsyiSzCU2jFCEBteuJGrmDF+4nczm5J2DJoXt
hABKaBtgWXHlW9bfOpieAJX3EUbJJfkjnCZmXmyrNyfTMCwp5F3W6WJK+ugI
J651wYcI/JdmJa0CITl7mMQZiiT/W0N2gOX2YCgq9TuK+8SwxAHnvtRcAzAF
usKYN2Fq5As3PU0zeJQPLCallvSVXvAub8jCNpCvk2Vz7WaYLIbaS6V6GM3O
Bim0wWV+azdNCKlFpNqv4K/Ga4Xf0HAItocwGJ3FO93SGC+//ykw29pcPYzw
FolaRtS2SN1nZgUdy9YTVaso2eoh2GoiQFQRgipSrTobzGa6OMEulRKEn06+
jaUNd6GEHQe+fwaw6a5OxFMBpcwQx8kGhp0lhi4hQilGIBP7/62YpiYKVUdk
iJzzhS5t2LX5UbchVTgxPflIYpCbztW4HOS+RcOfM9w1d8FnaRpHY/Gda6gq
p0ZzMKM6fu2t/qLNXe/7j5N8H6OSxdjfWhwFFC+ZOje7s7GaKESmHQ4O+Cd7
hLoaZ78GXb0JfY8ofTgArVxay3S8Wn+dBEWNCAYHfeCulC3vAxIEXk9a8AhX
kIVF6ELHnMwM9YVh+RNmQvqYSC8qhkPxrvAXV0kX6Tl1hHziz26j7uxI5cpq
cbLuQxKBhOsz/YKEYdQt4drh9LtFsii0nJgWETH7dMEJ6Hmwn1amQT3g7cXb
a6HOu57bZYl9aYYVSRHMNLJCd42zcfHk3YtpssU0TtUwIMFDTVKRUjqrVheE
4Itrd/UDr+rTB7KFNu2+D81/Ejd0cFVriGnmdUAJcNAPed0sj6XXQJ0dcOLy
lSyEHUgvmJzCvnXrEjuPP+EltqUjvb7F0mobEtgTGkt6PmWyanUrngkRSFSk
1PPrTJ43wOgpekd6yCL1S8ZbjqELQ5w46AbPbRycP1d+VI2knN7xL2ltMCuk
wTSB5fGngWNQbN4QN1Bf+l6lBNOoe/t7GuL/c/JsUe8HtKoJvWZ+I3X5+NZL
MjARXLfVXFho1BEqyQbiUOlGIxd1dASVgFN4KBPT/HpEBhHu7ILaMROA1OU+
K2j+rHj0I9YXZ/hfplUip0Nc2aJnMcZ5JTd4iZ3B/Zz+w9I/Aj7BPv6gNUfu
QihwL48Q/4XlIGuT7Pt73Mn5PPH6ZSx0lEgzRPMzPCtgxPD8cgslcMdM8scJ
D7oiS4VRYw3nc11Kuy1BM/4ROoofItWLGNbsVqNoyfpHpKQSQ2FvMuy4nsCJ
krc5kJLXJvJIu93rlTA2zcFZecxk/CA1+B6xz+t7o0LcIxnUUeOmYwkVAwzR
4DncSMglDZkUJa/zFPS6cJ5gMquzZ4Pt4cQ8RZRETuGKGR1/Sxg27YRapjn8
0odGRwPz+9myvpWASdf7E51kDU2+7zAxJ7+saIJfGceLETUcMbeQJZnwjz0Q
iGJ1LrY52poCVnzSELFxiqWq14pvQIOYP5jjVAjPubIn2WgVRiHeuSMBLWLM
3gIUH4QHbde8w8MF+Ruc2VE07vhxkKW1o+FQugBRCZfcNKfiQyJDE2NVZtGK
j7rIBdmeh/T2t7/aMqVCzgeyNuGeuh7CWLB+Kp3t18fMuFdJUyZ2f1E1xfMJ
oRJqjT7461LvAKiPrU8Dm9jDgBg4JomaBeqMaatkIabn6Y61R7BCbuLXC1x1
XGwYRV2pRaBHlA1CIHJoYwx/C6n5ZEjPBOjyOowMtxRU+1nzDtNPk7DOSvAY
fGKZMcPHsLoAyvBgkrrvu9+2ck9bMNICz6N75191K0OcKqMejnwBZh0A0LbC
WhfXaf4IqOhQSXTwIQhAQnvZjw4swQVbOxb3X1FerzDanTHMgdrBeX9855Lk
D3FzlTWiwMbixx1WpytPVsrWH9iMmvaURR5zLlrEse6+7ufpixa71kIAh1lC
UH1j9PEeupDu0gTqrIiWE8SzBJQ7NqntqzunDTbrjSbR0V2sEMqmjU2FmThO
+F65VmrQVHlf0LJHI5j0IhOuJ5a6MHtg8OwZ9fH9udRxNfwPUOUCVpEI7put
2EKGdgUXTOd+OP1JprpEVzQhiv0ie93o7TMSFwhnZjn6XFRtBUaDuW/RMABh
y9AmzWjA/ZILAqjeG80RCCkGWguTFPXrSiER35fevckTqcR49B3BLsvXStiq
zMTZFVKglKmvM0xiLb4vD8QLCn5EUcBA8B3NX3r8XGAKgzOpnHGHh0nuKbDe
44pYySTUUEMDlhWVq0EY2HpSWiEfBJtS+J8bmRExC67wioZThQ7pd4I1Tk91
x9XjTV2lWERFzoi/8UhX2MKz/R/VuqjWTGU8nYrsfVEVFwpZxflRMQDF8/2e
aBAWQH75tgqkmHW9dehzmHXhzAvv2lBSHeVkhES8AKzI0rdaIJGG0qGt85Ph
88zewAAPgNeCUsMzMsUZV4s6UV2XEARfAuc73Jt2GOknVjwC5QRn7UHh6AlV
MiKZtaFg9B/LdXekz7B0kDp5v6KnV8l8FQEYiHU3Wx6UIl9TYiC5NU/4gd6y
uacdgdJxps84WBrrcS/M25/lpTulOssCYwrynpaNW0mSekGyMVA4Ydi5UJdg
hU+9F1+gVNjHIAAURtNDfbXD2L5LGmKo+X9pe2BqeQj6ivavxF4PaMPagKi2
y6bDQPuEWdlbm8s745jL9BZJNssEXerbKcWDkDKMaj6njKvb68pWRA8yDN70
7o/k04aA0D0IhoJEER92NJ5Zkqi/+DihcLd/tOZRhQ2HZRYEbHyMXlrdzYKO
40iNRttXNPbsabPQIpLvkbgBg+yZMjbegOL72KH6f8GWFLK4Id4TZj21+LU4
BPM5Cw7expA2KTkzGLoqkD8je3uKQVU06YsrU4HLYEu6g77J7+xxXXdSLr5e
VVAfsImSEFj8pmDoSf8mjqKVfSKA9qxAsqs//bLagfjOof32KT+8xa9/7VL1
MmCr2RImVsH06hSiRAB2zGyR3OWNNs69aOueB2V/pipOWp8I8BqQR0liECXp
5A1mG2sCwvC0m49L4GAHRT8oYT/8inUKF6vd39TTR0g/idJ3j5oRcld9S741
9CQSX0S+czMihPsHZfHqJol+NS94knQtlOKNlWgdkq+lHDpvtCCvvp0oLv3r
vSvnHgyjsmq0vgu/q6xJbLydS0Zil0VpXUxr1tfTe+TaH8pcVYOYJ7acRsXF
Mn3Ej7sxwc1QtaexmU6MOh68LkKbOEN+ePQp3/NPfrx0ab2yOAhQSPxdhqCn
eNqWOpXUmQZFeoCZ3W1pNOQv7GzQwkftls3Ykh9QdlIPW0G0+lM3fywebriU
RaWNhtjiJzefP7f+wjyyuHy1EBF4sWu+0VQGeD0QXx/7vC1/ouiYWGBfia5A
eDNn2fjp2dKMbxOt5v8UXIYFtMCPumnfIxxvuYzIvc3k1daauealp3ppQzlO
mvss2gBZr0nYkNCgagWgKUs5KZuAsk8WpdQf7WRAtouAgzrqWdN3ba2nOo5c
3Gi+T0uvy2mDoe6FVbf9s9NZlQdZguzmlX6QRHpLFoLDkcNPWKOD6HZr7Sxq
wjnCU3boNrfnrwhVDVHcysWh49oEwmrgWrktM/D5fm5dGl345XjD9JuzLpiE
wU/EiPYSbNsGzRhu0CeeW1y6RsmEd4XpQ7m2q/h8u60XJJLmA5CCJuYUguM0
7TXwYXmL7UkySMBbv2AQGJCk4JoEBLa0UcxjVY+frkRyVrCCxYIvjZxPbV+/
1KxOp0Ny0YN/nmPDv6ccI0Mkr+BMo/5pUMIIw97eJ9dpwQHRVFvCdPb+zsUB
1R2WVFsf8GSI7GS3vVcbhE4uzXI8h01yiixbQ6lqAz9qDKuFBuuTSXjtBrT5
i+VUBX0m5syAxZLez3fdsJcGBGW1nDltBC5EWMrBOS8kPVS5E2pq3sf/mUmU
ogeB14siP6E2xbSofavplNHRCZhtoL7tqDquKkLc6Dyvfki80CKZGfQJOgWh
adVyIJLxvGpkwNyAdK9x4GGWqTfZj6FL1BqRkkoz9osdz6bgozr6wMjZVEWo
2CKdH+iARjTh420lYXH1puCbbYr7SgJhUnahJT4FMnNrrhz45aya2EZ45hEl
iAM+aiQL9v5bmPzNudh1qMAWAz0ldxgjlEEctYQCPxd6tayELG8KStPamm/b
TuZ3xJPJl0Asf4VE6csNvRPezfm3OWX5l9QI0zOzLotxuZ4/g4LBPU6kJTYa
ElNKCTKL0Au9mZWHpXplH/MDFW9BmkxMXAVVebOM2wy0evvWPwzmmDBb3ANd
OWKQxk5W6nbAhAYdjYnsU2TSs/9ejY0+oGvEjtvPZ9tRk17SO2XupIg5gztd
VbGbFsNHf1otqIV9rxd8/MfalNdNvBHirIv7HrABvGwlxYKcb81RDXvb4HZ8
jwzteFqgr7ZiBPz6ZC4UzdlPSoS7HinIo40g70Es9BEmBzaCCUgrbyVU83Yb
Dy3qrn2QV9fDyN/rwUdZ2DYWApVVaBfAYSGijtauCml7Aw9rKEmXRnu5E96Q
4b9tSbnDHqcS6U8JtaTe6Wd/+istuSjkEdq9lv3eWxgyZuPVWyd1oAwAnn5n
sWEaWWvq3G20vmPfvSQpdvMZeeEyNJMmFQgwoV8Q0SW/dcoy6IJCGre6xIra
v0ExBhF+M6nbwHlTdb8O0iV5gXgw6EtNYbZVGE0j8+0TjGOGTaMu0moSPhXm
KKooJdG5J6xq5dzlydFb3lag+KsIe3WgYl3hLayWt04PR9X0nd5suNmHfBKU
RuyLoPbVUih6E8I4bEhi37uEuTTiy+Uvchj1OhPicsrS4UGKMv4MSq6k1C83
89tVyggxrr5AvCRpQRA/2LsVv1CYt1zm0NVNfodCQu+XVQ8wv9Rd5KJFjMbH
gTF7zXwb3ZL+F+V9AEDvoxkDEUA1Kii0xqp1j/7+dQ819k/nDOWAj2mjg20o
PgY6lZV89gxCBxpWXtgpqgDIFVlyIFTkAuBuvWio6f8dr46arKV1MUJmh3Ns
0r6PF25TYzdtvEQt2K+RzT6kRXpUNZ8J6GMNAF0CPRwyp0nms/hGzMKs3goc
DdbUeX4PyquvY+6MYCmopHqp7ay7WjHMzjXbvaL4KJvvMSaHZ+uwF3X+oYz0
mASJFStJ0ON8YEvfm+1SD+0ehxEll1HFHyjAfltskJxDuba47G9+O4jceoEM
LQc+6AN/00i5KSX3SaYXWIyHxJSc6oErQ7G9hQlzlzFPRsLjB99a1UXG1Psf
UawoWszyceqMDFq3FteFrpEA5KQqhJ3s7dmcIobeGlP/L4y6GZdS/rdx2rFe
Fl84RgXmC8XFJIt53+amyvF0KoX0IMxp7JXsfuPUqJk7yFfLZizMR4BXQzo2
UEsR6V5yVOLOZCj8vXGrMTvnVBKmbP+wFM1FgAmqefsF7aDenb7OlV3uwewZ
Jhmwf+t7PEpxp/cYKDK2Ly3rU6Dhf3QHlT0OO4/XTzO7xbXc+V6SGZddnigI
CBr+JDlVi9OQAzYW5yPzw2VjkdTw3vrSQN2Crsa1FTlc6oAwQ0rdhtEopsW4
7qqaVym+qy3Fd6QMN2FaOErmQqeZlRvvrrp2KT4OrjPlXRq8sTc5vmYJVh2R
h3dnA0zEL/anbZaqCR9+Owh8wmykQFeSiP5JMAV9hpZdqT21buQDvyFZG1Lh
ZC7prLWqLvN2RKzXRwjzTdvzgcdWMLf8LkRhc5pAYMOb2dhH214JfM9wYrA4
2YdUj5ICO+UkV9+W0AEN4C5g79LRRfzUvDm9Z3kjiks6AL8FTcjVCwClJlbM
JPieyaFeVRJBxDT9MEE3wj/oHP04JY3qKuLy+jEC8DuE37vaqyTqJBMHk4Gt
DT8bYn0ubOT6hZCFqS4ntspz2GUbvxhwWsxrsiH/r7QN/MNebH2Kj/sD2pgn
C1rRyXnmXDU2NJD2kiJrKS4YvtwO4kfWEn9Wdad0RL1VX74jYc7owMI692ZZ
x40FVB/Ps5cHvxNeQy12Gjj2/pd5QEcZCB8w/MNhhA2/fh1/kwoAl+uXLmkt
sJyUK+sVpcfpb/Ry2aL1Mu7D2JnG9zciQDg9R/xyoah1A9jo7lFYLL+gXbzE
bewyEs3YsDNTscC89JO8P6/ycPn+FqhcztE/I1cvyjRc6RZKXM38z/wH7abT
eriuHI5fwBtFdi9xvl64NgUzXVRtPuBZq8igsjQW6UduLA0XdfwWg6zs+3vS
3LiHH8IU9ISRMKDB+VOzGz/ZbKFt6Jr7zIJeFGTtyW9p42DD+ceQ6DYHHq+B
YreEtMkkLjsFr1eMvxKn9w8+/AC9TvZHjVbsZopoVmk1I/fNEssuYKYcyHvm
Y+dltJOqRuvAmbpbLJ+bb0qJ263V4hko++ij03yqBU4aocBrrfnrwtwdK3fR
M33o52hHNSqxNig8N0/Brly5vTsLawx25Z1FngEgEOBop9EliB8wTZUQYS2a
ZWhFM68HiB98szY51EIffnxYOEtD9/jtPOe+VoXrSd/CjPi74w8pF9Wb8kcJ
Jc+t+kWPoV7DUDePpcZ/RfLTaJ94yWAyNdVxGbNuUnv1r97o7loLkMZ7WoN4
Q+TlHfhBNzPOuiuCnNOUwlB3YzofQn/KVZsU2Xgm5aKmmj/6JS8bs7mMrfUd
ZHxNC20nraifgYPo/r0FzhPwPgqTMAffCHzltdPTrPfmgIG1dvNGaGH/hZ2i
SKFAp+4xodO5BDgRF0U1S4AnBaiUTu+UU04lHVYxQjkwad0vDvbw6w6kV4RP
XrwAkDZhDOqF/u/NUZhUQiU8RdiGM21acGmq/xjOSJXOew1BWitKlsvCyanE
b8JRaPLa5ehh+osx/peXDHkqIJDjih4hMSkMgc1mMQe0FWaNGnaDRu52m4RR
YH/Cs0/7VHdBj5I4JRTFkzr8ZNiiGHcDs03l0YBMXyB1++NDiPWnODqymqQn
gjLOFU1ozqztEoFK3liDFnzUgwxhCk34SQqcFbSNE3gDicuBFb8S3SsCoD1G
PmOTjC5Zlkj70ayCTLBF+d3B3UfF3IvBouE1tz0crVDM2ZU+ngcFZUcifJjO
vfVmkCHZi9lOUgO7H9L7gasvaoFe72EVYJ5j+9zK5bk1W0BZu7e26pVEhVSE
jpnB8PXIHIrOIW3sNAx46D+DFdKQpxeGEu3a0P6LhWBsyeQNr75V7kAhVl8P
Os0Yd/HHMbmR5YbQ8Uw4ypb9Xs7VLf9eOjHS8qp7nrOn7aM9wkTPkJi2ikTw
sTaWRhGFWxfeJ7NGqNrqQVn8zoss+hY1cw8CiyRLn/qvJoQePNGg75tqEnZM
kQCbT0jPKMD+Ih6cyEmEqle1tsX3fUjNXIeOxS9E0+yG47Rvg0IWIYiarMlm
2TcrFfjW19Ty40Zw1ro8ou81E98bAxVpFZtsHjLwSZ6fysz+e73Wa3bfvZWe
E1QoYzs6qnv4zsT8d1YtSlO//bBWG0U/zdJc5PR7YU/1zodwjDQ1RelS0Cpn
3HahmIANzj5flW9z3Uer2gPKIupv76JqZrWzZC6/efFMHDLoF4mg6PKW7iCB
Qtg9cxGemfIRHjbZLzAe34oY6UFVVkb9vEzamM2bwMtmtpKQbK+6BX+UV74h
X9naQdMDDscPJZy53ave9RpMsFurwlJIed0kITmH9TE35zGu4fjft9vibi2y
PepXrHYD+gR+VKNVgMyWelz2cRWBod4K17OXv5pix9lsFV68/2CGE30KPZG4
u4RpbRPgPFOHWTmuooABnDbOhv9By+vWoGBlHKncuwV5/IWnzc4F9Ab7U+1/
v8d8/tyTU8b2EOoO1A0xiLByvRhiKf98KmPGgrIt2UpC3cJOXUtu9KpeD+Cs
Pg0GSgd3bHijOc9y+fd8EGRyhUXEzCuvWpf9hFF2aK3w5mRMWf6OYN90ysiK
iu9P+g88CyUXjG1Rfm7aNBwJ20bbxW4yTCd2auhGk0QvJSbNCz4eIsXhCXBw
gJfg2neqJfhZ7ax6Zn2cXuatxEf3+CF8sgPMZbryfXiv7bB7Fy2A+GKPRBiM
1Usx4+BBYHRz7d0xgsP3ultwJ4BE+DFVELZpXqwpuTIqL4vJEXTOANuNjipK
XEfJ3dmEc2TEh13MsD+8W17uAnbY8qOzkpbHgTCWTZ0PBP12T3S1dnqCfrjK
0CGLx0mjLcXjfCdbSOYXc5aDBX1LuKFOZzvbCb7D1TptycwVVfFMTspNKgn3
4k+oL3rGyz3vxJOPYSy5lTloh2dr9QoCaK6Mpczidb+RUEbtBsN+queRyCof
QPdG5efNWplLKd4ftEh4Q9eTN95k8ohi9gAdcn22ox8KK7MzlDTUUslq9T/P
aqbdzXSLGOGBbgF5gBJ1cjp4O2eSuIu5UsrWUQ7FL4JxbmNF5E/LTGIg+wLT
wGCahJ+3TS0qc/Dj7SsHJCk/+6T0mp9WM3H+6rfYTYdaMfQZi493YzNlPaEa
LFBXND2XkhOJD775AjxjOObspJSpeotA7JFiNgSl7nKV5kqZVT63tnCb0NQk
vwbqjCsQ5iqHDUkbHRb6Y5imDkvo7HNidkgTofTI2dxsYWibdZ4IdEA/Xq0W
P/6im/TWbwi3il0K9iZChY45EophKQXa1EdMfDBoQZrOL4bDv4k4DSloT5Dx
XKfhBILd5thI0nUkAcU110BIc2E7XeWn87dVhADqSjvRWwpUbzfZpG67oary
8ZkYf2+7fi8xbRbs9ZucA8NYJf1gM4UzQ6dvwQClG+NTDoYvLOu8ILiHJbMN
XzvterZu0ZO8dKEhOVXGPTHDjwgKXl5fws3nLm1oiymSLZVLYDdgW3uBwVzW
v8TZMdu3VI/f++EYp5Gnk/dQ3SWjD43IVY55SZpOVA6ic89zwNqFh75LbOOz
lvHh0z40ij/MqoXkdFJqcssbYzfr/kqKi6fAnSOnva+zoxmvsb+LrDVpHuMQ
H+CVIaMjHDMM4BZvwBa1Q5+zgCtrz0ozQCa9EuOCzVkEGRS1cQtuU5gP++Lo
9niCdonoUwDIFyH8eEgZGTHKLDT2ZmKICVPcAwy7hwpD+klqMcCLtZPwlbG2
AHyfzwXk04N2lOMVQTtr/jjdUAvCUb3YcSVPbsfsyBNTpKaD+Mdr+ehS8RWW
YSfNPfC4IHyRHBmIAi1QzAYarMClvt0J+xj8qqFWYb+d+2UHKp/siF9uRiyv
RW3Z3Qhh0ETyfu8l4VKExPPI2Z9P0PMBCKtgRKQ+HoenqJ4K/HgzQpmzI84p
B8vDlqG/qUxSmzITSNR4ocb2K63cWaATQ1eplz0G75u8Ti6j3PnoRiqq6V4v
nv8hzipyR+8a0NCqiCkuV20AIIb/7ClHnw4Ani5FAzx/5cQJ0XLBXiw3lCbD
ylTdnmEe0KaUTp8HQRlmafbYhdpkefylP6oydeSt+aNeWLrQmVWui3dJ62eG
kY7i25uuUCUBsFugfbLHnPhYPSXiCBb1VU262D3cak0c3S3trpg7W+a/p70g
qsXLUH/lP/Sn2EgRaOyVDfso8d8cyYefW9HsMPJd/SWWBICkJmj9hjYgxyWF
e19P7U70lrYy7Y3KvFNn/rZlD6c3pq5fafrN83L0/otRXf3UuAfN6JM7PdwR
bSZMqCPC3w7k7JwpfUU3DrAJwActclTcsNKjxsFbgx06ZyIMdVDYWtWpoxQu
3EqnZF1MGTvR7lY8m06NBWJBRHPl+8nEKQt9Vgbens3OvUyY25/7mBswBc+d
PXomSoOpb2oFQMUqNIvwoLWd2OSVN+1zcNncOBs/lNMi/3k+Jf3X1CqvI4ym
xlFRZ/eVILZeReKECLgKxgvd+4gwh4KM8LkaW+uSu2F93hafNpSzMeZANb4C
B1Nt46IeyTl3akwHuQE4EQlLwkv2Nh/NQvFO5IAITmlJu/wYftf9a/8RS/SO
os+dEIX7cgRW/tvjMzjrZO7hoqXMtDUkx46ZwggEoo/W/hTYj6shFTnLLzGw
INW9/PE7ZSEFwmZmZodStuZgk27uk2oKxMBHluWz4We1fPJ+uY7CcAcNPur+
78thVjH8KK5TykTRNhkYrvoZptgKChOBFhXXmKKkPOQU0eXum9zUsLAoDO5k
s0XG/HyKPfKvL/Pb/0ac9EtsGHNKTLev089MjxgIbW3uI7C8s0jraVe3ALrZ
llKlrWqOk4E//U/PnwMLGHDkxBChDAiIK4VfdagvUzqXpw/3nAiLJP7Vdkrt
ipItTsv8IkZzNwO4zxjfBt2t183sizabSnH0zJfO0DQv8tefiCR7GrwC1zrd
0bFucPgF7PCxLGfjhckz4FHeIidcoRWXBt7hlbva92sDVCbLlHAe22xaeVtf
RKNJ728MEV4jNTlv3RMBJ4oun7N1Xi1mQlmM1vHkB3W0n1JaprDt0intd2Ct
MNXh4U6bOBnIbtlSktNQAMrL3l0EttaralSR/SAC9mAoGRXLI9td6VvmsvZA
YBCZXJwCsu6BCyRw0/oQuulPndbcbUGQskPkcCEMd+ywoD29RDNG2wvI5INH
Qh521iubolrrE2aBfekK3oMi2BNk8sROgkjNp7ifdPVGtUwFCgygdSznbw6z
ai32K0pTboxax6RRyUx+uRahcHUwuo/KKfe5RMh8UYWt8ifjBbp5aDRjnqiQ
GN7hCQ92jm/diWXDaMKl08F1tnU++DcNV8ZP63cde9QAHKqx/ShPUNs7g7t5
blDU1yh1rGx2e3Aw20NSFNOqF6tzBp8YtQQNVjSYW5qMbCs6Xt++BD0MhPpQ
FfJfHS3vmmE01Uz3zIDVNQXcjhsOR/OPKctncX9cX1jV1Keab9HX0db4wLQ0
QHgRIE9000uVariaBAYDCFv2sjWSd+pxhu05QBoF0SrfbDMcjH5wIaac9J1g
81sXGREd0Rjz4n+KqAZb+tI+bEq/cIElhqUIK0ijTyreYQxBf+clZoOrEK1C
O8qDHPzmlje3S2IyyOtQXu6IWOLmBrG7YdzTILCqod82i5K30xhrI0sr4ktU
neB9SFR+Wq33TmSNpbfQ/ZxMvM146ziDvhR83NdyXFNu2YoEqHGbEoFDAfSl
ipaDZb+hycMx5LvAx5FD5X4syihIEtuFq2ikevZBdNeKyGjAEyassESt/OCL
RdEbmU7jqQGJp2YxaHQ+6Oc3Tli+kNgPd7nNZUL8ADkdRjikktNPZkSjOlLU
dddfixdhFiyrsSHDl+cs3kHOmM6crDdOKlO6m06Y8XbhLTDq1izbsCvAQBTG
IR74/93G/4bBs5eIu8G6d488uqL92Qo/5Ln20k6As5dbkp+inocq3FzalHlE
RLNk7tVxKQMYcQmVkZx6udh0i2OnsAZn7ck2oADPsKNSUeizGCvRrx8Je9QF
eeu7ayCVUidLfK5ZsVoSq15vdrV58Q+8hLBy2yvZIZavIbuWALjDmNKrTqKn
o3OQeyoOA4FBAG5CQ87DCiiNJSFOdEXmyPetRmAOYwdRts6HiPff+3+D7IU5
5/ad19ylC9tKysZWhlgOvVBdRGAx7Z81hMArm647Fe5pQetJ2XOFLjzZ6Ysk
L3rMcF8dbhwCr4njfKflhZcmzzo8LCkSdwO3IGwlp7tL4nuKUAfpEyeU/QW9
WSAaXuVr4yRQzMwndGwrSPik0okIHzbFH6PfbozsbhmKyEmBO2b320/bVidD
pUmrqFWF5ASleZmrTDhi/Zl4SaZSIES37j7lrg3BkmAWg0mACzI86P4pdgqI
bJzLJRxPHURv4lBv9koue7lggcfwwoHMiBThqJ79RuqENVOw3pkPnCq8857C
TRbqz5diU+nPrrf7YMguRmnII+5nLAyGDktZfFhR+dDbFyiF7kdlqLsPcETY
r9kN9HtdihD8sjZmy0BDArIkIjzQCpr4+AXeTUl8ND5XiuNp4l+jIdJ9Khx2
plxg4ckNDcP4DnIPYOwgwLUidvth9IQt5hIIfumER46lUn0Pn53A31hj6knF
tRkgvCpMS4atU9oEd/i+NpVOtXNTQVivjQQRoYxU5vhgbsWq2blCL7xd4LFt
XPYAgkMu018EAer99q3onyP7EajEztLHGa6FBPqYDF3eM29Nenz5b7FDoe2q
JK361vXkEWl33GkhiwBdMz+A8Udkal5MipxvlRfKRWdQKsbGCjJng5HQdw44
aOggz/sDNzQBzcZfM1ClVaW0uI3beDJZ9bA5pv5WB0Vs8fJq4FxIbj/UDIvG
LRJhmMd7ywATAkTtxBbKL5sjhcbDauDly6P3PKN+oMWGEgzp8Sojwi3AXn2V
2OxCJXJVqo/wngN+zRrdSKCr8u7F5qaMP0CyM1qBVKdo5kXZpqzDQ9fvzEIU
rfagJwMyoqnOuBvJbu4omKIINOnlT78LFvqHCiirKTIEA4iAjXUUn33M1qtw
8z1T6HKFgVulBw7lkQAF0NvxgQdPQ9Vfw3UgDZw8f1rjdkli8DExtD/YMdcI
mNW16qXkC7RW3uT0gP5oXtMe0F5HZPUNc7TwdNG6xJXiP07LEVwMTFxhaFjP
9OMHXVSKbrS1Bh24PiJCmvQuNhvMZc9Udrmok8yO7MkOmVLr+A+jwFQyC2Z7
OnW/LCmjd+v7BLCAfsydxncGDh7vYOEspeUoOmC/pt0KEGhj23RI5cfKsc5Q
/LmJeX3WEy1NNiiAexiw7M2TY7YwO1Kkf+D1kydy1NtfkyMWOVkIj5YrOmeI
OgXPyauyPD647mPYh3+o7T580Vpa6MIez90D0DNhWXjlaKeGBjAu33at6Pmh
oj80qH0C344dvkWa699K5ddpt4yOCodTjj2Izgl7mfjR6OaBniDAAttXC+ZA
0mXjH9LzRDuC1EaWocrCR+xtMFZ5QGjsaParR+/DPgTj3xVugeZf+gKWoyqy
fITN1W1DjbSjZI9sgUSVw8pxX/KHKQmcfKSDZDsGfDXl68VUKm9Q2kt8WDfD
TWbnMNH+yT/6Jw1a7I9YISYmbMywYJeUn+kxbYWVDru24+V4j5n9UZBmdgyd
K+ULDXAPsIRREVEKYUAXSqLKZZXbHYs+cG2goCL3VPmyKFRzJyRzgMSFxUAi
efHSY9aA9xi+ou36YP06/3IM6LOvV4RYehUOKuAYpItIrJu+KjzN+IsYYsKJ
G9Txa7PWMZOZ+0lEwJTMKfm34jQM9SHNQje18g5HRyXMQ33hfvkFzCQw2xC7
50WhcgOAlnlGh6LKRVEAgTVCMaUcLW56lOuY4ZqUmZ4pE1rKYrBF6WGxlNp4
3M63DSXV/tBBOG1DFsnca1yeARA3WIRZYLbWMYFBKvo1+T8jc7tKO8OHsusf
ymW8oTPRQP9kmB8yDExBrkicbqi4dUkf6lG/Bd+iIhx+Ahz/7x1BB0o7Wc0m
eAoaSk+qamVKIqfsUu3DpHKYtAKtfiy1QHLtSwP+CNXHKujxR7BwCuqkDvrw
/mkkSNX8nqVhRgX78nIu93DLIRjKifVPNjFKKR2eQd71mBD8D89+8owqWO2a
dfPqyvKul6iHqUTblRwuSgozJR3MyFJUEqFcuDllAJSoIdWdTl0w3WJ9hCgR
MCnR3hORhNlnfZgQR1ttQVA9BSpiZA4ENnHQ0nJvN3qAVF2TIz7DYKupnoNn
aYNy+6oMZJFkUmFP6jGUOsTb6ug59P1u7oqlso20DUGZpslgKGe5Ts+v8GPB
9wp7b12AQhZkB93DU0TTCNgK2t7NJshRYUlcKE/5ffO9ks9lddkV5viNlPZ/
aBJHmTL4MQDcLnA16psyOWPLXIuDcf//Jfrel+z2AK1XBuJ6jZbwqrsSkK25
Ev1+9wKJfgn/0jB3xT9DbTJ5jcFpbqyFvNgTVghHHvSGEbenCZfh6hoN7aAz
sg8zYJGKF4Y+A8/0okb++heXQi+W3mh4SojzDLicLCsYKRW7JKKGW95F5tKR
3mt6o5Crr4QL89QAy6AYG1xMgyDxD+xDbowCt7AbaZD3g6CD2Px5SYREZdzc
9kkN4nOdm2GyEWuoPvrPQufmyNiSVXKE/jOVhNHfz0XpQfvYHb5l8UXJpPK6
KxvBKDOHlM+EWeyLDkKDklp5TaOt62ycRuOa5g7E5MvTwQEg7dNvZ+T664pb
k2KyGMmCaNifEN1yRMIvEsSYZq6MUYotELR3++wAK8KhxNKQNjofB7EYCprm
QV6j5nDz811isHKDrhh7h+si3TIfe7vfjnulkKXkReL3IBCYKYvWVOqCl59O
TZ3wIhMV7K/zCagTZZBY5Jzk2IGW3xptpJZTtPaB58PVL/TFZSgtsN9sgM1E
VAJ49oqJxdJtLbIv8dOhpvwU8QYoTAXq3M6UC8EvSfJxq8Kp0IkN5dnYjo1A
4U5yGlfygeEhCFMHM0bn887ju8SW0V0bWTvdbI3RxEMlQtJOFP/Gg1TFzhgo
/FZQGAYNiKJQ7inJ5rpxoO7LVN4Sw24OvJMKfDhYqtsD+NgifZ3W9xcTk4bi
YmqaBOpcg0JMceHklW55pjdJUMWigsHnFGue6wuqx+oDPTG17ANbuj2gNZot
53COvR+rfOXuNfkIb64gqDq7Fxn9yEAC7rC7Mf03AYA5kw0rOEuSDqGuK40j
EugvpmYi5rUl/Y1Fm25kxlyN2drvEJcV0qbV0moCrVQnNzwLs+Q7QsXWP6+j
8/lJhSnLbNG9y9yDJZcMDdSHNA4CvXDQ1uNBEwym2/o9yKSwi/4tBNJKW3HX
q2hqk0MCqFkczXkH7RM3QdTLRMXjiyoDD3nyqLgXRLR5eqFa/gHOE/XLD2w/
0tu5yXZ+0y/oKSCkuaCbgSN0Vulj/pyMCVqHWAI/LC5KzAzNBv5NnMbbG62d
grwAmUF4SJSWhHUc7ZGrSjDuqQkxNs2r20G/qPsZdVw8Kg2GV1tMGm/Rc8ww
Ufj0Hcm8kyq9gHS9rxhulUPWIoqAaHMwwhJtU2CH3tOMmHleYwSfiPVBZ06n
fTRX1DSKnu1sMqZgqteYBJ9Bkjxtq00JxAHMYWtzehqnghunwYnFPgF4YHcq
7rQRpwbiO+R1HL9z6+ugCprroq+lrqGqij+KwSCb1BqenU0OB57erkjhAAuj
SFC8L28a5shTdk+wA+cPgIriEg97ipK51RHp2V7ni3gSINMkYg2H0IxhugA6
B8xBRIsVdpksQgdNr8hZZl86rrvhDK6At7f4UAyuUR60wOhZ6DGSTI1+oeEf
D9rc+2AdBn910H41Hu4moPN0JE4GiYfSg8t9UDUYGkDnK3DeEkUFYHkYnTcx
23zjA7q3RwIbvIDUSJcT/wHTHjKRULC+XX8ignLpIrvnzyH9g764BrseEfZR
ZRD0qxBeWURnKuLLXTCWoUCTQApBHZfn5V4ovvRx2o2Je3sU9Q4WkRzCern6
Jo9nB5qBPWVkVvXA+v40pOEpzEMmt4fzeWim4FGDuW4XRYCXdcif2ayO+c8V
C5HPFfwDsVYHdhurTM+2NMyK5LGZwZ/Fc7v+ZnYwxY0blQ36quzmKnaA+RuD
2n97vLGd+W+wKZ+Ylx0zExw5oTZJxD/gSVGtQoTAZNg3nTmoJptZEu6Pxr8l
AH+H2rWR6GsTlopc2WR/jpGuyiESsyGdZyxCl2dDwMbdoafxWqdRy5fLgGFj
MmLWh19Mkf7REB5Md5ZPAtjYXskeFZM8gYZWrSjyFjPyoVSk9zy13jyVroLu
FuogROOR34ojR42q/e6IhVO3BDgHnQt9kEaycBqONVkzaFbfMAhkiJk0ybYu
Q+dGcrLafwMk0YMdg82Keu+/25nrMEhLHZzkUfdikdDRluURAwl9jTob971m
uYZ7gYQzwlKr7OT3r2lfMruu7BLwYCtMemkTL5pqON7Zq+B09G0XIv0/9nak
zZSa+Rxy/pP+OpPizIYXBzNxlgIMTj9YcbioQtJni5urbfJLmXhM0XOIUp0v
sgz/bUUnE642h+DTIJiB0kldjrmopIAu/Bto9gDMQnoSi9dMztajLSLfnrEd
EQz9/H87T/XO04+OGtdv+CLOMyyxfvAHuuh24RDQNaiRqcO1hihvbgPg5Jpi
hOz4faXq37MR+1vMJwiLHbB+aknTFXfZv8xx7z5+aI0RTGGr1Ngjk+mJ2pK9
tg8vuSIzRCaBH6OTSlxFxHo1y+fp9N5uuL7sWdBMfFBN0KdCJAJqqFNXfAZa
FeJv0JionaFgN33q+VztmowdzeNJabWLhuBWvwFzFHrMFhLFWIZnZEAOAptM
cIfa4gKEQx38+KI7G9XiOd8Ed7IStuRgld1TDLXA3NxfQGrOwkHJqz5rxZ98
uEECw1S2mbBIoGiQK5ScMttQY/pP0Qm916v5vVkP2DAxeHRUv6Oe2/uSLEF6
EBAcmlEkNwUeDdAuUjVP5MQK6pfxDO4e4/nYqBzrrnrEOWV+MnCxKk5lNVCD
aKd7tXwMmh+tOj05Ya4I/s++mnxx5lXdb5+CGiJ/lfNFuswqNG84QZyEQiAt
mmcBzkyPOhQuimRAV524DZWFzhJvAvy+WjlMfjeGReN+895hrcFQKEjmayl7
ibvdCmB+mSPRKIllGfOc4YWeDyUcTuY6DEliFoJhpH6RuHWpe2MLDhwbuW9Z
rrZGQ6wBbqiIZByqrIQh5UwcmkcPDmfZ9p5MCWVMFmWvWNJOwpMDgqJ0LynP
jhd4oVX0NB0GCpy5I7yUkmdmLXJCDjcQyMiqg2auONoKxU7RGvGvYIzWlCkL
pCwlVL9Zc5VZK8w2P4+jq5bOVdqv1sLJVUnNi4l5maN9w1XVSRzBwn2he2xo
3ffJQETK+YKxMakmqM/Y3oy2KWJg4sLFmJPExzDYfXSzwqq9qvuprZwLDX2F
gzzZZoDVr0XuqccQmNl8vLS53rxQbQMuZ5jU0tObp33sA8ujT1EZ97xhGLSl
VNes5p/LnptbUKRBaTKJB19WWS8TH/cD/ZdiJY4usOYngtPuPBiT4gwN9gpt
EiTPW2w2Xn6U6RDOXzYNxV7Y27KBap95aDF+6fqYwTbzKyOKmMUFBYYSdJOK
7BQ3n6Nq0ToDM/UTBmwamT61KYRWp2ZWXvuZE9OTnhOO34k9XXScoxMfT8o6
DONqDdllxIaRREiZWNjDMUoedMC0rIprPwdlZAsb9tK0zLPF2slkcQ465vQe
Emx0WWv2dF4xn4+PRp/O0tMyLP84QkVCJqrgiCiv/haZ/5FGZP5l2fPfA9Cu
8dEBepU21h5dqRbO7tpYfxSv69AjoazQ8VflvGo4wNgMZNQjzel8y0Bsk8xo
iRRYe44rl5Ag0nAuuBCE327Rpd+U084UBFH1/3HxO7NlcxK2rPl1aTNg5zFK
glFs38RX8zMVVffiH2BMKyB+X539JDMcFvx8BGScBt2Lyq+azqwdbqtA3k4c
kQx6wfJn6QBHtkwZCu06mZQb5SbfQfzGTnLKXPGLGT4WBk0jfWf0geDdn2cG
jrPxVZomwc8zVq9j+bDSPrKYyM91TuIoigocBhuIdVwApadoPyR8JjEGQ6Z3
64LbwZMb3OvfDmVY57HS4j6cjbtCHt9OPGPpSVGaFAE1WHB5W+F6So6n56Bd
QizOrVWd/dhqE0jBHRa91R9UgfRgRLMMtK9702VPH9zZ6CfRBv4FPhoSdhsi
p+ZaJDvmxfg3vM6lD2HVC7FLqZO9Xfk9oaSTFqJqDgBAOdAdr8sRzFVjLAdF
bgidLPkWUfOcgrlFGCXEL4JVsnZ/hWIpCN+z1+4Qbnoy6gFfflEun41HgtKG
1XlL53obKGTZXlv5cuzNGMfYO1PvO9xj6ey/LF/p6xkorbuU37Us55okZMUI
meS/JFxTmE6gV96ZEaFBCIgSuVxNmAxlXLEtDXH1Jfsu606vKKWXJCnN2NQh
bQWKa9L9+22uX12H7iYckiCi/pXwmZtVrisd2WTWofqpLNc0wiIOE1ZKkzB+
KPQUfpfg+jOC2gBuZF6sTuSGQzDa44LnVHZmnzOqGRfFp9Vt+7TblpJV9/ms
aVKKRZHrmwTg7w5OZ52uFTF4UqGcYPcazpcDL76fF1VnSRCrTIKivNTUbcWc
A5Uwx6PNxhmWbPkhKt90Cd9fIFomXZcPNr/QGJMxzBLrE2kVczob+RQaMa+L
MFWy5ue/5VppnSxgKaNsZ804vIQ2Rt1yBnh1pDzNJMLLF9uyU1N6TRQi9xQ8
skN9H7D+ns5W13JVLPmBHcmK2hi/gQahztfdYgNlrr9Q6OUDkbkSkGQXU+Ar
M3bm2OmzH5ZFK+78TU6BYr6dV/Ef2cNMSthDMM6ynHANlyE5V9BUbgi2lwFI
GneH9K6A4qtKcpLYAw0LfZOK9qV//iZ7e9rAxTvOg5xngvtW2vDK6cPItzgV
yO8NR2SpfOHUQAWT76HYaGFy/zrwUsxbgbNWL0t1hxqx82KNoXEwQQa5KYSD
VJIf7Hbrzuz1fjD796XbaYNKFAq9CO/Ub25CWdY0CcChSO1NCJRMwxC+mkVy
uvK/BtUZTRu3a26VssuJxumJFRHMI9NRjEKVHR2NzwD3O4lMPcIztJi6ut66
9awNM56SMFrSbMHHD3QUXC8YDlb4u87bv/c05JH4lpCOcV+IWbHs1UW0O3fr
bR8XbvOAUXLKblpY/8ONwOne+8FElC1M/OYoJlIBh1JWvu41jfDSJCE6Olnj
rKd6tZ1ZujYiRX23E2FdfpxxsnG1wAC7L6gY7tfCksQJKw8LNBniwdqzJXN3
vBa4N4Dpn6MFNA04ZIW+rDEF5FSofO7eGnQtcHnB9QgYXKQseUrZ0CIrxsqL
emN5LwOBoI6vzMPWHsjVO4Mp1wVl4BpCvNTnO/pct0/NBMzoG4A4rIq9H8PQ
+A9CgYlqFhpayvtKh5eHffDg8+yf8uQDcIAh+ytXuR9LbkA4Gng6QxDdlsKI
6eCyjSLb3gOgkgCJUJSxkqm1ybL3KOxqAUu/237F0j2VGc94TXjML98/MZhz
nTG/hiftNiOv8n50IF3F8wKIBriQW6kDXk70H2WpjtGCENpDbR3CjgvDx+KV
TrBE5Ecub1XQjnR+yYnLFAyigem7n0hz3KyspWAmWJQmchOT00OXI4UAwrOC
owSGcKL/tlRsTEKbWzUjFeYC+GriLnJ96sYw1ltDvRQeJhgROCFIK/NZ4qLr
zp6GOGWWxlOFdhY82ArF3cd1bbIeL6Ccafl4XfLJttrcjuoLKcuh1UfRtiwa
4wQNWFTH5lmMFquTrfwEau2vL/sMqXsUJZBaZuU9V3/6UezRdPsB53Z5/YNA
lIj9eZrDYXVpVAscZhe0qCeJn+mFKWB/kmCUHt0mmhJbDHHNgYdhdvtfxfJx
kj6eZGOeafb/NfDFqscDQnKip7pBis76LbonKnjwH9SDgrO0kwmKOqQgds8m
MsdXguKgrdtIvHz04EU6yn/p0urOmnREHcQS0/GX59hqBtqLG/fsJblXvsEh
Rwz44uOA6aQFkTmCVfHLdBHZi2mKRKKaxv0HwMzjJkBb0XE8lxIovv0vgjHO
0TaRYgpovOFso1TrV0H672bjfBmyZShG+MUgocE1sZAurSB+NI+FsE8Md4r0
z9GZ2kFF+PEMiC7banlwvAi6Y5LPjWysIDzKxqb8V2ysbuqCm7LYYp820Hir
NU270cu945iiVgx66tyOb3Spmw3uGhqV9KF/3LMg9N821OCKO9ZPu1C36/oE
g6MOsYvjtP5+uGs8rZp3fL4rHP5DKjhjBjcsrlgoLWnT5MemDtGvSHxReLTQ
fY2NKDlavfcvkmtk6eCNCYA3bMQFAU9Vw3t4qSu+/GulYjGDzTdAZChwm2nT
F1p4VV2r6VPzXYOpJ39lhAe/PtJGgteM/MXWiZUV0BN49wmbhwvTbLfqV6Cc
/FiruoIU181SJ7ygBitPBayKB4x26lDI5kni+IIh/+5wNxzx76Kgj9vjj/6Y
lCcFHOjUCAyt3IIWkvMM3IYMP6JyXyVsOij+4Vky1YdtjTJlbc6GPYLw7z2t
8H7zdk/W7dRLDSbmBVFXlgCEjDrCksJ/H9OgWq3KWBUKrN1+2mz19clkhuWo
vFGJP8hPCDBS32XHBXKNYe0qTFFmBaBkt8Opf/IRuh/mP6gv5Fda/kCcjPfy
gwRwvsA5zFu9rhlRHXpkXjG3znTIw1kC6RmyGJ3sBdljGFHl2Dy7WFepuziE
SjMESmYc12BI/3COm5OthFMiIk/OCh5Qi0rUWV9b9kiq5Ed0xLM7AbwQOft5
RhU/jZ0imA4a5yyNkwGVJOJsnmA3e8cnrrs5rQEid4LJSIbvghMJLSGXTRR3
spIwdqI5Tt1KhSAKa6aRRDtbEBfTaQztjxglX0vjil6ApL5B6d4cY1g/T5HA
/krbhzmkbvjAt6WTZHcC2IW9+ZB17W/d9q59T0ImaGSXzEdT4wb0HKL4ihan
3AJbwxVlinUJ5RL0O4KantJoYanvbXpZnEkAGNRW2kG3pZ1PydLIe8ZY/zhC
MAjKzTlExROuNs8DiD9iBUN+zlTHySR91zegEgdmNBNrLLjfz5lhJZp53HtD
UfiD1qa8+oxR4Ro+10UrcAGL4X1zIRsGNbiRzDRhnCi36xnBFoHm9WHSDw9Z
eh/txclavEzqd5ShDqOdTiPZrOyZfaFn/0txmOgzgiT01+jC/dZJj4nMXhso
vHxmA7jet4b+UEhiia4yNnOniheoHsEL4J6cxSSF5dfo19ckrExqWnwjSxR1
VOjvbFf2izsMIQmtpdYJnAIxJ2X6bSbqTKzQLv+dTmF+GFVSoebhmXXEKzBs
9elqnwQaywLWabopQ0M0VcawWxAhUQfnqMubvzj+thDemMxZHTfGR+qyFpgB
xI3v1WnJqHkkOHXZ8ho/uKIrZOdvLXDReDSDqTjP5D2hFlO1ywQExVgXKgtj
YjkiVDZ8ySLXOi5S28AbNdjSHgzgyf5WaDUK/0UmUQF/xfJwVanufoou23sz
e2Bp8XrTIOJPF98Id79rLLTUnftwtF4REP6iNl6RgurjCRMkYho1l1rAMZz7
UtlUA1F1+6MiXhofR4T7/HDNUfO6Ay0LamXMT24PP+qYudm8RRIz5cRoUkLa
3BM5I4F90kjnOa5jJ08KT8L787gK5KuijoeAEJh9dowq0jYCFd/UOwjW8MYw
6gBPasLz7OAarGXGkkfao/k0dek3GXR0nfHQRVmVBOl0raP9wIqm2V1pWZP2
jCikkWj+1PARkVFF5bbdVA9qxgnh8gZ0g8zL9H5rn0AXMOk/TQSlp77oRzRu
56oCKEP0b5oVTbwa12dnHhsY9SltkWkwdZjAE/Pyx3c1cIAS8lGe7S6koyeS
TWZV7BmHeoBw7Md0vu2fm6zBlt5kBgINq+CuMFf2HflLc2dKlrzC4Z5NEmVV
T9R5t1HU9RfWHZyZLTFF3MOdLwSx3LcW+OElI+NmuAjvEUqM9WInz4h4PZ7H
8LG8CL5OkcgJak+mjlSD3VudV0Y3QIuj/V1ysy9Nd8kinE42EUjYA0uMxh9F
hZQOe1D7zw4cdY4Z0VWkV3BAavbvg70RelSTtuoJG1qeAl4ITJgZvbhbVwFa
QZOS17XDVKysyM2f8lNYneNrymvE4Ys8awuVPzgLggdZy9SFJNN3OqPdYa9X
pLccJNu2pgcHWE9qLpvl0SQkBgk0KHlBhr37MJZ7+qgZFDZnaXlkaA6q9nOE
fk5hXcihhiBfIcMm2vsjsDlqylFN5Nu8TF1bH2YWBXNkyyE0rTd1s4RWgAd9
pCiyB/yUK1ecOG2j2za8FCEmKkoPIqYpqwPwSkZVMZOXP17WS1Ljha7xWqFF
GDbS4soz0IKKTkwJk+zcCmd1pmjnFBX2Hqvv2a5rMtbbf9ksT/88jWiU0pV0
tlBoQfWfNe/bWkmlZQPfv2o1sgVb1iQR+hldNd40MJxFj2HVjmXpMgkPruU7
TnKhPftvuNPyqD82XxPDkASOa1Emp8Sd7Zsy8xdDUCss0jL8BJFppnfRDXJZ
hFiQWW3NPu2XfEvC9ZKzya7XdRrKqc5zBB5QJousf2sks2MLhHvqxLDTyBxc
Ky9DPvvhmm2yT2l1EsdO7OQEa8YLaWHmiKjwjQWG7zVxRgREb15r0w/4EOP+
j2Niva+jpBGLZJSekwMFS1AuTRVgSHgOtkO2cXYhhGbYSw2UC8Uol1jNnmCd
ets5xG92vzXBMLUMlRBx/6vG/0mcm8bIC54IYSTmjTfQf1wraYsQ8i1B46lI
dOVyJlJTRybOQ7VP5FE4aHzA87EKd4xVwPlQECWBb+KqGee8TWOppe+9Y1AG
XPDY29HE+9Pae5D05XIo1tZYvE9tneQJgAHh0oSNhEUACFPqujATtIe3a2Sr
AIFqqL5L3WpNHB0BtPukvDZMToEGcpHCRrIdqIXKz6WxKLw4XwIWNaSScyV2
2RGlCCnOs2kZMFV2Djt3J6+4R+HAyM9BSEzERHmpfboW+JR+IgUwdOA4Fb8i
mAegfhVspSmCNTEjcMBbDqHj4hOGE6rVmMqAIzIVP5QLRD6zRibvE9SCfUwa
7AwHs+91k8397lCU6K/hPXLHlbLM0++LRRMT8+agt9fTrXx//wExQZ88bGWa
+AflYk1+oFGCG9q26QbPHUpPZv4Bb2V6fizMMkx0z63rY84toI30ThWSU7WV
2m9d3/toP/bXKDLgI321/p6W6BR1I3Tk+/wCDBIn0icjLM2edLla8cnH5GpZ
KhVt/ikNV5psymDSdSGWDQ/mPpEEN1hQP3tNoweHKpkWgNicbq6DSL/+MCIB
kzFgxuIpCTQtYhz/me3C2FB9ctDMxQb5c7vg5bJKwqrCge64xDaE8mBVfha/
+Uex8abAXO0m7qJuZx9nIWlBlhCOHIT54QVvcDYOW21TiIRSv+Ml+rIu7tDT
0hkAua2RFlmi4xq8YSDrr3dQcoju4LcE3WD/e9d1E+QZZ/W6LgGTeYWztLCd
Oso/qndsJnuHiK7BYV8ZLnGeADbgJjw+1HyL9bjLKxN7n25atDgXcxSg7ixp
zrlORzjSYBx92Q63wmzUAsrjqZrwTdoh19s7EtVi5nQ3e0INdS3lJPcn/B+c
jbwlLf0PadPCLFwjj+awNemY4C7dfwdzLjXvDCrihDQmtjoz7zaA51DIhi+l
91OGtwG8qs86VmPtFKHEd1Z45v+z8M7hLA7LmQIb9tQD10uBo7nNr4vPO6BQ
dMAkAIN3QbunBCCouXAhAoudf0xoB+dAx5NAcQZ7bIjsI6JKizQ3aQimyKqY
pNV8fpidoC/RuUUX9s278ECVcct55KdFke4owH69ZNHACRs9wDilAHSv6g0R
7g3B64OaIdR672PCxRmphKdj39q7OkCN13DXtcxuMcfu/oqVpHImBNhB7I2h
PxScbACG92upevgR24mniFf7AWGbJ40PQtD6R+k6Mz6uxN0spHRZzZ/5vcXh
6xTJ6yLftol4mIyMtPGZkEU2bDahJzAxbfBrtXssXnIW4X8QdTSse3c/nrxt
Jve2gcuMKLd+JL3pkxMCYkW4Vf4++FF2zyi3FYA+Wf77wYalEBO5GctMx9HR
Gc9+pFKkLvolbl3XsETRz8/5sI2pfZx1SIYTO1CT1hDLKLkURiop3irOlqCd
STAtUYUzKzKlq12qjKo9GynnwzyR+bgozw3QpmHk/w7+VIg6gThjKJSGW9OA
UGk9191NWtwJSu/qocJBekkmm+iZ9ZxErQaCAB3hC5N25RhpKb896yEdvRtq
rHfIrJ4SpoxwKzyGrikqP4fS6li+rmomFSCdqVWeHiHyR98F9ehlBEqRHcmN
bOY1zrfYn9jH0dF9nvA9Ev5653ZDz/oHBa+mYumoMK2MAlwE88OeGfLNCDGk
IoEz01ePbiAzzLqnJ/Bngb5re2KINH8MJkPFM8KnG2T7HmjqelhK60vb73wz
4u+mGQVue1HIg83Z46B5ziypXl503xGxrtUUQIZxtqOvVaM7tjWTFjv1XKsW
tG0EpKhO04J8KcX8KXfpZUE4eAKilMfdDMua88Cd0diSXw88B8Q6pR0hGWeP
gi9N6UAZmCcgOMr8s7WXO86zwXRRRsfncAuhBe6BpkX9B45UIQczce9urHJD
093YjBdPbo9udeIDC6QSbJeuMz7tQ5oNn/VJ2UH1adkesce+i37+0QWTKG40
PgffpdDmL0QpcAdTB4KtY0gOi5S7KW3fEUNJuZYPLNICKQTm0e2h9TDbMxMV
dKSsSKTY2XYMYNCZyxkUAhDx9oQItCxxcxAB7dvrhM3lGRJIPTYHT+IAC+0a
WRLV+HxCYiJvA4rKOptwhVtfEi9PzoKDwfk30ROLe2YRsAYSvCnlRv8yxjVT
f0+gzPyAi8T6WWejEQa9SD322Kp0o280d/QcxJ2DVZw1ZyJ7ucvRUHoM/lGm
fEJohlfV+GpuCTDsGjLx0iSBCQfWM9OG1vgFUY46OYtFxSKAWenrT25z+/3j
2x6RqLbEjSQ7esHHoaGbQlAbFlLQaiSUmwBU9Mc6UucimNTkFCInEGic0LhB
Ie9oAvagEYau13+kmLsM8Vwxgnkya1vcj2HJPUeC6x+6uRJsZorqNSeQVaT1
RdjrSStRQCr2x77P52rO5b+hF78QXbuww2enAPK3TKghfqUHKW3QcPFhrLb2
PSMASrCChcz74zaHcEZ2zG09mdl+dE9bgF16tD2EpU/B5WWnNnRF2zFAdPmh
AELEd3tfQckRzdHkEQwfymaEYlVystQVVdQzDzNXZqEthxRpScJg5AOIcMut
LSBN1OS1E4OiGNzA6lzw6QKOaiJuH0hwXk6pPR2vcVDufA1xPU6+56vU2vzK
T0LEhVn7isWwGfmS86H/eXcrus4yAmZ+tMCbN5MDCUHsI+ss8EfFfHL+Bf5s
EEWhsFC/rRW0dbOHEf0lLGKGtfdhMDyr/xIsE9p+jifz6r/OnuCqauWZ7fcj
egQ2o3bEo7ur70Xnt3lnz5sErYZvasRxTW1DMOD0z8sSWwbRwtnPJxLTUd6v
juDaQ1yaIdAJOclVzDe+kyh4iK9l4+BoLsuskjJ21yQFDbA4kDre6qi+adi7
//nm8DyQN/Kzmn1QH4eFNOfvMJ754xYdg7wKTbKPrjzEjto/ACDD6tMECxI9
SRDEC8hoi0NjiM55Fywl6vURZ4Rc14/ArTFFiCo7CNOzLgppUHRenBF+ql4d
SEi8Dwe8pZkKDVqy7igrAUa/u7i4C4c9gOMWvLhW6ywMrNMEbr2nl1+eakzK
AmL9hWDL/kBmpiab14wAs+NFfZ1SkbT7L/n8NCK4Olz6ew5VzPzG3axvCOKt
yLSuBbNX6vXBhU6GLNKtkMKsL7GMjwY1SLlDdbo5btyUgV+8PH2fjfJlef4O
q2aYZt2Ja9Vu6Xofoa/0twrE+6Tm3E9VSwlsxu7QjApotlYMsiaUUDB6VjBs
WAbHYMYtLjHTLLiJsbsD9jhbdKmjxhVJxIvloMvSk08epIuj7Jrv/RzJWWD9
oZvzMEKGf8iPtaJisYzsJbzyJZk5HhJGvX3Ib0zZzNWvBELgABCDWCJgTRne
ds0GhQkARdjKZCFa2l2ONrzVx9yrTVrLWeHGOEpXZFnuWZELhL8f4aL6K5Ie
GlE36/k8N8a9llS4oQ6ZVoumXkmjVtnjQXTnLkv0D7szeQpKOUyQJPLAFHLH
CGILV42DBJ8cuv3YZaaTXrTOOHiGmH+Ci1r3bpJhmfEgvinfihHdsOOJs6ST
zHv7PAZrhvpFH9XZKAQHosIamrhFx1M5XwfakgcH7gg5ibLbwR12/reUEMwt
owq/SEHFfmrlInb4rTzgldcnU7FAOcg/ka6kvjNlJXZ9r4tVGUcLlbK3lEAE
73cTJgHeGut85c6MiAKhfvKKC7t3XrlpULD2NB4bkYucxbpnT5i+mxja/NnN
hT7SVWiGjVflhxbozMpCBnLtb+7+73nKduiBO8+UhaRbC+OvJHioz2AJVRGf
0wgv7z4Oci/9Xg5q/g2VaDhaSVfIQjRDpKyRmd4bed5fSDRoS0Z6WKJOefB8
PDiCxtGDyNtj5EFMoOcyVzlcgZjTsMVaDzWfBrSJMB0XDO5OTaZ79JaNwjUv
L+O6CHY7sZ/TvRc8ApK3fSQ1lpbkdO1lGp7d6ejiqYeMrN1h7IiXtX0tocL1
zrsCuu8inUXvM/jRf+Y9PL14mV4vF/s3ToUDn0IEkEuqo2JB66tQAP6r2e6d
2lhSGPAmhbD53Xv5w57AiSBkrrV4mxaSGsP7OjQ86QaKID938f4ZkFYufB+8
OPP9HK/VCU/Xyc99le+hHn7UbJcaxQw5SyExjrO/T4VCMzlKCrIvN3UcTJsu
N3gZlxkcT3MgkaCZo6l5+pKA8EOcuV0h2RzlHnvya6uZ5aYueDo2HAD2seGa
mOgdWpf0Luvf0QuBsCtapYtnvlhu229xgs6Ud5budFK5oJxL0KsKupYgc/7z
PzsRdUuFroO8KtFI6T15qbTe1yN1e1Z6kXZg867GySXDclozij8hQ2sMVt5V
nPXC12MB4NH1/65H4sMXCdqSfnk1YClwL/FfKyaJnSTIg2YLLZVw5LMIGeou
nwiJz9uPvBSXQuft5k1DOBRTQuejP90wqw5d16OxbL3BKWjjJbkVOt5NgGS+
1cR53w+rCPPryMa9gnmOEmAM68Quh6XJjMxprEjyiDvOG8zoRzyTDDFRU2dG
d0YxpnwQ4jE5aROS4ztIjNPyJIx2RdeqJMb63tt11ZwPaMlL0KAmCBvHWpCR
s0mFVz1ozQN0hLS5InMVAFXuaeds1uCkDwGc8yGZ3N2XSe9PVrSRkCQNMuV7
P9/i8X2tleJL01jA7Q2XPTgbRFY1XoTN7ifZKEfiDps+F7WIJHhmpMeqg7Aw
IZPEhA3/guvv9x9V77khZwWpJ2aDBaK3l54oTCPvCOs9dPIYKClqC/4Gy32t
I+eU5XqMiEBGZhYQ7ID1uS3oytcakwBN/fqh6ZRokFjYzMwSD1NPxL4X9Qm8
Ggn0Lv6tqhj1jjyAYvM6/KtPBUdBA87zT3Wvfwu1JmW89OoUSvNuZph2G9Gu
fC0UZAdL5gB+yFtJIGS7lrn0YcKcDhDnG+UjJHG7OdlK9wUPrrzAHgJegQGR
l9frghDedSiv9k66diPFGdRuAaFl28JBZQmskT20lSU71FrR/oBWksbk30LJ
kkpJmeW1X7EYx2w7a2H19WmgGLWQJL/Q/3deqGj3VCOb7KhsH+16kHZCnaXT
7iYl1NOBKghYgjOKGpkIawpHygIyXqH1UpgRdWEESono2E4Je3awTjGyUAym
dYhcOVaCHht9jWGvXuBF2LzYBcjA4o9V9B05bSIGBz5VR8N5kTwPxBLU0Zh1
80GuumT28eM2F4RWJJQXr2D19ozyBUzLFz+SvN6dH3+0BNbPk7/2rzczavHM
7tFAPKUSNWDfLnZAXIrrn8K/eCTV/wh0fgPPbSjr9Jkk0XjUG98iEBDQ3PH4
mQ4fA5kVserWQR5IR+3TtHjg2DzOYhiFnRb2zvG1JWiMV63OJNVCXKkX7UdI
D++Q6M3yXEAO7L75J8IE9RFgoU8L94M6xPP1wWkytGX/J/53xFdbbbd2urZz
C6pJXT9ioyaUzP3A2PiO2eOoX/K8b1QjVmtaxfBBxTAFTxKGoiCfVe0WBzZH
fTRh3qjAj4fclk4wuWAWnRsC60ywtZ/4JDNY3fzDv0vtyhLTXqm7qOLk/Oqy
NRm//IdfVegYvlN6AzmpQ7uQosg/+Nmw6KGyRpMAh+X5t3eEpRamRJ8jee1t
lDYVWTu/uFi0ePPgM7BLghw6qnlDp3PEnOV7SIcyPICZONaVmkHtQ3WkVb4K
0+pBUGBQ2JIMhzfrNhsUTy8CvgF5gp5XWjIUvHTM4uwP9/zcvVp8xrJxoNi5
mrAbkGuPW3bP+x/hqqy5yUJ7CGqDW7PT8CSemjT2YBzaHAUiM5BE6xwjOcyu
iQ9qzIfWB9Rjo0wKpbl4RBd3DD0esmSNcm6AuPejx2o2e0xJKvnbAZ7gDFde
SCbkLVY6f4KVJAgybgpwViTwicfNGSXmvJwE6FO/iQDr0HY3rp6ZsS5TekuZ
WnJGl9y0jfRU/74hPHlNu2lbyXjt5gNE/oP1lKuNOrZKbJv+uK74CYmMHxcA
S1uO1Xy1MoZ3nFpRZnJcNQ8kaXqa2hEjVu5SzlbsjfZwTrvu9ehj3cFci6ku
79Htwh6BVfHZw6JnW5vXg6xPjZMc2cCOp5GxU1Dvax7kbK9eTHSOeyJRY9zC
Pzy0+7eBiLb4IYm1oU46lO2wMNzgRCEBvtk0pa9CdPpRgr5wist25knfTV8D
k3XmD896eIytuIXPdgh3T5wkFH6kf1FV9SDPK7qEqG5+ZF1k1YJTDP6xshz4
teHGb3JNIV/4fdjKRlQHzRBUJjN9lxGNIHYz4SQaRzBWXJX5OJslk/pT3gLv
qHYK3N/B/Zt+CPDslXHRkyX2Ge7tgM9iIAJQ+a8Q2hF1NVidygdFJVZDNXbs
VuGKUgBsR8+//XReyoJLcckIWqe///KndVTEQgNKfZpNxno7xkMxVBNEE/vg
1jZftpjrgPRqxtIWeidzXHSVk0KVqOGHng1ZYQQdlf8lxDwPLVnJbCTOzFHW
dSkrtbipPRmbJhuHGlunACvJ43sVu3cfB1aJZwPcN57fHLzyGk1id3F6kEuO
xq5BRU/K9ABecY2dhZWPA4zp2/S4MNpUlkMJcD7Ola8hhRNi+jV+EiqDC58w
qtBbAPGiDL7v9azV1p5qUEHPt7QIwWwZnsDQKyL7C4p5iqQK4Up3I4lCOAvz
4+10PmBrHPnCK5kviGQc+D0CKrqiC5aBANtQUz6zlD+uhH/8WN24i2S9eCo9
OUvdtaS4QOp6WUhHKF5N5qpKiaE1IxuFUrZ2tekeMGWbaYdUtsLK4ttuVQ3g
uK5vkMaw7SXE1vJUPU6ivg9IjzZZ1JuDOIGKncADW7upObbp0D+kL0CDFAhG
vp7MAVYvtnoBCJEwRFf7sA60e0fBa1Q6Wa4wOACSE8X9qtsGxdS6VCavvb8H
0V9a936RRu7qd7DqABIH4D5XqIkxKU40Pv2wrq2KAmpEEp/STsnJliZLrb5Q
OXPSKJQI2QqCKmaNZnwt702bowcGut5tlx8wMwdnNc6RVL92t3RYosqY4oWc
puQeWsJ4DjLoC7dw3cFGK4b9A8FjDSI7ZM+X4+QEIENKRqm7qgzfyOm56otB
OygfwBRfYPwQlK/pipzBDDRe/BryV3HgJy094UxiwAlfo+1cqCPeWfDKvbNX
cPHDR9YUvkadhf1zNKd2niLEsRCcV3VBlvZ3QkYa2wSPeSJED5u+ygc7whq/
r5o1ytIZzwNP+QwUavbn9qUSNrScnZZ2wS9cS69Ie6scFtMtJoFQLp1xO2S9
Fup40QJH8/fdcuictRfKQ2uVfy2UHTt2ufu+HvkNh5t89KOJyzOGLd40VJfh
1yJgJOqvfwAJv4jN3n2+QvOfwfBkM7Bk097l2TKxgqgaKJcbzP066jBhllm9
NhGnYbiodR9RGUPmnaZXK+Qwc7MNz9gnmaEwmXSmbEZfZoNLlwRzJ5mrAkd8
rOjRczO2mlKCMvz5igdELog8G749FQKJMjQLXG4ARhpiivl0TMui+dO4M7Bj
93grR7WP49lO0xvRQ9e1XQd8wl1y6Q3E2mGjyc5V8aH+NxdA8/txLXqN79Wc
XvSLyoB+dLCwvK0fqEKRCR2ODPbF5PJj6Z4PLX9z2XNrwsADY0Kw/VG39DZQ
RrCtfQ1jw69E5DvKdsDJv3vwa4aslOI8zPzFpNgi9QLsGEwhiW3QWIsyl+gF
h3d6pD0gk9YJIGKOV4YqVfhLHuMBsvzlSMXAPOBUghsvPPZAES93DfUQBVis
iN/FEh4zCu5W7yGNNhVcoNuTREdmtyWnERUcvUbjIPRk+15GZLzJKbxSM2AF
KHXTUc3imPbdXJhgz8JZXgh5OphmkIxsFWs+H6W/+85NkVDA1KEuejgGCzyN
p6uByAyzE6TkDc6YcleHobG3K9edZDMtqyO9XKMFTpcficIY/uzGa7nD4oHh
6YD+JAdq9kc/Ki1ocyZYBv4AKUf+HUWGlBa6vP2He26n59Wdn4wsCS5J0tTk
m28S0+qOJud8IGZ1LzgI+eW2vTW1TCFikOZCS7E/nFDQ7B9qq609WkUdugkd
q5IQfkVJSXCUMwcgm02AXz5TzgCS+1Po7Z9p1vnDqMcBqCkW8oJSsEMsObl6
6DlBNWiSJhTIdVPgzvBT/FsKev/BXPanf3ONZ9PVEe722EBTKAqNWMMbJEDJ
lI65BLhXH3K6Gkl/AqFk7CuM8FPsVkrLWiryWdd0XD2wEE7ILoWV7uy2EDKH
sJwNpUTLi74QvgVn5Nw9vTfa9tMZ8wabqLq4Ip8detHHRHGg31yBUNHXYpaU
VNaSdutGs7iH/x08uJ0sL8odrJOhMjOzPKgUTzvivriJ/Rp7NnPCAXcle75u
YwEM0IEYlKe+O8XmimXWIU/IYE3NOX7u0M5DtNDoXpr+vODGoZB9KlcJ///I
uA/p9YXk1W1gjxoyHcMuHpS1HLOxPksWWkZKM1NzYb0DvcfJenN8lJfQVlaR
fZkIj8twQ+qdd9kwp5tCoz4/SlaX5rtW3EXCcc5SkkzcAwqUwoEOncW4GO20
PlBRnKh60TjxdbBJHCCyiAZoBZ7woeqKi4XlrBR/zn2kAWZ7EI1eaK+/WRrF
K+bb+0eUyyKPDJdvK95uuZY4J6yg5WIJT5KmeR9K9uY9IcghFdUDmaH06P92
qaZzx4gKtH3u6jjpsDU4kqb0wmlRLDPr9C1Kv5D20wvyN8CXSQ2hncahvpBl
AA6Vpsj6YHiYuy3PwG+CceuM1VrR8GGw18y0WhcnGeJRJ4NsubheCHi+0ZdS
hDYD0W8cf2grB5CEhiYlfbl/5ITcAIZ2sZ0/usaD0uBTHCSTn5TXYMkM97T9
9FALIcP6E7icZ6VDHkYru08gozmU3TGzx7k9NhCNGZN8XI0nt0LlUdShRAXC
W43WiNAj6RTFdXpY58nhmOvVvAqEk/NErLVH467VmvHemOO02TsDYNkLsmGy
4JPQ4Z/rbiUQi66MlOlRYUmWNq3oM/mb6DP/qyLzSxRyCS7cQC+/Qps79uNv
E/mBMkqsv0mOVyAQc3UOzqEKAukiL4SRYuRHiKZ6z8I0+kcHS2ILtMdtrEuq
5lsdEZNPZL+JegaO28JXvNHy0szLeCZU/ESJxLwtqHEq9aLNyVlbiFy1g4SU
P1qbg0KhFYUirZpHP/EvQ4+a1fSlBb20auGoCArFwfvv/44eMFdRpPXVSrQq
sV7U9VA2yqoQrNEsRWv+qyKl/xcorzPMp4OrGxn2/Cq96SkqzGkjd1noJzYB
GL/sWpOfzNccA1jBSKpizrpVkcM4wVtPnl0BtdLSbrugbZu3DxHw6opCvsUy
cv3JXdvIutFoG/o/scopGcfsopT1Wd3byG6wUs2d09n1hWNiH8hBuNWcjql2
4YpEBLMUUbS/gjOj0S+4eODvysC3yfp7Jn1F5NTmbovbZttjSpUVDJ2VzykN
fInLCtFhoQds+iNmKA5RAtMV1ey+JX5pLMn98WZkqj531yjUBbr8PaRxldXB
+UsiitWnR2rYOxZxt8m2uRN6WoxRjLoS5vhmYj+wM6Zsh3w2DrHfczop9Vxi
4+qFebTjOzG/2S4x1yejqe1bAjEOeRd0LifA8wcYozJn4SVDJucVGRqbScQi
bkAKd3705LOl0AinsgNqeTgmNG+w1UmeTmPM9zXmb0ElsTesqoMOAXFinz+k
VhKVhE3WrwhmWlKZjTu/UFcRMDatqV2vRCZ9dNz5S6J97nHNZ98702SO3Zkf
2lq5OZX3ju8l1mqSYpPLNlfXOx6EMS+DJ2w/7DIz0PnzzI4Zz/NEUUMntOvi
9qbN7R6Dxwy1Fez6ADvyKl57BO0malkmpCUVGvXms13ZDgFcP+AK2Db715Cg
qe3uarsy8eTpWKEm1k27hfSHqa0M+zQDwRT3cgcDlpVN6OSp3ygoqNngsxya
L3S61DCUC22vsjAPa/Z5JrMYnbWQ6xWwZbH6dzNMgUAUWDekbQwAYuoJYSCX
j/5qWjDuELnPlYWdyDgzlQZulz2m4eAVB+qbUYinXUsS2vhQY+t8tqXPJAEf
ndhVxwJb8MjnM2KhXn4VouQyVSNA5JSgyjoxflL2otwZ0+yHUl2TX69ObO85
/rtB38QU+0l88uHjE6YzL1Ppj8sISEf3au9cSp0/fcK2cS6O1mOY47OhP7Hs
rIs4Ivrs0VndTyRbwuwJmH5Xu4mbINOtlO4GAXEAdkIvOgKbR7vIWNUmWS55
3RSz0jaqTUeF8YXQiKG3XmiGkZ29yfKxcaOaLSz9r8FDVerSCHTcubVShKDY
dXnGxeXPtb72EdjE4QBCLTmAY8SlmdX/R9euGXy4dNcmXaOS62sZ+Mjz59Ns
msK3DvRL9F5cvEMThHVwCvFgwejQdX1BDxWC0qdaOPV+UMpBHSRWOtj1IJMc
I18c6gGsUCq74OwgQphzsEuBJ/KDHbR5vEs+j1CYyDjSzrIEXnxKg4KYfMMl
4HCmaka2rJfQf/U0gfLLg0yAIllr25Fh40n1es8wZYzsw477nm+7j2bFptwJ
G+6pdrqhfOmk1S5uysxa/wf4PCJUkV6f2nytX0fLI9uZq4nmfbPdMiYwDh6m
f+l7pUsDoLTAv6LBZ2LMohovx8PjlwSoll4cSS58QDTefHR4Hu3Y9G9tCX2B
bSebigKYdLA5WL2KsY2Uw++9AEYA5EjbA2LzW8gDZEO+jFmRRp3Dt0zWxpXu
DDTuouTwbdRq0F4BeSHiT29H32cJUIgwRceEYrShwI8UzfVw/hbeKq70+fme
0THWczPkXb7kN5lgzqkcEo/39J9n9fh7VU5VW0GsXWQJl0neBSHmu7JJT9Qo
sdRzC7CK/Q1/LzCWLyjNu8EuO09kxfPt55HlF4C/69BT9UX65Y4X6SsHQ8wp
gqyJvYPMw+nT/6imsOXxfPfh+B2cWcGZ3EJYK9vb4fCm3XJGG6sD4Qg/iiJK
z/EcoluGoS5pMd4mTnxZ+/Tx9GBEy1uIxEegYiyZ7/zWcc0/a4NGSzHD5lBx
1RtGpjIRYyYk7DlwciAdVdpHm6dxqBJp+jmsY7NfzizRhCoL73l6y14ydqzA
RyD/qbuYbfoIMbJ8sIrwiZhF6GnigNbkiriRo1MtNBebteKxAWXLZdLMnvir
sO7IEge6MvoWmXL4SrRiqT6lYoqPSbMdc4tZwwSdL/Nyh7qk2wfCQo74k3CZ
op5VUWtaX8nMiy3BgDNWbWWjNk5EACnHFZ6pYzJwjiv9Y/a1sr7i1e64/p9h
TlrHjogmhuae/RTvK4+BrsOnzrrYWr3MZcrFbWgmJgZq5vVZdi6d1zLplq5S
5c78+U825nL35TJ2OMgYk+W6ZVBKgxBliquyr3n2vfAE9AB4ybrW3oxnoQux
IloeQzQmpfFydr70HGDdxSPQ/oPHhUdEIW8v0JOrO/rJM7EMRtku/4RskxWZ
HvmzgPRwCvcGCsSAr/Fv6tam/3088Ci/0B+4w6OacnaeSRLKQcvej0n3gLZy
XZzfv1bahFE+NdkAj2PgbB7CPSeh3I/L5vwnaN2KjKzB1PR/SXgBqKGE6fwZ
40pLzlRKSJJneuyrvWftxr2CwGFyG05kpC1oZ5YLfQvCOjZc+sMZOJeYew4T
C9Qr1gEPAx0G90BulgS+KlEs0XdApuoEyGfys5FeMOi/xdjo+rUipWz3HrSh
RZblyPea+IlDVx2nDAlz0ngeuSNgoAjzir+XwPUpuYCCnNkbiTQugLWJFLsa
ry39nxTrTIMRjUC6xoMXza/eczR47Pcgrt+ptP205W1i+BfqRhqMQsqvqYCJ
LALTpMYXuBr7zfOHFwqbiirWoHIIvNbsD6nOooq53mR1o5NX8E4lrDyaXDnE
28vLRqEs2vZwfA4bo1ZYIHpAeOjbEnsFrrrSEHTaw1X8I5DtbetpSQuTyklB
2de6Hw1nFw60sPr9vxB4c0XLXrnpgxmEEy6je83WXf5Z4UFbLQNuJ9wS/1Eu
7/qzZMFhAjRhOJDrz3NRR/oh1zzR13IfhwdhyTrS3aXTL0bpGbID5ufBsLzG
E2gdVGlWAkQ28xVOqBWZPOapGS7yV+vWjwt0AR7lP5IV25WwG3qH9QmWVDsR
l3+fD7GwGkAhMdl9PynrUBAA8dAsNJrve9hEqK90lereDe0hwOuZ9dFlh8WW
zhIhyVmo41rxAR23MTvdxE0B0sjW2rr8vT4GqYLHcJJbS9wa4oOmxuNUMghv
iSET/Dq0lkfrm3btsQnFqNXhsEc7csqmDSIQrbKG8Ur7pogcCyVCKxNDo3t8
vF5gKrIKOzL94EtdKOTkFDszQbDcRLFqa6hNO+t38dkv8MIRyeiw1ID2Wnot
ZWOTgN02oOFNdrGYBBKUS5XCcE3YWBs8pNqaghCwNntCUZIHkDWDo/vMhAqf
Li2dJJyvXtKkTctTbJrfkiK9uZHdZ1GSIoxKGPijM9/cyjLxFBrOEGdPbdt0
Ksg41RNx5W7hA7cQ397TS2cHhI2YVOYuDXqWNa6eBqXi7d12ckwugSUoypPL
GjYQ2PXeZd5M4p2QDkee0+2TLcBEEvJgjAVgSgOh1qbPpcqqyTUTVcveyOKa
HZxmcg50ND0q1gM4otDRlb/WrENLpcmshvRJJe/h+gP6yEx7rKssv0gduY+p
1sMFQp5fgyhDJi2Sd2vaCMY6Vaww6hvbNLPOJOstB+bxal5uwdNgbst42X1Q
rG0ja8O4P+oEyO6mqE4Sd2Qcoi/AYe+wJxNDO6zvatsTM5lHoC6yMALbpStk
G+u3vGlgD5OWlYKDC0BasnyKQYrJ6PTfVVZAZK/Vq2LzH4XBAseTe3veqmVf
+VBMODfEfAaHsundnEiR1WHT7hjnCeg1fbLkRlKT+ez9T8YuVeNNIJO2sm9u
sNIP7Mv0Rgs1TfYrA6ZW4ylf3sYnLvWfJ6m4m8OlC50NY8Qq6ufGxQXe+pd/
w3Vwar4xdV9qXVEuvzL6QJQawxn/yMeRWFuJKuKj0/2vyZ6svMlqP2eb0JC1
YbXHh8+2NfqnukSgaQtI1MzbqlELn4BsrA3TPP99Y3b47HnmLxjS/LIAyYoc
HtGNnUlTpIaxrYQ6GUFfBAqQHky74bOgTu+A1dA0gxtwgOyf48BAS4rbYDVf
kes5lJaWzL0MQ8jhei2b8fZl7jDIXjZr5vCgNs7s7Qi8FApwyS/3am4lywLu
+A9kXg4nSva02YGOlr7+iJ2pHP/sdEVQ45y7HuRUdJEofT18jle0pB/03eUV
8HVbzY76PVAxkfHyZH3OsGbDSGzUYtCGsH/gP6+Xa57rbfn7KjrfFn1ChGkX
GwsozDy9sQ2PrdTJPhH1rh5ansbxSwxhdHwozMDPI+ZfgzZrqFEyM1/g0KSc
K6Gzlq5jonLvMDSl4ssYwd/vhiso98xmtly+TuS29/Md/ix3PoctKGqRrAkc
VVKnWmOSI8/ehrXBotK3rQduXUXazdLEniD7S/yUNXKgEQsAyCOxX/AfsonR
mU4qLOksUCfeXc0a7wTToD2JQWj6f68oQqDMU/4UGemlRalmn/NKXU9Xidiv
8gnMJgBDZn5R5Vv37pPHnifIxI4JcrkLQaQSvdK8/7oFzubuzGAngjOGuIC8
IZufAZu5obLa/ZzqrXryszhAQjW3rfOeZPJDIEXEFscSMXD5IoZjT9WUQwjS
j31v0jcZGNX3qYdGo9cs9cG01B3bLstKI2JOcTRxQEZJAg6drfZs0nKwAiG8
GMjDd6MI1tNu+Vk84FCFxNjS6iwy/x0sHDNikXu7PuAjXYJ4QazkxEVRwtHU
gwJzMIRHwlYtflJ8KxfLwLREkE3PovA+7kNHnEdmf0vCh4bw6F19+TT3GWyK
plvklTCKyo05L30S4LYBIbzcRz5H0m7c6qLTMWC2O6YRtjXKdrTqiu4/5bt+
aGhS8pwkFTuAPLfwEKhLtFkGIAOEsWesD+dxuk9KNcKJnPMACFGwBXmcF4WF
A+KZNmoFNOFPJXHO+k03p6H7iet1cmwrGwlQyxf0Mz9vknYkgv1KtHYzBw4+
QJITAkG/ILYdD85IVJOi8jYecuD4/Xsv+p/BKdhwTI9HxJQsh/vKqZXFUjHw
O3U7697hoCDWROMfb9Wr2Z6OwRFJfg4uVBE1hkRXHxCvEBMiApl1EdBIAOIg
P22tHDKCqIB20gRIb7YT8McSWWMhTeUppf80OHMcbQ9eHvjpA68KDld+Cqen
Eza9XeZ/aJ85Si3Dj0Lj9Hx0YsmM3WKajlormOdk7hZKixCLijtM5Trlnv2u
ccwFCO+zN7z1PQgp8B5PF+uE+MNi6fBPrC8/ea2+7t7Foj+C2YKrzwpJdi5l
mjX+fM5KmahIG1azBrWk9idgh8rWo1X5Xu2RHJB56xlx3QOGfDSm1CtjVpYP
m66XFuidMeekAh8v9JYVaUdnFNQvo4SCL8gQ6UW6N2A6VFaV6HHLKC5ukimq
Wbyr9CzDSl+pmn6fk9/WjHkM6oi60edeaZnb8wDmPjbg6vV4xqtQk4P4hnFr
rbOjoQf52mACUR/0/XnaSVINl1mv98Xuf/U+9QuqPvo/UNRf85E/n1eaSDRa
XI2yGPQo38e5b6CTd8p3MS1rsggtjFYkjBJgqWjQt/a06FSxj/DeD+V9esiL
nkWaPVbdvfvyQKwINS2uqyOUugXnb2355opkehmdEdB91huwB4xOZnU6D20N
y/d8RGbB2O4omBVDGUXoYodMg8yfftzRXWwdTv8m6d4m77DTghMl3srOtg7C
Fhb883zFGQPee2cV7rJJbS1Y44rGIp7w43QKg2wOBpX0NDhSSPH688btz47u
mS7Zun8mZA0SP4NkqRwJNUkZw8n9cneKj3y86hB2lQUNS7RinlOPXIv10Ck9
JXrFuxZSGjuMd62TwGOK9rgBGzcovcDvuodBlV4rYVmlG7w3nTrTod1pxv8Q
/EyWKGwqd5ZzWMuxQ5FFj4HxNAHYfOqJffxm0o+MIlnTxkvepQZPPienzDAY
+8hw+wD2ZkgAA/EKq3rukruRlO0QOVsTLFf+RzIK9tqZNGfegbGsmK5VbmNP
MiGWmTzjwNuU2E/n4Bc/O4fV/JsZloYQOHhssCYZk2ELsZrLiMSaQdqQjQob
CSGHd36ubwZzlF8sbEqdzvszhBXOOQIqt/OOPTTLgV+6SPUKBGRxY0LUzB9+
C2lSDX7Hu5JLSB+akvLH/dLn8tuNxjf26def9BVRoDAT/FYNSAOLqfVVoX9B
Xl08a3bF5NHLbPTprh9t4/cpn+i+3WizeTNGk7XqE8cvWfUYqCSEishcwlHA
NHSQCrOv/H7sXhSBIstogjAQIwUceG7EWc8yr5iqL+w7WVqRJeh6lWbtHjRq
X7wWOYXB37j7xwohdV/oJEho6B7+DtN337W70qa/maDyVsiOuCULHZtWdLuu
LXap8nT6n8lUsyF1aoPUqPuJy55WdSpwdPLvQIudaiti65bwl7hIM2dQWbf8
YMzit24YVapgsjeUCNpq+6hhYrF2oO/HFos0V+v3pKtHmNgypCmRH4+KxQUQ
rEethiiHiyg3XIM1MNoTvDpBQBufdCbE7QSZvdF52VtohpDXmx1fxuJ243wu
bYYcPOMO1qdFOI1O+Nm9Tiscp3B7OlRVpPcOxmgDeIg2JoruJuAECm7OsSCM
L07GKl5UZZT7bmxj3mOGnIu/bDP3WwpRDMEwVxspJujADl91+HtcDlcL3589
J44aMS8kdK2loEw+jwt0yA95A160T/JevK+AtM/Uv2WNkNn2vXGp4SrOQDsm
A98bQBqTdQYm7Iae31bM+y5GWnQDpLah99ZfkIemTaKVb1rDKtzgK1zmdb60
NXQGH1nh8r3CMN2Dl1PwIRn7GgawBzsGD/3CtiNqN9ApQ8N7vckme1ksyfh+
kpVQXym7Q9CLLdVePWXiYawgOgxxMiiZVMgF9BU1pqofzGi3WQw60L58RG+G
WhiUddL+yvH1luet/+WMV18FzfYybfBkcV/gy1sgCGiUrW85LBoqLoA7xA2j
o1HgfIQ8MsPY7PvzaqmBUgjB0XC+PouzYHrPZYoLac6QHFPUjemBVVKZ26ts
8vnrmFKnO7wDcGeN6xbnUHzljW4Yc2hNfjo7RGlVK+SzBRu0B5eBqPLoWzaD
ideJKtLnGgGk64ohfRXd1WA/ZvmosTDXLcsA1ZPXT02/WSYC05sXnJtY8oY6
+lh+KJq5YwQrJtn2rhApjchjflhpud9T1DYJA2NNLGf0Vj2U7YGybBqOaKG1
Ym17vgRUCRx2oS7Tj6k0Oh3PJTgPceQX68yJ1O7bWL8W9i/C2tZlYhFUi94l
oFwN1QEnkUHIOiuknducjxNUBYnfGP8XPK0WYd56PffWo+wMdMG2W4Tq7KAR
++PECUkhsRvgNC1H7Rd9uo9wLUaJUHpnlMsQoZNPOr2Yb5rsdcu+KNJpF7lX
qXsRao7ptyl9JS8mIFHoaiysZsQQN8oCCQiHUAiQKJzx3QxEi2UVfo6yjUt6
K4LBqZ3OxIWg+MZYhJGNyveN1Nl3zeXC+fH37wUa/POxRbkethy9BunJGhy4
hcLwVGfa3K+aHse8o1fxGNYQStuYaF9YMfm61KyQAVKNBy/ugzrQ4fTZATYz
7t71BOLQ1x2U3dx/7tJzZYpxSPCVO+TYruPZRfxkiuAQKYzr1aLptGCL5d37
wnCsMI4bHZDkPeV/gme5EoUAIq9E9ZJEa8RsADSEZRgXzFYvFv6LbK+hsarL
N7ramCkKfbfUZ0Dq6vZyTKHK1quqXmkJGWj7G7tYfp9OGJ4Zc4Q7e4reuhr7
zoEJRT7GOgYGn216cdA9G8vhK4w4oN5sXHyXfMlkWnT5cZk3e42zPptHVEdC
n+S194RBkCsuaovJsCy4ObrS73TX2QNqfxS1mI6K4RLpZDgzQNiy1E9OMS1G
IQpeskWYs02/y2wkvhCTXlULOc5MjPHEZASRTGQNgTrEpU9tBTMbhmcODKUV
ETk2RNG1ocXVxyeAWd182yREhsBR+73LNiJfdFMZGH+XqhDNDOEo7IUQJYJY
mr+LjY6+8hi0s11K1Klhi6qs8zV8HU+ZfPB9mrrJCNJjTeXeYbnAl8oHMRdK
8STwHvJ3y0nQVMPR0jQpzLXDZ8OvqSFiIUfVTluGpyvCQd72txqlE851sMdx
qNvUdsnS4B698k+fW1yE+foxujdE5wUaoESq6f00XshrBRT9DT4RoPmt4snm
vmrkptOojdPjequaNA0iCZsSYR6EhJCp9GVXGxw7Hut7FfgsKG8JJmPiUNuX
rZQKr5Zs3CPmTf+O4HyoBcHIsQY6TWWH9b6buFe6uM7V8Tr7kU/spSQDJCR9
ak983rkGdZDNk2LoCZbHtkzZJQMgSzV6145wfc/n9FVRFFFch1Gxd57Z8/Ib
ESMvF/bDj8JT/nVbyILdCZNCwsF9HWVMttkGbO35eADrjUlfqrHPrI+P+W+B
THgrtuj/rBY+WZ/cMuxn6LGcAfqPlTj9L30XiLet4hMJOzki82fnarkv+jDJ
6JZmR5k4D8xkzKwHl+AQj4NSy3DMroOSKSH68wFTXY2yg07HHa8ten6J7fZV
lScrIgP8nb1GckNSs1wg0luf8kwzBC9SvZLVc+lJkHp/rOpHugtwysv6LxAS
EpZA68o/uof8v8LfFybFmPyq9ifbc7+XPO+Hu3SSjuJGVjfWiBhAe4OztogH
FvlUwUiDqoIjOhi1vjKHdOAfyS51Qyly7c4DEBWd9fdJ/e9CeR4OQZtxpyxB
j3ymOKu4zWTlYPpq/DFZFOFY8lctzH0Vn4CMEvQELJvANPupKEz0b/9Ozgko
MzCBsIZpIOZpawGienXNpcoD83GT1Jb5vaQOD4GafuLlagL3AfJ9e7PyUcka
8CdOTYzlrbG7SjPmvvk3HKl2VR2a8mw6CaELjDmpA5964qFJW9hBNY6+HN4a
y7f2npz4rHHKGIKOVbtpn+vUug+ESoZdR4AhVgFzkGxrWnsPQ8J62Zvg/yMS
3N6zfaEczw+lQZz1SMJNPt++ARmkKlP135ZWSSKNbhiypnbD5AtTjd8cn9sB
/3s2ru+7orT8c3KW4Iix5lW6vPSSnLoDc+rkOyo9GsqSSV3C42ccnJ3s226t
iEQQsGJ+6nL7g3U9cqJ5AGxI9U5SVX33xBbACGpfgmF1T/IDLwAfRQv0egJQ
GoQbllGw/WtmBa1mOlJ24Aum33YHT9ZivLIDVDoIS5YzGItED4Ui6O3elEjy
L5ws587zmIeUVUE4ydK3JCVGyIVZ0ZGb8PvCABVeVeuC4iBGlqjBPNy6VFJ/
0TmqCXh+356YwY9TSLUDB30OaYvj7h9IaZYWND3tHeQWZk2FY/xusn/erGMS
gRWzX7v8Nldd/kFb/v/sjsAG5A0M08ZbjS32mGEXzwrUJD727gh+IUSsCtJu
oGAKUfb80d+5ShzVTR7t1WlJWmUCh4LpqgIasORHi54kKh0s8/zqxYIOx9I8
lXBButy6mORLm9r894O1FwryHqb7sz26yDhPufQaGl++itqImpVQBAV6tD/O
/8TLa7O1ZNJp2ZrP8uHju3LtC+3R10LQHXqTowyZwP6O1123dcRcCmSxKp9G
LSdxjeZqtrJnLKInIfxTTmJZMypy4/pIVfqVVRlo0YXgSmsSZoP7L5vaC8rj
9Skjosd0wjbQGhnppiXiCI9cG3lpATcDIq3zgBv5JEwfqOcY3PnrrmulDZKn
XscLZlRfdU59qSL3h6uEotNYt8RTTVH+IomJodWE4ULCZmiB/3BKw+TAqvgI
Ur+oUUg+jlm7+sCVpirxSpNeeJDKiS2luihMf8H6Uu3Ekv8etli2e6vdg0Vg
FYvhP1KbgDepPiPvuyTX6CwEst8DJI5GvaMksO0PQkK3dO6N/UzSuOzGEmJB
EIWhSfDuBX0At+E+mTRNeF4ZaPouM/UFgiDmSonhTK+jxxf5v6AN2VkZeXfR
nqm8lF/SXkq3vsYvAL/+Jd0DpWwoWjVBL57SPr0WeS4r1jsbh6Jav1U1P7l9
YMwHrBsDIyflLVMI6vrS+pVg4n88kBfFNjtUASeLfWptCov1CY1Qh7N8ZJ/e
+Uz2SbOhf7iaRInS0k9Q7549b+sUaRS0Q34GUqZBkk+1olkirmQYNJeWk4Wp
ZgMcST3zVrEJ7B8ViGzn+vEIeRL7WaeVa/csHyls5dptC8JxX2JiS9FgjwOG
h+tH7mePzcgW/lIgQvWG7MCw7TQDKoFw7oKf10F9/sYUatlClQo5gcSPaV8v
9Iiho07kxASgjkRuYS0ZgksPPCudWH4p4y0Max6xX1Wj9ePe2wbkc5Fdp1Jx
tDiPc4MKraXQ4G2Qyc7fFN+XnpI4iYCiicI/BykLTvHKrxynryQLtrZNALze
LAUosD0Yr/5ZCIBiZh61PXIml9Rhp6+763iq5qAOJmHJxdlhZWM5rx5vnwOj
RmspAMtcYE+5sI3ycJjdNJeFx5EVd9M53dbo5WmZnkiEwMckVfkktmTmY9HB
//CkMwkJpq3Mz4SsMFmcF6BgA2d9zSXhEyfOhtLTUqzohE/Xu5rtpPNlNdJ1
1nebn/I2Ldx5sSqG7rJC6Pl+2l0wCb006Nk3Rjlvr14dwF/s2VWM8MJ5sxaV
6xNk9OgkRMmTJJIoSpVlr/rU0OV45KwzWGDjwPDY/hzXKeGh5PkobgKYM42a
dhfsQbYzCHcDO8fnq8KRkEl4883w5/341BmRkdLSoOW01PJE4qhdQC89FqxH
rf68nz6s5moZJ6+S7szHHcMT2QD5vmaz7iGxvGWgBtCIsxv7wksMPet8pllb
Wy/0FhoclHg5WLPLR95ThXop9K5wC3IPjjgBqa5KCC7lR4e3VPCtc0kgaQb+
/v5OE1md2YweM8mJ67CypnpJEJ+eKXPV15jexsZNnrst9JKgFLZONCibYMcA
r2WC6WGBiaO8hqCwNJ2ywkorRqfY4NiJBw5LNfIIjA/z/LmOsYZ4nPwvMqk6
vN/es4g8LqVa0gQfg0NEhwrM6V0ZLLN/VKzD/01gMIjr3a37K9qd98AqByzo
CWaUdEg/1+BHpeQiqWNaC1CYfz4StErq4wrjH4BDjtIT85dpsrBCnUqyo7AT
05ymInMc3RGX0yND36f7k2beSmsYU7nZXalWdpJEnpN99Z2W1/DegHWmwt7B
+UEgsJCM42AM6trtnFy+M+KetpvK32zdWdYv2fuqor8xAykXMXnv0VPDSL6q
RV5uM27jFv1XvlGK5MvaJI3OC77eVIzvw/b4hxn4O9YWOC2NSoMPBT4M++Ka
wdon/giSCQx4x6wT2lhVaPmHO6dl431LMaJxQ2HGxBC0VUFS/IjoG+vLoGlt
IHQRDKX/WkDgLjwohBBPBSfgxOMEbgW9XExMT5ExtHG3ArrqCgmQhk8+/YsZ
Egz4cL1zm3+7m/DvjkWv8vgA6Y73K3j67/ibKSraOFTabjThBpdlSrLcHsiQ
dJxz8S8idqrL4ynxRC/410dYMiA1RtGjTUeO1g0I8aqQUtkmErnrPDLi06g9
i8G93E9jszz56JXUq6cBSchhqCOnXkqBNiKb+gbQZOCts8CFZJ7PqnT01SVj
bP0q6kNl14xmH/x9cfx6mCnpbrJ8HqWgQC+IU+W2FdMJof6yfUG3H96DFico
j+WgfffoaxxrkW6u85R9UoQ8BBE0vTWmjGxc+aHl/+e8kprm20lIfZxOuKJN
CblDnNP9WgsmiyFb/tZ7dwnplv03e1SkR0EE3rrPs6gN9BNYy9gJPga0t553
o/UYBOeu9OzcvbpDgzDSpRttPkuM9MjrbiyGxPkQWM/Cc29DwUvCHX2s3p+s
9r+A5/sMDf9j7Fh0bsdtsawHAoIVdYq3IYSJAhLqwElWPXbWuoXCsbKILIuf
S3YeF/3gDyM3Tl3+riyv7GsQfne5/SWEnGma0L/JwhuJRX/ZGWn845grInMG
cA2Piq+ObUqMGEghyYd+0GaJSQOjUGaP2juu3n2aYCZzYBTHqYZGBmAzuv5X
enAFntw5zBq4dye8OP5rYsehMiDGivNHZfHhJnopfmZ8Xgsy55pIDppNQneK
fXOGpTISyU6YeqOpmKg24fzzyvgbeEndL1dihSqQGbhFnYW+IdUekuV7VNeX
7dIXoNeoLhk/ugwOZBWtvaXg7/MiSrMAe6H95vDL2QMSWQueGxT+hOw1PfWx
8rQCHIUStH6xDIpPJ405WOsIRCwCHUlfPN+5XCVMYrk1hbAZ8iYGrCQGiXRM
yRXD1WHkBALMnah2t4+T45xNp38+dj0xzgj2s4yu8KO4AzOb+VAcH76z1nLd
FfxqDzZGnzhRdghkoYQQcMk3hTr9NG5Cj6WIVxqXtmB2uLN0mc2J+UXYmWcF
UUHOjYExBdYg5c8wSUWMi0m73Ju4yTb/ZXT285MSivKKyyZVMCN0lIussBOw
NXCkWUvLMmzMTEJ/Zut82SzED5mEL23soNr6RmXrdAhxxAKsQU1SUNhwjhFM
vNmLTdls3V8dJ/hVntMSTni160/8QD4i/X509LtmK5WWffP6lnwWi5N+lGEh
ScNUVGUa2nCHpGHAJTJgL6GhF0PWrH2MF1P3I+hE2twWaYoFn8qnvDM9vPrx
K81l/MbCyYVro7APnbPstUYGtRlAyYAoOoar+6fCkBgPfWLvgA4F6VBO1Rnz
GisboCcmaAn2pJDBiA7Qo8mhebhUbHNTYNFfQ0dNLxZ08dir53X75299yB86
r46iw/lcbOORIeUKgON7sPm94556MzAsA+ch/5npZGJPzeZh8e2As6AZO0Qn
EdIR1Agbj6Lxhyj7KgGnBvC6fdIzgEHMXLqSJ0DhUhbW14pvCbNnWFgxfNo5
CGlOErXs9jGhElbEUj87Hxxxwk9vOEhQoLGif/NCgn5QjI3gKKVoEyNAT8gB
uepiNmGQgBDVftpahFLFoVevpXk260jMSUIuksVGsLF18GpK9lnHRf6U32KC
bb5o5MiXrmdkKjs5tp61o0bxJxE+47OIRa76iMQKUJQdxZHgOW+7uvLBzUMd
ZL7w4B1OY9Mvvo2xUqOp11rO34N2jOyAmDYaIQUyLsnOZLhgR+rDp/q21MtE
JJiLpscyJ9w38K+txUtcO0YgK9iFVpdGgXqRR73U4c6KpfLJcdzaUYtjvDwo
zGIXhFD89p2jXxY7+j9JMtaI/bFslU2Exb+mWYUo/RJTI8Y9vHjo+qmIYyA0
7202/F0wi/DHdOm7fm2lWQabYaD8owiDmnZQTIKCJeQ34W9IpLaj/lAdy4g5
jHaDQelx2wGbyPEWEP421h2D1lTrrKeB2VUCYHeFZGynCFPp6B8wRcDXdjau
K5axSPRDofqkw0Cy6erny7IYy0bvO7P9IU9uxdI2kqskZUe9vN+LdgGiLt0q
eLvTHdVkNEd87Z0BkjmodDjDrOhEShXQqKwhxoGhf8955asy4KbDtTS+pihb
Z1ONB3H1TyPdtWt5fpoH+A5vkS8pS2X4vsnpnkQogihz1vLUeFU6oIKKb8eB
cfgJ0PL1KHI8BsN7agd4niudtChiGrCllSPPpy2XEgN21y2t1EVOAa2PXC2F
u2b7ZDO7ZiTpLEwP/dpZFjL0PQDk8s/zckUM9YUY9E3gTsAAQTr6x1mbKRTf
tk5mgBI7xSWpXFHfuK/PhcL5xDbkULPOCNRxeW05ysJgjrasA4D9Pv9jVIP3
vf1ANDeNGgPC0dPZfKvH+VI1sfcgxf8kC9vTJ9VWUrEFrjorAPrYNnNmbhoM
mpQg30fhGvNdbGnIoMY3dZ1ATqscTge8jF+Rd72d+AtEbMgiyrp0HRlHntnx
FYrDETn5OH60go6dnNaJZBUf6+PokeJzcVeFXMd80rTdd8M1r5zYseFf4psn
gBwARfF73RaKESorhc+GstgnBvml+zLoQ9ncvHhhEh0zwgzROOheuFLQMwg2
86tVAN5h4ZKWp2GUFtWyIgAKQMgMJJle5odlcKMl8y5NMEL44HK3z9khL3Fi
Y6DuK0yGxZQirEzbrWSo3NZ6MErgZPr2XzlP6SnYh/AaiL6dDX9DylaB42Mb
e3wg7PJbEHaSo+kdXDMzRnoM8VNRiMeokKmNOUVRgXLNH4eijv4IToAwZsN5
rlSv9wz4TdRo8q1y3Py3fa5C9M1YXKAPjpkbv4AlweRu6XRgwa21lF4A589l
Hk30lwA31X/Dk9juqcc5Hz0C8bfgaD7SPqxCkIfR0h+IbcD+9DYSpVpdBsjl
w/ubOg35EmRjwbUrMPvwRef0FT12Zj2Lms8hXAdOAs9/LkWwSV7fEXtoMI+x
FNRTHigpQtWWx63lW6Cv+ahrOeaQMST3rPzXvKyBwqDDezNuKApH2N14kZCW
/+4MqLcjEqV3sBsn+lfh6S0fAGQZES9R5EmjZvGrkv1vP/m4ZenTu+AEuJ7h
nq8sMDwEB0yjZ0ZLwczrqcituj3QfEjXduU2BEzCJ+QiLJy79CATSfPsaMZ+
dNYdkeGObjPAkhvjoKoWzOw82e8jY+P83r2ZN3mPqEbuQ+mYgAuVPg2oBDhP
G900ClyIB8U8LQASojLkKnbXPjtkZs0MrHZoWodvRQtjWZyWsySNGYYfHUsh
8UFJyYMaQh3CmghTDxwikpIFPmc1ThkWH2TH3hAoJ+0SYVSXo5YDr5VfFX9T
DPhU7otBL2BxVkMgkzh8RX8707OOJUcYgo9xNiM0zhg8yaKkz2dB+mFVRgGf
bodyroeUVp7KbQkXMfUcP8Cz5jRE4WFbt5bAqeJ6Kq75p6AHxFLoCAI6MhdG
MnXB7Ag7s6GGE2M1kNaM8x5yuS2EzpeMT5Ak8JMU2d1qcqNFaPinKiVdQSN9
+IZS20UqaEntAfwek1B73a+h7v37IzPjVBhnFUGRMa2Wl2zAQ35OJeBzaBwY
qiYWm0QKzI3IeB0rSs4XQBJ+x0cZuJdB9a22HVpeb+bCxZajUHPuX8RQ2iih
Ns2L+EjBr04SzaYcMuv5pmaFAM4UEA+BJaHrDAFzeTmCdVdhZbuG4IkLs6IG
5nQleQoySM8sflyo+TzhXEsXHdOtnVGSL8aoYDpge7kGTDN21kGaAfJcHDZ7
ARgCwtk6a4C/dKnZlul5N8w8NTTeWxJkUBD2wa04yhuzKlSZsO0r245jXqel
7jfa/uJjD2A7Y8QZsHuHFhL24WkwM/ZDrR7pAYlgzMVqowC67gPBsAtRVonx
mSAgUt3LXdKNthjmuZdbv8LW0MgjLzC9Lg71wWh6FaJ6t3izOvYIxHrdIgUv
RpH3jXzSlhmh+Wa/IjupjIpg9o4l4RA49ZGSlciy406bfkMNPotPQyydvT03
bBKOVWdYg2kbitwhxa5sJnRIhXQRtRxd21hu4OMg/rBnonIn8YIeGzU4/TeU
g1CUAw9005sHnd8E0/qhfjKa27BsY2Jtw+Y2hE2Eg2G9v1vQGFtws8IWliCn
IvexOnqe+HtDUCNAcreuJLZMEz7riJVJxBCfIA7+MpEGKcRMWfR0oq85ozrx
Ik2NKROvPjTPtmksp+r9a48Wfyn6RPXvJFq7AScRIRmIdTt1BR6wcKexgwg+
SdR1b0RlvtVnXa8VywdZsRaAqxb0N+qOIpbox7ciQNuP1n27kQN20thqd7+z
vqzXzp/pKpGPou3nehjhCji2dHqNRKSO20DojNnDwIimyjhLV0UTKsu+EH6U
HhQdJWloISrE6X5WhnoE4S7jf6YZQtyY0A3adb2zzEykvwTy6zYBikL+p9Ax
I0erIv0p2GBpH82I4J9b9FXDI/ycLPTgIFMe74snxbfdZQb9SqkgfRS1j6Ks
Ye3XtwqFnpfN9UrbQMrKmUIELdUHMmAo06avZ2o6uBA7ePXOUBxaoGdOzf3p
sKARr08hiF28yBA9FPDQ6SyzwwE4cTPN/Txoqvab0uaqu8ewlynu4UZsANxU
7mQ7nT1oyX7ERniLi8Z87GRAgXMoSwoWRRslA+VCOY3RaqO3Vc8LjOjPa68B
YfIAWtWDnQXileB1A+DeMvQvaS2rOVR4g0K/Qaa5UA6+Az0uhwlehlnQFw4B
OjOF/2jkZbtcXncZGdv6l2G5ACcMjRvGoNOvuNH0l7ngqobzLP62hPlqfDxH
qlWxtC5OQUFTe7c9YQc4Z6Ge7b9L55gf8PGNIm1NBbhZipzhqP6sbjmj+/wD
VnnqEc/niS0oTQBLWADLFN4YEXnb+XSk9VG21E8oKIitOP8bYh7+VjEs6ySr
WHZAGYCqSFDkdxu6WxOEoWVKoH0YPMWBcjVzagbEY/lNnk7ERaiU05J+Wlby
7FVv0dEwtxp9TdGKdRRClxfUcoq/cOC83NeOzvr4nUH3xpzWMlktD/ntGe6L
ddSBMg2JiaPoJUgNAUU0nvZAUE5PgTJNNxrQ4FzgWI96maO2S19lYNHRy7SP
e86qHJF4wo9ILgpqaNNQcn/Zv0ejLiA1f5ihd8VlZmR40EyHWZiC80WZROGk
lFhJIbQelwulcAkpmC13/6IkKsnjqiGu1ZS4uZDW5UOrBWVzoRtvRm7OzSnG
iBrl59QkInZqEgvXNj45T2yqgo447amNM8RPrwYxAmP3zyeeQd1boiiN7Adx
u/KUScwesHfEnTKZdkruSz0624V2KScz7jhoTUit76xTj8svmxfJC6JGhXIX
K0hBPyEc7aLTelhMtac3HgeXkQ6CydoIL72dZqJRA5Mugv7V7JIx+kRTw+QH
6otvgAwPaGN9WbVodxA+wSzSBuChvdxTPviOxjz+8cIgroHhBMensJ34KGDX
i2UaIW/Dy3MXNaOZgtWK7bDckCBRQbeuj3cPoD6yXGe1fNAqbLzo8T31+w9v
1b/mCarLDKbvzbSmxzJyD5T6tuyN0FnIhCaZBlJ5mK/odhRLkaWd1oikDCjp
GFpWNJnkgZxzbe8FoLXCqSq3GNcmBxaSPjdXMytxgZ/bevydHdoFHdTogAut
Z0o8XmS7OVFEZl0IynsNw6j/Ph4TXIozLOd08hJEamKx6kr0vhp2DuTOueYB
suDUVIbb5YRtaZkY8G16MrhQ016oRZo6A9w4fihTr6yOOgj4/WRBCwfx/9O0
YvnHsMi+QrjKORl/OmO+7r/OK15/+MkiECTDoDZWJ5gXb+4kqQQSTnhbdZ6k
ruOJ8WN59ctefKIlmSGjFncwrzTsqD6tWlQBAcWaUdkCJovMGlDsoKRVN5x3
auQ6QZ18mzMTGTtTEeNyMVPZiqsd3S3F9hDRX9qDG/kwAIFzRer5pCd1133I
VpDPtttmHSlAtTEo7JgaIp4EPcy0ca+TjDHcpfoY03xMWDlSYuai7ROIkxmJ
mHq3eZkFmhsKEKTy23XHNG62OfS/ITu0fm2CMQCepgBZ3RlHZtWDym1WVRiC
nk7430tgSSG8uU+Trf15Y5DZ9KbnwQ2e3hGS0zlNyyFA6c0b6wK8piCcI02o
f+GvZ2SuOVrU88AUQd2sB/pIXFIwAaB6LqT/OjQoYXNTHnCsSXrdKSAlBzzq
EyQxtqlBuUpfc1+zfwEZeB9ri8wEYONoh7OutYltB6Cz6m475ec/WhZnw0F5
0PSWIYtzZNzjUZcY8GRb8FQcCrfFR2IbvtayK9WxqpsVgMkWij+qOm2R7A7/
QlFkCfUsj0tg+YKoKnjGZKQHWTpKX3Tw5cH3i3VuGBSvAev32foZU1E9S/K/
o1W/SyxjxdP31fh2/Op3zKSTnQKBEKd1g9n8YXnxGQPsTJCr/ECQyu24wy33
LTCAxn9vMpE0lDsrPJzp0R++8pWYr+LpthEInTZLeQmnXjyKYYijF/AecKDq
Gl4etBTEyLnfq0M2CPlGV040jRNuIBxX4EJfPJJPgQLzQVE88y6bQOX9fvxw
bSLZnFfo95pCK4ThE34n2lEL9c3bET/nrygepUPD4CIpxPJZvbMOlWsuFTEF
sZ/Z8btnITQxzLszamVZxFkaAgHhINm5oPQJGGCngHFNoWf72COxDm1nftiZ
iKgKUKjNoPGu67BKTMVRgAfnGrGYuUtElY3KcRvaGOQyNoRIDU2tYurI+6sz
NJIaYZf/cOFhuOjq3H/4jBnzuQUN/bBTtymCjBuQbpBACPGq8sRFtk9brhdq
EV2T14abJXGGbnfWkD/9RDOLBoJrhsYA1F50gSFwFJIAB/hex9QCzF80TSJd
+ENFz/Kh84NWbkPpchFgCB10dzcBLIqFvfTNOkZ8ailB14hSkAKMBU7ptu67
IFMvv+6+u5vhP6b5RnUyPg/xgKcDpMup2URZctsNS8e2XR65UbSvDNsv93Mu
mihUwcfibxHUaDoi2XcN5iF6dceF9AzMNKSdYcR+DjD65OBmW6zHZ0TD3uBX
hsG6NRTzMy/q81FGW+abiCaG2Hkc3YQTtvhn67syoXgAzrZwK81tyP49uKHV
bnWOiPDnBuVJhGNZegOk546pGTylklwbNJldsgD6gRu0tCye+rfL93besYsR
zKXbKs/IQMW+2iuG/kKOi7FPDu4sOVhD0V/OR38lThfS/JgQO14HNH81g0zP
C6gt9FVYtmxgE+61Y6USsRskgNDZAIuuYdZITfoqHBOlyOhxOj+exmZAzT5Q
TTQiiGFb9ClvttgTH81fTyDZpK0hz/xfwFU3A4V/uh9bRDYDgP+/d01OmXwr
hhh/MWBsoMlDl9mhkHm8/zm0N0z+giML+nUM4qvKI16yB7bpsukzCQ+dnchq
Gx3LQqbQ/BhGukr35irbCMwpn+JlA5ud5zLOZTANVv44GNZ1hacXOf7wM0lk
Q/2mha3wGHZxXBnZ92hxZZoGZplO5afThd1eHOUrRKPicjF+9bHpfAY7Ilsu
Gv9bvcRJcKZPXhvNjr3GFBJpCrCHjjid34QjzHtZE2McHB317kZl6o/3CGjC
pA+2968ilc4bKUiwTrxLrBO595KKFClmZZ9ohTR63Vhkl115W/TLlEvfN4ML
rlI1fpsDjDAskkwx48TP2JJsXEyFB6vOSRIMQZEFoTRkZocOsMgFh3+XAMyW
7oTALKwG5LdcZbt0Y/V4BE7+Vmr+YXime40U7v/ukJ44coMBDvqQBXxFgthK
Of6VO7O8NcrzmMcZuEMJV6BIyrQCp9DD4Jc97g/Nu9KD+3xToQ62aMT1HNDo
OJDzKN936SpjzZhH0IwUbivd+9sD0OxEUZK6a2+nofnoKm/0nzAPs5pY0GVV
M0UTK1wGPIGpl3Ov0zdy7p2MQFYXXwlk8iRiOzRp7PatAYFJ4R6f2LkiOWdc
izTehE4LDca9siNL2VEXT1UUzJdunA9In2Rh2ZH1hGhv/mAegPzJF7FlLXqI
foKpFsPhJLeAqMCiSoNRgD3Kc4UnF0Adu1/rFUm64t2A4EX9KkgKIY/YH7hS
gsQF7jlRfWaGe7zbOZanEHm0LC4PcQjSl3oFMv8q1KN+IgMkXDCUrc76c+Z6
nQWdjLLuxyzp+NLQGdBYZWiOL8GMcEvkk+C4OsbyClXAVuBQGsKCg3M6/QdS
jdGr7PJLpuzZYV2oyDgJ9LRuDfoQu8pFcfOTsG1A3tEUC9gKcRbQIUl4rBS3
7fnF7NGujD0PyafS22hk8iTcKjTMsH/lx5TF+tt7bR5esGvUsjP2sEAp8YfC
GuEZp2KXa4XHR088Bh26DIew1KRigZCudfgfgsjkTJ1hZ2M2o929V5OlN/2G
Oq58ntFVSjMHlgsLSYiVolXznF/3/XOH83dg2L5WDTex6KZIlRBKFXmRNaat
DMBqXmP+kr+KxDjBD8lWBsvwHWV1aUdTDJcu10k+dtmJBX4C/mL7qCIxrY/7
gLsJQvjKMugf/NGGp/Y0cJ2GKRWT/X311gSbsmYBb1DjIejBfO0dYWsxlqKY
Sbgn07xyDTqyRQT4oKvFiQ0CrTOU7dCNmdegJNX+YUbjCAqKYmqwVZJwpqiO
HBHt3/sjGCCRzY7EPhqW2CxOcsayaIT4/aFQvJCGa2EROi7qwAQho+07AkA3
L434Va3vrWuIFJ6McSB8GOVtbMbGR09gQdTuXU4c+kV8NssCkH4bc+TzJvzH
mNl48gYBOucdo1iAd8j1gvKuBnEze0RoL+fV/qg7GCTTdoLDugrB3pOneO0u
zhnUUcvpsfxyzCDEtVT58MwX6jnToMnLLzxdvrmaYogkaCkSAy00euB1u7+u
WgIRNbiUjMPTgPYJd1hH8BzecYNfCGsGbC53Y3vylxw3WJHh2sHAmqhBVPxM
WT+QgKFCz0wdNHpmjKsyJLiNPBvaccCP100vVFjw9cdum36fckyRpYHXfc6j
83RTwn/GduhVDlEW/gnOr/vHroN3FRLIO7Y8yY1wFN5y2CYrVWvFTVszvhFx
/mIKTY68SrjKj8nJiDmi+7LEA4aHjUIoHW43nhRfCHIE/ws6deiHju4aPENi
yDc3hSdj0Ycj4HNRJbNxCyROjNJguwQzVh4iMOkru960WZgNmiTw+KQ/6vUZ
9+30cQy+tJhFYbSNrcbAWstlZRj0PG6GviF2FUFmOx27koxNqkna3Y3tSMfP
/2Csh8NtCBzC8UBuVWOgDA35MIhgiJIooT1uOB9dbWZGx/Mba2P+dtTaC3Mo
DzFKa21j67Umu+l06f9FidS3gr0Qi2pNus0ca4TqZrRbB98nZUd4OkKlDaCq
TPJrt4ybB52PNmZQJW7oRfdEDE0JoMskZdNLJxs4++IWwpc46sBLbGRNbxTJ
xHWWfZfMEbIZZS80erTH8Ht9HPESPiXCN5XrBkIVoPfmm/+nJE/FM/Dw7tON
1Csbn1W/+wCL9lYQwGgmRpgocgQ8T0t5QxLwAuRUui20K1vG8caX2wSmOJN5
bsSEwdAYP1pRlQf4UY+866dLgsDFVlHHgVG33Nw9bXzWf7BpWlS4vBtD2Q/E
PyaQh9tk6MsFU4XW779+GTb6CH0ZlZgIWmPoBJL+QGKgaeMgv73OkA38v0nT
OxYqh3QUpOTkRVBwb/7eDM25ywZtIHzzeuQUFJSA+wj1F4huDrtwxpcBlgaM
pzr1iodkntjKWo7W1bL4iXSBgss3KIpznQH3FoO4ACUl6Q07KeYw0XntarQ8
DE/hd2f6DbHHVlC+K5fxf6GBmGsRfK8mB1EwSmodBzZCvwn9PmIpgCzbsdtw
ozGMG1ycoDFgckOHtWTzyW54QQBbZ74ROls+m/NZF0oC05Iu8eweLhbW5WgM
dNkoM67Q/gemkvLIIMntik/ONfXFogzQtGr1nOGsdoFgXbi4VK5921386fz8
51xVNhantzDz2xJDU78YCfAVFzTF5KJRlWqpqE/iIqxlA2M61lw/o6xBdJfu
k//VLF4DvDH3NbTIs1IN6HL8lZUDXfpxP+Kez0whEm9MfVAJOKK4tJt0OmBI
iLvSlTjMQMnv+CuFP1+bDJci9cH8guIyYwFLWcAqsjhyM98NYpDvIqCxXKtP
d//dRpl0XFroRfBheuuCjA8eXVpCSOf0rV+X8r9HExRo46+w5oT8gwVxnw54
F2Js3Xn6dpfhBHfAIx8d9/G4oCXYIcY/DlgbGsn/6kqBzv6IBBVnlllOzMfo
mguLOX8LvtHw1lokinf049HDWahTqr/Ah9LF/8V9O2o3IYGq2EZ9b+9C9+A6
vLhQuf5s9NvDvyzD0kH5F9E/e3s91a0SvM54Zog4wJqbCMK8XE6+gfPtxr5F
U7Qy2YHoWOTw+J82cgSKlsfBELgRKJgyAwbwx9CE0w4U+O+zvGmtNhFt4aSN
Cat/31KXw9C1iTW7gMMX24T25B6SdKyckkzwwESiJ1xiGRT6nbTPMiTmH2G4
DA9s9JMy7d6fbdHFeRmfvSbtgcUjEdXLIe00ISMdZjbcvEhDKuxA7rcb14LO
EMjBS12rIVGodpjPh0B77RZkb//5XXnfD70WVROFXznqiNduT9sKOrIeZiEz
sxhN09TgGw2G25mtB7wGhsDeDI1crZhch44wwFZbz4O/pnYiPSePxUzWWriA
FOKnuFkK7TbYrhjgskGAUgldX7KhZvL5nJ5C0RvLCRnU7FOqaQR2v13OMAAd
EWwEapi2lnR6XENqng+nr7SzPDKrmN/u7DrFkZBETot1VaX10x+LCdKMFOyR
mj5S/NgW0buJGfnHDi0LghW7FeE4M2oLPmJJ/jV8E3FA99o1rzi/Zh/QV0Gt
LE0ABv8NkYD080EGLBF5ZPlB+bJ94FklFsYQhfqEbxxmF/dnNd/spF8/00Uh
6PLTUEx9tjG+WgQrYC7J2CocoUl7BIkV+6xxiJiS8qug+V+iHzkNys4LPsvr
YxfmRm02If2kpKmtZbkS6c4+LZpitZabNCJ0LDdFK5QAUZZtnfE9QUy2k8jh
7ccvcKF/89+LqEkRBoEcAlOPeL3efiSC4VgIPvPwUjwy5pvoiXevcPEz9R3h
zDrv/7gXr1Ud9Jrq319/I6pqlJWbCjX/NJb1lZmtdRLTrU3Gh5f+3uZboFli
CFxzdoi9r0TkQ9lmsA3N0mIvyV8Y+1CPd5rXQQpLMFpRjnvrAGRGqNKs7Y7T
FZZj73Na6yzbF79aGCSKt6iqaQYbQ14AGtyVKN/AWnqyncqAVLApKsPblM2V
o1Q37zFR9YEnqKuwijynInUkKhhuo8gC2dbRPlUVf8XGvX7xvii0+HUbNKn3
PS20v16HMPP2SGWBFhfdAtHeC6OAYiSJTGn1TSeO4DShgAPtkfG1eYXOkuQ4
n4SLguyUfjwnCpFZ/VkHQFEGU1xucA88tPI/4GuPpTag7JzEQ2TcMA0T4qzT
7Jv+LB8n2bD4R7mAjvfjWdpwKGt0DKoZXkwjvpsNS/BGouiu0zNhLkLSynmn
YXNsIh5l7jacpEum8YoClg7+k9vhNQqpfyDN37JL+59v/JWDRc/9cno3nUcm
bK2tn3hY7a0QMC16AVqrRTJC8VaY9YCutiXCPJ0RmUBvCAeWh8lBLw0yBKOz
VDYufSbEg+wR62pwGmTFZt72+CQch3YV94NrZGewjK2CsgH8E9JDA0ju8RJH
D+wkdtFa4jhBSXyAgWU4IV0yUS7GgCdrTfj/iem4yiPhlV7YhpseRxLx3Csq
2K0P8l41I53pRTStxgM3us5cVuxWb+FKjQodRG1bDIOqjm4MTlFq1f76C42C
9km/GMVGKCk94+XoT4u0kpJFPaIb3ZaDRX7hZYkI19YRAqn8Epwt2Z1gxF62
x7AEktgAJ+Vuzrvy0DmDJoE1WzGFC/XzppHV4SAOPSljZW+WuJlhp5fh5I0r
IFzdqHQiL4Q6rPGv8D4owiiO23Hqt/2MoY1deOoRTBX9Jiq1nTcq2/otYD0n
3O7c3Pev+ewxPfnsUUHuMKXC3BaPTL6IbTKx8pISM1yCTIAqzFhVvRis1Kuy
kVWhpwsSWeLoEWS/+vK474kigzORy1BM9xE/NTTyx84OMAMr5cK343LurGLj
6/EasrBGLwSN1cX/kIZso/kb77Ktml49eZpQ5aN2nB6loXinqg3PTWLV9uJP
pulS2/gHNekw2xfxl4fXWV4zViwiikl3Ix1MVI/s8JVRyBnOazZY5axNRxjy
2PHxoSiVNPoft/XvbmTtil3e2dn2zEpGPXcwvc0lZ65OiEaGxjW1DOgYZAol
xasF0d40VuuZaDBe24iqyS3NgpSvyOXSFnwXZwhycmSbzuoQ2pd3ZAaWMqLu
jYl2Z+RLYoGnzb5yqWqWfY1RrIgFPXHQuYkWFZTbhFVVixNKmQ5rBPf0PYlI
elzbNtPV661anfFfjzNopfCwhshCs1PIj5azAMrKb8uq28aXFC02fTorLTAy
tekDfpQlwE9+PKubl0Xv410mGl6Y3nSFW33VTMYbQ+lwIY1XZUM1P65X0rGL
9uiLZeICdYSW9pU83GxtnSFGqbeu6BSoPxUoPNZjOTSwFXaOfBL2MDQ3if7M
o+DCFNHQaCnAMjQhnh9oXgWn2M47sinE0ADy0ozsZ8Oh4sTLFB7ILXHRzzSc
yO85k+qtx4i/Nb7v9NcL5MgsXpEmYQRiq5kJCXvsIPE5yCiT/3fOL1sSWxaC
jZ65lDASG6YdxXaMhYaoRX8aRR0m2DYrkGksJ8+9tg8FnxCUdmYqeh6KeXaq
ttS6+4a4Y8InAYjwgx145Y3glO4AfDSvGse7v8uwR1g1JMl9AJOpVj1wHST/
M6Kofn4qdaO0sULkYWGvZHZ2mmW9SRSKUkrmUf3hwzHPzM7dDQhp606WVzjj
+yoMqwVS+AcjTWVii5Y1ollnTEx/wU1kPWXHAy4x5hcemJrbqY/0SLk0Qm8h
FQcdtqY12QZSsXfXe+mXrCo+IF1uZYR67xKCC9Ahz+KpLE/eT/oFnMVOLJvE
vUcyyRQM27uJ5SkavBB0bRzMnmXOk30EdYA/Z5BEQIBCNJVEcF9IOFpR7Kmb
MBbrkleJB2BNksOPSGmJGUaKgddtZt8RxkzHolKJHW/EareoYngWlZ+Hp1Ub
oTUIJ/IaU9uCuqYBMqvKi/nJS5hggO6CXOL2nlLWAwwE7TLTYWtKXv4HKgJv
MLzPbOyHHXzUMdj1NbDRXjmcLPzD9Z15ZiXeqF6ug9ogOVJI8nQ7wAzRaOpR
YnuwtQWORiOejY80UDj6QJut9l/c8CN1BnkIpQxWh/NCYtVuwRj7nbMGG0o3
2XHGN4hVmZTtTdqiMe03G1A+/oO8LR1YfBpz/G3JbjDxZZpqAO9SS6CIBpQM
in6WrAIwi3cmqiX6sFqK1aT48NuNGHT3x3zZBu3/omGw1v0WaiJOhK/zdLyt
ReVx5+2A9xSVEjATv/W3J+JY1M7fTaMWSMfG0qLVYQoJ1qgbDQ864d0IDKOv
PQQW8nS+cm7n/rduf58qahnchoGetkE4oMQcIFmFzEoWf7JMvVZvk2Yrilso
t7F3aNMEaCl9swFhae32EPhuBpSVDlK+Kd0xx9sylf/uTh0IPye/xAwQfRq+
u5g3K229vj/wxq+HkQqO6X1agtdGxx5X4ptUGGnTwvZEw8u6hWD0ZAOLcSa3
VNt66cpQgAI/4qd4EYACOfqgbogIXPobZIIdCuByxATk2zrTfG98lU7+RHQs
RLv8h6otjojb+pgkr7fvQcAMZwCkjg9J1jsnJ7iiT1Go+d3KPMuRPZ+i3FQO
Ec2Oc43d8mhelUYZBvJKcEUTNNEr0W7B5UL8N7drWLN1slYFkSDOa42A3SD3
/FNhKR/75Cm1lNQrX5oxXgOn1LaHZQSc3hiNZ04W0jPj6GIYZv1R26Nr6bYu
ObdH8mQr8z8Kx+PIF7zxE3YCmTXwWC7E4Y3QHftUNckWVsbeh8z1xmPyeSy0
tv4N6wgYa7cF61XqLTQzznaGP3ssm6+hdMI3C0qFoOjf6BCc+hsFcy7pLmDY
Zn31paL8Tk/uFuIuw4Wr16GHUcZ/QohweiFiG/EnhWSQOt/XGOc5HbeWx2aK
O3rsALFBFuwfvQLY2X/fYhjDJFmWn/boxMuj7zcPDVhZjw7Dorihi7+WQmkw
4UKpB1jMWOYVop1wPCV3vPI5tJoQGNMaAVvaVvTTi7UlhHnfERA1tF3biyg3
ajyKgqKZb1zbIsrsYWmcB4O9YQ7dqv3xM/M53CcEexdWD4B1o04G0+I4CJrh
dAk9P6qaVDej9aZ93KifV91uG7XTc6DYQeFzXg49HfswhWprVNO5IUoR1x6U
kXftoHQg27QrUtRdc+j37lNRm694wvFIj973vuIAD4bueSHcWDwx/kBzQwqV
zRo2QYZho5QYL8iGpMyiblOMJXm23TD6c3td0iLolabKuxGLHDjfotIMbF0D
3tnJMG2hNomjjMQS9M5Z5EodJwVc2oLXtvA3M1yFIIO8Jfu9bPM2r6AtlOAY
4WsCiI6Oa6PddeqvwVga2jx2RNALwm0BCdMzet3kB+15UbCJf2oJalU5PA5W
X1AVQI7IWq0bvVYbr0hdyAWYNUnvIOhrPyRsXI30RJS/cYUy78o23IrU3GEx
KnifdIj0oenz4HwdiD7RndzqYvOkeUoG7qkG2+KiSWxTKaMEjbuix1cbILyX
j8uItKHltcbb2j3/dobXsdakbOxDFSH68UVWhzH22Fkg46uZKhsCLWHocjLj
Bx2NTB64WYEj+DIivvZRhBJFHKmN8zYUXwa/FoTBoZ0txJ9osOd7RXYTqSCH
4q6IN2mLbMqDiHJb9tfLka9zBxebTpRqKpMEqYmoGJkysYrh+6Bx0mG7iTgk
PvdO0OPjrS8PkELJTyz84mgOuZLiPSGXLwYBRqnLE01Y3clDgIRvtmYIOwJd
iztzVkAfVTLB35r3JyAfxjxYY2WM+A4tyiR6/jfeGBlpmvMqVKuLwXbyKrT0
VO2AnHZySyaYzOF8STiiUIWKiF+oKx7KrZYfbFINw1qHWIDlGOm+VFLwVJIO
5KmVrvxsCMUeCOoZjdz2PjoMcYzY5C7mRqdaqj2ic0TyBYbSiQsA4txnyxBr
hpWNmN6MA99kvfDerRd0Jd54qh19koF2cRdJ+NP/v/VDmRARfIUZfEjgSg90
uytG+9pb+cehaIx0weQEUVxWNOUjmhLNwPHRSER1ATAW1gTDldfFHy5Sjl4c
mJ4R6fqvygSV3i+hOGj8yCec25/noojXTGhHn8V+oX5Dyf2PCHr9IW6H3Xb5
oER49C+spTsK2H8HGm/wYqt+z3Ot5is0YbugmU9NCvvC4HVPEn1pSvvZJxK4
NNaWqVVOtDCiLyZERGjycnfQJxRyIHPxa/kqU4J5LDTTBNA85KQjaKY5MFHy
hQhKq+ugzHr0NW1KkBqEvRBcEaJLqqAi0MT70k0kSE6KcObLtd9DOQ7VLpXh
XQOlSMUMi7tYx0CGq5edG8ex1XRQeQ+hXJ0LB9ivliAyMfJrJi5s0HqxTpOO
Es8gU1DOkBDhHivd/Y3bokVTzhrLGypR2Z0autKnXA1tYcalvMWkI3QF/Qgi
BEPVZ/JXcXs18s0tEZmYmRnFcrZfxdSIuG/AcyO5ku+hQvKecJEZy/IQj/ZV
b80emAhYvVJFamjHfAc5rQ7DMwNeKeNlCx02YOmOBIk5oYDgym4SbXXQcpCl
S3B+ErSkQf2pI4E4JK7FEEPL8R9y8GdPJtu4/Ti7gHaHat370iCq17rmhl6U
+Gxom6aYfB+ZoNSJ+z8pJR2zD5/6c2sla3VnLX+ueBfZXcqQk3aHS13lWYWn
oppCkLCpNOxHvj6EHs9KGNWthGDGGFxHpceFgnFxzZOxBIkE9u+26j2d/LVi
x01fPT4GvQF5PqlNs++74ABSnV0K9uOX+ZXvy0/cD/n2+GHA50W1dn/qWSjE
aJRs5D5K5eufcVJXSKW3bU8rKV8Im4jPohz9cNmE7M27W+ePPVdIT8qx2mEn
vBORoT3FBF4BHv9iNce7sFzzHtH/A6PjfLblEmOFbsG03QX7lCivvr4nojF6
g09p+8TuHdCcgTrZj5Ec7hCddFiBfOXWC5tmMLagrE198b2VFEA6clUaHXsk
nGMOOX1+NO7wLfxdBxKQQERwee6jfkw1ebE6Daii81PoCHpq/AGe9Yxu6oE8
pywV7SdOwW6AYCDo0sfTYwBvdgscF8NxUg3N1J6Ldgbtapb5hb2tCxyJQTT2
ZwaypWLtaAazgAHRlJ/ixZRvcZtuq6CJfncBRre6dw/GuEERrrgJjb938RRA
n14awVdTrC9fst5xcux1pG9P5cEqHD+2dCsWqlgidfgHAq8W/Cc4DRGqdTYQ
TLzvOMJAqnWaulV+d8imnD6xzd7dCr3nbig0yto7UC1Xeh2rDxLWYKLo1NSq
3YpcbBwYeEtTJTVxspl+NvPit93DxeiTcl0a2phONkU1vypaGEjITyCqC/lS
vt3Q1XZ89N/twRRUdUFNP0GEcsaB5/Pl4grkj5+oP9N4qjT2XL9CkBur5RDv
oMz1UaQCxFdchjQIuIPPhKf7nylwJrS/Doe0QT6iJYJP+wh+JVCnhCd/A2jj
0+qcReuUHYZOFae1QWWURawkkhN8KjPVlHs5OX1nt7nqFipsGC47ZMMU7FlP
+I0NpDv3bQJp0dby2luoQ5ZxqgX1xTWZs5QZi4xV6hT2fQN771Rpzwi3f7rP
pKaRI5JQ4ce+II3SvNmr2mKY+Ljwb1yPXUPsR2BnrhiYwKuQtwa6C1dcIcql
yaCvM7FCiV/eLEwotndoen1w2eP/vMyngPdKvUHAocq9XAydljjkwYaiY2gX
h5wyQvgAGOvEBUN07vWj74vY9glcdhgYFv3Tu8ZLWSPBWL/M30m1VSFZ6Ylk
Pb5Q/rMHaI9kbkIPaJsm/wXQ5mfi+8wwwMXkKo4Gv1IaCtJ9F1TvSTzuwM5q
ZTWtEftbY0pB7e79Zk/C+M5ulQ2FybH9G3zE1EpCwrTCmmjraxKHygF1rYSN
4yOlfkThOBqWHTPQ7S2Hvz5U/j/MH9r0wF+idmoDD7Kuk4QNd08zJYMWJoUR
Ys2HPjJqCC/NvYRWUkPY4i2KuqF5a7gxm2sONcR0thf7END8KE5fQAycWRn4
VOpPjF8O8NEEy77MKr2ogh/DtGuSBMC4hcYIvPv1K2y4yfDBJwkSM0sqTo8N
REO1nxP8jFnGsA3nfYQFaqSSI+PTaUznucG4dEnS+AHbQb1wBEulGLHFG97W
osYNqbtiAzWl54TIHu4yRg8PcjF5KprOX3+NkwevjfQT4jJxSinTGgLw/fHz
HcVDD+vVGa2UDtmSnGeVT7wv19TorC89UoIWCydY6Z9I0JdUXejcs3YbfsEx
9d8o+XEfG7jwz/JuXO2TKC7sFRciKMpMFvlHkMTASRADYscZ3AVolVmvB5jG
CkYXVq1qmNTDXRwTfBzo8I+gXvZkKWfMTLsmkHIfFEu7s2WBa/xd9KCEK7L3
BoXJ3rx1bIsx2vn0FCiVLkdoUW0jQxUD/StAXAcgDjebg1uvz2acxqlCz0HZ
HTXFjiBkS9bYZsARLyRAmOem5EVwx6dplr4+1amGh5jsbOOIDJfDRgFA/InM
f+9inDNd28DIo43OCXo9P0+KJg42NWzXSTBEbSuJPSatuc83xrleC66khUGe
R9IHMvpfEY72VXeuVl5W6IZxN1Cz0kE3TtIbFsVrlwZC79tq4Lg+uilZlPqc
2p1ktW0F11ZEbFsRQ/rQN1vohoeRXZavaN3l22sIVggjYmx2B+4m6DPV/KEd
ITwK8zEe1MZvm5zFqEeu2Wu8tZrVk2jMS+Dvr4ZDAeWJd8i71zZvU1zVbvYn
dU4vUSISyw6iQa4VJFEoFtiVUnVMnt45omtYL3duzDrUOZuhtuhhlVjKJVrc
O63s78uRDVsPRdgjvhEj2166qB01/8n8US9WK3nKg1vJ9DpRnQpUOy/k7k69
Ev79fAlYGm2yMKJOam7/OhfxERxcfT7wQ3giCRcniSbNiHs6LcbSoxyRqywr
sZSoZ9rCsmO2rbHkMJf4biBRD2NbeOf4o/m9v1lcY36+PdyGXERF/39wr4zx
T5Bm9FtMybWBDZepVpzEA5ppnLtLM8Z9q3bmiIF7jxFiFIosFcTvJTvtJHf3
8fDRrdYxea+ifixx7O7sKuavJgZQlp9AlOCosaNHvR5Uj9Mbidra/ySXVFYX
Kow4Cw6JXwa2+q2MELdgh6O2XqF9yEfygXVisuLMkp2hv7nrQrIXSRPPKcr4
rE19xq05nc5dAYgd/oquBPQ6Ov/tw5cQb4rcQqOzpNP9nE7yvzN3/Z7zDS7O
/hYqL3QfDcArFddycK0k45/kJqw8Qi9P0PI4dp3VCXoQ5mRT5v8TejPoEP+R
SlrP6J3N74Zm5FnN9mvAzDdGTmH/q5mw0291H7U4lmwwQddjLaAUQqWCDwnf
vjQ4631ehqBScrkKwPHwg1Ck4RqL/XRAqG6kyT+7cJI8guZW9x0MWtA2f1vf
phzAcRGaVPRg0vx/iEtwIAn6DPcvlsTQsNtKraVPhzK3+b7qmjXYq7z9nfb9
Y4jpc/H95NueNvQmjv1eNwELfJ78yJ5q0doB73sYgCBkRCnoJmwEqU4aLb2Q
l7KPgadnYDvCBHK6PrFzf8AOzfHAEPCU7xs5Sq5Qw1CF4n+2tcijTJQFPh+D
yuwZIytfjB4htcrAIYLp0HYs08IK8w0Oe6XdXtbccaSCEbeedSIEMrbjGnPS
m5jtPYImwITJ97beoN0SAU76iVGrcukdvzGbHhTgY7F5ra5G4FjEZ6nEyhDB
vCaqR4eGXA0cZLfh0kuiTpUj2TBR7h6fRMhc11xdwxOiVvaP/+MrII5zoZBz
CELta09SO3dBFC0nR/MGmQG7hdyusgObQCyRYdbYKpO7jpwfBqRbEMrBXDvm
hnoVYWNaxrQ7WmqdtpY37oki2qp5uCGoe5/YqLXX1uJhxorCZOLZ3GL9jWZh
ybsz9p8zlgK0PSTGNcKJnTVHyeXKFXG8/FyQ0dgmV3ehieDVzu/8zgi4qmwo
JLlyMjIYkua4Tt4CZfMNXNERt0d3lBNvYfSgY/xAjrxxnz7XyJ5Z6ihxbrkr
uYRMTXIQR1aH/U5dUguYHDdE7B8zBMdPoJ2By3De/wUlJ6uxk5RvRARPoqsV
uvSdTQwXGIP8ckaEV14hVq/NCIRufqS/mnLJOE86h/z4PIN8gOjoiHVbPYF+
axwMl3LaNdBu1XJMsXgLLet1XwHb7Slvp+rEjQ1GpGWkmugMxNoJO88GQSnB
aaDB3fuGL4qumoF2mZtkmuLNsbUDc4CP+BumrtSv+0EYCLOcA6aHyEvTDE9l
Dz8Sq9Jex5C95YNQrmaFUdka+7DZ7ZwslWy71VlNZ85gC5rqz2CqL67JkiN5
nqiDHPPFltAJQR2x8H3i0Ew2ye2BwjHbSL73IDDaa12rySqAvMVbBoAO+oc9
+UDhVlNMbdWj7l9pujPxBVbb/O8HIOxMqHdsnUmAFrjqyegGD/CUwRmtshS6
/w7CPl3t7Mvg9gR5Q7GduNPbHs5+gyU0k5VUzZy9o5wQ+3IXuWG7SxM8bH8K
CsmWWYeGXZOuXWUEbmznNKMBqW/sDdQ0job57RS5yn4Y3n1HNE61H4cCcG9R
56SY+sYX4NRE9+l5ge8EPIU2mbhVnGOg78nYL+9M0g3BbkZY/KFoUCKhXsTr
4HU5KKnJLdY//6SIjohi0skdumzzoenRUEcyfMexsMLile9T9iWp3j5rM7cK
XQqaQDz19T+sIcr2ua7uAhoIG2ao7478WhEmGhqJlsfpJdJBsacsobhdP/yD
Q2yJFxE74D0qZhCUQV4nP24xcvRcZNX4k8/6e0/ERlQt9KNCmucygEVnwNkg
QqcxHygSbz3YCMdcmO213cuEhBHNFThoB+5suwp8GCAkLBfSwjAiOjzyS0dC
2LDU9/DYcUaaTIw1KlZbLvuKollVkIuqoPN+pIb/lBodV2+Us8LPwm+cmG2y
4nxoOmYo+eddGcNSo6WZG+Jt2tyV/xbLkz+e2vh7ff/ys2v7jlOcx99H9eg3
y8E/7VBnxd1TqzKE2O4zDAk9fgi/Lz7Owfn5KXtPWCw+PkC4NItAF4Xxg3gq
BvV/f50ZvT5LqV757ePJpxhhu4xE2b2rZ9xv6vllRaDgpNkqYOOdNsKUY+J3
YparUT3jy1XGruO2DDph5cyXclCfmY30TS3Rj5fdER2DeCywQ9bvDFHoCA4b
gLdYkJBapgGQwzoFNErSvpnZeE8heNX5U982NsugJKnlSGA56sVxOYznVuaL
nu+lo+i1MjKyJJ8wj230W9fhU2dUBhc2aBb7aUCtPXZGs6MDUMLTxYpMi7vw
DXCavz+g6JtMH82TTCl+O88MPwQ+Rh+Et4dTdwvGl5xQsCEzGiA3yPiMoKCD
UvMzwzFFSOl/WiogYPYTuaq8sCvzxiRAtMpynXVscIhge4n6vvznIIB9gDzI
xkNR34bzBezDdyRtW7eqoy8Nr1GcIy/BXQIZajaKtkQI7isc/Ra+KW9qRV4C
0JVdyu9ZIdc1B2o8TLMWYGZxEJYNWIujL2ikTWJK2QtTUe3mVrbQV8nxXqkt
oToDOrjG/WFxwLa8p/PNB1tbDC1XGjey4ieYkCl39VegTxtH4Cqns7zelCYq
hRK8gCj567Ap4jJluD199UGaU2midFhaeCnOhBLeeR4tRbZv6UrmQng/KiC5
Sdfx45FVy3RBBEMMn6lKA9YAf7XVN67eVDwBjGcDd7ujv0dKui9IqcHleMK8
cYPf4U7ihp5tJ08HkBxfWSEOgCJPHK1Xtg/zBiztf2R3AIefSUs/ET7sJapr
0dtYtiO/alLoaGfQWPs54q99f2BOB9GUPd1WOWDiRS4Y988zhGbP29YP4Vvc
/XpHWwvjNF4Mnt7HslwKF+7fnkRcrzp8urNm85R35aR462nViI4G1AvBMdVy
aIuXUZNk6ffRDqiW2/yvm2FZ+pBnlDFEp/4RyYZ+ibQLl6pH+INgp4o3HMjy
/YP54Y226DxsYrAgWEs9WyAU6Nz6gHLvVmfAsQzQCnTJwAvn85U1xcAgiDGj
dD1WOS2YhAFAmIaFo8TmGAWgta2IRNOAO60Vil2Nk+oAiE+BYUOJJWd8IXl7
Rb9HqfEoz+HNFSuibX8I4WhG0/kfKA2ZrZXd7xJ4053OfvEgwEDAH4gsLbgY
bhj0Ti4cgyymmX5mgWaGbLfrtTf8wjvNnyxfN2u/f9nGsJjmj5U6gFaO8F3f
pMEg7ICSKAcMOp9kuIop3MgbcvauhrrLjW9cgzZ6pMuP/PvpFE6nArAYtBv+
DjDeL2tDDlZveog+TkF8svQcJQbePWo7Hcw1CyghSz4rbOP0Z0u2vx34lODl
l870Ln2tFHVyz8T26QO8e3dVttauh6agVgNIaRFbBGJqDTdINgudLiWOVAGN
uXvXMPdsr/9yJeOvSurBn/o5/KBehS4WHQS1qtE1gerRNUtStTXkFLzitZ1l
I0aLeTs50poalnSYFtrOTU3yp7KexALfXdF4J8KXfDW+dSDagYok2d2RTdtc
D1La/nHRlrThS1IhZesmX435vvV4kS3EwyopApa+4LwTbGqpmWusiVtHIu6F
IIR4fBLRA/8QN/pd70+QIisEKhZeErbesFBkk2C0nqdH/WKCG46no4BwX4lb
HKep4GoUhNeaCskykewXuZoo1WsKLQ7ij1WKnl20gl8EB94N+/A/MFR2Nd8z
EFAm1u2INgdeNYkxY995hz4Sljtrc/E8rbpGF8zyojkpP5iNPJH74uuUmCPt
DGaj4gMWs/Wv2DJdlMwGSU2UHpX/r2YfDuR3pyiyigPyWmx17SSAZaO4R+yu
a4dS2MNP4ljMg0YcSaj7+L9oJxpWHR0Q2zJgocIm31U51dHUj5J9cpzCuA28
SdSjGPtcUYnnTUVQ7ZYG+IF909fyi9wGQtzthyO70s+yL9Hd+I/6yYk6qfpx
LPliDdNKg6eP+bJCnL3+zwqu+X1brqIxOTW+yYY9Fr0sy3Mw24KXVails/Eo
HnZUx8ywSgN+a/tlp1ZXn4WVGrJD+RjhvmwkL/IjFeBhxqLZvjgrHXUdkqT4
j19y2mVmD4a+LobYzXDLAmnkeC4O94W0y7V+2IhdXkP3KQP+hhdWt+Nu956O
LS9eAcCh9iBT3k3qNEso+NPGWTB4nsy5ct0ZY1BeCeMT0OxmDR/76MRVnoQr
TKLNHhNK7euL8yrgjA3YRW/BAv9+t400y5C+kb2qL0PWA3Z9cTahSYpbWuVm
xxLanl/Irr8Lc7d9qEDD2FjCd3spP6m8F5cJ8XcqGpcL6iLn7ArVChBfWeg2
wgcnow7qA+zYYv1PYTHbk1Rc/D1dNfifNGYYSR0LeZGAyTUyZxNyGovMfSYK
mmMiB9m5W8/eobuIAtOOXMkNlOCSUUHaWQq4tvvG8QeUS2TjxPDy8CVudEvG
xhx19b3fPjuODvh3UxYDe6uLjGF421bVITcv1bU+1Pb1Y0u67PUCH4NUF0KM
Evfj5IhW27YhLTnj7MMBFwO6UZ0M4l/JCaOEd1bvDScTEo0S8FRvOVtM8uZ4
DRus8A9ytl6QGX2/BJ/A/b37pMnFm/lErq6Qb3yNSvpLwP4YHQTDK7skQtlJ
CJOcZhGROJYnddUeH0Z/YzmevYyfTO8prXDuiKos2eVnPJQlcBFXHUk5lOys
L566s307KuvvLaRAAx1GJnwUWTqKR97iUMJ160kzzYvZuXUxn3OXJlGwPj42
SDOVDJjB/sb1+Uk3bnTOrpvXRCinGbj3IG7z89hUFyRZs/j+8nK7k+OFfc5V
n54N9beY2bbe9WBmx1fnauui/ey38+JemH8mur576ObbsJG8YhcwIDWunIyB
an4DEcpYreBO2/y5UedZMtrUiQs79OeSPA5/jt+1wjYBhCcldSrOdXiJqXA5
9KXKSpk0HeVnyfXKjfycCy2JppPwXGx9fOJp96Z4oXRd4rrcfyH9Rn+vPj7b
cE7KxOQlNspZeY7OcSMBiNh7n0C4tYDw9jyUHcGCxqXf0CKkPWDTYc5q6nBW
8+pURq0FQyrLFr3cRiRZItQ0lh6k8BXTtiUEPoK10GyKR8k0UKV/jzE0qbXe
SJSQERKybg8MiI588uEhi94bB6FJwhVoc37MxfQml+xzcEIF965TL8HLJlGh
wEnd2VuD28b0upgsCR0VDTfYGFWVQcfVtZsf8Ub48iJIxydEHqu5eOnZY31y
2TlLfLSe4iyE4NzT539i2nqa7YHCPlIKegavsfNhyzLDN5WAsVfXfR9TNiLb
rApR4oXTr+fmHmq+DksuWCEHI7+1TC2/dUoMLDJchVjqEha6VqlQaw3pC9v0
9iQUPdlJWsdPPcdUEWaSoYMNSnkEgqPmR43Q/w7aINrj5aUoJFfmN+mLrFJ7
AR2x9PfZCsJYSH3Z3dldcswZwNkoXbKSSXUUEg+l9c/YgpjmDclitcqFXtSI
EO+NtrQ/4Gjb2xsIK2njeyEze91Tj83gesGMoPBwtNC9edI6kBLgWeCg6PrT
f2iWkPEU6be6zZjK/H9RyHwNCJeOY73DQd9dAIHOmVl4YmK4m+5SPYYrHbmh
3pO7jfiDG5wQObv3c2mXjzLjvEyGWIbe9acNzkKCS1R6p7IbqBoL459BS3cH
RKZiww2BkFXETlwFuHtWt2wP5SObeJpCaEWScRhR1lHhqRrDkt4zT5hRHGFJ
0DqNRnKXWl7a7diWUlIZ622rPaUU4R1DjT08VYOpQEv4zG4veWQ3NawBrRHX
dm1WdjdunYUuH76LDzbL922XOVzsCOd8pSWFWXD3cWcXce/ZPh5IMRk4m+Mo
lmXlGnHtVGmjaj8EYwfhlnTRLds3cmim4dlGmGLUcVxyVTzcH22Yy+Msh7Ep
ostjp5Rp2bxhc6t7DmxFAupOtklSyIOPEq9s0hzlz3aUjWvIB+YT+9voSeqa
mELH/viTP/dVf24RX1AWyhtIh7cmdQUXlzzw34TC9cE2sPzRlpAmqIfocDTA
SBSNSEX903Piv31BBsAwYAAUf814qIajHfTdRB9EdtyzMFxbUVnkw5qx752w
/JvDsQvCse0TwFLCwZZvzZEEDy395HexvRlztqDO/D71/IIK6mvlmE1NKeSd
9vefahnybInH6CvpJXX2OSDe8ccT40rVBJ8HWg5DijmxIEd+S2xzl/v8YQ5J
AQ8Fw9I1uaMfYPKSm7H4r1sFfUkwpiq6Dr2upWk1xV9w6MDMZwBJ4LNFfG5+
tEoMiquflhS1gt98EsmZ2PYTRCSfbx/yI5VE9rVkh2f6qcGHq7h2TcC/EAOS
vw7lNsaDsRDZRnIR62PIPovAXMZr2F7qOJ1jEH+GsOv4HYRHjSqsDFV2/pdH
Jevg2i++vl2EtYNrG0bgXj+0CAEGaNDjAARGMlX9yurcZW6fml101O1JRZvu
LE9kyQDZpuxNejbXt1LIxUSVP3ZQoN1ETyv37Vi9hzIgl+2D67LKxkTBRSbz
4+Jg+7v2i/wKx6HGXC0wRKPvRVwqUHzH6BVPVU8ukDvfFaFDV9ZqMB8l6sgb
Bnw6IOGuJf60pAWevq/4DMPYAe1ttc5xdFG0CUAr992tk+o79kR7k1Cj/Kvo
3rMzBpX25aEAaoc4mC095BH+4fTGBYSRIrgMZwFQHLZ5lVz88/4dUM0vvKyr
fTDS77VdDkYk/5GTbn31NMfE4SMcpZeBliOFa/2fCMKf4hC6pHtXanNwWkKH
TS6eFk982K5jFmKvvmHNZFInbFZNSTmLmlUz+fxVcXejYOBYJnEDqmiG9J6B
ti0qrwfZ/mPNirkAdxexLk4UHhdC0IvYks2a6f9RlxqYxIOWJOi3PB1EkNR8
uz7P3F+fXspaAoZb6hvhfdo9x0Je3OT16yEryocu+Ie+x4i0Fbi9Djry9M3K
WnPNix4pZcMY7PCZZi9NiOu78sX8a8y9QcffARy2ziLFp6ODmQ+JhERVWoQR
XPLSmgbO5z6qNii2l3ES4tql4zCrO69AvWBwBeeLDBEWUvoVCXOJNAINt7CE
zkgiO9/Mm8RxIrnn5dRtxcJvtrGtkKdtytvDzvwX0gsb+8j1WL6K2suH9UXi
skOGUS8yxhWftvSapYvumbI/KEbAmUESVdpvW4776NYIGzp010ZM/CIR6XLo
LzaehbXSRXO+482NH2VNoR+dXBi0VQEVCYF/MoOxqTT1g732ZROkrV1Q/aWG
URh5aV58AxSe8aLUVobO4VcOhNbi77F7uznpp8Tl/JyiBpmutL355yKKWdJb
NmSB3vMRJQWxv50Bu1lB86UqaMLNyyUejbBE22ULxO9xHEn6HB1FUmn0OXb4
r2zmAmvGtu9kot2Yjm4i6adUcxr1RZb9MkoQjZhSHqwztNlTi91aNoakA5qv
7ly9GWNd4O5HJfOoUJuRIgDdOTFVkoezb/ppuX82UJpL42kFHtRrk4axFM7r
kOmaRNH5UfkDRdDxX4t3fNgdMsm/Yzd6SSksBlIxpvaKW/xgKhNiZQLszwxg
JvGFt6Hc/nkFg8M2KwVVy9jKu6HNg1s7FY3CgIh0iL6f1epKDwnBQuaOZ4pA
ZacaAjERuubBJnpdSW0PI0DONoUg46W3A4tQVfQfVfHnicoKZD/S8pK4NPtI
mMqxRGZyZQyGAxKZPchQ+n7crEAepKxbwvJhLSrNrIoc3APvruHkJ2QWsdNk
cHB4bKg+SMwG/uFBXBmvnrEj1yuPoZsaaPh2KoKuYB0ku2nQVz7yzaLmkS0V
9k2/rbGwG6xx1m/vRFzpTe1joEinosX2fE6ZP5PzZfTDYJ5zYTJFJyLEjS4M
+Wdpf1cDeRvgr4BV0mTD/3fABb/aeRzgWlvV6PsJjFNO0sVPmYHRmemOzVIo
HvjmP8/gJn9A9WaW3iSpOUOZbQuwkwYsYqY7i/ZAy3iu7RRMNZJ4xvBBBUQj
cmKR6SfkxjPOuWRT7FzX+9XGO8wovScWG/abtEohPy1gDBleXRnJA9A+O4Fx
JbC0kKXDia4zvPmDad/Z2Y6LN4gLkoxCE2gpG7BDp90IFIR/BY1iN0MKDz6U
PwQP/vt7FBB3ZE5QTiuze3cyPvcQYfJiOwGwvwtL/T6E9IILoEARBejbEShP
Ec9xQL1ek+MdLN7J2KkL3N8vEf0pp1wZ7Uwx491U8Ix2LfHZ2oTR0RmTXRlQ
UbDo/2oeEfCtfF1lfTjNvuoUa5hpL+C+rgAuZ7wGOnmad6ZzFSlt7jMjBmCW
Mn1YUMqyN0ZxcPfhohfh4TnGtUl61bLnulIeOGSXfYokpujFYAGIvbZf9TKj
Gr0l1DzmCv1uexKibUsdshh8Z4EzoFtYURTGJ0/dicJMMjF1W8t/u1bXY3vE
FbVOZNgdEqmUoNE9q2/y2JHtcTTWMSRcwHYf/cd5iplPG3JoJw/abAGAUQkr
Q3EkCnOIkulflgsgtzH65XsWk+F14fRSxvKpKtoKYslF59sk7WnLIVflLJEX
j1gL5SYpVAkR++s5rm3TW7eGVJBB175euNR8imBjZ2AB55JbezgyOVJO7bEf
ze0yMsc6cEdoN9PZ0nyde6MHbPdbZCAdrfuDyDvjnrWBsx5bLzHVUy5Vkdhm
kyhFXKtia5dmSKxHrI2QNDGP+sEd3EBTCCH3JU3LNg7hOrKm7Go9KOp3VArZ
qHo8IcwDmkK58zEBOfDx+NDtuqiCDnelhnjQwRAfTrjzndkiF1maZXDYPnF3
ulDDa3R13qrk0/U8Ky4RZYKGhWV6WrGWeKIta1kdd3f7QWtIanGepaUxgBjR
Dr7Yk5I0UyoJHlJoYEGg+IgKnp2loXv+B2svO9t8tTeEmfdhPi+rALn9uE/i
ihilKaQt7jwLzVFwgpeq7nRWm+YOa0ix+3jmDfuEnpxkZqCM16zz+MBv0XCX
2gK/DmGd1lLFRmjH5AzuID5LEo2Rr8hyjTYDsil73GBYHW5Y8x2KJ407Uiix
La6XA4O0UpMdrRHXa7WLmVQW2wZJYU78pWJddqDcTMFGGssNKluGhaau3UPd
JaTV9cnVWfLg+kbryFEqa4RpemKcum1MD3JsX2k9NGynoHxsXaI5k8qUe5IZ
AC1EVsWdSdZlbvxybpdnhYBzB+qR3+dhmDfFbhwSmJGuC3QWvYVniz2FkCzk
GRuVXymobDQBG7dBSGTFFxVAfnd3Gii1BG3u6fKFO+V9jyP9oz6ipzygkC9k
rgh+i/jgg9w9Yo/ukdl2fiUQHMBoBsWv+DZteArarQ8zm55RtCSxvgtkdGIL
CJjFHSq9DsrrKZ+5T/RVs+QVq91rE32MNXAKakfOiMpaKqFsGg5m9k/9OBrq
wCW4GGOg6l+ZlnLyN2l4BBvtLoFji05KrX92scfSXo2PmMELbdkWDMGWDF25
Rs8S8Kx5AALGA0UtmCMdi5B8QLbJvG12sU2oR5PUy6hdnAWVDMJMF0CSKjh5
8jHYraguMEsfRc1gg2ZCYp+2HNlqOvPXML7IX+9LZ8RNtTwhLMUaIjRA36mB
ZvQA4Vu5W8ECThy75HPDzdzh6UYFnQ3jLtdkd4fSfExKsbrsAM3eVXS2Esi8
6kYO1oUpykgs72VxeKrFmi8F55mTKxv4UqKgtj81gkrOsvwJ/bAJYgvqxVfJ
jqGrcC1Pjd9kGoF5DcOvGNvZF/kDTIDZrjLzdQJdPdRiH4cHYq9JqCScB+3I
sxEvKMeLea0iq6ZQQ+FIr+hkHwFeQSJcQOM55dLl6RbrVxxk55KSN42Rii86
ZzlOWusPsuKvmYhK7VUwZdLl0Z6HMjonkaFV0sGtfWIH/q4JIDEeUospx7og
NRdCzWZxlk+bGB6r7ggOpnrSHGDMtJ0yeXUK+GuNGiWTpRFWm4gIXNvqmXwR
Z1u8OAITpLlQQtv4VEKwPO92kxv7sV3eE0rFLJChwovFdtBgUO6iCNr8fMvY
ysxZouwiZ1I4X1guzSr1o5fvBx/5z1+e5Zm0K+/j+FwjGGxJJuaTEAtWPXpc
ESdOFdvj839IQ3whtJd/8ntWFmlEVUB9VpSLryZvVzgTMYfBoaIAN6MaqjVr
KUrAnO9pkayyu/Q26oZTk2v7ivVlqZU8H6tzgbxZeyvjLyI+mAwnr0eYCy4I
T+5OuJRPyDfWmuYWN9d/FtMv/FaiVqkmxLOFv7TfdDQjLRhAMkFy2sC8va6Z
SatS43aOFqsAQSMTPkQwUIPGw8vlf96PxfssTwuZNpLikV8KRo1GzMCq2h93
842f4Zye02+iZvsBiU3bnJnlMJ1i+IO4WIV59yR+74sku9jmkUwTrh9NLdqi
kEAtJ+CaRFqvbbhuS5iVE5ftTLqg1NjsUiN+FqaF9s92q0rJVqPHIWtktCAk
XjWKDc1Yr27Sv2ERMo7aq7BO/0LMzsvB/mYS8UkPv/PN/iC5URmed71l/t99
dkA9aQcB3g2z0qnwAqfMjlcuj2sp98v9kdGsYnE0VuQz6Oj7r6Gg1EH1n3bJ
jaORhAQrJa3eCmXk2gvpyWptmRrP9moKskIC79FgRAIF+jjEVAK8qk+uL32S
qvlSMoxeK7e7bJ7Vxngw8GqI1HwH1+DgBk2v01+t4zmmHpFQRVHrqQyX1E/1
U9Ll/ARjOOj29vMtWnTlvFoZB7A1p8GGz+9gpO9sCPlwZIaNddXOapCbfkfE
ADZVG8kG6wJCq7WxTgNeKq+vk70NtrR+or+PQaCVoW57JBkyGsrZTcFCqQAP
FIqYUlirLPOXM05mW67lIe4s7P9Vj9qNKDiREhmm4K+l2MMGbTEahGahXwQz
6qarR3TWsGGYEfM5e1Dprs+oocef1Ip8fUdhbyR6spZ1+aaIY5Xjtu5h5zSb
jOZdRujFiG6WZL6vExamly7aI3BpoWu9PanoLh/IMQN8ozL74fu2SLR8YMct
CdK7DqPZpguomVqXC3veXabEufRaEdd+8ONBOKg8eTxFSTdFzGRRKHB/TKtR
jdjOJQcqEDo727rsLebNS/0Pmns0jW61V+9donrMa8j2kOe/YDsLT0W0fMrW
hEjhGaHPihlo7GCIoiti6DtOyLt37VxR10fVPSckr8YJhH6nxNPyQ4VRIoam
xhuJ/F8ZJGFPXTcqAnRFyYRMtarWtjhwK+eft3cHm+x+2BnIzWgF2kBlSho1
AoygwotHsBRFeV99JAcButq6ValTxaHG83Tia8Z8ZeGkLDfthNhThO7tf2+z
2dFdBGGSmlFtEINSy28wlPEVZpVCozM98IZIV4GpmCrKG/92moBp1gLLkXhF
gCuCA+f0zN4vRKR4yo5eNoIakzESMeIYhITmrAzZILWBYW/Kp5JBW09+d0Vo
8jxJOM+lf5JvFS63m7pMjx3+u6rohnztnyvO5k+wVe9YiYB3ysokzAENQoww
g4YiFvaD+3V2teN42nopzWI94oHq9aGZ1ey+MGYhZkngGOqQNb511HWOSBHX
yInfq3t8G2WGYLyz1DOBKeLar4ug3BgixVNutMJOQyBvdLvSgKUyDxd5g+Hq
cNzJH7Ia0AM1orBy50s64589FLCmFbyYFkBNvr3HS/jU6m9pOdb9QdyvCUYn
txYzD0HmmB0KvCkzaK5oe1GbHjorBI1mV9irCcp/GQI0ZR7YzPVBICp4Sr9v
aCO+fglqiTXR2WPwU4QgjoDvLoKsqZ8qmX+4VJZcX4eaOao4qRyb95mxEQ0t
t++N75dElFHoZQtiMjQlKPYhX2sPVPTigg9u4W3nnLatoxMSEz/NfjRevwwU
cCViOswph0/pyIoIbSYd429djDTgvp1M3H4lr25/rnQ4TMg5sFGHlbcNW6J5
U1KCehtPisAapQH4A21zrXr29WNx8oD9RDRv4j+dkE9qa84DIT5q3KXcLp6+
jUZv5mIvZpiHEe7t6wkonGwGg24zwYcIbu6BVbGAr9T0UDVdlfAM2DR0zYnx
SFYsrn6X7AHwWo0yw3rJ0RtXNd9tgVJ6OdlrsVJvFo6dirF/+PsV84r/uxEP
eQR9MXIvX4ZriJ1bdNuOd9Zwkw+xvkWIAYFXV0wg9VPGpTYdKzLql9blPyWo
jIeCHKc5Zep6cyz4XLAB6GSsLo+WA+VrWXrqUlw3wgbekCOTQvWd3cahdrLS
JTWe1rM1LinBfQOSKhoJLCD6f/beIFosIxwNvp/5qA3/aa6CEhHlptY601t8
I4uzpmQkrkK2bTNfvedljjEGC3SIfe/HNZqY3M2SI9+l7FtIUGb4atHXrRrf
qASDppAQptDDtUK9dKHDfs7IsY5xzeCscyMJklZ+lTR6nNevQUrZ38cuvsI+
Pnur61QXpVVvkG7Mb3q45kxJoawib/BhovcZiIiZpdapbRGtqV09weOV0ORo
SlloMOktQb7alkpk91DffO3qiHWXULMTzju7dTaAev4cyOw9VgvaNNFKMYtE
pDsGxAASsywE2zl6cvVV1J4Y61PSN4EgC6mqdQKKJ11g42NSc+jJ4Ib/Eaza
XuAVA5evlUzfQHc64dlBBetsuU1umIJD5odHKMrX8WTkLG1QpcJQE16Nl00w
L54Jzw3O+CUx5Vr1+t+z0+7rP9rzHEvueMLAf4zoX9XL7LqvC/TiGDUkaqFl
/f3PtKjdEg3apsU7ICJxJVZKQYn2SR/lCVqegvQB4zVM24rAeBP/Cprriv27
2lWzMxQ9lC/aSFGpJmztX8W4YicuW6hHZJB0g73Kwt1YOvyMMneiVXErOnqL
1F4xUAmqT4ZfK6rmpyE8Wwr9NephWCm0kgfbqJHh1z5iNiXbmPef0DeS7o+C
grTq+HVMuMCmuIJbiJIK1Kt00oscTOMsER0Dn9cU+7wsChq+QrIP7tCHOmen
qqDUmysfWr2AR69jrBt9Abutx73At3q/idUAL/S6/scQE4SNizkoBSzg9Doh
W1VwkfUvv4+bsnPBCBD7QH50Xua+JQkljmQJ/MOwHMB/Nnrwqb1d+JdOFiKD
VVKoOSC3Wx7OBLO9CfZwb+/xPpdFCCpURSPI2k+FLpRsUBqLMi2DwzDgT1SA
lqr9QIUl1Kqw97Q5UutVfsWmU830VA18qt6khRHE64JJjwkEQ6cLQuVvurOP
mhPQpyH91STBYsnl8sPOpUQCxFoIArv7wiuBuDWDu8tit21dd616BEc7loDm
jKCL4CCu0YYnEbOfe001cWFnZvjdvkAJaPv2HUrc3rnafcJZrMIiByQDWJg9
I5rxMhMrF6Ne9+hgMjOgxmG4eHo2UXg3bdraA1lLzz1jPV8Us2BlqYowA0Bm
AeU4oJd/gPLlu8kqSeI7fEFemZFRvAzcB3bbd6+vllpcsEbaNjChcydcT5rC
J8NGppfLLRqx47vZWXnn2aRSlN7taLKk2sjzBOcddrqBduv4dThVsM1MuW7N
ly1Nzbe2dxI6mH8gDVkAaYl6wpYSqEPgYAMkE1XBFGlBfFdCQYxIMZQdVN5T
bHSNB4Y9R3BCPZ2s+KWiN4L81XXwmq2oZVcAvSqKV0Goo0nsz++RZOg0xYZs
tFWh7OyqxWWvpWkVLV/H1ymWFaqLGp1rD+BFtLAnt7q5LfczJTV+2X1Yn5/W
N2Abo0IHcmrkpH4aWtet3roug16pLL+hBKP4N4QpBKvQZ9KwyjDeA+QuTUbJ
b/TFv5d2s53cZjryfpooC+rhbyEVhwTTob51MLmN/LXr8iABSJ/SIK2sch2e
8hRVULf3jA80E/dTQ9xcrQYwXT2yI7dnGr8HcNnnLC06834vTmZOraAKhP+M
Ms0PgXqcrntuV8GTqGkID1DH1okhTWi6kEqPKpuY3AIkB6qc8brW0R6iDojz
f9cfuVSMqGyVIdGmeYVcg705Lz6kip5RBUk2a5LDsSQ1wDNNH/yEtVGK6+bD
wLDQ11nNBjgoN7AlJ1s117b2b+3uUNZ9ZKIxxXI3lfZvZdS13m1GQRpGgEzz
zw1RXsvKBJwtFL2nmWZpokTIpVhrraWUTNgaeuzOFboA+G9VnCSWMnJNQ6HD
92gNQ27r0rWQAKPk3XHC9FsPaw9mGxeEOeJi5BlWZKdtBicPOX/jWF/7Giem
uVA2vfA0YMuKMQvwzl6R0AlXG/2W037IJK16MIfeGfnHhLryZ1/W3n6Sqj3T
4J8zNOA7eeNB7hJ3scVaDrTzYhQaq9rGzXGBjOk7lhlsXwgy4OyNc0hUddxA
qD8bKMClorRnN7WwkJ31RXEauua2ii3/VzOH8Rwy2BOE9cDSEUgrPamHg+yM
A2tPgJKzBzKXTQRxFKHeOJ/UjbAWApyciOkGVYZSwfXfeejb+FTJEQ6mNSL3
PoBz44wybcAA083N/DAJJcJXgbnYbdKo9sumigmEASVC9ZvHkDm04xTNilIV
ZBYaaLPLJ+iwJfigfVYRm45GNc6JE9V5IqpcXB9la545eIJH1703pocVJWas
Hx6s+61AUIccTzfO0UUhnPMYPxwzCLzzL0R68Sygu66CWfrvb5tz306KCGoW
2p+JJYb9eu4S08sAJhy7j2VcUX7fTicA4aZttZkLCmithoFHFa9ZMyFmdEZX
6omkLcZoiqrHFH7R7g74GOxRQWKCq5qIb6If8LiTBmrdiZLV1a9QZwIZXgSq
Qm5EUU7AAKl+4U8DDeqWc38W+XV7Kyr0wUcXQY0Xea41O6SewhklaRZFL0l4
Ik8+FFfJLHx0BNn04p7qb0mJj6tbm7rOjpXe9CjnIMzsHrFhCWz6G+rr08To
Kk4pHqvrvqbOBvJ50MeQ8eG06MgU9OVnWSDFV4N3ZkX76oxy+b3qNBFKEq4K
hkCsUgNn4WtvdNu5HdhNRa/JjRqydJFaJQx9pEcspSSeKJzjr7jnm6g+tcNK
x2KYgIO4ywckdUA46gNeBlsNNWfJkz+r02ONBwmcC96O6MbfYzjnn2yk7c9I
eZLg8VDoeyepvcXiSwn1rlHiwr8jWD6hwrBWZF5zvr1Gq7POXWTf5An9RnUy
eKui5qh1IAhnWqPnqqB+7VbslVNVKRBkWfXhXCicPxjB7H7PrOCvC9DrGRkA
zjRx8fI7wffBAqbS3DoI2SHNwsKeWRNN2vCTD55jhXUKUXrVm/whHYnvzPjo
7/Hb5yKn8R5HN0lkyletBlcYun1ZFUyXN2KmUU/yFackwPNxCKfaqLEYAblk
G6MsByzHBSH5ieQ/xneUoUEkXbJUxPA9j3t7fwe6NeaoOCzIbysvI61UPopp
vb4DW2EOgfW4lL+ZtB9kT+lRAbCxfT8s0yOpcYz5+OSS7lxDemJnpmEEgy9v
+jltotS7TKkfIhUgLU6O1Pt9SuKap/1Wn0jD/2bRauwOSbta1Guy7O5HjdY1
KdXKEey+6KExjlsCB7my3CjVfPSNVAEEndH962WifGYEeTsgpLj+ZumlIcVf
WLd6+4SgNpqxxNFFqIbWIyK5CJSQBnqoQ12uxqlMIXcecxgGe92m4k4HsJm9
FXY3r3+JGoN1aLreu2xo2pR3DLime4BGDUBUrtdn/yaV56EJLkmLEWV/DV6E
UIly1jj9h9RMeslmkWgYX/b6UlayHOXDEYqH/rUsnOOdLiXIKcGVZPhB8/RP
xnw+Qbs0u0G5JERnDr5XR/tpGMuRPvbNLtm810G4YsoFpUZ03kwF/zB5m96t
r+FKV7Zik1zbMd9ztNQWrYIFYi3nsc0QKCdTxNKp3kwPw1uIiyYaGF2yl+c2
di7owKmqZ7BVexDxI9Ub8kVbNycjfuZ8IchZKgZ53YDwT5q4mHTCHGNCYNDI
+LTArrw+tJkSU6O0Qq1ZEr+1ELE4EexUXzynP5nn/0lS5d/Dw9tg1yFUZ6zq
zh/kP4L6qVZSHmVyZh3/E4YlpQuVzqI5Z7AI8VBKiFnk78arR7qRlGBJahv3
VgSGQqwu6wxoj8uiHM2n101o0P7ur8yMPokRfyckChctIKYm/T7ZDIl/dH8k
3cIIU5dHTKwjAzu/mRo5rtLvDCAz2YQbeWziDHVywyrf42qrGP2+dL1Nh58v
n59gSUA2Qk7xPfs6s0g00fYqJI8xm7OHL+P0Ml3WT+mVJLBtKZHm9LUxTawA
lk3C5E2E78UD/y4chV5+cg6hHyIPBZefLw+HNAZqpYjdQY/rG1h6lm5yn4V+
d1pMywEKdcignmaQGZ+2Fc3+AE2CNq2P7/QGQ830T8zK+5gs8ghIMs2efOOr
hucc/Ep3RINXUrjqzkh1450VQynR31s+iM7G+zgx9ycOXtuWN0Zn243UazNn
YH0IJEhb8Ffy9MOVinEAYPO+C6l+SczhpupzJq4uXLY089+RTYToN4x6T8Rh
af/H1sgDS4dADCE6gyj10QvuiOZXojF/kKcMwHJ9JDdY7zBXxwIUAMJixd5d
urVfk9jvmTGq7e/HD3hExy970JJcEhXqAGDlBRdgdQSrQIMSplFMp5ab1o9I
KBvtjvXKyHIn3WJVQ5tVdnPk+6AW765Rnm1sUw1ZddVz4I/SvNNHq3dfpjra
phWhtC8X0OZlNPkBkHr1KTqdMzSZDiITU1GxpibDaOtGOHikd8QYn0jHsQHP
5tMuSqCf/QEuZYDdrOFBFRl/ZEkDq7CyrWfjvmhYoQc+azwJ/TtamPTaJ44i
HGHhFgf+RIC6QBPgFim+RLybPJxyswvxegEgS+Z8BObBhiZnCUNfsLSWW2U+
+ces1ijjmycjiRrxlh3nlWFykjmfoG31+cypQsWta/zCAJ3a4kpB4stl79Zf
OQ7W1JHl4QfT7abaIPYCeDn9Dz0c35Y3MjAKitPKRzsysBAORG/9LuSbqFT9
6MK2G2FV+McRAa+6AMUTg8JemRSvKASMmt//0Bskd2g17iYZLdXP/2maBWO7
jQIQDaaKQmqy3oqsfNQdjf7VyKYrjOJwW1IsNxiffkB+jDk5d2iXbMQx73q7
xLU8HFR+Q8YhNtsmWKsuveUzx2Vqmblj+gZDiAYIbsHCj+198dra2Cc8UhZL
h/XToFSNwEGeCA2NLib4N1SY5OekUHCiGSrxCiSuFzSWZHKlJ+bTWBHSAZdW
lyyFf5F2vFp5mplsfoMGbK0639OSnRWJi85+/ZSdjrnu5UQJduB//WzM4Yga
mNQ+eEFgTDy6YwifQMecMfeQ5ItJuxhL0bdMwe+ImmVVwoXVGf2dW8orzMBG
vGCieddOc/z9yC7lUbBdP6gvReLZdQZESMQiOanzrIo+VDsF5mPa02dtRuSH
Bj9kAYLw5q7dC6WJboaL/eC9J4BBwGb/9Og4YJK6B1+ZwJAwFVTGNmCWA8zH
C0vFZz68QwMELaZ3xagLLYzjEiPixGWcpaSeQAQ4mH5noa6nnYygRqhDe55G
BWpGgl02H3fOgOrSvUFvFovlnPveksEU2xdbWJaqD9RQC6qK5D5/QuXehanJ
VM4YYo7L9XQqqldwTAwHobwIhDkgaz6r0n0N/tMau7kjcZbY1V3ANlSHnZ26
vzjmf+Zc7zQP4obXSlvJ25wjJzW8WJYtksP07rrhyF/zccqAhpYmxm3XFLlk
Dyo81eJQbyoXUC/A5wjh/YC9RFptLiJVp6TFTTPdeMOfxwI+amp03bwC8H/0
GShroLVjsdkmow3cHkM1nP27bJYrX9rrC6Seia1vWzVWeEQhW8E/uQI5pYfq
ETC3NVqH5dMKVvmPoebiXLxQQxPl2t787DvAuIkE1mhnPejILkKSm48qGHvh
hsmUI2lcWTRevvos7r2vqYONnNJkt2dxaF70dP5J94lLdc/ZBYFIaO60JIB5
VB43eiPqG0e3spH+NwBXQzuYs2AIT4cO3Cko15ciC+r7r4/n4VQNYmKO1J2A
nECW07aSiB/fQXQ4oWHyvo9VqpToxN5qukwFsmLK3zbluY8S1QPUniB1MXFu
yR2SFyWz9BObRlRtuwT/f3oiRfywr0OMqbkW+Te5oV2aOqI9qYK87iHCwHQC
escLgYR6yPTUKcssGpHBPcwlMz2Vcr43P45N8AZC4wWqzBEZ7wizASTImfid
ruWifAFJjmxYiA8hnXl3V1IhpgWWPoM3JnQBeV2yFvm2jgwghULDPclr2+3p
Nc8ZnIM8Zl6Msyui8hKyCMd9QVc6s53Is3VcH0zbqI3GeVU2lFJwlmt5Q8zo
8BCMI9GEJaJUCAGq2EqaTjhGw249OrVnQPcAaKA0AxgPBtt27ZBctHLqnSPf
a7CvDhzgmhD3eYZrZJr/nEx2rup3ev5AfL8D6Bdyv19Fis5c36uOudbnlOun
zZYGDApp8MYoMd69M7bACZxQujy/YEWgvVsSPOkjPGQb7ShtbUWa3+8b3cxG
tXwdcNMlLVNSUI+a3ijfUhXLMJM0F3kRlxEy3Ka+E7+De7TRpeVcFvoWp/FM
v1WcY0qZ1xm5bQVHwjwmM0EAw2yC8AGA29zB8/hUkRikHRQnHcI2sGOxVe5p
ytxgaowe0uuqqdeUIkcy1H5/eb4wpVclYx8kAQOwBzVYLUrbgNlFrd9exavn
VZoj7MyzrhSTVMUgfsnuZJL4flY5/aL/j/AgY/VXWnBnfousGvMQSKlLhVf2
KB1b1OSV6Gl0FtsOi1yzi7ya0pCVVHZYv6HYC4m0uh69yR9B3iwqLWUWagYF
0RDgj1FxV3ORnExmbEerWpjah4HqJJOaRiWrREHf6R799LNsyHeSFQ/mO4JD
2L4LIPRMjBRu7lzYF1YQaUUqyXgPkNecVnmTB6uKz8/dpr3sTlls+8SkXa9N
F9Pt2ziraaYoWdk8bpSFlPm2wXke9E6BN/R3eDJCjs4SbpWhL52DRvmaWyIh
BDKsq+MmxK1WbhGAr8DdsP1Qh3m9v42hObkQq2WXQ1XwTza1t3gcPZbkPzZV
9z2Fk70DZNWNWa72R7MKgCRI0v+9zBl1myoJ8W10v+P/3l0n2ccjIAmWrXAg
VjI8VB5Bwapc1O6rzLIouOwUgoWXLNyhb/l6HM0D8l1ihXwwoa8If7ULh/qe
VsdPutbz+pYch0QB1jv42FomaBuN2UqJ9L8leprDRpdRNCMmbdF48+yb6tkM
2sH8A2i8CiIK/TKTxTjXxi29xXrlKgyILglIGTOPxEA2YTv9ReRLzcOJ5gjZ
u+KLQw0MQInAcEgR7PuQ6UN0tFifcNhHujoX+8Q92fnBfh6lJ/2GWdDPzpjo
1xGRkVazFaj/IwykNi3rZl/dIhQKW8+dRjghd+4P9/WeFylmekH0Wjgo1m70
E97fwV4XJ7N1Ft52pBE/+JqBXcBPQTQu8xOzbIiUKTGkcxDwI30C2FPqBBDx
x102rnw3IOCLVGmBrIeDvRUaJ1IRfYBin3TPPGtr4Ej21tpPAxcDunI1DcXL
geuRp0phDkcmXg9kz2Xs4PQtT+TudPSY0WuFwskfCZn4aQBmVOyfBf5+q4Vp
l5a6N0bniJ2earFuA8B7XxHtnH1P0g5HhPrCVkWwPp/Ct4CBN6Nqw0achkGf
EXHjb3yHSYq0UTC0saLlIGN2mBNBgQQasLH9idD+7zEnrJ1A/1592YbDxwKg
5vGxstEU1UNL7bGXljd4lAogpSSJx7Sy80JxZgQznV+wOhXHEz0XlXMn4/2N
doPWeb28YZG7kptgVT98sgob+qlYE/CTtEplvJmqAq4DFsmyubJFZPVd+lp+
byPj3gK7EOP4GwkU9/qA1fqXGQF6lcSzJZbHHaQixT7NhCuuBb+6KWzFjjl5
Ur6XlstATpMQWQW59FdsThJukbegBdsW5bIGyyNpy24jkD9AWCGd77mDSvKm
n4AZU1O61/IE3iheleFmhKR4meSNGnYALlZd0UGi608wL6CkoHRgoE/DB8Bn
AsKS3KpTEMznfbAmTglsyALigzbP8q4mrR+MpdV6bWPw5Xu2Qg95mELybjai
2BC5BUZW5H83PRTtJZL83l6UEC9o24lPHTz97QZf1p5KPWeQt+UVvhEHt+r7
9y0DBEcIy1auxLiDvF4ThWpf10jrL2fyoxbFY+VSFiM+6+pRfUDMvUjt2k6K
04ychVMWMWEj3BvxcIYveDbPMVo+10xKskGtWKQh1cCY0aR6hD2DF6Z6MQ/W
4fl0eJOF8FlDqdugHRMMdWI9eDG+yUNjuWcNKO2LV/OhBU+it1zsfAqKS5eu
QDbSSrbuI5JHtwzj8o7Soz1PpNVdTLpip0OI14pMWHsl2wPsKl3t2h8G/lKX
m4KS2vCBCJkaorWZVbWU8jaB0QSj8rhZNSHD/B78Vyss9rJgytzOwIHV+Ydf
rOcfbdGtCkyLCs8yAH0/4quE9wwngC6A7kFSwC1Nlim27C0J4Kkth/01jPqD
iVUcFuvvKOADWl4cGpBBDaxeBjHGaHVnlwZ6ETz4v7cAUonCNi9Rmw19EpO7
D6UmRHDLMOv3UIZ7YjvV8Ts3j1LPTHwpckNhPoriFi0TUAyl3VHzfhr/t7z7
TQVm2JgnSsgv+wV+MuznZe7mJPx9SK7uwzERz/ciDRrgGrLXoh1HaGXmOwzz
oWZpZiXoE0r0LAD7ZkKBnfhOGcGS1tWeEDI/pwrt/IitDLWhgRO5ImqcHpvs
LkGjdDdOsMv5HVw+kGgGN6pM7li/48kwPxrF48NcoRp1CchQCwL5JWjOX44H
LSj788hNrK3S8ZyVWlD1euGhJrr7OAo8vUKnayR+8qHAHUr5cTZqdLYr1I7L
7QpL7/8mUcHztPKsiiEmdsw7Cxe37Pjlomr9D+c/nX+Pi3cpAGVOssCnbJtS
lpr7dQz7cK9TMr6kD0rSScemMQfpnArz4TTfGPqtTFfpPcg4MPzIUfnDDWg9
68bcfgwnQep9h9pGBTwVFKLinBRzx6x7/jwJTtn+Z4NDbhgdWwqQ0Fts9eZ6
SARaqtiaLzGzvOYdQiUZ7kDePPxLlXJq/z+27GWD04y+2nBTimRSB8FeSXXl
YafjRPASvCWMxTW34McyX6LzzX+RLKeI9aRaMiWaxTcnbU7EbsYcDn/Og/P1
xr9Jgz9KMwtH0Z2Sc17bxUePNeF0mPJnVAHOASQOHaJHkZ4tQ/pvtdrpispq
V4qUkOUY7qyWX3ryWUhCBYeDM0end3JbcDopmYxHES2W9uAktbHeLl1tF0H6
zdWWdeEVQyaO3ITorbLDXeTw4/HaJhma9/uo0uHA5DEfxX/PujOM/Rm8hQPd
2HMW95kTSFVdLLPRwv8k6TCNOPcy91IGdb06hU4PWdElDSiGQVATFLREiQqp
i1BFvJJP+JIVUVk5jiDmul7zVNRz+HWQLRNYmPChYy0zv1RJNSyWF3KJQwh+
m5CtKvmMQFTnDSp8/supHN4OjAaGuPvMAgPfzW9Z6QfZ19UaLLZESvjP3s9P
mfm15UDtKyVC1TM529Pn2HRmcWZp78NuphmB/2Hezh+7UcAhWhw90KUy00l5
kyl8R+lVnW3jmriQy1SpVQ93tLU53eRqyPK7ZTnFJ8hyDw8qnC2B30KzPrkz
9nu+9KSo9woz0gkw2vzQSPJwu4MDbwaxkygTNVHET+d9gMkZHDfUHnmjxfjN
VOXB/8nzucSbmetDBi/FzoMhxxcUKLjQeEzMd0oZ/h2Qjk/KV/Iozbbaz3Qa
AwGY75Y5k+DtucTMnrgGSErvYlmtd0O458OK8mJE6JEzZj2M3eQPVMHv7lYu
WenIAX7XkOcW+CVZxYTY4X3gE6De6QjXBog31FH1jxygXwoIuE2wFQ7Ez1w9
gOn+44c4Ow5+kIMkm+TPbu7ZLuV8TAI6Afg4LgeTuyj3LtnPB3sx/79Bxyvp
iaXTgWKff/SjsUe8v1Gmtcqh7EbIEFhEsdtxdee5ZIjZozACvitmAW4UQU2l
KGdaC8EqswAu6W5unjDdemMUxHmyHCQIZ8P40kIKL3XBuYq9hy3PcMejDpTF
UeG4GxZyalM4eMajwMrN248Cki8EVwvkZl8afXxmLFFDxf9Ef8GPX3Hr+I1Q
J1FyjpqUjfNjQopAuWA01t3Q8i67ENF2UePj1dDKql8bZ+0hB0DMhCck5aHb
MkjBV0wQYQXTITsw286zaJp2daH7imGtlKuxDClstm+frs0D+OiPdfl3010T
7crZil2qDMwZZPAz26odGEF+l4YY2j/0FwIS55KiGs4otmrsDnPc0zi5H6QO
uNRu4RCXO3NZWJNmr6gV9oiBHc81ejYGertisUr2HlGEyBikbHUUXgHrQay4
kUmll/2na0rBDQaBX9dthXAopoH2198ZQE4gHHJ3HYJsXRdIuG9tQ4MUE2gg
3eSBxVTEgXvAkzdomnHWL5n12Y1Gz+sADVFa7ApfzcfhpqOwl5VrOoHsQ7VA
91NSKjFafHiIbxRa7e/jUNWeKhG6GGbLdMuHfn0nzDWeU0v4nzI3usb0ibWB
tTdYziXBxe4Zex70vMDGBnw//oi1SKy5s9zQpYiRDnrSdSb0+mOVCrPYIsLO
8qvn20wRS2gdfI3+8o8fGKkKSZc3DlZoAsGru/B6l5ilnLU2Bl5J6JbPHji2
+qtOzeb/d7wuU/y47zM8UzeA31553Sm6HZ/o8CyVkwGCb6UVtiEG/SD2z0YG
tQuGFfpRsyA5rcYJ1nHAtGnb8NyZ8zCKRockntIrJbLF7v3mR7evfdPxCXsW
PcPdldiSFLbanUfi56Qr9WbHtqNVu0r1kp1oeCJH4RAFIYAVTPqTf1mFlNT7
etfetESKFnLShWVetrPBZI+Hts18uFHVkIx/9pgMFAuXkKxZNIpxNVuwED/k
g7IIM2IPcybP/e6nLqjC8d83qCg0oGU/V6rS3gjrcUbmtfw5/ZPAgT2jnbx5
Ay/aAkJFz8IxI6Rx3y6mHEfiXKXCfJt6EHSQIYbOJhbQQlVex04nbVBGUF6j
6LnSXgMqUgy1xUC5iaAoibi20Lj0OLhpFcFhubLt14SBFxOp1WGR1Z3VQQ97
b9lyoZbwZeWH8qZB6E1RGtodWlEjUDDho/aweOc0XoUpVCFqfsJGng25PuQj
lS3awjHqiZ+9lvq7QPj4Qz4yeEUJCD6MKmShvja92LXq+dgIvMZlRW8G+l/0
8qrwAb5azKFL+beABrZ6UwRTOFhnXcz6L7ZOIXTRLSMCJ6j6+z2GdNOYJ4u5
ODC3wQOI1MChd+HqXPERr8HLopXqRxgDRrBtcLH2DYWPpJDf0Tly2N10/h7R
K2+taigJH2HV4jQ6yaBH/NmNGKYy8ODAIzcSyUFnihczSvO8/RS0XMZAZoms
p+xLOtCUlV2x2Tk5PsGtVCWDRS9TIlt+4R99G9t6x6e70CQ7fMSK53dPwDMH
P9/rOFoHDufncVG5VWm0XIrA3gplpRs3qOlwsmOt3yavnT5TFzpSsvdpJ5a9
kxNEWTf9MWhdHfL5ULFgYRmNKxg1pNRbsyeKbATpZFNLwADANO108gNqDGTx
oyzSUunjC/GQwIHGudzC2OF3skByeu7PCfYqpYv1Tykcv87mRbDOV29tPzCN
i8QgnUk+1JspLJa0Wg8/ffVJJZ4H61wjxbEaRGlPJicCzhsKmzC1Vf9rTpQ9
aPslD4jeVfhQySON4ST0S+fSL8nmtGdW997qnM+LQMbyTg4w31d/fdoHwooS
/Qw8ZugWd6j7Ke5g+O51h1JDSTLhjVTCEBQcyvBsJQ5BCVU64zQXo9+7FRfU
f+JyEWzaCoxfYAiWYPfHBNyzkYKUCYP+Pj5Wfg0tdbDXjrryPjAuEAtyk8rP
jpOs3JmM+1Ji7aQkQS2W3j8gOJdZhIcAjwo9IkNurjC6g6CS+WRLzFqLYD3U
wruCU1XBUjh6LN0oadAHWj1QkAN7CA96TBirwgJreAAIVSsqhjrxBasJZarC
6JooVfSIxlg/g57TIl/P5dzWN2/PRoOWC2Yxe1pznlt7noflqj1dLejbeoeo
FfoFIDRtr/6FvCzpi1ZHLR+3jCRfLsJhtfjtH0/9eRWBOqZDc1vtAIjHdV4g
hrlLoG1fMa7S2WUmpaceOzmAMqABla/sdggnztEZbLZJW94GDEiQBWPsmg/5
Pl+hMh/XjZYrdXqNvPjmt6yojkvwCCay/I6sYGxJ8DLMsi66VEpBH6pqfo9E
Enj91ikNdS0zT80AEN+QNR0s1TMsIt/w4E0cxz4kQF+yqtNom3LJzdP6JG68
+kCkBrMUWKia0TCJnzvgofVzrL9WRoABTB7k27VsjIpue80873y21nxAFOOu
tOwdY3K4lF2iieSKzTc8oee8exu/N6jpzB36peBLzhAeO7yPW7aEL0OgL3SP
BkzBsGG/5jV5d0wC3ZoaqLhDfLYz9j9bhmFUrW17LclzEu5W0n8xllfTQkJ2
MQitCnV4De0TPq0uuZqmq5uKQKS7gnsO6+toNEnbXh1YEok1qjS4LUXU3sbn
vgpj+XAmBx14QTmbsD9xbfUwyGjiQwnbYYsnYBkGoFJ9RDFjGBFw4nodD1ql
enkw6fic1gGDTqSv7ItaOWHX+W4+MrokVenzki41YkapmKV3D2J8Sb4Vj+iD
rTll2YQNhH5ELDDnfq2aSKr3mTWRuRg37uyiIJgZkHvVCBmpsOOZL3npYL+8
lY3ixLlJD5aoQOg122+gHRUX5NYicAtUsSZCbNv0eq53xPPaZIKmuq4R/zuM
rQoL2Pd5I0GVJZQhXcJaG1h5AL/48Tg3DRmuiwFjQVA8wXhJeO1/c4VSgK23
aJYFA+6t77RNlM6C0b4qrjjclpt6LaOl+QYXhY2WBxYT2qMxN1FvOiC3gTRP
LGGei3mRPy3j3J6imxyJp+rTmFJmE2m6tCQuaHF6QrWCekN8SO1R3Yn/HQoT
FXzr9HFOlpcDlqn8SPLfiwyBywBrIe7wffjeHFLkTKUQUmhbXzDJ77jzY6D5
dM/rP3oSJOaAm80EsaCq9NTZY0r2/gwRVKCUd68nh6cIPDANfyhxrV/jLPnM
hnoNMz2clC0BVdADXLC1+25mnslz7VfjMkxm2AtlsKlPgtOX5UmIT7lKWbCF
hLYwsI06/Bp1Xz8bot6SH/ZtU98t5/eNh3I8npeMdJhG2jW4e9vpD0qI7oiY
3ux+EPpYR8R0e4WT0USlSIqlCue4gDz/9m3hKjOV02edF3dBwgoFnkBiTO42
yN+EOJ3RYwudzZNCD9Hse9TlSraNWVyhkvY+P7EQdOFdjBJE5mArYSsr6otV
HQ8tA5WqvSNPJHT5HrZ86Rw7iZaoCMAiQksVFKBg/Xw7DtMEitLJDDKTG07h
dB2fyfHmaqbZid/1IcNYrY1q1hNt50Z3hk7EnetJUc9tH5vhln3ajxc5glrx
7skppAha8BhW3o2PYzexRXnRdohrRCfYnfMBMglBWTO/oosJC3FL0xMlobYJ
25XrCr0ludxVVqjersazy+thJVHKUObO1+6dxWu/5HM5lDMp0ywMagz+kKLp
IFOUcK2b/gEIk7KoUI7DxKW5DSavSiTP69Lst4/FNrZ2DRAc9kFj6gkvcyND
EFoF/cYCE2Nf65v6zDojDevJENfEmaa8zdXUboJ8VsCWBvrogiIZUDhVidlz
tvT1LV8k2gTj0yYeO8Ipu1Ap/Qkq5+6ZQynru/4lg7XdWhw54bacuivjGvFp
n7cgqYEWv6wk+2Rodqo5z3gtLVdv/0IE3IwR9FRpWGHx07tXBxHU+tOYvcCV
2XaBFQlwhAursXZ/RqAoh080+6qWJBvMkoNzgZvshsMN9PowGQVq4ZNVBERS
DnXdxQ0sHtN/fL7ogCOc6b1xPvizf+T2dxtxL4BDjvzrujWu9WRyjnSO0BIx
2QSSTUYE6F80ZvCMbf7skdxa6m9+muKnZolIZ6f2ZgI9vU3cik53vc6sdsdz
KUyL7ZRHpk/9sc09vEonsgK7WZNbEsS0sr38I603Y+5nT6bOToZGgtN1pGmL
4A/sPnGlgcvm5iY/JYzO6+wsj1WQyALlkXv+CYPTOhnfSbv5i1UM6Z/k8xsP
OMjcUsa/8LoRA4kUK0l+zAihfgYroOZJwFHh7eKS7eOszsL1/GD8yv3toigG
FnMhxBTmLSW0UR4DQjoSB6k6NagQpHrSwJUCAycQWnoFN9gnE30TdDIJMrns
NftAdgNxPWHBcwiyRGjnSNk/LncuPCdqsFNMnrCw8GVABLo9UuLKCwuToxrG
0kIx7+ux/lvW0Hz4RBv0o6hktTkq818k8h0bM6Raf4Uas2ziStt9xuTPuf09
ffd4z2xwnnGoYfsr0+ci6RI1OHwDhikFFkltXyBHiUsWn4koCGdXsM5IQswg
/WL0K1RURsbqepfnFzRFXnQXF9TVlTiiaN3TeSdKbjHaL4A4d7UidLRLy8a4
E/VR2yurr3dUx8i4TsiJHVX+R/i9bGWGlQbA5KuIPzECPh8SEDQGfOwmctfk
viCWnwjfaOyq3WLJsPDfLSJPZ0HK5sSb5SVA0Tp+HzHOIkoKZ3GHePj/ExlW
dr7qMPGbS2KzFGf5NfAiWZXbk62wpJ+y323XeYV3hk0lSjAcOffAZ2d4EX9G
meFQVNaHOPQaw4MrkadxrIBUGSAiMYIAn+ASGUbKZ01Qhy6YwSkIQSMLUKxH
5VNwTGKcQV6LiUBgUOQfnTLuW1t/TFtul10HjoVcB2Km7MekHjUQp008y3ET
IWzSPeKBbG36bRgejHudEuXAjD65MCBzmkhdNlGApAgfX+7Nc8KgsysemYOF
LmO61kKEAqn+7FXPdwDlppPARyTjp3sCTHxFC3b1dcx3GlkwOLdphshT1vv2
OhyuahZ230y0KPJGniuHI9hYEdDTc9ohAhwthHfdePeLEmFeRsqKZZoKtiAN
OEiIE9EJ8Qm+j3eecfYkNTM2a0lA0LWBXQL+kPgnOqoldQ+vJrEDYjPnX52H
nhcuNaTGJ5ZBalRES1Oem6LTo2M752M60J1eoJCtVtpjj1Fe/8ifRs/ejyP4
meNAbCPBC4MyUNWj/A2Wc9WvRSKJs3ehFGnrjuQdIkHqXGsk5omCRgEMqPMo
MlSJ2aMmYWnJVAVQk5L/udzg4I6AHjrlMF8Rv/bJLr1+12+HtPzgZzT9UR2J
2Gx0UV8Q7WPyjKS5ujOhTwCsTSq9dzfPZxQLDE1QhOhG1cvepbVGErTMpGBW
g7boYr5krZmFDYlyRaW9OHlFmomocT1sa3fiv73vP9GJ1JolhuNxiIi5UUfg
qUU0RU/jWq4+rdhitbUqU+xWQE6zbpEISiRLxP3wsZpcyV2ZDhX+iIPvBX50
ppOWhN3XJy0jMhr5qUPQCDPv7twpTu1fqvNbPp1x4OgEtd1YAGE774l4R7m4
XkiJ6M0qhDVBbbM95QGC6lP7X8SUwXnZV+sa8q/n6sP+H3ai08n20UX+VfCX
tBIin+xQrMsVx/Z1WtBdvnVaelrmlQi+QZlofmXzYAnEZh4rbjfXsx5i/CAj
eFk2t0zVtinsjkXk22TjN6OYE9si0aLws/v3iNR72KX8ThGECbLa8pkKEAB/
PAzKPf8S/Ck/d1jJDML/EF/PF4ejHIpOkV+HcMgMNyXDlcitV6HDKYfqolJl
bZtjtFx5TlsX7Xq0ZJaHE1orKvb4uqmrxnNhQr+rsnWSUHlpqj3dedmQ1G44
PeVWQkm8/L3+CYyHKxOcngEVnpyBiECJSWtn4jcaEZWNWAkX+S6d9yANJmYf
HwC4+yta1fpnQC5BQa/raMq1ECA5ingg1jBBC4tDqMk6fqJ0ZvWIGxLqht27
jHQ6HALwcbNaa8js/IPjHgmp70QDbmj0hSpO4CKMBSDq3ubux2oylKPbKeaL
NH4KCgDAxf7pd+eIL5iPlsPvC5eiWpWihTHaupKtRE8SzxcygSMXV8fQWU1p
/PkIhqPIetBeS+YfKUGfsQvdACxU3NzwC1ClsqkQXcwlwptq6VPMbH4uMC9D
0YqRDDm4azmIpYttuDjdbyFq3o+xU3rXbJhusoOoTlWLM1/fqL+kVEIziLx2
+5rW/pUjuzgBMdjJnnqZtaisyT4Y+oCagpaw7J/g0zpOQf7Iqmm1O4uYpicH
K3JtKg2O3c19noTHTXfDLoUl8kGy+r2iqWnQjQBViorSMlLKbjaPS6zYyw5L
5bifzK4xg1Eyfu6UnBk1Mo4cG7czA3QjQnC7tTMrqOK138JvSezrxAs/e4k6
3lNbKKOHI+30iT244Rqh4NAGM75ZLFnqNUI/05ENxBTAY9/CkffQJlYB6QhG
m/Fk8SgSq/oMKSiVpzR7+7NlV1VYW7w4bX5ieY1kwjQQB4tfLFk/r1cE/VrH
zLNOU/0iJ7VnCNDIvSxDLW1257kD5+xNYepaG7fL48PdXdf2ij3QAKVDYNG6
L4kLmqqMfbQnRYsIavfcuE+q3tB6ymlL4fmpVS+V4veBYzfiagyBJuJAyLC+
sRuTy9LySpgXUmExhSY1jcDWtpI35drp8D5qAfviR8q/pXEN6hYHmhZg4m3w
uFJbpUpNfURSi27anpU3TBeAsVaqc7DlYixtyktVGBpCVBE1JTgrEfNrF0e7
Io7e+iT+k4YHeEZLh0bU+RfTp6UL4qUAeU263lbODyc9b50SEFEjmMxb+VcB
eIambMne+eyV6KTSBrgDb6Uc5/6yNSzdYLyaj0evauJeRaQ5oDpU/vEvPMTP
UxzxSvg9u6A4Y4Hh20hWhd/8B0UGbeF5on+/5Ze2qguSlMdxA0BgA1zOMElN
xfjoT/wVggwegINt21/Dw6v5TDWuuWIX6pgVISZEXfvTwUh11OR+kTfH/6jL
yLuMPHBjMdSNcfiyesfPIDQfXVnJbbXdEwfyTGIc1JfAPoLp9qwFuvVidDGm
fgsFWpLwbGNrWLpjAklTIteObMZd/5fgPnnpOAiTXRP2BJnJ15vFEV1ODxgD
5zl49BMvbyzX/rb9uBR243R908XMXA5/2QOzz/e9yCH7ShRx909AXUHqEBcb
KZk5duby/cCtYxFGcLhStTPy1s+3H+ILAKym2u5eOa7LWLw6DPSno1Opc1XJ
Dw0hpN37l7M71qUWkwsSWSS6uhyt7l0SVA3hJF/fvJIfrdeeGVyd0lYNwN6E
AQRJXSs/eLiWeX8b3+bhMHtcWjYqOjzfWP1Mh9siV4GORTJ5to3QTW+FD4nk
UTuycGVbVzNlGPpT6Tt1q13YEVYr8JiDwWVNfaO83Eq4ibuD5YUADjKhyLzu
3hbKW8V1IUHLmtzGhG6x55IK6I428ILVDEwNXCKeMA1w14IUdM/usBWIlu2D
9pY9CEwME3eaglqJbeTa32ffW5eKebeeVzDHs0AYb/Hegs/h0M9i0nMRhImf
QDGGovByFwWqaawbPoVd8oP/OgOwSqsnmVxhrx48vsmJnQ7ueuIYF4yzvVL4
SzuCsWoIMU5sVn1JIqRxIiBpxGhS7QoBnn09B2lyrBtKiWQNKKZUC+gHxWy/
Vn7EsyrE9TMvuTdenX/KcAS81bmWy5aIA3r67Zl9nJZXvFi/glONQURDu66P
ImD6nZW3BDpP8L+EfO/HVUZ31J6hVZ805Vbt2RBkgihBxiMBthQRCrNHKkKj
Pa6soIQAa67/8Xq0eXvapgOCvi9WTMvrRtD/PoVoySzVT2L2S/emR6GopMI9
kqUUSUfVq3XXU+9e19ge1QdY7ZFaXhZXqw6tW7v7Dp17DrGK70CgOKEif3fx
6TqW+of/yfHr5GaNfkIZt79jn8jL0L+4LvtCBB1YNSwvw6KM6ajX91A8eofj
yjfV1wEniStCv3N8hmdLH1zuLVq7hjIl7OHMczVMDIj3KugHanm+APwnTKMF
FOJ7tGqtgGGcPqxTjAQ8OdJI/FdicalOv22tt6Aa4Qz1SRNA1ZRdXX4kpQle
Bar+HAV30ln2EfDW2ESAvf+aMSzUxbEWPBm0z25J+1X/rqHsealhp8J2a7hL
kyk44XUWLK23uBs5rjzriaQRL0yMUQ8I7URnQbK3AwNdEMhYkC1nNaMq5Rla
F0JHL0ogRzAPRH8zLopUVhj1KbUjxgpHCh03F7rz0DEly6LICdsLRSdh6cyy
1tGN7K1eVVFYxGQlmI/+9YvWUi9r4ZmPHZtPfEzTp/kCjX5M7lhD9B9QbFNA
jZ2avGBgVQGyXA9ooENSqoT8UOVzaYfRJqOjRXKZ8uJzzI6Rxuc620x6NaB8
ztApBGPEsBX0Hubwg+aEuK/fn8JyZCXnpGGVD0usGUnyCVjpCTFy+Ht8HgKP
Zos2eXlNqkqmsj/hCf78Wg5Qlo+dFdzvSxO2cE6sTNnkbnHFtmNDDaQ4PqKM
oMVTJH2r3u4/stiMdWl1EJlZvxJY3xS5+V6d5s0HgvxiGKZ/GJrPjDlVE/ew
z5h2mPWYccRVPxdas44lDGBbepCmUn50Qpd/y83Yw8Ig+nYSQanMa0DxJgMv
b923+hQf20PzqVuAagFz/ZGqjmMSvLawdWTAe8wiJviCel6hkxDB0WDm9iiu
olKXDLvKpNxyRnWLor+wr2PDYyaAhM+jANny4Ec69RmO9A7mzvufQCD5vkkg
wOTEMseSORzAVu+XNnXP4Ryn1KyAcdkbgF5eiMsnhOynvWhtibcF8TaalToh
cC3bFFVLuUY1wGNjq7Cv5XUgk2r1KbXRqJkGw/Nsgz6Zv1cK2RrUax8BlIhz
CLjSFihveHvM9UoF2Ndg9mDxho95tGKqlppxAxk6qhab5YCgCbyVL8tFb9Cx
DlBPEOE9clbos4Qy8H4pxkm5y+zftlyGOoph3Fs4Ib3D4Jh3HCOCz8eLivL8
ir05EKuASLYQQqF4i+SacidGD/RG+fXe1g4rewAI29XwVIT/vEy9qMlJqUcj
06jAUR5ryO57Asv2DTD5YUc9U/HuK9tbWPwyALO/epMaiP4zueRItUpViN+j
RAHCC99ZK0lPP2NaetopujgBZgj7wa75ZuPU8CriwaikMsGRx4ze66aY+May
+Ixl2j9I79x6+T2OLVzB8TuaN4U7NRG9Jv57L4pnlWOFeLLmsASdPL9W80tD
tnLV2zyME9jhaX+duZEiItvVxHAdlLjfA8Z68nEIgYIB/R3twAydb+BCwC6z
fk3ldyDbkm5pn8hRHpzCsxdMb/wyc1qQew2K8sMa2JhpzcMRlmoUnNfiQFMw
AOXMWTPx8TvNOqlbkbkJPNquh3UHQygGS2uPwvQDzezUEEM2mFk0os+FQa73
S+USVD5ZgL0BV7eM2QEx07w5oiOQXYtpbJ/R9aFXgrrKJkyH7v7e6LiYh7pz
J9VdMVkyjG9WRjXa4URJmOk7+XN5bqLM6GiGVJRYeewKhifcnwj4ZZACKnei
Bi4K2zjxXNxdMtJwyEEFbKU4JXmTHb+Klg7QH5ZoMYpsGoJD8++dS5ZYor7x
2HqO3KNj1b4UBniQuBpwhHUqjFviersAhk971Wx5M8vGzurem+oC5tVGlqq2
lS2w2IZlRxAnr/S44PqoPrH4LZHX4ozUrNLCnqtaZyla6YacXq3UeyTQL7ld
RzmLhazRR5QIwVN3iz1Ayhm1C7+8Rq06MAmPYk1UoIP4+zavyQwkEikqqG9f
OYXwS2oaRqy2sobR/wn7qHWhlVTejkD6HLg9plnX/wYb2dFo61ogB3MxFO4z
RyqrZkPBEfg4Km67g0QJcChQ7KTMKXu0D+cuGL1inLxzU/NH+rlt2ZGB65sp
23TOj3NnCkjJ7zP48m4pQZ8onT6mollinORQpvtjcK6o03If563x72wUp7Qa
Rl+WQLJGk9edtwkgk25xPP3RlcSh7XaoCa1NubvSJSZbdZLVNoF3Znv1WSAR
lEMsPKOejbvOC/IPqWsWEAihsRS/lYcMkIpmTSszQpo+OaPaTIQ5eVRvd/ll
PNICHOLhVTDz3e5SlAVWDF2tBb87JEfzeqPZ2Gr1jZ4RwJrTwID9jz66zBzu
MEDXaTHSuUfYRJmfH7arTqp1B5V8/9xFT3JpCHla/0IjZ98/jO+FA3nOmcVd
sIqBVsntDaP3g9/8VCkzszHCw9maPhQacWYnldOLy58h6CMAb7ICtErBOoJA
Rwwg8CC3p6NT4v2Pyi6aVwcEZbVuxKvpEkGRensC6RLpDB7/YcnzZvI4QxqW
HPLxj0LpgfD1NXR7kv8Lhc+tyd3BtJ9/sOCRHlkP6Zs9Q3rUBa8nQ0EOEAHH
rE9k4/y2gzByXmPDUshNhHMIvTdbydNbqyu4mQnwxpEsSxxlLNI0Mzrw7+NI
Xx9/jEBfWtSog6+ugl68uF6L+hRHRwxlxL+90DWktqNF4iOmJNuaQKovw9oc
ps61AZb3FBqAWlD2Fsk3rn2Po3SDEq/khvAj0g1hcl3RYzCcuRK/Hdw4tJ8n
18ML4ECSVNO9XKBgp8dd8fDYjF78x2S3XNko6i7qHB3y0NF/Y6rGhsv9a7B7
QGa+Ndf9BPNBzTwz+w4sHG4M6e7WfmY26tBVIVNzz4tjiyDjnLm+tZDGfI8z
xAabhypOLnw370VG7Qn/K3OOJnsvw3TiYowtc5+hi5vaNA0UDLN8Jciv6BKZ
5Nwoh8dYJo3/McYQbxfBqcS0wJsdZmE54fqp42zzPWcdVUCa8AMGdorPS/tz
eZG/JCmE6qX49wg6aH3QVRpq32WwxXRfOtIeKbvHYHEJedI0+J/S5w4/EL5z
25RAoGTGxEHq80c2Q4NEjDI2xKLSAgv9ObGFtuLHQoVmmSv9PpWovoYqbrMA
rrzJveOmzuL1YaprtpQ+4DeZ4Iykx+VA2JbAelofqa5x/dJW6ymHRkRwFb7x
vNB49kRqnHYout6vVkZoOK9ghT/fhn758XM9qR2yF2wehS3yt8pzmyZ1EEuz
bylXu1msr42EtFZgexMiL+EJ8oRznAQBZBEOl3k9ECIZbfKPQm46Xz623RMV
ZZYDtyYOGLrS7S97cRrmNAHOybTD6W8FYzw9Puo+tnwSYYZPoT54GnuB8MEo
DAKGtVkGXZr8Tj+1M5UT4+PliTGdvKshS7jueEIvCDhUOWuiU0BKvHKvUSe3
1qROlvTCOi4/0lWjomwHPYs9Vk/2itiwAY8TAUuT5RGzAqE/blhMhh+S7OPX
y/Rw8Sr/jRpWpQVJUOEk1VdQdg83qARYyiAb9WCWZaZjEWVpplZWuHBxiQs7
pcibrQ2CLH1wCBUOZhLnzSgESp/IdK82CECP6dCa1Tr+BbLdYqy+FUejcTfL
41LMwBETjegWSAJ4CdfqH4t7M5DjAiewY76DLZp8LvDM5wxD8jMHNHT1XSQc
F1bC1jl0PdUE0vYXVVzl43oI3pu8alZk4qvuAT3DwkQM1FS0aCCu5Qrldpj2
ZKejf4mK7Cz8LYotJHf8M+uBGIQBCqvBYDi4DwtwQfeXkYCcOt5ffEum4do1
a134GZ9pIqgkX+iePQZOfDNIunb3+qD2n3L9fqPcyaAo0Kn6AdG7mhLe9NWJ
kE+DWcSgo9i5jPfBEqLiryldWmHInf7Dmr+G7ZwpbquJDS/tHBYCIpkMcONw
OweEDR1HLwWMJDR6wBvw3usPzNDcPaCAC3spgdOJAgY08Ht4JppVec4nlkq+
9rsnS0D8r/qtZCSWQJ/ijOBFmHEkfA2cS/8psQ4rWoLMIq4B4gIWkAlfWrQg
gKGa/hX5gZHLvaaVqxggep9ux5aY2FKxOggKnG3HMlLH3wKVHNZnYl/xIdSz
VpnD8u7KcHwiHELCqG/UU+cG/WWLgvQFixmP2rca31/x05abSWR2WvHVYfi1
zTnYSLea14dwkuYFvIypyQxIsdsEHJfmup5vCcisTDqDijLZSl1bO3gkvdQ+
ti+wlihvw1EsaI96ll+vZ2ipugU1M69E1+P5JtALJNro7MlJvlbw+gjfx+aC
zS98+cXw/EfGzhJJsKYBso+QV7zCOEMg6UsOST24wCeXnWjSyepm+YJQOxJW
DO1rEV6GIZEi8AzORaSq2VfRcRjMA9AO9E3wLJDmn4qVgf4yVX+9R2W6mKvX
ELD9iSDYp8D0uiuUk9SKlR7Wu0ARzv3iw8osUq/5gXy2RAl3BOH/J38pTlqO
t6WPvW4fBjNzbp5EUoScqNLXKgrC31jZ1Ygn1+W8Hty1k/arFnccBsYDtFgG
EEs1Wf6MgrmG3ang5blpA3kC5hLJy5EljFiDrfs1zPvcqiCYUAjyuPk9TMNQ
DIyzC2avCCcy6de4BfZWUIB27Bae3/hk+F1iMrorYTok0wCV57W1zwK8+4Pu
H/2NGPr43BIMFR68NcybMmbYHwec83rkpW5CNjXXNiHG9yLFJ/YDfVu9TwUd
x9B3Nut9WOTv1wWUQR4YKhYolyrR/x4CH6Rb1rXzgLu9bqfyzq3bj0qH+wJs
rTjllS2HtDu+ZI9wrNAjqV3zkIWVfKYOxbAerP03F++59CJ26++zvpF3N9W8
rdK0ujkRsgfXTxo45I862tcex8Ri2QIUH2WmjxreWRqZQ1n0DgHr8Mb7iy65
wSLt+CeG3Q37Wi1SL0pJiKqefivuEol+VGscHtIO+zn0vQ+IqBBXAIRJZY2z
QxTby36/Xz6oCfxx/GMMg8on7yrc+O0keM50ZMdsKiR5NjsWIROsXl43iRi8
WLLT7nEmkhB/UV/Auq24CqkZUCgoQKnEHl9obJcjPNZdOSUsnoUZOr/8/7uh
BiQyE1QCM8W+AOB/JAxhT061Qr61pQQRQc/nGHFh91kZCFzo7t8RG8w0A13D
xThTESLpqRctlm4I5ha/3dWW2jmbiKJSpU2oJ2xtX2CKaV2Ojt4PIOON1rOX
u5PoH+7NB6LQECuOIHbrQtX5KT62vxYT7sCumKT5pZc7zwKzMXEXObqE+YFg
hempFsLogPNIxDMxgXDe/WlwNgkGOHI6M1d2GGhh/EXimaJcDmF/jDgtm+J9
3DrEtMe/+eOcwRwLaZDawKgich48WjyH+sYa5XfBzttWsFScpbP2DrBTq6x/
c2CndTyMEH3aUlnHhLfCLhDdYPFjxDh2syYbw47PrBAG+x5qur8e751X/2tV
3IUYZKzidBJfW8T2a485/z1PGztU7cNhvr2BBX8djfgT9I9qPWqa4rFkzBOm
wzpZ6sh8/a6joHO6w0fu/BXoCRZIk7oyOCmHGfBdlmiPrysLzT8Dhs9UyNml
OXpz9uz4FoedEYUNRKaal33G12phmWl+TSry0KXai6xFEOQGpDORkG9ZNGKA
kcLwQvdGOYpdjPWgqaN1gdgw4YGFQt+Fi4TQyU/qDmxyvDBLgM2mH+ty+sy8
oULaa69VwvfYHeVg+/gYQvNXcDsNeKDF2rdf+xj0Qn6RwLqUz9AI47OVkd12
eIzgVPqlUmk4x4JEzaV4tHa1NLnYcA1pxpnXAfTcs2+39u4+5GdRhvqxCXK9
zle0pHFvtvnFIcS9HKdKN4bRM7WVfB+ObULFx0gYu0qc1PFXe8KCfJRi1DT3
wxNrkEIz9wqp7hyRxaokhs2zs9BhPUXlQ7VM1Gb5Go/5VpT/btEacpHrda9t
zmpoS8Dacvseo8EMsCTjSqUHFBl8od/hrTqii1zng6TFMJ4tTC4af42KpCl1
FzQgSzNAtfLuwb83E34vi06uNKl/W68DNileUU3CospW5RCGFT4A7pTRxxuu
WY9x8dj+1raY49yJhwZ8i7gvcOw74wky6eonKEweUhUtgnu5zppbJcMzpfE8
+KNj00rERA+QlFr/iFiK4oMOt4/XszuMJWQVpvbaZy57Ep/5hhDDG384U+rK
Oc9rXLXQzEPsj1dx16sk/egPl7s+XvdmdNLQWgMcSBLU9ZIH30m4zyYVjx30
0nOyyRR3Zxf8nynXqLNUmRj4j7r+lReDH47vy0co36dn7CV8MoEBcJnskNox
6mZUayX9rlFfAh9TRuCuitSzgZ9K2F/ku1zUyBuxEyIekWFc/Ljx8+y5U6dq
7/gQHyO3fIw84lFoySdQfRgKUz0k7Veu6vA2jE3DamjnzvlQdhCLRL22Niiw
g3DSpEa7aBQJc9IRvg6BbgjDsIepXsBo0lAvMzBC2YupIc1vP6d4aEVe3/gi
TdKJTWz8LjdugqjBFeSO4RX8B+YFp1Lw3yKYt8QQ5obeNv8Pu9X3cM4jKcyh
4wx/LLoU4OwLxxfzQalq6wTVjGP2CkYN6L8yIuke8IkN6axdeyd6Rvt07mZT
ihptM/ubSizsQuOQmLL0Kn+EztMB1c3eGpxaL2qZP8Ufs3Hqt9b0TIOEe4lZ
S2J27SDlaM8SxaU5QumlahgN2coO3Igb5Scvku/ENUHBIyk4cy6/s0nxtpa8
L0Ki+XNDIczokpoG3KkLGgts94O0E+WX0LvYdVhUsYXpHWHKEckXV5mGaVNh
GSuxNH15LwjJeNQzhg11UTd2Toy8qGZcdFchkMNLd8ioNZY0oNdjT9EESbbo
ZCF7mY6dFczsoEKRiiaCXhEJ54lw67ekI/UClyDrZGNDhcpi7usbnIpVO8Wq
umc8C41734BwvzXPtZ7qv6d2VCRS5N1ACCwf2SdHMuGoNuWY4UtYD8nc3Kvd
tThMcjvVn6p8EOrQJa6ZVdIwAgbKPr6+c77tLGv0z/VMCIb+lhw5HIWizdQB
/Be/KVA7goI52ANrtBBerRzzgHtOtGKkfKY/9mel11LKVCZhDl1rMl6Ny1oH
xNRW2o7O2lDIwwh0FCy1o9Dx+9XFvfP52YbMZc9S4kVXwh48XsdrSdZgC7ed
dKcZsVevXBZnaJYhxVJKiX5CifE8TMZHERJD89e4WJOag/H9awfsuVH2PCej
G+PCcN3b6rfnnCIKtVdWPSgFGiwTks+MCo/arL5OYnWPVhuJJWUlVLeoeSm5
ZTq/apsbav7pQV1I8QQVh0Z6Mq495ED8tqHjCPduL1E5vHeFH2HbsVhGVrL9
TSE+4ZYqk2ySOpEO32I2M1+HVxijTHhZOzhnXx9N1XTFiJoauH41/ZF7wtMl
7h4JlxoT54IaSCETMeRL0bl5GLmZIlMLMjiSQtke9xCjBnRo24Vy7BJryCwH
mtqxeqRVWyTUkknc/1COahfMtsBYih4z/2h7/SzmRUmW/zL+fPeFjacZbFOg
v00c6DcQ2YDgi2tcy7lSBxVWK7iGCLnQXnKJb9lJd62pqhWbCpfOu1xn6xP9
xszGxUcm2O36++Cqy8eYdWL2Ad8ZODEmhvugbQ33UEqFM10DMieXolJzTIi1
TCWwnCu/ySD4LZBvm2QcOTsD6svdZo04YS5RfRCFCQlxOav87cxWo/Okq4pA
8AV6O704D3zjYIixD1e0vC2gNWgw+rRgB8rjg3jJmTls6qBVLG5quYR+wkvp
/jKBDB0Gy3zE3dspeHholJblXL1uuKehfRCKCzBENA2+WOa0Ro+ok8PvF0mZ
SRMNC8MYOIWsG7v9oZo6sf2+xql+XEbOonuX6+qUOqYX7KodLqnlQtm1E1IZ
K8NPdtifeg/CXamYjCSJin3/dDY/rNl3COLdYnbyKimD0RBgM1LQT1IDwKQY
Tuu6jAJUsR9F8sP6MraTph28nfXBkjgf/Bcz3km9TaK09s9trRDSQENB5bhi
OeM8wv4Z65stBsbOAcPDWZqjG3bNWHSJ/5ddtIrCfwGE77joDbzaXRyXbj1b
yWF7MWiwEwWptwZiOGp2Q6OpN2YQdiOeQUlsUlO+6y9mie3zpvfYXJ4ZXJZw
ktH0OtPAmXito5Z5QyBRT79a1Yrcv4bjTa9OKHDrfciMi0HrngyAoQeWzGLF
soxoYWN40o6SMgRxO2X7b8YPOy4yp94of6GmpfO0u19g29M5+7cKSEvPwFJD
oktKre6gQepapyh2FzCkOCha2G2QRGn8UDu9hBWL1RGniW7GhpKZwTQZc82u
x2NugnXJArt6jshatbG2bvpSrmYYq936SOuE4DqeSSJXPRVTwukezOHBEu7R
5qktUWW1esH3gHlNIOX/olpQYdu9TG9ii5j/jlnpe8AtlJ+P8bxWiLFsszQF
cgGGmwGuza0WZ7dO55r+o4dwJXaldWdUkhlgKClHmGkR+uWt4CvJ3SvaWFa4
cb+sT96r9ztgdzRQ7v+qy+T3EHgY9mRn+D2ek4TVVI6VAqT4kJ/26IedE414
/MuB6yrcqcd7nlgSZbKdv7gHMxiZmWTL+yf881xF7anaaMaLPtzz0/xH/b6B
oE6YLmTJFxJADVsyfHO4B5Hfpf2byi4+wUYFdxJpTOVCi7PlsXi+Zz26mLoS
lcv8iyjf8m4zFG+TVJSjBMyGQTiZpuGiDbYMbaIMv0KW5a2EfvfpuGWVgMaX
4TE6o6HT0CqSPVsM/QgscE4PG9Pzs0xFzMpP9Ilb+qTnZPF8cy8aK4464JaZ
5mvbINDR9y3Wmfl6GlvEHIJDcGgSKfz8VrBfJTRUcCI4yRfFEA/ssYt4xMnb
e1AGCc0fPwASMCukiyu2seul6a9iyDIndC1qkRG2jxexo3TsuqK+x6PWM0o3
uFEUb26UtHrInFaeHRrWlkMk0fHMEfXxGAlaY2RncdnOg4CVEAcIMh8boh+k
cq5DT1kI8PJP7XzQtU7RxmKAp7Zdi1kFoWn91QcjdVnWHQ2qIlQ/Ma4PzHY6
T024TAtvwpR290ReiG95WWHrZ7lGmA5JQVdHj45wVNpDQwbHXNKYXul7Lbur
iYHtVeyU7GMo/FyZZ/IQp8ZXrMfuShnanVLrdr68IMqosCtegDS42bvndReo
Xu3cGA5PoZYCNzUVTbgdC90oMAwdsyv2E+PXVO06Qk+F4jEA+y8gEUr6gqRo
ZQLQdHbeHrwmeKMSJxJpYmDIgja4d1p5Wm3ij2uM7L+aXrRiugyAe1RlmlAb
J19DA9ZiK/JNbxitFGOUhvfTvg4g6pj+6kVv9bt3ZBdyELrHD0tFY+/5jhlN
QVV2KtGMBROwGGPaGezefbR/FTphYE7j+hG2TwWui3n7y5ezXdGdPgWK5DQu
B3lQvhGvqR6EpDzfXXvNG+Tte1kmo5rEO1wNcVuaA4tyIfM7ECIHwZMsf+bl
+I/CFNvxZe+afNL1qAjJTGs0thJAZpp7m2CiWE9ZdKiqaVj90wCbaSD8KDOT
Nb3K+SItXjQbFfChVm+YYIsF9WZn92eJzZOTncPWA2o8K8iINTL2TlOxE17f
bK9rVmVeuWSHOth9xh06VVyFCzZ7jVJng7yujpRvplwz6d1hzflHUtjpAVEB
oZniHAIlTYJc3va469LhpHlQYjbfKza8wCmBC/GPen1gZXZJfuCAZo5YN9Zk
ETF6HmrVitOPhaHdw8X+BB63zSRHNZIUm4WGlcfOUJ9NMmHVyc3+C+X9YIr2
0+ReHEsIbgVTU0zFZQmZYVqsuSjX/aw2cxh/WrVyMDUGXDgBh/8fTaHAO3g9
AcQYPWZq1YDHRLkKlsIWhETHL05RqVM+QEVehAcXZFo3QvT1P0Cf9InXzf3A
C284aOlwwoDPvhAkKU/jslvZ5f0PLRxrd5wySJf4gt0e1YBgNknO5U4QsK6B
FNOUj7HEJodVE8L6zqKomJbEIiDDeX043c9wYNm5wX/wsvmdWkMD70/We/np
AIdTPloIUlC5lHdUpwLWeAFfRomWJV/shCY0U9OslRiR/qaB4UcRDgxOFm/9
VcKQSn5TMVonnpmmWwGWgb2SDgRGDQwnFcWQeFk9+kEKAWHwfo8KsFcgnGvb
qIhqNjE+A9+ujdeJ1mI1MKsDVsKj/E4bqO9Gn7X5IkuAfeAMl9fDqIcAHOKG
LF6h5DpHjDsr+bqZ13EE/pfRjhl9Od8n8EraPIN3dckIoyk2Oh7/ugTsmfXl
Czz3k7cA9ol2+E6ZejJDVCOnFEH/LAHxdWV0A2Q7WRu5MC1Y4NyvDtFv0ca5
5zuI1eUG5N/4CLfE5tO34ASTr5quQd2F0c25dPiahIcWM81D95w705d1vvQQ
gu0xgIG/FYFds+qxONwFfeHcNTfJp45Hh35OJ5L3x0961kbuNH8GN/JXmMFP
JB6iyYOO+n83H7WyyQwNfj3nGLlZg5siBOFyrCol8f6DrZnittaQDZE/K9Fg
UXXJhpj6ZUfZfWEKEnMumoMXcf25yToE2fv218yE1nV5G67opZp7wzVlJToR
F7b5wu9Ls9DSzBpsXq8yFMecDKVk9aE6fk3n4pRFrVmg3I5FDJgyz1Pdbqj9
VM9EMTWxnJqyrOFUJMyORXSwGAUF2AwAr4680ghhMdZR9eCiWGkkLD6bS680
WBMSuNv8WPtrNnwHjr9uqBKdfopifA2GpibrE2nMvsn4ai1XWmWLKcglnBbB
JneA5VtvWPt2aNa7FLDFn/GJsWWcnPgQtvxcvcwd3OdkiZsnkconO66xmo8A
khEhatslZXAHf6bl8yL5y+3FGcMTTU5QQ/UE1AdXL/lhhm/3JGT/oeYPA0AD
JfCz7TCYbXAzJ/F7POzRh2ITUeCEbMkGNMElpiPt/UC1DVmzuRFGblXskZB/
yUOC2LpkQpD0cEeZnsl+nB8SFcN/f1Mf4Q0ESPwT60nhZjEVNkIlPraVnlYs
q7rb5M57O/Z/+/+fOzLI3LGzu6ViaTMXN2Ww3+T/0YFwOr3q5yJgST8cuMg7
lvMqQNFsDrfKlGJ8gCQ9/7yAcns6AD2cd68HeQ8LQx6d8+DWQ8yGYxyGQB1s
2duocuORlJ94DhS4XIl5b1tkl24L7sihqYPtdegdUYcumTplkh/xNX/lCl6c
OQIF8FbEBiavBPcKzgYMricMVETl1MhOub83LxglPOfn7PZsoQ14OdmUTNg+
tTNOu7dA7R4crKJS9ENjvSPf4gtqpQ+bILps5yITKPZ3/tgd+DYP1DXnQovz
jPEWPfQVWiw4rSo2fv6C6nGjh4qWDb9N8P/RcP+vrXytvuiq8V/YEZuuQwXB
cI16LQIUjkt9JK9z8uEVRlg1tnRG6zR+iaW4QQHgsD+IzjWlrCAWrmVy0UhY
cU75XRnFJP/90kVlRXLCBYZI7kFToOOhXfpIMy7Hgq4wgqeEQZhKfN4LrPMn
vIDUmlPVB8y/tRfcSB/3BG2U5NaXJ/97bBa7fGQdTkNFgW+EYyM/p8a0obVL
Hs2QwLeHd9d2JhBazdhXDzo7nFUCFjk3Pa1NETcoGVish2F3j+XmnpfvyewZ
9NZ9V/LAtjau501YE4hSXqb7EVsx869gh7qrEUEkptsTgPUebUIAWHwRIhME
ohb94Nck9z3cuS8X1x8aWNELppTMK8sMUoWi6LV7MWoIHeoMn0N4kPnfE1GN
VkKK0txfACFM8GNEbemMENn1uZ4LgZj4m5Py4GL3lHiYlYxdyFNBERvXUMwW
9z7jnlj2rrEghby4p4kSnwYeEm4QtEYDHmF4LQ+rrg2cjjtPX6mmLUUAsAb0
/+kS6PHLm+HjshzurV+v8M11+MiZVA7JLjz1DZQugh+oznN5GSau+/9vTUCq
rozHldgJuFDCFiXexoNaxj07pggVvBJfYAd8phGKoMflUDbmx377YdHkWrHD
fje7BqPVLSaAu4aNrqtZnqJge4Q6veTZU40xnENgWp+6sye8yxxzyCeDX3aw
K+yNqFj4ICApO9jRQlBifboZecJ0H92tAaqOMcCvq2ufwLuLtCG0bIrFMr9Y
G/KjNpwTbZL0cq4FZgV7RKQhD2/JJWoM8xUkj7L4VgnP4TfZSj7vwc5t9iPh
U5UTdRx7S5Xqio8qT+fhPcd/gycn0qmniwN8mRsYE0Fthy6AGYX/YYp+ZBA1
RB+Gte6x7udkNWz/r0jEC3RbU3fo5R42l4Y9yTnmhT29tNyPGoHibGSLrpQc
LAy+rcyta0pP0R0jEd6TGgRql0U65FQm41nEUErVqDBiEBObLwwHtmEXV+Xy
rBVAQ3T5KrO0o33yTR/J9kNSGoOx9kTx4YaqjW7AndtsF61ZQej5yQS/xCJW
ebbEaU4uFBwDJFmnlQFP2oECib1Aryj2i1s+rSTGMG2TvyaWCRDXvVVdV77U
MFOFRzyRs17mr3hzYz4cEb5/UdtwhCQy0JvdkmoN7369E9IMpK59jCA43+WI
2SV2FPEACnudWfSTqojTTT0wqnp+ke98YPgleSVHAEvpJn/m9bNyIdDrMUyH
sozan96zIDuywS/Rq7x/mgjtG42Z9CfMeO5poVI/SBeazwvJ4Juw1zIsVwFS
rbpYTMhAVF616ZXwVxEONjVKoPjmjo4GADY414rcLYlr/4xCFvsakI6dgw0s
0cevmJPwVfveBOR0/d1FbkAPGfVxY83xRHOPDbhJPtLkV/SeYyOs6M7+TUrV
AagMNTze+lAup8GnXPlQaS7jKHCFe8JYBRWjYaHk9o+y8IFKa84JCohX+5vt
pH8R6ft4IOwwUmrNQIxhdcBMt0d2c/WBiWKnehl9J23Q9FImiIltSER9sLlM
3iCBEMAFcvibJkqjI89t8X/t8vNs7lzSoFw6P8czf8lP4L86htKALMyVNa+z
Mo/8Zk9n5UuyRCXYUp4cCnovCBq2UG0djyY7DPDib3WIxi3a6PJsXkTVOd1I
Gb2Lr4zLB2FQfKdHI73wrTdyqTABjZsd/r4duKxaPT0tjum2HKNQYyhmL0uK
+KHhle1KdEVyeIm6DXAPNqcCoIVa/bVcaVZ9Bxl1EcWFwp7MMhn3yoi0PQ7C
sJgrkrvte8qcqj4ydtOfAPH04bSHZL8xZBJZQ7vc/UPphScWRz4+YGWD921C
RYAtfGrFQNudhZdPIugpiCg4JGW7ZbC+ba0xaXrEHaK9yKAAQHDAciiM4Pip
ttKP9K/nJsV+geq/LFDCknQ7yxLfBFZMrfiMAgtNo9Z3RarkTo6FdQwitb4o
HCGJsAP8z7aE3HezBZvVtRew4L69v69lrNVjNU1335EB43bIhYCgCX0JHxvN
dEJNowbdqFiizQV6qqy9y4E9ijkhdwPheLFUfUZa/02cjtvKp4V6abd7gXEf
/PcRNu9h9D4cwD6t6xeT9LKoTbS6I1yTIVBCw9LMabdWdU4DX7BRnHJQ/3/x
HFX+ERJPM1rYn9qIwf+9xyEgvpHI7ifmabtPDEoyGKp7XmZ7ewS5KbFn/52p
xIguOrAhUj36aFgevwALWlzQS5s4C4oQlZeIDfdeksJVOVy0Ga/jqQSTvN+x
V4UdHNP1bYSiLbrxTeerv9vSFfw8TkSPney0ISBLJKGuon/ZSFp0Zr8oXXJC
hrPF2l49c9TAIYzmTkxgdG2u2Y8Y7JLLR7aMoR7RkdBlzV7W4ninYEYBQzys
4X8nME2PXQwlP6/jj+LY2Q2GOTgtOom3PiuQpDATfg3F+bsSTjWwwhsMQjmQ
lbWz+HhBpGBR1mykGCI5dZ1GnoCluHXilX7w+jxXYniyouhhrp5/l9UGrfIk
mWhxGOg4Wc16HVLwN5n0iVNn44t3N8stAf3IpKx/zi0OmHCbLJoxoTEZuJye
UQTUUb/FWGWh+Y4ropNyJ+xisPVFaxvcfbWBvPTw/s0vvupFTNZEu00RsBuC
wy2yL+/hVDaULxL1YiyqoZ38enP/DKi0CKBg2qbtEDzdbNxnuuBJwxP3oVfu
UHdEGjvEAvWDhzPMONceiYSxorOBoQ2P6SohfdfYoROmpr3mHsdoO33/pz/R
t4XU4Pd03CBgJCdpqW2cPIgp4qYIgBx115IDGtMA5mbsQJfRPLvimPtvESfY
xXlVa+tTpmwrHAatF8yFGl5iOLDAitfLLju4EerzJ83nozZUs/2aifprgJwD
CeBvcmE+kkB5T9uXI3RfmdOjtDN1pTtjyzmWEWGLZgfugKzbcvjL2h7YS+en
4UPkHs8qAh2HY0Ew3/qDtVlqCIAGiridx+a7BTNs8CQ2avnrGalQYL+DOnSA
qrPBCOFDJPDWi/zBopmz6RkI9g0AY3z6Xrot5a9mvcRKQID1wO2AAj9UC8o7
doWEvFXRPhSMidU1gcY9Vgp2sZmf2Eh54EWq1/Sd80fzyX9e5jpYIqid+mpa
uu2I4D4mD8IA1HnofeYUukQnHJztDmYArxOn3pqErhR7KewzMqIlR+9AuIkc
0UsXVM9vCnZ5lGj7+5E3wmjZgwGexT0x58zVpb9IPExrEgcA7Z3NiamZZsdq
9W01Ua0ehxqqd7FZCLbEmunHMRT3SOns3oVNmHMvYaf900Wjv3bstnb/tttA
Egj5F9/Y7gQcksnGWmcatPAYyWspvuxkWxLEwJ3yavIlcIpBzM6e2BFwIG5/
H0SbV1r2Qq3A4OC848Ql6yAVfJtkv5LM36fFTxZPvgX2Ro+nGBJ/RyobOH9t
OOKOlYizuvImFnjx+rChUXaP20zlB9MXieMNhJWXgMxgmEdGIPuBsCiDS0bb
hQCz3uEf6IbDo5avkXA3sE9c9vZBVGt91Z8Lc9itPDmYq5+AeApOCh5mLWOD
y1u0vXYdiTOrePiWbLTMAtrQ9UwRozYFL3IQCXuJXVHoPbP74sP2iXeAJ8bw
EiZYx3t9YaStYsOVPiazPJ3xZDIlp9PL/U6oazMVHeAIlOeC9z5z97I9xB0k
RJpcFtp1kzioRM6QnjhJQGu3Gp/bO/0Gwd3X/2B1mX/HqjDViaI5tDQ/jNGr
e9loI8ErYxzZHFs1pjrgxtKCX+ogIrnEqjmvF4L4FNBpwXmrbNoC34UYv245
W7c6xncDw1w7gL4cWebXSfTgiVTNST8axPujqfAacaaNbaHO4bLPb77UIZda
ZtH9M3o6AAHVWzA8Mj5ygSwVU0ri307APJz/7BpghV1lh2FdWNNbCE6yAwwI
fhL1foLL/FM9brMSSPBmTFMoW5kHUJodOzrm5V9QKU9rqOCcgp/rOmb0NED7
ll0T+r0nXl0SnJ6DzENZFpH+BOOMpeetGaF/a/fRN087L3+shUFOWUuS3x6P
QKGZyZILzRzrsxiADzqUHT13B/f9NPSjr0xBtHrRbzFWPPUOy1AJqSqe9Ui6
snai9dT6RyVngll9KWcjV49wlm0lwIwLDKrcA6hkjjW7OOHWF8oR2Rn7Mj3A
KRt655M2TKMgAlanCc6uWjZlK77NVcruTdl9UVWqu+R3dlq4cd5h7JmN2Hg/
bQj+pxTHAML35iO9yaA9e6TSvb9lQHd5ciSI+71GK/ULhGrMBT5YDB/g6cgq
/4ApoxayVhBU/MbwSuSLKpYXzPATXmR+9IifUvKjv3PllEiWuX7FDZpBj/qP
Eq+q5srQay99TkSWWplFVcEJMW4WMQ49uxN8PNPbJ3uPTRPIpx7qw37SRGql
a8cxIdCCpF7ZJWs7XG6iEuGXz1d4YDJoSoZgW24/6xrrybcGaDcfkuArgi5L
Tn7rqTa/PuPWKXO7d1Kpxk7B5fhkxlJU2ZuqSokqDeHHA+2CYhIjogkvSYUF
wZB9bIC67GhnJWFVJI33p2NE2uFA/xUQI4mDCvpU3prddOP76AZnCu4eCfsW
ILYwwC6Hucv8ASUlgtgIq80NNwdKY1wGqIetj8U80NzUz9gQ01up5jOnexDi
2izETo1z/RCvAvRNKslWbzHoIoqkC/eCIjjp1IltPi1n+m7C2uorRVmVcoo/
6ylXLTCeTPZNYqrfXoR2xyMwj9fsLxPpkmf6ogBO7Um0JGu8Jn1QQVzlB5NI
G9jqeP9eO0L8AMOHTYn3XfovEp2Md/B6DhCm4MmAO70ohQ45SNeUOdQhKnGp
GGGT3SzRtzF9fNLTyCQQ5O1LUNjCIwddG88t5EdsmuzyGbhk5nIpj3xfQY1x
OQLHR2eyQHI4SmDqGZ0B56mUTse6UEv9N9LcK7IJGLFVKvswEZ7JlKXTAjW5
GrpgJR8jj/NnOw1VoqpbG9E/yQC/xFQaKSWrJGXASWGH2XWwNzZ9WIG1lnt6
ntARVyd0MGMg3Bt720/2kgA5KMQV9/2L5U3e+OAp6NcAElgkQ8nSS5G4MaRc
vrc4cl4zRaTBz/kt9DfFJZNkK9z7iDabhZW5H0VzvrfRpy2SlxeMcasq8nW5
1N+6pACclerKxZGmXRmU8YiYLlfRjPTzIMBZshjuVHM0nk3IIX+AoWDpNWNd
0OrABab3nzBIiD2c0ImBqUb8VPHoJVOhfnewYltnkAwurAM73GJOzj1/G7Ur
RPRGna5TaGILzq1raS07+d5/lHuj7qrmjCs+NU5XDq96kaxrm4+IpzhggdQc
RX2gTY+3UdO6v2O1ZO6C/hTVzZHylITlDk746DvRbshCPU5sxucYEarKjPED
oyMTBhmMdrDt6YZDDIJ4BIP5jKi61XWYMhhwvdvimeT6QMetqbSXhd3xNFAM
jozH4GGEBQUD80cDEq9GI0MCZkBR3TTofdUmD5ODlgUK+8RC/4KdzKckj+5k
lVHytiz98Drvl0eyYkR/wAmGwsmlah2TM/mq3+2nB1owGg7kdWbxs4OMfbIg
FQjog5ATv+yT4d/9jMLG20kImvKgm1LZAhTAo4mC/rXg20UF/E6+T7mw7s2+
a64ximfLFj8s7/6InD391Rk88zR6QXHTr7siqmDGegPQ1wQD4r2vcMjDZzct
oKiDjrBuTQUhOTftOHnoZqNJVMhVJLlqmubX7ZhlY9T54BeIRgJs2amnf3tu
bnFjT+GUWwOxR+OaZXKa/JZNi1uLbnsHgENDXX9vt7LCGUBPCIhpwMVRiXzE
ijvoREg1ZNBTrzrD+OJPgm80fBwh8A1ATDLbc9bvmieM+h0UFGcuQ0CzpQ0c
C1IjeB3MlkRyY+B9sxUtBrJaANb8gD8vFxRJ99yFbw/eSm4k0bKC45eiZFCN
U8BVnzfqbUBShnqSmaJ+TOQUUNKb/D+gjXT2Of2+mIQKzvDgGo5CgrP70SqW
xgbS5Zrl8QE7wZsFhJKbLMMTJ4tw7H33D/NdnOUJB+2pVYPjte6odzvkR7e+
/LZf9E6pXJPkvAumpGeT+HAqB6JotNKliQbPSubcXfL/HP7uYCEBO1/XsNzE
g73jnj0zNRYhvXEcFK1h0Wk35qMagSWCdHX58T9q9xBui88e0dRd19R8UKgr
twIkza/sUAxTwbinavplo5dDveYg3Q6BHXDLVOPN+cRZWoZjkIZJLIp7XlN3
dMjUSjMLfAJP/+AbONC2ec/SLYtyaKIfLnX3SNAIjky9z786OPzihB1VBwLh
KpntL38PTUIXkL+ogKKaiYPTg19KPHESv8smAKVD9+eqMNwmBJHdfI3G7dcb
QE2zy9B0eG4a52JkIAYktDoTXBE8UwAEpK5N3u+ZYyEuQuHub4iOu9STAbrv
AdG5Xigt5ezCFXHPbdtr1b0ujEwlMkBk6QwF5smdkEohqPldrAcA89DZ7eu2
N0NCCFgQHGIsP6rMF3FoFoYJ7Sf9wtG09c+kN5xYapkvVX64bok8/k3LWqS7
dL/kLaZ3oyHXubREBpmNifs1JLw7PzwC7y/8Zu/eTOTMqOygRrrBa1KfxdHF
YgnAr7VaZf+hNRFL4EjABQjRHlGh0hc9f8J48cV00A2DO9Y/YFtHRbWYtYm0
eUv9Yt3ELZ1SQ2ygcFTnECv6WC30QeoPtXJPyRMhRnaPmj11ljmAMTpHDxi8
gvosIJSilbXKfu57nAn9o3IMjvYBRTz9Poh9/rmokY37ysLm966aQZ/Pp4BK
2c7vB78BABw75OnHuyIW//XA0wnGEF6I79lCdFXtoXsvAp3BcYG4WX63l0ru
XhKbkhOfVj3GHTtFbhojV2UJc6R8dtq3tmSZxWfG/mkSi7nR2etrq9ewvK50
cgbMVuHM7soWQm0qcJBHNjTon2OfawMubHaBbIgbaM83E6lF1UMShN9aN3iF
pz5cwPIA54cDe73Iha4jVI9RHVAJNBlYndgvtKQsg7Na/Gw/z1nb7/LUDHnX
8hnospmRZ4iGnvTGnk/iBEZGqU4odzgNM2/hySDL7PlctD4pz/qQFzf9UquA
UtLlhBs+E0QPhAJrsy4rjGLWz546FyTt16twQqGqn576hDJdf+n6mbBYBoRO
KL2B9RJ/mFoYPOf7zcLgrve2IKyLl+qqHFcP48zOuci5ZpLngCkCT1gxDeiE
hnLAxRZRZDVnRS9CC+KNggpsnHQwlMjam77ZEiBCPNvCmcRdekEi3FYb0qUj
9UJh6I7JLGJZMNTCsehZLTChOBA131GsIpy1RnNBG8qs+FMh4jmZkNYfHc+K
fAkRbAneAx/LMlbOZrzp0O4F135pIXt/BQwYnscjUldlDLA8znRF29IBcnPb
xvg6qa+C7jnjWZc8ucHeqzXhg3/6hJKwwnxuLBdhYv3Ws8USebhKcxCemct7
UEtNi16U11F/zlBr8cw8UopkfVidn890A3fKhVLuxuax5npLdeRTy6KoPFiL
Mn0l3Y99X/RcF7tCcKu248QCuKJ4fNnmO7W4gUvRpQetZhdtgIRlV/BJJSq1
hIYq8YrZA9kv3Zxx4QaJtky/XY/ohyFjjsvLJ2OrdD77utpPKMm+tdJoXjCG
HuC91hKEY0RmBMhhwcp+95dGlc4depvwiN7b09wOXienZshjsnEHVd1yxJBN
ddG/oBqtbtzu29dDBzReM0BhfDZAqg8Sk3DNH+G5xZKkt0wq7CMpNLYvgYt/
Kn542U+icOjvWpI2ykdUFCHASWRRI5hNTECBEAsaIXqUqoRkV2MS2a2yYdVx
fWHrhoVGIfSzFJWy/atINdT/2gB3gZ8rsubtsw3GPNNOQHquqVtUT5JE2xLp
DGn5W5eUBjJgGR3Skld5WGJVW4MJe4KRwTG0P6zL0iEDZOitZ8Cn95a3rfzc
hY2eK3SQ01tSzm8eVk1DJnUJntvo2//Z6ZPBbwh1H6M5FVxH1u6V/rc6oR0T
iOemHneg8LjLNG9z9j9vLvbdV66OZ9Hl8xMSzpwn5uiLM4SRBqEWUxN/B8ZE
syOa1JQlZ2H0B0KVy98y4a+5ANwc7sCOtTvbB1ua19XIMIlACGStbsv8rggl
MOKvJ6fo1LcqNI78U+WjSn20rOew3COnWjQWjsnSe7OaWF8/uA0pnXPeCHU1
I0bViCJYKSw8WyDugSwRE0oPUMQUUk5z03FzUiHZKnFMJlWEzSebQIrfnM9x
Jx9wKx1X1bSk5Sx1pz8jBMxchHt6WfZyUAz0N67dvCrm+rMAnOrDM1oK7kyh
vPfj0WXElJTCvaov2Vt0tqZuJO7lAm1IeFKn2KtQ8Eswyww1+N5ZKxjk4L/o
QoWLXcA6yu8XPVpeWK8BMM081qD7Vfc9ddfXqCP8bgdP1rwsdczgdL5+EIzr
OGg6Q2uvp7ghOUqawo2AlrCtpB2vgG7k8exyeDsTo4VRFvqDngFSc/VZZLh8
6R3hiVFd7ZaSEz0tfUCzv/ljhrYvodHDIVHdwi2DKhKOzHMJp9Sy/yRWTi3U
UcCCGb1hey+F5Yw1XzLTrWnH5fNP+HmcCIlcIrcDNL+ERnYbzwlpsE5cWlsr
knQxG5KXMzd54pDzMplU+qKhhdln8qNsE/a35i1Mm0AMfR4hEUp5OVHE5tvc
rNHuGAc6gjOUh2SnclLcTDzGEoc09aLbenj9baOVY/Z3n1GxyOyzzj7Nctwd
qec0CO+paD9wtCCJmFHTlWZsUm2adiFjtBhh6CHa2smMeI++WkokKmQBESTl
hibvaAWwTy6qrJ0a3RKeBWzGlBfqG20Z3JWYuACZysZixYc20wHGq9ux/v95
L3wGd2TvpQD6N0afMS7v0OH62R0npwzyrwgBBGiB8XMuJCUFhonRtzlYzEYV
WLaY2ZP4rTIgRVyGG2bubFWB202GcGK0QJixosPr9WytzwoIfENMdAiJZmmm
X0Os6LhAjP/dcZomohr9kgHQR1jwRgbe2nPfJzz3ApGYpjDgAPItzGTuiWQc
/BaJO2lSSe/KipILZneSA9rjkIUdmVZZ9Mttuq/5BHNwThVJXr7q8y2sLHrK
iGcOWBiV1OlY8qP5ub3yTfurpWb/vcUruRqDqpr/FF5Fjd98SCTVk+Xu6Hid
Ala6POrVGwj1zTrZuSiTAQFEyi4I32HfFWDce7KRs9TYJhuUYUOePU3l57Ln
xWh9lflZXeOl4cw+NKQ3zevXElzoX0x8zdaYKh0LmAaw759Anc6DiBM1XDHa
LzTUK2Wb3tnlo9ZmULwmVlo8zpMmtVe6LdOGvqFUtJClKViEH2DmOqFMRwrF
2egIi6X72DD2xAGyIHuTWhr0/l5oTJWp7MdsOlsVJ7bSemzeLxuGJ5MJAvec
57cT6lbZMbtne7fZCOilu9BZKHsqMVqn05XOEJFfV+Ooli1KNAswg3eQSDkr
u0jzZT4utW1vpeKTDYYjumbGprw6tq95rHplM8OXJ5szJk/PkTwe/+wLcjD9
wetsnSIFho3Gi8JpZBZyEC0O6yn8h3MrNo5CBqnGco2iGjjoa+feEUM3Lsh+
OCoMCq75WmfmqmHZEYoGkEWv8sPRwgFtnRubyIZJHzbu6XAxJ5RyOnzizKEP
5tKcPRtK+kVUS/5subKscQdKAtFeykdSMlIfhCV000DJq1YSqvalGHAnTJ6F
kDGOLAVW05OBEEpyXyq3pZwOrCP6+S2UbAPF1i0kmA8M2tSYRa7CKheI6Rim
vboG0F9K2IEghYoU2BJRLtMlm0TfPNCktDEI2A5DKqChdGnHBKBrRJ+cLaTG
dwgpkhEYsQuti0noy4WW+l/9Ko1NVdSCEE+URJiIcNxk2F3xaH6wKjZ0B8J8
EC6l6Y0XdZVqS9tIH38CH7hogzxFvJgvJl5I+YeZSEL7HwauA+CUqy2Nj7Xl
e4h5BaxdNfpRZ7k9OX7oxg+2ufzK6vBYtV0ZJsIcuXe+nDghIHKs7ScUs98r
xFfTQqtsQnFNMQmvLWm0pz41gzpPLoGmztrFTGXwu/jaQh2ZnKnrKg1/Kcvh
OSgj4ytVGzLGSVM5QLzY/bYQZ8GOeQUnYrtQRwVIgRVc8XYxl1Ix+jdvu7nE
r86ii5c03bWeyPqGXlWH7j1LluM1liIzn3gQX98APuEBax3a1nQUoY3YzfDu
0ilQr9bfhLviRAXvayd2nvWQAoGlLXve97/XfkixFlnod8gTzkpDeW4R7tCt
+yXaEp51iXRxeZaIUFf07qDUTjpyaM1eXVIUFmxn+Acfb3wPySzbpmIW+fhI
/dL7BRN171htJfF2poRoAtlFYXqOoohvkX6DutUHzGXUECMpS0oH5781Swt0
gDL9FBwVtU0aq9+HLo4iNn8GHnfWIX6/28aHbQHHO/iSTQg7pMBkbhV1I2Vj
dX8fSR4rhvYlop+72PzrTM7j0MoesvrtnImA5Q/LzT7PQ5LQIf4VfFT2X+EW
NEuz37c9re75C9/TBMtINyTlyifB5v5CXBtR7zKJ1PLEKroNescymPLW3OZZ
Eu9EJzqxXOCpxqCLoPrTDiyLhxPGUHnXzHMKxBWYW4xum3PTuhBYskTgBbrt
FOir+dvdxa9INI3l+W9LZUSoAFuFf4TOxkvxUSrXz8dYh0MVFW4KP5hgiyrS
V3iDQocvrsXGUECK0lvZHt5xvLxGZ7KBlSXJcMYwBMBXBAYbpNHcx72u0Hda
B1eOpZTdlRnpgWrS1/MsZZqQmFlNlZbsZff7CmOAcTXOUrUDaRUzzsvmxVnY
2YzZbBfAdQ2jGL9JktB+WutVFXVA48kdQWqEF4Sk75+bFycZ6gFfDAq+XUEt
EvDAlTzLco6wxSpUdbfedtpdNjIHh4cniakfbd0jZ55HbJmHf/XEIpWsyJxf
WgAESMgekWJhqY3qYzcZUuaocyJ1oXZflpjOOt9w+X64bqxzgaimxNbmA7Ay
FsYPallcR9vBz5QOxnopxUMmBCLoT7Qs8RR6jEGZAmOlmdbzVLfkQ/1pSLOe
vnfvssOLnDzKSOKYP7uA2FGA3qlxG8svaXhF5RYvn9TMzGwdemnqWNOmPoK5
g+yHRzDax6pJekn8RdnqiIqKDTYXMZq4cKXzETjcyNcgTqXJHuuLi6h7rpyD
2eVks8Ww78l6w5o9T0N+jSB6sqxX5VV7Xcn3yzc5pvtzlhuvszRO3BVZFaQ3
n9nsPkM4LT41MzioO8vu3RgXkMXTwgL7+J9c38PqdyBzJryrA3E5KM/chfCb
xCeTFOrTJJHMBiX3RkQluyPKMCED+uM3rKDa2F6UgJkvxhvvqQ1qQe1Z5Oxd
XE/BoyT1B9gtLrzqKGRBmnhJJOQ7V3Fy6atuCnGk8/yZHZFGje1qWdNEXjIo
LjBeFyNotkdRk2i82YSfx2eOemocrPs7ZINzcEZfr4Z0W/4THSp1blGGxauW
x7YyBUBUHzmgklmQaV1v9O4ehx9HvCnpE9fiIcoTTKIK0KI1S+DxRIYU482L
WF8Z8ie2V92Dwv4g3+zf76E3dX532309nD3NdQSE7rvWsHWyUhS1qXx/cl3J
N32Xg2A5faTXUACNLQ7SR3n0QzLyTcGYvdP3htX6bhlQaxWaYNkpWoih5L1H
hZqBlJGIApy9fby4eWAuzSvMxL5fQEjtHqhy19LBqA5X1QAdDvVIvgkXupKm
dCdFIvF+iCK9mokk1NLdJ4qUbdxnDh/0nkGevW2QSz3zeOOd2xakE/JKxhsw
8aMIIBrE2oDaoq4J9bmcZelbyLPuRDUhtZxZcyasDWmg6bIj5QHhhG6pRweW
AOthX7PQfUKRrA2DvCZcOWwcQKvSMJTI4pH64wFC9r9kXqJrjKgT+EjnlSH+
mPancVY2mbndypgMnvt3GAdg5zbHiT+w9TU4BzUr7kXAsfkw9fDWB2dOFs4V
AIYAZtDWksXwmrzGhEyypsyHSA0j4+xoHuTEuvxgvOvRtaxpxENkX7UkyGwg
Zw0fDV6I4fnkJhSei3voXKJUuH6Q6a37gTF139RgSYHsnatg9eWyFlnnmeyR
yeHKl4lR/kGawVAX30GVtaspB/x7oRb4ShhgrV0yayHnObxXQmlwrmB8F+rQ
egPXWnu/qZJ9rixz9bnHVuXCsiZBRSoB1mdhigv2azSqw/mowNZ1ntUTjsNL
NHqhEIIy+mydoEIygH5+V68/3RnCRhnBZv/Mb9srSW0lDIXfZzFOXeXkVlbS
hCsGSPM4gr7jkBtXF3hYdiRDDI7uCYOIZUsnumB+L3XqffvaUZwHfiMAZdKH
5jWlfp9ZcwomncfKGhfAFoNwV6dXiqBDXsxWAljhh20/k7zWROFHHmQ0t0Jr
peM8CeP9Gl7ldoYNrcM3FU9KtYWLXOfeltsSIykq5ek0QRm12I1g9iJyWKQP
KD2PCKzjPhVGOh/bvZ7UgFdxiNNQcLoIjzEGdaD/a7LAjakh/D8x7923/b1r
k46GoXmAVcN+rtEHcGKRmwZX/ZrKM6Oa1YZY6VK3h4c2jjJyiHNhuvr2eHHh
Vz23TrO12qOA8SsR+s75P0iRx+Ws7I2lJq1Vjs3X1OggJ7tRvvftcJ7gxdrt
cs9kTVWT+dlG0p5bmuyDaaBejXY9yfmnbI5iey77RAJxsUd7Jtov5svQ9NbS
pNfzzrP/Q0HAZK1LPn6COTVbAAVjc8BEn8oAwWNpaLACuY5PsZw8iZJpD6fC
uq3Sgr68nMEo9KN7CDvjqtHJLJowkTUvqb8pCSRhi3fjtrjJeK3G1qQWGkfW
2FNpXHP0cIGuaDvm5VJSYVJXMJCww3YmUgu+ZgoAtHE2EzEdIo+Fjz0dGNWg
IJ70Gi3yczO26Q7+MH7FPOU57/4NG/ysD7X0xT4CUD74Sgdk0DrRn0BLCUMU
GQOvpl5IG4Grpju4ZPQioQV6bdMdy7ygbAi0IgmjvpeEPApSsySo94CBoRfn
vKTuIKsi1cFDgnGKdzvnpdFR71HWuOhj0pWjtIDTkwKwvMfUgVpZBx1IdAKh
w7qkuwg599JMItv2yDCDv/R2OYhwi/GOJgZ4JATlc7Nnaj7R1f7NQKZ0xpQb
J5SDIJsbVVi7xKtJP7FqLdp9q3Urq8BqYDFzC7QW+qrMbG867ififKJOPtJf
WCfGVYRWRfk1Qy0RDhE+DoG2DAJiClsSFptaQ+pbDGRZ8vaHTG9FcEeoRqvF
Ozb6jnEO+OGR4+QyAtzq5EX4GuIh3Edato8zufgNM05VPvtC1z3pxyKUJM8O
afSgunBs7jW8QZ+1L1bJpG1i7bSaRC4lOoomhCGDfHUoceyiQZxQDclwhvfl
rsoxAQyqVwUQGeG6EVLlgBI8S/lrlturgv+Y7qcax0o1WYCotp8/6BLghxW8
7iQkrIEI6dg84OSGfXtAYeCtD2WkrQ34O5Z3iOHZX4pdgPbcZ3WkkkcWVGpn
8jKcXRQbQ1RwFiXHx7U2YJ0TvtW+T242sjTMoZMXKDQxb4/3+RpHAir77Boj
wUVzcEqJyey5drxeur+SwZ6u8YEUqqFIo9laWaDrQNrXWnZiFDR8hCqlwjIy
PQFIbIeMpPjwtVbQ87HNMjrycf8orASIt2KmH/xC1P+KeiOWfYkOLSV2YOou
cJEKljuucXhyqE0QCtjqeVReSH8+n1tc0Yi+x1Ql+8Jv3SF8dgOMkpndGWiK
en1RBDp6pVQpyiHj/WJpnWMAj6IFdXrvLSRN6HMipySzCSayyETfVPpDHXpa
H2KUCY56tAWztbouwGCT6NRfAFwX6JEQkBkuBOI3C8YiBdNA9o+55y/kjZfs
Bp0sThkQtDpCB9Cb6eV4O9uEHqgx3VgeCpPra6txo3lTND5KQg8yN/1kja+W
wKhqPSdR3+URO8CEMfubK5Q/Ua714T6e7dUxTBjmlEpcHRRL0Y/jYQicm9w3
Jlg9NsYRQVvYalVP1btaTF/MfeYT3SuvpgpNTOjEMoEcEwjyzqS/qcheZiLX
3+N1vw886e0rxzxnlwD9ozi1fWhV3/pUlQ/LLJroa76fny62V1BQ1wq6dU5u
ePWrGzzuVDIK6eYHm3GmCteEyNbtndQREp6Vg1V1l4B0nHVGfxh2uwtEavf/
vQHNAZcmjUBuTo0vmChnbiSu16xETtokKEulkheFTXut9mDjQS8zwv1smR5h
Z5pskX0BE5S6fTExgS9eS3kv/FKIqs2qlk6ebvJpMVwWdWkHGiS7XIl8CSGL
Fkvvuiw4PPFtxHRDAOXgbvKkEHnfw9IUHp1rmXXxSpYgidGQcifX8JI4ON+H
L3w0yFu1m0rs99rXB+jrp3Zn5ImmKyW0tDpMcMcQbC7ITg4RTFykZTwh2PSJ
rEs9Uuuv63zeq/guLq8E9saSnuUfEVB+94RoihAIuqsb5FjdAAKFIuSjl/dj
oMmENDRWpdAN1W4NFmlIjwHb48JDO4nS5huyVOVHil/jAcsBugHpBr0jxa4L
kqWr73IAmiUpO5I0fWS2RZokdPSSFjF8nXTXv/V6bpg0DxLasMX0a7N3eECy
J7d09nzoLzsRPUF8OA25NzBxgwkN9/Zw0HDW0in3yNaDdPfVtWfrhwAHJhYI
+4PZauvon5Hl1VhOD4WvgRBpWmN+xLubC7UjXzNzuIOE/tcJa811g9ekPC80
G85mVY9U+qzVIADmcRmnvsClqKIdN433RPG7OCBHHzhyXYI4d6fOeKw8mh5i
hu8Ev0QgIe/EirnR0UTQfbkgNUsax4FefHvOmOA0xl4HgIjVOu+BzimOGh4W
gVoPSWouWAknwY6JX9L3bzP/qsEQz190JtYiD4lexRtzyR3sUf7hhepyAwVT
ttxKJ+y5tnkuPj+PzyrIM1OHwq+LD8z1FmWT2bd2Funi3Pdog57haC74WYq6
wF+KGKKTxC1TnjaqvKPuE2RlZyo6LSo0cSfOWk7YPAte87QmxLloHQh93jyg
/kg090dMHXSzR+k2xvWU9n7jw8g8Y/Ba0aTNmeihqG+5mhDCjoTpiJEYOH2p
YzxLc5deGWdusUq7l8LEqg7HXWSBcB2C5TTAQApD+Awh+WkNuGtT6RGPsDQn
Usj0ERi5qFPGKy51VzSgJaOYylLJ6g5aziJITAO5Qli6BVC0EaxUxb/e9/Hm
KKeLhf3+zyRNw/hXwJ7XH7CmZDnnadt4cpdDc/nMCcVq5SrX4VpfKWGNElGX
2vLPbWi/ksJW523MTjDdNBkTekDRss5iDiW9XnBLS/0N24ccGqKdMdyGu7Fk
3i7bMlA/5guXiGDLvgzM9iJ9rrD94T2k8AWMSQ8RFxJYN+t3v8ml6LVCw0d9
78y7WWkBNZqzHfWVGDPfdw0UIp/neJomvo0fDlALRKxP0hskwdapi3ZE26/2
Xbvnjvcp5HWaSCM84nwbcqhocIsZHJYeu8s8v7jktBj3s4nmX33ZxX7luVfI
l8zLCtzsNcXHnTtaujzelLgzRhf7vfWhPLL/tcO9hDmlnj+/Plnj5I+56ogl
iqt89TH2+YxhsObvu5UMzVEvUz4afGnhMpi53BAgK8SwYVOswwDM2rEd2odG
ZREhVgvjo3D6SzMXaIGXOmLpfAiFc/rQ0M1IJ4h/KaVpIbvYUFT0r0s3Z6Mf
GY9MHNQcxB0DO3WRYqAY9zjtudJejyieb7o7RH2M/wOcVvHO4nFF3coUmR7R
1kEbn0hetLCxuv39dDSjIWPFp1RGdZ5JGybIHOvZ/7tVdtKLD/eFsb8kUAsK
ZrBXS1uDXFVSzO8AWgc0s1G2z4XXCSjbLQJSRlgYSEMQYMhWOHAjQSisqi4l
bZShck9LJ4rkFf6w3w3i6fyOP7gKdNw32qO/xq6cK0cmQbMXKkz1mseA0p2R
K5HyxNrgRmb/rhZqzzT1knLmDaEevonHOKR87mNdpIWsSIWvID6Dy4V/xewq
sp5nnIpjZ1WLFuzPAm7OhiDJh997LKtggmq/7YCjsMWfutFb9YIX7UP7O9/V
cGobqQu0/T6OTKxdYlrGYzINoQ9Tr4fT/HNWxa3/KCOR59su4kV3EI+ISAuH
AkH505EMmBw2m4r8PPvwqKWiBw+2yMR/pEjBF/h39pPhEaOyn/yh0X7Lp/Xz
ry3yp+1KKRwewoFqw7nYfR2or8ljd9ePDKZYYqKhS4K+1pTMQ2WtlGuPGgao
tNUWsjgsD9mOLE8n1I9JKuZPQopB5N+T7cIPuBQaNJRIjJPrX3j3OfVnqxZY
jvgg5HpHc8qI6tsnP3p+4GNK2jihjh8ZcHEPjEE9jJ58enGt2Ol2MtOvwXAG
8KyNU/FxDJhLPA2T7h9Q5d8aOjErXhhGTYgtajUuVgZPj7AgvSp88axmRwdL
vpsX/3xOv1eNmnYiszQl1Atagm9SYrBp9Jx6stwtOyQ8+9RyMvVnXCrFd/xm
Y7Y/oNs9rVHMpv0ApIzuYRZHDP1jBefcpejgAC1eYKQ1A4Q3i/D0LaKiaDlu
c13RyKbfm0gc80vGRlEoZI+RKnIHj5Yi75IbVxpex+sB/SYylx7c4aa8y2rN
lszPJKbapvZ8hP6vBPLfIK+XF+pIkMl0MH6InKljZXUjqoLxS5xtKFRK17l0
VEcDsRsytuO5KEaM+RTw+TX/za+bZCs2UWI1oD3gHJbgrh36wY63zwSGV85C
215ivVz2/omulGqrWSTd9KaGXFlEPd8u0G4hzP0+Uj1RITzAd2Cuhsi32KHP
5dlbvuX0y3DxEWYTwAxgVbuHwxESNgFtSpbseQXRLh19G6WmfaXtocdcHpHH
QLlCkB4U82CIY/b7NgD/dF+h1DhR4KcW4wz4+Y8E6EXLrMMiB4+JiCoPGQ05
67cugAl4uoLENR5xx0m6xUZedKcwaIQMFJq3+UsiAY6Gph/427Q1J3zddxKo
3SJ8My3xJzjHnFGessBBxjCvsulXatyrI+FHGwlDXhmTf/2TAsGeVqIZJcK6
c72xo5UxJSSfTFbvRCvpkwGVsoHMuKc0r4kq+D3NbmjXCAWCnZG7LVjrTRtk
CylWIm+/8lkx1vrjOBfKjpAcuEL2qYWPUA4b5IC+GhGC8iwAuUdjA994Nd9z
audP4LAOWpPniZtCDrCn6wAf3dqyjYZDtTfPO6SjhI0EsNTVxkl2hIKMD7DO
A2JGFk0mLuHlnONYcNxYt96NMqmuQU7lEp+K7wqK1lH02SM5mqHk7Xrjw5nh
ex8n8/GkMNrFEQLshaR9NCeTVwWgl8eUKz1ecbB15sRaD7fDCKb9f09tWEju
6sMZldC5HdfUsZTAs+KDBPDNaxmPT+3z81X8BLfNlN0lFWj/vZLQoIjlsNw4
fA/JjRQU3CsrvpGbXInULPu3YGBza9GaxpPrLBrliSd0mKcv4A3N1J9ZVbJ5
dUyqwlXJ78V1zssZVGcJprCLMmxSvmxj3soKEpKKdx8FLbhtnoomp7LM21DC
8TPfAvNC/t2ffTwNyMwKpLtkMuaK/rmxM/3GprEwK/JOIkNgqPMKz0Hz1O+a
jrZBzGzvWNNpYE3+bAurskKGxFQxtLfbIG+uAV3+oYBJPnMIw+LjcrPCTLY+
NvUGKxfIMLZtLIn5u9PjnO6lSg+qNd/HHjkmesaGLkvfTHWi1adYG1mvwvYs
1nTrksAursyJsbCAFIZRA1gbLFkdeUAHApMKDV74je6H7SL3lcTnSXFMXRol
AACBSD1WWv/Z3oPqN2EhPaLHE3bsafOA9jJAnwbzBcbjNgSQ4MlVOJ8gcu51
O8w8Vf+U6qtLvpKwkuGOOYG/vg1ajPKQ1tkRxukXHlVJljBM7h1jQWGX0CZP
KNHqATcOTZj1q5kOfyDiM3QMNjH9su76EnMP6b9csGeAR8mzc3urM8GLo0TZ
VdijWWwNsjpu5IV01P7UZ4sLe1V1aXdgE3FActiYiOaNmKZYe4vXqMHyW2Wi
geqAG7vEMm61N+T1t4UIihM17co9eb1RAUYUPv5DKFKkGI3oH7SFcwqa4JV2
oy1DtRACBDSnQ8ptBZ2aJz/PrpkKoVENxhmBJitHcVuG1/rdVasYeZXtDlNr
tYUA3F/nlQ6CgoN7onPd6GY6VePe5uAHRW9vYw4pLZOvb20d0t9w7D+yjaKW
PS3MFhhx1N8d54CuS1QUgOyV+JnmpOfGZXLwagBQzPlKfttaHDZrAkr5pR2K
FL/1F5gbaTfpyx0LR3gRU4RuzgD8DhxS4IZ+RCQ2L7hyetjdExqJjvv+n6nC
kZJTgsOAOqmgFoJQ07P6O3nxaGGK7dLUyoO1V6XQZv/XfSUDzXMXoZZF+1RE
bu2bgeurKvaMVPHr3J3FBfpcwk0IC26bDepjWA9Aat84Zxv7Tk12HQffli19
azX2yEM8znCBkodHcZHVvdBne5k6llse/sl5s8jNBBhr0vUaE2J4ay/Ae+iR
J5tkw3dT0IilzCjqtrgpfIJOznYXPcQS8uEWMtEF0R1WDHzS96SRoneNrXqL
n6MDv4Lf/RWGEJ2HjravoS76vxTXX/7bAG001OftMLNTxZg8L+CndLzUmZYx
vFqvGxRTnMuwbBmDqbcTHkDf7ryQvyJfS3oe2Rl3XgK4FDfiFYi8UsYkqAev
8LeYQi+M+2roBmyul0dLs7aTnYqZbl69aPgQ+QVcP9jgTT9/+gPkGGCVWmk2
9sHSfBsYtoKWpn6kconW/1UORYXNaV+DA6BL6H/KCX1Bs1oFrIkd65bTts79
N6oS34P+1mkIOVMMvH274K3TifvrFPtGGrrGGUbWXXoLF0sIvMNobS1M9gvF
bNEmUEvsAETjhqKSbn3DN0J0a9Fgs9rp0wlCpZWYbIujUxWkmhraKCJ+8k+p
X1foqU1mdoCOBi8wF9m4PYG9oMSJ8+DYb+99KxGi3TLH1HAOM3OmqoxA+D88
FN9YfsXZ0jI7V1r0uRHfcQHvfuql7B2e/5RtchKWLdqiWbNA9aVptuZGUsgz
zXF00R02huVLVFzMBOQmc1atihBgNNROZphxoCsArChUn2yvBgh2kOyI2kDi
7a06n+BA6qO9qbc7CwyOcd+jIlmSKCWyCDOJ8MnaCRD4Wv71T2ELd4NyMpYA
05DO47CQu44JifSm392Eemp44zNTmT6Gt/UcKDQvBgz91P/Mi/7rORQia6ah
uFitIr0jv872u0HrM6Qipc3PXw6CwhOnLP57yEGCyd5j96tDTlTNq/Ls7U5g
0TSArbljoUtD98Xl9dQWifrlZF1o3BvCVNRx701IXCdQAOX+KYkEDK+5LNT8
fGjdkMEgE3DUWu6xF0Sox6jl8jQmNVA2Kl4LMd0H7XQqsHr6vIcSCj1M0FUr
CHT5ZwjUcMdcswcBLItvT2GO6SPWLK1Rg5/GZzs1sRxRRGWDi/tXB9RZeSCs
vUzBoTixV4PAkZ3Ntl8vLt4bGGiOEecKBSXxrn1n0Dw9BftEtl+9BM07ru+S
NQZm+2/QzfuxiW8UYjovbhes4hHSEG54Lpmfa4lbwIaUvApMvKrY/qyPF2n3
CyCj2Epen7opKcPJfx0jDL9+D7Bqzcc/w3yW91ubp1tdSQOadsDVDzd1ljN0
JY4VMFXSAoSB4owCIRGladO1NVJcpLBxHHv9whNd2F8t/d/oQ+vWaoVM6xwU
hOtrMOTl2N9Pro4wbX3+Wuqfau7ZEkLxjTybd+7weMeBSjMxNF5o1ZPmp2hZ
tyygr933ib4JqlFkZmWSQ2wtlLcfBeSe0pFziUqgM0Qr4t9hatK5WHf7zqBS
KK4j1lW7+dhsDPlw6HEOJd2Rf8yaWdHmH7OZj/IHWiUBwPyfihit2MHlTQJq
RRfPn8MrjeHwac1Tv++sGNnO0DLTCQBMhzWZe0vpIam13zli3y0PLPapIOQc
dZJIkfbxI+IpHmxjzFtHBidQ1+gyVAoigUhewCedD6kKK8mIlNp7T8sfAWJm
R9IjZ8B84Vk2nSRcRfx1YqR4U3Sf7Uu1c/V6bqufkdYA/HfFpKM/as6w36xt
RwIDxY+eI7PtVpYMiSn55udd5n6m79hYswsYDW7sVuQxL4XInnw3IodVvdxj
goizBqq9u1Z8RNUFKLmuiJMJGDplwrGUERMIJmt5TxpPf2SVIUmagNP/YjWe
Wo4zZ5YFGER6hhHKgIkmyulHeatM2AUrGL/vIJGqWEk1XVsQkqqvYcLLrsew
Qrv+EdZwvNP4QKuEsTgeufHpdz299Y80+6WvvgERjRl+ybCYhgazIbiN9e98
OOd3z0ZZ+Kpm1xbuhCAodpB32jV/4KgUsjeIcZE+3bOOKEshD3SjcfuqYsHd
gp5oroHIuL1Q+TEwJfJfLuaSeho/hMzubEZISawCAQOvzy35DSA1vS7SfFP6
Mj5IMKj6tOB+JHx13SkDq3HDkNGL5UpSJ2Uwn7UFYodcvrw/7B3Km29rUf8Q
ZI+x/ISLXPiShmL7ZhHJoIIM2vlXTHEQ6audJTtvh+8wKq6FvrHlesEl6m8V
gMsS2ph1LI6aVpjIBtncz9gsKeUXAkg0bWvNmHAeVz6jvoB4xiQRpA0QGCHD
7Fl1eO3Dfu05co71l9u4aQMmZciAJYQRrnR9DA3Q70BsE63RGsXjL0p5Oc6O
FBKJySLTbRKBx2u8GKpIMQyM4x7wH1rP8cjiJz6dtEMR36m1juX4HaSeIF2o
4jus0rXMqhZyXpeZvMbaGKkMbDWvvf6j4DuRLLHrL8hwf0gw5gXRS8Q2yRa/
IctqA2n+Fjy7jJ9jUcRT6PVSNbhQEG2VJ4YvMM5+Hn1wJkw7yW/O30L/T74O
etu+fR4NTjLY1MyhciYc6v+Q8LjEkAZuvq4gvy7FT1ObH191yhutSLuMUM7N
kheECnzDMbfru6k+jzhI7Vi4Mw7izs14Fx/r6lkpEmg+7Jh87i5NP1x7U/mq
CGhjL8uzwzrm/RptOGR4w5RAplKK5lthhOPMqQT32H2Xp+zUyeN2/GyGbPVO
d42AuMTS6RFIKSP1qnuM9OTGEJAc1k+toNNykUOb2Y/r16KqiTZTTCRrDb1N
ER+5fILG1gVipSG/i+TeNztb2tzHis1l17TSBvFPzq6Bx2nrz+a5dMZTlvEG
Q57V4WPjzsuf5a22PNQ2wtvhz0/DRRFZbJ9zLLjSz4A7OyiIQzw/x04eCWQt
GnKCfDA8cIq1wnF4mkXsfELaKw1x97+OkIB95flkz5rP5kVtQwUQkr3NUWBV
kD3HFu5xALYdkR4faEHCWRN2jZ3PWu9wQD/ZA515i1FFWtb8KhEFALYcSj0h
R6ICoxr7o/4mAXvzWMXc2UL5wACUQtdzOE4stNl9lzsuSwTzK1eljK8ZsqJN
k25hQhjGRzKTu5xiICZ9k9Hild/SQn8EQMse9RmbHD14UeJlvniqrvkbnsku
Rl4x4ZzZTdHJfm8iC6gmmWPPfk3F2uOaFZa1yziYMewNZqoCGZfLjGZ3VwDO
Pg0J/TQGL0Pp3zNxHRJey8Fys2DTuEAd8F4g1WNFD+yIx55Z2kmS0VP0e6Mz
Tz9prUiHoEV68J118XAArm9LAzmdMgTD5EZro0SQ3rKvbxsNZuhicuM8geof
HC9U53uQ7Y4VrJBYJ9RD0p72o0Yp6wOPQntvmSLFGtcr7BB5FogodoCkgSSl
cRdXG/G1E0Nj5Mu98WpCjkTBfcuAAGBBkA9dhU9w9WQ5+gwPdFwRv7Cva4O3
KIi4zSRmgQqj+FfTLSJq7LseckLAUCUSFleBxpEuVvl4muL2qbVcWRtDShq3
huPiamz4gqH7/6dHaQZllY2P0CG0pD5BzMt3V5pLCFARmCFaMCfYaY/2TTc3
MQconCWwSOHQ0We0Fq3rNSsS3kdtRZcCL+qqPRzHFjrZp6rzdn26dxX1zgdV
5HmE3uFAiEzQxQznfpfCgy/IhQSjYFOqVcodYwQKr9BAdvS83kB05AzZ/mQp
SfEKOoKv8tR0luykomdCMyaqqjQ12ebgjQELOQUCrp5FCE5rC8CI30U7OlF0
PZE0d2DT0BQlbhjPLPFEpp8BvC76ONCEKcS8N07n/OxMu7S8HvMlA2F8HVdT
3o/gPILL83TzSVPKWgO1QtgAjJJxNrHO/5al1CUtifGQuUI1vbjtFNrdvjMz
ww+nLzH+nDoIrVkhHpaj1rbBTryBAW5yR4cT/h/7h5RsavfKmF+avGru15Ep
eFVOmsEjZUn+0Qthx85WmcgSboc5+pCWYMgaiwT9P6dnKcS4etOa6NQMuayw
vE//ZAGFRGdPfl6FSnp3H+fU2+WPo6Lo+BOVV3R5Xc/QvGikvxb99BSm3epI
FNBZ7ws+X/hmYKU1xi5eAetxRm96/N9aWOqtb3/d38nI6RM9t5Iz8LQSPdT2
Lyikjkv2yXtEIiCtZ9rnP1tA3/49RfFFZ7Jn2aVErpAgguo7O2m8eSQ2uXoL
9f3hkDPRBsGRUxG0ILKeMJ8SuHHy89FXC1Q/aYcxY0ewLq1Kr5bKwW5HXMkL
NOE8oSYvB9cY+kROdWmeMpn8pzhBPpRSNxazI7qxQZnLyM0Dl876HXEqr27a
Oz9fzB8So7FCENhQnxDNJLrTDqpCuS4f19xQGu1QMd2uBONv5JOOHzW3itXW
ZnI94vdxxILDb9WJhSYMnCB9po4rbmQpGh+BvGSa2nzvvErctJWIQNEvPHcV
dYOc35QlKwVRjk43bJuDlWo+wFbEkgzm+xZmB7gD83AZjQ3dOGRV8xcNAmQ8
wPVBEm/e0HvYju30V5U6Ae34sy2p1pcnQ7WYUMn0AAKcKGvnwTl1aom6Reds
UIPW20G2IaaT5kgUjSs75F9aMuNl0aJyJoQjyTDkDjjlHXfpht6BHrYeQzNb
gOdB3KLuZxDrKRlwOp/EN93xxgQn36HDFBk3o1EjPye4BmQ5jWjfzBRPqcvQ
Y+vUvuW3EK00kkCkTEKwDCVceyABrFSgOAdwU9eA5MjhGIk5JtKqkHGZPhR+
dDGI4G2aAGRWVYoTPdhfZq8eALWbu8vlEyqSseCE6K2PDYYFQHlFEeJtlWL1
Xffhd3OiIclov4wjhuWoo4cAWBtEdA1wYvfkSx1PviKA+Yg+dtdXKsQCbsOk
3e5HbRWY6+bosaLd/PotgdKcz539MPZa73iXIYMZGXFSwkrcsdhJcy6LzmIS
GAUDZwQujuHc03H9pU8/vjlZ1qof6T4mKINlyV7KutjQnJNYZt617SxHn8mN
DxSfj/S7xyiMSbXNkViEVHc4cygZIHNPqDHeyOjiYIb33egqX9Nx1mXc5CEc
q7Xcn1cNR4WxnoHR8Atw+mYEkUt0/6AtMjeyjpHpult9G86OE9iEgKqqYLBL
FMV0UU4OasKJHynqaCCnP3tLgjcIzweVAlTD8EydC2yLDQMX904eoyIL95zj
hjNtlHia8tDl4Yze6jotke04kJYSql8CY2zbQtHu2XplJbdlErviDMr4Ti57
bma5EUMlTMkTT5qkdjMh84j8IFBnvRPW7dOus5Mu1dSY4OqC3PNhTq9wpuwr
6Dk8uO+Xavg/YrafT8vw+i0TLYyjV5A9SkCKe749iOOud0AFCyIVfNb6YeNX
czR+3FwpL0yTiOKBl5iWaqDS/rddTzkwQNadX1eIzbL7PNn4btAkxkSYLQLy
oe/KPMwzXyyqeHVjJV013AWGwPWfz0Nt2ENXg2cYg2djCK4eXwemux0Cn5M0
tmY9otaFtIvCVZvPt23HCpqY0ttWc1fQQSz6t0L6X9bMq2NWFDPjlVqOnWd0
xFyXwBVW11s0LRfOjlmXcGSBKNu0yfnO1oGQOaRhi39YXSYMTWFaO2f+sT8b
KhVcQo0YS3XRJfbMz+Y3N6I9w9lnsDWyAMnUVnzrY+XZVFFaL9RBXIb2OoaU
VwYr3sUW3KRFLcTRmyaWQcVckc2dSt9QxDxE/18SyZ6TsJYtTQYs5dg9W7vV
5K7bJiOULZQWoqCEMX3NnN0ECrSf8APTV/ZlFFsHKYEbQ9uxEuOeq//FPl/5
WFmssnSjYV/zdZCqwSVdoqQ15T7oFuKwNHL4Jgas+LMTSzvnNQxdeuO2+oc4
sHh4AhpXWVEFdRid7OO2RwKeg1YrFkKKjUNxNhWPsOFzONAT93j7DZZCaTyn
4dhwlEnYBBRc0KGlYwcISG/b1PctnbE9/zVCDgFAUV15DX0DvxiVoekp9pvd
ZcAVoZOobXhoYhdLuYj4FX0xpKC6E4OHecSZOAeORPfNqDWmlE1BzLdoWclr
ffIyLJbzl9vQuO5ExVZaKbodR7qtR+bYCR2E/WVdgwqRQc44RXqQVkvir95H
odF0D0aGi8T1t6EtMaVatodXqH3bD/sF5wai/ADmi6dgVF/BCGDCXwRYoeBV
APEOihX2gUP7LbJX0MB5ceIg6vlV9a0g2lfk3TZIP+FR55b1PyPRcCA2dFHA
6rC1iZi5OWSMb1tAQ2Pqds0wnHu4YvH1qysBF5x8rz19xh2/UOt9uM/z3TR1
mmuf+db59ao50WZYhRB7E1Ir160/z/Wc1AGV6e+JRNlcZmKBcVY4ZvqKJWbj
XMd0a7U9tODsliMxhX3W9SIfSgDUW7S1cfQMcIcHrwb6EhXtWtZvzQ2XfNLZ
2JX+ECQCTlTRotMLG2HIx7CvoCGumvcirhI50OLGME/Vvv8aVzTjYCbbqMGG
2VsWGHSteTxIRN6qNspNSL238Ia4GfmRfs3Df0WO3aUSOtE2EhqypfEracmy
ftV9XHF3V+He78XkYTjrnYIbQPt7nm7F72wJpsVYzDOBAay7n4fj09cs6Qng
IHkE9bE41UD1nUBe9W4p1IE5GUpmX2cMa4aU6k0sHhdacGa9a5dTXbylbaQV
yw3pDfsLgJo2WCzu3+GpjfcqtdBBfzpjZE1h9LYcztoOgXQKh2vItV6Fibgc
2SKoMODSWi8waD5uL3CcEeHKUvYJIMMwbWNlGJQz+h9GFhsGp5m3S/LyKbgr
QtlpoD3WymOiPlo6HoFxJw4Z8jnVtu8nPfdFxNX144V3yqeadF7YGnJXayw/
4vun82WrYGnEI5+NuHu2nQxmO9gh9ubCZW52mKpqeGcKLw2UWYZJ1PFjXTPf
NEE7TXmZyMx8SBCZvByVQHqK81DE3JKd+zNZXVl0OdN0WoWtK4JY8yFgv6Gi
NW+wGouVm9Lsk8YeXmeJMMEAQaYYcWrf2udAVfNnTkxkqIHtIWduJNQCFzaH
SwVns49aKWfzytoHfxzDY0P9bsTwFXw6VEqXLyWq8jNqxNgC6AgUdgLlIGid
ehA5g5+hWSfVHpDmngTg/BbPf5msi+Nu++DPdsg7n1DeQcEfNc6pXww2+q/v
qH3tXTAMCUp3LNl6ZQFK+pIgmXsYeG2SzMhvy/Y9y8S12XLqcs0YOms96p2J
iagnfGHQ2WA4iTPXDyr5J8mblir93OVTQjGee3DPEwEWMiUh3NXinDmXv7/L
GV1YAP1txIKDw9FvapZNxXoZ4pRJFe7kouUIuhOPR+rwGbYOq/O/AfI8l69A
ISTMazEuntBliusvtdj52XNHqY7GKt38oaiwS84kAhd+DTfymXmO0UT+xtLn
+YAOV/TmGwX66wVTPuyuREsh0fk/mhoDvLuyjPgvGWrbBO3SZe80YDiu4t4c
41zl1MPH7ZeF6DW149dbmUsWB2YRQ6Zcce/++3Gb4qjdLkQ2d+R4kqmXZUk3
WqjWr+BuSZL3VRTwnltofOdKG+ZOPu6PNwe1xXZgLhdK2AKTqynWnPGNUmuT
bEf7d99YZiXSQT+kZUZZRjzoDXBr82VdBIhKs6sA93mCbLveFVs3XKbG07pc
wqfJwYRz7dJbQgLtZQaYoyFQFJUL6V0nowHVhuEI6rmH6Mz5ngcWBEqfdcqN
h6Cmvj6zGm9lrf7Jn9gDNPUUIuD7GqWJT5CEjLxt5ITJAAFP3ImaZpZ12Isr
Yp9JeBDy057ZlXkH6oibPoSfbZ81BZ1df2uLzer52Bl5RvzxR3IyJHhJHb4l
RaPpaKhskAtOTVvrW5Rbe3a4sLsjOLJlNwLAg2+p4ENHt5LjQZDN2UJmUUqq
gAjXHlBJnogXdNKWClgJaFgKsm3O7S8vRq9dFHdpPi2EKwWsQnN/Rn3T2Jcn
rgrCrP0NKirl6IRswfgqL0CebkPoghoCBIcaE2KbrCICVS5vZdwMlwXfvM02
nHqzKhZ3TeZtjfQl4qOL5toCAThTzQgfatuCPoHGbW0SakntONCV6t4EoJYE
gut3txaAFMDqWLSJjd8vBDxj9A/vU5VEnKHGSRNRJSZq6RNEIw8347/dOSph
qxI3qZN8kqtAAFmKajXh94y+7XyFKRGuY77cFn9Ua6rtT6tUozVd7/+Hspar
2mnmmT4XDx8nPiJb6HmKQz0xJFYjjhKZGcqzAp0vrCQRNT0aEQUFWooJ+mDV
8BZXGUzuxNQonE5Tb/5XtDoL5QUNGaJ34jzfrApe84ZaxICSVfZJAnztWUvQ
juoBY82VylBHj6F14UL3zAxXEL6paHXB5zVivU9nGVLEmfChWcymLWLDnbie
gFOvBZSPRma7NrShSa2qqQagdnMBc6vKhBN/8+ubG3/UoGIgEHheEHbGaIFd
xv8DsXasYRfsRPL/PCEw12orsOOJCOlKzh9C77tsAI96hZS+rU0D2GiOwEk4
FkbTKX3l5A6P1QDCwJmKSopLCSIvoI8JGJx2vDRDEFWSK1uRj7luiXYmQLsM
CaSxYwxhxeJv/d2oqLXsqRpvM1Im+PAS9rBtJMRmZD+ZQrXezLTLzfSfFwog
rgp3+T1mtZSoPAwFCtpsi+np9qwFtVpmNV2N4ykVQJcTx6gNFTppZPkvmlO2
ZBrC50wDFT3hXkjSD+/EKHZvb+0Lv7+/3wCQZbeNvvYl23zGy4zig8tYNuX6
ASLdwbx0AQg5lMw56jo2ntQ8JzxVJyiWc/zHZtUc3ouktyCAUfVxWo+uhH/n
79Ev0EMKQLCtpGBs3hVVhCdVBvA8aZxwwds7zr9sGwkJ95xM/qPABBkfb9uf
w9BiB8hWLtEqfXIOhQv8BQH/adR2BzgET/Z9Wjwowycwn4vrmGn38YnAQyMl
MlXFYhealixstANgOeE5p6a8dnApRxPhYAWYNyKLU0k1TFYHuxsW13EAezhm
TZcFAPwElZPgBuc1o/HfB4o+w8W8Vw5c2ht5Ah/8l+7kPGgLdJOivLyWXgo/
S+I6E4wqgWcTcyG2z0JfWnCKa2ZOOdGE//X8y3Lp8uBgsMubqvVgQYatHYPH
Cl4qx/iYhP9CuYfz0slaHYq/SI8ZFIk74ctQX2XkLdzJdTzFeNIdmRhyzRKL
1BXfwEC6Kmx7yFWhcaJxXPHMKdj/5h3F7SLy3ViN45oWdDiL1la0mtNLN6/h
kE/ETvz05UMytQfxTj1lkEZhlP/yTZavL6LACaxxOGPLLGODGyXMQIzwMQEQ
ZqqHWEbuoUNlvcsh8GWYEN3mssXw2/9TSuvcRTc8RroFImL1GZJlXmcVpjxS
uC9SBS7M60DLMlSpS8UCFecSX3PUn7xsaOINYJ9qIa9mJALtiUg2FXvpa9Ck
XpFT1Gm9ssxDJYxVnqb3CgE4md3UAHK67HpQasJCXd0qssER9ezfnp9F6h2T
QUMMq65aJZa5mE5PnXjY7F92AI9ROUTwzKGQg0eIsjxerUAQouzmC5O0jQln
90iVBI9yixkhFVZMfJuONL2SySNB/Oled19eawIuxRaQ/vGN2JbjoJ1/+LWC
ot+t8ctI4BSuWWxqeTxRLl1aZmW4F6idAQaUfZQTF42VzFEln6hM9L1vsI2n
zhaZeLdWlsxMCyVn/sx6HEmPXDzQ2C6rVfGtthjjvSiX6yio7LJqj5MOZBm0
vKC5FGwBe4em7lOqWBfNdiBbD1egNasS0rx8sA9Y3fi0dOnEvwtX88tRVlXf
t+02hJ78LVtBgAITGEJCwdVsOBJ6nKxT8hCG+Er1we8ogMfpW07Kkftf1d5a
6uMgPlbWXzsthyIoWvPTCDPE487j7oMAaCP1hXUqU298UP1JigqGfoKGiaHn
SMXPtEc+7BMaEdOQdOp9MR/9YdttiYUUQSL83/DMLF/OfPMDwKKoNMOCxTu6
bcXoXYS26G6B3dPx3VlD4YkruVMgdCs3brz1xmm47/TFDHF3TBsEVO0Kx+fY
BWdLstuFVN84O7W4GlsJi0Ds8Je0wErcxh7Pf4V351pujyLJKfrKtIkkb8qa
0chxTt2LOC9g7B7iRRvCnnJfsXamT98bpk1warhfcl8sO4UIh5mw8uB1K8b4
vPbKJV/nLpU5lc7spJ9ZJnTQP12HNONhHeVnz9QuukMVW17i2aSfgIINSHxu
jKsMy2Z93BtQSH5cWp0XvcleTLo6hG0PGRAIpO4DnGF/qZmISBeN/zPYxPNO
5zFpxBvipia/PTD7VdFlBdpWmXV0IPFK7D7a1l1gkP1a8sMlca0Xxj5MWGF9
cfPdWuZfYmasfqfJdXFzo73kryQgav7/GkHMMzVFIUjoIdAbnRKQWnl0UEUI
HSrMDhIRovGhRCC3xIUy+TVIT6ry4418TzhFtGYxzPxMvI7zN2hUrMEl9+yn
gEHalhoC6kyLGJvlPnVLtWzZWxa5CTiZ1BPg3+HXOmhMGq4XDBx5kPI9shYK
v/5RSHlNO2ycAlM2EZxkbHXI/5+8rCTyWcJaDVDKbbwKB94PuVA7UnTXUz7G
rA37yHQ8zBpv/bGT/fbS7oda9N+fnV/CS6NlMcWAU8YFAqvD8wxjALIteZG3
jCGQOpEBHmaS8NdWZgVoHXZKZXKdmjrhZ+AYzTcggAEWJUP/G+ccRHLnRF0m
ncuvCivo/bYSX26n8RhsbTpbV4ymFxBlUOTUNuTQ3zR4E1c/0Z3Rt8j92df6
2ynYpiiJt/fIitlRt4i88Bud9DhS3PnYTnyZwyWbiDAim251Y+XjjQXDP4HX
tLv/Kb95Z8OrAdZHC/G774c4HTNWt0E+i3qh3Nd+5ABnlD+qdB50Kg3oy7Ih
LPSXLLSk/IKYx1bu6AR1Eh1NKLsIw/2skwd4eDsst+UlzCWDCuSV08m0HEzx
C4RB7q/lSXK3liArz8Ovvo3xRnc85SGLQUFa4oDss2vLKsj/30GbKoS3I+2A
4+Vr7I4emtqH2ZehCQicMZX2rsSteW+G0uroqt+X0BiI+hrvcQigWfYvrsi9
6u9+5m3pieg5c9xL9wnq9UV9rebmwU0WYT8dmy1UREqRk4lp1Aj8T0XtJjaJ
Q8NdrFMr7i322O0egi1cV5DMNkjSkwzuhTQlmXxa0gGG//c0bbRif8e2DmzK
8/08bcgOoo1Tos1Ae2F/3aQCZDL0qWKavVNZIpZDR8KlY/911nJKf8zrwZZy
vJK6W1dmlDA5jYe44T6QAMdqsQMHl3Md6HfS3jn65vRUbhOHDBmabxqDTXxd
rWnxODDyUhDkczlQGa7DtQYiCdXbeUO7Y6UBJXGe6DSuor+DsOYuTCQckmXP
lGpmPtg2T5svt3A5QB8vlRH80o9nwnZRqhrNPhqTusFQ7rDOMb7Tap66IDvp
G1SsmDqDttzx7vtpgJeBmmqPY7GE0ngccP07QdnrzsF2Z1VmaE+gI0LBQzfv
uWQgdNEQHKMjBVf4R49FyJDwZ40PWrZs9qD/ewMAbnLWdet7jx14g1y+VC3H
cwb5f8DQOnKULT670Xb6A2C0iClBcTX0XzXl57fh9p1fiNmzcknb3eCgqZzh
8oWACdsJkwzBETsyf8vHxCw99Z9wyFH0Ldao+bXNrG5nGSNifTxzptNa+NIf
h6JXI9aIyiG5b+ZZ1Gu8k4FAY/vy9MiQj1r1Xh7+GWY11r7K1Pa057dezjiG
HW9JVMbyXtdS6CdtI6sKd7Fm0Xck2g62PNMB1SvlrsyneTb2R5ue/4Iw/pb/
W7LSuLh+I7/Nnc4uqWgzzwysa3s+q/NqTCnrWQiFsI9L7sxMszoEyEIou8gK
/at/NVox5CfKAklANQxIYO/5MhSSEcY9eqpJnfpJgMN7a9GIT6wLZInO8gXV
oahlQNFIkmew2mdMJkOVnggW2f+kQBfrY3nD2l8tea8ZNaQLpSwYngIs6zu6
ewJ9uiivxTReW0bXyql+Wb8O6m5EiVz+L/j5JKVuapxu684CUKIpfuTVW38j
OXoM0aIuMTGyOpuQthOD9dPQqsoFbEzpZe2CwrnLXhUwQlXd6Vqv+hhMmim0
MhVcV3OrQSREsGcBYH+94eG2dww+SHnRodTwi9X4Ld6Bp4TRYz782KFgvIfN
zgmOOGv5EdeFDLK2DNfoEz20oX50Ua/0y31tpJMHA+9IcXoH7xbPdIVJrMER
+N3yr1qUw1kDJrS+HwVcDME88TDw7QHxhrDM8caTuYTR61zLxkxS6HIQjTyV
iT36cHVHQyur34a5ir2s8u2OUvAzkPtf8dklAb8vgtADac7UJYmDiDTcPs0I
iVZcpHPq6pWJtMPsLxoLUH+Ia+gda9vlvuGFd7vrLRLMTpCOhQkBvRK74eTS
mURtZCbxiLzUl/H5jGZARmwQPT1aiHyJ1k9U5eG1kteLwJeyB5v8mtnbO+tL
QP9C5OtrXRCNkvwhIAKzkWEq0Q7q2/manV2VjWpgXRumgCtzbHApOo7ZgiZ0
k2fKRNYZjYYhCiIHcLMs+aVNjiCrPbp8PLIlQbbkeuRaPvzXm/UMHWuuuyU+
oqAaQVbHIUqlKc7f7bH4MNg10mVY0Y0vmfBneoFWBydynO3Flu+tQCdDKK/r
H8A1AivNQga9yP9llLxOp2Sr25V0wdB2kx5ZVOTqH5KNGK6H0QQaeXpxxnEs
6QiTd9rbkPsLWKEexufdGhcG6oXd8wW+jdJMh6xXGLecDTDXTBOicOTjuLFx
Kidy39y5L9JUqck8IM57CJ21ET9K35HHz9Itpiivqa/kzzqQxibs8JJfPCv5
HS62GgtJaqenZl5Wl/WWfcGkw91DgbcNKBL7lVEyH8xT7/FKjqZWnLlJXEK9
NNj/wlgY/jJSs12u9CblySBowXp80ivNDRO3qPpUqbG0Q/yRHrCDBpn7AIRd
9D8ODUZx55muQSL0/doHqKHZCCEnLPXtvI8ZicJzQld0rTqOXI73E14A46DB
UE0rTOdL/jCoDbz/gd5VMnd0nVkidtYCP500E3jog9qhlMAVLVuEdRcAxqUm
/WuwWOAv9egKsaPPpfd8henFlA5p7mKYnI7xS1KeNgDhAS0ybdh+R+AL+9Bo
DZIZ4OsLSI7M/aarjV3hVb3EKMcaz8P27kxDKF/yxfFNUw+Sz7zyiy/S0nOp
KOyDkh+wwX8olJm/vMSlYNpyAUCFB6MAq+UfqQxl2cEEY5lNhng8sUY1jNhW
MBb3lxadCzRpxHDcyesrqTXaHSoBF6R0D1uSPyKwEDuh23wxMV6Z5UEZRZyy
8Oeaa/lm7aDbHnQWql/uQTWkI2iQEwnx89vUf7S6ByVY6e36PPEnt/bdUFld
zsqwlCZqVdf6VA6UuWSZbwMjNvJAQ4VFdm0tTMsQSn2yXNw3ZoXtPO7KUCYe
u6Do8f08QOq9K72AgiTlZp1TkJet65fdBl8f3pC7q52DEQpZrThd7/mzfKEY
XWZ1vV3kg2f+Pcwm4kAc5ncSiUT5YbLfjZDoPENcd7vbzrXeegl0ys/ZAFBc
6phLzeosbB7vPVBtMEzJedejBT8Mon1EkyVAfqcWoCO+RwoD56Jf4TjVaVFm
jw5HjI/YwduE0dub474PhWfR0A2/o+ZzM2gkMQwKfYZSdMNwNDRjskUvtPBF
lYzENZheY8yeGPf1Nq+JIbhOYbG85jtcbJ6R229BAFRvyS+527Qbolwrbi+b
DWFnoPPN8t6Svfgqgg/I2E6YRK/CivgBqG/CyP+D14qbwSd1PkNl3TvFYliq
gi9y92rW1PsdM2icfV5OgyygZd9lWZmfDAY/8yLUY0PieLgZjlkTKesAXX8l
MOihctJWWIj60CD2cC89ea1nzetbpJ65uor/yiCU1Swi4QGf0GHwIKrLV4in
QbXyHD/pAB/vsIblbxmd8LmJSBMRCv4fITJtytApbF7/bda3Sen5UNoFQ5t9
zxySQBXSzfOovhnmtyltkiaLTNWsftqtQlSzrvl15lOVbmKca2CewrAI5yqY
vWi7zhpcMXyO7TV9sUSe/BGXFc/lMXqxMYLP9THJtPjXjvj8iRnKeUoHjAeW
yEOhUH8VbwCv2uwNfCIkKFZQPWOl+eMgewTDJNWsaT6pHOG8qXRgW9apaDTM
yu04b2yxks2QsekG+h83bFam4w00whQM/X2kIVPv1APec9+RtlMd6uCGfjjo
IiuZ7iil7FxymEBjLtlS55zAP890fwroO1Gvenf0lK7C51z7C2MgeW9xUrQW
fGLDIum+cGj8BOeZulZdeTldrCGWHr8e+m6aGkJt88Dec6q6OwVzicHs63K/
IkZIxA2lDvObPg0jtwTCGTYg72KyOZuxi5PvcbvEkUcljdkP5iqThNj61huL
ly1k/I5Pk7xpmbIGMbimF2j9+5puVK0wvcVv16wcOn8nR47lKXeUm2cbQ8u8
tkumYbHkn1K3cRRIpxLdDrz05KW3IuUjZeLkSWTqAmwDquQGIB77MaH8Twmq
Y4yGTJM206pSMneDwCRLdAsvzP0CGHH/jHFFqs3RZCmZ2VENZjEZBt4dBZci
vmZGN3tK5AVlxNCLqWGstIUbA94Wv/qGB1t8wmgPj4E7B3QTttyBrFh4P41c
eBXnwwd2NPcluuhhYC3amkpeoFSM0NJae2WqvLdA4JRl0yTvIsK1WMl9Cd66
TCuY0sN0OKkjyLPNJU9RGgPJurRDbIldycbXQ/6Is4MitIUEaP1Zi4vcsZ3x
aYQHTCGDO7S9jCSuGzDB7IUIJ7nWCA6KCFQJAUj9BvfoNLQzO1S9KtGC+jWA
ZtAS4hxBOXrud7kL/CNE6AGt0dUYsmt0inV4rjmDflwKs2Jw4Ilcgrcp0BVS
iiIUXzU8mEz+vwfGpdgcOxA5hjXjO08tmgJIKzBAnQTQVLS7T6jQA10IIEIT
fCD2YUJRBCuwCt52jd73JvVyFTaxsp//K3Ec6idx4+QApBUwo3S1p1cG4jsa
M4RFjrD1sUIjC5GtSsOjLoUoNSyN4pKFQzQQKE10K6rvjd2dQ1c+GORvQY9r
jQeqszbOJFDyUXACraKtAtt+5o8xMxBa4UvxAhUjGYIfGlk3zQRKaOmuVnDN
dMxknaf2DSipoNxR6km3iSngCboY4EHHzooi7cPaTQKwQOD9J6U3m5hf9zCn
LVr/KrkgZEk/v25AFfZaVElLAC9DqSNRpxdc8Vwl1xxORueZr2dfjTHtLlXe
jOIcfSjpQAdiP2ebuRQUj4bfECQvyFJQdXVeB2NyF+foMcdhnVGMGFfnurIq
UQ0+URYgN5ye0NyvRG4FOyRqFM4sQAtymiwPmc0/wmVdMg5zAor5YusVn1XX
z2m30SjIv1QTmwqSpKPR3uVFmuegudVEd5gPi/2RzXN9u/VBcttZY97jeTh8
tUX6Xdca4VNJj23y29Yqw4hzx0yX8SSfHRv8AFhoBpFqsRvTko4bD0NsL5bW
AO1bT71xsxU3PO2RjcauRVqRhEnqXVxbSA5X8S8tb/7iJaEVH0jBLKtlcXpw
dYjrGPleOmCb9eoZxGjX7hXpl2xv5Ax3zhPaUodlkoGi09xAD0g7l4eoOw69
fhOIzsnl5XyDMD5Ry6YKnH0iYjPXS1Zl9LhgCx27COF+PTpMlv8pTDqwwgTI
xsVsibHFONjUk6Ipnk069WocDzUhBFuC6rbASQds66wsB83c4xh/MLebY3Ae
S0ay9Tdk+nS8U7wA/89YdFHPIsyDY2chMBBWlJSWdw8Rda242+rcZxGnzTwz
o22ASKim03iW7jYMDdpBqEIsuk6O6Z3EdaY+eOUQALuWOzq+kEYN5LA+4hiX
IHVDM2cdEANEyDZTW4nry1u5dH17igpcImbV9cguhiqvBNKe73lOPzQJsuQf
vD9R6fFZQAMlfxlJpQT4wGuTt/oJ5zRfZGyH/2hX7S3XFbKZS7iUFSo2l39g
55hl8TH8WIy9sm76d542sTNf4QKs5z26VRKf+qCcIs4rlpUz3NBgSBe3Pbmz
cDjUMe2KmlhwqxiP8DD9foawYfMtFdckmGjD9LcII843fKt4S5dfctNjSxbT
V6CVqpPnemnw8t3g0ALfkwsxAYzKJkB+C6QrbjC0tAi59Q6TI6rNW0bXPHqF
8btg0ytNkjaardRPatLpKs+caXuWHgqxgImmr1NRGtDBtuhH5ae6K2BtxU6M
N14QEiJ/mXp0pS1TbggGhBqdMRYEHcBeMPcsz2I7ZcP/oq8ZAdaHZ0c4joMw
fbX/zruDW0+Q50SmC1BsL9/BBmky1WTKHahi6L1OW7eTNUMOidORvobjfgsb
V/Zr27pvOwSbwVDsKoN7Uad6eQel3iqtIfg68wjPFCCozGuZffNOjJoCv5Mx
U7Hv4QqXW+TLz/sQ82hNnupLO9HmEUTl5999MMKEWadahPTzQOXS8w0LQL0q
lx3nCa6nO1+9+AR5vdw2rkocI1VsS/7YHESQprSNf4iWss6n3moalABBpagx
JiG2EFeMNWUEZvJNUljJD5ZI4K+7NFGX8uWNAcbc60Ij6GB2nG7P3TjeDotI
dGHlK0D23MLjzG9CQHFQDWNhynehArITux+4hVzu/u5dPbptlv+pEl40BPEY
zfdmIL+kgLInLLQPTzHs2U7/awcW2O3s4MzvxB0AOiM3UboM5JBG4RID+15j
Tu/Uj0KfYINkMJ5EjQqeJcexKyCOC66oBJ1lo4RcSt0WvJTMnR5hWSfyPZqD
Kob38crBSLkfopN3g7Mk/r4gpZCW9dpM/Pj6fyae/SwewE5c9ahdJCmuvyZP
I1/cDLUVNb617KuU/vwO7v1WcIcATJXpEyaWtiwRve1D+4acdLHNZjTH25gk
QrpSxGBCwUjBMzn8EOHpL5oVf9mUVnPSJHJ2FWP5srZDWvf8F1sSRkdYGsHL
2FxOkqzD3FjsfgujPiV7nSlWAqTorYsy2jYCXtcsirQkpRz60jqvkLxxUQuO
No0cxOlAvTT1xDt3CNNz7ioJu9viXl5irPRfESViyBFWI4nIFI1R/+bJh6KX
MnHj37gGejR2+DeEVNq6a5+/Ut3rdARikwJOTp5e31CRt381GMMMZyLvXOet
tPB7Fp9X0CdYrFuEv7RedRdM0L0XgFyJGu8735c3GhBHOm3fyCogg6wjumhW
xrIrCBUF8R8eV6ALj41NcrGpXQSRNv52se+c8ZHZKs2Zg7kMlWJkMNzvEM+j
gfsbZmmhEZ4WxnLQFrIaoI2HVr8gj/GJ+CsyErm6V4/Yk+9mT3IGodHAhva6
Ub1l8mffUfyEIoBTodt1ooVTL3diJbmdtiJ6f+sVgLqcFbiQbiw4UREC4lSa
mMPaUtklmRTsmTqNdBX/lIGFGpa9sZdk3aLOoc2eawabBxul+BiXRX7VToij
kwLYAnxjzgEbltUtSFkioVO4rp3JRYAiJhzJLApKHCmkp8iyKa02IuReOYnQ
XTtXmBY11tlFckngH1s+TAOUrVHa4YdiMofR9xQrYqvLWpBidGt0VPlgGw6m
RaFPtePevsEQOuP7IE65FF7zer9nIdcwP/000PDHxKirPATKRvpMB5RjxlrP
F6ZnxrmXqhqwaSf5SukTwofJGsBoKy5TxdAYjiRwNER92CcfJg0JU0/p3kzF
sDFMwIHrn2G2SYHHGGQOjWzigmXHvM3XeY3pvC2PfyFelZb2g4cg8eHuRsPW
hL7StEy3zKF3g10AgnsHWmwwuoA8UqvYh7JRk5SpiqbVhbSyhZMMnM9T+Ob4
+/Dh1Y5IP55jNYhefgYusPuVhMccK0hkhVphJRDhGSiwmDGSpT8nYFbjC3Sg
lC2LbFGJ8ylJQypbil6uINsntSDZbEBAfULu9O3GH17OYMwq9aydijG4i/wD
hyL9z+DqB1Goz4+Taxqp5gAyFQkvHsWX/yZ68IwZhfVK11Ub44J/JQkj+sv+
wqWPPovHe4WGq2zXYYrZsOIc6OH1CodCkt/ikWYgUdRBPozOBdBQb5IWz6pY
ugo+C1xFG7o95gFUS2CrDhBaPSuXb1fuEbTKGjQxo/PAXuLFC+f/pQsQ3727
+uLeTWiXU0ECH71Ph1t46vb4qFD+x/c4YCWNDSGvPW5MVJerP+lFto7v56Cn
S/caoInE5LAJPWSQb68QN2ojn+tt7n+P9H6DooCJqFqCXXIzkMZLLJ/qN/Bq
QmrOaNd8g1N6qBBuqQDfsSvl+dntIRBZ5YqAurWN7ivixweBLtgeccrcb4Mn
c/6eB11CfB5aAz6TZS3zK7Zic4CuJdH43IuTYc2Ls+t9aOsvgvYegEd6PoyK
HH1bZX2PqOo8NwN+ZE8ZF6hXIy8Bwg7g+stqXo/UOPH/67Rix1VWLFYFIi8J
4p+9cnOLiPdhpCx8IeEix8p3totUueVuoBoWE85I5jU38CtMm9Xl/MeqrDNM
MkDL3IY/dtmCqrlOvgfKRJBkLHUuuK6osdAmvXnnI39o0IwMZxtK32IxcYe4
L0KT/S7DQbwoFASJYRcZdoWI5WqYThOrxVfFpxT1rjNm7S5rcJCUVun5EUTW
bndcm67ACt9u4n1PkRVZPYKiSoffvMzuYa78t4qn2ep2bp5IjpIaxMBBnEvi
6ofbqWy4wJrQag+hfWRno3HXqV/vDiy7ImoNyq5u5WfIH/X0+TdDU8yxZRqM
nfZpq4mVZxO9weNf/S+bD39qOIvoMlJ7MSXW8HqXk+/oddzDhsDJub/fTUOu
PTq4VYwSuQAvSsoNm5WLXVWINJpgaUhZ6+d94w0lhbr2bi/NJ+iRwVcJY677
fy8ZYPjnupheeSltpPbVQ1vXxgcIX3v8RXA8tjmDM/AwtT52SjEliQclQ97c
wuv8LBzEHjj1W9mIkHNQYkHadK29z4idly2PgOSo4MTdsy3h+Jiq6EmfontJ
Yd2WCSFetkSfKLfiFHgU+x3PkAyXw3pMsRy1e/O7uLMF80ibx6SfYZ5tK4Vp
uTuGCT7B/TMb5mEM1Ay5HRxiFlrhO3B5mIg0F+iPGqiqunQqn+TLLchwKNxm
Qqb+wDqZH7a2Hk6bXd2VyW+qgAEE8wpRnuIFQYuCetup1d61FbADF9wp1TXj
BCI01usOc73gOhAWxNv/+CoPd4mvXujs5ytoqgmTNX3+WSt969k4h8hiGeXM
73UVOxeyDMzPlrTrWYBMb9perGWYkQRozhlC2GVPrMrPkS/8MI7vtgVjZvgm
S2rHB75uMu1YSQ34m3kir7FY1TnfvRhTY15LYPs6qngI1J1F9B0itT4hv7AT
ci+vD78XqZTGcY9ARl+twB6OU31Q4D9eFpTrnxq9XVHPBn08AETXfeYFZeNS
L8CkHztgPxybj+YGGCpes62qO2b03ciTfguJ803orszLzJtwtP9Qi2Q8MrkZ
oBbT+QJkasXL5d94nYpKIAd9ARR99+OpyM8uJksxhymo99pmvEgRSotRLrR/
4er+Vt/bUJT8Q/LiFviYRs2R2b84Xf8tSXH/b6g3qncKYJKruQaiZBTnTsxK
HMzJxpL3DxnvoDpi0cH6LzAv3VMYYZ5Vrt69oTUaIWAxba9pqnewfBuFF2Kg
b4N501EzBw47rAEKhJ0+vL8yZPA/asGXkjY+7+uCabawyza8bqiiuMr2ywQD
HnrynClPi76h2W5TBqpU9n6CGJCJ44Fo6w18UribQgts2v3IGj94AxpPnYBJ
6kPIM03/xCBKd+6cWoYDdU0+tBQbCmwwPrz6xSvfWFOP4Wnb4fNXLLdNLoQ0
r4sLFjKOG68zPWgJ3PaaZAtc6PtcuQTgkItisLREGJjVsXbja/4h1l82hySN
HChq3mlyz3x5NEukDP8f9yzbMFehawMVYzMCszqpNKFiMRnoj2s6BREUx8qz
R516+9T0qgFlvfZDYwkrg0pkLMKdBh4YtlAqdz8hstW9u1oJ3K7zmfnHIQjc
yr3GwqFrdEnO5zDClkxbK434jMu8K1gN2IWbdy8pUq5WKV8qn6yKMb/fQF0+
jnG5PNBO39qPED6e/Cx6AAQeIM9FSSa51gljKdRZ7F2Mgc3N0e+0cCc60WgB
vIfAUvUrDR+Y+2doPa3VFrDx5UIjsFbijZd2H8fft7FvRvrlRvjgui008PWf
UIWfDCeYkOAfAm0RptXjndYMfBgUzZayA6Vdb4EoJRbj6uwn6IssnIIhFmFD
PrOXLv0W2Mdoq+59Rcfyt2TwhtgVHcFzeElPp/8uhrnAdjOtIS73djQz0XGp
62V9HGxaFneXlqlMk84z8eTNNEHoprfaUIQ9MHV4si+qp24W2SWy/xYOMwpe
6JKVw93OXcVrBcYk9yV5o0NuHiAnge6sf+Vm7OkXNDufqTcqhKxc5Na36Zl9
upo60AOHgzCz9wfUhMFqzY8Qj7vCls8dB1Y30/py+gO8iD23TIlhPo+5+GoX
+Q1ODn7oFEkrMafQPtik6hlLnPhBeN5OsoaI3+reDWXL50DWTskoxAPi2el3
TWsXjVHVhjpZ8lAiyoL86RvIaltNmXh8KhgzTHKDI0dt9qTdaVYh3egM1aPY
gQPnXznyZ0tO/qDdFhnuQ5Lezaa0Bb70XUS1qaxw56tDlfvChHXYxlEn3oER
v0knwTj3UWztFAmbYbfE6YI5CthyZXYWvEkJeSmRYXXOGU7rN3gFoPr5WjWA
AadyBn+i2mrs0R2FywEKhiaoXLg+V2j+6AHx66+DbkLhtqevAx/3P/ne9LU9
qr6hRpw5rfTDkOi0Lk+k6LK9aWZ/El+ZjovEUnfUHg++iEPAGieh5Zlk+5ge
7i3H2qU129SKL3AibrJWgurl8OoN6eeyNTfyk2Ffaq//4OS5cq8eJ0g7EMrL
1DCrfPqruF0syvoA5Gmzx/wF+vGRKZ1ylXT8ywo/19br7RdYKWTtQi5L2yny
dgilbC1IoDehajddjQaEiSmoJNybm+3I698AE/WeHCgd7awkWyc/sFWzLPut
VEji0UPPcIJatw4vCg259oJI4OhshxvCRNtbXXNUSxAe06Snf+J6PVQIETtd
EOmNTsAEinXPCa8ps9+wTcS5vJ8l49RHX4gJVEFuIh5hsEVuR90YO7J6fTyY
1a9ZCFfUpVcNV2mB+uDMKfo5J2LoRc9XpbRfs9WYjoNXljaFVBq+878S2xV8
wpt1C+zH9PQj9hu6DmU1hrQcCn/CiGEdDWsAaNi12AmBv2Q+yLBqAOGNKSKe
dZx83Xx/YYZSBSj9mBZhM9wEUNmR5Wgpde8jGb1K9BYgP4dZW2gpt4WJ5wDd
hPJTu5z9Xg6RbPYNtOPeaMNcR5VMnP/BArDcnlSxXmG/foVBC0xkqkapFo0S
Sl8Y/iCMP9CVOaMyQR6Jvv0jOq0+MGSRlsF3RahOkBYeZJ6RuTeXZBNLHgoG
ju3uHAs4yF6POh4K5xYI3Ja76GdnqHuqLNb79+7GSc7SMGdDJZ/1rde4DoBU
VgMK0hgYdMRBxWfiBtNM5UTMh50h477yVIkfOZyFb2deF83VtEg9x2n0ejJY
WIueqP3PULcm4LhA6AYbhK9uIFIFE6vegEsaXVEkUZgZsxxazCUZ9m33yC2D
wWcJuV1u2PvVIbbVhhRlghhfn79Mrb1g7XfyY6uIejaiLQ88eGTNJhmX0Ezv
SW80Y/GekDs0Ide9EzGjczVMgZPqh7K8O9DFwrgXPLnON4oxQzecMJRgOgpZ
zokraQfrbHWtms1rQd+Dt+pn+tIgViywBZYbEuJ1Hk+5sfpoH6WJw8+o5gbj
F9Ah7+oAuAblTn8v9rcUeW3YAOuHVv7gr87/4B3wlQd7Kkqiftnm6bJ2D7MY
QP8fcMwubiuTKhgujDUvmHr1EUFj9BIt48Ci8RfaWkIiWycCc0G68XDRE9ND
a4IRJpnFfnCgx9WfzjAQ3w/YkLZbh5re5qczCskzcrlnCpIVQcGucvLnX1vC
SXwHbgnyX7qbmgcy5ZQNtIO1guH4Nk8/md+ZaNihAI0t7Ia4219yEodQc6i2
q/sWM8X+l/iXj/00w267995R/bNh1r4CNn77HtLsrHb3Tznsv6GRm8n8deYS
NrZdcEfqB9Q2BV4VOOAmq3kRC+oul5XlJPipWZbEnoLlLNSodjlkz/Q617kF
N5DMTuFvPiBPaYP2g0LI/kbtqKye1xNe/hwRO7ZPUCu5Jx7djLtKnyFp8LSc
BjILl5z+RnNblBCHBNbG26btfNypgyC7U072/i1srFz5v5PUYRxTAWFgLGJS
yrf1QDK93JDb4CQ2YCj4DHxqk6Svmhh8AB1UK4Kwq3XRfhSaI594G03tNkvV
HY88zNMXC9FO3JwWopGVFcPsQsrqaJkgQghFKTr5udeh7mA/JPlB54uEd3G3
kArPXAQoYQB9IEtnoIu02tgbYQytoMU/M6Ltiot8qLQSTzu5GM6Jw/bI5I5O
O1Jhno8RIPkKXcrCMujhaUsEXlQ+I4H1n8qjokXd7XVNgdiDwV/S/f9RF4ue
qAQMtmyAUTvoMlCr0sQpnQ/qavTsn+XCNakf27iX2yQONuG13WfFXB8NOH3d
v4AiPbxfBmGe9av9JdiU0fXih8/9/0NmYEjaa8rKM50/00RCX8IuS4NT3nTa
Ba7V7IpolVJIcG9hgLLUpQFJHiV+mFqYROLu8LZnybMKcsGhOu785SfDNtOG
Zt1W+pLtuNTigl4tH7m6c7C+RTmtxCUJCiI81BKIBQ/EtJXTFKDTLnMRzqz3
N1S3UGh5OjyswKngV64AxqrCBS6FLk/X+Kn7jFiM3PpMd2DQDE2jC+vgIT9S
vFt3sp2Do4xPYgZJgwIGpYCXUKbuXuGG/u6Ouq8uq05rCg5XhfRBOVxFYUNT
Lg7DSFNX3ukbXXe7gVXPYkLmzrQzuOZd3tF+V2VudaH/89qYCuMuyMrUkG8x
77eV32N7U/I05QRL25Vq44XqMJma4HP9GP90GzUPkwIcLbQmAk3NQwQWguj+
yy1bpdNZxOq1aW5vnoRW52k+2K1wCniOkrPFAC7yn1gQcrlAf3/V8D2i1l0f
7Omf4TyyiCWyyNWWQBlwKG8fKCnsOc38oTkRBv04SWhBcOQAOGuSQLG5xzwV
NKXm0Zt1px43VtIyvw3gsmAXAwlRrCC/ubQHB9Wf95/q/EpIZlpNpJMk6QOO
9PPt548s+objw/M9eN2bZjVrgLUJouwieQnny3jJKMyKq+MpKftTzTppyYVe
Vot8pZOHQUt18TBzhx56L0qQ9ePzq/HbkfvaSt0XoQsy+RU7UEzh0X5SdDh8
auDbyW+M4yVQeSMo49m/yd3Ppzf+8oRKvNn76k1dBZeXsPqn4y9cOzNSICIQ
A6l5VS9mD64C7PdFB19uWm6Cqu/P6c65XSWwQ3Kfqf0xhQv9hVl9E93oIRzE
JnO2M/9O88k+YCTI0ZFBnOdgW0rPd1hiZlSLs8R7+N+NbR/WjK/ygyI7RlzZ
LpM0DxeUngRVe0E676c0NRJ5hqNVPiEoKoDxE2LcYzx5yj27nm9ep+JT455j
Q6c1b3LAIIQctwCXzddnOOGsKiyX1zza1FKq7rPl0ssYpP90HAvUMPhGarS6
Xm5I0SGwh2HzQJ4BFi+lYHJkeecJ7rKKL2dsWfSvC0Sk0YaRPM+/ylINeLpo
umq9oDlOS1LHjb2p1HN/0KnWs9B3VXEVn5qfuJWXUhp+qHXttDTE7HDuN8r0
s19Jiud33mf7WBoOTJnoG025BwbBPBrHm18N5ObN/t77ULXp2Q4Y/lUd2n2o
82OF4WV+l8eYFwFbwjFTxjrAMBoPeVce098/NVWVqMJkRMc2Nc9FmBh3ipOe
l/5Pex1lBtXtyYGdKO6ZwQ8EguR/XiEQeJA5Hn+r4GeM87AOztNzx+IpvLq1
0L76nwIRfe+R9UmkjmoOr4TV/sFm/LD95JWp+WDZEodth5SGdF7Y82GVEbF8
0sUQFsFyzXHisBMZuVgYg2ektgYW/5Wk88mdjenBjpKvmCHg2suNzGuc8tY1
BtDl+IG1YhZD9AUgbZ2JrmPKUGqdG4paKVwqFbqy9e8+uJfztY8Sdl6Iv+DX
lA503OBgssoyLn0609fI1YMjnlKBg9o+uexAwlsmjI8KqVNhMrcOlIpZpNow
OpjSev7DIJdJn4yCKI0C8KPfiP6agc5w4GCvpemUQX51sMSQksiOglOoVNfB
he8O/nvcPNyH1O/jgwf0jrj69M3nVdbTDb+HBhSVOn2Db6fc6Bv8en3v9rE+
hKvyavJaTDP177Q5Z6+/QYMosoHuuhIFXtrQXubkB5eHw5Y2uvIb4aiHRJpx
htNQcEYEmRxYn0e0ZHtXNp3OJnV7BFOeQsKJuV9aV7NVToc/4pJUnm1kou9f
aVGvWHzILlKq0+7lxwXz+21sIAFXC67BI8cHS2rLqu//hfD3pLUPwrCTAJa2
VfQkjHTIVkdjslGJHkh3pX04Zns/aMyk+wzf6w5ZlwOxB+R5S2UjhVWGgQ04
H/QwvEgvV9IoyrQIElwVSEa07X16dkR6l3Y6V0TJzTbu1fxAS8dGr5mB9U0s
OtvOLcAUYnKV1vE9e4nqXVdvlGPI/fgTgJD6mkANbKzhZCD4PoJBb179/ZS+
Tc3MS4xI+xGI/Ju9CXy/VuipqVQakuAxsHM8FRTCDnFmOqH0DrrETAEc6R0U
yP+0H/OQe4zmm5qh1Ojg3ZxQJRUYoHR4uJCSiEPcwihV3Kl7NTNq3p5bKVKd
Pt9CLeCOxvwtJipi/t2nRde/EHDW9gQrTvaBIuqiVaA7gpPcVOkgl7a05Cf1
aREcjBCX1S9XjdPu217ufrvE4Yoi6+jKWbgVxGdApOlngbxEZmx8staQSCAp
zPwXTKgmBD8o3IMyr+A0TQp0OgMeZ86uKxQejZP7J+vT/1GbK9MyAtR0v6MU
yGNOwZ29l6Rjp20ZYzIZsSY5pkrm3lKJP0MvbeAtgY/p53CJ0NJjWjfwTTsf
kJbbnDvab4QE/yfTrEwgsqC/QFtJspe+LX8v96fl98uFpsUv/+ji9FZAOvXL
vbkeyKDWFeDnslvlLI9J/mZGr+4hraOpC1TSMo88ZqsjbIqZDbC24ror0EL0
I905hIRirn3RlYdHpZjXBAb10rJOewtHKPENJFC+1BCBMjd0y/4w8JO0F0PH
OvtueLAo+MvuVLu6bxXbS9ky0PjjV8ywdiA98+68C7FG/jQUxvNYhaSgbQNB
52Ya8wRTreH1eMLVDXwqLZwLicbKanI+MHgH6cHOQyUrMi9S1C9uYrkDe5As
7jYc6tcEUsmNexPxTdyOcgu6zowIsZ68hpyxeaSr4zXx9fV/QdOVL6V2ZrS9
Nu4GI2+X+EqhgS0UM4JRUOZXhNo/eBeP3EjkebtRohFhmTyD9gUuUNXlJuSj
1i1B+TuRg2DDVkOkPftDvFZ4W3RSQqhFalMXw2rMzImeqI8VrPw5Aqv6E3J8
jREvEXYPtGJD3xf3E8lghFsZTC1vZFoTYTuhFr+4IN3rHn2slVjNMIOW4kaW
C335rFt1eQFYrSt+9HiIk3uMdGpIaqFTxUnZmR6vNsFuDkTvmQEjegY51EcH
BjVnAnM8im/X3J6quqbv1Dd0sG2w4msxJBU5TuwhesIPGzJPWQDukkKTkVFT
8c3rjuhtPDr/Q4bNcABOotOoix8w3KUlZIXpA8aS9pieG7su8a8rxTF6Is7U
Qnh9JNcgGyUEBkJrbyiAjqO54uvZhYwtZn2bpMjMUNXEEXo6CPgjuwAAwjUi
zs8PM9cCFmUxXD3az7TUyXEPhdOrcK1t2HqEYigLmo2Gd9MFLvsaDqRL6LZ6
C2E7QYwZjmwN0+XPbXoo0jnJIMmWegmqhIUTpbxToxq2M/r/DPrQRpGdDlHo
zEXgsiMgsj9eLKnnUgHZloxn7Wmj1JL9UURmqeP3wJ4yAAoYZWzphQbQqIXu
KGkdjnhKX1n8RK7H5jbDCUzTRX1DtSImm0KxzhaIzP9QPWZVuG7xWb4hr5yC
Hwnm1gzOPQwGpbM1VsjA9bacLUoiv12JnM+mMP28OE/sjxvhki/IVLukftzK
Z84l7OJ/xcNyi/ptf/2asy1RkGbhyp3Gvy/oDgbxQ5p/S9mCXeYzGadFsAQj
qz8pL6q7lCHZRkHO57pCuhlg/O8L6mvT32EH4/p1ASeNC7jqwTJUBtcz+Xi/
Le18akPGXV6tAiSAf/3cNfYcWpzKT21umWo2/8dqxVLoJ8Htb6vHuj6zhhlq
n4M3Rp9xGag/RDJWmLEG7amMg2iw4eK0t1TLUt3VhaeePADC7z2Q6kmJLZ8o
FcmadWHOFssrJjkzbfUI/0pXv23OLx61w1MGImUGBjq0O9GK3+3kd2VfSVXz
id2NCByRAm3NaQylCfHtzUsH6QLqPIXcbaqOkD6cdqQzipuKfWpDCfmTT/oe
Nj53rM5hKDzrn/+yIydZbf4qT+AIZ0rw/XLUakS5KOabeCJfIWtTUO1tVTkp
ZHHrds8QTN3K8m5ZuA3paTco0LWCZd+r/AzT4RM79gaA6IXqsWxEqY/OPTjI
buxTfRkARJQnwe8nVRtmzSOSBDLK8H44U37XAUIqiDEFA16YaC1ajkukraCl
NeG1ezrx/PxhHezpX+fM+6Bagpascs8JrVY9zDIM8Zerp9FJsBDI//bQuqrb
xXoVcaqzVbBp6t+uknGQMDOwiEV0RYV/WTpNS8kpJ9ACfW2Ecwb8wReaaJ7h
nB9Cb+jpcG9h0LLi/Y26gu2yFCUO5ukEFgP1Rs5Uht2GkSujj3upIU0CfW2/
t6bPA/O07KiJ8d7ree+huD0Fqwh/KRxAK/J/YkSYJF3sL7L02MJBIApFsGvY
SHeWfrKLrImqm2fLR3nd8MdNwbClckRt9cTMu8+ZoQ2Rwyj02gRrn+oJbgWa
vOWN4X9eM8GIWFCh8iSewYaYBAQXTrTDeVJ1ye9fTEVzv02uVtpXVLR22/az
BqsOpPp1HV95a2nLO0a7cnoj+JYl45uaJhwI0q8tIYeZwPMCyDurn+aeSP99
X5V25RnEg8RneAmiM6LZ/zjNW2JUvwO3cMPPcGWjVPBr4m2c6/RfTprgkw5j
qPwVEnwEFPJzpAMoE2O9v2Nc+DSXoSd1f2uxefnHTdiKsW+AMM+pBb//Vv/k
odmKnX8RQvDCzlvNX8syqQ6HGeEURAfcsTX7f2Pg9vlpRHRDYqLHnt9ki1iN
SEqAEtlmls2/8eGGD+q9S/adyp446LMadjPa/EnoKQKdw3JjGyhjzpcdRye5
g1koLrnq/O4wiDRHNhbIBGRawzlu7uQ6wkOdmPSQ7bJRg27okEdS7J7km6tv
aQPHbkEYa7RgFjAYYsXiZfvZyek6sGcik2RdA+G8OienbVvcuqPghlIlt6LJ
s1HiuROzi8zBJgtAX8Jniha4RyCnROkWNualeLTnchfmkI7SWYew908q0eQh
ApYCexxkaYqpRNITzcniZw9gtWtd8OZdrKuTnXwONktK9IhkE1sl302hNeXa
P7qQZaDOeo3cpBUI2+DOPls9aZaiof/R27K9dYFwqVgrniv5Z6C3oS3ALrDq
OyMD/W/HfIHMIBtZCHPoVeyuuG2EKx9bWLtmpaS6b2HXw+ZuVquiMkBCyjiX
+w4A1OamjDWaQy6sUvfGW/BdI3N38O8GHyRhzmUUtl155OCmIinq0cDioF1N
fJHuYRnkw4YVE1gmKE3urul4U2+wwoZW5lnVAfpaCMCMCl9fO1DgarhRnEjK
vP4WkNkoyt3rtzfh1cO6DJr7BKdTp2WyfEWmPpLX0SEurpXIUsMMUwf4aUIF
mU2duwVRdnHtR8gv3wuisosunUIpuM/DRS0JXDZ1bEIj9mVCQEtefzlmAjYO
oporaYVqtxAoDYXHjvobMI3sIAmzyX9ZjpXZUbh/K4sgF3F51cQVs7UG/tle
2tV6iJJTa6IfP+s1pjVggK3LIsQBZyrfEJmNkfU+aIGIZ9bJZX5z8lqx134q
uk9xDsYUI7OkxsBW4gRBv0tHHXjBeF3zAGDADmUh4DUBHKQI6gfhL69BeFQK
P/82vdOhlHtK7s+3ZXoCocBjFb6p1UTA9sNXn0A34mBYjLDIPggIA0LEdEOb
RTkho7COmu+8Twx726/FcBLIYDtaJdw0EW4g8DhtX49pCUmeGvDBaiUhgXqZ
nQUaI55NLlcrtYxPMVvLhxh4RyFG+2OJRlWTVvAiy+3Y/NDwwCd1uZpyG4dl
7Et6gWzDqBx6Z3TVUw07JBFGCVIM8/Dt/Eld4VnfXi5QFGn/jq0kdVQ6gHl0
i7AF5EjK5OYeISz3oYfhusdV5wjldXjrVubkR6AY2/wpvZZ6Sw3spcTCzUTi
WfvgW7+iiutTqW5RwChnSScMxXUMnWIXHOeMGBjEbP/RNINcr/V3D0ot26gp
tFTtFJrfxDHyXDRwz/+6yVCTqV/fV78LzEEr5f2S8VBsCp/7OYwy2WFjyWfs
X1BUxRjUPj1ughFxZUK/WPK4lYbrn4jeM/SXI1ZNQ3GseO7T0RUTJahoCOJH
qEFjcVxils/MXc6zN7i9zkJrTKmvvA/CxjsX3c6hkw2/FHruK/5PenqaiBYJ
wD+v5oNYEhfLs0YEUlWjIHh/cmjtHGmiHKneN0ZEGIwuxQvcl3zzXnjg3cix
ykGd9ikRpd0U/1NARFcbxmwZkI9H7VXQ1HCrwusZqsJUmVsTM+B/S1p6Ip7/
2iKE6r4JlbSMFeVZci2BWQ9cohhw1XhbIwBSbUlpBRIV9cfbkqs03ti68A9c
B40Y/sIupxrwj42r/7W+9SHh97GGrxOA6lviWNgJZM/JoHu1yrbuDtYNdOU0
nkKFoYSMX0LOvZU6aOWhGiBeCCcDQPJatj37KJNMz/wTZ26bbU4hGtmiYNCx
nztP4F6or86sFoVK5qIXq+XyPhnqe/+h5DyJ7ySoQkmdlEieFUJ9AmgqytpQ
H4oo4FqP96PsPrysUFMQv243oUlS4M6I//s+cJ+b+VabsaRvkFHfGYJUgV2k
4zcpcFBT5F1LiNHMOsQlbsAhIefi0xVtwNhS1A74V3rlghO2vUapF43qm0gm
dpx5pOvu8Ha1PHMJsrfDWeO96SErgAs2h/kkvL9GJ0WFm8wEjWll7XJjE+PP
t+ZEblOoB6hYqWyYql9mKSft85pk1hF3p0ZFPcx0q3KEG9qJB38vzzW7Ml8C
a4Oaft8aXZ+eEX7nXAeHmASUuwkBKfw0AdHNNz9DBdqH7xv53p/1eNxGoaQD
6DmCWGIkVRDlcRPJEyLk3u2H2lpDp1R1x+qsuU1e1QjV9epcurQOJfu9EYDO
5JpAsgI/xTdBqjhYcfYIHoY9kLqlhjsU7YXMO3tB2S8u8gVFuJ+mfviDb8n1
lz+ASyoP+cLiAvb2bxYtSJFm8cU8y6uQQ1yc1UcepEHB50K8/fQaxtjAw/lO
H8Rxo4C9p9oZCx051vtS7GFMdA6blwPJqQwKCd8MCCHVKjU/IQoDDN67grO8
KYsV6ncMrrwDjojBpvR5oVgtRPpdo6H+neHZn/J8i7neNqomx8BtB6T6lvcT
UwVRcDcrAybB9iiwd05EviF+OH/p+5Pd2k/YEztVQKQka+XyUKzwvCJqUHWe
xanzSmQoAhg4+p1NUwLLEP31FfGgbRl2y+EvpuWCnC+et5mYBvABvCkKBzD9
hHICzZk6xYWocFp9IPmd5YXTtqxyo4lK2xE7S/B6iiXnC5ZwgpXplMihMytX
3nN4nZdnWKBa5jqLOUzNeV2X/ZyPx3EzItZ/4SY87fZQw/J+isCNRY8A1d4g
dBrypHNI+ooEF9LqO832smRYnm8N0bSEfudNPwFlNHiLn/GnM9hqxCbf4/Z6
8wNJO15D4iI1jxKv1LNUozQ8UAZC3iM5WmMtCDqxzFo7J2qqUhWN1Vz47YX2
YvzYNmim7ivJw5QiY5lnyzAL4BNq9MtuzWMeKY9Z/p8Unq/BCAP3mkmcJI0J
FUJpjG5CZPBwD1PERe+hyGOxAWIghRMHZMZYpe3WbXuTm+b2cCWehD13xTA4
vQKb86fOwKOgWl5VJXtua9Xbd3Gqpw5PuK5xUIyXXfsNVpd/9tG2fJha3Y4O
OioWP7GoW0JcHadrycMcQSV1omt32pG96SzGkApU54ckcW3hgdVar1UM5yii
sRrXRRhdJTDRT/L6fb0zLDdwBwsqzK9CKTAFHN1BO5gb0e3h+kUsJUxmAhoK
mvOnS89XGYXlCQYVdtkjjjU3n0ZjfJGQRep3wFnHYIqDIhFBmpNjEuDgcQn4
yQJ7+j4B8fo8HGBpI9VOKzKAG6Sa3PIYVBlvIciM+1C1cQQtx4vrobHCQD0H
PaMkNMI3N11TY38fVGcT8IfR+iSV75SMc85A/eD3p1bBI6FRtRJXW4vntTMh
YxDz8tNiaTEY1Ufi4/1UYCIxrD+84WEOyj4minknCtMoZ5Mc/moo/s9zSEcl
ZBIiehuJb+4ccxm/QwIcOq2mtbvB5o/GcwwVdpCcFVjUSl+1MyJCIVIc+4Jn
tSST0OOdkdGyf/WLaD4QlBb00akcpL6lIdPHPaYsv/BeXtsNX3lRpqVjN62c
ueRiGrCh8Q3BmlIew5T4nMCDSM9x7AzwtrxKxQmAQxkep0jFs/QG49HJam0U
mnUroWipL+Cq7AoaLkTufNOfgKKnHJarXyaJlxwlzQ9GXJgnXaK4UUPR0W4P
usaiWD0he4K7Mi3DGQHNjv9VRbMjGVv6W7qF/3/cFrNpaMri0npQGRBKGNrL
ujO9k4NZ2QdrNnAPNBB1LhLu0Dmv22Ko5hCaqs5Hq3ZMvr5KGixCcYjsgKZ3
YqwAfysrJiuefF0MIy+gCDzDYem4jq5XMSw3fkUuRxMOiFyHKlNL9UFpQm09
7r0F8YJO3lxlS36oyo04F1wqnNXlecd2DjhWQgYceAOgNpC76Ep4P5vH48JC
9YxJdxjsWqjdoZRLzE1bi9XF7vIRzcgh0x1DuJVLvzqw4AdRxGQDECwFsaYM
UFTwY6VmTfPrYX4bALPEr03qHlC89niRN9pqMadD8kGNVft4WCP+6ZYJSD7e
2wj/bPWEE3cH6h44BBGJ1Tv1hn53HZRO0TPQAofY0RVNZkyQPkcBlVS0P2+W
S+9zePEAxviVwuYvGRWO/xDED56ko07Xk/P8gtqm1YG9bQVUaK/e7Qmt6V85
/frUb+wbKu9JelfdXtJCPomzHZEWR71yKrEPTg72sULyFzmCSbXYohm/hJfZ
L28uXlNsn2AnagzZENFC7UOFF/Miq7tI/twVkubdLx3u5cAtmPFJoe2Akd9G
VWS1ktwpbgcD0y1BmZf8bZPnt5v099rZDpwNNAzWcAfVhdSXyXN7EDpCW7nL
2jFdAe03oex/Q6GM0c5wxhJdQ1Uj//szDeAehse4iicxSnkyPdfRpdMD+eWR
sdBRyr4mOO82ccfnc+YWCYOPjT41R0ypvKPGVEm9y6ql8mDuqjRb326d4lJ7
il7xVipw38kC+eU+DY52jqKyPsEI5RITdmK5w+KYm6dfu4VWlzgbLedjzPUM
N8fbI57Z3ZiSJW9SiqTa1X+3BcxJqKNfuYLbbD6kn5BjA7SP6uKme2RdiWpI
m4TCG/Nyk5dLV+04iXBvsuPpr30RQZZQKuP+H58FOlX7H30gJjb+17d5+QaB
rgnTccrCGfHrhjzg/RpI6chfH3pPU2pWaSWhHWj4asnM5aTtZkNJEOjW9IV3
+qWB7gvXcnxrot/R4lZbfNsST+bwP7BOlJ1lLFjBP1JVm7It5+6uynhggttK
7YNzpyvbHQfGzXxRPdBAS7CTYE8QHgVV9ZsuM4yxp4IExqWin7rJDZEgXBlT
UcCRLj3DUYsAkVpeqJqX0/3UNkjpF2rDY+B7e+rM7Oyh1jUZaTPeOqgZeV1q
vi9jf+Y2dMe4NzzKrthTtCiI9wvyOpfLnQWo36UJh0gHo/mj8HjjUh7YfsyS
l+wSkBikoi5lM0Szs9uuC0+GinQ8AxrFXKFDOvqWWufNmqT4NztjlZQAkIsa
4/zTHFXVkMZ+K72CyWM4a1PUyqWCLxYnwHFeNuGHMU/GXhKhdlTpMuqMaWhW
MxPsURB74f3ilZAdNLgg/XvhdhpCkqRNdAPrvMQ+eMT6Vp/pbXid8vUohb+O
uMskOs75ULhiAkLaBOl1UEXBVQZXsxFaMnJ1EJ2rZAQKCsquEbe/vovhLwns
5aMu96e0LOap+pzYa58lWTqnF1NUZk5qskQVdJi9kmGvy34DJShdeNG9b4f0
+45YnC0SgZEDpHmiMLxysNs2iYlmhPPazWB2ghqMqDw7Lwl1MyHeKnFboElD
w8jH8GD8eENoBZkzGLSdjWFY5WzCi0audeo7cf1Pou/x6ZuSXYJ4IEk7gZsp
FRXJSWGXbFlNAZHYqNs18QkwXDYCoZ0hMTu/WBKhmRKTjQFJx1bebtDZOEfx
hKmti7UX1xDFMy9HJ0ARi38M1P7TwhpStphsk3Y0e19sWFbfNO2XlACzBUeK
p9+qsDhclMEjJqxx/zrPwr7nbl7yv10zhxf1TITWiC1CWSdlKixkyeOc84YO
RheE2GUkw+DOOl3JRU77vGljm4giZazMEkbAiR20F3uLnohdc2voPSt6tD3P
8y4jjbRuGE7/j2vhquB6NcXtgTZsEi6J0lMAgJcSGIWqDICD71s/j5Lth1cL
iK/oB75sCCjQxvry1Tqarf02o37H1KHj/sUclgPpzNH7/yhXwskYa3wlHBdX
7ARRMwGjb/ljsdA+TYTQvfocjDt+UEchb0ODyzXba5zPAJfqgTmOiQXuizvY
prJK3sNmK6+D3nPp6XVQIvVpsaLlQJGljhplnT1jdtixZx3XiIaTikMsyCFZ
qWUIe5606R02LWFvIKYPJUr6tGkE4KZ+5J8I1X8Bp+9BYqS1Lr4yehDSJaT7
/S5Em8WQLiY8UShb5ye3twlVkI2/LiTEB4d4dK2dOtp68OZPHkW2+/vT1b+H
h6Dq4tbABW8doZY4t86Lu/De+DzzzjEdipXQVAHuw7yWxb2W+sGj3E3JaFCl
Y/CxqD1v+lUKzbCxoYCat4Qh1S7qglKdZMu/Hg+KustGQRZN6JXts8ytlDFx
A/zFSUl4vXiB6HLHR0vbZ0R25KBpCvSzPa/0M0VZZdeFh+rPdcLFINKmCofF
6Xpfd/lnTYeY27Ux3SG2hMzssUrod7R+5mAtI8Nu0SZoz2vjLZYXU8m2zd/T
KvvYsgl5EvY7sukKGVDoQhwwQrm+IC66UPVC+7EwOSyRaLHcdj7qLVUNfkHR
LZ9J7NGuRJB9zqu8i1cjd9i04EFaqMOg4d4D3V3FldBeJX9EuAl77RH8oWSe
u5+tjAZ0asgARVb1fH90ZsUsORV7rJ4w1pjNO4PdOj8KRZvEHbCtx5EeU5uD
x/CNDdG0oVGjkwe3D1BTr+NjDC4uRC98eIij1v7EFsG8kjQ29v8oF/uiVf9w
/8FM5ZsvobUKZilNjl1ItNHCy+0GbPDHIGcCYhAI0etvi2//RLqZ7MsBuw8B
rjmCswt/LFWWKeKZ8fBu/euCYF9ZEPS41eTKQk5VLDr1LiwfXjhyeIDCpzJp
V2Q8HoX11s6uUNVtNF9SsxtGo2CfAH+I/IyIlCYhStQLK3bqhgWRAPDRCi6H
wenvymt2GCoQPHHHKTEjhUBi+kwjf7+5lT0jtPGiJM9C2nUnabTNSyauOmMd
UpRYXuY+WPIzpdVBL0I9sZLyIdL/i3miASfIrRYECfbBzGUqcP7Pzu9TOKav
LgdtxgfLP80dAoSrJpzHsHGZa819rZjdImdFSLcZsahLCh4QL1xasBqjJKpX
+mBzYdTFO2lsuxAwerF5mjQvzEedHudnbfeSnEOJENbSYO4zzmvcQYa06Hec
PnLV9WntJRRgTUxAEzVsRUp7rq2A8ZWF4dzcHyRXlObaOhg5VKFlHaVHur5k
LuY1x1Xm3VMbAaAGEdWIY8JRpDBWvzrOYNYNfXE91fnoInxYhvP1I7jxpI9P
zKN/3T1vq2gdmDMpqUdIBQMsYKEDgpJZs44wIT3WvRMqKo+X4UMJ06MKli+f
QjhTPtjjWBVL2SEpO55SJemz264zawK0hXIRsHNqYvSJ3zz94oEqhsGH06Gv
dCvaVll9Y1yrOf/sGq9vL2Trq5WXU2ICZJfpk/GhYzC1sThmBzGWQ762/reV
tvlCjtpt43Svwp72v8gPHg88IFFry0QVOMRw6fMz6UNBfH443uFknJIo6PiF
7i6drZTmSt7/3vFamS98zaKFfdLfiUV76P9fUI/zndZ2IqvsclgaOrEtOq7M
G60RYh+PBo8svPV92a3+Sih7DdYYIIfX6AeQ8g1ijQG3Lg5fxAxaCArsmI/C
Ves8JuPy6WawaclLfxq02Roon1zsa8R8Ep6HNFRNCQx4NcdszJLa6tWVHJwh
4g5nmDXrg5Mv2GXN/hIP3NTuCmz3Ix/uLf3RHdgOwS7NUKJxSdxynA9MVpTq
zviz0aWL3KS860i+7pgXkD7yCy6tnG+qZoxzA2vXyqNMN5IWVtlQ/ZACnILG
z9qcMASHZocejA+opWo40jaFOKD8bCN8YU63DZ+qul1enXfqh1cgdUtxmviX
zyHNGWeKAX2ndjiUjS58ZLEqo4efH2OFUP7qHNtQD/FOFsKSi5YS+aZp973Y
MMLvsBTtJa6t17hZxED9zpDG7wjYNd/TLLHGQMGqMVPlQErKDwBo5YPBVxQM
AOsZKvD2O4jR+nHKBV/4a7i8wYx3qWCgGAyGDTZRVfDvD1PEyXt9KZDB1YOS
HWx6TMUGj5uVm2TbqyEhdyTFdU0CIt58nWBztAlNCugXKqrDJlGK0pH3EQNg
720Ts196Inh7DGwNUDt3HWJ7gP5SyPSFGo04A2vITwguaDgSrlcIN6Mas6su
r3MEGHm/200HIeJo9SYSlJmK0O87z/2JcIxC2x3+e+jceM622Xi/wzXhIh62
cszMq8R7xRH2dPbrEXOR7XC1Mr5pjoZOvZNNeud9R90Nk13J/d/Yfl4KzDy+
I/69MpyZBFrQzyG8h/eaMpYRebh7YxDY8quK9XJv9Zss+DdgDpoWklLTdkSE
EC4639KhvxXQP2oQRgQq+7Qo641AjSL66DTGcyjEpK+V27LDLOnttmEq12jC
Nvqq8Q9F0B0ZbNpx1nqPE/NRGv62MaG77lzMusyE9xNHGSjUhC2LHjuVN0sv
HGrMNoqqKTj+oqOgFVRaAaknvL8FMBvVO/qM51nQLibCdu2m9x/ho4n4Lbh1
LpXeWeueuBi19LcmGvP446Cnu34BWIZ/uWVB75Zgw1mg6kdU8gxPxDPFymHC
Rkda0EULP1hA0mdIvQTDOgohaghvzAE8wEsY79zPoD7WLrrZFJ9itBnXiAzm
FJQvTrYo6Gry56AP/WqbZuPY3WLJD8dH1Ipg38eCi+CzabIHFD54QIszfRXf
J6GTE+erx3NAv/d+LIyd2Mv2xGZolJwhXeuviYwrRYkwQRVYNZ6MJf5FPS6Q
jG3y+TWKF0QdZvUn6HUHajUZMLtK/SdKdNcF41ga2q91MBJQHE/2swhOw5Uq
5f3AoiUIEb2mGwk6NUfB1iZwz5EupeJNy3LTXcpjGxlnf5tDwtWLVosgyWdA
QAiHR+jxloITYv5wliwX7OthU/mN1VtpUM8KyDcDnOmPQjpPfqjGrpgS6N2g
dBLBXGiTFHkC6mzicgnpblol0otTQwXJbRdQBAJ0A61s1Vyq7Z8mqNll/Yjf
ohEMnefO5OBS2d6aeUNQX0xuSUsImDok2Qc7UdVzO+NmtI5OzvTZNH26RpmE
hNaTDqW2DwZLDWO780IUJe/0FpygqL83IX1Ho567GOsb+qcX8v3pN/2+h0c8
BkcET1+m27POVNopq2K6ON6gFTmvHu42OQXciOmIlC3v1EUoqS9KL9HOZ9dB
Rh+aTeXjcT14xr44C2Zf1xhItNmwYDrn5NgYYUfUiQau4dCTTs6Wf9W3wxUX
BZ3oVm7P4OjTty0F+UgQF0y0Z9fkT13Fhx9Ksr30dOb25rsezsBzLjyI8yld
AZnRpsnrOaSuRJm4X9I2tnouItcEqx5yLFKnOXABiWF4FcNpkLpMe12QanJ3
K5dkOoRc06C1nV/GbP4IuHePeIB+kE8Ziy9KT7jsBNmgCCyrE/ZWJl3NrI7G
a+9jPxpLQPlKD5oB7N7iWNqSWE3g7k1WglkLy3rFhif2PwK394SptSDo0eU+
tRiOQAnnRQ9Hgi2lTG1gIIE5Dw0tG5xQRLNBS2dKHVVCt82LwPvVpRJcSMuM
uiVhr+x83BQNhUlRvcpY7q14kBGwLTMsGgXtzIrgaFCURDi8ZHMjDvlShpgR
BVtcbqU8BCpQHtHWuZ3zPtHrNa3svD5iziJRz3GCOvpa2sY+7lRp43pPxmZE
W50keSZgYWajMVhGan3dKWRFWsEYN8c/PPQ18GrblZOxRAotpVbTuDQW6RbX
i99aBz3fjK7+s1eWMYYxPQFYKYWd2gcamkmNQ4h6OoYQXWaJH2TcPm5Tqpzv
V7V9VMH2Zur8hejDHKdZjv4QByD8Pfrf38yu5SLrt5rEZQCxgKwF65hTKf54
As5iKI7Y3mZ713laP2u7qlqchtfoJ/c8ilFCL8KCZA1XfPsG6uzL8HjK1L+d
ysvi31d2wDvB4aMLZqdnSjLnoKHAkyeHETXaMdDJu7jzxSr1a+VLQGKzGkez
y3V/oH4nJ8WW1nkuJdgoK8odku+SL6GLbOMOlGjEx97OHVB+avuusK7E5Aa8
88XnZHCbXdLGnXNJya6QQSzKkCJv364rh4rQoJLWRH3BaYLRgUVkGz3sFHA1
u/UipR+hh1H/JqOovKAA4be3Nqfx9SHy0/UrmElxBXp1Pqv8Xxcz83zvWjSe
GbxufGdPtZM4MWQqb0B7cY7VlJ0qdA9TNR0fCB1LSxQOxg6I4Yb+JTz6P877
ZA79B7ZsmQJbR9rWo+U/qN+oFhsLbuKig2y3/yoZGWjos2bjyS6pJvX85Xc6
CsO3O00DRcpbwjCF2UePTZMNvUrU5zWj21iRadthzBeB6PyYV+KOP9JPY2fb
hetKCMZN971sh9oTjJLOEzKCMh3dMC93UCcpvFx1/tdvy745mJT2iNfckKnX
SRizvHnbTDuMGaqQyidfAJ4VmxfUlqgKeDvMzdVSkegZSRIEimdZtG0GnhZm
kTjGY1Y6LWlpTSCh42KWL0/ZuqivXFisQP2LHKWGOK09aAubixLbGR2yVWWs
a4YLEJAEA2P5bco4zKvemeE4Xellha3Wna/aP/fh29CpQgmpzTLuWtvDXMze
xDz8qeUGpHa6luMRiziCPwhCYVsAr44LeC5ZOFTdiRjgDh3zklmNl3l//E0C
j3B4nYdHvsPspSQh4b+Une4OeIYmho7hRl2QPJKjcH1glie8HLd1RZukQA3x
Rly2fD7hhRAvE4rh28oYqpK3guore8rKD6S9yrkn4t42eDnAiHWyvP3Syhoh
HOwKVlkE3JyjFdqFY0L8pENpJfWMDUxVUJPQqrBHuxg6AcVag4OL5z6NKPk/
JBQwMsxX/5Mjz98SLURY1ZWgPCDSSQj+qiE3miwfCOsmosJ268xHn08Z9w4i
TsK53wDpiaZ54PmgJ6XmF0mnoYXlCstIOsBvF4Ou9OfBeqqZ/GBrOwSTxHV1
LLn0AkfflugXeI5ajqSbTrwqAXQ6eRmRKdlyBrUv0A63FAOm4PXWregRlzFU
DJSGOkl4p9E3AsBiaU10JmiCkCCnN7EU7LuBvmoQmPi8I/OvaQG4PeVWwEPJ
My0/x6/TKpFhuitmOCgjWHHF3lNaD2PraDF4tU3E/lBsoR70lSTrgOoyCWX7
tItk6ef4Ngac4TZazgpUghwognH8H6A0qQGEwC1aglvfQlz24ZTmW1Pi3zuf
XEjYKrXOxJx9/cvzUQcxWS0nE0u4ARKbsi3rTZNSbAozABWho9iNgjkT+4bG
7lZjVLNs9/OtLuUyMrmULVhZmkYx88XrmTVfCDwrcJfadBbk9+qVz2meo3yI
JdWxTylWVuVV1DVApWfFD5AuXASAKDf5wSRFaZ5uDoC6ueYAb016S2n18T7h
prItuQuLIhiAb9WiCLt7SCqQbgpEDtqGqR1WThFQYkSmbFSnaZT4q12iSzO5
c4cLB51zDL+6cOHfHhnrZX01zQMTm3XSY5YZpOcxfCBAqdOGZGXBug2Ib0iF
SzJ3XzEChTloXs83dlmhlREoS5L6nOK5bG69rJ8d4qfBEs+4dl9teYABwEZB
6isFlHYcIS3FQWTRKzGiCZ9o2OdM+hMrjBS3rUiN+EYt+NYBnRMeAorhNPMd
+NFvxcG52Mm56Qshprp9Lq92zijyOCRYlDvNA5BKeF52lilr9kNJ/KRoXLKs
1MJHYEsS/TZLfc8Nkiou36RGluLFLdo/nu5/mIMc4iaErvc2vXChj5+u2i5f
BfSPKtpktMxf+jF2j67gYC3X065fSkEnmjiyWpKv0OmzpkytcBfddiVXzKln
HEWIQ+qNzd08cpLrvq/UzIGsqcKXpxL6chEGSK2uKftyB2fEkAdRzagWEOUi
QoGfYDMdcqj2RzEBCwr8EdB6s9YIZsfqSnTnXCXhQcUUM0YBzkYRfkRTbmwv
HSrqZz4o7qvweVjWqvgSvuJMmYzPPsfV7XYAMiEHrEgDaO2+qVjJ52W2oFMf
tRv7MiEbRplDKPscPaAqPNXey2S/qkwzZtqUIS1W4AFNTrSllnl68/FuJWou
oYJcIDke7W83F+th1qDSa647ukHfc8Vv8Sg7vHdbbAFX6KttbIZO82HLc8iv
srgeM4W3NggkCdkcD1vWOHoljcxT2xY9kFTEBs/5VJlHXIeT7bMd95QDCVoz
kPl9UMDfjYc/H6PQKP85o3dU3Ywr+tjnYc/qdp1a3XeDsQqHqcwj58r5vPUW
mgzrIui6e2gAFuGswdJfrBRTO9a2SHLZRHEh0/TiWrfxp0OnXMWMjhz+S6hs
67D29Du0qToXhjb1acCPhPHz92FGPgKE9Ca43E5FUhmfXM4BhW65UkCyr+FC
SO1z2AgyRBT3KKxa32rgorVC6tfAnzboPcGYme0kXc6UoJFzyEVNFgiN4X6R
mJy5dOGTgFR6DFQv31Vn0/jfUWaqhN3CWJTHk1akKGweGNfeXLtNc/Xk9T7B
laQGjkSKo17Gn8n7+S5uPcL38EjnfOtfZ1oyyTBdqn9DsFrRDV1NrEfIsIcX
Eh8C/6shPUIuUz28MeVPqtPZXCnIzC8RPEVKJUpksKXr3p4cifT+9KP/DuLI
u9jEeWldGi5LnXibxFtoilhmvd3TFo9mzBxv0Mv2k9EU4a1GpNX6KYzZc1GV
n/ddHh1LLLp4Hus+2H2t/vjSor0FpXRkvxZ37qraZe11AdHW85/9+T3PxGzj
nfRfibp8qdgKTt9VTUj4QXZh9FNQJieJkyXki3n/JGyCnbBKLvZSBDR8zL2p
MENkPmcCu6DYSqOqBtic0E7265t0kVWm8jj+gHyz9OdHZm5qVLEWIIU322rP
A1Kw+1ZBbP1Gsb1GctKrrb8C2/TXZ7gpcp+76nmRlYYMvlSrYGC2hB519tGF
RdzLxbL/SavpZmWTGcCYHwQMKef2ZeRVOVpo3iuucpPQkG7zoJ9rI7YZmCfx
uS4l5bdUmrIuy1j1kk/iZjJIsIwKQp6phgt0iRwdoPn1TWZinZ6FXkkC//Dv
QDoZ6MK3ZEhnzg/b/egUR1oUpSMrQLJLAtJaz+qp9dZJPdya3rIUmN8O90FZ
gcvTJWPMPqvfvUdHoYsuBcEDpfNO/6/QWqNKGp5Do1wvgY9/BwOUkO55mQvW
G9Mn2qd4QDa6OzTHVsOEC6yXOLoQcHZzxeRjMSkx96JWwaYTGgodaS4UAbJ2
obetKzlnAY9tgT48ljukVY+t7cZjLXam+AV9HpJYr05WcLRe7KTWer0fB+kM
hJmGfi4Hy/YitwpmCEeaz0GIqcWFfgBzAJ82nYuhwHE5UizSKrjq3ou5DUFb
mKx5CAz+ZePbgo4HhYFMvMmIyKE7LXIT9YcwOB+KfkMz8yPsyNPU/YFrvMLX
aTbq8vZIgxwmxoSy6b90J/cRh6reEfniFToey5jd15TNtZ11f0hYu8UO/vGB
8LOMSnmzBN1XxwMpY+/NIhi5wg+NBSTeSAn4VndnzroLpl92EhPkwPC6x28/
7E3VYtdUd9J14U/84LihcyECdOqEbvY/iDGzyNCjcswBqYlsrDTHSrXOJJbQ
1YGfn0eVv1I6fje2VnmLNI/dZbVBBXwLd2rZxxr7aEbwJ4qIa0LZ779ItgaD
C7HPzyqH0dTgU3xAVrJHHG/ZiIcaYuor7IyRE68gFY11uJ0jwR+YrmfNh+OE
k27ZrQXgFZbpLxZx8Jh39NGxv26vOq56NoMaI94j0At3TVgmGWQYC/lAa/gD
G9j3FzucvmuLHWHtKrJzBYHaJjqqLTbV8PCItVpFyqt+oz2DlhK1JU0HBsf3
E963Upz+JqLSR6wB5q3+/Sm7H84h150WM1TDshvM8lot7OXdI6PSS1FU7K7n
/H+nZA488t3O8zsmpYPO15gUA6yXHcdhGcG1ox0YhqTSjfZMDmWr0RRKsIfF
apWV6pSFjIJWTeBAdc44+2H6EEwwzPnSOm71e2l4yCPZ4NmfZJRLIfrEILBD
/UlS56D037LQyUaG0WExfcCarE/zjctMdeH7TLF0TmQckqLJ4NrvCdx8HSz3
g7MZpNj5DsXVLAbxOkbi7kLL305tIOczcvzcneHRf4UynaTtPDoxWvGrbOR6
us70IfRa10tyYifmPogwss8uS89sau6SKu+rNWihkuvPHrt5A0KPIhQ5DLh2
Utr7rm4k6Rbmf8+yTcSk2R9GAMGathg1qQ9yP6FXQSgSH6/0Y8b5b2gy19Ji
YCJxCnNrImWs03mjV/Uz6tF1u8gWThgoaE0miAhCHt6fH0jp/51CcENhvwpa
e0vU48VXNrHL+R8IcGSf6ua5/WwtjsETVKrVAQZwtAVA10RO8nwR1+ynysVn
xIpTzGO8dtJFMEqI5h+WhDzzGQWP0Pg/AMcu3Tqtura4U3vIxJZtK3Z5GIyP
SkuN8kYBvSoIQaoDaVzjgNZtg4qyF7uJzj8GrZ8GpU1WZmCI5zQKogJl6WAi
9nVIsKvtqNDwhVvVpQOspwaN4yOe3CGzMGk0lf6URPUZ0F/Ur1qG5Al43L60
CAs/zw62Wgm2Bn8JrSNfM5D4eS6AbW4TcdkArwoWMvvDrJL9fDPerhmVu0kL
C50wICE9VXXNSYHuOpssyYHObSUqdOJJpXkepiowK53zkUhmW1mJSkrtYNyy
pQ2gSe8ZO2Cdugwb0tI5Ff3LuXtXX1wDkrZRWjz+DMCGGsET22POEhS06kXq
NiyT22ioJPdblBeHZ20Z3qCCOjHvghgNKwKWkjm4i6eJRr2kMiCxda1mWJ99
mS9HTOMviMw44FEZoVk8IMBiAQNkMKFNNNL6WRv1ICgPL7+9HfDLS/65Pt00
3lF12251WcYTw8rhNbo7kFEVMIIfFHgWY+V/+X/BzAn3rS2o3rn+yMGG/sQs
F6JQkQzVZgcZ2LT6xaTyN4QKt2iA3uNumfTj2p1IHbBLjCVtHClMJxca3j3U
r4dhKpUjmEXzaGv7Tf+FJ4X5trD59GZ/+UqiUb3uRWwLM0JiUjxMXfpOdLd/
5yz23PYtqLJSDLRrOzPpSLWB8hub3RBlwrpagPJHQHQv/b93xS4jGgTTvMKK
sE9Bx2e8UICphmfAHww5XoMIfRi1FtFrO04fuSHV6Qic7s99KW20jC16JvYi
MmL8hdaIczCBSV35c4YCU3IG2VEl3bSEZ/6eOKojSlx2s8QsJ2O0cscHW8Uo
GkSv31xsFs7FV52goji04rWSXZcJkxMOT0iqw7uNEm2vNWVFL480hhMETdMk
Gy+ecVx+eFR9GC+RWPztrMA8InPJnSGyoRa86lfsAy/IreFmUqvlvo/Vs4tz
yNtwcYrUnqTaoUpkp6GH/Ft8OneQlX+h6akZA4YYYHeWzxJzxLAo+sxraXkn
MN7eMjkY2voDzEclzaFDbUX2TovWnAeUe+pLxhwAmQZWddYRetjlodMhAvh4
/p+p2tuDNdz6W9edJ4mWLZT0HJ2l9IUULKphuIG+Wm3SYZ5zDdpJ1B9jTOBF
3ZmvoHYZKVLyGMPIPovwFuxBix95kln1RraV/wt9Me98tS1F385x29i1q634
Y4kyPgp0RzvuW1QZToIjT7i43MquchD7DMfnSIWtPEJvPaBMt+WkMo2WX8dj
pG0ceNpbNwxgazx6YjBy1b9XI4lTtboT8BCMaT85cS5I6go0Ou2aXZQ3t8S+
W8qtQKdRZ0hDZYOKZSj51bI3C2ihZIMqLr9EGd7tBn3uzfxkAMhTm/lGsRx/
Ww5DxfGkZkGSn9J1yOAfICS/SgIiIIQblNyrh0C22fbmRmID+45lTAM6honY
O4gXPSQdSGYowd06p1myz2yJTn3Twg7ZaQgby2gks0TK3uE0ipag3GGh67Zx
o32kmQY+t/mf0hheMjoorn7qJq7KatqO/Uq4nr0+nvuHhX9Moxws42PybFbT
Jp0t9SjUcKLvF1UCvUmp1EZRZgi5/t/2ZhVqb12uOq0MDUgjzZ4K3S4yM0PG
UEDLisCJuEg7pZcW4Ruc3SutIAo5R1qE6V3zSIRl/zCbiSy1vYuoNh9n47l4
8MPvjetXf4YIFgNLmg2ubUKXTvstKCjDy8SA+ElFPuySocc20q761+ykf9Vs
FZErUuJIjAyHlFunV00V+uI88ZfdZvVQFfh/Q0V+cnDESUd0cLnhvHCoarE4
Idl1g2XfQUjj2r9mQYMgD2yWSDXdNHx518MxHUCICAooQ+xmAR69UqOKeUm1
QHjMWiRz3BYC/yDeL4GbOiMMOeYL/R5/ybzKQtnLQBwjGaa5yTicDZWmJxnW
FOC0YD6f6rA6ns+nQXtoGylBdmQDkDqgJFjabtj4wFlbzC0KrrKNMRvxH309
7/zvZFNdD/sVVHzB/JxA4BgAbFnu3+WLJpFLa+Mj/thKnrFrVWdRM42oZnK5
Z22LMYzvpNTJew/7HSJvNDtI23ZgdOM3tATbQGDwRPnxuw+9Ne2lqFMHh9th
e7G8JQ8od1EjHy6n7qVvJmNVsY0B7rNqJoVAFEnQ11LOgIHNlBPAfoe0awa3
gyXZUxWk/5Qg0eEA4skBIe44xTS5zeCeLK+L07Bzxct5CB/5ksZYS610ZbIc
m3D+3V2rxIc0VUW+NgwKUEw5z/VCQ1t9TCi5b60uGpmm/kRZLIbdIYtaMdJc
ENC5mtknUY2wIwcFjaoUb4IsTmOYYAPCwuslRLMFCK8wCpKjyHJ30ozd6ELQ
ndAhR5Y3jHxHiAHCB6qRgOTyVhaeTCzngGA4LhShJ4XVQ4hwlw+9fGQ0nZPl
ZLiEwtK6mRlxByDPicA0yhl4ZPg7aWIE4CJr0ChyJOsMwJp97/qCUzB7994D
IHT6VS5C7VAHgyMMEmML3WX4i5hT5Ycqp9nsd+3+5XXFBCrBsuA8k1P5FZEY
es8oASx9aLJB11ZooYcARialgCQUm/uB7utNrYKSr3aZDHZgpUxkBJie9JxW
MQMlRjRfWO8YZ3EONl7ErDbl3mb1321Pgah1xS+VNztR0uDvwUlrhVw3a6hc
jw7VGh9kRoJWL2+5TKwKShr4AKor23a6+R1Ya7hSPHZ9KKJQ82BGmHJAkCD7
gEko3jYdM9ndidvm/xW+iw1lD3ElE3ydRLvRfpY8XhnCDT5/ozDVno5GyRCN
kBjyDWGypLbgXOwde7DPBU2DdgKUzt79te8xTga9F7ioo2L1wbeLqUTl6LRv
t0xd/LV63WTKAzZdUqWlXxlDLgepC0OW9lDPc8DxIT2uuZYYdJcvMENsoYie
HSi6VACl60e/Y90Zpz/OcZVcW7xjaQtF6272jadC23o7i6OiS/TMj0cv5q75
T4PCJpEl5t0TIRhNkKBXcwV5kfslTxRdHpQDNr1RyUhCIdzamtVRvsp5tWBy
7RIXFhEWJ7sl85Tn1z0EEABjRoxHfs6yHI4Lbxrc2ot5bkeIbotp9VuBTucM
rHDiHMKftIhEu8nircv06Ji7/bOjlFOWf7IDTSFQzMzD9SPgInzImrA7T1yF
9Yv0qxIM0gUZIeEcTu/ZIjgFqm7o0t4EgKbyLII75I23hn1K82ffMJVafF3k
rNtLhjfhkjjEnBlZ09vhfzI0zWaA8jQOHASWsesb+YWtKDP4cPzbPYjcuAX3
DfUBuOKGtV7ecBhxpEqQCXTrR3U4x/9g7XxFGKqFzeA2rm9h8To3VIV8y56n
FUqIcv+SEcGHVJgQ8HBqQaGn9Blv7vSy3kE0yL9zDNJSJ9dHfRkrsw114qyp
iUX53PeMhS7XcEugbWpJx6Wmd/i2IpAbg7X7YHcbzhPVvfWWDMkAloPiL5fX
ERWNPO4noVrlDTVQeCUEdluzUWTb5iHjoJ+rMycPAEElVjVvwqsqFaH9tG3b
Mm6zFNlAY3MVN7l7xuueXFzPuGaPd6ZejzfzOFHFH5SGGexYqZA/Nt1Yvu8o
GMBl8GSbJos55Tn/X09kFgirpHZCzRiRSggBHdXUkfY9ahnhNR75bmwmJJs5
tPtzMIM6Mt2/7c/fivn8L0MwPEJDXMrVeTtqfkm//8XRHB0/j9kXbv2sT1iX
TpqaHPjrEg+oI1wEUZbZAFWmMCdXqatA/QekTBuoCvLoYv/9vAgw6e3W0O3a
+D6f6qKfT6OJBfkZKrKIdZpIOjpP0hlEYfig8Rds14klnlFcmgorJDlQN6rc
GvWsc7qSWVNp5Z/Mhvlum6kkemdhMxlFWdVe9EZzF/+82KcC6iAOX1S3leP1
ABPRyerDOBsDN++rwfbyb/M7WZ9rKLLiXowj6LEdCtR+pe7+UIfYgaSChSw9
izeom3TL3qq7vhAzqhFjKH9DObppA/vuORx9+wIVX3Dp7K8Ki+iM3GkJQmDd
401y9jnEOmK45VpX+F1vejwhuKMI7Xb8+2ig2LqwfkZ99WmHYMOvZKqcqemR
cszfN6SIT0vKlpjruzOanu1TdaLimMEbJyLo6BRIPB0z3dioBWZqYwUfEclZ
FtVAody4FmU5ttT+DAYuF40W1tJjFomqNwaXZtGwVcMnWVnTFi04osrSDL1t
1QkwigZgHe27n9AIsvQu3hfj+UJIHt1OrJASKjwPb0q5ffaKFgn4Nj0zHUL9
Qv5AYODHnqBjZvR9R91qvG1+BPYwKzg8XRhck1fLHM68bZ3MX1a52xRiYWZt
Iq57WTmDly7sFjJ+r6Otf63h3iAVRsByDvYetEX/Ck0U5ABhbTXVMYKXJbTz
M5j0m4UeBkED1m26DpLX0d7deV4a3DCFliTDAzi/oOZUq5Kt24LP0ilVc2Jl
V0/UMg36ywLCtbSQeWQ9HaFagt3hgkPzQ1tzqTf4114ZcKpUvMFyMEsEPbbU
Ed3DIb6k2krIeUDAjP/Zr5pH5LiVy0MuCdoGgmUZnyj/2xfHbWg4iWU5JE2v
YNuaSUk0SzSylQTbYTXoVQSiyeZXqFAifqbtu/jSVM3KHoc/9hVHA2aLqMzi
GxZKbnk0wApWE71sUc6Ynv5zDgsosyKIBK6jv1THKpVAm+bsE8Qs0tLOkuK1
a4WJbgysjIVazZzZ4SI4HDa9mY/NF4Hfm+MfCUkcVUf8YYn0mdOzcTg1PPib
TfRCxf8CJrjIia5KoQbhiYBXEtw9P1WCcHU6BaH63L0NR8TWHJUF0fikJUN4
vrtVQRgT5JtlOo0H8FcTlYnOB0ffXj1lm1p+yxAlnmvMnlCtBgTxd4z6gt9U
Bf1NU7j12YlLW/vfyTfRQ1PEhyVW2mAKhxxbM3wT5Lkhds1R66cbxO8eiPKC
fEiBAmJmww7gUVI7CSM0zj7zGjU8JJ/eZ0PXkd32Wue5BmHO3CtG98psCZRf
4jmcX/QjcFfhMM8lNQTc8CEwxu+9A6X9D76rQUU6dcZ21EZbUE9loRSXIonI
JpDs+6PxV5pLRo6LW68ASlCegAd6DCQbE7rZzctI4WdVHTNqV4C7Hjv+8kuV
HY0WrxFCXWbyMbrl2AZS6C299W3mkX+mUZPy83KqAxTr9bglDAA4JXa7dx6K
x0f772yJsrf5yU1p7mTXiB6cxDGU9lL//EaWVSZdFXu6GdFnAv8jAAUSl7CR
aEV79FjKobyFgDt2G9XyKlEyhnIQZhU3Vkcat49GcCZYC1l+Sys9bFcRk7H8
YFsrdJnbDgQx6nPOlEiFR9Qz7SzxHgGJWtUz9WHcLGmSsbM7V/lvxk/WV+5S
uuUa8Zc014L+rAXDqFmvHUqYNdMkDjs4osruS/BADr6V9uD/L8cs7TQ/hGaP
N073fpFho+dr1Gd2YYk6H3naJNWoHfuyMVJAyl0v+RZ3yKWkcHfFu+EB3rdm
Ftx/nyGmzYOcPPg1meWiVr/KuhcaSb9fre2H49jwShTIBqCShI8uG89oN+qL
55XrFB2yE88hubEQcMXMy+qYgexxGyNpfNxTgTZSlfFFV4T3bjhuYdTMX1q6
+fAn2esbospCpPVDhGSlec36nBWOvooxbZwlx9mkHvSmiTSNo/nmUN2Z3r+r
i4uTzVXqCyzhxv4AbinIvnR7pDgogJgriFxSiGen2TGgOyb8VhhepeIfAveb
sCfUwjuMFIyMD9iF/5TmMETfbhQmV9aLCk3dciEeo+QvEKBZ9JqH5agbc4Si
QN2J9E7/KSuGygjy3UTLqwnrfoij/80TtZduHdpU5g42Vu2rYjSvYLiigy0f
3AwlbKp5QZfzTou01sML4MGbxlPTlzfa7WYPmluVQfmvSJY5dB53aVNGZeHc
jEd8MkGKEuVNUZ4x9g+MMUatZZTeAtLai6jl2kn40GHXVxm48ww9la16ULKl
NUqNHDovuIHx3nJrcxil+GcjSnWEmG7S7SKrcUQqbMoBmrLWjIiTMixWkThd
SStlf8RDyZvNb8pJU1q+pO/NedZap6hsNBR+SooAJs18AdZX57aB7plWiKdF
hh6ZVdc31YlTJKykUfU5BimUwKfmMS18IE+dtLraCeRn7jjeLlS8sk92x0Bm
eGIYableF0u/iF9/+vPl/1jFPM4I5gwsbN4KGiwlqCND5/MD3hyXi68kMbsW
afh5NqI4ZRTGWRQOuxGF3VZ3KpaMBb6RYQIPPqxYg3gKSJo6dPpBHB4c5bbX
2WWoPLg/FmUxo4bTuGQ1H4rduD4/I5pSD+cGzSu3STLbrIx9/5c6dIiG5d0q
EVfThKO0NOKpzBN9ty62lSo6bbsAq+arFRLXLhymeESQbVNwQ5yKv7b7vc/G
0wAYpk3FHYMCCH1+fjNolUUDI4hTPwJatDTUKrKJNs9P63YmH2ASzbGHwag/
sB8PMvayt8MSsv9lwKraD+iL/v+DKm+Xs51AFQDf1iaqp2XupSdAOV3KnXOy
g7BrW/k40Ddk8C6QGXNHR21byL9xG2QMy9Kb2ZldGdgzOdFpceK3+YRfOReu
J3p3JUTYffWXb6CdoQfgVfK67rIiAlR6XvGx/+UQenaEuteEgyMcNyUWG8Rg
RUePNO6BzLXQ1dKl+TAL0PsugA08FMzQeo9d28/7A2oL9SqQx+WZ5NC5ghMM
iAX/Nr6/3kfLoL6rqZkEXaU4N6izTvOypb61eTLiMlmjWowckHa7rkE1Oo1p
KexzBSTVeObx0u1+wI/KMGA31Us6k2l6XXToYFW8rDWshtzqlk6Gp/5aNdHS
5cnIlKQtxtuavl94VuzbxrAAOTtvKvSUaet/Ewzdkoy2/avASCNAz8cDFo5A
O5Og2B7kHXs64oxil3GC64PRk+Ouv4xjPrZ/Ucc9npA+wyYcSARomFgSjrEj
52ey28oSgybYN+JADBT2TigIkpOs1zeo9v5B3HOcxYZ/BMoVlcDJIotJyFWW
2TJhBMnG2IPqu5YvOLmB+Stc1/9MdEnvM2GhEdjAzbB1XuG1A3rFwpUUobYS
uY2koFXn8zvJe3Er2NfgQByyv4BvxNCkuuc40ClLmLWmspv0KCYVUiF5jgzm
zykt/hY5erMk3Mm74KWMVhhF1qDGf+pBOl0pbI4JFGHCFSURWCYILufmSTkv
xW6Em1kwNBy/rjoMveuYSw9TXLJZcfOa5LHLE7QBOn96mQCh5MU+8Et2NVgB
1UChA1VLn8N6qblkTfwPKCd96LVmLrVTUbQ9jwu0Dy+M039Z8fWzOYARPSMg
l2csWb+7HGpJkI3K//HSlJKXuKuwqNBpCtHEjWy8JjYmR/Yx+2LTHwBxoY1L
WYiP/m52AiLdVcJetD7zBqiFOaI0y+W0eEk8rG8PzOB3mbjQ1X0ANxHF10pC
fAltpJ6q7nSDksltsj8gwunEwWdL3SNc6zrFD2FKOp1UvUT9A6Aw4lqpKj6I
AWhIENCflpshvzhXHDxZOeect7Wki25gZyZmw+3FuwJS0nEQrRNtBcdoICRv
uP+jaiTa3guu8B4DrA/d/zmn6bljd5R97xhZ7unmQ8MH4g3NkF5v9/UVKEaM
ZjMWeNIkqkAucn1b5USyuaDRlKgOXIKIW0/0xWVCpw7YFpV0x/Fze5m0tqvl
o9aMMYUlQF+RJIzbp9C3zX5HeI24nck6sfr3lPD3TpW6YGyH+2xSNlsT1Xmp
N48wiOu77mg4kosjzM+7/kOdbBJPu/lw/bCQJ00tHe1DtEyHzqNQ8RxbEkor
zeGiLi118bkPrXjnz96Pj8KEIEc/cWpCrVJOViT/12uD9LN1UZ7wA4G8tKhP
WxvYFt/9mawfLyRP7n6+AfOLeGjKRaAhttBgh32J72fRE2opFKDLiHKQwUL/
XShfatEyBcqp25fZrQVo1Rzz2a/7Tf9AfAuxABm2LffdxkXbnLq0PHmqmxFd
h9LFPVLzKr3zyAHfIltJb4jd5mC8xzbiGXX3VMlSjhbdnPcmpQm0TsY3lR64
wtgAYBdI3ro71zEiUVmX/2E7CY3JkfPYWdioka7CJgT1LXYC2lzjCM3o951F
fcBvxJL2lrDqh/UQFrCRZZ/k9NxlPiuh5zyHSTMi7pDarg3FQoCFMbPiDWh4
GzlNI0diwcsaVTMOYXhL+V0wkGUFNz/abQeUh2HciT95UpoeF9JSVmzjo+Da
29bAFVZwYF6XsYEuieQtiuny8ygzF+86Bql7zhQ9xch6NLyQ32rTK08IH272
NoLki/qDG/2ypz5cPlj8pKKWHZIqOkHFn5FhIeNSUP/iLrkeIem04yk+A+GL
jqzqHkNjkkRHKQjSIIk4ZSFfStpxhaKTiE+atCRT6JK90cH8bVptMx1N2fFN
XVCKKKGwhUmsRbo23H9NAp291/Bs47fWueyjVlCREyftyql9Uof7QPluzq2Q
GIpONZ26iaQ9VgZGMv5THtviozp3J96JZis2wvQZCvkXwhGkcpnFawqMM91G
ZgsdXToa8JojbK4eQNCEZo6D1vD9db1PtIorFZiuPJ1omYgyCuhwU3v4zxBh
xUkgFb0KTpulK4gmA9NDDfl9aksgKpV7uzwLH+ejZHy99filBrVU589vKkdm
wNsi/2B4twOtx2UaBKq998D1m7lT54xnjtOcyjrtxkiV5YN2GqNTOEQxDm5Z
8UlznUxobbcn7WIv5u3cMCEGTv6PANxuFIPvswKzkllXhdKy3lVfaxPi5dO5
OUwhvFVvZQPh+ZZU/exXVM6LArQzDlzfXSMJCtC6XtBz3E/YiLdmbym6vmUq
3hxEA5/+TDoxnApd/wJWyMTkVnG649IQyC+mzsoYtf3dZlXmkhk3rk9g0+r3
EPO1ZetxMmKqMAwcxa5oeQC975UjFhIaXfTO+P7lNrI0gfC2l6GjNjHmQL5g
WjybivBTMhWTcw1D3nUoq/Z1Bj5rWcSC9wYSQ83+xufquQCm9egd2hwedh15
CY3+OoOUE1Ao/JDG3yOKD1ypTsPy1ogWsOWr1wveserYBF7lvUrNo+2DJaDC
9wUNLPi2g9ftvxF0oolFqBKZiGAs3J8nVu63SpHrFgzmxS2SxgIfOPHcSSkD
Hha8esP3DDw6zymxQt9t9TqvJpcDHslv565+uoGPyb5KxZy6h8+PQ+oqQMyO
JzsLnKqiDbDmdIppJ3YCCfRwxt2bnmS+GWelI/yIqiAH2SVMX9JBkhfbQzzn
NSsEI1krC31Tm3eJdzuA6WvSHiqfq4sAAEH+pYiMmMS7eidBzBjfzoYuXnir
yg2Rf5b11LizRJDj3u12jK0WyHDzxHBJ8vd3DZk1klHzPLRPca5b8nXsusdo
OFRtrmD/AlrMNdXbIBGaOUuk71MHeHwa6XyuRMOT7zuNwasVBxYGmkW8Tw1L
yNmrY+lSPo0fbmzusEGycNKrUXZFNsgGeciSpha84rhSyqfcBSqr4KQpHCsn
TOcqXT7xfdg5yWaE4q2Pti4ZYSYKke1BkWlSG9g3quXuS8x4rkfO/Dfiv4Sx
/7c0fzKDAVN3/pD10Qi0+gR5hY17Sks0FiZSO9U5EYmPt8DUiWZmc2qKnzwd
zN7LWI1Mbk9w/tib3O8/uaJUAA8QgW4uP1iwj2X9fjmL8/7COiVFvXZjvKn9
digxCvBHwgfaAp+U8EHvx3/8HXA/CJb6RFjHRsYlN7Yo69Yr3lYNZd7VIYXY
K+0e8UnlTFIRZvFiCzuht+Ihd7YKFRzqOshvmSYRqJMdkRd3Nt0oSv++bqWh
EBCweqX9++nML4FQzC/b/fFYvH19H/PR9C7sY1dg5fFjWm9hBDVcNxvWiOvA
V6RhU9Z60HNQWnDgrusWrgx5NcrnLCRWhmRkG3OYcsW758Adxj2xTRmWk7nP
79/jlFxzZdk4C0S48d95N1nQ8asEAR25S4b+Ke2zti9gEBRW+K6hJrpKNhFo
nyvj5RjP6xr9ifGFS89YT5AyST7T1P59k9vlgIqs0oXOLH4zprZz41RDCqhI
q/5u8uglQmFJdLJy4JW36z44uO+H+A5v7wGfZZHqYO9OfWY9izb04/I6fjfO
7tb7q+JelpKe0R4pzDInoIk5PLofO5WQnt8QDdz7XiLC6Zqajc4X5x7Co+sc
DPPkn/kMdPXbqvFsr/Lw0tO/p7bsaFJN4SEWdEgISp7s9hX4OuahDCSD8gbo
w4o+UtEADFneXyaH3g8GOCurmgVBP+3U7rRafz1hNSAKz7m+L74ttGBoFeVL
JqiEFOwoutA+eq5kJGiAIktWNStQes3yR8UM8ZqDziDmf9w6VfSh3dO06vSL
UL+U/FW1yackrIpDVHyafzukcVzCByvp0M38cyAsDKzjvUIN1KwO962iiXLm
eH/EI2qgELpbT8mMIPTiu3nyySJNE8Lq4XVR6653D6gUfCk+x83q72Zewe8s
YirFoplwwrQEPj4SaExsgWjJCjCTSBbCJGCl5MApqTMgpJszlLBf24qSgXhJ
Qbl34VoUvlNRLYZCul9qzLmz0tJBPAJyic5bSN+oUrM3+sbUrEN+93tc03Tp
Wabc7TreYJATbejzb2Sq+ZWoE89EGFgvhXkrKs4uw36Ir8qdY3zir1bpSzQ3
/E+K9CsaEN/jZKdL/Eam3K9RptEYLZlFwM6KVkHsQH/yM9J7qwTbUoPfbyu4
H+JEZwnSL08HYeMMGrVN9wT0OVGtyRO/iumlbo+ga+wG5prCtX/U5fBShgql
MKCII4xG8eJPszXt88UjaXmbrufq63ynSjp9FSbWnf8TIo6pq0D5x5QBDUeh
kGD/AnNcUyCegNfyORKc8KglS1cys+B7/V5Yow/Iz4TlD8dvqXntjF4ERxXR
pUZVL7TDwJuEioXNAe2zazTu+q3LmLk/sIi0ozG4zGEf5zDNKOIWz3HSt//i
WKeUKg84obxXNmKx1CWM/AC5Z28T+T02Lkc6zKe8IpSswiHZsCMLzWGLGPmN
bYoNyWozgN7fHOs5V9DdwZJcgeDVveL972nzhRtsxxJu+wMN3lK++2jKLf7j
97LbRHQiQxdJErvSZDfC3Q0inHA2fnca2TKJVl0na8lsvvLeTPJEEkbwA1Ti
QFYzBSFn6qfBYtROVzzO+a63UplFiEb47bp/mpHfDmwgcPwWnyouJWPRuTcu
1GYXvM+PbstxSYSbNX2MOg1U6AFd1EqQl10YQu4MhIE4Q3imCHZJRqxVScHa
jflXOoCasmVjIWvEiHH7F4v+1QZUpQMAt2s/uyJrwwT+Rw/TAxwMIq3N7chm
rutvPSSwTGh96Q67UxqFU5/l7/oabk9narWlQnl7R9MgGU8Hjq7vNgkoXCpk
5pQNJeS3TQO31RHOINIiPxxZKVFAvLcR67oKv/rx6koKXwOL3LpA59B9MyKb
MfMsAte/JthcIL/9n5Gdj9k5vEYR/p2Y3gs6NHwKBtvH9u4PAEY6OFnuk+Jy
RaFPzTCrQPGhE55E3I5fnDUirVFlqQXj62Zub6++7mUQGGapv8mw6WnFef8J
lxf1VSg1pjX+MiT5hh+eYPRByYBFEqie0vAgbOKDUICO5iLENnBh2pEnJylt
mv5NyoUnhe05XNXuS+lZrcVy1Ro2MKF3wSMcEFX5iRjdZuaMdaFwt5NfC+ga
Ljz5H3SBv4ttjxThuWkWz2Btn8xPXLk7IJ+WBRPg5ttT25pzr+94F6foFELg
drAQmEgrieIxq9i2kLbHerfGcX48+u08gkhsdo5YhA/W5Uu1/AE78XSzLVCn
sMCA94oCCJHfOHRQ0RabW14TAvQ3KHfOYwOUg8rOo85dQVkl1VB5NnmcfUdc
0ES6M9VAhocGN7Kvbp3EMiofCcbZQz7Ff56OM7lfGrKVARqT9zjVyR3cZX5q
QWPTLAcfVbqHyyfP+gvA2jv1If6JtAL177GPbN2Ywo70IcvaYSEKWu0S7ukI
iwHi6gT6EuoxCFQyzuEVDPx+J3z/nRgqabBW8JB7dMA5idEC5ibIfRG26PCB
W25vG8deraFXFCP4e5TXzGuq+KBfSErwCiw9gyg2ppeCw1gomyafd6gNaFCo
xjs2bd4xSAi8SppBBAKrdphyU77KujFnGytuQGoQf/xEyscQQJcKGhP43oOQ
pW16W4Z4PKKDX2EavbJNF6OuM0BG6OYayrhRVVChLaUXhjRo2Qll8oolm7R4
EM0hn6NaEr6BT71UzHumMJtPyN49cVXZ49YxxUbu0xvuDuOP1DaEx8TpF8Yd
2BBj617TrnHOhykUO6Xg8a9Upi5AWWbISFBB2d53ewJ3eodOAbVClZWgzNbY
Ns15R+uFZypwDQ+c7UKJ2X8DBp0dVO2ObiknL+UEVi5jf1fP1hBDqA25UheK
63gq4zvhnfbSMb2VKljyAN4uv+WiPaXUJppPVyVCi7EXiEu/xED2BkdKFi8Y
/RCDo/bbRDvEA0/19Xsjmf0YjGxx6NlUux35v0FbNVv6gCpPOKjirAecNi8h
/GApJxvweMOkDIjxzDTklIAwkzXoTJ2zIfNmteyf/V997eQQ/+MrQm8sO3JH
KbPDCRF3jFq0Vv2CqwRifaDzHPdThlOzh8Su7B4+/UjfgRg9gE8MO10rfuz+
gBW9S5DEfYnWs8N0uGrzRw4kFll9QWuiM6Ie0TtHZxY3ELu40E6fhWPX+CYW
KvOgQq3F2iX9fZzkgHz9yHLAczqCsPShnO99yJ9OOI/wSU6oRDwOwvrgx1Xp
zvBRJIod0m+b7EMpUPktz6ZDgBbqDneP7ANRUw4z59DzT1coUABCkHAmaixK
CrDQSbgEUJQ/fYMV27iCzIVBFiHniqwqXfVg8qtCMC6/NvlX10munI3Xn24T
44owblgwy2F7CSF3swL2QGiKRYGYQmvOzPf2FA5jBUGcEOQY3ti+cvwML3Vh
+Ri84Wpzav+LVuQwF7av9GENXAgHHtkYBZWAwvezY58BSUbPaLQqnBZlUZEK
eMKuKJnk3leNNP761l0D1TUyt0w4dR8dZQEuDVj1k3eMoXOePXfy0ocP/kgt
08VPVmZcBVJS66X53+cE15U5sIjma515cOLyHK6lGtpbZnxTd3fV11bIYqju
tVehjAlxvYJYIhvYbigMouNr/xg793xXY2IcmCRJoZKw6w49oBWsWke2h78I
wPtEZUkV5BzeB4SnWZuZ59lf7lyXhr31FJAPzLAxHknMGVc3hfIL4g4MtajA
QGb0rPBZndIjkrmtVkNFq0t1GBNxszSyJVwZNS0AO+lfcd5xw3oKubzJ8QMS
M0SwRAOkcLJmGgxCFSQngX77uvJh5HXWq33C2HLrkK+HbEoUxRIe5yUnoiRZ
hKUjedxuV+QtxnIjPPgXtMKxwC53uHNoACHac3ZjWTNaChuop63llm+xSEbS
G2RheO0nFlyRJ4of942isH+S0tCqJIaIDunJ4W8SmDBBJqSKH7ZVteZUi1aP
bNKKOk22Q/4IZqm75IwFHkuJJi9Obc6mPAJMQKZ+aVpEnpbVYJhxgn5Iapnh
EW6Qsdw9GVRloUHh7+hhjH/luYII0bsltow0BaIe/jr/USvBp/k4Yv9GFT6w
c0wSCuPEGytqc7ybkSsNYJQHTmuRhQr9iuZNqG5KwP07Mso/E/REjxoFUysB
lvgiEwSemtm5Fzac8E456IqNrcFDLaeJG+Er0AvbmoaWEC5tvQ7yhB6eM0w9
VJqNWNEWIP8XVw7zGQMompWCwv9etWLIBtaGsmzQ9+cK/4iECrPkDr/ttH4z
Ohk3qXa4siXjeLCowSvoY6ZA3312rEfZs5MgnWe8zHUnx3LoyW3JXcp39GbU
156JZQDJ42o//ZQaI2NYrfKghEC4mVUBffHG0kZK4zpJxmZMCwMoHdHB+QUH
9nPyc9h8Rx6ZiWaVeHe5m7KJMDRBdmbU5Jm7o0DnVos1o3AjZXao2CAS8Ght
gTPJSnA4C/Lb5UP1ZjyDnAS0B8aWCVWnwqnWTgMPDA7x+swUunAFHxYHNA5r
bsvCMZvsi1MXn5SrZwrcEA2qBspyZ73SOnPIyUNqAe7pie3wIWhAzr6rQv0F
E1OirC4JosIWxGnmedPhYYAojWRB7pwWf223k8avlXrS6dDSNE8C+JRE60YX
PlWNMBliDk2RriLngsDXFxQn7qgUrC5cBw11pM8VaFLB7pCnh0TpbQb257/Q
Mb31jiYYUO4ghKK6d+ZAx+mnDT5Z7aeFoUSZxtK3VD8T+nf25wytQ+3J5l+C
BqtktbXzrmCIWTaI6ErOgcrSrZMWkovof7EjyztOw6OCwYpShgiYr4UH0adm
vD23wxgq7jwFfLlg+kFmFkTZ1MNUkhqXWsF1S8vh0mxF4CJd2TWON7/Q54cM
xBpQ+VXzjUzszfcI6OO+e19y9LLxpIvtiALUehaMtANkBDNQlUj9685VsoyK
f2zvca/hgl9CsKf1Aj3daZIei5+xXITP5znwjcT2YcQvfR14v0xq8nbgDlWG
Lse8t5whI34qGkaa0mKtN7L8dbgmywT/gpK2R7EpTCO5gzK7S0IkPR6bvb9X
MzwIFLC52aMX0ixHuo7ixPbJxXgMJawGPutjnlwsqf7Y8Kz4mwxAZLqI65Xn
5hZoqAw2crHUwVL8cXViSWaJRos79wQx11n1Ha5SgxToZYVRisd/CwNtB66z
2q60VS2AaGssMm/YmiomyZl5HpiTWNAoC6rsWuTzpkgULV+rkkUs0kLsPtTA
6+PZxJlouzqpTRfacWXteyOlJ3ExmEHaWqTa8thvsvva1VxpL+HNkVP/gvHo
+l+0JYAJWtO2fDVL56wagkK+oNi4lqEUwqoveVHiyQ2bQKXt93r5rQA76MEx
QuNk+b/Ti9dCEp1ogOrSt8OrWvCGdALA3tT0Ibu5x7P6uWPoAbAVb1tg3owU
Ewq769gvxAcW8tK38VR/BHBTHuxEbkrcVMjBCSz5XmnkNWVXK7L13WbzcnmT
UDHxgVoUZpZ7VH0tJQOCbNVtikXmlOSqwI1qS6t5A6Fe60GEnjeIruDHZYIY
f9mTU3nWN/ZZGpJj3nlB6ROXGWozFbMFmkzt/SdhCPVi1GQWbvs6OsfU0RNE
hfeuTI++Exh+OScVFwXXL7Ay5QAtV4yPyxrtDGLpDMtsoJuG9+L7yvdMx2ra
qlEC8cRXDu5tFZYmy9OP/Kt93Xe9jgiDJA7wcTNoucl6HAXtABlj5o4srUV6
Z/F8yVRFcZsrPTy2E/2GBd0lWKsCd/RVPpmuP+r/TSZfH7OJ0AQIPA7d11iz
uLTABfLAB170gibP5Q+ygCMuLkoQab37V1oaFUxi9ta00148KlM47jZlouIY
a+aUsAeqVb2ujA7cqZRmkpkux5/7czsoFs/bcZP1ZnQNLyJSQVYjCXkRZrda
c8jXslvNxeLR6OVzSSZyRvTFGev1swTDQup41vyprmHwZOSyOHmPvlLH6wwR
+uYtO4h/CpZzROj8qeRaKyglFDxzZ/omhVdoLvsiaZ3sWvA41RTAjlpl+7+h
cfc4w7ERvTNuYdR3j+Qdi2/DWyET2NDNZmz27oVCc/bCNHU73wN3xGRJIZuA
x/TXWIKwpUJ4uMGsmYkEVLzwLl+ckq7qHO5d5VcAtcznltuqMdjYglzxXGcn
j5Jx6qpdzc3ix2ATmKYPj7R1X8d8hBl9o4mbJLYLAp9460Ni+pFHKGi7C8nk
FglA3RIB/fhGN0slP9ctBEQFaOU5QrGWVsgSnLO52u+uOX2YU/3duus3hx1R
qZ3xMmZeMGBFa99FEpwjzcOEmSMgfufN+yUAVtCjXnNES36wp00XQoZOg4uS
iEeDEibVkHPw3ChXJtjNFyNd8D2ZRgN4KGooS+mPNk4eSoVJ13uLHRl824HW
x2QedzwFkXoZAUW7N3EWJ4qA7lDI7i6aTg2/LelS9INtcCCVM5PFeiiee+/v
I/JPnnwfgLvQL8wQD9/PHFBLbpmN4bd2DwBxYbbn+XycDALOVvWmWy2rMoit
v3yO/n4WCK5+/xVklYGM6gC0E6SwgaiHWOVtEWRYz9LOAilYBeEAbOhmmgcd
Rs2Lh+MtNsrAeCKnRrQ+NFihr9UID6QNTysyibV7h53DYOh9merRDPOlpmyE
Vv16n8zdcveT+BfHHHhPRjFoXPhU53G9i/WZv5ZP8SEhn/P0v2b8XaPPpWSk
5rRJN3vWnoN36cZITI8mCEbfd0yJWerba/o3dMkBcT1tlZx34FwVfLfpDaf1
0v5lBgS3onOtCH1rnrqTTKloZA4aJ8LXPDhjgmITNl29W/L/CTI/BsQF0e30
Rb1KyiNEcUxWx4ilOAk1y7WwM4cK1xxY9s+MSprzfMuhDELkpX460GmtIQPf
NXrzZRT++aO3mRtL/jngnf57vPCLENAmTHcDlB0xdNrInCo3G7m0yiElZDeP
dcn19UZ9EnnIKxQWKOXcI4YXmplqajvWL75Udng4+9UhMKZUg16iUTw2pGdY
eAC1hpXeT8s9aDrpjgm4huTM3h3Bz7ooeVE0adXFZihyNt4etMZPokh/hC54
Hy3n8ZefUjYfCJmDSkTsKbV0yBIrB8J7DtbaLudVS0wzAYWW2m0ouYXIoZr4
mrkT53+S0i0owOH9DBhfSKmDqzUfJyswqyFRS0lSR4yWEgGsIdLuHyjo+FyN
XkIxRP5DwgyxdY08rxngRIbhYgojdZRtMx5rO7DLZ462xx8NyVu+zW3C3Etv
LOwqMbglCJ6Wp2usnI4iek9UjDYFcjxMwwFLqtBQd/iRMZ1oy1nd4LhCbkIG
C7AFAMK8mWI1AH/mTKwIw1eNOvKPJ07s5U2nDv9fwkpYY6+SGsku7WS4sgtD
a3NZaK34mnpGFDrGYglCeELTxqSQrG0prCIsDlsd8xJaiBDzuFr+29ITitZ4
kTUmM1lHQAjBpHC01/Kp43Ffd1FeUAOSZHQqw/NoQSepc60GHnLFAGPmzb7j
zG7jGOyt7BQeLIvIKTrok8sg1HQYozHv/anwkNgVZ+jdA6l7Q2hmQv4WM4/I
/vC62nNMSKcZA9Sz+tAVi0q/GTdg79mEBh0j/Ox4/JpwjsiWV7Ou618gr6uw
CVFfvxXD4Ury8gs1nl67dHDYxYMAixzLfw+wvnxhwbGEo06+6Pcj0GJXH6wi
bY6n956ap0POR9ugAw6daCOqit6m9kI5R08t2s1/uzqIDeNqrXmlC9gF/700
/26d0cgJD4XyOsqnt2bEO7MGBxemnWtUK2sqTGCLfwIxJi9DCpda5/Yo8siB
2zGhcE54Ijttb2YomuaF/46mMsqNn7y74PUrMFIMLn40r0OIP/+Uz5ao8l/R
JocBH8NqKzR+T8ixXzfUnlVBCo/r7ixivlCppUOwmyZBUxyS+JH5QQHVLwqb
XTgdvKOi137oYsLqQhFdGur1YVj8b70HG6nSaw9CBQ+Fw+BuuPz4gFdamQkb
CnxQSAGvpQpplNgffyBEAtScm+/sqqg1aNvk4BBC+KnlmWRTGulz4ipyBQtY
8md/dDrnJ3zqDFdNW4Opo9ePyOPJjMz3Ygq2HAI9R/8HL50ZSW4z7RQ6rPub
nNrKSXv2kVDSyJfGkkq71Ks7unQSPzJV1fvxtaCVFxdCXzIbfRKv+YOQ7LXQ
m4Z9ePcitIdjo2QYP/egghT4IU99CvQFhMnmcb2CxvQuGFPI7qI/0EJC645i
fYzyqfwhJoS1CbDoLXtCQx0Ozvu1nPWWAfv7KNFGc1cEBxDvCYy0S9tUk2ls
IlCSlIhDPAks/8o0X6fyWmpu1A6tTZqzNOPrkrliGaZ1ZMtxUjnBf4Mpw4z6
1k3AmfnTd2M8v5L3ArgquEhzwezAzDqdeZu5847iKa/8cBBw5ErYzehKyGvz
y591LK3Wfk+TWgbyAm6bJHHQ72NvbGi1ErZVvBw7o9oocOkAdj8e0OuGMt1H
BMZyQmrM+RFg4YzePiDfgaa6Sg7o9j0tqXWdYk9RnkPDy+s3H9pmYhdfLG8m
nvi8I3FXjm6j8m9qNroCyK7PGC0KnV0jlnlVwn0NGYkkzD/vTXmrSYEpWLlj
LReWneEh69JUECdiTwpBTidJs59wrdwya1sJ+LiGweq5xd7ov3I6HWPvTVda
wqERi5dw5hm8U4QvaP9afdCLk1vLnglbYl8qUxjJ37U5eoGl+blAanJ80E6E
s678zuxXlcDhPTJPKkOu0YBoloU/MLSLqIMqYDlTkdbCaCO1j0ohy9xc+/GC
mITFoGZTqVOyqlp36pKM4Rd17n12Q//xZO6zAC+0b+3xEqb+dP83r06QosX/
nVjX4taqoAgc5Z+h3xVSIS55kvwbCyIaRC2rCbQeiGhO9dSiArCpG780l6Li
UPll91idIARyXZOtcC4kPQh9hwZ5kEtCp8OiTArY2ikuiI+mCZCSdbgCn/Cx
ssuolskdN9XgIQjcDUHtJK+qpka31DIu0Ls5QMjrV0s39swttKXLetqArDlZ
hurfr4QL3lxxUn8S7lmmuETUBh+onujVUELmYcQEcw++tjkYSOsoA2eVATR1
h3A4i3HwbLv7383mQ8tsfFqESHQFinulAeSU/ID7WPAQ6HqaQvEmry2P6yNk
/TtLAejDfzadZ5rNHUOdMeNDzn0GNn9uR4QEAVWJr7yhBijjLLgz20DYHeOy
cZuN8+YtkcbLxIe6pjttxTBU1sKkJZVRKTefMRYMVq/1pk4mZD/l6bfkE4jV
BB+kWHl/zNNUeTlJ+DOsL8pt0yvYj8H/2n9dG6dABraZLTW7VmyXNhBvvFxk
7R3YMNHKEk8jltWW3y6eI34WarhQaAYGcDHfUBji6EMmK/Je1Hln425m4NU0
IeRcoGPhVOrweRHUINmsHdo3fghmxJ4ZKP22cHfcE2x/tgsG3p1yJuT67P3a
Kw54TfcxwIqqeJ13bR6aG5DWhusvpwmumkGjShzPC0U4UrRDFUPujvPf/2zT
dyXN6JtscF3daWzZmmmJtqINymBsoc1twmFtutrIy+dge6Z4iUBZQth0a396
wZTC7IYTAdDJGiLNqdIbUwGjxnmANYhH1IwEf3fN4XHKkNHXaktCYuONpoV6
uYuLqNGKdZSGPLtd7hgB9d0n0CwDjSLk46OtsvN2/5zR7WDU2L3wdpr4Sedh
rKkVCMt3whrOPkYEjabAvoHyMiLeKyqyznxbnkvfvHvsfJWXzcUOYgk+042a
7HYKEhf2MhQ83tGybuB16CP8+KhX5xV7y5DzlSFM5Qghz5CbOHHhf7NqPRIl
rGRV417Fzt2OTDk6kXMulVfNsZ/Z/vSvKvS+a8oh58EJkgY6xsUWG7sdCMgw
+VZCLRgg+wNv4z6b3mrVbJaJjgfQLkf5+6pq2GNuQZ/prWLIK0EAunPdVysM
kfzD4vfwjdO8vxdA+osZDEU77x5CPo1u18ot28pM7qs2c6eGElqM8avCjR21
7smSsWOKbXQddlWimAGabd4gZ4awBSbCgZ3M4j6boeBjSn8aAu1RylUz/n5r
Pce+LFKQxJ8kiZRaaSs+zBGR147A7vs8K40BUw3oDDnbdVg6ScAKleqGAk2y
xPY75dbP6VWIbtQiRMsUnctUfPEdNotK62Y1mUlgWIAhLi9N/BjdWLUZ4wrS
j2kG93Fxtc7OYavCEjkB/+yf7UYCB4FJXIj2I0xKx3JfsdT3i2MzvgAeSd4d
6bn7UBm+hhJxUtHsV7Shb1bPulrnTn1uuNnLQno7DveehTqdiJM7A24xhxEv
1vLNDy2DKkMCuNhUWR0K1yeFDOWNga8sDaxgbbHmjRCQbpD+NpQ/kvAX6C6y
3OEdDoI47nT1gDiVJFKw+L+0aaV/VCjtRdSF2f1RiyXvWHgVDrBp+tidkoTI
DBNpZ8XxsHv7PR2QvPQZdYCb06UiBbZY90wCc97XrXDsOeqDva9L7+RiPfvq
xeXyGQNLm3uZ19Tkpox0HAq/Lzmf4VLTWlRQ0kyaFRJ/Arx6pFwo9CvHd20F
bNeP4g/K0OH0+uZcVkGqvila66BHnQJtUfLThhVO0rxSUieYcawsGQBXutl/
1j8AH4+0fxSkKcTxEfWukfWahv0R6xZnqCxsRpQI1FYSNDNZI5/Vh36ZT+XY
vFzjwrLwsYsInqDoTunHJS/acJju1BvA8QUdT07jjmhmEopfz3pPVGMGoPl7
HwPV2s95W71e3oE6n4Ba0qp45UDiCaA8uifVo7bPSWLCdKSROzyTX5TArF7l
v7pGsjHgQAlEqOzfYkPTwR3/zqUl1YX3djSot/p0Wmq/ZqGwXWE+PAoiyYd8
m7gbDxO90PyOmLz60TeOQm1Sej3A7+ecDwRA4zjKjUp69blgorsFKW/IYN82
3ZWF7+mlanvfWq8NFIFiUduXmR0xObi4UZbf0KNNGK7lxzFrNcHfAo6vmsT4
jzWu/fMxzFh8PEx/Vkc1HhA17wfRa2FM21xYdyDAmueXV1vtoNugcI8HLtFo
gRKmaDnKO9TGDPaUHuk6GDED3e6Dxer1yak1JVf7VtVMoIEhn/YsEQJiqICb
tozWbdiGGiHRJaOIdWZiqBK5TFcuEbn40xQM65ODyhhNqGqdDHpdX7YlS4pb
v12nKbcQV6I7IZzRPspsOp6lDVgYcfRElUaylcXj84Dmvw/a0VMlHK5WAKQd
ofXJkFsL6VbCnlBekw1hM+aRRxgPUllAxsjHwJgdEWWfNnSHn3XTaAZeOB4B
BigbZFBTT5OZikCn3HCZ6vug0BeNGyHDH71sVl86lIRHwoCTlb4Ar75cGl7l
Ur4Dfyg6MsViITPDjanpildLsgGJV1HM+9mbs5IaKnYYsqrnY7qpTdORyzvy
nQN52p6CYiNOHmStiYQ19uw+qJDH7/nAH1DDmuENqt/2dbO4sldQcKgTLtT+
5CgocPNNQuU7PmqmUoJNCMDkqyMyufKNVNgfO4Am5S/DFd6g+lx4SGqG+EDw
0m1Dlb7wD549oX5sumCp42QYtyzLlkxOkKCP3KHHMrgiHxrUUNsf491FLL+H
++lXNWdHyiUV4Kz0G4SMdOdNLairI3MCa/5/nkUuySXytgNbVqvHladABESM
YZp01XyINRFikS2whzSQ8aHf1UTyomT1Ihqc3BxPzrfwGZx6GoNSnH84cpHp
b1Zi0QHG4z3ljdsg5uFDE9gBnaI0dWN8sG+4EIkAG+TUXkOloQG/Y4NOFwKl
TLtuVHrjipwiQ6gTerJwKyaCdZKfb/F6tYGxb+9dKFlMCHiS9RhZQXTHeSq4
qpt62NodFAXTyT2T8NKKQiblgG81rOZIsufG2GsxQCHFM/lhw2Pe/tXFRX86
e0wysnn89HTpSQNK9fxElX8fC06sXFgLMIylhvaTs+ZCLRXPkgEu5JDmcQIl
4z1qDMfbojybxrP8DKG7LFD7+LEZ9vmXs0espd5qkl7WxLAr09CS2drERxWm
RzwJtLiiKeVCfdDTBSCBf4EXPu0MEg/r48W5DW4lPYXbipU0BXD3jB/2HnPC
BIGkJ7+DV9x/poCM+tEJOTBIDJ7W9cZ9wgI7H9SSDb2+82Fov5S22CaFb/Ku
fzsJOdtnhpPwgbMMQEk/PJ5BlwArVsSVUnjV8T6KInRVtKaCcwNNP8t/S+iq
Ir7EUYsV4SF4PGOQWMaZmCoMDLzTiYKB4RCOUwZfyv+UwhaJ5TOkvuawL0aG
dnj8a6P5ti9i4J8odeI90v7p/1FTN9SX5EOq6IbK4KFCVJ9ymAG9fV4hzTGC
ffAUG7MGvznlljriA1Fz60RMMuJrrm4ZGkcj1vAv6Q58JO+xWQqjzV32LTl2
dlbwS0ADf6+pQj6n8OOqj68elc0q1HJRDN5MvKoOMjNcMSvWI6Ub24R+ERu6
l2DFgq4zY1W+/IjousZuCc643c1yy3F6N00mRYMDIGLi26+elj7y5B6ZmiCZ
/ANebjxvXK1y6XFpB/p77hWJPaFJcuAgKlKbeAPw5XHgJzjVgxAACv14akYn
pjCRZn/mH2r60L7Z+jLNzArKRKyiYqpSgiaeydZr1mGSSSYilVPxwfHAHoFF
2QUx39Y8yHoVDG0HOYRIrHqE/YQV8l1Lcfllelye/cnFJQxPEqgp9yUrGF8q
AboOgMbCrcpVBz1HBsnz5JLjYDiqEuNZibppsXZvkU5Plrh2QeKAMp1UGIEL
wehTzTE5YPz6WiXq/J1WSa05v6pUZlWm40E1o1K6dM7tR1eDhy0TzEmL7blL
shJuLiHFWxZm5l8lrrXmRXfQPeMULlN3ayvIvE8XGs37u96cs+xfycprhAeZ
hrq5jMcRcVYDQXmPsL3oeY2EQm4hLq4CeWvuq1a95pv/ve4Groewq+crxYSr
VDmQQZ9zmcqJ+mizbI8VfTKRPaxtq6lXhvpismomF51pfTIiNZJ0jUwvBL+M
wRCyImlbQUr3TdPQqaqtHGC2J2V1vPjuHPgWDC0wi1+HweOOo2RhdVuP/t3m
PCU05WzdlWVjJ3oehZ4O6QLCSjDaknHzfypaYCcKr+T8JByUlNfnMKOLLOLB
GW1M4UsVVkHPGIMyULrO9k4EFuhjQ33+EIEb97D3UcLQnw9aR7/6FlZpTggq
vsVVLUbAUf+ZzpB0DALVVhNB9hHa9+LtmmsMKSr9jdP+nGTCj1s6UVHUqHpQ
JrWPYEUTBR7Yfl5vuQiu3GjJrrLPUgtwJe0E/oODfZeDCM4lay8apnnIaGsE
TewAXUOw7AKrL/o236kp67jQ6TAfTuvzm4pkBQ5akkl+bCsefRFbbY6R2Zdg
N6717j3QQn+tQ72wEYQJ4Fa61ssfju1Xcq+4FZHnRXpngpz6O3SRyvZ5qCZj
rwftZW0pFUSuM5tiagAfsmZhQy5hVry2GKfQkSHVmddZGH/5cE/v3ei85ZON
lKykZSPmyypJfxv5dyU9sj6s7QruWacENcLbt/vyWdudpDeAjWTdx1tbapsH
Uxy4YPntiLlG75HqpzZTVQ70fF0ZrIyfl4aHa4TZqbv4IShmuc5PsLNqzSFQ
/0EmLRyGqkT2fwvs/wi4jeyjjlCYbxQDZEcRaTP6KwAb8CD3idrMvqQPN5y2
Tqnmd9CbxMmeH3vtpwk6WSmAJZ08Cxl+3+iW+TPT/7M1XcYdIr4kI0A9UaF9
0x35jqstFASLPVwkJ3MW13sV5eDnMUbkmEjDB0wEWOAc8yNQb97HucQGgmzv
bYhfpsh/jSMXecGqi9fLFy1D4cmkOJCe7VS7zhDU8l9XKpDWHkitHMSf3PlZ
Hyj63Wkda7H8Mp6RjKq1mLn8B7QjCIqGY/fDt2e1gVBFh69zN8/FuRwByafX
S9beYNFfbtXxZ2KXxINRGk3/dTQldxV6HKnxV6b4GsKWXPBB5s9A0kwQcv4W
bNY58ZQTZoYOhWjXarzREFESTFV3Ij1mBdYtATdbx7PqJG9Vok2iRkcUJA80
jU8a4VGHqFRVlYLJEmv49h3dQeQ81ksTNmv4AxlyhfYmH9HVOMbeHIdW9w/j
gerFQitl/JcJh0XthuNG5xH5VVPZLaufvXHBQAOwm6J8zoWH+k013En6YiPG
A8eusURp7H08O6PwKqZMe41AnCYT15Z7qYmZ5o5ZtxZkIML4pMRTOOD5R/OZ
ncl+dHuNbnVECeQB+iEBz+ZbaMCBW2cgqerYcmuOM/7GHd5fWo+XTYs/ooaN
FnE5mZ+/r/1tNiEfx8FMxszh7umzmtwJrfd/1JmKKMW2IQVk9DDiVNxH/MIC
kEvOl570254ld7tBVwuRnQl5f+bqGjDrZq48MQ8q6kA//hTaaLQ1QphxT3bp
Z2r+2nk+mPJoX3kn+Pd2nC7y9UcGLLcmB+zSEhGGK/Lbmz6mmiDRGcsG/6RD
LCZB5A1/2b3Ca2BDcrvSVTNUt4h4FABiZj3NPyVRRZn//gKRnHXLaOIrXh1w
D/ZqVXZEoABHdhlxZZuAqsdsn37L0EwQWKzXjxjtiT1BK7E/TYjxC+SzvN/9
nKmQz/d+XZ42Jp2XhhIOjNn3cU5BusvxPrqIJynUmeIvShpAbgQy7h5kMbFS
pExtri49Ti4rJAuBtwepn1UqHFicqlbEZM1wMV7Okf4IC531pmEmbPSyjBZ8
HGkHSpM0xIeL9MdL9GB/SOl2CQArM9Ta06DoKvPd5Q9jER/DUcum3gi0mkoS
ykBpL8K57Khhf9mjrINf7CdeRqPFTINqhzGI/ObYGOSbiYJkxRRcYPv0KE/Z
5jq2W1A49I1LyPc1nVIM27XWqKJ7lzJaOMexCYNp/EstWkCXzhwk3U0M+cqF
b8sEzqexr0Z50+EjnptyUlPVmoo2uQF1NO6/srYdjrrRSJI+YMM24Gu5/Uoa
tLx3/Z+zab0pkV6j6aTSHMyEfhNcmf/eFokhiDziVEHEq2l0VifxRKCKT41h
cCdaCil5/+fCmqCrm+xzdciOYOxK4NiU+dpX0E60wsvbqhHCEf5R5hNd4Mi5
NKvbfMCuc4+lx/rG94VOvY3T12/AIG39vm5TX3W36pC16mabqdYXJy3Lk1q9
RwnzwU/c9aSe6OxQKU3npe5I+oCVFF3U/RSlqqOZGnLeVnfopCgHK7FMf84r
E33DbTKYR+BhfURvHb5lPqn+7iQiNZzQx23Ht6DC2a09+SLIKFpByTzrLqeJ
lTIPNARhY8q0YBoxYcb3mDVk3lM3ZKAZ7xzyT0m8JGL0mOug8NxoTUOuJFXb
5M13AETrMctWLPZ88gGApPwA+GKVRDCMFZq/90OMlK2ZfuwH58oPed3+chnu
Now9BnNi7k8VDmY/hXCNhlvXNtlDg8naNjrkrMH4i4e7YEHjHQvNx9VK7rAl
dYMsWfuFIXGdXhNnxh4SvIafCtBT4O9XNlKvzdKfUnRLHDrIp7JzadakoLau
MdQl6/b6V4ocJSnUsiRam3aASSiS76sOuwuz9HaT9rW+JTrhPBh0A41cnyhi
VnR7GCozn7FXFA59mkuJTTROGzmKO6jBEVuwoay2rpliPYbQuxrQOktgmxdJ
Iy7EpekDtamDtLV/p0aXO4MgN5zd/25bZVaZDTZSYZr/TgXsDwizd2+1GxuX
9Ly0sBtPQPkVITvAt5mQLI5w7NQOGB0S/IIjvgmlBM8elcctobnkLCf5+5sD
Kpdg2nYchzKkOVbzRCHuqAkcFETKmv6cdFzz/G+33p237HwjyJ1DMisp9IvR
l6FUwpaSNOSJPzJNoS+Vx/nlP+oq11MspCnzYi8wDioEtx4a0it0toEpt9IB
N84s+J8QuNVtQX+32g4wf6SNRaw/oUWZR/kFAUX71wGBftnSyHAtoOdTERd6
6HzEV9ZfoFJCXnQwH+ZI79cEw4kZPtKOjAm7nNNlJJirHH01aksyOBw6VqFR
mFDdspGcpPRr+UmzFIGFnOV3cY+hZfQpuELseyg+93uOUciudTXbZNV5UN1x
OCqKTelGsNF59I6ToL4A2mzdXw4ldO7X7sEWbyVwyOZ1/b/rjO/WbPrxi9Qq
Heqcqrxh+x9eakHqtdAURO0K5cbBFZ50F3VfK7O6P2mHMgSbCeFskWGyINod
NmuRu7+y0Weh/p7vVWV2z90kB5750LGcWcKSdRtBUvN6/zXRyh/Gusi/bKi0
yP9BNZRxdVaBnnXXQpfccKlc5S0Y+TQ/0O2U4OZOfcV960Lc/qWMG3vh57sK
t2LyykqYkTK0iKablryh4ePi/6cQiFTlxo9aIPIcfXyUsctSzagweEo8RoID
aiIXekfyPzcHuQZlARodJlt8XFWPRz7L1E6PRb6fOQYbBVanUUwsHu3uHScI
eDctcc9lxkILwr/QaXosb7fD9yj+fhEq/IUn9D8DrrCu5mQcVsr6XieaxJVV
fwGAA7OrOr8/Oz8G6GL3P53lChS2AsvgTsU6wQo+iZ1pV5enS8Zs2JSdfyKu
rsK/bnXe75XKn5Rsh/pXyGjNrJavVb8zui+8MEsiTwathWG681JNR8KxMRih
QhxN8jrSSDeYUEIOobmvw5pvYMzZqmem0qt1WDFZS7A2vOweEdtPQ4IvgdQf
umvc7m0pBrCuTXK5aqXdQkn38L/3EBOEUF+3vzRHso2ztQH7sDai6wdwwINE
5+pJnhV5u5Q7jhm0dKEHWuJhygLiw05te/fIq9x2B7x9ffB/+Jk5+j6C3Ge1
bFSWxrN7V/OIZs7P5KZM2zeErdLPX9AhN+mQR9vuCmktmTSCWpltBR2iyQiM
bdQI/PjQ8vurYo8S80+oyu3CyQr53SRQPODWaJnWAqQKlmGiMzlaPBN1m2P8
OtsnpJnOrCGVy4539ukvy/aWWTjhvUcXXgOXBp5t2dT8p6HwY18lGyMhmk2f
ph9CgA3cdhI2etN1O35yh/tSoZ/7JooDueoxi9uLKGAN3NspTpLqX4nmjmI3
JDClkI38TTbdX6ByIaax5dhkSAlRs1At3a/WFpFkwBNFYGwFzqbWpq5U2w94
wu+qVIbfCUtgRjkOeosvwy137UyPTj3kcmQbaGibu43qDuhJQVfFBKFLeOsp
rUgx/9XV7q+cgpJXmttvJ646dCuttja7ESIfTE0egXrW3kScyboSd/+4vWqk
zsEkJhFZEGiJ6ayGcRxYOypi8c0E981ol8kGcOJtkKZErk+QY46HTED9Mw9R
bR+n+0KCUxDFdfATM27NtxmgV45GXbcwxFqCWT/U7khhycjKNoUVYQIOVF4T
hTjFQlpiIsjSVLi7553kwx4G3HOd7aexjlJYP/MUsOlEp6UXEgqhCuKw4PCW
+XxiH0Oak+rNOBXOrOq3jCKSOL4R1Pq7EnOQkn7uPwjhNHqlOGH6wtM8VGwd
mfrJbjb9jLPOZw6fX3BgObO9AHb87NDRkC3tM5ti41hhfbr2dlFiFD94QHGi
PbRlgTR0KgC8FY5WF8b0d2B4OkfVk8reUmx8nd8rw+/jrdLiUaTCVBdTRA0e
h1QWLcc+jx58ihq40tGnYF9/q9D8EDFyFuWqnSAX6gojElQuozMHw6Zmv0wF
C09pqkLtf5H8WIvdQtUGOPFmdK8ULdKb6g4Ho8RRtAPtHjlwoIrRSs+PwWZO
LcxLKY/lrCYFDVVFJ1wYnpDFw/dTaEdpJsz78ifY2P5Qpm2x/XUcjc2p1vg4
dkPB7S4Gvi/q4w2FLgiB+bQ+BdARbG4c/+B/XJsi3RjrrcvIQs3W/da0vnTl
FRw6ZBf4+NmRtxWjJz1WbYP/mQ7ukDq2i5umlDk7++8PNOcdeN4wXlsVFmVY
tC+96ATATSw8QqZxGLj5qQBee6/0yuQ3t93vtnHg8v2VPTaf0KiwmMLBd23E
AsBPXijG6rtv8W3zzXpbblNV9tyTV7cVnNp6ZRFop8VOTqIQnXiUr/D/ZyMr
/ms1OEONq0Bvnu6bOh6C663H8go/uskfrCztmvmSeN1a1OeYt/QA1cRMahdl
lAAkqBrBWC2hSH1JyeOtweWeFHGkNvQiFvJozTnXzeL0T/DlgpHKs5tBOa5e
6uEfbqY34RkCTCHpIuWqSeECwJ6+WPbo10430lmA6rzdI5uOh0dldg/YqlTx
KF5S7Q6q+a6x+kG9b2GlEUBVGXwGp/utIHOxlbbEz5dgAX/zEleM3JKMqmZ6
PsfWJVskoF0S9QfL/z56PGYHDgMYcedbOA4G6n5OgoQnD/kA3knfHzU8g+jw
13WxAU/XrgdnD2NHJLdK+mwyHExmqHQe3okLy9q2+5zTDSh86271g//nLtvR
4c5+DQVRMNzGNGwtA6BdRnVNFNHsEzE6pgdGtdw/1N0FrWWsAqYYmG+huO1Z
miVPRR7KbyYRAJRHek96Ng8AsBjMOICOIdKm8OxlYX6wnFkod9x4wfYZYhgD
STmjPmSbZ41RohNhfCjUYGk7D3I0iq5qerFZrk3gU5jaT5Z6BRie7IIgmYVW
06w5cSq+UODUpTy3bmDwALtX+/0zP0pQ+hX24ufw8Diz1v7wVBbnEB+Cq7V8
+bi6QqFDuhQnuZ1H+cWBX/MCAkENkuRCjurCCoL8BEIoEb8U1LvzKA16c+Ye
zeiNs9Q30/qd2aRr0yxk9oHXei/gxd1Oa2Ae4M5fUimJCGhg38jHOU10TJPV
rpgEohiLFVfkO16pPWtNyX1ZA04bh0DJic0Lq09s9lX6hL61B9KzLEFvPi9c
VTeBEUr0+2V+mgv6HPSu+LfZ4jwtmSIc8ckVMMj22epAooW/E6DFZTZcU7cR
yNm1NC1aQY/QuVHSCm6so/Xz5K0sLqq7+dpVI4vilsGDp5/+6V4pRoNTXHym
X1xKmAS06peMLR6psbSO07UbiHdFgfmOGQsDt6YB/SI+AcQMXaMWIodmn24Y
ATvTyjwYwcLjz/PZ7O5JGFPAXHdJ+AInCgRTJj+XXEfcqiRxDgDSyfsik7ph
8hX2Loy3MN1Vo3ws8UZ08IE3QIy4+T03QAnewCpWbkn0CPHKTgjNL2fVkUAd
74qxHd3RBMOdi2vmcEV9iNrYoYbnjZcGEOWpD2C4KJk0ABM+++oP3SnGoY0l
kQAnScODkkk3TtYSDxtKhf+a4VGa3FTIimARMLhjGjz7ZS+i/6DrXNOfhkx4
BBYf2ZdzCa2H76qeRMZ06nK03064DyfJDTis/7tb3W7XujeTXgasmSNJZH+B
HcNW2zvWpJEElgClbj3q62rJr3IMXP0w/DBTrZa5gxh1JLke7t1tbTVAkYqM
PBPynSZyJJP8Bq9y9LC44m8StsBZBotLz14yDV+K7djN6y5zvlzJHMdk/IX6
pxPf+irwtx+/DUzuKK33IPXxzAvcJ7BB8LXI7dyLYGzXdEjSKj71+G4HuKXg
Yqcgv73CnPruakCecdImjTlFyMJUtEkKj09r7hR5fymboatMrgpGlEjGDNAy
SkvgW1XkI4dgstkeXc3zGeBAiODngCp/r9FoUtBuyXeokIW1ZCp7WzG83yc2
WLNaJCutSYQpStmuLZOWhObO6vBzlpKtJrttRDM5G1xcq1ON8UjLGs5CVDIv
OrWjXtxtyZtAPjFle8Oy97ERsI+La1LpJsWYCd4nKhmUrEto3vog/iack3+n
XlL5AHuwZ8fXl3RpXPSrqnlFowrH6ZDYxiLKs3Vl/9zzpNZjTiArb8dUQXKU
CxZNDsH/xBpsvk/r8PAajv7Z9jpPmzpx2fsJsjea3t5x8bWCLKDvj+lNNO8O
amv0Cyrs2v2dbEXiRHg3ybOJq1LGwStT1f6ca1MfrN8FHrmTsfbA4WIH8OrB
egLgbwX/g/EtVuL9wdnbRYYi3vIKHkVjCs2dr5igE//1g11KN9r88ndo18pn
05C4X12S//7r+RbKJrS0kvjV06nA2snuQifuJLxPLRjRmSvtOv2kPv+ImdtX
w2KTvpRSGULgSi9dVEwVyLCWG/NZSlk7g/34/3k4x1kgLSVfEHJdqO1O6Gr1
KswKMxyKc7P/Vumzz6YV+SgAkasF4PFiSCKAQ7EBkKajwTF0D3r9zj7uivjo
Ur0SfQ0iAWdUZ+ZPEehN1krLB5v5k/c2sAAE0gG+Msk2RvIA+YtmYhBAygUc
RANjOpDw7psXSZPvFtsr5mkOhIHOGY1jnIJVb09mJM0XMvrs5oyigmtKmncG
f2uu3/ZbNxUSu9t2a9CTVnLiTu4LvAtjMSkVUSyNJbo4EYNNCod/O2VEPNiV
aNuS0f89m5zhrkOuxlyQPhqmmsPENlRBnX1i0cOe5gBy4nZMf09Hs+1VYdIG
jl14jWk3+X4PMVa7uLAuda426KUQs2oroSTviNWY1lfWYIYDoFpIcES8Tecj
mtPzhWKxOu4yJvr+4icuFDGQZZWEA5ZHUfi3XDglrJRf02fDlDnhI9sArEH1
ZGNa/ouNMUGjXj1tJVu8IJcpgLWGhuNzWXPWHfCa1h1GGEI0rlZmZfVE1qg0
EjAQ7E1j3djn9guxSY/YX9KibI14KOkBHzgYBOQtkhYm7V1D21Fr8Oll6wRg
i65KgBJj8r9U+dix6p5NbKjfeeJfiRrLCeo17UfGBklDfjtOIF6U6HTMSRvk
tWyqwC+8/+LPbAWWs3anXd8RwsdxSItBysAP4rvyIzVYLeADuYIcGm4TWaSW
WjsYLXWq3sMyteeQcg+yDM3+mlnWAZfhZ9I+I01erdallhVIuKGtoaH6Oesm
9nimbTJ9QlKMuVPokpKAPVCOGcYs3B0TAuEc7I6yCcyDEtSj9a5Bk/W9SvsS
97KkgzMfhTqaK32KEG/6TvdAKju0LRYH4v3Ocf91zLqdog2XeAcOitElRnK2
PCi88SMEWd6GWl2Y9RB8HTJZf/bfpX7a3KXk2pa++gFNuE9HwHKR/PQaALaf
OHCg1ojKmaC7owMSplpCNCdkHcKfk6uMXoMmI1ZIVa51X9t5yYZRlnO9Y0bv
v1FMXv6Uy6JtDzX+gGxRy2Hk9oCNekiovFGNIZchlcwqS3wmS1sEBwrscijM
jsWSjCp+YXHwlLDkh+wDfJYjXaG1G7Jw4jleI/O9p/i4eXvqwf/++jSYtaka
sPZmXrMKwYiCJO/tkYuVFzwFeGs32eH5foKDmNNg3vH6+ew/lLa3y5vTaXiK
BGRsexOJ+9lH/z3xLFxkN9FyWo8tKwp7t/hm31iWJYmDZAdRz1kcTIWf5alJ
E7UO+W318nH06PUWo9VPYZX8Q+o+OMOAkzruKK+SRNvrLfjtP9Fu0uTx6xTw
6RTh03d1KSGr6NpL3/RMMmFGRFrih4Se7BDqvF2ALi+z36qa2uaiJIb5KqnO
wPE/ypdMdvyUZme5OZAXXwd+8um1IlNiIW8uhkFOXyAKBvuHffeBZaCmqcAB
dCyHczSeL5k0MjPWEq+ss6rwAXoPqN0BaWHQW0zU44lgDuzQJCg1TxmnHQSJ
OAErFcKwbLvvpvhv85jSX/cvHnYyvN2jwiZdiMsMBm7Suy6nS8fddFej+Cjz
sJtNCRBqkdEp3QLACoHIy9JTDys1D9RasUCg1YwfqIY7jTVq82CmxDpNJv1c
wsE3xDT6wDfOHnhOZURZC3R7qGCB3H6EduJhsNAc74dN/DYDSuCkc3OoU8tQ
oraPPT+e1RMJDvUnI1S9akiRDLyYSJ57wPpljb3E5wKHsfiXlWZ5wiCzFpL1
uZZ2eHvtovctcXQevFZFo8uCSZAYVRlM5aGJ6l/PyjgcASMUrhaawObhcsRQ
EZI1ivq6vObGOtutcM47xxY51+k9t6oJYRgfvAVU2E/ULz8IurbcIA5cn20o
AvRUbFIVF4BulNw0X6UwlIFvtPtJEwRfvFx3euCl6tNUyHCUqRzrry3EO6Hb
3Z5jXKuDc8jlQexdwh306u9ZnwtZAqOZLDkwnhF7RPaZkzr2zBEen9LYQQv9
qWCG/2VWJ9RgajTtD2OXUamfB7k2XthhXx82QxzpvKbhOH9Wv2BcS33iH1u2
OKpL60KiwkYHgQBDyNDAFSJ5UC9OARtCeI7E9Wls9zYgQtlDI9ZShqOURvBh
lF6EblENTYEDKkpoLMn3bwVWNla1Cwxllq+/TunlQ4HVPOe0BFwrQBWpPX3O
SM2I8vgUvKFYvTX0CePCxdNB/bjnQvkAfAfGI2vmOy8AvftxYmo5yzD86SW3
f9cpcZwfkKBWuOJ/Bt7cjx34DCgswZ5xWy291xHDkdSw8XD8D9d/wXrlNM2/
wAsgo6rBvb6lXJsn3w0HpSI+o/1QrD9j6mcGHBXfNuXLO5cK4z7Jb68t9ZuL
CZEgDtV9SwBarq+4Qt1iw+1a3F9AITysA1r0HfPclRWZAPkGpNCenGos2B1O
zvyMYMWwMlhev/XGgvLFuHNSyaj7Y9uLXqEc4GDFVQuQSV5AI2dKGNmhO56n
9N/tcEIWmHvAkPsOn9kUY7/Za4s6iJu2OpRBcPVaDzviLs0+tY/0ihjy8VsY
bujoV8ayUlYH7s8wCFAl6aDTii0R5QHENoqqXjYhEv8rqwYR3cHYZxRU1ifd
FiDFc0olnIIBY2+dvpH2/Dw6ZLLcR7LA9vvVk1RDvU66ZKI76G6RRtc9wkf2
AATC6gyfjVA7pldoRGq29vPW4POHI2Y6Sh8AIOtfpptX8ZT+LOcpd67VA643
oH2R0NxgmJagPWqYWhxARwbDxJuadSU2PzkKPucF7Jlyxpg0CqdJ+PQbEMy+
EOqZUu4JZ9nCHe/j966CMzk8uReM0dXSOxSlmeRlAOFrhUReTnnnUck1uAUP
QUKbXxwGyYpY2xkPHcCDap2dWVMlWEpmq0u4/KpbRP2Wrcj7KoQ2fDRgDqoh
ec6LCwLGdICdBXZzX+t/jj2kHsiXXeTLTKTG7ZjgFxsrDJMSBC83j2LAfINh
jhQwDytHfRbynUaPHKZRe/tBQLIPfA/IbOFrYI2r1/UaOHGt05pyhLvlXjFm
v6LTdZ/7n9IboIKHTpcfJ9YDIsxDcdFChnVAeBa9QTCBehn07wlqW4wwDKhm
Uc4gYLRgHVq/uRu1VjCAFDMW0ZRXA9PQMafkaF1XoeSwA9E8vknoYLPnM0/5
q/LvQ04cC8v7BdBSuflwc7OivzVRykVPNMT/ZUrkHpqBi74G/BZXgS3AMtKR
6WNOlDpsHkV8GJwF4aroTwYRiATlzs2FF4DXH+fyttXkIZN0Iusm7pS+QU0k
BQMsydibTgcw7hh8co0XMHxUDn3mHyJJyR4Dlrtrg5R12hXjRlr5K43LCYw/
FB+HPe7PbI2ZMDxOmj9goPs+PJ/fwr9IEPtMoMQJsxnQF50xerdZbcRhHzmL
ewrTacEE6x7ksBsaqlVSOAMs5XhOq870kRRpARmfqQprqr7uABgBJoQWOoMb
NhCEjwnElvob/Ilty1fK7ULn7oKevoghs+OwxJiz6hYxYQC48u+DxybRKzS0
xLjvmrJ+7JV7zUslMy2X5b6vqAfirhpAH9vnZkR3KO9hZ/N6PehG0YUMQePT
kC7vayGDIxGVEuCkjcQCJiYA4dFzBxrxpIeLDBd5SDaFWeX558dlTmK8c4Ex
xHbMer/MxVVZP/0etFQrDsM7LIEh5l3Y0vNv9eAn4AQuzessgSsUsfok00mF
MNxQombavB0TtIATzqdPgtduoykxcDuNo4IuKgKt3yEqJ+MRBzgeLPSiSmSU
PI20xwYsuzT0J6/hhJZXF0m+Z9Z59A8Yallzr9Bvrw+lWwVYJK+8EbZSgVf1
G60hzPqZxUAti0XW0rvA7Kagb7PsOSgEn4zKfjRyq4BGGCVaRGzv4ncOhvBv
lf7i2oF362mb8Qo+hTZDOW/kyU94vp4l1ijaU06pNkpCNwFYRXHTV7l2KPhX
mopKDCqaQH5UWF0b74KpwY7EO2D074eLrWos88a8fbMJda8A4xG2GeG41bFG
rkPHz9MnWtiEEZWfl1VlFv7EdobitFGhS1DkQOWEWXUmAouRJI4i/pCCIzrN
GwTKSzTJz8+lp0IEMey+YrZ36eE+w9tFodyDixzJx0icx3oTbtoHN82BmMVt
YzwyfbAQdCSjbOdhrMvQOQ+b/KfY4bJ22pz7cytvkZ7tnaqSQmkZvyvmuGKb
1lpj7rLE2vfQHdtsGEq4tEcKhER9iyJzd0NVdx9sQQA0hakSSA7j3VKhWF3h
Ym/CKCd1F0UxtWUz7fOlAWG5UJocEn+l2D4WCkLYohFXLt7Pda/DJwaqch1U
QLlh9b7clxmWYVkcADphViuSU4yhNmuj0LgDTDPyCfydFdfpMr6d9TezywEX
ccguEBUr7tZkKLRhQGF6FPruLtSLetAqiq3o4KVfNelhMsmAV1JboHJyPZk9
gMom2UGqyz9Axu9HVPxWsqzAPneyd9qqG5Inp4IOTdz+M0W8fNweRHygiRmq
W9HwLSxBSidwm1obPsMFTB7x186aVQshd/P8vdU4GweOIN2AN84Iof43qp1t
mk4jVlOMh73Q6MHF3i3rw8oe2WhySWu9TO9Uuu3dV6KvR6UDApH1bLJkIXsG
ZG7h2gifgcbB9mCAdlQOZN/Cb6UFBOAAwQYBrZ/+QttapsvW3nmR3xz9QVDj
mfRIbk1Tzig+eO5kZ6a6O6ZdpDu5CzM8BN3aBVH+VBj/chlQ7UF3wGt5k9Cz
xhszMN3XSvjUJ/mNQiOoC5KJ8E20tPALPle3wwJS8pmDdQwzX+UmhvfaUXj5
ULs1vY+9rTKC7jbu5BpRoEFCARFTn3nsD4XaHy/FLzZoYMrsXl5fi9F6eDB8
bAboOjeDh6Ep/wkafH+W9S+fydJiJeRNIg8PckYsB7H4iUuSNZl5kzChlsqD
Tw3tYXKMYXaVnjz/cPpumzWXAfXcFljt1xZitShP4tdPUMzF4dB4c7QUiv5b
YDHP/xME31f6/9nA6ija/pwl7lhgXwUWCGYKFMlcKfde8huXItE4LGjD6izd
s5UniwT6BcCrdLYbkXJVnBcrMDIcMeBANdHXWpCEgU9QcZAJ6gAZTjJBpalO
ddkJB2XN83KVDKv3Igmfo6L8fNskldSDYZN8Uz5tMeSMFpgUE+vMRN24F5il
sf3U1VL1VsaLPh4gnfngGHkBh2uPNTnjjeW7UpJM8NxK/t9gNGwXc3Rgepv8
+oYB3eap7d2ynEefVeX6LeuPAGGtskznRTLIz3s4gUkE8+mLCkuB/fvB/Mld
rTmzXwSGpWR3QBKakO8zDOOwVaim/YjJ9mtAgZDoKYX863fUH0qmUt4eYo4u
MynIeecayyedWqNJgfGKwiF8TGUthaxgd8VpVGsKy1ikvvzzgqaO+ptS7TE+
w+D7m2YiRQvdtXufUle7pDemQ8cWXHrVg6ceb8RvKQkPzkETuIyrYXsj5nEE
JnNwiilbOkh/OIWjH7+/8JFC77Z41lcknu0hSaLdV0jDA7L7eKDZyn5Ooibe
dotsrgUHSb8hX/GADrvSeAHts8xnQrJNMR/EJZr+orrQqxQUEj+ig0Nc+WHJ
eNidlej8idDo0uKxXBhPuv0S9+k3b2jL3pkE/pt68RDtOeWNdRqdYCquxMJS
8Lwki7MQ/OOXexoXpy32B8tiaMMBSCK+4OUrIA+vlNq1fWjmBUudVmIpDAcr
u/PTcd753VI4/6vLwYiX73E0Odf4W5xVY6IPvO19/vnwcJQUSHcCLr9DpmmM
eydQ4bnOs/8n9NSt80F6cilDbHMVuqAelx0AIuZj0W3HJzlZnO14YtI3Chag
pwin4nStlGB7l448yUm3P9kYfFsN5V7FELqJGbF3oe6VjVdlYZi7XNq3M36k
tSgoHanK+mVTcrwJa4y+f0SXYdo/Yh+IBjsnEamTAvPangLuty0BtA6uEgW0
aLgEgTF0AykPzK/ajEBTB6eqgDwLAoA1DQnILCr1mXBy/5NhRZ97iERj4HCe
ItnEkVWpem4EeZ799fn5rZZ9vCn31Z+f4wndZ0Q182Jt3cMftn9NVdoYOdmZ
7JjAYgjxgTfjS54hLK4LwM+/+FYW7ftOguJf68MMSEWdok7Eu3+jPNY42EAJ
2JDfOmd71X97BqHTBpQaoSODXk92P57DzHFnHtG5Put7/HwfLjWchxLVLnmu
gO/JWBT031U191NpncJJW6jPt8CyqzQi8cnDC4FpAuBuazBC2njbAIN54wf2
HNX1OLowaB9w/Ls6jRPHm39v+N5yEfYCxRxxP2fEHiW2VajBGBFSyXM4oXdb
AXaJpMSTLjFWyIqhE3wmRNjgdjOvGcmbiWUCCuo+4BHtw2ts+AGx2Gt5nI4M
EIoKOUHq3PwlZwFVPM3nI8zrTmCrGDNu+GrLXbl+LjpJKHJDBF7RKB6SYLbx
XydvtC8wft0Gb+O7CT1psKC9BXujsqwTpUstZX7mhojszYSsoj1NCytFxC6E
MNW7PzdnIC/D+BAyBdlzeRDViLeryBB7crILGgsIRNRNbK+Gchib4qazOG8a
qnAf5dy9Ip6CnR2dsJOYFnXVQzV0ncLUlaGdmMcXU9iUpIm/XCB6xHAUTEZl
RX+VYxmPW6xmGqDMrOSpOSd5f1e7MGtYbx04IpdTcsPrTHts5UxLuxNM3MRS
8DN1SJI31HcEvbFmH/YxlK31HAYsDge+wkHFdKoAZUGVEyGaFtvQzySSEMVM
c0s1q0OoJ502NUGsj7UbRTKuKg0T6VNraWupLo8llRKz/8ou9nAl0vAhftzI
jVHGUZjxKD66C74VhFnUBhypO7n5fcBNgz4arMr8DspoxIQ/LWvu2dfcO/Ct
dDLcw/fP0BQqo6L2rvCwsS6LyZXGMz+Iu//LrughX81hfgMah1rafgf0a1KC
IUKatXwgRacqmTAh9/6xXHCynXqU2w5w/Jo5JbIWTIne4oCig+l83TE2kAT4
iM7MM01gof83hQlpu9tmMb6hSy+W1QK0zEeVHKkI8ktomTIehmfEIBuBOywj
lmJvumKYdEkriHPl/c5PGwOcKNUPrh4wzN2u+fZM9egY2WO8J0Aw/6ft7E4+
VXDvxDbDfLxC4Yb//5iNlcsM6bpf37kGqlytWA3/zLwwsbFYG3TjLBESim1o
NsyFEzPAD8r1h/2fIIk8j1txP00gajnLaLj0t6FeThJ3Vtmroip3HGBrwibq
nRnig+ZUwkU9uIK8bMBQ+oIUK1MH14WD4CR8ywz4F9eYVipnk3mt+ijFuFuo
jl7+M+HX1mM8E9WCpdxv+F6IxlTYedOw2AydzCY+FQln3SBd46Hf4qVB502q
Zwgm+Gy+6Gssx161FGZu3FOJhGoCHiZpV/fcg2YYAUqffj1O20Gquz29TP4K
W3oVP3HLUDSzNPfE2G0lWyDBm9LUP0fmhmCbg4gBJGZvAncCol+DvDwJJIx9
j3xiaI0hQ5aR7Ogwk5XIiPdpchdjYFmgWACaLFhL5nJjYOYq3XsF3FpT2bD5
S4tkp6+/8+gpmQ/p1Ydx437n0FD7T9PhJDHUJi0QEewUFOLMIZNKi2I/eaw9
XG6xSQcGveSFIEd7fGn3U6hJdC81VeR3Pi/e+TIfxImxuuIQ4OD2BGu8EO5B
ajtMXA+5UMXXa1hqG8Yf8Q6s9WjtS/1bMJvcls6yIyNJk0Z76PZ1orM6g4Hh
DTPOCKVNH2t1zWTekkA61LCB3UGRVmkKnoUevvSqAoXCZMdHS5YOSWx7Vz/z
u/vEa/8yk53KDsXNZvAPO6uGlLnnJmFkslJ6H4ZsGR/CXND3/xSpoN33pp/o
5R1uD65+/5eXveFm4p3BDcof0c1z29N7ECRcqvDfhWjGEoJAC2hP1s8i+QTM
F7Ggd+oXv9TjfIrIS4rU+lEq6aHzxPyvBrrQtsko2ozV1FQG/a7xmOkTOf7j
jWRSDgV3PvUVzzw1JYGdpnfrITSJndqt/f8JjvXHh+guT8fHBtTKO0y3FBPz
UjcHnmqSZRXrlL+xIxZJbgOr1UCEHN7bH6TMODQbzBgkbFZTy5sXz2MG9akW
aJVogUWdwb0aqsZUHsCacPpVtyj20XGvpHtSdzg/wytAWwEppnxvbf1HMN3y
mHI6VnxNSjnLdNQpUXgnFPQq6+ex2YsrQ607u/1HYVjp0r9AkT19Wcy79RBq
Cxcv1wd3WX8nW5aRuFiqBcgPjxcdVq3K1sFPpjQVO1U4d0NyReFanXAjwlVS
Ita0PBlOSq0EupZqVOuaqBymP+ZAcG9753hFEXwgOjhRrqBKLoXq2afpUENh
c+ejKQNMxPyWV/w+1jHt/NopcKFs5JnaSnu7v5TRPmBk6a72eB9dQ0R3XPc8
kHrkVnECpCLhq9LCegfqBJsVunTCUAy6EjNXmEDwgIdfmX57Wh2YRA5O7Zy2
2MQhKjKp4xnvnpy7yq7VhOfe0Do7I1p2B/LY/xQM4B59yGiR0QCK3W8EkiYL
ywAY5k6eNpFybh3Y5eJXLVrBX7zxpiY9sK/1q/RC7z4E0J8BXDWPuHMEz3Yq
1ZzNhWs669mRzU4H3vXDZkWNH6GSAzO/6HAyrHYUxQc7U25ai7wurKF/ipKf
hs3UCuEXjFz1B8y4KxcXnyKmc1W5CF2zKCWr422MOABygHd3Hmvrg/mrZBq7
xSg9oQjrPBrNxFu6pWHgDRbLjCVMYWfryMjEWtMWhjthDYTYPaFZlfxfT/By
/O+N/oTJ3z1bPHGAPDRxRfpurVu9VkCBcb1ES+lFVJzKJF4sU+GjmrPTKMfU
OcAvk4DgBT/ShMUay94vkFy+G/qRexIro2lJ5grSg3tTNNs0ibaKVbDxUviq
jO7benN+ETr5JEMm1I7U+oWsRiFTVhktc2JShIf2FV84MJ2oWDYxNr1yL4lj
zgWT51wWlmihPquCtsxOpv05hifq8EUDGgbEwH1IfQrsa7nfUtVC5SQfnT4B
TTQFp4Yxw+iJZWJ/QKwe/PsEd04E7RHtlBp/GeftmQ+GawABo0c7ynR2TTxp
RNK/7DyuiZ6nMuVUJ+UBPxlsHxtk+PyVV7ARi+/c63xWPENf/+F8LwEFHMyx
WODLXJlD2HLK2BpVzc1yZVLSeAjHEKYhYsX4+Jf0cYg07VJgR6clPj1L6qSQ
Lcz1kWz+1OTTNhgrHyxOfdAFTW/Qd4iPTGpg/A5JRtN0xpwclYrziU+CBuzp
/NUkczCp128dmzeqtREdEgrnJuUDUn8q9J4miv4GS8lCuzP1bLEF03OKSt+J
VL55cWRwUKYhgmcji8vujqLmVmSSe/1gWH6L9u55UhtcYdkeooQ8D4ncmg0j
zLaZDSMxJHZGSRU1DiOAZ9PfmvFd6gZrrUcaejyP4FUYozXvF/dd5HmsWDoy
8GB8i8inhqMmtOIeIqll0PyFrNY3fDcIt+XwXIRROoLLB7TXL4VyEmReFmO0
VGnc5eaMI5bp7GS0eJE2Xyr59FzNiyn2Bgm8ecjftuq7dv8fOZtTZKBur28e
tzb2wQv+YX9KIsAt5cKiGvtMoB6vae3RX+PPQxpl3Qf6soPPeJrdIQa7UBpQ
11UOaErxzjl22BGAp4aIHy41viGxeOMoDbXBRTR/Xfv18H+pd7rlG/uvA7L2
sXgzvE5pxuSJ4e7c/hnt1mNZecrirGX129EKPUxSbTifaf0U2BUU93yV5WDZ
RviAM/eM8gmvo2LYCXxIQEfx+j5TPrheV3NuX2mvbOsKKwAzjCfMWBwWpA91
JLal6mp0n9ir0CiUbr2vVpvP8+Y7iq3oEKU8HfzvTZwN2yY1vMm7EVN5U/lC
Zx7B/VxhIcB3C/eusoWqzoRrkN7Plnop9Sex+ykVjQigncy3bMqUduO9gggx
mUTwyouw6RU8Ak8PmroL2ImtOWT9OuO3ydu3t+pl/+0K4MRtFTy0WCJDdUUQ
GTjuIL27xg434Fc7QDY7ewrpLu3M6HDM+ZlurWWStaMAlfbVP+DPpCrFaI2Y
wt3Y0/5H0FWpS17Wkf7px+gen8KUeXjx9xQ8DK4ybksOqSqWjU83Lrst6kgb
jhm2YFsU2lF+VgtQNgI+g2Ixh+Ya1umHOM/cu7fwfD47sOBNxR+FFgBziXf4
b6rzp16GqVEWLNDSpaRcdRebS8JK+EM5wbSW+kti3m1CkztCnQO8QO3OZGE2
eV3KA2p/ib7V+G5g51bUuXw/ib6T0gWB0t/uT0XiSg5KqfhPh6H8JzwOu7mL
6dlHrnBeaj+EG/N6MkIhsaGUBoqqdcxDCrwE/Sz0cEvCVIIlbB5BJiWSmyLX
m8kh/+rS3tROWxCAm7f5jjGXqOsy6fHdBGI8L7aLDU3w5dtkFz7xhxn+bOHD
sKXJkQt8OvBKGzJMcMHG99CbDuETRycQS059HrfkP6o/VV9H6NHle2lPwl9n
LcEYAougqvhJQ3i1eG2ppZIa20G0edUsM0o913vJq0L6fXqAdvMNaAUHbDlJ
OKDfDQGrzyqfYYKwKA0+IXE2jgSi4PB9FZ1F6ZTTGCwpFU4OKlcVGsw/dEQU
76IakHA5/hXwb16wz+JlE/EK07KTJC1MXzZCiulJkk0X0sZUgoYFlqN9WbMG
SEftZRv8E8nP5tzL1hACHevvguwOMbygRpgwVgym073XyaVnrzCTxohXaVUT
hA2PCsaYH9BtBQ09oZe/nRGGvOgCWgL5CohxEjmc2AhC9apZ9biAPGVrmjtS
bA+063NDUN5OjkFuT36xcygDxi8MklGdCSjzhW3gW+iYxblAyO+qlpUPxiA1
qAJkNt2dQJ76qHiUEuxsFWQGwRycJuIFV1QHZXhGSsTIyfH9o+eVF1Se5jBu
53dJB0GFbSLAPvwYHe7pcQuI9v+mXpDfCg0hS3Dj3nie+psE64jX9LNUbn61
vS+uaarbMq9fdU402hKw7O3PLcGXDkraYy7AyDnU1QoV7aUJ9kK0LbD+K/Nt
VLQDC6XiyaQyHJOFcK6FOSYPlTEyjsOdrzjYpfyE4cv25RB9miERolLbcwtU
SilV8AGhmB9Zm7o66lO8QHE8kJkDM90car9W/Qzqi7fTQq6fDCBNjR7oqGdE
JeGRO78T104kepovDmc/nGrR1RlX92ecRN78xTgCqqfoX4PCDQYUpZ2aecyq
Qe7gnWeNRZCaKmQcjOu2+4sdkA5FF9KXygmQ2Pb1IpOoEwlBxCLIVYN9ZEeZ
OQkjESjmcdwUTnlxgdD8SZ4E0onUSOHjjpmDCiNTwr7ZCmJMR8sLt8NRohG+
i8C5WG1IMsEYdYApj9Wnh14VXBzLNCs8yh2W50lRHzFynW8d3kWhLs1Onqc+
4neHyVXljW9YByogu4D4mraOQGfgJD04DrsSlcTweVm6YHOHEtwyVly+oxqg
nYK0DuJn54fTys8X9rHijuaJtlJB1Js1AY66uSLKA4UkUK4kTcQAIHMWRQcA
8POee9jFmSSBoEEfsUaPAnqrooxoZYhx4lthj/mC2dqmeXknQ4Kx8gAuHGYH
3fPqOQq0kdY37SP3sIfG8HCMJbPH1IuIDe779EYze3UaUxiASWXMjIbg7Q5w
Zzc3kpI2A4kBJTl6SE3N4ai4K6l770axADu2Su/R4aN4FVfVP8e5gPq7tzyq
Hk2vWjcqfQtgmOVjaXAFuSBM86BMKV12LRhtBAhRzvz1DhKlOlFQQSE2EilW
OiOoRQrEcNJFHdxesVleMaULHhqEBEj4nQ7ZflTCbQGO/OcQmGINW9NgvRio
M6xlUe7QyTxZQMwGvArcs3fEYncd9D0NWXNEwWeURBnaMT4kWxz+LDux7vcL
3MUGl2hd7n8RNkbD3Uylg8rLXXdl+aJ9oCS4rtixqbumXVLr46VdQBIctLqV
Avs0ZyEj60eTee9FZgDvhHP1eVPR/9YOBXStYubwjROGKkd2Ucov1Q+XFUC0
bz2wgYWmFYqhfJSE2d8687opOoMT5qs+n32Znsarzz+LFUtTCNQ9pW2TPIlS
0NBBze+i12yR5oj+Y/SZYthfE3mXx/rsJvwnPNTS7lRQecQEGwN5IAPC2BYH
KpUIFaeyTgUyzQE/Rjcx5V+NZDD6XIb4DNjIIKFRXgUT3Nro55fIfSurCBo9
MJRq7Ylt9mKTOd1cYuIfi6JevIH+f3mfkZBnjfC0I19+Oeru3zwRv/MYNjev
zVHBtvQNY0Yx056LIvh0zkN4YWETSwaSWekYb+vjid71peKHxJjFr9kwGsUy
471eKOrdWf4pZ4gt0Jw7NJk6bAqGew8iFV0ojRT7o/i3ZOR3MQejDW4l5f6D
GFGQcHGjYKHxIo7b7Xgf2uKKwT20vqNZeLMF44DO+pUQG9K1GtWpMYfI50Fv
VWLNBjJWaxDglLxrPKWIPrW+6l5TCke8nWqzmGFaGsEohmpqeS99N77stLjP
Wi2z04UcTM3O98/mTxuEnWRrGv7Ad1wer3i1cAqqdc6B18tJuc7HbiuY6bkd
mLtoz6dTxJGhyPVzUo+cEHc4sdGMIQP5WyB+31vogUTFZ9Cy9uvOZ0YpqC0g
Ne/WzpWdEcugZ0jhm+megxLs0rr4RV6r2u5jjWj13DQjaY2ZXasGZR8P8kLL
hHFdax1hidAFT6JZ/bTBX4WJdTu0FiYljt88Xd4IE3/ukFMtqz1OTiGOZG7b
HpG7oKyXubvw86n5BRpaawt9ZRDDt1KgQn1ifrwT2Qi/GGTlZxM2qDSYa1/s
dOiaB91+cqSnKPMzebrUKaS/UTEp0A+m8hoLStmDK5BU5NHAWaqfE/ZhtaeV
OEyAjLWrSd7mW2ct7qoPJsIrOCLVZv0M416FAuiOCaCiNDohSS4YI6ZOcUHv
C1ELKry0RYjEK5uK2TW9tWwoBatrUBKkRZVoYtpKYr7Pc+8bh3xPEetRCk/j
kvcJ5n35Wv+PVbfog4O/yG5VoCHN8kxYgFi67FTImU2mqgF7gb4cOHwweIE0
wjTy5GtMtaVnN91n+/cnjdjsBsPREpxzxrQlpFrkBBWCYUrnc7jjCPY+G9Ay
5w2CmV34l5esby9LRMygc2et1cO6xJbajbIOSQCj+gm/1M1i2cPSldNJHPgm
HZWgp7dol3XwWKLAuqGb12pyovZnA36+qqokNjT93FrVTT96A4k2B878WzDy
Iag1Upj5Ko0FnE3wz7/659ICrvyzNCskt7gm36kyuks0VvK4dY5Dm2yKvWVR
lSABIEPLCLx0rstgBHOmHJKi3VO41BCuDondF0PqUTtBnEd3dL+sv/NAJQ34
+MIsF4o+grkPbOUP6qNdpJccIYzoAZc2lSUq7prMkczB4QgzEUYi87jksmR1
NkLJM9l8S0Xrr/ol/9ob9sqTGjyHyaoSB+ontYLRL5OCCyDJ8fjJUlmGvrFH
nateOiUNGD31UFQz+AqFaxiDLyXaU78bLPSu7ogV8Xg1qd4pqw2tZVHal9lw
Z4rRToLjJi9dq9B1uMukbk1G5RdbxMtFNakt9kFC+oFC8h2zrr+w2yicyeWn
z37+psZB1khHzfEtc93flh0q7lmqVUBI6OgZJJprZi8e0E5Snva0ty/ngD2S
Qawk0tLeiJUIS7nnMearlS/q49WB6pCCIZ+SG2Q4nhRYJHZT/YDL7r8yzI0A
6iFiIIq7D9uvWFQkoK97iDDHR5QcXCAqBluqvYGd9h5A1VI5mGitN9prJE1m
1A9QTntrfNb5vzbca1dLq+3bSePHneYFVlpAgJgROKYBF36Skm6CZyUAR0/r
9QHxmZeadhGB7b6FogVzc4PcffXIKAKmbtc9Q92Fr2xZ+DNT7MmDDn7j/vdZ
sghgvD5e8fc92FkgZeXbtnK9TbsnHKaGiPjUDMNsMJCb9vNkLf2aFTRW+Ttl
Sdvb/NqTmyfMneRbL9OoerOpN0XJsxomf7t/BWsFBOKeIAGE3fiv6RIk5nZo
9YFxRz9xY7alAtoB+ilWjye07xEnOD6kff0gQQGBrYuusDUCM1TjG0I6mqSh
wSOGLAkY69+pHW7/c9B92dVQPfyBgj71pSVKJXgRz+XBjemt6fHws5Ah4UjU
Z/PBtfTsyYftVZgL9Lr5uIhvxnNciBWq5vv6M5SkdlVH9kWxTigwP3z7QdTv
KhjgEoBz/G0RTTboQni9mNHHX9Jp5zaubVEj55flsQsBp59AnA09IorKbWBA
XqRlS7aKhfNu5iFmB3g9RZUp0eaMG3oc0YEWWAAkamAqHZA0LFSxBggL8Up9
qiKoyhc9Eh4tYiWNhx+a/sv8Jsk3mRloQGqCo9KLdKf3K6pwb/GNHNXTjxVP
dMGJEmZQEa6X532K0xwH2Qd8GXzxu++6LUhwrmI3kfd1QxRNSR52u+RirwUK
+MuaoquE+8xtUl6VI4I+lUBaoMiiluEBjhE1XjFWD3AOWwbBqDSeHCD2VUCs
gOy4+fGh/yIJiWi+1NOdr7GV1lqVptX9MKlVkef4zQL0CeMqmrNC706/GhHl
MbYkODLBtMqll2CryegCJL0JZ63PBbJu9p5zQF15iywwBpkKhIcRQysB6maJ
6nl7kTiAT3xrOETf3HyiQ0FBe/0h6JDCeG6fpdaxzcGkHUvB5rLWRKvJnlGc
fz5QW++gmAA8KQpbnGHh1lDWHr/Dj8PiPSxxN37Vix4AXbJP+AE0ueDPLwz+
+EwKpHdrcXeZxj3cowhwq8pSAO8dAOj1uSKciLLTMGrrXtxL/VQMYRDjxxOJ
MhZ5KPk3MNjhQMa6c1llPZBq+Qq6RzE7nGEFw/8u5ms7+WjgY21qZ+g4nxvp
WSwfPMGCsdF+Alq6OaMfIhjkBjClyaYpDZAzgGgwrns3oeZLKWa1q+tXNZLB
1AAj+VNwG/G/8fStBwIKik56Q0RwoCpOzp60Lx9FWX1fqv7c0ZSAM1Gm8dsf
W3H2vnxCJDWzfAbjFux3lA7Tx6iiLcsuJVqB4H3PrfswSpIcCnfLOqeH7DNH
mczlcvTQJ3sIM2XcH3sx6MYmW9GuJHhMNxKBx6tvxLjTdVfsPMySSAH1mP6T
bjX5kDSihcAHKi3E7epZXNQ8XmUwRfQjAqTAJnH4CnaiKm3y3luNX1FhWftO
IC8JFn4l7DBfeooBk6GIUsTj6LYwcUqDoTBRz+dvopt7MO1rNJ0ycpvjLQjH
Ef0Q7hoZythGKCBea3wiUDzai7Y4DGks8LmLcZFucIoMRM53VyAFayT/+W9z
mXQBfcp6kBHChDjXceGL6JzPWQcOnE6cr0+ATAia+5Rt2NeBGKN/Cmx2j5cT
ZEMJaxEOOuJKDCeH+6TL0duAT6aaOxV101ot2ls2ZpGNARxkfb9ewiPp8FZj
lZObfq67BO3c++eVqbL1nZZ/VD7U7YJZTWmpOsip9Y/InY+dMb204zKVesYq
zSUhb3AYW+YsEuzno9PYHWdB32DFxgZ3+tif1x8aEUsADbclkWozsGfHiNu7
0kZWIVGHNOo/6ldwqAleTq11uj00ahlnS770WXzkizQ3lnp195wN4PLPiabP
XH0roPzxiPfRQAx3BzKirdsb0WqGCWsSXbzU4kqZjcw0NlSYcvEPkCocVjZw
MzotQOC2r5r/NkxHhVCS+03x+K0bS1fZ1RnmH19ZqOg/t9eFFU/tNuRWSr7p
yOZK9xULhi6e8PRZ2PUJElAWH5y4S6bKjy/UACmTDTT6O+9Il182KYihq9sK
uxLfEhGu4vNx6pRHvII+DirytyDoOp+0Hr5wXM3ruMCunAyjF9h9CrQkitvb
HpP4rH7rFQxNcCQ/Q4WEUVGXnWz+QNSSWn4peC1NXDzVcdBW9yT/Ehb6cYny
L1kIqyYBf82dChRA1sgD8vo4w33qmoNGIeyp0NC3Bxi/IEwG1ROJGOm6Iq/R
Tii/xYI2EIBrLZ1ezW8Xvp6szxV80gbQ04Gc90dDjM13OtWkvqc7LIvE0q8D
u9CyPUHMtNWSdrI+dUhzaUnJiB60xNS4dM8Usn0lh52Rb0Ob3wh0E1iLzRen
HvLellS0RNkXeEfjdOjyhZ1t43JmBEBRcNkYGZJKWE1MlQBLQvriKXMU7fn+
XQ2Xz0BIs06vVJ2SlVczkH3z4qkl8M+rZEeyfYZ38XW6mkGp7fxZtTZwvK0+
ar0Jzipk4i3nX+pkSCNMTui4vWvpMn+LvoSVfBk8cRbTjAEv1ZPAiVygZcmK
vB/scNxH/fkkStbkKDQVBh2Xf0fnV3MrRD8oJu9Sta4+Gmjczjyl2xmw51v2
Q+D3bvODmymXXZvNuB265lZdevYOeR34s6dyH2CR/kLlT0ETyr2yUVCCe2zw
Pk9Pxgs/7d7DSLa4dxLyfljehAYpvEoOCWMF267acc0AIa5I1f4VG73+xBCp
bJmAZPOEkXqrs2kfdxeNyQNi0PP2c1rOiZny4bwi2YZMVj2vn/zuHQ7K1knk
+ZWuPKe4A0lz0T8zMc+AADowlpW/+0KUvVyf7y/8D3iyCgPzb2F4C+SpO/H/
VPRfZ3pp7oCw2H74SUoWyVbyKEX55wgN3iyjP5bbkQN5+FSYxG3S5ORolf6b
DJZ5xA0wm1Z4ohAfglqtG3gcIlU+0+4wOPyxtBJmut9kI+5BkXraBp74g4mZ
5WaAkIxmV9J54f8xc9KgiG6Pyd/yYkDWZo6/SqouGZxdH7bdHfFnW1rFMast
gpiR8v49ysD0PX2W9wtGOOwO9wyW7xzyhQc6HQC08FZdcJfATsRFIw60zjsO
tnuEKn+4R4g4uSGbQNBBrI1WQXXnx0liOKpKNMSRAtVOba502gtpenIkd+5a
Du9W1w+c9oEtIgiGYjprR9v4H21Z++lWqMuzG1y/sD6MICTG1ujp5rMR3KiI
+z1mMQRVXV19kY28Ugpne+fykBslXCUhU5ix8VHRLiVHsP5szTH1n7N+sPgN
2jHmiw9JIsnnI7sC0hY6MQkX92o6xAmYvtNBOC3OXaL6J4xcqp4LSF00xWKN
bgDxvB3sXbQcAiS2jRSOmujoPlmPXnSkx18FQeP1EmoIJPf5mb43mMDPcUcq
CoNBbhQt15gFrjfBuyHST5GEz7mA1uQken6OkJ0R73eUdlc4E0Itn4Vee85h
JvKrPg6QajTWy2cyBZbExHuBJMFlHeJ1TnQkG99WZX1g7XeuL9ruIXirwfg3
dvcKHfZsaqTOg7ucnuR2kk2ItKl9hhr76vsV9mQAayd5g1SiPwA243Mp5m74
enEyz5zQSa8TUG8RXDDkHrt2L0nvbwDHXXaUvE2xxpX/6PivpVdqQaXJoJsm
QlHqhtxxmOGbzrOKIpjvALQfly9p1koE931cOahPkFaAjx+7+e++Ad3XrrUk
UJgYpUSnMvfLZMDKepbqOM7oCakkDOTGPRNA/NZAUevre1RTC3ePTnU+X/Oy
WAPq3epfWPJ/ifNIevOH4OXRPEdPKt5YJA6mWdgpnWMfc8fSWUrmFNCYPdQS
6fy5ZqAPsL53OelzFUibWqY/SuXZTJEMg9szHAJ7x28Gn+pGT+x+SwnlIUNA
CLRsqGvyD43bhFi6h2YOK8dAp5Ra3R2/f1OrJs4j+blyhqdruXfxt/BR4b4t
WGvtHmzmCAXhvJHWYQVQh9F4Z6GwRlQDESzhtiUD9pnIwlORiWsUm1oP0pCJ
moaZQB16vNusnlsgeXoqX6v64TF3/q3ql8dQovozGrj71ZXotIjCvqyg1SCA
FORnffLNKymGULKSblwTe+YgdZp0DrPZgyy/2+K9+gHxSG8Fw5Kc4rRHFZUa
bs4gxfa3sYgtipT4EraZYl0rnu1VavG+295H0kF65fnR8NuMAyaB/gAXJUpV
Q4WUgKlUbl/ele5rt7JM7mgOhSqvOS/EFTbjuuHi5nAnP19az1eRcSwPgSIN
LaymlJ42im3ZI3uY15PhNd8JoH7M+R6l0sSzwVSex/Vb+CIXaMHhEttmre4l
pWcRab4YnZt2qNhM+8XYD1Ef1Hu7esxjoigVosgkIsGx/SPdOPdlPiPP+SRH
MziyS0CDlo+F0iNz0BMa9uDroR4+Fn5YlL/UptnQp4xstB+OBQ5tgzObV8Zl
amKMF7OdwkRmrB6YPkxwoNiKTnGNmvIhWmOc9ht/JqOOeLPf3Iz66AZ+GC6m
guulldKbOrEiSzYWyCQmI6qVrfEQyuZlbTWJu214ATSGk8EV7WqhuGDRvpar
qVuEJPO1UwHZiQjYoleHCTSwOjkdrpYVSx65sRTDC8+g2eSNnV1y4JcEo1T6
mKN1E7HYLQusaK1Tw/kPZWJr+9dR2j/eJdl98fIxNRpiQ0/XR97CaXfdFOtz
V2RmspjZ07mUU0ae6NO3TpRc4GLUAc7uudR2R2aEd2Lpio5OIuLdU+8GbTvb
M53P2C+gBKgNsPwtnkWRdXVs6hqk7z7MgTUw+M/E1KS0aYz4tKjQfBwELCb3
c+Sf224XYn++tsLi+5J2QjFrpDkecb0nh5cw7ht4Emxd2xdHaZfVIe3smwbB
F3P+21wYX9SfuWeFX1vdUfOfL0wp+QFo1ypnVrC10NPjG54SPPuW01/3FfGK
wtC7QtLwtbd1Y5qbicntarAisAG7pDjp6hQpd1kWO2jL1i2Y3UayeZqGO14U
yYMx0yeaTZ2afIp7+KhQ9z5RFDlwwuj+RzyY8Lx6fEZvqyFyDrV2NhjDBb2v
wcCmeQ7jiJr0wQy28EeBzdW0X3ed97yuHW8lcjOgIq23BYFpEIXSw1wvDZf/
OeAUuJ22Iwb0B2oAUbn3Eiqc8TqRunZ3s8bpGl1uYWrYCgWsH8pJtVcZWQeK
TJ+WbHAWcLpwo7Ucp2u4qms1RPod1/uFR50GK1IRaTQXo8YK7S9pxSJntqVC
V6Xmy7AAWnWlQgbOnOYvDz2vvVzPA9qmXpeJ4WUVs+rxKt7bXpwJ6fDDvNKo
6xIBmVGPe/jRpV5yO7e+XdgcZTYvHp5s/ZQqkxt6vEMIaM2D++9DvMMMR0kd
5EU3SypLedDlrTca9UStptgOUb65+Ux/08LElNT3qRImVkGD3qmSuW6y5z15
Fte4yBsyVvqMfPXDU24ryzw3RHF1iE9fRBk7bKRVmZARyKbIIequmK4uYNDn
bV9Sg3feWgcmT3faERYWbc9VxWrYBy5U9zc6oV2gesUVs0yhRcIOULgUDQNN
jtuG6mMLWRd/LazFUCXBXmyheyfjT9MROvchSihrO8lL7Ngm7kYTkeqF51W4
eH6rOeIX5mFqYSCe83byhQFSkZ02D3fGSu29ootsujpWptrbqoi6hjKYtR7Z
/hQrDCAhgs+7rFhhuTLw2lWM6VGltRORxZTGGgnQP0pxWEME5SN8/TTJp1je
Hq24u5VRpw6FbRgjfcPxJG3HzcBTfLdFXa/nCM+jxfFFO+R72efyWPmkFRud
8LQudePP3oT2KetmuMsgEiN7WlPNsXdqDQDbiUxBoiax32G5fkW3s7C74v/D
0bnaxOSjyM2XTkZEkPTMIQ5c2zg8iHGG8/v9UHgCICpJZqOwhqFMSjfRGeth
omzO2b4iBuYx0dzeafPbNPb4SzMrg+739Nbde4xSPU5RBpkEqukY9pabnNcs
DmzzwUEiqryldzkZwvb2iCutkslwoRRGaJUnLoFN9Od+/71ugUcUttaNK4sD
7cXxDkatvx2JV6xtxc75/Cmqb2KaAqUuEYYB++tSHEKqMtTIWMGE3SFT55tM
utEp4+HG2yambLIh4s+OyIbtK41dpYerNEyJa8B9+ApynxhdeNjzvl5j7MHX
H4eL4Bq0s8XBwgHOQW8zUXlCnVS0nx2dn6EcV1uHjkJzOduIlWcObQjYj+K9
7VFhm4yKsZQgy6Kheg6tS38yfOu9sgt/+6T5yaT+Glc/HNiatbqeRlTfAJBW
Y+JbO6DFgDoVeos7FV2mz3j+o6nnTIkbcjGC5lxnbj4xjM749K74S/zhYz1n
ogsUKRzMUR2oeLb3Lycmrr2PJ0YLCJFr6zPf3J6vcVD7BCBwa2gpEKkTXLS5
NWa/D9n381sr1L5FNJto9OUrHyMeCyqWunJ1q0sgrSMfilUQvI0RBSetcJd0
9vwczhfVSFtD52em0T5EmNwlCqia+rvDh6fBb2GhTgNywCCTaYG0TLJg2mNu
KvhyhNcc8E++KEB48aMJrPG2EHlb0yodceZia6/V0q0klORclTfVC0G99HLv
a6VxNrqvdTWD0EylCS4x8N9qUq7iswwpn/d6CIzHLA5KaSM/Am5si7IwUc/i
dSYN1wKSzmnflyPVZ0zalTCwRsX1EL8yqOpyJDKv95D42cyBbE1kikdCYubn
JEH0UqNb2Lg/n13iBVv7qP19xtke+ZGbLzdzKS+oRnq3WdkYWskPC9XudNL/
e1Jkcg0SKCvvkJObrZif1q/qQDwZAHGX5Qthkl1dyVIUBQlgAbfJKGdSIr9w
eO0ZSXM1vm0+7ENaVOt3NxRSxJwZMpsSp5MVt2ah3NrGEU+4Bmb3E+jpahi+
RAnzKuJmZxqcEYXNufOahKb45mOqs6M5rbM/cmucWYJiZHXrgswkSmYLYvex
eQo/QHYvRMI4KOZog+FFBPzByvi+oSa3zK2JwAdOq33Tf6sRC2FV5zLZ4MqL
VqPtF/47DLHevHbl40lhZ0WrBmFukk10x3UFPI9zTWMYwe10uEAZpEZSne4y
jM8k63cEFuYD89Bui0nSMDECHdjAF5sXs6Kv2GdOg5GyqwWdYOxDjGsaIWnq
8c38pOpeUkCO7xJ8L7+dtEnHzFeKZuOZouYZWYkab3yqDW0Az2VIlm3STR4q
9IV/EyQaYLAU4yyIBc2GXTckiStKffFLN/UtNBws8sqAJ2bb74J5ySem30il
JR68fAA5kwKCmv2sdhlsoludawLwDBFlC91FpZNjOM0tPC1c+seRQsurrEpM
3S+tFlKDUEIXHUZBpGjQRxw19Zeio8hOqqhlEZ1Jfh6ud1qT9DMb2CFuhjcv
poUenBWLVMqke3NzjZWUcr9HaMB2E9/+JE7vyXFS921dq/NMEGt1bMHgRnp6
xB6zCA0fLDFGHeQW1vKxCOT82PKm6BhD5b6j3JR61o+5Vt5QSegubIx0HCF6
T3pQCjdcvg/2Psa0POSbyPivpR2W+Sl+rh+AxNFcHM6g0rUuL5+CYtF+EMia
XlBiTYlaFcq+ot6HbtxMeb08Vz0z7qVUkHqvNVvCRNaeaR2YrVSyM+oCQmBa
bBE7zZGOXK79SnvmgdO1mG5l5c2FqVzZ2kZ6YtuY3ys7YSeM+HB3WNsJCvm3
MkttXbL3WplbAkIzlERlhH6vfxcm/Z0CeUFPNR90S4gzfX5AoGRNr3qMwXo5
mAnN4DAf8XawfJ4GCEBKQlX6R1Ha5qgYGgrEyS7Zi1eBOnFnasNUgn/HRPmT
9NbNEAsM9HxqT8x0j6eEl1hD6XUPzq6zeIghQD3zlaxtYSM5EdZCk1W4SGda
Lsh+TtvwIB75gON5vab6Q1DnSHqUNsblQABO4G9BVJ5H4qOTqOKGmW48Wbxl
kjbc3Vt09D+4rTqbvy1m77wwJAxJIY9WMr6GQhDOyaQOmxosHpliBnf3EJFB
fPHK3G6wOJSRRDYW61t3ZSjn3LyR29UHcJtd0wXIhn+TsoziLW+luqCSp1pP
/J+9XOuhzHwYm1Oy8OnrYKWweR2sLE19uHEx3/d1SDhuZgODDRUKcfT9mmp9
TrzVns95GNWP/1flLzpij8roxasnOKYwS6cbKVT1eGRlqn5K8mZZxeF2pWTK
86S1Muyt/j0MJ0U0dvuDiVtc2kgOS6/zl4J/JH3QdFagqwCXpfYcZSIIxNlj
EmXjVMGDQZeTAoyPciG0hOQgz9udz8QHrxjA4Kurqu9zQss0yeX/TAbK31XJ
4Rlh3LvY4Ymnl2Eq/fuCivqRNemeTwK0TXB4GH/ADmwbLeZFfdJtNPxqvIQZ
3Rb8THMSJdhNlUzElAPYJUBOXPIDpIN6NnKiLf2g5ClJahMb+IVcukPBRksC
Gb61vYBv7a5a8Ua8j6iB+UvCdnr5bH1qXWVxxNSuA77D89Khf+Uv+PjD7Czk
H/6oSu20GNdjw8ggc3SxDkJivkX21Cb1WDVeF9FrUWJ1+j1iXO8J7kwf9S/A
L8fQI/u/WLQ/SuE8PwTJ4465AuitPrFNw7ywA1IUOFutLXauvqavnB/zaucT
GD6DjbgklzA8+cnSksSNoeRAA5GQZZETvfBD6dxnqdAXfQ1Sv1oRpLQnrQDp
vPULAjxTVTwifY1xJOQYnMV6uWNpOy1TuNbKZBo/U9TTwHwOXDVxr7vjVXCP
P+a4GAl35XgKW9Ql4lgkbimTfNTjSNMgF7vIjAdw144TsyIeHQfcTV/EB/5a
CWSxnGHFvWHw8NNy/mLvlydRNW79WOV66de4j3GsEimxjYiRvyHTerx7P/dU
om8PY/qHoJcyuryndGbhkZGuWP7CiOmPRm1wzALfpacbcYVM0vGpOuDGcoZI
VasMirlxOh0GstOM79CJdtIwa6hkDBkC4fuJL2B8koWHo234oaqZSrhy3Po4
+LabtMXHiVy/5nVckAiA78xaqb+dHbdsI55/Zv05y1KwPu4/LT1RQ9dw3BP1
+bwqIxKMkMrhvCXfnvdN37lHoeEpADeOQmBf82izBliowhJgkEzp3knDvxLz
BeyIhet5+EpabyBTZoRXNKT9LvlUaIzPGjpkUx9Gf76PsPTFfA3vS/KEM7DD
kviFn3qvcC9ikpJMrY7m+lBiK+HbW8DoX/GdEge/GjvFeS31aP22zbOuQ+XP
nJJ8enTjtYfrYjzpq4nROz5Hb1owPjR/HFa7/joqM/1+SyLzzOWXu+J7L7RD
yvI9nKdbJblYLCQ1Mvb/XDkkGFHrj6hJdeku/RcuziyY1fH5u/bOEZ2fQLsp
kN9vpdWvHilyRcv07K04HF+ikLolw7sA+ZBVPVeg2+GPtRIKie+ohmn/qU1L
ZmZus1nN3cKX529qm5wofe3cul1Gxrzwe5Qb4/7iGfu4uuBPW2dOw46/osQt
vFGMfUCiCv7eeRQo8P+YEXBwA8UXPiFP2HfWUIZW6LEcEtNo4WXD9xOXhtSf
/YCFCHa0HqN8Z5/vn1lpcWcRwlMwPx8T7ZEu0WLuDvqE0Kda8j4ni1zFjSck
tXo+UHXTngz0AXKl/MOBq6/2xfNPVoVmuPPS2Hq+bbKp7AEwZSCwA83aRBRF
yQG9ozBbm2KGCq38ms9PKgju1vBMxCGik4eEaImKyx7AhpWwCMZRuOfo3D2U
TP9OBQO7Lqs6Cxr8kF8QR74/szM7B8rplTi4/mQgE60R6etccd1icebpHA6B
OxDcjwriPy2ti9mquUUXAuhawPnBz0upwG1d/+nAP5AC5axndPSfeUVFmVIw
8oMirGNBw3aAWxTgyGvu96JGrRrdq3JX4gH94krfFOZKnyH9xUxVO+JjPEcE
OheujkwndM3uRBpSiMJhbi0uascpo4VFXWbEOrTXC7mNeoEXYfj0hw7kSqBO
ZBgCuXp8tN03FmiITXzNJL0GkYyOHg+e6r+n8naldrMeBFYVVzHtuHxPeDeu
YdKwcq9ul6/73aCrFK/7tBtB/8hMpvhEDYe0AHVmg4xmuAGdcUQlb6T0j8IY
Dziqwp5KuYrTGYx9G3qsK4vW2J8Yth3XAsUG0kRDXvV2P99KMk5lg0RcSBPm
w1LAXl39fH6AaRbXYXA+MZuC2b5op8S//RLIXSc+qHDQre/5J4Ub2Ajs+5eH
3gmxxeTdMxFNL+DQOx/TbHQAx89Z8EVXPt2301gWaKusk8VIFsYac2h1j7e/
RahhfBGeXJ0ly2kcfStHiVE7ifTMxEinzcvOf9PwhcgogSkL0CY0bcpL1ifM
Pvf1NnP04rs0KssQi7KFmALqDgFlHcXeq2KC5NX4TBOmPqw0RMmDoo0Ow6EA
fscvdx8o/D2gvFHUTI9G9ZSNV0kG3KadHrTZAkZZowAFvZu1C8Ahx5kP9R3F
IEbp3ajKXk6ZrNop8w2yADj0dQkTMIhucTlXcLvX2xy8VuVp8sJCCbe6Nkmm
m5Nqc4VBdO6DrNkjHzUF7sZQ1Eznsg6Z+Gnm57Wb2xyeA6dY8NSMowndzID4
7D9eoe2kcGx222jhbafYcYpzV66lcpLXULzNioVZSlOM6X0/PMwhzLR3A+j1
DqIiO9X/iGzS7QwDqs3q/1eCLtPamamFpPShfX+bRuMPSlArDTfZS1K45AbL
MahlT0rkItLvAoShyPkGJ1o9ei7EhCqo7IpSMzC6WrMIdwAbagHptOZMxaN5
GTeY0ZiHbKL99oWUMjs2c+KPoPyHW6HdWC7e1ogeJCqLTd+0BzaOMfjTswH4
Bd3ak0lThekKKpkuHeOoxy4s9pBWxEP+z2gbvOw899yaM6x8pDk7PQnc8/Hu
+2pUlD1puHoepc6ADc4eSEZYTO19Z/vCLp9Ce2U+PzOaKGxUvkveOLUrPiff
OLUN9E6/gDKKV6cG0CmkeCNo3t0tb/R+UyxYnyuzWidAHnNsOVGFRQ72FRTJ
5Y8v9vtYc6I5KFQqoAukOzBJVVg55BaCMqDlCuk+zYUny6UiXLILftQQ1atJ
4eQK8/OadFOQFFEYDbrVxy70VVFgO0q/m239mvH46Hz/O/Av9WoB8QfJOIl2
FepUz/mLXyao1d1FXWOmb1sy3AexsDStU5FZOmIA804xtxuiiQbmqIAEfv6I
m5liwLbdhOm8WP7YusmTHOF6HikpVh2rP7F3rcXiaotwLu/l3zpVqUcktyIC
0+R1DTwZULccGgRHxOlCMFHBwDGgyIvpdin27PK2EJeVwSTqlN7AvzLIVmKw
rxbMewdW8hlLeyTzdXChPybkrV440K/CxULC2MTqd0V9cVR2N1vSoXfhiiWs
EaT6d2muEMt1le8IGlKb9JonGl9BW3hecqIeKNND2iKUM8roaMBLDmpGUC8w
/XcNw7uo9Fq0CXqA4/3Mq6BXHDj1ankGgz6gbzbjge2uAylGrgOE0L1Dhgp3
J/0cSFVY4nKPkVJ25SsIa+sfy2a9RcgzVlP6wNRZRnwx8o6/nWoqry3l9wbN
8FdUfne0rXjupaR2YmR6C9m6BmP5Yu/tHqHf9WVDg8o4cUn8dx5jRxGi7dzU
lgXENtuA3ljJtX1aY/ULl3oyQZbA8WGLp/8iar1XoLRoGF1D8xdvN4opAq89
J/3dLyHoO8du20qmrSMntgdKOKUCKFcK/6g1UVKf/QA2q2m/aCM7yFa0dAwl
aBsbSiqju1CVG3RCOxIheixp9KHZmtL/SEt6mx+8/VC+suRBLhQCgKhBOxEM
IBIdzV8o/KTwQpvE5b7ZLmchJarOvcTo8AIQL53wcCzbLGUXe8WBtFpaW9US
19zCNCmuF5lK5gQO2xtHaJt/TlaaatQf4EBe+g8vQZhtzvAst6k1sGcGY+FT
VCrxh0Kdq8WyYq3UD/bEMMY2gZ3LrraM2Y5GdbfcMj89e0Hqj4PjG+d3ymaJ
ixmsAdSsCvH+Xe7279qnFs27hxc5sFzx01rDIrEtgGTe7L8g0XgxGTv6e3s8
z92f+DwGJKivmFoi09GP+J0RQoW21F1T+uliqnoqIDg7a3Gi3Z1nVYucdts/
a6LHUFNXbYDQnYm4gOV8kLD9Zf0x+x6rnJo0ZU0NGWLcPnnff5jNsltZSOiO
9hNLwH6uu/K1gTX1kW9bS8SMsSZWqfgtLM2dH+lzhkWX+flmBwCVNmZaNrSs
Hn47CWa2XennbzBrJgHObNlykxI1m1kJAEekzRUasb/L8dLXXqNnfOdhhWf5
opkOHOJSwdb5jZbhm4SBA9xmqrnwIQKTAxiEsvfoegEEw6/LReDylivj/Bcg
7ocHGnaQ24x4taywqSmyDfBipGA8dmlGeLwPZImIPiWXsFrssa78by2njOe+
gVbTnQ8okX0z002HmMwZQEhQ6HjOIMd0YTO65tfoCe7DYHwVCjM0PCePH4bx
NYr+ukiUTNaYC0tNDidIZJUImtQToF006WJEduGMbxEORFzv97vSOXUTd9Lc
4XWUigVEAChY+pzVR824kkgkLI2ZuPOLdlHQBIdGUtscv2yVpcRLrWHaMjvr
yIcDLoa2VaB0DbCMfk/UzqaCcyFy8YyS/Dt8E28zj9ekAzXKt4z2zvL/PVGa
aTVd8bHscXDWp5kJgtknlzYuglOh+lZwq2KebFmaexuBsHFe00j1YVvcz8H0
pbQEh3hRSvNw1TWl008iKeNUAsAqDPfpyr/uE76ebiuukOqgYulZNpnK+V5Z
zReS/pLhOLdel3cM29agxNYA04H5qbTAZJKPwkthLkKC6bplMTovRQ7kxbjE
ZT4kVYlv5WiZi5vXi71/RcywaF2ABRThTXpO+7LdAMBf0g/LsG9bSK9UBi2R
yeNuaKTuPKH1eZNzQMX1O1pI8sD1xD4w/fko0wiQlG+CGfgeUEnoJZ2fqQ7b
CO0TcccIbXw3R0li96XoN6sEQomu8d/DYYOCW1wQ2iFhVf36Vb0Y/zlQxfXX
P9jU8LoEpyYJ95w67XIQqQlwNkTFPc+DSjvO6QudEnHc1dzld4idnwTazHEP
CfuBlqwAbLAFI1kuJw1M3JGgnNOxjKbiGsxetfame6Fimsy96yCIFdQGzZCg
s7u5jNZg/sxBCjQdhf8jVRz36ML3pFpkA3N9ziBhP/z+xDT/PSuqLb4A7cTi
4ytDG1i+G4ikJe9tCBKQQ7RfCIv/X1x3EPEUraEgEOjvgDkRkjHVDcldKxNu
mHeptUaP4IkJqLHcbjsWdqEFw10UjirgqqWQ9EN3U+Bvk/QjAG4OCBRSU5En
WlJwRYF+3zDq13JsCLfPm/JR8ycTpstk8QT0OWxdI2fIEpcjdfONreDprzEz
RBp7RKzj147p2keFA80zE41Uk2eLeneIqQioaeOgqv3rZzDiDwzSL1CtMzin
0aQDSMMPiXu7KVvgPHNaJb44OtvB3TvazvRiEwKvSg8eH/xY+4QEGURlFRJf
CcL89o+A7lHXA5LmUkwKVnmcirUuTwiDBlTF8mXdpv5JelmrfFLKn7ZsKaWe
ObPf5SNl5A9/1zM1vrI4gWxhjaoGQH4VTqtMezDDux3rlCl0EfqTQ/KsZe3E
3exbXkJUTuHggECcvXv5c5d4xsoHAZjJM3wp4873QDn5JeWSomQoC8FbQkye
/pRV0s4Nvhplw+lOU0D9YEl6hlLQDb/HvGj73tKBOP37H4LMdJWKY5kzPSfG
ZLy5m4a2oe6OhwaLgfNlOGHB8Yi7amCyFfk+oWkt+J1kpPgn89oEC2NEwGp/
80cfuMIzVL0vX2auFmmjaKmqOi9ZZBPHmDBoidXYlwB8Gbq4getz3PlU3ftB
liEl/7jL7jrDWSPmRpN/sWfHEr5ojV0FlpvqF50ALih4wwPZLh3EUEFMYVJP
DPsnurhqF6WN55G7zsNtCyY8IuaOHH26V0hYB7Inx2Z1bHdWbd40Jg4r/D+w
ZgEpJ6dwoM/LtxcJMBFxFkU1ajnfmAuRM4laDowj3/Um1nkyz3vWbubN7tOo
rwEcL/9b6d0IMUBzhnvK15BizldmtW/DXpaZCU3e7dqy2JBJLDQJfmKd2Xe9
e3Aq2uI4RyE1zv9ZIwWegZnul4N4jSiiLnjBakkayp0yKYui/aobImwPu5y1
fcuKXKTmN6ERZkzNG0tmsjnAwH0DhQyVcTkYjIYZRmlAYtFG15nJSlWxA2Z1
xgx/fGtuhfh9OyLU7Ta6JvqXXQDySybY33FAYyBPM8isLvltc3Iaa4JpsS+m
0/4SvqGl1ve8kf5mgqVK/ykrlUzKG4I6mD7/B8hyGLKEfnMjoF6Szo0xuSkI
WjQbmVeG8sLncKGDSZYflLU3AV4v5W5nllQ79z1xfMFbhapwZP+EBC7nctY3
3R4jxQVR2icubOFyoehd5SK9xKINVhehgOgF1UVa8QRmmkVS68Xa9G7C02WK
F/FeB5tlaGONn8llTVLy0sJwN3GitgQAsX2/5w1iFizxKwqLYAMts3+tOwVN
4YAcjsgO4+Yd+ZGwjJZEFkPy3/vM/PDb0lRZhw/0PRPEA3vmSBtfY8DwHNPj
RZkmPh0HWvOsziz1Icjas6goxpnJkj+hBOpnsrdfuSRKuE18Yj/jXLM9Pbnu
ZLBNLJrSFtdrId2FIrHAh2e5HsbI1YQdhA8oQDT+f99K1W41kJF5GT/Vz7bp
OeI0TJ9OXMrRmebWwstLuICk/mnMZxTmg+IHweVjRglgoPLjNeaXpaTur8tK
6sdPJiDuHDWC0wCksBqABYgw08gUZN8JtOiQeKiRMHgZY/J9HwRMV9Q3IJCA
MOXnowmIeZuDiAXij8+G2CK5LRRNzhLxj7L4Qyaz5sfN2ZaWZuSU68UvQH4j
ClAjEWXFAzCUdgKv58ntfXoma/Ieo3YssOEMWl7oXMA2cKcfXrIA2MG9X5nu
boi9IU0I67RliktofAi8kG1zSaTEfSYShDkhR7hbNumv4M9uova1+XMdVOSd
WSu9/udpnzndpK8uCHDLW3RE5oT9pV93m4Os5jmekNh49ZXSjZxIWDQOk9no
UEo/4NIQlQitp9qNSdEf/PD474gnxAwsUOdU9ifmVAYBI5mpUPR99NZ/DmTX
fEVcCg0f9jXwc/CpJCY97OwFvLUEuSXCYK+Vz/q62LDJO0ZBMIeIOtlSIqDq
mx0D++1zJSS5I/LhB2YTkPv+ROjOFFelPGas5l1JXzfV3/NtPvLEtBxg6l7i
bNKj+2zrqgYWLKBvNC8165NjqnPwjggFeLX3MDklemnb28CDtGIr9j6MT+fu
5GYuw3dBIx0CW7402p1pEadilTMb89ekrEosB244pCJt+gMIN+vvEW1jZ8ds
P8aZvcqTN22MYwPSUO4DRDixSOxcSfWUembGZhNQRH0rqzuRRcNoqUPtvFCc
Ea2YbUkWLE6tyXDbarRnPRV25CrtUmwypzPb0x8KqkkvgFe6LcHoXqcRP722
wePoWZuBnbdiYGn+d9qdSyG6XHda97qgmVZ7jyU+1akUG7v49pR/9crokcvT
CmJSXpossam5xI26lDWoOUsY4n+WB+EcOBTuvi9dKMnCCaaskSGN08um56+U
lO7v1HaWALlYuffopqeLsBdz82nO4xcbWnxzJsI2taBLWcDHvuClUKOyFG3j
PNF+p4lwtHWf0h1ORYfTEVbif0NmRpRn2jlkhUr89GkeLEB+BIUyujq0zfTn
G25SFntyHC20YiTeQeJ5C2MjV6Y0fjGZKtXHCaliWo69vqMzcodge1huLIO3
DKHYPBnOzCixHiH9qSsRWDGlTcc0/6+WaMPy5wHHKhy9UOMDIslvARwEdtv6
SZGey+OK3e+dGoVho9exPln6WaOcoKf2O8j37496pjmWwhPlHGbJrWlPpeRq
ysrjF8ldZHHcWehDi75os69wThuYUS2zOes2NSJhNUqFOsxFgN373F7VlMAr
zfjyssopTNthviwPDpHEgn+Z/qGwpzDZ+g1DnvJr2qsFAZAgaCvj89/Z/trG
5XVPW6Dvi9AqrJ6oyL9jzIxe3AnjVH6zYDLlVWz20oFIIS8aaeAZlaH6y/0L
g+l+bMqr6K0yOVG4R1S4WWXjNtQjcwux/GZ9R6aHE1SCPSi56MrenfaqcEKI
XzO2W0IW63atgGi67KS9XQcL7v0yTcpheGMbNqAvIp50BIm0oLqpP/xJE3aX
orqVz22SXtIPwd/oDs7ijv5JQAkqgYCHBVtr8PljMrEZlKVHZcKPIAtXCjTO
A6e+MMPkk1+adaQRTVG3SJuAU9nP4odnNrZtkMPdf9XVAVUBaCmUmcV2ewXj
fFGBwhuRCA2jaH7Ut/vKW7DiDe9pSNcGyDG1+SyuFywdwbieDIyq2fmGmHS+
sWjskNnGDEyZbkVEme/2jjLlf4Uvo6OgyXmGIqI3l/m2i4T+Rq/yxQ330n4i
wTMxKyg5lcEXwPUwxGqMssRr7MO35WWTDrfYbeaCv3ZjuZTRkGmSRC+80d/T
8fz4Z1wyGgv8NCSM2Xf5ygywAxFm66N+Mkdgz4GMc/+3TzEk1Sk4DN3gt+Ch
0LvTX9hzt++k6ya1g2W6utLXlsz58LmPhgstrg194po1ozTlU5FMb+KhCw1O
Xd1p4M9hHhI5ALJWoaFJApq7+kY0TnAFBeN0A1ZKwmJmF8m2AHoGwZxYAoos
B7R6PEy0F2mlrHKAx+YTMxBb3E9XXqqhZmkS5JniMhtGS9Kzwa8YmmaHLFp0
QZf2lGiT3McGp89Kntd6XgMO8waZkp257WSo05LBN70LJtR4oAFMeLebF1Ge
dvhbnOCMeqC58yfyIhFMrhqUT5mboJMH6w9s7enspRIlvQHB2mIvKs/JRoml
MpaOdArrlbpfqLKy7382qZY/dQTNGppFaSovQL6uoj5tjzX4JLPZSsWR6iKg
ox04lbeKdTdqBk9tOGZkQg1bqFfx8NOFUNFyCYMHcGhNPvzVQycPkNTPvQia
pT6k8auerOzMFnXaTfMjxglNK5+9kBHQ4wb8twuP/rz062yobj+CR5gi2l/Q
3vw6XcnAFAsTSXiyvGa6JQ1qnIkYekkcryp3UrW0CcxYcaCik9aLT9UjGG0w
vaZkGRwqhK1bCPtts+EmO3yKX+Jbd8CgoNcHzawyeo+1mkImZIzxSl2OpUBv
4bYgiaPhIM4p8+35SjX+FaNsWKsucNgjlSi8h1F7ebu/olnfeTkUmkcu3sct
ohFgjFA+lxm9TamXjmwEGjMH7LD0Am3raYqjaH1uFVii3lgxxUX6YeeADT34
KS+NY1AeU+vePCvarN068AtIwTEBKUDUGGX+auSM2TH9jHrNckeiFosGRxWT
fb1PCoRq1+EdVAuFkAKpRVpYSXZM9GqSPnUgMvHbiayMj5VnKv2k6uv0hOD+
z6fAWHbzhi/n9FjPqg12IPx2oT5Vp7TfDw0q1kyhfM2+76AVOGYeimmfBiEL
qYfdCTzqkm0calxvKbT4qB1lyhZAhq2XNPWXr9P/6CYk4mus6ajeqQbqsmK7
YBtO/MGgktmZVZXDD3sHqmPQ3zhl8RACCkBaSUIKtMK7KJX+VG/yM4yAn6HT
LG2dl5rrtpv7VrQWwhTbJtsaiZBD9bj4GFHd5t5E4/97jiAtcKl9li/+fo3e
Rd8bfdJGGReKh+4K5cRcEoyjun/N7hLmcZa/Kun7WLLqRlV+zGDcDKG5jr7X
hhn2LWFHQSzXzE/g9UIK82zWmVK9uWXRlLWgeJh++5R8mtEjo0VlxNL6V0FI
4IjhnIthCuYHh4bASvRab3f5l/s4KYFca5E1NfZteYZqtFhrhuRF3v9NW03Y
UnxqH+PeLycyxZzSV1ELlGr4uyPqlEicCECfhlZ59g9DeJj0sAxvl9tlK84M
1CyzyCOJFvV2S3nhFybADu8HuD5n98kN2zx3+GdQq1n6NIoPJxnL0v2riMJO
xEW6YwE5eiKEP2JB9UGMfBugKu87Lf+A93ZbOTiTa01lffiikFlxKEz2C1jw
Hhdvu+Bgw8dS8rs6e8GID2N+7Wt/2+evGW5WfyPXMrOijrPTeKFM9OvhUTlj
B2MPJMNo72S4tyJ5Xl2Dptudd5ErdLIIFRSPQ7/BkBfq2GRJMSmdMZEmC2YJ
qHENgBAo/vUBSySphv2025/A0yPM7U9S9sXPn5QRgI6r9KbvykSSVKSod+sM
OR7tTo2lwQ7Abw4VpTnxgYWGOhuxroeBgXGLTewJZeaYTQO3iZg1V8ZwPkee
VRTTXwoZxbm+b/lTyoEcuJTcx3HBYTPCAAWb8jFZoM/Ax+KiTBJan6bAD8IC
Yq/S+3HSGKlebs6kvK5i7vdjFYbIpS68qZsqRkLz2rnXaj7Vc6jYS/0AdwAs
4d5XHa7edVspmPL3gYxgl1hmBF8AA86loqUjnbGp+Dko6iwXY3hIrL5GAyVY
tRjWKvFwTTwgtiVxJJFPozA2kvvdK2ZcoP+c+OFgyUUSNZJTQvuuVWuROvpR
foRzs5DTc9/p/KVt9zrJ2pS+S+QatOkbYZa46lHhI2wUiDiMZU2Q5fcg8biQ
wtECHAwo7Q+R7elGY+Oud6GadymsV6nNaNorp0Q6VlGWA7lYjZijcv70RJaU
XkYWa9vJe5NqqxXW0DIOTgPip+6sloydpC7qRoOzqOknoltuC0EYcglVKrdI
Qc3dREV8rPm6hkyWBSI9eGvZCD8iauX6V4Z32wKF8FpvBZyoQT1lQEww2SuZ
zBAk3rSfgWd/eRzbB5bFBysdq+dmeEsG4zLNbiC/ufRnF8z8LYv129SndgYx
zMWkkHkgXFGbGdLvMQN8j3hc5qSuUlizYycOIzXwKKLl4qPeMf0sz1Q4yU4b
hbQvKNqoUXVR1Pe/N2K9OkmHRGkp1rjqEyE4Ja5g4pqG40gMZd2muvEciax6
ir/a973eveGK9/ZyvJWg9EL5PWWh2JTZSbz2dink7z+zFSzn/l0dA60W3zqd
1EYWiUANnQv0bo1Aua1TGWXWCOeEuApDkggOVohEp7hV6nXLg80sh0MBEODv
JXvZSS/WS0Zh/cuqf9gHxsj/e9TguVx7uqHJT+MmK9c1VqbPZSGjEKfhMPgZ
xpnioipRT5Fq4P4Xsu/36HQwzB+mv8cMaZuI1SYnQJP7wat5/VF0NbYZmbqx
YgDhMJyqP0DlIguVSDQpNH6SX21nazSwjKbpColYyaWkEG+h44iLyclyX/dD
dTxM5R2iTCt9WSFgnLJzf84GRCNHbi8ujHsRme+g0jKjZ+fM+rSWS0cAfxk9
iSzqXk+0fZnwdbsGkF4OrKrv5MDW2FkLSGKUddhci2q/Xf7iOQ4XjlZvqQ1B
UXDi/JWAmJD0d8SH4v0EeggDfKF0j2dNS0lUw8XpZm6L4BL20o8LqUVmFyRz
o5LV+ijchMhXD9zDiItS8a2Jd44qEce6MXtxZ3tFIY47kVoaCtzd4KLN5c4g
K9/SRUhZY1XkT5Cpa/2vwp1CT//ev+WkaYoXaCYs9DW1EmJp07ataTEuXByP
sgkO0S4YBN50UYCQdTfAA6yfbRjHlz2JsOlCvlHdo0w/QRb1yDy1kDNrNOU8
lYhobpZXF8QVpdFcGcf96mf9Lzn/CwPFCzK1GRBCGJOMB55aSn5nIapqV6JM
oI3Mcz7oTEHl+kCz7e5lkWY3l6/oIIvELI2afFLtPootdKRwAR9qMw2FyKMf
rSOZ5wXYxbeZABbPWuLjGMQXxNeZcUAsvg0cpQ+wHB1izhMx66O3o8FoKmQP
/J32c7IpLCE9N2kyVXt4fWByDXY6rq8Tuor4z1fFdPbi1IGeQGs6Q/+8/nIF
DUy+SNHwRQfNWSrAykW9DK1ZPWmm59KRzNH3TEF1Df7hClSedYVgaoRdYuGS
VkUSzhgpO80SiUtR1AXuRG1CdNeGKakUyZ/YAbPgP75Qrix/1lOJ6sDoshl6
C03EoS3Z8ZtpeATUbXvubVXXvMlAoIivy1WUK/W0JsS+S3WPS1Q7c7fRF0OA
DArOBRo+Ry5LjzJvZ2DBIUgw79wm/b6kpPq5+lDA0Qf7uQ4c7vioCgi/8QgS
1Bi1P0fReXpZ4BGP3WGg2JDT93b8BN2mVbsPoYoZ0u7hDQ+O9hI0wZWgjwia
TLz9hlruZ0SI/P+TrqFHJDu5W6wA6LkuqNignkIDUPzabdNC72DjFlTsuSeR
ASq2aePnPMgHqkOTcCQJivpZoAFe/aMp0eZyUSBu2KRftatiEa2kRC19Vz3j
Xam+hWzJ9jUKDQP7AihZfTxi0HgDHiMr9D5UZulDH80I8rM5Jovi66TaFSy9
530V0mXkGBbkdFSyoCPVUb/kvNlT5ISNkeHs3Rl6tktcwiifJc1jmzSo5nA0
z1pVtNQrgan+93lUv1yM96gUIQR7UcBTGteAB/duCDlacmk62EGyqBx3tDKV
eozWxTApXor69rghaG/LBolxeEotrKUwoC/zG1D79HkfcWZSrLI/6ZHeok8b
pkCs+UDLdPiMkgMoqBpnrK2YvjHoP7++TOCtD+AhyMAODKMgcRGxitydY+6b
hSQ9d7K4Th+KrI/dPcVp0rPjO42kQhFYnl28O2RBtAXHr942mwk4UmgSjKzE
Vv3UdIaNAinev+Jv56hTzZWvW2JYE0UXcNupumQqhSwWQwyhFyWywpTHlJj/
YqaukZ4S66lHGtloX26wsCJte/Bh5oK2V6Gm0duVpTr1dn96lYsb1MRFNYz0
T9VBwas0W73bBUfL7TqKK6qK5zxF5F+eM5z3vxy5fFjqDIDDI9jLhgI1vY7v
h9BWU4/4lYsoKoXHRtC7fvZ/mLQjj1kMKhOWn5aPnD1k5Qp2NmE9F+/WcHD+
GXPTUm0TxOAQv88CXGZwERE4u6E4Tz4UnoXbqSgRSQcNHuoS4Fj5MgnLjmLd
lOFkrVyCt5IUGSygq1kF6CNq5ZDnzPoKTF13B2PzdvjvbemCFQqRxycfudLM
qeXE/sPg09N7ooHvuQNTTrx4p34Am3jZW2ZF9DkYebvVnkWWTD6v6UpczrA7
/ift/w+JeJdWMmBWReO8sjjgPacasclcq3PsnbPep0d3PDGlMhpN9aF69pNy
dd14k5APefT6xeqJX/KLKr6PK8CExEtgG43sHXlNu5ObyJ6it0Pu+2+khlKb
aSqwU3t/MqzLTX1Ac8oKto3c297LkPNjINACXfi7EXWukFNctXiZD1Hnd3O4
j1lpJmR1w5y+A0walLdgQGYLv8//vCY3j7n/mEFs5tQW8F/kp79MzBXLhwmF
D760bF06uzDXhpqc8Zfi5ueUUcavHeNs/b3oUmhTXAnSepV0nBBInBThWOos
5y4bE1oxkuLGbCGY5OohCGDXiBOV/eh6neLi2Xfn+XCNRfNthV5K8JSEWIAi
ofRMHicOj+MKCp/obbj7vwYMCbnvNZ65czfgOPSdXqdlnEH5c2rjGiQJNOb4
qlyEenWkSk2EZkGEbf2gLksqg8CkUs9jsU6A5Y+/wggzJk2pxO0oxFizHlol
nSdP5OptwhuGdl3oaXARzVAgTEe/OgwiYyzpULVEmAUnloQVgykBsVSn0ySz
MEfURWuBRHLGVWXlLcL0eW8VtssanMxSlicuR1WI6ZaC6WkzkUdzxJQkLhEz
swSDjtD5/ZY6XJ5QxJwoTGM09Ms4zoFA6MfBPzFmZB2T7PvHLFmvUbCIbwby
jgnXc42929E6ChNfFBMwLXtMZJ9Ju/ZgJKB7fwMG2xCBwYzZaw3b+451E8s7
uaZ+LjgAKvkFsp/HlUa7Rasi4S0jyR3ku4GE+RiataW7v1n5XKK4njHlby95
n3a3s2muZg8Hrfq63nFlb/FqmLeldWK/D42DSvrCKM/XmNuAU+hg34xVTAmE
XF8NA5GqUJ/khBYUAlOKPabRXxSE+G4gBCmYVCaUri/by2W50a0OLj50pyqS
gWmsLrV0X/nFymjqDriOKxYFu4CkqVC346i9W7zz/uw6NJxNZ7avoPxc/m36
/PY7hZH6ER3kT6h3VKSwraYkJo8emXoTd7Vq8ACYY4VY3CZ4ZSEoZEJmO8Xa
MDDZbQ1LhQCm5DgLMBvex8vNP41+NViQRjsMc8Lq0/HAJqniprUrSmD0JzHQ
oMsi0yTFo3H2Q3NyaNhNc/1OPlN5h+p7g7532Pp9SMSzq9ZrIMazq0zuvlMa
SB+ZTup5ixBtI+Z3ufxHJoZvFKJS4/UTtruf9yUOa+lgLjOWKw9YiG2kQhPF
3YP0Fhx4utJlrQlqm3sUpDzEn71URfgS/hqgi6J92ogKqDH9XL5ptfp2gICT
b4EI9C07h/A2e4C52Yg20SB02gcBe71+wiQA7Dnh0s9ciy/L1rQTz/W/iAu7
2zn16M0xi3FQDME/eodj9XfzuV2DXM63O12Nh29f3F8oW4K4YiQ34WQLMN85
8hT3VZNrAVa54mwv6wr5/dsV7Xt1NMfl4q4m7V3g1j14u00JO4I+h8Q+q8Cb
bo+AigVvrLBok7BTFNAPQwCSfdv1CL9Glf7Mjpj2RvnKHHCWsr7respzXSOJ
ZaceePC5Cs/T9UpLaUvsWQPjwLiRXe/p+DmFA0fvB1mUTw8s0bZHXIB6dv0/
G/ES5joXAS25U2lhnAX+AlrajI1SA08wC5SKXHMSuNGwZ/Nalzff+mUZbmGf
pULgRSSGC/mz9fsOHqyVnxsADk4GM8oR6iNNQmLOWBzBTvAWfDshYN1Tpm4i
7IflQ6u5r7w1v9132wjJbVQmBCgVOYtTy/fNfkY2iFbHwbf7wR2ngZBUBiYf
FiOgKxYtc6qw3wyAyZeIrFQI1/kX/shd8zAe1mf0lQgDi/50UYWlkvgw0C7s
z6pVOXa2clhaP3kJLTVpGC0NhUKCscCtcUdqBxO5n5d7KaFx8jNfFMld15Gk
DFvFkd58H5ouVGgjp4AzsHYCCdARIQS9ZJCJayIUSx+nQJOKb95780z8t3EM
HT/8YcpK82uAZ6uMKJIGBHY1o62NdchMW8/ONZhAQSfRc6fTJe/g1PE/gVmf
uRYhIXoheDDYhjnozuk3GoC/La3qWA2oa5XW3JrjU20vf85ZIpRr7l3l6U7A
za9GlXov1hZAn3GXwOAGMI+m+5gZyO/K+pBr8J7xDZrxRaZ6v0Igvnw7JP82
36uis+vLpIvfY0A40hPsY6BuRq70QpUtokEiT+5oLj9+MzRyh6iK6KSK0t8X
PchdPvrOE79GR2fj9s582hH44CzbjvD819riBUbPDFwS/GLpU15UhD92ufjt
60t7hNP2gB4iZQQtNtA7XEHv8zUlXqLUkxT4QI+qlTWtc1+h57NTvco/O0q1
LEfds2m27Ve3FjZBH+EcDkIu9fE5hB6Rb9vCqRUhi/W6KVoMeGx1KavOhWEv
Mc9p58W8sb5CWCcY8RLrijDmHQ0ndeYytdaI1CS5QpwVfOwSQjwk25ng5ow9
Cyav7HL5ImS5viMSQv08HFEsTA2kySWGqSUShLuPJfmqYjrYbo/buC6GXOIa
eUXSKL4AjGVKSumfMXixNQeHIUl8mpQWuCZ2YOCmfdss9CL9ZblxeRy+2peF
FbfLjO5vpaub6d0ghduKonrT/F6SwX0Lx4Euwq9//U8Hk6l9s6HD+oJUFhYL
S2bDQ/6HLcjhGxCGKCDjbHkzfe/DrzhZKYn/4mrxc+Bvt9CgJ+wHoGJJdthX
wFtvBXfNHkvVVlrxBhhRH2vkhSSaSkhH7IqP/cHZo08Hl6X+NN/O83xYxnrW
hAOl3ZjAZ5EY6+IITAYRhp1q0hSlrM4MGnM2ypyVTt8bA/94Z7xt1qqahjtb
0RMjazYdHhB+NR8VzjBAj/fkMHiDWAUUyCwKTTby3YW4/15p3KjV++Gbqf8v
cKr0EU+wrVwgAj8Nslokv2czAmCqCsKw86VoroDrUbtjKuPyxL+Y7QF90Eet
eOsM9bpmJP/b8IWXVDPY4pjOP840GrHNNI7cbfr1hN4XtQuyiKLbWbAUYF0o
7xW7fL6DGRxWinft0uquw+Gvt6jDWQ2rUmkWNWMSCWi1W3Hzm0p+FlmT9gFI
KzUrdyCzMVGw8VtEHywOhe4CzTWuwimYSi4ZXXWp0PapQeNPCqlKXnw26b3f
Nb2A+yYgHrVcjER7T7Tuv5Gh+544SgbQX7RrBlY2GbC64eKhiAPiVCQnHWnt
pI1/IuCVBf6uIvuqK47rwBpFMQ8UwCcdpIgFqd+45zMCWKel8q7FBh/zle4w
qp9Ag1YVDbToZ7tladx7CmIK7F2jcjp/eR/7bzlcn5m/X5X5R9SI4ZRf7Jac
OT7phZbc8mATuJcFc5Ozn7WFJtWWjztE4K2KR64YXMp7Z6MzjN5AQE9rfZcp
ua3VROU1dYdqqMuXunIxJbd/rynY1QJJNwa+e0buU01PBIzv0zwBiW0Ejz8o
a6bxs4iIcLUeE0K3GP0siqEQYpZK5ng6gRWHiD13MreMDeVM0TabZQaIVBOh
B1XpXjJCJU/zJnmrydIbC5jJKyuEewGW+DyKOqweBvS2LQ09iaK+rJjUM8Y0
bfldk1wZuInDZOO88VKlSeB0eaXG3GMzQ1rq7mj467l4Ps+pzEl0jn5ixdBJ
IucuwGEfzpR6H4k3sWZhPgBjbF2Z425AEXgFf6jmEMo2Cm71XiRWYNPHfyhq
Gp+r7SpPWkrHDYWv+aJttP3ixr6v8wDcq8XNzDJm9d7Gs4CpMq5uIGlMzFlm
GZz0vS6A0AgxID1ByZbtJbIqzKks1CP+KcINt+4VZpzy9CWPFybRvIwu9UCq
Hfkhg+K4kZ+7uNFfj4FlWwiiYBzwuCRV4H5Ly3po6+EQId9JtBhmeT1H32sE
AAEgGGiIiOU36IoflxGg2k1wC4vedFeggIkbAA9FJupRAWcoA2Jo7h2clkGw
yJqRKDB9/sm125C2AFpz54SUW/PZaKcRBdz7MLAmqrZSNEuiU5sr6i//+Q3H
nAMNJv+m0b6MlbGC06OgO3y14Dnn9jcWx6OaxYOhjSGCvPr9LhAtsW2uTVfO
hlEfQ58nf8Rk1VySqextOiAiFcFa8lTl9ggke5FksZYGybRguTClKDOPUbOZ
MWQAm61FxqC2vA/Os/aJJSFpdkDzJGbGxHdQLz5qkIDeegOBHUT8mTYIzY5j
6i22u87RYVhYngiwHtnBc6BiYZbjDJcloaRX2+jf6GOK07ktdwscnW/AA9Lq
vyVTdz0ocQxT06XSkbsed14Q/mx/2r5ePFCdD/NOGa+K61VzKCIZIWX098Ms
n6AQujyAfImAtUMxcjZxhMx8/yv95kehhmarXWPGlcXXCzc/cCVI4osRw6rN
nJxq8EefD8lSsIqd4OmPSMELyzY+2qRUNox/OpJg2XuYHeYKwl15fcMpuTZ0
I18TRinkOznaDa8XA70XZTJA0I0mMpRhATI4t1yH6WU174o5gqxZI2xrzaBB
/1pB3Gqjzzaw9s+crij7uahvR+ttU6157XsUtlRtBpEW0XD+/fI0cRh7VEKG
FWPrqFcZICw1OitcQlZHuZ33yj/QQnLNyxzlmVmgwJCbE9c92D7Y0UmMq8KU
XoZZbetTjHUFIWyq704LfTU16uwWfoNt/eZCHIoTFrpckJO+cOd/MJgn+bbl
jlZbfuw3xJLTRZfZQuQFzW326MfKRBat5CV+yUYsMUYYT15cL+zbIqGOZcHl
C7Pi9zJw5z454NDfLEip5IhseX3hAGpKEYl6PXRqn5K0fLW1HN7qEcA5z7J3
A71nYry28oy+QXlQRCxiAa/kRTh+dCPoGQjDWPX/fD6+6v7RcLmbJ0IV0GDb
Ht48O+MOsTKVspfsi9SaEzz2q8l616MiGBWBnkDMXQlp7GkoRIfAipdLfb5C
U3Z0Kgzxf2KGMTCQy+LXNINBiPpBkpNyMjbe2P1+x0RwQC2UfsAKUaduTL8d
MH9cvyZIAkVWllnfjzxgjXVyEOByL+7BwvMvT6D0BgpA712rN6lsJ9gP3oF2
HFCXgq40UvXRkk1Pr2foC19itUr0l2xktPdJ7MwpuAFEGn+35wqP9aYJji5O
k4dRHXj2hEzl4iIv6RWH76jMl4ZmAoaZzun4iT4unFJCPWiufQT5xbWDuWeE
KNoGPRgpyA6wWHyqUh0R9YcCG5FLRS3dV90rQNTzoX1AHXT+Gc1H2J04sfio
DoCcckx/ii81YOyJB/GDPvKzsKMPPFav4JlGXTMCn0xZFOpvmjPgJkk9kb3p
oF0q/BOuovYg+82p8mE8SYF2qhb5t+X7UZWgAcfKA+WtdSnqljeWWirTRor+
qNanWs8VcZVcY20Yfu1gqYp3wEtBP+0dGwCS+LJjE5CmUsOJs1MRoPFZFpOd
0Wqxcpha+B85i2wb+j6b5Z1/HDH03+D7SFEXHQ9Yevs7E8Gbnm8pLbXIVCdT
k0ZysuSbTH/YKUMszrYrkTGCGqhjdXI4xv7Hrnoksl/5iDjJtD82G0KDjkkT
N0xrtbSjQQvM8fONOkokV56VBo5Yq1RLcKJHxCYJae7kG7DcrpND6/3hPvPV
1RJoS5MQdHwip9KjzaETEyyTnT5/5C8BRqH9xq+V/DwAi5osNdZ/elMH2aF3
cdfnLISe//L88fwV1dPHJkkso1SXu/uJ7DkGOGj3SxMovwdQqSC7nV7mXqFx
l/RYu8qViVAj2TFtN/nlfqkVK7grfH8TRdGlsZoc+DpMF/FtajXl6B1er7R1
GHZHpMtHnGw8Wc+UsS2lp687gJEd5OXy8Gkl762pchilhKbznMECf263R+CC
1EfpWRZ6QpD6ewVWBSsWgUaSyBrdeW9SLv5lwDoEVYzuqIBnZ1C/dUqRF1c1
t3FKLSejXpVK3eOxEq0DLMPA059FMkc9j2dPOn9EKsXA2QhXxkiqafEJwael
9n/lbM4g03aKj+1SXGE/w3ABiJQu/xg3GitQffthB4i8vuRTxl1l4UjyPFxn
Y7aJ2Ao7urpZL4cTaK7vvXuIqPVBp2UsiDkAt5iwk4mJ2dlTDC63/Ji87/nj
yyQ9aRyZUlaGf4HPh9W6vqbHBnzSI+IK8PJ8lyD/HG7JkrBE4EOM6LPZsT8f
lwMM/LU3XSVjZNMe26mKyZn5QuCHqZ9Nz+OrwGMqkcKjwZHlbTL//vEkF19g
+QXFE3soTYFbpnR3MZRX9D2LtiHLUGlOpZm9z32Ly/FKuCtow6lP5wusMEkF
mu7o1CfaSZJvYGj6uaOOvO7Y1PCAHH/mIdlHiiE66c7pVe+3HW1HVjktgGVU
gpF7rNOC3qWKIoRBljTomfPbFR8w0/9ZXPZLX6lpr4ctLTTb6One9faB02uI
5nWT4ZvD7LdxL9OMR3YIepVOxco/uN9XQxfqEFftLGbB36TRomghLFJAYKtb
fW6xaWY6aH9VfKVkwq/O3XEi82UYjSMNvmV7qEzCd/zNLFfjipQ9Q0pfRMpb
Rdq8JSzsdTzcKnhNNG3udcmAqE2LodMsMKy00LiLGr41orDM8Wel5EGQzkeJ
03rMPNWTK/M8ahzKEnDA1Y6rtloiLe31Msh3ztQYcaRsY5hUMLniAzjyBC9A
5/e+rBuF9JFJo5SvuoSHJ5BxxWEm+LLjmMqhwxvcA14/Gx5MpZxV24/kvB8E
xeqmi2QH81HnbSRIBQwh7kXAR3y3cgPwKxl5+jFvcl1RfMybvHyEwmCjP0RM
HXk8GnRdao/J3hD0eCIRSL62qUJI6K8pkuKdl2Zc72sYtUURo78VO+NKjsjI
jr+xIYcuIkgaCXs/DQahv9Wv0UAknzsVuZCnLg34k0hSES8caJ7m8CcS6Q16
Mb9wkgZZOu/SuH1S486R7J83ntyDnQolViFghDkvLl7Za8TCjqtnBM2H8GsK
KsMMzcP/7SQfPbAfEYwUTlJ2DPEYVLg7SbKd/mKH3I8yffz3RQeaSaWmKIVa
RBA1MgsVp9C5IpVSd3eYaolgTpTNCRfPQ1ol6PmbsYcgRcB7j3jqchkFp2OC
uQufFgDr+DnbXL9l2MEFVIl4wTb/EQW0nXemmWC3HEIL49+Z7HyP+Cp9/JHs
KQW2vWQHnDVvPzi7qUv/pQnXdjHazeR/RrztuDIdJ1NpJcRmvChdgbKALRsf
LvawTX4S8BfgDCpmURsxZyLIgY5xsy3R8ck5JAvJbCHK2rJGep/qmpT52LPU
jHvo0Nldn6OO2b8dFoE/JelOEMfeYc4s+TmuZ+nfyxgblUqLiXaMCBPFJ7mF
Fdynb7nAcvy5SwgfqfWSN+c39O7QJs4RH7IFsmMo0EmckrGXwbEqrWjTJWke
pdVBgab1zbmRR2qxtVb0YY3G+yEdrWy+nrzXbH7DFwrsLmA3EG0NIt++6leP
/zMzncuvoBXFZhEE1yQA6gW8ynxQzmuDjKOnxftoYC+SraWQtxAzWWMMw93O
KmMcQ8svk5preTkAj0An47uBPTXJoEWP8EW3thIzM4bqCAAajauf0m3luoKG
b5Ya8z9g0FGVeU1rfv059CsvMGuh5epAiriY9hqWjPyN69988i8HE3pUmziD
5Zmaqsv9P5wJcZxqTK2bd1MSBIBpTQNONWMLoIAj0du2r1VXJjBtRZ9Cjs8x
dI9MsPqYF+bRaQ8shG61me/h1WZMaM4zxSa/s3VIAaoi5Rzi9Aj4dld8xCHM
h7PKDpWUa5Tm/s1MgiKBSb80T5bKmhxUssK0bRjmn8sLgkZmysswa6uQ8K7y
BhAmAO1WQJlzxxy5XwzfbNqfLjj+VuJjomfLf1zowMPbOKh7I6wGQUJj6nXS
G9X45VDkYclKy+cteZX9WXETSiMwyU4wVnon3mrgf349kOvHd4OU4Q67B4v9
HfbfHbHCZmjxC9EcwqiSMeNBLlu5qBqun3PNYUsOhz5U5cls3ABg/zseHqdX
gvNZA9sg0cdA6/PKDZw3JdUJ6N96xoLR92hTX+hdqlPoZGm8AqS2iTGce0gU
I3LpiUGrjuGuTWKepaFx3Ap0jPiYhV7Ex83WuXlkDIaGEcvjnsGU6fUXz35j
zLxVB+EhOA5Eg9fVUe0KdealVSHM4tRC/TEOtePYX1ofbIKT8EM1aS/69/Aq
P0Ryv8+YsS8VIt2uZxiVjbizbH+OXiIS31U1/IMz3ehU8pgasaVa66f1oXQ8
TTe8rlteEj0nTKS1P+vPh8l1+K3/CMgKuBC1u9MqDxD0KUkvUWB6KyNUepOI
Kf/kJCAWmOI0UisbFfF/XrKqxDyEXTvQsFOyF/69gJJ70K1cI4gSFWMdcQWb
mLgqri54tOv8HMdEoRFzfozmkRKNboLpnjNZnkm0mUhYQ22dPiC8SJfCO6ca
qQ9GHbwWObDcT29vzCw2UZdzNQu11xWv3ERca4l+dim8fYrzyR4G48A6GUYc
sTgKwPV2jkxZr2kgGVXZ6A89qHmEyQn2JZugWeXZNAtB8Umee4e3MwOL3gaD
A295ehF9jQBV65zYVyUIfcnBVRd/camnM54KuJC9LP0Zo+1MorX12xDMeYDW
ch7GGgtr7POtphQ08WEFxO93OQQNzq7lfpEESi//L1Km60+gM+BSKU3qUECx
OTiFQ8eIRcObhRw8znK8ahQGrgAuZJbyyjDy0A9WdWp3SuoTpuUNkFX+RejO
KO8LykbvYvYXAf/K7YLwRRxvEJZw5FMZsP1gbNUYHnb0i03dgqCu86M3MnEe
ryG3w/0ksuBeSSZxACtk0GkhjZ2ep1FQCkeOAErA9tMH2UzcOonkyAAtTg6z
8+PJVieviaBbNbZ1aUCSIuX71gYUy8vhw8PbvgkulUCAVewW5umUvpFGq6ka
mtQCKwvVe4ycAm8WF9Xu1MjlmUS+umUS8B8N1D2EbBt8iSObWFA205QaGCZD
JVZUulP3ZuR7Ign2b37N+5GO5m0aO2QP+QCzIg9VcRngq/iBPWownxjZf4Bf
y3eB/tzNo6FWC/V+Q2WgUtOYwGzpeUX/b+0nrG0K8XEQBfdTABd5pcS5WgZq
za4VcxoXVtHQmpz2/CYMABsatj/PG1tdlv410RVgD5eAkJW7YzrkwCqcp6Sx
qTCmAehLhzSdXy8tTTReoPXEW9XdpVLHV5V2trGqnmXMNOl1YPKyyd9FgTPx
YWSIGras3dOYL7gtSCL7eLKcJLU5RG64YLwquG0QUH+i9VooHsiUmt+8Ag8t
KfzhQHkouevRFBg3lMfiPQnIsXrrCurmejAwQm3Ecse7DZsjcm6Pv67xaMG8
vUDNy02K9lcx5JreqKfeVXon+84GZE2HOcqW3itBQhW/ipJOZRLSKyAvAjkJ
nzmvssZGqO4IRXprCLfkq4v3F6J1xRvEcV1+DIWu92NnADQc1GNiFTjBDeLq
ZtquKbUw7SKZU7IsawhWpSoyX5s8qpXs1qOdbBxB+uKAOhsAxgJW1gPZuPVU
Q75uVBexFZbnYFdY+BAwkSVzUPQAZujqwmSHJ/zFsTuqGvweKdJvWePHiloR
t3V+6YEzpg/2Xp06JPlhuug3DpqMmQ996SXqHdYiN9zPczIIbglC9Rl/vU6M
FEFmVC8kQ8H9kGVYz4kQ57e9YBbPp+mmjZFCBg1hqX8Zt8bYlx/6tIfduQwa
mvjl5ZEq3+zJ9UiBWrQxjO172gMAXeoM7gRmerADGs3YmGqglFzvYuH5GgYw
6pEfUR1u4/mrS04aZU26zkbXDwMkTfp4VUY6dwxV8QtcDiJlNCszVTHS5q2I
FUptBC9IHy0gBwnzka78REYitQvBHsuZmdtDJaJqMn+l6VFjBUg09n2PDBj7
w8Zs1w++vKTqbdJ96smp2605CSCgzL12Z/AT+StOB2qisPvt8s8g63ztc7sj
c8IaCJ7bbTLvSGRNMl9+GMYr+VrXWyT0XEW24Xc4HL7mt6Lmba1c+eAQKoTy
TUzK8kOEpITo4AlVmdUxpciQA/16K53mmA5iOKJHL63BgRed6h0UBQZo9x0n
CAvHdXrlN2sxlhxJwWT1X0UG2NnroAh7NPwEQIJDGzuVIQf+9a//izp6BahE
DLA13VuwEsfYb1KZmJmQa0hLlqizcB62bX3y3i3XbAZdILqCSuDubGHTY2yf
CKVAy13TFNaVmv4EUwg4vR3USgpLSRNwZPN2PJZjnJ7bku7nqCiglJDoTzaY
ZF/B/qaKmJWWZJfvQiLhgV5MPeC+Kf8CCVfjl/GRO2D3fa1UKXM+Moh0WrWE
iQeVj2h30viE+I+Hc+2rfMlz9LfsjDz8/BtRRj4HXlg7+6OYfbaoO7pfPMON
4b8WoKeIhMwrxlpnGjSVsOibWx9PADDs31awlBnAS/cOZTLOiq/7ilJOsKsy
JIrCMoRa5S+lb8ADqXFaXEtbkaiGjpcicoMKP/n0AtNybznvnszn4w3l0ztZ
9kQIQzAQYA3kU0g6hFsGFckycbjHbQHMBw788vGcPo+4k4HN9XN89DbLEFAx
8SKEmI5CuxGwcUzwXWvRZRX77a2Nk++1mYM9enl/i3xT0qMT5BvUnN8y+whj
nHserppeCkSHWO8QoHCXJI3pSV7PQi9pjUaPApAaS0Xr6rLOZe4j4H2i9MYS
GbM2rQNOajSwL1H5tYfEXICoJ5F+FEkFmRINDIQcpYJB94/5lqhfyu1B2lqX
dL0cZrP+QfNanpgQ5gHPcJREsVqD0AZarzYii5W+AYj6v+dCHFCmM+jAzFm3
uuWU4m68Cx0ZgG8d0QLSYeCy507WPPx1+il2qN2VQsTiIsYwTtkY37ScCoQG
JF6DdT9vTAkl9bgCfS/c3NeVDLIY/M65Qq8XYsIw4DE8bjImapWyVkzDyw/X
cLQxcyNaPgUoPabqbcEfBq6oLvzPDmANmADXwklypkCiUXafiDKRlYin9Any
X0G325T0OAUhznzUKRd/LpUiqzBXPZa1LiSdnZ/20C7sZhbKFEyJHBCR8XFX
GrBJVNLpQiW1RgriCJPV4iOL9MihE03iNAnNKmmOSwxF6Y2NEXeo1THniRBF
2orQYwuyprcplrhznIcZVAz5m/FoIzP+8xF0j8f6cBhPXyy3/0ONulvWEIlN
7gTRW6G20AYssdp6fkFMc0QKutEQweGpPwIqLCw0SiD0Djly6N4++j5OEjnS
U9RUO+LFFi3KlfIXd/z4ge/ERptNTLQaQcFY3I/9p4bNGTFEKSYXCUMFMT+J
EYNV8I4HJMcrnJ/bJseCtts5fHooMIIqTY9YUoLXTunIKCvsu9PX4CHcjVcd
xsBw7Ts6Wgt5lybZzDjA9OpIsqBC5nsYYzX6sFOBbeGo72j/E8q65gmGDA3i
ikoqAe4YH9dqO2BZU6sXnscT9yApsy2cE61+l+K4/dsRU3eZjViy1KQsfpAT
ezEb1otB13XU4Okg6TIcPzcFLdskLmUBZbR5JpSmPg3YMgAwGsb1q1MIF8zJ
sxrYr4VJiJ8PaUQNtVGSCKuJsKpLs9ipKuC3K/IbBt5wGrIts3s0czTJg7IG
0IQnffclLKsjtTo6j8Q8pe0kLHTCzSqg/l+XcPsRW7fp/2hwdUqcvS9Tnu0m
KSVP1ZkmvH24Rj4fLsGtN2k742MN/Ql/dpVtG80SosEK7mf5TljuhYRQEhOw
LRSNK2tBz0NNzZGwhOKsvEJux7HAJ2FynCDQ6XR2vNoyHxOycOs12d7/+hgq
ZKvlSqtoEgzsY1OpdKNlWhHGFd43vsr9F/jGC4A2UHEJHI4LSmxpvrnPZbdt
iEIIU4WLS3VsiU5gx1Obu4qkuWgmD5QnBsYe1n+W7pPyBWRmTxso+AHVLXUt
K84Y9k1mjzSy1nHajPFLsvyPz7pmAxHzotv/rQiZ2gqr/2ImHgdk24lrE0Ks
B5/MOM6OV0dHghZtI2Rhc7c800H/NCL3nMMYoN2A8klD4U8PgtaSrIz/5V6Z
GjuOS0ibgCr6Vkg8GFjIHpO8gigLSRWKVxJ8K/pmGyYrTRdLE8Lfbjz2KqBZ
DAO8EAaLbtBzZjqquKCI+wRUZU4q4Oqgl3pvxUhJoaVrgOuC+txC3Hq2nXyD
y/rXqMFo+McL5O8ines3fzlBqcrYNew+TeMYfVIDoUSHsS1DpUU7mC9vPKwR
45b2/4Gw+4deWyqqbWDVt/JZQoWd51ACy1KJrQcUtHssSnMNBScAledbCOcm
ciFm8yXiZJCHmGXKxrAMG3sl8Iz/qanYf9E6NRIaTuFqO3Q255qOR3+zJfU3
8u6+CRnpjd5XJ24HXOw1HT/bHOocm2VFjbV8LIv02JuH9sosBOXcBc6U1OyZ
EKSl3SZ/X5SHBoljZ802AFYIcpnLPNe/T+NdD0oGVx5soJR3yjUG+RgWVKKa
J40aNnawXUQkRJQTV2mfMJj4baOcGbiQ8Aynjuqk9u4L+SPJ1vLV0WWVO7D+
MH4fiKDyQZ4xc9SsaEY9EmBoc/W8dkgJysnOlkAZHBOQ/GfSdKog2OTuu2M3
sonpwseLAFdeoQZwTI4aQWUUbNYVk8aXasDW6GzJj1899aT3ztaQ9sHpgOTA
h4Vq3OZWtAbgHeD6IAGkEYz9GkIJDanrck0NY3MrikevbOK8dCVAdIljguAr
tzTsf8KGES+muMSPZnBQYBX/YPLmhGBU8QpoRievccogz9y2HqjmWsEZ6WAI
nBo71IlgAfSZqp5Z3SF8O6Z2IoDwOQh7uWch/TOJ0NEb6BD6Xxnq+Hm+6Qe/
dg6YzWl+pedn6o2AgH5Mw4EmST5gmXo5HwMx+vhdrMa0SpZ0cwIs1I/L5DPw
EarekTevsmWCc8QrpAl8aG8S2SiX9B01DCYsUMePs5AzJXoGuliCq2T+O4O+
DaQMSdE+Lh2/++GfPB/lLiCTZW7AElOV8wsjVwmv8xdjy0LA9+twmFYYvs2J
amJTx6bejwynRJtqkLNemEy1BqGcomUM6gDhnH5nF64nKGTe3yWhlKCRogGu
WX4W5dzubSj6vfQwQ11B4dmQRdMmhccPLkImf/aMiXeQPNbTlOJxXRwtKwhF
vLshx3aFkUykpdvpUFvalP5Hoy5nornkJWDAfnKCrsVPTK6nFGrOpDMgTs2k
CKiZ98BZWeP/aul3osbd0KwIavL2vMLIvemh+pn2Qi24aqqa7zW1Oxbbq14r
giZn6y8/uyRdxrmvO33Jg4YYe6v3/r57Xk2zikTMo9Ro0uk0u7X1RwL3Rgfb
Fd3bDFUL1HHdV/e55NoM/PhjtOQpjI2CThAGSfyakVn5QyYAjE4rSni8TLJQ
2cQYWk+O+azcVZm51Lhh6ckbU8Y6WgbFf3kq+2yrVwARhkj1gPWdu7+Xis6z
IkU24NwEOa24gABB9EWIuLSTiVYKEBVL9l2MNlC64CEfNf+lQlYZv1eKtQT2
8d/YhchOSDY1Vao4Cvoth5LD1L0dt045wcNhFiigM9wx2qXsiZabiN9uEqJj
h9V2Y6t0ffDVIu5Mcb5AKzWj902neUX4D2DHn9zPGvI2P2L8h8m1kYl8l4w9
68RkTlpjWHvdZSe8EpPUbN8ZQwfbfGWMozQsdQarDMHdMzWbEiPi/r0uYSVU
2dHaPOjb0ALQ802eLI2jwtfvU6TccI20en4oTc8uR0Pk8FvozYKqYTd6dIom
ZpEG8QdFhu+EsbcdarUeSJkagmlWuCjG8u4ztVH54Zj7kD++vcn9fLKO8QZn
GbnJWUXfKeLlsZAxxlqgdcmjm2hobAtS04WJWXunDpAbTU6Vr1p6y2o2SFvH
HPlmEcTkjm84XXUk6+WwsTj5ZOgcX90w4G+2jpgVkm940+XmyqZjvnMPMKBk
Y6mN7oxDTc4Gut6sdDF0Zw1QIZ+J2GCEfCeiMyPcuZ2D0TfVkz80PHP/HVDM
1pHlkwDJwAc7u4ygw4/73VRgtP3AoUkX1dClji5joUw1r19zbwodTsSJxUi1
kMnuj5ztspTkYAlXsNDgZ+quL1WSB4ODeuzWcw4b6mSyPGu/3H1Yzc8nXdb4
18u6phgP+3HJKCovxJAIhrbz8l1aP550XBabIT1+3Sa7jpTOy88lBapiOohi
mwGZMtnjnhFplL6gbeXTG1ui0iZlLWRw2XTb19CbcZXIIC9XTmjoJv4FUhdz
Gp1oPV7yVUOlCfz91aQm5GTra9Pdd3JcmKc5hjYrqqC7ygBTMxDThJivgDmb
Qafid/nHmrCH+TuEpbj9N6l+1oUZfguaF5zTw1zu8RfQiGQqdI84+Ui1FB6B
j3auZiodU/zkmLOpVWUdoXX/QCzLEY6w232P7DIvSm8vjO+6DGTaa4OVuXIU
+77209/XROAQ0Tr3TkDsXymjvMGrD3J9UQ2lZ41RqjozIOFJWqp8oG+OGzG9
lpjt/+eYV5rDI3Qd8IKMIx6wgVOqLhnqmzvB+wW39TX7MvxH26Nhxk3swkJk
9fxqjHlrGNPizy2MAeDvT6gi7l0/FxbXYhcD8Hxs5pRFlYnCiwSyRaFKzZ8y
BKJBR+NIcqAfWhARdcj4RL/+E8URqA7f0qqh/thsIbrOMUsZTJScTlRWEWBF
jJGJcoIrxkU/n2BuNgnRzcFUk6mS5seDFY2CRC5+bOQ8VdMbED8uCCstYLw7
lmHoTF6Ii4aY7KXDDcn88kX147ylF2FFt7fDI+oH1X3QQGzgQ00jcyNQdmRq
fJp4G+kq+142gUg8e75pqsg04nU3W99c9PxpWUdkGzEYgWII38ntvxbRdV4s
RyeUGLe7ChQDVxOfruhDTDjtTyrFYDGGNPpFjrw+2FfcE510FRXHkn8+f8qX
8puiWa7r0cPwIq8YTdd/zYJCC6Sw3mftGO6S/zcEYz1ycUbwicd33N000rXq
n83lj9FYmpW1rtMYoqpRdlmgY/33Vsv7+Yk74vr8TAC/485W6jNQZvMKRimD
P9JZNfeEQihNSH3pl84kNW23lXdokvs7vkLYrxWXjVuiyrxVBEqGggyaJPmq
5xFkvLp0f+1O51no9NeHP4Kv14gW/LMaRXP8HkrkzmN36xVY8oq1rebdU4dG
xrNLtNmxiaqJRKETdvLwnGglxqRKADX+aAMqiGcJnx1DnpKdvNKoxjR4RviW
SbR6jSzqFfPV28Jg5Y/MCE8GmZyWkR6z4dXFy0qftfyhyDGa/IwbouRSyKoR
/04oLGBufMlZQNJTvW3Q5XnCpz/w0JRNgd0bG98vGZkhTYtnh+7zqtWHuq/S
F1opwEwZUN5koyLwRQLvsQEIa44a3QTEfi8f1weEURsGr/wwt41SDqB/n7ZJ
PdTGIhmnfCF6+Txmqw1nyuNCtwS0UmijmeCp66K8juTLOP+Q+2fF+eMshH6Y
GaMaUUs4AVie/9iSnIokvYJYe2zimHQZBuqmsbbJMKAeEq9NgkyVA93xYd/T
7/uDGrnQfkfT/DgE/9TX3LaUncFg7tSlhU3M4z3e3wUvYrQEF++P6FPuqMLX
A6s2MNYSsKiGS+07ed0L03QR+oIU3pM0i1fcwFpsEE9jFjt8pdx8inzTxkuE
O7/PleA8ZWVJKT3lIF3pNh+/6P2UjHEXN49fS6WVmKIWmDqEC2Uhwc7cV8KB
Ln3Vb5NoNY0NhLY4iA2SOHWVGftF1dnId7quqGfWHSmlB/ICAQcJ4o/wqS5X
vNIXVT3lUrnH+xCS6mJsAE8JPJbpc9Z4quN4oX2X1HnU8Vo4o4j0S0MOpp5I
MF+0Ic/7vWViLCJP9lEqTlCsAHdpNr62W94FDdzYmC1sMps10WLamNcSBurZ
X7qCv+O1hFZ4OyMLFwtd+vJIk/nafgv3oAUVno1Csschk5NW1VYso0hf62VV
LGUf7iPVNrQBkhIrtjFEAmx0E4o9ypxk+N5dqnFhBpHU7j4mHjZ+qoQU/3ud
tM+izXagAOyjXii/Z7hiYfQVyMuAStZsGeCUp+OQVR9DCoA8QxZBUah0+F9D
g97XctEnzJLj4qyHyL+tTIMuL9jdfKMN81jcsFplecuXT2vLdcsVsFHkK0TY
ly9lPcA0NTKC1f4hBXqpXB+Q2wgM0IWE7vYes0Bb3vZdL0B9Ep5l8eN70WT5
WKyJjGnUAwWAzdjGaNCBTIqKI+G9q69P0gJkGzWiNM67G3FokqfgMhvWU/C4
TDRBck1AjH+e4rJE16vADzLOhU+jGjKUjYml3YsPEebsAVYxOrx6bJXhS49k
ApPXkuE8NenrduacSdBVCAllytzfhHrtuth8kI+i9JGoQ9n7Y7mUtT1FMY0I
9/zdmSgczyZqIhtC7bJiTbxoHRJwmmJRyugKkv0RS313LofuKZoj6Y5S/Wec
/2XtfBjOaoM5WFKyXawDEz7/sw/bwdOt8KAtwSU6DxJ9fhVafnpzrZFwmA97
XUDTKkKdZzINk8F18Fa1aGoH9D79sYf8kjbiHDblR0urhte1jJfl94ZHOXbt
k3v6XpsVGkI/lXFPUUvL0cVwuvSmv2rD4e2gfpotzye0Fstz8XjR/guFfi0f
NKfrIHlBRIC8aMgteOWbwOwjLZI586YZyGxuTjF0/eJWHWH4tHhWSgqDc8tJ
1DzCis9Nm2SSHNjG4+bv/vYQDdvq7EjfhIkirJMumg+N0Ev9BMgtafOeP+EV
zpSzqTEIAitCU/AbtUzfNupvKUBsTlRn+9RnQ37A4ixaDQsIjYoCWlbTdZkx
3jVm7YmReNMpjsn1dRUNYybf933lHclKFPZ7TxPyBMf9dXzTvGD75hnG4/FZ
56xN72JkSVuoITL+Qgf/Uhthvy5DpNIyQeugn6X0Chq7hMS3a7sCk35k6ybh
daryQjmUtSV9Hr3Sqtg2VZnVRXVdX4p+zPnrsMyRf+2a9F/QBR3rZbZ9ZpFu
9HhL5fyO4e96akv2294gHOeYklD4DbPDjXyoniaCMDfKyGrd5Rkw0i2OgWNw
6DfMcv4RaJR4XoUE9PYw9qpBCDKm2omNXQMJBW1v6JAbyMNpMoQ/IlGIfxyC
8d/VxZ1FBws6p+x+jX1RSdIb7uVoHMfPLePmKy5/y7tELW73iZjIFCRiaRrn
3oQ80wlbNNd2Ggf5ao1HPOnIAcZfRI4oS1ISxWlb8bBnRbVv2ftpAZBsoBCe
50EFg814mq2bqqCQTksZQGA+8y0FgJ0OcZC33qvpN32JHH0Vjjz1fTCEAEz0
ZtsR2sBdzGFFgDOWg9kGSn/zPhqd3YKhuKHOER5TIAxdE39uADFEV2wd/ivD
EJXUUnjSRcC2V6x0TJkOs8bOHvTccDn+zjxFYkxaxC2yPnzp2/m+y7G4fyt3
3w/kK5QYBIpecLiJTphEdNmat1nOPf7cJI20U+9yYTt9KASYs2r2D7agwVNN
Lyz/UyuSN3+tMX5Ni++DadKZUdQww5id1M49VoFg2/wX4e5scw+Zud1SFcJT
nNDePpI30QpCST6/jyJcGzOv+OM8P4YyPpAlWO2jvKJYsbijRLKLApwMVPhD
GdHPZ7XDqebSUmbchN6JgWr9hl7fPLMFb9w+eU56ssLb7bzovleZD0tA8VbS
8p4+uFR4BPBMzQG4RDDgaJByV+baI0wjbfR0rQdP9m+vPN0uDJg9GJI8N98o
XtT4qKI89MSQIH/bFvC5q7IjxuKLltzQVvXnchxtXMt+D4jDg4VczjxYfsEk
utKLQfMwZO23htztzw+IWdoxy+qEb8z0G/NOwlCkh35cZ00IP/Mgb5lkrPGH
goxrxYBTvA4JsGQsE5tquiQZ5yHWqfoCdI6w7db9yphtB2ol+0JsDzcCUIuG
2m4EAjN58f0VOQZlQDVt752XUxXbtiL5CtayP1anbIHlQJ1qb2duUhcbZzm+
Jwfv3wbXlKvlef7vxp9MOmZXcRptG5v6tSNLLDqPXzGI0IrZ5Kaaouj/dLhO
3DpHGyYPoL3MC5Sa1zGBZIh/RbxGEdfddRvQbGeIC6bXp58sw0CfC7NsUs7I
XlOVi83yfKLxGvfrMoxd8Bl1tb994fPi2VM+jlI2G0jar3zjcOPq+wYc4Iry
ohwvDOZzY/lU3ogybOBQo709NwSspwKRJcpFfFv298Y1h9DkpO3HLWVk5Xkh
PYqFGIlBwHIYYIXhB+NmChPZHfuVmPAV3/1wJHPEQaTFcVYVJm8tAv9UxgMQ
zJ/4ai/q8oHHlYYllSv5wU1B4tDPAvaL/ZwKYCc44gW+hWU+RP6FLZAbTVxL
byZxv1MmxcWm3snher7/yli6xdQZiRPUeZliFxTxQzyfbqfS4yMUARFE0uAA
1RyXaOpv2+JWdt+02tzWCWes9wCTCTMoYTPoMV04Y2N8WOw1OT9px9Go0Xvt
LvpXlzZ78v71LAZK/LA7FWJkdmWoN79iT2SurWbEsVJAmyq7rAz/uWt926k2
kJ8boMP/J2gnY/YxlTyUBXFN0kqvxn++ikbEmaqRj94yOEXviYcL1cNmUIGn
OTayPMOXccpcmHhFp+QEoNdcAMHGgIxuPhPaC7hwfYj8UFg1F/JkC5skZ8Zc
SDrw4w6YiF8FHZd0Knpt27qh80Ezj/zx0RNsdZiE4oLN9IXVh4hfAHHEBA5z
ufFa92O219bsMWhGLrS8ejYv7BFQoQL1vghowSRRFERPiGdqeuCgIGpOyheB
Hflwc5lOb6WbhQ8O1sYU/HD3rwE6NyZ1Eh8mkKmYn+PeZRhk6UivoW/bZsmK
sbV1lP8u9sBpdnDnhiXpf1HMH+sYMEvYOaIR8JMlE0dIEuZyXCMHVb7v3V1+
/sb8DNVV5QxiZMKRhsLsyYnDLs7naiyz5oHKSJlVyOFKPtv5jtdphFNEjiB/
BLp7yMlz7kSG+EEOGBmzVlGtfwR/rOgOjRPUHicBWiOuvzPVT3CundqDRmQG
XemTNnaw6BNdE4dribZIVyNcpyULmII9V7/jDi7Wjsb3NSPmOsbdOjxleq5g
RGG0vL1Yd3+bApmspJ9ooibXu/kemq/SxsHerw5xELG314oaS6vnxYIxw2Oq
AfuoUBrZQd7GZgHkc5SBmBW/Dfy1tTXrn7iCd5XfMsfRQWrVLf0NHiaYCrBc
QMC9gNYA2KvjUjq9YTiEaNCWsKYgia1b6R41HJO+/Fd54CZZ0xNXwlXWuH/c
JmlVpAexkc8DutOez2Dvb0Ff1WsVlScprzGLu5Mqxh2hmgeT91OmCqnsyTNI
P7Xb9RkjnRAmLlcHTip2sVrRYtusMyLdVG+ScGZ7M5809ydwvCg0wUYFAvVW
/MFZIvy2SZvrsDSclFiDzqfHHIJmunHKlU8e4C2nA+bSBv7ROrwqEHUkkTlq
P6ZsuMiuobFf8hqWuQ9g9eKbLDRhEnGYvTyc97JfwHOVJktn6inSfz9/r2fR
BeOPAy7pTCpG6KI8NvQzsg5wmpc/ym30v6h2N5NTfRGAHVc7pddyxw7byCLb
TR8CGuTeOXmBoDhf9zNaxM3ooGN4kNfAE4WYfsgAsWwoXPt03NAx3mSnio4i
NXY5cQ93owajEHPvK8G89z7CsQAHvploSP9apJfoXIa+csEJ2INpMYLrS9D6
sWFW++xJQprGlKTLIQ87dU5eoUiyAnewSYFFUO2QlP7gaQyAg6iTu5J6as1i
vo8EqnaGlUeJrCxw4gmsLuKmDYuFRwbf4NclhYE9QCFFO1zOppHzUmmgWm3a
dCsxV7e9k7scTvHtOkz1nHd1q0oOX1NHCUYi87tZBK6IHjT6rq+PvPhU/mzp
ytRZU198c36yU0FxupwZlqUXbNM6WYfu2LUt1rc6zJ3ce58nI4gDO9iNg0xJ
B6AIUe73zS2y+aW4uyjxvP2sGOgYy6LDeljGEGdUeyeKyJFQci9iNui5JU1o
n+WSjV3xqL1S2CJsHhAnHdsJpiuNBMUqQygy2zLZtZ3SXBvf31hhQ/5tOgvE
aEOIwoI1PY/JodXaBtBieaIssUay547oKQTP8U6A1+STMX+jIk8BinCypPUh
SmARHURxTbyVWRiaekKRJ5WyEKBnfvHvNQBqLQJcHFIG2BstxYafegUcqY5W
4DJO5b7XuYa8H1OnhVzPGJpfp5OrYEy53STEL3nONEex4chaYr1veinqUMEK
DIF+r683vkFOp4/IVhIO1CEPZpEWvh3UCwaN2UOi3/PGR/JSBN6uIZblmilf
gnGvfT+ccoLxSXp51r1bJbxxC0XQI6k0Eaii3kgUi76AKmgp00uF3mtEXFh2
BKkZxjCqoeJHceiMmAn+MvRwQogbIhoYNni6n81iNqFsvBqBPfXHYusU1vzg
tsuQ3EGtwalc83OMDxaYRQnhpksv2J1jf6wmjdapKwfG1r7chB8MJGkIO8es
yKWINQSEJ689k2Db9susRquXgPh7aajXEawGLqWhZnmo07z3XzsKhzcS6jGa
2arqeerEu5YeIMyeyCWNtyRYaWyJRnezfSvFYrr37/FFGlZNrlow5hSwl1J1
1qEDXbZrCVw80svyf32Nr8EduDhJjN2rjhFSiaEp3LaG82xLbDZnExfcdayU
9Qbvgmw6rllcfMmgjX+bF97oUNW5jQuwp5jQ9aU3m5tQb6M9G8ib5AFGpQjp
FlBSbw69TOZHK8LtxjvCx1+5b1q7yfGODwGPmlRkIA2XjQsKxbJgbuw+t9bQ
jjKs/yVei/4O2ngNOfFgI6+vkww30W9KFOKWIe18nUW9CRTdzly4UN/KzYSp
klwMD6AdiT+QeMtjBjYKTcR7L26ThfA1ypQESworMlGdHl6++ZwNhysJFoIH
618H8xvqm8lIBr47lHZjUUbQAfihpuHJ0JnEfRhZiSLHG4p3O/f/mfWYCMph
VKgwyKot/EaVsRF+aMPZ0lUs/0/NSqA3FopLkoMgqYNTt03DQT+hTsEAXEyz
FUvJ1kdweuT1CIkY0/LzHox0Spq4q7YBQMtvG+V5w7hShNmBZvSyEthpAlZh
TH38sfKQ9lxAONLGuZCYMh+A12wnY/mArU+4HnBy3K5Pm6MB2OSuNU0AqCYa
1q4t71QuBMgtuIbJalmdO+e90FIHrc0zi8g0kYmSHllDjbtA1qSkSPG+o0aI
0GZ7oWM8C+w9DSjHirFkzbARyPu4AOhLvUo5ogSOsrY63nTtWIPFuemtwc9e
cwFlg4BOIZJPzUebAbpIGT+5sDxk3EdP7HgI8I56PeJ/uDr4K2eYlzSLL4ZG
yVXynbVZJ57j3BbUISdd2jmQA06n4udycMJT+1nUxX0sXb21huw5I1xygPoQ
HNFeayf6CCqIuqZY44omoiI+cFURMSKGEw2wAqDezIo6fVoudK7+qIEG5Wka
DZ49yCEVTJkqBMBMj7U6Cict1otLDpl59tIzalviRrDvEycjsI/vhQiPOwo3
ZdLiTnUpAZpmAgwe1UUxa+qUgwz68yturnXBZ9fKOItKJpalQSK0U9AyMfRg
5ursEnvJzGkuFaAsCML9hvin/yL8Y+G1/CZYEq9ZjQDjn/ghkBP2YcisIi5z
DB3bXhY8zq27fxF7AsN2PUCnMHrvyIHx61keIdhXtpJGd3twHjnmFaFEXOOD
SzvVy22QX7juDK6Zb5UvYTawqw7oz2xijDkFJtkV9jSPyey4RRa3yxXDIfk3
f2GYXMxhM5OPw2quHTJkqzeALeVU5W2uxVmnboxN23eHjBeW05yYZZqwRBxg
FEUPbfwLPZ0LLUduLKUf9B+9RmIbD8ydl6pTmFHoB2nVHBGIZsvAFlGkr+WH
TQCFDX51EsfMcUhYXCIqODgw8JdIxX/Sro5nV5HWzkN0jjMRmlXaQFsNUqen
vTsved56chK7zxcznwASLajwC54prgrnXvGByXjJexvBRht4UnSknE9ss8/3
buHffj57s28SWpzavhJ2vNpuV1kazJ9d3fL2qqOTlllGqbQ29rbCNGu81OUE
yKWLshLWocA65tTCdwAMfvkQu7QQZRQ1t1hESb6EHtLWO/2HZOH0bD8tNHI+
zyIc6HgXw1XWTHtu8IZ3HgVWF1Kdh7oR/beVXZ6pyQ3KuYpWRr1MOFAE7N+C
pJwzAvvNJF0WIpq/im7kuLS06VK+3A3iV/vcYi1ycA824fcTSF2B0WiM0A10
CaJi0Uug5OcdmyZWE97ZbENSLJ5tlYY9qKzCue137ERbnTFqnGkhr/0ODNBq
p6qsPyH0yCBP0B6jYVCR1eC1lHtyaeFlR2o9m6PF8lErq2V/YSJPJufV3jxP
kq4weAGCXVzwxz9l+IIjWEUVUMidt742Pk88atneaAUkZ1WbsPOi4g1Zr5T4
V5jDEdaqKg7IW6kmdWRSLuOCE//kMxy14vCHyv5h76cdePGKfAY8fsKZeISM
c7mdvIgk6+P6PWMuRbMNbOMhr2ppxZAvj9AC8O7rRnbm7rktU9qiUouc2lKq
x0Nuem88//XSa0cmqgSHK159/yQhI56oq46FrUTXSd62+pXKFp62VSiBRBiZ
hakDHt98QqV2AvBLZvVPFH4P/eG08JNFSYpZpaJpPudVJdosqbJzoP8Ql0zV
o8VB6Ok4uHhtpqUIWbscEeKaHMxsjZ6Lt+tguPx+4+VhzHAEbQQwMrGHuo8W
TfI7lVf+yL5aK0naQjCqUgg7UeGWmi92CWK2zZG/9KEV77KtJZo+BTiUdQK4
wCofoInxJjVFHRaHzKGzqQ7X8jYLg5eJgWYq7sobML5MbZkeUFq9kfW7ft9b
O93tsdvQom7aQd2biL7SDR8qUpfoMFMxNVsZkUKv+d+BjtG4s/SKWFa1wvF6
9u/zN0Zx6Rb7WHPjAs+LG8Oc+MSYsQR9qjQAyt6iw3SFOmyGe3gK74JkUePN
vu+KHIXrcKCJu6Br1HJQkhZ118livUV2ASBTHTcPOh1MZXskcB9998B2w3pA
12eqV5f3DyulZtTIJiMxCc0m8mV3hRefLyWatquwW44ESW012kPkaG9bcgeF
G96rnkFiVAAYVWBPFvF911fs8eT0YqgylVYkxhTr78MC7IEa9Dgmj3SZQQGg
9Zvxrv43nAPYqi/YH4hZ0HGDMc/Bjvd6aishovVQs3ituuaNYuqr0zE/5xxt
gYzvYfeGI2YKSI3HDVLgqlkXOCGeSUalpprM1wzYvwXSn3QypzvKOnrYJY57
i8ITswGY/v1Yg+etz5E2uyVihf8hVe1K1DrmZqfaxU6KYKsZZN6/969le95i
w/rKE3gxFm6miHTp9Z1p815d/nDwcPpTMr/LWtVJjgZBoU+QBPpvwo3WeMXP
itqbRMShhxEnkDYMYO/kk4CHgWBPqdOW9haROXJ5HjEYfeZwb31BAawKQv79
Af3uZcsplED9zVhsAqyjZN+Kz+1+1NAIIVoxAfGCt/n3/7e0NjySdthVRxca
tcAIKWG9aNi1f3FT/y56TsnaT9WULrCvnVF1iNGF7xV5Aq/yeh2FX/bw+wsP
4cajrxmMOwD+M4FDZq+i7gemtXYdFzwgQbZWa+89itPxo4UadE6tGmIq28cK
jE3dEyfvjGRJMDNym/9N7Kk1gaa7/TbEAJtXKYIm8OtnoM8t63KMmreiQt4C
giJct3Ij/uAOgikw6/YszWIgvPPJZhzZM9tKjkg9ZypcaQzhV0cPp/u+8nTV
lU13uxSDiF3T6oxtOZqOoxRDSiUQr3p7P/k/aVlIJLeiS5p8xPwsWmI0jDRS
RAv58gLBeRkm5eSePce6IRNljWwDWzmfJWasHxHJPUI2+lNODGytY/xMO5r7
Fb7aSg4s3K9fbxFOBYeTFWKdj/C/esRN3TFJm9smDAI5PxyLZnXkDV9FO121
rjxS2hHfhLdHwNZcz9Y9lwCsVMPz1rR3GgaS6fU0xyPSnMgPCPcz8HVX01WD
sGSoJdIRsG3FKVS7ZT3lvJsnKsz70ESpL6NSfn2YpEXcR9sBSMkuYfuIyvU3
SfZFAbzAcIxypyo07ElqOBStudk3umwkldJ09jK5/iZ3Fz1ONEnhYNCGd5eb
0j+masuzIiVp9FQkhQnEsCvjGAnCU8g7xWW1Wt3EZbNhHCrM0P9/1EE/9Xfh
DzzPcewHrXMXPuYHu466y1G0KOXizyye3OTYekr/BlJtVjTr3T1/FemPsgPv
Ba6LJPkpllzOZqkowW1jMmvf7wx0rVYWyC0tEM4Qwufi27GT/VyJEZoLiNQ+
wNjYugQ1D0J+fQaQM+l9xz+WOEPKmHWxQNrVq92ErHi6+qWksqyapncgw/zJ
mdO3FmjxGKtLHuBcXZsq/qrz+Lp4vfPYF0fVo90sNUYMVHxenEsLOL7mk8hM
Mf+hkr6PjnvTRFVG27QA5GuOQ+iVU83qBLaz6yWVJ6cWMF+/E31A6FMo+5AN
SrV6kNgCIMwyvkvYt+kOQwemr0qs/KUVHF453QoyLQaRNZKzeWPgBlExzgQB
B4YVmHEAje6Aelh9TF3cqOb00ABPeGbkQ2llI2CLLUWB3tRNrSnqHfOqGpnJ
TZcKmqy1OZRcpNy4BC1aDfJYibNKsAY4QUM77wtXMaY+zyk1FdmMviPLz6e3
U1MjauLIh7TELt19xtxyZoIYIo7JrTF93ZGqRPstEkunwNzoDON+Z0+d0Yt6
7Eqt1MPo2FCH4JFP1f3KT8zCP8YGZYWF3pMBc+1oD5X4xDX3jIjkeZuMPyR+
MEFyT0ZKpufmewMQ9FQDPyGGYeocYe6u7H50RQ1L7MwAAkjAxirqxn66aIoM
cleZvY79Q7OpErcaCA7u78ojMrUYSobsf9oCX/yjuXbvIKnh0NQQbOtJE3ZK
8RGIbIiOKJZo34MPT6OGAijNXolg0aheZThnYeMHyaphQXHAX3CHAMFM6xkL
Mhqh2fVawZWe5Y0ka/NW75OT3VTFlfGV4Aa9eNr1790q0PAapQliB4vIr6HP
4s0kfq4kt3guHx+K9c6xslWKRQbMLb7/4ueQcMgxK+zlbsS+/zpZBgkvqYDS
kjGSO09qWqkWGASQTWRe8V0Uqzh5XF85L77ZwTRYgAGUy1UDxhra9YB8dDMy
zpATEC+/1kEZvWXrx201gg0MLrQEuBORmkogtdHHZ0PObRIRigdkltNvoaVD
wZO3iXvZ7eK9t9zW0VagLsizJ1TSotKUnKc39FVOMOTumuwh3jLo/UTxmVZn
/m5a8Mq8PhukWFbqjIGlQXbHzpV7+1MdFiSZnfCSq4eOiXfg8bTRMbiPhHw5
8jRRl/pk+VRQ7SLGYoQuLY+DWxXDcDAwCZX+E+/eiiZyW9AxMEN4UXSnV9YM
jGOhIAmboeFQFljNNvAZ8qjPdj7PP+MdzeoxW3yeQSmD735QNbGSvALF7yGF
+Jtil1ne/g6aA/+ae2pkkgZ/7Fj6z3oW01Myx7+yshY22UoR9bDNDzbWlYZ9
TCq4EqivqhOMB0CL5TEPLInzncmrTCEEs41DSZRA3fT9ujz0aJp6J2SVCzlU
gCY5EsVHpY5vlcyX0Jf/Ki13RSy8WZyZBvyLNMQttbvhcjaLeEqb0nO78Sxg
QETwMjv+xhboP+72Cy+1hOglhTkXv25oUCaSGe2+5PcuOgh9legJc8o2R/gt
ta7NQMj/4NWMwzPZzU1wVVBZtuA2d9O1cMj2fG6fWQpD7YzAxAh+U0gyjrXF
0fuPAGsTKJGmNa8EjVZgHVGs87MATdE8KAZgIVG1cECENNINJNpY1L5YEv3q
iZHJku+nJsLp7Sux+vLJY7nj1jIaqD5PtBeiWB8Bd0WZEvBNALKkz/6DDvDi
J17NjX5Bnq3Ays7POCBA+a/WXsHKuSptNjm89ra+FbBMHmSUEcfYqkwp47F6
jZth4WVaomgLetf0GJnDNTxNAjEEOs/dJ1nHu4DEKAzZB0CU0RVMN/B6svia
8+xdpNyVBDPKOCN6/5s+raFGTBp239d7M4FF96/3Fykqn1rR2b9CFXZzmZSZ
/WHeuip9HbJaidUySeqeD+n44/dDVJy4gigtj2gmbXnweTe6sVRHvnMBvtJw
GI71jrGkYBwzxHD8JkHNo+jomhkr1/7zBsI6FyEAtXz4WiqBwQmddbr9ecgY
XMEIu6OlsY3mEyF3PgE2hfmNdBynd3ZWks/N3s/uAu0fJ6EyllJdz/eCFLR5
TGDAHkjbYxGE6kectt40t/V7Mf5d3F6/ivrRVJTyjWOeRHAxK1tXhc2y/MuX
FMQy8y6pt/qfGCOG4ZiIKVzgKwgFvhpTbmexxE1NkJC3BRd3UhSFanoYdqsS
e5zHghntd1U8deHsYGBYbfcJpE4GeTt3ZNPgcC/f2XBG2Xa/ykFCfLct/mmr
zQ4WYFnM4gzXpQd3BsxDKapX2p9pfohJcfNzoDccAiCghru5cOFZ1Fq96Q+s
jf/lbPUB1QvJEvPkVdFxy/Fq2um/zVIYqi8bBFEgoredhmmJbYAQ/1HLENHK
SdILHqiy6oaRz2S16QZZLIzAhd3Ci5eJMlIo7/Jo/YQOOxFGQqa0nJeIKOAi
ZPxn3er4fOPSc4OT3Vqjv6/TSgU0zGzUndDDEdhA/U4Gu221hOA6UlBPzlZw
32XZEtRcuj/KJUzmyVeOfYUUZy0sbk4EkliPGecKt2OQ0FuFMGdsdaoe18v4
z5TztE4tw/BI6EvpvaZaZK5zvns+A/s4//QmLbt+PR/d+qMFWy6j6akJPYbF
AHu8iwdpCAD7N41OiVCjfbeS1qIYhZ2NJU/GeCEPKVioJAWBbv8aV7QUxJXk
YKB8FtpxrWwRvlQ4Pn2CZOFd3kWMohFJwh45FRBh4SsbCAhEyarfw2horOOH
/d9JCJO3NajPnyO5hfMxl+UXZERTkKWAfafNf1esZLr1/JGt53VCabXUYG4+
a1L/MvCD0PXK6DxJ6xN+cEWmki8IRoYOMyVKnE7raRg8gZwWxgD/YIXHxFPI
W/jnx6imYjHLOBvtoV8dQClOo5LFYbCRldsXi91dtuZ22CJNpkOh1T1+gDRw
zEIHu7qb2F4SinxN00uz7HVisoDbYk6Qq8Ak0TPqiXQ1BlVyArU/YY3gqTxt
nhIQe13SoMErBp31frZN4c/zb9BQyf7opViISr4nGVzrYVdCkXFI9y2TzDht
4qX4FcdKNwafArTnZ48FKlYL/+qSjuavqRKMelbhQ+uvxqSSOaNJqfzDUFP4
kww4P4gYTlClZyCuxBV9ahagl6wk8tt0B/ldbXnagvC20gMsHEUdwgqDzxJa
LSTTF3nTdUAIjBdBm2P2TITtb3KCRmnLcCoBv/Y6a3zHG55Ifw5ix3UQ2JqL
E0pq2mp4C9KF7+A4/Hyw+ve5tm1VRueU9hpFHYoTintoLHUIaOv2mSWAvLzk
/tQt0B18m9/26znOy++cxk9z9ikcTexI3A5wpH6AdOhWyDbx2SmSJ7rl2/wq
QKfm7N9/aOQ11qKoyj6OqKlyKR81p95rYqhmYqWVpEzocfL2NbrdgxoLWP1t
/HlG8Sjr9KQ1jsiDpsxGio/rCj8xViC5z5c6h/mxK+uL+1OCuBSdia2DcaYi
ipWpXJCgnTLurlgKOy/A6hW4paYppeORGjknYPT6VF0cfdfsrOk2bqqB+Pwi
PZ+uAttfilBf8YSwuW7+SXf0b4LqLRhTRyCPWJKMbpJjY12kyoPe2CWxKGEK
PH0NmVrjZxLYGsgbgKMf0hBU7hDTy+ixD51uOlJrGrn2x5wqTGcjtUKA0I8d
YpZzhNvq1uFArZFLbN2DCCaoM/dVuy853KtvDFAehIKF5rBTSPQJ3spLwmGL
ul8edkV27mppRlvndsIhVkRBVC2IIEW8ajbNHbsOQHDEZg1jLXITxgKDODKH
TEI62AcsmRCsBMIBbK2DQgF2GWzPH5IAxEGYfVvzonx/Mc5+WOraOS4nzPsQ
YuHmvX/gFg0tTXhc1mpmlOfDqrLDTo6PICgJUg3/QqjZH5WTi5FkNYD6OaVa
zvciNGdWhU8fBHcG/KNCAlc3y4MTI8f9y+zzkO0ujq61pOshcIGGrmq6tt57
TPovhH3PEsAYyG0AkHvAwQfG09vlu+DoQHSarHoPClzssClDT9ZU4cOzy3PX
i3GFoxN3Tee10oKpBokyS1RZRHOD9JArb0Dctqm/X9ZZ4JSfV03Fb/GV6yST
BwSWZVNqU2L2CyRoWJCNgYwPeDoB8eXvCOMk5trTTY/ZQGhLtnmh5CDohrtg
FtBs+17ECSxqDgjh72eOHkZZUWWIZdxEiRvxXWTQqFI/Mj6Gly5Uo+TyZMnX
8MXuSh9tWTxBKIMvtkbnDSCylrSy2AW8EaJGEKwgL4L9bvCwfYx8jfYZKiu/
YanmrzwffIFl3smxace35KNc+5/K0r1O5JzfP94654xt+MLpbPeR7CJeRTlg
aXb1IFeQ49+1uscG3Lexs2Sfw1yXRrdmh6mQuVchhHxwAWcgJU3C3v4oAdBw
yDss+SouyF+qITqWJP46W9nXj+wTfqIsKrHr0mTQUumJapvGDnIQBcFp4W+b
WVJWdsNXqLiMfhcvS0sfjupEkE1hmBBZv7/eElkvW3XPYAnzAcH50AOWjBpB
Hof326S6jxi9swybpM8ZM61r5/WVy6CH9fdCp7AODx+cu9OEnKjjYSGcixQx
ciwa+RA443jp8y4MGS4FjeiEGZNftwM4hZ5Ng4biYw9MIZxGYsEbOoZmQu0Q
GC8FkzAd6dw7fgjTZTf8lE5H92ZnIQfbuy8ItmUeTrXgB7aUtL67Cpcbbivi
lAa96fHGWUqa2WYtz95+j9x1zj9mrcOR9CSZE8Gp44XqvN6PDRIkhor+QIbK
VqkfaNpnnP29AH4UnhTDELuHA4nlmOkjRTMRxcoQguO+Ys2yNq4shQNWuow3
TjXXQJJPLkPYnGMRszOoFn2rtmSXoyVDUz9NPsshx9bpnCC9uH8rs76M/EHZ
pXc7HYeeN7MtYID7ws0xoebtpojyU+T0dMcrim8WgOCkYFNKudYJOVjBpgVK
NQVdidBhxLUDkdlHb7mU3xNRd2XF4m/yGDmrWt5qEziqYiusgziXnrhSxmXd
qWHsgyvnauMKRfBDXefw9uBgGKJLNSa9Ky565v9d9ms3mHFYodhJm/Cpz/E3
fB/0Lyq+ERcT6cxk0B5pijJHwGgnuOG8Y18NbJI/XZBDaZgpsvoVXyoFkbBB
s0nqdSKHHjCgAwul8WMCN8e9dexI0t/rbEVl0tZ/qHvVtORLGVmvGnufnvJv
6CO4+fbU+j0wF8RrYAjGGFEP0j99T8iKKilbV1G48rFiGQrmPlSgZE74nBT2
AohWkh3uAImHwEBM2O0f8d3GIgoq4drLNkQxMlCqi5o4rqlN7M7r2y3Ff6hQ
8FqInDlPELNzoQWDWyxl1DCPgUSokuzOteDaYCT4uA6cXUhDrpQ/qz6CvlVd
iYYksqaCoo1mlomd78cDIhvWGCZTK265Lo/lXbBegKsNCi/VEhuxyGBv/KDh
rkdyNvG7G/LxPonL4SVeXRAoeZ48bu2iz0hj+O5MhyTQrWUJ80X+Kjr+72Eo
ezNXT9pLAspXPhJBx+Y/BUZQmIXTzD6DajWYNecId1OMo4DTyfDqn37Peo4t
eiDp0F4iyuuGe+5rWpIWWEkI8NBcZjT1aJSB28xrA1O5w6I9p4R0B8foM/SB
Zrx+HtBTRp9Jco62RafR5+Fj5re26T7QaNvlZ7nFsINZOVFFjHWKV1BcnITr
Ot4O/kW+pjhD3towRKSmos+Q4Ji4umkj07Uzs2OtqA9acnZlwgttlsrQmK8e
FZMtigC+g2g0NdyV4f8HwEcsOjYK3W/oeTtnuEMR4pbdmTPpRkYeBCnHEaTB
NGp+HAe+/vZ6I6TpORapzFVp8J2QuB5ShlCZSO2XHfsHPVb/VZJrU8Iafb/f
ZgnoHgOJXw1Xjx6+MUQnnhJKQmorJErz0dCYOBQ03iUV6kIYn1+7IDQRRGAh
7r9VSwRed0jabv4OuDj5MI7pPJiwHiA9DporTdu3CMa5u42D+nHR1xRg+CKb
U/7r399qCA60cCQwUTmiOsXPjs2lR2BQB8yMGWadjHoWwwH+fnlGqyoHqxr6
VQLQME7HQGNjJfWSoFJ/VrdS8sjjaHsDwwTx2QgdYlsKgjxlo7bA+1EZUhHw
UCLw9cNkaRZlHsH9U3LQ/K/7zAv4kdFKMN1GzOjQu83pX3r91QsaYkszxdGc
+6CHoVKdXHVC+IMKx9wMOr5pzR9ilGNbeqgVkirj4rtVHR0rHUXoYQDMhexA
ZWm3neA5/s6cF5eQcahqqU/5whrp6c4k++22jg4K+kIzNz8HWRhTseXVin8d
vdDK2/dfzRKlJb38bw2dQH13uV+29q2g3ysZ9UpMQnIIH0/KNKBn4YosjjNu
Gh2czJn+57K/NtkYOKATC5BEePAsEpuaghu6xx6X1l8yHX5IZcSepRvtNDiu
rYShXUqBqo7tqmL0xD/x+dijMVg3i5ybDhZWGO9yGgbOgT7XV+KR1WQk0ZPk
i3w+IbHs8j5/DGUxbfIeuWapz+KmwnWzgWfsM46LO2/jyvk27CUoF9T/rhFV
EDfPFnsFgBOlsSh7lVU3Gw2TH1x3IRzRcrE+qKNJqA0333KfTYU7QMV8v1Ac
l7BrGP+1zlQ2IDr9tMkzcUOI8N6FBahRVkbeLi6d3B3p1HMR8hWl3bLEFcG8
cyCPF/zW9a0hbSYRfVsUyoAkf5S34eTep4K8AtKjqQgvl4yDy4m4V270aLfN
MqMUk7+cANEaUopYu4zJbR493BUR0Rnv2tmMrjcYIACPK1eWzUNR4xamYmTw
m9wmxjXMswAcOx7W7gPvOnp3nwc/91TVrXgx3A0zaVJUufZ1J4SG5ggrIMh5
P6dRxi+BR8MDD+nEoTtJB9bUxtmOJ03VR6sx1tg/00K/rOhQ/VP/W67uJ1jr
jZWkcCztHLpStXLYPCOUL6N//B6DQEmAsVaXsDIvOETkmtPtNn44cN8VgXwu
vItFrOrO7eRnLKTXhUgGEbP/n1zTEFiwJgwVydeNsRulj2PbzCoFsZkTYGSf
Gv4K/qztB4Pz9o7Gmf2CGNiez4AKb9+yr81sIhiddszl5vY+LHD/8odRGxXM
AQgXeND9URE+la9jvekCbv0dvxp46sil4x3FAehLGx5Yr8N1TQ9aisWb7DVo
RCLXVs4cygQW8Cf3+G/h6F1/CZrdm9SJ8cG8ah4uMwpwa86dT2GTrpTbRYdz
cZi3zKCJ7yS64grvc6H8D6s0dlFbTTZt2AhF3/8JmarGhX4sumwUR3ngFJHo
NwA4vs4YWQBVGeyotZIx/mWchuRj/2A6jx9LOGMsTshHb5mrSTPWLtevKd0T
ieDRHjMrwGv9PT5lgtNcSKr5XjIJ6+V7eRw4s9nG4LCXngwRLHLES6jxiLtj
ud4Rf13EZ2cJTEr91EXBvx8abTUidbdjksJ/W0xgQkEmE9nQmz/II06DPpHF
m1+KbItd+tnRV0V287OcEW+SGttogHpukd7OMGD5GtXiY88ml3QkPnpggL/m
fQU6pk6QLDEqVI8F9rW9POC7tMduduBYFci/RF5HpU6mkB8oj0xPme2OLyiB
0Erdq/oTz2OnN0G6XfjakXXhwFP+2MhZ/s6Uu20+A8vh9R7BlEQPux3JfIOz
35H8eCgsAsttIRfTsIaCQFhanp2D5cDEXtImhzYeWNUDTf2yzBFdVgSuBye+
TMaJS8wAVJZJYU1B0WZHlHhPPOH1begDBFH0ZUxcKO4zlC2GfH2mINQVIHwf
Oqn5nSLZoSYep6TT+Wdnl9JsbBuCCygnwnwya8YYQO1uEx96nLANh/UWsJyu
qMA1n9+jw8UGaQ9cYvvegnvnjWSdry6hQKf3wq+dzPJ7EJTYbUpgzSeP5+Oc
9N43hwqnJ/6N49DyuEijM1Lud5sKEcnSoot6bI+v9uTwhGs2PZni/cxOLQaQ
Dbt8SaymRjdNVs7ARiUe4uOW8N8Szr+YVLjMv3HaVpRBKOa86h3tLXMzV/45
Du40vChVuOVAFhz0KGp7AYYS8fpep85M6ukiJjB2XjMrUiggF1dzqDG03Qlo
T6JxtYJsg4WrCEh4McNJhvZT7KPrb/nBRXDGLy7EWPVGS1OOncCKZvUCaztK
srO1/rdUT06vj1dbChvEAa7NQtpFfVZexZ5EImZ0lInW5hc7wP5Y0ZdwxfHx
I/8OpPNA4chB0Pk2QstVYbyIpQDa2JuHquH5fpUPWw+yQu4J1wAyzlgt2Hlk
/MBYtZa/oi2edYiHYv2FRAXuKNq7l+pJ/g3+Y/sNeVGziNUBBWbaGmOcUk/w
p4bITtYNt6GI418onbtCzHm2l0AO5lJ7BgtR8i9es8pwaIR4fExeMjoOoS+f
omKa+SlUNCRz2N71pWD+cSYk/lB/wQxmZTh5YtIqwZuCKFkyDbGl7neif2X/
vso9XrXYnVA/mZXwmW2Vuv99P9LNgpaFVQuod+wCQfmxNFZg+GNuOUxDhPWn
/097Nd+BGVxEOINmIyMOhCxrq1wKo/olcD6BZ4JWSomtE3m2E5TC2bun/OnL
vozdIQCH+isN26YB1y2c+xgqyL7r7nlSzY8kITz3kz0ooIrMCUbU4clLOUF0
Kev42wIIMBOLGFRcRDtJuiHa0PMw4tMCQZ6Rk76XoIX6EwRxElMNqhW1Rirz
mKjek0Yv+qGzQObCUEBDi0J6Ec+MqxfQI3kzHLkkowKhmE/qoEb4zqTvWE0B
X9xrb4YFbcGMZA7SBQBAiPybC8wOIq/VuDNt62+VI5zzOjC9BYWS4nsPaSXT
HKoQkuEcemAJjnlFAukAYcRtRGyHpTkh82ZqqmxApla/z/hTE5U8LRtg93Mz
M5UK5J5RrMVHBKI0KDRonLexPGryMkoXolATnoHz9xBkJ30EVp56rqFkwxpc
BhUzSEfC9m25WOQ4MpBaapZrza3YFXg20KiMeOnuvflskxmJa0denwssewkz
qe8jre6EXjkddjGbHnfuZaVoX/xJgkvjESlcIlB+4nEBvxLqjxehxjqWQBvk
sfURhf6gDLyfE1S++DkEBA0y5SLA1HtqmryJiLBUCmZkZN3MAVO7bhdEnAiz
uo5pugNLAHyd7YDKGmc98RZeNmlcsmF+E8d8syeiJU7AXjBaC2Vr+npIMrZn
azPMVJHrKOWmrBLxt97e3dNkLrH3kK1GQVE3vKw8/PcgsvjHdxMgps5b1Hj2
uxhkToEZiDpDYlNvZ5smHxX5P0QhuqJAk9+1qUMjDuwrlDMHvMXMn/7NQLPV
8qpfQGnrzMbBysUkoesI04PR55v2KzpA+HwJLzj29oxlKJ5fIzI3YbeVSHcg
E4FRY1UOfvSENLaJEPH548fiG0olh47CFG9P141+XnQYrAECJOS9maWzDW+M
PJMSOalzXQ5JzVKByGTzC8IyZPpXki/sMm8vaS6wxTGZbQrp4q9blpRdNsTT
x0CKzeMTSSk8egnwQA5cvRMzr+B+kfdDgDuRIT1fB3sVuPRYPgjHx9LvdN+Q
OAB49s52zZ4oAXK/+ls65pii9pU1wGkKdqaFhOfskf4dS1I8FFgv6Axcdro7
nyJ+vdNDnuj6hy7fAULfwzJ5Xx2g60G1oxcFAnttRQlKtrAROY1f+518eMVR
tzrikn2N63Kxo54lrq/VnUhEGZWY/yn8h55waFk16is01FInyPiTrmwCU3mr
47fkFByFaqVTeOaTLqT9Ur/1OuuTdWWck9K2NouKv6mh8oHAdMkzNRA3PGd4
7EW6dvWpLLEQ17y38ZsPvGy8BKowLiIBVbyDFoc1Jsyk13L/26+wPgEmlVyZ
VGVN0JJkRJ8+hNRn14RZlpp7QNvU7fXh2vMe7poQ2qvzrwhwvb3yB8Mm1lW9
Kc6sRxaQWCdZoiRA18Mt4oIo/V7q3fheWMprqElACt0Tts1otqlTn7TT7WpQ
w7KDeq66TuBvrRBt+CB826oDZZ1Izm7Ux6ZYq/ggqxjC0E47rtUiCLxpLfGm
PvyCKO88y7CtSE2702AGtHSXaoH9cgQdGMzd01CelMs+GvhPKJun+gpc1G9I
cHi7Lt3aFv7JN1oMnXaNwaQoRZUMPk0M+ptkjLPzis+F8bwl4lSpMMk3PNvn
GAdDRZ5zNYwFlwE9+IgY07XXZcbNfReMYLq4jwPe0tTfaSJQWZfM89Mk0fUZ
l9BZ108J/pM/vPp8WO+eiSreLDl2Nn0gM3n+UwD/YRO1A4R1b0Z6qUQZZisO
fxlbgWyS0aFb7MeqKf4B9A0yyDcsGeHVNPbxCxLDhFLdRCg2oSQ6nGB7F8sD
ovWZMqSbiUwirocQ8aRtz6JAJGPA3G4nmpYGXUhMAZHnr7/9AygcWwi0OdHG
Illxu1v0A7YnAu/bl04OkW+JK/tASrm8p4OMLnRdq10bRev1vBT4IxyB+JP6
ISSBE9wPWvQgJ8nwrzai18x4BzfR/AFpYuWcoUda25LlphxGiEg/WOx+c8CS
SexXUNSy69brR2qi/jtdZAPtNXcik79uj0+a9OvU0uID5Hu9xuOdEhK8OPiR
gIWaKId60GBYeKiJtRz33MwtyrBBP4+sstveCa9IPKkWDSzQXb88P9TDKfoQ
1x+sV4KyoebX/33WvlVBi8tuj5Usm8ghFyjsGK0DLfHHAWWwVzfUFHLGIZf7
LZD4Z+V/r6WcRMv6dHwdeKhWtFihyijPGD4pH4OMZ5ashsUIX2k/L0h71S+S
jKvsPX/I1rfu8WpoDMcI0qMhieXVAjBVO5Ugk6x0pw2lG6bg0AfOdCqmvt0M
wzMPTjWxuDjYI+KeI3VHKx7G1hmS0iDOCqzXTLeIwTGs1XspYwjhUB0+1ktV
j2paGbRRmHN5rHWO3Vc2rZNAXdnhEB1cgOhELBC2B1n8qA0CaSzKQQZtS6RN
7zaSWjD/1Aa4ll6jOOCAuxRHmTWQrZeW+isS7jUIpknQpwdxGsJ5oRhKuP31
AwHbjydAWCfj2KXDqhdT1N7ZYPTibeDet5AynKwb7u+RRJsF2uJx5pMvbhMB
c+CwBiDQ4ZyPnIOLgwZDnUgEWAy7dAcqRWlkQZpG20CsU0qvvoBck52tRt+/
U3XAdC7T15Lir+l5Ei2cz4ixfKYPzTWf9VKnePPPI5IKhRtoeHGLbtKhg8ae
QHExtkHKriaK81dIhojM4z0R1W9Ha8PEbSGDVGwnFxuhGgDSA/YOa334BKlg
L+kS3UF7Dqf1TIa7+ZN/B7fnzQmw6PbJ+ycUXshD86YDhmDoYcz0iZvCCTGL
D+3BB/nzQ+PSWi0j/ZUV7mkXwNqjKLlcXqIryWRDyJYQ5d+xYxyEFBrzRyRv
U5x5rLQJTtcboq/k0L/GtN6Cw7Q/GjLwyTsS6KgeLFOEtTVhI6nlpHxp+/pq
rw33e9CaO0opwC80qXtDyQl+XAol+yp7GFtVZV01u7tZXeeI4CYueAyqYrY+
nKQhvH7YM13/FlB41aL2TIlrhhY9Wa4TaGu2DVkdn6RGzKTaWReyR4CMDsZI
8djoOGrD28v5eobHiWPr2lT7/EZLWdyWnsS0VJymrla28ZaoRKCheiMdAVP4
nl9RKXK59PEct2G/X93ZD6ZoiFND7OEoeh+ZRUBQENqJK1x8EQO4LX5HIlZP
9yj5mGUFh/FJpCnXBSE0V+awvuRy63ED0clZZbcjHX14vVnWRnFLEfwEw0ks
4bnbn6Is7HCrbzPx68jQZx2CrkpfzMlMWNR42ymZzm/Wo7cwkcw99VnzPPSu
eaxpEajUJ2I3H5ZlGuX+GeFipD6u9h723R8kgrNBZY4tbPaJ1RXMoa5aiaXT
pCbGTbn2uy8vA1ssYTvDFA0mJwWOFjS1ujpil53Yigp8LTWS1M0O0dIx/t84
L2O733QLsZ7g1NiwOQ7ErbdG6PrDHpUd/3SuXs7g0wAz2BQUtzsUk98no5TC
kaPKSBG4hqeb3X3t+uC2Hp0LbN2unMBi4+uhephGrih3W+d0nwtN4MNdVgMb
dWMdtTfkcGy2CIV7ARXkOsqdg0lqJ5BWiiWceEDvmotdFqhlcdy6/m8ebY/k
n/6PVf0JxcmfDU/7Brv+fGq7+bto2mAob91WpYTbsFjhrYtCoQYXOu+Op5ri
PIB83PORnGOD7wo2v4GClJd11+5bzPws6b5bSZj2zMQsatG+pqYJrbyJQzKy
FE9KExrTgbtgJpZGSPeuA9WJUbSsa7ALC/l8PN+cQ6Y1zhqiTUGOOoxkCiUi
h5JljgdWgNn98ujuVr8XSBG3lGCSYekvQv4GOAG5LAO/7ORqztLcAG6BdvWs
vBqvQOorvdX0ZAEb9Lb/H1wrPVXmgEsGEIWubIDvurAU7H4ywFPBaK7iIC4E
AuIoG2EweJC91UgRhL+AGH0Us5Kt7LTKxuhIQ9yTtoZWgFVzbVdii3/FSa4O
DeFUOaIkYM27zNj9AzUEZffMP5eJQPsaGJprE0DNIKNNbrd5x/Tr8ZjOgrPD
dT7AWVAk+Rod/uZWXgB1wADDl/9J1oEE0e5f04I6UyQ5IrPml17/O2C/zntz
g/JqGDgvVj4KBi2UebV0QedZVb/RXxdPmkOjbhgsv/B3gQo1FYEv3ySR9087
xNfoETf551p3jLkAIMMlJN5J5qWtEfIUyqxdcnA8kafzVRpu7mC0r3m5uJ1/
hpsmMbWrTA61t4BKQsN31qgmykO/2V7ayzgJ4jeAtGvuu603DMhLN4qnC+Tl
H9W+tmb99dS6d0uF+H1R94pOFO9H/oM0EfSwzLHDGaNvtr6K2BY64bgMPbwG
DLBJzMzM0kCuuKdSji9/gXFHZdrwxma6LXZ4W8TBIK8LcD4b1LUpAgxFeyBH
KWC8ZnDhPryBNWrKUo2DGLrrhC5f/2MbyTCWgWdb7/xA/CyKHMrW+ADnaKk5
euWB75SmAIjn7cagHgS4zitUHmpmBD4hExibcdQTLabZZKeW3brh3/73Lqeu
nsImjSP6ejG6FrQH565pNxBIQhvqBaUsidPYr664j4NF3RHm2e999IZ/Ykpj
CB9TGRhfZr/Cjkg4EhmaaBod09GhnrMYSK5B8/XjflXAB0nk4AW2wYX58kzq
iwjWyAXg2OgH8Yku92D6yoX7ibF2XM7KEBWCQwekM5IEiDDT2Aj4NGKgbWFd
ve4PBos89o+eTvV9T7gpZ/Jew28bJghMaWfukVvPSwKgcFxepye1Ft2u6egz
9Dq1NhHfWuNyCMa3EcSrGIQQkwHaayaVPeCtj5Z9XB6qOXlLLV6/lP93E95O
8NyBdMtonkboe/k/hYRvupKjXRNghcBHCuySg2Z0BS7KqDJjvYJVljxFWD3c
CXmW7haopEDXh0kM3QuhnEdSJJ8hM/DE3d7my4uJnMidkVRIZQMryPdV/N88
qu/vGnb3BV9bHzWvsKK8BSfFSVx0tqyvCGfzMRxi6f/dENOvOtb4XHwPl5lY
y7jh4BXDiik6+xIjonMF4zOK/sUzqvYhQNw4fWTmsnMSUvMPjWc90YXbCgJ7
HVlWjTipB4ojBahkYNF6dw5L2iFmu897Ptw3FOUhZgsBo+A8IbTD+leUAjJm
5cMzIBOMavEKIw6ZqDx33xJA4VNR9QIUGH7s56u8hd4XUS57b+O+POizFkGH
9VNmw1LIdxvwFhqLRQ+fzPOiPTpZDNyKaIz+r4XfDvbV5NMMXHZIzlGhye2C
HYwwVyjQWDV/zOdvR9oWmhMQfPPLtW9M70cy+xhxkcnHw3cliuVyzqp7zf/c
d4chZieiNvycvsM3oJ214pewYFG6X6IppIdits8y3nZ8J6rBkFXGD/NyhQtH
uPDTiGY4OJwp4EPJHrjXapkW+EWeboO+buamz0mocpszrJXSGuNVIOTcpztO
SBlFduTTSRSUWx0LYw8bFDmVPboMrSAt1167gYQrYFjhLNLJxr216U1WNzuf
6WyMbTDssyn+R3iQwC+5UkzEd0efmDWwwXFxHxplDpz8qAn7G/RasZYqsAGg
LJOyRKfJiMG+CmehFnRhEbWsufTXeYaFxloMjl/o+d/WOTU2wDWa3xzh5u8G
WYJ9ZrsM6foHl6IjCxpND4uSBUIqnaZaYVKpmgpV5AVSaH2c5Ro1OG1GxgbT
dXZCO386CR+uKpGLkpPYKQPeR6KHmzqN1Q/QcPcfQ6Szs0nGDMwaZLqzygAm
QmK5tSrTMxVYL/T1+K8oRJWHaZDuqhZV382ZhrGJKzfWkSWyKukPtDemNrVW
8SX0mVVqx3GLNqx8dIsThJt0YjVZ9Ge2UZ/9g0Y0MouxNMCfaAqs8QqQx48v
57JrDs/nf4b9SiHMAMJAAYABtt57+v4KBsS3AtOwB058Giwc+5KUzE5rc5KG
0WQVyuS1Bcf50vDznEzEjBvARV5udAa8gKy4QrRYeJ/11ulyL9Bx9CNKJZtm
LDobjaOGmpQ/0MwbPFCwegxRnvbT/cIuLZxiIuIe+AdorMZ7t1uwrv+f0sRi
B/9tzUopEZYkwdeQmEn4/lfWfM/yHgjRCZXfUnJ3ltHWIT4R2l7nvTIrUFdL
ibXnz1AIG8VlIbBPWtEMm2Zm+MfBvZvnwQXm5rgiDj4Tovu7G0HCb+lKheX0
gP1Fbu3ftzHMspYzDVM/8to29ydQalz7CtznSsTvrQaHSj0yAZtgazPvi8fp
7S+c8WRHIpR8GSJpCvfrDMbsqOzGlJsPPVtiSA//nBJAFedvy8fWWRBzMXTy
f/DoDXzNDo+Bc8ed1jTTMYZU82Dy6wGnqdG0HplpwVD9s6V/ztaHhdxpF9UD
6ldlGQ/ASSoBhsRkdxoo8irjzVP93A/0uU09Fo01K5aQ3zTjRY5swcirwzXc
lnkABI144Y6ZPHk9U+qs24pumowsMtbf7EUFlrIVNXEK5ErrsgjExhLlH2yK
Z4kAkERQ0LIf0sbqfCl1unfpXJ0u+YuEpqHI/vUARYi5N06rvxjyvUacmwhi
ohU6xTvmOxllmD/a/gB5fOwx65WqkWAL5Blc9YxBWo5GPWDdhWxPOmG1YH6U
6FIn1kNJVX9pK6KrGW/h51QRW76xj9tpazW7Pi+KTJGpX3xgSQRh1ayCBlqe
UtsVVOBWEEeIQoGXJPeS4/lHqANjhcSgL4hrLWu/WH0jNsZP+J6VfrYY0FsM
fuAnWxo4HeJSaypPJyaLpDDYVVHC5p5K7VZy5QhV8nT93eySYXt+T/WI3Buj
SX99UWpk5xX3OkqPvWc3ChPJQTk2ZHfNDdg8uyIbJwVmTTGD/y5zcClEBGsy
/9XAEAOJOxFeLepEC22sgne/57W5JrZYF3RP9DnMB54hl0tp6kThaoq8zGZz
/lRMdq0g+k8WiK41nLXW/sEbelD3fnvWiChUw7kNfKzQhWiohPj/P+eL9d94
OaTr4F6SYv8HpfMcXoRUfufPJtdc2rPTY1Pu7iRtiMhtjD21rwrBerlncswx
sygcR7r4nDMHgtVKWuEey7b+gj7w6WZj4/rTWr6lCgSjzttS0uzkFQD5cFsZ
4vhqBQKqFO2aw5Se7H6dcQt/uyintgxslMenmX5euWvojXfe5hb0BnB53GSl
QzziB2IVOYGOVPYJO+P/aIlcR35XZ1/JoPUM1TdrhI93dLrnz5AhNOMh7TG/
6gdwTm1bDuM0E8aub6eX815An2FvD8AAvk7xmcM/dlJeNGrDxQKbsra4JDDx
ppVO0tH0aXQ5Hdn9kZ8o0zdkdaTY6bF+LsO3XLpIs6imb9haeQqW69SBdYAf
ti5/zzXZ2zVegu1qyJ/umut6srlXItqFZgVYTi1eRJIlzEZRwrm5eruHQN0d
dMrDcdahCCImB6h2PjOXqbfyO3jMMK/R+dUfrWvTADFnQuFOW/civws3P7md
JsCmdmm7lMAQDQf2RsGNbE1aqKH3MWsuyN6QTwiQAisVbJIz99X2nBPbBmsH
IojO2qLke5z8swjADaYeCs2gproIE6r7IB6p3ocAH85ttmAzMfF6/DY5Nrnw
XpbpJIyGxDOQenpup2z9pb2NUvojZ274BaWlnABraMoHM5RBZqfZbuF/52Za
hq1c3zxem/K6lhL0AoiViqWdecrad7VIem6yrgRPcJtwPkJKRtFtrx/gg2mp
TqgSPh/FKDM1VnjLpgma6oFqxNhy6P0yUOFTyeT1KPUPN4xmWBxVWBce2sOO
Nc6Vz22dsHIU0Btsf73+ipVTdIKkmoZVtE5HwVWy3OAaEfRTRXcCVLaC9aaR
zQktC4zrPS9P11AwSV69QeFYkYtjJR1AUbzRAR+4ZMmiPBkC4NstrkeU0ef9
1zHfrFVFPOgCyhVmT03Aa6Tnkg+QjrzUTt89/BG8uI8CauvKrmfbXKnl2nj8
U3bzp5udcr2L883KO+xTWGBFXj8X4x6zkmuKGdEYdXAcIO2X8qG7UR7Kdr1W
ebRSY7vk6O4CfjZPi1HWG4y7u8CIBrPhFgncWIKLRv3DbOwb+KmViKDfXum4
6i1cVbMwpPWBgGOCr99n8OiOVT7qPiQIXusQXM3BsJX/xLW1ED0u+VaJlOem
rLsvTVqBkQz4B5kePxbhhsQ9FfD3IdusdETiokTTB1avxumBzcnz5iLunoQt
n8GQa02Oa3mxgsOvZR52I5h7wYIRo9LFaP4OsxuUqwKIb/MQDSlgfvc0VKOy
5NLU97FAJbDxfn2NJTpCCErpm5A02YEzm7J1kSPKfwXF6gkewZJSzrqZ3yCP
zBcvi7MN9DgxjxKQIGX/l30TRI28z3ey/xCLm0cxOVrH+5hq6tiarbSUMG3p
2TStIjJ8hMKDt4OrKh7oBTdd7m0vyvpxR8EIByllgmHHvFfs52dDy5XOXAj/
pPhhq2cNvuronJw0mfHlFZ2V8XZYv2t0fIiTpjRmZ8pceQUpOHNZSsh2Sf2S
QjId2ffTbAdYBp/Fg/kSRUMcGYiCnjnyp4rEf930TBVE9DiDj+MAomRCRhpA
azJzoDpUWPQwNR/5nQ1yWG8jo/ZtG8o3pAaq9Zvvyrn1/v0yPWjA2g18XINW
FoSHqPIadKwjB3KPeacw+ST3AJXzbHXposESBbAFuiPcLuWF8GR+GT+M6elC
Z0I2QN9yTqeEg8vhOFU9NvKksNTxHGeIMBKNbCYUQlOHO7/9TzDHk9G/OPYK
HJcwWqjJJKJ5yTrh/5iFvU8NOqDUC1iimg4YSeL5W4VtYFWKZ2Igl+vFbKEK
f5dEaa5SPGC/dq5N3SL7/rKz7OPc1dilquZZ32+sijc9EkzcAC98wpuZh++R
aNBY+7t8CcP+2dVXtJ7AB1Jqoer3uI73GUh5XWD6LbuLbBO7EqW5i3iG2ora
ulqJnW5rtQztz+0m3T6/W8jq5OP8SgOAiBmklTLP+GCcFTEAqMnC4nfClArS
mAqXvJanZKCaKZ0AzoEMxAX0i7Cahn2+5JwcZVgGxcALsLj7GrM1iboynv9y
+wfDWAnS23YgiPsed7LvlYAIWZZAegWM1PLeB1MFuIGujf71826gSAFc6YJf
PdIIeC5DZti5DFum/KxEdmiVkVkoVqdh3uHsmGJSgwPFunpSwejGQVepzhHy
C+RmjniEny7WSUyzoliP9n/J0arCTz/7Ex7WvG+TDPtbR3czENRWhPwL7pnm
7i46DEAkMSD3uEV3gmXNx9Pu+wy5zoTHEnHWNEs2O/UV6pnaVoJRi8OLZ5Yi
Thj9tcPu5sjZ2/Fa4DHyCyJOr7rtqPh9GOdoWbfF/XzHJ0JWIg/GAzNngDbk
umSrDIYuffgT5KStlnru78jMSUiJmRgWw0uEupLsGS9Qv96gxfr7W8f5Aan6
fsYHCzDlOENIlpimH17nJ24SN6yKgxF6h2tuJYm3qRCQIICXtmImONqJKVpg
yyY0B+dJUGdCwrzqr3S1nmUxwrWgkCiO4o7acrNF+G4Mzto3OEWlHrEezDwV
e+H0gAjhSI3aQmPOxLtmLIghjdK5AJlmyKJL5OtKdvHuyfVmGCOApuq0YZZ4
2Eo51X4spGPVzG0dLM4mn0OyVXMEnCtQkpvZ9XiN73NK9PoVzhokmzDOTzqj
vIgcd1wa828lErai0LFJOlddrhoOz+W9DNFy/4o9cxk0lWhEVAAS48K3Vaa+
6bVyKnxnpT6VOFq9PJjskT/2X1fRFGinLkfRX2aZxo7l3scdeh/AeKY7wdIH
lJdKfqRs3uAfm64hYJy118w872mYwsQAPwyNtLxw+N8gS9G2ILqs3dYGcd0k
4GnQQvb8R3c4MVYTTUpKoSgXpeno/epf5esH68FQmuM7Bh+JJGW0czpQaDra
ySu3x4ICeZoEHF5M6S7w93IQPWiTkJoc/5IFWzV9u9BlCUbYlPZf+akfrq9V
PdkxAO0CW2e2yvpFpC0h86Ti6KRUSnzsFGaNkGO75CPzSW41nYeKuuoXo1Ep
sy3q0OIJo5SCRnzuaWNxnAx7rVWfdXYV6ViShFEB4QPKNuyBTgk6E8emOHde
D1oZjb9Kdz4db69Y6Nqs9Tbg8qeMu8l5lLP8xNZV2atmovQXHxkQMHDfjGLq
Ro9TZ/SfQW0doJGGsfidRbcyKP+xaeVeHBFtcWfhO2P1znklhOmJVVv5e98X
I3UQeEfLwNf3YwTmPTw6T0H2jheubHVHgMaLQROnJ0D3Y8RmNYrd5ZcvwbPM
3uhKBkUgvzuUj14f+KE2xNEm6KDUIi37hZe8qBaZhUGwOjXfThCGLFdjDFoe
UMELjVPuCTsV7hwkBn49Yvk1Ax5CdORDLVeHdxLTdYdDmhoSZrSbxTzYd0G8
sk/X2hV8EENOJr3YPmF9URBFrovxiBEqzRUWm9IXOEmboUGeeZkzsH7RXvzZ
pkwixxkhSAN0zlHOH49Oci8f+nbgqUdIBxJNd05yDU6S/s2HFGHnteiSlk+D
x7wHvUhRIiSZZDTtD2nU8TlddUSC2OteGDwOof11D4xW9jCdDHT5yW/4s89F
KTAGxDUqt5vmWZVtyw/cE0RC/1rilNcFQbi68IUrYLrYBntpRwYYMQJ+Hd2S
4H2K6+aMoFAsKW0ENL0kukJAxUjjtK3FrXo2wqDiZBFHSDa0KZRmZX80jpLH
7D/tLwPXCSU4qsDLrjThWgGq2aoceE4hVgEAJQuGZ4DeJyzBmVCYehPQhHK2
6je8jRuQw9DKh2auLBy9aWtll/D8B9E/SKeJOt5qBr6RUFKvYYTzENQo4+1K
jOkRUEy0CtDJN4cytBT4X0Q5xm5RBXrpmyG/3MQ4R9tkwxwJ2Kk3Q9Xf68Ld
NwiwKnc9LXtGrwCgCUUsJaAklib0keu/v3JEFNclNy7Q+/djWnHAPRqCOTTX
nQ7CuIDMIgc8F+dAEBhvw2EDYo6Vwb+lo/82hjIyBTDABuUFp7W1e/52Gx3y
ywgpHeYrOo5JaTGk2L4QkOhEIfBkFSZeUqhvgf8THc4ZDqrBeTuxRBKDu3rJ
t2p/S7hDZpSWjz7kFPo9WHVt4Z2DSYyFdy8KCkt9QXYCvKwQlkjcRc5oQRNT
QuDj4WnOozaDWamhBU0kYdIU6Ewr2mK1ze5yZR++Pw1E8fXyksCgbfmkX6o+
mpX1QYlKaLecFA9DCFf8rEXvimVmcnomGMuJHxzupZcQSoKWy1VJ87btrzQC
vjBFhjDJQXOKtjNeT5TNLVmHg32Ylow5GoYAG/4Xuqz2pwOov6iu/1G33SbX
emkmkm5vQlPiZ+vvyPzu0nOoBPz3W6FehCUIJwjxPCBO7TCC7yQSmIJRcZp3
+Qyk6weuRq+1qDiJvBF6lswNTG6CQLFLyscD/64WAio2kiNuWcAc3UDCfCA8
KMZake/MJRoijtCICK2/J3tWevCojTywPaqDEdUiKfvgwaW656MOmeB6kZlP
rgb5O7K+6qDqxAbMw8JZMlzA36IEv0s/Kq452wFM9hhQ8RDN/gxcZR7xZDy1
GrTsj6bAyywuJX5RiGwcJcToQ9CZBXvgX6lhwjwq+Bk3Uwb5x1RNUmuTEmWx
Emn85qAp2UsuzWwkuLyfr6Xs7vtL4YHOCno0LzwEPH8dqhO4+4ID4sverOZU
4dTwgiubwj1Dxl6jyDkMK8C11bvOu0epsbD4FFWKL9YoSrPuOPPsPgeLKFLZ
X5Zyjk+EFv4vozqEBcyFL5nylxhOetlZw0L+MQFZVuENIOLEvIxT9uYy2FeN
HD7M6hIgkpoUKN88g0ikYAevPUP2jLEEX2Mbp8q8pWW+yZsR3gkK703pIHlb
hnp8AR0bXMJJOCXGuWb1L6AOrXuUi5OzCfULQRs0VcohguMaT+P/vCqDTGD6
vxoOOvpfryOg6OsFUNBHc3vDpZ8pps6Ezc64zL/IB7B5CLLxm2DqeU0ziO+Q
uVR6U709lgU2xZgnWMJlw9IRNvB/T1ZfS/ACU0l/CQnxUl6EEGMUGud0M2K/
CLzp8FoVFaC2a/zPmLcef4yGulJX4gyOo2P/2m05DZ5vp4d3Y4MYuEeAPuva
xqKmu00IGI/Eq7mDlO2E3/bBQ6IAeQuOxZyLC2HrfMn1H8aVcL3OPVXB4Zhb
3h+ZNAWnrR8aVp814/mXoKHMB11xE5tj1pIu3FIwDjNpAEVkbup32vZHN+DI
OrS8HDX5cRPT87bps5uHbqMF5TNGarut6FxE8p5sj6M3+QSaZUwH/OeGXuwq
2e1LDwWkLrTHSXc3fi6MJG+NhkjsvryqrA0i/aNjxn5DCa4S/3H64Z3AM8IK
ie9nVYZAjmzB6vsULnfmty0jsKiXlbQSDhbpO4/rKOkqBRq4ttLFNPcmn0ij
MNhR9Jm091R4C4A1SE0YrxkQTWT9843/BFT1InF2CnvmvsDIb5jsKqo/HEW0
H/SMHnLaucFsQmcDEOqh70+wYw2Tt2G/m34AQ4qJLwNrHjawnpsrnOYoTfYU
+z3nN+U7SNCVczvJjYWhvXfmBddLhYK2YF04NtJ6zpHKrAI8alYvXeFEu07x
F3Bv25TuHxMWF6/7kArA4NDJEQIfL0V07IdYxUxL5auzCamX+azucFUYilNS
dLeCZ4Y/W2cf1VXGi1Qo3leJYCaHxblw80fraMYASgMcS4Et5BFknLcRuSOK
uob4fx7qXlw4mCvcz7bQPPfZm+Jy6kZeAFjjSbfEm8HA7N2R/fkZIjbpQZr9
SQce+7ul5/scxKpx6BCkFUtSwcS8PLWN4+0pSmmO0BJLL3e93pZZWjFNMScp
xdo8GV7ipZkDOcRtT38ebE+tz2l49Nwy08TWgj/na8FqTIE0b/fRNb/owSzC
ogZ+fh9H3rl+Y4dJGpz8Ejixm8/jrZkSO/dtbJqGoMht3IfG1FxJaIIsY0+/
y2HPz/4DtWEOQbjLjd2weYo3+QQBtX6wkcu0LREsUZpsKICEk4kl/bZSoK7T
I7E7t23FuODyfLOvOJzL6iZ8JlizyvZ+OEQQanG9TJo+13B+sX5S9VgnJ5vJ
DzglNl3CCI9MdEG1sYFDkbhImFZlOj4Qm4cQszkXKiOR4gU53r3egGSzUyJQ
3KKh8HxleEo0afSw1rmh9IKivpXGXPaa6N8c2C3dCB4SLxLKxBlAYzVYLmZw
FLmIapU+m9qEzrVPyOuKBH1VE7cOLnk1flcTKA9PC5ONgpeNDHB3QoY9OQxp
hBUDJcBvNW31gG954Kg6f9tAvhQhUH+Pmqv9tkp2whSBgvxj8/w3jnI3Nmf8
bYXD272kNfg1x/V4GDzoEzeJ7jsPCBT/5l/mSLJrhwqGR2mLjVJqMVgT6UDp
iPy9/3aRaKNbzRJByMmBL5ONJOhKAexBPtkW/gAvanSd2tc1hRoK9y2g361w
BVS4M6XBenBqpCh3dE0N6rKIayDtcHFtxoJvHeidhDBlZSw3I/nEs+GmR/Rf
x+Ke33at1SmL4lNicnAgcw+J/NxN26k2y+BVlEhjUbPjYthEb6jH+vgqsBfe
aKupnGGFDzkgHpxZwmbeuzKVFdxuUpKvG6pGlPJDXq4vcPusdEHpHCHhTw3v
1RPCDPjqafmDZ5lhPovlvmIBT6R7xAAMy+BzYcHzZ5llk7LyZj6ay70Hn4D+
rwlZM2V0oJF1Q3hz1Z3AMwvmyaP1mUFPG6Hz+ixhwc0u3KgmKPfr7obyNHMR
vzTiYX/27VfqiYpDQ5LQeGDBLwj02KKQLnhpnhD4A6jABAcOz8Ocgn8Y44gu
HhNszbSyRjcJ/+YL7etitMo405SIJ0d939mZ6eOVvTB6BUVJ/rM69Ks8VVLU
RlRcQIGlVcndyOX5+5ZY0e0sn9KZnIrORtlxUU0e/5fnkShNMhaC2kU4ni0S
rN5l5UWfVqRy+xiDO7ZSpVNCK4cwOs6go2WduTyIDXBqzy2HCfsMyNDVrtqZ
TBS/uSE9xh9+OZ1P4+rVKzm6LxKJsHR4fy61OWRFzoJ4t/2BwjeDVaQPrRVF
2h8tVo9g/rcJVCdROSYNvz6Gid2Z7Mo+yLOFsTkBUvcFav0brVohYkbBGhis
ntyjsdkQCTHkkzVbUxnYXgnxIjQbUf7qEBcz+TBPy4zAOicpLdJ9iuJBzfHj
ET8Kf3hd/yPElWp6hCLlZGctX/BdNhV73VOz1WzypF76UnpckuaIig/IaD9X
335jyzDeyPbKzS08SwuIn48yGAQCA8JylGPlfc5gw9blW7d4sBkkyHoRP0Gn
k+2wqxH7u8gkxsJNcSTg3lT0XdzzjPxyjsMcqEh6t1K4xbQvBzaBptc1CRkh
TlMS+iEPPRAoQbgzFifLz3lOMY/NRnVaVJYr0devVRx/2EOlDLNjHNFP5iE6
Gz2qRa9dPigE/uDxn1gPPqNu3GGIMEgbVauQbtkAgP+2pGB5m7ybiiB9Husn
oeXbiUVQkElDqo3PJJJ/JaanThZwQNl30Zo8rqXfqLSBMwDvhNRaMWP/Midt
d5dzpshePLDCEyQ5K5xXbU/pSooztGXDnkFg/lp6f2PrOWNAHfDGKI1V/2gv
wRSLdb12TpvxY6NVMfYudGy2jVQGFNOF8XLtANxwdpN7fiO666qbKUi44nBw
N1tMCHiA2f9crMSF5j4WFSE+vfuaGorkL+zmtJeMIDZYL0bxYzugTLFVE3dZ
DZV32qzb9dIAdccQXNtYETWKZYzZyuscQGEN6tMB78xxoqmjufTzzKfpMGcb
UQw7br6hTZgYIS/vW7hpkkoZMq3y5d/ECvIlUURcKEMaOK1cPnkuwQIkqFx+
/PJh6yVoyW2+Wq046VfvSbdX0eoFbv6EyTG9Dx4fvJfpLri57wDFAeU2Fwso
djjL3OGSMabsPFaqrDYG0/IPcnHpy1GGVtHOjLMrdVGcU31CFtFwODsBrQzI
3Hp9XMV+fq5H5cp0W594l/SX6XcVnmwBkfvq8RtdDgggLuEsn6HwGg7hbcb7
djPIOoniTjYrJ1+Zki8iIq3dCZiBeI8yrX8TUKFj95sFtNExgyFZ+iS86koF
GdvV6p6MT9srSpMa4g+pWx8pj9IOiJbCjdrVglU3eCpF4spsfKRpUi9Ie9Cv
hZLb8e/KiVdcgrrEticljXVYU3mS30MXMq5203AZZQjWzCwJ/yg2dJ2iJf5/
wzZeDQTApJ8FSuXP0f+bVZOMySqgb7CyppWMJCW2Aqw/2jwlDP6jxOsILUMS
DzpZ08OUMpLiuc8rkcl7MFXSkX2mU1FWpy+y3eYYpSO5Ff4t/KC77S7gIK5m
Ub32y01ayjKFtMa7zZxIaWO5W5Jth2Kqmt+9IIM/153tAg9PT/j2aydCPZ3H
WIuUX6nc/Ls0im/u7v5ib9Ava1lfLV2NTctl1cV9ejxc/U28bM/ip2w9KZZt
g6b9bsKO2STeMaUlvHhyUzkFa6k/RhmW1FSEzz/2oQ0mGjXxgew8PipMK1L8
Dcxy4tJZhXw0A+dw8luIuP2P6FUa8m8iBelBRQBoLCr+YghT+5PJnzxTuNdV
hStNwXNa1qNF3+SyMxu2QbAjYj6FnkMpQb7414YCdGcA/+Juqjm6X0yKFnNZ
0x7zhAIdtMQuYCo2SFbcLRCouHEkFB4mvQAn0rrVyiVTAORkwquIHsANHKL3
+Y4ivLCh+aIXX0ghj2tEOwl5FWLbLDvubJ2K48wPWXFNE9tFG27s8xqrMpdX
qAEbkl8IUnJo6yyX0W9JV2ln3bIdHl8tO05ltLBCKWCUdneXtTqhBcJlUmaE
7MNyvJZ+LW29p1yocrKLn5Y6a5ntNHoUXl8oH1Z9kZayxos+ff8eEkkUjdQO
3gti44Q2Gl3FpPp1J0s+DQdNuMd4qhTgahkxx4dyOhd2sUPFooYbpl7JWWvq
HtO+IIlhkQks27j1qIUCdZY9QeVz9b9ZE+edaPqmZwkWSCBJognpXn1gn/I1
wqnz6G8ou2KLl7l6givlOAfqwEHZjW+zVsyEqd3e3Rk2bsKLxyg5pLMTFI4L
jpd6iTyBBEJZKnZt4TA9gjMH2jOr++8ec0dNlfBMzjESO3MmQluP2MZkhWlV
wOMkAwa351QTOd/NAL4g99KBLpcinoG/SmMiwlnC7HP3ywmY/e72d0omZFiq
+XQG67ZJmnu+8ooOldwiGJZiuo1hSh2WCnj6PEFP6Feyt6K77KGHTcFwqBwq
YyrtOjQbPP5nVjlrHM8asEZ5Me3vSSBpgmB5vXFnIOFfhQwvDWZ9HAiKugJH
7hoVtib+LkFTKTLFaAnfu0jj3dNXE/W0H2pR++v/mmkc/FcmWN6fyg5Dyl33
aFvbHM1ccKCGsz6CCI45C/Esl18Z8JUGiHqHJ37toNFblo50dByEo7jw197J
cPhfvYXSfZXAZJ+FPlB8b/kK8jmcMW5zyfvLlsehltHh7gEnpvA8tzesQBgr
O4yMVvNLpspdm7r8J23hZSGLeh3yfS2i762aiI11qeMW8xo5t1wcFAtFTTLY
eoEbYoIVWmDZeVh5A3pSvFDpEi/Tk0me2hbEN25w/uQAuBqw6VZcqnJYeTqY
EDx9o+DYySaITKfj0lxMzOdBdmVooByyBJub0SXLgoyDKY564s4DZpj3a30O
i6ObiqlIGc+qzlGRKViMh13H5rZOsZmTFENJW4tc2bR0HCl1ZF7XFkboQ7/z
5zEulePAb3gHtB08YLWoFvSxhk4AKSBzojm1keSv035VclOoh33fEThyVZ2z
boaWzFp287CKeCiRflTK8+IvW6bWVZVUICM57UFdeZKPeGHVUGvaKP8zYvzE
2G6VIVbrSFCZDee1YkaIXH2otj25ol60IzI65wPFdlLKvTk97TzW58wJBtJZ
dY+HhoUMtR4VZ/TyWPbGz7q2AvrZ9ZcdoUigT8aBaMddNUpW+SaXFFocLctM
hQKiPOduB1JV244KCFsE2jObGmT9IWwbHoVG4uMrxWv3nt6uBwNldi1ADJoc
Pp4dEdcAETXCnOMiMcb4/ThE224DCYSAJBRDJnbSEDn/C2VfqbPDKedG+mg/
j+EJ93ULVY1JWzVqP91iIXrdIvZ3Hbz9hWWQ4X75Ckq14zIciPblZLhLz17k
kjJQtlcRMigMcXSO2hkZiiLLeIdBqOWV2YB5yj6tzggLj5YwKODY6SlcILJe
Gdfe4EEfpD8lj/eS6RwHWASSFkpQhbt/9ZaRKJ72TMPecwIXjzt+1Bl6fk/e
NSjS4GdO1iMRFA2PCJerCG2M+jtKXpf1Ee46/epNkvrh9oMR2zfw+jFRzoRH
uCcQIZSNwBGQSc9qEOGdZ6K0GCdjTYbd941SoEfv+kl87HTdtH6L9p6iFMDb
epX+genHmxsqLLRSzSdgXs70DTduTYyhFi/AeaXMDK5gim5k0gYQsrJPffqQ
eJ98shFuKT6ACD4UD5YQyCcycA8dWrETO2b1+OZKTn/MOgDQdSgqa5swWChU
GFUtu/nV7GQXvpEMmhbEwNUUBQ4lGdG2jAt1hDjmfX6EXNrpe73h0K+SGALe
SHd8lkr4vQAPti6ZVilXDQj7kBeoUREn0fXT8fy4MehkQ/fiaXIuczOZW+ch
tdiJ/qZtVA3pT9dMrzD/3acgKuAu1GM4qLF3rkZtB0eVnvf15oOjkff13naS
AaODKE91SVQpEooC45qhujjkTLbNuZdJaA8xPJMjrX3vduxlT0YGFRK0OM9V
ipGr6zQkKK7w4+5s6F1MyIwqjOr+BsJNXskfO1wk+xDcc+MarTAUPcFCxabV
MGRKKlr+5DyZS0nFCFpBJEsX5uebh/vP4oYr/Z6muMdUizX9PBFj3bqYIrz3
F+u9AQZjGr90k1tknFVIPHJgFRMbLOcvmIi+mGVIj0sC1d6iDiDYM8WAQ4Xe
b6qK1+sIKJAbssf3iWbdQa06j2iiagvfDzcKOptLJGN9vRCsUewzH2+yotE+
i2VSROFj8jpcExS1zwJi7cjbcgp/7M/Fxs+wNijhnyuXzIkUhzDnoA+1eIMp
o+oTMIDGweA5dEbPh/ycl4dG8MVWN2ilJNzDsKnMWFKeXmzRNX5d4fzs0QhM
ZN9xfcTHH3L+a1r29ea9FTOKh0yOsWQltNLzd4uShKzO1SCfDrJfWg9oba6R
mLcXPmsBxnGXqf1jSsysW4NjBIq/X3PzMqgUdlg/1YkPpYH4AnPeA9eJJF78
FLo6S9gHr/FbdrG4PPiurR9TmX908lzIYrkm7jNVMllsKIS2SUUVJdXZLqoE
kEEkxyrD0z0ai/b5DxCsmCF7KhIpF00oOEFva5JlwU2mZTMVAZtFmnJN+hf1
YWuNJQUOPUD32Gme223QKao+cK+hN+Df4MU90wNwd9y2S0XBIYrDZetHuXq3
oUm6juQ197OvzJ8JbXunePGQEMHzz+Bao4Ro9Qkavtkz7NzysylGAsmXunLv
v0kq/BfqSRp91XPd6XNnUcERQS+WomNqxx24IAA4cFKKVfUT83NTnh+nEqqa
l8ied5rZtcqoLmBuX2Ej1rioTxsO6P1Ye6VW4jzrrXefDQ5HTR9WHrZpKplF
yQyyyWJGhFKGB3bpf1AXQPpkxgBuMZXGJQ063kWUH2veOELG/tVEGZXhQ9P1
KQneGqL7V6JFyFOcC4h1cXf/X5ojRAE2AB81aguqFxs1f3JXTmjCdqpkdPdn
/d73QISK0OKDMMubGct+j8RGsMJZDXVtSnd7vu6BTQy4qT0RiJb3TnM00HVz
WzLV3jekfokK64ZFX1iN3pMzxDtx2xpCrLXPP6Yny8iVPtEfVylEwzRAzIb4
DwjAI/YQjtMzAWMCbwpo2SG7H6YL6txml9de2eZTQDPQiwOueiiL6wN6zIty
MnIJ2MbTfFNy2VnshYGAH/XguLF27mHs5DQki29AHV5ZJtNrCFU2bt7LWUKS
NSO8BCde+s9/uWdAsUGgiFxs8qiyCtMGPo5tBQNPkgoIRYkoD9RB3gF0Lalv
AGAfzQJwDTVRarmX1fxAVntC65BQTwqLPE3P2lpl05mBpLx41vyMEfpM3++a
KB0IyXYwdOtmmwxBTxIAyJLXwtOkeNGM0QcjMw6ThixHV89bI4WpX+G2F0Tp
nNTelqGougIG2XCildOb7foGnXKyAF9Aowayclv345l0KKP5PN0KtDOkNxpe
ssricWMLke7p7N/XLyphvknc45LrtYIrp+Xk628Vk46/S00YVKYJJ14/o2du
zbTj6jtIqH74SsJVuX8ToncwySLoKsd7GFwGRPjPwdqjFjVjhcO5/5/9z9W5
0E7VOGL+fAYllBIDZxhQMRenWDOHvj96XjEyStCIsjcJmqfxi2Ge8dcYDpRK
FTEMOZoYrKqdqi90nUyUqrzvkCP0xJf8gWqBUkOoKY2+iq71gR/7/zx99PMA
jygWHk7Ica5XpFBzehlL7rIQ2qDC0TjeQszrz6vIEsvgU9j9tv9drmqyoNZ0
CdkLkqwcw0IOPApsHIf3u/inLsfYbNThWQ2Oa98RmDWybU6ApLSQTQuM3ynD
+zFREkWm1fsce6XKLYT3LDESc/egz0UOpDKs5SZJJftudv2lQCbGl3SnouQj
Jn2nWjeENOcbl+XdBhFps62mX1LErlTr4TsRMhVlC52GxfECcLyOrtujCt2y
XmoX9bLaLvuo+3YJE0NTXwJ1Dc/1ZctjxFm7MsrEm0hap/qztGtdkXH4ANfZ
VOJ4T9iwBeKIF4Iq0HNDTypELLbFBV5H9ay7DXre3u4FLQxEX/qyxj2jml3G
fYZAMPHDilYZvFASS00c4LIJXQB7hnGPcMxhc6f/ZE+Bal1Z6D47oqAawSK4
2BQkAybwbi3ZrGSaAc9up09I+oXF+4bFYif/Rk3JSjDvwCSHP0CmpbfXWlxZ
ddz6y4Ac/ANRB4KPKSci8zDY4nfO2MuwCRr25g86+tMzWhd3IQT1RW6T1ljy
/iv+ZaIDl5XsDcPAHJm07sHHNIW8FojRCbyccnflWEbVYc2WOQvVaTR76YaR
aOHB9P4LXht8uz0ABTO3utunkFwsqXvnX7SP9W0M+oH6GrL/h7DAW7mP3Yvr
o8NxyHTGVwRHepyhrol+D8q1wU4z8UZG+6w/aqI950e8TuX/Cn8Bj8Zc7ZOK
ThrguPdH7gfetwR3UF9vLfmpC4iCkaBJl7BkcLtbc1q9TdSTRwLQoX8A9U04
akUhf3c4cK6kbe10dXRIiyLNUENqJFBzSEDqCw/Vh3MmofPZoypCZkgbir9k
3DNCpLuydzkCkNvN6apKYY9Ld813J7/1qN0c/ohLhdcOdd3vB6XyEbCg8RHc
iKjoDlr5ha0kK5swiTrkpo+FfnqKVxeQyS56BIRKT6VaVARnVTSxLdAC+Lg2
BvQ5zpYGARlqId8alf4AMrxJVRprH54p2OW5qfI3Oq3sC1fKSsVhb9Fz/ZU8
JDzyl7aselWVr3JhZrspH2/ElMroqWsR0rT/Zc0EDKgfZIbBrq2JgPfr918i
eOfbS/JIt1EmrC7U8AMDFsJ3wtasCyA81JiENFTog9Iv61G3D8QaKDru9q1v
hlg0HC31iUzsyMSPtyvYBENITTISPm4JOKl4j1XDGEmJdTmWDAGywWiuPRLb
2t9uww9ebhSQUD/u4U1WFEejUrjVcCFiolfJm6s1tyQMcUrO6Bqwp2r+DCT9
4WnefcmsIvvW96UV7Y8hOdsFHuBHEOjEHC+MuGDq1h5SkWsJNXEqugD4jxQh
dfKLm55KvcBWbO5H21mJEchu3AKhVKithBoZLQp0GIKz23ZsuzpDJwSIIs8T
GVYydjC6wvQjgdCNVRx3+A5F1bgNiRKfwG2CCK3oOj7RVpMiuOoKwYFCoUmY
C2E9zKeHhpg6olj9eSJTKYKnKTyr1PcdjDu8t0MAKSdxaX9My4brM8OVeB+4
zsID+rNMF5Ad2kpqYX4L6HO8t9zrnsbjPsPTPWWFtRm3tIEYPYj99F47o6tK
nGpzrkVMoImOaiyS/B5vvdeJ5RUozHv/7pfN1Hx54WV98Q7BWRA6A4wSZURI
W96manvUc1c0TZxLL+d2Z7PTCezckNllFlX6/J12D8MPJ61nwhZISMfnrM9X
SZgrdylJ/LUG0Bdb45Dlena/1lRCwKJzoWrHveC+nDIZHAoNfEQkcCXKEQz0
hpI4ZdDosBOQ1+rzujXBxV4HaeyoJ+/RLlUJNCQtlT8VrQ88pZMOby/4zBx9
YH8xomo9ln+grvTSGmV3kESb9SLA8rOSovSlMF1fqdV+Yd03SntDCPxpyuTf
jo/DY2/d8xqMik2vDn+1RU5S+eW7QVF78vcy+nzrXX07MQAhPKmp+zrNCJz7
+4bRNeaZEpRVhGaz7V4Ge2H5ZHnLBDiDMys7V72RSJ22cLGLtuejGgXe2rz7
bPafXaVPeKF2+geERWUPRzDLVrwia9YHIKnmRZu1aZaHe6GG8mdgIH7CU0mD
Ro3+d+jlyRc6kOCyl3i3UzMjaMmdE1Ek7I1gyUaxNSZ7fbAQFcYOITxVBx0r
qNa+6ZPPbo9fr8fKfKcenwdn3Lk+YkrfJD3HdRxGGtm5IHj9OL2PWSjtubT/
G0JOfyqKEcbKnGK77jdFgsJAK6YvtRjOXhbtHC3EDmNPhWt7fvzqW2NO5229
FxIgU/KtnVqZzIEwt/a4HDO4MUJbF5P5JKDcNdtjoIgPGyXei3Ryd8MsOiIJ
ijILkP0cUQwipXxoajRAK++Eyjj+F0xah3y9aHHr9NlfY8BxlYdI1zbNE1Vb
z7XQWmVWZbrlhZCVpsv8rNThr7+2Fep4wuVmBIct0tXf1ikzga+7WyGocB4I
jQxeTVqiZWvkR4iCBBZirJJOVsio+T/Ws0OEMDVps71I7SH+ykR227dt40Ly
Cm+cLQJQ1i7GZBl9ZCj5msXWwDM0n0+O1Ys7OWzsO6tus4h0L41rxkhLtDwi
EMzOr3bjeOrMhYfeWnv4+I010KbJXHlMp1zm3MwigLkjcRVUA4TKfY+zVGUK
hIRXXccRbz6Z+08Ngd0C3kPHt+Cw66Yh+aerNGFqdRlLTPMvqMZwbfdNkhig
73d1FG7G4yL+ZWu44qyvqyztNTKdFNU81JRZ9YSBIUqCnQkJQUJrnw40I+ga
8zz1dfqdeaNNgZxXMjeKDXo+fq+xG+M9KxY//ZsfHwEj/zjD7et+NVhTBnIV
8cJE15OXpQZWQxu5BVmNK5r94oSbYVcKg6rsOPkP1/kS5G5IhI2ErGBaVM1g
/MNopnQmG5EQl6niVLjpf7LuuDMUCiyEk6qbF9CUZTOlfGY+7Yjrz4Tzl0rJ
PmlaXZgSxs9CXg+O/INk6e6uVBKO9Rjjaxs29kjWde9gyFRgaoNSx6SN5TJ+
eidJCYMUCQ+GUEjlBerAGOwFpkQuabKEZVNsYZs6hB+dCF0jOr27Wj1s0cXl
pRWcG4jxWEsfew1A206N0wpSusnLJOZVryH1/ECWPMRF92avU9sAagYa7RGh
N3MLIsLAJ7DlzLeXVhzmugFpUt5Ba+icOuhsePf3+uzR8GVrtxtFhaoIDwXb
UvXfb0sYTvh7UEWrAPlp8l34i6tuFdwP2mxXc4kQAgE7BkEsKAOAeo7q0JS5
D4JBORdsFtrxMiNuOcwSULmdyuAeNuYsmrlzL4BgKQTmb8nJ5d5WDI0SIbQr
LLvgXAZchnFIXYXxWBQ2wf09dpyUqhvuI2n6ttmiSYNhGQWqpPZxFxx1AUli
YIkK3PFd+KjlQ4rX11troaKZjbWnkzXVdS5I9zPqJeGvT4tThQ/f18msjfs6
op1DL9mhlvNHmV1S3VBHd5BXQBp4gmwYNeN0oNHfhIzVMOEcCk3+v5sAiBEY
W31UJ0V90jhmWv4hL0Plow6Ax80fhBEueOXOuhX83VW7HlgrhKIpLh5/OQYl
EE+5YtRK7FY9HI9VU+72x5Ps5epyUZJ4L684w5DbtlUyB/48MPkvE8iQDHya
9q39JBwx9X4nJpAHAOlBWln6ScZdyilxp2xxNSSGme3nvjZL2HdRuV9vlpDS
u2FyHehayF+khwF06gu9ccRd1R8yunA0zk+eCtPD5E7Wl54UyTDs4VSP/Pua
GheVC5QQMArplKykimXv1wIAReib9bfrhm7cU9kC59jC4IRC6IqWdYOgWowq
m1CmigG6N1diaQdXsIZ4X0r4APSUeJSLsbf+kxrzRvowTKC+Tt154lBcAajF
ry5ok6tx2sOK3tk1AfPwkSSy7g2IonKN+DmUqO1T9AIasr3AQh6RaQwEc7JD
9dvYqCiqDqnW5out8Zmdp06Lsn5tOekpmDFkmZ5XunqBG+lqPsYawbjCIFtr
GaGtTD/LaeTZevNEkH9ywKxZFK3EyYcv010pMvu4jB5lZxrdZIlLgj8if59X
QxIOMaQdyfktmlQP34UbVJOkfIVXK1httqjFwiEVvHK8ruCO9ArdQTWKbqha
DMKtlUQKJf/hjQqX2bxPK7EjNd9rjy5GXMEFUraZ1upTgnmaSeAxNYarXZtJ
BF1dN6rZQe/nIZdm3D4pdJPTzMownUxdEBABvVKQ0TC+qbOlkUdMWBs+Syb1
QleY9NagHEO1VHAIcUb3cvTtH7Zz+iayV3LjVFU/XWXD87ikOGKzVCbvIqfm
evBb5hUPDIZYJxHerxx2Nok+fmk7WQx1CzKdTQ0DqF9k+YssjYrrjs8jjo3M
btHMJLy8mus3TurZjDk7Awn7b1Fo6mlnkWvMxXgD+10uNK0kQl9XpVV0A5f7
lh9JE7AlqacSoExOHie6/OZfDNQDEHviodSlmR/6YBDeM419YwdoEfu8SfMd
6OGaNyCsFZU1FQjHN/7iIr+xjhrrTXl8CSyE5fmAnkg6CW/aclZaULplRFgG
VZejTND06kZnH0L+8NHUeMCzQ/NMeOC1ALdQ1nYDKh2GIrBaXvPDQSLN+Zk4
5uNCJ/6zewH8j00FhS+lZZUhXxHFs6b4w+HLWt7K62SRL4dqePobDlun33Zl
xdp19kxy+SqO4lwbTYMBlBRv6raWGmLz1Q9Ll7G1hwFm1LrXesrcW8kSjPNC
m4GlAyftIjI0p32VEw4KBstG38MtYUc0CdRSteJ3gJbiYh43eHTZvI+Mwnn9
3EniR67ngpedC42flmNgvLrwtEgqZ/Yw7JWGtikcxmr6iq8BF60qfW0rJC2E
KTSD59+QnvrbVof7MPEdtvipD+8zqJeBUStd8+K+LChwoJikA8NWi1ywEP85
LPizFD4ZZ3AORsszm3ykPEEY2IU5wQJ61cLzLVUmglo7kC4Y+t0nkhlgZM8X
gCIu7z+v82eQvcpThhXFthLmTSQ1nVJGKi7QFQ0UCVX+WQWTOWyMW6OO8wmv
qZOPFZRqv6VFvvxqn/Smquv61XXUxv7jGtK/ZsDE0cwD3rwaifbLg54TsnbA
ueta7KrK1dClCTbtxsJVP4pgETHaHq0slKQ8mEpC3vOIWOnansux97IyIX+y
lc1hGZZCEU7G3pjzZzfdGHZ360bSsWRTUHObkyO/jHYA8R+b/78YQR7RSin3
MJHlc+k0BGXS7ShBAzxsKUzxVuzVSTO5RGVm7jAPsNk+SUqkpZfjYNlCH8v1
+1gRqunMsfFdjVn9belVvFTWb9qVb5/RDMOxMlKN/xZL1c6cDHB2LTcpOUPu
4Db8TVirXmqH24dDQhHO7nROb7G0FDspnlrolxWzcDN1WoCEbXWa3WLQoJo4
I7tmBswGH5/nvBQVJRnYz5O8fdPbUPQcpGzfoa6BYLDPNl7M7OKZv4brw5B9
8/P+aqPjiWZRv3VOxKpcx6pjcKbFl04XX3VYLqgxZdsUxB5/qaOolfIgwwvs
oGNY3cLESyLYIAsH8Ed3p5S6QfKVZwT0cjQLKgC9owKj8Hu5F6DdSHtUIMcb
zxHP0ZUHQv7vYGKLJdKUsR4vGZIICPBfh+DepHAJpmHOfryr7PWpOvlmB3j1
YrjGkCaPX+IrbBneswSB2EHDceBx04kLwX7QOhVabYPQc4bxcBkxghAlka5g
81yVbdcMBsjS6VXJSuo5AdfL2tzLzj76ZNuvHD8Wt5Md+1V7nTszgSHwmw0f
VunPg3CTvzKQa0zLFCTIVA4MfF9pTBaxGBt27WyRYoOfF5MpBVlsjBduQgea
iyB5MUjaix7WfxEZWYc0o8r3bthhcTWzJ9bIhPJGlL9d+TzgdvlAprVHVAmp
+ywKXLWUf26rpI2hLDUSusIeQ1AtACH913r9eO49oTKNQjiu1DfZX3HRjEQT
Gai3eHqCk5yuy4QWHG6PkvS0nc13IOK1+OK0qGbo23rvWcHPuJi/NnGomLbD
vk3YsD1LAkm4QtKD7V10ptiXHxIBHeY5a/j6WVK5yoIVAFgRIeoeSUlWS5cy
MYV3Tr3JzGbC4RaCJdi6BAbIDLiMamPcfrO9xRdtnAWc225BtEkLqqexZxeO
HGTyBBUnj9gCDeCVf4DnovIDBtjk7Y+EccRJAO1MXgPP5/eEJ3q1N71tXEJh
gFibF9jEQn+DQNYfiCff+weo3aqjQiX1Ijf88OvRu+Mx6yS8tE4Rx/Z/hNnV
ADPegQ4Xvo7NNFF4+xXELZAUcuh8TfkuWFoW9x/5Pj01V5BOcUL9dRDdAPhZ
LPS0EpIrtz7t7ghDTDOC5RvZ+tK3lh/NI4JAES1lMjex8gfwfzIn/zPfjfYg
hdiXCzpNXfg8Fzl7wMsl/JKFGzB0XYUqeTVWtruvRJ1A4bEOiHXfUSnpuKAP
HEwP0kxfYvm7dVNCxg3cOq31qdReudAe8uZWVxHzXH4imET+/MQnjjb5dfFk
/0qX7xeuGPvSNKigwqROyV8vLuYXiIjFHwdYORlDEjlS5Eesag5cfPgfO/vT
01ztkocbpx+hKOLbiXJwxvNaIfxlJOzFj741mY5Wgp4O62re0wQiAtz/PxC9
oVqvXZOU+Axkevws9nmds71hjdwankebmiXG1xra1elgNNrt0aYXK1/r14nu
PHrIbpe9h6rfkiaQWaB7GssMAQyC+gy970AbrHC4UBttgYAuWQnXbCenryEF
poyuwx/ddGKDLgU8xNXwvj8zm4LDjD/Ojgb07xuIP2+egqVwmeV+rxt5nOAX
ourR3NxlO8AGb82oFER42dBXWkGI3xBKYHk5HfWwG4OTNVJwUry00kWtMT3J
/tv5pUJOR8w4GsvcfIHZAQi1UIlcIRV2a7u8BtApME4V10pBzn/22ZnxZ6Fa
oVbcsuIApBTT4MWlVlNjvLw1FX1Unlw6o1xEDpVEKGquzD5bK3ZvbEGaZfgx
KHUaMwyX17BkA7NwDBKC60o7D5QXkv20Fm9erSns15yaTpA9WExKRvTtlKyX
gVd928cOkGiUoxUFjC71zVEEEi7Ee2vG7+LUQ0v+uUTVOoRK73eWU01DojBr
/715xEQneiaJ/jEzOENIQAKXuRwy2w1CtHv10DYAQTU6tElz6TMwYWliycQU
lP/e8eNAmz7yZ2kNVqhkW4i1cOToZpYHhJcq3v6IJVPCvcC9KUJkY9/w1A0i
q3maSLryVdFhBdQbN/RuAFbLlHvolU6v7kErraXIHX29nGQayIG1bP4thHP6
cai1gLcQGk76fdCV2478KAovfxMso8qD0wFVWW364NYy5mS3EroeIUxSLIqI
1isW19piA1bB7GGRHKY1Xbgwz+AuXjgYD/c8ZQ8JIAYC5haw5OXibuZLkMYJ
w8CeqvRrOL75cjhXAIgxWKiRV3OmSPurgib4prRKh0vnn1UfqoW9B+/OLWAr
QDZfoyqEaACwA1B3iCOpgIcKzc3+am0/XDiWCeFT5YgR8HIMEF/krns9wFSR
P0CnUmcYp9SX3SKWzBLOrdS28ejyLjAqBerqAAkCdkJZGLFjKEExlmZEiXSj
zG5trC03RZ90yS0Ka0OlH2gyU2VSgQpb/EmYRqKhXNHllDo6RnhX/gzdZ+fZ
wRPx4Tsz+SEPFeLHJGLeT/RwzXdB+Yp90/5LMD4sgnDxpE4woBSFCb08O85E
IvS2Uqij1sF1upGIaumjNL4Be7VJPqJXomZOamNZbUGf4j25T9s1B/xqSaaO
Hlts3BoQPz65Zn4hPwIVScqGqGxCV/gIehKPlw6RhGDixPyof/W5mRGoQFH3
MO+zyjM29XZkrOHYSaFaZGwt8xHzLfZSip1JwPn5Nhz3hPdM23lVCnWdKklg
7/BHqgfvixOyLfOKUKZuVAhUTuN9wOaTHT09ZGdHnSa9XU1p7/LDUYcgi6En
+Am0AHtairOnsvydvIK3lBgAd/sWaw4g3zHQWiF+kt3HHGppGoRb4o6BIxXl
oBrORZnmJcWRBS6Sq6nxbpFiAghVSGqRcctS+jKaiouIN0EcrI+7ZJ56TiTq
+bYv6nL5OhzSmoBW7nsuifQMIMDtrPbErAZSnyZQ6AELq/MD0VmNAdWzNLil
QKVh8QPLIT9XZ3LndFQhTh53yVW2r7RdNnCvB/orbBk8rS3wmx+LfqF6mU11
j86x25TcKSG1ySuUfz4mAW1rDIk9IC/No24tKZDHZ3X+krB1Xjc1ggxZvfE0
ixRCI3OO1jZXw1a6CQ/1IbuGwCJ7Z7h4C4H6zIbh3QVmmiSfOx59iBcfkEHw
Iqt8uZ3yHdw5dWekL/2dDkW+aYRKgbVckrDYFNjTIPu9r6LRfs4DRDWvJYa1
mRSRbmQ+eCyqGu9BJA0/B6bbIfNCAeZCs+q/y826LEmO//UrH2G2qMvOPO0g
I3OVHMyPiCZZjhp7YcaDf8FpjOGsTaV8/j0bo9ZTqVSHjctZZSkfWNnTHBDk
EWo+PTMuYx5WQ9/mucvCafDABTvZ9KnHotKeWofogjRMZLILMd+oa0gMQez8
HpY2VN7X9P+2giy9SLw8SCx4LM3hjTZqA9MtgFrm7EpazxHRkWIZ3IKuDxR5
dqTDd3omHQJMbJgghnmtcXVhMhivY997OCQGnOTorj2ZhlIy16cM3oRPFO+5
OJFcMq89SNHCHn/vfAiiOKAJCejZe6ceTuri9mkphpRZGqzwXYhURk7VhbqI
TIcoR9yw4/IpMi//RqC2I4MahqUPh/X5cw58mjDErjCqw6ZsIy3Vbi/IK/fY
p6vxIFKpM/12hP9CW8sgsACnbMhnq0+mN0UCCmaQWjvlkWDFBYdLYeHvP+tG
HMvj41me+MAp6zBpptRHs7qCem3GGgiQ1DI3DyLpRQ/v5YsE+J6pw91+OeGU
YB8PZ/D3MgcnFjfXUxz7Xnd6CjaW+kXItuy8QgCOhVDDAyOqJYwlEI7mGJIA
hiAn0Q33PnGvHo4DqTmlxZJeZvNu4Dk4BdCCQgPhhoqsagayQI5Nxoe/sphN
tPde88DinyqndJQVUokYee9NDJsVjw4UaOfigvQkP8GQSyV9UaKDPdv7Nq9G
39PS9ujrUyWDJF/QzGY12z5wEUb7zes7GfR+T2YavRI8r4TfUAHWdtYXyR/Z
29xZzt7gTkL/EopFs1QLde3fqMBZ1Ve/74+vAdW9++wn8kz3ANtTGYSkIMJC
N02KTrd+HIBHjtjh27C3VPHL53FFnfFr5Sx9VtRkYciER+s37X50ZLS+y/Tu
SiHbIA1iZpOe7tlvHUR+fY2dLRifLStdixyI0YLmJcluazLpyMDb1hiWsz5m
s+fnyPVqty8Qx5gI2BeZb4k8FqEfo6VRiyhNeeZjR8wLQAMEoyce9+GDa82R
lSV19NqiVlRTjn93PQqOB1YAE/xUvs9obDKTHONVjLpXpLVNiaDXZVAnEzbA
GQyE5OxuhsOnQNcyfp6v14nmguEXKpYshtMYMf2ajHH5iO3tm+HeAkzRGsL7
rlXjNT2GHM+JRudlMRb+si8X+GVyVGnX1TyVDsdXIpc2i2DW0gqjIWZm0B4B
puKKjpYwT7bgEBowNn9v1jqBiYVtnbOdbcJVDdJqBa2V9ocq5hYT23oWeBSo
+Ge5W3miH3NaLgv9+xNd3Up3Y5dv5cIM2P3hNcQq9mS3voibAclFzENg3D7G
nKO1oO712xo8j9cWUKSmnLfY5tQySwgbeERQyerj48aohMhikCOF5rCoFP3b
++JG6OwgAf1C2YW+QUZhR6EbsKSnIMIcaxV8gQzMMn4cJdFF4UZAIjt8QWz2
KOrHlbKdq5I7OInnPf8zvwFij7e2K0+yjBeIgkaWD8+vnf5QDkKkruY3CjQz
6SakRFBatkFGgmYYomZSbQeRdtyOEo+qYTAatznR2zJC1OU0O6KMQGkRDZ36
ZQj8jV/FxDqqZn+0dmO+5pEy9/TGb2GfLL2LMwKAfHPJiWe/Wz8AWQ/x3+1L
Z3gCD++O5j7W2J3h38y3CxT7AKG+FhuvaJ/3YsY3mCHLJ741Mb3Snx6dwA9d
k/XaPEIL+9dP5SDkN+CrwuJuJK4Bs1VHByQX/wqBQy4zaXXOpvtwseqaEnFa
5rh3DOwDm3ZcVq6agIuRG8pPV+oRlUycySoJOJ6wljjprBKYOl0UckfHpLRc
i0BeihddNYnRkOsxhyr9DLeT+mLzebE9PVupjgM2Zt1eK8cINyOdwLVHA9DN
LvpxkkYs8BLhKf74nW4ntoDBlxkHT1t6miix6Ympkl1lIijOQmvXrYw1Y/gM
W1Hq+zJmb80yq5ZMVyMiUdq5pAbZdx5tEqHmqvnBHFi2qllkntxq+sBz8Tz2
20gna+Eo3ovKs4BDkyoMuptXTtr6dHEE6Drc9VOoWwTXKYjJ85jAzODru3a5
HWPsZv3x2fjWh6uVb5Nu2cqMPB0qmaF4i537+CgAnheKCiimKCn3CVOIXAxv
2XHarDv8DgQWrj3l2DuEtKTtZ8CijfCvWa2mBCkTT/RRDqJH1PNDbx9vSPWW
HKYsNZbR44Bd8c1vUbK1Fb0W22TopunZABkTVYB9e9gVXYu6hvTLET38F8eq
2pZk2HgJl95T1aycC1BRhHKmaaafVVqCHMdw91pKZLfg09cmUH58X4ZT6I+0
IUhtVRZ0S5/2CEL8QuK07OkSEuvx/NPe+7rK68rIas7Op8xM7qxkHg44QajL
TqGlGPqe4OJD+1Wh9CRyLVS4VATg5/nBGz0Cqw3RwWOgQfT8s88Fd88tEEXx
JYHUn1YK8vdNjRb56K9KtXlv+kT4VHTqobv3dsmNJuLEakjUYWC0uMYLcd2r
IIHMx4YLvTT1ftqtOy6L4qW28TmyLsbpmc64l96SD6GlsrPRW77UC5P6Myfb
zM7R7qn8ogXnco4H9hYOJDeTxw1Jgh6bmZ7lCTsy5x1JWYIZ/+DxwzxZ4Gaw
qOOLln70iJShDkuDFgCe9g8u9cOQg05UtA68k+8AX8bR5C0R0VtjLBtrzISn
mGIXYiHXSn7icBuiYIt2qILVKIDq877LkvmvVKmozMNMW1sDieGnO/vtStk7
aoHFGLTF5NYzVGX37qOCGkgepPfn+pIq5lQDLiPNsVj776QivLhEjVbttLvi
3TfSKy+fRUPZySIxJFva6/TgrIP/stMpvyiqHwB7+sEuCqzpqZWXPF9sOU11
8Ak0DcnuuihnJl21JMfUOs6y8Fb8kX2e7usAVqVv/4JSeyazjC5DdoAl7bfM
K8DQx77w+50DSZPaWJp1f1qn6TjCKpGhUrqiD0nlBEcIGubwOlBvDXmAGwle
i0LCiWP/NQBgb1nEzpKSzuEfrE4TIvr8PXlg/q7gybH/C5OcntLSej4HXHK6
OuEDGfDUgImwTtk/YHL/8OTSJRKSvEbAXurhXc2QkxoK/MT6md1v1BLl0vst
Lwjlb4LIypUWbn821pItOEImYPqYwcb2h6aYniKsLSPdpzOEcQTRAm2QzNUA
Wx4Ropz37AgDcIeV6yv8q9ynThXhgrLNwQua8hfTxQp6MjIOk7OInyV6MHPI
33OVRMs9cqa+qvFIcnuuHDTAaFfOon+oA/02xghsvSFPdCjrzDDV7kMcDyZN
KxoCALITTZDO/ueRwuURwioNJoa9idZWdS10YLHmES+bZeWW0JxCbK1Axss0
iQjZaDX2kHbhbEM1Gc4DprKHy8dx4BurBNgg6piYrhrHmhtfltQaAKIX2fsw
XQBxmpMQzSkzAKnQj/e8FmvbMiUJNA0GhiMFew7UPRiXJvZobG/51CqxQPrW
aISV15pKzvVX0KOSIDBfqZ18Ce8kvMY6wdtpQOSdqCvxiMPTzFvyXgGNNYCY
dQgYr2oyKYXZ6kS8YgHPB2ksbU9r5Yq/3pfhI1u0TC5oairkz6tMwmxAE2bt
zKPhUo7BAeLbWCGU4EFfzIick2G4b3j92YasI5WmJjTB7+TW4d/TweixQzOS
dGNAjKgMasU6tK5j80LtuPWyyDusjdoPLfSvE+aIwdtYJONxA4Nb6XgGum+B
RqWSyCPZLTIWdSOq9IrXLNbRbjlf8MotymQo2IZitj4Ejxky24eQQdOQXGTe
1m9R+8hT4so52JowO01I01IvndKKL/MlvIzeZecOA2Yj+sABJts8mVHl3nQM
fLImqbf5GfFsrRyeAYeLPmUAkeM+T/N3/qg9jPuM4m1hdLCS88+B6zdHMF1C
gCzHYPMLBH+j1DQwiWE/tUEm+Fk5WheQe7IeHw8ijGcM43YLuQwobtLhJE0+
eBrgcBMVOlr5l6gDexe0Ikeh5UgJXEEonB8GjzDHiorT8v/f+225kl66ezrR
ta2oVH23Owa0B33Ej3uvzIJCJB6nUzSqkOoZKakrmRc1dqiQxC35MaeNNULp
RAPZASNOEQd3xx/jPrfgL2XOQDga0oicC3U2dYCqJ/CPK6a8Dh2iJE44WYiK
OC9Knxeg/Wr5cqbEx/Eh5q4eqTUNOnnwLPR+eQY09UrjWLHLl3DIykPQV0QA
tbNW5VZsjEwPWc5ab6um5Giv5X+D3UuCLViUAgVecn5moOgOH8e35mhuy7Z1
94CY0rW7YiL150WzipYDBpvtFQFTQ910iV8Ppd3SgCeo2IHMfjNLQOZerh6Q
NfQRiqjMMXfg0/1svGpVf64OgQ4p2CUdmuF6nqz2TlQ2dLVsDHS2wwIA0MDM
lN9eUWdz7ZvKmXMgg8XvSQvetBIWlfNKZL6bxY6W7sw8jPvmeLvGiRr3EXCR
6tg3lZcXEQxelxoE8be/MgYvhy369xqpZ6xb0kPicVel0wlQDBAwuNB3wv0s
xxFrySse+FJKUJezVOsLBBgy9gLqfOQe03VMDIuXDHnZB4Fp30mAumMDLgZb
MnH+Imyy1FmI3Zlxl3O7wB8G/Qeb9wCpTSay24OrAFhvpontQaxqf6l4MgN+
SbJ9NuVqC3QloAgEDAaa1W18hbFQ9VwbjZ1ur52we/UtLVedDe03u3xwchCf
mz9jmKLCY6GjT6YM27hg5VqWwF2uCLeJsqA5sU6srh/RMz8KAaLZisfWb34s
8DK6/uHbGNOVYlhZbVaba90VhfSfAG99C31Rc4bupn55gY/GMiQYB4UnrL3n
uPgKIz+gDO43I0FMWbv3NKIaUATteXNzOHswm5PGMZq/Euuaw2i45DEN48hA
+0+pqQkLLnI9MVjZ5PPBMK2saZMoEdtHZupkWF0ACSTv4Ugl8Wc9L+Cfodim
F4hQ9rJqYgR1jJITUlD5Q5JIinuiaouUzNvjE1EJWkAfjUFJ3JFfN4m98uYp
KxMEt4832m2654dhpAGTOuS7LfIjvcg3FU0/NGR/mcs0obd4zTYSs6XyNOFY
munVKDRoeqjnquwAp/R8/xiEGg2VbdDahmSt7AZU4DIYMw/pg+buqr87Pyde
Lq+E3GeoShOmNd3CHE/rsD624uGAyMkot6+mitr1I9HP54qhxEu81fEKFatB
owERd9lH+uCRaGz69imw4HwzvvOehhJsLA9RNJqntRH949c4qJ8eW8I3qHgR
oAkaMvq5GsgYoe1L82QSNM3XggNr6GV6WjcAEC5GArBLiowy2vaCeeWsA7FX
wTCIZDJMRQ4AicZ0K0hA/p1Rm2oSn6hGtfcHPI/nQUbmjZgM/TsaYsCYpaVT
hiuEs4RSw73mnb0QeWGOvhLvjDihFEO4JHgZLxjHqZLw6qOez5RCu7XFPiem
B2i/Me2Hs8rRkbN8qzVcQOmNJYOZUg+Hyn4xcaJSnBZuKj2q6yokfuPZ5icm
J37hdQ4jmfBTILOt625dK4Cxy5o4Et87UOquiTp3TmmWcm9XAnLM+S6PSwii
Yo7mZGlRppWvnnga0ez2qvFuBSYOfUiOgfuDL8KMxzxsgnmN0hb8YX3JJi2E
BgCVA7cI6Sgdts0MdbRfo6PTAh6eIVunvEHEb/vtXnYxpYz2zQPt+vS4XgiK
ttIlEnJXy+rAiNzU1HfHbbQl16ECn13M67wdyMj9Ykm9sQkBWhagZ4/Ayeye
WA0/KiX0atRz5M5Bpnwpmmd4FA4Jv5XPlgjlwRhJdHFVS1d8GYn8zQolG8oC
hms/HpFtC2LLfM8YKhy/Ezb/g5khMI3szWdl5fkHjafQxR+LtREL8pCn5Mc6
jZfcIG+2rvHp0VEkv6r3tZTzFqgKKb8an7GcYW/isooPugnMghJR9bWbCE4J
J90u7r73Lt08UzzP+CYeQORmJnqL5xFyAwFwjr+uHCHCpn8mBS3xiUG1z3d4
TFEWFp3UhvLfWcOKSihqdPNskpxBcT3x/sXzZftZffWxRRqt/2vTvH30HVE8
A3r+oVl64XwiHpQmN8r/zdz2CEjlURCybsjbtikWLpt22XTXwbOhFGb/5e3h
uJq06IR1Rkug160f7Kjcy35IFaj2DWijpZGj/6o79zhPBhK/qy1GEEbsm9SC
jIjvPARusWsYixNi9YJe8fg76kWZi+DbS4gfmSVYd9lURcqoiY4ID6FzrXT7
X6w8qM9kUiVGfLguuEg8WKPkBMkxN4flqIfZ6/oijxTbElik7xWwNHF5zjqj
IYob25e3mGeJsdQPsbfGoL/9yPanOx1ibfdWGxjsIX6vpbiDzIjBbDpJjiBe
1Lmubi+oe2HZHACPizPL5hiULKkdJ0nGsRazGWjGa/5BqSrLv+P7cqSMhqSs
vOsu5awcPiW3GiNe0TTk50Nlm0HUS883Fin34n9XFIG8W5D4oY1mhk3y2YTJ
5tDyh8lVgxnmfV9AzfvWkevekYuoKjfX4tYgIdvYpRY2yIvNC3OSSPM4KMj+
PXKI1c0hHKRFyFpY1UH1WdBxyT2cYpLRZA4TklTbZwpAYAzxQihpmgg2ffK2
u7N5kY4O3xeufvjvopCo4CUMvlezGza02hcghe2ElagBkxWbQyJI7Jxr7FtA
64wResAqYDQR1hbuN/ocZsse/0J0lkjuvHgrhoiTOlUyiAIr4rCZExQ2TCw1
npQYaaEapvXoDNWwt+h3B2Fm2FhqgWWHmwQQUxIa7FnRArYTebf0ucba9Ytw
SI+oWaSW6NyL1vhmLYXDickqBWNImNB0deyGE+CM5UJJuXb4MjoarScVAbU9
GDhIKdb9gZecobzkN/Io3NETkRQSKziZ3SdIuAsoQ49lCIeBKiWZSbZXI7S6
QKSnk65nmSRQcYInexQ45WyBPIFJbeKcGLV/g1ojxXwxj/Ie8rnzvw6D53O8
Jc+R2CL8iVhOXBO9ArBCuCR0ZfwpQh5UYlkLbXQ4bfAyG2UnpyDYww1fq87A
E7DfUeGLgNBKqHaKHv30/4lp3LI8SEryneaWd2KCMnBAsHUS3mdJPqq3c6XO
pj6xtvNzJSFay7gqpVS4t27DOY6icr+TFYtgmIzYnrE0hkYegZCBP7oiD6Lh
PHHerTRoj1Vymlwtqm4Rk73uAEuhnndY1qVWOCOBrPOxWi1mTDXJUEhh/AQy
KQaz4zjYJctZmnDvE169/OV8CrU9xKND10QAIJgY/hrb821FALJg2PLt3pYd
Za4Q4b+GAhwoKCAZto3krM7v75PGFsFX0WoULaq2zjaGPlw6qFrqUFhLvzz8
bt4Em2bU2X4SnC4Do2kgB0hrAHAcz72gGMm1BZuCXrnW8OqSQNWQOVOG9d1y
cYXvVc1FfmbYysbTBcRVYxOGl7YE/1Z2hG2bYEAriDwkZIafzvzVNoTLuppC
itnC4uG/jTIIxbkOThTVi0vNpT9fe8jd3lhb3sEuA4GJI5M5ihYb+QEeECCz
ep/dgfwZ26K5GxHIdxJKj62pJ6uezi+CCVyFwEHHcLxmimSp6bQ55ah526MM
nW5n0ETTPKw07jrl+3202vqaLGDS0MN5Fbm2Hmzw2Wt8+O7Fvihjn2dbzN9x
O0MY7ie8WVbfqA1ejjmWp4lt+steVZ9Zje10hAnj3oS+iOWWu0VV0WuRAG30
CkYz+1NQekld+zYhwHiZMjpBJvPukBZUtRmfUGa5ySDEE6aNdm6JqZpVKCpY
xYw0KZOD06nejlZPebYBtKDoCkRe4syB9vSzR9NtQwnQPOjWjXlkWH6XMbR5
uu0Cz4hLf+duXpux0mpMc5Q8BOFGIAtj799z66pPA8OpGQp9ZaGwShGc22bN
knDlvOrby49FY98tXfMIQslVprvIFb3oYgp/d1ZnNZ+JrX8vpYk81kp2fN7c
Qrn3hof6WYkB+E0X4a8xn8v7RQeOe59OlbPvV8R6byUTg6GgVhXufzrYjwWD
2baurYJVjLJu/ro5lfhmCgFZ7bjMkGvLimZ5fBauflYyIlHNUoLvf20Hx6GO
uS8K0dv+wbEKxwrThVEZYlnU3lAG1a5jXI7y/QmJfLLZHkvWw1F4d1c9rwIZ
sH2kNXkfB6Ioxhhce54Q/CQETMTuURTzMbhJM3INf6sC5q8FClxG3SIGhG0C
0wBAyoapabM7XEvjkQmBWrHPKvTlFGi+EEH7B2yi1BUV9RQtalag34gz9c97
8MzBCxIXDIiqv71a04BgmwMoidg3KebuXt1ANSS1okpRicuKn9FOyWUtav5V
WhDBG9rOh0JRQgLY8RkCHUqqWP4ELLZqWgDCdQvMqo4aF5X0M33ctecpEdXz
MPvx0G/yMVTWUriYYa764Ej2Q/xRoTQPdKNqx9+znXJMaMp+BTyXw0c8ssSO
rgbOtMiZjchvCsmdLhxkIl33pGDHP5I0jl3JHEH/nq8P0F3czFBqPC3xEg98
UuKxokQi94xUZNJ4dbbT8SzNto91fBolp8iJbVvgC6QfjeZxQASndLUfMjYh
OhZKwwhgsOQT7EoSpTzo+VnhVGCgwZZinDc53cJpAjUrOeMDICFJeiJjaljq
+/xMn+oQCV6p3rGWgRGUCj8Qik33TeAeb2LcosqLHqi812PsKM+pgrVdA6yo
vLmhQGGK6FuDwpjZbZPuz/YspHat4GNafj1bQ53zJEVL2jaTwB4kNBnrzNj8
BbPg/IaCdmelocu/clq0tflo5HvteJdMtRHo77z5zA7ImN2lnV82zVhReIQG
bWUJCfPSOhIFksj9ETnu8ocycbszLRAC/CVUNTRzXStBhIAci7VL+sz9CtzB
lTQCoy91tXLb1Yj9/XevqazSPIrVH3xeWj1/qdm9NcbHS3fgp18h/AEKWt6A
gaA1zRv7iHuRz9BUaVewWeFZhzhO6+elG+Iqx64KMpvZl5ohIXfGXc3vUTzt
I13DSg5rU/+oKOOkP5iZVfiYZLIK/HQqrK+nYrEuj60DdE3LJ0GXSppcyy2k
Gcm/OnIDXUQtiWSsNpf4FXuZuv/sXrdwp4BWQLrGY3zQH+0jcI0ZHiJo7B6Q
i8c7JiaHer/trFPUwJLanJDj/VRCYK5ARno4ikMyjDaT5dVlvzv67wPIbxjd
260BrDTVTnJKTM8xvkf181h6aMBJQF6g8InHuH0153aYjjWw9gBC0ql+IQ0i
0rODDuCzXBv9xnYJ+ys6ZVIPv38Kq1h2SiK6yZNKOp7XCp7mdHHN29IBviIY
muqh16hdg2ghAO56mPtqflsGD+RLLwhIyHuBR4rWO85cTEZ9W8Nor69fkB+5
ZaZCT9JPpGDL1unuZhTN9vhIOxs+sSvBpSVzC83VahDbRZqSbVz3KqXARMUy
583tC6uTrigoiMHo7lmUK6uPxeOVmsq3jjsrgn0+bolze+l+efBm3xiNz+es
NvgsphJJYdrNdDInbERm8fJQqNJU/deZ8gS1SUy+seKVVr+KBVXjJ/5nGSHW
s92yEm39quf26iizeL3R3uYPowqyrrTYbFipPQeByAI3jWqtYRHPxUhN8O77
ahzfpAWeLgAVsvGWEV4aexlLWUaXkdrROQMfEi2eq4C51PbXCEgFmWQNDd8x
PMrLxx7Yib0zIoz1mv93YHVmhiC2srQwf3NLhy635wpCc2vpzWJEgfEcnb9j
I7PP7GjnWYxPYpZVl783oMd1mjErnaEsjPrNB3psNXXPEXDKL6dNEEWbiLpa
/wP6dAiBKLZRW72EA0Xs8NXPKPJw0vsXTiWGNGMQGvZeSPcxN0Igq9hmwWID
R/w9jNnAxJpGX+9aHzoW5ZL4Je0D/TrZL7jbvNvDj07tcxoV198GpplpNTQB
/zMmbnelaqIXpIDCxdl0ixM7X/ecBIE1m6ra+HZGUFEzTebCa4IO2es1EgZi
pN80Bi++xTd4Wxbm/kRqf37u7tmwiTX14Acs/IDXasKJ6NG9Djg1mOuP8QEX
AUOHQRUDBrtd7laAbRIwgxftspnLWG5wDBcdajFIg8UDbtY26CQ6Wlo8Mdz2
VHi0qo34P0vNgo5B6moq9pW+1HJm3AdmrflL2Hn/fUhnV1AhasHJD38X0Hgc
0JeX2hh7BHUGN0U3N+7a4WqoWcVp0isUpHbcD/XxbQU1vKSKUvQ2/f540r8u
o0cIB3P2ztvBemnbpZ+dQzUKote3Ug4tnGjvcMw/8Ijrv9Oaqhdc562VGWIx
DQIMvZpzZxKyKxOtxv+tpMErPMOG0uiMuIX9jop2Hp+k6jjH/SCC+4Lf1DzD
7s4ixXNVerKCMhtTR1fZ84zKJAjtIfB8UaXh2bRk65lTsg/LN9do9jz+VBkj
N6SvQd0rFd/ha+9E9hIDowr7izwUjWdMkYZXtZsnf4z/TgDg/GaKqdgVMKb4
DsDgyBEoDxMOZD0RBOHd6muNmT93+R94wY2A0pgb/4QIs6qLb7R8svKypvW5
x4UdMZI6mXic0hEAYq7j9hAt1d5bFxSjSe+2XHKUEcM5jp/mt+eYI4a2sgL3
P0YBeEE/4iA71j8O/vXAquKzEJiXpUOylTcWbrvRDugfdTTmOJhGzEvx7uQa
Bm2NZN9ziI1+ek6c9IV9Yb22Q5iRw84vezPYo5ULGd9ogaB0QHlLzfLsRTMT
x0/8lxWxAhBZxctSYeIOgC5JWc3g++6CKmQfGPXl/A5MoLc+6n9WGPIhupU4
Nj6TOU+iytDjpTFOIMqQPliYwZK5+Ga67r14T9ONHdUmLEDIKlmntYp9y/Mw
mPQ33GdzuCAjlYkzkUgMFBEagIb5pkAjpPqXM+qanQXVZMEkPovswtYQcWLH
zR/FiCNXgwEbmWgA8MhWfXgfJaBjqhPr2Y6m6sfcDR71yIV0GPnHhfPnsjZ9
WXEKgPrR4euYgdTiK05gBRnxRp0JXZUvnHF/DKsxonx/DTkzIkhj9VsU5eCa
AB4f/qgmZ5MXxaUqtUJ3WH1ywcUQBdJ0GLHYrAyrwMqlxXFMqVIbM8DV2Net
VHJJKP2oe+FMQxTVTtZlqiz9olbdbfF7+yUuEJxC7YkukBHRAqCYSbb588GU
6chkTE9SnS9+v7ddAWGrr1VfTO535P/diJUpi9CN8lFE7CVGThHd7j7pinBH
0o5UrCXfD2LNcdzXW97eTKuVT6Fi2Av8wWuonvg8szfoFdWUeK16h3CPrTiw
jmIP/I0PmGzlzgHgMjsPFjRvftUk1vcSeIEWVvR/6AX0O0VmVFEj6HSqJHpx
CrVnH5ixtr6QZmfhfYEyqkFKn9y5+C3TCJU4nP9cUtXnmTDVi9y9pMtHzglU
BImo0tjnwJxPKniVErUhkTF3xr4pJEY8kY2yKB6uhrT6B90WvdHeTZ+YqCrp
e8G5uIuOn9zPuNyhqwT+6hJFbhP0hmwX+du2TPm+o2a9FS7ElTQTREUNL81h
8FAzT7JP6lgpvv3Tt2cdfATpbrm4wYqBDbIhegIzqMImSZuQkpQ3rbo6Nwi6
V/HOFwCWpIbr+nd8oYlPtZ3cOCixBuaDWgH+N81jhNIJPrflP0WTLVwtZG8P
ce5i9FYdxv0VkvgAMnNofYDcQt5BStIkKJBzYN6aOpuCo8x6bEE9xK/BMwIx
vmjqjO7u8a8qSvMjS47QqA4kMwymrz6f33A5I2kJX66kl6xt995UMURBZ2Sr
uA/NNSBHfWzl9zLaZ0hxDQp/Uo+giTiBUI0spGlQgDaZq4ld7ge+K4aM6jjC
EAvF/xqW7zBH0onu8z/YR0jHvG3ouQS+Rk4cV4Gk2iRx1Zb3Pk/hyaCq9nq9
24qpv2HfoWFELvVcRUJy7t58XQyJKqxEW20cYycZ+k2kjIcODVVGNAnDRDhR
4PLX+GUOwPyRDY9SwPxgehBsrdcYJ2OCu40EhJW4VtcBvYe2AkPHkloE8KsV
wSbUPxlM0EtEPDELx6IuOG54acJ5quklrPbla5yucp8Rz3U00/GF4EqOh3jM
ViOx+t0JBiMfYiyc7nCpOU+Z+025HFeGx3p9X5Dl4iiWbmuCNsQpQCfVi3xi
OKvF+8tkL4s9kGPXvNl7uPy/0x1gCFVOBeMMGh9GOqBtyRcBWmpmRhFyF5eW
w8CT2OzDESuB5p2G1je/MagoOI8Tf+PCDVDZyaKoPBFDoO6aeoOQCH5BjoU3
gGG5zOp0fEaNyVY4vUUAKYGoYOf3mV/9VtU+dyAD+Jk5E5fm2pMQDwaBKuQ8
Fb+Yc6BiC+ija+PJfVJBqgcIUVU7sEWWDGml9PbBbEenIMUl3EY8bjVAidJu
iTX2TWXb/FTlWzUaGV637x4hmCim4ynRRt39bTpjXwn38lsM3RlNtDZ3kQVQ
rZZp7/6+ypnZIOv7Msf+KMpdsiRH3b+TnB2BXH8ZYcjD8dCdLm77Ctg704BO
2beNJ9ufkg5xuLPYsX0QsHZfMGR1HRf++D7EDpQCvJou5asWses59OQxMsC2
jZbfAq/MoNRLVn39UZDKCZcwII1Ov7DoA7IuecJquOhkiinymFDznF1i5ixd
trlCIsmav6LuymJYrC9soUw4r2HqoZ68XBVkyI3feC1pvn3zoanJ3txyoZ2t
pyRxgSoEiAiba/g//z9ArSQR8k0PHzwuykJ3OOHhbAQxzOHyTC11h75vIao8
zVFoPhxXlI4nZo4sS4a6aHeqgqyYHPxo420GbIdB39fkx+ah05RYAI2po2BN
nIKGeRsLraTmj2mOAYdmG2FI68wM7Pi30OCBJBv5IxKH+m1ZdO4oQcPkrN/r
rWOSudyP4ki+GwX7JEgBm87QKAu0AD5gycrfecOAX4QSn4P7JoVIO0iqQhHP
3Y4p768FNW8XH3CmJeIfAGA/qZCTaeCZiRVfrOtpzAQSxLlfMvDPWGC4W5xi
k1uK/dygCCcKmh4YFDuhzq6APtqmY8GvfePuS5m+7FYYWtxJiR34wNwjau7h
H6bK8OxLXIiM99UUXUR4t/rfHMZewVl+RB7el/2payossW8+5y66XRPMuYW/
ft2gnhGIyfAjbPJUILWxkz459+BjCD+pqdreXc97ja/S9VS8LMo+m45yZmsF
23d6aJ2FOclLs25aas3tzO37g5bfcTsUlCn6uN7dXXKfQtJx8efybKFo+Sas
MOTzFKSitQ8TCtAHVvT5FrRJ+IS2IqmL79Q11DTONGlfBQx2VOhbtlUxfoQm
c7ldK6JbiEDxGagADuOU/P90n8fK61G5UqiWyT6gt3PeA/eQwj4/OMSnFX9k
o2vWSskDGafMV2HpuYCi7d4IsIfOdrgbodfrydX8MhTnjK00Nhs+FLOK/dvr
R+td4KbtLv0EMK8hiqZbTa9rZ6zTqwnD1OitrkkY1J8mKtCsTn1b5i/zK6uf
l+YS46ZTy0ipDVgHHojPyu9Leb5hiTLFI25wyWQc7CHbNsRJa/BjtfU0DCxh
PrVYykD6Otzs5cpUGW3Ei3nZeDWC9xUb8DbLVaAMln9tLQf3ZHykxUG0gWE8
+VKwSgFAFzWLX4h54B4FeVMO8FCMdkoM280W+46RJjZ83b24Ag/05yCdYc1g
/bP0G0VWgpAVEZI3NL6iGd7VhxMr0drXcdmHvbrc8K3XL4sZ4QduZwThLUN0
QdfRCVqB62fZU0vawvb3cOqrDMkQf45nFpA1eXNXuTPweA6yy5IAlS53z3re
q6a0znh2sbniDCTx+rPTw26+qaMEC7USQEv2g9+GqmOZtCk5+i4+GM5ZfHiD
rgPRUAQW5jbyMlYSLljd1kmaoMkqKOLL8V2N7QfS45ROonXLHPLP+NLXCopr
8pnSfpjPlQrAgTvWiUXlUrlbbKfnAmPD9jod3gTT0P0RcNJDLelIB/XdOe7z
9ZUXgKZpzgWmUEZ+PUeNHm5SDNyyapvfPQ27V3AM6QJX9nHSC9f4nBPzm57k
+EkW1nLUtal9V7TPbTD2RNwIjvVrkFPWEo0h+3UfeN60K/pletOt02g1XPTS
3p0W6XfEH029q9COMKx2VVt5beNtViw4S+FkzgGF2Z1kOlBh5JimCTbURWG/
jegRINq8S6RsGQ8yhT504BPQ1PT47e59/wf6GKg9knrbGP/LxHBw/OMJwvF1
pIqJxlEYSlzq1bkxKdMydQHezUp5d0sk31KBKsEJMgfK3Qrhd4pnMJI/ScPX
/LLIiqMxCitQFFF3/Ym/hUj9z+CnK84CeJRowx5b7laP7G8j8V/zYZPQL7Lc
2vJ1gok/KHsxhsa4K5O7UeQEmTHVy9JHJWj59PaGIONGjNhDnTujnTdTjYhd
03bL4u15KQqw1C+ilspoHjvXzVInjzCR/9VcBfzp+OLnaUaLZDV7JiarckZY
aEAV9VxcvFW/J2YK3CxkH6wXUigGlxFgB9uLNUWBpiLC1NmcWTw0CKKWHYVd
npiQzcTvOR1I8dUrmehVVM03Ay00JLOWNA61Nn70QgnlVhm7pTNam9CtOryG
MBzW/pwyKiXniFm9H+sPV/i7z6bN+LgRLnLz4qWcZQ6E6aqnqw0AdM7hAcMQ
s1L9ChfTJYCh2nqmhpnO7dNDdbqqRPrxYt+LjzYvnIKJNhI5FihILI6FYr11
C5sYxUn0TvDHEq4pyKOk7glZN+jhCgv2FvcQqbY7M1RKLCT8T85QlP/lgANK
8e2fxvadV2XrQMsgk4CFUnKwMj3G8UBnAvoQiW3hELzrBt7X4mi5qELuSAsm
z76bBrpMgehFFOJpBiLnd93a59lC5FIudWbh2tICjTcWopw7zUpZVBEFzGCm
058ChZj/3CBBmigoh9noISeUf47vJaboZnJQMw+lZy25MUkQl50t8IlPf56W
/Pw+oVAgu/jtuEqMadzwwwux+S7PEGJMD8OMLLNOxnPjtjMqG4KhXWGDNPiH
ai0y9wZ+Nf7r5+JiEjLr2U0MBvMQ9sYE6TLDnZcYqxHDY4U7kwkH0RotUszS
EWCSdLRh9XEnuQ/5D211mzIzuTP1PdaYcktKBEO2N6hj/Ne3ff02hjkxUZGc
kMuFlYMKYV78biMB5/dGjX7y/WsT11HpAcNKJO5LiCQ3gUPuU/zC42znqie2
jEJ2FokPe3Q0Ee2eY/XEvzXTK/2hBGAQrGxIGdiu/d66juWiH6wPitKUQNaO
dBqAhxpIlhYgP0KysNZS/mzpy6rXylEvW4kODM4pQxEpMXBm+5XrAkGuY8Bb
iZ3WhyqrMYjTFcPmmH5Q9/3bEV3svUGppU43+DtOk9QexxNHeyra8Q+/jD1o
b93UrkK6z2x77vbp4RImo1SDNqiSOlpC0hgmwtTVB2MICM3SonVu10npStuU
xBlND6N2ombeW3o/o/KPSC+8a6uX/3NiIypRX97uEDzCzHg0TfMgqiak89dV
r6Acs15N3VPAk/QsKoaMoR0oaey1ZBBJ/82K7nMzRL11NFHf67E0XO9fpGEE
vmsTJPMvJ+/JymlMT3ZDQzt0lPCp+KEKEMZ9ItqgrvCivXj9NcuUFZEhNuaL
z+KFuGNZw1LMRB74AafvIDgDOt4sa3UlGdcRZC4m4Tyi0a2QTB4MBzELRVhl
ADiElmKhsQ20f0oADnKZce89YqRLTb6T5rDFXOt3abXdUWzHG4nIFwD7PRjB
o4TWeghtfXSiB7RPPgw0pbSLe6iWdrU4R5EJI7JlJTgW9UBpZv+Nrg6c0h6C
XTFXyAS3j2aFyHa4BAsQeTo1f/7Bu0UlSfrDV/17IG1NNkP40I2Oi8vyCGvO
qjnUxu31E4wi0mi9tzjr/AZ+iSQWhgIuI5wr3/NUD0QhB9ca/jwkVzQWrZE7
H4FX3R6PqYun2os5BTTTnMSdZFtEtaZYQfTeLnLwsvKTNcAel1cSPyeXufY+
IZs0l3zYVpZJ5klLwaYIbLFYcS/i6QPrnkRjPXC9qSSkt6d6pTsYA1txsW2d
PEwYfjQydsJiwDwzN47PgI29/KU+liOTNearvZXbwH1opLRRrhIw4axoDqhb
z2U6gOnlcDBy06L7weWHe8ZU4ab5m2rmXP5YPxUoBXs36I8dUxwADfkPlyT0
Kkf/wjqjB54AnCeVOOLU7AnWj9v9TiIQkQBPIQseo/7RNPZSGvEyJVlZPeCY
osPfMQCIYLMGOBgurAKZxG9An3XHKkJPWev1KsuRqNcQ+bvstoe3T4yghio0
g2DgWjPxqx/I+MKXkHKCDOZep41UuDNxaOgzfvuNKWd/eaFyzwfgDB8YNv8J
jEb9c9PEIiddwQNXnkFRbpSrX0IUX7AVCHjO58B7anvb/Ji4EmkVhDNo8THS
+vawepYGQbnhNFi4c1JlofFKKSsHEloU+PJb7aWQTVbmvaOGAggjuFxRhe4f
9pdhftimUFW3aWyXiAKjlUK6htXPxZ3dGg5gbu4MCRxiqEo+/R0LEjdYWOTZ
WesnaVuALYhsz4R1sW/FW9IcYGzf6lGpDkIEXOnmZQdwEz4zQbA11w8fJwcV
nMQF5uAk2jyOHXjCcuGwCuW3N+r3GvsUgoJnWDihRHzciugSI3ND/TmzBUQT
gVnJHHaDW/v7B0Ix+szlYbU3CGMDj43PdPamroyLkfRqPWm3+u4kxF9dLw2Z
bsxfo6/KiLF4yWHNoDCFBrlWWC4G0NiXmHf5JbqT2yR1/cDPiBsQSIOaCGpt
pkk7yrbZgAfR+n/p6Mv/GYTKCYi+A1ntf8LTwzTzh+hRfSe2YQft/rbFMLFy
wucnu1jyZPpwY7m/5J43Wo4fIYwl/3pL/MtxII44ZWLiBGLwmD14yMQDkV2y
yR+IDrjnuZmdOxZOFloUDXeJfcc0Izri/J+c0JhCdCApJNswVM24vOZ+D0EC
T7ud/dMC0Yhc7KjeTuuMRS8gfQV6OcuUFzdt8mCuJOmF7PpB9jx0zO/HN5n/
n7u+cmj4eN3LNg+WpYtPdVfA41+/dgg+Jut5jjcO10+p0h47JeSDikv6a7JK
qUexRDCISXus2JDJbl1+cfjtO4FpimGsdOVO8p1HgzJxT0FLKTZfK7o+u+KS
xalvsw4uzgl/e/qFH+KJpkWvo7hlgt/LjxwhVPBYpC7iW9kRdeJOCh33prXM
n79sUyq2SfKfGeK7HztRAHYF0Q//Xr5me1dpWftfb0ip1ZKmyBhPVo6W9XDz
ce0OdvfmGFC00m/PyF6PRjnxIR/h6ZlgK+BHGVSA1tSob1sPBi9Xl7zAeRRL
Q2NdAejdIP6SOwqiwfgp+pfeoskFl70eAAksVgw+R3m1QPXySUEHaNg1fRFN
1QLdnlh7VFei9l4+nZwACry1Jkdm8dL6dtTxaAETXPUVoQ5IF+sd5ib0hfb6
aFHut+sWVIgwprjXOWnDiLwuMXYAWRdJLhZKdtDQeHbhVX60Qyt38oUh5Udy
t2aIFRWv3UUKYtyFi9mrbxNoZe9xHNElHhtpWOaH1oiFiuVaPWVfv3IX+KTf
5ZVXgAEdeoJKzoybjBWhJPk/ppxG/W6zpKFDastjmD/nVim2phxZBfXqFPS7
H0y2wEojvfsRsKwRQ7ziNXzT1z9XBtLNSDtb8guxCWmlAUK8oIvHy/VFMSUR
vNCIpFbeuBUrEu1D6H6zFae+1K7RJBqfSSzYkzWaa0QuPSluet6xO6oRh0K2
FwWwUxlFS5Rw3gMHSHf2nUK+qejvhMoLbXzhySxsF1AXeGddX2cvpntiz6n0
G9mYMWRp0q8XMjUcUFsPbls1fvRqmGuNEVbu8LPnwOw5jtUbZH9PE75gim+N
/TUNMVPIM3xGTrBgsG9UR/VmlPIhULqYGOhOKE0GRZgfcOgS0zYubISv3qKi
NKscpX11WAjOqp4Z3uS+0b1jMGzhVzjkxXFNWxXK+tLXpF1n1rq5FQNrv94L
Gk+Yg/HdKeGgQKz9VYrrU2bYZh3zl5u23Da8IxZ41T/IRjYYk966UHIKqt90
P/tTfERRo2kxLMZxr36c7MQZtLic2K2zWvB4tnsk48+L4VNvty7OSQHmXmW9
WBufxV7Z1ysaJTqnnezm0mU+AN302cPDzyOBXBjOBjX9gOgBJ7hfgZG06r95
ph/gKT3yn3zKp2oUqlaRizp64mO71uDv10SIlV9nRLsktKV8SsOPxw8dCxak
IkRoz0Q6YaQIFrWw1aCE2V7cKGR/UtdyzMN9h6Oim5CspH14izEeadsPwa1H
D0iO5L5jj4LdKjUbGJzQvifansWijT1W6KAMThFQsMaLiwQX8cp7WTybcBYQ
6nEEww23K0u3r8J0096YHs4fBmFH3hgspX9QFka5aeibjsFxhZsn6H7JTiuH
A+g6/MOwtxHgQnnkDwM4vbU9252MONZf0KELuzORzBl5FKqRj8TiagzUM9w2
fe3zvbFDMnadnJOVGmy5Yha/SJyAACXbPAOlezjFloe+nGZSP3hQNOyvrzF3
3MTLhcjKCfMGjqZhuUIE6i6hsEz9uqQKBpeSQiXxug/2TZJvqqUoAXS5YDow
/ik6xImoqNAXJeF7eiEfsXMBf83dRAQy8ShlPkbv0TvBNOlGREX142vgUjGZ
OD3896vE65jhkVrnBtUkhRULVqKHWKMrhIaFZaaNDnY/avLOvMxfT2Xe58sK
nnj8sjFKewmDM2JUm/pkBIjaObYmDxycPXF1KvwCaa//39sB/O06366NCpVb
Q43AfEvcTbqqp0ErPZM5z02f2zhzVuEmxuaIH+Dhc3Fgwt2bs2WX2Dkt4vs7
e1oYZW9SmLoWSugwMvWjiSQfh0BEIZlaYIUq8fg+AZhDAXc1UpIdIOtJXntA
79qS6QE1toXFYnNaQK3ZwXPRbZwbt2C2TdGSe1v+sJrg6UhWT3/dy8ahy1KV
9m25hT6kMHnrk+Lte4HUHZjb3cQE1UNTyZ3iPo5b0+F6inYUHanec67H3krN
bIPgp7iqgMsS3UyYVsYEWpaSx4LE6TO4wu4E3o1N0IkqTW9Xx+zdQ0imOKmU
FPNAYvAsPgLUf/vszsyPp7BfjgaKwhj1M18EtVrIvBJwgMDshT82sMSJO469
CN1U9nBPzewmNPqTAkvxwLyrWWqKrhmfBKgtRjCkxdJNow+J5ysFCKcy4PD1
d9ixQdv9fNnvbpeA2NTlDFTYIJSJmahz41pweJz0FvotDbqwB7/Ka0Xlvthl
J/IMeczDfNq5j5rdVch6eUFatzG6r4tP5fA9qCvAcBCbnDI7V/7xE9WGvkmo
7J152Ww60qlurdSzm2wHKQ7IzNBahHIWy9pR38ByQthdvKF+TnP8vKGvdin9
uhX4+MxAhR+66+6AOBj+BKwGD7Aq0Hn7iYbSZmt6i3jjCBYWtorjzKV2hAa7
iZYaezSJPb5CR124mDM8CUMlO1pU2BuWtWbVYSopCvm43WW2kjMLgUrrzxHU
2BxhRczNfZsZxZNI9adj/yh0y8LA4XInkBKrkX7AKd9bLKI+CMpIzNvEubN/
We+lRf/CCISS2w5PeXXdu3bTglE5nmxreZHYGdv2a4jkc6f3LU2P8eQdEl9w
zV16Jtu3xCCkWnlG2i3lv1Qiu/ffzs0EXhGi6FA0eGo6ltoyHQhYO91uJu9V
k5Cvd5yo4y492SzX8P//lEc425pNnPy/HdT+ZEdhJEEW3Y8B+2AX8USNWofa
CdlS5sdUKEclJ2u0noZFLurYcj4P6aDlm6Cs7YzUfd6Suzjc5pMvIrXDDgpL
vR1OmgCGhF0vcwWGTpTZ3mPDAd/Kz8+q67fxyfAKsh7O1ReYX08T9qkk+MEM
uUOvN6Mt2vrIFC+XAJzgHQKP2l1TCCKm1B0kOD5/6IZkQZDa86k1jbSNs6B8
0P15x/Z2fPKVZpI4ePXfaqizbwkeTGE1mTlGNdIly07j6StHhitAd9piuVUu
6DSlGUtsQ93bxgrFoKE9f5SGJiDYA3mb0gogWOJVZ8NYzZrGOUKR1gPdXEbG
MKProXLmf60FTzzLllaBCFyiE4y4LQbBpzlt/iywEzbo498BqHSbIXxxklDo
TAALblgxMPDQiAs8shA0ASC4CImBCHmOH8mtq4jzgUrhPHrCpwOXDAdEv6ew
HwnEETk5JfIAHMbso8WfYsM4Jj7j0JZa0XqSshXvKqapU5k6g/tphsKxTQqm
2qOTMvccXPBKUaKIItNcG673aknMGJ20/9DAB1Y51NFic4yszFeJE/RqeS03
anmA/BdoYzwIFn+cVNDsU35tjM9N638lKrUuL7mOpLkPIDH7+1cx/3Srb5x8
RwxinQYTKq1P+G9+iTM8kP7ohZuq9J3lM40N9/kqkKwK5Jfz2hl7EwDb+4B0
Tsgk8uEqGjNWfT4wyzwiRc6HasivJEoNP3wQy4bHmocBYdpsf0RaYLzEdf7b
ZCIKERkxCFhjXXOqHcNg7A63VCkOqrsWNnKN+xk3EzeQl1b2Ts0MIpwsR50C
bdG3w7F4ZBmcAnEd6hLC61zCHUgBHUP/QBEW5C9Z6lMMXH9LKQeDqA2AuqfK
iFEUADtdxw2uYAEMbv6rFm9265sRoF7AiGKVw3yz+FPQUBUYPS329JMAioHX
/JLU3A/YRuymOKNo8eDU4P8BAFK4nY1xpIvfY9O3qFDOY7ccIwEUSeBta4iW
OHpMiVRrGRS4GxwTwPH5VXFyXwczFHHUMtEZZEslMC+dXmJGkTdZq4us38iE
crl0U0XovVUZFf6QSbBd83hqHwHAFsdQdbYCS4fvT0IzGhRWyLITs+FsiItg
FyB1BkzVJjgId4hJmeg/j+32gpD6bhOUjGzZ9OmshhoPozvBaa30rKyPmuid
7KbSs6hXgffy7N2tEiUK57nOS1m/Zca4UfVEvsS3VOpMW0JDeukvEgx/IIB/
7XpvNK8zhyiwn8QYzID6AcDYiH0ZKS3LEqYHn4JetX2OxjJ2xScbzQyUfcOm
FffTFou+PIFLnkHQb1WRV7a4n+qZ0G9fbnsmdJbwmkMtYx9dauFAW6/TalKh
z7VGPeRH3lAqUbkJL2PkNaarU5KlYnuO2C6cm/BQtUbVaeeSV2yPG4liTtX/
uMc++UvXH9A6Opdk/vgNckGsfTZZOxhKwpi4E8pYA1ls7Ur2JDa5scvxETq3
4SY/OvCWpz2k+2WoroL1KE8pPGPUzQ0MINxtqruIPCKeVJV2Zbdw1RtaiQdf
uMq8YrfNum08XDXiSNZ+6PaKqwhcqSsV2y9+xVFAK5LBgeoRUMRdoXAMdiDN
u77FrF1bU7zJYEcYqy1bpTJm7LGAYBzcPrQKHr6O09fxq5Ohph2xE6BX9rYb
akDxR+YP7owPON05V93HVO6wnh5rrvznl6jmZownYEOhU5oUF5g6T9vee2Ba
ztV1gzAosUZ0U0pRZLK4zEhqURHdiSrYEM8QhmKiSaRAsDLvBpjmrCI5Mbej
qunyP+NTbIroBVxFhReM3TBF/78hg2lARKj8Ae3b6lLnlQ+Ca09BKyRoTE7G
R6ic3lTvayTeq0gOUdaLU5dzfdjZQX7mvf0rbnzzDufIAHc2h1Ml4igyU7Np
MwSGHygcYZaEErcaPEShPX7Q16nMeGqz12v9UAMoMXJvxgUT2qFBbra42oHA
RILsSdMbGlV2EwUda0z57DRrlE9Xd82BuzVeDMiAa+ecshS9pg+1NkYmDyyC
0ise9PA6G/CY6TiWAhmMivwBu+4q4pSBf5s9jxzjLwk4S0nIpYnmqjTsp7SN
lljG1UaxALNLjwYJ2PQhNuXK9wwpxeNNZkqki8yX7bjDjlrTJZLGS74ad1Ny
I4JqAmkd+FuSj48st2uaPL3eeTWDS8Drjg2BCNT2dCZPLjAcQIz0x777y4jk
jRXO1lHuGOIwsulxxK2bNjUWb+FyBOSjTZ4W3p+nQSbAWNSekas8JrVI2XT0
snA8uSF33jo+UhbRm5cnBv89plpdGieTM4eAnYX/3kx7eBXJ/Qh+XuWrytE4
S3OM5eGPSa5J8VGKjneEHA6U0Ua7UVsQuyHfPBWFl0xVXZpHYy+h4nrovYt1
my8DF5RMFhr+ufa5YThckFAzOEgNm1CiQP7wr8YBhfIZUrLl+4HfMk4RYHZb
EAvAlSepdd39ltiSCwiFmnpdLG82AadcG9vkryQrmoY5UwMaIiz/XEpTUEJP
qahXYm8+9V1j8bgADTX4GRVefmFyKvjlBrABgPqTSXuMZF+V/p0D2lbiaZLH
MHwrbkE3HWVkWE6wrRoowIPfBMVVN+Ie+v3xKqMoeFZY7VCDTcwAWuwqj7FA
Hnw5kSIhWz9STNbLcNFSCh9w9GaZHr3b2SMt5GXalj6TZCMsOJGK307H083S
ubRHTXTiFHmKAdjmW4BYYwEkFCBYEf8v8jr5cxYLECwISpbOzsqdIKI+Slu1
D8dS/DFmxg6pMcQfp0OXav2sr7cvuKYFMgFGpzKi59EHVr5zhM5tTJ24jIDJ
hawBJSgli/T9wHa0meSsevEOeMcn5/N49zb+O65bgCCNvdy7SX2iL29lqRBi
8RjmUg6VYHl2sNHAg4TvHjhSt+y096k7nhW9RWTSOhNmyB+vK3BKsBfRYv5v
WTFybRat2cCPctCgKGXYtst8YybR8xlswVcz+wq/9ojncxClzQknZwGA7Zn9
k+dFb33CZSG2Tj1rx+zkSvCwHOqUDo1RWuWCftVwSJ0+N8EXSM0rvuh0Q/8X
sjtrQsjCNazjeMApwvhy962Z+P6r5s3sKaHGpKINYY3pYsMxqP/wVYFozGe5
glczkGfJXrkPT96SC0vwSbAa6VDKoNbkGHGM2UgXCTrYvrjGKaQp9VBkmTth
qOOMEw3fcHjieQKPLtLwDVHdcMHg26cTKtJUxGntmiVVhnWwutnv1cadtHIi
AKLyHSCW7R4X+mx4KR0qAtVnq8AQTVOtiMNsqxwAGiDbrbIaMM75SvUjXFKN
Vz59Si3yxK35AXu1BjcbYwTHU5T5I30jzHKqEK/ApWM+qe2JPQouMz0t7CaV
HWgvNePv/EYn9mo+0T7NnoMiO434eGqU1pyrjnBj0MIDpb/KKZwx6ONQ0uMY
y2JAfv/guVRlhmXmBt99mnN2Ldtbx/+1NUy9+hLtEBJNv9SwdOaqltGi+E+7
89u8IHUOFtyVz8ZzyyhtyqfLpl5eq4E0xXD9aimu7VHHglYAmLH9hfnRSaTR
Xd/o/yt/hirqupbyrF4zq/OfggRZY2o6NGXXHvkI72Y5pkUyzv0DZyyO4icU
ghfcBH4xyIEcCcP7+hoUUmkzWRJYCFRM3bBzZmW1pT2e9O7ajXpkUYgGjohb
H4QNyuW9gM9AJGeyRLYrGUj87XRCx0qFvZbCx4lY2kiPPles4B8kjqGynree
T9vsqtYAZR718aq9wNLeeopgktx/pNVar0ADmYs5yLqZPb0hMV4+kKv5VRr/
HuDaXoEqyZSyIwMKuujAeB3bxj/KtOCdL5gIGD7qZvH5rLXiBRSBXKKtGwBg
NxXF7dr4qVU9UKOV4u8s5MNQc3ftcTNn2+U3LYe+i114+KnKiYslDuqapJvb
jhvjI+zokLCjyTgX2hPa9SfkU74/oqUD7D7hpTesW6FfAa+HrmxESF7EdBgS
nwK1Yc4zC0ezBYE/e+lFgjudMiVqi9cYUyX7M8zmrfb4Uq3QGSbjIVJRKlhV
6IJB545aJcRuIbd6cGyJmdE7o4g9xQJrtAWmLHvZ86uccRZ5A/dtp5g7o4+6
bVGNwWa5c95rvEU8rteH35KE35LQ8V0tE73bH/K3e24zHQwPi9R6aRZ/Bl2q
ZyzTnTaf5gxXTv4Y+FYGyJmvrZtle5nILHCyU3QLmAU+SOf9O8DEhn5iu4Mj
6SSS23KmacNxqwZSjADlklsVYHDV8KniZSy1GqeDI631v1jcg2AoL4YDDHrA
LS5RXJIFnTn7Ckj5gTX0PQuolak1ZXjmFFrS1qSvLP4LaU7Djzk9k5kJ2IpH
j/hfPK9gpEujmpH1eTkhmXaB+IdXk7O8YJbJcgmFFput5gXiKGhVpeDfsDLQ
8a6mo+Sol7E4m/rGXtcfaOq6g3wYtnMra0p1Dm0vgNvR20fcmvN2Aj/sEgId
jLpuuH14+MIwMGa2rvYZG5HNSpDveS4Lxqx/dTfMVkQaMpflkXxLg7yQaFlq
Je9+VjgnVg1PJ07BF6Q/aHXxVk2e5iJMzA5n4DHdE2v5JSMcnwIY6kvNSbo7
MhqDujFB303Fz44fLFSE+wAVRnkzeW4s8FsFxuwu/s5qqpgRiEC9RoIXVfl6
RAvbpknNjTBJBRPwRGiak0sowXn9LFzU63Hyl/6acf6DrCyBgY0UifaAZrvX
5PDy9AGLvKLTlRJaZcgNyM6mFYudju7h+mqsCOIYOF1pk2+bvwAH0PgRX/gz
ucAgZtt1PAxo7h6MYc2+IB3eDaDGD31YUZRSpknRL1xHMnNJJThZmiEpa5iM
gScGEiBFS5p7TXqv9JK2kf4OG9k9BvyVe6PxzorOk+xUUCEnhFVVH90Q2jTT
/kCHoCCfVIx3Pl9oYhhj065uZCg3yhZNPwYwllO52rVlOh5C7EgLfgI00JI9
K7iqKwGdHgapywTfvwUpTuaRHbJL/4yloDmsXMJpX5pAj5/Bb7UkJEkjDW3S
b5vYfE3P8WVCcFlIdXvzfRDqWuqHLEPtZ0GA5vRh8PPz2lt3z1giFmM1E5hR
NoYB7voFZVFNKrUPWddDt4+R9s3lM8VRT98WnQ2ODY1Od7cpR6C1Y6am6v0h
B1/0YeMD8GvN2ywFgJeficTA5md+RCNbRhA//kqqZia4V5WDG1GTula71EO6
GBoEzaMluwVsLXoCdX73wgJ3+S+bAdyimhAsKGdjOWC+lgsdLWQvZwfACVFf
ITEMcz3B+OPdUUweWdzPljf8B5L5r0fp86mABbW3nVRnAgMpeQTeH/uxdJBe
+hYX1A0LhN4ddn2nbbzzATIfcjuY1mpG5VTBBJ+hbB0ROdX26nZvrV0UAQkc
/EqtF369eWguuN9HbpNQKNzlzUtPJTNx5+PXNCL0sVb2ONvlU1N4AR2FJqQZ
lmqFEzL23ibLgxG2MmYQ8ivzRaOAIPUbSUy4Bkf8m/eYxy+uVaWCM/OsSFhp
+r4uToRr6y6E0/tSdqGWtF9XHAiDV/WtHjgpTu5LEBjH1NRz648YeONR8R8T
5M6kvXir6bt/fNuHWCqr1pcTmCblOLgyMxjujcvDM9X+YCUrln7QBJjHEdQP
em7TIyYsHxpufts1Yj2pWoN+jNw5H6P2mr1uJ6YHcDLs0J3UgWxrC7MaqE4k
cebISfw84T+x6cuy8bSFDoyHlK7+MY1faTYuNaDUdG/hI3OWkTfxgJ8qLIWK
hrTzQEHUTC36X83Z0UTEnMunBc4oK4gn6H4AXdoFK5O4RGS8OY/y2m5CcUlw
a7sJPvbz4j6VtfawQfDX0IfxZ248Msc2y/2i1wZSu942yvao8s8y2CQLguH/
3ct3V91161DMSUd++5NvrrgoCp+xbOTx9r+LNLzPdijbhhRJc6y1WxATL92b
bNidc3ku23gso/GyrKE2h8vEfJIVxGBhmlFS36xm9046roBWUf5OtgjTZWNS
WrYkwuPiMG71kmhL25nM3R1wqSjUwZLWDoDYlKUo66gYk0xIVktXun/7e8sA
3K0EVpJwHkXVwHRW3wJRTXPQdZFipoMr7Vf+bU5fZOu87bxJ/mDXSGT97p0E
HgiA8CHdkjGypHD75h3EHIR6qDdDDwAP5VJts6NWUJSj5BUacrQcyOOV+SSc
fk215UZBxjZsDreS3xYm2xWIfHRmuDEwemTaDyegTcGpesFDH7gJnnjlLCSY
4FE8d+1RSR/UxNUN+jMX2y8MapmUYCgdY+pMU0T1F5ugFVnh0VYJ4ABizNvX
8lDEP+f9RHzjpCc1Bbp1OQqZnMdQLYg0edia5PpNVuvw8OWEF4QRXPQSkuVF
D0dHhmX94ILLdXAXa1vfFJiciPOtqqxq62giMAMvC2x8QfA/XLqW0ESwTBL/
jjY3zrOqOLFYu8Gh2q1SqUui/KfsbQhnaFZcuzel2og+j13vnQanKbrqPaXq
CP2WvQrlpus1Wieb3ObKIekBjctG3ocT61PsAyYNzYz+XBe8gIfGLxSf1UkN
7RGLuTE2mmYuaktRJ+XUD3uDoERlbd604sKRpfi/I56rF3+xKq+H9sfc5KKk
f+ge5L1xoMCva65GZT2oab7jxnmzK9K+qGjY029lus3sQlJCmpnOJuaV+3Bd
uC2Y2Hn+kpqlbk4/GZ1eeKCTva3m6Y+jnfOgeTCCn8Ut5wurcaxSHVfD6EmH
nE1ZYNv6qAbh8u7hY2lamgxhwSHinB80Zo98rVNQduhTvVFz7bGddG6ozPhk
yQihd2+n/6c/g14CwkYICZVCrl6fJQhtasAfgRMjMpKUSQv/nqhUB7i096j7
fdJvdrV3mUw3gL9iuG0IToMNanAo1FmDbErrRE0VgAOzOP3qugmY3GWorLNb
tBGFnJQh1f8UzG0LztESFh0Ns896tg1VcUXjr92Ncz71AMKwvqGUgfGvv5dh
oHLCMaA19DHLEWWbcSreuVI9OflpkaclrzULtRXPZUJFXDaeKMwCJyvzOuuI
AwA8/A1UTGKoGovzn5UEQLP2ULUXXKsqu1G1vcabYgdwIckIAYw6rCqDQO6s
cgTLpsMmt+1eL60UceaYy6eIiwyibjTyuOzQ7qz0HCQ7gBxCmhUkE0kB7Dg6
E7eGHaBVAm6kT7nGAXJPkiwB4TUIqCqWFjb4ztrYsSoMeCWyDzF2vvcbD5Ss
FEqvjTREKo204WYR45b9lrBrxx2MpyfgfoVV05nV3a5Z5sBEptPGcbz0qjFM
HtmScxNDv34Ypuhf0qtqK16DUaryO/aLBQH/dpubTjwGDJhIqWPP4Fv7ovsD
OaIltmDSZhy8uCoAbt0lYf9psnyfyn6AtVR59wfmW8ytlUpKK7/0ZH7erA8C
Go08GaWeZNM2mkT5Rsg79bUuXFJAMKXBc0/IhuoYIiC6GNrtFmpEoa9PFrvl
ol+nvmVg2ifO4C2vaaBKZucTlaXMPMFO1ry9XxDJNdsEx72k7k9wAPSrG8YJ
Hzr+hG2Bs1oW+LqtacImAs+mzl+w6a4F4teXk08r5F/sxubHYq/Y3+8/+/EA
7ygO/2LeMJeJbznDFfOXN4zYrfaSviaFTLXvHCeVRonv+2eQPuJ7BqLKUlRx
gJfgaa9JfvODp1Bmh+2vVqHkwWESZIyKuXS9L1x2U+g6qZ5AIgXAUHa9ww/5
tAHlIH+MGQ4gmQw7Q8waeOQPHZRIgswZmN6HspMm2QcSXK0digfNrjsMjRJB
1Jn9+wWT/9XRVicEitcJpGQyRz2xeXr9UvRpaBlNKPh9Iiy1oPi5kHu77sFQ
4z0Z0kWKefExndd8I5pNG5SJKQANwEhqzGll81DuwKcbdijQ9uw2Z34tGJPf
uzvuHm6cPRi65s+UD4fhnalPcbEC8n78XObkFYGyM+NNWagxw+2f0b8Zy3Io
MNgGlpqPjIcnETdlmNVTxwd0uHtBDBi3QlZVeAakT0VJHdCPLLP8Fz6zvsc+
rWzBlEUBWpVPT0zlqgbnu8925+b17IAop38WaEal0GRCxNeyzU/jFp2NmGZa
XtZ2nIwk6I10FL+KuVzgTHJCwyW/D5f3UWSAJBkgXn6+snVGuPSBTU9cj8cQ
1PKSsBtDu1gq7w4pe1dQfc2YmHX28ufHbZM7gRlQBOcxQRoE6SYkv3zYluIJ
dTE26z5hTYvlgx2eQZdNpuktHG6CTq+MI5nlBktOHI1kBLE1p/n0mK+3kVWx
Uj2FMNCoDW3wMm+Pij9bOC6HU7TrPk7K8B3eYJ0WC0Jk9J+Zi64MDT7Hqofj
yKTB2Wi4qBtt9l9bZJPzZlRTkvqM9veG5DK3Gv+EjACg6IzVA2ljMmuKo7TD
l4UQkvDC4RCNWmAF5fOzqGiBsrkQ2TrCak1Zk+s6mGTzrjdcOZvZXDSGkPvK
vySkm3Fpbi6GA1/cCP5nqGgZkrw/ognjaq9G7nrY69PECsKwKdTMa9WAwxGU
g+BJ5S8ylF1JT4cYO2Y5u3MHxsEZNCDEiS8FSrccsMx7BlHs7Xh+C38VCaB4
sq6nM081GBNibJgIpbyp/blAZ8+O7pOOC5aqr38L13rSIeJpGshdr3/E95eQ
Ygc3Yj6cwX5O/QVV474dizMPm2XahSUQtBCzdXbYLwVI7HCjLy2DaarNMvxi
XesTA8/6fKEkF3BgH04qeB5hzSqUDDfMBJmK3aj89qKxRFLCAX8GbOkBDq5U
ZZrFhMHoJhNeUDPn2cle2k5pa1K4jtY41NkMwYVQy2yj7rzHn8MtLs+/Adbc
sgRt2Pi58iupvVf5Ca8cNDn0WTMUgofo+aGCJ2JaXxVf59MXv+4pUyOWf482
9aEpIGJ0hExFKRUYfDmapjaaHqfOetqGThcGPSNRAR3BsF/3Rffd6V0aa9Fw
FyeLamsCF0La4QhnxzyqCOeJ7dOOXxP5uyKy0fHs1eg8qB+291YstC9JDaQ4
h/BD/PjArRahgbZnUkHFBj1X0C/juHpfGTZ1SvA1KHrbhaWNoTri3Pi76ltH
v0C7//aTDbW8RpHI4kScDMDWvVOlbIaQOWR/hD9krhjhfUlyETtCT01jO/nI
cIbTiYFDCMlaXgTabOCSkR8u/BBXyVE36dR09doFUhVf8hCO04I+ipcZaKfT
ALFgz+YQiVbkK58xY/iHp38mrlNTKQvgG22pJUvSWOEHO0nMpnw32mIsQUse
Ae/fp7FoQ/m816yoaHf/SRDjczZ8OmUEc23LI8/ZJeR9zgsLzchhoyTTGPir
ZLi+DKylv0J8b1mhCFzbEnRlTO9jaTAaf5K0Vf1N9Zri4d87OPtcNRl9PjfP
7mQApzqC1C5pFIQTR0Lj5QqPWc1y6+tHNsCg0Tw6HFB3/y1GtUxojCJv7NQ+
CvZIpflNH0j3umanOd0PdK+jLzOkxydU8RJwOywzpYICLak4HgzOiqG8YHni
j27u5kWf7MIc0EKHc+m+bn64jUbt1rn9c6KoTthNVxpsny0s5/m2sm5gTk0M
WHxFSlMzVLsX2r5WXEB0QZlPz+zZuPQTZq60faQxuQ67tUv/7dz0X5oVqdIT
03+abC7/tmADwp342Tv/+W2bPc14Ev8MuAaUq5q9j1492BrVXWKf/VUYh6dq
uVywZ5LbfpAL5haUWyemCMBdHFgSTfT8zL/9DE+CfqwL8KNbhHR4DQbr1nms
OedkVvkqtU7tCf/jWvK6sgRZwlGVyw9FNyuHsrjKihJSERo1Kfw6TvDrjirK
J3sdchLJfhzLo5se3hATuP/ANWfT6fVHypOtsRftRkZXYkUu9YY6odACWnQ5
/gXaaC5o9+0nuya+Lpk+Na6la068eD4w9N/0OBPYssyCUCrVjjOLZPfDoXhF
1p/bynKih+v0vq4FUtXUTVrXolmkWzXkX0eGc7wmUAmY4FnW23fLmrJWXD37
q4D2nWM5RBCve8ELI8uadPZ9LOY8KK/SBt6sG2EmdrqUJtWKl9iOZRVuneSt
KOJtYsAPsFaDYdyvTnd9x22auOhEij32wxJgcjx4EQVFFHVLjC5FrK6isL/m
vZIHFIW6Uekh0JcalU1ku0vVbI3RL+tBxQSv0xADjL/ms66HaZdgU03J6i7Q
4oArfC8wDPxY+/UqUltd02kgROA+kmCCTpA1CVVvFF/tcqbGFhCcAuXPPyrY
DDz+3cXXGtgys1TMfckRnqQ0V9V16nns+ucjWkq2vV9gECQ/6jDJdrC6oY/Q
4rRCu0BbXqnohSpiiJIf8Bd+9T01xNPepz1nwbChR9sSPgZgrVsHHL9oEhoF
EFBO54w4uG5+EEg+Xnane3QzpMgav6DGH0UgNXlcmUEkJ8WkiyUev6qhcxCB
ppmSrdLQHt8SlNfzQFHMwnsv6jFSWnMr3kITqfO9AcPAU3io8SD2tqb5mi2J
ek1QQHlUTOFkQOSKqdYtDE2J7lkPDyNhl2ic95Xr0voMYaE8swG/50tMmxyn
BWm3v+Vzk62uG7q5Uvnp6DmHl9K3vRrGs3rMHd+a986CPVcODOIqHOCpMj2+
E9R4BqOXGfY/YkVdk3oiKLdiCZcmgaLhEB+TcHf+g/f56JsAq33pNYkRN+Fm
1q9Vy+7NL6mBr3FEM40hFobOO1QS+WQL/GJwMaCMA2Eg2yFuGrbYt7woOgL5
5wuUb23I2Nx/ZjRVPgX7pOThKqSUr2pdvd9c5qOUtRE712x/VQjvXXRaYs3v
qoZSBiH3bI3xzS0cnoYieC/rS+ktm50nH13xn3qg1EL6T0fcfgXpLMp7Q2iw
uN6Yyun9OtY4/Q/fKC1yzutCdb+1FvLKS9vKnM0bKzeaQfiVbjsMTL+/91JH
QYOr3+wxDICoSh/zP86uzUjqpCpLrHqtn0k096nCLdXTdcMGJhF0LN4ucBh9
9WPLU2xEJfitFvYlQJhUUuuWG6fX0m6/yVb8Tx7zx7gTlhJ7asBoPtrZOm5r
WAN4uCQ5V4e3xwJC+7xtzPyp171Xe3XGF0lpTfvC/1AAYu/WAjt43OU1Jttx
Es94PygBlUvDJUCAWFAI5UlRXWYQbCjF+KHBaBy5IeANJGWFWBoQhHHxnou4
6cBEoIThxpjwsWIXXSK7P8iFpmFCrPE+rCNqOokskMSPXWlGNL4UK3N6Q1nJ
eIqGT5fm9deDGmnTfvj8ez8epONnQwGeRcIkoKJqqC8kiPRkYIuO4qASKl5U
6DmBhDPXO0ELKK3nlTYk2AqUNFruSEwJhsOB0Bbgy7c4q7ALsu9WCiuvAu1v
PP1EFx/L8doSHnK8VYsm/S9C5vXEgNIcMLqtKfETtm3Q65ieKUUrU9WFn8n+
NN/zMDDPfAKbGkYhNlIM42DUpsGyTni+CUKPT8uul/2mqDN9unnBks4tij2y
iKG1ND8afF4gHaB94Y28XDSxnmZwq33IXbrEJN85q45kzv6pHgHTKAIR1BnB
2FTGrj8hr58U7CMKBtWzTgN6GRN2sKzlEe/mf2AEVZaoFSiMxiiYz9Wp4asH
rGdHxy5Ecav+gUCyToeWskp1WMTz95SneSRIc2jmLScT42fObXZ3QLgP+1o1
vRcxJ2KYr7yl6LBmU3QCkMnkHzA1gXaAfyGg1hwYknR7Kj44QMwE9eUGBRG9
xToPJxoVwEDdM3xQ7QrHQUi0b3WU0pAgna5kXEtMe32EqXgZORgsqwWbR7j0
9u0OozPyS33+UMWU60+1U0sLeqlhXNpGcUEOgFQYJ445XDdZbnr8cLBXaYbl
n3v/c1BtWpvU4lJsw6EFosysx8tDIrVXwYYwxrg5GGvYi1POnPdXlALpSoyQ
i6PO8GI17bU7KXl/WPvpSzTgiNZ/nkAbF2pq9iNhWZ4tLzRaGmUbHFnT+nSZ
1rt64lnRNKJNBZpyxFZ3Um+du8RFnlVTehy1g/l7Ydaa+u49Xdj6U78qvLIf
+ztimBHHR4sR1/XiTPvdHRovr7H4IyTS7rVPRiwjaVaoCAqC8C1J4JBg4aF+
cAKvvWxRaQwJznJZzfDyuflEkOkqmiOvDPD+v++icoeERJeksDJEnMSiuTUI
hmzDHQ3apBtFmJMWZvQfiQK+GqjFb9ZMsj2pzNVS6i7hZsgWyKXCXu8RxozP
JSRDPpxtkhi1lFY93hQRrv/46BrSmLXPWE7fo8lYrUOox7bL1kbIqq1CNW9T
dsUToayUOqSpsjZiXXmHE25ayAJRMXaZJ3s03ZZCXdKGjgHODA9Pt/8bx4KA
HcQI6zUMj/tYsDRO0/ft1M/8N1m1HR3anU8QYqImtbRnXjTzP9B3VhELzy0m
sUFkTpVzciQDt6EYjGk7IdxpLJwicWhR3j1fNNI5Oi0Ce234cygUlmgIT0ZF
WEJHy44qkQruFjKOwK/BeQjN3FkwbyYe/c4/21+Ku30b45X9v9HdUDGzlfKp
SaQO8TviqtATC0w5UoVvaWYCG5b9Fusad6s1fv0kub7Czjhz4AVYWanigf6h
opNHoSP8vb4oV7eo8srwkW4sSj5R1gJoBguu6NTXaVuP2gM5/XJTzTAoXdFd
4itN9RYHNx1OIqqC+uIqYtNYz8pQZA2XFiq3jFFNJfrKmvT5QG06GTchWfg5
ThPkheWb0/VshhiYuj+dmOufmV3ws3ByGG77/UGNbq8WotMhswQu+6mGCcZS
JXiT/lY8GV00Iqmvqc0MYvaYBl+i/LFPN5pdGIERg59S6XYfefJpt/lTKSy7
EgBTm9XCuli97YWzriX2bSY788weGvhT6rby9kiZf/MiIPIKgRJnzCcBkGFf
ygX/eIuRcnRIX5Ag3deUNxCHTorEVkAguXzAT95qjq0JLZaXv1ycEqBTrsOX
xLJBqo8fI/Yxe4tRf15GZdkMMP0s8CkaYLOvg9CghkYltbWKQRpym1fi0fm1
/CFbXCz+f0fcgUhy5kwiiaJpf9CZB7bZX3NoZMTXQESG2hdVRO5+5N7RegxV
r1XSGT1vyubzBA9DvbvOvYWDshiGtFB630bJPHStNHXAQNmA4UtIqFajSuqZ
mPswMjaVnTcn/FpR6tc53PNzcjbc/h4wQZwOBKptA+zHmatPgBgjAxPRi2Pq
k62SJfwCoB9eFkPfU/VE7GcFhwrfE4kNkcFiYN34OVuvUZzf+PtwMI+mOVFi
SeettwTtgwJhlxQMkrh3KcmkxSEjxq6BibxeWaoAkG9s71r+s2pVExiA4pkc
dS3IP+Mk2bzZOE9NwkZG1MHS2wUTHfsDiXZkLROTKmoAiDpymolhUQ7+DSoD
i5ORoibVi/0k8McBecb0GcyJpjCMm0sd7FqrFEskwYJMs/dAEJW5dLOUHrkr
NFdZarHhcda9iMpHCgaS97YYQI2i55/fQ3fIon9c8nGxvs7Cm2WUNPlY0sBg
HxgQKg5PwKaWY0acWeiy7J+xbqk0+nLHywSG8i7R+f1MR0T4EW3YeuyrwAS7
wURcHNdTtOGlCAwJyskP7wWCLocn7RCvIAInkvbcS+XDDk3Nohc5k9d9KCqk
l5lz5hkIYj5qs3KlnzDB/A9ehOuSapzN1X8XO7/wUZ+z30fNkVzZHD24P+7t
G7qkC/92LTJQ15BXxXyh9fiRDocl25PLFHe2DfS25hLZThOigdSzfBVOeiEm
tXGftzEAB+3HXHV8g7uWrY4CXPuw7myq+pCI5/RuJgqbGIw31rcRUMWDB4OI
WQxW8uZvibdDkWC+f98CTWWoTjTKhJEsIfKLULZy8Jo8agLp1VHos75vWA5d
ptve2y3hRIqmfqf7PnTOLfA9onAXId4i9XqPN33SwD4Tf4ukOLDM6KFMm4Bn
TUNgHoDdJJfOdiEN3AGOGE7OertKs3omH7d5c2cL1MluzAMcVyesGqiLPdXn
wr1gnnjR/qM6omnui8z5cTGQWrii+E6+HEGzww2AFCg8LkuG9BhbYNlHaFE0
S22Z4268lx6NttsVjb3xDleA3sCatPM8sN0Qq3LoSNB8dayJe42UqEi9fH0b
e6cQhGNe0W41s1BAJX32NLn5HRGM2emevUZvD8iOitZDVNhg5JilVoFTZdB9
U5NneylHAknM9y3hXP7hgwN/JtFGKaDYok1qjyhnaaRJu4pHzbdCAQN9jufP
zgicAJ4tTGCVC6TF2nvfSwkaq9oJkEine1ubDK8D/dJtEIYfolKVJCs24f4l
p6B9NJGVtqbAJ+cKJaXAeMkBF7bPUvtdH6rH6hKUEhZNK8XY9qLgMoRXeKQH
iT3bydw9PFjW9LeLGBoHv3/AHByVi/iCmkXCjFytEVPbPh6AEnZlJOwPBKhx
HocPaYCLxWzXFFv/KGQunRu265VY6OpM260q65uPgBMNDjCUxVdK19zhseVw
5d84L5cuTbBaaCXtUCnqf1xVAFKjvlALXwszfjJ2LLb/hOQ2W7Dca2DaApKJ
sdB7TqLLRZJJyaKYs+t5At3BLQUtLdjQdpsJAayuZnIDWlaupV9G8OkgPdVV
zbzwSsRNkM0bo37PNXXisNvza2NWpqCgXBhOkyEN0mKy6U7/Em8rAtP1Fxt+
0F8Mn7y4SjlqyeWzlV8Z8wnsOFQumj3pM851URNZ88WjRT9iGypHSZ3uxdnR
UO9ZYvAW+wVZ2lqZyfCND3hq9muXq7Xi1TbqnTOs56qHZVCQm4e9P1B9osrf
bDwUBN7iMgTSvcVgc4quhEMIFNvFCTcArH3uSHjz1h7jdYnKMQ04c+Y7ENoc
e+eYKAVmMHjS0R3dEbfVjh59AINxl8dwcmVawrG63lnsizDLn1lyp6gtQjDG
jL7kuyS6cyCtHB2n8oLF0PGvy5S+At4ipkbgJIlkO+zouCjxOlE8hzZXTY1J
455cz010t+hsoz9+NEGqQ/6O88SwQ9hQQnKeOVRROyLKRXldV3rDkmHYs0YL
ZYM+RBjcYEK7KqBroEvlPVRoC3kwc8kWOFXfZ5quQIb/Fjl1ftp78ocnfWRf
ahwXFrjg1/vcNMJUhFQXcAubniPRrgTpF9aZkF4G9o4gRsxGmrzziJXthwwc
n008XSKzOO8Gq2XTpLYcRcp6Af0AndTsSiv7pIep9pBc/jKmih1oM0OKo4zj
C57gXA7TGET9DM1rm3AkB1RM0P4TAK0QAbB9TqgMI+meSQizrIXv7sifUQHx
rKd2zR1YsoKqNsVM7G5qS4H69pC44Fn/2SDqTCTZmhnzpPtaWDPGYwhwgfq+
MwptbhYFY4KaAWxGofLslhSDMEZnpmUZh7C6R981jtEaHHWCR1gFI7tYpVQd
85AJRGh1Q2aJesc85o21ijXjytsRg/Oa43vp+QByHT3iITC9IlvLUUcG8fmq
FNszyESYdXOpgqduiV8y7jOXmBpNXyR+vz8bJcbhYUK57aQ4AKLc45nVoV+k
Lp1sGMsN8wEBrM/02PaduwmWWeIyh5DyZawLHzYkkL6lGbhp2spn/nwIkzWl
q0pEG/u0CFTm5odK6WC0s713TYzo9tmOsh7rS4DDDOYEm+TF/UDEe5jbI4On
LUi879mMKV/5yzZKjMlUvhoYXi2Cdjf1jF1WBfX6w9VFexzwhK0Yh0Zfj6P9
qXo5uIt4s1mFI1YhfpBPx7cMfTqTY4UYjvJibhhppus+MQwkSRtzKfpiAMYH
uEyDVK4jZBnSg2QEp2qsTyTP5U5i69uaR3969wuQ1JrVEjDQDq10vEHToG2I
w8F79bAB4aU3VaczeTOdoTOFwdBIa+EncYjsbCJhoNFYuXbvPNQfeyHFYHZk
NlCVD7DtQRu6CP7KCqp6PfTwpeLLv0iQh6qd1MUFXGnUZI5KNMtYXEuTCV4q
jLWvbeT1S5az0yJQcQE91SCQ9sV5v23wAOiGkcbUz1TNOzzy15LiT5Pcfjdq
lM9eUI/LHdymCPVAUPQec9Wz7ZWJ83bY0uL2295VV/4iZs8h+cudil8mK0Wg
cRFS2NDsNt5NYF40vUerWDP6/x3T6OLFOCwzI9e8IG6vEU5k2si5Gzlz22Lz
87tQMGe6FTNk5CVThVhlBcTGUq5+Yo5yztbjw+9nBC45O7IkBU8WdHmQUli5
rC4wbQLl+8FJ2ZyFY5t0xbpc18Z8CX6jXHx89uH19U+bycRdKdTVJABI8DVQ
nyM+setkck0aN7khytvL7StxdGJLn2EecHgR8RDhT2RBJSd/bjCbnfAgaJ3+
Lt8KZmZTXGoqdPVTYUiRRmvgEWfYh018EmePgbFYZy07RRTlIWh2j1pUiGw/
9CyObBbHui4p0jx/n+vYPEf/HQsK1c5t6izW9A++Mk6QDFVGhCCdGhyIiiWy
rGLu11AwSMjWbwHr7UbtPQqoCPXKaqSoLLoLWK3vxWzFsvFbxIgz90+fZE2X
H+CGamf6NXcvIKwYk+0ml7+uAVxb3xc+Y+jJrpPlPw+Q7aIAv2fPBzpYL2xP
hSl3Tl1IYq9F4DB1fZ/8vMCkfn+MhStxpRXYDVx/8vFKuaAGrFbEGSULvuDC
UrDTUMQWViThQDd4dFtU40fM+5lZRwMtCy3y+xzoDyioTgUQTTr+wWeKz5Jp
eGzVZZIAD8WL/bp1e9PfFs4aLkzCQBuBz/hgdpyjhSjpJdvZmYH2eVk+kl4V
SRbzy/mKNDGHGBGs+M88fjUN0KcLfzHOvzP5PWjWMjSuxTxbyPLEylyz8A7n
5+CRUHk66/tURz0LnB6UxXKIsIKSwPrR4ra/u8SF9lnus11xhLm8E+dS8vmf
RQnb+18uuSrVzMvNMitNQEkFJbjtJo+L+UM7IYoRT6xeI+EBg+nHdNKCOF8u
/PMgsa5YPvlCYIX208DIBRbWeh1eViwEVLTMnPSHuQgrUlyo+pafr5/posfq
J2mCvsmrci7zaXA/a6ycMGINqBq8p74A4m5mX3xIooW/RVwfuMst9XaqqPGC
QMwVAaDNgR3DKP0uiOpb8XoBriJhaT6DLt/IQo9qG5iXRZyc5uXBZFTdKVnX
PTBYE6JpkakqCctXvHo/ZWORLlT4oQaFYnGD2vZUfBHX3MGtsxv0nScPIDsV
jzf4JfM/zfetnIi/ca3xedRlK6q/sflvgAOIyVVZfXUdqJAMZHOWQJLR9Ors
PzEfx18GQtJtvEMBUyxLe4gVf7Ghv9jlruXku8BOWouVBNXED7rTiQgh4dHE
R+gyh2dvjOL8s78QZdoMfl6fM32uT8rjyQTRXItFQWFpXrRzJ7GOUdPB9YFL
FxWnQ2W8ZQs2FxaS50CNRfgiWmG8LaNiVOg2O/IIpcGUs9EQ7sJuVnW334zo
2ugorl+QeiMcJ7owSDzzyLLivcBA0QAPi8wX2pD0sZXCRdR2eo2rjs3JYqib
aAD4hvGP3YacJBaZVnhG4sq3ZAGnJsAPk25gHZmyyGHpLG3W7qz3OK/eYfss
w6OQW58vFm5Tdesb0JfoL4efYxRL8F/OnzM6Wk0NcyPu1b0wYxjC9cxhyM46
t59U+SGhpCLwA5iTk4X+FO1SWurD0VsBBtaqkNxALpCcsx+Q21k1EHpa/G+p
Oru59YALpLcimq6EpIg+l5/d3xsOd12VGwqJrxsR0zsHRK5Wrmky3MYFzZLo
TirxEhrszhPXzFGSkQWQIE912q6WI2L40UeRRBtwDAhLZogwpSFo4ObyLEJK
svizh8Tc2Yp/z6p1cSip36wKr9Ur6dmIOvObej3oUHNIbfjyZr6P8do6xIQ3
RKS2ntdFuUqtMRU4QWhhGKsYVmbt7h6RM1SUG8+SqdgRlf16n5AbTlG0AILl
8OTb1BEXIzkTuNaM85BqeX0Etz4hYvGlT9bCcq4foH0rR0cUwJLlhLuXvXMD
X6BMwIrRDDTo2Q1cDMvbzwdJzhTVRyFxyfcIRWyQxZc/igViE+UVNfkiUK6f
dBLwv2MynXkopU6d6Ekqsc+FbDvpSUTXgMPUnhdRaAtLtOVUL6AYiOw989Hw
YaUs8xnj7CKbvc4UORzRkOBYzMOYmmO00fJJmu6qzj1eoZuLfG9yPnz4NAQC
FlFfImNiYt+Diue4pcEh9G65F8DDXlzFmZOzyjnpr+vxKN3e0NWct4icPXrU
syQ4TSDJydQtbMi9DvvkkCUvOsZkovgSzWfA8AA9MtA/uxCIHbij0bfVCkIo
Re6l3gB+COolJ36zabuvdEpj6BUqMwOPY7QjkAWRiBjHoZoMI3Stg3yQFqeC
mQnPh53pGwsDEVX7INLrjAU8xRJR2CXiKX7/Vwu7q/sWApOqhnxMtRdBrI4A
//oipQddfrwZEXC3U2xOcjjTvdpIksiwsbydRF0U4TmUIuESib1ckRs0xMJQ
5jZ6+XLzvd/2HO4dkK7MKSXnXbBjQBvkxnLkL5SSYO1/vpQ72yGfu/bcz3vN
KgglMobt/Ly9mgspVu8tdX4ElAj6kK6skRvbooJS4ytX2mZrEBXFgx3L4+0d
vpM2Y+y49vFhjvoEIXrxqvd3v3C2EpbtUdURvWMGUPN4ijDWtQa2quSjxENj
I39gBvIRbSIxSMD3EABXRsNOVTIeCh5Ke4jz7sf/Pv0qjLMqGI/bjgq1NfHP
juIi33Wqto3LYvf2M6rvmAoO8F0iM5tO4yNJhRR390Mwb660UfS3ib6Rx06g
f6tiR+vLD60mpAVmmOPYCiyuLMlQhJ18kTWLkuxJ45Ws8WPDWigHIDe5FkfM
jPbWK8hltOCNnObvaZqtDLz0d1pev1y++5iaAASlvDDdl36AbXj52k31ciVy
JkYrmVQMg/YxVPN5UINGU0p7knNMdt8aVIOUHY1sxY7gZU+a+cd4+j0WwGlS
11i2To+tIcJ71N6B3irSUC5HSLQzsnvrPeyVrMGrjYKn1M//nX01yUA15gwM
Imokpqh4w1I+CoxK6u/fyiz6/I0fBI8DglQBgWLTJs8OAN0XSvR47/Ks+ltU
+uDZp/lemJestUsqTLRCR2UVgTRv18Ya+1RUFYmp1dUR0WIIYPcAdkojufZy
J6YK7JeYkaLvkvXwxSuxSuJEcN++C59xWTwfhAHl1+gbfaoOyAKvg5vRPd5x
ppiFtTuD54etJGBfw/QnDyxMstmCHg3MktQ41V72Y026tmnlRCEPU32+5WVf
YOVLx4DpEhh7CledWe4zpCMjXZTrJsX4yU+W/mYtnXebbjU9GfEzg33inseJ
+IC+aHLvR604ShzxjgcaClxPhQFo+5PYC0FOnjHCi5ioeWJOSMSN5HDvE15V
HvZ1fzvwBJ6IG3yE0aIEbhMhu1QX2XRoYMOl7MxWoRJxXhsyCZwEyca6RDzw
b68u9NjfEHN29H3uza2AgJNDs5rvmA97wboly8HP0moXy0RxdnU35DGuRqX8
pF3oOaM+9tTQoyzXozHf+O8MuEWibnNNZLs5mAb0W35ijvKpWofvoXxeyM7G
k/C3/rt0yaQJFwdUwpZEqON1gemR6GPonhgXOmTth3yQUgfJhiLcUjSaNk3z
pcbTd5nFshkLLWLisrVRytG536CaiUqWWzYk3z4G8L3YUdyLOK04c1sh6YD2
ly6PcBqnrAGgSPBo/DHMxIbIriXNytoVKEdHWVdDjJYlGeMq3bx3u0gdry5Q
I0hMkicUBvm3+rcuwDqeAPVQxJmevktNJjZk/IgS6p2vtuX/B/LWRzaFSfpg
55t5Er7n/IeeOaQPCaXaWCpqSnIh+ArresJyjgxnCNdw3b0MzO4SvHvqmMvI
KPO+N+pnQldNIBVYJa2cixdPbDKKngUl4MI/Del1Dy+fz0le0iRemLGcoTSR
z2cjssUhM2X1r0Lv9wveM9KNMeUYBSEcGoERWwv2lLMU8u3hJP0WIgpt3uxC
x7+p7FXC7TLASy+OrohUoPhc16epEBZLO+vOk77d+9ngslCBfw0fXtZzlfhA
R5JxkcU+2bsFSufM3W7Gkw40x2zq1CuJo3IysIXrkxTTTMhH6opBAoTR6Z6p
0hQE/RVFAije/gVbBwBEPGxOFIEyBr4++oweuYkdRFJwd8W/jja7tfQihIxq
C04I70IyU7c+U+OKewGpf2PGwa5uECRMs35ya8VZrWeJc9IrxeNekgjw80ku
g4WpQHQKkltMFV+abRSlLrqYbRj1/KMmmdzNQJ8/gnTucBSdSgwkqSMvwvre
kCfeNL0d7hAR+xq2FV5Mg2oT/tCTIBMKgho63jx8xHemJbM2a8772m/xH+VJ
NQx2zCv2LVTKXc4/qnAsz9aGtVRH2v+6PGnZnawedQxDE5bTWC+fjwZ1ztqc
AJrDHHTdNIQC/tPkkTFTCZ8nRLEEYDZykVrgj7zwqYZGdM/3fMBVdm2oXvaB
+GjO338dCc3fivCTK8dSblqZz62T2Dhhfy65gw22So4QOfDDosZH59EUlrdh
poRqUYHyICJAzUnEcjHZIGYLlhubqNrWOppxaDfkzPkoupVTFTq8CspBMxnw
0SqcboEEGqI+gLYO3GGJ3xCV9ezWbU/0QVCBQZwmxfFmVMuYz5YYIfTf8iK8
KCAXRC7AYBEBlsioxD5TqJgKrN31oBv99Bs+zKV3KDstjNc2xlMEzFKKqVWn
rhqa84HYejqo3KboCqRbvPAcN3amsh3ujkBHtuWzebGPCUM2HgGK9RDBtxbP
bwaEV81La+VnKhqCCOrXRTj1DedM3A7rYuGp6fYq/l7v+JgFxF6CQcmnDJwo
Fq5PCQ/oFbZm7uw7Xd+Lz0lLuRsW7QBig14929D5hxgoRFtNsnW0574Bh7xT
WMjEDJHXHs/7TCxn0DKxq63CWiD62a5rt57UNxgvrZrJlHyj4vpkgxtcuGHz
qxOvwnPuKskfYbnODNwM6nTmfZuWs5abEn1nsHW6JNTNz+gN9Jlc767HAeHB
3WnRK3btnUdxbPtsUc6LljkklJzlh6GKErePWz/RC/k5wwyHSF+XuBpjuzW9
tuFLJkShErYyDichoLdDdrdWnr6ywgb4AGG4CAaw6pj91JUPiWXLdundl+Dj
D2XEN4lHk9MFR/7aQhYnoDf7skGutvR8IxyFFj8HUlyZj754O/PyTJ5fGxS+
Q0JgaEyd0dyrmAvSaON7vbxlgTRSuS8rLrqCvDX8+5sTXwM5ECcMyee0eAOw
x6xugNkR2Wg59xR21SocC3NYii7D4L1O7zV/2CPqGn11D0JUWLC0KFz0jU10
UdUGsxrwm6WqwbxF1Q+IDAUZHzoNYKgILfLUfky+xik4jdKVG0dVB+0Qnlsn
cCicXigDRF5vYzL5+llMSbHPMif6EU3z6a2NbPwm7xbShZ4qZ5CA4FNF3p+2
R3muDsLlA88dR1X0/HPxT5CQo2uLU7AVitz8z9CL047walQ4pDFrYo4ZFu2w
f+MCLrUag23xwc7WNo4weEEAcOs6HMZu8qTy5j582h9BW8Q4QWmGuFu9Qdx3
iK3FOlGRgC5GHMiHX1M8vXTW8vYi4a717TG1vX8vivSJwnBMt8hjz7Z4QnK5
sotHG9+LIScD/R6tmlzj1QsMfm9Awc6K8tCeVUFjeimtaBRBrlsnb8gbze5K
kKm1Ff1iw1D1pH6gdXlV8ey28BBtxBIiREpYwiLmJoiYkI/1JNhYXvSIvgYO
GUmuBrI0P6qiDLWtkpToPW+t9TA9a+9x5k+IGUh/OOjTDr/1/usLEcGRUvOr
vvs1vJlFE2xrbZSI5nwTIc3XfUVAl9QkVtNHMYH9wlq6NTuhWvBfWfPr3s12
DMtpXFfaMM8RyE00EZH6kR7OvSTGYmoXeg22CA98JCjLf+uOJxMQVpTVWcUk
9YuG/E0kLHQrjKJ5J/qLpYDcrzGj03Pqt7famq94YDyffjINcGu8tvcfuzFP
zgOJs4TaW6BkTgCWq9U3oMG2qXblxANei67cMAkw41alO+ZLFVmJlX17g63g
/LZH3Dlz+HuPwdKk+f9lUU1LLpj4lC5Pf4r3RJ9mZ6kaGmI17pK2UhtXMaq1
P3CGcZY1QGYwFis4CycgxxgpCoKZi/zvGAXpXikDLi1dL0zE4tkKmONouTC+
lem7P8boLEuOaXi0xi/25tqwH/dGebcByzf3cB7nP+0z2+J7jIAktLAldfC8
8BErBx+44c4BrjbtBz9GdbaVDgFc0465i43JJ15UDq4GSCL8pQ6EKImKKIih
ZifpbrRYEmYcN8zPkr2KGPTNmg8FdaFNbTN7bVSMRU5o+9sLH2DJ5ey/Ob9i
18GlscFze0U3RSjwrlt/7mV18/n3t0+FAr0Woc+B7USTnl9AL1nlTcB8r1kZ
vcfjbWCQ5zAxSANQUZY4ZyXsW6o0FPe38vUUR5YCtXk3siuYbci8pCgdeOov
yQFdieYkhjXppVslTYgCIoqSyfoUr6qW+NbG+PGFOW7KhAxR2o1bwxZ00EJA
5A2WXaP+xlYWu0+LeKXSTbDD2OrkZ4BBQITiXU77hU8YcpztRtG7R31qG8SI
vstybESfpPMheCRWnwZna3vza85lvJnA7+pDBu6RI9RYDb+KrrVgV9zJ5uVf
GHVF1yu8kyi8HxV8GHfZIRBMg0RUfBkqXS0yuTRvdRpEEaSsL2Q5GMrxPuF4
I2XuHisG4SSJuaw0lroHrQCSxPYv+5jVVpklP9Xxoe3TBh81RWWfw+A4AF8w
z6CPPLpjbEdVRKWrwRVt3LgwQER3bCLkvpVzwmdvHBn4JsFop3CQpvoWmuvn
3+WbARpoUMNQrZttyrVmc8uNz8mYonDoraeeoJSNCOVNICkA0+jXAcZcSkmg
07oHBGESyPAqeQCWEO6i19L4RTMg4tPUYpWysIWiM+1px8fTXb8uE3vJlvFP
QwIhgrd+64KrT2g2jNiwvitxJJ+k2RXzMuJYGpOE0fK6xeCa31JuzOVMHYt+
cIcFWht9FiRpBQlAghRG+048X/+To6J7wlYZSdxemADOr81fMe+tw3pq8kWI
tBKJsDAf/WkF21sx8OTXoCRv5wTfweFK1bnJ0lz7WbBEh3DXza03Or/PTQQu
cdNUaoAdEr1TG48KUcM34w0qTopJrvDJJmWI5N98FNY7WBwX6Ph0AvvqqcIm
SUBncJc+dn2ixfvl2dnn4l7XFNXuXQ19sLS7p3uCZY62TgeWwdpXEKe9t851
VlijdMO3z8IADcDUIMg8ZxdzmMjyrqmgzd/+2moQNgBW6f5WQwkbms8I6x01
5ftQUfY7nF8uq+OJtjP/SRr/h+a17QgON1+9zqD0RIRoFDdrWUduX67cyFx+
MF1aikGTaucmR9EI5pUmkssPd39FuDBQu5JC64a4hBBPDOF4yHNa2scaPGdt
Ii2IjxfaJlhYzdBjCL32yugc4sn52hz14dkmPPfGDC3+MOtKic8JkJEvKYuS
IEGqp0LqpdJDbfNc6fI00gTmGwsFsq+6NwH33fBxDw2aT88Shak0nUVGnPjl
v2FHtI5nimTKr+NvwJhhaUPFsyS4d343Wl53e8Aau0qC86APJNG+gknRaqSa
VKR36FEAb4ptBB0CnVijRcXEwJEAzZPqfos8lCy0ypUloC6lb2bI/xaaP5Dx
thsBsYhJkaF+7RGT6+gNSX44C6FiOT+kHwupbXv/NLG+6sF8wfqBnHbGjM8n
edZ5oeUhO8JwE7SMn5qZH3ulHw1xLq5lCas/M4BUWwowAw1woxcvW7OyvVGj
zO991VxQVqM/G4haa+3g95JmhlzDOkWb+/eoBGiFCZ2uPV4Lyxa7PK1uR40/
GNr/Pwbb9tkbPznVEKtEMM/KC+LxKNl8cGHQh4GWoZ0xEmjw9x57in3FTd1e
0wdIYX1s8baY54+F1o4neerRNRLzP/nEk1wfpWPqkKRgF/ORVfyAD2tRbDyO
a+KQs9ei/8b4pJQhKkV319qZcl9tmXfyUuQdqNAMns1rLTQ1shv4WkyBsoEf
66u6up7DL+i3cHLNEk8Y8kuAvUf6okh2KKE/pwtaYa4Dw4mQrmmowIu60nw2
Zy0A53ilY2BYXPELXOi5On308WnTZwkfOORt9d3aHhIdCb5285ZkoxqqtgBv
eOVF7IKmps+lC+hbmgBPgT0mvSjZj8lVm7bflBgrvz1XimvpVLO8KqIgqNyL
Vbdyw5/ByjhW8n/j40lkAzv4dIaOshhNkl1nIB86L3AEU9fwB1QkjbBtDdTO
2+02WW0SFXndEMPy4egmQeunBE2KExG+Mvl+7ADPwasl1G3VxasUQQnO23fp
kEn5b4bK0DutmF3k5O2KwykY+YbsEGDqBuY4fNAiiGtE8O2L4oChg2ca2/WW
nDfu6feZnPKeeeHFD/Gc0/UVPe3WIKM8uUpDJj7xevL+6SGdAAGk2QvlFsdX
nYa8KN3C2D+4dC6/Dp85kJiVF0tV3ixC9fHZ5H+xsCkaFap8j240vcEXVo0e
PmIXUGI1kYBcoH2FBBsmDAkwEjeHGl/27iiV0NPxtonAH77h07T4kv4MTyly
8DiusnPDs8ezsQJCTF20DJBpsmPziM08WpLFTIKg/uYS2dL3jHTRoYVr0ItD
uHiOiRJ1gVyixhJJQN/q/gBI+nI8YUJ3K5MeHysORIfr4quPKDJq+QsBUYNo
GfTKSoKf24YWGg+Bbix+FHwPBLzhMR/bW4JJACQAZiZNRmiO+nA+neLMdtbn
9NHCNVXUrRztRjO9FYKItU3olOI2WKLTDSL+4UhRcWhvgND2i3BpH7Ttja7O
iw9Y0OKm2dbL2QEq9C/zA1PllYOISHqMQJqcm4/0wjz2O2CFU0o/cCChGXMR
9yvLXILMmalvqM5rbTI/SCcYJ9nUqAQqmwD69lpMTYgiRhw4727kWcYyOX81
UDgUUjYFmDZ/qiaaFIk9R/klXRwfsucomUeKyYWSt4hqdDimLqxYxD4RciDU
KsK5Lvqzrx1hC6/mgafRRJrFl7y4kydsZ2hPFm0Wt9iXx4hl/RzCI0/v8OpS
ZH9ttLXJvjA77Exar8sBaaITjKH3JvNuXnPJjPiDDo1PN/EaGM2DdLzqUnnD
2fB97e4aFZtPdRm76YlIsCcvXjmT4Xkl4A6SvAk/VGVbVT/wywZA656YOGVC
vnbSLVhGrwawBzDvN2B93WyZD6cv6mTadEOtnIPtw8IGZ4RquUNbQT3cPcmj
6iiOdFmWV06emezvpF4vOAph6A3UkIl0GTsxuMuu91LNQ8giNDrfNYuxwFYZ
ho20vFpyss4fBXwbkB/jaXA4vqPva3MddAoDCpR4EGtXuxY1ZU3ntR0yXtuR
v0aDjAF/WVWS88oA23KquRZVLsCBBI7OZbIPfC0B4ot4eKkuG17sQlZQpPP4
Lb+2C/OYuawAlVo3ioRVYVf7HyKl9FHBHYDA8tWGkkWHBozkltuuqtMcCUWI
XPDcAJ+dX6MMSxtjeNle0WfsLLb+bm6LqOUKuwj5cQ1vQUs+AJKhdgW/JyRt
Hv4t6vYNruAvg9JCCWM5yzutBKKTFqHMAEIxYuBMvzesG3NJwuoelUGC4iEf
A+iVjw6Gnb5uoPXvj/TwB1U9fYzzZeesjDeBoOyWJv+pWvgUrh3eaByfqcsJ
9RuUL9AIEgCyn9XfQs0kzO+YOTb+Ku4kPoLwCL3dl70NZHB3OaGPUwbbjb/1
ezPg03fUj299X6TkDUiN1t7AofzfNErxXnk7jussdQB3xt7vRQefffIzZujj
pzk0fm+DTk1A3i7zSZ6gEqWDJt4a1Wj9l1c6hXXhxyApU+pwh6kWo+h9dYzk
i0m9X2kGf23RClVTuCokui8+BUrNQ4dkyrAh8ZBsJqUtOY3RXLb/oAbLAgh0
gWgW8hNCdR3bHIHutZCJhutwCL2o1Z22064/yQ79qljscMgTGGHB4jnbNYZI
Xjeccy/yyq1XIgaVClSuUZuslllbX3c23+jIrI0u6QxUrL3YIe8+P4FLJmKc
Yfk9HjqgMtEyNOvVC8yc97sGeE7Ztt8Xt5ON8cc4bcrHu4PI6aDxCTL6UQqd
UOflqruNLu8PLEdzw+m9kRrhmnzJC90vO64valkveR/Dn0yU18Njjp/mhJ9/
FhmiBoqKmZMzhdgnQjqEUjQE7F0aiTPo8LUKrf0/PgIaJhEUKEG9/feOtQHk
1rxZJz3ckdjVymGaTtDwYdJ4phnpVexGFXDDXLgofXzJz7MM84BkBhBY7dWM
0tysmxvr0ZAPukKOzb+pZKSc/N+DysDnvEI/FLEOaB37MAr1xdwH09FR5R2A
NoLEn7OueTOgI+92G+As2nwsUlLXJaGGUA2mh5MYd4XsANRioVzCEgq/OQwP
Wq4VZbYjiixQwQAy1znG2jgDWLbqWx/FF+OG9Y/AnYRQcHWDoBDbR6MWRmPp
MfHppwPlU0As/to5IpLmxE7Gchf+AHd4KVWtq0Z7AaiHJ1Tk9OhD0hr1SiW8
aR9LDD+QsA4deUC05B7FeTe4tF6z0ys2bHBbxitHSqAilptMYdTTvgmOktAE
NLtt1VakSeQ0uSzN8Pv+Vh+3+1JcJ8TGMpcGNX6eKiFkNQLfwk5paILtmLoV
Rej4dmt/mqlAptU5zJBP2D0EE2njSVydbhVcMSPYZn0PSKEozueLOGkwC+33
qaILjfFR5K2SjstK535EVVG8Oz7YyGvrWob0DoIDmlgz//T+l6iWWV4ltQZO
4NcamBj3WeQ/ouksxTvu59ZCFW8F7sKxvnpxjPGTebiueyRB1Az4WeuFjqu3
SYfhVwWpqWBXfh/bZ6uUk1ZAFeh+lJkWXqD3Ydl/opS1GfWybG257WnTIWP8
qUK5SCn5Ah5weq3wEa670Ms4ejtpJ8QpYX8W21SceyonDgPKvNXgvEeyDgtj
JmjDEjCzYv5TynaaOr5xUk0WedgILW1JzC9mLppUXBHi27K44Kly9sNQ93/h
pVtYRchx3c29PDZT0GDtqc6KGKzZbbsjkC3h7fzWRXR8qAuIM5wDCrl8Jvrc
/wYCSacHyqGq2tTuPUUurdQGJ+GevZO9mBZhT8Item+tkq/t+WXltERaLJ4c
x0rDJRPjDMcSJwouQGXWHoOTBnMIF4u6PTuVlalzXeFOMFQbB/6e2unv4LNJ
ID3v+dwOKB25vJ2Gp7dh4MqHE+Zyj4AFTdqjIYPUGa0IbzIz+LFQRMBNRMXb
qEmadVfU/pRIU7rQ0bm4xKobCnNy5Id/lSR2/NhoNebivPrcMyMp+VstFTFY
USV8epZVExY5yKPdhr0N3KpGwinB202ppLWlD4eBIZTExt5uDCv5ZAEW7AB2
Wedf0C/+Fm9bZjwLasAAD8gJvc0QVQ4YZELr+VWxVOOidHpyDcCdQSykg/QP
TXuGeG7iCeLWc+pl6dLsBGOno1MzneqD1hq+rQ41BkhuShCd7Z5hPwhsv0BE
2Jm0lUyosT+2SfogTBPN6+9JUuMe9N9hlbwfMH+IU1MneyHA5jxurvFIP0Lq
uBEbZHL42x3oG/hIneND99WCjuSz33neyQdNYWA0/9ZnKbMg2eglxP3VlMsS
g4Yo9VWwmQhihtwiSyfE7jK7MBpCEaA+yFQWGbCtL6DrRUKycDoJvf/z5qUa
GAJq5Akv65OhLgyaTcole5NsbDQovIgw293gCnAMed46wHBZ0Dogu12WzvCw
3qG+MDfoNLi26bdK6fNyK3b6nZ32pS8rohVbUtq5gnhtTHdLFZOLKakIrDS+
sIoMUvxeS1z7DvFFeYsFOAGInNOwjZYlh9vMK0e7Sv93qQsAxpGbrYA0setp
WURX5SjCopRCQmLEt5HJwTRt6akZnBU2DtD5uByUauNXYpBsoLrovPrVXaFw
rXnuqdBcbf4E+bBCt0nsxh3IYR9ymAVN/jk0GG2t3sIMRadZHsiW6HB0JavG
r69XSDwHEkLSY7sW894jxZwCCgrcENlCGqijg6GGuQpZIja9Qtixb5Ole/mh
jK8dkMrpWrOhdd0MTQncmSiBbFzNfuDl+rt0UyTjV20rdDBtC0iv7c4BhA3L
RRqNN3XMD8EIr5FP331Xw/tPIvb8cqv7kjRzZmuAuFTfqF2qqhjX78pm87Jv
H955sEGqiwzlByb+P+32cWYsYDslDnHbEoDA0JTRjk5XJzSpb7sPM+CeiR09
WmveP2bnp2Uu7mfR+WcMVC+bQEyQc8YngaqpEI/VPYWgmX2fSBh0bMQIY6sw
mzB0SZ7Kp2rOrmUBIV+y+5vBOvgccXjCnOhxcySuUdH3+Ol0pXPun8dAZH6B
XaUzSY3cPzsBga1Hr1dC1yGN3lEC3cRFhH6QJTZ3E2Vcd6G0ySe5IlrKGISH
7OW1prjFUvhIVUVhZCSG5EayrMYVO10IA7QBJ8kUas0eRwJ8lCnenyl670Ga
7ODyT6TetcFQ+1O0xfTJK4ngPaZMcK9kncld9PPRCOXNiJTgH4PHxjladR4S
/v/IrOGE3WcjMunCIduZfi6WQPgOFjbKkAf2M6VY79s8XBkbYrAeDUZR2cq7
ysQTudrilOh13E7OVnCPGODjvZJi9RBbXfoq871t3XvkEXcl0BrODPjDtkQz
zYs7IlxLM6iA0QElgwboWzqeWd/cB/nCGF8ZqqxzIwHPoBHwCOTWethLEdRc
Rr1NDZePcR2DBjMeoVBnveD+Cm3M6YTk3VEm9rU1OBTKs0E4hjyuJ48LXPwO
qt4gbQMAhgplqWV/YZOaJ1LTzKX0p2eH+o2qAddQ2eXwPiG0eSTzd2NpZSEp
3+g60BcufNAtvglNe622MhHUh5wVBqBOtQ7zhZJowkSI/JLwe2KvqknqkHZE
TMZg4xcgo4Rd+LOXSH8dXdXY7nPFcDsHlO8aQxsJpm/musDI37nsZPelvWIw
Zp9YUFmMz1lE67w3r7yfMJLW13w+N6YTp8PZr+9l+qA+ck4KEuWwd7ADfpBl
7P9zqwnniIuLntrT3wkgz/yCWlq09nLVbVw+HgXALy0FXMHTOehUFy+3LH6Y
UaLHz9etnL7LvwNI7GRjCsULU2Aalu8hJz1xyJQNABeVNex0VJ4wi76QRXKc
aVbDvjD1KT+27sy5jPfPskJdUiley10qLqYdhC2YTtrLcBdNxDnZbx7mJZRK
BQKj9scSZKtIqLkkVlIRDGFKxCGOWi4pWLO7lGUaEXpa1TxMzfN3NREAUyMi
J3CTJBOJ2HSZRZ6YsErMQw4XGk5WrXIVYF9Me3sWgOB6jS5VxMWrTjDPQFij
HvTQsrW1Q1KnYQ0qbSp9jA5SP6q6eKvdBYOOVfJn9VydsfqHSmu1YqCR8Cny
NkHGB+96qkmBmgvY47p4f2Doa7sEpEcMHlsBAlQB2yDCLeGdJ6YGdOQtQm/i
0Kk9ayKbN4Asy5ur5GPi7FautO1t3nBbWCqwIPpMzFxrGxRrSQV4v5zsOCEh
L9vM3bRQqaKvp7FMyvTTo5i4lyRnXhgPLfzn8eC688sC3zaCOTdUgzD9dWYp
SuUXKzBWoy3rgN2FbitjpBQNMQahTqXfHGgErUXvytLWD0ZqyRTLgmuuaZ/B
Moti/ilWAKbqQr7ApDkEOhu/Bjg1LF/JPQFn9p8Hk/DT/aK6npseJztFH5+1
Kb140VWBm+kfifYRjVEIN0c7gGE9G/TbXxxI2fEfKbexkrrxZ3T6whtE+OTt
k6xrG4zsVVqEIqWH04fatxyJItW9sYsekPW6imLr4an/uKDGWuTksDNTeXA+
WOmno+5Brg2FIJExNPelYUM9Xi7FtMa4QhR7/XTN+nvnveWfandEl1T5Akeh
AugTyLO1nCaeJ5UT6OMMtsi3dBp5I/jm3elOLrLyPwxrsq3VOcNtBWroQ90P
ErUSlIM928m1nC/mNFD0/wu3c+qBV3NKf4b1e09dbQbKXF3ThLL4SI/zs14g
A34dzeCZIHW9Gz3IRU0qbcNNlrXw2aLX/pPCSX+h9r6w3pSiqN6+7wEOzwBl
56akt87O8mHxxDnA4HYCnPUBb6VTQnhsd6n/4FOo9NghunVY0Oee7h8/ugpI
XQa7fkyrsvWQOoYECuJtnQUAGdqQ3KQ0oD2wkWKQW9UhiBIbSQFnRyLeJGyK
Cn9DNTSEjJf83kLYOV2oKVqJnADwrrMbOYGX7ZLpUyDeREAgGIiVlQmufM5U
rIo0QzVCsxSF//a0XfY4Jng5XkXJ8REeBCqD+4s5c5kHpgZ+JXuhS1mUS8U+
qgXFlVRUGOYhvcsMuzIQ+8+ZLOjCpHD8ChgDifiW8ZIILHGoRHaLxRbGEdTh
3rF40T9thg3pwqCtT/wn2QV8PkYTWjEIuElctHXVBf+ZBoRtC3z7MojPRKTy
VTKLsQLh/v9dqHMf8dSaxjMPlcf2b9OtK5RVWkdKVn+s9Y0OgfMygTof/T7J
ZxHslgOo6hGAAe1+gBUY7nZvvQWrfiSEW8T3B3BssiPoa/devXtTa59+aPuY
CqcVvdjIxilG1NRE/hectsYx6fazCAlK96EMLkR/2E950mrDwyK2RPGp9dGa
e9yetyQZhVD6NcQB6SXaaucmmXGs9t17gApl9EVVNyTv1YiaQhZAKFHgtATW
meD7OqDsJrkmsY9eCAseaoal/8Z8QKfNkZMisicZXH6mfTtDFh45t0KROwob
9DGqFxSVO2e6ov9ychfyXZYnIEb4a/RL04f7/nHZ2UunZ0s1resBjI4Td+rb
i9xGP5a6KYFhnZhVtvaM5o4CbywsVVkzHDYcLmf3XidsbOCKEWauG9mbi8WC
brrXpiiOZMbleYqK6tou2nLX2AYHGCn8FRUDij0ylZPxNM4o5oL5jrlq91MS
1oDvRsH7fE95hqlI3U3KKL391rwZyczQYTZeMrhamaFPShRuDf+drThJWFGW
Dcb3uvpcSxhMG/CRhVGfCrJg0TsnH+Lkcl97wa4EdYXRq1jJe4/x1jLi+kWF
AEQv5qu1ZLw62k6SKfBQtzrefV0SGg2LuqqrpBvoLWuYL5LR7y7XdwLU7QFr
oDEI7UufAEw6PTIcopoVXmWZaevxqUEmHNgKIh8qr6J0QO0tYX0oiFOw1lR7
uzTy7UdPy1VXZFpJ1Zc2rRFae3zt30GOO4/XxoRb0kePDPWLbmeRUfbzKoAs
16lVJdsn8eY0zES+3x6A4zL18+Cd+UpVlPojNTYMlRDj5ibvhY419HIuYq4x
8+gUe9ONMpTUz+D2cGczhXeRecg56GZEVcGmjlKErnqqN4wI+WTQpvsDkQ52
U23UE8D99C1lQnA8pBjxUXP5+TRgJM9pN6BhtnHI8Zdu7mRLcUe6BP7KTyV/
QhkGTeEPhbAAEtiU4U+U5sf/HANT/oIOWyu/QSTuPgc+z5DF+mMpfCovLDrD
i+z5FWT79eU7lY4oXRjN345KNpqSsOirFRLoMRPQH2kfPkqY4E96ZkbkDkqE
xv2HdH3LT1DXY2vSWDeKDwA6HTR3vy0yqn5OkuHmUwMZ2gxv6fVRFAbRZsQP
am0r4N1xHJDHBnzlDk5ZXdqjCiCMqWeIunoTaufdIFly8HqahR237rGG00T8
kxlPLX9s7mGyFXuAWT2zLpxS4hyGObMUkf3oIx8xgRk0mlAB6yswBt0OM3yK
uuEnbevvnoAgV2DFCL23bdfEaZHZbiYh2Xa9ebKDuxY6DqkuIQTBwmHQo7LN
tWmIbAE2DjjuchwPCisZDZtHnfRO/OQI9GMFh36L5w5oua2tlKWgt1kaR8u9
IXjvxLsIrWDrMqD5rVKkGEMmZEFMhR8aAiSwgCEeHyy+W1eof8xuR6mukEoG
nFZhuhN37NVbbHe2bO79DnAFyF/fGy+rbElgMRus6N5iIPQBh3RAo8t7KpGN
qrwvCmQLksNuvKRx8WMegYIvqb9pzPgP8bQuTPyigCh94rjPEM38HybfSIMK
JwM3uql7oMQ4a7wmvvs+tyOj1Of+CuPCTnTAxMupyO/YdsuQW2CnjzdeMx1I
dAFGJWKsAjklvW3bSj/aupbjSRBP08V3r/pLjPSuf6AHkyZm8pnrxTqyctiJ
DdOnHgqyqGbzgZp0rj5wIdpUl5wVGNVEzCUeIanJ3FK0TZZJdqbq/YiEIPlY
wd0YynWAR6QsLwnDTOpy5moL/cvflRJGFFjGpbCnYjQnFYaIT+j1mKAVBF75
IL60/YThTA7ZofM8KOfvHbBW/2sDCSxTjBK+YliOCxaq+F1blcFFE1QULHmx
VwatA0KJoHhRaoQmCo4VNbrL6lM6C+UohYFG5bX2VgOQ8S8chJzyLXeai3Sw
PQVLaw/lcnX5yOtcIaHjAxHvX7Ajax3BmI9beQoRMBpqsGyPS2ugij0hL4Bw
IhtG3970+d9vCeFTs9G2L9GGY6oBRXgNPO55qXjpGqVPSH8xnaoGg39Z4AS4
x0o5eHhbhlrVADFs6VECuIeqAZfXnkGVYCP8ZMBTgTR1uqeJYxdAm1ivA76P
nSUZ1uh+yLTt8SuEpWPZLRYwrnQro1JHOfr5Kk8wlVb35+qK+cWKMti3lvvF
dVLIkq6+HD3qPf+bdiKnHPOcoG8t5PX/yVc2BBpd+Eqh6vkzmXJGM07l9Yeg
ok27r1Yb4r7KHkBG7pgBLWyqzqls8ROhZ0b9ddwwCsudM349npe2G5F/2ceI
6IDXwcro9z63/O4i68q87/IQGKWa/EWgO8mx9j6oXgA/w0dQLTiWbba2968L
NkrlPyfvYJJm2afF/qccNniCGevkUIb+HYjj4nuXZ4ReiYj2IJoCdbwGOek5
UfBlDf8qlVZyTVD31Y+SJUiIeT6lv5FN9E2nATkSy7ttf7lVM8Hax8DB31/l
sAz67uIxHnnWSIEzEn4FVlmAbK+r6Dgp5Y2G5bz4ddvO9/opwiDGM7YyU0kV
GREjmdVVjOygT2hPsRITIn4OHlEygeVva+mxe0VLPb7gyWRyii8+maR3AwkM
ERsUlyW47XX+7maMIy+svGdhdncGMuxsUWhYJCG4wde48H6PP93mmu97h4Ve
VtHSSFHHYTGmNL++QWdEXUjenFD+ByGagb/09Q91VOz3v8atCe1sIZxq1bFK
xIoF0cjjtPLmh6t7VAL30ced8PaRI7w25g0iTDVSehvfx3LXF0QAAdgUwcVv
vyPR7tHxrPaTOCKdJ0lh3qGdNQ3WpH4eyOz7+Zfp3dQw5obenOPz3I8GMRIx
DbMdp/R17u/OZl2iDbvaa6/gJUgoUwLNoBQxvy/mQu+d43pyJx1/ph1jbJ2T
eHWZ30YoQEwFbXe0cPD7u71OBm+/CcgEtIigp6ErMTGFYqVOJe69pZS2yZSz
LthqylSgHv7pRUgKJBi0MALT+Z/ikvZdvTeawx6nJlrVJpyExn/rI71GJASQ
5Hx3iSyyBZkg2zmoilcwvbg1lYb638oNGdnL1+LGby31X4Z+tFwGxZmyCFir
V+JreSRH/sYxxxnqyqH7feAicCPmt9cKEC6SeSoY8DNh0PRN1M9HJGiknoXE
uui0O6GwIUhBcO4vpigEgrqnAeydb+uXcSnOdez2GZ6BuIWB1toSpFVcXdlo
ny7SBR/StLOqMYnltPS047GYeD4sum8NlgvHVP6zQfcRDNFl0NxtbXa9HmJd
FDXDTn5eIzKF1Xv4H7W1yeB/CR4VQIU8EUWSBMzjJaBkffAjbwHxr7f5g16I
5Yjjc2B+l4CQ1hZfF6KwGel+2lKRP/fwMGQ6IqFr6QdrsYSNpTco9767rRqP
5lZUQYAoqt+PzbqoaBqv5Z48OhPm6WtzATGCleGAA/c0VWwNWn/0Lx/GXDKB
4z6aK+esTpF3cYidBGUULkJ6HM0K63lzRu5L38khse7C3ch5qZwP99uVpa5C
g7sK5OqoRG5Jqef/Tcy/MIpD7HMoQ0c0FjxFDQ6p7m8kWHCtkIWNo2r/SZJY
1bkdP3N/RZATjvL32ZOQCTgw/lMZC3B8UWb00KgiW+70smnRhhLEpvWwGG68
oTssVDAg12vd0paIKjHPHqxFRuOsSwp36H/iIid/47p9aNheDwY3NykhquJs
TH+Bn/M8hLIdR8v4iQZ205UU8YS94XDdx1KzT0flNznlJ3tf3oHjjAzAWtbA
a3+/nDi7Haz3++Pvm1kNfjj69Lx61As5cM/hXg8Gs7xlGG74wiAF0OiwSwoZ
x1q3jx+xf4+swPv5wOT9xWaBcDwwyZ6K/hstFdxcJFSPZctkwwkO/uSv8lOe
eflUSGca6QDF2P4zUJjdLmA2u9mSEVjsjQ6+8ShhY5zZT4fw65Jl7EmfJgqY
rPwSHVLc1Vk9rniLvwcmXHpZcKyC4hkNN9qWWCrfxHPhdvUL7HDzg3hhqmK1
ppUGXETLkYh4b4d9/isfiRQ7XPmQnVHo6tFFHAM71PEGHKo2FY13wey9e74V
67lfCKNe2A77EyDfZrDrZvv3suT/gugYTqN+MQUg+gdGppajbD8RPcKqJkQ/
t4GB3HKnbNxnmPhv1Hl+ILAyFIg7OyQoF0lVA6TangMnsTGdPmD3g49zBpHV
1mRBGVkdMte/1WHXZWJ6f26vB2r7NAyTb0ummX/IXHR0uoTQHaJhZYBUVoIT
Dc0KEcXJHn5MJMILQ/Cs9Etk6zYsV9JsM3qFVuH/3gN6SUk51llQmLNTglFP
/IsswMlb3de1T8X4vvbEqmHcXUMgixtsNtFXYUZ0Hlxx9gV5K8LM0aJ3y6+7
3ScbamPt9NDCgpQ3k4FXgQZR5DYJ69SmKd3CFWpGAm2ufZO2dcG7Wtox+xCE
DLJF2Z2q6doBNqqStrIrehC9JBlPt75BLeXKH9Lz+WD/JVvTOJaGUxR3XSNR
rCVj6p7tt9AvV7Af9fo3oPsjT+TvyfumMGPyEty4hWrcmE0Ri351kSd3y6OK
fuUmZlvGthOwMqEseHjwns7+zLHFRYRub2+k5XlzlEEfNBIXuwhSrQMg+rnj
/UILfPyj9XgiIxMjP2Kmgoqt0OW5si/t4yQzGA3mFNdXC788M0CvZwDAMuo0
l0A8tY4l0jjIz/m3eS5ld8zXcdVbaCfiDWVwuRpyFeA85/o4ugiXmqFIqCHk
YEI/Qlkd8ukl2Omkci8mHtB7GOPw+PU+w63QWHxU8stpIIWEwLCy2RpqpxDv
SiZyEpVX6D36QFBHRHd6APJ2kw0aWBxeqxwWdE7IpvpTwWKoUnwzyHrk8N3A
nJCTHAV/9JvK4dG1vEFq/D6KzafKfM6oQAm9zp8CiqOwgzly2cXc8HFaJRkP
/YEH8TEHymubo5kwcTEHAIAEi+/aU06tHS5WIUYadjBE6wL5LoXMfUeCeA50
DsBQyW1kaozX8XFzeE7gLIbYdzGLA9tOgz9lBJpefQyAtBklt1wMIt3JMsUB
yze6movF67dZTGYliW4Z014OoXOQ1wVdCKk4n1cIl5O5Xb2qmv3i+dY3qUDQ
R3koAj41+8Z/bE77mdDNA2nFfGNRGtmYqbHOQBcbACaCegRuvKcbLS+26k6z
H79E9XhkB97azFIXKceEr24ksF+livFARXN8WX+ngX5+9Nx8cxX/NZuCi21G
QZNSZKZRwGimZpOD/p10y43DSYrRgvMpQFtOMxUHAnNJezRujzbUop9OoioX
Qt9tjtchXRmE7QmYeRJHT4Z9wbSstqqL4KKv0KsnzvFXmLhwRENU86NCXdrx
DI/M44wwq1WQ34uUoHeOpY/Or5cigv0Wt1oK4cHjO1FZGKmtDeqONlWP5YxK
EPyAUiC6t1ytEQB6xz03iAxpQbM3CaUzcC5rTa3OF2S0e+MB4yIys8WAAt1U
7vHXqDnf8xvfeBB5qnzVNeYkMsGy3O51ceNJqlSAYZN7xYmjTZo7aTmMQAaA
j14RNuTClh6SGfBguS24RrTQ1QcAH0q+VLtXAU5U+71zZ5OjltDwK4ZeBeDa
FHBWGrwoP+lMysRBTo7jKuVkrjcmKacd4iu2vjHj4OOXGWlpWoqKvQM19Mac
ttzXEoNN9GssCUo/tPbczfkwaMiKHM4NVyyvVodbpmcmyrI+C5PfCg4zQly4
D4eoY6BLrFN2/76HP0723wa/D5JSWiyO8vtBmujoCmzkBnpkd4/MU7de52nO
948N7sIdOo50VEkxbBKXjD0RsmiJPnJY3HaFe97aW2ymc1fz+HhJIDbdatGf
OWKNi7vHB/y0LOnjvbZem7xoQJVLDnyd2D4eF1CQtFABJw4BUvyWbcEQCs+n
US8Psf75I5d6/exsDVciDTF6IQH8TT1uLVLXRewTVU9wW1gdj1SElz+1q875
Ul6sF7YTrBTYcGeI4v5OTfoiJxU7gSBANKblR5NsLfQY0pd34S2TrWIgWOOF
Iu5LshdHVEDnotvDhQTSlEXKYmqiT5YjK+HOQmMEdYBlxc0D/7r1Dq/Z8awf
CJIjE7hwBWIg+Ml9hylZemPuCgpaOd8Ma05Awi8cthQCmaHlnEFU6XDZg1/y
yX5kFpvkgy0ITtp0cqMJZBqw0sr0jvdOOOC/0Rhmq6I00swzLsdMp6AY1+4L
HmUpo/iu7Ht4Xa0gV2kKVrXE4vCxvqTiIUdtQTpeO7U5kjGhaRkokca7Manp
cgULVZbGre0oGfwR6KLTV5B8lweG40s1EtATla8idvJWG2WWnciM2zWnqS+Q
U7A4ay947nwP7Mq0bblC0gvQQv/JNqy8aev3N3xZb8HC6K02InaQKf+TWpfa
ztrNCoDcnIZgiOrjiW+NWn9Uqej3ix/1BNXT4Q5aIxHnj5vfKVPdO2r2ZlH2
p+FlRV12nmKlaGG1EHjJiLuXc570TwD4uSYuHLtIMPWBa5Baif2c9WfpGXHz
K8saEYgatMYPzyJRyn7PAyTyi+izKnMVmkumyZTp6eU3DhW9kfSH1dQKn0MV
dWTP9K54J/ZZjJ5/WI6wvQIdfNpwgftpDLx+o0Eapd6S5SRjumJv8PiHUyBL
BuM99pePdH1PLu5xwOH1CG0qqf5B/wZqLd327BWGK1MzE+yIpX5H1hKOkST+
MTaGdRAzQnLGH8WEoMoHMT/RgLE1SRcHYjfd2ifkHyk3nZSVMT+jGJaaFeDB
bFuBV9aQzg/9LYig6IUHemSglRuz9SJ6lZl1BFOAazssHxRgtgyryjajA5B/
z68FuO5C/U7KfeWEaPcL64ZiTwxcPOBHXNNsIuCoupF8jsvJTAgJ2Mcu0pBp
tx7d59Jy87IWuPKALGJKU+mC5aXqmdf+vALhw41qg8EyV+ZdCJeC0hFGB2ip
auy5vSFM7eJc4PiN3m/r4ZHn30pT+8JmRC9Y/hHx8itauu5aMnN1fAeTi4C2
gbuWAT0hX3sId45hSNY8wr4HBW1aV0+CwG6G1nAfBJiyA9IZDVzj53K1+J0a
buCRGjOqpnf69YvJZXI2v2P7Du3DQ82JWpvhTrBCMcbsWGP3wKxXxy9YKV+E
yViFeODwPW5v2KYTAh7+DCqUq1EUoMlL9Xhb4G2oaVrNDHpc+p43uQDCqR0c
cyeymNnCLGJvuorR8s1fNf7yt9uc8B2zEiKUVLgCUQlrvLH4WKoor6laCmpv
5OxzBLyKt1TJyAK9fTjyWfQYEzKMZta0XriGOfG+rdZSPhQHXMPs8DIjOfHC
X8d0aujvFS27u2nruUYEaDWpU1/+4aHU8EZS2cz08Bqxs+B2m0LFtTyXVspO
ZZ5iHoVgvGLjvNi1VJmQrQDjJsWPrrIy2GCs02xycjpJexeb7esnww3OCAUL
WG2Kux4no2vtyopFz/ENXWa60atu7JCEQSVzqeuF0JOrtfSumXWXypy8/k3G
8fgQCnCK9TNrnfGxQuIhIXavKZQdzNdRZeLKcbPmIhGFMpAmnjZEbj3KRNAI
lqJbTZw6c8OnZjVkEln7hXm7jqbVMImlzC5mc+SEOLD/ApysktgeYmcsLli8
xgXg85pX8ejDw/9VdysqOG4F3IA1rmH/MjLuGQ2nc1NrtI0x4LDyOmK8MMZ7
B3212ZmHWxAvHLjQJlp2Rum2DWD1Y81J+1rVEZvLzDgZZDI4ceBj1ON6YLu8
OKYIlDJAZ+cFfdDvMerJd6DY8AGI9MO3mR2lUkbi/w9rRzJf7t90XdCJgr6v
I0Gph4Q4q+YcSLZ8TwX2z+xPIB4l49DXHK0+Xtn2RGPZKW34qeCAbD4bECnY
2m3Rc4hkmHvc8+7B6mAhJyRCIOG+hoQdcO3+u1A5zGJSSOmdbab+2ZeBs1Fx
zOoqZNe+xxotuzLhpi0OFql2Q/w5YC+hARe4It3XQ0ZmanGqK8Q07xy2BipX
PGlnnpp+6SH6m1F26cMMJcYlFoo40KAYdmYBQspjA9AZ4Dt5jmVSC2K8dzvZ
2lul5VTYBPBFXIpBRaKrbWF6/WNHt1t+ElrE4d1ZN7sEYBZ/V/H7kIJ3bfI5
rsDn54w8COlRGTfDiwXOQ1zWfeKbK6vAfIvH+gKURMlP+HXh4nN0kmazPYZ/
oRHp8Kb0hhyP8tRwruVtk5LsgbyPfRxHvO+CQQyU+JIYk4gFT5aMX1z5EGLu
UivkHDaGg20QkjZcA3wYlE//l3ACt4HjJiVH2SFpGQ13SNnjyZlqQdehbFQv
q1EPOEArUBGZ1ECgu8neUa2sWkEXZrbFiHA3zQvaLxNWcGcJ6x5kj3Xy0wdd
1A8Cfdo3IaZXEyDo4cvQ07kiPv1IKxWUK8ks14vPoYieNWH0w0FwyDe6Bm+i
HTZfRXLV5F7nRMYC+JBoLV/Mpmq30r6FVfHZBPeJpZa0lMKdPIZixKR5RI2X
vBqlz9eDsfujyL3IqhwQrezFxNARXPsEdcBjyX9iMlN+gmb3ENQ1zBF+0fmQ
QlD8/ISV9ErKurvmTpVF2zn3gioZhijJngXHLNVat7LL3Gwvf2/FHltvBHGc
CCRqY0U+IXdZYzATtcYpvxNIon5+3kAprgWI78HgphFkTNom+HgYTCyjnIv4
0Kwv5/HMgZRJaoRmVmiFIniXgSiSt331QjOpq/cL64Tm6mUJVsfrTn3KRH00
tNbysjYsmYrNRgZFAkCzFS4CNRJkKd00zEjUHw6zo10U2d3aymQz46nC3PoI
oc4KRbmv+6y0aG0rPtYDaoontrWEcQylA3sOoP6OvsyHvtKaSQLhAYYxo1qa
lrSlc3KlrPf5A+PCEmlldvzYq7205p+AZLSVCNrU/YmxHCnte9DEMc9AFUcV
YLDwsy9jIIingZXq/MZ3D57a/cIckQXEjTimAgMMfj33Zssa+pmOaERuBiSn
v43MBk1pbspVYtUDLuRxtMjCOOEp+3u8ZevJMQRrDH7XSSQr4EfwY+b7FI2X
ojxm9PuX+WvqXLAp0zVe/0xTlp+WkE6xeHFr8Cm/gnYWxeBroJYfhHnKjh0e
EvNsnxuOZtleK2Td6GqNNt94j5IhmI5v3cPBFX+mpi5O8l6MQquNqWeyZatf
JyEKbtkpu5PlNsbDiY/amawt+E+rP10JAfR52YIYjrPzmjD81QDCIxJbQezt
SghQ5PQmaPa6UTm3yvFUuCF9RYHhEmeF/VvhwTuoWqpDabi2yxptM9FHeyaO
gpfaEn9PKal785c2Ji797fP6peAu/QSpsEm26oTVP0M9JaPpqnzFmn/YCJJj
pfcGWiM5AgQd+4nWIzn013Ktao+GAUsHLOS6eByTd3Xj2yd/NCTt8wxWnG/v
H2oM8yAu3yIiOeeYD2PfH39/asDE+U62B5iX0rnuaEqbAxo3MZB7+yc4kw2m
MzUHGrLO46D/y95fwu+Bk1sTn5eEM/LeAs66ATXDIh8XiSfNYcGdnmKIm8xd
sdp70qI2At7236buKqPb7TKmXa5/i9E09oaPErnI/BrKycHa7jOM0pCEoQ6o
IeWS5Iz2wk4bN4MCk7JqNYHBZdcDjz+LF9NDE+Q7z+SGTX3n+H2eFlhNPE2S
J7uehDwEi8ndIKFq8cfnBlcTiGrEIKktHTtOVFUW75FzVtgir7PWSGbyOTV+
CPG3V+irBRYs8igDK7lk1yyqTu9i6V21CZTw0JRsFMpuUUu70J0o/ZTOXLXj
n+wJj9/Osaur3GDGYbkbL9teahPiOQ0ZKbMSODCGO8HTmRIfvAmYIiwRp01/
KOQmmsrBZovMJX0HRS9sqRBA2OyRSFOizycTJqgMtuloy1PKIEt0tBtPjj+i
B0BkCa7cUCJ82ee00IVwiLwl3pgeCUJfmkBSVEPylLaBrqAif+5YUYGOW27B
HFYZpUByp80Hs2jnP/8KAgoU+cf7+bxKTZ5CEK2KQRx6SEBG0XQUUwqkcSoS
BCn3kvhTTAQryQSHFcs2W3qjviB4nXrmRF3Jw1636HL/ie2l+KFglUs7bp/I
JGdKBGS1I4al4SgOg4YLLrTgoHbknSLNHskNqYWpZzqzA9mKFp8kzioY5tVL
fTG/0N/ILlYzAIdgyktdiJJbnQsmnY8r5DGeFTxZzye0I1woRywhXbSkAdDT
WLlIIF3YdVi3qrRK8K+OIODx+uvDjj2r+Tn9l67ejjVkZfmVq7QiiR7reJUd
tPofwDIACsr0DgtENTGt9mw/e5vhM5MZRLwqUUEOhHnkPov1dPaeP5y1ut46
XxFyNPhVkai/CMmNty+tnIBmcLy3YyklaRuHelkk8no9hMBA9HVR9mznIQIW
tuvWSzwcf5OydP8wZgFKDCOGae4l/2+k8+eTaieRUJd/4ZcVY1S0LZXhG0Lj
3WwMEG+zru00IoxCzwMoNlluJTbjA42iPk2C3FYnYDqPGEey6naKQyn9YY+X
1sA1IfKof+uOtQzi53eCDS2FWp0aDX3MjNmCSW05hgFRsy8TfqKSgeG/TIGC
8C0LqLWpCa4VKjT0UHA+ZtTdSGtDx0ELBU7bKcZBbtDXYFgLSJIiAeYuLmG9
SsLiWsm3pP6ub/iws0wt8w89Km6I1YzcLPvlIWh0Iu6cOyyolm2T/xrYXSLE
pUiVsfWsbR/YL95MVjXdeDiL8aEgak5wSmAEmu7Dv34Gc9hRH3QVDPt0Tl2f
8JlwL7DQPko0DCM5U8nRXlqCRtw3OwUu5FWBydJuXxcUz//oB8hbjC2oTFE/
2re1Dz9KaXtwA67xK1X33tSFJwVzspWkNGabhmtV3ut2Q6xEI7eR4AZA3FgW
Ll/pG1So2QnrmDqTiMMPzB6fvtd5ZzhS4I39TqsNX2Y4tE1E/0++xc47GrvB
A+HmKQ75EYI+XT8sfsw4mf6bg+NYrHiNHWLjqX62OHB3oF3Lo8qe0UnQLCM0
Yi+wsR7H7wZBL4UBeIaHVcWV00OlkvNUBjsg2ogCYpBfYO3WbS0QpuPDuFWy
DdUsR3mXLl6NWZesw4EwmeXEOuBCVcgdsxsOllrfL7Jcn5lyy7G8N1i03n32
QonRcciHwD0Cq9BU1JrPLh5ydEHas9KNQ9zQ05FAB3wo6YUSFtJEjgej96wi
vwhT4UzeuLUd3N4+8kyFzTYS/FIhfPWqUylEUiUbGbtDEXryE5z3poWKZHVG
K4Z7Xj7DblQ5W00nLVDAjaqQQueE78ZcKbTkOsxlqta3wnrd1cFqbalSYhB1
U58k6oaZK1/v/j/5YuluFFf3/cYmGsovhY00RgEKJBH0qvxico0KDp4x+dRo
51mC9JaBgLWX78i60SLITgZ9836D0SSHIsLRhI97dGMKV1agWf8Ea87szEC3
O571PfqYK0iEKtmYP+BWP6qeaZ/ieCngyvF5w9pmF89n7Y740JkLxlWBsES8
kal5RcypC84CeZFEgp6kI187yrVNyS8dxrk/Tfl2OfH0oz2du/sW2RqP4XQs
cbCITsKHxnIvfMQ2zwT0v6s6GOtPhetNDHQNGPl0BzQZyoAJ09ZQtNqUNaXG
ZLo13m4yy9XA36iCZqIDdGDXvpmDP/A/eKV8WQs41/tn1MP4hI2caB2fHv/t
eR8CtklxOrbSSmUHzXm9caxWx/xH0Ik9ExPb6naq1X0zRVsie0ZYndSd1mw6
Ok8P07pU2ME5rCs0r/HQPtiRUBRXpApk4H2NEFW4xCRMWQP06Lkbc7vPQMfT
y1/NhKKHmcOsfO/Azo3omMFz+6Z6GCola0r2uWdW6zTf4Kr2rIP+BhP1nx9T
iq8qEcbWBry8kx/JxQtPp57PjPUBR93EVCQPaPTX2u22kfRvhZjYgeEOZh9s
lYcxX+05R8jFy2snGNkCjvdP89oWgWVRi1YgxEPhCCj/mmm4ikacJHUujsNA
IKVu0VLxMAg1ksgvDjIGjjGtng+AAzHwdzSyVi9exZXSXKmK+Ig4Cnihc5y3
r57LUdwWMbkJRT5sdJnsekoaPKKUroMkM3SLwdEiFgUbRC9x5+Magb3pnOjo
sDrOInrN0r3C7ToTNDuuV2T4CQhZQMF+8MG6CYLoQj6iTd4xQ16xF3Waafug
UrAJT7MKCVKCoVivFY7fTjkAVN6OjXSrb3ge6gHayT0Ye0870j9zf7a/Hey2
wMJDzKGP7aKVEKDWCPFU6bvaAC+sqUQRuON5R5fb9LKX3536z4+7Sb1PvCVj
1WIq1AMylk/mxIPEXBtXq1Dja9yMu2IxFTrQiZsQ3Ckc7QMroSz4c0PM+u5X
vtuk34vcAUhOolvLAj1h8/9XyoqtLC3seAp+Etfr/SjaXvaFagk8jdxtcW34
hPCrU/1aDyNL6tygFq4j45UzlkIRE3gP+l2KPaG5SOmnEpxxmxJHHfRCxnWr
Zv4LX+SA14PruLoWju7rBNdhnMZZkcclxzJdk6eQGuaIKRzK08ggZSFjNOez
TnzSHrCC0SKlsknk35lJiGdCNk46zQ2UVJi1UaYBWFlJxCzOtG+4EFe4IbES
WeEZ6zH1+Z/KMC6ZhCGJN8AUaG2hACXccQqghNIXD9xlnZDRBC2SXgRJm1Im
/H6fM+bwRMwmdYztC2UgCP2S9fjsLGX4nRJ+ERbImZigGQCd7OYrw3JKdbFN
Dl84s1s49oFdbe1FjSoy8xxQfRm/kZd0syN2J71ATwQ2YKRdCdtDgoSMl9mB
ZVMlohi2SKWbqQK5YPTu9Y/zAx/GMF6UC0atwNNyizqOSIkSuRRjYnO0sroy
oPQxGZ139ETUQngUqobEc7VNSanU1mlmESId7EToo9PpE71FrXrrLPmWtLaM
zswrnYjn7HSVqTw69XERlvXNTxba+9yCCZY8mmKoNQ3tvBDW0tnXVzhnS0tn
Gy8AzHNYpzW7ry41/MWauk4ZdCbx3BlJqsg2jRyMUmfKcAClIAu7nKr/jUgT
gvJbo90mKnflMFyew1rboXMU0nFnKe0F2gba1bPt/DNdgybJPIKr6gqmcfDG
Lrh+MlZ5Kp5/6iUE+dWKXiK5YMULe68id3B0KsebiYZZy6qgzYxNNB7wm0lT
NAoaIJo8LK6qIY3fvlC5vNShRWeRyU71aW94f507tnB4tj2RM+ibdaGzhkF0
1+iG7f3xn9Wef4dw4ilb7x8L2hRhxX5iMNBog+LIuqwP1mA2z+oPMj4cMRzZ
FoqC1DBgGWVZdbKdo2pwB+qyXJYAEDpTO7W7ra3FcJOHQfhFdLok18OSj3CU
Pg5gd5su8YIgfzZjdxCPgK4FhcI0lmkVrJQS20GCiLMK+rwEZTzN5OeyN+pV
hX39jNI1iqnP0h/E1/Y0VB2pWF9tJI6mAqxR38fM8iI5FlEIwSkwJj84cM4B
DYnv9YaVVp77P9/3Kc0MXOKRSdEaPOowayz/M58E1wtTtOrlEKN2os6yk7VU
Sf7G8CzAC8xmKO0M1G6gTGbk9MHQv3vkh7qwqCxeATuUFHt5XXCAEK6rmoOc
n5rTlZZrVoTAn2DKydgfx3XiuxMK2R54s1DZotq8cKjge9eReiZu+Vk6tFmT
25MKU9ZioMad/Hw4iaBqzudRmbpgn6c5NTppOo5B922NB6KFWTGfuxM7IwK8
88wYpNHicd7ET0+uAoy6dVjQaNi2cQ/sas63euAD0nq7UDdgJOOnns0Jtl/8
G01Oc8ZxlFOuqUAqvkoQHulLw+8Kl6FNzUHAWbtD9BC9xRGNy/eQh33GcE60
MdOflAPkfoMiz2DYDSaCraXyboHlb6TztPcPDRye74+9YiAf+MmA5IWNNOP/
kcQy3/+hNKjrhsXACqIptx7Pw9yvBA7/jPSiJbaLLVkAIrOTZ3CzVpEf1sap
t4qC5XDBgqYZQrIVXOds/MWddRlFHvlPy2St2bOL76ivJ+QIgmGHnmFdnBif
ocSkmzuWrlL0IYwBDAGRTMGhB8sSB0DTbelyG2Hye/xfypf+s8ZbJudO6BnP
ZowTvjUMKjyfN0ASQzfgCMnWo5ksPQyy8L1Ukx2nVR4+IKJk6cPg5jEzCRG0
C9GVWo6Hi0r92XqnJuNP0gItYXK2LU3x6EEeDn/u7ePswccI4chYA8qZAnWA
eybeUR0bnWkk13InJK1YHfs2KFJawBeCjMyVawWXu885GRCU408Pa2ndhV+W
aZliBJ4xgPfcetik5ve3dZEqBEgQg6tjbveQ5XieIjZee0brLy9QSKHo4DMx
wN+YSdU03HSiARlgyzkLJ8g9BECIDI8phX3/cgtBmOlZa8tKcFQShCL+u9Xj
L6CPdl3RAJha9+MZMSj5DJqoO7Mo8PN4Js0IRNduT4ARTfORufYDZ44lp70A
roKWmD/ePknHMuifLHKBUHbfqIHVF93iXm6FCcVpuLn7mpployYdPBzgHQAG
TyzQiMwCaTby1/ZOhZrPv0wYzQLdLGarzczbTDc9Z0qqaNciem9dBjzce0O8
2602ZD13kP6FCr7hZw8Ofah5YUqmxe/QlfuTIRGe0KFrnfeFSpxtzJIcmA6y
tY5d8wi4g3nKfubBhDt+p/XnikRyefaIvzd1nDpPGot1ZNKCP7Dgj/DPM6vm
li7JYUmtql83kxcThjatLHq2BdGo64l80SBDmes6NMjWqKbJ2TKojdR0l4aC
IAa2m5z6d0ETZAX4jAE3gLn3dJe+5ijdaU2oXx7Sw9rcSXTATMQ/kI3wdnlE
SfpWxt1v6Mno0GmfrZfib0m41DWfaABJalxNbCd5ZJL5djOTtTMfi6uUvVvs
9L/W2ICvJIYXHKlE/9lEv2du3/L0YoCuys+bXd2TTtzhyF/folhm/Oc1D8cU
0zoo2Ygb00m9KgOQOxAg+loRRWqO1GtjnnCNDzDb13BBWD8X4YDbar/UmsGq
ag2EnyRWTMCTS4rxiKXYZpnYmIRcJN7Dq9sBE3F7Ks6ESobzxIwhWlSGb15e
l0jKf8PzfMqDHjvUrw8rRzYH1QpQ3dGyY8s6UlMcfyJJ1DNmXP55SfbisFrg
vmD3eKcwgqkGAneZEU2hMfgWWbtsvu1Rdm14PIYVY8vgD7H3ySuB90ZugPD4
lflDaV+HP43ZA5ZP39crLNw0oYrz6f2qL2iCPmpHZ+8Z/oasnf8xPKJsHwgg
xefyd8e3dxBvxhCHe5yKwqd2ja2WxWpjeyuTDLwYrI3GFh5OE2CvpQdOhdqn
4+XgPNPEaQsBXL3ZGXhwGxQQm3q/oeh8rGMFaewtNUSFHvz67JNjQp/AYlep
05Du7dsfDjxCwPbs6Om0219RSfcd2pRlpikAYxoDQ6GnVtoRRv5CU98br+OJ
+bNHxdJmTORZnotiTICNlE2earjYxjEshKR7hZdedtR4OOMVOcfmSYtE6GRL
IzFYar8VatOMK5FT00BfTGWBNkovBdcsm4al3XG7fpX01U1atNw4bEaarM6+
7Tv5GtHTQbIskcgzsz7pu+FkiltQwUYksQIPx/XkrKpXC9IWoibqj84FzL0+
+wKZ2LeCOQdTCB2vgnG/F45Nu3fPlBeQHN4gfGNBRwmaTGK6X3rCzTVOnkdk
GDSqyBIGO8lLN1vsjlOLB5BBKoP2bAnp7aBZsuIuwFeJBQc0lD/aiwPLUwuH
ES1yVhFMhRiY63EhpsH8nHd1WlmyRMugsxSjQVW3O8OnlTMG4nHmydRHkpDO
IG6/k0QO9dv9lzCAucqrj5bnoSxLgB8EI35xJihKqc36ozqs3G3peqdYxY8J
Ne+WOBvgGJn9/Wb8UvEo2mLvO0NLoVsoq/OPEG2tMitI1JN3OXYLYfcJno3w
ATWTaDR0VAuQJp5fJDNbg5WF3vzKs7Xt/Tc/82eIWpL4Idwn7muQvjH3hHcG
CMyj4SOgA1pwCYYxaAqyf/DiA4+wBA2pBIFPVfzHatNXN8NKLzciNwzdrQlo
1OYLrGNJvzB2v9uw2zC8aiT8AATKmqJ57UUSJ5/sKz7Ji0SGVL1HeP1t4gxT
iqJtTQ2R37wzXg8B8tMmF6dKujMd3URS3AtN5givZrMJ4ZhS/7YL3Gy6n6XS
Csr1x9lA4xEAkQ2p99MKYh8QYBzDbvq9BC5TwnLu5OnNiF+E+caBxSoMmSrR
NLFnArMWS08xS4bwzeZ8awEiAdzaGGZzEHuqR1RxHZEDiem9PFdPYLMrqMqz
Q2721pxjkfaGyRv9qy0Bs5b2OPMnD2w0e+4Aod8HeeTMpPmFmyOKZBwbmnv6
JuDVgvVJLW+XMD3LwK46w4Z2N6yzXSbKElyjEazX4pFK1U7KhyJe5pWp1/iQ
GlsOUofDVI3fJluFla1VruSPziJKYz+ZHzHtqRJ3Op/Odc/1+CTWCbg4zUwM
Z0KppQjL6E/ryR6zAYnvjeAKkmid+gwucrdc4RFgE8pfPBS1UwdahTYx30w3
u+h95K5RV0LuMv3DqbMGm/hyvFrzoKLq53rztrMgKQDRiOpN6IS1QRpdp2/r
AvvABkJjXveA3oGlkNGRIr/rYGGW4VRIE/5pXEKvKnQp3HQ7WAI65LXEdFYJ
GkrDouU6qth6LOzbIeLj/L3m8mnsiJU0/6Iv90096ni1ECiEZBqkonlc31Lk
eIOBwDG9yHc1BJrvasB8XTpy84dUwaOFscTJg9qLXoZkTHg2s+AsSrzpbkNF
NYmDkeuQ5j+rSaPptohjFMmkGwxZRM8J9by7UtxJrpeQc07wZWdZzhknPnX5
F8XU+F8SVNQCh8SgGEfLIunflL1p6Iw/0MpzOTux57adKyx7tgejd8XHxmnL
N+zOYmVe26dk34JOj+HqLQ2rL/e3530WTxb0y2f25nfiFdbmMOBTh1UweZhg
/+C9yRyJg1woh5mqrZZZAuSLfk74DDMGkgJqSLm0aHjz+E3oU1Ct3O3F04aa
5L0GTv1a/iqwxqxPLKLEoSBxNnkqmN/thuUGxeAoIZPMsmUQn/lsgtu/yKUm
fnQw+Sr5oELS958epPekw2v7S4OU0UywrCJG1mdlyC3z4jIOCQ4iiq2eJcEV
8uZIePNGM2vIwt3GHhtNvDdKkSNzgJ6knaAyDtqMawYXz86XiWh/hOPX2trM
pXQGoSyW0tKVOlVaehS3mRYdu87isKL+rxdgp2f0P7X57ghtqaqSFHdBGRY1
ROhApK0qy93rjinus4N2/2VVysGaYDrfNa+a3Zru7+wuV1Hz6PmT1YVKJk9a
t1efPeRWxShjUxKvM3aMYWyHsSQFZg7n1pOFfKVcLgp4kKFmqJt4ZWA2JydP
5VreuEX5OuwbtLN/qUzDu0piViDbT6MXGePlcetjLhY1Z7sTtU+8GInZJLcT
ihBiYx+BMq/g5rCIuLqX4sNmf9ISv/33rUCTilwpLb8lHa1NSa4HfEi2OJnE
8F+gSGt5joUDyCNkyDupfKu2VEY+cslQVJIqqJv6D2C8iuTJq8jOjb+6nl4b
n4quNPGGUcxVEzAGHoIzRxl4iFX8ht71N0+p/zjtE4tiZY1Tcoagy2P9iynu
E12haV9jaWIwyOSv5exGhg/hUw5ks0C9HvZZOlerI/VOr/hH9ZV0pLZaGMbP
3mXPiNVAzB5683tOWQ1xvWaH3u3T+91zyJeB45u5GywieztnMYAcL8g53T98
XsVrbakGbyOb89cD4R2pyyX/h5z2mjD1um67RCAEIIGr/vcYldk3r5zcJ0yt
dZ5vz4sWUj2WVapDyiCdVZLnNA51gNypCmuGbB/HmFsKc/xXtX77JopJ8rkp
uqSqbpN3H5H4tqa4yszuQc8gN2y2Wp5uJlBNujoIzmIiUJeKn82z7JFQoBQW
ktZRDiHgGVk0Xf9ogtXiiAhuF59oW4M/ZM7Y88CtOaMmnmtrav/y2yAfmN0V
FlOSfU8Y6FlCDHHh0ZtHdB2cvngHq14FmIjg06VI1ajGEa9jlaomg72VXsLP
QqJXoYVGEsnIARLGg78UR5pxaASZ9BVB6ISDMhEN+4OqSSWab8M1qZHDHNKK
ZERZFsjH5krH6tRrGejQdVOsUGpsVUQ2KLm7VcgaMTA+bdT0lAjOB7J6kp3u
MPctf3hmZzH+PjYuDEkS+/swEEPZAjMSIj9afGTpBr38xooqJHGsTtW5GFYy
BSYO8cNgDhhK84UYlF8hViBOWAQ9AqKhH7Z/i+9mp4optw0gLoVC03Xj77BS
ANKC49hxckYKGGgQdukfNpXcI2ZApIl2rxi6ah0EOsgHsj6Tw44n4AFPMjQG
7tmgOWGBUUSK5ydnhVEYSfUsgmHNfiozesrUOmFKJhAEsH3pllL308eJLux+
GETif8axzziPRIj7pNc5XHZ6m5GocgPvwCo7UR02pabaPlkftqUSvEel2rnN
Od1r+MqoEzFbHinNaqmzhK5tg1oLTn8NUbcpvvW7dMMiDXSFW4Tb/hJ+sROf
gcl4YjUChompW9GPO5bPop4oLwGaHM27ShqmUTETzr43ALxLkPbOvxtNHdSu
4SHdmVrOvCe8+mXFnW/uObc1Xza0moeRiaS2JqJo6SbaCGZA9y0FADLgM1WI
PVd/+kjpiBJ7RbchazZ1b/b7MI8y42rNeg+s0wme+ywssNOmYvOqJ7YJIf1t
dl4slSfcxigkOGM1pTLkLa2+N11jqAfZ1Q0w00YASMVT1w//XLMx8pfm+lRr
fQritkTyBwFJ6N/5H05VhrmcYUmi9Y0q85Bt+/HXxeaNYIQ5tHobsTUFB8as
9N5JxUDjN0Ly5CdMagSAGR/4/l7naFILRUlZy3qseaWtYQbOz+fbtujt9NIA
gbrjw9CShM6JhxMRjPQLzB5p7BwjxIQ5FB2ztIxxDybb3ZD8zPei8LuTB9U0
sPbSUAmVy+Y/lQoPcpzwAmswoL/5Y3u0X8leTkbMCdN2xn/7JPcJpPdWYixQ
bCXN1Kh5feiN8TEbv3tLv2dWk37Eddbk4C8wVeVgn+ahlYhMtP88KYROxy7L
QKp1z0iA4RWFCWWpSwhdb6/lQ89L6GYwTinpmFOXAGgkxWO7EaAvmNZWggb9
yIkjgJHM7qqpA7K5GWkg+JluSRLaMqdQqRKTl7O9EOvvqKuHfRqODzWEFv1q
3RdXCoYE1cBy2k7BWefgeuiJ7N7jBHN0cnhDPFgxw+Qn4g2mcuAn3hrFJ+4c
/1bLydsuRQ/3SChnANSGqdBXCQgRWKAlDfVLVW1pRZ1eqpmYlZT/ujKml56c
dNgsr5FCNZXSK0xX4TjABBxlHriSQjgEsNdQBGQjO7HgBiCIASkld+1LT0wr
dbE/cwz76xZMjVMRjUqM1yOVhgedi1Nd72CFWJGa/hSrkDkTINrXxI1H6ZBZ
8yVm34zfMXeSPWl8ijWIfFlfn4u3HMlRGWAsC6PcInASMgoNX5wZqVH4hav/
e7hSY8h+xlpHFSdya/T/YVsbhK45GTsLrJg412N26HFB9SM0WxTyiRt7q9cS
DgJ7yWDUqQr5ZKq0/fJgZWMScZfEZCnrLPjYrXYRE7OhMDPhb0PvZTGVUShV
blxRjW5OWFanHhyszgWlWSHioz4PGF+USH9sDgXRG7R54FmkS4Zn3cMTCbab
V3pPmKiKJiJeuESlf9hx9kPc468Hbl9d7savGH0vdFV+SiDrSxsYA7m06e5V
aQCTzS/6LMzAXljBf97A3YXVAtuqOKGx89LZ2hjreWAZMfYhlnhEM/n+YBnD
d9/9Mkx4K4iC6xf19qbiO5FfyHsuggwqWj3nqNYFZarGlhvkhG2mfSD/fvD+
KlHPqOB7kPog1IJVrsmM0g348qzxdkyZYTBnmpbcC4T/XiNVHLP9/xcjfZWU
74DloiIVlY3xKOz9b4bOQ/XKycONvCtZG2cIYP8B5JfDA3UTCByC6ROKIV8Q
PjxqBqLT9RfPJ5ee88v25G6X+b9pR4tdchXKQkWS/DN78h6KSD43SHzor2A8
4Gs37DGaf+pAkvdqzjKiWo1Xhx0M1xj6N63QDG3zjMZj+2znvTHnDXBOHXhK
EcAx4KMnkmsPCpelhD52iRXqV5uaUTwTSJA/LSFincJggjcWHx+ztSvPWZAV
XZpxvHPherOnC0WQuDLbflPdDGzA01iWKTFNNCiGQ85G3fg838ntLHgIMZH0
8H2antcpIi/KmJS/r4rKRk8aQR4mrxAE8HSFQbu5jVxoTTA6OGfWpsuHtBpN
QA1ZYv2gK42qkP3tvIkfTaaIO4c9cdiX6OCoXgtb9QIPExc4d0MGUkj75tP/
wGKkHL/fprnc7PZZHx3JoJyfYtURFfvBUklqDCKcaN/oQJ5Glk/iGFxVyVDE
zZuedJoNwut973cDuGLrn7T6VJjJoUARCi+yhw2ghA1WR/cnD+thhS0jIgIx
//jeahcFF1njqokphqFAqbIf6EuzM2nCB4TnikNgDYHLwsdFsUAdzh/AG/X2
hrKoGj9bVRZM/INalU5LpPwCp5EVSEcrytXglC0ZaN1TA+FUMywnsl+MWhLu
CAvMlk0ecXcwyPn/t6+UUHEPizVSg2bBqiKzBBLg9kTUihcsCfe9/6mljgFK
//umcnuNiffEgvWXgHDLX9q/lo3T8g7VijNi+SGkjzS2Or8i6jEnl+0vkTw2
Vau3tGQOxjQqBhKaSGEfZOTU3N3caeVvW4WfIbQG8DDgs9i0DvBnQ+nkAYmE
+NF0LAJrdhMa+H/EqijnkSee+9cV7UNtwwj4wOmYd7vfkHGJl7FinyolqzZf
99+GLfaVljLoqDtVS5xwGM2aZjtKemKm71V1QS3N5U0oH8AUAaiGsbYdBdqc
mCJBJ+FqJgpX0XEEQnKZFr0lXasZommE8dDyynewbEf4uJ6ZnJBM6o4n6dng
RkEiyT8T9j2y0AVebJo6XYX5uTb2ETBUdnsmMYyqduf7wxDgdzUFEeD4hGgk
kZW7RF0QCd2q2zJrPu9lm630J7s/JazqtdQ0oMrEkCHsabCyRxtbil8F8fV1
XfMn7UC/pWPfF3VhPi0tE7g/mvjm1UGeQ7ONneccvOs5Yrd3YeBfe9rPr4G+
sw/gH7JVfxT6oMhdl5UldY03nd2TjofkV2idCNDPGLpxt8Om2vARKg7TqilD
eB7NdC3MeO6VgQHf3HN6y75UuvQFykwqVRvPIwNR6BEl9z543CfCE9PUKX5Z
O5v2lH/Vp1RoNXXX5/LQNKWGJTY5nxdBJAvblHoYeHCbiL8X9k2iSRJBNOsz
QZP6zkw3fY3SnptRlyRN3CPdyXfsMPKemx0VGunut7LQI8xjtY80q7rrPxHD
eljk8EpCSRzldqZzjiZINtpTOEwiS3aowi5fHP46lsrGSGNu4x/BnI6idgne
FZZald2fXTRTGuTPk1W7yQTyXzYprC4Ek14fuopgZRaie2y0yfd17aigKSMB
Kt92KPxXnoSIihnpPK5auBvZMXSZ+QtMWsCKF50G7s77XaeATIhiJEEEUCMK
2ZSeMeZPECvveQhlW3HW4wxgLu+fhV/T7SQ8YyJ13RIShL5NxmWaL8lQuzW6
sNDMvdDuaQ6YHkfu2qhfHlNn5PHgyp9TaHMWdLpGtetW8AzCJfpQt4UlADpZ
af5NkZLdOUzh50zk5QdFklSx9eNVEwk9WcZm7DMT2aDoIClNDuUKBfNfYqWX
bXf/yEFeMXCwnAFa48rDLf4mc/Ps1c8QStKizsSCixS005xAeHkNmJMEr/cU
GMtA+CkU8YyIsmLoJSw7rLPQ8dvt1rU+Dclio8Ckifo7uM7hbfpNtgaFB/2h
Q5kFgwEWI7z8DBs8ji/LWNfNa3dwP2VWpGo7GsxtHc/LtZRyMmqSruxD8McH
QJj+3qewrydDq0qOOYAhXws0FdogqDKLJNY/XMM7e77A8nw+HBv9ttnCf9Ra
pVzzokehKl6goWLVFx32GoUR7vq3KhWVdnjugxuVvyMtu/HfOo2viOVDRgSe
TuGNMwPZ8bpN7bbBzZws3DxnqP7XmFZ2d5HIItE/Xmh/nybza6NrO91349Ca
150tBdSvNp3DRejqRt/GE3hgWfo+dWK2bBPPIacESn7QD9anK6C+Bg8ufQ3f
QtWybcahSwChUTP5HPUIJnmqSD5EhJ7o8NfVD+uRB9Y5DcRWDDrfaPYapwH8
s5k7f9OKQR1k3fqVBGdUMOqteELdHobl178O5vZqv4CJyOPBCz/qpEpWeRaP
4kD28blABl6M3oV+M7V3+4ZIn2i3YRP/ZHhZEE7JyfOFxzVWGlhiB7S22DLA
fb8OBylVynOL9QmPWwRwBElBz1th1SxFhIK5iAhKQKSShTaSZYeveHsMHOlJ
xBTQ4s2COAkfFsOH53OstMIYOQGVWmHFlcWMzgMeVqzBqcvqUreFTgTPUsJj
HNYsHFc3mZxrSI8T3+jMYqnpbdJSCQ/n1YVqeUqy8aL3EwGQGKCJbmns4Pvt
jthc+T1Uqj9LYs7U23Q3iP+fgkxRcEruRPRibj3QyWIauBLZVXMhOOsw7C8z
QDHHF7QrVdctWLIHq16qlNoh9mIvl5fGzZzWxF+duvxYFq34MYLQzIpLLuPB
jWeH5n6wiLxeHvqIlOQAtMyAmcfKpXtNbkg+tkwlE2BsLtD2J8b0+nGskLXy
350D0d1qKx/FbcJwJcrEnG4mnJ7b4SMzFlgUHi+AjVScI2ye+fvwhNvtXENs
aup72hd87Rf4XMMBaL9/5b1Nyxk1+B3pXhbclmTR/bFY8skeFZtK9T2MyzkN
hrfp8EUlfVV2sHQp73UyfoCGJC6sIqkpc8N3pksZ+cwssPIagEhLEoCtke71
wTEBB8/8OMyXZZ8YQDFjpkWPCc6ULZpUbqrZqYbdFyDXqgzqOT5W81XoPqM+
6r8f8ZMsOTLa99BmP/SE4o9jfDZXfkhLP0RTR8IPhTOQlj4cbTsTMmgEKKEq
prJNxKfQcsmDKJgYg6aWpy68PxWZQ2mtGMamaxmEqIgUH95WbCcCn1NoSw4v
n9JvToMzr/HeNNgPbzoLEibsi5RWmFhdN6hjRCmflBTmB6CY7x8P0aqOGHT5
sOPdQfSaEc74WDh9TQvhdNQItoX0cyjRdCxBltb1MvkGio8vCpBOJprdlXyn
WyLyCadpQKFiQ08ouPGvKbES+Xe4i9cBdL7787GdUfk4XOD4fLUmZldqhzzp
+tnDIMQnHO7DKCuuzyAJIkgtvdom9CpqkalQzKV3Z1CUJEXobTzDUWEoisVt
KlRttYHohy/I+PqtLPHrKFj6dDzHwM5ZEA9LNEbrhHLLNzrDmMex/VRaSoOv
WKDN1o4O0OcV30N5CBwIjLJhEd5Qx122xD/iUpHgaw0Hv8xoUdOcEc5NclU4
ZTxu+38ShWtmlcEL8vYIbzEtFbSZKPkcVv8JyABF3CF7XgctvVloBZdVDglS
PNGJJNOAuV7JkDzlcP8dHL7JfKehUfzSsasO3p6hT94TOsjqG5IQ3cSIYSas
+xA1uVzVCJNiXVaxccsswJff8TF4fCpvY8NdvQGpISTXBdnEmdUaTqFhpsXQ
T9tBpwryTtLwIM7WuXmR+EeXRoLAmd1RihNKg5VG/v7sNbGhCZ8FYaaLoALS
LqIB8oBMdq7wyhHhSKMiHB42OveIQk8f+G6Hwd6dIVxTD3pAM/gBHaJbk9aS
hlPHDEgr9/qbv+h/6XEUfz+9Cn5lUBnib3wHtYztJMAEIxcGRy0vGdkDmQgB
tufKSS8eYqgG8BO1/udjldV5H9IMVHPh78OgI/NJckL9b6syeWVeoGPJQc/V
KvoY+hLIOeLF38zUinp/cBtOSI50iF3B9HjLQW+FzvXHLwH4ymmkXLd7BoNl
qmqTa9DAJEBEitOw+RLhlIbcoU26sCprGQ2ydUjVRwmTlvpsgBOKvEM7scaQ
CP9HmXpllaEK9rT85/bx5LMPRJJbjbPGAbjYl1gIS9JvnxYaYDIRRnjF/Ejh
VOp1+N5gcY0c1YND55rhThlUEwXdLL1kuvmB9d9bcS3zL7fUrbkDzwLA/x5f
fWqFl+aEHFbxS9p3NE9DeBLVbOnie6xprYHwaDY1yVBHwudc5rrneNHRiMhf
N9py/qS9W0cd71vu2WNJ+TiQLkstLJ/U04gT4VIUZAnvwI/wM2Zs1mVWUXi1
ma6oj/7m3E5gzPKl3U6EO+jPeJbS+BJuIoMyk/q+jgQqtL5pMZCsBfdYwLOE
06P5KgYTfNMFVJCRZGoo4yP4XHtR7FaxrKBe+u7xPiwo/nzd2AG3PUK/8hrQ
cw2X+f+iOMd89wrn47w1TRf4hVvXBdQwd8WR/vZaLks52rYa3CGJnvvgl/Ew
XlIt0yDJbnYNflJDghyXOLLFvTOf8ap2f+tlGlAcaCRCdOyGrKWwO3lYxuRW
39GVfRIFNM5H6Hf8yeMi/UOrICyFhpi1LSgtdoOOA/dtK6dGjauN3CP1k5TS
STs9Kctt7USbcFXXxlX9ZSIJ1CVwBNogVlIh0QV1P80/2na90/TdnkxzDGKB
TEHXu9O53W5Zt/7swHFPr/OG49lA6xn/dCZMif59VApNsxu3nJQiy/VY9gMv
j+ltpejAfwCyiaQc7jy6KO+UXbKvWVuvxBmNQjzEruBdBW5fHrBTAlueMFoK
kv51xDQY6mbwcJVr+PE4kwKEHWJ2wjG4B+ceekqI8ocBV4SB46JysUREvyo3
imdIQGD/Rq1BDdQ1BYqPRhvt0kyyoaGRjTsFw3XFA9r0cYOwsDMrirpNKb/+
ahSg36dBbO3oFIrrSSuG176v2rHz8TSwDMz3gN5fWn0oyS4Bgn+geUkbSoah
543z0rcdPBv7oLVqMl+b8TFLcEDBlrxWLS7HXtGthfrL7zr19yO7oKqR5VZA
DScOqJyyXChtwGtm34S3uKTtkIPyArbcItgRASB3gKLKxjix0WaFaU5BxfRx
yuSmsop6xI2D0jklybRUpsXszNMm6jRupVmH02Ur2UGIQZ46A8MTzyEi/qGF
0GD+/aUvajqACGwzfI8nw2/YSdPU2j900zUxTAfWXor8xsYerXbzGd/knwNd
ASzd1Y9QZjyhdPUB3MCbn5K42RKdqIK6cTfElj9rSQfP2kn+ipqaQ+3+WJ7b
C7DdwCdmy8+ii57+FN/WOEmJQNOwgc1tgPLXKV356BzbIP10e0Z4nWoEpYp2
I0HjlmW0fQc7mbs3znI0bZ4vrCnpW/uaKBee5AB56O/dLzjYFC5mXtMnjx/a
TWz7K0SosSY+dq8+tmxbun6N0WIl7h3sG4DwN/biA3YoEaQ5gnhbngQuaLO2
A8XtA7tV13YgT2vd3p+H4+WqfMn9lhz+19xJVl32b3vqFKION9DtdxaAxnTe
pIYMiuke+ayHGSyt/5KfmlUYZd9e3lD/Lrcmoq+JwHDu+PhpCswyc9Rb2GGo
AuR+aKd4ufH9kmPlYk9HunSFOTKmL2aifxXX1mpmYvxmKeb7+iDVHtqeajSm
4a0ZLI3iCXz4TjeZiufwV3vj1OySpqqUJb9jsKsb0OMI/xclNWxD8oX5SR01
GmORH5suZJ2JlDPMxGhE11Op21QlJNStIid4ynd0hOKaWyfggs0P29qckSj/
t+ioptfOrFudQUgEgDDU4z26JuJ4ht8rakTmSCNYmMFG9UxRS126boFbK7iq
RcJCH9Li6e04P7wfEyClSROTvsUEn4+bU8JdrCQAE1NAcx14li3g+wSzy8eX
rSQR0c9EnPAuv1vCB3tr6AJSRzI6mQQRnCoIaGy8yNWFT9o1iwwXjxfzJISg
TkvbVn4wGUvUjgY7HSBR4CSZcMpW23QbWQ7fT59UX0NGjN5UtCJ60xtCoeDN
f3kxSu60YetLsUx/ueW2D4iG96JEv+lDFWKtTdswikgVMh0ZV/oLTmftw9hG
m0rKdBCl8+aLeYajhfuMKWIbQRGkS0uH+YdWLxk6c3X1GNhwrhtMVIzBB386
jdRHQIgA6/sP4nzUMV3ncqKoN+q9JVyaETsPR2oJWdwCpPJg08dSYf5wHwQv
2zQXFt6LAKy4RcfiLA8W1kbzEHYOT4z3JmjI7jpQ+jIEJdfYI3+lCzGHY0Ho
x1aTWc15HOPl2dniu/XrG3JMhGV74iWEQSh1uB7sas10yVw/qRTd+FN6HGhh
Xn2+jyqHfFNrfDPpQ2wFrd2qxqT+y6PaGQOyF6iQNip31WneHo3Wb8Duxu1F
Eh/i15ZgzNefDIu8JAHexszNsKTqDsfKkFteXod6q/Xw+iAsF/XfsQYjk+sy
9oWhk4OL9mqjtqdKU+CTOpB7I4blbgrTPxr9JtmED/vBo7ox/RJ1AZbIi/Z2
SNkpVqeXQkA+sSA0/jyCRjfYfwjiwKS3PWnm2xlxJxZ1uzQJk+rGOtUU3v6N
TlwGIIx97SfdPnRtWXhEBVu7BIqUS/buQT0JTYkfrd/jfGlCZuzzDLcafYj7
yuwrGcTGYf1YNIa6iTaEPfTYulk119pXKLWSQM0DhunljW+xvMi3srDkBY7C
dhA1PCPhV8+gSwJgqaMtgoUtXW+9Oafj89HHdKCaC7Rw6gRruO2ADsKh3AOD
YxXnzT8RDnOXdc27SYg+MVPxMH60o/0U454KROThsMDBQXG+B4XMi8HJyGRu
6Y9YOSZCQ2SosnjKpnJvm9HH56g0/Y2bEXe+YPiBSAhiRzMEv2r4O0Fh5OZJ
MEF8bVHpJR+ffEMF6V/IWZnnveSxj/QlxoaWbSrEq61ByP/n0/sjz9BpTLBZ
PzwUSQ1pwCIt24mGPmQXZqd4qPQ2BiG3cUJ00E0j2OReo+Id615Ksbcm0gXR
wQWiA7GE8ZM2XNyBDAWUH/dMqLjN6QtjgnqOz6TM0/qUGf0eOsL+iCUWQ0+s
kZVsXKQDxQG6GpV6JCocswIRWDfpbSASlJgpCLpsah7NJhGAiXIuG5PhQbaS
WrejvHhm+qIhVs9fCnYv20lrGav8FL/3JNQKn61ekynKFAO091aU6ujSnZJe
gPswn3Jd8qPNUOrRCJ8pNrR1FsH3dCIlW9LafyVmkrTNNyYMrqykm4nHIFUS
9aShsu6JY62cv5DLqcEoU4gaeeLFhRLy64ROzhpixdb7XmsQzYY/qBLS6GVR
nC88EucqkZjecWZA+0jtNItFiCN4JuU+pNzSKMHbj5bcjKZcxQbjCjvPAAmR
W52N6cj2fLTV7hBuwsT75dcX/yhCwHqOBerLq96XGBPncKkEvZapfu3nzD7s
5S4ho0i94L5PrMD3DsMKhkwLNop/q/teGejI0KWpyeksLGJgufYF/HlMtRRl
9vJqvN9x4XNjzMOA2GEuyMt6UvmJ7p+dc7TyhMDkOMZSzTEbfOu8GXkIlGdz
CAgRdEss9vLtr0Hqo+WkzckudwyfhJGj0kcDkL3EopFQhQ2SWd+/ARpBkEs1
bjO1UAvjBPflGfT60vnNa4IGKfJ6Lf2i440PaZXwahDKoyrqFqEJE+kmsV1S
qPWkjjGgu/xrwBJJavu/zi+J5MxaBvYhNxWPw1ZlyIxJj745pmOZFGqHNSnJ
I0UB+F5qbYkhwaOnGVwPi306ogfeD30Ex7knQq8SP4KaF3SA/O+hAg0edM1i
YJ9hj8g48R1spEouNFu2PBFTMUtsIE46+jYFthDdl42GTuoT3SuTkv+EkgDC
IDfjMlH9ovRIDes4Ka/X/y4Px67b7VQNc4BdAFzVZap2kQYqUvLxONbzpqjc
z046JNCGl5/EvFYZGFuj91ObDy+dYlnFTOtGNTW3m091Q5qkkkX/W3a6SEk4
1rxjHpHPtrPcZ1CkfoI4/WkChAirlrvLBTQEaHPPGsPBAq1QYXDMtUjLO8f2
j/Z/6+/OfGf7SCIR8QzPB4mwnXLsYb0dEVk1oACYHRgoMBFieWatO81Pcy22
QyDWeDV3EbswXyYapltNgywYiaK+PpkskCozd5Hw6fZvDVL2coPZVIprZ3mq
DsqsayM2b2iumqJoj3hvP9vfk17VDOdzSpZK2G+BFpK5kRdxWvwIY2RHaN8c
23Lab9Ote/TmCIFsm22D9Lw7FYWhzomEyWOT8dYMY+f2+gt90Orzj9PveJPb
AnBjD+ZmD1Ij1ny67f3iLiLXPCRgVe3HzRIckkrLCO6j7AV6NCA9dQKDf4WO
BtAuw9Cez+CgXGQjc7bH3pFuxjboifNc0IYtvqETTJNf4DDExDnFaVboAcKN
W7VutjZFKM0bue0JdWCL9Y+dhNhp/NnvCQNjo4+WFnCKFcXckoshm/+z1Buk
D3XpXeKKVHRn9VsLzBPr13qFreefnqSjG+DPWVpR40KuQnmKMScCblvVY4tv
uQB/uD3/h6lC1648RvEyBIRHi+vyGWnWNh6t4n3x2Uiw5EgZG1ymVe9lCD+8
lsdPhaYC7TZuOHXeeC/hObdLL3uUqOEXt3M/rTmAnrUrqBHGS3drpc2fr/kH
QNhPcz2itJJhiiUsWdtQjjz1lvib1OWZ4evW+PNfqRNkCm2B0FJ1sEhHr1Es
ep35lUNyvLjenCWnEdPUEntngZlmHSUSfiamJWBYKTUpLe0x7SAIbofFAsuJ
7V4zcDFbgt7DNQZAP1euyy2ar8nSsl3Lr+IxGW28dkap2uf+wBSg+RtVIYgO
HtYgil0TkdSlgZWZwoIZ/WfvyG4G/IgShakyCzqJbxsAtW9EA3iviXc93Lsz
TUL08kdkx6PWOdrpxNIAQbv9r1GDrGn1vCzBzDlZ0Ai+gEH0FIdEwB0xU0I8
IByfft+UpQjwfV3lP4rNDK2+KeXXdvw45Q9xxDDXInnc5F7cr9oF/ZEco9cI
qrnjcMjRG0H4570h7x7DgaOWBXO9i8c7khl+TeeIzqhEl4BQWTUVAifB9eh8
UPN2wT8wBHEx2OWeiO8J5lfWyi9Y5Qpsq6Elw3Mvst5bEzC1db6obEKT5nl6
lADA6CAiq8TK5H3n8q0a1arraR9+l9MBxZYe56Ahx2gjV+shDdAnqfQmNE1T
ozjihdb8ho63FYuVcKKXvAo+JKI27hKMeIjmrA5tBzMGzuuqLcEBMytytrB5
997/e/hdIlaCM1n2ZT8M5xaA29mFIRScFSiSP6O4T0u5tBwGgjSBx/eI+Bqa
h3SkmLOd5MTy3GZS41g+8NGjgY2iAIVcU4QTlQHRThDHDb+0/zI1bovz9yVP
lpXnopQDHA6ZNKXJGTC7J4o3Pk67Rn+xqWqMsqmJFJfqvoZ4FfWRUfnZQLzc
cXIlsbVN3dvRFLGCiIKP/O5E8Tthi0E7xIqincX4xSY09P+BrJHczt2UVVBr
PYkJsStc2MhcUKV01qFWLOCrThMcW2Qn+n70bny18bODT+8fVeyLNQaZcs6Z
KirHIFlFtQsM/uP+OuTHVk+U3aKaFN11QTB30tR2Gwc/YFriMjPmlbel79id
+j0+flftEQkf7KCY9pLpcSorWzUmBe2eWO96fytx9rA56IRkW74DyQkykx/x
AH6TDGXhnm3K60tfetu/CXrPC9kt9uSc3W9UNXnm09QYuPbjHr1Wvhxu8vFu
dR4MxkCQF60B1VVsMCnsElBihm56qbzodwsUYiT/Xf6ms3ddqcRpWg/pssyk
EJkysXZPFqvWfgzWsDoAGXQs7WXKxzyh/QGygL0NvwKuDYhS8Zx6fE7Cat0x
fP/i/ZWHVJD+hlACN9G2j2P1W2cuhft7SX51zJb1WZZcBFFh+O19RWzILGH3
d5m/5rgYsVtMr/iP7ZTB/HuQjpAezO34d7rWD/CThPfG/5euFuRzkEak0f3w
xglp0kwczg71pz/9/3QJKHcKDOQc6DxrxFyjoCEhQvYApIdLFcHzT1SNkR7v
swZtsrfnl7GLxY1DMrUFlx/AAfSQpHo/ungxLK28IzAX7TgmfFuXB8MsbkJh
jEiza3xcPhpO2kF0xgDfCGt50MYN3u83VbUwYJC03ZuPYDex6q/sZi0C0iRB
im+Tvw5i6WbSVAtbZWdpsw6XDsjUm8jt7YGP7Qvx6FCsTyegQvOe6gRCulBF
/G82Zn+ybL4FiMbOfinmjgKDs0Cr20+u9g2b0fKmb1axtRsizRPoetgeZD1d
3GY2TY1672aKT6GGhGc7QkIFxVkC4FgYcitQJLUHOthD7LvDIIWfR8YrioS7
rPYVljWUCRyq/YMtkgWhVLeKgoznAuZcGKS8Uqb+hSFKIi9g0Du55OpjsoOl
TuUEr0jsRc1n+3PdM+3deJBKrHqbDzHHAJ9qoqvFkRkLO6bkF6Yzn5YUaPDo
XFJ/4HXyZjZhpgEyXi/AfSz5O68NHxb3WBhZCgO/KBjaPRY+AojLmdkQA0yD
VXRVjjkAuRl786evhFabplkLbalsnVhiYcPUSWMQ+QBqP1IpoB9BWOzm5Kve
kkEAXmiKL0HCQ0RHc44e9Zip4dnW5WChlR26ACY6zfzst66FfNBMenwtOdiM
QAUrcvGujCWVga+wbYAciSByZ9fh+D1sXz3q+kpgSO53W+UYLkkz2yQTLw25
1LdO8L+ExG24fHxKnYv//IL90kwQbfVfruSDQHNQlKEDsb71nAEXgvTmIVJk
26xvd/jc54xKKDsQWiLLBFR+Dt70dlfDSv17UfkqPzVBhR40EdnSDumbSiSV
LsaLqEcOmmd+o6LOKDMJWG0Shh6mWxFH6lzDmKP2HB+ZjjGJ8ad1D9nQ/+sE
aU44SFkG2iIml5Jz3k4sJXzCthbYQWaP0Ol8Xvic9e+9GR0Otg8of9gh8wF9
IkUjyERiJkdaGjJ1KwzUYhVcb2CskzjqnTDiuuCA/U3k7sVlIglSURoGOn3V
9Lodnj26kuo9JvyeMbDpBcLZXDADCTOhAIvf2y6mbSyf7MnQ2eBKjQYfFqtD
3/zFmGgrDC/9lr1rCp8LwFbWjDD98qpSGWn5eowSPgqcScXstRYtGASDRTXL
U7q3SA8vM/Xrufl/03drQ8Y8P7MKqYh5ognfA6pAtrq8jdfAdslKGcCkmL+S
v4SQYNKOziR2HF1uB3pc7XiHQ5zE9y1l1p4Ompkf/a3avZlO37zP1AOzgyc7
2uw3fqydn0Qn8M0F0FOLOObE1d0Msm8AdMDRA6pEIuofvss+V3CkLl6qRFu+
XOFhSQZMd/HDDOB+uH5+5WGtVNv/1r8PPfGnzphlQNQFFOh3znAEUqytbs+y
pnIsOb59YrW2kbaSF+C6nNyGA5FTDWenDtXEDbEClPBcTtoWLHu5QaKpfk0F
zmUr4Z1VbKU/j+hOy3m8Pq3xHP7Ih1GbTmHHZtR4a07sTUUdlTnOqJ4iA+tv
SnwP0uS/OREqcRZKnFqYKj5Sfa+4ZLdn3X90m2xlryzXzmkpWzkIlCUL75Yx
A9Zds6fel4cyB3wAYaUqE57wYq8skoJSYgpCsUl61LxwIO7nIp0gEWBswVMM
GHZayQlNBeAVk830WP6VWyAIaTXcohJdL1qdXpvA98gr5ldVElRcF5CVV/Ds
HUTm9ucFmFh2/RFt7V0ssRVLbUeDMIUsLveLni7z5hahqnwvWCJEu4//G2fN
C31gm2wI7L6ubojqZ1ybagOVKxtJZu2xSEsKBH85t3rSosIa3qIx5agstRDg
AsnHEX3XnDZMP8X5KWGnjLPGgUYmRHJRjIyG+1GRzdVyPSfsSAPGJbiaOcAw
rRbA1n00lHlSic5Mn803POtw5ibO1jLTtFdMuDXxA32gqcD4bVVp9DtYOKXb
D/IBZ5AqHnYjtTwJx/daIZEE0oR1fJgAmtBm8BPYq+Mrf/KdUnPyJL3ALJjs
lzp+lKX3DXSkQh/i4GZZCptbW7iIuQCI2Ff3MpOdwtsMdlKx1ikYT501qnJd
Mehsu1LCs3ujpjIhNlwPHhF1EeXnrnYwCe8W8cqnQs6t4yCCwhcGJTakWW0s
pKPTqyE5GVJtJOF6c/vvBXyB3q5+z7IS9CIVk0dfZrk5xNpHgJCQidEBZ+TE
G9UtD/TouyRonQQtqE0r7w0f1CPRur3w63mjvfU38U/tFtyzWn+BgaaPGAEs
odqa/qcytdpkF60WybeLsfe1eCnnicc6uPkROkR4OAP0ZzeQMDoAyYDS945k
/Glq6RLYPPNlbNLPvFbjQR7fIUlf4YuTHMCLuyGmzO5/hYY5D8MiT8MHnGvH
juDactAFqmnl/tCsT6AQD7cOULx/AFJwKhuJhEmkyqWKqV/NYzcgwOky1NaQ
UdtEx2SvYkxYfr6vBAkHUIvnhHbiO/LhhxCLHfGdomoAOoC6zDs32S9M7VZ9
CYbBG+xjACGjdWuKv4rrlbFRyQSST3/X+rliipJFWrnNVnmdPel1aXM9cM/V
1VL0ut1BdZZrh79+tju13MY2Tgn7bK3j7bwgQHAAcOS3oL8CQ0AVzE0jgHUr
s9GvQGlniBSzuARE9z9igB0uuqt839vJMiC1Z5s/AuOFan/1hm8GmuRcPf89
3XPO/thvKkmuRw9AnzmpwRtQbkUbCOUpdcytKYUvKvT7fSlNZAV6B8sqYOao
kOxt+h6qhMfL4lAs7gI8o+T7AdaCa6V8WQaTzBGsSyCCk54g6xcE0pfJ/0Dt
YRtwL8zUgsfwFvhTqt/rN36JmvzJy45V6t+D+r6H4GF+bmOzbBzFiIFfjniN
F8wkX+aFiHRDYKwzJp88I/zbsy3GGx/sM0kZXYvBj6E1CkCgK3upzCq2hrbT
a1dXsPtEtL/v3FGMvB7fxqM8veYT3ufelq2AWJq/pZLf+wYitI1hxM4b8aUt
oMe3OZnSPiflaXeJ4SOuWmg0obg4TsV46ZC3yeVpBezlPfAQGRjDWUnbau6m
p6fK2yGYPwLMQmS76k43KIpNuESxHbt+r7TNX4wMLptUKpBgs7Z/lhaE7iRG
NVE86DBtFoqRoPqYzI3Sxg/okVUBHpt3qkHX8vosP9u2x4mbyTuTReIdMSw5
jbmfiTO/k+VQUOZ8FHlM9UC8Sl7t/gyd92dIg1Zj1hSr0xJnhQDKLK+EtqB4
6FL5VC9JjFftVqlUq7mtkaXfc6Cf23lvVb23TTFJvLpqkKbTP3rmlUqz1Dtc
S6TATuekUM84Fj8hzkrv1f4EFleIAMO3b8/SYoKbQNcarBFtt4Je1F9C/JMB
fk8SaIvtBnYMMfGFVa5CQZkqlWb+/PyOY8BF4xpI6p+MJYB05NUH3yyvXkQY
+cXQ4ivPhbWVZzyGPVRvCnICERc3i7z3KJ8/WuV9ARQ+csI/7JCtvr3+a4vm
GotiNVhwWuGtWpEWn5fHLdRHSAxJwl079wX4oUs2hPbK72KELJ86FtgUsSbg
x8WACDpmgkM4BZ+pfFqmQMKM1yVP3aoFhWEAAb8Y1ApmOXhikA/ZYKEIre3Q
H/yeaq/EZZ6IVYy5y7XQrHGs+WplYXELgUUlN+VCprY3BUT9OPhQ33FhQuyR
/QYy6X1u3SUmiWHinromHqDLgobIgDFClHIpBNvTTiRoOF4nkCfooAVDm0gI
8qOWRIefbjI05z2HxuLc3oQqMCE1fsVoFRw6XPt47F7/XtFRbXPuLV1ISBYw
ruG5Ht5WRnvits5AwOm0aqIfhkFz5/DIF2amQmBaL28BTpMaH87+KnCXaDmI
szgb443vFWkC3Kp09vFbCPMc22FOVQ4JgH0AjFS5nYyrOBbKbA36JvQvs0zP
F04rCGJ9uVSS5JV8lKQW2kSdm5rQnT/3VSqCutqKY7Ao9hDClucGOK+r9JGq
i7Js28tlROwL7iCfCURuhVr2HPtKtqwQ0OGqJNheCZSuV8A5WzRTdMUQWycq
mopALrKQ91iBiMFtg1/aZ7CHIgHy+ePlJRC4O17DRlNIFv0bD0tAbsfp5Ov/
sLFb15qdOumXl4KoA+XF/yEXmVr5BXcL4G7zjqistNhBB5dpE3VMoBh6NJpJ
QEI/FZJPxSSM00Fkp/b0q8Y4HOAvJNxTbehfFgCLQfQhxREXB7vzSWJjcJ5g
2QY0SYDolv3/yxlIWWKWGYO4tfSJS2kjyYjXhB7fAqofNiAY1k6TnXDvqY0N
BaHsaAuOMSi5njkKaXNn+p9Y6amf9/k6ylCfolyzCnxoWW3RWHC1WPAWqxIV
9VfU+VvmmBxfqI57uGWo0E2jHCZcDqI1YoNw8xOh/2l8+5iD/c1Nyf8KeAu7
gSkyNyCeSOqDOxyIYyDNMVJ3fC9Xoc3f7OMn6C7J5b2E2xYwbBTW3RqEF+Dh
YWxxryyKBFPQgaCTIp/XwZ/Z4nocg3qmHax9WOdGNLckJ7Znxcf73Ckt5E7s
eP0P8lTa0DpiCbt54gn0bbknhwwOTw56ewu3V338z2Fom0sVqVmluw2s+/RU
9pUdPEsEFuqrpKUduR0e1I36CGVDbxhGBL8Xl0hA0dudfwHKTxKFss15eNU1
sli3Gre6pJqXsUsiWf98XfaarCxFzCvaPd+pE3N5LLsCzvLiPFsgh0A6OjU9
eiUUJaAWdt6hwoaB4D8+KHrIVFnAriyLOtRuvHaFuSrapHdoubf1TM30uLfy
vZWEI/hyRb2VoKKstNco4mBp1LJwnBPGC+4WhiBXg9lh/w9qbM/z2V2MpkVB
tbAHLt8EiuulTm/Ljo1+HPrc7lJLUNEVuHun3H9nzDSmHEYnTIYeRoclWpOd
vw9fi068YwIVEn3Wyv6pLI6lebKDkl/rkYgPoKBOk7BoFqONPE2EXBocM/EC
N5wsSnY1ITDlSjjMFPVzTSsF60123v9DPsn5QHmtHXEY2xItnv4FZo0z9XwS
4x38WWUcftFnh4PIviRIL18jcGNiUvq8VTw+Dnmw7y2ZgCTwumWh7B2si2t+
6P7J6dWq7EkmvHCgF9O2kHnKsQwyCMQwKDZGlCPW6Meod72dKZnhL9uPTscw
91lcoD28qv9RUlL9PWjQX6vO8nfJgYkFWfp9zsI3+XALwXf89LL4XPeDKheo
j216E8w0PCq9NUlcfT0MZQU3lmt38RwxgB5Cr0xksFT1kwDvInqkyO9GQsSM
PvOmKu6SZ77KHmSn0hma/w6USl31R8LgTkN6FF3kg/IFO9xN2gWJz/pp1sqe
fTUC14wrDAL6chOoBOhZwvsYFSAbTaCnKjg1uDb7whO50wQhk1EHnHvdcua1
3nGX5RJqQgCNHAZpyu27mHFQe+puGOfLyZq8+iaY3Kiwo2Xr0pSU+XmVWE6P
SxJDcFVm1aOzPRMw0VSFZLyBiwPwBfDMkJ0MsmhC8c+Lp6MuWm0LMG09X9KM
UQi7xUKWQVffMZ4zJGlIeNalHvltT0nivos3NTa72eSaObgImjF4xeDGjCkE
jY440Hp+sxkZfQsWjXN8IArNXmRwgaP1YKbjrqTTO3v4h31EUyzYEZ9DgyHz
gVFF3ztmAUobKCrG8+gg66kdDXsgvCuEIuNMMHE3pVDwP+94fHAuBS+H+blv
7qtdDRq+iaIsLun3F0YiQ9uc5ClGgCawOURn6PtUOa4k6nUIOzhjxkJG7xxX
GxNr4NPVsKecPyBPG18T5A6B0Pd7r1Iy7wUEpWeLMO61Ncl8LE2U1v6tPbmn
ZfdRff5Jk2g1WtZzC+XtMgIYh4ANwj0Wu0FeMX0jL8DRT0twB8CVgFrDpxHv
srbQWaOVCjUD3AYpckGC0+scuy9FmOPdCW/JH0LU9arQU9VMjPpheAdGzZq3
v6wXChK+febN1IOoQNmi1RHU8cfQ2386xPyx30QACrwJPvZP4vsicPMlTwuf
xhYjM6+xmwQAzlAoG/tNsIFxS8Yuh93JJMYS8Iw/SBsvcFDT8F6YGsjUHvqB
Tyyjs3FWDTMQI3JdCcba9JGg2nE96d/XUwxob+i4vKpzvduHwaxWY2E+fJYV
34CWkAA9X5/fulfBteOcMiJ44VqeZugEaC1oyD4r+0H/9vAHH8cIvNgH0UMP
lUuyoaYFN6cDH1KnA1OoL5conz2FAqHtapC6RjENR42W2Oq6zyBbTD3ylpAU
JWK2RdpcymPSMEDWyg7Ty3/O7QV268+AJYZ1GCPm7OqtWY0xUaJoNqJmcUOt
4RBrkDCbkalFhOORGx1Gpq8JILd7JL4wdnr9nBC3vjCjHvQGes05jX599dzQ
6W65r9lX0Zyued3HMQgK2reoQaS1dzP1Y1tEq+Q4VIClH9xkUoZxPH9h5Jqk
CU1XeezQFmSZoWbYlT/pvw1PwEIBZV0ip61s5+qcFwiNnvj0OxEZ0o176m13
eHeEy50YCGPdh5SF106QsePxc0RMO94qUOnaOegs4mc369oJ2RB9L9NRC6Sw
s+wlen3854+NnH17BCFS8ppnkk8nYuD3HDOPeVG2b2MIswBpmZx8mns/j1rZ
s3pG7yZzOeGIEaHc7ovlZ77tAqX8qmSfHqXL4MD1f6IvJKo5NlgrQsY2FBCv
Ufino7UVZUJ0wosnfpSkrbC7fofY1fj2ZLjvUSyw/0QZZPQLl0+yO4PFs4Se
nFhjKRcaj7HLeyPTdb8cVd5fY1FQevpI3rBABtSAfAUF6h9LJgUVrmvtM87B
xcoOtJ3TBzH4dIBO83jbn6+dA5yFvlof3ilKf0JtxWCe9nFhCDhF71wikD8n
bFbOE2i6zT5TMfhKa/hzGG6CEmNBSIstvKEEbXuUHRZaUj3bQSn8RVWSArEw
GlT9LfwB3lpVK8IkIEuBycReGGzU1A2o1Tolw3l++JX2u1YEUJBJaiNfTe/1
Mh4j6St6gvcQN2tChlXd9CRxyhH9IDprnPoRqANH2wIAgRY1e6caW6hsuEAv
uTuo/7AVrpmBbVtCwbmYBXn+voiOOUbkNZL2KAoEYB0/IAyRodkA3hzSYq84
x90f6mdbVRl+T3Ou0XMdSyIn+NCBd7zQw/5dmJsXOgPwvukhxHfsJIVjfhQ2
dOfuM3XxAT7xkhigHoNea85YlYQGbntsa2HDiu01dcUI6TIt2nkCgE+4lC4Y
x5LzijLUb+Bg4m0J4b9kJnOjCCyzgycQc1CSr2LEEeKSJ3BjFvpyfeafDqot
T+WJ32FT0jyMkiMXW42h7FZJjIabgCSJcVM1Dk3M5xq5j5F/Ms81fq+S+mm6
mBebugkrXZ10kn7TysubFFk3DzIV1OkLf9YnV2MyjMoM+KqLLh7yQ6sbSy66
XOk84lBJyqSpzQ4Ay8TJnYFCJG9N/OqWsQoG0Vz7qJyEdmFM8cbGMCwArLXZ
uubkugbf841WWzG+WGPc38ly+IBrHzNPKaQ+7oG/ISea7CDWBaJe/L7qg0e3
7RG3lPErK00vnBI5SzthCArg3chA7PLvabQjm+cJK8HjJE6bs/dRG1eWl8GT
TiNfIB1IForE9Ni+vJBnQS0xgQo89fjx4W/D6+CoBTpD3131emNEjoEbdbm2
t/nu+g+ZT6jW3SRIyGDKeDKSWUMQu53L92wNgJIkY3taO9zSWxYm/3PA+MFl
I6JJiMILvyKsv5G+6Y0QDuVmZt8X9Ipn74R9Bk0ZhPAJJNVxwpBgs/XCg/yw
KaG/R75n8vs0FH9lvLbi80Ccwv5FKMbr/gfUAkmK9XZr2qk/QNtj3HEXWpvJ
QROYrFw95JIu/UBuFT/bCa+saKANFSZvDi8X/avmPPHM/RB39CaLtxmVDOwl
yOFZ3oiO2rFUxKRit6HgCTMuWmf+Ih2ruCdxN5M7SssfCzJUnGteC/s6vL52
wGHAqTT5nY+T4fnVCaCDca+0sMRAZudjKQAomt57wVJjVFZE789+OfmBCiw+
PLed5u5+fNcW+49SHLoygWM4leJ1b6XyAwWIrPTJF+dtWrDJqFn+9jXJvRiZ
PYvfwvKf4kPARkuyDJ9882cju0+3ON3AjB2M1WSzGdpxK40wq+o/fckGLmxg
woS/rvs0AVT2//Mf5yEKVO2zCFCfggL4SxnVd6nVN78oSBajk8/TNWQP7UMh
KtPPrxcPS3MGQT/yMY7h0+pg154dEoh+9VOINohKVbDRc+afUAV+WmBl3oYH
9cdhzmW6r0ICfNv+4lX6qmdF3v4PZRWI1V5NM4gHBhLblMKj+SnHbBGNRwbR
KeanqUeDDZsC/GureBcy9Vdqskdx98d18XFNc8gBTxHHPoB+LU0VVk+MQ17f
QNXUTUVQ7ompAyACdR+CIJEGnRacTwTOlf+810puk5UIOwy6JpuhdZw/b6DI
W4wn4REEsEkXeAPW0ln6RekvaQclh4P+JzgpymyUP1E1gWFY8oknSrI7N20L
R3YDroVQb9+6NDubXFWHFM9JHoJasruARidoPJGeh66mRLllp678WU0/vcx8
SCR2vP9S8IFvyzr81RDmywWzAyoElFvLaMVEFZTDTSO4ObYFgngGYN6+KuzH
d7JV0J8UG22RN7gDQDhvxfjS52FGRkTO/I4mVH5UfAmjv5nUXopEIV5uht1L
hUGIaUM5t2ZBIK9bxa2frd3Su755vHe3SkM86UznPWx/ZhaGukjGCTsuIIRm
+hwm7GmG1U+UORhWoIx/8RTKB45XEK9efe4gA8R9Uaxyk9D/SC+uD/Jjadvt
VCyZN8nYOXmQNQubv6/VE4ECjEcDbx9hKNtBuVq8TKUscNecJ4gJdZHX3ORZ
ZvBMUIAbBlgcJU9HIUl+dJcsUej3bjYbsrOenuQU0IfuLMXZ9R9w852TryQt
5jZVhGawoMiwU4DYEmI9GTtZ+B0fTpGH/VeC6xWKB8smVWJVB/UuSb6K+LQm
76N01n+YpvMnHBWEbxdwgHMWf16BzJk4oK5XDUmkI+wPnRatBIfM5zNf9CA/
vjdAuTCRR18Lu3KVdZ+cl5Wa4eihOhwHJH7cUn5ePrsxNFsa/Og3jE6IugQR
fslVr7UuCaiTejaRDkCuxiP7OmkNzQLJhc6MReQEvcE3hbIxndwLtkYrkwd4
KdvhNmKmNqRBC4io7rwINFATakakZcrZ3RerVSPIEheXyt1g7d88EsiaR7aF
L8Iq8EQKdGrQXDw4ZvLHj15v8Lt4SKX2c0Z18c4JeshxDFd0trBtwI0gt8GD
xs8yuK45+2dlgumoIDOTySIW1GYorY4W/lbxL2NQ8FfkLd6YiHNfczAdWQnC
qnws69zq0qnWNGAyPt7koAkt2RF2PDW7N0m41ZXYUBRJcteQs/XXj2VdgTro
c8NXfFje2lVbF2pieM/TgM+fne1Q04NNEiD9st9JjpEm6Yir8ZkScoIk8tta
Sc98BU4L5PLw0elzIMzlfwAxT2MViZ9SbcXm2P0YM6EJKND4IxLDGSZlhHgE
9Mtywpmnkt86ZBjuLyO34xpEyrAvL5OB4hWuhrEuBq/6zPWA9rgKHlR9qBiJ
jJfobpPjgw2wBkAhARLzBn2OdGk0i3to2E0g2Ebpl4O2L1OXVh+zqeqtdZ6J
LC27Dc7xCNCKECIxLMMj5n48b/dM9vMPnvtnw2gkqnZUPgINxttwugZCQP1Y
KXJ7CMS7OtzX+FHRtHHE0M9+Sg74iGVcKurxQGu0dP4ixK7r0+RIhChbwjnA
xJskHMdFN2yYbQKhatKSMowtXAUmzjYnk1f5NB+pqtrgHMf0EgZggNqUFhz9
fofx5M8NJr/iCBJm5vcHpLjMhXoeF9AlPG9Gj2tvKbQskidEG0wbfF1OyT3L
KrBEM0GJrF0XuXQhHVu0UIGqNtJUdkSdBhsCRzXpfeWtIDQNybXigWg743oo
2aSFcoP3SxeI71ikKDItha+dSCwwL10LSVtIp5k9dqP+54AInEyWMVZB/o16
6FREoEB0lY9YhgkMraeCQhljhUZJNONQITKhybtkowWwEWyrwSSaR3GAs4iG
EHtfKsbL6qU//zzX0mKIK602Gnf17pT4D8naunViSknwEHxycaxbZ1sDeINv
t13CV+AGZOA28+UPVVPw87j3bagwTyL/JeTEjuZZVxEWLjP9m8lcqp9QRS99
vzdr6MbUm5IZdYdmFNWjliwznDLMD3d+EABTfXcj9JyClJhYiLje/OyOo+l4
SVDzFfUeUTK4IiR3IY7TjX0PLw+0AtLBnPgG1Ae1OoiZg6SIVPV5pQs+bF8f
gar2ej5n4Ti6rDrsTZxe8DQRVRDkkK8nOu1PEhh964PMy4UTdC+0tgIOpcHx
PCV+IlyNwfv5E52jzjRQ7rP2vCMemjU+qzx4DhBn97g7fHQ8Tla4Gtt3XbDK
g7UVlB0izD5AQrYgG6HeEezAP5MQbpSI5nXof64Ivcj7Cs2asTCfdGZEcier
dc4LLutPmAdPI92TI9UGKunm+jL/B/FqmptheNNufH+cwsHMljem3vVPEecH
jwVPLB1GqBeJYo5YThM1B/t2oZ4GsBT3eG7ZA038yHOrqND1kgvLUWWjs7PA
cKCSsgaQRsEH+Eo3v+xrZsP6FvsRakKSHYXHfOt4Fm04vU+pEk2AOfHroFo0
ZlON06g6nZ60imq6CLSZr/y0q4/h+KoxsOfetqSHm6CdgBvhtMJhCtuJ+yWi
AFII/2D7ad2S5f/a1hINxq6RdPVdWJFjctYEFbZrfEC4DqA9PnjtsQShFxfq
51Oplu3KBrswfn92wufb2I/Dm1GeSEa4gAgxp0XolF2VlhosM0CPLpGBCTTR
g99PB9BoGMOGVpfD7Z10MwmpfT22G6Fnt8jXxJNsqZrHFr1ghzeuTTVI6TkC
sToLrMFnbObP3WNwGQ2SvY2g3ALHnQS9jnA953/LIicdfyT4NeObVjh+Icva
NGjPAv+8k96l+BFLdGX2D5nRtxwCsVmjNyCxeH1ccuyd5L0iByyvJpSWNHDL
vYhKnjksPkhOTSvldbs29rmcnfvi9avQTZaXAh+yMt2PByEV1kGd+GJlC2xX
x4VX9HF+xkvWra6a6ORV9508E+XBJ3yHH3s80W7o0u2C84RrmjvNP+EZXx7A
j6K/41Lu5BPOjfPOnW7LTRnmRB8XO9/dDkFCj6lneLBQKyvIeHVaA1sNaF+S
nUaDRxuUkIbBqqlqyhX7XkYqeoUdi6fElV3CGYTXM93W0088CDd80MnWWSrm
gN53LycNXXOTwHpSAdiByMV9Owr2F9mOS8h4IhN0JyzcuGw/yL3i+mcDHWwS
bu860CTQJVWn3EC0MtbBHbvpzdUDZ6HyYtmyI9V0E0bIITNjfl6Do1vU80or
c3aTPTqViJUDwnKvGUhW2GEaZ2p6OODfFSIFwFZy6g3h1G632lq5b3ZC8LIn
rV2qZPGjfoBMLEI6LDcfF7XXLNOYAdprriOEc3Ztze9wtmqq69Bdfa/rzYUi
aZtrD7y0rW3DDpbUxes9N8bNyLU2UrrsXozrGQDVTsjXEBCCvS/NrmZ57riV
s7KVJXbpPjzG9p4yv5FqMcZEQW87B9iAT1otQehZuJSzaTPj4gXadxtEdHr/
3dvfUssPI7teBCUUcEQvhnMEevbY+wn+BUej+RyrbDu34MOl3B0iIs6YL48c
+IPbR5MiL3b90Y/tEg9qTmMmm3EAmweRs/VPVqgxt9mz8AAV25Lr689oTHst
6WRTUX+ueK4zij6r85A4XAV7ST/lKyA6YxHJNuZWfBHmHTPCYhHkzH0fPBDg
ZkqvP6kgVHkq6sUko90mOD5/4AjbLD5BqxGn6+3u57OXz7GPWPnqh77acuN8
jbXtGl+aZgnyPWueOYCeNf0oYyY1nsz9jOgCxxrs+Srrx3hOwdBWT07524Hm
PB/1WAd4W3WzsaeCF8beQ2Ows47kQ/oAj7xBKFpb7pReJsqZTDXbL96htL79
+A05WaeUmHvv8kfwhMkUPgsnuOXnDqYI8oBw3Qi6nwqYjl6xxLCbjB3oGEMT
p2X7mdTJQvNTj1xagsr6HvPwVllSOjneagqjypE9hRJeNf3VHV+va8OCT6aM
fup96OdnvUNLGCub4aNOO4ujzGZYwTAUcayL1lBh46MghHxvUFF8bQrHfAvw
44frsIxzqbAMzRnG3v3NCqbSF3e3oJC2LA49H+OreF9LtHk031UZbXv0P7Ky
qI9l5qX/n6b7v7o1fDLCx217O/0jY9ECwLSfWAvpnq8Qh//JBChtL+GajLxJ
pjglX+pSzV88ssvG9LAuKp/0ebp5OlT2rr7G1qDxnUjpsvgAZPBukMDFkwyn
2+Dd0qlXJf/UGHoYhfwbVbX7tuFqYiw/MFmBVONf0Q/dBXw3SIqXZm+wBzqX
HR12FDGZO7rGn2uoPJFXBmU/OSrsJcxDleVYa5NO61IRZwf76+xMTI3fvVNt
pxtAFzBUToFpmbDPbwZzNLGHNgLg9liYq+yxT3mZRc06wRLBL2PDuJKsb2Tk
GHwksRIrobkJ2MecLc+9J+DSnbut15kFWvQYBU4xC+PTq1cJzwraqKKXmaCA
WijgXwreOgA+2eEhT9iq9k61nZRm7Blu9tp140IRa6MXbt6MNFERfW8Px/Ww
kAahDRc1+K9OUr/VPxxGn3q2D+z/nISLvpHxZJ6y1xG7t0kzYW2FwoSr0O3W
++L4mZemv3HDR7UlcAxgBnagU55+dJIDbob/L+mRWBRzAtlfSKbP5Vbzdlg6
gJ0uBPrIA/ZroIKs9ljTL4/A1QH4JAMTzAg++JF5F15eo2YIrELc2uQCeOSn
bJHBrDNsb7DibqbK/Gp6r22BNdnGjuxVp1SpmyOZlX+rL0ZfUQOXoo1Fd2yG
cWw3pHEimaSoy/wioE17AzaTZ9LWPe5JdLgWe/e+p2LDPuLrRawxphJHVlzk
S+XZFAc2eynKXdmE5GcVhyK0u5AGUAgWKE9RYcBB7KTWXpD4xpfUBKN3VMh9
amMVFizKDpk9/6LuoaACaBDO+xnDdB5RDNWa8IJte1tRYrtjTJC7F5yoHCu7
+7mWJHE4a0/5tumQvR+/WDwan4adS6kBc7vTotVr6qnWPbUXDlWPN/JVTN/k
+g7hLeqAC2YZqewyuU0oL1W0d6abCbNFbsfG3k37wdvCewdZWWGCMjIngEMq
vL/6zI6UvmHhNX5TirpOi+x0hozpof6g02+88xWaRmOeeP5fIFmCDu6e3hSX
D9uvLqRjWBJt6NLuDIYj+P/ZDKdqK9l1h1LLqt0bKzM9aXq0CZDk9/Vz20Y8
C3rqn46QsDPzfVZaHO19+9fhvAZh2uq0lUIiMI6HLp0a1iAksPs7454OFyZ1
5Cgg/Jey2IcWpM7Ln7NrP2p0D8pn+OPuD2MtS8fWbRHAuz2X5t8J/eic+ej2
jo04ZD8du/7nB3YRdmJkUUaJ7tLlCRXh7DivARaF/iMoj09S31pm9AVrLmnb
j7kLFxa0J8zO86p5gY2KCjMJiOvlUUIP3eHvogiC1cbnWqNR15H8axtCUQmY
+rpj1ks2D4rzi3FpIgatTanm2fnBYmmTzBjMtGK7ov+z1Y17RzJgnChjrJGP
BvBJAjjGtrY7oqHfoMaVbC302mpf4nDlI9hDBC42+z3G4ypGpU64hKbTM/HW
NocUcQhVQ3783ZnJIHEwJe1btM4+sIouH3XIRYrG/xhv4y2kFIXsRO5wPlv6
B6BiAwDh3EVaLTPB397GnfguosxnQlVinncPP/OjxvL1zD8G4ozRT0ImM+Qr
02KDPuZirZxz7jSfEEuWOyagMvcjHM206KQXYOXvvjF2F8xsCZBkdODht3vt
S09KpxeGntYOMx7Y5qaE9WgbJFhbh4vT41Hdfxkhx5uAHRlUYu7glDWsH/wE
pjmQXVzAHAAKzhPiffzejckc+/jjT23VdP5Y6W0aFyk+47yaFIORoJ7QYV1u
cVX8/jFfZoJeuGFQL4Zjab1VujezuRb6ndU1gWlXCdxTy0B8HBWCHSunsLNj
81g0BWaIuhLOAm738oY6SqCZhej3pqWYZy+rtsmr99ZoWguNn5mT7VGzzCv/
Xi8WLCC+EtC9aevkfBgqemLCxNQETj6uE8duhORER4auBHmnRweZQJATJfiU
acFV19h7S0bKoWiQos5/Mpg2VTgBfLXIKAC26TQmEf44VL/3GgeqJp1yYyr9
I1qw8EoJsR/xhLU2/8Pc5Do446zthu0qTW51R71lOYgYa555mjpHgVBryIWC
+XYLxIq4+j3RT4feuJus2ilpRnYDYqExfOQhH/hXO4hQhCXe7/pd4+6BNvK7
s5/73tEwLxl0xT1Ff5vQhhUwcsU2/dr8ldXtPYy8ovSKoSEauZNMcvWlWD2H
hv4DVrE4Zo4GHBfTGHDo3SgIjhdcEox0eRH+GVHiP9WCfPXAZIw7jPpvFjPp
klCB0MqinNSKGziu91PD+DDEMoftUbTulgYZrw8Xnr91ZHfGgXkrgbZWjXgC
4GQ0bw31vtU38fbDYqG2qUe2Cejh5Tns7YlyLon4WYvTHEf38E0tuH+vW+GZ
ALoCWnOP212SYsKIXtdmPl6PcoqyusAffPpAkp6kIg/B/tjv4Il4ZwpPllGg
Ckm7Bkxq+g3VyAftKubfgwXXI7O1BzIGrTw54tdftRVbc+mFSXhT7QlpCYp+
7RUpzogMbq/junFADmbOBGN2qSzRdcy3nIXMZ54eeB3bB3qn/8vWO6FoaTfC
ZNeK0nmCUH0RXZcU3W0EFfeUPE18ZetEbqfw2wSDedVOz6SlcaZ6LBf03g4r
UodePFnkqZQOvypcFpoCAygZAWLeo6AxX0kK0TeW8vQ111giQXNX6XJXyhqF
nzbPftTMgFQrJKOtek3Z76lnPRfFPP93D7DT5FVG7d3VSrNJk7WVTB+R2AnY
Daja5uwMd5ZFMEnHumrzdXyIb8vq9YdvFKDtJCjbt5q5Hp/b58lIe6kkMk3B
fy7vALXg5SvA4E86yNAZr9t3pqSpvt2ErLfj88wwilmnHshcIbjYtzEgeL0K
cuYrrvhaCVYQahovYhTFYvcaR6207B6klo625eytcGs1BRS+bFHCxnCbBlw8
jZNgVZLftwFl6mQBR6Jikcmh8tejUa1XTl9YZJom05OcnjvXlkzVhmogUc1O
TOGvNTGliIjF6+gT/v6Z/CeZFfaWAar3EhsxiQr2rQFItR4bKhYXaxLooD4k
cQ6aIxFtg+2pNEZVH6KlxZbLK81abPkMGFTrApXabz4A9m8Fqv2M4lOmfW3s
7eVbdMGNsot0hOA+iIibnN/3CjP3XORIxBc5UFHH1rEI9OWrb9FS81aQJEms
DN1tgNiwo5ysC6N8T+FQCs96nJVHZNVnFS/Y0Gs9Wrqi2FM5bCy08TzIoDU2
04GUrSh/aqm2HO0rBLVCuurxwDZA0fZuRRQGOnE1kw/OY6JmJu4JSTbOv7C7
I18AksegqI8ffkQmPxtyg+7ZrA7a08wLn5nRsjE9WK5vQ97MLsM48Gj3nNhb
iqXE6+JIk9Sn0ZPxGGhLRGM7nv8ncgIXEUtCR1TiWpLUY0G5tXvKTG2PdGTB
94gCQJA/+sAizPE9qWxyo502FI4T7XkYhlEKKAzHl8D393Y+ZDxbTrJdU4Nx
TF3mUWVApn+QPaYbgaawYcYIyCyFos7iPv0NE8HR6BhANdEi/kZ4g+JsORVi
2tYtXsrSkfVWBMpjdCY1TFUwnJF/lTUx9+CU50jtBqikjUflYkjavp/Wxgl4
EhKaU8kk39i2n7jBc51DXCWPwLGsyyIq5zK17xJqFSrbAcN3XOX918TzvhBU
i4SxMa1UeMdGVvnlpAGVls/y3abrP2Lpsxd+rUJ+Ln6ernrlNawi7PQBC3Ib
4NbL5t+064rHwxyCr+XYAQuWvLt/kg6EYY3/YedbzZmY+FXv6nAUmMpZjPYI
06/NY9NLj+zUixfQ+LCHOfstYb6vBBlN4XyU27zJ9qjoBnAD1aI/07hxJNY9
tjLPh6UMW5sCcMve2Iw/5kBZr42Xz9zBn+KQWElblU2MdQFapme744GI3wG9
kuCoU6034Cb7o2r+s/swAgdUyrxWnClH71DOtroereL+jysw71EJxiBEmytQ
KPUpW6LImXhed1JxMtFii0Shs+JKc/c86OJWk06yw7P7zpECYKxTe88nWNo2
1P0cgLArgGHQLgmpkPdB1DtV8NgmUR6Q8xhZE4Na8eI68TnBImkxT4HYDoMB
3k8Y2YDHNMl+CIs+wuvq2Rf+FZHtWzI/mdcGSUYROxrhqpVvEljfXnC5Z8XQ
/tnwbLeEUyHJcV9Jb4kdedDnDH5ODQ7KX6LnXwnFJXV8+1b1EiTM/s2wTRu9
jcsPa6gy5IIoIiLjdb12HxaIJXBiZ7sfmxnrA5Dp1hh2kA7ZzTByvsDSbw1L
oo3TuLtxB7c2eNkmkdnP1pkqpkzpzf3uHPW7urKKAlq6L5NzdSpowJAuiEGK
vlTMvDymUnP2XNvcL5RPmtZ50OHNIN7UHPGngvskWIpo/nk5JLlI3HQZdaXh
+LqV+a7KkBPKGSmnhVHryHMcY+F4KOklGzOb4dOdEREI3+hiw4Vt2glRMfYl
ZSLf0bR4zXP8LOxd+tPOfKBkMa0gxCt750Fps5LEtO/y5WhT0KQWPhlvfsWf
YzFFYsJX5pCzobC4VHyItuWEqVYTEU376WRJY7g+C+mn4u6+vGtDr23Vs1mU
R+v6+x6g+iUSGkfHp1CoDtB2JInj8D0FJgZgo3m2/Hqx5ABPkxkkbWyTIl0t
oncIYje2qhi6tqZHtqGBn3IA9fvlI62SeHQYB0VP+w+e9mOOdygHQlPrOVlf
tXRzecjj8j+LF+KAf+yZfOuo1W+Ome4E8Zb9opgIFuJonGObRDezH7CowJZD
YPTwKV/DhVd7OlnElr2aYIyLth6WCBGlGtnpKQ8Y1BusKLmzX0K4hCX1iHoH
4qvujIY85BcncDbj3HYU71brOAWeQmx4M3uULYpezkKs2tDq7ljNnBjSbyvu
/brnOd0TlzWrqtsBLnJw65ONNGjsx1R90yjBJIYOZtlX3/KN1y1JlifsGjwV
iiPTbv+Jj0fUKu+ohoFI8tWYImjvDZW22w+NH+tF/xVHCR/b7TyvgIjct23a
bPi0fa7//4cLEbQrbJ9+7hgZXfqcYqIjSYez8+/nwfZBUist5m8VP5KHzV6g
vUYewtzLrIF3/AAvBZYcvSR3cvVNq7695PW2c2sMRtcS5juvNzcznsen9CA/
psll2xbujY+fA/gtpeRJ6Bkde2Q79fHkvbl9fDZWKsSiQL0uMJUKqXxpRV5t
u7ZnpCDZTJVv/dFgUHDnFV6Uu9QukUOa7rN8YLCF1RIN9YWqZAT5wT8hOGoa
GzOHhP71O3uL7NqFhgA3Xk/LS1G8dymz9NvP8r4+yoXwl1VcMbwchfyvM+zS
6MNL614UbACcwjw/GOFt0SfpoPaTZ5ZupcK9C1rpq7nbrBDmOf9KWs0jzyqh
5BBZ5f9XUmOzO0LAhbvWVSIjh0RnA6vBnVcsWx7ovSxrOYGCBAXFSHflmVXM
RNm7l0fCbZNKOab0XoQ0VQKAcr5Rs6eoV6TwhrREsXr/YkbB0Zq5KzQ8Sl6N
ftaIjjAJ/YsEvwp3mir0GaBDL1UYAWFYTb0tcDDCjTb32iCoUVxDSESeoMq0
TszTJLmhddqWlo6jv0vf2o7HQGhWUd3/ED9+nhwzO5dd5gwrBkkGFOOTDdAg
lShLRm4mn2o03E+4z+ouPiX/skahtmNZuslXlgOlS8ew9nofGMFXRKNN/hhJ
ouRYSTsNKWClsIqybHUuzjDCZC2ptqfEhaafO6uSNsjU1ANj8d1L9fXyHMbH
hJjPaTbePT1BGwM8bEwbfT3BnWkgrtoUrsp/GHa0FfpR92TKRzYBmaNxjpM+
856KIsA9tC76pUCoJ6qieDATiSCZNW2GGdhFqCEzO5t1RRis4Y+4WJKfVF7i
Hu0u8BkgaPPKrEbOc8OP/OHoZAkLbTSQbTk12TxM4tvByOIY4dDNs50uDcdC
wqUZISaJ6l0trbybY1pCJGAfP7HezVk2KL2aoUISR1ab1HXXBgPBs1ztv781
WrEgPXNC1NHaMJdH5JLevYajUdcZ7Ywx4DLq8hpOk1sKi5lZkwC5rDyVBVjA
ywxmwa/k+U7E5XluhDNSqvgLmTQLKH5E1Y3VBqFIJ5uqyB9CPXkQqIVel23W
6h/DS9QxvS4ht0x7POhMikC9nt+4a4Of7KdhT/W3XhtdmvR2v6EjyKqAVCx+
bHpsSnfDr5D38paU5V1eVArBBukfaLb1zERkUa4FH43h3mgusnXN002cmrL4
fSg+wUFr9z5nNDB1pB+GSlY03+NiLlnDkl0YFsPwJ2iaGIKNFOBT24mvVe/F
8Wkdbvmj175DF8C+xHuFkJYmF+fIsNkTv+GD+cXO9wbPVmhr9bJpQEraQ+53
JQaqDv+fJdsjyI9K+FBkzetP4jQpeXe2o1jnnDGvq+JRi2okLyHa8aCkcK4Y
cSyQbpfZJO1AniFJO+Dx1roAtbB8maptO1CRhk+szJqD2BAkdEfKR0qAU4hz
5xOoWswPykQKfV6ApdkalimczewrZL9ZXcb5+ijFNnNdQHT0dRAnnLQBf/eW
+n4LOMm4Veu2Rb4yNmWxPOTcMkpPK6iznXpmRXSTsmKOz2qcqAQo+jM2Zllh
g7mF6xZ1h6x4QSXf3dHy7FeaHrmZgXBg62/B1hTw2oPvQ4vm4BOKTaaIeHgC
aKo9t1l1Pq38uAwBr0/a47pCpABG1uFpdlokCr6LzC/Hm0e19Aw3DxQQfrnu
4KORk3Io5hERpNWY0MoY1ZF3J9hntM1H+sA09esvAIWmvy6PY4uOrJaStjOi
vA8lplAmqnjgHw0ik6OJK4C7f9GZb6yecAoHIm44Mtzxpqn5ytx0fc8pKsjc
AUrK9LdenmthESr8ebc2fRGQq6QI6xSzf5bNhYY/NwxxPWR3J2Prsk8KUQ7t
Imex0HLvkoCNKI9T+/q6qjT8BdTmo16EnR57xiGowDDwe2ot0xalRTWqEgiW
QjmpNd4nHfco+akj1L+xJIqyf/vbvXWbyjMUSemgQT30YvXoLvwpAr3fkwA/
m3b+P30z9/IQHQbrD4+LKtd/SrGmG7bjaj4NzEXZ1xilxXfevx62HHnqsqMq
Ih63GdISWpjiew/3i48uxDQ8Ecc+fKxaac77ZQ96rIeJMCs5wENfUvzHkNiD
yuTXJATRAWMoLRME1Y9Jgn3mnr9v0x+EZhSJz1oY5YnONkCoUBYS6GZWpKAa
qHsyH+tUa1cJiI90pYXT5CTxhkKKTXF3KFD9w6X/e/fd5tz8Ds6o+YMw3dsT
z8nr05MoUazzasikJwmzzfov47GK958qbYBgGvd+YrZrJ+h8kAd7v7MXlwGU
Dvopx+F6y83ohgLkL+oCIDiEzFTMLrBjkxmfn/IKlkH51xWEP+Uslsz/2IHT
cUbyxoTlIIal9KyNVDAro9r0km/bfpxaSmE+6MBjEK2Xukyi8U7bOznWlcHr
J02Z8zJR2wu0DxuS2lwNZ3UoAPBNU5D6xC0mRWCy9LKjYpQiaaKe/BKJC5UQ
uvJ7S+UstaC+AQ4ebKc0lxgi3tn0N+5LHG7R0S7eR8ovgKHy6+51KJq53s4d
Lbg8NbBK02e1dbFec9/rLwDXEBy424JGVsEA8POje7PBQE9IMbjjCwY9Qbdv
XebNcdlDFhP6WxLBzRPZE6vSFf+mA7y/BG8q5up/0VhxPLPcG++zRzYF/tpL
KGf7IWQGC3yhnAc9U7gTaocFSazD4ysB/8sGbK3AIa492fquY5XfITsekb6A
CzHOOzpTRP9FQJ9W0OSHTKwnIxcJKbbVrKGDhjs6Q/4bshleK5HaBHiJcLgM
b5lPKEQZFyokn60Y+JA5KiCxZle2Jhd/8nFaElnKzdlKhiwr/vcin31KkojT
SR1pmNDH78PnYtpNNnUH6p14veom6wyLGMIBrng3+oQpELYd9HE+gF4n4CAU
Yit3+avGHy2F47gITyLuoAdzYE/BbhYJIPDPJ29OdipQ/IqdnW0h20ww1H2v
4k3jtEEsi0ts4h/Se2aKNMBKyQgSh22Yau5mHTUOH7MPfYYypQ1upRfEWGP6
HLjynkIxeyjaANiq/qlCNczAPJUa7NTxMyXgdiEIt16JWq6kA6DE6yYUn57e
CS+MECzqMGDe0mEyIPGCSdqXdlIcriOPRlMquTMnxyz1J36mTyMGR7VDJisG
J9JfBJGnQGogQB0zfw03jIDo31nPDKakFnNcpEn0JHVlpzv9iVzMe1CnoiF7
3WpjvaGXfZcSZDy/a2iW0Ns3nSeZ4aFmnbvpauWSOwtk9ToZNuMnWUoFD4u7
2z5kQJGkw0+SQWgkVI5RqGHwN/hn++DexbtFmbxbtd7eKZHbh0blDlPU33pN
hQPvAt9/lMFmR8eoDj5vDS4NGP3TFkuiIpN/Ll3/NNyEFBzRtH8+O5HMle01
aeFjERwtgDLC8UTTvBhUc5tSHqndwckrIIGKeeAecWwpf48alQl+Xz/3FX6Y
ioK6FXE0NEjo3P3ewiZHkvkxpxBOiAOc+3MgF9EJdwHSOV9kOeWwAwpYaX+j
+N8jf1IKvidsscjVijmnIVjMBOB07eg/L0N0/oid0bdckaw8NtXRa3W07vst
AUZ/OB337rkPlpPy9XzMQqpRa8iUiMG8jNwpDGFAyXA7/zDw99QIFF7n3p4y
CkIapXf/lR/9Byo/JnOYz9vwgCmdY5gUD0I10S9JujMg0iiyeAl3yA4Bwnms
16r3XtNo2srGP+UWnUJmEclVTcdKN0hHhjnfU3JkoO1Y5kDI96M3joxTTyVO
8rJml20VG6sybK6RbH/EwBd6hhHB2iEBAi9ChsXfbcVQ59jGjwH6SIZpQrU8
bEi8iB8QgfIqzahvE1U2QwkbslK5OhgTqeSToSoW128URaDf4DRPFIVONuYf
7VKR54R72QwyklZxM6YEvkipMjpyPEkehFejQFir85ZRmby/SZB2bba8Ai+N
Op7zm8dYwaAP2hmY74/gs+aDf7LnSv1JdyYCPVwrTY+3GBwKoo9trGc75TuR
6kMvjCDAc16rkEzWc7q1LZrDrU0vbE+mL/ug9wq+0XHOD7utLITE8oHyUjbi
xSX7qf9eBIsuDs6gJjscjbN3b1uTW/5XhUMa6IxaCKT8we9vTOM8OJatgWoq
55l0jQEWZhmFObCEvA19MrB9HQfcXDOR9EBWgpvbA78u5R8ZpjxUxazLosHJ
rpUN6xXpW8HxLQVAbQWcU1GhD1YCbYkypkSFsGBjx621GN20nKwwtQBf3Z1C
+LfAMlK6bqdzt4BJS1uiB8OXIDNw6X+U3rw4uhzCoYZznyfzyGM9XkvFz80s
7zRwB0im4FeIT8fJmuJcyZgtAm4wsrZYJE2TJkTrxuXJd6eYibZEmIU9343I
P+tORt4m4sA2nIcC3mKE46rJi2E2LMluuk71KnfObTz5LMJ/ND1IiwNeKGrQ
VEmloo9NMfuQ3nLZObeYm8Wj/fd7XQ/LU5vy+JZyQVcEOC6X7UtA2h9swR5E
p2hs7m4UuMBg2lXfHGChqwIOdo0+93PRycTKyEafH0ckTmqIeRYjgK/tQUJR
A0BxQmjatTse23whr8Ke3E8umo0L7Es+RqZYrFyjntBXXHY4VroNoiCltLMs
h0rwZ+CO5wfgoceVpDg9I3/VmsK4m7htrAJ6QRElpI/fW9hrWvcGZ8kcLUcZ
jrzCatZ9kkBQd++uhTLF0h4K2YoOVvZwZIbPxXCsoJ+FFJjtETuom/yaCmbx
0ybd+LsB0xbB3zVVdNYUFlmnMsyNg0LZBjFDiFL6pB0N8gfW1Lrx1iJMgMoM
zQnfR4VxQqHvZwb0qoRGDBZgwDQeQU1pEiRPJmp2Hj54NuJLdADWDMKGTcrk
RHf++q7YbzaHGexwOENFfKClUfTBHB8XjMr41tw1rGmndjUMyuX2YPOoHGE9
KiQK2+1ATuW6hjgCuCsTrt79RisIgSE6r/lkpWcTt9bEMcuc9CU9fs8NKfM+
rJG249/dNkORx5SkaGh0sIfTpndt3YwHmWd2/NpbkJd2Hyc7C+oXEOzHmEB1
URw2DpjbRs+w+YmntqnERm40dFbj6dd0/zZmg7kasKjkWYO2Eh/WXr61FNEr
fBFJkYMMQO8VuSNTgXz5PAhq9X/ATWGheUuhdzrJzWDLRbIqG9YBF82lm33L
syS4YMPmJngHJTDyEkB/2RArcA8gV31/FExa4DrzeB4RN4RFy234M2MfrnnA
UQgSDFCxMZFEZq+2AOC5fCn1QLvgymwf4KDr5GC900cUVX5bXqxk9A1F0X95
x7oDXoc5fcHPFjiV61plAvQzV8/JsQAgE0phOQEMJ9WT+KzDy3Cu46dorGi3
P1golrKcn2YP0ByQdyOkPhZeqqDufAq6+GypWdL1furhKX0bsRJ5UEcOP9r8
qcftsjlgYUK0eR6chiBq5UFwMpFOMa92X3lnbY5iDPK7OmS1gsZIod3TzvQP
/OwZvQCzuzMKGiDN35RfvfTkjpPxRdPJQnZ7Cs9ed7TQ9L9+0sYm+DI4/u9k
GbYxFRHufdKvK4dtLdDeK4bpIIcPGyNAQyO5aSEqiCPRY/AHzV54OCJYAODg
d/jdo1E03zxNUebj1KtcDBYxtIXLKBzPe+6XdvxvdtACpgSVRY1V6ZxJSa9r
3IpkWkCuNhuFDfJNWDGWDSKtAZqEmkSwjzr0JG/3J189mQAkD1y4f9zCd3Kn
XFU9WgZhlJ3jSae8sl/ZFmBN3WofPd4AR94ThVeguGeMm7jwIyRDUXimNXpH
i6RutOUPI+NBIu2qoBp6mSn+/c8qzJigUZzOSSBqQuEO0XdknOuMUJpF935P
kUYq1Io7MKTxnC6pbVMMLoXBORRpigcRWZMF31NRdcmNaVV5cHl8WxSKcPQo
Xf8MT/PCdm4tgSMd4xCFQ01HT/0B8xmttco2LH5w4++g4lEcN75zYoeYWTO+
sb7JcB3fJPs376U00l9uIZGbx2aIASpCcH2JCr+PzCCg3sbH/YueF0vCWW1b
qT5fb1GGUVniXeC4AdYm/2N12gyChJJZFgJbZUujcGkWi1QqJgkN3Cvq4C8S
ay01VHHJ4qaC6kfkiERgVfGPciBM5bxb4H511kg+wQwjeFzwG3bJyrLaT8Dc
nmpFa/3tMNFapYuhaXndhFhZMxNTWqkHKYswyPprutfRTQYaR6KAn8PFKZkC
RG5U7h1GMmwRLbQtCwiPA527h413X3IJq3W0wPEIQK6O4ml9IaRTwC55dHgq
ElAQJ36hxc3xxZGrfqJ1ASWh8B/Ft1sDsGVhnyQqZfbM4bBajtdMESZtA8+D
0S4CiI3hTZyOM5EtKIDOKOnbm9+gCVf6P8BTz5sn9/JcJ6dmJiif3qX4FOde
iluUHpPBOIvfyVTlSSc6D2/HZa0tY28nx/x5nbzfD5E3AcY4Van43JrVcUV3
o2zD2ELuO7sykg3zfiiUrBP9QciXrAK/3GcmbZiQTDbgu9cANKA9PewIFRWo
Wl/1yZJ7xzDiW2mV2W09BWaRWYI+V6DbAF7B+WWV3MCm5S9j8T8iOw4OclnK
fyP8O0euNJtyQ5cZ9qElC5QZki+VOP6tlLJ/EfS5KuGneuLlp6h782HChh+h
a9iprVAvYo67Zyi+ZKiq1q5ApOov3d23cy6194f6lZaxHYdLRH+gxpoEAh1q
ErI/qrpCuk2FgsMv+pr5LqpZppJDlQatq6C1duq0RZKPF/jM2nZ03THH+Eh/
qST/Avv6PY4kRq6TiJkj9YzbZKus4C84iRKHdINx15FXuc8hb5dGuqiXdmbv
4CNUkQMfSLw0CR/FSAdYPttA216Il8XXIXzW0C1M5IW/HG9eq6f7Aq2cCnhN
jCf4JvU75TejQbIxQhI2mAbjhcf6aPm6kTokJYiqZd41abvBDjA8rHg5mL1I
yemt0XNDzFUnfeIcJZcLl0ij/4/tBwKiUNNDtVP3Ko5agq0PB0q4SmYIvTDw
Z03jqTTNWlbo0EDvnTl/mjJswE1Kg8uIrtaWuZS0NLy3jVnUCj7sP/mCpmf1
9Y9HUw0lu8dJaDWCfAeSs7hLe0NyMQUyTiCj2IOBeQcjsTCBkZYQtH8ClwS0
DDfTpv8eWk30E6B2HpcEeHFkkEblmeIcwAipq0AvH2D6FntUx3niNouJGZuc
rwyreTW5ATBfS8/bq+adQ2le6iremP8+b/iDSzKtALlamYj9hQ8nPTGSfFud
7WkZ+PeTmY30PzKguKSZEM+EgNP85vl5ix65+A6K3RdbTHP3RkKvZ79bw1Zb
wr1aCDYCOvZgmkzIjXEEJrLehAa6Bu3kcXdW0SUcZUB4rfLqZ57sX4w0XxtK
1kUBTL5fXtx9Mtel7Smzy3+cBq8H+VFiHb63boJlsHDwW3hZeKi90oe4ve3Y
kB+3rDCTqSA1MFA+Q/4BwLMyM4H0zGBCwIq/AFDsRynLubyggvseL9hBOoi2
lt4Ulv2cd+jDvgjvxafHDxP8NZKowvLzOejs6DaStQoP0LLmZW7ru+8JIL3t
ZVYOlI1Y8xLQ+pmL2y+XfEHSIs8+iS4CJYcAuZlvnqnqxIi5pA+TeJ703V97
LChew3Hw42qlhW8mJiwgFAv7fcWmuJ5dOBzTiRssAMrngCpKBSM3idRtFIZf
PHQ2z8n48e/jYXX4tj4ELW2BqGgAyPhh/ssehTR2f+RsZcMaG6JwMMbU+EMD
/q+W/L/CDRvqwilWQ9cGs/3c+s3FgkbKfp7/0sKnZIn9rNDA1bEZOOZq+CPB
YWfvmyEk5eyamgayo/I2IoWoN57NB5oh0g7FyD4mqY91T2ANfv5YimPzuPei
7cGQ+ZGxt26w0uWNyp6UochxMRF1I2DiWTKuOxpUdnzD+PGquGzDKy99sLVp
e0Nw2qv5QWYvxn52kVucCM++/c0iBi9nMVKGDDV/MkkMYp/NdUamuTxaFJdA
B7jfgNlpupX46jeK6T1W0G3ZRJZfAYN43Ci+mcj0eV8xqaJVQcBogzPzGXja
hIii0xiMSEMePCB+0B+cWMuVaC9ZcgPvlav4ms6BGx2gqNm3NKITkepVILJ+
eRuvixsX2vo/iqKiUWZT0ASU26eN1ddHHahTp+l+cRZ3wbrbbRi8fh7EPyvI
8InaZJWwQf1G50qD9cbv1QaK/8+57GtL1aI0g6jNJkSO3CC5AK3dn77baY7I
VDVVsq9SICuDQY3Ahakzchaxi0QFS/7Du1Hb4/wBUwSBYUkORm6M0n3X6eDh
hodz9k8sfCK+3l7Dpsjy0hIQej0YQnVI6CxHVHxqXJq+lzMP86gL6wXZRNGj
XK5QE3i6SkPedOYAOGXz32gOJs08lEqbak30X54zKpI89yH2enJWf7dLDf7J
YblW/zXrq+gPVKw2qvEq2n+GzZjPj+jBCuSfpkc+SrkxYPJavhbiN2+Hzg4a
SMwGpOUtAJmNDvt/MoVLnxqr3LK54sjQBEIqnq4DzLywIRSe5maYUg3UUmDJ
Gkogdw2+duN8lYR1c1rs0lZQNUUZBX66N+5eg640ElV0knirRYS7VAA511gu
XWnqW0JcxjXvds4L7q36iDVRwVB2VreqdMgmtxn7ff1HZSganW2JvOuWrWmg
ziWU8vHfKsLbOAiMtcMpYSVDH9/DjHPjbb7z6yWcwkeJhQ0XbgFaZPBveJqJ
pHUuS3Wg8LmHNlmdF1fagFKvgsq5n6cfXzi3YlNjbhi6TLlxQ/ElklRomyAZ
PN/V/M41vA4Vc7KFWCuSdTOoECtUwDobJ+Oh2A9Ssnj7f8wYzZVqQBEIwyNm
/t9MZ94yTpvSKn552iYKUoMy3lwRJnT22HZ2zVzYeGZVVf6R+fbCemqGBofW
oN6IYn8MHLkMQTMtKo2UKPUBUaBHPSjLek7Ra65Zxr/mX3dSojk8bxU8eQUT
vhOaLSk3TQoDU38kXCNREQf4CC++wJM8OOtmWCDaRNMvJwj51KYD88LR1vmm
moVw6K+oK0RCTP66AT7oiVDIBL9U6Y8y+aLl76orTbtHNJxfWtQ7OLIn2yOK
OTMSeeQ4v50fQAh7xNSZafqp6ao8j0RRuijTLHYPZ1eKtuFQaEa0oqWig21W
z7NVxoPQofEP0pr4d4cJp/SMlnI2dm6gWKMRzMze3FI89ucNcNXE1hqhc03o
PTjOqC7+uVN2TygUZ244Yvxdnw3CxsjGALbchdjzacAWz2UrWHhaMIKDqvSh
UkoLYp//AxaGrBDTEvnfOQZZ6/t+QA2YcSglVR5obkaxSj10fqZ3UrE+x9H1
nkkd30s4GhkpGpOD6aFeWYb90PSUiFdMYWrj+ZZsb2BJON2sc38y5NH3L4gH
nd0aEtrpBMefoDd63qPgM0u78HtcFcIF96wpP5XuNFh4+3FG3UNXiMqxpAvG
daCgfz07IDue00onzb1trZa1O4sL+t5r9EdcpaOWeWY1VrdSM8AdnkkXwTDo
ik6I1LY1x5y50wbN+VgrsghbdNcHQzOkIChihVQI+5S/duE02UgcFuD3h7Xi
sftRg9UAB+3D3EZhNgeeJ3MC9luOQixDeiCb/qvVLHqYb9HM34Nak4Ds5Wb9
gQzEI6o6mkb5huhV6z0QnWdfZJbSUs/yRpa2bfv+Td3qEw+lu3JMLVco34bK
1PpH38qmV2clPxHyW1KAEQisj3g6a0i70neIO0Wr1IVKCeXRLIce6z6Cy4Cq
k2DyFmAZY/Rtb/JA+TpzaJ/YaA++71QuQsnW7ygceclh2tpVPak6Ii2vgxja
BumOpoubnCkZlQFxFqB3//8bs0Xq4Zw9FWSedyaxgpL8kdDwo6KnTNa3rE8/
E3H/JExMqi1YRwhc5GP1C9hEAaf5jtG1IMfvRt4bw/5OKXBCN8x8drvmEwZP
4FpefBSLngDiT//CFFrM0zY9hhKnaPhG2jROm16OeR3pYV5VOOUY+EX9yauz
pdlCiD9o8wfE7DofsORzjRhmjb1ora2He2LNwkbU0u+iVQih5Qyn2yhCIhjR
P5xw4UhfyF7w4Iw5TKn2SJ5ovOOAoYD9426+3uwtSW3kTFrLNFTKTa69uQnB
b7iC3f5Ida7HMxXcDLplByAGry6ScE1TJk6Uhzl7N+hix5GbhY+IXozRHSPy
tls6Mb2QZzj7dDPwqLXda6n4mupYJ/tpOre61N8F4TvuzOedHOj+dlKqPLmZ
DeiM9lRcxX9GLw8mKCq9Kpariy3Tra72IafUYjXqNbNVfxNYKa0BlsFknwnG
2qZ40eKJ81FurbbYaXyvV2IKYPyVH1DL9Qc/A4UCEuWFa5CINFf1ldmM3K0F
rdbkTOP2v2CLCw8ubPR71nJHjDW1C3b5aLH1uGrU0rWYJjEBj505W9dAf2q/
aYvCGZu9Hip6DbvlCEUy8/Hg4kc07We8BiyxoEwZ+StUU01G1OgxSuwTJ2hU
Bvp9B09tcYW64fd4Er8Qxhot++9iUAY3wONes+Um6bT6LG4BUVfSuSXjdrxQ
eTDiHf0H2zIRx/1RTh1Q0DRUlYR4Qi9CFBOgqOUP6cXW43q5vb6xZ70iG52I
bCMVvXdG4H7+3Kfq6Q+aI5e/0bmlJDUkhMB3/JNWP6tSZHM5HVeIPObRi5Bd
lbJLB4XsG7zgDYW+G8Z45NHe9y2V3bpp/+cCMr3QCJktv5bXPZe0zJQ1YfBK
NwykZ5LembUxz2dv4uOPtbbNFGJXLtMGt8McBMDZnVAzvek4qJpff5pXL72H
hr00YlXq9jFg8X2gNzyEEzFIlYfGe5vM/56F0kb0TxoNDJpbL/o3Dp27aANn
qA3j42d+RHePOqXKPf5XITWBtJf2pTMCOVQXULIdZEziForA66dMod20tqlu
ctm42E/eXh2w/1MNjDDY3138Na5d23uG4jAaVfCEWvoboq+wX4ZEXiIiIrfg
qJE2yYuKJw9Xd4uUaOPSXNsIPzPI0hpXcWB07hv5bk2lFSiD+QDRX67F63M4
VYsWtZAVQThnBVvNFoqxffZ8Mo2Po4ZBjykwRglllPr5nQ/ecz0g8RQBbF3o
TunN2tiu0jPSDI66VXNPtk9vCD/quRH4GT7xDnb+2GwzFJNll5joxdhb4Eg3
42FEcgngUssn7anplgJZvzPhVGk7KXjsUaWgFa03p4ujPqXAFv73SCJ4pr9l
8Y+MhcMSV/hGJ+CuUjU/5TzjMAkOwxuJ/fOXUoefwiOApsNdUPV87NJpjBxy
2Lvsbvn076r22t8EKuYYkTTi8OzhWUYyHgDbZI83oIJ9J7ieEO4ohQIq6XH5
pbbfkiv1QvOt+tqFWzqHWw7HCRw+XvzPjow3G8wbbI7qh3ltp6YooIaT1t1V
fXLw3xstgeBsFdYL/lmtEdApyMf8fIupujQylegqk8EKosYxnvpcHBzS/TM4
EeBRG6RSK/GdJ7IxO6uW/bMhk346U7fFZjeL8NVsAIePjtrEJKmw+th9CX6e
ri77NW23YuhZ6olBqOBlwSSIZpy7FWZYqqWfzdOXuQljla+W8n1cRYVpwwgN
EDqS1UKdh6okHastxyJygd6hhImAY8qcJ5qFPQTOurNpzUGzQVB8CD7i2K+g
aLwRFkyFs+GIiY0yAJ6ZSi27AQOR+YzURiCIFbaLvGDnST9+wtamcEtuRkzf
g9zipb9PfCYJo+MPOZFCRXDJx8DurUesr96GKzfESX5pCgSMTU1k7D9ZnjFV
3t9pDWUiFkcxyp4PxIjxBLHi1FigMQKAjS/XnyIRWwYsJ43YvL7N9IMxMEkz
dFGdnYNooPXpZy7itu3jRaWnMcu0ITEWiFkUAMF66OHatHIIahs1lrU65fZQ
+k2i5BL9Fy6IAYZ3JFhdwzKCJ5/N8UrWEHAq70aP5mheOaWHqm8FXl2/OBi7
NPScQytiF74+47GxHhKkhOwMcHBBRGakHwWCOzbcDRbu06iaX1wWyHdjwZJk
dnHwx50TCucF8GYQ8MLxO9VJLabeZNSgoL6x+HEE1nE8Ynl+Lqpd5AywEBrJ
N4tg3sAIpu9GB+zaEh2s8wbCsS7IZ0Hkto8/ectGPDPwnqCYjUq18gdFxhp7
rIF/u0ii++xCCe7IwHkvS2fSyd72NNslxhJd16m8Re9LV19l39oT2oyNh8Ja
rWZcyPV+5J1HOa2YFogLofbwqoDpD4vOwbc4hI4oyq8Ywa9IYLsw2Z/kZqPM
UYMdkJKpsl0S0Jj/okSwbjPH1STNy4poA4xHoxGGiR/nBkqAFuxDaXHqlkzE
SCSwKozyT8D2Msgz8mPM7kiQfIuGqjrikTeaUbJxLJh9njCoUwiS0b3RO7bE
03el2ALXPKB1dpPg7NQCUoglmJlveclspm930wh4rhoCHA2yWG+vhAtYIqdG
AlI7wF55laK8ElEt/VAuE1gBNe52WsBieGpNwKoaXpl7iyWzWuj4TS8qNPb7
MXmFb8DCw3RkmvksgS336bHQGQApUMWAGncsGFUZrQhqRhrNMh9yuFG7hJZF
0PtE3NN8WaOfIn6aYPaWb2yLfTHragtJkhnbIgFfnZ9T33JXFkrDna2/Vq14
AA5eV500XfuyNbG2/jpxixZ6C+jiULSM2nKm/HrY12tdCWl98AkwofsKrZpC
FmkajNuUL56bvO0NwTvgq5fTY6/3YQmjsMx7EmcZcrBggPb28ORw6GHUjqPy
gdOU4CZShN0IHqEpL1GwABlvNF9dtReqjV2o3z6QXNGWO19aLtek6Vj8oD3U
OtKu0y4gQusCS8hFreUmbCbtTU+hugYRhuF7YwYNL5WZ8ncULh7YObjdEZjH
zBJ3Cgtr7RCQJbm0IIsxT/FcVKmFDk1LoUH4lZPIzRlej++ybuobfdjPoS76
ZUUBkVavOepBSIagLW7MxeKcMgdgQrCoKpOmP64s4dVX/2ysixM3RGSwkVLD
d5lz0NfqRC4f7bQtlwPcgd5xjHueSz68tYmlMpmS5co6p+aFAdQPJa3jPuuL
UhryeTn2mFCA32PP1rHPKh664T3Y13xjak8IVfoOo2yOmVOHZEtWnHKievpO
hhL7ePXnbS4q6CJV3hsSND6Qp7+LBzDFe1qTsF1tNHMZfMWYlahYxJ7+yWiV
pibSfZf1Vj2lP1+7lBzAelM6cPhAG6NfiwRl1IBj3mSFW1UNGfjNgb6+95W9
+CRoEIgGMfReGSVkvQO6OuDc/p0umR/JQ1B2e5cv5k4TuAradj7smYhn3YJ8
q/iNqftNpWvZp/O/UtyWxFwBOJ50MW2SAGLsK8NwUl+2oclSfUbb9jhLAy0G
VY0ExIVp+YqVnZAxxJuDoI4HLaHeR6pMX65pxfAWjggPAtS5bHshoGk8kB/M
YxL21k+kRNisJ8t/ChgOM/C2iQoaeQZKWHOKLXs/VOLRWKADT/EbuR4Q3NNt
rMenMJGHYVJ+f0xJ1dXAjZNaJeXQvdbUwyI2MXE+8i5lANY7YmxxSBUr5/xe
mk7VNTrD6pjyCMm9EQXi5JercE0ASjT1ajpMvN8dvNzILucmdQY1PLQbSRLa
b/F+rIaPJOq59MA6bsxn21rMFUU9FwBub2ElqlsUdBFPJ4ntz8yTyD2DGGHq
86dXc5/Kvxr/DqlLG1lkq1c0W6RUzYKGhlhE8zl3XVreoict+MVHEOR+wsfj
eN5Jf+1tODHVmXbg3vT7moldCXUR/4u8q1Fzs4DUOi6e3H0HwglCmqvROt6Z
g5FIy0PgdhheMW7CJhZ4aMYfaMU/hviQzBCtEzI5+RAobTQgVBBeNFmIuEd1
Qj3gIEtHS0CG3ofcZZK03sqLgBZ8+QCRap2v/8Ipk1SKd2yDs1xaJzHRorio
PKV+a6zo49y06mzNBwIFxGNqEt/v2xDgEuFG6YjuU9Ua4XfNlnymUPNlkwmH
VLwQL1ghhg8wHk1liTlkrjCNSq/4rixOfyriADspNh2VzHsRTay7tnH6w9Ee
UE9uNpA/pYuj6C1wIMPX7eIpA95Yb0bw1jxFA+kwPso8ckuOpF5wlztAo58T
UC2giOeWVDIy3S6gIAY7kN38wbyRrKB++t1qiZH/+LMD8iWUv3c8taBoIqbM
+bC7aHSLC+MdKHkKtibGEicl5nMFJhMfpGaGdV+Vm8l3hpg0ocgqgxtahaQ4
wAc1vmcpecFVSjErWoceqPelTTFbD57zWhHebfCGyF+u7A9KDt9A1uCI09eK
pShnPIP76d403ollOzRWjnrHndjZrinMlbYhJh4V54Y1A7Q8UImUAOzBcLv0
zrIivzodbzNDZOqXKtliUY/Ozigaatg7RQVqDapb75fnsWbJyosnNTBtD5nA
dfm5CewnwgxHepL0asHuG1xJEnu9zT1ibJ1sx3wtfOzfOnxIaG1NCDAdwpXS
DDjjlil1CAc/wxGegga+bLaolawpnxhfFbxIZAFlDwyODxwMwjguT7kWvp4w
5iecOPHnKVkHm7AO0mrslN9fGG29gvvLdhHDwHsifT/KAeywpuH2jQmRtxuY
iVyLQbml0lIFkJLh2aQQSgGftnULXpPihsJnwN2xie92KF/6XRDfKZni8lYb
TkB7EuLFVu5AP2TiaBEkd0MtrgS4TEtSg6oQQRZCld4NXlkMr0bQTIHufv2L
q/oqdslCAFE0nE8bUM6NiovLS6ZuYdP/iOqS1/+tvxv3suwLf1vRJo/PfFRa
kbJS64WI4/wTk5pjrlSuvUtNtMXbQ9KjRCs7vlURDk+ciGjFIRKFzGyR7ITz
TXMOvSw9DFWtPzZWs9IUt+4GsT6MdH1CSjHK6h1lnuuVpAhEqEpKFLQXdo7e
xZwB3f2nJ7dvdn/NvvOEtWOOX+6bqg11ncv+09NxKgSW5Ovr28WKqHPtFn9W
TSV9LaCqiNTFvAW9xq5clx5JHWcgJ1+O3rkdUaJh31QFraVDHRp6tdub7IxZ
ZCHLuWGhFQm2LIyhovtk5sAlOcbaAqpBbSudBHLUh9pr6GcFnMtS1Kx0xNp5
hpYL18kzPPtVyYCw7BgnKCUXi5cR9u6mMwvbeimLp/0W0lcL9SOgXZEbmEqz
IcImHoEp5drJD0JbrYtqOrMN9XWbzLCQV8r+kkSNp13Y0we4PyqdohVemfk5
Epi1nlfCMhxD7ckoYiRt54N1e92833idAwLE3HWBty7wM2pI+h4fEtlxEUYB
MIVFb8rkl6mI+A4OaCqnqnGJ21UDO6uasszrweFbeagUVImpbsfG98lTkq58
/XA0xc42hOjRywangxVwmm7RxYZaStAUUOMQz7h7aTuIIj0ZiePkYrTupP//
y/9i3ENuldTDBQngHc+9pKHqxGP4/WsMn4fEmt6+4biQ5MpQkW2YcW1ZL53W
B3m2cOcamQIdKgSnnPUUWc9mfBz8GiALfKUqmInX+ImTwHmMnhJMVNkWG2A3
AtcGMq/vjzSVH5z3OPWHum2GNcyBN3hq9KVwiPxc9C6V7E3OUtaG4t1Oy+qq
kep12yuYMFOWkQGHmgoN+jwRBuVFH1u8HNyq8ebSnvPnwfci99AfUXNIGLao
ZQbNtQX5EPQXMUMgWZ0aaEZ8yoGNeutwuG2PytjgAwSYBVh/qCViReW4c+r0
N6cmXAYUoue1ZDoKHZ46dv0p3xU571Z/5kgy3qOQOcbd5ipS8uKN9tCB5t9+
c7dXg5dNArDb306jUcgrPK19evSgLNwM6BSO5z1mUg07YN+VZjLrYOCe8/li
kYqmnZoWAODFwcVmBngjdPoMHQpSujWqXHVnIq1bV5IF+VPk5YL++K3xLqIi
zJYdVyO6D05aqRaoP9JFGkwiZSYDyysyZYwCkvDgPIyb9TJCxaMUA1jH7BeC
uSpURerCVxkCq4qSeae59BKSgSSuNopzz/U2J0d/96x3Tb/qLmjvxt8hiuQU
cz18D7MhbQ5c+A7OmKExSA3SR8/Eu/ITTk+zpp2T/q5KSQbTzpG7P50QA3gF
TReT4wq5EzVrmiI5m74v2zs9SrS9p8dM+7Q6ZWEaJZZeELP4f/jlW/1Pb9zw
PDpFnSTBfKPgqeVJEb2vryA4jMF/J9H33ok3yBweUhVq1CEfKthaXK+V7Ciu
8gixpewC3rEjC4HH2S0bgfZA7dHUJ6ILwkOJV666IncIaxDHyBQV4kGii2UC
L3JEM/792ttgPnaq6sTGHY4HSfM2CW+cvJvfqFjnp5b6VwRgJxyumZrCZUpq
gfnuNkNCm0D4LVPsFm7TsdL1t68nSMrtF5bRG9gJGdSoFkJkgTiLzw60f49O
a77uTVdS9KrDzdbwATkXtFEF/5WKKrTFhE5J8uWmPA3JIkIljITdI+bcVb/i
rJOigluogy39KE4zm2/ZP+jBdmzGACwbju05LK9ZHDSuKd4WNSJP013Ip/Xw
57yXEECu4zdQWqDC53w5UJ11OXXHhw2rSjbzTRYx0DDokOq18OV5la+kz4mI
wgNc/KIjZQoq5ROiRcl69OjllaKRCfKfpH3JL9AsPc0/egcQjj3BriTZGX25
gynR1UTcMdT7LZllUcTP1XYxlB4Detywtbr5G/GRZfO4EL30pkDS3qH37xqv
WejjWp05oyNc7IFf2PQNrbHW7fias6L7xEPQzCsitV6Z+7sRJu3y4G0g77bo
GcvD3XrikbpVmUaRFkC6ziAidQxJLx5W6sN8P9fwUMIMM5DH4tcmWdSNtT2B
kX7ZIY6dIn4lBr5u68KvKFb34c0WezWSppB9zU3vAJ9cQvAGr9BAJej9eSzp
YBQYsoeN7dKevpNV/DNnbVe+DLNEmodhpNonhJTGTiX6dFcUq42fVKujBoil
qXCanQQVGTq1+MK1TOM9278u/YxxoeZxn2Ak0yrLY92DuYE8Qj8R8b3SM8d0
xkTQ0ahKydTwWFaO03kzibngL+dRC4UmW10NPjSLtgj0G/QOKMdjNuGb+QDB
Sddg8UgA5ybbf3DU3FrYaLIoZ3NB87f9PV/PS+fqsdvI3TvwXPJkaU/Mjfuy
fNz2veA0PbDNK6uYOTfSMalKdmRuaWNVjGACsTJP4M4H4Mdkyazltex3JvYc
4fzRcRrQI5Lo0Hhmm7Ts125tRrsbkfK2vaggcICta8dVqk8zswcoF4D5pWLW
NgR/SK8eMNCdIz6BLyQzQ0pUDxgoL+hkqSU51D0jfQMkjzDt2VhDyBvhaOoR
YXjlUPQLU6kKo4PLERf2UL9x9w5ZD6VhAZurKXhln/Rhq2nB7y+aKdvz9QiN
fot8Wfx+D0D0N5LGqjk1lQ2XcuGFXa+EpH4uNNjkoRXQSvdp6E0j19tWGZ1D
ACpK+7pPWLhbpC4GSbsb6WXk1/x/8CQoVgxtksqyl+LuOft6JLQkCGsZLwwh
/c3yc6sMCsxeZUv8eRBGsBTWkosvI1nF6H0pMykI9MGXGpi6/WnDq3QbLIJw
ufUgBFMhpsW8BIzEzTFayRqWacBj6tYtw9c3O2t56jLMh9LmXAv/W75HvUIG
1Le8EOpyLlG/AUqjxH0jLO0FwjPJz9HJX9IgM2WYalAb53G3dRvagTMCMNya
u8vhpWx6R6z62WLTaHaVOeP00+GkJEkfwUMSsKXTT5iYURjRL5Bf7hs/djX0
TPtQ0d1wrXG/FCqDlWLAickygCuPvjV1tOlOlVChsSEWIIAmuHQglG99UHAr
o4EQlkWf+7yRhwSYdlwFGJ8Lj1fze4aA5wl+ifMXUJaJMixLN381HyxJjz4G
zMFEHcETfq5vh6igN9d/dYsuOWbGKi7eNsP8XraOh/to4EQ/4pVrr+4LTbLV
ktUVaHeOO2lgX3yGAPeX0zyVupxGiTvj9gifAMgC7R1QkCD46/fGTLSzkTd/
lOeV7EwsSQPFUKErISD7XffuoJrreY8aQIy8IqwE4wzXzFgLm/HUjIWNnoLN
QC8YbZjG0s4X7HmAbN/Wb2WByjc1yIe2YcTlvPSHe0vJ2kdFa0vBlPrhiku7
3i7eEo8aMcvbNeLLY4rEaOx7oZMx4/oZWYaDSjeBAYJxAvmfifgkkAP6UdVe
HLSyr90SXUV7zYf6XSyUrKnGhh/l+uQjzKxZ2uOz9uWKFvl6nksuubd9OUUn
gzilqEAkKP68ilEVPqqvfvf+2mrGhl0eF78NAoB2zMMw+EMBe2jCqOghzr7A
+GN8PQBhE8nDf769/VUOp0WbnX0J/+D8fdAM1xkNHW0439WbZ3LB/XxkmOtu
BZ+pQ06riWea+CJrZDeJ8qiBX7Usu1XdnFd8mG4DTSIQ6wxXE4RvDustestx
DhEMeui9n0jAkblgirx4xGfkZT3WGBj/Yk4bYAIA0lsu3thCed4Kwxa1pwnT
+XJ+ritjKqRIY+UE1/LnBbIlIKZGE23VOS7IxjknB1lGGZsPQyOBDY89D1Nh
R2p7CNoeLUPCFxcTPgoXr6zBqHhSSmeRn542ctvuMjbTIUqrMLEBJK/AvDE7
SNISL9XxzKNoHna5aTSOlCLJj2/N0ucmicqGwGCnWR91JDCqxyPX31qYmT9h
moSQVM350K37IeK6y81I6y9aQzY4JDSFSCI798BjfvA2NW/M0/u2+qicP4p6
6h565URHlrffwoOZ46b1f5M/utv2TG/AadCLzQA/SZVIHDOAw1yqG7MZihki
B9p1TqQKTLzK9Xp6eq94LPfdB5Rz0teWi/x45L5+00kTR0rBzoLrwiRdEg45
stTIp4ODpsQjWN0LqXoY1ZKo7/9Fst51gc+9vw1NhCbQJ2TDZ4utNlgvtd63
SP+YqiqEN/QbRSgE97kdxPRdP8+FfosTy9TCBSStZIV4+3nIhkxBXYdg9TPV
ybxjhAHjzNVEaCy7ooCfmhs8EOv8b/TE4AFICz623qW6N/F1uX9aBogromVM
yq33GiiajNVxrvZTZGNmgfb7dbCO9iibEH0MS/IAgr61GY8CEpzYO8WzxU2R
Dsb+Tj8wpoz928sUzrz3OaxJRhTAlo/Lrzmow09n0Ioy8483jEPSpuUYV5Rg
+40ih2rxZxWra1048vz888qRBRNC6pzvr19gOj20rfkofiv1UmA7/4ZtvfIh
sgncrV/IJIBwxV/9y4teNL6FQaTQKDuqm7lSpZUiNrCMkKEi2Wk0FaVwwOl7
R9k2cJUcM503IDZNjinv/Rcl9LG4DmzDI7LNmTfiyPqRO9uOG+A0VK8S+ll2
2WXYmMn4581KWo8x4fZeV38BQl6D5t7z+725B3BBBCyKHlN//obFAK2QCQoe
6WJIjckBKDjnYHLku+nza9/IuqqpCS7JzQO4JYPORgHdSDTqkmsaEdbBxe/h
Olz9/5jsfr0nzFWo4Kkd/vXxcZ1qd86pagqhKxezo53Bu3+jUqyA/ExOEYD8
Zy17S5vtfkHic6wR//VlrkLwm/hKeWH8NXokq8DtbW6zWIoCWgv6VvKpc910
79CK1O/8rtlIqI3dK61Lt2YnWj0yr4HJRt/7PbErRt37ebyO7o19ERWyEGqY
1BZFYV39nZgDeXOSJoWsPfubBTnOHs2nmWLfJE7NuAyLdgZ2MSZaGeR4DACx
HnBj53Xe0eE+SbveQe4LXpvqThJOb3NpZoBx9k3L+Rz2ft8Sh3x685dYCzPm
m2D9jsWeP5YsXtNFtCd4goOo1hFGJV2KPCF4G8XGt4GVAGU+20eY0pFCuOX7
GyM7MuGOst9cMcRHtdDMEOOcu9x8M7Uk+8YLrFUDghODaNxxZmrE6hl4kDJj
rLNI3pwIkuQ5GWWIkaVHj36hFNtpDCWAl0noe2y31h0VTPpFqD02QO4a5jtW
BrvYoCCWwocmROVtONWH084CAu/CZbJNO6HK/x5/5GAYiinLQPFukRvwyXCe
JTc374dM1mW7YGN4RnVNT4xQKi+O0YVTjoLCD6nINv53lQNfLWORpT7M3Ua7
HBgiE1fcZCMSyK9/EjRiNle9pzRiQo3ZNaAGwvb1+2+l7WuK5bhJEz32VB02
tCnDIx1N90K9xh1CeB5KuowTAaYctJp43jK21IO9ILoopcAxYdAoXru5Q41s
UMh/zHAD+vdRhlYDsS9jNhE6bqJpTDBCGEarHkCaLxG1s6BO+SoUPGISe5KW
sjZWabEBD+daDL4o5pWb0EY+O8S3QbHl211lPtJzm5Z3Chvyqc/wyyxmGYUP
NH+1ocbkU/I0/mTf1EYc//eaYoSgM/TIpmuK99srePiSYLfN7t4IwVqfH+sk
6LhrLjYoqw+mR4mejsKxp4bugGNj73Gc3nYxDStcibNyOomcA1RASpQVAe8A
auyCIGVUPuWW2WPzz8aGzdbzweeNGQlGYOnawH+49RnSJuVBPhSwyAiJanKS
DnN3EtHAQyKeTfrn6u/g2Vc7Fp9kXRskx/f2Si6lbv3OLUofQBaIlRRAousX
M4bDU+sdRuYBjscnLT6gYm317cjWfqcKL/3SSqeARlZlSo+VJs2gHoiipa4P
9JgJNCMkn/mNUvWhminfg56IAau3cVr8lgIMA5vQiZp50+DKbskhmRx6C25o
LCkARoLLe4LiQwTGGQsaCZHWMe558txYHUFzUMvcWbIqPIARVQG9FhKkdU4c
LGkyrfc2Fc40jJyoIOFq1ubQa1Us47ycZDjRJNGxF/7FiPHBAJVFzF1LWCBb
El3KXLvtPLfv4aurYRdEfjE3X5y+m00u8H8/VpU6JA6/jHJt4ETBZzGv7Uzb
nsSyVTbWUAt+d+rxjVwIbVVyWD8mI8v6taTmPoXYjN8WF0atrlfpDktBDliP
pqh5/J0zSM07Sk3QGefghrElM9Wzr/nuugWjBOjlvYA5v3nAh+jo2AiY37JL
pB+qg5K+HDtg3meG6gFKMRG9ZSUUPKcXI4Aia+eEYneQqDypwUjCjPhSSmeg
GCeLlTEiYD1kpJYS4D7hfhaK/azTQtCX4vQF5b+qE1yVWaNuXWULdcfmPkQD
rSdTN+4sSjmctcObGBirIz1h+ZNOhJiDhJLNKuXVGk8/H9R+Aw7Fs9g+/emB
mbMv0/J7AwDqw9DCzrVVmvcnzxfgHJH+FSb91Bg6KpCNthbXsvmHB15RugTR
5hWTTGNNPmhtc0Uyy0t2MZwthti8ToytDWyoUvwskLS+8G87sxgSgI8yqfNc
3yocEFw4m+6a9KWoSalmzelNli/0um3z2vgqLqDWgdwXmfASXPAW4bXJQov5
kGDQNLqW6qANmYiCUJNO2qqDBpO8TJTbPjt8H9yhCbUqVyQ0Wv0zK6Jfo2z+
6pSHN3Eb0zZAMJeW3k/ciR2BVCWjG4lEDQKWfaWTSwHliB0doy7fPFdKu5Rl
52JCkiM2o96XoafFx6ef0HpHrqv7VnsQf/dtL4BNHWrcuc3rYaLgYzjMn66q
IH9kI5B3jknZCItNGwzNLd1OBRCgaFuZ5cdlNu8raVtQcjWvtd3UTeUGH7vf
5tsdLz4j6D2OIZIMeImJUU/TYf7Z4xEgC1NbK8S/JGYvuzjbz180rbVKCkTn
29kSoOvfn14TYy/DTIz8Wu24sr6/QJx31+WsOszAljINlgjnxWSSeFs5ktjV
EYwHFfFC/LAzahmH6Q3EX8cz9HAXlJjvd/5EYf3RIJjf6HuCfkbLHN3Eh1aA
VhS8Xd61fV8Ad+cruK0Lxbolbdg7DJE4QjVlV7lC9vBQ7n+Ann6486IfZSr7
10zq979gANTSi/2KP47gKg3qSOtaIE4tiuoaaB7j4Uwrs5+O639g4ZWtXyzN
sH1z3TakqxyErCIfi1NzJHxmSxV9DRrtfb06aFtIbC857ZlIOMz13KwCCmY0
N0B2txLR8ojLqo/z+tw9QC3CIcBke7+OkHxBG4ufEO7RgiQavqO2FzxiWnYX
S6oKY7gKELytmajUq0Nn06jydpWnxxya13b5duayDRxBkAFH1Nq8FSkZ/goW
Y5SKRH1LAZRqEo5Ax+KcYcdYw5pH6nP4fOHfQnu64BUymfKxsriI37bKmaXp
VMGMMEk7VTbsrhSJ7yF3qtbXcDic1usrh4TEKUHDwAIuos73LRr7OfvtTDiU
VZb7Ph2z3wBVT1cbtekKYuHMPmI+b/Ds6yt8PxRJfwRoLTYPApGElvwdPyi8
bHjg75JIu7x8kS9OUAckxs8nTxIWjyAClJjNtWZv5ml2dP1PHlVfEdUPcdUx
21x3PwbTCedLOc37SaZfwshEz2XYr2SpiU+lpQnwuUS0jzcg/Iwo4A9KkhBY
4AyaCg9p2uJt3cIpNWKxwWz80rYKTTVURYzvpIidDdZ1u1WS6UxnvBsC08QC
SfVzcg+xPf++AzHNl7AbP1k4dIuGDjEE9PwCvbQ3LHxzGNaqGR10CNgpbBSa
ELZH/h5LhVvtdkwKq67HEddINhFxl2Var4AYFHcwpbHQJx9ZmcL+19/qBXw3
9G0hvObOcthInt8wUgUxBCpm7G7BT6D+8FjU3bY9TDbun9B8A3KBQGFVDP1O
W18zxRzZt3klBTSU2/5uo03BAdMBOtwCFxSa/I9Z0ODinnAZ9RFNcz5m11xW
pPnqTf1cySwtDs5Sh2ldI5+hy4hRuFQvp9zeEh021f33ZES9odkf0MXlrGii
B574KjwweJdTKE82PBSDaoQvboxRmJE/9W6QwLHVDuU/YjFaIQX4VsyEA1qw
2hQZA5EK0zntV3+baLd1WxwJyxjIN1cRBlmG0hUfjL+veWg7b12LNNAP7ypZ
mrTEh960cNn8aJVPpX5NFGRmN7HD0+IJ/ZdJ7Dx/s6dCsk4g9jPtxyrdRLrd
c8BIOJXX+lWQCjlj7tbT5BMYOHhO8pjS0+uON6m3frYpNiryppiMm7hcUC/0
H87vvtsXv5kLR0AvPjaxKoRJFIgKJhhIg/GULscRlFosiNcXxLFhn5QRK/fn
I77gSMHZlCZr3w1rRvagBzzCJvAAtRNP4QnbXuaUJlWGZAhOFr/tsadmU5an
4LR2LqG8Azq30/QGT0i0Wq7uIqJj6Tjj2F+q4C6fzKZKFHuXn8BTlMF96jdu
sPKOrpncVje65mI4Lx92BPpmn6ofOYLFyfoEkif2p/YyrYHZp3W40kP+FzvF
kYkfQF7V+I0sWsCQZD6wsNZjGR5PAFJLoK4fI0nECecBzT7hc+bJgv38YEle
DozT/rFWgSjtqz69RXUG8SwE5TKh2mxaoDm9ZMav+twMJckLDL81ZomRrJ9M
md2kMVnDN3pIvUtoRKpA8RAJAuXW2ZZuU6xKTTCLPlpVSIcos0c3wJdcthWy
VLhGQAs09ojIvT7ZFRk9djPGyh7qe3XfE1fedFWX6868wPOvQQyF/4RT2hur
bVvu6ZjAxGl7Aajh3W2Rk0gwpG6X3LUDtf13DFamr9B5wXo78Hrr/F9Q4VCP
VPHj46y5AyeE6aXq3u+b+A/XvXZ551jgX4doCTvzpAyxYCgqxAAaBHKhBLRs
ppKTsSzJhNngMb35t7quIZj8P4MLlVCyr1RUeW2BmO/MFNOvwUQVKzGRXb3B
qsEScMFoZxVkNPfvcG/bwZ7ev8S3uWR2oqR5EXu7x2o70aLW6Bn2Aiw/7SsF
zitKTYzKW5fpPC6Y9rF250u+2RUwkSB1kPR3/gSqjXnzBLWNJVMYiVZjls9L
+D/bQrA2h2TVBOYW9+eYQdyo3DGVnS9Q/CnzAXzxDfShzO+I7tNwmb3tq5Ai
8VVt6bHRffa6X86A1ZI9LHjtcP1BHGKFZ5/c2v0o9Nl3o7+dq/IjQ64+wYHR
rcJyUrMIbLVvT5/JKcNpmpS6wuqa93em43kJAFPclJjqy4m1KqhR3b3HVeFs
j17/Nx5RW/mezcXC1VDouN92S2UypC0L1Iwq4jwJ+prItDv+oSA2ygL7AjgI
Oe04Q7Koum3hdCKmg0qoGWhXQ/2x9fNhPPOmerssfV2CC6TyCusg0O6urKvg
roUXou1LG/rpDSz15PajDtjgz2XSKXp0hOuTEniiNn9w5uKTEuHS43PhcWow
skULYIbghfPTrugb/fL2PAPm5yoR1XVBgWUbQI+HD10qCi1R2FoaCD/Q6xiG
RDf7xSF7xBdURSGLW24EzggjJobUwjbGDwbfpTtMa/RDNQ2v5bRjkgVuMgvB
jAl+T7greGfl0ahQ1g3IfD97sAUJhyg0x0K4vnbLZOG2DToOPpEyr5W3JszU
c/MxRdWMw5xfc4YroviU5E2t+ffzd4WLyaf3t3IvsB0wkJYlqpzag6memxkC
2keof9kcZW1eEvLTrWX0gkKd/s5PtcqdKINWJn3oirw6o8MB9uziMayC3qOh
5QAK05X7WN0xzkkLhypbsxaVwu9Nl0kivPStw/F88kMCa7PcOpss1EE1vzhu
75cW7HrUV0zhccbTQPsJW5yULcYAgGM13DLuFQNiSoWuCv04NAungtCMwfd/
YsZRbtBhN132wefIol/Sb4zgmwLRrdPT55ZAviaR0TtaXCOaYyuqm+QgEwlH
+ciyiR4tPKhijfAOZXazch4iReYAx5jFsQYz2Fl4x9f+//rOk73o6FLpwOOu
m7/3jYYULyM3qrVerXfY5RiHN/5A5sW8tdBW3Exvtb3ke8FIEcL/VawknIq2
bBlZ9dK8mu1fJVG34Swdx0idx9O/W020Z/sKEtMBMvYtqc2rINr4bzn640dg
phyvxtb+1/jT6+Arauoa0KrOdy9JERmfWuzribRu8qSmc5hhSQEirNm+rpoT
UVjvwwI2taI9FaVlxlxiNlW7osU80GAGqCMtBu3c1OqISpxu6xsbcQSf0p2B
QjXsOXVFuXYeqBzVcva0KDCQty/zPbxixgi7p2vb3EzlCCEcC5hNuMirKcz2
DWr83lHLDSUur9wAcV2yqLFBEQOVktVh0FTHB73vBDiB0Cb0ZJBXhQfi7pcP
oeKNRvGwGzvzBbXGkYzOjo/54M3VU8fR9b+f2lwtjqeEObre8QB720FcoIJZ
sMI4/KVmpKTBKBsaL3fVDOf7cUZ9D11ctFWAWFPH6YBt3PimdLZQIIJGDnRV
u9St0aHIWfgDEmtyG9pRllvFXtyR8s1dwJztNnLhPDaxW+DbNIBp/SBjkNL1
m2SGkus8IKSFVu1kpEgjn1fnFnFdx5GFjdnHna5QHlAWxIe+r2qkTb/m7u/U
g5vZpcY3mnL/kZVWc+xoaKOuxMfMHP9nXucEzc7ZdQ0DmBcHdvxeZGCG3m59
10UwagsY+LAnlXRGc86o/tp5KXQHw8rJAanZAGgF7ppaFNvZ3Khx2kHk5iKp
ObkBMlqHSbFm3S2M8GKB3s5OkBcB/l2M1hEvZ4MTsMuiAiuEi+YWR3X0W15e
HtIpuNRisBUUCIz50m3gfbDdOF6XX2r694B0hsC415c28b2qBmWUn143MIDi
h/hzx6keamUbFWWeEW66pv+9eW8XUwH9g/7dlpZI+egKWl8rJG357yCckupF
W4NyVzceigtAe3pjl05SpJDvPMOhcfoO77S2kcOmKjkVmnehonjNrRiNgzIO
PJYYI4NyPwfOen5m62GrBHla6fQWPzIWvURzyIQm3AsHJtufIAEU/vJdeIvE
5dKps9d925LDo8kiWGYXpquQpP9kdiwKgL4p2Oi1291hTE3SzhggU3eYCNB3
owL4gXxj70W/WnFAdydNXPtpVSMvMM4PVd8E51CRgxQ2/F8cHbQBDnssTJvq
0ztdwgThQ0WBj6JuC5/+K/+pkYBFhXRGOxniL20oZvHsdyh1IRtbaEiUv3Z4
J5MaVZ4m0UGfd4C8XYXxnsiq5CyLp50Yd9kGXswgGaFv/R+GXJNJC2ZewKxN
6sPNEgtm5f0/JeAzJs/MLTWxrTUVU9JyzMOCqulOd/cEnFy4tF34IAAhUCu5
jTIjW1gdkT+7abHfaDlS3I2hQXhrIjqkp0ZxO07U1YnYTB4s9wgB0u7d0NSI
RUxscz86Q/ApiKC7AfTakbF9xCTORK7RsTa/EvGcHAypfdSSeIcsN6Kx+Ud2
B80x2dL/TZ9dp9Jgc+FcuKuIKFvNVH6spazp5ta1AVuZfT8rO7WfdZsozypv
IdJBn74V/7DsOf9fRfvH/jG9k1DqYFX/xndJ25BN3u7Q+UHhcr7PEXp7koxs
pbI+be/qVRj5bK6xPLl51V2vZrVnvsGykNqCvW0gIHdmPsovPEvHf3KxjArU
8Ij0kP+3Z+gbVGmJoSSEC3R4jC9rSz7Ikh4enaWQy1humXnO0cyThzWP1DPB
6vAo8/r6qqu8PLx1QozMatdftKAVqbtHvaG8q3glbZNrSuGs5TMAl02BE/EW
37/Qabc8DHYHZ0gswv3RuMf2Z1HTvAJWL5fUqSm0FTVu6DKVglcDHyor/7vl
3dlUzq8d530PTSn+/yO+BM8lmE+aG2h3i58AwGVAxCQIW7tqii4uE4JfoQI0
SNkaCGJzJa7/budUJOU2Pn/3k6zK2U+WnbhrXv48AvM97ErIZ4eFkrqKhVt/
OmHYsZ2IEsc4UCnPI9Ex4e/AOeNNp26XJ5h85j9WerWyHkfgYdaLbkJgOXoQ
4Qhfa5fXur/K2V9gXhk17KvnwrQILrkdIU++1ThhOqtk7L3PlO/VUjhlkWMb
EALIz0L3fjhut+E5YKFgvnjaE1TpAGwO1sTi/d2cYfTTEJK2s3ZN4x97TW5P
xMFe3V78lutBaNsq80ZYb79T+IglQ8jkiGeCyC8JoXl5xp4XywzOLVVF2U8t
1NHQAKk8F8jEnaNxEpiQ+tFjVv7BaN30jsTB79VBWH2EAouxlFFM+7nEfvIL
h3kUz57K24YTboDfyBI6XCyt64Bate/bYCQDiaxVZmbnx9iXXTNm7MsBYFR6
4gPP7lxpqJRU0qGT9C3o4PD/Iitl2ZjuXfEs5JiqbfnbklFBxgCt4J/TGzoD
HsK7je9wTRsO++M3T1p0vtVY2F89MaH8W2ztcLsqgPnK+Sw8loTppxvBNhYv
FFve5IT6SRF/QZhU+zbSRLJ+VCQm/S7vQ4d7NFmvkVcqjoEfojQU4MaxxksY
4FT3CLpgigpStIL80gByQVYiUB/nlL6sSmSY7uk+IRE9iTRxg/pDlytusn/r
hjVNMxw/TrWKaJ8XqfcWfk7d3YbAiAu3UxTt6MFhey0mDah+a3E5ISksl7Dm
yR0Z4l96rq/QmzPe7tDd3BpG+9kZsmFNmI/sXnf16EJ/RhwvgaeVCaX9ep4g
nlNKxsWbbKnCthMnkeaehP7dt2hoEu9GvSp76Y1B8Aabtrzp6BRqFRkti0SH
le759AD76bZF/zDwFpt28O3Ml0FKEBJ6/wtC7Yhrb7RVuclWAsRQieaDt970
eRLshEl1KIbW4SC8rGt0Mgq8Gv2mb+8lgtp+4O8eiTBDgq7KE9g1oMacJuOY
D2WJ9gVQPMaXdnRjyeGgem5JqCFNdIpAfX4rZdE5lRpG+ukeyN3m5U8I01e7
JW88knIJiawUnr4knnF6dW4Lyo4M7ybzHGvRHRgjx7T3mNGNStnjfZ79hug9
cj7EDGrV/o5vUsCvi99LMxNs71SbRE1jD8HQBhKFz1cWRF5V4SPVfL9YBcjj
fUx7GGcEpVVZv0dvXl9kjpcVbdL6+D1NLX2YoLCIYVSa5+bYpNebIPmXBNLN
uhq0Fr45Hii9A8m4edOOyMQ3ByBRQ/J4T35ppxLJ8PC394NtYUOGtkqm0FT8
aD1PSPzhGVC61imFzaSkQmEe2mrLM6SyYeKirp/dNo6O6FlHJs2JI0yA+Lzh
ufycLvikhiW1JvMQi0vieCptq2lg5DvwFQ7KovaO76mYT1tjhDZh1VbPHDX5
8OERYw9Brb6NnRf+2yXwBG7f7TiVmD0yQfUvGwSQQIKnCn6e98cR99Pv8P0j
UP1r/4kONXhVRLMUuMZLKIjxSwLQB4BHg2AxCstq0zhoGa1WF3svaoxqfRaH
/GIqibMeml5IFH+f83XXGhd2n3iwQz30JrDb2/e781FLIirlkOQBwI71XMU7
c94ceqKpMsGf05ryoz6dJhI7Xti0t5X5a8Avi8YtedocRoVfWsfnEGGdESIR
8nbYkb9aAehql3EAFupZrqUehY6CTS6/P+mTj6OGhMBQmouJ00Zh2mwm8oWU
a144TVkPhfkFGg4TqzHXGC+rheGUeo1UH4LvsdC2raAWdZrrt92aVF76j54c
OEkpSAxdalVy2uAqBWGhsRe2rOGIC57SKl+pNgcUfwYMG2bplljaVMYEe5On
ICGtLO4j1U+MApTs76HFDMMdUcizpaWS9v5UyRo1iKQfvxEIY5kOAFrNWCJU
NIbzS+Hx+/jhCN+3CYFOHvEQlRgx861G5Q2oLTKge566MG9fmpfy1+zpd+Jj
CBxDul7anz1o/GVUAm9z60FM/NOb8/i46UFrMAgD7tDQAAmszpSdCwcpa8cu
1Cvm/fuOGeTAoSnBViJErGcafO2JBmjmmC4p3rrn3NDgWTUdqRsh7/K9Ceme
9h3V1CZD6A2hBdvAKWZ0aD0pz2bHaxUQmE5mF5BAvW0qqtRmPv5pCkOo59Av
sD+LNdV83UttMLCQhZcdsWP0YQsjNRKhRw/jOZvRKuOJJUZHKO9pB8by0rVk
KsIbb4fC8DCGXmi3jhELKUq9gvvEYC5daBjSmC77fymN+Yu15eHuU8FVSK6T
CunJW53LLqF/NJd+fO7LmhzCeJbBD/GnggdtPOO8d44MWH0HGbMz+CGbr5gP
7Aj7uj6UmhBUsblI0znlHibufl+/GALrfjT3yFbpSd1jepntbIIO/MPCBCKT
C38NhYUXFt2tTyUfhInwo6fVyf0dTOWyEHFZY9UszhIGDdsVgL19kKGeO9FY
V5jq/eOnXRPLjdjKIVCWm90NEbOatLyvwunJN23RhPOtisQQKPpR1MmQRy/r
9vUqaDc3E8ChYg5/4J2BDn1Y3MRCd3vxxyPykcaX9w0FhKAORTh81sLAoz+2
+NhrnyaBy6h7Pa+7DtAUw1CCM+dx4ssYu0cIXvQhXYzSh6hF0S1xxebuHv1U
Z74NvrAqyTq2Ea6iyg/vqondyOJru4H2lYQeiPFEd54378SKyUpaR4qPP9b5
8JfD0BqEi4Z/DloRTi5Q6ZyRcgN01Bcf9/CFN80yjjvWtuG0gSRUYfxR5u+M
T0LYGitsuTQk1rbL3YgSn8EcWLnU9BYN7RRNGreE47NlGV+bhK4AReNPy+ZR
08lqKkZdUvvpWwCm5IiauflpGj73rbFPjTcykC+NbYIspJN757Z7jAAD2krl
SVZJMLn8r7mQCXFaVat5oGoKv69ZGmbwvDBmy7seBDnnTB9tuMkQqJW1OnOt
/iqcd3VNb+EpDNZtnwhtDCbFa5PdgOEW/CGKwTZCC/gooq9me7koneHJlNNx
IxPCg/TirxehZb0kw+NGqEEiIR20hxuAFeihRzVuV+FVYgCGAm+z4M+qKPTb
66dO0Ju1JMTdF6VCuZ0nQS9H90AZ3FmUW3wCbcTFJ4qUPO+VY0DNwGQhm8p9
8rxWFy3zd059/U+ZzSH0k551ZhgnO5y005BFi9bX/EzPVJ6lr3Bs3wjJ0RoR
f9wAxRtW/sYq36uTYFRLcdRIW/SWlPjv7v+4hjFWtsMwesRqeQdjckt51Jo/
uynQGxhISdIWUl0MIXCdb1ZJkXSJxcjaHSVuR3Hq8p5BK6L5SecztSIBNvjb
LT+hT1C8dS2VkwNiTWHbuAhv3aWKAHoJXwGH4mK3v9CQxODPNCU1DUy2Urg+
jQVVOt/bonnO8URUoH8dp+csd6y2MvfT5s/E/EThurYA11JjJXsZH1doG24Z
slhHorXTWTqdG+3FW0hPD+SBKhx+xUSO0i1zk+Tlspb+BFZ0dysBlc0InjqX
VhTg5L0o0LGADKSUJEaSKCKSbuyuosegryIeze8siZS9ZMpEqbOMJiBe1a8/
6xwRQYKInp/Qhi4ATyXMxPMDhnPiQ40xqVJrnGk39avEI/0AbkTABRbf0C1E
O4vEEb8R0zzDdUKFo16HBXy5IEaabvkIQiL4yrwifm8twD2DejGnOo9fXKBq
tSlbJRCKFxFbpxxKQcm4SQQUrIvlXMWVqtsod/Oa39154iVwBVaBGypnHDRu
s4MMipxc2jeqId8Eyh2kcYOEUQl+jRWUmX56YweMCpQpWd8DD+jg4fBx4q2r
GXBGJuNZ+Zuh3uE8zoPx2pYwmXUeZs1tLTNS6ujnT3a6dwmvWeXculyytGYm
8MIno/qK/F+ISXiN8g+9x6N1JLAiioYZP9rXP9BJKNJyHKWv7GTt3p1SY+TN
Qm0oxUZRGcuh0s7wqsvHgnOwxDWGnVKfiUoYv/RgYjWrk99ZSr/T3Zy1qMjb
06CiNe8eZ4RgjWkBdgIfGcHu8cJRkxpYPbjVnQV+OhSezrrqquP3xVITitdu
W3acEc7oVXDyneUIzthGx+XU/UttBlgf21Vf9Fw8TIIlM2yi8WOuZLbUAnX7
UQtQTM6B7Kr1bdyBEDSziftdEOYl+yy8tKLQLtCidAPxOtmo0Mq2dPIr/y/O
BuiINxS5Ue5xHDMQ9F9l27GtCQcY2a7r+kKLrv2QQXZmss9XysTBEK9Xuquv
VI5iFSw2lVrLOE1Rs1/HGq76RDCAC14CupSClEmLj8+ZdTUJcefYXiYLgiO7
INMFXIVU6A2n6Rnl150OaF+G+TPkCDB3kQn0dsPVtpTSL3xFQ3/uIyyaquDo
ITfeujRKH1MxME1EtWwxeKCibjti25Oj91LC8snhRYZ+K/laXzErbZC8H7b9
j+nbqXDfXtmSEGEgj6EldNn8zduncIsF30RlwZb/qroX+5NOjn5hTdIx8PT+
nNlzEQ3r6JoGw1pQq6OYSSD+MX+xlRiQdykn7TVLHLsgxHMrKk6k0wbDIzgT
tXGAQvGkZwJ7/BjWG5M1Dqv9mUUgZ39AtL6WdTCvYh7xvS0C3e1jOJ+881Wl
IRbt391Yng2k/0J0s7AIKVmz1S47yYv9zfWoQumLxg57q62g+N6/f7eltfjH
+lQOl3MBlOB+rmTZ74cP9+AMpJc2pgG59xUhesnPbzOxmQfgRbCiwwGHdm9C
UNlxsDNRAg0Lr+OtScIX49IPOclWQZHc+G3Vf423tace92w7l1hE43mvS5f1
tbZm4vwePivP8YSrUfVRzlxfhQVicm2Ac8xR9hee5LJozn9f/hK8NXpK9TOK
RksA3AuGMomYTqxtJk/f4dbUArKYtDJbKPvqC2dZ7De1UeL9C+ZKRaJDsNZ0
jysM5E1m9IoTvx+N9rd+pqBhA81jG8x6CbKCyAKzo9anGCMtbZp7DT55zhYg
Ygym04Tgn2jqMfUu5/hWuMfOem71w+Oe+meAP0jpdaW9/4VcYTh9ylytuaHL
voCWygvLl8hSMj1zK9OE27BZB9sGBw/ZqQY6/5sVGx5ZhyPoVsSbZsE33ChB
u9vQAJaFB4J3JjP5OHWxUM4tw5XGAfFLWEL6+tuSnev0w0rsf41DLMsxenYj
q0AYi7IDS9DnmlOVR/2BTuMgYpXmHUb+J/3mlf1QvwUujzu2J+xVxspBUx+p
7nq5gkkToZRGqyrC9+ruu6EqGuWWC5Lm4fXj8RWK/ceMAVCKkF95KSPRN394
UltzyHslNc/9SoMckw4HdKRh0h/IOPwct2/Qxn8aj0E2A1IqkAiWGTbaNNpi
Q57h2G1SliURf9+lgwadUCfLr004xZMaW5R4qrMlU0amyzfjzaXF4isnQ3HY
N7lAvdYPx6L3gLuKOjam9/1f7P36hiiK9S6qn1cWEEuj/VzcpocB/QVPy5tk
8TCyPNL9EocXkH0cuCiu88cNN4SAHqKjmi5d/OdufWwOkJc8NPLiJGZOMAPm
ut63zTW6ywZOz7rgm+ubiY3HM1GU9yUxebcdasIh4daypmjmKXTworp78Xvm
hhfqW8yi/9boyCcscYuHlJ76i19Sp2XNCTS2XiPq8Jn7mFMbpwmuvAi7d26P
1QORRaOPlVbv0LVIZsdlD6X9jLDz1CE0Rudr2j2MCA4cB7S+7qKinq/xBi1n
/TtA1rCO82rHlxvxftBTOF3pq/6z2IuKhOErSUCHPdoUCitUyCvZrzDE4nR2
fdN4fqqOpr9LXO6YOHcM+VxnC58fesqvGQt3fnk5FwJiUGHhRtEsx5CwAU4W
/rLCbu6kVxzvpZu5vCAhkFoHV1VN5Ytm7/8BmJJ6PDosCcZHHvqRUvBjvQGh
ljwUNjjMmp2F1pGCFAp8k+NfbOO8u1ev975pqglmZH6Ov/IzjJvT9djmA4J7
sbGcLtWOJ9xS+nIjiOxy1z93L49jxOMPHv+iyoTubli9WKOY3VqSsMchdn1N
e41kBM5mDHEkY3n9WALE4VXW56O96fCduHieMAJHArmvIw9oZD8xAWNk8uhr
070yfB8xJ24RTEbrJniUgUCxJuOjTfpB1VjVAd3b5+p9Av26YpGN1D5FCxpM
OSedhWN+zJ0PiYyuFzs+6kZMq/740qDvuH1EbXXJq5JUtkS5k5dTs0Br23uH
F7XnaQ72motjIuRuJudKdYZr/14PbHZ+5IwgqkBakgDQrecMjGrgaa5e3r4m
GCwzC6X3kYgAzAZ6teprnRPsWijat5W+0GD5Z0DcRlm0GTzxuG//hsVG0QpU
vo42JRMrPIavzFlbSgvZChnEyzihyjJ4kXNNyGuGlI/xsb0K7FHIKaJTFHpl
Y+6e1tJkLr6nyXR2T5VGcn9tfPt77gVouGOxJnirBHWvGhg7jC/vKmC0tQ0O
LxzCH4Y//7dGZ919t7YVxGugTeWXYKzqLoMej3E3f2x0X5bvDBCujcfLr+ol
b3wovIwBrxllvt+SrH7KeEmvl95wjIE9NE65ccRA/8a4R+gDabUqPzkdHmk3
eQ1BtBwDPho90VZw8y2cckcQuTf2AJy0tdEUG/zWhuEvz0B/i4sch7oGtEux
Z6v0LNdfXHicdlyLZng2fCFDURuU8HAw0xXQfbCBJwGD0GJ4Gvp+q7fdeU2g
vJs9rPZNWXnb8zZtNQnE0+fBbqoGLzpmf6AepaDPTjmaYnH7fTdqFjAzwJoQ
ZFPOLBqaxyYIYrcO8LgzQF2momqa/16MduNTopKPZMuatqUdINfqa8hfTEyj
c469IfYkNucqFJO6FcJqjT8p9aHdOimTj4S9sgDOTKPACJNyQNg4tqZcNx/e
CbHQKfhgyyv/03PxQLjFI9VI7eJkOuAUOt3yTltNyg/ygJOruzmTXTdo6PPY
+5WDdWfuYs/1dkniPz38vytvWRLRkdn3eTcYNO9wsRpTOS6/YsiYvOANCLk2
Bx8rs1/g6d4G4CcgE8JZzkdvTTW9PsodvSQelp07wEGfuDP9bSoIzhF3FroS
UQ2oVgPrNUsqC3nhDLJz6lxDbB3+S69W0fOrtNnk5axr5W9ghK4G+bLENhI+
Lr6oDYcCDOs+oCB4JEjcw5NDmFG+fTg0ls16zj2L82cxOgQCy2kOenaHtvRc
r4xWpmOaQQmvUJY9ZscRyCVlrZCt8JDNMrfhzbtyzKcL2S5FhW0Iv3G39SLa
s7IhEc08Ltiu2EdwBQO1ebPfnfDwshHcbpcF505o/TYljp3d6KHZcdePmwtP
p/DN5yB8oAl99oypQl+k9zYvJmbKaDgKz4ozNypnwaL4R+KLFcaXsihthtWI
Z/Ox1i9viDHvIOHlaSPK3KV/vEwDscn/MxxE0UlvWOV8/ywbzTiJR80GGHFi
vffRUfNjLp/Dm89d1KCUesQXJ6EsndWmGS5G1voIAIo5hfZ6E091kDTLIu6R
538w1v4/+Mubd3f78wzObX1H8Xc22JR6Ro5/vuy7ujxIpV8JyLb3KbiURe8D
coDVCWjqoUmTeLDXZzWbpsmHQ7YozdaRGJbH6IAmXem8fR7Nf2uF6nFTSE6B
DfhdzWV7B0brq8yI1BTIa5bggHo28Mb0dW0eVJuDExJrBNbQugtKH0S583bu
TljR/QRq37gqu2Vkz6MZJtJDcwNhOnThoVXo34YRjLm1fdLsaSyd4Ew6gjs9
vGDsjVr+8PstXAOmXehG2Fbmtk1sZWSjOAwW39iz2x91h3t6HfL0jAGoOejm
JbPl2n5C5qI8f24wEDFNUp9W8abYgjnBs+X3SEdU4Z8hp3vHOEptdmpNv5VE
KXE9Ucbm4WA0clirpyDqeMeRO7tQpoHvq/ZgMD/pemoTLixCvah3JqFGPEA1
1/SLR4Jj2tvAkZIGmi0pbKN2Em/zENrktgEw67ClPuu2ZE4rl7ey/1e1N3Vo
WMVEyeTXrTR3f8Sk+IWv5+VlvzWFSWYUQ0o10rt6MKYZMUElntR9N6rd9NIM
q1APyZrr9idT8xPPqkofXKaAG6CcNM9CqMgIP2wuDsIXKWgQRXmWMaOCKoS1
+7G/RVvD5vYKWV4Z+ri34VvGvHyAyVyzhbA3QoA65AI/IIOr3vzlUinEr3id
kqnLCv4DzDjYRvGaC7QavS+VS5ac896WzjsP/7+n4OSVDe6aikRbTZywKkF6
Qu9YTNsNkCZLxZgTjw7Y0c4mul19kh4BTgUZ0uJtPI/9Q9kDCHzf3s723LLg
GOM3fcXAOuCRMLuHc/n2407P7ewrKdEiRFA6SO0XMLU0NjdL8W9QuQqnAKuN
1N4JPgs4mrEHCYZA443bP5TmqacWMdPNtoqzP+iTUYDnveFwhhGeIqQP/ND1
VSeV2EgQQhg9t52qNlIz9IMP5qQwxzqDbdhsKHbg3no4M4Pd7RWgfROnzPJh
iW3BqN18WnKXUJJRZMKjyW05XCedd6FjzHchVVKxqCiH2VGZKOerQgpLF1bn
4g1RZNf/3PQfn2x4fGQ2CTQACDU8S84hzyeTeZ0myiyY2vueqDd072LrVV5m
pmruiWqnRsAvN9vBHygl197JtIqOJFgOdHgo1n/hJ3xWIw9k2knT4jVhlHDr
iWXphWEp37F17GBxObwuIanskJGreA2o0OjGcPFyCQTNMgjXYOjUpOrnpIM0
eMIGCULrVRZHOFXSisyoi5SmCE/qY2VZC4zd3JAQGpkPf12smqGo+XQHnpjv
8X2l7rYIqPAQmGB7yE2JlAmjrqaNtf7du2kKtfbXSB+h7e2F/g5KHeMn9H3V
VtZLLRNorDB9YkLRK8/dHQ5ve7J6w6URKC5bflDb6UeS0b24T9U5GjRxHFLc
j2qT69Pa8axTxE48tgRkr606IzZX99GltxK2X0STHFEeGZNcEUFSitXAMViL
oV5XR8N4v+LkOLkPgl7tQJDrF6r2PO729kcErcUnybeDshreaJLzXW6rc6yB
3JeFRxqAQCp/Bu+/YbUIVgXmH4seRVMXEAz6/DpIyh/4KBJfVunv6CLipzSj
qJN5uQzCZI+Ga6PNGAb9QRkccWKWjZviqP/2r9tQdzNsMknyxWjkBevYo2PG
dysinrvOCuD24LM/f3UPBI9gwDusQo8xZD0Cx0TTgK/CN8gpH3psM2JS/aG7
9E6p4hfrDzv9LcJSB9PHTyy/laCQZWKUdcMqrP8EKofM6DGVOkZ3325VSxQD
BIxK7mnUvQZtG0HEaOcTILytVbazrukK5p6XRbY3rJCmmHuBnmEpddHvvK3G
q4sn2C3Jvab21uRocvXlgWb2DtuA4fW/BC71q1Vbu2hFuNAwh59otJgl7qZN
CXX7AYmRwIibE9v84SEhw4vzIQgYCAmpmom8RPPGjbykj37b1/MhjiGgIolr
1EWaNbkp2/XGhCaxJTSKRmqL0xfoCwWPe2+BbrFIutd7jTH8tJ/uAhvX0Fpa
qval7FIqjj4IN+xpCsWRzIPUhYWl0dpIbsoXJJdXFAZ/iUd12q1sXlVtWM3Y
j6yWEWaD+9ZzVlXPmqDSLcdG0Ra/ChueMZFXgX4ki0AJHdjwOMnL0Za13+nt
bDrZnUdbUh38dif/dNtcY0RkbVx6ee2dWgs8pHK31WNAUmZsOQ/CpGIJq3DN
uabo3zcnY1h1XGKmuBLUItKHtgJQNHXhF9+h84FORgvWa3qXjPHULlVz6cP8
QnQ3kIuT9auFTQxGq7J9zVxGUeXb7aEyjKtV05GbKdMOY7mNYkOzjJt+D2W/
3hF2BTsewE/Q6HZeorGeswFjQu6qzFmQEIdbYaWAc0+WtVx6XPLlf2iBibeY
YsUY7L3R7Pi1p6juAo0jYRoC1y4Y3eWN4H7XNC9SwICR8nJhFsqFZgDYG3rk
gvzo5AoG3uo3hsmp3XglFRaQ4xI3lMEVefJZkMgMsTlp5IwslOdfQhGLM0Sk
cSL606nXGxnQQ06WH4SJLsMcPYCRkmHa9DFOIxiCbiS/xfKooIc0gvybYMiN
qvUIYK5kSqxVzwWY3989405otzFm61CjSkXyM1Ggjs4yWAu57SVhmnOsPOvd
n9sJy5JwhWmQc2ZF7x3raBV8bnx4WkDzqhRB5TTx1F84UrwtuH28feT2fMXt
xB4yFw+C4srrsxKf2hrjvk35KLULB3lPczuCDorhqqr+vcQaKVdZHdfitwJu
9ebnpKKhFdhCFGcb6VAVaopsgTz76Aw3ISk596OKjNMTRcUwaqq3ybSdH1S8
a+0SBxwkEBa3kAG1gXACyPM6wnA6cIHuL7gN+JUGW43My6Sbn75MnY9AuRJG
XHRp/2he/t3P/SMNAcvCXGL7vN4xedvxz+3oQKsZyH1ZtzaqSfT3oY9TjKWl
H0ToY8zxjzIWeHht/rLdqaz4FdXy2QvEM+CXbn29X9dfdQjjOYBVxwtebA0f
8v/UJG1ONlFd8oKJj9r9FkcwivjvyV28fp1m9VEC2+xyy1OFtJLgm78e6zPE
uoZ5s6cgu/sVzs7/x1z1zb+8rlnngBDXa6iltZmcQEf0x6aePRJkQwBWTFNw
0Njn7Q0RvY4ZWW/AI6nzQaTSEANfXu4KnUnALf4/ox50U5GJ0BJ4iWDJZDdr
7odk0HCAJpw1m86T5sCxEwnxY7GNbbwnMv1I55I45f9v5Tisib3z4AF4c+rH
YAZ7Iy4mNKZQV8RBlI18KY6Aj3pgTmat+qBSQSLFBmiGQsUN/oVbXpGcfKxQ
quyhQAbfi0O9pTUvjHkLC4mCrdnDrvkC0C5XYkpF8squxYVkdfZH73iLvl30
eB6P1X12EhP6NtfvnA41QIhc0aHLS7mOf6Ki3gwOKiRJKutoiZjJ7XJfzqOQ
bGo3j0N0ecaz+ahl8/u2L9mr5AUOQp9tjmSCq44BgN6pEA5dGzPpob7LgvdV
NyLk8maihnp5RYq3xDEjEARrmvHcFnV/YJ7RXZESyZh828UHUNtW+tjSaSJ3
Xq113kxJRQd90ayJD9/9AanB4vTPT00rDonxXd+3yj+Z0oIfZPhgmzo9n0YK
7JQAoAYYnMJa9aKjzMMm9ASJMlbWLJBhfSsVYacNTocOY60Szfg8hvpbfq9F
R9+bzK7XTHPb4JsVxxpraKJbJWlx/vUTwbtd8GiFRDeN1fUOX8Sxp4MjVreM
C+Gmo/suSiE1xOrZRGvuXFhTzIaJ726z1gr4Jlgm8yHlMzu6jHdPn9JCTEZI
Po97G7gWhZCN1WILFOBr0APct1a2JmShdaqLfWC0FLOs/GPwZjx5CwojByfi
GioDLXDSGZPeKDLTWG5z9ekdPucpblDcG1rY/sYzBUJf3zfkumti1DDSyeyp
v6GbPiGgS1mPlFr+6vlEkCHS1Je9P3QZke2N51rwOXJduJk8Ydbt8Xtvi2D6
SLstySK3MRfXdW4mTZD7z0/6j0J5pm3epzvaqD9Fjqz+8jTjtB3HLH00waPu
0eFAk00W+VhEVdm0gadzZHpFWQjw569Hzbi1L37BwJltZcw87D6Q4qjyc50U
uuqPblNk52TwhQd+WQd4DW/bUWUX3WKYVT/vtVdmCe/f28GkRL4OI9U/wbKM
7fBCyJIoQ3x62TsD2NHwRNTUbLrSVw6ZnYFaXwE7hr1wDXBRKV8PeOfaL23G
8cceKZMTSxVklNH9K8FnNLXveefEOtJuD9H333dAA6zxzmytHPzfJRNWu+yd
DYbrbK+tY1H6CZ+Z1ywh90//vR0hSdNbnYt1+SMebFF52HcQHDxYzysulVWR
WffqGEx1sn49x5H48G6ugk4WR1LRg9WXllE1f1P1v2h4YRfyseMe3zGAzRTi
oL2axHtc+acsfPNCGHvbgqaAiSPJC76nz6EdmwMMW0Y4XUpt/mAQEbNjT6vQ
Bi3hNAaVYlPv0bp7NvsVFiztLCR2SvPWf4jSHph8Tp6BLuc6nl5MaJqZld4W
UJkAamLugohSDp2alONE68ymGyCm1SaGAq9+mYMPNg64k3JYnHbyUR0dR3Nt
EmqtRZUlZpJN+ojpcgWx7XJO56+/SFxV2uuDDlEcFFqUeM25HmZyPgtruaM/
2JGD82gU8YvpGgomymeOstMeGMzlMCAItdP90aVWib6Fw/vHDj3FEcr71rJm
wPzsTjVtHauMuAxqdlm/vE5UT8WyB5AKGlriNmF/wyFa9nhbuiX6E9IiA6fJ
mwJbun7OCurj556uA96U7e5a+4sTaNwILTn9JCRk8+P0Z+8Rh5UBzAbrxor2
xveoednjqM95OOtYS78rJ1oINT1nKYz2KvxEVJLFf8YpeZzFtLKKY6gF4nc0
tieiTG3p5b7QsFEeqtx200DlgKsWa4q7tvL44sQLt1CxDt56UfQ0uKYWWQ+o
1JQRoBqx3Tbd+mwrvT3YAt9pvW0z3E5mdk+oWm05jscG7HnzI/oklGvGq40+
5MjnMaqbvSTmbLgdvQbYYqPAtJFCjDmqrTQTcCtTB2jQxymqEKnbOJf8Y9ly
O3ZSuvQXs7D491ERNh+Pl0tZ9Lmy55+rdZGVKK6Xyekg78uPMtASl9MuqeqI
M/I3JsLuon9v4k61oTGdGEhKjkO92m+g6skOa8Bbr5u219Jb9brnkIK5BA/s
RqlgozZWvrKy22HoYf5m6VddRyX10aPOC6rJv2QTAq5TY2UCDYczYxIvEwQ6
s+kQ/6pP6D7A9Cf7JUPo/XTNu3eN4IPLTPsAWhyn/2R2LiNcGBljWCTDUB8M
akH3PSNTEu5f+KFTQ2hVPbyIRhzWr0d6d29DLHRNLJUcccW2QXM/ta52IXeb
mc+V4Fxkpz9P2QtZyrvIfV4ZkL5lp2GFT7SOquKCERo89frMb6uRw7y0dBBh
+RfK+YrwnkW7+sXgYmGnaEjeIg749j3ELySJDCelQiqozukWiLJWCu6OjRtH
ZTAosLdkvZXpXyTHSVYLLg4AO+l8AAXvxiQgseO5dwCBkH73eS2Y1wIpKh2F
SJe4lA8AhcfVC0YqMJb9vazlKq0gb7EZdfGDRb1GlsViaFBVEvaNLokfJkOa
Q8NCyamixcOiYCSk2UxCt7u9O96LKKj1fz8Yq+wmaLKb3Zxrv5Xte3AboGJN
6+RqdlSuDxhomQhRpmiNTS81lPA+DdGAZdXI4wr2BwTN+wSAVYSJ2rvPUquI
9WdQPthgchepZ3PRMhOoorRuc80rdRMFofkitSEO6xa8sPA2MfCQnrZS10H8
nYBj5v3Vb5Dj2Xu0BUvEzwO67INkqdDlZXig2GT8BOVeL7B2zFrmy00yOYPD
ztuJMbnfs8qlD2A5bhxZ9f8Mps/J7+d0RtnFEb3XSdRMzUZde2jQ/6j86p1b
iDkWnUibhphgaCU5xS9mETBh6/QKC0enPCxuBC+wCeUkL2clWmB79aItBUUz
1cUgH0P5j24x1xEB8qWPagr0jyv2RW54qi/B2EnnNFCSOMIwZo5fG9pmsB40
5xR5WutAhhWSDLGt1rMaUjbhdsCY79fxzXhcf0SzRRSYxFZ9ywhptSmlleZm
vGLn2GgByOqW1AvXXB830j4pQCvAB5qTmO8FxZKegPtcP0hDJmA9ExQjO9bM
Y1DLtscmpIU59sonjq+mM7DTUF6oxdCUb76RVwUdBCZlwnu0cHGa1RKQqb71
u0BE5h3NdV/tCG4kdCoKsT4AJuMSy5SgCC1GmQGV0OyJEoFeG6DtpECOQcBB
P0AfNUm3SQNsz/E3hcU4luz0RXRhISfxr6nDPVsoKw5WwITaUIlTpBJ+f8j3
xkT2b7I/Mjr1E51P7PVbCIqMRka3Thbk95w/D8BTwUrrsjzz/UPBpmUuLOn7
p/sRvRzQuo84TIVOkb1SqKK3RCbejoDabDfxQ6yNV0UEokjmIXkG1T+iTmfH
uPjGpD8JhYFp4E3Y++E1OvhOLS85qyWuIB+BiYUADm2R/6NpnK7ozmDIzskQ
SF/WJdEjHTbldUgGWTI3paJDhsA2XMMYk1qyRvFBduohZAoEL55VHxHratDi
lrPtI5/WnR8ZihkmpO3kOIgA+hnRgsn3sFWn9Spfmte+lqeqkleJ2OulnljO
69mhcStR3+s90viG6e6Bh6Bhl1+ft+b6ovA5F53LwvCjYR+Cp6IBsCEbMTfP
hByFt4bD2reayjXzliLveAzSmHlAGfw6Ny5IsBbyARUQ7DMk7ndUqAqkGcyQ
hhqpt1EoqflpWPol11izJhHeyBrzqVFPdx1aX393wE7VveL2q9kipSvPZESC
4FACYhbnfWHWu2WRM/sTP6OQIDned2ok0xZmLTpGBq69WgOnILBmMX/KnVjW
i9E9oSIzpC8GqDgLQgzkZdV5Mc/JEyHp36mzGellWcbbXlgHavQo1Hk21ToX
QEM+E9ij5bZwqRfuMKtKThdcX/r/EzXXsmUTl+FJzCLkGd7YhEBVICVINwcb
G+n4I+nmUsUokwyvGoHDClK9G11WkRcnmBtHx1R8Ifrm5faiJCu69xjnU9LZ
69vJoI5axf0EwiY5HIebfwAqpPVQbS8aa+TUUBSPkObtY11Vj0ZZ8DSRVBRP
irHnL6RmlY01MHHaQkh2Yla5l9n6bi/uDFSlRMOH0mxpJlvIPmech2+2UK7F
yJ887sjAPS6yEjjxizNLtajoa3ARXmNlTUktcEMdKUkhUp1wnedfdcCYd+YU
f4NXO4wJIW+DycnjNRDxuRZ8PaAXBnYNoni7zL5trU5wsaiWv3eA6fn9UxxX
wObSCWpMMnLjLMLk/mZSw3Gx9lCp/9gv73Tgf8lAQTTygXLvVa8S//OGdDhi
KjfhinG9PB45c7zzId7gmma86++JpB3W17i+QDmr3qeBtjAtOI3rqxmZrhY1
3aDcNNqGyR24Qg1Zf5z6YAfqCRZk1RQbUUIT6mzyedNfsBE37X8d/OOeDdR1
TJRlNW+xiaecmnvQEkIm85Xgmcsbr5aRfw67xC3R0XXLCqT7zin2DFQJjLMP
gPk11bsLCMdt7KGqKnES35E3oiX/cuQ/PmQydMohBn0CuxnmicP5B8nnPBdE
C1jJ0cp4IzQleN/11RHmSDt5g0kTB2WZ4NWJR8eWe/4yXLeucx2/VqdB6Qc7
qJRnUb1+Rk4dG7CM5DV1b/PwW2CUaelGD+K2JFbjdnucvFXDT0kDRrz5qhb0
moGRujgplsNkHqz13ru7ZgQid97abvHpthFi6x5w5fOTkBK1mmRCUCdi4LlE
JJqVUL7ambdp1BwUdBQJ8TxiqPwt6sS1m3TLr2q7nc1DTBRbnQ0yhpP9MmCh
D6xPpcm+5bIeLpeE/1jsGPyKiaSoTre9cyeeMLLJocaJRQYQOf8BeAovOPJg
xtIYc1Y2nAP4/bhPZ+qjFVlh+2uH/1LzOtJjWo6mBfEYnWoh0ksmosD3QAM+
Y92N7NAt/8aM4UV7/xYyl/OxwEDE2Q0YcjHYbHla6VDQyo/8wtC6qG+jvVgQ
+F79O+UnpoEHRuA9r565OPPjHvjPRPQHL/s4ePMhsVM5ItrzDIJN0xw2LMiV
JOivpO1mF7G3CrbdS3MDMhK/6wI63Wm1zF8MPWAHGqPZdhTsGf8nlYU9CiI/
Yt+Ezc1o/Za3N0dtqN9rcwbM3LXM9RlImrd6/Q8jpMZsXlMSJCUQ+JjuE+71
3WXcOEa6nhXgZD89LnKqjLghjcYnXUvjPP6yxwZhY/ATXD3rZk8jZHmj5YyL
FO7pkkXSdb19mFc2CGdS+hilJkjRLDp0Z8+lTND8kApES7iKa0Xz5cKObEoS
3ith6p3LWd6QhrCbgsnulnAq8g2BfODP+Bpnt1XLZyLtJz/I5lOUsMdYYhl0
wCd/IiTRU89ysVOfbZe6lQXAjoHh1DipuToSyVAeXkjn3CTKv5fkrdeSu9fe
JI9u0hT1P/9Io0LKuu/HMJMLhMKa2k/QGnU1doPHXEl0NF0fy3izJv1dJ8Mo
yFu6X/ujp8r7bd7KJi/QTvuFbtkXpUqWmCHihrZLMNrjyGUNt8y0mmzPrxxQ
pijeIhJ9nHN5LJNC8uASy5uDh2kDMHzLQA5+4hKr6ASYqhXKiYIC9x3vQuyR
tsAiTwcwhN/gTAWPBY4nXSVYQIF8wezqH2ugqtgAQZBWn7ycnTeuzWsWxp4M
MyYcc3ryimK126dB4HvNN4GPfO2TZ/fFn56WJGxYWdub5Lr5k1mW0csSD+Ym
c+g6FDkrQLqVTYF/HwcNASXFOghzIYMcpoKJto8cHmaehwXYA1Ra+Sgk0NV3
AO0ffnblh1tuRpMu7w+3Z45tmeNEBPy1CPMaxU2g9D57g2jUuHRPh8Sfdt3p
tGBD+eLXoYn/URXicO/ZCLodLk1+qOrqTFynoUGl8ebfNwJjs+vF/M6WC52B
MXuD0BJGreenhiTlSusFehpEnW2P/tRIbgy1xffR/SopWMjoSJOkYxvAkmRz
LcV/DXwi46dHrgAoeElVPxEqr2xkvIEXtyC5F+YEUEI/vQCKgt4h7a8+aWpo
dyJEIDqN7GvIz0l2BISw8LzO8OA1tvEdRxuew7bSmfb8KmQ0dqzWxFHHodq4
HnwQHAlOe0LzcnsyHvO4Gnxu6WL6ZJ0oWWlruK9fLGP8rcClflOC9LF7oWGT
Og0tw1rATGMTe4WBVhjE16CRJRMwelWttfPI8hrjjYvsnJ9d/1JKJ9DyujcL
hZ/mMwIcLEE9/9leLZNGZOxiPtY5rCSh5g9oydz/t0WvFAk6W1XO9PcHK6SJ
vYcpb1E5NiOPfaDihPSPm8wST54JOjhrz5UXULFvPiZ4hnUszgewsGsl2si+
MSIQKSGaiREmfDpcwC925m4CHlAWnfxlblwoLFO96OaDKglcKkVZKeof59Au
gIylG1AWO978/s5kzLlkqjEssgdKJgqbzYefCEl8GAPosHeydr01z08Rz/ZA
VOQIVXCE45mqcdGrowWhBlGMgMrXnWipzo8aTF/YCd92FfxUhUJ4/IWLLMh+
KLAyMzFWzyl1sG4Y5tK2N0s8oD5jwUTaYMdqfMdr5Por6hiF0ITw2YjNl/hq
r3hm94IsNRMnrmzCQu0IxwXbqgS0rO99rEUzkw0n1RLKqTKyzP/cIcbDaoev
SglgmB5mcoT9Up2bo9rrDtZLnwiCmCcixbQZnS6aTzmu7INTmStoZd1RfnI1
fnBAechunfHGGLMFR0XEKDH9ibgsRWGXPh++OHo3886hamDvwzEtwK8rS938
77QF3P9TDHaDVCu7cV9yFI4WyAAHXZHyT3DiU/D+QXI7WQ6IFtbf+AeuGH38
NMSiodaKRLSitHqa8RJTLBzFz/I7vUDjFKKk7uQzLGdF9iravi44KmjOd2q/
yNaZqF9gN7yxcLJMQEuX1gcv0dD2STZBumZuv7L3u3mCs+BHgonA8xiFiGMQ
L/bAuDbbOt45uhXHN0JFKV4s9nQwc74kJu2tvC7DP3IrJkXvaW5U5fAchdmc
m/pKuzZhB3BntiTx6EamvvTSdRWlR7sZLwO/NrzuVNmZjIPYqyc6uZZjKL6E
56L/SFINbdTqZ5T2wii1uGRtbHQqfGkDKxqgB4AMuJxvHxgRbZ0aQ1UelB3V
b9Gl8naQXVOjUif3jZRJBseQmlKjSsv0iH4P/Lpuxvz+ipnDGLUOoozdoRPy
ep/g0MEXAUX3rFtgQJjkiR4f7N8AeQhokEwBDTCxL6UTR9u7XXQpMmpFQT0e
UiycZo3Udb3a5AEETs3nDVYNAWsSrmN5WB3x2BcAyyMrs/7p8IM759Ug5OPF
qQVoTUqdf/3Kjs2kbrXnLZqscGkxnASVxlhXk1lIXuS3ymrj8Kq3iwwwl6UR
tKjGigugpf2DY13sOU61VBThS9IOUK7Sv2bxzppz58PzbaRm4cq2iCkwoxJ9
+rZtJXzT1/aR6nlO6bOcpp9zYSTufc5LVec9ru96Ws40iPMuRe1vq6xJNYoH
29Ya8FLMBsyw+ibeIz3V/4GaZT8g2MorrKkEIYRoyDtg9CPqTOuioUiOqPIF
NuO5AHw15Me2FtQNhD6pP+VIEMx5iub2A6YdvUhgiWF1WM0IhHaIeLzdSSqD
NrxQW6CetB+eoBtnDBSrX/eZqxgwIq/QhoClrIz5kTZhh6MWijBrk+8QWDkn
jmz+36q09OXOxr64wCEk3JN4JOiG9zzZvAqkXldhurn0Q84sIG7WEGBvMLVi
QwtjMZGciqOlqrnRpPqaxQTkXiSU8cmTDHoZLB848aWQQ3k6fsNNN3NACnAD
zqbucWV8geLzIgltkh00BlFPNX1Dhayi0Z4CB0s3L+AqsdpSAiRufuz7y/Du
9qpaD9N44BqS1P0O4pH/TI8Ve+PRgQ1uBgVfGhJYEgmzb4bwfMvt/C4hIrSH
d+ngp7pj3vhrmS5zAoy1Hw5kGXKxHsh4L95LOW8xlNIvawRg5TVAoQ80v3hv
HSAtux30CiYJh5wlMta1eDG/apGjkId+kgAqd2jJe4aIPJWDtTVt8/C6gaaG
JF9w/mnO/Neu80vRD6ceeuuhwBpUdFhJ6HS+VvpLeJpPOoiGGlKZRn7s6FIY
v5F54bu1+lqUksP7PcbkjBqVOyLRuzPY0RL7uAUgbuI5iqh8qBqrFpHPusFN
cJE8CYL1TYw2erLXz/XYaWgDHGOS14BjANA6EK3PRzu4H2VK/jxRQKc9fDl2
G2D2OU1XmyWV7elBlFBxLu3KsXEcd/ZBxzWxI1E3MhVCyH/bqSRzbfqs1JOR
WwDPuHheXevBecUczE5V4h39vO5zaT83ppWoK6caLxM8X5a6H7An3MlaVg7r
/eahzqe+l2/jx5IVtXRZOzNm/WuOzeJE9mDM03QcWUbM3BCvaOPnXu8gNdzQ
/A6lA1QEviFXP0gy7Toz9XzhqPKGiQ9Wk4VxG8IxxKRj3TP/udk5g9ZD0Ucc
262KGSzK5CE/TL2AwWCecfvv3gwSNDXwWvxw1uUBhyjlv5LDn4/rOZ36Uaos
OwN2AEbRt+zh9LB7qn3p/QvqwswUDZdAr3jDPwni5ozTUfo3fOLNedUcNTBy
ugxYdPO4Wk0I4lU4rGQ/vQDiiP9AIbtik1dkeX9B+lMVyCUcexBjLbfR6Hmn
5p/TL00YMV3TAmu3f40dKd6UEV9qsgubz9RfQBvR2YXku+//D7AlE28t8OWb
HPZCEPONMTqWwVoufktM5zodwxgtz3dpksrsyWRj20e8r1yyad/ibk0ksX68
PCLXWZLKWuMbBU6itBKXDMscRgXR0BCTUpQG5HNqvQ1KtG8OYL5zoenl+LSj
RBQ1VntJnyCXCNLxS1mLWFTl3YXgIVSXxZkTJkpbPCp13Tn7NmVWuoWQX/VY
ADLGQT/Zx0z23YHPCDWwyQ3N/U6NBxUROwrrfGgmVX8czNjs6TB2+qYShi3/
hvPJMQugym7PgMcHGbAtKCOSw7fdesyCVCt/gsjqPW+atydjblrKTOtgweF7
EnaVmKlfEJplKZiCyMMDycx7+WPFO/eOxdFaL0fjm7Duzt7f8yLeEz9Jg+rt
FdAEONdv5mcYZWMtSJSlLoouZkLbJIvqI9+Pb/ffeRNy47FFlH2K4a3UqUc8
sCym/vzOhfj7ZTTzL748G4zt12l4yL0Jr4fcIi1nurc0KG7I6AtyAAqvE7+z
OFoSuUmZaRQ8OaayrxFn5aQ97ceAcVUhYD6GdBAhifxEfBNxm0scgNO+mkHA
K1+s1Zf2vFvqN6tIfD4YtFohxHaa11bmEzi2wuVkco6M8trBn+iXJ7TD4egI
0arolj4VouneSu2ZJ/+dWbBDPYBjRuY3pYoX9uHlIvXsvhnSPZWo1Yy6vuPn
VsRMeei+iuD+GU79PLkdcllCORO2iW9iagTb9UJl3Wg5DJBtSqTRA/hCxotx
tWjCTzbJTa/r8TrFq81afyoCUT+wy25w0raPGqdBr7YDCJwtyQfDDOO+gFC9
radnHb9dK8+XCddN9n/aTPdrNA3cGebf3x/0RMu3ebdYOetJsEGCxPlDjAsx
MchD4Nxf+sNP33YwivvGXofqnO2mmqQB58Fz87UghpfvDELJBvvMgisKEIwf
Vcuk9UafDTYRU2/pAxIh9TpggaZQjhBO5UJknASkSZoR9jPL4CE5F9/Txmmq
oLsypjy8LOH/rYugyijaBPlAqo44ZFortEYhqx2zp4pxwFPjLSpSYguFzu3M
cRO6LiLsHIwLpchojdyccyajSArR6nmKh+Oi9XIv9WIzqQF1DrF4JLriH1aQ
EbgzYyBqJveRXiiRP9OVvTLiPvMIk5FvULZOeoCdy+28LACZ5AL+Do5wGuLs
1hFCRC4vZ6CqxT0ors+xNBZlfqLFrOxLtjUFBAdfrE6mmBfb62N477kf6xCs
faD8TwjxnzIFMOR1AhO64PUAns5z7v0HAsTDKYzX9eeMgVa+MaCE7OMPNnWC
eXnQgn54jDZnuRH9ScrKbxLnVjiWS4nymUtHbzgG345V4JgU4nKy8fmbvUKy
PJ4PisSBmA3j9FmTaZZ5qE+ASq41P7yrMQHzEORUZjQPQHKvdig64tseI2q1
qHyNwd2BjPaQMYpixIwl46OsdqEmi2/z9Zzt143Ky7JsW7ZxxlJURqzK0tau
IdjdHb0Z3rE/VFOxVGas/JEjKlIWJZi0hJVqvrfigDqyb8/4jr4cTtUelk67
B1JiFoQAflIsjIhVVmuV/+TlyNjMfCuUJPA5boxo7vfyOMcNMBoNI2rnYQ+Z
aQsFykuQ7Djj53nm6WDUcAWi+EC7ZhK03Ma5ijEzB7r7P+fM8osphnlNikA+
OhMAH/pSBldjNQ57PY6b0ulj5fuvgICnWPDmpOwQH27WB8PWTeguKxh2BwlR
f66gDFZF+y5FmAaDLT2FHhILSXG5pAxSlDYDrDj+gqDWNxp9WQFeqcq/z/pj
K/C3R+7DgySjvyLlt/2zKkiLevPUmlWwIxTy+9QJH4VheRjZ8EALhj5xdkef
lJnE4fNHcivEuYdLHQ/yMjKuRpCJqfTfpm2Tbgjb0F5VINyk1y8plZbX6WiM
dkiXmm0NxFhYwqjulVXdb/1uXTtW1bJVpkDtlDpHieRXLXhyBD0ro4HTOkta
6varUTxteqpi2ELXKNC8gaFJGI6gnl9MxmPy6g8zzWXpey3mcABgHKd+BiTQ
SsGKvlZiIh78kOgL1E0vz259NtZvLJLDYrm0I03TFyqt0T1Uk0oelgXMdWk3
kukDdsubtfy9xSLKygWQqdzuyOuYaPa9M8FwTArOAw7aEvwrH+RjzehyY6i+
7ypYq7+tKsBpWO/Ich0h5yh5/7qgj4b0LLqUpXy9t0dZTG2LPo3ew29TdI7G
Hxw8u9+w3qi/3FBmoyoaFN6YFD8Rjts4we8/lq4qD2f6+1OYJRrrTutdMhtH
nahBSEO3CcSmUKds9Vt0/JGKXT7DhK1Fd9KpYsKh9eFL6btE8lBWI37TLooh
OGq1gPa/X2oH5Qk7iSbpYIrLktWoFXwZx2y06/Qif81FlO8j9jY7kWvL1/QF
Dkjx/qt4TvrY2Ux2QHye8AOP90mo0z1QCevV8BbY/1XP0Yq/TY33yHqTjqOd
7ku4/9yjz74k11A7G1xGtzIvuJD5lecNBNNGtFQ3JHUYAvjlA7rZwiGq3uBf
xejgfiBdKuZDDp83xcaj5QSHjDMhJ+Jb1oArB9fJgCPVKi1NahuywIFxsGeK
sGeqBZlsFQFbLCq/eZPcwXGkBfi7WifPox39sPD1XBqcr9D1FOYwSJ/sS/10
+NGT7D/fZvaacpXFLort+AgAd6bDda1R4bke9hl+j98jJ+C+c9mZj0jz6+fz
a4yfk99JpOG/izZ4Szbh0Dz6etNUBUwUEptnAeaaUfE4CxdoRDuiY344GGKh
4qexWtPUq7Uo9hBXvA2k/wtiW3R0hahEV2hR2rOvD8kzvp1GoOYKiJk7T4He
QEJAh8H4cyiCpO9ZqrDlsolVw4o0U88DzkP/qgeRij7AfpzPOr0LQbpIZ3nA
/b4nbLe/mu1jd4ZSF1dlaLpIHJOEFZhDwvExkM6DnwTnUjIMZSzMueIz5FcB
i1nRLD+/6zKQK5WiGZWAu3PQCilAQ/5LnyH2hs3XBVK80/bMxQWnW5Vt64mZ
GEx10x9fc0L4rjJpfqiu+WxqlTpKBEFcbEX6BSgHmVMsVRXtbKIo0c67lPys
KYWoOLdLhkkZ2IVB27BXBhMOMKHXzjfXjmHSRTjz+QqGFGH6B2APHzFh0NYu
qiUbpk4E6zqx72Ortlys7GSUck5+GrA1zryH7dfCiOIV6N+4M9Iwv85wE83U
WcGOZcIhVyLZKheYOBv2qrxc49pyxZZnFCuMHxBslNrpuuzA90fmI26CF7u8
w0HIRT8tY7BxrI23X2RwSQuR6XMTvA32CZrBk9DdLdE4LXKA0QFbOFs2Bplk
Tqh+V1dpu8Lz1b+gfaJvMTGdSWoXuHUom+8L3YOjELufN7zL71c7Xtkx3rSs
omxDIxV/vz9kccaxnybByseYsHE7RQ6uVQsjiCmlJ154RFIN+EEHLlWsWiQX
6gIxyJilEQxcKSwI9Jve0xK/lczKbwmx12KqlbUDLthGTlUyUSbWpG7Yx0CZ
qDHerXFmejeCnASi6H8MsFmJTbuIpOPAGmGkSZqIB50LAYea/iNF9VcvQEdd
Bi/6QxqGa8uXdhJXkHxYNn8HNljfdyMIMnUqMgPKbRj2Fw0aPA/qQrFdHmoA
MEzN5o+/sGHMAE2jeXPfic9l4S3xwRO4xgc+NIdr9nQaMzB9ljGnYED7x9yj
FFj6Pu2rlRp8gAI/4l5jdbFcXxm/UhkOL2BfVXXRreQmRnkhvccaFbrYGVCO
WyNXdssJF4JOjeuQxVn1ofQp/Gt0PP3/1nOaLIkHW0YlJOqqrrn8b5L3akUE
Bjw1cUOvRrv40YTq4Lk3j+3QLW/5QopiHwVLoQLJcaZip4N8cxQVOocNqNls
KoQXtdX2dAzlRyAStsT+HOVx7eMYIOZiNNbieHemrd0cpQhizhN3f7dK1fyq
x8fsr5su9AA5hXgfaasUifr2yvIxM3Ht/WGRA8PkfYnPyjuZF38BjvvForY7
ZsBkTElL+EZWUelACXIB1L/49TUYt5eaWJIyXZ2Ud4GL09+S92sxJQ98d0MA
2DnWVhsM+urHyRyc98uaU2aOJes0jc/UV759dSpWSJBEglCbsBNs+R4xPQuz
LS78s/rHvWKJKt8JyXWjyzAQ6kaSoTwYIIjkjDcQ/MvuUZBtuKGP0oMpysmK
l8e3LOsx3QpwT0SLQosAgt16rhi7qVh+XpDj9ycEI6qswflP+pKQlIAY8aEK
vqXSdilKYv0EXxBxNjNomeFvQUp/PsW7C+afoLuzvx8TLrfgyZKmKqyAYvZN
hNQNbamaSPHJYV/2cTJQdIzukdrV4aoNrEbletqlsYTYfmJMuL8rn9+obwSn
xV6pjQDijYzVB1JFucfOWC/cAKsov8F7ASWzdh5Jt+8dAhDod+NRsfkE8tAq
L7m4aREi/XV4oroich/Yl+e+DNbKVzN07wSrEnTUmKpos4G8NrkV6ChszBPe
5/finFub5+HzMRwWZWuLsOlFfaUhxyaJYA9t2MG5zH8RECuuPx1nJ7I65qa+
TLqck8WIHIAkPKh1Bc4o6eeZfUSgPg+KIov+a3w6CXYe4ucHh+5fubCO/1Sy
YVSEkpU9oyqt+eyc63w7RQdYpYV8pkuat2uYO6tljaJQ79Agozs5L9qjUTBZ
51tfdXQsM5GX5ZygtULufgjz5w/YyytPiNIPX0dc5ClzPmZc4g9wiveLDe+3
tcWl27vguQuzmn71Eqeh1M9PZi+KnB9/Necls7T6TuagJ3bFXgdqJd1+axPW
l/1Vkl+vLBYkHgBW7tTe1rbOUhPu/lM7GAqvonA7yGPAwW7rJrT8zp7g5x3f
7N7780Gxu8VyHWcVi8Z2nkZ5RBhwbt+fECaXuJ2/pNka/Hsx1NumJGShesyX
d1Ta08KMDiALJxaYxHoyuxZ5JMdX9+v5LKDE8HMiscf6xWwnFcABKdI93yfr
syclmvYnCb3szPZE45dldBsjrovIjgo0zD4+qzyNlPQSBP89+TDvp38PQ9s4
nhExugmyzthenGCoT38LZ+Ip5oGNKJbeLoq+iuHlxgiz3SJ5i3iF4fwqL7zD
aY4zv+L/cEMqepCJ25NGi2pyMIa8wHzg6zlWqCXISu3LnC+iOibsP8b9nsfL
19+iUu+eVv2Ey+XAcqjokySl3rOyjskSGN9Wu7bSG3U5ZqYGrPCJRdpeqEwu
V/x4YorM7LTw7coh4mZuC5ZT+tZ4a3hTK32oHZjDly//QsZbwnDsJoGKFTmC
f81W+uuvbjAa1T9oExzVK+jGsL0/tRg7QBVW+EuZ7LbdcgwGRf/dMdgEaNk0
lgRGNPhLx+B7r1DHJ6HfNwGyAYxadOm9MCzkw7aGMM5DDuISl8cEVfAc7iBq
zK7dmxqz37zorfo3SvFcC+F1UtWR1On3bGHavYdgL0WTYHDLv/5aXIHrAMan
YjP4oQvxRfQgCgM+lvUhfrtGQVRN169ZP0OQ+lgx2WJ9PzfLlXAjKumFIDVH
6V/6YvFUTIMNNCa4MUEJGIRZEsX+eiJbQl0TtaTlksZgrvrNfMrciydrtQHK
63sjOEkrue+toiIgTxJhoKA4vSFJDsLJSZPHbmiMz3WajoTaIV7u01Ixg1UP
EYtv7yO2/F+MAy0V762pzudZv+I1JSBfqiOXVct3hL2/oOR8bq/+z2AOZlyg
YU0taCPMf9nKwkzc3+meccZUvdgh4O/P7nKkgi8VaxHaoZKPXNctLotJmnC9
K2zaOudKlFJWZlGe6GxAnqTB0QeGF565ZeaX6eodtU4DW/BPq+pd7NBBQmdt
5qFGdcVoP0d7wH8oO9FJkghvzOgu+SHlPrMdC8f9oL6q2ETbg6XNqS+kTXNZ
BXoJVCJNvMhz4gBoz3lLT1lF9/pxCf3UmL5BqlW404Nsl4invJGFB6C1i/o3
0vOp43fBfHliUQO+qXbKDhT8R6CTX2ME6CyqsTVEjNxCxwRelGHUrMtU0U9j
tJC3pXDEJ/my8KgjpufTfJG9UnQnxSdXk72RDxV03kz1jgiqT3jptxWRp/aE
/d4vAuIXH/5EFtPSqc61ugzsA5l3WQDSwS8ttvLSkj4vTqAx62NQljORqv/F
OqU/t5RJRaTu0YVL+9DMxLqakvx6ygXDF5xbF/TLxDq/Xy7Bfzb3WHVj29P0
fJdpHCOWh8YQUsE8y80jY1JTEAJlISEkYtee/Ni007urQ9d7aTHMjMDezCDu
v74x5cTjdkWL6sGgbv9juNuILUwoTI6NLu6gNb7St1vhVA8FuwXFYOs2jiex
qdmw5ET9AZhQZG7fwtYMvu0vIvJz0t0YySc7C8tBYTrq62B+cAu5eXXzFql7
gvPTuVEwAk/31bZTb07/9MaNUZipvxvjdtr53mlCEf2NNCXQQ1AZIj3QAJkJ
tycGoqfdR/4RylX4mJj1S5Qn5xqJFa4gTb2xU0CQmGkT2Xj8n59ETkXDgDzh
cP6KViHFptWV75KyuKDVBjPo19q36WIUMJHOXSAwIpH3guTcjPbA3yHaCqRC
ek5GpmeIQznyLVCocTBuR7wgWzFZe1RKZGyxz5lIoRbg/F8FJBy/9lkmXub0
wJH6ozd/WZR/2xjK990umAlzF+6GbgJkDVyfCQF3PcCan/me3vCdoyRxD874
K9ei3L84S1VTreW3M/CyxxVV/VQ6SqHtn/q7XGC0DBYNgw1/1rax+Vj8NdFs
i3ZvNOlH9lekj5xZ5bRJWQlB6DiToWr0JgEkEf6w/I/znnR/2fkRVw83NkAU
Jnc2/MjDuCussHDMBka6LefW6aa8nbS4WVTtgJU5vLDDq7/61u70KARZV+da
Q9SO+nxxwGogo2y2ZSGi9ghSV5IjmwsVjZwIt/BugyL2TviYf1wzkj2ZhN5L
bXOeCGskz+dQHIi50JFgqnon6Vayor2+dO5pGlOnK/HYUzobCGEuIywd9HEJ
DQtsYKTYIWTs1y+zjeCHrpplMz020WjTwqZGmq8l6CLd47Zuqk/bjp0+IzYr
ttAPLBStkN2CwVS/s4UKWl1zXWOfYpOEkRUzWPYGxwu6Jv93uBKtF8x1HWWV
bc1OBGkUT3FwGP4nzZv72v+Kh0NReiR8Ed3bu/gKuj+i4VW5shvqokv4WEw5
xInusOiKiDQsizNuMhUqSa70jsWdWZRqRMeDYnVnKb3J4MavFAj+Gn5ENZHf
gaJXRtduqY89xOaPBv17lZEwYrZusyZ94O5oYjhSXPz1xQZzagSvmzEflmc/
6kjmnHaMz6vkWfT5TIkno/Ioq0jAXbAolSIo8PxMrHgeJ4DDQdweSpuNxTjQ
2oPIOixLCrY6UuRuYQzOAE7VtQGSrxo4ofzOh7dwvXeXVb6b4gJdfoQrlXRk
V8gcMw/KuJp2BnUwiApeUZF9TB+KS9i6UMpg7Gd618AvWU8XoxThhKWcVwSs
99s/pz1+ls2v0zFMQWXo8a4sLPAL2plv3j+nnnCqN9SHLjaExgCNX8CCYLI6
d74RwGJ2uQzZcRf0JtaT3kihTopKIy25qfQaHzj+NM/xldhbGJDc4k7kQC+k
OJEJn4GY9SZ9qWkKyb6KIIjeVaWEBCdM0sAAH2m35Krw1CwMq9AOPJ6eqTqr
53y5fC+WJRzdSQbbdwk8dKlgTV/4/1IYWd9KH4fKPPNVOUgqgdirSaP7W15r
5eUpTeZPt3KXE9LsJstFZEVgQ2nXE6Gli1iu3IQTczIK3bJLaifnnAx+efGG
X95hpmGfRXlgyljDAlbGDOppMFeqqTt+bblQzKngaHXGTuiPMXUmLCH8c+Sj
LA+XHh1/376HwIfuWZ4YPSoXYDL4GmnKU3zHwDSnKwFMUtdAslAfRSkZLLOP
alzRMI8Kc3c9bEAaCwHtAPJOJ1tQyCQutEv81JUEo/VvyKsMPN3b98TH8LIT
H1UxiS3Yx6Ive11fT6W1W7l0ZFa4pvsXYe/OvV0owPZ1bnNVYmBO4aHO0VV0
qO8p9KQZCvYaO844v4pDL838uw7JpQtNItG07VG1HESQvOWEHX0BKnJWwdsU
U1Yx5ck9VhNd7bgTKLwDxNtjn9wmnN6Bacrk4iYrp2Sr2yNE14GctCTdoygp
u8eYMdE3QQ6B3VbvoSioszEzOIUcC5u47vBj1yTzyfwDqA30+tZQYDku6gKy
bghZJyO37jqCNQGfh8aNLlk0xKdylfiV37iUPVqCZeyg2zvfpGqW2oBAkDXO
CzQpPzrdhmvpYxp8pPfonZZMPKwmjVft+lUAKlmulH03w7oWHSypo9XdRRYk
WCFkn/EO3q+L2ZTtJLhGmeDPApoddkUpXjluUanIUoeemtGdSoFVYV2F0Mob
lRtuXybF6Qs5JVhiUp3/1M+YZW/AG+6ew1t5v+M4jZtk5f6jqaETkqrJOfJO
T2ylL18fOQDVDlh4srjjnVu00YKAx8FxvlbKbVChSNhct0OHTfqh7AukCjwm
7g0J8RCu7P05b+na1LrqCVODAnBLFhhm5shIHtK+ESkX9BNUmTAg2gzAwd/r
aIzWOx4nAtd7tozHuMrtbtNKtSy0p9ohPFwoCxBe/lkSmsmp4cTDHBeCt/qz
pwGn9zGZqp76kX+vWuAnTWAqWkozCDa2xcbS6Z7/8CXk6g35c9jNkXixMC1P
DCTnFhGPGyNfRfUD0zIfnwA2HZbfTyv7IXX+aOslIl5r6Tya3qSr5cMsnyn2
tXXqRTTQzpbJRR2i9odVr8K/z166SB7VrVHhRsvNxKgj66TCu4SSjWfTibz2
+qlypB9fewWI3cf5VhHHlu6IsFtaZohiH4LROCMrEF70qwTGRe18xiNYXJOd
k2Dvu6iEeoENOxjLNPXw3CFdbUTcHltOzX0bWaWLPZglmqnNhu8myV7p0yy5
S4ZBu+zXCHmjw//KdTCLesx1RBUY6+UgBdMiApqP/mbBNgq5a/QYDeuOYMr3
2LofqOiUPk8bDfd0La9vVJn4xGxWUeOToyAfck4N82eBdciclQM//UtaBVEn
EC8QC/1zml2rCxRsfNxVuhAwZ26dSl+VepHmheXpm0snHcA9AodSHtk3UEJJ
YO/zcMcrlpYQOYewzKOay1J3VWBr3PpKyVughghFPgKeuXm5BoNjmP0wcY/g
vX90z33DMJE4hPT7jx3OyNW07tHF/FRPpUagfgK+tM2kxoGcc3KfWEc/Wrjp
PZ5wKXpEzCH4ZlQnBMzVkMHAJgfbUw/381Dt/daDRcLBmeBpo1QkhjSHQ+Yx
mLNinLpREoZZ1vIdnPJv/c/Uck7E7cWWaKiqQLIwf59MAXAFGSkOOsaf2a6P
4OniMgYMjDiF85d2+Sbf26EuPHnOUwhLpMlW30x4g3iXEYL6GXi3T42nCdQH
6de6F26Yn8BC+e/Qjeindd5ZzARiLvDPuFvgXwmYbGhSS0cmjCJdAlQ2KHJL
Ry9VYCNhNxDDgSzXSNQYxjJwdiykKCmEMcz6BokM5D+VyeAYwlLMQFQ1nfVu
dHvRSy0ADUZglmqpCfIdtdzoXasGXeMbwq838dlMvD4nq21nLu49Ocq/Ex/O
m0FloULAKod/s+axWv0RjL5KiCl9sv2PQKvygTdjHhHD52+hgohr88q2QY2p
/e5eN8nFZBytnwF6QzvawdIOqVa8TzuK9a79gzWKOUMF6sVHSufw8gPXMWHN
Hpy12SpMOiw1Jx0jeGhW8KyOhaQUqyIRwpS/stScQNvBxZsd9xUnUHT6nW6+
mNEk2l9jxzCwM1BYttK6C2UA7Fb7GlBES6zjY65fpVenBgQk6031NbFEvJdH
cOuR2q2vFfftmrgMej/FB+EGxsgM+dY2MMT6QL547Qlb1KW9O7l12M9G8QjN
yfI3ZoYsTT3Zr2ZreCP8fQNtZZSI6swRtgnSpW0AKwQxyKc4CgmdcyKNlUom
2q1Kymk7dm7CC61FZGTTDWwFht/hBjOZ5s9ZHO6WbxGK/CNzK7SwoVs9ha/o
yDMYLtAYHqzqPN/T4qvT9PoPwkGb+xDvSvQRSt+9UzL6G4c4sjTEAYLXZK0V
i71VFQN7cdLrc1X94IBJjvZ7q1M8COm+9QDkYdoTMIJ5GyrCUoXHLRRojXrd
MgOMqRS4i/Ke4HYj9S1yKG781Wo+7y+y8CEnpaLKGNqjfupvg8UklIg4DFmH
I7lnxn3xz22WBif44cHPRBPdq0hfp+rzSKxZrwvYq2xJIF64/ZluJp6qmGXC
FMKhSuWLHXJtLRNGUzf7j1VwQFECvYPDl8ynDH7njmjuDwItd+JR6FpDDrup
DdxJepnzO1sLMP3Ih0qwrJV8MCk46QSE0oqxQbNLJDsu1zFzhef8/MJSpjtw
En0vfd4DSDHPmgHxweEXHMMHIn22UTetI5buOzEZSfRY7z9J8C8VwAQvk8d1
5kxonINCcEOfegMTcxOn/4HeTVQrNPCJrRuBJsL46y6aq1jCbKaUx523vL4I
lePjc8RT2YFirMv2zt+HnwZlRdG89T+Kl6VLnn0jN/xQA1X/KU9+MVH+trL/
YrNDytJtF0EcAL4sUXjTD8256QHE4tlehgDTUzA+hpewHmd8DTvNKMzbDcUg
buLWiybYXiQiVN4YVgJofbtJsAXKKh9iRWlEwMiuyzSWBT+UMcqSe5C2CDjC
C2e5JR5IczaZi3oA5d6RPzwf/WG8UY0rtmwRZg4tELyzo1ZcviRKasdYXem0
kykZE44lHtCULYEGnLaUWUYo0WjqVH4beC9Ywqj+HMqTcapWVmntNgRO1HKg
YvsfTEAkmSmQvYaX5ixu9J0mPrqSwe8vRV23sbdvQPayAhw/lQgpo0UdGN3+
gDqAaYuUxkEPXg/W+4jfJBRlR2qwWxHyOiUKjyI9CtZnxevJRxzyRHUKWhmV
DDKabr6QqFH6CeOHrhDTNP/aduF+k6Q2t3L+pRlq9+g5fqSkDOCLAsb070ba
mk1XLfoG6BV9g2cu1txf9Q/optzP6sEDXoT/PapIlOlfZAU+vfVcMR39ikwl
0/lfGe1SVMAmyXfR6PXqxfpcCBHiZXclKz/rR6w5auRDAxuB0wkYRlgPo12o
y0iFXjpj0b419qBkgMkSnV6aaOZw4IanewoYSUw5fvl3zb15KyyhTvAQTVgn
Cc0sCH3nL5DLhplgifBgcCJMQ3GBrba2XYV2ghc4TtGAKSwEevMBF89kgxEo
/47KjCGDJYdcCP2nbr6e9rJzpo7o1h202U2WF9GhSLVuduTJGdya7I11EUWW
y/lNlugXcC70ADgKYfJ7dIvLFNQCXCs4+LmnbHgj2xdVWadEBKA7ia2QH+Bu
ln/zoHR7wm09b6A+gabBLcxhWtxCjE+XWYKvu3x9ZE28WUxSht9XqZaJqhWL
2VlxUSvoVBMBpx3XoTyOvPjTMI09LDrQnbTdSZhTa9XAT+ODErHzNY+BGLmD
yYk/49k2cEOhuUgjYAPigE/3340ljdSLFWCEQ/ifQoa20Y0IFUVXueGV9PEG
DwksOVMeJgJPIlkPCUBC5ZAH+ZOTKtIAx/eDJmtuVk262aCQGJqcz2Qbswrx
UxaLlQAyG9TQuqdCpxh1Q9JT9COlw9p3kCJFQrPHJTgesulUx1vR5zJk49DO
0UczNebZVxg66j2HBAuZaz1oYWs179gD01dvS+6O0ursBkEYQIJJzJSEw8ln
FpX9PJ1afhONM9xd+n8FwM4H7pOTKY+v1fnOXroPe3DVZ7WXhoLgPQ7ahNHw
1TnBjSwU5ktBtNu1y0jdr+yyHLMGIFBjjlEZFW4i3NE/g+w5GGGp9m5pp9Ca
HGesmr1/9/2pYJHZ5k7yS2NdbZ+SM3BWCcSPjBI4M1E1cIKVtRUaGHRrrVWo
de2uTHaetljeX1UWA7NVIg6aLP9fSbilYC32s11Rr4kXFnxBj4BZGkgfjdoe
3cwsKSAozS11d/4KRb4UvRUEeTEQ0jyi8vJfNTG4vbvbakuorPORuODRbC49
+SUBkxH7lUQOAih76LM+fyQmywXUaeiO8ZLb7zPUbgIuoR9iNZLb3iFxVoM/
oSTKRDh40shOXgTOClp3POqBg/zTBiY62u749QAzw/0CttbTgpZKH1qPFIBz
LaJLlmkM+8csR4xxDyoS5rm7kXmz0GHkV01DqQ2FtqvYE/WFSWrVYlh+Z4eY
pS2y+SV380Pkk44i4oVBmdWUUMS6ljxzJzrMtl4by4CHuG8WTAIk8j0lXKw0
Q5PQHB92HiouE6Kw4d6+RwsSh0X0eIqdHkVnvEMa0SnscF+A1ujQBBJFNHaH
uJGwCb4gH73V/zM8HJoWtvOfjzWGIRLVpMl4/aHplaZUbCc06t9+NyPevZOd
jvI66iUhOl+cIQK3dtnsEjl6Tp8fFlC5G2LXtCj52QOEQrQHKzztTewfj4rr
326i3nZ7e5104vp7lbjlEogGJ169pzmxJx+DeMApgnDx2fnRgtXr0wCXDdnB
Z/o2h79tt6JsU6yXmqK3xT3xrw5bZONOdd+nPaREI6yl0aAt0q0i25eahrTX
GiHztGvsD9BOd2n+x7Fdw2Bw0k6JfU9DAjISh6jvl2GUm/YUIX701HQkHcGZ
8eblSzFK/9wr0APLfishEjPNKUUkT4NLxMbXd0hhyhxYp4MFHKQGCrRTruNf
i3Xt/j3Hs+4OXPQOyPIfk4gUgFhD9S/V5TVbdXJ0mae5HrkaDTUWknG8dcLw
5VppVDV74ImEbmJP4+UgBOHJq0cP/B+MZQ9W7t+ICjcv0yJBr/kzPFwcm3Og
26ADrUV2CVUhqJdgocFlAlRhDRzKStMhPYuq2xggvk2SeZImzbn2OsAE5Nx6
tAgATXv7kThetT6FXI8JRGQCmKe9tmqTm3JcoqbYrcG5JOn/yG5uqypi/VVT
UKw6yOKHV1rNm2kWqTRG3sKKvMxPUBIthdgGB8TIJqDc3IceGNStvF8Cqxm3
ROa66LwaExkirhafI9MI0ZpCYYo2WIwG/bSUaFTa92NnTHI1NIGqycGsnmeS
tpmGsi0wSMLOyDPKY/qiuXeDjZv8Nd9HAH62dvNLM5Gimp6kUokpcAVkrhfu
kVLZpQ5r7fNXryOnVwcY1J14vefZmwLzS0F0szS8/EuIrUw0y57bNzd8q5RM
dibXTEJhAmYhOR0TPFWHsVCSSOZS+JKr0DZQlUQW75++HKCmB5MVH0ceGil/
KL5iZ3B/sloWbSZd/5eC0L0nzMnP4DS0dcwI49q4EX98E0K2sDgAb0tkH772
LGqsaTGbuDSe40OnjqRalOD4qH6mSn1mcwVvMHS3M6vD4rzxGBhQOjMA5Qfp
BM7TZJWJWE+e0YKbpIPJdyu4rLK7sAMyLW7o7cVrdDtyIoz7L80/lPX3EVv8
xTWcba6sbwhw1gsG+PEARnAzHwXgFXr6T1OAwZ4sf4QCEBRwRhbtfoPyaUfA
Ejd1INEAwieUMDdfp0Y2uk2T9cEGrF6aNJYFFu/tirTYJeaNfdxsExRKNdAi
JlThrMDjIBsw/NX1Q4kRZISczKAFis2CokpTTyVPKE+IVNpucQqN/GEAALY2
b6yas5N+npfFZ9SNhReTkjvfKqLLBDJJDQ5INdmY4+0XQvy7ie7w3PRlTcLm
GwC0RrwpRuMoF29ZezTZnkTAqDu1OJi3wUxKi4zCZu6PRngjoks9ULzhPdSa
rY3H4uoXPss9rwxo0+kxzYWwdPQykgpr1Ww81y217pG1+Y5K/UcEuQDsB7oL
Egj702Q317x+Q2i3W0YBaXT55qNFfUNR5cjtqa+UDP/zWiY7IwBD5wOH5xJ/
j5WIJClwa/ewqFZkHriY2O5nMnprfUCqTz+9pQMc5aSKfOK5k9VExR/cQsRb
ZMd2+cIa1yPbgJsvv+lbITr0P8XfP6ukSy8kFfFJE/sMHDgi5HUFt1pojnRU
/G+YVSp4Wnv588sEKRbFfZi+ec+4mAEcQU/78wqDGmgCgRFC2psiPmlgIU8C
gkoIeKT+OVM5q3ZgqYAJlzK+0q4izsk1HSjbixlzJBC9pjvH6ynyRjUA33X3
bydwsT9EWfqaceEpe2zEWY7WfpX600PbNYlqite3zo1Gk0Nos8dL/l7ehz6S
wiqtCXeltW0wMnWSYn8l3QWY5LcJCgG3d5+g1MCtq+KLN8vJO8H8w/JL4mzr
jSORT3UyipgQY/HkDujfh/1heiMcrMW3qT8bGV3PHOAnV5SfXyta7EY/2SaE
J8SeJcKAXCd2z8Jm5v+kJkihJJ299rj8HkshKBBwaRhv2Dtt+x6GIWNlrRm3
khUFBGx7Cnqe32fi3/TlA7+zMu3EfX34SLxjY63y+ryx34U7bpz9llgVFNls
7spuDl/gIUhAsHemKeUlzK/8p6eLgbAMJkYKZ6jDjLAePYBq8Nh3xkmJiJ9U
x+9Xie/+1KurWVsENeLghKX8bl7a9ndMRHcQziD7iCJMmDN5EvURqjqUBolA
LCMvssn4LNcxBatCN8zsA4AXXnM4Q3/w4oS92h7u5Xo6Y6+UsKHukWBQVOFJ
L4mc0Lx6YLFaYD7Pz4JEm/isbXxWtoWKvlidSC3QujYAclCy8nV99YgPDnzB
uF2y0DTr0fLg9W36uPX3RqPnxeXMuSlD5M+6FsMV1Fct/JTXgaInyMdjpox4
8zHU0l4oj9PwmYta4/7bgSlWXHjyao94ke3COxux75ZWIdz+UiEzLmC6tMv1
IDDDuhfTspEUWP/Wab7EwduoEndyAKkABcyA/SiQ9w6CvBkB/zi590bQwQO/
MQfL4Olc18ivL3pEzBesPsv13M2Z5de5kSBUCg/YcMS5kXjycN1fbAi4TNvn
xY1HQTb9bhYeCG5/KSJbOaYnCYLVicaLIVug1Mfk2Fqhz5vKrWLeWGpCm0Zz
WRSLCt5GeGvQQgl1Pr/GqZpbL8KfE7tBdWKmh6tmm4/9r8Rt6B+0MD73DJBe
MQ4r2fHrM/f+KZu64yQkQzr9/yDqEz8TRGS+OuKuhF7atnoSJFgTGlkyhitk
PI5g3t4wsXZQLITYEsHJqzDqtRy2e+nvR/97xkqM95GIkPk4d/W2N4rym2Am
hSSMAcyxhnQ3H8fl4dxFbQ04SmGM2ua/jPGP/HOoRQorDh1/QFqKu8m7HQt+
SiEwpk5QRLQx5js8orMfW7M6YqwbS2D2bxhHFsY6LTUPv/JD0see92cDdsx1
aA2bYoMWuX+T951ILF1Rxs+ATtEJuL8LVjmUGYS20frLLPIi0FiFQZDV+sL5
hzzhgIZZsrEGlJActzZe8MkkyZlPiffpT8GowruCkBWXXrhHnJMRYs1PsfS/
LUQD0kkoqGCd2IrhrLnbYgZbBzBb1CmQrNRYiPzSqrlgkWHIodQk65FDsemQ
db6gXx3nlTH098ggHFlK+QlTrUvJ0PAMcWvUmsF7No30oP76x1j5CA7ADx14
3PaPzxWOYba1o6QZ5S4u8Y+53vXHHLYV7K0oSnO2AyvGabXkDcXlJJfwQKvr
WQBLgrnfv3kzjjHu9V1fUpNBiJyS/cu6UsPY/BSR9zalMCq+WKqKybtYEw+n
Fmq59acXT05SO/2Lf6F+WkLZj4IoFJpddPJzpwiEcp2UbM4T3cXBjI2/wLxW
m+CTtvPP8HRvVmJGe/1nJ4FGaWWMmsJaMaPOKMGhfCb3uYgoQPnhAotlb9eQ
aFCtK+2gYOUVmZT+KYXIbUL2WKqXbxZNm7uKncjDYCmus4kI2w4VukPjtevC
QofC2DCD3kKTYgD2ivQJrQc7ukRGcExkFPxtPvAQ7elzR+3B7D5GFaoBQJZB
GtBBQB2ROEVS/HI9pUx9N07KSct6DdSmOQaL2am3wq/ozlcSUmS9qdvnioSo
zf5NvTiCj0BA91gA/QDKlq428cfSM599G9L9b8lUhsuuzGNoxgeXQQbXtwnl
XDPnE0Yj8VQoBSTYCS9lfbs6AvODiFX//a+e1O6eMRe7/g/H2MwGzNrmChK8
1ft4RVD4J3+wjLDcDbZaxb1DRMv4okdmyj0T9JKVFslHOlOxuqjUZaGB19CO
na3rb/TpGvDezXI5NLi1W1RFTpkOvrURP3++bwlv7/5gARFuUEQuUzSbDeDM
i+kkvFT2itLyvKWSZbFSzZTGdDsBLyo/ZgRs26mBYI4nG9uAtKofPFLjSOKq
kwarNYe2OipLrxy0l7spMdjfp6wXCZ2YdtoUT5z+2fKsM+oNr5oz5UwhdCxA
MrZRDlzQLzUSSQEXnyGwK9t8eU7I5F2OByUQ/s3VNj9JYXx+AZnxbnQErg6X
0G5x/71DzfRpyy4tO1z/zdd6eXSXR6CzIl6cLIGGYb7ovyJsneTDlWL0YYrO
xCwF/k4ui7uI7dyoq/k0AVI2bNM20h+cl5nQiIjV0WguL+TK1E7NaDbNVH9H
N7ZCjXq9dKtTLnfV7q694cEMdjaD/9ZLT7EAdtjiPQvyIOkTtg8a5wc/ACtD
IzGS7FeQBi57pVYSgaWeYO2go18UU9wIyky31C/b0jf3awMt9zdlLFe6N2g9
rfKVAE54f6rL78G8YB8RmD/cJJcTcNwPbTJbJykOkaNFhhvV7ApVsF9MBJtY
c965sAYnbmLal3TuCgUxh36o61Zz9DxWfxwqXb19h3QGZqo0Y5Dj8mYpV5a8
TsihN9Zz1b10blqO9RtyWKcsjvP2sKg1F9crldgouFNoHPMrToAyFADFWz93
1T1FWlrzDOekZ0Q3rjW0dITSBBcrAhXqtRlC5DLJFlVsDfKOs8KU++11KQ8U
lx3yiD2kPP5xOymCN5SZWveod4xDtbix8K2h8YDcoe1ShndPdcIiYc676gHp
WHkT/2ZVw8LMNRt4Dokz+9FBrjPdH3IsZh3KMw+fsG847QWVHlr6PxFwGuI2
WBv6FkPoIXEpQ39GjbE/Myah/lmbUU4PCEPbwSinjDYzJXCZPluQg53xPaWb
SKfZU3SbDoxIaDhjFTzxYF3q5VuXBz4nBrQ7nGZRrGqvhrESnMZVi464WGaF
LFaHhAbBR8pCPSKxQvwGQcO9bf5AjnuuuvYmZh47EtfIVvMWeo2eYRp61kAF
FaDx4m84p0xWGmjzezBfw9KXCzLz4W9lntzHjrIfBSqzMnZbcJfa0hDU+0j+
zmdXeObmJnFyqWd/3GBdaFDHavb61wJMrsPLk9JsjAm+LM375XXnJW5OxIIp
/8/HwtBq/KXlIMl7McyXXFNewaJitGl0lKI7GNINZWDdLXyMSKsnRy1NIrLa
pOCGw53QXKBNfhL5cPYyfPGR5VXx1ayAF0IX3oSl3tFa8dXJXnj23c53JHdo
8zNhdhU8LTsNfuxuhmpaWobAQiVWj2BGmeRh3uMIvleXvTU3B+adEhypyFiP
Z7dDGqj7CkXWWE8+IVTp8+a8cbQjNUqMpzvBsHy60ug8GOqNwJ03xo5PKdY9
fbkOuz/0qHQwfxIezgzlBVUkqGp0UnR/C1Tb3o+YS+FVOCDrxcE0pKCs+fLM
A2Nk0yL5agKsGGNZ80D+KDmxK9jmpJWSonmfZFpNQ2IoMvkWV8Ab178SH6ge
Ap8DIN8IsVloDxndZKsuJyafiuQipakKhWGVPxbubGkWUAgFuT0so1AseoMy
8xEMU5tqhwt5wTI21nHAm8JYzcExY1L8HQFEULscJDL8O4sJNAOM3z+3zZ+N
Vj8VVf1uLmf3hMXpa2YzQN+ApcWFtT24zYOr2ezTliP8b/P+qESipcu+KCnt
iQlhZOSSVYR6+Wr/TptSIyYcEK36qak++phpsl57vgl2L9VkHZfnjWn0+EMh
7FXCzPqq0pzTxLXvMlaYPEb4HWi0UGEQsAWXQ2K62bg9djS3gsDLrWXNPuih
yfY/HFXnpylGuGnAz5rfn4MRBsdadp0e4inw7PrpxgKHZTqwzBFNnIN7KVz6
E9FGVxZxRrjYifcxto9kj46zgEhMex2iBW0NCNQcunVpQG85ZOiTply2MWwP
DNaUkQ8PjBK0WhzGYXsmQESlRO1OmNKjFNRiKPtU6RaOPI5cSB1PqsYbKyKw
e/N6QPjrE9lXLUkPBcMSZXV25HVsyL+vfJiTqcRqW80W0fCiPp6tGJE3z76Q
bwXWvfNkUcLOhKHGuD85KJN1waV7Ixh99uEyYxh0zQz1ICLU2Oc+vjfl6afI
fHcKYuVRsIDBpKoMAtNVRB7fLMe02638TVegyQVwL/53e4+tw+bGT2Hr+iAu
LnAaf8X7kGzw00GMdIgidrlggIWGZsccdmIWbKEyemnM+zQoEpMWLyuspA2O
RFfO3Bpje00Ps9LsP775e4bC91xDxzY4lgjcX5xkAaN14Vp+IUku7D13PXIS
CKWuyPTtmVwozakHTm1r1NeljcL+2KQJ1wvlVHk0tGQxTDEpWPfo9J7BjcSd
UF+hheDJ5wJslnJS/pGjSNBrcppcJGTngc9sDS9a9nmLAAqCsy2AuAoJm4Nr
MCim9PAHpS6tKuGWhazEUpsne5hfSn59KTVYHm5tGZWgQ04TK1EcIStt+tqT
2/Eq6Bgs+o+tmYem8e6Fg262T2o70fEa+6QevacFrMFRr2ZdeeJQ2xTsURbh
ctS6p5/yQhoIerHLFHPSVCaTAqGIv2iB+Fl96x7A43cAhOY9JgKbKrSTeP+j
i2mGxjCp4SxYzJU0leDJJHHEXRKsl1lINtq+n5ffILwt0NNGqEEV7TBtmNl3
ulZKdh9aAitnAiSuCQN6sxPpzvEKEGaD8XDT54anrazf+k1mKZOVVXx0B2cf
DmTeMdf8pVoQRr/TjP8tWlwJL9o5Mq/+oFpwMfJlI3UqLN4iKV0Baqh7ukA0
C9Dp/Dj0jUo1ctxBWJVAW+VtLrDeoNGMwLvwmb8v0GBWD5DyCt3EdKZqPb1N
TrerF7OrKbn2q+NSs0bwqKmqFaKhgUGWwD6X5GJYAWkAemmDrihOpNLm4n/X
47XSQ+ACKFzxjL9vGfpQJ4qx7KUpmh8d5U6RGigENfYCMhgYObGs5T7LBek0
CDkgNlEq+B6d8+Hc5xAC6/o/ZU6L8Y2qFk3BNwcTxauc3NhQzFc8N1ClaOBP
rh0FvzHEuglrrkhQzQv/pNqauI4mcaglqKc6M9iFOgnEbs5tBww3krRY5wIN
7HC3Or28H2f5JrLKQhPfTGqcLEakNsuQTrwKN++zD50jKmL7XLRoDtvAlpkH
I7UennIfZ/onUyHrLGYeg7BjrJ1/Ag1vdQ6HEYMuEI94vGTCxdZd5Wzx0rPp
VyhUm0Ig8KXIPBnonhOr35bQF40W2mEJhzKbbqlYSw1Z4r49/oBt4AnKR8kJ
m8o0COq87Pk9fpZruJHFT1PoV1RJDGRZWBQzLqIM4ceyN+UYgqcURxl1XBLy
1LU2C+1iN5Wmr/7xsUhT/BlaLIUTES0qUKhMJ+TStYBaBO5a+9UzzHcywhtI
8jo/36CFf+AwVj3OTEkVhKNK0RFAc4LsOpaWwq0s3KeRsOWZiIIwcaGb7SnH
fmvzrGKkOfQG6H186ENYV4gKrJZg0fPO0zlqLc1Vv/Phmrb4shGpQAX6Dqc7
fbHr2QZeDVtXpBJ/wmAnhKXN0oCVM6SOwmnQ1+aFpsS+DXqVDgN2yrDB2z1A
7L/DYF9G8q1ybo3jNTAcFaUBpHk7kzW8wxs6fT/mw6GhIwIXpGofTwrnBNK0
mdCqQw47G9kAJzZ8fNaHxW8FA1pNT14XlJ6qLexBEjrZDrZW2cc77H6oYvfg
VHVvNbutyB55S+IBB8JDPr78LAt838tniwxO+Ohlw6PkifrfjeNqXPl6+6cC
RSaaEnRqB9QtFlJZPrhVjemANOAbBmTSMo+OhvQTmHxmQwcW0+nj2Z5ZTDxs
F7X7Gcn6wnfwpkd0qcDVqYAtD23nfOjF2uypoa2+gW70/9hcSVH8rYqM07wO
+XNmqPA9kQ65YQAoAHu8g5Ksu8ODB1Q+5PfRN3XZiOkdR/HMjnXr4dgXk/Bg
EYeexjmtw5CfeHoCha+OmijlShA0lz3By6wcz43jTv9YChcjgklsr5oizBeD
sa2y/qn3gX9lJFCJS1tCM2aXnwtRSipiz8GUDp20BOcBNWLbeu1/wh6PhP3w
OISFKGhwU1so13/5t1VjGnuwDS7vWsYr/tTvUzGc0sXY1fb43HX1oBG7Hn7d
BZMFiRqYmkQr2WfWLQolAg6ccS+m2QB3uzcliKRpjn0JeLjeyABxKzepcZj8
L56youpBQXEDL8Uz17tOZ/l73II7Jjod809dFwKv371pcL5HiZb5VhsepKNp
8B+q7fN1KIDQREv0q2kHGEN4AGACm3HgbyAVWZNQPDKelqQRjYrQCdbCeOu1
NbOGU6DB7FmY0gJ1/opcBYgFU6KYvfLR9eXEUptA4qzVK7f2tYZpIB67MFFC
C6fkQpFtVnbyd7UILoK2E1EM349aYV3HhK07PHgKIJhO6OcIstzB4q+Gi/Ii
DMN8eB6DcTH9q2UzR4qDXnElO3wCYyGyhCl63wrhqkeFiuoujwQqy6xWWoAy
+5oCgCKP9H6KOeRo1/WCE57WVOWHHMuPWtKfbVs+moTkjyPvxW96pUgg1Hct
nfkp0iiSG4X2OiIZ9JjvIQpYriE7BXw3N1JraZn4y13wJ/PFb35hJX3tScwd
aVCnST4TasWY3NcQN5sn3ausNUugdKou0C9OsLcckyjSUuROljCXK1ldiiP3
uVFcbl797Q9Zv6LGn0aJlVyHP4yworJYGG7ik8P0Pm4OyDJDr9RlddJFbbgo
wKPKLBGmcc+2QRJkgB2Nz04bhv9r5mg1SZG8vg+hFaVMzvUOhTRSSoZDDuIl
k9zG+IexoSTyMmhHJflJqmjBpFr/uMo9J0i20o3SsBnpQKc2hxKaW3sqFVOS
b0EvM7cughXN/8oGLA1uInok1Rj6xUow0rOwP/gBn+gQM6yoyRyvTFVu7fj6
+VrMw9tFzJW2FVmeJvQSHpjlIaVtduJtrrSl0PwdvO9O2GPR4oGYcuJD5nbE
AS3iBC1EO96BR9dJ14L4aZ2U1VYOjcVsKLiaBFht0gcOd21Utl5qZ5DKe7kI
yTcg+3au6Uos2/gy++Q+P25MxAkOfjogxgLDswEQ8yhY6dfpjgLUrHfoZDzw
4GyhuT/gwftNICL6TiHDhwawhQp7xlFt2sEcx1VdtIb3eAKo6Umt60Y29hFD
rgbrj8q5vK2k1HQ+8OdpsoziAmk+c2JpGveXjsYoZDAJzplvoGyUNUplWQV9
khBX0v873ckJybMM6KCX2SXAwwmuDM7jVCvaCGi5sC2Vklz6BS1OXnjZso5Q
JW+he9cHzRdjFANzO8PCfkIZYToiF7U18ooD867OObAhZ9mDAPfREHuvTkdE
S7vc319Ryq6WpKMItULv+3RLVMW1LpsbcPX0a27NJvnaYXeo73kTLvQTvN7O
1sSCuChsAKFuQE665rjRVI9KImZpcN4SGD85KHoYW9WxoPlUiser6pFzqRg1
2yFZRyM0py1c+9yYMRzlRAxxXWQoUzWraYHFI7be12iyHKDn//UmjrmmYVJl
8mmTdsi/Xs1kULGcFVGaWe93omv5B7GygTwO5NxBU99ZP/SAToXFrTNQ8W9S
R2Rdh06JH3dCJNqtB83KgFIzcCEPYdoZi5bSpYRUAp29NPekVHOqR0EqpTQM
sF6KkSoafsi7dhmaPcZt2yhbdGocknsONnvDetPXadDUZwxhQ+ek1BRF4me2
/wzRzV9mjXGV8rP75Ezw7g59w4bLRhyrpDy7lYMRtmrWEoN8FjhWroHt3xim
9aEjMrFOEWt8pe25HyBJrlbKa1P2NcsXdudujnkWDwt+C8OxmIpuef4wMkad
bXPG5VxY25DfjdfMTSEGXJXbzrfXUc2EaL77yoVPwv8HAbyxRfOlLfajq74/
B6cKJf2GX86th8Gyp49uxwNFEHFtGxIsJxHe/ucZpZzChtzbzsiI78pnNLKe
X12hXrGAbcBoYXHWO9/J937q9PZLLEh4d9L8jMIpx9py8dvBt+Muxt7++MJD
FWfonz6BzTRANdWWAFq2gRrp4Y/YHFtzOv5tvGmMUrDQwkoQ5BDxxgsnPEyb
Zea0fDJd7BIZxfAvxRmAde2B47+TD8ppgXbixSafaq9aMnI7wJJPyEkADhyO
xVEJwsLPc+wWyf1HZTz6oasnRk3EctgPYH8NVlOo6YKSCdF5WEe/EBVOHZtx
corLB3KegVtbRLOYZNMsZAajt/zeEip9HfURz3JWhVfyhR9Ruqh74SiWbL4N
20qaqxpitPrJGokjlVJ7G/AAXv0c9su1NOaGdudzFV5z8JaxLCKKEuk/rfMM
V4uf2f2Z8WBhPOveNjas1tI17DDRv5QdA7OJgJKvFCRDmRs9lZI5j2W9kjgL
RKr86YK6gvbQAtmPV8S+bXlTCuHeabzAgL6qgLz6Wuis2m/s5/bG7nYh4Q+N
aYiCx7FFreZSK+7+OEEkp1jMsIkMh95v54FK35tSocA5mgtdbCXACqgDLDRX
W43pw7egs6juSdXavAwvLfrt8a8kNKkSX7fX3HKqLlHE01OHGu0zMhlChXOF
I+9zv20Z7Pym5F5BrTfdE0CN0YupEgoTZPv0VDoyzv6PWQ0yO83zpjRgT1gB
6smvzfbrl/f8jCVX92p2TJKrV83k0dUfd90rKRcA3FNaLwyKG94CSfBPRois
o5M9/ysTWdsc91zNwmXla5AZA6e6a6pkIRgp+4tHbKu8bzJiWEs2PWYUA/JM
g8jDTlkNNzliNE3v0SdVhq4R+VGcOJfellkWcvbmZvZ7THYQf2x7TjAiI4Lf
JdlRFI61UWHj/wfeBFx7jTvbYoHmHSOGT0pMHcK3Ji1GW0ocAp5r3gIDYPpQ
jpyVNj7xUFyRKKEid565/UaXZY/i4uumbbeGx5hodHl+fpdbvGTp3w5q7W+k
Xtl5D2sbpSCd63O5O9Jl0lKd4Ynp6w9DcxBVGKPnqNeG9MzQ1rtSImcMaV+Z
+QiXEfuHm4xzrH6g0Zrq6qXlg64UxAlqOweUeot+kMS8UoWyboRv4noUDbHX
tLo/PHew0NQo3Z9g9dJzP7TI6eY4pRJANlHrAFh7k6miDQQ7GO7uzTGC2Zv6
/yukDJtQNvG9C0DvDUCFJqfcohp9Z7hX0H/lOxHhMUnBgNaKosye0tmRMx+H
vrQrU2ugDlK3MxxDWSubBO4JytnjkmxixWGHT7oQfDteoZ8Zh/T2Hoc6V6lb
EJvcFMCE2g/oy/edBOm4rNswl4+8H2kEUr3+QG+jv44Ac6NsHi4uV1Z0aEjn
VLeP7LB4yDGP+q3zjVecqLH93L0uO2hZs5PZcPjISNTYR2F1enMSdMIjiKi/
4U675mjj552V8em7N9+2HTi3k3BmcA52zhchRPRHlcc60S18rKxMnRgxI3es
qT4cjM2CTjZyYy7rwOG4cr7RvAs1VvgdMvNL3LsybZXuJ3B0zU+tkxBFL4p5
VDMWIXUhyRTkGLjlz1FOy5eeJWRqQZjn4G/Z2ZY4sycT6B2v3fZVetRyB920
UpqolKp0Mjw3/+Vv8RwQAq/XVJRSVrwpcOZEwkYNSOAtYzibF/ql7z2A18Lx
cOGC6QSyt6G6awgIkWIfHJGaOUDbFydPvTw7GC28NMy9k0GCQJLQxMwQ3R6R
kTOdidQwjpNKJULz465tbcAcklPPc0Q4deLtHnxDfDGT/eisg9SsqSFblrd2
/YZ/3z1G2ST5UxMPyHSICMD7cj0Hesq8jY7DV/Z9qhsMGmrj69tXRkHlrAdQ
h05zdWqrzH+KSgz7HaPb7J7MaH4hoo6PSvQqDD/LkhrwNwCw9up/5ivOMxHI
6nlUzUFk81ejKBSqZP451A8GZhPv1e4u/CZ+VlzKhRxAW/LiidO29DkKdC3P
B4hiCndQMRUD/24WwQNRUdJk3r3qbRADmySVRQJpgHwvkc45c+YYLYs6tZ0y
YCqU23KDObJK7d3WtBww0w9xheO6zeFRMF01WO6eiEx13HHcXGpD/OIyDqfT
vlDRMLFSLeukboSd+S/PNz8jbJHSnbXKGoJL4+swUEVWegasuR2CHS5NiTdh
MYtoM3w5FQAxMs6CGPzmoDcg27AP05YEHuEoPnzTgb3Gu3ClhMcorrucYdvV
E87sLxR+/PkAhRfYYhHWC0cPhDzLmghIg5wGtC/+N7pmJ8I5ZhBRawY/qlUe
cajRxEsSJPZ1mBtCebXVihD1AMAJRFw689nuEgUZ2bhwvrhkDMTzGBqrfN5B
/VvI/qRrueWq+P9Iyr19o0rQFzVNoAy1qibCFp7YXkkpu41OgOh7A8PGA1dO
HaxB16oGjLvm5F9RfP1w58RGdyytP6vO0+ANXYhLAVYYnAjd0dAxUF8FPikx
wQZphzeH31AH0Vo8wB7HSncIjmTxNp1Hand0wZeKCmUPvO/L5kHxxwnDj/Op
ThTEb1SuNw8w903hjaSEITOX+AwZ+UcvaYj2S+zA0JEvI8RTLYrUy/IseFoe
xSenObUhQxA7NbrouUNjjaxPKFKPiUqtU2q1y0gGnfGrc4eMvaQ+xA8taY1g
3QdVQD6aPYqgaZsI+wnNbSjtzd47Cy3khZoV69XHCnepC7R6wXVa9MNTQACd
4h8RKbgRarPTQjy0PjXUNRK9jq5fUDotwmnrTuB3L0zE4Jv10hTAcUuCFQIC
f9XGji2mX0yvZXHfyDuOvwJXMB/cb/y8t7GUdBbDaK4M8maLp12Ta2A+XYAi
kbKNGgddfCw8fUp9B4DgYhwr5b7lpDbs9G3pbx9oqxSNuIgJQAsZMzv3fgWx
lgdMECssjYg1rlssdiCqMisivu6Z13vZz3K5xEEVAAalpgC3hbNrhCmgbIhR
pSxv2jusTqxJJ+Kkb+A7SbDHjNYPCpJG9zInb4mBA9ON/thz+0tkcNi6CpuZ
jWniVplAT1w5Z56aDz8M/Seuxtem5oAX2dVpq2O/IuuEMe7L4DU1qJo8nTz4
qcMZWx4pkEj9fZOB5IiKwOmGJ3ijdWGHnX96J+DHnuj34Qxm+B8IrxTxFahL
xFGZTQ3J8J1RTnIk+Q86LFary8jVIV5vlrUHNPJ8YdH7hYBlCY8qMY9cbej9
arfmNllmb84ZTmZKknebcR3xSH0FPW7juahQjCsp+H+GLLbfIuKerGlexh38
qYb88tmaOH5QAOY3r5XvmmBv5B2RhNtKDoQ7Gfv+y9apeL9eHZcbqVB8f6up
9B8GRWUG2P7eyEFnO+bc/LloVJWOgttQH95zifMpOBU/gMnXjF8Np1pDvula
AQalXrnzqHMQNJW0qtPI/McBFrEBlIrYsOUNx5rEXk6ld1moW8ISrxItbF8g
PU3pikDSjOe/XP7Vi+0rb5fTE6ujXEktksI0wnbzYl2hmLot6h6WKnKoZWym
8Bf1gmMbxYSDNconx7Cies4jpbt1AvfVSbWjishzQhoNfs3q3cULPN4IsMiJ
ePNSViqgSea6u52gtzBiyRkVuJhHiLwOR+sv+QX7ffeVWBmSCUNGkrwyJc1j
NanB1Awh0qicbKtqLGkG8wB7swGn+rkhfZlytDp5c/nTOHKAJvS5Vm82HgWJ
26iJGtVNsW7qK/Gv24Rs+PhQVwzv4iPLOnA8lhSlesKwBGjHaweCzWfx0OCl
/xOMBzZ7oAqs0R53aTCa8Cws5qzeO12qszJHrhPw18af9Eiz3j/YSxE2uPZn
j/KlAHriSuUhuHOA8/s4Xk5NNZUipC9YHowXTtr150gXdHuTfbuRq55ysDFg
HiZz2q6Mli9+c/snbUD2Dy03efqKM4gMivGgqSi4cWmGX4Xi/urj9E21D0Tq
PLjamVHc+LcjuEIWgdnYM3Sy0w+4Dmb7MVBQ9/F3cSE7lwr3n3ToePWd/99G
eSrPhB0EXYex8mG0hLvZS8T5OHXVd6HtdjtqMZFw/p2DYL2xURV7SeZhN5/Q
0My9jfaYDe5s6JyNXrZnfGQXvvxKHWcpjJNNKB6ak7O0sMl8PJB5iCIbCqls
2iCOSkLdKPlnxFWaYiR5d5ZyrHa26sVGTV3MS0WPD6I0Z5k8EhSh1zikk3nc
qm7YxPRJCiggPmiXbU62AQzCGc4HL+laZF0fMYM2SBT6BqBvAlpsDhHO+bss
U5DtR4UVwC9CzEoLRTvgfZ27MfE9PJdqqjrMO8uf7nuxi6MoCIed3lanZW+F
l+umdwIEVAdJ9dqUnBUWEmllXgb/nYubl57AjX8cUAzpUnh9hVSP8By8LUw8
9RBN3nh/AbrvZyXV0DTpLjn291JKIZy8ZI0K8vVLTCbR1SCq/nxOng6SLGre
gprAbJ8mQP8MBxfpElIRwY9dCJ/wFizBeA/AUCDmx5uEvfghYY3L3DOy8ldm
EbfIrCzq99HhAE/F3SpnONfkSAvUJOut2g5w6eN4DUY4gW6d691ZihR97OBG
HEhr/WMxY9ANO7tCMegUdBlWTmP6Evt7+YmCeGX4eVnl0pgBPh2TM3OO7fnN
PGjS4rqfLvXYDGzE7WrKu1ufVxD/mkU8ey7O7f9HnqHrNr70inzGpC53+BOi
taSXCUX6fEBGUqOxs22ogva3RrU+w5Wxxn770+uhaRmHlBet/BqT4OcyM/+J
5ey6gDSU2s5X6fdqdCZK4wKiG0HD8x2u0mgxI9Q4YzHxD+RyYcTYLw9TIuiQ
rgJCo9Nmj2SkPBRdVaM9wONRXnhROlYPClyFVUnD6NDFTI33HmrObVk8z39y
B/ir/WUJJ/x78Y3SB/etUyjsnDBbIjzYYSD/RRBL/0zhG1Iyt88ISPoPohEf
8JWAZSiCZtB0k0ERv/D7fUHyAeQVimlo5OnqcduC/ewW5ERDBpTDBHtRqAL1
8ZG/o7M84cwLjO8IU4znh5vGRC3VIbTwt+BuBSwZUC3rTjP8s2nguW8jMr3n
xsBLRj09+6nXHgY/znVryTAbyq3ndGsg95DuO47s4IawlAVlfryeqqgg3XQI
3zntvqHWXUEEqHcPcckoLTtl9d9os1VBXA5o8lmJmB9mtmo50ndYz4bjI+DK
NFwQ5DE6V7ODXSjCMtdHFkJmcdTAH8A+k6aoipgBKBgDggo6x3S7U8n4xfnE
ggE5kGaZUeusOxtdIZWoywglotap2kyc6KA7yYjwzhQ90bybhiGfzPCqUX5o
M7lEbZ8KKKwfq8X56bolvjE9i9n2skfsrRj3fRGlaF6S4beSnJsOdx3lII1G
9npjp0J/cVjvYQr3W/lv2YLXBClVOA3ZJ+e28dCxIm1VJYG7N5LQ8VbjeBZQ
Il907+gWjLuYjB8MMA2FU9TYIJ0Obj8nL9MnullftE7jzTIIuRyafWMLbg9J
AKR266gLNE0oZC5+kvkMtDCgfwECvP+jdW6ihbsA68Kke2zsK2JaNWZe6zOd
OO1OLvBf6hZaWsL1aIFkEBFfc4Ink3v3gWpH11IZffTKNTyV++QalkLxwsSy
Q1H/oRvIxb1yiiQSMkz1wAW3bIRhk2KKDd4ok8mvauUDBXQIyDGrT+ITQsRQ
OtgAcwQqRQt3iKPc8g+LuE5oYG3tRlUAIbPLKZWOKJOWjd5SgTnJB1RJu42u
MP+XlmZObZ+hJTecLHkyu+l8vFmZJhhGpdIjYa3abdWpksfZoHpgEiGIQZAL
ktZz+nrxVHosgLrX7eKd6xuG/I1roOZBemsxW7PtiNetXsYmQlRT9EopebbW
NeHlwFEnlaCUH6Dnc+LGM/Ma5jUHyKZWWh5SPSgYTftqVKaVXehr4wjSP8DH
6F0pJvlWrcpYzuClo/A/xuZCwORzWa6Crpv562aVqC5X3Klc35XcnkC5pZ0X
FrHyMERRB1YEMnjISWSHyPF3tcU/9VfsTD5KybdkgdVYdocEiCsgvflWTekl
FwM3jBgo3KanOMwTWLOk79O3TDD3yO76H22ZEDENWrzmASSFi5fuMPQAJWhS
ndAE1PQ+I025nKFULBR1g2rAuPt9cu1YPXKAnsuW5pTJZ7SV7Bp++BgEwL5w
/bH6MjUEnSdDP34SnMmYUthpgTqLpUCYQ3R6eyv75e37S+xR5oaHJxXSpDW9
YdbOeqiynFM7//ycOArWv3L/HDX2D051bgxwBpOuxzxdKfz6hVWhNXP2b4AF
qKZk8Y4d8WLwPCqToTcfeRDzDBKb5M9MPEvQd0FAu2cA5xbl8hOuD6nfoXcp
KCAMKdcbVIsJfB9t6P7qj6I79XTRwBxVAC3EtizkMyzJlBytWOBs8cJWQoQN
kbaHPU5BgS/rjD3LG9k7SUvyz0CaqRoXvwtqjM4Kyj8tSJ1YzJ4AcJUyJbD8
rcZnISiw3+iGpl75uqVMZm6lHi3aB7xAd1NsTitMja5jW80DDQoZf7gtO2dB
UON7g+estK0E1fu7CzFPGoNuWVRDydoSVKgXBZBepyVjGNNST3J8x11eCzW8
16+kxrx9Bju+sCrL+R2A1ST4isacAGyHPPaJlWo0tV7hcMkQ+WoxzCOsRSwS
8dIZCvtIxD+EK+w6HYYrim7xHqHcz2Fd0LV0sSbia5Odwk1K0k66OkvF9YPt
7pXXuyuHwGhwSyC7OL2U9/SaW+0rlNPCX++TUvL7XUMS3KGN8R2TNqUCFQi0
pG2hkyyAp3lelhNoRmn9P0iWid8+8JoZQSfvIM9AHs0qljJ35IV5qnoilelN
6hdnvPUNzyR2KrumqgqJuDsdl/B+84aib1WBdiCkn2MVkx+M8KQ4nbihd6y4
51qcB50FvGTYq4yrnd4L602YE40FEDig0co9JdVgCCXSGVNlpq6fgg7D0mdm
4cncW0+FNaM+rzyt4g1WzjfP8mJ2IwxwV5sg2+/0lZjfozHzb9hlcvWcDnxD
kjlS55+N2lTG50H67AawvXw3YfTYmziyv2vETSCDO8/Y7/BzNyFn8qh2K5FD
YXjNAACepsMg1rExhon19Eqqt2IbYv0WUU8SbmWDp8vVkkzKMapLMpH/FAbv
LAmMPazGNDqgfbMhoOx9RM4YMgHeW3FTof20mQLJRzwvzL66AY4bsLSK0Yoq
gg7YI3XiPfo7qf8jKJMbfMvNF+YOHDL1H1aZOUvX9orrtEg3L7UmWygouQVy
GN76ixgko/Ji2kEEfyeWaAguin23cZwAeuBQ5n3hQ9mzseE3dN975f7tqPfh
8c0LBwMxs7LGMcytE/RCh51nIXGEdvPSmsMg9QcxaRDp3ckG/ly3JvLZKWN4
e4C6OzVsYHoYfRQ3QlvLnXNZYOGA/91gzecdnAeJzKoH3Lqj+GcEgNA5i76M
PSNJXtqqes6INSZU1xa1pcfWH4b8VeOgDRpyxFgtPb7LT8lz8UMpVsI1z7MS
bkYtqzPniqwbtLtQPHxosuAl9LBl7Cy1rp7dzAllGr2jEtjPeyb97NM6M70K
jzaNQws0UqdCxCUY9Doa6NM6yZZUDvM72l3L+VLTdnq1mnPca7uZYRPm7xts
RatZhHwKcCL2MSwfaTKnbsGzdqLIZIQWeGbc75cOF+9mMOtfYoWw1Jh5xYz8
QBr4488WecAGoHwC5dAA2lY/X3B04aBlZ8MnCTFHRWUTFYBBYUpWbZbnU6ot
E9holjgU102YgXTmBnNw2eklhJrXqNGbGsFR17tUtBBTzfZLo5pshi6JtZEX
+gVQhIbURlGtrRT4oGU4W7VMgW3xY/9EuuINrafF5zBQLneFY3jy1UMu7rlV
9b4Pzas7VR0DLCbU+JU8V5DIrAqQnNMe4dam3jNrr8nS+jYsrHxzj1YLwWR6
PEkwmg8jk1+XabgbpKvgmcKexwY1nVBu4eYWNJVFo5gtsqYjbf2ROGQkwOlt
zpCD6bfNc9KmmfzVHDxZgstPWOOr+F3tQB3Zapf9R/lapd6cC+1fBaiB3K/Z
n0hdIAZ3AWWLLworLrwZn7qEY/Jft5R2ocV/LoRpRqDmNoujk/qEZ8Kd/sBB
1VMo18DZ2HrAGGcEDdjZNkymW8eLGuhX8/zvjWmjpdK8W3q3W12hT8m4Gc4D
PW3N+eCX9W5zEOZvWvCZAwBCjNrsfhPtij3KkJR0IiauC19P5flM1WRfkAAF
vgtAaKjL4Or4lNCxcNqWSTjUb7UX4Bgsu/JdsYhEcs0a/Z9Yk4egYvLT7XiU
1vb0nEKIDBBWra1amu+pKDkgnCFKK1xd7dzIiIqeNt06FLEE6IT9ebhirbFC
skdHNQ7M2vls6fteLiOyUcbeodVlJFc8Xlqc4TYJ6Naa93Tm0ihDyKYC3ZvV
YU16OQePlyWKE07d3E0s2I6iBADe0GfPUAFIvw/RbAXQOet1femDYKiaLrTH
M5o6lcDS9KRNoQYesHTUbFMlbEWExPLzsfXgI5niAHy2jbpyeDwj+9rtJjNU
qrjHHMmcKDdQ8n1eYJNhKqZVBXlu6vEf//9t90adECrvcY5dd1I7WqKS5S3P
SJGrFFhlQyUlUT1tfsMjFBiRJ82bNz2uSbMG5l2EhY9h5rRUQooWPJIe6VbX
65unqQVhpNhlzlCUE12bSTE/WWxUJztJvmX3VEHHaGkieAu9tK+Ffk9qYQL/
BSRLU/xO7q7LY/mP1WqZk49uIJRXHOYTTMVSicKdrG/lPulIMCwZgYAtqPjU
FbGQtbPYH1tpolzxKADT+Ec8G64iRXV8aZCIqKL4ltKK+9XxtsVMxcUXrL9b
Gz9psnWTV0gea/R7fuo7waB0yPcmQQ4MtUYsX7TQ9VR/SiYEdgmDyDA/J+y5
pF0HBYGSuFX8B9RsawGrSJHKKH5m1Zczrp3jkxDgRDa6ms+gHjESvqdJN3eM
63tI8YysB11ISxtrfkD0O73XY1eFLuy1d+InJJokaYLxycetcKPWrWg+o0n3
2L6S/8pYNYWRaULfS/NG1nWP6Pm9eVpf8iwV+l4dhWc9iPSqqMhNSeI2qJWY
L+BiIcff8O9IWQVQMwhnn8Jj+Vzpi7v3dk571NY4DG5A9QrIzOjo7bYkmg2D
d6bsdevx0PsJs70zMT3A0VK4O1LKIfkSxSpKapBYIlohUeZLqUKL9FilhUt8
ikDLoixr/PWtNIqAxT68FiQRBIhUxnhisNa1lXhU9OGgHLakZldmKzfAVdl0
6e3Hi6T6XjjSJxg/Qb8ayq1+nAya4QzT3pg4o2dLT+K+y9fGf+c6dSzjQXn1
dWwJYn7m76h40oWcq1WOAriElDARRgzyyJv9hPpkhav5yhNZUwyi+4h7oVdO
DhxSnOTy7r41MavIWtp1sNy3Jy8S5FO8qcvDQrZPLhEhkUHr0p/ViiDMzrL2
Ca0QOKe00MiwWA0hPE85KgmHfE0eVBmkNFDiEldKSBBNt2Pw62Sf8PBjKcjI
3/amuSzuXSDSyGG4GTROXnW1Vg4k0Rngd3AhIsscj5PwkjkQ4FtimeN6tLr5
N4uYtF2EJbaPHnapmLO1KyHMdvmISpMOc1FdR6/islDln7i9Js3ipQPMIF0P
hucEsJ96t+ShEYE5NbYgpkgZAgOeQTsoqFudQWw6LDlfafB3yukH3a8LXJCl
2mSFZ1tcrZqhFYy+KwuOhuSA1/P00YqK5OIiJOYhVy0T2K6Vpq8loWzx5SBZ
yHQV4biPCuM92ivoI0e40BBnVCKUQuzk0gpaY2qmqsPSk1oY8oyPVt6pjZfO
MnGjfvcF//Pb2oMHpTReLqzxoOmWb1NaEL+Gnbo/OcTAdc2myUsgtRyUf9zp
DnvdWOYAXbuLnhhh8ckqge0iIJNS2TSjpPY150Pfc0Fx+ZIHCHSGAmy72RJu
thHTgnPMzw/MdZtzaqk6bIa1/QyMKuqnH+muBJ8vydMwZR1OmHYe7XvnMfB+
52g6AeVzrLHAxEeApG5c6uOwlXoL2Q9j3FN11JkL1FfEAT0sF7q0wAd1siVv
ekSEXDuxcayXyhBvlBa9fubz9zgXO/+wBF8yhOEEJkwYq3323huOgxIjwAkW
taAucN4e3X9Rku/+X6EL7HHQF3hFOgTTyjP+T49UGwL72pEEfCb/UoH/4Sg5
dwtW4Do+8jk/bmWZc3z3FsfE0TkSeUk38mt1+lfZ5PZVh2ww1IKpbQRn7bku
9YR7uIM6YxtkRuUjQomtk91KOzTDKElYOObNVoODDz5qY7ZPKJif+wY7eaxv
cVkKZJGwwfdzlxmgXlRo2IUEv+VCxzzX65ax7nI4rKTZJW+AH//FLEHa4tW+
0CUgH/AHDMNAUXRMzduP0ciiP5gxnQlz26BtCmwgPfo9B3D5fVnDatieIBtY
wpnnLRVckBJ81ju+8ESgit4hnWVUbDmeakbKjMUlgtADn4KLK4dZmGe+kgkZ
N/l12TtXhEDzab5zHbuju2XHVjzC/pJ4G1BdRB+qmJy6DmdJzZ+nFOC+73Qy
VP/IuFxXBVEQ3jSTh8hiQmrgSbTR+gCquMCKuZEfxTxu2GPipnc7/cx9TeWL
6dItt1mZjYZZEZwVaRmyr3DH47Blx+CWpEWtLI+HYvUHe7eHLab2p3kplXxc
uPiF0ACR096dcTgyQ1IO5DM0rZ4bUDubkArKqfkX54FcW/VY5njRbihdckBY
F7B+HDq4GlwBn4xD2Na1GEO5T+T6Qg46yZC5c4RBcLTjsL9uWacO5on+GYcT
9i3fVRxOQ9P6iEpGr9tH60yI9PlRQVujxdzEwirBeAQa9BJQ34OAIDcqM63m
HhdiXT31bEVva90qgushvrxqL2Y1fYEWYn/Cn/RwkNQ9SIgM65SwNGGiruGP
2uRO/94mOBIBuiYXypRSNDjoP1wRo3c43H1IgU0JAi6ZOExmMWXVazo3BRZn
RBDzQ1lnT0WKlwcRB05GKR3hymbCvddz5qE2saQ3Y5x2kgBjFXlNPWM2BF83
fRE+xDEav3/gNE5szekyltJfgIIHLx6iNj3l1W1ZYeLvKdQ+hpheMS9d1PXG
rP6lug8QAYMkR24Rj92xUaAhz8fzwLEtdT+NyMBvkCa2aVKSc23sXHW8OmIg
H0oEVDTL58M0QSKAZo3Nzje+t3Ti8LJbFbnsKra63SZ2qjvWanSFLwZUDzQP
2pT1p8FgnQ6gk3WpfY6C1cVK/HqwktBcXI5IOX89zg3v1tnPk3Y/07VPK2QS
hbsIenzWnglerOSX7DhxaWVAsTU5CFZE8NvdTY1jlHR2jR3UALZ2jPiUyFxN
3AZGHJgASPvWhjLgkWp0mfundCiWuBfom4KQdarT4XtQQn6THVSNhXqHqoSf
hmCN/rZgpn1HBfZs50KdF7jmn2eTj8MMFM4OWIWkB8Uh//zY/EuCoP5CiLVF
pZNZsWgaXa0xMeJ47ZIODQHHMIEjIUdNCY6K0Hsrhe7b0x38hLQ2oUO7IhtJ
Wm8k//KTAT9t56AvcYVZCTBqXFzN5+RuXWTCxSB2UzrW45MDh7ZJdM0ku3TR
Nm4AasQSFjFU/NgUN1yrFmw2jM+KfIgZhQu0TI7yFLEEW153hvwn4UZqAdwV
N2EiA2rPi9LpMjoA1OMFzV3lv2gcHTfm1LsTBI3O62VB/b1hGalHeZ4JL97h
3SyBWsRnH1uf/WZgDBUsMe78aVejQ2ZUHRmdjshTINIOLqteisJrxIBA8FDc
RDtDObu2cbrAQ7WlhkNkzQ8tCZQjcUrzn5vDn8ZCxjllJs1gAiKCGqsBNiFQ
DNwKEq9rfmEj6iMr6UabkymS+vM1LXlDuuSwbSyvfocFQfEmlMZPoSq/18Uh
xhp8V+TDMpoyFeN9rY0R3JpszJ7uwnxT0PytBVH1lEG7dZC1wWZ0o5y7NCXl
J5BzeduczJKTYFaz3VreGC2bVCDdUrdXDGqVRQaJ/O8gsENFfw79TSQFWzZ6
y93SSU+feLlLWc6VQSnrSQI0TlkXypTuaNOkQbh2fLyZrZKzV1FBdIzrX0+y
Fl8w22XO7ySMm+fvLhvG1poE4ltcIkcmOTMGxn0ABEoPJHDeV5t2CNmZa/i2
3ajKBE9GI6qVliuTE32smGGU1JCkXKhzlD3dRHBDgQWUaCV6qjHONO5zysc6
DjHXuWjK8umrmFqWez3Mo2g5hKgt7IkbKMLZ267zsaYh6/SnddJxh0YuryA9
KNScUTiV9Qb7b+KVPNDchEjcieVjyivTRn7krnlk/KmGG9Ekl4iHfK4SrpAN
Dp18ollk/u/WzomAkAyG4SoJlqYTBBDeJZj5Te7ZRjTNTGrVsKOEZzm7gKLK
jpVRL5OUXEEGKFdOa+xRcBPmza0eN+zKKwj2WRFB8fys1bMe0WXiMhN9Ni28
wPbJ3KLsKJMpQ17jH4QyF9phbO3f6TwyhBOlbToI1afP9jInQI1mgqM7v2uB
G31w15CvuQcyfcoS10NyT23aofqCcyFoIdwr5X5vMCIVA3GCrlRJtfKs7hHt
2T7O/qKFPrmjzjwlWCyy9tT2U0Xb0F77HMxoO+sUfXmP+cSgIixDIJViflfr
fCTeFnuGpzvt1Ou1K1qN8ag9OE52CxG0QsuLyG1dGFICCCAFPUEved46SbF4
ML671CzOI1iZe44s8N9lHNeIjowj/x5RhNrLjLEMkPJuUSg3/XFlDrn9Lm1d
igkuKtl5ylSmrKPCeG+QKmtQDHKTW7bExMrM7XYQCAWegn9kCFpr5E+m4h1v
dkhxsLgU2INDjXN1ChBLyFsTjC42D/UkMTU5ZIHllVoWJZDE8i4Xk2/A/I3Y
VBeRhN8pmiMbQtI5G5Szos6T3YPa0mV3PuP9n2xvJ23IMBeqSjsirRhpDOuR
+uM+sCrY6ODZie9wOAb+rjqhUPondo8OIHF+3M6EBdbRFUZlxzguLz2nuSCR
llpB8RGJJFXesQuR7r8fGvd42CydZis8WaMj0TqEwB9OlbyrXLUx+sLzkbVU
Fj1g4q9UhES/550Lv00eajutGS4ZRmvM/kELFDdcse+Apit/imx135sI+M2f
CouxoOa13dvm4t/jZQGln2VS02b7KsIpNe9uZUGROGvR6jjiHmE8/wudG9qm
GHtLLaSQ5TjEfX6G/dlUVLfiLFBxp648gsrViMmng42+5ALFENMAiTB+Ig85
zsMZhcZXItwq3EcPAv1rO04S6MCVhaEpjzvyRDCdyHSn7+gr64/z3MWhsAJF
lyo8iyKRmNBEoRpkyva+b3z4psHsqZMuHx4OnyK5dCcDAoQ1/wSIA4nrMHnb
V+VuPxQ9aodUhg1sFiCTAnNsaKvhXrA41iaxroh1uIY31j3sLpFxWTyKgPHc
zmSZQZdscWfW13sF3yx56sbyzKdni4t5CKhWFbLdWNfo2/jn2BLF6Go2GNui
PoBaDH1meKQCQn1jCrA6NtTGuwrwcYq9IJgTnRbdoaUs9jUO/PnXw6me0vZA
wvya0tCCFWO3VM0YldvVFRiFC+gZzfCt10GwMMql/u0kF+yZZTiUvIKqEKRc
bCSAtaK1/nTmVo5z1qQCcR/9os4Sqa9PMy6HSJaT1PVTWOdFB9UT79mDy7n6
xRlgoV1JcXqsEBeQEunxU2cMnURO3jLzTiOURbso7+sfEdwiUVAeewjfbrBh
CiToGZeAzp/QmBSk4yQTS5ZH+orgXeZQOaKOwmodnDXhEDKPYncZugcqK1ks
hqk1Mq/UUu1L9nuT7vMOqzmVDJFDNo8AYFeqE7ApUtfz/g/qQIRyJUja1OlG
UrpVmpDrWN6xwT5lFk95T3+ApI/DbpXPOwXuvm7qnzol+TYPSj/3h6+k8gHd
aAAGgBfNMP+itTqUUz3h+aiW5d+1J+vEeW3vCxHQQqoLyh0NWtMGS9I9axYM
AGYtiugh6wmVL1XdGc4dJ5p8k/drC/NNB+Sn33s0Z14b69p4BsOcnzGY2itx
NuJ4ZTGjSrE9v4RkGQCKUaHcdk2W1fkH0z6X2HH2tAT9aeuGzo7BnUmlaJPF
5FL4QBSo3eZ0ms/VQTldiQ8L34sPRkM96HsrN4yS15T+0H9FLR5YMm2UXjeS
0qL+LqJkmmVRb1I63+UtQJWrgcszptblri6MxveCzZq4uTrd3e5QEDw2o001
s5qAkS+i1YMhKmC4oKHcXjYD2sryh8QwbPMQ8y8IHerWjb3YKba0pTMQ4viD
Bgl0RD7jwKMvV+cbwrbQKRNDybH5e3SnzlkUfvA4OWvq/FPVfOLxIi3CpJV6
uNFUdsegCXb+nAE9OCTs/UY5SK0HPDcymTqjQBD3w5vuHVl4o1BvDP2FQFv0
6wegaRd4oL+YB6x3wbBxEZhB1x6qYcYgmEgTws6dhugyFt5aX/BEeiebgB9H
v6+r1DIzXH9qrpp3aGBT3YDASguNW7FoH9AIkkjRKGTuQ3TIqfBx4torKfy1
GaiCPOyaoi2/iljzoNiWcNn8kNOrUnH0PhohpFjia95WuL4qsnXoklMSX86X
idhOdMdujMiWUpHoHQzLY+TRVQYSUEZ57HPuE8x0mLX6pB3wcnv77tJUw+Oq
k5yOY/szI/8kAzAQX/A10wFm9DoXKRkr3dhaBU637HP9utny4KjVaDlPAp92
LmOHZBaelAEcen4IMSE2Pti0YFE9aTO8qzHUZ9gst66IKVkx0rVi9hO9EW/t
olZvzuSxWNiZea84Ts1Pt4fncXcfH9hrH5YuETb/65p3iN/MoRF0QChq/OmJ
TujjfJJ7vs76Q3pmx1EOHZLFHADCcxApQxuBa05bSXvVQFWcZJfZMneBYgk1
6nBgvbiPZB8900mfUWiuPgpdKhQ2AybBAEZKgxhDgOpnPZDYT8wCV1i7T7gC
gxZdOSIHPci0e06w34CFjCa4WkGhWO+Kw7lc3Mkozuy5PL022c8gI81cZIYI
BSjqXiA01s8MgBvEfvAK+61yQ/7YiW90uw03p//fSwXvrutTFqbWZHfBK5Gr
N2JkzLPT7AVkTiKgpQXww+JX4oftGHB746yIXe9K+7AfeyU/sHnPUGOr6rBk
jml1/lXzQ3sUYD8ryRFSNVqm3ryWxd20kAiAVRdYD+28QqUlfObiIKxhPbAJ
IqGO4+rzbTcM541r+2SOdR9h9ojnIjPD68TABoHTz8FAe5wf42u5E2JaZ+J4
UlWXg9yRUbQgEHk/xmlxVLIPAN0/iaAK17QjNMLCyx0ifFEaHMQrMoNiUh5P
I+/eUs3Ug9eOybTWrnwuYn+Jx4xyF8eBMx73dWnKkp41c2i3PXEngku6UM9Y
lwq/DndBztrWmCQnYKl6GGlMXgKlF0jmcD2WhtaoO8KBewZ54dzA7VHna51h
/DmSl5yzvtZDdJB6Yk+ltKHb1/5XxIdS6cjrLoiksWfrqLK4M7ooE0f7aKQm
5t/5alFHI7Rezg8ttE+aUZNtwRQln+D0yij3AAXi9Jw5uSuT0AujTMLs/tsb
V0Zokot0RKGVroBIdQf2WdmbupLcJsSKg2wYfA7wMr8KLq+cu6SbhLjyA13m
pIvCsT3j3ybv2xJnimEMlplr3MstHI9NRV+m8+UV5P3cLN5+///PmQLJbEPN
eB+RqwyuY7c3Gp/xjRYazRMIXHJ8rTcFvLIcDa/pAsnDEqpKhJvbgOrt5Fiw
/aN1iT1uFHqK/d8KowP3TMqNlbWA0v/9cdC7pSy4ph7KNFNgvfeChMXoA8D+
BfNJ5fHY3KPhG9HGUVKnTahiy6n1XBtgXFruefKH0W9iI8c1WetcG1LB5C+x
+0rhYLY5s3CqoNyeq1tHtNbKb2wA3D330B1LedtKWl/gm/2htBT4T1qThcHZ
aUD09Pc/L9wW2r2GGI47PVkI748JGzqts7Uey8m3hVmdh4UZxTVQ2/BLcgsu
HO+f8P26D2ZR7zNgMmQeXL+jGM6z3pNtQ7gFN/VEPJeYeX2SuQS8ykDv/4xa
tIkhneGj5a6fU66f+TuESj8k+twwy2Zl11dGO5fRoviGnQymwAaQgHDIIxpy
rUr56kK282AUjoRDOM3x6j+OELu3UhgYAVjiVfNNJ0PxDqBpYNvRm8mfSqQk
okVE9PTs04yneJMMlvtZmeHLbEGM2DzzAPn/Qs2kXrhogZEBRFeSlJaJUxL+
+FjLNBbgbybC/LjLqjKaJvzfU6JzkIyFKadeYz2/tIxntVkRU7QH6/ZfJ5J5
8B3BGebXa1ba1vmbMAOx8htbsnBQUNlfMxadMD7JjEZpGICifcalVrJGEglX
2uLA4lHLLtA4NzmtfgO5gt78iQ3xqXc3DfqxRkdzxJHg++yMbweyjs0NRhv4
ZMn4p3DeL/xGFnTiGTj9iNQ5eCHYTXFQpTbODlzVXyA7UJg1S9NkLVcMB1Ws
eKVBWt2I6sxhJsQGgIcGzwnxJMk7HUg2u15sHehjPjgyjl+FbE1cwNm9VIpG
HQ/WV3HdDUrpdXJqMvLQBn6PCttpP+f9kkQ9c0i15l3jNEANyxRjm3MX8+VN
Oo3h3FCABVIcK2r7GR8HbS1WUlSnawSIDlxCEsfvsXR3F2+vKyKQkWwZZsOP
syKkrlaQmBd1Dqavoi5gttCfx1wPvueEvVTTn9eFbptsgRZuDuHqCokH2WTk
HDwODh4+UI2yJyw7pLPP5B9CHkpmv9/rUUDUU1ZpeW2Sq7uz0NQYRD4iM0Na
2/PhyXH0deqhmwy+BMD8Xm1QYohsw+EcMxKnTulr5bBWDvjriGsJU9zRwQdu
0S+m/qeGm0KIHLL9Jm/eLju9N9JYWDv+tKSKq4I0+IA1Hpm/Wnal5aKxYRx/
WmnhoXmZ19aHkUivOdbEsC2Lr1/BC2bBorxveIXB1KBIusv404kcl9tptJTy
s5DJfhDHsG8gxHzlYCnVlKSAGCiW/CJ3qGjRlsPdRPFhUROpZlk8qP/5/9sR
/G6qZ0Qcu6001tWjmokBgdRqWazKhRDeMYQ059tXY4WMsWoowa2aXPgnr3Q/
osN1yui4TeIwrvSjJAPfDbeehNJZfCUugfF9mM83D6zJ3/+A4dqjdCvsG5J6
vkJFvhf5rOQDZldeDYb2S/uOHCqlHFGd+qZILKk63mfadm1S7fN+pDDL2NHZ
uIvtBApP9NdKdV431PYclRxSvKT6S2Y2xzFNHepA0jivvMgvFmF8XApS2ila
h7ua4cjRVfWukJmyEASjuHU6RTZ68lTnmHyfgwBn8pLz6BbEFEpZjs2ZEGV1
6W+IM1JsDcaIdlozZkq+YHa/l4gcR594gV6Zbm+RwRi7JsFtSWfCsw5bT9pH
ohCaDxvvyfEmluUafHtVmtT8637V28t5YS0sPGM0+8HEWkdwU6HosMYPjAcl
QAwRzpU3s0YkOFNlwSIhpr0d7iYAby83kwg9V8Pb89FLkj7vdlLkUacP+aoz
s8WJ8xiaX+EqeX9222AJVlnlpYc8Z1C9gFKjDStKHAyYy5GT4RXP42U7k6z3
EwkoankCCrqGl68lQgKku8JOBGBhUN//GimvpjiurNb9ElU75vlpu0z1d5dP
Vpsg8zOyhYodpLLAYlicufLazQmnyTEmuArsUa6iohLP8fZZcYAD00kwL71R
hwDDl5xPprt2IQUS8qPrTlEPCJaprWB2KWhUlNF1OO7Qu8j+KNChXPlYWQBK
9IBgYbchwGBitA/51+kVaYpGkpAF8M2b/AA8xOcMXPWMD3J7nbUBndedcLi/
UhvmiKzRr39mwT4nljq8oWvNRUpGGIHVLqgs0KfK/BhIMB4+lFG5MtWJ9HMc
kDSjA4wVS1sRpgYc6ayz0Oi5d/IRVu1dLj4B1N5PMR42Q3M3qg9LDrTdxQ20
r/8m3+L7ueRgl+7vHY4kCiDlNkThHJCNGbW4ZLqTnh/UG8tsoFxvNM1R62f5
t/+8wDI1W4YFFlTT94icXUDWPUWJce+yoMGY/YHBMskMZcFMtPXITiy0mecT
WyivC5xZ3BGlHFihke4NeSDPIw0uRlnemlQk+K+ZIv0S8KUjf3kzOLkPeXrX
1yVPff/254oHdtIcrXsVKgstYu63D5N8Oz4kboeN76DBdLeX++xJTqEqXOkS
6rfRNy3oF7Gk0rZo7jFYHCf+xtpdlHqDlG9YhB0EGbDJYwf7kTZi0vIdpbr+
cjTq0+kNyzI+o59pBl1kcTwLJBt1RTt3rnfwJcS8yUCV0ecj9w62CRwG0Rrn
03WNstSrvtlcWaBl8+nrcN+TnU+AxQcB7WF6Gl641eZvp8FMGBX1QK3Vzlr6
AP9dHpcjW5Em2XaXU3/t0ctC7U9pQWZ/okioDlII53vm7fzv795D4OpO1BPs
A1O1nui0swNqXT3V+6Kdx+ZIUoMw5NzE7vecH2ipfa+N6ZyzP9fQC/kKs5Xb
ZLMHST8xwOdkShKoMV67zGxtQCSsrkJW3twfcZMKaRqYuiD6Vczg8kXDZo0Q
t0Yv8FilJVdjJ5Sx75ualWfEclYoP9KxAe9UCg/E3Y9dqt1sX9AUxbv2uphB
WzOfGVH/xtLnGSPnnKCGXmQoQqzkaQILjYa+emxmqmOH16ujJlCbuOSj6CDh
jsDJ3bnP0Z5mmoJLJqlXOZhpQ5vuQj7/R3jAEGHTl6RqgOj8ur3tT7nwdETr
twPb0PUkOJzjRN0CNHw8TbOOAnRHXBHoW/NWF54vf16T9TLxswdezTmTdRD/
6aNG4s4xXLK9ngjP0jcmvj/+a9CA8FG5yyo0n8O9IaB9abW5DLqdb/XKTsCN
h0aH52tYZPxompnlw1GucfA6+R9OthkzswOivOVl/Y9Bmc2n7IBIwiM8zOc5
vIE4wPDBa7PrZGkcRpUTYCChS86d2fnuO3IuKAcTAlY2BKmSwXBaPhwt8X5+
03D8SUFUsefr5pBt+6iwU5ianMBuPpvuhAsgAb6SSDT3QfPrQXDTxzgh9X3u
R2jQBgp3p+gtQea2w8WZpTmbphMjj/2S9e+ZRfwbF1jq+HX2AoCTQth5jnqK
QQSTXsIUGeIVg6EBaQWFVMh6ea44F3fqYDjfQMdTif3FYf1pF50wKh12asBt
w5J09g4/ar97q/RGisH8xj4gdHInFArIQmPaBWDq7AXzTb04lrLAuEA+VmzX
4dtMH+a+/x5E7i+dTQ3WIrwcE4O9b9VajFIEx6z4yVbK1Rb0dhDD0UWP26XW
faV2QAb0ATauV0niVsdlPifIAH6mZTl0kXLR1uW3iML5lcRq5TS3P3cFSzkV
ZPoNiuPhFqrDEQCiKzGjQnVyXJQxVD+Go7F6FD9+oFSQoj2Z/PvEhE0fM6I2
eby/KTLTtlA627PoOoPK2ICqNgxx7n9xrlLh3L0r1rjpWT7luZpYg5zEfriF
O9v2Cg00OogcjoACt2i3Ws+dj0G60c8Jdb13t4/8w9U8JU6EPCh9IYBBCZwy
aw2s8LxG7A4cAGZMVgHicnz25fUeSrveWllcWDlnsIylkFY22/bMOV9jp3mQ
5I9jPInDRjazRvDZDTeb5v46J637zqcjkBOxAOdauzPS693KiTLByA31+its
UVRSZRX56xAkMtNHUadgLBHEpMhKjE/nK94ZHvpjcC3KAY0du59qmzYjjWA8
sdqYaFzBkPoI72NMhtRmZTa5NtWgqBUafaNr7+IcVARmGO57Z/7D/8lDvsJe
2crAe/coXiQeWiyaLGx7L7BadjYv9q1woxuzrML1teOAbcpJuA//u4RI1lRA
le8+nfrDVZe3xtWhvj8G4IopMdoBKdkdMc9yt9eKMJnJsYyYzyV3NaCGi4dt
o+HuZtAcNLZSoD71RjVdNtBsO9aJuisasjxjTENWuklA4noI8N1TSIdxt96Z
j3si1Jf9qMQbZ38kps+knpNzkIatANZQOmroGeHBrSkLxqzMHfPQ1QO6goF6
lmZlFKlAT2ANSPoOIrdUE30WC0/MkEhAqwYQyDMtFQmzKGgHRGLHIDWY33im
1NGy8KLJtmxrS6fOoMr3bRmelle33zhF8INhLEwkSk0QQ4j7EyFf6RYqMp1o
3UJVtPDuD3xQ3iWQqi3RXAPIVhT8LBmyTh4Z8VW/6akc1obZBGD8K+GmHA8K
s4QwDIKHbjLPzIlGcWPhcfaU8yE88ciRWNCtTiEAeZdT88nhNm4k9tV7njtA
xufoNMqcI6oox9mYUsOnGOku4/8x/cTwuYerCt+szI0IGbHu3XvNqUzTy1Up
3auH/0JuqoDIcAdQFp8bG3xgE96pEAbOyYZwsaSICH3df7bnIUofWaa7Auuz
01Zjkl4oM0nzhyfpOqSstIPAKNfVhx2FRXr9EAkdb544f5LLzdQf4+o1/E2B
39NupXZDhFL3ciaZCbNldLvo/UleLDB9vAHepljn1JSU2eb5c4gN3ZpfrB45
bpZ+WexizMlVhV5cxv59LiI3g6dsxyu5BuGngbt7zSO7WCdpDdIsPLL8oLo3
g3AUfs/tDm7hxKHvMHW2N6Q+KSEZw0NBGbqqB16EF2M+accN6SqCubR3u3Jx
ZPJQ5FdtiMpSBK07fvVpY2J9A4KSVSGCbOTaYL5LOMKnM4jXw6o7xNOc/VCw
BZ2p1CpAoddC7/sf0S1xMI133ru2+1XBh8Eqkc7p2hNlYWew+/7ifEM3Mpa2
1n6UpQOph/M8JkPcM3y0nMj+vhj6ubYSV+K2+MTrjMIde3AOqFZkmDwcVkl6
b5bDgkzMRShlIa9iv/hsFphBK344sT/h5b+PY0exB7nhrsrZVA3WEmEm6ZS9
ccyi/wV07/GDi5meqB2ptuerbmNN7iJKKALCZKZHhK251IhpehbNmrjEzw6N
2fKRHkmCl4uh6cmvBAiSR5WId7j2u59BRWGO1EaYeZgBByHwpLSrQud3ms+H
eoJgAnDxgjG5p5FcyzcwWYr0NADWmI1VuQoP6TUw6WMbY1lXGRtnR91r3owt
i5du3fMpkADdq/3bteYbB9J06RqeA3SMtfaEmFOdT6nS2VPAe5lE4nYsUkgM
a7yRgs3NbFXuDjNOVoDNL12Er5i+vBAoebu2IRKvb9bCS/ijgAIrComEHv1F
IgUl0YBg4O+MhKeR4qgPl1mz7vnmZ++JZ8Sf1v0rEWOSw9c+ASXgT34LGrw/
MdFecncB2Mj60wvG6P6N/VvGcD6aMikK8JWCjb9ubnF7k60I3nYea8+txkJ+
0dlMuMM1JpoTWZmm9Z1YiY64ZeAyH8abrtackQ88zh7nipxGm7oASLEEGGPp
zQBKvwrQDsOhwlIVq9bT75HqsKr8AoiHBu0o2cVRiY00cA5VIX956Sn9+46m
6t9n6f7pPFoBeckto1dj35nvRxSlpSMaDiZi6PYNQRQ+AerKRPvoHkDDiZsz
WcGzGqWZN7ao5ccY1xebJvCEF/DLrlSSEBbLOot+Pyp9nYfcm6ZYTVOKHGMv
sBtQg9jwihr8c2SCnZZZAUft9ub7mr08Zfgjp6Ptb5t9pE65JP5+iWbhahRN
bcxUPMr5X7UvKxhJgirkkjY9m9Z6LZKP/DFC9gwY/5T4Mr2vGYqmExrvLgO1
gnO6K+b4JG9YOCc1cl5+wjGPbguxEmTiGnOy/ISJYhhB6U9wKZ46Wr5pPHn4
vOTg7qmXUMDUeywDSaOUt537D0guQEz90xcUWcEUUm2AeIK+AX9Efz2rcawm
aaN0zM4SCgGJb4QJ7OvyutJfP9gsxY0iu+7pxQhH4m4mT3xkpJhj+U3eRo3m
rLvKjVCEftxTOoEJclw4dKfsQYNmlmXXic2psWpETjshiJxYyszQIy2AzNeG
2Ri7Yfn/m2xahdhFrANBsftgiIW44k80lTQ7lakNolDe2afh7jW5tG9J4XD9
PSqevphAf3OygBA5aY+lkADLReYWjcVTRSC2BOfYPwkTnvM5bprxifUhHhTq
DP3Beehf1AIprYEbghw++DjPl1uUVz9Ezhv5l034DeNyQli6tdY9uACfIeJv
a5RYHvc88BF4JuRyMEi50tV4vXlgwFlnk4Emtvbw4/+qwFyW0Ev8fgBxbkJq
L4nyDojWVCU4AU6UL8Y3TWRV3+b/Y9inmLwJWkiHxMlWPaRQo+rmxRFCvnW0
LzSr8/4pZw4UalwkrHF6g/z9sCFqRDo8D3zEBS9B03TWkl7FmGVQIXVWcPL8
B2ej7blfxG32+gNEn9LYBXiYgyDVdy9iXQ1hxWGw3gZyljZfJToqLwTslAcJ
bNiJPXGj0+5F56zSOFK/NzKxiBW7PKcX8ivbrwS/9o6ubULysRZAn0+CsiTX
QDqYaj85mrC0ipftVuNk80U7iTZ6lnb3M4YmZ6lJnZxBtF8g3G0Ix/G5spzD
wFF9ZIHof6UbeE9tvQabYOczT7aTeA5RqW9vj/VFx219FW/MeAUpt8iACNMy
g8+czUWEmIqw+6N5s9HsfHyx47glzu8YvPxXkYjQjuamjknb+d9RKLdWxwjc
jVaSMpmQrsZyaYSq3C9ALbMYU0s2+MeJVP0eTmZNpKyvOA8Rj38Ox5RusL/2
osaEFMBmkPRlAKFA8YyWBILK/f/TDGSoUtOLGhsRC1dkINlxdhsvTDvMm7MC
jJJGZNJzHvZ9dm4pnHntH9XTTeLqH67Ri8kGOMCFFbybkSOC715hCCooJGxu
2/AWOI3/Y0qTTlsdYfa5vND+gYkNDQ3sgEBE3FE2HzTadntR2nIdkWe9vVzw
lFFHlVfY6e7uwGoTfl5pb5UCVZ6U8LG8vYca/dBvaIqCnUc6Ont9u4sW1R6D
dnJ7xQXE1QzCFW/sC+aqp54mzzlDfdrYY8P6jgJ8kFpPrp4RumvxvBtotF+l
ygxKJO8M8laUkemAHXMTrvt216gd+IoXTOIJ1LTlo9I1a/QfM/k2vvZunfDX
P+WFeHJjJsKg0aWuRfzks0Ig8vU7D9ctXGxxXPRNiDFJqdwpQNod/6LcDHQr
T6ZyJACh69RtAeCPddx9TyV5OgVmyiAkqHpN+MuZtrKuZyEgxCfA2w+tyXfh
Xe5WCGsEzqiOPdggURnmKxcxfyTuoQaCKEIYVWwOBRAy87y362UzD6iFjwXa
PF8r//mRbXT4JUyz5YInwEjRycyxaqxvhWORABzFilQ3ulvLL4eix+f8Vacf
9a9X0cnmZ3PKYlufbZ5sGxilaBOj3Eun/hfK3qeylc3tmXywpV8o5+LN/sjQ
KkdRBLVLUYSc4zmmPvEXRAXT33CZ/IZ+XlFxUDHq+76aJNxlB7+YEOZHVHZt
edR1eiZc9jldTH7yPl0NwHzjM/SzkGTWHx+uRH59sTkWsHf5r2CddZJAlWdz
BYSXbJosppYFS17GnqIYE1mMKUG8f+WTu6rFPItUW8RFHMO0sXH1neaOdOq2
Uf2QGEecCNOAlI7TroOOX4Fcq+Qu5w9I/aPO4XcWMfqPoTwVZNMqzvQxl4SC
RNVntX2PvIEWFTGDhogYJqa7N4QAW44wq4vHsAYWRU2LEuN46BWaA8MJPMfy
4I+V3OfjXbbJ+GX8fRCCvVYFV5Lfc8+33De2VuvkWiik8M0rs2DLaJOZFVbp
pGFS+KCXlW1eC4E+nPvQfhAdthSRYW/G3c7MxPNEddQzmGlfYjT43uQ8psgk
TRtwGMBJmUKjvRXcrUvLZa0r+Ora7pwJ03Rox8SCEVW9P/q4Tqnh81DusQsF
+1UzAXrs370nkjoTEZUsHXLBkrPZFOg2iyYUvhZaSbF/9ZJw6uaobqwp1Org
LjkkiCzULca41Ht4/+JsxMS+HbJYpg2MRGu++clzGe+nuvjjFy13qWDR1hXY
vUlQHBg8qJdlmKHE0q1xXaPkA25wVMVfxD3ewzmChWsQK3Qo7Ps92aJbhtjg
bMhVsdMo11kFYH2AYkQi26NG79iJVAPg3Z6rDFXCAdWdPuTcEtkEt5GBApSn
atf+zySYGnaSHTJq9R4rhRmK7I82U7K5xj0r1S32d+LIhti/Qnyoyfo3jLic
1olBfode/wkTOohSdukFh5PcNizLGGqLkfiOfn2KDqLKirbfEGNIXYHottT7
KPKVOf366VcJkC+32/9qN7RkSllDw75ku8gIqhZQMiCOcXQuwH1z1WJRDYty
S2mVBgorEaoM7yK1G+L09/JNDaqellMoDRmxxi9aGNfcPBtA1+FhwASpkcLw
6G+8Inv7fhLxMtc0qbSIjdKRF10+WmbsBiuJH3mSIN8cKB4C5F3NWNQ7PMb6
Q0AZEewPq3jevyb2NeYYyaXdgr+KXhen8GZ6Cfvi/3BsGviPcuImbKOYmwXY
ozSI74vDSEHbM3O3eEN2UlVfUjhVVJ7AemEErInVclr+v+je8aMa+37yv6TU
XS7R4qMT9jUlGapJMuv+XHmOgQvs7erWRmd2HFhRo+oiiNPcEGKDeqpGA3+u
0Nr8p402JFM7N+8U4XWs9d2vD6eYB3ISM3flWVzXaUsZETWHtludoVke1sZf
Uuj3JLNfh78RUxL0IL+0Jud2AoDa3b71e+wFB6C/dEKhQNEOJVM1n/93QHWg
Lwz5f7YRcj+fQVzyg1Oj6T4NVAcU1qvDYwhDK0TWyk74aAwqE2KcRPlc0FLI
kldxEqWbptkkgoS5PDnNG/twFzkNcju3K3MgQGucB+KcYwkEa3tet6+dLIzn
+Rpxlo52dJSpilfqloLBpTxB2c3Mz+PW/hhA25R2o/77YYpcFwGiEwwq/CUi
dS1Q643+KhG6GGPvV5qSnfoVbIpas7aNTH3+Fla+ao4yD+8WZp6eqEpB9Czx
iv75ZRwBAb3/XikwrK9lR2/azd3mNMzd9b0qMGmk04YzDn01YLTVX3G2Mjt6
meKLLOXlSIEGmy56OvApJ8sfx25tKkK7iMRIPw/CZg74XdNUlgTZiEOAArSO
BE37N8IqvIGJLUvigY5nTu2tnp/qZJQsiwlimzQnkyu+LxNHI3A7191JgaG+
pi3k8C+ssvOni9YNW4pM73o7a3D608jkRFlAXsnbzkbFMsdiVps+ENMtXIrB
DKeY1he+uwRHp6+LEL6GR1JEncQmAZUlyPvn/m1UcH6XHzHMyWdHecFQ5KUZ
duopuNxpPs1E1MT2eIZrF2AZj5aL4JIx8Z8VhqCP4koe+T1Sh9SToXE9IoBO
Yh0cb0PImm3o7bRQ/IwlKlQNE+npyMFFpszEbM6sSoXg2n3+m3tgYAcBT1jF
mzuJOtYqf23MeSS3JIzaCAyzxKgP14Y93jsOGCFB8+g6Fdi+o2ONILxBjWwj
5mERDOg9zXdD6S6PeINya14J1H60gWa5mwQVJYPQv+ZNzJ/ru4s2IvOW3j7g
7VzB/2I/yCRXKg2wkVNSeh4W6wt/kfTkzwJGgTepYnEnmysdTpgX8VRQ83mw
gyqAwdtrZttDo8rqCX0FYRzUm1zsXZY/k93hB1OS2B/D/3ndKulAUSphMF31
z1gYSKdrFI3JRoXUahLOE9glIXYtiYKn5s3MKGIBp65M+nqIZxhSykG2zI+O
zujuqG4F/nn3sr8z1G+rSH/a3znzarxivXSpx1KMfUm0I0XkEYg5PWtHH9Ts
27VsdrfaMgjelna361aK/gsRQ5D6YVzIoA1U9wLqjhBiA6QQKYKNYYo1Kk2u
5s2j1LEUF9QZlVCaBpWODVdIz7u+Fi6EpXgl1tgEHZM9Wte0cYlfD+zFgU8v
LzWAt3TtPWA3OzH2TGtIecAy6cPqwyX2uUv6glMQ/sS+TjYtkejqfh5ny1Tm
/cJk/x0Z4bqjBvfrcwXxnDfMH9TMehbNTEejYw09TGuLo7VuCcOFZG/MdpT5
huMwihbeI9xFex/RV+8SLUML9b3ghM+RsASJiypPXzHdLCZwzVhAsjclEnJM
efFlJqFwdxuVChMRfO5mvuwCpuLSRY8lMTJWIO6GVjSzj0QbWQFRkHo5SYfy
NTVHzaG/3un15PuyLtM3v5tfmZ5boh1YaouyR4JvtpVnDXSqkO9HzQYkxXC7
dHLoZSOKuX07bWb6BvfAp0G5BJtpB0dCLwoe5yrv3rHQ+LADypbZhrDoPaQQ
34pEaf6NEyFtkpGMDw/BPb5z48/8jcXIPjhxEo5Pc65j8JRSdZWWbJQIuXxD
bvYhGMwL/2vdDOsGqJ7tzsP6IwlJQSpn6Th/FL3DIqvWnlLBMg9PkH3okyMA
Q0yQ7nOLprPajN0eAGtPvKn30mymUnC2cS32hIcLhnu0w8dR2+4+zoHc6e3y
EFZ7jMJAeV1flWtUHN2aVjhH9QS9XtkuWiT4zNJDDHBeDfV+zBpIb7kpx2Sq
dRZY/pQ1oAk+tXwY/pVhB4XJ7Tk07b3DzKpbMYrz1UlOw9/O7caqUvgjJx8T
IluzWJJHuBO2Jf4E1gKZBCZnM3KjU8daJDUoNAuYgsB+BDq58+c4giTwfTCo
9mcUhp/BRRJ5YKmczPUhpb6IIfjN7XYyN4dV31k0aqlwJXk34BnPO9dQNvqr
9vxaOMkNAGZ2D/L/yHIgeqqNkZX/+uwNh+oS5N10uhRJLsKbftg1OkjOFWVW
PR8L9A0/hLpU0C7DLZg7xAOfXQDsEOJIdEQFDLFceGL2Y2WoMI+ZvAX6QGfO
t4M21Z28WDOz5oLM1VwGY6eDUEhuL/3UcEiYGA864Q564dcGRxJclS32xCDU
FyQL/dNZ8t7mKtcCOdyXgS24Cjajg88kFXJKJx3lttU9AUC8lRVXS0mbORcw
mMp2qE6KucoWtLjk6lp+ULxPQrfwdE0jkmSe5dM9i1hHDJNAIWaMismB6mD4
WQewvNcIOkPVMGCz56mKPdvqE7jKvWapmxbUG7h4uiLU8z4wqexWOkI0TS26
RLqskIj8+lbR8DACemSKf+sMNb1tu3+el5JzPhE/HrQ9s0VbOC67/T5TC5IR
OCgLP6DrOoKimIomDUaObxoWms2F2J5jbnqvrYacLTjrbKleknhtCA4duJLp
TCutKfWfACrjtBfPhsVQKwunSl3mQxL8hwgPsQsSU1sC8M/ycztsFYHQHJ12
lZQPrHaKvraV/T3/uHitPz6VJGFuALbz7m9dtiJYT3x+oFNCeGh94z5dkzTF
IaQ6xY60P93CJfhbf1pKTi974TN1mAkCs/iit6AnEapDyUm+MndlBaYm4oSj
6cyRsAO1YWOn/PLRml5BFs/VaLMlThKEe6MX5Lt0W1gt1nGwVKCWN+QZAcUh
IivB+JVxaTvQj0Bydlg1FAWBpUVW0KdA1oJ1Xs3LEvFMD6xGxTNJuK/BkT+O
2CvVEOZ7fZl5qSxFQT0Kxdn+7SqnyE3Bg9LuQpGaDWurvCgZOeykvdrTkOGz
y6cQc+/QkwEejOuqMFymHoCQuvIz6FlqsD3g/LH7IUcM/EvZo4XqdBvzggHE
OuqO/u6WjgzTb5thGLJMI5qEd4dqtNuF22iVF6WnTzGI4oz9g9gteX6LI9OD
B3JSL4HwZWxWjgK4wy8DGZ5McMP7A/Qk72SomHTb6g6CWroXB583tgEpDTVl
XGlJBIuP9piup/6YQyq8S2nOMcqBfNXdHzlg/Avk2e9u0fi16BPcCLamzL+y
gBZxKxEPoR+v5PVOr1MuuFeWmeIuPcteckO8cTKOD8sbSxYeRZQkybCD322p
SULWAaEkUKDHa5VXFzxarvr5YzyILs+hlD5Gv9c+MKXuM0/sVsykdUgUn4BS
nnfPMyRHLIv0HR7ZKdYuYcMCARaV9GdCt+RF3c26tPe9IJ20bBbnDuah8+QX
UeDcdq0cmRKxZfUd6Iaaes68driH31uq5Y2jrwPHQ5eIqMpeBwNft4KDaMdd
VJyj10fP74XAcRX/tWTRzMqctZ1W6wVGTfQ4eSV+NWIBv9BUISDdJQ3lLIBC
kkDCsWqCi0YPrqAzLQpKkO1H/gjgK9QRJnML7xXd/dOkHbjtQRnVRJU2V+A0
HJyyD4fQgfDr0jhNf0zUZxqqkjTKP4AQ1anOSEahNp0Hk37SPOGP+g7hGfXB
OgIAZQkkKieZ2uojfbrtcH4gVbpXcRz9EZHXFPlrKmp/ywltmm6KjmBykMwp
DVQ5vncru4QDsqy2yejETNyIXili93haNO4TV7Tt4c1FSU8004HvnwOhBHal
OiD7zgDp3umvXPObnSinylR8NYoMhe07EzLP+G9kleir6Q8L4TowBwBkp3M4
B7nqeomCpeQoyHrK1Ky4JV6z8Dd2NL63N8e2hRC6zEoPzypVoDNxQDHFi85o
AwIp1muF6+v0Lx31UXqpR72uCbAs99TTNf9R3nZ8p5HxXnith5oGh2w5HN0y
WQmvDr3bp/OiOmwsdBhO/ndntrJeeV1ts/ir9f4bRMEzNeqNHgHN8GGfEe42
55FTYwoxNyfS0RZnNyEq/4HRG0SqxFwsR0Uj+xhGElodb/ze0Ala3o4A+sDH
+pyJwZ1bAkpLC1Kxc1zPHTRztqwPFhQ4Xq674O/n9f94y98awnBb4ws5lo+g
Fb0oARAby7liyUIkiR6ZTmmzrbwKp6q/5lnR2F00CcZSoMfcYr/Ml+mfHcqN
ZjTyA/rXCQaEQwbjvB1Lz7lL/cxGMo10fgE+3ebf82pByEmgXcQycLPg2Fyn
F11JHDRAABfnSJPfr7VqHVS7ZmLKYgrHxeb9YsPWsEYXBQA5ZM0QQSavuc3T
YunT0P5nP/Z0GZYgvFQJVJxZ7vk5nV3QCm1aa/YyNQ9XEbWvjveL7OrZcRr1
jy2h/Co0IH4ljRsZLne+0GMK1qT39fidFgnus2MmDe7ZWITKhx70+9sCLss8
eMSHhQgozwidaPNwGnab6hLU764SPCcxSaTiuZjIDxFY5qgUN3onSgL1w5MD
nWf42IVF2s7tbLVlJwLSXGWb7YeO9Qb3PPU2nbEIyvhbftoyZ0TWf1bwHNgm
U8bilkyPBJA1ZQNVYCDzAeLyWnswerMgPY0bAkmYPhH5he9v3h3a9/NF7FU5
05M5tqusMEJADJRw2a6xNKfWsDP0edkXGzeJyeS8JPeIn/sq/8Yezn6Oa8tD
k5WZ9S2vfFesvncNHUbwEt/XGMzJZABhxyZe9VHH1BlFj+4+LLKLCcERHige
K2plkrPG3e5qGDR2fW6j53eo3rttemZm7W68yWX9mfFsjMLVegAHovChMlVR
ViQpv+ylskye9ihHdXWpRAOL/yB9iYu3AXY8HeeKCojQB02igqOwTtuhNBWJ
ShhT5FOyDFAApVU18Al0dFRQheuNKwWzOg3mtKFWhWjpG8KTW8tuID4nNouT
eGbwjvyiFYLbYl6iMcvRnpKBxxS0oPNGmOU9vmeF/fUn2TF6Q6EFxwbqeUcj
X8TKFDkV622a/SgdUNmZ4/Y2M2pkZC11pMnQzShZU3hSXBqJBKerPKIevhGw
YFEvmV+NN2rIaViFjPi46bIQGQCXOEKK9fQS8tsHGgCly6dLeShnXixCnK0P
+Y9PWEMYjYCBz0k03cyiKjT3J2SjozPA94IFKTy/kbjypDkO4AtIKmEmE0KL
48w9OC0OO9sPProbxWebmmjktH5h+Dj0aQZ7TkszSWgNAqu6WhEfTuwBK4vO
SOOqOjMdBCyniiMFxGcR9TZ5T5H8NtdWXaPXL/TaCfjrJLhTctZxPHk6l2ud
ljQpQU9xfhimeumXB9QZCtrjmHP4FGv910ps4sHiQO/zndXscaSNUXmyWl0e
wEBXuBQIaqKE3S6bvjdRudru+JziS9mIGKG68NmiqjI5y1XUQKSWtcIj2zmn
SBNA1P2p4z3BXevv9QnD9hvEXvyBT2GqT/LzNZgRsMW+IDann8A8sGno+sSp
2AGQMpcGTnLQIQtTL+NAy9yfpz4x9na9kYLsik+n5I5ZkUWzRCaUhmXtKlJW
EUqeJj2+2ftDQhJ5ze2/BmkmXX2ibRPlHrflvgcJJaQvkvU4Yz4e7eu+wr2B
C6ZN9EXIf/BmZx7XBpP1cdzfl173Ict7e4C3+sdFjZQ8XO0rmaw+ivorD8ln
S52V4J1ToX/wTrPVeYhcf5I1CgQ6CGFCd4sV0MwGDBonFOvjDeui+iLzjm1A
qn7Kt1mCgy7g8OhWiOsADOvKzeYsXGjWCIDP24Y2PI1z+ODZSsqe4IZH4y+d
dP5DjgmCF4VrfrpcuLD9ht5MaHpQS6w0+BhFyXB8LVpCAvZih3Zt+zHe4pO7
1mhtn9NcDxniJfGQPK4JfJSZObqy3lU3dOIOmH0FOOAU3iv5FHddMswkgyA4
nIvoErYo6jdvcxVXkAsNQ3UFBvjv2vl3MyC0NztcyqHyyRrGkDE2RjUpbGWq
8IILfJLOC/ReW8Mu/AvBZLpDrJIRvQLAkjVhYGTQK1cPDygsF8afS99Xc7Eq
54HkfTyfnUD4k9h9awFN3EcwbKMYZbUb4ossKy/rLq+dkySjtvAFb4BoxBj/
/FZhw7acO0jbjnXitTgxG3O5fZs4yXICVM/IwPAq/rfgCaXun8JFJihqL7nV
kE6rRuczWrMQ0t9e2SJ0DSkRN4mb0/PkYsnuZrrKuutfD3tth6BT/2l8rfe2
LfRHs/91tmtpcenTv5hUHgK/UFNSFTCSX0aSLC6dO3fKTy9roPtI2v4eaNMX
1jeL9eNQjxEvmQXN3mpJIJfFFXAE6ENmxqsYYC1Eqe0tzTrcza3qAcp+O1PE
tkTXOWfUigZdTM4Rg3xiwoX17QUhwt6yAx1LzfkP7fxQHKr2c03YbJ7z6LwP
jnCYvT2ifp7asQnQCUZdbhkrMm1fnBEXmSFJzB3Swqz9CFi7eLZqiQ2kllnp
miZsHvNTeslTSIIVx5oXjqy+uFMlniW1aNwfLvOW/fAaN76qplYPQCnWSWqc
CEFcGuWOtsgH1vgm9jm/2YTFbcn7ntTLMK1sQ4pxIf3MVe9xfBXo6SHoAcVt
T/KO/JdNu2AAlCkGHrL+eVGRPR6FCJqo6iZiQAzgRvTqeO/4wth1heQ4WbOp
l6qnmNtAK34vsfPNSGAC/HZFxRjM+VAN3Jev9Xr5On+UWJTNMaqKsmabAQf6
yhXmLvdNkvCJDLjk3BRZFanlWE9UyFHBCbqd+rNoxCw7iiSMW9mUeGY1Lx4C
owwyLqhoMOMc6+NSMld7h0PKfsE5JX04KJ3/JXpZ1RGpju0wSnwDOs4D13tF
IRrRJLW6L3LfGh3nKup+Hk2I+s8Z0WqpihDLDlNUVe4+welUcGMVAtwGenKA
Hwx4GPzZtuNp9AC1tBHY4ZtOKXQVRIaMWicz/K+Nd+MUbcD7JvvoGuQo6xqx
zfYdzDrao967320A8atobcVTZjLkbXq9lPKFx+ATW/olqbQxeCzYRmXYSIHm
mwHaU+U3g8YWXZdG/JZvorxsVE61HO2kWVf+FRGnMBvtEyO3F5cdN4xNPIBW
TRLKKT6MBPMAdDuHGz8jnwVhTYPUhYtRKCzdqgIRfCacwbLRfOf4H9tXn8rG
a0HB1XN8BcSDU+Kp8JRptojFFhh9r+CfDeUAFICU4Ra0wMiKsVwbV2VJUUa2
Vna08DwJtoSwSzcB0t9JNR4NsbWlvd64fCtmz9SWH7ThqdPKcpzBzNC/YIWQ
6r15p1vDFgvb8LdWNTdB2g+TxFTR6ubU+t4sjqm+wNfCwvOb3qIVT2wyB2hu
FJJhT9IThCjrlesewg+OoegXZiyRJb/Qvki6G0ZCDJyK7lxRwc3pAZRI6qC3
IHiQU0qsg8A344ZpCqu65jyxURJ5VM1/KOyhK2lb7SjC+ENdoii2zvUlaz5e
FSvHK2IifDppF4evKghsCLoDc4xI/fPfSk4Qh9kEML7eiNIfqdCSymWy4gI6
CHJy43TUZBgS1QRCTEhM37o1AjiyI2MEywEeVYgEjWMvJZnyLDmnDdy/gGS5
HL+K8u/EiTJoi/LebVpUEeweEfZkxjSYaanPLHJvyEFs5ed57qDDpVLZy/TJ
WCToqXvDMm8lL68rTR/yr8s3qEpcLryWivCauoi3V0P9SGFZb/TBOjWky3/W
SF2HHUrZVhAoq1ak4Fu+wVYUO2J/AXUv6QSipHZwd+0VDeobX8/zTeInbsS3
vgNiahbxpACjrZaoYxfvcQiAOmD/gAO10iB8CChs7Mj9V+cKgYBISTRuvnVS
vAUXAeHGeHu/3JDtWS9vonnp2oJHvhW4X+XoRejeWMltI2+TveS71JBS67Mj
iNU/OfIkpJbhLvidurU+k2C1NOZVNfBCzTnHY+FCNM8A/ZBTYWtWUrmkJs9w
RwJ82oYfKtirb/rrOKyppiB2oPduvxtSIQQRC+OaGUrbdwDQFkszGu3Fa38V
ImmQOEGSeBqRm4rZCs78uUIi8pKJ96XW27NOicv7TkalVDdOzbfS8jCx7ED7
IcIkYsyocqIpIHkgRTa7ilEbaV8kRhYWqKZqJMa48Vs0A7wWSPFoR8bDN3bX
gujfpYMhQQFUi5vuqTPrmI2zjKB74tB94TcV2P3D6Cjgt/a+0Fz/Htz7GQj2
3cmrJdps3OznfDcziY2bzjXD02itMmNGUyRWR9W9V2Evzfuc5oXx9c57yZq+
id9w76TlDH/8A7po0dw5NEpuBZgwULf+Sbce5mc9JQAowqB5N0NOUez4dvWT
O0FNVylbM3RvHkhXjOfE8JSpGm/bxvYYBoP2MlZiVXJ5/ztc3hkFgPTlRYsG
yOgCpVnvRvDOEY8nXKFgOEnu1Q1boyNa5kyN7cPIzqCGAJOn0I8A9Z6mZBum
w5FL97f2a3RIxcpSKKB3CYR3faGVea5AYrU+ClLyyUcgNN22kAWdxSehQar1
q1KgQbU5Xt0Kbsh/MfrayERVRmuTqsyhc0fkTgSVF/PxVBcLbgfDh+ddICE5
lareXiYH5VVPipkQ6AQ3UTXa/Mo1kyZ/rErp3YG2GFcllN17nTJUXFLl676F
G/ozmH9XLCJx1dS6PzqOkIemMFTM7ViopFaMl3w2qgxQpywRrhFHRt+MB9Oi
Jz/huRprxBljdcLLD+JZa2Lg6JIBW5ooYuDb8hBEi3vhm6ZCiWx8M8H7s4uU
UgRR9O/3iX1uuv4AreL4q9HXyAuNFpk6iO0O8Wv/xYXQKis//QpJhZOMgcZ0
CHJoRwcIZW5QO4q01D72qeyqecWJTlSGLQqJFLUNMzdh7O5hSgytlY2jzibQ
+kbkoIqR4tHu0Sj15tKHentuK+k+GK0/hEC47WeQ+QvknxgV/5yckAswtfOz
M2igsngObfVAbDjZuHVQgvyzFNDbpsft3PIG4doo/g+DOMIf403Cnd2V29dH
JC/BvGgr/AKHoYaMOQ7SmDAq+ZFGm8lA1/VdJnoJjVXobIvlAk99IZKHnfkE
eBEPLsf+259oVP+PlYnnOI6y5ppFK6YcFYwzJVRr9SOqP2xUcD7hoZdIcTgb
YXWllyC+wTo2ge/gObHtIYToYt0rlc6ddsQIlck2KLpVeOjT063gT2lPJIrH
hsyCKhD+A8/YtWoxJgYT9WbV3Nif16UtNaYiiLyqsWNyq5O2v8vG2KdOKdmU
p7OCBzPPZ2hSP4bzIU52dRJzzMnex1msrD1u3Jka5zMykF4t/hNXTH5q8eZ5
bTby0kNsitBMDTe1dNcUbhRLBwbCKmWAHCvWhVMvrhctRxkYq87HMFSRyxvu
A1VQh/0u6GOyHCxS1qu9cLiOTL4K4orGAaBWkYqE65vs6vjpxouMnlUMYjIi
WEtWKWLAtN2HrbfFxZkIIMEkblmHTelQqTwVKB8ncrvie7/e3+3cRM/hzSmI
8rPtgm2ISmM/FcHmWYkM3A1WGAyNXkJfXahyy3Z2TkBUj3AxkFlF+z0eHPBT
fbAtE8lJ6pnzqZEOuYx85cYL0EUPfxUGVwm7NntT7qj40FXW0VZ8our9t0aX
VzwFQbcO4A6TCIi/jKVA9lkhT1QrkwFsZFgFcf1M2ZrHGpsRw+9psXLOvJvS
WgYiGJbxKT0TWOtv4SviglfhTC8jCVHllogIGOZcTMk7uc3IGreS0U9k1qHy
+JRmO6BNt93bv46kcHkAjFNGiYH48kLzhYIQMYa2H3gKQqVVfY0Y9ZBtMf6o
ENupQOlI3XLC1F0HWsPadNPWdYmHgWnmfLpn5CbSdU/ry3H+Omp/hhlIE+4W
9jIgGdogChEURb8J1ft8eApUWFB1wFYvCxHHx5Xe51SOxxuvACM3D5FSccWt
PVKhPbWXuW0GEEMAYSG5OZkFy+/pkVp3q1/mQEHJNijcYhKXlBD/JIEhWtkW
NDeurVY3pkyuDypkfjc68juCA6i8iCK6pr+5hjbL29Q8zSfIZxWpOoTzQMmU
0z1jZghn9YAjHLOIS/TRbVszNLvrcfungZQ0bcCGxciQxr6C3mb2PUmfx1l8
Lsopfjq5kDJf7ax/6LxGxOzG/O58VVoDKswWSxpGbVP7C0W3Rv5cbX8Xrhxm
efp6HDINEdqEGmaSh5lAaZvJoomIGq5iJy0W/+7rFps3bjwBg+/IeW0mlQcy
84gL16cI6vJWs42GWKLO1/QfC0735ENBZgWTaV2NylHummMv4Yn5F0CApVRO
T83e5uBAcJ6LZkqWYM6FW0rkQ+2azVp5UeN7Z4ajSgTuWD8x9Z/IK1/1BOh/
xjpUJPBy++U9DyRb3a0u1Y5DYuql9HQbC90L8hTNV+lxAnmoJL5j+bH087k6
/frqPpMKER3kp490gqH6g1OcygNYp76c0Vd9Jx6VUWJxDqzZPqE647pnK6XP
mmsqncgJ4yboY8f2pWK0arQH+aHQaCVkveyxudbxcsREPB3QApgIhAHXID0X
P+AGPbJOpUprdEkBS2a+Nm825ZIvuRRCAEJwXwTFzmq5TRDA0xIW6Utc4HNw
+oiKa6syI4e+pn4QCGC83YN2hzr5vDlRWTZorIL7gaVjrQ4HRJerT0JY6Snh
1tCqJfP5oE+Q4fd0mOE10MNxGj3PI6dcj0Qmu0OMXec+cOtuCtCPuP2Ixofj
DtdjJ11EEP6NXIB/tT3Kv2ofmESqpMW2XYropKX8spstCHFabnMoxRgYDu9C
4IRl6pdhMvBdp0LzHjUaq8kMIRn+QP9QaZ4ILsyuLCuXbuSQeCTDPuA/AGw5
aSOlX757QVvjY+qAUntZ7J2ybtu29zjqIqN67tuU8HiinaU8jpIIGskovL3i
uvh9+4MpJEVCwA9FNE9213FaRi2bCgGURWdUiSuSa5MNN+Pw31BDF99NB7cZ
pKT7QV0P8HdEzGfpsLLkZRDgne1IGItVJ79COZ78TP1aHZG8/Jj04eUSbShY
AXj8RUIXimqRmMU3VP4ZTUO48zZG9CyF1TQBJg9r9YdxD+KYzbjCOOOik0+G
6ASFg7WdjJ3KWHL4rnFWG3E1QeVqmdMfnJLPm2zEDWLszKmUUqz9cMGumxVb
DNLEg3t/Qir9/7a8IAiEDHYkp+qPdRsJlnXdrqV2t2g4tHI0DlDutodml4Rp
Lf1Y6xv3c6zAOn7azR2QDHtebMgQmh2yjNFNsJrx6u/qYtwKJCqw23Yd3//N
4aFq35I8RfSgNJ+vNdRreviMFD9du9to6jr/ma6kKEu9xgYNoh9e8/+OcfwT
PCkt/2ZT0gRtGptUjFAxNT8m8Sv26r580bfkVRgSjRdxub5Tt3/b7PFfgIQX
92Q1yxmKQL6VhSiGF9i7CiZ+ulgYVapYZ7iCAzZZYN/0pmNnG3AEom2D8iWS
oAdwntLspbH2K78VC/E31XZ/U2iikYUIQe66WYYvu70K3nQzlcF81okiHJMs
ANc+G1nS1GG7Xu6QeSvqTbt8f9rbgX/70UpFdqkzxbKZraqmKTvQQccfR6fh
dJuC5a401GBGYFk4zRstMkLLO0AlYbmSbe5uf6RJZV19yhxsZUaw8uSLkcIq
KcGWqNk9jxaGXoHKv4Jzhlokt5+gdbP2nIDObOkYPCmonlucTE76sdDoo/Up
BoRjwns6N/l6v6HK4tK1zm1U2xGpUy1iI376BDIJEcWsXIK184t8cc4EwMoe
lv12XyrtURaKOxH7ZBpokQdTFFsQ3uMOemCkWPSANjoCcjqMNFILH6M3ec6a
cRLI9anoveQtTLAqEeR8GSAoYLYDTHf+q2/VKQvyikQZ/xQ4M4ZA7oQvyy//
zWDp/E9ENH8tcXi3bo/i0CKy5himuaqAml8XU8RuIBpJdu8FS6hLkW9vipdS
wLMgIPXFpwl8wI7b/C26dDvzfqhFSEmDeOppb0LLJWnNX4PwM9YNvsxF2gh+
em9mdUdQvAHj1kH3RLGcrOwEXhJGiGMS7U4EVaPHgvVQvng6HDJcLVd3Z66a
9w0de0muESsT1/Z51SQDjd9gLCxMjt5oYeFoLQj17tshd9es9NQowKCZWSV+
w9so34b3iS1FgpHCseecrHbTMyFERH5AyjnHUeRdzrWhuSTeFamKh2vS8s+j
X/kpInT7/URohzCbRE1k1gZ4IOoY0k2giCAtBbjvw0XSZkVcCdYmOzmDu/g5
j2kkqOLv6WFQSIiSK3TsTHQF6g07iDo7sSfdshEashPQHMAYqa+xeUWV5QQj
N9kol63LJnwSbSIKmwI1YsmbBf8StYA0qgHNV+onUFKXgf6vldaEv8hLe4YN
ydcSG7RNjeHU9DcbOO0eTQ8eDl60/NJbA92YPimjfZDqgDJD7UEOWS8hUi9L
VBAhEnydpgrAEl4XWjw4fWZfPMwtIbXt8fd4g3m3eOgKdIhooR8EXoVPm3sN
uSCtLm6GcEyhRef1U0siKwGMJnuY8ATSzAY87WS1MUR/vGNN1z1QJaJhtRYo
L/421wL0UzcJBDa5jRK+ymUvklHQK6QUWoGsZGOIPDJzjlqKpl4a8jkYBLYK
B4pJpRz0RfK4aQ6KrWc45DzoSpS7V57bJR5ZQK9bKAuRjz5Edlis55oURJUX
LDbu6ZhLDC/sSE63agPCxcGOLbQA2ebRhA6SyNrx4WHesNSjq8AQyvPP6dky
1R3GcS1O+VKL7THLOwPKPe2w3Sqpu3zT0gV3xJvLfpE/3ruqIc8wMGOVb2Kt
w+XPtvPp3kkM4fsCUzXTfxpI1cNTbDbmA2UmXWdvd6IlPUuCZSgYwhPnhDOk
ScVNOEB+8QAkP0kNLq+X/yOyfKz10kblDzTYIRwyqFNkZFbpOx/eqr8lClkD
rJ6wyOTRu9d6GxMcxHHtbiW9xQq80q5CchMS0czr28YBByte3wfrMvDXUWMQ
Oo1tkjCX4r+wEkiyAF5TXn6TxB/xXr2UgG9cfcgcI5IGA3nf9aNQXqmfNV0d
zUH29/mEHfNLH5Hz3b7B8JUsbLlhdWySNVRFCMZWOIE3bVhmD9dLkuVpX/S4
KEcQtHmeK3USisBOeycN2ev1arK/u+mAoRmLqtw1OJz/WiAxPKVF65Isc1RQ
zoa0Bvm51Bf194CrWD9RB4kLtHPVlZAynOjS9rFO4ky/JRou1E4N5a0LpHjp
HlLB67y1BsUnOvppIMf4EYbJstZm/vReEhfO2LGkpzh0zmiOe6TLrADt6Lpf
HG0lm4l18MgCxSn7HTrivLwecav/lddkmaKZ8msghE98YjdJLX4lbE5HgwQv
gilDZDQSzejAzRQ8rjY9oj1tb6KmLUtjIvenlQmJccMwgooviCJBGf8J+0Uk
xCTvdEyR/HKbLAckXAikrJIdbZ5TM0T4IxRhidlnVTl8b7wRhCDolxA1h1g9
muFnUUMCvcFpQUi0Q6u+KaQaW/xA7Dxu0NAXbll4S/+urak25PTeRBnd3o2c
a9VRlKSsRIP8bxA3AOS9xrJQobZgCphjh0CGDIJuelyzQ7utZAqwRcGQRGCU
ZzvrOepsczlnk7DLteERaAKStbZcdms9zuK3fIW4/zfXmKuUHzdLazyve/9v
i3mxsFYKVz8mD94tlRBrRAvXaBvBbWtISeGEyiwavld1Im/ztRk4y0Ua0IFS
wuEpuqv7f4ZCJNYWBOZ6hxnyZmn4yJMejxDsEF3wKUPKzrBXf10WHG0z4vUj
wfg/U10Z8HA/kw2LerhNEh5KwB8GKQbAL/1bGzF501CEpZ0QF3Uu92UYwV4i
4W8L22V/Jm2Y9GFw01H+Z7IjcXuTWKPlcWBOTXuOvGMY4B3O1RUxNfiSp95N
iUfV2he67DiyGoLYoiJucIJ61jfPLFtVvxhy7Qj49R/t9N0MBzwtiFEMlqbB
HOCMQuN0lbX015ALdJY9hahuBKKXnmZpgn4syp8RXrZ8K+EWdzJ9qctiZKCk
71TEAwMU6ijDkLeYRTmAT3FN/xZMiz3OmJsMa4+9jMJ2+XurA13Hm6mZ1pZ3
2fYQ0qIWn7v5BnjRMOAnSML6uO6NiUDX6o1hNgQnyAQ5CaO8uwHNGuokQvHv
I+3Qeeonif8bM3MWeOKW6ViVRwFwHUwkJNCY0L7iyCMvQQTR8ERxcxzeUkZS
bHgIb1e9SgGt6P4FEVTEKS5PuB3Oc+0zACS1MpEfWnOPzY/rNDsn7tLaCxTM
D5nCIqvn5xygLzB5fEkaFw65m7bnihVKdpuJbDnu2hxQPMxo4HN4cW2DIqKj
FSXf1JQCR7I0akJBjm8G+2cj8xQ0a4bc5vXOHNSBmjKmahR3d2hmX1a5e7hH
tFd1U4xqXDZdXmbEYEafwuhiT4gCURXBaWvL2pa2dWUrwk6dM1pmJOHpTiKE
8fSSps3N6d9UfVj+HMRKuCrnLx5uHBx+stJHaSoj5nIsBeAsxemDJ9U/YlQJ
bnV1Ti6qFmH1nMirW22Sh9b6NBZdP7YsNY3XqjCY/Hj6z3uzY6Ure3fmp52s
k/ZHvKNH3g5m+7Y1FtAN83c/bNYw8hO3NhiIQ9gZ+QPXoHONjg/jHuUZQv9k
H+Zx3eijM3FBqwe2tpSHq8WD+TlQWpb1Uk3qxNQsZM0xnsDbC4cP/tNCurwM
WOe8vjQhvcjlcOkKC1EgMGpu8gvLZl2xITeg86lZJxpmUULS6aE3oY+74QiX
tczfZCyqRqnSgDDnX+AEotKzfLT/yPuHgg0LSnHCtUTwrAoyp7N5h9XNAHTS
y2iY9oqlI5abMDXMLvltQHFjSZSjJu0Gz2TtBnDoKUXcuS33oRPzASJjZEci
MBfoQVboprhgt+lHSBfjvwsK/etJAM2x7Akf25pGbLujDdDKaf27u2AcfW3O
rJ3+ta4mTW3MoulP7OIUFB6H4geLBSCrq7oY1HHcedD2IgQB4S7hqUpjG5ib
RAJZV/iKyp+sCAjuAnB83gmji0T2VYShkfEn2wef/vcnP2eG5kUeWtWoEIv5
bwnBuk0D9Cm1sl0QLuepLD7wWDkdTi5ZAaryRrZwLw8qhrBfYOE+gyZ23U9m
61JAG1cy71Cm2XL21Gm6TiuceVb4Mh6AKvILLey7HT6mnNEZkHMS6A1BMhnv
UqFx8iWuK3olOK0hUtwj0alLg8LJYficLKtbu4MlZZGBQ5TJjgpjDybTG4kA
5ChYzNOev+RppWRW5mQS65ob9TmZgNpPgE65Uu1PYH2L0KfF5yYyUCw7r5hK
STFKF6PlwOAzuv9aGq6PjObCgrmLQuwISJWwKMmcnzA4DGWK5gGCmy5dj3Cd
hS+8FGeuOTOjDBX4Wna+bQ9wrr7RgoyJAdQvxT3pmkQFfvzIUvnLdCTSuc1Z
rPRmhSiCD+F+hJNoD11/mtOoNDR6zAso2VV7TNXlkvoU6/MX3mVxl2SGS+K5
YIzzpUU06wXyQADJnYsiX1QwFdPAU82eD6RDgFmFsMv8+RdDo10wG4YgM17/
zDArHVqfh1ZzxQlKM/RCVHfF1Q9hfJCQHt1I7rzm8AGTIiqBlnKXVuynfEtQ
vHd0LgBoc5rMSlCLu8cPQ5smLEp057cPpZldn4METwHdpL/dOEYnXDTK2Pem
dx60ieRBQfdo3PiYSL/z3UCzI6fzaQ9hp6E/8PqIADWe8pp/EDquyLI2dPu2
ZAE0ShQj/QuJw6Pcd/3pAhmO6YxQv3qFH2d1QpRyveA1SzkCwtcx3ml6XVAI
5oH0mHaBqOIfZqjfSWY3YJRmXXVTD8hJCKMiuDkwn0fBAjrBcVuFX1OCnFWk
zEt/NeCMZjXCPAr0kB0PSynNm1T9AHfLpz/wHyFq19h4ZCRo1ju6RGf7Q25f
HvlhH7c60CCVPI8oBpb2eclhmZJmnvigzMMCFkYURPLA5uBHKGx3guzbTlDa
J8pSOHmIOYLmmi0cTyOnDo+3x2bBIJ/CrRbC76QavaHTuOoVujx2V8qrLVlV
ucsz9x89MT0Ar/xLOZhm9QpVHL48upwvoxGnae5aGfJ1j2bGtJu/xQvwLpjq
fgJKfvYGOV/WtnBpF89TaMAFdvplU3vlTsaI35nx2yJU8UQ0vY5lSeRSrEKb
9MJscs/UXCTN7a8TY9pCqvUpkPfnwEwNyAIo5szEXzaK21GQ6SO6OB8zjDXH
1UNJCukR1QdY3RlvDAGibB3720qcobIB+EqC5ApXpAbBiy5AyKSJjo6qCQHK
8VGDfGZq1ohNXnhPVKF052KO+/hJzfYym5KIRaKWIKVioAOYQLZqO9hz87jS
DJVXYwSLZrwrgLy5sP9Lg0Z+X2EO/itjVmEtzKikaRKioseZHMBs28COPqJs
O+X/t3MkAPxNzl7vZBiDbKOCAxRc28vMkgNQFFpPtxDJyb1LfR80TaK8HPiZ
Fn0A0qfxRFFPqDrlgdJBj81BUnFbHtBWiaNzJzjfKczmfCAlF6iJV4ALybLl
c+P8mQYgnx2i2msoUw+ZQ+j55v28yOMa6HNhY4JrwWAP1v382jMNjtaziXb3
wh+egujboPwOi1r1/RXc+R9iw34Rq/AJf8OXvonUfOzm0PNhSe+GCieF+YNk
BaSjy4KMK06BPxupfiFQf05AbP1LGVAd7jom9ap4NaVgHDzWdrclfXNOaUoI
7Qo/uaqy/0FScKM4dNQ64Rqvh64GeiVvvOO/3Ts506wZP4xosJU1ZkGXVrBx
AYhqJikUQhg8swnC9AcJVJearEUQajONnN8egDO3BtHUGUOSrPuC7YJZ2zHJ
cbL6y/vhYw6BJmfB/Iuzl5kCEsmFRGcfCFZWEJogcFk1I/KSoIBW8ibHBjFy
MC/fn0/V+xYu9yjnmTTbNpH3NhsWLz1cZaPVEdGnLf5kkC0DGxo5xQAddt4m
iD0IoAWHgewkf7VYSef7xaulHe/vVKhi9eQiqIxbgwmpkf3ykIxj7/KZX1Hg
tTpRHnnlWHtl9u9lIqPCpUkXOsC7tEySQMNMXIvQJLhoHKZKhg7+mmuAS5GV
EQiIGE9mopqcK4hUvMjriQ+86MCVATcSHn/jih6mQLMQ86wWhZtfWA8h93O4
lI2RDmIpyIIEuJ995tMSjPzi2JfgQR/lcgwQYEtOfowc3+DsI17lznbVRUcq
dC7PjPnHKC9O9TRcG8tdi8YItTFDATu/PePg7+aeslqXJ7KaLN5MVz7IlFfU
eWdu9XpXw79seE/j9LImRy17/AYSC63beJsZI/2kaV9X/mhe50TrqE6sxKJ7
k+fY/oNCB3bsPKm38YffdTneBSSaUW/voRS/n5ESuRgU2w4Nq5PPbFT6TcwQ
D51mipqMrgcsC/r1GplMDByBhGpnfR78zgcc3R4aQoRse/8bqNNm+ZQPHoyB
zLMV2HDWOYyY5KXR4kf+UwSZs6Bg6fUidX/qAYziQJ+7kFot31yu2hFQoi2d
CGryDQI6lkJzLh0I7INdPnFhsER03C+VBG+sAxMH2mfDJIEBDPJ2luLp742r
8RfabWAw3cFKI5IBLz1i02srQQiw5BPbTjBskSCAd0arAA/LALHQwoQJztA0
gMlNh5cbN+UGrpIyrPft7EosImbiiqZWWMgUZfl1mESRUP0x8Ww3ex5fiEGd
ISgxQyTVOmhk7v5e1kucFCcqvZTkY2rhf6HnH04TgEr3Dts18T2fdy/MYvE7
UJxeX58PtbuSB6RdKRx4wKeMfXcIXZDPa19EyjZmoWe5EqrMDpc1bzaAxFmv
WsOAS++RAm5RV3RLISF9LWPmVNf9apjGBVxkLtVJaZphoFBvadT9tTUnIFbw
4kqPz3PpYlcNhxwYVrv8sYHL3+jjmCzlGk2OVqF5g2uqc/iailPDEXxCU1zT
ZLR4g22/ZeE4kiWC7NtOcAU+lS8fhRytEKKvEn2zDygSJ5EvgbvemsxhilVT
pkY5mjUBHUUGvMDaVWmG9IyjA2CqNpdmp0zPShmH//FjqG3Otvd9F8Xj2P9b
UBzwJw2WWgEzkRYSgQ79SquxCAY7qh5tNN7v3PqWb0wgl1RUGcq6n/cVV8Ex
miITyb9emUJMfSOeZmLc/MZmb39uPZmPNKqbbdobB+ln+7gGCPge4lNIvWAX
UWunbVDTNIAAEvBpSlIHoe67SAihvNgjyKRlwGmiO+tvaz53kMqSCipPoaT8
XhHopImfET6ruhtYqXQMytt8rSrjB2dp2+ViB6WYtKiPqBneuc0ef/tlgnAF
C20XS+YVMBm3zxDl+SLqxU+RKoEYTIb+2jKWRCNr0BryiqhNZEWpEQhnyX4Z
1/Q4TzRbLrKOuMfGktFa+uJET8hJvh+P/gtEeSS/5Z3VPqGX459dGpQigB9O
Tnlf1r/Nij3bM3By3e34qbrsnsRmvIggnSDVMZE58KMoI8xXAbVh7gJ0+L8I
3PQZ3Ui66AZv7uYVfUv2In6SF5yPdaaeuYJaOgaRycxDhTp94xzd3ZICvZ0D
HG1j4LTUVLsB0YiurM6CilUzGKi5zHT0MeBd0BwncOcv3YsRTUpaqk7fesa/
fjvYemX965cIMeQWq63/KQuDbgYU0urCgRX6qATkG0l+AfNHEnOMtCynjDhg
IVsQnFu+eXlRs3EB5RguKdoEP6KRaaM0bzOfLks99b7RFPmn0TRIICMB+oh7
qT0eC1fHc/2Nv8hgA7gra7/Wjh6HjRDC/vgOWZUg5HWq8qzamI9Ou+JrIjnf
Si/2EA3dZh1E/lWqwuad90+ktAWjEwmtZNaT2cx3dactJCanAGlp8m2d5DPl
9PZg0NOzOzenGKCLrALNJcCGEqAZgUtNKAZJ9MpRIhXRKpq+6D6jkWWSF9ws
9BcwMjnaCfCn4XJxYDsGe/uiKKtrnieq7VoKbdRSYXOjy2Ahs4iELxUVp+6p
8NGiOdU3OVz96CB15XpfZSa40FNKQQS+ugvHd6w+rNF6Ygl65DOXud+BiUV6
KmNm+nXmsQX83m7d1Oxec0JO+Uw+u+uY8cmSxXGqhkYCan97R8cJW5P9F2DE
tupzWp9gzJCHyecd3PPQVhN3zirIJe0Ywo1XnYQ0uBmEs7Xv3f5OILtdnHqR
9SuX2Mj0LKNLlIGkmwBPpNIVOfXc29QmMm3kmVb8f3nLNPEd01VLDpVez7VP
tfD82l3IKm55I6xH3+bvrLtm2pC4RlLQgPgyzFqGFgptYo+wWa3d+afZWuJi
vv0/xWJeOlSmNTkUE0Cp9a4V0LaxH48OPD0c9P1+YTrJwMw7iqA7hAsbwBHY
iDnaqVHWufwrqV/mr6mHsSxM5Yiau9wRVVOzcid+MSVSda40hbOz4JTT+Spp
ij3oVCyoopVDu6iE7rvDoq1g0hZ2XSj4QURTXdAqFXYRU3gfCrvtulinExKh
3tV8KO8y8mXJtQaawh/JyHkRwJH94Tn6Y+ANoHCL1fFqmil4M9vMKYAv+bRg
/uv2Ny8X18IHW3xpXpiUuy+Zl6z40DDOKQXo1qK8jaPabzSs/cfYep9t1bgs
7dQYQc6COViZq+2WuFd4RN6FmOv+59Z+5Qpj5/sB74TyygBrEaGZYQDK+MIl
7/ETXgQZD79bJ75ZtFXEN6dfKYeEYozUvjoTBcSz/pyIYX991QhVuGnketr9
mDkxCnN6Rwzj5Z7tzTl72mBc9zUgiooxPlRIvT1OLN51tAUzMKil92Umr84L
+SRYh9AB8zT5pgeIIO4Y2CV3l3Zl/8+ZVQ2bgWN5Psq0TdbhAx/jr2EcYvcd
PThA8BCq4kA/V7cxz4IP/gUfpCCn+w54UOyfAHTxwidS1HAAaufD8AmCmidm
VIibsdFBx0bUd10Hj+qnPOIm5tefKdGXkd3uJXVsQne4exJiGJSB5KwbzrdB
QHs56WpCMD7QStwRDl5QN4fhlt/xnLlmbpBAIsPbPS4uhboCNpQzGZMy8BZG
TiBkuz8fLVpueR88BX6ZM0tIKrS/OvUAZh2Jm6/Wn6qF8IrD6/TDc7pukSm3
7ypnDbVTh3rWhD5+8TaaqoJVJOVjlhNF5FIilQGs1WrIBobsAh2PkgAf/ldu
zA6OGz8YZRnRG8FwvTTYJmcVFc5b42h1dRYCS8i4L+YstNCCMpdCxQ3Yz6Bs
8oIWIfkaCIR8oGqYrO/fOKtmGuD69xB0HrRblf9TblGIExTDT1u/YyET/t9r
ETiDrQZEWwP68f8+WySQeHzqT+pkXa0lEWUQhxQtipU8blG8N33VS+CCrQ37
JzV6XqTEgOs4cyuTBxM2JWFDVAf8fuoLedatGe2UwM89DVXuhxIFvQ7QwduZ
4zT9FbtoiLpW8xaesQi5eW4jWs3azAlMxqy4AQFO8mveu+KoIpM0eUh9xBJl
jULHxSXrQ/hZ9Z+ghZhF6pii2gqafL+CiFaNqfoIZGcZ+c+nvBOGpYrynwyd
266hW9amzTxiRfCZw7ryvw7hSHkRGqzHXoDr52U2GAI56dh0P2B/9MbigPck
BScUIl35O1lAINPlZ1dHFkUuM5iWaA76eo4jWRfXRSaUyLtQlG2x7u9t8I8j
DzoNgHQVxEOqBipk9PHDJpQn6oIy6N0hlqgaL/mHro8gawM1Cy5hUUsjXiWP
FQjjda4J2S/JxcpEBhlb1eN9/YzWFDSELpmUFKSwdsZLsT7yj3QyNIfYrafq
EYGgsErSvoy+nS55MJlhdxm0ntndafiQS2IlS0FYNdS9diAq574IxjHCpMZJ
mtRP3HW8KZvB4Z1Riky4r/zfltViAcaKxkVXQ+RD2n2vNPv+yTcDmni0ygdE
8fP/hawSUzYLpFnKJT689Kts0CYT7CSwFOCmHOLIQIsPmGCmWIyAg2ATBijD
nVokAWL/12YCIR7yIoKbJeDz2qaJHhzPVYDcnqrPokK1T1taeLFyfh3tMs1z
yeVBWTmJxHRUtya1msvuKA+7hePI4Vbo/x7x7W215kGT+TAtTG40oIrGe6WF
nrquJdvYAEKknlR9XG7nSxmXlXPWgpkLjIdIibfBM0y2aJ48LDabgCl0bXHU
lf4bZloGKaRuBlzTdPydRQar0sAMrxgn7SGccjYf7+GjpKcWnn7O5dt+l7qk
iK4HBN6cguwsyTHgzi1CZtVGFzfcXnaDrPXYjcObWXJOjmzsADEUNsSN+7PR
7EdSGruAIGUgQwEwfHulfyfl/P1SvtatvB6Z96G9tAaXzeZfhOC8uGyZLGRp
Jc8a4CiZQt8YhirmslEGg0bOFUCARUgksMRFT1cvGPRETmcVY1lkLy36Ty5f
XS9UQkd5GYMK53bcm39dJgJK99CH0c0TTwXOEEnjmlY/vDdreIo78gWXV1rt
3YMb2cVk2jYVCJUatvPeVEpjj+RTUbUIyexKbBCzfs86DoO5pd6lthI764SU
r8Z+4yYmsCdNrhgboeKbCjVebCFziLsEaNEibFUMS8vzvEQV+b87Z64vWvvi
PQ8r4esrc06ArCAowTDCZX1F2WbCXuM755rTWkpexgEPoz7uGv8G71hntRhm
kzbhhZ6rhjlnNGukIm5+E19c5oApPUCVUBuvQPPW9ZwX5IYkxdHJTygIVGjW
NxY1m6JqbwxzuCYE0MLWRWT5QayTKs2jMrJjvuf3VfpA3qXU1L+E0JqaSa6G
VGcCyZGrsiDeZ940+YJoVVV/HWjwzEhfBRWRLJ49YZnSIeS3dlJsoc8IbZFZ
810pbrprpUkNa9hDF5g41y9PxEF1nWy9Nm9WHvH6BVImq29DV4PHmsqz+83T
O9/F1J6L4bAzbyROIbiXR9ct2aXZPfgPvkkzuhtMC+AU9H5p2Frs71J5w4vT
WiS2tTZHR2n52G/MgKSHDPZDF0373vv+xX8c0PMSb/a1V1xHssTdRgIB+uVB
GBRCsv5mvltFJ+eq0umOlfFSBmJ7K6qLVA4he2zwsAyfl5vdBpovKlVWH5Yd
rtvaw1K2fI4dgYbgW66Vb+spCbKjNFWjz3IxzF8ssefcT4X6PF9zL8x9pQmA
F5uLRKz5Okim1kiW0LMf6I1aPmVMYdb3UPeu4FI3mIoDHu++gEmNi0b114d7
crkKDmo8+kKwA+sZ11UoDiv5frnpFIPDtifixNDtekYmgNfshvt+ttyY+3jx
wM811y29//sdGf7Tr0o3oQW4IgottzJCeygiEjZrAqRiJ1sKosK3tuhWTqC+
fijczlRabXPNp1wdH5QADu0iw6T6q/o6BsSOgpXuo4vexHe+wWc2Eyiis2+Z
A/H25AOVH32rRpyQS3cFSaS5LWUlCe64X3go6/CpnWIY0PpsvRzxKKFN7bxt
Ic0uJJPUdXhZYneTwsjlGA8dh3BvUoZEADDIJJxtHZ04vIE3sM1GcPsyEYZm
pAy4509zuk+xFl+FS3JCGl0uT3yRJmLKB66lPZ4p4aQMeOE4Z0JX1D4HCt13
Qwlw4kFa4C0ucM+//xNIrYKkX5NW7t6GcfiX5Ok9DrSkeI0nXN1CAdwTnEJY
la41C3fg9HEumyXscV0AoYapi5WjH+3vnxhgghiCDQKfCMRWx9pMA/jI7iEE
H9hH4JvpO6cIAIk7rrcXQJLGURZoDjdSl20z9nCOVaK1PdY0C2TmnEqc2GIr
ymu75fqJ21Wy0J76LQRTmK1khUISUrBZkW3fv7tMitbHtOyaJ2iuSYwQMiiR
M7V551E7zVqJYzava2LKvfdnMTQiGqiETf6wfQjkaR9y1JlKrWTHVY6fq4Aj
E8fzfp6CeiqvxaIH7gOoNZa7Cosm8B+3FDclNMOvBXAeQKxH6KNH+EFLjiDB
yRymB7q6IfFbq4O1M7Fb+0+1GqzO22HBoP42OOTP3yCnz6x1VPhulnuBplGp
A3QysmpDWdVvfvQr36ULJT4B83RTWtY3LA6b6WgZbf33MojrP6L6mgT93v1g
yC//35BvgLc8rP57AoDa+8UaQMZ2aHpZR06u4D6f/A6M1ssEnBNy9yWZoULj
p0+Ns5/5ba7YVNny6xxMFWQjFuBdjpITwBD/r7TuNdoIYRRMTqd9f16B4Ly+
ohqUxEPIrPM/7+pcYElwmlizq4GSMXWT8pw0H+4NFnUF/6KjqdsEVkGFU12E
MAw/KQXvi755vGHgm6EI9J1nvlb0q3OdlfhsbvTKslXi9PJJo5QCTs2JrCWk
kIwBCShq+MvEB2xwxk4tDlFnzelNo4lDIU0TrPRvbVs/ctCkvmCF8nzNIh/C
qsGScslC8jbZzuVfDPzx5M07/LtUJLE5yee/3OCXOu3nycL/YlDxR6S9Z+lK
BG0QaCsWqadEW5ZPSlq85lwL9zoMqHaxJfrv+rIwEG+mdHSo9tiVY9bpbrEK
lCdzyAv30hq/aRoSAtz+eGBLY91SbTwX00QPm/YEx7k93w5MS6nYHC5cg/dM
PvF4L8XSFDJxdBLizhSUf5U4wwpsVeV89X9ki7xw3Hj/9z7lFFCgkkcxV8yP
o4mzP+Ul2GjDY1VEu/kB9812yDvbF+duo/z3SDQDfce+zs3f316GM8JTw8Of
/CMwpAmcOpyY2N0EraCuAons/X43zNMZlnPMU3kiBYMLEb8x7aBCul+qhO9c
dz17k7+028kOhnIBak1lIQT2Du82F4XbbTOjXUd/lZjxl3+JKTRqaGbmn3MX
8gYAszeSEO/DoovX6RsvlKGIWmqDL/Q56Bif2w/GP7p2rd7Jp2D5qMyatk2g
QXeUesbZGNV2nijz6UJfJ3ilTr9CR55V7/d6jaXQeCYs1IjF8zR8J46wW7ys
BOokqnn1GFnezR3pQwcqxn0pSM3XX36NvuV6yauELZdftoaCGR9KHNHumAbw
R1HvSbL31l0nF/yd6Rr/ppr8w3LCd/W+a3bM4Dj/fnXztTcrAvrRfKEYLGCH
W0EtUSyeUBR18PQpszDjAvDxEe7k0x4kLZtgO5Szm4CVl9NS7MRVJB1LnH9s
pQ4bHHq/iwN4SdQObD++iDoxgC2F7jDY0qdGzXoQeKpk5RNAnGT1JaEGVOfr
lM5rSl3QGi7+OYdvm7eSS0pTmjEt3tDOBipUMImBVOdvqGi4etTNVwoMd3uI
7gul9Ll5tlo7xp5Wi8quq8KkrYHqH7wvjBtPII+QtvQW7x0/82vHQDSoxPC6
BPH/6CD1mxHxo7crNW/IrXRITIbC9B4vCnEL7SXwLivjtnnKp5Jz+R8T8Jwn
gShas3ME9Emw1kYzaOYJ6JIQvygEA/Tjg3TCu9BXLhZeV14Eb1GriQTVlTiH
e2eMVy/mmT1AEdWsJQoV2JX3R4lvZCn/HNgB2a6Jk9Nwd14hN6TIrKhuVdka
F8y/Ee0kUvBk796ceh8aKsWSHGIsWDPHkzY7f3VK3RLutppi8isZD3ZgBq/y
MTRPMMmB/JgoG+EKR2+kzPKBDoTC6AmSLaDYHljwpnkLHRpc2Q95juicCgpa
ieHPkpNJza1YOH5JypMHqb2VPtfyhK4x5Lp4ZCpbExvXuvnC9dbia+eDVtW8
Ab5Ja+QZENBvBfRPlffiWDOo65xSWAgZyfch5qqdKwD/1RCbcgwraXTOLeEc
t5oUXSrUazwx3IW1QckRAKFN6rJ8pE4YeiyAZyGhCdfc42gSxyctuHmk/o3V
hrG5zhsoNyLX1uFnkgu+87bmhFqfJh7E7+XSNuJfzmUkB757PqN8IY1P7g8R
7rIp9E2a2SA0EMmkFimpvIneIhSqSMPpn5II2zs3o6ndyJ5nL10YQCG0Dv3F
4L2hicLoDNkaUBlHCAjoC5nsPy+44PXo429gJyyKSmvULc3s+Rrun4kAEs3C
SU6MN4ii/hzROQVnCGYxGYubh+2oFeeY78jTAIMXuYCh9dUfJGRD2QLSFEN3
HW5naiIQhlnDv70uLQvdy0sPAUXCvCEB9vL/F8bGAj7uyXcfe4GSr1OuqpBA
1guGNvtqruy8tpoQd1laJJJZ/SZOmFe6gVVjsuhjJ56hzSaXJYvrRiISdvEP
As8kDe7quFcQRk5EpsKUGVrKIHSCGHT2CI5HpEcFIa8Yq42+fxePACT6F0hU
7Z5a+y5zohhPVLQMJHzIdWcPEKgFwEy9Tpnn3EGCxa+U389YQIE35eMyqkBM
LkY5XpnUeMDodnlD+P5+7v3KxKgyZnJzg+BRGad8ZMWBQWviogj4sYSaIQPd
1iCROZpYZA4mzqbsvnlItbCheHg/eckUgC2Z03u/azh5MaasNaih7bWgyGgn
msUKLyTohgrOni96G0ahI0Ae5mrP/Sxbm9yQSCDsu9hxB5Q0kJsmqMa/ZwGD
U5h5ZqBdfu7Jie+0k8Lf2Y4k4v+Dfub2GWSLoVoM+rWnIWjaHCsfHOi/4D7B
DTrwMQht6XLyAEEy0GATAK4Y0vD7ZWnJOO1iCNNOrRMruq98C0nP35SuXEDC
+6Rf0shXVZMyCRmss1/jEf1giRpYaS7H9/by2haKVguUsUfx79gwjx2uC3jL
yDvVWgYSqX7Rkr8/QuHIfODysY4QxYsRfUGmAnPe4uHuhZbGCWLNB18Txwcy
ZqGuH4q+8nimnw6eDqVCbUmdhPU+Gz6wVFrGQXTHYNzXIuBIFlPWTsmkh3r4
OXl2l8oKjMqZopviz1+fIKQOSETpullrVkT1i/drNe2L2zlR0+NqBcnfo0vN
U89toCOQZE+sjtV5WW6Xm938FKUjOltG2XeHwUNR+o2jimgkswSljs8/R5wu
HEGRT5NUjOCx+SwXglJz6y8url1pLCH+KAYAauSiVbFDmmkZcTeDbaR1Q82i
DhXYAFo3RMUOvxDgeSC28dKw/f09foTmSY/nk+DhdAnYNMVUNR3wmTBdMx+N
ytl5pifKvIToAn1S2tty2ROCM2Pb4T6VqMkLD+d39tyzTOdEfotPEGZCubFE
bjifN1GJ8WWd2+U7mRJDXCJ0YAnIdQC7qV3gI+ltRrBVTn9+iqBNEFIbLhOq
BnEwbDV9FsVO99RGIrVhT19jfL+rfa+7CLMezwsqorDmxmSKma8XW6M3jmwY
z0A0EoWNGGwwFIAz2Qwxkis2CxDEbR4EbsPYaduuuJlZy12YNk81mJRdi/r9
+FqKE2KYvaqp9JHB9MONpfZOdOEP0neLYUu0jOkS5HhRhanOrgJmdcL05jrD
YwqD0kTeWQeaN1pV8h7pNmgNaHj3KbaA+zMIDx8awkpKSBnR3T6lMqFdxPep
lC/+MePIqCRRWaIWzQvPsnf7dcz22nRAuQ+mGoGYLShzY9ElAb6iAju3PI1M
tIIx8s9UeKEIKyfM9HehY6euyh5G1NEFQpsssyHNSRxOSsfBHLb1omo+ZvxP
KRVwhTq/qfcVCm+voszs3ZgwiVhZxCahkEg1/aOQtm/DJ5eSManGo6/JiCcv
hWCPtrlPweizmYJ3JhvZH6UX+nZ+lMpahWwG7ViiKrAZIFF1Umgegy/JEPlk
E3A2tNCSgMPXbfmRtnt25Di2aikvWpxH6CC+sjLYgagcQ4f3LEzfDnqBU4/d
1K0s+w7hq6xLo/nIfOqdOo8AAzinLABqBJJOxdBChIl0pbk9mVqdNhgxUpej
Z0Y+ZX0QuQXSSFd5oXl4pcM9i+YJKDj9DJOhAW/uBxtl68lv5p/p6xKdt2Hw
taSwAeMe8WI321Yla46HVRtK5fPZknKtA1256PBffzaTdDx1a6U+vLv5lpEl
HQYRYeG5vTnehnsQXsEu2F96C/y99eBjvd60EKme9QYrgkjGs0In2ac0MpoA
i+wSocX1/hEHsx+MViQIEQ4rzEoQCDNCnZCLlpkeQ6OqAQk2oRfrr2Q9xl0A
aoH/wzVY78RzsHr9aDocqMhPp7GscIfS3ijYk3QYPZxkZ/W13GIPqPYnQzmZ
YT5i9qZse2gQuulmZFm43uY2q6XP191WTi36/uxX1GIWHyzyIYNMaI0DNr9l
5H97IBEoviMRJWh7NylyjETsF/aJJ7jA/VLbagb52BRFUWyTBbfwnyyhNxu6
wAxCtC7fQHSdQ88IaOTtC76iGlE5P96+DLN65TH2suOE6Z3PBkGImfNKPCM9
DAG+MWZarPVVZXlJDrR/pugILcL+Fd1t8t+oYRdjJA0wttmBh6NemebKbb+z
HRBT0NT4yoJoRhSjI76NJgCWPXu/y+/50vCy7H+HcQLWb577O2ROUC2KghWi
40feLyz2YLm/R8AWOGSDBy4ekpJDdBiX3DrvNAnvRdXtoRO6+R7c6jrj098k
bKEGSmps7RTlvzNoKqwCayMKw2v9I64XPU96kF4luDtNrWxQ+CLHBE57yYCq
dflwnVsQWSUgyThJFAg66rNnP7ESCYP/8zWcnMpzgliftd+M7YxnjHjzKCYK
HZj9aAA2KNGpjCjTjNBjarkWvrY/6Al2vxyIpByw4PHfIRXFd21QXTGh/A6w
+lKUp+L0HCD+nIg6P4/s4xlVBF7egkPgPdLB790Lt0vROyZyJzwPwfha2DWB
qRguhlP2soqV/8RLiEiiBvyXWYgiMiOsTuvjxg+vSed9Kvyo7a9ozw7/0kUS
Cm6uMCJuAWBhQoq8ZXE0t1KT1rjepfd6pj6xczYzJoPmOll6aS4Be1CbbUzb
TENh3Nw52TBh6ZyHMMNgj0oyPqlpiHHKW/NX0lOTSBTMwNf1/DHM5s7+x4Tt
T1US6bzVDsvA9PWPBmwp9H//FRjl+uBAxvdoxgWSJf1SggrMSGE4/eZzRwoc
20GDQpHUz5L6NO9LtT1t9ddvXOJ9blTTU7Oe/WJQNH9P1b6rBUUZnMDTKHcP
HnmAepxPCHSnlzIEOsoVCtDE13w7MyagzqiE9JtCAhY/SKxj+QnLZgmc/YCe
w0F51am3WOs6ms+Z3m5wXk9o2KkgIlU+1I6dgv05+ENz2X3IlLRIPK2m9ghm
V9wS5yyCduX5Eoqhr8DIsz43QSW5is2TcC9ZMZU0U8DoIW6rydOmKrfmgqjp
igazvpHXdHpQsozH4cUa9IkCFZeWE3br2RqWGEqUBI4aBhWyC14Uo5D0Hu43
JeFtPuspt4pXmIRPhvWGjcKFzX7UtBdqBp1hHwYc6po49E2HRVRhqdnUElAr
b1ft0PYuYlrVWKfVkuU0ZNlSG9saZ/vjCZEdHvGnFr4qt/QNGcTwiVsmpbo2
xMtZHHpBCVSUy58jyL2vwKqUJA8vVVFU6YVPvLH/A2Y28xoWLHR8MIY8eL8d
0Z3qNaOaoMbI7y9utqurJkQGGYzYBuzConwGR7W8bYQag7Rhuh17nF3/qpgz
R4iwzxDn0oteL+B+q0pg0Md564+oglRgJMcw7BuPSXMYzy2pbeAqc3z3LIHH
6uVj6Sh6a2QfUuchHbcmbkL6R0huEQRGXHM77LJTGuDc2RPkg6JBodsVJI/k
8U/i1LLTxiWw6PqR8IAdvk7nwWPCYHVzs4Ew3w9KJ8kRWMzMQghIglt/g6vp
qh5fUkOuTNJJY3AHIQN6T4EDClgD8RTZ6wNWkoLM8MHtI9xMeJCSvkSPtIs3
aiV+laYWZLpB7fZz06oWMbZfMKME30eIpYEWpwHGU//0vW7BM6MzlB0Msh01
xrdFKHoZrLHw+57d5vhXjChsjLQFLV4AZkJ2A9UUBe6l5UeIGeT2GDPNVLgI
pQBhzMpkzY1ic5Spmi/hASa743/eV/H3eSKs4XMWVgBh4ew6RGCH76EaAxRL
Rn19KIWBfBL3DKfO6XKrDr6vUTTj/rd9mBDBu/EGH6V5XEAE0rH3B/H1iexY
j+l9ZgVU2DEn2nrsGovMQ7pVDWoCK4qePbI2SldA59eY4C2gpVu9RmOGjB1t
Y6+LffzSZPdHu6RQaKUttDhA7SgYDRBo1NDuWvo5WNBvKXYKmSohCcq+LrXh
azoW4w+D+lARCX9R46+ssCyLEhG27PCCMo3LV/d8EZOntTVMgekbMKoYhiBE
rsv6O2Ma6EiXCR1RN/Nyojta8y4h204ls26ePEful+QGmvDvMnBl0xFZkLS9
PXb9m0MRdhNxnI5/Se8TsuOuqH+GAnkwlNG0qFuBIe8IZPBHormffCpY5eDf
Cq5LyzAwk1m1GwyiBGEoPnow1S/9NC1nf/d/LJdqQAGyI+jxv4PFm+7sAMMk
HAWUexlrI7Cv311bVEl6URaogmE/gxDUHrZiQqivYYU87rf93VIZtQ/amfZn
LBw+SfVMG6tKkUPw+89Dd2cJV8s2pSjyZdpqA/y5WqJrMXd3O2hASD8QEfyU
UehKWcGlMzVNcfmumXuMCm6AGeMQnraPh7jJtR4k+o6swXqkVXWK0T5a7ddJ
3pzqaIuYfJjGDqR9Ke/rysBmRO7A2We77duzX2ZSYYCuLKZLn4SZxyRJtbt+
uKYywEHV7ncweSsBfBvJTQNTxRc2yzLKnIs9H+vUo/+7CHF63lOZSSFqnf/2
TMapgGnz81lGx04sppnkp9DpFN7gORa81DAYxh3uxY8qC3j75sobkNhNucf1
MxG8k7ZdEsFTmleREfDfsKj5lZpd/Dec+eG6uP71ZR8KbMn9ReVs2m33WGk2
o+qw9vfWGt2IzpvRpCHO/83gkt5nGKtUAWpmB/GOur0Sr4xvEPaVj00vRzcV
Cs9aIlgVg5/16XP3Va2O1l5XjpTY54xG0GqWSExp5KLHBbuJcHDmVFr+WzCg
Fl20GKkPljosMPhjo+54yLKE1bPOKqhZxTLdpuJQ8s/g3/2tQqTY3plXPI+q
31l9fbzLmliE4Qt6ugYvyOBtG8m6qrsa5vBkmTvO5TZURvZvVLFWhHmBENUC
10qvt7ARNPSgaRM5u14yXtmkBFm8pFnNmN3Gi42eKMjrl2GdpOoHcpABSRpI
lrKp2LVVg7wXKogTLIKPuJ/RaUyYmzgEAi+LZef2vgn31VrXQsilePW3u/6y
VupVVmkKCxZO1iYIQWXxS1pLwQfpOYueP+LaWGrfOJKe1UGJ0kOIoRP0Xmgc
qRRHSsPss5qqbTIRJlak3LEHhp2Rd6w97BEg/pyYEbnSonX+ipnyOfY2PFZ4
umlB97b5MZ+ukUNGbw/L7jz4R28td0owQPdkFw/hsA7FBzvHkszKSI1Dgr4d
4aG8FvWF1NQd+nAG3/o77VqWDhE7pT0FPsLObvMcMdf23H3mQV8shhQqGe4d
VSnP4jxee96zt9FWOhVhZ33LoON7qluNQHPm4NZgXMptB+56FX3UhMdh8D+r
ZG6oKE7sIJVDagugimG27Tqp+YwFlfDRgr0Ck/964wKAxx/gEIaj3zbOJA0u
ijby2d8XI8RM1cmDllnidA5SHbDGaQQwIuqel9ZC7qXXLsr4EE6cPDZZbvWW
C4ae40xvJB0coCGRO0JId2wGKiutmTQ4fd8xfLNY/AfDLSZGmXBKU2Ht2yUe
8YA1MYRiYZMNBy+OABQzXHVjAO46G9WqlNL/ecuUjOD81wwEFU4AuYig8Wq7
Cg/K2t+VAqpeHxcGS6RFWP9xaAtavX7TWiwIIP5f0gtFBGLOhR/9G+QFWjl8
G2Msa6zGZ6YvtghaUZItEx9rOvN6DsMqQxPICwVrjNf58ht+v3RwIcq/jEXE
TorDknGoEVNuWDcsb12xTWjMexvc3XMQc/iLm2RBLBWDIBZDFPytdngFDD9R
0Q24+sS/2/MEnwRA/DZ5f0oUwUKr9cCaNs8Sat2a3cdFWPGiYQ9qhhRbaWo6
Eecd1XJAMwsiCAWIrBMF/Niqt779m+NUjxDYbEbOHPx/s2+Rgusjk6PswyhF
C6enta6o1a2s1I6FzXqlAhChEFqM4HN7i9JzCWc5O1PbWTAFj4lE3nWbynjh
Q9rylTqk4q1OXYrlodBjzZZxXLe6qzv9xp6HrXvs5eN0HXRro5/izyMIW9mw
Z/HOSa0a5zsCby0UrQf4+quDTdL+1QyzgSjaH65G7qZW5lDlA7mIwpET0wdz
l2nd7k3w4T7PE9L6cGnG28Wf/QRZSFtsQ4RQk3SwAqqwU6lZg0LJSa/aaYTA
dBN5lbwn20gVrpmWXfZywzwFoLw1eB5Zp2a1Uz8rmRTL3ERgr4/4ZP5UCmQq
QpcD+yDhM+6ATKRNgxsXktp6qweBcVwidJhdrWkNbvpJAqn1R3VcXV3OMxQx
c1YpQTSCeYaWHf4Fci4rKsDff765XMgn7k8KQ8EdyOtTIEdoigkAj38toWz8
jhAx07TcEMxX6wPZY7ZZu2sFOES78zvRo6f9jvs0yqEI1Fgp2jLBkXaL81kh
D4jyFBAY17W4hRaUKkXqzILxPZD6adbu5jZwun5wCY2sg++7bdqmeNlU+sIN
2jO9h7t7CrczMh4Rp3sUV/MXcCtBhsPMGerO3vKTteNAv3zQ+Q22S77PR6HL
DyppL4qx8FypJjqkyT0f4CyBDXEWjeWctKBsDl124Mzts7GPVFJ7zHT/gasw
eIit3JDtceE6qXc/u+JGJwTw6QF+QJ53agR4i4+GPatt1UcpIpdbO7NbfAil
ZcWKtBk4QpdhdTINEgWbiT7UTt5IuTClsFRsc+Jna6sE5P+1Y3jz0hAI0ek9
/SLVS9hodO3Z62nZ9qQvTH7QgPSpIbFGYDOq6LKjqAqU/N4tigCWjX7+I2vw
Fd0bfZCdTxGYHC0P8qWBUSrQl11Y32EbtD/2rNEI9gN6FqdzTQqHKPOcT1MV
GUG2UWA0xNUvoRDnChiNIEt2cX3FPUmdoMNdDijYsvFD6keET67wfRUYNCuY
/3h3d9cqfpQ+/XTpGk5j5KofmV7XCNHBP391bmpQq1DKhvgq8eJS2OY6bBK3
+FwT/662qHgu038Aqe5adkyxTYWZ8DE4UQCEw15+4AOxPxKzkGDFlaenZb/R
xiFMgbrLKMtUpyTbVkV8jm9Lr1A0RNyaW+irha+zYgcMe29bLfkmD94tO98i
7tQCLHjlgxB2MCfMzmwVTKNRsFxbPfL9QIYEW2r+IgOH6SRjrxsl7MVGs1zy
mzB6f0CXWtJib+ondwX6x5GpF2KcWagn+LsNHJtCysl1kp+Ym1s2daBh0yrn
EShGJu3cS3P1Vbkzv/IZhTPiF/UtAJXW9fsAsZV+JVzM4F3ie8WjzaHo7Qvj
jif+RCIvbT/+4SgTuhrsIBJoiT6DGJPpKhzp5unbTwH0ArO5zHx5TbOseZ1P
jsE5wcWXfEwtj4ZZbr7feIcNnH7RBJCUfzx7JalEdEVdEhkJrMpx6ADTa5pB
1ke3ODrbmS12Ki1iDDDpl9AkB613lhEwCJXRv/FVJStIAWM9Qvru+hcwCKnr
Z+9Y9XccvZcUNX1y185yQTnR8ytPm8qo01DI7n7ddYaINimbde2kJFJ/Au5l
RadXUAu0Rvyp6so0v41Pnb1WBOTfDZ+I2BbshXEmIUexLFXhaQwB4oL4BpkD
t8Ph/BcmktYmDb3FDW+Qq57qSnGfmUSA9EtnOBoUNFK29gRfYpPUsPfEf4Tf
ny/BaNtVLUHp4CYkamkOzeazZ7HMbowbbe7BdNh7NPBETu+Wxun+ouJPkufQ
m8ltcHxXFxJNVEjmoQ5ctKuahffMc/wEWQpLwmUs7BdUEUSNvfhopKaYtsWu
rCVwg1LXqCxO9gUNkSJ9jP1aRGESjDlp46HlS2LoCvd8+As0ZPjH3lTcXEaa
zzWYotYa9WkZPefI1TvCVIGqfblLGrT3qxq1wt7nc4W8gQhv7ACaP6Rkf2AJ
hdsooaIIgQ1E7Ao7TyYasIihCLZUNRnYk2w6+5HAsQKu1FeyDsFZxW40dtyv
3lcSX7Xrdo4xbnOwxcZ6L+/Ph1iQRegXo7MWorEV/POlznxwHXa0zj7qW/kT
DDAzy0jb/6TaeeuFbEA1lOS2U6aztbn62c8qWfTIY6XcLK2/XOk2C5mJUUJZ
b/QvZtepCBKx1hhiIBUN4avqIkOOW37hZNyRYgqrXYesotBekGM9/AsjcWzc
CBUrlOWSTvLVce1wGVxZ4/MyvMdzlZOWEYWXZnIJo46uPbIBWJ+iQ0T5RBEo
L5k9Yw0RvLfKyRPvYsx7T06ytf4lCxD2PFwejv88/DIMthuhiYD3zrxjB+wN
5Ju2hfDSKHMMRSt1g5jsTby4DqLrVUbcTDZsuaGzPiVftoN9DtYKmieuJ0YU
Z2W454Wvb2hVYyw+NRlmzJ3hfDRtC34npQEUEsbQqVcZKqzDKrV3VpLJvrRm
XiOakFJ+LKv7oILDVa68ZOBYEsuXuhAIZjfZ+8exop3WWymqW+mlWBu7d+jv
TAk6jFdZFLAq3BVu2oKHKuaWSBpbqsBGROLk+t7SsvRccXIkr3PTy4bTu7xc
U670aVZukflP84cUR/ecNWyZixmQ6ZyzjfRAf8yLPjcHvuD4eua9pRxmdN7V
9kvUjLW/t2IjB5xDjqeH9ebx16wplPjGbMf+aJg/NYRS31kbMsdPXyKKYHRb
5zaVSU3NNVNhP8WgK2gDy/d3xFn6rRPrsRc4bDPNxpR5tV2cm/yYXOdVIZRq
xV80McoBzjxc+Mi+sbTjqe9yI26r1zoA0Px1/caUvj/DyDlJXM1UCnxk3ALM
6/n5F/O6e+2WM77eP3Cu1tRa47UobyvWJZW/gIIwJ0Stp6COE5l8K6awyyau
mQAV31BKA0UvOCBX+AlUhjaYQYUfFbL1Tju3JmYbOCOX9gqxyigCaQJ8zAUf
FZ4zvrT8ER7eFoUiT3wKT4oU8kh7hj721yCEXyi3CAq7HQZ522mPl/n/rUbt
hfS4/CQkQTFe4He13K1CQVvArZIy4F4mdu5Vg95GXWjJf7kdhGjSUCYYFeqr
nLUBmstEL64LnfQZHdGHzJvrpmwMcC7hKTk64FoK45Q071d1ztQXAhxvyUMl
4O8N9TG4Fy4cy/NhC2dPpeKRu4bAllyN4nSNl1TbM5wlxwpO/WI9pmeguhNx
aWuwMPtkVv9u2BCPV/eA6VafvWK1ncTWitPuou+elX0Ve+82doppi/wS/LmP
O3vlKFa4uFku/aWIqYOU84Ld1OGdrdEBeZcmmzoe2JA/8Fn/tiCZ5yWPt5X+
EufGIPgZmh22voZO0t9w70FRxeNaOu9B/nuodwNuNdty1BcIUTU32XiWZ1SZ
7DGyMVEHZ3mCaKaOFEw+9xIcKQhjtOfA/+QnfYaLLRJ5W0JNNLywbsoMGuWL
28XdlirIs5jRncs7+c8V2uNaXN9OhBxCBKdci6Bfq+dZW2QXx8UrBd0R4evg
ffLtiOtB6Ui6BcaSUi2ZMdwb945IoC6du1LKIjEgBPG01jy8bxbthGJcHPup
uPeIz828a4we0DBRt1lZL7zQjwARpiZcc1W6y1YEXtatfw2IswgJII1ZszXv
AuzEpnoiW7GWlhJls7pExrrg84S44I+WPPJpaW4oOterswLGccbYyChd5pRF
ZMyHJ4AilRdZ9LWehJvz7E4KsDRee4VOa2tAL6tsHHVBbH7CimwxPAKrh++3
8+aRLuaMgRmgAK3e0M5Uj5xE8NwKlR1v9RabJcO9Hzclp/3LY3IkgxgD5IYn
R0P8b/o2FRicfqhILaUX82nSZiW/O02Z7bvWzVwwXklb1tWnnOJa4ZI0qRCZ
YIv1A2Zs8t9r3EzzsPuqrKr0M+TUkRV+YmKOSeqa1iyN9pFd60AqwYHgrcch
c1MF33/gsJfjmwLZeFg1Kj/j4bOvSOU1wcxUIRthfFFJJfxR9iytxcvL6aKH
5z9HNwFIc27uKAHY7rRF8Wz+Dv8Zxo1nweoR0abKP2SEt/cn4oqiejlRw7wM
lNZXq6IQ43MGJ5ToAmkT62KD9isFh5DzSZWu4zYf4Kf0H9Rn/wC3PN6k8i/h
W1PmUMTLHjc42iBPgLon5LOI0yUKl+9TgNHQm9z0t2bqXgvF6lvi4ttdwRmB
sRtzKtWSU1GT0w5cnagO4Iyw2eqJFV62JMqbVvIkQrp+rVvMu6aLKrkaexa/
l3tV/cvu9LIVN1jCS20ZFuC1i2m7ZF0z6+TbyuBYOTAHKF3UzyAgIiZJo0Ta
48rVYwlc9h1fBUQ2CfPsSK3AAHlgNJdf9aMugEGHnOX6cOfhyC5/3lnVHxxa
SfQJxbB5GX8tSR7uqvjUyAMfLiUkv5EtPiFO/n8Qq3DGJK6CRiyTdcj7JG2z
k2y1pK33ls7fK8tBnVwuiGtnTUf6juHxkjSpSf1ZkwzU+H/O6pzG2KzQ1B+y
Wj5lkB6W65G+6Q/dsldY5hXfwhmqPTv36bcx2BtqmyBh+0VzhuBCCWkQgBCG
SEI0l6ot3gEtEFlvdNz4t2qYlMCooKXP6jtjzh1yQPRaXw1f7aQnf0ChoOUz
suv8vEbRnqFt6cmEQKoxB7RV8ONSVpSPTVtMoe6kh33MErLO8VHZ750xNkDB
eGHLYJFmTYNLT0j31KQLSQmopzuUfVEbkDBEjbcmJRlhbq4dNwvBTNoUAokN
oewpswxxXReZc2t8AzZiFBv2ifdG6uaqVZB9hO97884sHX8wmDFz/wAba4zy
zruzItG1crP86/YVMKyce+kf9ppFJDbUExCJ5cgoV5y005tTO1sFc90xMWdY
gvYWx4lxUigEVwQgVhFYW87YZWapPsZKo9K83rthaMT0NGOqCGQlB6cLKhI1
Ex9HIxOuKXfWafWNYLgjNlFEEW76aDA6FyP140UKk8Ssy7UuUTl2VVlIGWHl
X1sraZMVEtLUyfB8Nl9oFUSR2cr3uCuCTy8uW4CVjoWDPKtGhfWc932c/1+b
73v0AmqqY9KGqSUD/hlWzjnOU4ABSHtdKY1pUdDrYy6HbYjQiTjMyglvgcSA
Eh28uwgrcFIUdqlnk0uOEYkY+lkcWKQjWO0BG3Amp2L2hAjl98eQzjd8vSm0
iv7xpZ6hAmb8r0FtJr5WNo5sN51DnpSsm2uzKWezIdRDJNAe1TLS3CilsULw
1fczGYNH+bcJf0Zfz04btF+zVnkma4iY9dJpQpTiUVJGicQNGQB9CA/dxcSv
eZkU+Mno6/wes8Bs+IWbdeGxbs1s5VGxRpHWp0Ied1gwRGXXLW+ee1oWN7W/
YH4zbB6OQyk+UTwNKelDUvU5OwFCbehCImgAxtVl3nu2XK5MK7pjLOM5/SfI
5DP1HjP0R2jIkQ05HVEgMWfaOb5rtnbYvH30xgdtE0lhoiLjubHMJ7crzwqn
ni8VF1pQ23HtuP3k8kdENDB6b952AJdctRk7ApHtL1rPhl4W51QlM4XswD6A
46jUMDnUJMZgT8fed65RhSZRc4mptT3CnMWAOvC9XOcbrvfG1iWvGfMKSJ+q
xkoUXIUiejXCAM4nIPu8V1Qbt3daGGRX2M4MZVI4M9EzR3ODG6d18/oa90Co
rMMMwzU3ZvUEoqP67eGa/Vcztx7ZHABzAYuU71saIIls/Zd7thu54n4kz5IY
mzS3xv8wYgXJV5Nq6xb0L5vNsrsgVAHwAT0m6c26NAqaXG9vDbBep+RHSf4G
GZxMPLc5Oiu3ZeGqijJ3Wea50kiuGmovHWqbHjNCLJFZYX6UEaqFTxDD8Msp
L92UPrqfgR0LeGEHca51P3yPHglktKU4JajfLFojoJ7aNNYV6rjn4hZXf1AL
hMqs3uHmpe2LsPX+9yYzcA3oyBJLd9t8PGERpPz84DELLBQqXpPcCPijke1y
WF1B82ZAnkLvoGWYvanmwyHlPGpTKwS3NqxyB3Z8CZJq5EQ/ox5ptIFLn83F
ZsJ90Jbi6mdLmnA6vLZakJOmzaJeH8X1qE2VwpFMgVSMTzWwFHHhX39IhEoB
oj6eCSkrGmM7/EsfxbF2+ngqRmNnKR39kOwIAIWVoiw+2EjxSHaZ2W3zgAen
KPQwcEGsYzY7uhgqMucucMRjJr5/P3j8rhdi52oXX0BPGUbh6oBUyhOAXF5R
CxciKVn7Xhb1UxoK0OEc3pdYmn/MKrhBhqFS+lt+fs4yhhl33iKcaWLAJz+U
kIw2Xlt85XnpLJMBeux2YAHg1rlQmAD1mbtUHJD3W+JXaXnzVF8aRGrfqWKB
YPUdWScUZh622tIp6oQ2pLrNLgPLSRS3rdkbEZE/GCM6PYe6DsIH/s94R7WD
aEJwcBCr7HjbEBz1Yg/KKoEq1KrAdKnNk2tyCjxAVujrsZHIyC7q17biWctr
7oOI5dqMAN0J9NRp6pync3+713sC89YHbFFdpzRDFeGa98ZchXLEZ6k8u/Bt
YwAo2KtvDyoA6R3W00biEIjNvtvoQkXtzlEYt4/nixAjJ8Tp5Em7XmnX5t2W
4I4XN0BHOSRqrxfj92qV4yV8O5k4yeqyxfY/VXzjaXI59Vy4Ox06Ke2lTSBc
S+A0Tl3WwpLeMIY5iNB8pFK6vzQLBdpKQKyC66U11TFleeGSaxTD12Sr0+q3
jHQUuBcqaxQKNjb0S98Bf9IM56kqkVccobg5deWM8/rJkJNJwRUbL0yFtetq
ExVzNQkW8or+C61crE1OadBaosiy2c9raVNqn/qbifWNbFWZiGTur4Ujz8by
ZNAjBcFBJmI3hjs0NHrLjAEL6GHPAi/0uQ6dPUBEHfvsthqk1w8cPONCfgQJ
twRpIP1M/4GWg+fG7yYPRlOguwLyLyySGkQm5mYQgeyBYwCpV2KAnlisqJPT
qeqBb5gZ+kACkXCipfivhlDBK8u9MD7SHQFFU6yMQMmfqSoer4wLU3EyYjdt
kibSOjXPJKaxbJE/t7rH7OchTEf/e69NM77lbVnbz9oAGJcneZL8w6o+HB00
raPmQ51hlxAO6N+5vN4OgW9nr8x1GHrSmKG6eSVq7QroiCBxK51BqIes3Coa
PcNiO9vRbXTwXtdWzKd3FhMFjuKD3Aryp833U9TQxCBRg3uAzLHji5LB2Gsm
kUY8EnPnxSJteWlmiqyPnkPakFhRe8myrmONeuHZjsGX9Td7rQi3kMIGQ3KI
ZypzkyOkLXO4ppvGFO6nTYRhICL4cShZTeyrbQVszJjyKvs4fVKxc9g+aQU8
J+BoJSETKYr8qQLTgzLdhCF+kRb2AdrHbg1ShhJuvA1Y0fc36UPRIoPlo782
CFYJNuM72aZoGPi5gq3s/ui/mAusLLaUH/ZXnl1ESWRxepIeuTGmexpZA/vI
3zF7MzLI30Vf8KMzuVi+wHtjbVDCaD1REGnKw134NnZ5GewHh9sz8gqUN0wT
HoKeww1GxaDvW8PLBAVF2BwFFBJxIjoSGGtCSyytC/CIQsm47cCDZV6uj7p7
XdFwCVXaepmlNfy4FyCwNPmMR0GnyXgmo7Yan0l4x0U66p58A6Ggwa79dtDm
qz7hIg3+g+UVTTTWS7KysYa8ZDbXdkwiP2bxMyfZ2/G7+ocCDVMjIyBEaOb1
qJbn7y7rCWYWCWL3cX9zdHKTrgwuO/+k6bYKyXodsA7i/XVWO06sY6hlp2hN
LigJjSFZzwl9WJsuNdZXjFUA6nl6mq42CSMcOCdm1cU3aUbJsDIWXW7/m8Sn
1JwhxKGz+PJsml5+Zg5dH2sMp4Q3t5qk+bzcrItVnXmtQDbvzNI7XTLcYxpc
ahPsr5PxgYYc2bqf6teH124C/jtz1tqfT6js63QsSDe4K/Fu+EV/tgFRZNr5
IARMpSH+CP6+yujYHzwagSqFXgPG2Hy+nf7UcMxzsbM5MIPonnDCwn0g+hl0
CmBE5sBzw6Do4IRiaDcUEvaioqaMmLK6F8XVR1XOt2Tv6sUohhMgr3KBgyuC
hkvIxfPZQBMWooltiBnQ03cnL7Tvfng0FTsOMY/J1jm+qnn+CD7ZibX7ZO25
RtxpHeI9mRcoEdyW3c+6oPDuRcDqCzfH+3KrYukuWbBIGQ4awhpaW91gUpsa
lJLjEvdWbFjuwFw0zJqC9OQxRuVXr+IFtQqn4OQRDwfZKI+8v5+BBSDTRzLY
rYo7nXQ3jZ0vGhRwX+7VvvoX/RMAFP6e5R4BbeOjCy5QIoU8jaVJh/sg7WJX
MkHdnmfH9HyotmcpJ+okfIDGAS0mbP+Gsq89sHuv/FzOgOXfvMV9HbHTEEtL
3PCXnNZr5wYjM+uRR2lzp0cTfwOeov6RgZOkienD0iT9E99SUpsSuXnI/aiw
nXQEcJXV2bI8ZnNesFl9mJYv1KgfgGJsBYv4O+zR672HsMAJ0aOzma1XBMCc
UnJO+FKF3AUW8TNbKJoMPtle6/2ryoHgU9Kmlu8Iujch86GcbGOzHlIrcOBI
+0cnEON+a7Fkf1WaJAG39a3fwfprSuJRSB0tPwYMV789mMWTdJebqimmTIN9
MEev8jlyTAHUPbjTcnHUDPK0lK8JYNgiIPFbyFtAPYMsJx5QuPAtR6OmV22D
onaTB8SZ79YYqDNNLDw5IfMBJZ9bhI/CYwcVFUn8/PTx9XPuuQ+F+K4mBvdG
EZQk6EEj66HUdJBmaPJBKlw6XeRoUoxzkY4SbkfFOkC7mYLMZBshSA3WCHcf
u+obLJyairab8PKPK9qrdJw/CmL8MQScuNP3Xy8zaT8U190RqBk+4QE7DoxO
4I5TF6lW9TqibsU+5ceZfI2hvUTXSRHj3EwVOaDrT+/2C0z4XNokbz6KBWoE
dzPtmhdmAM3JLSbvx1wab3IP8t4t+xUYb6u+TOZkrwvJAuXiLlRkm5d3d0jK
R14dqFAz/cL2GAdiKk9jpDRQrKsqyceUKJXfsZU7ky4Cs87ZGFZ5QcjEYhOX
/MkLCnKG2CHIrUuWP2btXJYwDd8RH0fIIa4JnyUQ6uR3zRGJsN3ISy04995H
po3qxO1iIcZuOJIeP9CE/+dDbRuXJ4dDxmnxI9KymO8UixDPuGnCQq7oxOf5
TNDnsNr8oZCE7ncoSnhXIUQTKW1oC2yD6CmfWVFCRsb3A5JVvSF8EGNYjFzE
PReF+nTKsc1+tjhJFH5nx3m2F0wiqyUBboCllpn2iOb9+nonXMi5ic9Ep99Y
vCigNKTkySNuOWjbW38w+WGeJi6efXDI/vm9Ue1XlR9Wn9AfxtOsG6+cgCuf
/oQibd1ObkWQ/WgnewsvDmX3xXjYKUVKLrPiFyk0GE8aJZiJMAZjhsOVO5W/
C12JE4EWhn01laHs/T3MSwpPym0mN/jjI+oQE+/pBU3Sh9oGCPE48aEfVJ/Q
ou9ZDjSkFBcA++LbQB5jn06i6hxCbTHEna+i0zEZQnuiPQG6sEyHk0FHvHac
fptvYDXUx0RldfJfcDY9BMYkibd8OnK0lVUPVVkvzp3K9k1PdzWsj/Q70T9L
sAQOZMVlCeqg9hJSo7uSRpBaZP5c285LLk0uuk/GaxF+/IL7binYlTqZBLAJ
9BgaLQ7UIC96bbC1hI3gx9h6mxWTM3WPdcPLTLuHEwD/XW9NTjoEVGclHC6l
A+G4PP81Zdl0RRifiRBdeMXMW+8DTGnuexbbsr+u52ukuXocML2Tb+6Uvrfi
NkEkOxaG0xx3ruem5bMoXylG310UdXBrKEb8izDK3qQ5yJLSPeC98yQqu67v
sVyy7AU+jc6ww17jUjJ8ICqqLYq2qi7R97TZixIPh2ZNQV5aIIZT9Wtx6cET
uFpO3u97OSi4qCaebPQ5gHVMJ83XkgPhGKKZppn4U1TNupraoPBkUSMNEgtm
yJM19B/oPemtrqWAqAmGfQTORRRuJtGnoQJI+OXa1QBOPbNfKWhLVYdyzfE9
9kVD6hHrCWOE9510ZVDpeFZt4K7cvjrAj0k6xcfjpo2EBqgJ5q9a/JyuREDn
FvwnNdeaNt78KGz3OBOYdv3pq7MUtlCNfTVcLrrG7QsBrVGaXcqoiHvCAzpD
UJEt5FUHZzXUkFVXzb1B02V4FxosXgRRQ+0hDSlPWzH6N8WMvqu/u/Ngx/Lc
2/k/yxsNkKD0VujcMXjzGghpEyqwEqJ8DMkL5G/Q+8gMqYyNn5yDDSa7QIAR
4XH/pFsZlPjKuxx4abNZq5oplz9tR/Zc/HpJf2R5aCdZ1KFEQgPUSZQ6diJd
g+0YfFHRFXPZFnIvNgQG13tA9RGfE8q+uoNLC6xftDUbNPGSQRbTzUVZS57G
DyTVUttdXHWmivMiI/Wd81Gn8c4nussPuYUdt8RUZUOI/uRNk6C0Yuz0FEnH
pUUwQ1c9asYdX9uLjcozHP5/ANtiTLMn93WPPrSuDMUfe1IC9U9898vyRJOL
XseEnrqITutE9Y1epmAlW1WpcTXbPX8lT9/RTWdwaX4jMMqKabarDzCQgNFL
KWb1I+I6V6K504k6OPNu2YEqdyMoLBKFPtkDUB9/caV1i5X2d41rjfgZ8zwH
EhLcpb9bnPzlBkB/Wf2h2BWX0g/Yr5Kx/VHR8TpwOE9UOg+Hst+j+atgEG6i
MhwLcQGucbsbQ1+F8qtbMqMvAtJiADQgmzcZI28MG3tKB0/tmXGl4eMej580
FBg+W8Jivuv9J7FBKGAUbbkNtRUvmIO4Kx7yWabhx410A4oTmYAuap9NNhxJ
f8Teh8xtCN+6bXYKnPUiGQvtoy/7PL7dDS10d7vpPPH6mBDfMAQXv2/g2D3I
kcHcCFgbzjczQBQ3MqECP2u/HrCdcA87BkFM1OaE832xGKbCV8moEarT3cRA
4HR6v1qeW7vg1PGkt1VUnwVj4WW1FSjIUwfdOBju5ePmIKR8a0bfYdBnzCFZ
GRz/gtge/FHAbPQ8E2oe5hYv/B9AmoTbUxlHxoLBvql6KNBjBTtM4i4FqIEI
d+ui2EQnelu/yVwc5ImK6Hpdbinm6aJN5h+A0eBF0thgaGSvMNtJapU0y+8h
fWDRn3CLqVzYsYjY1ESYOuU9r4wIxi4B4tiOF4MrvcbNvHPjnmudPxWHEZFF
nWnHFoLSV0qim2eGERT8owkzLSv+aZlTqJUw+roz9fbtmmh3VPRhaw760ycn
PL4rcywkDhgzYqj58LtHOGLmeSoGNNVWSTbYc/p59M2hp/rkeKgQCw9Weiw/
kbVkV5GYZcKWp/278tSmHCG+3Km1JsvbdXHnBiWXkGoZ2y9g2tvC98lzqLzx
m54x2LvUggQQ/woVdUmZfXkxhsnSwTKzBycJgzwIRmrvC/7CPBwkwW2DpJjZ
P1Xd1fJqxPn5dsO6UC2qZTcwGGrLUl/W5gzD5dDrQ+NsuXtNODcRKAiHjLsc
rG1RAEH4Fg+Emq8yGIhjvpXK8jHKXGjgsIww9A056C3ppLtEgTq7/8fTW9vr
pOmLz/neAJzDS1S9inYvXlV0AsNjhXr1yKfdSx5RDAWffrXcVdQOs0VF1v4x
0CnxJ92qaF481D4uYXRO21qOEAXeckzg/GlCNOeVyDQ9+xhB/Mxz9CIpK8p7
1TazvjtoOD3aYCL3q4TDe8W0BVWyHNjuT5bIxZGWhAtLqwug/ftqmU/nMvLB
xZ3+n2NpGj7Lc6J5Hw3Y1nRR/YOzc40v40MW/u9jCG8XVZ3Dc9e8+KmXDYRq
o/hjVGRS2yoKSaA1yJGXZ6ww99ckN7dS0WZ+V52VTSsUQC6BXP3lZiHdV60B
+HIOFr1+VH/LV3T/d3Ly3QfgoTjKKeEUI2lUTF7LJdW8SPC9xNxwXmvLtDDQ
nZwAORipC2L60BYMQLOkPLMdQAwmdagRrHyR6IRF9lgK0CCZQrL6Mro/1Plq
s8JDL5TVnBEffVU5PnevuJ79+o50RBdRCoiav9SasiftGT5+dWTOE46WM/7t
2ioz8CVRvSVbyK6ciAVn6eRteT2tB0yvXMyPTTS68vkr+sjaRcXAhhcjssyw
AtQWuOL0e3Ne5XnqS3MKPR7nusWZdRiwug+Afm+AF2uOL5tkRVF2Vj99H3du
L5u9PtAp5FhAKflbSlRppYf5B2JUf47IFceO3tBFQhZXRegNS8Sx/TSd1Vxd
7MFOkmiD18CNkpVsvOBWk6nGnXg4uflhrSROrKjQg2rhqXnXxBOoQh5Qo7RB
I+SlDZFhftyCkCoi9jxKmUrfMarklGnQnWMHmwVmCScyCezIkWrwGp1vQyO6
qukgkdovYirQtQLLIl8j6kjg4KVP8rYo6vuNdrDaNmE2CA6Hkj505SqN8Gi7
PN6FKAbgcFxUxETxg6/GV9Uqs71codL5+v/wxnixzy/D5S9J04BLj3imFAcv
sDn8lM8HZ3rNm35GMdU94qlJsf9ZAnzaG1fcD3JTJmONdQVSSGL4iTm0y9bZ
A4z90y7HlQPlbSME0bKqk6YZyJyFJl/xTjW4O0MZAcHS+kI9UE1HXH6hO18Q
o1tEj7QvSinN0ob4Ew8iT7WC8wDFgqrcNRlxAKqEl29QL7oDgPDxUL4505qO
aBifvbIVrClPEN8n6OcUrFT44QuWcxe6qhJ0oMW5J9hw2rJ/bJaD/r2cARND
3krtULAvZ0L5EhXnUxQNJ+se8WK1/110JkRajjGjS4pNwigZha3MmKNev/qK
dox5xTHAJeIxIPEabttDDZyuzK2eYljNxkJcDtQi8wU2ioDAxuTyruvZ9f4/
uL2HyRd/RJm5avHBUIqoWn6GM1wQoMium6nZ74nMhvyscF2d08+7QmhyHusr
mphJdOOQrEpFJVzu7PUwg38XqENoFCzQWGGm+f1ufxQ63iHiJVWqA1Gw2J4Z
c4+y70HXMo4g+ltPZU6aHoWVJj4Y8uKBQ5by3vL6uJBW7qyNMeuHpJzvekxe
1qSmkOmMlmWy2LXH5+Htvqskp5kHbIdWE+pN/8/UK+fiETPLNbOWaaJ1jnyx
JRPNamWCV2k4OFsjjQa+Iq9XG5UCz0SdZp/Okbxe8++PG358gVh9eRxkFOME
SCT/c/BSSUsOn2o0GMF40Iln2t8xzlX1ANu/LAvAq5nnnlqV2TUnR9JNlOE3
YrY7p8gZ2lOdu+44KKcjWr9ol1EfIDA7OCkOjk1j+CHQlSUQEqUBvkT6fFWg
EGNEo6QA1QZMRvlote+ygb/PUkXnQBXNhG/Lp/gHwPXyTYTyqJh3YOD/1lcM
PAyvBpK6S7IcTSJX28hDTkRyLnKBloN6dwOynREcJbErHZ+elMuMK7G9QTAB
WX6LMkRaWkeAfs5VBO3dZGYAIhnHpX65n14kd6lKcrm6EuijvixnFq1B/zKo
6m3gkX6T7bihkUaSW8jQPKe6SVYGtrMT/0tNMsD3QCaUHqQi2QMZ9rVq7gIj
R06GLksjnJyN1Icq585k+4R0fVm0265IsFStgSgmkOpHkEdgXgh4jNCfvVAL
B4MhLr5iQxtcwC9zcQMO32FW8OtPd3ubBVHw+Pb7tJRM9whZQBd1BQqj3WVQ
0ZWX4n0d53cPaeI3qq9WilvK1/+bysZ5Qt1+hlmIungTs04+ynXO2MGUE6cg
U3Y5X+K8xidZQ7SL2dvxPGsQ7wkL+Ga6Uasr1pAPuF/AB3xYuxnAsv/MnqEU
1mWAwL9rV9dQsoRgvGbDTyxGipMNrlofidcu+obJ05kL0bAu23JmW38F8kZU
PIH7YWaat3Sl+GEaZOmYAC8HQ6FJDQ1/W1uo9OgiYSuV/JQh2Mh3be/k8QLR
BKxFxnLVM7WWg8vH6K741A4Ipi7HalNwG0v26UuyjZu/HsLh+cBcADOIE4za
r8LacqX8B+ktXQhpsaPvoVFT8algc1WnnOVHBF3JveeFks6C34D3vOlOzGCZ
e2MaPKFw+ozNMRuPAgwEtvrWiSwTAivhxPIkpsKqcl4ogDYLTt0yrVZXmP+6
WM2hCqhe7MaThUDVJlytIsvxB1v6yYGHCVy45ULBCk5BCJjFHgOOgUGorZY2
4eesFn55mns0BZJazymv3YWDUUzT1ACLtA3UYN0bvjc00XpUst0GwuM2wPnv
d8EM5hfqNdNWMxalqe+eV+yPeoZcUAj3FzMhkgOZHCC+36xQejxv5munjxHG
EjOiAnOf8rT43cIKEtwePa/IkuX1iD04T/yS3cLBb5KU2urzmDsNse8K4mu9
gcvY1tOMOZ5HgnuRF7X8sM0NNf5xB0t0u6nCNKnXwwN0yz0hg4x/e/Ob+M1K
SX/avOtuch5j09TvVwDaxAzHD7E3uFprZRO5NczLWzWpwtGLtw46YcQzQ0Hg
GjgVweHKzgrQ+KEb8N01hQmFrlgJZpNyy4cZ/2MFUQvzEaxNoq+uOdz2xn2E
BPAYnA/5IsW4pQ7QLCuXPVrRzvPaXyOHLAZDtkl5bvh3T/cIcr3tmwfvpwzw
5m1HTnXvG8SColOGX/UaMEE/d4mhdCtbOTtnuVVHG6Oxm6zDLzXgsJvIOoLb
X867WbP/HMMD+ihaNCBUNOkisjerd5YUxeQ80oGZi78qLxcR+l91UKlTHJNs
UlJRr3L7nshhTOk653fACmTMFtLpPHCk7Cvtwv33HVEVrTms3nOKofXGFPzf
lV2ELPc7lM+c+lABZwKK0fB8Udt5P+5f9WVIJCo2NeFWXcVnJKe8N4KWQnY2
WPLFMxHFbTzXV7O+i9qIHnlnybMe7XrYNCfokzzmknDPz6yjTooyZWsNJWsx
Ai4FesNclFhuYZ2GM92lPubGniZjx74HwbBEOwHlXPD9RyXTYDyqJLQynWR0
hmiX2VHNTS/jA/Z5H2uN+lIQg1PTIG2Eh/OGq+aRiZklIZqwdFfSRzvOO39p
N35e7wNZw8KX5QyTvsuVtp8zBhQE4dEukGE/4JzXlUBX/Qt5AaUTIC8H3Czs
J9B3F+WvGXU/hY/WJV4QhETDZrg0QCIdv9+PH2E2i9ej8glMX9cLu7zjitGS
v7l54zzcsE2UVbkhlpaQdx9yy2i+UMbztCLwEAux2uX39a5zFqyO8A1ASS8g
cvEVw8e0jFSge0+RoacOKg9gz/ePweKZ1qqCB3dvRzqGHsMCOjCzodwgLk0d
UVd0oW4FvZ0MsA6YUs/Hl03zvBRoBPTaHv/y29PtNCIjZz5qKLSPKLDUTvUp
S6ITASOGPy7Nyd3Ws6MgdrsCEHnMRzBkyxUuDkPtTfd7UUidbzRpc1up67f7
I+x/FxglUF6K/22sCqA1UX3Oh68qamgDCoO3cG6amLuXMbjpUXIIHg63Z9sZ
zjkOFtzndv9tcnBanzOWc7v3ar5IgLgHwEGw7BKEHp8nYfWWEWgwp/eQy3Uf
VHzj5oFwsyplTFXtJHjfV1fHc3eQHAHQ7/mNNLyrCzyPeNlAbh2fLX3dKtqT
yxMn77e7tTY0tPaSmDdGnqS7nSRTx4V9kPmQOtZx9OyF9LlBJOwbbUAB0lXZ
lxnLFCj9nyijQqG1ircfIcDm8n/Nah8Z7LuD2nmY4EC4vyCA15beVFvThZkd
q2zxyAfEN7MxW10e8z1tzmSfCRhXTPFA/6Rs7+Ervyq4d+7xrfSWIYCsNBva
OlEttNlR6Ze+xyy0zaORWPd+WIaQKF6KCU4uuMuJI3RW/LsETJ9oJLzIrS+e
xwhKjcPMo7sfUN3NOxTmue5gZXdnBB+wyzsOT7/LsNP3WWO9tcuRql2NQRwj
mgpJsXbyG7D59KaxrxfCucg1YwE5YmicvpSvXsyUen48R+ZRwTOftN2ot3+I
uDh401JWmNr6MwRvbZ9F1URwpy734lW+MC17XrahSK8/jhsHrQO2RmXC+yca
Dr8cWeMfQ/ac9IYFPOpw4J1nF6Rmk+SZ17bxd/WKK3E4pPatdMDiyPj9geJU
EwfmyrRjfPhcg5vu23rppKnF8pTXJFGKhhYQtFujLUGzvmjyID5sYUNUJOZ/
vqXXqDiitGXN32uwGeU8y7qTCLRfII3yF89qj0WN/acJiGseCQznnAOPe3zZ
op8HdrNzFSwZJfLxMGuWEGBGt3HYiubAOyPpBl1ZZ0NkEEULG36oCrXVTfNa
jHoSOITwEAGExlNNb0TD7SbhBAr0AzuO7TngUM22VxM5rwxnNo5djhOJR6qj
vzDUmEQeqRH+Do0D9YjtQv+IXG1i07gfqEgdltAMiPJOBDmZ9OU/zgyurMLG
Y8bzJD2joj4oKlwSxQRfrTriXs8/+2+4L7QkC3ew4S9OelyD8zjQWrKQ3+kZ
hOErg6N3k9CXPhxpuoqgiq+XQS4vCLIEjOl75ExsQJMSS8zFEZ0SRhl7kxlx
G+eCS3g2FIsfNrlQxNdVILi3Y3+DTNNZcPwVxTQbrb40xQGrxzUtTDVBvE3O
w/rwRlew4UsWejZckN+ftH6z7JqhB1K7Bw33qOcx30I3D4GKq5KNzRLQDuVp
6F//yC9AozE30/RmhUE+z9EyU0Ws/aobibXYnWUZVAYX5u2/ny7E1sbwQRiL
zIYSRpm17vvq0i6S15+b4WXE7ANf8CkyBC4eiTuwcLMuKtDLM5+vegzZgsN1
PyzvbwgUztf4UubDBpHG4N/Q+qRBje3Ij8smOUEjuxV+L7155CrqsS8z4Znu
zZQplYM3EVybZBQ9OepKLgo+tmZAsT/kYw9PfJfTKeXRVF/SLVTUkPtnvP8Q
XmMCW3G17kXL4GDgmnGgCih/uOdpwK5Wn+vcI9Zng2ZSnlyMYZGRrMDZlt3N
7Acy/Pqzzw1DILw2WSoIM0FK6x+BzjYMDDXwugn4MoBRvkhLajwBHPONprph
dQtn/PUcqnKudUEkVMUsVe8Uq0zXRyxbBQO2kXBNZVgO6fC7NewjZiiVRAQO
5JYJwLLKy7dQpGshqFZwVw+SDW6lP+1XXeR70kMyyK7Ml/kI51c+LUUIA0+M
6HOTCqorOhDIdA6TZWgWRPcRe64Yy2hfR/4CKf8+I/vpiex42SAbzsMLMuWC
6SWIkSeuw8iSXwlm7nRDiEwCrsRiUxG7W0G1omN3yUjufrumW/ZnldO32EKA
l+15ev8QoxY9uXMjWtYMtUO/xdH3B05vPACMy99Duh0+uGS2qaxKRw4/Clkr
ejKjCr8dh19xxCpsNlIHkAAw6Ydslg94gbySUZGiumvx73vFXhhvUUap9Q/C
y2EKlgjCICpHpb81cUm4q8LOuiVmbYAS1GBZHIoMoIB8w9rpOqgvC5ioANMh
W3GS37Ot+q/LEuLqH7O2EfpkgUfS2pgpOtRaEik8HaL9D6CdZ79Yy/LTE7uj
0OkByxfJd48w5WKVXkP4R9PNlWHxzN+1BunLo4Amk/5ZAzWkb3N6M+79p3CV
mwx7KwCaktRHdbU4bSe9hXUjS4NI978IJkpyeAfzcEyQQS4m7obT4ikhvjUe
xEFjCBoPyPLzwjkOu64Nk6X3qi9B7rhIFXgMg09xEELCrGCfpMpsj+U9Prjv
GB+3RPNqf42K/QSB0wKJyu5R5YiLOHfMAAcuHR43ybdTfZ2bN3NORihyxQrW
ubqyEQ8+qIodMNbtLogN0fo+w4b+D1ANeSumG7wN3tGhuBBgLKAFxN1epoQb
X+64n8Ov9uvUNCuh5LUkYccINTB/7Tp6ehO+91kgM+rtEOrlWCwRsU/rWocW
rcmd0tL61h/S9Z+mRwstNFELaT3Vuzy0P00errj41CJa4LORN99P4CqddU6q
0ha7P/DWgW7x9Scq0uQBECnBMqD15kdt4en8vF/qWiFmuQvRzVe0j6zt6HVJ
xH5CzjXoFoDZbFEyxnEtZpcz4s3i3cXqCVrFhR3PVy6xjz5oDlrPSQ2xg6tU
gBoAOtLZuzGHHrXGU8YnbiPQy1Ixv7EjJQNZM9NMP+p9IPzrzvXQNK+F9kLt
u+ueKSk+P0H4c093GgczTt7qAqbajSzA6txzgBSKyfr4IKBDQA8/J1d56g/F
NLIsFB/aUWMCy5d6miUSUTX4Ys2MDRjVD/cmTawRzR1QxPRRjOhLfqFszScN
sAc2M7DxMBkdLLo1G092d5QnHpPGldzZ7H9YIFtERK+EuN4hwsswME2dSdeF
UqZY172/1DWB0aGL7+su5ngeuElhHEARP9Bg2SpEulAsr5X9uOM4Zn1T1z2w
8R+yVHERxNThZWc9GkguwvQ6U9N/+x+Tw8NpuAplh8M7SpEpAIh3qAq12rrK
b8oa8YQb37z39DLCQoggCoybijSfGemcxLTTVdeg0PScvgEFhLnBgCOUY9Ke
pl1OytjPk/wF/2ROL/RCKIlS+XFk22EGgrz9/VPLKe9RA3cF0Y/KC/t/WAhn
Ty4cR/BVfjI4RI/koBfmbPaHdudT0x4hxABwXURoPdCc6ugyXf1M+XfTA+AU
pwYsw6WiXIVhJ4cMiCc443AFuy7ynCJ1PK5RjTmw0iio/iBSveShkDhlN8d2
2PTlff2q+DWn73VxK/kV+rxjVIbcRfSSiU+6kxSDOdJko/lfcT8nXl7Yy4LC
iQEK/3PlLf0SzqS4UsnJJdESJz7ColYfuAk/6JRyyRV5FRb9y+6V1HPMyeUQ
dN24Ocwae6OLP49ePPRqOoc8ecORt99p5a7hajgVgSWVLilOPpjivq9dQiKr
2t18j5M04pmXbnCaKbjIEn680QjimmoQscad9TTfyw8YmpEsmx056WuMrgzV
LeEGiODK3IzKNQ7PZnZsjv58RZFjwxxOYyc+JWDWSOuUElsmyt50tp1iVEzN
RYKoosxcp19K3tos7BCPpfwGP1vhm1chHhkhnVj81UAv+BDmLrhAltmwZjSJ
B04vgW6bfqqQkUvm4DIDWG4F2UVbLwCXOnEQNNoho4s1fGocvtnIhOLwayOR
6VuGi2RIVsMa30m+bavvttIINTyijRVhVwzc2xnwyjfveDBGSO5Tb/Q8/HBn
wj8aewidks/y5AtL/E6+heRQ1RQOls3rP3VUwsGVR1Mu3y6jNETqX4s3alqA
c4ZqcCsO2hW/+EjEzJ5S+FOMeXdeysJfXI2FhNW3zpPwAShnwWcivxeFEMEV
uuo+EC4SAPvpa/xg9uihUA8N/7mJ0lM6UMHJhjSnwUWEUcCCsJE0W/m6zTHu
eRWshwCrx1NwQT7UwQY7oFU9WjJsSfbymzz3RrQCpL38gNRWdIgAnIcETTAP
TvJGAWKYSshJrzbR5ZCVLT5wIQI5ZEjD6XnjjhlbBXT5kRt2ALEi+zyXCekr
HaZR2bjPjzXimCX4wrvYvoLaX3Vxel5OSBf4fXWDLBURKeolNL7L1Ptx5Jcw
4uAemBhgpdR1edqBA7qhCpyecgi4PwjqzNGCJZZHxsZGwB3eE1sCfJiIdmfb
jo12DSnIi/e56+VL8TrkXm5+5QA4e4PWgU1EW7LHyhfgWFJpTq8LigldmDLI
y+FDrxLk/eP3hNR/pQDnxTDgSglI3EIIIbcyCnaxAkL4ZlY36BsZPGvNzK83
4l7AeYcbf5dmIEw4AzjMXMHzzmluMXvxwLteEHvXHmJ5sZcO/SrqBLpfwqwR
V/KlcMN463gY+7jtUp9YHIFeBjX+/N4AImlFSiVx5oRPE5pWpZP1cvojS2BM
o0qm5syQVPgsnfsvZtgf79XRDGAgYWnWTed19ckmwTJZfSqmHSUzwnssrfUv
IfFY0/pOrYFsXPU0PeThMJpFUtjeglznxK8Ceq7kONvGXHzSm1ps85dkqJ0j
X4NA52taUD+9hMGNOwAvOBVNDGW+uKnw52K14VfcEpiczyCZtBGfJd79Mdxm
f7x5wDUaRJWjN9RP6xQ3Md6X8DN7vYLdUDzBW3SqiqLgLfzRSuzVz8wE2Stv
qwg3njb5xlqBfM62I9NdVuG12RpU2zwAjJO4swLhWe+HDm69aNUfaKBJT0fP
JfVmDFRHgv/196wa3hLLzwHfy9WcCzcFkuKJCUA5oogP5SGx5+KL0wJSq8/f
Pwqvd48fJbpAlz2WGw7n1AYaCo1UBQMfNTcamgQENiV5dJ+qm1sCBoeIU9sP
iWpmAFHTti9Y6WqnJzK+AAfYUDGVnpCMKAwE9quQ+0+3STMlKJvr2nGRE+gh
qEk0AyUfW5ivnRdrEUeUP3/Qx1hlFTIrNoZU9FTokMQqv2JB9ze4rAWQTUm3
y+DwXCRiQbqdptzH3sX7epDmFM6s/hfm782ObC7ipon3Bs7gNSphwKsoRBRC
FYL/eDNb9sRYOpJBFlXyd2is3iSpaFMmn0VsSirSUGAiMq+lVkZHLqXdExXn
z7YFeYfssjL4rmfTJHv5sn9zzu3Q5yKVUCgYni3d+axAZjhbJwPCVe1Xmap1
UZzawx50pmABDsWZTTJaTs/diRMRUAu2a2lagG6QtaioccL8ZenVSVFc2/LY
Z8wU8STEFNLQDncrzrpN6hb29zRkaXoDFWFVT2nyFTErJFQaw+FZgZGRX9YA
EbfsPNG6NCiQSLwpR605X/WTtujSZB4eCJg4cay6h+H/28ea4wFztUl48JR2
/X4FHJ04hHOBMZoQzeYXXerW0OaFmZ7ZZH0YHzYXSb5WnnDRAGZ5DuOkxYf3
rrab/4TCFwQ92eWOtWyoC6imC+ZUWryiYoYH2kS2ASfMiqTxLaeL4dmjVpMm
vlEp7/DON2Z1Bwnpe4gEEEItpRHX1jvYpMtgHI/BJGiMnGBQaP0zpExNIm/i
yE2H7zWdYX8dY+D3pDEtngHsL1t1w3iLikbwZ1/z4WZ7xhU2M8ZbM27SZ7nl
0ZnWZn5tVMgVP3k5gTofdEAUpS3yWPnWCNkRGAz3QMapBKXGS6N2VMo1tzoE
KhwfVBvSvvAhdVuiZzzjmf6wYt739+8ImPyZz4B4OXJsIcoCGZkCTEv1u5Sb
O3zLbFtIQ8uB87/m7lTv5pb728hTteTP9XemoKBmyl0pPzCT2dksyBvn3HbJ
HqtnuNDFcctkQe6xuyrVDE+gBWBA/eOS9yleYO35NrydFDiZu5qD2aXLZnOf
B+YloU3J3HjzXZ/6cMLh6yWmoAfNeaTb8vxI/kXU2zm8hTMNuFrf5XYSajae
eutsmun8oMu9UdYJnh6ZSY/Msj3i0TOi/HPwis1PblTelXM/N4JcThm3vAvZ
AT0TJWwAYQ3vSuh84fmVKsAVap6DsdDav0nFTOvSr2kTFaeNfBBsvWz7bnVh
SUisxG24wmtFy7chauzP52jcQkwgNsiqJ9DbYfKHE+3D8hyKQmMGPvlO21d+
nYpSgz+S4Dc/7jEsmvzZk4W+yYu6KiOmnlt8EAaf8GqBsUbAYTFFjZwOrwIt
TNsJzgv65lMd4dUAqMbcYc8fwAGSkUIhCJ4yEoCcOi4YvXmOuMmMTQ2Clt3C
ys/JOCqha/a0ayGhdk6T/YHbzXvju5ArSDBpgr5pKtWIy68p+x5JG9dKtOqw
SsLKpy6vp0gUw/VrifHmyhkjb7BUXs/vz8cUzUIxqyKiQhhw0x+B+RKTrA6q
960lGR8Aqb2O2S/OV4stJJHgu1VeNvkcFBmaVZTxwsW/prGIhsoGvYuSigab
t5jUUrEncz9rG0PH/ZfTRjd0WXC6eIp8fpRKgucpprZVdSpyHSkQ5Ow3D2lx
QKI++dwbp28oU7Lka6ot4avlIIWi6iqbZk/bVTUTj0yjNgt5OdYTCfIFXL5f
cDIB6Ym8HmWWCipienb0ou5Xk/RFdTOx4rMVBuUzZ0wwghHk8YDnIyF0Yvsd
NVF0ksVoO8FcI1Jb27m3npXCUWRmp5MFUKaJl14ok2LrN6Mbb5RCChU9/nig
Bzocz0HJBjVS2ZigBg6gz2sZsQyoG92WL6/97F+mu3q5tG8dtCEaGDel9+aS
vb5HtO7hjk8SPVwbgpBGJQzss8BQ7XJRd3fsKRrnIERjjPqmoHwGVvDR5GKp
4dr2aWmtdehGHtRv/BMpQwFZgpnkUc41qpaqq7sh7Sozgcbs9x/ggnmnizdo
mH94jbxaLP4roP1Jc6ut9YqC1yAEBnOMOoM57T+535AU9NWtXV4MTrLjGblO
oWekr+28waR7/ZcJSkP8O8IGzmugIGQOCynnH1Bnet6nEWnDjdCiSZi/P+7D
B/egrf2zn+WwBeWv8cjWCGN6LnPRXOm82KM3qOHzZw6Zojt37TI6pqAXaS7j
6ZgUCT+nkBsbWEs+biPrI1LoVc7ynImpr7ELIvfv6L9QcqSFfAbQYl5iSOki
cXH6r41HcaGV7ZzTdN8oeVmZv+qNRI2gMP1dQWn48z+YvdQTSIv4TX7lBrYs
0VQJyWb9anlKR2FlsT5Ck6ITNi/R/SHK9M+4yQeLNOUZxrzBjjtfP68K4QwI
OyaV4f9OcebK5Y+rQTIGKC6McGUrZCSSuoSa2sNDbufrlioq1+mHMwQ29UtC
GqbwNC2zVLh/RmfNuLi4LU+w4rm82wW8X6ToMpbZUmE5wuAz95kawnwMPJxl
Fr/8/hxu7kPOeIX5BhrXqr020jgnFXr6+rjfuRpkB7exZMJsjIpY1mYrhvTm
qxhzQmKC8FZOFImSPnhpcqNMXn4n4d8nQr2Ltd5d5XSFaXqltloFHVIu/Wcp
XmoqtO0BDqJ+bbnKVF3xqnTu1D2UZqvDNt/qUn9GhxdzC9ZPIajMJnqmLuuh
ALh2jonZKEu4TYpJ9i/x62dznADM2K8T5IPt2p8U1tXQlRjU/31/a/hl0Pdf
KkL28zlC+uCmvjKCXWnEzy1RyxBNKusqibPqwqi6XopupONvQPsxwROxr6/s
ZKOfhmaLXKZHfNLJ7Np0S2MgBr4SPONnfhZd0PqDN9FhZJK/JKhdxDp1uz22
ZqLX0ooMnSAeLeIgsYllNpXZsJdbTui4gnGN7vrk6fo797KT/32tE6b0pg0G
wzg3H58fPswIbWF7pf7wDUghT25vY4K1OLntj+ga6VdROds5t1UTjSaUwjiD
N+pDJqAdDSd7r9CggEQDfsONkNAw5HH6Q5j/cliwYj73iDMw8ehLT3EJYyC+
prlSHyPJjPsJMenuHES+bZha/QDHGdY+FFO0m49+rXDVpK0B8SRHw995rrdz
gaL0c9xQXBYdaVEUMzjvrLHr2Rrq73UBInBxouORwwpdQSyc2npkQxAuzeVN
EF++AEK36SY8sujMmKrx0JSRyZXxf61o3v4/UtRRi8FidutU3CUhOJb5+2Ms
1u3MfsLWz60tUMrB8FUmD+5NMzLpWLtKJAgpaEaJ5aCYpw0k13aSTy2aczy0
Fx3tRlSCzVdqTKFrSjF8EKkcAj0JslYsKPCyd8egY5W+BUsFIQF8x8eRthXf
ZRZusVLJBlA9SGQwf8jvUOzm7jNuW1xxc5n0R066sYvyawfyjI94n60aOOAD
rEnZv/CBvN5lHdByxo/IOIZHdNhBtPNltajhexmVhUm+KumTzJfVZuVT89wp
bJoCCldfkuGbFJ9fHmy60QdATkwRXQ05hqXWeZCY09pbYhtjFFf5r1lnjrf/
NaIbmx32rY3TucxDzy3c9aKfm9Op2+HPcATsxE3G846GJODZluE/4LSH1Dwy
FK6y133JLoHXVRq5leK/1As/T8g4tp99M6lZp76tNjnKYH6437nvePwisLer
XMcupGBLP42geN0O+Fdz29WlaSP7LYwk0jzZFdgomXZV/XJS5SS/W7ao5Dlr
TG1Nr+QV9RtJBanHSm6wjB3bi/fl3bZUverifKVX9YvGPHnwPIkengf4UeHt
VQFqMoGUfBquvkR2RhUc9XipXsxfDzxYorJIGEqHBFxnHRurWW3tyOUgcLf+
VJsNSzH94bUPxXz2G+ibc40AJWPZzDCWQBLN+lh1q+8Zvnh4EEQydnp6MRgT
YzbQH+VoC9uPjeB4s687pNCJnbFZyrywhfJ4ukZPNyNLk2D4c0UTyvrBtZzf
S9H5uCppC2Ml+7XxPJ62gvZvdVy5yVw+XLNKBsc880dkX/cHuU4BnHOZpSpG
KSSAzNKHFAWMSOzb4l3gg4jHjoDIxlka5W+cRJsOIVZoemmb4nHHDJzg9WUs
xOp1Nv7/CoWnCDpS9BvkldhL4NSjmoZYbVcGxsR7H1Pr6a39R//SQWNrrrxY
SnQXVEAVCqfk3lS8ew0SNS4FKFXicb6O0TOYm+u7UUZx27d+gAT2xe2xEy+v
/nTHTy1TrIKxbGaeHWqsW0Uwf5Re6zH1k43NSS/6FCBz71IgicWwLKlGzATi
QtVIn31YVPeAbmSKh7a7cgcPpi5fmeQkbnfsZyR4EwKhUnRCCYqdvKS6ES7Q
fwmCyU7QfuWEWrMbL8R1ZyZLpiE3t3QXzT4b97ahGtjtAMgbQdmNN/w0uEbc
Rd0jWXjEx5pv4OJzMWhhcd9Jza4j+gEiLI6qLiJnw7bc/CoY5X8nDypl/0NG
oNpKs4jJr5Yv8ZeKBJapJTuLuz+Jhugh+5FGvD2iLvMsxzezJVvgLbEoqho5
jhdPkQ9nRPHahGM72IaQSaSjFVLMrnTCHIL9bY0+1xqvxbFgZxV6lxmRcWIn
iGdNvOdjMRYgQOkFrQ5Um5Cjqpc/dymsfbXUVHINkBaN335p/Eyuv1VCsWq1
ReKjYleGps29t3hLwgq56sqJ8Ks3OcehCpGKEqh1U7MkUSvhVGr1rTnwS22Q
1wptKnVlz+1aT/EF0Ys+9vQ3KKARma3ERUcTous28THIQJ0QRjwMVKNhnCiT
ihKdDO+GNmrvP8tnv06leB0n2S0p6YGz3F0ugOTw1OiZwH0fInyRHqcsEII/
XtbUTRxHMIVMtkbU8jkLsMXu6jcRvjB86LQOINaVjijcaXoT8rP8NzONC6/C
Vt2CPzJTloVjslq0+2tgrz+6QQbETRPO5U1iFATItnVoOqRgNwbgHUTG8+tN
o1pno4tnnDyPpVH9ntMr95EUekcQ+/Qxjj5SZQBUibv0UzEqdCJ/SXdVHm2M
Lq072j1YJuXR2ql7A2qLlj2WyfLB2KnEmQLdqDjv6nQYRJpAVNEfhbvQSTSr
g9o+2FAekLtWdqzh0SBlrzw1CLPyZhQFrn4pseabnOkIvPyWRHkyqrWHJcjr
R4mbLCTqSmZGMHDyYeEGRTs9l7rhUp29jKl+OipmimXJyceMi/tQTvt7U00D
w99nxqlfTa+cjq8ktH6Ak/DcXFxOci31EA2f2FoNWnvp2fgZzmKWlYEc6pWN
rMNUZ4rYA4/0qHsOnXgasILdNXHiA7a5L8VMBO+eqJQAI3NgxGURlLSSkFY0
MsFsgKVrZMJd/WtGH0CfDAhOCOuveUHWCUiZVkeSR/aSdfT/xCwjVbxL9W1P
V3/306HQH7sLZ4QRJSjGAgDeHIUgml8oaGK6FpjrVRWlcYvj3jhl97DOFmgM
Z8RkP7OEejdakKws1it8Efluu2lTRcMyzQlzVfLJJEA4+ej+4KA8AYmTUn8D
ZIXuzoBQXSOu6QZGbzPXotXd3GRIXRdlQj9BlgZjlvojGLOIc7sreJCVmiK4
dXGe7mMwX7TqTEgtCPub0P6rWyN7iwxYMezUHBE3wB++0NZtoWbxu0I61/s9
36rS/ZD/0Ddrujn0+WWvI8CFrhpehvnICExLnvjh99RE+Qk+Zyi9HeCvEL8U
m3bo3XK2ZwNE6V56XFPcSrHEAsZKEDrb3q8PjvUt2HTIDNx411jRu8PvP1s4
MMYsKnkJTPURKVNRYcz9vz4PjNqDt7Slf5cjKUzOxi+5GeZVwNsmBhzUCCfn
CQs8Zqeek4IiywJjV3ilnI3YpKAUoKAc4mhCOaRk3BC8TlCq4F4fa34Xjnnw
Do9hs312e3Lgc7KGZMDHp5aBgmzuvWiMdnGheej+3YZIPh/VJ730B4yXV2Fw
NV8nrQaJ9i10JO1xSFG3iM1J6IoqbOZTUd+MtYJokolaHXZFI9MRRb6WoFCG
UT9t6QOs9+T985C0ExGSLHIQ6u+gxR/IvOTmgA8fce51z8ziBTMMsFndkvg0
TEhoAhJ/FzslcMljVGrUf9hkCss1h8EUOAgKNeQlusOv2QREFKexzbjGtsUL
fk7lSAAF/GbevABNoR1ov5+cMeSefoT/irhBtHJRFFb9QW13136wURcTS7Pg
i+mCss+lA9d5iiNa5TWxrnO+QMg4iiv/KcYyX6wtM6WMtlotRcefT+1WxDkd
j82W7CV6lVv8PAxU+e5X1Nmk8HkGuU7MuijhIz13EXkxJGHp5BKF0BbXDbAb
ruof/iRXOhr9MnTuvoNfYPnTQPw/zss3/zONBaBujXz2xvym6hdRA5yRRWG1
st5Cd48HoBq5h1LjKFv42FBE1Wma9yGxDsJ0NOg5zE/iGkZqdFD6ZZUP7JX2
LgFvBiJ1IYkMy0XPKPQ7Mp0LBusBBtXVjwo1jMWBu4TAXHghCviOGUb4YFoA
DKoka8S4gIUepvb/c2m9zWmSeg+LwOMHVlVVamngAZM7nn+L+xOwcjRuzNst
1mUM+R0AC2jZCxOF0WlkJ4KrPvHi5ZKzkwzN4vrzimsPVlELGyrDG/4Cebos
qeiFxphf8KzvY1J+9xdH+bj0xXUs27G+g/MAahpdU9pMyrc6FEXiXEyYJxpz
utoR4HccJd4SjEe+J4yFUET6sE7Z0BU9vDnoeNlJbFzqGGb077Txre/3iT9n
jTEyucTnhqnKL6rtnyvP9h7cL4Jgx/08qkvIeOA0Wo7t8y6xJ7gPHtOsja8/
4e0UcLVl+2uTnFRxlj9kn8EhpeGuYqRK7P21Y5wwB/AGHfLGQ7iUp0wwwjg2
/Ch3xiFbRO5iNlZcJZMYveimLjLyHU/aSKzRzQnKt8CEFpw/lCegoMTvgl20
Twieqb4AGf19zsK1bmWOO6RYYrU7FL360ItTDyljUFBNOojLlo0XQ6ikjjnZ
sWlyL4QGiyghuN0VPmVHA6ac3e8pD1hjaDEXGD7sVgsAAuZMnvm1UWlLMMW8
ZiUD6UqSl+TNU8w64dIa8ti0ohi6oPXn5r/P6KjF0gvhz9ISrpYh1l9DQkHa
p386VupV3crGZ7nkjwA1ZRAMGWcPZyqHBX45VkeatwEBllwEbxPZ5oXI6RHJ
Hwi2NN5euNSNdKwQtAYyXz/8hYfdTaBPxHYWGyNBRE3fN2gMo9GMjETxNgz0
kPEsJaox45/9BLj+QM/bHnF+XSx7UdOwCZ5quaIuAkYG0mb2Fi9JJXiCtNhg
8Vx0N5T14dYEsy8vVqx/uhxeazBcj5IIGKJLMjeriY9x0TDnieQ0WBGuyAJF
whTmlsjZUD85zNSrM1T6U3ouLaODU3vDbTp9M99RB/0pdmO8UizAFz8yZO+z
kwqYLrAZfqFeG5KRGgcdQVysrR6QDVEuXj9X7o4hXBUd5dKN1fbv8zCCzhRs
qz0FbKIZCRQ92DVgT3OoWoMWQpeuKH7X5IHqIhjXI8mBT8/YUlFnhWS0p+Jg
sku82D/rSwmuyenNEauINWnZzZDkIv1rrxKX2LwzvqtP51wYPsDbr3xX2n4Z
tAVvqAVfA4qzTFeXT4n5cv9XWvsh91FilC0W1eebKBTNtbOJQ2d+zJegUnjm
0hxrg63Rr6C+eZcmwB8ByQoBcZhcmR+qtTLPH1y6Ubj3/MQaTN7PbmtWJzsH
ECm7shUuOanaFnEP0I6v09Q8HOWHaTXmjHKk3gIYhHz7avOUhmcxtJu4RJbA
e+zofT+cAF6ifLG3JXEiWlMqOrWGhDmylj/fNlmiBKAtYN/0iBHd0NRIdBvw
4UhtPG5RBB13JO6CGk0iRT9jQR6SpzOjYQYL3ruT72mmiwThsbCSIt3yGNWg
KP6dHy2hOhf3R7JW8oD513cjWGAwJbLzLZ9D3gSqR2I9Whjav4CLhCAXSPPS
poKzsDogkPkrDU4xOKhqbQOPJ+EqIhuiOBBv6OVrztMJzPzLVFtiUZxdNwna
gWF99m52CCUnvjDMZG9ts736tT/8zdfKCZVxUXBcpqsv9+OXQm/w0iFKKj/P
ner3zgfDDe/KVmPFDKY5CJOE2ZexfwJ0caQyq9tWTFksuIOlgd7BQ0EIyL4M
MB18YmpCP9UWfoNm6aqrR6X+kn2auu4d74y9XkWnAzSd/hNzOXD0m9Cx4/HY
eVrJSEaW8shHVV9PDOu+uAl82sgWMtE1ZodBK6hcDmr2GQcziLaEUqy5ZYDy
91+GfL8j5gdN6XPvqyxCtF7BIKG0JoGoaioiiVORBtQ7pf2WKm/fZptbhhW3
HVINOwgmYG7PqJJTIbZ7XXjDMh7UxBt3rIYYbAtHis/zT8BMfxFf2zR1fL4T
vzr1U8eLYyQs+lsQEZ3IPtT+SAx5CWrxjbGoN+mmszJ2/ScDLb9pCs7wznjk
Saa1/z6hR+XhnjNOq7H5X7XrgLbC5ov6HyJ8Nykm+4QcDDZnXvk7I7hWbNx5
UCu2MIYX0x7E6PASE4Qjt9/ODtbSQlijv5AN9sL32wQDc6TxiT6PLwQiLhDy
WM2IMYpuzgY2HDhxZ2PXwwp2+s0ZJ88CQ2ks7JSFxtbWbwauWAWledNstOWd
LVpY0Xm5PqTLKmq8LHb7Jyds0qeCZX8i+kxro1sJZ5FSnzZpmhX1ZqZMX/Xh
jzpHf80ffbmWlbgOkluihn78IIqQwjsvBuI5nJSihajNJo4HVqEB/J0ia6rf
p9cv/JcU10jRDyjHtYRDAFopOlfHGXEN0gFuMKHXwP8HSDdpc9BasIXSwt6a
2wCxWtuZcSQHb+VtJSzD7Vmz2JzRQYB7XoNdHkq7G1dTG4iEWzDpxTn1gIsT
lkybfIpBDr5lK6n1tgqZacwyksggkaAZt5vvXpZLl41sK70x9hJ+r37CdKau
NN/Q8eaXMGS0t9K0q9+TNuu8o7SNYAehkhMtXZ9mMMrGpTxXH6Np6hQG2oCd
k6zme2u4/n7wljebM5e37Gcz1/+GKodd1tGzoa5eUtN6DJhG2vUBNOPAn6D0
RHDO8okF4CckpjRM3dQ5Wk8IXQx9Q3hU0DXAkVnMtxfxu2AatTS/f/tV9/1K
FDJBZWqAqJM2cSl0B6C6LfHBbdtjlIeCdXkBCBp0PtrMiKCHgWcKRcVCJUYI
D3kPQNmJwWWny4gdjbIFdQOLJD97INsgLhem8XaH8qBkgPzmQqdfG45qUzkj
ErIHPwf234iFY69sZMDo1lV21p5aNQr66bP3UIodXLchylNoVbHYJmChyYjt
+SUu+FQWEAknVOlAZj1qFBV/1FQRxSo9iBvcXsHeyqVQK6YziFFY/nZQ620/
6uh6P5NgqLIdnT/eYWJsO8+q7fzAF+yjUuyvBo3f4lEU+UCZ/2lno5oG7peI
EvQflnAyKwvSX5saE5KGN125Aga2Mwf1PGIU0mT31Z1Y+4TIJsFCXBH51b1q
II9ouBWQnbdmqsmGlWZs+8n4lAHiEp8I5BSaPv3IuhQ8Y6QYWdK6G6mqdRK3
lF7JjS626e5GdpeFrOwHnXNuYXBXxjfo4n1szcHCoraIiV2jND++DGoYDwyg
sKLbidAwc9acOAnnuWTEwcivc4BYeFa0IJAW3+T5Nu5yowaLtui/duc0O00m
KpHqWiQZRuLUMJWLDXFeuzLpJw/5GYkC5bCfLi5HpHrzjOc6NoyqKFP8Ug5b
h+uT7VcWjLKyvcbxq3j/bUdBvJZozpikq9WAgEm2EcMJLlXQfx5Gq+Ep4ilt
z5Kca5G/jlDFsslyAfFV7OdMTrbYaJr83Cl/s+Kx1WDvJFuHEozDJqUUfSHF
GT40Kl2pwcYONiC+IGY8/UIS/fO6g/c2URADhALkUWeKPY4dkIbBgZIlo5h6
fKCjKDohjMe4FUSjRPLIDXQXKq5iBNywwNI0LME4wTy3mEjPhG8Sjlm6Nw9N
FtpR9TxMNYxnKhAB4lC1TDkdBELDv9SwhDz3E7+5UltLVBvt7kBDx5oUv0ge
m5eX7m+tfWTWgfoFD6wXFnoZQq4sFTYjYQzBPA8Uoor1RDiAq/vRzyVsR3gJ
xwo7J/rOencKFccczC16n1+FRVIwl9He2A+vbRQviUpcn/T7kRtjDyfIKw0J
4a8mumOOoC9Lsv10FBq9LVP/D9tL1E1ERQoBReCwZGqFHq6CSpnNvX1+LuTF
KgnvCVIFO8kkWYFf9hbUfD8vRm0de2NBlBa1C15plR9U2dHabXFlJSOOy/+D
HaJFV2e4nJ6U/+WqQGZNO1KPDc5WH0TFiOgsXZsTiQDwB9E1LA1P+4XBDkm/
S7uRonPt9nxBAlECpqrOpOBEeIbqq+nA+U7xZVKKsh770Kg6nNGjyHpYxzjj
d5CPWze0dfrgYzkuC0jVYMJ4R0QCfOeIkZp9rVXCE6PXteWoGgA2fjKe/zJ2
pyAggU5ixuoRVgkkQC2n2kfbiLDhiwUWORE32hXesYPleIMHhD6KggWwHU+5
8D9YmNJ0SITc49x2GqFLEg7AUP2+YM9HGtVqLkTNqjZOgCupnbZ6wg85y4He
4ePahat9GssHKjre7aT8Yu+77rMc8Ji5wIEqNtY2/V6BPMTk5r97SL8BcxMk
t1hWbM3DyfQd+3sQQqV5QhwbOhAHfFW+ZQg9CqyGxdTgJTNt6MGRI86QCErZ
9Uw3kxol4eeh2tZStFM98r86hIxsQddj0FXwl6Eukg+3XffqQ4aXzrXijdD9
m1R/nSMVle2M8Ke8wFOUYXxaY4DN27zXjFnaIgNYmxAwO9i5SwQkMjezRea1
h9vRKvRF9ACU1ICuiUnJKQqXrUry7YXWCMItgPASe+3UIh5/B/jo7xzKe8lZ
H+9PpfjN9HOdKpTWepUpHXzfnf+PMhpMan1/fBdkCEXhgz2zJaGjNxFKikXb
u7P+dsWi85V1glPC6DjRBWG0rAjnavzeyh+SaSbfg2T1f0yuLZOPTOB8VI7u
TYfOv/Z+1yXMlN/RHpSykTMswaRAzXYQzrcP2ccmTAOxQ0hHUP0BoV+PZMvS
GN4yPFg8DsOdpi/SzpG/FUA1XffNn1C/EVRyJsaEizjflRvz9I7FOWfPO4lr
5xxBfI9SsVsGsB6Cvc8UbcMvap/BUm0kWAII5bZDhKMJFfdGN0Ac269MORWC
5Yx+1FuRxMQqm3UNw/q1RoKsY6uQ4JsKagtdiQ55o5zDnVcdKUPWR1qGKI2g
0J1BZukvFtiiZrTi/o03Iu0+xPB6hQcnl+TV1OxBmOHdLqrQRet6rFPb0v5k
tVYpkcVKMa6WFhUnoencqDAtwLrauuro1htSMOkuYhoOu467bCeaJy0z3lbN
VbD8pezhvVAhqAXQzZsSXSnTWoJQQ7GX5TFqxtm+h5TBwb1icvuEVLQdgg2D
UFyyOh68ufQUzWar6w1zhyqydb6df5IqTIxL+sX7xEqrtLzWTetW4OAbWX8W
A5IjKEaXt9BJr8lelaG4sm9zHbi7QmKcSMAAENJauk4qiTxpJVJ0kEbrU/pn
AaJciVcYYzIqGY32Xs5sIP23pGeVuQrZvuLz/zA0Jof2H04lPrLktaKjNuyR
oo2aIYgB6upDmp7yybw9LsVDp4TNV9IhMFGRasBBEFBv7wZy/qL574KAyyYX
bh++xcyNZFaixIv6FBnJyQ6JWoORDpY+fYrx10QX4kfTve7gCetmRjR643Wx
fus81Y0la0jDEWFo9yg9Ooy+luUAVKdDSMuRlueqIM1/VTr1j3rSG9pQLWnS
FDeg792bmKvAVzbBVbu8L3jniIj3RUrV7I2uuA44U6oJo62yYPF3n5Iuolqm
Hiw0oGHyfVBpkBZM/U3KuYVH/vW++jusVb1/Q1YUjysXYvzIE9AMPju+BVb7
3KcqnMRs17gVtdAUX38SSGK/ywKBKsJHiTuFSc5roSl/Eb2rYlp5LPZKJgnt
OUVUey41JGAKbCrkUNf9it303Tm6Q1P1mmpjIXs78Er9FSHS94U9V7Q19KQ8
HFOqJ97+/p1plVCvbmjahhcEW8w8EXzJkffEfgzi87D6yoEkwiVdFD0/RdNg
JqtcxXf1cgEzrjbl7TzmTiqK+P6blcU7lm9u9g5vHnQtek+tTRpUORt3Ey9v
bJQcKgtII9WzL7HCrWbQ0dDP3NB5FFZgvZm/lIG2RDih1dbqPRBvlP8Xtf0X
ZVUWpNO67vM7xDROgHWGaD0GvmvuRh9gpFTJccPaDLbTuwRd0f4MuH6mFOqm
XGlARP4C4TplyP2FsIxwKAtdykObstT1HTDH0vpEjRPnNaL0F2DqZrOjKKNd
vqykjohLdhWWIp/5gtSr6s6mPhR2WK4d+xPAHALPgP00gTiHXNwQxO14Fquz
C/vvs4Ni9LAGsq8oxmbTzfYgla4TqY4w6bQceHa2+Cvog5A6ylMgsITUYMz2
iWwcF1S+yeNTDz4Iu9HljCjFyNWZ6+wcfZJBvMZfmpRDh5LOXJwb51ciQA3h
LB9jtIxYsdL4rp6kqATgFFDdpPVxnwvA7c0gBdqBbC4heAe06OYgRFaawJGc
1ySu979c++Enc5HnyxrGMX0kw7awlDeSdMP2ia4b1yPHKFMYFPhHdOut8/wG
BbaZokwstW55C83/uxP56KDxVLkgmDwxuRJEpJUrOZmxS6z9bqcjuM5ex01S
3JChnaZz0tpAzkWu4f4R4v/n52Soezw/7hJuWT4L922x/rYfkMROtYPrhic4
ARRfkf0cfEBiBZCUhOc3FJtSUNuz0S4utT4oz8OdU4UvuSeREeg66a3KImNH
65RMn6Urqx6gK5YszWIo97W9cvv2gk2sNrbhwvCD+jdmeDOOtVOcJwSbo4dO
l1dGg+E+bxjIo0DWD4NqHnaCpxvao/6QoyLKoaCDLfawk2DjXGmTSLZbnzX5
8ouZHAK/5RKXi4pIL2nN0z9U++s1YVtynEV6pXXnOTt6/QymBLuyhdymwmLt
ScxXNcWsmDuukxqTX+t/Zx3Zks296hZlSq6oHmfmmjheb+tfd5/eszLi04/+
BXisf7DBljDp13Kt46hUCmL3dBFm+EzryZjhTZDe4bC5da5kOV54EAPW0RzN
WpkFT68pOBgO/fdXT6DCa9zOxEi6IWIzKvHP1JcHnKAkpt7R2NetVK/yrtwJ
SszDyhPT1jWFPM6ES6BfH7DQaE8EMFnn+zom7oWN37NmdyJ0CxVZ7Xnm5kMw
Xk42M+X2pK0nPyALOirSBQ8V0NcuKRIiA59Vw46/QJXXgDSltVnLmwylIkug
2iVvmJ6bkiVyLKCNH0NUeH7FHkciGN0jq63jWkl7u1uGDJ865QMO9hc3ClvU
ofwrP/snny5GBIbr06T8dOSSS426r4eqvRmS86M7rChajlIK7yXNDLtRAqs9
ouqLrYuLWNVLvzeREvQrFZ7M04AqVTxUcpu4GdqyzoYswvbxS2sNd7Hy5AjT
tIA0BdGGHQnTgPUhaAcQDOQd8t8txEF3fU0FR0VlCSYy69FQQ9Z2bHQ2WWam
wQWyqh6kTqMlC/j+cdswkRMI/dCWzwK5htRcBEIkrSqYTI1i07B1UNpRp28K
/MeCUqAUQWvoVo/vGfjTuw4ApG4GZ6hW2ko1euggBxx3tCA8mYm5QT5RxDdk
J7U8X10LsP7/D0c6Wc29lnXYLQ+ZZCg1c4qtnP/DCEN5rJ/m6aKZVWDhKa5w
zyL9KxK0XRX8WLgQGqf+wb+9Xefrf98SGNQi8IR2tvuyPpFsy1Mt/WdyphGt
OEg5bFCoQxUzPjuh76BnMdSrLW2tarTHzvGn7pOon8mb5wkFML6zm1r3hmlT
h2SjAyPf8D8xMFUsp382OKrvqQhWDfYam76/ckoXwFIjGJGXdpFPUHDiyahb
EBdREzAn++xDlXq9UwAXOKr3seDG28ei2lfK6byDkqvo96dnlXb61auNZGvd
4ktMy05U02EuQdnWgwWykXMbXVePyhCo+Izq/I5ichMh+qIdMiH6Yso7fjGQ
koQ8fkOY1hkb5Qp/9C1D7y5ub9VcfUSwFhKZXn2xXjS9XbUAltNdu+U7BQqc
tpKFZSiQI1PJUNeo/1KCaiIa1KPbgwthwNGTPpR4gkh95O/Fmm0ngWEUA8gW
RccLkkV0nPsZ3Z7Lg+wW2NCr/J831I6zxbQN3XepMv9ZpLLwjYR3CqykDso/
JaoxqUQJGP7rHjeUMyJ+3Y3gylSeHYaaRdRWzTqUs+RhjNuVsBzu0Ll9vX4T
ujF4xaMGWtarZvhl8gEKNR9R/QFZ8fqabLi4nVcJ+ugrPeYwNX9RCCCZEipI
xrZ5ev+bznnFA4zOR3e6LQUcTXvUxuav7saxG7vATr4McossQW6MZm1fjfOO
MpZIKH59+NdBu6sRqprhKR7wQaYO/ytIJuIF2E/QrF7mbCxStQ4tDi03kt56
HN0exrjNTw/BIprTeL0XUzqnQiSCzIKB/IswzJiuPnkFP3/xqvD/TEa6TRjn
ew9CbrpcS+RFqDxL334dJD+RIpTYV1AXtWrFJoxpROAIDmeApEDJ0fgUcvJ/
kBJPrqzlJPqNRZ7EWwuENqihP1J42j4kK13lvhTde/+A+txVIgZRRqEpyKvf
3/ge5mVmEzM9HOPAfycw567U3CEgl5gql5SYfaAWHS1PWgXivqmGch9qxS/V
6v4tPvCwz9RviUioXKbaz7+08W920ReASa73hx/jK2ZAK1poFM6UpLh+593F
1qjOTQCYUo2g+Up8A5YFOU9g5BkAZer6TT6+8VRWJ0f+3BcFjbMLJ9SyS5bl
R2LUAjNd+heJ3b4IgDSKXAcE7ZgJ1Zr6wnfXp4SlPX6e44CVZx4GfLtKNdJA
GRxG6hW3P/SD4ttNuRfmwS6w5zbH/SVH/YRt3oz+j/6dRwgT5lME9GNf9Dth
qrbUEEA3IjUg9ZumorS1ZXd37KEZHz2exBkpbqWuO05sG1mLBJHnd6oFCLWB
xHPyxY0VP89ywDYicNAWaAM+hRHOwycxtt9WwvoQAgLiyLhmv0E7uwijAq0u
2P9avDtZGQ5TJtOBIc3Tm1cOAFMCaJLi3tTX5yVPR+qy91YITQu9EqogJu8n
6kyjzfbgOpjOtWLiruWm4ShMgl7u+1oZL8f4M46+141HAbOq96Lbf0KoVK5B
wjMGg265ZoCRIDA0KePuzGqMPhSDOjCyyhvMgNbg8XxbC+e4xvNdoJSWoq1s
apquH9sgyXKCvd13L3lNwlFV43p/YMNrWTBZ7/dLyubx5zKYm8JjRNLhiXyW
M3H5zZnDcUqy3eWr3r1DsnGExwQ9hUVVUee9IOJfR59kWtnhJSLWydZERS0X
RwiWeiXPUs3I5uWj4ovJ0m6PwOtoSycBROnYr3yvTEvRsZ0GNbG2BMu8Z0Ec
RjfddaA+HBHXJzf0ekIeZAjsGFIA8wbb1W6uX7/3XCPsCyE2TD5GxTKbfIuH
XQd9PJXQ071q9cInOOjQ1lr6bAa2glYfxey/grCqZ9yWXAaemzK9BNCQqbtd
3RpaksCW6uNBRHe6OYam2KAL/sALHPrfVhNZrz9POwtJFswZFSAgXd2T8eRY
K+3pXTZCjTloEDrmlV6in7wmePsLGjW8QFoL5ua0wWneDmwCkX7XE6LhQ99s
zcCJtS8ga9zHgNhQbvciZmMEmH3ra1mjRJpGWymAbgIbdbw+tq/DX+Th4oEY
DDZggSyOPrbtUq1DiaXmL4AhmEBU9716Gtix1gmLek9FKPKLEeSxELl5Pvzy
hpHoAu6UXMyL06kzlmJckItIHs4lhMNpKVL2iL+MoVJ2tTsWgfCYIuZ2CDdR
+ivQKGFgkBPH62V5ckLqSd0v3NMg0E4bYQhOvUYe66BGuY90OJ9yX+iTP41s
H6xoj0drCgPavFVkF7s16009eUfm2CJ9iAoMnMBkT3PG6udWv4JFee1qfImT
O8R8VuMpCWna80zCBXjqIXLhUSsbhPqAmZSwhC0TCPKvzYUaBxNKmzuKaqUE
awHf9SoaWLS2VIFtnWbmcuYtOGntCbF19SS/mxHxI+C1HOI2rZalBBbIrSSd
C2a3c+kvIptTRBe+ELgLxdgJVu4BKoMweqJkxl+Zty3z9QboYFt4MMRRazPH
0nWsuXEZ4/0NOSL6r+7wk20BqBgYmsIe8jo65vqcLSKL6ROt1bzY3Xqujkcs
b1by4PBwK0dvmVBaPiWL6j3MPmrVybbB6IJZKS9tgDAtXt/bJyyAd2aKqluI
5S1C6PrbvSAqsLSzevuyiTcyKvXlRexQ2A2gdyt0m7h8X2lKjswYj0kSoS2u
IHeB9xQ2s/cO5QGDdtiVIlyDEJkJt0iq8QP4tGJrieUdWGCkkBrnGJ8an9ZO
7o1vKD+DP+Wo43oRWUKszaswmFSsSF4r7VHLQM8vovHvdGAm6yzqNRGVB7la
CG3YOiBQeHtQa+vXMrH3IYyf3xXDJDcuCQvAZXTt05MVzySEzOwNw3vLDZQP
aRrW6/06qn0S+nwPzl7Rn2L0wH9YxQc2HH2ymr4wEAQJJY3zb68LOo5JqmY/
ozcZhU9uRHU7s2WORXJ9OWr9ThLq9Vo//fbmhrcDWLR2/8/Tj911ajV20p9p
5BqnVEqa0Bf73zqRPgV0xp3t4WKPABRnnEOojFXg5kk/QopHr9BPfKiR6cPT
HbJUKHqrGkmWv2Q5rFLybQAq/Z7WNi93zkwPcXU7ChkAMQs96v4/h/P9JX1r
KhHGIGDs1gcS0wBoNrGurItmdLJDwRyb8UU1J4p0Asv5cnKKf7JdnXMY3giU
djNMxUf675GDiVjvTy6Iytlb1hjISbkOA19ZM+fxYNrU7AIIx1VDVEBDW0su
QWwrTyUc+zTEoI5BsCzVUO8mBrUCxz48yQ3kZctcAGwXuyMOAFYvwWMKOAIR
S9Fnema95WCbLH4NhOGPgmiaxZT95DBP2c67FFa/vbkOFpCKKeIb4+gSqlIX
6tMacF+ED26vs54Y9iR/nChQAnB4HUYtr59qTTINhakYFBJclvxGFt9+1YTp
IbX/jDoh2jUSLBz1GRXpieebfBF0vnzmVCzHWnmPoL7ckDZbGHhY4PK1+yIR
YhFc+QjMTkcYzX9kFmoH2o0NFA92/p/kyrS53nv04TEBGLQU8Hgjgp0d1GpD
OOHFI3yCuxWjp9Q0kFn0ID3IzuqPQ0vLQwWqge07t7+OW3ttXSs7Zs+3s5sr
7k86fKhZd+jeinNfgF8UsN2kzwo+zNEK3Ho2QSF/eVWY7g7oS0o5PQgMi9Vk
OcYQ40k4u8UmMGfdur6qqqoC6JxURyzqbZbLEo6boBmZcwiHV4egN5GIO1gT
3A5QZdcU3y7mKl/9jAhW0u38fY/V+B68cGSl+qtUsgNNbQDTGdjiqOQX4a97
i/Dz3K1i5eb7C6K7tHKDOwdIy7tPwXBBXwFunfs5jPuOMaKCwROa7LDRqtqe
c25MoG3ivs2m5O/SGrcx5P8Ugny2s2mQpXWumaVjXqB5W8+Pi1kKlIUTvr+7
Ej1tidMg/NKwCa638FTGIINLJcxSwgPyyqrceQnB5jO8dpjC+zdO0+mY+xAt
GoGdqVWINwEBJBtNOK3o22cW+6QEsz0MUDuDzVYhx7CluvvyrwguKWsqxw0d
uj4sR/HxYVSCqPR8MWxYqcMIkPzqxnG8jguSk7aVFAVOYJ6Vo8R1aaVGibX/
5MqsxY9fEzh1p25P8CJlkHlOOtG49nIIw5neED3/yW8o0e+rU34EL4Bgkhtp
s5Zx9qkNXBLW+XG+DCWoBrJff4+g3T1JHsvzsmCe/mcCrt/5giQii9yW5Vtu
A0iRM+o/sptYMdgwsjZ0JwSPcwdz78OkfksfOeMw/R8XUlTXBCsyB89Axh1z
yBmA2/TUQNX1+iaPjq3n0RxHXrcD8bF1j/95zfCtVIE6xLPYNIwgc4KYHSyZ
qT5jkba9zXZY8EzOPN71rEpJQKyzsyBPWvplyjILmwV8FyBBHS/cGWBibqlm
RkN0MqjASFCxaVMFPaM1sDSHueBj+J4O2xh6jnfZ63e9UgCcOMgwEQ9pwx02
B4uYq0SB5JCzTBDRPq+0Svwvp0vWUHfEyOv6iLkDhKdtGX8c8sKtk8lpPwM2
1sMxukD/FP2j7AWtRyRaUgEAYzH3w1+l+RIBSzB/cZzYVXCKVWZ0dF2GDTmd
g+zOj7m2jKJ7e14zIg08ZMUzfX78DGPS+h7LuunYqEDdyP6xp6CBQiy1/bXe
BmXA7OO/0ptkqFJ7ud3ZCYgZPuHO615F+TrJ1NjjVk02xlNMH+7UuywChPS3
YQhWYrXixysg+4lOQ2eKj3pxJ7LAtvxZ0UEBBRrLJMj6UhJ03Qp6zutD/UPh
sQmNd4c/99IfndVhgvpEP34HJOxMBNqCpe0Ur6H30Ot++L2xfRATRoLjNL4+
3zh7WalbKAUa2bHp+2EO3ZuoffZjg6Lr0RubxFsYezDGWTulC4EC9+N0Oi0E
0S6KIHT1La4wv+isnosLfPJn52JL1sFUm3ilb3jx4fJOY5rvP7otRtRfWOoy
crEhFVu3XMtaDkYev1COPWP4i2pxM/EzEkVThWc5BSiCCN5FY/7G7zrr/W0I
61iBgt1Kl5ecpyOZzEwCcklaLGMGxWQZmSuJfW5ZSt6gjagW25qkQGOARIuF
nsp6CNJ8FfErxZh77S/SekTGak8280TDB1gDRK3XDpv3odEAchEACFd03cIC
e9/bbNVUvT8xabBMAijYRoJZKO3v9fPBqhtdIgiP8NfohRXyZD9DCiQgnezL
gcMDeI6eYNVn3VbGw0xeLhKfIuEnQnqEETp2q7Rhy8UyBsBTLXvQQyTdPOwP
0wppRvmos2j89p9l0Qcr6fgFfdTnAEkfy2NtkEModMmhWvjUSPrQ+KaTKvl8
SzoZZa6suXOrLdDfiHxq62ptPPaBuGtalUdgKiCeQ66/ZZJGLFHy34S9vH1H
izmkgyVyBGB3+4JqDc1cx79MN7ViEy/tKCCSUUYBm+5gWL5JWu4Y+yyX9uQN
U9LF9wTc2PPbJNkH/zpP6tMhMXYS5aFLZglB1Ff0r29oeOzMnZ+hhMFK9g2M
UwMa81V5ER68ht4ywais7Exf/uH/VDmWyV79NgFaqCsn/XaM1VknzzGO+cTp
bw3kFkwjxhkTu7xKff84KXXUDSA7YY/fOlrYK6Wyaj8ooRcxuKKA1dCLPk8K
oshRWXtl4PVxW5k49tl8vNCUVf0flmKsNAlA7+wyKEicuLOKfzuDdDGWaDab
YwbpxcXv52mCj7rScS8siwG65ahKzlFglYViw5BqapRS3qHoxDwOJu5G4e9N
8GRWxMlsq4jM7JlUM8X172ZfhItboAyxttkInaASK0wD9qYdzzaAPUDuNX7O
wHzekJXx44Nf1475YC7frS7rcSlLxNF0bcGpERU6PFRRWfTlk+VntnjEYPkO
01t45Bj1Rm5DoukfNzjbBHfst3Bzy42Jk29aZw4OKS2G0sUoEy43GIvcUtQR
NWOtwjXpU6VJdzLt2KOAZ28/NNo7TXHwJjUE4flaWrh5TB5SspJ+76TNcbrl
rQNlxF1+38nfAvDhnpma5mFA1v0OhtprCqtM1gKNrnrPtm5N12E0ZJuQwCUY
njDGUF2i8Kodub7RCVUkbxg1UDiwh2Bg+UT+hlyeIE1CesJbCdmfdzGSp8pk
uYuWVHlOpW60IUkZKhGvDw/EH2RHeCefzI3i8Nsu6VgbWXEp08rRootSrw5Z
hMvQ025flqJYN4a+mhWfgY6REDxr3E5ipt0OyqxKvN/IC9Pdp8HDPutV01UM
ZbZTyFMNW+odhrtVyxz1dgXNfGnQltnQ/3zh4JvG4zRZXmCp1m1TBW5cIMZI
oGhdOnY1p/nmTH9WaiSqD+bcKowuwzZKBw0XEDQd3nrj5VJjm9dqRN4U2Os7
V1Zb4cI+s5JZwOeoXekTu9upr0/wXVGHFVB7flhwm4KEP9cHBibS0TPbCbH0
Hi6k00eMKM04G8L+3c+Kqfdl7Ma7D2AX4WdnwtPjiaZfFV43bZ9zyjjFhM4D
QMEejB7ViN0j51MLtW4VB76rYhhae+r4bWGzqfbcv2On5NzQj7dFxl+bWV6e
8NQR9zCSiMWtCbY0xnreXChqzYWposC3k9IQ4uoP/NC/9QjjDGBE1PNmaUCo
46iJk+0i90onpjrhCbIhMbeblpB212qrB8MRl06g+npl6IIUCet3t1xt356B
dP8cgPbBqeZny6ugHRvsnfU3TSxDXByRiRb3mGhNkOIhnYL1Xc5q/Tsy3EMg
0hOoYW35Lf0M8xML5xiVtbnEEEHRFR1hRTcRR3iQrmI3mUDpXjfv8JZIuQqo
GFWYaesQTuUIFfhGM75S42bjZJbhCuZp5lBoL1PGADeyoSPzZR1mIgPguiPL
ftVZnjNSh3fjEQIDVqLEVechGvURUql6OfuW/Nv/LKx8kaFskiIQz1pHs3RG
kUbCZ+LSJPyqwtZuibys+IGN/DkiTk0GYqz0J1XfSmdKmJZPZfdUzFCYkFrB
EPg/eHTzBKmGT9VoJjmGHe4zob6XlfcbIhYq857JkUxz4In9/tmJpPUIAmrz
tCCTBYFLhzikzGR8UZ18+Mohkpa/zECZ2Ug2Nij6/rgEqf0EpheVeLMOiSLU
UC3+o7uHqG7zAJ89EJu2V0sFSEO78/8SujSXtsxqPwJ3i3vOB7GLe9myhE4q
EknY9rsGhKry4lS1A9nSXPStreKGfWPygRUcW1gYDkqNQ4jIEwmlKp3SFtJZ
5ioC5iPsvMGpi3MuqFyWm9qO8sqoJpO8X0EFYdBeYdEDd7+TDmTvkSmYY4Xj
qDLIche7BTHy/4yOZMbzZ+4vLsGUfRWtNCNWRZQoqFLjQ2cuq8J1q4zn6hh9
lm3TN5RWTohU6/eWqoEJOiYYcwDqDdEFNzUw9ZL+OHa6LrWNC0Jm9+tyZESO
V/v1G045mUsl2gaZ/L3C1f6gEtL6WvkYmudY634uhmKucSd68CA0sifRrw0i
DazwnQdi7GWvnVpSqXDxIPGz0QB6PSwyGKNk3eLCNCnajkWI1HUDupyb0/Z9
Mkszm9Iv5Ypk4DSfOpA06Flo+A7oOvFGJzF/yFhquERFcit9lAQNRX6ONtw4
YLqvkj3lTi9c0eDTL+eniL6TKoECbNDKmSxnJzsEaS8+xuFmj0Ari6ThYlO3
t9HOM0DJx6LJB/AcVPbisD03m0L/sgkxM9i0WDLXL9ppR2T3H52KGyW91JxN
26tFaHhUILQPWnBT2Bg5FP2cDbb/3d3geft/R2NH/eZErq9fNy+xEOzEtkY6
q6tQnZ1X/Ets/+AL3P8TjPixaOn9eddZJBahj096Jjus5XwWEW9OCflNMuyK
rrRAZRpAK6pnIzj+208iTTo6mwdpplvfsD4P6v6xmqCnCPaEMjqSFaTTMSEv
hVZaiEQUoD7HehE+VEM9qr0AO3kx3pzcSiCt+N40cprbbBryeeQaqSiBi5Lq
lrU4SkQUdxgLEPKGpcMe0xKZy79Usm4Ektu21QJXE7MCUpM4U4fa7yP+XyR0
K6LFwjsOGPqmoTjySwi0tk/KcHmwzTP1/EtvFgO/ccMd2DKg8dA9JGPxH2tp
mojVpt1oakgxuKvyZelGB67QM3Gph+15u/gbB+XxRvRqQR5tgBFvqQM2FNcT
m3jhHs36HdEY4uZiuy76ybvcpqMnDSdgy4k/cBIJbCPYZSjXTTtatJ3niQz/
B5Vpn6Ahfxv4UzrElfVb34e1BImQ1RZt7w6paT2w3ccsYdP5SlElza89sL+l
QQnGKF0MXE67r9ehFlo32no1E2uV1oA/zu1N0vSNVwlfpYgJTN3bfG9+lwe4
XTIk8LusQOGoUyX8q4Al68fRF+ANP0szc13Bo7ekNLHgXHU+/rrFpf0Y1eZ0
aIkG6msjaiFrXr9UrhoEkgnTPJSsEuHUJ4Z7DPdtC52k0gwOwrJma4Bumstk
GaWdlR5QsYp3ozd6M5kEveBfAxmKceXM6B8vF7qfUxwnIx+d6uYD8OYVaKn/
sR+PlXnTQzmOfKDydc+MD1yJW/hodRjW1Mdur3Vysh6wLo4xARTFliSlBIx9
BtzLY5gEAcfmERTcxypl2gXSjAm5dWwYbvJi3KX1x378hhEG0IIZqkYZaQsE
um2FH/QOlVax4ET6SmD+VVNo6B/JSMg1iHLBNMrlY/V5Nz80o6YD27jfr/Hz
VxG9gIHhaHB4Ja/rzti6hvj+d4A3G6mROrwo0T3KzhcnhZ+RwIHwld4IOkAr
lDr/rpdJZsGK1bJ4/Eq2n1RAnd9U2CRAy9WE47z0Hu8MJBobtUlDt3JcyhBv
1BxoNtA/MoczTJJ6U3UcCY+S9zHyketjLMDBGnDnIjEfWckBVR28aoLAN9Fb
b8UlrIjegVd5AWwZ1U7+tk11uCUl3CJRiLKKLb+l9Pdc71gksoQA5GQqxU6t
l/adRmnCfY3d9Nuqug+j/0GZRZOYnmFjqve0JtwHmrvD28YPJO6PfHJoRuGV
fY/Pi5aBjvHCc8o219gW8H2sDX9lWC0yBQthaUQRp/A9/I9WsYynTngfcO00
/QMYCLex2iPI6PvRD14vC2rDPsQJ1k9Jx+eZGznPaplSzhwukAp5Hyu3HT5+
RbrXl5E9VQG8T+/i8iFulJEJdoLJgWAXDEdkh9KcEKe5wdBfNkxOdKNTOgPt
IjZkaUf+Ttu5NYPUheT1LHe5Wl5RIrJAVAjI5/kqbV2joN2Ll97uS960U064
sJEaR8YqdcK/qpraLrAOSUbgpkCFfvry7VAxpWBbrpPTkDYppycZahYvJjqO
tVRxuzHe/ky92k4FFMCs7a7eMPGjW2YiGJyn8onut2iCVGdNegrCmdb7r3NH
3uANqb/9VPIG/O1dWKrBCH/BUr0I2trRZTJPiE5J/bzjD1T2xYLxzvMqX8km
KxglfThejyVI6wANBBiM7CGvd+EAA+XJmBM3Zuax1aPpzbjEMsKQfAZ/gvYa
0iMir7Y6HF6pPZm0Z2gECddb3/v5I2ULno/nV4kJkcaLEMMAcx8+GU0v6oIe
cKFUKwqOTQJ8Tm4XaQAHZAI1v6wvtQKq8fHnmDqZYbjNB1aVgiCnjrIGZLQZ
MN3/zENs3xkKnOHJqWDVmLVfFYUKjUjvyfDYI89YtgGSzssRa+SGoR8olABA
XnSzkYNz62ZJRCHMb66LmEYnvX4on3iJuXdCFZkHdQarHKRvuDpNnteb4TTp
92jA5oOgZRpr2LT+pWFEs+eo/jEcPoENqZAOKsm6QFh2oi4QkVXLRfmRAK7V
AvkA19b+X9z8+54okrB6/YJ66X3A6dQ6hFfSBxE8jHqG/4TSAcS18PfySoR5
Dekuh8UOm6LbxIkpYKkFnck7NyH6ix+bgJ1AU819kTwDJq7YZ2ShzwV+K+Vg
wzzt4MGix4t0dnDp592iC5CBFMcmWGdxtJcrATXkghobKb5EjtdZeZZx2iBi
m/Wp1EK9m/gObAiZ0MKR/wlybgxP+sNuczwd3isCyNOdzcmCYR81MEi3hw/f
4id3ZVDQGHAw7mwpIxiWXAH86GURDdcDIgyanTI/XxjAB1EoALWAhItGaOEN
UYl0k+0UobAZq/YubAVTCs0keKnNlA72ugbtwUc5+TpClcifVLivUHZfJ8yr
rlgYk4Z37VErrGsSywD/U7RCC3QN/aGQUUdw2qh0g2jOGKfkwqZ3jZY4rWBO
rQp4xH00z9im8ZMCqBqO3sYc7ffijn91/P2QufUJk6RD4+YUxusGDM7BtB2f
QcA3S3rCRedJIFtiG40XqW5VrzzqEfrHl8sBw1AUySwOevEqQkRqFsW+bMju
ZQKA7tY3ubvaWZcAbjomMlNNf2NXFlwBHavZZly2OkBHeRvoy4ydg5A7r8Ly
SgXUVlDP1oLZZwzMrEBfsIUUBG+HSz+XTchErguK+piLlJZdO9DEwyfoGAK+
OkYlI5DQbtwhDsRHvxcHJ3qDRrFJ82hqY/fotp9KQqMsGzczebMjJqCsP8zT
7h3kkd8aptgf8CCvPLBIaeaeWvNoQ470UkV5V/2nI7nEL9gipskSHe4lrsz8
Ri8L+kbCSR2qNHluRI5Np7Rj/yegSyJbdbyBR5yJrKl5RlyTYhsVb9ErDHcO
dNY6DAq3o4YpCeVkP86zJrVsv9bXehCZA5KicTHNbYdcEzt/MM0rtot5nAKV
TDBzMJOZz+dIUzyEv1J3E6ASojA62mxRrHiulcjyZwATsTOrlqbz/HRMhSth
XI8sE+T4zjphbfAksOfHjRAeIkxCT7VoHf1yK1VpPKRdlOx24wkGEk/IEPzE
T8ImSuUQyjMfw/M3OyhOeANlIVNMdcMxYI8l+aGYvU2yoWUKJwP+51h7PBGv
avqOljj1TJRz5B+u+CLv+ei6aXddOiA4UqIuz2PYR3neBriVnLZa4R4cEd44
VsNk8//b/1QUUuQ8BaUPmF/kxPPuclz3VR80mRCsN4WbU7al3CJMcSN0kEj2
iBew/VhqkU+PTg2ZqBiMbNDZ8wvs7lSruROA5Elqne/tuhheJpjuefg6j5a8
i700Oy7pTsyI1uB9EJip+kLCy81TKRpmhsnct+ifuUF3HNGep4MTKHM867Qo
w2BzzfiXOXwOiEuGVFIXJwAcAdoYapHXcsFvO8mZ/wlTlr99TZ1LfEyTm2yI
sWJic6Z21RQ02B/Pfb22oaiSiMsWwepH0Bn9RV0DyN6/+puFJuHjyU7OoCiZ
WktXw8HzQNAf0urFEJGERoFkUVu2OI2ASoY8ieq0tMZ8S7WHDh9e31wiGlpi
J+R5iAPvU4K9Ngo8fhW27PLV+gfRWYGTko/eNZK3lRyL0nGkWJPN/7/7bjnL
1YNWGKJSVdZpbdIs+j7wtwNXAeyhV32g+efMVG02qOhei1gSVHRN/QiBqEOC
p6g9GCzGQ+brdFpzIvuNvGgNn+8reAHRsEfN7/5Tq5Irkic2px0zX/ukS7Hq
lCma1PP/rLTkhW0w9l74UmTsW40Y9JtlM++H1PbDaga/pWTEKrNYlfE/8AWi
HfKb7fYrzG0lvFC7p6Q24lnfT+KO44a6NmlpyOeLNbB8992Rxbrb6HKTTnK8
OEtZW+Rg2oYqinMBuJ/agVJ2ofoLDlNE/iYHcQynb6n1aeOev1dHH9HTwWY6
ZP5dyoZ3ECOOBbUfqAWEXrjPAe5uprWNymQaoEqh28Jh6R/KePFSvqchD+c5
a8H3rZdS1FfyXnJd3S1r+vcibZLOM7PCu8nYiEAtCJ8I2+vB7xdzz3G17gdx
4OLyGrQeOF6fZbmt5qMgsLbQza32GsOztA+CWfu1pPAAl3/dG2FomPQZ51Ok
3/3lmuDwgK2M9BGU01wGN1AuSsVOl92m90Kz6CmjPTV4JfKm3/UBC62RPleW
krga6QxtUXlN2RUouMNeKdDgIng7Dpjt6zT92prNchz2tle8cub2YQyJGC9G
Lk4e/D3DvYVEtRB8900DRIxPaqeg+mtg/lBDXzSyEcEvBeBcbPkeqH5Xd/AB
lKiTy27Gn3iKH+0cs5t6KpJSu17LQtK9HgE/PeJ9zcfAHAPrfRYvtm3eCrA+
6QtbVFdt9g6RHTY9FUc0A6c9e+ZAacpHPb+IW4YQ+wjO3AbtyawP6bFtXWcv
0gQXdf/yG9Fzrvj+r+V32qWjF1mEAYUkn37sMGrAeF/pzDDca2uA8tafYHr9
EqcJrrmUwMa06U++txKWoKoLyN4vXLCMsZHBs2FPxp1VWXNa6Za0aCskQCEw
2NKtRYafR7Qh0qzwmMge1Z4nwEk7DShD2YgBvgEkn+Yz8xdsQQj13PJqlsX+
Ia4tZPrYQO8lEKar67YNDnvcGgo7BpB2xjiaOd5ZduJ6tXtM/0+vDCWH0K9p
2I7JxkGfO5yLKcrhHTWj9qGym3uNoXokKTPUpX8NhiswPA8mg6yRahp3Zg5C
0z5n9RFRQAefZTNeJYAV6Dib0m2y/wwCzFK7GNDYBhvARjadpNIG2DsjBXID
tTAuZo3iJyuITUUa9AnDmwWlem10yYpEVP9vcPvHbXAA43OiVD9vdVA9CPPe
GCcZEFO2Jp+f2sJzLtdd2BgYlcRtocF1Q+AlSnwkeRqC/zJvhYD15OzP/Vdp
2QeOG2MUqyjs75W5HMwNEJZeuMf98zOBbTjHWgiivOF4oDdwN5bE0BaiTv4S
3cgVyxCUEECpX13n5z9e1ZTHt+IPzwhBP7lJZ6IZncliXB+DzV9WVUqj2rbE
MDM8LFH7qh4UfyKw5yqZx2ef87/ImwTh21JTZ6izLCct4mEVG4q6/kef1h2X
TXFEEVJ0XPOkDKRCI4Po1iYu6nCKye9C9Jvjgt/AE/UFaWONBRJmdU8BOpJX
MBaBQP370V4dut0ZtOpdibrUdhMjf0/ClfvwtpNAOn7X3QOrQjIeXygFi6v5
amjssUwSdiJy570E+rcNg6RKeDd0LGE0SGHKtTt0viDGLXQ+f/zsOGNzEOum
EjgXeXSgVnppppB/TmvL8ner9RcUd28k+2CLTGbC0Joo4fzmVIwB4sodvQSL
zoFQYTP0yCcriCWmnPvGLDwz91qrhyPTRari94k/5Hq25ilDNGLJkBDf0hAc
QFOsw+kv15YU/rqeUL/oYCHwBCQJnRWmPmryGdPogRWWhlpwe9k1fgMhsg5c
AuLEY3/8kNzvgeZ1fOxSu8MOzeQznsdgbMwiA8HM/zVTTxz9I2SNjBa9JwQa
Q5hae6MHzdq2tuaC/mQf2GzZIddp6kwNY1H6t+q46QdOlsRfHE345VkC2Zof
ZWfVh2VK2o5GbaZcsW5Jps0p4FdLLYdoma2PFySEBJLxv76YkwwzFBpND4nC
0NdYgU5W65TZImJXXiFjFG/bAiNxAtpsqVhMtvCKwpYFIpSzWpHMPu8Xh63E
yfJ+8kxR9YSEGlL6bpmp77n/5YpsxK/Uy9DlT3ZE0w2zf7P68DUOeHuz0JYP
IfORAPPyrcvsVshP3EQ5xnPPo9yzUKfPkZQb85uhXBZ/9VpvgOyLP3sB99Q6
+zuuimKhyXpWpipvoT/SgqEHBG+bt9zLARdUlDTeH9fMG+mPO4VoY4hJSiQf
CNzroKCzPhg0C68g/US/qSn84SJmopyX7+tqdXChF1x87wWLCd0f85qPhOfy
KqM17J6aDM4A5Mfwd3shGUlvHY/5uEVHMMUpee9Sl3LtQLjdE8y2TfE59r8e
4tMNJuyaEpD4ymsWh2viUA7N1/3ilBmL9UoX+3+JWlOcw3l1yBwKjvrpNY52
On9c5cVSIL2Tc6ILE9YVg+owZ2Q6ElYx6nKLgR6iXDG7/a5TTEVdgwgAQqka
Uny8c4zNEsx6Fyx5CitQrBGefV/IXA1984xIFk8jWCr2DFXz3zoOF7Bxw/td
ZRj7/dG07UxHaJUp/j6hvW0QCE6KMKGhfgdgciz+XmIgMU24RvyxLbNOWoDP
u4GQoIKsWq+xzi2JqHSFhaWjb313MABE+m+UP8eKw/OAH3E7F0foUw6QDFr7
1D51UJltA82x2Pt//+Jn99OK7CZgT3gaCTPO0xwLQaQtVOLkyg5nWenY17dS
3fwpcc8UFrNE1Ndgm136IfUCyPhXgBCthCSwJr4zxX/f6masGV3SiQEfgLgT
lULvVx/+dMad+xAnr2Ta6tNiEMkicibL6aeHvCiErK2E56uFUJTq0Bn9Hxof
AAVlYlhIU3NxyCstzoooTFIpAgkfxJhtpTwsNWvyU2wPf2dhUKKh1o/agqkO
NqXmxSXBwGrj3Z8u8Ezg5FQOp3DVulE5WpSzRH8ocmj1crAfvQWQDJUnE4gJ
4CXteHtmiNperpnGb2fZq34GXXlRx+/P5A+fEjyotFGL8JnJGwmKhdXBLvyu
jYVabqhaGBVKxGX8/p/s3EujSKWkFcGHKdzDQv3dLyh6fGfkh/Ssc+GbNsGn
W3RQA/cijqnluiDx91lgoPk+xkkp8Ap+eDLWoI4DkQPH24UW33F/Fno8Syx2
VUlxb+2nFbQNC8vS30JPOn997q1ioZYFkmVst8DtXAJ9QdLSg1ywPyaSnj9I
JCOqD4SMsoCII85XvyZoh3YhVYHiap7cYFZbR/ruYxBdIT8981ZTDgztS/ph
ojPDav8IR6dKso5/kYLDuGDbg8XQQx91sbWGYXUOQkDUthzh3QHpfl7qsiFk
euviS1Mkv51Lt6Op/8+5vDsD/UrSEaImLcAxoL+FQerzC4cAO/DsV3LMp/zt
oCO+OZOvV+LfhVsyZKvHER3xCuh/8OcAfSoCjopCrZwqsRTSlW/7KvHfeCTg
dXtea9AS3PN5RzAlzXLxYmc99WKg3q68te6qdHhPhUpAQkHUrWpFV9JEMPa6
RzDbcOLksa4100BFlQGNh0nWjnLYPndVRyb7IZRqonQdOqT6XEwOlAGmefl2
0NMZ6XjfU9L+KtRDsNC7X05Z57FJxLJz222fpxkDMfxnAIW5bnM7/MYEO8XX
pbqhYLU0RSOUHQOh201ic8nSPyvtCB2puS+cGv3bg885Xl7dbQT+LUQVWLSQ
rg4PAVkJErRO62+XzFAC2f/2OfXSd54a16T9GWGO838FadjUbs7E/TkkNMoc
UwsS3gR5MWiDyvPzsWMAeqq8hq1Zfq4ec4Jje2QUSlfWr/n4a5REfMM19JQN
+DHJbE5kT2eYxxNTriBERl4x8lRAnUUI1ZC4AMpCxNqEpFwOSKOjkTU2JTXo
rCKXu5UCh46vgUek3ezlcbgrNsCQ/EiwuMcealaJXrcojMMhmIzhbFL1h1AF
13felyMUJLByne9M/S66wNBBsTi/ZBHWT7j5e5ZtIacIbqHT1jL01cufOWYp
UVdAkRCyqNjCIcymxjy+MfWLX8Jv2DoOLUYOawq4JwtbkCESzgA78/gLKgTN
hoZf9BFMxMA6opIcD9oTupM8XyMB9d26Lpy5eh8nNvQ6P+qIG8W9BDqUbTzS
sQQKSBhVDPi8S3BuguUKh83bunmhkDVK/z0Dw02HwY5ox/WiG4iaQVBpvUsp
5DLbgkP71bvq9zHOeSns3ji+cetyuYYG9ETsHpU4EIYZkp0fYCxiwXjbcvEv
XcCTZaZrPauc1LD5fNn8YojixW/oP3KO6VSgb+I7D7ulJQOjVZqi71q2aCIs
bjLHOqrHEiUGoLlCE7c5ooLCXq7mwnIpVYhTL39RLWsiBdiklOUgUcyuhsKX
MV/fJFVZcuPf4C92sw51dPlu1Iqrp3WSdqWGm5tsYGPYf/lvd4R8O1t+QlYn
hNl2eb76C4ybZa9GC8HrHlD8SUqSlcxqMgNkORdB7TZRsLTu6VgXmtRFnOsm
H+1hHWzktbubQJGLXXxRJtI8B629DecQkB+/RKwIk8TKmo6Hw+jwkpFXqog7
zwI1kRZoNJso1nrja9f4r09m2ak6KrS/mO+EH7Nobwi8ZuwWTRpTn0NWZYBS
34xDjEWeOj102HhOpHtTKP/iDU/QI2VkQME+aJ61rUgOi5CNrwh2DtNvMVI4
9NwcwT8uNKoeUbHx6aXCLLtY2F4ypWQWn6VZ68WbquNl/IvPaR5N2p7bbk8y
GD9VwIN0hvESgrjW1vcoCbRCewdOkF9Ew/wqGOxiTn+hCer9YoREgggttg9w
xt/H4A6Wiuls3fvoelzVybhHNZ39DcA5Lioo4knFZFUOaqwKzY8ZqJ/xC3Vi
rbbQVhkn06sXMbuzX6/lQYWtjEi07l9rC0+za04m8FivAvgjzn3dUWq0YdSt
qAC6UXnXuouREZJ56Gee3hCXyRea3qqmtavPGRV4bcB92iWLlgcB/pb70/vg
58N+QLR8CW328y3paLpPoIUn3zQTKqULH5DnwTfn9yD7LgKnOGAoESoMdyRv
0IdgfAj7hase/5+sokmgBtdKdMNjBUvisxlxa6RSGZTmPd1rnKO3fT+E8QLh
0JjXuR0JTG+GW6PlKh0U1+4FvSzpP97Le+hETZ3N/2S4fgZ36luJl6ujSVn8
ZmwxDGB504jFqvPA/8nIrhuvnH08BQKT4LDDBjWzrpGwYigZm5j3RdkSVkM1
l6IkltjeC+eoMDpDB6tyMEKpgMz/5tJSpkaCBy81/yF5e5VdRyHo62VkE1rX
a7QFGRQWQn/TUF6DI30rvu8VAUK9Y8tP1loBc0BqUHawVet9gBIgcVpODzx+
iwmgRVCy/pBoVNNJHQslxlulzLJTKD6uA/M5Gw3S1dT6UWKRWlQgAA8kXfRt
qPArmhoDGhVXl8mKP+hvzGTLA8rPmQ+uASB9pYe+MOQ6EeDX9B66gBQmaVgU
seFqj8Nezowua89eOSPuFz9nYE3bSfsILR83WsrGwLeZcuV8Ja53kDfk0Vtx
33+Sd2BmfN2NcSeh5O/qUTp/OBhMwCa/3NQgq2f25cUKPPv8jgv3Owx5XvIk
wlX3OzRBmPEyuAum1Pbm7BPjfLP6GDtQWfm9hpznP9b40YY/RB8IL3jdF2s3
Zbr4tat6+XyBpYpDjvt4wwS/HT3ThwwqpJI2OXT+BIUT730OItAjfdYtsP5I
G+t/hnd37khFAUbMDy5BmnPWveZhZI+dk9z/ReW7HnxEq/g0vJbjJZTrAF3d
ZUw5NWwXduKu9ejvuGeQN3XhK2xeXqjcIi0R6iAb001X3lLb6QGdhc94VFSB
JH7LL853103bXDw6G9yppXWd7KEhnQI54kMeVmYLi4u9/45TDgLEmT0sasQu
sWw90d74QcxrUWKvwhJKTTmst4DsCKqjp63cB+7G0no6T/XQ5LaTKhy5CwGR
eGUw9shucMbrZScQuxxEhiGfj3P38IZevyqRzxHhKoun/FXKheDGKYAloPyi
3FSzAlzk0j3EPOoBpFU6mnBb1rUGx/k4NKMa+D2aKzhKhmHbbUyqPZy8Z2ye
d6oNQNMZiBuwfxYBtp2xYAAS7OZVGq41X3u/N5DG425Dz4Fzw171ZhFmcrFJ
JafhzlLbT0rbZS5zmC4V1WCw9jlQFjz6Tdce5vK+N+acTnPFKNgPRcipb8OL
cD+WB+YmLkQ7dbIq9F4dcUGuguFvxLM7RDpej6p784nXHIRvhqmEojglkX/o
rPvpLXr4J+xsWLO5JQFRlx2GBhvg8T5HlDi3TDBFBP0ofBaIyet6JkqdXWTt
fZPFRCYqpeZxTvKWlWycCWRmvxw6Xd7mNt9C33ZUotblCI69UxExnL342tXb
kzzLcAMayAz/8l+jVv3O+G5187bzNXxMNxQPKJbjEMXU77BGiAC1Gb+5JhDL
EEA8a488oRyYBVqapaJlqZ9CchUmlRvaPdudj3CsVHsoqzrkz4EQ1MqCRh8h
CugZIf0hsV8qNqMpkJI6Sq1tQRMIGTjncgt+bFAndZy6NR41G4u6vZJ1fTCt
8A7AdbbbSMRY1i+IGyNAbOtfC6l7M9VuIzS6TmbDrEAvhFKpu1uVZjLtkd6A
Ee6QqGQ5EgLyfSzc0SoIiteWtEUXw7/Sm7nhF22zysf/f1pzzL3SYmRZd9WZ
DzktmcSbjKNmSOw6E+UdCgOXTRn67hD/cYUkkWx97o2HWqTRKnnMUw1DWd+n
MiEIdofdrbCDqgDQSPVBrap1sf6M9OeSFo/DpSmHnqR3W09UtqgwUA94Fti6
agsvFYfqd3QFMv2Qh0naIks1hYMptO9Pxuo1yBqQxApyWncamiiQDTR9iN5w
GtlwhmUYHOa/H6tick/G1uQz/dY2e0HYxcAoC9ICmcOH02bUSXs/Bgqs1zmD
FHQYDA0JDhh/cWvYLN55qRmH4Uo+6SS+b0S8mnk23F10c8BzmeqPT38xqsti
dT/6PejGGlUOQWxMkmXSZiYZcWB7t9AVv/VP/NwCJcgu73/T2/hxxSPwueBW
BMeBf1qpQi/bTHTzgNUzCMIfaTRA+9aS8D0lmweHHlAyHwqWuG29CJlfx7vx
7oTKvLCFLy7aMwm0ZyoR21ly1Vi2A8WyaqzAGhHu1u687O4szhU2f+bOnewa
Bqa2uXsarQy1AHuvg19Bb+YyCH4pJcjsjOD2Tx3ufWm57YUrWDFV0/HSD5qv
RY+1R9nGlT/dWeFFU2evv/GEBm6mYKbfgDVupRJucMKedvvvCSn8lGBhFc6G
Aaa+WWH2p+GDkFqZZ++EcXI9iC7gmdcQVEyHYyRDfd+BdaY7I2WIdor983Mg
ln/tVn87RDUZPgQ07PfKprA1Wj9cNEt4+06DdLpgfEzw1cHE9LAoYzrel5UD
osO9AcGPTg3lNGA2eZHXImw31Y4GXr0Uw/K+G2JvjVVu9SLMN8g4eGCItxwA
XvVBPJuS5/wZAfiCpw6kAy5Bj2XQwn6tLfINbDR+OCQJ3YLNdpUpUcqLzqB2
05mzAemBe94UH0RkY5LBcTylX2EFaqIjAjsf/WYgPyYySDpCi50fzp+X4ktX
uJOvEU5usNHFcW6kSDauOlxdvsCJ1Fok8iiCIBmliCu243189zkugpafkdi0
UIr1FIpHBugYdtkWgAQCI8VK17sNHoP+pVuQeuRDIF5A6ZPK2WEpDCDayqTi
7oqkkzc58Y6qna35A9UxrryP0A8h9GvWtN1AFt3e9D0AlvEyRJydPyldny+C
YpNwdDPnku+Q32huDsGH6m3rNsSTwt0z9AfzYer8ZLqBudNWsNa7n+B4T+pD
iioIe38lt4l7Zj071B9NIShnb3TGRCOy3q2GHItni1Z2lm/4VA0Np7d22woi
BzA9+oBCF7qVrmCwPYUB8SlAqY4XtKOPEOX8vqLxbyQ/ZspvrmWjbI/kKP1T
ZCqNTSSxlh3Cxgv9duvQnP2uUR7vRyrgalmL1dLBymczOevfm7hixkFcQZxC
LeVUITmhxlJTEtMfrnTFqaHodYGflsjWLrE1ztAMo5eKgtuFbqz7JZNyUtn4
MBnh3QrnoSLPefT++GLDQhWXn9gE4PdiTf4eF01mfU50b2ZaJdvgPj7Giy8I
58sqrmjn5PuKkl3r1OAo/6lbBlq4zpQp77/k8AwswMpCRfqrFKv60GNyHJ5Q
vmvkchdKyVV1y+boETtatM8nvvnB7SF6zs60SEU7PTocqJtKyCsMNmwemqZl
2wwsOd9qQj4EvtGGixH5el3PT3uNrZqbcdew0JHf/sqOcXx0rpQe+uWWs2bd
bxArXM5FR3RRXhdM70scXeTKcDdS7ulRkqjypth0XAZodcbP2J2c6VKVQYqa
Tv97v0yVRyY3Td4HYUQVKkLvWdeha/I/0134i6anvgEiOX9cRT1h6kvSwVBH
lDkcUL4Zzl6Tn9NfqmJhj9cr4icS5rcb/WsGl3bPpQQELdIsuJJ9ub7j/aD4
imlC9x1SmZEK72P4AJfla776z9Lop90RRtSvzOKZXLWQZaqV0ejc4mbBdrP2
oLUSaI01TdH4NzZFn004w99rUb9/HYvvbCCyfl7rKGuDR9t6AsSKtAFuy7Ay
QNReqb9XFbn+4tvZ8AxbloYwkmcJ5LcPp1mPTKFbct/oJOIY0lQko2h9hQ5/
C5UpxZzsMs92uKG/fQs5+J9bJ/E77W2OJCFvFcWXM5RCW+2mD0yAg8zonapV
U9c0As07FNJsISpPKQYVkhFtg1lp9kk4VbnPkrz3Rb8fO3Siqe7rKf9TKufQ
XP6G/AS7nt/69VGlT8AmGse2zAO55nvGnqQo6XY/q++KuHZ0iu53/d2QtYYF
XS6rUy6OnE/YQNOJsuznyJgwt/UT8mUlYu5NHRrUa3sr5MvB9Rtu7S0Pxmmx
k9E6o09Aua79oqGEapWx/kcfetc/8fXPbKyzMLoTUgAeFwiuIt74vqqeUNjM
O76Q2hQdMO5r2IeFgIIEAocLihQ8SDbPKm6LlseGaXxoI1lN4yiNOQuJB7ii
ZbkhvJcmNOVPdsi1Lyc6LIvqDAU11fJhhTtaiihjbuNF0QaOS8pT+IrXqL7H
DETZpGfC6t6wKp90edeDlQ4BHG6GRo5CVZIJYS4TtIkmvfYPtPFEsSJhddXV
9DROCUNtL+3ZHkzbbZtxXTCYMVGXcmfDkGeJE/mMlvMeQt61h0tVo5yTJ1h0
4g5iAZffYLenzjvTlOMYbpIck/zwgQm5Ti5EgMaWVXHq4dSjQwE3QrpkDIfu
9q7UlsNKcVtucJdjYif8U4zgw5u10QD3lfs3fEdWdf6GxE2igyaLlBKwksfB
nDc83RvJjnLsJntjslddZH8djfJ23pmczzvPCbKSkfkhJUVthzzpbfVqb27S
Te7AjtV976k3MsNKUT9oS0VWJY/Z1yqovfychukIKANfG4h6jQE02Pqc2Qwq
WoF++G7nAAKxQb1dY3S8ldvGOzfOZsesjeu3SPdcyM/+lVvVl+vsQc9wUZ1w
fiDE2oUsW+Cqtb2YWSqnRh3KNhOy/0FAFq/lYLa75lrYwR1NjZWEhPIB9uz1
8TeyZauFCN6F3D71JL7JcyTXKPdBXLK3anLTrDicC2QmMQayz763jcKbl9hR
Ob0NegTXbPM79s+x7o3+FMBAhaaPPPMAzunZWQC3ACYCTuEidfqrxCeobUhs
2TOPOqIDwlj3Dnd1psyL5CHbMQ1uTREvA5R6TPm/3ZVej7qcq8qpcG55ztG6
2sPgGxMlKtN9ZA/y7bwsZC9dMqky86242C21XpkKSMVCpw3HgqKvUB3df3Jy
ErB5YYoluAQu4tdNojjKeLsvVOIi10G4YdTf1k5Q1NqcQNGofIHxEa8AQEeX
nDBstrNdOmdfC4s7l/NMaUyv1rHLN9E0ZtiqT1mnjM1J+hiS72BGg99I+1DC
oPvfRJ0ntBR4vTwc/XaNa4pEDe4jjZhA9S1R/A6mYYNF1TS7oZs13h7adWky
uQcTyqUpPByKe8GUeS2meIzbM/5xyCeORokkp3t4hhUus1GX1FVKHTuK2FGV
VZDulSHSOhubnSckDVp/8TD/2wYnr1OQ0wuzJgYXExyvuQwX9iFowCGynezL
T4hcbPMYTQtcE3ZJ128c9UUqfaTt3DoEBHdoUQwXPTamCQXqoH3gK1WAPL2L
AKqERlBaAta38W87O4+WLdOVoe7aFVpn8qT2N8Plg2iClmR2m6G6LKoQvNGL
8oSHJZIsTgNfoHITNoiR/OZ/lnX+40MOVAXBSF22GzGvic63Z322Qqfb9SUR
hT4aT6IQ6dbNg9kmvlcpHbTKgYhPNnQ2EwBxWC60X0fDKAKf5+6QNNsAicbU
s0SusHYEPdSWh9p3e1pHqDbygjdwUBN3U2M7gx+eKiXgpzwURBHxplCgRRNe
yAMGP9dkubBb/4vLxAFCBZWRi6z5oxx0PEjIol/CK5S7MrlPljsK3eeegKwa
mdfONCiaDigb19ZahhfrZhi9A8pp/NGLiHMee+Kr8LlNPOt6qL6oSq4DaIEI
aELYdgWWYSjaDQxCNUiHyQ1ieYf8NiDEgYDcOQ9+h1kyxreOz3mMvueP1b+T
Wxiivtl4LZpujhNZZaJy/Shtp6hK23DC6bz3M883ZBRdjMNBojhRiu+Difm3
aTD1M8psEL6+EBXnY0gX5D6T8wP/DDGEIDWFJQTPueUILN9VfAN4qvSUyx7B
0hg3HPJLfyZV5mARoQYx4HF6+MjIDAyHzc2tzCi1Zn3L1iDQc3853nSEeiJR
F+/xDYoekMCcCBt+NsoeLL4WRZA3hfdgnavyupzMNzp6RWhipge3A1b8yiAp
NUovpSs3dN4E6tlipLD5i1rBUiY0E3BbjzMXOYPMWbsztAnfQvglFB1JFFCI
WxNNGJeFD6BmFZD+tBAU4+YH3/z48OYzCRDDoUlBAMc6XgcessvqYDF6YR8R
DhSle16vGhfOhGiHXJhLDVDfbw/2fHgTooilh8EKmlR+qPHzacLKaQfQhRJl
LCSGYq6KM1a2MwIJaZjIBQW/SzUHfjSTzRi5EgESR11Eve/ujN/Kd9hD7aCR
RjutJ7eLaflNEKEMJqAmxXe48tU2j7yCqCGXMtT9riaErztyukoXLaBVxvYq
t+wq15bauE2BRmWg2PB0L+MieefY62FrvodN+IW098zaQ7gVwmSHNAJMLzwy
g63gTnJ8Y+axhbpzmaLhPqZmNx2WbrFuX+YtbFEE0gUZvMkmeges6h3wIwHk
k7TO5ayNkDGKE5yZqmbVbeDGXs3tyyTw/K3c/xYnc+kjIr2jkEOk+eqxPxOF
SL2j+RoB1KymnaPx66v2beY9c/JwXANTYwhgtCDhnMj/N5oaWwDRYUMH3X4L
N1enekAtEQY2bNcoBV//M77a5FUBsV4j/VWIY/D4ap7sbQzgOQXRHQaF0zZH
5ogWkXgRDyrgL/ziRsvUVyTKiFWNd/fNMtMoimUKuFhJJvD56EtJHQTPl4Vv
QXfIjoSSaiqkJEOtCj9WG+C1Tk0yuj4EC828by06uybbkFfI1vyC/ulyTM3s
cmMJKHWQyT0jcF90pxRLVukJFzEQUHoflqWDyJeCBYfeDe2InFMjJUhtljI2
O6MiBaeIpHBOHoD6bOT5G+DgvrWP2dDEUn0IbpPkFcyjN8+sBzyUJh5bIkzr
pRmCFaws8pN/KGM0mXza9OKeVi/NyRR/csWZE+EAZ9CM+5URFIODtyCecpzJ
De6dVv4mQeBU2uBY0POWx4yGjnJlpscLuxtfwdIIL0lECWv2DSj5Bwy40qk5
V+3L9ykbUg7DyYXN3/nLzUZuW1CGmTJh04f+cfIB8rGmW985cwJmj2z0MWYs
KlZtt9hdWrzoyd7ZtXI3e+iAVJi4OT1e2ETBzK5txCDRq9I2/O6OHMurhR5B
341l2kWhfuarnTQqCCg328KaMMzxPIYRNQQbzjPYMjhs6JT5a6iPpJ1JGRY/
mlyycFUqTzY2jBdqZdyY0U4nni5UKt5o/3Qd4VtIrbDgK0FxPZ1AVpiqZw41
xXuTCNY+mg7YZUpdVNjEuW1Ja7IRp8I7ddmnu4p5RePSmf/D6CW67xB6C9o3
KnY/YjXkoR8b0gitXnBGVQ+bg3sljb07w/VIN7WlsyBdrih8uzh5bkkJOP+E
kFumeOyjptj3bV6VbjodsoKCq+Tx3pkWdseqK7MVUAFnoRPXYFQj3bO/9Paz
jq2B9jqLtx7xY8rCOkmDV2myXX9CILGS1718iVoUJL4QzTsmzg698KG1jAe5
I+xK0Tyk23ca+4n11s7jnLMuNS/suURbVgz6hzsBhVqKI5FDWYeEoKhz+1rS
zdF+P0U/x5JsuPKqlx4axEsm0DiswGCfBWl9OLTAYaJzJL6+3tiwjWvoCpaG
1rxR6G4oYiw0Entk0x76IDPN5V8vPGt7h87MuEEzBGALCgYn9bvwyyBWmHUc
9PePIXh0puu/HM6JCq6kCncSCfbXBKVUHBPdG3QstzJjvYC0/uU2i6tCCbuL
/+mdAgcuIckDlmBDsIKcMmmOr15dCyP7fApSl48CQIxlRRbWoNn000SxpxMC
Fgq4EPJTrxhoaMSvEyFO00iUxyo4+WpCA9ngs8LaoOnUkiDrQrA8v3uL1e8O
2WBS8bE8FXYnz0WidRhy6QutRj33KyXOlwEY76/Dr3bnYNUy26YlpdK1taUs
io7P3JsuQY1k+uWnXhN2obf6E0kTUrBNFkFo4fOmWwfYhWDz/EpGQUJpFhRs
bsfmyIwWkFS9IFvUrNEYng1j+4paS/z7SBrAfrN2GDe03CytHr08/vhJXcot
LaYPhCI7kw11rV09Amdubv0CKrNQ2wqog7UWFMp64HESBARMDrBPF+CUsguN
OL+0hDav6xaT2u/2DUqI60iF456jufxT7sVO/pH2L/BPQ0brEkhYU+TM5lXT
lIF9ivgJbpqEBsmXGORtgVyElPWXrevuTfxgrVETU3kHgX2S436h1OE1KLKL
oQSEjHF9tv0qG6YF1DbBd30yIaRTQnBPMYDvbg9IV3P3RLbqZfcWXaZuwGw1
QIUPjoyka6Rfu/pY7QTiNQw1VPGiK1Wup9PJuoNXW/JsN2CvhlauXC/1nQKV
IvtLf/NCQIKYcWQdUw7DzGvJ3Hf2JS0D/+WPd7ermRkVYJBWDH82WrZTYXD7
kTKFF/HUTyqxSQVytsTUgdS5Oy8o6n+tWEOZLGja0ySBk8lPD/q8+lNOI4ot
kZ1HOuoS16R8U1tGKEvqdLC+Qi6LAFry+ehbr2kfsm0u5Ndcp686PUbUuFYb
+IojFtrwzcWih2YF8SG/46S/N4BDYfi+AO9WqY2vF7esBb4x712WPDgGZGQl
ZSYoq7GMPt8XMipfcL+HNlYNVMFlSC7Y1tTdQ3rr7cGSj7MBVQxQWWl3r8J6
tWuvdPLsjCmyL153gWRxzcP8SLvdUN4LDbxB58mypzkMHO/waXFupexwRSqx
BBWV0OI6hZQIBDnXlv9otd+IRY0Eg0jInmzrcjJyxUXsKiNq+GpnLkiHgIH0
rNluykWrufmXydT5qAWyFjJZaHN+Lgkm15jFPqYXEiS25qTgTNvIIdwvGplg
WFIz7EoIXtrs9sk3/qhbm+hcQWnAK/RfUSiN7cFc5VZY0gvktqJCPhrrJdvR
JXjnxwwR81DzByxMlVxzME/In+XRxdnG3GCFZFxB+xeepI2Vpraup1p07SY+
XT8mzukpMhkbMWbCu4n0gB9NkUMXeTyDS8KhW+ELCW4KWzxu3g38hDU9TsOz
RFi8MwpOdACXIvo+XANCLUCxYBBWkJf4zCsgCAy4kqGpTQoAoJcOSu4p9Ec2
4HrGJCswCQvjBAoBJdPmEG9CAGQ33zNHqfHQoVDZ2tH7l5wz22g97fsjMLMK
RhubComeo8xjKdv+UTSKZPxM85AoYI9+u8hnQhNHAyoi+8Mbzc6kLHCD8Bsa
4RxhQhvvZGhwycBR08H1lbJgRjkVBYE5uJ4iLJ21OqJocwvTNPxG2T08uHWQ
4StBA1tJXyEqbmDpQ6v9GQxxvmvyBXUA05LoFqtA4+cZZj2cyoEK+clygNif
8MMMmXY6Ml1L+J5pqRGf5KMNpdbKtxvdpIvWauPFjkGA9/D122h4H7KtYCum
XAhnLL3BdED7bOV1wbAWiHyCn0JMayBtZiE654pkOwtRjCHHS8n3jFhuQAQ9
Omgw/cFbPayhe+cizodOlp7uFYPB8dmFD/qKbAMSpUcCkEDkaHv0o58VWrBc
Dvvnebyu0YeWO2KaJ1UuPREXbB30A2PLUShtWPUC0z8ygojLm5GohDlITV2+
KYJ6nz4iPVWPPcn6pNqDnEocRQd7KNr7U4llsqBoVMLIOp3qxSunOeNp8Jq9
qi2KGMvSy8q7Ox9kAy/GPNoRh77QmRUvHwzKxtf9OY0TUYv85RmXstCYISct
E21bQyrDdpiJaIzYWg9h+FrVIMtfDGPgA04OUiCB2WqKvZUP36tzz6LrSQAu
bIrS2BzjZwcieDJq9HGFqGlefz4fSjEtPKUFlLsrr26WVydBkcFVsF2+KsGN
U5G+N1DWLpX45XCSd0bBB5PtSbbTd+Dvs37cpjcS5onCTBM6EAc9qGyR/eV+
XVdYeMrYNtdM65xQAQorqiEuk1DGZxKx1maDO2sqHqF928ASuKKE95Dtl6vi
24YueK2oD09HozQEDDOEBnwRuiNlbNQLUNpxZN5RpJFo7utjBgVGStMUp1ko
j9YhRLMM/LNbxSmodXsoi7gD/icezxw9a7HLeuPcWtcxTZyqiw+S+cfG09HW
HRt6IwNJuHaF7r83CEMGW6iDS6p5PL8T0XDSBxnvZiyd6lAeNpuaJ+B1zQV7
lDQ2S69TZvy5JZSrCiCWfaH96MXfsahIc2H3xmJa1dI2QzLrzpGms5U95yzS
pHDHWx+QCanlNP40foscC2+Da6AXw7ZSARPkEP/jwOsbb7RCp8y2UHyqlvyX
yKKJ9NNTw09eRfqh/ZwKA1kgDHX7lAT6+fd/IsMEmB9DqAFbHfP2U3ZjsyzM
b1qjs6c/tqEZUbkm9++VsUjCtOa3r7WwbEV2IGP/NireXvq5Gvz7Th14xFE6
MaQje8fZN9MUjo5NaxBgdbQF1t9cCTR3AmAsY1otd82fMw5qvizJajVJCJYT
2g8bsp4VbfAOsc59QMVmsBA+fGZqAcmI45hrq37FJp8K7qWHDxpVv5umCgo2
xGy/v0MEAtS0wGtrOQxqCske10jqZrhkizViUfsqZ2I4tOG6guaWgkzwAuGv
9Or5/X1wJeHP16jxgwdpcyvNzgHAiT/EUc1nJNuYYTt44rG3848c9yLkQaEs
mPKp9Egj5qZOpt02JfQgg0s7HIiFkr/FO6vw9TamlqxPB7F+dcd+dJjBlL3L
Xi5B4h/lBNpHkr194n28bn9wV18U28mVXi7N+Vu75arVPzJEGkZFzt1/xgxx
7dD9MolHw9EYj+4VYcGJU9lV8P9cTDPmwAR93A1Ro7G2tpMmi3890f5/eipK
v3T/o2Kyz765QFN83WEurmLyJ1823gm3KIX22IVVcDfKQLhj0Cx+UvKGCIs9
1ezzy7Ab/g7+IgG/6YSBwAym3fqHrqziEzsSStHque57hZJ8F32RXLtY+c7G
+RV8KcJxDuVp339A2q4uVJaf0aaF1Kjz60iTLj+0gqvssjHXJCZJkMIFZ9pY
OpjHrJ2+gNpfviT1eZZ5oyprWvQKwNZQovuGvlg9Hdrj72P3ABItqWjFoAgL
evACZvU0VJC02+OC0RDSVgXT42Kp5ynxEJujSmfxtu40NLGhCID02EdzDTsB
wVfSf3HRF17Qgbm41S7DBDlViHOoMdoyT2/U+diVqwqDkZ9E9fCtaKb0UX76
X9C8uWN35Vp7iuo8iwLqbKEqvNGRqg90M52MS0MqzYQx1nCn7gXcIXBmqHNX
Ruj0hVOoXtUx6hAw3m6B+1R+hmKdpRaFa8EJ04WUCUr8BnYd9QxcOLD0izM7
558lAOQW30CY0PgfEG9I4p4VFGUor/yLKMwtVW0jFBxvn5PpBt1/bnauRU47
2L6pb6skX0UZsNngMmPQqAlTjHgYAwRFsLFODNpqW/908x2CwSNLk0YdhAVc
KLCvtMWACT1FFoZjFFdR00QK5rTwPmaUZUzIDI7Cm88XClZf1wJSyK+FCH47
493VeMLHRmxqCXdmhviU5dZz1m1kakWw22ueEqvutVRJVEnNt7/EHvgVTPjz
5D2xyI61Aem5wbO58oMvYySV2XPhwdniCdX7xuemnn41DeA72/N+JNq4aClR
zHezXyOPoXKX4N9EvyodHPMc/tj3jKiVq5ZJnuW/ZiDSrucoMUzLokr47mlT
YvXM+SF9SBmrE2epTy0dmTFZyXqiM4TjFSTk6TSb/12iA1Xhn9Hl5E7WBQ9r
TCcJ/MCARQFFISqcfbf9KsG3+nI7U9YJ1K76/YOogqBt40kvLWlEs/aALLOv
7esthoFukGgPYr9AkJHEoaxWjJZiVbZXGSzYKBRVmj1Cw4cv3qepDizAWDIa
SPYdl6qWMkPvt++juyscq09PKZQLkrEEr6ErgbjQ1qp/ND3ztxcNReP821fE
D41IxrHjFMj5iXHUuSuRUY219nmf994JvfkFbSHymJ3ysXYQprVRtx9LLUNi
O8vxOidhgl9ta0af8yJoGQd8RWgRkiowu8aSAqnqRzg8klezueVwW0utHFI1
s4zaiRso3Kd34ZCgBmFW5Qm7qoRNNMKdRrUHR5LZYtv+u4MHCloifvy1XJyN
eiMjmuDuA+dgoFXxM0Q2T0JGiSGeUqZuiaXIfZfagEouiX6Kj5X6WuZ4Yb4E
HmJ6xCznpdDPjklDtjMsCnVVl7daVhYmyGtTBbfxdz2+LyrRShS3IoGge8+6
6SzJZlPN/5NHxx/vRQXoPcI8yPkBp61fmsIRAxKYL4GKiz6mrpfDELXkQjo1
qdMJl1CybzHrLaCl3DAANzn4XhlfrVW/VMdtJWK4RcnBr0AQ439NUwbiG1aq
lPLENmp1Vl1uFyjuxHsrgD3U8eu4Iv5k5x4SEmZKs942ARhZRfDk01jY/O+4
G/BFsUqJWLKsNYUkwRZuZAmP3B0/9eFbay5OkD0xRcLAL7fLqUxih16NhNIb
QADlrILxNPzfAbsVdAM+/h9c/3VD8YpFGs+/oDyha9kBEJPMEKAUcBbC5L+k
JhwuJM7a4DRJqh4fmlGS3LS30vA2IXgH/5iZ6nR+/1RVp65f0qe0j8Nv/+y7
55xwEb/7x49qW33fxkopPw+EOXWKYA9g0xYbdQ7ibAFrZrtTtpmCbzB2CtNG
z7wxi6mWLdwd0FAUBjLBtqOsIAhKCsz2JFoe3/wGvzsgMOfpvAwGKJgQQros
D3Awwvduq6eAZOatDCuDjNX+p6bGtt6JGCYFUjuNt5WERfe8LJy4dkhEhwCE
BM2DJ9Nm5vbOA7gFPATh2t5N4VDLsrK4WdKfBDDJJ13jPJ9C9QoNLXL/hum8
NERcLxFnR5jaUe0KcP/UXBMFt2gsABeOsfVBGk2JiZTRu9Vs+vwfGUWtXddN
/Ex8zBXJh+fy5t+Te52tpwvVN2CnbHp9fhsdIvuXql0YonnKcp6j4lfNt9XF
tv2723BvL6ZnHPs4SoTLdCeE0U8bVEcuduV9P64TILYMWvJMRWMWTayqvNm+
sXk3QKcNL7mpRGFLlmKrePR/pFTUnfKrAfzSZ97Hb1zGMyIcifN9vjj8ufPD
fDWWnCvaI2I+F4o8bbCA9FlTYyOcoCi4oz5iqZJ1mT4eWpmJCrT+dAnYJPLv
SiG7l/67tjRckIgZpEzv+8CcYPQC7PpTvA+G8rPgGPqvIXskMVxEB9KhpdeP
1NQZ2ii9s6SaCKwuyqh3vz6nDa7XzDqhPCQ0rsECQnRKN+43cgJYKOMXgOCd
7WiUsZenMVLxMAmm4FyQjmW6gwO1jy27oaxvExZbhRR45ksW78qWYEqGVYC/
sQRrJsCRRXeLzZp8VQCvpUKe+9t/psHwRwLGEw1NBgoDaSm2gwiv58OG7rSE
Y7gDlIBgOTkoV4EB9zgr1e6pr4mPFaKHbiRqpzJbvIiPrfnv9hmahhOJfht/
Xemte+6/VDG8I/yFZZcO3J/kLt7vTEfBxG5y8XIFq6eJYR9b8Lc7xQ61HeMU
Crtqw/ltYJiIN1NaL7tW97dx8OrnGUXiAG4fpL8ge+PIXdOxoeKHIZm17IOm
a6fS9DN8n7CHWARHC3rPWINh196r0hG+q6RcfkF7vbPkaUzQN8yyCFmoYl3Y
19FYH/4YinMJSRlbASn61nGCqz/Q+ozcE6lb+RKZFewTeD5zsqxSfZdGY3yT
72Ger30FMaDxJkFPqX64nzUC05FMk1Kx6tie8n4GLHPp2Wp+Q9I8M75K+gf8
2FLhqLi4ypZoH4g+D4JkVoGnorwcGLSHi4aBAMBuepwzuqJj6QztpHpVvJHL
fXWazSV/VvlbdQ7U6mH5mXgEHT3ONq+3KEnXb/heXWThktlku7ZelobkhJ0z
/tZcejUVAJnqqlRA9ufUNWHFndkbPh/GW9fF6QMEDaMAmJDtl8XFP/VJlUTM
y301ykQMaIq9X4o8Njzpv2SAagyzaeOiaQaXoKMdiruY1Yhf8M1UeeeE6TYk
oqy7zb42QJS+eCtvQthU3xQvnQt5zj/TQRbNyxCNes0s52Rw6TFq3I1PJ52a
B59sXrKaq3xHD8Q/65sNmk0c7Rbgho4Fi9Dhg/kJjOEzCr6SlmElaojEcMEI
1AX5Xfgvy3TvknoZhd7MM6PWaNASLT9dAkaY/yRCIJfAfaSKVXL0vHOa3dTs
R1o3wHRLPozIeEC+Ko7nTXGtZZ2irSSzSJ6ySXLMnh4HU3FMp08621ZUZmo1
RNENf5rMF/nTcdSgyj649orIp0ds6oHazIB8rp+HXIAM0yD7Tkr2SanNX6Uy
L4ft9ylB3/7sxg/cIdtu8VadkxzUKlxQxnkydMXPBEBgxoSixegMJdgPEtAA
FzypRviMFY96Nei5cjIJR9C3D46IU5P+pfs1ltNz9jmu9SYbm2Fwx7Ehtxbr
nzchG+1t+MUB1JoyZdOA9nrlyyRDjn5H0hdE5Yr3/fmgKkPR8MXrj8RVcyXy
BMhYqlzKvt8XYJFQouNvZMzssvJk6I/9ShZzVvlDuE0+q7482V9uIBD4uzAH
Gph7/AnQIBSoqR3NhC/MUpb396/VWzrZmZDGlwMM3vqnrNDcjJ8UTR9DoRcV
BWMrp24p2Joz+XivHank7s31s2FcZcaaFSt2lcL7Xw0aEEWU7rR/TnxGOJf0
DTXkElg1SbS1YhOOVTXjGxGzVA7oAtPKc7ZiGTX17R2VfTqfq9llQONa89rv
xV2qId7Zyb47wJZ0Dzm/iZ1QrVrDZcFl2OLNgkrChxovo1pOdCAE/xNmGe+n
JEL28oMe1/HcD8u7HDDQsYSccn/YDExdrk1J832ECZmaLV7lw1Cqzfoagoc5
Mv6IkQQgqTyCs3Cv4H58WwqQIQEcH15IlZDH27EAqA76XgbtnU7y+TCD8CbU
IYoMxralH7pVjiWbnDKx5Q8Vjh0qCM1WhWCAqi1QnDXfizLndXHiWZljlYam
p6Igjt66iYgJF78FjLBsjWxnjRmMx/NASltY5NatcfzjKvwp2lHo56gn2/0Y
BrucBU9o6ppzF3GU/kDYyBT8UvK6mVpVZGlhjDRLMrf08bFhIkqY+ztp1sBm
cQgiPOwhw4eunsV7l0tdpoFFYVXzwS59+ZME6ficdrMPQdKP5Oq5t3BSSVSn
ouJRceJaMG0HoqihIddZV5S2NN9XLYjc1GOSI+sI9DsHr2LsOZi8hD63Im3d
C7xqTklX6gC9zH4lafS/PYmOycm2DRSimbql26ZuT9yF8g9ts8vpc8sT2gzx
ljAf72q55iOrzngUjA8gQfjrlNB2hhE3VGiWIVkYTQdqRkHxZCKRYc/MXLLu
aLL7DrzEUmnAkuXIHOJ7qZbbXk7S/i8wmzpUpNtM1o0J+9KI4JiFaoXIddPh
CV2R72ku1blZvbpo2oddcDSbeKmvsUbpMJGBg6FyVWiIH6ZPYGT5lWGeM5Za
/NgOuzP/PQYxEeZq0ifdV0UK8MfEzMT+xU2AQ7naAsmuAPcnEYjAFmNJqVZP
1k/Fj9QxqxanjEKETOL4MlAuN/YsAsceMmZSJugVB5hulqCNX+CvnpQsIRjd
RJy5+T8p01Y8K0ih/xfz8Lpbkai8WUYTw2cPINX43aVcxwideZPaNNQkf1V2
Kd9JOmC3bxbG3kCMj/MJeQIQFwIUGMOYmPgAidw7M47IBVDpYpjxkazf+0GT
iv1hqpqWMOa7x0blFIjC7iC0SMBU3NqezGCUcAGQnkZgafjfyXkbK6NRge5i
qjqaXEf89WY5+Va7dqwVdVZ2B0sD5z9CGuSL151qaSu/nJPLvFqRwCSnmJHU
AuEicalZxipdCgd/Iiw7vhgsi11c3jFXrKgxhyLIjOQKI1OmcebhRVZ13umr
rlFOHp63keKP0jdKf36jWAzQyS87bqVcQ3q996LS82lrUOuz4at644BNvRK5
V7Je3ykwSJF0u/vxQbKDGT3kbv04qih2ziXMKo/7jebf1UIbURBdMMoIdbFu
YBlbtUVZ5rXyHb/r8Qi3VK2kyvLmCY85PfFKd8AqmwoBMhFTrjgJKSp5mwbi
wzpjYBpaR/B4/3ciMa3N3N4IRMxF3Jkux/aQ9LKF2qfw77Sgp9CUXcm1keVK
kGlFE09wxaSKiKBse7E+paBX5PlndCNcnHVbYc2YrPg9kNrUZjPree5gj+z1
ino8kRl7DCYEB+mJr8gVeALcyjZJESg3m068w6ICpAent9uP3WULC/+CKaUh
YRVaGMgoJM8GxySSX2jNFfcz63c+Gazb9D/F/2SYopUaxXQrNH87Y2teTmag
Z+POs3wb2dwq9aqvm4tSXdiaMGHQuwj653c8PeIiInUxNzNdJGMq3eqdOU5K
9Su94TBggk2mnbcScyNLUn1mDIoWrtvLns2zwue/4Ie03gULVOPSWFeVQ5FJ
/CKDI0841QRD+334eTznNz0KF/sztkFn3hjZOg3NklboUMwiTYKCMfZCNlTo
0BPI+SiyqzVxd4z5QV+xpm8ZP/TKfLKcGr6KHuUCmZMTtTjyxODEqu/T1XSQ
f9Dwd4RmXiJvxDqyi/kRreWEpX3kNJmYra3DuFGGbUfjejZpU/pQ3FbQwT4X
DzL1e4jWBIG/xqp6UFBY6vx9pPlhc0cTAptgnEPvPrJSwi9Ke+HN1Sa48s6q
mQhxGSG+IvIQeD75c5uK9Sjg13ZWNiJ6/R0fzDwuem81qfeQNAWphCasfWUe
+3Kayro2wetEnaGkliU3LTojuDMncyKsFMZ3Lr6QOlMLWS4JGpvjXkVpYJ87
TYrTspvRSFpl4AK2TsNOwO/n6YKF1Wtxad80kZyD77V4d7h22euVLUvPdixz
4aNy3c+Zb1T5QT/BO0rU6aKtgP/bN0cXSs4zmqH02DiNDoOLyr+E4rCA9akM
/qz/FM8IdBMd6wM3F+6/bebKm97hpMBZc20VFQie9MpD3b0aV93VzvEQuN7n
8VlUzpCHSAl3Qua7wv3kkiKOU2UzoFwJPZ5qaFPvDcESFNzld6eXorRkA9Ue
pEqAVSiib35f39NMtKopJdHbGVHkEJl0D1GonjkBjNj+hr0137/OEljsbppF
THObKooP/Av75kaLRRD6PwWOpOzDNFe0utkFoEMC2Yi3D4WnWafTv4zJU8Tx
52BUwrowyPmSrkCfxQNH6ma+Uhss7wT7LomArm8I5roCOqCeT8rYo9v1+90C
d+51Tz2VUb6h2SvomHmit9KeJam8/BWBuQF+2sYZoqOs9KqOygo7jBWvna3F
HX1687OkRZ1NOM5Pq3G58QkUUYQrMNwk4BwE+iLoQwDJg/alFoArlLr5fd8t
tmVFmhdmOdAHLx1HWOpt1BNGbYELgDD+GJL1SohHGj3qKOY1WqMSYH0iK7jN
n1+QFpP0HhxGOKzoQV/8LbwJAhfo58qjMwZgXI5b2svXeDs2Ohmtjf/WEyO/
v+q0ZnHlERSZ+SawmTVyRcQdOctXYhxjWVBVGDv/BnDr8sRCIYFE4RTsVO/P
sctnM/9pSXl5b6npPOZ/vC2FEiI63DS3lYW8nrlJdjL0Hk1LYb9MppdZnJPg
Fi4Rf0JQaagqgxrlzOjEjJARlKzPNoH8J58mNkQ86WiRzLFuIdX+hOLjCW7k
70FBrAS44DOff879VRpwmH+ZB0PK/R6QLEOlMVDDnIYf1h+UwVY6ZAYRQ4iL
No9VOIhOIRlAmR4cqNwJGkrCjn6E9K0uOO0ywWhKqJAcSoU8roC14OY9YSXG
4KPDQsXlase8WP9e0WemXVRu7Uxxi7or/jvKPqc8jsbHtRDrMT1/TAgZW0eV
AJOMBQcsXGEB4HoT2+DOiiRPJEDlIv4rGwtlQrfsslzYF7mMyIekQAojwjh7
32mSISQUu1uysvSr+K3B3zj0nvGbk/bwms6Lb35DUkM/x1YiyoIwmPfA+vXw
m95/apuT0pO2pQSDtQcyLmwqzr5SHlmH4ofFjKQmdxYzUzpKyeOkgKX1HBhZ
hsaJs1ebJy6LoVHWFAwQLu8dY6HLSDzXAC2/UET7sWbsV1L2pXXImpgcfuyS
r+UUkyGHKBKlh4bYUFWkjwjFCCNgdJjHwrJ2YgUgVhB5NNZEXIOi67rXyuso
6Q8O+uZgU1ViLzW9+1UQdS3/hdnxhLfkQe3uzfJ0X80/qqWkwb8XKMWb1Hsa
sei/KnNFVx3BCsvuNPenDkHgJ7+43seO4IHdssl0jsYaSd5cva6j13REnhAM
xgdcdYC4QUfaDiu8BmRInA53Ucbbh1vM1lQIoAwbC4HmolR6Y3s6ESOTvksr
mZCf1L9Lxer0RlTpfoJfxWRK88Ry+fq9WvqrndmTk3RLZ4FigI94B8TIrVav
HYIYOcvlZTz6TN1dZLAzHwYSZPOjLC9s0Admk7CIG9VjH/jgLkE9rp4BLnuy
Y3ukpRHJmciYHHuJHVX8dx7JAoETpAc0ojCZjM4BXuuNlsYk0NtVfLxznm0s
KC6i821ewBOr63HabenAI20tonBRuHnFmgjYTnDvquvB8Qsf9jCvSIOrL2js
fWKL63FCXm7Sr9UsfDLkgH9zfPO138AgWc1gEOLaQQN5TukYC9ctVIWx9rpa
/WztWUlFwS0ko1e2EhVnVvd07bNNxRyDsWI8NzyfYzLRKW0+qkD9rKYYL+xd
IEo69OZX+vEsZYr+iGwENOqwN1AJIs0Z9MnwWc4brNj6qI+DtxuHZHrPDx4f
Q337gh8vdCnS9icyZar+xrvYqPZpN5tMRIHTC6adI3lZqyJYxe6qHxUFGm7X
pDbeqtqHDRid+1zG/8Bve56ohpq8A9hQrrsXz91TXNdzrySmMJ84XO7IgfHT
zJBf3eBUPOn0yFS+11pIpU2bY0RwQtS0PFRUXaKjZBVEa59WAyw3qXRZ/s9Z
gdkNjK6zI3OQMVhfS9+v2guG/sWu5Jwf5wEzbb7ngr3RuLRRZTNxgSBAq32X
bPEmZEXDFUIEOzON9yq305DLLDxPX0zmshbaJspjXiSvRtgyMrCEHHKVDtlW
jLmnmOfzLDVcNbaHiwvWUqaz+hteS0PKN574Iqj1U1539qp3567jR9kut7Ri
3xQUdsF33suhpooMb4bQkCZI7YFvc9IgSo6RFACBiova9wGrH40QvJ2PFm/r
DxR1JDv/QlRxoyey4cNUkTGkhfI8DP5lfotE7nEZr2Fxu88OGFsL/AM1ycmo
5QK0iYY7kjYqAunQWKquOgS7JeTEO9MRYSsOZ2+JEZ6CPHtG7UHQXHEEV33b
BJVIYBFvvOzYYBGaZqwqmMurInQ7MtjJvwPQ8gh4MclOsSuEiqyzNLBCjdro
60aL3qjqIufSZs8ikoQVsN1ahaJmoOKF33/jAPK5pmtgbYXB8SqwriyDar2g
8E6+SilajwSyf0U1J4rupGVVdLy+Qp6AOMDuLPQK04f+j4qVMO3ZWkomX8HJ
S0Y8ph+KxowisJ7ZCsxAoQwlf95d97CcXbU348fX5Dt/ITsN9Nkxm+oql3w1
YmKxLjkdgtSDTGsKaxa52BaFDswN8R4ZwbzJjHVBM1GZiueMdGbU6x/mUjeQ
gvaCfq9kQ5HGM2moBrSW1aul4b5TXGQQ0sQ5s8BNytv7d49u7Q/ZK/vXgwQH
B8laXPI00uCO7rOYQ/YlwMw6XivBPb97nrggwpoONhkdBVv1scfDF5U9iwPc
cVU2em+SrfAcl8Jj/GZcgarieFLCNPA7Tel7Al2GoWKmefpWRvAAqq6bJpSP
Dq5APZ05C9eLLVlIv2x1s19wAnSpz4HrY1gG6k5HJONrjuYFbfPAdKANBJBM
vjV6sgGBLiTn0viXtHVaPv63oGdBWUWKU4oj/2XYOx/EtWA9Bg+qz55Huj6G
HK4kIspMCZMv3vNCIdynbnI3lOLEAyJ+PqNZNBHHgEY0bwx0Zgze2YYAMsjT
MN4YdgTFsxk05T0f1phDONZ2KLHhiUao5b5QRrQe0+kqHs0bOSrOlLT/Fz7b
q+7btuURgLS4GakKQWPWpiAaZFffIcXtnkLa0vBn5ZsyRk4vxyL6MG2Y+6ny
yl4mB5DAwO+VC/ibcwU0k/LnwTDUOwBzjOe7LrK5QyszOrzuO/2H6NYxs/tw
ox3+ah4LFAvqVk7WJQYoLLD4XzXMwi5RaI/HVllRCiOlBn8Z0KkBl5mlweQO
tYAkbfJqNw5F/8hLtGzNpXDw/LQxCFOOxiNWJ+BCduPhBDNTIYLDWCbsWIIh
9rMWfmYWpIZCTLG7bdFdLey7kbAbgHvLpVnclYehutGBUm9rf03w4ATq4lCb
iw+e9i3j8OdlNTZe+nG4XUO6746sXCI4ezd2E+wO10q5tiKFMni0UWSOXEPY
1yr9Ow1eb7xdqlk+3fR178cJIaaiNqrUvdlOUYRwYkPfSL6yYHSo0o3Z2E5H
Okv5rKfxDQVnn8+iTIpUUjsbM9swWRiRriDRAJS9GVeXNoTOeQ19nQ3fLY2z
Tr4FihBT0BQqOz5pyuRN5o1+LzMKbXk2Qknzls73UNp2/oTb0WW2sawU/xOw
/0bL/riWSa+5xKgZOw6vSm95gCK8xSbgveRTvjcJupb1MgEQycr+vTYv5q0H
QPNmKI4fhpvG0gyG8CdegtIvmHl8rtrhe1fKUda/KNmXsb/OesowV8A6qXba
JsU0yS0iQbcyfZV374WrmIim6gn3m2FRhlxvNMMbQfN4H3Op/Tw/ibY8wmZM
wWJukSesItcvIVJlBS6mo/qR/vPnlRLXqBnXDy/hOF2/gsCCGCvPP/UWRqr1
wTtC+LHPb5lRzuXxXOUTLbYlAdabsUZ4i/py3U7Swzjs8MHkS5Hd1wtRp2C+
grKyepyVjxtjOgQYptLkuRTZfE9rku0SDBGn52o6vdtxAzbpciYdMNF7q1no
+TMhjZgaDpQfrvIhRQznBwXDwSPF4DtIGoC8lhaCdfPj/05/Xi8JX+gsQREv
q8de5uGsXVtoqqSrBBwR9NMSjDAveQgKGznfAvtrmOpceVogKpOgy6f52yHd
Mr0ibFC0eHXmTR204MMBNozbXiMa9NefbhLhWjtGJC3jf5ulZjqXd5+G5UJ7
FQ+xMsDXM9hYd3bJ4cUQWHdm8EF/UKxvQfq31/1w482b53JCY4dLC5/8Qghl
5Kh7CxhsKxmOl095nI/msEFCZ/x+/r0aB2R4e+BcGMgE76k9BtX6THtjoL8d
m1fpFYfkaLwBqkgcSrnnCB8FGKybMocloQq9utIU5HDl8OcqQDBxlUZiEcCW
U+l1ekpHgl6aUHxAdn/mZVEG/kydgiTzlu4cRlg4AJadqcT7oopTk0Lh5Zcv
IEkV7tIX6UKyMIA5kDmLfoffmoi9RPYKE3Frqvf4led/BdzWL/ncWFLv7VHm
2Wc5epMBrlQwwGKACWR65HGzbk7qtsTvmunH1kJUI1v4L62iE4jelm2ZS1E1
jq3XsTTC4IHm3tvw9INGZ1WE0+L66hKP9qFClEHe5uQmS7KaJYknqVS6ujhY
Mke+85YEVNwMOUCTwoFhxXtoA3K9FTo640DO1hb20HD1Dycq7qThlaEQ3VcP
VwrvRNmFFoCphOEgu+79vdLJ+i4jrbDcgAJ04MqKKiKs2ahTHNo+jpWL58j/
44J3Di7cNG646V0/a246Vz01uujQQPiPIY0rx66LodAxuiTasGoXNu9vjiJy
CYJBJyGb1syJU4eulMdKOgERZUpOPlmdkxeuVAmtM+7Lc1kSQemZeXsd+s0X
4EJHIOoo3VijzPxAZFNhXMIDuE1HbSKicx26OL+oHqoUjrbgNWTny3iG50hp
bIlWzrCYcaqyP9O8X4X+v3o4CKCwDZDKUsB88S2HU50y5kRpgO1e0IEY01vi
NgWVAHi8qRF4iAGgZLaYOARWGLa9IDBmlWD0aqLr8QAU2aw56Lxgoi0tkwFY
AvLxXdJWn4PEE9GKE+RkAftPoqKNn+HcS3EYdJ5lpwswb1MlFDCzOZJ6/cBa
mt5RvsTfD6dZdUL/SI3otXqOEXkaMjT4kYjlwRS09f1s8xBSgJ1nn1BBYvM0
RBWr3KhvEKDt1UXnkB9/tkPuHAUpLSIhQ4YSTET/J6HDhRbPbpK4+0TvYvOr
tKonE2ZQinArEdmYX7bjY3uLIfB/Giqs+wxlg4cuq36t5Dyi6pnIQ7ckOjEm
JATh94Mdh7VjTWYRbZECBdS5uGPcEwFM4KqgKVby4AHOHfU25Urdp4uR1p/q
6cFsthB5jNnfmxuQ2pKK+5R1OLvkDMacOVDSiYN5G/61pIX/+6o5Hrb2+JsG
FvY348aHZ++pScD6nysHxP6IuAkrylRga7I5u9a2HQITO+dd1YB/WuwBveNO
yTo+58ekOHVleTh0MDayAlVR0D3iyW9o0ajwuLilpXepLWVjruyMKpd0sRqj
I37njANNx7Ju7F2mx9lHAsA5CYRyNyHpdLEu0DOj+jO7fETVYSY+tej0aiv5
4OGz07UzkLoNqmO1p1+RlkbsVf6RLC7C0b5ixnoZEMAkqT8cJT/Jc87Xg7/G
4zkCF+oGL4w5DP8vWexOqPUfDVvRpfnARUCfca6XJtFOcvZTaK/Vc0BHxKgD
DGjKncIDdlG9vsSr9+MWA2C5ACxBmNYHWnfoPucE1XDGFS9UyMHYLcJJTp+j
ikdIYPwgIrqCk6oQSEqqm3PhEcLVhoVN8AAHK4nRIBkGfjpcP1/X2tIEZn19
daKkrJPkG6C3/Rz5nJYWYfyKY8NE19SCt5lEt1GkN5XaSsYjIAnRMQR5j3/M
TUoBwFjoWsu1n3/skXiNieWHDq9/w5ZVoxKWE7ZdLc6nSnz/U4xFTYdoBYp8
9qpWJ1/N1EEdSY3BNyEWwutWNNgCkUjndNpQRECeeuo+86lL3vSXMxLinnC+
LvBw9iTc4rYf711dxS+l5HlwpwoKhAEp74EtsUbqoLcezDQo4BzaezCSoJS9
7n15XC9HWefmn5QUjtyIqFWd7QgontMIJQPWovcH/HkPLH+6a241eX4f82ul
4fzp/e2Dc+4Aj+WZm8GhpDhi3u+Yv3K8Gji88G5VdQjtwyI9Kwbbmsz3UB/w
loT/k4bdlnALBShFklm5XnmsG0K1fEpBjlrLxSRur11JAe0Yk2pTwAz4JECZ
xJD4Q7lPUKs9rGRkJAanifCwf/RUv63jjB/14smC2v5MTT/ukMJxHxzxz0IJ
QpgT7YDS4s5LlWacFvBBGU0nXlYHkURa6fL1sJX6BIwX+76sLLpZevdneGZv
Za9xfDTB+EVnIXFkx45M1DAeFvWHZgKeR3cGyBpAHljqRClTMJhQDQgekgmU
DXtg4WG+7Pe+N3Gp9ZLp8y5FgPribHNfEehjNxK6wSvTx0ZDV6dI+mOsECIQ
RC/mrt0FFoJmc9KWsxZLTQuOYdXfCg6+gTwgHT3nh1qubTwxtG+EDBVoQtFt
n0k8wGEk1P0Z1bgxZOfuO2udm3Ew/nxp6yrAw1OAtUTPEswL7W7prqcXuPpI
0lVzxFkW1tec1WG13Vpk2WFR3M/JqzP+WNRZNvzVaYmZLt9U/TFmLKF7sJrq
GfZirsPJs2yvBVr5+3DnN5r3lJQTtV1oEhZFUXkoJMpn0b9+OchQyxQr2xWf
TdFhipCUobfxlXKou9SrEiVEmT5ZdNi+tdJ7a4oT8uquVg/YxJ/cfiMFdkQ8
iBlxd6Qstlr4gNTrbOxYx7+PsUxBUuL2wHVBPZXQdmGPTJDPv/u4SPBn+RQo
6RyWdfKLsgCmNYLLiNVwJ5+nn5CMbeWlqsHtNxvhbxvLnX9kBUkIlO/AIHk6
4fu++TMZ7ns1QFhjY/JdUiAQdwwjUuSZptLP5SATN0GnEPI9uvbEK3xLIGCQ
BnS7cUucePToihjksFsIsUBSQCrBZ342CoNrulmg6KsxgZrAeuYSB+2+9J9j
QYBNLvy8l7Q8OEF4v3dCdmgPvprNXbMDpnspx1SAD/lG3YtxrwVtSx5hjDCq
PY5plnkLnZpzJa4wn3fu/KGWQtBcTaS6Pbwh9yqPIXvW/uzhwArv6pknvIMQ
8zXYHwsIEzEG8nYCEW6vttoGr7iphd/9Y1xu8oRunY+ACmBSuIw5Shl8T7lC
gyETlf7Cm9Q1QPNLJ77R1G1tF2CGv/ljo+0DWkrwTP31yAQb8U+iyP6V0F6V
D64EYKg5mI7bzuLV/1unkCotykXiunwi/EDCkhZ5Y61vyjPu0BNqQxF96FWC
vvJGVAsWvVMIwepoCDAZJWf25sV+IXghmUiHsJPL0wMszLdJglYn/ACO+8bG
QFUp0kB5YWZ650koOYIcVO+etFFM9Nqg5s+gkTo6bXKfAkaRmQonAcfBGXKz
rPNiMonr3pxBU1VkSqEr3723Nxr+LRBg3BrBW7eSGat9hS8c1zSj44ITQScR
GLyKitqTz5dOb4hCXbKUj34IE2EmPRUDBl9zNtxM3DFVQF+0jF5lVTrbTFH0
/qhPRE3Mq1bx3OGcl/QAIepiZyk/7FDUjrgDqB3HHWe7PqhOm2t8q7mnyYY7
KHRAAm0WwT+JvfIuBqoKIFyQOaXuQtl3QobPcF5+mnoHCHydcalEcitJYu7D
CkM3Cbk4Vwzm9WfccSz/OBMf0FH+dpJZUoHxSe9tz8yOFxKxEFAFWWcJ+125
RRXWM9Tpop2mdLBXfXZpOIW1b4POnak3b9Sgi6wIM1L7VeiZKFSvDlvC5fa/
rKolJNrWMfVjwgPBkfOaQFzuH/ievZZBFjX4V9W9mcEr6rkwo5Kmk7tTnqLQ
oLvkJ46bQI3Y2doH1ebpJ/9KrEUcQQuZe3vYzeCfTLH3A5HT/RTAIwHCFZ3f
25p9PL8tcE9eOZzygNI8Y8GoilWxGKo01Y0wAGGOPyX7KgmBuYWkvkANpWwG
4Xz1AmyQ5EqyKzh8MSfqizGuOggHKPxMbwxQmUZhH9PtRD43IUAxEJuVPqPX
NwWMjLh1M0d7CK5jUewdW/W8EHNuy3guCvLJpTnNFrt4cJnnmz7o0S3OpdZI
ZirEb5ccw/t02fkb1nrSJ3t6LFlmmUVV8cl1eVp0wSUgYf/PLIP47G/lGQ0v
a7uvfQl6h3NSfD6Jq0NYzHN4yrwkKlOglflILQ6qV8cdWyaj4pASOIONj+XE
ct03g0UA1X5+T1T8k696JSYSwFuHx4hOypfsihDVTOHIU/gD93Ezik4leaEV
QAvdeTU/m2KHnLQ/VmcZz9xBcMuKsmQDKejR7ViL8Mxyln5CtUJ27vf+UoZa
mTKdQc8jC18Sb6MPliIxthdIjB2+lCzeBze50vZ943zcm4Opa2/zW35Ac0yf
y0FNmYJxEn3UqZkNSDqTGYKFnTpr/BuHgcIDXZhOYS8ECRXBwH695LZliXXa
+edHA/KxM8zP5QNN8w0KKMe3GQ/vERKhA+jvqh8/iCLgTpL80qln99nr+8Ih
yyV+caukAfaa0kQmETp93nl4v7Qfr7kwrMgvN0qSdoHVLIg3loobic71sWCw
AUu7arcPFi0ZjLH70ZswBzVjtWaoQ06AEtiaOQYorNNk9/bE3UdHyvU3x+wE
30jeOKR54YXv4e0bKA7Fe1irzU7T6E0qrnLlx8CkVC321aENo2NZq/jPSKsa
h177wJYQ4te49cs0QlNbSIxLCtlNqLfzw6ENfkL8RYX0qp54cqCUaeBEUPKi
8wuiNA8HG0Z0eUadJ8Yc3nnCsBi2zQbNWGEEcSy5dSBkATrKO3oBmYxfqJqM
G5isTcb5bQbj2mXhE6mIMYs3CBnqX39bgG0HqsLwPAof921tbjxnp8TDCc3T
feI4KPTeBe1o8cTP/5GDUv8GcQrYoJ+c6x369JWkLdFSkfNlMsQr37m5mn4u
IdJo4TkuQc3hYB8uRRKkFacD8cktmkAX9lBCXDMqsvi8aGQ/CuFkEulAFkOt
C2mYu8QwJ7vgTdTxaUEzHnjb9GWNQEfPkiFOczerxQ8ywpUZEafECCl+F0oi
8p+Tl0YGti2KO6wRb5c+0RG5WOlMEfC0gbRwlh93+DK9NNVI2/hXkWFtZPHV
VkyVIAcJYwRj8TX1jToKfA1Oce/WYnVXDrWds4zWLfGQ9qsim7gzEi5NFlVp
x0iZAwoSrcszJZEnURjc5VvmAUzRIqzVY2uQMTsSD9sHX2izg5W5o1dvWaCw
KBtg/x9WOiaIsCiQ7LWA0Ncl15ObgMxHZlFJk7FMZoShgVp+7hLPFfdbqElw
/KJpcMogA8HbTt1Ql15Jh9Lzi5h7HJ8kOzs2Qe5TB2Bf/UJcsV9t+NouN2S4
I7HsiUUTCjLfpcDpaSTNHigRt0RL1oQRl6lxGTwHpjg7i1uxNGovw95cdsZU
Z8AStFCJIAhLjXDaw1iteojQWbxNWKC+YhK8vK+XFtDbKoEYYQbZP7kqdIsu
snJQtRAzWlYrfpyJlUty48eYJVTXesRImGJuGs+tI/tCPmiSDiXs00Zy/Nyx
/U2Z9gXjq3xdzpvFHLrpTdATEVhMnqX18NuKynh3fjOMjH4O7cBEVjFMMUW9
OQVrgAzFdWzD/b7a7WrMf4URCNr2KoFw1lsk0Vf+zmj0xrfbKdb0Ldu4TZSA
5pNfCuKlXNvD8qnKkjAB20Tn34FdiF6wiUm+7DiKkzLPd5LUkI6Wrvp1QQai
ib6jQHTIDLE1VvIbWDphOLLNy/fib0DSvAGIJNlSFnATG8PhTUdWV1NAGP9d
c8r3Pf+QVsV4rvFoFHTxytWHnI8tW36HFa9E9oR6xrbJ4C0Qj8pdamGpj2hM
jtMI/Mg18JulXsXAkq2BFE4lPb9LdktOJ1J3C4LM4s97sR6veB/Cr2G0x6cU
8i0ynYZeYp+2cjKerw4qvd9GX/HJvPqUbd7pyZ+GUnnbjw7LIK6yp4ISXH4l
IhS7+riSRbpi6rFElIymBcwCtH9jVBKp4SrBmNk1Ahn77vikDVsVa5iBIfYv
WFr2oe6XVYum5Om6aT+YEVaBa8b0rc1VLuOUXBS9WrVbiVSptc0pyvt/sUTq
55d4lVQGjwLwJvR5itLDV9GG8gpGEMEBDxnnq87/JPGo8givR/+Q2vDkYkP/
OhojHEYPOxMEOptEXZ7Ebo6ku9WzGEDSCSJ/g1BwIJ7svev1EEckUcSXptxP
peLoxfGvdT3h5ACp6qW0Flf3mwIuAN/GNELq7MWsdNH01wAsB/7JJulaBIkE
iEG/ONWajKws6cM7IIIxL63CHPJVHL6jAuLSld0fELEhFN6VdywhaOgopamL
1nCeNC59hcP5g+4jfagqSnE4sFDaR4PYgAbPnCMhoqkoz3m6P0iSR0+ysamY
8HpvayOUUBps36g0Bv86fLlajiu9jIIGzkqTIilrpRqFY4rLBt732toLXq3J
URRqAPvnDgB8n0iVttxnA8Plie0HpbfXVk7Jzg0+IcfZWc+Je0jTUa3Ww1OK
4Bq1Ivz7luvSNLtsp1KM2kXCvbrCweuutJHJtGsFL3ZQ2ZEmFS726DVPud5l
lkIvb/3dRXf4dbLb9RCRIeLHvyz3hAz+VFp5f/3YSSPEFmszjKFa9vFrcIWQ
LRBr0gjvh6BdysHpwQj3O4tu5Ie302FXYOSJNmRtutI7IifGJveuaWt0Q0oV
/cfoF4g9QDFp0ZlozH/od8rbMVgr8/RnXeQMwz1fCIX1gPAkV/kQKeYWJm3I
n6UZW5BJrBfJHfGy5nEudu6jw3MqKjYC8k36+6wl+Nu3c9hJ7p3xmucKiJtT
oNHiWgKLqMh8pySdGsn6Eu+c0U1YuWrB5s/jtmyYtbMv8qPB60kq4DcHyIyI
XOF64oAThU+1x1V84P1LouLtED89QBhqS+VCKMDaW+wy0s+EvihvRJpFqoY9
6eKf3kBbl4Q8l+TUN/Il8cZ1uDcFbAWiGXXWED2Ijdkr56/PunXG03+Al3wG
GA0SotOQrxpk+o0nvCKhiHkKHNatKxw1du7RfuOKyiZkrJYUS2tbzUEnm4gh
5RHFDAMR1ecFuabRzfb47ZMZS58kQJno9BQ+CMLTjvKGk+SVtCYu9LkIHlxT
l+17QL8uyAinvLcH9c2UgKwo4NU3q1DtA7at44gfnHSSi3F033yVHcf/8g2V
1R20lZ5ICVR/sL4CI/LxThmNKmbohWdxiWxRh58JyRsgCX1AFBQLkI/zkJ7m
sZpBOTTbbvsZt313uXQR0p9Mz/gEwbockVpKg0UDYDxNwk6pikkrfP2XQ2sb
7tVh+3eBy2xN/EAHsBGOaUnmZEQfgEkDKZlO7lgxL0U1vkFpkwaTdhRIcBsM
44N2ogdHKBs4SMZWwuxldbUU7D30hHsHV6TnFTUx8YskgISSR8Y+59g10BCb
TFbUmSK9KyrC5FM+kk7XFCcdp/RKW+ISXNkT9uJm0bXc7XoOI4teFsMfOhFF
EvgzBI0IqCxULOHlLkbVcXi2KO98lgUKQ0CBAQjLouOjqqooD94dFWydW8TU
U+Fzkb4xhGwa2lUwa4EeR26ev1f/cee7EKwwmeDL9T++j2ol3dc7Z/zwB0h2
faxt1weO47/RbBFMZji+d2vo04d5jG5X1/JAjdefzSPDxF8/cB59/SpjFFzx
ykiwhU6/4iJ/cIk5q8ynMFDS9HlOjfBYGoEcd1ODDGCsbGghBtqwsYuZ8jAc
/uvKqI0Li6wOtP1xfrDB5++Ttq+TpBzr43xB2KHSiHOdP7EKpox3b0HnVPyZ
nhpTR10EioDP4uV6x60eFjNO1OSM5HxrJMocvFf/JI2spkiXDpycC02ipdEN
LcZ8+kab8KYVJ+DVyucXSABefc0eaUdmNNPI0/R93mcIBzZ2RffUV1bL5Yl6
NsM79MvOUo2coucXWclRXTXupqb2PkAvU50naEB535mDogD4x8nf+4F6hXLk
jjHQlHwvER/ryB3S0PFqh9dLcw21s/h6cixxxZGDfkDbHdeAXZmVF9SxQwVw
9WyHD5UxFMWCWq0R0m7RGsrYSBZjxabKdaB2CcTm2A4Ieq3L92pCDmXP2cBm
T6sTmUo7sKFj9penjuh44YMY+7sFhG397QSOf8A6NUVqPsCc7i8a7R1MwqCq
9mn/vQq+6m5kPieHK81N08ZOXcPl/wEOq3EaC8QrwhMfU+95a80uJf6GYTaN
vVeQLhXvqh+xY1XInWdO/CIxu3mGuTMupgPnCo5hEBrZ3XZPAjqKJ1C5ZbEV
si5Rmg6ZcqpGr+1fvk25EkO8+1/JUM8fFVDZiBgshtXvysWshpX8roUvNTao
WRdrkyqj4nPeHLpMBT2Wu0LJkaaq2jQwNiyau4Dg2ftFlTZdYA6WdQuJX9wM
8NMAbdQMsFNqiCY47LdRQXCe+i8hlEGZSLWnoom1ZHZi+5bIzY1izZ2X06jF
uPtXceEKpOIdhH7hiPvTi5jnGPeRk6MviFRrxamU02i8fnIH75hJOHKHXsM0
hCR4ixt9PLr0YoIy3IC24ZlyDivEISbqIlqvUQnrMLlu0PwJCBR9sxKjAQbk
BQoi6cVepOZM1khhsHTA2e99pWSP89CqngixWP06xLBvZ3KHJCl0MWN99bps
w0GATggEdLBxF0HreIKozZD/oq2x/f4twjP8oQd9qtIsLkmufHGEHW0ohqdl
IlhLyTn8EX07PxcVVx7Vd28uguoCggvh/F2de6kiB4tAKh2BWN8FLR0r3Xvh
QovAPP0X3hlC0AEWo0SgsbbzKXKhlnkf4BI78uPWO4bYVbwrkikvBm8NdaIq
JuYDsSAOHlLsf1o/2Hqh6Pqr4QALGPS4Te5FVAGnmOvpgnrp2tLgLJEAIxYq
aHmvGhvnmh+0S4zSoWRnbB63vn8k2IRw+iDQ+3CqTQpINgZmHl35ay6INV6B
uEtHv+zZmYyJTjN5PuJ5dEQzGnfBINym2IbGZcnkSvqguYYp4ghqQX/XM9sr
Z01e/cHxenwC2FeuKbGC8HpMOu6KOWBhsMLUkKFR5ofn8/iDces8Y7zGixSs
tdeAqH8ulI2RP2WUEarLPNysAFcivfzWVBF/fad26uMefXdK0d/vZyv1VJZf
31aTYzxqYbSnYb6t8MvHrojz3iWVR7iusOJz/ZgTQHThj/1WTZFvr+GWVlye
m3t7fl9X5a5G+61YnQbNm0EQ/fIUKU+cYbrn/z0/5DsFaSkdLFzuMclIATha
5QiXQEJzWjxsE/IN1FkCFQpCgvIPCsvMMvskzYTnsNGTlgF7YixUZt69h2Yt
itvaqnGT3XNHQBKizsjfq26Vxna1lJDzOVGZ+Td7doxuh1KQb+WRct5mWH6I
r5QG6DWBl0r5fR5/GJnl6KpkwVCKdaLllfoH2hrd9mT/ETFjRNTifU7b3bCb
sB1HWQIfPkn32Dj18wbWtq1VIHQMVQk76CWQlXRr2Gyx8q74cv97yOxdhb9W
61NZmwBPoWZW0GwWCQ7D8yAK2SudEwkwQDrdSazovXjHWFcyZOIWF2cVfe5b
4YJNWIaoSh6ysF31xgKKIxmqfztT4WS/2wTvIRG/xe5xZUj7ipsJ84EN7yW7
xX9GKAN73p5+lL/8WbXfJ7lgpeeYkmXxf2IoTU7yTyYtdsqUUEHeP33P8HEE
9ZwSCZI1+Nkc6feiPgphJjZ7DuX5EyzoTbI/y3EmiMG6j81A7AHJ9dyMnlLw
gZ82sXUbj1tDne2RZNtpnK1TRnMktNGU13VNdnmurumbrqmIVVdr9w1Z/NGJ
KZHCF3yLGQEos0QVxlS7lfLd3klWLSbgjszv2jiR0K8RRhmwl7uiMBnhNNyy
zpN45lfffp/vyQUwBRuAoapamdCdnc5JtD+pv5+jWvUnJ05b7FnkHRPxBND2
61E+kclW5rwHGVUSbJbIntjgqTCbUiFM2l6NPCx1esTHEXB/SHQSaWNbLWFA
RlXZ6BgdP+2KzR4F5sdPWY4QvgWtTwxITd1C5vM/A8OPG9XMn06TZOri+coI
phYwTR/PDyfczcr9W6eQgMz+JVrfm0JEgEd2Wws31eCVedcDDe+HOx+v0kRq
oYHqU964PidYTZI7X8BIfl/V23t3p/Nz8U8I5OtqrclXsVKddNbrlu14NYIo
Jqn31ZRw7deQv7xM8c4WRr1TC9TuJQmkSVAQiyRcIzuDVFBKr0vmb45Q33Fq
31qBn94NPS+bMlBR9at84WV/k+cufqwHxxcCvY9Ssd2eQwY4Xhz4jH3kOzXi
f8lzVIiBzDvRng8RmHDVmsetOQcMVwuxvnpGTdzuFhTfQUFrKJTP7p4PpjQj
DS1+KOr4/gRj9WP5Rq6KfSqZIEPhdIMn9rCEjfUwE9CtR1KoK4F7ayadtu5p
PPNF/smo5ATI/EcH4S6ZfMKKgIXcNeVc226h+WbwAds1BAWYzbOg+6vabEHN
vHTJnTgGyIR5KeU5ydpQ2Z9vm3RhOiuciOGZIXLH0Pop87oTVsJE8icfuUDW
J5H/MlabPbWNLMEM+TL0VeoFq8Dgieny0BOQxYC0TUusywO8+bHbOSYGQwiP
rj6adi7fiwNmtVecV6wGjI2w4lVKinfO9Nx98koK1FCXt+4L1PUKVbfVsYcV
sQmA39KykYU+a+oo934Fz72D44BxmS9TqWC0PY3Ln/9t179BAV7zxEM0XKae
Mt2LICSgeGcOM2y+dLHfi/AaExlGCC5WL2sJEXAT2fwLweUR22srxWm7h9C0
1st8XasWRkt7GwUwb/BsC+neCcMv53+b3BAH/YVojwMV3kPaY10+0492kIsY
k+/RWfMtn835gY4ACeMP2QkpIWX/d0WamQ5vCmlADZDRQHUHYxofT0bgdHSq
Ayug2889lLoAbSZJCsKw45nKdekGRVxpiQHC6QPB3AbmrMb4jAc3It5uVvyA
SsS0LC/NX2ayEM4rXXDgBAvM4yZwPW8KKcMd5+y/L40pMAnLx9oBcvqa4aaU
r/Fz6TZwG2OZXQnJBbLYub6v1oiM25j2gn0rwSuuuv6dg037h3s99HLHwAYj
b1IHKiW0eltfy0y5xa53Q/mTQPnqCz/sayLDNMxEFE+Wfs5Na37kisHJtkOg
gS1fCuUD++K6YGyyB5oC7pVozH2aWJl9lZKDzU15U388A4Df8AJ2cmR2QZqv
ZInokIMXMk8NgTZDvQwntpbF0NNV3oFw9mXL1/jVmE3bVp49NuCIzoc/H2An
f0XmQ60p7QXgDS4nJmRmI0WUlgnh65flFkaaN2tPRs8zhRLyr9WE++AFvdN3
5C+yPiaA0Llv+ZFBm3Xgc1mpWwF3r1f1NfDkA7ap9tnQH2M/qLe7UXX3EQwt
XHRZhP6jI0inEaT5BOxTq9cGGevf0qrnFwN9xhYIs1ANDfaGOp6tgiaauQrD
eASZtXuYTzYNoukWxliCycTtmt0g0X/uTtjqLkQBJbNPVbZkWHyZ6I4QvPEJ
yiNavzGjokRjCrQPq58N+3wjweEFCGbiso1hFO5ZXKFk5ij4gzX58BW6dchY
fL/5GDxFKRBUe8bns/sQJW6cO94WoAMqwO8/Ua6RnBztd7emMy7hSIkN3zrr
4s4S48xIJ3Yh6cK1Rp1BZyOvWET6ZmU66GpoYguH5W+J3k40TmhSGfmoOF85
un6RZKILxXNJZBy2PW+r4HF5txc0CJknHUUfQiUgK672EB8V41tB0b2cj59y
7IEn8c3uwTE9eeYObxjJDuLu7+e75m5Nm3QGHvN81Ku50a83g6hm/9RXLjGi
KDx42x17bWqaCT2+oPsB1ND5bif5BQWw/afc1EpwmebMXWlzhC1WMkHrF4GF
NWOYcVdXquwkvIasbujoxeGgcvYP3KzNZK1MK+OQenS4j8aEtWE+frVNfWfW
C2FCuYTzef4KXiuDvHog+8DG4fBi0fi80pFTF8oLK2rZ5QfZcGQChFqDGb9Y
jPjuhDV/36HNxaCByh/YVew/j3TrqaAE66vdQl40GHD1kaihBGPZhAooWBH1
mdZSkfdpKbsPZBb15Q7jXN5ys11NazcAnKOu/8YfwAGgkOgsm3IVYOX4H8vU
o7rUr1osLCR0Z4eJt+2G4Bz2tJ2Y8Vcix6WOHxKuxx1txWcTVf1IbZiozKHJ
qwFF8Pqn4whkz2CxTTbX8/3CaATnyKbw4WHC/TPqNqTyzBIHOaBwiojT4T/2
j0Lajdi7qNiej+B/Q0xVhvEWuxCgCLD5shjBtdSukAZNrRlOTHNqBJc4Y2F5
GPJlPKlKOzAZ1NhcrsykbLmisn43r08G94gBG3y3GM5cBJjg6xxzzOEVRxR8
Wl0w0g4ZputFhHk1TZlgDGjh8Eqe4ChN8EN8AXtLuT6MN6KtV13P1V5WhUZ3
XzP5WOoAbHDKgQVbEZXw52qE9FcfOTCg3R9CW7vva+5XsjbdPEDgFAIdXuaQ
s8OqWp7LfUtR28J3P0sUS/hI0fglHK1GMc9gIjZj1dSxhxugHTVDGSLWv5uU
585xGmObrlTwtbv7Pe4LOIqXKOerPrQ94qVheAnM/pYHgldzKAxLKBQq7tD3
AcYFIunkKhmCuxUSnlgZBR/gB0olPeWvqTOz1JdRQxo3UV2eks4IrohurAfO
DfAxZ4JmFQC33uJl7H7rDolfFMOFIemjWKsJF1I/MSn3ct+GxnqGWR01OGCa
PJ/jR7TzyvxhkrAIRgJEMu/vaEKZOUWsGwS4CasPznWxLtFMqePHYjCsdVhy
/aFue45VQGGUrEd1oUQrygrxm70B0BsTcT2QN++WomVFNEM/cBXNw3JpQ+PQ
GmjL81YvRnyyv8rUJrQBAiSVRitiu7nGZcux6DVhHb7QzfT5KJRg+epoMAQf
GEhr432gqBw01Zel1NjBWYkGtVYTUvAT/1DJI2KqU0zc3XDN81uCABUNOMWE
dMXxMbYyno1Ypqnk+X1YtF0xuVlhYHJhQBza4cFDnMsr1zWfn7p02iwX7Yf0
NS+t3DluKlNPtt7nZDmN7AYBRHf3ZJvQLjCXkv3NsNSlo39JTXTuTewqfutR
CPOitOPvdXnAp8p1nU8Z0z+8rgEwz+k7flC0+7gRKTZohXSLMmJ1QFNZOX+n
L7UEesv6fXKWqWx8WsXl/NPHOpMLzhRlE/fJ2eeNPv4zw1zAE0B8wao+I2js
T+gHs1JKXu3lozOW9300dmE4HQOdghrAz+AvjLKigIDO4B7x9gygQ62V26p9
hjcAJ4r5TrteSCndr0r+S6AXtpf6lORgj24m5YNOpyyI78VVwvEIy01kzT8Z
H0TlCu8Wzi6zwe9gLSvjlGnBj9HBpl1WMuHnOR/l2ZBlgMTUheOif4gLSaD1
I9DuaqWSmlg7YOKyEXL0BPrgvOVmu6u6OIUzr0lW+6XBPw2gB074g5dHEf2c
ia3MMBP+tXTcTZPGmq7jJiRiqwsdrDfLOwZ4l4JAxy4CFonj9YOHNC5192yp
EMxC5K1uDiy/humEsac628nrgku07zsJ+as7hQYtKNpLtYY7ylleuuAAosh+
FcjeN1WqLRGOHzgnlDa7DiHeV/3cHoXA1b9dAxwpRCv1yxyt0fUtC9VRq5tW
ZIQzrMjGIWSWD/wQpVl5fQY/9k9scl+SUYJuX1YvHlQxFNSb5/B0VcllP3wl
+imxgjY1lQ80efHEdsJtpxKnCrmVFO/lB29q15fZ889lilNg5oAQXrpxI0W9
/K3q/bDytVgrHgwqDkLkv6I5jpnCQPdVGdiRRKOsLBZd8Ic0J2BjK6FbTkzU
ur6tL4KbfFXT29luDkjbIfqWOYS1/xxETiP4qW8Na9YbHvTuvwYEggCNpANO
qxUP6gkRNPl+zXeFHsDTnV0i5BzZsqsHasrbNKCqSstNmNBdofy5aGfDkNhJ
JFHhYN4XEYx/kV5aUp51NpzAMN9uOzbXv6jnKicp7/x53eEywOZVRbOsJKKe
FuTalpmS0WrWd/b6Rs6SxBBycPnMOTvQQN3d8tZi269owLjvq0I1oURcJc9x
ELvBjML93hG7lFZdyTwh8S6J9sYWhnsBSN/74cx4UaejwfRTrNJVdXuU8Bwh
qu45sO/TxYs/PtitbCBpDJw4GtbPyWp6RI8AZONtJnAjXFzPCw/CUWtH89Uh
dJWz8Z4yxmOL7CijAs+2ldHLp0cJ2xBHyqSoBCxRoOKjwA8pCJvhOzyZy6ER
ezDiigZrHh8ztBPgVTcPPRxvzJ7Td/oyaetdALn+GdILyaDaD1Sh+OFePNSl
w1QcTVZDs0VpmYltc/EeSbiPDKZk1DaoIVQS10JSSqHkLGardpA1jbBEeydc
TGylg4euMjGjj9xzxVgfjLeW0YRNgIEHXJccLnZX+qYs9iQZRKXkg0oCsqjR
5sDXZffwn7fUQvSOIJhV+PwiXt9k84LbxvwxzKUZuyalZ9x9sDvooK1Ef+yO
rNy/qWLQbFbfAhU0QvV1Wc+FKUnMeh7TVjuuHeztjpZ+r+D9BHbFMXTRM2ce
CKHHMmYAKLegvJ2Vv/fU7z+D6HCI+RJ+Si+GOznjNRJVWSe8jG4DswzrKdp/
5M/UdmfWRyxlyBpDGLkcJpa/T6N/nd6bwS356qii1Mk4nyvnSZML7Qe6tuJd
4HUdstbhS1BF1G4GVw/XaaKQibFKb/+pviDQkQ0+dCKRF2R3rM8ML8lVewE/
LnmyqiLV88WMGKNxPxz5Lyh2XUILv7dUbIdezbCg8X4wQuctnp2RkdC6Ba/d
xX/Nam1PFSqJYh59nMAUSVQyf7nmc410/NaJ3oijYuIokcD668th04wOrDL8
T/STxcmlRJQscu3RFbPcmaanuWLl7M+f6/0gDybX0dMFwkOI/CKB1uGJ0PNz
UQmBKB1sxBxxM0qH+WtZ0tSJO+Gngi5SNebUFeN471mAM2TVwNLZDDG1eWB2
mK5SZSP/9LnUiQyWIkD261KasFRbR7Owu4mnuPSSECktvrpHgsOdKbw72BmN
c/B1l03UV7+m5PjCM61jm3iTN9Hi2QvgtP+nXoQQ395NTEzEh13kYH61WOaV
dusOOAQnFbdiHqYUeerC6pLOlChi0ZTgqGS6V7uDisnx/CTXJhWOcdKH0aOK
kmJnKJkjgZYteUpyYj6mZjkWvai7TpXeeAp0jass05aTh37xP/QRF0+4rbsA
wYgX1VN52noI2/sRxZbRA4BJOm1KobGLyXhFtTPzjdXfqhGz2scLVkMfVAur
zOSB7anISIdL/FEQv9/28ZDJgzcMdXiAO4kphZQ/1iYIpvf+P6WEzwtRs/g5
LVj9Z6d3EpdaEMleqZEwb8u+S4JwuMrEDLzGwZH/XIs2rFtRmQ9PMM6KV7k8
u5OPFIhUqtzFtrrPVoKYUyFtRHiuWevuP4nbBLLVmimdWr14tvj17UH0aptm
IYht3/jBIOeY7xsdo4B7y1h2wxgIN0nICEERlWKK/uj8eWkSTPiSKgUXafzI
NkzoszN1Z5skDuiYcr4YT+SU3I8IpjuzygJgMCs4hh0P/fMBtkysgP0UUjib
tzK/YrxwexC1DJCzE8tkqqDQjSVvCevKZtSuAAC8tZNDL0HFVK369e+77qfs
dMNIhUaP6xlZLWYZ/HSg5ggLLSIpPdZh81UR/DBDbZ3q7xoQprzw7jOLbntL
5PpUOuPRQzprIFn7UPaQSudm6v7jlChnX8Dtl6ubF2/zYlwz+5jKcF7yex+V
xdOWdqrFFJMdF95tvWGKUh7gw4fruqz1bBB8MUYnu9M5r+pZxWuUfJ9xayk7
opOIt93GXiI4bK86HoL9/JGqgnpFtowRY6Yvq5A124+M+mFC2yYJBnQPYBAq
ZLYpoB+UsPaPkE+DC82daEfEMTrI2l+Hz6rsrP8l1kJrimJzTQzo6AJXlr0i
iC3kaQbLRBI4C5JhGT8YVjX7ARV+cUCYcuLNyiFKW9GcmnqGGQgbUCwH/Dmm
+rEetEuT2DEg7/BioomztE5+WHSXwImrfnbAHo/LGyhgWqNEb6YExE4HxdqZ
tODMIHG2ySeVBl3lVL8jEAfqVRM/6YA8f4ujLJmCmW1LPsZLbz6k676sxd2E
IxFmWqBs5SGTTJnskuBxgqNccrPA9AINbvwz2QK3dGba/kbZ5SoeN3r1p5Sh
IOAQXxSfEsBS+noQxCUVecuN4SnUrec72AaLXuEwewPiLqX53biRmbvp4a0N
qtw9WIMaK1QpTjxgK+3Z4yalOisuFbcfI2Gr+vgPJ4DYSLJs/w4/RY8rVnEM
tewZFfNzAkaXa1Dx0quKp0xYgDEuAOZX2d33uvk/ruyvxPe3F40ne+92XbYZ
xobXf0cjCI3DJHBwATpyp8Oh4yS4BrpG8wriErYbIdczVt/NUFoCNLJ5ZhKu
DkW2c20ybE+B+CImMbP8Oq9qmmIQfbFx5Try90z5q4XHjJazu5MvsZx8n0vO
EW3T53/0e+RM70mP95LbLrhvPZb6anPYUG36y1LpwBC4IBqI+/tYx81h/237
H/EkjfhFeOQ6WOlQbU5b5QoB1Jz2v4X0HyfI3CC2t6jCHUUEe4VOIt2Dcvga
6E+7wG8jhUoKyxwxj63st3qLepY5+rhEUvqJ2OnHCfWVk4EXunSVRdfDEhox
qqR2jb4xDQGDmpMnMnN18P21B9IQutWGgld4Z3nqRfr/fxRKW3q/qQO8iUFd
evFaRoO1E6ATvKzMYPnRjvlvAgqHp7RRu8KZSJRDpgt4Ua8gG8mhcfR45rHW
20ccFoAmFToFnBmwPdqT+/nPuN2PRF+I0WKDnzuDXROrIFGpXnQO/9ppQpEm
EAsWGwIjFfn1USqurZCBn0D1GiY4BFmHkXLI0RfUV5RHeZ6nUNMFqnl1i2pW
IIo1+//DWaLYyntv1XzawPvFVQKJZnJo6z7FGKhPi0QJ/0KEYPg8q7qMXwvI
dpcrctQUUO7Ms0VePYlitM9qSWAgJal1KMWdy7iwX5iZnTpnS3uEEB9+lSU2
gnGwIV80iucLDByM2n3BALIvYjh7uhiLy5Bql8f6K6mup/D1O88RhPvvpxnJ
zMPVK0Zh+0yFtxaJ0J5JtqZMASOIg85Rk5fTTFoffGPT9uDwxAeTzqVbi7vj
8jgIR3lwhH8gyLFt6oM0x3EzptdlJMoS5ehqQr8cWWcomu97QWNZqQDV9lMr
Xmie35q9ecJLYfV1KhnBtoUCxw4LxDzQKZH1yV8Tp0LLcuYgIu+4fvuivd62
Ogtyt0xxWXkx2Pzdsk493vwoUPL6Y8YgNCXECiHbZkVp8xA3+B5zrHVDheDm
I8m4X+UbclVHMr8y0slvmT7JW34cNwfqitFvbrJPm7kI2zuh8N1VciuRI8ll
c34O0R5bU4aPXpH95G+NyJc4nP4xQOxcaIhFb3xSPdLpZJ16bQTpgsLBLw2e
AO+HqT0lc2AterQt7uDHbEuPH2/qA8tQWk6qcILDgXfXV1QY7aDn65Q6l4W3
w1PVHXPFNKakUEcsAtjuON+10G1hhnfHIntSfvB6YPJaXTU63opCMZdTunSR
0e9of7xlIwhppKd0zXroRDBh6t2TU4f0bYn1+IeYDmCiswjmGVK83QIi9Dmq
YEfGsf4wpg7QlIiSYOx7HGsWY5wGuW376qtGIok1Ga9vQW9BQq8Op+PgSVjT
lpy3WTTFT+4rARmFOd5peXsurjDhZWY9YCpNEWYdi372VGoNYPBSflggQhLq
aYohAusp3fV/p2v1TTp3w/zF7uXr+g5AC9jJB78anhy6Snbe1tLiEmg0xjvG
4RBmZB/gWUJ4PVXpn7AoMpXv59t4scI9OYzLoUFip90emEtNByOYZJVm7DPx
HieCgbVCW6xrArdHPxec9EyfHIvAoIQjf6LXx/oFBVrV0xsEnPe0GvWOkQnS
oTqUk46mJwjpYIWAIdOGYi8QId0lV5e32QoRTiyMOi5vGRjkLu5BycOV63PA
gw0GMZaw5dJh6DMzCws2vBmxy5KvkbVKvNJdsPAJjjrda5Eh530UVaWgkwAG
LFX9NMzqFNtFbEAgxcebeDOXWe6zX3YBeWf5m66udKHPa9KzH/c2etxI16LK
11Qq4pJzWIgSiT6gwldIc9H9agEhTfPR8FAUvpGT5xrq35c5NUGjs4jzkL6F
REpyAdwZJKU7NFIwxunSmfN0EouVKunZskidq31NpQOLRf6wFzBPCFGDXJ2W
vwtwvK8h8XBH1Lo0lMf4hOYk5equTnwZWl4C+1K291C6Ua6rDLi99rVD+Lj4
n/I0E1RVOOfDwFZzP7loC2k9rwa7+S7YKsUhTFfJtgVgGctqlW/HkcNObhKV
LWsVpEE16MMQKv/tsZcrAUpEEIbZ42KV89+hjAawewgcEG0VEm1Sk2JIHPJ+
n7i5WFJlhvd56AJ2+zOvIFx+y0jy+VznuhXOCb2sHQBrN4wd3/MQLogOhUrX
S1pFgTK7nNc8kX7/c/bqk5OE7Z3nYcgMmbXjUIDJbLmearTbYT3YjE/NsgVA
0u8Herchm8cL2yL2mn5Y+9u1sHR2BsQZKvrysUs02Z6ig0Ib9lcnik62pdgH
VXGmBePSF//KD51OqGiMpi0FfWlAci3PcaQxiPCg57nvCGqAiQ3iC1w0wrLx
HYAmXfgYrCCKHujun+NZjSbPGfR282VSqQjAlgfIroA0HzF7AMCZMy2TrvFf
VhTN8YlrOsaqmiprDbV/IHwJUnnnUZa2Baa0XmzTrest9WwWsVgYSqTV2uyu
cuSg0h0Q3b18hwmHNgFZuTA/2vRUrUGDOF4+nMHfYHfXeMgXOgWsrQ9gBSrI
4nIgVQgdvjxDmc7fW8j2cQaXHTnWQ68/J+BGC4esLgImTjkm4wj5npPNFFDF
vrcHGwoLrx9YLW3+Fke017FkSE3fdPUt6nOkjr1FsFWsrT7OVESrahf/uNM8
982tCJYBJnXRhjobpAmCgjkIwl9zRb7Bxshv/Dc/hmILINPQEHQutZnuHJay
8yWZ1/zvJhcaFQRQ/fNinc7Pw3f1vaMS9sEYf1fkDE4+KYin7YR1wXPlShb1
PCvAKWDWaXuArjKCVgd4ESvN4+Vw3rtT0+ESp4nqi51eJiqR2kFmV49NphST
NqQ//B14rtmVgPsY6QDHM0MCapdgOdy3ABaY59kzCG/fsSoJM9AYwUV0RIQA
5SLZeANMb63+1AUqVQvmzYEm/uNG8LDQ+5QrYvcvM8QiclUzbderpCRS9vnS
VVKSGf/8k9ptAhGZq28EsCWWvAZ7ZdKrYHbcs0LVmkmg198pyx2r+ShJdAh8
k7mld++/xJQJxTd2hDrjIZLqDxmrokNplYaS/o7v64AE7O8coZ28RSAjB0Uy
IdXPWQWCXGI/j3fEI25KtSJFOQYoFVu5UzAuuvSPNBndlkJP2o0AmqduzIAF
UHUpN2VtLBDYrJjTZv9LrjbMQGiXOw1HcOUTk25uR6SeNQk1CQXFT88RPlDP
IYDRrTUqaaQqAGwHR7MhUoQVJ4PHqlhUckB0STD6nesQCHHbrUviAaWJrFOu
S0SELWyE2rb34QHA7KisYgICHlJUMfX5LdztLz+orm8I+fp5aAMg2vo0I6HP
1frMZ/7e6ngoNhM5Gf5d8NwRRoB/zmEcZ/w9h1uE82wm5UXEcZLpqbDR63it
jLFCMPi0GdJCXfesvrOX/5Oosy3jZLsVD1ZHztOAj2U2zIh6v9RjKO5vt+i6
i7oG7CWDkkaLlOFBNF9fE50cSV0obQb21iTVnV02l9sM/YFJFaGAxuadh9Fo
Hv++Fr2Csw6u5zok3owmVh3BUcZyuPa3HyKZ8miR2Zdwynrx1lgjUhTndTxV
FBoe/xvVb+AnrOwRgmwZfz6tk5yJzAGnRgtoB4nzbAJbOOKNNokyCJHZR4tO
o7sowLTlFYPvk0fY9d8AJoW7owJN3SCNxj2V/XNkSoqnKXeJ9TW2ewVXHOw6
B/y0xnkv7xzcVGI8cN1Klp70blv72XEYL45qw2jfdAIKIt+EgG2p7hLbLqZ6
Ixk7fSjTo0blWDnoqgjby1rO8KIuN8HcjbGVJGFXB0AuY5Qx4S29gJiB+NON
Puz/Cespa7xyOO6NQ7limEkIv6XdSl614QUwBU433i2MKpKBjuwCip+iROCP
B7RVwscQwom71wdLD4y91VsLgIZffxqmrQk4qPHlBmQsu9rUKJcpLwzI9kDc
RfEp+Hck4OD3D570Ni4u7HXyu3AZlFNgOTEJlwhAXILWYChnpuCMpj2jO+y3
P5Qr4SDai5qqK695YqdbiB06Am/PXQ/ml60ntuek4hXXV3DJEzvJPHolPMAR
DRxCw9758fZ+KKAA/94oVlcP0W1yCwzSsESeNIcJkAqMZzJci/vCwu4n6K0s
QMJIXaZzeuCMafBRfwvc+1+Yp2RffrWMqcJ1pmd2Ap1YncVlOBk1J0VZKGHo
kWXj77xPTNNIMndU07gP+3kPogIH8uVasu9gA8en6ICfdKVVihJZ9tovA0iS
1e1h87/niUUTDta+rlNHwnsne46NS0I7V1cbSfxqsRRpRtIyyIt0AGHeoK/c
DfJr/n/YHoRdIdwnn/iX1+o48ascbC7P3FOoZduEPUr+lcOS+yAJp+eypAQY
kksq77ZXw53m0RupoSI1gl+JabOrMRg4HucHAq0z5DbUkdRww46H2T+6j7ZK
0nDo/Q8Kh3M70WKyDayEIsJFF+ejmR3qxXx27ZxhSxl7lIC0b/6vwF0ab21U
W55Cgn6F9FFRZIK7+tOgIBvcW/7yaJuEPo58eoOGEsJhphexCcKqNSZwF+zq
jyJKj20pAs+Oc1YUMu69UOz6iPYqudEtXWFVrydUhW/pH7tIj/jsZSReOZxJ
Unov9HmMSYJ8RmaG8tUo52H5Q7NqkYvw7XEMqhwzWHRUl6XcMf6e7blsw6mY
aW4SSgHOoYeJ1zS9KlZoubHAR8UVhmUMxxcHL6ak9ZttC1qBFM4P2GPeAxK/
p1h7sTYUPTGOka4XcVCKWRggoCMogGc60ePefWNSENzjMC+PgIl12oPC9pmy
sRshhQXtXsknc80Tl3i87+w6P3tx5tR/5uzh9rJOgT75QKdv/cdkGSqzfLGp
Vg42kkdXvqclA2blrv5JElSozugzEfFeisQ07oVYS5pCdVxIhOdngaZO+iU0
raxjDiCq90A30fWBpEkRg0XdJl0y82rfzBX2W2nGzQ2sDMcEZy1nlSQ1shKq
W5oxlm8nfaJeQdA/C0+M39y+3TmhX182ZEhL4L4rW64or7mYsHTkGSCB5Ytc
pH6QobPbVbVg+p8CPioCOcL8tmhhDxkvvDVsNa1MKg3ZfahDWpKkCQ0JAUnU
HgkJtJlxC6eA56FGLzu7WgmxGaBDJLAElORWJ2usXuZ0JHmikFbFbVW3ibVP
D4uGFUkmikLhUROGE786l7/gpUpnkctbWmvDbM7s7s1Mxbc1vG96qLUxDAOb
Z1KQiaAp4ksdJaPSrCAGl5sUmMYZhnh9OvARuDdrDB4Bwcpgpo9sIspuZ2cQ
A9nBQCzXNOJg2+NP2uCn8McqLgHsO7t9eYFOt+OkyH6OvJ0frNateUIzorfz
iC0V2uqnnJ0X7drUaKVXhUqDSO5quTKLPplB93Z9Es+YmI1JtAWe+ICgZjGd
/2assybWKmdZRIBnPK+ECUK/jwQEF8ZDaBIueMR5MeKluL3hm8K3e6XO6rw2
QlTg/zQffS6GFg+JI3vBel4VSsg2JUq4920TLN56TlPw8KNkSfOjVf9WMpuU
Y1ZfS/4n73M2fzl/l7KpzQfeUfFO+OWWwpurPjaaRTmj/Gf9IbUpZiPokpuM
Fxo4zOwVGGp2ew2oBVOrXXo+RQbtQbbFe7sKEtEFUrAc07EoynPWl9JP5EZW
JfL0h8l4D9L4gDlqzhm5nfvJt4Tcg8pANOVFOe1YzqmfJFOl4jJ2T/+tlVZE
OIP3ieAAHfamAE84FqKwRsBKhK9Ww/fnsB7qeFCE1SYDHVqNUS5SmFC/vc0M
sF/veSm7GsUstTfgMzS4G8xlrJA7/hcIqbuvRlw4O9qMWm5jEqKKLo09B3Ws
DtIK1REp04vQ1MpaXLBp1TEdPNMbBDgvCd5EuWSEYXjI1/GwlN0iZefSazgy
3gnY+oJBeZqWFWGwHR4gCvA2rf1ajhk4b6ygiUFbU9l6hBG/DeIx3uc5PMmF
7iKrl6oO6Wmq2BhkRKPwNmbIlEZF2orYtZ9e51zF5tg5ZMJ3p2vCcOC4CQqb
1Xo0O+m4nm/j5RgxObOn6rtCxMxIonjcvnunayg7Sgh0RuuqcrRQgLaogy5y
L+oRCBige5PjNMep5s3nnbslAEXIeVodMEGNL9VY2+7KsUYUE/dcB5qvzvv/
auMWVr8BpakHx7x/8TqZkZGL7wx+l1Nj5OF57g5fvWU4HIRDjnxrbTzRXbJZ
nvs2RTiyshQm8qoJILTLszqwFpEQb/Llds00lk4i4F5b8efLS5Zu491TQNzh
j2OqjsLPEfbE/vUZZjdN1yzkF8uMURXxNjUZriVP6YY12U3L80pmMbrdtsGl
Xn7/Ijm5AzFYAG2kKrmLCECQpNxUqBF1GlWCa19vdPRe5mmYnUVKOWBBB7a7
YPwAMgipk8neeOIAdnVBedW3cnISzB4rJ8x/x22KNG4gInrvBdUam2hHoQzq
l4S8sD6TIaqHqLGx3hJFhBRqLUMgea49VbxuaDJoJ+bmhNB8WA611oyq+Hmj
TbkIy0QGcIWDX6H1I7x+5BousRw6Y/nWuo8028AVRH93SD6wCA4gqMk/pyPn
quiZKUSudEdGy9RGTiNMCUGyl0/PAy74Spu55D3xCX+xQ+0opiazTqllHari
9nQ+Ui45SdhupKqdugIh/dEwlY6Xn09fKY/ebC2Qp9npYP/T6wMW2g8gypr7
LfztIWMk6/KgOCxW80lymQ0lI7qjJBmSYpDbs6+Zw8fhjJkvdUDluCVfdbo3
jEPoNZJH2x1F8UvVPc/isqT/EHvnGqYJAqXnoHawgb8Maa5CC+/5OeLHcTSG
4SP3/715SIvg6ubqRgh6YT1jy83uPRHHcYJB64ga0AAJhhoJH95rHQA+jAje
SJk3rFCBDhMenGWgTLy/ROm5XhM69AC6TUyuPi5Mn04M5t5oiRg+s3DTaB+U
uheqxRA7HrEoIgiyUlwLBe7ObdJf8KelkV4nPAjMwD2XxfP7knvXXZ4bYZuq
EhWXrVaCwzx1tPCSpddNwW3yQGYckrScLz+JKhVr5NDzw7SBXU7AXtGUJ0zv
7RAiwHD9M36tWL2I4YW13BZxjxKO36+zsACBA67j5aKLP2+SxFS4Du/xlrn3
om5h4ehElZ9PxcBLIA6GsN2r92HKFtdYvmId3WLXSQAW2qEmLx/NQClpVAc8
KrQ/Wdsu2ia2R/rcnN93yVeeLArZwt67AN7qlgrian6RuPATG3jo5hfh8Qnh
k7zIFqJF7c7qYYyyHPL1LmUYwH1y2stEIPFHKyq+/h0c2VvPZ2TqOYnVcsqV
Gm8xXhy6zmzyDK0gDnNwyAtDmT4+VW/FLF+FMQTjKfejvDuDd/JLfcLeTRMz
6c1waGOgaOr7UBxOSaeAvvxxbs8eIxtMWzqbNpGpLa0m+AVkDjDHoXX5sW6/
ZX0Kv9WhYNVgoyE1RMeodJ5eUngN7whNOiUc0jGv+ipeI5BP0c/0SZrldCuD
yApLdxrPDLqfUHICifu6/8qcEdIUkGilpn5yFV/DK7kY5cYxv+ErBequeTH6
gXjEkhAwLe+w1d4GnFWGwFyBxeBUIGb0UzRrCWtbqYkI6ablje7YnX0RP0LJ
gPSGYtDEXJpF3LBXDBWtXQsRpc2/koadoeU+QoochTwQMbWp97kGttn3MFku
EUjo4kP2kNHt4qcY8n0pMpQ/at0pt+BmhI/zWOwpCXlGAf32788D1PokrfP7
5/jIIg3cg0UJjTzWrvtox20MQyP9QO1h6sKnkJlYC7p3JfpWSodShAZdT1kb
QjLzjR5Khh/KXHDf/CEOOA3JzOfzChwuzKw4W7ZN8aX6jQ4jbMSJB1iZS5BH
qtBIKe1rWtvdy/vw6b5HlK90lZ9IKvMNQONNrmVsriVJPhTqhGlYLoV6rZQq
v+llvgzD0Cb88rm7wPgUAeO8WvwRgEAmInoSPLrzFcfzfgvA9Ta8CUKLcKzS
lKbhLb8c+6ybeE3j0qcVriXE6IHzAgmz4xvR6SZmFZlkTjy+UcdA8SbjRFmm
P/XZmDUqIEMy36ugAj4lj5eqidps+AFX5QuBbXyhE0ZWIHeXYIk6Ho4jDugm
ikJbkChUA19AywW6c65mu3kk766c8hXFx4DhdoI9rtCioLKiItl9XmNt9ZYv
CZn5c7Gn0DLIYbJS8/miROacqlOzN4XDuPhvRYAigzjiVALfyuWJprZ62ilR
Aq+rDO2ZJz7Q1xGw6XDYOq6K4rIhS0kFK0ajJQC7H1WVcWKurdVneAqJVX5L
ROVB6ZcTbWbCp+2g9NxcsR3qYVc57E/e8Y8QAG+ei7iNXQz9VXHP0cdaHRiU
DlMioiLEQ9yYJWubDhdn1bvI8fs18h5nfUFMSU4YHMQoNY2AD45K4i5UZKEB
eCP4PhoTGaspa/+s0TTicpJR0u7lyr36R3MvqhxVK+X5SzNJU1DD79MdizwW
piMcdudSS00onsZH/aTf2r/mbNoEQRUJhrTTrYcNgg7ZvsAD2aHcutyyLwG+
dplGGw8sxcZeKxbMRR1VS3KOEnPGMVpjtDet7z/3GdPBuOxFgslRzglaYBiQ
DnlWpP7XDknvoxRt960GaCcU2uThg32oTr0bybsoOtzYjIjFyGgeZEeRexrO
erG4Z5nb+cW4mYrBB91rgZnyC1fZe7iduaCPrcLraRBMfpaYm79qfIchvS/g
t+1JkKMitUoZ/C+Alyp77wrVNq5JX6WnOZWcmab11FPfFkuJP+M7XKJ0QLln
hNXhcHsFm8j+elhCXBlYzWmGDu99KhYRhSyAmHFOJ3vMHXXYG2ufeCeLMgYM
k+h/3owq10s+Lg8Z1f8Wq7abJveIvrlZOYfotlgLeKliuHV/ryKk6AR6NC5V
G+d6vrEIP4YLcFX8AXGqk508neOfBb5Odq1UZU0UqhMy6IUyzobDzdPY+2Le
snrVO+taCYUXzeMLbMOygO//thYFmiBur7KCs1qs+4m3906sevY5SDaTjuHM
kWk+2WMurHXxVc36cNAAg361uktGWQmZ5n8GLlPK3g4ayz5YTcZUAXdl52nR
2K5UEgtV5JLOXx9+9kPzIyoxyNZhIiU1EMhydox3J6ekmT31GSrLKn2rNDom
lqDjP3Q3I3PLDZuZ4H1tv0W2/CyqB9lyqerlGR0QOoJOQrFwhw2o3CU5ggdN
h7jO5a1D9tQQV6tPENKs5dZ0GK+G34A2q9bK0XDp9WtN5tFP3isxvt3ACKMl
VThDEY0HBhkwZ5VwdpFtRepCizvz6EDNUZuYWIAyheAFUrt+7ZQ/tiIdwB9w
6qQesjt8/jNoXj9XGW5uOGGhKZXDK1tHP2J171keRw1VXNa7gZRVuLq26Iyo
TeN83nJNIwok2b/qGrhDbDd3biv3jP8T3RKsNNaoJr5Fb4bEEA/NGt3YVrgr
fWAMLc/Sx/rDVOIiQUYeek7Qz/f6cyi3ACEfDdiH8R/ZQLBXq7IIlRQe2QDA
U0AiYxAbQ9KKEM7ANUcB/0f2XcPHgDVCfOUa870S8EZWtG5qobvvfxhIuF+S
WhrPekyrEnBnAlzBJtu+X5PeCArVvCAzEG+5IpRD0of8r0cM6opWpRd88rvX
NS191+iIHHxtOsk5DUkrFZW1tAeAWRuV5GtMJFyqdu9BS21ON9LlZa85aO97
G7FxW6FgerVyzCb0UExphr2+Y5OKAmd5cpY9r2Swj0cE8GOg/1PGuNHcXBoV
cajKIALpRNdjF3c/01VrOu1WvbVIqEJkefX42W+ILbq+j9R8h+loBDMxX1fR
d2Pxsct9ClM4zbM/p/Egdzob1kPcTzsjX45XCzqITJik+yJqc8nKyYFkzoxI
6+ENOwL7Ow+lZtdWH71yV5HxfA6Q5QckKQyOoT5VPhWM/c8762yjUqUPxIJq
PA+dEdc/uIfgz1VXcEqCuTFZmTqUSsRVnwJqLgre53v+PF6usHH+iVar5og2
7e9hJ9ERmJ7SjpD9Q1c+y0QsUSKeXYZv2armryt/xRp9izySJ/alo/1oo/Z8
7b4Dbphx8yQscEQLyZy5cZzmszihsgm5u/Od4EXuEsJsHjoWy6Yq1CctsbFF
ftWEi/nGhPuMIieguoGwOglHJRj3Musa8OyCttz8K1lU3KTUcNNj6JykDmdF
pCsd9tUHfBCGYx04Onpsg58kLGiv+FSdC2jf6Iyn9ydQUNV993xkYHLrPnfE
iRxX/KX9HpZijXQoZg9tWOUXQk3AO0YAxKRWVnQKchgXrjuZKyC2tdGObGVy
T07FF2hgi0PFK6E3kVU7SBDiHQQFmfhSamZ9O4+SVbiuwZDwrSEJT6jGVObf
Y7yrwVfrf0CiCOgu1GQvF9MyIeuKzA9IK5dPcT1K20KXW+fL8YM088wn+pFp
QdXB84czBP6IMctCfdqX77PV6/BkTt/G50pbBJYML0xL0ZIRU1CMQdk2Eaht
q3KupxD1S4oMRP4wPQSeYWaE82NDOntG8He2G5yWJG23zRUss781yE4GFdyj
+HWZuXUbWTGnqo0xNhgd7hmmFKH2FesoAeQ9SD27EHeeUjN44Oack1hLMkht
RoH9BydZwkP3ZFy7TYOdiUWGATalHU7MR1JizI3xJ2jj48AA3/NAtWPhSSGo
d4FUGwFsvKK9ieC4UywYOrkoivduOH2KzUpJU+f1KHFdzr0DJ+G4L0r++lv4
x04T+eqAVnWimRcvrrjVii/hNx8zlBVL76Tf6GQE5GJklWxdyXO8Rl51TuMt
GtETLtYvrKSW/bNtVPotYd69AXxy9r4bKMTD4qosy5HHlUmnWyq6xaPNn2dr
UYkzlBa85U60qKf7KMKP2tcNULAWqIVcJpIM+wHZXq8/ZSB6ntmM5o0HSFcg
XDZwP0W/XYhZZ+nQXKcQGm5sc9wt4tfRhZGPEyw4fIDL25iUW0fFAxxK3N3N
l2UcHtS3l3KF7P+n3fgURcyiwq2uUlAW0A5II8XTUlNpQiX5U3QpNFlyAWvf
PMam5qxYC2ksLuixKjvI76T9v4a0YewahbBnnInrPLJOsLDaKK90v7LQuCAj
QPGtngf5rM/RPeNWTeQl7t6GjjlDjEW5CESLPnrhPB01bEFpdJ0glnZiLS5U
KPO6BUPz6C8VN1PXVX73aOoEIx5eJShaUuYSs32Miw4X63+cxUdZsc656cRx
WLivXzB11Lc6gfBeB6vHI+DTj8kMTlbC/ePoPQPF+t2l7Ayh7TYAEcWbywtp
YWGpDBEIiAq29uFPEq72ju/imMzMbA9yDB+peiog89bmN8/yD6Uc/D6Y6dm8
aeP5eKU8SysFjo6eDeoZ84Tyo9nIzyJ0y2xI/SthYAbfuDvpJj/8gGeOKt73
LD+lBh6M03UA1rW4UorO4OClWtDrXmUMZuPUR/493s+RKgoGSVnLvItAzoWA
luw/Q4GRxh/x78etWa4lwuZbw8TxUNyKdfeE8yKTJeKh0g+azL8dWaW6kt02
v7WMDLJh9LwMOdtioiu0H4r8Tf1S+PssRjNBzP7wv9YrpSrg32tuzWnI3QrN
/tFtVXp5LfNJvlvnwblNIELj5PMBkT1duVZ655RozbeWeQRCYPdHTpjYeJIO
KQkHQlCcnakKSLmqIwEWNAWk73uFcYbr69xeMNM8fP6jZ5i9uHGLtlvWleEM
L9cTh0Ep6yFVzz0QakvVRI9rOjBf3XpaCc0wPkicVCwKoYBpaNgxQUiEBKGn
rqOdfNp11urCAYuTgDc5QKebPqhZALnEkU02QAeyL+4YBhXlRXYdjfxMBexe
6h0oFg8k3DzljMd2pSOiBnP2hdU9tJBScdjA29T+yO2TS8s0MqQmZ7BanAE7
0AA3dd0FU5fAY006OxKRV2dLfTP5iEob9iDB0hbxLWXcOo+qy3Hp8TVvZBEy
wWgDEa48D2AvrbMOcBXUpzT0C/EYU9Uos7ppBINEuPR+iho8HsaZ0Ddo9Tmw
orCfK/dCnbGlZgfvNtst3XipYX9h6VaLRz0pbqOlVxof7LlCuQJ2+4RomwI6
/c3gulsLpdF4D4cBAyhKAB2Qu6KpM1xwv67ErKQyuI/zsQzfYsgKUmrGN/lx
JwK1QohXGmkTo05o//K531QTyRAQ0B3bWSEu2yu6jTiN8Fo255k18q6oKM3h
61r/SwTl97Emq7I7XmOM9+p6trBL5ACmKJpgM/OM/2k/lbkWI4tdT2RyQ3E4
F43GyjkDVQn02lV960h1hdGT+JfKe3xX90MPejtVlU6cUuhntwavStpu9H4t
IehZlh6r+B4I9F5HSwsue3hpn8tyTrNfsYcHKg+wqnlkPFWCSDvVKep1hztr
/TG54CgKMlTiSsFTeTqHCuHIxesmheBe0hi1VgwEq7Qr3F7oSOt8wO30WYrb
W4D76u5m1Z8shIiGvRXKAbaTBYwYNiUI1VrO3XKDzJ4lPaTvK03GyfBZ2PyE
88xulIG32NyJ2rnccDr2PIITSbAmfkITSMXUh/kwRTRoVW/BX/RMTP/ULs4v
wLw2tv5HvvjNvgfXLCZ8t17b9KdP5dEIs7OJfVBPNKkZKBT2WbL8936okV0g
SPPxUu7a7OcPyVxTsY21hvAt3tvQch2VN97oewv3As1CkFMxolHQ7K6nspXT
CA7n/XIgIRZUMkGGA3eqIsS33jaCRSKpvnCapbtWE5rKfai278LJYeZ0d7Ii
SrGFX6ffxpoWqQutAVFadIxfCBD/gr/PTEIHiR2X2Bym5/OFp0QSMpLRHNwy
8ZO92QRxZjsggMj32NZVChn1WzqeIy1ao6kdx5qAdkPHDYFw2kEId4mueSeR
+PYBjZKfsukcoQeIYUzVlDl4lYeHIREfuw2ydyCE7mwD2AP7/77tLb3AGOO1
Fa0bJNWCBsrnny7dx3P4Z+ZijXjaYDn+Nv0N9W3iQeaLkajHJse0Zkx4Fs1o
Q27Z+yjdkSW5zDuSLxCl3faeCM0wUbeHNkDAb3RP/oQ1oKBNDi/Lt9YyQ3Jm
3ee+uAdiVk43hFog/Hf279jXHrRmLx60E0PpgT/m2oBXSh+N+tdzPkiZRHrB
6EF2awl6luYrk8WgeC/aabQg6/GumMKst74DWcv7uUTfj/N72uC5jrwh17eX
vs5mdp/pcMuGuCEF4zGlgOcNqo3pPFb+cpI+AaqaU5c4bBT8UJbt7hD6CDgN
fBysPOgdJJlYfRYfoSdS8Rz0maaVKpAmubt1XWZbNZ5MLyL8wygoiSwb2HM7
h4q4Og/2+BRWv+bcQbteoLAL5GmL2P4FqyUNVeDBWYfPBZoIE/p4gxkq/RnH
VceSIJzAzLFpLcgUEqSgen7kOiqRUS8XRi9OazLO/SnFolmep3BF0p+iZduH
ArlaRH5rRbKUj2NllmYND8iHibwyQ1T0tjHuSSVHTHurEnklhgdHmzXj8A0g
vruAaLZF3SiHNKlRboqzeJzPm53BbscDQ9RLBSfm9H0NCg86r8jSuN1VG4wd
hJiVOZTP8N3SJqD/6T52h9VLXO3/UuZZ61LmSdxwWZxHyw3ghq1XNTgiEMcK
FWweG7C/ftMa3sE9pEzRHqtup5iBzGBY6ARH9l9UEGeZl1loeTRhp1/X5hoU
AMQaclEf7MYPs97LfdsLapqgTA1hfV9sGbSF/AbmTN5Dq2Wxdd6HEJDf7ItQ
nKirLgcm5gvmy1YLryaCEz5+RkLUIukOYdLZv6G2FF9AF6546BqLDJgSdJfK
27zWlI5SK4JyMoymA0mz8BQtF5tSXAm/URSI5uaeFiI1cxauMbGi4woZSSRl
/fUHYnQV1Co51Z5NLnqlUtRl5Z3HjDTt3NyThqHqgWuIsDb4gFdTfR7oyx/X
+2TuSL4HMmKF14m7m74303UdjSN4PPtzZVntKu9Mx8819OD6epbEFcCB4TbU
oIwfT7RP+q8dXCBScRjDEoNSDmE7CZ5rsVNyAx31Kvb+4cGz2eBeEGhIWl1E
Wpod4NpDj+pzHx/1tMY4thLYyNT9Td2KbnPilS+zIRML1/XCI9YJPF1ktRgv
QqxLOxZskOfYKWUN5gpeKRR7U25NoZnQsoj3zgpdmoFK1KcdU4lib4dtTm5b
PW1S33TMkv34vG9Rites3KPPAVWKb3eGLcYlfeylKSz618WlhpOh0FQ1auSn
ItCN5mJw9Mt1TMaOvAjEIKtnYVSmJ2Dkl/z8UjJM62rQ4nyelCWA5ft8fTmW
U0XvEdNCs+6T9TxAtTOmDjhX0PBCAJ7MuNYe5hbWTtkSbnnfdc0II5Pc3GHC
j5a2uwSC9L9QF46IwF6aUazQviz+FcVXpURvMvtN01PQNSKCzSXPfy3WeZ2u
RbKbpkMXIYZpq2Kbn3VWVmWP9e6lIDB4n6ba5LQK7BuzmPNYvQ/LIZNsY2TT
XFV8mkzlDqRi4bs+/qr/Ozi18RuTMJXl16FnnLe/n+lttGqPW8BCY2LogXE7
00t5r8bWiT9C4WgE+suSBjSGxRYgzEyEeN5VGNCLPHA/8OxBCeaREzyNeYNS
9EbOkrcIqubZP5ExndQFcZn90nNWXPSdKW+vLDS6bsT8t2YxICPQ2E0XAV9r
2rXAPPBI8QIGv+9hMw9W5OIvonl2G3xDQ1r5ENFkONva5xobnq+94/NwqeHa
QsJkW+K4SGxYtXU5RQ9tAA+9JOh7fa1F9h2/ldhZQ232G8prI3+rBcWZfnsn
UvF8PdbqvpO/sFbUaqUCahGUFekuVdbUBJnrsJNFKcGPUmLnJpjZFNBZ+jRN
xWjwI1qII6pnlRKduCcuUxTdaalELG0vHfCbxWRpHV/IMFf10Rflqk6vcS1p
IkBeBcyBXqZ0inH26bR0F9N49uNU4T1E7cCykDupKUJNhiclBOVau6/G6U/B
8eY0VxGJNgDrmFrh/KsY8cqu6Dfiip3NvGAoPjP3t79ZfFOPrLqWuZA8x4it
Xcjw1RErBljieGuTw1VxeDwfV8+hUzi/UBD7onul2icJgLBFBbUEOGKfCCWL
nmPHTrPdQqelfLH6JkJLzIL4e46lFFt50f/2z9xZAsJLWuvG4FVqR7EjmoDL
3vUFoC0wn4QRyEQXv8cLCPuLyZ6E2xWIY35Ar7KMNGhfdxrieaDa+lVLX+bq
NDe2Q0CLTOKDYi0MxzWrhI2jYtDSctmrp8Qmz7APkbMi7VtE1ar0FH9ariJf
I8M5T+tRhW4/OXb+IwT2i5nJo7kQQ0XLLCkO3vAcjCwPS3zqVv3D2PkVkYxD
YreGMzjrFaeg1DfXZuAQC1EHHEALWc8KsceMjm0TUFWOnuWVK1oAQsnVDuIB
Tt2wMuXD/uGYCpPgTRrmxQwQAGzpGXwzGKAcSQ5CQoV/SQ4VDbk/stNgI1nW
Ce6bRVrpuaXps8qkmokDsNIQeAO/agoiaGhy/j5geTdpBrhGbm4rDrdDZb+K
dFeWIFICIao5wY84lamsoiaC7z0HOfS8Wvfyd1mx8hYYaDuu9Oh7zfC1MPhJ
yY1c0A5q50tWDt/4zSN22YJ0Cgl1zDNacts0fDHv8dc6FkgpD7Lv1PmpMazy
68KBL/T77fotp0ovIucJM4IIni3sWjWpicNddvnOyM5CmQfNDK8cie5mHoGk
n7FQQX1p0aTCky4G6RIHWGfrIS2JeDt1d4vmEUu7E7RhGDrJPTWmwppiKWWk
YZUFTjQGCkQm9MzD+J6j/zvOIOE8wtY/iPiKiEtjT2YH5Xv/0mWWdD9hmuhB
ZEOZJbh+nAFC0gwGtEYga5ZpgjjKkdMs1qyiYzO3qXlL2IKUvTV8YAvd3Wa5
PcNN1r4Hx1kn9yUtZeKHC+0YDQBYlXbDXpirvKiIyYo9Kj2sHXsgNVFPMISk
IDeZAuRcEd6n+wsj0puDISc5wYzjL8OUE5D+dGpWmxqmxxQJ45zvgKsfbvPB
3VBPIuYRUryO3JxaDJpN9w3Fc9HXNgPxmBb1idTu9HHItKVtmBjkg3Z7bwt5
+AIl25SwpZWvWyrLwl1zr+fqTX8mr1KLSKZ+KzPhf6/USOYkgHCU9BpFCdBP
lKh7xutOe/YZ7/OEv0h5xj3GudJTGiKzHr0Vfqdp0FS1OhFMyfjO0pq7qwiv
Usr0WRAoRH1ZFW4lSr5k7uSOjjd4e/bmU7ltlGVDesdNezl9CCYyCUsdLxDj
PHC8wWs96xd7pPYyGgbbLD3ZJ8tAy3Qa9Hyp/qoe/7EeEr7ZtKzh5iOLQd7B
A3sOD0mxtj7JijagIozLWqZCdRSkeAXff80HPl1lCg3p1z1EH9b+atvBvxGe
oONv60U4WDqOfEFfrjAQVSOsKiC4QNbYGnGc2vHokTqoGnO8dtHQlsAEA5Kj
j8lqM5BMjRCZWjB8XG7sGeNJoQaMd6ucJw1Zy6Deexo58H+S7ULqgLmr9TKL
cAacMedlyyYLuJK9aAXiYp0wrmCsKoYQRWp0hBuBNdpijHw8PSOyuk4eHtHw
oKj7LkNIRwmPUVA39M2oGFkz+yrjt2GrLB8PrMlA0yf7Rn9Eh55bPIi65YWZ
PmdohlkKkfCJiwDw6H2UHM6etfYXjx9ur/beef/2qPYrs0xa8EPhmngucJm7
QvtX1D03E72Pey0kG644SEa8/1UZu2PSq/175xaYKMxQBL5/FxW8BeSzwlo3
4BOXNPgswyZ6yEXXdbpzrY0U9cm7fXXZVAAbe4c+UDz/zcoHD5wCwsqrKArI
LGLivcfOQBwSR4d1tRutk63+ZZHdveLhG3hyMrPHa8nApug1LhAQ0TAYDHY3
8w0oNNeBjBbCSi7ggseAtATLwgY/hW9J6+DHJl6vn6zPJ/NZSHopa18MkMoZ
J7ZUSR786k5lA14XVdua6rawHJ5z2zIsEjntgAP0/ZKN/2VW8VkkJsOzKUTg
Ui82UUyzE12FRW4BHO2tGjE6qfbLQw3dGbIAdcAH3cR3H3DjpI97UB4I5hC/
NikWGtKhSVRbqjgN6gGZNylTdttlQDXtDkCHffAjr3WJH1Jp3Iu9EV+0NTrE
kYDUt69ZIMWIDZGPWTmORxOuQdFgVAWq8fjrqN9tgXeOCkbg0okiHQfU4/cI
b7QtPd7k4Te1BBAwBqcgoLHiX8qpvoaMcxrGPkzPtbFFblcbnA1ZYYNjoj5U
EnjQPz06x98xkB5pJ5RG4aqrP5808Wqbbd6NlbmXBhAo8007+xEN1NJHE0S0
T+fGsNvxHY5A5SRkCfoPFRV0jNoMiwERd3HySSXwqkXK5Vn/eFJSW6nbIH3I
hkof3lyBupm2q6VHOEb1hfTpiWUr07IzoZryS+8AgEcPDV7thv/S39uzbq4q
YxGQtkBFvoatMsOCOVPKf+nFQIEnd49WNz5HHQwv1Jva8L8UVgcOWxB4O0Mp
L+WHGeELluMC65LQF9Dn/vIO0WNT6xgkJBH2OmLlIaTKZpsjrw1op6fuuaVS
oVPGYZR2itokOVpkfqdH2e3XGr+wbkYoQU2uLhlpHb+0RqN+HPINkhrlDgLl
I1xrB2H9O6ITw12tSkfG7b7noIuZ9eca6qLNTzxjIqcRCZz03kkt6jSET4QJ
MT9eDw+aFwefkgnLbfKnjdxHurCXtPTzFNCm0JJDU8ovYyzJTt316BPPzgvR
/HlH8xApWi+v8cNgtVz3bcYJZV9eCKydhhQWDfAn6s9TbxnT0jM1DC6f5dM6
ZzUJ1wZErfI5qa19DRqhbdLAK/3LnNtpg4gYM1hT5/bjXNPNQJ+1KF9GySS7
o058wbqgN5ZTm78FHJCUNH0wol+5nIex/SagHVQDXkky/xbloXIAqGtIfHut
SS1TuHSa5l175ey6O7v9uPSfJiN964ytJCAMeIw8wjOZfZ5zQmM9cM8u315V
DSWfMJsDzeUTm6GLvdvPxCxklXpOkVD0lmmwXG7Sn6zjF4S8xDbR1Pik0AXo
qryk1XjdNnIdtujczAPGJOniIV15pgMlf4BJAuLL2wQpaqqCfz4A0GiQ/Sf4
u1Z4N2tmk64jnl3JRyTpKgHRKyTomlezENVBQTO3U1Kzy2kfyTmEwC0U+EpO
RPh/uhpI66A+t7z/6ChszsMb9L6olkc04bxtxxGBtOLjDNtiSfhZBa1xTsXA
OQw+37n8uPVWGkVgcOOO0pZfhjri9srzGWCcDv6kldUmeyuSwPwi+evxfl6z
Ad4/ug1HlYZIYrapOxbnI7/kEcCN5nQsqsITF0OxSS70iLUxsrm5bbFG5apU
C7Jj/NTAHXRB0dGUsUkmar28CXvOCXZcK58ZfXppV4XfTaSz4bvJ3KhMZOXK
RwLjg/mjXfLj6JM1WNPnBTbn52GheL9vdg67mwm6qomWsKk16nNmMfCIadxe
v394YZRMBY0nyjEwBn0VB7rSLxX+U30QSLgDaK4IYcrj53dfRScc7WbcjB/K
FsTTPju6cqTEH7m+RoSBD5m+ZTO31AtWeeWEmFB9zktI5AkPU6rlgo8x6pnb
rwj28sPnVRAymSpsHRBzzV6Zubo1RWyMxGgb+1/qE4Ly0VSPQJPSddn8xATr
MSQgWBOkN9qs1JGjv8yZP4EDuvmny4uS8chcYutbi7PnayQzbbD7J2pV2tJ4
WB3VWP+xCz2K8ml6cfOwdgwvSaUSJZr2+PT9v0xMAo6FOz7m7n2ZvcShZ5ul
6/hQsSWW8CAi67ytdp+Vfr8h/o0JgOQIU+XadAYPpjkKRqKj2hRjWhF4m+3k
I2B1xzrixB9ekaxRY4mLeyuQbRTk+59CRHjaQhut/cBSbv92eunoV5/ebr4o
WgEOzzIl0trGORou9c99S+5UU9hRUpu3bYQRGmHoB/b5RKsr8VZfOa+1LWaT
L06V9PdyRIwCHZbwvm+w9lZ1u3BRybF2XkZJRuVw+Pe5dkMDTQPFMQTmMPbI
xyYBPgdy2g0L+pXT2vyhDW++zYQA+X2Rimet/kTEfFGz/KA6A+aMmHFxTwHp
ZZK0G2daJjeotBp2YIm7OqUhwxRfqgDJN1WwtOAGMQKFpd9nwzHeXyIZGEXO
0LFd1WJkxEZdGjfXlNpqtrt9nu7GnXbjQLA3obn+QRdNU9WXTicwZfhmJszx
Wm8jUVfuUGheb4t1g/DY3fsGVu4lZFDmgJuafD9mTBIAbrH+U4dSF8exE52H
ohGOgs6tO7YyJmw0GbUBD+SQBS+4FYHnOCdSBvYJDwBk+NOZ8L9nn41ZZAGx
IR1fQ6urvLkoiZmj24clyNI9574w7zN4bBZu2uEBdLPttLegY0kcdkWggaCE
ePAGWdI0tvloolAwL8ZwBE4GcHdVbqCA1AohNmR1F97uAZYPl/g5dQC5pKJU
crjEJPuVCbwScc/QZD6EmczVpthJJyZVzKIwnjtyDIUm0t4Ah0oLAtfdKr9O
jr0InfMkG2UOgbYYhFF+6ScAaPtJ+C/h4lPqpnSmF/UbLVEpN0VSZ7XZtPiG
/s7zMQtNQFOm3nMnBntzX52Xx8FGr5q/wpETQrR2qjrhu9ZHYeQMs0NVJ7rq
3BQt/wVgddt8zOPeXEUFBA5iBNpWX/LkuGmxEth3GDLA4pBHkSOBqXOndGnF
X90EA40QBogGVzPfOJHjwAztGneoAz5SRb1SZqLcpsLMkAsNeZT5oIsAPiWR
AjFUO+6H8zaioetmg+w1/yAqGsJ2vljB4l2TF30KAa3hNMN5Kubds8bfsOVt
LNfNw9iPaQzaA/zQO0p46hZxYuQWTkbaReU5/Gu5r6895jBhUaO1oOENjuSW
MqU98Cc2ScmvgzzxyLmr0ULk2sfQa5PwldwvK4BEIq9GxUr6aM5ZhuCZGJvl
vm++k1JCX2WQqTY+Qe4xu4Q7cSbpTsupYumhqq9MzTzwFtBG9K5d5Oj9DkpV
YjTh4ao/LVi7beoCbucQb70P9JS/pLkUH3aZoQn7wkn+NbqyKaI5z7iUP/Ze
gMSfthvEAvRYGBNvcU2pWlcKm3dcyzqvDfAm0juZeCyJkEtEOr3MCnwu54+b
R7Psb4GfiItL6HPrTDYqX23wtH1MQvFIowLErwHxdpJ2f9jBEvBKk/T2immn
RDwT9wslvaD+aQhbvpEk+V3xiNSsueVi6T/2vN254cOrkpzZ81jlB3bRDAbI
kBrcXcANOIxwdwjNctKj64U/l31lU06kw/sfAxVctxwv6TRrghK0A9Q0Nudp
0NpYEMKJE0j9qZQbufaZOiuQW1yjWijHAKL3era2Vw0g6tQmeh0x/00bq12a
cjztlOKsufkTdDs2ulwp9AoiDMQ84QsnzxSD7TUmEWX2/1Vb5tlDKNj91zcn
668SY1vCaxezVrhbi6QZFG8c2qb+OV+yxLsL5HyutqRPIBvXX9pLCqZijDtt
3J3ZdiY73M30NITEQ1UhIXLuMRPnIB7S1WG1FgSCTSUxbVeHYAaOvXQfYxUG
WyGqsBUEEWwHZwT9hxUXdhpsgGKpzrlve21F2qRCB3rjzv125UnMkaCjW/a8
NMagVmKbUwLDos1eo80KtY9wkoc5SsV3JVesI+1btXhq2g4n/EXtlgu7ZHm+
CR4sNbV+z2Fx3f96su1IRPTTu9DvOXDRD7mW9djQgXtHuArYwADXb3Or81UL
+93NTLbBu0NPDFcImkm/5HpyeCtbS+ykvKx8ZIGOkb9ZVkMJTV53g9jVKNv3
SZ4Y7c3bsrXbd56ehAAZEqPAaYbsbDnEHA0r6ac7lMuCHADtxfbK1xvA8rMG
Iy21Rpnnvj5yINls8qE59mpQm0agHcAnRcvfCTU7JeP172DQZ3+flu5W29Tx
XSnHbyS/CA7ahbjLUruu2kmcJxuAfJlD8/liM9ho8ddreoyklKaslGnqUKMc
9VUrG/ZLiKcxccT0vgnvF6GXqIIgwjvRZ6AyrwMOxVmHv+OJSANvRsBV6En3
kf8wNzyalchtg36iMSNFgzGVZrZ8SYYat9jXBYamL4/DJzOmK0fT9MWoM2LO
WEMp+jDGhvHfhyoJ8q1DytR+93er4ibfnEQfEEmdWeikybQFVHeBW/N41yj9
Ke9U+Qu9NOi7+oqrYrK7P63REjKBi8KinwVKTqFGD/RhkMhdGgfVXZda2aKd
gG2q1md2fHm0rWm0VT9Am7O+7Q2zqyCG2X6rA7e0+OnxRRajR4n5ZKLmnZv8
rShxt2caF8zBoOhD5lQTD8Dfo0ppR8UFp9g9+nULUlrCdT6XAVitB3wfTXJS
s6GMsBK6GT37cgWoX5RaMP87ftL3mrG3foA9//aJ6wUznJUu82OcIIUaQx3w
2VLxgyuI9nBJhKb6Ji/QpPi7SiQH7uHFCH9YKWbP7x4Ov++irkg9jQgrjTev
gxDEkcdejTozulQHUjBGHH24kBjdod9sYikwawKPa8Wu2EJPd8bUzxBVXLR0
Q6uULT8oFgGSdI4gOCFdaWQoSW1gdgcTmgEw2FDrmYre0aYgjzq9iYwEZ8H5
Fhuj/nfNUAEoG78W0DzFMh9XZ5VYPBCWWAPYODa2pjrT366L6rlViW5zIjJX
6vkRCnbXVEvPRAtDVKa5/HenIL3i9cR4KCg3l6TXL3uF5WOIfUvHHtv/BGZk
a0PT9dFoR7/Z2a0hOKiqoVVbMQS0I5v8ppw+Wk3x3h/sOFgmT8HNzBHboHO1
s98NzHyadeMli002hAU7Om+XvLGzNZVJ6BOQrp8MPhwwRplJNmgT7FUa8cvp
+FNlwND3/4RVBO0RYcppcHx1Gv6HfKq/xchak5tlUs6GXtGz186ujSGD3V2I
Rhj9tFc+FApT+8c5rANk8Ci6TZ5xpE3sbzc1oOP439PaZn77T0MLKaSvZ8qX
8Wyq7neqsf8EVlUv7Dxzy3hloo6iGufckssaXIQiCHBSBHMxlSBLU3RWqy+m
E+ZAKK2iQbRFENbFL0F1n/ZM4yve4LNIKvHhgJ8AWKLxk2CUweGkkLRhaJUg
ciqK+8aWuRoq6eRilj9zJBV2s5FFMUo/yrfEV199jiE8rgXVcJQWBD22sHVH
ExoqtY5w3KZ5P5CMMpCwpRIRQKo3q/4rZq6W6yVgUyyWk78WneepHm0tr7Yi
ujgzaS92y5SZMa2xVRxfRkQoeO7OEEDfZ8BOmAjd+J4gDu7E12kya3XuW8WT
T+ddLdbANiwV8GZxW62kZh3FkQdSybIVhpg7mrGl7xaILbsWQWILGSA6B1aJ
26f2SECd5WoXV+g9ptTlp/n2dpiKZ2ctAbp5d3v34Z87Sp2dPfx1/xXzlziO
/hGZYN3soNtugDUIB59YyLAsm4UQIw3ij//ec4Hpsevz/rFJWDMOCrEThdRV
JNEd5QwqfDpf+23KOKj/XWUXnv+KzXwGqFLygs51eHa0a4Pw+W3XKmhZ8Wvx
IjWEdZGtE+WuV3JlLa9ekzlJxD411OjEVEdZ/4enQ/9lXYx7/kWSdxBhPJhS
wrZEYvm1jG3Dz2RPu19WeZsjkiAOhbGZUVvyG45z0JT3nJnZTCBXWsGry9v5
7UjWdl2aJZvyX94jd50/zrZTTD9XNSQSAPWvYKGv1m+UQOvrVoiEaisWnLsZ
pT8OpIBV4hrt5t5b1Xudd9j8eEbjS9zicf8JJQr+M9dsy/+dnyd5WsBrEHOV
ryc1Fvl00dh1ZN9WZezzvPTSADgzyKoA+cSXnGWA5aPUB2dn2FyUgkJzJ6vx
hsf9b0KPVp74hKLi00Hr67dfBt8RVkfEhIL6vk2gAK2Mv7yF0Im22wrvlBkH
7pBXjj81a2Nz/OwCYM84CaP9rgt6yE61dES6Ek299fcd/ivH2XfWlzttENI7
yoTXmybR0XhtNxRoj6N2dtBJOHLx3e7+mPhWHaciodZONSs2Ow/1y/lTn9pB
gINja/F8EKWFJd2WXuugoP2miBs2l7o/Pk8l9YmduSuBQy9haz9ES94SwdU0
mCviXi9ZPajsZrjRU5Dg2DtktqOCZgbaCVb46lx0RpqLZTKKlGSm7/AtjwPV
qJEjqg2tzPad3OOU7PW669SmaRkD32M6GCi/vcn+e+9jaBkf1FN/0IXsDFPf
xQ+Wqnh/jyhiq2ZfJvj9r8Fwg3GCrkVB2bmzXqbYJUsJznAHIYXnBScIuGOR
Pgo6X7MW/t0o5zHLyESaec9e+JX0d4v4WG20k9PJFSCFmXYmJOHP4/oeT06v
BtVuGCbY+K+cR1ZaeLbGuY2JtIRfX/ZlN6aT+986Vjeiqrr8bRqaK8F3XLoH
A7XV3MCIVTrC/818hg8OIkL5I+flx4kmR0DaYdVs2j+mF2J5nZuJmO2b+wP1
k7krVcSj0q3UfxFfst0g0YnrFSCdPVRl9JjQ1bENCvJc6PC4WJhGrXgRbj4X
vTo2+fpXXrGEwEYFepQhaqzxGsT+rMfhct8K2sgJ2QxXd4Of0yKC/oczKiK3
19uqpQfGJZ677+Gj+g+5EsjlGxSObzswq+lZK0SdhAztEu6ixWpqkt06D2yB
o7H5csrs6ypi7LBdZhCZ3g1ARMXpkwiSXOeHGU9HLiimlKVYgPiH2ZrSRDZH
hb/u3mOMxmv2ZVICMDjco8SSbBso8w/O2oLgwPXqBO5uwUWhTQDm81ZJiHnq
uMQNXnPrUk/NDtrEBoEfzuxYJTI7aGO1+j17tuPDyvWqWekwY7/21jht4AWA
w3fh4ojYBKpb8SisBM958+iAzWuZ7lOP0xwqOQJbHDZDoIDsWFJ1TnV4eTE7
2FKJTgTlMYlx8iUm3ClZ6issUtm9/C58R8BzI2giDXVJ7Ix7GVcFqFRN2N1e
V0vdhWk64ck/EG9bRI4+jzz+0fwkkunjkYUpn6NlK46H1uZZ/S2y1p3IRh3k
re4svUTjD/aEVS7grzuZ2L2j8xcuZ+Kdkf5hA2/yZ2EPWE/nF7sk8M8Jm+tJ
32DKjVRN3WpTZtLhz6xWnJBJ6V98i+08nUKoUtcXqLM2TNEwulLUR5OTyKfv
0p+4fKOLkgLjwb/w19ET8cLgEzL+a7SvseoBgBfqixKNzh8SPH0+bj4ef36c
p7gjWzMEJiZPY6U2du6/dvQMY+Hs7QNZ17qWWbA1gVhYdlyt4A6nKnBWQ9uj
OhzlSSEyI8yjS1yEOjfJeyxeX6AeaadUddLGelM9v0zmc1zjTICPc4nzKrF0
AuE0xe4ZN2f7TVahIdkffNPcpEnr/SUIu03+m4aYT57UnrL+jwGWoq9VGbJo
C9trP30uymPDOIEn4NF/0iQRjDWTAvsmUvf4MoVJMY9BE8ZWZD/C0yy0u723
YG9m3lncXVelpoUbeYlwToToSQo7YkyLUO4VF5tazDU6p+J/MNn9bunHi2PU
64i/cLH/uWAvU9PXjPYuS5AdB17V4IyRTunwXZOx8L0ZunxjA8JSuANhP8R3
m9RYD5QxQVn/oDlCfN0e9EHVzdhIG0mZjvi2IqunfrkofbB4CwTKYJ4byS5p
6BO9zl0gJSP9LHuE2inMJ+7Jg2ODhS227URJIyj+H4c24WLtusz4QGp0YuPT
oulpXTpZgPlGz4Gxx6IvSqMhTfBHeqXM3B1qOdC9zqE/bmhNnZPYphd8f71L
+6bUeBNZkVQBpi4CML2g7PVxVbkTXo4epDtsD1j+DAXSCv/q0BwZOCVH4CHr
zHoGyQ5EFOf0l6hsxA1t3VY5xYEtANnXqZch+p5xWDD5dKdzUTJ5NUSsw0fb
SYL7P+F1ctUvkJviwzPjtP6RvfRJGq9znqP0t81gmxTwf4swSTi55pBh2YlL
2X7Vp4joX3MuRAq3jNUlgY9wkXwyQiHOUf03p7sb3KiGIbuB2XwZZ6YeMRRU
SpZqd2C3C+JJCOUwlefefV60B9CrsONnJdsdu+y3IQXqgb0oVOmPCcBYypOo
mC8gCPGmLpJt8mq2HamhiWtZTqO6OmRRXW0ZuMxvr3bHjvSfHsBegJWMQkNa
F9JBZ5Uf3XSHmNBndQt3GJ0OVOuH5Q/tH5ki1tz1sVBpwCeExoErliYcyeYh
UEZaHFU7imocFxJwSjZW9Jtu/ap99saH7HqjAkvI0/RjjxgPthVF0S8tOrvw
S/Um2KqApt3HoXqLub3xo7eznRmDf16ry25jiI4Lk07ueeaZRi0ktvb6syfT
MQoaSMhVYAd9pB74mQFu26HnbUE7KqQ2A/xmoYL2LFjn+9aCLixPMlXatg2I
qHpeY3F2y9YafrXWmnVffGJIdps4SYOOPUmTv2+hx6nY6/iUz3pGlEATpQo9
4dtJug2DhXVN0jhcpgttSUbebIbjTHbq2iy/902YqIacD0w3cVQ1FcJrwM/U
o/5FwwIiQ9KxkBjKXLUioa20hiLesFSC64pXebHtgkFtxP5ucy7OXpnZm0QE
7bsdY11cRualLC4t9CA5SEcvnWBV4s8dkqlupNmTAyGtr181OV/x9ovRWkrl
sJAnA4SbAWbPmYuCHzUlOQkbZvbxo8vB/0amijT5v7YTtY7tTTP3dktOu9gV
KdQUn1YmVVjv3UvFvZSxeVHePirLXtYb4/agW34EkYHBqNCf2JT2I7MXxpZd
blwQioXjSfQHqJpFQ564BgOfrxXzFzGHuhWc1ZfUUAgG+C74GiKW/owaxluI
ZTo+VgpnrV/EsrloP5/HlJ3WYYENANwOu7iwLrz1sELt+n7tv016VuQ2NJTQ
SdgvsQ7FETiObZj6i3lyQMBae8pXcA+AWQhSusTjT/eOLJyXSbgiMZfdO2o8
IVfHRsaKxDg8NELKLfuKLMZDMygVuVC93C6T7vjI65hhFwJemTNn+gJ7FpnS
xXpUECFkiwKp03MN5HOJvgPnXKIHSGEv5LOucYK3eC5W8Z5URU7dLY+tSj1T
8oG5Y3fNzZSNrtQ2wADx15LrwHAp8Jr4z9nLsVdzWGTnwr0LekpGKDd4BnWj
0ELnkxIs+Yg5yBVkV7rBWTKfW7Nbm8WGYDUm+94oik8nPefqFnsHaTA0UHb7
wXEG3zuIVAyeMCMKq2JvU4g8wE1gN71XIencHqD/vICyFkw/xB3lb7ppw6Rr
G379upwhiwQM2/2mNEuyG7XNAOJ5KWVNpoGDIP0Ev0G9JYLkWEig3t2HE+nc
YbFaaMEpwOp4lqgBmMtBTQ3QhdkW3y9MG9qy9iNAOABakjyeoGZ6zVdFFD9k
MvgTjyhH1ZWoVYArDfxhP7ft5AbJuU9aIQfMzp+mI7GuAqFIwYDOaLurkrkM
rIR4EqO9/0Z4yIVVC8PBJUJlAGJ3xzNXb+vlGd/BQkzEY6CDHaJgiw6c7tmA
MLT0L0bUa38JqXs3L5IlvZXHNLp/85bdbXMO1DlClHu2iIG4TDiZmQW+iSiW
7wE52o/YNIJ8oHRLBDtE/tfFXYc+UFGcGdQMrsOHTvyxqzJVgtx7xHxl1fWR
WuH5Rq6sQ7V4AfLBi3dPUgZ2KAwppKYc5iq6CKVe2ydJoatr2PUGDZcQ0OQj
w52DuY0P55ZQfHHhkIZv42mCzZHMmvbdw1dvUNFdR0R6i6dFw0EJ2qaRC6nF
BkeBswFmwchzC/W0Fdf6ebq4Cv3DVo0iD8lIfLEQux+qeRBPLmsYAeb9MTIA
FmpC/ZhfkB7RmG8bWEcfxTs0UTKWPRWw6lves0YtHfqVFIWN/xYBYTUuT37l
pYJQGrM3hvX51c4zs7deViFzVlmvYmtMdBbvrZv5fXkpwxExQNARgLcOqB1J
BqRONtDWXf48wXREuAEXMiN0JcWTjrqfqv71O3rCLazb7T2c0UAfFiYvDs2p
TEUoj3v8GZAJw/M5WaKsUKi1xa1cz6AZk9DT49QHoLB4aRVnTdPhyyCgC0dB
mYfNdUrxSdKaSocu/97NXZ9chbp6Q2vUy/llnEadEIJy8gVLSTtJMDEyzz9a
3A7bHgtbNt8v7g1wAYBbTDdDpCLXOW+byVeQdBdUeuuRbaS25yGB/Om1CmgW
qaHAx5zpxseiHno0B7ZmwEMc13ch7KfYkGEBnKy0CosOZJsZILvw9gyIiHDc
dJH8FZNFS8gmqjWDghD59r45tQapPMxQ8iVTL+RJ0NDF9x4xG7etuicyC3yw
xXLlAbzNYyg9Gzr2UBQzYFLVRfDFbXWlBrPYw6U0iUxqn+hj+EXUJQhZugrF
Gy6qqFWCL4r04KTHgnS47DrwyEwFUWf6Od+BmQ0wO8wImzEpRYzFoAdBaeno
TIviCOwFwmkv2LCcHAFS80cc4sJCUeXYr/HeXT1B0jV2Os3+y8Dmc8JAOL7g
YNtoGe6pjptTAggBFVus9tBv4Z7fTxneQ3vQU9Xog0gsOka6ZmxYxr423fbv
QKb7dH8vwCQl5ltlKtIDB2ewFaSJqagxFNEVrPeqqWDMBBg0qDkOJYK3QjqA
7eHPLSnjiGwNlGjGCWtskDs71YKWEicknn2rINGfHhXQGAscrXCHpUC5PVRX
siH044+yYjc395L3vTmfzMmcFYz88Rzgzjv0x0SqGYD1o6SrMZUhneZRkONK
CpESblzeMGg7ed1aXRITYRSw+pvschfn7djue73OpcZ9mT241dHp804inad5
GA8mNThYlIW/FkqqDQu1dVil0DUIHPtPgr0jfdFjgKTbC9/RjwTF3eJDnvQN
F163Ez/U22h51bIb/YV39bIBtxqL/7SPAZ+GI3w2IRO/kjY6AcszVBctP6z8
TSQ9gGga6SWSALkw/My4uec/fyCe3O1QknA0yzzsyRwT39oxj3nk6wqPXwe+
UfXbc4xphMScfODG9dN9+SJGgq0iDkFo7ZyLIHa6DPRuAeb+fvxYl8YCYUCW
9TgVtsxTm6PlFYZir1iblgET0DmIl89QSvNLG6hR0hbJdr1nskimoo9vgMTx
FG4L4hdQCdM+gED08DK3haWFhoVNLQ7vEJAsFbVgYnId1yLA7wn55j2BHzjx
6fjt579TUNpSEnBzDOaraCZI6kTIxGBIPc14epQBkRDsnLRzjHEFLsx29Pm4
cYS6yYsQeKYOOzgAqqR6S8PsVXiyuspZOOgFPYKphcdK5y4m0adg/S0V51s9
my33BslqO3lrwrK0S47bJZ984zc3x29EiZDBXjBgVJ9Xto0xYFBjvXjhzTVQ
vRVyZDKu94pLoQnh8qRj0ki8sLN6l1PCbeJYJutXitIDnhunjNwXRyhBBjLW
DMPmHY2EwsTOPIc1G7mFAFclzGYFpxM1R391QrOpY21R93btH7tGqTMGsHVR
BUgk1C731qc0+k7Baxru7wb129eq6Rb7+boFnP/CGj/hKP7K1afTtNvH2I6t
ROs9SNMX4kRxyGHQdozWtxSbvrIQNyiWSxBa7hibJYFW9JIU2HaNjjuXBoXu
9d41KJGbDQznCbAc0i31JxaLz1kWTi0GXMcD8R50ZjyFvG49uAzmyG+yVE/O
Bnb5YPVleDxcDKgDcaUKNlH87WegJcR1g/NYq42eQFwpsMn66yLIsiWCa5oT
5dzlkyKEN+fA/Cnz9CFAMgQkO9Q5nP4PnPmcb2buE6NjuIHkQSGG/RgLp1sE
XMy0xUP0bcj1Mftd3fWwtzWv6ND4vHh0t59p83/Wy9gCiZEh+/rPPzzAeHxa
KRIshJMA9NhP9OyvsAxPqhYxii0HG5dJrPtZqYcnWlJIt/4amLUOcGE4ML7w
MaE0TWEaRxKFtObtKzU259BY8ryIiYYfSASew/N2CpX9Jt9gDk3jbwWgluuQ
3M9B5tYCKyRhDUrUGjJqC2hc6WUFurUaaIy7kax+ExG6P3aTouBgPgG0EmRC
D19hkxNwHFaYp6MuaF06A7zAgwugSo2NSMpLCWSHWskyH7j4Ak4MmphUNk9r
ofjmthRyFLquu8RCD40CR6fSXxElhYYZDat7srtAFXZQUSKkCMpw2n4Ys1Ho
rnk6HKf3j+nN1Q0EQc7UD1IUHrPg1GG2uHo8LjpaFAA1UC2shcgDM6YcTcuh
KuWwMX/WucNklljmbXCZbb3GUu8vI7KgIM5XFdpS6FJgN8tOqT16rk+nc2uu
4XivNYnD1+7RRg0uFQJ5Cy9q3d0XYYwcgmUH4ULq9j5F3Tmdav5SlyFWCzlB
2oun30TdHzXnrb2VvBGTsc+aGEDq8Ci+iRq02yk2+UqWnvYKeBW9/VlCctrT
JNl080trfQVjZEyCah8DwseMdFJuLemal8YrekMmwKPc3U/wV3DYBveXWUkM
jeRSsPelcNP6xlzmoT1ZBGTjJ+NJqyd3YKw1x+FsWkjwY3uoE9KdUjXn77zK
Yk87H9n71xui9Gohu3d7lk+CZX1v7Xto0XV+fNIO5RlbGfQbnCJkX5ZmoMrK
38pgPgtrl/SHwLxtkxV/hT47ZYOCI5TAqFUdFdPVeTDhY8LADwcUdPPaUGU7
I04H0diYGCRf6C57wqGPQsFCCm1P2bsrAABuJjrZzv80ASoUCH2zy/zN8UL/
27n8XsVWanbcbyR7ALAANa5jhaxQ57h5uNlaKU5s+se0jL59KWxNtrbvm+1E
W/d+qbybIIpW5y8/lvr5vQxU3swAcP53404+9N/dETFdRUiUR43Mq66MXwfF
VEfwzVlqnv4lso+1DfonK9HMC9o2Amgx978ouGY9u32lf+jzAmm0WZObdw3V
hrULgYOWb9NxnofBbf1wkbH/Tgea7L179i5Qvni7Igj0fK2CUd+VxyMJGwv5
RZvP16aVAUrc5xDxC3rQlH4rb1ZUDuIO7V0hcRgcU1VEOGoRFqcnGENc5cHn
mceLCh4t4UJMl4eWZkrI8QLVtj0F/cvzADAtthE3UvkhM33VRnK+dK4cBYvv
h+nRhQTzvXOvw9P1EdxdZLPBwAbY0mngk+EpFwm+4EdNhhzg3PK/+X/Dtly9
yQyQvc2dn071OXqZEVV3DPowVROpu9ifg1RgSbgGeXwfwS4Pv9cfcR7J4S0T
M+1TQ6+1qV5eWtbwtNrAjgf9hDorvlsiTjX6wuk2+HWBNqUYr3232N3m7HK2
mGlPS0H0yy8H0Qs+o/EAX5W3qYrUe9y8aHxT2aeGBi/3jPcTxX+gJgMmC2Mz
o1yBc73FSn18LQmlz6S0VeKW/vmK4gF6K7qWi1FZUarPyoBJEiGHQkuH45RW
RxKPsxKy51+Ljom+dZBhZl5aW8VpFm6DcUsUgGjZ3wSDKyPD8xevE89SWugC
PlnNTOSrI8peHhhmAqBjpyUuaWuxLOpwlzu0XDzqsB8ZUtb0fieERUuG2HEI
rcFbIqJg3vtX7b0qu1vkK5Sptw34zSe0Jo8m9JgnXSZr3D5sDVK0avdY4gRo
yQGokF2nXDLBw1a3v3LmvICeSHBLQfoTNlvsex9n9LASsEQgOeRhr/7gTT7r
OImD0FwgXJjoTSBNHPZ/5Zj4pTaClN1wqmmHbfV6/usjpCweLEGx8vdlp/jg
CKq6YnMQMefzrpJJSpNTlvMaO1YD8/nffCtKhNRlXG1BsQT54hCnPgpbk5eQ
Gbl/C8v5II8kzmcm2R9PIa67FvZEfiMXPW2hcGgNckFh9BE7kuzXFT432Qcq
ZMF/tWDVgceIgOMwhMy9SSnU9QjYz1s5nLmCXOnLiwg9IEILr2cPgEA4acRs
wOE18Q99M+y7YSDDF8gdCm6i2Lr7a9RfffofQVl/CfkM5JxV3+yUice1X19+
RDJk7pZ9NUeWjSbA0BGr6tcz8FAztLJFifwJdOD4ZUSPZKhCKC5tZyKR4chJ
7o44BzDfBvaDJjIpUk16cqhTGFgm1uxc3D1bpNbjLwyeWaIS4YzXNkMEoDXs
8gF16bAT7iHnh8hHRSAow111BPYjekzaf1UG2GME6+liXwMUD+v25aIVk3Er
dJ0YgvtL79T20VbOMxoo+xCczeC9fRNCrV0JFN/izTGokwFkfF6rzGeZPf0z
YI46FCZ5SrLS5ZKBDU3i154O5Q1EGxJTUIiQzOb6MFRHz4xB/uLjQnyGP0h7
ui6KtSeScaHCyeIA6nz01RM/EsHo42WCIKDFhXkbStoMiM9sliLjUiswrUW5
egNIgqh6Jga4cfDJFpeBUr1lc8TSJrt+5Hcpe2VnQ/sl+JsrEAzimXkDUJWp
UQJUi/RL5r8w0VfMfprZTGNZ7jqmw+8Q3FmR1Y+iekUhyKKQq8k5mgVyQJKZ
wq6M+OlTTTByagN9gQwbB3DxBQ4nN113BIqlPAWuf7TR4Z7xyeNTatFX/u/G
K69i+xcN/i2tQ5gXNpTa8G+Xgx43wITguX6GTpWhPKleBw4hWXzRWDrygpA9
VzD5thTC7ow8etsWBOoAxlDL8vvT124pMLLnDYULwWwkaOkZXynF0QcVY/m0
nh9e2THnvqJjoU/UOJf+zyGhsQpCzWY5bT+1HTDpgD1c3e1P/LwALgO+QwYP
UEoG2RE2io0RfkACYzGslASSNiReC13QuI0kOdQQYvo4Y0tHq8Tli9qzrFSm
s6bhIWCAsg1W+U576vKfdI8NQlaHrbtKJlJGvxtwonlLPuL5mpO1ZV2+Q+zf
VxhhNuTkLv/lRT3j+daWPyfxxQlXiSmHGsDk+CVwip5VCsvtFexsb3JBdjov
tc09JRQF0kHAtzV4ImXwqMuzO2M1i8l2bXsQhEzXn65PNXMGq/Es4Ah5+Esp
8ZCv8HPcl8+z+eDH3bMi/0X7Cra9S2g9r4+Oz6EvonNl8GnqlJyoZDHowcq2
I0Y1gAFpL9yvgZdwnntSVNKqe7f/uiQiC50Q8b9SZ0DdlqGEikW9QJUQjMrV
FxFtOSaQa+l2S1cnd3PqqFyCAr3KDZeBQyr0FSCa9KT0yg/WACMCxZhm0nPF
U3DsVZtVuhiwuDxCMCbeCtb0ozu9/0c4bfSl97FnUyc+EZV507XpaCqLf6Ds
oS63TZr22eClNn5JxQWVztLDP0/wE1fpkBuWf8dewd60p8wK2xVJZdDtxlwO
lbAAM+qYAO2jH5kHaXobVpX6BOoUIau5CzyIuPSNBLWBNFoB9pVkjhul6TXb
tU46uM3NfIKuwDmtbvj5dqKgIZlBpcYVj4OzKwWvhgPUYbmbNoCSsJE60J5F
z2q4BOSxExtv0EFFlMeW2X8yR0921tX6WvO+ypk+/4VBV40Q+vmUvTVCW72l
ul0LTYP5brhqdODxSRPXeFFyapcSZJb1Ra/5PDGZhxmOeP2tbPTKghC6SwKj
ckC1BcWAe0ib0lB7lcxAW6FcwKhIrBOw6+wxKtxr1bQ1C1d2Nhnfy1sA3Mw4
mZQ0AvldVCmgtrCqEGb9lZNHod2ejE8dwaZV9W1199FWczXirO8Pa7VSaWng
DTYHjKxXm/NhJQlzX9lEvBQz+Gf8uIORIAVMwL9H6SiFPcsoLMAUh5yethxv
CSEOP6RgJ8dnhs77UZDCNgnp2sQLRlv/zlnIlGbU36+tKATGUZogONYjp/O8
pr0fwG1r7kcvWE2D2YYRCLB9p3fAyP6QVp7bp9ohe5mr29j6WSUDMkAu/6Eq
5XVEr7Onk0WZ1fvVgj582NTPGBmHDutsYDFpxBLmP570FKCRlaZZpCDKfEDI
ipkKHi14vF/q7Xp1VFFOAHgIDajHr9DjlZ1MLKTr82FPY3nvmm25IBMHgFmp
0h5PcMF0A1jfX4+eWsQX8rToHJVXmAlu7pq7lV3DTwkJAo52QxBo+Wrodupv
e/fBeNlneVf9F4QNNBeF0+OWJgCdA1mkKJ1E9303MJinGx15FTvw9Xc6/b/Y
rBuyxZEx9EItIISZcGsZ6ODuJQLRo6vkCgM7S76MJVJB9Eq6PxsLC0TYSlUT
bA5Hv9nFZHDnAK7OaV7H3xUpY8PGq27aFP0aEDaxNk1Aq3uL+6pYLDSwwsER
5APgJoe4qDog/R+Lb8m93B7xCZ9jX5sG0hM+X3+kbAC3cPXsH5i1ixEoa6Od
cR9yIDX40FqVKvY9M4NoyJYXGskFSLaA+3JRFiKAokgXZJWHpU6qulB1g/8w
Hart+Q3NbkXXC+avs56tTf7F6Gn439U3zyK6cfFPQ8LSuV17hOkA7aIyO9cG
2gaz0DeROshkg4MSbZqweHL2ispjNfa8z6BraQb6Y0ONtlv6Qa3asDcttpb/
0MJ7x5TAqZOiFkBRsCEV65SRbVVMkyLB88OpZcZcxWOdc34XtrUG9Kf9Re5/
ejHuwbRZjqMIvLrIxlmyvqlBrTqtzQMXGK7gotcIjcdb0hYVS/PRD1dlrYJ2
Nd2hjs8oXIa0pQ0F56oFmIm2AGqqFcnbLreqgi0hffoUNIVBbW/nOnj7XRwy
YjRS3Gl2UzxeBYD85dTH8tSLIr+2J0rKGl48R6MoOKEEg2z7Di0whfiOs6xP
lOjUkfKesjmpajxvyCUJkBBkpLZuISIvX1tfkbop+TFdI7N+f4QdFeDms3+w
4uEHIp5R6YAOoRrCUtehSKvpVFFgUQRnqLeVaNSuj7lEk+6gZQUJ84KbrTOr
eDm6TBQz8iTeawnPTiKkjz8X2Ec9BRRzxjuz69Y38fkCmXFA685LMwjgeyXX
kuXKnstXh9K4LrvlzaiyI2EsO2StXiBhW1wavbvjHGToeCRcyIdA6pedIh/6
xlDb/cZVpRZ3in7td7ISm6m/JiCG9q2/aad173tGIxfOfxWevdfvq4cMxFQ+
cDDjde4fVAKsLOs7nHPrUaTp6yvhiRys6napHU1z8FZSKQinWXrrDLD7LbPQ
fiOQC2vqMjrKO3o5kyL5j0avbYv6hpQjhAIyAbl3cNV8o4vn5WcB8ewsCuSp
/rJ2LkftC8xJexzu9ARzP0YbLbBgbjhZ01UcI0r7rpu8oEudeLCHoV+kXxbq
3V/5mYcOcMImd6TGdYHztbVsGG4nox3wc2OFgWfr/IblZQB62YuN/Tj0e42G
R1UznoNLOFvciVkh/vWElvj/d18lN5fonoRsdvbSCoA0Cx35Tu5kkfUcJg+R
MDMoPEA9oDNS+qy4z0FrBqT5xO1E9ArpviHs6svKDWN5gZixWPoFACMlr0Le
hT1unfAyvu3U14R4OJjDAJsXHvy7uJZ9a1kjIWK71qzXT1qcUT5e4EH1njhv
PDphIOI92Kt4fmSUf3SMM9hMS4cD4ncLYiLV7jnBL1vGxJW+RcuZeX05HBcw
HesCBVBCfmMQKVMNX0Arl6q/2yy9tKeQ4pc5p4o5tfepmQZe/iCkwNh0jhCb
eXsCQsuoG7EbjXgXRX64ddD4dXlxgeWRkorbRJwI+KEa8eSI/c4Ho3Sf2jp2
DqQD+wE0fzlGoNVVmpGZJ4pW2Rso+xsWRsYLcTzfb2wwt6Lu24ve5zUvl8eR
SdQ3fGuZwX67ms8LiGNsFpwrF2DhA0olyh4WYjWSHkOrReeVBmKv9WEmLa54
8nJs7owkeh0f737Mn+lJsqImcQmBRRS2dSo+WsryU6DTdK2r8J/1q/Ofh25H
rgBpXqf4vZubMUWRk6ZERzZsNuXGwS9x0VDShpmkkAMpbiiURSnZb3Mh08Ha
7geLIO9BwP4gjPyOhg0TnubP6ORskj+DP/F4L3tYsomw6bmqeBLLM+abzK4e
D7nenHdyVwVEsqUsMdW8kgreyGjCwf21MEld8dYrucLpfo7WbeuOd0bJhD21
sJHZHT0g923CsIptQYdfHKtOdnqAp/wVALzYicKlv4Ot1mNGUacSWe4PZ7Xz
PkbHIy+favHraP/YRUbz++oUxVai3D3XqMVMyPQVIMULDtS+IS9a5aUKlNzT
8+Bwhqzu9jprFFxNA1puw/T7W4IYbA/tStUK+B1eZ1xMmMbxpiEAJhz+CALf
G7+o8LyJby7mf4ENDV8dmNGAV2EgJ5/ZQ8S8JQDJTbwTNqFYz4f1z0rHjHsj
TpoQIDP5Kl9E1BIhkHZrZJfwmYkjJbkZl4W0u5Y4wPaUvxdkXtI1e/2jt4+H
s/hJ1VNVjV8Y7mp+EHTRfLzG3VIiOkU+t6S+DBa23BBNkcRWBft4eBixaMbi
WDaLG47u8g3H3O4/pcasyi6LRVaOhF1o9gMVto8YafqEibEPNe4EQ2ui7rrC
Rbp6O/FYhxtkxV2YMULJeD7RAQ8qK7DlQEc4F5DWfCa88T+kqhU7C+8xGW+6
jEZWLPmsVdm61bT6JhNlsxFWWcs4aF4wPFyFe0SbieYNWTFkg4zF+x2ls6bI
UwUHfPfU3LJuMkoHTg/Pi5Ieadw87dcyZvbxXY/s1QMKoZeHb/0XgcQ+52BX
ZL6+DcPxBBnm8OMp4RHcrXwuR97fsQmjKVkfPbFcg8P0yUoksZxJa2GLYkV1
ODTSJEmMfS7mYaloEpNPgW5/ayA+fHVhWsD1q0qzlUA9eBV6Jqj4rFdQ+Wav
q574VmoLgTL4Eu3unbWB9MiBVwAT84k44wuTfNLU1P/GzdR5DCn+e6JjDRVE
E3G9OiCXjp8GjhGuq8e9/IfGpKnw5yOzHdPX8T2mQJwRJyKLGj/A8x0C85qp
AVOCU6w/qUGphCO9A4ZW2QpA90b1wngkyQcs8o1OE/5fqhStaG17Xq2xxAxy
q4PSmls5SV+SQWDkHbXPAhawOH2JxDL+JUlO2hvHCf/DX1NDCNDsWZ//KZ4l
J+CgErYI5woShrwpKlFbG4NxQR2POq36FPYFzdwkTKmKEQaBj7Hc5O4be+Vt
pMySn/WQEevv4h34Y7nkCJ1HNEs7f2l7D2w7avEFBgqqrXacltWrxSvDGrBf
5ynCs/GYw/6Di+1/wDetMEeQKjmlB8Er0EjBRUYRTUyzkyE3MvZCNW9Uv4XV
IbVZWXdW50hvtNSyPASYE6RBBiVLq/c4FLQmnpmtxXJ1R2eq79mfa7bSPDeU
C4bHrSe5yhkuhME1v46MiY8Vf0e3/S2kItd45S6pu/LHGHDp8cn5iq3C/fFp
lyTsOJsWLwQs/sKuahw2Z5TL3e1XOd8e0HJ8WlZqhlsNXdI+P30icH1I4ehR
/EdjN3ZUZPQZidLEmw+a6hnyUqfglzRcM4gvefOIJGsv3Is/NZllbTWJgxNO
41aEKBeGWwbIS4vphCGwLQsY/X6ebEDdZ2rSG698Wn32tDC3tDrcG4kUpXwx
tq3wZiykgmhwyCEsHEtN8V98R11W4CAzWAfXsCFKjuAdOq5n83yeINLp5HQm
eLznrwaVxzhJ1b//VaIqj0+eMCJ098JrLxomKKj8bh4RLcIH8dxf3OsMH15i
nm+dyyB1Uh+lIYPa245GbQRyczBHgl5aEC7yZc5ffPb3PZjey6JepOJnP5tE
VfCW9xz1L5XfgqYH7dEr6UHg7vYWlQfTDSxquDA7RjWor8wiSLdPEqhsM6WH
5J07b3D7aOrzXKuwfYRLsbGyOgeYAcTFZPIvtJX2rLulMuj2MikShuM/Vo+r
b5HVBCu8ksxIcq6qageTCjQLYw3tGxFOyHt3pngfqqME2rLtntKm0w15n4BJ
gfNghejuf6cQCFi7g/0ZQpI0NDkdvNtknWD1wTejqfXd35+PuNjgp0UKPKm9
yqaMzjKwUZNCDxXfLiS7+BuRcUhQXutiuXHP38C3i5kozt34DrvcqkUaviKO
n1Vfh8CvopptEB2k0VLUoO0uynix9JLW8+XZt4CfYpxXpPi3ozCoCtAJT00o
TfajczNneJPUuoDuzekb0iC8E39vys+Wz6ObUJ+dRAPjO2oDZ4RyVAKdJXrC
FQQkG2mE72r0JOfyjrswe6BvJbYe3rrvFBfxRQXcg+0QVJfmig3Xn1s+2iLX
YfNuewNhcyn+vmCPRlpiskEahEvqxofh/FO5BBb8NOPPbKTwKbExc7dcpIOB
WoP40gA+fyCU8ecBSoBbxzmXMtwIqQoYfPvE5zNx7q2w0uKhl7g5zzZ1B093
HLs61CzeyQqCI3+kh7ZJEsYGzjuz3V9F+OZAdAboufdb3abLSuD5P93J6AZ3
Z12R2NLhG8D7z+A/apkSsJMgLxXQ+0p+uIbJt/rgTSo4V3ujNF0bNaelE+sm
cNELK6ePBov3TVsCtXB0OzMWtuWpPJ4DgKHZgPSDswMdC16xTGBR4jjkBYzn
XPBRI6B33xlz5RD8rLvDd6Zwr2vzvB/jcNqzbBUWD3YSmFDoAEwEz9wwF+xu
IKy+ZD2a2l9s/bjKIeas7hutQjQ1btpChhM/jotESzpuJmx+GEZoMH7IYtsR
vvYoOpETvWl3S//hvha9ZMzsbPVY9n4M4JZmOpWpn9id5Nr54NAExr298/PP
95UzMbkDpzhL/xbXM7iX2jj214xPj5VYNm3jgUrA7us4tSF3Ax+6jjvtW1c6
HdnpIhfCo6OT5zGUFsiAJhW2AqT3PzPOU2LraGktSsPVz8m45FNOW8FVrfTR
zL1El1uyEQ+DWMwHCmHhkbRl1eMx7bDPw2XTvYTRRmIxhaKN4clFS6Sv6ex/
2F2UuRl0aQhV8t7rdUX38o67Crl4j8IUMZcEJLY0HQ011H5SYnKkAKjUqN/x
KhLCQKBXHNg97e6p3i9BRfgh84x3hbn0HvhX6QfaygcKa2PM+OtrsoEdWLzE
d4kxGZcsDDXEM4eo8mm1ai7LCRDke4qjx63Lr/pYXScT4SWOuKAFrYSDVBOG
cTqZFvX6i4xe8yzmq4vI+zhVIPwX09EMZg2/c7wkm+F91ywwk89E0exi4azd
8e5P2MI4GgFS66OUxnH0DfssL1/GmOBzGdGlMRarcehJggalgy8zqlBBqhia
5N5Bmmnv5751x8vm33Pf2BAL/NE3dFOGbGpPMTHVE3rEGZaZcLepeNwhd8rV
LQfeu2v+kZxfW8dzKMrvZ5J1exp1f6huQPv8njFZ2kLZMg/q/O+EK6BQY/zd
V1K5ws9esWneB2VBAXhVXn54PU1YzJvqDQlVM6aqqIJq3SZT6zZN0TCU2Dvb
VShGziLSPebHUrkMhugJtt0apFnx5GItv6Tt6wG8EIzxvnQUaCGKfLXH/B8S
DpLyPQ8tjpJwTpKqtX0X1FM1VhmiOEWJa/o0/DjMiK9mArn7IY/Z9ox+PZKS
nWQg+Iv8+MDAZqQlyEfpu4Axx2JQyQ1ld/Bj6zIPmdB+pAX/6GJzIWcksJOI
Sr6TiCl5JMCEziTU/XFykXGb5jrzwEDhaG+W8UejYDzdx3gxOSf8ewXyVzNC
BZD2z2SZ64zmuq9DozF5ArQwe4Cncv6RQucKTM8Bl+1tzZhk3PKP8eQxubzB
vwN92YyeLS9KxBuIEaP3yCsN388XyKZPZch9887ymzhaz8EWeleOcP0+n6ca
mmozaz+xp+DFehfsHcJAODsfqkfvGEADlGN7NrYmZ8XgNiS5jvynh7G/oWAL
rn4TyVyKGYEpnXm3MGu/L51PkVE5DuU69r8jUdAQTQQNO0oNPxAoajrNooS/
xIZwZZBhwqc1jVf9cTB+YqiW7IeVlWJM2ZWcocPutOXTPACkuvS7HQt3KpCP
v0isXYqniEJj68kFjoTZe2efynOEStGCWyFZh0bsPE5FN4mJP8j9rVv1VB8T
eNBx3pYJiBZH3mD8qhVZAFnJtabQmknf4cWiyq+gPJ4Mht6gglGxrvx+lOwk
UEuq2lDOxiJ414Lg4pMGDoU+Pc+Pypl61r2tHjePWrnZpuk0xXuil6tj7IWa
It+rfarwvRaOrBILABpHPGG9tc+NUd/AN8aYbo0WrziFt+NDzVRoqnw6tatF
RiJVuULvwgFgHoknKj7s4dkq90ysChEcwYTf6YsGE+/IuxMZCP3o2HSnSVoz
FWmWQuv5/xAdxRDkvfr9IKx8ptM1NpTP76cd/RYR2nKRU0LQlOeFxzKRos1o
D7eHMA2KeduBlzFYyH4579b/3dr+eCflw7RD6DHQJWKyCjAmuyJGH4C0hW+c
QlxcerqsP+D06zkgtQ8NIa8Kvn/tUZTtYOdL0wV4SyAh1YA+ygeY+XrGvz/w
UAcNK4krT1kWkc+Rv0xhsA5FMbYSd4J5+wtsws9LdpHf6DFnkNBtitJaCP4e
Hp5OtOH5qbQ4b/DBgvZwSk/PrNZ0sUYEiEpESAi96AALzdXKHc3ecBIoRjw8
F89z6Aygl+byV0HLzVvRqlTfxLJZJPNG1U46BkkqQlQCiA4YYgVFVENu6XJM
BHNQoFDknDOGwRjzZYj2o3g+KZoinm//ZAXw7qAiRGckiOy31NsMk1htp9Jh
u2QWLFLUAndz1rwYvzSFAG2HLkpIJnhnTx/kQxn8WLu3p/uUfG9GH0Nnu+ev
EJejzUix4yndommyhD6cV8/PpPfL3/hiuqwIvxZYs6wRhlw+STafGoByG/AP
JFoQMy3hX7s6PsQzRpOaY7HbQ94NLZuQSp2AsUEbbzD0VMdGjBNp6a+qCoJn
gzXUz9DFs1D1Jtqq/IIW9RhudVe1WOaKJvpCE3yGSy173gxX2l97hhptc+pl
GyrUMMXTpcIc1COxBhyoEnAZS2tImslM5JYXtQ8e/0miAg/kgN+xBH6/6RJk
A9JXcBRUiHHk/SV154ntbr2pCn/GbuIyuIYI/0fTlYLwxrEXhqRdjEa1DSWg
FNacCVB5mqXjex7ICcrkCXnU4MJO5CDIIwn9yZNxKgUnawuyvDRINWzyXAZD
f1Ev00C9yOgHmHDFn7RITqyaA8WmwQ7Wud8CclpAGNWI0KbT3v1I6UBnAzXL
HWEBuhdeX9s04MgQ/5n3OhrpjmhoW9zzgmfZXJFuCSDIKMv1j2bo9smKpe2J
BbXd+TH5ecgBUVLG30VxzxXLwhm0BrFTbsqH/3gV0Osm66WQoQYMdlQ+XlLG
VTTOyFhCbBQMIF4/pwNMtEx49kSPCs/D0apnZVPxiNM4VLk+3t3O98lJMuwT
M4EXpAqZ2djM7Yl9vKqk8o6W7gSOWT3UviiIKrSfRrihWxk4zT3PTedH0M+9
HBjtQoHWahRi6T2OD7OTIvObyPb8zO4tKi1a0QcsVy1QdDsq/WMP/SbsqOW8
1jlE2NEX7A9tzXChrqAlZkQqfSyrezEMyRP57pLeabWE5GXBLRfh6PfrRD4/
ZM+/7znjsnj+Jm/Qq+Rkgbko23QRHG/BSjA6AhoDvJbD+gTWK3Ch+RVSJHSm
ByfsKZHTYPexDwobnMR3j55QcytzCA2RnXnOCYCXUpwjAfITuAffUcpVjEgT
y3CDxJv5oZjOfYIBzN2Km1qTqlcPwDqWzG5tXGSBgGIpNKRmVwOiBi83jhdj
B5xRHAjRGgGzdMJLOj1j84UDBxCO+WVLNAT7gYyQdcjyuKnnu2ouq724Utso
dhZKcjgYU9RcMcAI22KjHm6lbwMdh7MvsYaOa49B1zgorpcFsO61mo8Te2Dy
X1szYeseBQBH4bA1evryJDew3wfr9H0M2KftOwER0h+dQiOaUzU/D5g8WHJ+
fLtRxHwROJ6ORel3v3I++blIv5c3F6jAJ8Pf6AEPNre9AlpZU6CSegeJQxT5
s1r5mHHdOedJEk6tB9SlObd7RZCMslbWgN1zrugqrKQduMsA/bS4bGNVmHV6
J+LKjG8SdlJyaOdi1VnpspjWk5PVupFYJe75yiWOLDNQeMhjveZ2UCcJzf49
6PRLZrAcCPezgD1IudDGopBa5N/SfxGITmhv+lOPhOXZFL0GYygqJbWHi+5e
gzcIYte2Vg+eDGIfO3L1WporThv1lc1+O6oAs5X5TqWw/MWwExCRPInXORJi
2ZeJGDOwi79dCmzYAXrATErTy2o2QUNs4sjCu/t9HjpIVLV4BqZYPlozcP5S
DOcto/s5KTfZP+kiRhxA/R7OTi8gi1j88Qw+CBxNG/vMc9s3kulBo7hz9Z/i
UOEQW8r2I9L4LXh0k9m7g7AR4602DDOUi9IURLod//ybok0iSiHPC9MwklMd
KIM+FwXyzM1RIRYb9tHcXBQru4pwn7FDJmplYrWq0s11HIWYYR353JF9E6ea
4+QR5+6XXdusk59twOweIL8eVsVqtsiz+Po5/V6YkPgEx5spnschi3UHJCoO
q28N7n+rtKxhnik7bF59odDUJSwv9eL/ED07zNg7FXQaL4TRsk0fxDKoZ6El
uRP389xG22IZSBVmC5iVNFdKyOijE05PYef8P4kSLDvzGAmXFmV5VMhXeV3P
w671y0QKUydMZT2lNhsmkVXgLFH63zuKjt+WNyJMyyRwRveKjeZwVu8h6dyq
VNKaXyzoMuYqJUL6KGE1i5Aew1JnAGG9mTZ6i6A0XtywUxXX+zwSdGJNCRIt
C8mFr9jOwACNhlMfphlV5dTtCaDrgqo7A1uoySYAx28oD2z8qCF8tqlfiZC8
tlgNxhlzvSgNkc8r/RQkddSOl3ikXBaWGHsvByZEWuNUJydkoPpPIhrxA94V
gGXFXukW2kh8Cz7K/5gWU6CtfXiFHw9i+SAlXOSbKkHQvT/r5mUrkDosjmrO
J9lVdX9OotxXLinWp/gPS4EZFO6W064GfMIxrMt2v5sP7O624KCP/skS1IQz
PcldN6rHSLOmMdSYSutxzgKNyIK1d3VoDmd8NlqUKE78GLiJ0nGW32uVe07W
AlhPsRvK8HaMh4XE06fAapL8ybz0qEqOztHGbr9p6XhW884XyiXBv2LxKiIB
N7B0SP6QWFpVwkixwxqDVZWFs0bnm8xP48MKvm/vdWAaKXKaJ8wHc8ksoOMJ
eb9oI5va8wFaNQvcJ2qg4MNwXbEWo4TcoNIDkIgoJjSEvu9556mh1EvJnlo8
9Yw7+bSdpCK55Isqbnjs8DDyuVPErRvVjzAVMM0gEONpNXz23ANjP0cgQgCT
ktqTLzrFbbyMx4umf2FQuLEwzyxkRyKvLinBiUMH3psjeOcGlstdv0Vg5JJ9
xxIhChChgPNyXqYfvXL6i5Y6Nj95d+aNOHW2CfqqxrwFWgHymuw2SI1A/ABt
EJBT/9hW3dwLyEpDpyVP/JduRtomxb8mVDI5TuO8bgNdSjB20JdY5vebl7bq
4rqzJ8y4HKOvWIKmhkokUgAdADbYVlONtry1ezYUJfJ01vKPr/fSB6IvKiIn
INkRvgbEMpLWU5isalB9xey0GUzbJKfO7m1u8OCntcjjnVZoItVHEMVpsb10
o3kRtbUgVUdbAGIxt8mOgTqPoqOVSY1T9rOZ4GeHvCHA4hipZ3Fq+t6zSL1I
6lZ0stgrbSxbFky68EAahvaqFPMuavhpYqOTY15CrzMPUSyE94oq9JGgIEX4
6bF+4p9YATjIodeZTg6gG6mKRI7b7QceY2pfJbIYvgyeh8OxC05htTvGYbYC
SMu72LhmPHDW/pap0/GRrXNrVSLEAQAbJ/TbB3hgEyvgnUYiNq5kWJu1sUJu
4SnUjbHNkHNeJpBUWmFLSQSZnHTys5AIgPnk3sxMSILTWRNEqcqrBc6cfi4I
CHoP3C4XUBXBLoG26Ta+BwjmwaBquNtF+xEnKToAbtMPT5enfpo1TQE5xp6V
Cz9P2e78UBEWgEkLgOr9Po6x1qZzuF++aBAu7xaW+cUmCyXWuAnXLuCe+KPk
ls9pb37SBEnnONYN7lB41iS7v+w9/yT9Z6aQDoFFsn63gYjf+qiERfrDwDOs
C1W/3YFv5R4HbAZYu2S8IVnMaX8hl/+9KzsCykey5BfIFqibDgBxxaJjj1FU
ABS9mUBdFNFsvGZoVE9m2qJlFv6uLGaqTa2maPnpUMucNP7AtArUd9vecWoc
qHfTn8yIt7b5tvTO0wxzZD598kOl41pjEP4U3+RklPwu6TcBc+Y5Z36mOOT3
bpE77qiSeoJcnprLubFaCmlOq6mhpx5uDWMbnUjw/4rcgN9RhtFjaBnj/7Vu
3KALT/eOwtTyW/VeMHXawjTcOOUzr1Q2h/jSwTWdj5V9XWxIR/OFaj2rfVRR
g+D9h7rjgIbk44xBy36qWdTx5UdDrZSWal8EBRPmSW0W66+qwCCx+3Ds0qde
j0fbx8qZSAGDmOVfh5PwQ/owl9r8vDSIDH2OpRogrGGbKaMja/qsmKorymSb
T5KkGqD4g9kLMMLL2MrwXP3fYfSey4ycCO55k7UBk+fmDkH18VwFwZgF6OKX
pOH8CQB1beZuaatgADdgjEIMqFpguWdnqLAlbfIxFlKaEW2ejCetplVmgrUg
I2Yow/9KlZkCnWQoh9usLjClXZsKc+GPxKAGGPYOjdweGDLMycYol9EuZsAw
MOv9NiNUuGN4gdDiO4+QsUZfT30PVuXMjWXqTi89Fp59QKQu+puymkWGqIQ8
/8Su5cGxtrTXBwvel+QNclgaQ2lln/27C6/lw8nnEE+n/LK8kgbLb40gJMU+
HF1uqryOaiP+DrLa2ikwTAdvhHiExIdHV0AuNByK7eoY8XR1KlfLUv0kXXKw
y3Ru8PwJr/V+USct9TktZKdU+N2KsN71DGA+W606kTecVk8S3s3I43wCmHqS
7KYnngJMO14hwyt+7YbA9Bv8gDJSAgSYtHpkoWOM4mBMF/pBJZPxXylHn+n0
72ftVU+3+Iv4EXNLPzuyhEvhlMNz0liP1T3FdqWsUxwELfddVt5HW/SAkF2L
KgP/fRKI1qVhOSJbPIc2IdhHn//MoQtUytreZ77/0JK8VzMv4y8ftJmWliD/
Mm/G1ZnhdcUI/1yK+/1Zms5J76wqxmHh47EdnpeaDVrWOjXexUuBCnxRDldF
MAB803R4+xzXUXB4HfL7ux6LDThoM00MVSTMA5UUUBtlYoZ1lgTWu0hImEyT
O/zRqNrFJDPsWpoMs85/nPE3v820LZj1T8s9han2ZVcBpEDC+/0IviOBVveC
Kyh31b2OBilozvQui4ZHSV+8KosVI+q/G8khGizo8FP21lZ9B135+eb4VG9w
a8ZoXaX0+Zgy+lzBPyferhfijeW9IyDfgEXaeUtoUvxeuPjy1nR5Mvu2i+zN
2e+EPCkeDUE4Shzv6lKueAfWlhIe5IXAlvAXhS+fPOGVoAZkgiDLyhyg9v+h
IrvtPcn8X2mK0TkEfCAkMcIR6BCm4MIwDWmYPFcNVXKlkEAU/B/cJCkCw9UY
FgOgYNSEV6KrK2mE7oUX3rBpZthExym2ZNGNfsQELINPbZLKMwZyoNBfVF4z
BRwFraZ56xl9acBJpglpJaftJZN2EvuSEHCD5he6VCRXpGhTGET9JL7y/kgq
g1ta8kGferXxirLRxrHJP5U2CMVRWHdw/bvW0DDQAOas0Z7SooCbrhhUJV2l
FPYDhVGuacJOylMnF/IlkcQFEAIUfOPAKvGN/v+DCuhDGfzR44w1Vd9WwX8G
GRcDaZbXPhthdTAEBpnCr0dAwqr5BBw9Wi3SFOS4K0fvxfXksJwKB8hB+h6w
bc0PGT19NK1S3ZVQIpjNJ07qxMihHemj2jDGj3SVV8xK94PGDQeYfCfVP4pO
ofKzCTtst39fYkceLvk8ahZUK5DjSs8sAkLjCtuPz06qg2kELKL1COC/vNWp
Tu7MgHNisA5inVBPec7h6PrOS0OIiv7bl/BdrsOAShHD9Bjxg2nxhTXepbAa
hdC+iYV2rgruDEq7MEguqMr5wvfDFg528nkC46lHwl30MSQ/4yyNsc1qL6fG
ctUFAChsy9dG6HGsQO/9o2jR6BWnXYvDGPeR7Uu+9WhsA+nSpAPyVVYlcc4Z
xqyWt3+1Q0Ag2T3fmKRmYq7JRoNv/u4vQG+Yrg5nE7OB+mNxpUR50AjIHMfG
mBiyp+NcJBBmGvX1Yy8BYsO5gX5j/cOAZ+90AsHWbgFw/f0meXCa2/FOUA/7
3ZRdkOPAjoNFgmSNPRS/3U5uD1hV1XKot/xSIvm4z+f9PF+YWHLz3W57ZQsw
AEVh5IvX7Kc4EK/BjNAmNY1RYCDZuM4I/mDPg9BSI2p1AMqAxCXBrTHF95WE
cUd8Pf/876DNOBCC96BiDt6snglwIxN8r3GD/ql7PbsH6HA0wxz0YEtsUqCM
jSAXqH6H2h14qcQgoQbHH2OF2YFBx5xyB+vFEGayOr0xgpiLGJWiLC2/jDil
8xenIeMoAkUx72HJpAKUknEtO1xYEPBxStk1RBtt+Exu4Ms7gTJIL+Bza6tN
2u85rRqLL0vmV1zKwpNSbqVOJpGYFOw6y9hpMFpTb3eFpDuHl9huFzW8G9/F
KwHjAVFJ5wxmndw5HEDQF9uc2ZD7BmqfHz3ox/DovYrLNX2vsyKmDcohW8g7
XvthfBOxw6mqj/Vn7GoplFA5SYOJgYOfn3focSj5acGLOsmZkJpO+DmVDFWS
F9ZG6wLii7vhySccqpZpnyhraA3zL0Ji8rB8OYvWntIbIUzboFFq7CmALeOu
b0Sr9HGtYwvd65XWhEF7mvSRunWLcPGMxMutOVRJxa0J9nxDUeLg302pEakP
+pZzX3g3m7RqtJYoEuVnPTRSl4hKP4CF7n5gJeq73uxF/+wpWle7LMytS1vb
Jkou5gyI25rEe4GG8GW/fh/kQgiKqquktRIKznOPKHiA3wzM/AoBsWu/QCST
Ecltjzlxg3cQgXhmaPo7Fvlb9ty9e10gUbK2L5Bfrj+Sta1vM8YHcVJgmaWe
K5C14z4sNAZqXOOiKoAJ2S5RXrKk8U9zEOYmKvD+xDeMmqujJHPbu8JWKQX6
lll7NTLhSZfaRjg/g/vaZJ0cCne06teHsdjLxzz5TwQuThVRZNbA3ILVMkZT
Qca2wsuP1KUVh/8TBa4/0i+x0CtK7kuJE+SOtWfK4yjNpQn5vqKqlPji4hQK
D9pyMyWBQqE6PHaMcf/+ggP9hONjOweMi+S83UeLEnUcs511kJSaplyA1loi
HbyiSKVGeuOZPQNWKYlg0trH1kG7PzDYb6kLg51t67lgfl7EUwXBVAJzYwjr
cEGmOYjmD0svbsyjZTMSBJX+B9hRkrUzGMBXawB2Zv0V8xDgPqqHKGmMXef1
5T/RutB8EFqfgKY7gfFfW3HXbeK0tuuRL/jcGxN9KSjklc7MsCg1AuK533Uw
/bIUiNv/pSyf+nqw5Axsb5FnfH7Sxk9J+TMMEH+X83b8gStUcWZzMP6Ziuw9
AY9p1N3eKeXD4PGDzAmsGdMdUMwO7/6dy92L3eJGyFNHoIOEpu7+t3nFWwKX
3YdHx5ZRRRes5Hm0jFNDzyUv2e+A1OIPEhC6pLJL5JwwuQflNSDX89FFiN5i
YoN8Tsm+6nApuFwy6x7wVqKTuswpiQ2HjkPADxhuV0U9vdiIv3JgSGDItEON
JU0bJ1EsrdqOJj8S0E8CV0sy1iwnjfgOSBPM8O8H0sO7VzcVFvKY6TXXc3gQ
hSuB3hOa2dFj4nA7EMSFVqvUr1ESNnTpiD1lllMB+BradPRnEyz/PZQpWKHE
Sz+R94ZcLVV2edWHsLMl1jUugbenF+e2AX5/ac5uAtHXiqDOx3yH1QtYTvI9
md+gAFTGC24F5TaqQgTfavFnHSzS5XHQfR39YBy+V+3uSCb7v58olq3v22xW
/4U0cbBrjzo92FAlqdHeO+94P8fEhcUW1hnn12GtsZOPWNHYIZPdfKndz48w
Tu9SEQ33OPtMPiv5CED9fUwQ+TAPp85I3mPylbnR1rI2RVRGaTiRR+e/5cm4
Dj/Zbgf0Vsucu2a07yc1weWhVjRmmHgPPfdTL38DtFl3OPs19SUHv+0gp+/g
LQpRHteCU2l/5nWvfiQd2kmNl2Km2iwtCRsD4Gi7GqaZnpzaduLMNG7Vi67l
FE3qsonnfGmDMmmxVuSbKZ3FZFczmXNbXC+M2OkbThNOeCw7RlcXg/ygATBA
QMej7Vl5CP/DIX8jKaq/kKxbEB2KPA7CINq2x/maICWnIB+k6CLycyieN/yj
mscOhhH8+Qfp0NLf5ZrM8lmZ3rsDsOFl0774O0aCgBUUOvTsN5/fCa3uv1SN
kHjmSB20yYFmmt1B9MD4KJkCFYgl90FNY/12ybzjost7ZSe3Za3WSLCvSZdB
zGrLwpr5ePjpalBiTp28qEuuugnW5AIIVgqwdqYxWEL68bLiqz9m0/noi+py
a4aCVBAm/K4BVYtjpEtk60+TvpIyRxGoGy9MZJ/oeZ8vQx6Xwid8FepG2VPK
5eRShICDMXAhLXBiU5prCK3zGsZLQvFCHMRbuFfQBXTHAgjIeSAwGGMO6kwb
tDAVuFzlV80joKqAnnS3VJlSkKWkrP4eYxaHwASt9B3kGSseqVLne0PAwS9t
l2sTkxmuOiJX8urjsUpOKcRzWtIsySp/x1mBvDEjCA2xieLifEgUCiG0nkgW
wqAJbwY/6Ryy9b0IYGmN6lime5gBbOikB7IZ/nV8QenNGPX6tSTxK3m/qxX+
2twjZemrCqempkrXUpsSZpN44IfNT09KFEE2pvBnuVRLwsO2zlZ1OM61QiqY
PSSjBcE0NtTGvGsmVGTNvLF1GHEATQRN9WyOTPTnaR0KlaWvYBmPcNUyD04e
0ZD8LF3e6E/gPFOSJ09KfOYMvnNbIz8fF1IIB/F/LCvQZa0nnShynvAEAjr4
nTer1MMIAMwnfkG8CHujurvEl4M7GTj/f6bYm/JEDmaAph7neQ0jwaTLlR2/
x6t60NZw5VAPAfagLuditSWj9Z5LqKKfP/kZ6Jpby/K8JiGNgjsoFRrOHKXe
fbljxhj37o3TZ6QKBWNsC1SOB0cBKBiouPwExNQ1PCN4nRQcFCXowqZBeRqH
ynXuAdAJcnJMJkLmJX3SaU5jcTsq0vnTRsRadRHJ2S6pUypIbakr/eFrnxx0
VhqTjACB6G+MNAYJuqVT10RiZtx1uF1k1WTQ46PLAFLd1tBHlVsWBwGc50Gc
fBV/eJmDw7DogJBnM3zBGF49pfsCOUDWGKSZSHfiMNekjA0WpZRGa+/1NKiW
xe71GqcRdrArrrUoWlRJrA5f2pH0J7+U8qI6VfbNqyPzWAaTKAM8GNyL2AN/
HxTN9UwqpImDET5t1ks7w4jO7xuZA3o8S3IP/Csrq6wk0v5EqlWhqTQ//04W
Sm9MAH1R7Ze4HK4QT4NUaIfuvxJ2BhdBUqCN+CW1fCPeJCHaZo+OK7RFxa5g
uT65gU+OWH5aqQcCXTysWSKixNsQhc148jsZ0zrZ5FgHvD2Db7rJnkjhPWHJ
iYctJEgdbu4w4NKbJwtWLX7IVbc8pP0oAvBS0Lz0TDLOMh80n5ULTYPnhpEI
/9giinZDVmEKi3cGCWYJuG1QGF6SQeM+iWFH7o1IR9QKC8/1MYFvu1YZlJH3
w0dwWg7barhrlbctnFnnxMp2i5Hgi9xlVxAfRW/ocNglrptuaWRu5lfIgjSq
pMOgct2rcr1rDQ90jHielk7WGoo7NK23IbipQFdlXag72Vuu1U2L1IuMh2rA
nHeov533X06a0cSbzXwCztuJPW6MqkdC0UTZTEVWrZaB8gZpmsdHocDOcolK
UNPG9pl25MEY9ZW3Ym+nXNRUdjJFs7hSHDqKZmdKAMxTRd1lA1aKcq71U3xG
6no08iMvlJqRJi+A8Td2mBmmGomXNPCJhkKz7UD45jYdBZNTQH2btoctcFbs
B9vIkjsC8uSBgvnnYOt2cuIVeKE4LD3yjfQaIbtrDmLYK2sSezkN8gisT+gn
9udUdCQo1mi8oHAMK4LZ24bQEW17VsvDb67cEQwU4aFNxcKUE2IYTUSOAfGB
cCIHgenQo12rB+iHJY0lPr3h1zCnpP8qa8Uaq7M5z9HH9ycY9ILWSpI8wDc+
0b2xo4kvS13ax7ukU5b21q+5M8Cz4phGF1QpfyeKpiVCy4Wt6L5RBLJshjaO
TeWHkEXpXIM3vRuMIsijzzp8idpaJqyOTEzeFYwQ9v8T+JZIg8ohztGR+zct
3OuNVlO2q4rpqs8kiIjX8KT6b+SkXb/6S+l7thQnAWOd8SBm6L2CqzKniU06
+sCAok8nnHQv49qttLhT7eL7Z/vhyz71kN8ngSYZ9iHYWtldPQjuMLGyERb9
I9UM9oZ8731XYpSJ10qyf+U/0Qkz2Ovi5ke/LYWU2ZIchXVzU1LS10DSgwM0
3KzgE6YZ2D+t74CCD7VLm7cZfGsmku/YIfKztgGgsujpD2wDDWe89eClW9Kx
ci8SEj+7R2zCjswOf2k+l9MvWHUzLzcGSzXXtv93xb1G+qBPTPx7CFLXeUfz
RT65KjX7dZZ59Lagqn8wqIM04pM18rKMXKdERg0OVrS4/Y3olxC8at4MjdSd
M4VskI3Ka/Op6kAPgGyzv9nDValfPUvRpp13Cr/CaaWfULCSSYJrPV1qkYkl
GMHTlOLfmAW6Iy82lKncKUrMnJZ9LNXDJCCB0IdwAGMZAH4InBDnx5DuDAeq
pVxorT8a87mLol7v/vnZuN8aVlUvYXAeX5Fy9qy0te7KcZekMt4t5l2WDCgo
zNRrDx9m2YeEWhoPTBeuofl8VOhRiUv+7q35u1awzslPbb6hnPUUl1A2ct++
Mgto90tdwsMZFDhma82sLrHjZpDR2cLePWnF5gjxajyRHdGXxdLWYlsOhbr6
WO3hOZb6ij9j5TGGyd3r9Aouu7Or1gHH43i4J3ZgHvr2k+M+pFpppwu8l/Ry
YACRrEi7KQiFmiSEscD3SlcEO2TyoJVcdtLHxBZkKrLMo6rqidShD9PKJWZm
nv+t/uFfEnUwYGtvfGcc2oBg430L0+qzb+PywVUWntP8kgBUrEmUcz7bHaPj
W6f2hM9Ime5XQl9WeezFlll4/FJZEGKtSxRIh0zLD3qwk+v5lstSH6wJihWH
JNJlSQMIVujMQmD91J+wxhOaYv6OiqQWZ5E22Wt7cI5L9J6P5fbURc5QZ3z9
AschNa8Gfy7b9AgWB3jrovTdR7I8F2JkXK/Fn99zWY2FWpx+fRUznB5nGuOf
8+xrGiDhubL24lnJ2PglGZn3JKt2+6Ir7JAdwtZkFR/2+EF/H1mvb9Z4v8wb
EqJnyQxrMULdPr8iY+Qn6J/hxIkGQfPGtUG7oiEXPsdeyJPusfWQc7gAXDoG
od0brg3Me5GyLI4YYA0eSlNaGZ11q3KK3OXu/Yv1SdNAGeG4aIBLdRB5r+c1
nsKzNKnzV7O8PLPqMWl42qo9DHPYQpYhEKYdE/EhRvxu/PQZCV2vEuw/Ea61
P2aYYWSI1KLv78H5SVlSmDj2JYLa2iqEomU3rTv69e+jk0/YbRsICWdwUnga
YARq6vbXqq9uJC95+IOgGX2XRQq2vCq95LN8Ks1/xTVk7FdUvX59Ectp/QkM
PqIbSnF2s/VQXpzsphU4fWBZHxFtjIK27qUM/N9RoW0skrSsSMAklmBSn0au
Xa2ncuKtE1n0pL6imkgGD+G+hq28RsGmFklQTy0aqe8al3tIrDeZUtWMrnas
da0QIrjd4yxw0ZZbBcxs9owzoz74WfirAQquQccHyYh0CAcbSiJUoICUIGyF
Gs+hqPX0XmuBWRZInRe7/N5IbWEZ5RlXGvPNHbQIZ0Wui4CT404lfLbf1aAd
hOmnNUBWCvof+cYsZTTG9Jj8ctnUywidMXahix1QlkyBvVBLqHZL+k2UNXli
Mz4Jmib3KFUlgQ4d/oJRA62OzB6biSL3NvLA6tj2agvRw2AGLzmf035V+O15
z0dSGHM1Lq82G195ZYLcpjQZT/YHIiQbnIhK7lbjenV8UOE9K7vGC5fzFPs3
JGe4nSX6ACPGmnlDzzcMYV5dI8AnFlWpz3ftw4D2e25d5/JpLmRa/8KDKC17
vuPRRRmTIvIw2Ukc9PKl0wEAjvDA96f0LErm5l8EJr5J0PRRBPjftXZ5vc8R
7C1UF/wpVrvAxFCYhNeYu6Dj4+aEnn3ysySaoeJEIhgvWUzM9adI9D4jLIRA
moYu2Kb42CohlMc/HHpLfxrHQe0w1fdUCNnbPU0UiHtBMVyrJ+MQw1b9uQzz
SwTy4NyFn5Tbux6xubWL6f6BNDh/9DL/c/6ab7RTjEr/5ieJcpCzIV7Pdrqa
c9y79Q5FTq1lG9dAnn79Q9VcWDJ1HnZ0vYiD1eNGFYgFj9PFppWgxnhZRKG3
rLly/BW6Yvj2GhWW7ITy5F4Q2b5BxdqiaOlau+0eUWIQoCXaGwKbGo48x32+
8jFSaIYwy/K6mBHd9il5TuNv27TxLUdQAeUzyqJjbxUedv3EkcC9sNQT1J7m
RyYaEN83sKfkQh5P2Nz6cjFXzyYaFkkJAw9Qf5Rja88PLw7dOkGU2OASdvkA
R/9m3vW2ZPO901g20GH7bf8nXd+rnZYSuRd/HRj56mfx0DZEx8DmWLxMTWc9
oaWjd0PgU0AkUA7g5sM04mWdPnfjzgo82vSKZdAJc13Yis/5s7IbLYiG+VZ3
5ebhPedyMKSMEGnNbnrE8QX2mQ4l0FPoln8Qh0JN1k5ZTrppS55LLaEIaUwo
o9bWX2p/syJUONFZEGhsMx6hSRa5kruhXclO/sWOrRq+kjyg/Oh/6nyqWP0a
J0xW59R718kfVt5Ac2u6j8bKkrzbY2Hb1TB7EXDlcSMYLzQ0zTOGWF0I1I0P
LdYEoUN1xuXJymUF2juZEF4mgu2yoJRr5Sa0DRRAsB+zf0pSG+gOhaJ/TrkC
yjC+UCfhMaya8kfgDNtHacuKC/WS9obLZP9wxRkaC+tHcC9pzUczKTIz7oWD
MfO7Ws5VIL0Sd/FCt76T3nFEcZiBSnK6LepwFaA9x7xG8OiBiPGPpwfSSTuA
pDi/eCSqowtFW1S23zGjH4givItRj1c1CIdA4iGQ7oGLU+O/M670JdQQwOY2
IsFbxfk0kQ2YMxQHmmP0xhx6v9ItvTCkyJiW65xOg1lWz7bnv04wbApZLhdO
gFTmYN74yBbf/l3MZFngPk0wXI8KULaWi/gjii8ui0PKY0Alnl0qv0ThJKfT
cxYljfRkPMNbi1vYQb9xM05BRVQpraNRxflLApC5824i22CVKz8gxYrJJjXT
8saXHR0Ez4/+M1hNkCiYWD2krAyvWpijGDM/hNEFjAK2aVlhqsbxUuSus9vz
nTwc/DzGUVcaEJDFxImhtNyL9Vgczqm9b39YujDnShKKr/DT7LiSkqNiR8TN
2Zah8MvFyQScrDHzEd1n+Obp2FbksWHLmzepkRCKtRCK00Wf1sxXU39/5Y4K
gHJBXFnxY4FbP2mRTIutSlwX0DvaMpQ15YT1puxrbf+55BWTKfWZebzUsmPZ
K41jllGpgfo0U80SbvaYA+wTbNAN4mg76dRRBQa8x2jH40leanjcul5HBEKF
5DLV67CTqEL1m7phgiR7PHtgjiWzQj34sLjBAZy61DYHfwmsqxmgPECISstg
F5u8TT4QZAmN01fucGCmTi4AYI0cjR/E/ebiZ/uewrHf/fSYtJ6ezu0D11un
6U+Jji2xMDJ7TlXbHUEG34iG8Ut5RwTv91qMpppbiUu6JtL4eczy2ADEzhJK
BiJmSwGYJzQLTTkJ19CaysJr1sKcU/sF/iVmhYiidqflhS1Jc0awNZtZ6qBB
BK8yXMlLMA24GPXhoUteLaMqF0flPY/vClXunxW1qWhHsuTn65p6tHDQnk9A
dfbz4uYKU68eTnGqeIGaxE8T2aVzacH6WVdLQzmzF/Z3uGFtoXvaqlKNmPvw
EKIMUJx6iZBZpss1poN/XP5rQBUM5/RlgPUoWwm8oZBYMw3uhMy+7DNnB6lG
sdrnXkm7dmzeNYV/AthPI+1cCkJMIt3sQGGAM+pue6yBiApxLrX8oH6FFmLi
o+sUMWjG4b36+JhX74QpKJVD7GpVcJZuJWmepil+Li3mKRPhs1YrdRg98Pc0
mFuXLL69i5iQhGskpAVeAgomJKHcdFaVPtKoDp71bSH87nqQRHJ8m5NakFGM
ns6uaZrYYrVXZ3Bs4/ujavNdfz/sZ1W2hcS81l+CN5myzhEfZ45JfoWFfagi
Pz16JD5M8Ay08q+FeC5LrfwI5tOABhPeD1XCcwOTh0sStP1F385G8dWqeaLB
gqGAK7SSkB9qRlw/rDbj3vPiR3ivhTIQ0ar0NJrWn9WOX0KawrjkWK8huZoT
NXxjju4u9xM2M1zyZRIkDUsUfnRgGgmM8gWdcEfUO71YgXL/V7Xy3NNr5iJ7
OuumiW/AAzRRmGx9MZhl8mBmlzPRtVIcqi9aW+EQyHoGXLWIIps6XExXJ5CP
J3vhz6ii0pyYpIF34wrXV0LTJm5nnMqC2FdGLqDfkbOkIjkUjyAXtGUtwj96
fzQg5EFwwR8ZYDxuqtSnVWFlvGy2aYdpogXu54qeksdV9kcJuAbV+ICI4uNP
rpSBCTRCHp+KtCj8RsGJCLNJdV2UFOS7Aop5ZEukR0QOV6Tco9oBSCSzyHUg
p29J+5/Q3ohEIWNWgzjSxk6rcx2YL+st99CEnWVaUiOAPzDfcfCmXpI7qin/
p/psyEY7euyc00d55/BKhKtf/dFLDg1tMw0bvU/LeUrJ45+mkVzJHV+dUdGj
uZl2peKTAsKrkqcQ/dvJ/2b/dd9P559tF/oLTyUM4e6DEZOErlH6H52NT6AG
XyFvA4LT7dEsInn0dv2GmUtERpJAFMyrg471p7xKDplPOzgk8+sOr3pgUxhE
fV6enVaC6xYH//rjv5TkwU+WE9q2xkwpdiYTan/F6yDxQ6j7jilbf/dhI1fW
m1q2N3svlT/fZRDbQPK8zXsYepVcmHocmhQtm60nPDg5cPgnxQlon9EpOoN2
k7yDIgHKVyK1+6P009wN1yrCQenTKFgVyAFs+UQ3tMt97tt/LLv+VcKkoKEP
D28WUwq8EPOrT39bEdbHMe1TsbwUGxEOO4zb12LwvTi/GnRHEQkvYvJBme+9
zF0d20oYFDXeGTvqDM+2t9eU/PSJ2pDZqEMZYPWBR4gKuUHX+tsZKsTRxW36
IoHEGdSvBzuxeKgTRNGaaS9LSzdx7Xci8eM0Fu4Giir32pYx4aMLg5rM+oSZ
TSmUr0pDx4ch7wuIUoAYuAesrVTU1qWb96jrd/LNuv/xYAPTMMqNrBXlJy+H
dmZxT1DVykH3uPumy3M1AGdOen55hwNU9mCLcbc5rF7hYeJTH33DCLdhRsEn
3VSNuXWauVhhRPO+6BtbB27gHjoT3CIEbBmYhVfQIz+8Zq+9WroF0xe1YlG8
3gGAu6VCy7XEquvMWAYgdEA6CKq8yJxalD/qHd73AqUcnfAlChZqhTKlbjUc
UvxXH6ApX6sbPF4Tq0s7YYz5DrIW9iDE6CDF4Eu+zzN+REVri1qa4H7VNRsp
TS7o1AnGOXxg9ErIxIM4XTHxZXddVVBYdBXhiOUzGYWhfjNvLktuQ5T5wq1s
hPWO3LObFbVYDdJUIP1BUlrc+1OlTtuyajqLx+8UrL0zRzwxz7HHsr9eP0iS
MeQq0kpniGuxdN6407oB9ogHgglQrf8s64rWWhy93WlMTrndGxq9aF2W/bin
GN8sJTt3rCq67q7aCheyLa6EKEgdKExg/qGjdT5AFvp8TAwKs//CzfcK7Ces
mpSWwdvz/tCqzkXxAIqa8IGFMXfZ0taBsdlBg0PR29J6cWPrspWeT6z0Iyhk
BxX4R/Ig5C6mCG5YUJBNDww7hz14IoGtEGEINXXRiczTPhetVG14QrxuTOmc
G76eRwBTrTrlJlSQtLDtj216+a02KZ3Eu3gtSUYze+5DHLh7qMTZhxiPwCBJ
kmadftadb6Elym+QRbtlbP3FWQ2AmqNBxutIuZUBZxygBsn/Wqhehn1qH4hk
xx4Kpd8qaDl+l4miDiix1Z2RDq9cI6MRIxji0HT6CQB0/49cGfiru7DZG9vj
GVIo8nGKmP4O9Rk32/9Fmuv6xRlgLx4mZmONuzqRuAllcn78ItS7docRWklH
yk7wqzEI81wSslj4/Owz6ksli6Zl7K21bIWV3LC046UbHwUL+3zt6CWF2i37
F+tS9kC7hSmpEaTiD8l02qNLwF6m8iKHkgiONqDi22hVOYkllJ9RDdcvpozj
kmjr79wW4t/w7Pz9Q1y2aqd2IzQM+pQ6LPbHw8SPKI9I0wsUpr77gidXitQj
q6XTgbKK7aCU6JJ7gIzGkR0mXjRddWzmjBxA4w67VXotJTYJd+egBy7Z0D/w
Tk7nUdvNSj+bOF5o9jbHx0P8zhy/Ih6PgoB6EEaNyaCQy7lf1KsiwUeW3C0n
Jsim2k7GxFvQW0T/6/hP0jMoIKuweZxNdTbRLPKqB94h71lyMnUHCQGMCne5
9rvyYDH3Hmrzf3I/T0+uwrNPxvqzMSpXXk4RxOQ5ibzPhLBB2Uma1qhH58bu
lGZaviQwUL0zPDiYcElApTG0RlaOf41NKDrPvM3B7Qhstq+y7fibm7b9Z1eF
TI5yDmlTjVSN8Y315IW6t/yLlv/o6VEAPHoLXrCAeQANdpBJy+7scZca8g9L
CKMzUThwgM/KWLTMHvLcFall9EENuqn4TXBlMvnkNCaYP5YZq3k7+0PUwVJH
d5LrQD7yHso+3XicTVOYn8epA5yX6A3sgnLTicVR0yTeU61HQww0dzBDQiA3
TlIHh8HO1lafXSlKVfF8XlhluotxlMn6XjStO5U/+J5zKyb/4RhokveKnG2E
DLjOtM2FWc/OLWk56ZeK+IjfcSexnP6XiQ0U+r2hewDmqutrIIRHWoc8hxK9
gJSlh/Mij8CfddKBuLR24wlrGcGBUm3l2HT8hEKVFDFEn3uZHxgSG0BBPxXr
2yP2/eJbpycXsssBaQyaN+7ljh8gipsde/tjJAkAZvjp7nYzjBg1dmP3sn8c
vRRn8tJ7FAxTIXqQWKx0RfQckg81UPBbpGX8cAWb/z7zhunPozSmWgk+3S+d
xQcwITTY6Z13zXz6B7sNhRjUSPJ7ig4S+y1nPPQGFakXJ1rzXl5v+0pjbycu
4bEPe9/3lXzdTRtkJbH+Am/VYlv98R7htrzwbu1JzQpbQFzT+UzkkDXJcXVb
DqhFCPks6jUXU2/GkKoDI6sS3rkNC+OQ4ux3L3L+HwUGIzl+HbEkKZ4vHGx9
+lY96sGwGm+XjST8aYvQ7tio71wY7dLmhwL533+iJHMAMCuphmcW3XMj7iWT
HnDgbnszf1fjRNhkb7O8jEqFer5VR6x7sts5BQ5DZ5iqmE8A6qkbOjXcuFGH
lI2ucBK4lnTdU+B3HeI+etipOEY2bThdKqXodz3xZDP9wN630CNMrAyw79y+
417ZJ7n08CoA781T1otdjG+M7rKo45laBc1oeExofpl5fp7S0wFKepYslb8V
8hVVB6V6Ao1y0eZl7b8oHhuicJhbQouFumLjXM48iVEFFD3v9bzGojnuuqth
E3BPNJp1Xp1UBQhXzBM83awYumrEv0dgH26MVKPq6asgFhxMlX6T4a74sgFo
js+dEtJTS0DguaJq3BIuuCX9dCtuppTyCMDb6muy1vdrRyuYFWyaoewePWcd
5cFejW6Q9uq4HhiG+uOrfzCw2K+iRih8QEWUM7jYkwhMpvyoFSmqYQ72Mua6
fJsrmrBHxYWxHlmfWO8AHnZ2eUFI4Z7QG0L1VeMZyDNcW7MRYM7S4mYeSPnb
hG9fQP7wdoeNwr13mct5KDhgw6TpIeU4M9g3MTTOXAtXUBSL6bnrLH0hx2x0
3aaRuYTc9XsSQkIZZtliQqqxUrNvVP2enDR2Q4MnPnozpGSMRq5qLnKzMo6h
wg/T8nJcSi6eO6Wd2eUKPXPzKLbTobme88pBQGPsahwaGZ3YssM0fFsDdH+0
WrwnSBiWpksSmjMGBW95hTrsSJDe6h6+DZh6sBGfUevA2CTJ3itl24hFL2MV
dZPxrKCjMhcn0dmjcTrgGMkVa7xvFf/Q0sMmRRPloupRHNKeiivCbpKGNXXq
8Pp8+erXUhKxJiIAvw6JJtA6jlnmY7vOZoQVWzTpfC2nyAGDfp88cAfKbJ+0
kXPO474Vv/JnKq81dC0MwQqm1QIzHf12TeCOQUNFc1ivnMBcBrGTWh331ubA
FMckpSFiuAMAZx6fdhjjGdv82Gd5nnBzVqak/23vJTVbI611N95P7lDusaeL
0P7BkhtMr46RjvFhoPlwlm0Bf/HCJxrd5PiuPqQd8copXeTkeZwtCf6choz0
Ac4DdwJ7At7O+1ph+3+vCq/BwHx6nAc74VRHflszCdP2Po9N+NGf6UySPQWT
Jcl1VI6JeBD7w/UF6/m8AKEt+mpz8WAI+3jHzLITwRxNwR07H83qwSki2s0W
2COghTFLsucfUiPvii1nY26Nk4hPrmC0gIfyoxRlPAh22qgAuFdZgA0SBqsM
HjxpovC5rlQDl97UTO+h3njHfAEnKrYybELE1k4c6gSYudEviciw4FPyP1xF
MM6Y512fMgc6PrUwxZNnEMdwJePNj0+CTk/D7mn7mln1NODYzbtZUBp201Tg
15dgJnp3AEuHGCm99beGKZHqoxcwtu8+xdA9OBDPyeaVh03MH1Og0yTGPRcb
nFQGJAf4psQTvt+jUgpoHc5mwUMET6d55Bng7IOC19YUisx0z0VNFX9Vzdzf
iXlyoWNEKkOUxoGyCQuOMwrlW4EcRBQmz3M50ZSBe4utNoOS3dVxV83uy/YU
+oJ0N2ooXMHRmHiDIZpSLOc9jtuu/bMs3vnPU8umyduOcBF4q3Ub/jfnm33A
VaZYL5vBkTXfMWo+FuL0ayg+OCn0/0lhbhR6cj0l7iPdfDqOkOsizLb84Vu9
Tbb6aTPRkwu4+FFsTyjZIN5u/U6+TY9JwRZqZGXUKZzQX9em9RBPK4wrVdbD
HkL6hUvzL71c4KI+3irw9osLrYpMQ0BpWfKaF46twfvHrgYLxfr994OPVdKH
/qDAyH86CU3hcSrmMNstlfFnONfFQSFgpDqyIqJRKNISI+dvVq7k95KikCSu
wd0Zd4UoQKnc0QaNiv212o4Q3YJeMmWWiq64OFhf8SktvltrA0Ooro/fsTs/
Xo4uHiTE5/cHeH6ty+LWm6qNAzZ8lewt+ReEbJS8MsxKOy9gu+7XjcWYzyI8
qht3uA0jdQa+L/eJdOlVsIeex5r1W0SLUGx0bQM+/dE+obGeqx01vVXezL8Q
wCf/BIHzqyYyO3bpqp/qAOUn5+RBW0d2Tv0Feh7SNtXgkk8cLwHr4OILVuey
l4/kpyuLioMMJxA9+7bnKoRyAHQ0Rd0CyGK4iRu/GAHsaqoqXXpQ28u0fYDn
ITmBLQFFnl+wNGKc0TAed9oGeXgq2LKZR3IR/WHKTw7er0Swb0+9Lot7Q8hp
+JYKzh1s98PhBKor3BUpol7Y+QV6dfTsJfxClcNgn6WscwVxGHnSf6MPBMAe
6WNcjvcsfXYoB/P4cmqajENqtCvU4ZvftuIaCBlUIQ5Ox6nj2wnHaBqrX+rn
bKOoja/9iBVEaH7i8Db/HpeG20HWKBL6hvdsXMydjcWZ7BfvyHlrdJXM6Hj6
xw5lgWGjfJjLnhLLhCLIseEbi84VG9D3BVtYh7MIJhOX6CU6gLgu+SQ/q4L5
jdgXJTbK84T3AgF7TNS2iGvtARU/+gLRW6AqvY1ACZ2wOmCx8hgoKNPcMnBv
ltth6LGK7pd1nhIqShK2IFJ4bHcYsNYk4BaNZZJ0ZPMifflFR2GjLYPdhbwQ
wpunobuRw7kflr03Rn6gDGTYsyZ5QMWL5MHNZg/pQ0hry0d966r70t91glOx
kAEbBOAHlcrYRonyUGwhb13QPS7DDCgnosaC9Rn6IINCWRqb1UvgAOX8J+us
wTIi+kKFY3F6B3gR0lhGFl6bpw9TCs+io/jg33UDm+yGreIXPj5dbCGcK28W
OOaHCLEqw438LW98gNzQsaeOTdmnmaJqaaRqjY3f2/N6Yqcq78pvZ7JkQ2Rd
GoAQuH094lN6tiD/DxmkmC0UlgsRZiVa2JvMrGrZYvZBPG6U5y16SefOztWm
WlEtlRzkFL8OcsxaE9kXFNE1KldKUHBG0j/1R/drR8gpez7g6GAzODzMxNpa
MPO9xe2M45484snS+9k5u2gI77695hEmfEtrjJu6hhxzyQW3jIzWbiHpysf3
f7iPgwcYlVvObhngupGENgS3mu1fZuva5zkSv7h+addZ8GktkmZn8a9kGIhS
CYqqw5VhRe2So8hLJAQf3x6+XHpuWheMkJLNAzIEn+NvwVOk65tEq3gobVas
HG+6wwcz8a9+ELSMR6ti/d2DqdMqS/fWWtREWRycjY2viw5TJlQCmGDBZNnl
5/EQT8sn7CkEFoDsgljZQegFdFww4tSaHY8KMTLZtFHPDU2t2QG6EmAZLsiI
9e1PQInxq+Mu+KbqFc5pQmLX+7h4G5BT3oF9lKO8tBOtLIESYxL3MMp2Dwbf
7LIWAX7hSD436Fsv2fmY71UOPkRCRO0XeoAhE0Xkotm0jV3vhpUA3QRFi+4W
6/eB9whjnWMvtK6XbpHufu5otdC43nt/dv+bQ3MkeQdu0pyrIiZXNxCJbOSg
TlDCi6SyqubeectG2Sb1vzkr6lbhus5rYXDT3XGs9WDGUKuv1HDKYzzF1nH8
dFX2sRVqUjwJ+4XWXbBwB2jUD6CE1WKAJuOXp3Ciq6zalBROC5E7ndum7Sa5
90xelCA3iCygoI5WK7Lebw19vagqE91LeIBnTRePJ/ZerZDREob2jLMgnIDn
EXaMtvaGK8TxCmz/Cxg26VbzSg6WhHdxHX2tEJ9J5ENNoi9345CRwUPL5+js
t0fViKjH0gSGKfNmnmHz7s31fhzrOqH6Ypz/OxGFZ8WfQ4fPIlZLPXZUHZky
av06vB8XYKFZcIvQGwC15/b9fQkCm3n5yWUlWM5f2CUJquGU+cIalRK9Cc6H
SUIhXQN8X0oHFz8Ra03wBw2vby2ipNOUF7ueC+IZOBldYMlTJzizib1MHRr4
JiUceEx322iU6vwXnfiVvXaFpmi/ivmhPzXG6DwKef/3LnAIDKQ50m/+FNaB
/W0KgPUoV0gAB1xGW2Q1Q0qlsictKgy9xPRb3zRIvHzafq5Knt7O/2uSJOVb
ShKq7nB2Vm37iZrL96DZVkyit3ft0iX77OKyJLmMFUYAnjhyxObE/4bl4jNM
l0Fsh2ba4o7c//0ycmKj53TeaQmCez2eGwuhNygNq51353N6QP8JqfHksRU3
Bo4PtM3cWJJACy5wwRzljMCPdnvWfHOr0N3abBZOOrAWIoeDD4TWSe36e77p
NBwM+m0a/7jOucpo+80+IrR2zzX25d6gWCTEuyqpKsENEY9gbLWVVS6QCcPX
RrtDgHBUxMlxc4OaddVek1rr4mYgrkTMCgtmhnv5Bpnu5u2gDiEXVuRJzB3G
xSm3my/PdzNXRxj/mN2i5fD+PWOwoWLclllqxCu8iKV+R6GCXxVxsamhI5Tl
iCuEqOqikFPo/eNq4Xb8bQskCjMxqqQuZTK0eDOnrbQx1WQCAT0efNtlCsvE
qfc4ouFqEA8t6TDZPLshd6qydOQE5TNnn7m+WwV+pWGCR/wYlxxkLK355oiH
oLWx4vyver/lEIdRyUZTbciPhxpX9f1e6myg2Muo1dH1enGe4Jvx+uVxIujh
GPqzyT3WISpEuydmzptuOw1Ga3NehLMFCuKANTt+Ea3JG8A8e+PCIczGhX3s
/ZXkKeXDK/Jg9cKwN9cNaFx0IuPMBYQfDKvJWs51XwMF2l2+Je/d9HomPexo
gytxZjmy9UB5FzvGnY1IWV9ST0ALtGl3f1OTAoYTe8wn2u16CQY/JpcqXECk
eh2nju2jU6sxYIkOBW+GJKcHhvfe/36rMMKPNngYJ4XxMaDMoPyQ1PSsnBxm
fp7PzgGBcGHGxe7TsDeh0qz4XoAqcRGHOwgMU7DzLB2JIshE7YtLivpSm+2g
+fqkmpIYX6m6MHWUJHqo6vOfEUILw0cVQJjSy2pnPTa2Ke0h2nOnilUgQA0m
rQ0Wvb8CrgyFvS32cbZo7LNDciu6U39sBzKh39rv+12S2HrmLI5FH0b6Zm9z
sqE/PKxHc8DxPpqF3uEhK3dU0Nxj4PtGj18nSCopnmjs7s09gvieLsMqTd9m
4HxQnwqvBXwIAadSHXGBMSKL5ceJmoKKVXahVV1SkM1jf0q2O97Bw61aCDp3
f8EePA1X0gXnKK9AmcaLICa4X8DFWh6BVwM5mGE9e3+5HyavkknKnlBgchRD
sVdlpVO3k7zfuVWKxlqRWgEFxQty+REiWdX2nHYiiEouXaTxWCwOMUXUxp1L
uxRSy+9IwBBC0oqvFG+W1SzBn4VaJUh0wlB0FpZ5RIaMZRJvPcUBtRuqWFhh
uK36UYtpb7XYJBqVlZQ0gyOTuUeIL/882Dn/FWonofQETsQ98w7FJu8UkGYJ
68cNobFxPSKZDP4znW11UzCvPY1QSJ9DsHPybKryZ/RbzmH2RNYhQ0pPu+cb
l1NsYH4kP14h1r5DrojeI/EOsOKFIVhtxgM89G/3bApWF6iimbkB3moZwrNz
WZM65Hm+6IHf+bGMOxbYONNRBuO8vwAHxy1G7fMyF4lFKaGPG32G0jSf1jSs
MBG163FWPpwYKed4c0prgaedPzP7uHXzm3VODvdIXCKw1KqLdmpWFtdzVt8N
BeE41jvvotnehQ2e0ixVUEeJ5Pf2JyJphEtHaSTu+TgFxUwkbVxqjeF5Teny
LQZ+CwS3jyQUkMcqTT0m8KdHqWR51Ui/77YoP0xBjT651zvFsJNY8FvVSExD
u9SGBxV6Jvfw4aq4wL+TDkbvJkG/PZeG+xL/zdaTwHhJVB3AFq+R5jmlJaes
zlcxNTsYWihfKIvL2BNUP7RBhYIwdNRWanvVjHp8lEsEs53Llr0cFikKSUZO
O4SBTX2DqQ2/O10EmYE8hKz9ctILUggz78NVfjJgmOBaUUpymAw7niLlhKJq
hRhASJW+4dbr0fY4rShRe2v843gucu+bK83xOox9XXKdGjyv/VoOZRAX3D/b
Ie68r7KIuxtL/piw3moe9khy/NM9j1zLfXWfx1TjYqKz5aCdN/EviU/bt+wz
+arChYQdQeRl4/lCKCjn9U5d+04UDnDDUPjSgCaj/Te8IE6gVapBH2WSdEBb
SjNY1A+aLxvxMHsdQ8tqFygDOO/Z0B4b0wh3KloGhfcGudN5iU74bH5+0tn9
acewxJyRNI6pXOOZqOXSrmN5N2R4DN9avzTAdTnGo83xFt91JVs/n0y4cYQQ
UyXZM/CVkDOac+u6v6NSQVCPPMpor/etRsyRbiLQfMeEPvBkQQxlaqu61ppS
PUyUjtbdQOx+5dj+LSpSytZL3CE/1+mKy+EK3DnCz/J7c9l7NEw+aSCImLeC
HuPqPKRqZayoN/1T9YHfC6RQ+BxLjcMr4mHm6BjyAxcb3I3eN4YgfSoE5wvO
YcZst74XTvF/dDjGRv05RMJws2jof0lXqqaGOZtWVDMnbI0/NDNXn0naVfqk
sRpsepmz5CHqM81oEhbnPAm4Ztt+FF7wwUu7kkLEvs27V4RaYkJ4uIUHVwUf
VKgks30K5niWRZNi+h48hvoNGtcF4pPUaYzLDm5aYJ1/AAUREC24MJihoqRI
AWTdAmTOrLVHip5MCwtXBNnmRJI4KFVH0LHYvwT272ufVibYbsp6RXqMSHo7
VSfjYfgWsCpuG/dGRWK+1zY3ay08YVNw1kdtAIUDp3p8LjcoaBhOA/mjUgpg
OiraL4YoK85E2AfmJM7jBrT8G62tAOD/hF6pUTaMMikjyTlYdbpbMFANH4VG
9btv6UL8PM3wJRRdAoal9FFCY9TUUUszn43rWXGmLwt5kd9vxNg//gb0AMRI
yjIUeX+iV4qRqNJDq7bu9CORlmDII6ETJI9ypPKbyVn1D+PcuVpxWXlYAZ/Q
72lGAD6tJTcp7sQPXNpRLNvhEo6PR5pBMKk5oBl8hcCojGePXTqiGTWPZfOn
X5QtyMejO/L7x+/IjhFeSZPnl3Ex5TWH25XaT3JnsY08elBA03JxkdS75noR
vXzvpnfYvThGH1XD8KWHJLX+9eK+M2buejmk2BUelaJ9nsXM/+Y39cgDYNwn
6xiWBnfrxENkifJaQRBQsM5zR8KL1vfuuAlPAhk/xDL1+SKp/4Min4VEpmD8
6jrp7E8MtSF3rsqLVPAHIrTEgEX2II/13uLkXNGFNE+Uv26uUprgVzYnWx49
qU37EcDMk6/x8Us4EsPYbHyLBjUOqYK+zTPk9eUD9d06uGHpRHK82LW2YZCa
UPZvFot2OY7/pNSy1GMabYQUi9ZigIlOdnZAuWqAVy6MUf3Lxd2yQgbTSn3J
3Bj6yBm7CyX6yiKLVwU2HSWdL8QeXZjK/RSqyfsR0YpPSSbxvCjkvYUp4Mow
L4ZHjFu/YTcbyorIvXrxuhUzGLp/pgwkXGBFzMVMXzHJRE/E0HZlCnSCV0qM
TaWa/LbXKADtVXJALslnOx9WLJc8t+OXzv9j2oT8/f1jE6c1sodTa3bsYUC4
aqKGp6UdysUb/fB0Cfp9f5WZ8tyyPoB1PzKlk/MZzh2UAtGh09eUXNJpQyVU
GSc+96XU1thTT+NTewJee8f2iSZcr1lv7bO+uycJ0YRZaXOvqoNJelAHnvLp
iw/HmxG33e6Eq+aBNAij9TXTiSbuzvAqmx98A0Aafh5kvnCmLyUN6muOcr1i
QlhgLwKHA/nxpm3iwbd6y9UhROq7Lu8I0CrL28yNtP2EVgPipJPeQxn2FExK
gh8RKeXPwSg2D5Sk9QgFbuQjM2qEO6Hb5jIavNSbjkis/FGuOt7FuMCKEyyQ
6W7fzWL3CZQ3s8jLqEc6q6ATP4B37snZz91gYpJnL806+JzcJ31xk8YyYqH5
AefPi573v1tU/WihVych8JyalHAvG87CqzWDtB0AyxFoSSCNq47HyYGZRkwv
2LigBW0Uvo1oPW4PARM2y1OKIevZWAH6h2zMnmO2qWdsjvvDRBPFBsgQEr7E
AKDOBaCvQh5tNQDCqxbMbfnkjvFZfiaugQbkRxLJEZjajPWUiGTgbuR1XMXN
MDOQ0uVZhY6fCLwPOrwBj6DxeEFx7UKRRoD+UT4Mx279mvrQtLveKRBsfjxD
cVqZRzndU1XWf0p9gpgpZd0/nQNu5RYBlAT+Ak5+U9R9jKWUKALsypmuvlra
U1CUIOdhzNAz6ZUiyGH2CZKCb5zGmy1jF7/FSl7opo6p+HnCqLVabC/LdWHr
dKqSRT0K0+EhK78Y2kmdYxF3EvoP+Wzbndkxy8nt6uJWtYHtScaDm9HoTiOz
epUafwMu9dKaJ2JpHTqAZ0a9cu7F3o2Dueq0qZziA5qmCwnMi5n7a7BBDcBN
51RxQDC9hRlpeDuSIwIMIn4qBZ1EjsLprnIcfPqLQWM6sflG4k3Ym9Cj28h+
tEaZMHYJN6CCiv/wT8ss0lyYX4416UDLHTsZc1lKcpXaacBBpkDoH8/uNwAq
99iMK4uGzbcvQp/61qqOocBSvwQHUJYaqaNecUGEswwhOebj63dHPV9NCLBz
6xkPlpmlMcn8e+8uzB9I2PNirimW+JpzAs2lxBjftAQA+637zV5AXwOhXD9x
89uPe3nfncb6/oVKm06gZk76uvAcdtKO//4DMYy1C8Z51W0NuUW9cIYekCbX
bDurSmhWfVKKyaYnL6BoBwl3ySMpA7h4Th04pLCs3jDQ6FFKrZlidbxnaI+c
RC1bBx76RaF+9jII+OX5r3I7OOvlLN3cuiH2pd9Eg7fxgIyBmyiW88VzYoxG
x2QDrr6h3zBFKatp6TXr2hIZ+wh2DYy3JqqAL7i8vMVQh4ef4jKHm2tbZtBc
yrMwVKyfjEqvG33tqm6+AmYNmufbD8YNvphLPvAjoRSSsNRaYs0v9P3VWfWQ
AI7RF07Il8Jr3ujpqDS/ckrM+lpBmRqkx36MbM3t+GMECivxbb+8TMhvBu9+
aC8GiiZy8z/walZOxNbZ/2qNUKzKnkTo8uWYR5hjVr29g/3Z8pv8YeTzJIbo
NTJYbMgBLPvxIU2RMc421SC0Q/oi31818neYKU0e6ypqppZhQiUHjH/RL101
ktmjazyoUfc28eDEMY51AKBtwO8/WMIsAuqTnpXdUxKLzXgblXuzp4N+h++5
VpUrCE6krp/qj1TmKizXlbguEyMPkBnM/XY8sYhjuWJs5EgTOSJj2RSK8lX1
lm0HuUqlvM9J9ukCMRKebwNeooOp1nJ+yoM54+cT9F0L/oHPiKXLvDeH13Li
9jjlZhRP4gocN00jZ9+ZuOM+9xcy1aGh5sfX7CX9q7GG9KNvh1EtCCCb9E6v
fjM+va5l0wv/QLZ0lZk6GaVBWtW6hvxPhzxoP27dNXD0619li3bEcR81vp8a
V3xPtV1SKt5K/JTwtbWALjvFKj77sRnbm/V8ES5S51qWZPs7L0N2J+uy2smj
vBGwntOW9Y7cHR0q5FsmkHD/O1/iCYIE2f7DDZJsoOtZwfQmCSfKPO3xJNuI
9ix18vs9GiyFuI/fUlb0iqKHxg1/wL+RMkJ1j6WXpvY4kEbXDdFAI2qyFJjU
lVS35gfOOr6babRWD8qd+j8l3KpCs7xsWeZghGqiuv1vuKbB6xgOsBatj8Tq
PYjVL7dBlIkM+JZEYWpaP9hDOpetLY40lbId+ZGrU4K3Vg39tHYmhjenRMsk
qjC5vjUDTZD0xdO5VQS7jsXYJba1XNyXGrhkTx5Zg7DQB6XEpktAZP/rzDrE
CEvXDiB7aiI/GYpvXhoQGPbiabbFuvWWTPBZHTLkjgVk8VrWtVDYZnoVP15T
RB/0zEGJnWSo8bcU2B2Wb11yHvAmh3ewgSMrHevQsFNxNyWCGwN7QMRytfLR
nImKBFU9BBr2UI8UhO4y/S/bTVS0+biygtkYSzhJYQO1bGzSLjktQgpPp8eq
WKMamPqD5n72FrtBzfIkoJS97gL/fX0I2GNGib+ZOK3Hcojjvzd7Fadl+IRt
cwgYdFCVxnRtFroIiE9A9PQZ8jLk4RmGgM7g2bKJbwfyJOlSfPbyPA7MbUh1
Q+nYqbX6BDlI3odIuLsPoOAKQL/LKLkqc7jMuS7hywyKwBzPTxzcp7bYak7J
ah+yCNVzxYjNPohhg4HHiMc6i4XRJN6iedsSMdprh1uuobnhysQk7mR/3HOF
TGXzoTw5CcqUYN/sOdy+iomXYotOZp8bMG8sAM2l0h+IX4o0lAFPkE8b7HfH
yYQoFqWUB1AZ3jleLm3xvacrArOtUiedGPIoqdrZ1u1K5z2wNAZaER9SHjVk
9TqV72rXfC3Y5c4sbK0/iAVZfyRuyOtcQfQeJMUbg+sLzwOMH0zSEBSACAHW
KqsQk6OU9YDHEOqxc5egnhIFO4nbc+NpORpqB+MDYEDGY7syJfVMN+/a309x
RYU7l0iQaRdDsOOIcTt60ZILCzPN2uQxMt0/5qvhAGdbIwXNMFi14Z4lo9mq
Ld9BDg4rDSC3U7vjxag03RsVzlk4/HRSKes1uLk8DxJzQniT9s3YzWR6yL3v
s3C2+1N8KrzmAvtAQtUadBx9F9ZhmomwdzDv6KxiCiRYBHd84A4krm+4Kt5a
Pnmy2pNG8gmYSu+rMd9Yh+3En3SFaCZKgYqqxO302c0XRuYKK8mm0H9plSVh
rIopiow3Tf0Mw8GvTBT9jxewBkzD/9w8cl3F5omL3YervtgfjtCpR7QUYsRm
c9F0BivOwqFEgWUAa00vJ9RL3V7otouDRU56LuGGKmysy1ivvUGBs9/gl3CH
ZXoQc3ZRoVnXX1fs+3tKuSazp5px6r1O0C2S0LNxCCCsS9GuyieT/dGTWBea
41PIlTGGCv5/17Yoin/H3UHXTKNfevOgucreY71Ik2nLxAMBjlVctcRBAZwq
NVYSB3jeZds6MXgH5l3OXVd6lSI3BgKKw+biETZfNh00fFpteDyD36sIsVAj
x8rBzB+xScp1xLAVpaNw8NtVxooAZXCTfUY6olU2H86rpCBojHM6ScEWH3GV
FPOb1ab4fS2JO+2qn8juYIaNbSiU42cMwCd4GPa82JYYOvLbOE6ulqlepu8Z
qYgitW1+GkAcaDtKd/VG8wSCKdyS2hH49sXSrWzpgIOZM0GdZ1z5s6bLckV0
MffWAWg7IvJKLdeWPfi4yIdlBG9Z2ezrxcHlpGMGrb6hiYF6zF03HqNyzrOC
BP+epU+y/RiKnqK4pP0SventSUbc4anyAVxwqnCM77Og1iJkCfgzgyUeeKKh
/d3v45bl5bA/D9+znjNb5M+lcUUfcH6pwXTBJChieCyDTS/vYuU7y7ntIUAf
W27NsV1H5kCespiBodJgVZvRXznmlA7clAkrkN/TYPkBV2/307UrGtxXO160
BtlyvL2uMZtDUpDL7bdRSuB30HsSc6zbnDt2tuG2M0yHdOpsDEo9wUhsWf+r
CJWokc9P2V5IILfsRjM2yktMVgZdGUSwxxPI8hftTWWR+4FIcM2sxJakY34g
pjAyukpdUS47J+vkDq+Vq+bK3U5ZqpBI2kjvwLY9w4F7us1ICIJvJ0MVLDFd
42WVYXX8x/SQYkXE763k/tToXk5LcTtgJjkX4DL8p5vRBQYw4MzUNgsEJ3jH
g5yqjGKx3g8jz/R477KYNTnArY1ml4giadNN0rBcXOHz/hYgtn7Vj5gk5xsK
kcv+K2awIiKEtSTERVeDYhRuD3HATWsDOgTOKh+ovSc8aVgN1U1DIcQGTLvv
6DOmJatHYDI6vQKq4Mji7NuCM/uI7SDO0gbfJXQv0fbUN//6Nord6nmEEFre
qwoXKTgeDe3hgq4vuPs/curWr9Yv2yKeaB9PNdd59i/cIUvAUIxn+vPPKPQs
ZqppPdbHNB20+J87kM4KAcq4VfNuAjQE+nMastnKre8dtwrnN3y/hQlW9IgJ
Ln7XRq978cZCi9BUTvGbKJVH+bJJiF89XoMC7V9+qVLEdJB9efAA6V2FGvCQ
j4pDq9DP2X+Ox8Qp0oERPfGiuQIdeydGQoldQulfASdgOeA8KmRx9MbK3CYy
uAzyDDxYqCRflt17f4JlrANTtelBmCltHTatDibE3yCh+A9Ve5E6/FlP82zx
vQudWFabj6d8ltMkqYREcuzzF5KmKBwT+G4+rNm5nclcXVqR0ygDk+oNTuDN
BBaOTTRIRrAsfx6KzdsvskYF44btA87OK1pcV4u2Jgk7NQQhyv3NbkvrvEqA
2nhF1v0XrEG6AmDSCyVo/0xs3ZxzZK0x5Wr+amBJ4VciwPNlms1hv1SElTuQ
rk4qMETAmsY4Ju+V8IehLq30dqLoEYTGbCNESQCxJyndR42mftr9wdoBpMZS
pn5wk2ByOwbkVbFl9kHRpN3j/SG3kYoBU0ftG+2Kt8ddh4SNOQAQ5MgEN+wL
PpccpIX1aJTWqaGhtZN+6HgH+fShCktPp8CrlYIP+F0dSaUwKduy+QJrYcFA
KLTyw/NJO+VP900qHLuheyN2f3EBs19inK1xjQobX5pyABVuPBsxGU4lYH3m
uY2I+Dv6zSzfHi5J/5cNnYavAFb/2XEE7Ml/pTJcn8ABJeJzW880/XV0DT4D
uOMYoQUhVr/78sUDKgbD6L9jweGIai8voTY58/2ccJSxA/sLmaiWO8G5Q+d3
re7i2Jb5Y/yLbNe1tpnJbXHbVdi5w3nrCxoo9FYWdFPUdIAun3dXwiOH5X0W
rYAeskgOltYTv76J0+4rJGgYpV9Glbs58+4Z1CWmuDGxNWGoVFseF5QSzdtw
HFuXu+knqHfq6r9448wNpig/WJxxU+bcaTpsuxoDHNgQogFeLEQK7qJt2C8T
Koqj54opS5DQimUOocL3WxKMfKBnp7sij6jtDWpjbV7Dwg0PDzH1AdtVo/jD
g1BIM1MivBTtC3hERGqs8Ox8e43+hpwsHRGLgRtNSAbmNTsfY2bDua6TLQDH
m2M6+6hbN1TFBkj2i3VRFzHEumjJ7CcjMIclfq1iZnVmcjG1e2XPW0g9C7Af
+fqpxMGZA8YOciUdM8zne2pBmJrsLScQDlJwZEgxBfSkdFFgLAK1UTY4W7j/
jrOenSRNdWnx4VeCQX7yWICpBX9p018GhCPzhBjULQyDTorOcr2G0iWQ/OEj
6stpZ9m4KCQRKeBSR1BMrwpBLJ3Im7MCBXthQgAVMCd7ay9oR2Ohvet2EaQz
+s+VQWQpjERB7k/ZnIBjnkm3yI2swI0PuQm395GtMUX0SGjS3ZIC7dTJmy1E
GyoOUpnb1W/y6EQuBP/TBYB0mMV+He/q1I/Mp5tmr+zkJaVAPM4gU92v+aO0
TL16z6atbXEptJcpqaFPbDnSmWjaZ+HDTsASJdujezs+yYH/NHNgYn1ndYph
dvgyAEOoOzSmfDp+zg02/InC5p4yb7SmmCcDjQspywGtyKWn7dXY3D8n0Qgm
gg8WCLG+7tl7EECfjD4K/GnvmT21VXo5FJLSiiEtbEEkfoCtd9YF5sEf/ztB
kgcsF1wRBawVxRFHXhBASZAMutcLH3jxZ5c3Mei99lPeUJUb92XHjn1ZeJB/
PGWbMx5WV/ELFI8CkmjMFGF4N4A/K7UYjKHvPE0sXakyEStCJEB5bb5jrKw5
e3WQbRzi9Fg6zIJhT5o1ndbESL81Pv8q67HXWrxXgRQwx/izQJ8qmlTFEX+L
3A2FdB6FdVv5/1CmXGC5zmgNS8z3I0daa6jrYmnc3NpwA9m7jpo7TAPLS898
xE3m1vSe9603exiNngtyzW2xPvRIEN04Ld9P7c2K8FeQhDZYeia8glFFFN15
6P0/RhxF6XfI1ThSyAHs2zg8rY7Y0AJmRRDhZDnmeDm8XyWrssAn+o4FA+hP
bag7g/D+68K6cJ9gzxgBUFrqQn40HsRiW/flEofGFUkJgMNIy+LTcDgdLurT
zEb/ohz0fNe9BWlCIpt2HJRCr6DN5YMSaN923wu+Cy+yIaKo9NuwpnGNknyn
l9XUi61KP64O5Q36R2lqkTie483ONd1xVQBbocXN0VYlk1bE1ZzqGr9i/oT1
QlM5yAnPdTeDOy9oYzEbyAObZ6+6+XouO2fcjDGt0l6RDEQ+rChVmGBaTSqQ
FRTUSMk+8XTWtKyimGVfBziZGVaWWqOK9gOJYQpm681VeuhWUQsiMnAWxjlj
wdhK47ew+6uWFfffKixznTYIU8sJDoWZ1oUZNSQifm14BouNCahBXYlTh7vC
oN1l5hDvXSKDaXt3qT2NYhfLMZv8cQLP/No9SfDzPyg4wQn7rbmunworHwBl
rQ3JpjvnbAZbDNhrcP68GEvw03Rs/U/d/dlhHe/ywOtE05oJ5ezuB0b4c4g8
tTp90uWhMezlwy8xBZtnC7VNX0VBTDud32BBp+UJZ5pwslj1s9kD4dp4ktOd
DUGMlhGX4x46PmUUC+h5052JWSrRxwoFep+ks84uYLicdCVY+2jhtB955gbl
J7f19qhVNpUS8blRITiC5Y9sd9R0r+CMD2FccDD3aWZ2OU8rFtIbCzBllC1g
lVYTZm6CTNbcjkB3jgaVc960tB03Qlkqeid4/iHyFq9Jc9njeSVEwTl+ZB/1
mZBBjznSyFqFcobF8bTzlNBfrAkquB3jGpTib571vh10piXYOadNLCHV9wnf
C5a5EJpEefB0Oa5wkRJaLg7QR4dZrXxuOfdwKF8i1DYeIg5kQ6ZiocvfTWRJ
8YlR8Ejw3sNA8MOPAsVV7K6syfNgMANymht/jaifAZdqO28EzKjSy6x9aBIb
erW37a2FgdPjuw237zWWWhz8oyfTlfObLa8G3OI3oQe+N9WJj8f6zyUh1KAM
HgMzvvZKA/NLXF1TcQdNFQhu3YPC0ZdnJoL+0YGPuiBWCKtim7Oj6pLeDmLd
SJpa27fVB8PT1d6Rrk0T/Fj+ca8ifd0m18zXi3HLtsVruezpMEIZ6xGmxD4G
GxGpoA07xjiP+kBG4nBF5Gn3zZRnTieAUfjjA5Vdv4w6LKw1w0NYvUtQ50OM
HRo5Ad3hCcYsmApkax2DdZKQcwaqB91028MarXosMPhDQm6TqH8qXJ0DhI0/
7aRRSQa0SAfO+QmUPc4denYDxcP/cC8tN/odgXcDc70ZU6ZXdQO/F6nhJ4ym
PH3BIgxs22NFYEa1tWrROtusGTb2JusEYpgPj1Z7rDD4zNic4FFkv8i7PXHM
8t5INJI/zP7IuKibxg+uGFWUI51H404xAyk+WPqNznkz8aPvBGuwMVAsGgnX
I1RMpZJKit3Cw7vAl8Jpuw49Ybct8WVvEISo8F6wOK1yg4JW4+V+Whmy8iin
3oFdW6WQCD+yh/qQWZiAWiAY6sXPiMBwinHkEb3TafulZSq7B4Lm0xpFrNxl
Lu2iFW9CFnDyPiskmQRcmmxw4Klqp2rqPUc524RDHcbNuLeM1dN1UKntdjmg
we2jRzLQeL/otAPoeYJvBbE+YN+KkGAwWzF/stlmOGgVJPEIPYpLZxb4kAOY
BkOk37kQok6HJRwPVtKmAavn4PIcmzTkq+cAOZ1HDztgc8hWZqzDHAF91c5u
+y87Ww0kQYIvgQjSMqEmzai80abRL6yusjd0nQLjeDgbYBXWgrikhnAVxKCy
//jpL3HqwmrrwB8RsTlTlUomUz3hGCF79Y95UuILj6KocrRqhtOwmlKojsbF
UkqWSgG0w41rzIDg0XaLMlVd0M6NQwTauL3VYlrJwWoIWSfshi5uPnZU0b+O
23dl1hn0VS3CYSKrOuU/IoSKc3laX+qN2spTSA416p09tbFAP1F1l3x2eSnb
9yhPZxV7/iRUQvSTo3P1vNZmtr1Mdwritomjri+7iI+0bVB2Yv5Qaan0S9Pd
p33xLHE6hhNEPOcpwgqr9vHUH+4XEIReQ2nxeQPkFaIg9GaQsw5Fx1ZhKNa9
Ip9qPoy66yg36csFoLbJJa/mjVIkfsrIf151tvs1M9W+assDRBQuiqmmjTrP
En6dbQwjZIFFvSYz4mKqd9sgL3FoVZIbV4s1L6xxnNn8s9ARyn+thdQcOaDo
6fxPLw/ewGx168vNtCXcBYq91jiNWYeOmh0Obnf2L/kqsq5UK7lC4WsMpfep
60QfuaJJ8Q80OehaIAoWjMJh8Q9cKGc9GpaOM7BnwxIS1suzeaLI7YFqR7dN
2pgfsDUGh67mnJkyB+1iF+vu1PtCwOEVBvR92pJU/sGSTSeUq6lcIutCoSJz
LGe/Akgs3nXpIaXoUvRjwSnePurdi15xaq5pkiESLSXwb4vPp+YU4ejo+jeU
VzL85Nurt39sFGR1GyIzcCs98bawo5QYW+R5up4xbVLLglTX4gZH/7FrMcVr
T2dbThw4oAPiq093KrxvTE7Q2jvM2FFOz2WrdXEBV3r6uVUOTQ5x2BF8uHtU
k9wc49yLbdMaSlg4EiwoHH6y/29V1Cauj88NhOJf6VA38H4WYtDH1hEwfeO0
3T8lvz0/zw48iBG3XtsvEImm2JMu/U5UssNkJ5CDl8vFF9k/SD9+Ah3HibVu
gL+sl/TsUSkMmENYt8SEw3taaPbJUSguPPlQciQ+ySacA71DmpKMHNN0Lhcn
/93x4AtikJ4La3+lfWC+v0VOUULgx0/fTcLKa5ukQkqe41TyI9YKsVlD5MSt
znGJ/PjWJQGbQx3uxn5gD+NHIPTjCUGYMh7nNXjXyl4WVDNmS4DRC22E6BVn
hfcrgvJ3+/knCqTY7/Z4rKWWs6imnjv7GZaTaTm3s1JsfLVN2NakTrvadtVU
puj853sdiU5aDbDEAT39qEqC/YGnpYU4W+Nx+JiM1VI8Lc42F7atPI8ZV5EQ
E+0bY2/3uALmwiVdXxEjR8JoZa1V3fq9nvrjCWa4KZ8/eVLdUIl6xP5gauvm
Ub1aQQ7ORWz0JJw39LDetSXI1y18UsBHa1UN93v4eG0AME8czCrJLiqqrLUr
f5JHZnWepPpfKLjJos6VZAhsge4jm/xJ07NaMMZ5XPsJv77kuS+15I0RrOnu
aFzMXdHL+53yzSZmQzCcUvTto3UghPnfn/9v/7M4aBNSXBSaEoWE5w+FAylD
A0xvPxRtt3t/9RrVi9W7tSRcKSF6vWKicIHRkvqEm0ojo6sj8vTfEB+I39Zb
xTzjDeUTiNgDx0icZPCgsjWU+Zr3zNhb80OZWfJWi5Tgro42JPFpNOt8WEWn
XEhAwjeQVLdCjLSaILKOZzpovNp6ONeeSwUQIoglmn2H3KTSlW8F5kgO1Idc
k6FhKUQy7pbEb2o9VSSA0LGH1Ix4W1xWulj3TSTrGWVTetuV7+UGO374KnFl
rWKK/hGz0jMdYyokw52ZJKEQO7nQaQ/hyqWgm9/i9L1XDWKvO7U3ogCMC0LQ
XWX36n7aGp8C3R0XpUQ8W7iMzcr/Atq2IcyYxFxRfmzyVvOG88PxQekmPiKN
keFqvkRLWAxqYcIr/1zZyN0fLawG0mqTr/glXWCPI2RINLS/hBZJ8lUntv0Y
/wjH4/UB3OPxbWcZq5lrIILqqZETkm0YnXCsZT4yN3wk9XWql9VTpeQ8Qr1X
tmG1t4xYTwUeI0deV9tn9J2QR3X/qUatMQO+BQRV+WXCukDDjDbieyMGnwvt
+QhvV2lxd7H85PDYnpZxQ2x1XaWPXDPL7N+yqJp1Iu7c8HonNPfvdpRrYeFY
kV1f8k3LnOGAE7KCcNprkwJk2Fuy3SK4gp4EiRueNxaiyypD094bGO2aH4hl
MWifiz+nViIdaeo5gq9Ac3pcwKSQHk4LcvcE41DY8vQAxBD/7Tcg0duW0r5Q
o8A0Vt1q1kc2CWYAPX2OPG9U2ETwAURh8pldUO9aUODeeUFIt9DojPczDbv8
6CmUx0YinbvZS1jUrmBhbtbrRVcjV3IP2ySeMTtYQ8QV6gmsmGfrz137siUg
/fAyIMGoPsiCIE31mEZda0WOD4Xi8CX9jxbHN/nAJ0zUIhjdxNZ2yVTapUiS
FnNBqyzNekTFSOYgoy7K+JM764bpDUhheR6Gbx1IOchJUEDJ8Ed/rvsLjoS7
MaN0vsGywCFVCB7m7M7xKxqQjl3IHga71jTdLEDz+7gHx6nrMXi40YDLvpR+
Fe2Ypb2hbY5E3k0YnePNEYcQkmSNjMij3hy20hg6m2aN7+bVWaqu7JvqZ0LJ
rnCopyk8GV7APWhzhTXIgg1VqMETWr2gAqvwkYXLYCN7hAZnlFi804I6OroD
p0/ZpadJxga2fnQOFP0aV4vLCyVQA2p8PJ/LPm4X9dqEuXXpu/TpQBhMOrpl
6AtNr7BpAwDrRDRTTCeNf0CkvtPfXJmDma53sQs2cYmCkLmCuyu9QjzSgQUK
5Hi2FWuIK2yGTR6kPGdCgjzS9HqFvzkDXMci9BuOUF47vEYY9jioGCEqMhgy
AfPSDBuR+uk1i95OtxDoXz/6h6Sa7l8y+S+IQhc5y36EsQiNyGHSahr7LayC
9v40jLBgJQXvFgoui9MyB5lrFPb1u6YTtcoY4Q6HHjEFW5i6WIL5BllQAHqt
U+wIuwJHoStPpujgpNK+diP839fGMP89oVlQM23BChl5FWLN+Bwj3fwg13bI
u+mrUjn2c4h8fDK3q9Ak3yS43vNKlEpl6Y0I2QBIfJZl2cFpeqe+OMD25y6Q
LH0cNi4cCZ6WmKsqPV4uJToLpRCU+vSKxDi78XeRYSgkvJIYdUuGCLgjcQye
jYjBzfHRP15VKjXiCc+vHptsNHfteKt+LhHWWZM4XyrMBVgI9Dbtlr+TfH58
ArIXdwdEui5IEvImSH4oEbSdQo2Z3ViEUweZtTVl/JvvsTh2r8RL1+56ottM
kn5bTOYr18yviJO38xgrdsLbOyuRtDwX+QRZRqjtmHuMZ1uAYL2Gr7IZnkX/
PjfaXba1ZnLFZKx7hSYExUrG/Pa7Gi18uSHWRv1JGoE5WV7AKg/FR8f/BBuy
+tI7dy6wzMB2o+1I+0ylpb8bT3qyCgGurR9WXVo+fBjeWH9Z82SKhyZujtsY
zN+hfCxsoJUozbpptNS5BiPJ9I7JHqkYKrlrfrK19n8Qp05iDbX/CNiFZdsG
9FHzm2+WnBLaztrefK4Kw2Bt5rMlOlUvEhBBhJ8plI+sxxN7E/DHcvfJyTNw
cM52ya/ogUH6kKiIBpB+dksYd9n95BDqqClZEOWwIJEk7rOpWq/25hWBpFKB
tGYZfg27c6vgfkXYXUVFqgwHAaf918ZkQVNnjZgUWqz390UNENnR7QED6m7R
NXO3OKgmGhnsNtZus30IL8E8Fo78ptjgKO9jsumeeqRBvm/m49umLmxeVLAb
e37+oZtzRuPD5ZyUBcXhlq3KZeB0Rie9WA5XHSpD7Y0q0wt4jLSAEMioL4ng
I05KMBxD4gSb/NahM5ov2YOJacjc6rsm0cjlNJs3YFak2gqcLztfqXhPnREm
rws5VGAC7xyutuFFdHUabmtnhnXv+sMLVUjIis2csyH48moIY/d/BuC7emqB
tQXDGAlZE+L4USwoMHYrJUwDVfndSZh71gKdFdYQ4MZX3MfRdU5vUJIWR0ND
faZCJ3C9Q4lkit5U1TH0sRQfViKmb1DqsKsliqg8VaIh/tvsMejj9RNpmsJ/
6tPcrfhr8VbTChkVZZ143pYYp7UfxNhZchGhIz+nFHhWy8Q+DbtLZ6+OTI6x
KRMEax/6BBkI5Wr6bsUj1wh+ykz8DLn9G6abCanjsSeuUgQpw9ZSYVEG3Jo3
/mFAQfdSDzmCYTzNyOVHQo/Vy8tCdY+OY/GMCs9STPMUpQDHK8/aPqm+T6Kq
1b+GEdlFFetRv6w0ChY3vZfliYtS8qWO5Xhk2K8/HYnSMbmvPIDu/pHYA9LQ
Do7LyB0dloAU7gLQaCvu6HigKZQbmSFGAcQn3Fbjp9+myCF2RpzZaPR9uOCS
1dMamahBxb0nUFAAToTJW3JDuKQVUoE/Pg/ZU15F6kdXoz2ZItLdSVXqbHq6
hviLcmgNfaqmYusvowt6s/8SaUl/mJBFKs5bV/Zd6QbU1fm2MrDYPw7v7uj6
+1STcZNtAO1crYeFJ9MNVbwJaDdSUZchfD+1fSWF/vMJFEVVBNzvEOgoZ7cI
MMa7ndQwV8MtoRIBNPJtm2iK+eZTWN1boJfiQIMfw2DHHSNzbMHzdC32528D
ETBGZHFYX5xKIJsw3Nmy+kzZ62jOCdJYmksDUhBUOki6mxVBVonkFJdnGIgB
qcPXBZrb1sGunw85VTXBhcM8ePDk2Zt/1VrRq1dG3GYFsApH68/mZu+FK/aM
ujGu82h+9MYthBYElVdJZKS5g5FqSmU8ugX5BDTD/0emCu04j47jo2soGPtb
JrCk+DRNVx949pyGP+yAQN5bV/9hjkEV8viXjqWg7qgxY/rnJHbAa5XMEXWo
9zH87GaxeT2vhB1o04PoqR5NX0IL8+7VgcQxtmE5Iik1l2WZDOB/iTzl10eN
VFq8ZgXRxbU4SB5T57lT+RcQYrr5BvEfSRx4HOax9nBfXVVsccZ/iQW6i7ct
hor6FscAwG/aQn2ThMzpOZw/seNLZeeyuVyxMXv6t3PG3xlkguvbhP5ObL8P
YQB9cGjTdWZ4HxgFjhinK0bZPyDn1A0RX8H5IrXX+MCTOKRdorIGJHiPebTo
0wvXxmwR0RoMTnKOcpzzje9+yt3OGCZgUAVPUGZ6Pn8tEB/k4OJgdwhO6G7F
b7rH0p5q5MrOx8QI9o5/2zpn+DSGvaz1t8Vdaw9JnddMmNx4TUCw/YqWNVG6
fDGtXvcsllibBund5/kG6oheDdvP+lCEPAlkmI7c4F8u48Dtft4ueT90R+h5
saJfb5UOb2033dIUdZk4cNUzUaCQe16Jhe6/hrAGCRnfnvmu5MsleQZ+3VKM
dRsNRLkgKT2cnPaJJpIEOiJw+7LGQRvxm48RZ3LqN9fo9hlU5w4RGK6gOIsK
JWM9+32nwiUefsL7PIGUEJ5zm3byuuA/YghJ80IVdubqXw6XJ7DZNweyrYt1
NU7QWuaBy3NwXQOhDpTzPdzqOiDZ9rIhWsnsmWtKlfcEwDEmlkfIK6iXMGqx
dBGG9Iof6ebwhsCNFTTwkVlJ83cRyXrT9Kgt4mlcDc/7J2zPk8cu99lV5zOn
2Dh8dzGCQMGNgJ/3yfiB+McXezuQCLV6diWalHcxSQzfs2FtpjnIHgM+0pJD
8qcZ0IH/Ovw0dUM2UOPJvE6V7CcUANq7sQDWXu0ZFBxmFPFKzaaDEIZbIgAj
dM+JuPBeHx0CS7SZWtB2yzMFjm6PVVsth3g+wBL7zcIvwqGju05/kGA2DQJ0
M6TlRHQR32WM7jM5sURqZ4sTsPlGee0X8wLYV+kLAi/+Kc+AY+qNeH+Pa9qr
gPuyoOpmfQ+OeIC9j3qDoAD+0NNpQOlBvlc8Eb/k/cjbZ6rbZwTOUHAJZfnR
bh5i+aeukx618qf3K26Z4wREVqNPcr7sqkmdy2cNjMeo4d/81j43GVnqlCl8
B+pw9VQo+2blCkJf4Q93WsYFKFC4lHBZV1Th7t+dDvL1I/DywALTe3tKOkny
X9XzXHv0ns8Xgft2+/y/+dZW51qdnboAFcLP02qoYe/JyYfmMAw9wMMLwezG
5o4obhvq6cU8Oobqx5vXe1XStdKrge2o+XbgMO5QpaRc2h+P8sCSYUOC1IPR
IMsljhQZ9Vam28yHYdwZrKMj4WE7eZgqD710jN/I7H/3Nvb1sIoB4USw9S8m
ftuu90fRifrIFYFHZI3ELthHPFAHGCy/XbNneeO7Dd6Oq0ilqUk4Yq522KLn
2R2OF29cQr6FtAZD9maEX2VdiwdrGZBv2jRvsgYrtrWThl3rTkMXF4BQpmC2
Trvx5E8u40iE7nOCDMOHtgAKgJqv7ivP5T7bDRQ4/0tKsoFoCiOtf7OuKSkZ
IG12nJSRJUS0inSp55wtQkkNiZ7e1Cg4eg3R+YonpMEuf2vRpCyRuRSbnLtE
YyPn+/4H05MR7eZ/a4VrF74EkItb0f2904nSmV+9n8dSBaCqJuAKG1ZQ6pyV
V1hMY5m1IYE1Ha6sJvc95b3pjjiHcYJgJ4mbb2W4506iAZ0OLVoFwWMxerd1
5+tqNhmuEkPqybB57nSM9X75Ptr6PtFfY/ohffXwGVKi3L8t2TX3+I7MKwxR
PdT7iSqyi9mv1pu0+9m6mR4XgW1E+s9iuSEKp/4OqZTZji8BcaX+/70d5ej5
QUaeMvP/ddeyLP4JsOlDUHR7KdqA3SNZJvu/C9BmiOii70RDulGpDjP4gmr0
LqE34zKgXl7RUTt8mXBVbEpDSW+uGb6ujuB6OhDk0FuZAAd5hJOhuQ3WzXmR
ciiJJxfw5nphM647g+AeAfiOmq08UMK59htx0knc4D89VBr9FE3ASytjz04k
Nk3pJN7E2UdX2jF13CgAs3YWfarak1q48AwMTfZb9HGt8fXMf7AUeJsNoNHM
LzHdO5hTAy/5mPCZEzaQXmm1UC1MXtklAL65oXtI0HrwBaKyDNXtpUUaNJxp
ZDM73WSauJThsl2Rhoj0OXWGRxYhBxeZ7zcm0kVjl4uzNAkwkwwW6KHOIu0X
T+4AU9aJVWdgdHKQDBlNCr6mvy6dPe1rC2gZaTVsYzwhdDBVqz4BnqNAhGEk
Dg6IpCj23374OpKb7kBLoxpfg/NaAG+TchQNwQL+KAcuA9mhc17KqW/ClHhv
ym7SsUB/4qOxj5fD8+pKywqNdTBpNcgbEvpFkW4hSnIcLS271b3FXD55abAi
apuq/Mfwnd/0sroR0fhHDcgMKjmjM9m833+3qYJjtbhsUSewLbeHRxYh94WF
6cSTFD7+9HFbcQUFGtjDcR/VAmmBe7QL8MqwQJk7vPUtMGCphRl5QiDZC7Ux
dygw10M+F3zamwj3wcAnMQKd3QGK7NCyIZM3mNmUGcKl0rmUICjVRu6KBIOL
nwlS8kKcMgcoP3H1lJx/ULrijC2cDGbP2vZc4C43+WVfa8rZ3ING9/5BwfuP
8F6GcyTM5HVioCjANRUQEGEULx+7jH6nE5mD/i6E7a00tCbWDBuuKMgZEQ2e
vYy5rnNNJ4THngy3OhiNudH25MeP7CmNKylZLKxTXLnu857gz9eNV6EFQCvG
5y08REFllps7m+pXUvl/tJ/v6faqFYAEFloid20c0o/yCzkK8xGA5W0zTyqE
jyU7gfh+25cTtQVee30oHPuj5BzcKWDxgYQYe9tb0ztE8AUjE6APxQrKYHr9
4P60yWpfVLQtGwfZob0z8CWWLh0F4Yyoe74x6dv551qOu1bdmjPLgK7SsM3S
NAUwUZkYwJ7W5+BVc5YkVUvOS1OGNV4iSlW35u0pL8cEs5aWQTygyIB8b8oJ
AAIfcWP+CMN8256TqJ8A/+/Z1aep9OKYb2TfqpNRwna+/okbmECu6weTluzq
uAJn86syOpaN8TNZMx9p/bOYj2Vf4wRxXnA+4j/+Pil+MZuD1j1ivBMtoz+4
Vsp/W9r8zexP2l3FkeyXVjL+Y1SpZ2nQq0gjNfX1lb0fCO39VC/dElOMIhlW
ZswPUZJ4m/ZM0zO2ULRfkmkpKGeMuDd61NxTwgwV+L+MhFPGi2BvV2CVhLWw
due1wAtuJWuBi0kPRLT+OHP7XL3z160hTC11Ax0SBK8WNcHvxwvigkacSL1E
u81qw9vyO+rz6uj63vIrDMA7ylo6CLcV6dKt/1MPcHsVf+lGDQf+fovPRnMp
V/kIzyQtd9KysyqcnrBgYiSCjpKl9qChNUtd8XTFKQSI/O57PI/DlaWxG5ln
8mVEizvPiJACSFtNJbIcvrrUCUorFrQDynXkCEWVbUFSVkCWEfPp5CSbscFY
W5JfPJVDDhhxJOFR0O5I8hGMeCBvd6HKzfHEZZbmm58VSPRLFMJ9R9VDac2T
St6FcN///jDWggxmYnvDNgUN3Ro7adRMWG1MjML/Sw/aklnhdNjHw7dfWL+d
UhTwApuxT+pFYZr6sOKlIECNy0boh1UbMgBSXZTMApOaQu/Pj4tgUvkxhYXc
EY8H04DW6LHjtqEFXz6hMymH5h5ndFfLu2XWhlORONE41YvpTQNmUrp9T9bH
tke2V4QMxsI5BMkboECHUP5gsscj6jMcWPCK2DIHCdtsOIXhMo7hFh2dCcEA
PdwwPMgH4A8AtdRDTpf3qGE5H8oY0hIg36OBfg/ttLHLgROM/leC/8k0z1X5
PrdE4e8TzXjjnPhriMg8d5y3hoCMmzEXF7651HPKjkrMBe3skwMvBp931vmG
TA4NyDo8Cfh6H+x1ZkoSFuIOq2ko2UGuOYH51/ChOSF9IWpWPYjqWsPhD2rc
GTmj8HhPTvt0+SM6VBlg7w63TQ2cIKPqAXJ6BMkE6yXjaIlDYX1xH82z9eYf
BFNi8I+c0KNzOMUJbRjBcnnIyz/R+HqX+jxHflvh3+S5+HcJpFOIF3Fa8BaG
/bDxkGwjDNb612IuRQiHw7yFDAJaBsjdMnSkGjUoFiQ85BV0KJVgKoa2QH1V
ZZjxuTU6T/KOhumouVuydJ5qu86/H8vyfg1WkiZPBvCay3MgnFqWiPjguA6s
HnLXcXCDrB7WPNlDOB3N8SSJjaZrnpS9NGE7S8LU1QCUEdDlPzcVchxO/76V
mECZ1Rs/l8XHIorYCrMoMuI9uuEJBIRYLYkPwldjulpIh/c95QmrUa2MBTOB
aPDpGhkWnQTwW9gouQ+jfcNu2YdC7ELh2Hgq3lq3oJ9ygrFJqac4MARCKCBY
tPRoNNDLS74LTX4dTsOlj698R52xqD1s3Lwi9olVC2XoBgEDDu2EFsPJYIdE
6xTCpgwBzdqBYrKCX7K5jHF2F1SIppHdIiOITAuutNi2/a5dvql4gf7K/EXR
h1BKV0j4lDME4zMvwZ/YLkR1lTV8JacIfp028GmtwwGKx4/LRFCxGjnV+qj1
DsrZVsv3o9MS1b42zUEFSMSx/MEL+74REvZZCII8UJ6WMeo+qZk7TGfVC+Js
9xNbw2U06gRh1zYaz8brQJNasAb66P2sAoCf9WEV/VBI/FtXLnFzVW9gRodJ
zl/lhnAhcW4oEOe+Yrj7vjRJ5CgHbpVvy+JV6gEfeN2vIy+YQnU3YSib9Bq6
C1fm8WfHIvPTA6usE+t5tpOC/ifVD4/qZ+TAjHXUOQjHmH51OOAm1cPXimhM
4MZRJcty5uKzm7nE7iP6BKTWz7mTbIN4+PZzrrj+Igf5SOLsF2q0dGK0hs2d
Z7hbIsXFN1qHL1xtZK0k9u7TqlgGOlQ1IsY6sY2hTmZ4L0CBtF4y4dUqE0Ca
eixnwvkg2EX/91LqoHD8RmWrDOUCIFolgb7lvB5+86HlL161IK7BvVOb11nz
RohRbV/ywF2Epzm54CClC0wSNhVzvOh6GR3m9zTryThEIA/vMoIMF+dje0Hc
jWjMX3e7b+2iXwFjG66SeNpWzyMkHZoSKJy0+CPP375lhIWBgadI1n+NuzX3
K1UJPorHceIGYXtp7/h2evDXmC4a5U7vJETtdcEJGm1ELxGo5+K4+TmzJUT2
Yrg6Dg4eACzril5XlBi7RaiojqwMxKqbnzYjwBtYJuiYhCYXj3by2/sSzNG8
+h/aBYkWTBE0muGcuC/HAaQEg2f0xOEm+19m8xajkYJLNw7UvmnI6P85ri0E
tKPvTYXFp71m102KB0slWPvw68WIxEmzm3WayICypKT++jgYo0p06EIyfVOc
4GWd2I7PmSOmQoFi2bRyztrYAGtdwTS3Upxq76nnAtPyHNClfaDxDmh4D/r4
G1X+cAPjIz4W4MtBZgXqD1FsedyGh902/4hUb26uGUJnQ9BYGLPqI9PeeQHD
MXWclV+5GAtiwJmgM3pnLq1r8rlVV9He4FdHwC7Kdo6wORFh6j7N+Y4cUMss
yTIbX1ibsaCXXVuixSNl4cXnBxNhBVM8lKbqB5Pr19g7em2wz9ux4ZYsGx2K
UxuMaZG5ElcAq/6Du51efs+4RDMZYB/yhACMYTRRXo7Qaq2yn78bJlzsTVJT
QMGfOUrqz/Y56Q+MXnWc6/2AdXn4iRVyjKn/NH+46kReez6TlTAwE+Q2XQmA
a/s4ASDmKOxfYECHz/0ggHUDZ1AY/2DUKnsIuWQpHfnB5q+BV0mKq0gQiZpy
OHW1LNiM9SNb5drJ6fCc5WaunSD3tw2DVYpp4wPX6FkiP5HjGuLEALpeus1D
jHHhWVhE3en5heGbAglf2GE+a1SM3mIykyevLk5ra7WVhgPQ0TwuI7OM+Yjg
gABipbBtUseMWNnwO7lnD5lnA6xEaa+lSKONU7+Ota2pC2fpYNHMq3NeNaB1
ni/B91iGc8ktJLepa5xhX79FNpmQecAZvOIvy6r372QAUxNcmip2Px6jOiKu
/FWBAFh1oO70eJXKaE0RlosXN5t8mNaoLtw9eObbqrIpi6yBLJ3ptAK+bhoc
qHn40ZX5dMXK8hsBxXShOmKBmkKwLbHp2mDGJNA4YMIOzfu2kI4RuLBOyz7L
GkGuUiDhvdKIGGjCiqu4w9OdUyo/WQlaUtA+GubFQ1NJgSuIHRt88bdo+90Z
Dp94Tpyf6dJOlA8SYmEWwZtVaR788RxeTN327qyOdeO1jaq1VQmw9cI6rb1r
/4Aqc+flyP9d9NFolFD5TETyga1N1UitzolBtpGJwLKL0uJAEsuk+Hb3XeoP
UndxtfzeeA4KW0i2f0g2oe9CIPpd4WloW/AxQKtNlS4nOszM+0aW3cCQxj2I
p7qqgQiLHnt6L+IrQOEs3S1deO3TPJOio274m5UpUdA+ng2JTgL70BKp6NM4
sG1LVR5XMSkTpHaRooLu3ZvdtcRo4tvpmPZCWwlYYVKkmcJe0/dxxAWbi1d4
Innz5PiGOzr521HxwjPSQAlqAadvWGpkgaYFRXjnNyOA48Z8YZSGnHZFQoQY
Tb+b+2QUq7qdxLYecyMU72uINBWcFb0R/WlQJVe0LuA/8mzgDzjqkBVD0bSc
a8akNjS+DR+ix3WwNbg3gPixN4EXTliZ0ejjVpsZFtPqyhi6Mhx74giD5b7z
ef7S/kI/a1Wd/nHqr+FoJEadxq31axwDLUDG2m/QoBbnj9cx+9l2jLpd/Ied
zJXnAlrBtYKALONw1yjArPVpOwwfmpgK3o8aUtik/MvP7QdVYzZM5G83Ha2x
WhkqXxh28RQ360sXtrof7GPsK6hStFdy4VrsoUwXKUBu7hUsWBYCg6fVxOAY
Z0auSaHRaZhxgL77qMzMCHd4GNRPfx5LurnCSU7+rKZ15Eg0KcJp17QV+bnk
dMObaf+1PxlS4/Nzx4FzHT9q6IpkgrqVB1b0ZewVwlLmBMAQgUIRBKZiUo5g
SLF2u4UehIO2dVy03A7CSUvy54ZHgjwAzJ158rtPP8fp2He7iObPZQddyPQH
Urjz67tB4//fccZWyLTeRlW4CC1gDj6hfk+ed5Gfmb9uNFda0+lqm/0TkIfK
MGsvOoK0K0SIJuuuF1KRcTzjg0IpYs3e4+GayP2LmCF2ujLIQk0r7n1F4BCe
etlSSdWubibtkf40d3dtSlb3kDTmwP8VLuFQmLNybqq9A7r/SXlVe86XLLSa
uyR0/PjXkhRQWJUAQ/Vw6yEjx4YAwX2OqxMG0P9GsglCEHkxwjAKweJRneSq
hreV8f5JqlC+uKagehymdIdWUI0OcsKQgGUcBWy6QFh+ltSemQRAkxs7Cwii
sITOGQvBcwkcKjYbDbotwYLNDAlIZetjEudrc51Dtl2c7mkEgrKhD9xH6F29
PrldUacuZ84xZJT0AOvTBHmwQ2W1vikFXSaeLLqE/mAilOMSWTVsRdZqBJeO
GzIeOMMnfz7Pq+9Z0rqOLlVdW7RiwqeALuINZoEgBqv6ZHug8TXAprBc3BUY
mh+Z+HEpcX198R20QhD4xpXZIc7ftKv7nrQr8CMSawZw7bnkjxiMrmZ/qGPj
lHFfuwa+nuQoEDknpG/WdKQ/Z3PRLiwK4DWfFSKE+Wl3nThJIesrSqzi1Akp
N3+5EyusHSbIX2zaSV2sGu4HlXGebPxciMQYMNn7AsfRG0DpGetzK/z4wH+g
iM33DCgOV3vIgltOY735ht4BaL1ibC1Qxc/ZUQBrKMo8BEZdKx9ya9QUvvv+
KhV7Cus7grPGqJ89iHzYnKXMD//rxEGX1mWHgKKG13iNCNV6I6JgxHGZW52j
lcIlujIkH5EkO5FAdqWC8vAxDRVDpCVx1uoIoqXXddO3AfG1fw3r82l5Xvrl
cFN4a4EV7OsFfPTQWAQk78jyYibqZlIendkm9p9pHQsMMd4dDoJXSpapMQsN
E5QTkz3k29N6avX1+SDkZiYexLfJxgqAlulzDsh64UwCIdlTbH8pR4ejyuHX
QafFBnM7DlnQY4qmFVOdaN9v4sk9VykpQlga0Wub+OQj54jwncWlV4Yl3oxw
790rq5OBH4jFLBwaOhrrumgBa7hhForPT2wLQHOCuvCClnVVaw6JtjrdO/F7
O5soVugfnNMYjjRzoVUDNKtScCH5W8zSQecFxiZTTvRMY5hWUkAcI9Fo5EZw
TppuJ7LMFN/8OwLYMyC4V0n75JIniXD+Y83C3zFXCdfYQbrqY4L0Ysfj//Lt
uEZc09yxoaX3CLzo05QT/ip2WFi7pmexl+RChcFT6/PmDJSpWTPV85NM77xC
/VFQs6z5E8LKPYN2hpz5KMJhqJDnpaW/QVtr2FuToFs5ZjqPZwNE8WnvvZoN
nNRs8yDWw9ryKGgbUQB7U00xsDcDO70Naxga1/XiMAWPhy5wFQdWS6Q0s87F
45WtCjlvDw2iP03t6/JIxz2IRZu7npstGeiDR8iU64mw68iYjXVx5FtZwNJx
iwZwtoWeRPlWBOcM8nIP0bQJls82efeSWByZh0dB3wAlFPYWY+36aRrUfU54
3owXFlAKZi9slVZEkLoHGDjOW/cAJ7VL7Qy4cGMc7fvHQ77QFjKlFmUWQNCu
/4owDDvJXi0uBPD4Fdv1VEu6fQVC7qSojeI8jrrMWoIdzLssAM9yabOQSEY9
g7xTDARR7dtHStXQlXK8xRmqAyLBmq2sWevmHHPV+hlQE1uZi0kKvQYGqgaD
P9BDxVMRzq4R9bmea73MK/FaHEJKru3t4/Jo3bnWddM+uP2Q20qaWjNxD3uw
/tFFqNl+iu0fRehStLT9r3LJheRVqkyMAIyzKXil8KMVuVM0QA0vDjUFjMy0
Lz4Elm6H3TfksrUfqYT9lfi0XK1wSuaOgDplk0aa8K3TIw5mvb8GEI37e4NE
OW7HfRcqyQJ2lG8WKnhKqzjZsUM2eD3m5JMzf9wTd67rF/PWnvJb22csSJ5y
NpZXhPakkzRzRHrFAp8f0YWebXv5dsGicwyWIUA6laLuG6YW0SGr17GM63GW
ID7qWm+BcmfYz2DTo5DAODkKYNkegyF81wwSMqTWzpUMMONeazv05cfDRVOa
lXExCgCMSKoraYl1Sc33bT9AoVfqzRmC6INeUuR0o1D4+Hyyt1kC+fMXg5ZJ
yZDWqucYtTCPk49QEqbUBMsNmzRml+1aadOIl6IxA2NfsCrlcatOojP7mpaG
EO4njJXlCPIZW97on/d9gArsDtqHt/2c21/seI6ovegA7qNpe0IvznykmaEZ
Nw4GC1qt7E6aiImu+CFJPMI+WRGn86PmZ/EW9+YurdNy4TxJZ1N+JdwN7On6
DOjV6l92ySprVXmnmOcvRb99DCa/BeoVQ5Igu2E4dXml7+iRXKIlKX7yG+t8
tyHLTJ+H6It3ldCutgOpQbSXUELwL3fWMfCr+VgSuKdxY0lUuYCh2zRlydXQ
w0SLzid8ar2xUAQIFoViFd0xA3O+menVAvfJXB6UuhJkmS9qmYwjOCAI4xeF
zserqHjgQEWUHb6S7DQCEYSOXQOHFJ2iKdzrIkEYuiMB2gGZAIveZGhdD5+I
Dv00OE1vmPkrlRS6IuX1BTmT6g63hc+trS58NRSvPDzcPpW7dO7BCuz+WDc8
UKLbpVaLxEIqhZAI6r+NsbNBMzpSRQfxNATNNU61MlKTXwhcrUs4KlAVKYBQ
vgx83ix+6v1SEh3hAEGFOLS9n3f0zNoe8z0iizfIvoNDSBRYW/FCUMqxI9Yh
4cccxJMeM+KBlK9KmQOUeQ02L/40OtfW2qblBTVmMkty+bKNVBdfj6VY+jaU
8t6rg9LpdSezkL7CQHnr/xKzWw6rMzDkHq4Rny8T3sg79qmDVTPmXin8YDxs
6FmVxRmFpxSsAaIyChDNW/2afpjw1N4sZFfmOZdTIsydN8Zk3q12BgWXuG1D
VELZwT1/TUy81rOvF5N5UZWIv4nDjUgl/tUQKdCrz6i/2QW8B5MhenNGI0wS
sKoTHVqDvH/Z+BjtKvEY0MW9L3CLjrJaEu28WWXyTBkLgZJQiZlXnpXaA2ii
wDlVwfENfiUQG8rCMtbpJD/IGieF01n6E53gx9VTXA5VZSndAwP0wy9qzGt5
BwkM0vGMMZGxq5lVpW134JrHr04ouLHPd0JuL3rgCG1En8kaAA5kNNt0eG1P
vuhfRO4IUtGVrUMI8IfBk2/Dm/f1q/EJ1X6plf19T2WAZk5UYpl5/Iwa7SB2
wPLfawwK28ZIn8RBb3XGU+EkN6bJUGpQacRkPvNB4kMLMvN126JtkxQD3hsr
pBQ1ke+lbY/Dlo36gShZORV5S1VD8O2qlBlQshXGZ9FuANb63/+vwrFeopMK
iD9oFfNrnQpA38xMb7B901U+HRhPcF1UkUX5vLkqqqOeYMtEUJPxIIzERbNy
q3SgSakFsHvtArNJwA14mujBfVEWD9NR59bqEsz355hFNS8ys3VpJNmNTdJb
DDtez4dKnl9Sf9eyz/3o/C4r2PTYmxz+PQdMt0/5LfFulGayIWbbREzG9FbQ
zlkicVBCuK0VjkJZvbTlof1SWl7n06aTT7k4A0/XFSaWG5NJTo3ZT8igOSLX
ViUuBgATIIEx4kb3PGv3QEKTl2NtkfCEnl81udUMsePkJ17Pj7lGB6DNMkdv
rPldhJp0Lzy8WA+p8+p+o75rOBcdl1lYFsQWpom1GMj5+9JBFCXmbYmgfYKy
/ALRfA2JhyD3qnfrxtoRFQGAwm6OUYYo5lPBEJrVPJ2cjQ4WbXemmfGCOKn9
5CHCCoXzbTZhy/dHNbwSwW8tO7nrnQKuIAaNGugdE8+q4nkzJJX0jzVIC+ni
TOq2tA88yGDmaBiXr8ZisAwpGYH9rQ4OqVlL8YwJJqjsTfWVXHQOsWcEX8Pb
1/aAX8Z2xn/7duFCjjY9tUGjulRU9DAoO4an8NevaRYPixfPrLEUDaMdgUQV
yeOkTKL9h9mk31O0n2QwdbHwX/yxGceMxd2mrVbrlfM2w+m8bdrB3XI/cHHq
20CwauKLxtdEL5ezJj/Ah7kBYpqDAGYFInqj/wSbZnl+bgQcbs2VCCFk+ZOy
68rxiXW0K+MN9P0LjfNWexZhsffc1/kB76NdZe9qW7PQFzXpHOx52KxSzdFi
hZLvoQ8/z2w8/und39o5PJ0iU46O+CiiZNOfMM72kmxnMhFkw+RFCzRX5/Td
4nNT6DnCBJ+Z7Jlv6BP12Zm3gHHEtmeYHXiuN2fksfC9S9e5V+1Af4eS+CFq
44lvfISOE3cStFuVVCU40CATEcJFOyBgIQRPid2ktj0mh6viJoHc+I2k6EeM
uJiOGB3pFvDDiGcKlo+31J0N3yf+Ayr2or0JpiqOAKMOsmuYBLQ+YzinylQm
Et0GG5BNY8M1Ohfj5LI6BFKTWvkUu6LegbaUr2FVdY8wMAWPyDvVCf2U4H3S
GX/jVpAE2XRbFM0o9LG5cZfCN+oPN36Z88v34kXr9o3iR+8BsSZtkmGsXzY3
rkvwLi6DGt12mAZmTyJcNkgpE6J4nlDSzS9UE9MS/vU+AldhUi6oDQNtobgz
5roinfEZpjfKxsHHJDs1/iCc201I40s15iuDhAlCVtz+l/rhnCLuAPUgDWcM
ZeeFh+wZKZfE/FUtM1NrIe7dUNcFWJWygNjyNE2keN+jQ5e0M8e8Obwg1yfZ
0JcAyIC62ISHdCbwL7OkddR+e5iUbpLytWdUAfp+u+JuMRpvAcX6Yf4mIONo
dvDgqCMEANuPb6qPvmu7EPXAh97IimVRyEx9cdH8v57CugUceHWyrb+juMZo
hKjaNqu/ZdnXz6HUE7Pglcks7oXSNzJcSbvxbVSVopGcAyEJGeoMs156iE2P
5D/he32JzJN4UroY2iix00cmSsA5nelhhwm9zWIXXhX/pLFHe/+drI719BXn
LUisaoaeJiIFcGjcWsJZpcw1eX1PqNgQbcvlYFT27pGye50kevkmd195TVgp
FX7S1Yn9BFC2SDN6BvEAd0GZysS2Q4VmfDvLbwJgakZaQnTEEaj+THQ8FiL3
rqL/fjjHXhfzdyDlabkvZiwMP8rXBEfDLK7zGL5mt3rEiKETCdKyqAJst+r2
TjwtgEA1Ubrt0nww8aYW36QtniKWqUj1Egf4mIh3wq395M2IapoPA7b9iXFq
JcCBu13HDreZsqpKgB7t6Ycq72M+YTun46d0Gu58RaBTzRwC1kY3iPbDcMsp
obybq7pL3voemmL6dYUBcKgjgMvPANtj74r+rP9v1qSYLSu2RGNp24++I1pN
L9D70A+Shugb1Dbzsn/qlgJFW3NkMxg25Z4yN/26bC20XBDzBuB98VP40YyV
2Ed7cQwhYkYHdvIv3iJ7F7zTMf+5EGodxz/Z9gB12+oZH6BV3Xt20ZTG0Mcj
1WxUtgewF9GtS1jrs4e+fLrwmIGvvXm8unSJS54fV6qNNsJkOrqvozoN66fQ
4qRjaIMZ0f7Fp0TXoEJGKVsnK0pkoryzEpMjWGdODtasO0ksZF5upCosFd0Z
PLu+nX5E/20HbzEi2nFBgP6WJMKIWLwaRM/VXggGXorWpFOPgNNSMIFbIJRE
mceSfdUIvWdES6yISJEbgz2zLPN/FgiRg3e0sPhNYPnys9+RyuefItte7ppV
OXyeA6+LrR4i2UV5UvSesvjN7WCrMHruqIfS4ocbsnaOoGHx6jWUEghkxoIO
vgJPf9gZkqm9/HL4p0yEWmljW8ls5Yltg0lT22J/Xwq49wEzgmG1N4//yxtD
EfQnvhcUwsR7J5qLZqjMg9nzmaOrdTmEV77gEJ4B7P7EpupKK6wAiyECFqGU
nlzOZc9Dc7Z672y73IrsuGw2/mDn5LFn51rV0kt/8RB9Qas0SOf8KKSbFov+
GsKMPffOLl1hcGJbrOWM1QNWz37ozScwLHTcw7YQ6GU2qxBCH4w9a6RjSjo+
MLvBWNUodMIpQULjO5mlIyzrJhYqOl8rPaDFrcZlgl1AorntFtA/pPPu8Akp
2bKP7SdNHPKNbf636atBruHIlpmXD/1b06MW/avIoJu6OHElOzFfzvDouq3p
9b8Gb3tcqi66OzRghCu4joaguEIsbCkMuKzWCsvrWoPOjgOIYb7ZaPmcBddZ
4EEJRJJMflEEKbudJ4eJY0+90lFL0zatdml1IPEIsgNhoSJQnJY2noBgEOq6
x7ystlvCfY5NWC291gMVRfXfxwO8q8IbVVJgm0NzVEcvo598X0PjF00XqSCz
+Iuuc/fDQF8N2q6qM0ZQOFWNgflCV98uBfDxJvIQivXsRA6kHNeeyU8x5AG4
31D0NVTNPyfotpndAKwjq9Ui8SZ7ZVbwAado+kJWsMFmDfCfZP9ggAlZIKp5
1AW/zU3sSRKQ6iVT1XILniqzo7hqrinrmR9NzHeSLLsV/uXAmA8vu2gD7BHJ
sH3q4RS/o4PSCigGVuNHjvI9OKa3+mqfn/qynP/oXgQiqKje2JNDSoP8SSMr
wFCcIyPfj36YMDJ4CEfU6Bn2gbVG59nsj5lXKD9mZ9X345XRAduPPnr088Zy
9Y9LGSrgVg0tKLbyjfAzpNxwDgB2eJuYW6hUINPfqWEa8emfsoOK7P2m/icU
ixss2BGsFL/QDKnMZheJPhprEvxcmH+4BeOBQFIEvwt6YCZUq+O+Jcd2uTjp
gS0OVv5Twb5rKeikT0f/ujb0xRFpoLvGkRUZ+tWUpGA8U0TkYVs78ryLb2v7
PTWhSUYkJHRdV1cDhbPvSApz0JnMN9UjMtl8tMdwuUGJQ/Q/5ZFzKbr8eB3P
1oED0MUcYI4ZLXabgKn/ORk4BIGm75QKMCdK2jx8JHFOW90o2pkNlkdjEuK6
EYhJsr0+oLbEehei2JC8SkbgU9y21Sqx2eN0Aa0oBQ/8IquB9EakcmqH0n6g
LCMVlfh8Nyl/zEnWu1UjFfQhfiHZ0UB9Jxyncm/cqnRYxdbq//mpOgFxx6Ru
Lo+KZrfeY/4u+jp3AytHQQQ80/Ys2SV14Z2mEBi/q+Lnq105hQcD5BdMC5r1
XkFSBEVTz9wmUcwk6u5biMjR96bcb7KGfUfgYwZk60xrBW51S4VDDKbfxp1v
xIoICYYCpEx1GT+V4rXPcUM8sFJsl5V/NpL2SDGWttLBLBVB1zUSXaGeHO4q
KkZPDPgUOHnp3RwWWuLp6vnUXnbt2+r0pH6u/j9PwnKO1tTOVJI27u7YSVfc
WgJxwKuODLAoztF1EEVvFuZm0wtfUsSCC5XOFtEsfdEq4bp+Q1MDL70pSR3R
jQYvbVkgEisNI+2bEB4unpnPMbIF/TZHFQXDjbvwSbP+MKnY6Cxo2nuhCydx
SgWb3SqC2h0C4+inGIX2UZ7lC6CrtS0/9oPkekSp66Hg/vSjWlUb1d8DFDKU
KLzdkZcoZKcG+2E2qO2aU2ULB9WTHuJDz1LNW9aZPpSgDyzEmdQ/mAnZjhSP
i1JFSUHPF/Pw/DrGeckK1fFbDqcqLBVtkhzDq2bxNd91nhK2qJOYLZ7hrjUN
kr8ZxDzeHcArCukl4Wln5xA8spIjG+IsRzICbrPt7yE/tPYsXDPIEjSFSVNO
7HrHLry1vCaH4+W6Nh4Ry4C9kC7bDNzWNLvPtcO+Jnz/zC6V4zI9k8fYvF1t
xS1vMXb9i4pw+jxokXM9KBJu6tnug1QvJeghzpaDp2q87QrBmHa0sPC5WWOJ
IBWrSkYFGXBMG/jT1jc6+O9j1jYr87h8Ol4uSNTq2tZ43TdB2jvXdeDjgupF
J6HB1xjg6a9e1loTJI6KiDQpyPpXvQhORuSV6H3oN9j3Vd7z/snk/RQe9PHD
vbXFctUHcuRqBQc+BRO25pSTxXHEvEutfQwv4o0x6PGXxpYND8gSC9MjgGjj
J7C04ZYoQyK7Tilmt7kZQ6oHd12Nz31fwuOQNAYmGUOYNtAJYQ+vQMQtcVAp
cM/BOI1og009PcawMAaXZ5e+KVtBLWgNJ+0hvCpgvr46jVKRDr6xXSV153jQ
XswXuRmRuU4rUHvZ3x2Af3HhnlLzZ4dQAKkLS6f7l0VruHbscC8BZPoOSQ0I
YMO7Cmq/ML3sxaSelfrUzXlpA3c1DvrQKWFFQwX79o6SbeU2Tski0eJviYrl
BBt4M0LQT5ytul8yoZkSYn0zmwm8tFG4yrcb0Op6WFwgyym4oNWA2jl0Gogc
laivB8dFwF4CdK2lRUE36+ED/q5lYzv8cbk1Kva82fu78QArdXqO80Xk5Ihv
nGI1h/VkxEexuOQvZ4nLKyb6v8N1jvT+MpZ/kKdkdV7UmwZwuf15sfxsEJED
2tbAhxYVb0qEsG5Ix11m2uqUak4Ag+/rIq1syjuza+oyMxfywBJo6gJmn5Lr
BRKbuNmQeW8c7bIMVNz74C3xbV4yuXvolBb+qiZdSRH0Pk/82gC3WbisdAkW
YRtIAAQJJrCIIfkPz2kFNL2U0vGbYV5dJb2JARcpuMEzBde7qSPoT9Dbz17r
DjAKqJ8DZMKsvGwLoSkt8JjOuQEGrNTqeqTjZNj9GoFGayaxHCGGcax++VNj
HXCOHxS8n+uHGAGG3z6Tq6K2SrUJe0NtvSINBmpqcrbc6IC+VvCYJAV68TXD
nOzvZxfZmRaL0rnpwl/FmAd+YLnzWPZYmwFh4/SgqCYG+d3EBp75pxGcmu4s
OT6I4m/j+p23kwwkk5iRsYKX5Zao6a56B4KrXjl2ZkDegSkC3mtXJymsOHCo
zjhXGTHxF90b9JYKGd1UUee+4bmZX7QoSDm82x0qcZ+WkDCUq66H0GnLbMIl
qYFqnUzw4t8MiKs7BVQETDtIkdIyytXNW1dFUrRM/AltvXNs7AOgAY9jD4xs
fYAHsSlaGxmiwg1bT6YmNxdAEU6Ofuri42t4vqJt2i5oheMlJ/KZCB2IpanQ
chLlM9UB/q9FpHiF6YrLRYAnqcjKjGmoV9IOHOzQYapH2UukzbzKDHbvNaqO
P2osxOltGTa0+heGeMQxG3nHmguSQXYWaUtgx7KZ1kJZ5imINTkTf9Neamje
EV6mhYAH/R9ZUc8g46dNUZ5HXGT94MVcWuKhpfSceghy4/aA+Z+3bGjRnXu0
AJtsredqEsdaXAeBfTzW17hfMV7xCTJT1PfcVKiaDUJGI+MHs9amFk4C+6EU
pocR2qCTWIXe09i7wK6Eyo2xOjo+QSB475Rhxc+SzAu8YCz4X33Z2BZZq8vG
ISy+KKhQwY14F7WKRc5R3y96fEwPW8ZXAHq7jtjb+BLEHvq0Z6LNigVOYtEl
H7W71v5JVW4NEfZ7zJRVfhmRlznEv4CK8WRcQBrMU5SfsoHS2mxhbcgJ6Qy2
4UymXe/d+bxrCGRKeGb1m7QuvuzLPciSTmzM+bnEhCb7qKNtiU0blmdC4FpE
39Py8KM49VVLB91sE+CWfkU35BDNZfv85J0I0b+KqwGdpJY7CkIqjOaDmmV0
oedelagoxxiBFLmJth8qa180lQuwUKIIZ1RqvKe+k4KKUlmnbmxXgREwvDFE
kmEUnvYeqBGfm1+dIrrauDD5aaFDNlA28tQKPNs6NUl1KgotX+hyrPM1yHgo
PMyCohpiE2Gsq5ysl02K2ErVKOWZ7P/7a9Tj1dTkap7IB3gs26JAtBQlGcDM
cWuJkWpvCFvqSqVpd7khwK8VQCP9jByaJiYEutVrjRe2jDlpw1Q3xBVdM/m+
Nu3LdWmDfR0oJoEqQbXn9Zbek9yympmWP+SnheMPYZaEVoIX0+w2Up4/TLgU
aUQ//xchEdTGnzt/Mc3KsPlCbYlVetg+EF+2ybiuHylMWkUlUoj8JVDSXjLI
VrjSg7Ykv9N98gdF0aznL8MXb5vai7rgIp4+nTltxzlRYpj2/icVJw34Np7d
zgNRCjDVQI4QvfCraM4MTkX6wN5bGTWRXLLNQR53tU/xRR3JZhsJVpfcLVcO
WmF4t/gE/zmsn1YMA5XtqvugGlV4Jey7FGKU8Yx/hugSg8Bi5OMInERFfGV6
lkOSuPMnEjl0ko5ikOeuOCkjiAL4R/iCpNR9sgvr6qE+H+cOiV0nbw/yXnhi
k8m0TmiWSLK16sSrjjjd5eQB51nb1/IYXGUngZjzADKRBxq+oJFek1qkqw7J
whxGAJygrljxBA/se2gj33BKpJjY3mAUtqmGfMfl5u0xWMfAvskg6BOK37sz
ONbSijxd5ScP94kFEsp3HBaCIgKa0jOl47DqAy7PlH1Kfan9pNy3XUnnsak7
sDsAtWljeyPa1B1Tg5LHJdejMX2VVAA4uIRsgYCe+bOIQ+2E5JLjdauhM/Az
F+Sca47+vax/g1QD7lJTk/zSUigbjdlXXnmvnMUhexEYLpr2fSVIP5h6qg/C
DLJwRQZHQCiJ4a8wFzjb9rmqXrC4cWy2Bu+jPKG8eNMGr9HaMGEzNDTWfXWQ
rn1NaVsSOT5waJyZv6q5bmJ8GAGcgCwVgS2D9bzE+vU4KPUiWEB33aYrCStj
BigY6/YsYEyHOEm03N+cSYU3ss8OBxfVdfV9zZzdGwlXkgbMW/5iF5AkC/L2
MydhRdB8x4mmqAftM0iA3VVMXOJgGqn8wGOSjAc7CGGx4qM4Es50dxMNH/HC
6sPJMZh4z/LLO9erh7YXq5k/Y8hnpCg7TEjw15lpCkT9PYLvFcuEPbR/J6X1
SShupE9Dy0C2UGId6EDd5QNE0f2gXd27FuyuSf6xss28EatylziiZTeTbs1X
HfrB9wezI00fp0T81uT9rBMbwyE7wF2Eht2i1mN0WWBZKafkG/rAo99BMSBK
uWYmdCVpq4n38bgSs0K0rfImNf4jz/zIlJOURhSely6/5hw9K5PaZ6Tf5+IY
8ZIgc/dIw2eNdHff1gwctnEJEfeQIOqLjw0XElqWuBrMBR90II2+3CF4qO6m
0s0XFb06EoMfQ5MUsCMpne0fx0pxLH9jHyDdA4FhAXR3vRx05Q39SXzs6ceg
yKolTVCgVsF2+2RoZAAyNRNQuaRv836ImbkbDjfCkERfgB1DP9JRR00irQub
r08GyyX80Z1sZUwCW/ctYxKWNlVrt5D6ZZWMC3iHXGF5vdOpTqpxx3TVXaup
XuA5eDEwh6eNsU4jbfLc/xKiXr1hoYP7kVHtnYk0LLUqVjJILThVRRbq43CK
2hrz1qp/qfu1ZQWnZTENIiUcOSMghIC00QgXa5JC1jY/ha1zaTAldDI0XSi7
Ua6/8js6XrjF7GxD0s3/m9EW5OTnf0Jnb5waPF7hdacS7OdZx3zjzU1Sbpk1
31fMyEEbKIpFhy6xNyU7Ms3UAH53nUHTzOMvO2qt+YwcdjlfsJaVFi6BcWAY
ffW0NgyIZbLNwnMlGlyA5q3R9m1TdiY+b6QTCCRALR1rjVRG2aOgedZJNLbZ
WHMGGWt3PIcWnhh7H/wSGMEnYxTQAaaOllbMo7mzhM6+rjlwn0MabZmRrWig
OKERYqh6tCP+4yLKQMBSm/xthMU9ehc+GUoFnqQZk/P7E4YjQbiYWgg8oquk
WyqXj/H5X8g2YeWv88ngui9YcJbRM6IQy8Q3txh7iJPheF/RnlMQuhvn/51y
KTAv8wgQIDZe4kymty+kvVbq9Nc8YQuV4j8B5fu8NyzRzNV7pt7sUBeoE18v
qv/y8SEsC0sx2lMw+/vzX7cjiZt1Ynhgyu/bb2mK28hnk1thckR5M/nUQWsY
E6pC/+gybz2dfOx//OwTnvXEXDnoIf/wG0SOgdhDGTA4ckSKjITBzlcgpSy0
V6VJbVA0UoXAwOGIBekEd/s+h6Yga3+kFAKqEsCVD8zbQKVi7i9BmLXupqQl
NP9/8wICs+34DTOT5I+b2kvPLAZ7BWRAZAaWCAPxwCuPYRzlERBaaKwMAiz5
XHfMA1Kl7FmsxwvtQnleQOc0SdYaJK+LTZg5IKW1wjnAWW73IG1EYeOL0rpA
MByNu/9F8wcK2JMZoNS/NoZ4KCJbtCiITVUpKtiDblfZhjXLKx3EQlQEuNQu
YGUBj32I+aTyZm0Gys97a+dKTo4QnF4HLHmhVSl9jj/ek0/+0Ihw/tYS918b
49/RKhSyG7NyXLr+cYrBP3yTAMTF+EL+QrTyk2cyD8pLlRU9wCDLccPCAq1p
Y+KwCtpao+E0OkPDSuT/iM5ntdgFL617zV7yrSoegBUP7FrnlrBS6s1DnAh7
8zCV+KBmliQyonQjxWLUgU+Aqq8gei3y5tts9Nv84QtM342YzvatyLnExVwO
siig6NZCuDIfSR4zyvXVbmeVRsan2ry54SMonhSSuSEHcQPD1+afazLumtr+
zdfZJ4QUtadyRNs0Rp3GItpr6PshQW/avwgm897yB1aybwI2lHAOFbw/wJmN
myPcIvMNhK9JYlNr9lKn2mK2och8CKWoIHpPEhwF26OlFrBwtCXOj+a6KxRT
iCLnkrCoukFQhtSeebsKxLdD8NHSzj15Fg48rdViWK0hvVZP0rFHBOTNK5Ln
l+PDN2FHGJ/IVSMg6XNRkXgs/zDtGzysxRVvwSNMSbl6MDBjaVpG9GXy5Dpr
Si3hiTgWY9AjM0MUq5Ajenr9DU4C7rfpGqOhUuP/WaIFfC2TJztFNq8J2PVz
Pdu/CIWB6ZkmAmDjrnKelZ63glVkp89h+OOe4rF2+DlMWYPeB8mmlXTptYbc
mbmdGywCaXP2geuTEwiK48C4Tw6+pOhIqLwnW9KL+vARnTqhyK8hkINDY56a
OR5fkuylAgJEMPu/Vavx6+UZuSqFI4POZeyfGhYTuV7PlXiAWSM0DyxyhLJ2
yRVMJKdqgil3FGXUnk8lFMDTBfYMEeY4e8ilERZGt95eA+Qr8X1cti9zCet+
n2MjARaQhnhs+QiDeHEiuOEydZpWA3Qzm1wmf3Q+9OACxaGpm/eMb44DnGTZ
6Kh3Lqj2qftc2MkayrIs9PKbWz6RKx31fwRRW63TI+saS21SAFXdH6dqQot/
AuwpWli6AbrEYUbDFblPg5xkh1ZbZ4Cduyp5MAWiclfz2RiggNkvHB96QYfM
VkwFMZKsAeZf2bygMGnmFGVfsxmL/WKwbAuKcAH0FJToijIKmn0JgiEU4ffU
Xtg5N/w9r7AxN+jihEb4hWjIEyXSKyovwI+/g6wLaSYVhjaZTUdWBw1+NS9W
FNg/Tr281pmBi4gV7Jc0gVsgNx+AGqtFrXCR6Tbo81PATguQ85Igv56XAioj
osHrW9oQkGskcccb4sIWGBF+UYVSrOxdu4mevnUGCFR+zRO9fIKFwQ/isWX8
jzaxDTzwcF58KNJ86VH5sgThTKwuizCvXguw9EK41fFwWywCT+hLHHIs6Ckl
0p7OPrV4w3Q8bdJzoJ5i9EGpuoYUn1ssXlOg4HNwh1S98/NQAOAiatYjBqnF
S4p/AEc7FSvcYzaHbUNMJtV6Joslh4nv9labfE94SvdGAZOmlKVqWOf+nO2W
6Wj4Q08PNAi4c+cx/0jP0QvByKmX3LBQcgMlv8ZfIPGpiPafaJlJedUeCbq2
TAHrtvASIAZ3yCV0h70+GiKN7QVBFM92lObq/GgGYapuoRPv84KBNb0TiNX4
LI8ZSlWWUQ4hdQIAlXFGu6VqJsntycXzluFrxX7lff9iQ/5Du0CjKqKmQNNA
JyzoL2+GOg4uwQm/cteRyN+kvgt9ktgcw98KlHgPSkGclhhINVcIACLhqUy7
XdjwsbYij63kZDf01fWgl7yXl33qEQWGcBBgtD7zwwY7Jx0D/YCls0t0e4rv
+3ri4ootawVB+/SIgIYlqQzuoYklZAdbc7Lw8O0ERaFkzwdJP4sVUMGNnMv9
gbDIHwfDCXc/XSEaFFE+O+dQdVWYU9ehvDcffujzi6JnEKgg9zY5qb4C2I28
qvoiNdr07xoe1fis9oOORNia3PrfcHPhYMmGWlPtCrZPcPkzykkTUdSVYBT8
S2MXMQqDWPbtMu3ZkEjwZyBmGr8jPCEZE1B9FUNYVdaa0M99BxKrk/kAnfU3
eysCvfjRPClAnrKV7mWwKL8yvnkgOkrwrdUTdCXElnjv3B76FIfilXfkFFi9
OmxxGtFOM5On1SOinxOtlgEFcWNe5rn9baO15pY4Ve6qWpUzMtXO/Rzt8zR1
5ur6fr8UEZgMpgfwiid4FuviYr0HGKUFWNkOBXmyw+kunHivZeob8e2xvSm4
dVJw8P9zJQVShVDmSYyAptEpEYQdizzFwOnkg44PDNEYx0/jXSq3z+Ju+qUn
4E0Wkw54ML53pfiTR6qzHwpoJPBwck5XEecGqrreG2mq83al1pXiKnfyv0Sx
Mgqfm+2Dxqk4SzZDT35wRb2zs2+PIuFUahjKDGm/fSNPT4esozh2RYHpTFAq
hjCXKmdxSe822XxyPc6xbvCeDXQZlum1+H5ROiNfkioG0PplQyl3ExjKAp5H
xvi/QlF+n+6nMZuIisKYU/eoZaQ6txS9P8/qxYuFE6qIiXe1oHpQ/fhOqb8t
ixPdMQRAnCNT0h8pMGDGNiuhP7eqR1mHZewWuesGrHDpeXuLznDH8QfLLnWl
b3GaFiBp8ZHIPf53dn6RyDPjmXsAobWD4GfF/YInDnZrvmdcqTuXq431SErt
82w8L5s6IuDSo5hPoGw5Enk909ZwlsWRugD+7pOjS3IzBl2g5SBtmNM2yn3x
SuQcF28/rRYUtoP2m5wLsfI6vnVFM8tJYTaZzvbE0I9wemyA/GqK7TwSTAYn
sf8x1mDMY9uZsBvJNfy7auhUQuga6/BjHH4gExfJP15455Ci3IDyvxTb2mZ2
V0+P/ySfAA4GKo3hX85GNHKY6tSYEUhP65mazZnQN9325iBvKhDNx/4vKUxO
breIkx07Ip16yT7odp1a36p3kH7ZlCRJFn8Rj5ejk/cz4g3TPkel8/pAIN9J
ch0+w0bvSepTO3WuDwkjep9fyieDCA0AtaCNAwzyNSBKB4XtHl302+CeAgYy
Xl539lbivK+bfpSMAuBdw48mvAkkAjWmR+HoxVkGFC2/4TofmdX5nB5bC6DM
tMlJjeZBdnibcVvr9z27fFQp+RfLPdLlfi6D3BvKwxyTmgCK911WPxtWr1wg
bNugW1ZSEnbnLwWzmtendv7VOErIpGcHh8oiO120ZdBOC3AdD0m3BVmHq3xx
NwwXZ4SmWo3t+oyx0774rLkua9Lovt65djWUz7K0Dodqt+U+/uUqKGIdrhlz
yA4Fl9sa3fQt5aE2zLVKClpuD9raSPCuaDJkwBc1NdJOZ6VIIYKUgqae6neH
ffxvR1fmvchm6Y2b34qIGHqADhAWxV7xnphWcqo8gnyumXN+LuP034DD0jvC
Xw+tFaeze2VbrmKX+beIb7+IXnPsEvgeLuMl0DgY9gpd0JQ+ErVlDbZnA8fq
x08ew26C3THSbZpQtGYsJQ5tr6s6X5rzx5sfgDRisq3V0o20p/bEpM4UE+wk
TwVs9WtN9RxfwKO2sJkDZ3mjDLA6/ROZJbmwfCTYetS5TT9Tt09aPlISXNzd
Xg7bdoaYv5opxcZAYC2ZOMxqMCwi4PA1yCzJFRs6e3gU6xoIjQOH6FREeeG9
nRwrUMtX8QXWuXIQZHKYAQCu/4ILR9Owse4U79+foFZob1UUqRC07RhcCs+f
U8OcGpVXyipnepKds4DJFLx/i+9Yb/+90VEu+KZrw5U+v23MwzPwv9LnVLnK
lq3nnlfD+blxvoDZ8jz33I9950TBKZ9siuYNbOsNgc/gRV4WvcJZrappy4aw
GrrpoZcUdch/4zzCRMOZu2gvzG+/KFUHfpK3Fz0LfVxvAd5nc2459Kf9TwQr
7KkVBGehEJHmYOHBrMgNTMMgAce2m8FbpDw2R4rZ9OKaM516RvilWsMLg0AQ
FvGKakqfEdOwRAyhvMAAiUnlxtaohJxdQkEPZSHg5Hiy6/6q88SCJ7LeTw2C
Y/InBussAMgP1en/FM3pm2PvAXZ9H5cdVDyi2E8NJ6y3PsTSqy61VGGYgpDL
PgCiSo5unlwgoVMTtR/3vdjFtcCADejBtBzR4OAE7DormxGoxXJ1/FjNqFrB
UDsSX2SVi9IQ1wYSV3rwWiXzAZ0XAo/8oQMfnuXlvVohJPK59N3LOHW/Rsvx
iBqfJm8zQoxVeqJHQqWPhONyxqFtG1DEnUhj+0j3IF/GfDQ6/nyUmwCFdOYR
1KoIU45RoaDktgNCsWECbrdZLGDHYWJKe06qBy8pSncAPAZhGGv0WwCuFT+Y
l92kODnhbdXcagRStVPUFdVMRJfGw3LzLXJeNgAxuC0T0nYHqO/sjRsBf/ZC
kruoXWIcRq6i+QgxN5hM0tG6ydPdE5Vfat27V59IByinRkV4W7CXJA8MofgF
V/y4rKoEd3adBKsgA5O89g1oDPfEOQba/eCIHqAFsHGxRbM5oRMqhjOaJHHc
6qe4DNNzsCJgAX7s0Lh75mo7yMP7RrilPKd+HNvDFw/s/pPkn+Eiivi34IXG
mn5sBoBtO7smJ12GJ6fJSQdAWnhkQI2xqcCyrX82mkwckZru/20AwkbTewi5
RP5UPCmGW3ELZzvud4J5P1no7cjZkk8xa+6iKGY7P9dfMgGXGqS88gpJllK5
DBNBD4/tl6lhiY4jCq+stByEWIx+DQhJoSXU1un2f+p/tAEQTBqCYgbaNHV0
AlM//jH0uigVGOwToweHjYQDEX3ey1MWnhsuUoU+THBy+SR3dIhcrFfZORdz
CqJwh7/Fix6P/BHodsm0vAPLFK6h4mS8//8hG8CyDK7URURs94l9Ei1FfXon
2nj0UIohuvCJre95B74XdQzkJtv4CXgOAYoED2hFlLUBokT5MtCrz4+fn+ao
SpScH+ewQq8tnEPs1Q/IlQOxKlOZd0RD1K2vHMqAwB3gkIP7f0FlCNFUm9km
/k2pE7ai4t/6dmY1kRZueWzUG540woiydqoTHSBeNk57bXqVpavhcrxigZVu
jzqrPH2aDKKwSHjrvzaJxpspitraOpWWtHr1/xXARmcSsLnJrOMrG0bk5U5s
V8rGzdkvf/5eK0vmpoYvYQ6Srd+R5KMBYpsELTP67DXuhL4Oyf2L5Bt/bIqS
0qfy8jRL1P2LhDCHJZalBDijn+alt4tHY8TeVIGVbVCY7WqIBvCM/ild1w7d
v4sxf05bhlkkiNXdAcHWApAHbO4pr/DiaolJzMJ9gqGTuVgfneFJ1hbza/2G
iKJ8HIg/SuSpC1d4xN9I6OCvuC/oX+coyp2gCds2UHirAutX2aY6fkO9WmoE
JjEUSHPDGNbOUcQYnrPQuIN/L0J7GaJ2pqiKedK/XqXmSnXm/qQO0ZY3rIfk
Xk5W/rBOBn7S6aGxeaT1pBJnxgBQOlthRECqoakW07JcaVPQFDBEiaGjxXkO
ElxeWyi9G623IyCVDinx4wIh0R0AVlA6zY9l7iTpunNPTSJR+yOWh7gi87wR
Evdzm07S70eiyZr6KgbieOE3rCeqI9GnHC6a+xWUPOqkqDGtlGMSF4UCx/9l
IBaxopXc2Lvfow/zeWXzDKMhLGqgP0u7jfySD91iFHovD0C8VaV/MUZwnQ1t
mB2QHdbSwBd7GfjYGyuaL1XrPL54JGDVNaNYZjayXQNwSPtk1H6MdjLr/2tj
XEtpjv3kP3DYCRoaBo5eSyarl5YPoj2fk1RiGsW8t0fFtf38MptJE2K4yq4N
g/xxsNEbigx/7KbIaur5NZs0gnpEGoCgfoYtbBEtKogt99jLx/QvafxxPqKj
OzfiP6Xh5JCC4EZDqQUElttBwKFVv4W+aOMYhvNWez4FW9hpJF8CUjkk4A7G
9COx7kM2ThKAJNSa9FlgOK9cbF1/3VXrjshjw8j+7pY0MNt3ppOAyzEMONvP
GycaOpvzvsJsfpoD1/qCFOKL81V0N4we7KmNSK8RFkPo8FXomeXSUKpE7H2o
jcArApu6vxPRN3dCpQaL/j8zrOFnWNywIeZRmJjm9x6nKLvSyNwGqLeLb4sD
rNwyITCUFcLN/eB1kWpwzXkNxD/l4Te7ozEKocXE8oDutvmsO+Q6uXH2BnrT
LbiIcYtI+MoYmIqm37pm0az9M5jwY7FjkcFNX9yPKEOcfa/970cl7Sm3yPsz
VWhVMXjzoVjAYoHmXe5Ug5Nk8cJ/+6HlBn6ahRBrKBh8Qrf3yhjiYznO+R6R
CFKxyiYT4wXWnC8JL8jDGrC4fRxNfBCBbHKkl46ORsQHstdUmtwj0EvgAyn7
zdXpoFygXd7eVGdYsowbZANVPMSXcOu7d9q7a9cI7jF/LXFc2PnvfkLOPkuh
cm/qb2ffzHQ8AZoIgATuLXk2YAhfuxLWCPiRjQhjci+hJas/9mDCdtaBW5RQ
tcWLR1bix5U6lMhgpUn+C27oW40jAWDriICxgKKWBDWAWbYjZmh+niFvnj6X
/wI0ieKdH7xtLltzKufIofIK/rgKsu+RGVQwIp2s18gpNd2MZyfTHAL6MEhK
0QPyojrveikPuX/h/3sYSlICqWOIOKQ4Zrl5i6Sm8QmNGq1i4/Ef9aJxXY5o
StD2XMiwxODgMaZm91PA5kyp5C4ZUgHxiTLMPHET6V/YnUu7fZ5ztTiXp+2w
LERzvJ+LzyUKp1ZOGh9yJpMzw6M1+i9/mf+MvpHxociGJkFbJMahCr30mohG
yBkn0rP9z0XxjnehKurJytrHccLY+BO+fHjQWnhcOy7buXvf28UdzTA4DjpL
UFdsLryLAqd3TXcF+3Ryed+ZFj684SpNJlyP2WrCFPqexgVuuSf4xKSDjPki
AjaN5yisj2cb6+BCDWS39PCbQ7W+K2HfFw6G87Hsj9yBrfd9cIYzoWImXxqv
+GOMT7HNrPISLMD1djcOVZ/95B8LEPTTSJzIbJAbC5LEXM+v1/vyRpNYIhIS
vWCusIjNNdfAGmEO8lnnH7SFZXPVSZa1THXiMtfDfByawxlRyhecP1iUQfNo
leorxswVpKhDJmqX9PmdRKFbzvpgAWPrrlMatPQcU9fMG52qxLReql4ImdSk
+MoVn+d0Q2wcZbR6yaia2iDWNau3lJg2fe+GOg9ZlECbdG/IzjbyLYZr6OTe
4Sd7JdcvrWIO8N9NWDG+xSs9v+UnpvBHwbpv8fUnobkT1i94wMqCQSUNrqEr
CgzAPqva45r+29d60GsJs72jTfQw1T1/5UYauMm/4+mmupWSojpZFUW1ZLqz
s+fjgQIDxy/QI7sGrGLdpc4bVeL93Sn1luypNjiiW0m5KzT7//n5ILtLbcDw
Um1pMgGSqLKosBne1ArRkdV1z+pBnd1o3oifCKUmQlX4Q2vMrX39YElZZlAa
DIVvyA8Wf9UoxuVtfS48gNKP54aYPTBoOCpHIluCjarowpFe4IRnB6cQR9EQ
4ufBOQDaNOXuZrpEmitvNaRvaDs5geBndfwO1cS79/3GhaAW1ndI+jUTm/2/
p5xOZIIH1HcxcY2Yd006fAjRmC8LgPG87tMLStVxIhJ4D/hrN5B9xOAI6FcT
BOl280MlMAeYnf0i4MrimSEJMStFG2f4hVm4+px05qPWt6y7qAQ/MJxA6maq
Hk9yjLXj6ZekKQ34SXFezvzcTNd7ZigsFhZAWHmHzj2FE3RlabunE46pZZgF
my7rTyl5rnCnsteikG0Tkp6ZMIUd3J9KbprL5+PHnZ0qS73zJFPg/N+yhcvS
XVXCb+x5CIACl+F9BM/E1kNPzSqBvZYNldPMtlN/NGd+49qVKck3MinD2Lmy
PQqPc+M/7mD0aMe76g/3Mt1h8siMXhHvxd6IqcHT/fPRB0l1a0Nz0X9Ty/Um
v7tTdZZTAdm4ne8YMzFGnMm9Uju/wlGEMcfvzHhc+jLbga6XkFrPAbXEpDOw
zrz5+hqHj7X/8VyVmD+VaQPJVjQtHJnFD9h/ThVw9ui17RfUwnQ7eFP1SB1B
F1fhJB17Ekz990UTJTsRVA1O023KtECfLRrS3tdMdZU926RUN4WAGcEoUbh2
SufTLXF/ifNCAUJSb7ZEUzQKVPZLTN91WduZ3UPmh7UO7CDD5a2LNWoWtoZk
lWcJCZJ1B5LAnWr1K2qk5dtpnbXIuQp+HLLp7szdh9cUDZVqZ3WsdSIWimW0
zz/S0KSc16/QxHs3sX7A5b1gN2hQhKZRmSQX6SQoLAAvmzqWM2Narmivvx/6
fLs5/LXutfmBGGK+X7rnf3Oirv7Gfg2Ef1cUmIx/qrRvvlXut2G1nLBkTOxZ
TpJqDAyz5JT17AckKko3WVpU4GYvaJVcV/gHZM/t+B+3m0CC6jwrJOsy45xw
r6YOjSeaYuEAXc2tONshXQ1K43yIsZ+tNBpjO3hTyFfwGQ0cQ4U6l8AJ470e
i4C5xEvXpG07j7We+E1ENACufqlPwH9HvXSfMqwpm1qBB7MQCyTMDkUnkkxk
e9VkpNi5AjjwnETgX4CKxkw0ZveTCn8TTjmnBGm5alX/ikMJA9MPEYg6kFMA
ccTCWw1hrBUknACVCfG1EIjd4FeokijIjclH5Szz+JHtpzfFnC7FMToVNHWZ
l9JIg3C0PAYsLSt08TRvjg5lnYsVsYagUGIlb7WXInIi2oABlqGJDVXH/Ac0
do+a4CRB53Lz7BH+3tKHQMpefdt/GrhGZZQEU0XsVbpmbDx9O5+hzOesZEhK
CWS5H5oBctuyFGn0H9CskGzv/0/8L0uwOuxXDhhz9Vgx+p2qsr7ilDBzwKIU
GAdjfWN44r6N5rMD0hb5xlragNnVRndAXL6Jm+voTLAm7yLAMWcJEcLEhKho
7l5bTKkG1kNeA3WA8/gR6jCuKJSLse5xLQ1qwW4WQdJHkJz++Ore5gpD+EbL
jGZ6GpApCgwupUpxzk0Q0kzDrwO5L8jPHrYOwEHhkV7Z0VbDRVnRvdHaMP/g
ZQ8bzPKB3omSsB42x5cmtAhPuND1Jw3xiYuVj7W6Ch37PI7JuelAL3GTHnJ3
wJI1abKi9mdJikfWSL+8g5r3CH88jKcjILPx9ZE3mEPYsBdH8MKv0PJwTxBt
A/1Y2hSnIdfnx1vioNT9J0Ewk8ULX0qlph+5G2P7KLN8JvcLkVYxAt1qci5K
g+iS7ZKjfHG4cjLyvY8gFnTcVtVYjXOxgiFkx28lYbodN6EbrSr+y6ypY/AJ
BMJFCgDtUw2YZ0ZJTK6bTnt3MOEh7gRHCXQnxlWRskFAdxKy/QU6yCcKNKHC
SNmYeHedvfFHSohb0Fd0YmOyy5FrLprwkEDSa/wJhZyKTB1VhOfdkcA9DMoO
cHujeNGi8lw/KdqKMzu5fBltQAofmG9wtX5bp1eJ0L8BTJJqF1EdSYbCIShF
BXoQ4JM2T7p8NubQ+LHX3LeyWAcu2pNM/v4VbAZvlXffZJqBwriz32fbhowY
gC5pR0FDIS9qKzGwREZKYIGNTZh2PBEJA9W7FuUKFP2jdbKCT7DybwyJsEKq
igCAY9U3X2plbaf7jIrGfkzvU4Cu6HfVMySUSkaelUN03R0rXwyY8ih4/xKj
4X2r8iI5VAqO82ib/BdZi6xulpX+lYrItdAGOiaphUIHY3cdue/FTuG8gP26
2bqvd1fXxjIHMwL2GSTUaMNyHdSNuk/p7FuSWLttYepGwGCr4lIMq4eZmcqv
yTV8DfmZSRca1n/l1XGDSn8Icv0Oa68tdlbKCEBfj+QIAYSchUVhpMZExklD
WIk1pl+hfEvwLVENlqbl0Ik4Wc1V7s+6b2K0UWn1dTC9fOj3vj7jPQKz1P5J
peCsEBRW9pNIUOqFkfQr7KCvfw7fvxCkNGUqp+pvJ+zywJM2TqspiMgTJXSw
L9GPAE+asCm+xJf4bf5log/TqadtcRrETgDNITLoiN7gkrH8nOGCoHjW6Mp9
mO+tOIYs9fFz/q8ExtNcPy7g6OlFqv020d+Ro3THKdvYVdlF4OP1SEvHa/9/
GcpYkeE+MoBZ8PMjnG9qfzi/OM27qI4nWfhjs8xLKLRj04KMY5+TCH2Dfyxh
vsDJTQx4BRfwnwFRhUh8nJgih8qgKkiWtkIbEehhSpmMuGPgNl+U8Vb+ogT2
zVmlf4GfUqPnMscBqM/eSoAB/nEHg+mD/avuitI/50ZDNA6Vv4Eg+jz+6mUr
LsjstWYOprVwIzoq2luMb3vDx6q7ZvSETEtosNA033YGRFDptF2Klk1i9cLI
rUGpDqS4iHotKX18u9KMopt85grW9kACtVo6Cv54jzd7jI3Mp7iFs9JEsK40
/PZdY++BTMXuuvpKZT/cvlcqriq3NorM7fwb/qZUj5x6owX4KrDJ1NP1Igk+
r/1G5jGpNcl9liOqO/tncA41B5Byaxnwx74OBXR8pEFLmGmTgoYtIOVlHxuH
vAgFR9hiNJ2TsxNG3I5TaaV0et/kr+ntR584LOheZFtjoeGv2rb4gJFiquOH
QHe0StsmnmzwRlZ9ey8blnAiomncgmu6i+qrQUbRoWJjfQm8dVCz7J2BfNTH
iHEsIIKSlWhw7Y3iiQlM+W5tiFAo/ZCJZBcIiYMZHGhHzXKImbP3J4PrkMol
mkoS3i/OYAeh4Lg1IhFcFfN7fLdINSQR3t1YFepksqqUrDYbJBg8bcb6XrV6
qwOj82kfBN2qPxLRLimXlsr7qD3AXlMqUalC7y+BMd/fIGiYiKxEI7Y8LRj6
joiggJmNlGPIb4+5JU06ia5HW6N1lgMylDBQeLH5D8Y6yURi/yv3P92p1vjN
voNv1vyU6Hm0qfLNe0ZreS+Pbbq92988juz9qZbZPMLHrhuznL47qJ+gZcY1
9LwAm2v0xTyv3IbIl5D0856OtzuxvyfkS6BfkFzhrYo0ihPa0qR4kk3wRzHC
2RpqJDGddGozYIcvZ04K4fajnrBuWqoxlTVfMHPTHJjiun5WXzVcCRDnX30e
WMri5AmR6lREu0Zny8lKkTOmNh0yOOPdt+Tbnl1qo69mNw1/KLZOGy9sCo7R
kQip/9u7y0VUErsD3XuJp4d1H33jd1FGMnBdqJYZx7btTbiUptmvjkh+qeoZ
D0h0RZNSfa7j42V8EPES6xaGZkSsw7pAWzFLMH1/BFid7pfCAuktGdAjACEk
xDjxa4QGwdm/AfIMYSHRkBfHSQoCWsGAFTRgLI2bzGIB9pj9JcSzkq5MCbE/
SA/C39NgaZfvC3MuX2kFiqYj1o3uHRpiJR5BvAjefAysVbvRaiUiNNt+KLxe
ZdFiwRXMkgM8lI0uJ50/d93sDFUo+EMhd/wCJLcDw7AJIPZD27fNL34USdpm
+Uwy05miaEd1/aXg1x4oD2SlMQElL3ZqiXDwSrbDIUmbYTSfbZCPt5w2Mt/3
wAnOHgBYmlUBawt8sgOEydahQHi/iao1C7hnlqqiz82w1VVKuo7/5S0gmJoq
uqXtg9SnIJ3U1GNBHO7C5dD26NC8upHo93DWNmhWrY9cxUNLqg3mK5kqmZqc
dQ1goorMT7xD3PRFkDKGNAfqIi6xTgkJIe7n6hoX0833UOGok6dw/nMrDL9u
xsuJPAZmm28KXWY+ZmLIedSX7dfNTvyf+k5Xdk6oKgdq4HfoOCcprhGpBbPi
CITBWntMkzOHH6iffZ2fmNpX9RN5PNW9x7g9XE6ad9HCniWcbrKpIS3/5qsJ
EyZYWgAyPJdR9EmU8GQlApirJ+JfZBc8ui/LDXkb7KbVD0Xfcgg4EQOfg8dU
XkHbLDacYCzx/3dugYFGn61o8qE58LmN5qM7ISIJDBNdpFpjruXR82OKvtQ0
q6H0iZjZf6S9nqEiiAL0j6mq0OwfAw/zCMSSO8kIOBpi8nemseyPQw8Q4jni
wgj8Tk9YHeGAgKY7Bt80IM1NUUtD+Nr26Wb8eTYAbFMRFI8nNm53ddUH6G98
NWPdnaeu7tezBRWruS31PGIxmvsdCGbdrJrGcE/zeJdh00khs+jU2VjNmzTv
6B+t8RCBOj6fvUsw0NcdBPCseOH6++l5f7zmMRf5oZZS58zyXUkPIRGbsdSo
D+YzsLF4wjgz2cPErDf83A725SHVXMU73eF+XtxZG6u57xOjbfv1vDj6569l
u1oqHDlOgmJuHBR/tR0GDEcW5e9N/oI/MMmJjpplcilfa9SYPTtqPh5NSRtb
key8TEMyzav2+8fHdfsi1/Xr3UbsHHNMj54BgQmRf1fo+/Sl+fSaV3DFLNKf
RMXB8+xxOirQhTORzDM2UnViTym9wjsL4saYgN9Zgv9NeVhott1DKxcp3cjZ
bRIFtuMd7iik4+g1S8L7jwaZyEiOYfVCNI/VmpX9vhsvkDUFAMZXGs6KNIp5
PY4h0SFwZPj7oeER9gvyLz4AXo/KbOPa1O/g+cND4XYp2AlFMgXFpFsFUbMX
eKySDdoLNHOyoffupu8R9R3OD7g3/6pnajxJqziQj1urq4Wx4Ayw1Ij7QnxP
CEKMEt2xv6ny8ObpxLVqDNmkRIZwmJnSmFIYxYTCK8hy/sTSRmU2D+d1vJIS
pUpDgYLWDeGfPhVvkYar9BM+Fi6ls3UXoZv3qH4s2hnzQ31TEzdCwk1N03tp
PFNDundo+EFrSGU0F/FXtVGyaERCvZSef6eGNg2t06KPAth5s7DoKe1GcIeu
0KPSpr2XroMFkVYYY5XKvsOW0rSzgBdhF/MkEIxsApQ8twB8mMIQbX3YX0bL
RBngkGheF54V4PCsIPLZ8Sz0GE1rrosZNBsTN9TuZ6bvulaLE44+Xl/UzR8n
ajQcR1ajRKx6DMBVSvdQjhanx+EB83iZ9Nvk0bNIpYZOGeHhcK3KPq7CDi/o
YN1ze0JkHI2crTtpFfe1P01BG0glyFMe6bxvhh3l4b4L+Lq9KUIO0+bENwXV
J6MuOgL4zI83TBXRn6pUp1O4RPahQ615ahcndbwdCd/pNILvCpORQ0DfxxH8
TElWv3A/8DRJVNCx7Y+lyokBkVxuA1Llx25vw6p7t/X8w2a8yrw1xXA/FnAa
R4aFvoSJ3SF6llgsTjQ5t7lzORRMzSfkwrRjdxx3DHvZmlKyUNiX0lkuk36v
alFvUdE8qu9JiXST8m/jKXid9AHBEEvZrX/gbKlORVouLyVAjq8PHP6FvHAB
xCIUX0Ww9eNQHU6tCfkO7XkNOhhGUxG3wnbI0s6W9oxSQqRd+jtRIhB8QzzJ
Juc7OhJ1/Wb+Z1XM7QSKzVSS1ETDatBVafhQD+9ddYl/Y0ObKTImlyqlpo8h
Jh6YLA35uWOJzTLRHLOofpYd1pLVcnICyHBCQFiryf3WuEnND8OQ3Sy8RflT
ICH1izDMp6pYnjFCxLj0DMhCuR0q7FGck7iiVu3BbmDx2gl01bFv0MbapmNY
NZKhCX4lAjBswKLbb2rInR5isx6vsOOiVzv1Yu3DlrHxvjlCVEFdqMVrKazM
VfPS2fuyH/KJwtNT4mRDW3+hCf61LC8ciNtMApUBktqD4pvzoYZjCEVdTROn
T0rvKd17PNr5SsjO58P+SSocUM3brwxVTrny3QEZxFJlC84e25wQusgJxxTc
ktpLc4LxygRUTlIIAXjDbz9DuGjwOBuQV2tH67dp1WJ03ldoH4gWsmZxoR73
Pcmhhu1FkVoKMmXiGmtDfCCBWTapQz6DuBJg9itfkNdjhBkyZtyg127o/8wT
wzJwJGdNkwvlE2oJIClDgkwik1Fm/ZdSEYbs0dASYinXDeE4KCSYsiV80NU/
asu7ds/OYzsbeudnQkuoiBr38mKthGYP6ozQBoqS2KIkLQbceirFu5mi5ghP
PNMRJF0EfySBRtt+OzPCe/ilGWnT2NB18wsA2Fo+tcVm9C+17nklzm04mI08
TtLWMqECuIeMIX4x1ikjz1BFxUZoOwHPHzeOMrNSSjBwNvL42teV1Cdq6XtE
iIE7L2OJjnnmXa86XofkwKJDAYkvOk6CJdc/0fo57AB5wKhjid9eHa26wneR
dEK6jQZLT/pAUcrSs11MKYB5IsZ/RO+CBeULSlsoSuRYoS+th/E2Yz9591S7
cGtE34TvGpT9jof9PYGU9TxoZPtU6ghJWLdswGRXjhTOv+r80cfNbyEvQaX3
1odLpb7umJU9ktEyujnbJQM/23VNrPoh2DuYPO6fypdv13Ie1QuVbpyIVo9o
2A99A7YZXSrClpAWMZaPV5YGlSBYyfWjbvsxekCyHuwxb4qpA+Cye1U9f6Kn
GKk+Pm1u8zch0mZB+gnSZmLbBihC0EBFs2AxgnTr27TPOT2t89mmYtyFwyX1
6rAN7ksqD1G9ZfFJnheCi4RADXVzuXgLZUqh55aCd2epF7Audy0GveLbAc4M
qUP886Y8F/kUuPSBkTRSaikZTuMRl1mIMKVg+FR20Fp3w0ExDzqQFW2+5hhd
5EZ31zSnUlppMJthwbhfIobCZjf8+XRpclv/t5bXQ0w3Sx5gfQnMoxVfabYk
3fmi2w79Ni2oL+MY/YNHy/EGcCHUsybLcEPNJXu/beRJwPgPzxfEWu7w6o/e
sVmM3rJeNemqXOY1idUyPrhLfKBXpbK9o0nixI4peeTJBRf2CTqdeWMV8QPT
kjaxR6ga2xWTEQ2yfs8UbF0qfTyFkmwy7BxGRY5KzLimNQefmMUXJ72toPdE
/XIfDJgI/7YQgTK3yxoFUeTPrqUViNpNkQJOvyX+3LKxYZjuokLEWv0CWVgn
WOL/8GAzch6mgp1Lbn8/bFNCzdoeTeIlmnomExVRcL/6NV0Dtl+556UwF5nl
hZOhHXo9Okn4M4hVDPeu/CKGRACCCmcKonZcM/8V1CYqanENt0TQZR7y6Mmk
Hs5rQ+P3qKgfV03cij1gaa/dhUZtoyfKK3fxBZ7UvpLB3NARLkubUk1+JACL
RFdVsm1mIgNkgo95AIYydAk2SQA19kjXo9SZ4kP1jjzXEbBfddm4EVBRgFJ/
ymAaKr7kYdcvivCb9xmZLWbBLpKK+PqjiXrGh/tOTfX3riBFSzl1y4WfczpC
K0GYJGgrgctLl1H9IUJ+OwUT8hP9qFOtW/gA/rkkbmXARpyKRjl7MI3pOPHY
0Ag7h5Y2mwkK3BqfIkjAbNka2pjOjZs3sIoWns1vdelxCdFFgijWGDpsDdei
+mSCCSA6STenNB42OoWJ8bOid8IeUVJWEOX6j4khJsuWTCntdPCrqHYBKya0
Rf4AEFzMBpbH58As1oxwhxmoKiPcZeU2y0v5vFSAMMPfc3a5wGTwJI4QdxZF
7WDZnl09xZbSIyMk4baktkXNqRE4p7rzOap4HSEi3Yz7IE6PAIeNS78HA16k
ftVAf/jeSQQ5+7VaWYBRRCH9eXupWPWxiTZQMgLtLC2k2/axHVRN6LzoKly7
5sKztZDihZOqcqSEHT00TJkn/Rf/M5SZxrvhsogkFtnulc/qV+9ErUPhNfex
8u46r/sIRPC2Zet/UEfK6RsgJAgBiIOa5cz7rSSqnY91wLJtC5ZmDkyzhJAP
3WcYVILAh+2rY1blBJTQJye0Bx3CAnbelKSkKpEfvdnNEDfmyMtyP+Vj6Upe
P3QZVSOG/MIQ8v7t4gMowH+ZuVEx4dmygeQgWxexmuMyj9n0sIkK6TBQddGT
4PVAQ9PLiRXsesn+sDaYkt3cExya03srHR8CZHGI6uT9FycuE1fbRRHX+Y+8
JyDJZICj1pI/8wXnAq/pWdXiyIlJIjG0GZ1gt3BPMYcZuIfbSjBjeVCCGiLS
vpA+L3TayQXcAWM8TIHtkCvDersbTdi+j2ehnzqpSiB9iYgBJ1TsfHP5i5C9
fPW6Mp34CCsdxhrIeLDjHJOZ1uNYaY+fNSSswe3CXZpOFDrWQGvvuvCufOl7
ZYtYYbWFRrV3NV87zocYRcH582fELqcYIRaET8Z3PnNjCvq55TGrZNXTcU0d
88IgLLCgnOQ8/HVWTMTivepUEqCfK9R1hnCP/sCjgv7X3ydEseOkDQPBUGBc
UbYa/rkFCFQ5oqTv4Pstz+iDFwwWWB0OX4Y/LHYKzN/zu2ZvP4Agnn2w1GuV
2dd3TlZIRrQNsxgfRfZd7xShFS+4rLH8qAQWNNG2EeNllJeprboz2Oa5Iuue
SuO6oIY+7JouIg1RrVhFx2h1RWRh94tTcZ0W8TxmhlVQOmG/jDMruoqUI6lV
keER+oCHhbB1oy+8QbR0sWHp9wzt5H2WruDCkmqqLmlg+t+8pyAizrU2OdVU
5CnYShVZP8PeEl99UuCYCJhqGsD2Cosq//axCEusst7rSCnF0i2UllKlmJfY
LW56ZMIUV4aQK/kAYFabNGQogqVCs0LHoqUbEQtY4MsmeBJKH988aASo/8Xu
WbdO5/X1prlb78IfIH1X0ic4VtNIqVAFIRLsDVlLQJZNwWp6eTvA1Sqp2Utl
dix5spXCubzdFnXwqOXNLJqCaayY0kKRxkiDHp8fwbitxt1tjvqEWeW0VN8e
/ZQDjRdFovkn+uWIaCgeHwaKIuW64r7CgJFV7iA6ZAk5L53fTkFIV3tCgUhW
3sB0b84rBGtdFWqPa+ik6T18FyoS54FBstqO2r1khgwj78XC90Df84YpvcSA
tsxGcxZH3BpfDrOgiBB2N1L87oqPemKK0jD71gHIbr96gWEa0tnU7D+AjK82
zWAmjE9on6vaLNWVuqpOCfOa9z7A4CsLS9Fs475yjRT+vvroAaFQUvhPQRjw
mMWOmGEOOm2ejcDxUrgE/H+4QFInuknrtOqKiAQsdr9qZYU3pKQnj/kdFdhb
n7ceFHRaU5E8EVIL+LYl57ecv0ClpM8cQRBlGKx0mHFUBLxaiGkUaEU/RkUx
uHOcWdwBPbE+8gy9IGW/kgpLRPqzJFJzNAnHmg++M4UcZ2UxxgwXKnyWgVw6
fbCcTBcKwpvljFu3PQjvQdWIWrxVpr/xWw9mXddTL+rVeaiJGCDd5KkkcAiG
HkOMEwyarnBQz6KoWxWYO9kMgJ72uj1uJLOBscLqPBQ+gBVSFdNQl+Fjh77t
EE/Ft6/wurBRxrGbc0d6sW07qsf0L6CrilGaqNkilkGj9RPu08RfAME65mYg
L7vl9f2vS9xmHGxNgEF5Qu2tHw52fW3MdPH/oaVDnOOGY5S2cryQ5Cjc+mQe
UPZr3BO46URXgOeVEsiA229u0/8WttnLTEHWTWGiq4tHoEhldASyLMzgigmI
zjiO617jVJla43WLmJrsm6sdGdVuQzZqqJEDUuGJD02aPvGbKHZZvYR4u8fS
T6X+Lq2korW1hVx0BGfRnQTW1wIohMLayNYjMB73zNC2+leapXncixCUYosz
MhAouAHxzhQiey1GhxEdZbTzcIP3M+76wPs076AAlwppAElNM0t65tmDuBUK
mN0Cf4kEWxUylx8MqRxW2AXq7aRqp6shxgJ2Jo5sIfi25prhGU8xQ+Ew18ow
/39caKUpdXz/ftAnAqJGkHzGYV22wKFsFILFJXIr5msMVlIv3T6jObDGHRds
Jv65rTIAjg53WD2gY911aX18XyuyP4Mxg9x1TDFk/ucWlfqlSXK3LatowDEd
KjA7qLUjaAa6kPcjU9y2bLkNVMUS8LSrfM1hqJOes8C4VGxza4kxRxbGvblt
DEihHFUcwHCsgpLKgzciiimeFeiHGXCn055bdWqW2VOcLo9BQVt5wIDfjUmu
zFW+cY9RdF3XOz1i1YSLzW+3Ay1fchqzHC3X98awIYUPn8QZwToH/a3C/QrP
jL5dAygr5vmgsP6/93ojNelqPwLE+/emhYzAMEJRcdZTYA6qNcAnoYXr2x/1
YySsd1ZGG3WDcVQGqU6oGjt7adID71v4QFZLyVQS3T2h9qFK/sra6EB2OO7t
ZekFLpH6WLcRY/vvx4NlaB5InoWx4F7rwPql1kPKBgatpk5Wj8SsepqThtf/
dqD6R68PvIdkaGzhgV5enhTzgdiuBAraeQJ+s6FxE5/2LxzpKEEVNszmiPk+
qL1Znq6AvFKCEJOxufmpIjPfKMNrmIzXPJ0w/EsXx9gGOIqTK4n9bDc99gEL
8SEfYlIea1N4wMRpM8kqmBjSwYs7BtQLiui8qZ8DXVKvfUCOiN4fE42uTSVe
C+iloZpEGjT6lj5ss6nLdG9tYmHN4w5cMUJJwD8DxZuRPgMVIypHpjMBt6mj
Tagd+RgNIuNujDhEIIfXvsPrAtmnYdf2Bk6Sbj1M+y4nV8C5Njoee0m8FN/l
M1JWiyfObC4sGgK3Hj2d2odXw4ytyB+Lf8K9FQusr8VBO6cOV5dQD+cVGGPV
YqoOGeBrqpjvNDgdjFo2Sr/IPM5/Q/3mqs8//xZ+tfLhVZiaBVXKMKevU1XR
P637ICjQPa50ih7Xi7C8JddODdV+Sw1tEKXNcPg7FY2uC3U/uLogtCCdqXWJ
G+uOsFJiYtP7ptkrrf7Czpp3cP6AJsyz/T25NXBMIVQlC+LnRfpd0+Dmt6Pb
z3KSuO7TbaZ4hkZtmKzjIErkz+H05bFmGwOo9bLgeU/Vs4q5qObZB5hchSxR
LZbZECNLYqWHbjakfRoYtoaMPzozLH6c2ma3esUkCuM505ZYZw69Ji/adJkQ
g74mOYbOJ/zJ1ocFjT7ELPlXUGE5AjbXOQhQSiLdfmtQLis8itrw9Hf5mIWJ
bhlzBM67s7Ep3aGNj+NB/IUhNkWnvC2D5nLUzS5frDysQlBU/1wVr9TTfgAO
5d/qP8wsnm2GxEFgqEBEQ8ysT6AaHQmWqK48NWIZVd9CFQ3qcvFxSnjl12x8
SWww2ffrva7OvxkTXFlSP3Hm7RfmTSP/EII8ClXFg4igpDo/dC2n91CmNnKB
Nh/cCgJRf8zDeHS4zfJ+WoFpRf77lOsMpwQdbDSl7E53wBwHlXV4bbe9Xxlz
rNvtjWfzWU+xlASjFiXERBzuBRApUFzvk2LI+JpVgtaecGCLGYBFrR+wWv3v
drCm+XDrGT6xAuLrQF2gdgkZteh2rMu6JtA7OXuq9JC2obrY2xipfQvj/PRs
CIVCznqA/D0PTCxFwNHx6riZy90VM0WlKHcazK4TiiIjOCjpPa8WD1/VknTm
uaZw6qIxiABC1S3zzLNS0anVxgdpEZTPMZwEqI8vAa9T9K5g9K8MuDsaSodg
Elb0/WN8hDCZzklTT1othq2HgBqLKKF52mgUVx1NsEyb6599CDaYoERqQKSt
PmECveUEiyqSkc3w0Qlb0PqM9f8XvzmUqWFqdvUNjMsWVVYSWztX4hYA+tqT
CYCnx5cDEg+z7Kx/8307NZdtFIeBWRE21ysvZMvHr40l/aAoTGk4bD7uRSdJ
r1adiACr8BZjoIZJFXiQ0ioIhdCBF+3KvdOCuT/N0nvECEkZ+OVBjk/vR4+I
1vPQe2tVj4dkokYF2D/bBxFDhNZqMZ3e4TiuPju4CpBxzGs8rIJG1S3L/9NC
MqvztP8RLPnyQin9rNuMJ2VQtctrSrTrdmPXijrHXHWtwAr7bsHXHw71P80t
tW2byGQvr4a/kca2JmNrAoynpuMH8M1D8vYcWu9xqxs6XCi4o16WUwk/ljPr
SO/VM9E7CSvf8a0NTEi8csHR5bGHvuHhMFvxAOV7l3GpHxBg0CXFq575yxu5
fM5EXmGU5/6BoRdNu0ttFDYEN2sV+LtgbfJku6Fkizb2lfDP8yAcwhU1ZL53
bzIhi70ozQcS5Dm/67OtPPR/p/UWX/rTOzUnyjk8pR6agfbiSIaYR6pxODHA
8Wtb9y/gbNoIbkgeNQ6eAlacTCbULRZPsgfdLpwRsO1gbE8NLGxIREe6MJyq
3hy0lSvc1AXmKZUkj0GrlxhInxfJPr6/aV6rMgND8ZS1zfFJuzOM6WxRF8lU
99lnVswQ0lQ1J1UdES2SCUROSWhdw/fz3UeUA0S5vgVH9Iqft0pPCwqnjW6M
cUaGYtMtFelURBmOEQOCxcgNvyCJ1VusjbdgoMnp7X99BTsNB0NnGmuu9d8R
HxswJaMGNa6xM5+LVbk/BOgUN5ADKxMYYNva11I5gxURe5pJ1eFewf9x8kQU
6MWfU/4dRz3fv59E2jppgmWOSyQuEIPcJXQjQOwEx0ATXqUaFbefk29B0d7I
FKoMm94IqNj9++lN1mx8tNcJZfXiFmlD8A2gizjv0a1rtSPWm3PyY2eEaos6
aGscEjLCWnHWR62MD7L0nvSQwF1DfZ2XA+Wzi9Hhu0orE5gh93dh7+zqm8wW
U0r6lmqMqdIumpQmQS3F9O1rpq/FyleiN6kaSEySkZcBgKp0RiH6WzDJdfSp
UouKLxUE0VIRYLh14L3uWAekJ+eWYF7s7gWwuoCSKOHKDOnVlSX2/c46uYUy
X6j+amGrq4uwNL2zzwJRyv6J92PoGa6hSSWkEAHY2A1jwppXTcB6+DmeAAy9
aIDOmqJb5zydUCaGywhMG+Z/2pSpyaBlUw1ccTPVVjsy/Z+TXxwPt902MQmw
VLSRcv9JzXwKGp2Cr9wIF5LHtMwE89tyG7YoKWcgUf9uNSjaRisTuvSQsYhe
p6ipTQ7aI/n7mt4TgeWM+lmd0taDUOGrKl9wBIVdusGXhxVTTPyO3EnMCYx1
X+6odVhFjOes6IZk9IUxYfzSyj6/YRKZLapBTsL/GydSKy/NWCdACrFHZPzb
Eb5VJDpXHis1fiHoolgJoSMbqVpXBEWE9fQvETXBuC1uBfORwCaEVqA8e/t8
sNJ1r2ryobPRNdukhDWjdHJm1I58cbCCFOb62zaCIPLkV8w4QlSPVaroq0gE
AOBju+NmYBus3vHadSG0vva+A10vUmFF37TrhF5zUPt0ggbt5aD+4ak8ox6s
Lx7ghwXzBOKm0l9tGdMY/zqAf5HHC5wQPqgpuCDgf6Sp6qK/9hubnJaZAUHI
qwWRiQjY3OTprL4tvEFZHAfdeo36E0gESZDiclWKuyaXL3yEzX1xU7gGKLPC
NtKr/AtzUJjhsPzYdUfvDFsBB7ia3W9HTTpkh3OOEdbRQXo0kqVba9xQMPuJ
xbHv4bt7NvJxMCoaVZyWeRgP798azn1hSF71Kz3uEnqpYglIfwXQDpx03Bm7
kFxrokLdx4RENXmao2JExgUuyElMvl+id/y2GYEyap2WG0xtJ7sX5uvZxvPc
ibdvYy8/xqpB6i7aS53vcSd+VN1CNKgvC4O7YyyFnOwwnZYPsXQ4NuvggD3C
mfOAm8RYEQdL5UID808Tr7F7uqyJg4t73KTQFGGQPb2gdwbfQzmsgU2F6Ivd
X291YLYZF1P3mw2jh2trPTBsjXWYa5SwQGs6Gei+FGSVG/dHr4lIENRf/BJ0
VSNTrA+Y8lT2xwm6qMONatIS8h2i0/8dNoGAhqyOA66xHJ2pHveiAEqP3Sr1
Zm5cNJ5zjhMn+iCSximPYR+8LI01U23VLjrPPHnQ3OI8D4erByZv+kSBaVj2
mVYPr9SX0WTH+msBDO9aqhUAYWDBQnNoutHdjuB9hAJfp2a5ZyL/P9VDKPVK
OiulE+IiPGxB6ZzQaqNMzfahTdWO+fFPrSQLhWdaE8ixxiu+oYGB45LR+O2d
OewA6NDmThc4f1DTHXd5NGvFa21DJcM8m1cj0vRsCbL5I7lljtXpNdGfsdHo
hgwjDy6xVB14wk02uWoQ4j52ePG4hwfcHqk51cGTzYARFADGpYdkOOMnAqrw
2LkzxLoGK4XpBwjvQYCCUKvhQI4EqgULazy4AsRhvBrkvK3lydIbuuz7ImOz
MsEEZ1rTgXbUVV8HCHXw7RPGtVBL974oC1onFMaZMiS1r4QzsCaOHuLHxgHJ
dq2G5GX0EpcxuQjMMvg4J8FUJjUQtNBKKwgVxlRPN/tr95ivs2s2eNpwBdr9
PCs79YYC0hymAluJ3K2n6gKGj8RoZ6WH6Ns+/h5U33BGODP8QtkMAYkGkmbX
CsmCYdy4e2CNp1hzen0UrsdMs7a53VNNnFDpHumWmYh0p9X3bjPruc5kCtoX
Uo8pd1fkTbebw23R+oSIvh/NVc2x2go+jSymtZAA5Z/iMdJfv3RmQGvotcJq
AQTNRButQW1RRd9kFBxppsVbmv2LcJJsNj51EJg/tHckJUxNm6MBxqJlwtqF
7T5MURgZPNK64iduYGEvjJL/DCmz/2X+KktaKjVajL8Y2c8PskNIfMew0MdN
KqlktMz2vW+SozAFPUJMLsbDqozUwmONvt9KQxrSlnDYofhlQYsQB88bD0oY
GZei5E5BhfQVM94KxJ70pKQwTGu6jgXPnXLe+jVo5VUpR4pBLj3ujE2UooEE
jxklhIwukyRZX0AFw8XXzDKtvVBKBYDLEoyjiKwPpQXa745eRJ3XMHt/qUHP
aOnqyVmOWPRw1xtzJz3yQSEAVod5lGKDpBKecXKRqOCOPmlQtXZwvkdrJL4z
Fx5XZHcNrcse1N7V/bTye8YC8fga1vIPKgwQ3PnIzD/mnn6VCKW+3DyLNgwK
eBGqnt3QDf8zzx3sHjnUOmzzNzxzpANP5YNLvmzh6Aa37DL8sHH8B7qS4Ufq
sWMlE1di+ZDAp9X1dC+Wn7aQfiv8yyosjgVSvjMrqZQwe0AmOHIuiMAJazMG
sTfYEhdbSfSJjX+lqWBuCVGMVm6MzR/GWzpPWA4EFyZK+Gw/7pVjlLgL3lbv
d4gBAB86/ynuhnwcABuhfQYIP17+MJR3OD/zLm18O6gHEDnBhw0zRm9j4j8Q
2sEwuzVClZv0qf6TrIRcaC+crM3yhErOiwkhqAHUJsku5/4kjvFFWcAU9GpT
Xqmf+uzP/Qs8UpICeCtHmhbWE1uCR7lBvxqHBXRrqsRiy2eLSl9Pm1F1F9hD
77w16kDnOjRItOHqcm8Ro2VE50a7T7JcpHTOExD9H4l7vBgPvx21QHHkxg0X
fN+PUDh1BwjhRSD1kME2KWvjz4l6eGY3T5ltS50TnTQUsCo6vXemTCdlBxKT
Y67SfV5ibNHed16FM6PDuYUUKbeslqu2VeuUWbnj4QYI5FrzSNyncv1bxIFr
J1gVuMdMdfIPh+r4aMDWepgu8R5E+h9hasJvbepzRi9J+9iavSeD/2M1W06c
YLyFgG4mM0fzrcDcrD8k+4an6xtIZPeTJUxSzwHG72sZo28AV9HBeKsoNtkV
mgCtXV2C7qBK8GgOrPGJMNgln63mqInFZETGjagS5XRtIYVIrpxpkTsjWOmm
jySbNIBox6FjZhNsgNt8m6OoMmGy05Uq3UqR61j5uHe9abZbe1f1FHBfQ1tQ
0GzpWb84NwP7S6fdEQxALXIiTsmWF1f/gDFk2q6dr3YXzVk5EQCZLqQlOUCp
P631s4WCGuLq0Ufo3F2MGzNUEDGhq3oQqMPYCGPA25hQ1s7YojBDUVVN+hlB
da34kPYC3PM8f4zTh9AU3nuMnrr9pvJ5IPYblnPuzQjnc2I5Ha6Lx4fxkpEg
J2QQPBJjCoAJxat79EC2PNxdBFdEmRPav70ApNViye5bMY60xWtYeXSWMuYS
Il1Qn2OloeeoEaOjINiJerTDBeaBTAreEMlHQMebSOzL3VSwdbpTv191h8nZ
S9t4gpxJAnbIYrdYg9h4Wrjurif2QHrqNmpG45HpTbdqI2cuPv4KOINYNlp4
RKhxxdEDl5yXo5u5ykr9waYB/YwJTL+3fXZ6pCHCR8FHxcOwbX0SB1DqsK/0
HMQ4damdPklDqMhCUm7zuihbrgeGJIjyZYTQzRhCKVrAbgE3HPyZ0MFjNJNo
skkFdmdeuASWpwbL0bF9dEAOKvk92erPOp4ucIjDcqiPkVdXxcl/KHLg2kjH
6C0GLSmbHpN9NKAnhzlh4skDcTrDvxL7wnaCoU5W8hJYdVo43KGZsBqGWqcA
831cuOzGpvimZyTFZl8fUtd2Q+llUMpNEOKUrLsEqsLI6VAwEugNoQ5rMTbu
dHc7DHBD9Yim9om2dYGyXo6Z2amBFfYSLx7yc+fZSa9Qpb5UbvQYBfRwe7Sc
uhnjlejRP5hh7WR7fKzKOwiVxlY+P+IQWsSfEeahYcP9Tjdyjw7tX5Q5rD+E
em8h7N+jxhM6M4EXWn2CuMy398XxnpfXgPTxhQawrTFhuMDFmRYjA1NG44If
+EG/mRXydQQREXsYMe4j5ZyfJU6mZ5G8kWzwyhJNa4pELG8quRN3tFmLdsDj
iIRUeyuxV75ueYNIp0M49gs2XDjR/g2NhrOg4RywdgYjiKUDdMg2UuPQ4rqe
utgDZ0u4v+K/eiY40pnlXBthNIcBHkGfQTLHVjHrboDcQoxJsywxAJRbXOIE
UOzEZmN9wJuoiOifH3tYIBAOHjDYywctSxwrtfTz4TvxbYxg2SboRqUY9g/p
ziDClV6h1TGt/XEDmnMQGb09hip7MHrUq2DV7SORad0VbMmjN4QsWTDfDxs0
KgzDRKNAP+wrtA1b31H7dL9360qdyGb0AURMyNchrYpT8z9iYmSKfq8p3ccy
pW7w3Y2+BYAMzKG2xfK+f80AzqxCqHAyzYXWDDPlCdkORqMpqUaqAOIlLh/c
EqgaWloTnHqfKXVpDguEvRlAY7SCjwPd3OXLRBUgdBSalT51oqm7bxBMZvlN
TINrmn8K951bx7LBj+GdM0M2iV5EhnFpTCMLtu4NJ67l7SQRYLDDcFvOpR0C
fPTIQXLWOpjInslVm2UjHyxL9zkCUKBf1Ea3UqsNUrkmzucaMoLodLgVRogf
YCzC1E/BQvPsP+mg59yjJ9ATIZ7Yb5P0PF5dKo2TccZsyJvNsc6R5qCpJQie
pkHgN2s4bB+/4nQqtLR1x9kflCyP8rIkAJTN1BQrchs0ZZZiSjWjIIQ3cHgK
Xm2D2RnLBQnnl0YKkRhhVRtfyEopeUmiTtTIjGVL+/IRvdL9mpmBl0WWMzlB
5zS0Xb5Fv5RpoITxzWemE/XWRpBGKlWRAh3FzSeeB6N8CaBDmZMxrnQqT2iS
DLlKK9Np4dyugKdPZDLPx+na1gLN1bbTHPlqJXocJlha3plVoZI6LtebEZ9b
Qq1rmQ4RlFmwVKG0GG2AddsXAc9aYjw5DLYq/d2zYHjrdD+qFs5A//zJFKx4
cVhYrFR8S27DCHW5yeY6st5fPxGSeCwSj458y/9vp8/b8nv2+0L4RSJ0z8/7
Vvd8EO8I8Kxgft7qPBvWKGe+xG8FbFWUW95L5m3czEsBR4plDUjHsByvWe16
lVRFKE1cjDKEad6fMoqnS8khEVi7Tuy57is/x9bHMojnmVkt2GtGnMI3Psbd
AO4g4U+8dT3uyTteDdKdrEPCunYFL8FZBtOlwqPNjdBtIAG8y9U9wZa11AgJ
lEdTlPxutmavmqhCHyLFAqAhvXLStg/ryMXlj6LocQtkGEkLz3tsE3Psl2A5
mUSPqLKkKuG/q/nTiISKDF9CgSyQ+DZ0TvO0XPL7a9eg9x57vTlvQl/oIziA
UoLd8HkP0PZhj15H5+AjVH4AWlfF4+CHpIGQPMM2HYVCYxThMDOfKmdgz7qE
DIOt4N7z0OY9JxOQbY0euMub1ih9nbtjqt+YSxoUmKBXSE3fdTpOS2dnfP0Y
qNNf8QXSIIymbgJZKJ8i4kQq17NqXdEjK4JyX7ty+18NgKFAE+kX0LbVitBp
/46K1zIMmPVYBm0DNUtDYg4b3kYa/GHI9LYAnLuwjA7H6a+quGhD33UdzRAS
+vHV++z39UI9uUo3dmIiUgBbgI7UCe5W8xJ54+oRegA7kF3DClpvDi5bpUnF
6l8nlB++wFW2jgythLYX2z96hgyI9daFxuJRoIQGWcEwB4DOuicPxLuQD7Ch
LQdpGuVR8196dPLkmgz+7iAnL5xbYKo0i9SAVK2H+gvPVoObZ5SAuR0YIC/1
2ezz6x375m6Lfjau+cpxQ0gqvvi+hkdkDUUfmwoxRtfSdYps/R5opYG/b95b
dZspIprpweYrfiSD3Qt9Nw5yyENartCqagT4HT7UR3TetHK0IRpJnmBWvydy
+B5fWniDrMFg4WjHR+W88fbt+XW6NnXB7BjvbSED5ltfnjro5ELDKLzj0+WT
N3aNznyGhy+RrkpSOPE4nyTyWZss4V7QIoYt8ygWnnU2E3K+wyg3AW6xN7Fx
8X6cB8bUv4i/hYzVDQlhApeWbLzp9Fnas9FmIJhjIw/Q018bMP9T/YiqfcwA
qMRKPPCaJerY/H6bIVUTdrthiiPuu8X8LnuFlnr8lGp1nORdWq8cEUFeyeCX
pp3HDercANoTeZbp/s5K4CPAdnWqF3OHgsUGlFlVPcxX+9A6XsD62n6n8OJF
Nljat9BdIAe/y1s/dUelT+EQJD2B1EaXE7fCNnD1uicepdZIf0aNOGthwxcw
jMLjPFbip1mMmBkYLScz3lrG5ZcYkUROmWt6qedZSbCyhG++14iQ1RvwPX3o
JEQAWtU9cW7SRmEN1qENYpYHYZhU8pfQnjAeh0I8M8PrfG6PoopyJoOiG3wt
/y7HdtJgj4xGMTiFzdTbGVtZ9EYuc+cB+z3lQ63U5siXxrXe3c4uwLYTs+23
6p2UcykNGJBYXkUtTddFhY/1ZVavfx5yy/p3IIfeEFsZOOt0nAF8RdUzug18
v9hPc3OTDhGb+5Ez3Qy4ilbgfNiNA45sKRa++b6VcuHlb9TegzX6lrs8vY2f
xznTCLT+ujFnk7uDx67TnmbFTDrR2G5Z+L6M9vkj2SZFGqpfqkkhl48K0dlH
QUvG4evGulbSO1gSPVxQaDZF1L1nLovdzpSiIZZZ3NGx4fQX2slCQU2bEGJe
M/dp03hkFgIJVLtZrzX8jiKqybvq+XUO4onqb/HDPU/MD7XdIGZxIt9XT8CQ
Fkr3+uJmsqjUasAxobqEyT+DzPbt3jIPp0zLV6hawN3h9TuHDm0OuzJ0pFT4
oPV0iK/T4W4YSeYev56HJ8Ntf7kI/mbqpmwN6L+nKMvBhF5YepTdLrrNdAXb
zG+kER50EXoe4WcQUULkOZNmV+S2rCC4bHPYhaZ1Okf91WIz721b5MgVIl1o
ajOt4WGKZ819LNMJMbhQzgUO7kBFeAjJc5A00bc1QwsFVbiQn80A+nPepcxI
44FABFPvRllp8hmtsB4ODW6kgPxda9DIWHu1UqFzTP6cOxdBqammxTs4f7ce
x/6RPNYkffC7nH5sA2YMsd85Jf53LJQCjw/uXNY+56TDJrAeDJMab7x5F/gl
hCefxAr9G76chfbekxpwF+Wf5q7mUO+OHlSj8650A8cXeFRUce1+RIMwm1l6
5NQHdu6BwMt1LtS/yG65ha4qMlTNa6cCsCRbpP6QWvM6/y4FTOye2Q1UvAVc
GeYKz7+r5HKhM1+6wyHkCk6yygz9X5sGdioVOJZyOBcSW93aOVEPF4+dn0NP
Ni6W6Q9uW2vvkFBoVK75H4YR4IlUygwp6vbPmqSPn/ITBQvVG0rW61vDN4Yb
O1Gbz0hg1juEs4Ry8UqduNuZO+uXlklJxzyw0t7V9xS2Qxw9BcmOCezuqeMk
n2HnEY05awqxZwZjcf4iWSoXVJYER6gff7i6zbH4vVl1Fwh+S261U6biueeA
pcxnL9XTYnXFuvuSHkV1P+GSif57Citf5YSwW1xed8K59H61ZeSimzv+PwGB
znsuHC7m+vWBWNF0QmgcBWZ9feuQ/g3lP1/ownEGEAHIrskG2lN+vIDDbtGi
k3FXkrKctD3+JPK7TJFSm/aJMoI8IkXP0QgoHrqn4f3JpelkafnpQ7eNJV+W
rsWyK6L7DaqKgnUffLp0mnAg8kwstROldK/Sn7z1MW3WkzMFDvhgvuyIXz4s
3lbBqaSBY8sG3O504lir4ZbmsVamtcW4tYxjdSR1oqAqHk7NEn2c7XhdWkIp
t3ykAj7JB3iLlJgbtlkSAuYa5YwzjDI0ob8YrzsLyg0RU+X32qD5naeiPai5
sM4e2bPZKnFg0Xo7H0YKmESnwHdWzJZp5QYEBgjBsi2BBhtqFYR/vqJ3fiK0
3YBIZuR/Xccysh2PKOw5t6pDr5q5hzB2L+O6U57LnuMVvqR3SgoFXkPwN8E5
7bxIgvmx8JTUjXGxiwpkFZ7dBJtfx8zGrmSnPX8OBonlCE3lbNlUmvUbWeWj
UeX+grclBlZaafnpqDni4OL5Sg2QdeipAQ6EtPXEP/W+7x/hEjG+9OQhmv4/
g1LtlbRCYgDxazdS6XLiROF2n6fuc7kP3/sl3sr6bw+VwrHntF3NYzZYMac8
yVgTtrGKtoNXCkoSBudxFpN1hMjRkZ9rABBPcQy0zkUyy3/60z3IBFwUtmF3
Qh8sSAjcURY6xvF2tb4t5O/X8m08bVOPSRaJPzIsiUVK43w4b4R47ygEFIaX
2YEGpNPjh6dP5Ib+F2B58wc/aKL2L1PZIF/HmMBf4ysxUEYaoDahZ3NZdK3+
A+xR3i+WLhSXwE68/lDcxbjGhNEX9q/qdP2NG4a631QxfxCWbT+C71lUyXWJ
Iakd7DbUooHIbxLk3s5O6XMU47lWG6bqNjoierWOakq2MWBq75+LDugnIoGx
h70VDT/6HK6y+I7VYbkatLZel0jmRhX2eAuZc6WusUcnuvyaq65Q5uc11jik
QMyjPzuC/zIawTwJchfC5+Hs5WfZyHqeJlqNcgA18QSrs9gvb9j0Y5EmPvWe
BkUCDT4wJvDZyLBYBtHN11KHRHex8itCDYtD7XVsdOw9Wyx8CU4qHA7thI5V
c1GAsOnXRwX41mqytHAJ93SJTbAQ+x0kz3ihWG9TQThJ4Clh4Z6wb+Rmmi4m
VQEJbd1nNJlBcUU4G3M8lm4y34fvnIlSKZT+xGuy2svFGggWb2IKbWqZHFvy
Com9MRijKK5NI7ORAHx/4K8x3qTPADA9vVW2lvHpSHljFB+Gl53jIEutQWVo
3TemVr9cCmftvvUKj1bo7JKerNoCSJzhVHKSHe8yIXDqhldX+vKt3BJDHbLp
briJuNvdRtP8N4jCRczpeGFewjybkAu6jtiubvCsYWfEyF1nBunRhJvTGWnd
UMOEGEWkQrVfBKY7yJc7A0sahyPmpyBQBoWRM7rozlMk5Gw2IGLpSuFeHu78
KyeSApWTesGNLqkQahplButxyh+NZYGeJLWnWf9M5KlPMRuaicPvreZ7INbG
8OtGiLbaivKQZOsK07dDHGzbkVm51d+M1GHdvQFG6OyZd25+4PjFqfgQ9owP
UW/0j6G3kxkxxJruhhwJCQse8rbKJcW5VeVsz2IV+u4eDuCHMLsAlgj2UXo+
SAsR17a75KAO0SnI/a0RLYcINNP9XG+R32lkOuTDZQVVs+OjFFfq4lEg/+9Y
gdbTliwJqv3SxOkiiV1zGcAkT2GEvgTvOoZW81CRuqyiR9Ip7jy/tW9kwNVZ
uQ66FLNHdtgq7rr3XxNTL0u5GtaF3WjZHo8yoACnBxAM/tH44X0Oga65SI+r
TOgQnTytNvq9uCaCkflaovQdhA9eVGWiCILJ9r6SaU7RFo4/Smbr6Cq+rK1r
0W95bGh3eWWfCPZa5drzAfmkm5wETd8x+R3MMNMoXQizV2yseEYn6Acmoy2e
x/Hdu0gCqmxOIBWJDMfIeX8PwzqLc8WzUILbGNub+ZUd/7uVukHDa8MM7BkZ
73vXAIO+e3OO3uWuhmfh6bHlizeP8GekD80k1HVoC10SAVy5LvtXIjcO1gSG
3Ma9VdozolWX2Tl7teIJAtNZ0YefSIMy67WnSk0yCLPsnhif7yu+JRsPRdK1
UF5myWonss9TYv369m24C43SBTo6xpgWTlwa0366iFw4ZN18wihnc0zLQZ4l
rJZd6igywVJkzzPjuqgJEpnTiv7CYJNZj/Hnn6bBKa0O8mLHu2teBrhGu2DA
cf+gUAjJReM72/yAKwLbMeMvQ843+BJ45JGKjxnLiT5cNMWxYUPLPJ5CQSFw
88f20gIbPruXuxLTRSH3geMQdQcidkdPu5D89gq23Qx8BRwKozpcKYPSnvvC
Sz3CzpklJGeNdhtFVMmSq9VBYvADyIMAeqDfLdNY1ZtLu7Lc8udeHQHJlsXj
uNPWTgG7MD1xmLgqCFLPlX/E37dgT07OYpTbcdv4l0gOsQjF8eRJHdLYkUCO
g6VYA0hlBCWhCqulUvj+ggRzdxWcsLbg8E43YD/UvPVH3kIpKLTbbU5OWCAR
v7b3GNw2n4hvduA1HVcif7yFIHZLuJXUm8rtYHRT19+k0anwMYIor2WwGEu4
yeVmbP4BbsTB5DfdHApvW8to60KuCPrgmoIxeqPkhCy6FB411TnXCCMG0C67
6pwEgadOIo+Uc3NxJqMxElxBa4p1eKR3rIML0MD2V/AutS9pju3z8L7mw3hv
uoZsBpC961xUn0HAW1mnaDAysxg5r5sAuTtTo5GWUU/25n0x3I4xTtky/4Qj
K4uccgzLpEYb1n/8WHg0GMVsJ005QWSaXmTVlUiAA6kg35CZaP52b04nQtdO
tH4gPKnOzYbKQW6eqMiBJwISWw0T3x6t6j3akViPDMmUelZHjo4LTAqJlqm7
O4qkIj5va8Ok6Nm0Z32nIGViNRPdz6/cT/UAiEUOt1pZz67Afo56jvZDuHmV
YCRXxmlr1FX82b8YZ0FXJoZQAMHZQ4TgI7GGzV/8A67cfItYdjFQwQr/+wGy
rzKC2AgePU0XspBF+lZ4o8S55k4AqphDut5B54HbWvSFq8+C4ABBkL3AbiSA
7zdf0ewIVBHo+V9W6//Byt61I/qPHlE2dz+MObwqnDN9Qkem6YmPZ7o4CbhC
0v6wWUIUQZJtkRQV/HLuCUofmrg5kWR4SinSoJj107tdTjUZw9cOR3PR0/jw
MW3EsO24lkCYaj5nLwHTzG1+3CutKmtk8hvdxnHsnj6lZumnvpTc3ARqiSEi
GCur7tMX337jrDASHdtwKbzTdTifXlaeyvCb5CHraXZziKH/u8VU3GEYZW7+
vmY8HLXgMjMofw420Dtf9+FhE3fOdXmvEvPYwxqf22DkjzHl8h+U9MQmCH/A
+mRO29PghF0xYzbJOIFfesQeIjcnRa9/SN7Irv1qrw9UhrPaoXGYWruwohV9
ytsj2TTOa1kjFJjYRCbgOxkM2qJ04/+uaK72s4NoLvQd5yj6S0QtCsCEGJJI
+5a51K1N0rRfzrQQ2S96mn4tIihe55Uij8bzkeKcGcctAVr3M0zmyCDWvW04
DfNYSBBRUF1JoArL35FnvKdQEodwP2KXQl395gO+DUIcKjA3cuFnn11N095N
Q0trQA1Mo4j8nrFGS9BHY0vfdHSTgFRpUTeyKQSExXWqcHAhxg/aM0Ez705g
8/o8s2tNZ2epD8/4Tp6y/Q995F5wDoY8YINOh08DPRgkqjE4MDybgZ3pEaNJ
PBgqS5jNOAzwk47m83cStF+PGmiZpNvAfMFFwec1IQNGAjQNa1KiCyg2TkRT
mRpyZ8qk2hJyO1zDTNlVFYJItiXF4uHd0HoOIFGm76EbVSGBJX4nn26c5QrY
3lQyd33/whnLpymaniEHvtHTfIHaFJT2DkvfTlhf7UKnaVZyyW3wfkjhnjpn
Fan1jde/Qg/oWw2wjwMoNjPOscEgTbZS/BZ6nwTAuKcgjuJmhgP5hxwWF+mB
920vuQL55YXi9agaVL2A7kjoARy0WsmJKCZEAM57ibmdQ1uPzJJRKA+dW5ik
88JJzw9NhccK0dlEYgfvEFWdNaVQi2MT5FNOph5uYO5pVrWMEL/POEZSJI2R
NB+WED/2vZ0bYiKPV8oX6GHMyMR/N2/HYiNV4s0PWdTZUnV/kdrRSEnjaYmC
kZuHL7EgixnZXqe9HJt0ktCMkmjnz2jNyL7VYUpfXYdUec9VteBUxUsfNgB6
nQDtdx843JLwC8l2oV3SWtI9dgaIJ9Vw2U+A5BWiNnvFAEdEU/vW9JYQXuQ0
UmAZogpY7nBHx4+9G7IlGe21ql6EpafpiV7nU3kyyvOLWj7aQm9F3CDngeO3
jRvv66jzy4KIKKIzImD2yqu7LYCdFTKct8skr6V2Z7jmRcZz+XUY+fyYiH8P
8IkxtKTgrOhyGYXS2JuihJl0Auup7wzTTx96rQswKkdJPrTy3kQL/pXo23/l
7Yl04lMx7JltEkyYQwpTlGqfNaYngKgLZkX67svZ7KcrLE30VPC3afmdabZ1
j7hFec6EW3zoLkKucw+Drx3Z7kpX6nNZgdHZPmropNAhqTk19FixImBLrqTv
rY7FxrmCkFFy0QsdhW69FXEIYvb0o/UAAOXssWnl1zomryJ9KOhffkF5KsEg
uhj07VkxsX3U6JsA4pT55mTDeoOCcInXpRhC0YRgzk63klrLVtIOwbmM3t+Q
eBmyZ1AbDqcou1h6nC7cOi4sv9/WnkOFRzJHgZnWf6LuC5qu2NY6p3bmvzvN
fXrEGfDW+pIe5tcbUF+y6N3T/HM449Yb2cKryyOq5YrERu7/+7W3K3C57ERm
2wGd5JpGzyPeUrNpGU3k5zFuuR9PeJF5SA+sPrdv3pQEydWuATBdLPwKZ2Ez
/tCNl0hcscKnHUGJfudxo1OVHuOImU+L0kVS/exbLX94s5Voc9iWoTo4SpN0
dhx0TzS5qK6Abw95uX4DZlAnwG2BSclCLJdACk4irlGJA5svrny3N/sjJkYB
Egasns6xu3GeXCiSrsqC2KFAnpNHpSDUFT7Eg9BBv5or1ODt+OpjkUO8sMoe
1395VBQHpSQzm2bNPXFBJ/HnS9djrfcuBUdXKJ+udwsjjuZgh/s8xAzvQaXZ
vdY1VofOfBRjug2TKHU6QRG4Wjq5TBI3IlK6i5v10U0+LKMGKgNQkFbzbqB8
LvWlW1Uz0ayqTOCh8Ie/L9NnIYZ/kXQaQLIahIrsE73SbrY8K6G0FinPmEoH
4nydFnELU1+WebML5gND/Rp9FAaoiJ/jOdPyFZNMpTodkwpK+gckhaQd0Wki
3Sa2ejaVGOdlCcu9TMC9+/MEkTUgWeLoFDv4bCmuYLv+Tip6bxY7gVWTforx
vRkV9on0sPe/uhzCQU8lNvNRkYVqw1Up1VKh4Bt62/z0SZ/0UcewxWmdm9a3
DI9l7wUAvlG+XCGHk/hfZyxuE0DKqsFwhv2lhFabSDafnzur6V67tt1TA3j0
N1RUnEc82zm2qtNLUbaCIOnolJ4b5Ni7eosjzd/PqN7JYLaWgZVkzyKyIax3
tErWsRZuuBq0UvcmCLt+izeemWqcLZ+g55+UlAzuyHpUAlcJCNbZJygWvz9M
lIDEw3DlqOsvdQQ7FmGK1disI2ZtiXMFUknoSszDBACYdOTg4ism8d/V+Zul
Dqo+WksswiaLNfzh2UDempwnSbBoQweFVWihRtYsN6Fbw7yOdhgdmQ4tfq2Q
DrWcoWq95xzYCCxVY5lp81udx0lJm62nF9f5Ixppiqys9E1FYhmYZEZkGXpB
qX/PCxlggEaGm/R9weJKmC5n4Y935K7NXNIIHM/U5ICWzODh3Ecdjo5HuZ9r
hMHJlWiPkUbgRrytGD+gcz7KD8GeoEGGqQmSmyie85uJ+Wc+7UwvJj4HYRT/
EyxCUJAghMnAbebNVPlcGQDpJw+KwjMoa0CUp5Wl154yI/KSGo3J7TBCsmil
0PfzeFvh33Tnr8TYhz9cDbYIfUP0RvrTuRAtia0DLhifL6MFFnEieUHTkxDV
bxO2PoszZgHX0mSnY3V/LqeSdjzJbyE/NpwyIw7a7HYLdsVd6IwZPWQa23uv
zceJH1uF7q62Yl6CoDRxEnCBQ8RPR7SPbSjVEyNvdgjwSF/zCfyA0x2tB476
/wMhZZFimQWwwks4H0WI3seqc9c2aSik/lPRh43Nhv6kd7UhHrNSwIz1BNOM
bvqoBCH4bdzrVYMarBaQ/B1wqAODs3tSoN4ki30MjzWfdjFEfDYizxAQagv5
XHH6hGxJNGjfeRSZ+ICaynZciW4HKe1wUnFZu7GKmbjBdQFhv0/s/kH+6BAq
TsjYWJo9o/4i0vv9a3InZbJOWaxw1ByhCzADsOC1gjEIkd8sSgEt7s1GX0Z2
J4nYM3k+WOpyxo/XmuwTxYlAj2DqqjDIsvgdFlwTB+2d7bA8bol3K5kkkVua
qVVJJYDwSQI0jS1SoVcRkVpn6StqFJltzfT1JJbnMbmmnFhHkwrHIoPkb9Yr
4PFCAyG370p3KjqXiNNyQ67bmioUJhKlEEyfsMkAmIQXVRTVRP5qK4/5o5BD
TFfrXf7Uhnm6BKXwnJA2kkPZhYS9N6gD/M/+HjQCLkRzN53XsP+VE8d+OuIe
Fx6tw5hGaJuewMPCunZxASDu36qydPu/Gr2tXXAGVpbGncHqT0YKuebAB7fO
NKPHQ2PtoEFH23L0G3L2LjCKrsPC6owHkhDQzCQB0IHi81wkXdgj2NpNLxjM
xeKwOqxnHXO2t7CO9QqtRuWKUsPbhiB6qKOUbfmdZfrnlO+15trheIDuGF0q
oab1/8+R+hMPe7IS1rw5EezzCPGgSwRfnWfs2YSw9IGM3o8HrwUa/R2TaZxc
2oIAn0z9Bw188tdfLGRKFAlYx5ZHjHvpYSV5xI6oLLijylOVd+vBEGVmTtgY
HF8+HkOTyahcD2fKzJLEJcp6YQyb1chlFUBdHsDVrFUR4jfToqDHTMEyaIGI
6YEGR6ZmOMrH2mK1tO18ELzSLl8nxyIJFOosV9xIvOUbvG9K8jDF3nbTLE7N
m32ZxFNqMvd0qG1ExtP5myg6+g7FQ1Ihs9Ir0hcc2KCSHl9q2OGuehMrAX/O
5Eg3Eexb2NeR4o8ppTypPijWBZe6VeDt6Pv6J7XiMaXBgV52z5aOBDGSx/EU
nULNiComEJHELhrPcE21nCF3XMWCkideqBYn+LxVnkPql7faOOLLaCF5YuFb
Vnd/NqWgPN3SkUSW07qVO2oYij+7Hk0jwwIJHZhu8yEJAvW2xoH/rYWyeaDX
y49EQ6dNzq1QZZd73It01ZpJmJorNvQUmKldmHizVF6KWGyb9VDn+6Fr/bzP
eL0YFm+A934hbXWyN0cTfqzhfmVWvdgYUDVy26lPFgVXDIK19QnDorfrc+jf
MhVK5wywwMTA+4R/6Azvi+UMo2DYJX2oTH4LGDnXeODMu9kWHPDmE6ToFJvp
AG2rVWD4TiXLtBZJUlxZK0uC3VKc1PkIrQDybnWGi/0qAPcQ8zGk1y6bEnKz
8bSsUTJ0MBvpip1p8ixXpPn6eJnBUhw7jA66H/4xbVTSWifm5pG0tZjRax2G
QrqNic8Hl0BrDEz8ZgX+z9vC9f2Dop9jKV887iLykRX1k1iX+Bn0fXB9YT5B
7ycMW1D//kwYbA9CyIDleS1q+hJzkmgw7WQ5YVQCec3fI8uA93j8U1hYCRv4
E2g3iYGzPBB03NDvbn6qoL+gjY+fpI39aR4Q+OcgLBRMr8hKHVFN8sjiz1g8
BuYlCcUW4n24Xbk68zLNZiC0r7VufM5g1Hq1BwyO6HI1pLPFjOru1mPk2LFN
GNBCQvXSihJStXF+6d+p+1v7g0mKGMqODntVuk8+AwNjOm8FUMKfmC28Qo8D
1/TqvwPA+kNoU6VE9GkWsvtzXPTks0eiKJnNQvzSId+eNqX9u2FeMFNTHLNy
UY7ha3CL3pwCV9VPHnKdi/BV1C4g9ZLdjNQBmUM3d2nm9yxTP3yVusC1UVqq
iBCxQBQqA4TN4NlyS+x6I1ddZM63lVXz/00Aw6T5Vyl4DWWYuZhDRPj30OkM
M2ukaSEBHsVFgL+1zGr8lD/2oKIOduAtccQydYRHEirCidfpCPtxdtenCxZY
llHs98FcwdBD4dpw7nJcGAMjSpwllodtpinf/7AnLL2U5FGWDE/A1skJ/972
5TbJ4izLXSK4MLpQBUQufYCoeOrIkSPlmwpcUQmAPtMZdYKotbPMffMuGgwm
j9quEVP8fT+9LVuUzPJOWqq7Dz6ah8Kh0VH3GVOarQM1mBxEVpyBKs5SPeGv
xKGXO/vZndXYAtsL7PgEtxGFGpnl6Jx/3YTuM3H0hhwmZ3cLPfbSSIRWmo8U
uVTKJ3bjNo3OCLqXZVKY/7tdR3rVomUxq5bfVVJ6pBwQ8IWI11plbi6OhPd9
9lte94hJlNqgNFKmYYzVz5Ks//H5M2AaKCYifGr3RLIIwj0jzBh9+wItWcWO
Q7f6KyiwWYKqgxK8tJuyAXd5iEDHHFd3ocv7u1Xob2l/MSemTFHvQvPsZqkt
/TAAFSdL2XwVonAG0Wp2bV6t7rcO0CCkIW9zQkkvy8tYmtxYd/IFFdqOcW6C
WqLMW2g/I/vGZF9B7doewwwj8oLLijJv6aecg7eXURvORTlgMgmL8JuuvexG
atmAhFK/iJOc+vT2cBBuwGdgg5SSGtMCxP/8m+Kxmbnk1gjJ5taMehqPUC5b
b7vj43iQu97wIGTBqevUcStw6RASaXMyDsFWzf/2mlEeAW9FKv64MkgHOHJj
T7eOQBirosV+0SO5eKjCPWwF+OVJUaIKM8xOu/b2f47ly3fB0Umg1PE7IyAQ
ljYIaE0dO2pwutgq960X7P4erJh7yYrWkjB0ah9fw/6K7YdU5RsYyh9AhcID
53aH7zTHqo8YguneevVkKx8OnR1szOEPakX18XZp69mSbGuIKs0cmb2UgMKp
kYjSiO/kBVQ2wRibmOlPEKl3o+l0drFCMHjMb+ozRHa3/BFkavhZ8L1um/Qa
IN4HCzgHXevKbwN9Zc1Xg48pcIkhUNMkGxBV7R05ozcliyfI734iNmusOBW3
vXLIPoyUw4Vee7n7gq0Qxe++BS+WSY1uW2t76JQIEouQdcy4gIdoh/Kqb41O
nLOK/QnnXHGKDxIY+38jUvqXyqLs++xQwXciNNIQO5scohXtTVFya1c5S3OB
NVP2WXffqNDF9xQUmg/HZH7l+rJp2lHo03JB0g40PlfBsTv/acvzddahuni3
3b4SfRQC6AJfKX/KnGjV0V8VxY/ulUMTNuKTamMpcY2d9xOrn6EA5xND8krQ
oFlj5Db58o79Xj/jMd4SjsfrLujUDeZStgckL7WeyVK4oOAYbg5+lqg5EdO6
uuwxxxg/7vMzBtuE/dSHj5mym6ajtsZGPiR2WEEmb8nk065P7i2p9RRaPXHP
39vjK7L2HLpxTzHGJGiMRj1gxwaxDAPK4J0lunkCcZHbxJ07KWwpgBa0glBQ
vWJoSOP4k1m/TVCRERNWDH7lLe3t2YKH16tJBIvYWCWMPiEFWdTiAKrfLd5t
LrBRJElZ36bezr9fNK4Q4p5rbH1wfzDDLtOu9sgu8rzKb67Ih+udew8ZxZYo
Z2Os0yWqGLufLEdZuDdjI81KYcIaO/6IxMCcv4JWSrYCi5WB9KWEFpN87G6w
Bcyi5hLVWa+zY0JW1rguxeL9J5hgfvFNLKqvhwYARnF1nE07MX2tTPmH5w8o
zq91on23hWBnq/QtkBoAgg+aHKAdBnADiAuU29NdgCD+N5nitnymckRv4N5A
DvJzpGJDB0NigxysibRwy/SnBYwEmtgNYA9S9eFQ3z+uRf027hYZXYEaCCNZ
xH6U2Zs41jPJYnj/bCYbn/y8hybNTyWj0p57wUwo2PoXjY1ayEnsJOewePfW
D5ZJnQG4CuAp1Rue1lxu/toqc6wF/Q6CkUl7SSOUISQOZt2Bv3Tr5K5gwWL6
03XsPCN3HbGqynSTQok/wJ784jVvwTzeuuUvh8j1CKW6iFoXrKBJK6cn1JZm
yziXyrcux3YjFs7gDdHEYkcAZaYar9BRGeuswWYMLXxqz73/G3KZvnlF3g87
XjlSxDU0uPdJ2UfEsBRI5pQqvAa7VlOWRuNvROaa7KE9AW3afoBVYzbCtYK/
Y5ctqILtQTLVs8OSJbj+GACNomN1fBsvJ+cheWHuzuppsgkAYmZdJE2hdJ50
miSCMO/Kns118/vpqEkuovQ0jBMuO8N6dygsjpBxa3MfyAlPjsLMSW4Gxhmb
tTY2Cv6/jKgM6nR789dfmlpfakPcVNf+svj73MBMhxWfGAq7z4hO8L6der/Y
YlIhTVLHnD+DY3eL6NcrHALJ54fj4cUf+NQrDXn0idmdL3wiRoGpjR86KJ/C
Mr9KMRJ1qOdQLHfp7T+04tDCwEo4QTPPHjJsv8u6ETJqpgiiit1Ix/BkDWYl
HO6/+pM9xO41hkYZu0mZT7qjWwgM15bQEKypVaSgUIOTXwi2bNJuqK7w3/Nm
73Ooh3SSgj6qTWKfsqmk3sTuTJ+VVTIaC433HfU8T+URbIkbh53vutHMLr+F
Fg1NEGBBxg7P4lgehxXKczWiXpQBU2Stjf+02stDi2f0VFVVtpCqHpkmP28X
x491mUHTAL8kH1kulgrd47z9SNoAWr+6/wHCAKaFuV39GNjU8Ga+Yind5wbn
EQJ4/t1ItgMFp98oLm0TnKnMru1XYU90/q/3tzxvoCKZegZmFDKjQiGMNjCE
xkzZGV1keBwvxOKa1u5/AWOrM9aoYEqlUmqyQKrsbr99y6r6DN5PDoK+mxMx
JH5+47H79Np9oecTfG2G1/fZG2Yc/tXxE7updxGOjSbFCZtmK03kSK4I2NIj
roJQn4InTBKB3Z2aPODxyikQGCPG1V+2uDGwJ4Za9NrsQbYmPOWaOmp3uCRK
yxxSNa7tUNFv11ubAtK+kACc9+P4lHf7zaeEvRKSpMZPrbXBvRrQ4puSszO1
o6HhzFQZ7lLvMUOFTkelm0SkLeYzoz/rUaOxnwM2mj56RYFhwDPq95NqfFlT
T/fo2pTI+NrpLNC55CYiWxa8FjZguzJZxrMXNY8zQUyQPsKj01NGFp2TWB7P
hXp8GgPDxwu9C6VTgx4JmhQ/q2xbaftWHjhCv+B5DVB5l9fQie4dSH/aPDcO
sdAZJd9QOljl4n4weXoNhz17nUcpn7gDedaoHTTwBM8HNYEJ/2Cwn/ekhzh/
GXnsEPAhPSPEYTOfgF9DeIvu6GmnnViJv1jEslI/PDxa5UJJGiauVgNPb7zn
gzYA+uJ84cKX7JD+00AR1Zc/YiVYxGrMBM4eNoRbvJQvj4oGvz6994PNX122
iqn2z9y5KuYO4yFjIuqqNSjGSqIUlWow4orBFYST0fnkGCuDV/pH75G7wa46
RY6X2UECN3Dm7wVf9FQrZlZT1UKojHiDba5cd+5sKRTSFZ8qzq4Ih+kWDBzj
v9nUdNHx79W9/pOGkc6g2T9amt9Y9zLQRBNTudNoYS2AaKTzyG19+kbzbG3i
xDG324e19tqCmHjKBXi9oDKkG3U5ho6R43mu6eoW9LHud2lkyFxxEgXAWmYm
tJWB2SyEawT0o2vIiJVdUQJUvcuDAD252KLHunAqSNhuSKNuh+Yhc7BPylc6
we0+GLLxeFuVOigGKSCdIEK+7wBGJyyVFDTUNsBuZuzk1DiHYVfU6RDiiFIK
4jGN6dD450qH3SzHP/u22b4LZs5B1i3frmMuIr2zCIlScu4lNJGuCNALqTFw
hS1Ube5LVjphylYrciMP7Crd7xV8sO/WC8+ZxXqbP9gtTmqPQPDC9zpaJegO
Msp6eMYrpvfk/m2d+pktxfw8RfY69bGAfufQb492iNcMBasHCh4ID2pL7L0M
/FzwIqrPnO/BZCUWpGh9i2UvaygrftWOujW/p02uSOYR8tZ/TdtzqDA1az62
KN5GUjQS+GYmBSx+iZkZ084wsKCaNMDppXpgwrVOMUjTPrGckTq5G2aBdM+S
EGW1JC7RHgtQlJGkCk2mArVyO6Li7XBHzZ4H1spgXC6KdNohCM2P2cUTzp7v
2iA5NzlAR4DEgdGDGBp108i10q2Tnr61Nw2re9hjpHOSC7+pCJlW7TkIbEPF
ZJ8P0g5jRzbN0jUXRGC3F74KcSTLepQBuU3gzRhu2vQTgJ32CxE5DfXLKZvH
y4SOEUyB7A0XsRI68KGn/TENevMQuSzF+u6QS02W2kT9a87kIeN0EtjJs17i
f9drG1hqbmXfpruMV5EqZPR8cqYbOe5G12oYrXE1X88t+zRYv9qu6QP6YNt1
1TcPXf6jURnkpWODJkvercoHzRPKcukU6IHcdpy/6Gms9xWe7cehnuzL0mQe
mae4ncixmxS2sLSibH7rr1yHUBCXbROLnoPmpIu6h8z20E3w11Fv8Wq4jd3l
k+a6/ueeJF0Z1H9zD3FVZp5Jass/DNzo2mF1648h4L7iYMg2XMqKNiGlsw6f
FPucREFujcItaz5kdtpW3TOFcqGoutqWIC81s7J6xyJ+0vN+l136LvDbZl2+
8TMsnO9WZrbEcZ3PT0m3GiKjVdJVj5SCALISA/szOzQchPdixXfI+oASgYSJ
L+PDg6ReIQQgt1Km1i1XbRvYXprYgbxgL5trhVTknBhY/Gi5vcFyJaEVNPN3
9ZiWDoozaxu304Iu4WjUIOxmhwSux8XalOqTO0F7pbd4Gr13nHOCgl2td6q0
Ej4hELL5YzmLXsCikKz8gaADdEajTGFjS012miRv+aacjteiz/IZv4hgC8sz
QGWlMlug0d6f3OqPE9uWDWI6e0agWrC9vEYibjP7tCrXEMojpp+Lc/YHmaYR
9Qm2g1JbNh9l8fpL52/5NNYoilPuS8nsH7P18bty2qhoKYcOAA6NLDTTtUwL
XTx5fJ4zyP+5FDrQ7hO+NMfxdjYxnOP/P7utoaqpBzoCvAGKUceNgZjngnhj
lg7tyHGRZNdoRzCtnXI92dNo7qU3kr+Hs6l43dEGNovuGatW05oMfJjlTXVj
VLoxaPcOTsHUtz/NLIYz8IVquapA/R0itwtqwMIto67/lRdUdXrOrm3fUbBM
saz9I7p2icIpKYKd5l4gCGVLQR2gf96noAnAagnVCdV9L9sxbATi8Ixjp9mO
BhUQnT0IjbrsCStxqzjU27+MISRR9NA/EwwAcVpvPnwkpkJl86Ebwmx43/k9
37wOwfBZAVDW1XZW8gTKA2/DBZXF3d0rCmneIka+tlT/UAY3zFqghqSpAdcP
p3TQJYEb6tW/v7Mqey5ETv+lSDV8GO+V56ujSGQlYJf+gCC/VSj50i4MFes0
Eqg9SwFrSs7dysASJaNJxU+JqTBPVecieeX+2UPl/w4XWywqazouHl27Zw+7
quh6RP82IIoUBbL4Mz12aZ2shN76GTW0QhKRfsH3eiiL6MFvVK5KtnX5tcws
yj3/QBOB+92MKTWNZg5P+PEg1tAx6yHgitVVIJ3Sh+ay9e6cpSpgVx76dIfK
Tt9jH8VeDC2hfdlempIXgzKSq/SaojEeCsDp5vdymMEDgzKswkr2HnLKQoYe
WCQMlEPaVsP47df/ojUJBJcRbUBKY4GKCVV4Lv32kf9foE2W2iu6lbyRatKF
Pq/Amy2cv277DTTYFA7FiH+HXGPjQGt+1LNaBdjjoNv96e+Hi72CFtxQ92sQ
rJ3JypW3zvO2eNKxYoBsQu2BivaMrHAMypsKQ0gY0+rbm6vbR1QdLkW4qNbL
z8UQz9MeJcUVJa2dLU9hNMelyuD3T6K81PISvX18qQ0KWDuRE1XCipREPgU5
iMZTUS+lWJQxy10d4AZafcFAmGT60QFQKfX2hyyj561UdMUx2AeeZWYeWxz3
waiNDL1ZfG7LIGYsHucnVVcY4bivT7jUAg8fs7G4ccwv6SJ/Ubsnd7vzpKpL
0S65Le3xUxkCNU4Yw4674NCRBKZ6C6/OQI5kzK31rPgiRO4lOVFVy91KzpL3
D5gRFOnBiGT9mCEehksqVMUtNnWHNXhfCnvWe/UyIgySUo231DN8EX+FbEpR
1HEJYVyWz78DDnK5HTavXB8J/5dlNUI9guBTX3nV/H3NIOcAG7ujwBFtoS55
A/RDS8qU1TS6gPO2Abi2kETbRyHwLk/RYKM5t/n1gmXfkmQOYjKlun7zko9X
c2bj16dAqSiVkiVxhsHWpzEfSLX9ytO+Uv+VsFIrJ0iNK2KqvBUGbTIIgqBJ
ASqgsDecuY+giwfdJY0DHcVSP76HpoTMdhX3DIRcTYlAAfiUC9HNiMNyAGi0
FaWcR3rzrj66ffgdV5u7SXvQ0511Mhy7vU6x/2IQmEsFbdh3OMpr17KkoO6R
Gmwn9Dnap0tIm+hYYMuKmp+32B6tLh/Kb8CzlB2E0GFW6zlV2Juhh1AomX/E
Rmpd31VE29jX7UmLfdCrS7SHZKaVJ53h+bpK8j56D/VKrC7hdfn4GWqzHfEq
bsfhBJmZggO4EWRDAASXBEEVWlI9OT0ZPaq2dbbK0GYEpy6ZREwgjjAP+3R5
lDxrLidJAdV2wFErs6NjwnR3OdCdDqcpnBSyWMrDKOuLtUeGhK5C0L0MAmca
YceKBQUQ2/F7tNAxLxsd+QBlksJyIUZc0wJ1T5ZnyLVp3S8QHPdvOho0fPwD
8+G5rPW2HTyUiokcD2o7nJeqZsqVpj5arCeYFl2WmrF25t8WXI+RrylEO/9P
1EAtT9RwA+9AoDnuZXUETLL1DZiT2aTSqHFlTJumMZRwgC7fRD5dwupbAk3y
FhVb+IVjXJuSpFk5jEhDmehFIcXn762L7pj+0JRv27TmPt01Y+5I5iK08o7n
gzUKy4OzC0zdFhmO34IJV9xvBL5ElRbBPsckB780mITpB48D+mZ3s8ZtGx6e
r3pzOcBlnwMqACfJsh+DQFJFWB6Qvvjxc8QWXQVq2WK/b0HvXyApxWioYSy7
xw5S2sPCLorFiq1H76MX//jLZZ+TDcwWI7GFTWuF1R29mc0YMsUprdBzMq8w
8/MUl9Z+kuT6x7nmojV3Kb03GLrpp2ZnU0lRCX+LnFvgdlL9dsXyi9hhle92
2r9J2s3/aQoSF6B1AuNeOVMIXmp6m/sIAR+EASM1Wcpmigq9FN0la8IjK5iS
Hu1o7bO2tVcjPI5IBEQQoeDePW0F4oyXzt3AZpajDjEHAl64/J6P7mvm0Hte
jwj2+ZgOnN/OWjKib0C/WTkRa1fQEzj/9n0DPV0tNnHNYVUmpbxekR8av2TT
IIYexn6hWA5j+t1gvPgk+TJa+NbTVAgHgiGmjgWuVBV4GDflNAgFZtYihj26
AN0GxIx518HnN+9/VnPSc24ab9GFqMJfKImuTZSwDJGN01IlsSH8IQkZi/76
uN6VgYKkpRjmwk/ZeHOfDc98JqlF5ct8twgIDa6dTqVBiXrqHh9LovjkAlEc
kJsA6SEdTVswANejLml8SVuLohIEePsy9++U+uj0K6x9CFtiD/u0iEyLZx0f
P49b+Qrw6AB2oLP9ux+6q13IRwtDNGmVgkMOYw6Axou6rFspImIKImKJMFke
Q6H+cmKNfiefpU5z0VxWvcCxSWCiHhVFlzOK3TjSorVjxkUnrZJArd45KBNz
0oL5pN0O64iv9et35vPAhaT+5F1qKWBI7ph2W7rxxhSZxzF3rKuZfuIIDKGg
R87xBr9eFcWP56wndoThYk9s1r4zGxLsoZgWc6MjJDuC3+t1OvDPZm6Y8Len
nFKX6irVw7iVCKwJZ4qCdfEhvgfixuBGviqCjTWgWPxMmBqn7HBIf76hyRF3
BzqvD+b0Hr0rr4BSDCxSvMPeVIECUG9WXaS+yMMe65V1yOFHZqk23fa+5RLx
JRhUiTwbrn46elx06esxPFDgyJc9K7vmpzqxMrKxXwi7KUTi2oUb28DUuBd1
FWleHIeJMaX4E3KV2HMvZ2frGDYl8Za/5YTV/1J2pMAWETcl448B2wsHv743
TWPSY6q7QVVHb9qEtlmB/x4imCkZIs1KDFr6ofTx/LLl5mpojBY7noBnS445
8hathNvoXkHNFONlSmcDBcGPPkLreEJFcowldD76SOchTe9L0jS9wGSciuPv
i0Oha4cEDMKnndQnTCwZSUbJ3oNXj2bIaRqRcUvvM7H4sOKJPUBWMw9otJsv
+enaof98zJ3fQ5WJTf8lDM6O0uUUw2TA0QClCl6tTZe4xVcY7MZh3/9+a4ex
k8oeQgkWVcfoJOWtnfwbggXhk9i2di0WsOMQjDyAbBUvtfJWaOBNsQTKQuzV
PdQew0rES5EmABZj65SD+ey4CXlYoL3kEK9lc5A8HCeiASttAcjWFmpreacA
phV+HOQh21xFzSNZobGURark0EO6MUGqukOaV+/YHxRJluk1T+rUU0Z53cER
PlO2TrXvFOzC2wmStYw3qkLz7vYlizk2mwoLFCXkAdSeeczsrC5lbrZ0z1wz
fciN8sEl9Tl8Zh/jeeR0EYwDO/HdGG0yDHk4yz6FYFfBzqreBW0xOo9w5h/s
8D4tVFUmCxGXB0U8M/tHpdnZUmoQ45r7AFfPSzuo3itx+icS4X1bOn+y/WFk
PDwIyj6Z+jXPiSPfZxizdRkXlgWLGZhLu74xKnGX9WWB4k2EGDU8kV+VUbWe
33ZZXoKwewdO9wp5nG0834XTeU1gkFFTeGgiyrgiLnTUdEvpNlcBZ9JSTfDg
E0VuLh6KWUK+y2/wkalmJxbxPNq0w5aGfdXuoWIHMO3FiFQ7NJAhd2whEQ/m
jnMI0gvFYs6bAgHPzD+qshA1R+VY7IXGVliRoiTHqhIRQBj0xVPxEMBpOnKi
QVH4oOlHjLMuaRnItJCsNyB3yxTtwNr8Rm02pwVNUZlkj2Im0dytvniwJ2lu
LT3CJs5dSZBT75bxcHTWQnpoSY4cVXdhH1oxLCGBYRhaa6sFRk9mcMf+kwtT
CbQ44ksJG/3QRR3dbzG4YVb0KfUShNRH12THB7fu457yjjX+K9hBGnxu9BGO
K6Sp9+FP19uYXqcPt26DoXENO/DY/QW+6IFN07dFTZkWwGPpLiyOT3kaPKFt
l4yJm2pLrgl67GJ+4w9S3licPXpZfTvT+vvcQ0uIxOBiZjX+YS2CYXSjqYyr
oCojlUv/+6Yo0Vx9qJVQr4QNwAVzfZEg91yoUQ3AiAWEqc60wb6DTjeDqTJR
b39zSLxNXqPtXLmUybdyrb/H0l3C04/teWfxVcaXbBKnc2QC3zcDftsv0b09
I8Twh9hoysx1bnUk9jbqXti3yQMs++1au6BY83AfPurMQ8q9x6JS5s9vIQwf
uLyaC8WPJCHjacaiyI5kVYUGyHM0yJN+v4Y61eN7wD0/vQhRFAKfoam0BtT6
LXSMheMaVatDuQkxo39QUCZHUvauo7JXi2xIJi19jHUBbE3Fi+Ryt3HyNdBI
f8A6qs+XLhASNHtyoK6E3dsyYolqsgNUB0KN+7i5KWzE87asYvFP5/QgASWP
BvyynvMH/2ShmQhs3NcLrIKqC6XSESyfrq5ROFSt4F2aaLrp6oL4l27+KW+R
4i+WAb15siXR8qGIsQ1uRYfcIF2F/UL9ce+/84VSKMqY1LIylPhHDBSsE5aK
l5pYemWzyqx4OOjP1kK1tpYRt9lOk12j/SuyBNOglWnpk+8fmSvfbpbErb7A
WZP5bz+FKrwahqX6GFd1AjhRtnpsPdeaJztURhab30xDnRfduGbsVAke9suR
FT4DIS53yXme4xKf81ISxNfQMEV64qIA6BqXY9qvWTpDWqHuhTcfRIx1apL1
27mYbLcdNijVjCS4zzFlPenDpWAzxBmcNKL0hCH+qo2KLtlKMrkCWplCBUwv
pyEUgZ8l0MJr1Ia7CzOqkxRhnoyia7/V0NBqxxPma1eGs2zlzvZnTJ9zAifi
hXHBYYmNHuQ31WVD7pHGusfs+AuRTz4Pb8GZrLrxyoQPOGsPT9GaWOCIuffq
z9VxzC/L8cHFiPc6ErcDwQ2QiWJj4O8Uovl5o7fbHAePs1eU9RvZf93eBdK8
8asodwzv5XK5lbda3qbd0mhxKY4mA9WNwvWPdExrRIfwDuwcDDVkgtYQZ4rp
y5Xo76ngmuRDnRjA+TtWMP3c6VOYfyIsujlP+OeyGysS7cF63Pyzft/a/prA
wOOWiq8I09Os089yQrbKDSsw3nAlvxVj0zQE4dP8L+rw88DtJ96ay+ETHzO0
MdHtpSV45mojm8mw7FPWzFay7je9JEbPmyCvLtnZiI3eJ2PpM+UHkdxuasD0
R1+ec2o/KCHoJNgKJjAh73GbFCqpZo17Lcf5wEUcCefg1LgjLvMWHifrKn0H
1BaAZlkJjxewZLtT1C72bXkvw0+jm657uzpdS4DgtA5djIoKSQpB5VR9zFgj
jEQO6SRcvW8icjppTZxuf7/BDBiLGB81PFyqp3pe9BXHww8yurju5+N3M+hr
Sa4s8450GKXIWCJMVNqsyFanbV8g0/C+lytqusaXoQeFlE2VE//dqupTCE3z
/w03H9dd9I3GHmIeBAYQZudRefO6IcxInhFCziPTuzhjf47R/ys5IJsywtS4
FXYU+0NYB/j4hc9KM2UgWsN9RITFAmYKD0X9aqRyAB2rSJcM43KRtIfwocRS
5BypMmYRA74CifXt6u6jzJsRj1HfsO6B/HxCQ5DElZfmasVRq22ZlfeoJxox
XNPU5kgwePwE1T+/SupGbpCc8YwHIdnC7mB5WhV0NCDk3fHjbOrW8IJ5DvsN
B6tqce4OCmxrdcSNDzgBwo/iRotSEznbF4pJPFIzPPcth+2B1wSe+ydey2pI
LEZgEz31ucgswizR7N2ITwNeRFoZbwKN8jXWFT7Fl/iAwocAmDQ8VeHOlqfK
k2ZmXS2ixuytcYs/ncSz2ho33jSEv9Flg1MwY4BmZWR6+51PY07V8j0YV3qq
05MWcL3MsbMcmFMIx9WhRt8r+iaSM+RgSk3wILkGlwhYRDyc3PSGZy/s/LoT
NBFWV1pUH8QlqawfNHp0BBZsR/k9hYjUtM0XwcgKtqwrbCbkjwXsEIapVX40
lw86bF4Pl/mJM/21p1Jsq0/HQvlP7pP806SCmVOmJptSC12dijenuet1ITaW
mMidYiuR/yBdgLQ5cPJOnE4nK5ttgyYLKZ1N9tSD8t/RDEIgGSqCZYmOmYRJ
1TmEEtZY8TlOVQWGrRiIzCWW9uQAOaUrM7xo8gfVbWS9nDzijRjuC59qjgy0
Kj51vcTHC63s53FDNm7gttqMhxYtJpwWTYfAS3KI7/bDO0rSR01YNBthAVaS
ByMtHEsM1eD9aXGyYXEj9xQKXuXgPHAGddqf837jWbJ+w46K/GYU/kvWk+r2
IKi3f//YpUkqK/hHJV8jDtwT8nmtA+ZW4PNpdziL1VqWnjQVYXEl1hz+uWXe
+f3P9fJJ/v85lzP0RiCfd4Ijh0YfvIrDmILS2tgjNcRbRVZetmx1tZFJVcRO
GCx6eToWDjksIlyKsJiCUnvw6L7hf0xU8hqj+0dUvpFu8Dyvrv9qRDvOvLwo
baifM7IpepZTGPDjdnvcHA2gzgrqDYHNW25XEY0DhDia399QLhk8jEiu1Ot6
rkCWxMWx0AfaXUtaV9IfPKhTlGO0ZJsYjJc7PCRs6T0P7MvlWm5m5Q74sv2d
fF7KfazHlPFSXJSF1ciV15SJeVJyWUxTh+gWW/lWL8YK5rxH/QuQRPRn4wL/
IbceoJ2eQNvM4Iv9ROqLU92ajHy/EScCcI/GPrdCykK9gAL4F8E+Bb3UY4nJ
mbABFX4IyGKtFuff0QFIeMfpdPlCPfX/gctAQ1be+zlZ1ERuIpmZfFqZO8By
BkE+zaUgSZ+b6pInRk4mpdlp6D5CRrYlvrRex5HLS2LMR8mkTdGdfniUnver
OQHyj5vE1YDLTG4N6HBcuZJKEpb2jeZ/jpzawbZV5QKcBBIoiYyFW0D8G3yH
FD45sSzrXscwbVSxoKNCW8A3L53miJQkCG0hpwFp4B5VYn6q5aFMXgLTDVGS
b2SN862p3Sllvo16yXHDfLwL89ARUUsnFqTeokkA/vDQUieNBAWul+LlfAnI
w2UfLreGPSSYUiKUoFgMGYgXwN9W27aMKEKpHzu77tJ96uvTfk2Ph5//y7DZ
jzSXMruI0LVOddinH3x9lcCzEUPcvbUM3G82uVI/+Takzc3YWAOSWplGc2a2
4rJqyXBGYJkzZ21hQBpj5AuPzod6fFXh+szUFUldvuiY/+mZMwaMpFO8eVda
usFfNlySnGFyWDgaOn28nJ8b/xqupOhoiCN1BO+iyvbcCSrz1qeqa/wUoC3e
RA/R3VRlXrZVF8Qhx0/wxqI4JNFMQHdX1mZdgWyGpRHIl+kS7pLNfWnxfip3
y0hbzidLymz6K3rbZG+WzlnnoYwIGkSOW0wkePrROD0atkvABqUq7/m9fhcH
vzXh4/Wb1vqmxH8wUk9qe3de0DNzZXgB7/W5hCow7UMqfWa0jwBffWIzEoQt
cGObFHPBhICzPz36LbJjjItbJjc5jtMkHb8fvEXe7dRw0U1UrUslRaTzVzO4
qsAiwsOhx2NBEoLRJ6GSU9jF/rDYyPuAvYHrrQ9hpKCC+mLOZvYYftrN+6A7
B+gpJirsucdF9+ovRMgncdjGXaywqWzzpz8m9tAffXnY0Fqi+eYCyC6oUvxO
VVyhEMYIDCoYSRH+ZC3Pk9DFocbXhQrNu2rWZBP+BAF9rJK4QlccH6l7HKGH
pfT88vxyVHOeWeV1s5X97yX4RvgRrbfpEjmGb6iCNqQvOPAjidXBI1USRM9r
7AEdnfHywB/BOxKOwnscH5AkCY7J1IjSRGz0xVUYKQxIVYaGabmPBR74SS+7
b5BSiW8t3QIBpIlCElJXBaClgECjU4lH3WRX2uOu9ZV6TUkeTqkJk+G1IFbO
sSsA6mt3S8/RwBeRHs09xUTUF2RpeqFF4csEUZcw2LH4M0pnYTplAFdOqoT/
CkELDwe1anegxKk0gT0+5wLstbKNEKPoHPNWbH6vgE+/OgfokU8tJIvoKUjr
Pib3nObtlcf2o7nnnVyObYyrYzIEWG1TATaj36L8jfEmXqT200bwKlB1S31U
EcUOSvpLWAK2DFBCTVupuIyVAUQoV4ZfTe3kAV8zfM3nI9N4WaXODYgyj+NH
vP6uvYjxyLfH1q0XDKaSRXLkgGj2SxeZWdTlcma5b4cEf3h709lGUuff9AhB
7ROyV6rUhHQFWMZiAZZQxQ9SzZdGugB7SLnyU1VTFotvi9Y07qNmyay4yJdm
CWplU5eSmp3qaA3LmA3NQ2vrWiwezAMdOWLsq6qUPCm7JyYwyM73C2FLY2wY
qEVDLMBB9QFTvLjhfBs0ZgynHG9T/pEWr6DTKnEjKlyL9WMAzuhI/olfeu3J
CWTR4a1kvvG1HxubJv20siei/ggIYPyKj0wm7iKRLxM6M0y/wkmNLceN08uH
PMCTHkRVYjWuU/rNADwLnVM6HqEnl7DGqGsWqpquIFDEsvRKDxAavvqBujqC
qZQerCW0IUJXE4OsDJFIRtQRFcR0vPzjnrxHvgKVI/qwzVtvzkoQ1JzGawcy
/n0udVehn1PJ8nZOEFRpCHehAAQt2U+EGwyhe7M03VjWYWbOUuVg42bMQZ2P
1gkZ4o1ZKrkLkkiTHTf22LpvVs+atRtPXcFbN3UHEwrAOs/m0VF0IRrHB/hr
KphKkE8o0DsarJmlePVbnlI0vNvsOShXbc8oloj+CXr5mHTUOgznPTlBPPwg
5qme4uV7VERo2RNQaDHr2qqxR5GAlIhLzwn+CR/R9TJT7AP/wrhK5KLNfjjA
SeIsml8Dr2t/5yF2ziU1+ptYoaEcQ4u2BEkw5kpN0BJsrs+1vKogepIU/6bG
otSakQmp6/rtjf6h87u8h24l6Lrv82Qcs3YgaHy4NI0KqVkudFBMQ+bQZlnM
alrvDK3l9VZM+cTwGf1FzyS51QkQtSnMQ6OCh0qsixWbMUDL/RuJU4a7uFtN
Wl9VnJbWqVx97VRkkjmxheWX4+HwIiA4/KBDLMwGAE9IsiVQEO37cgn4w1g0
GLfHh3A2OMswrGAHLr8V2gyo570ZGnin31ZnqcKvur2hLyDyIxE/S9a2JNfL
/A7+txkI9hb7+xcjCSxX21pu7SrnM9yaVEOPSyh4h/BPVGPuX9Lq3YC7/b5f
MwjQhIwn0h5ZOvKrjdsOOGqE7JFkORKAz8lBbPgU8uW1XfkHc9x5F+0pFCPh
nTNxIwyodU2wRcLiuXPNIC5itXNUvzvKbQoafnpNK6HfQWAWrmS7xaFb9Jda
qpneZMlNLHgB2+A/HM7CXyK3XW4KuqT/e2kDxxJzOU26qAPZKooP5WrbiiuX
X+6vJ7AP/4bM9MtMhZIH5kNIBil/9Y+UcAuKhjIDLK8t+wbQtHk5cOU+uXjB
MMq100cQJzgtfL1WnWf2hf/jxvBVUyo4l95V/r1iAB99vDwgmlxKN5Dnbags
2vWBnWrhcttl6Wx30BGS1K1S7S0R4jGILEUeF6nX82HN6rQqvlYRZhm8vuOd
JQTtFGvPq0O90UUb+486cvOXKSue/+CxIxc0BXYSwZ3qlIKEGenGzpUz4qY7
gXP+HRGIoSuxZOA7kMAQlcoDUyRxmafMkPfwzYRzHq3pvy0ey/Wha2Fg9m2U
QPIB6tpNSPVG+k6N43610KL6iEDq4aHxKexzXCBjV6fClxgZ3xVdRwdiDHPT
ADyr9qA8uBSzebD3rjvwoce63Hlqykn7sDD/GpL3uUeNxhPtAtqUjmNnkHHy
AHrKOpDWwDZ8S0TYgxGYfhTms64IRp+cwRxSNx3s5xsQAjWHj07i/u70N8Ap
5obyBYjGoWFQV/IJ3g3EmHOXUHf8y5O7ZxGlDITk8krnRrPP8xJS9j3afGlL
/tXroN2kRoV5m3B6Vj3Kg/oSSywhb1neiFcSuxkZIZ/KEqnD/a9LKtL5YbYO
uXZTCFA117F+qYTnEEgZVUQK1MJRfoy3HtUUAxfuuRSFQNrgV8fuLgYb7Jr7
P72Yo0eg4wIFcqFrGjGR559YBuIMBPGwrGJjb42gJTqd7okws24XPW8Wl0xF
c50VJ9BmMTDP0hlE5zpqm6fNC/HSZjhdd+gzL8wlFnIfE6Dz2B1n0M5nYB2C
hiW9H9hEpK9ETxiVPZ6gl/JYBbJbpA/dyUL1s9WcchaaEs8JBdIyDbDGvk2m
ChGkXXLWjN509/DW3kGNHZaQxTWxQmP57g9OY9I4lRUztXbsF970BNXC6ZrO
2PUDi2ZHvzgUOnQEcCMGhnjXhjRRcf8VAS4LwONHm5UKIfT1t15Zlb4l4ZgB
2zJCxC1vs6u1DYHF5GrrnpTBAgN2OqTjFBSh2Hb30SzmFnIB5uh204DlTr9t
Qc1uyADtd9+RGZ2vuG9B/Kws10a1M2GyH2OxGJv7t/wgbb1/b4lv2YfwxiqF
uJVmvPz87ih5piwI8rRm/MmX20pm+LiubFd5p9kf9QbE4uAgOsjKvwO5IN3L
0G0iMRQjO8bA39UIUwyijY4flPzRhNfxXXPH83j8n0sT9P2PowLm6+CxX9o5
rqUl5Jo4SENreJNgSXg3nLmMbkVaH4rCDaE+vshUUTkWMx6oei6KFjpXfGLj
ZuGdGADaT6Q+wezF3udB90wUYOONm9kBpWAQaB5GQxnQz6Le/QnT4H+jEyQe
RfpYZAVOJ3drkGnm4aRoG+x2fNXzSTO+gh7CBmEQ3iXr3fIETs+6r6/GDZHf
YN55mXrMS6arJtxCTfq8S09C+KLsV8Xt9plKzmWi8gE328w9Ip20Yms7LNic
AB+t05YvwCWiPDwjzy3LOiTmEZkN2Bij4i5W27nyMLmKsWC7Ss8gWKdOSHqJ
MP7VykpW+Eviu0d08/T0hmPzT/xNnMQkWsdkITYnN++IOedmIsJOPJ1ZGE4A
Gn8joBnBNgt+knnKmtCFeffoaWd20fn0h9yccwdFODK+N9XLp9ZzhQDCGLGu
kqyTJmOOsWKVC13gbDEzUiULTCoDuYG3cn9k5Nd0McDIXLsEVa92/kgAzUNh
mSnaPyC/rYN2wLNf141HxKg5S2mlAJFUTyeM54VmcPFYbx1uU9mn/MMIYEEo
i4mzQcEuf1KzZE9KEOxcbTKAXXwvByoYZpUg3TDFusgBvzSZBW6PSrCb+Dkn
RGsFk7nflut7lY0e3IVnWoSdSIeVUiPJb24PyelBI0EfR+W7o3+HEi4nfN1j
j8oJAz7JXksSdJymXxDH6FMyVov1AHNmzAtEqsaA5wDgsYYsTsWOg46wxhHx
V2fg9kGGSJzPYgRCYM5d+7xY32US9i/edLNKqNv67v/h5CH3JKiswEuNeJhm
UIljKcB1DQp1haHIOeAnTjNIaOevmflpVbLub7swj191+OI2XtC+2f+3bWHO
Lh/aU1PLuADlwDGWV2whnuriDnXZyfDHpg1k1KRMoz/ZFfL5TU5umsBPe35g
k6S18YGHq+KdTHyKH5sFTGJzX/q2qvc3PO7oVb/MuIvnS1tmD8lAQhVqJDqj
a9GE/kwSUjwqcNyCtqR/DBtcuaxySlTxPZ38S6IBPSNV92wMYnynn8Oe1GS6
LmIDo7s08yVCQ7CLdKbqRie9ldgt6bUNYmi5PHYrpGWDhv8w1luka8jMBQOD
vUM8LynWVqLcdJJP6YAI/9PRobiKGlGc7D5+bNes/rQcF8zx1uruFC1bdw2V
BGfbv+OfnB5Zuz7xv/eOla+kLI7SVfzdtsB25NMYPiNqNvaNt0vVIZj3BjVo
4LOdZfWfaeZPTLz8p72xRIeqXym6jPmQD5O9nQxzzitv4Gmf5IAas0uDqegn
uIzc8SQ/gdLhr65H6dvASh4wuY/4/8uqDPKm9tgWjFbhCSxkgLp6ZN+xvYM7
J6h/fOO583PArH9EMLSQP9sqXHwG6CQjBcswSM2KJbpYDCepzOpSyt9mjlZl
Eju7i8oDygkX2O6+NJ29q93W+TG90EReqjX4N6SbYcvDci2KPzoCqrz61dtq
ZTjcG95Df2B3W9b9j9z22LopvSofwq+hRjmGDgdKIGG7Yv8EggC2vM7Ea1TI
SIfgbIjTt6lUlntcSJ8tp5DglNf/fdE9sbJorq6WnILPZZF/WHobHKEreQv5
LGCUddZQTOc8PmsA0zweDMM4dUnisqRfN1G7U35IL/q4uPXhs6F8/G3FnFPs
aTrJzkz9gCSM7mceYXN6O8KUxsTyETGiie6Fuq29LgErPzNS4mvHIzC4BLYF
Filauq8x+puRfZrToSK8jYFnK/Vkn0QhdYv2RFoKutGKL7w6epCuovrdfmHA
U5G10hvceE56PCvzQfrdFHCoq9mPrcNy0YOs7uR42hdXmeCuYa9nd3rwZrEU
QVymrPbjqyNsJSq39+n6BV46CD3tQuE6LCd+LaA5fbgGb0nkcF5DMIKQF5X4
dDmepoED05kh13Z+bRTUH8sY5y1qlROfcrqykKcNUY4OwSbNR1rpbU1VJGWw
rkEVSauXuBsuok/6of8pIKnQBdHmZH6XgI5jEME9Lb6Eko+YUDL0dkJFGSTD
/wQ7Uat7jN9EpPyrlSOEpbLsQRm1KQIwsSFZWo5NQ6PNJ9Lbiw5a4daRnzA5
m0sxx/psoud1g+3RqXAYXcjqzcK3/Oe/sGXRacyZzTYhQ2h9VcfENGb05lTz
YNCdxXQG1jKGiVnXx2z5EB7yF+3NJ8U29lfg+2viLyk5OaTjXFVqi5kLkYWJ
/SQBlh6WHAevvUCEjaEf5LuDsA9tjWFQxaj+UTe1NPRU9XIyYNgDNp4oJt7A
g9wv/fx8US+3BiEFf+lPBiYszaX3/YpITVLkeVA6VazuIfDUT64NPS6bT8xt
+RCDHGi/K3aAEvSPYa/ZKLDbZUCkSI1qrPGtISaSG0Q8cbw5JNXXwkX4pMTK
ShwilwRnARklXqkV91UA3Lreb7+zo/dJX9QUwh811o2pmMafoo63Dcwrx4ct
CM5sZVLqATxspbtkGmaPQAbXL6m1r2jZIxaz0S7tUm1hDqHR2FRmW+SgneuB
aCB7ZIDjpODbXSaQNut5dxgYowDXfGshcAvXC+BraaRrjWvaAwpkUe5uVbrN
+lETKweA5gVecZGcEqlEp+bRYuUei9v+N06kj4dqhFCflxtIXQDslI8MbPJP
CPIZpWsdVyJ4pa5DhGOwFxfA4FqP2TAgWu8myVNwesWitpr4/q+QYVr0aDIG
bgs5gc0Q4mND6Gkd7R8sBVaEtYtNfzND4R3VmYmxAop5FPF3uUMCUwfil28z
4q+gy+YhwQ4mjQf7ZBslXCvHR8VwoUr9mOps/fIolrctahpCkFK0G9ifFf7s
gEQWhpEIfyJiXq+PkSpJABhN6cUybxs4x6OM4PAy+2U7PC5UsHi7mVreu0Rh
LE83IrSAJwOiLtlwfLP4qkOzNyQPaU5Tk25Mr2sQbKKjuTcqDL1IAyWDtvF8
tcvEyHnnNF7KokP5worn8/cPbTmAigVy5d2MoGnWbrxrYQhhY42vzrj9CQbR
SNxjJ+plxe2MD3ywLKdtpXlCP9yYblxqKS1dWMGgO+FyUvHqF5ag+pVYjOk+
b0lqvwtB60MOdjG5+1EobXSlYkPGT65e+qb/e6x81taIwCk/nz94+zN868dY
4Zro2EMnFIFLp9+7ftzerdKu//Hajgp++S9f5eLvD8MP0Etl8FUHEHfstZnk
PIxIXE2t/Q7M3L1NnqVMNPUNbSQknULUo1J1/qM6P8cLnIJpad4DGPMI4W0V
VJt6h8LluYwSGN6jQcP1CnYNrmmvBJK/T2jICzzsEK407Uv7J7h6g++KmyLG
FEJj5TThWJhWw0fB26PeQw6I+WAhMBDEQTYGc2AS9NZqOTi3U4o906GCvcbL
YRAn0I+ZuH/ngvLxT0mkGKxpJ9feN5oGwHRFn/ryIxNp060PwtWNzTaVgexc
RPLe1Qo0/jmWOD0Pn+5cFwNm682Up6u8fmTOHUhi/oBf4FLMOv15eXT056tr
UHbkB1OrSgMqTU/yyH4d4LE9B0P4lFNbXAp+bj7AW6nY962Sp+xGnKxNtVZy
VPSryOZVoebE7umvfT7AKGCCp/Sh6kiFOD3kWrCKtXeYm2coDsq/I5cPkvmK
0xYo69El4GyGDmMXXetB3rTYj4ntn6jnkt9VRkSCXUs6H7r54Li14zxEVczb
OINMY9kzhYu2z21F40Fga2nN2jDmNEUZqfl2N69+08X9Rgj35SU9Zua9ko7I
nriGGm1X/nDOcquawfOlLh3GK7bVJpiNsU1OgwJ7Pp6NsgbhxK3VIySZ9IcJ
UUudM1aLQ9T900KBV9qZMiZRxNbSwnpZk6ke6+2incALL1GBscKS9ur6siS2
sMAI4zWoyxI4RbS7fhyf3sM/mP4SD3Uvex1op3C1ouFZpOh/nejvq56LaTJq
sQl0ZC/CBS+c3qFc4hg2I/hOMaprbam2H5uxzY5sWyJ67AE1nAquAG3rTRS/
FaW3ajRsV992T0hEUtooYiePDcEgK36qSn9TMM0M9JaA8/EYXekdRcnngfhn
U0+tC0MgvaYX3CsFwjF7yIHN/zcfx82xG21EAbT9GGTTAkbDNOxHGjOcBN7+
uduvv9fIKHLDqyTXqANjpDMjGaYasqCw/iWlgHmi1BUi4cO2h5ZLfErQJVpf
HP8PeYRHsZTVlRokZb40gDaAEKNMeyaU099mUFMKDT6zPdT8xF2kYTtHtoJG
lMCivFU+ahwzvK6ZQ0adkJdtvxKMIWLNIXdIfzunFCMVl/ObZ8QKkTDOZd2j
lUo8PTFLH9QC2A2l8ZiJKHlxayHBcwWlfWCkgBXWauJjcjYOjkNVC0Xz3fFY
q+axJtZR/Jm8vum8Lm1nrouURMv3wL1q8ld0yRl2bIL5Xg220IOLfeJZonCZ
xN67n8s65bfdKOVZBRN32f6R1H5wCUHTzDj7/Vr/Bb3P3Z7CulDyGBxceuWE
j+i3xdA8E3hGbiS0jsVoPP7xj0PKbYd6N41VZBvDfC02Zt5ZQCD7TR4Q00ki
ZGhhjt3p0CyORRMuF3BtKyfczCI4oMhw9CzbMLx+FFYfB54ithsMHlvqVJB6
QHDc+kt4LZKzCmG4DW+KpiTuLD76UoNkcFNGwhKqDjfXugkraCB+97JRR4QP
v3cYQ18SvAcISNw+pnc1Gr/YP94nuCcnan3mAYMQSY4MzUyX+QoeVUGno7sj
wA1d24rqQZsNXNd/J5qoSI6q4e0jqHCM8JroUzlviB3gbcesCzvJK1tzlxzL
dck6k8yZ5etcHMZkuEt8yv3Y/MK8MTinbzTJn7q4bHNGWt6D1LDpZa60+PsR
4wtNUh6Zj5sA43+TVSmwKFfKr17UAPGnUmFVQwo47PTeedRpBB5lXe7SN+ap
uVvSNIJmfhmYeNKrFQRjGtm2GXMIf65kwXFFEy4NVeKvOmai26DQyu0VH79K
UzUn9Jt5WDE7f+LPL0z/U/x6GGjm75luyfgUv7JlPnKbWw9etYEQVt1pEGfU
lYJOc1qYLwgFxPtXL+FDosVLVQzyhmc9v9E8TPjWBhRM5mSkTPBY91FB9Y86
nMaaJAKLdw3NIW2UNFINLidEhYrE6jpopMw5q9aKLgtQYNg9vCyFd+jNeibR
G/VELX9yN8HSJt1gIyVUJaW+o8gq4HjnAng71ZM0hcsIuj6baRKgmE8oDcC0
ubpERyXOy13oWfkPUDw6VR+eNcRs4gadMfVSp8c+k/foFVxivPcIfQy8bNyi
RTzRrExPOHrIdqQQ8ml/i/vwY3LcehPsYl8kpVKAyn6QepuoGx7s5PZZRldV
52BLIFBXjZTR+c2t+KIbhVZWtzBXfEocT0RJ/NFnGhhfIVOyRZs05CZdQKs1
WVWMR+Rb17h0VrbrQvGu+6NhgJ0xZofzTGQsJz9qWiHfmgkLgFfG81h5M/jN
Mvs3JR8AtE4MiiboKTNFAE4umoj4pTrDK+pVETQp5PMoTOmt2krKLeUf9TLn
0DrWHltXfoQF0BsTqNnIiLuehbliy+/S8NG44bmW/5mZZ6tS/crmdPegu7/+
9PJqeHUHDI3ccvjuNSPI5ZOvrDLiudgKpUl3aHMogoYAzPB4fojkLHW8dutC
ekDWBDAAT9GaWV9oVPio9n5mVVCzl0EJD5UphG8JF19Op+nwjKMYKA9EjUBO
aUdwMNAbAr2fn2e9afW9goWVKM0GONq5mJ9vvSlqyueb97zjrmJT3IbSte0/
VHkzMJjr/kUpYCPoDyY/uxUmG5oupWdO6jqxivrfjZAuNdKRRzU43vFoCwWi
HYs3pdbgl56HpURPJxjy9zuGw9rA90xW1+m0cAMIuleV3p6xmf1OcCJCUIeB
F2jP8HhS+xuyFPYyP1vbO6xIOtCMGSIBaq5LpGOJwT2T4g3EuEywTWjkBQBl
OhGrI6IOu04n9SiBBcmkzvlYACt7yUhQXk/a6p26JDMPWsZ16qvU8Zb0kGai
O5h5UABkaR2sLkBx8uo5Gz6lBD27V8NCmS2qo1XjGq8OGi7LAJjchYZBcT/B
CG46r8K80Aay7ox7qBiIOtYwcoxgCf9WiufeKB4Eqoo1GMb7JRZNlGkLkub2
DFmr+aBEiBjPddMKjMfMaSxEnXo4dmlajWM4TKlg8vSwt9H4tjmQ/Tey18bp
itnlZAfSLjLbMfMUwTUUBDoqQ99mK5dNKEauiTJYwF6nDxshiQunRI/CS+pB
EAs7xCy8pS0Y7AL5lKURgm6J+efe5HW4SO6gVAU4bYHv3H2h9dfkxLIyT2/J
vrXHcAJNmTIZLCvrJasbF/9vnjpaeCyY0LnEB1RnJTOsBkEoyQduCkM698ro
kk8K/tFFfBNzNhIOoLOFtukJWWKJiBC9Iir7KHGY6g5HZSRMkV/mtC1WQh3g
4AiN732RoeflprVRmLInZ7Foj1rm4eScQw8NCjipjFQQXYQbUD+9/KXSCsQb
WfTq5FhvjM3u8L8LQeyVRJgXJuPP3kv90m9lWEaEpYB/Tc7lwHjrJ0LJrtco
refuRgsqAR56SPqZDwgdQ6W8F0jsvnNLWeOiFJHYaP6WA4LA1DAq5dF3iiKy
aKcbUcOhBVG4ERl30YtZGL86X4VMy5odJ78LBkhEBS2SwFlr+AbEtMJ3y8Vx
8RLOQUkUYREEUje5DI2/v0nFYsYzyG35gBPkEvBm4t/aEx/8OMcL1Hu+VjG2
rQR2/9Up+PUlGpJYVn8uNuVvB4XWGYOE//dKgmHTcyaSBoQMEu4b13g0LBsw
wL+Jt11HA0Y3WRfkztCgDNnn9c8+WS2zGdAaII3WUzBAedYRm5HUF+7PeAER
VZ9UDvTKXq6ecbGAMnlEJ1bKWiqfVvgHxhDV6BdmZBX1KBa6U9fp4HbGkOKk
H0OWajrSgoYdwuTrQXw6Gok9SJzeupwrIE1b/v/1z/jkqlIGNQoddyVNHVTZ
boZ0xLoerDtjCG3uTE8wFwDU7cNPox7yexs+YcesOYe/qp2A2UXLmaDRJ/HK
iQfhNyD9BK661mlXyt5Dnt5bZzgNYoafGTg2pL1a7tDityGpx5K11CcB9zgO
dbsk9pCMUg7nKAqzavYyecAEqBX1NwyS3Zl3AeUwCdPuErWKM6xbUxCpsqHH
eZJMIX53VwK7PC7/Do3NCthBuL6wy7Xw69WeDeCiD/9oOjEA7amu0PIZfAYt
uBmr+kw/2NaUV8S74AtUXoJq3664sBT3enAzBqgDrQfIamofrEbPCspX11ec
F4CZi/uEn+h/YJL9NJsb+aB+PCsAtLLmDDowegopOdkvFKMb2MbY+AyW9r9j
wEsvMLK1DodNxshzz30rFC1HZJv2nqbpmMEEZwjPHrO8j2i0yBrELVnNUyvF
9JgI3KJtq6WH7CT3PZrJGFpQNqLiOVhMW6s5oQsORjQtuo22NbcV51weNMZE
v0gSNmAnowDMXUHErDzagDTRMJBEt4vB5wlnldSW8HKMw7E0eB+BPBL+fZ97
pMEf+Ai4l1tyBUduU/Iov+KZgfk+Vpf+dlAAma+ytvqeMkd2FeDSrhRUkRzr
oOluuiKeVf0rIhdjVtcz+9dy3m2o0A7tssRp5V6GZWo9wyslXQCaft2uATMJ
F6har1RbbG9ymxadEx/2e5XA5NsWAHN/GtkmHddrWstZWC0gxct1uN9zM3eN
C1tqHy1m8PhYKTPMw/8HIpbJA2gqXybWID4qWClOaDylrCBIeflk7gbMT2XB
L3l4XX0M6Vb+lZpMtHqfwzpObAwWQJDtiufemglBoh+eW3l/vI+uoErMpdz9
eEboL2mcu5ZlnRwt1eW8yulmKcqI61roiBZ59nwADM3DWW9xJ0lzKlttd9gP
My70Eddn8aLEIgGeQBlHt0c2IbG6CwpwUG9Eijw6pPmxQVNaihm2W9eMDfGY
lXJuV63WxyF6uWHzW3xnJgwS+xyu+xqjf9qbDEjzaXpRdgu9PaQbV6N/EmQM
gijBTrKNvRrUob03Llv5Il3aK4l/dzCQUdxO90vd5lFJ4Y4xwzEPju1W+jZj
sqCtjeEQjXTvNIa1Tc6yEmdVGzCgK/2G5YopVZ1YTGlp/JcaTiYNYGnl0U2I
q00kxaP5c7iS3twqzuyZLbC2z0N57Vfel0Q/G3xKAsXyYmN6gj6Jrfm5JanF
4kHKTJo1Co9wHW5zQB/pmq+7F8aTOdRPzmVZ5mJJp0o0TrXPLBtPrOTi9ttc
5jZ/4ARygn9gZpYNHnLe5K5J0LsjDxNcCVKhqARAEokH4Avc/9RtrFTs2Rkr
ERx6zMyVfDmQQyzTgHlaKZMyMr1u+3IPqsbbHJ+4uP4HJtBecPkWnJ5NkCGe
cQMwnHiVbFkEHUnL0uCY5IMWsIVHEgFWurXuy+u1/gBlrwSWyELphDwj+Ig2
t3zbNnGogFnR1DBh7AKhOZzcEyb8gZ1eAopwoPL2c7afFtkrbiQ/OuxloCaG
EsAy2e2WJEZhbgoNfGAC9WCVrhzaqb8UZp3ytIVln1dtZOXujy9QyUvx4xnM
E25SQSGrDDinobmZom9Oycy1ojbVDCRq8G2q2Y3rebXy96UciyRDy0DhReMW
NOIta4tDBMrJ7bl0tsysXxdb1yxb9gEyqRUaf7erbzphOXuU6NJtOoMMmQ7N
XiKtHe3XynmPzPh06INj1hTaeWqdl+DvAq/qEKavUIeO8BUUT3p1H8V9brC8
XaUvLVI36QzF2dIzIrvSYhRiag0YSb5yDO0PFj+GgmEg37zl8OenTBYucO7a
+nF5zqLWiFGJD/2WsywNuDXNmFuozaACisc0lKJ7IxlkpTyAaiAC/Z8eaJlI
Fvb/NcNZpFwwG5tkZ//Oa571cye21N+nzqmiygy7c0UGcK72G2rEDRjrNyvq
nyCws6t52EwZDBZTm+Ayl4C4/8Q1TcsZC6lOe2fDWJgUhC92Ux2RxdYHWNLF
SvT/ckSuHTakVfJuH0b6ECQINNaw2VVnKDteaQnM1RuCg9bi7koQW5R8u2RG
yR+TyXNZATo5tbr7ErHbOz0VYR5UQr8y/wa0IBm26t/48MBHtGRw/4JjRWLs
JK0mSDEtciH23SH6Cg4F0s3dNdiFwx4dcHJOMKuN1dUMLU/tF96XjRb+T8Q9
Gq/mpNxORMUqlfgeV57DI0sQ0eUIRi1ZaT/0Kp92MQ4DwlFVwKQ574BFwYpH
vHlRShcz2zQ2nkelHlPPZcc6MMpSBa2yuXEg1ChrUOH1/86Pn5vdIRGRTxue
WigtoKGyzZG+sTh3EbYIo6IjcOEp2XRes+Ll5aceS8BTkzYPZlOoq+iqa3RE
Jd5i84Ty6vb8gujCTbIwzH47kl4NbymM8pVFE9IqnXmllcBCJoPCtQQq3ymh
7dl9+pl8/45f/Pnme7dB7TeulZ5IIEVimezNJfrofUL6/XNdSp1Wq7wSKQsH
6K+e+rpbyrNgoz8JgD8mN94x6SoLa2q02weMDy9N6hnA3BxUQUG/RIeiBfKE
cNICF7IO6b3rDp53oYNzNhPemYjue2jm8Lw9ePI2raF60e10S0z/MZ7smn4C
aBShqC/bUx9wHACFh6H3HNSicQz6BaEPMrjifX/utrtDqyjgBwGRh1BGuWO/
RRyVy3gtE7iBsH0FjHC8TMxe1JaHzH9AmN0jkKkvh1OuMtNAXpCCpDsL8bG0
2hINoPlNKNeDVwIFI+8jrFlQI046iceD/diSI697fOUFDcw31NtvPGjUm3Ep
IBKUsUqDFAAtcFaVr2l+61nvDj/BcQcob62fjppDkc7WqsfmtUTz9PBCKhJ8
ttP1upA5rCx3EBbz4cArsuhzpPwtBpFLe5XHe+s57im5zDF/ws870sywq6VO
tm4Xh9taNl91AdgVe7pVxX7QNoeGI77Q78A47cJWdBpBBe+ayLfAECGsbJPk
8FBzVALHcf+50rq3DVm5zC9nsr7RSxSUk6DK4WGOXoErnhuHcA+ktSnunTNf
NKujFyVF9IbyIRgHlK0guk9o6MEkzonEdh6PRGHU8lYDcs7qcooMHiQDnpnr
ITNSvtpIDxmOThkRD4MBFd4gN67/RbtZX8XBjtOvZVn621J/3t4MTggesAos
WoV+JMVXezP88IzE9M9dsLVvcjMhwEzJ+MkA4R0E6akSjI67tX1HL3HYy6KI
r44SDO11khsGxp/IvhrAIqfwjj8unpqfDOILP+oLnBa6kqP5PDsj+sEEd4+Q
quVUk/hGCeqJDleDcHPiDlK+EyiDrpOOSKl8Zj8NfHhKz2gYg2FD5KGsncEd
0HHmkTM9VytRTByK5dClCiI1cTpK10I9RP+2cCv1l/0iV3BSdBkZ2KmpXym/
TKumv8RU6RR8y7CWHW5nKewEFfDMMNm5nwLDX6csQQL91Ooj6pgYXOI07ZCv
yXww1HsSvwU3Wvrcm9TBjOh78wjhHqnxHrGZhgGyA9PXCEM4NRKXQjtM3ST7
8E0LJO2SUot2B8GGVE359yFV7rBqF84cz7u2pFSc8y1u1GrXO1jHhtrWfE6I
s/R29gal9L4FMNObYQMN3gKEHUuZ6ZSM3aR6H5oUxSv2Wyqq+B3SAvhrI/GA
tKMjcatGoTf7UcAYlgsUg/NhRpsVtSg0sjngbpBG9sa27emB0YzesS42jdf2
uIbswxS8Hgkzz81wxYj628onGhw7WfIocoHqyPs9ag+2/yQQdhQ2COOlIysm
jjZPo1sUy9ex7H4kypq/jjl1FwAfy+dllVXuhsnwmn+0Z/q9QvKEAOZtTrqW
cQ2ZAgEZcvNuXqyFjXdPzLxM+VoVY+95dt9ysTt8K1j9WNd6kwzW6E2195Yn
C1Yg4pLsMnKuaIFpKKt+f+OmranbGrpWuG3k3VYUVRY3TgR40gXCXrL5k3xA
RpooZ+KJUmYYFkzoP9+xIBphPNuoqHY8MEQKeoccFemoftdGFPysS6lsVTUe
WmujgtsdCjsVOBrAZjA60OZJj3JMUWzm3vHzjjjbM9YO+QfA/QXINQEpzK2+
2c43v4T/L8KF1vFNg4OIpJsYtMtvE866Mep86jroiykn76roEVaomnQm1/Pt
RdXBjufy5tN3PLYd9vbatUX0bHGZVArWgzorotk8ZO0CD+7Vx9y/n+e54y7W
h28+BC9UUv/ncDyL3MVJDjPEP0m52iSUuukrIb57K6tos78UwCJUsMudzhXH
CKNQWsA5ZlaYh48Neby8Pih58PjOPtLV3nN5CIhu9kPeKhVeF4Y/MsphdJPZ
PQm2llA1meCjCcTEsDZzp/JoQgRQXAXExF5pLI68P8nT+k4w1wtdo8fHMR54
4U654+jc9AIDYyF/F1ii5JmEu7PuOuWPSTW//WBfHllO63mKSBuw6Dkmbt4z
JMOfUvNs1sT7mS/yTqRqfDISJIY31/jZ3DNoB1XtH09/5Cf4UoiBBkzqyNe/
leRKOmooBaPLBKlvYn8ROPasl97BJ0sZsfxiOZSBEOGL2oF5PafHq5MlPnwZ
woCVIj9f2UeZm8LkHCIRmYC4oQj2a/XpOoLit3b+u6vqpaw86GzUX/UkLlx9
u5iUVXKFDn0UGS9t6ILdO/UTsHKcwXy2eafb083bKnm58hbyeC+uYvqklv16
bwzCze5o7NFkSFH3M3iJft4Ie6CRvf5f6iVqajbAdE25SJ8sbtve5EZmB108
sJ6OqEb4y1ojlTOlzgkBsFiz+K8u8m9yKfK6NivYOfm2u/ta+NKpV5eJO/FB
mjcYDtOJTS9PlFGVQLn1/+p039itBqfJzX6mEa/mP+MbtSVgmldakZSjFYAI
mO9BhP8z0SoOhtgeZhxsQ30e+OOpqBCQojMVKxlvyW9PYtbHzYzK/caaVBIM
GJpy/5SFE3jobFHhV7EiRiafZIIp66yRvZtx+yc/WR20dHH/x/sdoD0DdXi4
s6rIMYuwREKbMzKUqe4cFCJoOx+/IMhDc51zIAsqdT7KTdDE5usNA0fKD/wv
iAKBKkFz20bBJ2NsVluR93oHH+WUY7U4+MkTW8/8dQ7cvfD3/oXHnpW7dJOw
EE0ozYBx5oZqgStbVYRAIUEtM7NpsSpbtKHwGdCOquBWUcP05lNKydUGgJz1
d3sBJL5dtecnwPrblWsJLy1sol7qYJNV56c5UU0ePO1F/Tg03Y2ocX2pfWaM
zCAZEv0DwCLisqQN+rH0npcO2eJnIEiJx11QoSkdrvVpajehJ1ekATWAVHln
LNv5F0DdyJjp2gQhDV4YAN26BEWD2odls+WNiJ8H36KHiSZOrRTlb0YsxORC
qDx/jIhNBmZ8jE5PeBT5QkbdspSI/+Tz1on4sm3JBDCqBeblVQDstH89w6QU
TP457rCS3xXk9Lbh/AdAmLtYim8CZm6VXUryxzFWNxZhlLfJmui3ej6kGTQC
kOur6wUx8N75KBLtQY3CPrBbm5AqvvHWSsxeXdoP9Hrj5+/0Ho8zsHCh4/6L
QH8h0/6x+neaKYRfkHiYVx6iEbbekoBum+LRKOOsNodvbEGvke2GFTrSy+0a
qyEmdTZUcbCNGhfm/qOvT2sG6CfJqC7aBhMZkKRGwE+u46748/djdpsYR09h
eE6DAQCQIqjybG4ukz9bCzI/HrR4RWdyUcKqws8ZMpKU5qsHsPJNTl2iR2/y
LtIZJoHmDLMCh4LoYbKgRjOyYrKUpAP9bMqbk47IkqPEkWSgl6OaZhqc4hiV
sMnW+xt3Gu4hIbGa9yR/LmdZaQsjdhCWO8VrYNvJMHaHLK3BFrgyZ9zx+erc
g1tQSsXPwzcIo59goAvK3mlUof2z19aRlIYhh8JBsrWA+ZgidZki8ZaQQcWB
PLSS8gNlgJ3yS2+SQ+KzpmxjpJctzVGZqUW45/990k9ZrJmGD3AQz68mNbaD
5sJktolX72vJ0Gpf12uJO9hrwN4pIQlgTuw6m3j07oC8ehIkLBC53lSaWkJD
fThiICz2KyAVWRFL328wpANgHR0DkamJFjSCkdyeSPiRTWxFOzEuUkk+rcXy
XQaDT3REHB5Ychp4n3EAuwdfUymmdZmpjHQtKB2X3Uq7h9i3KWgISTWht53r
eXdKgQ/WgywYlPLUB59FIz7caXAim8Wy/uOBpbDwilBFIEDt8rl0hhH6o8sR
eeGuvCxLTCjePfNYJaX5iYj0sBddnzqC+2FgZejqtbCtYWPdNXDS+17psyrR
JrDrOWYgfkU7NQ7sPn8pgDUTvoK1rodNu61MEx2JQ0wFYZawSvV15P3NIqcA
nSPkkabsOpYZR4ocH4brvJ4e4A83msnZLVzT2FT3/fpEgsOeZAvhpflAwm/j
6Kii7A1+VK6NvjswnNTD8ZmVt57XFkcJ+zLftOnt3frKV25FUR18aUiXslAk
IvI5YeVvgy4AGuUKDAk41m+3AQwc7Mpo47go1IJmaKXNf9mlTnRW36cJTIZA
zGo3LlalFbnAaDCqGdrVUdwolg/1Ojg1WG6VL4TZKidZrWnn9lY780gFkANh
fVpH9K/ae33Bmyj8zvNAubsJW054dh+QZMYtSiNV/JwLn87lw8dQQ0/MyExc
YGsO+GSG/ysRNYh8cQ4R23ipVZPGmNi5QYpftk57DSpFBjvCbyrJWMknnONy
rNbk42ficM896ttL1pGGQKZQ+1KWEvG8sv8dnhQ1rIDBvRxQL0MgAtFLUmo+
jagc4Ri0pYOOtKNHpqTLvNUpKspkWpVjqaVtZI+O7yrJZ+5136XJIbYqsOid
xYMN44JzxAbdEscRee+XwDr52HbD5oUuSu8VpygYBI78JkvOpruSrouzPShv
emDL/yr4De/JagssdEtTWVEI7adbZDndBWtfLgjdE1tmmEZqkD1jo0nRI0P9
HZhNfBdKUSl0+3fILjRTT2jHs7CWLOzLqpsm0wf5KUkDEht7fP9GIsnIJsUJ
EVrCZ82tGONn+VmyKaHeSJqH7tHEvR+xnsobyfVTo9/IR1QO7LzSlwEgjqXf
QDfrcewtHy6LfcyX9u5yqirnDc5OM0RUdoPwrnbyjf8yfNxUPAjcAVJ2IDff
RGrywCBxaOfmCkoHUC7/SXLbn6alCLTXaCZBgUFeAuy7YuQ6NGshgVtr0i85
rNG43NXMCtbN/sAzw/aGAJeepwwt0Pgc8Ll9SzzXgiZroehk75VaX4XU5+hj
AijqEsjZ35tRW9MolDpx6KZfzg4z1WcjIur+IdjKo+wW9CwNRbv6pCLrubeK
xy5ykb3UH5v8aAgHcUYp8ajdfz/AyAPSblDOzuxSDDmgb2Tp0u53000wdtRH
7dW0ZQovIqiWvzSfufdl7QxzB/3O9q2YXDVfCHyK3Lk22mXU9hcWE+tJAOLE
ynt6QEZyZfDdjvX76vMQxGlvhbf5XifMOYbJN1z1HJWp0EmAJO0iiTmrUCiK
m8sdE9tIl27G82iHgPQ4xtj0SVbfQQ3WFzCtIS5Z+fP1y8pFpcl++3na0VKt
/p8kad2EJomqp0+CkfbEcJAjp3I5JPbanAZWmEAYBJBX6nuAeIP9T9ZUkUx9
oA36QWpixf0ggVfoRHML8Hf7W280EMh2ZUsh8TWKaHE3SUIagREDltzNnJTV
lFEIyX2aCT36ekwjVHt2BTeiFOlr6Lpmqj0YWHZWPKZiPq8bZLB9vlrFHkBk
U98unP3Xioth+ujkVIa67S2f6H94bYwMQIoDn4cYc9tCDwstD8/nwevKbDSu
LOvGiE2SuuLotYqGy4vNQP7TrGGB0rQVNFbwGGkCJpXkA2HEgr8+9pLlpQnn
+rIdQu4NwQEWtFeVhEnO0DqQrEkP2mE5LqLArWUce3FbuLrCRnWOyCon97q6
i5FFP7GIpTsJFk1U2mCrXS0tMEa96AN3mKs3PDa1ziGvUspuWj/ydkSZm4DD
T78qsJZNaLOQ+k+1Kn7J97spoMQmn1954fKxfU1C50F3Fd5o21uYCY38CAtC
rIATSbjMq/NQAzt2ovFqFwXUkk3PCiZXND6E/JItUmq6TV5gFJdBekhIWDoS
OOptPRkw41A9/i5GHD5ydRjdXn7jofF9RZjTrFeczWrRmLetefI0bYXAkAVm
WjXb4KsLBUbZvmMZ9IuNMSvkx7MBo/GEwySQdnX5m7D816PKWfHcnMExhVxO
UBOUxYZog2wjKoOawqhbJgLnYE9l/LqotXb2DINHt8HMFTxONFtK+tEyrOWK
ApTtUVMEQeBq/AoBo7IOHsTQjh9JbzBju5gSKDfrQg/tGA6k1Dyo3zcrRKdI
k2/Y1lz7YykVMacczaqFw7g2EcaJBMg9WOy90lvGN142MAdsf8QUiaQILrkF
Q9S6tE50xXYMxyGFuGlFUqmWJr/5taOZR5XkDIB3z+q2XEw+z9MN1sgsSfC6
pBqj/wP0poHCukiPqIcnzNm/6vXuNoIdjCkxGC8q73V08hTW+JdcziPAZi/w
fWeyRZOALSqTS19dWUeNDbRuEoh0/sWapxEYjlYiST5CLeO3mOTZOShf+o8i
ONhMA3F9b5VnYsrfP9C6qZ0cJow9OAge8KNJs7p3wBfFaBPfZgap1gErU3MI
e+z/N/LJYQEEKyFxmOr5FA/4ERxeTAilqCqaQVWIXHb+5U178u8CQ146XuJF
O254ciudTffZHD85cuFXLJXuYL0sV5S3j90uPIEpsAYXvMz1lcNSLKBjks+y
WS7Wlf47xJnfSgE574lQwVFPDWFgMQzDCk8af6znU8vNTbdQRoLfqhl74V4d
hESbuF6oatiuwL+QUcMeKDearOmek34lm8sXcy6MWshN5FyzjsI5QkJEIPXw
UuWjKl1FAI/z63dZ1L6PSDlE4luWzxsYzfoqO9tvpCktf5hpQ6SmCqH35bp8
Sk3JKpVjy+1RqMKIc4qhGbAg70a3kROEDCCjVIRAS1VXmOADLMlbayU/1YZz
BlRkZWRdoZcLY76Q/KMrJp7BISciVqQlOdBNSb+ITgAUq8zoh3itGALMUIG2
z5ikmSPnmqiS3uD+G2xk9LXk+GztMqUkQLxmp0bRKvJmol5bjdvTcDDDUbBH
dW8N6HVfMYAJGCMv/tKnikHLXBm9KeE3mojaS+6ycavG+e4E+XJ3gS1Qn4B0
MIasY8hirSUx2cNIfPC9/N5zPmEn8FRP7sW3SktALcOWGBEtD28A37VZoK/L
uUko8YmtCrzP8xE0fXZOV8/OmOCZ/QIbAwmgGZd0TGxGmeE3pj9rbyj7ndCY
gHnHU7GV+GI29AVhB70pj2gOVFxUHIRoekSGRBOe1X7OLnEfhiFlh3vtjPcR
qg1YZ7YsxmKA9piTr486dYPh62Pbg3dEctzdHjUdF5QlEdZsB59KRaTNZ0VQ
jrxX7OVvUtBq71JS5um9nmgpwua7YhypD/4ezHQ4ojzdeViucxQ4gAYwPqWy
T/NsLGBCsH3RxQlDUPYQp3JwXlhANmn57A2FFFuRZur9LlyQ8wK7iANVdO8p
nw50AVSM9B6Z7A2cLl8PQPlNlFUFHtqdPCGWWFMPeJQQA1QRfqU2aKVOmgQQ
aV02Kt8nVJJ2xxDdLBCicCjd66JRXOQqPvox8lRWe1k+L+ghKbzvxY2WIbQ0
L44srCHXlMkYy/PJbNNJNKVg+R8xORuStriO1dVj7RoUESYfJI+1f3R+mr6R
a71kRlwuwZQecf1l9pFPCY3eQjLuWIlUMeqEiNJoottjmPHclkaue9szWSaA
xSL6C/hNUtwcpsefaG+UxoaEPZhvDac3huyzfaI+KhQRURIu6jyFlXF6JXq4
HRrFg+D40gLbuTtI0flNS8PCwPf2b3MK/0icXTE9Qdo3zCw4pGBDJXqrQib8
B90FmEMiDxRLpke7iCcZ+IEICY0P5sXLe5YJlBGx1RZSCEBqtkXYAEzhiJWu
f7It/aw7zd9GB0ottaRgr1a9IYqMfP/XytpNBY+9IokpU0VBWxu83x8eVNnp
KQ3J37f0D3xg46QVb76HBC0Pencjc0FZVzZ8G/BLdrqE8deh5zgU98FdrUXH
7WH2zeERoWIYawYDuUbbhYvipYkJB2ZaOsQEo/hsuho02D7QlevUPobzToLd
JCxLTwtoei6cLXMjXlgz2MHzKQuYSqEm9/5+/3K6BQcAGoB82EfdGW4JQm7d
3yrb/t3bnpaJfdl2M2H9F+Jy8KREapiNxtdJHNLTeFOn4Q7dhv/Cyd2CBcUr
zS5LCXKDcEDyrF7DVUBE3VkYcsq8YxHX1/ipQC0/njBuELLGY5QprANGm9aY
rxnqIPaDH2x9/vN2ROFxvqx24N2fcwd6vfIv6Ji+FuLRA+5CkrU2Hz2d+DJ2
j6Eb6DcSl3TMKQYx99+66uiqI3cNLQGH7+nnZXyFQNMill3VBjgAz1jFMy5u
I8MF5KGdXShR68v3c2tVJ37OvLbUbWpxaCnso5YVzeXNZYddzEly/7GCBuQS
qYgDHDuAoN6u1wHbgK4td+J0tYKAoJzYUtEcQtYMbiXne/5WR0Rj8DgOS8l9
EGhU9uij/I5rem8wOD8gIw7dhezPjctUZ0QKRUpMvXW994qn+TGoa17CnwXO
1pYKSsU3S20wrjtMCxQGBmfUIQVpFtK3eZumyiUxueyIk1rIvNcJRYwItzmi
9bZZ9fu/fEE7nIcfP+9T8a6FoN4lnHampPUjeZp1n9HuUiMcqP0bXukRXqr2
zGYEtGl3qMmFiJwJTEAV0/TeDNQRDEBNbqbcnNiX4AlwHrq9Laib9qoSxRK2
n8lQ4fCZ1v8HHdDe8yAWHammrlgJXTZ+iaAUf7v4Q9mghac97C1gym0nx3dS
n2KpXxVN08KGrsJHS0YtGMs8JLi9V3WwOmPo1OAXZj7cX00byOAShKZbvcgO
rtzn1ohP/1li2UTl8LSlh5PMaf697GFrIWWZjmXjKmxcxey+WuIY8tcey24K
jRsxMi3MThKVeKAjYoCprhNmzDE5X1aptAwVr361fC3kht0c/Vluj6UZSq7o
+5xP668tl1wqDqNHHaNlF3OBnd40EJi8qszfaWlkobIJtVHcTPmEz8WJmeCr
6/jCn/3IfXnzANL3o52UMi/cqVeHkLJ81z7x0udbG7PdXp/j43k2zhSx8dAw
h10oWpC4sv0pLdk1dU/K16wapEzVUqXSOHJjvmxvdOZlzx4xj7pgFlU8Lltw
IAQUQjJrLKawypNNykp89vNyl56GMjuHOYInATtfeTguoUp8vXw/T5OwhU81
e2hbnRFL6AsLTMR7ViV3QVCCHhZt/11a9TVVmJib0WQJmtwp0iDfFcN0kKJN
+FN/HQrUcUv950ujWL77fjLVZ7xPC6DhhAOP8RWq8gCms9iOs3zmuIi54l81
nzlbHQZPGXMz0XbP1wiyNuBM9Z1ZVH0yd5wmoAKs4Umk7czWpxDxcUKEjU4g
Wd1rLojFXPVq8MZkT0Y/SRN1Ho8BOKGCQk6NntZbHLpcaxNXldzrR/6jb+FV
uaIagwiHWZNxUPi7GlPqXuzux7woBibIKXVvbVsfJ0pNBC1sw6uh2ZHf65Gz
bqrb2hLv9ZBxBR5oTVg5PtgK4WAMJw9GVlZvZ9BCen6P+J/I423m5fkJdEk2
Fh8Mh7SgS00D1zrlsizALscHsAKDxRHU+P6nbXAXb/oBvzWl4p5LnEiu6EJo
pR7MT1gSIz9XggMoTO91XZjdQrE4myXLhOVusnSqFaK/bgp/5MDp+waseZ40
1Gal1q0IvvQ6u02YBA4FHWU7eHecIpR01TZ97m1wnh7IRBwsDNjmZcacqemX
BQlP1g3BBnz73NlW9lm+CVkmGpMDm7HnK2TtrdBHrzXgI+aT1nNs3b+qKatq
kGRkv+elzK3NXXyu2W3PScQSuz+H3H7fVbCAS2ybXV6esIleI85OayGVbc1U
kewUUCZjUHvMYsoQNbSJF0+AsSW/ATNK4mrAxw4hP9trzemRbQc+GCM0lHP4
+eSjIR2uOFk8zj/SyGvYneRi6+R/Lv5R8DYTFNtai4GKqZfAL3vScUkR9a4N
qyOA1UtVcOP+7mGu+JjX8AEH/Oq6SaY+BD2lJbtrSTjXMuWNEtJSglQg5ZJB
DiNHl4lSk2bDuryLg+scKy7LpQ/nyPmIf3Lw37ilbLMpmewaqQM1GS9VPZoK
yAAAm05AniZ0io1WcTlNKTrpjmYb4g29dcpVXzEZmnd+2ByM9qb2G7UhHwNS
ulWqPJb+hg+oY6Q42IjCGHpqfLARQ4yqKdzoNoQCGV19yzfPYe6kqpVRrvsZ
PaZyhNNhxFQZmZKJP+tuVS6DtE9Ppgj4HgO7NEThfUeHjzO+sA9PSvAtNdTa
NwScgDzZqmvvxE03/W/3rW2IfFhFfUqjzF0xTBpLSp7xAXs7/YEpiQ6x4J51
/nALHy4ioeWTb2DEm4rWrwJFSVc7WmklebhC0I/HqLeOCprYiR17MYJcW8Ak
ZsYBDpBRiHqQVcV8cODDVvaig8XRXxBHGiJ1z94O8t1WVxeVRIuhuIjwJR38
KRWNCzS/uzZ6uX1GLAx1D1SAKxd1NbKGLVYrNK44Fc66kHThU6NUX/+zR3vJ
MTvUv/ghrYKddMADw0j31/YnVzs0WmXcXCrIb9JHd1PJSlGE4JoFaVGb4h8w
WMOhkPbJdBzk+xax5EHWAqEWl/RCvroUEYJRLhv73HiipBH50CRul44A4UFQ
y5Xh2oYsEuGf+SioQRvnPj8D5JTzSOwIHybVS/C7gRcusyw9ydTEcWCOSvVN
XKG0xTHnPEsX+YlTbxXgTrx+Wy959jMyybjxj7Dnv5ACyKUSiM4dww9d5RNf
AUp9SlzufMswr9Yk3L0MeAiBe2jAzn89J1z7roc8ocjICvOeFh3RDGkkYo/h
dshAsZEmnYuoq5kUosLn+3kaPyZO1iU+fkcDrAkXHJjjoglzlRifsvhZSs7r
uP+46RyAr+t1nk3BZ86GNh4NsGSUqTaaoyjtK4h3K4HN6mT3vDZ0OGmYNMF4
8T5M/VRw+WU38XxOgBJv7R8eagir430W5e0tIJMwTDHmUiJO0Dr6uz5rwKiX
yh0c7rZzEIuMCHhIglB10th7jto94VaBlLm1h5ixp3rlcwYobyfScWCp3Uof
LqlURVZOiWEvcWaPy6cgt6UnVCL292V+hrzRC3JzPj7XGoVtTpwOWRy+ayDo
I/j8XfZ1rICNUTq1+36giFOm6Gn7z24nC64D5DhBfEcmHH91zK75Mz2eumrS
TA5I93XEP9z3XT0fRjp05nPAPDUdh9bCscwYPIjj+ACOYmmp3XfOw4DBWs+X
MQnD4G1JhBUkQJgw3IHMwkmW29Slts1uKOqxqGQjXDpXjX1jwVL4DpzgF3zf
no7VA6A0QzrYBo8ffDcUs8Wrvr+E5zEE20cQnlTL9Ez1j+R1AhO+BcAsbXmj
MYy0Ent7j/UvUEcAkOYm3vbHEcHXoCrbRgPdqW0WGfTDenpja3rWBCnD2Yw6
ulnLB4PrqdMVK9+kThhcBKj+R1f/7aWF+q97EzmQ8+ry3bK1VMO/4JPyLoJq
svx7p3BfMFwEhvxKvW6+gHdG8hYwSzbqBpUZDzlhpCu/qEM9F9OaTcjEpJhX
7QmFkpR1v12Q3kTMApr2wypL5nDzh/kmDofxLJw13M/GZ/l7Ok6a5qMxyMi/
G4uWYqv8Eg1YS52tbBxe9I2p4Rja9eyCiQ0KOOGqTVvdVtVwm3vKpLjrx0tG
SycJKbdjeSSeQy+n3oDNMIEJFOKN+LEYgI0HEkgHgDo1M422FA8iyi6ZQr9d
w2zxl7Z/zZmACenvWhz2fc4vhTPI4+pcVy+p22SuH9CxsKq+5swx5iqzR9qU
oIPbH4z0kIeFd4V2gMCNSUBxRPDuglHqU3Mj6pg2IwWPSmXeSjat7Eggiywl
px/TDn5yMkbXABW6200WCWxl/wUlI+8ZNDWTivTTRS9Z7M4GOSUNSaWuxFIM
uYER3UvyxWEOVWrvQ42nVQJPz4Sr71sZMAOtLiRhEpQUpygd9+3SLhb3c0Qq
QNKEaSA0KKEA6m+GC1EGT8mTD2qICECBWQXcVwXsT0n9ZXTnRu6cRTM4UzIt
RgyKsZYt9q7DOPDbU8W6DTw4C5+d4mwrHFJneXMAajiK1cOs+8nkNqGkTgsh
Lx7SafpM4R/bSiNZvGPalE6NLF0kZxdhhgNd+/bNWehK4sqHKCiZr1iEos4Z
ZICKiXNLHfntVSIc6Nq2VSdV0qAyhAl553JssCCJh6celK996RGR6yrHl3/t
SL+aDoCD/lztX2W4+N7o33z4Eanlr0G06/Dw9TJ0InQvzV5Zj0CrCsir/jyR
YKv9H4wa353ElwRIj7sh3fgbBgnioQOwDYZ3G89Or6jNiJdjioglihSwhcuC
GolkJGon+z6vLwfyz/6iXgeM3sORTj5hxb/CJjHs9dAEcriFZI3tLtbhnTRV
mPDretPGb4Js6sLJ8MHilIwzQt+oxzBpoA3Qn3BS/7BKQnETKpgb7orTu0mi
QI8/As4G1Ty9JdweDbuTNKtUkqbaQgQoB9ZfS6r9PwBJ4LNKCVF8L6HOGRXd
rgo4hm1rk/mWHanhzEzh2OWFS19dWD17hXdaRkCnAcNHV6LocRs3qe5WPGRT
2uIRWcBG2P3dYPcGkZ4rXYEO8RTdjFtj0Bt2pCkLWBe2fIrxx+2/TDaAcZSu
KaHagsWempfJEyj0Vh/b2ZCkbcU2NdnUnC/6WqjG+mi7zISr/SPjaMa/k1B2
5VbEUGP/l/d2UhmDWo8xUlK1oGqP2OomXrMl5WWdsAO0KX8WvOV115bm6Zrs
imbmH96emlF02tCWxLF6kyOOJjpGVjBBu7GE7Iah+fi2yI6QYITqR0Hv/V0t
Yb61wYrQDqPP/n/za1SAI6o0SlDZ+x2J/dp7sY3tXYeibV3lYybseENSAIyt
LWe2FVzw/ZI5PZnb3aa7Yxl0aev0Ed6WkplRfHljl60Xa5fBGDgILvd68qUT
Ub15p0c+oraI1y8hFP0hsycClCa1si0QBVriJ0tAIS6mW5B5LCTSacP55VqX
Bosvf5zt8ZWGFsT6cvgavBtJHQ8sc1t/Iw41m872cXckNXoniTjyEG1AgJ/5
MAroCT1WIDYFpug+7wworksjLBvo5SMcIQ5W47GfQtjG+zkttijpTIh4GxTR
gzhjjU3A2UBMbh/qVU2BKIfVnRiJNbER25K/KefYb+8QLk7Atayn4ZBl78jz
iqeE4yEo5vEvLcaDf1b0Dz/8UzMfhc25eduQD2uG8hZ2hsgElcNT5mxHrt/L
OTXgC3ah1/NSZVSI1P55ji9uCPLcFU6oxkcPIm/kkfAsowlyFHNjj9zMOu76
qDL/oFXOvrXZ5CD42GHyFAd6rz5FYLuEpkjZuhGWkyXjIubKuw3zaJbReZPe
8JoQqxrGX/jLSXaNstfyga4+qiijsTAPG5KkgxfQayXDh84LJ8ov6DuwWwbX
TsqGd9dD+SsK1hv1zkmKyiCxIhNuZhlhNi2aAGxapXPsR+x3LIVqLqXE3vyH
mpsnUOi8FN4d/tZf1b05wrETBTx+9vMjMg4HoBb6blPj+3s+wUR/fBgz+1fw
y/fgRhDwHwpy0kM8bcgFC08qjAzfN0zIfkmemy3s+dgiDRlRaKkKYGubxt+j
F9JQCFADglSU3vl+CvP5awyRgctF3mDO7Olc48A42YMXR9eQsgvSgWPTNSMm
sP/CCdAaGVdyFcdQL9BmZguHdYK13WV+oCj8Q7cGka7qtlQ7qA7T3NY+wFpL
zrlBtHcgyqF6Abx+R2n0WVPrAwZAAcatD5VJtwHA8XXmsXJJpg0txujLLTjl
dI2xlhzUaOV0aY4c16R8oYdm/Nban7p2pk8DsCJbwSxXX074N2uiC+1xmZ7A
8KDyhgdCvQ0DyGPwYTwYuVQErvCiIgreiQwf9gfKpNTgjPRjFY2DkfteKniP
X0I/EeW5J+uRcPJUddHOawePTmR2wPXLY6TStRZIBhD3BE6LryUHzCE0zH58
aM5Lm6XIsgA0vfuqxnRWGj3335Crr5dZ0YAgPQpt+0wlsAGGj71mCvlA6+08
ozEeBbh4I/q3bn25k71OJUt792GdZb7cG/Xnwu93E7DBarFGzQ89s0kKeDvm
/soVwM5YRQ5+e2feqHPP7xz5SQ+G3++rGYGF0A03/mePBqAOU4XYb5JEOzQs
BRLh9hCdcki+dTrIrPR2kaKOrelc/rkO5RB15Z4AcyGI9DCAa9MhZ3TddPCv
tENpMK72QYdkq0ohJSIizVADYcctxV9T+542uJvnfNIjYfPk5yk9Dtyh4w1T
rSwplEU3Gumy0Qg4BZHuF3/nLYJhI9mrIfmvWH+B+EmE9nz55NYLqt2t/LZA
HrlFP1YheLyjsIExt/Ku2mMdG3lanh0m+dPtVasN9j22WDKyemDnzfbFT9sw
OWnxSXt6zUmMkK38/z0CVQuNoMiSXgUh3KZmchpQ4zDlQMnNFCCszTfHiv2P
n2XFDG8ubiBuPNKla3fVBEl/+Wwn0I+fLb7jU2Wb4YgQ/Yoxhd1YfqZODi9Q
QMvrfxkSYMm1a//YPzQZmEXKYAN3ib3k8Y2xm1RRLXQfvL+CNA6AN2Oyw61r
iL/f8XGeLnpDCPOjyK+82EShE9iSXc7289jL9EEFDJPCpNSchHtI+6Dp8HGR
dVseIsjtuOkvk1OMkqFkvSR+Jp13kGDFxfcsy/qm1++uISHtaVc+K7J3KA9W
tsNprggR2c3oQ+fbwUOsrcHC9VqELN+R7hm5aCCEIiWNA53H7a2N4ohReyq4
b0tMCApOiT9sJ5SC44qSiu8vwb3uGgt4W5dWAKaqOfcwj2yPVMdHCiDCZ4Gq
xdpOp/pDqxLDnNJIoY7Os6PckzGB2G3Y5DL5sDvc83Fn5haBQqrNwaQICWhV
qkv7/7lWTAB/ihdXbFM/gFomNOlHQVaWB5VNBL3fSqpNUum2Q6bw7Ke0kkBF
8WCghR6bq3aR3bz19LnrwGAG9skuBlj+gnIVnesl1AteKPBuwqZmRTw4+3Cy
mqzOYKzyWwIqF015j5V1t8T6CTDywlPDH/F6Mq7LPXnZ8iyVHyOImk1rznPz
Kgso3DEnE64D9W3WiZP+G74o1pF6faZRAWZS311OdVVzzRATXwogpetPa+J3
TX919w+8fFNJrAgz5AGAwF4Zmrf+Bw/jnAqWBpZ5dWC7AS1Yn98uAq+WGmf5
EqGKThoO7WdbTAhR0FX/jJ0HgL3RV5bGkJWdjYdM/SWg2tLTpdV4tiwyxqhG
9NiAc/Px4Tr2iLfyTcLyLgv6M8MhxsqPs6WHbTG7q7JHJoJrTwlBSKJwxWy3
vOq3aiGOvENWotdUXhzdOnOu+cFRJo1/DSJ+bYvwpoMJDxrw1tazj+4Zh4kh
9rnLDlHHWa4uOLh/50WksXrOfvhEqRrUkqpQO10OOKHw0qUjzYMKmeKpnawp
LrZ/V2Av9v7BqVwD9Tzh2D6Y8zJXSM027nUengnk9hSCarLlBj55dfUKN2TP
0ysNDmy9EESuN8lS08nxv3CZgYdG4JKcrPbP7DE31I2w/7SWGloukbKYtCGp
M57cN4SCXn4Pg2a0kLpfKVo91MWFqGCaF8/QKu+6zBcEKeRSAgELVs3KM7YJ
s8lnnJSxjea0pB+Z9qaUmDznIQJMhO7suhk6ykU76F/n9ZBOiduhXCCwTl7V
Ex0DCCcF9P5oa0TrZ844dCnN3Dh8fgP1UrLyOE+Zhja9zBUysIpBctGFC5Ju
UGsLD4gFA3qvX8V+3MlBFT0GCPuRQcxjpIyJJex/wLZN+xVu/xey9BWlKXvv
eiCzINaT1NwlEYflZoOgWiSNpmtYJ5IxxA94nIlIgw+AF2csHQMoNoj6+1g4
jh649slxp+lRPDCWaNx1UxKThHFC7fB2tBumDkeflYxHpSXFSxAGkca0iHn2
5Xk6COSVnsfvJ6vujBV6eVC1uJoFSoUsisVx+vD/jG+Am1Nv6xz9O1FbFGiv
k8JGqBc5mhg/d7fAujBSZwiKyJ5Q20h06RjbqW41tbGfPqTRzxzt8mJal1HF
BJqbVYRnkKsFucJSQO0er15Kx7kjpm2d4pq/pSbeIvoJG5yNRdV0dfzwyt9H
8pEw0Lo5rxIRZVmMO28g/UUgy9yD2QeZg426mUvCbDlBwi40KD87if7coVXz
pMDg+X+ey5SwRiIjZKDjlLrZxrcE7uG4JPnESOLPWhfxPCg9L0fOxJ7wVf7W
sBA2EpqOihgHTGEviH4TYS88s8CAmXXZHU3gm/WMSgk5GBY2I9UQwVryUo/m
v9SMDtcrRTe6zuPtTLr+Py2QABXFXSoCxtgjCKSUqLtq1CCmLSoeebETKFTh
meyV+Ph4pyj2ni3yvxmUv+NhLc+LDFy0A3kXd3VOL8qW8ehFQwkGH1ZEXPUh
tmxQHQ+eD1ioHtopKMNmaGC1MZGwDXKzEgJ5LYE3AduSkV8Tg+lBg/0Db0ve
ubJJ39/VJ/tforLLg2muFzCcsGK2RqbfBa+ydX759ihMXo+0xmNbMKl+HQ6z
3f39m2keoYllLrZYQa8Balz5NYmdGKETEdCLgdP7yhIoNyxyqERAjfSPePLu
goPJHZJrMEsRl1Zart//LJndyy5dDc6nNGD/STYd5TabUZqnPQsVptlXN1Dg
u3F1vFsP1WpTGH/NNxKUEZ9/m+D/5TsSwgyn6wmK60Bxi3K2IqF16YPs5GwT
pTvsRADNZiMg1rW8deWxyzelCfHEY4tR946VTHPHvgVE5zz7VetdpJQhcRLV
QsuHy25pwUb81It9JLXjz508nTy5a6wBiM9bIC9tD655AmcE4HCcBf34MvTE
iUafrPY7XrKTnS2vyrhR8JYWA3FH5rLlYDJ+Nk2HKzeHcZeOMIY5ULBbvbb9
s4cucs+85hU73QsR8XpU/jU2BfyICenMCg28h+5yKZbI67cfuEyG404qYiRn
R5Cj8S0vXuh90VwmSSy0TLh5mvblJuXXHSWZ3l3OJ2jFscUEdmilmuFCHRfY
DJNrf6NmuL9GPThzXm8mlH+/gWB8RLKprEDVmcCV0tvRfteI5KsnKlOOp0Y+
yI2pCLPXK3iwlZhzmViIKqP465D3w28FhtPl+CWT+GReiI4/50wbqgF4xhrR
dXZysZKj0hQXZsKlYHOnUo/4UgWC8yzVppCkFUqwo/vn8Eg2M1FN2N0VY7ZE
MErD/IFpvkLVlG7rxQwsr4oo/qHW54bwRaMoOA5bB1/sVNo+9alhMdmox8ud
z0PzV06sBopnoa4n25m7C779jUCRQccreaVNZ1+aZGucinILxJazpHi0X6jF
3tEsvMZva4beinyAtoZYWn1NFYmI/c/BtyIGStJtfLibHwoDZHWI97XXPrr6
iHp3CPSdOob9BrLRe83LgNIOHCf9AHkLUVGsQ8tTQaEIKnZH2E6KJFlvqAsq
IoUnwzwE+yZfhp9BnEqRh1x2QugFCoils/BoYq4cFRdl8ovUNiJuqN3sqPIz
f8Fqkjm0iLwl4/Hz5U/BGhoTA9idwfB+ef3jEc8hMSvfVvsfv+o/21mFYm9r
qbUrCyDSFpE8yTeDRzjEkEkqxIK7l//SLPNMi+hhG+cx3E2PFVYsH0Q80tUl
TuMyGMWq00TmYxHcKUWrzKtHfPn2UlYUx8YaadQxcVv6SAGG6xnPUEV5Kx1o
1ILhpTMt2eWJbxji5np41sJ1hK0kDQQcso2fAdXgcAotxcUP1ftLspwLnL/Q
xftQVvY1HUpURoF4gxFiU6uRcd+AhyE6zHYvpEfrxZPKvOYgb9/GUQXxlh42
ELFBfhwjsazPvApAwa6Ji8VM4vBfmvuLZg0EKG0mgXK1vIQYa2KlXS3BWg0a
MJ6XbZM7lt2nuQgtimqQ67t9bot/LYeW/S766o+TQcoyyNDBAdKZb+K6V2Cm
wC4B+prFYif3MTAqvx141qx1LjE0sNWde4jyuB/rd+27WuFxN2g84FUB+eua
ayzfZq+N5k5LW8VyHxiICGe6uwndMuXWelNOeODIGUcM09BuTPrcaasWj/z+
YhJNwnJKOsXslPVpSVLPvpb2tL+EmB5Ou/WrZ+NA80uY5Xol5urWq6TDCr53
A8YmznduYWVReocAyHnrbNfxgpB7XE23Ubzzn64rt+zELt/bzmnGtg2sSEyh
I9KOGjrbt0ZyYoTynyVVzNShBoV8zqO2rXfzPxH/TXZrqZRllpyoAlQoMDQW
iqQe4kMZ3plghXSpgWQfxPV+zlHLSWyYRLrIfHoF3TMhdIrmwKGhNt5zvFOY
EaAllCJU5spHjZqpdoeSh1Zna9AakXLgy0T8IAiVFjzMrLLyBhZVTqEjujD5
dQrEEvF8zYZk5HR13Vf2N2nKk8OgXfpseJ1pu5Fiv7Eq99tgoDPmXtqAcx5b
1nLdUPPdsXqLU/Od42Vghf3jBy2ebW6l/1FM5mF+UUmjNyQkF1Elg++OuYYU
pSkBokao/PMVVxsNZMD337BIH0ge+LUmS12lM1py64tjhhtlY/X37HffYWC7
XlpZbZGrPIMjalypOxGsV4co0sj21OjMdAiIDXIxZSYpkpyxBf6bXL5QD6qm
TGAYMPcLy+Ocye3jRfkiv0Ho+9LKkcxt0vDCihYc4OlHBYjj+sthNWRIA1FX
CXe7NkwKCmZ+DJ5Q0e86k5v7H6OSlvyeNSoMHpJpdw4r45WZ2fREPRhij2BG
yh158YQOmCNNrU7YYi2/HEI8BuXk4HYZNw4qTi861hblVGO32SqXK1D3shWo
w4pghsSV+u7X349cmVssTYWP8Me+zzJOrJQddOfwG3kYwMgQQa4ex92GBfzg
u7R6jEfCyVK6gyCXlDGXg822cH2smm12lRRLtqSJRl3pSJppCEzytNNa0ZFT
29KMyhrDXcw23a1fgRdmB/FbtJnk5aTSOc5ISKv6HKMPgsoGAswYZjwl4aY/
MnHCMeXlkm1bBupCWeMXBaSBXUBulItHEZytKk8bvuPUF8fBhsDrHxMTimHs
UFrjQZij6HGE1ePKcIYbC8S0WhI5728g8JJE0aKGRtnkkQLu++oJUB+WgyGu
vdCESu5IxLpYqTUScpcd+NDv9nE/tRQCA9L3GnNGUbcyzRo0IPKD+fNuONMT
+S9sF/E6u8N0muMtFcrVFSDgf35JoYjH88fLFHJstS5+Y7JLwU5lA9Hx2ES6
hXx5ViBszUVOiY1DErKQyooA9YDdYN+lZCxFREsLAz6LuK6yGCWQm4I2pfxZ
7nmUHI3zkw29vpKLy4JdJQgt0YiCIzdgFI0NxHsUri3xpj8oN/iBJ8pYPMC4
x0tU3pLhoqtd4smiFvmN3yhI2nc4L9TFqKD9OJgk4ajlsaatU2SrX0f0sT+4
pfGxdkYcaTdwSOlSV0/7uOYS//NYHeze/09HpG9hHz3M7BXOaYPVNKXuOgG0
cRj+NZJSElUiOZ2fkCbJl6XdFVvgGgTEL6pBe2cW+rHJlvCMLZH7nEOR9FMp
mZJFzRUWLyZB2wJ/JCI5lQCL9eQGhIGXTTfKAZuZR/NWcoLqF17Hk5AK3qSz
KItaqITzm90OUWimPds5GlNSs4j6YVoUOfnTIURZoMDEfKP1fcXkp+xgh9GB
ZRKI7H/eWGm9YhlQPkNxbj6bUj+XpDR+OoBIr1CGLpelvOU4StOg3HENXAHk
fqpj+owxbsK/tUKXXbgQNUudKKlDsOzlBYQ5mgHez2gMbZf2ZdKA7ypWeIde
1VOMDsLuPgse47oEBsQDrtLnNCHQ2hpLLnf7FNLNyUza97SN82VuWOaytWNl
M9NWV3SPxixhC+RIYZWtQAQlqH4N/oPl2hYic7c7DFmxgKLI/1owExu5p+VB
JMQUzb/ZTgB/Y41F8zZiR/6mZw3sATK3NoF8YcMSV7hjTYVs/a8jT/zPnaJG
Io5ly485brC+Lyis7DTKt6LLvNt64Es+6Mlyao6lKx7lis3sPrP0waitdo7w
xlb3zwpIp7bAQZ3/gXunN8i2G7LHi1ofUqqWsvVjqFQvWjp4FkoqYZ97w6fg
QccKDo85D0AmueCCdfCNaf/VDd8RtFy++b+IgKOL4JGDiTKhmFp5GbrJgokE
61mZvraRYub+gFgE0zja6df7qiVQEkpiibKnlR6Xzr0NUQmLxoiL2H3fLedG
a46CBrhspp4qTcmCifd/YS3retyRev5CBmKebdfb+iECFXYJj7EOxrXndcRa
2i4EHhdTKGN5LSp64MNJEHliw/HVSON4U8g2Wiuamv6qLLTd2kfxGQjNfLtp
bK3utkHPMibZXDyJrvEWIWILnx05KfY2Bm0biHrOeJmkK+hN2u2uewftOmY2
twLM/fNDzFjBniyIlB3oJAL6HOEzMH6wwvRReB2NkGf4BvURPclqjfEHCpC6
yPWWHwS9xu0VzDcBaeaSbfZAyLaU2YJmb1I5vXuuFT9fnnuI0NdBe4c8e/+s
+tI55W4VFT5fJMcqZ0uYZ69Igkf0esTCDXzv0gUNAnIPeT1eok6TvnFSLHxe
qhv4KvCbC4CZRlX/Wk2p+xSZ07MvUIkffaaO4rxbAkaMbcV7yQHNsBmR/N1w
mvRo0YbbKmSVFOfHc2nI0OPopyMuoFPCjGlIrwZ0tXgct4V9RpkSnWbL5SjN
x/11u8eCpEdB/Q6VrKIV9BkbxKyYNwBKEWoY4ZtsFvVsMEbgSkvBm//DGref
9wEdoR1oAwW8NfAf222Yg2uGBjmRsElOTCasVJyXEnMGEL5o7sl2YtVk2DEu
kTN2ayY6Lmoo1GetvjLi0IgG4BJk61SvAHEddS+JTCpqSzFWyjHAUtNTJPxN
nLTxDYlsUejUpCovNoiY1+7M2LEJzoFysd7s5rZ4kxSj+2p7aY4DPf0q37Z/
Qfckof+SBuYdBZy7fFPEmB15VXRF95CbdXoxjx2S6sDp4JPjQOOWxcjc0R22
rRXUmfT4c9ivrTKKneEAnM1IIl0RZpuj9dTiN3vYa2XIknLSyVea3r4EqL4c
Ff++wYqlHdqeayYyc1mwaU6D4fv4HSdgwt6xMKr+mY84WtdPNimsAxiJOolN
DSSGFkZdKaSH0+Lp5AsSN6w6AvSVM+IdlyyHeuR9xLZvvm+c14x30AX9a/fC
2E4Rbz2gci/d+Dh7nBMuqq842J6mU7iIGQlYCu8Sr3M3rNQtmETk/HhsykuP
LkX76NwVfgDFm3y6ZJp80oel2xc4E2/mdcp/WByRcDJqvh//bEWx+c3yfMtW
lgC1vUjQQrIQLAxEkjsrpDM1GwbtNdYMu9mhTpgXKBnuSaI4Y/7YQYTkTbh0
etyIDdCKtmtfxozRhchb2xifN9ujrAZuPPkrRiMcrQ483kcAMwTeEo3lbmfm
PQJ0r4abFYoc/iCHOqHpN0g3K+S1VRvQVpgonClOqyeEjvdd9EoSa9HUjvYx
EsjT/S6Tu54lSy2LBRuJvIXOss7rqQeA3bDiXnJFp2WMe2uBD0pCbMYwtgkj
xQNs+zYL1Wo8EZlmXkf/xJn/HRICJ9vfK/mD5A/QYxqo7HH0rCtZWAVrsc7v
AKvi9DCv/l0oUuHsn2DVjfUsL0I2Qls56XAR56fD8cvnc60tc7dVUA6fyKAr
BakttQVP2i9ie6yuSRWhUt9H4ZrUbhx96wHlj6JzH1P4Fdc9K3RLHG8DsSlz
mjecavEEA5iCx3zeGCz1uaCPHy/Dlnj3bTliRdxHyVmoCdaugKdJe8wTqxCN
nchxocM6xTwhrAhwkr43t0I7NfpkL08jmUjqF7dRnolRzSKMvxezXUIZrhUR
glMVpkA5zqATmYre/fBeBjNTUWRjbnkGNjWTDcm/whaw+ovJ3wVrw4YRcknM
ZhnUO2PACp23Y54I3DHZGbZDmjWbPlB+6XHhJDpwMSnFjTrOC+AaVptm94hH
gnvo8TNhFZcA9JOsODVE4fWjTriXGIMdgQqj7K0wLzzImWrEd99KT2M8Gy9G
BJv8kmkSPlubBTn1wmBC++lvqAjB/xnmSXrBgSbFxgZc5pN92ARwUq+P12bS
XKcrwR8Djo4/ARv/5wV+xntu1Mu3rg8zLCeB2t4d4Qx4OKU/xX334TQJU8Sv
9lyb7TWzl52X7XLCTcyss+Q6Dq78ZyEPfNY5h8bQfU307w8pZs4M+2oL+dCD
0RvdIir4ASqeZ7PR5fL9UOikQ14Hqvmt6Y9n56+jfEOiLX/lBQM99ey7rJGQ
3zNzkacLYidLbAuy/9QfnTUKrBXpRqF7DpyAxYMWOJCLHE7EaOD3BjY8eCik
BmKfsmTLUnwBVE5XRGRRRs32MECuVoivBpYgKObJ3uH7tsRiGMsBEOQhSAtB
T+3Y5lXoygln/THw/HU0W0imHbym9M138l5JDHuUrLux1kBkENta/Fvs4pfS
v2poGVMHTGBtCvkmXmT1eISeHzXL4t769pJQuN7Q3Uz8nNmYIxfKG8zYCdZb
D2UbBCDFE5cD2NtNn++osNnneSn1MUhaV22SoetXpzKMxmUp3+4R0oJ2Z9cr
ObiePi1ARH5j07Vlzw3R9l4XhGFsBGV9dG9+07TDzPKTmtmTwCOFcrwyPcau
yaVwsc9rIJDdAxq5FvUf2Y5ZkI4orNLzHYtf3RJgoHKGu40RkrfALy+348xZ
0WYf1zctsdEHHGPk6hD79kbpj4NuIjwIPn4VyVppMl9eOHZ0gOShlAJfYpxm
Y/0JTTHcJMRb9O3LB5q2XNOmtf/IMwtzRSisOXlvfdyadwbfc2bsD6w1boWZ
4synjOFb9b19rq9x7jBg4eSriV2JY/kWYmcCgKWiSQShTEoMjJR3Q6FgNNRp
bz76y6tl3Rvbt1m4sbNO4lYIO+6lcLjdJfiIO3lbu1gYjxX3i8tk2/xNxpQ3
6cQbwXtl49UgjA/ZYahEo+RQ5kkwQ9D/RvH+XkWtFpdfX5oiJy5Tl46hlHSY
PEEbOXhP4zcPrSceYbmEtMuDFMl6fDtR9p3Fcs3ApnNQzVX5wVS6NVIuNn4T
xuV6xybqp/FEAay9ok5t9L4bKtJa2nvT8Kkofk5x/UutrRgM/2PZE8GBvgxn
K5dYMZbXlKvLNELtoXnt3uVcjlaQRLGGkU7tjtW7agMXb7X+34DqH3gGtUWM
+z0m5TQSkXGTZPvfRyeIUiKHVeWCBWcK9TdB7eumktTsfpzXuRQQDLArykgR
Eb2skrJd3t5Y2aDTElZEdiIUOoAjFg2oIHlNUysoPn+FrBrYjGFl4c/RvTJO
V1eNdoLVe36RA9wbjMvEpODhB0c3cG7XhMCTRHsIGl5pXwZJm3EkO3sYdfCk
iFanEAB2J1FIrH21KewYe8ZkvI8Kw1W0HG2HFG6i7KY33TwpYpMVUEdCcz32
DzDMVeHi5UMnYXWeKiQiLSDoXUsjhNxUKFCWG4RLr6v/b0W6T7SU9JiNSxcH
eVnaAtLNkiJG8Y14oyrNZXt1kEeC9V7Gv95k/jBMQGrdSeC7IT9pwKzAgaCb
VB6+4Auaq6M6Ef3rouBb4JcuOPPwANGowyfoZhdaixxj14YiIyx5Gnavvjd5
9FSdEDQFY2TL8PBqIWAgYsNpWBus3BBEI1kk0z2qKV5yzk0ZQmazcTRIgm6N
6dSN2Zm96qTcFUcXRqOdv/A6XvbIS54pYVfXxNfFfiIuVOcpdhZ78QYoixR5
0yMU9owd+3m2oVvgj7PZeBTPle2mTVvwcxK2iCa4OQ2+IzdwoPE+HC7b33OQ
9cGMEOKRaEbyUFnFeQ717Vgz1wSpMKtNvnsGNrFc3F8J+CrCnclX2Hu7D1Mx
E7azXQbxj0cGVkCbsEYGFqQZIC1Ld93P3VNLBpHT8sXJ373cJdJKHO994672
aLv1rl8olhj5Gm9DmL0B/SgJnd3vQyFlmLfjcPETeCzgEcfOq51m80FXEUKi
AvkJnM/a1BnDTE3DGkgNr8p6hn3IyCNTwEXxdAgWCAbToXuLmVsLFiR0Isux
7AVX725Ks8Jyc8SH78KVkpoA6ZqJpjGw/WYZAmSNco/vfN2CcWC+VHo2QOON
E162n/AGacqkWSJpqTskH3r/w34UC3Uh411ZFz8je76LF4i3Fpj86w5xb/OE
VP91g0Bilxv5/JQz/ugUk6xsS3XSYSUhIhyMingy5UkLFTHjZ05kL0B+mvZK
ewpJ2QObZhuqLSNhlfWEjhoR7B/MolsELI9L08+D5pfGF9kVjPW85IOUN9Iw
e9npjllO0jqoGLrFb/grHUJGW9txTf2ZpuXlQjcWfjLF0d4uRVoZ7c5VFBgx
rfVh9YxYf+o1taL27Ga/GvERBKD/xEfiVwFyz5i26ar/zCuBfvEIDYccJnYD
BR87ooTQAJI69918vwvKoipmTz/vUJsmEVa9QdPGD+mSSX+tVpVE8Sifozik
7CGvEjY7eWTbUXoU+pR6O58srZuUGckA+5/JDYiSdSt+MbYjljC67bKfNRNx
Dyxjde1UQkxyvl9erJhJjuM//30QIeoahmHA/CG9N8xl6HexOuVtze6M3Yai
mZPQuOsn5+jToaFIvnUDVimDiBdvYevzOae3o8hgxewdFzvSs14Veecm6HVX
YunrZqNM3fvwOKHT5F8XXvkAq/b7+VrZSRfjGW2+DIb31cf8NuYIGLfoSESY
AnJW5zgTxf5yzQmRs3h7Vi5fvzutKFI3gnd1KzhYYQoeuqrLEgO2220LVQpS
gks+aHVeXjIuRfiz9T1isv70Ock8CEItId4f2M1ynJpn2IoahoqM1wyysP2Y
azJkn1mrpEi0mB++W8rr9CpPSUz88PTDiGjD8Z19OgFsxSWxUEfHh/1Bbanp
B+eX7enEb6aih6NGaK91hx3RQsAVx9t2JgpE8bV7xIQC+NHZM4ZTYQJmGh6m
68kMnYF1TDSenLxhdhWArs32ZQ6eEKkRKLWsEiUqmu1puNwbvnxJ/kERiepV
jj2Jz6PfZ3Z2TUZr/Ka2LGzGucjn2NSG1Tut87+V39IiEA1dVgQ9QwIalDfF
9qjgUFJZI5AyG/94OpVFtP3aCbMd6kKv41yiu5wZp6OOI+Z2IOkYFTTJM5RM
6n+iMJbpdpWq1DO3Zs5bJHq/VgdmJr/nvoUL5T44zLFBxrGPiyACns4Dk8rQ
5Y8ejBX1jtViA/qBIOCD1lmIB0tOGJ+/hz94gTwke4j95ZJk2C7jpr3togmV
8N3CKkUq5uumcgDjf5s2cWaKimEOOjOvNjPBsUysI69O3aASrN/92RD88NMw
/waBrWRzN6IRTopGv7/866AaXwDVDatuszPR0y8gW2+NSmvOe8ZLLq5ogRXK
7YDxiGhciHsrZgIMUkm8HnWHlyj7zeh1etaWo9p+fug+ASJlBEdaNEfe0kej
2CaLpI4wt4Q4KMnnZ7HIjllUNvsc4SOsqvzr4Ouikhx+p14CzZjDtj9/9kUR
eFnIpMJiTzrcaWGitKMNjoASJa6v1BRw2rGzjSmTQSXSm8+dUvsCnbs5xl2Z
D+hBeiLGV4Jw1UksltCxUroilT3tg6MWMydM9bDH9nhJ82xRI54dKNKdDFb6
mjZ3/QH4z/OH/CVR7ndlqSyQK2UOYt8eqhMtVvsgonuQp3fB9CJ8dF+ZoTf/
mID1nzjaNmy4UrC9SudpUrSQrDngBXBxC4EUj+Zl+HOQuB1KRtIEdNkQ9J8t
ZupCHCehfq1DtX3i8a9keVMh1LKjuhrYK7SG2zvWat5f3JjOae4tY/Nr0YYt
inrnOYUINdvP2mS82DpE/YqjH3a+W5VSrR6la9rp/clbf4gDFKFkzs/b92Aa
ha649GPFGgoYj+1SQCfP9/6gvQSCAgrttHeapDOZJMonlIi/3olOMmFu+RRC
eyjyfojaIjSo1AoaKbkpw9JnOlrF4fQM0wKRK+IUmprA/HZxllcZDFWMoFX+
nwIQwbO4jSafLBsAnUmiCGOj/ZUgdhGZYJS4SzsPu2lDtmdmIdwtrYLMpN5h
9ea1iOrw27lPQ6lANA/m0J5zzA7sicLVS7gln/IOEQT9v8GiqS9Pue6LsYTs
pPm0nJR1Z/ICN7NZDpGUDL+O65WsQdjc9jox8ZTGIHT2H9jPXo8edkYfw8re
1EaXfbDQ03lsYiwJUE6HM+abW6fsr0cX1Eo7NV7qC3OZMC0m/dKbaxtANY27
xl3Gxifqqj9UYaqs3OBO0ThCH003IiixS1RPtB4KTqKFqJtXujUEz5irwP10
mP9tBWBlT0N9AMOpE0WLBPSCxbrQmcQ44tEo6UPpapPvsCWBUplK7ItIckiP
squVHR63pkXkUU05w16b28zWfsjO6gW6X+GEZM+licfIUIdIWcrEkjtvLVzb
/8jX1P5nGio7UflZ4w/pOSN9pnGhss8Pm/nnEQy1cq9OBIYkkz0IM2aA2YCX
AkVx0TLyx3XDDgA7cIEx5iy2mDUa89YT5QTWY1eQyXctsPf1ycPEI2kG//fD
Tr/YbMwfA0f7mflqFvxd3vIdz18XvKu1P3kftI0h83SO4BA0crfdiSKNhV7a
jBR+qH6w7vaoUSgYDjGe27xMRvCK4Jw6JZurbFarx6XV4wsUdos1S83Bgmj0
YQWls7l5+zEr4OEfmxNIb9uLLlb94lHI0k0QWkXMijzRdKHeYZTKtmtmosxS
c/ZHpznoX6B+5CuDDsRqjYtx6EKII/pB99AIvFqhTfDyUhMMCxOp4wqdqiZA
+oqnzwaoMY10TUI2DjLdIeNi9Qs+x18kPER2QR6YJCmBIFEsz/cazpbR5Klv
umY0O84xh+WtoxqTjYiAbTQ10rDGk+PSyKhcoW3xqZ4JlGvaLldtB+aHbvB2
n1cJJfBuQJ9LrdydgSZVhgz0Gt8Cq80Kr7WFOAlYkHoZMCE9syucM/QfEvdc
ZA18bjIdLFsFUOdWZ75ynpcoc9xUUYWvP38fMnExXWIrZpm5ftJ3z1JQKGMt
73vTSPGIR5nUBp7Irlpy9lZ+QRSq61/VI+vRyWGfgmDcgzyp/M+7XfwYGjJa
ej8G2kRjqoctHid7xpKGSJM9Yq9Ot19UNu+/AvRecZa6sP59mnMg5j2aEK12
jH2ov+EieGAl68WfT1bWXvEquQQ2Ll8xvze93EUBP7eDzV4dmqhCs69fPdvm
a1R4ZvOcCGX8heRA+Xd65DIhBBPUri1eYDDt9344joavU8gjzbozWXvfEwd8
mZsKt2EfRny7kfVN/h21loQrXiHUZudAQX94JtwCGTlsgemb+H48U39pe+Kw
yf6AFj4907pIS0xWrTk2CJOciNABLeZnYpOYgtKzGqeJ1zb85F1HDKzAT2av
9Sa2p/yHU4s7UOcO5KjY3BS/7c9V7RkMiGr27yzXB+BD0hH6wbZ6T2xpyOrq
+hUIshfnusQk+d8bowvCJkfn1WxYcY5BO8KSjpp1KEoj5LdJ1BODuSuXWLoN
kE47hgKCSX8Uv9U24K8/MgY8N3VDrVksIhJacIyYNpXLDSroGHQDOjgbBBpA
2VAFRRIktv+em3Xf5Ju6ev817o02mGMklYQDDZrtz64AIoTX9wTWH3HMNW0T
V4x59o6zkIXdCEccTV+WHcLiEU6XcnO3nON3CmEelTShvq3zLuCs5nn0i9w1
KWJRT9ctwXHGoBShWh90nDf9hSgfzmkM/g6rk/VQ3nQOGv1fVvM6BNTo30oR
I7lJ1400ObtMY0gFpCtujqRHzXYIEoQlXplsqCmZIvK94XtpG1amD5vmvAF5
dPn/y6IHhnWsRCFzKNzM7KVLaep/rIKoZE5QSQGCGq2D7FiIxWIZ+JUvJ5fM
4HPt1SkZdNevjCxRjS91s+skYWN+s1Ctq35Toh5YtzmPcIzaeT9fZbfZJZSv
WYv2GvYWDOW4GisG1uMFHsn5RoBCmIK/no/WjxFORxzccgPrYpfovE2VtztA
uedxTcI3kRwadImmfze4cshUzgcXNX1NJnMxABXuS7teUnb3AeibqxUaASHy
17gas17ldFLe9fPyCOqu0X8xRSeUGo6v8YsJBUuer9P/R9bnEug8a11RL5Qu
BvXrLlNQQ5IZaPVCIrlqe2Q/S0d6OnaSp7cNgwWUZ9RPpi5GkpFexor9iBLF
q5EJrdRgQJz8lyyfl7TvQA7AQ83VsFlv2/E4Quu/9ud5NVPX63Li5GWN2uv3
LaeVZU3l4JZU+pwBfGmfZ4TGhRkcMVheb4+EZbZ9+XKzPXm9DcuK78N/FvKT
hEsMA28DbXhk/KSOlSzOhX3zizE3bstWaXOoiKKnRMJqEscp1Cwd+mtQCQ0E
lqoUs6RLlFRfJUeSHGQqg47L+PWZz3QYOKKtNx6R3FcVZlY5n5z0CziNZZuc
niIezxjp5mf409cl7XiBYVtRrGprPvEuEQfOkCCDqiWAtTGGUHo2lLsT6wUf
sTi0zRCQpZsvy9LaKMzZ6fJsJIqOQvTI3n2wJjPY30PHYKWBWAZSeslGzodS
gwBAtdkTjVyQUz7g79as4sDQmooI2FNmCiv7lsfmXnwCFBoLi/K9hPILTVkB
CP/+9Jz1w16PKhA7Gc/fRxmmOSzWWmmm09TYe1mTCnJMoBGnFJClT6DENKk4
y4AnsCv9HveTV8hsCT7S7NgNonDIiGgfgf1TT5Lk0Aoxdeb5HGfHBR6vuMB1
FcXPS+ubCA9JXA49ximrAKBxowKvdEIg4Xqcf2cO1lrUcBKrLxR7IO39VZF4
UVvPj2/2evmhXF+otbGEGOhr2o+JBh0BL9akjzJBwsZE9VY6z4p3hBPblPs8
LUJrGwjT0NPRCaslE31zWriET3iiGehlUHI/aFeJ9kCoMrPJJ5Tql483gBti
kzDdhEqHdHa9oJpxcgJkIkKzenBK+SjHEKlQcSsZJDSma2qKIK+Ssrd5IlDe
Y4i8gsY9GcIuGqRNrX63E3vgRBp0x7gFq3NTA7O7cMQT4QxH5otiXhvFDUyu
5Zfw0vF1Bh/59a0k3fg17/mz5Y+1W/yxzRFRMfdpZp6GcfLSLRECdQUnWpqM
/Ao0PPEnBl4JQeBxwMdNWzu7VTb0LX7wEosA1dSQxMLNLI33v33K0NgpWwhJ
HB7Z8/iuBpjGuHAy37MjhBNAXHUnx0ugbyNhPGUFS+//fpMgcc1uA0Xy6JE1
3RYWy6S5G9ze6aGLiLuPh0DkTWrMvGyl9OG18Y9XmLc+fqX4jhuc7PbM8TGK
jWAm9lIpLqBBl0mLi+xLIGwX+NMPbk4YcuX+Fd2goNeDeRdoACP4GbbcKHct
vU57TORGL9uRa9xF3YNB3gC/4pQX9qgTO5tEi90peUBiWlstxgMjbbfeYYVi
IXO2a0RgTvdpSda6enFBh15KF3EHy/A6WnHJQDp1YRYKP3rndy4wUcNFk07K
g4JkcMJux2QiP6jZmgJZyDIVlEbT+7hYlpBfgooHyGbEOUyxKrbw/6OaWped
I9e00t6joHEBw/4r8RxXmcqRLcZVhKWiTADDxCDnu0BzQGTfX17gO9Qn8W/c
bmPf6cks1EV4e+hIAetUggHgNMORKJHqIfNgJMSS8NFjbMTVzClY8WNQSIQD
FAWpgk8XxtlMEun+/8+TeEKqIDLuNUFp2QNlHvBSkfuMMg0/90gF8yEJqgNb
5VHgylRs32S6EcTMSRwS6xFrHPgaRpT6I8g+j+bLqKAv0Qn9+2lETvhceQhx
r9czobLKRQmo/D427ICsUZskNs8Wwwu9Iyfk6Em26AaM+Swo6v2jLAbIUmbZ
9T4QOkb2FRTJSRTnx1YUBo+BJk3uHRhBq2pz7cOyDCDhb6J/HBV1WprNuHkh
NFTdsW4QsJGOj0lPYCe9N7NTYL+rwhvPQULZmeznIetAIVoDroO+0O+ZXHVx
8l+AOfzz7jOxhD2J/t3JcxzRjDK2PZthsWjC3MF+0HjSBATA2rmcURDPvshc
eU224yseRwdtPoo6JQWrbN79K8m+7+Df9FRGF9NFiYQmtP7lF3OcHb+UC8Ks
WgKENO6hEpMf0mZR9VMcPIYyWobS/N9Rs/Om02aibTI7vmk4qM/dQOc+W9se
UmKptCgPhdvAdK+MlIY/6fAq8SFe6qbCH9mlhBfZlc6330B4poqXQItHPqhu
llaWWCmUvsKPsVUc+Q7n7GfLjLGco3kg3dvSXttAEpLtTOmMt7Uc0ClZt8Ud
0Ndb6hU86xeKj01VIbc3TG0flkGZBTPbj36hYT49z+SVCyBl6frr20hvcb/w
k2k0OGzQskwM6XkvkR3OjwjcTscTZk/DaqhdWHdfSTknmEgUE3KCq41RaSup
dQTOfVdNaiL+kUH4U4Q1zzlsxpctjKwpdbxzCjKcT1LBRR5wj5TDi56CahF7
RPdKrGNjOz5X3Mo8Y5k/D9OFyiifma96AvHGgpUjHxL24myPbD6VYrzdEPSK
YI/8sVo4w+EXF2g3APk0WKiyGAFZOzCBSHaMrGu7dlQ8y081vzyhQKIUdiIw
ZAPvEZ1yHEdJgo71pjQAewX3WOsr+z4034PQbbLvVmPaeXKUHQURMRQqPgAJ
XeSCXAZo7ErSjpymoQR6VwnFex2g0853iEYEfqsweU88/P1Ug5VjI0m0dy3C
2hmXXGvygVRVLntaaRhcim7keHkXdBiN9w6ktfApFQ4L51fRSDh2hkCVhv72
0px9lhLGVREQ5y1oLpseSXXQ143IYdc4RHi0dkMd5MRbcT0fV5HrBcvCH+IP
Zydv7YrrD47Bh+DDv+McMr5hgNN2+0xleIEzQCwEi5iOAIs0laUROwsYopW7
5eaMvttVBoeNNKVd5A90/VVywKNN8AOL2jRe7An3IcVrClHfZ264vqslVk+V
OZ5xf3d9MbAjYEvkjtqwr2YD99aQhO9WeEzlaUGkAggqEjDWISiSNajup1yO
sGdnKzumXcBPAFYGUljZ5nh+cVqx6NL/ulLVpguEHwJGFnOzIf5sXU6DPmQ9
3rO2FYtN7TGNfbW0P5SCvWqd2lQ7o9suhzwIDTiSsRU3cVCj8+y/zXxGxdcx
nDHFoNFyj+Zq6TwegzvWX28bEsL6B9XxCxaV4QNnBP0T9Qgvpgs5uioss+YL
lLvvcGo/O4PhrSTxRB64Ff18cBoTyPZKp8pp740Da2u6KAUePjBQyHXUhhYe
rxMLAIDWZ/SUv80yRRakg2hxYVepiFg7ZqsTocGD6985Oyn97LlmK6zcwQ4O
+CEpTwt3DFc2UzP6NGkNx3WXO0uzdWHfuy/domYtVLu078E89VIYK/abPuKE
YrSljeGNYh3pjc8Ih1tY0tlwr2uhtQuqThmuneX5azEudH0e5aKM5VzDjYER
5og+Grl9XYa6aizSG8SeSQLTQWGwSpFudKhNNPeY3ccB653xm+RXeQ48is9p
LvUwvPoxsC2ncEnsv4ume+ORGnHdFHNE9+8ULClEnzUH/rP8zjKoJOPMV/kk
2tOJ0Bcr4CbA6vmTvWamnzsW1r7rDvf3VJl8Ig28j6r4wF5Z9sI0bTmpio7f
U8fGCO5m18yG//87/snF+gcfMBTN5HbcwY7xVFzsGsj999yYpXMB+8b7bfdN
yi69Dss5HDkJh2wi+5dpSWVh8SUTaG+FCMEGYqhTjFfT2nwhFUA0S53rPLdx
T9nNPL8ltScqZh4FHQjWZV9R33Nc2efsGZevClHZmngPGz41q4dj9sUrgvLW
bVGoz8CehHGjPosQ3fcBVXXPkbd4Pijuvcru4ZPEV3usCNcGEHC1R23+5/Gb
0S2xJsHtERTmnoSaw2O2a37dmQjFBhRg6f4qHAGE6AcjZUTV2/BQOcSjDuhP
aSIPg60VMUd0pp2DC7BPLjsyp9wO7dGiYPdwra/OKjLjNZaAwJiyX/nNZft5
HTi5nUqTb2JNd4ooZhpQQapqimE2lNIht/dupAZmhMLr4yOtE7RMw32ipbOi
35AXBbVLHGB3WmbjSWiW+DNnDQzfQkG4i9/P92RFVloJnNfF6+KI9q5/rWnY
2dUf0FYfMfmiNIjjWTiAHVQ6e5Bt8AeP6Q8mFCr7FFe3sx1jjVNpPEhmFmTb
uTtfAXpJHgIwpxEVMO0PXD52sxCx2JOelMoBlE/CTcCsInvadXJTOpIHVYba
UFdUO4hiibyPBxaTKs5mS6oMPiHSCDuvU1+KxzRoHJobyCWb39P6yG6SyR3J
wrZG7C46PYndq2idK+3c5UWs8RC245acWwAP/n2yd+YQjLSec5jMjGynuz7B
hxFQsQxioy24KnmbcawH8WnZ1Sc2kwCYlBwbaE35Am3E5nNjWh6ziPqMHNDA
FNUejkZacJjSuqZDE+HBWDGAop2CVoTFBvjtbEwvEpuookm+1Zjz8jcgQT8o
WGgp2jeO3aF50689HTXSelcQ71scc9OBeup5BYvdnC68cnB69CP9TARJ/ElQ
96B7vNK8eqY237Em5B4an5uMqlF84CbgGSkoYzkr2nLpdWwVrbF0jkFgSA8K
y/H+CosPERBFW4ZSbFWrYhaql32esNtY9IFTf+0SJmMfj/eHLMcH+7A/CY/R
iTilncdaBL2eUyInZI50Ag4dpJWrtNfE9nfRnwSnqSgayyOGoSxYSGual4G+
YYW3sByg7Zw1Fy5AO2xlFgzTM8BnZEYPuGAVCYn4gLlyb7+aZl4MsIx0Ih00
d9uBB1gPhVs2we2hb3QJ1bRiNsq9d/ekFi0FCwL4gVFiBLjhoaLZNnjmKBeI
eJ24J+tO3TirluXZ1+HEV72t7kwl34a2Fzk0eyB/+EZa2P097XBDmzXVn3Bb
VNyGdp1STZ2vh44qDsTgfdyU2lr3MOop8C0rhjeNaDNrUdVliX85CdaYIp2m
ZKXlpzk4DziuKnJgDUiz4IGWejCQMWiHr+MdTscAsTyFyA0dwhSP5kq3n7z4
5eZxy6MfbCBC6EwqUf0lc03Vv3XhtdiM91BPCR2UAa2/nz41oGnWAoq7Rt+N
Zs3CSqrABYOBpRI31npWfu/Ylvp7saSmlnf7Tq9oLSDOzehpnFr8z1LNrc06
faZr95Lvj9iFfp1dHhVIGH2MRBURKS3fdddDTdjWY2hjNLwq8Mvz93Imiah1
owmym3EPMOWxfQ9CwEyKGwRESdUEgmDd25xbeRWT19kcglLHY4cTnGNh0KVR
VY+3E/twnQadW/yzj03CClzL6W+JLflubGXsLGVyPBT7TmaAQZnPupfq7jCP
hrdQLcuBcsKG0xp6RXMjdoaC2xIKfD75vEbgqQvD3W1wM2ZoaPowkNLxaol6
LpTmiLxlqizSapRyyu4G+qH4IWXUGjiygPNDK2OF+oTsfXzUOo3s8GOFXZ0g
5Y7h0ZcTUj03gINkkbzVbyzx7y/amS1RnxXhx2ftjjI56it0j6erzxD+7U+w
ZioH93tLH3Ec2nLEfCvN0XMqbNxFT6zX2QlhiE/HqopjvOqQTxTRDC+tVslX
2xW8IwnkuB2Fr+PW28iMglnmhcmnWRHWSKzX4r06LBqMpZoXwDvkBfuxHsf5
te+pXr2tWouc4uPuA46kw7LQwhm622nf/S3hBHc3bDqgTH/2Gm+kwtie/P3n
hY/IxOt1+YQHfAjJT6ZcYM2dUTllmCB6KwsrBNQ7CrZqL/ydqTxiC9iXGSaE
sno42qKQNI7KE/LpEpcMvlOzpJxBgqO/12A3WctnR3EBF4iSNxGcmGNIcaPY
mMzEkztOxUNo5Gdt1yyuuIXNrkolulyF8uvFGrsDZNr2xnaEe3NXbr1trEJO
BN3AEYsolD1SAmUGXV70LZDI5935nwa5aHQL8QsQ2dqcV/ccVeuCK1vxuHU4
CN3fgHbZ+uN1aDzLYbN1PuwZNee7SELveRHuRtXRrLUtfEVZWS7SpmrToQuU
CWRFhe6lPQSxVMz25x5vyJ0mZGVvsExvUg/NhKYe5/JPkkGr11ero5osZLvA
7YCoTThkNuUzq6m77SIzTSDOSpLIWa/yeTtDxXTyEu+iAfkvgLIV4lHNSEkS
hMHNnIvFA4qmobJIl/nQTV3SxT2/NdH7qYmcoiyMCT6Er/IR0Ylk+g468FZc
UWjLQALYhGAcyu2Qtmt/PxzBsy19bRoKtfT5O4oKDUpKB+JgJcuj3dOx81PA
akDCUkX07eQgYPz7sEPcQ6HkaNUV0cJEt3kEpA+1YT9FRxDv7Q37PGW0tvzU
Cn/0MM/xkklqMPX0nVg5J9uZnjr3HAuLE+jUGbySVtW7YbEuf7jyOqZPWvj/
u2fRzjKiRxYbC6XbR8qE9Hgf/aHabiCKZknSEmigIu6bfQJsVy8mgx6vPfcv
jlqLE1XXwhJ9teJoSYZTHCTqL5W2zMXySJSIHR1Lz4L+UXpkfxV3MiKSwlo6
QINYYWsUBJPMjVexNZ3occAseqcjGOomAt6WAXcXk7W6H3pAbmFAgHJ+fo4r
KqE/sQ4EslL50awvq6/oj/VLQFlwwEwFFzU1nnaTqYsPItLzppCDHoWblKxn
b4gklEgZla7OltFntS7BkQGTb2F03Ofd66C5v8+PH47pQuUrUb1YdBj+pG/p
5h432ULOF6EgNyUvPhZFfUVjd7HGAQeoH6Kjah314QHN0YMA0ajxt2nyKuj8
kIxJZxkAG91NDU1Jnj9RtcwwoowVRxwvprMPillMHsXqAaAnLhHI+9cUG6Zd
au4cx/GauXusSZX94xVT/ijjNNR6+i7VSjQBCuqCO00N6NIuReNVxkNxzFtf
AdVRlhEraIs5hPDXYca5Oe8BykFruB/zem3dlLZQ99F/YvuuWbHMqeQaO5qO
S+vmf90YzjMo79MJAPwC7vKpQg1Q/xxmUmpbpEpor8ot5NK0YvvDlXqKUwKz
0VMepJeHhfwms4fm7dqTnTyiyCoyp8ZXxLDrp5RPdAgc5Sr1RX0n0Ty8tcA+
GOicgjRjCsvX9xIaeyy+WBV/hfMflXgUFprruMDxBPdg0t7LI0TLr1DxiyhI
MGoFk6NBDgS7z4iD5C56G9dXpKAmhJed06EQLkgH3lN3EoqVBxPULpx68IvW
b5nMKfzCxn3s3p4poDtFeAP2euYRNeLBAsTi/ukiaONWmjYcQ6RWjz9yxnCf
B+yKu0ghFm8mzew5ML70C8Q1REEnV2GJTrzrgHG7W/c9lZ6hxC5TVdWi6meU
etxf0fHoge8xy2mbzj5UpB41OjKUlBEyoCkOfWRmZS0O7ihZEibiFSTzDsA6
g5Z/D8k69zJuke2I0CFmJaiHVu1jHWD8prRe891LfVfzildlHxGvqjmIGCGc
NmncZQ8M7PjHbnZ3eMbt8ZIFDr0n58lG4O7WmAxaiaeKuJkRc/BdZVy5yAQn
oLCka56SrpRjx9k+Le0+NqQytbrtT18jDxThxPpmNKBRj5jpargTJDoVyJKK
4Gq0S6tZKRCkfJdT743IDPRWeAJZS6jIT2bXwC7P7K/KHNURsmipqOUcO8W7
bBYYJg89xS2tTTaeS3Yg1C8N0MDaWtugpzZkwtsFCy8Vw0rfB2+20xHOd9Xq
TElyd5ESbaQBREr0lGpL53IN6fluic/rkgQHC2+mYE29+rrQVOaUsmJzRgpK
Wk6xHr+LCYuIv5qfrK9sy0SGt4RZF8Vb11IbvAiJTAdtNQ6k+fxuobgJKqSB
bQ1ZBFbpejo0RuTc9YKazKSVu+QJ/zPcc+7iwNBUbh8XGwIZKb2F9JS9ndGF
CTcNqspnMtkFZw4LuGYxuuCvBzy8Z1vgcUmNYPMIjCZfYblkjzrQfwv5M9p4
juZ1E/o36CfUnBgguuPaDSZEvoX2li6OGGpfTPd5I/4DZ5qg1C/BFuVa8qyU
+MGPuFOksRKvpeQrktMWhO0bsuCZiDCaeHMINhzS404HIt8eZF06ly/K+qZn
bvTiKQY6wCV3MYKjFgmP1FpzZZOznlNpS3P/zZlFSBxyGwT6z54aHR/DfOgX
E4nhOlPOrK53jZ1vbPi0H45+wIPB085q/MMWaCJZRj+ka6r/P+ArSQnBvO5m
dlRFEnzfIywDtAyJdMfAQi2lS1KzOUSel9TMvecCX41Qv+NkmBBCJIzu+StS
n6OC0oKTad5u/cXX+uZz5eD9kNbjTwVTiaI6wuROcx7tDiKxfPpFXwlEeKxR
XNfhr+pPGEnFP/nv+nVdZefnZWj33S4RFmg/pLb+eFBf7DKsJ+HfxrRdvrMD
Je9TPUChuqVjzxT6KZabKWL4StFYZJDP+4vD8gnlpT+C71xgFyXgBOHiaa8a
7qJxtESRznHY3dnh05TM6Kiw0NGhMKo8B2g0AIutC+tXmh4a3bNu3Z+0bNGD
66tRsilxWjNC4M/jUapaBFuljsZrAAW0uEtPRJxDAUg58EprTRf9+kPz/wAo
aU5cwckf0GEQodI/NrI62zYXzBXBVcY3NVTZx92ZOQrZWFUosHyMYEQ5yoAG
pDz7IiiYkpQIDObgGELu+z/Bdxt9NHsfNSZMlYYeZ551aU87pbPzCsKJpAZn
7E479StXNjDGLRr+ufRprTe3K50+v1tpwj17ZX9YIL6Sh0d0fzeZQDrar5zR
DzRksr7dDiK9LMSWyzZFDP6WTJd0R3O1Wr1hyLsLZZSZYpwu4+RpWWxIvUOK
wl8qpZK2qZEYgW1dvaOXNAiZqNUzfO42rAPx645E4MM3blKOytR7Eh00Ih0U
D61zsJYYg4j7e6v3yDEJXnPHLYSo7DG3AEBz4J3si5MiZ8ur8Sq2qHmVMhYo
9bvIpH17GqQ0BshB1qZvP5PbMzUORZ3O61DLoEa9YMvdm8PIcbT9szoAdnYJ
tTnLzFRTr+PzTQVEXAZgc/LXY22CUtGvIs3Ey1NJiZqq71ZMqqNzcWoCdLH9
l+NKgFX9Q7ekmP1MLpPTgP1BndwoGRoGJEm2jkP2Ngi5imgEQA7B4BEp2IR8
uZAmhu7owdnvn10MLb8VbZ3bd/dzHJ0ZtSrSUu/UCPw//kyXFdwc+S2abYDe
YhAFOdLpjh2pOJmnrUOm/OfA+Y7s+yvG/HhJqJAbbnfvxWr8vXUkFPmWoZO9
C7DjoPjm1f76+JrOmwI4Ke8RWg+WJ+sfF1REhHQUtI0mg8bD3d8CEMX5PXtS
xCUL02sJW+UHPcFv+SXa9MlIoFq3L5pkG0MYBnrjk/Z+bsMNm9/RK2EcbCRa
er9cQ5zbBVmIpPQ2eezwY7q8M7xFuDNqkvYm4CvaO7HrqNE1xgXJyP/rcZq6
Yx9Ru729XD3ded7BWELklOF7ceI5iuep+7nF5NEGXchvyXs4ngeCpBBj57oO
1wx23LCfr52XViPSOu0A73c2Y0FP7H7wNnE9Ja7ZgmKbJ7Sj28AIBY8cSGUh
+A0U9/UPun08vOhE5wzwjkDJr+30oCS1ZMxCqN1c8IN/UOMGe0G4/6hhFKo2
RkGBvOegWVLxiXUJDERDQnOgacLQ/kEL96GB4NMoA48WeT3fSB9Q5ejPJ4BW
btMbjv5eVwPxErKi+QdZX2WbnexPLgDDfxKwJQNiBr6kIay360W4Bjd0nZNc
ucaHSexF+xIlkCKx9e4I6Nekqw6H9eY/gif0FzYBhlgaEbO2UBKEjnt7DcSi
RZbFrhFf0XaXkDdTb4rV4rQDXQqiSX3BBI/NhxCEURw+sjGoLvC35E5aNfXZ
5T3XCY0upVTWj4bCfuA1WyryrOKhSxjDh69hHCSVxKvqKq/wAHXhPWQLi+yo
ti40S8ZnMRne9ulCxfZCy5av27mnLVynnlZ3n6gcUKyRu7fFYSEKdS3Z938u
57riyqVg8VQvEWZgn7DgBelThi8yYlqm4dJzi9njPIZN2ryZwvjNs4QdgX8C
0q9EbPJLlDreyRFDSiMYXBQl21RSXx+bUasmemf8wPhCv0I9/4jcI4shfvjX
UOff7FUkUjm8gajsxVuu+CKu+PCKV4aKPlnQgICPa4f72fjVPYG7G3kPiq/A
THpbpVUx4o2rGv71Vk3p+1PCuzjrw1ssemsBApuQ/qrLorO29qDom6mLMdDu
s2lU/u91CQb2Z9xEXZ7HcvpBtM7XDhw3a3rvnSQ817G7WZ+qNGejm+IDohID
SM29a/8m0MNggJa3v0NnZMCIvDF6OX/CX/snMh4GdMg9/d3Y8L3fSkrJKP3g
OJRCOy3XhK3T4s2fWRly7SXwYkMSydI60uwjisoNuWlPjOg3IsE2eGnEHzt9
JYm/m2iFG3EtbHLSpkmB09h1ecRamEfGGGSysjb72VySvSVIO6xsTNe4Qr0Q
mL7PRn3fBGiMXlsT0kOXrrVihoPOJqgBYFTPS7WIxbngzetgEnSlRk+ax0cT
9Riv51MGqH2yp8gwAQhFlW76xgCwIbSqS0EZoL0JPvy3+Ri/scBPqDW0xQo5
KpFCU/8ncZPwyNEECGzgKpXcarfYXcJJn5qCN9M8wXUlZcY5rInbTMzF4OIz
fAOdsG9yDDLzfNQqPordlZ3pe3fMMQrN+QjvhU2QHkTIZQA4O6ZyMchjtg3e
BEyVSY8iU1m0PoMJIbmg45IwnxQzimFUxzQ0bZFC++93CsAB1lqAQzZN/J4O
72SvF9NZgEVZ+hNne4wIPkPhAG+IFLSYlXxXDCKqXUSBM52G3Y8ORqm96yn8
+k4DK1b5BUtRNo8opcEqo4N4Geo/ml3cLTO3t1KPv6aIv7Uko3YqFqBBJxei
qpdB+43jatQr+tAb4bIxwx89CSwGSWZ30qzSNgv8Nvcs7gccoeaZNnUklmkW
jhsXv6evNjESAZ7zwa4ptIxotCk+Qb8QyUxaYSXZ/ah/GAAvTu+DehkGywxQ
xP5ZvM4IjBRrAsmfkptuodkiulEr6KP8pvkkGsjxz1X+MImJWtP9sjzoXwyY
hh+QvPPBE3YHjDPxJ+1HUcgWiy3ycIQN3wAWehUsPEETFeE+vf9RfeGWx8Hp
NmfQeAb4+qp1EQj+daoERJZp0SWyeG9gzvqv0lg4KKk8JeTQg0W5sSPNqT09
MZoFqpi7bOqHc/7zUwzbCWNTP01AM0qjKA7xplEUN2kjE7gAYvfP+Cvij4lX
Lmu7bUUatH9kIHmy5C4c4nq1xnis4O1YpCdSIWXZtvtq9CS2bJB2VAzFQElD
xy6QpKtwbg3FAjYlMvM+DlviSPEMoETkXlm7BeH0X52lL4yJ8zTygk1dYFj2
aUYZTyeNwdp+XBtuxwMaCKaAXdsirfZjk5mHZxfXO9mIM8z+WXZX862JEdPR
vMHEa020wQWkiO6lMrc+9jHcHa7RciRtC7vlkB4RMgP8daXz8zv4ov7SURRi
Nzk+Em55QXncmU4VjMhIaZT9jBeEKnQwraEL7uWXHSxDTpA0IPa2qB6+7pwS
pj2zzJ4eHh0tSBpU7RGrCwnFP/xLwHgLWR4TznJx1q2aXONHI3H9YndFEsSF
Iy/RJzArhnDYS/WjJ+wi21DiktIWN67CvEpAhdqFQFVTElUl8h50mosx+1Gq
ZgiLT32paoV6QIS7hnyXfffeAcZul1LIgXlMeNmBzmTIPS9Oo74zAq0KnoXF
SXhWvioEyuwjaJPrWSzDcqGg1smmk8euX2hDs37Nzdj6VVi1Z8mhzcCKUGtJ
BmF2z4r6eVCJjAxdY7hOEu9IzL0RcvaixZGfI5yU9QJaS7uFXlmllPcO2iCY
t5KgkGbrIVIC75201CBdSLsIQ2VmPRNPfna8+WbGx0S5LYj9cggpvpY0MhVQ
3y3ZK10LEYVIMhAvczSMkceAkKEALz5dY7OUB7xIU3TX/A6Bktz68m4BKjK4
j7QEjiZFBCFyO6YiYPCbBviKLmgHUfPD/y1+FO6yot4pP93DsUSj4WsLUYBL
gxrpZNFjnE5v4CdhGW9NMJX7mrAtyIRxwu/IAqWJBKY3qDztc6ZzajYLG4ao
e+D7zOJybL+6xRyHtMWNQGgZPYqvpGARp96IpHZlbp+tcJltzzxii6Fdm/e0
zhseUWAU+q3siZNoGB1dRs/VHhN9nLTR6uB+fJy39T0YyqCIJ4WkU8KZ5pp8
oFg0UtfDPkSlIroKGeXeevkiGDnH0ff5m7hyMQS2QdY4aqSrzrKtJJNtCYqC
UEc9InuDmAGukRtBdKeLjehohMN1BBJKlnW7nms6XgkuJLihp1d8Ih2c2hS2
uNqP3rJRh+6frTYfPw2I61pngjK5G1gB2ssPqjl/jikRcENYQR6lLr7pZ5ep
CJX8hmcLONH1LPHjP4O3hJr2P62lW1d0lIQ4n57ZX0MOjpfDG9FrjEmIzoed
8tI4mPfkFYbdB09MpsO6PtMJtYZ3puAFrOiid2QjT9MaP+7RfO5AJRYuIdv1
ZX8d+hgdfeMMdTC7Y3P5sUDL6XqTo9qFtI38bY1NcgGKw/8+Q/CF/nSxZJWd
2TBmVXGXMPQz02vXqbRL62d5FkB9NwecxfZ5cjBIO7a0jRV/+ny4BlVTt/ZB
9DDnczsT8GoVpFO+vU6lFFSjrIeTEMLGLGWq4xysrG78p5HZTgnzppQFlxNh
H8X2Rf5ghnligQ+AQ6vDQa9KCH8YwWKkqv2E1lmXsyVN4H5CQXiGfnTDovZh
pguN5F+0m7jKON7Q+QDMSUG/94eKiEzXoQGK+fT8EppGi9zDAC/ObYcMlQ7j
/QMD47VvigXYBg4UVaiOzd1qgvRvosco4Y+CyTVnNBRPWcvgMIV3Vj8zLT6U
KM863DMnTFrqlMYyt06nayezVUpuvykx2dAF6kt78Ysy7/lVJVw4l487QMSh
MrHG5oP4K+tGR7SwIJQum+Ybdxj/ZfyVsuQBfjwy28hYzJOId4sscOrqDCH7
4bODHTYYfvdjONCnDfSZ4UelY3OTzGHOy2cZEk3jCe+XaHKPgYd7fdl3FvOU
TjUl51RqhqghFM0kjsPaRapnFrLy+1r/RLutkyxZChQSGxLtiyCKba9FWPh0
CHiG5VYw1xN19oEimDnq2fcnGDWxKcJraCKa8DUgyDY2blPfCO/VgrDVxTwL
tNHj7u3GeMw0GlFBq4rL1bOdF+CYRMUNjmKu35+9QMhecz52hmCsV//QLB4W
z8vwwzOts+CQPRevCrZNFCcFFAAffcTln088I821OZ+jCfoHTd5RrlxwTlth
a/yXqmvTTzVnSmHLZm2Ud2a23sMxQkRrbAkXSFW4xJ9r4GDuFAvcsGHcmqk2
LuhvHx1e5e92xRC0DQciFxZYcN2qUIEE2HYw0XP13QePOg2M5e4FSSlsG3fD
TBB+MTyGrdWOCPXV9OQH9ocDihgUKix8XaOWdqjB4+y8e2GYhHl8qVgqFmeT
MAE+C9+j9KwV/ZuJQ5jGC7zkeDg52N2BZc06UFCERsM1pjqFg45yZM0kp6Cy
MZBm8H/xajPXj+TkS9Rm9Xg+8LjeHZ8NATmjaf3xRccuKxXcELgBSVpoN9Gs
cQSpGcx8sh0h5Nbz8aDN6zmWlzMCXE4nj6DQLEctw3TI0m0qPQvVkUmM6oMC
50zX95D688P5+JhqN5DoK6yo5nMp4oFDo9nupwELz/Zy8UHgiVE2CY21dFxs
LMVvKXfJlQycD7X0nbf2eGSATh/uS7LjYrVdadhF3GJcd2kM2GJMQhqyagT+
DD0IT6rukPAajeYFAcmGKislGtqB4GVe9PqKbJeHjXUqhIuK0vYK+kNf4yaL
QvAJcvFnhjJk7LXJDyTl8KbNhHouEgjyN2w0+1LyHUSjwTt4Qdc7vyCwoaqB
IYDSm78/Jz82IL8q3wgnSKk5NvBbb5Q8yXUs97p8JC90kjV4qv/ZSEpCTdoo
63WWqsxuATPSK+fPphiL+UUyqLoBc1XWawxV7HHcIJ6P90WlTp6NwBFMj9hX
ayUAqzEwBiP09076Y3b0i7rteM1d9wvKHNhsXiTwF+SSN/uoS6/ZQBj/Bg53
jo6OOjNV1VlIBMkG7XwTRC15N9THDvNmyZlGMTyvAPO90hwzD1IbZpIDDMqD
UsCi/Ur2dCgGMufAUigFlOoVFIg2rD27KL2nQ9XOFifG1tjpERn9ifVRamrB
erOgif+uh9HbRBL0RkYUSvy9qnci9e2CCYd8FEV8d2Q8XThoXSjS+dZKmc7G
XGHSWBP6Tacs0LERsKLK643pxj7QZWeIzcv6qWyUe5WqJq8tDoGOditPefZX
VPBZDiUW4gnrzPtWvdKnABSkDLAMrU61QrevYOvDPLUIWr2+Y8EPGUKVGsnR
pyiEi9AhD2L4/rkazXHwpHKsbuxY1jDi32SKTLVPZU2WNMIH1njRSH2xRm1C
BuPvVYIpU13WDfnnPRKeOckTkuR8svUeeyxSfKruZrpI0Au12ob/2ziXf+Ij
AN/luyel3lmot59yTw+el0Frkteg0/k9FGFTDJ/UQwHqF71b5L29uZHFd9Xr
XJUCupF8EDger3Xd+54lEF16faQ6KroEJPHo2NX/fkoelpzBJLabXcPRxruY
3CuRwY/hmEUzhNT9mPhX9TXCgtYnHj9HoR44FOg62HscbgadJ8s+8NcIM0BD
o7X1Jyo81sltstRamZiGazM0VNjO0OaADaR1BSDz42mISgy/gLOwGEwo//wk
+ocskeR+ikTpO9GJ4oCJmmjBhIw6XnEoGUP31bZC6qG59vYlKvDHZx0ws5Vs
1sxwpRBF3sLHmdCSA3kwHCBFQ2Xle37veh/ki0rDFk8C8kilYejhNNhdMp9t
Cdr2Z5WTfvM9gLg18qcMWdG44Y5/3lAfGm9OpwQH7WXFVxLF5/SDf1/5YyOB
b3JT2CLUY2lcn2MFBge8I+73o+pn3nKR7qbMLE022Q9jGhhnjqKQ9zWyaiEk
Fwv9WfiwXlhvM317MidFF7D/VQhuBTEGdXxwXOU/VAhxEJ6ItjfHTSXlN0D1
3EhrTQqgGQEVOnzS4jZQmmMKKvRTw9M1t+j/zbcDWzft8SAdYX0euEww9Mqu
N4hNceGr2LV+I1exrhnUBJFX5fm7HAJLvQN6ekYxg9oQdArf5I5fm4T6jDsD
b1e7VRWWHMCWyvibvgecYaXA78gbj5IdfQczAaCSkJ9WfbCpfpbhCxpQH2Kn
XHAaugPqOvXYUeIs0RySROyib4Nj17gp+SLEUahVvKcyWaAyrZLqcLM7myT2
jIMsvSZRCWPo7r+pR1LSkWBPk4tLoG1/G8TTA/6S3T7OwvI6qbt+4hQF+RFx
Zz3yrq97sbxOskFXBs+7w/TpoThUXJHEfN3b5KwvUTeXUVmHKb+a+tgKej2A
OwBq9DtfFVDne5Yc2ksO68E5H3mv5q52qIsB6GnyRYmjd5oZTb+4kbyy69d4
gzcgftm2lJ/+AtyxO/RGeb7ntZ4HqSuTNvg4a/kLzzGRYYLuU/EVr8g7AWxL
c1h78N97xxrfXj1uxQ2Lhm2Ov/cA6axmgmC19qelsihXtowM6oMGpYeItZ6y
2QQ7YfcXj1HzI991LgGhv6ofxDqG11tG+zi/jnQDHlVd9ovMOcx0sFzLjYvJ
cC+Apa2AobR6iJbESVo6D5a/QfF4V+RjSEahHmV6dpdFr/TviNR4OGzQjXcC
yNL0CPvflhrzmveqf/ov2wh0v6rdsqTzGepYzfJslB2wRN6niqgOCptqe3Ar
x0lrfwDU+K6YT2dHJk8BLlvB+UZqYSFkSbaAwL+UT0DYO2+9mty5/fuLL4d9
Z3NPqHRGZJVUqjI0c6VyEWdJqREIAWivl4/Ked4OWrhCaiy/6uobdOwqzMvN
AU7m1lSx5DFFBg/y3l6vfxa38499AO4bXbA9N+sqWej94QrDTVWB2HaO5qi4
MVge/zNUxWJs9lXhsCFcI9urjEiLWVq/EX1hyhGWPK1mv2nncZIEYtGgd1o1
XdlFiqL70K+4RK1WX+xx28znzJSNboYoUQDxXlVJI7XOuP+KGg4hhnX8HJZe
rXOJiXthB6jbfA0r0nHNVTISiGjfQHQ0r+hwsVT7OTUQBxwsF9t/DB5erclB
8xbgC+zfedtIugj850mExQAivT8YsqlSLGUG6gEDbDH15Tuepn8X+y3a7cvi
x5vdMZwou1cilnCHOEAeOOEqBB6PxEKE9J4Kj2Q46Z+MD+YHc9ZmMFBqWTME
V5hd7tFkdmUMQHunbLV81hAIXcs7hQ4BXgWX98eI+zZDQTcgGKv4sJySt2lg
IpFmZSuPm2ZgsVsIfNX0auIvMTyS0CqHlV4NfUYXO1htjYq9qWlDPqA/tDKz
DF/r/HSgOIEiDj6iSrtVpi1gbu0NgAMHN983ZqKqZ5PBVarMqBFENOF2eMeE
/jDGs4brJA3QHECHG79FKXfpUUIXx9DGY5Z2M5R6uUaBMWl883J1ZxFWTTEB
ZY0ovs4SYfrM9AR6b1AmKUUCHZExzMekc2TONUvRY54zk8GvLbvuhJGcFRjB
svsXtO1iaxSYgIJZ90qUZ/03rFpGIc7lNp4W8V3+bGVacIQVnqfCXnp0JiqR
g13yC+AhQOH3BFl3bZitURcdyE1WLoOuH0AASXzWTL8YXh/a5AL+guyoGo/I
jYXUInZxV8acQJKoZOy1FC4mFF/5S9bjI9y0nze1LLGaF3CPPc1ZyuRtHjuu
ZckRKtK89SpuMDyFwYXZrxc9LPOqbunNDGDx5ZeOcKh3p+40xlaxoSq2fJIQ
YA+tNKO494Ww25TI1EprATOPlR94dsnbRqtoy3Cbd0V1L4yGWF7TnCVThaJR
NSHPs3GLz2ogxuD2Wd9d8Pv/g5qRefA42u4IqHs0jANDkKRTchvCyfo/pCC2
jnw1eZZ91Fe3FdylAO9LW08zZcnE4TTXhizgVCrIPfWR4j+exCNr5JfAwLBQ
FBIULBcAf+eiOefhXGs2RQHSDOUULkqD9bIf58nRRAXfKyND4atXXgeHo5Sx
UmBOfvMpS9jO4wTM5A66dQj9rm5ex1IRplQXYAGZU13eEYR4YIwjFITWaC6T
tIM2MXDu9ZjsGFffuZAvGYoISkMlt0d4xjqmMAzHDJ5N12h8Jiu4H067FnCX
6VXYsr9KEKFJQjhqIfCgkVhgGFE7LVfp1q9wC8MI+lDFERVflN0QvCw95mcK
aHteJapzpS31AfNkFCX3mDYDgQ3XJQAWbrF8yGEuPfCFlK3IY0elLQ5AD5iq
TYzxBGzaPEki+3PfNeTsnT0NlaOpvhPNvfOX+lHZ+yf45DjUxnd+gY/3+6ya
dhh1CICnEeL7qygutM1HVfqiutKHg9Kw61G1SVwbPdZ3EZiFV0+bj+leF+IJ
gp0PlMjOJIvxDpMlOCkAt11x/ovEVxfsZbOWmoFKrfv98ffKN8gjnOwArBQI
BD9kZBSoOa6DhShz9e5B6yEHfcBiEDw+5pSDExJVXDNa8tRXq1J1VfqwqL7v
D4XJ+7VyDQCd08Mxdsj6LLok3byynnBMtAZOQef5TlbbP2/4rgNG//fixaEq
+o0jurRQSHVJ6cVtOrKBZPqNT/NXTT4b144cZR3zW8UTSD4yJtZdPBn8bHBL
AMS4Spcm+mMIdsPqOtEkP75jMSZYdafWQnw9DkcLYyTvF4DGXi6FeuwWfSsP
m5TYY/IykFZDxcD4sFsy1eZGNQ5NuFcbtMjPFJtdgVDRGWb18MdXjVG6oALe
szNg4zHXo4XvMcqSrGNK4SJ5jnRinjYxzrb6fee1hTlxqkU9Uh2fDUg8LFA4
dFgcHgBZPssCr2MyaqYmnUDhzmwSeX6q70/2Wi7cjRH2MjDWxJmbiGczSKtb
dPBI6B+BefbqceBGo7YNpK5H95MgRTftAnmRKFcxUB9u6LHLiFnsho45WyMh
mvbrvqR07kjBkE3AwHvEdwjSkN2nGu1K1GCGiR50Q8EOLJqZBUtvKRPpiQXv
fBv19jizC/ZdY58ZyrT6VrRx5rnLnKc+ePv6t3hYlxA4TtBz4SnfsigGk1lr
W5Bewg/t4L8y6d5CAo0Js9JxcjnnYV2EfwD84hkrfokQur+mTJuVzFM2W+bT
YMb3HXWENGyOtw/BScZIdNP4pvSl/oK8YZT1fdAfOOxIVy4OZf+hlV0cFSHE
rCo6pxGOcsYk/xs/AwmCZkE2ZXoNSnhlQqD/eRbJ+iw0iOsqXu7Q/U2SDCFp
jVMMCModbqVlGgHO1yvyxvptJn4ssuN1WN5tx9u3IRIn1Tq76YtowUXyGFJW
IwQI7astnlHOVDdIrJAxFx1fStxpnjY+Au+M35n8mIRJrp3oGRdIkWflgjn+
Cfl+OgDMdQ3caknaja2ZlsJ/n8SG7HhL7NfU0/1L92iipkMgYmn0+dnFsu6n
g5LHS5+tN1jag0A33850uzcBZUdqpw2LXeCU6GZS+drc7erXSvwQFBhQU+Qk
4VEGR5iq9ws24fJ0m8YCypBXSmvLFgyjjeTaRirIbcJVvUGyFgnGpqtzFHJM
7yXBcZWrG7qtvRTM837sbxJEFxyIozYYjRHIfj8jt2bgUcqBIbgF0dVyHWKb
dyCCwme5zoNREgr2ApHbyJj4SPLfov/dbDgEnICMhTkOjWNcPz2pXXdM9n5o
70atWy3jB5B263O2ylvn/7gIesfWad4kPQ7JWQfPa//1gQFXX3u+QDfBT9LB
VMVDGY21H+l8bBK9D9joGymB80meA8avoXAJduZcv6dJJQkXIK0xHncXqxsZ
v6ehKrmcFtw0Corzbhx0gwCiz8uCOysYQCk5nLhj2IRDwjenWfArjhrq/cam
izl9/htxZktOm/nCfEE78/zSo0NJfijf+cRJOXyzgGyS3Dyd1RQwcOkt1YHs
18njijN3hOtRe7JKPOzdMFbwNyQks7xXeStJ9+Ec8jmJCmq2MSQgN0cwNxKs
ny+fG9hXVFrFMNRahGeKLP1T6KSsyT/o32xt8jvXWAqfbbCP2ScPc89SVQXU
yihlIAMHjXNG3JixBuepjhDZUQTB23Cav2J/PHmOt+iEVzmSwyArl0OgExzS
IfXQWZ4oDbAe85qcYXRuVWaAw2etYb0HTpd5j2Zymg0TkaS5CKlIsBhFV1D7
9XLYkSXu+6WTf5cS6vZC26x+f7K+icf9GkMwasJhrKUTzwAEjKAHZIB7mPz9
h9LvBqLSpARLgu8ZR3WpeCodjrZ9WbW3k1y0p82961yrywVRf13B6QPSOWYc
7yUY9ExDEcHKnH97Nh5/opkRrOF1z+OPYpLms2X4uMJNpMESAc++F3zLWOmD
OlXEKFaYlwpVtV85jLTjct8jF+xCZsw7VTl9yA2n0lC1P/z0wgzMgwUY+Dpx
MtAg9EpiGmSg6WXuD8PZiE+qj8U7+mO8o7+pRkqPPOps3akz/NkloGmi9eCX
IE8v3p1S6xbuY4ehC9RjzrU/Y7q5zLZ4VoidOzTEhEDd3MpqekCmGkCCx3UD
nim2ckOkja4OMHOOflS4kTLXnm6xp4pj4ZDpd8y58G/V5FcYqrUl4bYqmqri
T04rLvSVtxsgzJqXWxX4Y0p5rif+v9XxxG8vJxeYo2PnoREBLcDGVSNiD7kb
7j1ATZdoT1sWcPnwk4yp6Sxw+tjdbCBGhQshIzcOjNjSOyhuR1hbJVsrm/vI
y4VwS1k1xP7tQnOHugZj/rdRBKeZ37//BwQp1vJAQLIJq6uAuMSvYXWSFez7
RruOMu8K73SkHGX+pl1+HfEVH1gUjjs5trJN2AIU2rRNMtNuMEjD1zAUpyAU
2ir78lTfULCFD0xxEC+awuk8vnV5g9HQ/DVOp8HrfCb2XDQseqeAguL98Hj9
UQEINJb80kzWPCq25kWN43y8sW+K8tiD2V5Ewv76hInJQJMaMj04OVPeos/G
19k3H/+L7WPElCBSLLy0rV+zoBrHhs9aKG8Jc0G/a06kJ8fqM2Nu+cgSlQfG
Z8ezNYgt3kbuqa0E+nG75eI4FTMUC2UzpICQWhtGVnyTrZiLs1g1dVIo1I7B
TnA/JefZGfL7UOLMTUNygahqgD1OLbsOlB50HA+2C86qziE/dO4ugfwvFHoR
cQ1C2fg7yODE6/knn+g6+DDgZZPyqRGQzERmmGEwsY7tQU2d1O4IOWk6gufw
2/CIJA3iH7MHMffvs06mC33Xb1xh5pZsd0IiKXly53AXD7bREttCzBX2b7Ch
I/cZAAGUrq84OOOzU6OC9jszCskesnhwdOyryOkWNfphimxJq4gQ17GSNwmv
9YdCeh6Iku9eYMrRqBho2O6/PiQUZAuImQVodkIeoTGzV6pkSsIAClKNDFI2
aSoPXNo0YYcWzuETrSfw7RxWTTg5Da7dRylMc/BE1M4//n+8MhV/OU83CtnM
AwyrwifEojz/TqwG2jvAxDRyIuwyhmJsaUv4cGmW0otzW0/FsdLh3QrqF6Ea
Wck6X3r6Ix8w21toPIu7V8JWMvpFpy7MWLDJdwSXgiTT1ofMsMatZ4P5zqMx
bDoSuISRML9UoI49Fkm1BIlKbdlNaFohathCtJZGjSELwjO4n+ph3UaFLmga
d/RbjBMV7pvwJ2KLMun4MGmPnL3MbmXH0lFxS+w0mriuJs0O0yLTmBTw/lJR
1TYQV4umZ6qVzVL1B/D6AhcqjGUtNqEK3WHerADOX+F/MVv0qn/CcizUrVTt
3qf+Kq9eLuth2dnwJYLfGCenIXjv8BP6ILYBlw3h5Lk1N9n2HXXoQOwB8lgo
e46UBRA5osuiDbpN3H7YA8jSU9JcayE9u/mO7Yf7EeCMJqGJKc/ACupRvX6W
3B39nVxXvuzV4zyRk77AwGWn511s9fKPCXn2TWtmZTgImjN88A3A7wR0hmGg
53so1kkwdADeeVMfJwTOqcW1zcUNGsfJzzPJMtrl4VmvtYnndy/lfVY9twlr
QGjJmP99c5uUzCeiZrVGQVznl36sBjPEgAnsNWpjSLmWrYnushtJ7+90J1E8
1Xm4x+OtdkJq3QawMrX5FAnKAuVrRysEeJYNyZxvGmeJ4jGRPHUOz8r3jL5M
HEcj6++kKmlmfS4UDI3VRAfiL6dIHA+prS0riIJpP9maGtFu46SGtqSRUdOG
tuu66n4SgPTLvjOMlzyS9wdk0OGAbGKG8UTBv81k2l7Rcf17zQfpkmyPA4Ca
ijVR0n40XwFayBAznjbNV3Q5YqHYNYhxtwuvzv2xV0x44J89Y5ZXa8rRloYB
MxEVutkNqsiL3mIwnAwP3pr977NzpOjCAvb9nplpPDU26TePhKHlYEdow6nq
H9jFJo6xNOV1FrvXrP/x7LVtwYuQk3Bg4kUCmdY09CZkkslpZj546Qf88Z8L
yoQQnDD2ZOPgb1D028myuO+ed2QCO9o/0JH9Unkd+8A052X6Szks6qRr2u2M
16WIugY8Fg9R6Tr5++t/uhsSaifsd65pQFEK+po51of/CikW9L6aHQ2XJgNz
cfcpvsGnCcn0OcbR2Es0o70BYc/pIrJgsc4f9CfdEc6XNkNruh8gBUdmoU/C
23FWsb3kG0y3rDEaUxDMu7Cu6kxXAROhtS40Hi5FeyJgRiyRHFH0w0WOl4ch
vMgFlOL7N0OTljQWHbCWSUUQpnwANvsReQJb61spAsGqVoxlB+HKQ0FF6Uct
7+1LMTtUsfuGdkQ3lbrQFHMu+4djMEHFSu8jVZ5L6p2VYEHm3gseZujf0aP7
D+lEnkbx15+ZVNJ+7VRI9B+LF100JFh/xz93hMegZ1y1YWLcPXsiSdsLn6jA
OiNXAp2HG7b9w/xnubokBX/05Z7n2AR3ZncL1QPfTsqq61B1MsLcIkusgtLY
tQb8IwEQgtSuDfj0Yhe06O/xstP1bl5Ti8tqOK99v3YSK9ltqmCQQYxtDK8g
OUTsmq7QLNDiPar8Ax70G0I7MkCYBLxHAof/XDQqNUidlNONInC3F1+xRb4V
gWObd1tcmmROKjNJtKW3mlng97nw8GgWuJZeqRrPQ4COFWK1NTBh5s7npQA/
eaBGK/GE+O9ek6DKuY6PEFRGTkrBBA7VzmfRk1nI+5KHsmZVNPK5xS4ucT7a
YJlW2ONE6u95VlKUWRbIIRClRt5RKkiwMCUlngmkh0Is/0xk9QhrdHwCqErI
NnGByPzIJqeTGfZy71H8Zino+XAgOyrcnXur8CMNKuks+RQvbuwARkIR++dR
P/UmfFlT/H48iWjPLFEoG4b+9RQO7FEj4gG5V5cikmPvTiEJcUlMupdSAaej
d366/senf0/wW7Jfy1SWpCvrduJgio1hmGqI1HEpJU9av80592SW7HuiGyAr
Nck/5I0K5fZWXwKvVc8vcXvnoaslTP78wvXThg8rrZgeg4ilIbKYPmeY2TOV
nXXFauXfXAbbXETQYvTwWAkYm62vpnvhSQ1OKTigmNsswu83Tt84CvUBfNK5
6aLZdANo3btKopbt6+FbTmETXusfGCK3ldaM61JzmFFytzHKewIqR3rAmf5l
3Ot29XW3SlLdS9xNUjeRr8V+gmBJFTm9wTPKaX4bxcL0tG5yj2ZqKPlwnIcQ
T/y4kLmCHApBoTF7EjOwIJx6ZB+hBSYisKMXgm3oo+BgVLPiaHbUyd0eZnq1
hx/UuPx7q587E9Z2Zpqocij8Y9Ug+jKuoQ6FIrCDRItcrTKHcyYUBEY7wnc2
cuT8aMzonRZwTXKYkjyRWIn7bAIF1eIRkCUiNWU2M4fcP0GXWboO1qLOQXPY
W5Io9QFMxdc5L85z6LfqGMcyauUg/P2k52JbNsP+9g1Osq3lPG3OrgBEAYMc
ZwIXTP8Vp5DYBnPx/Sria91bx0BJG6OxHYYknV2Wq9/R/ACNPBGMZj1F+40+
JAepmM3yoh5k3F8mFJ7QZ3i8zluwA1EaMF51atj3aLdjhNCgJTPj+gsGXzkV
kkZ2WPP62mCALCBTQqdK498em3fcy8VPPRgUSbb41xb/FPYobhszvhNLjXRC
Zh3NapQV1LnNMLcB2tpQtqzu23boQfbEgA4jqTpQzKKIEpEx4ef6s60uv0if
QUjBBZGWED3DsUJAcqlH8XyrN34LjfCNHYVCKaGNQM252YjHr7Bnnty+P2vx
9GFB8xXwi3A60Bwju50SPl1KmFzo6syO6VmKzOWKaciBlHsO9MqedetIng2+
R2y0+CqHatb42dcherqdJL76F/h3XRW3KNb8P8ip/2c11XKGleiiB14x42/q
Our2HH41Kcd1pNjZtYmakIk+WrRPCsrzp7JUFnFKIMjVsTJ20uTjGeruyhof
U/Jiz9Klhvur5JGxKaDkaCSEc12TGth/Uw20+trwmACabjOq4AuGlTxLlG7H
58fw/qMdz42NQqLkl7E6kNNh80hM+TH9+va0pWhv61dbjmw06hCMDK+4MfRz
sCMFBtcl3AdSzLCne4E6im9fnEQgt4SUkxORk08plOh8V+kUeW8ygxdV6B8b
FO53qMxP0P6Y2UScavPduL1QKxWBdJX0RvE/8cbDAK3lurdjhWFXYF08nRoU
OHj7G+glHHgUQ4JNs1lSQP9/1n6++E2iR8JVmC/NZg4d9VSYBAqGvXWX/jnp
7LRy+FZir87UmYRBHklchfOGW+vqCmFB4ILyY31Ma5A3X2vT7F/5HtMa3es5
mQSAcENj1TPbsHX5lRf7f5SrLm4yKvB/LOi1scWEtL1d3QTADW5dUNTDCBZC
IMfj4RILDeTH4LWNNjpvrRYjEGUkpFHbfFZp4Da58Q6RAwBXvaFK2hy6PqPn
tXCrK8oRzlRobcuXe4m8XAfpLOBWLHYpKY0VzA/9RlfoNhm7ZjKgDJ4kArxZ
EBbVLiyY3we/gG1nyhhgwP/sXZ2pKfE0Zzg5RmHotHz7RMU+ZktMoPuHWy/m
XvTLaVptqlEIP9rwDuSR/GJdmqLyjwhoY+q8xtR+E14udaajDLPrqqAxoJiL
b77lOx9lvJTp490vDpt1E0yChfx40B99RFHaJbfZ1uqscHf09kdlOMpHM4Q+
vVfWbUTYBIViICrltos70VskHx5hKngAtZZRqM7XjnU7/56u9i7TpX8emHvm
8jH64pkZECdDPT0fLc265AY0opwjxnERmMgtYzVJF72gIueFucYTCFvVuanP
iz4fIhUmwwpJ08MJHwa/F154WxTscVxdkkFQ+AwPAFm+8T/lMTHWo8KxVViS
ZymyVC2HEOA4/GxBnL5gWaV7+eiOlkDtuCisK9adsRzIFDJiiHuk1+UEjBmK
0sr/srydaIQ7eF82azGE9WxvDdRZighomgq8mC3IBn99HJuL6X2BdfuAPWYE
Ic7Iyrm/GAb5O7+Iyw5F++cJDVEygVQjbB/st/aDoemtT3c9l58JtkY8+C/J
vLswkP2s4hCWRgMf1qF6IceeEOrcTuIDQYUA+0pf7vjDkfVDT3czPTXbJsHo
T9pQFE9V4pavQvCrrPbhwQd33XHv4JdJ0Th7sktpVGa/TRQLSEScat5TGUXM
BuaokbWcjifEkIqsTdXynCyto2wIisv3p5KJtBVUckMgqwI4CSqchHoJvYmr
687Ki74py2iyFW2gIK1ZrfBDEjUFclsnAhI3CD/zha8LGXGrRpXKWkzOAH+R
8InWsyj03XA7+4F19AQ1Lk/wy84NkxW4kgMP26RGd4nYGLC3JbGHzFiv1Pa7
/sCMcD8i/cEhoo9yuM62ZoJqz7F/kLyD0FuCSn4L5Nq16NKPGeiANJsm2hM8
j7y/SWR5qh91ZOWDiRoqiC1goPlOSc6jMPwSDcZPaBghrtJWQ02hmKIte9mp
QL7HTP9sGz2KwQoSF/Ws38jOMlM11x/SCDCQ5M9ttoCixOg3T98n72l8GZVR
K5c7LiSzaNlw7u6DOvoS7YUf/wqDQXZ7z5vYaurtFZK+LnFq8AyvQteDRChz
hA5BbWYufFtAg8GvMGn/sz+qYWNNVELxK+sLEFwENDPRm2QF3NOZtzY2jGS2
mxUxNRLJiKUjw8pkUxXd2hFVU2vObK7RM9rpz/H4aXU1xy7BH0KjLeAJ+yc7
Zze1AkhYWlvTCvf/oRqTEcdx+wgtUXvNcnzABWs2skFKjVVfdl4WJD7M05pO
xnkpVsHHEDNGDoQ6484dp+3CbeeUp6fGH43DAhOgEPJngHCfqmrMqxzyK7Nl
WqjtgLCsLORokqY+Vm8JNCzC4zsY4ZgNJXib2WZhZqM/LmJvtF+Hlt+cXieM
tm8s5VyOp57RmhbIvcWqRZP8g8V53MbQ8c1tXPVG49hwT83/yaipyFMuYpk7
u9DAWfuPu7I0epi08ACao88x5hmhsJiP5vyxBTQI6UFuk8IrPcSYwiQ0j3yd
1IBDX4XD+x0JCqXyomF+QxGIQzMsuiEroVevFmaPOErdbxO5S4lRIUs9LMHO
6RSO50WTfOYAJv4RPIRlJBX8svH2h7iS+Lj4O2UfEvYeZR/aShytdyPcQoNn
2e63owvUnaedzd8JdrFVSMctyeAoahrnDtIVSEs//QeFA2MmSxLM8Z+UXm84
r+8FiuAqUeCChrel4rztMbNeQ9O+bi063jlCUIaOWQjlK9qWTDvVdcGr0vLo
DgdLVfNoa7EBM1JpWNBPteUY4rkERvOomyjpqUvT9LsHoQ73NT5o4l9EANhN
ggVEo8GtKrfAGu5dflZh6ax5w09EFWRLLURRNtoERi+v8khqd4yO9bMd8wrt
rvS6WsQsXzjHdXTbneGViBEOcb+jgJv1UVePzpS2MRiQrzZoBk80EUQPv5aL
cpdEpej2qw6N0Xpv5r3G+oKnPjl5bA2ICc5BazB2fQ+82MOAGip5+9nqPQZ1
vVbJ1Tgw4qI167Rqr4oHbYKO0gHz+5omC0U2bxQ6aBx7QSLH3lAqCToJgW7V
FUxlejXMQW6G48ekQtZuKwiZhf/Cr2bjKz1lXyS+hoBgIS2epih18TihZDlM
EpiZL3Rt52JLenYQvs9674ICzFZwwvbR2oP+6VfNjKF3qFgVdZ2/0GU4OZX1
h42AbTBDxoiPXjZNs9d8Ecq5tBCEu/RWNQNM6my1RCWi+bN3RnTc3z7W4v80
ATWEFhGtJwPMidBltvp1GxcPq5jiVjEeed7AjmUM8y99/GkDkRO2Vv50SOyq
M13Ora1feqK3aQKlHkYWJZC9z1Uo3DJE4mNswY8FSrtzYI/qQFEFoLc1JxrH
n87iPmhn/GcSdAsQOf9l3yuEsXOh+D2MidNDlna5whVsIEL6qJCxQdq8/ziw
XwqIGFtfJAAQrN9j7AGWNeSnYiS+/AB0+UrWqJxKrYtVV14iosj+NSHw7ld8
A6dXv00+5GA2NGqpmrTvmo554rs5OyL2vbHy8LFr5Q+Rg7oTNtWrw1rTL5yC
pJkPwNQuDo46GsCiSKIEvO9EGnlcYSIboMqujyJA3B77LgULPjSJrIHNeaYs
Rd27REczaLjunA0xlnIh1a3pzzRC5Lz7d377eNkTWLEkn8PdKGP8F9VIfqME
o7zgY2TJJ+qKIDjhQGsvbQzwTlI7E1iaFoLr43vRrWYiSJK1ZFPwJy6BHa3K
t3W9QjM6nGc8oJnbqy3NB556NachnTC9E5860FQDVmJ0vlwvLaoBLp4B8SL8
3ZpaxKrwohSAnQ9N5Eu2vq5E3iMw8wmeCOhNsZKrW55/fizETlmzNPqVx7ec
sa6FzKj2b0yEZrBmh/6dlkKr0Eer56jdGrlshjbjgwPvN1I5lHCyv9TyKBfk
a/sPrZ26FE1y7AK6Gs5AG+z7CRcjTMQtkuLUnqHbb5/o9lEk54JYgDzBhAzX
J2uwbWy4XC38g0CeCkhRX3eP/9RdE9rLp3YjQ7med5oj1ISkAJdmygEV2PuC
lA/nGHgih/9gItwcx01Q/yI5cwGsAF1fHw5r7XX3hxZLeoDJKjHmRq+zKLYr
UdEOwVvhXxwSxfw5nmZGk2vlwx/taUN3JdnZ2dw1pp956zMUTwStBQ1UAhIA
7/ditnqWbI9byBxqy5DLFW0ZbIJ1f1/z3dHc6kD1CEPdWdxOII0q17Z57+3G
Wf6sWTwj+GkiNvoukLoJcuade07Xt4QH094JhmRG+t3dZa6pN/Nx6mvRKW/7
CaZVau7ztbthRfDSnSbfXmg3pwaLPEfDLQn+tvhQOuEQNdCAnRtlAbQ/Vm9V
tro1Td8+e3JATrwz1BLEGw+23KV1hdn8i7M4hNyUqBDEmo1Wt82x5g/YBcsA
rc+rpdK8W2ZnFcnEiF9+LuMaOH2ZVnq7d2mImqHt0RvcrDp2FyMAKFn4ILH8
fi/ISMR6tV/imyQdsX1uZ7MGjkMiHgQY9BHYiguJ8XER4u2sQdb+BN98tUxY
FO8dGpASGRAFnBWcHvcuDOl+S7CO7kH2gLiNfqlhHgfBmpIpUipkf4GMI+7C
UKLPpYPgHWMnih9NWgXnKBtU8TBrxIvAmH+Tzo71AE+FZ7eVX9Y1WMsvoClF
MbSRI6ziXKx3V180J75JSq8afdloqtboBytQfjQDQeHaFukBYc/xVSdr2oYE
+rHG1VlpbbhSLwINGSDoTH9d98IYT+lLs95Otu9jLdvZrOhA0aKvCpxeft9u
ytqihFOhtbY/fkTpIZIglg3XhNjrvQ+4WgtjDdREAmnoyqQACcjUoZgJ7ZsI
pODFjt2YBSUd/KwAEZQj50vW71bG5fp4Jk1tCjqOVkCU60UaFyd964ewxOhB
6efasqNn7mKS5IR7A5WBGC6NxDBCStlp5eVwmN/kN0DAfoABUDXqDxMBYk76
/YwuPPB6Cr3L4EIniA8Y4f/9aCbKf9h8hSeZxfuU27SR5nMPuiPlEfEeNzqk
U3iyBkxGVu0PNr4pDpd65jl4qTnV5RPwitufSG9IwMKzvlE6YQHOzyjz5jMA
NSe96UJ+ZftaaZEiYukyAK9ybZAa+kFT6hbibfm2Fx5P6xARGe83hTwvIc4d
5Qwm7PSK5SkblfNqfiWFvKYSLBQyNsceeWGLcoLMI/tBMBcfua6Voblb+ITx
+qrwavkVP8xAo29/BxHFuElcfowZ8r4dRZ7znkvQ2vNdhf1GYIWKUQTY8e2D
WkSBjagVk03/MwPtmULPuJiDVgqgtQwE5C9YvBnppOVYWB5RMl46B5eMsUwx
EIc5fjSVubfs5j7G1qOUPGP1pegoPt65JfmLsEHKW+0ODR+662wbIJBY8Sv9
dWniu3JsCkztCpkDF3jg1/VfJRk0RUiTzqErptE95jGhsWXZRBZa8SnLZPFS
v5XIK6bWwMMs+HYbTzetRaEKW9I7362zWtgsit7/XD2UPrGcHpOygNFGp7X+
O1VsJj5SvDgOuX+ge+NfVhEwo63b6z7/dNwtk8w7HI9417l0VnN+9cLKNE9z
SuO6oe0DTAelH+Gs7GWTAmVzY+P/vsK9iuYVN+uZnPzJd8T2OUsZk0VS2W0K
c+Q5lXf7cBQINyWO07+Shy8wj9USFnsZ/owPlC64tjXtqdJTEKapgCphdKW7
RZ8uNnaOV/gBovuwhdGWV0huEuIzFsQCWY/vJ6iKFz6jaAXFYOplHJ6bihcV
kne8IqWrh5sUWuMd7DWHbFkJIanA1jU7lylbo23cThSzvDB3lIH8UE+JZg/H
JIxsYbu4KYuN/TnDMOEh/NKgvBoVRs+gJO76dam+wC8d7FF890F6Js5lRQPN
29gOZUpFc2hqH+SnwgrJH3jRgyI86+qYRp4mEpduXfLvFzKu/ESzLMmkxfTM
za/gkbTeWddJ+meIUDtEVSOUiFpj5RCl58Y4KNh6KooZyF1IhjwnIbXbqNhB
aEfqoJ6KZAOQwLj2pcNaDhiH8yX71Iou8vIR8lSN3kZF3wIHdPw9NTkIjYma
mYsDsHhNXw1mCqZL/BdSjXw76/2praBC3AoqC4k5yroLdueJZmRWgdHpvX+h
v8a721zYn/9eKzEEORFP0GnIZrrjRTQYFkZp+xkaLfwxmm8DbZbv0GCEHQeG
9OrDX+mb1V8Th03NvW7xn3rwMUtsLorXUux3pCGX1K5l2DRZb+9Y9toZxUvk
PW81bFsHr2rq1HJDdIO+kkak1v0oAzCvUPSscW6+goMCSfDnWoamlTu87Svr
WmAG72thNR3phIbdUolKA2JIspmXtzbJTqfJwDSSyp1mybY3cEv+MlS/jTH+
oXEz4csrHfdMzHgXyasAEVMNr9CtVJU95xlSXFDCQZNJuqMSyvKqxNhHn7cy
S8D4cdtPnrKH2bW8jn+8cMpTzHU32xoUn6WxaFXVYcM/9om5ELffX8wPFc1d
jI0uq3mzBbo5x4xqERd1ugvKSaHrzNsUiVYa+ya8ORAUYnm7V5CZutgfjctZ
5ZQtJMkRvMyeBKNoW0HQR7l4Ldo2d/f4SnH4vhPsc26iIsEGZ54eHx/xKJ5k
YcbU8akf0q6SQlrijz2u4Yp04VJaB1LMi48a09QqsU9dFPW5pkTk+5TgzDTc
UZhdEDd997/tLrBs4rjtDFTmGZRAcimywxUsw22ZUjziKr18YI93Vn/sMorO
phIH+lWA7foi3WbTK2xtNoynO3exby/Vn/3Y3B9FFHmGIBsHRJBoaGZ4Td2f
2sKEH6rqJmmppYel9zAlfaKfhk68mOHmttMX5p/YhTW5ZtwcdvbVZtmdK2xJ
ci37vPbquFWTRFt4QKnW9e4spmeqy+oAoDaw9kuq74/qZmPaFWycik6NgSEY
lrGCVPAAkIg6QBjRSu9LhMVID+2Lx2XfAThcoaSh1SfwHPw0FJ8JVU4Smvcq
DPicMEmgRXQhoRxf4a2nCIbuBQsbHbHtulDkMIiwykUKbiIVe0I9PIAUtwbl
Be8f33tlvO5wROJdgIusFCB0u073tUkZMJSF1vWfD87Mgrq+Q2zfuOSAjLVr
4b73pXstWQaVYqw8h68EO01xX7tiK/Va3z+2W6KjeiC8CdKsEELZAAho68eU
KKOd6+F+b3uTd3y02W9MMYnueqM0K0Q6+zwdsegEagh8OMHFigwhQwvPIDtR
hAsQdMLMoY9hemfQ7UGETkVTc+xO1QPxGlm7DwAzSBaP7JuREuQihq5YMqtA
LmTAqQUadAeW/AqiTZ1A3PvIXgLi5G0wnhF/anET94SCicDaRf/fQ2ly5pcB
AkV4Sk18IVtjEGBtV5kcumx6ttlKAjmlumCj7RjmLQikRtqd3eYkFpda+mIa
u5eNroASeYM2eHiU5jzjQ+1mGWqj18/HByq6dw4LSnCIA9vFPkELkBehhBZv
U+Grb7Fb2dcOZTatFqPv42PGZT0ecxNxPoMto2jyxZ2QmuVuvbugGjGV2kp2
P01UBZftTVy1KzgXhKufC5UaT3wu1nBvMRcdipGTaF3/gSkIsvrzY3mDOGhn
66dyh4Yp43ojKIsudbg4dkmJJrB0sDlBhrHnqNIZouRQOnIYwzsCoMxtJVM4
UdZzCzmAVupvgM9xPE4lkICN/NK0Q8pj05Bcmt8Pohf5xosyqaS7uz7QaXQ8
EqStj3Aknc/chO/lumORtqdmF+EbMk0GfrxzBtfx6jFXRPCfhaDwCUez3zXf
GolKHP5UufKwXfJzjm8z9RupLyDsfUzlxo2a4ZCKRgl+KNU8eiJjz0r4Y67b
H/o5/MwvnXLeBx6kXXDaFUztCXhssB4v4aySYc2KHay18zDkYJvYn27FWGd1
LKqEWDb7a+4Z0VExt6HCpzI0meqWZHUzIWbOysC4mnjWDeCqOVYzlWpV1yha
INi65GX47QljTP2w07eQ8hPggZOTU+c8kI+SXhk4e1xejrnAEySNpkJ9yLkI
euRhkc/B8FnkTA9zKo8TRQD4rvMv/oCcOpuM2oUPNTgSdigqFv3UBDg0nsL3
wLFHQFZthaKUeob3tZXSmfEMsE6C5THfzX+SyMDK9y8tKLKjRG5mXAFQRHLs
knxfbxV+x/XLVFikUI3OQGHzA5DYr17QTwXYJmva4WZcgFkdcN2jl2EYmIaX
HUWcqY0U4PIJH0lEKhcNb6H8pluvey4tA9NqXamSwdDt8k/OhW3SIMjmV0nr
h5s87oFcb+oCTTX7U+2dGgelpvLBTmky9DAIaCPAbc7dq64ROSvBEvigmVWK
O2wweVKcijwC2SUMkyZOkqHYtQme2Q4XJJkOjzvRdOM5nLFfl5thRvNZmceF
eq8dJSYnNYL7gJLWdUpjJyqZLBbS19ECCY/dUfzFnTApSit5s8sfkOnMBDqt
KhN1ml1YWaDDydTsExR4Oo9N6YEcQUFN6l5dPkVZlmZMfhXIQoiedPWa2vQI
DwndllPhtltu1BWJfTwuQivECgdWitqx4NCfh0KV8UXLT3EE0T9J43bubfqP
XBT0xso+cLmRfnjyq2RhB2pOzbPPCz/DU2Wly8oEfefimccYxYsI/CahQoNK
qA4pAhEE7PfvIEmr5h1J7agj8F21fY8NPpDbzBmd7ExqZjvOxrbjWVc6OAR+
r1bdGUiGpggFLNMIKxLWcZDUl7GdO8xH1w3fry+9cDKaJ/LvNa9ZpQZN279Y
sNWNKveQQlh3scqOPx8qE1SDjm90xKrxkIgdcrM1ULz5X6M09LW/9MlU5dIk
J8khgVktWDXVes5HEUG+FS85E4nY3nhaHTIGArwWMpo1lriKJwCfVFPUT2d5
O1ygB7M3/yyaqEUG1JkYoe9YLyP2I21c2M4975zpr0xVIzjNtB7KL5qSQHxn
Xwl5kG/o48agbLxeDFavN26Wc7aowc4jfS5IcQcPtuivvHy8VfEubfWSZzt+
PtKHAY6Ay6XPO7677z1Ope/pNvBklF/nFnxJuA2BCcWT8Cx3xYHTOL0k7iOy
X6FTNm7rbHH0swnd7h4cl2EZOzKESqhStbAyPXxqVQSBg/jQhAkL0xrl36SY
subXU/sTfkOgiicQSgXkxOxxoaT7xyxMuTR5nIKsStGL0aJ9FiqKz9lT1QUq
oiRag6hAqwKc2KPHnuGpcQmHqfkFROZP9tjgKmlOD+RAr4jpbEatJ1Y9fxPq
hsw2jcHcfdXe9jMvBx5PU2YDE3ci4iiKgKkg8unSCqG9Jcqu1M/OqLc8H50q
FIqvRvBz0LrNEetolUfSShRouo2UOM4RHHWbwG+9RBa3viuKiJz6deHk97ey
bGF4S7XCtV2RKlDQ2xh7q2KD+7xu/EVqBhyfAOINBBkaTi9t4NX99MNmvXCx
3+vRGshMo0cnmJoFuAVH/IAvMJcdlQH2Xh9207q801yogcJGbS/QVQOGpHxU
wCiymhHcKhCjmriAtG8l7723BTNS6Rpq3iT6jluWxPqAgN2ffp/Ukw9CvgIc
UUYGFJ6P7xqpvZazGk+pTM0A4QBb7quCjSCA5Xq131E5p+lnQ/PLAV0meO0O
QgozPG/xRzXOd0afJwwmI0EawluTsbpflu4gL5QBTfOmg4UaMo5uwel4+fna
OXRLOlza+GNaysvcr9X10EaNMXsssg7Tzi8SXbi6CnX/H3QW75ch1SAhg227
DmbjzccbTC0AqF9iSnlnYNyGjW8280ygdGesd2no7HQWUDrkIB4ltXc3ezr4
K5SBJbS0quoGVmW/CQCPfV/W81UYWanRNLkD8/SsYrwJvZHOM2KaoaZ/+toY
WHp3epWp36CgJ4q733XSBi1k/KuujUk8BruJO4hjPbSZfaygYzT7yjOgxiEJ
oL+WCj9EG+KU/CqqLbwB9GfRyPGh2wEKKPXMkrIxUab75lu8BuB+/fpytR0l
cqGiP0mS5qDtaSyMEnnCFQHmtQN7CTaBFJKDlbPrbM8AsSsfR179+i4lWjTS
UpZI+ICfkVwH/5faYqtUB2Oq1Toy2+XhrdCWlXFxAjI7XnN9nrJzF7dPBuXx
ViWPedJcDOTeeK+y5mdv1QnURH2qsRE0l030GscLEAapsqYWxH4SlRuGouVr
ie+ZbF+zE+6qyQEVE14ACe5S7vUy4kLFeoqjunXnsL7vVkAC7eIpHLTGV0ws
VUKN3T3c27sYEbgGb7F6zbeZk68/R2s1AIIjqPi5VSWFcxEYVs/VxTtHrjKw
Ila1XEU5g2WVeP/QsfvKZgm84jGCaFlF2T0cO9n3TP8UJlWRPb/68dgNrb7R
MF+C5JZ0E8YyXtVt2VTC7qMQHoij20UnZKVUXX4zS0P5MBwife9KA4wEyNeP
vwGl81j3buBvrIM4oqAlK0/uPou2RNeWHfE1+UNxg/Wmwhc+hSwLGhdpxice
xyEkZuF//6kSddcwMmmee8khOKlc7JpxjCm9u8e3fykOVoSEovrwo61zWmRL
ETCdFtsuROVZFVMfog87lpKhrg9nwxwF3ommsN/a1adZc8o0QNB/2JbaOvuA
Qo/gSJLk+tNfgK42PIqVFTbKevgQvT6CHmMxPsyqb3JCUzLX8TxjVyn2g51m
0cGIz2eATUlhlX5AlsvIsBvlj/T9D+nZWINGY3s7XJVBXAk62+X+RT+OWe8p
6vQxC+vXYqK9FQFA6vuzeEm/VRZGvo2qEYaqVp8HYnlkPLMRhDMnzneCwmjL
K+zOEbuAXWDKNgOlbZJFzmVFR5oHzjFXHQ1FRURQG0VPj1wkImdetizPnMUN
C8pHselyNd5jdzOX1qIrsItVf11OvOpMpliHnZ9+5NUsYD7xGSAPRlwKppk6
dLH8vBNWiUkNEaNdd3kMflBOR8BhvSo6jycG9wBkBewhQWlKx+PnDnCQZERV
MJ5eZTOIt1QfSDXd0XeHEjyuaJyG7PABH/wU7DAj073uYs7tls+wZBoyJH9z
uFOhxneel6RfuZMphhaP3+l6hNnRPdWqHG2glELuc2Zcbg9CZi0GUgRAt5in
djmHaLqD9TdmguHdnQ6HpAqkBsumgSPs9Q0wsIReVFnSr8XVj29TmGKf7M7V
vl0675KT7klzqzXLU26+d9JJxYBOWfg0JDOTXDRPMh9UteA9EowHWAY8BnMP
SdsFPoWIdSGHNZDSfccPGh7nFE/Wdh3upPtsvQfhyg3lKPqVrW9NrnZ/lWMl
8pMeZQYTbTtGXiuenzUjmNviArg8w8vOsUwp9Gg072jMtJdAKiyXYdDCvGMr
jKx1L2fIx6ZdwYC8+Ua/7V/0vmIcv2cX4Wa+HAtE5wT5tGVjQ8sGrQjaNgOn
VrD4keWb1PR8qlhS3WQidQXk2qTpeJV3woCbgNa9g+oYZwpNIYZfJMaPj5Mh
x97Xd6fbsmgR+ONuCzbAdOKkINe9bORfVzxD82dA52q/C0wHNjIj+T4knuze
vZ7FbpP34rCg/d5URDwJl0TBi/qYOIItoh6o9/w7+6LPpKES4eTDzoUt4t0y
BlGfEG8uX5TA6J+Dw08VBf2FVlfNamKvis9CtJ7aLQmq88gNC4FyyVRZE/qn
c684yVmCX3IFZDQcB8lpz6MZ+iqnenTyxsIB4RS0BxPMvk+GOULAhW2LBbuP
rXEuCzDflh1vV91TV+HyWLxSma7uvyFlEIaiEr1YMeZ0BcV9aV/0n48+qTG8
qz0DFesLh1AE3vBarWNnu1nhEQVXYLeSxmfTDGpYZeKPy3mAm9/9k2zvT9Ys
58IbFXZ1tm9sJ7b76Zzd3QBtBD7gAet+ntdLM0t663b7r6puj7RQU0Bn6ZW1
MENdkAaoJvbVv3PIMf/KyZwuS5PlWAj6uhi4ndcvMfhAPu4+8hvGjG8ZS0m6
hejuNosmDzmxicJSsaOFNWn6rpEFydOzl77oB0/du5ebEtQ5ytDNPExieClQ
210vnODksFugf3AhgnGZqZI7dUq+mwfdxxtupW7TnVcW3c7N9m+eFnUVWnHT
oA0nmRkzI7mkpdSFXNJ+SUnui50XIpQpJcurrF74norSGzzK53BieThZaVsp
58BYMzJ57tM047jWKW2QeyrTlDiVI+HvTpSAmqRCvK9psSgsWe6UoI650gw7
lhPxndV4zqtmtRB/lToZEC6CYNuRB2E50RVS6sd1RxLdT4xzCm9GOgUgnJhO
/jyRqe7TbY2BURg/Rvu+TZCjp/o2CZ3MvZdtAjfJUFv2Lbngwe6LtzRsivFJ
wNS5JjotVEEAA/U8IxcJoPGbeDUGQKor1wOM3Ie9vJpzSk44hkKLf5zB9KDi
isXGW5Mrut6vMzaEKvdqBcorYpTZ3uF8TacSXaAhnGx9GWnKV6t3wd7W9zY0
bJviZ2eIhj1LZzG6fDsMsnlAb86J5TkXPNyOF+kTS+kaFnqCH7mNygfSn3hm
ZvSsDGvd94JboQ5QtXIGNQU7f1N01TIsdJC4oOQurRvHZwllNPqRnlSu1Y4B
ArPKcDnpu41AlLeEwH13A485NFhO3TubwhA+2RXtvMUGAKDeC4F8dVBhE94/
yWV97GWzUszT8pZLS1iDOO0vV6mkskRPYbpHXZSuSKcpO11FkKWYQiiO7ef1
ifm+vGcBGkV+T+l7Ec9WphtvfFGav/MM604xefMQ8ScwUw+gO3eHVWoCrSlq
psCwO6qmU+F2C6EmrYYx1BJt8KxGND/fZa7bmX/UoVH4jLQeci6SLHepvbxm
A3w/PZ2nnBBMv/8OURbO5RTZOmraNd6o0oDCdp4xFRRor4wmG6svOBKKy8ta
FrQnaOlNmT3aay4aKWhSRto3k+z7UgbBQaUGxT7WkAgeTrk8YP8STy0b7/7r
XCWkT6pbDacmekYUpckZeTx9ypA3gVnC0blqekXHc1Bi2oA7X61R7pr6LA+2
CsSABAJoVRWTIdPZrCXWB1ggeR4cRoXEjTDsowBZNkLjRWPNVRicAM44Xq/b
6QIHObjaOjl40eU7VWCJBuZXrao+I1Yi3n81otIgRNReITkTfsAuFhhZGv7f
KU2iChDIPvYnw2+H3hPMs5AhqSZoS39xEtoRPyO73KagDK3w/u9lc43n6r+4
YYM9++r4idKaA/y2nT7gLJ7awXEA0ERupHBEixwxdxGGG+Yvl8b8FwAJ2YvQ
+a8maT3YUDo4O9+m6QPRMJV6RmnyR0J+2t872sjvQqO2vV3akIgJ0zRLDOCZ
bEp4myeMJ0qz3pHCYHlKTw+32AbqukLIQpwrc7d543+0xJBKUrF3Z9TVZlkp
s0Ct71qFjEpvGDA8htZ3zRASm7cX1iqKGmtpGznKPc6kcD1eREPkcHp5/u3A
ikSuaOt4xinJsW/3G6XsVkdnRps+SkL+vFy4mbN/xKzOCrtt269UksRa74Kn
CWsKNKHuhc8WGVNmR7p2tPsU4SCnhu687dDU2nO1ciSFwE12yfOWZblmPom3
MGfg0ykLGDn78TITQqwEHb32N76WEYJYlaEPS3fKRkYrblPZyhpgT0XamExo
5WGesLtLIkbCkRvNcTAoL09/Abn6vbc65zrJ53qAOk7VJT96fcYc9+O0pKOZ
UoBl7hxWmD2gnJEYhEO8Btj41P5c9GvoLZJpDtRwFsaZubatHSaek/NWmnyB
2Yb/dYEAmozrJzrHyndGB0NRi3YRPDKaiR5SAN7VAPhpYeR3ljfmirRAjXhw
5f+sH3GaGNbyXThC3ehe9Ga7zSUkJ83/SgaMxNIC2NTTRo2fY5L6EBjviXqy
upRUh3YkmuUpMnjyBmOrDRF4MIy+gWLD7t43FGdp5DfL3gSQwKO7Rn+R5Gqu
JKX/Xy4eT+ekGlnzb++YvXeQabJ3audPBe6Ko2Trt6Glpycjk7rMflTjvdEI
A8f+n7c7ap0zvS9+7cj5oOqju0sGnVcyCmoQkubJXIoBaVTXzLcXoYIve88G
2kHLuikFxEIA+VViJXJ5L1oAWjfsc9d2bLXJB0aSWOVBLnBasDzGcCuapWYj
3Ad+EmQyVR0uI7rpumypaHzrZ3uRSRGpWKlCK/ZCs/4ikiFE7ce7YRmvCen+
59x05ACTrIkauW0pTX7/qDTAjdreedW3tAhkV7BHA3Emuhlk5v2oBLNFly2P
lHkxplrvLnPMj02E6N9uwCYKDlpCpvxsdVSR/ENxqwHoBSfIm+iCcBIOij3u
yfAsnb1udMMxNbLlkOyTwRi5GMC4swK9oF0uUxCjiYmENZNUO+3tyBuEmtAW
Q19W+wd+Qlan3XP3P1H1/oSFUApGg6IkWRz7nrsTTJpL3BKLxShTbC7LYGqW
Smo8LsR2CL8lQTe7fCSY274U4DgLvSpJbN7mvnc+JbJaF2hZJTIith6IagOE
jzfGkhPtJdrZDNq40oICM7NSmhqTIZixi0ZJLwzbc1eFAdaNPJElIPg5a9j+
vIAALRwGkgRDtNIf9CeVnghfSfts24vX0fh5wMeyYLnflH08sx7qfx+QDAeU
zXpa4msOJ8+ZgKynGKLoMjX1gV/0Yk5+BYrkiHFQ1QSBto0zeHF+2plPE7Sm
0z97A9bsEo7Xnc3jCeYiMOJuVXmPrRHSD+ckV/kQtfWaIzUQQleee8dl01XF
KQnllZaHIZlzUFPPA+TCS3BhXpXPHJ0vAhcSTZ6Y7wCQd0VOpMWhv3Hfk+Du
uBya5xRtzx0n6IDJ19Gmh3+6ovTBs4+UoyP5EVM5qAS+Im2kYDkcAyAvB+t4
rhjiciug0frkW4eNcsaqZpWhxu8WEy0/lZ0wjmvWH9Ti81Sop+4pHW1Cuo+o
sveXmykkNAfkXKUYo004bdqgrWAuVy50ou21+ngFI46x3fNb2p4qCIBg0eHH
wd6xDQCS2UXnTRCbGQbG0b7bYSGRg9jNMtz70yGOwGOnQar49ilZDigft4nI
nWSH7nXEKpD6X5uYoexbfqQDXmPDyAjy4DwpDqp8dwdnE9uXUuhg2gs3mBtT
k3pZgdxb87sG10bhhi/7a4DdGt8Evd/mV77stR4SgoLMEsqZN+tCadt2GnXO
DskrQMm0CE9f+oz7qtENKV+Doix3GX0fnhauuZ9JELQvkoVMbla++fNZP1K6
/ZS0gMleSn6gp8MPcfoz3S1Wl4P/uX4OSWw6iSmdKuqVksUEUH4y/vQPdCe8
GcQ2/+6iNxAsdToFsrkDV56zTQZR+4atlN9RjjdvYTXzuTiP45cJBA1cAWJk
q0I3xzno61CmkQigL3ndTmN7whSd2QHLhgNPKVvhK+2XxFhA0nnhuM/ogyM6
D/EOCeNN8GMswJYyV6cPIqgmoVgr0sVqYjBWRRYI61VoxwxSOwLWyET9fCfP
UN1uCNRT4n+LdatPyBxIlP5Hy/t/I0fcbAdOH6U63BBVG5peY7LC4ZMD1Yek
Dcqv7jDBX/dJBPVanJqbtkAw8m1y1UjFklEV46FCTYJ+vIXjvK8jbEFTTiK+
WZokZ63Wi6uWOMATmgoPDkw85ssyx0lXUijAii/pXPJ4PigBiQ6OhJFzE245
C6sOFinv80K1wYf7TGvIFl6WYTzfJy+pWBF6IVh2euTk2aLvMJUeaO6u5KvA
qGks2dJcDrd35NzYIhDXbP5IDHkeUgj2eeZW68pEMn7FwX/n400oyzoRyz7B
ytfOsffGEaiIRI4J5sO0k6QeVMRLW22JunO+AP7foq0q9s1yfH1XMGEF3kDR
Qe6+/89/8lQ0mBYep3uKK9iiFF9A5TFlqyJe6PUJ+MbJwDbPGndUJhbPviER
3GdEnwLLF5J/0gabWjafOe7eWFpyq2qrNWzJ8U5AF+jRlQHDFXw6qa0fW9E0
nyM90AO/aTqo5Tn0I3azmdZGQjHTZXX2QfCk+5B1iDfmOaSMCzaxNbZKdVeU
JD+1oWyDB6YEI3k7VqkjzfJ3XrdT7QshYE/gDSwmVhdqcjTe5Vw/fIDPVHoF
WvCdsNM4BdmqfTSZTV0cfIeMFv6HSgpvQVnAUlRTQfc48M7LEAA29G+hxrLS
AgqD+VmIq4JW1lR5udGvq08KNQONIDJ5QAQL1bCg1oJRMvIdbwFlnCvvK3US
C3ERuDYTLvCHKzhtG4yHqnXjM8haT4l6vuopII8aj5Nn6L8daUM5gW4DF5q9
E89ILJv2S300wAdYRmBtg8VpaaEE0sDZt4SAx6NfeH0qoYDUGrCP4Xpn/KlZ
HEWorOY1sYA3iMGTvQvwcLRG3tfX/86Vvsp3aBS8vvY9mfy8q5kAror9YKVQ
sOROxNwL+elADEp4mAXV/tITRj8f0gBkJCFE9gTyeN5INyWMcvWcgc0C8zc6
oDKBZu0upnEuCKWjnGh3LLsJFthYIcYnbeR+zpJbr97JE84b97yWM6TycO+V
bPF41+gigafNvkTXBoaxWswclfc7sxS/p14pT1dw+pGez1LMdgmkZoL1T3KZ
kxw0K6IC2cCWg1fbf9q4yWo/mQvp3LCZlr57JOSu3P3BR9rMwJp/zBh0WX/K
GB9rWIZNYXZjyKpLykONpQobfmHCtxsyLACP8/3vjNkZ8AjIw8hSAbBiiXOm
3P6dyGwtoaW1VCgIAJxYgHjAA1cjjTDnybXzACvTcxGKLETHIY0dPGPhulIG
mcVIljGqQ//Q0D2xdY9akZA/gQ+dHcMDGmfSzq4bVhNhVSA3q0dQUvQmClAb
jTQSEAATufqOkqYpLDkeNqihR97n/UoN43q3qJX/2LGcxGgLFkagzz+gpD7e
wQ1mIRVOzXzbIB8IQBK3E8yPifKMfhF9aDzAQ0zDyCsSI0UNh7n4Wqb2Yi5R
sFvDEIQZPFQV5Mrhf6f4DlZ1TL/Ram6xHFdMIowaDET+FiQtG1Bm6RbYJRNW
Qaw79d+YiufYZLAvTdH9o61xezUAthn/+PspQ0c6PvvAOJR740CwV20QTkgv
oLYDoiLtiTecNAidIanpfngQpv62tJhNKy7rmyO0qdzqSV/IC/EDqBseO4f0
LhmPhttXFnMYsBcz1L0FW54s4Uk5dfSyINBIbt7xY/b7PFlv81kspBennqNy
PXWc7balYkWAfIOcdweIVm7jOb3zGvqAM0WEFcMa+wGVPfQaHyvnqjVdaP+h
Ky5quzeJWEmDBmKlPjzxy110t5nxiakzqO1KwoezhIxEPuOt9v/w08PbTbO4
vB9Gw7rMlKh2WmlelOAMvSCGRwgSjcL9rOmVOPzTmzwsos0HcZZeSGl1JEco
iKXBmgKI3JY70R/1H9rlYD8js5m5Bg4mMMsiyFkUCAoX9oZL380xVEDNYGUm
8+YsSj+SYzoe5sonXOUj4Cd2ME/4JgP1qtEP9vMoAYaGjd6WpZg2QfWAGiEv
Jd7WQwjo4ohP1gzHdQ9QSaflbwfqcKdkRP0wV5YmjZ6GfeV2TzNr9HzZEMm7
fNJgphOEFJw2Bca2tqczZUdgPVySrZDP0/7I9kTJGxzJps4/xqdNYHLZ6emB
6qRz6/hovrBRPZPNO86uRTP/h/aD/JVFeoTbm5yDFUzHNMP3otVA2VNyHqcF
yQ4UJPOlREUuVuZihv3Ru2y9KbC96bxUrNAVYoeByEDRr4+0v1WnVQP+UTGZ
5zE5IHznxu718XIaM2yXSVuF1C5bYTix1ptx0iHur1ThpvDtlqNBp/Lho0zS
iRxPmiQ+dtIwNrVLrC2PUmU0rpeay6cFKMF2ruiCWrYoq/IHlQNUQIrsrVw6
eHBTFykTNQ7QubXW+fFhwbnkWKp8ErQzVzi2KluXLjK91Pe9bBqO6xYCj0mq
ZY/B3Z4huQZ0ss55gx7eA8z/yvPjZMYRZUDMxRd+JoSi7prGmgEt5XyAyozU
SNWIkLRG0tPdBTdVYcCihRLHGyl1K6uHl2oQzW9HSbXvBE+vpxkPt0jlUM4B
HNQu8BVy++8DawokpGDvIgz8DgDEU/ao9sTwduNOB6Fd29IjxXAZrsN425yM
f1sKpKT+8j6qQ0BGv7HbBcKLgdYdd+seboYlC2GUR1NY8VhG+nmjPEh/K25e
xBGCDdeYucaJFNILpZwAQ6sLetiliZj69DlPeCGNF54/gSpxJluAf0YmkAgC
dpPhSScDq+hRsoJqfDkUSAc2/QwVuJz6fqgfUj1PbYKgTa9C0wt/+vBH+RAC
6rgEGp/n89xoDbmy/3VmiDYVqK2O0/kIYH3Ge9RYFQehoiNSKYrYBDBNcn3d
7qCy7flgcfVhRulUzoa0MSfcu5P8pWTWiYSL0NxLcGEkLq39b+ORQRTuETWw
nshgdr0aGKNXBldg9ZrGNR1362GbndA0JM3DWSnBYXgJ37eYM9obBXGH6Sty
RvkIoqS5Hz9QPMNocQ6OBUmdN3aqnnbcXIck/KcxUQaDLpccXyRgaixhXo4z
ZTcl50mILeYTvUt0cQyS1XAoiORgdhIXCJQX9GL+hj5IhXjPLsknNgfjNn1i
sEYeUonwEISmeCP+bhSuqPKWjicEaxrhWpy0OFlZZ7Tmoe4HT4NQZkVg8Jg8
kOHYC4AVeGybjyCUwjvPtpkkAbXmZ6oBBTgmai5dgvM2JSUye4B+CMqj0O1a
fhUpV0Evegc67XSFCo9MKFUXOJYqzUdYpOBhs1HoruZi9qN37AwHVy5LuvlO
vnZuj4TBzYct0OR3w2IPq9vLj1L51gT25Ocz9edbGMqqa90D7cCW1ZoYeIOP
lTi/S3/R6r4qsbY1uOWDCFfRJsGyTLkezlrDBUMMKPr1NaoBv/8ACEYF4d3k
lDWDg1Sb2FKyBFeyEJ5Dj+zfyJc8DWZbg4U4y56XUCLq1vASsWWhhjV7efub
oT5ewXGC4UKLYNneLc8Y02EHPTXt3D1ZAMarvv+qhP3W6+mP1lxqKB8yM/gW
notXftFepmBVNsBlyJb6dJZU0VntIWMJZxKda1tIuntoYnDNbIVaddXrdfLm
JtnaiNU4gOhMN89VssqnVSqxVq6ipyTvv6/5/cdfxIl+y+RGmaVJuOw52y8n
uu5BD/4AJeC1PP45DgsRUsEftxnAbq01l8Z5VOP/2xcc4OgpgdSDSIB2Xy/o
G4Azj3gLiAxk7NgeYQ+Tx4gTIAgR4Dj7kfZhaud4q0Qw3zdN4ActD82CHGsW
aa6HtaVRVbEdrXRMxPJKpYVzmzb5Cd/ozt8Ou0O40lsc/hDOf+FUA1x00GxV
Ii2lbQGh6+VdKUOXnbEIcLPn3waNGTNMWrXtf8UMqgySyhMHGHyKlGWAnCWS
HnRc7TxVm9eLIW5NtOroJqXyGMV7ZBUx6pkRzuA5/ZBSrG3f9VNUfjZ/Enr0
Dln1+DrbBzRCvWM95DMZGAO1NNbzdpF72LEQeXyvbf+3uDpvmIrMmNpdvgnb
QXaCFuNJKWcNBR0PNttk/Nl9oILB4n9FxD2+8DQXFb2hRd+snS2M4jrWnloa
vr/c3Hr40NW8IyuQJbvn1VmjVTzZpTue4RCavA9fbHtyFUWqNDaSrZVJssXN
PamnnMS02v6j6QolTX3AaY9VngjEpvNHmX2n9ta/vfpZ3b0y9fUIOadW3W0d
SPe8LpswuB/Waq4eadnnTSAK4ut0wY2fuDTSML2XxLiNWkzkUnNeyzUgdV1y
i5zbA3LQw+Pedc7iYgt+H4Qx1fySoSlLnc8Fo8GK8NgxoPnPflJWbjrKS3Ql
anKbwIJ1Sbu61/oUvyCfLaZRukdJHQbRMGYciJnkU8t11mgVMR8yFYGvpKT+
Z/5MOkl+Kbtm4N0pbH8f4WRtywkL8u9BRJDii2nFO7HO68PJd4v23Ojpw0zO
e1uKpUkBxaUc19HROs20S/tD16jInSipfWWQHcpKEHEvZbvZWl/jvgsraQbh
bBI66aPth9d04tYAvOwlkpxfD+ZvWLRTuqixxekhUtJzaTY15Bt1bHNJw9eN
Nae659GlKN+t2ixB8E3KVy62iDdR4oJwzuVQEOqj9iiE0wSdDpAi37XOHirJ
gr4FiOSqTVCapks6j/C1BcERSM9119ZfcmPhXiwT2AuOC4n8nQUCKB51Azec
wnhNS1uIpmlT8Xa1hrjZTgMB50HetTavrTv+KfaLscc8VIKcWa6Jz0AjBMR3
grjsMBIxlzePkJCroerp4wjZTj2OUca4jXrrHHf/b9IYoj+8koSuCcYtLdkC
XTF/+nyTH8SII7niRqgCucFUVgHzstvCv11AJq8163BEP9boKYHurSVLGgFd
c2C/a3FOjDvlmnwXY6UZ8RGGWtDX78S2uXI+XwaG5sKcxrAtiLvm39Bnkmyd
d5kRC/FqsQWJ5Jzz/9cI/mqLuGjsayYC1BmxieEfJaTantF5olxRvloriWz9
kfVhXeW0UYF1JOoMbzIm8/Q1WwLZg/qkI+wKtzzGl4CwK2I/weEvh28JZjcU
RYfgmUIsF5ILu20y4vjVfLXSNMjDW9PEIgn4DcCc32Cy0P/GcL+/IHDXCgx7
9VwNmtFSeVfcyqwwW6fMvN0RweY0QaLiSc8+XbJBUiRxvdBWkAsCMv8AmtHs
a7VjDVdKUZMQBU1hRR34uHugfX3H6/vKX7M5n66yJL+KbLLrR4lPNrOM2Esd
8xcsdceYKYh1ovAVI5AqB4wfvHVMv9k0EJSYWBZIRHcEfDSOBWmxJzTP4AL3
D2+YA7iQLeK7KEXOm9fJkLvj2iY5kpm3WYD9cO+k+jsgjqH6NMJR0zGSK2hH
z3OhgFeZPGuFOTML+AW93i0NbswT9gPQWjog/7YHU+0MINSgDP6ZnRKZbkAp
pHgA9H+DAKLZ6+mhDa7lEUe89NEdGv4RaDLDG5QCZshvnUFn08vKm//HfKv0
1zRWl5uJIVOM5kpWIuVwp1QjbEujZySt16UM4kF4M6fKX/SWH51i6Z0AvejY
S6udU6nIPMMtJN0NKoVWnu6S/cb8pxjln5Dr2N/RKEdekyTD7/ibwKRcHi07
whTBKZE5GtpVs17/YRX+mGqyd8osRhWFgoGwhlQPKAgTUuwI4qkZmWS7UxGH
vcTx+T3ZGRjpKux+e7lMwUm8a0EhilArBfCoB71hSPQLjXA1qzOHoC48vfgq
WVgZ5tKnSxNkLljtz2bRUha7cysiZWwbUupophvrDte3mjHUzfkBLGCoBSRc
slmU7qVr1U6NP+9gylnToFKGJ2msovH/Z43XawTcQTIXJu9F8dRstc2q0DmV
Bal6GZ8TSZIIuDsSiHzFCValVr8veMVQlWgmMjEmbuVd5uaiSxIV177mX8FD
h7BqYaAHRSZEeIr+SfFZc8/vBqWp1847FvsA9p7nYg8P2bmzGpH0OihXZ/wF
oW1Jtd4JE6FnFXk9v8PY5GiiRiE2ChxfeRrc4TVaSDzP7LXkdLtD1NO0evd4
/0APv3oPZ49uxp3YOkGrLg7REhKOeY3i5I6/T8vUQs8nhexGSeMe0FfRV1mI
H7uXAwbDvcpSsFaZ9uubRhIRIrW6+x7a79KQRf3t4E1KfDcgiQCRQs/un27s
H7KrgrgBQX38kioZH3TIQEZ70p9fD/WbFcRyq3Z1vEaU4FeRB+gJK2pr0739
SaV1XzQD4CAquxIuUzgTewPI4aAjLoMOREEse5HlK5l2QjNgNuAing+zamX8
3zAeS1v9wAumG/hZ3sVJa6dKUyDNxgoKtFv//soEOQyFua3DfCGFcB4ELWL3
l/VZpVfyFzynkwrNDaLNyKGpwhtiV8fg1K0Xxgno2ed64utqQCGmHqGoaP+2
XB2mig3vCw9aGOasHeULFo/+UMx57XEBP5Kys9v2MIUxocb8S7cE0ZZUkj+4
hbQHaXXdp0+iqiRNwSwUmfInDdpagKlOj2pmDs515hJREVEf0RLQzUDTWYwX
+YhkesB++3KSlSijcBhynyIijq6n9l3Bss/UbBUxvxrejJ9/+t+0ZbVx3tZ0
RwAWQWgLi55Q0M1Uu+BlWNtzm5cVNtM0k1OeV4JlG23ek+MbiIzaZL7vXw5Y
pfLkFYNDAD3cMDYmsF6fv7cZujYqjdsV092G2wF827og/Rb4zirEThcjauB3
ZtU3bHSk2bQNF3nb2IamswIdtxPpYh1u5Gp5MMLvwVR07e/9Yz7sHVKLZn9d
wMAxlo/KczOJdImuqtpcJ4ipR4sVsfwH4xOa3ReRnz77/wyQNqECYH46Ip2t
KdPkSqu0z2YK7FYYZgNwaZMSR2gnAJD2nFzOBs0ksBXwR/k0ltH2zMVtCNNO
UIovRO3T5gL+wShI+jFjnq7zG5QaH3vDlNq0XciWuq8Bt8ZXsmY4DbOGhrlf
26WRStKL5skyNvLBB0CfsayyosEvnKI+6zLoNX6dZAKcb3fdHztzuX2GF1jf
CQErp0vi0APDoWgFNZbo07MO8NT7BalTlWaNxxzOSk8brK9N4NyGwTJzfdei
KRd4TbwQPEG/YK80CCjex1zA4uQOqEika5LpzzTDDL+fqN7P4/l5dB3zAmwW
7Cn0fWjj7aSt/bGgWO0QO2qSKL11uVG4KZqmEY7pDt6szyeJoxfsAiNn7iZO
g+vJ6OaQZfMgq/wPuqVn3p5gUGsAWmtBi6guORXFDNWd4n908ibRb833LKvT
3LYa2brNA0tnoEb8yUDobH6t/Om28ijbrBn9GHtFfPXnpnKy7YovkB1HME3u
rmcjf8DhCByon/58NC4cu4k1zE7TAOa2telOqBfbDTIN8/vCeb11bsbcC0dj
1IonoutA3zfm3Huamt2hNv/rovvBeTo0L/qQlPWamdi4J/BDybZ3uupOj1yo
EH1K7aS4Z9zuLXPHph31irKceC4m7dqYxnD7zg8a8gT4bDN8VqTTuB2LnBFQ
WWvytBMXxzqtq8aWE79Suo7NgWVhVVEgTLZnaRAC1VsX2gEqzHUlVDMpZEa7
+tXN5KiyzfonGkOHIGbKfxkT2dXh+AgPv5ybikbDLuTQDS2sZmVKd3/qenZT
GaHAd09HWnBJbSEmvu1CmO3sewhaS7R4df6ANKU9GD4Z38/N5jvb27MS3EIH
vKYJ5kC8Btcze1kO9Z23cAtUAuJCykE5Pzd0diM6l3ZDuUFpqfWHOmSXXmnu
AZ0NnyMkLcrLmDrGg/8Jj6Zl9qDcMEHwMskYBxRUaNB/ASKIj18UluLF6epB
+QW8rUABDDn+kP5M6GPTiN/hQU6mZtOPLHWGARgRu2klavug6cHnpmr4p6dH
uT3wWVZOVjAVKVD1x05ZmCQ3udxIkCTU4ND5a5ox054FhrxLuvoBHl1g/pO7
NxBlT9lwQct5axb7+jyrfiBNzGiR0VufxXAJsoPexrlafjxL6NbT9U6qxkn/
hc77perscSPIOQasMl69XLyUoPHUneLDee1+lJr7OaxZgtM2ok5umABng7lR
RjIfRKrOzc0JPj9qkcwBKOWt/rc5hH9y2XCN9akhcL5rL39COdgIY8HaLlLK
AZlXwTkxPBjOh0rPmRP2muIHhq4PeqyTCIZbClHrCHP3+Su7WE8UFE58qacl
60RQy+UhAiusKAxiGogBZ8MMaUPsof9WuxiEGUUBaBqBTwyMtRMegp7Ff/ss
qULLdxU7B1RpEwqE6dHGiyoLzPoTnotDP1gSIUmA2ptHeo6kGXe2BPZBTRC0
ef6LcbJkB3pn+8txwwR45SUoWmB+XENUL2qtwj0fJE6PCDlmzweHPlRPdNOW
H2T5Avxufg1su+cSuBRH30ambMaoqBKS1m/5QVpTV1RRQvkmj7COAug1J6w9
Cv2QQrPWfHAtPmVd1IDhsbo87SlPVxjSXZCMUqmsOSFmhQ0cg1gAZ4CCqAtY
/py3mYlZrxXfEvgdX5qoXaZpFW71Mh5E3YOdX0pZPLxNarybBLC6j2MQKZUx
R70XB+iNGB8fW2pNIw1NJc5iO8gU+ckGxCjcRJEe5Owdgoq+q9lRt0s/UssX
Kna856wEAJWl1/3sq/8Q1bh+ZkiOBL6IKvNYZjBFCiq36LKaOEStZ5Fr1Zok
nEdi4PgXiLsAeJeuZ+T97L7sHQQef0BJ+B4e1YtqlrLQYgXrD+4FSmAgSHcs
z3l4ihQ5jM7ZXl9e/fq0Orc12HbRJiPBbRxymOPegBHWQ9d5QzMtW/Yeuu/K
NJ1d92jwG1J+ZmZZ+AKpZN0YqSFmwRnJXx21W4237RaMt568k/HFzhx3c8ui
AJav+g57Njuoi3CJPkdEj/ZkZ1XPQ16bCNQ65qlxwJbOUKg1FzVaIdQkM+CO
3xQM+ePJDWhbcgF8xTzhOSq7e1dDnow33ZUejVCUssKkYndyToxz4IhasRMq
w+KUAzKO/EKWIOCbInMAS8Un5rSxLM1HmU/Rg/EcweZHeNv3ceGckgzrGvzh
ndWpu+xu6zRdRXsStKjJvW+MNK2RgpXKflfZ6yroDLTM2Z9UzmIkz9/DOAZr
xFNPe7VnYqBM9JzkgE/pgdVx4vGUVilQ3zPjy+LjfFKt3i519vrImEOn4/QV
gHYlsQbxLaE+gliVXCUsILymVyXaMmWjSSdZVeeHvBOwoh0l8T1KFTe6V28E
bUEAaDnOffKoUQkWTZt8sjMq5/u7Qn7LmJTXvnBeYFS7aJr6Epio8U/Ks6Pe
WA44gsHWl0Vj5k83U1HrdklBPAi5glGcfY18GKXThCGarLWOaWtQARJMrAUh
QOlFkUI3/P46T+v2yL2p+fVqTzrMS46jdqzHYBndKxbzirt8fZO0GprG7Guf
CbhRozK2tJaZZkUfrqG9O6P1121rb31up0ShNaP61iMBl+fZSWDY2iuVX6fb
4sTjgLF9Gm7FK9be53K2WoKnUibDQiDHs71JxYNgZMsonsy/YP9Wuzws6ktG
msJPWXoeTcp8ELnzlxbdW2x504Gwqq0GXzHxdvQaR+plA43YYN9joCtPjOZk
Pp96I3a7rjUMFRXPia02uz0QYMfisTiujjyPwTGPQDi7hpNmYTBbnRJIutJp
dRFPZPKu5eADxREOQfZLmr6h+v2NPJsX4gx2DM2qUjZQ43JhLSt6TlJhgGrS
iONsGV+cDfGEFwKmxiEawYk0UGxNIvm59u0rOUcLSWPQkE07LxGMvbR1sgRU
TGM0v2TxSUsOeg/g+rwyxksH4qe1Gu3xg4uyFRjbHKk1A/HOqLQYQmWbXtb8
z4zT3ajyYUi3fetMaGD4LjoJIwEkPI/RX1tAxvgXpi+O3QN68R63vLm6kkVg
6Qc+vl/EatA+sxMtE/TCR0F02A2pyKa1RSm+i4JANWcI9/NbGEQDBwLCCFKF
r+DecMfbegz2+D5maAeS/G4PkTOeXCtlYTXYJLDMBSWj0dIJv0mVtD05tFcc
KBhicakQdVr3kD1Ai09+PM8m3oncQkloV6dBmh1vI3A7gu6gfYADbPR4nCsh
Fx6vLl74jJKk781q1NIvRyKKjynujAzITfUPpoFjFSai6RRZsBKUsVgL/V+y
NZzFkvAWSEPvNr9C8jUUanvbwriGkp/1bo1hvobGASRzvlJRzex/HAj2hZUB
wf+ATHrOItzpopB/itQxAm5VHcPChfg+N0rx3vH8cjGRyvpKa4B4a8g984uP
nu3iBnehdFNrbaJO2/p6XYq90uCLxw2HcdxJ86Ak3uUGA/tohe6RzdXHdmr2
jA/BvDUByINYUwPndXZFVSqNK62n8nLTCwtvYZEa7zpaUVxsGJdlgvB+1/Xp
dkqDp/B2Cw64SKpAMOwPZXrESujqa5tW5iUS6yvww3zq2pTIsNfcWtFNBGAs
hgIl9CS0S5Q3X/NngU9wRHxr9uIgy7RtHGqn8aAxa9exQGoGpAGLrCuxVrYa
l+nM9VpKIjhAINltS1uRQefqOvOsgsnzsS4WsmebVbBGbT5C11F6uDJlKBK5
I7l+QES0VeaTb8Q0frOf3SdxDAeJDC/+okmyw0rWFZKxI7J4S+RWqitdsl2m
wWeYJgIPoFH0Dcq2DRSzK6a0RvtnwVa1JKA0B930fSFy85OwhxLFeWE8Ym2+
2rtf1rmJoPSMTWzdu4Nz9Nlh0sg9kyvvQubz8hSmeVxHWRwF5pToMXLR1Em8
VHbO1RAVp/EngU5+ekIow4gpv2SVBe6bOTnV94bYwqVg3tqt6opSJ6mpvta+
JFTvwS/xUV9GuCiCKuUTZyIS7pRaZ0DEOMFxHqKO+mZh8JIJUzCXxRtuiDeq
oemUuiINOO6vMVqAT+LkEe84Kq1O9h0gan9L71PdBG7uUQ5WF4Z63ztOAv4a
GoF6BhkB8TN20qXNdT4/Le+ml5YqYG6s3BQpkNlGh6fVE7/9UO9t+Nb0YKib
HVGZb0oLMDJSF3b7yQDs0HtzOCEVtcxhuFiqdrHHTNATnBt/nHIuCs3hJR1+
4jR6lRNe96k7eUke+2RqozRgwISBPb5vn8CdKU3DXEKL0Zab+gkvGRsGMZK+
x1S7L5r3fj0d9KMBXBnTZlwH1dWxK+MdhnZ7gRlp0uSIIBNDZz5S6MUiZUx+
mG1XcUED1e11TDnoylExV5cZgUf38Q0CrkthFZaP5TNbNZVJqUEWGlMtogq4
CPqqoPg/tsUehNVGHPsnAFhWupCTco7i/J62wCYR/tVIxeGg5HBeZvmi4LSg
CmadDPISEEzMhdgGz+0mGhJYSzgoEgw4FUOVdgXP/1/yIrZpzzh/reT2ftyB
j7GcTEChlHUCvbmWIta5KoLKTRXCnao0MnlDv8bJbiuCK5FgzznZExx+eCVl
WAX/YgFzBytnUuM112G+NcobMRmhc9/THPOBUI+mdFGClZGZNXSV/eghDgqm
d+J9+UcUre3X060NoYTKLCAMVa6wUXl5K1ggpT+jsndPfTWlsUldZlxFbp0p
zT6ouLITC7mzYLNp7UnHMjx7MbxTt6sNaGTyBDfNqC5gOfw/CzaMhkbIhTvb
X9tb9U64cDscs815F4aWKAqqNzWcPLRayxX3xe2W2xD6zAoC3pgORHu8YMg0
IIqiHR/4Q14W234jf/pBHHXgSrjbRcsBcCzHb1lS6cB+UBAox0E/ctD2uKqV
3B6Bcs0mHB31Bx3kQomoQOOkm1EOGLtcfrua7fRj1R0GMc9ag8knBiSVY4Br
qTxBXuYOcdIur9pNEXn64zpv1c8M1IPqa2SmBRC9F6D/viYTCfJAQQqdHU2F
BW/wpAnCJcOerJPlooBa/kb0KUEXxInihXeXQ2suE9yfFp4rAp2kJZOGBa2J
qe52x87DFra01nq6OrcvnulmzYuT/Rf5O9pVgLMSF7trBZ/VtvmAX+zaEpMd
GIishHcHl0bWfVO8SJABrD9yTnzERBTmyCGY7nP4cG+QQGoiYlWxsfz8GiC1
+ypLzwlYmB3+YbPivr495MrwR9dDW5QQjxUkoaKSKIefkavv/Hz2RrqlEfTA
ahkPHquYuk0HtZiCpJxHJbTYHIIIKfBKo8JFT7+nLTTMW9bjNfxxeoFnkytj
Pu+xy3D1V38pHOvaMumQqm7T15lutcKB4Z4rMIAh1wKrq7kU1EjDbGJpp3BQ
hAtt1IOmZqKX7P6Nir1tUHkp6dF5xaAPzATijpbamgiT//BWG8b94WPkC0Ui
7CkwjSEqn7LGEZ93ufsRHOFq2Blbkua8OYi4R68H9PNNymfV1SVXhm/xILdv
q595IM5O+64ADFuUhVy++tT5wBIrYX3xXCRmO9t4CBtpizVSdyjXfoGEXFFS
B8ij+AWjgNX7kzbD2tTX6/1+0wF89DGU+SxKcMhr7/BjhoQmw7EG3BEkwd2u
Bu2UYr0WH3JKayWqZ2QxXO+sR/iVl+xjeUY3sRfLrt+Qj/Wc1cX+fGJqyVS+
j5gHO1QwptEDTIPuCTJEZEfW8GjZGw5v2zA2intss9uH6pJ53DjdOBkrv/kZ
zNdwBq611JfJY1LV369mar2wxu3cVmjS8deBCNLXInHcqt6hMji7BC2GYdHN
SK0a5efsYPIuHpVEzG4AEQewyfmATMj0ezRXRW3Wj0XI5EnZVOPK7uXxWTQP
3Ss2kiaTRtOc5YKv2CprAMC/1JymhXHvBUgcFPP9y6LCK/N/xFO6ig2aFOoi
Z8frrQkHqfVsEw7hzbZpGbE6C/fMx1muMoJhDqQ08pRhvvnrZ+ET0Id4TedD
XuAG3M1fjY1xVNi3TtUauZLoy09umcKQtwNMrjminT/2U0OnholOcZI8FnLN
4WPXRmx08e8qKRtOqlH2XCKtOB2+5VuKubCKa2pWP1x75FsIgOrpGxEaVguD
J4FCylHB+mqQ4jbcIQVBzPoidsDoTrTlJ6RkVrGGAIpK/y9QCTS4OMeM4vnF
QSi/jg4gKTbVkhJLxbD7rpRBe1QcJjRSbSkiAUFGXqw+cpDfiSct6dUYbePe
8YLOmYV9vX9kV7aOpf+5uwESPSi6v0Z+8+BBX1EYEtxdRV7S/PaNKOHtBF+6
jihQpXON2LNjUBn2qbjOOw+4A2sAc80pQxTmhSwctTwGPndlpGLqBFg9Pi1W
mYhKWIYE4kSI8G80mB+65+sXuOmI9I26hHfEPXwOlUuY5QV4N0JbQfEzDp2y
Cp7+DeCDASFqh+X8l6UkUleKvKway0g2cEZ2vWbRw1SmrfvrCoIdir1xU2NV
+FJ5SvR15yiYrtM8/O+tnWM7NrakAKMmsN7r1J//beG2jWEVa64zRUvJWiBo
lzj9yyCbvDWKLZZtwA+BkdjK+pHswoC2SKkLuvQKaFlBGgBMlk8yawaMKh7H
wMIp0Xh8Cgz8IJxEyoELAN7g1UXw8wZnp0rpQK1dAVvpijIBV8WV9nzf4fP5
/v7IFriFrTTMV61JGUHbVvLrxZbdySnHpxEObWXobqvGwaIw2ac5+1E0hGz1
tYeVKogI2A7KZC6d1YlPDpuIVBZQL+XpwIUJLybhPmHilnbyyEXcTSXtQoKS
h+A1wartfO9+lWp7dJY/ZEqk92eG8wgd+Y4Ao9h95zd+VsP25iaCzh9C0t0Z
JFewqXdOwG33wVhuXJZ8Jrv5OWyzxyx1rLjRZoCuJTTcr8R3VREv3OvOaWMx
vWF2jjLiPKZFSoyGgaZ5qBpZ+spwceiXoc3FN7wFCWd5LTGHPrVyhBAnqYJ6
EO8kwWZK3nb4ANWEXFhmh1PrNiomzjMrGRX54hyBYA+8yaeMBozP0dT/EGZs
pU1lrqFzQYUCIC3bVLQiJ8rAEuqb8hcI+2c+bS8KKdJpOhjw/7QQAki8DWSI
Yce5qr2o1umum2yREXav9c4h9VGnd0qeKZ5C5GNtka2dgZYptmr3nMEwbuBw
E2XQhlEmvkO6N+Vavlu03LggtORoy3MB5BMpiaBa0Yq8MT9HCbmJ5oxDJ+fi
gn1rtU0SAgr7W+XtXdPxRUNoPDfdJAT8AVnFXn+F0FLWThV+dU4i/q2aB9Oz
aSUZQ8eeGFg2r6u3bovyAXE6ko7kvd1/POfKbiMb77JeWGqM3SrF40gfL2ME
DeJEPqIMv1BqCmrcfDJxm8czYc2npiLIBpX16IwuGl0bpu/5Eh1sPC+1UpxL
C/kLBtBwqLRXVEuN57lvorQ/S5Feghq+oh/9KsDE2Uhd5X+/9aZRbFDHN8GY
v4n3TXB450tn5+cIClCClcZQW6QIp/z6iPsE449Ek43HUTUlL52FGRhhKfSt
hP1doP5HLQWT4YV3Xbsyg449XqZdWHLGkKtUTEN9KhRfyEj4k/I8lWku9i3e
NnsFR89EfghvDaqSCoFyHcVsTuPS3zNNeW+WhGRbrn46lSpBg6/rOoIM9/6p
KJJyDnMtbZ2U2zYJoS+b/alST/hghXE4Jd6q0kC+1Idn7QO/al2F/JAisJEr
6CxS9MS130S5pCUmjbtnlksRCXEA8v99A/fN/qG/Iae9honuyZvkfMRMUV9v
tBhStkZ2IObqTqAqPoUDp+nVu6rDFGWlOg4m3VgWZ+0AQw0r9YRdK7KG9Fxi
L9HRE0WLZZIGwRaLMCcl5i+abM5r/3lDyqb8mtmTIIhQzeRiaw7aTik6pdi9
CtUhmlsSshzihgQdpzeY+zdJfG2T6PPEO+ZbokVgk0p/YnRLr8mPby9SvEvl
5zhGRzet69oPSFyAlVDBHEACfUIghE1Io/mKHOIYP/2mdsHPhUYWzjwkGc4t
1qC62jtOJd+VP6XCsQTdk4YsCp6ey55d9iQmm4JR0Rr7LG61IHZ35mv5dMLK
lz7KfO91YCfXwCA1tntRFXDISYfm30LFeKIpACt3WwxcHARUWX+xBjfkVHyM
DZoXupkYd7cMxwcs5OHwKkdnjRHskX/sCb/ra49z0slvUewjwpM32LmhhzXE
InKvu9bs/vvgE8Ouf29Y6Pgk4S1CTM9FaEDkWrzmUg/x07kEmTL2YsdwmLC/
8kyWdDKBQxnG7xKCbcEqYXZ8b27/TPa+8Pl0UvwHOBsBx39DI5tUIKO7RlMw
s5Ff0qJVV7WyxEAmEzJEk7a7F8rv7ld9g1Gr4QKQOXQH5GG6OcGzqFuyJSXD
24zBRnK0WjuwFbNIcYCuelLN6PgVXDDJmwy0PiCTGZ3nkKb2nSw8tL1YWPSS
j/BdwBz8wx3LAkzWuiEsR7eDtns41KMeV6DL8nC1JtR+bnHr1ak19I8pukmQ
jMRkkb0a14iynPzs/bCSWrs/4iWdbNEgINuFc8rer7veRtgGeOIrGDqf2bCn
V/zd1o3GyCwaMlfeZq1fDwvBc/PThakeV1Qmo7T4oYcFmQDTczxWZPuakcxj
XF6lBCJraccQz+aO4akGDTx2k/ygZR6w1W4Xf1QpDON8Cbm7eFwyKvJglInC
sxUL8TUGbQq+yNUVK41LaJAGGBQy9zVKsrK6h6bdthKi5OL+jx/udteQ0VcY
C6RxBZ88INvyNn5UPuw0GS0nt3C4if/qeIu3rjKjKkWGSlJWbM/xd2kXZYco
v+jafqCFqtbDY6p0q0XQsymehXCnwljAp20f8PnkyExqMGpOKukWBc0MKs+D
MLYmBD33yaOjuxYm5n9gt6rPsMdmXU4zeisr86oPPuE1cPD7E41gk6dsRSmO
7dhNEj5qfBQxecnLojqelfTO1DQuYXI+bauIb2yg6LfbpCW4F2c9ZGUahqxz
kNmmk6ODWXWDpFwJ5B/aefPOUzrtl5pgoav3l8V90VCC+EGzvTs1t95XHyIB
nwfugp6/6xOi/ruNDEOvCt1f+S6nOYN9V2rp0Huu/t7IYy6R0TI3ct/GFI7i
CvY2wGBN7ziVc+TNeK5dPo+FgTyfSb+gmFclvO0fqwoDJa0rQRvbhZIYDY7j
43G4e9gym0MQ9m05s6odR9n4G9AhV/LsCL1q5kVBBci7Lsgov5JkqmWXewLW
m6hsrCaEohB1+K7bxA+aTBBJfIS0ps1s8VhJNczHO9T44B8/+sXCgHW2YwaX
kTmRxmC/Y3HZkXmfiCpwiyqL2xcBiLIqhm9g0LP+Q6msySqjNJYkt0LIiAGI
32MiDtmZLp/sPci/m2WfTyjImhVZIbnsvpHur4r3i2yz0AMc8QHc9BaX6Uxg
qBQwYFaU536zK/5MLA8SAcwgAHkcWxfxYfbbI6INA1klK2TvEDruoNeVt+ww
AhX2w35z1BYfMg726B1K8NRfFgG3ki+obe1AYATpyCcd05lxK18GNUcz21Fd
vZEQQEtiqpB6BU3PbN9RCJfSb4lvZYvJkWR3vq0DBk3074jydFyOLZZ9KuB2
1c94hhu71TzeNfPwQnTZfuNbTBgkNx+dGgLqlLxSFoklE4NqX58CaaSDayQj
i4bFsjWHRTx9Uxm0P5o63Mm3sJ65NPtwKdA4hRjh69VmV6V2vINqHpcWQBCx
b2Ukl7stA4xQqdXaTwlNZVCcEAgTOdvzrTotRzo1YceT+O+wv1ixafaXu2+2
gN47H2ANV1mWDBav5Ocj6r5KV8fAKmFoY71R5+wkyyP6j+ljbzL7oUnjMAJf
uXXe5NlxX8JvDPCi9V1Uff+yeQLwPhSDB0vsrPJZOHKZ8K5vHCIeyJIsAoaj
EpMnzfd4HkWTjMgYUIbEn1ZV7UbfTNlel2OPH1dkpBDGKQE/jse9/515wp2m
W5mrT72vkH5WIGBuS7E+ihtP5zVgUSihyRib4BADKeVgL3t3w79/MXZugiQ4
tsHSRr1BPWY6cXPU0CM0JLr2elGlWnVqSu0qdX1D4J8T68QINWAEk1v3cw/e
mWmekVRg0NxAQVLzFOzDw47YJ3nUIH5jySQxTFjD0SPnt+EraNO6uJOSBLJU
wcPE5cxgTSW04plUsKlcHqkDZBiMYwLCod0VDACbdwHxJPi9C7WrauyTVSvt
rqwVmwqpTjH6KHgclojW8VtiJ3YltSPk5cGKhin2rIASqQ9v/xMm+C2Eq0HU
mXAlZjaXpvJX3XrRhjIUfIjGfdjcujFCcyaQqUTklcWwBIsQa7Gavu+prwSo
YzSrdgD6zmVcrXHUaRg9smp45l+qGoCH71/5KBgn9U4QcSgBrP2yKRPbwrNR
4trgOC8kZ8AhVYgU1dLphdBIzwQJwufPzpp5Hd3YYA1G9WvdKbF9f6cuXKR5
pJx15DVsYDmNW8o+SYUpWtCogpg9QekGB5DpwHFLAwJ7FLH1U+9NF6/iLu+c
Rz8Tq5q0DrCu7blRt67Z5KS5FFPSoUoBXpZDmHd5JN12DecJMikRcLOgIWYw
D0BSzBScmVzjo37AvMXW/TSg9gRuWgKcvONDBqkdOtKzC3zsrzo62DvzDf+b
vlui7PqEsiSrVcBcn+BV+a0eYBFO3wFaLHvV8CgkwPnD7H1QmGbiD4DJ37sJ
iRQhQ7JOLXgZZmohQbDfXrNu5tVuD0JpDmMY09payb07c4FiIuVNvbqOS19Y
u2DJlW5GqfQMiapZEi6nYq/hwdzRs2EyFGANpotfdO0FB/s6nxbdirW//Lle
LTXmQpnfulM3PKXBVOJPf+YT7PK2SKIC/esq+mdZO3uyYY3UwDMK5Sqs2xDX
zOsPuKXNcmPGHlvuSU5AxkdwwuqSTJHLsapiHAlZb/cy0T9xjJMyLTYiuDM0
nvBb5vW+SwRRdd2dZUBf6ZKw2nwWkTrjSknqzCbo1sNrG5SGS35vh7x4WcMG
hz4ig9F0XdRRgOg2W6La8Hkn5ZIR6Kvk8he/wLtlE+eqhZuhPhNLqMJhB1DP
ZhDxkE4D23W1T+1n9WofnHl5DJadwxHH9xtTY99vfVxd6ulZq2kM4aaYheqP
DDnQobnqdzNMrxoCB+n+LZ03Bxeq6xfR3IIHkKazqOISVwKZu2a4GaGuncYD
43rMenzIwyVfwfiaCU0Pv7tUUyVzaJkSycZFpqC/O+lD+9QRMh2B+Cqj45C7
GrHmPUc9PJZT6AAfRqy7T2aGs6Ya/YqQqn6iK4rxH5aynpIuaCNRwpKNTXWK
2c62iaNFlHVJiwmi8CeM3C+qqBmKV2+eA/yNBNRi7AYDgFfe6RpvX8mXraeL
lIWwyb3FE2scraX1wNrx5iOtUhA8gmxZAjcQcfo/OLvbn5sXvH5hrhlZlscT
OxVTnQ1zzKDX+9p84WGKt28tqcZamSOWsD1uUx7mrWBjI1F5d749vlFZvhv7
dOrkSZWJEJWyeuZX6kR/gbFBds17Sr38kjXJwkcqVVPdwKFOdgToSC8rqMV6
BZpinhTVmhXDRr2mfNORscoaoegiwlbQRdrYGr0t43GJ598lPivMs1L/B/MF
ASHyi/Y8h29oqfjJEjcUJR48ks+LCighImA2WWMhN+OoJECx8VvkrR+Q0P6C
6KaAaQHOTCpOY72Q1KFBB+pqyFvr7HC12ftLupIHPIKzJnj4TCAIYUC95VeF
FI4ZL0EeY7Dp+yIbDyGA76E8SJTR102uL5hous/hfFjqWBYYiiTnoFOEahFl
zRV+U6Owp7CmiFEtQmIznKCdSIOs+gXwfOcZTvZlWH6sQSNRjGL+FxoxZS1a
kySS4hVx+A5K1lMr7EAQCxC6fvBb9ngl94S9V5kCvEIqJaXmWNBU0bg1tpDT
8dUpbzfolBLDT8Nxn2mJWn76jZQ+eI3UNrx1VmMGJW+wO/H7zeM7LGHPur0d
3BZsIHDSS9xXIcS4EQq03sscEkdodcpCp4HXN/WhiAX/SkJkM5VuYL+BQEzm
lsOuaZGDlW5QPb3xwbYCIIbO4BtirAIyOfoeDUcHMhWFTdUyjRCkcVgg5X7P
tZy2+0qjwlFkzcezNdXFibaR29BaFdi+m7JFQovTaARZw4shh2f9mjPYDj68
ahpdWsEKc0zcxO8frp2CEY69NAkgCKTPZ9kk2HglUsrk3X9GA/GIftNpSy3q
h4bR+grxagQWsy02jqT9nYev75VQGJo6YMGxOSL0JchSbnlsHSQQfPxABbz0
Ov4JPY7HQV3do5X48PqyUa0NX1bXR/iVpF/c7BX4idKpkGfG3oFyK5A3jGO+
G2QMyZMU4JtYxjXQ2NnIB80E4qPWTUKVIf9Ar69SW6BK5+SVORxzUxz7zIY2
Nofh3WZmLwP61xFnienjzgE62RSgrt3vg7krbkPljfz8YsI4iNChaT8FMiTh
6FuOQ5omw0d8Od0LLLg9OsE5X/N0m/3oNm9s7n/fggLNZbLesKiJ1hxq1g2s
0sLxclUIAk+6cDxVlsgDmyq/0h3IiAMRFSMdxQPASLhkD+suzUfwqQzmR9mX
iul4v0JvFhqNO1X75h0Z8b2gF6LCTtNmMiTT+kGfkc4EKlDjXwxIDc76OfF1
Oub7uSssf3ALDZfAJ9EpenerI5vaNBBJyM2KeTktm2qsTC0fM1SkMytCz7Vh
A1ONZt0imv9qZ/j0fujvTVWLoN+FQb/EY4UxmBS/bhKzjBQ4WaG0XMkhzP7M
fkXI2q6l0zmhl/r8/fo3Ku9pdA/uDnmjS7/WLF5sxUxORzjloWfjYtFq4mwM
TQKxXFjiICYRaR/9zhIjxSjYPPRPubvwT7SL/x1zogRJsr3cu9WMPI0IgOYO
sTR6nVQp/15D6Q3sa+io/Y28vzxKUNwcmlzTkn5cdo4o59p7zzX7EmaCqEwR
S9tU5jgLbsjcnGh+QFmD8BqQ16aXuWpmUJAyTTeoRvLx5LqnyFxc0SWgCoaU
LCLiBOazMgSJozw+IgXxePqsx1/AIlDLUjhgLHtATn51Nled5+Xd6Jp2pMZ+
8OcobWMiIlCbyBgPi5qk+Lapeuyelr941Ghz2Q6h0bPIhlL7BUZ9As7jJCEe
7Tjw6bH5L60m/Dt0GJ6BAhJ9Obt7sZIs3LZmQtuas3gvk4sBjqv20nK0zVon
ZUCuoguj4HopihB/gM8IHw1ThiG5i79cgdYAGA6FmAfXfzp0Rtq72vydqyLY
CG1pyqmmxSBup8u3KUfxi9PbGzqcZks/GqeI8KgOi0TyITdOyTbxr23cg/59
ASZavM4lxZyAKirB4Et6Uj7MoT3GL6VNNJ5WQyjgBscU/TfXOJZl0apQ2CVo
f3hUsCr+Nq6JA1UDBI4kVmvn8aVBb7++EhX5QtfogpQX+nCA8B/xcS7eDhjb
gY22N4rTw2vYw2ut2IH1tzTjZFG7Z2aeUCMTqIR5WZirdolcPeHQVtJSFF93
wO2561RjEiwnkimbGE0th830+m8BDSI449/6FRe0dMSRWYXVjttMm0xK5ptN
7LncK/V67cW/TjMIRf8lirGx3cbRW3FbUxBeD+eRmuJIX2RNfg5fwfPWp5Eo
NbDfNSEjmyOmgKaLJ/FBzYVKq7Y7gnah6jZslQb0dlo0rFqL1yRoX5n8xspi
hBwD8Yi3KA4NegMb9sJZwKxQ1tsv3c5+Ow97EkltDSFDbiYYzW7zQJb12ANd
yK2PstmIk3nKuDVTYMUg/ArpxcpxhoLM73egjM0CgkWh9X5WZaPvxishNhmQ
tIOzKjBMUAhtPWdSrAZHPIm7cRTBN+4f/IHA0zB/TGQVjneInTMWOW2Z5cSZ
zGHFUHaBlAPca9x5wtcGNDKRRgvLtg2Tdj+iABY/nn8ov/adCTH4rzGvWNcX
r4WX2vflpGDTYNFIqWaag0QVD/N+GS+Uiffqs7vVQ1elsQlfSTT7cmklzkE1
WuKsD/3fQ4orY7o9zG5uigbK+vXh1FGTp9uizj42ZJKSjL6yk6wtSkOsY8JJ
kWl804kl+WjCVJ4RdgT70lg4adWQabivEL16dd7T52W/MysGyZKkd31kNpZG
tHfobJwd+RDb0tTXut96nJu8sW9FkW7IQ4aEuAqsW44pAxGj43/Etaqa1LD8
ZaJrueqdeTGiI39GxcziLwgrgsZ3MGly2mrxnRqJravMN7+ijbOJi+q0RUXd
NhEDW77hWaFE1VJrA/0zkKVmoQxJTxvrb+uP8S+mKgzKkUV+kz9fdzihTvAZ
LmjiT8PGChb1JG63Z8O8xUGD1o6qvzUVquzpRlTzcy3/qsXsoe3bp2B4pkR9
C1j5F2/S9CI+L44VuFR+qpbhM3Mg/jzd1gDuhjhrVSo53M0usleaNRobqaL0
gcVK0Q+hdvKaNFvuqKkEhv0qZeh44FSV7GFjysBleDs2tFmfBwmbOtWqoWWV
vQkKtCBWV+r2U3IzvgQOI/h++TqR7GTzsDlzkeNVvWxKcY3d9oBltdPp5JgL
g6ZyEjiEAHq/l4FL0dj3wZW8rwvZLeWotkF7IsOdS+Gdi4dvLWFAqurenjDf
vx4kdgD/ikcljGIRAqFKrYSO3J4jm71Z/OCIc1yHE3etBVXEcUgpn23tXwTT
7OVEsnRZbrJVH30T0cW/rULxwgA2Wirv1meBTSBTTQIYSk14H9BvrsFuBrAK
LBvKhOliIgfOhDz4VOS+sJV/P08b35pxvYKFNRiwbHtD8DfOYdC/aDNitFRT
j/5vON0DRZIiRUc5ndtmED0ViZmbjk6pHip1b78DQ2CsZxU3mX93gdcUx7wI
YPEYrp4pHUkgTtiAKhPJe15ype+NcUv96/DxLqYvu2JDMrCcDNlBLNRO0lYs
Kz0HyZm7HVBocM7BgqboaqnwR6ID1ASnXjErAXB5I499vvzMzm8h4MgGg/3/
tZ3ljvLGvXjgmEtmqgWoQ1nikkYRM9P3y+5W/V85BrdpOY5Q+NzjfSQP4w4y
XIkFFPd9m2qO4FOBnzF3mDAla8UTERGgmU5dnQqFJRXHyMiRavAo/t+yh4Wk
rIKG0DAnJKzpZFkjdDcBbzCj2kYmeJWvAAaofAxr+KmEXb2jP3rJ6Xiv4Iuh
jsjSkjMvUSe4SspTGP0v/RBYyRn6mDUv970WxDikQPyVc+MvFjPR4R5wTx4g
AYeJtkb2RlSf6HSU2ur2c8ObquQA9DPvO969rTZVuKAev/yJJsRq2eehe3og
i0q7jRAFK4AQnTmuDX9rB48GmxQhSEFPrWTrcncN5Z7cdBVtI3zJd+dE7A55
DD7MZLy3YfOaqoQSFCc+3pVF9Bqopz/WOUsDZ7JGvEp6JWmkVDLT9BNG70hr
jfmQDpTotOElb7tGGQd1tstTd4UA6EE8V/WjGErq/2L3LPVgHEDVgjJlTfsp
3s/K2Ku/yjiprcADy9308YcAKm/0IdA4OrHitU5aKWornlv2SK3OTWnqx3m0
/FRwFoOM7XDaH14PcqXxSMq1wW35FO5bnJJKE8p7U8Xcgx9g2FBxT1NlPSyT
gMSGBCEp3iI1skmAHD25fCHWSXQ5N3X5ER07mjcRJJCcPJF/3SdcHQQ+wYxs
bAHd9tsEzz6xdqt4/HKXb5mi1L48SuZZYX278GfSf0w0e76tpjo3N7zAy6Dw
7IsBD+STNr8VYBYYqzbGV5tfYRh/iJ+uwQINaqe8WfUsgs1jOrpXmLACnDaU
TSffNJcQHaSLcCViKxtNZSn+S9v6aX49HsA1hzH2frlc88neZ9kUZyzViXYf
QA9Rk06Kwyd2Wbq5uAUx1HDIJigUUT68Ip4gukp9GPjLDz0MSD1JgV7vBqUn
XdBuRo04n34yat9sQiiDHeiXfm1Icrf41mRXljE0tgLMWyGaX/QmMHchWl2Z
mrr09OFp7y5hkWzlwzF2jS4tF/4U3I9pC2Z0nnevQNpJAof5/aNirCa8V4Wo
laE9OinzrFJpGeQ+0RXjR+5qmmjVzme5WVZOfpktLL74tQIk8lj4taQ2sb5e
xQFz+EY6TWEqYyjzkYq4e8vAhlrXn1oOennqgANdR7wjpCpLAGtGLI2F+a/m
sO1MUEuY8jfE3ZEmV+pSiurvVkj/IzDwSjrRXSqpwejhOhgJAXgSwNYFQL3l
avN//hwuLIlt0uJxhEGCnAv3aKwh26mK1D9zr4RuOoc4iIVfhMyj8JOngvWQ
KaBtfn5gBYfku5shxohMMEeSI9dkG8KDZKjWA72EwU+DP0WWfByFPEuPoX+s
PcvYnDp9+AzbM8+9TCwLFJmg0REJyMpyp7gvBWu7pJZ4fiomJPxUdMa9uXe8
xm9baA8/x5tzZoctVfzVbebKW9vRWVieDINbEBUE6wC7CEkR7NTQNbotV+tb
eGsVrRs3twlWHNhMl0BbO05nFWn62T6a4knFWFOzI8eos7r5nza7fruArs59
Rfv2NQD1a+iwgDr/4CVyku9m7lHFGu6GvzDNP1el2fQ9jo7IfH97GtLKKUQ1
XJXPkG+HNEdX316XU8ImBZ2oxPNatXhYoWoXFAt/X2AsEc2Kh+M7NtQB3gwO
g2cstOwKtWXccxmBjklCFQLjYkIvpBRKN54uYc4FEv1c6wWv1PwsMMH/tT08
Y6LuU1pRyOUxz1nTaS1dF8JVMt1meOqY4Zo5yfphIedJvrZbVrCliOd3savC
K2IQ3KBFqmI/8AM3SPhdVvfphDy+AmhnFmpoaoClPh8ezesjg5EFxD0Uxm5o
8IZUwapFKUfTWn1Pv1LbtKovzbvaocbWIzy7/BLLqZJbhlNo2LSSZWgUT0C0
iKQHSs6h4FU3eZYwwWAn5wWhCjYDQh4VUIEmHv27LrYjLCX/7g6C8HmwXF3I
Zl0YJMqJqNWMs7KXd2RihiRtb4ML3YEIFoH3RMMHl+W0WmwiSa4UzY4OZ2Ym
ebcW51pXsjZba2EZ+LYSZKgmkSMa0qrEn1L5HZ5rKwMJHYcie3mjP4ihzYme
BbqXXRFDPZInzg3LpDvelS+XILk3EvgFiUq803Ewtr1EaIXJ3PXh9SSzIVgH
Xzp4FrLZHpFpIvmyCfUpw6UIAG6ioCFky5W9aVv3IKmOMg31vvWK8Od2f4I9
C02tnB5faIVGINo1CzXT5Y67B5DtaCY09AkmbudRUje/WWPXtXC7VDZdLYZl
/2C5G7d4bZfyGgyLovr5Nk320/8nxvuLFYjk/J8Mt9OtV5PVWjwtBfWEkRg4
4Pve33g8nMVfBjxqqsQ01M6w8GT0zz1LATS00kP9MdL0Juh2Jnc7FZIjgwpr
eAiUho2C6ZjtbIIg7JLbJKNzfdqxcL+vlUUlRwWSSbxvRo1syNi3vBtM1hEh
QSt/fs3LsZ4kb2tIyf3XwcffTbXoWwhx5DzFEA1TuT4eDrfh2n3GyBhnkBg8
hEc7SlQvoLGlj8v5y2RYwCvpOwQw4N84d97EOwXgyJ121ErbdykDtY2r+Hze
t+/5+V8xDnKSMPu0h5NjxbfBuA6v9/rEVMkaJdG4rRHWBVROHLhBKQXkZd5o
r554nWqgoXSMlqBXryACYAM5TvOS2qkI37qaC3cX+cTcq/dU73A9Gxwh1byW
lVtkcVW+aPF5QeH8ZUQxkcrG4bFS3c5VCQdbdS79+zewEMUnAc9GWVdGIEib
Ls43CU5OElgF9mqp30hZz2t9GWWoURzZb0ZS9lpE+yRQtJ8aKLxJrYb0V4AI
m6wPHj8KSuZ+xjeJxUOP2iEuBno4WmWzg9FP7okPLmLFrHA3/AGeCR6ZPnNT
v/uNsbwbQEXMcQb5jPa6JZYb1kCuaKzT14SBjH/YDfklWBUYjymZBPgnv9Vg
kAkIRieb1w8loP7DHnOwjuZ0NZhGbogg8Qm8wiYxFjhO13K3dqM1nwFd235B
6J3SEXbqalPICuZ71CqHCF6lg/C1AkpZON9zV29Fswtc+3b4j2xzNY+I30rc
s36/EVBtc/lUhx4kqftNvJAlWMXGstPYtdu/QGIThGxAF/pGY3YaNY5Aqska
yGQywLv+QTgkq4Cd2hBG27FdZeGQ/F8onsh3JnvYZn6BiF9Ve/uexe9PErt0
0yezmnxAkYqTYGZjSImDC86JUsNTzJgivyz46k7xDs8xJtozseIbHo27jRxP
mBqzfinfnYlwe+/meoErUnMoWxOEXqB56XYHBR0PGymp7qHNkl/8eY9XWt5z
tAxyiJ76KXRh4K/7I4pEa2dfE2su6utrwa+Ht1LKDApD+BJ0z1D/Zd8OOSHw
lwUMT9HaX6/wIj7EwsrOEFSoe32FJYUZzW6kljmN5Z+bQvr/RMGqjLnM2dyg
DMLt/r+dK+LO5SYGtD0KOqOKDvSGripba4WiaT0wtHht8EameumNNbbCz191
qhdUXW2KwFkrL2xxP3T8PZoKhtSqUwMu/DUBu0FW2ftZ093W875HYWnj5NU5
Tk5wYtERso+aa0iXy1AxkX2KQ2Lm1yvDIpFtQ29FHlRs4lkB8p2B0Ox8sEF4
wxuHIAeoKRmCe43Ug7SK94tJ3l46USiYcuzvfbSBMmDysJBj2kcz/PWYtUvw
h0tuJBa7ZTR9fZ/im2Jw+90Qq8JCrI5F3L0/EgJsGtWSfGr6M8vnjphQ77cx
6RblE9UmMcXcDHyIcn7/JKNb+nNwn+vbwTH4dA+IVPC7WDKc4tkcFTSyv1yo
kBErF9Mo4tAO3LvsOrukaN9yBSI8BGm+MreG3EgNGECQyypZ2gNWB6F7dCNm
yk4SGZ5Prlqm4IHIS9fcv1C8cBRfeOh6AlheN4THiBBh6BqcCdqetggqlE4i
1FelUgxicgmC8q6xP/JI8g1YVY2HpgVDsP+2Gkt1nI4PDE25wUzr7e/1OT5W
8SsB1ErgGKk/jrMbBrx9TBliaCu3Pfu9jmqI4cFeBWUK2JEZBZePnb4gkoOk
9uhjyGqjR6QcqJ3dSpCcAR4ygAQNWoABVlPZLzEJBhEYsNmMWm+bAUD2yn/M
DUr1wMWEnl3WtQdMnmGDEcvH8/vMIHT42NXOM8ugSKPTFUBO7JJGBFsqT908
YppYbOYnRPY1zDJXInwA6R5jRj91JYGKRfBLQX6iRMk5uUWOkTXNaO2QDlkz
+xABu6ApFAHh3QDzBUmgIPvgAYKYc9ItXoIjRL0zBBwtobP0HEwOvXCAba8x
ZPXziEGyLU8ATqajXNrbWdwyi8t+cJMcBxzB6pBuXVJEcEJdhsVSyGTpram0
ZgcGOX1UP9S1qqwBx81XV/QbekTB7STWzdTHTshsNkKV7UnTtbKsnK1Qsc5r
+3I+sjDKlKm5ZN8VLtcre4HpH9AlTvcy77PPYuKNLU4UWGihEJ70XEe/ri2F
+2pZcfkP9/0ewfAjQMMtHyBn0GrSaGbNPbiK3vkF5N/U4er0BYt5xXVQWThK
sKQeLr7vdTgKN3eON6Hfk6y/Nnp2vvtftJbtphSW7CkdYDZ1BDx+OAS1HWvE
9l3pI7i3gi+Oo8VnpmzJVk3klVARIIeQdBsQBj9VCqDUuPNtP6ZFP64pxwwU
QfF4UiNXSYPg9fR2/7s0ykX24XF3dwOsjkGcPabVA/+iv3Jj0a9aj/wKeg3t
QtNXZvPg9QNHDQ+DCvMgUXWLceOKA49srhVJlh1ysGCwkUYNSCpNYWKdbRA7
4XgITnOfURC+SmeabAReIkPKDrnVskQlqbUKDEEDWg2qfnYPVqbgvRsvIUn2
C/7iYAF8aZAcCWqCAfPD1/iKgQl8KeIQQ8Bs9ilzamHQKE4zyeKtF4Ee3LOj
UHY8cn3fIIK1XlEO09xCLgDnUIvNgiGzDk35OEkPdSLYCr3RjZOmC53P5N5i
i+Y89oLhvJxH5O4DSEDgsHV4zToU3R7j80dIGdBFlZWODEaAZif5ffqli877
yzREL/ntxejIhJouLlwJrbQTLO8G3DnNe4Pg+/5eAiywLZ3D2gvVTqklWSl5
HJRW47Ke1Zh4v/brXATNsI/4t/FxXBHUIdMUM6hYtVHvF+GeXPd6HD0DUQzh
vzHiffTjCm9MRF9PLXcQhE2VpeYOuudF6K72ZMrnzq6qny2HVM5a5PHBN9NS
+wTjyn2NPfi/fe65cRBNNWfTWcrHapgRDirP/FCTUitaylnUGPm0QkIH600k
dWINAHkE7mpP7u4KLtjLJIZn/+jrJJpV9N+YI1X2/E1JtPZMvZo5Oj7Dk9ZI
Irc6PmCJkuSrwHpJw2Tv5G5o0HLF0HRWKQgdY8fnEJzclqaHblTpmX3eR3oX
nOfZLkJkRg12rY55yWgkF8jymmg2A2vUiI8Aou4KY7hYoc99OO+cxuJ876VU
OrJ3trvvIhwfHQcbWNJXHhq4vbW1ALwEJ6MHV6c7H/Imjn7UnedgbqNcJ61K
WDO1y+nUGkbnYXjNkoxhTizM5GL/uDZyA+em6aEHRcgzVrNdh75aXbKKqV02
y6n0pNd96ewWttJAFgmyguuXQ7t97Dbedd77I7d9lidiVbVCnWyOi6xzWFkN
fNycTAdVUzjjFut1+HX1rId96CLYCWk7S44XEiKPDKnEyvRm4mVxDGYlba2k
AUZWIubWx7t8BsTT/pVMseWrMb8r0Ya175foMwm6LISZDz5fKfNouYeoiv7c
uhAIhQ+MI958GaK9HuwY/BlangJcdqvpRbW4K2QGk8hcTB0pfAR5QQEKkNjd
WSIkjcZ7/btZP9p6Z4ng3vlgd4alF2Uw3pDQz1NH7/nUHoqOiksAcJkvMUNu
OicKthiLbJbwjRveXF42CS4F3U23jv5jNtRb17CcQiy+wiF790MxalV3utED
vCi6wiJ4MgYf2g5cHWeCWtp6HgyjNIsdkzr1na2dZ7YER8AIYrrj+GL4cL97
zx1XvnDx+Qszx/V96WtOnVvOFuL90hMMUdxD89Q2v8BklGTfYJL4NiOD5hJ0
96hyt4q0xv3lPR+nXMxcmnfecG8mA2cydA96XORlnBoS/4L16bN+4HGGAXVn
7NvzNvpaClvjGh4zjn5B3/IRoZVuBe0VjVu7bfgOZtoojT83jXvJrkM4jeC/
nYdKZ97fsl4qhoWd2v6Rt8Spe98V8chy7uMABDm5NQOAY5l1XS8EDpxy6FMZ
3RXYowHE5r1f1X6ohwhOis8rsWV25AVzvqe+E+Kd/F9rKQ27zndgOrYArajv
h4QhsH+0Cu67diVPZdCodKd2F0GSKY74Pv5w8bf9+HyuMWc9i1qduwf0xJfp
/3w/nEEXRLpSdtK5Geg7wLKETt72RC0TZD9R4Xyd8XHz+UpJh2IKI9tUEAvy
Odfwr04+gX62faXIvH4c+wy4/3nQXX8mCaA+er1RVTjMTAGeRW9/ewqrYayX
BtUaE2dMHj0xTPoZyJtUjbMwBzBJI97yexk2H9vNHATs+tsL13q88DmM6gB+
85yTG4ze+7548PtobkDO4yGUulmki1n883fl0g2IwPAiVZXZgrElM1nM9MtJ
hbxkyEaztTk2bPDn3lbJdNpKsvp4raHunZDuYGWGTtEOxBCZnxw2vo74Wctg
/5OEx3FTjJVOpbJCnf6cn4THOy3BkK1S5HFUeDFRUtlPEU89/m4ND1K4tj5o
+jSdHtX7X5/oFmKxkBuOiwq2+F9/mYVtksWG5oqkao9NhL4XtEaNj5AxlEMl
1pvkb6+CEuYd18UWPbMGfIRMTxB+kzm+kbEUzt8jCSKwTZD9Dm6xixY7iuq0
Ev95CYyGXQgjbsVx+5jT3ISrEKaA1neF0u019P6YuQBfRX1L5iiOQc5/dkBi
OLrqLtzLKlD2DXqkTbh3cDiDMgSc1LyvEvusAwbEUkT4h6Lg0Ed1n7tao3fp
n6DXK6lSdhNVF7YInj6WSu2vc/eIK/bdZtFQR3CXvkUm0pSojf0i2CrtmaG8
gxFfvanK7O9CmLhX51quR5zXvhuOLfds0ESIs2eedAhPDJ3hKll3oepfH6Yz
ouLm2aLQcE67PPJq/48kTipEtonw3Dg8JzerMR12SUoQzK/xLtKOJE+08oom
lthQTodZ+2OZ+7eWnNSCFGeNmgiZgK7Q7EPma23v3sQQZbQJM61lIl8Vof/H
tQc4ByS5a+H8XoP25bpMGXOmmVG9RSMuWV5UT9R/GOcvBDsBVlDJReZxjnxS
uA9407xo9hZMGr4FP1uEGV2vdwS96YayCaRHPIg8g0uGsln7DQwWiaZzYCN6
81L1FKtm+zjeQXU2V4UddfanVQ1QomfQZ1TxXEMDUnFxEPX/P4KXrJztoL68
9MjX5MJFwQesEsOQkjxxTUR2D6kaFHHhhapGYZvH5vad0g6TG40G5XaFEt+b
n0ffuISJ2RqxEJ5s9RXoJ9+LyC6W/BXhP4FPxMrPo9VEOSUpOhUioTWZXvPz
3LXuJ/IYJc2yy+PUCWxPJuPHoOD11WyOApvLovsRJ3qX+8ZQ+2ffwCwWHlH8
d3Vx0dI2AEKabMHjrIFwummbT0rKixJCd6+eS35sXVSE9SC83lKd4Z455ubp
O0x60lr6Dayw22DndpM6gVrTj/fjKKmgh8ygkuuBNU4I8nfKesLpYoIFav68
hyqf9p9IAKwrW1YeRHw0GJusiyRj3RjbzPI03Jmyv2Tm1JWGTtI9XDDcuaY6
+3hf6SSXNancwuZd+yeieSKLNeES6kreXQMpSN5L1v+UFvLdxmfse1uxt6ph
g+OqXKRHgbnQ7KSfrTSaZpNGnfvg+QynIFWoc6++OA8hLBb+xdk9mSoaS1nO
w6EXpPuFarl10a9t0JWDyc5rQ13E846dyfSUuvw9b/IOEz1XVztlFpaCnaBh
9pO7wBb7YkkG5izfo42Q5xsVy/HSO4QFozFO78K/E3pFnBHlIFs10guYYhr6
u8h5Lz373oKtH+7/7VAS7bQkJQECDKIx7+nsfhmi9d/jjc2e2rF/jAYHsDvZ
8SvA/xzokLctU/olkT/BVjqPLQcDixitNKBtHKPap1+/93m9DsUo+k2GggDF
2RyCuGD7sZR3L4FnX5EyJEfr5VQkvV8dSNNEbxaXU4fyy23iXfLzwsnjJUIb
LIV4DtAAcRSXQae8EHOpLB3SUgl8rH+zpyydSZ1omd0WrgaSNFWsFid44j/K
UrYaOO0/S1dlMNCF9FkDiME+7LK2o0SSKLimnJLxrsAz+42q1nwQa1Rk44iU
78IZ7zKfBr7HQgi7rkdqeJgqEgIGb8hYMEJCP2aZjIDvazSJiWqw4LYCdl3a
W9na/DgDV2+hmnyl8oWWA5750lkAv2wraMvQAxRdC5njm0L5usukqfW/KR8V
EWM7ym43IT5o5DmDfSLybL6nh7Z7ASFKCG+hXbKElfYuia/+35P0kyS4VR8N
w0+pt/K0p7oEkIYQzi/tU9LKEql5HHm7tsyXNVHOD02iEH12T69td7zz3ysz
cOt6pIjkFBGkJDKVfkIQJelA7JXvLofpd8X8NCSYnix2JvWY/BrZeQqEnFUP
eli6YzNshaRXo+G+3cqP9VmbYtdIUr3vHOFVpc8ZzdcrHIbwbX70UsiZb0+u
3n2c9wlkhsDsUGMjBzWQCbCIzlc1cVl0aDYj0Og3lX8jNGHzb1x0z/01n7xo
ZrYOdokTopVrtk3HMaRyIsIFivYPUuRbzuif1SCniIpeRuU24nWnjmuWsKBg
1Fmyz1vz413GJMEFljVGNlOZDcSUyG3NEgKpIF7yi5/CKN0lsETeyxwKw10n
z3ixhDwWjytc3FuXov25s5WLA1oIHaTkouQdNYPUGszD9t1Rhp4zQxuLE7e6
+VfidSFoB/Ex4CbyDqoRU6+4tcarbrX4rWJgHZ/dNfw2hcclY6xXU/NWZ+NO
rm0Y1iwIbEp6YFAX4zhnTtVlSpJw6c9Ah9sqI67dJXAK0ezC3p2DvVxh3XWD
JJbnl+nYYZwg06ALyANkp4UaPuZ86b4ZK1IQJfoedKAoNrjvCc8bltyQ6hKA
7W1oPCm3uXFmFddOOZFKaoX3PE/TVpD/0oWU/vcOzBYzbJNtiwN1Ligr+Uv6
rbMRVZz3Ylly6DmWLlr4XIWk6VtSIVdQM0WDEyj4QsDH7v57GB7/ZEuvEJYs
W/Bey2abqvQwVmqu7XM6NnHv8288AP5rUk+l0+oIX6gIq0Fj/UTt4sAHi/AP
yi2W8Zwcga9aWZA8mLfC9/S+a+zw2k7CvZyPbuKJNr6LPP+Kq7/07/+3Gagc
JHEKfyaWwFK92SZSTlMycnK6hnkMNtd/eXs9efNbKdsYdMS2MmuG2ObNnjKe
7KyhWQZDmSEuyDKdTHuYUQycUOrcSEO10uHQZHZpeRpSokI/xEkEHibVz6kc
QftXCqse4seU5SvtalfNlKx5eqOnxrESWIzzgKhrrkqJ7A7qkpsvxrfy0Vp/
FtDVctZ4xZbzvoBk2jRbVnch7LQm34oIdS0mGrXtlSJCORqlPKOUUUHi9/v8
+5rZj5Q0hkuSB8v8x1KHHEPtF0CJ9mtM/4N6JWlSOgCsgL/JI4n7WHqZBSx5
yhGKFQeZ4cUVPWn/0nXqguixmDYywd6KYrh6c2IH88qFmaYOnEb1apqXoBhu
IqztW6c+SAOJoCWH+hfmYuIKf03yAmi3QVYJ5hYFnnFxsBmJ2Bly1kPcW7Yw
SYej6DlK6UqNTvauA4Q9lA1Q9EMxhC69Vb4PUER5ZUS8bnfTgrQmJA8f6FH5
9MDRYLuLsi2cUQWS/1SIiguv52pSq8G+qGu2GVvWJWxTcvWQF+OJWsOJiBBt
pe2eyvogKI72cRBnlw505h7AaQg8eZdsVxx6wgED8e/Ob4t/f0jt9vefy0gu
IwUwnhNjpUxq6dTKGFL8cAILhJw47Vs+B/9k9Gu/iML6Z79O1PTtJRDNOTAB
CreGri0o+/ZaOqqhQqhPs9t3S7SXmFYYLwcITjqw9a4T3BD9il1+Zax+HdZe
AQV6lJS3O3iXdGCU0RUB9kMVnfkz7GUyXE8xugML+rlsRMNqOlbq62mclLeH
uIYlU1rWkZaTNGYL74cGU43bQgKFC3dgmD8XBtzkupydcW1js6tGHrHjfiUL
+pbTsLI61YA7yy/pfDzzciSRyh4wuh3Kc6oQItQ33VtHcDvg6C9kWTDKcLHk
RPwnI6XYd6kgIKeSsRCkn+Nhyuz5GixojQp5skfrShMSyXb+q4uk2OKtGCuy
pZnsT6sn5ozjhSvrFsLEarzoEX3ujxF3cHoxPh7oOFLzwZAv86rIxfr0wGQU
yBBczaCGJxqRx4PcXHw1jPtQx3cPKVn1ELZp8zDNkciGb33hA/1olrHcvkF5
Y0nwMwM3eAos263tXqJfteAoa3tbzYfmIu41J27PFvh4+eYFu2WZW0HTWsdy
8hNtTo9dFHOiWxh4OPL0cGjrg02HnfCuXFkA3sVaueKdiI0DpajuQ/K4MdfU
HsAQIcy0o5tD9epZgbz5DN2fnkd6jr3+Ui6sgsSckvwuFcO/uBsjr9ZFviFu
Y78XUC0vwJvkeMCBUvd/VHjy+Jao3C6kVspfsf33UAZfNie96k3vcTwRffpM
loa/c/QEQ7gJJqq47D9BlGg4dc4ARNMF5W/0ou3KgbHLn2lEKylCIPd5PEO9
mnXIZYRaksV0LU8qpusMDD4l7BxpP5JDUVxETIJGhFP2SUMBhMwzwT+S5Fgs
DeS4p/mHxxTcfuwr3ldb9Y2qsCQulyb7Qh/qkvfpj01cKJYPdDWdOlpTATTV
eGGkirqFy9p6w6DJyD4Q+PNyqPDcAuIiYqDjeS1OkTGNQokw0hkYqLvpLz3L
ZkqsuYq2I4PD0HDPFEzggRrwPQhYVUUaIYSw9fLx9qLcHMkKj2RpY8DVgl63
8e/yD5W/u5NE2syP5QDGemQQ6LVbRNUu4f43z25mVed29iBtUZq58Qk2QG9+
RHWGl3qAicqA204XiL2+kSsSdtnguO5OgnS3MJ4raEiALMG9I5BMswMpwZwT
6oIxE3cf3A92KWGvw9b9yjeHwnBNZKeOQlw6909HxX2inPgTyq/mw3444dJ+
0plYxCZ/cW/dXBCOdH89oQ8tPWTn/vu3q6AZjtisl/qM6d3AelTV6oLid+N1
PxiPq3AQWJi9tvdMWUyYhnAqySWJOR1BcSOIDU8DZA7hWeRO628x8yHUhFlU
aeSEMD/BW/a0vPwmR+7CmqWCTENV28a/nhX2miG6IGwZaDQB1RnnOI2z4KiJ
dF+qgN/2NaLEespP43cpGEa+2MaDW9NmhxjW4znX3KP7rlzPpug/thoKtD3e
1fhSFcLwcFMYmOOYundSwUlcrubW8RJklo2pFeeSJd7CpvqN79MrV0nxeYHK
AqTaqtDRxiUaA6jvdlMqICMt4cn4RXepfKN04VEPzjhTcr3NgbNvnqOo8Kbq
gbxKNtMuIgr/y7ZBcU3GpYNmGwd1Ie1g1eq/5ddJCTBMwIX7romVGU6/4K+1
wTGjgdQ8EaXoLakACceu4JxJhN4aXSs1/C876nN24rmIgAdoiiWedaJDDnCf
Pw9FECFZnwDPsZC6nFrgny21xfPhKPDgnZq/47OP5fr/jJOsnofZKq6x8Uja
WZ1IFkYQy7dezRB/V98GcOaxUhG6TyKQ7NEcdCnc2L4apr9gLf3fXAv3BEhk
zY4IFIJ7igAnf1qK61tpH7lOc8k8YrmHhaRladFHQIIY0OCAMn7qEovvm0xv
xPj9jq3Yg01cieqXOiwBQ82WojzKD1eRGFFvlMot+GVxWGnvlGPVPjC/DQ7F
d/F+870J3IlV3tNab6iFEC28IikkdRe+Dc/qCPCk94L1X1AjgnZEYMd5Fv29
LnsIt9fmrrsUlCbJznBmV+koyFBfB6vWAK7cxc6XwXjKPvAsNNys+baK3enA
051jKB+88lhCrm9M47PgsIpg+4HoClXMT2yUlYjHMUTKwfnuh+Zq+2cnQc5f
AdYfZpP/563RADQ4xJqr9x94USM47lfRI6tpRzIyZtoA5hMalvq145MfAzMH
VOWusdgOrOj3c/dH/KtWfTYG/SLRoz7X5/ipTCZt/7aDH639P1IGcT5GrAJd
YrN+6YEmZChBPv902HaY+hXCBNMbFIdn8ClzSZLDg2JjpU+nW5F54PX2Q+ME
W6y+21hA0Nv/MdZPWGM/V1PHx6JQtfx/p4VnBTSKiWBgzBNUh2KeNVU3k9fY
vTiZVqcZPSH4jihKrzkl7kn7MxnUUmQ9CdHPd+mQ4yq56Xqmg7ANVWDc1WQR
X/OmOUhzpxn4to6M3McKXBDq6KYjqSzd7ZP1Ik9+jz0HiqlH2i8AfKhCa/S0
+Qfv7qGxuqg3OUebcdHk1x3un7YanzvMboQXtGBVlj1ObqJG3/VCUw5OXDkN
bvQQhpfRwz5gZKcHYwETEEHnTHSSmxxtAPr6hzvPFMFjUfMycqwinFZDez2d
dtUA3M4Jy6ScH0jEMyHqUhbLne5T4Cuxzjd54rdXHuVY4PbPwLB47TpLPUVF
oDrYdy4gAo/Y1rfux/a0tNmqPcTSoyju4MB44J9oaB/elvLj/L9K/+I6Np3S
YQCs3LIc+FjUs5t6KVgmcO0RmGPYUjdZb6A8d60U1kQ3O7YiBVJOIU3znP6Z
+jrmG8Q+kDNKrQB0lVCoo7fw1TLXdFh7DBv7LM5g9Ui9zmM65dA5a5JxypPr
ATB3B3vMjVdgucUhx3C70juCJ+0HzpxxD7fTZvWo3+wfQYVUtiObZjJmSdHG
9KOedWHjVnV1HhVB0EaWTl4I3wtND3JN4agFsLf4PZM/Knme8rfeXlmDyCZN
7NGgcZkOjetV6glqkUsGZPiN06mHGlalKC1ovy0CNnlwHeWMt/kiWfO5DWAB
TjwGf4FyG/asjZXVI95frW5xrtM45l/I17dgJGd380018qyA8W40btsq7oSp
nLlniv2aKxXnMys4yqbycj75ql4UcmO6tC7HfGVIkmwzJPGYL1dJYKicRfHd
k5rzc1z2xgbIs2cJwY7WUxp99rIrjWyf3P6Cfh3AVqVvh1gUgcaGa9rZBvwe
TFd/kk8sGmLDF5D9iwXn0+Y4PoZpVAUSKUn/RkG3skI1467+R7eYObpgGQ1v
72tq/ZHR+QgH52+YoeoQ7u96E6e4emRTnV6wq0x5SgmdTNMeGCkceCfJ0tKr
Hz9744qQrPqhpwCreTmtRgwp0nU4O0pIwlYCjkGzO/Hh3f1GUzxEfJHH4l4K
fBJYEZdJVs0nVtqXqeM9Esy3CIJp9HmkeOg243wXaJLd6sNDmjQQg7vww2TY
x0mgS1SeS5xI8VbVFzppgaMUWdKiJP1zgfew470XYSvvEjYPTjIie9ez/6JT
DlBsLIYaTNKOo/z5ruINtYjMPkGxu94PWVMUd+NZj7cnGotzuIYSIjvwM6kM
X90w5Cikb3KcJiPhPckDlHxRcGclcOpDRk8Ok8kAPGfmDOoT5DmeCc2qZl4h
7+BSW9+oeBkCaSYefw24OmGWeqOqCsTJU5A2rhJRH5XCvps5md0HUx3wRPp+
grWj8RYOY+RXMV14EsrCWiVzyOV1MTWpBqLI62PIdHa6GT4Be+LRIJnbGVRl
tKND0IulmRaOJphS1iOm0IDnsk2nczdgenorBrkLAObUcmEx+ZYmBaMs+uuk
loEjm5huZaA0YYN0/C30cknfHoSTj92hKSEmxINMxYIHDQX0K41dWd4WWJjt
ep/2zhdLTbct3BiZc2B3nll2yVpcO4p1WlTCOCF6cdyvTyhBQEqf5iPh6OOP
R7qkLGvkMNlMiOreuBx/dSbE1ShmMkY7ijfYWF5jDG+pbj2w6FdsevJzuHOI
PGiZRBMSdlXMRJyQyHGmh69hiuaGgYoGEXQQzCPZXir5qr/eZ656q5QDg5sb
9bElF2hW0SI7uGH+47yKcQpjCB9WSukZ+9Ve/9z9709spqAm0F8kE4XYr+sp
2uhJ3rvdVxEOaab/h2WgKJ3AgAuvSDQAsxv9jY3uvQga1J9ubwNQ4bJQFkAL
GYcnIGkkzytTiWnLjP5XdPRPkYIzpPIQioFwEEgI6qyHwwEwHFYDJlTpQlhB
d2q1DbFuOUwvzex61xASE6NEfg2049/JIWSgj+jJDWi/eOPJVO/VYaiiXpXt
X4gawpqlm7BJkTVukyPIxlZLhwbnbLONV59cf7cdrj9cSPYMQDRL48i2/lR8
azEn+MK8nSr/Ks8c54ksQxK5WbahZWUi6mDGAfs+sE3oZwMz+D9AdMDylqWc
rI9jXIFJ0DXkt9nMymztYyGzr77uYdhsXIAhsSl3AvJaG/Fi3XNAXT7djjb7
OQXlEHslQXsoAgk6rDb3YnZbLkF4r3b+ey5pyAIuokcMySk7yPNXhKcB3NT9
RzQBq0fUGFfDZfTgZs+/MFPYt5JSpC84pxkQAAtN+v+5aqQ/x0AmcM83fSQO
n03EPZrrjk3qNLEVpG/J9+/BN3uS7PI24hR3+Sv8mCNAu+UOxxUpjYdy3usW
neWR9f9Zuu4IF9sHX6FopnPFqrh+kSjvAl1j4B3i3ZaI3f/eGEUvzTdRngHh
JxaZx3rldf80WWT/aWVtNMWUSaghZTa5x+/8TTfei+1ifaexfx39hg6yA8tq
rmyqv+vgfS7RQKYXD4j0v+B8c84xG3G2ZpYHi3aqH755xu/gNOc7lylNjR6F
z+D3BBZzX9j3gC0Qs2cn502ShXWepTZB1s2xFvvRHU0tXOYq3AjucnsDDhy9
3bLJeU0qD9WxCLeb6Zdh1JfePAcNvGIRXMlnCkyRVXCi2SL2hLh/jfv1vRql
rxesGtCAyH4ZTLzr4NaJHlzbCt9oe1dEd8hqyrQGVa+JN2ZWj4fXUbB56N+W
YcNnYh1Z4Dk2w8FZ1+JpD7JG82En/P2t6J+X9aNRLQw+zkcV4u6Zw0kliQEv
xIa+G0QKeJPGwUE5H/KNLqNGvcSEN7g9RuJuBe0zl/vXh3bKDfpNdUq/xtb2
woIGeqkkwxtwb0qzP38pxOmX6BzmRRkoFFq8rLyuDINuWts4VnNt0w0tMW8b
dBbkJdGbKMXNhpk8bweVIlNsdnfrC4iVz7XiHkuwQzbKt0hnmrLkGE7xLm78
G80l6RicAn0MGYjlCs/sHAZ378GyLQY1Nz7xzcyLgUpLuWxVAOybHMuW9c9L
t8Pt+roXvdmmir3am5v2SpyXISKcxkBacIxXYuoYE65yxlHPjcqiCu/U3vU2
gvQor02Xy7h7YQukAebiixUNkV9kM8TcT1VbcE7dhyyvk9pDMtn0EYUGSj9r
tPYBek0ykFSfDAfbzi3Zqf3Bw0fJpsPWZxBIlmEjeoSNrhKTY4Vt46nJV8uz
/s9WwIyxp983FDuYP7mCV9RFGy4Rp/xSdKRXcqRBNSXZ/V+IA8xAkhGqI2As
Y+yD3NRDe3m8fd5SQaHPibaj2MZqfk4LcKEEfJuPKg+evMhI8PU6PVinbtAC
xFL+QmvcFkaRFvueKBKW8JyRsaqSBxi7woAl5yR4F29EF3l5T3ht6T29df87
WM4emk3/hA1IfQ618dqmxrn3FVCbfD+/GOGtyr6po1cWEWKTxysMwpHWfM9f
20WfASLdGrU4f0l1y+/o6SnbMcO9EPgPC/9Bk9m63aZeFmpsU0JzNKRJIcOg
FNJ2IotSPGzdNCUHZDfbF/hO1yXe1P+1BIjqe5ELas8qt2esW6P+P1Jh9T/u
jp53KpIVrtj9TPn3wihr8c70KCzpSlEGladVY5pPsz+dAFGXy2/ZDlxRmUXI
dRtELZNKWjEcEb1/foaN7NvtIZe9wF2cbk4NfRi0O4OpnPMKwg48A7WTk/aV
1yVtAm0iizAogMwpNvRamIlfyhogLgWOctRuaTmawehzj3DbBSM/Wo99pRdR
lTBgcy3WBhu64/SPl9zbgkSOASgzNEKlw+ujsyhyFqZVdmuVuq7yZsKZYZaT
xenMAfdE2QOjSWRQb7GaBPUN5RXg3ij30PyuivJvPhlaCYR9Ie21HQdSZOs8
00osgG6W6Cr7D9uHPBeiascEkzBgbzVKj9MOjKWgmCthZjCPAFl8haqXH4iN
V5JjYSj0Ee/kQfE+cUNwCF7yHUmUyLY6Le37TOh1CBrUbJ848obWNC7362Tz
6YKpJ9wtRDe0YY+mFK84VGfEvcY4+iMN4vr71C9XScKeZahh0fAFmP/OaHZP
4EONLx4ZmuPd2tBS6S/dpZLMuj5iyN4TJHbBtfULgTykL2oON9U4pnKVnLse
Dkwshh63S1F3p9Ddc+SQ7jntNBpamteN9rF40vtnrjh7vIRY+9SKO1ed8NrJ
D1wf5JibicbYqh4UnL1LwX6I3jWrHO5pb3TafKD/mINt6B7GemfpPDOjrcsz
jR2YMWa+GWwSDvKvCMp+dAiKEY14ij39Aa27RErnS14Nf/do728zY4MDiFwU
DXHsj9tjKGszAPAXb4jelYIM3+yIWFvBRjGpx7zJkphyra9/LJ9ZWlF7FbtD
BE5falUsxNlb7Hc6iGV15gxwT2HMmYT+Yqor+9BuMces3FXsS/e+NslKNd7z
7VG8FjY6FZv09LwJootN5bPntMYWDWo0kpzP6bASFqLWoNcnnpCpSKuWGyOC
W5BbAMrkC4EI6dkdbgiVa3Q3bSKHDyPC/Il4LkSKLWo5Tfo0/Q2JcsUHAPiN
/Lv8RLxXDkfyML+sF8lbiRxlYGnf/iqW5t0fge7PiUvBkHUVMSNER6pIfYLz
LrWmKz0UcnzOrbSzO4BnOaP606EBGLDVeZcjdTMad31rYpZkG6VQSKKjw3u+
F3HKO6GrmvEbY9EePR62GYL/Le+bxGpx77kKVHKb8VLQH4qxsR6RJKd5fK2C
Dxpz3UfWg3x9adAU97xs9mxOYLCLuqboL62Lfmt9hQiTfP8Eb1Q7yBlPaFUH
MsodBW/n4c5T0ca6wyZ7swENfXek1eKiigawGFCEmGLN0UBS4upvT7Ionoe8
Kxm+uM2DAMM4x6+A8DLRQajybFAsH6TEFksEVzQjsFQd3YsUPO9l4RRn9AlH
+XjXyaJ2hAGVBCPhOWxew0nTCeu2VxV/7rUP0r0MSHDjD8e39mP0Bw3FXh2R
cPU7AYHDU3Mwidd4NexleOKuMhWgsFunnpu7DEMok4qnyC5T45SuGbmLgePf
ry1Px6QITAqn8DNI1Wd3UTiaMfvu+dlEE1/VHkV1UEzA4Jd9Q/RZCZknRwLK
/SxwBAarTESUPhuGgVpZV33rH6RToHpDgK7FlRnzM1SjBvXrFJEJb012038r
WAuK37lw2+kfaXvq2NVf2MC1vjl+mgsRdq3lc53+N25BneiwOw0+vNotWknV
WDGr65UyYNNM7bcV/ie4k1IxlE/U3btp7y8c6eMYDFS4z1VxQEgph3Ak56SW
JaLTVHSEZ9n6oOMTyEW2gxOKF7hGr6Qv0QUFXHS7nF4IZErSMPlczIaEEH9s
lAcLrB7qiQ089KjhnCjctA6YwltGzzaJEWZAEbLVBIK76siYd8LI3qSiyt9X
WJnsTmhvBMK12dx6RSO7YzzHlXoXw9/vKNJ5A02lESpuD0PZgQSkEL0VLOrN
dlOY1mqpPjDqh4fQL3FwC9bHNyliawUeDDpSUgmvOv8dy1Swp4klnJUFgD5I
G6RdYb4RnhD4bH05q4rIV+INoBJfr/EYX6wviSVIZ0UChVME5tx2y0WKyZCg
KfSJgsxN6KeCyyeJBZH76hcKV46VRgVOUuY4uqVvKRbC7tqzwE7DgDaAaDFh
IZFpczzCP6uijIJu5K4q95mu3WP4Hiue64r36Lxiu6a7ATjMwBHWyZDOMJYa
8V4qHQlyJlgM+soFTiwo+mMJRNkTHeUdsmL480K3v078jVFfyPQXyp1jvViG
aBw1IdyLo/sBhAzMwnzo0eRnqZEOrSWYyq4lemTi08HdvGuPamZs37rBOiU+
9ttCHi+wLBBC4GW0Q89tIKGOtD9I0GGe6bR5GNz2sbCn3VKCHjeobbeoEhM9
mYlzH91fEwaH9P3O6xhIbD4OkaSEmTdcMgTaYAJfz8kqPTUFnGkLDlw6qxuv
vXVbc8NawylJr/9O/1b3oYlLuJ/UVWGZv3DWPvrrKlWx/iOiR7Aomw4oLRx9
25z7qC3VwCW9scMea66SsuMczZQh0nHJD7q9xwhC48Gjz1TxyPbWL2EXLAZj
TAQlsBi3OUCw/RBsGtoMF+SpSKVLpZTU9yGHPNtV8CL83JN3rWu78Fldybli
dPi05vkkhmNBaP6kYvQrGDLpwck+1S/ZfjtwkVssc7nKbpKVdkl3aji9Ztw8
/JGP5jcPN4MaNjYOl7Fwqn+vt1hRXjJDk86wOdZJm+dBRKdIBTWAUi5o8SSs
23P+P6R/wPiOXikdJ5zQaEeBT3auwPCeTEnWFgpwROILusosHEjKspJdx9s9
cW3LPNujQAzC+bDweAEDk2LP35wDzf9o1597M1AagctC7szEMARfbKNeHgv2
4j92Px65BqGFTbbhmgGqfqev9qG77LTZEl90TqkykDfVw+sZvprQ9w6ZasuQ
hHDbIyIFnMCPG215KG5hXrbzYYKaeeVXP4B/xZTVXhwbk9sinIi6OP4X5Y9O
7qRDArftyrDKiqeWlCgAoR8qvkFQK+ZcnKH+LxmIiVPp0X/JCm1hMOH52mUf
NpZgcroK5TnkNttDJbfAVoGIIeHp7h2f3fLsayECptW3a/pUpaYfTLZKtrar
RymVpQV5wp+NrOzPx9htqEntZ77O/Q5uDi4qNdgE1P7iDruspWB6gddY87YN
+tOtw30GvWLe8u6vbgmftHRg9xLnCL8HhQ3n4ywPnEQo6jApX4b8mXLJjbV5
tAvUMZMGUfaRfnIQMBv8b27YL4FL+9SUSP2WhUhhbHCnF/rbt1pqWzMgRgEw
7SDzM8WfS9rys25Pq1SwvERLu4DjqmIgasSC8LEgvU9tpRiC5XQ36CvDKKIJ
G4nxDcwz0LeP6d26kai0uCduGNdAqkev+nMSxtazni/OtR9iK/pzBpeK5rXs
peNZUt7ZsU2rIS2YJmtx5LlhDv5BtPu7/wnhC7Upq7ahRp3yYM4iXwvPbsq0
9YVKavvNj2g40jhVxQEiN8JsrtqXIbdg9fbQZlCmbTKlOnYILCqVWzWUo+4r
usim//4tuSOuynmGfN/P2axosGkdPDYyzqgnFe/ksi3+yWHGnAoRACxNOaQI
o5S+/rnjWs3qTRBYjXWhQ4dApg3QNB79ER2iBkWrsuZeHZ+ntJfOfAOdjH+H
ks4//9ptJ02v85cNt2CHg/RRmnRpF7pfESuAy70DzRFSfu5+4M/Gns7BaWyu
EOnwaDAyuF15XWNq2hA7fNKbIihaJE7Lj4K7vYaBYF4KRjKAfB1MlCTjHSOd
MuPkpwRewEoV4Q/X8HSXPSyoBbz6kZ/JWpM6lrONQ7foYPBdw8XV3SR18JNj
KP7flOLiDEGrYr4Nb0X0XR+j5hWayHniFbGKcIMlJg/QgTVpa4+rLOt0+e1W
79w3qFX7JsWPXWH9tZ6w1vzkzsIV0TzQxXkEyJZHNtU0rIJTx8zYrsplLF5L
7ZzK1eUVVtpUSyv6cLcRFdQGFG48Ih6gyXUr0GgvDqZOZ8zpCnG+VfCNxbzN
8fQv2yznIQQblNaU9wZcbvzCo/2SYIyFeL1DD/M6JnzJxtbGyA/i4UPqLt1T
pTLS3HD6BzQ3Tvh+BsHAPiPfjyg3KBCMjt07YTpT1A5MEWXDTcELiuTSY71/
HiP7U/H9ee+fh8Y6EcP/twkPkAhAjc436UWVkT5xjvLj8IsSB9r/dW2B+8DN
14GYcxkxFEnhMB5AI5xs7lgRrD8ib2ASNk5QrtNo7hpoGyX2hVNoGhOWgz9D
qexwgTqY9gcVLNlxiRnnaP8wFAshKMyRrQ4aSfeqR4/sdQOrhLRGsRSI0b9Q
ePowP3vZugoechADWIChUy643rlJ+Tmbw7l4KhWVGfB06/pzuye2Qpx+RmF1
LbfS3HdbC2CGK+6dKqIrlwkI7KaMV6lmm4uhAmXgKjxUa3esJGfm8+ELE3GY
AyzbXK1Z+b4Z4sQOirXxSDQKnvpQQv7upV3Ega+7LhWyAdYR4jtwxnLgM4o4
G5lKBizTj6wgEXafotgNIBzrY47o3cAseERE8gXbGZpQXwXszRKJbK7nyCKg
OyIaOm1Na2/rcBHBxCqYfq0DWvKYzXy3yZmBuzQ57ADJS4ZsJy/vU0farYxh
ObYYqe2+eDb3A/YarEujMHxSzQ+/K/mW6l/ovoYzc5KCGLBEzOWYoYbAcmsx
aCwDGEgesNuzFmDxmRo8+N/tBjArMe6ABACdjvBNuhutIF7SSkLSXBCjCbM3
53n89nVMbFDlvfXP926MrHAr4/RYt6FJDV78aUwuMi+tfBR8uGoomS2r2o+F
861Tu60ERrr13GPClVclVkEpYLFGBEVIlAOsvg6ho5y8Qjh6laOD9gJOAeRi
uTqiF7PQ80wG0gW3hWhJNb+BIorMcOWeOf15I3vTNzhZ6nY9/aVGAxjSb/hs
+I6ypAzGS40MqqCmwUbYZagdGHv3UMZguf6I3LvrQZeWCUkTu4niVfXoSgsq
uXF2cH/RlEJZN8VPgcz/92q97a6WA4JCJw5A8PZVSiO7N4USvy9BHu5ufDW6
xv9kPqA7psb5bCKMko41gw32DqAS0nTNw9BFYAu7RQSxWzC/os5Use1R9bP/
Cc4aZgINl01+lbr9VuFEqMH9RSyyGUsfmMLi7+7IcbbfsoTxKdAT+hOrwa0/
BkKnVopVlidJ6rxFAOKvEXDjUh1slvMwFjwRF5i9QRVSZ++RVhmCHLvSo+Tu
hNWS4cLvFDLjBVW1UPj1GpBmRd0aDoG0Jj9MHMPqw5aaDf/VVWRQuRqQHMUD
pnoElWad1d/EfE282jUZ/MY92ca/Kb4wWmQDAK62GhbG7pDjvoQS3zxGnU5p
WYQhGibVBInvbuUYnPxN32Ir/0FvK+r46iO0TJ8HbUPrc0XKfLO1KovHpdLX
9/Sp9gW2LgO4DwNaSitzOk0ICZIuwGWXNsLQVWIt99ZaDjptWKDnYaWXyGUB
c81T+e+Z+ywWeWT1Qwtd1GEKGaCxvSES8rsmZkDo9Wwge8qHbqx/miotpwfy
S0VZFJEPv/QcDvzcHgcK3MIM56gCM6bTqWbzMadf8v9W1VJolmWwXNVzfG9b
ox6gYUYeQE7KwUlVvPT677RUtCTHXgqqbp003EWqdGWwuObg35i1OV1KUMu1
1tyO4bmxymd0rJKcQzhqpZxmsQ5QZf6Ak3h6ijCoD9p8abuHIj5dmCEfOlrP
G/GL6vDueHTqftBBFPlgO4cpjmXNbgONdTXXMUoEDus9XaGNDyBF6MfAKu+S
bpj5HLVDcTjzTlAxZja0O2B5Hxk1V+3Q4PMYrWjfIQx8nGATRkxX98UVRYif
7TurHL/Kf08VI9hUKRo9dy+J80u0koJtGPBk5IZRekkOUnWqG0l88TU+70eq
JY9w76Q+VXYfQRly0K3Ov+yll1w+l4KM+ZAOK7V2USlrDS9BFNvSOln+Ovuj
NwxN1eiXhpdEWuPLZU4xeBbeBYRGUJWZT9Q+4l5pjMpd4FhDjY2hkPA4g0zN
8KR+HLLGU/cHIjlIjEUmUFUktJh6eaCpl3JHP16ulsrBm6i4sp8ojL4fD3Jz
F6cFQnIhjwXkuvOwm47AQgk2iKvJjKKhhsUVVNuhZV1ju9UTNdDH7WwQ0LyC
PvZihp6O05CexaviTpZQuqqfD7hMGX6w2d1PhYDi1RR18n/kuA3huq2nUlno
FsAwq20uEahNbsEHq8cbbO8rgmXVKaOxuQfChNqRJi43YQJ0hI3ozAPeGIxi
/9Q4mazy42tuQEP2gWLzBuKOSCI13mp9zbGmas4UOwFmAcgqudfcm9fd2JZ7
NtNqQkUIbvTIHHuTblINzpVX6beUQW20Fcq5N4wQD5hKh0pbzGxwtw+kX2t/
eyyFs654oYbV4TI734a5LeO3+jBesS8G/htawyABIUHV+3Uqjq3Y5VqbMiY4
VkbfjIQCJCpdbfmheEYIgwS50UXpNYmcWTZOaVTc/lA0652rZ3wHHcHwSo1t
BRt496pCbVWNDNtg2/qV9pFT2Q7aMOCmQ+63c+e+WGGuCdVggvipfC7glZ1k
AbkhJtshagVk/k89JvvOr1YI/lsVG6xVhk1k1TPoivgu+edu+kTVzSRdb9To
aAGUVVWnTbW4YYDcefp6HPb0MYCPpGWajQek4CgvsZN4+I18+rKUEQLMPVmy
o6Is1/xtz7OkiISseZ4Da50sbMnloXwqWKVj+KrKGptHn6SpL0i5kn985KNu
z8JMr1YKmgwHsT7NQ7rdfdAXcUxU6fdZcZ8nE2Yajz47v75Yingkg8fRht+S
LQ29CtHvmItmaF/+jCBRtQtNthQGtNSRMQBZnHPFE8c4+l6xLsbA8uztyTkb
uVIhLAOg7t8yO0Q3CSQD9mKqYi9A3PxA4f2YsduKEhv8Orlr5qWjOWMS+XMq
roAWh3tPKY2z8EonUWzSX0f9szGgZgOFHd126k4szTfPYDvhl02B9JMHHQhU
4xxCl7ig02HvhHIGWJG81e5xBDnWOr7KcojNdW0OEmFUewv0e6TJlE/8cgvF
l5vbQNDpqvQp8h3I2tmznd1MmshGTAb86FGNJr2KAP48ygzmGj/F5/KjOTny
u/VlywJpwl/1eYL656fBJSHWjHqSuTzxwOQ6zOxCZtMYpkJP7/a9sXI+RFZT
pFeRXfKq123UxSdTdRtnjn5IipzgwuZYbCPrmqT1AHfkbGPeRTK7hw6VGt3+
BSn4pEtu4IETVEEltveHpk3ili5BZ5eRW5hPFlaiRDs4VYN6oFsvmGidzOvq
FBcFdRSrs5ODKkqXTozCpjNB0dzSQ/zC1je7lHV1+MLpvfqGj1lCQXiTUvtv
4L8M9yef8szaulitYpvmllgXZun64l66exfGOR6YKhidJQZ4AwSwQUOGkg9E
e7Gq6i8I+U3SG6WaVUz2A/2vd22E5zNJwxP1iOm6TWXAPr+4mEcOX8znGm3X
x+TQy+K0HEcH0SyTNJtb1Be/ap8ANzxLhKzWOUxFmAtmceqreL6lsHPD6iVu
L1UP9+cIN89Pf6NEcptrQZc4ar+HJoE+1BlS1zMIXSKzbPzR2Xc2LCIuZPol
bKDjSCwJ6zx5JyLucA/pK/aIftDCUkK+S9puR0RLmh2FtQhobumqjde3SLFw
jQ/WqujlDbRarIxJsvT4VVFrfiDl37ewz1g4MT7RMApGOzj0c2rbjDmz3IFz
/2cd+alt/l5QhoweGYe1s5m42WZNGTJjRaTElkDDEak+lkdroMv7qb/cgYzW
n8wKVZkT27XrN3MsPcLUaTdM32/yXvaMVJ+1VjTCVM8kgGQC2Js8uh0PO7O+
y3h2ZndYcSNA9TrVNSaoDMKDy+mpyfdgjWFfrU3O/3NuhywRuxXmz694FWb8
w85A1G7DB19f9l7x7yRJY4BPenzLb5YB+7YZ7EH1/J0bBg45ACPBF7b5YaZg
OyMUIleYy2ts3/2HRvzSd3v78SM6eq/9OmN2yDbZTwwakNYEXKWrSTa1j/w3
rPuIbW8+ZO64fwbjQsvKzaYTYaRRq17I0tvOy+xQuxTCpP9qaZsUSqgwy03v
Q+DlXfKD/CewEr0g7S+VKmQGGhYLkZ4uD9gIkToPNmILthvBYquFmIol5jkd
Z10uIW6IusGqiiTEvh+epTsQ62Pwk67aYeq61BCivNPpHOgtI4zvOti3FBDX
LYvvI27jkuIPegFW+JfKcyMzT32guFmpHq+blXm7WlpJjvQyVdlK7SwHw90Y
OJLH0WydwU0szKO6JFLrvsfxw9eltjUxTMV9Qk3nWm0jgZ3sCG39rGWibrRt
2aKe8b9ugq6WiW1/6g/Z4vMVNS8BTaUQc8vgTZf9u3AOGmN7xKuIk1FY023U
vdpv+g3fQbQTMS3g3afNOLCdVf5pgAw9XwJr2TKt/QIdQI2MKA6nlQ5bQWu+
x0r9WqjJCAE6qwAeKoRfVyz++Lpk4PpP377wLTFKtpnRX6w4Wc/ot4EhNBHy
UwYSGFsw9ggsZtX0z4hbnrRHcmK2ICFq8KXaEZNTV4lz/hWpVOoqG/G33fsr
VmUBXglaCNIeRqaSyS7UPNOG8Lk4npINU/8c0LlSAJzauw9oYBMxa8169hMi
sS2CrgpviAXLLw7wDH9LJJ1B9Conk+5BmSybFI8wVKZPEx422jIqRoMXaRpN
P1tIHHlSQzofbMvl41zkXMuslsWWwaxORpw7tXtr3AQcI2d5NrI5p1URyZ44
rU5BexM5J1DIFkox1VU3W2v0lGxRVyGJD0BE35GAxEnGQ4aZxGNFgJYrXNG6
VtwVNR+IMYLl1hDke6hJXBVLcThIEz4/IZrJbAmxi1D+XxdHCR4BARhIecMC
BsdN4mIq2TmTWV6+H3D4TgG8rcof1gC5/BG64x5frm2AC0yp5b2xFPI82X+h
bFdqKvr9MORjPykg+t7S8GgXhbyEuLURzW1JHHaqIQUxbeyALKZBotVUuRZF
KlyMhCrybifX8nYwlJup3GvLvOIF8qYPDMyrVc+q/86PGk4+z9bFNkRakS/U
Nqo8uOP6XERLSRtTDK2Hgq5EjWOEssttBIVKAxhAIYqRXRi9T6tc65sA/oMw
7Px1dzBEfKwlYFE4tSGiaKSkdZZiVz3GR3LwsAY/+a5vBxobCeaKTbnh7xm8
ShajVWBVLkFn8vFWrYrTahXqAiCT6PidhHEvnMn6PH/u6Ine9mUQEhpf+9Fz
uRA4EYgBMai+N7N7utzypXTstyhBhrN2d7zKsGtitY/qJQtWwbQN8K1UeXZ1
FXaz5uuVLQOyIMYrHHf6K+4J4hpqCaSwHZupmorDCoIFi0uZVmz37AbF3DV9
MHg6V6bgAwXqD/pu0bmcBqHEdpC1NoCD9aqWmGknlSRRjmgQKuUGLYPbJMrP
0ECz0O0uYTv0LQp4h3bms/Sl1iPNzv6hz0ofn17f1SEcA+KuzZCpaMdID8/G
Ua2cHZFyvczWObeE7qH2hhHso02TIA2SXMhLcY5B9DQOdz3Ly4j8PZ2P7m8Y
qGSQImfY9YFgIcXNriwZthA7Y2HXwIA63Wp4LoO1L3YdU5NRggOz+sxrga36
0DXBkiKiHwqhUzwPmMqtF4ROtunpeCQO9yOu1+szzSpVYiS2DPrjvmpo/Bfw
ejCeeTwOzvkRfdSGzUOqBsEUg1xqtdfn5ONuZF9rFXBBRErmhZcmIbRE0c77
Ec+lMwvsu8DLDdlT71JeGrZRkI7xkuRK45wDm1PfGQ8OaiQMXomi8igEIb2u
jkAvapDak6JIJrorXC4Z9SSAMrsyke7NnuOa7p+5jWupvPzoCpX5Q+djh9Dc
r5kWB+JIEXZT3yytPGFfbWWEFzOUnnVJIJpozsJgMV93ZJdmZusgOubmfa1m
Egzn++2H0CdulXgnSZsEjYyN/o1LxBkd06r+f6wtzQLD5dk1yNDV4Y4AIC59
Z8hTvaC/FFf1w4pQ/USpY107wA4Ofnb5apjk4+aWtCqJucu9hz9zMQXdwhiO
VcnbSdedq8oMiprM971yl55Om0SVOPlGsfIx4m3GKLc2Z/3vFMJLovyDbYNN
oYYg1VkVlivjSytHanxdVIXg8uXBcrQOn02GbIaYfzd/XCF7SLccF3fYyO8t
XmcnPOhpWR1R4WOTwDvAkhXQiXAFemb/7F37w+GKJhvF94lbr/30vpLXvahm
MalnAXd1JMX0n0XGvNQEf4N2wHJ58hhSCmAxzhdOlwfZTSIeQMbG1EVx4xKq
QiJIp5l9Hi78wPHaeud7CPVHNqH/kHhMi3w/ixb6bYCtll/vUPYb1dIZJ1Tf
CYN8PII1B/kjWyBRMQAVxze4A9jQ5h5jj7vMSbSGzEjLkktrUyY8txwugoBP
hv48SPDVYbQDEqKSaVKzK05lOag/A+pYp5naiOPdMQYhPRtTL2MW46o58Mb3
QAsJElFueEN/AgYj726/4xnrQoF27UKym72C4EtY7LX99Mu2TL3aohqbAU7R
vIMpwg8gBhOtXfxhMetlNXo2tp73IX3EE9rvuIBzmqUPMhBpuvKQlNPFWi3L
lG2jDNm+N5xQsm+xJl/mEaBjYT/EUSLRYi7kAo+ds9XUY4PIs/znZf8BwkEY
sKy9kYE9BL6o1pnX8OfxH4CQR1JqUuxMP2xhThk78U4BXgVKarcD+IzuuxsZ
QwtAMzsakuwEi0ZgBw4LQpc+RXQQB3UAAEDER53vtR5+s2UnA/ivFx48IXHN
PNTVVBF6tnpI78vAfsfHKak2ubdn2wWeAn4a8h6np1tHvB7uys1fPlfHVgYB
kdnOMVzB0Ho8Av87k+pLLPW3rVtyIgqu3woM6P5L03lhkS5KVzpYPMnLHjk3
CzTrOTNmL0pYc+inm2dPGoCp7LY0yvNCZe/DkEKrunUU1Fe6BpmR+NWSV/Cd
fZhw4X/nZZ8tCo0g8jPF3dU7AwOu9qmZjP30AT4bj1M/T1wCtoS0jQlZk5LL
LxlBghfutpS4Fh17QTcwTm7DqZrHMZdn8RJcaK0eeETuLBnTNhY9meotEWSp
/q0ejxdJTc9z5UBBH5/baAIN/ylL/bo3OFe5NKs16hzjSF+kvZWXjP2SFwuV
Nu3e9HKQY3PmyruahIUaj+YKFjymVPjBA623GScI7FMtTmj+pSpoSLp2Ue7l
+GxsXPo9329eQXhJ5n4wL7OjvyIrny5r1ZZGXocXg15FV//oKv/VBLHpPxFg
6NOsyfiH3p9XnjreZuD4Cp1KDBaaajuWSTz45BRj3G9+7/UEZkzEtCOboa5F
DdOxw9zyO8kqL3+99djx6Hgv2Sim0S96dg91h5Xfamy8zxjzWbQdjmV3NcKz
+gkF/sGSOq+ynlmvIvpLMtJGylOvfid+WVDhFD2ZeeJkbmfzU/QwCh8G0DFA
s8GC4BZZdQYOzWtjTn3/GB6cdaLibbwSnjUo9KCAJWHvBjNrrvVpK4QE0oLu
21e7gGp89sR2W9hbQkAxxkmh0FIrE7qFbffYjaLq71lElttK1AVJ8zqGfG/F
e7ASO9YaJUy1+fP4BJn7vXBRZ3vHNEf5arrWsv42iAwvj/LZ53Rm/PJKp681
UGao8mlGqq1ErMFC5HdrgqIhfaWYBsVK9geDFCyzHQvuk44ps4wZesNrDIkq
zafIgDo7YuPeXYFXCTJG/+Aq7avlBTYctxZx09gt+yy0xiuYkhGlr+5UhZ06
hCQKZeHJQIJKpCKH5tA7WLF3FV52+7tRqwT+sJWh3Au1Z2rMmwNe16deIpMr
AzcqfCP326NZwMnERcGdTfZcaONhPdxACo5MyJui6Au31qLp/SoUaYhO+IQe
GgcPXHE3+ANPq2BTowfRjvH4CL8Bj+9o4c2C6oB+ub95IJoh67/zfrLE23sN
dMuzjYJqDr2WYQLmTqlcDUuxTzIa2O35KECbYH4P8zkn3eA1nhRQayzKLqch
PqHKUb62RYR4tYrXtf8lDAS1RH/lb+M5A/gBN30zWncfvD8kfD4MNEruPjQl
9l3tnitd3VX+CbpCOLMOD5YxJZddbOdPUjuJFbzANID3j7ExQg4XND/8lv99
XlZewtxg9jhwYkkgJBjjNRBp9qau9uys1f+z235VF0Ez++H123EQnON+j5ju
alOwHmbNTGST2EzhJJhg405hFE5x7xbHV7XwgyfHTfi7x/5y2qRgLaR86hpA
19s00AqgLK/xcXeuD9FuEYx7ljJHHewHQPGaD4FTggg21wA3Uyb3Qv/JdcGf
k8hoBjUJ4lS7Tz9rcP0RCqiw389GA3Nz1OhgFal6MZTzqhleXC4tb/80dXb4
jFmlzycdSiyD2jWwpfpoG8EeWSU4qjzydTjJ3yiRcN72d1RvCw7xVpj9hQMu
T2A0lv9xHLeKLJAKtW3iKAmMXe9l9q7iMcy6NqSzQG/PAKlFkB7QRV4xob3R
ePXEBVA4XDrjPikPEWqW8gB92whnzw5dnxmpYSdBQ2LgH3ESlNFBLpeRs1yi
ywMvPe/oX1QO6NSRCqS7X6E5ZlmHzr/bxE9lLp35u5HJKea8sOyDZ20A7VQH
YgcvW7awxTf8WWxDACFPyhM/GlECN0qQxQN9aLTPVpaorsx/XI42e/ajXQpI
S+w8jc3OezkLF1Wd0JFOWK0gJIU4VEovdJLGcZs4o0h6bpeQaR4NLucqJVbM
ERvCeuIhxTN2kk8TsGqDM4OSg7e9pEY8y3QDkBT8J4Xm0MxKVIFVg1kltcji
n9JSCoYREZx5TS4GSLnK6CMEHbmmGIVKy9WNH7JBNJ2AFYGZ/v9+3qF3pTav
ULdFxqdVdiUZCWsFoN2inJMeAqvlhc3HyFFG27MIJQEmPRibTo2ThNU5roMh
PspiCShr4Pjn6X7hag7fIZ3YMcUV8pETXi5kWQWPoB1qHJeWBNIIoG9eKWOy
7pLgH9D/kkdJ50z3dr1znlXAdaEuswzteFfFBo+jC/JjvAEdqf4ABoLfLQbX
pSucjilCPSvVZFU26dWsxnfCEMBH/emzn/HlBWPyFilXem8mO2jCrvUc+hKC
8CjsITW1fLShUn2ThTzN+vKTb0kHD8t6sE4BKVWX9kQqQxN+7HPqet065G4s
On2b/kRxmR8hY/AjPlQZs6UtR5ZDNfqfjBicYmonxYx+r2YvVrUzSrZXD3B6
r1z4vybxByFaYC9cEdeJ+SwPNBYvLShg3QMaBFv+bYR7W5X+CC9WM4T54eJD
WBKaJG4zINzN2D/bqS+LtmeouEUl8gsJR7J/d7bwx/Pq0UvhiYvBDpeMPpdB
CHQJzij64D27HDEQrYkmvG3sdb2xlgqJ6r9u0Ye00BXH1n14s4zNQjLL7Ol6
LZR+u4y4GuB8A5ltwmexafOnRLkKLgXYVpAzxPjnF1pvg8/D3zMy8yHy3hdI
yO7Ss+rxnvzfYCj2AWe2VBt/w0O6/ySOMeOITyvIy3HWZ7uoelHjyZDGnmle
8Q9BjXI4Q6b+GqhBYrDgqpJntRnSBvI8o2mCYg1z4x3Bxwpx2+vRx502YC5O
R9RurQ2h8n8fkTMPBBfGYqAumGqAGEmUYJi+DGGKsaSbJrgojhk+sR78IPyg
6PbLOUm5FUOMZGzsiouXTVqKnO3WS7xxBuXuzEmOj2orC6LeZpGODhrWjnQj
aoKJLH1I1W5jm85Jz2zTZXSPix8SlF2GHaprd+BQ07ZYvjmkuo8gZGypueSW
xd/8JIdW32exaiGwAF6uvt/A6EoVztmORYrchl8IJds0YTeGNsD0Ahq2KOO8
BNDW3Zu9Lj8Rd6o7GX5RiXsmAM4N/yyIJrQi3zl8ZRcY/rsVg/XLvjYzqYzF
BhzaW1PmDysEc/gllUoaMxTIi4YmnTHno4cO+wnByXKx/E4vxdqiO7pmbRZP
cDj5qleVfo6VoaMbVHxB9onidq+jKe/eIpXjtnf9Fv/2pQ5ujDybpspS3LwN
gXXxwxXo4KseCbpK5sHer2FBOFsf09a3zN3G6suzqD/fy/iX25LRsmfVGbvZ
HgJv0EsB25LtPE/IGVN56zOEnq9aHE78WOKLJGLtTr5p5OmyWtS15xBv3RH6
lAwJCRtH7u1p3/hNzXHyCDP9tTPxzLX9XXTJvwcA4eW2GnVRc5M+pxirG615
z+Vl10Yv92IQCxLSlNI77eTf9uqjLLf+fQTDugUB9MG1ofxTS/y5ABjOWWrC
VBqCQm2DhfYaP6T8Nbbg0AWXspihnAbjD7qh00a8dKnIDnD1O47yJjSfN/jm
LD36ZQUzPoqArD3FLVImPQOu/c9fYhTGA9uSlDcMLhKIxMgTnf+7mpVAyvLf
hhE6WepTOWj09E9PWbIbaEIs2mDkNdZWaK6fd04+xGyqAm0oYSMh4xAdX3cM
NZEh6/FCXeyPKm3U0wqR2Lc/h8XiI9b4VT19gCOnKKRAhgki5XoQG+VKOO0+
qmt6Goj3riAhbSRjk9gv8YOx2Jnu2Ztbl/cj3B7J2s+TrN5ve8Ou930nrTpe
d+DUncu3nH4ujfO1lusb96REygZPRmUl43FCPSLca6WjRcdfPQB0nN1DxVI4
pzJjH4rKLkMMa9lxGQ6XmudRssTucG5KEGMc368Bj3Ee5r93W1Cab5KIoTxg
dGrjSu3Yo13PD1AmffVyGEv1ygf8AW/VkMFjFAFqGFXHY+qQcXuud3BkdJCY
CqdUDlcoXWXAuUdYh7czDG/r0NRpZsbhwgX7HErNrVhU9ld8lMLMQQZcdfbr
yOzRhE6h0z7vjSiYjaMPEmAMIhutbRlUWdqxP/0z7K+VJcw8izBe8Jr8meQ6
1Pr84HL6kNk7MJj7CD3LQLc9WFkMGfjaEymE221PjZR3a2LVPPB9ozrmwnlA
j/Dq9enEFHgXRaA3R+JYQWHEpa6R9C6Kr38CV2x6DEO74m49ULGizPYr+pmy
AHTR0HCxejiiYRjmCMqIYMHfQXEh8s79ArhUmhv9i+rrDkCJtZJn8o9ASl/Q
e8EwEgq87twEhMh40Du0j0yF+e/nZaihtl5pIPoFVmDStYjbvPM3CFMEtDhn
N7brLeFt9yA7nxxM5JNBvjq5I0P2ZqT2B9kOxCFmkhkF+vUqShB2OydydJc5
Q37YRLayDM163pK3pho7d3iCAyuogaBBNBBLmojKqBm5n/MKOY4a7He6pZVb
6lceKRD7TwxpraKis4/9SVVywl4JNfwvQ/ZoxdnPRNP1JOxaxQmzHhFqAgBj
1leQ7LMlvFBqKroe+uHiSdXM7cTcYZBaUN8l1by/WTqpZBGT+IblVk2WJfgy
oK5yErehFwfRLWLP3OS7yOlesbfRy3eNT3CFmQCEI+GvkYyeIPuH8XEAjIEh
OyBwjWAAgshdHWW/CcUCYZnlkIZOmUhF4Qk1+cHQ50oIiW4i3TNZanu/bEaD
c4WDvPTMcGKqymRGd03IuARF3YK4jpkVzCqQF3zItHDMlBsdCOKriq2C44z+
77xt+cDEyF0851+6nGmBjKbBqK+txhj6ck1fFlB4IBSfZYGicQlqHxG+uwlE
ouiZxT5zbeNtaAfvRGBdcd4JVYSTjVziHYuLMOnfK6C8PFUzscnjJY2C72M/
Sv3iTG1OLpetlGgnshbQLfeUVwufjpLjOhUSXAciDbrTGbI8kvU+cb1BXFXp
7+qcc7kcPb60kzNKiflkMwmzL+iiBowtzsU+oKmKdzlxa8ZxF61krXAZZWsq
QCAd5XZaBuVrl8xw16lrwIAuYLENwa3ZUF84Sa7zvG7ol2jDWx75Y8eaQP/6
j7m03tUqS/9MUquFfbsYZTVwpmctQ80YxeJnqMNbM68DgRlzKaR2TVdRDYha
O8AWMXH1hFgMyjMX/u4469gxxbY9zqo/kSXNm7hUStNBAhIY5Q0+YfGBk0eX
1pzZjtebt2JDKSiOf6HyKZ+lZCiUeI8Zmmd7FK4T+O/7ISYa0FYsi6jt+rCd
yW2LqclTo7cIiEKZ+JSqVh29IJ9B1uaCX2sF8a2Wdaquh9hDfiGXVMnvu3G5
2Xo8OWWOn5k7VGKgrGWmZC8WfPv6NooLt7lZ2bLpE3qEWoAZSqeqWkzU7EK1
Bai2XEYHh9mJvf8X6ULZbQAodd5VuhODRbwuIVt5fvEC6Y2HoFn4Ctq0QCJN
i/7NVn98TvyyR0uISpgEoGknJ0CIWO+2IyKtr71aF0aS3pZSg0ZpLQOkVFiu
USTaSh1R93UFBtu0Hy9vmP3KmUjxCIJ0s0Boq/MiSXat4zCK4WKfwnhW07GV
7owTrSX0Q3CNbLEBPlGhuNvI5rCrzJv6yO+vrd3MujaqLGBirUBNjLYqRHvh
d6NMUbRr7l5oSr3BlsG4t3JZGCAZfgZKxo+gBvt4uniG+KC1TZi2LAL9txUT
tCbzpGE9IUJK/id+svUPd7ix3h0FlaQG2HOck1Ed0Ol9fqtQ94NSkGEDvUzZ
mkzKfVo2rcVESxDt7HE0uxPR+fYUgCFlPD/mCn6i192m9OCIou5JhgyyFRZd
R3KxfhND3U0GYRx4stugOpwL8h88IMEHPrSw695MMTNfW7kJ/5MuicoUjTDJ
6fPGo8ypXvodmryjoU13TDyMCFmZyUSrDUqxjgTUoSC4gjy25S/Bi6Ke6Xqg
MF6xuo+CtI4QKe4B+FaylHDT/GO6udbUmeX9+Juy72RyS8BgpXBCY5Xo6lVV
MCEKja1pcnWQqHDcZWO2yN+hT2rw9p0GxxhUtyX/kfmqOlpVxpmtRSw9RHNm
E/Vct3cPl3issH/vQ1uPe1hO71iM5zs+GPXlHbAp+jbaF68VlIBn8wm/5ZCR
Nnsf3vXSPqSQMN0XbqhCBM3f1Fpe3/3u+Zqh8yb5dYzH6gQBrLkZ94NesMat
kFcLl32yEAlNhjD6HZryupIQw9ulElV7qMFMc5jcOrfm7V/8I70DPGeJ9mwx
//ZP5er0XpiCZrp1y1x+NNuug1MZ64lyrKDDT4dHCYHeH7aPEvHkPD/uq8Sm
YjyW7+XpCFyRz49jo105lRvOqcIcloyJGY4/KwFeoGePq8JcsMX6kz+HmeDF
yM+fveQw37mf+QQAV9+Yt/pKieYP/T2o3rPAH4ur+YjNY2PryscsSLzD++GT
TwB3brDju17mcqwo8+edRWC6H3NutdLbALGnPI2/FeO6b7Ngtt46pRuQPU+0
oi94osHlCz00TwvWyLdnWxLZXaJmrGtuZUGWXeQtnYBxbhxM7wR9qSPAJjnV
DPmgIVWi3GqKKn2oTq8SbZlAdTNe5i1mV4B/wEYo6ZsZfAmLgA6eF4TtbOmN
+zrFnvTZJrpSaM9VApi7vrGze8IdxOPyYmPn/X8YUxSi52DE44Tb2HFZccbP
qpTbbs4uVuzqmrF9C7imNKnsNQQhrrmVcwxE+VgXn4tPd7vIQ/zAIJA3pjWk
1PHsZN2tHjfLpNBwsuQauXGw+oyKVBfpqRU6C6EHWEM4wPMyFc7A+YSEQFmj
IG5cAtdDym2EX80WpUroufjMBD9NbNBnCSYWMDSmUz4bMPNAQJ0Ert5EWjTC
CLxiikg5fccvCg5DTfkz7DhwysFiZYK6hB+L3ufsA8ol4687kwPMjHIeR2uP
YkAYPXOd0os4TwQY5LhOFp4PBrCbsAUwwbpMY7Y5lIqbMlvx49AmZfC1sGq2
8AJ7/xiL9/D/aCDYX5+z9vluj3e2zXxrtztoJW2g1N/Rcf52ecRMb3wXK0t5
lsph+MzWjq/yHxfmlzzLpnwdTe98GPSLPR15ZeCmj+GJtsy5cvpWSr8Ivnp0
RQASEryIlckTKcDb3tPK1tnzqmJ4uZOwajvKHScvB7qX+aeCyzQ0IoqvIlnC
ix9in5GGPmHTAeozysW9rv/gZineaEsJ6V/LJvsc8csC2fEpQStDeB/Xg4NN
ICnZGjz4Cc0a8pq3r6095Q6EBdfH02tUTl4SfB1xv9j15M2B/0y14YZ4oA7q
9o4KsWeMvL3foXX/7cEVsueQIFoXQDTCO1VWbmVaqKgHYNjgGatCXp1LOaEr
GZJexG0ZrHgA+wa/+KpFYWEMKFAV7UobxoczqOrDouHGOz+Bal3/Vx9pRYbH
13sANxmIlJVrC1WLUyItTg7XxQ6e38HMm2/YsvX3Lhvj6ZfEVgMdY6E6+lEr
FRfRz5KMhYnmAka1H7RISbVN0X7XuevDFDaG8Ks89tTPGMwSKAo2sSuBJrUJ
4Berq1AvYbYE81ssr1YNtjyB9otQJmMGO8EQB2yymVH+Xmhr31WY8mch5m3h
WIHkH27EckqyGsOabwq9Tv9RjzcQMP7TpnNL0sV/SmDy+h6NPq5iYnV+hUQM
xA1P806irXRrYnE++TSBDjORYtjgOmh4TnC2cpiJOR0X/uXJATjfT1bsFCob
m0uOuyLG3UB5aiyyk26MJ6Cprd1viz7qu7UvZA0+n2cm5V7/mfd6bhdzSfjh
Ceq7RqJTJf6mrrm7uDx9TZjwVXyWu3PzhsdSnjtnS9PxOxhdeGM7+awPuVt+
uxFtM8CmjLtDzmsHlhQg0kP8cad0s91JxXs4Uw3XlUEraztO1q7zkTDRQh0E
9SxJGMzcTMz7tXJ2IrF3vZP3haCRKz2KVYPhoxYUxIDIzZ0vDegLlnJdu5t9
E/LVYKgoowb2aWGD5rl3zmspY1V7j7yC3asJuvdD+yCO2Lttx/k7yUZ697A6
1AQB0s6E52bUWsU13pu6tMSBgY8TTqwtqzn/crEvC3bS/4mfKQB8YYA7XK/2
qS++/vOrFUvap0yfZfaMsWhQaxc5rkU7rjnMwRXI2k8zh8ru1UvGDpcFZwmL
iKcRXo3HaDks2dWJDMzK4BPFmB6z5+ozN6G3zMcpFH5QSYxX4M6FdSA6U6js
r2uZPjKXs9BkTYynj3/HXo68EbnR3mJRp3dnl3ndFFjh7tHVDSXTYg7Iv9OK
7RYu5Q2g3olvsWGVvg88fEJKZ7S8Z8qSbSmgFEwkkkYaTFVdDdqvyZt5HIUl
bdZk/gRK0rrCjtZmIW9RwfUSXEUSE9rNkrq1S6XIlUTNkrm+PDwuIapdDRng
oWvhXHNTl7M+Z5xrnDvScQQvQd5Ucp7oNa0GDECz3sZCD5cBjOe1tQloNTw1
Y/tdsHXZIfeKFYMBowxz05eKjrx7NwERzZfwpv2jm2cqsOr7SqPDDKNESt+H
Nmd51MsnaWbWjcjaSep59dnxE9sVwd8D/8PL4vkXbdAC3poR6UMFaitgeHLd
EaI0DJNqICE/6M+uwcKFBjSIH0klv7iTjv0I84UOlmTPCNcQmy3Sq2OmUarR
ruVZoUbw+BOobdnhT9Q0ZQD0ddw+sKF5OUikkEFk6Dd5L76DaIlM6zniH8MI
9fq+7WwaRAoLvubBwFsSg5/EZ5klXf9o/rciCOovLrGXcnMD4yttjtyr0HEw
jkZc2gVrG/S/LzU+YndFpbzO0b6gqRKr5rm5sc7sKpBeuNPXyheSYEGIxUJN
2gPNaULsxtgCN/WrX+4Q3giOu4iQieOUctpPvNRyfCP0C2VzdXGuizVFjwHW
KDrTHK4Z1hcXnrYuI5hE4QRzxeuI1AVHkbQsZuwOIMj5slgjpO4jwX0h66DU
fZgdx06gy16+2fOozccCUw/jdYmoHVb8StDQmswFOnp9FTvSyA9KUwIceEk1
dm5jtZyehJZJWw2zjvLg7a2429vsqVfGoDQiyPEmelS0n1fK41y41xgsE07z
/VSq9sT3LBk5xd5zB/hJ6/6/KAyHSWQU6dkNjls6zrRKPHs+MRRkNRPPccwO
5ixvpvTrVJ7JzYLg2lI+WOz78/oEKBg9Bn05sx8TnIGzSfL6BSws1d4TxpBT
aSFJ/T+ibMFQ1/a5VQ6axWry3M4jX2SUW3skztKwBOrW5Vp5CvsmZ47aZoo3
U0CTDY7rFmzfYjdqqnD67fpAGXZ6E0hUaPsy07+Edngfkr5B0PW95R22bCNr
aLPnOTeOVj+1622Dt+QskieU/6Sqk2sx9Sruq8WpT7yBJHkGUsKQEctZgokl
OxlVpekOGnivGr9iJUrWDLJ1vX3Culym+Y4F7q7fDhuwkFTu3DM9qaj7e59/
rTThijCWAMGPbSvNIXO5Md1umymNvO8GOJCMGcG0Q3zR/pgtYLZEK4/Xb0uj
sMdGZZxLHqN280OVinyDAQwAIaZMvLa3SmkM3L1olM9L3iAhluDncmBcFEcV
8v46IhT15BrbNEOeUb+vnezzgfjGpevK40m9tbJglwUK3JPLFTo7S9BfKsEX
nsGlQKNrwTZKLha70S6oY836+xndmL6PBX+1o1d43RDPeygn1Vkl7mMlRYHh
TQ6JvDbbokoa1/q6euo2ksKA16otSrOV+EGQCfvDqvR8wHA5BsCtau5VSiz5
gBUwssHXgbKoNyVz/XO0x+R9VKG5spFWofedymZYhFCIvZUk7Hr8J8mijhLV
ISLm9O+Ypuu0HQBjUT9yCqfIhh8zpj3N0CYkjNGkRAbJQy2mHlGhewG3FUW+
00b2eFzDGIYvfe40ipfbbkecokVxsvkMJmH8nvg9VcQY8bMq8oemMa+IM6N7
UL/lqtHO/ROJHeW0vgXsGhDdixs/zAXUWOq4h2yJo92ueHn83sOnmVifGaCb
NtfVybplGH3cCAR9mMhmEI3vUcxhyItDZ7g72XlFpai0HHQwQ9NrE42gx1RH
lPWgwzWCg3tWk2aQB3sWYzXjv/R9YoWwaC4+uQFsZUsjXnM+k7nk1m1Zk/zv
TdpTd8YcsOWl7k15YWUtQukHxP5RzBid6Wuq54x0ZDYiZ95ixj6DEKHrl2zW
/u5SN0eY1upkIfC4YsPEGGLWBUOrxUxgV7EmS75TNO8VcgJu7J1omR+4Qd8f
3Lh7vW5hXsrIgBlA/QcZUxst/qpZiSfiOvLyFj5Iwno3+0bk2M/muUXteT29
lE4GySeDK2XwhSjgei7d2FlcsIrH0LW0mebIoQgA3VNWrImqR/rEnwL+fmZA
CvfT1r6bCiByfFchvFx4kAz2nbBxk130V6jZCZ/51lFz32YmLQ0zyuTQ8rNh
eeVe9uy4mqxPV9xogvlHuP9mqh59WHmvlLz9xrJW1swCYxkcATwmPyvLlyBD
WjhHZQqNsO0OOW9/QkYv3Hh+bcnjJeC+EC5lD+EWPs7ts+O/fLbNWIXWbF9l
JW9OybwBnuw/kymrraA8B8S/88SG6zpYQKhIPM2gRk9xFdfEDxkYQw6Fw1nw
50PRaWFrGk26ogOCR8prUNDXwwPqC8ELjVVczswMWCAIMEI5U0nEbZ1ziCEe
oqgzExgRLepIa7sqTrvG05eiZQoKFNl+W5NcVrQhh6EUvjRIFCt5vFNc8R2S
0hX148LWdGHHq5GWkbC40IetSQQ3ld0fweeCVvQ3/KffCqLzeNXdObzJORqX
xcNfv0wNiGkL5GOMPv/zLbjm5KjGP0oH/khym5efX2zNBfKNxn960RtFLdBj
5PLr7pITh7PKuNChthA5a8uTLVWjL3x3bGEYtsymZc0Bk5IeX7cHOhkX05m2
d+pFBkLLQ66BYxABD+KXbKyX+oAjnnUrVrEEujN7heyKcIdZOcNpx3w03sC9
Ytqt8vgYEEo7cLQ7dND+TU0MOT+z7uOQpPASxO+sARo9hlapPlLxuE4nA3BW
TsZnrhXDPx5pAwDwughtCyhpu3DUfUtRqhcAgzHK37DB236ZVwGUwEHTWTjc
5mRZbbQsJfhNoniimF15gxEjlAhEc5KoQGLfA0ykxDsyyVU4f99UbqebCDsf
I2s8EAA0+1VvqYLoEaNxl9UOtoOLPE/gtJVP4NSc4sOHo8uFHGz2m3gRENrm
xD63K4nmT5lnwPeDVcWX/N3R78SaM5nA4Qp6TQ3TCjpgjRIuxKiU9PpYccrf
VNVTDcMQnVwgg7sgQtZia5hwDbzoCxAVirrxGdhuG9VmGxvp2xrMFLmeNaJc
AsU/lz/ZIUVIhnaSPaayYlOhm8SdCLts1rGXOLhpD6SwjbO05WOFefTiNo72
JvggsKSi5OAY30JnDwU2yLzt7KQkq1B6pCi/f8idC5609Gw+vFoHuzGK33FU
OpeuEpMN09Bc6rxuJobJbxPdh2FLmQQMNfCKs2G9NlcgkE4FLHiT2WSJIscN
/vt8evgibSb0/6mPiiVpdja1qWiS2Pp/z3pu0/CPpVViOirizxpGuS0OQe3z
ghf1eRbYxD8Zuiy/han2RYMNRIJzIpRdFhqin4domQft/wCxE7GNgz+13jJW
fUjWDBnO5fQGPHwYZUhkeg2bBnqrqOEjLKROANZo0qk1O6+8oUSGcAQBcbRZ
bHEYhMKC2PeHeIob5PJfkL9lYzwGiJIn//qT/5avCfSybDWOH8Ei0NE93II2
lgMQjaXJSxr+xLvSNih+L1etjky6FK8upI41EpmfcxAe0kWlnBVLTxDUHttx
MGQT1hnSzmtC2k1w+DckBicL7/QLHj9Bcn6UTIEuMDj4MiSGSGwGvrkmJ3LA
Qg/p7czaqzFaZfdD1Ip5R8xD7m1hAlFHhIgNnlDuweWOWddIxRea0rsstHLI
sBc+LaT4UtiLy9x4FD82PqXEvcz33NsYFtpLWPQyYqONMhyxN0FzKFUJOsEt
w0/oyyMxiYHevmqyAsUTh1wSOEUfnnwh7ZPdsZ5MOUdHERoKgX8+07g1qU7d
qebM3V3loIhkfsCW5/o4H8DVbk+xzUINHaPn05h7O2rDwOqWkdPKLS3SW8Ji
EMEQZ6Q0eFVqyBoT+T8TVQNFzpQGvesE86NFcf1ANvPwWtDWoJlVwXvZsjJ4
RwTcZlGlfDoMNCJwplW7TlDLJTDJUO+plpFpxY3X8ouI99bEMy+i1qaRGjO6
HXG89/T4eQH0CSqJsM6Fy8vZucQaMXoCT5KfvYp/x+PNrCZg7JfM01GUlyaq
mPAV/bQ6cCxxjPf/HcvrPUzvXX1nlTuxyhbdR5nVFforslzu/rPYxsU56PRa
EPqX/zpbS8OdJ2jsDSgcDXjqbyColB6tbuOkkWE/hIALPDUIojh1fjQ9W7oH
tEK6T6RUGZHGWWwwGLkUhJpqpse0iWHCiipmjpsi6BDmdwD2Fn/Z6np7zSf+
9F54miB2gJgPmq1i4lmwHh9JOTFzgEFWSX6Hn7MG1C5cP51vB2WaogtU4Fj1
9OfncBz6NqZ4v/qi/nrEFHiNRmMiIODpOvKR6Hlg1iER+UjP2alwx7sppFxQ
/dTHg+ydFVe8KkE0WUA0T/SgeKAdOE2LDBSCqTNWqsDsnlZ5lD3HCzYCu/IP
/5yaUh7lxWW/MZHDQPJaI3K/AAQQW29kcnAXL/3nN6/VEK+cJ06gstEJYD3r
/fgdAXJ8CPBmqQbU1i0Ke8Vkz+rZJ1VpFnDPq97zG/nXdOinwmMqA9lEa5Mv
PF/tcQ1W1Jb/wdEj1xSUwdd04LM3U+VCWkrQ6/0Qf5Kl0799b1o6oNHtA07M
NG11bJZx4ng4C44lwG3haEc+E7WiG6AGFIf6fMeyZ2fwWKGa3WtpUuAXpCGI
BDNpdOOEXxKu9U8bNknGOwYJrVA1kV0vl66zHYQCqk8V6Qx7rW9ZXGZknr5z
GbPi85QTALejXgg4Zt5C9UMa+KE1IKZSndTK+N15ZeNmS8p6iGceprMll0Z0
rqiDAOS4K+e1oKFGze0bQ9KjMWPNJ/3geOTBQAkQ0oo38DoJEjDVlD/E1gAb
qLvRpEr010Q2ibkodugD6ok+d//orz9OrD38Db4BKGtOqCD8Xmv901ddB6aU
8zeHWVVIhfoXk3UHtyDDBDkQWsQf0CazfmIX4QdmwV31OFcIZPPxrhAfigFv
fIdD14y7wL7Sbf1gLdUx4tZiYrFIqjQy0gPWPSF/eMwP6N+HEugB6lhfSM6f
/jGyg5bFdZF7RYv2Aii356ldP/MhOv4ww1kzWFiuXRVgjZxFEcb7rxaglRfS
xcRv9WTGH5uU5fhpNHudt+qfM8TG+KvNJXf7IcC3STXaeb88xkyT1JmRFAKT
vtzw+Rri5wMUDyxLLEsRgOr3AedB9OqB+qxZ9u8pPGY78DcXJv6+6RMSsCAO
0CP4UvOMMHICqgm731LdYSM85kL8S9AD72jdGB5vqKHnzYcMGAbxqMzjQqWE
94tEAlt7yyBcFmQu677Z6CeuyIpPxdQG5oan3ZY0clqNW19Q1sgwMbUlRgi7
y+zGtR+lL5wg8PY6jx1KallUV8rDEVO8uzg6hdi5DYeXVhwUSbL8itcRpKAZ
ZweQj59gF+w2uYQRF30Qz6PN8XbqeF+zNryvRUJUSS23XWEOi8PEUGAlRrdj
qKmCpuReLuQcHMrMMs7mxCmHRvr7zM8JV0mcAOPbFqIa5ys9gDPKGyOicHpz
A9SMnP0vksSv6bzFlQthGbGCB9TCBCZIGJUXgbnB3DgKDZInLX6ER6cg1BWU
cGuXQ6BmqVSG8jarS3+zYQSWYc/TTKtpW6x+JfdB8mWZUX9aACQ8uGn0f2Sd
o7Wtq469MGUJiqbsAmTiAvcpumVZYQQ2MsEWq9D1nSl7sR6eYm2W52XyYL+C
phLAIcz8EhM79T1qAfPF2CKV+Q4kzDctGgO5wcAv6mWGrCNLdx+GQ6SZW3k+
503o4VyTgUZAmwnifp0zBCRNpLtLnJGh6cuDTEUsiceqtwBKOMIWm346mYLn
vd99FAZkpfkyJQUcBPUHO1g3AD0uVjcrGmWNj8yWlyEWFmm3/AGNbRQho/Cl
iqL78DlZB29a+Up71TOK2p0Nx4vpc6T8w5fiZ50kdOboi3vaB+8B9om1+Azq
ovWUgSleDmC56LU4U+EPaobes4tsUGgM4mfIR/K/qoOyfnn2aokSzlp8kaZX
+0ZvRO0V43kkxxfObyReyX0+GtU5NW/eCx+NKHP5pUlLn3PVpgqKe1fWH47L
5512XnBBOIW/3G3uMjACKEeUJyJzKm1IfovoOTbj4Q1aXrsoIngH+M3N8Mxb
SJldZf/4crDVg8W7fxQcpRWrYbwFVFsjGbYwflUaBRjFNhAUy85WsrXieBC3
RWH3MzsNlc9rrZ4aAoQYG9o5z1E0NqPxIqxJ5+x5dvAypmuPzcPFT6eVa8k6
CRC4fWnwrP43Bcp5T+uKoICHIJz7iIpK5JrmsqzT+MeP4I9kjsbK6inbwO3h
397qb3lo+yEeJJvR6jNHasIcQOWKynxvU+2rgTEEGJ8VXZIoEklszFSmXA8y
fe5+uoq+rIDEzy2kL7k1k+qYLuN6bNPlnRYP16Q/WcnAZ94v1uQP6auPdmK/
6Zijqgp7IpzJjoPcY8RQzF6nGHrP9YnurMrEl2khOJUMpPCBxg/CwKoGWsh8
Zhm/CCy/chyHRQKy4yC6jTXSZVcpXclOqM3Q+zSVv6d9V8GiHr9yfgSdJtx6
IadpLFkrWCzWtXqVZRdxZ3qJl4PvwrcFy/evqOkba21nTYrYwOYXs9DxAeme
Nmzar8OCy9+oL91OJxzi10D4wGz1NZKw/BWV2Zbh3wW70rSMCT7aC1kESpMQ
L4tzYR0KNUVM8t2pPBwdOq/d/69I1RfkaXVaohzgqkUbsGPxq0rSoS4Fremp
SCkFZnjV/g+t1BWdc/r210gM3TA3d2tOreeR3E65ocK0qzHD3NYMnuR2BAUl
V5tfnF94RdXcnO+BDrF14zCLfnHxIkoZdwEEG+WINtzV4Av1C6Dz/k6G+QSH
V+shc0kG3NHuiZYoJJ0i7ZzfAZtFkz5MSeqeK6dmnvI6/R+FVQ+Ta3wheKtJ
vLJnnVwVhgDjqz5SdPyfJAleeG2tNVetvrw7PLX1zMA2ttSD0ImkrKi9HWb3
b4PoWdhjodJ4lwYI2MDn9VklqkXq8EaR6OunRLGkEpEiMo6Ok4fda8HdTcP0
zRaYCUR1BHoQct2Fkv3wRmaEDIfPbqxKPaN+wca9AompxL9hOUHHnyIuTcDP
E16C9v7C0GliGFps/hbmnbQ7zOy/mA5MPVBMPzWN9tHbVIX4GnE+Ddl99okp
a62eEiQJu9F+7yDdKpmBFly33efY8aumcgLVvXcEl9APo4Spv86wlnEBjrRP
WoYZTSIDJuJk/RICgDi5P5VmHCIVPkHqw2XVK14RZhiLCJFFJmM9fFlEi64l
cxlXb0HBAyNmR1Qdqi/pKpFFIe76ZBz//CAlkt7W48bStcWRjVdsRddLkxVi
JjclkP0FiSazD8n+sDCkW12XKJI+w6vzDHwJ4zo2K5Y/Fzm4txpjyMB0Dj3B
MyDeteAt/0BbSuT6MOFrXUH1LxrL3JXy9UkPV1CpxXjaQ9FSaM+FrQgLuLGW
xDrcfyZs66h5Gb2TwpTCAyYlNdF1lQnGRz8R7Lkk2oYJuJ0+hOTfztDnWTq/
k9YTKpjzd/DUtptNDe6IiQt8/IiFF0aKBIERLUjlnEErr7mWgqpuJPWLNVhL
JjKhSUvZ5iFTJ4caLw6Vnn5amssYMuPknqwwrGVqXT7J7wYyH3eX+baTLHJV
wZH0cZZOLauM5y2RhVmHS0SxfLyD3Hvjwzvw1yXiEk1LI5ULYwvqbTc5ltx+
nG1mxuHW6d7dw+W8rB8qcGFuBMs8bUxe64YNIo2w3ByDbc3EvTNf/t7p/MLK
kh8XR2FNeLQjUJYZjdS9Bkp6SnsdHxYUqa8zqYh637HOTlPVbq+2Cp6C2JR2
XoKyDoM0uUSd4ktTbvxjlCF/RUQPp9j0w8KRSm19ChUFe99eG1PS2orEnZdN
If3U81drTpckZtI/daH9auA6I3Q0N7HLUpShEUgUcVrS7Nx0CBoMO1PwJDrO
d/1zZwnWXUabjqQSNVeF50uYZeBxSLJPYUmr+v7tjUr2z7TYPLrmqj+kB+m8
g8LoFASHx3kJhbtYmgFhbYOnzWxwu1qqEavgosOBQ0CTE6zY4N9CM0SlDnzc
k0M1K2YV8Hg71u5SdmCJuYx/WEICfDvj3kMICsDEqg2ai3lyw5/z+9X+JDOb
c5i9xHRqgaEb8K96BBxhjt89a8E61wJySBJfa4SP0tTnzqYFc4NOiTX36wT9
8gkHGJRA3dRyqT3r2Qmf8f2W0eRrcDR2GEDDpdmiNhmXxS4JdyhnXQzvU5BI
7GpHyp+DTbjZDtn20XCWJc23LwqDWEsS5IB/Y1bgi0GUDjdiBV7y3k6ZBHB7
AYIz/BJYCSd42BJCKUWSrWFAaSL5T4kjlnY74M2i2uKOV9SzWoPV2A/rE7XH
O3hBQbR6Al4XoX4ifQhHcFGH/R2MQTrss2UcYE43vsjTyjRxcq8ujxcj/rPg
YGTpAZiUj2x+wtT/WHYCUmOo+IwPDo2uLfeRHDVtgLdGMDXSLvbZB8aY+tt+
xHZ8Y4eUkQgxVPIq3btB5IJpJrL6snkvLh2Desqk2bq/XsQXH9Fwtw9f6DSG
SU7mK52RBZNv/vtnQwzR9rHuolQ9fSgIjz4YhT6xSOKl9+LG+V1Scn2bbOqx
ZMDxuoT+Sy//utQADjtYtqLoCd4RXi/nt5sPpzj6SqneXl80t8WxSh+Cx3we
C7BsPrECtqjjQbwhH2CPTrSk+yO3rSMFSRno0xz2T90dNan/yvaK0tLBr1vM
OFE5UZa1/47zQJTAY1irBosfIwH9o8guJqAlS4G8EN+nq26aZY8PPajJfd3A
OkxK4emkUhFFwIkLv7tpc/aFZ9Y6PDnpamXEYVlIHWUy4a0tF3dqlSgDhQ4e
PiEIG+7uKhcJOziFITqWYtr78utPy2d1kj6B4IlcIDlRxGDiPLGFqnkUDZv4
QTicWw/eNQ5B+rmszvUetgFav9d1Wp4cMt4cFiyFLfPt3qVIDi8XaRNqfqZ9
CLWjuXYSrZX7r7kjrZCbvY/vcVYWxIObXyvlhPtzevSPRybqfz+SbSmPs7Lw
5OcveVVHai26SV+F7cwgoFgdGUZx4Dugfy7UbxF1JJRKH/CmyhVje7W4Unqn
M9eHSK2hqBjojD8K+1ni9UOCbnxuhMYAMyBG459UMFXT1ZCKSXBuflK5POu9
/90FB0nwtiGfe7zMk2YAADNYfo2Z7qw0bk+pIttJVoR/n3KTpMSmL71xuNw2
M/hwJCWN1sNg5eqVKgnbYMco6fj1yhv/UErYoTLePfCyjHni21XmPQaB4Pgf
XYe1gnRZJz/kh24GG+Suj5OQYsHkxAzfoLsg49hcPKzkQmeJABLsT1hJ4iFV
TTWAkGM7xenqN7iKLupjSDajJ81msKV39FDwYKbpb4vyRV7XTnTLPn77Vxg2
rNuu7wKBfXdStVhw3YjQEkKVSaqdk4aFWwC9PiljFPg+8GuzIM2AQDN745sY
mvaaLzELJy5Ccw58ArDjX+uVvkeBlPwU6+jtr74JtycedrY5U3I5js8CBaz8
GnkqoNNfqfG6Op0zhMImhMevJF6bTRaR0fsfnsIA7tWAorLIyV+LRNToBpbg
/NPJVk6mxdWTIglKa/VEQ9tNbYmnzmz2hbXTP/4mQk0bYrC7e2j6yNaFRVRs
+CP/K4hrkTFKdpeXBg7bSvZjBqIOq+c+DjHVieNfUrzt+FnMu58wuYwLpOVG
3Z0A/FuJjmMfUQzswgFknhgM7lC2CfqzEZQTE95FSOxuxMWJGU1vpG9Cgwu9
dlfZvdn+yhexenQmZt6pIVsK2o1NwbRqFtnIIuEz3CsBsSLziEKdQf+MphDa
xHA4Pd2xGYsNiDZB99sc6HTrDVhugdby3HV0rmjchJdvoAumUSh5GjoA5zuB
nueVRIOtUfcZg53UGkeWVC7SBaXV7/nEAMSZh1m0st/xJshEJcRDuq+u6XIE
NktZVVSf/6hSB/9nSPBkFFrA1dngl6HmXAOXx7sRZO9bHXVzurWpTPAX9DOZ
50BAtyowulyYXewCa4ilZ4t2AQOsgiLBWuCwgc215E26543rIdne9vYM02gJ
0gkU9pOQFJoHtxEbUOeL/oBWPvJ6TRdj50DCxPgxTm0+2gITCqXOoWQcPCTW
H5i+4r/72YmOzqg9QH8VUH+aiCBw9O7HpLM6y8MuF+0WupcUFHHTpYIniYAm
YRoc3HPe4NtJDGuwFC5uSSunXI9iS5p9lea5HLAZeERrBQN2gsPqywSrUw7M
piJ8J+PyG0FOToYJVpZxMlOTS9FX21YkKLmMinuh9A6HRLeYuxtgt/ppf6H1
0omutRyTFJpN/TTHqa0yotVz/2QtVaeLvO6s0QF5hOQPiYSow82YTxkWV8vY
JuzncZrZuc8taoT0Yvu2jPdPqOqMoXK8l2c18a1Dddcor+K6Uqt2KXqg7hBt
3CrpmP5Cx7S7M52mDPVVMWy6z8rsVhRzJNuKrBUgoYst5ak/FZWUSgKvbNrd
zsZwbx8QBj1j0W2Qq0Y+i0r0WLLyyZ5pzWsJKRlncmtNyP1O8IOAlasaxeD+
a8XZfRJIOLZ0FFGznghGaIZ84kB5o+uAOp66EnVtIOGz6VIgCkwy1rKs3pzp
ZQigz5wviJfBtPtCFBbzUihb/b9HH/gC2GhDuuq8GfFyFUafB2pmv2JX2Oub
64mpvu9r82NxI7wb/xOCwPZz1+2ccJHw+eOYhyiwYz4XMGZQ21c3bHNkGSXl
KEBc8RTO2VXsTiXxz4XeLcWn1QedyzOL7YNE7sMMlYCnV8AAOjj1lniIP+iB
X0S0orF2AIqAReeRUpzAVI9iVEe+glVH/BJ9Y4CphV/WfkUKUMcBRNsFos/5
VqAlEqKoJactbRftE04zzKWQzDGiec1hObnCVcKz3RQxypXvwxG9sioBm+pD
a028Rrmbky11Y2NBoka/tewAbSMS7oENaRKqImZdv+7BRJpTsrR3vwlIZpbi
XIRu/OcPiPRaPp88K3alsSh7sVXSqNBpz96t/dAeUhxx7uzqOX9hHa3LBBKe
1dKSwGFl0Ae3xjTXFIA3iV4HwoM3iW3iL3Uq6hXFJnPFhhAeq4iUamFB21Aw
dOUIzFtfmo6r9vyH2om20Kc3G0QUaiXM54ghBW0MXGa58U/SPUahKAZDcQjr
rcFrkFcK9RblmJxQ8lDpKM5x6fa2UVgY5zAH2qUEoPOBuZ7KX/EhUOXZyQmT
kavDIToRGjPn7VbNY1G8arr4MwqgTw+Na8wC1B4DjKT1s8Ea58WCWxjaDeNs
ZqNMS/QG5CCNf/6WrQmedUX5j1ZrQk6db33fYFL9cxytYlk50c6yCPl7fLtN
qTuxP1i2Iplgewk3DJJ9eNNSW4lsO9yzqMOi6DkpwGp/j4VxmRehDn9i4X8H
/s6MF8hSSeHeNAlMAGw2ZgsKj7s8hRsq3e94WKNvr5/4MhWhCZSiBB86dmzY
YmoEceb5uN6tjPKn7loFgP9QfE6dXfbxBFmWkofKtWa3/hYqwcW9DDPKFGfe
f0ruL+EMzY/fiayoYrqjTWdFNZRLuabjgzckiKrBhrFdfU4qzm+AIWnZ+n2m
L197EeCV3micVXcfVgX5GxUR8WG3mt3mqOIyY5BcjhjCefQEpZlfRJvzsYba
ArICl43aYASS+O0/D4ddalQqdDp1ZpBRoNWY3JkaS8SJfyD8UgOVhUWPDEHh
UVDyHGskLGpKoRTr79kh4CIJPt3eqfVzfNFdMLelxUXnp3c6rC0MupMoQCxX
hekwiOARRUm3CMOujeAeeCCvLck3sW7Vq8XECyGDXsGge0foAyuGsz4NF+bI
AsIpvnuWxyeK9Kln6387uXbVR5pvOPxozq76Ppgc/Qqqoqt2PMqtGvZL1lUN
0CEioErC5kgN3/blGfEnHtQsqHk/RuwHo/b9N9wlSIVx3SQM9rgO8dUhC3cR
aSVMbtv9oS0fRNDyr5y0ns3Hn30/td7dhmLJyP+u73PesyA+1UTSuMU0m0Q+
G6QJXcNcvZLatEJkRMDx1HcjxDRHoyJrOOVNSL6jbttEfvGeTCC7uGKCTPQ2
ewU6u8O0kvjmZPNKDbsO5M6N/L/snpbX0l/H4xXFpi0Wodll4Kjye1arPrgM
8JVzB+jeW03+nODubI2Z68IRooLIOi0A27noSRuGPIkBRAMtqkTTk1fKfiwL
Cbq5KxJ+KsIX2LLUv45/JL/Bhy3SJmqdSfVRFHIog2zaS3UuRD3ojSZh2ghG
S2Zbb98cZP0r+00bDfwJk0eNRCP4RcXQ2jWOXA1owJ5x6L3b29IjelNpzHH8
JeqEO+vQYBhG6yXTOHCTVbLMRhq/Edl9JUKakm5JiuUNY06F21/NP7t3HFgd
Mrb9SdZ1e0pFfuEV13hjYx1pk9Z0wxpOk7fl9/W2WXmGNAHme3j3Z3hvRj1Q
nTHANsP3CCat3a0OPTPKV6Wx7sWodeV6sbdzQ+K3j38WY5rrFZaG51X5aN4P
2tHrdkRJTdgK2OCE8b3HHhCZ+gkv69IAfYO9YL6YIpK+NyLUFxBUk3w2hhrm
VybmkewYBD/cTjgzrk/Czy5qujM9eWbj9nioVhxSrRAHNTeSzrDUOTkuQ9lX
cDHBACA4ZC6efja1L/GMUh1pmSioFboPzqHvK2q+X8yAywUh1AeWc7dLD1JP
/rj4CQBR/VfjVfyp6hrvL6ScB7HaO1unpD7aHcECbkPvbenj8AwKQObcqam3
8BQY0sc4fq6PJxIZzzkxg6/P3qqBoj1Gx3ehFUKNk+uZUcG8kePRRGWNwxdN
fLZMsS6mmyfuVc4J73qigRL+1txbYHg0STjAffK67FYCGv6DVznDKI0W28ZA
tQ6LZ99XJzICpffX+oZkm0fxrbFXD9b0bXE2AkU+SGSA1aA2Wn7Cei8+WHyh
ov9AN1LuB6PzNlQnCcg6Hn3gHSNmTwXP+QtH3FxwVIVqWruqoJ/Z06fd1kga
cbVP7jFpUj/sxhFLRLI0TtH/Emk38mtEtda1mkKnfu2k0XL7cKMaJIccZ3p7
hKaPSUArx+XdOeT/v6mvcWDUu5/MKYgI6dom6qm2v0kqKkeAk5eJUp3ZMiEq
2bIghqnutEP2ymLp+kIRJgVI3ndld5Iv75wOZEe2KUK3s1D6Ma23L48TlE1p
SPkanlqGu8C6jyVNAOuu1PrrNc1XTSvwYZMOjf7Wv+jK5dZbqiujyAyCgFPM
hsUzSWZCsKroCGLrd8LAtHsKOxGPbw2NnzV5NjB/p9aA0HFLhChit7qk8IKr
SM/OCdiTTK2eMKIrPrItRCCFI4nIpQy4uF1ckl/+AWxQkA/ZanOXMOEeSxoe
hhKSZe/uU4H+hJNlpxEhhbPUaQ8xufbv+lbghBjltczKv87J3gkjHXogV41l
ZP6sHkuVef9RgD2Wd78PTeS6I4K6BZRsikXB9gMlOn3vhaJ/dngd16txjK/q
SvFPfRoAvZdoi8XrU1q+6MifdHE4lP5W6Be5GVyRcnTofN+zgIyYSjofHj6M
Nr7A1asGi9sI3dC2qHaUx4szlUS63uP0RSDgitbvOpe3+TUVi3Th9UqFv8lo
xOo9uC4BDeQhUKFbfDYYiVf9k2T7e70XZo3op/9HnhgUIHZG0fiHFZDD0ET8
srwXvjYNS4W9pXA9TKxbPobLWH2K4ola1Bn5nFiihfV6/NfS7R3dgpnpxs1h
p1gK3CrjK4zkGBZkHcFQezxF3HhEzYzeDF2bgokPMgnUDqMjLdZi80zOSUTN
/hVeQnyurIXczY+7aRQ789rN5MGvKdS6YNKTF6hjljOBCN6Q7I3dTlZ3ROjS
eAxBpGQzB9QzI1K50j5U9o3yi/ky3ZMEMhWCrIxFMUagoqe6lNTI7YSCBpdc
OGD4rlZSxVSeNV8XQ9S6i8dO2PcrUgPlRRdwg3hQVLwXF0Ovg310OJUeF4HY
wTRA+DTZA388CLglZyELcm+P/t4K7NT29FqeycLP/IPOhk8518hMc78le7Q9
3daELatL7ky5Nduk7E8iKMBfa9G2lOEwhE8BfgiYxCLzK92IzeTSdWQ6gouE
fqGKxeW4s/Z/p4Hd3KVGe1OdPDRkIo+mubCd7/RpqGenWK0pC97sheEJVw2S
4QslQaxMMvHXfnLWCwG2gK0wPSL5F7vv7guwzvJdICMeJe/nhG7B2da4teGA
AXDpvnnh1eYhdGYXrj/lENcQnyQzDsdLz77H4bx1zfGMPt4W6v9dqeDZoNWF
t0zQ/TsEdhlUxLwPMcYaS3xM6eikH/s/A0CHCnMPrn2LzlIk6o4Dl6N65L/n
w++X4Z/NwFptZolPAvp96nK1/JDLB3/e3AdMGmDIHLJzc6MuF3p33blaiqdt
HXWmyk2PM4W+tUIVEpv6j63rP/YsgEPtKG+AYsWGpOHvYBIPhy66on4UhEdo
0s5t3ArzcfoBZ2nqUDVyjyZ+huvKFYrGPfMnFtyrxm8ImiHw8YbQcb/fMoEB
45MQMIdInzep4nRBC3wuytP6SznvzCLWzJO6ieUafNADZ9x9M6UjE4utrj8y
tTqKLPdW4IMI88guOlBHYjRnSIs3QSCyM1GKpci00aYN2i9UCmCvdcItfKWS
NRC92BcJ0kfMxiB/2tQOCdNxcje0bQ3xkOSXDilQHWoWZuJPiIm4ngC93c0G
2FjED4RTXSw3Jyomk0nazNgKEYJONuTCt9bkkPOPWTPbpSi7A1Vdeni2Fddp
euT/OkOQwXHub1Ow1TZNMrjTxUCTUOSE72whhFJjQ9FH9W+Amijwg/io3eVw
1Uu6gl7ZvRNB1iOLZDFwjUmxxxAoJbeLU5KRYSPM/RvyMFMt0nn6LSKJvXUS
4FZL13fNKcMWv/lYTRLQEXCXcoGEsCp+83nELhS4qyxqodpE/0BtGFG9ZoTa
ouv61bdJIsjOdkr4C83GelMyYxnJZsXujPh6UWQ0bC5TIKifSsIi+UDv3cYB
9otxysHdbE7aPfDKntELLS7QAOjNc2r94Jwp1RB1VlwaO00/jb1sVRFCO8z8
9tKGlPsYsi9NRcdyAJLWpdiVfVarB88fLERQfnCLqpH9iV1J9AJIXZCxPFuc
CajamYUFKviT+2WpVypvSzVFawkf/OvIJjiuqGh50H8eHiy3co1YNO5lzpVO
P6meAzOCEgHl5CpoJ1FUtY4CalaBIuKdaDi6XnmSQcFfROXxKJuIpb+Frecy
yDdpp8BhrW2Ce+YAa1EGd6HbVxy6n3QMc6LNBRx1RMdwHd9l73kBQc0rgl7+
LzFInVhAKQ68YqPPKZsdOcP8JVTjPEZa2zkkDY4w/xi2IDm/+RNT0eOOGt1i
gvFtEyis+tfGQnBpvpTpuJiStbRQbBVrqbb5U18V6faae1dIZrNhvasK05ia
HM1L6GHxB+pZM1gcdLMYeQ4CmI5vJvi5zc43k78Vkc0QA8x9NJZTAK8IRimA
Wqk9lFdAPLlcWTcJBgm0CMguLtRARDUg9k56keBwzfzggalw+Ck4qNSvWPUj
Tf/PUiYfsDa0SLi1WjGg4CBm4L+IcOa4TNn3Eu6/1lHSBvMAcbtdWHj0Jkry
g+AEaH274yZoIJvQ2gjrAG1hAIHx5ofzaTIAqgMyyg0Q+6QH0fz5lx6A74Ow
D/p8OFOuLSFPY2yBclIf4DS0MwjgtLq/DWuD+F/eZWIekbOaq0nQUxkVgUkB
8AVrNjNr6JzEk1sOe1B9pWpfVCv85+BzVbrGgR9i8iAtMQT2lC7DCeUff/sO
kfJMVB4lUefRGRNW886ZWCJGsG8fgGcWFNARgR+MfA3kolGFox9EA2chNDcx
Oue4W014aef9uHbHM2bQ15w7dPjaC30Mhus4c9RPrTScDxQJl2k0afE/yBiX
23d/lYoJ8BNXhypQgsE1UyFLwUtuAy3I2QhJ0fv2Gi5Wt9cnIbm2xnEsrwLO
rUCf2YiWFd452fK29LapjLTWcjl0AwWeqos6wCV9MHJQqEd/1RWjOqinBxb3
VZJiZNDJkOrjmaend9Szo21LBxO2oS5OY4d8A0tDiM30pC0wBFpqOIc8l+PQ
+lPbFP/8IyzKysX/ldgarf7XDJLTb+OlDpgxnxzCDI47Eqwp2iO5/d4wlrBc
Mp9UXfruEflJNWGV6fkOLI+w28yz5PIQfqMsRBgnIeae/QU4utUPOBfS/Fmq
2qRRbtaVN19T5mUmk8enXLa0V7SEl1MbM2p7ksVRRuA2MtYpiq6VcxQsVNCU
l/DmIZsOz+Hc/QvGzdrjjwWBJOWbqD0eUZXyUqaKnatR3Bf325V/2CHTOth4
I2G8JJWMmtlulPg1EPhTs956VfszSzf71LU+D6NZQ/VwCAKe55F5LLVo8ytb
KVv6LfddH1lRK9CpK6887g2/6M8j7PMSV17NhvD0JWGcSXQSBcVB3xHNtcEX
26nF8v4W42QFiamtFvHThegxTR8bq1iPX3RkpFZQPOyvIr8+KdUr8iDAd2aZ
PHRvhybbl1yB627QPrt7YLDs1nE+08N925YkbkLs/awk85kiM4A+vG7UptP/
llU6ocPve2dL9BHk4ni38FSuRl+MMJAEm58+HJ1HV/39/s8WihJlxCDrkUhs
B0pR1xYby3HE/QpdH4vT0/jUc87ZXCp75DHUZu/1OZBvpzCNqrlXuOYssp1r
phT+g9FDIL2flilGFbgJ8z7KR+3W1L4w8udBfDRYdvLiLuqMjI6G+d00MYI+
QkpDL7jdZQ0fXbpkV0aqVxkiKSDkLXu+EVCDUM6BAfyJtJkcBNSoBDc2aEQn
48PrUhfFbTLloTwz62xbMDZfJ0rzcsn43J10k2ZE9Ike7LZTGF92gepz7mQb
ZYDjTClXrcLJrqIG9lXlJLTqXx4VMVkJ5Rz+j3CR4FSGdJ5piOZ4yH09ixJQ
SN/tVm3D/Onj5qziSTRm4eb7F73RNDOs3HJH9HI/puEZXEur/mlssDQD3KkQ
b4HRfTdKazMxkvTn6VGNyf3rrUTVE3psanqp/4Trxii4cJhMOQz/AayLa5FP
aj04tZzHQK4/G5iT9kCXrI6fagpAfcW+qpxsIgQalp7lKnpRp/ylmT79uU+t
MkDYdSh1xG4MXsog9zTdBVeqyjtsJURjfyryjx7VeEW1akaqa7TIMjEVZL7Y
kA27FmvZxBT7p9QduG8sr1+nHBCq2T9VQqiQmwI9Ll5wGqtiOkyd9OON3Hy4
6uhmkZR+4Vlse3bjMxFQtyL6ckWw6vL7ycLQ78fPAnAlrvwk5Uy7Bai6IsDS
JHrw2rY+0w6/jgSHhvFJCqZvO3AajW3t60xCjOm2raouUNEfZYnwDmbOhEU7
82jQ/XkGswshzawD0PLIkNIHwLlw2HfLUCCFT6NC5EgUgDEQs+nlCeieQ8Td
wi+mL7kDNr/kqMek1DmlLBso2khRKOoHxDjJmVC16w0EGMRgMxkutM0z0ZVZ
yruuKZAnqAJWdkzExL5tA+cuS/YoxBiOoW0mzIoycJqNmzjiXbJ6oA6w7HwF
ef5Grsx1Ihs1BmCAf//IIx3Z2qewcfKQYza1qeyDyS36FfL3oyvvZ5DJhW/2
elror76bDYswdKZ6RH0HXrFcgQ9tk8NB/BwuGw2vcyZohGS66/Ibo8KPvRQa
H91WHewKDi1PimudVBYzuD7RDecAowim19IM0wrSLaRWW7BwERYQcghbn48v
JSLHoUT45CyrJkWiL/DDLq5+UWuCB9vd5wqdygvYEDRlreTBgGiCprgQ3UrE
U7f1Ldk0aX47Lhc1BFStcnzHupyCkJWJ+tsFee3hb6RTEwDd/kBupgb6t2j8
Du4nD0OpnCB4lte/TxM6aTCTL97RUF18Z0CjdNss7uuhZw85SQx0QdiqDhEd
I/8nmFH7n8ZXMUiiEWCgbYituwHAUYWzwQ6x2GxA+fw/d7fFb9MgCC1KCNDZ
JqyKnV+SYO8QLgzm/8ZoLaStNJxts6CDLuBtDXj9RQfJEzanLnrAKpRlMrpW
xMxLfFiFpsmJjHaGAkk7FM7YFPBdRt6y2vbGgE1ZHYh6YKGOBiS51aOL/5yV
3skRXx4NJk99ogj/7zdrEh1f1iRq2oVv4MNALuGtFWeE+Qkkz2la+/qkNGy3
xIgTZHrtCU9lb4aeBWrg/s0XDRioQ/+W1bdR8TbkAUoUymrFSQSu/qy5XYt3
4idOb3qWS1zfElPtM0tklcm+zdxe2qgtEWY5z+9SzvDHXPhkgx0hi/W5xGex
aWzvaoVqki/DtiltSRpeEi/3Z6Bcy+4LHOxMaSWTuFsUjtB1NNqdE1oS6Ygr
0UeWJyD/6sAGdtlrGVzpnxeEnT8ClGBS2BLjiKZbnGUR0tLVvDaiSmpsNkh7
lH6/KUuiLtp1czUn1c5szHsx+vkddgBgJ1Am+Y9G5+S5azBfKCuh1fOCAmhz
klGU9TymuWOMVk5lHpmYf9kFkQTnYDsC9HZa9raRa9uJlwmE/5ywbNqvLa69
RVxNhJhbdHGplvuGgACoOU6/6dRiG8cxunksUvEScm+Pqk5EGg7cMtTMTcem
n7H596/EQ4N0StvpZScrosOOVNSvsdIRlAv0rLP10SDxouMBICcz80iMhwts
T65CfhFfAdvu5D4mXmSK6JCuCFRjEu1/oUCMyWy0EW1wAcniJ2NeLSW7/7vk
/h2LhsA26uQzpdVNjiO1q0prFTIJL1jhGesdBxBPQZbU6eYOu0WGcT7WumFN
B58ojn/IiboLsjJ4+e8FFUHLYVLI976xMObYPXYwr8wd7Fs/MPm6j9LEvjVm
Cl/XCnFZ29Q9YIGEuRB5zucBW2Y9+RCS1uf6u9y2+pwFCnz1bHNGBWsJVqXn
sSWWt2Nu2etIRcIvBlOKTB0RIVSWvd+C7Dh5kn3Tsxj2IqxrtT03RUSod2Zp
R5MSK4tv7TMRqYVxrwo2p0YYEoOBsWFYEQ6CJhQ1jnpAIIt7rmd27/gTwkAc
aMRp0mr/B/gnbH0W76+87vhV9XmgJpCKwmFWrjAj1MFb+RAlrgfwHvlBAe5c
bQhQZDgI0Wa1ETIssw6KiCXLZss4scRF09zgg2KTzxnQqLBpHUfXtBjXCCXf
qbbKhxDuM/xc2XQYDf3ak6aPtBqmLIKOujfFVpQCZP+sWuM5rV6etKCwChUV
MgrCNdd23V94XrsF3IbYqYawOcvi0Jx0iOCAjQpDXmPB1sQv80T59qs6CU9U
2RpI+BtiI4lb38WlLwrtwWy8vqeC1D4kb9NQAk8cAMNlPqcplU7r3me94bYR
Hs48XVPBq78fCmcMZ+upJYp+6pw18V7mSz/eCRwgD4fSs5plHAxMbl3cnkid
j2Dw2NECKfsl6UA2ujrsxLxpbfUebAe/GM5W7kq7lezNbwANDsPGW6hbpTj3
QUbiXbcePxx1yAp+jxX32+FoPo8Lbxs4+e02l4IxYpOl8HVPi6DMyF+gJP7m
TSoCcaOFNP3riKmFKYllR8fe2ub1p1PGOpcULl46IxpmjOSSrwQ0THyqzjzz
p+zlVwIEJ6dr1HbqLKFQXavhl2Crd5OeJ4Lz8K3g/mJawIvuY3BNow8vTvR1
LEvjHoY3IgBx0d4PitpIRDywtV4IoQ5TxFq+soarg+HY1T5isj6CJeFPr9hF
3uMr+1E2G6LhcFaLrMib3cVLtEGE8EG1KofvouU8yuv33NEa2zM+Gv799YMl
noDnbITOYLnbYvXAgaMw78b15Gw/COGPpe2yc5dUZLzMK24G38w1+moBWJ23
AT6YkR/iSPWvoG2H7GlBDzNNuAbPiTe2+3d7zXvKIHOkjUezORmcsAMfq5r7
G8mXgTev9Iwo6TEqsAgVWARfwtrAm6wRVr64Qv1aWX9spKOXgOoLXFG5T8bT
AiAMhHCeAoGMRTixrvwoWYJ/nA2kTaBmwzGj+AYO9e236xtIFQwf1HGfTXEO
Jv0bvzkvfL+uR5R21K8JjC8zsDPcPNFFvOsufkCsxT3HzEPRxefY5eTFpua2
mwQ0lnLjf3HEdLitowxffHox66TAzY9p1R/ydhzBb6IPMBsNyBVE0+w+RbBi
g1fYfBp312+7LMecSTQPKtQ6OAZDKzYITkkbElt4HYsDCiw9sAOILa8z72AX
jtU+cz4+sw9v47AKC3mP/Ujo9DRNy9a6enPjqpi42y0CntC2MqHGMIPALdz1
6xUF2GsWUJg473UndC64obqKlBPEr/6jKHSyaX+Dih+XK3jWuGmlQOkZg4xh
yUFxwdQKpSApUnx6F0xGKW17uX83hgbfsF3brlUT+/A5H/RXyVtdYdEQPfxD
sww6o06MlDot1PaELXbgvEcu3RsxlvRn0zZVxG5noWAC/BOvTAj5kY0xmifD
gArNYBJ8ExmCUVC2HYeYlmHcONI067vCCERVNEMfuVjlU6UA8sWMzFECMpr+
tTVKGZ85T6FVBFehH08QmoJQshbe62SbNgs0/ORGpZPxZ33nHK0hoswf1xpf
MH0Ja/UvYt2oE1AmS4PyvHrE5ecwZGpr7Sg4iTWe0EHjwVz3fOCCwVhkfwla
bozaZspKg1dMB9Ux+bFfzU1CH5YSEkIFGzY3DxpeFN7xY+gOXJ4dvHxURM+r
Z5tVxJjP/1VF5+SLAIOiqJA2ttYAGeE8LOHVyUUYUiGoWxugkoIq7FUoaZkC
NQQO3GxvhtUJm/1e2R9UhSeQaV3QJQbRnGZOIfudi6McxTVZ8NFAOFfaQo7R
xjNETFlzxmcG4H3t+CnmMRwIXAfZ0tnHNtU5AXPJe0ZKHlpijjvrMc7MntGW
XLaImbFZn3UysBXpEdCQ5FcQ0apxZBsj77FC35oKnMWnJBQKR5Q2Og8X+356
MLUxTqvto4wirw+cGMs6ZevQc4abpzbVnyXnPsufPyHnp6JnXft41bRX3lEx
M2+4VgCzq0agPUou7N/3Z2Zn/5lC0JxFjWtTPe2uVyqNBns6IpR5Raam3AH+
S/4ifQgj0zqbnP1NTsdqkoLgNd8TUtSKijyTUx/gHxLmxLe3eczd1jF4g+8V
3v2qNf/vdkk9+xuSUKt3WP4bEHUhVau0/e4sp7d8Oo7+Y/h+JjGfF2P1V3XD
rlbYoowPhI9+J//jzxTq5hAm8KztUTrAqOFDiZ+J4Ld/hRxWqRC7ORoyLesW
7bRaq3KZBjBlpodaISFfVKDgCW8Wf4BPpaN09oAgCrfwOrYjVM1ljXcdPPo9
ulYlYEzfPzFHSScYRLe6yfzIfHYPbuHyd/HmIl99mWmFh6C11tG0uI7wDrEK
kgbbJQDJp8odBqW+tbBU4jhKmUUIed9w8YD0TqFmHsHDYu7r/q5MPMhwV8I2
Jcw3JUK8M30B/CaU0mfZJP1G7X+dYNf1s/boB2sjofKw3f+d8ycP//GVQIeF
3qahdQDQP2P1OEAAWABRZnXETNIu88+G8JbIwEpIBki6DO86uHhzX0OCz2y2
3KY/JXW0LIaj+7xXGaltkuDEvrPIG+P3ieTopH6LNFZd0t7lyiicZeNX4DIC
GEHzT6kGFQeAjnj49xM5MAsGTf6MyQdMGzrCd6rgO39TqfJNb6PxfxzsP708
DZ8Wj6HKopRMqSgtqLqJdybWnjnunjHvYfQqw+mEqJSCWu9wPh5sJ7NGACZZ
wcDBS+gt2LOwX3Jwe4xlAWjUaxn94YBqIFvSSyiHjr8HXgXoRcPMaGHLPfzU
c+fdkc3pJPhpa85U6HhG7PBoA03RYzFO/zmV1c3QoGvoTtXHx+MQo/71E9YY
gepSH5qLMi5EeikmctO5Kfy9Q0gJNF3fEetK95oq84wt42y5oxiDyd75gcR6
shkjdJZy6aU8FE+3ED0owqIWVVrFQBQS9ZW4zDvvfHzJcceAc8gPvRsZGzVy
/YUqkm52wlnqYj8m0QKqodLEZPe0HzxlJue+oARPpVJq/ltUXBohA9puRosQ
4Z0HvDPIE/cxxBRLaUBtAnjbBi2pXNegaq/Z9LFwowQrhWcWNF4I/nWRdHmj
xssQuwvKv+yfMQvTdcY+xEtjon8cz9ZL+AVDcM0irXyPaPPPZ3+fVqtJjipU
q59iA+cn4vqWQdwzHlbhMRWxUlBKRp/Hip6i14vEkgg5Dhe1U1vYXeZMP+By
SRiODnSgJpca6KgWZpmHT/GC0UwmSGjZuc1XqNTpqjEvkW+vT3AWgty54MBt
SOCt8T107ZBwHephrLvcVmC7uwRQ8tbgZ0UjdVsnD0qbh9v/iDKaGLi3RmOk
eNHb3HARfSdMq8TrZuBYMMVsWEgi4GQ3n5IUWTBQrBh8ZkBwpm4Qh9NQWKCm
OPNKqvtmAMTXXP2aa9jzGXFXwYEZhItEiriVdpnb5VJDqxuFgu1yVO8Z+aNa
WyKi4TtX3JwSewl4+FNrnoF4EzMiK/uE5xo+yzUBSDII/W7cCSZ8L7SmEUHk
wmfy26eXsEGOSddX6xQU9RbICTddJkCFpxMYD6uPv+tEdWKSMFQHAalTPBEa
50RKV4beAhsXGw69B5763vglUMFVQbj3jYdLbLWqPJ+g1gXYumzXBmLesvEG
INXf6nUVjZxa5Pi05e25nd3ivr8zEby1Dhd6yEwa3htLT1PNgcZ43iiba4M0
n+yT9TdDwMbRrcpJF+F8yTOk61Xg9Z2UVDQgjpdJVOErdNgc2kuzQ9nmhU4I
xdwN9rsZCiRJ1o0RSiDqic+7qx7cGUiZAIOR9VwHzIeLdJFfKaEczW6DpSrM
DLeSuSMU+7saanGOSo95uLBlObyczmuawCK85RAg8Yqb07p4okAm+61A5eLa
2oS3lug/1JtP+wpADvrhzxMxl69Klc4CK64nS66DEgpaxsbZKPTgU26B1bCD
NJaWfOZgah909dY+R7kYJKRgBmUVPv7SB8qT+/BMcn137BAmx1HyF5nNJ1aO
i9L3OO7HCk/Es3k+CCgX047AfC723d+BOHBrk94BTkoJifdn7Tj5cRffow8o
y4eosU31itolWiJ4l3JxF8Wcm+1Ho0imeNIR8cgTO+gZn4NEEnvI3YYikdQ/
aGzxuQ3Zv4v7QXm5LSPJ06lOXroDQGGf30xjQ/VDjwl0x3r8dCCkVAzZ4JZm
vTjkRO9UkCptGv+lkGat5vr8i31a8AQnXxL2Ai+sWlfLsl8j1Yz0AsjEd6N/
WsuvRGyW+RCEbAF5/ZN98Y5pLQXDajdIsxB2dhgxI0Wtdc0vRvYxIbsUTAU5
tb+NK8gctakO5gJiDUPEhQ3aY1P1RBZnoWkP3RSjQzXA1Rm1JBxb+A1hSPzg
eVMMu3eU2C26PdC2tO3gQz6JYwWagLw7XtERTxYwv/Kxv2QoKVqzb5X4m2M8
keoE2V4XahUeOY6oFK6OPH5Up468CRCzPvypEPDPJly71WOzfSQ+3+aK9gZG
eAuTLpyqzKK4F+PeRj8BscSkkPjH3+viv2Tdjdf5Xn39S9D6IGxb+GNjEyiM
3ql7YQqgeFkvIiRi5V7vPi80fvRacEjgh0ae8+gSovKYQkFIIOAWigKAfvDW
2kHH737vyJYliI76V33jF4FJFA6bvEwnFeKB9Yqkymd65cNaWt04j9kO3Lu3
fPVf2f8RKdKZHZI7Q+TK1Kr2mIL/AeDhez5FAeV8ZM0B42hFQMOzVm7vltMM
HfjLprzYlML72Al/yK0uGCB/fIQU+FMsiBTE6GZ0sM2MOtEethWjtsVDkJOK
nmqWFbwtjVg5laJEKoRxKP7BFrJI7MWZQp1+u+QEQW8O1CIBX5TYca5uAlKL
RwxWV6XLsD5SnmgmHNs2vkfGgC38Xr7UiVIrW6LtpsiuH7q62/aIj25X1DqJ
Z6rwbtuEeQ1UWzgkgEePY8djswVNa6WPTPlVKodCRGj3MMi4ljxEditty/mR
6elOSy94pZGxeotzv2ZkXc697Gb5NGc485XOfLrWbOFoOLAFklWc9HMGIQxh
fTaChJmcR0+VxkDT2gdAkefsTe2Iku+uoO+ppUb6I4PYooKh17Q8PffYatJA
ycVkRe3Y5/oXqirciih8VKJy0Eph7zcaH+OyaztkWc88gF2CL1Cr0WKKW1/9
He+v9o3ir9nxYyu+u6QoZsrxDafaQ96Fk6dOPGJ0qBSk8zqVBNb3ZoD7OOWD
FSKllFvJVFDTr9IlDGDpmuapQ85PmXyQy2qbWsk5bo/c1gSy0TW6Wa91k68J
bG5uLv0fKg2iK4GNFcJI2QIFgTyqx+nMykUzYFBDCvOvkEqbwYqXbMBZdFn3
8U7kLi2qUxbl1w3y0ZKM7+Ynn223Z3ApMFFfZ1PAOhVKaVV3h35OgIfeHfBm
pSGHVC47YEaPAFbp33i3uda2ayuE9L6IKA6ejxXotCkbIPa0WDGl7q0o+86b
WdQy0W5PuzJ2R/OX3UtK2cNav2C8s7C2hi6Mz5nyQU1w//J3R9H7dKVKIaFt
NPWlYqt8kv2dqUNQudCZ1Sjhx0aiWZIPHNIhp44Ta7o5+JUrpDN+H+21u7nv
BX+3D7gfgrH/A5WOVtfrmyUSun2kJI1kjiw/gVO9KCDvIQfUfsJJnk9GU9TC
8yUUZ8nmSZm024I0V/2OjvabknqvuGnqUhPftSO0T4r/xfMOtfSt0/IwnN4z
RlEQUnKnf3+R+iZqxBbDnTmn4GfEjFi0T9MgQb3TwmbkZZ8Rb8B5tAlYgtNX
C6trFtj5BP19r0hSdXtvP4il91LA5L4qSlN0edahtleFnhWxk8sX7NtmoFBv
yVlDDV+vb/8A5yiaN6UcnExhZ3CCjfNeMfeeu3zqg2Q17V06R+qjWioMy0Yi
PeRXleD/PmS0BFn6/Y55xzzjwFQgcn9YckinG3pXIr2YHtwdPp++vlavx/j5
J4OskxNoMA0+SE/LVrZytYjMzaMB5b0utat8TjNsgDv3SRUrq7FICS+mwECR
Bfm26UwNu/GyNTTGR4HjJclGwnD3pj8pk9RBQLz5uVfsV5IWZ6VUxV0xptXG
dpXoj+rnrAAVLil3IvOuYRbCLBhAlF7jm2wWZYAAXAlz2omRxzPhOdzWf2zQ
3ZAcWYhaKWknShonWyc0CEGoUBQTaucy+Gl/M/Z7nsW4WWJaYef562qXK0Bl
/VnfnkjwkO6yogh6DiHHhfV67l/G2O/DvD/rnt284PdI8Ua8Irnyen/AYDhO
fZZDquuMGr1xwLFR9ufUJJne4HTjUrcYikYg9f60zd7K61w2RyOrAuxCGghC
gx3RKZ/dBvFxH6eLpBYUx/feEbUFC+I3HLoLDnknQp9JcoJLwGwCah80IbvZ
e34CrqoaHrFnk/D8/4fJY+xgWAOa8OXAIQbJ0NYrkvZm8taBsHWG/eQGHOFg
agtbG7/Jrp4ml80/ZQlhYeg3+V5y0GTemm0DFga533hnvAQ+hoUDcIgxzyyi
sFnnQ1JHo8pxcqdIJ/PSb4mYmJMInoynwGccZ5oHXRGW8pCJRtHjzLeJAWlk
7z8HdNfhT1uPKvvlAHBb4QXlqd6D1lg6hx+lQmDYSh7omzF2pGiWVSXrAaIU
wo00nBojZ3WRCD+qfDacr7tC534MawMltYB53M7BKX5bchHRyFMwSZwl71rJ
XV+t5R2cLKqrptD/zt6yfilCi5flBlVepBkau2kThANb6BJQtn59s4EGy1EN
Qbg8F6bsiCKVq2w3fllmuN5h6+fM2gy9vzilV9Et6B9gmf57oOvlhrDeU2MW
cOB5kvTCDS4MazrD/EAElKpUV67jAUUv9tDME3uy6JlXhi5A/328PH9G3LG/
b72G1v3TCebL0hhFCXIJ8+XQVcY5fefnJoUzCU5ySbhtZPgvAvoVXWVId5uI
3wS9WMdSvAoCherEhgrauaFBuxSUrV9rjDx34wEj94LXLJBhp9ynViC7Zc+W
j903cp/gcNPL6tDdJOmz5OFHBvqhlfYemrCiwT9UrCLwDux9hp9AgQVSXLUD
pLDyXwNCXZ9OdFrPo1+aLCnMwOzezuPXlb16t3DAkWjir9JFgKx7jmHUnf/l
/zuam6/GuVjXpU1WX1GeEpfR6QH/Z0ExqTznCB5VNrSeJpnG75/cmuZTxhtS
mdQzOVHz0hteo0JyiZR7piKRrlpWWjF14RDpSgEMgSrjSwBcLUbUNoo/uh2U
TUXQ7kV60ImKI0jLieNMQauvaBXN0UVK1a5rdiHwcraKgOj0bzhTBUwM6keM
8Yj7ZBiiJd4zNVatkaHMG2gyEqqGhuCC/Kb92WNV4AAkVGKRyvuLp7ej8haI
0Xriz2qFAfHtLOG7YLa4DihQUU/zKMcxxeG5Wp3CTynHjLJ7UQWE1JxVZvLI
6gpBiVbyYKavfNk9Ov1YjVRUwdeF/1Q62Xj7KpxaKxhUyPOHEbK4bqhlV8Re
fl7pCqbmlYJriA01pxovRIOUibScPmHgpm2xK5UMCz2AeltkutM4QKL9gP4Q
TIlfAm06L8P5CTy0V2KqA3gXNKENjp2dPlVldiRcp44K4hMbv+AsMkdb1H4M
W+ehpcSnuVcc9zQWcKNTEdcPAY+fS8GEMjxm4p19A+pO8WSL0xvng7/1JjPQ
p+JQ1khjOTInfXm+KfBhfUExfQCmJ+stlAoQHyLpbyibfQ34dw/9QmoCkacK
tFYTLOzER0pzAljvdUCYZlSX8YwM/1/JzHe03w7oK/Ek95W/meWC1LNhnCUM
RexKikV5FhAUtM/301LrbEscInZtB8SbW0EMzEoGy0l5CqIkuYRHPMLwJTqQ
KHOGkxUtNK4IofB/66WTTSUleseGtOA/OdZsqJb+Nslm6TWfPNwcC418ukTK
w7VIJ0Ni5NwVUAp5Vh3Y/nZ1HOElpv68VvsCshSbHoyridGD/MX0POmKSlpl
c7a6iwvKRzyNZVQMPRMX+d0TOfCUDrHiXlSEnY8Uw1G2NaV0sNgSqA90wjki
fCXxYDaBns11GFKgwWGWp3slncLdIEJBcmP/A5HPC4nRBe5lTSpEyUanA8gO
iCf3rmNllGBWWIw+mMMlgkhk2yNVP+w06o77h6fq7dcLyZ0vgMDGn3XIdQYe
/jIEHesZRKCQo6dtcOl6VRd157QNKgzqa2j4cx0B3/he0bt5SGuAp7DqbmJ+
1O7vbpSW3B1gqDbAHkI37zQb8XIBasaJsHBf5azRCGh/l4pxVl87nKnoWO8b
NN0sfEKMA6RhrsFbOxFzJXZDdSwN88TW5ocW7BKwQum9zM7v457LMzooo2Zt
L3Nyr+BYaRWS+yzVfWyCs7WDVo9uq8NzZmZz4lOd7EBZm0sOHOlJZpSOMhl9
xSS/Jsf3aajayGMpZ387D+i34duQdDduwowmQMYPzlvfwaZYAphiZfrKd0z1
A/Y+6tEkX+t7T4q8rdZ+lot6GgbvTrMy4+8RlevN3KbchepOrke1u0CW/VoM
rByya0Uc8HSoC/unhR9V2Q8gVOUkQDGj2ri5Ul0I9lp51Ws73gCRpo90N1ao
SA5pDHWjOY7D0Uo7otM//Im8X75jgIzayG+9vIvsael1AOyyzLq+T9tyq1L3
a9Yjkbitvg40Zne4+sgLEAA+xcdxn4FmXsvQPFkVHEq52a/6cEnzQxBgwVmJ
WtuOX/vqYhKzGvxtxaHD2mGKV4dEqju9KvwKiYq+T8TFuUAKKgpppVaqV8DH
I4prgeVZ9gDNAzMpAJ5D2ce0Mfi/tcAQBHwSH5b9DGQe16yyJ2a+eI+fWPiK
NvuZ7KVHIbkibXKjmDvjAezcPgAaT1Mioz5qEorcNWxDCuC4Q9PrkrRuG/S2
qSW434lBQdLgbcHrQeGDcii0maGuaYqvHrP6jItw49kr3k/zGHuR74GNd0zT
PYI07CqE+L1t0zntpTSnB0OPR2dPfIV0NBu6IuO9um8FPl2E6EkO/a2agCZH
k6o111+R6xHBFPXwmSLYfYfuJiY348Z38rqJVBl288spHr7Xsk476LDfHZoo
2UZKlujZ1lljKLJz6bd02AE6Enjj82PDSN8KGKXU0MxosAMxRa9xoH2bQ9zT
fqUEeHSe50oTbY7EOGr7m0FZ7OsBvdwZpXT+Weqs11b91dUfJ2tkQEkZkJRt
xpiUpfDSBdwYycVsQu3i0v6q0fCyEZ/fJZqdw+X/lm+QmRtUgUfZD6DAwC+A
ztJZ7vDsd2h0xazqaKyt9pmz1nx5CcdNZOXS5TVXnAE/n9PWwbXHrfr3lS68
VJw9KxurAXAfui2vJcMe58ZPeRusOROy2CzFcQ8lo9L6QLokOuZE/FxsvZS7
9P/+cKP4b0qjrQk37gvalNQWPrxEEALArmrxWcGN5iavqVxFnxNVBFQFDBJt
IvtPHToLawEec0YHmtMVz2MOgxXHQtQlqr9zn/3XJqj/7l9s8IPbH5bJonHi
JYXLuXN7zKV0WSbiHdSlo12pM5OQ/PvXFgagVqKU6+SVhzVnRwa4ovPsbiAk
seGxWrZMX/wx96JN9PbDpLifhfvnBkh+xO6avQn80dyPPgj7Jc0YdNjwfNSq
7WnMztsteiuwiVui2ZgUKFyz7oHMvFw6BSMo9TNun5BLgvToMhbn98Tbg36X
OT15oFflbLUvkg4Q1CwxrAqiblkd9L3jSNCtqSsGqUhiwLlvd3gPxw7CgFLp
mMO/5JSs8pFf5iemwlxcy+i2xZQ9OAir/ZgBO4HVLDtoU67+N71n+PYI8tlo
95fAKgbtkffgniFwjE/+za+39QNnrJe8bic59kI67j76vJfAx8Ny5wIer3uz
Yytbx8d4JYhBe9rZXTN4I7VgYKNdU8rR2a18GYtllegq31DHWaVqq7mTSDpM
JjLZDcb/OzaYiX0Tj/9bCaRcLi+AUtsv2RY5j4rdvlvfn5VQaCxwB44AbWzc
dGNy5IL9X7HXMl47bBAZ6uMDEckVbK6Uae+RX6Nun36TWOP7vIKZe5FsUzk0
4RNWAyqdUGTrohce4hOJuq2FJWYxFDFYbu8VaejEeZ785ZviR0Bgfqwag0pA
xPYkX1vJ/Op+kAxkQnw82iTLR9g/jIYZJS7dpjpzp4JPH+Y/GV0+6HEOIB88
Gj+XDW3i6wIwQBZWgSAvUUAz1xY1Hy8qLTgsQ7FbrJeWjNu5XRbQGDemBn5m
6RrN07qpbS4dGW9GbTlHRbYsDtB+Bz6BD4yE5lxqnkwxNs0ceNpcnOFKUJgM
odOzddpSvpzT3AGdqYQN4bIQbrsppMgXQBPeQEvRlz4zp0iFxv/s3gzgWuVC
uWAA4WzIzxfGpiNKJcXsdEDxCBVzo2D4vbP0p/FKg++5XUwZtu0E3B+QTrp2
pD0ypxVr8vCRwf+sAnRatCSy7bNvyb9fkCPaU8tKvHyxJ+86CfjGUd1nPCwA
emQpYWTxwLaAXdlahQPODQOjYv7vkRcMT5eWMv1qarn5OWobZfCJqTE3B+on
f4piphZ++D+gMleivEiC30VQEfi4IRgEHVN4lT0Y/bV5zRUO+RmJ0FK6WGYL
nIsygi20HVRNITL24V/ZgSCNjXa0v2+74T5MIJ/Gl6Y/qdmweYQA0DHMm4nG
As5s3QfpQUMAKj0Z5K/Ozp61AsGyR1YQAmp0jHLPU+GbastXJLJ0nuMyvG4+
VMllpKHFgZ3+mxWM7/IEtm4pZPnuNH3tOfYnJaKhUeQ+Ys9Ok8R4pxnHuJDC
ySNgyEKkUdeCIOnBF5h4vfMjyz59LZH9GcKJnQdtP5i+QFpIIdu39yhwz2Vu
XVB0rmALcOlpvNinO8s6QZBfw+LT222xDmxPXDarMphTYof0fF8lt8laS9Dh
6GmXCkA8qGr4wzlx+7vR5/X8fNuSq75Uom+lhr19Ffo93Q+qOJFooFBx0tHD
QHLhgQRaXwToEjcAsJsOhs+aYuSRx5HWNQKeRnlZwmug/yAKaZjZR++/5cl2
RWEBUkWBQnzXC0MNkJvhKrTRJuJMDlb5jJz9L8Iw4LlddHmW16SInAnog8SX
ozrAQok7uHayq8SYRFB/FRZpUVBmxRZOJMHkQphW9KJBkLm8Cv5v2U7ZuIEH
ccOjofo19T0oVb1zuxd3nhtOVLOSWyfsCBOg/+tUFqYhq0E2zuPBrG3wCy+7
FNJAgZ8H8UjQp0JrZhfN67h+cNzWSoaITrsBVr5NqZjRhvtz8ayr2As0W3RF
b/JRsBk7cPEmjMym7Dw8ujbMlLEGCYQe0Of2+SAD7vtqM2wucF/LyHHHIVZB
A4NyIe+uTS59elDzBHHL4/So3ryNJRUsP+EgHk5qsGv8yvDYKfoNC8a++S48
9Uw0FKcHqFlkNmLKFnKMXdf64uWGgdx0wHLDUReVz+0lMmrQ5SjrHI5r3Zk5
LppxUTj1qCSFyOQvMzoNFmyIDg58tO4A9NM01cZywpRsJRsgDd8LBb7JRROb
uqJlU82NSgwmr+n9hKxPs9e+JlmhUq5tH/KXx5/CkjauGWJzvyjDKlmVVF3E
dbGc0ABfyo6fB86aWWAwKVj6xj0ADH8pd7NIMJwPmfm6ZAsUx7Jx+USA1Oqy
wsMLrKJvJ4SBU4vzD7nM4JU1CQh3AlFnz8/lf3pNDAV+OdAaIWPwW/liohIH
f6ISq/TP5Wy9rdsy7bpEuxoMSug2bQ95etYClpLOIyjzaNt+s3JOmSMLA90I
9P/pf/l/FaRxFx3SKAOKeLQ1mRq/xIYjsn+7kKm9+Lwb9d9VmbccYDPsMybm
fHQ9hp26eQRrBV+9YTWSwV3z//ycD2tg1x72wcff23gaTwu8Dn6LB75Gnqgp
8kOdstKDBhmV1zvjYEiL8lnX7ZCJ1nGuKFmdK2IODIQ0Bz+mapvxjQ8vb0ul
BZrDofJsEr4ArQhKdulVd8AewWjVQRIIjSey9DeMFU7089e9ZPNExTQGD328
eG4dCHlCMze6tYJM4eO7x808Yh2pe/d7FcrI2/V0smhW2dBhbi9Qt45ctwkY
U06s8MI3CclJqByVTFZ4czhbFVizJldMYzuedDhXhGgWBRmTLYSlxw7/eMFe
LAJ2Mk/a0F16ZBJneM2ZAEi+8UTbwgD0YG+imP6fe57OXYW8tgF/NSph0VMG
Y+PV1k4eAXT6vhpxauv66gDcMWDL/wQJex3WaRL7P099hDZVpd5alIrl5k5C
+7CgE3ak4DYZblKfVPce0N93DA+IiL3ZoQAHTWCoCHwUJdeD3UF88A+/ubHF
WmwUGf96pTGrRhm0akKrT0k4ZoW6RdGMsLEAVAws3AJXKQAF60eNrYtW2vdf
WoPnI1j9UgIS2Bzlim9P9iX91Unfw5LHj4R91ZwF4CEsegNo4eDj553CGJFl
GytM03pY3IRFSQoI2CwYrPlFssrqLqBQhhcAtctRkLvroEh6w5ljbHktG8ht
SBphBJ2kzGeG8l9rqjDHxMYsV+Hbby1gjCuWEd4byGkoRD9DF/413FScsROV
KBzafbfZkU3gh8Q3rgif0XSaYO/phFJ0nYul2MpfKXnFjz7Hlbf6qY3xjuye
KuPen0rsRrZLWU+m29Sypgkl0qvgFqblZLKej7fT8ajJhsRxk8aXRc4xz88o
xEH0FEE8AHBWBfmOMSsCQF1xEzRI+KolyIzn0U3e9jhHh9ZE9TR5YY91Shk7
FXyBjHXpdZuzO2s/7ims/Yk9OtuANcDXzhXUqFPol9lP1+Akbsl/cGYFC+ZX
kQyS+VY4Xmux4ucBOTsiDwXlHMrtDBG3il4E7OekDaHjBetRpdMAl4oT+nq4
1j8WWudGQs2nQymvPNDcSWECrf+ZC2tdFuVzpzBwpNxVgCuWGQBju8TMA/HI
7bwXGysgQZYSQADKt3VrSzAF+fZwqaYcjnwH4VoVzTHMpygI3ZjMlw0J8fyY
dk62AHWCYwEyOZ7VhnIbS9991MQkyJY+zLZCqmMdPKS/l3DjON8krw1Eb7S5
7UDkpHBf9UbjLZx/G86PcszubLIeWlXxfXmFb0cBS/WQnmjQD8AAksyJ3thG
XStYfRKaQzhAih6gd1oYuFKOnkegjsr3d9GsmhLcyyb8N95lRYIyzFPA2n5B
0Uzh8Ag1lTIufz6DsIUsqs6G5KgbBb5BPw/5sBARXpNFt818rc2VbMXzJY85
5wTalrkzM51RZczSTUPAmd0lM4hzPef/cLWQ3uhan16oJ1v0S/p5HjxBQszy
rdAFSAcasENLnXn0ROGocjC0/q88QbY7kAeg3ACoDSgxYJganihVGxqLFSos
n+WT7VxWUXKaI1IiYmig6rEdeFYUu+BbcnC22qkkaX7vAkk4qQyyvR0oNpsJ
on79Hpiwq3bkTOykaS+yfCvL9OQ0iTcol4WeMGavHlNNMgBAGF0upC4SIijP
F2fjMiDmoKnQmTwYEII9s/jrTm5P2TkjpsXqCQE+MjhWgrQqdCUJnOso6Qyw
0K5tre5hzzzLMvc54Mrwiu9mzruzooLc5KY/JSIItS7DJSoNPrEA+uL2+u+w
ukxrhQkos0MTpP+Jgl45q7iiOu5AA6k44JYj7OzvnFXikU6kKt4/kyDLZuDQ
cA8bbVC0Z1GMygTEttCqTeHEb+NQM54WnjbLDMCgovR1//3DGy9BGWlgDzto
JP6C67NtobFDHQ8WBKqsctutUMVG3EUPKxTaTGlmHU3edERqKfw/st8+98vV
SrE7ADSbPNQ/Yui1++YZ8cTgK+TRj3M1KPLNzs8QDxLZE2euYnyzcbSXL/E3
yVo5HNXSeKGg62qvRKibvMvdzgSCsmk2kaxnEl9R5MY8qpDJzzq67LFKpxje
eo5X0JNameaFuf6o2pB9E0NqNdBlXDv+KWodRFkO3PuK0juF0Mm+ezLvecYa
9TN92gT8nmmpuIdndXEazAhIT7DgadJXfCvyJCBdSYcgpXcN5cwXweTr+J9/
4jAMPgrgzRUNWTFqaAI4Vcq229ZWQKD3LdxKyjbtT/4dpMgde8+JiHz8kgtu
8oVf77gD5Myp1967xfoJVlTg4lkN8XqOHCL36Yk1S+jmsyKNErsSCTEYY1ig
j0S9yKJE04oYvbGaKtfmfjgz5Bbmcrgwmg42GzsXBLI37/7v+MyxySE6M7qC
yVI0GTw4noKKP2O+TxR/AClD1jnbXDytCfKLjCzJJaRSs6AJzCq69uCDvyM4
pOgfYBpccYYtrPmvjhO0p9L/wo9sMX9WRQ4AfTZS075H+jVKVT2LiBnBqKx0
PUqcZHnMs0/H3IX1zUfk1+SlG71+DM2Mp/MXpCbXGacnkSPTm5qNo4Sfalu8
8wZWO0gvroUwy391Jg5/tZNXfNtLR5DkkRWYkNnWdeDlJKHwKdcJm8BFEQ9G
ar/xfU0zD2el3b6WL+K4mMYwQ9jbp2Ts0Yns1Ps4p6Vhu3wWGojTyPIs5wYE
xSdtHqEPULoUatO2ICDwWEZ+REzfXOEw9iJgiZ4RSklxRMjqlV/RTVAOP2ha
j1KESrqhc3/n3oszPuBfmHHG69kaESZoxBNAc+WC6MSi5393bvtyY/Jj71ke
9Mj0WjDPYVDlLo6DCBgxnBBNkLmvUHhlJ6YwLKBJrZh5AtjjVvEu5mjev7B9
pmeXfhvwCfCVOZTHluXWf33Ra+VOmfiyfevM1Xqt16ecBpYDBnv/cSCPY4es
JOqPbSuY2IovwktDNkEicq779peE06BSKex4Su+XmjkrPk8jmlLoHSE8qqZ8
tH28GYvgSfDGzyC/bGKp8TpWNHK0YIqcW7GqPnXDpdVC9+rVAwS2kUBF8SjI
uGAU2xlgCKhVbmqBXY6ks9dXOc7kcGf2a//RngOFLwrjIxNH6eRmbeekThmV
bEHmO78YhpiGz9merMXrz+773inNcnMS3btpBj+bdZQhQXjVKhvoRmXHeadU
luB0R8iwakE0FLtHcvq4crVXT8AKyHhEotMkJZ6oAjsVOnft2ZeONSWmQGdp
PUIif93nSr+gfUANAzH71PVU0wi2YKOmiu7A/7c4bfMVT23W1iPQLv54n3ME
b7ViGP1YNy9L2es+5nyuGkd3IHC8QubTrHsh/++R2vWlGHlCN8e2ZRzLPL+N
TXE+mTBwlAmwWDVkvV+7YjhwYUlK0MW1Brlw9GSAvN6QYPtqpfgEn1uceACR
td1Tp1NO8Tv1ZRJs1DAm9CVaY1Ldo5oFhABAJguiCGMZMlFDkg3gS8wVMbcK
SfI7OKhIDB5+4sqqaZxNYpa0lVjqIYXUV6pyqTM1D2oaB3KdZL2bSAR8lbR9
ghN8KlXwM2aThDHi0udcMvE5Q82mw0ABlq3K0O2FQJqMYNfZ25jw2Culzzww
eN+7BARM8OLMuTFCE+C51onNRoqutazJhyQ1oHfO+e8/12O2AN1VYPJIISTw
CcyjsOSziwbIGeFVZQihUy7tYzVBnk10jpeRsxBWqcLC4/2xn7TnEkxKQoQK
znxHRvYHNEXMFLVl58gD/HVCDywGBDKZg6dA7P4dXUNJpp30Ef6uaLfboOE+
ReNFbwt9OCFVetGCJ5/4rfOsJDdpH+pDWhxbmn8TmK+a1Rq3tLIi6bGDG1pP
ZDU4mUk7iL4KjllGmro9ZjaQ+2xyYfT6X4ZHdqdeirZHadjT9OU5NfJyMOVl
y5qcWiKJZ72cyPqEcyTBnfvcsib/v/5wrAbiNsPsJFL41gVZZioRDguvdbkw
dSTU50PWkYQpRjwRaq6KbCeeq1Zd//YRMcH2wfUzLxiDevnriMCZeAsQ0FNF
pFYbk5/R24g6O0IZskH9WqWG9/MNl9+alQER8BIln/jBV0o+/9BAcyXQOeYk
LUxgCQnC564xtHvaAcZmIqaowFKfXMKwB01ZMwBOjU9qyGakgkLl761WKHUh
f45n7FkJg/SSeg6scCcBoW7p/slXJcCQ0FWqmec1v8cv3m6M+ZoHb+k8NftG
7kyHuTgAqJty2aHvvR+6WdtBKTJ+b/T40BBQQt2Bh9XSabOcwxgMHlf2qyps
eQpOu1iBF3uvMsnRh70o/d7W/5djZHoL2DwONsegTf06ibtV1uqwkJ/tI+nN
wBtFLpN5pZ3yuAumnVLMLvFFlce5lGqR1VKI5NR7Ku4ATrPKPvIVaq4ecemy
/gstrqTyvDMguyVqkl2iZNbiQ/HVuIonTBl6wI+jNGXZEOzzNmDgGOeVO4Jy
roJCD/QiMECdrcu7ztZ7RQ40gq7i1nHWIJf4Bljf41SLkAcFJvJV6uwEcP88
oL/pkXaLyu3rsOSsGfYE4a5DC+JFqSwBG2z+2qg1OWvDYdWUUKH7EcW2l8eh
oL68oNRM2xAxwSv0XQE4Q8tp5Lc2Ig1U/AwqMsjMaEDWDxOrB7oSS7+Ku9x9
jpCQ0GxVuKO0wbGonrtX9+1ewzGTNLk90+t6JD89CO1/syMzikx2ZUq4B+EI
TrKGWo9XJuiMAKQ+POm2kokevtkcWWZnUxXwfn4nGh2nyT0Ey0e275NnxC7x
gm88HyhOWhuJKfbcj3POaUpnRHFp7Bej/T4fC7x37CTlrWYmnir3vuiVWBn6
VpZn7esMLKcWbaadkhj9U9ZRFh21qR9DqUtZduZrBhnt/X8HkoM54suwO9qN
l2qfMtgTb58zRBX9WRfUY44yvEIvZyNaeFZCCUpisQAMyRsoMD23WTAnEhoB
Y7Axj89mAjU91mam8z9sV20DTroeL01lII76rZgQrU/iGAIc+xZwdBcJISHs
KQ2zJE6efSCAcAU0r/CV6UBz7d9vym2LbODIx1EvMVd0yzz/3E0+8UDQ0YkE
IJ+I5Y8g7/VN0oBHGod7e9WM4SO76xb4I2P6F+RBYAOzahxzyrzsS4Z4yFY/
LV/aiNK9CBo1R5jgemPZTCOpeZK1tLnjzVeTGM9GFDIuU5zN4odUpYhvHcwX
WGgfJc7HouMUT4T6Z45ViekoGlITxDwi4VTG309nYNHsybFKXkntl+YI9sTp
Td5FPXN8yMkZw5fBYjcWixJegU4Aiq/F03QnciSSO7ykL3ax34zCBaV+iktn
x9qw4U7C8R35KPqt0XMmdZVrG7c7FJZsag7KzxHTTGHomNbeCEI6Ladg05nV
nIrWKv1pDn+YZOblnYDZO1y9fsj07mgC/gg078LJjR0JCCpRUvgoM7eI3vMT
XRhXanQ/bJ+GbK54/ozNqrkK8mJivgObdjKejdb0cPopyXCYM2IgMNvrMaw3
eNY0h3DfdD2YjNLST8GMnsq7qiudg+CvH5cfrp5ezYcURqttynRQep7PPh32
zzMUgfD1ZRm2eU3cQzK+6qWIpTgN9ilcDnXnjN+ycXPoNolhyho4vhrmCXcW
8BViliAn9uZuSnc+RDWF8obTbmhYXg7nV+rNZdBWqzlMoGqVgtXqB4gAXIzt
psXoODfm3v/H2yL0gdATJF7xNhwMzSkWdRTWJpjofWDuwdieyK1+CWiGhar/
GPaBZJ4SBXDfFDZxSEWrPiRn5znwYjwy/h4M3bMTjCJJRT2PX37Gx0oVN50Z
NWtg7Wu0L/JWDkg8iwQJ+UPRyWc+mS2u1/KZzK5Wvih6J6j5a9YZ7px2sbpO
HF3lkN1O4TXLrukFEH8ECXa1A9Tga01X1GbmdxZPMslpXxiaNd0ZIBodwDEA
990U87iEj3MGmPqsefXzBUPbj3T/YMUq9h2qGwxGshwl9y9ukskCeRY0QgzU
umwv3OYdG6BCeK3nv+Ht/bJoz4jJAq5KTqdB/8A7CgFAkOYxsNuRRTt+v/1b
Tr9fkF/hzAKkfhOcmpHN3SLLCyCj4cxY4CzQf84GwSdFkgOdDjbZGiVxBzsw
RGljkhHFT63CpryV56DuxI/id79kXR1QT4apOITemGeIH1dkf3hhlEjVsPjq
mOAQMfTIFi4hNGRNCUUwJUXzLlj788/Whmf+lI0I27bLWZf2xr33QLpGtKZe
d0Y5EZeqEGR5E6U5yXGjecMBHz/GFk4eowBLi2bMnXkmdLfDvfr/YrpMg6FY
MlcU5JEcmgPgoIiWyA5NRGmj1Q5snU6No1FW9MxSIeGobLF2anyjGufBeBaW
WGs6FzB6QWzXVz+7osXplS3RwRTW0rKoJ+cGUYqTxPAQnyDNRaz0f0sxhuH0
37R+0MIE2eAdWt8Zv8aYo0XqBCxqq5ATo438g7W1eo5Z0k9FniTQqDdgfamw
xaboJebxpzUqCaUfN2MrjsiKAYBpZJfUY5T1YqFJwhzoIYnwksEzuGv3LJtM
0sCCyLkRf+2DDwV7imbmz77KgNZRwByFKIjD7euQoNAm55iZb/UnpFPXULbX
Ggap7GBkC9VWSaNXEu9ryQhX5Vb5tdwdeftQf5Wt1xsBRN8sIcc6QxgYVoQk
qA9bQ8eddeAGD1MkV+HdoJa3ObAq2D2X11vpujwLAsAoc6MHdagJJhmgsida
9E+uMQ+ziOmkrrAGP7Dwyc8bLrsLmvBix/ErmoGZk87Pp7UiQAn2QxUazgXV
v0Q518nHTaIg3XkhWh1xaN/5lh3aT74/yc1bRTHwEvk8XLYbphej8ko3qZN1
BUmsuib4kaKd1a0yyq5dn/7oBkR5TEnLbakg4355Lo8kYcVyt28dVDiQy/Mk
KdzKeFXvJMb9QSug6pFANOERQk1hc+z2WOLAsfljU6R9ERtZbJDeefq7M1gX
NWNPVfrFTBV7VY8gfZEEBgkqYpGe+7q1K9pj+aooWNrKh+KiOqJZCYkfoVa2
QV28mm6VxIkrC3jfAzO8uWmkO7niXDRtZj6yX3svmMl9WVgsyhfGJ/vZn+wH
pXcCmDSfbLgyQoGKEM7auc2Z52r4Pd9CfJX3P3nBEa9R6N8wsR9Y4vPOrNw4
FFIV3rwUJuUIfQHmcmC3mQjXyNFvf2ofcVlJCYPCf/eW9TrirOuWjJ/u3Sr4
MpmDq7znO+oC5CorFsOm09WEddohD/WD5OYgNU4yMsWXvWw58NaXMctEPzXX
+ueUk3horsNeBMVDM79JWWE++OvrkF+TrmTUfn4600QfE1F261aemGK/xB4i
9UwVloLDcsIu9tHZwmdf6Gc0B+a/HW7xHV4lIl+xwhopKsQJsJ5/WoM/C3E8
6g0QVqMyjcWdIVXhnGuBt9z+SE7DzCflrmApaHM1b4PPTbzkeoQo/uveN723
mXzawu6wO+fUwHxQmj5+7FQmlJ1I2WJ4m6ulfECj9LqsTVDX4yhLdtT9wasv
LH8uTXrV8pW6FR+SSXmvfNlFr5o4YWUKVX0+EjkZcEJM2H3zWQ4yuCEvhXtV
qxU872USVaxntYFLvIidjK+J686v8L2FIJY1AzXVzvbq3Sgof+uV/42aRfvV
XoLBtnlcu90I1aj3T5/S7cO0zTHY4cOW7SrWgrk6bh+eSte0sT8x8XaHkMi6
kDY2QmNo/lGgKFiXERNihzVtmBAcbrp0MbS/pDzUWo5aWz09NvGsunsLKp5K
pNXfPRqKUSHx5P7iOsxJOIrtY96rSLq1713hV8dJdGYcIzp6GwJzaOa1tdBZ
e2v7NbjGVLHuwrVrQUomuwdvHRq7+1yJDerHfv0q2iOEWxsTZWl6TWAsgeS2
TZUevmyxKRT687srNcboviD6YL32NNJ4eAciOOjPsBDlsH6zy63+ntihvtBH
EaBhIovQbwDtmymw0tS2M+5WBJ5JnG2mSOEk/jqj2mGwA9Lmm7qIUDBpaPwB
i+bTJ9HiaknQkcS8nO3X0V5KRN46f9YHuHO787UqAQAlOwsl9TTaiDHPkPIP
pBUFjRxnJdc2YaHyVgPCP8zDlga3H5gm3AfyHYfVvIKXmGqwwdpc9XU6lH8Y
hGhEL+I8QtfvpKjsLPOgnAvET0P6nnfw+s2fOlu+r9QCQsbbcIDa13ijH51E
QTnp1UQR3okoo9ZCajKwArXgAKMe18Pkq6Fh7jSsh9SH9c1uU8Y5IgkLrtxY
DzISzG3t/HQk4ORfItS8bNhQBUWF9pzOms/0gUALoWVBIb/J8Wdwww1h8Sph
oXKKuRlQQeCur3IHnA23r5bhxKqZNaw04eq8ApnzT0ASSD3zUYnZJUJ+R4Bx
oJOWzrlPlWuczAvPLIQ5dsv7ic23DkVcz09Syu1yQbCsLjyXPEQ+Smb6nXNz
+6VeTbn3Rb9Kx78cII5iiGqwbPgnVMaxKSzvVZCA+t+Brxc4l2KiOwUEGVn5
ZuovjEStgdGk8VkPRs2Z3SjyBhrArj6gsHKsvB3Zct+93iezlCY0yJtFL5K4
bVU1FMEUgvnpvaDnS0Rib1jKF9lsU0QMGUzzjZgLVgZ5YUD/ArWDyJZOb3Ov
VAEvbUKTvzzoOQIY6heTtIdU1kUmClp8ouZqEi/HPftKr2lYlYp55n/VQoku
TuxEhBEOVmW4HvVpmYdcd/qp8G1QCM99FR4XYjkuBq5R4aQujEoBSVqRN1dZ
KNNT5u1HuCQkbniMLP6j6hleiOcpobEAW1Ou25GoU6vmYb90xFFZIy8rDMuP
YW83Kq/FTZGz7L5Fr4PMcqev2z6hwWd+IrXB8WVK26mXGuZ1hIBLqZilYTdB
yORCMojpiY4hqUFWL6jyqPTP4rGwxxzIsP+3OZx5bki4mIGvgGoT+//g9EeJ
AbN+gMt1OTEQnLOV2I766gvX4qaEp/mg2KJ7Andge7llURBJozELfdOSM4Lk
m8gjeJHrlTdgP3MPRyZdJrcp1SGLBiWA2hwypwOowS4samv5xUEkgF1EUaSh
mDkmMuS3p4Iq+pL8x+MYzGgGp+RllgoU3T/zeAIzzr5EU6kSliXUw3EiOWQw
knoikCtW/ltxht77jfJ/41Q3T1YhcljgIT8nw6jmA00/0dC3KD7fhjX5CaO0
XKA+Y5v1xksFMtM3ptfRcUkOq6Zc+Sxjp2x5czaH20o9A4XGPnRP7MOWYMD7
ck10PPgHKy7G8Tqzqv8xfFZCOC6/4ItfLeS7tsdb/YojDdJaW/6pLfYXz9Gj
qoMzVIIi7sKkoFDD9cGTLdDuzJq53x/fAjS5hb5eLjf8+nywDi11dmbnk6sb
a1IUcF5e+Pui7zu/HHxSYy3azKHBc/IHaUGiG9hafYRNL7X/sRMuWxQYbKzg
69HOWZzp/3uIJhJIckRGg0a6DcGFNlpBUiMhPltZQctWTeOkqx3Jb+oPetud
A5qFSWtIgPiIuDuhW2yvZcQPEogOZSvy2pE6LPxHZbluN8Pv+SkE36DThEVu
XuwSuUA4f1jx7fTyMIH3uixIEMXo9rol0Nu4N2vs/LW9ePlT/paDYtHnIoCp
nSPt6SYY7ZksYs4KlDAv9G1oRRrof0oiiySet2xWSO/tTTsLDkxHMOWwUcbO
HDWnXqLbERTopbftzLw40hiExY0/O3R+bIAIW0NRgVDdAHCviQwJ2ZC8WOHS
1WEW4AE9DzbxAR9ZfLFWUCqw45fNN1z7+wSOJYoFqv4LREiKUuLtpuzOk5BS
x4cTSHudp4DWLsr3IpcQkt0FP9BHOEc9ZjY4GC+ydPJe+bdTI+JAVlsrEt2T
vTWwf4MOD8Z0D4opSn3D2dd8jhmw9PaiGLLhEsm5yBQVqXYaZ4kncMkr9hCJ
CpoMDWUxjmHCrLfSU/WdL6p+IteLJ4plcX/XoValA2xecS7oY1wwHYkapsu1
uFMlXXc7TPsrPBsOjtvHPr8pK5GfskoRAbGsP1yq+oORLeIc5x3pu0EwF9J/
G10pp7JNvKkQoRx2IXf/zc2HxwmI+nYiCBwnc21IQySY4qllyWd/ZmMuvTvx
W9NB6A8f9HY0PKcJg2AQmDtOQbI2smxTeEr7phJYDlEraPq/aTH/rLGy0DN+
cMXy1bGuV297Iatc9eEBoQ4MapTZ7FfemFPC/XglObegsT3/Ek/Hy6jcQO0N
VaZdoGhL5nROcixFg31V3mQBvGk1iGmayLmD99Blr165vmnrQ23VBnKcd9Te
iJB0V5sDmq8IQp/XycNFcAM2x5/2AWMxnAKV53dB4yZE1s5T90hxLT0jw1uJ
RG0r/v1PaGoTTKKNjibLnZTwitY9MncqLuD8ZtvaWwxePCZNcdacy80T3OgJ
ww6n8N5MAko0hqwg034bPcKHBzah8JvXsG+TO6WweQ+M66UxBGxBNaJ5B1R2
Jz/Q/PZaDPc/sLno9zgrl7ntar4T3KDPB1krGlcyIc89GYplsUV1ajSlEQJQ
aOlEAhoRDftcELn0GtY4oPw9DtPTEmx70Uh8i+JE4/ACqTI7daZzEhb/5s01
TKK2aEudkCmH92BfEsS+C2jHvCdOewR2EOZ4TKwogXAlqn46QPPynJRplgXH
1IG3h3fKoBrKHqsHtLKvoixuNE1sWrkFv/v1JWEWJwvh1xmR2FJNhRwyOytF
a7hutjKt5HfHYrODpFTU+trjrCS9fPj0whSgM5mdntpW1a+aFQe3FdoWezcv
mbvt82gMycUgZ77VOQKu8EOzM4aKcT1sJly+RueclQjJ3gGHYTM6CxjBRola
DqyEm+NrvIRu1rXCnxOUzHx+fBp2e7PsALYz5kbswMJUi1P9G9IFJu2hXl4n
nTU12ErXqf9S5ky9Hgu4SgkVZ56jIqxGbEuGSa95j8xnWL3XPakCVwZYSgUh
fc+RZpcZdnoVyYUaiJgwTwmb8xz9SQRkN0KZZlw0Gx/yN2R/fznVP7E/i3sW
ZNXByQWwp9bx6KfGh530DbrGfQRGwzCaqm8e9ubmHdvmOuZUnCVLD11igfVl
8TeKJtuKSqI4qsQzIiW0KvjTWoO6AxRHhdK1lhqMOA6teLZFEMa8kYBRQ2/H
cHqMWJ5vPTBivqCfR8cJcT0F0KxI7Ehj1gn73eS/6fMbhLPrPh5RXjf1Edcr
SPVTufEo6ZNKDKAj+P1E9RPMW3UDfxWhvwLw9k/C6LzpuYvKXBy2nizCwPIT
c0JqV7U0PirXRrxIqoPN4AWok2oQsdU4NFW+8yloDf1xNFhMM5ODZrumd0q+
it5PB5WQfCqMvQg3VMw/D9NYZ7n5PvXeHA6TsJPLA1KALAH6iUKSuls1NtB6
eRiMZYyW1VPBNBQlSFkt/wJPDaRlI5tLNiK30Wy98DCxPfZMHKUsjhzuanQW
djAsSSVGAqx6IPQ/Np9nch29H74OiYduffDSxGCvAjK4HYoebo6R9oSh42PG
S0jhSCMPLm+hsNhDawgG17I2FO1hixn6doXsfuhbRI7Tg8mo4rGuG9bkZLqn
6lSpetCHPLEkPmZuSTkUuVMDFK8syZA7vnzvpjETLqb93Ooxz2OqtK9LlmPK
3I9ZqYlxAku+KxDCNAQOfpVQ3dRShB/cwtRn57Jhb/QwaVSE88HmBE9V1vM3
XBXz2eyDliwYGhrotzXrhS6aCaVS/7yVmbgBn3NYM74St60AV4Y/cg/eC/FC
Z/yvi3+L08ITiLHWovynJ7MtK5BtcJs76VClMTdkdS25NkL8kiZw+Dx7gt2E
sitwWeKc5O2/cqRWg19ws/qB75QDV1cgBqkZxEJY7z+kAxhyQ9yfmX8Ye5bA
3pazLUKBoy5zEIpUP99/fAg682UV42kCgpgZ0wEaYlj/XnW/SuurrD8LnZWG
5t7ZBZbTwSUwif0zNhrd+z4HwKTmQOODKZm4bPhhPvygDYEFKxdIyhe+2xbM
OmwUIVbI/clJunzcvSgQBuqBuSd/51pVKXQyiEbDcJwearDB4zSDXcsociCB
geQSOfdXTsyDCSfDujqQYEFFfOqHPh+EC9Z/+UV7ZVHZ/NGgAKKh3+1QeueX
PqYT/BTC82nTnWRyO9ZD4ogMyNJi12zLzJal0fqblqMow+EvX6PYtFHjaFie
h0vbdAuuxpeO+IQfPfSuMt4+LjLTGvOLf4l1drXOd6PArObIrjsbDbvf2WFa
GR/vj5jxFpnwiUX+shRs38/44APh9ccgOkRik7E94h2jdNvOSTdCdZVdJsHM
zYV7swK8wta1IVxX+4shGYFbJHjVwZIQnCt2DCYXHd64eEChqVQ+6gmWagmf
FsskTKfe28bc6wwzA4gD6L0m/TVCfMInGEaLYW3/FOppnp3RovKZCvJg7D5T
FyJ8hQcVD4fgwd1BascVDf8qhKscHjDTVkXZMJifzcxRlbgdxgPoTGJivZBG
WrjXFqjCDkQ3DCDj2UCJa9vF3yxjt0rGAUboyzNpEGIapWlnBpbrWUM+RCqR
u4K0lSE0FiBD1sndVXBxu6f6O/F8DZcF6RSJHG9x67mw2hnPB98GOnekycjx
lf3xiw4eCv+AreKnIkMTpvPNfbv/fEZ+8P9sYV7HAVyTAoUI2DPZQoKBR+EV
5Oi+rSsXE82wNp40wEiYkfAkCcFQBSrR5iuDchSsPOYbyiLzZC+JbiCCARPj
Qev+aKpPVIL9sRFdMcrmhtDNTeFh/zAbqPykAUPvD3/p/6fKAV6rC2AQCk8A
LqJzySMEiCVCgyfArHAUWPbv/aaMUjhwI7rrA7ZEeF3UGeyfrJxCLwAHdMpZ
fnQ+1j+S/IDb2drkFr0oOAHBw1k/GHVc6/njHg9XDJRuXJU75gWLzU8jZhRr
esdJog5d76SXxDBYGjd2Q0L/4JnDE4th61M7DMHc+s0gmErMxv1vGpFSbOZI
p0Yx/kgSF4+buXwUfGfHrCFJWsTSU3THS4KlzS6ac94Q5Ntt6fv0YsST5ofL
SvnGUchZF2Som++r0pVRoKL/wg7Q/VCUnndTRwVnxcE/FqL/s3txxluiShlv
v3negOwwfZ05U2hzeQD3gcukjComg2ShT4rCbugtoydMvwqjC0TxH82Cuxpj
TS/2JdPfOp8J0UP0a5VDuT7NTFGRcIbvh9r69PEE+gafzlOAin0FAX4G8E7b
BttgxqwPHUH0bvpGZlO4ssvI9MX21lx7SYYcMY+gnjaOSTrJd/4ltlz0oXzO
6kz9Q07+HF+SHTcfFL6fphRLTSzIfQ9WZF2vbnENs0vkrPFJSlbsQQEFiAfY
xxCkEilwKe2NYhiOR6ZBhMHJW/9Z4To/15x+mGNhJwv2FhnVdVDYr4DUh15G
/RrzpfiLkMKX+Trtcijesmkh/TyQQsHNWFgC9IHZuJFTqG/3DGr6Leki6B6w
q41tc2EI8H+1HVsZRv/t2/cB1ErViwbd8RSrbTp+z+nBFZCaFAZ4eh8BgBlR
MHMEhDw0tsz1pLt6dDpLX+a2ckGP+Daa5uWpG44tl3U4sJ4kFhNVA+/NgXX8
lCCoN/I9+LVLcu5R9u1Y2K3i1WZkJuxjzxMkrtIkEoTHk8frleG+cJp7PskI
+dKULmxj0cge9dMyaQ/L51C9kaqrIPCaAxTDSsZp/o0eRc9wAZcwYqUYrEE6
BKAKRmTXQo+0399zWaZWCNyNKx7MHSGj4gmTsjEHHY3QL8omA4t8S8f7etqE
HtqsjI9x3Cu+5SqAODtpZkXVJQhdL8Kizp9Zhse+kr8uMOZxoj8+Zg53NIjl
W3gkkQcdG6Uqgx69UlSGFwEa6vrt4087UogL5DhgUrFYJAueUdxQ1iiL1Pl/
FQl3Nngjh8GGZmp8ZurNMWYXUMElZ7Eea105YVkxRtFhCCHQ3SV3bFg/tjfb
vuUNY0M3Magc5NWfL9WVTKBzAWXz+Qwz27jdcKh5/I++ZOcZktYOEq/M8U5E
4g2wC+vABcXohxGSzfuG+nGfopFI9RYh/3NcmvY9G65l8xbauMUB42fFiUT2
FU/RWH+yVDOPtA55b+sXAvhjlEu9+/GACWfpmTevgjah+5vyGrT9HxoDpQYp
F5l0zz/pyg2RqexIOcJdSfNp/Js9DNjQ3QklIWSy0najTkGdRpcqb0vgBYlg
iWLPqomJEGV0G4QLy4GAEfGjci53b3ke0rKL7RSaXSvaTHCFv/2AEjMICzpa
hfizVISZb/YQsvlL2xb+PJAZrK7w/oxbtsqTeTYO4E5HQCzy9tvaCWgcy8Q8
keVlMNE8nrZnmaN2ng7zjBa6EXhF96xx0RX+5msJzsCjvy111ntxs80cWnC9
WQW/7bIc9T808k4f+lXvx3LztO31x6YAUZRupKiOQGjHn6kqOFI+tlPKCYyy
M40wIOB57MDPvLkbad8UvFjDH3VgYgN8GnK/nDAGMcZ1TiGjAfxzR1jVk5C0
RJIq/uVrtN0gIY8pTmMk/FHxTr0q9bYwNuyvQNeOPQWiIHBI3rq/Yg5XEp8h
b46jQMnidT2zP+849U+Mj2qNctzo/GEMW+gUcpKi8KyomYv2uQgu0OGvnjFg
AXVVLym0UjWtWpQsudOtgFNzn+ls6pMi0NZFhJe1IdXu+Kqo+KFeKiev+l+A
4hzvLwZS+cUBMvO1fuYXfFXPScV6YbbU9YwgmcWK8m+tUpmrT0Ot06vXvZCe
8GVEQgo5wNZON3/Jp3BFBLvxYbck2ttNaCrKqIbwOM1c7IUBhIC3JGLH8VUN
ycNFoA6xPe6agZECU02ffQl5OEX+f/1lsJHIWZhtj84ybUD70SpkwYcK9r+U
EIaJm55d+BcisYMfDLyk7QBtf0xzLYrhTrmc5OFfhXcvSlVyXVmqUJfCcL1w
hlYm7ZwCcekTZSIBiQo/pAJs+Rmt40VAGaaACIjTT0UU1SkeSVaGTpmBtdJb
l4m/dH6HHqXpxlWC+YGbKCZvS14+p4w0K9JatqeUWo9sS0SQHFLhRXG/2Ww4
mbecKDg2PZWkieXU+hu2NLGCd5goRMEvnQ1BMNNuzdnRmJVThhOCJ0UM/nPB
d8pKT9E/Fqbp9xMNe5Y0jZDRmyzznFF5pMl3kVtYtOgdrNEE3iS0DHRXcL+M
03k8C5pNveuGUporvwdJN29K1TanzyVfapkcBPzpXI51qiXEfTsRyEjPvcaG
clj2GQb1sVu9vsOPfsjaIwfGonjfLbFEjpLfvbp22Db1fkkCbcVq4wmaXJK4
3LR1HFTrTMZvf4J+IIhjl+CmPx07QyunAZbvqEQGhNy+3gsbKLYE85eurn62
IZDgkwYB6kxOJx44jxo4RoAcMt9GYNKZwqmBIQqhsybHuMCSaebqtump4R0x
VGt/3JiUXKzGaVzzw763f7vDGnqvrvD+mkbJnqqUMhFN6HHvJjMtCtP3SNKN
pgwQcfkj51KlwM6ooI5nId08zQ9v2N5ACX0fDBGDjFvDPS1KDFO8S38bCr2X
MLBecmvqAUaFZIzqA6Hx0zMkUBMMENi5I/uAiNDEkqvE5MoQQQtfK/UdSCMi
tJiQOKDOuGgewGoCmCCPDdnTmsVUm92Rs8x1MXyIuG03rTpeDvU6h34f/JQS
HhrWOD+jqWV7TSUDOQA+WdiOLHdfXX/gx607/QYIuVcn3DlzD/zz/jrQRiOF
8bKZJ0Efc42Ng4sG8dIkrv8L+gaSA72nzTx7GhOjIYp71oEH0KkG28dgVI22
FTKeWZk7VeQx9LLZrh16nGyYsiYBcC6rNjqtC2oS1eEj5nYiMf3pZRFFvMHf
WnDRP/+QfRxs3wb9/rJAEV2XVOoE6ltKXQc06AuxffVLsfKhVIJvBFQDvkpq
dGACWWIgWZtxnWV7S/fXU+Ab97phL5uIpTx5pZtalaKYedo1hMjjBH8vQcBk
sIxId84Rx7ohQ8m7TQTTJlG11nBTZZDejbxaut66zU8Fj/9yKFeujcYPynqi
6H9RwHux79fZhzOUwHRV4zuf+oMX+P0YiH8Wh1fw0piN0vCJ0PrLumE3BPQv
UAZNiXQeuXPfKPd3baSZmk6afKKH7C/jfxzYn00MOQP4SFzwjmJushcTzKDg
csBYR5jVRcN2UNAx20UdoSg8dNNG/9G7EyL8V6aFXepubge2jZaFFRP69q5g
bLTzoAG4eAMQHNFYAFwTKxtPmfOlnvxBDbTzApK12p99xY4Y4OU5QdWKp2N0
vZRlJebpiogTcx3TxsGpQxhg+WPIPpYArHXvGKOUF/9KgGuPFclRvZyuNFsd
8TrhwuLgaE3QeMMlJ0wWvt/8RRHcZ5ix6/NKYo3+JUT252FiuQEkMdQ+/wH+
GRThPQ1AqVGnbnCCnecEokH0pGDfwWs13rrtNeOMfbSjC50NgUDpZ7rHqZra
yz2JcrYOsl6AE18LoV4HbjIHDTA5zw4HKKQ4ivs10nKjR13ghmyXnvaIoOC/
aGrezdVl5lWal1c0xc5rAFNrF39lqxozoSedm8YDykHcOddtqZuSnXeYR/D1
0zxKkUadGtaO9MmVPgMZ5d9LBfsHVbC75uYVeaG6aDlMYTkC/cZVfoVnXoCO
bJxp9mDG+HGYoXBcliYls15UiKFPXIhuOKXFhlU3i1DmwVpsG77Sn+P9E2WV
yG3zcgHM5odHkvq8Zv4MD2FzCL5IBbMcM93gv2DxgWga4LcII0RPgrWTgzbe
vtUt+zF6N2PhvWlKRGjcJJ5mN9Yyt+r5bLMRJJDtoWYoP0m/uqtzY93SN4gT
ocuTfaO3cSFIwmsH6z7/iMdoHUi/S7CmuVrukD7pObwpcJKqxXHPOXSYu5DC
0ZMqIFHZCoE5mzFd076vgS8BgGfJiJsHzcUFBOKlEL7YftVr5WAxjyjAmnpC
fwyK6xise/TMjCQUfqpdp8gMO4SEeFmY/EedQcX7QmkrZZ4suD4uqgKEAtDJ
OIW2EOOllfMO1l0a+WeP4w5+6ywQX7eW+3jnkx6TyDMJPfVX0Qsu8hlrokGw
dbRq0s0T3K/v8yjo2j4haVAnOEC99Noho9KSZWIbDS8Dw82AR2Pr0cXXTdyO
LCk5VJ9bF41Ax/Jw+gJadInCyDnDm3HwTzhWJw3H2Y/sipqXJdwqjTQXVky0
WsfNxfqEdSuc2bXh8wa0u117LM/8co/bu4+nNdm/25DuxCl51kZAO9HAcgdB
b2TVzWvacrMN9S3NREKDcupTLM4QncxJDrBQyDT1ORpHYYstdTJXZv4xoy9G
8ktDZrkb8DRPdIiKpy9tkFYeR33SWQGP9iTSqQaJSAJogapAsqYMQ3cgYf0w
qwFsEFW4YJWNfz79tnjX5vaYIZ/q72s6hdsV3Ru0ePeacUB1hYmYAY0wQbv5
ctU2avoUMsXwgbA6z8vz37b5h2h2W2Tsh5DybGv0AvhHnH9nVMlSBrDUDKXl
Msi6YD0kHyFQuWI69inUajJi2T3wqacQRfHFLGTKBkLrMl42xn9arLVBF0Rr
ZNPeypRmeylBK++9uchygKss9Omr/jnlwnL1LnkGLEIc2d027Avqjiwf8+QU
0usLg+i37jl/AKRnj7m8+8P7g+zwByZrc0r5+vWyyJzBuh30nQJhjGzuuoKT
dhnN/nEKLAICFQkcvL6cSz14sxPYMJUGR0F7t9EFE8KsRvoV1KkGuRkiJdT6
zHA3/hhPEhFQ/rOuzMDUEGcImxT4NYHOeOOcb0MLuNiA00GEEvFwJmTO8yDl
P7bPDC15zLvi026hZbKiRGUl80QHf9ELqJGSKBxzXJW4FfAXR0AIOfJfxuId
/PraI0zOljg7S711n3RDqgMM2fQUZYyCAQ5SeqTBltgsTaRsQ4Nm4v1dccdP
ZygZSTwVkyEAd1pRgSrATauYVWlTZOcMBPu83f+8WTWoVohqk+thLvwEJmqy
pdycoazyT+7Wd1681kBWkdIoXItiVcXhTfSG4/N6UVmeN0G255pFUKj70ZLY
AYit9263+09NiRPrKywkdGn+nLbl2YHuiZLcU5ir6l94tugSXuLpQSGATkQq
zQOtSbXY32BY0Nh+sjWTealZ+e3/rGEQUaeumHD26mCT2bL4Wkp9Nfh0Qxuc
1c6YdS0uwUm0uEdulMGHYy3+4VWvYdHS+9G+kQj6Mm23WERv2ETKv3YI0y5t
qMXO2Q6eio28jdWaT8v+YM3itD+7rgsNCVQGy6sIxIrCBd7N9EBxuQXjbYm2
iO+EVvOCJrA2QZ5s50mh+Z5+t1TkE4/76pVPUDCPq1fUmpIpksDUsBtBSoxu
12p7lGNlPGYdNw98XOdQgRkJGeYsCPxQMtwQl0lTPtSNN6/9LEb32/Dqdyfo
HoJKSxwgFw+r3QruX8whQqkHXbJUiqe8lUt76zmDNouY4Iy1/sDZUaByYw6/
hJqz6eIu4iPAVT0o+T8MTjgyN2aKvWv9MDel8RkP0wkXyEF/37Zzc5vYABvb
oRS0SFcuNGr2+itMrezJIsB3v1WRJ1TkZa4fO1jY4UhzumnuOfRiPZZxbyX9
3pAEhFo27OL7q5KhE7sWmOI2uVQtZ9NjDQRIIii0IlIhht1Efb//u1kckGg6
zhzTe+efeXBSAjyPE23GP2+RCXFv0tlbdEYM0ydLlROlLdmj3rXGUkBhqzkg
I9oSlp8BFDtCJxOijN6a23TD9Y8ReH2xZH2UbEEDIcsoc15WQTKJMirgYE50
c5owixOvlPzKi2LthR5WVRsEhhns170C8mc/5RGQG8quxy2NXwM7BJMKcHF/
KCggeGSOP7Jt3o3G7Ln6UtRVh8oNVIW2cWYvdfkw2LxFosF76Mey+E5Iy/zL
SJvPa9N9TjuAas8iVv2ygcZV+0dEBxIxu+RgxMPbFUbcwutY2E/UW4UCicdh
g3sJz5LnYua83kEMjcIUis50GsPAIo5P5+8ZFq7jSYgcY70+MYUb0Ny1EYBs
ggcaxVGeGdf7cMBpEOwvzCCNYTvBBfvC6vQi6QEBJ8WjKeUcLenUXJAMqxzB
cV+8ESAMsIG6EwXA7FZqPISElnJvwfjXlT22EQy4j2mkWTfd1SnsM7XdHMU7
2N01eiT010giQwWIoD2o0PN13X0ccfjZisqZssbgM5OiLWBTT1E2F+n65XO2
8pFQTJFsdO1AgOpxu1r26dLNu9jPsQ7iQjoxTC1dtbq85yZ7y56KCpn0kRi8
nRL0/2HHPGaU0DXlsZpHzXcWSRx6ECZGB6Mn4Wj0zTfP1/W5KXqwiaIo/gjU
9XJSatllHyh7Lv5658BiVpIWg1xTfl7QvTTC2kb3jHUX9v0Z6gOhub4M0TxK
zFm8+AbT/xkJt58US2PnJ1tnMhRvSdsONWeax9IpGl8sFMb4jeiqIGcnNARf
7TZS1hK1VUBZ5qvgAVinXjAAwlP7awbMr+u7UHg5T5vOcyGyU8NiDl3wd2Zw
Ry954VtQJXrMNL9XwHjbCnDGihje3V4G7+Vq+U9YJYHXEdG1cTj5qEGV4jog
75bPJFAnP+jkong4hFRoVdW40HDPjvF+x6OHgiGYTmcVz/pwsh6jBnlbQRBG
ghfp6UsMWSMCY5zlhhInVrq/tQEJ549yAMsFU02VJOQJpAwWEWXPbIzOlqCx
gahPEV0Z2Mm64ETGdhupxUhE40CWHroG5gX0b+VdB8+fCvWl0D/uhgTxe9r5
yUxrzzLFrhYwwcEq4C/2bi09NmM2abzOEA4w+b2sP3JsL0db3rC8bsTGvtMH
eR8UdZB+qK3yDxwWMZAU4wcZ+Omq4iMoLbRU+us0WaHLJhL5MLVOv7Z/KirZ
xFHVoJxEO6Ro6tnWse8Kec4FQWqdozshu5yIP7KY2hCnr4Tx9ZZFYIQXSvhu
IVcpWkBYQwWMQU5dMn3ouivxtjmvWxsFjM7D4luIbgb9fpo8ouni8ME62BFh
qv7abUmjTS/1myytQSszP/DGSuX4MDrHLH+oXJDU1HK871l/7ZoYwdktV74D
LUvYPCmu2xMdw63I1iwD/q1AP5hcOvSb8JlXsxApog8m5Uf76WV+HbUGcluc
VF8SYRnpqR4nSJhqADYqWJCQlfBZBK5+tcDQELY0NxblfxzS1w+g0643N3+3
7lkWIeqmTiQAALAwqEeZfvgq1Os0V1RfA6+Eisbli8RHA1k4UYcIHuXAZU+/
zkLcDypNXP+tNCeOOnP5N8VkplfyaOLj3UCaJBsgHwhSezwHPWaY6gzCZdHb
y78byBnHCOnQnAGnGxOgzBd33UU2YcHmnDQ2pXKesd46HfBiF0Tjay+h+++e
ixhig6HuHULzzdZLV9r9ADQMFmCUvdUdBaHQCjZspz0Gc6aC0LzNHwNbs2d/
o9eV5v3nu9ngYMlRJz8/vv47kRGlmsVGIkZSzRUY8s5xpqyzebq2B9Gi6yv3
zkgibn/6kZHR0JLZG3FKrit8WmpJtCJJjoINJJKskINpksc0TuSS5tTLP8QQ
xLPTYyQ5D43txM4D6XKaBpYFktAwTta7e62fjbb8vO5QEsoqjH1Ywbwpst6R
OU41cH0ywHrhE4j9uRAqB+MhtahU7Ji4D+pils2QYVzIvOy2vovQ753Hpm1+
7ef6PVfIkQC+XCJ6Aty2UO2KXO6XZUjU1LupScb7pI+vEteIRIlzSCCyGY+B
iD2qtzU0sgEmsy8bFY/vDhfvWUl54O/AsOtVqYD3pFOkvtBvVVOZfk+0Uujk
UAZDq+jyLZiTWPG1+eCgYF6bmS0r6nHTrlQwQs/4vB+OZ8qV663bLocLjmUa
mEUjNTbqlyuYTmGh8ywfkec0onTqFCZReeqlgvd8mQyzPvG8LLsYMtPfw/Za
BlnmxmnS4hpAu+SMZqQ60LLvbgqgPaW/6aUJcJsg/jrIuLF5IGZUVJ4+Uxeh
zbfwlTNR4c7Jri2cwLNvQvbRmLSAShFPbdJBCGc+lmV99VNRzPG+4LpcW8Gl
BI9AQ5PvenZa5BAOYe+OU2W7p/qh4T2aKan8qoUvVwEmBedoD2g4XkSrR51z
GEynRcHXdoBr4+YzjZVR3jCPqzZXD5JLc+jXQvXCwOB9fb6WRVa/8bGveOIh
x4aZuqWUyHpVtiR1ITpC4hp+TSFm9HEXbT6QeE2jVVAvkGis/g3xpHQtZzUu
9+U5cCZx9MlwEx6FUnmILN+rWkQ17lKJs406AkuBT4n6qynhCfp4rPQW/0U6
CpWkFrb9X1WsSURCb8T8FQLGiyphEo3nOiDLxOpVozPDucaOHnn5wmzsePxz
IhSQ3niPkr6nytiK7N6eMjAfmK8K/RsIWp+sXL9MMEfKEBN8DoTFXuPqHCH3
dm9ZE2mldVQcw4AhburfQxpKOveicT6GyKwDDEIXQZZ/klChlW6l2JJzNWT1
QBMvvY5Fz8D6rSUfDtS7d3oCskwYkmqVy+kLZVIcnoHXOJJF+8rh/Hvx47p9
PFVlaashZDi35h5/LHz2Ze6yn0iWY+GMoy6ky9KZoLigbbSvfpEge4xV7WEx
IrueJ5PIzMutCapewHvmjkYmcOM8nc1KxVxJK1FWZkQ7f1zNdgyfIoTA94YQ
d1rKEPKcBCmxVvlKVSX5i/TnDzRunuIDBpaN9Oc17e84i3tp1hVQPhBg2fdd
zFeidMtsL5oC9745aqcAhiVue6sMFfARMqTt2tWA9HI8d5+TBPzwS+r3Q+3X
9pFOCneHLBZOn9CMnirhHTnfJ2YmUBTJfsliD5HIvTrJM1WhKjB3+9odRUDo
+86k0FUJHZrPXZaa0DHU1Cei6GGSB4dCurPxdvfMrtpb4S7ad9NkqTqDm6u3
lWh8VdyhFXCL569b9TfwWsPA7VVpJ1rHhKM0Nc70wRLpEwfnRyF1cilBYtNM
wzgdZ+dF1h12EiGeIOXMkSVIXVja+Dk9nHgMFEmRxg46dItndqnmj729tHtQ
Kd2x0JJMxcBGnZNiH0Sezi4hVQqaI+RbdcLjysoOd+NBVkKDiGPMqfaANBkR
kyf+r7HMR80ybkr1RnGgcJr4F0W1RN+RkDiogMrOOUxpUPwcnS7xVjBG8mhy
gLiBjtVCbYOdyiVxW6RszMdOQB1gAVZaTsFVwz4qt48VRl2l8NT78OVohlF5
rwduUqY3fl8FOiSUhmqn9AVT4DJ7jhRQItpThCa2jY9UR314Uzc3ujTZupoX
/PqS6KfBqCMJmk7kw+Hbomt4sunVtjSCvDaQ3Wt5OlYpZlZ2lesA0faJIg1L
z5qaQqAKOZQsTUQkj0s/VogLqnu8AWYkuwGjPyGCglGdb/OLjQoZXJ/CRBrw
LOC64AXz9AZkaZPWJAal///HqL9yCPzDiM6D3oeWNnqQ5RBeGodInAwv/HhT
QRVqhzOsjDhZVB9nm8Obyw/OmYY8v191D0EDnzK6ofBWk9n+6fcBcu0ASbyK
1mfohGDmrgCsoqytHeLmoDjSaqhQRu3b967ChJmxkXkzSfPxwtDrfPMOYztb
Zwd9RF+xy2yH2bH66VKC+dhyp1MKq0RcsKEkR2+JwRYCYoLReAjWuS4lsY6e
t1iO7gwShqc7iGiF69fCwqBaQhS39EavlNsjp5FveL62OTw9TUv2hzGNaCYj
RWXM9CJ0CTRTvFpHSYoHHfdqiMVv/zUdD1Z9uULM1mXlwrXMt/S5GUjLrkCf
VrCUvJRyK6aJmbDhCyzgdh8LogzFdlwMpKZS11xWvlRFhQ2MXKtZ6XDyCihk
zZtM2nR+MeCnDWsBvGwCLT4RWucpYqn5NOZsHEBYzZVWmuCPI4LxlqPyWPAX
uPQx4IpWsBeQMJXAU4kcxh8inpyBu9L2fYdjmdHf5yprFk6DW0Kq3kwLM3xf
1qe5JG4fAk3Hv/UO5rzDG1Ot+5/lZVHRA/QE/SCurcwGiLXhq4ZmBsbEoFVC
S+o1RJUJIzoIujqOV5v82lUZrhlAXPZWOA2Z1qRIm4DCjxjA4Q2B7ZEOJldH
171Gqi6r4gMHoS2Bwuihr11qZJ4G5wOEzyssLlqWPV/W+/H5oEGJx9fpU4Uk
DD6vjQEh539qCxzoc0aP3xOdk46TnuFYdPuwVH+2R2/Sx4cAmG2DyGwq68zr
SxNhkn2tBUuVVRxSlD/a9WGk/UhkRNmj3PPddTqW52Bt1Ve7PhozRSzri9t+
SExReZYRvejB7QHSr9K0x14xYk2X49nJFW1bIW1YMboFD5s35EYlrduIQrDW
LO5AIGpDWM+IjswNDE4cySIvQ132UDfndd3bCnHdyjdMHmyuUKL+3ph1k7Rd
WYR3BAUhqrCn7yPol21Y2VzadUYweNHxC/bRXYgUnjaXEEHrxachdba5NxdE
QbEOBmXWkYESkxZq9lvuW2j8GBaYI/LrMHpm8Oe89IrW+tsMWInILKdTC6LG
YcKasRkGur5+9aL/yvmAmmorws8xfo3eJlQv7WRbhfVXX3d5jLEKT75qRjjf
p3sHklMBap+vPLGw4fqglbFutrHzzwsnwhmSk6xbVKWZ4L/ptpWTD2YuV7Vi
//xVUkLL2Au6TdcgI/lmb4F6yAwv2Op6Ro72YAfPThB2JAuWzlvJsnYoZl0i
wlB0sT1veKvyRVJP2wTGOwKerLS8iCKHUduaswdunDepO/JRe68fYPk6lqsR
aBgwdgJwSILPAAYgouqmF2Nt4jF/0qaT2oPb7I1A4xpUZNs7h8ziJ8S+MmmO
fg5XKeJxuMDSMwz6X6xddUqy2lqDv7Mjv8mMrFMtZAgayJkOKivVt701hSw0
VDYbR1tm+u0XhohXvW38P9KxJxDIOJNX/LEkJTr/J8gsaVU0mebvZS8Z7X2L
p/c3m6WjNbyJf4tF0uRVzRqrLxebzPqWliaU0QMtzCzHN+3Amvg3L3ILkWWs
wy93yhHz4W8BIdbXUWvBymroC6FPEAvHh3MqpadpAgBqCUxaW7N97hQzz/sT
wgZ+s4/hfTSiHTpFENYWtsfjWLU1WIX1zn9PNCKokae0ZSZS5qqNAAG2/kas
MHLuu8bj0VO7arYca+IngJh6jYFEKRthg2/z9cvWeMGGnHWGbOB8IcKRkguq
ailq6T4L0FVgXow9gcpwhJxQDsRKz7yYueTN1AOvDBebJL7q7SGD5wxGuIlT
yvdoRVR/MatwR2l0vyPzU8j0FjvOXJ51KhMHZGGworMEC9/EPVxUNrqqAK92
IpYbU2kVujrPsRTEwZnZa2yYT0wgz/8G7JNA22qA4LTVhB5SjFBSD14QYttj
rcSYfX/DpNwNhWnfHwstx57GUAMKQvRAEVUmKJyQT8wtYJO0/EkjaIrSVqG6
muoRQfaLKfhC97NSDhxT6wAysqJ4rT6PQwU+onTLbaloTxvF4DI7HITizxhZ
+ugRzs5Mi6x3s0AW8cADQK71YpSQCfo3z/sZ/OhxwGF3e0lsdhbgSnE0qFUG
1eWyr4+efIVKFcwybD63Suw1IzSzPQ4UbHTGaoXk4m5vWZbX9HCwllqc3xmK
vZwmUGEn3CWOnxR+QFat0GjqRzTsJGTQ1x7iPSYIPDjxCKaMkA7eAcqTSBGC
FWEQKVCl8XPz0Ie9JhxLSmErJo0RUA4RAwWEXZKRaGP7jkFEhTSm822347qj
0id10xYHiE7UQ/OaTUxVqYpmGgip//zr95Ui2NyO8x36rcMFKJpiuNiwQAzy
1L3SV9aJY9oowojZMJ/Zv+E+g7LMvKqLOc1u2LQqgWaBOxfVBs8jP9nEntyU
60VueC02tMJ2B/KA78LtUDTShcVq5kS2ZzHGYEpIh6/BBYEx7//j1p8qlo1j
1bP7MLvsxGp03w0AR/fmYzAHTqtIwFcSv/skif+JTuLfjqablMePhuh4Jdik
5k3fAtLFLAtId62ZD1o/MnjyyGp4lgokGtjzUfUpQfALWnv9b++OzG7mOlrK
+s9XFAkCSEk5bwcBJBoH9oiNyANdqC7oIMyl+54K1dRVeqQLzF/uwFSI+kJo
E6jt+t0AB1q36FQvRM0uxavowiZzxR7uiVJQG/KLj71nym7v0wVouRFaLG//
2bp8xGRSSIyYxfnx7M8flZKrSjZXEqoMEiKkI4P1OapVr2H3Rr88aJxYP7GQ
REPVG2rFA1MXJDpfUTNAh+8w3CDcAZDXpE2/T718tTUkpDO4uXdGlxusH3Vc
udzBuUqMUfFGE2YcJkAJe82P89rWiEPf872HBe41TmjRapR7a29H6ZT89RIO
DVQ4CivCm34tadynK819nfCD83Nr34JT9uKsEwrt/b5GG6C9HHS4UeCIAUlS
pZKnv5V+JH/6rtbiq3uJPpvf23IfOwYq1ZawI+I1aa/XjukQAi2LQf6xIWSi
vAnzhlX7Y0UCaUOSvwp6aMDUrORYUblw5OQKaoxMsi+5/E7HsThzXHs5jUEK
L/ceqAwRSGSf9gg/cCEEm/71zBDiwi5kT3r6xgp04FPEP3tehHAo77MEGsva
0kt7dlg6yz6IaNHth4phsUNU2vzYGLO1GLjX6ektPLgo3irxiEbpQ6trXJWo
9Kr/8Tnry/HP4iJkE1NqmIo4YySHf1TI17IFA858ml6eg6yFO+tHo2dl+TGp
VGCyRLMU9iwMqEoTaScZnIRZ9pRED6G+xus378znemqG98Hnjwy+Rdo//egP
KR9+A8y+3nKi//vL49Z/ML5PqSoB+aUGnWQuooKxVX610YkSLQjEBzQ81omb
/1WeEUke17I5PN2ZNPPBPvLyD4irdO0mzqsJG4dYBUzuByKifWPlc21lQTf2
lmHHXYw2SwPeaMduX7C73NsPpivlouWiets3391JJPCLH0AS5BbFBSlYleNJ
0SByv1wqc0X/GP3wnm0gd2pxst6llqSrEk1+Bi6+CEscbucm2bWwRLdfr5nr
/kBjc/FACf9UlCATKVwljpMXFc+SX+pCFsbM4vkzpYrBLf5ZI5xs9vVBuYVT
yNx71xQHORJMnTdPlUGXJfjd+SBI4JJnKdeeXNfgOQ+WTXJNfaLQFv6zg2xK
7n75UTOKYP+PS3HRPqC9KXMnpT0NBKlNulgJQdpRpe+WBA/Re7WbWgagjeeS
0ZiKg74g5dFOXzdKu0MJPhIpV2wZM6v2MgxHj6ovC4g9NpqFypvQjLJooi66
gLh7j8mPqPyvnKg33mk6ElK/On3Do1QTjxUR7mEabu4ZU9mh6rwFIWXzlfTr
yWAor1n9urdWRCokE+VtuknKz2ajXaFecWUNg1aXvrWVsPkU3Ucbx3F88fM0
2MT3MIbGorNr9l3CSocR3U/USUzFbj0W7+JcLlQelJaxExuVahTQWsEiMSyq
Jhe5C6n61bv59q+Ir5ntTV1XwW37+yaUErSn93+FAaJqnAiSgYwRKtNnGl0l
YIwuCOob1DXn8PUYEFVndFi1ijuoCIF+nEDbfo5MZMkB71PA9dpxleqyAFjL
fo4iXo0dEqXo/5QfFRNvdrXqJ53fuRtuAZHpkMIefbFOMElC7qKkuI+qp5qd
6mejs4nibx0bl9aGhQbXLzBwi6iKjjJCmrydHWvgASrds3/ZqRW1FxBObCVa
X4b/bG9/YKn7n+8e3ESYZSl97jqxG0bmD4I0uUsLFjJmZSLYLT+LBAyHj3lf
lD1D4zbjTIY0C7zkCnpNrw1IC96QYz+zH3EvDwUyKKnUJGXtxUGioNetnME7
K+1omICHVEAuFT7dvEOVylW5VstHe6lmC9CtyDhDksaElc49NIEDU+IVf2bJ
2yKpVT3i267LjgfPQ9AUMyUV793J67981AdlkshedLhMV3SJ0c4Q8+Jou0Vz
WBrKfe74QtqB3rSnoxol6kikqF6uEUN5XfqWVPcAWdSZgqTph0sqHEYrVs4V
pc0vpcwcX5m8m9WoXAKIVOhPGOPgn+KDbdJtl84rE6IQG0mXaIuI0HK03cQs
V0yNPo6nrnINnkDxizX4MCpKXFK/nDcKr3nRPeBwbiWJvf8gcWdSA+DJ7adt
qaTiD35DSeO218XFCzkwAo3wk1eknvG1RdwySDKFxaYR04pAejGuFEcYi/SI
vnDH/oyiWHmgMmiPKggeNmhIJTNtIvk2NFESOLQzBNJ/TuPoOoj91e20RUdP
vFE4ZxN0Hp2kwCYDYjAKP9N3Jh/JxHl+SaKUujd5sqYEIp5XZqhyZWnyHVt1
jVrZRUNgHJ5mje0Eu07Cc7HwzJPR8HqGLyCaWraR5z3aY26j9kXnkkG7evQe
PLJbTdK58+UzE60eC2tOZWXCoy8PpgUzkUzY5ecSOFktzrnCbjaekvCjyNZi
aM8os8+REiOshq1SUcGLWCqgsH1JK86WiXNCjuRPa9ZB2/fQclbYrfXPM3kE
yVMlpC8nU+UG33dYGPRaXj5ejJH/j5OwxRkR6yOrJ8ObR+neSoLVbSEqoAP6
p2QixWcT6pzCUy3887268NsG8XehrJhewopsRJ/Zra0DT1M+RWmMwCc5tniQ
WDONeNqtLM14qy1EnEUbPbFxXt8aiem0TdXHggCzH5P8BPNLdq+4+lrx1UZl
g19D6iSln75IxG2hQFoDjJ3tb7bZSnaGZT/YJQ127YCqRg1++RqZ8Lpwb1RY
pBLT8liim7+OvmQXyI0FfWPumIc/Z6ZsX2fYO9+jFZRy/be15XWoJsZ0eYOv
hXIavM+0fT29N4URJHPS0pZdkQ7j42mjvMgdOiwIFb5xteBWsY73ngqzyetD
zuKVo3kL5KFy6HH0r4clMn0bTiFZUvKuqOfsmt5hU5+1PeiDWUofA7qgDRMo
vbzqfoEvdyht/aa0BodniRQjooWAI1B2jVxUxzWC/1p8AKXN8FIeWLNRdP8+
xoYqVv4vy+5FvP1da2RhF2Y2KwvsfCNXSGhVb5M9dbH7N/NL76qsXxlrTI+J
Ni64iG48jjYvlFuKJv2HeMc8d5rnUZFkd0I7ZDWoB8TIHbEcbna2+aQ/w70f
Xu5Yu9T9euVUCu+wku16+60WCRM1TW7cefduzTROSL7v234lGt7eiGajH9Wq
HQ0dwk+GQAqoCEWGgnfFRoAN/wVMDx2+AyXxRna+1/qKJtt0ovDGWIGAFChO
zKSYEzJRZ+lAWCVZ5vqti8JMfQkucsX88amkwbxn5g3UITPOUH3nwc6wYm83
ULIpYXZ3wmp7509ErrRPw5Tl8ffhJDfvaFJ0Jf7xc7+SesqilZ76ugQx6hXV
/HxxO3JKBfT1YL4EDCPDGvqgtvoXKIfj4VPFnOYoeOnoLXDruKyr0AjlCRgS
6jJ0l7VC+1Kx2Pjobf76VvER0wlS/56xsu4JKMnhtb2UEqxGqkQeaURIrvgy
A/jJUBgCGXOCPXJtMzKzLjeb4LNyDC979NfkyjNZBabghyPbZ7/9i/WiztnQ
P7pzaMTFKr9l2vjRuc1NfCu/qAiH/oIXAoNSDW+CEhIOPj941q17jQtMdFR6
AfnWhx1fOezALykKYUtQnDaepH5TBjSMH3Oz+Rdoc+MpygqK9FFgnDzw5N2X
/8YiI4Jm0JOdCZ+fmKQOzyHxlJePqvdTecCwYboiNtvjdbI4u/GCW1Kuz+Ok
6Pbkvrpa3vJN8XJ78QpITCEucTf/cczrELgL19abbnQcPySR63OBMehccRNH
Y6VBkgbKFmHZudnbUmEGQgFrwg0XHg0S2Wil4UtshUGgpUrthpcTJotqnBLl
x4zCMDhNSAcbvd5mGti7aN2z5pQEJcWgkqIojvc2Rv37sUzmhtQJT9A2MHgr
0fUbEGodEG9bYKClYHuRaXgPyE23fod/lASVsXvBHPitz85I3tvoPGSOCVLJ
0o4T7+MLEHz+whiaE3MdGKqR4WEJHRHRswuXhdWxccE0AG3AkNL5imEhuIHm
IwabzNWL7qzvcr4DchHRjS3l14+yrMn8O0nx+nD1ZAShwfOH2fEVu2HZ+eif
QtSVnt2Dkvr7AD6GAJ3acpspQmCprSL5CV3BgkeY8gpgLki2rr1Zy/sJ1vcs
6AEQZukKmolf1Z775D99C7JOy3KrPQOC7A/klKdwWwSOxKUsw7rkc5dEJnRc
0O1Z1+zZC4zK41EOVF+wb5Op8bMNvLrOOZeeTKU5r2DyLcklUUbUUjsbWYId
ii4PWfIeuevSmj/uRmxmGmGzQLvFsk1urcjBrzbyGwhs89xyVM3I6VrytL5g
+3tb+m6BjLxDKdwLyiHT1QaaxnJDruTbuwaZItd31BcFq2W2kyR5BKIRDeMx
sl6PoTNdp8rVyhqgeWrYvRozYDjWkpnJDhvOCsbNutDl6F9HXq7HwHZuWo93
QIFExhHKD6YC5f9c8eB3akOXCPQrMfvOLRrOoqoVf1UnmsPBozip5cVLz+5C
m/qZtYkUBfL0B+6MaTw1jUkJC6HAWwtDXbED3whjvaHm2117bpnwU3wchVpZ
JQ2KVSduLw26qGp9nKlE8beVMHKNUFR6/eF0auNa2//+h50ja7r/D1M8A24j
70KNbdVoitwK6TPaICxzkmumd8FlqxTDcJmvMEsrKaKeQ6hhWewCfMPyRYXh
KZ3zc3r93CxNg5Co/SKEhR6ZajO3ZoBYJHyllYcuyvUR32zoqAxUWZd5cFzL
WE0aG54P+gqUgawcgRAp5Z9eumGxknvWiISfHTW5DmYPRlARPP5tTMser7Fk
WlCp+ojla2+z6Hy5h8pkKuNx2lRZgCQqutipU71p3VTs3pPtHWzq4UAjTM7Q
54HjFUkCteLLqQQqOWo9sr6rXC2lQMJv8L20HRZn/8eMj77VaaPH0NEqxwYv
qRhecV1FSXWHlmim9iMLt4C7xV9cuXxaLM+GnSBHX+EanBj3am0mYdm7K8NM
ojgxNARpuVPprK5iVPqEIU9rI8XhKaNl0KTG4CnrTna3UAl1eWJc8kOegkRH
y+tW/uRXsm02K5vxWWe8SxMJes6euUraNL6cDmZOP5upXd/pQU7umgYAIYKR
2bjEBSIdEZ/SsFXB1uRyZZ1Dz7IW3bO6Tkd1Q5VxjWUPSJ/WEWFeRmVO3MhQ
q6JKARx2R5hG1/4MYkg4ngL660VGrIT7uAIqE+PRgPS2P9oOCk6Di+pF4mps
nLZJuIOBTLQhI2stXoA0nHCOyoWmUgk7y/mSNjI8AWSeCDVR0nutl8+wqkmD
GiqTuW3AxxeC5YFczZdqTgs9qX54qdT0KlXT3tkfjFfv9mmuAAwPyC1at+Gn
PEM7QOMMdRSWWukHLe67+n+J3O/Hq2THJ9yIrOwU0igH0IB9pAosPbNT8zn0
1Q5L3FC5zHJqK8JBJnMgxcv4r508MGlUxjXARuHO47MERJX1lTZ1ESBsuUbS
/1j40X1YvzVd8L5+3RPGqlUGr9nMyrSSTq9BGLRMsoXXNHOv9B9EY4w+lsO6
0Ij9caC7KhBgIB3lWCqs3F1qO7vrSX+d3OUkFG/RY7ifjZKxJw/gJWuulhFq
wMSxYR1IF2OZCUS5SNP2ACc6YtHTIYCH9fICEYZ7tFh5MIqUO4D5Yf/ODcTJ
+7WINFjXwA3NiB4XciluDlOa/4Iwt4fwPaXz+QvZfaLwSTO0E1TR9eWgCWhm
oiv6sP/61T8uSG4l6h8+4RuxIJejMvkiop/1yQWmUXERJ0crOdc03yFquoHO
twITKh24+Q+y47CXk5+Ra8fhN6rQEceE8KaKtkdQeQlM8tg0+7AE1U2safkj
EUd4vlo0QFD2v6b7lej+yTma0jrjZ1L00Z939gV8sh9u4DYltjTCnqbyuzB9
t7m5UpIajCVeZyjRYVCtrYXTExVR+2xY3AZZZ6lRtjFHJdQtqFX/nYUqMtG6
YBXGwkew0D12cEqpr6PNqzrKFc2a7JvwvBzyuoHs/AJ6nDJ7PcID18jVwf4i
wNi6S8iLFz7pLQsxzRNqLIScgcgQocS3ueFQqMgBRArX9KBr3N0jdDi/mf0J
q6ly90YwARriV7B/4gSVyWzLn8UzbGee2k744x3eta4F2BR/4iRe4HTCoIGy
pbpkbEbneKxMxs6K8igBVRsoAB/HQcBAdnNU9IpePGdq6LhJN6RQz9IlL7xF
1sxNKLlqeBczGn1GQ6Ii+6BvGToylhQLF9NvFuV3GG/kbX2sSHIjCLnnAKzW
IcvQ4Ff6YTJkr5TctK9wRpDiCzP1hcj7n6N6nKGuN7PSN7P0MeH20J8zyQ+3
Met1t9boa7GRTGuIEz+6RbTwGXe0UsoATbFBHT9PucflCLnI63z40G0KM0m0
WiGpuqJpHZkcsuWOsRcjYo/fF9kYOWKgfBCcijxUhZy05V0q3xTHEWWoOT3T
0xq50V69al5j0o1ewoW9C0lRqYKGEVOMM5CW7SWtUho+nYbCdXfbZnC3VnLG
E1UWRy0xf3aFXGukpwP+hI+bg3bH5CVCx4RNeFOZ8FavHT4M2gW7/8i8pNEu
tc4yTTMJ4EizDM99hNu2l8Vvb3znZdXmXjwiwYzL+d3vu7wqOxQDaOAD/H93
rJixbUxXPjWKAhaOsg9rCb0FfM3RXpnnW0ju0kVl5VjZlDbMQygIBI5i0Osq
brfY7LdSRTbNsEgJTS5QH92NsfJktuHbjoty0X9EhH7rMFAtex+KpAhZXvRb
woQuHii3K3JR8z8hjHfmja4JxS3aAfayo57Piuu3MKNnm5Bc5Tc9sNLdIlS/
7cVpt3+sYLUbxLQ+osuELCmppJJIH77iJRXbivUeSx/BQ90DKze0/GliYxyP
pLxIXNMfjoN5SRzTgLAxQ/nUuoFIkUMpWjB3xBZJ5zPWKPWppxpPIpSVGeN4
Q2N0+Cqk/mV0WCvFuKyV1e9decmc8EDvjVVcagpUnut/Gu1uzqLGvT+ed4+Y
oxLxk8KewXc3yond2+TRFDY5u3+P/beozSeOaNB8HxL1wEbtViF4SWL/1vb+
aeaDNidRh/Hv6UrnQKhhiriSO5S+mxvJsf8fiWP6C0LFhX6VvJBFbv5eX9Hx
P5fpRaBlsaDyQEpFGHiub/4pk34G0vUq8oVVap1FlNQWaeQcGNa2fUWkOR1i
tr7Cg9L3e3VHEluX6z5PzWKTnECk1JWNXukfXT+3ooG55sgK+ZpIVYQ7w2Fn
WM3r6eWWg0MqGw9/EejwiFsuhjvb/REphyREed9/7CfhWIB2jN7aMaPHNOoV
NFi+5wpmgXM4mSocKwbqbjk/9a96OBprWPTV32h/xU3lJs2+U0Vkg+COKLRV
BlI8I2c7tXX/3wNJ7rDj/XcdbMDy3SrPU7V+9QcuNITW8eVPREctoNR8DMNd
GhRzlYOi0WOORj7bGFoCZwpA7KI83c8rh86NOndGu5aBEDlpwKTpqy4YUpQp
XQcqL2//0jXc8B54p7HBUc/ZwZzJ6z1S9yytgTusFmZkvSLYfkLE7nEKAUQz
8Q7WUFr8+jKWLurdUhKTr+oOVunZp/EQGeTbnL2rR7U3cUglS8s0iv4X/euF
WKMjyngTbsMlYTgcC5J0gKuGNIKNQQaWjotXRDO8C4rl/URuYcxHWpDKTeFU
i5ALbGh+8pgSBO+GRUhvCLk7DXvSz8N9Qh0E3E1OEeePOIcGGSdHbw2uKLyN
PgQtf0dXkpz5+v+CzGUKM7WbvW6tqzoElwQ8u+DWS+yzj1oUFXJnvpUrcG+4
W32zeDh+b5mEoWvfd8Y4RGHc5QnfmXN2QDGwCEMzldnfLS9gAWu8UhYCswh6
95gDfFr0vVSIBLpax7gSpLGKzMUM1+YExnZzMbbVrttx239S9vJ+5D0xYikk
zJ0DH07c+DdN+zAsRHa7k7eSAU723VXra3prPLlUFMNhTwyWwVLBnTbZ69Kn
7vWFPhbzY+cgnWm1NUicuHayFOChJnDRf+CGH747FpPdcybVF1glVZ2OinAp
TftSUyMaIipEWIEb+Q+FIKwsIP8rRavOmG1m6WaDXPWGLnuHvUFfU7B3J81B
XwFLQ5/1zt1ucocRC+QauiP8KmGtLMESfLlAUH6fSllWGsdo1UwUl54BKRJu
pFsg7Z/cajDGubvnk3KEyNccb0ZSa8VUJ258oig2A/QwadhYRI0DVrXLcsO1
rLFJDoXb1b/mBINhLiCGZsUu14UtyLCbOU87iRKFX8/FivtCg0OsbDadVtgi
YysX21YgSWJjByKcbB+DZyy43/x2qTn95SD0hVDUjRGGzTMF34GcCbBjhE9G
PZpzLt4SM3V+0nDAf4XkC8dIgVntwWZpVBhJvlyu5MnCBur7hrCVimW9GpXr
uK5VLhuxSiVyE68TgehVhuJP6KKM6vS3ycBAXHny17BmgZ4ZVBThyV0YY3Gy
qUBVZj7dW2OpducGFKIc9b9ctma86bp0vK9JP0irQAWs96ArB6LbjfyeMR71
TePV7L6AkG6KTAWJ/iIIOZZv+T1xIzFCwk4dXpzWlpCqgb4WxQyr4Rx9fc4A
laWI2nvXnFK3TAW5ty9SpyY1D2tEzU5gJfPK/JCdeZWCH5LTuU+zK4yOwKoD
yrZD/qQqXjIpB/gnrkTJTRM7Do37NCZYoSKoK0Ym05omGeUTdopJdoSow4qH
04hDxYA74dBC9nVTGRP6i6jR+HYo3r43q+HkDyf+h5JWuU7n/IvbujBQqoz+
DAaUuIG6c+Kuxn4kSQoj4+kd/Nuu0KRDMuAEW45W3HyTZ55lrjJFtLnXMlGS
HoAFeF9uNrHI+m6E7uYIME6yRQY5a2T+3L/394PZM0phGE3T5jpDuDSm8Y/p
xbHAm16El3ccRx7UuWTIufvZCgrAPFTpP9yIKvSSo/vOapY6Eomha19pfc5V
AUa9gR2eEWTjXBidqXzxx2lC+CQovOKMuYJgYBqbQQDumtteAcpgEsevMp26
E018He7BtLFEnF4xDsNmt07FoApoFJBl4zSkY0HVmSiB08TbMAtbcwIeAVXH
VLd7/AXAAPrGbwFWQXHrOL85mI2ZgS5u0FGwD3vEkAH9PbCu8P1QzdBi8OyQ
2D31Eod7B5rrgE2HWq8fS8LTFDdZbOr1RYHxG3zea/n7+NzkdNH+GAQdTR7q
DHJFFk7e1VvldgKtT+8775rc3YiGJjwuAJnPbK+7enpqyHGXKK+uHPGw6inx
M5NMS50vo5RuuRq6aERFsmmNwuC7LcFajuminChZ6CyaYPGZGeB/etvbpz2k
0u3zRnUphx62wPe6bu3Rbyh1+R+93NyKAoJjfhuN46HLwOww1HLc9iD97gJB
oQ2AAYescD3SAsKO6cRZQF4FSCtUnV1CEWrbhZv39KYUzLKyjgb8raH+gb1c
48Xs/phRcXGvG4UVi9jVirWXdqWM7TJ4GzZ1ISTNZIYhseYK3DiOnk0FJbqr
YzVeWJzig+uxNuaIskWz6xvYVLOQVEAJ51dCG/ucW1n7+rk6Wkn4r/afrLZl
rQ5TAFxZR0ntmu9jOGi/N5VMI+mf+g7V/goHsJWR6O0ByFh78tvtWOcBhONv
QcD6UktMaGTfCn3qSBDxsKNoP9RSEvCtHU4RknisVFzFQi+kYEyTCg8Wu2ux
IrOq+xNHf7hGWmn9ldbbN/zzgqQ/7TdfYCSwQn3t/La8C3TnTMKQPe+PSCIX
8lxGhNw80aB54IUl2MwQ/zM+ANgkhOAty6HgUmQuOlWPiH35cKiciEDLXkvZ
KzzOJMHrGGeaqNpnUqlQK3Q1J91Xtk5VOmS0hJcRgNiz4OnrVsLxZyWhe+o5
jSI0xXTpXk6PQkx35MoC4vdmYIRYzh0nHZDuA/pHctMnyf1PKntB6ZuNZkJ/
x6+Zxn0arWW9wb4C5i+UmTkRUshr6vodB4rD9YtuDtIVHwFwfjzYWEPqHbQD
ioAhvgGqkEVydFpp3Mfqwi5V3ffO5qzWkODxJ/46hAEtojc9lurQXyVspr4s
5VRYUBLh1/4hl6m3A02L9j2WeAsG2jVZeFrUBZMGEJz4ctjHPEKw34m7ti5D
aKyVWgrPeML/ikpsQnljjrx9L6uYpFevPyNFATFwkuisZrEui4bxZgxF484B
4u2dJ1WYUyjbGHrtvdiNE/qEzug1t5de5Mntfc/q3TqhuvQx0faI4sBn4B5L
RFrUKCxWnBSokT8l8zjHbDJUBHlQ6xe2MMpo6PHfRAN8s2HHmwG8tKZd9Kl9
P/ZVntbYHiLrpSF0tEjXodVcitY/ujf+ZqV5ztW1xppeCvSRiXahazQU0UFe
hMdTHlN79C6Ejr1RNVoQcMwgqNty1yNZ7H/sHCa02lYLnCeBmqHiivcXLjD1
LCxLz0C3HREOWZrt5NBstJ2rCLQG4uMUUmHVp73JpvqO2WXN29gqo5Z/f00l
gkRgAcVIbo8cX5uRTPOCwahIsara3vAeUN9N9KEDn7vHrJ+wasjF5seKZHBI
SdEq57srtqkCa6WdyZHnOGgRprcM+TqdwLm+3AneiQiInKHWOoktpJRHGptO
PS8TAoQRluDVPeAhMHaYIWBn4lfPV2OE1TqIF/foskue63NBC6MiFxnZY6uw
Tapsi5AR/weVAXVEp86VYQC+o0+vz8++fy/8WRilnka2DUzsa9of+Vig02yS
8gCpLzgb5osFXyUA4ZHrj6hIcJSUA6b3L5lrBOFlfHo9DISbaBcCPO8lKl/u
cAtxtPecbdyoDqBnmmN3MYllzfjeqxE1TpX7CduVyw6FlZ78xw9r7DdDDwGL
Pel0mpA0m2K2yVi+9fPUIZcRAd6Z+ZytuppnaYT7H/NQvAoIHDvS6upUQGlg
tfsCCiD5IaSKXfE4yjGB9dV0XgUVA8IZ//WkXgEy6gYlm9MCUog6DMtEaYKA
3UDef4FYLAZfk+E09emDUmvz6MrrJrDCXatZ4asALQlMrNgMzs7hUPk/Tl8C
04Pg/xuO1Q7mY6RYnr0OmkWnzoWsRBQeeFo1ar1bLmzQnySsPtNMrgK9+j3O
yIqLB+sFjlFg+G78v5ycEKV1EoJIInMi1A2Cw7C+491uI34SJgav/mRqEnYh
JKDgUAaFEOLt5jiut7MkrsTwrs2IBJxfrJVEL45filr5A+/2MC00JdxBF+cO
XzgNqYkR/XTzHCUzwOhD0xDTMJXM69+biVclf+WGljljoR7/qNqon3XYCvfF
wMTbXsjuQ1T6RttSbHTJ0KVm3pu8CDu3eWOlQ6PPM5c7FinGKthwjt6ajUFN
v9V8ZiOC0xwD2pceRxdVKr+prqKCFiBAMvyMMWq2ArQ/497WCVeHvco4sAdB
eevAtcqttnMiluECMM8Y5jZGHvtFrViD/rO6qDp1nPh7TYqjOSwmuDpAci6n
FX8/dLMLEiy0Cr1xf4NzTo6XAYR7iytDe4kdinIwlNb8WZxMxJs2H050zJ6p
AIRhRisMAVN1IoA4ihu+YKUNYNgU9Wb8ULX8tviqPOnN1puRoFMS4ukFHtp5
0bqxxiTcEv2LFYoSXfTPYipK5wwUEkxpQrY8OlsfWyCUnlrkWH3mYb4YChFH
iwpOuz+TAqasgexQaNgFhwH/NthejwHqihOX4sn85H08e7NsRoFpnnD/JXlu
VGKDcUOKNcLlCz1kCAjMFolRN+CdplKDtSkRKsFumIm3CIEfJJEQ98/86Y2F
O/tLnZSFX6HwvLKKFbQfnyHCvU3MVU3dX13bmIi4aG0oDu3crNfQhy8NnILP
AxedFGhu45zWJt8wAUnOcVDX9pqEAnG9Yv27O/FNz/UPxtH8TDkQ/4+51Js6
6ODc68m9Oo4oCjoDtT7bhRMzPud9tv92roYhv8MW2C+feDyf9X5eAXCL5tW4
yGzBvGw2gWiYlKNJMuyUeLfBvPqHhorjUmj38EYtqsLapTijKi0LYAs1kdvP
cbmImDrxMn4htnkYQ6zq9uOMZFNJ4CL1B0ebmHvklI7Tbz0wno6Y1l4QCXx6
i8MZl5J99LenXkLE0s1gt0Pltl0WmprdeW/J2H+fBVviURFtJVG8ck2xwxGa
j/C7IQKbo1bn6c0m2f+uD45gCkPJRwk9LZ23/h9JPnBIHz/AZLrTcfzCEfUk
E6aWCp4CpktEK1J3ABno1gl9s3EONru/K2AEBx8CrldPTZcp1sxf1BCAfSLB
Rn6SSlXUXeoWB6Zn8OUqpZKUGqRy5Gi5ln53tKWOeJD3aeWaa98NaLT3PkWD
5Ny3Hjx1ZhU6jYaBZbaW39eEpdgNUPt6sQWu0x2+SVZufRwed31cwqUwL+Pq
KwFXLdP8I2DOhEr75tlc9tN8dUU+UjFP2JM2B7NCi9VBB7RraPedixDltG7e
7hxJDwr9mY+OtUyMVcSJSwR0L3DaIJ1TEfq0dtCUnuwE7IsdGzBR4kvdETVg
hTaUVuOvKsdQb+Wa1yWx0oiwFhmbZUSx74aAd3F9sBQbXEor5961/Z7OgIjP
zuoO61TWuytfOrVhoQNYsw6NkD+zycBJQOWYcp4DSMoEQDrPsT8z94MIuh8i
l4QxhBNpZXKr9/ObfVid8okuEVxpEBKDfVwlrhS5RYvnQ/fI/N9uJXaC7aQu
nOeFiqDeerVdyEEoSAZhFgFSxYCLxGMKrlv0+Dd2Zs5xI4sFAOCjMV4C1EF2
dZwrVXqABVmn/ZdHS70mCHGnCrFbl8ZA5AbpaeRJCRyk/kFi8o0a/6ilVlOx
/Hr69283yTrrXN/vRbbCksTb58lAvF7GUXFf2DhHsQhwqupY2UOC0csA8e03
PAOHFGaFAqph8dGC9/gIKJ7X76LOEQC0Sf+/iGYNpejIuaQVNDGRPpS+F5v2
BQ1968cSD31nq+YxaD2WId89StFQSGuzQXOFaSiKP+q9oRtHAyyl2wnX1g5A
ImlPjqGBcdyeqdK2+mWHxijb4D8Y3RXuwGMA8HVy1XNCDiZCj0xEQmgo2VSc
kOrER+1FhPozy5jJCWcSoZigPm8sHtoDxUj4b75AJTGExurgA0J4d2m5I94f
pAenOq0mvlPiDEbCbc3D1lku9U2He8lzMt5GjLll4kTAPA+DnvqEV2f/G5Uu
i0xWlCnwOn2mnmoEbeqTadSquYBLDMdCCHIK/aHxxXU8cFkSOKZE3bn+FZ/3
OvUe3fjB3Nk95Al5E3yUOTLanuR3oFgQMc3qGN4ZCah5f6GCxnDHN4fL+YeB
eZuKwYC677vcUmQFQTLe5ZqACN6Bt8sWpJfekMwq1GrXTd0V2UM9TDNlU81V
9wwx+HnSZJ3mXVqoGwjUn20s38E+EjfOboE0AIPqZpTycl3FAiChJI6mR7+v
26b3CNXTB31yjBHOeT7ASJMOCqb1itV9ACdUX0WEuOfIEqVzfWYsPbzidt7c
UBP4cMbZ1DoE7swRDRsq4W5pnOAcbHMbXJzXWcB+wzckweKRTx4Q4m+rxiMz
7MzpyhR+8qZziSpQ3DovAGxFMrPC3XjHooNNDuARINo9jlmnOx2lpRtCYTLb
iSfci2nWEz8JX9W8Kr1EkcaROVlPb/10JsoEcqGsDygg0qUO1ELJxlcM61Sq
EVw3cL4nEqnjNADwN3kRM3ZBupmLBchr47dPmqW2+B4JgfMcEm1F1emO+3Y8
7ky1HXibefxyf3lic6vkvNQ8DJxmP02194QlcGXmVx7I1f2AKWXbjxB2cnEh
CGmKT14pGmDMgpFQ0oroxAFk1esg2P4zc09UTBAPtxj+y7AYfpRXe6iecyv8
rNzTVZlSiuWfpXacXDTz0i9AsvvWaVo456WisBW1/375mFmNtKdydpE8lEee
584gP+4bI/wct36EW4IM9f9zqpyWgCBbCC+hCijAyB2+e6f3rvPJvZlISZIt
2JgiTZbLkMwTz8n3auL+RQ1AmtuqWan685ghmTJ+P/FQuqfs7RbZW39u6cc8
w6YSnYxcbc3DmpMpSC/88hX5YU5/5/FlT5qC25IuA/crRD+hKnWrGhJhv7/1
MBOO/gnzKJy5pIo9AJ9VTrhCWc+d1MyiLswF+57iHZBKE7hoMuiDklIWt3SB
E8YckY46rq7bD06Tvp1BIZktO62/ryoTBx/hX6CsRDlY0gJrn5AWMBM9LqqR
4GlYb4OVSOnugrYFYVCO68U2SujzLL04LWHP2QSbS9tKzZKJx6kryXkAex7N
GWBFHYG316XjtqEJOvunEE2ODCydSidLHgLNL35Imf24AN5xh50y77r6Bfkv
j88TITZAyVPjl+rw2Xb4fq+PBhDpMsLSfByezbrgV8uVyHyqYyfK9lOTGc6c
6dQINcSAlaHjaZmhyTk/nbLIzmMnfptDNyyrsvKl+kfMHBEnO0vgLe36GC8S
0lBI6pkbsvgLPc3OMwjhaaZk9iL0Vz9NFoZUMb7C/1UVlvGjeFOkqOMSw2qn
bNxx8n+b1svTzKp6y1SN5jeP+8lW3+EPRS4bh/jYsYwGoOWIsDYejc26PryM
XuTURo61rP04Byo3EU8TwOoNrMbsbVRJlaUdbW9gBcv1EGhONY8iCNU3N0Gj
mvyV0G3HIeqG3J3H+xAl6OqgEW9PYqfmzfA+qtlXoT7y4hDrcoJU0ySw6QgE
4xEaaNlF3udexAAlNhMLJgJPvWBfpVJqezYtjNggMvoPdRNq7zkufdcC4Se8
HiC/aIV6d7pFor+iJU55ca4PKpz5eJastyarHDlVPtTqfnAMfD3lP8Bogclh
WN/cHWgkqH9DnCryPs/QEpWsiud0k/jUxGNYuLYFMzQCmzjeVgv+jnS+YbHn
CZCoE02coi8yVvfweO03slaD9myMem1qtBdzadrIgMmkly3qDnJabXYvH0lO
Z8ey52FFiUiBq0ezivo7u6GL7TLP2fp4mpHpG+lPBrr//LR3zf6zEKU0jyzB
7QHxHZT9EkDCrKInktbI/LXH1vaTpB7upOjNbJ0DfMnTOZ8c0S2Bpum5dkxj
BkAohIomhRTrNNcTLUjhSZEZFRFI7le6brhpWWotFqmVzDD7/BYaiZBrEcAd
rZ86pX+09ZnlFTDJURid2uPdFdHHMSVdcXLgHf5dgPzm2/AllF1xCTH++7uT
X+j+ljs91ftyXa7EwqANMoNNPpQWVH1ZjQyDCuLybH+yusIue8/jRFtIqu7o
ZdavDj3vz+RCiapDln/u5j6h6vumg72QCRRe5PLBvV0XTABM/CCyCURBCcDY
BwpjeiJGLqOPeSk4LHU/aMkh1yD31aoAkguH7MfhtdVCiPoAaFmf97dj6/d6
qR4IGpbvMPrgBW6wZ95Em0/QqZA7LrTDw8jzYEZyAWCnsktFY8ceFhpCgO0X
+VEpKZEw54VwCu3/Hs2xDO8XG8+5Ipbj3y1FXHXIsRBm/zs+XL53HMvviyln
09wh947mmmIk/7V4NoPhupNZt0Pc9TUZVcnd+EDdyOsycTyM6ahIha/b0EQR
KVysnvpN25QoH6qhExQ737hFd/ltMLXRVOk5/IRe8iAJ17sNOgpVQu8ik0dz
zVFr2VtgejDHUUP7piEQdzqhzfbU/7N8FzTC18qQzj4P7dviMPB9oN75Xh7A
wnjrNdvUZmcG0uDpgXasY7jkXEsKuKdtcY4LHAlYdMdfdmZNryiQTzopy4Cu
q+vqmgqWRyMwZmHuttricvEQq1wtUHHSFO9djoSYS/O+prL9LPwrlZJEj+jF
bPBCWkVxkQj5IMwpz2ugxieq2ecVe8RsFKyFKAJzkT/kRiDpvR5uIkvTghWX
oc3R5vHTseMHaoEvBg/o0tuPeRAG4jK7fT/23Rpgvgj89E7zZE/2VLi9XzK5
2npNqjqeLtlGP1lo9zpIrXcWlB4IjVBdxgIvfAj7H30Ti8XA8UiFSkVu964L
RcFqbWTd70iI7LFsgR+9Mrh5v3ZIK1QGYIpVHelF1F3fifSWKaUg0sbFmzXu
CKI/h6oxzJEfX73sGahnf+l2Np+ER9x4rUUh+c/s5lHukBLd5KgzLJR1XhH0
n0O4hRQB5mXGGETsDL3cqyB6yPg96wodGYbjy5381DDmlq6sM2QC4zYrXjyQ
KK1qZodYhdT2ECabAEc4wmZW7WmYIu4kwnLkdK0JNPFWv4E2Fp16fAZWHFSI
GwZqevoCyv5jTxQLkd/JrQ5195TZP+x25id1Tn+SoJVy/t4JXj8MOxw8z/L1
puB5aYh8EVr4DP97ze0uMhUHQVink+xQshUqMWF411j2UMlOu1spoThIFmh8
jTjHpC883nJETWPEsN3VfVLiNC4IyHNa2a7wnbBP3jPoRtwmZXKjax07lB1/
DWzfBua16MQYWS+4ct+dh1VGm0C1cPXy+EqsnCkrNRs8mSRQhF8p/YYt98Ky
BkZSrOHz1SplglByx+CmAThl3bxgnGslWVNdjv/YdxmiOd5Ywxq2EhdJO/qF
R8pcHjCvc8mu5UxT93iCwKeHQnT9DqwXeNmHH1Hy/AKRcSDkwQ5q282Iy+Xo
gCdgjitNldUEi7OS+o6tTN2V1WDpIkLzZWPwJC7vfJoaAdQeYvT8HqEFcfL2
qffHmZ3bFNSVBVq50Sy0zoGHIAo42wxby/Tpe3bM9fkC5F+O0H/dPwwKR0fh
ZICI6mpGid2i6TlhZi4RFMGc4aAu1Z7ClFX6laXDisFEn1RE7mYBeb2VFLzK
myTIn8pwxTEmjLPWrIS9w/CpHyr5KGypPGTjCTxbOc0+4MbeMCuW3v1xuqBf
5f1xS2DGNK2VKWgIDgnkzO59WdiFKDWO6/OiniXaLBD3bqdlaSF51FbGE9xF
F3JQD9YJppFkDJJmN+23oM1fUV/oAqsd8ztn22V4YiZA0TJ2iBwIv1NU2M2D
0JlXOt4iCrD5q+YdTTgHS8ncqNPEUhJANFds7+3A35pYzvikgOGTmPamWu8Y
O9+fKDIaZ7Ay4Pg5R1A2i7m5Q1/hNW6tP4LSV3FS53JBz3jMrG5a4Nk8ORXO
1LMdAH1ujqGVoDiftBwvWj8/nycvSNSGAQbT8PHiLsM3T2laU9fhyUz6asgg
EE600SbgmeUprBHXThelElhbrgM6Q2SD6WoKqBL8euoaI7PuzdkBkyNkgtGx
EDA4tMLuo+Ku6rzBHgcnT67MwnU35a9wz+E69Tnv+uZQooiS8o+eYC7vpKkc
dYQ+gUhDZYpjFr9leYfqqRVTj6r5xM1P1egFXU/AqpENVeF7iJm985VeBOYu
0rmufyyrMQ65jd8HowukFFmBXWmbIMqwB0JL4rOTUlHYgkqh/pFjaG2oM1Ev
fTQMu0rM674/ijHWO4EkqjCO+xeHkejL1mRQn18rSZtrxUIDKoi07ujaNFO1
2D6joE7vdTVSCSc1BML2chWzwoLuX+UqVa8aTiaGBA0rWc1CucaG1OxLhQDS
TJD8RfYmn7quYkfWbm/m263kFVVvBoEarn59Hbstyb8qjdhtY0Beo69q3akb
AKugJMrp1NMr0cK9cMXizu5oG492wGDgF4y6AnYTkM9ZOkwsR05y4kM5Vlyn
e6kX+1W07DsBs2x8EXNLS8nyux0f98PIA0XmCkntp9h/B3dt8jAeD8enMS1F
VUKNtBBYMYQNtfU1/frvVlcnVZKDxqo6pU12egnMNvuDbwZM08J+zIMAWfaQ
+MKf7X4NHUk0Xt6L4fHGWtep+J/pV6YE6GjxbLg6+44ac+H9OojTeMqrahh5
5+rLMpATMtiGGakK7R9e3wL+hBGDEPuySZ1AOy1FWca5YhoPwOTsDUIqAP3A
LsYjMdc/4sJCiOW04/+i0k8IgAX2wUwu8RoNvIasg4Dnk98DMjG3wMR41tCE
RNCmGZkHdPN9DZAymIqnpbuxzq6ealfiISAzPBIBGQ3TNk5G2NrvbAtPkPGy
3iVYbEKo3nS8+Ui2pk/k3VCqzBF2J7+ZAI44TWdru73sK7cfHWplY2MyILEK
LfwX3BqYq4irkUX4EUtZyfFf5G+ug1oF7WjLoGXVFlx3YcZUwmEgV/GXISpB
x6QNuHVucK6p6LH167JlxXf1d13qELxubiTintHaiCswStuNbKvsZQE46OO3
EbHa//rTvBuQ3m6Rfr6eK7tQGnJ/yowYYSQ6arg54eCLnyIF1KWJ+EOQ9HrH
FGpHmb2sWAh41ZoQQZs38ZkA2M/3ougV7URDS+1mdcSV3hXl48MQ8IiuexSg
MbC1gZ+UitoWzkGkitQLWyxWSGv1yY1ve7SEWtMarORaXrI9yALMCVwTzPBz
LNar4xg6iHKwd+nneMUq+7VxvSrJX3zfUdz4qML9Ebfrwy5+MSL1DdPi7DAz
w/e2RzCVTN4WgiGOqLm9kVXK1chDKytlAnwxJZY6MQB5qARsDqb89klAehCz
4CiCBGulhroGJkBU+wsblSkpcrDPVGh44QLsz9cP06sjNtp0bukf0LalqoG6
6Kkt7+Y90QQofo4YiPZOpQ1Qf5NoyMtXfiLPl4UOdVnCUWaEyfIJAOc4oj4e
cPqE8fjWv6XV9uygXL5C0WE05/98XTiHocEUSpiGrR4oZoKOUn0cahpYUieI
F99feqKpGJQr2TGNOaENrWC2snLGNLxmPOcxK99BXJrilj1cjqR4EyPx10MO
/e6GPGEL0BdMpH5oepCzfibP1AP0taCUTusrEAbXfd9MNSTuP3ENWlrXHJIJ
bY99UgX2XkqfsV48C4TEILA3AtkFi75LwKEoDgpSNf7LqwWaNmy0GHCiN4A8
IV1WPQnv9fFoSluYquN0+Mr9546pdhEE7YhUWlQu6FVtHXfgaOMrIJmYlWUj
Ic5l2JFFvvCode9XWHiPVvEEpKEe25iHZtZGYjXqa9NdfBTcJC1B+hXGl4+n
loVOQ5g0ry/bTkKumFZY/FBpV/KZ68XCphytTMD0aXBF955HdMJSKrHq4IKW
YISNWO2vBzZwL0ceQ3lVL/FzvIqWUyw8ZOD9VaTzSsxxE6GTZEh0l9Ckfl1c
iQka8d7fUgkfKS2Fe2GStc9ZA84eQ1VUvvT939nJ9aO8B2f+fh7SbxsRVNgq
LA2AAXuMsDh7OKv6CrubuwjZ2HLYlkt8mFvyk7dRu8EEjlXLJ7/di2XffEXO
K2+X4YVs27YmzLAj3oSRIviewy5mmsvGkh8P6tNdVQxOVZnQT8MB3P6jJk5I
meGVUp22rS6+Eie4BpEyhyJop4J3o7gzSyGbR7ABaTDh2TdnF1NoQwpBLHFH
+W0fQoWJiPSvl9qJxgJk3HBOQ09mT35GEMYADI6PhfZwS391hZJEf7HSDBHU
lhZ7mUtG7UI9ABKg7HCt7IMyVsa/NyjoJ+9JWMLgvMiCI4636iSYM3GRbQds
NwfKe2OxT9e7QsaFMr6IfJa0m6eT58RGfPc1ZeV70SlbxlAK5UBvPMGUXkOT
CmmMrWXhHb11n1G9b8Nr+QJSnmz5PHZENNxmTE4QMY4A+6g+VwvXOj/MqEI8
DoXGKZiP9ZJ+hbVwxPvfbVzRGNyTpR+C+GA9wUBAknqMvCm375Ui3D6++ctn
2lmdJAxWl5YcnG+BrLHuZDsYK3e/8ZBXNUr0I3iuAyMz7utiJtk30JHFLIJk
zQuRHgqMtnNd/RUc6d3x3fHgD05jBwEqn0WB9yqIRPdFSV/jWFuviGzxQzgm
TXMeI6chYQziotGX02Wmpn2OcNcSlMIGALIBPa72VywAnW0Ums/mbgCB8+J5
Y/+1NbRCbk7AMI4yF67JrrVUjW9ndSEhElJ06z8cJPty/i72gl7yGRfxi21T
ik7yWDGMUMTPeFz/eKqjDNsWQOL8N7ZA49LUj9PH3+C9zWaDnFCsZ4mJqCzc
5KLZN8gHGTXHnKsrRdAVE0ezCSLqWnZRzNEoTUkoWZDYr5U0U6jxw931DU/f
UyjDZoE5gUbSc652XC8d9jiM0VG0S9DSd0qaQNNltgr/zJmflRqu7YvUyxTZ
4qnwgo3qElSJLYmwnXeSR03zziK+SGeOcdg97sI6zOj64Gn7FoESAxbQVrv2
EHEwdarLLZ9HjzjRREoPOMjaJU1CiW9ennSHdVsr2eaXt5/cw+0VfNWInwY4
jrNYRDrmxPTU8EZDaiL97G8LF99M1iDOLYBghejdAcLe7zdk5sY6EPkXgpVs
r3I1geUHPOOoHmHw+dX/yLWn/aC5yreIwrtx73wx/POyp0nSf6y1/RdIax3S
w+267jsjOvWaOiryeWGVoRFhvfHFZdIc7qOjNB2d6IdJVRBE4oCwp8X5Avro
YF3P9DQYj2DL9ViAXSkdfrerG+UOUUVyAr1/tj0g+M2pyQGbBt0u6h0fkyUF
Sj2SJB/FXlXKNj8NykOfEXjWIs0sA11k2P/BpdGWualIWodCw/hTCZEOIb2M
pSwb0ZqG0ARoMsJJOFbgEjkcNictUsfG6mAI34ISYYXm4AmtqUHpAJvvrzcU
3i/6Tnye/zZTATYZa6QpyJ3ibrND86jPzTXKEKmwQwS3xua9xuseQdtH2foT
Z/I7rQElF+iP+UJz86Ma65kMZ4HHJFKhKei3DF1uhEyv4n1QI+jkyHRh6HDY
AGP/XFaxxz4eKchvEVAGovlmuqipJv2kJHfJeNB+tuug7OtFT+y0Sz3fW/9Q
GL/bnWQfjBtj7OKfvZKioU6+21Scc3eZct6gtpJ1kEQbWMUz4/qR/nhTikKF
1rvigGGv9SiRtYG3OncLBkagocVu9tQveRnCwJA92wlAkJ3tSUDq9UZ5z4JX
wceC77wNpaSomBE9EMYnErVT5HniACZN7arQMH82eZxmdhxNI7Yg866p0VGs
Qr4H2wFfqB/Q5C5K1y0yalTopE2dZEU9NkobBZLzbOZ0q1TfDPybQMaCsn3C
OMCU3Re+9TvddD7IZ8pWRBsJWy+sy7a2CCpZIWP+UqyUHXH3zODSMSVBHHEM
zqWxAKYwCU9Zrt7ZSq5BX/bJyMwq9nrU0NKVN79curYnR7Vg7nuhs9Ydhee/
KIDMMqSVE/hZIMd7duR1Gf4H5uazhOX5SsibgHPu1F21labcrahnhuNuUdE2
1RAi8qecdomx0rg9g65n5mPnoRpHD+lgzil5ebRRKjmZZBTVA4hSqpw/zIAM
A2Za+ko8JG6RkxuZ/q4JZ1IH052utH+sUJtUviL6fFwk2OTAs3ZOr0//Mbl2
ZelvmU2RrT5YCmGf+jbK2MtJwQ6mvF9ofBY1Or3r7lzfbs/v1VEkFez4aVpv
hxpFOEr1rQKN5PvoSgLZv24BCfIW0RJkYA8uZJFc3IgzrsKviQujajF3m1Py
t4fmbCDT7koKibgB0kuazchuQJBJ4sdhvK/S+fu9GhKGHgDZIotnn7UhX27v
kor5CR13Geb7QcjUDg6g8LKCAGpuGp6sylBYBhpPBYtKbRzyEWHgUtb5Kz29
lj0fz5qpUwLlEkyozQnOu4CV2QkVEsd2Oos/R2UoeJsl3ocl6X4ZyAGxRd9S
bo3tKi9SVylgHMnzAHJW4rGyT8VGwzWsWg4zdDhUWeu+H8qbcGhYatFdT9An
4WIo5mIN30cY/9m5kerClwi0ExlnZxvkQjFcw/aeTbs8wpws+TOQbvxfk0L0
wlQ7DIak5RBP8Aza4v0np8J9MqUOH/bNZ8UgriBZWhxP1hPvc3wvX8Iov4nU
6KyANJ1+0WgIVwZWqZHMy9shpDh9a3fv7LvcZ36iYVdQG3lxlj3h0uXVmH4r
bxJGE2xTLaJP/WEHwH13nNTvxmn466nokqycaaUSUtJfEab0sZj87hVhb7SR
Zo1V8C0SzopSjFnmQ+X7lD2eHvWVL7VNhjWhLOc+Dc3qWvgnqq3AR+WgJlNU
HABSlp37UaKabvT0E+9iVfiy6UrlUxBPORZMSInwCz6CZhvfW/cBq59n5MRb
Recbv6rK1LggGAVodXNRgSiGFFH05Ns5nwXxi7d6asAbbMWk1xN9qBAuNpEB
r9juZD8kyKEwhoIoEDFnsY89c8rMI0789QgD7QQKEO17e0GKZ1wSiB67CS7R
DzUGgl/fRsm09zRObNDbffD45WSBPXACIS+S1FHJp7IG4XLmLrwVEfUP6zGM
LehU4oXTBSJ/q73iJaBl1aCgfylQ+aDIBfZpTEBF63kbSiFACK66U9EOF2le
eZ1a/nOvAKY/frZn3kUSzBmiIXh1K9mqGgZCVnUwR2dxBwFlukbWSbsCpJCz
Y4jG3eDPhc2LRJHZz1OcPrL0dJYVdub3rvkClQlO3Uc8ytvNqSJMfC/mD2sT
cdQcsLPgKeth7MW/VWSYGh0YgiwVbLH7g/x5+NFNCsgX+KYi/L8WXojoF1fY
Mn1qx8FPYaoDRc9dAiELJxI68QA6no4bWYqyuX8lJm72Jb1nF4vsZUXkKhf2
Cns6Gvh4/jkvVXbRFhDD7qJrOSQkFJSokiFxpnLSzk3Mbx0HgPAWED2tp4A2
tz75R6HzVm544EFGue1b4xMpJTymfEBmScsC63yVA1UjPAum64x/PyiltWBQ
PewFVU4fuc5q4K0MY82jeA2BSaxDyOwKvTpXVdg8Z8MuKZ9aFsXnagmgsE/X
l16bgmECjoz7yxIkV5UxkltENmTuNTOtIGmqq6cdsNsGbdzvMZZoi8l965oN
I8W9WMntiFI6RahfMywtHOkjUUuIf2Sa81BkY2+B0hE2rVtf14oDQWZ1++mk
XM3jT7G/hsbxMILCqQen+l3PiEwUu0mIdgIXfsesAFa+7MS1vIxO1TAG5cR6
zU0yRyQ9UnYiL9dtO5jWAxP66Ohgf3xVa9cD2tG1Q256cs7rNWR4tdEuWtMZ
dSGUyVuA8WLIXZS68x2TUnZ/YZmUgO8VTDOCyeJ7HUlk7AOfFAJfdjNAWsHN
Yln8vGU0nlGOCRGqAxqwu5qq7leVV2Jn5MbUsDlJITrLcoMy22A9y8RV8Ksl
2PFdhsXQ9KStd2bLXCPk3FTyMnMxoYaMTjPMIpSGoqQVmHmkPMBTe4p3RZ19
AVs1b6mP0YcjSJxpW0U9wxlOztRqOOUME14tZvoVbuRm/4hybPyChSNQTPmK
Sq35g6CtifftzWhydVLnIYjrFET2DVZ7Y+6u1uW22/Eq2Qnf9SwFxvconiSJ
Z9o64nOHWCLhgJ1K38GHOeqQPHFSwbOiq7C2oApuF5W0FLSDzD6AzzoAmGId
H/+E2HZOLtvcdHMCoQRq/XXrwe47sW7nSzqMsYCYLCkUejY7CqiFWXSkFHWc
j3MOZtLp9/njKUusTQtIyGexRW3Sw9jelvCH14I4FKkwoVUCdFyYSWD6+izx
8g+VfWNXJEzVWymlgiR2nW5TWLGYGH5/t+DWTDEmcolDGz+7HD0/pCESi6Vw
rugG0gmSda+9F60kULGTpcfYiaABAa2VETUofyuQ3DhhjTSG7JKuhE0GIQLt
ZFFKXsVWPxyZTOb7EhD7YgOh3nXHxdewBnhY/dBSbFjIcbf61lWKo1a2bzAE
75xyyQp5tDlzrEzo3nsKcdEh3pTL3GM38PW0HTeI4MZRcG9a5WwMgMDGQjCl
k7sbFlA4fGpdBFVejlZrnfG9YoLwL7hIV2lRDKaUf2PnW1IfBi5y/HEfE0hr
//9YVKq/je2by+UIuTrhkzfUyiJ5g/eXJ7k0dWurI9BlL8V3GYBHrnPXL2jc
2qktSqDzjgb1MByUJpicQK/daFH8xYlp/4UItKRiCUW435LEIPxNeSPhz8nX
0OA3hlgu/mUSH7/DZK/FCAppgFUHXyaMsZmYt+zUZbrYKc0jDAJf9mUV7HyU
UP8uQqpLpMD3FT3t0rgTqm/iXo23lejOSJsTjH1OKFFGi38rbdj53pPBpoiR
oLqEWvX3Sux0Vb7gTnUC19TAgCpyjhf8OZdjfYehuSJDrMfL4mGO70mta8it
Y+WvqWuHGQPgRTgSNETX4Bw7i/qYEBHd3gjT86d5x+bmT1T82um0Ifl9UnBG
KMMDPZ9xex4LhxHX1tUNhkNew6hZkYRKcdZ3FhbnYaK6yU6rgMzWm54qQtm2
kYjKpQFIZ21vH/U+3Q2/d6eZcsV/GzMg0eaOsCoko0fUE0Ip6tWvY20XvZ3t
zVuxL2rzT+B02krPHWJO7k1nr9DZw+QB1WTOXkLEKxcwJZOPX0xxOPnf3ssu
AJzsto0RCyxE5Q0QZ8A7pqQqkO1vSHsSlsDeDmedR7wEvZYeh6ndiLj0FedV
cEjSQeorXhhlpmP8ns2Dlkr68eyYEsOahwr636vxkGZbvfdjLM6IRj+Edopg
+x6o2mKbjqVuKCEIPyh2/TuxWG9lAkTtLCu8wRYlFql0gfzh2NC/7EKYm9gY
B2XdOgFMBGBTct/EDR0BIIXBqVHEsrDRVhWEGGlNgwUSFckw05KO0u72iacB
v9mLiGvvkeoJG5FgLep2RwIvPNQ7exAUHwWafZUnSV1QQ+2E0FRD0S8I2Wao
Sze+Gvb23lol+txhyBac1ngq+rCntaQCV2DXQPdOTkyot/M8xfElpgUCo2xb
n0Vlq9qokgHgsrq/joOnMFmA29EcnzwCT1PqKTxD0lVIUnrXe4ekiEqf6iJU
FK2BusE66bBkOsUQEJdT/aX1M8D0PB6S5E3jJtiXnaVcLzHjsWXYC51MVCLe
Zwkw3CN0rRzKrrdozbagV6yrsHSCxik6sjPv71H7pJ24Hlj91Yll4zSgpLg9
RSyr4B5NysFEOw6q9zhH0woOyWuNlv/xkmdNzJQb65LQUIzbtswPHq5zTEXz
JAoe449zM8qZvMaEQD3qvdgrVcVk4kOE0THkNjOT+zjrGPTHPsj5BVPMabkk
4QMyv9hqc/aAmKlH3yRXuBsA8ZdooNGgdihxYfVtGbDhq4wipGh8kjv6ahUI
rAeeF0d+Ve+zpSbELpGsAP8N6nrqSDxpLclqGmSx5BNEsBIKlwVA1xesfPda
KEJe3d7vmO9ZfFojhUbPs0W5Yehq481BcULo+brllU+lAPFXmLtW+Tog8zdM
9Uov2kaX3bN20ezTDP3rGr5o3GHRt/jzF31mq9iEVpdJyv0uI9hX9+wb7v4C
nbS8R8BuT4rfCstZDx/s5x96onwX0yNea98erPXaSlhobctcceB0j5LnnGig
bQl2MBc8wd0vF7HCo7JLYdTP6g/j9Bu7EL1JdlaFmHQoyjoleofSqTkueaPa
ABRoEdyeIa3MuxgEYnFZBIflod2hzolKZTCSWqtcgyGHwTUbeMl5+8agQJaa
Gujo/pbWYVMSfCG5IXMOcocCCUOYLW3Wq5j1YcadmLzJPyh9+O8SVuiVnE1F
W4KxdpdqKTsUtPWn/VfD/1nkbocThvHElTpKhhuqTZzd/QAQWh00rb4PzZK3
MQuBjLCKd295gSY9s5Z7qVA2RTd7nhONc+rQPg97zcr5iNYYEkys3jmQ0oGP
5/OH6nmlkkjh/7+XjXnoCCgIPaFivLiz9e9CPOjn3SH5r+vD1IEb4vRwbOCQ
FqBGCz3YjXANWPj/cE1w0q4+CuezlSAppN8gWGYd6GdMlLOwc5WBL+x0VDJg
v/gcVZpwsIHtfV9Lk0cyK8/QLB6abMkU1XgNZ+4QeMD6be8/EgX47r1MRyYT
12tDaAyhHuTI2derwdpKwDza6kam9iajjiXodE/WvSb9tKLyRLgAk23WXoON
hXuOdwFIU6YVa5kQxu6CbaFdCZ942GipfJlk9igKTgasW4fFt2P2VJ9UC/Sd
hcJm7fN9y7xGRbBMpDGe70DI+bLioCeQV/yBAydQAAhUhh1Rv9Rkfj8nh0Ny
m1nSp3I4BE1MuPY24jzEZUroGuDuudEK6i9si4GYnqL1Qg9hts3aadzKygn1
Y76GqV6XNWFf5ORTLQDWK0gLRI8qJcqSKCqws+MGIGzrB3L9TM2mRK+rhMEq
/9AZKaRUBBivr1RUWbDdW6vHskzJz+SEIVTneBbJXv4iimPe2Eac0A2Zh2R5
utzBPZlBX400zvX5itl5D6vQqEAFmy/mQQyUfV1R53m7rq3QiPHUmA7vTTkn
oefYseppf3kJutpExLw6wahiK8DQeKBmLEE7AvePe68PXCfrEFjT6jXTtBOn
BjPgsIh9bhe7ZFNupW7AvPIS8B/s2Yrz5kP7ptk1pJ7HstX7yaDZCVDksOxa
Z752dkPWZ/LTD38DBYbxTxZ5B+cdF58RfGa6CUCMPrf8xgMt+8AerJUNvC2B
kQvH785cGI+KPCgTSW4l7VE/4Q52F4KX5eUFYSHlIRK9xef9gAbCyqeoXtEY
9IEwaI+Ufjf7NqzEpUl+Riu99qzyd5I9v5L/i/u/XzVssiEIwnMc4UeyzFOl
O4IXYGaQePBcp8IZuLPblGkmHBbYtY46Hiixxq08ff9T5H7HXVtnAB3XEaD/
DwIUc0Ixm95Xs1N86Gq/4gC3ZElLWSXBC9cGKifua6MCukQ9uSxUNUt0bmZW
rt3VZVQHz/REeXKL/hG3RPx76l45jwJDmEyrD3iKTI8NT7kET7GmZcJDJith
+7c40Iuhch9er5zf+u0G9i3+CJNFBd3GixH9PhF9tnbN6Euxf7UmaO8mmGjQ
VGf+DCS/LMDoJq8OphK8WHgE4ibfNMmwkjeUmXuS/7jy9f0gqdqa5LwHMsUl
Eo2iHvj55X0nUqampmJzROYgCtMCLlDmxfHvi5Tq8TfSsnafiISKh85MXueu
hgGjrBZSDl2+ehmeDC2BaFo97PXlj7jHbVLT1PsImJtcbt4WiG0VqmbWtcns
x8X5rr1IXiOE6fkGsdoqj+UE37t64bE1OF6Y0vCGRD1f399wW7EgAuaBW7Qv
4YDWu79dekCw7JDekCeFe33/v8i5P+JTy9syNHwkIaZQ6K49w4grfaRmnfNz
SPi+95luEFlW0r9C0ZMsfUl6958utS1ERTIGSNVCans7a/eXEreiIi9Wuv1N
2qqcKJDIk417wPJEFYQZgpOYEIvfmq4NfLPsHvKNmdnmyJfOOtEAz6taoWUe
J0bBFleAXOKgfR0vEbWYvKlMcnt9CvGJas2LHrQcEQU5GxWlYfn54hj3fCFX
eMV8tEhe06wJhI+Ze2s/ETP73s6dEWOOjpnEEuG9OmgtHi2BD3O2g+RkE1g6
C0hhjn/2BoTIiozYUbtpb78rBurk1kh7iYq3h0E6lGfm66hN1QaWXXGuVO2h
GNp03+dPzb2i28eAOAwf7VbZPvX/NRsgjtDzhuSxYEErcAVus5AMAhv/Zgl9
xwYKv0FlNpWrw2bkCIEf3RrOWmb0mkrJSrjhaBnsb53cWnCJRGaMvcqekALm
gGpQdPPiIOjPEoc0I7VfgQ0aKkDpR9E7wIcD+UQKbIgvRxiqadxbd/OjMUAl
RQEk93hHfqh/suTxo/h2fVIyIVXs5udRFDuEa5Ljy4rkufmZDTtRrUEHRmcq
/DnIT7uGQJlPGIvctdC/ClgiEv8pK4kRyA0/NWM/QrQoEO71niv/pbiBvuK4
YP82bSd3+G0Hbnkf+EoDAdNb2zDEOC1ybfTblkZBE8yKRKM1DMxrklh1MHsj
HYYrZ/Ctzc7GCEAseXoZSH/3pyp2jiblMDwt1Ok3lLsc/td+i3VjbXWYORvU
u7Te3tqaA5kDrwaY4HKxrkAOe+aPytBoBVlkt6Cbh+1qdgQM0yUG+zC53k9U
aKnKe2PHqW6vWLp8dUUlDAD+dVpPSK+ttKIBo36rRSwbKrVTVE9xlklwttOn
T2d22OouDNlNq2PhHbFGmyI3Qfm9Qb0+DaP3nQVynIg2JXvmOzUkIj+SuMp+
GRcUbta53UFiUzAitwK3Lqk96GXDjyDN8Lwnr8iHAtnpYK82KJYoafxML3wN
JAWJtss/A3SAH0AFKKkIWStwWUseIoT1CLxvLB2CfSlwSSjL1UP7cf2mvJ/Y
wRiLCL1A5iW3enDR5yAKd0JaAmxInIpbZNF0zhgtB+dooDVfGiqbDek9K6mA
kMJXc53eB8rfoy1xFEInTN0qmohkYA5FU9uuUlGZcWPMiWUzmEsmOgwFnonY
9gk/BwaUUH4sxRBZLJaCHckTZynPzsWExQAiwhRPARAFzEAm8N8FH6LodlTZ
dP8UgsoLo0eOUymqr/luauPMEXLeWx47WrUfxmGMzamlnkwJ6LzaivBkGfQe
uJrdWvv5B2KoLgnG5evCAmwAhBMzg4Cwd+RwZXL9dW6zPJlyxJLASgMWX1Lh
oTWWBH2h/9+XYrIe2fGBxdrUjPIIZ85eIFeil7bz5T5bk/Th3nxNyIIDuLVn
hY8/kK4QYsV4NA0xLEGCdk7SvpfZTkuuRZPa6yJWCCsVKLa8Y966b427qrfE
NqGfWf+cmJ9eJrA0d3/rRYeGF0An2BtjXjcJWZhDoajcfsPNb657bX2CJEdV
2A0V16+q3pMKrPuIduLyx2qRGFXScsmLFyZQAIo6LG/bST+SSZg7cLVCEmdE
RYNiePc5FzWpfMy8quRA8zZJXxdAfC/Da+Pl7M4gyZjaR3JUtXpaixUD/UnO
HxlTFYXq4wuir+PbFmhEU6z9+JT+mfDYPZgMNGl+2y49fd3B3AMXOoFOpRjW
4kDKfdpevp+Iv/0eSRHLc+xdBPfEych+ly+xuwzoOjt+uih1ICO/xS3KmIxU
4v1VM6IqQFk+pqzmL6wzVgAPnTDmN1ZSOoyrIAAZvJA0iTZyv5mEcC4OMqJ5
u8i2391FjJvs/Z0zowF3MTNm1ygNI+FeS4xRutoMB8yVsIOoqW9V1DtjJlQt
DcfAkxPRhYro8s1iS3uYR4ftBlmivDReRdesjEuF/FzvQFB/R56ZFd4WjbdR
B+oGzl7K/tfg9J+lEd/qrO0jzxU3wkdCi2oWLPomJKcht9uUIoFTXXWtIH8U
LWQeWBKhfiVwYj1t7Kv3xoQ5umk9NOx+xRUUwvb01ljm3PU6JER7cr48J/0R
dOiSA0te7ZbL4nx8QuKSlIPIehWAJEFCW4EdLh3fR+ZrrXKipaQW1Ftkleg4
udql/HT9K4XFyZcNUCZIiIx10XaumbO5RfMIrFwSrZIr0/9enO6D4oAw5wji
1YILzUpv/lcgnbytwrHHu7JbpbX7/fQjudswOs9pJGDIMVOke6taMiaz8WyA
V0gJXQrzWCEnlYkSTm9SsvctJNsGYpW+lptVEltwJrL0gowKIQ5V9n7BVvwa
ZiJkqfsSVP7bZWv5ubWuj2FeHp5GV8ZBC4nWErDDoUXRuptKr8AqU3uzPGFW
gdN6B/BhYysZ8iURCR2gMUrG+jgGWnmem6uxfglNl8YqGsm2BcgZ7J3/TjjP
Bx1dfWgKhg0eW3HcqGykxA5UXnEu8xg1tLYDjnJRFjKqoxjz7jVk+1xO60Yz
dsgxONaT6J4B1oC06sn+tYinsEX4QkCXiDnk8ZVsxZbIfhMoUZtCxk0bozpO
EqICTYMmTydu71nz4cueROnEPBJnr5d5QYwkzaLo32Og6YEq8m9PBH3pHbnR
bAUGw6piSXKXxik0bZ2HzyWk1fMZyg5KzFyu/7VX8IuGslkk9hRjwegb4Kea
ZSd3iHcnutOOvuflf9S9FRfsA5MvFkpudnGsF0wAh42jiCq+s05VsH3Y5gSW
8mdpr4J+dp7iXVaQZroPBkMj5fPL2uge02aHBCvPFCPOj4mgHlE0BidFcw2A
61M5C0HXImXNyAGFTLFCj3pDDnF0/LHWXyUlqIrn3/uu4Fk1SPppPXO1RwOn
Wq5Dq73gE/HSG0JililM+X0fPxP+0U1DRsOfKrddDFX27xNeIifEG9veZWIF
cziJsIkAswCdmXGSdWIu2XBQ1/f+UZ6HAkt752x5ypb2h2CJY43GhDieLIaH
ikQ4Hti6TwkOzFEvq+R9m2gTJvO3taKMKmHzpORTTCAPB6aCbBY2BZ9IVC/4
SQVUMAW2vx3lgWSYBEQjW7tFBlIR2YoRDVGPuqd08VlcWfeCgBhf/wk9T6P4
4N722p+FTnG7t8wXrJ4BpUAhBtFRMTFZLWjhHHvBxoFFSuHczHfDJy0r5zuj
uY2cC9Zz1BJJgAj66ucTdqe7g96yfmzfAafwiHdRWfDhAtDfvUDvsdkRcgkB
/nsaeKwfaK+wLagNeIDkDv2+g1litwNWqwhPZ/OdyIV7hmytwCnR1BpATL+v
Kax6krrcxDZe82FoIQLO7jOOm+RUwI1xl95KfCRWRI5x2QNsGb6R7E9euryV
vxZ6inEiKo0G1ArQEeT0p6pLDcSK9O9c9489A+lvhLy36JbDFwZ/tZN5CTcs
th3gRN8D1jCGPmTHwSBriEzkyHydZr372ttJVND3tzYp9R2x74nFGugKYhcI
09bu57fSi0+zxyJzS1E5bXNV4/7dv5qPsLNoTrhDHdq4NFqXH/WARR+TC5HH
XsMDxf1SyVqEO2xZcB0K6gGb4cWjItuzGGHA2BtZOpiy5BzYrxwwkfQ4kcU/
jqvyIPUY2pE9nMo5lYbx0PUwQKD7UL19zfjNAt8XxPhU4Wet0SpiJ1o4W31y
QAPUBv7lMAg9+FOqiiMew/YBDk+phwPRNn32gYf2DvBT9t32n4wz3a5WrlTK
mTMfPAXNgiMWQELqZjMN3L+UsvvcYMKGwEKAI4l3s1a+dNLB2MlYzTgolem3
8pKtVWWa4CycLpvTAMDG+tjK8CeaZ+RDluQMVORXQsHh+F1hhEaVstX3pCP4
opvtDS4yZqtJADZaR5uXOHoWJfexuYvloLgOtD0LMhutnuELsdheWm/8R2oX
I1pg/QPKKz+KOdzfoUynqbuyaxnzWyX/cNekR+JEfIEJxs3oxcn+gI5Y3DS0
sI1w8HWWziDbfQ7rMP/AhRoOaQ+OI3oX5GOOz2MU3Jk4LoNh/ZPBNu1VFORn
YRZNAnkNxV6e0tUFslyKxc64nRv9A7A4QK7dQNs+mf0qKklwUgnS3/u92E+/
hP9TPJ/TNx2yYf/Lpbg/05He8zvpwezVrgMPBKCS3WYGfHPlg2vhVcUAfK/l
RmGZjagDP8gwl3yKiBhTVGezO1I3VtEUO/Kx5JgB5mgQiu5IFMFffDdjim0Q
L8RUuPtLxLr05LF/E9RwoapYrwydfbxwcOAOi77bKboyWZ2gCTScMMOrpOBB
iLV13qeQm5jI2/BRo8uImWeJVHH0txv8Z5OHpi8bVudt9QrHtblEPcivlZHh
78DhMCVB997mN7XcAYaA2gmycEti1wWMo9hpeyNia4m9vYwi22aKcNlWs/BH
PmxfAHkrZFeJrVCTdRUDurkGpd0yaADd4yeltMU1DmVQqL2zEjQRtR/t9u4r
yjnpfct+e2F8KjP8zg8t9ORbZr3+th1BrFWrJ73lmXCDR+Xb3GfQxQI3leHn
68t6zJjgMS297fBi08JlRNXrk6oj+L1dweG86tRiKc45jcKRlyth8VHWRvAB
ARIKQPATRRlNqRSJyWRd59H8/gwGN4Kd5ZtX/8/fqDD/qW/kd9eqwbfTZkTJ
43NSboRJ1ZRk5+bZwTJ8X2pEAgmA7GqT5pEaO+hoT520hCBysgN6NGONkoOo
RFvzzEqGsKjHW2efGCU8rpnS9Qfidc445HG3stW/PzOXHWpn/ref+PnEo8X/
USzJwFycXYx0F4IzCLTGfyep/wk8wEYG1GZQb9yeytCWfUVClby1d2uNZV6y
f2nkKiY120TUrAT0NghGiAFYFXgKtD1a4Ip2aPSJHx353XYlyaOgbPZlSkHc
UZXguufYvEZviEtNAqKzcq6E9d9pxizWUfdUWKxFNvN7ayVqhMz3gELmMhCe
d5RrcKGvF3v2viUdOvktaCgkfavUNyBhFFzN/vdPcFkvRhWZXT2sBnNNCR4B
nHw9UxFu10LD3HqbXDwUwEXFHHPQXQnhcGChfkLqOjDRXqO/N009qgnw2dPg
Uac775m3cow6deIbRLSrqZX1nfOcCBelV7XUwAo8tvFsFbQGRCc77XOwIbye
gvSTEPaBW374vbi8z1DsGzrJxN5ECQ4RhAbdlyWqpEnnjC7udGTkAdhgmLcH
NR1RtTNBltowPNfwzoQ+6LGruis3FgNVGlLOJCJUw5wTuRIv0Slp1cjIEw2S
bkzijtll/bWEvUiOOta8nB67rWL+8K1U+8vqCmfZDE9qXEaCj/lzwbIbwl7+
kolpkOI5+TXTm+D3FWXTmX8IeFuPL+xstezJvQNOfKlhO69EUqIFleBCR7L9
YB94swjV7jExIivAlaXwORn6/XLDYrFoYWsssXquSSqcJX0Q5z8aEHNKESER
3lhAUuJFrJ6/iUpyN18jB51bEnJtd6P5Mp06U1Nm/SDio7fJvxDA3JDOwPBT
om8AvS3BD6n3fCMEfvraSfaDZKeBLmau13fp20VCO15i4wkM7yj6v2N61uQq
Jee7+Nqwp4y1k2qqwIIn0MnjYTgq2TAkmQexYia7i69B01Q5mrrytlz7bWEd
aJIn0/lsNCE1c2esiWsUhft79uUWHE2FglJoR01Js5rpXcMCPuqnrh52nd4p
8ylpHtkPhTDz6scVrqB+pD9TlEXFaFxButj1P2llpOdgUyl2PBVqciU5sXWl
h/4EvLyvaF7x62tjIacrsf1nt7yuqnfDEl3WhTen/jaj/nzWhTgBWyCsZWgu
FptWsiy0wUzdVeEvmNAjmxkCzNYHN2/aPAr+ycvyRPfRWHVKU6VkTgbWNQ1V
IWDYTr3KuJO4PbqHQ8IPxBfTQ7jo6xvKDr/m+Ymw0TtZVR6MBhRgVs+ofy33
XwF5ouHLM3sUshJKX3WVWParOv7pWbXcQvuHiBD9BKePkyEa7Gidt3Zupmjk
/xBDLxCniD+WxApdDWIAhB5tKunGivMiSVM6HpLfmEv3eNf1Oh0puZXowAm5
RbTWAjJsPZbHB1PJC6m7g79wtUYhq7EQDL09LLleB+KMdYof8G7on8x21eM8
0XyLc21Bu0qMIHA/dzwdAQeIfQABDSJQCT3y8JGR8IHSI4DhwfnMxD+RZsRB
20Cc26HjB+tKQkHsQKLZjp2JvRGuBPMj8ukOD+tpmn7W45VtG4Omk+qiSfBA
11Hw7QHurpl5yM8tgXF8lv9KVFKWgZw+PNOkMKDWeZXRJ9GHHaxG9OQmnA8g
IklAN+5NvI4q6slU5KOzlRLmUItpx4FrhKOYuqZvy2ga1tW43U3n1HZ7qAIQ
ecqb1FS3X4OCWXchZL6SPFGJmXjDYaUdGAZmZP0dm01XYUBwnppPxcbLq/tr
gFu5Ddr48HAj1w1CyIVE+tw2Wu6EXPUdY7LZBw8ocKlwwdjk03TrVAChXLxY
/Yhvwk735273jEm/l+rn1IhrG/JBOO1S/1aJrPFy420SYubM6e/n81s2dO0W
wZx+mig+hWvT6dTqE9w03kwFUhh7k+zib7kkKzS8Gi4qQvFKK6ZQJbDdYGyG
/CiJYFg/Lav3+OcXH1dtO1Qkj8i9KE+8vLToX8E9IJyKtqVB63eJfIPIA7sO
De7lgKKT24y8PCLCLybeC3sA5YZEe8k0O8RAVkjSlWYf8zDjODagyTWHItbU
RfDPywqp97ElzDR+j0XI0obV3Ij1/p8Syj3s86ssn07KynO6AHLpgk/4HLXi
RNjlHO3npeB+3zxcUejti6jTk66yO/eUTy9/fXnX0XhMt2+ptP/cvLsG8mB/
nd6KBe8EyPirnDh7YPL6wPYQ3nTk6n7+nIUcPvkVImj1ibscaRLcu2w5qSzX
B5svSiogSohjyHIzvTMO15FipL5ksWwLm3Ea5RVJwlspdlRNtW2LS2pdFlCO
NG2Pz4lCMqhWfIUh7UEul9MEoZEn4uuPp3IMZjb41TrGs4r58e422c0JtCkP
RmS63EGXrK1lSyc+GUik0A2omFmD8GGOS3VgudHg9vUh/i3rfFZvNLu/egXv
k9qS0MqOCZoKvmnB8piUDWPK4nSWnGseaToJ2PJMa4NNSFzWS4RWoae8swKB
LsBhUiPBgfrwLfIrzISNCqBZGkAD7ROfmwpU+a369U62YR6qjZ5QYA7Suetp
SWD8QYEnkLI60m2OHNJuHTIYTbzdVIbrJs14S/lhnFLEFdkSUVLAacstsulX
gIikEUpXtraTzWU7ulZEvqvETSH4gROvtDYyZjwTgr1hGhY6gA8xwrOf85hE
MFGrXXeaEdOOJOscydPP+BWNjO/oZGw59Zu+gm0Nd2anJ0pIv2xhZbhLDQnu
tvgv0KwWMH/3Cp1tFJA7XD0lEdsNgRZfIF1qpXrJR1Ntb6UPorzVSqdaefEC
hyKz7DDyyxFLzF2pLDEC/+9P/S740CjOPuaR3GafifmRijJUILwMJ+kzhy7m
1DMP0sKZTnym6FCWFIB0l+TeoKK2xBfCX3yWIfdO8isf/Utmj/uaSfsHnn3M
yD7Hw4wkxaoOHVvX68vTcbg5m61MqeSsnqkAaTuZmB8aDHtIp9zP1KzpB40J
26dmvvT11mPGb8QaMsggFqR4aNBg2X2nNACaxkhrpKc6MHAzQ/rVvwgHUefE
qidhWXjl+hxpkxxmr7LAzAzsRT3raB5NWaSi3zlafjVPdrF4mKiJbNd+2HSv
iR+rDYIGNq4mv7rNClRiGN4itxL4yoYxCePdaaw4ChRrJ/yg8en7iLljjOgD
wI9UlUUWyVpekVBYctYf6P4U1tOTRGx4AsJyKN1NmLQj17HoSA5vS8TUKiGN
QGii1OCy5IXEh0VTK3QqGEVrDdg6YTFHRxg18X2jJnCQSAzK32rcK/iPO1SR
8fKh+FVCyP9dVOXod/eCHu90sxnv2kpQAMGvn0H2bijDAWeKHZOzp9uEks++
HjdOcuCP0AF8K7AKi3n8cmo0/ccTT/tncBIdthvIExoQJ88wS6QPf924noIs
0a6fGhrXdQa/VcbheN635Tc9tiYwXI/R298AY5XUEMSgSvfc9E3nE58ieAuv
+t8BNpTUg1aOE+sr0Ugn0BZD7SBY0i/lH9WqRd+XsuZ6Wnw0NabRE4Wp5SfB
k/WAYfhCvaKOKeK6yC+IbsaHXeK4WMtWeKMnHn9jwkVPbG9PtooZpEgo6484
dlRaisKi0sBM0z+j0HRvyzVc9zbZoPZK97O9C9iL5J+19zFMFwDbJSDxc5Bh
samC7x8buiyltzMgg/2wca+fBFKCDmZU64l+yHCpLgg2+fvWQKzWlSWLR22h
sXb7VAcnthR/RIie0+mZau8FJTrTeMCyNdaUUr+7QStqRxXP3v2+ftCWxczi
L6U9qkrb8MGHWFuz3JMrQB4MPeszrRGQ9eqf43CnJZlZS/b5TIFrO6/gDIyZ
NOj41NHlk5c4ABSOlVvZA7X4g80RTJ7szG8T9KvMEqMxAOxYxDItB/KglvWt
LLc1fui5MrH+nNJvhrTbgyvwANmo9S1k96aj8oRiEWXx/TVsBlih2ap8Zl2a
izKZ34CY0mGj8/ydOUZ/iGzc+RUil3Z3QatjF8eCFKPfohEXMUoauJntVIOM
nW2IBewJJpmNfWU/lzxOdeSDMGeQWaE+sz1LYt/GnFjH6VX8UhRQuFtpeI6i
6DbOlW9yhC58A5JHrP7syk+v2qU3j8jyhw/A78AXvcklzKXQcaihWxjSJ9Kc
E9BwTrLFkndM/OhgAQAdeZTWtwy5LMX9ygg1c7UvCxAk2+K2cA/eNq//cASJ
NG5WrqOv1w9BsnmXwH7KWjJCY78ecB7DeIk/SEIyUTuw+y+cTlQtSIEPhqTB
FHrN4RZuYm/liwThhq5mED4IMQ5Q92PcTyWgl4qwksAZTvNiX0GcMu1PP9+k
zf+UfctSyoSAg+EB0BUsfzhdT+/xX3NBThPYwDXHD7VCAzp1TZb47OXw1tzb
uubViybcxWFp42Veg0Ndljx1Uo3nkjB60HFZkn3fXhzlpdkJgVlIIG+Rkik2
gqWYl50NDjOLkC/dUBxk+2g34NqKW+6NbdPgRCm6Daxqbr/K6EtFknCeXaY8
dYf5gI1X9BxBU/j2QCKUQi4OVcIBql8xfziH6B9Ux8mwiXvFmMb4AtxqesJ6
93O5jk1w4iDyE//vRgyx5xKxE3TvrjFNvkXtX2II+nY+jRr11MLvb1oQlOsx
XLln6Q3bH9BBuNuZORaaqGgyd7ZVhNDRW1ZIRIyOWrlOEVUGMY+G0YGnic6s
Fvi3BHH/Ey36z+RZc4crVkDbBtV86cCBbvaJ+TXquoy9AIwaZmY62onb/GML
HoIcU6jTEavBbyoiY2Zog//fUXWey1jwpKjK4WqNiH2PFLzcP/O7Khax4YOR
BKtHSQJyAnNQ3WYhA6axmdDDR42POdNY9QcYLrVy6wxPgtO8k3/ATCn2u2Bb
kGRj+VOt4oxGJ/z/rTfqj7KUW9BejkI02g42NWF8N/0cINy4dwNqXeOyqvvB
+jxDfIPVut0F5sNcd5J6sxtEXPl8oIrLS/S2a+p06Q5ImDRIa09l4lvBt9y/
vQeYqYfChv3UbHy9j4EmUFsxHmuYAdFPGEO8WpVvY/IDnFQ3d7DvMm3hA6Bt
9UEFm6eIMUpEH+FEKnng6CSM1sXLTyyOCD+5VaJf07h2F0bNFLeSeIQqHWAS
5m1o2ObxDdCYu7opkQmvQRTuDISO4uQQsNEhzkaZqw6TdWHRgKaFSxFK5w/B
gboBDUZ+ZMWEPEBKklb19QkWv007/WhsdroPQ+tuvuTe9rlgiOBKKahVpeOs
+IoXpuHrMoJxrtJ5+872tA7t1c8INTTZObUPhcjJ9mHqpH4pjHqszdH85mGL
0YAx3Ymwvs9unIrWW2cgOZQZ3z7WVuepHjSfl+3ctqSVFoobR9zune1BA4eH
HroDAsvM0kdS06Z2+WBpuxlAuWT40zphlvU/8YeZj+MT7jZbEl0MEl1pZ8+P
dcpNSnbgr6HjhsOsjKixE+ekllKBkuhiZd6GKyIIfGFeBJiG+tVNzAvpv8Zw
AgF72jxLUUoxL46kOXO5NUL8uVKSINqbCiV1Wt1Fb8nA8JYV3SV1t+z5rkJc
t5l8Zx7gbYaN2WIouMUYKc3WTbrC1n5R6ju6sStA3LzYAbJ8LpGx4ul1FbE9
skMqRTvJeM7Q0h1A2COZRm3Ks0O7C7EG7FylIiv9gaBWiaLWWjrdqnC8E4KN
2JtQgwL1Suwxni3eJgqDyy0/DUYlMZzGrw/lewj2FqN/oqNDRoTMPLREa7DT
XJ06luKvqZ3/iBlrzS+25pzm9IO3opd98tDVWGDMw6AytOejwtcHsnWIpMd1
he8FJSR9UJ4g7mpEr65h3QURhAcm+wH0wauCa+ZwCIMHex8aW4Ly6okFbs3Y
NrebFNobyyQYap5NwpjxAVoXpBPpVzc+QC62868dSH9c/+/XGnNxuKu2Q3JO
jT6zegJcLVyv8hXqscfsH+PlCX6HkzsEjijQnmLqF8CVbCRbTru6sY8zxljj
PdHVwKo0wV2gwA/M+EA37YnErHfHyVEPD9o9j37pwNiZnDyM2f9EOoIYqjGh
iFGwzMIya6o8mhOV3adHxfa1b4H8bZ1b5rNRebWgnVIg3ELkwmJIp3y53jY5
jVFUCeJ/sC7/xpSQy8dDFNP2foi1xC1HYf6X4Y60qdJCHeEHkqUrQ9JNd9Ub
PXvlRd7l9DVJF1aQi7hMmV9aQaeQ9ONEzKWMB1pQAsNjtolIOsf96vjwx1Mn
Bvsgg0ihFih4/L1kPiCcLpkz7MjUHoiubOjiMckLwCLh9MM4PXTOhCwVnamX
7azSh+mlHGkqPc/niIF5qC6OjeWREuO+z3kMzWJzWHV/JHPaeBhOOQWFPJnB
rh66Vm/Ln8RfwdL51G1bUjLx1T31RSszvpHhPDZv3UmnuKCsOxXHe9MUfFFn
9EP9Nqqc1dpktWm5UG9rMY9iHZWvkGfBX4Eb0GRjZ4XPn4txYO6h7QXOg82M
zEyRhE+dSDY28h8zUcGmH0LNAgU7wnU5622qxIAaCEbaKrJaNJGqJwsYGwOP
KmffKPfkGQoKXGk8VEh7DC3IRiZVMBSN/M25ci72NFPI0RBcAEie20YKZQfO
jgSzIq7zv+DWcVVgEi/QCt7OMXwgq80ayjMHCxuU+vqpEaI939Xh9+a9gc+8
73GVMebFjYXIxei5IrTiAJ5KxjIogBQaHnPuVTKAi1eTTUSq4HIMqWcHYVPs
rL8+dFOpznz9PU5c9R4s4tOgbUsRKX7tPRy8oxFwPmo3VMYhHhkA20qrbAAy
9QcEC9WK0RSU4t7OJ4kUL3L0jAmQKCLBVMABXybDMq+pL5gJJYHGCbjez/bA
HqSnnJO46B3dWZ9FOY957IXF64v9MCeIrxNikKfe6kkLtoYUEicHRaMcpipS
XNHHPsogrAaNL7+UEs83lU4OqJGmT3YgI8zOtwI04A4DLD2t2cqmwfH4NYzQ
vNV4hht1IvE2dOelt+DQfuhxoR8dJ/ZXY2JPlXDWdN9LMVaVFslDI7kqY3qj
5ckLlZvAZwNofUCoUP4/QFAV0r3UUMcycU3n814mXmTx0/7QqqP66vT8xjKY
mKVj3H+OPjdzdRZoFex0Xq1zpVdzcJkqFXNxSDa3U27GRLqhoFLJRKuB8ofK
HEmzVHfRf7wp28AiqAubWlelDgji8hzbmHZb9FrTXWJ1yS1PDbmBeEcKOUNC
bzfHLBZ/SYXv1SfRLAzASrPY7pd0WFHhCuA9IvnsYifZGvR4goiUD5g43yLn
H7BAoLll5ugVEW9670SHOVDXZ5MDEeJ8ftHuZfgnAoqAmL2BEh05P9fluG1y
5kVpZhuxeFjTFuZy94BcolHGGx38CRnPnHCsYfoKu2yc6QbYKEnTuBiyaWuD
CGsabb1wY89WG52WLk0RTcnSILfJMQzO1KyTLTLD3ibGpUEHShpRkBSKFKOL
Zy4rdO5UmLrkCtcxhjNTM3OJD+57yqRMhGUJwvIRbooSyrRbxokVOsi8JYsU
C0qZqCQWi5lLeYQuZ5OUS80065qaPclBnymCNfns1X9lliYUJCo2C8UISeMt
EqknRcZHBCRtHfRNwjByjMRQIKIUxp/1Vgtu4UgrxKlLpB8HLF01s4j6zv7J
ywZnppQbjqnoUoT2wBXRfvGrfIUH/PrhVMefHDwgyFYsslFHZohSsaYClVUa
dgnRSWEGAfoghKjCMIhsknKzm/yd7V4NUOyqLaS/IDXcw/Hr7vAq3RH+I1La
n0NvNHWW9FytLuq8av/Z7svO9Ax1lf8Ta6jBuARrBzzIYeGFYoGNAszgZSrb
axn/7613nP8f0vmcrn/B2gylZXUmMXDilrgUTdtuR1mNitVJhKWUIkB0Skq1
4Wv2NYV7LK691sQ4kRfjVy9aUPF1O/rg16bLXTgDnQRWINN11tUg/ZZHneEF
O+ROS3HusTNqVfJqHo4xV3BV6o8iAKvPYJCHC2kitoZm6VEUiklH5HCG2o3c
TMdapCh0sU23zjtXiaLMR/cAl7GbWZtxQuCeIpK3s/HPBE7Cum7vGNoRQuO0
vsqVaAf9s5+NyPfaDb+oQVNyVuaXHKObtoPDRCbroNRCqgk97EnvpYdoDZei
60IY/a8A5wOM1GiELVeObqr5eC3z7D9xgwpG9xHf7YBd2Do2//VX8n7526IJ
Yw1Z0oKCxaZzzaER1HwLFqSmu0BYsfz0Cce6zp45xIWygFumiNmHNNum1AAr
nMIS0RCM0/OTbcxNijb8PSJJhyl+KzXFO7ImP3iSx6FffHAdr1x9Btinr4Al
2EHvp3uoFzZQfBtkNSD2NZFuOJWx8L4uH45ghInnOhIAGjosHimzCGFYgt8N
oXt9nBG7YgSdQzIFUtuQWQJtaujGl6HNo+zDc7KLB4zWYqoBQ6ZPYX3qWl7P
0VuT2HZpQOh0ISzHDbP1bCU0xEeCoYi+USyg+uOh7bxa+PJzC9zp0h4bVChY
3pwzHExz8rVipF2jg2NqJ5HRwv3m5P0uefhnqfWvv6PaCPE7ZoDjapdEqA7p
1IJd4Hbdd/axRVjORWr4eTwu6taUmpkATj8XvcmGoLt7a0s3SNDHfxYvGKJA
4EixPDOjAA7+E24wNWsbxs8jkdsDWrUOgufIQDKkV3ozdr6ZDXbpj59Sa6uL
aM8qXJ843p5Aj+aWiCU6mX0L1NjOVr8VHTPKDZTa1A2H+5L9wONUeO9JV41R
wM493EBYoBCCkrkCoGbUtjJ737FkLH6NQI0v8DO42/3ahIAIrLSaazma3oQQ
hR1HbfkCiWPCnaF7vLpJLUwglyu+qBzxICfrERIkv5TFG8xBl5zbs5atOhKw
nS/2xj16FiXwAavv0Iwdcj+mON2jDWO513clp+pGwrKC9VHwTIlu8PLeryqC
v9jhRnN+HG6m5rlO//3tN53HifLfkbShJuEczt7LJFAZTRDR5wz6YDbHnA1+
I01CuotmfZ4QvdZYIDUxIKDsuO7VxT6XAlk1JAjsb/S7mjElatXaYvq+3Dte
lckhH8UOI25b/naZ3s0TYUsH+Lz3cGDu4QB0xYdQx69zqD4/STwP9mRVTA2k
AdyAf/eUUxNrXyW3u8lQUBiE5Yp2jbtSJHqeL6wbp9htfOySdyQvlVkre/LN
5BQg/qwH5C9fN+sEHi1rEXWwiqURUk0HiKAO44bthZR97rcVKyu5qxSAo8vz
PLfFq0wauExryxa95ZIAogsGtzWm2TS1sLf6qmjpo67NumRI0vgj+/Lbu1/D
zcUjVKYxy2m1yXbLrcLKqdNV8KawN6jMb6HXVJ37288UOZn9gNTdK/rVdltS
g/DlqZ0z/DInajwn1SkcGsN3e+j4zs4IqGUCGvJbb1mcymqlZppRmw1Gfpg5
98yDN4ZNM3hyhj1lplj6BIB0BDmQ2Le9MoBtMyQAfl4tfkSPrIhauwSsNwrE
btbhIUsYyQwiLgd0TugNuTZvIat4ZgZfYMBGHFjtQTTCANc9N5ooQDIrYw6q
zKzG1ewItpayc36EY6m24qsdbiYXffQLQHep09SSaK0EPQzTZLm7aqQvJ8zY
0qxMEwUb1JfVIiW+pxNILcCYowWyAGgVtmut0silQKnOihIq5BKqq1EUfE9s
ejniwbDDk01S9xlLQrz3PD2jDRJYG8zCGFZgZCtL68ejIBr3gCe7lma3IdYA
Fy0SKblI91hVig6AaSfbsSN4G8xCQB+M8nP1dFmK3CpASm+PV1r3SCON1A80
nlEcZ7nPOUE1ITx3AccN6LnZPnlqcCWYRRaIEg2M2X3rwH8TDzeXMOF/HQyO
AZUH8Ufzx+zmpiwFZVPQnEMD0DrJxQl3obMDFaDUeHMRRelu3OgXkgqQUy8v
dPl4BbqClCLlZlQlZ54lV15asrTrywWsYXictNpgWQlHlPqUAm7OC0TmqrVE
W57jXH+xWo899sIEIL4B0+ZreMOZZC0t1LDPom6OCT8PHHKUAFwfz5tZQ1lC
xcnN6hEs1b3TxzMvjv4kQOxf8i359VmHo2FnF+FJTddUsiGoAoUjv+IEIFIS
8bjhqNLONqzLFq8t9d7C3xULAziB6/dKpm2e+UT7BWy6siB2BsuhHW2E+/3V
mQvEnF5KukJus/FG0HQlwGAJmHq9DyDn15OkkbjMuuYLIUGEWQaUzCE00DTt
Ck8B9adsemXVcG7M63BSveJqLNVCD8mgj1JiThClvy0vmOhj73DVx9w4jzMu
MRguUcyZCnpVti1JD9crCpkiMCAa/3flcuQDXJ83o7+uiLllxpQm4gJL+l2y
dK5J/mT+YBHTS9dRGvGfo4UXqgCL4JPOL0b7C4+GRibGL6ZXuTz1MRCTs785
kdfphdTCQTf3fPgs97XSfSEEfd2wolLDxF/bu4GT4nZw9vIG8cfgeYEWEs2m
vIH+zOASCLbqlrjdYr99tUm9GeY8iHj0zDFPxhyxNlKkqJEwo2D8qc1hap2g
0rpfbddyCoVY5vkzQELJl7ux7awQbWNWUyTvKjGL2wo7Cj02D7XvT/oJR92m
AR7m0w6mj6QnstN0L7Mc+YHKhyc2d42TsfNtStVubJ+IEozbDAKsdqBBe+sH
5Re7Bbpk1D8Z8LYLURq1a/dl/+6rWr5juZLjG39QmewAHjPxoxtznoGkycjh
JDae4hGhZrhskll6yPbNaVaoHPMr/ZhV3t7AbEVqRP//6+USgxjcKjdiQz/Z
NDz8n0pT5rnQMr3I8/yv2KXzSLbdNugdzOI0GXINPTb4tkPo3zOAVPa79S7+
VeV5bwJnHbg1EX8nPU9WRRmpJhUO90nsqSLASjgog3HZcEioOcf5fdBvx/zl
R9faROFyM5CvNl42P/dSlrIPdzCaPJA9co62dqkVGyuE3YouIUkfJu2DPrbp
4iOspUDtEoD6Tga0ui0SEp2AYb/hCKMA0p7e9gSoYjWKWXdv5rZgQWq68kAX
lnekww91zpGfL7pz25Vp15lH/bP++zG1w+qOxiJjhhzE3jh+r6hAbmlA5dz+
dGqlk1AIG0cVo6SeThULCcmXgbCKXe6ddJ3X8dTbk54U8slYr0ZnAUbvtxZ1
jZOX4iNtlfvrBUiHb8uSNRf5A7WrE9sPPb+uuTiqhU7Bm4746RojeXTSPUVR
gnZHbjFrAr11RIK0oetZQH2xh96rgABAMh7XEm819E/6zNYJy/ZQWrNVlHV7
jBvG1GHliyHiTgoBT3LbqoD1/M94J6+TBpZJ03uSjqXO7etDtTlj0YhhDbnQ
faJ5vGQI9mWf18KLHHY39h/aBKeKbOoLzwqOkPZTCw8VKFSHFqtEGCRAuj6S
wVtZ+cIg3b+dROmaakJQfleASZwuDpxmeQa9ggPky3k9ZZ0anNRgL0bv89DB
QEmifQywJQ8kfRdR6erRpl8B+I0txGWtjnWt7VUevtBm09B0osSUhGjvZv3g
/c8vSebHQVFHTBV29tk6PmQu+xBJpxbNg9NzbQWG/IONofZMHnCAqlWzVEXV
sL899/RVnOMDLKIT6vdtEk/Nju08iTE7e0bhan6g61l5lPF/zCvAbv1OOk1W
yAKzppAfiWQ80I6Rr3LkPmCQZqVew0a5AQnnxsNy/P4aM1Bie+ACWK7kCkeG
M3dNZ1170aTEzYDhbCE5zlTnGLLOEfAytrnVa8TXTLqmpTGlGDLg9e/JPZ2t
L65PZ9BdYAiu1BG1htXiURLLY6tVUkYd3EpFOz1FgQozYFQEjnc7ifjhuDia
VKPD7SddPRpVccZS8LI3J0mV2iw7WnoJsIYzItG2RTEsMsxRDV1OvkxOb10h
mlrBOuk/eM4GskdEMlHYS+Qwc5aCKhWZ+0Z5CRHWW9JkJpkHfy2e1IA2Pu4M
EY2mleHWPBKoGLOOUCoVo9idV1ReC94pTfwj667VwT0LOL5fPzJGw1HVjKoi
+zf9fWgwyu6yPhgeoh7j+Q6kXvEb0SGHeQCjQA7UTjKqTfM3jv0VGJMh9HkU
XCUQVH7DEo6VHH3jF09k1amT0jbswl+aEvRwcm+SKM/RDK9O7qtc3i7e+I6h
1a2zml3V4F5InD05yPhYZop1VwtyjUJ83O3Rwwg7lKzROGt8sSrqvtpIvSIV
kiY+dtIQWZeYuUMY/+fee0hAJkz3kojRc6I07ZLXlQS8BwNR9xg9qHpaZNFL
qZAQivaiZxU/vSWk5H3u4ltks9zBqra//coyq93sl6yhl7BTsKmWHcCGOfN+
aYNuZzqfXnO7dgYzRhJ3ZLHTR5LhS5gQBOcXAe8hlaot8zz/GU/gO94phADq
pnlwajhJIlpK9Ab2kL0Tw7QYGMSwyPCMPr9NJWuUjFjYsqa70hqjq4L55VV4
vBuI0JFBso7e57M3gpRJv+qQOX6eO7J/uHVxRGMqyVXdHTGmYoq70P89vBQc
7Xl4Yck7qvqyVtUHenXw1nGuJvZCo7eJXu6EMQZPSiWmZa3FeYZNeh1aq8UL
sVxhxMylCopjG+doNR3fOFclD3bTaLc1kp3kpzahPgU4uPx+Hi4adbfmdv/h
4l6jpf3SXpIto+Plp3ARn/+laTk/rVs0XlOz21zpxofc4MEkizU8cRwSTmn6
eeu9in9dyhT62ZVTwl0dVRVmGMhrysaEAy/z5qd3AK43bpk9NdjNCqXNM7aK
9OU1A+SQrJIbwPm8j3TyvMbIe1cA6EG8sle3QQBOCgLSV2edQ43o/lWRZfEx
Yd0N6JUjhfJQtOvYEgrYfzlBYVG/dFDw8sMWjd93mSt9TxJhyi+hjntP+uJI
1L4poI+oiuzlef+11WjqN2YUS5GEwuOPXVJeJhGCgmxAfk/6+UcuakYeFGaZ
EoVhyd5PuAiFjXNpDCnvxuHDGQnPKsQaeTsBScI+q3ZFiABNAvXS7fwuXfmz
BgFX+KwSaSvd9nejaXDdTLVc8VX3XpJYteOIEWD8Cjwexiohd/VQO0RLYrzN
xaEPXZ5Do57lJ21J7P+HVkPodsfc6FfvCGUw346sOPSpZ02qL8dgOk4oIIXn
j5FgCoZAEzOlYfufxco+oDYIeGajICx1BI01L7KwHyovPzIW15hAnyUPxugY
quXsdb1z/zB7pnwQXo3EmQv2Nm9CwmccOjae7lD95RRbdYeTld/Jhg47P89n
Gz2UAZzp+Yhi5HJ6rHfQ2tbTXCNm/M9yjX0FLjXquR0vvBPNzmpzJStPtul7
NvamrpnXR7RrYk+rvrHTgqYimr2+0KOm9gWfguzyNf8fmFTkox4f+arMxe/S
lO7YV3txFQNbMnOIAiQMp04V/SRY0p2AEHW68TeVYx3z0EaAxFlTtssipmAn
RHHKBDzVYMKVeJsKSGxzKkUMEiVbpmM3WK9G0BRv8fYElpT2LVlGLyr8sY4U
XF94dqid2yQ0vHt2EvDYlWuo+2WWriETWL/60AlnGqYKfykovQ/alKZ5eRpd
0E9BA+oobqpSk6O1jL19eSZwjfakXeSodYf01GGKYmKJK4wQ/azTj9PymHML
7MYA8BNiH7islgAvmP8i3IShXIzlg6r41HgDkeFfHiyjNYul7bqM558TVdFP
ncOhO2Un8RonwK2NtcyoNVyUwYyx5HQ6pkhMTY51HhK9/Ci7Ui8Ywo/OlKZ8
MJqwJHdT4Z+1UZmzOtbmHU61YorPcbcULVIMhhxUnC7XUf7vIVNf33Dv4JPc
K6D8+qANOplsaba2evKc3ej3IwJYRB2S0KqlzsvIh4+zZDmGwrcg5a3tgm/M
SJF1jbPVl7fWloqsUI/ff6qWeb36skxIawPGa0d9ha9J7F/ouC01+5Zq7uCG
OaRXuVjAgxEM8Gg0nvicL3p8ruaEOnn/fIulHcvCQzKygDzNouh6h/ZtfXx5
b0WwFabtCx4/esZUgackkrW7IxwlLVWdnM3bHahiF0uUU0AawdSG9EA/p3Yg
uPYl/hZ2tqYUOsTxijNBPracQuGfCdDF7MVFH694On7UkyRaxf88tMZSO430
wBmYhPXxABUgsm5+hQ2LPKqgolxH7S0fuk7z3a0oiPvm8bTF1LvLj/Khh686
JY7koBs/0PqSc5fyxSXJn20HjYc459J1CwRBZEvyfBqBXrExrZ/bAovKjDur
DDPUyE25MLeYEQ6xTsw6UtUBXYkaqX72dZp9EBMROSGXW3YycCnvj7czfptD
YvxQXI1J6ogw3MD77UIj7AKOZwByNNHgVVi5PvSotYAeYoYCH+QWApncBvVu
jwQUNpK3QhtY4OOsnalXs2mLzclQBEheyl8eZu9CvvX7ERnXi1SnwbThFFiz
Dc9OnplB9xBwg9VTKBHB/sy8w0JewsnufqDdrJY44NwteDEPCTpOUibjqohi
Jit50nbq7fKpMvPnslg8FWJwo9rphXis6J2qLGqKfY4/Rt4HIef152TEeEaA
XMmuk1Oix0BIPqqFAjXuzY2jWoTeqLwB/GTNnmm6dH18h5/sTm/sHfsABbGx
flEoWYIodeGxmPWhYRbN7jKOPExS5uBbihuIkDqSHaT8vX+Z2XAP5sBxFAU8
45K4gt502sVw46qwTCR2OxKvLIYC+evOXzJ0bW1KoekfrqErm+umoV7aK1/b
6V7vigFx2oxxB0pIc+5L6nrMv8X6hRrOg43cqVjsp2Z3WImgi2zOmOZfsA3a
40tXzI41h9GF4FGdAzSVmnIOYbGRXETn/oxgsUy87zaPJB4U0NWX1FBkHTtG
a/z3lHVunq9U4y7j4393t+HMDLgxYzSp1qtb2QN8Y9bCaeKYrxOmUIwZu+lo
9ojVxcyyVewMsd1y4No19atOi7rJ+AbHsHrCxc6ceRPFnAl+OPKi1diixHnS
eDZls293p2bLSO80xjuD5GHJ6NPGMHOW80HmpDvFV9KDyNTNxxAfQ4UH4KuM
/PzlRcgUwK90i0NS5/ymjnqP792vL1b+SulckC0qX/e5UWCowP8YknoAKoeJ
3O+uqAvPzEjQYgpgc78CKvGBtr0rDRke1UmhGP28twkLV9p9HWnVx0qKYD2a
N7WOT4IqoyobwA8G9JEyJMB+vnOodkU/zBFGhjzjTX3vNJADkAsi1k4DTeB5
ipk1rzzuYoo8dPEiGx9nzqlL6HL//ajUkWWDYGjOu7PhCfQe1cimPCmttBJk
aZ8vf5lKbzl9r8zNXB7uo0i6rHn9tLNwLQSacqH9MN5ejzMboq1eWgfR9suY
dRdibKJIf2010l7GDAI4YoEIFil7utNGeVWHIPCauoe68MRDJqKbVZ0c4LpU
rdLaK62r0MN8V861VGNbqsb9H/JH4IiAZdYkVXuD+Wfzg9AeB30zgmST3Ia8
04F5Hxd4F8mltsWWhD7r87T9B1xAJKf30Kh74anT2oA89Okbg2n9vDNE/MY2
we98JVaYb9/TNOHx0w/CIsfV+Ch9X5eYxmBhROpCoKyZXlsBkS37/Xv1DnKS
WByOije0XF8MQ0cRevnAbe7iFPMUIcLlJmxpVT/Wj7i2EBunp17gpiZ0ajNO
37yaa4mb73BE6MU32Nr3v/wVdMGvgN/KyfmZCSbSjmISrW5MHcT3wCdatpee
7QxzcEMjDxwYXZmZ+x0QS6Ho8+y9ZTEw2J+BfaVOiOybTphNaItPAr/QG+sz
zwKugECK74scD9KNOARr3Yf4/UDe4613whyZghYVaGpxv54FoGkrO1cHx6V+
DgJR9OWgfRGTfkS/e6xxI4FIy/YWRc6SnQea4t/hEasln4VtI68aNiB/Nb+E
KWN1veM2vagao//0dw3H6Oaa1Acn7gpu2FXAbxgA6LtYxYZHqdQ+2Tye8AEU
3Fam2o7ie6MFElBwuuurzKSA+brPkuKUaM2K2fQTwJjzHGcHQ2Bm7UeOmuSz
Jgm6CEzX0QJ6YRaIgn89C6c+JSVoTmznfqrweC8ZWlaXoSw2422rMsGjEZIJ
D5mgs1N1Njljw73Tqd1KnYrsnSqy72zISkoWmTiaPuDrj4IfOGmWeCyS5L2j
gVYkdQmUiGhV3ldrbLLB/h48Euxsq4C1tfpaabi6wWr6Jr5wI1E/zFUdmAFY
Wzih7r5gdnr6aqvpNkCtcwthbhkNsW1q0eeSrZT4Cx+hOnXzVIVMTqFWOuG0
8Ijd7bwZIscAwkWcRqSPscHwcSDFxMQyTEKiHzxZNVKXzb/g6Q6RaK3yP+Tz
rwvVxOMVZUMIrAqmJMrMEiMuGgOXdvB+O/8JMMiYyrYgnqqs5F8hHsRvYCFI
DYKfG80BjL0KEPo1Ho7teQbmAm93IlPbsVB3AbJBnf+yDXlc+S+jjlRJND4E
G+XHLBgN1l1wW0anKpSYAp9zqQfuko4fCweOmIFkY2GG32f0RGl68iY8XGUE
2Ha+HjGiIcQNqz+xDJdHJ5Y0KLe28rIDr24w8y5ncMQJ81jjZVQcWCkB0hy/
Z6+3UOuwrO2ncwQR5PfjLnpKXMwMBZ1aBL/54EiSbCPDEDhEa2v3x85jnbIi
jpcilJ741OWFMaZvXfHgyGKAFCNDE2oruFqjskc4dlMeAl7KkYhOeq7wOe76
ZHz4D27jwiOMXtVOi6X/CjyUemX8W5Fu0VBCMbHFHiYPnHo2117g1D5AQWMu
E+qzj9XFeALRkxqlRqDGj6CgEy0WYsoXLXdcXhfNZIq+MuC0ogddrpj1HM4i
wlt8AUwdqcP0qEsBbdcDvzOUVvMp/JnyyEIhRSorWXWV2Aq9VRka83cqgjJP
zEjkJaV9pfIbROqPPSA0u4QUUlJ2opabY0pYYreGu0vT5G2C2pILiY36Zg6R
eqWxmap9Tnh5qvzO+7OLFNulVciKncsbKOcvV23oGfKbwJxGgaul9Lkhmtaq
+ib5qoFis11mSQ9a7bo+KnQPJjjCSKC1nEMkpntaPWjmvNn32jaEJ3qE5qTK
v0ceI5cxTefWF5LjSWHTod4h7HQlnqmmlN0JUqo6ufA0CDvYSDH/cGjqMzk5
GcKiJWI5WwAFo+IMLa2G12Atqv57iVAKKG1ZeFR32v9ZIeYO+GcIocPZ1NGZ
B9Wxo6VmDAoPnGeb74svcKy3Aw/Ek1uPwf9fSiNljOCef+RFAvc8WV7EVBOP
hvhB5P/JmRexViI0lSdasM7JN0xpdj6x04NlTsDIyZfIzExOFy3ZKh5KlqkU
G8Xt/iDOOKDSZ1MmmjMtND3RUzliQNG41CktF2sHnvti0P38kQljD7xxGmkL
RVmOUSfUOhOW/XS9xSIuns7G0NyHpTzt7TTm9zVJ26h9wdwGc9yfBp4+gJjm
6CMGF8F9dsOGjLtNGWfr3l3+a5eEE86LFXTF8Q8OKqjZtHt9jC7GrR5S7is5
VEUHos39zMJNic1+iOTFwqnC2YRuhXCb1bUF4adjabuhJfphDUZH0uZp05wi
ME0Yg3fBZ7mw3tq4qZtY47vAwIeSr40qIQ/jdWNF04s6bCWwT0cRjyF8G11D
9y6bYXzWbBgbFA9Zyj1O9s01tzeExv1FlKcN7MtlFwJFqamZR1LhnoSfwyYJ
4QvBTjGsQe5EAzf4AnAuzsqRGBNgbeiIRnC5VDCkE8Q03LgO9N7hhFG2aGvx
PTig44wwjL9OrjY9v91dMaTZ21D32rHGFq5NtnuuDJ87Pp1g4QMPkdtMLFel
3Z7AkvbmS8+hlGFXrGGrLB8YeSDKqsr8QvWZFm60A/JsMltbeV/3X7JsdygJ
Og6XTeR4WE9M3PZVu0UBDIOE5+0zBFozhJiRbVuUqL0Ote91uLYXn1WsyGlO
vXezfJZEc4dMKTIUxjg2NULXEtujoeUGL9X7KpTtikkPk44pAXPMosvgBUoK
+zIe/+OcIW6XLeCpHo8UghjVj2Fd7x0tt95IKV0l25aB+agDrIYDe5Pbq5x1
JGITzVmPq3xnnkGP+CiRxkcySQumPve9MiYYQS4RUt2do0+IfRKsuPbJka33
j53J4fAlTbACo6DT8uMEeoAuG0kVyW8BB/FENdxrGBhcUcnTjHod7Fy2GBOZ
fT1ZXuQjLnmRNUN/jtidsSuJtc/x3QkwrlE2GeUkB+pgOVHSGFqd7h/+b3f8
Q8AlGMQAJL4oRpe/Hyziy4uO47a3QzlQdDtSCyomKRgE6Nl75hdvgJG66KMk
mh/FgrvtnBikbJOD8g/lWRCBm8uC9ijcv9k/j2s3MAh4bDOwJXkohmwP5E4b
PyYq9LWlR0WzP1IhNT5gfCP9PABdw7nmSWMyUrRf2+no5Wg6UkQc7vy0SVRn
6eJK2F/tt7WlFqlDqyUmv0RkzwXIvXLAAmEtAn54LOpFlbB6H6jXKTg7BgUC
E0bWQHSSVN8OBSCNu6pC2kX5NPSuoWkERypQ6GSrgiTZzNHLMmjFukcNYp9q
E86Trh1ntFdTa31c5y06NACr0oO9fY/Vaujhlqp2ER5Qqg071sWO1IEn6VB0
ZJJolxQ3Q+ecR0FRR1Q4cwjGN3Wkc5nG4QOyV0NAhbxA9jdaW341vI5yXY47
4oXIvYE/rKI7irNhsjv9gnGkewcm4sEG/eyRYW6h4Jz3qHNkMty2udCR3n7l
X4o3gizgETzzBNJtjEndSGwciog2fPv5P8XvUjsEe0AC+tgfT0rA7jQ9hxgB
ugJOiVY5jzuGqIbsZDyBxDuFn3raY8NqwJ6qaZsUUCNGHZjsEJnJaG7NvMmR
b7WctN/Jb1NitmtEYotJoOJsMIuh+0Yxp6ym8pJheDQ8jZKeU/NzwyrYnoY3
Hm1P/x+R7ploNmqMXNs4wK5+ogRmSxHBP0nukdAjTTf4Euu8I7QeYj+XXw0+
7SCLMzUiOJerImlBC1FVJVcDwoMqlXJD4tGlEvL2OElJy74YYexLt8kuvPI0
2YJ6mNROuUjL5A98GBLdq8vYH/cfbV9W8Df0FXjeiUrJAGSuS22BBQVLHgkT
ZvzKbbCA5yk/tpJ6muicwCB4DKFXmcYAcZXEG2FK2NbN8x6566xDoHopOtnF
uY8TRX4Fdv8pz0xXj97cUbGboZSCjTX+UEFeW/fS3ZejiL/JJOd9XF00j1t9
scoGcXO6S9Vbd8KA0gDEGXVnpXSV8Mm/rSfbruRYgrLnQ5FbfJU1PyZ5d1GI
S2iMvvslJFzheWBK9d7Z6dadCO1Nip2qCuQf9SkT6e+R6Q7sX77x5VYozUoy
xDfZ4r3w9HdJM8lh8itQIxTU3JomTyBCEaGwSk/LlhD3NUpAtGsiOWGvxv3u
mJ3VaNbZ+Iim0IZYfN4zOAA6ONIrW2bbvFH9oY1QGeNNAyAyekcTwqqRpcZ3
w8aK27Gltga6PkTTepDMpq9Jy0Hbg54MTd7Ej9unu6lXjPDiBFDjaT9suhFG
EEjX+5Jb8Yg7sFRr0aDlhGZUv9+f5cGqYyDHo9fbTkXngEpMCTyIjlCxYi0h
FSBVlrMXF5HzZSXAhI2zbEXpXwYH8sEBJqnio5vDeZGhUCxqrQX+FoEsc5mD
PlbOyz6SXx9Ot9IZJJB5VqvWnwIWg2WBLROv9OehDqFcTlX8l8Khhlql/iY+
zdJf1uERrfiQizQrxiqNj12dZpdvHNfXyCLYf0a3OLfe6FPmKAkcPSvarVho
L3kmK3YLeNsO5ZZKAoc7LcR+8r6mJzafzt6mtpX6Ldj342Xr1oN9q+B6HXfo
uqXnl+B2L1Bg30o8gaFd1nwGrDCUyrCJjVlMbKwiz+bR7wGy/8NAXng6rVP0
/XfeeRvIwxSmHwh9jRQBtqBI4Di63K/AchjLdRKLqgvlp0bdcfnve+iFBjxB
XzBOXpAxT/Fuj9GkELGznmUNVx7ox406snQwUqK0XxqUVcHfxZSNmBTtmVyc
H0Cyp73ib7Hkx/lmoXYNTavZ3oCJ/APti/2m6fCGC2BRrm2lP16WwEXyVtrC
0LwTVDsCCF1Kteg+169XlTZDEmQIwGNmaks70k4Lf1mg0qsN50f7Ur7LSxT8
P1Z+vWCnwCPeOYapuUod6Vi8M/zfZM/2oAIZsVBFguheu1h9V8OBExU47a17
jikLyhSO01wc0BVngJdZznkcokxMt+BDRRJ9/A40BlCHBI8zKGW5J5gzhKXQ
RB0B21mRrRVja5kr+MzVJ42yr4NvqDvxCF/UbFG523zVCPHkPLYfFCwfIq3d
WG4nhh8z6ESAurt+qo1K8tV0qzf4fw6o6mcpaK+uPF17jiQKpshwAnu5CV4a
6s5mgjF2LfrCyp38L8Bn2uvrQ7DvrXFV+gZc+c28BI1wv/wLrECzE7fif7SK
LHofXdmZvuw8kGrjlwccDaTC7VWlh7E1N6alvhXJm4C5Ib7+0otLXY6HD/yJ
eQr5+SY4SzNQ1/2pCyIioEEHjecvfVr25ibY/o2k073zvJgP63PAZF5ymuYa
GGaAoPjfnHzlWMuau6DeoeH9kUchKHJobYPaRAwawITXL4Y8reTnlVSqwPIj
64nzyhbcSTkUjO7Y4fVNPgcDEw91cueiL7jw2qWyjZjTVyX7Uy+Rn8AXUwIz
yvHf5WMZO4xpneLuIMMnkzi0GKB9GTEgmK6EFFw2WcEC16LiE+1Z0/BJcGeg
xgzzknvqQj4xiDQgE69yvbRy5eGrxQktM5vhzBzXW3JaEAGchq4VZTpTAvSO
m80UWaNFuP/Gb4Us70660r487sKpYevpaw54wO2imx2PR7LEjgr5/XjDnthO
EN0K5oJd6F8pmt+iezjzLkkhMl6+/VAwmrigwSK09Y47uqLGWoYrSL3Pg10P
ffjd86poAbz2z4+79oX0vMojSwQL5DwK8W8L+3o3dVPbQHGWsbVkb5PmJAHe
frK8Rho/5cNB/3LHGVSg8bQK5dLEMU1KnTJE0FKVupo549ZNiuViwC0rjcp0
tEM6r/1jCOCwkj6oLF9LYPWlJPkA8dvoD/bAPTqDWO20yE4bCCFihKqhWvtS
7ma9sNfy/Q04zVpNnaYx+Csa9NGGNm1GCFFvKDR4ejBSYh4wwqsUFEzkm4zY
l1X4QGKdszfq/XHp64ISOFshkdGFyCk72O+xxlqLaUy035Bztf7cdwyBMGcS
I52MNxSz6hI6CKA51HoluJyONeu4YAsYcQTgh6vVwTP4v7PgZwjNvm9BbWN+
tb9ul9OkFRnNoVdVMtcByWFn5iTUaHsT+wVrdhNYZ28AivyXBLQxdW7JlT9i
MjLCEmmKttbLX7Pt3E0XurGlSXwlXsx4dxkdO1+C91t1WZBPZa0qXzcLCwiN
RmFWo80kgGptr++zvBULVZVaRKWCiNfzRoi9eYgFbVj0vvLG+haKSTbOg3rb
KwiW9qO+zp8ZHqN9m5TAEIk+oB2X98bf9ERUFAy3IXy9McNTzuhx2Fu9/7nI
NEWB0ZMALCiVNnCse9o4X73V3qQ6WcivnuET6OAk2p3z80+f9KYU7eQfZDQm
YYmuBD5bIfYoKoAklnL+KoswbRPMvLGB6Bsd0GY9eudCJwTAVIgmYKwl4b2A
1UpNJcW/lcHW7+M6tTxGtAYlyKGd47/186ykz3C5gv1cAY+oGdMN3hhp02ib
xe7oDeHuHjH+WWdmOKkJyM8fFFGq8LpK5MAUmsuPck7WMxcAn1YEjhGL1ikF
X6KyBuhHzbmeNMnmM0nFdXWmFrCESKXrIPCDjzb9CQyDiTEBGWGgjtr0D/T0
sD5LbUzBAcdqiP2S/KZnI/AEtBTiPJeTXd5nV5pyG3py0zMw4FhCW1ZoSDPe
jQAUT2sCNynNhCIT7+MkNBjixpvyUpq/pTwR4DFX6n8PKvTRKpdJuHyYV5NK
ZHI7LjrLsxtgymloaJ0ZEu2DJ7Q0+Sp5Ay4AlDFIYpWJ+FhF6ceg2oTQSmtc
J1ehN76QLS/kmbyQ5bfj9YfoXAE9FbqP0Wm64xWoM0PGkVWEIyRY4alV/cDV
3I79cATYhjgVx/W/VL6cNnJHiXNq1qYmscbBJp3hYT4YyEbnadouvPCwo7Oz
sjQVUrB/vSCkRBOIkuYV8+1LTv8S3Ba6pkJP/3u/JxdU7S98tJhzGfb97Oky
577EIs0NQsL/gtHdciAR/CsF7wpjgopuvfGuBZRtARygX3jBUUuuKnM08dHW
xPMXH1/kqBj5d7It4efGpTNg71uftmlfPnYXz6HFf4TNTtWBU9cn8HbJeTF8
6xrAsps0qEO+aNQKRd1m8vmASXzsHLiAkBwxPdVEqXhyfZ7GVkRNTksuUgDY
w89tj0DCmUC/WnaqF1RdbKXsKsXnV5ShIhwNObiv2blv4VQIjNEsCavF6OTc
e9BOBn/0w2tWCtqitqUi/rZvrAnP4FZgc5BTGAYsCh9r+1xzgOvF5rJqpgbk
OY8xw0Wqf0xQ5MDVNsZSj3hWsBobdg0GS2Q8aRK9KEkpE6RG08rU+/xMotmu
ZoYkzjM27PxxyqGrxtMl87LDfgvqalUg2mCniOjpPLQtG5BSSdgxVDBFGQgW
03JTdMxnRcNaGHOm243ttGo+EXDySGm+cd3nROhE4ujeh6r5zUXTG5Jru4NK
0gdLYusyHfjejTMX3HRvMWugYS5rcnTetNmhM+We7QBh7uTwIR+d1VwxuO5l
9fh81/76eDw4DAito5KVQIMJwYDfUFC/VTB34UFeQYh/f26+n1aDZ/HKDYpe
OizsQqRs7dodUExw1FhWqV/5GgPlUb6RL2UPSao/Dho6ovDhxvhy6w6UyqL0
O5T3jx7qekGhpYcYxepRW3B9COOneYhS50VphxjADvZrbk4uR88P7oU5eKp4
oUka6G6EIKr6cU40Qummf+WynLQeLpTE+Mtfl6zb35y+PIiqIpRK6Bu4yM9k
cdYAF3Y3utswEuSeK12p8rZtZBQavMrzJDElJx2Y+BPUA7uBjRnNjkrdvzrH
W51ChRoymdp8HJum9J8l2pBiyNmC5B6Md6xtaziprVoynLBuhNvivtoW/fWM
MMtou2p0yN7Qdg1npkXua5wjPJy2lHTgNbmXmT74GuXSV4pOd/NqoTzVmlM0
CntYU2R6qJomD8droWP8t4IGsVC3G8+E1m0QXlJHQHtnfXX0QPzlpUW1pcGh
RAsGHJ6eg3zyM59te382OwquUHuN73e7QCpbCdPKYTBcThAfIY5LmeV2MjCg
5OnLeOrHMr+TIJv25MnSXNzhyk9gDaMVew2KCh+p5aO0x7eZoT7J+7RV0sGR
SQ+XXLAC43r0ch/v75eEsh3prcBj67GYJEddvs4FXraXGLbm26w58PVFt/Dd
YltsJpGZ6XSiCHSm+ASkKb+Qtw00IyR8ihu4zC2HKUo4Spya2l+87jjyMQ8s
+ygZBu6USRnl2veuTYqD0iAT0R+g8ZZsps93qjVIA7TWZZANSgHjZhpX6ePJ
EM/n59lSulrym+Rq0ew1T68eo7KY8WDmKO1AZ2bSkBdOxqZs2F/IOD74aThL
4lsrGfRu5D5lFCBiLODOZ9BW2I1HSK0P9uF9Fs/nJ2ZRz9BFTqtxQAY8RuHh
kVoInRCW6WLwta9/WUP/9y7ZQmsWYnukGJlspv1yG1i149XBvJVsSl41UAl0
S4o6MmsPfzH6YPCgr+JOpuQM7TWSJvlvzJ+0TZdSfbm0LI3K4KEcz5HRnD2d
R4OCQCM4zehbght/l8aSiqFfD6POyuTaHjHbOhPEQyxgOfyLVRA6RrhVxRaL
mEW39O2ufaAhr+JVSr2LFF5FvHVcjJJ51ggH7VQoIfk7i8ari/s73dT9AO+D
c2UlkN5pHTxgwuH6pPDUDGXG/ap6iXgJ112oGgI4wjrqbiT/zXe0gpPXHQFs
KPtJLsp9XBg4GKF1tJLdqC0Ye9s5nSZcbJYJ/YJ/2S4s84fzbNLNMxmFEN4X
sFBuKyOt1EOTVWzHgk11GlxLzosi4XZk0pzQ5vcUbjF9fzAqFCHkQ0vBoVVc
UByRuIQMLxu2K1TavsFwBCi14PTfncdGlu0JE5jTLbPhcu3wyZfqPwx2g+9D
dkHSvf0xqT4hF9BHQq247wqrFTBw7xCjjRnZNL339EtqwzepZ1Fa+8I+DLwn
GFmSi4Kifh/26OnWI1GArcMsXkaxUejrol+OzBNzmv6QK3admkJf8NNUIl45
2izoy9LJBZorgH1g07+dlnZcsoP+VUgCT5nv4c2EgbW/9aHdgbQvoYP2i2ch
CUwVy5x873EI62LLaRkM94GJRJ1GXCBOEjYGz587SS82BCxs7s4V32mHoB6I
UzeE4sy0YHBrria8Y2llq6c4P7ktzicblHWyj8o6HMxtAiRUhJC9FWZd8yms
CLQGslIjcbAVw9zwCof8pOrb/K+2eVTqAOI9NwFEcOFOILzWDFHX5koW+FTY
d87GVk1QdRvamjbcXl5nP8PuXwPj5RWcPkouMYxC2DoCOahyBVS6NvD36YEr
dE9HZRgSvQz6rHY99CD0Qf3b11aV1gOaF5LLKQPA32m5jWgF/d8IPGbspTlo
o8bEfYbNh0lN3iKPLxx1uo2i1gMCOqAeTuu8zqXTZIAOCG+zhR1zR2zBYU8C
zQTnDfDMQnvM+O1DMcHunNkQHS/LyA56lT2H27GgsFKVN55GYEv2GkNSif1O
Y8YA8RXkPBnwss+xNZy0s8m/oeiXw36If4QwQ8kNTyzc5Gxkd2mRC5Ew9cnN
/nNynbTpHPBctWEBcspSyNc5vpAZNH/p4AifqCH4n0rC7nbVpigK30bTLm1M
sh+r1+ybYIhML4ETyiOwJYyWF0dUk0IBvyJxZCZEb9nKBDIkD3M1AAaQHkbZ
4h//lyL/yL27xaCMhJ7zbNII5GAL+Ka+bevUJFOhQ+ObhkqvyIRtJwg9JNtg
SpQ0MDLC4EhUMhqSxSY+yCgRxqFVBmNh9yt8/iwj/zf7ROqQj8AecICE3Ldn
qF5ajRd16fmPqhGTIRaI0sBBYWhCigr/UrihSwH7/NUsRa/UY/afpYBgZC3O
ok8McC9kcq9WHIQ4VpECfzNPk2mSJB+BXeM2AlwsycrtQ/d8Ywdht0UbJulS
63VkIV3JURnK+NXwbtMUv1bb/AOyGLArks6XWIAzIW/5uk2xYb7GIX/X8Z4L
5J4Lz/2wT+irWlkAn85xEZ8VZk4xyYlyChD5rW0luCty2Xwm9myKSdcLB0hr
5L/yKIaDcrOmOoQsp7ucblSuMQWIzWREf5mDH/O5lF1w8YHteXtAW6C4hnY2
DBrAsQjH+YQLJQ8nKhv1swux7iHwZvpwlungePX+kDnLmp9kKyEPhs+yOGry
XPodEJvUKwGaLrfX5G3Bfnn2bzWpjTixVY9CnRf7Am9cocTfA5jWNYdmisCE
JyZdS4Yw+2EaaD+bA5V5fVIiYDMEz0MI2HeT1zIli5WyB+TEJZAVgodPK1DU
fKttDxXNejRwuW8TBX4nmToL/x82rlxzBtvI6oKdOUmHWbwPyVfqrnuifHIY
kBgDOMuZkXt50X/sfUeIeschscLVBqIcAsNdUP2yXXBMNb6jhA0159mlTr8Q
JS2pPoMoGUCQFe+gdc6LA8Dic54RYQT7gmm0BFf11p+zp95F+enoNkPeyE4c
zf0N/YqltumaH9h+f1dy2D+nl4cKJgSmVvGaB2aTY1H6qvA+GvSnBFPJsi1D
mVTe+iKiZGr3Xo0ejh8t5NsDij9cWk98YewpYqnyFaGFUWbMlWVpaV7IMxzD
39vCEiif4aMw5UtuR71UeIykKVmp+WBDKh9ARZYHkWGN1U/cf8FBISDLZtpO
khkHE2md2iwlErfRzFHAeg3EIUj+U02zB/gz7FIWgsZzHVj4q4yl5PWtsMvc
ma7rQrI+aaDfn5B9+WjkaP08zEe2tR1oPuVJJmbiF9ga8iVofG9FPFSMFweI
QGsIrM9HyQez/xVdhEWBxwEofq4HWaFXFizf0p1cFbMEB96q3iqk7TWPBf+h
qmm+DXazw/cs0n5DQWZ/X4VQsp8qknXIT1VBkWELmme6TWS3DJFP+Sbprs7U
Fy+J9l9D0SO2RBTDrNRT56DnI2GrRcLsTyVbPfY/hXIJrzAZC3WzCvsk7Mw0
rgGDg1HjxvUeNIBrht8ayMfx0Gpn8OjaoAtMcz3PVAeo20diEs6rJy8RYsRL
Pr7uJnfDjVhwYm+fa/0Bd1SnROTwIfNYFLHcL1msMhgtFr2b45mWTRMkzsiy
ocDSttUv64EdRyEqpOEq0IDgB0fzfXN+kJ+WlaBZ108xG59BeBiGAWmcep63
llpXJEC4GjTdWKImG/BcR6WnRzs+8OyoSG46dXR/BCRAXu4Q+pFBtImTDecc
vbHWNpzwu8UgOkeMCElyCuPsTKaxbfqQfpPbHEbntQXo9gPZv6pUpUHqnLwH
nMBjMZ4PxUDY1L5Toua3Kuu4I7xpkwzuQ/NjLZQY2OnAn7UcoZ5xotDM+Mu8
dzwTINSpztseUYs/1z/WKY162Q8qasBLBnE9cInhj6oRh/lz+6Qvy7MeATYG
EXRmnu5knpcakelpjC+L+10n1KIxuaeLu5xVh07yxYsn9XEp4rVf0e9gVR1e
+z9wE3Xwj1uCVt6pcgpixO3suamCQjyIxBaoBe59RdTbLnvPbzhBsB59Di3w
accHrEA+ZYOPvNC++uxlMdfFTmuqv1pQct9uoo1IsNxL9IQsDs1hMrvxF0tF
Xm40L/Y86XqSBSwXhTxVKR7tMwue4obSP2cna91K3j7P3HVLxx+ME4YK73oS
lEO3DRsoadPrK+SLum66NJc+RQruY9OS0z9RUqfuNh10p2fcGj/OzKWH3uaP
MN6zhsa07uIFDN6A/01wt3uttT/luKWcOrfd6MGAXODqtMfu7XLt8XVkhksw
vSCNbM2Em6cOQMOueuFCxa3XejNhGm/1ExfaMiwUrSHeTjiQ2vOw2Z8XkI1p
i3VRvHBUSlRiXsyP1BDNtcBGRwVY7SyquREXfCOwXjkAlEn3egozLxsA1dv7
Bam+MqHjqHFpPPRle31qbF80PQ6oc00EuqegQkhuQFRosUmCBoQaFCIoKxBj
6bmZ0HNbAWswbb1RPrzfNxoVXcn2njxZgWEKZekx4VDONl2POUt8DLW+tXrc
AkJZe4CHE0ZzSV8JJfXioaYZ5bjqmK33arNOzt4J9VuuoThgrTavdHGjJuHI
d02aLybLPvacvDFFJ7UwigvNpmtzbyKZMcYDA1wg7KP3vaZSWsfEOQD+zQPo
zJdKlkY0ip3dj3TEp5ZqTxijc5ERgFRUrwzIrspjTw0WxTTmrD+A/Wq/av7p
NJVSRmlukdPVaHi5Y4bGW0fprpc/hZSeOkMf6pny3YJ/cPK9RomuQO6bBNp7
puge2utsa3YZU741VeiitNbMxnX3CDWoO3OVhJupV52TPA0F/AMgTADzKP8J
miJvj3GOp5gGOQiw2oaQoL0COKIlaZmMxa5//5D7HA+ucb8eErNv8baCy96Z
WgzHTdW2EWALijLJSqKRfBrN+JqRlE1G/IfyldDLTwFvGvzY5PYLy1aOfGXI
E6EeQQ4AihssGEh9BSYgK9TqD0LxGtqoI8iorfTIwwjKvt68tzLDUACBu2Zl
mjDSOZm7fp5nn2iMR8AvmDlA1IuxiZ+q2Cn/Ll74/0tAs2k8QUfnW034VssH
ZSG3g8/2kHxXDC7638rr3RlPKxImggUbTpac0YcoUw8zHTPIajlg0jfRWLdo
lI2HBgEWJKgVLWDP7wJUoTuYvRyAk9qNQA8O+09ubSgbd4apezFAlQo/hyH9
j0n0GJyQDCMUK16D9SEUWvomslLUE1MIcNxhTZth7Y/XsARTZQFMVtgb854m
0ApLokCyehLJHg27jxFJVb5sue5VmsjNi+BgDMmiPdx7uMKOzO8ThUm7NswG
a3K4moL+V9lnvZa3F8PUGhFgCdgpn7s/0ib27BGWPdt6DMuxptoe3/s9sX+m
UdTNEe/TqR1gQb/ZpVREKpPUUSTBTKl9/sJA08IT3eb56F6FKIOr7N7Car1k
jDTatnQeLyhfElrVRZ508c3wtxlInc72vjgNDIxM/yfDqwY6d/CA1VGWs5eW
GFKKfLvgy5S9/pXZ2/+ontEmHJ9VpaPvg/fp9ToFlISEWhKuFa6AdUgLtduL
YtJ4AaypDTbjL9spV8FVkmKRgFwpAn/gTzbsyvXj4CfrQNaOS3jR3Gop5aTr
YSeK0MbgEElKSo5eOGCzOTbI/7ln5UnuaOGuaFrzMx9AVEPxdPH7EvmX/hpe
umGqvAdkRhAq68dZo2kXZSEt2fTKUrj56QMUuVTaOWlhhbSPdvOmwuu1/Rsm
3q+P3eP414rOwX93ND2o23Fjz5fDT69jS5R7rFyZGYtM/var9Dmk7rrjgwIS
HWVfQOBpszm2oS0/+NdRlbGwTIkYbHvGjPnag8JbI22hAMObzh17kGwzKvRo
RXfZWzJVUd/S+mZ5wrgBB/GbbplB+8pXOTn2lm5SDK/+Pun/0ofeyotBXJ6K
Ej9EONBzocd498/UHreiRZHKFBWXhd3aWKQUtfPF9/e0ysLRAt0wCOxjQ1fM
Ppq+6nu6BfRkzKSk3p85+6vG7wvIh/booRv5FNfguGQqF6qorro4siCzliws
ccQw+yNU2o6gwShBOWtgzwYKOfAmmcQZbJ9aIUqOYj0x5ypixXTgRDhCy8go
LSvpLwZVyJ/EVrujIN6yoGXN9scWoRZV5JuQdChYaSS+X1NwKHhTvjP1h+ZX
RJ4Jzy7TnTNygSfFEvdNKV7L/xh89zv+cdwhLMTiMHgNJfPTlYQ22JmVZVbA
cWqHDpQs13TVKt6kvN8NgYauS2qoEeV0OH6cxkRHWPMif6Li/Ee0iEy2IDPW
ZccB/lL8oAhMK9qivTRyxC0lTM2zVlQiVru152WP2PLYlQgpNB87p7lOT7Uq
pthJLlFe3nUJ6dpAM1RF92yRCICi8DRlNkXfXsFu1x3Q4sDwPFbTcwEOLehl
349ikQ1y2Obc94uXCjVu8TYhbY4JJ9I6WLSdwh5aFN9wzuooEqmmRH/17Rkz
gDs++cye29OQd0VI1AvWJ3xj/6XxlxiTaug+4+XCB9xTE3NTQe3c+6Q6C3lJ
USY40ZPV3w+SBmW1cAZIiMkZtd8DNAB2lSXhlxJN5uYua7eA7t/AtxF+GSuf
Fw0MSZ0sTSWTdwuH14D1D0mUgWdxQDkml37MwAoJJK0w66+qvEetFBmWQe/t
d5RBDxJ/uilLhgIjD9jo6dBMwqWwinu8yI4l02fK+wizrC6umzFsNWJiUYKM
L947/FLd34HxbqZuS/D7ZmIFQG+Ap4Nwp2NmNGw6uyQIvx1kYe8sIgBtEqS9
DKGz76p48pgPK8RokNVqRsL9uDf3gy97Ld+wJaAcY0usuKO4RRO9pESfwj9X
H2uf5Reqo9H+02rFWbAOqBrEvr3TNHYzJWY7dMtJ8MNN6oMtKVpZZ40TH/9+
24rJXn03T/ImW9D0XMOYJ3qpmREWFa7CTMlac2lb38ZoKz1QCFHlGAY0wiO5
FSLHvoAcXIbuXI+k+GTJWnnai2ZlnTZMemnQ1c1du830cNK7tNdPfN65UMqa
ZrHfEtOb4YYBaTs3c4rlD0yzyvAvoQrRjSqjlVbXJHw5ju5N2Zo0TkZWeh/h
sjR1yhYZ8gAkI73XBahZ2OgEKXlAlow60L+cNYGwGMizE3I+lzfe35Gi9GwG
kpgltcEKhiOh5CYhBNANVAzSxkDNShaUZdH3ql8M5IIr063ZO4za+n+B/Dgf
wTL2jhrTJw8/ATqxU6I6I9w9fR2sQBVYyO4iyGCZCpWQ3AFTbmGs9pWgrMha
qJg8NFaWytn9c1d1+EgZNEtpYgMX+TN59kFXUQnu3UM71ghwRIUWjJCwB8jg
OLgPXDKOJrdfFQeWgd+SY3H+29n4JQP8JNeKh7syB60KasGshBdU4zdkCNjr
CQhdXyQDKwK95VNT86kTfAAi29aLblHS2LC2g8EsnksVhe44y0ZOg+EP3oXx
wVCvZtIELSl+mbPe72eT7vTDlBpm4GGv0uUtbHNdSYaOAyYaoo3k0l1QF4y9
p5MOKeiNG6yQJkGtqnJ5w3vYp1g043ahB9sgf6nV7rLT/R+SRB8Z6hNFJNgP
6By1ZtFGEzd4AP1y75jiV+bmg02t8hiKd0Wv+wXCnosnaWCWtWa4FTXFq2a3
z91kBR+atns62a1/fFpkiLxew1GH9hulwwL7pcMhZBiLkYJnNa6f5a2swNXn
l7otwgt7WoNhZ8bdIsNVNHY5h10IsNXpElAF7jx+uy1s4DKGxa+GxzbSNF8B
xk/VhMC1BGouL9rvOsTJn77OeOoqct4+ZcF9p1YN8e5VWW7CDYnFr2pnDXlK
fdfpJsGuViAjgIvITdy10XVLxx8sPCiCwe5luySAOoGtx+buNTjSedx3mrWA
rDSRzRYVn17rFTU6itBGQZnE+Y6rui720YxLrV95WxEE8tuzHeWcvET2Reur
IdD8/CJvc+duK36KcHERovQp2rXjcLgxPfrVIGIuCfm9wZGKlhUqRgJlYddR
s8w+sZej/nmd/i89tgm+HZuEc7AklJQuCZla1mNd23baxhBP7/kq/dax3Cmc
hvKwSJbIkQ29PpdxQTLW4IDZs7cgKPsoll7KUVYXkOC2AW/GFJ8CdfjkbYdk
zLjWGub3zUwVEPhls7NF07dCfXWzNTTfpMoAMb3DUfq5tyMH78eUV0YvkJJz
tzbmZPIlva89d7jCT78wGfJlrKu3SbV09l1F3fiK1haRK1BsQp+RiSW/QIte
CZu898Eq9QC+3X8OJw57nqVm8VCB4oCTKH6kbIQSXLp1zIK/K0WossESu8Xe
K+DUCTsbUvbxyVdj0EGeF/5bKInpf7ga30cNMhsdvm8uLzMfTEd+azqqWOZJ
qXdA1JwJaVAfUponWSNVhqXgJ8cliKyD2ZAj78aKa19HgRJkMcCBgE7GffqV
FsvtPFIy6RNnitSZ6mURMikRce5R7p6vhWVBsmmtvl6tnnaG6rrdKTNb/oVp
O5B0chw1zJ6kHTLJpgHzM81ncNohNqZvsSrIm/ng6/It35nqD309g+uKJV4f
vsqE3C8SwIdNlBlqUYxNwdLcGlF3ADb9Poy29zhVMdOddTTSA3KgeiW6WvCJ
gkVhG0LBs3ZpHnx0Vz7eYDsCvENQWtjjoGmc7Oa5mNunxM4c+w/xJNzdlNFL
d9Zi/odwsTS52oVbF6KjMSc0jTR6rnIA2zTPo3Cwxnqzdp91eqjn9G0fKqSZ
ihl50U6bWsreGVFZWUZ5sosZvSpdSq8kXb7SHQ5JkzYQeEQdOWJVgJ2lQ2Ig
/H1+oBL2lacbfm7C/OrNVU1oobRr46eGZdO4j3sTkihjEu2qxDG+D0XvaiA2
NNy4D/ZP8a4JNviqQs8x5bujfKca0PPnJoJTL9sVpvJc6qfwlB7iX4y+XIdK
x1ZWL8W5j1M6w2fGWqa65ckCB+eQeAxGAS1SyLgXK/3vYfTpoQeQR4rvE087
qluDinFVmBLjjm7bw56RqJgBFnNcZHqW+t6cxz/jFp7FVS29UQPsnATxguLB
Efb0byzzMDYoxog4HSAkHrk/+9JEF8Nv3QoA7bDf2jaRoICTidDuXKH1iLf4
Y8Ru+6VQ3pRr+JtUuiXVB+ZOLattgmK2UbLSxGtT0d8hTay+M8Gza3qxlV84
AzMHwjysJKCc04rJ3eAQtk6APtMMrXTqDUVmFtfhjk/DMxPPzjW9wx1+49BH
77Tdanx3TCC/RyxgMsBM0kH9PACQUWRtPV9v52CDMMdNtUfJn2qGWKZoQdXv
wELKswGbXlYCSOsFp4lQIQasEe5GyDdwaiFZ5NFGsQdwo4glwBUoxSVQuTBo
ac51Ndh1lmgr4LCszkNlZXpWqUmULluWc6PUzQ6vHWWoLrfc8j0sgUtiW4SY
TAarxLSTWROfpkdVGo9OgQLHpkzr7Ixxq3Z00apGzLlBLoYbbvc4FU25aanp
eKbRkGBjKf8Rqvuil3M4MaovfLD6c7fvFItwYSwuuDcPvgjnWfTuUxlg+K4O
UDrF8wQxSuiX0+XDdCnc2+8aSu7h3fUtblhVpYnL3+dmm8D7Ww4qakw1gVmW
D7wa3tCivA2/QPZazPGyYNv+hTUj8shn1Uv9Gc5Yb+umdROAD90UBgJ2M//9
tC7M9YJHjC1on8yBDHXtRh0CMWOAU7P3CSHL94+jgVYQacX352LyAihvjnYc
tlMVvGxR1FrXOhVPyf6f1wTyiXFY2byyvUFkHThvNbaUhvJUI9NVchZbN6bz
HxvpY30kPWadYDvgNCxSnxNC+TPo33yHwDHs8HJUwGiMieXNCGBz7LXJH7hd
q/WLRY2Fs75hRtkwgv67pY2KNSu5TwWU6lZXMOoOscI5y1Ph3PCBQWPmgm2/
JQSQY32EcAX2UjRW7pii9c5ra5gouDo/cYDYDroMCZ5jKcVPpqipEnh34rUq
K4F4UIi6COfnv2Cot+77Ckv7JeBAiWEBJxL0XBdJGcO4Rxc5JeKSA1baYPO9
2mQfw7WDyCoKuDCuxZZEdG8TzSfIUJq/sBH85zkkm8yyiOBTquUtOF1W8TVI
VfM2n7UKVty7fPassFsgGjgel4pGr0FfusLh4Jc0X40+uv+twORDXlq0S2YW
DKyv0KzBiOfGET73vkMuEEcOAzj9fw1a2xJ1N2szm9NTWv43ji5OL/PnSz+8
8Zw5jFyv5Ye84Ldq0Yy4jKw6yNFglauLX1c3aU6XOQWlSr85EqRM9sxQ2SYH
kQoD/tMIJKsk5iKErjOx1LdCZxbxgf0WjpY2SA/M41tjTl2hhHLLdZD6k/UF
1I3jHtDM9oE/VjLqb6qvPYUIdh3F11MVqjcjf6itbs32HJPviCET4gXlpLXg
aa+sqFqmXAfN18WpOiHZtSz39rgsT2eUqG0cN1yzMrC+UEsTLX8yjnQmVhaT
FPzDwdZFw9lQyg40Ot614vk0RlTPIpYdS2SQreFwTHmcHGBHPzxzLKLmBkI/
VRQ8KqEo4rv5Xul+9W7NONbvWyrIAFLuEdwM2Fpo+5lAMqJZj5glIzghrA8u
kxIQa0gRoanP38RDraOYIjsbgD6bnq2OIQXt8Mz3gv1/t1AkWWL5VXUgw0vW
64ZcF52rod+f36Pb29ngHlwuWo+x4YtTmSVMLwhPSNLcwHLw+hgre3mAZsxG
55tk9TiSLLHJ+VzAdh5Sl19VjLgh2sTvd84WKaD94QjMA7Aod5f/gCMQeeJL
kLJRbd/AKhhrWVooqZrQTai5Qo68VAyuvQkQAbcatSZE7eRp8QiSr/EO4xNB
L8n7qkDxOBoOQyP4iH9nslCQ3lu8lBdPAhJvYApK1gVK2LWNzxBUa9bnQ9Hj
GaYo2ZBglikTsw7tP4O3hAkL+oKrKiTyvFP6ZfugFQyOrexSw+XzH3gJRMK2
bUu5zcUk/rX8lZgzenpdQ9A2yOiw47CHSY6y3jLXlEXPga2eIp+ldfMchqpR
l/jdgxWyWU5TaVc2+HaoVBNxjm/o05fpNbhqOZ3AoiVf9T1k99+g58JA/P1f
4QVs9LU3tJ6J+RgUEarBRQP8Vme8BgnygKnAYN4JJ7+ngFVgdSHRsxdd61Hm
lDpK2ve46t0xg1QJhAzDGlex34r12j30l/fftNL0DFllFnEOibN3oilYcnqT
4y5GO5Z7VYmbZ122AgLj2YKW64Bn09ml0vZaU2Fq9fNUl0D/ge6TSpRDN27F
ff5ioglkY3VDh+faUmB08PSx4ZhMcZZBv9pdYGdS7DVzVlwxgYPC7FwoqXwD
a/mXsmvVRUeoowMq1X5R98PmIKFWFlSZ12vEhk6GmHPpkv+c3AoOIxj8IAYg
MfWYYZEDHFyU+PTvM5gStAB+paxf0V8puBPYpvnLJnGzmn2+s29BKPI7xPCw
9HUGbYtLFhT6ycEcba3xv44m3e6ecydgr7scJ8E1tYDU9Wk6+5rxHMjWtWTc
f8RZq26rbhxCb/vBETdDSSXFYQmcT/R8qeYu/W4eKY4J8iPrSOdD4iepXnki
mdKycV8bHQvSeiqsy1Ctee2oJAEhafMPrHrqcT/0IAEFgz9PJQF3czLNq3Dy
3teoFTdenApd1yR1cVHGUgwlRUvp5pkYQ/cWtUKqv8hKg2Fbk/SKqxiPVuyT
Zlm68sD9pGIXLuRpr4r3QvkiCkOMsQzbf5xF8MNfbuhcesG0D5nd2rcIwJV7
IBsj1xSM7ilIFHt3pINfSRhWf1ZzcGqHRlhbJeSktB6rQNYs4zyL9qKjOxYi
ppz4tqZBw0j9whTnd9a/WFDO3AcmpxXL+bPYE25Wcg6m20beQeIqm+KHhbiR
iNjrKZbAB24Kj96qj2dPHhFz8XmVWJP7NBtpnMGSvnlyVMIixBs3mwwp+owM
Wrt7t6dizH0qMvtvOLcCGHvSlTcpjEuQm/r4zYFPdy11QGC7e2HIwwrZAXXU
hpKXsOZM5Bx7v5HdnBoY+FCTJccpapHjQUB36nFQI3XgMbdC4AWJVJLRvOnV
GcA2SI7m7s8ZCnXwc5k0tFhMKkhQNkXcD1UfWvoQnON1vsI751b5UzH3t/hx
hjcNMRsSQmJW6UOaheCsdRzxd+DHGmDcG865Wc7F0Nnk3gMiJ99frS+jEFAa
278emjAzDO3RJWX/VRQQTdkuJ4se8VcUNZkob8Rj8hwGuIJ8g2P2BBfFS7jf
ENgcItcjRMGFaMqro5O4pN0Iz/AD1n+xkBtrlYLA2PSCPHA9u7HTNVhUk7qu
vjAdJqzQo6d9bHrl7azSO0VZMO5qZFB3lZJctLRAyFG010HOZ2jEf1OQGit/
P2+qXFXgXRO7Ey2opNQGrO+xyWwNeWlK6knxCovP7b9AWYZBIyzCtZz+YLOT
LvqDhNDMp06ON5BmOStmwaP8PSq0cDHxgyVmM4/HzsfKWGQvtfn4qA1fLiq2
AyVC2RoqhvXkdotAg4vDXUhWhxQk7b2Zl8yf/uyzEhNz8Fso/plrBcNEXe9N
U6s7jcglXaaS+9Xd7bwKwkpu+EdVe+BwIQk2EP4CFlAsk1TZqLLr6WbaHdz5
uYzShwFcRsFONsdP4N4i/jNa1kGaG18czWoYoeUil1WnPDfqpvBPRmKQGj3b
YM5OyIJuq0jDm5UOgbAZf2gnQLNuSKaiI0Mu5/Aj8Yz2g2H/oiwBGD+UdooC
YfF1TaW0cSq5iG7rNVLGTQHyLqCyzhIqhk83lDvjfLUMw6Ga5cYYTITQQ2Kj
HKLXJiBY3Z+dK1N7IVWr+SOk0tdiq6FPT/42sf0NBETk4YRelq81EdLLhzKM
vnno+s7V9liNghO37iJHnuqdggrs84IyU5SXjLGDkPT+JuL6xjJkHbo+/Vmo
+TD77YOjCaz0jSr6UXHIoxsjhmi3mRqp6A2EIEi127ZjlCbvXvnDjFnAzK7T
ohlMbM8DVlfzKp4FzQoaeSMdZ8fVo7Ydld2nEk8oKC4anb7J5SMCNYaiVAe2
NzzlJXsTNonX22o4Vo1R07+oJ9tTWYI8D8UmAtHiUcpUws2jGwgR+7zcy4JU
4nd16Q+/Zm2bXK6RpJiKwnV3JC8dgXwzGJNXoY9jwLlBsA5sDPS3LZhMi7Aa
mDEBDDVeMBrsSyd4rn3wL0NIdn5pbYwo+HrobrJPWNvRU+lHP5sJeswBmzDD
FQ/xbjiU3YmoeNZcbbPy9nyP+YjLyKFq5Yw1JZfPREf/a1VSnIfBvPFp0L1S
lHLadPSrWqz3gAPtl+TBw4b/nrwStf6MV8ekzUZct4QWMoEtjz0bCs3XJaiD
v76wGVu17FvyM2KnXRL48Le+eY4t+29y7vK7KnOypHWqwoC5Ouek4rjoi7E4
k/bicVr9Y4nijHyj3E3UwOq1/CVm49fOzNlFdLU7CgJGiobbodU8Uif5NcXp
eeLA4L8XoDcIuEAXZrTAXGgmFkk/6b3SQf4+tXnUB8JbmcvaSv+Ks+20G03j
PMp1vV7LHyA675T8AGx8NSpeUj3N8ep8hBgbtXXM/zT+UqVz2Z3Kq8BRV/na
SA3zNR5A++mzBnbYJy5npbW2CujBTouNAx/MHZps6CY11L2ocFrgEYOP/6rD
vuQp2rfontB6ZND57VeiS/jknD1gztS45rxLdGq2/3RX6n9VDC8pLCcsF/S2
BLXLzKIkGLHl7hYLF3i1cWRHdMKNMMfePfCbWLRGWKkh+33KG23Z6g3KHD90
YiiK4/7xSama4IQSnZT5UE2S5V/NvpOwh5wJfb5u4iG23kooExvNcvrnW11i
hvae1aMgB8xx1Cbo6MLVt49gFogQ8225krJzDktoU+0OCV240R3cVnJDdl/9
cQJYB2vJUc/U7eMr+Sate7vUs9sCItNHYY4h0Ym+Eh63jqV6+MfddWr11SZu
j6DnAzpmcP4E5dT+xHj6R568H+ApCotZ+eRY58Wtm4IGj0YbMqfBS1kmMaAl
PjoeA4IX/KAeEMA8QmOXYXRNvUqEhWRMb0m6I+d7jk0GNld2kQNMSZw0QzPZ
yFBidAxMbGMPmhaszj4K3zEzfG52uXF8EjzdWMRFZ7Kr70ojDWm2/ouG3P5X
h9bHR33Syu0TTwjGYAUr4mtAt5TEWYzE/xQ/mspDAoqWNPT2E0MXG+BSEEnE
SD7O1hT7l2s9vEq2M/U6ZSDpvViplOqgjaTLGbKvVq53cMN8vunroRoRfUo8
UaAVyi0xLHbmqGzdCmfQcFBmvlP7BI+q2EMPsezIsO0j93OYNYW/p8msAZ08
ely/fG7K+s+ZjYWFWKA+O8LS5oZp/aLGs5Ygeh9DhxuLQDBZNgfUDvJbKYhz
jDeAx5u4JHMDKEHQ+oS/xiOnl3O2RRfE559f7qt+9SaV7K+240/6U4OPEBDE
P7TKZiCt6hu4XiAWL4ARxImz5Ds4hSC5v85glpJ92hRAyX4Xu7S0zxgn7xEs
iXMUh/Al8GWpSLyOxToZnB7e+8NKGOLzIbiDYZ0Gz6vqCkdb4BFLCE40+Cee
GvOwsWFFfkLYrUiWNiBA045b1zgcckAW56djkH7mhkY+qfaJHnBYzFBF4AbN
EemvA6jis+sdkT3piDTRKEvjib/+BjnlcIb4P0/TGbd2mkJwJ9ce7Sd+qprW
5qqD88wNvvOZjRgdJCP8cHzpDcXohhSudUI+EmafUBUngUllOP5L87EUoXgy
v7J+pMdE04TWF00u2r16ngTrRR8qavSPiPI1uQGzDPO+uVG7XifezDbSi8Vl
cpWTZNYMjxz8O9+CwIa8YWaTGT/Wg5XWhebU4kmrNhMPpcO/evL0s+ZqXrn5
HeB6yeN6tMBA/DeRrtbtuvQrX4d58yKXr+Sw/pZag6ZiVqg6S+ZSDlb0XWCj
HwdtsD5UctGB0vCS1V9bygUUnEtLa7JwAxQU/BUlyXEmNV+KiRAC6eAtsZNZ
YF/uasL3YVW99AjlQEDUdAmNXZptjduP8yWPxgz8vTMkDJnqjU6xy2TgLvJl
TG2csycJxJFip/EhSh0siE2aNE4XHTvtWV+lAuIzEFhZP5K8Uyq3rlefqljE
nAs5I/+JBH9lBToyh4rpWYYK0FDkLgYI6jf6BAcKFmV5fDoFJlM7dD4b3hm5
JtcRj3A/i10xfTuEIGbnbg4LUkVFUVG0XQe94Nt/Jqhk5gW2OKiOs8fI6Rtd
cNkbNsAQ2XjzEhR0xW5Y9q+82hYSao4zrKjn/bbl096eoAWsXfhEPVqRmAMc
V/fRFCY0lIPcwH9Hjs3Azy1JFaPyOrA4JAmN2Eb1mZCc/ohBARSatHdyaxvN
eDzkKS5alpE6WNU6+GvzYdNmO1szspbs0zRnevtljreOznpKoS/CwTfgsM5k
fMh4X+lXwIvcTyug4DrCnKLrnOFqD/r2/+AaQm6j2P/WK5aioF3zJOcrZqO0
tZlPNXDNk+i25JcEztPIxS/EzC5604wtiGrZ9wfKqUvaU169lpxREENQhpWT
2+h5gpaFBmIBXyxAj2u4/9tWbUGOcg5CNNLkzCwdBDIRuf/2C17Gtb4tH/Tg
fKGheoqDCXD/Jw6i25tVz3F1tyoPEKMQJH874rdYb/3v1MKiPtzVWifp7wyM
WUkUBA9uAvcvW6PuIUIobRMjMhwe8gE6kev/isv/GRNd5aynt+8fe76Kma6v
2asIO1wx6LIrj52+u5bboqW9PBiyaSqJYscBAiiE9Ii0aglWbh4Gt8zZrNC+
CCKP+3sgVJf6U7oXklioZshDG5HTv74PaZ7QdOi4YcJQeE9JoI+qMwsNux+m
oYwL/l3DHbT+hMaKFqv1gV/pE0MAEzkdN5KQOEYpeAqoRWjNUFwaK5cVJNYg
X8olZYHrscZguiEwB0sPTw6DW7qyl54bv5ophM66xcSxdQ/6PWtqwz+bmk4+
GPi5fFd42o2chtlLkvJ+uK6PZ9dhhBdSgEXCF47Hop4kaVTZ8bi000muZtEb
VaKNtsoOvA/Bda3cP3wzmLS1mmVgCONB/Ih0uUrtgxG98Ml/LR65J/8lbp0z
6j/qZNvJvrX2pbkja9yOuywbu5SfltfDpWGrqk2lke199MsjONsVX3ixVNzt
H0GsmSUf0dRX8Bw3TGFc9lreYePJurcwbzTk15U4kdF1RhdrvTTLKsg2RLHT
wzeTThh6zx3UHKqM2Kpv9loES0ErfbejHZyv4sGFKYiMQMFZRhJK8RpIY6Iu
wxlgvolMYNLo6PwdlzNnpbPmDT4eXbM+CXCDdyUfqmAeHKi6r3lOUSLYbvT2
8Qll6uJaJNPAAgkGG18yeAhBMpWALlTJyl5zMIEDTLswatCP5NFjfajH2/B2
w9lo+bjSEyS7rcngstt4wWZU5JFE9bwvc0seg549dM2N9gjuxDhhL93TzFxV
XcGyL67wwBdmL6oMDctpX2WCHplW2FSzCpWWdoXlxn8Wp91nOYUkNPOCckdZ
jlLC4NjM8f6zhPe+UYnyQAvN7fZ06uMaJ2rLrD7On6IWGDeOI026ZRJzRmJg
TPTDQy+eEuisN3XkzdlKFPInMwwYUHCU8lj0XHX4A7mKaI2uLPHD7ivjHtF1
vs3AXbPIXWErniBENZXGR72/DPbbUknO6C2o4/w+FtPBR+eHADvDUFUDT1PX
/8MMtx6VMpc7Fx0KQ9ChQ544+0Kq5oedAbLIAg7sQrty7BpVX4Gduv5KDvni
fteCDxiqsRgWAoQWIpjOkwBam5IbOY2uzSMk5Dxbq97ASu9xbn7PuPWKj4cN
fkuWVKmtursIc6RMbGD+pbTcqh2KnWaPLwkSBCXX1G7/jE/6hCRix/ugpxFH
o5aO/OzbHZ+jhkpsISUA9+l5mI2522Mzqupb3r+j/tzxD5UaYeOsg8T4MLkW
7Wd9AzO/kF1KVoj36eVcC0wqDw9b/YUcOaNYx5PVLxri0JPxhAEreRkwpRCK
2cDgiRleN+i9NlPa/ZuSjCQov64wyj0Tk3Sao1Nd/LpSVr4FYsljZfR0tV7Z
Q6PGFvwztMdFW+1/NMmJMatdWajDc8dikgXVophzEZnIHqxwn9a+FOVL5l92
WN3j3JZYTXHd3z+4qzklg38wrTP0EkTRmMoVQ2vf2tfMiinnBEZWaxhE4LeQ
WY1kkV2gQm9KAE6LpALmAdz2V6C8LwI6RUVSMSOo7HoaRXlA65mcwb1ps8KA
sd8qZdzupw6R3XyotRryD8n2i7PL3/uENOEV4Sutmej1BYQIdxpFwsKMJBHg
24U4f6/KBmaRF48ADBgLF+kQxdqvRT5MC9qxgSHLjUY5fnBdrydYNZgJmlFd
IlMQ0bN2FaGg2ccSedsjQUj5T8GSu+P478UIWZ+1XUgvBjeggLEM5Tws/BPG
7rHXQFi7xCYPtptKmCjRK7BpXJ0QcAmSnDsKdSm0Fe7CZloCLQXQeERaaYrO
LESmdyukI5IeniBy2Uze78p/r5MBt/G0e6/hr8sz2rRtRanIb3mEycI9DIeC
16Ukvrh3uzWN2YrgnRVw9xA4xrqxyUjN2rX3ZLHGvtbudDLBa6FYLD/mMMlo
di+YZWw9JuBlZ5auWSZYkpub+CJZLv2I/UHQSy/vWv8CbHY4dorc9zRSEwjc
XUkbZc5emi0eea4iA+UU6ZsIDlyU7j+U2lwa/fweqiqd/Mp5ff/8hWeNowa7
H/Ej9M+kJlTfLZJnXAcPhjIRNr2v6So7rwXeHqoA6jBux3C6VvCqsQGwtiRv
23sT2B6EbS2PtO1Gq99a/nEaF+2unX0bg9AdwdYbMrI8WkbjIpJOOPu5p66J
JPznGXeMQdmvRo6WX9QqUGushIBY9LvvIwLvQXbB0FfsfvXqLSTFwmDAWGUV
i2VFq3UQkJbaMnhHcceDbnIdmdVcckozBk8e55gLOdAww+sJUtHmPYLtfqU5
G7xtlHgCfe3A0IPe/+Ep0Ys651P9/MEVVhn0cZMJUSY47b+BQc75YQDs7LuL
yYnvZ6776BIG6BRHDTlPiANF0wzfME/j0qHj6tXoeVaJH3iwx9dHQGm7FAXl
sGPvBeKVTlB/4b8neAJ259BzHHGqQQ3nQIjBWPf1b8IfxPmrJUgwVP3Fc3GK
46HaKqxWetXTIWjGBX1Rv6QN0iYWNcqYULF31ci+DHTMiUGkjs84nd0A3ZF7
uUc0oOnOvzvMU5iSntocLEse8xj0vmP9iPWmeXX213Z+3Mfmwp/cjZojbw9Y
+xkuRvLbDTOZ57xX9D0v/6qLvkwbeMRn03M/GSlqLXMcqmwlKWB+vyjVvqjh
lFFEFvI9JbNFkl0lHQo0z8GVG1sFKvZZZRrp4rFehKiIIraEQCSWjFZjIPGS
bNk4Bf8d1Ka4GaxNkTOJ4K6M+T7Sb0zdBoDToipeP8JDqXnHGajwA/Pdnj8J
Ncp8o7hlkohKar5p5YbhIOFyfiH0PH9dH3ZuJUQd2SzHebx/xW5cWR0vMkYx
6R8twbgvK+ZY5P4K+hD4aiGoW8HOtsv/B6bTPS58yVrsP5u3MDeCISPFEDxL
LHWMJocaCxq0J4X1ToEiVuZM/yLvr+bEOeefmRQadcadnWqGYnfjsTZb42cu
V1g8OYbPUj3A55h3iP9XPUQMU6UmdZEv5DQphB+LMkSQP3ktxgfXd0DqBUV4
SyFS8K+VatKK2QtoDiidSWGQ3ZWTXZSFbbiRw9iexYScsqqGn1j+ZU63aM9i
53U0zCdCVTyt9E69iMMgb8fTojD1fZqfYhVqIWPN5psnttX8du/0oIRBRS6N
r6OP2Je0zem6p/Fusttmk66PhU64TKHgFL3Cyb03tRbzq/fkHXcnsKiAdYC9
zTXCRTjzO3cRhHE1UixPldr7uiJh1vrD1pByTfoEQ9tvy6O2ptX6wzsWDG/Y
uqE4JheviKxhwbZ7+dt6fb0R1cM6Q4qUSENQaOJGUpe9ZxGred2BQz/X0FC4
w3lui+9PI6VGTPdVPJz9Ad8drs9VpPIMpckI+z+jAOY+CE7PfINizgZ8GB9/
ke5OuOjasiZp5t8CHXknMdEfX5o/h9n505kkv9etFNHrMnN7yxybxDu7k/QN
Ldvx1J82YMcPxTEmHpIcHWboarE2os/3HYSr/YXtdn1CE/IAFy2rMMHc6UMu
ZVGJrDdFJGmwSge7yjyJ4ajb0UH/7Z0fzOxKNRc02FQAt4hd7/gy4ZaLARkW
Bv3NNK3K7NDhKuKy+9QQrOt6sogIiCpNCOBJsD58yL6uzpPLgklyMgfWwF+n
FOy+4bv/itqZIzIECFAwaK6qn5Luyvx8NG6sSBSBFmRn95AQ/vhJj2JRRxyP
hsffz5ezLcCfssGdq1tvzIxVjgQkWUQpmYgBCyTbzaA+XxDwVSeVpwW9s3YB
v3D6k8h7rh+xADUsE+PC9wCW19wL0BJoorfE9510dUfyGGm/SVTrSKAMvHPT
FwPA4LknUnfjd1ecfLZ5kV2zqCifae07Zoz1v5N0xqwFsxpCzDdVF4z5c2rr
8fDv1SRrjAbtlIZ6CZdw/Cq/FNpblwkNlpuN1nfhw4z2wCziwEW2voWqSw13
Y5ine0PVXe7SeBcEwanuYKAkqYjsfd2O3TId8cLMza/vdVXEO414mHG8CWK4
w0Qkkh6lJ3VdwVbebZdixtWhYd8ASXhFj1dJH5aE0JD8xYaJNeARHzdvxYBi
LgsqpuOYIUEjMeya8s2HOlWr9WN7Mp+6CkauszxJZ9N5o3K9VJY9xEGIFz7S
wcIqmq0POuW8N2ZQdsgwhzjo13HHldtClyhiK79sLgZE+8qz3MQYT5nlbls3
8TJPpM2Rp+UAQAMsDUpSI+GLVLHkc8xERxtITiWQODlpd7qZFUXc1tSWAoDV
q+nq8eTc2vFiJWMUUfRDCgYoWFs4s8VKCfBC6UexrF9w/ai09jjcBO5ob+UD
qPoBtgnvfbuoTEt8GdsxiWwycN42NodoIvvKv5H1qvJH2LmKmUcO3/fOlP1u
8OYfmDjTLD4QdtJ7eqmvoZr4VH1plah1pzKRJhsbbEbYjOILWGHSCJcQ+Jv6
C97Axqfgs57WYRnp8Aeq3i48zWe40EMMGhQr28MLJwTNYrFjV/Vxh2VSmmOr
flFCDnEj/9CX4+lvemCwwf6v8XJr6him2fA7AaWOqTeFW+W6kt5ataT+ACcV
V33wW5TvizvWZbtLXhYD77Lw3bm6g77EA6mbRWDue6IRlSedWuVjyayBfxau
wnddcowQUvaMk91R1EWd1kq/1LbuGVeHrd/EV7dQ/mMtYZ8BLx6/gmdNDMWb
gNOIa6ZR6sFMlsutPs83NztjRuSNcKTrI/lmSAoeqNIZ2StUrRNrMMU57WLE
2hyqQ4rFGpbro4LRs+0vAgHJMXCs+hicU2YjyW0RYB95rjr/j5P+wWUsd3hE
xmxQrQxA2ZLDtl+b7gQhdXNTGVN06osAjgAr8ibmeVrNI9zyBJ4GUHU6tGbK
ntg1nqc2GZ3475WSmeAUWR4COkG929J/IpIoCENvvDV9/ObWZv26XgIaVoct
bOPrlLYmcjTfQ0jNDtnQ20FQ0iHLQFf81ly80t/+61B925ub8K0RqlW5v9ne
cCFbUKmGUT/qD6llxE8kGb2LM8EaODhNjNMLZFSi6lmTPp6Z8RFi1F7yBrtF
wVWdw8Uld74+35D+udDNynZLUqVNz+x2TJwaHW+P5JZpq6WxtQHJnF8Cam8u
nWORybEhS9h/1dIfzAIGAISKhvdGp8bNyrPCU0ZWBINFh9PEb8LrABJJGbfp
x4PTdwKNzJXCnA75O3V5rQCjHmJ/k0p9/J3nqj6kmdzNzZLI1hazM6WBJVun
8QolIg/h3+b2KB8cd8ifZRx5GojFK16lEDAXh9IQuEKsjKlYr+w1JclWe9JC
m2SCcB8dcIuVsKBFUzA8SSawhyaJeosZttWbotTesPA3sx+KJCbkaJCwsygK
tvJzh7jReODuEaq0ln25f4Xk7BSbtn9ipQp9X9aFrtGV4aoTkGRaRfjlt7eI
wuyDWgKE6ABmtu7Np8DuPseHysJFCU3oMwdZL0bFDdKzFWsEMB5jJPp+GNTq
CTx2RcSihc7f7asRGZp+Qg51+sioUOqRC7zzCf81yYsX//V3oADvusOLu6Q3
gdOuM5Zl/QQZi1UsgXA8CGx6Fx8pQNHejiLCq9DglA5zumKKaUqbSIv3J3L+
wkIhH+KN0ht1rwbfNj/9F8yibmoqo33xPfuSdxXhCQYgx7fFLFPOApm1e/Xq
3pvpBl8ubsn5Q/ehqisoUJ3brGSMoJ2CQwKGFVtcgsQPYy1UqpVRB34GikyQ
AwMlqtPTfHt/aj0HY+DPzSDs53GE6sUxQ5qbn5K1tA5dyroefGTcAghG9HGh
In7MubKkInvAq7jFumqb5gEBzBBoxSuTfH4P9lSMzBwuxRe2/2dMXVQC9Jrj
U4MMra14s585gQrFdbDnSlgAVwvxTi2DOTJvoXvvikQT8R9P4nXfXNOIDMby
tB6Q1W3JL34rU1LduQOiXWDNKl5flbe3z/jB/Pg6ysgBfgC/psJyZNxgTrzN
K8t+R0iwj3KDW2uumF9cyx7ARs2uYTs3+hEHBwYMmiYntxq/MaIoVaBRnENt
Q75GC3Zzw901zscUiT0qtdQhA6LW5b71aZF3XvO+/qaSKZmRu7gEX/HzlAMb
0OfycNuwYwvMyOiyQdqTIbCeonIfRhWKqwqtiUbmroDogW3z8k3SYuZ5mtAq
YnuxRn8bn3C0CxQ0YarU84YtM2F6W5QENeuJFcui4qEvtYAkdmPu+YP8dCaL
vo/1b3ayCgl9L3LIBdJQHwVIR+nTXTQjaJvgLMcCkxLAty0BqG3G40u2oapx
/1wbTCOVZcm2SGXFzru75ljs/40N8lbFTduFwf+kBmQkVWfzZ00QL73K6s9w
A3IQFfpgyaCbcarvQXLorfrBE7tZOsQGwkMdkrFw38MVPQcpaa+zBNfv8YPl
6qOy6XnnYbyrNraBCNxSAcLj0d+FifcxadfTMyBiJ7OPolDzbCYnmr4HSArX
4DdVW2V2jpncaxzywxqssvJTTHzGM+9FfNZFhVSszguihzuDH7u0mwaNc5Kq
5kvqo+pXGvbPkR/pOCQOkg4ilLzpo7C71dLzCw7nEX8SVsXuwcF72jcyW7F0
eFptKkPkPsXzQ/19agsNHFUySqTZbKo5kbrzw54uyX/HINzhQGRxhqO+Q4jr
o4SasWCWmH02F/MCme/AikymPVG+1oLQKA6wwRAIx/Y2dK86ByNK8rF00wh5
SjJvaSpLEgyKp1JCl50C7O6OdDb1oLtk8nqdLRd+PVAQkaEgmHtEl5ytWTT/
EtbxDn6bZFQVfeJn0s34m8jofMDhd9DQF+RGrS9JzxzKdTV8iiagmz9O6ZpK
7K5HmcEfSD0n+HizTc4ndjwFF5u2cdwoNpH6yBJwnIz72InJiSmK/V56OSmP
JuKiyDyaUVpX7NvtEDfnw4/wvEtrOutyN2t/Lyw0zQPa7RU078uPNZe4rItD
0qMvKUcGLGEyDo+OoQ6fN+EDwMexFWM7RRPi5XnOcbSWMio4/Z8dw6SiaGIR
wwertsdPIN69pHaNwNYfsqbKO42XybKdJJs9/CkC/okioG+F7/5TuBeue/GH
SLZ1aF9NCfZsRFwi15ZB0pOs56e+zW5JpDcBd0XWjOQN2ZOfwmR1wnKhrLns
4hJTFSgUEKNH2NJdXBY2ADSTkfmd6K/lPEwe9QC86wXnNwK9wXFIWjKt6cOI
72YSGKWJr0qwEr2lsBTdpRncReg3e+L9FXjUlc7YFqcS7G+jcctMTAZelCX8
PwWRTjmTx3RF8r/F+c+z51Dk0SKK/rn2zuS51XvojT41uccolT4HddrTFdu2
uDej9lIDCT1EGqMs1AyT8wo42YZwMAYBk8DZMIOjbpYGlR/MGqFNnl3dQqTI
rjYjEJOo2bu2iqeRIzM31JzI5pprzmq65B1qT71B8h0jSuI36S4nO/wp1Ngg
QgveBvYNA/8W89ZhkVwuj0KwiATXR5YAHx6oiCeOe7VQ+LKCN+WmtZ+SAX0J
WA5af2Wn9WzaxFKujCWO+EZhQOUGPlHOrfhRCj8HoPIt2AQ2JQwiUIcFRNY0
eEWnf97lpf8CfY9u+jVYjZ3u3WUrSQ71Qy1KsF0qIZ+VjwFoJTwEo9Zmt6YO
48tin09orBjz4+L47Lo2X3Zrd9xOQ6LeyG+5C4R4AbjBj26VUOZ7nf+eGr3R
0oir8w7rlMQIcwnCjGKsIMU5BKiwwMzoxcFBwfG0CifEBpTxTpaxbYSXQG3n
5zgwbJZr50Oan8JBWv+yTkIV2ZnWLbvmRr8hgAMyjdpkisH8fwQdLCTUm2V1
hwNYQl6si99qdrBSpLLOVIwYLYJcZpaR9uBWrWPhnmykgqty9KXpluxQPBNh
J6t+9V/xbldcrjhh4cZDlqpscpkyWS7GDY0mqdRJz0j5xXezg1JaEMP1j9tq
LDkSY2BGilj/LffwfVXrEBw1wOZ5mCcR7oJiM6vJnPY6in4eFS92HbmWBf9I
9ZOQfNxyJQr8ooR7oBnBjTMT8s8MVJG86my34vraWxtX7+H+5hv5R5isc721
pgT/7F+ZIhjiVlzcXBjOJ2q17gSr5IGiJnKxjg8DKoJJNKXJdItiHPTcihIF
b5HvWA6C1aGCg++E53N//E0jZvOEcr3nbtlhrpBssv8TgtjiHikyUUlO5ae9
qbzF7oM++igY/zIr/GJ6Noz1BsEd6CyAV/hUx8ZttgvWMTwnaWp96vGaXKrT
zS5F4i9x4OWvtB41wnDtbuxtZeL2oDBGwaR9g4UFG82TaqQ7Br7pFZbNfOgG
EpisSir85NOyBb+WTeD401mXYKNP8iyc48tuLCgw8UaELtLWJMQ5YC/GbiHF
OUCA4ud6gMbEQgf4iZzvgA9EFHFvP4lOKsTvVFDYmLr/zzcBTpgd7gAUnmFo
JrXcGK63sh0ZNdew7SqmfO5OsCLLF0Td3P1zfgVzZaXDDbrIM4a6Wn46etD4
deVj8YJZ0TMWSd4HG70sBvKiyGWW+Uy7CSBFbatimMJqKBoaYw3xnuk9zUIp
JE5oPPPcxAULEtxguYyAr9dtB07OLuSbKPPoDtYSYHYgU4cRmB2jBQpkCDP1
GHbmMh85XmEjG89YSHu22xcLCQ5CxMAI4/BhK/coSHY+dtLL7MU6AWuYo2nl
+ExfUcmc+Vfl73B0JVVBH1Kg11orzRjZ71du6Bxeh/GKMW3ZEGCsXzVKvYLs
IFRgRpDGuvKCMjRfaXRWGDU9I7J3OlElSQAlEIK51aaQyIV0uEg28B75pi1a
tZz2YlMlugmRDmg+TMIn/D2t3G9zsxmqZMKU99vvlOIw9xryoER+yPNIQvYO
X7NMGTRkZBZUQ7ihC7+D/k5QsEy4IWFtvkas/n4MUyfduoIAFsg6ruSOwquU
8LbFQSAf43Dr7GQbsxF5PHanP7hQ0KODxKObkwdWx5GRpHS2dwNpfxn6PKD4
3WjTV4xkhl9AChuSee5oIFa0BiR4UOmhSmx/Nvn7+PR2kSHrgRpwqSUEy99a
qqaCntDwym0ykv9FuvePT6sq6IE8cOoPM08iI6ksTQ7O4CoVQkVffNEKCN1b
2cTal/9M4aCju2awPZleJBjEnFSH48PX5r1liyR5+yJFORUIijsDDEwgXGSJ
y2Y1KPdTlzw9vRsNLWAGUMZGGErf/tJ77WsbqrK2PwAU48MkGCYawnIhXVCO
B7E+MaRLsVDHIoGh5U/6NbzwmbU48VVILdwS6eirb0sZuaia7kxKJVuwRm75
xbqel1Mn+swi18Df4pyEihHyBMVwZrbulhNFGKfK3tyWObwfkhxsiveK48Sz
KH/uao2JHL+Ad31ROHZNt9RhD9C/0BtNR108lfl23oejpR40sOtBC+yh/7sI
4NKGABUcnUY8GnBetcTWRj4qhKna0kYxWVO/8K05p14dCiEAsxRbH7lSWv4Y
0JYyI1efsGi6krRtVESaN9NeTVfXM8k5i5x1YHlDPs8xUG4/qpWJW4o5ubQw
rFIkSOQU2pZIWeKO/UqFIi3P191eByVxb7y0SjE1bZ3vJPAf3KruEysdY2Kd
l/gxPIO0QSK02v4XKBYH21gH8cMN15hgCwwXKQOQJEXm5PjBRmGLzIvzb0xp
utPm3qXDONZNTkGE/SbBx5QYrMj8WdTn+f8QzBHcjMGzY/Plx1BojItGxUJ9
3p8UkTB9PkZATAdFTg2UvOwe0U3nwAG3/gYURDTQpieHCEorJDSgqYAk22Ez
e5MQ+iMH5pp6FY46rp3dh32XIrdJ0fMlXTZp9E3EfgP9Z819ZICjxn2Aqy6+
XWcBaisu4PRJ4AspxsoVlJEC+CN0fysH5FLQ1NGaHX3Jw6miwE4tVNmr1jaY
4iGqUoHIUDXfTQtRQn0inZ9eu0JyUvlrw9lzDPFEWkpXLo6JqCCcdYNtqYKW
jXPI9OXbeNbxg5nKcoYIRXPE5YTuH00hvx469j8XNO4241ARqU4IGhUKAIpu
4ItcrOy2TN+DSdYjxmQ2p/n57hud0kSlXVn7Sjq1ABPgZ2nPSLrAKXo/sKC5
VmVxqYyM4S8WmDRwcLaV9jlId2T4blsS8Qd3lF3LdKRfpgFpcEezAW/kNsK3
gCialdZwH/R2RSMBCtTaWiZ2XTy/4hDKizEjBMvBLId6eFQHUlIC9rep2HWV
q5wr7R2B9snaxhxNQGFSDmRp7Yji9S60mHEtNxVakDGHWXGbidXZwJey0LBD
lD+sMIs5dODxIt7/dgMAqbeFh9PsC6j3C9nL7cUmHuxU8YG8WaoJgQQszyz3
RuPDU2QuKk/1E5DaRYSQauAauCTEk0BJQ8MbObkD4A0uG+vrT751+EQMkuNy
b9wHq7xEnsWJ9/WS6Ay8aWjJdl3oQtGXshZcMM6wdbPeqwEzxTr2H8XikCgc
ZI31IjdfZux6jodWEyKqzrw445/EQI2CLyQYlOsDo5F5r4TxleWOOPRuvfjQ
ob5wt/wg9RxGGD4+/nqaQwdMB7kBRdj2aAMSgsSBzECMZwO6MACHYEoXVQIN
bKplwiqkXUS80X0Ip58hSsBiIPoP2WwAYqiTFlUaBHCYF4PkFH8RA0OYxZYF
4uMgG1Fieu00oAkkmNmPjOjshrCcq/lYA2pR+r9hZPcY1VDaZtdOziLrSWvb
SRPxVCw6xq0yqykhT1taOL2pxdVy65CZ8d9B5YSAzb6TlZgkcb+ayWtJukGa
/VcJxwVnkwHv2XE9G9bMeY23ezSSW0U9JiXj13x8MJUNIWrACHsAbLU8aoZ1
+Clg4yD5btXYrOPVCE6A1paiVdbl/O1jgfO0sYBU5crirEcHFqd78SZ20Q9p
qM4XsBzBHZqAJerww9Q8pTJ2pDYqenYNt5dOJkYYG0HyDAN/0E/+hNeIdM5k
1qxO7AnUTBua3HhDaFEWzs0vkFS/04uj5aBp8BJf+epVfc6HV/b0Rg03XMD9
i1h2dQGYSYa96mag9dcVN/pyeYIdXEk+sA2HiAeQtK4qcD4a20psX0i4lGkj
mGJyUjr4GOLS3PttZuITSwRTq69wyJZXdWIlTCgdrQ+4HEH62oI3w7NYsgFw
HCH78m0SibYmn0882fuGOxelODrU1hdo+OZAbA8ahnkwbGnmoghK7/GmIb1l
vgS4rzF0+x6nDqmvLDCVv94hSlr5YpJ/6nfiOwL2y3eyyHuc6yjd5sLMA8t6
MzgweljDiCZImDQaVJ/j4bK+UEPi+wX4Wu2AmDhw5lnGH2PnoGzD8a+TFtBy
Vpt254df2sbUOoyfP5Q+irwUK8vY+S82oNETkOwib0+94PYcgy/wrlTg30dR
2aPLDSYM/h3A+KHbCK7Q58LAbdHsQZZJsay1Nd6D/GSJ4nTEMetGAqTnn9tL
sTQrBceAyAuBd2wXG25yAikaN0G19AjJbC5WmEFl6mbAWB01Dd6UY0PLh37h
+CGqckW0CzlLQQz2pg3AqU4i2eAsi5MZ+yCmUcXV6awtXzakz8n8WA3ZcBk3
wzZf1iODUvT4itIyv2iBMsXzEtKIL6MPGLh3APKZcT5Iy/BaoFAlUCy6FZnX
g0PVp3blzQfVQ2k33f1oufKJcEjr2K3rAFOYXrtlq1q1VYTU3F2vHQJdqdQC
6T77ZzYOrx+81IiYtIDcJnh8s4yiz/ayo8+C5nb7ojtUvx6WhjdFibJ5LEAM
XgKC0FNJV4ETAGQSHjCKnq3aV+lE8DAaj87YNWaadU8/7Jlx0+8dDbGELXZN
6ZWF7BFm4B9a6AxcK4RrxyTk+1oiS5wbQN3l8qjD/Y6tS6x4AVBu5F7Yijaa
IPa/nT1s2x3QzRodwOwyqF+FVgMcUi4kAfOgj7j+wwkPtmXMDQnncljqhWh3
e4hUVObkAwcRSQ1JCMp8yWVDwZDaP2M8vI80DqsKZ6+A3RcY4vjCqPxG/CHw
9nIJVqxvmrd+qWTmFkQA7wmgulFmDFzzlvoZi7PdFudnoGJZxeY4R6iAcP4J
gqFj8FRSdj/uo8tbprUAeqGyh5HgVf5W7BRv3PcXB6AXAxNrmb0IZcOx0P3E
DPZuVdt5VOjcM+WXzhuFNcag331fo3/wdAJHW+SwHmlTtGT7XSV3F2FWdb/W
t1i4iS8x/LSFfOoZATR32UqJHf+pEkfR01HTp8SKA++cmAHs9cO6Y1jWPnpZ
xe0uXc1T0mSuv42QuGfZUKNFLM/x+4Jn2jw3W2K7MUtWDc0dAWf02uy4svCk
kIIGgw6yt9uPhYyGAEG3hOo+eZsYvE/hBap568FyVRYnmg3cyOuQXt3CmqyE
75zMnqUlyEvjRREp+AuSHzi8iHUYWP+08VGZR6rDygTCJ/ZeqSg17eCWHcgF
x0di0sNtFQrY6nvgz7E2J/2CL0T2CfZS5eMW/JNykMHaXswiNAA3ehiHMSUH
HlfcLcB/YJsRoHKf/bQ2uLFTt+i1qb4oLVj89c9F+cFtWBwbrPtm83aOc7Q6
WiIW5jeSQHdBN05zlkcYO16J+pgX0EXcs/z8Fajdo7zLyNE8JiX/l0ul7vnQ
CDa2rm0VETF6ORDeyad2o1CyDplAGxMGoQre+aZ5P7xEYpEi1rN96FpW8e/L
FHB2/QSKiKb0QpyO2PW/DDSXn6TEoaz2S/2Wf1R4XIeF5Vnm1SYaDyr2UzG+
ZHZc+2JuCSaUMBwnD1Bsc2FhmvHtetdcI7FaXJbQ05zCrVsqZMu/Ec4KZ2oO
VoxiXj4/mOWPmKJSefYvUYCdLsoR+jW1wUVXSST8B6jweBO1NDQWUyvJ5TKO
3D3nQuQ+1NaYyQ1h04l2apqSkzf62CyxVGmjqyRxTE4XdYSwBuwvlYv33iN1
LHk16dzHYaFBB0F14CQHwHYbAX0VkmfgJalfoaYff08tdSYfn5qdCUc7EkzC
gkwjpscZUDUB9iGZho3CFbEVshcmskBb9xtbdY8D/Cb4R2nMWLXPaVQ9KuHQ
nWIsVnzwiH8+cbxrmKGPmBXjq1qBkNtAnFyzpTO5XbRaQeWpyqQuu1Cenpzu
pF7VHyj4dvDsZQy0SATE1QpVq2t9QFzNJ6c6jFlXgX6PjlKgm9rAQwcw3NTX
xDnofmD/KvQa73i1/EI0FvOnyeWUP/uzZ1Uay2aqcWEPTUG9P/JLUgee9js8
jF7jyBBABGxuOXtUoC8poRvEFgTIQU8pmO0NPvp19s1oGshasV0+8OcyV7IB
gLBiGsEiqUmAmM6SQy5rGrqaxoeUzcy4arVc6h2R9LaTHbd+/LZmLBPPxBdS
DTRCFqwxKOl4fwgWJ3+11mmWqU60PxDPnCyiqqobuLacDi6OtYzHe7Za1dmf
hNBoAabeJHchxUqUwXhvpOHMr5I8hBKTKhVpdcLQAv/Bq8ap/NYyivajl9l3
Nr6jEfLVwe97FiDIopNcUZcuIWQeZ3vdJIttRzOVp3yqHo6zxrO/XjfymZtW
YsHAxAuVMF6GaQKxewymSXIQlrUQFJ0H/Jno039Ige4xbCH2gi2fcjP8BRzr
DZU9mzJ4pVF72mQ7OS50B+kzlKHdzwr3tv135R4mbc1GdpL6CD5GcG9oczjp
97et6+ByfFCrj1Ba6rMkPV65BpkMr3gC+AV5ao5OMDTf6d4lJbIjrsR2atcY
6mrSM2qhZzvNzALsNEZRB5QXKIbFHLMtW9hR+5l6H9QBJToFRX7e928DmTzk
xFLQfwEwpebM2LVHWM8A22Oo3XEMouJwGqajdDjI5T97FMgEZ/TPZuods/An
Kc9jYq5k+csbBiQ1WM3yPxPlbW28fMCiZFEYHXSDFK6ODiG7vpvZ+/1H9zLe
Ltau7XG2wf6ap6PjSzvddHWNGFwpPVRp4msqWiGa4nW8GzyBWF/0vehKVc+N
+v33hVgqcj9eMpUyo2XNvZPfXywaLY9woO2BdQUc+lKoqj1/g/uIgWN13/Ft
4Gz+YUePZkKGx9Ef8jRMXg2gFu8EXr4zYp/ptenjhV+jIxFTw8Dk/0vbyyky
ta0eTC+b/0ONZ0f2s0OktuIxe4KZYH9LM6N9q6qKDVyPIkmUEgiOTvRHXoki
X2svDQhieVf5qgGQqIkJHrToUvMp/1hJeaDC7mQEIz53wb+DPoZ8rBx0EIoB
YCXTNRqHEnNTwZsIBRBFs0K8s01lIhhHFuiog/vJFtmeHuUvtNrKouqu5sXc
FszNmPxULni0BcWrHXre/k6Z9uW6Kn5rbM1sueh1caGOst0/wdFTdFOKPqrE
LFH2bBVf9GcuxgbZtCJI72fDFzMab4K8EkBUwdcfJ742C0jAxYcmc0JDvQYd
Y2690J9ndNwaTAgKQO/LZfbT5g5kNxLstdsZzWZ2fZrCtA3b6wggoCi/B3D+
ErvCUOtduqRYA/gbUHlN728MOmzfYt1mi6yMXhzHSHq33xDSueDJdS9juaqJ
/pysmLH4S2XPlZr7bYo4yO/2XRTsQBeLa7kpnMXbiK+WnyShW6UdEi8tUFBG
v+V2hnMkBVTJkmxQRerO55XnFPqy7sdrQPWiRwovPWnOe2o+xQi8wsb7WiAG
guQxp8HN4NfqqOC/WjA0V6uRg+C0BnjVW6lZnkEfQedeOcXQF/XCNLZyZp3n
dqUZTmj73xc+kOAnpLutshTG0vBvsHgVgW3AbJ+dBeo1W3l4Umo9QslVS/Mh
LCtjGy6oJqQieWP7gnmSYGAzHBO+/ik/AlmIOAeM8ULxOcSLAYzr+xAGVTEw
pyjxT790DPfzqsF8ty1PAb48dytPgI5WgVyEZTGLdeURengqE+ALkO3X0IZb
CosLZVBZ+HZWR4TvL9V76b3LCiLFYmnRZKVZoCUBY0pzZvjmENStcwqcx3JZ
Etp6smlanAsISEA/xJ5XwBcTxUAbDMFtKmcIZnj0uXmQsN8OhV/UBb3RQe53
3KjhWTFAQtSsUBVtgPBWUB76dixN9ahkuvB0z32gegUE2TFtmO0np4jutG6z
5uedzOvTjDkV1qTx6DvK9P8X+WJArH/A+rL3Gskn0b/CWh64paB2SVw2KY7x
eXPXHOlX+YOuxDkpwwTgvxE2cpldFmhHjw1OJ/PQ7dELtusI6bMhDLM73wL8
5T3Bc8NlHveJdxrxdjx0/rEn9ZC5FS4K6RzO2OsZKaavkJijL5O2IbFVbX7v
T+3dl51Ccpx7+53di38nF5qlYco8vZ3SPbLFVMPmPLW/nrr2w2y3hqkolf77
eIQ3pSQIuOCfZE1Jhbm1zlQGtD5nsjeV1YQxTGPK2S1NkkzKxRkJMIGyUZVB
FoSME3AT8tVQP0I5tf4DGfOK4L3urdTT3XkRM8HKjY8O6ucedffCXRB92xqt
bKAArbQo+2UDvewhHs4jT3HJUgeiPuP1dlQMCCog9wtXr1Bo83zV5xvgROzo
8NYbGw+wN5NzCL9SgXTwyJGxT1y4j6vc6mkcQEnhZPN9Wj1mVxFI/c3ub0Mq
IxF21a/hGsOaKmG/t/OsiMtAwX+D6O5fj3QBfA4RLmbFRQCzBZwpWYAvg7/N
P2YJmvqa0W0CbR8n8tP+Z2DQv8JN2RMjBW3x/QekOmkvWlkhqwotyzbgz7RN
+gfdvvj3dZS788BUw3p375rDVadL/Oc82k5+Qq3aIZmcr/h7hLOCN7B6IFBb
2Lgqj1fGm/pzrknALg5RYRLGJtLbhuSsFUEVlTrt3WXnd0ZEfpcKvBTW8DOw
oAFkbC5q4em4B2xrNhy+8re1NqGQfZKqGnkw4Tl+qsKYqwO4oecoQSLRvHwW
a+z8cAJXlzIB7PWyhmEV+59nRW0YYKpJzNoTYWRi0utZfo8/5DxA0we/t0ww
B/0ND75V5n1BOY8PDnOnit6Wldso+gWGiXIYhsQOSmQJIOx7J0sDS8D+gAZL
7eANbLeV77QFFRQxhXOrz1Oiw/9eZIXSql82f0oq+jQvMRN54ZHJbOYKRfnn
AToR6QUJZ9gq0OXnaBus+yARr48CuwQ1YfHB+YNrSsqQWWSlKfkIPb+AF6oo
+NRqIXWLk2CAonG8oyrS7Rj6cXeogWjXD+x5Aqcacs22+VZc8ZMjNSqtRykA
JLEGq9JQpS2DlXI5ovjTsmLyQHYB2m2n8j49kXsJenLZkykRCc+dONwIXkI8
aUdaYYsYmdH7ICUbnPv6r665ODEc9qJNnfAvhqD+DXBT4yxRPXaG5y1YyFT3
dITV1uJEudoGOMxMeeQ4wZDvTbPYdRDEBgyDpNAPb4PIoxBCRwaOq4ik4+uq
VFpGhL3CWaEYZqsp5nURfDNnxszvW66f8vdT4shoqV5lWwjkoqPDYf/anPLq
G67wY94dmxmJ3BqJjN4pN9JJt5CmpnvVaendT+Nk5R4Wrzl2RLM4ql9sQUPM
3nfhFShDInZBNOu12pVTgdCTQ9pW2HUahiv4ONoLP5Bio36tlC2x0Rhzir+I
9YyLerbu1Ka1hdOMr2xhUx7GE1ZPhHAbxcILMwm3bTEAyshYS+IB845lhTIh
KePHGO5JqxZ5lpNy30xoIpHecJkGJlM+SY30w7wyfCIKTYaJiSw3p70JHrKJ
X4OlmtHPkeWYk3Fuvi8Qaj+iYBrnCkRHT+IgryK3GxN+6MNALeG5QM5hYBpp
YZ3wQ9E5AYYU/EcZi/81COObkFbaHhRFHJY4whjQ7LsTomFU9EK5qn12Wndu
3Sj2lBtC3zYfH72rJxGF2NicUDna1Z/AJoyknJTzS5nqpMwAlEJYHp3/0EUt
7ygA37n4TUlVOuQCRGYvUvOvYmEOfhoFyvJt/vTheJjKS6rFzvb/72PLt4RG
n8UUfR7yDIRCg9L9pATJaFstqZUajhgSVxRHcAXDBPOeJ7ZGAFoOcE+sv7Mf
b8sgH4hNBGMw+RJROBZfZLhZ69GUWCWT/A47d9UIpYHusqa3IdY8FVojZWUW
1yD0nJaoyxaCJboTkWla0vVa8OWzUvbccTH+2CsBoCr/J2hz1vgXJHjovW00
CTNICOWlOQqChGV11meqHDveotGxUr04YZkqzatBuZs88HbBbRbMi7RrqyTA
tSkOh9od0TL/UrNxueC5zpo5OdlsqA6zOrPdx0HW5YJFIcg4chgp7NfWpn62
zFg0765VW4vk7kDvFTWLR3YAoTVg5prx0fINkcTQ8EwtTQVVtqUg+tg4Q+tX
JuTbdxSwF1nFjJvRyGuwizxUOH3SDbJs8rTegBMXsh+jKMgDtXdHY86Lq6v5
iDEzJ8uZtcWfa4T/M5zlLW5QjrpQd/vxD15CUAXv9MZtM8dKE+KQ4RRRh0Rp
NirbhcO2TObUzFbT5nRE+n8CLkej259+7Ues28TpPOcaK3ptuQZ9P+RHYTUz
wkUPtg8gJFGwvGknX4Q+uEiTXgdK73/bXMDqsLcsLhUldx1tCB/kxi3SsQUT
vUXY0WjsDtvs+htwVliRuag5ilvpxwVOrroOLJwmEEkGTW61e6nAJ8JMcoK8
4HY2Xh965QBRr4+Le/eY9/K5RmrTPPzrZclOzPU7ONiW3v6gJ9K3cDaNmZIy
lzZkS2PJAEEpPkNiP70lAJhssfWwkbbeCMOVSNTAGXnHYfSWbkKypenm8rKH
1CFc5HG5+bIt3l6trDzgJXOHjOSvyrGJphzyvkL078A5u8N8PDRgFGNyqscC
5ibasVcyzI9vI31Etwz3EgiC93jOferRXI/e1jO9o8p8q5Kl8zVP6shvEf7b
RkuuKypp9h+/wlEJeVQnb+9a8G00AV4AC9VOBPKUpQILITK0EERug7JxtjYe
iMW6zW6KJ2sw+AbUpFP0o/ygSLJkZ4A1814JAH8WwWlplXVlxcxCZ2ix558O
+VYt3iApdTGHZR3uzNbTxYZEDDzcKshSWnwL1MFps0vGeTZogrHJGMVPNvcO
VMyqbzGy3pvx81uTcNU9TZ8axFxvYhU/ziclWEJkx6t5dCvsUxhvFwC/W6wF
Wy0TxkcPWVOuYsDIISQVU8VLy4cJeSlWnUJooC1HXy3ow/WUPJufi6tVMYFo
xgtg8NueIaJjUfTGevh8HwEBQzeAyx0b6YrCNfu5OPrOHVqeHXW4qsXqA8fU
HZGzyzwvjFiA7xodsSuPlQ94+KWY9mCkj3+0oDU7410NsAWQtjzIXQaVHLM+
/HLCJnfY2M5Q5iX2FqZtAlWe+FgUrXOGLmtbWpT6LPxVYSrgPNV+LHjvM+Zi
jozxFz+WCbieIyngEqfK1fKL5ySpEn0Er9TaUNbx5JeLI6dE55AkBFjQu/+2
nFG6SFCalBJezZbdCrvaMnr8n3lmZ4TzPIy7LOCJjZz72Zq9xQ1uaZfn4sdq
hZ+W75p6fq1F601CUbvC54ErENMqyN+EIeS4tRQheM8bisg+ew5fkmlJoe6c
HpTGyobHeECWHonoT/3u1ZEv3l9tzyj7QMiFvG/p290qToTmVDE2XHELRNGS
I14AYSBTu41MDErMzZZNGLbIL3AmVrpF2DdnkUClFR38tBRg2mTi5i96rPyi
4zuoALsFPht7/osyYson8rszuJrUjaUl3jnQpqi4oEjW+Q4vII540HarILCB
AhXb2Ce4lWcHmsIIGHg+bSU6tACzFHiXI3uHI01QzGribyaAkxE2b+fXaq+E
sb0OT1SPeposCo4E/Htisw5Ih9ei7veXLrIAyfqaR0ZQ19sJakMoPYMDG8Lj
xjdcxXeF7GSsihviuvbVm1WOUJFp2h1h9VxEHgWGRMjF6bxfztJEU79XPVv/
hRWshErvtYs7wog3ekbXkoNUwG3Gn5Em2wTzx2r6FxZwg+MqZlXKIyKrNKgr
ceZEQPAoSxd/DeZ24Rsrfx5tRSSJ66oMUOfrjJHNsf3UBBDl10wnlAGZdVJb
IHrgvbO1Apw1YYYBAB39+oWKxAKVLRjJQtmYKKjWhmpVoPdMiXHCQvD6WIni
aOuIGFeXhu6FGPAU+GTKG57YqHOPeEureXvTn6PfWmoOiOb9bHP+70i9i52j
DnFFCOj5CqHRNvkaSTIAYyw3WMRMJ44+ZVTGN+47zFF3awnNzAK84lLM1QgU
oNP3hAuU4MO/gKMG8uJqANnnUxUK/b2nXYdI1jnDwRdxEV8NDmuDRzfZg2tl
u45uiRajCQRlsNR3LgQ52KM1Ir5At3qvmpX1XvzdnpsnyR/2Ye/+QmQfvoSh
9PQu4SuaIQ7Ok4dod4KW+mxrhoa6g+T9wdTjT0bCRAI5aouwJsSznK1cQ4Rx
eCX/HhyYnYePJbZBfV2dI35ETNYRXV4/ftoz3nk7yuzvKkT5sCEL2sNsf+mS
gGFTUrfpz1Gm3wtjfEkr+ZZ8mH4nTPihVRMynYVTecO1kKJ/mMYDJUpj3fXT
l/zS1OHth0J8VCJpZPcLhfklLHy2c2Ij5MirCzQy8j7RYgBbLQZ3cIQpVlg5
3zuy2zAOgK2zMwtDPyCUblBXmV6HIeNEZZ8Lgrndp0GfKPBH5cTO8Y9ixlJM
lAZ4ne++m1NQe/u+xC8f3qvV3aYvQCSPl+E+mPR+BpyhO+QUaQ4vaYrbnCib
vMXuF1CJn+qY20lrS/eotQ6w5DR++qHwCFuSvogUwg3ctSYekgdTzAS/olvQ
K3o6xhkv26GB9M24DUeCMoTAozgV8MwXr5dFbD41J5z7IqwU9LB82LA3aqk9
lhoKiU09/mYjCtvOHGgzwFNOYXdLtjIR7ZquEwWPqh+d4qlI20N2A8qDF6ou
BA9YgwnabCOMtBCvgCM0Q+DWyZegX64BU2FC6WJO36pOzpRNyb6KioPNtUla
8v4S6cKh7+NuSBkMragm4QSkg7pKsk5GKcC74uVYsqnmXZKvJLwxJau1NaaQ
d0y3c5jbsnzwCbLCXtN6ElliT5csABPizczbYGMZIHntUBv/TVRchbmIucl+
rDKokwT+s2JznM/Ll8EYxUE08OJkMegvaTdFS8t3ta7uddGeAZhWPt3f4/bc
8RCnsAUj61ubQfDrYzi211Kwrlx6SDTnUDMQxJsnJ8bb1mVaDo4Qn2r8TZjh
FbV/4lwcG16GHH2XtwamVZnT/YepsvD7Wb85aIsL7RXQEd7XuyGAR42heAGQ
7w49S+aj38fsAlUmVTzQiKtYQGwYqTqL/nrVmv0LVnuCzorFrsGnR1nC1v4S
uXocnXkVtADAhuOfaj3AmyR0iiBQHJ0TY6RVwvVJWs1ZUnA32Hhbcb/9q2GA
5qglMQuThJhW1Qv2akD4k/MTv6yuXtIwvXIQRC0RXUrD6QeGAhS14BnZH441
uX5OyuHQmggH1Tk1KMGt7CP7SRhBptROM9Yh0BOfnbZ8vxDJ2SriNgwymj+N
2ZN8oGY05YHucU9H+kFBwF+WX5sUwHcu2felxGDWITi7Q+36n2BLy1L7PZMA
d1rGXCFBy7M9WepNsuCgcfZK/t6W2JymgYgzq62fCjHp1k9Wltc3G1+CSD2X
rhmDctNC4qB624bs2fg7lBiGgQEaguv07/QRiEI0lJwjP4P0SA9Sqr7KDaSl
uwt5YfsN0HyRjBFD7HhQB0b/2VbRY420wPlIvsRWkCDDVQ24JDkw2VtoEhsn
AYeX9f+Q1LT/s4umqTUdSJZEwJJt6AAhBPFxEOFzHWcqsx9i20HN11SYgDfG
SDnDcaKoVFk/0Part79pHM0GROapkrOfRH7YSyE43Ug/PntCgreOP0tTteTp
tjkNKX35cw+3Es8GtZgNUkoRkZolKzD5+V3GmGuZjpQbD0EirxuRIIKh0xrt
V0PF4crdLoSv76BuFJxhFxth2XS71tXZnKFawkdgPNV8bTm0L653+C/SVY9E
0AIOKZ0LMk2vdMWEkn/g5pSOXuBQ8/YfNlDkpFqgeC2SW+CDkJB8ck5yBquB
QcDqAhkf1EA+3p1rDhU+vXOQhtYClH+v9fV7O1CL5voEdcCMVSDh/WCptIgN
chFM0aQANXhpiJaisIWDn8azvCkXWPZCSs5Phtqv9VIu7R/oqqkiH10y+EXy
8sR8TF9ERszguHOBTOtDU4FUO3F8GJNAp9o2EHJ6xQM02zki7394ppJL4zJD
OBxSScqDOB60q9dvvhgVDdRfca4jI0UR40zh2R9G47JGZkh/qrkP+hgtzif5
aGdwuf7QweopaIw7Vj1dfz3FevJJV/FE6pumPdiDEcJipjn8QQ70EUPxz/FV
Bcs3ptngCmAp0S0TqjOa7M2AC5mzoTNHYq2O1aFLJu94g9ohXS4dD2CVAhs/
GE84OjUaLzoq40xMFjJTZUlz/SjTV6CM8ehYswIStehfx0KAzFs12OwNOejE
8ElUxgK5pCFqyMSYZ2XfhocimYAOMCNjKkUtAZASsLm1OGYDGOd4z5TmWIEi
82t0HT/kiKynyeP8ivtuQBZ3t1Il5cyT8jTEWupKcDO54kiSTFbvpreS/exW
a2EEunaDh8EmqTXuJygV9h6S2i065Ui6c6FXXlzSbx//sHUIKL6BjzIBHLxc
xMtKGCDuZnSSQ6cQsk1IjiFzn8Mikcal/iXA20l2h6Lif0Z+xTlYQGn8gxBi
NBqfvqe2o3stNo3uWpY78BzxOIZEEOWe8kiayBRkifKLbBSw7ZUhpvfWGJWW
o0bwijIOhLNKSL/cpmruHlY0TcZs6RFrZdarb23CS0AHMUMGT/oqVeHNyzh0
3rydxUZCv4y27ZDqqkZE6qA3kjcdC6NI3dzjHr7km9CSOAahdO0C4GoDWH2x
Z0uQVmiEm/Td27i+rEf2qFWUiqs3rkCipzRpRPZGdO1QAEOHfT7mLPV+hpoX
ta+g6l8p2fKVCBbTV0FSflDM0A3g4qMgOw1kRaP1eE+pgMTjajnBodmFStly
n385Vleg9MviSafMQqlfaNX/naYzuid9DcDMdrOpTT+sHApJtz/JnN8DXy8O
myDqE5h3i0OeZiIIfhk70LX23H/MSvKymnazRa5EI+a+k7yHlAptNrXD/U33
lmBwXVcUmKvU7ihGngHA7+nAc3Nqjesb26IHvFwhWK/pwpv+hAz33ESHEqjz
hxgAM3XwdqV/dQ5zHL3//eLFyqd80bQbMrqqn0LBqCriobmzeh+4/8GLR2eL
HEKW23LnuC9RSrfGDzPCWWPRJ7L4YzSkSWWTtEjQEixteVbMMAfwUxxuz8g2
b8EUweYPaGk5DFE0DJsD4dUZ6If9YTjAbPNF3DDjKoIms9kLahZ7zuCzWqVl
2ifbbvzAYYHSPwbUn+mFFTrHGFyj+ly3hCyCZGcQhhZl6SJYUCZ/UOgCr51S
86fdoPoQ7nU9r1Zzs6hS4e2d/C/1+EadjKt4sqbLiCkR3b8pMJbBXG/bOUkj
6V4SmzwAAxgVdoiopqzc4CQpXEdXAcL0c3H4D3jGUCBzU+633mbMtf01KmE+
Y+H4ACzC2hPZomxNmiIigU5XI1VaaznVPNY9Z3C0JrWWYwPv7EbK3JXns9cZ
pv3PcNQoFvjR12iZaU0hEzD2RoPVyATOdL2NltPnP4CW84B7qhaUqVqRMoPK
A/jbPXwENRr+jfYOBtiTPzQ/wg3dje9EqdbNtmDoRKW+D8VgJun+CFJZsTZA
sE+whTpz/qgYaEg0bTusw8ePtMA9cPT2l/dLGcvysnQYEIZK3f68yG+zZqPQ
4+VinyBUJ9Qa2APpptvk5RP47tb4L3KoheC5IwT9vrtEX+ll4mF7BXuFHkqV
dm+IzbKI+9wrjqw/2hKzu+Bu7+2PCzfMxQuRyreCls0KWCbZED9rVK3pYSIc
mNuG4vSMrKHpggPno+4ThKA/DequDVEiAnqD+t9Sw7M/0bU8gAa2HpyWAfbG
KwIovf9GP0KhvphwBxYBBC4HZVN6jNDLbSyijTofYl0o1neop7y74LvBnHad
tY8W6WBhn8xRboTqBJoGj+D1g5q+SuqadkFBG8lRm4oBfIFWsyfe9lc9S5Ju
QHXlhVntoXi0ktqo3PLFrkyYucQof3wxf5oSFRrjmudc9BDWoEcRYDnHpFXf
0SDRxIk0qqqwYCPAV288+MWLWGTbrohbjMXYRkziXjKSzwfUdtViUb0Nx+kH
onB1bnf/Cbp56nwd0YBL3us0MqkCahLYrKN3zjL/HBnjAoq7txwErcvmpXal
0a7HWtLhO+UQ4pvz+jH7rV/veVXvSsnjX60qkfY0v+rWMzXO9ayl9T8niUQe
VtjtLOZATmHsnvKRLOyfclkkcgMu3gmW+7nKCvoO5y9mpNhTQp3oFXcHxmlR
L2WMr5VknGWLUxxflLv1RWtn48mVofYdbtaMGXFBuIVEUeIxifM51vnRU5I2
jJV40o7QUsXAMY+a1RV7HYXzResE5ChpQOLAcupIZGKEMwa8JymZ9+vvAQRm
wXJa9UFy98drLhJHouzMYDvi+JMFosquKZAj9WxN149Adp+OClvDkJGakvKk
vPzInhkD2h9ruZse00vqZnPEjc8VjlvlTt6lfJKk2rHwi/8xodcaSyspbRSd
HKeJtZ2IzbYfazFeRyuJAFldh09d15j02nb0dVnlUJlnQrDq9u8kz7lMdPW0
yTL40tuRLNhu2me3wwB0b8ARLqOLtvwxOM39sbkzpmAWIo+GIRR9P2LnImkc
CmWU4+gnCZssTuhwXISgFhQO1gDyMs3ME7U+Q5LRI1Zxwaq+oPgZsB2k3BIX
j0aK4BuLCMbgKGjfGHU+IVn0kwg3H588ueL3+O/iqQ/jKpwAXfa8HfGwWM2l
XUc/SCSezQd11aJelqRU8bO3C1ElNa2El15Qsc3rlDOjKn2EDbEVMGGtFx7I
NTycsz1mNEVJlROQQVbA9B1JrFGeL4dpTmcI2WCQV1/SDU/kn+ks7QpOzwqe
yVbbDnogXlUjm/5scX3wIcgNPEmDOW5pqBXLSraZ1D7G0s4hJ2JfThKfbSaY
RrSk8c6T8c1YI9dbBxKpodhRp4OpYWpMGHC80sen+NJxa5C3jQc+sBMezm6e
zRSKgyRFmyuXQTki4T5/p7bI/+ey1aoy7nwex5/Z3VSJx353bfs9BEyO5sF6
zo93dgZgB8hBh2ZtFxGnpEM7wD147RtmwWuOJqMOHaRHN74oe12U/Klzazdt
f7R7G3zciu8FsSG8Bet+MCmvIAFrdVmmYrUlT2DVGjCg/ar41DZH2ORnoLJ9
Juwb2Vp2K9y1rrzeuVjJcRP30Gu5fA7AplSws29iEgHc/KF2rwtw75b91AiN
sh1IeDa07erq1Yfj3sTlUKny3nQxkrMRTGldNdLSqwcn/5aOoUjabUOUStjv
KxFAz0igX33jz84vClPrriyfG1lhdrweyrCCi+9RcVfaj0NNRCFG6xL6C/Xu
UcBAIpGmKkP3VrSHaDqqEhEWDP3HUq3G1FAk4PE3DFx30lb7hi3Q99dQVw4D
ehPXOdDBvgNet7qylEKDILp1pNMDQcKuJUuCTrgU6M6R6Sv4nggh1WX9W5bg
8XRPn26T0cHgpn0uVw3LIcb5JaKReaXi9sJ7IojfFvXhpylIVm/9zG78vMdh
6P4Mohwg6NczGkLoF8SgsOP99j3eJqueaPR3G7x87Im4evgwiQsiv2dFiMDo
iLT/JYOQ5m7jnGprJT5bzp9JUPm+nk+h4wUgDD6gl4ExdOJ6EnAE6mX/idz0
x5hEgnWJa4y5gnYRk4Lu9+xuzyw8vx9l8RhZnhP1/IdKUaGCTlao7+lrwiwC
/H0mzOybmk0ajhnAbJz1SGklg3gezcUCLwMUY+rELPkqSElzEzOILJEiykRE
PoOEdczscioDxdcxHvRGX3rUgk/kkvFz2rUH27xBXo6nfOWhKyjO5zEEM8tX
DytlIEBu+o1yqkBPhwByLK4NUJFGGpUp+/c4puH13m+KhZIcAp7jWkzUG4m0
fJaxfWxE4IbHFjmR1GJycsTanCpL9HclVpDc1c2GnveLpMLUpmXqfz7BjtSe
uX8NvgKBjFFfAcq/khfXBl+ASIo1JBuW7W3XDT6Ae4to0dpFqmYGt4+2GmPO
GaoY40ZM/Mri2VcQupgcnJh/AptFMwGpVGb4X0ooohy54LGL+2yKDW+QZPKv
4D/Jva6jXAQ9OnAtIJIAM8uOa402IHeKUDbZm0+pKfsGKeSPLyzUE1Qmtsbc
36upEpEo3MIqhy2X262CQiqKKCoNpEpkl+nDjXz7xDer1qEClANeeJvH82Rq
sL3mnsTob/ImkKjE3/QP0Kt4Eh5srbSjbreur1OCmnR+S/vtOIX+4zQ5RH4X
RKAG42EkLv5wGVZnhKVKVDoM5p//n+kvWScb+slj3t3c1bqWTL+ffmXfuWI6
7m06YZaRYHN2h0gUdKu3ykraWk0KkT3tVAuPQq/+md4Cs+SM8VA7taZto9u5
EBSXlgDmYp5EjI25ityhnEw4ZdhgOidkNs96B1iI6ulsfCaXQfJd5ye3YvOV
3ULe0vNs/MUZ/NeZw1+UYljyhL/RFlaKCf2Ufx+UKafemhceuSlRwW8eRrOG
eJnVdB6rVAgq/P0SxNya01OvuUZsNUM9ZUMo6TjXtodZpMeyJ6Zl/5p4pEE5
qt17hnHzjALcy5zrTBXbmWsZlN+aXfVMUi1GGk10PUXuDZutmiFbSi+3GGWV
G5CdvL2Vl/M+nEzrv5/ME9aZBfeIAXDb9r762dM+R4zYwXomu14efNuOpKcs
TFkNaCl5YI+JZKWrjJMuw+gNXR0DRi9QQmbaGJnWaZT9xAg1RFEuYTlkCww6
SFzfZW0+uwKwPBkjAYPjsVya/qwjhnSCKgTKxyB5hyJieJ4wHR7W4IZW0F9X
XmKwpPRR40DcPAaLt7BgSgrvVigliSwVXId4J3+0Dp6wdZnlNMCghk2dLtMI
BwvKGkp54AVJnrWgjCfhV0ytnP6AChRmbPeRsz7SdmeCaFfEA06DN7r1m/Qt
vAs4O1yNxz8vFJ5rrUeO1ZfRxPtBHWgq0+s5SWVGV3M4w8i4StV/0w1y/kPc
sVThcw4dhItTN0YNae1T/m6tSmvv1nrLr+5xvj69GkJbxQSF88oADwFvYSOg
ZaWmqzZ0wYLLyAGuMLk/MT0yK4aMuS6RRodO0UIsia5yXlyTHssE+iRjYyui
475uMYCKfL6PYCOCTXHKuz6upuQ8cfpw+VlBgqD3C3mztDg8uNpeC4tsrtBD
hPhu9tEr99AIxBKmgZH22k2z9u5yFhmqSh1F4KuakUUgGJ8wtetXt2Wy8NOi
JV99r5kIVKBd32t2s9hc6JVqwf42Wrwe/aZvulaLa7n4y1uy1Z2zgiQiZ1HT
5r3pil5A3XNmtRv359NtQiCxefNTTf6D9UtdiOHvlfbuybBe3ITJ1UvjbaVU
J3MNiHYmIgZc8SzPKULAci40G9gwrdZT3luW6yxzbx3LnZ15lPdarNZAm2/Z
i5LCN+JBZkLzcEsCUyDPSbhtiITWolqYdbqtXwCujx7PUNmy4RhDlcqnALyP
EbpGQewygogV4xR85suZaTRK1WEwukfuj3NXvS24HoyMVJ7YjAmdLISBG3gn
7vUfKICmMdHmJV6s5gi/32W9lGhfpvZNHQDKEyBa2vXiCAEnJEpqwo9mgBV1
ZzEGZrwp98mosO0RcWMkMUa1JgE7vKMnYrHUflzerkDZJOyMMeYuTAB20aiw
Z40KAiPoUq63vp2bWdekE+PV663TSyv4xgN+cDyLzmwx3VLVbG/BxZuWf3zl
G/Bayk3fwvOfw5hbWLGNTAcRfxpw/I/09XUjg8y8H+oR54mdvmJVBNaW3Wn7
8DYYHJhqQWpJTpvKifqrnJfAmTtELMY151fLmyo8A3+6zDiySV3Xfs5/DG1c
k8CBNDyClWYaDh5motHiRXxx8JbB+Q4zaXMnmysrV1mmgARh2bgUpLzbqAH/
Oio2EGqKdXtWJ6NQJ3U0GcTgMCcMYbEuUjndVLCJBYpZ+CosWev3Wgl7Tqtw
en196uSkkKOc8/6H6VwdNlK0ffDZKfdKhvttjPBs3yCmVDJgNmbUkyqwC58H
UiY4LwpakYCuqRKS3U4oj+FBZyWaw7o28dn8IgM9KhqAqb4uJyGVuxCgaGTR
ah7/h87BmiDXcm2jsNNZSpht5UmR5nyi1uGlo3ljXFmFqWbebh4jLWbXI8om
MGmgfqqkJAo8l1ZEdhnRuuPqp6VYgS3pq7DUZ+wrHSy7KTpm5OmpdXcmzC6+
jgsQWG41VqNsjb92/laxNvGRw3A8N2yTwtzQN+xJzhgcrENimf6yEtI8gKal
jZRM58aH8sx+G7Hsef9te3YVAh4j8ECyTDIdewyGOQ10NwzbjlBWXsMrl5Wn
hYWhan2yJwk/A70IinWI3ZCAYHvSmuJyhkdKHwwa1KvCmoFvxiefbNDp14Bs
Tut9cyxFvgHAxlWR/7DgCW+IOtDFIZ5RAcy2FugL8tAvMtIcsjEIM4qPVVR9
EklOOQrA9sOUWcUGtt/OTjvh0mm2jIVWW5av0cZbp23cZVtkmpha+piMDbWK
8medQPP6gr9K6rB4oy/Z8DB9e5yMNLO5R8HKvqB1qmYmb6Jc5e3doKtlzYGK
FolM+v5UGbviz2C6u/QeYv2H1CaxWxczEWD0F7NPRJ0fxjHHgVvM8zkZUlQJ
R+Qc/mqqHZzwWjZpaVpRk9vU/iXJVvoEUZb1MQXf2MCbMjv8oTsvyoHvEjeS
qTk4cWTH6eIj59WJxy/VlvGE6ZgFEDBhM4XWbLh2ROj9qmW075E5YWVcqL9F
hX9g1cSKEKArjp4b2CKBF0XloGY8uAv8jUpA0lNLNDJcH8LUlVIRCNMtqCDI
wPa87diRrlXJEK9w8u5x16GgjUGz5YnFYAvA6JiDF2BYpquChF/uyZT3vUGu
dxHlvc35wKAvnjcyWXiyOfPv20Ky48A9Xm7OXxf0r35xIW2r9gwvH2pOPQeO
JBD3yxMzJp5I5pHfMdx6dz/sViN378OWavkmygWxZGy72jCaEm+EzRRfx7P3
+8ss+mE/YEpHyq7IK0n+q2wKrxo0ug2QGdY8Mfn9i/deL6GaLJnZvsISZNQh
MiZEtekT5pgJS/QrLJNp3luWKBWUWk7WnXhkkXX1Q+VtaTZbOFItv3drava+
hqFyIgiQus0u0z4REri/bFTnmdCX6DEEDBjC8wa3Bmqw0Py34p4Q2pHymJOD
PGgzzjD6jsxTZlGUAUxpWLr2lfNySiKvERshqgS/bQECs3NznQ+isB0w/oVH
jcRhAQaiG9b//SOhipPpM9KWOQpxn/Qdl36Be+ML9M1fsd9CIh5Z7xC8Lygd
1+YNhtBlZsCuuyTeCdhIXuup6QK7l6CHGOPAQo/CeT78gfLoPZeSgLtMJiNL
EVBvOXhwgj3Ik4SL1APCkMalB4iqt7cdzWGfDRHhK5cndJOd505mDpC5uy5L
QjTLPiJRNkbQ/m0vKZxHGkqHL28gC6vgYgZiJplNs6lJREdoIklMBncIwCqz
EmDbar2SiL8lsuEtF473Kl8YVlAUfuDvvnciBM4XWLslRvGXuolQl05M0PjX
VyrRy04OtkqRHXnjkLyMeOqP0SrCVtS3Xqw39Psi82VvxX4wCPFbranX04s3
vhWgbfYHU20LLwV1EkVtnDspcbpLwXIPI4Pcf9XCBZi19TRAdProIpTiflHe
/hdNVEhMb6R3zzvy7Ja0O0rdSAUF5sN6V3cFNYSvrxPVN14I4lTGdbj89lyw
Ilpzxo1yTEQZvG0t5AE7biWaAE3fVMx9TgvoXutgWpnEX3m2HMMpfRgjhYvF
XJ2PCd1kW8onFAUFEYZMFyHsDwAg51yjkFslNOegKU5QZn75wKgyiryKakjn
mjP+6H9gTxo5oOdDyPC2rDarONUhQMAZImAi8vrLXoL0kdDfqmFQ7ji20nBf
B3nhT0Aq47zW2TNip4uxZr8ydb9g7gcUQ/IlLLgkC6p9g7k2F+q6Z2P116Ag
hmYSpF3ACpEGFrng9B9Sf+cU3Pt77z492n4jslPYb6Mbie8WtujXezpHtFd+
lXw/BpIRxuiC0Rqu0xD1XBtDq41mZe+tcss5sY8ImYQmynDcrr70Ij1+x8Yx
kAGRSm3OJLl5hnd6yF2PQdFowZ2SW+9nABrkKlWJ4EdUJYNRSJJ/7J1u+GN/
wDsRMUVSG9ZJyDBfQXlI53ViXQLjGAXwEnHCVcTa2Qwrfkkj1wmWC6XKqkJ2
1PZpVnWlOQ0wxlMt1STvKC4noqGNqpNQ73lbIENuzmlzwp6KyhZVOTsyJgIa
QU90UgHPWg4E7L1Tsf3/oIxaj+0bdHuPl9WRsnv0PXvWfnwBnn8/+A6enmPk
2kYBo2hWggJ7L0G+rn19QGXfoMY5UzPnwB2vagw/sAwRZS3vmkcuJYKLlsZ7
AmBaR6kF3ARoWD8pfmqmi3RyGy4B8LLoY3/1BozV/6/msJnTZ2FFtCSoMVMN
2ZcR33cbko4hLj5ZrQu7US06DN1AC2Go3pKJafHMIfjAmiQuHrJqbQCX7YPy
AJiKom9nI4sgcgvW4NjHZx2s8/LHtW6bCaksCcCtVoxynj1t1D9sJ7uy4tg6
3dYLz0L94sanKpBK12iOgNQ4utSeV2bw4RoR0mqH5imXbapcvbKJmlg5lmjm
85vrDBzXakxVUX19M+twKd1576v1mN5Og8WiqMtIm99W7hKiqbS49IDvLHuc
VzuPR8FYreotAhMp8NjGEZBy3XylAnA4C+QU+fa9vpfmxIALKTF4Bn/Rrh/s
p/GPeD9kWX1s64dJ+sBa+09mta6uEb6fC4ieHvWXRuEJtlwSLDBxAG135mgd
G15J2f7Xl63z6BtBwC3HLo3flPFL7XEqwCl4T2+0v3GEQX3pFZmf+ed5sFAa
fBC1NyXnpsT568ZffdN63Vb14v79bC2OTyN5uVbfN4FCSsfPxJiEXc6jYoqU
Dy/xMpLWmoNTgERCoDZiWMhR6+HZ+5TcjHtJphRHTcx2JCsAOucTBbKA77MS
wQvU58kEINlQIsvWa7F/Ra/BMTnxO01PlZVwF1LGjyVb3qW7M8gPHXzn7Gqt
gT8i7tK62h4qjfAC/LQcs54JF1burJoVqhh9t1as+OOogNeFkDfnzZN7n1g2
kSqhrnrT2Ai4wnKRY0sYyz0LxdWhNbOZZ977RNd0jyl9Yd5aVQXnJtJaY4t4
Fwr9ByN4vztQpNh6KK2dffWWL3JtpGtLXwZ+5iW8nkYvFtivBk6ePIxxNJvo
NrtqSZY7KVl5jQtuEn8MyNN8BV7qfp9NghH+1wETMqxR9ZgGRBvtaFO1GImY
lKovqkdl1qJJHP/6M3Pn6Ei42FpjPx6VL/B1OMdyPf0NnwsYYJ8DM8NUe/+w
wyNkpQmZDZxPXaVRv20/chB9223pyAtYRlVQ0uEfU5DgtpcEHi2xJq0qWjUy
HyKOl7HKN5ue8/2buRqSM9Eb2ZYhy0J/KiKDawN7PnacrTJb1XIlE8G4hw92
T56k6ZnASh/Q2d/TuP0SAmDFIpSrqPCxdli3Q4fttd3y9xQMIO5atN7Y0TA9
6XGSG8InLKYFbRK7Wb5NAhmLyTuLheTlQUJGHCIn4JnbIY1i4PrySv7gVV8y
eeUwC6lkf8Ufry8ieVgX2xNxsdFIqj92Pnh6zuBnffoeABxR1WAZSCE6wK7g
8VX7pP9w2qhguPV/K6X86tE5yS/t9u+zIiBVKja6WLASkgl958GLoHStfbif
8BJGQ60dy7fgQGoJ/eoQWZ7H2cY9rEPKtbtjGWkau8OXpT6XEaui1Gv91A5W
ZPWyo75XKpWIr7AQggxT7CQZ0F0LqlPjOLDM4EVYBqUkHcA3+edjyXXLapn1
s2thfWarMl4XPPTSD4hM8Id7ASd4AI+xUAQ8lOmqGE2MmFZDCbYUZPoy8/4g
lZE+E4PcuhbEk//2V1O7scPMbWkvKw2rCf2/0xtn1FxQpD1wNrbCsfAK2S0y
uRA0Mm44z4z0C+xCoXmb0IGUagmU0Y/qzDAbK+DUa9YMq85lSNQFzViRDrzm
oeVA9XY+l7sY9NsGNxNQvy6VSoTHvaqJEOoD310BxGICKcInyf1d6CJcJrfE
FTbHcuvRj7N4XZCnVmdyBSrB5F6ms5UUp+pyJf6CILD3+4gfbXSDmIW++qqJ
TwGuBHv27ZeQf/7wg/RmTwjyp7PAqJ/2KzbBAoel6YhE/uyaGwLZa5CPnw2Q
xhKHVPNBT8JEwb/T2BN9+l2bsgdj/+kBt6OI+lbvO7VI+BKqblp07WD7Hh6v
L27jvLblEw9KhwQxznC068JM6E76TCDNog9FVUHX+Q3r8PmsA6PpwrHjmRuP
2OdZ2STRaTvy6wPUmfOitg2mX+/hnFIFA3Iv1jsNPclLZFLzMYCWM1o68zGx
UNPnxLB4CbIkFtFrVStbLjQ+G7JRvob3cSyCoeY/otGVZzrZWbQGjNfQ/HQP
IQJB5WmQ1oE/R69r9GlqrKRoPNBlfOLRfa0uNZi6XEXaQ1j0wamda9yfuIUv
PnujhZvusLT+ppvlseBPZntDGxDlsKaA47s68NEiTtB51BEtJY+QHpfrp9R2
xF7OC1J9E9KFXyYmlhhaTCrbE4OZPrmRcKr8L1zzcA4ct6KBePHv6DGofEhM
9B/dIp2FmU4TH1VlzSZbpK+RZii274wGbut5qB4KvthNmXxV9pF9agM1Wwxi
fMT+iYb8kLC4y7kcq3Ob5JcF8LoaXtGwG8s1RlQqOVYiHT0QpQsgDrqPGS8A
R+iMKIONuOF1RrfBvSubCqlny74/ajvigGPvXtjpneAVENK+bZw6PgVgjUZm
1Ge4mkhZjA8+piCXjyL4IKJEphBsOZgx1/jROTU0UlS4RgzSs25jxVJkcaS7
x7XO39CNOufhTXtdGyF2d/Ujkjl0FoVneHeL0+7trCuMfCBc4KSF5+MD0Eix
JJHPITcqikU5PJwBmCx8gviZtgR+7WCmyrFJO2z2nO9bcOufSd+TXOe9ugEf
MX6zpbxNj0iYt65Ud+POXplugnmd+m5hB0/HPw97/r4GY2eh2t8Q+dvOl1m3
HyT3hoM5z7ZplkMqYTAswfqyrpz/PTpBjYpSfiCGgGdD6LctKdOHkD63ZiFr
L2CebEGnWcDUQ4RAoECebwFVsv75gL8GkovLUuCJ/rtb/rr8VaPIIDEnqCT9
4L5wKLis4nAkZ7BVhcxGiCo9DtwRPppwErgSWQcTR6GKdLYEWPHDadHKGVYE
VN2dsNBTdkrvecHVaOFUZAdkhpsYwCMOhhfQKpWqtT/idpgPIXmnDogZBR8k
iJys+EEXwLNNoVKJ96ZJL/rcOkv6elfwBkhU2EisRgLPH9WTwjn75ijAYFUk
Cf0CUTMimg16IotoU6xYGssi77jTfoCtR7BWDGvphoHg5+/3C4LsgJIlj2mz
hU1AHB8OE2ErEqL62c6q3VfnAMrFj3Grr2MHtEce9WOC1fmEkYwKRZJX2AQU
Zz+nvpEyQOF3AvDLmlC239sMP8fhD1quXSljZUfZyDzUaICtTWhJKxL4CC+a
VxAAh8EdUtN8npHPnuDLzT4fSQpXk58UQ1CDrSeYUgc0XdXC7pXs3ey0FbpU
RkUtuCB6I5+uXsZxur+WdnB+hWTaOAphMXnqgXt7Rl5yGGjs/SxLOTTprOlN
pkzwNBVdLK5l/5b0U+rL4q2/uPSbizPSuedglCd8F+p/MjpELiEJj6i9S3dr
mJ5/xLKMHJYwB0370Y0dCra3SX+9/C5s1LAt6NMa8vhSmgccsmQBicpM6+iM
iZkuRytL3chJBtRGIZolJddlduOyHwTt0MLGnjcA7+Fsm6kHhKHMSmKiEw44
Fp/E8KBAOCFMLb6yjh61Zpl9HO2WIqdJ9LbCMS/PzNe1pWUBU8U80WI3KYnc
Pac0WvRGl8QSJe0ASJwA+lid+5jcfiSspvuQrvKlkvuIDddWBtuV+G81BgS2
QFFUBcmS1AcKiSVaLUDaaTNQjLi197tPTVGdJm8yPTs0IVdZMV0MP7pCICdc
HTqPXhyjCw+DTrvtFyFgVxytodltECCsE1chuHskEanIjgXftH/CwJKLBSyq
hhj8ZoKXvYr9+hXNcx5NluRDN39RaiqoWWV1tftlYaAuZYoIm7JcdP1kcKv4
70NI9rrA40DU4lEXlAsqTWCfd1DvP29WJQsJceqaa6Qv1n4Q0r13r82hzmXL
sa86290lkmj2fT3LGDb9K5vi3OCcf+bxj/Pv6IovvNxgByMEvq70wUajiqHG
A4X6ki8OKR4WdMFl9/hbgEPpscMh8HgWqaUZ4tCdEPSjHvU3TYqZLIfS7RCE
fdeHATZnE/YfeDPBQWTxTZvA1jec4NagtYuF44+lV7t4GTv4JwXymuuXyztg
8i2IECsOk/YKmtnDPZ6oV5eVCvZwGPgEEU1axkXX3X8Csik1uovH9BPnwDgh
u/6yqlZCj5IltqVFPb5GhoJI0mh3wYStdrzBvc1nlVctEb4Vx9eU4qF/NglG
dEer4Hx5erdMwrzGmKk4eCi4bU9Jt9CIPbM1JF0cAlLOb/xHwNZjuN2ldXYU
FcQTP3+gcOEmE5yhfyJCF+i/+huwBswvtzd2G6CDasx94urDrFsSWgeab0p2
i7d3AhBX+DUwT68FVpoKzptL/982oNeDz11ngsN8vQybVJjC1pL/dpjC20uM
FJSxNHT1w1o1BeL7GbVphrE2L6HRuwTtRepA/IvfgjiG+A/aw5SgFSOu6Vek
3Djm5ruiXYn5V81Zvn9TvI9HG6VpgWUaRRLRNWnXev0koof7IhKc0v7Zb3m2
7cK9kYVK3F/Mcaer00zcOg2PgTRCbYGU+U+tx8d48UuvmFQZyV+6PI6FwVPr
1cOsSQoN7eGadSJSvI6ve+4wKPiJ8O3FE4mIzai0ljOMpyIxU7OyivfYIw4D
P3oLSKJ9JSU681hTHCvSHp7NNM3YydHNlZama1ry4NWpz2ueZwd/dPKx5QYd
W/37tzjE0cWq6mQNTnBMFjjqljxDtzTYXqEPUtbLrX3/uqTibGey3wP36vxl
FrvM6c8I/jGQt8Le8AALmiRkg0HnyHEd0aG3QVKX2LPuDer22f3gE4PPfBnO
Z5v1/9DAuc7HhAljeRF42nC1H+E51sQzu2kDsdoEBoxytCsgzquLOpQS14bv
+TdEhXoHZvutl6zbiBzad6SctJHfCRF4wr4XByfqkIS9DEQD6/DD49yHhNx3
U0fnWVkfLRXJQTSQtCjnUx8rOj4QM6iuFbqEbY1jweJ4lpy1kq2OA2ak1uum
ThfNXEccvEXha0uwWT1JkldcRWywwCb3qxj/JB8rflDRwUUawOQ1elUHSEV3
gBJ2n7ZWDcN6dBSyH+IMXnaRPWSg22LutYGRiCjciXmkAMmIZzzbUzjw4pUc
rMAwAkhsUqErTaO0hAdtUsyM1VSA8xpN/ywQkFLksDKiaMjrxZRngIEydKhU
9lP3JnJGE/RcakzGCpMfpBeBbc6xZU47C2TJ8W/ZVAY8AFoom8JTvQs509XE
tVR0/jumX0+6WlkgV9A2F16DagsJH2bU7hNVFIqZn20vlaXatU0IENmdHJd0
DZvplars7xyYam1WVJFvM34JY0jBkI6Z4kTu0lpgkfOtjF7BCgkTcrAr277z
GW7mzY6GheeCVIMEDdsGcAnlYU+FNcQT3X6c2TyCBRBhbpHt5G+lpobr+ec5
baTfy5zC9UcwZWyT+4sDM4GxeMHwwYdHNhDoQrlD/Q3SWF79kguOHH8NoEGP
RxpE6i8SqHNcuZyNKTAaQ9u5HP8E14L0StG/jH8ju1EsgKpYZMD4b25E0YEZ
avaUX5GrNJlDiqE0WVklXI6ZGjlcn+Tyu3lFXiU+VglNNRVrsrBiZ+9sQa1M
N0Kj4cxr90l/2cbGfWrC7cOkPfVUeHgz5sBwX8OyzbKfBQz9tWix0FCVpZf3
Sg/8tiiN+jzJMJW7uWkXq/R5HmQ02Wmo4ZuMLzg6skYH0nyGJAntRuuDEM3G
QRzzsZKy3Tta6ZKHe09SKGAuPxnPq6uf68CguU5bd/GwWH44vrpgeQo+0sUv
b7ySLhFedIDrgpYADtKWCeaS/YclrBtlRDLLdJDe9/5GYVOmAAwxyls7LFxI
IDp/sgrDGd2tF5W15oQUgAZmCsOuZAJWuvYPcAYE2F1ATzmxKheazB5mnblS
4iFOwMsPSKtAmixwn3y/a4OG2O0XW8edrwyGNlUDCIeS3tRXdc4KLq2waRke
g/TIsisLtOlTkcBNo3BPd91fxVoLTmuepo780baJ9VFEj57f6YNbF7nmx0kv
naJs68lknckyNJGAji32zAlYOf52Y1l4J3a0h1CqhQlpZBqeykzsjcTInsWR
vkNvZyGGIyh3F7zI4+mP3oMmG9C2dLegguPgiUdW1ZqUmL7B85Dz8l8LmpVB
taqK1SxhHDmCSJQGWO+mDva47rrVJKB78KiDyxiuTwZeilZIRPXjoz1F70Ea
/DpGZzoJmWSjSnyIjDrx0wo5ubiI7xdvk7fIM/B+WvFHWT5fQrqYR+Ms8XJC
cRM6UmjaS8voNdcmzo4FVt7bEOVVoJwqEnOxdi3m4iEeyoERwnGU7xSkH5O+
h3Br8A6R+jxbk5IP5RDUNeNrD8FP7cDB+l/CaL9T/F2fZw4VGlzr/SnhWFw6
xQEZE3CU49tf4L3LdwORNqovFcJ8EHiNdVxVNuNAXb431udey7Gm1/i7jR0F
l+YjWJxtCJGPhWONcHoXX5258ouIIu2Rw4EiI3VGYkvFXJmJ2EpPAfkfcbAo
zmJQFAXHjKTVdtb2y6uN9zXRD/fAK83QxofItByLAUxJ6/BoI0ZDdDvHR3TB
5rk7fVodwaY9Jaj9i7TBsWhzRsgRzbgiVYPqe0B4fMWrpDZmrN89u/R+xZlD
3pIE58zjkj8Z8ixWrFL7ywz7a8hLnyvt4UqSQ4rYmaoK/9fVm2eK/3549SYi
Th1hs+5imzmP1x2f3aA4uk/MhPdEITphdU60V1M0jGis0r+VDdqAUxv9HC2B
zDTGkA/3Ys3kgs4mSPTuPRfdXk5O6xau8MmG1RVdnE9mOi9BPIKudljH+4o8
YJDlgZv5D26Z7LCdsw0EvwgS64jLTMKdyKK8GlJHPKB2vK4FeYNsWukauKnt
zqLI1IJjRb1axCIwM0iYN/MPv3avnIpKFrqcAYhaQKN2bU+uWRy5AoM+2YBR
QlOKcDFyxLUynUyGZAk4d9z27xm0KRW81fluE/wPg9IF1SWcjsaPohDWcmwu
xtxWLR7TBehP7IvIJquMYNjeiyUUeo+X07hnIFZDCj77I1JRYQEW1l8sQGDz
DtesDQgI7grZNnIMfmGKS/N4sekOCYw35xKpoYbKBf5NGV2Ksn0sJvkPXYK/
7Km5cyyYci1vFMRTIAosO3mJKTpZWyMtheTcxwzEp+/D46oUPZ94bek5MaNj
cLxcbMYfDHcs/FqZG32s19OF//HaqvZ7nNwgGsbYq2/cLalhKXrUZFaX6vMM
TXIBWsvnzhykvRx5qTpX0rPqQOj36ce3X16mZC8N8fXWD2uBG44kvNX7XVq9
/Yj/t6rz1X9iJ0EPrj+wQ9/xlEup9KYpr4748dKGe5PY1i1Z9tXFzMSGOKmv
VUX8aBL83rrRcdAwJmEnbY3hHD0QC/SKyehyKt6zBfW5rXSgecFDUVSPpxdU
nvCQxAeyyBb6NEl2co9JZhJZ8BkZGVnPMJJ97hIJaED8X7OT9rrvmnIEv1Qr
DW9bWPLZXIoQ4ywnU/XHoYbAsMwTBy0Z3r62cw435zPbxOY/4Yg6/KhWMlvI
sh/ghUUVn8kenqQGLjAN/UsnIXhPQe3euDUYCj4HF69qDNNRyfMnXFA1CV6V
pmvhDwktMP136jIQKcQlsW3HX2ZNOV6OCnLLMYYcNtPGt4nhaPrNBW6teh4Q
cZj85cRRImXZBbB6xvMCp0r81HOmiIPpAvkVGTHNPPICCDstobyVQU2coDF0
Wy0CCFTozNC/TH1Ft+Xs5vrxz4HG5RTsTDQN6u5kTjCz7guWs3w4S8+mUnA5
QdXHcCp0j6P+FC1eRBbNBTYeAsPNClUN6jlK//Hg2AJlNeSXAgJBOb7+OALN
7P8iN83lBdgHl8h6H9elCwx5w9aQkCZjWO//Vv0lDmrZXCc8eavcNtKwI2e7
UP8edI31Yct/Qh/8rT29Q6PukL0sw8koQoE2h1YjVlLv4mUqJEt5jAC2xC9H
j1E4axmAkbKjFhfcpixLg274PfqUfga5YoAZwn27abHjJRpWTgVatXnVltB4
svCpaPRyJztkj51wtM1btY9qQ7dEaWWWFuoy7hdMRwoqofsGAPY2qV4rGriJ
E8RT+mnpYecLTMk3aJB5HaTAaRJIC4WdkLOh49kk8gtfK6fHuegLwIIWQpkm
nlPWR8ai6V42YetgU6oZ8O4NJjDVUkxm9cKE/LrDybNsVmrkOqxOcvX551JM
46Rk5Bg+iMpaVdXA8rHyHzeDWje7cHzoExNA6aQazNG42fmZk0xHowid5IG9
BsVm8HuyY0oOogdzS5Zspu/uU9urniT8HppQenGTa2o+1AgaYOh4dY8M8m/E
rSJBJysuA8w6cgAXNGU8FTWWeiw8d3+1KLw8GQMMwqqjXChDwYpWJ8K2a6/8
fLC7+p3HPjleNEfax85yJSlP1hYWsVKNUmQV85hkPkGrWZnoPqgD8CQLcWHY
JmZypRbXAzXBdrCQU7sddxpNomvBpOyMBXayOwZvx8l/GCcYGhbqVJy2TbG5
FUh2iJJBM3hJ/mC+sfYJgm9Vbo56obh/oyteA+lmssN9TKCA0+mzqRsd866Y
J9jm4SGFI55iKZ0iiWc51cQ18ORTZHOJqFXL6InoIQHSA1mYXm9X7sPeie0o
6gyAC28qIf6E786siNyOCWqpgpO/NjAFrc+p63iFosT69OIyT1Q2lUJMfLpP
CsbKBSVP8lpu2UYYBO9jKUvF2kiEaihtdBnQLJwOw6rnSxVfo1OsfjAZ64F5
Z4W6/sWn2g9aMO5KUEroxLy9RkmfU2sOqP3GznVLfDBQlYyLNICNxF93hdqJ
Dcu/327K8p6WyoaFwZ5BiI3Bo0kcRiV07cJdbA+mtPnugKHM0XHT64lRf9hE
7jfzzJd6qYmOSWRBjsQkgb4CibpNOHZj8hGuhclcecE6KjjU4sOB1a6hOJHN
s2OQusDK01W60Ko3qow5l1Q6pZ4nfClC0deV0+RghTp48kIrw0b7SKDR+ADu
xN2WzhFPK1OKjA0ijiBFHsO8h5ECUgo+RJqPlaZbG8LBmk83BDETzZzDpgUe
ZclkNAEZsv2sF4a9+O/JzEcZkKHUft4YQDqV1AN1AxWetZVyljjyE9mYsVJ6
1ER9bdgNA6LJxlywBAMAWkgD8UNqZmx7rPvSLiDMjMWO5RlzIfl6mSFuxZ/7
GKGDtMjnsIl9ye/bgBeNDwVh+QkEA0syFADktdHXD6J7/aUnu4yOzTHsMZ4j
oOkdGozvH+7y3OxfeFVv7hmv9MaUQuMJsx1zN86C7l+Qn8ZLzd1PKIhm1aGQ
4546WAZGLD98lMN1Ujs8UCJzdw20RdA76UIfvD/WRm01YWqa4Sv5j5lP7yVO
4WbQa9dr5YY5Afs74W13YrbyokIfSGXDBGuiBAxAqFABEW9MvovxbOFKhzT8
UKawiFKbHlOOINS5IeZXNiML+cUAsjP6+hQg9qmHyCnY0ftzFOVuDh1+CK8d
1hv9Jmwh58Z2XAAZYsfIEUBY6WdIdUVw0Rx3P83GBMRC8aShbOl5P1Q8rXnC
+jBKMjmr72TeetScRHiyJlKeJ9gzaqPRNCZkRRAR+pRFcYoUcJWLzLY5bXiC
wRQMRjzngodS0kx+AJN2UaZ9HHS0ttanmUjwCnwhUaMN1Fx87LuqD2wYiMOz
PZxLZyaUy4RwUPD0glBM50h7+FpNJmjb/uShc5JxbiUma4azoz+n8XOtSX6t
dtr2nibkfBLk90fy0s+mTKHN90t6UuaBsZJf+I6ezsiiGzIHMMU63gs2uafx
za9Ya5Vsugz8slEEMselX3j+c/DAi0/MC9zr3icUNe/8uAyd9dot1jteDo1X
8dUNN0Kwuq6UhQkYDU/5zc2+QB97Aw9anYxExOV/IylJWGAvENvTVDLgftZW
OAGQOOyFA97ZtcdBvdxJZ7qaruqo4gmLzyMILhyJ74sBIXDtUWm7bRoE/KZL
uo9r2MqnkprLPv8xCa+awett33Y5wSaSvVFjNqR10292fA6H5lLF1A6KENOU
SwGPqbiDTNO0J/JPgtEHy8294nS6nLxWaKlJJYbdijYfiZPWJrQ+S56iQFWa
/TwfmPza17hj0c8zycSySdTVAJrLSD0VZE6IH5rMp/RvGCxHLzjmrHXwN1zu
i01WWBSqh4PU1AOKie3x+W2Cv7k6o362Ktii9VJRz2pQ/ZfYzvKP7CmjfNT/
XxntsGiXcDSaVdKimGShZUdNidh9FC0Smw5wAM7tvIsHDv3hUPihrz/dsrH5
n4q0NIJxMUGRJspqDV5K/d6yWLeyGL1Wvz4LT/IybnzMU3+K5LbG77DL4Wdg
rESQRazjJsSVvE/ig7+BDMb4mMOuJJbrCf2mKl1dg3It+6jWyFUiZn5JFEkh
KycbKRFWCOa29X58nB7t9XjOlV3Yx5NBzkM43iOqco+eYuJpbKCEgZmgg8BY
BYQimzc4Z7F+kkHUpcr1uHbgo2SCxiw8BzO+kDLSXUOsO4adT60konDrEWe5
kUngPxTInZ06GhOxxbtIZH8oyOyvEUKC8DQ8FjqArxxas5BYr5Xofn9l6F5K
dcnwdSUr2cyaPPaPQQMcMy98no9mUziIzImbR2P2lrLxj/E9fhqgQ/zVByD/
GpPn0DY5d7LwqSzuekT5k5voqYQEuFZ5BXIZMejiHptXpVhy085TjOhmeaaV
JoRZfC5X88sh40mtGzrlWkxCCsp4rHkQ/DPq0yg5s8LOUCBHXNj9xoYjhF7V
YmfdeplMveTZSDdWTwVsAj3SpIQFSwYlKg/ghDKAQ0VUhMO7QHOZsJjkWqxZ
29oKmA2gtvaHnXbb5sXGIXpR42JI4X0Zuz6d3MCUnBZLvHZKNlD7JLgoAFbM
jOX1CcC10ZHfWiJewSUhiJ9tsJ6RpVWBTe9encsQZfUCt5GlupI2SSs3GELX
yjlsGZCZY6LUfJyTfS/ITgn+5VYMtBidA3bPb2DdOqN2t/mTJ/tXm3eGx0vW
uInYAsgj/gX4jmhDGvVKdzIcoA/2vxg+SSwI3SJ/K64ExYv4yXUcd9jceDTN
5ElleOnrV67OwyRq7vxTlV6kFLSUNIDMr1MCsztvQHzed7RtyeyYthEk99dv
bYHGdUxJYlgyKpqJosLYvoWGy/VoYBdr6Jq3tmzNyOykymeTMhNaz2EqDkvk
bpPfq1cp5s32R/Wd9E0BusyN+NpSgY2X8xJr8zOXUdFHQog4chnSviRn3QnF
EEUvMkpH9+ZiOgk2PACzRwjRGUBnF+ygNtsStb65++tUt2t8SHtbOzDwt0l1
xk3bwPL63RjmFjwMjKeeJ206/IF1YvQcU2yLwA2ndtzVPrh/kWPej0A9Dixr
C0LtcNDIhkAIJcx4u1LJzwEF4xH1IvAhEzk/eElw6AujjSiSC4OEhgP+1jWY
FAsK9UdheiAEi8hIIOuuY57wMOzUSBzZHhCiTcPoyqT2LH2t03A3rJd7V7eN
VBgdhx0FhJGzJNNIdFqHeB6GA8aTstySzv50E1H80iZ8GhG8Skdur/KDKr84
hWdjcPrZSgl0iFcvy/lMO/tVY5LaKQCyJ0sglBA9iQDn6IySu8OrcaLThgX9
Amj6os1CEgZ6w3HtdzAhv+AE6VhYuzRw2YSM2+7XRMD24BzuPbv3qU/fCKL/
zGkfPpWl0jDfc9Eyu1uSwtZtQQ7iduBV2iqvmYoAozBbvUmIqZqoKF2AN1Lb
JTY+EtBESepb0O59UCmekXXt/zP9Uo3RCIhxCxGrvJmHbzHG6Eu+wRpAXvbw
SdqjltV6cVAl7tz9+eSe9EnL2WPVBiLQwcCaVhpdydxwtBC9Hgfwh6lUnqLu
NDAbitmbHPgATPwxD0CzZQnpIZjboqh3VclCHN606wnahVW/ozYK3LZdBZxo
c48mENJ2HL1+J+58dFP4Liooj0hOK4o52rj9OY/N7ubQ5BpPmK5ShdqfKjDS
k0jDFtWj2N1hG73lv7Ps+uITC5kKBFYHb161H6uUMKcPHECLDF+vk7aZmXVP
pWuHeT28A3061Fe/+eJvJkqNkLoMJj0pi81M3GbrAbPQIZj/CfH8oG2vhpCG
gBKq5aBGUbu1wW8y/I/LVzej/+MX+PqpFvNDYyrPWkYIlh5NxHlBQqS3E3PH
tTl8gwkag+QgxNqJLfYCCkNeLyjEXaFDpuIwj6lIflxxiMvMhiSv9i90uJOk
RUWUhZolsoViMqGwP7RlBRLeX9PfiDdF+Csy8KbhxHpOXlA4eRF1sSwGlMSo
l4AGEeQ3stiB7qigZLWbboa5ah0uEDWYHGPmisEs3rkC5gntF1i84nmvpkpi
g9XpwH6800oxXmO2/9wihPrvMTKiLEGxCaaDLrcuPfugJbm6y61yEpUZBzrY
hzMQ8PdawRSrJHNWUjU32DJBUBq8F+/Pk/uNY3HIq46wBmhotH5cptUKVW+S
aStRANf7pcTKp+YlGIuAo/mEvHtw08KQoTqj9XvXoXBOyU8ZwJOE/GZeu9TT
SZiSP5/9QlFpxRpIBGtIpVvyQOAHVpvErs8uecHWZeBz9Oys1thcVD+WL6Og
U0yDBFgFwHl16GfBI+RjtIZ6Q24Z+tNd7oirCtTHtsTIdrC+0iNqMoc2SrRo
sEnDk/NmomAe/Qk6VkuKTxNcBaxNpwKdrzsZEgj3NBxb0S/lDEq+pH2IUlc/
5a7lngjjScoqJ41PnKOOYxFjW9hpkgiK5FX7u1Wy0olfvW4FfJmcQs/Ofdox
M8El2SSV68QUaVVAupDE6uRJU7HvEenaNytl7Q2a3NLuFvoLdzj9t/ZuoMzo
4JL4w2X70uQ8a7zfMIJfeom9lMQFt8vmo1yeoqO/nY4WWSojgiSstS8oK4qI
O6DE4LqXBi1TM3HbYrywfLVroU1tnlWn6Pwcd1GSipEBfNBMYpioYJsBuT0/
NksL3IIn4u/4xM+nf1Lk3EiQLTTUEPrgW8HtoMX72Uhvf/DrOOVE2k2VNe94
xIvshYgrJaJWjAv8K3LoNiyUdCb4+aPOZgP38QbuBXr+I26cFfPU4P3wd0VB
kPvYGlEEls7LD+CAKwERT6F+66euQn05mjbWGENXe+77kbACCFLoEKKhCXiP
lL1XwEWV2cRD74IE8CysdmVseG38KfyK8nYAvVP9uDdyaiKSAvZpHHHUJ6hR
iyL1bKC0Ydqg5RVIKq2m7hLI1W68vPJdAkE+g2Eux1nzgBm7AlYl1nI06Joi
Be+Up3q5R9o8sAFm2LhH1LihBXtqBmiB1c32Sj52UoiKSEKOHPwa2b4dl80/
mxoyQlDCVRX2K4IePdrn7fQWo/2KNxepGlFQuMt4HF0aUWhF7jNBA54JsIRg
sdijpmTOIv5srQxMxeZ7i3YURxciY57wPLiN4bI70aY+cUvmEqFEUldpIzEP
kinFsvCL4X77Nuke7XokfRSz4M9KxTjiratESwCwtfPWavljcag6CC08b+Cd
8ygl8yietgNhhuHg7OYKF1L7GTC1Als/wVvcIwNEHjrQKwPtuI5orzG5EVyn
WBJYx2/P9Qq2oRvjzisBx8HIKv35RDUaTjm+O+EtHzFkFk3klt+x3U7ATq8/
vznUHD22MG2zawoA/k7QYV2xKWvrfdnpq2caFul9YiEC43IDrfahjSRlJq/V
hfubRylRfDOTg2vd1edVT8rovv8c9Y4yrcO1W01Z5GL7TLuyVzkw+lOlKzKS
/1GnLYSnQus4O/hQ+g7WSE34Zfy03PL+tyT/id7Q2B8iScDmA450xAy2kOfH
4rG0nbFsgNxGvAcl6n6aQLcH4Zo02+54kmcK6FNRjJ1+6M4ffJcIfyenLZvJ
Vu9GHAYn3z7F8X4tbFRCy2YnI4sNj7hlaH30eoRE23121//CBKIWxZRfxIwl
EbXpiWhp11hfmgCJaNExLvEUUom7whRkW2cFG+qOhCXt35EAq1+lmc3/zRm5
de0W6y119YvVAy3Y72jx5fngO5skVfrtQjHnl8h1Gfrpao3efi/edhgDv4J2
1UGBA9Ivuu+zOqfI7lfZNA5R99PIotTYklS/egSNzLGUU1usgqaW8lY1eZww
7AglmZneRmZKndglBQV9GkJDIA1OKBzpqromf3NwAmzOvmSPk6upF6eMDlg8
hi3mGoJK7AX9S3Y3eiL3Te44UyOZcuq5hp7RtNwKPf/RnBIulglv8Gkm8Mk9
fvL3/KXYJO7t+0VFlpHSN9O3Ww8tHJ7czVljnHatetnViy10nhb6VgX7KU8d
1UL3xtuAoVBC+5mPp77Jc4xOP9NLFL3/NlNmhTJ+alqqNdD+eRNn+o5KQcyh
bfTDjCgtk1J8v+3HaXy1DnHwntef/YtrQ+9oWURgZC3sakP6ehVFbx8IdRAY
mG816zIxE+dTwCYeFrrQd3OOwqOGLhZTqn/qAlmOGsO8nsGbCBfT/xXmWouW
90dehDWVfJVswrIoVN0rw86tRwymEEYS1CRUKn1oQzFtM+PBGesPNgzO114y
zHcV5gZ6iCTyifE5VwiwY5q31T9uInV/1GbPc6m60+9gyerDiln/NQWz5Co+
WxcUnr/Vii0VITRnle1csyv2OSXHW3uVZKPP5ksSZhmONeDYvyTJEINFDOJc
2h3brmePs8AnuZM+9JXE6WOcRDxEZuXvIpLtnINQ3vAnrIJ3KTCoxdGQUWIg
djg+TL61p3L4FQFiSLu0nu9lZ+35BKfCvpY8lOrXRTW5DPqycA4SkvPyNy4Y
7M86mncAwbQYNQouT2E8KPLMYHNaJRs7C7UbBEaQs5BgbLwDUdm6PicOd0nn
AmgQEI0YWQ+f9kpPUsbFlN13TuWgV3PQvnkjHGe9mCE2XlRbhJXw5st3viVS
iRZUyZpwMU8IOXHujDl1MFPNgTXhKoKmQZitHBxTbenErtpNSScnM4/TMOz4
gsVSWcrshNh5AMXcjJHu0/6rWJ5YvHwtESrsVWcgAW4G1PM/ashFhfpiPqwY
rTyNcV/wEGjOeqL1EoLNoipzmDwGKsQLr5+3HgBwm8C4Hcp+Wpn2T2pTenNa
FVTn9KDM+NDMVvJQLoEEGP7j0tUk50JttcUX+STAVfu4weucyTvpJ2mDcDYo
bhx3szQLJJZGajyoq/C2q1YCnbPwo0B4bBr2q7Q1wEFBcZ0U0IQBJ+giEcVk
mVOrzWovhKHt38KQs2cFAft07uz3UwkpquivZPE8wPHeuhC141GuMMmIOTLa
AqCsWCpiVP9jyLUeAVw1cWQes18qUkgBI/NSwQnT1QdUYk6M8y6smOq6Ljsu
AfGx61v7IUukJaVWduEAEuAC1kTmhgHDfbWIsBa8zXJ35t+IAr8GDWuH4iN5
BbiBNPwn4qkbit8ZyALMthb2iLlTXxHHtO9FEdML1TKUKCG/6sVfQiFMKMtL
qCwtmxc63Ax20RDHLk72j+YkIgUuhaRm71LfksvusPGlI5cRatSQ1vFWlXBk
OfjEqUTbekoTzVKxVt7SksDrY1cxyjiTxSFvl4GE8ILjMGIyoYwfy5cADYb3
znIuUpLEdaretgIkoBGajXCHzUlfa+3LuukRXxqMKHRC0xx1n0oTJ2TAlrCv
zXVJ9swE3NpPKIaiKroUgV7VgZc5t+FWhyo7sgl3mLbHJZNzMGIBo2xLYZcw
lGffX/RDz4HddRjvnArmL2/KigHQmiLxsCdgPn1py/GCznTuCsTIpkyJO5ru
4b+GGqrDrb1dSh6l8a8VA6fQanHuPEtWd+grA2IY/nNQpILOJ8YA65uovfhp
H4Daj4kmZw2XYdzXdQdbLRffVt8iUloh0i1Tv1nv3jc1sEKRN0rMAz61w1Ni
xvidmxTuc9AzP9r0heWlqy6JlOKlm0oUMfWPXbz6yMQGVCJmfQgnXATaliFc
gTknElcp2KswBsFOQK4sdklTZj0t9sHGCZ9Mak2CrvijiWTpRdwzeswYO1mc
fKcTYxq4GwNgp5cfI/BaAdf1lJleR7DYMp+F2h+iz8z0of17s/JJZILQjvnK
gpR0tWQXNaA9zM7qcF+ncLNff1QtxIJSIl40rl+biXOKc5WhsgfUZmEjw42O
mAEt8pRcjeKUQwdwSnh73vCTLtpxJ9v1QXhrpZ6eLgGW6zKfl/x0J9OAcV5W
rh9MgZBf+nGuU9RmFw+6TeLoveAqNTC0I6PL5d4rwdCDLXXJI3JafeS0uD36
86ukwV3ERj6QM/etTIr0Uo3FJmKvr5HLanMQFVBBhMJUwwVvCXhSQP1lo4QI
HPzRjsD3+6uWU9JtTDmryBihevqzzmzr4P1TXa/k1zo4wRi03dzM5vT30zQ/
iblNWX5r6GCDWcKvLmQcnabzPWsn08qwztCDY5HfE9Tvjc4sSqaeDV74s5bT
8BQtzmkSOIH6IXuJXnAWtkdwMVKkuvBai5wIeuEckc8VhD6/iincaZx3Ku+R
jRHXjbvUmIQDt2KqPgDKSOlIzcQgHfCQ9LczZapyLd2Ll/lbi3t4Zh9ZLvO7
TEfNKtqfMMSSKUT3F4mWwEAUhIAUbfnRxTlcZhmbvbB8LWjUIl1j0Nf8f4KR
ITph0bnex3CSE7830UbOFr69WrgmplNzTAPcAQ0X1lV81uU/oS4RiJtAhruW
+XCfNA/VpDZP0oaRtUAcLJeMCjlN2ZkiLivC1goOXJ5LQwzBw2NzZS5BCaOZ
DTOmrcuuZ05WPeYVFqZTZXpjobf+dczoHHwD9AAFONPYfPykoVkeDIB5BxaO
4H4+Ojz2NmjknSlnH5HSMNoMxHmFmjklJeJvcHgrP2yDRn55B3cyKD1o2goX
ZlN/ZdvA6n1SkObnTXO8x+cytX7mwkFKByfPrxDNVQ8i3EBUUe9e/MJy1IY1
KcTYhZHSelu37TDzf4XqHCAmOFipghG8OjSoo+w9BB9vAJhWt1Nubp/b1mnb
W975DKQSzVGCnt2xGNhF8MKYUBt6hwbhQt+lqblJw1OjkJlbIABQh7H8qnur
qqKWclGVQaeYyrfK00hA2ytC6f6oRxT54T8MLVI9XnMnjhrY6jY2sPxth2Ic
n66ZT9n8NtvXMdY8ChdcsWg6Hpa/WM08n6Dz/MkpslnOAEEMky3GYp6EIAyS
72GmMV8z1PEB4OZNTwg5XZVFJ8YQRIXwTqEvHHg4Mb9dAGJJ1+GLvKUqOudr
LkF1ddQq6qj28qAx7s0rMnyzbk2xK/pbEgydye0hGNimPh695iHf2jRpbLZf
IX7/1SCExoEMVzEci67wWWE3kXY+dc729VzUScI6gCbl3tDDMqm7SSwvIFFz
ooHAV3oNSBk3Hatq3NXOw8Uahmpu2In84plki0uOILWyU5OYgYvoi+te2eh+
sMZp7OCiTIaECgDbpcAxMVNvIJp76wg54A5SDklTO5oSWv3pFV8SsZaRAqpN
Yd0+qmsw9UTggZps4JP+PqHzR0p1rqU55Xi8UZMgrafJM0Jk4gsIYPtQ1Usx
DLH8QFjjlKTEEteW6cthyGApY0qDdnEKg3WLkMVxffMlIM6A0TxEhZUFjI87
pqBWWvV49Shoc5E/qqnyKgNWSzD7w6WihPcJODwkGKEWBHj7MEtEDvxN2s8k
ImzxR4KCxac98gdanT3M0I6Un4IChqX44QwejMJPzd0kFsVdaJ+KOUSmYjsj
wwj+81hi8aChEEXlHEalHnEaif8fjiObAAYXVCggho68JMuGjzihdw8k7i1L
xuwO0SulECtGvuMr+127furnAnl/QtSpSvVactJCdcmJ2MdCGhszGQIaR5in
DUYAWqsUkpcS15nM9cdkhpd+Meyd4jeFsncDoo0Kqr3d1iouarNaQVjKwyc8
VAbuZEL8NcMNJKtXtWpbvcPswgjVLlk8H4H8NkBbZApGXPYSlNwGd+FTndBn
czoPUuSBKk2sq0enLm8dxSrgORWKl7ptoG0YXGhMpy86JBVdlfr5QK8TJbAx
9+sfR2JxqUYfZQSgo/Qvkja1HP6HrJa77ykjs26BmZYEfdKekVZDGWb1zPDq
xmTMweI5gF1yJqjKXsl+8BmlRoLQAWlNjINDHAjdMRPog5nGlM/+aZcItIZM
RISPsHNBKj9rPZNT+V9WcoBdkWFUyZ+qOVaqkrNZ8eN+3Q/bbYFkZ+oYZTX0
JjfI9glSUb3yYY1yHkmaubSvtvt1tyeFm8KcXiFO55yt+lWAUnvQ2PshQqg1
BnGvRTdFLeiyDVYOumwgLNtbxxCAMLpvf4SH5l8PT02v0gN/4aR14Mshqouq
XPPDXueSlax3Ppx+NSH+iTfV7XUyYM/tbm+3I8L7a/x6hN1fRwvjdzUf9oDk
r6FBmt70IgPNxP8Kdbi9PO2T/sOpgN/v18FApvVetUzUTHlqvaHu+h6aVSdJ
7UW/UAjQfv4XzoXxW0nI3cKKxAL5I+GFlH2nQFJtwwj0ggfBBFMU6YDBbiLM
qv+z+2tkT+dltI8rQ7vkG/Sgz+rN4lgIN4HPBiUZkljyHAV/NVwI2ccg3uvA
iCtkXAPXtmDOKv2M1XedvZ8XszPYXYrOLLWbbys95gXa0GPp3UekbB4BkhjH
Ft+vAwtSHjD21ukKNNeTO/0II3GWlXxtaBvu35/0ps4l7qYUM3dKhWWtTOVx
pzUYNuaOu8OtF6PZogMlqb+WAQsqZYdvREB1ped6wiU9QOoCZBcIGuPsMHNC
jjKywhl4vkO8BsgccEt0r8v9FiXmNNOvJn00scTD77FJiKUts1b2hnSQZDWq
T/Jn+y8fBjcc87+e3eAtBvNdUhFkuHzeHczRhpWwSJoBAjrKipaMeqhKaxub
dQWSO3pI4pDdd3eMcWVKnAeCgPpMrkT7tQV56qPteJz9klWgQu15aO/BpYHF
bBeaE7XAahm/a72mW8kuyY2t7AEawmDcOP7Xm+Accjn/1HWcHbFli/SiP/XS
9eeK3a++sWFCt8rKSWQaDehqd0zWNpaId7Y9yeWhqNQb4BMS3BuK9nSaDRBm
ectojOPiSGR728gI7pjHfR7IqqbszjWknK7qLUf/O7AZ/140OopJfMDyi1/U
Hxit+tf/eYvO2SqFdBUYHyyU6u/mNAt+4Z5OGN2j2rKmwND7uUbUuv7Fq/zl
Wow5c22Lu8JP6bdwDuoOwo1tN4W/v65Niim3TlZwLFLGtRBJX4EtugoCY++9
8ot25ZZz9hlsybMGzHsOOjHduO1IU5valOVZaCB7EicushBEs3gDSoKEkMTG
3OpWsrqlDqnnwF7sOnkDfHs+Q/qvEPeZa6qqr496nq1HDaxTZr/ZBu8zF6zD
x3U72qCTJrDgZw3KaSY+IchMACRmuIwqeJPD9mjcUBB7GOChCswI8rezHixc
cUHf8x6mmDD4g3Pzf5mvpsPJjtX9U2LTYGWmthFj2rIGfiK70i8/R63JL/W0
FTxCg0q0u1TNCyKKgjPzIRV3ZmxJ6+DGUfzWps5AKkX78WeEEXA0dRYkLWC0
eOU8rPhCM48rxshBswrCqXNgcZ70EkxFPGN+pHa94HFM1BRX63TkCyPmvE3C
F6hcprkT9L7fajxsCattLtN7X06piZdMyftlx/+WR9JNfJ2Mq4W3qPWloBBG
xgOzV847VjGfQ9E1eH1IRyjoNdytvK6kfYpHNfH1DfOR85lorpjwv8ocL8ia
iMXolR62P62hC70dNknw/0NMIlxqMgqeVGvggtZ0fb6ZpWCyRy1sq2easIon
wHC4BqqZP/aM3yjq8Kx5L1A4sMTA31qHcO+b9OaA1j7GIynYRaBfmzMl9Dm4
QdYeCFf1Pg79cWYVY3k0QxCjkb4HzDVHLTBVfm7gKDANXjIqMH4Zb4oPnz1U
llGLjwuw65R8YI9SbR9QQdR5uBZg/eRQlm9l/tobl1a++ax2dIXPifKyj/F0
RAke/67dJ8bWVDEG9tUyjPLETRgmq3c51TKLCcr04DddnHghOX6PyYc6Ybre
HCr4+05NGvJ0Pkk2PjLBuaD77MuyVxyCJw4X1NfzIn9gLCCOydIikchYsxbb
QQO5qDnmcpTg9fLvlAh7gnWRycXkAhUYB+Vk+BgfQKwO8Kfy2fZqn2a2NgiP
HecBVC522cHseKDRRUPhqpDYRI/d3Uybk8Xa9fFFOr3v6ib5gYSJPmZDIsoB
nmumJAVcqD/6M0RMwFeqaMpZTeFPln/1QQJGNW+cmlUMGneG9b5K74bwaRu+
yCGsYHd/spDP4bQ/9tqieXHt3khzmcSGwWYfEc54TmA3UHv1dYUbswMiZleT
ZiK6YT2Ry2owy3aIijW3NmzL8makyoYN5LiLBmN9TotBeVAK5e6DnOUcNeL0
JDGiMfmH744c9/VOl/usEuBEkt6G8cwZ/2ui6jebdQFLuaCUePTvYtDgaB0d
Qk5kt+pFWwRRk3SG38XyOkZ2NIk7z6O+JZMpshHnS9gWJwap+CJLSSvPv2xl
rbaAy2elWAH1qKCoGiAHulWCKY4/ldUYR6yNNkBtgzD7wL0O9K1RoVSccCIK
HB65H0EFDM/ux2X7w8+F2wtEvGKPDCj8MFcVkHA5EQ1NjPIg+9nZ/FY/5Ri7
bePw3FpddHnqsWcGoctywu10p/pY0pnPPZRzbxqNgSUem9OsKVcNKRU99qNx
iE53yvHXeeLO+Jj7MxzX1kYzkLB7ROyF+q+XsgKx41TVTKOxQWpuGKkVg1Rp
VDAJG+7aSnaGG0a0Hg4Ens21GLfkJYQmdNwj/je2shG7AWuxrMfVrJv9WMKu
KTZtCPXEwYtHs29Os2sFZexn3WWB1p49tWov3uE92pf2WbdTMkk3rIKa3vtJ
bvWIa7Jq0i1nmf10ZJcbu0H+2SjVVsPGGuTCGt4IZwdHHxZMNZ/Mh7pbQnnK
g0lHdJTAdh6CAAlGeu1G4kWYY1uTAzaiGRGOCxgEvWbxwOYk2DGX/U1EXeG5
3KONre1nyT/tlJ6QGlUQOTsM6iD3tnWLj3SplBtn/7gqBOPBPsY6QEpjrKAS
i5goXWlw4B2H8dfh/pThEPI/Bpu7/0dZkJthKlG6diRPC9kyF7vwWjvHu+PM
12eRP6zZfeIxaEIHaw+Z2l1GTESwSOvRYZ2u0g/Kd4OMzfmZskI4wcZmAzsO
reVui5K/A9BgEQJuNnyVjfkg67y28QNGGLrqWbfr2hFMb1xfhMwSjsCXQQte
zGA5Elk57odNuANPwtSaRQk/B1HCFKuuttEblQKNxyTaRGi/wGzVy5LpMuXa
ymLqpVI96BDnvjIfWAvGI/0EX4f8LIiXsBc+gvI7eefz3XCY+YbR/em1fOKu
3JGLTlpNbshwlRr4kXVLLqiGNESK0umFMtWKJpfxbWmZ2LxkKHZpvMZMxgjD
iCoIwQZRZ5le8SKBs9zj5BpUP4Sq/y1FSG0BJfHyKUhKebpNqkBSkwjxMShb
ZT34ylYdEe0zXKHH16j2gFuI515UtOKiM33rAbl8ajvwFoIV6pYcLTZ7P+J0
r27zvHqZrvvX2XzPfUHUi1Kj5YPDRORDNaVurw2ZJxRiWIUNJ9dSYCHNkqMB
hQKNQsKZGxRk9f/56v5/xC2N+YxQJslK4lNAEotUiqXTb6/GPLx96O7QfNXn
MTjfH2UDLx2jQ18D5ccdARAkzLcAdgIjf+Txo2P4ywBEGe8BYNFpJQDTHugL
M6EWXe7yKvM/E9wykvK2YGMKOC7ErUOuKye6j1xonxLUPraywCWKgd5pN1Je
xMKqhDaceqTP8LAovHAAzCm2nLTifZz2BjXyMOARxi9ziG+R+DJRIIV+0eLr
ebAyVSzxf3WeePCMRkVm1qXvlLlNEWX8Gcrb6EtjGyVrqcpBZUgDFKsUyS4G
SJI7lG/34/hYCZSsih1lRP0kxyenujdibjlnxIYajUy4/ZpO4OhEMRX1AueU
mabevsjqABd6catDTIK4otXwR1pb46pDbcB+L13GHoq3HGTqFIDGqKyRmUKV
VFcwObXX9357MXBo6CArE/Ed7mc97h22F4N0ZUT2uCwSPCMZpIsZ26onimoY
BO4PUgPS7qs51GhSyQktVziADd1gUYN7+1EDSfVtJO9JCnwjIybKWiftVh5E
6YYmJyKD0X0SBDkjrToQ0Q7uyUEPBZZV3dcJL5gqUy4sOS7t24jb6MQ+ttRZ
RbmszR+NAeupLBpNSfwKS6q0cvXk9NYg8LYhJ2l7/W+28jq8J+yZcZS7U5P/
2WQ3h77bDgv6BB5AfPbO4zUZ+JmC6GVBRp9Gn/NQglPGsdmpZpHDMlHNstXm
OfJMSzkpq5XnsonOkvf975p+q9cAIymj9YC5Ky6dGW542QMIBLEVUQTUR3sH
4h4Y6iLkMsxQkgdr25KWuV9R0PusdPNfvH8DgVKU3zQ2S5vOA8a7eFlKcJTn
Z4qI6rSygxBr9s87xx4CJWRSxR04Jf4OYxm3rwnyY4/fWaPW7aZdy0FI75cW
DmnjGeCqpqm56n39uEiRENN2J6GfB/4u1OGhLyGh9feUDqaL7IV6awHuHRSB
ay2u2Ng3qnRJce8dLCTvfyImtE4GSERgt9wcPUFmrOdhrUItQGQoBVINltF1
GjEAsnfK+QBNVMmoJ2H7cf8pUGT8wrLXvvbeEroZzuoMWubpvNHW7IcjDgYj
8f4w3gKjN8gvsoRCvw/zTW9i7fBDYxl9OuS1ai2HsCoxgOBvQjmDL7vubarB
TnI25jYrq8mWgxgcYJv4jVETMrSW5/vUthwD+bCsLWs7rxLXKaCRx+H/waju
Ys4dleO1hworaszYSjM9QUT8NDyXom53HnqcDRcLZyErihSLgUimsHhvK4jy
jTEL496rvPQuXVtg1QmGS3jKNSowXcVLwIb5t4AfHVyK21lqAOSLfplCVPHq
fLxM+LfrYz1MovU+EsLCd9fYHRaEtzuLcHQIQ0SKIWHtlLcdtWHZ+4jZ+4Dh
tYWUHY5UYFn2bpZxKl9NDEkKOFUERl8DyMSJCDTTRTk05gkvSSoFM59NxBOG
pX4pm7gEDPzOteqUc0sRAmtgzn4wZ5g/yqzYSqjv3KAmNFvgEAyAQZkzFmCe
lL3cHntKr4xxiACte/0WLDKBYpctrfANqvnBuD87AFsIkx5UyFh2Avcdne/S
7AxhsfWz5zPGJCRgXHI8gAXL+2+9q7m2YLr77pYXNj8mVZcVMqUD7suzdY7z
CsTe1Eu+Bn9feYcvhtN6MmhI7ZB0U06nrsnrGlPlWNqIYL+GYs7Y/3bqqzPN
2K2kTdCtYp3ncsMvauGb++2i/gVs09GOZaccKgmLqgavOJhy8Mhj/jUlN6Cl
A7U3opyAgtn0m7HFJzf6TRKOAF8U/Sm7wp+qEIqQao1zB6Iwh3XoHBmW/Mbc
2d/5MHmK0gCZQo7IH3XeMZ3dkJbqpYoJYWs5R2zo/Mh3p3jXWha+SG+vsmPl
yBFmOYhkBLAOW6wkyLH6U7rGfVHVzw7I2jYe575s9Iye4MK7CEPvLjTNPe2b
+S/4ISjckJngdCOx5/Mrp3q48Qf1OgPtgvFzdsxjsUTPwpQGxu+bQUsmxs2A
KzadYd6pJUTxPz1lHktEdPrDUHOsWyv7uySE5fEA2/4oWxNVUDOnp3FAigso
sQbaNfEa6e9EsLOxj+xgPiMUMPnkR8XhONla3FrIzZlyMDIz+hV851X5NJUJ
IKacnh9Z/IqLGkCH0EcBR0YwZ0dvidkLxqIjJuIkYOG5Baqe7Y014boS4osD
qon6qSYB7dSiQKj6X7B7pSGJTnChTKeE0A2/yyJ5XbmfkJpylyX472MORY7i
IvuE93j7jCO9Skntjwvtka67C8vby2U3o3gBU5rrUDgLOGZ5y2MqwoLhVknR
kwW5ckt7SAzfrFzUJt5CgkkGIJLbphbyb/BskXDoEk9HugogQxcWZL5FpFLx
3KDdGjkDgzfL9ykXZk6XJtLBgJClKXPqm7X2+ErwGU/HR5QJpDDV7onBTJtK
jy7o9l6kr4Ugd5WV2MF7jCyh3T21ulr9/r3tPqdumOMC/9JD3NKX6kyVE3yQ
NQJ1ffQx1nqjvq8byrjft1oh274szT95FA7nHcow4Nm0fAACCgQkueVAeS8x
1q19LoS++FGV1IQEkOyCEmL6pTkjQpl7oEQd0X+xNiynIjEOrEuFCqwxYddg
qj2gq3opwrL6mMvh+JH2hNC0xaUH+kk/pFJ7k2jwnbXM3yhCowEU5Gi/B4sl
bxFxgyWQD+Jn76Vo61RAw173RmZ4g1jWaXx99bxcqhVzMmPggeg87W1mXCq3
J7TtOFfJLVKfR6YeAXdXAeDXnMzPujq74QgdMjW+PSNc45crMzt/Lz5tULed
P408QRTFleIYte0wMLUvtUPQA+vsCmxVKwStF8dRZU8RMaX4sLs//ZK+YmwU
PxTYvMtW60Z/7FDt0sEURIi2eQClNeewqKf1CsZzDTpGQnluWRMtGCKZMXSV
tHjxvtufElYisaypwhriv2IelzgRG2cNyEVqRNWeUgRzIV5WHJql4P+kUNiM
CdFWnYsH8NJcOZzegOhzrYJRwgTl1Q82b7OihMasG5Y2cjqKc2eimp5TWf69
BSxqnafC8lM4+2GChMp9xqN52BNhcq2pRGlNISyI79DmBkh1bQlBdK/2IFN2
bD8FA03YQe8GMOE5NRJTe374+PZ292Dxc8vEwAlk4ff+Xnl4vB0ak/Jr7FOn
OTN1eLF/wWKl8U/WPzDnuXQn5uJZAyXmmYWnx6CQCXR/L3TVmrUI0EDFD1qH
AoBGkN56cT/y6y1ds4nvs9ZIFvgvw1GnfnLcPw5wq5DcfqRvMiyl2PHH+zkC
/erV0L1eQUToyRt9TOpyeyEBDa/3FRV1giTC5msMyCBAyTgz+hD81ia0gz+4
mSKSlp6IvXegr3r4olmXob1KN93zUMOjyQ+scNIOUqCM/j3bl8mBPZvF9JJm
MG2ZLnMOeSRh72GVkt4oYgWPEe/WVZEges7aHAQ/Hcf09Jg85BGhEiAY93Jq
BNK+bFe8N4Fe2TUrMLFdunhgxCcRhl9zuQ6CN8yWv7FbeAOr5gz+jEfH30EO
iyxAAXxw06qkULtdAQ4Pa8zgiAopzW9Aqku0rJUaYtSTwGr6/A8Ezz9QDKSv
g2KF8zdKWnmfIzlEdFFjN0k1W0LfkaYQ05jtXdS+ShIoKDtJ9KsI9vtTAri6
JE84PE9hF5flkoMgVCSJkHoeyeAF1mxYaInG7J7NRSzxFy8wwkpnNY7wGhxb
BIhFYg7SpOVsuVDGM68axOh9BEi7/mXao7P9gdeNBmZNPF5CAw1Z58sMT24u
xCgT+URu7+aksvMO03AP/ccZ0FgsnnIEsRqMZjcU80twP1uSn714gv1zZYqO
c1QNEo7jPRBJt07C+/96CQ5gX8ZmP/ptC+2pw2KobLgAdv102mhvNtiJWX9o
I0UvNUQ5HR17/hYtnuIBMlwmVCp/iq+h9TkCqJQDIhnygFxBoO1rSME5Kija
zbFDmA05efmzi+KKiWVYYySArOMATiBKfV0xqd6hiHrzJaixIyMFNhzbXrcZ
UpwudHHVV4QDTs/1u4SoRUHmkIDZnG0GGsfNeiU0iFa2yKDlC92P/UTE6TEc
j4pn0nVsGWXyz8eysAtVKUchi0yZ07IOCnAoS49zW3owkujS4b9WAIUTM0l/
Bmd2B6v5O5P7gGtw/2YZ2vyHBiSxS2+IjYsgKoHFn7q1P2nLE5ciBHZnowwF
4i+upxD1Lf+tg4tY0c5kd+FLpr4JyfwftPF8F2D03iwMYOO3NCyI+ztl7Gtw
3Nj9Cw0cehVVTQdJzU2tCd0VBYtcHPIBdLaRTgCOCSlhFrQNFIqM21hJlpkQ
U/NH2I4FzckPm/GHO1LyS16143Y/P549FYeF1rYJwRguqc1dSUJSwGu0xN2y
djK8l184FT9UmQ1eQ0HjQv1yr2ImopuAzGx43j7Y2JEeXJkABbpzI1ftsTwV
NUaU5aFqPvltQ19o14PtPvx8hHRqsckpVQQ4JqL+xCCxi+3bhuShh00dc0ih
zIkWCu3gHCNCg+RYj1YjEBgQYKtg4naBowuh74H2JH6VWPPTnptqo8FQ7kvT
bDDpEUHK3ZzVs4Sp9mTzNENUk4J8C10FRt3nE1PtC8O17jEUft+5tjGVNaME
bWwk1cn1FgCH393vi2UKpTEEJQFE/own8xht4cQOSFDQXjGVlVdmLx0vYZ/w
sKqfkbbfEQaeS/GdODfbXDLLiz8ZkkQzUy5FaUKf+bM2nxn8Lw4r6FoM3kkz
DtaA4ecqdpeQBynYtaddVFJ2tLtezEFvW04uuiUMgJe0fhq+KBxwv3W1QJwo
2GdkqxzktnxNJJyY/0i3PfOZwHu4/PLC2+7ZeNpzqtEF79xeZl/tDr44eUHd
ddPOF7hk+IMkXYf8UVT+tZGWYqSHKLTKIU3jT6jXFjz1iArApaTxQoBxxZXy
i8DPF7zTnVnkZ48P+aLYpaFinnJRZD6bSKytnkBGZxcs9idC+YSFq2NZEyaN
eGUVWO9Yqu+0ionFaZZUeH/1m1DfM0F+ohmagr4YZ1TuKyvEL353Matxbm5m
2gRAUPVm0fwXPcPa6PhyCaQ38w8PejywtzFGW6E726Np2GhwK5C3Hh9r0/kr
DMjIGaMeNU/bkJr6DW46I6Yx0Ni3b9vRt7A5H2k1bNELhXUqABOVP8lKz+8c
D+s4aOLVkC53Yj3NIK0jNWh3/sCZxSy1M0lMY2oLZJjNwHh4Tpx5ituzkM9x
f1CIE+bJFHEhKY2aTGlq43DZoPnlot+c1gc7ivwiA5JWmE3LzNXuf5NbiTO/
y2rteyChDRer0VEErvcFqdMhQgtrlwV7tQHZtzfnAnswLC2/odSm93+w/Wq7
OzTN/IEOGawPt3DC006gLsyx2IseL+o4CeAaulS83bLALUohWDk/GT034k4K
vuASM+rVDY018Fha2T23ffeJAF/vSyeBwaTKL2vy/fVIr5F1gOKcY+FsNsE9
oc4CvtNUi/c+LfUBhOGEBn6+jNYebPvxAA/rBXGCC37DCpNcsiBvR4uoybpF
sCcAU1e3I9aZuzoYK/bopov2kiV0j89EMiwM1K5XjwhwW7M7Kc+8VIN7Px45
qO9EeBANObdajjQylsn4pZAmMPBBDmR9F8PLNyUk8qjJlwFc15ftk4CxGRUE
tdgWDqV3qOnrmvhyJYBPmgCMy22fJspr3zz+Mp8e7aWeq9zi03Hm6D/QLNnI
/N/vAZhVYR/xoOAwvKFK/THoBR6fFrjeIo7ZmPI+addcwiLlUzsVGwKPDxG6
JB6Yaha92SrFt9bNnBSql9l3OF6iLMAaMkTdEFj9gUKzKU0UbC2Qctczt7VF
brgqMb7/K/3nPmzMtDfAFNAXZAEB/nCYgR60IybOOo3D005PNNmNnFsoSJNq
G8czFAiakat1fLecpqUFXOnUcmH4GNrJEkPcj54Jx/z+PzrlVvNSAuiB8+vJ
NpykIYTvqTlcycSvaVye5tXtoA9axg6Nob2JRdOdgCQQi6I/0yY9eME9jSom
EfY5Bt6TVaSliiXnzLL9F5sZMe1afX62vOd7fPcqgAmGs/0ZygOl+ROCxeud
Q2Lysq+ac8EMjHcrQ8FkDTWw4Ui2fq+YVY85U0s3PsSXUH7twd0NSiPw/P/m
h6r+TQZL3hwIw/USFZa24V6LZ4lNIksgyAow6HcACb8qeoeQedEg3ryjnXuj
tFeehtPCmI/sDAdc1NblZxdYA+PmeTMTOkQK7w84FheRXrgwWqSLcRiZH1h9
7Oz6ccF/rXopeN3qjRQ5mK5lzpaQi+Y63pOAhVg/zQFQUkBOAHR93gpfLf3Z
4s790ppgr4ajQAPnxf9KIUv47OR9hnQr+oJQ9L93fpSGZ4uBQ0BkYXfIyKrs
P+k64+Ln3Iu34zzNCruEZlNvtpvPjTQqif1VlfI5ygjrpeIdocFvEsPjeMLw
xmV/56qTCah2KVJgIA9qvChPlbjCtb5rPhd/BfPilJMD1RQayIiV8Z9UysfC
LJkVztkwdzCxUd6uDh2VfsU68ld0AJl/EzaNd3Dy3/5t9lsY5WCKiEpVTEd7
SakcvBp+UOSP38ZP6uSjJcOV7RYOFqAl/6aDg3tJro62oy2dTpegYBBUBSb/
uukLkIr2DRPGiLX+BXylpMr4gkDy1/m26ozwsJSbbx0l2/ZBPRCilZucoIz7
folhkt9hsVKiW3Oe3lrig5C1NFwPqnOass59X4/0D1bgcth9wLt4jISqfaqk
Y8jdp3/XtYFU8VSc20ivrkQxefiWFg1xMfDIyqy+tfbEdktRMSIVcz80VhTX
GZNsTmlQuubxOxKmSw68+C6BFsEDzf6aqR4Xad3zFBT71uaFI0PvMVzP8oIP
kOWKkym3kLDQowqg1/qMNWyjQZwG24YYqcnI6m8n2Lfk8y/CwRey5aw4AY99
psjwgO26U6g192giuyQl2yajK96dAoOqSgW/9tZjwXhl6/x4vdX1BiFIX2ro
x8JwQm/fy1uNX1BEBEEvVkfzxQk/x5caxK5Pm9fk865wtevPJSWZhkNe6hqT
2vbB1JWIua2IQDLV1FBvvVL99B/WD7OZWAus4HKMBV+eZ15oY93/fAM9ysyq
7OSfXA/BQQqhqVTPpJFzCh4u/1pHH3gQhRTCU70HoPnFNa6f4QZHI560OQYp
o84wGjDkBpntkqTic7FK8zTR2gxSHm40bXzQE+AVf08fgQG6ZUW5nYFEGNjP
eJ0y8Du00KAGPhleXI7FN/ptlNkCQVodNuE/scfgF8+//TN8Tn4wXTHQXGKh
fD70zQ8kSvJVeF2F3OhNAWZfCnA7La9ngT7y7DWhSmDoC02AGZ2R2cy5IbmG
BNhGGZnfTzExU+aarsCjc9XPsikh0n2FhPFERRwURLhg7x7UGAH4wrr7eDYE
31k6HbrV7OTNGCZo92PzaptQX88S3xmHeWWijeMyuxthj2hJw95YSaI2nCw5
/OCDHlG1fr2TPfbjpHTe5HRhSkIkGxUtCpF3veVFDlQyP66a0m1SPjkgxWRJ
AgmN4wohrpfaBIO7f3ciFYRZxHJTuZyRrO9yHvnfgJgUZygtc/eUG3KYZWC0
zGCQfpT5DGq6ttHfv/j+2+mPmFIHtQxrGFMSHM1YdhnXTMLodS8ZkXHu10sn
xKHPzcrpDP/fGaymhl/s/0dUUVL2mZUfNQ3jr4lkNrovaiwb83zcxip9Z70/
CC9F9xDdLqsj9oFFY6NNp6bpX6XeyLjeYwqtDGwKw/BaTcaz3BmRjNRgTVeM
f/ocG4eSwsqOPjlGvNkhftTG5yiSNfkVh4iaZujDxr1kOCiax+xoJxo7Md/P
lyNHlYsaX0GfQq5gUMMR2YW9lPvLlDdcOyCP+5LDaM+GVIFX6tDlRLj+tFpj
dMyQvkZMydZVUf5lvrQ4lJ8idCNdiuhADX5k9F5h+tMIQUfZzt7O+ESc5Po3
Gc9Tq+4PCtyK4ubAwkOV/I7Upo8nWYnVjZKaZbisVNbjT0uHsBfVmjku/ofn
izjtfgZ4EFFVFxYM3M4RIcijl4cLeWs/dI4tE4vbaO1lioVoopKF/JoHLl5z
CzS2XVpRIpkTdWF9SWczd90ONI77KGEQ/AeBVRYbrOXAmXkmiz/OCGJCO3so
FjTPtLad8LSxtKq68MGdiDxry5th3NWpmdqtJQ3rzO7KhXYduO5FBoQ0YkXF
DKkHy7IR9cHlAYkOb9daax27CdVC1EZbNBlfMg8zW5+VuFLCqcVyoWdAHfiE
shav7j/d3HHJs+TIZPs187cBcgSbctiFaIaOFoeBRpwtYb/GT1/eXwOEscVa
8fSCE85h6ifaV972EnUbgNcZso5gdXf7i6NSr9jZK5PkzzRGwofhy/QKiuGG
oSAjx6lczMvz2niRd5jUzpfaW/xaV1o3PQjM6Lne4JZEVpCi9vIxzfCjxWM0
+XGKvxLkF+359VSBXs/LIpY7wwWeGFOQDVEOmsNELtUBx4jNUtckM4qb8ayh
OU7xSrDHENyVmDVoTHIwQtwhvToHL/G7+FOsuhYet0YneM0PP5ZDIhCH8pbH
rqvqTVpbBRPp2PIXteZmwS8Ex5W0ElMXXCGVIMyA5Jf8ioTMVKZQTcumpOsr
BASsbGVcVDcOxjz5C7CwBlD+jDzH0w3y/jr95CgarAL0ivai+Px/GBqAJtSE
NGfE2UaJgvgOfqMRXIBYQmB/x5mgvrkYBhDlReXHtKhUTSAcsPb1tjW21y8E
nAYJGfxSsER6mWHhYqVhU5XZEsvlTMncELuO6BKENP56ScHdfyp6MAXH91Wp
Tpo/mkSqNn+WnZJM1pkl1QGgd4dsiZKRXO19jMpxV26lmszF8LHbkR9WlPdm
CH4F82eR1EHu+RwDkufRNSw+PZWsz1E51E409LzK36IwIhdsODYhBpK4fOh9
xjJr956h2v6jxXPL3e0GJ0Gvg/Z7mCfaWwncbqpIu4Y983k4vZy+V/rPuMM3
GdPA0N6Mc4HxHq3kuiKhDhfWBRu30Zp4JAhON7EWjM5TgvMK4yBFE3Ji4a0G
eomSaT1CW6E/0NCIq36BLvxzl6ouxP/Q3objZbMV/lhFbQZpK+QM/gRRuCia
zs8B0LGu/MLl+bPJsPHWQ6sHBxOWsrtqjRaWg7dtYwYCCDqcmsSMY4zWEr8k
g+z9Z9t5h/WSIA8ajmtFPQ8vFMphBCCJdtiuMJj4FCSRIKMb9+2YQV090q68
skZ5zS1GmGSawOhgVFSSwjr14a0V1Cw5j1zSPQOxaVhe0bqYPUTOnv1Y9oZW
mPTpzRshEFe/DuP3SCC9XZQbzMQYVLpLjTUoJFLkYwRGMkfW+hgK8IUrLhnd
GxqOzO/1kknIq8+EXqPBmIibkxARLMKosk9l1C8NwpCGaL0mWOt4HdKdvrE1
ZifuG89GJ71iiTxHeQkZ86hYY0yKx+B8J+HbJ5SEyq3WhRu7I5k8uTH2qHjR
xbPSfuY5GFEAExh2EC4lipgVLPIoYrIqeOYNTpuw6eq12ztWNGBoKQnBHNmO
iSUOBzBvkZLIU9wsay5ebE1ieS11ehu5kGi4mkCuSP1a2Gnua+nh+S41K4C9
u/xzzkgHe6g3WHWQ2CDikouLF2y7ctxSEjVwLO5cF4ekCj+an5Q+Tsr4nsoT
xuMy+VAi4rletd3GoLAUTeFnC6S/UY+hQSpi5zxrHg+wWjJ6K2KkkcbTKgpU
ZjGAbFSj46SdDcRG5jmBO8riwb5huRh7/UC6oZh9CKmdnv088ZY+WgWtpP+U
5Ra6Ea4COgU/m2oy18NCfavkrovynUTSfK1l9FktB3+YYQk6dqXor22O1NTn
rWheQ51wpbe57BuaN1QCE88ZR5TencTDtJxSte6AwpbouR956vzWpnTllu8n
VbRTmswW+d39qRla3eaLXp3sY21Fi/xe3nSuaZ3smGMjjZY7+miUoM9F5sf2
0BZJM1plxUK9qQAT8rV+qYwEXL2qnT/oFC5u/6pOSWtPDYwc1o2k/546y7jy
1jO3MYHaTerVANfP4KbdsjWeL4W2HLmHxlxpYs8x0GI9Dva1XO3aSS0P5kB3
F2EE26MvFPp+GZQ4qjcCE0nbtPpMFn2z13WJysEfk0XcJMamsQn9ta0+m+TJ
qOUHMDrTa3SF1aqnL+ZU2Y7ubL9m3LZBqn4vxRr0FXBQCFyGcYPS7foIEeUl
V4sAMswHg7OMSfZuWyVw3fU2cnE7q8+0xVXc5a3OdGRa/sIKutBEDL2wMdGg
WxP4wAYyloQUaz5Mov/2Z0gMIPOTWkxzeEn7Qsi9+hHY3jXoaljdW9n+dj2A
HldLXU1245YJYur3M7oQKngqk4MQaoezBtcgkMiokA53zcNd+L+uUpoKLMPD
ke+TYrQaO+cyPcwxLFXzNXNszlPAmp6lMUKjnnFYdQnl1RBnp5Nz9EIcQrFp
OTXlFlLny7t2WHYXnMGLtFj75gJ4pQhm19VDuZW8zNGUXFirFc3xmXE2JQFA
M3Wi8XivtIeU83nJmAhDtzO1+LGaeXabnusrtKwMtx9MTJ/BaLJvRG2R7DHQ
xt/XCwmJorsEURgLkPs6+HgRIMJiJfqKK0wSZCV0IXuEFsSEubRrsRHKMFWI
D2rWkENOgp3QUKvVUyjOORO/8i/IOgsoY0EKBhPKHEGCgJY9vtqEr/e0jt1K
1i0Z5p18VT5+KgaG+MU/yHIqwjCyS+33ZD5WJk1WbOVjXRbnM39ORsGpMb0Y
xqbTOVC43ip2OpibQhzn2oryqegudGHpFP1DLFu0kRlm++HEhvqUnvIDkwKL
2xnjKKV86xjbYil6+7jEtbmrJrWfufodRvu1FWdJFYPbs8+ojLO+f6kiqymH
wZ+cpe6mF5OX9zZprx5HMY/OAkTPllQBiaFeM5T7mkNl1RVLJ0nBzxB/FmAg
w0Ay8/LF256sGhTM7dxTVZloj9iAJbZaQ/vowK/sPVBZqI29r/47+NAkrEjK
J22/UWLPAhGVcA7GVlUOSm8To4DD08yaxdvAlRjyXCY4tze/1EcgohPnkQTV
f/IsshVjbzU38UTt+FuCSSf3gH6o0VYwmh8Hi04pHREf1KLKlxLgzetwJIGD
7//ZmiHAOTpcAlFgm61JVkWJhrTnhuwTOg1p9X5DBbGGZctabjxIqSXX5Vea
QlbCd9EK86hVl92Wl3u4lnChGJPlNL+RDoPCV6ioa/1ClKUADcBMlpwLeRDC
kNWN9uoz2rPrp8L1qIAMdPBLSnk38KrqP2icbf8GghuBzWafgOt11o39Djzk
O3mMBEuHv7e6HQHQngIXIo9cg+AyG7lU6SeGSA0IRORUS0QBR4pW1PYyI285
mb8JPNmwXnmEErjgbTdiaieOpuGZAwaoct6X4Ag7glHqguZprhtMXk1oOGLQ
sgnJTc0voHxvqMRy6qUucPQhqqj+6Wvjbt1UsABE5suwCp/hNyhIlgXSdgLe
QlqH/42YI91EPYASMw0u0+nCXNkD7drbPqcEw0v2TH4Czubih87dtTAE9jUd
SIOEvQiJPVggNlcATGCGzCavEXy1S5YZgQYCuJYsWK6zzb4W9O4u6TBGJl7a
dODzvd5ynD9IBhIWiSuszcGRBF6I+8evxQfBdedhOe2HprN3cA/F1UT4Sh1N
2WWBYAZSYNoU2LkT2n+9xN8cxZRFecKsy3HnDkBTg9kiax6UG7eRXPEN02D6
DFNDqs9c2pSgzaqFnUD3N1cdVKITaVdpOII08nW1kW7GlDmNrA3IiY7botM4
WTSH1fcvdBvLQBWTTR8ZNbQDLtBdCy4Vkb8bMW9pSDdfzZiaJjXb2JLe5pjm
A9aWYkEBdGw2ud8MxYUgEyV8kfbZ+BMTcl+D23YhoKo3fR1JhZfhpS1SI2TP
plFRnGU7mH1zs8Ee0EefY/+YvUcfdAmo5q5GgvaAtVMR5tFvEg4th+X0ktaM
xpPRO9imUlGb/dvl7sTg3V844qZ5v0RAodi4AWFEOg3O9nbl1KAj92/qIeQQ
/d2U/IyVxHDwWqp1DHW6t4/FyjUtKvWuNLcssiVSII3mMRCUr++6V7hXttl9
wTNPgE3BOhGP11/dT9Gc7SfpsUWMM/y2v/N8y7UR42Sl+4EGZHopVVGD3xSU
c8FAfAJHaprLwvZOT2VWv4tLsMUAbBCiv7GtMM2q8M5x3mJ+j7yulVEvF3+X
mRZgvl5RgYTh8dv2txZhS2a21Uv20umDdJ8VwK5j/euUTa2PqS+YuLnl7KPo
pzIR1i2YRBEZlPIN55yVMF4PyDobb0X0u1bp7n0TDVu7wNdDk6rw5TeqpB+H
iMP8suMk/snOPwiUmkHmg6z1LrJnTsuui8RvpFmrrpxucqVVa8U1rW/PdjTu
CB1VwIc66Qe3RMjEPA1WhU0a6PBMtHz4e5/Xd67pty+TENeFHf8C83EZQAvw
9Q1AwXSQunB7mkPfIFt5eJNo8s6QWsJkvSeNxvxFY1jGsBTT7J4SzSK0G6pO
Gs1Z9hEgjKc+YOhrHMSIV+uPhKY0fgSBf0BmDzHkAM2vn5uc6VuXchhBLPXk
K3CFfl6/x6nrCr3dE/oxUD45i9perAHsjWRG4Kfpy0JkgZNs7LZn0c/PVce+
eHrNoRCpCicYqn0/aV3pqP4SNpHzpk+zZUakog9MBwva0vlcO2le4AatW+6M
WfB27SzgYQmsKEmY3NXfOmmgroXgi77GhYdgkeMMsmhn7Qey+aTb33K+UZ4P
5PbuWsBDflZFlR+gQ9ZHlVPS26PSjrshEhxraQD4rNbWDlhTMXkt6b7cnxoP
NLy9QyfIFKjvCTcagf68eHwD7wNjI6/DtTnMmKBR2gFDx/CKzDlAYxnjYhBL
+4OOQSv2/lHabTOrSZH2QHbd4GFjuOF+jXvv4NbjJQy0zF+Xh0BWbCsTCtHb
2EVsBEVCHWFb8z7fqX1qIyJ7J2bTuKbMCOSUAU3Oa43OaN712B7dJJVse+z0
D1J5cxbLGqJDWJfksrDjTTpT9B1VmMdNThinoA+ierJEY01/QrYmimh8mXW9
XC5n/VZpixSXYDPcm0UI/nARRNapgIhazjUzjiPAPOYYC5B84LQDn2e8XRdl
V99gHaHHvuaJApATY7ZiAuf6TwitVCsMQS98YkWF9jU0yFkgncpkaaAWDqeL
isrYHzFPWEvWt3zbXfhfDC28rMlkL5yK+g/J0fosWzs41SBjtZvwKhP+m2JQ
V71bPktURWEp19hmLMcRU9EwWBZoPoebbsFKyfrv1XsH9y0OtPUSJcZhvSIK
t9bE1S6bS93ZrUxpxO0f2r0lzkx1WcbHNe1FkxosaqX0wzkjmiJl537KhS7e
rhwVKTHbjuD+OWLrqfvV8nCtmj3ZcSUg6YmvbOyoz+QV8gWr+VNM3Nt9+zc/
KaMatEWGmD3IBnX0To0Yc5K3T6qgTU4OP4z5y708jpumZ6NqxioTybjrO5LA
w1eadOWQcPR67gl2zhGqsndqqqBAPl7aLB7aDDImuGbdoz3QAPlKqXCnMbsu
nv3RD3XGj3zaZeBc6ViXuoznnM6ycUkhz4r/VuIASBliXS+BRSb6dc9OLnGa
5pfb2p3YNesrrh1ox59HV8lavW/qhqIefMlzh07axEellBwvIkL8uOj2XGR5
WQBB3JNI9D4HW2+/A9AuLGWBtNBRQ4Jm1eaPYA+vsLrMyDDyNl1gu5ZDK37X
UIt6ngjb6JP+Xxlv+6AB9montkAKMd+CaQNk3MwBH7cX2jhXYvaMgIEHfyZD
eNBYk8lhQsU+AuXigY3wM7f3r/6WmTndpPaO9KdX2sLGUynVYErOScOmBsub
RBjUCX+tFu6+YhGcxqI/JDJ/aHuhBsGo+FSkQl3TclGl3detXAO6UOo/W/iV
mE4DuPl/9dY5vz/l6Ib2h1/IxmBAAadmMGEZkY/GeS0RLQf3+qvBpKNIlhed
Sg0hpnO9nFYX6j/NWrPPyA8zlNpzgJSSPdpHTyLSLBuu1XVtQEltzQ4zbGWG
KdhNesF+Jr/EXLEjyBsxTtyhDquU7Zk0i7NeyJyEzxH3UTCA+6uNaN2vuF0y
6RZezPnOxRs3tRsmQd6hZ2rQm3HCTQqBwcqYrUjwbbTV3d2P3pUqPYIrcw52
rO0xCA+6pi88ZtP50lur1subUiqxdBfr7DlY9lwQu0sGG9NBgdtaZx3sAo5I
2C7176gsudOctYUZ5j8rAd+QzmcYcbppqrBhr82fWnPxxsR4OiHefNVZrkkO
xqRdeE2x0j+l9zpjtEZ3V13p+jRhuUGCMIswWKJS77VqFZSl1b7JpC3oELKt
va05BGtsHTnEKimH0cpNWO1u+jepTt+kQCI0aopn43DfPuv1lv9F9OYepKjj
A4nxNoMOEJ2S6EkLg3YS/B0KQfKCyQ8V4/z4k0JuPFsfjzsjwAIB/MdEO5Gw
MbGm6iaTmUnGkHwz2UwW8PtsQFxZEFyMxe+R967VgBX3d0QER5JvP+931PPV
NondbVFKXB3ZGdMaYLP/jqk1mQROcwDeeTOt9W5hKzwRBnygCuZW92HJn/A9
11jIg1Me0rYwxmIR0pT9ZIwScllusy24+z2PdZZnZyyqcnSFarbO3F3qr3sX
kp10Cj8W1M3blXKYR0KCqmZGvjuYqq6SEqagM6NWbaTSWltBsW+xwAegL33E
8XbSVBrFMzKyl35knLOKbaqSB7C1w0bOFMSQzLhYJcrsPqnpU04Z2uu9REbj
gpYdIXEgWlBO51Gn0opiE19CsIj2B8i88888qVraRmUyPup3NCmwPp4cWFqs
u6CBNQpIaShMNuvpjasKrlXkJr0Fi4mtAaUtrIiS2GZ2hLP7dWIMQJ0pJowg
36rEf2xZA1hukWfCEM+mFxVI+oixG85tZXmY6yEW43HXRgQEvKJSOEqi2RZI
C1YpyT8wmOeZxi91FBu/hgzs6sxr0TFyoUA/YzjPzfqKFRJ76tvbcniSSAPu
CPkxI8NQD2EU3l88WZVZok3NPtoRxUaXpY6KSz2M+RvjojXLs04ed96SnxPR
e5nA68lY2bG5aUHQHtBv5M1oHyXddNuwpSW10yB51vLTwlgnnd/jQZSLDbCW
xG6yHlD5MjQnFej1CJOKABQ5URVtwhga1VxwX9DaUQvE4ms/SgdRKn4jnZ9n
T5zb71zWJCbxfohIPqIThdcGXk47amqFIwmGZZBYEkD4mxTXaSKynB5nA2nD
tAfb4lokU5YH6nYP91oV7n18wCdgFyvZ2uv9tRGnGeQ2/WDGyBCebtKo47k2
EuDNgNdmwUIWDvo8JUs69BLqEdIqXLb6VuVcAQkkYft1PxP9Nqnw+w+hV6gQ
StDuOdj8yMIi6yLTVdC/s+60s/to21pnoBX0FfACu9POpcA+Ju9iqaV1KuLy
KM3eaTbu8UfLIx6JyTxcUfGDQ9eAXMpjCQZFubvOD8reV+KnCW9m2+qGj8Ee
XfsbVCEPfvcpsDp9tsHFXLuGIgnDza2bQ9CfzX2O4AE0NDU8C7ZDCAF3wJrh
nBWkASAQLlpVuAkJ4AuGbwTM0uBGX0siQO3e0lk1tyg5FCJxptcWzzdkUswt
m7dTadiXCKRaHrbksRiYqmq9yUgAJl/iUfofcH8NRQzm3wBYzMhsIj8uO/cQ
m8x/1+gwMpNbw1NRjT/UfenOe1QfA1yMom2UcnmoI8Zf6FOr3Rjy2lm2gMoW
nkDFhpBTkKxSZltet+tooEjseCyQtBeQpzhRNA0Up1eTdbI7cgsGnnOVfwmg
QoKFMFUOz9I3PDvmo5QKLU6O0xh9ApjbvExTwS0dqX92QhItSDjOXHsvvm4E
jXJjjieWG3Gu5OBDQ4k+Wc8u+chq6+XmCwNtYDsKbuxp86FZY7W6zQnyGPDM
iyu5awV5n/PtQt6XOutJr+38T1vycUBjYq1x9df996cyagqaJvvj9jCv57Tq
/psrTFYayqLWrqUWhdpwGPX/NTkeQbFNpaD690uttBWnYNW3xiV8QEC8vQK1
abkFAN7y9WtzTTVBnsXmQokUgN+CZTKKECAHvIx2zUUWBCFhxrEC8EAMaGA8
0K2oI/qDBZTOHFQkf4zAn0DJEllkyF201R8zhX37/MQHqNpNa22zXvx7FgmF
36YZJjeFLH8QO1Z9yrNLwNnarECvb+QUrMsPACNBmgQv6gEznyTkOUasJohO
kZCt6DhgglG+ZNtKZQxtshq7yx5Z4tudPXFyyCUbhSwGed2ZotMEqPaUSsyK
QYiRtmsWcjnHPLCftb37PdA4KJE5JtPe8weQa8xlB9+UfPcdjy3CDh4/p+gG
t/3sbVa3Lb/sUWp+YuCKG2zZolrBj2x6NLLBLZi8Kbgcm7cfPiaKYD5VK+0W
wVipZA6Kzr4sOMOw3wLOrboq+k5HrWlBeae+uMMeN74oLW4/G1KyMitQMebi
qZf/vP4AWGiQiv2baBU+yL7lqilEhkrCnv/bHN16k4XYLpraGVLCsP8fDGjQ
ux+y6wXnuGoEPQUNjIrPRJ3TLzyIsfed0ErvgUD9d5ZsPYbNjRhJc9SXrIod
V8VR76tFtjYtT4BEdT7SYXBI+XDzIoKlezlEOm4GDJelRe8pQpR5KYuAL+XB
JJXNdi5a837lrU+b6lu8z67uYDxDcax99gaTKqOQ8B5OFpviW+n4rIPsZDJ8
EEWZ9sZLqGbi2MI4mghYbpfWC4eiBRiWHROhRDyRO6+xa/h8B+sX5+ev6i8f
4HM2RyWHgbsv6NA5WOZEYvB/jmOgDdTRfBuuQOtE0yLxHrUD5Tr0/2NGM3VR
weMpIzJzkqC5ir/hkBaFg/jY3eIfiZDbv30Q+2k95dtGZSdMy+IDogZ0+g+t
xz8QhaYYHDT6OBWTIcPP6ihjRDWTyttYW+RBcZCKuQ647cuHYZ5Kwm68E0FP
PAbDPVl1U7/yqjLJksq+rTQMEkNNh1ShWH3WXHS3/M20npOi45pbnZQiaunW
51l4CG9l/QKyF59G5SFzsjHWWX5AasxTt784PZgyWfs0UKaes2vm9n0c3a9J
l2LymMMSyOW+b1Zb1vMV/5waRkOFxJQnSIbXYSZbSasZWbe/Qq4voM0SByS6
PEQFChYgHi2t+ZRPCeN3nB+oxjvXkaDyJWzEjnFMNXo1v/PhN7uelp5LykTQ
8OZrZW4FD3V8L/OgBCLn+qgdkzQQLRiz3jkwExbYardommY7Dz8jT5vQm3iG
6qJncOOjxxnnSycyELGo95xc1o2r/C75iWPbq23wvA4PI9xDGqt1p6FTM15Y
N724m6LO0kBlqKZj20TfVxO6Q8OCijNU2J1WCD4ooYOVpSpZvTv+XRVGNroD
mKKTiUSxC39xTzfIjxpIpuJg38KQm8MRVUm1pekEKlKd6gt1HPgAgH3io2ED
Yt+FYgqcFo/NK2ahX/DdVB81LnWfzYpN8OzVRXOcB/gGIe4gKM7hbB5Q8WSO
A4F11GW657HqWLFmRa3MgYEfuxqGbX/U3lOb5I//xHzMZbhxOXI/ROvkQDfW
m0lCCmGQhBAmZXW834H/Kph2VERwJ5IOy/VyUHpIeolmqKeL0TF8FDMI0K8e
dqfc6QqgD08rHvCPbL6Q+1tmFYUuH0vgx/rb1xms8kFiqwf3UYiNUHLwV7iG
ju8QN8AcWCoeJm9E1u7QOF31uKAmSEzh+A0aLAVU5TCkieNjq5TgAGRsKKzx
3N5brbreC/13YYUWyp1P61FIcfK/omFzoMzeTwij4R9JP03FAsDw5awYGMey
eMVtO/x+wbGdXVn+gRj0uI/qh366bYZMmBSHMIojHaTIgzuuMZcCHFw42Wrf
mbej3gQCju9M4BJperLp47HWaTfRblOGNEp1DDtfYibmpeQNTM2dWmgrG0Mt
gpfwAe2HoFKKHxAOdYGbwAfrakyMI+ar6aIguaVCEh4alDja0QI57fqlFh2R
sUJ280PF3wnuyvEjREsGIGrV7oPY09mkafkFzb6sLeFJB8lgPftSaWbhQISu
aKKzmfHp+8lsc3GuiEucxENLnhlu7iescnJA0j7LPo7XiCCYJ0rtZP3uf1uY
RDYl5IhOK9tOdp4ErsLQqHtAvOLtBr4m3Tmo9QKUXMAhzj4BbLEvfGgxRavk
DDpj3lE80b8BiVTc1SsBFfKMUUoQ8FGPO2leMWBpMwG5AP5ikr8cNecJQhp+
dWMpNFsz/d/gOap1OBM7YUL0HisQN+I0ofFohH93QKOrnUTOr8YY5a20TOFR
Udis1he3N6ToUHKfrXNA+43anUSgDS07EhJ0+xKi4zFKOpahtA7KmvfuAinD
Ta4wNi7C7u3qRhbsWQCFLurgh36hbF5P38wH3XlUkm/4H3BLDEqX9QWadf1f
g6XUrdwX7t/X0Ru+FNf2AOy1vn9ThClANwuqJXubOBrySzBduUqWa9F7RPZE
ZpvdeIgzhmfoST+WwDf2J/UVjOCtBwjwrzI3GNK7K11Dv/+lfJFuDRATlZGx
o+anpa2mWWDWDeINHDphQHhjLrKHESsdPZh1Ia6SgCssmyzY3fsYwYOD0Vu5
++iZouoXpRyugrsZ+LLvW3ed3T6nJut1+v+zN6/ol7gllxx5I7nN0Fy/oTLB
EsX6DqDiWjccZ44jwV8t6ULZfh2zLLZTfoCpg395qqrblJU0jYAKNeycz3Ky
9hIirZcve+siN3167yHWJ+sClEcc7rkQP+4dceyh16gDgcdGeLF4oSs0jOg7
SY5U2jmjN+35SDZlDmK745Kyn7O2BlHaYTe/oI8leQp9M7X/+4KPctEp32il
CLUPGW7iH9JjcHb8mrJWiM6+Hu5Cwrcj9PTDwp4mT09oO32nYlkmSHQOzgcG
uzJee/nLQ/Mz074u6jmGcDEVUFRunpJ2s/8TRMxD+LT0t0CnZ2FlReavElex
hvoeJemm8bzlXzQAyMzjsRS0y4aW231MflhGqB5+YzQaGM8wdllqicdGpH5E
dOu0Agux6DZ5pOuKTo7VyEsyCJ3B2FeZMiWsQP4deJgrUtBoPQCicRAXL0Z+
QiTY6I8dC4cKhIYFGByrmhwz18GAix3Om9dWJewFnZDwiypWCIn3IvmmZfEL
ztvsxON9ctHjN9hfSezEVQPH/e2H2guUVVkngxsWiatg9up51grQ+yfUK5Lh
JuciKRBP/tFFPXnRb6tq0MuWJD27W7rl6WzJ99Ud5P1t3KRis0p6sN9dalFe
36E2SOOJaC9weU5iAL6vvTfQEav5tMKjLn1eftdexEqMjpQstsY5/byaNE+2
4HV2qdvoKpUrPJqDjvaqMjKWDFUUdudnpE54M4efzaL8XM/zknmw58SI6t95
PmfYc/5cJAp2GhGDxYLx9RGUgM/6k5ci/VJUgtMbqXeWWx9odj0PkkhNZKel
74pd6OW6fStlIW/wnps23asD8piwku9q1aHg7KBRT37uK0Zd1ivjzXrxh4V4
ht2R3n+9w7FqtvHAS0QRTOo5Mikz5qZKdSvPQJq0YxiYUH07DsJW5+QMz2Vx
N65BepeEpwHev/lR3KCOrqBFy3cqHfOUO8r+2Dyx3Cyr2Y18JgyKMQkGwUHI
L3F5IsoK5oGR50+x27YqRMrNsqpGB+e+nF9bB3n5UzjBgqxllucuQyHta7oU
CF4RRMCAvCsWNnGxJfdkItvtUgD9oL9wJ3fUYwClAHtAGUdi4aG4AODK7N32
qXCjOOdRlX8SOgwp3X4hS4MQKW/qiaqBL81fDXzXRCf4vP7mqudl7oCZY808
gwy13mFYk9sIljManUs99iMnXS/jxK6G00tUhS3hPzz1hyHsFv5HGSpzZzxw
yQt4eJfODFDxB5j8zfRZ15a7p63gZZelub0mRT4TC2K2mfJNAK+j9u2iQjis
G3ivcZAWmO4tch2UcrRi8Er02xBoKsT6pacDno97MgawJ4K1rNwya+OGF2Hl
gCMqx38hpUbhk2toMB1kvyqRF6zmcfujoU5gquWUVmR5T38nH46FII9chb6s
53vnolr+gnLtEGgKim9OO61ySS+XVWDLuHVBgBx/n7erAige+uzinyTTaWoC
lzdYwkn1vm2FmLhKu8wZvNFDmqTqASj2w7KYSEL+z2oAF39r6EorLKWtuRGy
t0dhJjYG5z8IiP5y+SH+hy1nyJgdmFlT6Kt0WNinTahAQUzh3pOI0vzqY2Pm
rcuTzEmOfpByRNlDRWMaKnlVo8SKZ6u8TNEpissHx3RxdxYst50zU0FSjVPt
jj6r0N9z/RsnBIkw+U+282/EfFv41mIGxbve1IfQS7PGLPQJoPL9JioRKFhi
z2jHeo0wU/QeM/GvLHsDgKWtTAWqvNRjeoePuRHgX1oaqsqgjnnQ+LB2ypUU
GIkvNuWmbBTMsOCEWHGFZZM7UBo3xlOmvcKb9JPIT5+1A8Om9txGmWSccBQc
CWryXFGCxStFQMl2QRt/VCTUaGFmGYILd3UblmwwZR/vR8b9LTPd/X0TaZpb
Tv75y72vft8hRzse5WJ4LydhYB6s6n4YwDMYyDdt41zLvrA1JpmZsLy3N3dw
orFpiFiG5s8vrPqV81wG3S5h1w+zDQwr2w39kfncWZSRaT19e/FAlFWGIbdu
KgknMSPE52vv8+WnKDn1hE7X49byUcRhclkOKGxwhU+8BQEsxNBvZuJK656A
lMcBMJmIaPdYTas9WJSLgdR87uGFhdZxO/r7RCQcnv9fCXPzeYLnghaBtep6
6CKM7kC9CKKTdRoXc40G1VsYMyNbiZWx0YSqRffVPK66tjGRmnCQjI+k8VOu
mooKqEaTrYBhu30ypVEzlcCQe8psVfhh1IqN5InW8FZfEhSkySXTYYi9Mof9
ylq6ZXHofdlmriLV3L5aMVnQdS2f/fwr+vgLl04PqCY3AlRQvLyYpHzQBEkx
nm1Q8pi3MrpYC2eawdhaotWvWGNLTt0FSkM7ZvSKn7/3eBQjNxRiWrKAbUzt
Oe/ZrO5JvETBk+0FWrBWuamYl/vMJs1tU8yt+7TsSSlIcSkglftn1Ogzw/uW
Q9gqcwlwaf2SfApK9ilHwuszi3zrwfKRleCJ3cx01s6EglmCRMyo4I+2T8c7
QspceZn9otJ5CvZ2mtLfisnYXS4xiQ+PuZdgq0qHBT2lCD2suX7iRGsKRwFu
laAyqWYaWA9SrDL1YjtBmunEKqQqvPEM2O9pGwNK4LLjG2ZxG6hr8Nhj0wCZ
TwX76D28KE0WtB48UnQLQ6a+JYZk6fq58obWj/ILDqZs/6x6WCvx9owRxdJM
LLBLm0aXeCDf3DlpJyqBkXfM9/6URUl0uJHn19z+LmPgZa+JKok3KdKVfXIq
nkem5VhFpnx93dRmxQaX5ANrIMLYhrvbNmIPu5Cy30ys131rtMIFAXp/zczP
XCMGPv0HTRvYexR92sDp58Uc3MosJdqR6pJa+z61T57Dts2V6v7dqlA+R5DK
/exq71m3XnKwozJsznWXSAUk0WTcPpVi4fAgCbVJwBLtjxy4Jo99VPrTIlnR
72ZCW5zXIqkQTqKY8my8k101g+ZWT/HGJjhgJuac4bLpF8BH8FGcYZh6Mqce
Y6g+8MTKi/fQjG5qy1B0FMdx58bjlax8ltnjjniu5URoemhzKcYGzsOqrQzm
5Ln8ooOA1/rhJm9aLhOQG6UofR83lIPFI7CaitYPcbgsDhL2+UQza/KH1e1J
aE1qaDMFegkE/lsboq3N7B39PoT9ZE7fyXwsSeZ9ocZBk+yMG/Vz5RNaG10w
fc/6ZZ36PXF33daR1reFskFIaVUY/nkLna0Sy00liRaiIw5fWLJIcgeh9TQa
MadQ536HGVhqa7Nsdld2i5RfCena7f2LMpiTNNq2Zvl2T1Zrt0TN4Jqw8/vo
QTI9diP7XzLRHI9pscd17Y5FhjL9m57EUG40d7ln256NdGrtiw1A5op19DVT
A4GIY8w+nnRHPjkYGl76SN39OrZII4dMJXi12y8mfjz/03e8Xgc1F65nP05y
w6HMQpkGOumhzEMhf7oEllkpr+MAOvfKu+Bpim4nOSOD0CGv4lgyap6xIeVl
d8OA3k2seqjvIIL1fle9OpRVLOIOGhacupqB2Vmqu8j/u+coGUPbaLuOvps5
NvJ885E79emfKVk66+r6ht9mbPxgf/Dsz27Vif1kG9c+K/k08ASKtaaS74aQ
k8S/A4XbvHVnyWROOET3FLIqAIrDH7P1841/pXemf3Pk7czs8DsewFfYtp7e
GIB/FM1bLCjmbkhD3Tb5uXHbLeYg0iiE3YM0Rg9JO2tcxvsHl7vfGLgeydMF
XJ3k+Yc4WNRf7YOHYxVhLLFmbUrtN54WPWvWnzMDQGkVflRAd5i2M99QNLaw
BEX8N30cCEE9X/UefaKwNfXHiALsF58DRwhJKtEurTTMkF8L9hjsgIMhwUOL
0oestM0O1LtF4OmBlgFIaf10vJaCHPliQiivJuVD2Czo++EAOE+x1TQM0kFd
0e4y7BWQLn3FZAxhw0LOxt2beCj7aZkoPfBFMlgwrQadV8PB+HEU5oRx/7IC
4ezw9JGKB+ExX0jngcF5+2XPiTse0dK3dVZJTkLZxN/f63raM39+EsbqCuQU
jK8cmAgYt5LsSJiUQS3x4hc5ueI4YyQPnQbPQfl7cBJVDaY8kOgWPfgjYp3h
p7hsBEpZ1rwvVnHhiqQ4ok1hJd7bvVrtgBl4Nc4AbVXhPB0axFszmUJkfdkX
vuoV4kZJV7xvarsUz+C1Z46r4W+uiMCshdjDkr7DMi42U/WjW+qDVQrD8j6z
fWg2K4ETVn0LcA0r+CQcifxrzWFTGswZfOzgjxfgCD6PMArXj0dbM/708tCR
tzFw85tGRvVm2UDXwlM25kZRLR98u6TxjMQfjP/FWkn8HxEIR+gV9exAD4FI
9XubKLjHJCTIw++Ddv3N430Q9I1ARZkyLtAFOVoFTxpLf0DUa0f/EToxfPlS
J4FGY9HhRX5/kn1NcWECWAoPdGm0GuXschzG32tiHS4Pl5id4x/nvoSR62ut
XLcWxTQvMXt0egLamby83mr9ehleeJiiBo0cOUoyZWa0O53rJYyb0PaI94LS
i+MLIfZIkzH7AtJuJyhvzEkmwbEcZQwL78Az6qe3Qq6kUW/3q4i7P9O4e1+2
q7mZzdEea2DVoyYN67zTdH2cLT63gRmtGtRukDbKFe8PLCLRR1Lry4e2AgqJ
SjGkqcYD9KNRISRv4SSVInm7eb+e+KJ+6SPQmhgwh5GPj+XJFBuCSs4wLmIm
r/SPo8To3blZ6mGZw0gn1a3dShlaPmCGADmN9BWiVjpM5Cd6iWQGTHttv1Ul
f4PmGpTuFn4MlkP40htgL52kBbK5HAeOmbiQiTuNv1ShKagnD1lgjWxCJ+CM
5RLqKYh7pJtjtQ0YmSWfAnEjM4F+1FaEud5LsccPRJJZawNOoz/SlmS4TaXx
S0mb15JMQ09tNicPByJbPiThrag+mPC2HQcFPqzi5fCPmrVM1wFxPe63OGTW
XrO67ew1JY20fhnbEMt87XZ8SsIW0c1cW67D49FSCJGfgikGlBwKlhtt6N4+
ZKMw4LQm1wwBBVuyjppQIrkW4R3gOnfcqZq5uZDD+7SojKm6MV2A8d5iJaD8
+NO4OsyHoEqD5YOJAcDOEeK1t3gsoZUeqvINwQXC+P6cpf27sQRI0R/KBUHv
WTzqz30mEeTemwCIOpzctER6pPvFTwV+NsI8gcRSWcK8HqKdlvZ04hRYWK26
PGkNqLWPpKsWd+jVrnlu5jIICeXk8iP6Twlc/7Tk4jXsICACt0ryr4zJnCmC
zSU2xC86JQ9jpHt8TzDzd1lT7cblx4V25f/XsgqDBAK9UjBdzH8afWKCcLWL
yWNqobiKjYDx3D9hpRPo6f1M5tyT5NuIzhzxuPzhcWikHTaZcShH7Ezg+Zdv
BXw1zur1VmUPxOaYT/r139diAr5zAtIVOVc/gCmy2wAJjv8Fi9dNiwaXSEMK
oZ1+ogQFyzRRBJw2Xoz+VmQ7elp0dtw9cj/yJevbAxn8R+ZgmHGGe+qMK3Yi
zjTVgFz8a2pyVW814ZXwECZtckC/k+JTDxX5lZfegFsTPLJT3D3mJwaTz1YQ
Pwt3Hgzm3Ajn1viDzgeU3SHI4J5VsFvVeZta2ibKVJnpDDjB0eziipJh66wn
m7eKPh/c9rjAfNObLWXkp6e12SFwpoWEElqDyLTLQKB7YzwEY2fmi9I2ZWpx
TIlRg26ZuznkmOZFBv+CfyZ55c+xSxkq6+YrdBXSmjZdJa3zqCSt+4Gfg07B
8E7wMHQDfY2rulTRQhAi5yoPjchEWAWbB7Ftvczu79uhdgjwOUJ0J952cyaB
HMja3jHfx95XlXvZ7TiiX//t+pWcLhGn3nxkXJPjCz1P/i55W7ssXurJDOQO
zmcBMWB/9f5DSnDESBAvHbAQTP4sFwqAjQQwJy3BLumPGMnqiSZEohGjTii/
Fvcv6wR6mazF0g+dlbKvWLesf3wvLxav1HYHXjzF9h74NnSuFDPqDxBH+eKU
VLAzye5HwOASy3i+jaR+GfIMcQ3cFjzzmsbB8bR9pTqhtmgwaOnf+wrp5+g3
rqBCK6oKYwuti7AB0r6r4xnQZaQMoAzebRU5eeN7U0lpCNCFImDFuL/GB45j
/NL8naKA/F1tU7rBu5yQn2sUaY8JLkt3VH2+bb+8R9/vydqDbQD2dvi84SRy
HOiGAkhGPd/+FbSCd21XTPtCQbWPTcx6y54+SPGYnwF8aNTh9tBnAeMUSFF/
G0Ew3d12UCFiAfae20J3VGVDjlkRifrcKgqSr2MVXpKBD0JrSagfRkNHy3O7
W4FF30VYBVFhiqj2qhY8hh/U33DrQZVIDjJQMJUjIsDSD6PyYsIRT1bTyXO8
t12txKX3sQ52VDE0I8iL9+7nyf6C4OE1cq4bfEu8HBFJo4iuhJX0KiHHDqw9
Umi0R4ZFI9uy7BIhsym275YE+cXYaf6oVnfkpzuGyBHh9p3DIdjm6Szm6Cvm
xvwkJjbfQeRJf2fKSHMqye30DE2c6Xq6Rs7gJVBBA32OwwSSVagTP2Nlu0OT
93w9o2vVI1riVJHVN8oC4ffcz1mvsCAoxvdlRew0E3H/UUV4+o4mm0swaXnx
F5gkZ82HBtTwiI7XRYpBXHcGeUnz3rTSF/BLFlDS44waTvt2ZTHZvJQstRZe
eBYuLBnHWqEqh98PdxtKUiJSDhX2bfj/P0rZwnIJxPmUdo6QQ9pRiwkmKIRg
9kw8ki3JTpUxMbCA1emrJU2Omt5iD7kkluanSPZRlvX/AF4JmA7Y89Ig3AAR
bev/JYGCv1Q6RbPfX5OpVXRr/oCo1gH+Wjr5x0K4NGnG6Jg5RkSYAj5Vj2kz
lmFhuk+aZENcNoaMQD0mB1u8JAheQGy9b1/aQfl0n/9P0wDBGhphSra21W+N
kSuiP2t6CwoO/2O5hWJt+FZ4TDd5t1o3REgqIV+ed57c2Qzx7kLPykRuBrba
RFHY+MXii+r8PTmIxx2dfyIFIquFYc2Er1MPC1LQ9TgEMoHIFRPlCrmn60uB
p5k+UsOsXLfE7uFrnDqwAkzfyvRsJESVpu24NK8/2TyXe9SQ1Zcg/o9Lm9ce
n4AkvoAndHimxt67GI4zxCYqsu+bVnwNma0Q3TI+lh3FFLxRVgD0SX9X/M5M
HM85anbyk11Y78WUtcolsLICltk5TIDvrvZM74wQDnWa4J7DBEk4Xe8McAt6
RdJSf7cwJCnjO59kbF/4UqIIBPcTh9z6mXWJxpu6GP3VwQOuZ/OeBRXOiL+Y
mRn6KmFSepvBx3VtqFUQ+3Q/yFP2g0QKQRuDSKY5ouNI1SCwairc4AFxRUcp
05A/ZTp3oZuYyiRcybdmif+5AmYfE+IARZPhXCBS1V4UMqKt8HzaIa7/LbEK
8kea+gDlu8g94PadKzd9IqN5CURgnYYSizHJZ68fA6PmLkPJXxsFZyBi3GLZ
O8FRGVQZlTbyAYmMfUtaFZI9bnD4pEl0itEtLC64CNT00unN2MSoORmVhhp8
iLGf67ods1pZSeMspaPbmmnGJuIi4AREhVdxit/1R0xGJFdvW5UBTaA4EQQT
K8fSHxnjwf9Ja5P2WXzW0iHMtvHnDH68rI9Iw2yVqsT5aCiFv/ZTOaBV+wDv
Rz7G9U3cSVw5sSrJ0eXN2WdfTLcc1LYp8dFp1eRxFs4+NaoR/fD7J4UM5hzM
kBPIW78+e8/JtUj845yWAIDfinDKb7lqd+T+LhW9/MpyxR0gXErJpLfJAi5L
1HMwkAaEW2ivwcIFbi7eh5O/EOA6BLY4gJOqPi1N85V4yjghSQEmimNnnDnH
dW31aEO4ZHq0q2M/1YkV3AjBXLF9OvFiTNuLlZP0FG5fqvYf/9vsLZ0c/QUE
86Ry0U3CnFmfHcrVf9d0g/54b0Rp/MiJ44TZIIok5lELkamfsuX3RBeaglyW
zBHSJUGmATHJJU5ZsgTvdEFcnggGSvzLSt2zc4BQIl4BhnsPDG8gXIS7Le/g
MmSduF8oc3E0SK3Pe6O8SQYwxSTpyNBKqUu0FKjfsTreEyXeoaybPnlOp4l/
02/NEfY6YSe5huckCOfVUlvgFbdP7SnDDlFM+hWz7aaiWXiUVPpKXoLnxU4X
vM756MOuHzAiI4CcZIp1WkJ/nFE3VszqUtWS1Qmmyvga6K7LavJY66H03h2j
HLn/dk7WXl4A2umv6tbUPGVfZ7fdyfoHndU5cb9NFzyc0P2ueKymKzvtqxhA
d288ZSClPpO4HNuwj0G9xRySkbF659PKNW/jg7yiC6TmOzuKEuQ5Ar4lh45k
wzmxbiuh/5dJLeMXFDbC/lFA1PeZMRyHRhyoQkg8H3lsgC4Dn+TmzRV9ZCFr
NPwx5YpLbvOiXAAR1jNRGzBTARWnP5IhiaFTlp1roOzwg1yIoEMrEBfBTS7o
EVjWz5KcMZ+6NVlEHVIHCURO7PuomvVOYHsj0yKjwGzJdfNKT16MqCgtGUmr
IXKdvz5Tddohm5qKRmkepDbOt/MdCDyk4KMrMmjhiPxdfYjtwNkJQyLD1MuG
01YRBljQHQoU0f6QLEMHOJKFavJy+ceVESz3LakSss0e/0aOmsGnKQvr3+B6
bjk28AiwxuCI0goimXAOef0xg3LC2r/N4tlOm6l6MqGZBoWCOIHKlsU24pnr
xhjwIsoKmSDbpt4pBjqG2sMqpl9lv/L8IMRAOTFnAqYx6pMyMage9sI9sda4
Id5RjKSeN4hqaOAuwkxf+ZIAiqHCpy5oDFbpu6O6sN0HHQ7YdH3tVcngvxn5
uA/iyvueGCMms7YKbSp8iElpvoesJZobU4C418GiqOWKIgK0bCf4L3fDQLkq
yTquZsWg/ghpXip/J1JWzpenLuVGB/gwPXYoOHBf0q11OAqjyUksKsa5uN79
goyvCOhgVuUJEVHHVDns7RLZz3RmxrQ3oJuYBnZb+K7vxOSpOvP2LGmeuk2v
bzNk2YWa5+lxoQh5R+DWsAgttrFDf5oWrZ6xn1xhSbziC9cPIZpKN56B/3Qu
kJOUMPNKm+TjKtM5hfOoU51gEbXfJUsz/Ri/vi1TCgWfDQBgGG97WoTU1SeT
KTavEVwH7Q3i28doZ/qxbVKoXS5y/VIfZNwxZou/xPbRxNHEYXeMP1vcID7Z
eUt0fzoiaheLBLj5qQDWfWVjJJxzCRhft7LPOgL3R32WDVqhU7c8HjH8zctM
GzVKvYl2mXCASFj1I6ylWPcxQ62PiPx92POPrgotHyX09+3negaR3uo7LAty
JdtNo46pOvbUiRAp/J5oqal6TTbeDMYORpcqduIbS81R409z+4wXdmtUUKZ5
NPRORY4zoVImJDdJsrnPgNIRmdUAz5VC3h0RkrHuYoyANjI7yWKbg0XWPKED
CWiUuqJ3li1GtsiCEl+2pRSlFPso6Zt8gpRb3Lph7RAKVOgOnjgUxElVN5dr
0UGs/LL2uW+Pbxh9A72U0ZvGl2LL+ojZ64OpDj3KYR6pdbsOP1+XDxcKcRub
12ZTHD9yYbtng6tlww1PnQt9G/cVClZ4tAqk2XKj/tuDbo/PZsrQyO2gqN48
8wWazj1SGkuot7TSylwWEKjAf7BOXbkALiZInBle9zuUmTszEbchIWSfY/IH
SQu/yhgpxFTZPbcaLkqICghTNxk/9+yYCJSNV/ko8Rp/65uvPSq0EtC17KPK
BJeZnvj2DgUSV4Sly2eZqCzvhtOMuTX3xfaNKXb7jwDwHTbi0yDMosQvJIeY
8ecj6TBPY9K18gZ0Zj3bXu8RjW7++xHLiGA3k4IQqkRdE/8Ceqkv/gKVfPW+
K6P2QYLoBZ5P+gr5sKvMFtW7uXxQLgJpT9k7p9W1L+JuFxbqpayR5VAaNS9s
CN1m3UYnAbK/euaaIOg4v/5rmetsod0m2K/UhuG/agVU/RMxtnYOl1q5cAO/
Flqw8aB9D5TAN7uCDXSxDiHc3KV2xw4/smJl9OkqDVir0mTkOe4MOpe72+nt
lI/65BXOeiEn3va9zMGM1aJInZQAwzDxf+t8kxY8USeV3M5treXIcKrvVs1j
1bK1dxETL+4ik14epl/CMdwxMu8wU5+pB+EHeKoLBKTqPP4qaLhY84cBtb8K
acTD/7w29155N0STHupXTXrE0uVbKtHuxa5T01c1z7bVuXHFe93u52wvKG61
jutyUYQSEz1Hx+pIa/w22AHpd8fMD3Z5sI3M+lej7QJoul11Ndnm9KdNomiu
noboy5B0LOSFfYDIW13HcfwXEX6xtMw+oPBYu1O5mVJ7wl5hpa+soHfbRaNY
mveg9VqlP2tQDlJLKXLgY17snlkWiHKzxYLOLra/CtCx4ZzqECpkgHoQdbGh
idcSpQ9cAqqVMrm1fZCw3bpn3KgrW2FV8jK233SBlqQ0s01pcLjhz+2FmlAL
aMb4UB4odzwDLGkQisFsOGRazhgGtHIHCNM3bqTGcJ9kzqRhwjxwPEDgAkkK
MXe5jMcD9qjsw7CnrYuirVzsuXQyBKZho1SO/0BcjaxJfGwZNZ/c9dblnItl
4Ezv2Gl6cbt8Rhv9oo/oj46MNhJlGYru7RaU9KV6dpcaq5hHDgOnFpezLLwz
UGw4O5qM1kU/V0YM25u9+iF1UWS5/9MrqGM/jw0kBIwionAOmbSpalLYlPCb
iDItgFNAhToAuRKFWvFw8pO1CXmnd4Te442Z/oe6GBIbwxOBX1dEU+cgQ/xU
dlT7uLQVX3uJ2btcigSysrZ/viGy1WgPehxcmqn1lO7S7I4SWGpx8CRnzhKa
141aVFF3vbj9jfdOwO2x/t66050ArClF9mFdjFsJ/ORub/4yhJw6Eh/Ucvc6
nlyLrEawMUuzPXwOnbZ9zp9AI6J6AzdvyAebB7Fa1dDlEoeDxqZw95ewkQLA
C1AV3MlEfSar4bJ+E3vFhgphekE/B6y1Hm/urGTLA0wEGGvUiAZFLOeVEdvX
t4ZU0CuAwWG+zuGsxlcRyV+sPtk5UGs8HasWOroAW20NGX13fDZKXX3ZY3vN
WMUR3MxmiqW/Ej7x9+CbnhshmhqJBw2tq8QQEW39NOgZb8CtSw1Ejea95PVr
Z2TsYE5hFONR6tzVbretl/1GwcR2IpTek/8TDHD0KKgs8NvES4uorwjBNxnL
0qpr+9hg4bwf+JD85yoYjkjtsecTBLwZDVbsQi/Pj8J1VhkzhnV8CmZ5sa6J
ugubioYAuxHDml0xLc20JxjTz2XkKUMPbpyUz59Kd8fxNDsQbTgr2RXfHtnX
OuII4FelWRUxPOmR2NiQ7NRwXONdxJPV8EmjKhigLH+a5LYwASfv7RnmR8Oj
Z2S5k3TuRLF4fGQRTof0YnFYvZCxUFeDPc9vIGkJNnUIN3qg/GQAh5IYfQIQ
kjKC6hjTyHjFir0PGoVjUctU5OXNrWG1zw+ufXWZ/zLQjfGJ1zHPreo9npqv
ynZ/ya3bwWksCLGBZ5XsJt/BeVEjOGGCGzpY0jzTVJJ7jAdvjMirvckKn/b1
emJydbu2gT78WGgWIIyTQBkmAbCRGGcEnyQ4WC8Pj7Fob3nMqVHDz4Gxmq+a
xYW4Ga4XSlGMFlEwBQbr07JxG/3reyZ8VsKDJnLhF9CK00moCOUizEBgRi9t
rJLoOEvki6/BgAqPAThGck+xLy/GyWC9HBIiDq8onkyOR1OljevG7r4j51FU
l+kSiRnV8dEn2PDWj17WHlRFHNSHuO7fYWxaAIgndCTBvvOFCkVuMODu9AaW
aq69bSxVIHuKwLJfcJGh05oTYuGP0FcLoCtMmU+kEcLn5xQky6T1Dk0o8htK
MdhLDh/rEZkH5wFoimRI5Ar/o94z7Z0yiUXu6anwTwkPwzQ9/bHZxupgyxPZ
bbtFP8kmdIk1EXEiXzQz96l2byEEh6Qg8FcGW1GVrQd70kLstxrwL84L2QLl
gNzkqzG+pSBTGJLTcF40AZI9e9Mkq7l8Fl043DFIi0+sEoaCHDXcBxEb7+K1
5hK49qncWnLet+xp159qZbpWEdx4lKBGrQeZD94V9KQqR+nwTiovyuAdapGw
LxcHvedVaWO+7VT5wi9z2vovmAWmpSI+cLOwpHpBsky6TxfKp4TFnOFbXz0j
VMj0Ty0k3sGXPDfJU//6nVrIQlZl+K/4Gc2k3tsE1nask0yVUPv+I1Y5VDl3
r8eHw/yZatpKAlf5saC/0Xmxs1aUM4rUO/cdKVNzwRMsGroHc6BON+MovBwi
LVcHoZMEsBDPTb27IGixtk+f2SwyadOukIl5xPv/QGPdyfiBRJokOvfzI37c
i8580VT/1mmH7JLtiZDVTRua8BE/fPm74I8IEwkf1kIB5qIY4gF15TgwizCX
WS3g2dwiXq28vqHu+Tc1mKlVhtqmfJewyH6m2//7HMvxdzpAtSmdpBX3ckwF
tV1snClIafUovkHDzqIbrji9tRnWqL5ILqyNZ+0ZNoZqYk6hXs1rdPagENvv
gPnREl7rR34EctvYGD6XKR8sGMuxmjf3rtX2oOGzCnSu7CRlP3A7MqWx3Ks8
Oqkq2lf/nY6Rls0u0/0UikSLpkgb6UWPb00Lai+gYVI3qELtB4Yk3fkCrwej
suYLH9taF1uOxNXRQahTt01EIRSbSLRFT2OtnDeryVCOOfy5vPC6mnrs0th+
UUEZOPTRqX+xuiCl8T0TWlxa2hdEDkUws3dexqD5fpDfp9wGFOhPWazmAfTz
4+8yoHsOSyw0ApJoz0z+cC+b7uQSchWCkjUpdlQ2yQqPKkdCX1DXouM9MNop
4gUu+A75W2yyNdwnAxD3hUOdM9HxQ/pwJG1gfRcfDQGYmE/cSG3aXOK/wbJB
0q5U8f5dGG+KggZNWIi2SSKk0XKi5zhThsM7L9xub16aLIC/Y6BwmhtJ9Nmr
OXHWpO9zvNsEDCfXMXsvxUm5pYe5wieOVaTa/g55WWdh3bQu0uFcuC4xhuwA
RWp5j6LTnfJJbjdqbgzvPPUZcslccENAo4WfSeAp6S/d/zSuIzKhQxW/H0IZ
jb90vHHa0tCQiRst78R4Mc7p5kBht2kTaBtLW71x36k4yds8A8PtHpqpyd32
noZNc7NroVOwX84NuE3q4u2TS+BuRoZPmqk/26wfOFBC/S+yMPi8H9/urrU3
V3ABwQ2VfTBUsq/IYWjjXxPONptiP1EDfZ96MuQJPME3SC6SJ4RO6ECzKe2s
gDPXdrSa32Wzz8qmY0gsXWFkfLsOnNsKONPQhyXxpvrZ3svwJzArheAHzfLW
XkFR2e2nZq7ZMuPJnWOkLMu30WXiWnqeospsB5rKk087OccsNjaZ7WOmmZBP
RzPy0ZP1EBfg3OoNcjQNTVWdVgZUBduG3uzQdHBZ6CUucH+Sg1i4zRPhBKoE
UDMi2qf+YjgeUZjsxCxDi9TnSX8Q31LBX2T492JhxU8FtPpLlIzaVEaHXeIy
6GMLG81sc48kEOEkDtTLFwL4Y+gBp0JRS4oRx59h/6gJqedJoQM8YpFQXVMR
fjNHas5pKMLdMHOmfTG2/nY9eZ2JsNnI151hEMjd+j6FSDUHxlsZBkcmLUiA
hfUK/w8jg1bObNt2Qvy/BEZxqbpv3OKOVzy6FaOhTmIu97d/qZm1ySWm2+Nw
wrHQPrXqK4K37dhhUEva3HmR5REzF79PD9SErAJurw5QbCPcGTYZt1fp/WEt
M2QiyhgYxB0wXOw++BetoqFPLYsBA21ajp9bK1TEsSm79iTAr7JETX6n/zeo
zDjVhRCHiNy58gOaWxGR//JvPiktPS1PEymq8hoG2OxQyU5xL3xVOjWnJkpD
dXhfHYLSK/IHJ26R1GhQxdeKOwnld+uodct26keTw/hupa4q6f4K8ZT3h/Me
dsiQVmU3YzwY/OyjtY8AEYFdSlLXVrl4JdZzfH2ElmLgr9hhXJFGo90iyesP
7/MF8ft5DpgoHcZLpzQFlgWbOjkwmcLir5+Jz8rtrGrvFivJJ4/XdOSWYJNK
xglRhbpWBsxRBneTIsYwuch4oP1oVSrXADcrY8r0lh1XSfe8PMZg3puonRzU
Zb/YIqy8EPJ4Nd3j0B0a6FbBMClLSDakXfcdXKd8AmPJ9rtAj8FAfDv3lB3c
N9sWceFEwjbbZmY0GH6wflV1y+JTTju7OyxSGTVmSNLpJdhzy3u8RomzqZyl
tiCBpVxPuNRJNh1xK0RL4ZJdaaKZlUNCefsXkIP2rQU8f/d8eBOvQjx8mzbF
FFc88hnpiZ66kRrGsZ4QBZkZeyyxbKTr6viOCXVaFZrVoob1+L6y32gAudvU
xvxrwkOUMnW/6hCaJEuVFliOhdMkEKNS0ELpPG5gg7ctgfyhYXlAsCVDwOdu
Dtxxm2Mj4x5Gmd0CRF0Yr5QdX78Sp02qU4DUUdc1XFH7dX3s+GOOL9cmmPm5
rrrtai2NeYbat1HEogkw22Arub+ouo9iFAqTpgT8Ch3Bik8j/j0sS+IMYJv2
DwQpzbBhTTEeq6b4oj6nOpAMlqzkQe1qR888Kj7/6D3DHhwi12YjfytT2Vkj
hrZnhm5U6xGIZCcBgWh+tHqhEfWL7+N1xHfMRODvE0ERkc9IqEdyZ5A9m57w
UJkHJNR6ln7qIm5DqEzumOz6NOxAZB21BwNK4iSeBJX4t3xOlOswP5UoDew7
oqHdcx1iAB1TDbBCuQXLCj+3ewNYwBsfvCmf98NoyRNvNYGmcOVY9Ut+75OU
LNNxwkpoIa0ydQjkzGWbIbT2RyPq/1UCBwVQWwVPEXnFnkIdcUUy5GidyKko
RVKZOyTwHoUvizkwkASHKWkDr7fU6nX+p5mD30HvnB4QylXHluyDv/6N9Wb7
LdTW7bs6qaTRrWaMFOj7zvHBFQchvr0oyUrfMAzPaoTUmpCFumeKvlYzQwTp
rD8QEf0ihbkHtkogUnBA4smObuwCvyhPsQUoAsFA32UXYewxOD/MFxE4tDbq
j/hlStEtCoWTAtFdYLeVGSCEkF4NYO1gFMd11p42Y/KBYgJMb+taio9rd5uX
vChhkPsyqD1+pvGF1GZokvAqBCF9TvcGqp/1N/gJlRLNt1ctcIyBcQUT219r
t8gdimNiBjqlqk+gk6Zxp+gFDrUXimQ6yn3EHq6yxzNGi03VlFuqk4R5wFkI
HV1wT4t/QrRLk8Gsupauor1CTlhVNugiqRY3Odxf5KMAHj08+pdfYX2sB+kp
/5pfevvDcdFs7MjO0usFagA0UM/hiGbnxF/IFaDfvVlV+oLFN3GcihSGA4VS
sIv++Vo9oPD/jSnh8KEsPhYMc8wm4wqHREvjopYCV1BCWofwL0pOYLr+vEiB
mvoIzOyVLTWDmS/aoEQTNCaQneOAqeSOKqdE7gnTtECirdnsJgaysyXfBieV
dBu1E4wwkxN8c20VNsCP0O/OlGLs8vbdRE0q+Ei1KfKnY3GQeUb7+qxrZjqt
wdrkd73aXA4PGxMr4ZycI/TJX7vyg6Wq/CQS+BwVVS9VC5TQ/2glGA/s2Ky0
flZSrtn7474GKD5XVhLf8r0N45zFr+Ixh+p3+nfBdD6dt7Il9xFa9KNBD92K
2M9hAzJb85ckWYmUFVcauPoehaPh8Ld7gOXImQdW4KDJwkyqv3HLmQJjLhVJ
vrNulqIqmTJI0TvFT97cXncuR/j1cBzfV3QLrxzQeYm7q8+hkWhTxCNKJK3Z
1u6W9qXNekVlqydMGSeZmb/4GJiPojrD36ry64/r5FlcuqZB3s7qPQWFphHy
HYirDCOtHdR6tui0g0Zi7ngUJx5VLxNR2oYf32h61OPhBLOT4TJKco2CFEJn
jaJpi42ErcM44DDyn2UiXnQLXXBK2MutEq374xtDE+VPlDaFL9+ifLjCO0kU
wz1uGKIenVHtkij2NZxGEhaLIyRPgRzA5fI9bIRLFlzenKKTVXCJ+DOlgBE1
U9JAKClUvUUusKOMu3lh7ZEJpsZDQTwU8jiWfE3sok/PpGgQY7IcIvJKh4jg
mmeNCg0WsE2kT8D5W1B8Civ/S+dqp4bOIV6/bP3PBuVw19KYMQUsTxHgy3Q4
oWF78dR4HKmyjESuu+t1kRKk6B0+cgjb0HldRT38uc4c9uQRFZHNTLLiuWxZ
G4dB4kxH884/Ee7y+QYkGeUtNhMHI+OegCUMINg8zDVqDpAdLiS0j84V+FtL
7PNCD0xQG67qLDFJhF8PVP/Cqfx6NIJr3l5PnJagfyw3Lp/09d+iT2pfjGna
M+DCo3XyXP7DYC20VDrmF1rm8U+v1Pk+etcyfFRCjxIE8FejSpfepzoUewiT
wRXp7aQR65e+Jdy3rlnTH4hAYZ8XbbSdLEqfkvWG4m3qLII6QkdKrupDWjkg
hsJzWeB/8vFWLjrjvIRG6tTLCKqw9wVOzjJttcJ3l/2cgvP6/WVHZ0+wsKS4
dweGDy0PfO8lUaTpvjZcrGyNxgmCMGpeo9OPT0lJCOB20WnvOSaa0VHo8jdo
InR6L8aSP4e/yPQxEZ0p498kTqoqEnmrLCVcGa7w7CXue0IREK8hQs50Ejro
VsC5VfXZ/+ns2cbuc0AGds+u6eA+jnn1ma7H0uwYwjc53opgJpelFkSIh5Hy
rJNMHvZYj3DBcmQz/qEf8KjxLMWihVMoAa0XpTktv7A+ekfEcRM2CNmLvuFB
YGklQj5IYZdlAwJFso+edcPs4Q3AhcBR90Yxc5LlpxX/k1DWRd/5hmE9f3Xz
GD0Cft9IFLzCzbCYzJftfGVQeh1hpArQjsLiNwYDIoV5LN2xAAuTUJP6G5tz
CDctPQMCwAo205YxdFsnY27+ENMoDb6+2c+g0N+/yj38+V8mBOXnCfo9ptHD
PSG4YCiSNlgVI6bIayFGMDUGL60PoV1K5uTxokpHrVfej09+Ewx0dwn0XX7P
TA1VvCEr5t2Q88HJc8BJlbOZWu2dbHeW4Cci852KBCHG5xdCaqzHsC4FElXU
yWFthGXeDTmbp6a/55R8+oCuydSsZCYn/6zO2JWYp3VszGTdr0m79HvbGVxQ
0PY4A2perlb316KS63aCgchKFev+bfV9vaA+QhRdqX8c+5EsoRVVXehthgiK
4qRALjuwT4+vP9uPsZs3XKCa67pvAmspTkCyMN/PjuM/yCVLezg2UYQRhgKC
mQOqcuv3WF2hwLsvnITu7SRw7KwadJJSISGGtOnQ/SMt8/QgAta0FMBBSxkw
FO+VJfNdA35QX1rwLJ8RZWb1rST0f0BRl1DuUIVPI1CHsD1V1pcnqHEPcdw7
+FxSLLQdCF0bfuJuslHICI071l3jKdLxWhzwf8T9n9jRGzXL76NrbZnwt//R
kIeWuVXp2sHpWczFjjLxYaw20cM/iy9CMaGuNQPCOXao8MudIHI3+RyLazZ4
Ulk+woaTJVsymbJ9xX2j2kaTxghzNWlmjPImCccQrOWFuPU1XJ4AyJGNRU28
npMkb1TJ9LXySuOKLj891aaZcluMi4mhDeqo9CEciivSgxa1DgYzMaSQ08kF
H4fib74aSqrWvdVFbokNEpREcVdb44+HZFtDOe6+JsCkIa7x5bBLau1iGEmd
2mkfl/4SGqXUMJMydmv6+bMMt3IYaANKyewe72ZUURku5MgEoAUALxt4wr06
c3cUigFm3Ga1ktDrWJOrjil1yv+XOl0jAMFMYJJuJSWY/0ibG6zQEwQ/qjSO
eh7yGKAAp6T3HuIL3IQWFI6RisOW7Ft9Nhck2sb8JkbDTJw9N8RJlKZ26nWa
t7bFx+XpcWXHahTEkBMBEumIQkhjr8CnH98fDRxLn7GWFh/Kb5mEXPp/o/vF
cvQMnEbEeo/ncJ7xlkAq5U12aXcZlJCpjqUvia0GEZqjwDONgS5h48QLZWJF
sKj9b4vT84yTqLGLjbrF+lnFpLe+7Dyhx+DYwLpto0caUlD7mH3/NRa6VEi1
5GCX1knwpg9kVum1ETzykepiqqHK3E67UYdFtQb9SnGmceYiJ6NolrtwnHfl
doaFVPOZJkerqvygoR4Odl/TEXR0q2uAGgnKqsJZK2lXx2pWhuVJ4I2Y9duh
pf54VmBOEy+W+2UJ+igU+beiGmZ4H2py1DSvb3uEUJAd9pc8LuiJksagstnO
UC2DuUPCuRjox4bL21Ho6YNZ82foHU6rJQsoSYKxfSURkGUI0RBQ6KwIL0ku
o9/Z7s64k57RoFtGyqy8EZsNKTUkB4gdgBteA4uTdr2QEUTWEYQKQQs8mL2G
OJG/x5K+zP6fMu65Flo/rGKrenAnSfWBR5Nt94QNM1KeXoIilBm6WrjpRPCX
N4YU8uKW8EP5YKjHdi0sZaRDigoVMNhFycfq3xl+WXZHhccY+OsWAa2mdTsi
7i07vVZ5RQBxMZbkBE6d3BvMDLIcyu9wYRFdMeUAgqd1UoPly6tQUqGJ8jWk
CBwLZ5MP9+6h/4xhK2HVU1Q9lbD6/9seXOxUEkKjd7DxjgeTXOSpX8a38E0S
UNYjbbXCeigT2G3MDPMxnRjlc+aMFjGLbc4ZNqDjJOeyoNxgGiEuEZlj7qE0
Z/qxVqeZE6ZrTmsB4E5oo0CGgGeTkOfp/DvY2x9e55SXchCKESZePVay60M1
cGdMRQ7dmgk6g3fHc0GobC0wo8xXT7ceDHU3E8YGapSaXCKyKP2mGT+fhAyJ
ON3h7y5ndY589anzFiXwbPtaj42HR2mbARpIcLJJQVBIZ1pZnwnNVsJnzdBt
W0ZXY54l6XerrnV5pHppDP/Ye5s7pQAxpbtbVBKMt4W9qj3uM0QcPLnIzEws
JIDtiLbAvH0lzxFS/aAv+GVL80+yu9DggYcHZByodkGR+Uanl65ymrxEEqd6
lB3lAe9RMJ05q3wyg7afMtl0QsoxhappNW5eiOsLvSBJr6TB8xE9XfwAMxPl
Z8W1z65GqviNbYizWCkroBF6BGMkYp6yuDvYnGHlwducfMYrKzWlUiGnUGI9
a0X5k93C4y9+MuRxqtIIPH6if1xWTT5hxrE1Ac69qXYXc6DPrNTxaVxu89bD
aRBXXAqeik6IkbBBRPdH7fAPT4M3WmXXSqxPUI5vJrsQc97kQS1ETq2TPlR2
ehiDJVNTeRWhh+mSf2xpsgUP51JBOoXud/Uo6FZ9vrUwt5Of5p/7E49o5e7C
kAr0QZK93saf4n6/qz4e50XlTrVTdaMEGuUBZDtNMJsqCLde2lIjgGr5zDak
gsHB5nEk/Al0N5Usn7AFEis0ff/lSSu3j0h7WK61d1bgYj79YvXSXVh+/gHe
q5viVLoMLHPuoRQIKCEnANCldc/SRqRuRXeCNnUbby37uwVQHcqxUS4DSvhb
hQb3tNdAPz/y/b6Vg43VvfUwoQHFnneMW1q7Z02MimF37joKxq2S2DVoTouM
hFRGqmDChpYSGS4U+NINmwdXSRs6sqhtIEAn47GdN8LumiGHkf0/uQVfoDwX
tAg6osonF1DrYTPZ5dFEMhtYc62G+7NNsxsihoyknlwaqnSGzB/y1Bp+Jt3n
O7J8M8nKzhZnPaBN9JZr6YdjZu+YQJ7rPTLafllxzS6g0wwNNF4gNS7mx3+7
L45p5RtwQEgOy0Nf82MrRZZ65lksenEGAXPxqBYcVBVRoIwFzJp1CZ9aCttt
BgQEn6OyfoPzyvHpXMdFbU0tIgGjnCdIFcakNZcVwO1+/RDmGRCRIv0PkZ9L
69+mqdVzKPc48+QKqCUErmP47Q+IbIpJOps2cOgBcvGZd0nnIqdfN3v92v3U
lMeEMIJl3p/OvXViFxNiJt+eiiwh/M7JyC5mLSKzDlOFhDf8ONMcQWG9SXSW
/N630o+n7bNdHV0iZmzySYAY9GPbgTn+lvUWwnOHp1+z35xYDr/7oHQ7z9rg
vFsNdBV4aHwmDo9Z6vMZtiAa9tUtHsHFqytNs5JkvaDrb5zAsHCkperGuBgn
gLQpNGxTpmuTQns1ukKujePg+g0X3EDwn6zSgEeqIQ0X2V2VSEvPioS07o9n
Jeu1pRVFK/042kI6IFWgEA0peKquwily3XJwy6IOYRJaa6UY2lnlhWUBdo5c
oZdiiyR1JB6dh9QrQAV3Qe7Ej9rkME7VWZdlla3jiXVsmveiDK9vq9jBbPW0
B6bUv7pC9UedSFZXxJ/oBPs2bzNMdEkvidu9yBg+MXGLl5pGNBFR132F8IBw
6WB6DEEmRHGBoki/1CLqBeE6AZQWT3Dfe26x3m89a24lImzFbFeC2qhXALMJ
7PDcDe3X/m6Cqf5KRxLGhhCRv29fgaWagHojJg5KJj3VgC9ds6rZskjxzTX/
VsV5rFVhygYp4z49+Oi5lClZfbcbC8OLbfQl551+4W6SGoiGlmct4o5rVhu2
gRlfbqFtgtgLQ+Y+ij/pr7/XaF6x5Uq8/Jl0vRIAbZmNC28Y+nPpEE/fNkjq
sp0Bh81PUMqTsd8UM28fvvQ48DAxKGVu5tTbrOCQoH/DkHV/snlTVGoIoHBO
1W3mn/deHILXNHoywrkJHc4TOQjZr5/KHXoY1PE0gOnmtgDwcwltTjVHa+tE
v630PnGnQ9h8R+IDEmTcc0WnbCxftg91pIVKkDu4DQ2prLQIpAY3G/pBp8RV
YBV+AE4MZFLTgjS+SIM8HgVRCYC7pEQSgDxoJo5Yza5jGvD3VoN6cCa7Pwvx
h2uB1z564fm7HPQykSdFTs5qYkXzG3yTTsf4I4qXh2EIbFguu19YHaOU8AhQ
fj6uc66HG0fTDTfsgJ2ocd07wmIuFY7z9t8Gyj8OB2qeOZBO6iny0xYTXusZ
bN5TjL3UPbil7aWzwosuw7QeJuWl8BLzX1V81ddxw/MhUcpIwBBXgOQ4TEkW
V7FvGh5j2PgOfXyNHeIqO8QMTNk1X/UIotp6YVFnTlBlDLNyWsnRAz/Uqu7K
nYsd0PwAx2QQrFjNu6pE1uUoQ0+tN2KihLe0T3Ebyg2j8SRZgW4KKMXbcJJf
Mv8CKAm5jBZ2A+WdN1mwB/HcqtYna00dVjH66Kp2LrPSOtacp7g4wt6Vs8fq
NqYBZpW+YR2W92awl5Kuvk9Rx0LBmO/Zyd4KJs+iZYfXEP1dotGh2yL1nNjg
OdP308nDHAPUOB+NklU5IR+88hbg5AyRegMmUMKUdtChPblE/CzxPo3IXTfd
6VFt8YEQuFHAxXl3vCiSbGNE8MDQB5UyORXA8zjZWS/jKg4DY6X1DjG7KL5r
iruepRXIFVcILoXSzNjLoCUuNAY8b15rmQ//nisaflknh7CeY8ugrfXuHQI2
hdGD/grV+QTF3KU2zTo0xVAucQoHElmavo7x3HJdSLvRBaKEMKnHLbPZek9g
a9v1BF98kcfd8Hn4AzTe16DyLvQKsD1zrHJAkpJ5AVVoXDyGAraVyFxIPUJQ
2ibLqEtH7x1Qmanumh50DN13nzkFnWf9GHMuRWr/tfprPry/+OhHDjeOKNM8
AUsnA2fKJByUZjwH+hVlyuiaIArvzkpWdKMR9o1IyRIhJ09oJtOH0WCnIr+c
rBrkFqMvlsIqH+3fbYs6jowq8TpeTCVlBfyLIYdmxvw1ES3IX768KQMqYZ/y
YEY60/4reQXrtoWUIFZGLk0X6x/nnTjwnLUg/JoYvl8wZulFmQF/8VhA2o77
ES6X0GBRZplo4jy1uh+8rBy9PwQZWcJ5D6+iRQHQoyBZ7CPQ6or0KzSLvV9p
1q/GBYxKmq0ceAM8vCX5PJe74cK7cr4vCHoAUw/6szH5Mo6garchKe6N80y3
LctIoHjLKxaZU8GojRz4ecQWEZuo4xvYKE8QHtICcEHPlXsOVXDRzDsldjWO
nvhBZR1A3gNyJ63bGNsL/YqoTEDFcZO0HaNGQpdFpIJE/zDyp2P2R+oppatH
FnQa+tjudKqY4OT4x0eKNN5S5UVnX+u5J26Q8e+0+sUgKxP2afTox2y/NjaZ
XkFqjauiHTZhFbcVbf0nC3/MU9ef8WEER1SjM4eYNTkFkQeap2ygjZt/LcoW
b3/LBLjxfkjsUh2Ift0Q0/FBiU8AodYP6bYF08MN4/k8wMh6zkL+ZuPVl6N7
QQVeXGOHGMnwd+wZ3BfrhaCAavZ2Q9ZmCuC4d6mJrAjRSSLAVdU+TR3UcSVR
VqZnix+W25/upxfrI+Umt0AvmK85Yfip3NiOiutiqYrfLPJ7F6j2RF35HolQ
AvSEHXcs+Kt2RlIITq/navH2fap1WUGtPBkf+otO5mfibjs7J2S/rp/c83cM
NO65ABlZUeF/1fLMuqIYttANT9wskaCYrGFpFqcgK/vU/k+1fHabyUT9M0lX
wHrE7obMGt4bpmBbt65yVPIJy53ACUTfuczPsUQ1Zp8qp4+FqAjwrKOtqVmi
yEJhBMFEC/FcjZcVJDzCacDKSbKEBT+9hEMTS+FTa91tuvN1ZJ9kCH/GKubM
OnJBcx8h/QnLdUZp0ykHA2eFnW42mgvz0xQ/AdSe4YGxwmcbP/8Ucz0zdBmj
knFuYJkTQZLrJmSV1zMO+iJx+BJ7L1PpRbWwC/APPeJu+8nLirKcizYI1/7Z
yHKqqL3Ao4QX3xu0MvXUNo6WvnvOZsN5vBVrY7yaxzd3HkboiedV3DdLINRy
TYJFHVBDlCFoAnGyV4GZUlaPjTUZyjR2AfEAIF1Ta77nje1rayltAel5q3ub
tInnm9AP3dT8K9f/ee/FZKh+nxME/ESun26F+MBQqXfp2WHNhct5IY+9pSBt
sIWjmqlygsBBEgrdIV3+TQ14//m2uLsd/qk/s3z/YCrOfo2httTZ4OtGBpQ0
gNTUfAb9cgKF17E3D60M+LX+ZMgye/ZpiIZhyiqMsBpxfHmwX4QrXhE+efYs
qMiKLEB9p2a1VjcCicHwi2v6NPUUuYU1PigCR6zKSyRQS7TJLDR4GdPKoeN8
o80Hw9Q3cFKQuPzA+AMNkrHjYh+uyHl3iCoan/5Sy4O5rq1aHQlNTK1cLt/2
ZFZkn2fEUQMOiWRiAyDdRNSczOmg6a3knK/kB6gpQ8ffm3Un0v90WrXPjdrG
RUPRviusDxDNxQWSy+Zq0hMfJn935WITTl++45RMG3Wc3kV/kv3CYDsn4F/U
lBZJUzqMCRDpVON4rmvQnaggWYwM+k5tQ94axq5v3iL6lIWbxa3TMUR0M2Eq
G0H4EEU39RfuvGyKihy/dnfj8nHh1R43qHeamelJT63qDLzNC42HBPt5bQ3T
9S/Z1FwNsje1asg7HBR1SFd8iOngW0zf4vPGcrcu9yQz5ZgUfS30B7Sy5W+i
duAE8Th+0qlUgPw0Fqqi1OIBTCgQ1OlU54UkEP+sWxIkIBCHyawc8MBFbZ/G
fXpKgmJXY0SkCycKoFhcW9W+pJ2keOHSlp8in3AHLMupb1JLZXkca65XAO/W
OSSOIZpvVy8InZuUl9Ipg1HiCzIgfJgZg8OY3Vpdvyznq3xUj9lUqeu0b8Rs
IG+a5hDEWnAZjzfNXYSWRQ+tjaWs1VF1k0zOQl2l1LkD2mVV1Y582gPvbxcC
fDAiJy3pbZzy/0PMgkqDGiQsTSvz16MBnvxSSfSvxtP5YE2UPijGOgdwdYvU
mWwUblJVMujidOSzglY/C2Z6CRPZXQVizOf8QTQ6XyOEkNzzqOmyVeLjQUYh
4Qmrk5UWA5wVPcGN2i5YlfBX25vKugnjC3bmpodhMS7NIFzqN35FiwWIYSoD
Y17UVG7GehexqGekeB2lvH+bBBHIt9DOPcEef+ElRWKqlUPjrGDQA6/X9cgp
LSqDTmRSsefm+ctH56RXFNwVAa9uP/izOtJziSw1lDbc8SlHgap3lF5p9OZO
enMo2p7ySpejmgSddhtFtvSyS+6JGIHfNsjTzAHJDF0HY/mY/5D7wZj3OQxu
TfhzkeBRMTKkAnK/tPbs6aKhmw9HgDhrb+3F1EuVBn6mBBk9LgSPkrhaVwK0
xdpAO2t4Xb2BBaiPHJACKoKzYUP7yM4ZRYfCZAVzZblxnxQpV7mwxAH2QDJR
qsdMs1tvGrRMjzYt3JwYQeCgzAotvBUKC/5+CQs0NwdIMBgdNKmp+GBoeVmz
bNF1r8yOtSSB8gZPSlNtisCT3U9Nhnj9EgSVQ77xvLu/DAx+VctV9Eno0dLN
fGiKTMg+oFRKQi59j5yuBRRClUwobHONldcvryE+cY4TmqB/h9BCo34shljK
vBIMB+48sYsLmT5sStUV1t7+2fLr6szgSI/H5c13pnNxmvUYmJ8z+FuiY9g3
xYv0SxmCyIgk7rNHUZAiysJ6WtnhCXc29Pmj3Saa/nTt2xdW1etWrkzybpqy
ZNIiYF56qisB1MysyCrwBcoJye3tOwoiY1dM3Q24ZW3k4TAoq9gZkRS2h3Gn
d3tbZJ7eSFrykAKc2ydCL5L4LizwR8v6/OM4X1TWZp3roZFjZOD++vVbVfzK
PkEoq7jl8dA7HPFrHQjt8qwJE1ecz8dxqw+iI3TyAasblF06soQKv1eMYYqf
TFVsYZc7eSCKJQLMmsGlQ6R0+2hadudFTxuwTFZTgbu02lP1W4U/qBNOHluk
M3zz93bxuU/wqiN6uu9X3oB4ktuqC1tMzRo6PT4JpYGBBzSZf4Q3b3lDgtC3
FUjfIGBdSeituzU4H2uQoya8PXApbv5G1RpSt1yZhqPu8OWwBzlG2dcWK7TP
y32XQHvDUP1ONjeTMLyHMxHPF5bQ7shSMqbVi+sXnTCP+ivo1TxTQIHN1uHP
j/UK5Mw7gbQR9IpSQ9jSkNxbL+lN5HK22v1KgUpEf/F3gLsn0OEzLips7olG
d8iLFY4WnvJJGGSXNQZ3OwyN82lkNYlGSOQwtUxafVEjuUPs8834KRFkWki/
PZGbWmjY3VEJReWqlwN1OV0fdv4DF5bFRpOh1jRpihNOpaFOfNo5lOk1kTDK
qlbE/sW4s3Kg5vciTO3gftkoiACfEfHkal4ltB8V/PGiyzdtc1rO/+N+GXF1
KEljGprpFLPq6vV2Qzwrien2ALlQWKjrnl5YlUwiFqNoxdFkIpKqJp5eG6Gc
NLHWRk8Rvg/W8coJ+f+RMB4z+5COYsPkA2XnWxa48aFJm2t7BBnHmgADrYm0
TjcwGPSEdqag8iTSJjfsaXb0eSSxx29L5T0DjvqAlf+TemRPD9Y5N8QlTWD2
5y8SVAwOV3LTL8aqwbtzmGwUY5mAoBdwTmy0AlbBv2Fo1s1SELlfJDDsNcnD
qxBoFWatCzg+9SFDurWtKgY4lX4ElF5JHtVAONkUEhSDsCvY/vK+MzG8KjOH
Wu4QvlNBipi1DwcNBFHi8j0a4VfCpN2zOhUflM3avjTgeqw9fTrFE7WQSPeE
KuaFc8j3O1f3yYFRC2gfdjqwKfFt1dmZ1VkWu6j6BYw7BLTlSEZN9eJXMTOf
Z68kJjYsLZ/qGFUf5mmOZyQ3dS4jGsOXGMDjwKhAQqgYsnOzzvub+k/QWDgD
KuJzjDxn/+d61YxEfe9AzOa8hELoIehZBTM4gJr/X+N26RI3eEJ6pbx4aV3o
eo4O2AW7zljEK67DnNVdZQvsvGn+ZoUjmYdJqqnt4J65H/mclPWU7Ijx7IAD
nrGk4v7AG28YllZcgMCpkfOuwZJztuZ1bpL4fg6hkxPKhVxqVcxSmJYtURr5
sS+Fogr4XesCeL1TDZYAkns00d4eswlMf2WZiLik43eLBC6fpxZ9wPaPUZni
b47hEQcYvo82GeWGPWLwmTfrpz4xrx53uCU6k2HFreiBVAjfIhgQCTJSCnRS
vpVae86tXL/LB7fBVcUPUP+OOz9mFZjvRPGpkkRK4bHdBjq//NX2TcTuqiek
2UUVk3Dlo2ZPFckbXFp8sSZ/bOZG08ha1EscVMT7iQnj2F7+ApmGJtHS4ZNx
kdyy9FQPTPp7BWpR/g67pJhObzYxFgZmngn6v8icpsuZ/sxabISu36v3dOCT
s2PECjo2FQBuFOvbNLoDiev4vs4m99L8tjUndQ1wkuGkSF2UTn1Zq7jEUWVK
iUegF80Of+auB0TBemkdRgkrEu4AY7COV2IpY4uiuncmKxkN/KKLJj3f9CBy
NVVxOYPe/HlijejXonZpYRXM0gcm0JjzVmX916Y20O+aT+7kWgo5wwCpyQNZ
yYG63kDmZkPixOAnQpmf7DD6A4vKrZLbJWC07lsABcpPcwAFVIBVFfKL+VpW
3m0XPmoQm+4C59tF8FDenMYH3X3sdMQbg10szLeshu51VJJv7FYCDzMSMkER
TPPoyHlVMIz1lIFF/x/0Yz6B2fW1432Rbh1vOWQ2p+9m4jfZORdRQtnrOGQI
ute1NcDqN+7LfGbR3TVmgvjMhaYqN7Kg/yO4bLQ7IO9eoRgwpJ6OlPulpEHb
RToLQGfPL+mJiQrwMMdFcBuuP7Yaqq8L/uGjcdU0CHVa6dc3jKBMLzJ2O1+V
6ZiwRvqDmtHuhkYCKH2WDOUKjC2gfa0Chn5q3NU+ZWHfTFWohzQFIdAhOXKn
y4rmzlwJruRIgrMIMhrzHA+YkJS6mR+m/S7HCFqs0OJi71C6YqRuybsDcx+p
5ChuYLCedLW+fNXtQnKHdL4ybQY36fCTYHE33FEJcCHOibFPJHymfTuRHJJo
7kUBc61mxo6ATPR1nwK8UFnWICWbeXFY7ICuMVsDeM86C6cz4Tv8CvmC+nOI
jFK/JV9xQWU+ICmkPrQDAugTRtIsTHN4BFnIUQ0H/1jBIVAJDcXfsztYP8yM
ew/a21UvfERIipjwL0Mt6rrVsZqa05NJziqGKwSvBy8NFDtte5Bjb9UGwh3A
COHFFHJKRNQ52c5Yi+qLcPLg7I8T83nmiEnDddL83LTH81SiYBWLGoEAqEo4
nOPEyGwhx3skSxWRK+3F6oiNPTNQwm4Ebxcx5gUHNzfj5p2pF0RqLTuShlEi
djqKXY36pa6hll/e/NNaeVbdS+wGvloG9si8llVxtYzl2Ol3PnmsrFppqFVB
gve6z+Tru3QNW6IY/LWWVSVrkPY2FL/nC3/ZxCtBrI9tUVHrved59OCUW9Uu
hMWtsBOGxkiXHSS2CBKfTcCVuGzSsZoHHtxRBHG/pgdo9mTXEFl7kJmb81Qr
/pA/Na+8M4Lt6gWoXyHyE7t1cPP+JBiHFYL/dwIFVPIcmvosrrexyrW7FtiC
u+Bn69JZfJBY5E4SbcNDA8wGJ3VbriG6kZ4aDuy2y3GedgK36MI791v+IQ4s
nViUqlU3ITA2rHVQkARsWCqtYeInWxRLYSy/QDEMJLfi7BJAnr39OZofixLX
9VTDI73cRnc86XVNJ6AB2DQQbtZGTxmANk9UoNVACsYl86tFVzz/sM1/JNFB
WvIvxrH9sbqJGWc5LWgrhEheUqTuZJ8RNwVfTMIEuX7TbMOpaUDI/2tacL4I
nzaJADWceN5qrxWXtfT8JaVvDYH6cmg4VDcVKtMJGb1pM6N9494s+UVJ8oYK
s2gvmEefBWJxO/wwf1WOFfOltWcZHfsr5ZoaYxqnnFzRj0HVkKqA/sdzZpPE
0C83v3lRfmi5IqDgmqsBTCVQcneljOesuM3fWR8KxnrjPARbBe3UtH06jfMT
2M0eg/JSsz/inxpQknGUGawmXD6bsR2UD+No8aUeLnl3WTeRTO9gEimBUzl7
Xm/KqLbyoXC5IwHRH2dCt7Bpb6U4nnbXzkdToSd3iW0LH6z0r5z5yb9XyGmS
VeHdOMfwriEgPvN92YVBV8b7/SSVPo+w+3TR0CQT3cYkK5/Ykxso5ohoErZg
KqmKF93/gPapeMtmOkuSg2kXKtSDwUyv06igUkF71RsCMAHu7uu4YWr8GbFd
MKE8ZYi8faihq9Z8TxjSICeArKJzL9+vdzVWdzgydr+feg1L3Q5NzHwMpPJe
2WU6eo4NLxSZBCyfwG72oHgwdinuZT20AgikpjvCLfrp6ledVkjsokduHqBq
2TUzovW2a6O5To2KCsg2rpEf46nOR1B+PVCGDime3AMk/kIEqE7ZizTk47OD
2d/dIqxZN9Hrpiw5DdVFAQnxREIjEuGo4EEtC+nQtLr0Ei5jgFtorY9eU9tF
lU3chBZ9i+XDHctxCj83wUXq1eDXViCQHDbXTvitfnyPfbVBQum/qjJEQa/F
TNGyW2qqhp7AjYO4DlKLFN4HnriLerzBtnPV34Bw5Y+o0nBUNUr93oRA74ru
FtgMxsuiJn6VGp42c6bKPuS/At/DhcsNO6J3PMD2EW3hYvpTJ5okH8Y7RGdS
OrlVJSjANvbG8kbxqJi/ZkjuHiJSxR2TDwW+8uLvulaAV64THy/AFz94/+Xe
f8ZlBrQ5hO/e797O8DpIw58yJPrqztEc9Q4OqjCy7QGTx0Tl49M708Xy8j3q
W6woTRjw8WMm2QtXWqn+89ZYqPFw2qLr0FMq3CGM8YjvDDQsCkuD9H7HipiS
jnD/B/h2aXQw6lzkzdXI/nHcJCCrGncesSWqym8GpG3ETtjVZLGWe6Je/3F1
0FZUFKjRhSFvHRjrKuLPodo1EZl5PzXSsMIyedWYI52F9IoJ9mGpIbXayTxj
bJF5a09Bj097Po1jALbTZKlUIoe8sViDyr5CwA0Oj5SHsXAThPUL0BLZMj1I
6jQP6AjhYK83MV10M/RK5RFB/YLLIvz/nUsaacRCqSEqM5oY5ib5pm2BX1k/
RaagjTeCjuta74DnuAsibD9gdGpcm7DUFw1ML6TkJ6/mS9RwnS9Y5teoAuG3
VF2kuGykSZHXDCFHnxBJHJp6FBzgEPQabytIxP4FlYZ3EfebaaSOvWxbBkbK
vVqQay2PUstsbSGmWX3LWlPPy5/4qMY2NxisZN0rNoYBJOAuQoyMBgLhD6tl
Q4pKCcoYEt88nF9jt3NXndC9YNsGKEAdrPiMM8InIyWbY9GSwWzhOB2alifL
0ainzN4EIMk5QO/Vz9CI+Q43f5xaqMaAtgJfLVQZf/HWqjsvhaO0z8YmoJ5/
QM2mNWYf46N5FI0MfGXXUqOV1GRdu9L3acosgzUgk8wIKNm6zlx6i2Q+b17E
13LDXzdGh/I4TBTVyg6ggyqfSLIGkzshfMNQkDUQMBQ7wG2EyjQwErVH4tlY
PHYy6MNG/yjFyMX7wEKIde5M/couMV7mSi0GYLQwdih0EBZLptCLA7GbMjt+
7lfieYt/VK6AGQGDP0bSUiqeR5W7e1PTivk7lTeuGcecLlmN2ln4wJ3BHou1
jEV8UkhsSi2YE37+NNtEpJfeZPrf85kuH5yDNQoUgj6PqNzluAF51ZfjJJkh
/o+idqymu/z86wMvASbbvCoVx0g/K/t/8gaj0BMz2LxC1SI/ThkWaVYl4LAX
CsqCkIa0N2gacY3sE4rty7QLwLy6FvE8izJmZzUDqlVWPNz3QmKwXmOURevR
YKS3Cv1ZTIVfSGVVTSk9h5wyEhetGqO4cduau8oiwHHhfW3TumeAmNRUx2tm
4NVZ1ed1jtlHcpDCA3gpu0GiKtAu5SEdHuAUNv2naTHSbBBDAash+WyOicKH
uKllCsL3Tkagcn+gK4idBaR0iHuZ5Z0OZ8UK6Ef5HKrZ3dyhVRxe0uT14XFy
uQAQzHI1PJ/zKBWbe3aNqKXFEMNqKjKQ5SFW+J0H7MXAdyvl49f5MQE/oKpd
FDahvU0DyXeYaWfWrnCrzwS1Frqa/pCGu2Wqq5pGEZW08zmAZZoEUB2tFZ89
tnXjlyaFXkFQF9L0sWhSKX9jai83wb5SoBzD5WLUJZxMLRt3q12Ccbf6zkg9
b9etrzzOTSc23ywvwwJ/ICZYiAYLHtiPgCL6wfS3owT4Q3SfEvtEBW13S0fz
k7i87fDNtZfUJtusZOO7s6sq4zGnR2eewsnNyDa2KV0s3DD82R4tr4gC76wa
LzPOLsoC4vi/DMVyzLPP7FQU6kVzQnX6ZTCpO0zX2AbYm/4+8nMTGTL9IjIE
lOGzD310qPAB35FgUTx7+ffgDXxRSC9cTIihi0OBLgUAIHr+neej5JSMqFvq
5emE23Cbw68CiXeodhx/DiFduCuTsOvvfzZwVgk6VNxxN2DBCi+qhgXx4jn8
wcoTv9L4o0epMyUUmfkVGr14U4epSqYLMSFXJphqb/Ky8NiJoqlfJzxZPgAb
foEgo2+qVrNm6SSuE7NgiU2FUggeHEijtbRQmcY6DowgrCSCIaGdY/bxKnBy
lPQ+D7WW0R5DJ0gdYWh0/5G+pNmeCqmKOlr2wdTULlAGO+sbTd/XO+sqPhTS
/TQkeAEgaGjiA2pJYZEP/I9ffV+JOzY2HhOAr0k5jEC2UstK28UubBkFvzWX
4PTFR+QEYfxLqewaL1aSkIAfb3aE/CBdw31fg+2gWrsV2GPpgXifeyCllMX2
g/XU/YyDiHhWfwZg+aLjfatK+8uFg6+cAnxeG6+qMiCkbsaUfERd9Gx+CE5G
b53q5I2er2OhuSNTvDfsY/gRAO75Fr0a64OhQJVL3x++4P96ABvRhytllYgM
E8TsBywqFBsHhxZh8/VpkIZsHbx7+TLFGTyb0gBvRTo1sDKz/Usianmu/l1F
+4DPkY0xdsrExltY0X6BzZD2Z8uoPBHH3wgvUoBQmYDi/1ln45T8AwkNqYK7
v5FwxasRiy0emC9u9U02XyKZr/3UBqWWAfyz9qEuM5sGXw3BXHLyvTBz9WoV
8X7nRtFU9aABzZUrsAiecb4Z281Oov1YU97ugGjrdhe5uWlmmMG+2WHwQQdP
hf5wc/FEhhdJWLrW7i3sGEc6YBltlsGGQaEEEC4T6pkZM28vzJ1HvTH+lW0s
ChTbCqalcjdhTGBVZABzitMZX/AQ9b0nIh2y/wyivI8zduU6Fvor5Pqe9cPA
Q6rnjStEXRWZWPTPhbeIIow85spVvn0k0OiX8G+4NCnYvysWDKb9NaehLB+b
9R/mF8weWLILqw3O25lxXfFUDlkQ/XQenSxdqgHw1YHiRJarZ/kTEaeqYaOB
SAlypBpyZac9/PSth9b5Jz0WVHukCUonW6EloQToOEiKiKj7fcfoOgGPAKa8
2wfxIW4XuEYLoKwjyyQTflDFi1+jBxMcLUoDUoDGAVB0+ATJT81wCgB7sYXE
UEmqLXx+EV8sbOpc4oUkKAGg9cSikvUFzCfQejzGH1vfcHcWr7kPhdiuJNqr
LlDPBuIG70bHAzY+a9yQ21iUVjvqE5ktUxoF2YWWWcNpEhbvv92ZzlSs2OH5
Btxh6ktnvd052S3Cjgfoida9v58RuISMF5sZ28BTv/Jj0/Z6nbewUCc3K44j
ek2JKBLQ0CXt64t3Qo2JDBVvpoJDUMX93jk7tcEbcb29HgbW/sX7bHkeDQg7
giKUHj8zur7s+72QD6gg/pnIr9XMSw1PVZXnuQu+t8gew45B1VOAeuD+rMqQ
wYkkXtQuYLHjFE4nxUO9S0VXtP7qUadR9z4UsQxuZKLNI1wEgPZT5EHj8YGt
iJO1ifSxK3QHPqFJMWufhp8/WmpE37Pjedi40v6syYs9ZqphmeqnqceH97jl
TGLqmOwOpg2R7Ps34ybYswYIbK6okw7GMw3Tf7UxvzeqgMbyscq8bR6qbJ8i
zqbqrY/EdrPPgErhbwtt6oTOOtKXXZCoooLYbULDq9Yfh50DPAc22HRR9/G+
W5CLJDytee/FCkBpiuxn1rGM2qbBp8EjsgsU5XDYb64hwnK/xwm5BvOGAVid
SqV28uAdCiXjOsl5ehTSFAUCiwLjj0dBZ0Ntmf5A0zzF3FCe1f99wuN1ykaP
EKSmyrjCukuz+F6kRvT7MMcWkJTw7lUl+GdLkXJp3aSFRHPcdDkOv5UKz3t3
g/ezYD5WOuGhVtBdHWgG1HiaHVoJw3qGeVcTxKFOx1Sc4NeAFyOf8Jem2NZf
1uagdBJtWkELyA6L7PnpyRw3BbRUKxZVg8BTAg8U4hpUZ9i7oa++zPyRkyEP
7LdqMmFKCPojqvO3u0edXrPnkEh0qfjx771i1ks74UxJ2VyNTwih5jPOyeDi
l4oJKnQABlxYiMB1C9NFBI1nCZe3YDqzIUduycRREwffR3nUe1oLFM0iyMTE
GFmxF1ksvRZDP/E7PeYHS+IS5aUKwRd9uO8K0mK4/4Jk7ZXdG8H3WrmsrGHz
Ht7nuvlMlzYf5KrlHn+w+gk0WHdE35VoFWTd3TzWJyEZ1lNyKEKIbdbnw5yw
E2llyi5HSXGsgSDV6HZXQuWwVkqx3DT93sd+OStp58RzMsyNJu9eMV4ZpGRB
pXeg5R1SfTkf3l8UJWT/LHkCdB6Vgoy7b3BjTjHpISuxFkM2zArMznQJEL0e
rRubmMKUI8N7B40FBsfdyeIlqpbJUtOAdOFq4BF4SMshKA0mE3JOTcT5deN7
/6Y7VD49JWQ2mbTRnSdOdtl6xrGkNCLygkj0LpnLpdazj5NJa94CYjq8rRgX
knO72fRW+YSJK/gg1Tc1dKPpxQvyo32koqdIsQAkXyQvtjKmIDT/IEkWp/ng
rAjwmsYAMkd+Y52AiaOipsB7TDP+FcCJrBGJpJ/3isgctVtfitdqKGTuBTOv
9RXpW0vIuAH0Bq6OGsY+1wBxNDr+97ftXsiOR/3Xe7eOiiTaN1vjlRroYszx
jzz6XAhe1ScZCSJ7aVCC42n8UdIC8jU87LnjuEZ2kteJnHOI/tEpATog3u9B
qS94NMV8oRqwauK2Zf/KHLLikRz+RdUBi8zcbRrYrjBagJiJlkc7osNqTgoG
HzbNyoHWT2p+tFqQyINsajL8URUGRjObRlrdp0PEOyvUujrq3zPq15uaEnt0
Sz93XZlljVkHCzm1e/ExuUWEa2CVbvHjCiqnBSRv4Zcj86/ZUdEFVN092L4T
lzOfV2/2Dd6Vp3IEw0dD7uItwio1Uesxk4vpF7rklAFpxVkPVjZhEgbA5g5q
7USzr84mVC+jVJj7RCvy0YWihnnfKLXtMgG8UEqB5DT/d3uT2LLR18ZT3uUn
9kqQxyvs/ZKiukngRUuoVN/XQ3gzx31CgOJZAZGPQcO2STP+SNZo/vK4admx
cwF8AEeKgEJtKAkAWHdtB51wg4/evi0j9uK6uP1MkIT9RBkhqPtetXsLy7z9
rvVvIo2S7gJe9AAL/b07xzbU1Xj6zse0oYZzP+39LcYuee6V9K1ODfFJmIEz
PNU+CTUnBFglM7Jo/hXz+c2D9Xd2RWJ1x7k39kWtqLkgsFY/LcYZdeJyu7zx
K7SgDpLbpPHUJCWPjfXSCybD9bd82XS23bL8lHw0hrxlosNlRawQiEMceXW8
JH+0CFZYr3NSlsE85jvIqaK2WxCpwoIVph9G10m2/1TSow8vFbX2zia5pV1I
D0S8GHSu/zF9gfMwR7/9kJhpMSZvqMwngzyzY5SzOGDIGZQcCczP/npGOTs5
wkI++xybQApd22wz39AxylOxs+11ZH3XI5Er7e0F0jjWGJx1RAOhlUji2HjJ
PCZ3Oay/nyYEEND2b3n6DZtQb9vLkNez399yD95/h2paxQEljzrEO1RzfZo6
ujUz1qfxrXdvMcelgxda3dn28xCRtfnL3GklOqvzZFpWScsCdTm84qEbR8mq
KB2yIxIZziSxoFYl/EUeQrzZNAd5Z6gzwCdzaS0Um9l4dK1JKpoyCXkWpYiP
zMEb0D9Jhe+5gGj2vCaXzitnFyVPa/cEVFU5+0cs/kUM/81Eo/oQtLbiuDA7
d42Kp3GQ+ZXu6nCSY895VtGcmvQB+7j5d2keBCoxxyIX5loHM+PI8yv+LtzR
cCsSw5Pzu4HvE+kcbW0ejn+/a/VKSRt20GJTgsxUT0fS35LRDYaj0XxXMOX2
cOS9W0RK4CZe0/CU8IXkmkssi9HS0vTaNjlFoWeI4nHrTSqZYpByyYadSmqS
bXOwAZkR0yxeUa0S35P8PIPN3ZqIDgvHfA+96LzYy6N49nnPIv0Qu34w0cIv
YkXy/LTfWI2TXZtZubzx/42OfZ8PdwPtgPaazrUsyAr5MuwA0DkEUsdX8VP5
NySBhYUx0g9cMlsiQzUv+HU+d9jm7Dch14wDcaGgR+zK/NEeqOERI056z+bv
K9Nt1vzHxvvPNtKHOesxxYo3e3X1ksLvBi/aKl3BGP42QKWfzm2z0C7/lbev
or23ytzsjkjTswAKtAICv7/7iZMaQyZLfcRMRThRvu7lQxW6aXu1H2ZsLMqa
l2u0fu5Bi/5XFCiKwRZkIx+G7uqo9PogLrjn73aoGrirs4u7D3wVrOHKIqf6
3kK2urw4F9jNE3bVTvaefjEh9ltfgnsSAmgb2Q91tLPkSpX1uLOMmdPhr9oy
toyoupb4ADcpSRPjq8lY+iomwEaC8WZ7KyOhPl9Eu64BQFCY0V3HUU8ocm94
kMSxpDoYkIF4FQnoZz/ZUQTiMYv2/DYdM9S6+kWu4mGWgA7r16lXQJXj68hQ
mFbER03P8XFDqJsepB6TeT7tifhRMsXMj0VPhW0iKtrzrLBTs8bRDhusjTiM
kxavymGIwznOFweld+v+piuG1UGGgA7eDI72qN7euKPGYk+/10ii8g/3e9GV
wg01EikuLy56O7Ad9NfZKZTfkPSCMaOoMNnC+DcNWTjcHgbJTSo3kYYG40c5
EKegzehxZzQw5gO0Vw5VztuN4whGpZVhiQxBly48h6KVVWVxIweHFxtHn3Ha
PLoDtywlNQzzcbr9cuq4SuKmgTNsDVmRTDyNg81yq7JjUz63Bxx6PtDLWYeU
u0rhlLftSggl3PK5jCgh3gTXEiW961P/B6ZD7RFIUuj+yvWEH2aUgze0zPI5
AvKyFFZYMA98qXxq7wvb9FUGC572ajy1mYNTNMAeDHGMUwIc7EWRt60v/fUt
PFQ8banjddtr9XH2ioAq7WsJX9KGwyTOcbCc+2wLPjn5zc6Wcul5PcDE6I5P
LviDzQj67HxlQOavtox0KQE20/1QkklSF73JEqn/CAuS4Ny+sQVWT8RFLymd
gNZVaTU+iy0+p4h48OhWbQZDfvQfNIoknAXCCPu1gPJPkKMDBdYNjzDAPLZ+
IpTdkejT2wNiOnB0nRj1RVQB76pAbmE7nYUI07m9bQYeVmgtZ5D0ROIVkvll
EzcETb21khXFtqNkc+eBxlFWPpfJtH86gNcfNTw84YqXX0gkzEGYYdYZSR0t
RX9KggGZSrEvKEB+lCBWtwjRlsbJX291eV1kdOzAuSucHHWB/EoGhtJmwjLh
rbr+U9GZhjUY8hBmPVeFYGQ/jzWDaCNCulmehRYH7MTS+mva8OICboFobupz
qfGpH/jE9SjUgKYehe3V9p7kOfC1jfIyFbFDVfXpyCRgrme3LO7CGYStZevA
ICablODGZAgTdt35TXbjYrOjpCLuG1C1tNumL1SRDDw2ittDBkzcLp8yB72u
YHPcdKcy8P631nQkZPgCwsjoeK0kN1gPujHZ3TpZdjz4xEO/oqxy5sSDQhFN
Y5gF5YgbWx+spuhooxC8LpWIKXBoCRXCNoaq6Tv1tIqtpErx4n1zMLxLk4RT
tXSPROYQCs2jsRnMhpoBAtxWtRJXBMkpaAlZDIgxxQUzvrtBwfImjbx2CU/I
Op5Ag5ExWObHz96s/wh6QoXnjxfeS2vlaFQHaGdRDr997KIq22dqudwMTxEM
yfp1336iC7TnVNiQM2k6J0STklDmjsPvvbZp0FmWtZNTvydUI83BY3QkR/a7
nmPqgTrmMabfPV1N5W1gbUHunkaFHhy/Xb61hHY0PfY+cAJnEC5OFphyWY86
ixYIg0OA3mwqXlb95SM16ai8jf5YShK8erd7c1c/rHvNCcdedPCXtaLZszXG
Ih6M6RXuUOPO0LOUELdSRdY7p8o8gcCO67k8w5feyZSGyC9XT0566745txQt
zNMmyqYlsSDfJXUQ4Uadf//XN+NkB7YEQ+ISVm3aTE89fodhSD21VgbNqf07
md1sB8rTdndq8dLBdyhZvfckuVfDERv/Ld+4GKK1R4lprBcANsFjpoCqw+yn
7x8gqgEY2Os4k4mT/Z9MuoE7ib3anBy9u+/ezbDQ5OsmVBMMhiVbdzfNpjl1
e1OntXGghhtL8rlGYm9vB+BWVltxTd7AS5V/2/PNNutO+/YzJsj0AL0WUq6O
7tWH2Z1ujj4kG1Z4gZ5CwLBx9LDzsa3GqP3pIpXdVgU9PiZBLSmlquiioAlb
LyULWMLYwFMas9mlwgMVM/3rnbxyCDCXt8vE8pOk8jlCGhAiZQyj7XHgvUF0
ea9ySnnzUc0uKZwFtjOSGTp7WeX3YeHnI3C15NprwZuPJVNiO9NDNlTZz6zZ
MHYY6uO9Kx2RQlbMI+AYKUM1VtslUFcEbzePFepOzEts0XN20N0q4VB+9KNV
jhuQEiKSE4FINPN95lJHfKhW0J7oZdcsQo0Mivb43wra0n+nM2ezdpwbXAld
3OLFf5dGiKX18SZCXZn1Dd2Tn1DasfLbB6MTCbprmZNnxtIRXkA+c5Ir51w0
PX/zPwsL1wqXbEouF3KNqU54GpVKT12mHqh3sVnBoqlnHSU42LvCPe7ZdE1W
V60LaB63mxZ1Fxrd4uP8jb59i1tA3ZhCkg3YHInn8Rv54UJmWquIRt/z97YC
9VK2Ef+g+2SqdAW9UIsRGuaei4HQUMthlG6lX/nPRP5ROMtEYixAPdURqSCs
Os4JPp63Ql6D3hcEi3vgr8nGc5JjdViXtH2vNqfs0rTYezgdp/SyyPYjRdj2
pqyBnwRb/vfANfDtrZbkTDQBT+i06e74bcEuCNmTmgECZ0El811ops29OaV+
5fR6/EOIn8YYKENMKdseyykkFPnFkqXkpf2+Z7rxbbGdAkItJyazBYZrvUUz
XLxAde9HLmeO0eU39U4RQxLb5JOWDBd+ICd7jRoA0xHXJNwAH7RFfvZCJ8q/
MRsXmN+YmAg9pUXiMzKtlU3gu/thVy4HawvtS/yjANItkMGZuqWsXZBXqp/V
TR4ko9k8KGLZacu5+iM2gi9T+GZeU0AeAsF/nN9mm5tVKhgYRwmRAxmH9JfX
7dZn1ltZ9jiV2E2HqIl5uWHAhJxijRVHb8adIV6NSHq9BuPOFU+bEn5weadk
7C8yX4SHIay4Al4rYzs8qd3Fub84yVJSVb653Z1pISUygBOZws70kRes+C8r
sQBr4tVM/z6r44tveh+qmdFweSIB+P0spes9ALN+lbYH0xve9DB+RE4B+WER
UE6lyekybi6NHvdIzkGzXujZnsATFAPzqMm/ry7fWmhy8yVD8LIQVB6TUHvP
k/NMSAiZkjfWnY2NvqDgrv9CETfyE89/Gdcb1LsWbCJ2YQHgDo+iDqAJM8L2
5Jmb9sMjajt9R2Vn1d/pkp6kX50eZ+G05MM5jrYHrFNYtX5QL3KH10eyyuGX
GbhqmqraK0rdwrlFm8g49a37gWCF/KHvPTROLv6ziHzPbCDpe2S83psGXB8r
pdCXomzGNqqEbaW2ozc+7b7Ul5U2BIVBCOmXTGkXGMxBFXXIXIPU+TQJEl/3
pWBZtQeI0Fa/4R/wV9vyfCR73um60T1mmjAdTEtOZ9hw0ttIpm9IR/Q66zfH
486OXq7UI74eVxQYNrkgLOMG/kR+vk7i3VU7KCUJF2Oxk3L7aKmqenoCFjfN
GYLGxLEla4pLDnZ53qdbq/IDYw/VsIEaV5Fm134j7AV6w63ujhsi+PI22sXR
vh5YRpwiHUt+xYTKzwpOKg+rknh/4Y+XV/djl3axeN+V3vhgF8tglzq+rMdr
ttzc0dpChP11vbgYI3TArOqc1NayI+Usw2cFUEb3arNF3hYuCTahZWKrNzSY
SS4FYb9pRABG28p45O9/v5sKAA/TrS/LSH2uhmbSvY1OsNnUSBQ8fz2CQuqE
IGaWYqEBLClWARnKXuoqvms7uZRAxGUzddBFos7n6lZ1FUt/KEqR5EzyrUcP
HbCj5Jy1IbK/HpzERcgVgEiQYcDmwO6Ky9PDr43r55TVT3X04ma6k7HpeDCv
nYKIaj1aAZKsw91noz2GxgUfpySgcZzmRVkHaDjrw9mI+cN0nVDI24x1unoZ
O6kcKp+DTJj4ZDuRcy1bQJA8fR2Awg6yzZ/uxjvRXyzJgs1Gri56J7YZvWfl
R2pGSjim0UIgtTQUz4M8e8K9zVsUzTSMnCWvFfP79ahb2lBF7XCgg9K0UcYw
3pojaEMbJNYeph8EVHemih4pXEAauFzvaM6CvbZf9Z00u+CSKuKzQahTpYmh
WtiMwWtck7vxmkCKsMou3Pc6DLFVoxC+wvLkKDNBYE0foeEFzrfwEUQkny2h
PV2ekokyBoq88ya2/hODnhbK2vufBJ2xlFS1Aye9vMnnth6RLNEv+0whrH91
qJMXXT1G4P2FPERwXxfFzzAKenF3E8FUaz9TxWH067nW17Gh7j5EX1l2IM2J
Jf8jOVczeDG4fb2zfqYU9cdXAyQfutKfdZdfGVnPOJINC2N2CtfXSWGORogx
Zkbss3lOYh11bfKMB73uY+fRjiUhjvTULtgpCmrYMLHf5jh6FNO0HWlhgg0J
xnZBCQvzeq/Pi6ksMgzC5rH6ySi+7XqMPG7Dc6jPKyz63m+CsM5KueHx3AOF
a+NutfsigCqhP9CQaciHbLufLVh1NQ7fEZlmDdnvu60Y9VtOJrfhJ9PEzsuP
4cH2vV/WPbx5CluUrwnqKA+HZPR5vH39i4jsnkms7S2P7QjPX1UdW7KlZ37J
Ap1COKRQJ/LqnDBNSM6SOHYjS/udGXOE8fGCVXqt82eHSubfOCcVo55e0ZZ5
MMRCbEV211yaCA7VpSWHiQZxObturG1RUE02d93wSu+ennb9unj3o+eyPALt
h7TZlf2u/UmMANIfs6SeNWNmxZGCbFIGlBj0/mmVhkQ+IFteg/hAzvBSm7mt
AewuoyTTMgPHEOgKp7MsKnYmapj7/Tba9Vy0K5s/2KDTVkDl2nFeSWBk5gXb
AhxDYpzStZL5m5xJFn2bmQfod9XZxl9nNqcmg1+C1G7/MSdgRYI0qkqVYtSf
Rv+7uJmbupezvgE8jWS2oAjaTsoDBs5FyNKTSwXYz8IgKjHQfpRAdxxg0QVP
qGDBKtX4ySchNAYnqdzdoS3e3uzLe98mUOth9OnIyIu3CWe+D/divK/EOW2s
w7Jk04QTNUFoErTfpx8izDj+7YyO29o+ST9+Jpv+DQpA/dCiwpWkJUHH/our
hc3UnTZUrPW4c/o+/s26tHp5LVCax2bCFNh++I5dHIvYE7FqV3l4QzYUnq54
G1wGRLDz7s1yHRJIqDNdsoRNNc+h3WHk3mcoBmm+ybDyMK/vx+PsI40wRtnS
AiY8cIaEzWw1fGnCNccoyOdHbRSpE2Lu0HocriCBkxswE3AG4GkTNgknp28I
tXicC4XBcLoiMpI3eNNkrtn3SHK01c0yQ5eT9YPKG5fj/uFieg2fmOg5GvmA
07Ng5RD07W5rX/EhHXyxvXs4lIKzVF4rwxan4K2doWIUOlYtPUVCJ70Dnz5T
dBxePHi6qOvzss5EGEwPQj2j/sjUskTCP12wHPLsuUkQ9vDETLmb/rHZJkP/
+cJC6QBNawIflbxxSbFthh6iGpRhm+qn/R5LRWZTgoqxmBgrjA9JqHICo1s5
SR/C4M4bkig8XVcZVaEhjSkJxbx9eNkGg7E/96ovn5AWQIprukc86/Q4qU5e
2I88+f/ZOh0j75wbW4WLet5DEYEV08yTWjqY77aSaYjvB/Q0tLRJApjrvqjW
dtkkqlDNRNOAEr+yn4O6To4Y+rcYt9hQlxocE0cnW2WT+/Uv6OSqR95+fttZ
QtmlhLP7L3xRhEChlYTgvcMnwKXP8BDOcK4zZKysv5k21qMlQwPmI/gDDey2
PA/AwM73p4bbRdc70IN8bhWHyW6yvGuFWNJ6urzSjyTSt/Lt0dpCFRO4hZ/5
y55Db6zTE3JbRMc2cEUSZFJXG2uuFXu/NfE4MomA3yjT0qi6FmeGAd5xYSJA
GE7yEYRf2rGbK/uHWuBPlAgAc0E0xKfMyL4e0sXJxEfZfsW7EdTqrVtKxeIx
DVGEML+Mg+6SEnfPvM9GcrAz7RBSyRERkINgXVQxk7FF4QQY66Tb9XkdCjo0
2UxrZ+T9y8MKIbtcUOd6Jlc1ONCLHZHNfdDHGGyQ4MHqykCqRICsLOlNqJ02
xYZuywvl0bnWOXHdykkKLqyUKpG+9TylBKeumb8x6QhjBgylgH9ZAgSOB4W1
1UjFFbUmoQQ3KmqyYZIPeTOCwpFrVnnJgpWD7Uwukd2GDJcD+QOFdwpUgDb2
S2AkSY+jk5F157RpiohZkF2zgxoO8Kv+RuQgqzQ+g6GuFyO0iF4lhAmI3YLv
Uh9B66Z7YL+KqgDfh+EkOMfzOq6LRvYJsMb5I1811OiqBweTkwVOoBF6rvuG
aPoKdC8ZAcZ+0TrKW6Bc6mGK+SZrGzMoI9yagWC7Nn58TUrglCrOqMKu2dYO
WPqzBgQWwo5XBC9osssW22MBJAbGY5VLlmT340o908+W7GFh9xuQaHCOiO2s
HMwJ6MJvg+g+wQbL/M2Ofgnf0KvVeoAGyol0q3Iir5wVDEdowGeix6rEp0g4
l5Q3QBywbgdUnnEQ6aOguF6MSBk+ctVJjALbt2NMyCZOYMhDlqKZW24BZtHH
3XkrVjP7smvEdlOXtmTbm6MJoqpX8aGjN+b8llx1VWhg7YGbT6b/RE5TSBWx
JJjoUbsFsZCpc4kM9nYYFojET9cbgRSDSVYwce6IT919YZu5PPMHrtofm6Md
eftOLz0J8DvyddyLeiRCSsKA3Jk0L9ZULsGBTqE9tZZC/NU/GHhrxSPjY1/+
yKruQP1O9OALvHG90r8VL147FDnD1BVG8eV8Ix9LVxR9estcj57du088q63C
kNIqteLw5zvHM9j0PgFdqpIdp7az89FAWDKWBN3g9AQeNefojoLfeO2SHIdl
oaGoO8k9cBZkA4cC14+uBl/+7+wRk+qFVUA+dsXbApUHsknegaEJ1mQ119WQ
uILqdBtftVGjRc4KlgxIut/O9RBEEmZhWda0GvQEmHKn9ypww3uxlMPV9vN2
mGVQWyLXsiic4bBN8jWC+viyvPiVm+oi9mEORvx1s+Hhvx2pKKgnTROFTnON
w83XowrDXN9j6qPWK8lf/nBCmyXTTciUd8NPf/0JbhCdaqjEkQQSgh9VCb+I
0HD4WX/Gr8731D6IfSfC3KifGv2PTv+7I43euSeSvrDAA14wQkj8HDfiWVdB
BUFCcfb91i33kKpfHyDGkh9V3JD9n1MXRWy3wghw/hOwdLrP7oohV34ziCj/
fy5bSwQchdeuekOsRlsRRAL7UiIYKblO/yBnOnr6prXMyqhn1p62cOkwWnGP
1s3twRBVlm0G9zTXYcI2sUqsRoLCzz80A9EL5KNrKvGQkAVM3kK/lJOT1MXk
7lgdztrAgLttNtVdY+a+eiQZ57rb1bUi+SZgMwxFnpd4frfHghvyjfA5Ub61
dhl6JKyHmkuF3RHmOTl39YdVeChaKWa2HlsLV5MW/0+uyPRoqG6k+XpjjwNr
Oi2mqs8pCyVOb2yBjG7z/3z841/ED2QKUjoMc+iMcqS2MhPFRJxkbz6JnsjP
soCiOCpOHd6kDRR4PfgjTWQmmMK2RY7dBJ3FjT+r3or20BbY9DoXlx7XcY/t
qB7IaHU8ZJkVZxiIAvTP6QkuWfMEQUnSfhljNk/IisZAn+g/I7Fif6/mkbT/
UIxQgXK/VfbePEu60Tu4XvvnLrjoxw9Ut7zfDOIHiLEUfDCdZ8t1ZNJWPPqb
SX/wTUqaLN+1wuhYIlXhowtrApoa3TBZFNzyBNXX1jYXFKTs7QxNULNBehJ1
Ka9yIpH114B5b8JNL1uK7rtDpc0+vNwWFqQp8+YnRVcgkdw3wS2OH2KqdPMH
hPdSz2a66SMEZdIJfh4P2EIBpXiO47Fgz0Evh0dIi9UBhQYG1/y+pfHkxV0O
pftrB+f9Z9TI8PYKyIibfGVWsDKUlc0Vl0vHL4NMvRjR5sbWVcGrrxtgmVeA
5/FagESSJ5u6MpI2fEiSq3yJqfQAgg/favOAr/OCYmjaqyD09ITAWkuGYZ/m
879eRonlMWmClv4vwjx3L0XfmcLJW8L09xwIrC9fy7AItGKsk26t1rELmG1J
ydLB5PKdrb7ctRqWvqpI545TWAEp+uEn+MLle3Q2rlsmTyh5+1cNb/UydGf6
Ss6ygQ2DYDE0qmtTeNIeS/paff2D/IiZIzAYbuTK4frS7zkAMNqG+I4W54Cu
3BRJgM7/W04/ToyahPOw0UptdRLdvwIEMJh7Q7lqJpMPuBM6MIiy4wNY+O4t
eQ/ln0gyRHnSrcpoDhFf7h6P0qedzNZegv/YQgio1jLF8uqNxeLQ/qS1WdSS
bXkkqun4Q6Z4noLdtseE4HWi5uP1KT0zaWrtcnfSolI38z7BlSdTiDWlqwRE
1wzJT0C3bp7lIPi5A5ul96kCf/FJtdOBuOmREIFOk5h2eXyMi27fdf1WCR3q
gZtENxj/G7QF3boM8X27BoIQo4jmNuyWW7C0Ql7yf6WywQJxBEqk7iZyVryb
09YgJbBUR+aXVoT+ysksgzD75nxyVgYCdlULRoiMhT1Eoy3lWPnvaXdtbQOu
a5NExoTvafNsfrd2H08oWWONZgE5/WpBePUMaZyLpGze8/yc/FY/oFExswWZ
/ix5ytT+xai0v16202PBgnK6e8/RidFBMSWshkucvkIr8Y4HAaKvuZZXpISl
Z3HWopizXO3SlLBW8rkzk1lcaMf37VUMyBl8ULYsyNVU0q0Ids9v6zI/T2tK
V1YBlIFoEcVpFA3ZPiQVrTvjKRBJf9QeoomeUS9OIzk/5Eoh2rOKqTC6eHAG
vxu16z8B2CkJIoMkttHWjROVY+9ihSD/thUTXZ++Bk9IDRd7R/njK8wV0Ela
E0a9bhzd8yIem4TPdHaHtNQzyIcntlhd+sWhfK61+/DA0pm+HwBGkL/xPdhq
0TkD4RxsckXa+HX/X7Qdm5tPG3GAOX3hUrfqJdLuK2elTi+qm7TgZWtEV0yt
/5yXleKmxRWj3HoCgLF7L4i6+Z7J9uCEU+91VSmyZvfUGzHLaTgZ3vXGyL59
TlTJFU2Zn29uzNMh50adb+iQpi3OyJSaZW+z/UKEE7uro1rSYFOYCVDdyIvb
O/ZGOvkbObbt7Q1HE0pVwnF8UqcVu0AMpchifQUqB3cCNq2TqXi2mOMopYnv
7abh8VUxdFa1k/i4Aad3zP6t7XzP2QHGLUE4w8rKiWYiUmJ+4j2CrRVHTgXs
ZFjLSgsP7GEmOnsJ6C4OyMMHQBNsZezEGS9g+c05M2MUpWhJM7w/OSGzXDbb
dhglRp7zDqU1JxtRx3ViQ6O2ukkuFzjiDx7votJVmkKSi99gqqRpYIYotj6e
kN6rOBN/H0b7NgIk1LhPLsYmI0dDv5Ac2CvKSIQCCpSnaEM+QH1aSv7BWZO7
KGcdErM5i6YD/+1jQQpmmdBSiX1OSpypp/atNQLsgOnI3oSBOiAARVOi3pgZ
nvBjNWCFWrtn85TS9Fzg7MevPMoKLP+eGs6QEXMui3hnuj2VB2s9BWkx9/VD
ZhZDvu+ZpazWza40Tv/u3o/2ZmYA6+RJPpIF6CLJswCgU64MmGUgAwG6B9Zk
jJHz/TnAsZnGgPt6grDyAleZhr+UoRfik/Aks/QAYQoTzH12LNtuTK8ZvnV5
7B7dgdR+Jd39ucFKY6++3J5kpbGKkDKvqujHMN2A97sYozhdPatbEMhf6Rjp
+NrZp5uxor9kVYblU0Wx4leTLhkxKyCqEkUZFt2JdYP3yt83sUbOC6739pA/
jmY5Eg8iCRkxzAbVHwVYVonIk+NpgsMeQLzqOIdMedkX6hQP5ga+K92WN7za
p/G7wLKHJQ9xtckJCdwa31PvszsSfX9a71ndxLgrAItB5lxzk/E3M2G3DMbx
N+0wRPnr6wkSrlUGZPFAfGSGZhzNFv3DBP7gAMiCcbh4q6NIYec2JEgCrhpr
fm9bMObO1Kp72C1qcgm8GtbpObtcESCS4Yf/70Yxfqx8acC8YeuWZSGjubhf
okVp8p0g8OBa+np50CPPge4+1NJsNUq/bGSTC4fTZuv9PVbXb7pau6pnmHiE
DVs1H+ATDWu5J/2zsSNhS1NyyW1BR4TcVwJwkqXr4gsVQgUrFJRFxTSpU40e
yuc3XAhaZ/PwinPy+kGMiQkc8+pFnGY8QMq+wify7wCGfG8xykMBNc3fX3pu
yFVw+t4dRJEVko+NGJTpAXFESu6VnMEfq0UgT5sgkc6rjPS3ZLL/ek891QPc
9+TB+kBw99FogDYW8ItYj/p3YhEbcrAASfG7ArlczRMvihPwARlP6eaBaqTu
s8nC7qASK6VNF9pc9YuIHs/dwNEpw2QlsdRK+FUhiPWNSTK2yEpcVLPrY/5j
7y3oS6Kiv+NOqyIVHkej7ng+PXUjVLARG2Vo+H/pJnpNISCdhWIHSrVJWGSP
pgSnK86Work2qOxxX47W6pbzkez9r9jizrBUMVRQulufPaMLwVuOywR5Jva4
iZnIZI5rDgEktP5cRxUE27Ts4FlQh9fuqXK4Bv13oOwXc39P0MlGB1H+2tEY
OH1XrJEzx00UxHaRCGP3V/ulUGyIEMHvAogYO1NhJVHK8QMn4mI7TE1FODcz
B8YDzJFuX4/BZ3eJ/NgFsuSVVi04wvp+AAsNyiwR3I4Vj4fk5BJ7Q4CodxT3
NGyT1+w4ZYwWksr4FhShKULiGpFf7WJHGg1E3rDDF3gmwszRI02M2PqAY5MA
X7nYuT/YfLZDQW3wc01klIZC+PaUp7NcmNUpUy0CZh5hE4BOWscvSPdejH7G
UyDI1QzW7D/Oni/rAaH/W4AW0UoBBcQnZ9NUQbXRnZppsK2jqhI3rHTxG0NK
BQPTenPZA5I/GPeKvl9Yjxan9/rbw8WaBIXyWaNEvPKX5nXcYzhTjBWFV2WM
V+njcapLCckH4uHlDcyj1VnF2/8f+C7vrovZd+RnDijlgPdRDOQMmgjioAoa
xrkoUxm4PW3d67iXv9EC/uLiLzkqGR0yZZWwTEQ87fDTC958MD8h81h8neuC
K4czoXMRG9wPJbKwmeRcCA4hjomaFTbJ3FOoEH0KPGLrkoHN+8rjL5SkLIqN
FmYN5b5I8wMxTNuCwPgs+CC0mX4DjVcbtyhzkiz0XNI4jqaExwLJeIiLPsdO
/RId7xjhS/DDcvghRSVNhN+MhH1/+GLwxZbYn9FD72YZremVVZ6NI1txRrWU
m9FtGXKNADAMFPQT4i6uKtvgVN7edchsM/xBSVtS+0qoj7oY6lx3T01r2GxO
+bRZ894rh7EJ1UKIJrcxZ3QJTzPWC0jyMyPdCMOt7Gh1GkEZLqeYgTUVQ7ns
7dpoNoHRggClJdpl0ldo2vzlcpiEv9DLQwmEQmUufXxxTbi3kUkmjkjSAXL/
1qiJJly0Cpn2FNc4gipVinhr7tw82sdreTQYmjvKfxzACLGx9jqTLUdos96c
YXCVtEulsx2dNq9MoniV7AAZAMuEIBqD3yM9+r9J4ryA1UzyNxJoPU99uEa2
YncIFzNZwdtprBXy1EO1OWN06poCBN4Dw0OFiRyuiRAJqB/MpdYp6SQWy94z
UhXMMsNmqC5uMgMm2WnU+EaTbAsG9hYomKMQEsmJK4WXWEVFSqmM3rVEB9zQ
KLv/QS5/u8ncArH7WmxL82NypXudODLVNbFlu6W2KmzilYFr9J7tVFtr4SDE
dQpxoDqc7NmAbHqUvJCFZVHXWt8o34LqIrsDHCJgyLhSrmf23KnVMFB7EFFM
asb/gZ25+SM+p8dcQqQvp1ggQeJ17HNdjTtsOaDgG8LGSm2GelyQ3IczYtNP
D8auY/RvqtvXWycT/lZdCb/UBH8i2BM8IszpCNgr5R956XrIXwBqrvFqEBHk
JFdeg9DEhH6X/bb2lBH4CsxWYWlnMTdtQ5pfI3l441F6TEAJ0tS4Yss552xn
fWJsYrWUZDPpKEGwEMl0tsslepRQLlPl5RAH5WY5qzMdSQkTjcoyJZcwMVmN
Puk7lg8jFtUpKcOUfuXfZMj96F+lIgbmcSsQkNYxq9JAan+YmLe0w3gq6pLA
rXUulXDol5wNWcrfCRtHu8szMuro9hJmOXSHW0pbjR48x5dhNU9B5lKhRFTJ
DtUUaRuKuNgj8K2R1UhjZzr6/QHNGAQ05LML17wk3redJpBAT+0ycuMKwjrQ
zpSQt+NbBG6ZInJtgYYB9Bg9BKDkAE0UKCjmmFprqhTpg8Vn7due1mWRwsQp
pw+p2tjI/VaRC6WNt7gFZ+RBEpNZiQuJ7DWDfOGfmLk1hyp+AYkaIUjQCDYV
2M4knVQ7yoZGMdT4ddB3oKKAldi7c5kiHxznmotvKH8lW0z8c/qG/KMUewp3
IkR7yJKA/R52sRlMLeMsxo8/fLIt9KAvlMq+fsUAZoOqHo3qhVYLUGp4mbz1
5euCkbBGhhawxMUHnAAFoxTHYYed1RJwShTcZ1TxJ++nWJohRvYxuWnYVxos
pSDd60nz+40AcUYKA4jDbmZeRW6tU8joFfIDC6XoliMBUAOPBidGviVdr11u
r4v7G7ugDwViAkq9ej20l7AALkleF7nz9mOyy+Vn5DZpDpRoU95Dl0vxBxya
Ys30UdTokcZ0fk4xZAwwDDm0HTv4hvtf91vff9aOOlBhUnFK67Q65IYym57F
hl52Zyw0PfW0pK/q7/VAP47PRjtLwl8RNajpAp6T/RKPy0FGFfjsNYFTKJoq
z/UAW7f7rwFKTY6uC4RKwfyt6bVv8b9Mx0glnRPTJ/sx9matb4TBlGghC6u7
8wnorq0J7Rk7qYa/cU6cmmkceulFgCztH7vYQNyUZXfu3kw7aR56qxiHwqHw
p75g287/w4ZT0wEwMqw/DtYfa8w6+7hTYffLZDo7kJTq7qVP/riSzxFQQbj1
VDJECIeSdfWf1rKNubCtq71aNeJGwr5VsbB0Q9ZtynsProZHwpmwAnLnq+Kt
hADyoOUnwBXL8HOsvtR8ABFio45bkXv6vFquglTbgycbV/jTsMOTuU0UqcO6
R2p6dzLqoM2tgQ+etraDKKm3OBCC+z8RGLm+OjvC5WKHSxtHHYba+KA+c8z2
uvw3HPCrCloULrKnUtwTucpSalUkRB9PpKi6aJ2T8rh9vV6aiXnLdrNsqWHh
0wgX4dL6BMdHkJUJj6YonL376DrhAY16vcs3Srk+axSflVVdCofm933GQzxx
YoXN0CSZQ0pxKDHhTxpvCNij6XZ7QEzo/0L/pruyCm6JPjVqtKSFsSrfdxjX
C8zAktXwBbfhtH4prmjVDWi3ZCx9aISpmy1/oV2gq9pdqN9FAdeT8oQU+dJq
VXbbFTHEiSJwlF1sT8raM6kL3IHJG6hVcvt9oyZsTyqLVT3uVKv5ytVpYJdn
gbzb9yyJQPGmJ3hZMsbJJpwhxD0YEl3BTvgOKMT6B+WrKzvLmGrqefDZYaOG
Gxd06zhFk4Jw2zgG5dUYUj1erohjLcPAHHEJq48nwCidkEoAWPpKY9+U/DDG
VDxsHnaDGQJ/DbLaI+OoLfu3e+7XaWJcvoGW/SOU2PYe0dAQsNrVR+avubdx
tB2YWf1EEXalJDV+Gb9apUGOfe3WFuuL1X7lIL3SAMQgeozSAT2NzIGsRTcf
HgbUHOZMTyXpthnqSUGedt6FG2OYXHbJNTos32vqGasn9+txVPplI+uX4oRq
yp/qTVxC/yQvRoAF2FEcom9ZPjnfGS+hJhzH621g7a1M/V0vpZui0Aarz/VO
RbjTvP59A3YK1MC/OPlOA8BZmW6QAA7MOYjmbp77xWx8vV3qPwXl5w6V64K8
woGOsWgreVgNV4HTc0xLRxMW51giwCBRkY7LLQkQnJP0v3wNQ1LPQ5dsFxLM
HNPKQWIq+2yCt0T70e+7hwBBOx+4+lmYfN34HOmfrD2Nxdda0vy91b3BY3Lu
cwugytVvLzz0ja1UdH9TVWLE/TK02vE0apcv1Bf3k9mL5vtLzeFyXicjEn3j
S4hjfcu9vyOYjF4Bxt/161Q3KwuoBx+2kOEor0gvaCOVBB+iscREK1NG9um+
Evn8uaIA/gu7vWMkYPhSzRuA4Ttkhqm8LDGez0OEwcDuiMjfc+SnSNZUaWia
zT/Y5YjY3X8CfpdW+aSzd4jqY2hfa3gizgSkMhCg89XwkJFX7dEvDDdRJfAe
GaxGuGFXmUKc99KfEv4hQQhGR99JvyvjUdXKTeE7blAzQ+6/Zs101T4q9WxR
UThglH7cgY/WiNwL2MYudovaxEKgO2yBxahPXkEyssBiLerTkDJkSQ8fZOty
I5GcHY3cguP1lon2ACwFHLKujW5Mqx8hToFxb92g7ql9FUPYVqoKHAnBe8RB
ONBfL9+xJO2IjX+8os7N2Cb2xFTVqkAJkWA4p3bD8p/2ErLsYWKW54QtNb2i
HrQsWsR2mhojwCUQ/WQ5+OC5T2ZYvQdEZYld9Jq3nHe0tCQNdBCwZSP6jzAN
7iZehW0Em0los9ObmssetwiT6Y0mW0mNotqoxdgtsdeoxtQzk321CyIqRr3y
yZ8AhXHNnnlpeNWj7B7L1qmnKhb9Kpd+ZErc9ahhE3wqgjoJHzECpxHHGgvS
mI0JMrJvJrrndrAgk2zAXPnJ8JRz2/auIPJeubNFvrrQuAWSbYOchzvECtpk
Z1npYVHgzuRpr6r5uRedwmNJn4ZvA6wrTxbA4YTmBAU3I7eMoOg1hu/DsSjg
JpicjfZlOacuCpPPq8V2f6dF2lAzJvlLFfM2osFKIc0h8BqlOBUtsC8yKFcq
/V+UtYIZed0Q6FIK8yghH9lr2CI7RcLmC6BujADDkCGeSAa5J5R7G8KiqCj4
HM1AxNjQ9VNc+HJ4HodbH4JTVTJLl7+qmNut3T+GSNTwsuGmnzx5R9eRm1tH
7HS539pfD/LmYUVuEv8HvAL+3+b5a5zv8twBP5r+ADzjYY8awZAcQSDWoBqN
eHHuzYy615Uc9Ls61+kl/YB70yke1/D5U2oV39uDb8RKzwVtDUsaZ3ilGhRE
f9l3jgI928x2J3vQEjxI5prfI31dnAig5vfNy3gQi/IavRGPZFmkKQqH7ciQ
RDzHsx7Sl6aq9Qsv8NX1zi43RpBC7bL2l/PnrmyB+IYYaSufKxkl50VT+uPd
0u56zaEPw8FvZFPL0CopJONVpjth0UnnH/Dvj9h+1NyzpU27BjIqrSDCSffs
Fu4OxVS2Q8PgkhPlnm0Hxh1KyUQxhmVzMMBJrzbvuW2X+LzwuC4/8Mljfd7Z
rfYn7uNhoPfiZhtFRkYk9jAM3I1r4+sXrrsSCRxuYEOCfqvJHH9ewY8anFcz
JXyBbrcl7TE3ZgKTURlC2zEofr8pdCxey9QQax/ionFvJPjaJ/RLM6IL/goK
2su1eqfY5cJpkotClFBd1krtKhSsDcEdOenIxtHK7/k6EWqLEZlOpPuWNPqo
1PEbO5I92olCwE5Xq/Bc5P9+vG92VqXX4do2uwgFnC6DIq8w7EIcUfzJYGlh
zH8yZHaEGbmp9GtkXTZ0nUIHzZioLubLsf3vQZUFGQr97V9Xo3GZ/uuwLu7j
PFiqEu5nXH6x5y8ClRmv2hlhbtuyYg18iWHXavC6uBbHUJPCR6J+RrNgewB0
mOXctt0RoPBDEjVH2dyc04MNcy5yzaH+HVctVBVucVksvBKd9cFu8EUpoN/q
UnwtOZaScyHyrcpyUxrQUcNRUhMqWjwzlCStDnozDRKyD3wnx7+QLHMY75MU
sg/CSe6Yg9t+TNUgbgR8NDsJaKomoR/wLXt83UtgGL4bxLjzFwJonOn0wH/C
9SfqjqNC60L9haBpWPVfW2nOK0bPcp2RqZmLmKtXrBEafK/Y2AZGGfyp1OYS
wtnu7quoa8r6jpIuPj1SocQFqAYapGLUEDM8bKuzzAea7yT7Ysrj4wfAa5tC
MDLsjXwybyiCxcaXeMUZtp/6yZZUJ6kbqmUcMgRRfUiRdRN1CSIwn2/CBoKp
rpVrHklA+9fBxNPXwur1wJbJDf0BMvsaKuqHyrfgBkYVhe4IEPk4ccSNIfLs
QbNvfWpeTdsgfDHGSRgQ5V7tGEtmpVlxL2plcsH89AaZdxiaDuBsAdAm8HPO
1NhrNYpmQFHqyyhIo0YFqr/OXASBM2GI2reUDK+pltH/f3CiS8Ghqk4UTEUx
lcCdhHx6Ib39K7mUK2hNbgOF2jt/ygygFfFNZwHKnYjWMJ/oI4TPIbDMaVFP
PFFYMaCQ9SS7gqiWuT4uTIHZlP++MsrSIvCG7aFk55EzGgeAvsJ0iud/z+NA
P2xREJSXnu3kDhfnWH4mF86iial0Yfcm5+E7YHcfpE3bSeWQUCmZygpTy5mT
OC30HOhMOgJFpQF7w1pQY7J7iH4q2KWdaNlm0RAOWtQEStiGJkN1nv5lOngn
OriU0OZI+6NZNIOIosgg+gJ0S56JeHthyFT3UePmgOL8ufe9Tfd0g0bPJTJ8
IC78hYoEnC5M0p2x6ABz7mG7VUJh3RqXAtwwvHO0/HMK92TRcnwd25OzKuJh
/GMbs6wITvNWXtGbBHjTHUcsjgDbOuADAfr9qJmhU1pkehn0etfMlFS9Iukl
1jfPUzeUvotDDPt4jOzIVWYn9eK8JD/zkFT98cpWG9zgfJ+/16Hbi/fC9DSH
4sQZR7D6fM8mOVv35oaSaRb253NVELfJ1EZ4WRuDkJRTcp00Escx3IxhWXln
t42P2NCxGU6AvGOhGQ3wkgy+t19nEUKF+xDXKyqhRrZioZrgPODio0Crs+TC
Ya5+eEinZHMlSlO5LagwFVCifMwoi9jExVYbvG0o1P3mOzwLlX5wn8j/XUDs
nn+64KWSgW9Tlv3LR6gJy8nUZtwqNagSVRaT4vWoAgxMjz9GiTQNVJoYd3rP
1XOZnBtB/aez6uVoX/rswSW7AVdWanl3HTIq+1IRvpBPcxXWAIqPK/6zNhwI
hoDAYUhdr7Ts6lQlwGKizpagItQ3dgbsO5HOZMVBN8L9CsuQoSePLvuWEaRY
hMehuqsKXk/HnUkfpvuwEELUhlKZd5qe0YtYyndyLVoIjI+LW3EjZ59Z3Zty
k2dCkLWlDy4AOUsEwEc7yTM+Wq+UcKzFZFFwDf8be3T5oJNVJPtnLZ+wLhJw
j0Oar/MPPNfGQuR5vNSnuiTtDv+tOBc+EBN2kRnsSOGBXGoPI22fLEkPn+oX
Mo/7zGNY7/ZHb9773OcT7U5MKXMB1lQ9I7GpDH56+/jera2+wF0Jp0gS3/Ju
FvZrSsG1UDBZZ/OtKrJAh6PyFrLvi5Ha9+j+gvXz9gF9zhx+38Z5hN+MZ52Q
m1x7mqEPBW7bkMImUez+2ZZvZwzTcaavZP30e/MLuolXnV8Q5OgFfeOc1O6P
mudZ+6bKZPIVthhAVOlG+bt+5VCIC4vH/bGGFdATYQmbxePgpZm4JDYUuUWs
nt/1YMOIYVGOi1y28n78EGq3DxIOSLykmL2Bu2GmBW/pDCBLw1jBqD8xHsK8
SPMBKQtp2euQw9pEILzUTFSGUdalvzcoHp/5hm9TMwNvGDPwAITu6bgIWQNh
3Dj+yMJ9aAQ6Q0NMa+gzElrV593VgZ5urElfnHkSAN3XpRZ4+1VgZYTTtJ8m
1ro/Vzei4ykJ6WT6/7CnhFLV2L83EKfp5QM6YuqaNLQCRPCbNGzhWdHAA4w5
FQnYMp9bwsXRVw4eHbTLIxSAs9DX3TwRfBB7BWdJcmFPBHlc0HaBLVXHl+Rd
JXUcswjAVwkg/b1D3qJQZstNADMYsyAzL4PZGcpNqCVdJCFGq70yAkoHJEfc
CnaI7rOin7/nR88k23qjAfDDXWGi+5lb4dMpLYAi0yhPRMMKirQ84EURMeIc
B/5IzAGkfogyFDPDsdJyTTKjHPk/SuNMZ9w1F6vrqmwdg8akmZGw2u/97/CD
rvqskEJxtVK2YiqXkqaT5rdc22JtKBKFro7Ri6gf+w86uUlNZ+AWa8x40w56
YpLmXdMrMwnI25HJJLZEQLGWvieT7IGwT67/fUH+84HqegEooWjfHWhgwFX8
ZPKVxB+SuPhqY89nKPPmZKhswSFVllrVNns+ab3BA3gafTDgf36GItxNS3ru
YOcMGqofDNwR27Y+jMgIKH//mH3CvoqFFmmGMp0of+LqihIb7FM1BsABXcKp
sCsQiwy/1yM2ViXNPmpn0CHFA9ANjyTOmjzcggiQrWYFVSzF+v0Umc2SC6a2
Ed1YJBvz5Q2NidnpSKQ9wo2mYRF0tyMte5imsZ9/EhH586bxRqA+IjvIOZ0g
Z9eaaUehdjyjku91AJYaEd0gct35MtjP4jDsVahDgHJiTuL3uKj4oqWfCf5s
z41/07S41tE0+ug2T5T3j2QwN3LA8YOizWlzCseLkzfqIbx/ekgKqOhfhlnE
dEGQL7D/Iil4jayio7Zu72fVnQjGovS5W/e546xppeJWKdBps8ul46FBsLA5
VWUrUAj8Jm3R9R2BFpjTC93QpSzDhB5ANhMNNO127HMF3U9+uLf/Q4GE5kn0
qNS/F59DqfCGlBn8N5SOuKggpyQJwcxbgTWhiyLcoopag683LI0Qqk7H4Hht
cW0RzxsC7JzaoaTHEYuSlI4wpKc+Dbn/RGpMwfTpQteKM/MRNh/3i0TAnOoW
gvm9wiqtReanYN0qR5FXV0Wf+EuJCVnYVeM2z8VTF3MAWPC7QabEgoJXhnCd
QB6DI6V40t8+h8Z7XagMmK3QYhb/+Z20OLyQmcfdbc5rYPO38k2Hz+BiEcv+
kNQSc3nnixDnQWkbwBhZODrMxdcz642rkFmxbHYU7cR2uGxz01Bcq+OrOfgE
+AEin/jdzrpk5H0TBYWE0WxnnCGEq0gTc1eWTwwOfI7H2Zsr+r0aP2j1hVjL
6FlAT3u4Wu/LkvnHdFdOWvEOARwmySpmC93L1JzdX48JlWbufPJ0R7JEnJ2S
B9uRlEmfhgPHCps7wxUZBXa+I4J6MH9pc1XLv9mMuDtKf/Wgk8LsanGVgfp0
QvSIMAPEWeW/2PnPLMDwWOSc/XTzauHwsUTK/eFOJldH+m29OVzilU3o5qss
k6w42lU2diTesfDdDc80ScA3oX02lfqSigo5ED8xF3W7mmiE4U8CbeWFA8Y5
5eOn38ttmTlybLl8ojIfFKchE9Fv8Pty6ezyyeKNPo51djOCCPWLW+CiCmpN
S8QR15LE0ExeMV2m01ss78VYrMyB+jqq1qMEHL3pp+kiMAdALPsydeQQyWAm
IXLHn4QnqhoIs4Fynj7Pm3aXcNdQHe25OjWb8U/HICRDoSKOASJlnhr1KG6A
AqygDxFsNkBdr6NxjuITDP+aeFwa4iD40JMz6K+IncxglEfT9O+spMLO72VS
i7S8ijiQmBh3btJGbmDHia/eaP+3SFjnLupCqUKiIfZ2Vx2i6OT+mqFO4Hrr
hDFRXzkiyWQarLlqRx8PuDsMhu4Z1wlodpgUqVYQenxnjhLVdwMKpEh88pgB
n5OEc4yQqlLdhQ9e1nrbNwZOskxrro+u9FHJANT+HuEAJj47D1Gq1nnXO627
M5kn4+m8gYq4L1iCPuXKQACoq97Urcp1ZU785TZwJ5f/UJ0chR706tgxuviF
j9crR39441H22028FzCFEjarKlycDBo/GbDWH5XbUzBcItdZstavIoR0q7EU
dWJvf7eT1SGa8PXmm6fOlpfOCY4a5rb/wlPSInQovOSJsKagsdEpsivSrK2l
30lYaa7YdLvgFWTGdF17j2CjCbJ4egUSYE0lu+2EYBPD8k28Y3AJbpdrrtG3
O+TgyfGsV/qvLPyU0PnmgcwwTiuNWmvaeURFZG6EPOHdPQBqkQ7trLl5eMMB
bTjY/KCpEsQOlUMB0CZQ8iVuNV6P8DMi+abYNAerqvH3xdCPUsBxyBJlMMni
JYUkuikXRkS7EHgZ2kdfLNlTNyg/6vp/ppLu+AAVvuZm8bwLoWMGKP2bNGkI
NEfQ8cSbsnEA4TATObtZpeKSYmVdT/az6+nuR9IyFkBBtUvEMBZUUhE3mXws
lor+cVFVCj2loX65j5kAqSVoZgommSrGhe500NV26lX+UFRrYR8vbCCmaqBx
ZU7lryKUghUnkE4xDrEQjdwldJ8iK3M4QaflQQipustIt2Inio3W+DwMIlPR
W3Fg+twm4k11ahSabyNzgiAsDdeYrIyBznLzEfm8NhZ9+DhQe01cPmwvB7F7
COyAycQkgmalKavX30lsTHA4E5t4Wg4KfOIm0H4jqxd4gyTxbdp1+rY+98K8
efk1JTZtyzjISejp1mdfe7fFwmnEQbz2ivvmSB6KLxNjkam1WhGT45EevuJr
0euIuqxCVaSlEfUr90P6+HohOOCzaw/3xX1WrFthS9L+R62JnutRqC2zVPuf
oReyJZBO3iwbbxpMQiAMBa+TsCbjMPRlFFkoIb2/GPO9G9c0twCVi01wCuF1
8Utdot3V7X8r3R+rL1Zea1greM2rGTuB8sPv/BJUllnACWrciXmflsWSL1OL
imCG4A9yzQIpbCVg0ekScupcjAtwGntnMRiDHgwrF54ldrB5P2ayisYa0HNk
qb/Z1ii6tht2vvSjzqg9JHvKP8mTjVsSOjezDN41slVkKkkJW2fPCggQlSZG
ZJVKUOkoQ1L39qMJBvlq8vJRvZ3BqcmgUWmtAWM3mOUROgMsTy60Ta2ISCjR
tNw9E2LIoSAKTWUb34D1NbjG4uP31aCbeb7cxa6xkIZpVNmQy/67ma1HYHpJ
q+7fL4Hy15KDCSiyuMfwLT75T3p9oyyCPDJlNlF2W/cydMuPkGYYfWrtBn7s
0DPgVGfRBL/keQJ1bpN/yPOA5moDml2vgmZ+w3GdwJml7HW8ecOTRbk+gQDQ
gocqJDhA9Zfq6RSo22iYD7tyAjQ64Z05V5ffPgKC5whfH8ueimk+bDLU7lZY
kMIWphseKgHgiK6Wa1lmuSiVIxPpormwq6lpTeC+CmOIRThiL0eRLD42eULR
hL67VNeNuO0Wou9N50EghgnNkdVUDOOXaOxx4eAr4wItDTA3BxQWuSzg+2Oi
eJ95HRx23L6yF4Hn4B3HNHYoIPTQ951Wc6carK/UFWL911xJhtyT0CA+lEA5
fAxB7JPl3lEW/WCOBFCFkd9vosr16iTQxpRYZoJJ3BBt4tv2SmeExXNAYI+o
PKQucrJ7PzKAyLU1He4xbv4zzT45gFg3n2bSITTZ373DVnrKWUbDGtDkfHit
/D5ODb90Qdy0u8f1JQc6miGM9DW5UNYPCG1WK06ckqE9Qd47KhfKjh/rgoNL
J06kto9fixnBMkO60PH2jVzv/MQkWoi86h60j0iaiF8CjAnztmYZ8Yzv3j1c
GiCzSFWrN1esLHH4mgpsgt7hrrcD1vVjdyr5C5r+BFg2j4ufBMnehZxJvNSY
0r7idbnBxUpoRSGABasCGHvneWWoaN3uaMrj+SNtwVT0+q/Py13epE9K96YD
RhCxBCvlGKuFVfXZymlW2539J+LoN6493uP8PpVoJDP02DhVaABzCmA9oqZ5
jj7iG3R2YoUCDxtkV/twHObOQ7DVX/XAJxgcYuFtAE32I/6eeIi/a3DdsNaq
w6BuY1lG6JE2QknhioBuu3v8CwAQVQr03hMP5ZlJ7pKVD5qAwcaRYG1TNxyV
FxYDJCxXJzFkuB0GTk9LEa+xBMw0JWfglp7O3rGC6SykcOFHtXsawwMJ+N18
AJkyl2003wXpRG5CzZzIM3XomMsV/d/v+8flN6B2IcgNsznQ4hE2Bt8ycssk
KHdXQ0oiuuBOsl+nKbzFHkb9u7d/7PAktmoIfE/V+YqZM2jX6V6CNBxt4ZaL
3hmyHHwYRq1AP+1MSbjwksBAvqKBkba3bcGoywqduVgLcKpJ6DbIHoXVVTVy
+eIrL8K9FBNEcqVQduddWZy+53I9guJIUqlrGT8eP+B4elHQAc4trKKel5qF
E1jtMwLnDmc+4FFjSsxp+gu+J2dHys5k4wQxNzxlPtlZn2WCJwy/g8cmN3WU
xb3eL5OMdsQKGBQQ8KieF6HF2u+wuNPBwbWr1Dvmfa6zOGcwQyx0o1onhxqX
2btnvSAPwJWtOfUcwOOLFqoyMjJBSfxh5kWlAZCrhtLYGebi/MDKbzEbA42s
cSyEI347ocXngruQ1mnAiD3fVzGVEe4xq62Oocf56ZGH5Nk1lQkza6b4j8kk
NrghgROCbfmcd+a8PFtvURV10N9JoEUGEaaTWharotXdm8hN/nhG3JvxZ5h5
dxC3zqYtBIGMcBv4jRDq/4S/1g5jl77sTRkdzaDNvNypqX/QOR6KG8RmCGXH
RVAIFXKmHDiahp1xREyx53zR33lXO05bjP532j0xq9O60f+oeUsOKqmspxAz
M6G7Ct8veTjcvGc/pAtFHr8KuCcLeYD5M4WlUqiLbjDRYv7xfXbQIBBqq0zx
7AKBXzmOXTalN+Ckr4aBZ2/sDmNy2zBuK7ArwEbf6edXI1GnG/aBHGsVf3SJ
HdoistoOz9Jh4tBx0mBhSR5lrqnM3wtDtyW++3g2JfjhTlq6BC0opRZ8Ch4Y
VxkXnCmNmYry32hD13B8OffG5EhIIRmzRHF6YAF6IGAm5aJ8qosxt5iQ58mx
0+DUMf6yzVjBuvwgejpxQref0g+9c+sUjQ7tJi3++xxxj+f5TBsVRtmmgvgu
hPBIE9EIbnejG8kA6tOUGSnrLDVHG4DiPJqLVHw1igtiIN6BDqYsyLamIaol
uWyaP655pFNiSSNkkRKT1YA5q6l73pOFG8VCBzQoFm3Zg6MMP7fEPxzBEBxv
Hu7RlHpGre6y3WC0WCzIIZU4KpoWkIhK8mcjjTJwfxYq+PJfmaWhLjZB3WZh
blvnJZv2WOGKYcUSY1/6lgJEZwVeDET3eH6LbxXGXmPSIPi817Qq2eTfYVWD
J5Dyz+FqhRb6GtCJdn/D3+9nSb+RxX2EAe/ss8W1M/2gObjtPPl38lHxYTlo
tiRhXiaGkEDS4CzYW6LqKadiWZHs9mo6pXCFsjHNQK1rYEomzdZEfu63pqYq
GREMe/UdV5lCS7aIyqPkyXHQjbukrQrkhJYEc4yxI7pW8ah1scK/kaJBt5k2
jKWYtjdokL1pyYd8TKAcYsWY9FglJNgEcbaPxtnUFVmxwQi9PK9Bu7bdSU3w
RUe/23s0PNdkPBa7evRiKpSztfudIupXGhLpzL4zRKox6tfn3KR1WqEaYlTE
jRt6w1qF7tceeyjLUlBYYGOVwv/NAuPkxwfP0uCgKM1jV0OIOgsNxHUWEDWa
3wr5K1RNUg537AKBEXTVFkhDRjUgJ9j81rHkM9BMP7ZxbLD2Ox4jrysPsnzO
R1VbW7ZrHRlVqTNcSa4H/2J92TmscmSLCbXjGfJnYvEYg5E0EEMlZfdB7Ilv
2w6sHVAiml8FJeeaAPBQs3oE8vQcBufaBBuu8aK0/LRN4NTC7vi6+CzRmTcH
IwneEU2k7rtdOoxNza2qRXDQstBoqHX8Ze2lSXuge4i1/YwOH1mYjhGGIefl
1G+IeUFvSTTxPDURDk3TNJxtX5wwHKdpecA8oSfIxkrv8kbQrveC5R7E/Qnc
ZXCAe2gAplrJHcKs5m+guSKplPuH7yZTRjsGcNDHN3SV/jEK+U8quwWMBbhp
8TQseMH43YLWx7hCZgCoOHKxKmQhqChETLO3BJbX/ETd3IeMF/adTHjShNf/
Qs2Fwwupv7y9J+TqSGP7TA8br/PIZOlNV0SS83K+hu2mdefslaj5oCZkTZ1B
RJtAkaU09aiTTpMmVthd6p9J+YgPP2YdaPGpdGaTHkMupeE63+XvJVkjB+Et
kYQOKtvXRmXXXiLBAvq7kQgILqslwBeh0ism53m+xTO3IMgVv+06l/8EQ2vd
c3kYY4perXsMEZBVj4hi9A1awq+RXWWHp8FDWK/c5GElIkT7xYUoU9D5U9H+
u3qfrL+nmsAtmNX2iyDmSYm5yGwBIsDAN2pEC5gr7YpbWBNFY8KmeedVCNoR
6n4Be/i7uYKwBTGCmCtERimZ9bwC12SdIZ+SipQQNvUf0hy5kKeosFJGfegr
YzvFxYZ71iugGyl+9FJ5s656fn7y2hvqiLYxhwBRpyJKKQm0Sdbk4lBXO6zQ
/57ZvnjAubfSLc2jINtQZwQiFLQOKC1X55k8stgbnQtjPTc5GsiE5hqkYOlR
qj5L2bAurY4zdUnjF+wde9810ZN3qwiUaaUKqB8UMj0Hi8bwponFQz1aiQ+6
WpwKB/YjvMVj+NSLAGJ88od/Sk+SJiZZ6h9MW4kOp57MjwPtXaKR5LkNvf4n
1fkzxbvDMNUlGD74DpnBd5Ti00R23Z514nvjycBeobKG53aEP5BkPb6NWq5Z
UaWmNzTB9ZtDrlYsKIa9PcYowu7zd0ziggn3FOeCej2WDITrY5JgZx1+yDxj
Xy0ulstrtVlq11ucu5byMcsoeX71dC0QpPc0873LIeGdtW/dypOsw1A0kc6P
tSjB24Wsa4fgPhe7zLICIYKlKTsGDT+GWLW26FUAIZZotfQJL/p7ta8VrtKW
jYbgxmadiZYI24enQ/JB1b5yyZqla3XnZAdk/7jhSBBxRh/IKW57jVW4gKdb
i38PNpwsb0joOETgqMFptdpHPeyUP/8sFGydAE5033pZXyNtdx4l+TBIHqGd
VAQFqLXtFOUc+VybIGuavE8bzbH1PE37C4R9AVLCRExhB+r+KKx6HTiQpF2x
JJqa7Fx9/KD+VFRrUMZ+zcFveIJgtJ1Ry6amy0Ku0CclJ+rTeUOSrimW5Mch
59GgjCk/6/EqVeHAltDSVq9jUgS1vGsyLu0zJdKvNJP1/zQ644F391bdShvd
3XTCYGzbLsU0gDKePd3Sl5Q6+pswkyfWbJWngGDQ1WFUDhgZDrS1hMgzN+2K
+I2GtARFYqeZuFlVZTXbKjixPZi5Kklt2PnkkJ9tdJuisR5HY1MchU+4dRHa
BRHozVlsyQ+08/hFpFaVhBTlGTFuWPGERNq8ge9UGiRF67aowvaZR8KvDHRY
93FsBWR9fAt178VoBCSPcz8GzlxnlCPwg6UpK4kXPdtRjsJuVb6iaybO5/dp
1FJzeIuDJgJ4XW47pc4ovh64dt0wyYB7yUPKElkSbHtcTRTwcQE75Ve9LVpW
bjyUSNMNPwZ6xyZKVqxmfJyhNo9XrjfMCpavtMRn7lS4/1gQnwvgmSogzQGv
RzftGoGpB3LU7GAiJUWLPybiuBS2dvRmyUghsUGQ880ErYdQho5UjQrBgl4f
/ep729bUiNNS3zWXH96prdYdfpLf2j64EQrjw1lg2RBufoXRHHPWP9r1GnI7
NK8Oo/PKhHztuPNF/GykLfJuIHCW78J6XLQnZhMSzSgPL82bN8Elvz7rByAd
DEvwkBaTsfnkv0NAVYVEXY5WPfuu8mLw0nGuDJxHPuxQbJBtmkalGnQxdiuW
QLTL78XG60gnPDWzWv2uQbCYuvf417ZymGsQOTt40icTsIaCC4F0QNOU2AXc
Dpyl/EavTBfHU1u5G+RTGDqjePsDvj1w0AATSN1p3uMzmTQGHDgSekL5l+hT
aniejZFqz4TU82xJ1jtKBcyyZFctf5QV4ErJyx4hmDZ7RCjlBCWNaJCe9IdG
g6K9rxWIi+nyzpRp+3w47q1OL+OSQWSfCY5k7+sxc8E5nCDJukVWpCd8ouEq
9iiniAxoWDwncVnj2KpRslB3Rt9JLEFNq3x7V0C5+hyHD5qhiGD6SitSszbe
j4X4VbovB+b0OKk9fzRJS0r2uG17pZQoYgd2+HJgqLerW3xA54smr0SJxyoM
aXHR1xoEtHd735UZtiSacWlyIDTdAMB4Ni1+DpcGcYLkYOEk0EDhTQaRA2r7
tekJki9bwa8iMGZtvjg5usTP432txkaQ/ExcxVM/6wFma6GxLJUiDtNf4ekS
hAH1tZxDqvOe3kWh6wvkRSanGJh5NkTABOk7E9b9Rz/LF5wiDCsFd3q1DwJV
ma15+ueDN+Svn+eYkWvDn2fxhRkei6q+fw6y4wJgS4KkMxBg1I+OrIdijEQH
BA1IXv998cDy2uMSDL1xBSnyyohG+fKDHEf+oVooqSEeD51r46y1CA3572XN
1gnWOVlzKfIMwwjxtcyyHxuWPX1og6tTaaS1amDzC38hK4SUZMTPcGlCwC3O
fhr6l1qldyg+nK2V3l4vxZ6SqpwaN36US0Go2z+CdONWEkZ1CydWTcJi6C/e
9adqosWbnsTkwpvtu6FSbFkKR6V9Js+3d+SvdC+O/xB8E4/gtQsh/etmaxag
kL1umEOFcvNxJic10qx+SCfFJ9rEhZ6mzTDHH8IsxUFApE8BVuSRQ86XoMQ9
0LY4HEHzfIm0dQ+L6srx0GjwaB29nuV8mmBTgFhQ6tijbZZqcHmPwPETUt0X
pRNVGSOJzHFlYq6s/k0GcvrOHGpPWM+8vf+c9u+mjOm2oxtQEVKKSgGxHacE
yCcOsCwPQr5p2ZG13l0infzZPE2YNNj9o7GTdTgFfKgK4s2cGQ5NqIK5AdsY
y+f81wbtUs4ewrCThqkbVksmaMwJZMuhryOiRF0G4N1htoA8ZBJeEKuBId+X
Y2k7kdQDQ/yGuMFeJ28OP70OtWUJSdtsWVVie3JHL7nnyBvHq4XF3OKM7xfu
Sconv2n7oRJlE+MIHsJuFuM9A523SvXcDo+CobvyqdEhac8DoV9xMN8v9OzX
eTwAugwVSSp/RYaUVftWpLrgQCgfRZsb/4rgxe8gOaUtTaxizWWjI5beHtt0
pVg3Q1hju2ZMjJvAGeBKo5zAAVK5nUC+qxb3yhrDsUertpaCSDS7RdnIi0JU
B28meLcHlYzJ9yvcxKz8nNYLzBKqlgFbpo2Rj2m0tLJzJWdAoHulvQTIdv3x
JO3/B9UJzFsTa76Xy26vax9gTo+qouYDKu5Z6RCMBEnyAqsTcsoSarNiV7Mj
JhgiBl8M6Va2fHPhjnIYXQYw1uZhXEX2GQJvGurvlLYj00uWRnxbuN9WRTy6
TPa/spn798It4qQZNMSqV+pKzX0MNimv9fVqEzH9fzvdIWHfSHsHKma2wAEX
9yqE1upxGHmLpfy1k+4VZyPhePQ2FRIb5q9KmBkrgUrmQeQ+CIQrKA7Vl4n/
ff7XTmTEbTShV2LLbMbes0t3XG91amJt8Ty+VG/B1L3jadNNn5s6gypxRXbS
onuL3uNy9SyIJWDX5/LULFhHInj1AdJpes2Ctas7Pr+IsDD74dZ7KiwFlZtk
KLtiNNWsvpqkiXxhiuo6Ef8qBtDkuubO4r0qXk5Y5sDtcLavyEBAZA0t2MT3
WrXjRYsg3yMEwB0aEWY1l10qaJXE3ladGuchRYPgOBScrIm/zx83TFbdcWoc
MjoYuJKPonsLEa7tD4Frplhf7Dmvmx+mOA86D9ZYA4X2jhHVT4q/zao1CBPv
9biQF8FPSky+cI6KUGeYlXJcygz+mlCShq0xu0Rrd3q5XZOwzkv17GHGQwjO
0v5P/0GGVkArrA3pz/TcwTpldY993jFLrAziEgf4569ecihUm6KfXrT4wX/Q
D+Lp+bHNlwnQ4v3+On5chRQUVrCXuyqtebp9N9hJdLxr65+nNWcKR+r3C7Sk
yyRPx4uTlv88p266UuRAqwpoy41tCMV1Q7mWChg3sRvdQMgvBKtgqxoloMby
LrxWP5cH1xJDmIM5mlwDAinqR/EYpEjCd186C4K91mFDVy9f1tZ2f30ODr8t
jxTkh0vQkTn7hwKpnwXEmOO6Y9fUKo0CdL9ZCY2Mt0gKkVPDqL9/xt4Ue4ji
rZcfadvTiQrNG+XVk4UP90R+YoyjFANaRQ5v88S3+Z857/ZozjD3mLhPFYu6
MrTeutJnW5DGYo1UF2uiDMH+k4SO+zLKEhb/xYXsffLpRsQux6SH6YyeLDCH
FrpSzJnz/NT2J/hBjeXTfB1yFYzc80KaFvmcCmUT2VpsoVV8exTssZlMzpNH
wSbmN7aN/U9YCGFPLIIZLYED4JokCeF3ZeMkC7eVeDV/TzlldzQQGilc2EG2
/JNtCs4AI39Yd3SSsxrNwQIaCNPnagbr8jWjcMZgCb5D63BbpS48RU8pKCzq
72bd9eryQQhBis98aDXJEIiLEROcNQo7Nl4x28MwyHfa9MZ1eGcCJCF1/Cae
pROjjPeWmj/+ycaaJWk6VAu23GHbU56z2U0gZhkLwZ6rHk0vVLCG11xK8ZDg
Q7d1CtCH8eC0grCHn41Tw8LKxvRTc4rngMDGEjAEb0ytI7oXmygUkUyRkHXw
J9H41s+4QGyFxiVb3lUejXVp1Rf0iLqGwYFIxDmDSMWRHX2saw1TpKhPeQSl
f75FHKDwXvboYZmqBGpviJM7o3bu+GXRZXCS2C6k5P6KKARLNyvDaBoL5T6V
rG8lv3oAOck65dwY2qGIRfLvTztxhFRPLHWkeLyKz3M8gyJzIqFFOMj3ch+Y
H3LsJpP9/fHHuHZ77dYxRbKSChW7VymvU1h0MbByhQ2HWQU7nnzFWhU3Wfrn
IajmTW3TOhRB7aZlH5MAhg1n3rjFxIVqWRasx2kwdp4UXaW95Nsc6smjzFaz
4T/dwI63b9BZuH6alsPhm5uk+suLqrcn9lpdvQQdxn19NcDbqhqH3Z0IRuro
aRbD6rI22HQfJhdeQAhmmHr5eS84pgYlG0mKKJrpZJKjLSlh7KCDYYVc2UEn
ZOuXWSW93F+vqzT2WFVaYLY9i3OOzUuTP3B4pa3syOx6kh0xImfMSwdQ1fAK
zL2Kjw/M9oKRT1M26yxlVVEhWPI2jDxOapTTYkpcSYk1Wc+TFZd955isp5U+
cN0n1OL6nURPK/voQnXCDzeEM9/INJ4QUsY+99jxLR02QSnoN8+iA167ZmhR
C7A7vGeDawAm9nNg5yM9NrTfOtpMYKLdSzAV4k7W0i80MHtGSnVJiJwdVZQ/
Zf1pJMANDywUj4sIYDX4XJDjmBHU/JHLek+mWKzvImHbsSo7jNofqW5FBrbj
El7AgvBJ9uxTXUnalHh5EAqc23TxxkG/beODHwi2kzlY++1HKnW2B9Vn1aqa
xdBzHoDQC2SmSS3rneSbOnLeKics/odncuT31W76pWWLf5HBtPA3w6oZaOx0
3IM3+Umop7NXNwysIE3Uo0vW6KeSRy+B5Hlsc5a/gfAk8E9OcYHEh4ruTm3A
DDRpBJUN10qeogWzYEk29fBmBwRW99BeLpYO5SAISKoZwgWcyaMTifELdikX
tYaHRFB01NzU2sXs58K59eqZyfoPWvG4TvcAlhzf84OtnxozJUWQ3tmPonu2
RW26Msk+yOfBuTbH70PCo48I/xb4EKfTXV9nEZOFb2JRQFNOx7llH2OLyRLP
ON+UvuW7mOBxsSqfZdJcuDRcwRdAYpfAXWs/6gVfTmM/2RAmkS5orgUq4Hby
OoIBmZTFGn5mKDpMJJcyXsol8ul8HV5IYUVsNQDUtYYPrDAR5mnU/wZLKEjj
vtPb33e4gTxaH+ywiB/uUH7xZtCv2pZk/WUHu8KcHO12+SqAzhRa9wtcRLWy
7ZdjOuUshPv6xEuIeCaG4FdbwrNwdOsTkNfYBwp5hsLCvjUqovpM8ywjdfO0
KFitv5PPtYnz7eOvFh5rFNdhu56YOVGh8BOq5izZNk/hvPEWWQ2RZSDsk/b2
OLgTT9Wh2h8SPNvH6xYCgIESFFwXjXnpkCJS99+yNSzOzethhF5W09FGsYU5
T7MwYjNJUa5N588zfvWFSZhEtAPl0Y9UIzLjiET5P5zojOA/V8i8IpHswzbR
lijZVOoZeRRuJKef47B+LKbHi/+QkK8ei896TwASGCnkh+mc+bcBWiaqqEqW
Jk4xJsUjVURDWF+YhjTO4nhK6Y0PHONCHt7n6g0VzP99shDVLr7kZA79HOgA
vup5HzOIaPzQAVze9eVBuJ6hHZpGlwnRB9eF6dFz/GIoKgWEbev8Rr49/S+7
cGLgpveqNkrlBnUMBvkgMdoHQq9wn4mIlGjsM7jT3TxoqX9rsgCUnLJNgI67
r1sqQnl9sFvHRgDipghJQ8DgNHS1uZnlPwUD3kCrmwF5akXY/AN0hUDwylDW
cG3YFaw+hutKDd5YqQci8bjdjBO9xRHPdGPN3X4YtYX/R305Ffyo0kPCE8Jw
s32JF78Bz2Db145u4IBp01F2mOOSD/MZBXoOFmYZnro0MUKqE0FfIMkuHbsD
3Ytb09YpbSMw3p4G/MR74oj0iEMUokCHIyYRuVDqqwhrzmc9XkyvUtoS/ehq
qKuK47DpvWsw08GGRj7B3E/b4rCwlwL5xIx/1bJUUF6tV50a4w59fb1B3LSS
S4JSomOcbgzfSHHq3VOEKQ4ZCOSpYto5S6f9bHJxLZvIm3crgluLWoWTS6gm
v46fvuaTWz8Fv406/f10eMy5XZMO2FmVacU3CFXdvkatcCJFJ0/VKsUbrk7R
K2Y5iDute5aI29FLlSyr+t207FGQscwS4juGlFojl1TIsx/6akcM9zKQ1F4R
0f46R9laMOX5mTZaMCQwkmqfRDQ0c3mRvXLew7ZIkWcl75xMCnijOYrmASN/
jRayfUBNrknoa3rnVC6p7pfGPSXQ0nJBI9u/XJrMadufjOGGuVZKFIRbouLp
oMQqS/UIViA11ixKR2SKzY++TJ4qzl3MLfedSDSkeyUUlH8f9atbqLPKaJ02
ALh2H5teFj0Cw6PfZpyFxscBfOus0znBHugO1tF53NjSaZS/UQMHCFM/Ag0D
QwauTXg8VPRc7z7Hz1PXPlk87zP5B7Yj1DophnwvA8/RtxDLalA/QbOrVqyT
ULqwtZ6B87xNrdxkeApetFtbITM8KrPxbmhRf3jzqJac6tBgE5BYq9eb1+Xn
bCync5neq8aZR+AbapRkBFNUVToV6FL4m2MT17N3vyZH4kBAKW567tBV9BNW
H+eTsLcBHCHwDK6dqQ8vTwwwVkwkxoEsd63ByA71jcLi53kxXHTcp8JZceHp
H2KQODzdZCgwHcWY/fnFRlPlVrPeJ2vJPXBU2bx8m66tmgWYTEDaHU1w2JMo
EG8Tq7EyRKm986f791asSOgN2Eo6ZPBS9VC6/seVyTLPdCxwR2jOej7bBPJB
ZOsVScmT9Hoojv2Qxxx0N8dM4Z50WWgPxZaWSkb39AIduTznKu3OENZizBtP
nI4KP4v0ZeqYmRJScea9FGH4dhjMtKgLFRIoObHtAYWf65nPBxxnrBVmiRyY
Z4Qg1yEV/57DtzGixPaYqYnVXL3xJDkHFAzMvohtIfkOkSgYEVgbF+geyoBF
+s93O3r0qPVRXqwQm2paloL1mTKpI6f7UCDkiEGlOT47G/a1pE/9QSbXNO6H
V0bCkmmhaCLdxpTHzGry/W6Ui2LnQ2EvFGReddzsq25Np+XS7vUNsfSXFa3L
ZvXOxzKI1sc5QsjqUWY4lbz6AXhA2RQ7nLCppqR0aN0LgKFulzwhAqwa2PFx
gncaaFaAvBOIIvNjseq8PMM4i44Nqp2ocLQHpgphW5FeRlKZ8dRl5ciATQJi
NImJCi2Wgx7iXLn2mtw/X3D39hAkclFg2EgkiVbKNA8H1yk6oy3pdBK6wF4p
NExdufUE0lkeODBbtZ/fXPeNY/5F4eA3LjJXRQQdacYa108vm4J2cEwHo7zO
0WAaklVSIkcAZoGdcYdiW1YT/+a2qFaoJ/yrEvU1eZ1DAD6q1sJvKNc+059+
+De2bNiGPMsxqtePfqZv+Q5FvAAkhZu4QzuB7/sy9HYgD2NVICWU8lD8nc1f
Al4dRNpegqI0TlNnARKp/CSJ3J5joT7UoB9r5WPf3E4i1D0/GWK4w6ycjuAK
NM3sTW0Qa++bCyaxUEMF7e8bMh70WLNTfj+AnviaKvLnlwJph1gxy50f7diP
JKlTqy9cEgSRkZuIAro0ccHS1FRpm49ID0RG04rzjSg9HDDpnDY2KeT/bPBG
auFn9NEctgrNs3lm8PndNl/WMFs9tHu0X+DGEBI4l1sYXCH33YAgAUaTljAL
VtOqtMS2IZ4ItyPZcVJOAlQvBBuCJMphwj5J6Cp8+jVFzvUqJVyGwMlYzCet
BYRevaEf3KlzesnkuVYeJZ7kMoncurVYDjLvJUb7fa3/fGngYCPLLIOao053
Mh/rdBx70J27H9skOX3lwkcOVBANZgSQr21/P32jgEDkC3VD4v8wo4Hv5020
SVdA4h+rY3kwfCydUovPvzDNoWytwgjdF1KGBKVfObCUIJe7B8WBFcFHaqJz
LYr9JpJn9i0qBtilwoW1bOcRRBNfrVS3sZ4bMRNx3HC9xLLLp/oUsw8QHmG4
w49WkEEKFbxJuu3KEp1zawsNlg+y+NXtGemM6o8a16/4radp3EUlEk8gpj34
NfY5BfoYRLdgm92KMfZUZQ78mFtyjtbLVQY3I8WkfJMJjRx1k0vxmyBYBqJn
8dT4hG3kVtJcGhcP5geGgli0cR6+tp8XBFUDi3rCAS0efLBwJ5HAFmwDka/m
MdEN4QJVC7q4JB/dOc1el0P1cMJkYJOUmcbfFUI3C8Eakisd5+0pBsLFLqyy
THRnTNgVgmWW3zG3S9p7bCnMuvAqFOpe7D6pSZlCninErACGMzE7hx32CLH7
b8ZjHI+GE2mQEcRzkar5OQQmQvvIc2eL1fJSvaKGE5bigkk0Kn2HcAit6Kml
KFoZ2IdTh6Y+2+7OzlwtDE/RNjRV9HX3jACv9ZqMLqzcTKXRS4LyUvpJATBX
8C+v9TGzE9xtmSLW5JAmiOKnKvJ2aTtfKThtn1lvc5XojHbIfti6W+gAtrId
QiDfG4TFY06/BHpkroAFd1MPgDMncHaZ9YfxktBk8L5WPxjk5eIzdR2AG4E/
vHHP50PAW9TVxx6bnkniL/h5PS+2EntlcSGjalzfBYDxLJH6VsfZoQU1VBO9
RXaGx7JqZOQXcqRl+tZb2Mmr6ApRabGtMug6l8a921kknE9n4oBRzwGuH88T
Xr3lb4gUmAc1IwryGE69zihWAjfCksBaz+n39QL6CxcloUVFNwL2fstPXTYC
yEKtn4asfS5Irj30ZzT/sNOpkCf+GtCyizO5KJ3AP8m5Y9gkUs+QX7Wf/2lI
kt/PCJOw4C5f0OqFJQiWSbMXcjGf5bjrijY6b26mVRI3yWU5NKmdO+9onOBv
/h5qa7ngiBRcAMY2N3uR4eroEdfTY+UguizCTkR3uvMoF4cM7Y0vvVdLEdzD
7OGkOcheaZA+WLR8otz4syzHYmSpyU8YH/Moumpwp50dj6iFCj3sHC/2mBL9
m9b/IohFInJ2f9YOH6tnMWoHdXOzoCVtNyPTqztPDrpspbH84Wf3PkfNXlJn
inIz+428nky9UP6g77qNbmId6nzbzIiLb0Op5L3jKrWwoEMpw0LsVlZoFV3A
gijk08PS4JGsiLS0SoKReKKDTm5kZxsUP9Yhn843/R0wCTVLzyCnI+ERLyjO
cLok/akC9ruQxIpfWzuI8rh0L+gx/1inGBWAtO6NveBmXixkms6eoxe/JBVv
fnHVtuh9wEa56I1whFjdkUyguY/sQQSrGth95l0EzX5WyJ7y0imWNP3qZhhr
LTSRpbwCVslyDAe9KODhQPSEf0JgtGNibhvhb9TxKAp0MoItVYBE94LJzKX1
Vfc2rSrQJdFNo07SpHjBYBqDf+QAzsZWSgtx3PkdffjczfQSm01nJwc6HHyb
8tBQnaYwDAE5+L3PbvP4NAC3XEPszxpLMvjo4tpNPluwcnA3DiPQt26mDekC
os8qTklPLlAFSzcqb5WX2oN0UCYpbf5xrD1tLLC2K11HLDvrpSES4KrCbeqz
peyhJOZf+UUWW2FqhIgCLCYPdn47qKpDMXNEIQjyR87jNKbzFpkYmduMLspP
n5U/6oGsu8ht8ZM9659knyiLXYRp0q20G7VOnkQxf6BbXBqfws8pw2dwi9wK
PZZI8eXcghgfVX2WayYSx5M30/ByEMrR7BfIYwN7VlqE+OZrsopBpifWWOaB
6nlN/2JBYOUAUWIDQWYMasZ4Y9xF12PDX5sCsMDASUxKNtpTD2icjAUrjgGC
5nYcmD3PjS7KY9EKtQEYsGK0O6CCC/KkXgTT+hLT8q15nUdbLiwcY/EVGxMY
OT/T2sPIGmfTLev3Q0GHf1t2uYppwy1tXkUav0EJCdjgjtp3SCSlkkR9e8mc
+zcMRQIL21z9jpNasiqmFBk2qbexfr9nSNLN2NNQLiquctq1TTS7pKnmHG5P
4aUBJEHN7UuOQ5SrsAfpvB/rhtj4ipzuhBMfA9QAbmcauKdornj3B4m1ZLGz
TlXawIoft7ksMuZzI9rTs+3enPSkI4Hyo295YuD4Yl+7bziHns0cShekWRJ9
xzS/fNbzvIjN7MhfPe1FNpOxhC2JzTw+JgItPi08d2FgH/M7z0epgeq/FTKW
oztP47SGH+2Z1qXes8y1k2wXTBTgcgaHk85L+3iNLz1Qf/x6qPcNZwroLgs4
dPHwTIFDxp5D/FyOlldrG4ogmOvPFDT5Ptf62znU2G0ssr/cytnkBFkDHfpv
SWdGdulujwLC1c9cLDK2jaw5uO1TepAiXFZwpy1duSyBpx5Uu5r+Nh4K3lNL
iq5HiMnJz8146r32QA0a8K+nheBHg5b370QJSFjciYOb4qF+3pQZy8o0KsUK
E02OlQelxsQONIpMgZn27sXwr3TAyuDGJGQr4/R87eEw+4bePqcm7fP1qN9i
ByV9AXNudf67E9BtJGV8cfOfNjNVjAn/FQJVnyTdyNLZtpERtSMrYesLRh6N
Mjdah+gk9WZUkM4dWMh+6/O3nnAY6Tgiq3L7TmR50LnqrNAUPmwg4ce3KANA
2D7+sOtUG2OaoOoDmxzCyz9HF8xLappKw4+cv3tafwWdsXliH4PJxGLzgkmV
x23oz5kJ5TPlWc4Tk/g1DayOxXs/6e7MnsvH8quoYqwXdyr052Ak8FXajzDg
JgXZHIs12OKl/o+UzZc379i3ywxAurlewCbb2gtUDpmC5q8Qat56d7+jQ4KT
sNqSq0HFUZaHFU/CZUq6MnTs3uQW45aNkc+sPxfEh/jqFYqVXZVSIloga+cs
hIa0UWjqqZ6stPxscl9nQfc/+I3NEd6bxAs+zxTYE+Y5lvmN5QMVudzRsxR5
6ma5PfPEB1jt4ZE2cZdwcCivTLKB4CHEEgQp0tOW5snJyJ5GAbSyPGA3wESF
PRK8ZGJZNMNp0QWWyQ/gFnWC+EJqAydUOUSTM4d2wPosrVJ5ef66irx4GjDH
ToTnJ+1a0zP3k3AMwALCRUmiRqw4vRNx09QSVBlrY60eFEihH+sntqYmGM2s
kdFM5E6l5PMSvCmSHmg2kGRcl58AQl+kMu691yVsh2qdpl0ziKXuzUrtRz7T
d73ToVBIp1hmRx6dkRvdkvovHQiGunMXDiG6B11YdOXFde5PpOb5S2fEtQsS
H9MkiR+NxHZ8H6nV24uX/xUelsbRCbZAWV4iy+PnhBIduq8WsAZWP6c/3M08
qBu6/OBQe9zzmy2Jek+ttPjvUY17jmrlnLM2aqUaetEItxXKaHM1mg7ZmwQd
lhPymQd559olBxx75IeUikORjWrCr3ecBBt2FkIghmsrAS+qe09Ohd+xsdqY
hk+kZtomY2tXVl3JNkeVG5dOJIHwcbXKZTnVBPPiIDXYK1tQSdtlF2WZNkU/
8ec0I/QIkc5NoGiaepdvfLSObIzD/UpMZvTO7nSYa7aSIjyjjobLFq9DoG4M
uvo39wvofuGnK+aKQ9xfEKH8XISWRoMNxht0k8iLF/Q5ZZIAbtXxvsnhqpfi
lxzczTabvTwOk9qYjbhXWDO+fGNSQnGqdz43jx0aM24e25/GWWHayJTHRQqA
pG5Gf8LQfENZqy7EHME4iL/espBjk3qskSSvtwga9b8f9zBvkTjqbOLTsUJ7
FJwW0T6aiE7wEun8jJN0WhgNSCXYDuBWnNX8+oNVK04DTDGo9GEltIEhRua0
Uyj0s2jpYknaxB1lRqtHIC8oOFWPSDwPOFharCSpBSO1XtcUwThV5cZAJb7T
AqUY8D+e76/BjSrEg3uGOecoFQzE7LhYzoLURmybwvktVYmFrntK4Bg0xw5Q
hU/evXr5msLsFcsBMYydcQpA31PM7IpSVoM9jnZsh+YEazzjOarceNui6B+u
IQyEAY73Z0/ekWsOi/RjxN58W2M63sUU/TY+CpneMFmnf2Dg84wYfzcCV+Co
HC9QUw/qztcYXUQK7ibCZRL3taLidZri2TeAIrGB3doAkDBP7MWUd75N+Hnm
o68HPLZJE3hHQR4471kdcWZoi/cJmqgJwMquu7a7dDyxbm3hbOUcKngfN0q1
lYpkc+2GVhQJ1lXdm3Mu7bFMBc+3w111shO7K4McTI5+yvAcjoUAV8iThJmp
eq7Wxrla1UmwEcc5+ZYkcwgp3qwFT9BImwIdG9MhIfMNfo0eIgZ//6xVTKsW
0wy4szvVrBHvicI/J6aFco7CBD98yiWxnd+2SJ0w5eyHBN5Vvwqr65drFe3M
0e61aBChlphyGk6s+e6cMwJmcwhe7NKeS0katHt3CgL4PiFOevbHj7vpuN+l
hD7gYmjqpUhLt2S1tnfsBxBuWSBxyxEIRsAVCr802p6xbQc2Ci94iBqyAb1N
Q/8fpJBOqFug34s7CRheuN6+mCabDhhieSCFzRX9QyfGLj3eCqRtlFxg0nG9
nU8NrMG6s8IXpr48Ayl8KlZWSFwHJxDKr1L7Q0SOVRAUNmQ2fX856O0/x5GM
35PUPh9dHJGPeDvdYW+zOdzMvra6qzQ0cY8jLTgUJFcsTuZF8KGzQcA/9AqM
ZM8Lv7ECfnIZPQr4dYvEbfxqetDhC9b/i1luIY9CHpcLodu4NyZVUMKWTSBi
1Qc+1ToI8BGxS3bHRIOVT+kS6kpfjmN1XAIBx3IgSK3vBtb6XuvrQcr3CoSE
Mb8LY+w0bTfeJZ4QgLze1GelzeWSId75ovlW34peOFyIze8pu4PYjYgq/z7A
NYUgtAhuCXZnKTcw2DcV5m9BXreWY0N3dD1nBBZJkzIq5LKg71ggnumYDviF
PXnURyKMxcJXBpHwDDSBFqOp2vGLDvaq4FsA5UPcZNSiHK2I1zDhcdLfKaEf
Az4cMnPPQshjN3U9yODiNt/pcV9Vzmv/mqCyh4EKsAIgcVg8t+M4P0D+z7AM
rLnaKo5npVbo1v/l8GV747DI2mWJ4DdhA7mOuGMNc3iOdFkJBD9Sti4aTYDV
KedYPjh5cqWHRQ0Os9lacW0RBv5tVcfgGhhaRQVKxf5bJYcI5evPgRfnzRtF
E6crx17kXhTDEVUDrY2eaDGaNE9+2oNqIrcE2DBWO/T/PCBRG8jCEnRttB7C
SsqK4NQpCM5Auz2K9j7MrF6A2AFTYeR/YC5dy8TW4ebD5XbwXSdo8DUatFYU
RdW3QuvpDqW2djjwdbb59YP6e2m/RAhsHylDaBLSWXCiFtTj+akHjxKYekll
xjz+IIVlwzLmcyUwNjq76bjqJunUjMmg1Yk9W/aQdXRMhiz132+sNGDsqB9j
e6BDC1qRTRqNBoN5s53sJX9Lc/QPzTBC2YRvxu7HaHbfNL7R58O3Zd69Fx2m
vUXV7faqRsX1hun/Jwvv7JS5mJUqygNh80lNMBE+9HP8XHJ00/sgmM13gQb6
F98QBNSzGiuE1LUTFQgELViqsj7gprYelIQgx4RAeN9WQF6DyhrpdJxe0Whs
yPz3AB0+SiWAJK7x34X4bIpNv+ZQM7PKnIQD93XOo8+qAMsKHipjMeAowxyc
HISdE0VhGWZL3zQkCCtUcn9bPwC+CPt8DvqbH/QRLRjWnWoaYGDG363iNQa7
t5nyylGzE35LOJf2RbRMYBnrcrzeY/nTplD81qtV2ktgcAwFY8g5yTG5zjwF
k/ybpcpMG1VfZsDpn1Uh4+1h61N9A4O1bBiT7/dqd/M06d6Y16XtPThNrGA+
hLydu28Rv0mxR1DNCvyTHg/198+vJwdrNVSCwH5J8/ziOkQEGqdNY7j/asGX
lr9QhTdBD6L+LLojBpklNWQDJTt89B78IoF5iYufxQ8jz1yu4JfUsd4cMzWO
ZAgsaFB+xlT93l8mwqr0wTA++qaQ3sOPr9HVu+doZiUxLDDHxDM6KcJain+B
GHMNFhlUdOSuR06zXKNU5VgUohJ5FFM7fquyxJaiewZ8Dut1zb+U9BOhPrlL
baTJzSRgYjRvvOPSPN/7Kp08vbI9ZPBAXY98Is2HYHn36QA/owSuhYaFd5Kr
v4HS4od+BWRbM03oCsBBHZ7dqMkaaJvWAgzOKB7jOwptaLlfvZ08Ikj3m23e
7iJX2b0SW6Uv0Tse4Sh7za2egXkT8VwqhqEG04tMbOXlSjfdZIy8KOjeOtb6
wK6+8wE8EUmxK0dMfoNa7MqkyuNeH3m8E0RkA85dtgo+amXyk8KXz4KpoDAa
DI+Fajoihau2zDDhiyj0GuXSjn/lWxye/7MK8XH7TqbiVO4zYYzrIYywAx6f
Ji4RYX9tBCxTWGXoQQKVn1qcg5gKWpUnTAzv/scii9yk93uw4dxKkwRFLDBe
OykMAjORijvE2fX/cgQj5LyidWu/6i4H34GabKz64CWN8Xm418q5Q2wv7I8I
RUnXLv8GAj1gQ3vaZU1KOHxKnMNvznlWXZAHYyseKlTdJ9VFpw+pRmmo4mSt
lW9XCYR8d+VLb9XeFZo8AmuMhxv1gYZyFfDyBCxBOYMaZLMtPhQ/jIT5WFV8
gzRQoswo+poBRtfqplJBF/DbdcH4dXFRlcrMumBAg4/P89ChcJpkmkogDQnJ
VyXYitTreeWAewsnVXLL5hKOT12hEqTCENfX9nQkiTTqxEXyiwkfvjDxkHDY
uC/sRM3vAbx7vdADy5hIkHM5NWrmhzztMF3eNPRxAQNEKEs6e6bQvgLncDur
TjNiz6etEyYkZWECIRJi8Marf7jBmgFIrWFLWqMrni1uJBvWLcdur/mEiXuL
3o0zNz5uC7aPT20ZPjYVenXoej14zyt4/NpXz6cWY+6WFD11xY/wBiPsqTDw
eZGDD9zowMr3rsXDRxN5BwPdBG5NSM/BozJwSJellfx9lBgazwhcHXykmGgC
XvUJT0Ra34oTpLCcm+2yfKs9zG/Z6xwiGT4TSvmAT9sjc0sLS8ruxhJwdvHs
f3OEQKT5F8+ZHs9naijqp6tlu/qi9VYBza5i+xFQq2dx45WsgPtn47myDRwK
dmaVA2bzwCigaNJHtBUoT2qseU+z5V3ZIt3OE5tfXRXZFjVhz3gbu6I8V33x
M3nHrMfnZ7KtTeExI6JpK91n7JM+QWlvKIv0Mq6lQmodb+JpAqgAteKz+kG3
tcrt9GjXxC17mq4TcBkVjBlnPoM8MpLhfDf9cYOxvdZnKh6E18obBI3AE1Sw
GZlUKMK8CYOu8RnzwUhvSR6wCFrxsGGNiW78HJQm8Bia1znh/RLvak47YZS+
9tCQ9kx+DiHRzOPr3Muza/eEECGnrBayCTG17LQ1ZK0sKL9QwD8mD9eWGW5L
ztOR8WArl7170wKZwIIyO3pO4aeqSQZaV4oSJuB/r2Bjbi3xEb92oygxmNOE
LBk0rfK9if6htOQI2hGlPs8o8v/xWD4z980xG2z7Sy6gCjx8QydZtc3J7hW1
iQPh8ja9BRkKitK09vyLu+kE/UuXmlJYz3RDUQxBqtqzbgym/eSzhW+WsqR8
G/Dg2qtHJowC5xSRtD02cZy0hDMlPrjwHl6C0FFNKhfW6ih+mIDxIvkYNnXW
18RMBrQXs1n5Li2sBgR07x1cLyCTyOwihm1zA0kqrbA9dB7ancfvoOwwslw3
UiQDL6WjmIBNOKqNbqmaFV+WFmumtmf+dLOqaaR9V8/JZtm8l33mioZ8C3kv
b88RJyuqL3eqfwNxt3/2rkE54c3Xvo9DWX0f3W4EZOW4ruucmfKr0S3DC3O3
Ymglw5qDI+xEzNBP/o83vytgXpO402DYrm8+OvTsILFgyPm1BA5gp8IHEs4v
08+C1WYvnZf5NqDxh5DvQcsYbhJ5bZkxn2HQSNNZ9TMzZC+iw+2TVRPQq59a
EGqH1dMiT68IF0/7Cta5tJqWzd8x0Va+6jQ4il6TT5k2QMP5lC1kNR6dk48q
4+QutkKG+Vs2RXTH2tIjUAK0BL5kE7vQQ3TLyyFgHQXfOdQftV+FBvQPTl7l
wtkrD9qCOyUBITR+bz663AoWDbpOFPGhNQvAhjMBx2fQrVRUoc89w1HbkRk8
wMz7qjmbbVtHtjrYFu2Aj2KFleE2OPUAcbXahYzSUgqy2+w7cylAqeJ2IC60
8In5lCnudaxoCnNBeJ5ui/8VgNzZ7oEs9YAZIIlrFHcSirsTTMPxHuH2Y7Bb
czrggQL2lqVSaDv5Qi2ledVeOjDWPLfrMUQd0WYxUfSRVKPdWpBSxeg6UqyE
QgM40KKs0jYE/OSf6Zitb9WxdvykHEIpw+Wmgfm7/wfFVoSG2D2wTUiIdr6Q
VA2wIXE4GTg21F4s/2ou9bbT1TcZ+NCWf9VqzSIYLo7tZiEGFVwLCc9fnwS9
VMnW/U+9KVbAPMoskyMgmEzYUHtugmXLpYyRzRAueGHkoXjr2Xra6jmkEvs1
m2Gj7niXRxzDggqq/hjiCk/+aDuz9ieHdSQPtDBoPcpyYHOBvNBBzXqhHjt8
wE5g/IITt/OXfyT80UCZF0yqmWfF00sySQYQzwsGFAF+s2fyQDNjCCNRjMZx
dqrrpHhUOrCeY1XhlRVNcg81cR22CBw8U0rhOFmr8M6IEPoAm+HT+RFmMzY/
21LV1Ap7dtzyREayiHONWQ2rsJVNRwzlmbi04CiH/uEBYdmhL8OXgDpXYpcl
Ye96wVjCpxQ7xYa6XFsDDEoxsxtnLtn28Oa8vTzMGBba7t9WhTIgQWFNzm9y
m9fGZ4vvkbwObInZKakKa502cXstW3+Y7oGvQAMSiBK5c2BVrod3ChjVyp2t
SVSftUKUbMHCIsGOgP8nUdxcarNPcm94PJeM2lUJobq9e6ypuOvnDN5rSyP/
UvVV7qhIh+e7ejRErGJqg+AWg1iRmC5Lul3WIE+aTh7v86QjakLQiFuVM/lZ
0XzBPAuX4zDO+CSSK7kf8ODjMxU73RRgM5cw7xdBJJLfcQ8FPyWx+Mn5A+P1
Y8NH8w72aIfzVNhljJNwtcWDxzj0seYzxJzBragck9my8md4t1kRwP2wmsGG
8vF9IIT/g2WDFXNX42I3sAzxFh4lF79cdqRmZAnB9UDLxEcjdIr8y4Qcvy50
aOUwTQ/SvgpfPzABhp8SJ67IrXr/w3ng//WRXOEA2X84NjwM+BrBT0wKWjd9
DTVQwFt5zXSaEFRa0DhwiBZbNRyZWqsFXvC7xg+HwYFVYr/qXdfAx6BFkgQA
JGu7EYqCSmptIgA7UG8YBHem21ibw+u9VGGbWlMQ+8KOoubBWhKaeiD55WAc
MIBRyp8Z6DE1IngJ+atEqKcCIl1ffdWs1GndKIvNJpmacQ30k0sDZNq2r0gp
dH0legW9tDDpQ6733I2O0vVGcGtq9INuTsmyWeSRzY3slT6O0EzHpluqldCT
79vzo4ZV9iDLFE4I66NPR12F7PwDPf7rQWZs1sS2WnY7IpXAO56+3/NZPIQg
6AJG/vjct7G9Kwcd+tJC7S54mFT4RUsj/t0I+3Av+aENzJhKM4xnzfb0wnH/
lMoYwGkKpN8Pzl2VclsL9OqT/M9VAYTCW9ootcfkTSUq6fFnhzn0haoNcabO
KIF1xnIN53mOzthRLisIraGDSeA+eNGUNE+gJHA4YNOgvkp0u2XdpvM64L/X
T6dqUS5bS/DQ9MYLbIkg+C8ViG8r4bwawPNn1aIfqt327jTHYMDIwZbEwk67
meZHbLxRgyUSvLCR6rrzK6Sfyx1BzMw8Zp6EmLK8iSLklVl+BhPCamiMYDAa
aI0CzadyzBEhVIMdXhTV74PicIdJIOUHtqvlJrnluSXKVtcUbZT0ck6PkyJt
5s7fv/BjMuOl+ky/Yw+85DERokSbljNNZQfevs86frAM3hwEhdD5RS/A/UR3
ijcd/mM3ZG1GqBaYNBAw10HhE+sf+tyZoLC5WjxMoB2Bktfqg2fTz1JvhKdM
pk3S0imx/s8t1xdGu+mrYblB1MEKPgZr5grSjqS5imQJnj9aqwDcr1UaBOdZ
7aGPTwHtCq1EjMxT511xaZ7D9Y0YgYd2ddrmFWdqlxT5qxvBptY8PRQuy3mE
CnKk30Q1iecCkkbNQU13DRuw0MDNKvvGHovSJeqPW65Fr+AJ7pUje2X1ouOe
W3JRKn5zrmr/C0miEpuSHlv/iBafw0FPiSfHNzDRnLhE2sKiRMxNtEcsgsQd
zaU9SAatDsDFInGfONoe11ab9qGchzMe95ZG4zGnhgwQYaor2f99pE/jIc25
LzYq4pV8wWXMCyhUj6I6m2773JriTRFEkF9IYhneKdpRWbEwuB/Aqs27RzEI
LT3QQplfdddUzYxP/t/23DT6cUEExxhBKkS0as4gdW4mcjgW6dwCSH6sviB6
NBLMz1X191BXupkQK3jOQ7Y2TeRKJzz771FqGZerKq12DkjLF/z4Ey1Xih7P
NAVjJL8RBj2D4LM1lMrHu6rFzGGYwUHt3a5ZxgIxQ25ohTmVnhBjUMo8TfTv
E6CW9Vm9iWkhGCYU11GhrvvW1Ckut99Axjz1qCNK1apWReAeH2QJnsW1rOMQ
T7PgMwKr6VbEC109z2/sJ79d8bnQmBAKVKMOF7v2WV90r+R9ggownbDVuCMF
Fy6hq+SWh5V+RlTyBBi1GoYAhGAwuM9pwy5VgA+kq5q1TW0iA9VwgTZkEBqd
JfcVoWdUb10vQBay2n1J+tQ+fR26hqYg2cMnxr8Dk+7fumb+Wnkw0zhyLAid
Env8zMZIozNMLzlIR8DR2RRZtVrmsZv21V6MQFTv7RT7Aw2JGPVtJTDvvdm+
0cpjlxqUc49CXuFeke/eZjjY6lTOS9YygZG/Upp6SerKkzvZtzDIwxcQaVs8
wspxTMuSFaqkMZbR8iBbFa4iljJkjUVxJhGLo+ycYpAMgg9Q/PImgs+9m5Kf
WjtGF93dI/X/cIO9aPvvdW93VgjNuojoizmjoT5ipGmevI5p04CWVmLrfZg3
DOkHWyPPEZl4vu4UpecEQnGKBjSXPeUR+NAQ1YCY3SkgyeUeSGtMZtgn6XZk
qIUCBalUTiuPRqOIeUaIuBM/2fBIRMqdIJDRyFrJIz3P5d7g7uKjfWQp5NAH
GUaFCfKmDZb3V28bRp0ouuJJq5UnohE3D/Zi8Lf9sew699WQD7AVC6ZyevZc
tt2pLMs5QYyiDsPdSQ9/cu9+AVx8EJcgHpczHhqOxo2214wg9I/8+YldJp3P
PV03Ae6WuUjADM9G9nG8U56aMem/OHOEZ1yTaaGGrsEm2rrdWy3+WsA7fc0D
2FDP2uhkMAXdYa9Z9fLwBCcvPRLLcDv1/mAD5Q8kpcjfPPY3Cp3KdThh6HvI
RtyEP9Y4KjBygHGYUWEFPvaNcysDCGfEU9ukuJC7WaCCVM80WLJ080YhuDWI
jPAngkFLfdPopAMRW00BWMqW8uKnBQtGgI4aSbw9G/aCnIJf1OBQHsYJ4GUI
+ueNaFYRnXM6Phr3h4Zc0AwQ9Ao6zs+9YKQ3yK/ERGEdbgZEEZ8gYisriPE9
I2QnMCvIJxAhlRqtIGi5FvFVxE/8LGCJrqJNPsKQBaxHGLcbh4YdWybJaU8n
14QI6l0FlABD9Owdto1hdqeUNa+HBO7HWkFzmtDmpqpKejI4RSFgN9yGsS7j
AvVBuzAm6OTOFSZe/3pKya1wAWb3EBdCZAg91om2Wl+fBrHnySDL5EqC3JI6
UV87j+ovNyPUplxZdFXsf63F8nFHFfiiSOXxPC9xqQNySgn97AeuKYEohBrZ
WbKaFqhP8pnLmIZgnin2BAOjlkt2l5orYijukiuVqY1ZkuPQtUK0pLJuPqBl
g90ZPObM8W4AThSUTL6xiWC9lLg6PI5VzdlGwS6cOOrN23z6KBtFji8jojji
ydJN+3iAG7/ceUdaBIiPJGV2S2jfevT8hoL/m7fBc2Mx9FLAwOyOgKrS0+tk
STTDLmnBcYzeWXScum0Es2oR0QtNuH2H9aZlU+3XWmf5nlIEmcVC3nrLEzip
etAjvWPFP2fr7/h5x2WngeHB/42emODYwCUOrH9VlXifpOlcHKsEUEaDc1Sr
QUwfGsPlOTZ2MiLKM+0MC2Of5WjcXILY3Ax2+CYxUQqtWBStkTNzX4XWZ0/j
WBq6noj3+VRUTX0ZD7YQnDN5jSrY1VoEqAIEhsrupO87eqJ8lCaacOK1ccw1
mYK7Zbpby+bMdYbK9C1rGtG8detwzD8jKTAF0UA/cQs5kqPOfF3HmKPmQNNo
PdLcxCBkUfCvDIqma7iQ2hZiTSG4PobBifXhAQvquEAc6Kl//kZJu34grUBc
MwsDeqK/wbByp9QlBg/VAAwUaN+Z1sxEqM5inaQ1vnsHfC3k7M62Pq/SFuQ+
p1kwDLPSXQaQjVyrIcSFjHYMbfcCiiSua248Gc0yOQOC1Gdo8zFaEYBb23/r
vyUWmnA9WTHq5IshZR9M4i3X2S7VFNkjBiUUX8TQqPVWUgY45cFlMKCKxX3r
cfGG6U+YdzX/gZqDAwZtTu7NUht4V8U/kncILkOSVIfLJTgcTLHdO1fd5QNE
I4MEPkyguUeL484/Rt6f/wcNBO4pXYOGtCo62gd+KHGEm1jvl1RCj31MLXFi
9RZcZ4/WDx5KX2bMBfGfv0tUFEEGAaTb0wtkXSWZf7U7dRlLaVrZJdBJTExW
a367NPbi36J2qCh4GzpML5cAspoNtzs1um8DDpWb5N6yVYhnWEQ+U57XqeBY
t3ZTGCnbBAvecoJaZ2WRyFtrdPHhIrT1kn/6LNWHc48DQ9LZs1VZnyonc49j
J/PRNAWXuWpPeGBQYvQWSgHoQq6HcbKaD4yz6Og8T4s9cz3HJpskHKYOuFWF
i6IVqV4OufQYiPD1MFlHq/RYduilr5cKKsgNcR3tTUh9QxSds/EGE0rWck09
Rn/3kn4q7mzEM8kG7zQdLSjRuU+SBzUfUiWiOtGY0QqoLyvzFoj/Uqu/pWwj
FzcLlkSSb2kfk3dM4UZJIjBEOaDEH6oNg1uHCtxYhVv3iD3XHZyF3VmbEEQj
+I/DrbblvvO1/KEip6826QDYBVdYrzYgPPxeT6Y70jv8H+D0VbxO4Tz2p7en
A8Tjw0cbbAaxbuGZYZVoBI6Zh0l1qnTIugX1wL/vYoQzVFDTjxIGNdJxBKrx
KVz6DJYUXXqFhDbMYnhQPzW+uaDmFVI6G8GSJYJv5WNJJKFMxI6BKQeXA0q0
vj8PGXuvPkH2zzT+rr/gyX5qoFGt1ilnO3g4RfVK8pLY/G8EFMJwA4ONfU7d
8s7evLZuDU8VjtV+agJ4Md1fWlcnBY1yT/n9h8tHRqrKTcDterG1kZhzMuJH
nB57THAKJPOFBv/zpdlmCe+onuVpN99yfjPmw/c1US+R8Y86fCRajsURQo/e
gERW+WBWthSoFl8JaLyYLwxTIrjAOeGBgFlEBG5DTMe1JYPwaQF7cPTARmpm
CkWCfYwCNTo6L2Q+rHV/K9jlKyzHGyl2gw4g3A7RByTx4z6OUj6IStkAdlNV
BgKp0ldI7wwlq6m5g4iM3r/WduxLSUNHdHxQKdmEwcRYjB0PlJDef0TpERam
2bP0RGqLFg2q5NAkJBOMa/XjyP3/AnH/SzgDPNFElKaaohE9cWw0WvfAh8LE
m4X69j5qfYfEwPAXH+5Mqdz3PGLYl6C0eSJ1B3q8bDlV4oZefyfI2nwFcjIn
LwvY6E3alGPj2KA/voDR2u1qAi4jRF9ino9PmeiSRVe78WsF3ZXwoSYwI+3l
+pAwQxFXxPiRTq0FkijBXACaLAIU4dsMoWOmm0mXQgfi4jY+WVO4nKm93sdW
L9Du0hejSR1dS85kYa0JNc8U66/A8o+qTdU745vRmwPcFM5NSIhmmY7kFmtY
HdeRCSsL0ZmgVzvZkPKb5Xs7Me+5qsUrNJsezagUqbHXDu2bj7qSd0wsVg+X
hhjjP65bT7yJ1YsjC9jLaGP5a2CaxoX9l5Oak0XTrXQLhK9bmV157gEfTowp
/K4fJdkNkYtOt/HwBwjkmW1tqEsBqOtdeQQaXN2DG4T971RtFe6c7HjpQQjE
9Iw9gOC2Wk6OW5wJAKMBllfPYQVioCFkaSXLJwWrKJZbjiaP2oB4Qg+tv9bP
25FB3XvdMWOriCwxUX20ck33AFRRCs9mbQfQWRtLGMAKnDBnHSuMp9v0aQ60
/8V5ImIH4S1m/6K8j2y9nmQpQHon+8jRXaKlaYb6j0M89HX/L73cBefGAN0U
YJN/cbmkUQaBzRhdqKVzLXEMsy5jXVT7XHnAAgXXJvCpgFutsjO2dMNQ4Ftm
vIwIQp91iAnL65mCs2bM2fOpBVLpqRuFxlIX+mWJG6IFM1wLpn25wdjh4PpH
pUp1Rt3ACE5wPuzn0HxPajE3JEpRj7ERa4HaGCiBUzbh1CRfQqpRljQs79qn
ow7Lno3Es/rKcCoAh3PW29FV4jopRVyXniqoItgDDNE7ti5mpZyiaHp+ZnUx
vANznSBQU5WousnRalR7VSEdiiqADF7EwlIxHP/RX6fEJJJt8M8FyQYUIHhI
XlNUdxfFXh1VV0aQ/QTaFy4aV4ECE9cVY3hAnWqoIYA81d+hRi5+dk8YGK4q
sOwyh/AhY/j0sQC4dZToAimsH3oWLmnd55F8H3fbeV1PIue9xr6isBzxaLen
urMJA6j2GJWlEUOlIW8dMu1LfT7840AxDrhbBgSgMacE8J2MKGV1yistIrgO
RoRNTk5YrBZ25FOBq08Ptyrzwh8ojw/Zjlo6mbS3W/RrCyc9/XiKQyXHf6hg
qvsTWgbV+adOfDDn6RajtbIKoCMqe/acVkTKsZ5bdXlu+U43LjpvwjWb/ykx
5jqYQ2czrBpQ4iuhWwHUxA4ZP+xUdCgxdDPfBZhHjSgUhnaTSFCgwTm+wZBj
cL6OYt/Etz65Ke7REb1ZDNNy3U8o2m2PGcRyopmry26RoAQO3a5dkjF0F3e7
gqV2KWv39WvuwoLHIbo8AQF4gHurPTPt6hiqmapHGaNfj2FFoakAl0ZTZEJF
dG1WgLxeQ9fAWR4zTgDdrPXp/n9BQBc2QNhcP6n3U5IfjkPkbZQuOCHhJZ5Y
j6kqwBzgAzr9qgZE2oJR8078XEnYIZ9z7TxLXvWkdOM6FbIf2nkmY08QOuQH
FdKXY7vpRGANhCEwHwj2U4G5PNDGb6pIwZdfK8sgib3NR+rds/mxM63UAXPl
EnDA8Sny3AysqqixZTElerWaJv/+Z7+pa6WC8tPdFWIx16BNcrZ+5hiXRDMe
J6no5FqUPpT7ohsbePtZ1aKJMMX8TaHglpDvn4PWNp+hl2f/xN77SNzyq7Yf
OcWZX1lKEHScoQnJgzAG/wrxGHk09Q1NfZO+0PrRbaqEZ/GkNeskbLgz3vmG
4IW1C3+V1SzV4p4uNpHKKEHnjbUkungLjfzBDxfDJHca2zrwuFTyeNXqfmyZ
4nWz3SYfZoAq1+2kRPkUhJFHnLCyDNhvVLmF2j2EFFkl0zRcdujDDv9Pedvz
7KyfimzxSoitvb6LuSPoQ97Ef7/5b77EeJ+tEXBecR8Ud9aFg2SzezlKiTU0
X4qbNrquq4ef53pliUzvxSWal9JyB4UEtciG77qZUyU9k5IBbjH76S5VhRJl
drJzmAahSKN2jefJo24rDvNz95IDvj25KJwmSufnbFsj48VdcRzaohGAzU/k
aRhNv3EOP0RjJMpB8pJzajKiHSdp4ecsYvD4IrpFfc3G+FyFGll/vZdVdpiD
QjOhxksLvPuOJgNWA2Gab/HoSZTXfTHgjVsebX3FCVq50eIQ7elsURB0fEzT
jwySube9z3nmx2IP1gwviDsPTWdrAvYPvb+JUbd2g8NYNdeMq/lWrv5OA8Ri
Prn6NAGqEpAfTr58Ql16O7vkPinuVHxsK1cTXB6LMUCtT9put5c7HVidpPea
sU10qdg/WzT+uQ0g0M4cX2Pa/+b9zEiMRFmABWss4fcxHLk2wcqT4K+K68y0
zGYRaScmk9944MpaQmTHsaxBKUWTQ5oUk5hybxmUe+RCb4cnmYSnwaITwe0d
Ug7LWCY7vHZVc2e4OhGtkprjRyudSmNNDEZdWXXhYlklTxCwJi//sAmV13nb
uRLwCFmnqpPOaD+H6LnJGqCmOv/deY1CJlneDrZqyVAWr09pI+RJAzP90bWg
Xm/NpNb0/orNl83j5vPSZv5D6La+O+4bRlCIaw2XrnF+8aq3FDQV2zWKQtWH
pI9peo3JOW2FZYGhZFjhgoOvbHTqOXF8vYCFRRrP20KYCLF+UBvaRAM1UYji
olOSMqnz0nMUGJBssuk62lkhpIK7XkhiaToJPYYeDvfNjOf1YHGUbjlmmUyH
WXoeZnC4T1ylkRoRyW0iZHgmo0UKJnyu8Vu/x6oExFTtO2f8nI9FrbDTSzh/
TQUtX9qw6pQeJiwoQn3aCw4OHHLCOxbOygAg03WLjUY6ku8gDqOQp5cUUBqY
053T7kD41rMGbjqUGrUTCNpz9nvMXkVZ4MvSNWULSJL+3UdUPuwdX3+X3nCy
LdNMnZBOulhRsRlXstSEg2l6e3WyDf3z+dUGmbOOxYZ8Qvc9os3t87FkgMXi
e73oPPUOkNOCC8/YRVZQK6uZJreG0BYg3jYUL3CUR7+0Y1DvbetQWrtMEcot
rdABw63oNtOU1VzeIdCCsZwq+BHHRKBJKoXMVuazcnuWQnY9qhvmkixT09a3
i7I1EQn1DHp4l/WUoqI0AIIp5S0J0sy4AOEZeIPha9Mcdh8MxAVel5mq0xEZ
JVHgbVTmk3j6SGU0YWGGMGVX3mFsmFXwf8Df7dqvSU/dnLFKPUXkAU2dBinh
ZpGfexFLMVZZSEqdlo+ITxDvplb3yXi9UnKoYmog3LKuye54SQgX3ZRB3IMr
kjRVUkPnVVgeCptSVb6eY3J0zn/2Zs4z64EAfco18c7ubnPM2UBKRaEnkWbl
zvftOESh0sgRg/GKsXLs5nd7CPxVFu+9LQ9gTdC10CEFyTNDayeQfNSDoJnW
pX3bRErZr0kSkSjAANzTcruqjCEagE3oyDuUWSdBxg63qBvutfHt00hy8neA
8EA+4H9MMsqqK+hDxugIuQ31PrrfK1YajJ5vV/36dpn8G+6RwBE4d0Fq59k1
9Jaa1M7yFeRXd8Yevieym8dJrdcxTiocgBJCby08QZZ9q4CM7Ge/FLrlSywo
jOhU0DiVDiTyERje4pfqpRm5ZW69ubY0tmVrH8wZjfq4soiAredapeP9qqTS
3Yb8ljDmmPYCE686Ph85oVo99X7bguRzMhg2R1GA3435QsncTFQKLnQ1nYhQ
DRy7TqUuDXOZBAZTopO2lakCdvb1+RhtCobKiz9dgE22ax/+uLGt48i6n6FJ
n1DpaGw5vQK0IGL2bBhB8G9yTRM+6v0xe7MAoE4ohYHwuQ7a1JQOU0K3Vex1
4cYg7m87/aPz9T8B2rec5jYP807OmBXGvIhRRLj/65QfvnhBrmuTXdY7PmWD
2+ZRDdyMxa3aF03guTPNkW6FkGBK1KDz8t/CrfxwdTOhIm1qNEW3AhrZ4Ca8
ej6NgC67QBv5u2PD5GjgNZphb4xZC5Xxy6Cc39QaF1TNJdQ1sOLGQ9p3u9fC
VwwwXrlzuilg/x3D1d4X0mQBEbmeePxAgy0wBQt1vddI8Nv+Le2eHXNPjQTx
OfL7sij24hEOoTPTJ9CvW1zm3kxhu4T84OtYQspSUESVSTF/1fM7SS1vMv0v
y7YaeKffvKmQ8U7Un0EpVnlOa/7wr1c+3WVDZ84jxw/aoNnXFHyOluF3+fzy
TZ5z9abfVIgfTWQGL8aF2+IlGvzL6NcZPIl5lPeql05OpcYwpHWRRyNRgykv
OEdcRgY5RKJ8ZGn9t7z6XiTwNgciakg91DzY+nQVdt7ioUgKEHKqSPv2Z+Ea
C+fsB0Bgwl6ubKwDOnMyd9bMoEKs8vR7RLfSakko9lSYybA8drZ6N9xv8+G+
SSFetYtBmgYK4nihgoQlbLIFSKe/GQvDi6YWO5UqDGyGu6P3QrtQGnpuvGIw
pLqcAqGjJ2OxGFHBCOc4dTuVf6tLTaVuDzTiL3Lb9qs107h5jepiuwAfbUy0
tGYhBIOYYbj2UDzztBvW4SlOuPMrhxbTG+ulmyqBujqcyyw2pPwoEZhcVv4Z
zVT6ChDy312A+6R9O91uxIH/y0+xQzhLpSoitDIl2v1zuxPjYrVWrf1FVmRk
MHOAyEvNOn2D//yk/LM0aIOMFn7xYNJC0JD9hxFv6Mn1Sybqpsjj0UVIkjJX
NgVc3jPnU7EHeYSrUylI3GHfyjjD7l8hf3RkxRXiuqnEzqqNCU3Sxq97Tthb
WJ0AqDBlp5qZguFpCSZ+ZBWGBHdKDk2cn0AnVeKDuxwSx5PYH7GFSBh4Cw9E
IWpok7H4Lkp3va0Bk+wqSFFEl1zpgM25yiaU1402H1UHVJ0MEFilkJyfjZeD
teTMkObavk5DC9E+8XSnPcmpJYIHJjrr5x/TthMg0+FY2MjweQYRXagOs/8t
8H21LIhAGvThGugib/0MDDrm845U1b5UxFRsoCCgxk1CwQePJgAemilb32iA
uMAPAOGztJK8FJ/YGkFH1o2PlOQS7CNCgXHarjWK/zCkKnppp6DCAWyTjaJ1
wtirLNNZEfVsKnh8HGBWkfvp/ZpsQgBwsL2MkrD6SUCHLLSUDaVNW2aostOq
cGgL4l9w7BMfAmfyUS2qrwNoa8Tvf5VHxKkFWBapactsK00eCV9hENXmid2C
/iHUkHd6MvyKAGdBNLX3O+c+rg4tj9ulr5Oj97RcaFmBdgntIWXx8z8ShiPh
qapkr1Vxd48THCEkkXcQoHEiqnixa1KXln06qVaLifFJt0ONnp0mxn2t0lSW
uF3RojCH4BS1qPI2/8me9C3Y5jG7+xW4TN3KDOVsMeg6K5wRaPipvRllSO7d
JPFsfuEFq+0iv0E65pnlVl28l5QaBOP84suvaanyS74Ajq45RjKAjkSGC34i
3gYNzHA/jSMXIZxwbuajIrJC99DfaW1h4FT9PepRSUbJuUsWbCq569wAm4Z7
CKqKHi4egOE5quVVMcwP73jEaIdWfojVepN9wsJUtiprr3BRFqFgKvUNxzCo
ztWxMHnjRVnD6ZbCBW4OD+yZCUziLT7YrMpg4aDtnC2tvfKWSUFPkAj3ENhV
4s7qH0gHLdivHiUdFVXYoT0IUyYmE1ynpO3xIU+s6ebjB7IL6f3xZ+0KyIxS
lVPpldKJRO3UhyyF+sK9JihqNxPMpex4J5YpkHD+LxLCblMMDIoCv6b2sGdw
Lf8Or1C9/jon3zbIgXuXWSmunRPEO0Vz5X5rBrwuJhztE5/5k4axL8R7N00d
zIpdgrxe1YDHFmLva2gRnLVTHFfg1uH6kW4CFnwtOwbhoAl6z25lg3sdiqsq
CWrurSPDZI3fpTm+BbRKJtpIOAjh/UQfZhKqQeecTPjvS1tGQJ96G1zo8TGR
uU76SCZyr7w5Yjfid1ApnD1eeOYp+vPu6MJ9aMhIpef00cMTbpvlDjRyHode
Ezsqdx4xZ0dVYxkwOWa2z91CuW/ywjGmD58rSJHIrQ9sR3ppnwIPnG5bsloS
Kjv5ofDcYpmWpKV5QFJVhFY3DTVFY5IaA6Jn4JUkBW43/DMSumtSKZTjlOPK
554XzuP4eBPxj1rWy+AbqrEtlJ/Iovse1BsVkxjHFbJdQBx1vC+Um90c1j1U
3iDB21sAsOBg8qRdDoKCPV9/Ff/Xtd/QN7J+s5UINv1fYrvzfcNbmEKQNgUY
0kKHSJJRrsHmQx1GZ/n9JESkc0bsxe8+SGvo3QdOgtCo2xqPISbP55JNSP1o
fbjFthfpPBVA6g61GR4/a8beoBREHamvi1tHhFKq30qd3jG+UkGGZ+zfGN5S
fmjgHsoZs+gH8tqR+ekEeRHIWBbTN4fkzAg47+5m07VE04jf63j0Rsh2Zryo
A4h3Pe2pgjDM8GgbhqKb0nUcD7krvq8EzhTP11E7u24kAQMrko+y1HNb0djn
WTIkZbPeDG+VOWO+G/vc9YgDhJWLnTsqahnttzMphGcUrwcuWvo2Y+RqdJmt
zt2ACdOnmCwjn/ipnDYLR/K2oPz4reVv9ezNM4azI0STSaniazmJeMotp/ab
NqvZBbKXaJ6UxBnGXL+5vd9zveYl8JOktzSTujnTmwR42NvT6yy66lLhzQmV
E6Pvg16qB+F1O5ZdQxBUpqoH2vvW/dvKB3CdY5X3tD70+ejDuqlnDHg46KoT
ETBqowZeH1fH8UIlQPnKZeB7BQm3acVsHoO1K9rtIBJQMmD3LiFuvfGvwYIT
HN5gD/4xyHv+4+WSCI6PEP3gXGMCfLU/wJPvTNOoN/4HPH7Po3h1OFeWXK05
NVTyIp/Y/Xput0yMEYfgTogdtkrl38rJX4HP0ludHN1ICdlPSbMJPFl4vt7X
AxVtDwSe53q6K1gopCgBh7/4p338WYR5HNXI1iXs79tbZtcklq9i4QyBOH9z
oP4M+0EzZFq0yUEtgWc8ULQqsLbR5WdqDUt5Bu6zp7/AT7CfqrNcaeNLygo3
1t5+HSA2ANtIMZK2L2KV0vEckpcsxc7DUP+fqSVilYc2yY5GSWpkKiDXaF7w
bHYdgqb3S0eoBK/mVziKkbdfTq9AloPpJsjq4WgiFJRr4CR52kBbhXwbPHh7
eMWumx8FeeRAzccYRGlK+yRvn7SplACHe80AN4WCdqf7tFgFeRIkXl19YbpM
x/+3+glAHZZTYPaU+rmXCW1vb/x8GrFgvntfLpFEoCNEoI57EzAJWjmlqip5
boFBqd4ZxwWafkzZ4XW3nUpY+2odTujEwud+rIcG9M5RGwluHz7uV3XsF2gT
w6mXKZ/b3gdGqWaO+vFEb5UPAc3iEsxXuIHbAAKW37rb/G18DgyLYYtcKyKa
h75TXSUNJslWoS3Jv2a0FeSgs7wG06sqx0vVBGIdnW/S0ormwR3TGWsJnbOg
dWdwOUHPYTLw/TxFrCejlHfF4jmSKDf03ntp+uNNeL6eZp+w0v1Dgh4P3RGp
GCXqxXJAjAXnjOuDEw3xru8bGI+O9rs42fXsw1zK0TwbSyndOGVcTbfaDFFP
fZO87F0Q7VvpweOIGGtwWRn2eeD5swJ7uwytUPU+KVhlVerKpeQA/g8xR1XK
ZXC2TnwJ2oStXiuFurkfMRYNb6+bN7kyoNKNnf8Wa7FMN8fSASprt29Q534q
PHZrgPeNuuGUG9sQ/IySjJv8/XVJJ7xjAauxlIAMJ5ry11F1XRAsC1/MTpIT
1wOwPc39jmpKyHVNMT+grUv1Q8k7QKCNtBAUBZr1eKfLnpHtenTTIH8vkqH6
EeLO5KVkcI8Is7CziCE/nSRz4gJfRDUYHuhZSl4nqaG7+O6YGD/edMeLy3G3
YUQU5nWeJ0DWIq5Od3pwAQXQforvwsRoxXN/YZ9ZJ+U6H3/FvIeptL9reCPG
riAnkRXlQxYx/vBwlN9gjzf9D9sufhmcCNglNrbdrcxchAFqxkAXYjBNcoxY
ze2VmEtm8mRUJcmk5ca9XZKYPaDOFihP1CyYimxnk6zwjxM0NUSiz+6RG9M7
WAYGgctEbV0DsXMf6HZW+HRTVadnRscslRJ4nxz3+glgucHClouiKVeMWg8S
vq8CN12fk7OfP4twX3FrSf91fFpeZ8fFHcfeBpCuaj6JsU5b19D7KAs1Gnsf
mzlAND6AueMELVUdNf/XSGoUoasItf+doDFAcX5zC5Ewz8M52eTnzaEu91/K
TvswtvYGrZm1ncaJsHjaw1em0jiKWAZdZNqc4GobdElnGrneWLqWLd/X2vnN
7HuXz4hTUNqHUFo3mffVOrBVXQCt8gSZJt+50D3XfhTXdV/HaTjlPCdi1M88
neRgAXU+d98yp/5fnwQAW0uXJk/qTBiiQjMmBBnhxS09u8aM5qRTcojUL0wx
0JDPldEbJYnBjv/BW9j52AwQrCI4F3o7ZKvDlI0WO/VBTrjny/b13CukEzst
sYQ/BEAuWooCey8i7ZAo8f0NpDREXjMQOht7YqhrY1berXXi9evQOT8UsgIc
4NAr4LXbo12+Pi54fJiSif8HR9f9RlmOjKFZltwi8D+jrTQsudCvBtmNGjy7
eIf4ajjssO5WnqnUPKKxDq9vhICeIUjKW+Dpym4ookHLUaEFmSn9Lv0u4HE1
COPcVThZ7JhdiePH6g7l11yOnL0ffCt9Sqbwr+jKfYtt5DEwc05LaNySP3hW
h2+cgfkzlsaETxzY5cWkToZ7lvO6vs64uvzue3Zvl0/qliE1yEhJYorC/Gzr
o9+T31NkgDqw4YEaVTTKRtK15rEGYgrxw04nrnF95k4QVl686hyVIqX0De7I
iA3mEnz8HL2EKH4osLIurwDoDls6lIhY4z8VagWNWuYvY4i7rzqozF6NHPM4
hAgwy1tjC2a36XOiK50aoKS3lrmOxCrwO6d9I8F7Fziw1+KWNC7jBxBIq717
ITBuZC3dLIfPJklVS72cT+RymXlGABsD8i/rzX4mTlz1gNq3dXajdCOcTdW2
eS0dpQ4eTPHllPiPBoxtBHMjKdHNScVXdRP6eG5orC4qPCPOgURBTIE9pfVd
kw67Saajb+xaFVFtd5aYHV4H7mPGopf2UdYxhDTwpiWgKbVWrVHAmZSzTxET
xKtQ/YibziB/dLE46AFakl3OqcvfwnIcopl9o9Ne8XbrKSfxrxQfPirktPHW
nG1R1pfsTUe7mBER7sHp2e6PJMeQpGV93+C2N5QHrGyHHl4quUSQ7nmEcYSk
4gawHwzZfEUccLp5D2o8Qp8gacXvKpaX1nmxmW6sOq+WqV45gwN1JvlfVa1z
DXrQVLdjwMDcC0kwISK0myBHNhWXhOv0Hjf0coBbBEhk4krbEZEAlROC38Iu
dzPwH8/KNm18Xkh4jxq3SUrhCuIeg6VHHghhconqPWWIUJYmQ/dIdbiJsBYg
BJq4U+9YtKOIRDhuifQhNMoa86B8AM4xZQKX58HJaGLpedAHfU1R42gtYx53
yP0L41UQIVuWe6VfhJurk3nTNxfA8H1FWXqVJUMQwULQlOU50PEfcNhctl/9
xp6J1FNSkvszBnMETvAxALgYow3X2TTAu9KyQWoy5gmQ/5ufrwP/tl75oPv7
rn4B4P17F2ZTWr9nzPtBy2AghSTbM/jd2rLaQd5QxjtnihWMu3ZQgBBtOwWY
g2NP8p+11t5HdGa8jjEcBnAB1oRE3YFMQmScnKDBRDajOPwuXxrDqciAcDmB
aR8V9PT3EBf22qIia0YGJjvdTbGI9AyfSEzx55IUaZ0OAlKqCgOzvoRRIcRv
0h8jeSRYAwBw2l7ZHqLjPCXttMk/ItQOy8fakmPnJaKRx8dPOTohxOhBZuaR
ihALU0ThGFIb8mRWwG21dC5Q2s2cga+LgDWI3VFiK2camshVuHKkfSU0QOZD
+UswNRpvPBsILoAbW9UmHBOHnCtOcpuO3Qsx9eIl+GRi9O5W4FBM6MjWxLyz
3AUDEPXfgSQzJ0MGJhLXYzs7L96vHKEa8zwa4Vo7LAxtrOV9xhoSZBBLF9eS
2qFmR1A0nu9aw2vXBXkiuvJTN7DxW9tpVm258QrMePQUebElLUOI9W9FRItp
MHP6dWQKadfMvpgwJ8yF4xFlgZ0fwEurTAb0HcfvlvXRRv05T77P4YLxlhDE
C6GkmUYZKe/o+DtNMVBk9Cc1radHD79LcS/7C2Kui+x1eQ41Js+NhoWkD92G
C2NmMEq5FiUDpVxC7aNUU82ouXIuDeNaez1qR2hbFVGi1x1rIAoGepzYy4u2
mfLL0Gbo2mEKFjfpt18kkfbW3vdTv8xdutM9hsoCBbcuN6A9uZN2dRNgGhBt
NFGz9Rg/kG3YEjL7Cc/7giC7QApzqf1VgnrrsnIxayL8YERK6LK4la/aoFE/
P8YK3c3GjCNGYc8ica56TcBzPLYucKAcj1TqJ+VAe9SUuKtvKcRm1a9zLqNd
9ojjNj/abcRMNJk2iVnN4OIJQYHSU7yxCr2DIQfjexRtN/pNTaQjnlJLuuCA
ARMHuFZ5iBEeQraV8ODp3N36YCiEpsFy/cQHqcR3c2RiZzXWhI6XRESUBV2B
wtsayKVgDJYisMSQyDYd0cZnU2gEv0qlGjHTCI8TY7tnb3nztP3ijayVUtl+
aNM0C/+WCCH6ruwdckp59rzd5hRFgkrmUsv2SyPH2rmd5XIe17Jz/jdlfpSJ
kU+F9f8hiRasEVYH0rnyz3TfnnhPX8naG3g8WwB11jVXHuY3rkPELo5tX7o/
WR04Zh4eDn/dvvAMmq8fSlWXaOls270nvy48dTsf7PxnpJJYfLJm0v6wYU4D
YZUOMlNfK2J3bRtRgrL0kg2CkexfUT4p4cYAUwVAJbgPJ9T+MsAW9PstI15R
7gcHTWnPBMeMHqeC7g+r5Asf2JWGz8g3Ul8spCUcbh38DBgcXBZNzjKzn8Ud
EPbQZKrkkEoTWzS+wZaSEPzHq00WyjOgQNGh6TuZo71n52tGjTdraI82jJn7
9lTN38V3qsp9GU/279rOTh0USMG+XyZf1PxKClnpX9Ao1fm9YhgoBDCbvMbH
iyt2HKlCF2EifP0Hdifj7x/ehVy82xX3jHuvpVFTCEh9t6mwmaU4K9yxB1+o
zDWejIkBekxNDITXTqb5qlxyZU3fgJFv2w1wFjPz/k33bIAgYrmkupYJwfjO
gvs7e/1/fIZoo0eKGj69kf3Svel4PrDCtaiupy8kOJkf0w9UQLPBloBkOPae
sdGFuTPthiZ/ucP22MjanGfbFNi2650wPNGEWMjJj0dhAGDMyd9ZsPcvmrGs
eHZt7feN8hS5/DJcOabgel1e7XGBoGCm50vEe9IkFyLgfL4s0LjeiTJjU103
jmv+XRSyyX0irQZu0vZhrv4gxGSlMxfrQpTmgNTlMIbjHfNS/aA3hKvY6hio
rQy5eaJVeSGyakVDDZD2wwEsgyoe3cBoS4Xrro0qK1hx5PlrCstDJmAwtOtz
uzP1czzDKhyQ2clU0lnbMeM4GYK1jTOB6/w6BWLSVP8pdMK5MSWEuvGYfrmb
EHhiE/eAEVkqvgKUziROawKPGbCpbOiaHOOs3R+baRJC/6hSiugH9JrsCMNz
sPT9kQ8PRewvwqCnxCz9PKTQJ9iTIIV1NBfCis2f4MXOup8yJp7odBoXacQJ
R9WbjFrvLCFtVkAleJswrWAf3C7prQdCj1bNtdRqHXrNLgOaOCpWGAKa4Q7z
/PtC0HimQxH17xb0j3jv7TRZZXn+UJ/QZ/GLQgDVrRPq6LathchhRGwjuoDT
5xH58WgpEesn06RXz8/U8Cd3bA9ryHryqp1XruL+N2BAI+fQs/6EFOCD5qqQ
TGB0nsBanxvMIj9VLyZf7Vfikwm2jktwliG5kympwmrFI9ytKD5C22aVE2K0
HgAalyXvrucuSj0L9pEOEND0itU61sOnIRrVFZn459/b5WFzMmu3ehhQYsMg
TE4oMEnk67PtT3xk33fp+/JCf3La9BKqI+nB7J8hcdgvZAui5nRqkJg/Vjx1
BpQwyZKu0tisfvMgvyQwglqaI1uuJfoTz66AGR657dIQbZs45YpO1rBynQbn
L8eI2aGA5dwh8JghNTD77Azzi7wHenaYSIjBTXAUQZnvq8Dolkk70/+qxrEx
yQkJLECg0ZAC3UseLJIXcRCIsvWGSzoExB70J8of1eWeRJYkZpQ1GM0QYLuK
/aAlwEj4jYlYq331uOHHQu7Jt4yokPSyzUx119uREZPRE/dDdc5Q1zoaQR2h
XLFiBNWwd8XsEOQgzRWXox/0fu9g5/N93wxcZhH4Lm7Rdraok93pzlElkw2+
vC5q7M+fREWLO/khUzvRMvOb+9JiYBKRUPiceLb0j+v1p2J0Yf203jm4HjRd
6B4NUcdRmeRpm31KzksyDCQmFiTQ2p/ocMuR5SfUJlU7a7ahoWMkB+Q8WvjG
g/VGxNlwEEHkOR7N97iEGp0Eu6URSqV7SDPVMPhaijFtNpVizG6E5goX3yix
hsYxpdUkk6lvLXipATHW4GubU1B3zGvMcvHz/OtrqKu4SN0yjLlfgB0FrQ2B
e/EufSAbtoMgDcuAr0CTtPcgWEdleL2YXS8lWSSHl5o+6Ng1BT7t6YAgHwwT
ka/Sbx8STIBZ/W9YSaiMgxHVbEZRL9tSWtgvcUps9TVX1UxPHPdFZQOQ6Oj1
WCA0n0sGRftqTh8Z2nTpxnW9TGnIQ1Yd0r4smmfnyZk/I05E479u8lyimnmw
p2tlQeMUfoUhpVltyD9bi49FX5wG4hVfUlJt5Dj57iQujlt5lO4R9GnIyMdc
+6fUsZ5OiLIEcP9FlKzQy8/4NAoCPs4fKn+ujoMquFarRrzTJDJl2JexuXvb
cplY79aAeH693mDz1Lwwr9iR2bqfNJC9HTpGy+YEx7BXlHrMZ+PipkrJ2gKr
t/qpSsJVmb40xvhcMb0tn5d79VgRt5Ix4Z3iR359j1UvSo2UBW1Azvi+rx6i
mjFeWjD4kabWwfm8NytrN+inR/lLlDBQDidVi7nKm4T/hpzZHJEfQqJQbZ6l
yT1PF3KnWLwQJwbaLtCOwn9z365Gh4AUagzkm09tvaJV0dinnLzVqPPZJ6TC
Gw9EFA91hu1qCB7/+8AChYIbNGfWvWy0sQ8ANgKtwGohxpDc2P98shXNPGrg
x8wvydp9pscpudwSIPK6nqj7RYwDhCmlg0RTXD049dAIUH59S5ih3ZoDCsus
B9a/M0HJxCQg2D6nK85WHP96q8jLPcP2nWIuj5/3/OuhQgpPjO6ORnyy1sl2
Tqn7IFycDXLV5f/otVLfpiEmZJfwZR9qLoEFf99O1FexasOuwcxQI2BtCyWv
IVtuijXc1mblhpJ/fSwTI3T3SxufObHguEDiUKn4dlBomSVgYtvMCRYBpdIu
pADE4L4nUYM2k4s6QRgqyzZPXGKODYuLejg3MLweu3dXrVfGVwERX77HpWzx
NNDfe0kbvH1VfdmFW8irG8gWP8FQSHKfep3G2Tg1/p6aKILy7WvOJO9r5sz6
vBPAyUY747+VgX/gbma6JN45VRL6ve2i8hsiPNhBwEfqNmm5jPMW2Fw1VJ7A
gVnp4WN1kR2pasQphn/waig7L5Pi9isiJa4dPT0BOL7bZzr8218EcShLLoNA
U7EIhVktbK+aCIcFn4i3isqAOCqN0Xk5uC3+axAUxBczbSiGNNTftXFTm484
NABdcuCtYqqrd6uaYb3HtRiIWizrqCM50Tlp8KzUibkiPHQrWdWB5CgzwhPH
m1if3KeS3gBde0uaf5L8shrkMiPK5YKG7xvYnWFMP8WKmtNfsHplQCPsX9AV
cRdl3579Y8ZbuvBxQvfi+5ahHRV29aZLh3bT0zi8LaiBPLzV14QfOOt8xn/V
8SLgNoGjLlQ5/C1oMuM0/RAQBb3KdQpTkLvLNnLAtXL1SZ+MsL9eLctc193d
orUdAca956QklLtysLqrKqHKODGchjXxkaBm2Wa4f350sT1JJI2Izr4E0Co+
tDqQUMOrQWefXUqQAvK+dxQZvXkSjEVBrC/3cMOGQohnbtl3FXpKoXOW7nZa
xdnj650YFfqbtkiOZC1eMrfy7CjGyapaYxXkeJjp6kwLZCf2gaOhix9z3zYa
wVwenjnYbxpLGZI0o6kQtg6h7spOczbmy2aWvQoJI3p6eo9yYYPVX8wMiUim
PW+vAQUJY4BGA+UYx/GBy5yO9XKLmpzWF+fxbkxtdK2Pt8+t3Uqp06qiN42d
AchKJYAmjUYkCw0xYxuKLvZ2U57r9qro9+ouOxfuuXhrR5Xk0JeeWhJRpYt0
YmwyyBfyxzGgySb4LyZZuCE0gMqvwbmA/Gf9hg7338MB59bZ/zbhxTMHNm1L
L+igDjbkgapRETywEm8pIui6Q84n+eJLbc4fCUGGRtZrO6VDs4hoB4/yUi0c
dnNvzfAaeGWLJfuBZqUagEZpcacQmPBiAKFw/+ed9tTQhP9RxKk8tLG2uoQD
rv9DfnC7DN+80v/SfyKk2YU5XajdpYhpBJxmpTZz8xj250sMNxAjFEXMKzQT
1A1TdwMam020YZGG88P7IJubcaMYibGNxOrYjn7CsOqbUqiPuEgPko7lBp32
Ww7qXsezcbKiBZIVq5ZOIqgADU95Dt79sH0HodljTBeyCGV/2TW7TwvserAq
yfa1vJbhdBnzRpdMOlaBXoIGSlGUllaKp2OQXDNVedVbpQKv2cXJXAypFMZ7
MBoJgqE+gFCQnfKIARFQcGl25kBsFm4xAalTTVXYPWU6K+vXhDnMC2OwBmwo
C/FOMJsza+jRhqptgY6i31ia8VGfCqHNGVrD86oV+Hw5aTwpsL1f2EU/Ow08
OsxmwtODX96GqYdrDD1Hpcs9a2pGUzwMgCbk74K+YfkXjvyVAqv+RkMcBZ44
9HhA5jGDkO48AJPsHvfNdTL+hNMuzo5unOAaksgUXsjDamroh/yeHU40axW4
UsT/YKC+Oa+iRUH5Xs8rpy4wYLMaGVLdXB9Eu3CEKdo9OpNAgM+PAlVLWMqB
U3HV1lN1PZnLZpbOAg/Q+v6tLTaaphGFhwBC6HRjf33VsrDcE3R3bnqnFDkf
b/msA61qOipUyY0hZ+s0U6z0Kuf2+4NXSrTM3TOdwe2xlfxE+YE8xQqRA+1T
tFgDf/J0j2RaSb6jdqyx3TqeYKwtNb71/seuuXsPgc6aRJXTlg9X9pUNxw6P
Ga7KO3o0PLCezZqqQ573E2O73xuZ10IZgWP1XdwiGMfQj7Hrh2S3Wusw6PlH
jmQnRroUKnlVBKH9j74G9wt2cMweS60ZjOe7yPBh4q4PzWmWPbwk0IGIxgM3
1CmQ4rSONUKRJDUJPhgEfkENoUSMR/eOUF5xQOGYI1psWfboqAErPNbiDttA
oQjaUl0vLzbF6Spk0+PKcHgMtVTaWBP1Wb5dSQhe5SlAdu0xrtRnsGfBpOpY
lKYVxVUB1ppoLjj4MuwKeHkTvFSvK6QUNAfW0AfoVezz3/SSKUlYz19a9gxX
1YPgc3KiNN/NTFQv3X8Hzj7qZlT4atGISg4NCHvtpVbYRjm7xy6+C39pdeQC
URB2Pu1dbT4dL1/AAk2UcD/3Gr13CxgqGHqMrjRf+sKm/aW9yzNnzYyOu9I4
hmoo4/v+q/FKTHQafVhY3+0QhTmwWDZqRlrbKWEJz4Vtxo0fvz4ucSR0EQB4
UXYj/KVTUYvGpIJwnKcFCqECb9V5eOT1qqLanztzvOrhpelA5MRfBNMsS9ri
dVPg7dP0TcyD9A9r48t/ZjtWVDvbk6+squpSSvDZq6z3Q7c3mXGj0c9RXZBp
Mh0hBNOuldpWWfTDMONNvrQkSPhKeEWpDwUjNfpFLJbst+QJb6wIDdQWfCcb
1FLDfH/TihCMG5shnxJZ8FE3hdCvE46gQSYAxVuQVT1nZIWnEZpK/WhIN+Lo
206EcWT/pm9mdZ/u5qvKG1pYZn+yplvUk4d1upxdNV1rXqz4UnW63AJjgP2a
cY+0BPXLA89WO0HRl9XWEUAyqDP86IHJXxKg5037RsSdEvC2D6IfsMQ2eacT
Ra/z0E/skXxT1cbsP84wD/UbavB3rhNy7UHGQwUVb+Jx4uhaCAf8FWvIYLz6
54W+OeB5QTTPmqXMO6V5Jw42V39qXX3niPLerWW7UZWluJOYwMuS6olleKUc
fn5d0A2cVYEZlV5D/aMbxqSNv4duHQmbbWSZCRxHjae+YR2aahivpM9x4F7F
7Pk2B9OjRryuIGjGT1BXvAt48XeqBIO0l8P3g2rEHuXtwGE5RD5uMe/seINc
EyaafVhbijpDglhdaGrakBz3I6CwnJHzksV6cBlG268HWHeRlKrEsUyJwFHC
VTRrYReq8VCtoX2N6vEcExqiFAR3TaK1VVkH/IaarUERQGUsbfEt3Mq60Tiy
I8DwPF6K8qsaZT6OrudEaDR0hSca4sNPjdZyvMEJG5Ex/3U/WfbtWCR6fnL8
3E7sbnbeSq1AoOv+Kju8dmXfz2UyMpiSe/cYj6aJtVZelKwVsHG1wSK1u/qf
6JSyImbwM57fOuxMjodUAzzF8p9C7QH5Z8mfsq2Uo+MxIv9F/Qph3mWUbJCt
1+hX/VfAYgyA0zByc6OKEpFujXrIx+tzIcFRYOJ6rms1dm16HsMG+rjDpaJd
Gu40mRc0H5cP32KvazPnlxtFbCxN0cQH0XOeUK8/I2+vC7Vwp+aBsfXZF/6E
38OPG4WhBHH7yxf5mX6sSjNgxDL9i1HA30f8N8bUhpTRAasEC5VDbtulbCfK
1yM5RcTuyd4zWKRtS8W5O2T9GzMUZG8aBq9hBh5pamI/NARnAWqHKcNhzRwf
n5NjsFoItyKt8ecEf1j89cfvkMCYNDJ6DdAWYe9liQFJphWp3JSFvCkWzuL4
4tyV+qmk7meeS0MZUmIvu4kxpQ19yM4+PKF4gclgg+UC8+BvEN++y+mNUSsk
n9iyYIPps18A8fdCwubbSUSDUt8RpYyUvLLYK98d3Yeh0VqQwYDs3WyrrW/3
EYIgpFaP3OC0eo8kpBTyOrZ+GssRoj96nbvdDoSO51bqtMxuPJgV45hvmiYa
Xxk/9CRy+0MPpo7nynj/FODpnS6BDKzDMfu4D4fvlqA+dIg6+MsJSriu8j1G
L4KuqErw5NCfsB0TiSBNAuPrxa6Or5fn4Q4YY6By/WUbDIqU5L+AfP5ywKF8
A6JPSg/4u03b2QBLUTsiKKV4+wdtWEi91h4dpQ4H00BjVBj4x0FOwqWiZVTd
atnOoycOPyjVGpdeSxUXAvD1FH7tOOhoqS4oCJlVa5owhspSOLiB14F5zh1t
7TQFDjfkblclWUEDiuo3+ARgYN+mNXGqtSQVw+/Ok7KNE2WVicTqcCOHaQmz
SSgttPYkNJ364JCfz8i0F/gbOwdCeLcNPr1CF2tgGEH0hp6k87szA4WGmmJV
MXXYNWWocWuiZemEo0+Kl70DXs66rRXpFdtVP4tc1AV79fXExyVdZ4oxyrfv
fFRw2z4Vwe8j4Zo90ZOORIO5yQnl4pCMAk0s8KOCJSemADPENxB+2QXtbMbH
aeTYMyrCWT79faJutJZ/U6hopCdsf527xzYoTVx/kn6e/qmB4sFLQb3Q+U3X
wt6KkQdSKWmtq8xDBXdQu3UlwbNzwJpw1SbKeNzytfqYm26JhWNuJN2DHoCb
V3qf7vikgFNXZuag9B8DLvM2hXk4S7d4w/r/Gh69zEluWLP8BxEol7WTLcvJ
sAOKUnLhhVCV2EOISbv8txjnvoeBgfQWUD5l4T0a+r7bvQOrIsxDYy2DPtlJ
CX2XdaFpcz2cgdUg/J/9hIfCdkz4PH5kmWKT8JOUig10a99+FB5SUvn5Wneg
ou+uqumiSZF61BbbS8YEE2btudZBjuWxIXV1mOcuDei2Re4ru+3SYvzEnxx1
xxn0/k/D9BJyg7ILi1piFZWHDzbL7wU05K58ffSGvoLEiRCbdGhc5uOFf07h
oqKNn1M1MP6axkKXmh0GhzCtCkpxCEtqte88kNkhbYw6mIt8V1dztjXMY1vY
W6RJDyNV9oM5KBAtMudfHddXT8FsDhHuwYd4l/76erWJV5aPigjbdSSb/ESn
FYLWRW4VzQb2Y4SWBqWQBLV5/wd4hUcnS/SxAnVOdnlERoHLDZWOvoaAeYX/
aYkfwzhlkw7KBnO0w1ciCHrOnDFWhEB9JkpaQzxL/N1SyyUj9Bj9q+QBqVyX
CTyr3wgXjGY3x8WVrkVJVFPlJWM/tQlSM5MoVqrqOX6WIVK+i7j+yk8VxR2f
nYUnmwUe1Q8pWT38Q9egJD6qQ66O5Bz3qANaOGk76zDFOuYfmMF3ZHiisvyA
q6ldPVetYXDR/NQuh2JtJ2CB4HrMbTIe4JgojwsIdRG5vS4dMe+BCIrVF8oZ
/4d53ErKC2ioWoJLqBwuNg3eHeY+xgvZTfh/3aRXhK343cp3Z+jhgMw8iSFh
Ts78zP0ns4D/DmHgJSEclTFiQxEdCBK2aXHgrw8YPNJ3YGiXXHVRKUexaR4Y
XOLCDqU6gwfeNH1lv/UMBmJetzZKyb+RW7T1ABflBGPGpa7bI9Q6wreut37c
Q+8OBK+8AEkQsWD3Q7OCkaXpf9C9uBBp81ti7S+/shTFuKfShhIiLh2w51Z0
2R1as3pJfTivkxqIHRG67iw1cfYYlU8VOyJkhIkykyiKxtPT//xyjDijEioO
bmXnGI4jUz6cOe2DzLJqNiS/59UkCp97nm+6/u+XZwCd6UxPOJkJY1xnc4Hx
gAV7JXL0LSiq2vD+l057Tpy9BR39pLSGJlbTH04ArnOezJ1RkIEEQw0k8jQa
dogJJNFbCu5KPmrGdUTY/n0TFyJKtJKYsMG1NLtate59yDPOhZLno62CMWYQ
6PvXA+VBOlqAg4qAQOA7e9l5KUoG3tnrXuUX6gIw3Y4dqzKPgV4nOd/q8Rf4
mIe7haayB7A2Rjsko4W7EhsY1XHlStgb/sN6zsBN7XARb2QvYYYKBL2S4ULu
l+DGy/GnOdjdT7NXYBgkoInCbGKIKif8pNA3oLfQ6RAH9wWqmwMROS1hndy+
tOh5XADfRsy1xLMn5clxON8Q528gzHal1YRxQriWnieqNLr7F7aeQDFl7PUK
FXou2OENZHQmwZO6phdyS7wEYdQqDBOIrAke3ySUxJk5Fjj2DTzhxRQkWihc
lZEatWm3iKpXy606MdlEMfys3Q2Rpmz4TTy2Rl5SBceIdYEs4nMsqkoRLmWL
tFX8vUqViEpEXtjrUOgONHCCYDEA3dzOrE5BlYFnW+BHXVmgB6oM7J5U7Rms
FogwYA8IV/lXExoqkFh+YL4kyIs0plmYqnaj1JdOY8JafuYyVJwldbilsmGp
lOVkrWeQE4bjVyMzcqRCmaANhxhLWD/YWpL32gMfYXe2Xs3Qjixp+Ug/qcGx
P9DdVCmCjAnPdAXbc5m1TtDhvZrLNdhEjadjnaVng+8k/qbz4eeR9Iukp+IY
hV8udOWkrEt4xXIlJG2VScPHMGGRML2HLXLZnicVpJCPHtWzsPHemHfxHEtP
jzjvs3jxibt2GQNd2xvzvysLE54vYtufHnHc6tiaabqonGQ7MupCZZGBBGVE
unX2qAelt8X5XdhviumslwpcjaF0V88qSe0xARYB1o+I3+l47yOuo4jYLhU/
/CF5m7dOCz3FjbgRLyRs15m8UV1YN/L1DW8oJLAnGO9YYWDTpBDxET+7zDqm
igP6v4W64kuIb8S+HYb3IOoDgoHWKRfyW76NVXBQZEK2P/tzkPM0kdpm2fl4
pcM6EbtUYJ+P7cXG7QEqNpLChe4iPpNnMn/dQ7sI6KDzbLcdOmQjbhNxTFp6
mGzWAzqzdwu6s5tosI0GJyKAcTeJYu+S2+ihCudiZ+J87wb1IxQj4JDqPZme
tHZDY0HPkNrSLlz5gIwZhkC+TLnT6p4tiF//IJo2qa1HR7Hbd/v3Fnl+RUN2
sSWFUSATUvX6yNp/NVx0n3AuvUPgpyYdFIKnQHaBb2z4G5dIVOQ9NLe7wHHI
D8iG8N2/yhiqbRWMmE+TrZhGuWzvRTuaR48E0lxFeQAdl5eEYhnlzU//ISa9
TcdlAa8gocB50rS8uiBUTyDg81eax6pl5Dyx5AiXVnuPYb35zteVxh/H332A
vUrnvcmvdgGmpVraNoDUeT4fK1w3/0lzoX0RfeP+ndhVcMZNWit9grEovG3u
gk6rbx2GhrEHuePas5HSfRUAvLP+xs5xT8iGC0X7VwwFuiKnd4agjIoPrsTe
mJoa03AcVk/PL8TPHOyB37FENeGUmlVTFGHCfzjIZEyjtw9Kp/06mY/m5j7S
+Ame69gotA7/q86Yy7Icrdq1HERt5O/7J8RfRVe9/kTkbY8x93GkBzTLMFFh
2OaHUn34Zgl/vFSp13PShLAjzGUngQEw/ll7irbuaJEdMYvuMetd5F1WbU/i
ypbooc75dlIHBuu5k+VXKRp0PxbhBxfbjUy2skxYAql2ON6FdvPBN98ksgy6
5CuvtlUrZkZogiWpqH3W3kLH7g+LSUsyb/TSz/HWUTGnPZQdRk8GVle4j9Xr
FBv1dVKqbp2OSuq7JA+8wqB2ATl9iNNIUKpwGTEi+swJVcJQPIkI1CihCR8d
q/YBTOxJ+X1NlpLxGRw1uGnh6WkBiDsp+X1U/iNgCEKl6gFqCFQbUlWxFMvr
3W+ejt9XWXe1bMMEh8xP9YO/Iv4qvt8zUd33TU5HOAvn4jmLjib2l3//Hfql
dgYVjfT8su3R1AnGPWg9szuNOmlQ0T9XkSPRFMk8wX7cP+6UROxPLROBX7fR
WrawMWRZhusqZL0w76OtroqFL4ucb7OVTzE4K4MjYqL/NflGtuBnCBS0s4MM
3NOYjRw5h2DYt5cHELTj9zno8OEppxqeOJJuUJdKql1dRn/LftNl22QGhx2v
wsIDU90OFtCMilm/F0KxtrJTy86vioZamDJeMKnRzsKuVQAmlaC5Aw8V+6xc
HFAi9DhqRe7mFX0En7IQ6lCXHjlH7KR+caZGcIHrJ7H8G+GGPtpbqv7/v8Tr
DiF1wEaSoA1YZIKqRC1eUYtDTv7J9LOgXew9veheY902Ap/gBnKVvx3VXERo
G2wG1ZaBTG45+ny5u9yDxcDCyiwKmQRYAdzmLYVNBieaXBsTdwzounpFmX7s
PupuHoW4zQGEtj4kob2QVFr2tg3TCx459Rf9+r3zEpGfpOzfm5RYdN7GqnPK
CPatYL9wEbsb9SGStA1F5h04ycZWCG5phnJxkOkHcMmsbPDjSRKQavf5XHL2
ptfa+MZ+y49S1TVa3el2jD282c917kY4LMjaN8OD6YVHhHuXBZiecGOxlN4T
WrtODHLurpKUdq5QIig8ti+J0djPUC7IYUw3CP3XWV7lpIrCv5WT84PM09oV
KxrwG8hiKA+gYWF6672TXRidUfUUpFtExg5+WwEuMlKBB5IG5QetkqpwZeo8
jhN8RAe40JkqCFBTRLVIuBPZ9nnUYDj8VENGs1MJnOhybHPQ7V3xpkr/A0aR
kEvSan7Vsy+qLW1f5QktM202Xkp8QALwavkU8+vtewZgYILN+VirO4RD2akC
RRdyCfazpsnZUny5BPjyjlygxLFmej6t6w3NsXUiPY99qUne8Ji4APvGJgDF
IlJziiB6/T7ChZrmMf5u0xHqFkXHeN05p989QuMUqj5pIUJZJ4ieMIyp5lvD
jo0JdJoK4q0UzT3iLMy2HfbN0j5wYnS2mtC2RJdy+uMCYCuU3ae69WN3uS3Q
x4HDXqTz1TkYBeekoiTLlpdnKVJUkRqONUsYn68GC+aapafysWQFblZnsv7L
XuKsTAgMA0WNMg34uk6IdvFG5KJ7115a0cyBEiIv1b4YuA1nkNmITQVNA12W
MvGI9gksxRyTtXYNmY9b3SH+oMu+redmJPMG+Kq5gBj0t9Hc4jy0asS11oaL
2mvMB1ImQG2c43MpyfVRczE0YGR7n9eoATuQpWwaMezKXKW4OViaA32+38ug
u8c7cGbfkv/6pncPxgzs/36AV+4+tVNsw8j1EB/yv5RPE0aracmxJI214jx6
83ci4gPzSH19yP0xX+hy05HNu2W6nyZ1bX6rr4HY2fILAMD6hOLFjPq+PJGr
7LYak61wPrceAwsPQMrVadd8hYfjuABRaj+Vfp4irQm4rBysCVqm/y2DLtW/
MtdrW56cNJ5bDQ22/tawYxv16EBrSd9AFoDs57+xqDXlub69ijOzlaTWMwvR
DFRpMaEHI9SyaZJaePXctHR1V1/22YZcebYEX40gEM7zXrYFGOd2DOQDK0Cb
Rqh3DIQAZMrtFawpQhu2Sa4dmk1KAEBMQVtMMAS//5CyrKjRXawbhF3EUJa9
vRpaSctYIthxjTlFKwUH+8WgKIf8joZQHQDFuoZuW14ZdKU/sd20WhF4SvXm
gS3g1PA1UIetiAKg5vTSLOj11X25tzEZGLw+HYiId2yMTI/AaDzwZue7I0kI
N/WGGT8BlzsvWxfNyMU4/g7pOLXCv0ghZHUibcg/YhMmWtnVW+NSv/ik+M+m
OGmD+aUGEAKfNDopTORwC1UqOr/AyHJ59DF4U/zItgsucJg8DL9RDi/c+DI9
zkKteXq2uXKVf/F+auhJKmTJ0CNT46lxJWTaWLR3BHb8YrV2glznoZtG8giZ
mWlnjl6UFx/GhgT2H434SerDqqsxifvoZcBv6h/Cizw9Qs4nKarwEMSTomoV
p8LSnQpUR+xO6uPvrYapu4ZEINiQDFQ74cjm1l02kwvYJ5WUYMzUsv0Owv7f
a9ta17Ry4Vd4O752bKIgVVxKZqWedEdFj5mSA7Ayys2ifHx11vm0I/6iuig1
vQvnoWBUTdoFFJgNx06D7WwD9XdPHzMVQ9wMYqKYwtccd9rI4Qwj/b9WKh9D
6T52AIQsS29RToVfnpyChXZISfdFTXMrlVzUaDu40zMdkbeDnWYn1crDNkU3
s8ppIWSqusb3zESilM+3mc4vxN1dwLt2PY+b538bK4vCHyr/uSXDI27xDZSR
r1nrJIZ3BmvVP8hEtccF3VPB7EMTuTm22IBC3lny9rSTXTHhzkMgBnod0HQc
fs4FAaoeC7+THZJp+Zwop+fJjpjDrc0Uq/VLAUfA9a7PpdFqNJhH87Zlj81F
XVo/32InCev5ynpbADGUeqgGWYLPXlstJp7MQRF2Reyq/nmAIL7v1A5dhFET
8elOAAzKZW5ae8YiNFuQK7socQORXoxg0ZPa1+OyIiJl1SGcU3Gu0OeqjjqZ
6SfBl48H24h03PF/NN6r1uW/VZUWGmFNLnJMJNjZd+9g5UyqzaxHOO8v8uX9
sS1bg6Tt8WRs4f0s93Kt96zisv+PIPe8+qTiyFaBvuVqDOtkMHGHzK0eXS88
e4L9850bD5nR2S+nnzVOJ0/deJ7Oc9a9BRmUI3sPrPm1hk+nPbvIIjokbb/3
wuyeT4mQsCQCTy9g6loiJdUgI7zHp3MSFCXU52cdsV8Fr4YZ0gOV2yinK99T
vjCEZIOA+NP1PuLWVP0oY8hY5BdF0D9V2un3lZ11R4Ycm4t8SGp/avxlOrM7
3iZhqlBnxAFDtZrGdIrf6HUzkpQCaK5npJX2B7CRoeJxlYLt8IY3cDHVmRot
9l1plWK74ON0VsGiDKmjdVrGx+HZMMQmUb/F/3VPVJ7bYkUzDHL5MpiegaSh
aDkLyZEIUOLQktL78mMlfZ+1Q2rMFIDY0CjFuLf9JwGay+hRHM1Yhc8f90dy
m+rfADmOBjFGiLrDSfbOvK9wTtfLkXuDCZiLuF3MqUyNSutCCT40uN2f+g5Y
h/XiaG0A+ooStqvt3S6YUGBd/fdsTWqhHY0SJhfyq5iuRZPJe2oOypKEDHiA
s/MFe8GeJRTbuxqAel9MsLduzMjuMRn+WrYf6Lbd09qUZA2pjm/OZApx2qMZ
qhtnGDhbKCZg3alnmIGwA9TNDIuXBggcFv0S/IexMcjwrGvw0OutrGbkPxJJ
i5TE9UWAw4ZcMhnBSabTp8X7pjcemOTPHkqb7CF2c86jZISzc93njxUjJ0mT
K0I4r49Gx6dxK0UhVAU5sgyVgGrtp/5XBTd56QwuR7hGw7cUJBs31oHAWyVm
hH119mqAzX5s6LQG0brm0GzW+8w7pH73v3WrIgYdPVP1U1JMNpv+aZepL2U1
gYy2bBhmT3M7xDXKWo9Yhp9JZ6D6csMvaYlphBlwC0iRwJydwzWhW9a0Q369
Dax9VQ4jvA1Ljas9thxKtu1HIM2WfrgiihvBlWIb4e1xq1X0Ewk/D0kdIh4V
crbD5KPJLU2ZT18w3XSLP4Fg2VpSYcWbp5Gas6/ZBgNvJinSfgzBJGaxu4OQ
k2fMFLxgxOkdb4AWsD22I8bu5piIgMpy7ei/S1jcOMe3t5NWgkfXRLuaDDiH
0o1lYcQtxvMJmZX5ubTWGpZnsBV0U98VM9xvZg6mgW5Yt0W/cJ5KvfJm5M06
MHtCthEJ7CR+mb7GfBu6Y95RCj5jG0DYpKfa7qVvUt3OnLnYIMgPplpanCAN
Xdy/vR0pX6r6KhQZrgXnA44USH71+wWljaTQBzJwhMxwuRcFJOJQPReMBUpY
zD57QbyyiLX9rsKWyyvL+i83bAz5eG91EULebziYkkGxj2jCe5v72WOFYkPn
AbKNwRWhNneoPX6zlsJWG8JkfffTF6DriuM5zYdjfCBs0oegtOxtyFlwQOMa
aP/QZi6zBH7BPv4A/yQd8OQID0QTo0YPt6ojF6DV6xxc8xl9dGIN4OwoG36V
Jz/jB9B9EkLcg9WDE+KWZaUNJwqfXMQzOj/MwrDVpix7SraNE8760awiRRWj
E9tEkJLvda8dPHsqajP3VTy/z7fm1vAGdCf+tSqaZbwMgQ0U2DJ+TsnqC4/M
o1Qg+P1xYJZ9ejiAC9HTWrUeA0MmdbMNx1W8Lznzv0pgk+QhLL8bXxHl5/Xz
FO00C9dSDvCRcAK3JPdRR2g7uBzZEA1vy4cmCNvLmmm7tW73v7ZcTyCGUfv7
SMX4OE0IsvmGDoq3u0ny4JNL6TPPLCEN9hiB9Ep5jRIcu+wqi5iq6POxwYc4
yChJVvBkr7w++OMRsAAD7UER+q69WIuz6y8ZlZBhVtbDs0OfciddunJlpypH
EsUq8TkCcxCHnYZcn/9aYECMMVYeshuAL/eogj2JMFoT4vLn5TGPfpicWIRi
ROLiSoDkGbwGDEjnRbCtTrVbgcoF6KMEuMSYs7LYeDTp8OKYM4e/cg+WXHsC
tbTPdmAAQItjaqwGkpGDlvCtaqODta+qL/TGN7wswEpFQJwfwHgZtSoZ4Ns2
ZFXO6aCoBn1uL5q2JUUNWtosNap00z/NJMHSUfSgg0PH9mRb0v9CEphQfn6e
Q5g//t6lYIlqunNCH1bWrU6RmhYw42K15fd+4RWnSpyNH58AtBrDtjFd60il
305+WMyVE51WLcvYEJAWdKSy6qRq6RuZ1DNfzzz3+1I/lOlwwTu5EwSvu5A4
EcKveqpqbwqYpDpd71jh2JEFpRfP3sfKLCyI3dgBLT4hswm2Mrl/teJVgFpv
O7NAEEdfsdt5UPp29JoWpKPliSxx4nJxy3x0qAVktes/Zr5LjtJdeFmiP1dO
JeNsSG1m7lsbA88zKm9v/H/0+QSBdNniHwmZnUMuYvdc4RNt5Uj8fsikCJbW
5nitmNCOxUmdWfrWdLi/r4UUgBlxNRePjZLnIvGK8BBCzIMbdlwEYMkhN6Us
YFpHD8PADanrgMOFUNaI2q/CKXcu0Z24JnKsZWBn2gFsovOGS6ZqZtpOTXcT
uDT5g7hPF+9g+QrombzqARcaKyGkOhgwkkdzry+HfL98GlAenrt67eviIuwp
2+ncgoYdPxR3mXetMI+yVZlyRgo/+fKVN+wOVjV89irgF1lm/k2Bc/G/zZJK
JsfLQ7U9fujbItCl5Zl91LW/p31ZFAGloUGlUm+t8AyIldSxk/qwztPZUM/x
XjGM4LBSU44qDW1jDHcqfttbh0k5/WUeDJqGboaMSNZ3e1JXGRmjAEcqyw0C
ehsEDE/NzBc/zs+t6pOvmOkOSdH1x2mi+wNZeDNE/7Z6iy/TJX1Wvds37fyO
4fz3GLQ1KS0tq6QtjRsEp0WKJ6iLm6Pu2P/ayW/kMTWSBCzplN1af37jT1Rt
5PtGXDNEzfDqcDtT15WsACwAxfyyBcwLMZ5+lO+r7NqLDcDlYjw8cWbt2NIr
4wPQ/XXXQJz3JstCTvJ4B56vzH1O9oZEbfvRT3GlaFQ/AJ/WJyKDdDFbPySE
ZFJx84er3PuYVAyRbu7mkCSwK4Db/5MC6EYY2m2THja1vlzAJ3BoqPI7qLPT
nX+18N+UQemZK0jjrHazNAPopyJKJrOI9YIZLD88cAMJU9zaRhqw2/HtFgjb
tFVbjEV7z583uLLMOtLGsoNprTqZeRtfa8htJApsPOSS11io47QAnC54KwDB
bNqZT0p2E8xv/3BSQIcml1kKn6rjWHfFirGC/BAlag+MRjoEuTg+q+n96L/0
GVbvbRx/9/nzNO1M/EKRNE9hhFDnvS+MjjPs2ElTYWZpO376jfyjjB/ooW4c
B/8NToCo7+dCzmQQgcns8Lq4xfN3DVhhpD16QCRrASAqMSF5ASS8P+gwLoEj
7FSk3KqlknIB7l1Dhjz96FokPmMetbIRAphNFBeqmjXzJWZfID+bB/2eANQm
56EUF/Fmas98FyC7vqPRUKDZIRTcn/O5uWT0F2druXwP+i5XkiUooisSSh8d
BViqTp1NNRpUiNQmkE/DnrgK3jdS7rPeUFv2dRrM71YqAwSYO+Owvk1ibbey
w1fk3peTOFfmRyFOt7rl1peGhrHVb1/n3g1JwHiygvwguLCkILT4cORut5vm
whMplaomErpvRJ0bw0eqB+WrX/qDN/armZzAii3OoErtJlf8Y5jvBtYaMmR9
bgLhwSZ1eFs8/y2JZ/BkMHMRheu+CQE5mGyuOPADIIYZDMaRjq0eTL2iD9hy
Nerm1UXbK0RvHfakFWrnUeyGWHCGwK4gpdieJY7RQxZ6HusNKkw+af5dQ7CV
SoJgMoXLZ/fHZ+25B0xFdsB5uEGBTXm5O9PT0Z0xrcznVlWmSzSySoelMAqe
xAxtSo0g8TJXJGGbbrlwJ3xXzdbP1UDTiKUDp/64qeslvfMQTNAFIpg7XdpH
AYOvDobZSmyYQRCezeu9j+Xkh9PuZesT9qtIb0831gwRrOsU8bwbgwm/Qz8V
deU3NHvYMzbhKL3KhxwMd9R6HYJVU+r+20H/sgeGLKL/ojQnnNvg8/Z992O/
3DaFibHwwEPxnYuWER+Cu7ZXKdLu+6cSvFGJHfOaSn3BYwzIB5DYIHNaVsgk
nIeygs0NHEql/AxSsRzbW9Ea8AL6slZgNSWSqpnL9l25S43jwRehvOul2Ycu
stwqFZADBHLTuXROin1QXUBQyoupDdnSwlAvUoWBDhd0SAReLghtsfAfJFeJ
pTdRW9EDRt5sN4fEkgS6dnAa7LYynJBiFIQAwaDGl/wFLtYqWg0KtCaWuwbp
g6e55SFNU85b+qK7qTm5iT2LoAGraBj+r1UaWRqs9AnN6lprFLipCto8y9B+
gTr9IUSyB3YEoGAKnzDmJJV7ZPz/spUi7vU96f9uGHgU7OgPg6q1HhK2NsyL
I8za19T3A6vlCtZLCZ26GgZuDNy6BUOxoKqBpMk9Td/evoqMfi8JmD2rJkqY
qXJkMsofg1N7vHv3ivWfaQL08dt3p6PZ3Kgsg67P0VlyojY6qeU55gxqeRHf
rPin3WseCF3X2EDh54TSFb4KUILBNRrTTHFSg72SilnxCnw7GpSmyVlxn9uY
Maf+tUHCEq/pCTxCf2QXMBEIXMfwVg581rNhp72jRA6vAxIBH6wxi1mq0bF3
A2vKA1MTNs/JjgWCJJwqwXU3EWo0UPlNdhymJ2bdIXc/LNscdwIvxc9LrQZv
limAqMR6iKIA0oeI3BpkF5YMNRb1+FZVbOChlTtNmkXZx29hmBPXVeL+0Gum
jPiayt+HNImhziCWtrDX+Gq7G2erc2kRtSNkxSJn+qQMXQB/AXMwTmWfvTYg
z9Jmaa5LXdYeRVnoV5FTfYDqV5IUy8dei0nvzkWUoAYUIASHaz2gEOuiRLN9
fIzY8KBJxr7+46kcAy6tUMOlzZX+08ogoc9EXZWJT2/thbwNVDT/kRih3MPS
ZCyJgmclkX611hUDqdb34KykaXtSbXy8qbqSG9dPD91o2f1Qo6GtHlA7YQCj
2MlsnXzMA27oLhwFCEiD2zlclYzevndytscsP3vWPKBNgFWPek19xMHTFd1C
1lXECCsHnfPXgYIja3UD/39lLq4QoYwwHiBFLlbfPYrRHzne9cS4CWmpeiLY
UxE3/XoWOEsUiBGkY7AiPNhIp0MDbFYlLPu97ftOvLLaPC4hQeC0+5Yt2kAJ
O5v4325IORO56nK+vHNWbLtLccKpAH8QUmACmqpHM/lADnk8cwRBRyvlQ71F
+U0EG8Bh5EUotSNh21sUr2AY0iR0P5H9XVcz8thEINMqpoJVkSg2YTyNjC9m
FBC1+nXBUrmAtGbmYuy+wJkpdHma1erDFXx3LrV1mhYQA8j+WkWre7ZXVvlE
oxiJRtA7Vw/MX1yTBmEWBcYjPuqJK77OWV+xQCJZDepfd4RN4jYHBE0zpOBg
FR08V3CZWAbG27qIZT7Vly8nDg89XTX7+eEwwErWM0FvoU03iF8/3NyujB6C
1BBddKzHP6oSS68i8w0uVrrAJknZ5qaqGN6IoPXKjCSPwMjRAZXW+d+ZgEtO
yF9+qhvW0e/mdefvOvqjgtZAieHqQf/Aa4ZXmhRI5LeLtWhY/VzrOf5upd/3
6ocW2QR7VsvmHfdDKswrvAfYKhUVcjr+83/q5/3wUUZluTiYtZ+YRXvgIXBB
FvNpM6ltDEsv4L+cEoAcRTk7K92vHXH8uMSrCrzbbO12V8uwZ9jJPF7dGorT
t2xMTens01CybrNhrvZb4JdJ2jYgTMFiMVGmDhJEUlB0w5HIuwXvvaYOlR88
lIfjihR9hHdGcJQ9i0TJ+GJVTYc6hDSaJ5foQ/YBaiv7yYhDsC08d3q60e58
3MKUxnKLfXL524tYT1Nhh6R8oCuYgncldos7ekecpS+GCGhlUkRKrKpfkK+X
JDXfAO+55PbIaSl86/4fLwvUal3HCsxigo59wvRs2SJslqMe9cAuI/574yPP
4HS3el9ubyWrPda5tlMc09nyZoFhS0+/VVzBp7hggJBPUiRHAoE9S2uod47f
KcTxZ56/pmNHhNY8DTWY3iW7L9xV5CjRflsan4d1PGEvPV9EECYCIFgboxSD
1EZdzhLTf6w02BWe4muNNAVfvmpRNKBtvD916q1/ZGM5juprB6koP4HgMFy/
IQMqlTQEDm53HA8rIISPCxdLwt61hGn1DT5mkoNcwFZNxxq8lCWIQKgOY+Gr
CpdpOa3NtgyCGSXLsYq0nTNri4iifPW4MCmKHuX9t+Nxvi7rvquYS1v68PI+
2k8zODp0QoFKpe0xQEEMEROs7vZZCJwTEciNzM4bB167Sll8DKbBzkXMjxYz
0rIaBs9W5UChF49YSVcPqA6m5kpub0wZyoZWvfOs01t1CLsf1zeHMKebPP94
kVCGBWlMLO6Kn8MPlZKRBv2XclK+TUqrJ295YZ1CCqRaQlXFWWQ853h9sNM0
+MN96XrRN8omAJ78kTKjjLHkxfTjC7s8V48WOwuXh/MMVdW0s/vEJpFaRrp/
/6cnwkISUIR5eKB8T74x2whWuoZr1NqtDLGW05iOlvdT0lo2iS5RYu1aJ8n0
LAVoSGkNNXbQINo42V+9J63cqDeosmOvkrCkOyYk0Hx86ZctTo8pWwWLZEls
eW2ncJJ2seKjc5oFeh+R2sHQeKXfh/wWNuWToHvvcYCrbmXTZNHkw0XkOfwQ
sLzVnJzzQOjLve+V0jBapcTPHT8ED1sbwpV+JS04EW6b20N6zD5pqyoUx3Jz
P3/CFN7QZluCMfCU/6sHUsUSBna24mHjU1HmAAXixe8xjdfJCxgA8qeCiYap
SP4/4oPmFX7j2VygwUrQ7F6JvErbI21/REky3/6efJXZ76L4CzH3EOhsbwIe
g71PCRpVhNj8Cpq1nlA/JO7hMTLXstXK/ko/qMRGGWnJUZzZQkRHzRhExgWz
ViVvwWF31LpF69LP4Io/BZGQ7mHnmS4on2nKTxJajauQR+HCUFBM/TiNZnvt
mmmCr02gmKGRRdJsQJqARJKaz7zKkaJHvavbvntkGUPnbCeSMsUyIv90mq6T
+PVjKTZBMRlqx4CmXSJ1rEzXmvvFf/RMAyBvHJYadD4gF9FxREB6j/Emm16x
mPG7b+912Hki8QvAwjcMIKk5l9Ff8rWQZ5yTQC8cJaAyEvbLPVtsodgJ4ACx
qCRHB3V3zZOLlIkUfo7RVcfRABpZpxSpnGFTN+UBKixMptTGrJhbu+YC24Vg
r6+L94RTv/hJyaYhqX5oNjpvHntL5ayVa6Is2X7hBOGM+NgmBFbg8liYwxK1
+yJWr1RzCXjAxUXYQGUpudAvyn/rnEKit2WgHqJkzmNrhs1vVe9Ronlq5/gd
8rxw94xE6jvalm9+lHxjAKgb7LVFZF1hntGU0Yrqqxhl+JSUO1mEZJfc7w1n
3IRZcA+foGLNZnxqMBl6IaV3rcwSS10WeccMIfPT6M1diEk7KZxjD2V8skHC
v6JHGfCWppn8TFHDOTgmppz09WL4VtT7ThVX1kJHgiKBZY3lHWoQcK7Z9Qvz
9NvCA7T7J82wCQhd98WLR3fmlZtHUKZMyCFsdDSLtyMtk3gfpKlP12Ed8GkX
0zOJlLGk6moH3mV6susHLd0dQlPu9tFOOAz/8uNZyKZUiswgFxou3hQliFon
DoYyeiGlFg/QHPLbMDpVBkRl5YvxYShpPX3nZxg1CE+7+qMLju11lP1sg3oD
kZhh8yb7zD0Qr2kP/RQCk/uuqU71+4Ih87Yldrn/w3V92eCtZcmeBaKUewd0
AZc6D0lstoH3rc9OkVogxYBtnYZ4bGCep8T2L0YacSCQh4VVHZadul1HJKrj
JKeiG3TNM7uyiUJ/XXzyUjGUEjxnRTCYe2mhQqXegixjyUDIlhNkOpojPa0e
yCFeADt8tp8U30Cayqf+yJhBRNFmFstXJUSiXV+BeX2FNm3Fun4PEIf0D0sM
cYeSr96GNUT1dSRbLOIURTbytTLSUvtZjooVZ0jAP33ho2xin/ah0ivJqFRh
ifT/4mkMx+0RGndL5TBkpInkETHAyCF0OTGHlQWVcs+sMbZG0aPTSFEqLAv7
yqskKIfW5PCT1dTsaZlAW72UocgOuHhzHRAUVtpf4N6awCUegYmA334s2lnL
OYNL7EddKbdhv92TDlazI3W5HpSqN7jn2Zi4tdW8KyZWel87OodoH5rvUP7u
ZbJQqFXIpXDKqGt9B/4MwfQ/xfYR2a2q+8Am5pdZ+1fbZw9pU07BE1QhdMj/
V5t+Fj2uEMu42i2ep+MORjU6H3WqARmCeGJvZCqzq7lilo3vfKFIiop9dDSX
1IgzCqab3kUu4Z+s/lKK7Wush35zYX7z6UQsAF8QhnHbEpZhOsw+rdFiAIRj
NQlr8qnPahODKiyzO23B79lB0b0fmMi3zPppu7KQwlLZsN+u3YfUp6OqDclH
9txns0oPn+cBdtHICb8QNp1diWHDtwiVn/gR+Y1TsnALb6iPPRgKw7P4s4BN
i/2+RIGTyIdOixRRhJFhYhLbzXAr0c63ox3K5cp241iJ+TOWRoUApsdu18E0
vx583+6qijrGUSQcQTT1qL7Qb42hCVM3qZOZusJS4ND/miHG3wVQs9zynVv2
RoHzyzcnRBGRpHU+AJwYHBOkv0tU+GIJbLo+7HxHOc2SanpAp99/RF7xz7OL
E54MIfxIiF1xWj1SzMNp1pX7j8Akb9G1m31vERPKg0ziWGOBx8Dyv7U9EMf0
y7mMHnUHI/79hrAoch6gLCwZH/hF0UyfFuISySPpk5hjghmfigQc5htF67tN
gSHX5XSOFKZ5P+jNl9O6JWWo9g4pealMkKFGAYYekfv0NUr9OGbomp5svQKj
/aWJ9ze5kuc1ng0z8Rxz6hTOyZjwPfIMvuefTJ00CoYqcDcHgJO+0hjgPKwv
PW+Lifs+zLyIQ2GGO40jz7cHS7m9XcnNRXVMjuxuwUxAsMqz90jDVCiWLrbG
iW3MmM0HZOKAQmrHJxmRc3GSlK8MkeKd8RK19OPgn+pYwRoKMsnAnB3bs41r
ql4aHCrwjtxDE4sDrH2ISddVzvpwFaGiAE4otqlMibZf+OyVBLbZuTz8Lwyh
TmsvJ890Gy/D2iC8fbZ6yX41m1b4H2YO+W5At/FP6cYpFQacDYkiBKmYFdVJ
aWEdFnY1ynnB8Ato0zQJDnSNzLTFyjHYMworvnVFbpDvI3ZQRjX2Zbo+i0Xd
0p8U3t7Qv6cdZPoo6hL+9DiJMESqlNavkxROJeFiyEiFl85pGk3Tn8La5UUI
CyXmhiPk1DujkJ0HLETx6DS8paS0BNYCkUQOpv9ajg4R0itWo+PUSIMD6E43
w1H8wcIyDUGSscbd+tzIxMhbq4E+wosPjdhs5wJB3I8P/tHWBU+cb26sVH5/
/Wc8aoGDQA5Nu7f9M/MGepXgGuaEFUeOyQ8Ed7Ccs0gBr9tK31jG/HDqItDu
b8Nhg0HJC+HVhgLkvuMxLKvELyqT9nRMeGscVtEwjQbyznxjvQV9WOWX0Ord
JGIFe0PaREQns8TL9nAYFPse3KWIJc4dh16IMTMtPHpRaNfj4K9PyFI6xDmu
GEwueYFE2tRKYiBoXCj9Ro4VnqDUF6uJkEdwpAL7klg/t+6sQmS6gx3qsNdK
QQmHyqZWGcvnESBq+VXgUiEoHOjiQo1lNSwvvtoDTdd1xzksnXTzNGrjSLr0
3sLHRZvZYqrjMM9kqmbxGLC2k7CdtLhKwa2stvXQWQejUVC8jbctX2qHRnM8
M5tiX24h5Ew0BAZkRhilKsNU8KCutnXro4d1EUj6ad3YTpGzu9PSzfg9YdiB
WNcD3CaXvP8B3JkWG6t898zLge7OdCFDgCmnbcU88wrcFn3so0J/3pe+D9JP
xWjA3rVZcC9/5WviFK+xWiVGqyYPZf/gxEH9Y1Lkw9Gj+kYbP7/uXY8urm2E
Ks8AxoMZOxZOMdBs0z7c5+b6VaC0UqeT5hK6BhpyjcxN7lZEasgCDG55T8Hu
Mtls12jpD86BIsGe5VzJ6trTcY8IV4WdwNfdn/WWfVG+vIvKb7NPS4iE+MZt
6BK9vM4bUyubAztSiEZE6pT97ORgqvoHdM1QYcSr9NiDqlFXH+dlcHWGC4SL
sRcQ474xsSs3qdQH40kSxZ56hd+YpGkl3+a7nt1b3tiLs2zgKlhST6kngpng
LgKERUwM4HiIrW7GZWJ3L2YuT4pJNTQVuK0lU5aExEyNON06gcd0sFj40aiP
wtrk2OgiHofrnozeT4ZzZyOkz+t2WHWj/Xfq9mmUEj2bJFDhSvAUrIke8MKb
8sL0HfX+e7QRGe8roBjohK0Sw2bdi56MU7sKyiWNqudEpbiBcCnduTHbSqHO
jlbxEntNgncTVX4xcGNSMGZRFjjjvfbzFOKFlBRe+DWiUvJyhJ6Z1lHfqth5
9+RC3FmyQcH9t9cWsx+ShowJPPz2BW8Y5VHgF58UztVO1aQ4qpPrMKHf1aqm
JynhyadwTGFZY8i8weYJpJnoZqySiu4rJfH6R/9rDJRMT1vp6H8UmMK9W0E2
NcKdULl8Qi6Ag29Q6yQVKFuEmP38fPystqY1hUMUuP8nAGOwK129ow10Pwh7
yobTr0qrnh5uOMUKYN8GWxoRLWlPH2Z32F5v+VqbWEurSrVdTV057ysXL7GP
wuZGVfFImnm2Q6cX21Pi5x0g3cJAKd+ghlZqhNw3qQh9Kzs6hUxP5xAUktQg
0D3KdSf/w59p3GBDN1gZb+PwqiCh59Jk4BBbadfQIuzydhphvZIc+Iow4m+f
fmI3lrxqhTdVCwe/7V9xgFTZICDy3ZP8gsEX3ncU2YbO/wtq7teu6cHEom94
f/FllVhjEDHuupNP6VbvLYADEtwNvawu9xR/v4kqj9ZWP1kzUXTtcne7jyTr
SDm06ZT2wtUUIKD1ZYgNk+593CV9UvEqFK4Tro8Rj69xA0OkFYtvMEaY1gPk
TE08RErTuWWgT8V3aSHPcIjqxLjvtneza474i62Yi5ZHTRSeBtpcfZ+2jtRZ
tJRhFXEiMJ6LbrtPep70zor6uVNL2ILS5y++Mdm70MS2Qu5+rc1N/D7C5JqE
vEhL9nZwsFF2La/3Y7wkm+9a5qgHwTsasH2umQaDjeqNoRTlzlAcNL486xXk
YMaei1/C7Ye1RrVbHSqrHkfDCMVf83X4PK2l76HRulejUjB/s4AcTu0AquUl
+a4/JXWvmaKuX5Sxn8TZ5XhNwhDHd1B3ORCBQvkipu49tcL4t5tTB+faCI2b
zNiiVK1Aa5RYNA3dicTgeURRgOj0qXEvK6IQW+guGspfoCK7Vyf1QfPJ+hym
BL1Zl/6yXqCIOEnRgx8DEehw4jHsnFzrht7LVI6GZj2vwQCSdXRV/aL+uUtG
Jw65Cu/dHrUW3nKW1A5mEG05sqRLVUg4XPuPqZOCMvLtelE2JHqn3sufy8Ew
LxXMqnOdwtKMHlotpIiSHp0ftTuRs80GrZlYjx5L027+GK3Y0R+IifHSsG9j
j+w1qMP0P1goPvU21+KJOFPw/ogEAdTjtva62BOglvQW6fgklT5nR5gOiuq3
h9Q6BYb77oSxaDj27a1O5XqTuLKk+RC77+lEBpUI2FjsglQ+rpkaPLQ+n0Nj
kVGf8EhD5vtiJtk32FYdd+2iNWIqgpP/Er0PiPEMsctis9pU0foOITd6Kvmw
cGqXvwCFU1vBDMN9/V1Gy6VI+s6OB+FFa14feR9jsHiI4K+IScFaV1mR3LgF
4q/D6MOXELI20pY46pOD3E2rBYPmzwBg2It2bRTzNzk+KYPcKtVrfr3EsDxi
0lYKWDxRzpg2p/H5+7K90m/EBaX8equAWeZHsOlIxSxQhkaaEMw6GPTt8vql
pEIiKQ8tRHqo88EdA72cRrPXXXkwphq/BbUh2z4tRhyUjXEP+YhfQJPDYfTL
3sxtMOLxZmfswKlWMWAZPHUuaz+vVJA/opotiUKn4DDqtKYgFuuRXkBS+VjJ
bnRyW05PYsmy+9hwKGdU9gDkGS0NX73V9yWA3v9EJIBiYvmHgGZhZBv474vT
7FpSJBy2/Ky8/r15Z5keLvBPYKKNtny9amtPrS7WBGfkYRLmaUsGAutMAw18
7C7DB4g0u1KB6JqFcyxHnTb45qvH0zxSbxA07XtaUalUThWzzeYxLJ0HaPvA
8k0OiVd5WBTLOB7BMWvcjqKkS/z1DKZVe9x6QhcfGASfZqxsKtPGuVq91h/R
w8lZBOKBHlbyhMznBhrbfJu7CErFstlbgLjpcu2PSQ+ceSQ5LLdse/BnZznY
2H8lqnTeSBfgGpvaPwDZfNDBJPVXEZ1Z6isrIOSDRn7RQpbCTa3Lv+0tbcpk
9rL8jXmM1mU3h7BLhxcfRhenfDXMYfMYBj4SlMCEsf//TdKwkZPFfCACcx/U
MYuOwzE4wulR722/QyzbpDUOTrFl1mzYbZ++iVFc6TkU+8BNgOpjOYrOfkRB
SdjnuHSUlBcovTDFJUlk9Db72mHHh9pKKpLchrQIMW4ilPTlTCqmfNVukz/E
/J2ftPkLVfa3/PaBvKehFrN+VaibhQdOu7U6V5mSbv+G9P8wCXnwtkqO692H
kBviXAbh3M0yVWv6giGhmLHdyHh+7iOONsrrDUFT1tvP2xWBtPo2eS+u9m4M
Of+6oromG9nUmqxrE6kiyqD0BB3kRggzZuKBCaTQ29aiHgXUFg2lJH/Xx9bp
rZq3giXLTh9h0hLgWoJHECh0QbtL9vyJfqaPNmku5PKzstY33Ry5KLx9fCKT
teIpjqktKfZALuMrhG4qoU0uvb2npStePEEY/XV1NuTemiLO04a+aAQ82AtB
jlLqFo8N7qfgczlKAij4fGQimJeuT3MLtEH1wtx3ohKI4LtughNQ2WnchPw6
xxJV4Ro1Uo3fZ9keoi+W8pEzoqdS2Rv9C1uKIPouNDHNggZPVJOKG5IPwfuH
fi4thY/qnPtVhmbeVaUBpLq9S2RE5/yspxDjnjkmo77o1tgAATBuZwTENTEp
Wt7mqQwYwis8sBHN0KFddgiFi+xgGh19UlJ4xF2+2tjOotP1Nd+DNmY39e0Z
xaf6QI0irrsow1ZupX4tJQnAfuAePOzPWguV5gk3CFyYYkt7f6LFSkVWmBYO
9CvOY4L/Cj64RZNMbgth30S/tlCFFYJmcmWTrNCCMMl7nMFXQFQUYxpryx2e
4q4WMEek69k2zc6ZcJQbV1pVMRcAYk01sr8CVoa0cC684qtjgGivAZYqgNZ8
kD671Fcyq95fFYCrYyEO2quLiOqeuyqN3NehTtci2weTOj+KMI41tZS1Vdmr
rae5HdhykA6Xe9tZ09GUlUqv6cK7OcxobMpmn53RToircx9Lm7PfOPy9QJyZ
9Gbp6lVoAy8y2W5jf7RNzJHaNze0m7EU1uPOZ2X6DIKBbDLvSXvXpLAhKOCh
L3eznd7mXi0FEIubGA3jyTV9vvRePC7o7RUcFzkIuS2+Qu6fjxSkxmEg51zg
uF4EeL/7m50HTxYB+A53XQYoVlx3oe/+tMNI+dAbQxmvGwGwze3fzRp+IRgE
s3v7Pau7zXWe55EojyQuD+LemoTjPymZr8r7n6J7hR2APjEZXuFzErNwuMhP
9PtVpxq+urxOxnYgcXkx7iNjgCLW92mTLBaK5iPV/2rvxuM7jBcugrbMEZjN
OVzJE/8+s0AagU3qAwKTziTr+sxZ5cY9wVsrMT9ojDoqBayICWdMqr+vg5wK
fFDVIs1eZG1jQ594hE3etJljtjEfXFCrzes5chmQG5lYAmL4kLASGXHDTznF
Iqkfeoy90pBhUsIqB2jKsRVC7BA7Lf2B4q9D32FXoFWyxQ31+gwyM41+zeJZ
1UgnsMCFpsarXwxP9DFEH47+JOv81vzuqlNjLfgWBpKCM0vlZqxCat4tRLkQ
HiLR75cJtVNwyULZCgppNM8g0nqP6/08JvZWsBIwDM0XnQyotD53Y7DJuhfZ
FjDO4/b8GgqvbcdKFwPK2btyWH7zrPlElKUZiYDnpwHDbZV0DB288ODAyy7u
EA2bETPb00amYDs3PLqsoheeg3sfcWU00OW3YjF0qlWdJY3JrLureb0ADynt
G0IQVmc0jlSJIJaOxedR2rBKt8eEZN7S0FniPFhlr5ctO8NcfrVzo7LimIm4
fHzrE7Ayhs2DWuvOeyPawEda0gEzriECOpT3mKnMwfw/F4BzcB9m+ZDYO36J
mHzO7eXgPHJk/SHVAbjoE8pbx+kgcS2R4/9Vhz0voOHKaaChkE1mrpTt6utH
leX4Y+sHGPmWzF8BGjZrW2EZ3G5aNQlzlX9fMgyUlC2Zl2fcY0J7gaiZIJn4
SwkuKNYauLbmfr6mZVkVYtKujvfOx0oXayu+/O5Z5EUofzqIhHobwJDACiNm
wsws9vkJjMXct/aP0prc96QlQHZu3RoHEMD2qZHlRs5TMrcSd2dJv/fGkM6h
05JQ63nbpsbmg1NUkngZ3jxM5MPaRUaHHMGFxuHlGa2TbqFf/wsDgtZtK3Io
l1ODn6O2I+puLRzwEaAILwTw4o4KI9Gq2VgNbZg58TXAhMSkAkNHVu3NOPub
dTTIBZsH6MBHjlFWHwlyboR23M6jHbiq5Qk6I5eUUE9+Cv3FU0ff+iMd8hXg
Krc70g5XX1v/1iT5xdNiYXSFuyngDlzfRaynWQkMk08MMe3m3HnCoLmtzv7n
Yu4xN3uCxu5j2L3khp8MZRTKJ3iM/4FRp76IdosO3WNqH26bS0g+Ncm1JXgE
hoWA53FIyQyIx06IwQFGI/SLjPLXHM24Xe2aPN7gDs0kZpF6xXSitfd0Ny6M
ykL+0ZzMVNkhjZVa4wk5sVDMIWn6JiZT8hoeNdHe91h/M13r83rKnU1jImhB
WTSZe38CWX4Bq5cJ1Asddh7LIQQr4oP3Zx81LntNxem5++9wE/eWcz285Gei
MFl4Ymld9/+ntK+Yq6a5Y+M1jL+dQw3bGhYqs0Q9fTlRa/nM51xS7SVzzNxk
/NI4tMsXlUjlF+0KT4OgVT0VllQhbLFw+bsiDqlSsFR4KOS1z4lMsgjKOTsQ
ESHbM4bi4TyXGJLwETUDabImHIQv4A+E1lMq+4Xr+qKg5bkeUHccBGPi13lX
WtCcSRmmmQ21cViBaQOtNgyCLHqBtE9Zztjphcn6dOTXXV7kHO7ZM3Sckbzx
0kOaTpA17QYclEU8qWyUzTlkq6ZxMKQR8AtCtdFKmU2CH9xrxTHXT46M6He8
Gcs5EwCc4aAFbC7bMAaJQT+ueqU+5hTjfIsI20MHjuih+9oR7sVJhFhkWrEQ
scXTHH90oCy3E0b38Ju9BWrPLsLoPrq7at2n4b69ctaHCImCq2MwxOHpCK9e
2ZyaHg2oFNHw9WKe4smIltYNZkfJhv6E5CwoKIrkyGZXW/uohgYcQS4jJVaZ
t7wPQlVA70dbem+hmwph+AbE4e5MGbMMq0+7Jdb6QwIi9kbHQY+dVuWIRRLe
Za64pIOavK/LQ5CHWYl6NQCpWnWGtgGdrcXv86cir20TnM19Uw2MT5z73uiK
oBxMtnorRzjd7xoelcA2VfmfGxxaT81fPCmaOKAZ2ceinRSrk3DmvLeWgJnL
hCWQw8DDPKUGRNxjD9U1Gduf+HBv2aL5qQKVZqtE0T+FIBLZUQ/1SU9lOxRJ
wlAeH9BPZzRssCFwQYM1sROxFEpb8WoGiT5dHc7dzmgcrde0BtpsFklsgLae
L8MxJZeiKoXKJmQKbGUNBSpO6LjzvgBeQkTRqKgvd99N9/gaUFBNpjeFm+gC
fdmgK0IdbwekYGWfWY8QeiLAju/ZtZHKqj6jpuVCJ9SPgbvaTExSVX1Xo6IU
1Q0CiWay35ncrHjCxIQWer14FL3JbX0qtiPxFMRPPnAG6GFoWKtg/nLQLmG8
PE6KlsSo8IaYPfQsihnY8M/JriKO1xD4CNOQT8zEQNJbMSdXXajtzU/2MHto
vbb7APUz+cay5/YMSgssvhc5XUJQYxA91P376uzHUkknuGDc3497Z9avpl04
pRW8lKCftuFXG+372A9/2pkeBWW2+VxEgI2JEruR4zBslwWNHXhip8s1JNcU
acKEhmcuJKxU3eNgFqDG0T/XxwhO0ApvWYokM+Go/wseRIzCpxOfiU1gDrop
uci1TS+vcAhaldTVDtcLpMXCyQLXnGqZqSI4bNiNSdSMOjquUhjkLx5LiaAj
v3i729qYqlmeHAEKYz28pzGRZokSkWD3oixZsrTmBmmSOoEs0TyQazHeKDUK
CSD+o2g9grD7qbaOvUUbDZzaYiPQ0IPFjld+COTwDg9+80veW8yhxjGOPwsX
6BbYVQE81ThwyCm2+46X5cOPvM0Sr/qzeQBMNc02WwuGFnO+oHeeImCjIn/r
UjEJOu+3clIOalIemP9yKO+FhDa/P8oLFEZNerrWCX3JyR2AFb2IZPjGmwPo
KKGRV8nm4F26V7dVzDc8IYSE1JWvWrxtuXwe22wuDXAVcLaW7x8dU8WI7j4o
J9+UDORL6jbQuv6VwAOzkJYw+v9F2WRSJktGAM0YySV6TnxJdhDgqvJ9SYj+
ir/uJZKLEOhMbRwN6Hm5Ic7oQmH5MxYlba7EKd3ok2nnJilFw6YS3eeAn+AF
ePEBxzs7lBLuYE7nLapxnq5AQmHL7OI7nqWXpHyD1/JDKlNZVw6jnzXa6Q8N
ooqAfTxXac1FJeI6XLokIdZQXwxP9rUr5EbWfgOea2/oflKgdehqV5wXhOyN
Mhb06MZd5pNf6Itp5TqPpDrTYWiSq21pKZQFmlsMfqhOQXZ+le9yqNEri2QR
Xf7ZwBvEi/locU0tpJc1WsWQ93KW2ibi5KfMr92vaWT0+2YYc6P3WORQlv+F
YIIWwnS+1wi1v91Dd316XO5VvJ9+RrX7QyErvJ7fVRR6PVMWZSOUyj2Y1HLn
Tv3YmdmMW32albPg4uhtNUzcIKT4wziJFZCX0tQwm6TcR5byilPyB0A152iQ
6k5rxRSiSWVt75f/iuE9UC6xTBKn6jV0xU+qPEoIeX2yG3uQfcAPQz0gMrrC
VwGOch4bUN9OwRgXCd9gs5NZywN4UtBARiSOXwLKhrmathkOK4qhX3K3aI96
sPSCm4B34JA+LRacZqXgNIKlkaDws0zZ1+5naMtEB5gboC306dA7My6mTLsj
1rmuJFuWL2jifAkYWLw3adU/POX39/NWE4q4PUku/7NUudpA/VWfKd1m+gJF
8ZVj8v+eJW1EbIvmvpuAN7liciI2NHaEJx3jniqE4eZrv+6JIYpT5gvGJbIb
1Au4JFR9ITDseGbuuJ+ejC8Tv96DxrVPgMym+y4HWialpopX9FkCIIER4Fzj
++ULvT9xvxg4HUnYRpctQIWKMgMLB03w7uOZirWEYPRWDhz/vijVaf8+dXpz
2BsnrvvzzZyJeuRA62ZgGmmY5qvraDGG/Sl5UqzOgS5ODHEVrPSCXrsPFre4
v1E5P7mFegN+mICs9oct1BlO4LnDIicNUTs2vZyHBzP1bwWsbWJ8LOsCkSTc
bI+duzDosaPr4scpZC9GdCQkU3N0z3pv7AQTKdz+YHPULNC/mUYsaGxJ6ERF
YDo+HZnx492BUViMN8oTdNKnKAyQnwhBcQnK3WN6YeYKfPPRqgRbp4vH0dTP
As0TM7WCdbmuXrlq1rYz0bAdZqWcJ5UiNr+/0Cue4hby2in7YuX+FObjuicS
ztr1fiiNqAbsgBCmSYTJZnuaErmFUTsdAJRHKysOgpTgaLUfR2ZpObBNyQCB
S68ycD8DyhzaIr0RFpqrvr/UezHpw7/w5TlADa7vilkL+fskFWH2u8UPQe/A
EI1Nwk5CasCkgeeN/cLH6gRyoCmiIJ7JMzCrooL1LtPt3ZqIXfiKChF9qeI8
7nYo+vwA8ov4yNqsgV5Om3blkCOI9JeUbC1OEgHFWOErFyFeo0/FUxrWXOU/
+Q1wwU7x4MyRPmaOQvDlRLEVb4ZvaGceavklJ9dp3NMWgLAto63z8fR7lf5N
b4JOEbDjF83CG7Qfp3rrDXz1pJ6yq705XKUpuFcS901fa4tZd65LkTh6U4co
xMaF1wx0uyJSLEojy1aOm2clFYKEu4noV4MDcXWZrPsIYFVtKC5mSOfCh+i7
0AaLt9iCDFiyjj2maUM1U589kX/YVQsZA9BMcUpnDFG2orNMTs8DaaSc4Jb0
CQirms7wSZJ8AkC9KHF2bowYqGkrM+0XB/4weFTwmv6colX/3OgjJarS+FPA
uifpPEJL4tKtfxMa3nnt4Y5Qsme3IuhafUWV7wCMwMk35YKShkHppoTRfEow
pXZ+j8VljTWoiVLm983UT8cX8V9fBDTKTAE2XkhVuMhePX2Mnbp2YFm791m5
25/rLRzQpiCGil9EfpXPWIzDWrSK3FGGJMtDUyq2yJdmuLv8rkH0WEoA1VFX
RCOAKfODoxa+bGbSY9AdiPgN9NtLndBKnulqZEHGk3Mw2gFrTVz6/8hyFsZr
Fu4XGVzJIfQmZJVweWRA6vECieaUyayRvmMFA/p7RR6k1FpEYpWadDCu9385
zaGYsasx9kQg5m6FT31ZyTbwh6Fir4v20gzHRx+aJIQ7F63z1xhYNo+gWVPa
iXCtQ4IaXKXVCPaiEpOf/zL5gi9vQenlDEzhGdWkBKNHCj1VqszGbWNnkw+f
3JcQyE52bViMdkmbKsma5RVg/t/frChEDZ7/EltXldXyRR/oIPgDn/gnd22G
MIohjwGnAdGbi9Kf9LrgUv1SoGjBZnZo1h0SuEBejjfKRR/pv3M68+VyL+KU
Mnxn2l4GSAnuHrR23lz5Kqlm19qWZyY7R1J4ULBxOjPksjJqas55BRBmM36R
Hl1nUpuG8RKSKM8xS5Am7+JrBUAqXj+yDSVDL4n4D6P1T1DH4ANVFHhKzjW7
fyHV5E0n1ZE4XJxKQh2EgyCB1ptfN0OQTlYpIVtW7M6ZJvoEdDlPmMGTHvJL
SlEvJoku4x+dvzUhz1//JylZ7LOUjs0Jubr4F0hm9g5cP/zSSmJWOWURWy5c
ZcAoYEjN/jOMezkm/iJY2b58B3rN2jHvpPfN94BBASSFlbUVeFUNhD6T6g6l
eFiks0aCuKRN57tsvqmcodIZznuO+yt69HoXi/s2ed6i2y5E2txUjQk6U8VA
taqclZx0355AXjJpYL3B4IgM/eyqbgoibnHDC+TzEAFQqaLeqH84ebxTNv5B
gnOeRayh5YW9u/nlxW1cpoV2A0tH9KDQeuuSBC6H8UerpmS2q5rIel/wcL6q
75/JnJdcT/tJF++ukI2cp7vQ1wFUF3F8eMuYcg0YmHu5uRNXqaXNtWg3uLm+
sea0fFFyKKUCE/xgSoqNOCFoVCm/LNoWSSmTz6UNe4C2TZ+frfoG+UnPxQZQ
j6x2TIpQe7BV9dcc78BglyuEWpg3KvoTRMFY5hcDZKt8QbA4kprh3dh+qeGI
psi+t2Vnzhz4HFU84fsxkBFz2xF4zhaHSq1m4iAgM81h96yn/8M3+twK8avq
rwbb1IO+rnfnZHfx8SS1IMOiP7cTeJC2zzRrVgG5xANXqOD3os2pIQ0pDaOe
+JJL92rq0b6+t9x7StinLjp4K/0BJBCd9CLh2TOPSmRf4XVsoyMHmvRWdxMs
tt9M0Xne2o0Fo7flklkEm96FrM4FFFf6zZXf5gsUxTEasgU24d++kQXCNiKA
/iwUq3qHdKJugp0rEDzJwpIBfzLtRpDc9TlGJg4ami+jFoT3pvvUdPCb8HqP
TTmm8178lt1i1o1LbjCZvet5WDfDIbTMV3Vzb9702hobzkFo2vqOQ7S3XyW/
yPeUJESIWAvkpTNOd54cFS62ogp75CSoka/K6OA3qITuCKsZk4M/JeFcN4LL
Tw3oUCbn42hWG6SzG1hRjUPh5ENyq3D/7NxgGs23Z71uif3URL2KUjNBwBDU
y7mSm7OaO9WoWauk52qniJqc+QpL1FxOxKQgg+Gw1ljJMDoRA62fMl2/UkKQ
sbbrqPRE2iFPxuA3nj2MV9MIlsPy/O2uYMaSV4lV8noRxRijexQT9qwuu8F9
6/HfBB+3qqR8GOCrDLzmwDaRLaWow8gYmPFJ3BW/zgvaPg82HwfBnzVLIy8a
8SCD2+2nmoY2hf5hoFLkiEZuf9gAxF6/TXptM7o9UBAYGgb44wQ38rp8vg2D
STQmbWG/oI52g3b2IoKyEtisA9yerYA7b+HOF47ztzxkUr5C6+XEKnw35pW9
XU28V/r+5WfAdEH0hXlZulKBFuPUBJ+a3YIY8iEUv3yXqdnplGBHuO3Ghohv
yWhu7S8jJoALRT6A4bjeaSl8KCw19kFlSowN/2TXzKG2aKzVlCylFwvhlMQS
OhcOSHIR3JhrQDZxU8Gk28r4eozzRyK9Ro6JR0dI3WjGg51e7yYK+DH1Ok/z
wHM5qODv/rIsSHP3rlSFLy6rRjEmzi4h79W1FamY5xp4TK/q4aZBULqCqENZ
qWI7ocpc7uhnLp9X4KoFVknplquZj8PrRc9bXS1jPAQcrmiRBCQjKLa5eunt
nW6ca0Hrf4IJrCV2mvIw3XPgRHkvayg3yQ5PX5JjwXFH7GBULNxCsGKcnv4P
DyUMfTm5wAsCPEi2MChrGBk1Wco7dwl0ZKgxdNAhEHvBD1O2MXUFDEUe8Hsw
CbNBtNsQjSZNm/OBz0W2V9oxjWjOFQf4pFspw/1VGAumng0D6xBE5zZeO360
8KHqOTWO6EI29qqZXTt2hwZU5W9yoZfRo2aAuYkLTBXb3B8XnGN4W/A+qtrh
pU/PiT7Tvy1d+h78hJPaOJPNhySQbgeKn0YBL5kKWgOcXBVd70i7dTAC8GKW
5x9ys2vzAOK2yAwMDsj7mZgf+yb1bnG2gTtvwp+TaZouHA5yZUA05qMdLwlI
gV1Kdqj8+mpMOQkH0bH0vkWS7PTqyQkclVzIhWG6t18WkzUE7tVhuOSFF1Ip
d9oco0Ogc7lhtXLinNgFABi6kFFUH9sejNXOLKC9T90UaQz2EP/gWDxygEyl
ytAG3l4tjmPAPz67BNJk0nrWyhGlfYEH0tjIpJ+H2ybZ1QFnF55meh9+HkAZ
nwSk4QSzu3Og2cGBIbPCTleTFSwyT4DTLWHy3emJxKHQ35WoNkqRCUZlOBAk
HJsLLNXjPRFC3bTizVvzIlCgDCc9yAKZ5pCg9EZwBqKOUNnuBtk360gWXlMP
kRqS83erdLrnUsd/xprrQHIEQY8KWWljtFzCxjwiBwJG2qH2DYnVd8PHosL2
bwsPhywBJbEq27nXf194reDEzUiR3g0tYZ4XUv80xYnjMie2W9i8tJ3sMqmP
HBy0Jvq5QCejuHIEP+SJHdNkWv/3WXQNjwGKfXLKV7QW9GuY2f82NQNtrbil
BooSPlQq00SEy6596Njx4ky+FgCO3cI2XoioXMAGdw6gYJgpycit4zwcNw5P
LPDtlYDNPGlUoon5rWcKns5yDLxMYpK7rNaBRqDpIXYtbVhsmRu18aD/1jDP
gPtLX28Vw6OzUXqMmEPUGfkhb1Kr0FCOl4CycNx8V8aL5xdjoFBxtzAzl/6m
fiW3b62l9X23kz65XT3SpG/7jt2Q2CY6HH8ysI514lenP6d7cirhZSQ2MDVO
7C0QqHaR2v18SJ3SWrX94AGchVhzYnURVslE+rwTWCGYIGYtB1YoZH7sb4Gb
MJxaRl1e8SrI/UvTg6Ba7sew5CCWtA5CyhEPvisj0EqA5fn3TZ1Cjhnu2IX7
aSCadsvqaY1rjKIa07LxQIV0j6tAEyzRRkTwv9Y4BxGMBf2/vAu74SYxkDgu
myKdlfli1bL25yyCjIPt2giIFfii8m9dsAY2YQ9wzf1eytE8DAtOydXPobHV
lzcApKRWjqjYZxEd9haI0UqetkQjfCnYKnMhWDoNeGmyDhZNRtVs6VJ/SuiD
wbFLrDrDgIsfUbvF2GB7g5rHUZ7l2rjuQk985yUAKxgT27zHk5qWisq57N/I
+MyL5wPiObci/mImgXqMIyDew0y0Xs9DXjw+SIzuiTVatSoIorqboyQVhpX/
tB1t+7ZSjY/V9Gshx6jY3K8RPlfKt4KXewxguA/561jEKHSAIxiOTr0pcbl/
iLVSCyDvMPWsCLR0g9n/a7p5O36nIdZojv05dZcYNuPivdCgBYQdsO+gvU44
qRdlo4vhSXxS/o7HbGTDAVK1RhqwqxhSz8F8S6ty9FCl3GKO5zou2hi7mXwV
CIxAfcsk977Xg4WhJYjF8RsP8fUi4eRPc3QGCDiE7abEBAzy2wyWtLyF4Kde
FgECKpJPMj2LQIvnvWeAqVBuJKXeKazeTJyjllNKh2wLSObzeeV01hneWM38
MQ15tCafTQTzGheJVgaq/dp2gWGkQl1GV09wPPGnDMJv8Xn0c+Vdwt55Y/Pw
6MNE6XzwzHib5SzCHnwWExc0Of4k3AkbsOiNh5ffyO1Y2PYcGrT03/xiYmXx
L5ORt+xEk0Sz6RATiQDKn5w/CEgcqBjt8Mcx2cElQQYVPjyY+jK3GUI9QefF
Ep75QCWhKEzi7s/TOVJdbSsZ5224A2AoYmo0tit1jzmAmP5pnIp4axahal3R
5rdi1NtQeWzmLD571N+3BkeFvqJqdBl8HBLV+hae6CJtr8c+hG6pFjM9ovK0
31eVZOx7gGtQ2W4x4Uxk1U6PtzI0coK6EHdvjuMR2MocxttxmHDoRHDBYNfk
oDYW9hkY2bw354YRL+j8jp3LfBupEIBwvVz44gM9FUbNkR3NUfNWJxxAW+D6
EHPKn2ZJRL8rv2ZUMKkjgWA1TPBFF7Nt/hg64qWR93KcNwd4nn962Fo98VeP
aQnSvAmfQTUo9jf7w63Jl9Y49M35ECSLxJnDGXUWqcXNi3Z6P1JPdd2jULiq
4zxSeLLfKM7W+XpIZmWhc95q6ycvUkrOffgM91gRJRViYX5TWfXZTovqO5/8
R2PQ7aMNy3pjLP9LaeJ2Go3NQcwQwu8p9MHmrmHWrCNn/MRiFKp5X0E7BEWt
xpx9jFfrjR7OaYj1yvVF1Pq3tYKC4+ldX8B074Yn003NppGMrCkG4uRvfsuB
6dU86yfnrTuDyCzZ0BZ5+JmiS5GDY+H2LX4AeWxqs2IKNOTdx7Tx807xq61s
kKHtcqGszu/8gklpU1XraLM9dqSQvaaGAGkbYb4l3iAmk151L55/yaHJXFfm
C8HyP3XobwgDNeIRMtJvMO5mh+7MWh+DyvZy3/Jcb+oM86wUxAgvRQ24qG6z
26bCtBnG5F+/U/Bg50Wo32cGruTZFyohFiukc3WyQduRat4Xu/OhIErQltxb
AD4UTpjYq4g+HVFrnMlxlFSXOEhV6PTsEePl2GC3uIdByqnlEEDg0G8vO0nl
3rnVDfYXsvBep9oweRBbvsVwocRIEoH7A6CXvgQTd3CZDeHP+aR31DPp4hPt
EcQvIKjW1KIEfPyzk+ljQj+2EMjn1HtyXPYCakw69o20OLv/fsYRZ1o8rYeO
kQzwEnehBCidMppJ7MQqh4fxBST6hfl8IIrHg9z031aAsuzdTBS4/GfYzDf4
e5Y3HnXBsumo9+5cD0sUGEXwpG3w6M+W3lTOcyIV0n2KQ7Oyo2xBHxfTvHAx
isAHcCRX4vhHcwUpeUk1Qb+++ftjmysGhRG1NvuwMkWqJvjJP6DAcRHsk1qi
OPvpZ7njXggDGH04kVOFHDNqvH3I91m+BW8EmbB7eZD+PLIDxJhw8+x4615L
jbH2+FaiN7/zq6D8veVr6o0aj4KJE36vVViNgyxA5phpYqJG63HPcpH56YKY
PGyU4/8Sk0FQnMXRyOjenDBEUpIPh4lWKxa56UVWyiNsaKB6ygClYga1FUXM
RjsBTl5xkjFOkbfQ5sLtFmS5EgyLXJvf8uQG78YeAdx80Pu8iaiTzuQA0bSp
kBdOHxxbjsMx2LIEiu/n7dDkk5AuzpYuB8BrBccwIll0CwM5lNj4d63drRX0
eyp6LhU1SzNdwi09E2/kxN0av1Q90u5HkvWUcnFO5cuHcDP4SOzx1rY1BkKM
pSHmcXwdY8rzLRElAoUFmypdqpDaQSF1zDcbIKFOhLYcQ5ED7e+jzgWtS1Pw
1B5s0qmgcye8bI5mxWmjK2AzWRcnOBXNWjGBuaYCPsH9a+3QhI7gOhznO+n1
LbbDuf8Z3aeuBHhviBTwavGptLbPBWEtzfjybauzvKEafkBDQLiZ4naai6m2
2VpYPy/pxlitQuFZaYpjJrqERl2eI8t3l179dC7mblmjCXTz+QBHkokUpam3
J1VB/nWKWLwXPYjau0noolkNirTdjW9ti2+b5X3CsRhaC00wbcWZPXvX0Fxu
wTYShPalzRtHa3kOSOGR+9MXCIrnKzmSB+mw9KQR9ufzsRDvLja8LyHmkLri
arJrD9BI+v1xAHrVHBuQo771mDT/haPwu0dAgyI2CiDmj6BXxwLKZwB96AcA
9ge18/RTinLTiIuRMw/xOqs8u389YhCu+tq+U89NbMm+di+WTZzHjQdHjXq+
kU9pPPVbKwaazLvWg/Urywe7XEXo2Z8avk4amKdK1S2IQ+rXwzBkoA8618sA
sl0eOePL93WtENqJoSTT093X+fowf48zbBLBtm/x6mNbsRdanuCZnZ1G2KDO
v8PV3qfglG4ItP52+Rj1QQAVcm4REm6h5SVd8YP40hZ6mx/wtD8klxjMYFFG
jnlOgk6b8NPMsbSSffxzhli0zkj+cZnTtxlHJqZQ2QN0eQr2kbLRL/+L3LVo
kYfbk/lZi11iY4y/AyTAYMJaoWSyu02+Dz4isWrBEUGEOIhTIJlvvWGKDo0q
ugsgPcbOABFa5JUC2n0/21TCcuZxwHAaRr+uRo6pgoXUAoAx8jGvHz+v5sgj
Gf/sKaxYSCjf7DGuqZONQYYwo/QG5G4JrrdgyOL4g5Sbqp8TldPDae+dhHJV
sdYqiBic8Xg6BEFEIYOt3nFF8jw6w3aiYsLiI2VbXAjD/8uB7+8iTAWF4Ylc
WSZnx1BuQZ28WfgyGiu4uB2aGsvZjeoI7OBn95E+N6mZXfy6z4fGtq/zwtBq
gAY6nPDvzfZaZ9cQh1p9P0WAz6/vxtFylO+okyYE2dTWh3pjghO1m39aqqvI
I2rD/OFSRNIEtKmZT/V7bbxnCzGUZSMafPLznxSR4KIy4T7r9IU+KdHB9BEP
j9K3aMiG36Ch8fW2+d8fWn50j6wGOFjGrpm7mJrDzfBq86XVhZOXlAzvcbKx
MCKoY9K7dv7YUAQHUrHXUPr8D/LdHlxByAMQDrMnxgDVvqOtuSsu4Vx9rg1l
L901BgyZn6v8WnuBfLnTUWzGvL29E2/T1XOAkIsv3eWUagRFu+GoXFu5uQIm
S3QrVytYrO5SfLzD+VlxkWhjGQNfunik4uL6m8l3Zfcs2x6zI/hEZkVhLHQv
XEYFnhaXiVg5pMDhShiFhLmnpf64VgnhbD8OQrLxoxyw6DwWWPGUkGyb1SiU
f7Qx4eOZLJA+XcXoERmiDLcRa2GfA08k7RnZWxQvejQRGOkDPH2sKb7Rh+qI
tE5kjV+P1eINVKIz7hh4OiYGVZfzY2OFgfEbLaaDJtFRle5udwaCLgKOkHaD
yXFvIB4D8YmdvJTeQ+1Sp6RFcqLF5fuVBhQVLWiBYQKcBLP6gIUZ+FKDHTk4
Y6Wpo72YnuaWnAcKhCx+qBFOBTm4Ji+tTG/rG5EjFMuOK/jQXG0h75RO/Ze+
25oaWxDIsFbI+1iqytot5IJYiiE+RMfOFJjUrqPWbk39rVRynC7BCd4qjBqc
tVqZtAk/A6Qobx5cA5GtoKydZPctJzASFdSwczzlbk+aGqkyOsRUnYiczaBX
tGtD2IrQI/rAFjQKpvmrReA8pbM7AQdBiQdKqWgxORzoThvhR9aZ7zdXTutX
WPG0doS8x/hqxlNCjz88zRQjQWoXQm0T/AR0fm3oPnKF8EpU9bHitkucGapS
EzFhHcy/hvA9CIrJ1IMsBrbr51XQ3peowAdQ1e1nngCAJ6D7CcYHfcbgYdUO
P7Wh6IiqBDA8L1Qg3HFygqbhoX5n+bJgiYvTC/JOq2cWfFPudRKep7R+FvqJ
+J/Q9tlVAMA/pA8xsRgmqUF/xeg03/AB0kK2ZGIF4muJ3WMLV2axrah24qv7
mR/gtMjCjT0pibQV0IzMYUAcOvVKY4Ch/YmwEOULqYV/PfDisTZXYriDgQP3
hK33xWv8SSb05i7Eujjf76bITFg1ILcenrifePOUwdL8ohesUxOzyozavEjr
sTXhD926wUESZrW6MXlXnEfKOOoZNFP6dmg2gqLEnSn23rDDRaJK4DpI//u3
95m01bYPVtVBsVqUR2uWpMf5XLGSS2Y+h1JHLTYT8DD6opZer20ukVQlfgOo
u39mzXzCfKheCs95KhixGhWzgsQthl+HkUclGY3JcFbC7rWq/+cSIsIw/+6A
GzBMj+E3+KI4cL+wmE4AyHdPvs7phP9oXNuXNQ6AiyIoxR2m3NxtQib2ezcY
NwyrRqArb0q16Ur+8kXQhPg8hU0O0RpAJjV4iF0GApovpCqvaIi03UGm85U8
NEyILiqltixv/ba7IhRonh72C+pusAi+gS80jJRFlWJhf9yAcmsNkQda1OC9
CBoPrRBHMD6CtPlEU7OMql9I0aueDFj+nVqnvtJeo8VLr5iaHw1SntI/7/6u
xOG7RdxA8lO5sHlluKWPTGQEDr8d3bBChdWU57gPQEuqICe/ab6bQNw1a8Jn
gxQeugDfmFjfP56ZqunXXrF0OVJAFKreyZZMhaVy8rxc7na1BsjQsf/meW8v
nl+t5nXVg/0EHiJ1giiTgPeGyLXcp5XLRMNcHOqy5qZ1/oKHsb3q3EewkU2F
FOL0seQiI/NsIprkgbU/Ahgg9Oci51sqqvbNwn9DjWPU/FZV+sdZd3a1+7IR
Tv6P/nrZMtjM1lvfjkqbr9akXeCiTOcTOfOQETQn8nZwGSTzCo8VjSsIaKhc
bwjrkieX8B3zEyG2/MblGeKemlg8EuTktmONnHNKJEdYeTXzME42ZRr3Tdbo
Y/zLAKt5hKzIwCP6VKJc4ThrNOxdCWVSeBtnYxZU+vj7WogVCymIYpiugNRg
oSfaTbKQOG12YogQnlabzrSgtD30BBmoVt+GoJyM4PoaWjyiw7X6GPDfR1r7
S+v6dr/ZGrF9YJOUhtU+vg13F+rqfWDfXtPoCkTas1BDFqA9/GiAGMrQw/5X
vqfRawKKe/fAVqqH9pGHZs4ukMLDBpDNC5pJJkV5kKbsZDSECSBi9rXWZOvQ
oq4otunGOyFuxYN7Yp7zgAOX0bB1pEstG2yzGJCXPFzR9Dv9dzXF+3z0URCd
zeYYOchqCEi2wHq1w8AxuymcBYNH7EASuUsf8GLbTLE3VfdK6+20obd+1zXk
nP+VkDXDP2rqXRyIbEY/qu/1S6Efgq4UlZ1aGE8BmipaucknXgsQ6UtAht3A
Cwk7+Nv84n8uo1MdMU+D3e+wZwZy0zQgRT7a2sG2SWkiJb6dggIlQmZCZ/fS
mU270ncY0FcZ0P0kkkbhy8059u1Fck+kGuGmkPBmUiGm50O/EolZY2bcCxPW
mWTZ+zHhBZ51b4smllbd8iV2lteW/GlOj+FPueHivD5umK5Pvx6x5hxbcI9B
5+t8Ff3a52e3HSScG+NLN6eYnz/daCFfcfDAMLH7X/r8n5y4hG7eZCjNfuzw
vjDd3Yg1J+INIz4pe9N8Edy3kJ0A3WBcKB7daOQQXXwCKyBobU+4y5F0iYMX
C8LGLrU+7S8Aa7OWgmJwUf+cyyy2huC6naSUMoaI0GDjrJbVZb+EVHMMlNNy
Fdh0YcqInve0xz7goTxJYjtdoCjVV9y4Kc0Qg8rTb1Okzdt9qHtOaZFABtOl
5TDRaa8peTSiv/Q3xlIW9Wlgek88tvO46dwFB6UV9WI0YEtWuxjDQPNn5C5a
ZpfVjqL4hV9jHG3DGZ6e4RP7FFV6uw3ersz43RugtHrhBg41oZ/AcjEo99Yu
GwN459DsnZHB3BArgLAw3wLe+HT1ykf5jzLGL7zLWkw3MH90In+dLEpaVt/Y
yOw7aXB2Bd6LDkbJQc4HUOXQzbQGgVyfL01IoY4Vo5/T8qOcSNfzB7/mcMdr
F2l4133EVGIbRwHfJ/Jt1gdKkf+0qGQmxSVfqPeVNqlV2ZCflOXgm/uh63VQ
v3euNGqzt0Z0ps0C2MRkl/QFlWkHADclTrZn7eUm3igsmLrRzlPCsvW7rHLm
js5b8WBN+3mr5gTYbMgZdnJkDbJ85Cnmno2EuzkLGzIiW/hqQtXyG+nj25RH
QcmOAAQqdQkd7qIYkeWDL+9qSo2KbfxWuqQCsd2RvXAWY1PJjmh7iGRX3i1S
DZzya8S+ioYKiEQWmUaWydwmV2n5lgLlHhS759w2tpwCXRWYR9xsRsoTu75B
q7Uqflgx/gKtvdAUu81e13xH0Tpj5RnxSBW/5U8n7yWG22SuI4Rkix47EzGw
rZ7KO1o+INiQAWQNCUMPaeLes2+xtOV5zYdZPJe/k4d4IUbnXo5sNSzQOcCn
neSEsKEfiWmD89S9G7dlJlr+AhW1jKw02ynwt/wXB2oXhuTY20jbglXKHQWz
yZHesPk0of0jc/kOPdCQPMEcrzKtuaXESGAIOVWSq8tWfYH5jZSomkG+Xb17
UOKJr/JNDmCa3u9fRnM8CfhiLjhOK0wrNGZnQOoi9K3XOcOlpP0NXuOeDb4H
Jk04GCcBV6nTOcJR7aZYG5hIyWkzcLcVvPvGzagWAuD5OH2gRjFKYV0PiMbJ
zVIdeUr+G76CIruZXz2FaDja0Dcu+t2w+/yqmP/N+rrvT47Fqc2fgePkIvmA
c55EWFDzSZahytMXAgrxZ30QqeOOICcYzTbqAKGYf6W8GlkmhgcOTOEVdAsv
mwErCG4zfZ+sB23UN3rjb6WQHLOdZvT9a/aNuC0dZu0H9TSqH67/uyZze21E
0PV4gCmf+5G5TWhborEVYC8LZhMSPbu9VbGIQmOUcC0jfDArlJLNT0GLP1Zz
kZfMrbwYB8v0pjYjlrt+ow2Kbd1kqRx+mfrMU+VjwbG/svSYIPA1nrptflHh
lQ0d3kX5gvFdIifF8/Z6ZYbJkiISN0cM+C5E9DUbqbQGTgf/mIYWTFglXvzd
06+zoMV24DQJ8opAedwP89qSs8A8h6opP9qaHz432tpBe5M7QWXuQRm6wyDM
xEJ7XDbRCK3xnOJdQRooT4kdUUWbDAey+Rj26D+xNsMEKdyJbtJc2PKnQvR/
AeLTHDPvZpxd3iyDB4dSp4H92/i911bxReab5A6jWDx6medT08DLLXd/N1kN
bbbVYo295b5JoGzOhWu/enbdj/kj8pF/o055vkUaJJQLi4dR7ghAZ299WTy8
VTDpT3j25qlm23RhrbAgyaylSa6XteO2/l6RaoJqONIju46QNYGYG7htn5Y1
VO3HsJvyvjdUhwuoFrwSmSBlT1AFbxw4KOlKrBQtFe+a2UvS0JoqbenZvSS7
Ys7FwATJG2qy6P8PXzuZwJbz+nrskExPzzDiQKj4mz8EzVrBnmVgwu4kltAa
OoLVosPBPZlagYn2gZ4pY7UAHp/ObdFWCDJ47iFdiW6JbZkRsO1TKOGuNJBl
eoKGfUjcNLGEj0V/GDeZ6iLEta5/oYbs0cvXZTENFNcZ2UFcxZHISQW06aOe
4qcCsJwQCg8o8dRc2KtNAQargiw1NJ7SfhNVat8cS/O3cGgbavl3JBz3azni
w26fBa5JoBFoCo4s/sdtD+CuNw6+tR0Mf13dlMJ+8plLEppc+HfeQ7TC2Rlo
qnhgFE9GHoNKaTkxA1gh4RE4GWLd9wPm2VnLNSkA83wTWXJDgE63jWS4mvlY
5Cs10GPwyqvNetOi7BQuO+UrnVBDyyD3vgsyqmMsLwzS8JdG7vpVrQ6wQgGy
qM33sX6I4r8bZOqEIZEQKaN1y9j2GQNujI5//l6W6h+YqpJBn9W5bUlqsNv9
N37SOK3H5Bh4YrGJPlr4ovAqxI/LkwrgyL5RsmHs6lX8yG8Z82tVJkxLHSsb
SQ0tOETt8zm9MyIhyOkwazcHRlsxdMHWFPHt1u3xao16sKnfHBPRqFrVgUR4
ryy4rn67BvEhnE8tKY8RMAr6ciQK2dx2lwlipyI7fmUiPOOUezoairwXPtQw
LOgJZBtdEIdRIyoqtF45NwWpphRryGwl+NE2SiE3MZtCQkGODKUDyd7jnRns
yXL8Xd3oE8pKZtwADG6WkFcQO6puijKIy5WreiLXoMia2gfBVL6EFeSgVd4k
f61XbCA8E1Q7rUWEgSxaG21NjPeWl2HGNAPDEFf/CxnUS94Rd1N87jkGg+6j
RNi5vdBSkj8g4J0W8k/qbirrCtrZhdkRyn11/nCGccl6IZQSS9Qx5SJnXRwk
HAdHVZPiN/7LBR9ePcDTQFL9x6e0cEuEHlyBXSiypoNPSs1wnPndd9LVbsGK
4NfUz8ckEtBLKh3tVNUPZD17lHOBxHiomvUGJxkPSyY8LsBJSCG1PEHiJYht
S7V11P5Mprhhh34IuOar3LqcI+8KO6wGYa9/8tj+XOLfQ1X+fj4M31hteDGi
U52Eaeel+MvhoE5Chk1b0cZdGQ/y+VhMZA6T9UqX9aYG3CQ6BJ2DOMAbjnGa
PqtmfyV2TplOL5RurWrLJxVSkj4984GDD2h+aB4A+MW9nPj+sXJfasaHwbdP
4qO9ft1T/JurKwAdAwvHOgzJ0qOm8cek0D0HxNELG1esfF3GWmzjj2iua4sb
UA1Cx8kQEX9cceDL6nygeqOiYvcYEqbob8S9SsqJzlUcM2SeY42cebuw9TEb
8l0M4sPIuqEpQpCWSj4YBfWS8uoioA2fycvhir2aYt/KwDVKQo77KkJJzwBK
xJaJtJw/xP5Yis5pfH6Q751Kr9CKflUHY54pmDazaQDQng88IaQUdaHtJQbI
9JhZbTizw8A9OTnHZpc4AMzfHu02FEpMGV9AT8AwuTusb3R8kbdQ1HTLUkK9
IXaNbjXIICwLSEOVPO4H+eRISDqS0/NtKokAZWFFmpfrSwCNmxHLCZsGZrYL
O0LtKFVzYz5QMKQ6mekuDFwWOYO8oi02uAUlyh8qaZapJxnvSnyJCRAiw03j
Q4vpOG7iVN0MRfJt9//fKiVnXB2TVtVucHTiTjYiyNJyyXakrm2V26KTDPpL
+wvr6ya/QWf3tyxYycIWUikYYUlU5d1fd/KcNG06oe1HMvlQ2GszylAsELKX
EJFxNObd8UG8yf65iLCY+Wfz7kkaaBjQgD0hyrEVnglWEKo/6QJsGqJGI7S6
QJwyZmI+4Nq4Fqkt8icgFV7dJM6iJ3+z41b4LtDeXzsH0a2CqD8Lm45xS5Kv
hH1iVcgBcYyS2ZRNRaOApGQSkaKsMb8+wIWOvGbRE2WkVGqc8NNYtueCz1FY
iIw+AR0DgtwlQ3YvIsCtRwQL2vWuHx1ngZla5Qt2HOJXeMXwp9P5aFo5HF2N
lJ5uXkqLHXEo2nC6mZnxozUV2KYkEweZyE/61/KJtBxKyhceawK2qr41m6v4
VDs2xgMwIXM32nUrzNrmAwm1d4o47PJEvxk/R/KYHTOQu76Zb8LvQJ3pJ+GK
m7NBgkI5xD/vk5pRapu4MghgWj3wPP+5OvewBDpTXNScKW9lEU4HeQHAjf1r
Jg804FkQhVCha0XObhGc/DhMb9HzAiQceVL0jBOthIWxUv5qf9ip+LJx3xhb
bnjrwNlg2mvN0N3BUgFLloIb+CYztCq/ADRZ4HwcSFJeBWdxZwDRRnZ0EiqZ
fyjDIJpt9+Pl7Ga/mRTpx/R8dRSNP0ar6CL6tZcfioPm3RxLu/IxEDU2nzAq
TC+mvvfzrDdTHwHwA1yOb/oHhOYjJv8Zfpkkw9lNqMLFSZ/Y1N3SWQo1zr08
Mr6g8ueUyqfQIH6hbn8CoXzDj6uJmfnALQcjrzJBYao8EdlujjG0otqXDshR
owc3iweGgBPB6COXu1/n1pylfnN1oxlOWBmZzN344w8TV0uEhzd1VUJo1yUe
S8RrwNb0DNwbuzbOJmhLU7GKgrm4pYskVkZukgRFunAweo4sOEiEt18FfQXR
3V7Jqx2fzYKFeq72/YaGcUNq1IyFLW+znKfDhaQbJ8EenQiUgXQqNsk+W3m+
4UZObAZYijdDLZGgG4cPdtMTNCdYekTiF8T0KYDTAiLv8vbSnw5D3/O9YTNI
bgGGYT+pGEf8nbNQlu9KYYhUub8q7UrXLE4uq68RN6fbAL6mFVzF1SLVmdSE
E8EHi3LcaRSYzYNb+AAb2ek9xObcvJTP1KsJB0ex051lsnbB9SesSnvp6HA2
yU6STRxJ+Sh6U9bZz7jSbDZkyevG8wY4Oxi2o5oQ5RNalkjL0ZzbL3PZYDLG
K59WZ8GynVIoh2urWjsCSspzPwGXfu7MyzDlRGGM0A9W5Q46DGHdGjs5vuVn
t0oKxB1UnTPKEyDHzi8zgLhN980H4vVIF5LhXqWJz1o0w5YOzHhzvDkbdrMP
KDn3hubBAG7vCVBP9DomPtScqKr/uS8Jhws1TLKYeRUGgqoWhbP/G1BZ8X2u
Al2mbRlLqYi6S6SLV9l2ZXkllmvDu6PBIGetWSQG8BwaDSkvSy1/eB5BIC76
KD5d8DTOC2A98A3L20fkkOcNXHWSbbP444H+kONK8pR73nl8BVpfWl8kGDQW
yutou8X/8y7R/MJcytVUXiBlcncLg6THz5oYyS3DhPirs/2JMktEOBbzhVhy
0WtwAMju22fx7zoMnYkpNbRC818J7Q8RFu71wukUKLUnFXpFd/odymaDxNQB
I5ri9CUEQ0mMh9gwAPF6RY+EjBkyueWQzZp+asXOaIYHp6KYUfmk2VjNoiz5
wrthqiqcDQnXkZxPDE1hHheAb8pvL92mbyXfa8lzpIovSxA4xGcSccriggr2
GHLpLYSXuEFR4KYfOdDY8A8Q3cFLztsBzoV31SRwpxs9Ug9UT6re30HDHrmD
lc4YPoBOmsShixB9XQ9z4biksGvsIqGn3tYOe3WqRuJhyvL5iEzQvHItNZrL
vHNkl5kHyXVMGqT5reTqNZgH8+nEQOigLZLLvHpSkSDXJmc8PV/vE/9t1WeV
YAzXaNkY/0oLYvjger5hgJ1hBUp1kPGUfZz1O2PAjxbn6mTEJ8GNS1AhbG3I
sWj9Vn+6KV4zpnMfrEO8sjqO/lJ8seBM4rvboo418/VfAiGe3uzWZjqGEHqi
M11GVMXOgI4adu4eFURkVd+mHmuG9hgnNgUd+AsjJzNS5M1TL2aFNccQPGd8
HzJbDXEKWVQW93BGc9d3FHeL1U1hliffOrJiafluDa9mD8utyMyqbcuc8+0Q
kCoFuv+BfyDNhCp5Z0L7lT7Skat4kMgSGm1fYJzYYMspIM2C67SxZJZ+9yLj
sUFbraJUNGtIP5vzH0ZDsW00aOaTY/E1m3wifvWw6IVQdAVEn87MvrrEDjnB
lrU2veDDAqcheJYKRsiKli/H7oMKzkeqmm1UaVNNlQH7yvHcE6sN68Kg7v4o
3VNBMFm6RTIeiUToytczwh0BogKoCAF/Z8v2KXP6PQcnv5IqnDJAtAoOsn9b
ggXijTUoX7avH4ossR2uYVupmFkNtfkqOlT9THDoDtBHmNyokyby9Tagcpsk
A/WIbkBDEYppkVjK+iqH2HM4exu4bpgHbyWrdWiy4scCwKGUCo+ArczJ1Zu4
dQG3mUDtSmEc6NCNtawkSj9dYyeljKsvAusp8AHHJDM1pAoV24LC7J8MaTjK
uOdKGd7EgqjoLmhmT/IERAgV1MYgtCXMyG/9teLA1mHyWhRNzCaIvmvPpoae
uGQd2npzyvm2CdYqMyK3n6FsgJqurUO+X11t4RBN5ZqF+rSout7AOHZ+td19
Bei2nAuo3wDvHdBIySK8T6LhjEn9nNL/4a64SeIdUEevAK+oKi6t5yvw9Ewb
pCTANcVygnOaCCuPkMQvGbvJAdMvE2KL7deO21T+s9E4vnHfmH3a9Kr4uT3j
5O/nUBgylaGrsTa1VH71b9f1e3Zdab2F7jgvRHN43wNu6Wbd6GS2gpxzWCPT
sbTzy4L49apBne+ILQA7bFyKCpk+1Ts+YiRz30TcS0tL8Q+F0TOZ77m6gV/N
5/wzunVmCw2G1HXRbUYjtFU3OlzCSpywTFtiaIzkj25fFnzbhbBINkETV9xJ
vDOhc4HDjkv8rWb20FAI1M00snowcT0AguupaZlrotR4EYELCtgkfK22mF+y
QhQvee9LULV+KyhKxeP0xLYX1ekiMCogV7FZv53yDzL96BORyCKQV7B54VLd
hOoyKYw2ep0schS3SsdJ/upiW02oxtYZp+2V5sWgsHwv1zRaVv7+trGaz0/7
N5bxSx1mLFGmT+ue/oz01XAAez8AN7/GUC284nLqBwppLOZUH13sfXAhwPBG
mIYnknNkp1+U7nIImTHTr8QFPZc/KaiP9LYdHzDva0nPSfNETWoX7TGMLHoE
ZR+w7qQ9rTEbQWG9FBKrrhsf7FfvlFjf2vucWP5vtX/OgGWBJtEnN4/ZfU8f
ErXge3y1DVlBpdLxObE5g/mL9MfEabmxQS7IBM8AHbC0TJ2wE4rktnE4r1Jc
Osxal6rK0FGTy98qX7XGIjqzbaSGPnQR//yYrvL8MyBD5F1Mda9UWVWmPKvs
9er/XF+j7CGbq8lymHhalEPYsm+OBNT6gmEKFY7zVl2r8fVXk5j34F8hL2/y
pvCchf3sdVcO0hn8IQnO09sPykUvix/vZJkdbe/fWgYuxgsLUy7pp3X5wBAK
Q6XNfBiY3sOnLetvQzV2F50oEQKmxk9QwdKah8UK+ja9wvsFhEe09V4SYcNx
vwLOBitXs2MAea8xVyiR+jEQmMp0c9LNQ0e6rySF6+UFCv9kchRDyzlWQxBl
BQRSna1XVu9h3nRKzPxQMJniGOJcwIYc77Jidoo8W31oTTRFWVbT4Oc8mtpg
JX/RTzGM4odiSQl6ZqOMNEjZPNs4dH1yNlxWmbO1ah3/klO5S3TMQS2EWejr
NCJtlNSzZatcSNTMJ/PaHuQ3t3h7dp/+TSlC8TVDIQtGU3EERdMaZmtlM0lf
Nu9NrwRtiV5vsYSr1yT5iwdwV6L2S9uifRcwnzgSHj/W2PFqumw8eEYvU3cd
Is+4XWGJLbnbXFFXicKi0isU8v1mBz7j5xzQXKnu753Nr2aZesX+7bpE8Qvo
xFDe1tR3I89Fe+4NL3pbdAoETtOxectaPNmRKD/J90jzjLbAnFk+vaqDQSNo
2gFFkNDWLnm3U4WrZRBFYv98AtUV1Tl5IA9HoTFGBlw5nYZKwpr9VPWIYisr
dcnN1VEBxmF7PnBYVz2/zHLtfxnaH8mGuPuAjeSQAXWSUp5j0As1j8Wh5n4D
sc/8eBIk/Br+uIDFkNydao6AD4cS1Tfd8OKc4jP1Frsx/DDYiUp1igRasS4O
jtbNxp79SPyi8mjypZqhw7yiHua8ryhDD0I0BYh21ERc+7apyXMPdzN066Rz
uQxUZJ0wB0RWrcYRsmoq6bwS/Qu7TqYUFL9lnK6mykPlEEgxrLsJsi3nMKB9
9M7o8bkAU+bSN87DBvpWbqw4rWXBqT0v4L3YId82FwhLHaghOPtMcNCJ3URF
spI5PGiEn5EosT+GR6PWepXa48dlfXKPFTYC5fWKCFb+F2tRROgIAWNaWLyd
XiAhTjLX1ttvkD3JmAzSgjCPfJq6OvXojxvuBkkPBbiFsZ3w85OtnPq5FiML
ngXIU9WE0FL0uT28qWMTM+wUVwaRM02zUySiPft6sLAuuEks+yqx75gWRqku
oUv4ctjWszalmsEiSBZyoUCBaZBFXKQuvDj02xlqXSyb8OY4RlW3VgF+907X
xa1bp4icDUlRyQgmrD4Sx8m2DBnpGulkX8K6HbhQNnceK9lPkDxyz+jBZH54
3/IfIGhpxtIXHvyEKDnioInTea1RmRmbIfe6yNevK+wn8eqUOTQ2ZHEa5eEH
Zb1wtjXGb50hi6gXB1ghKK20MaWKn37hKOEtNO3xvEdAUvqsxzbV7fUJzJUj
BdltCF7eV6DorRCv3lbymq0ZWirav6IPeEFn3TnMNk6cYwSll4g8drBYXrpM
u+Zm6SKPfxTcLEi/FynyWp2L+TAIpNc9eQYb0xWrqCm6x8ylRJ9UUtmOXuVq
QnqSa3iLAgu1QXktccAA1XR4yFnIpUjrqg27Ru2JMEAJj3JuEQsv6GI42G0C
jIMKEvZRfV8cglWNow4Zaa+IjLVAP2urDewP0NxZ1gizb5M0eIUx29GRickL
8GHDlUx79WpI5Ckyb2L/wxgaJLlbHxaN+Brt3PiMys2LA2SuFIQr4JpCauUE
zsqdCHh5/YSTtux/T4NAO2rZ54gOtzUBqxqE0c9iJ34JvKYXiHc90s+KC0kZ
EQurL4hkp4x3zDg+c0Sjb8DwP9UHRGJ98+HbXWqOZkZasypL3BkdSesI7nY4
MIDirpObkJjeYkPjsUkZQFd40+UoqAri/xWCc6THVi8AtYIt80VjW+0q3rs6
tj4YTK1ghTJOYCzQrno1J/OGlqEta5Wd+GpYe0CXKt0EBkj0KBnQAVguDgxq
PElcSj46anOgtfV3T6BNgrJZYjU2qKz7NGH1Pa1qpDHzly+Ynl1jrtweCIpy
ATropMA/JmpQMok+Uvzjr+oy/xkwZ2ciKOkTWaP5iaveBiA8DwpJu7Kx9ET9
Ij2cMvQ46KYmCASHiBy6edFJMIpJYd9bpfgP/xsG/1RPSB5OrNaaMaN+NFDh
UMn66Elperr6vFYSl4VNW66Nrp8XbKW/2et53jkgpIeJL8a35B6jTx7UJy0+
k514li/Eu09jH32qyfEKAbd/b2oTPMNcAGIMfSULwckO4yM9z4D+88nCkMyI
IWslErcPYE99oDXhO9ydUhzwk1/WCmQg9I/Zm3qyDuJjpS0Eho6LH2QEzGjF
XBTU8BDTaK4/vJkxGDcQVAPbAQ/pIoDNfYTpplPd2nZ/z1lpWZgRsY/cHNAC
HeQhEvm6S1SE6AvVpMfLyhc6tg3AvDgHJGSWQvqj7kbFivbpMMLaJlbPGOW8
fBV+h26T7JANyqFsqTxtsomUfMzhX4Q8lSZxScCg7BeP86gtbiQ7L9dVglQV
CIUGJyqKjV1OG8pWiU7EMU+fzpSVvGiaHNrLheeLQtQ/mLaiox7w8p+P+xIz
IElkasMfzIpnUOjkS1eELD/wGpcZZ1rbDVzCb7zSPB6rSlwlwbWI/jSbcdMd
auXeTV8hfx9Psb1XGYOKKNvQLT4gkLlMKrGs8HjkC21nzJMj6WNBeh1lZsMN
XgxHLVMReALFT9SU4+/rIKcqc3ZdZmYUCMCaEJ1A5qsGwvtd9u9iscy0Hzc5
5ZW9gEzTea9cy/WfzO0cttr1nXo6FK3NWZ6sasyPIpBLYSALTpDI49vL2Vpc
pjRpOsSLXzig/f6Fhx/dQwy5Acv9+8xCqT0C0Scq/a5Jf16LhgabnrZusYIv
I/r+lr/UTAHrjeJuVchSZxeqaT6SqXI9A61oeQgAr0FvRdfWYXlgN3B32vwm
fS6SFlPRHuf9iJult1y1sq4/39MEo7wnizVu+hr3RrFtLgl193v+IKzCLc11
BRFlWwZoFL4CCv2dGokBemYy4gSOdMsUGqR8ixwNYfEb1PskMEHhbBD3ZjAk
SIL1HKmxQKhVJVDIpyjlcO0ArpTk2js5S/WJM+csheb1dbqcef80x5huUbR6
DI2MYc0kiokGqBaprdfD1CsVbi1zQt6yBVh3NND3+kt+2rj7mSgKFWjZ1XEJ
nADQm6yXAr1FFb1EZzG8Hu/M584ilLhPmNJ0ZBpjXag4jI44gjPCmWGKTy8i
TJPWd3k+OHWOsvE60z+2PcDff1rkGWK0lolV1RfWbp79Ej4clwdbL552bgTh
seRZWB/z0ao5HA7149fWa9r/iUeKAiqN/59v7Tw4XrAPz15qpp3ZmUGBiIol
/DdQaDgKciuZEcIwQxKzgDV6GEq8MEPdZ31hGiFabp6qPTXCxhsWbxG4gNoq
GnK87s0QRhcAZP4AEMzh1W35vTiBfHesbalZu2K5TyTrTsGsYFmtL7m0vZOa
K2s/NJKB1XzYj/rZHAnhjLODNj4nWSAB8SxeNEBLRgww7TU1u0h1d2AMNuhS
OvZ9kLfFqR7wHDij6MsyZEmHDhtND/vyY05uMSkqzPmN6VTlj7Lp1jkF9Ufw
OXTHwnopfGPd/5L1QqrL2JgcuELrz3jz1/wOk2hcpdCT6qhe1z8hW/inPeGG
xO1vuTWQ+wBrUkj8j7ZgwzUrd9Oi3FfMXEHcfKW3k8opb2FgXPnsIOg046si
5b73CdwMarZcXk9udmY7AJCUujPUYvYSUS2jrhtNi6r7S8tp8mDgIRl2tGGU
afXh0vqev4YfzCQqma9Wc//tq0FWWF0gH/vWhDYBWF+mR9SH8N60Tg8ud8P3
oFxYaXEHLSUEajDR4bXWt/JK3KApJSEH2EyKJUgl9Acd7vXofPumHdViuuN5
FVwg6zvuggdhfbWgOQ8foIyLmwTq2jiknFsClM8+8dIdik//Q1L1WsHjPeWh
GkfiVGHR0lUn0DTleAiXEWezA8Du2M9JdkqiktZikZypSAwAkvHw3rQU2+ev
/Qgg+6nenaTeAkpWYz9HN67lV6rSbVrLQMQX15+ne8s8qgm7SIKsi/oQFihx
i+fbjrzk+FZgfGCHh041XC4RYlwt9OK+uA95IXEbrICwTxucq7HYHX9bNQFz
DZFX6VAxPHvEwxRHYhIR8qch8DNrKUCyzaeelEX12vQ7i89HO7ni/KsDKDhH
fjTD++QqwPsWNUxZSvy3KiJjv0pg6ldGQ8VqDlcGOfOq1ctveGYZYLaLNDhI
smTAuzIUYhZteWWIPnrkHRCbLg3wTHu88SfRELASRlgZ80qk2bgllzP5bMoO
h1hX51aEz7wCQUqvVl2J/fXDhuHtNNlKFGMrUa9LP9nFQ8MdIiVejz6EBJAF
Bsu6jYhDCPScoKFWI3D3CtpvB/X/wy/ga7MweZuFlBJ6YlfJ2kJPvV7/LFDI
8MffWcbbt01IpwPjUDMvzlr+RXwvq9lWEnGBnWRna+GrBZttG5yW0Kh9WO3N
ma+Xn6gQlk44H7rr0F2e0CqJDrI1gyHTNik8w9InT7qPfXMLZ9vbRlB6YC0j
3GL32/oJcjxOQdku7BNwpJ5gmPmvAc2kXAFBnRz2qjnOR5AeCFvxi9RIoQ55
yg7/8OVFLL4lPdxt2Yci3BCvHSZX9H0aW7TsujTvATHOolj+kCSeeGftuFyY
Ma0o/X2e6kOpKCgQcJm5CbXO1A6+mOxP51aG46hbeHXNLKaMmcLI5FwhWabc
FTzG1f2Rsdzf1lQW2wmjuh2tUwkn08NRh8kBUTdDndmb/0f93vb3OhT2JGvp
sQnAO6ZXa5kEE+EPBwx+64buM+4Zm6e7Vt6aAjN2VuP22KwvxGz/VZByDvk4
xCQckBaS9VfxYewfUdwlcn/rWID4XUjN4eYE0dqXALJ+WpBNKHdJdwVzSYdX
YYPihTHshe4hZas0Sm2ZVwQ7IdrjXA4sIRge1k4JmU8zWA79mbu0++EwZmbw
ptqGOVW55PmvRi8JZjzjy5VYNRaeOs6C6F15KYq4pVVc+ZZsRAph6sHCQnAY
Nv3Ilnjb8zMuRKmpKRxsuWNIoT+CdgO6++dciCbECeMpt5GHd4YOyuHN4eXY
kDKvezCOklRKk7FyuA7QQjN2lZYHP988sonzWiO2W9Xw7xh0SXyw4bP/HUUE
24/6S9DNqHYLubC9itCPRXg4x2YV0Np99tfGVqWHILGgqRn9I2rI6j2EqdQJ
CTJim0r+JE2gzd7M4Qa+jMVVkecuTgkwSEazA6ox9BywyVi6Nu6X900ixyEA
/I/6yxHUxiUZhmYEuiYwZOgl156TkW7wEuo9Y07M/ftvMDLzcdmSKWxzk0Hr
o/8xbpjGsJ331WfMREOMt05LfbqHTwY8nglWkOnIVDBANhLDAuIlVnQgzkvS
KgeB75fcVJsXmXSwoVl4u+OUZe0NHw8wVxYXZt3dt0Jo+9Zmb63MSDDdZFzF
szr7WN+fUHLleT+jpI0dTU74l8NujPehRoDKkjjfJPBtcUJdnI7TNKO8nXOK
VSZ4UxDDmhP2veOBjNLpzvLV7w+sngggf+DrhR6/+wYCtRP2gDTVRvjH/mWz
45algYi+25XyiCzHODX67dhBx2NVGhSU2FIsijHUuTWugr6daztd3THa/Ox9
Stxv1TgrWKyRxV6hG4wJRCI13fjADwqcuiuVBzzyfgQmIwzqego8Gw7J1W5h
wz902Hy92YJIjepL0KOOOvZG2EzY9vM68PwptlPuw3kXv+7cd4oPPGCllCzW
o1nWlRTk8ZZASU2kC7fayxP3+0b528tyfkn2c/E6p3CFHrelDVTDez9MVf+T
Gwms9a+UEJLrIV74giRftGmu7EpIqw0IUEKVXU5tJFrZvLBIBeMFllsd8XEx
o/wg8/AuK/eFdmLVRLy7wbrTmgdEogiborF/lWSugcwIYGroHHw3FdQzIVzx
5tcGYvoivwVDE5DsSHXVTsbXLtAhRU2pBcQNoMA9x0XirHr2ip1RPtHHucu4
gYa8V+GzaEIjdm47R8ObxqZEDgAHqwVREPBNk4Lnu7x7ha5soBVndfwLHjU0
VCeCnCN3dvNgjXEFMF6Fu30+q1gdaA4d2Tbwlze/nA3cve6xIpWEEzAn5APb
IG1T9XmCZEh4ud5OE+zE4vZJbPq3CIIC5v8bYXyriz9XHSJiw1uZG+bAfcKZ
3OY1dlXbd8VOoe6/76KH9xvB3qQyBWy6zmVjLg0jiRmMrxI+V5V1FURJtsLb
yfG61xffD+bU8vrEz2OLwqAcCrQvmsNREqcpJzCCWVt9S0PtpPA6oRVRXbP+
mSJd3peiw+ZUCmy1u/FmVBjKifNlsb1cYgepwk4kApPtRNUxcmdkO255gZqc
XcK2eWv2CFU/OQ335HzdS+tOQp1Mqb7K6vbrnwhQwQ8ez9ssfQh/yTUr+SBG
CnVYJ9auBWG/LVcAzvHOplwVLtEm+L14nNYkzVlSKXQni4BxRh9lgSr9y/Ie
HnV4aLyp/dS1nxvi4G+DectrM80Jjafu3g8Htwe9casfGKkAEi7f8fVg2/9s
aVehyST8J3Nu3kTJMN/1ZCmb8352TxSjaHSqDXJDpQ4matx/yBppaFpFiy4s
KAi77r/hHXOMeMoYAc1cPqjWxNauHSB8f3U+FLgwW2qu/Fxemn3QdQ+o85sm
DLXoCaiZjUb+5s8ic86CBb/S+sN9w6VnUS8n/gO+xqX37BknPdujQHB3mhcE
fVsestlFDbGRg+75tgect2ffT3Ul4vjHdTEEPC41ZARMHemkc6165iWsZcYj
CTP9WIAx3nGQjqIqQUgLulxbEDZ73uPxcLV606DBXRqBj91GceFoE/ZPOHWB
IWJppH3jvBWkr3h9BJpuYpI96UtDyxxht8L3YH0Rz3IqTkPjKbGD5k9nuuBF
rYyI1iFjK0jIxx0jVo759u/lHxHsre0cehPJ9lWzNH4IWosNJn1Y27ktoeNC
bf543Q12OBE/Jc6YmqiPtspo6jNh2DnF2Mrna3J7CMvYUyJ3xGPjdjzt7mFm
RJmHe0GZiXqDTeyzA1ZgyLSd9obRWfoUXtojtNnWJlgcGtt0FPOHPiShCkKo
AXrq3+V2hvW119c/c9eVSFVWatHqaLrN4gTDs+MBPKTy5yZZDqPm8Z0eXU8R
igi9MvofE3gmiG7/rlgKwZP+PTqsjGxiACzNPPi+E5k6Gy2/tBzwO96fl6tz
ek6ycmNS3Wcyv6slhKASTAEHvtHpQkAJF17zImwKrk3m2b3jovo5RI0lC8JJ
AT0bHReBK9SzLhhjqZEEAEosgQr3ZzGKYPPojIA1UhfoTaAhMLbfYxvj6BWW
FDj+1mykUoZ9ouj5w5Nk8cXJ/6IeHsDSqwTC3LVWaYzdLugpXpzJXz+Z09oC
gjRDzbq9jJcR/RKEgOxSReNXAb1/5uDPIXXHL09D2RHOnEO/fLU+lJxCdxuP
eicMjmnfakQr1gHPwXZwStHYKtzDIIw83PflNxCJvNN8UGc53Z5FnPHT7pqG
K2ttgWqOPNH+U9G7d94PRUjsGKOH2S+GHg0t+9fjbrsBZKOnpGegy/4m1+FJ
82AebHioOnGiuQXq7dk18Z8JPLJoc0XyHUr65pYf6g0uQdraO5sXrAjX2R0n
rgaO4e19yskc8eteQ1Dj10aRsfk+oAhPUmOR2tsyI6kQaYb86eRP4yI6mJZQ
W7WoufJP6BgjJ6cVYyFJ3qEtK6HqzuCJ4lrVNWiDT089HtHrIkZKGf97Okvs
qKV8cfgWIf2Ry5fxKHKjh4DCrUaBLKQdS42m/Bs5Y7BRo/dh25bICnTflvdE
j7WkFflrKWPolxh6YoWYp4a1Pn95LNZFoXvHUhtAcJk9A8Em0XM8uPv6EIHR
HO90JIHJGVl3MfmJYtLILqOqcUqk+AjGR7oPGAvPjjsCFr0k/i2CjYWqLj5L
DgeSheH3rxfW0zRHphxJymlii+VDf1oEN3NS9ClNfE8MhpDlK1Ultgr2vGx/
ONgYjxsnSzxgrzrTsxm9Uv0hJSThnXc33XjdBQqX2CubPstZ+FSL3IQkya0C
KTqeKcKtoaV52YLs94AbRLZdXLvid4eR2gHkts7ElSl/zMipL6N0D16blrM0
OSRE0nGSAFrnxGNx4rbna8ZtUHV+zWBkExI7enXDK2nv8vherScP7ivbSV22
4298E2OwM8yHfY2ZZQw80TTpykTjmj+sOyc6+Tl5barO62w3oHEuTZGqIgE3
8HUgxMKzjWaSqFdvFchc1+i2aidkzzMruSKMAaHSTDKwVxhaTQEMDHCzjWXJ
IxMT1tbYFb72ucfj/E3X9dxTpUGKHQ4qiF1pLEpTQ1XSPrgtks+vpPbrS+qF
szmJBvcLQFv7ND2p2pUvtAclAwcFmeF50X5ZtT4jXqJG5HoAJyK9p39pLWJp
jnPTv96gScKDVtdx+1MibvM7wwFHcLfd0kry+khkVvZfYwF0cfmWRo8L22iD
1wSx48phUpd5mj6ETtvjUwTHX0Stpe0wn9e/vtDZjGJXllGP73Z+WDawfSgr
YmgCme4tIfmVoEArCqZuVzsZFB5XGwEDk+Pf7LtheO1LdErBv1Sn/AnrP+yD
5MOdSHqHi7n6EyDB6x02PBredcgRziq1WiZlMr+tERvNd6uz2y7R8Cj+OJBh
TxXKZfWQVh6gM9tyNQErifEJZncERnuktUYV1GwY9Mj/HwLaopjXwG6INhGE
EKugjSfBLM82hDuJqd63MPJI9VhvRR9eVwU1AAgCAAavpvzsBAEBfU7XzkCE
JzHdcvi6cqj0KC9r0ll19/bT/7Ur/eemmZ12NUBA08vBj/YVx+fXdatG+aEP
RQ5H4lfQQLTVVfddtQjm5tUEtoOwYw9BwzpiP45UQNyOq5FiEj8jPBCSM8ih
ZZq01XaG+Zm3s540nlfGuCa0mPg4jshkcL7wA+4QZmtk3DWIgDJH8j/CfDYn
wFzQ7TNLU+hksl3QE0j+M+koJuv5JNSfYcqNLXE1RT7hv8JQbUF0BNTAZfl7
TWvWoPEuYf0t3pMM+oY40KZDyGWSMwflodg2vlUhZomRLgY0lABP+Yygh03f
PyMtRjNVvtDcTlBupqi6iBmL6anCju5Qi+8oFku4om9mcYNycqiWB2pHqvol
DlzavEvft8XWnecmuVbi3e7CcFI+lYA/2Jix/oELff4+8gxpiJOTSPfC9JGy
iOQ79kf4jGHrKOfHssKZO9Zv8EM7kPR1lk7M14/Pm3MU5uqcFAqrH1aKoIyG
kqhiUZWVcLpaegzMvo+jrpQxqUYqIf4EflJgnPwFyfBPKgIwq0sze4BEAiw3
CQET7L8IcaPfuiqSHGaIOmzf42x3INXcLuWWXE2XjOwyGu+n883EQ8GY+6PV
MYe+HguEi17jsDNvAcxNSaVHJTe6wNkqqkEE6diugYXiGRYQ1D13oLmKdQUw
lr7Fotz0OwlcncKxc929Xfq4p5nrBiYH40jH/nb9oNipldkd6t18IXeWtrou
r54tnRQ/1AcsCMJOsjqAnH2eAWpUl0odrFm6VYkdhYl7Oc+P8Un1hzP4VY4o
rv6gXJ3rQqmtHF88EHCztqcdHEuNS/ciGHZ32Op5oNBZ+6xfWuMNrtgpar/C
x98yCLEsoRLQdlBcYfKidTsujNIftXcDvQbYX3qSYmsbE3laCVwD/ye+VOrp
Bt1JUmV2fv2TlptU6f5N1WNB0rXCLnAr+gLN1Mq72nhqrHPz2S94JUHIwb2A
6PTMkYLmQ3Chm9t8yrNr7kc0SYsUPnZSz6H7XSbcUV1ErVP0s7TixpgQPlaO
rG9GrYwTNI10UEai4j9y9NF4N5P2Ohy/Fml/x8/coZHRAGAembt+AACwbJqk
7qSg8REx0qxiGzN1e4Z9HryYqDpTQbRq1JMCM8vWaA/N89XwS1LzAR7MM+CK
oqvnq5Blnn7uLqePI2389z9O5DW7opqogDnMrX8FxrQ2zIimzeqNmH4WdeT7
kckZnQpZ9esU7jmLLRRSFyUID+YWScXxQrQcKOagg1mofvfyeK8XPLImOukI
whGQdn+jeERVY5nP9UicSbHlo0SM18lAsQokkT91OJ6OmBUIS39UudH6Pm/C
QBvRebUj8/nJd5sf3rAZIwQJKupR0vV+Em2bf1ds3Brj6omPb02VU9IDKrYE
1B4/a4q5RH+8G5odTDZTbBvAz0IXX19aSTdYHrGNqfBh70Bc9fAlTszuAWT6
9/9/R/dyvujHJBEY8dZHfAjuphf5DbuYIh6lMwBztBORboJwDbeHLcFxxdSE
sRjiLqYvwT/f5Uat7EhVrVGN0TA/nicYdsEvjR6pxfafuGaw/etd5w6gF4gM
Nn/0086K9aPkP4SR83dBa7ATtI5vlA4ji05Z8GmvEnW7M3OgKuznaWnPz5Fv
oEG6elmjolNqhGlpFkRSsYVS2Xjx6NnoQo0AcW95TBa+zLC99TYLZkU5d51x
FwErlFusiLQALyypiOWl/qIQTdN7YlyDq6EKm/ed0j3dNykOKOmZxe85lx4k
6P0HnCFtDhIAti/HPM2nMuECy48LZ1jfBtmuV74Kx68lO2I5ekYuR7KU/BHW
VFWNZ65kmJPBKh2WxlRQ+mocp4vQFqpSgIV1MAYeZloWpEly6CVseUJH+UTd
3wb7/4VTe9K+E/QLSqltgjPP3dfnBI1VhIcAW5Fe3nU225c9dFCJNlbJANQM
0U7p+FOZqQXPoKFga6AsCrWK7ihcu/GDzVx/kk7D6hvXp/P4vxywr/wwbEVP
8/MR0LfqiPw68f3U/uGckr8JxaSTMZBDw1TxCz1D2UO5deJeyqDuJJ+PXaPO
qt5yHL71Bngc/I1SuhIqu0nNRKizViunzaeVLRVtdG2Z1lQn/ICJRPjFHv5Q
F9bN5dK4Z05tovmPCUEPAQEIbzhwYZOiRJ9iR2DzXhN7+eZvOneIjfMM7bvp
c/KhS9T+0K0T6N6g595dGbtXkQfR9VspElEXgi5O8WqYmWYru7mUNQGpZsyl
WHMf1PgNM2a/crlA2n5ZQEdv+s/avTRSGWOklgmIIL/npebK3z1ES2Q0Sgma
uQHa1Q22SD4gLXT+QLs6xPtBXKkTPADsel866HVrhGPFpvr9U3xRciFgrv+m
Zk+nZfmOmolv/z3Tb/Zod5F/TaRN3zkGOQMdP6Cy2WtrMQnKQxnn51VQVFN/
wIHNh14m6vfao/Ays4BdbQYYacZ8FRMKqOSbSwIX7osTwNQFQIAbMSw3qFwa
Zc5CtFSlLdA2j+aMfid52yEEkVYicDGuHn+XksWfDN1VnBexNLVtScATirlb
xz6WjKfpgD2kBP5A/ZOXTp390cPjdDcBCUHUJzKCBmzA+0IL8NhrX10C147L
Xfv2tEIyjcrFJ0zVVfmE0aOAwhiBZcC6g0TZGPEDG3JzJN0U7SfTXsEqGPhe
/5MNGfBkViUNvkF1OOD88PvqwAvScSNWS0z241SrxDQtgBjSqridkPOL2Mxh
ppkUX3Ximss9BLpyd8RFqIJMy/oxhQb5vKlud5zqcNfoScGJsw6UhV8mLQ4f
+d0JMkRBfnwBbAS15/f9jExc2oaaFuRI1VX4JNBUsDinrBrzObFg2y6LvnP0
Ud338CbOWE8HrBwG37WSpouASlvKP+MLKVxqqMvUBGDbNDcV84xkHiDpULM2
/SFd4cB/5O0XW9pQLpsMQCNWJsysV/h1+3Ioe+BjgMe951GZQqGNNN4UkyLG
Tr6zTJakmDc3NzV7wtrxNBbdWjdyFQs7tf1nLzT5t5IvJJpRl7WiBLA722fE
txMMa7p1X1RETCWNTlZh/TlpM8vttmiH+ckO1nYi7bfFcpSNCRskbRbtLEvo
wN6UKcMSQ3Z/4nJP9GPXfhJ1pHyCOzrV/DZjh8HoObed1LfH+CcxXrArMxck
AM20P5WhbCCIKvxIjG4Kw5PVXyQxc7CXg1lxjTGQ8Us0zZ4HAK9fnxrz97PT
ATWJJ0KFtiTIHU5rlB5KMi3hFdbGLf/fVMUEkAxQIrdKgHHEaGifp8FttIeK
O83y8bcUKaxyEdoO1X6vk9LD8vEM1XeMDTdl1NFpADIgO/3LeLi2vAW+WUsC
QELjvLS6PtckQCPGEta47iOpcAVPcBxC0abCJozvx3XV7RvE682VDoM4WnbC
ok6plc9Nj5o9bHzN/rYV20oiw716hwJ7y2MWcCABwbYdQz0Rxkusa9uXCQuy
g3iNFja3Qhi3lVi7JthFcaKPQgW2/VHOhkJjWWkx9ZkUYmS0sIi9BHhZt+iF
+FrrsdkGqCzTOS8YE5daJ+0SuvvgD9NAOhdiAgS52JIsCMo9NEJ+jIqxrRIt
m0UzBBGIjx31MX7aK73vaGhbgrQ6Zn6Ef9VkOZrhNaULCpc2HPCnAgk1H8gL
IlYsTAHMJpX2A9de9SShixSbwek4HwEmBTEtWYcPOhVBT+wFYmo0QfNXYISn
whGw3R5+x25VqQpJusEm0UGpl5Ga1WtxOXV7ze0wY3i50OMWWvuTFJBb8i+K
j6q0JrTW2Dl95qyM+oD55LbCSJ3WxrgIt+heDhV1j4pi8i3VtwmZAm3cDS9G
LgQ/NO8HQPY4UfCF1tvjkm4C6SVgTWC/VCT3viKE7LCqQn5sUI+drbqMtZg6
Fqg5tLEnnKEGcot4uoBy1g7r08h29plWVFMcv5eDQG+xn9ftzrLSpeVTWduP
4XCY7FX0qYOXDDE3vmiJfvTGvVOaffRN8rk8QuM9yiuZQCORlR3Gvp40FAoA
8Gnh1Jqku59Y0QP1SwUEcTwEh5ZrnmHaLVlL77Xr2fiEFXqLbppJURIQz6ra
t8u/dsjrsvymxueIL/SHMSmUZOiBolZ+j+v6+64efSZo22IBlGblO0WpwDfU
MtV8MYT7AbyuTz1SnMxYhF0rEtzB0M3Rt8wY1PU0PeI7hNjbEyhb0uDqfPyf
MlAJjjoFBTkZh6vmKpIPPOgPc5i+HuZB+kahJVRrXAKVdlxLS9sDjg6fNM0m
gXu4RAB16ncWkQl1b3vNyUNdbGJf4Pa+nDTlmHKzQmt994Zw986DJ2m1UjiU
xQI3XBZBYpuZi0y/ZAp20poOCl8O/vxePjfZxiNvMkYArhGHY6mlaKy9Gyw7
XrxYDVnBRnHqAIKUHNC9V8cu39TsqI9slEhuCCTdGaUs1XQ9Sa589hjGuaSJ
gVHiv9br/AaeVR1h8HgnzvNHy9Ka4y5YDtbVRqyZhLCs895xKJuYjTPqUADd
LvwvZ5Zvc5o32lMPO5Jxg/BvxcGPXzoP8u7i4vSL5q66ctgzCze3UBMhFwps
l4zGWRnH1MXDB2mYID0L+2khxPH994QyyToWP+ZcJQRPYDcUrUZRDOWkVbp6
MmKQUojcmPbCdvGqF58MqOJjskWU4xv3wSZ2RhR2aNiu/su/7UEY21YlCx8D
tp5osNJe+uJl50jMBinlhEVsn496LNtefKuuDWcKsn6O7ki+vQXbuOMse8GC
Q0sbEZ5Eo8XaKCKRXcTyghlYEluQBWgRpc7qKD7fZccAYErCkwJzfF7Oj1sh
bj5Lt/Pz/RkDsPXRmjLiZZyuzWh4OWY/XuX7nytIqDk5fDBCYfw32SHF9bLo
gd2HCrQ+YG1TGtK5Gew+N3YGe3Ytowbkpn9/U4CSZDhzzW6CaL7fBlRr+Jof
okdEldeBQdYlbctfwR7Zq/d0by6NxN0tVmqjlMKoo/TlVI2bZj6Bj/+K1Q3a
/YYCSf/d5JDHFgFS93Iy2KFyHsFjtq7c6L1BvHGTIgok/eDN32LpOUXsEhab
2/DrWUPcDj6/TAtilJLqmzmUSqsV7FLhgbLC0EfiEYzmKVRebDXWOV+UIX8x
UxeR6CLpzkFGZFdXyH6hkmg1YEnRO5KAsJaZ6gJAewRupuQqwVLD4L+YFUm8
UIMwnEI9cg2KGoZ0qhOfKFGRUqq+6ZsM3vNlc+IibRSfXyjYHOwRu97H1vlP
VMYQbReY3R7Fdh1chCoM++bR8V3s3toTiq1svQERoCh2Tm72QppYdlIW96sR
d60hl3wAwphrhr9SI3V8W3m5crYjcH5TWak6uEpW8Jmhm+FQyRBfHEgfA6CN
Q1aFwng/9xHrDR+a2YIus1BC3Dk/OzJ2zNxWZ46+lpGlhF5hMrPrO0iZvyW6
9qpDKgmEV+rj0SRXyBCnz5Kjodh7edS+7kuRJnxCrotaQkYfoQr1cVbslDrL
NMRFzy/JKE5nDcmL8E4s74lCQqTRMlR0gg/F/wA9IKnsCWrr+EJM5RWGUeMh
+8/H6AiqjqpWXaHhwHThrWv9+G8v2nFxqhYbXiMBBnninEmOcuWMuOym4IPc
fuUBm+4mnikoQ/IMj+nezmoZVOT9OTAPjbYG58kCu4XgsVqscAmqBPJHzaP3
LXT3WLNjI757XwMHL/tGTboz6DhY1CpNWZSciajDbSW6lntEZm4QUP65r2A9
VgFY1Qfb1u4jdvdH0JipK6BIlk6RCtJ0UjBcanu3I4pliTJM+qDIVfKHNcCq
ue4YEMnqv4EdYr7+XtAVjKD5syIZPtI6iK3Ado1kh5cNj0XTjLmWZeoaWsAY
wJ2o+FaYwirekXs+uXLLudwS5saoahuS0UnXGSgNQxeCIwuykjl9e6PLS6Aq
TPqRT13a1RCtwF6rCXxkrxXINU1ZKTB1zBfW6h8x3OzHusp8OEqfkx+6tUZl
ii+zwi5dRxJm/h60GA962C0h0InMX9E6nxjcxwMul8Kvax+i7G6/AKWpiqF5
nhgmPWXZID0D9bZ2w9+nJ4vvb5w9bzXviIu0Y6ab4vZ2CxxbOSUDe/3cA+Vh
omr6D97eRjeZVq/w3WHUOO5/wlHRaUhcc8pI8wGfkvrdwm15Adk1ayWlpXho
yBOEFvThvwNieunGY4w2c/8gtodxtusFLjuPzo86UcYiT1GV2FkDTAlpb6kq
EN/c3SBHQh6MczjnSoUGPgtk6DMQb/wmJPa0rJtgGgW5d837vnd74vIhF9ej
CGhJa2JF2shimWt3Ub0AndY9XV8HjrKQWHEKkrlz3D9O+dLiy3GJQQQqVTHv
nsQxv8mWLXH5MTG8u639DY6dj8dHqTPXgQawXcR5nruKtc1qLUu102oQOP/7
JcI5r3IwYW8EBm9Jik+BhRQLCeT8v5ppYhq1+k71hwPtzYY8I51OhYdDK/te
jti37eluFA7yPTwP6PDfTEIN7+quWO/Z5WKDE9plOBIC9MvOskqp265fh56w
CYmvB0yXZmNo3i3ggT2oLF2lufmvVhmnDUYpDhBT+orLr+EAXgFY915Anh0J
QlT7fyIAYJb0BDIUJleazKDStiLBHaGoyZ6f3MehUbcEpTuHiY9yGZ9mkCJX
PKoRnAabHYLHeQa2z214qvrjBtYnmmh0z+A61lSD/XF4TtE1PT3eXpFvvKEp
OT7R3smiCDLhn83J8rGDRdnBjLMLh4MemuYfTt6NVlYuA7f2yizoZYhseSiw
SnULJLltnxZH/v2xLtTbQduGWFXKxAKAwqIgEJhbBFYcw2GiUOEPgnCAvR35
0eeGA41H/kxGc3LSx91bJDiLiKafHc0Tff9DyyoaPpLCPi97Ac32h8X++1k2
cswWI+K0WYTfeDJc4etISMalyt2pVHsqJn2kJBRY82435COKoT70/QNGQwh1
3NUi+6aKy3QSs0hXZU/tdUQBC7YUfRWPDeD397M5ONdqrj57iYK2xBZ3cPAY
lnA4EqTPJtM9w2bmxGe6DSJlajorJkasQf4sXzSCZisAtWF75HjJjrJNJR37
cr46WHx4JCma5FcCRWvx6bh+2oKMRz257IdFycOob7R3PJ44/UNlqHz11r6v
z2/Pw/4EMQ31NYtzmgbBLCpAkZuLT2j1vd98EHduPZWzo7j2k/Vl4K/Vm5u5
o0XWeT1FU5SoP49rPSCfvWNNTkVBc8tm16EYdBhsSrvhW3qhTxogGnI+EuBN
OfUJO68PL3LzpnWvCSnN7Ncfq5W5ljBSPOnD4tHNqY+PVugeh29vw6FQ5Kja
DDySF8e4SqeuKpw5Hl+b2g0tJ1xLb/RnpBLhPlylcEHXxN4Pm3mWYoJTFn5R
FAglbyZRTj6d8AIIg7M0VRABpHaIgqcv/tj4yeEvzDSGikm0Wfenpui1A5dR
ZlVAvAEjGmbCW2gDlX3at2gw2Rtqivs7Kvhw0V9M067H9fj0egDpY9CutXDz
YrrTiK5B00Q8eK5onfDZEpcQ8/4m1zx2YIjDw1UmJ6iQNLhNgXcrrGJ52EnV
iKUpGm3VRv/lVHd1n4tNQizQfiESIx4JQrtJq3O+47pArwxXKL8+JSKmNB7v
LIXR6FqatOfqvv9uykIY5VAgJILF54BgKoz56FMWfrMqaeJwP4qD+ekkmEmC
RXt3qY3Nu0SFHlFmOAhCpllM1wmNF+fQP/0dLTQvOL1KWja0uccIxzEob1eH
rKVI0aqfVmGm+O6ewlJZbl+STN6rhNLVxXt9kayUeiBm3Jad7YDdygd9clux
fnDPE8oL1ZiZOE794ucNbniSp1iqQJWUGHb6mBc041j+vwxOHSt1ox5NxnFx
B9JUS7EGUZi0yrImJz2pwcjXKtqsndjXAoZmuo6JcfkF5J75Nx0p5xxE/VfO
usWsFe6EFvBzcAm/NBnmiTFLcu/w12kaIMG0t/1B+dim9D14xtKJE7cbOMQj
L6VYEly3PTWvrCbQaEYPYyIIu4MxtZ6OoS/Sdlw0ON2Ol2ybHsB99Rbur5qv
Svqs9z1ymlI21MWqw/3pjST0XrpHn9ParQrocPIWPS52VKj0jC3BRbcJ4AaK
tWE8g4H8Je8P7+v7TAGFMeESUhn18qP2pP4JAwATou2ASw5peSCgXbX51nya
elPfg71oPSDoFFYRuEwGYBv0CmN5dbQADqdW+PcFSrtZGTM375OpVbB6//bf
fJpJ4OHq3R/BFwrZHGPL0r+P+2rbTmXYL2v2kdz2MLJYQdLGkR5LBoI5DxKX
YZHWU7jRrZDpVoJB3JTA6a5Cd6UlFa0WUvEZnRcQSKvVJpZ0QjTGqPkVRXHX
9+PoLnBh8mbVs5DFcz2HVBctCzraKqyQZYgmtTnbB2xOvCJvanKUGD5m3onC
yLnZNhA4/6RtMDBqAkPMeGUF3iYDkjQwIXVYuN3A0g01WBWBfW+gdTuOlkJG
2mo1Yj0jwTuVJPyvHBz/1drg/1gWYhZM/ofL9CxnDu+WmsEbEBGf25sTdrf1
cA9Guk7nUccGmXu9ncoyFHzQO7hQ2G0+T/idAFfMtJRTJEyKJTkZua0fpbPQ
/7/iHIBvRBV2U+9f6dPXfaq9k7ulFhElfjldEgtXFspraaP2U/I7Sk5BNEdf
iU94rbkiG2P62BJajV0uDbhbBiOXADguZCd0OLxfmyXRk3KQVpNGdINkLJbO
FaLerpP/gMknJqf65hrTpF3db71k2/159yABy+nd4xEO2rLO6+lBGugJLkAV
ThJol0X+pzVG1wVpenIrwXKJ/Fc4ZUKnT0LD9h3ciMcj8w6qVCB8+P0lEoCf
laflCZYfDR+z1AGFZ4JTmh8EQUtqkrGatz3JDiNMuqY4zMzDfLDV8mLXjfRR
INrdgDtM0rG1ipa1ba6AhB3cZ3Jnk1VfcBG4uz0y5d3vYRFlOF6vo6P148Ek
59TQ1jKvH606Ad52jfigU9XBzTWj0VowEbu6U+BP7F5LUc/vxcNZDqGOR/9v
ZHfUVHxq/mcy3NUyWs4nKTF36h8N1Qc/oYt5sRzRKUXIlY3vKjTfJM0TD+jS
xhBAJ48e5Yk8oy1/8Kkrtc5XKFO9gJ7tG/WSg+9ECOLEk0VuG8RlX5GPihMP
OH34FNDkL7eBJ/g/092aLjZuBLo+ADj34r6IfM2TNSgIQLFMSeh1HGKRdWCO
T0NqTcsbXZi5gtmKVZtTfUTF9SpAt5qx/Gz4QimPVBTUPI2OTOeUGD1POhaj
3+nK60qvfEmM7FFr2cJ75TKiXnARvt10h3tFJXQt2Rq0YIHBt0JFfs0W74Bv
hqnsIukm5JY1/3u5RlImAFEMdFZVROaxPWOagV200kxFOdIGDAvE5N0feS6s
4TBcJjZAtpJkX+YkIVC8uArXGek69IhQcy5vVIQia7AzmsqYeCCrBqEdSGug
LhyfKD0wZryebi1ZpMkBV/4ErerZFzriEBkSIV904jyLGhVXLCoHye+LlPzB
RMzvpZqKjK5RYZBAuCvb9oci2eDTS2NYknHMI6Sm7Tc0yTe780XftMYeAFM6
8qm5SthU+Aj+3H6obzFDuGHfSYAbaAN24ZbwM/+L0QxK6maQGBQT/gvDI+ac
XFD2mTo1odA0K66Jp/J1vAln5UJ1aIBP8Nw3oKULCn4gnZvBc2k9vVyEoS8O
q2w1SE8buQsIO5/4lHIjKsGYdcJgpjnBj3uv6Jk13cr0CM5z4UWe+6pDwSbz
Py2Ti0DBNXhye4yhY9V2k/G+kksMHVGhHp/FV60/0CTcruknhUAGmOI4+xYw
AjM8Jq3PWCpFDXtr+2Tt4B6Y+8i9cgbSnhUtVmTsSh1tVnRbbn3dhidspO5L
EFnSG4KtL1irdw/bfGFXo/yNvPginPf6F7GEo5diIOv/StHWt8WvG9q6MNw2
M3nmQ/n3bVTDg59pPHKBnNT6eYw4OaBHEWrpe38wTcXKWvuDmSqGZa5TNWiY
r9y4ITgB64sSzCjP0O10FgqKFccpPS87dhgXHEy+sw34V7AO+RX13etTfj2n
rYxxMx8kudf9sy8rz/WeZMPuvaRAttxztD3lznD8VSCnvUKoZnrqzG+l21lB
XciOgXg3yWtmpfXtzuO7m6dyYAnjwxQ2JALscWIsAUWybxXmadoPMziPNwd0
Weq1Hs8fRE0c8ctl9VttdBeDsA8zel3yX/VbnTzFlYv4PNWbv8krME0OvXVM
3g8FV6j1EgpNmn16yJwagrSbP6gU1QV+06IQh0Pk7ynTmdyScvyj32jrrgE1
CvYn+VePOCb/STlq1SGZqsMMfMZx8pvnRYEz2vkZIhgA83R+eu8sdPb78LB1
/gk0TIhOaLJWpd1srTXv+y4tOIhe2tDO1UO7OYhSgZr0s8UYJaZg4azJZzoo
xFrVKFKOHI5+vBnpKXdbNU+KR/CMTswpIRGnDHUSo0Gzy4IQuKpFjlsZfKR/
qD/jL84itWHahg0x3GDsroaBPsGGGG3XxeVlkK6GwBF1xwm0ypqCtdk6g5gu
aUMbAVcUXXqYXd06+wCsFTYxv9jHK07De5c0NkWLo7xPZxPF7XtHQF5S9Lt3
dRNxeuCMPMaBsG0kVBPblW4jS+K4MLKxll0SwROkf8oQkTKZFCujS7avKTmp
auzLvrwpVnTYNoX2G3EUhoY8XqD5SLDffRXHIwrZDDuBvsA5bQ6lf4NtNpH8
HP89TfCnZK0txeFc+jImNDKpwImI3003LuCjYv0/McWyCAGOUvmb+BEr9+nv
ICDxume11xOhx06j8Azjd1fVBvREf3r8Ym2jC9r1WqgnjS9+n8K0KV59kg4z
CxbZw+Wro3v9gsAQeevVyGrChQ0lJd5pizyCifjbvXyoLVyzH4gM28mItesQ
3MHZ8GG06vrEcdsAQTY9th+vBbA4KSw/1xJjt1Hqt3o6BpbPdPM8ixijaKdE
QJJapUGlI0MRjYLHHmAnZ5kQL6H8HfPKMqTxRwefgcW7eX76WDmDalRmxfvf
PJTHOfq6HM/JJuVp4OrClVdbOvsdMok4IWjYJjbEfD90Ka5ZAq+m7T27Plmi
3GVqcZRMdjWL0tqpEEbNbjfx1VJDhq80+lq8LaFwoCf6HpCBdiB6dKtUrp0M
X93beaEdLxnTfkNnwlcbjCb1IJ74cgIw5ReJBER83DHMkFgwqDN4AIocXnj8
hmJFhEz7a5SzsuPWnZN56IH7/jw+FaQdVC2j+VEi6ljSFcSejBE7Thd0bFce
zFAd1izNmy3uPvXodDK9gFI67DyLRaRnrcE22OgRaZvF71kVyRvg4fPwW15n
zZsay1vGuhmaEqxacltta6nzqNheMbBAGyoCNVfSc+jCH5mgGluRmy+Jb6Ts
8aSrdlfE67NX5QaiNscEM8ImQRfv6OHb/gllMUBJpATEuDDCZj6xPfyF97jr
E/BZ9RzbGwBZeptdtZlmUqGrpQq8Wuo5Mld66QLFV+3KYhEIeDLR552mqPbP
yCnGy9BCf8+JBCbBIDjSKviVShxxbPCv2tGovyGBKz+hji+/Myp5U0FOnn8P
CAf69aRTmfVQrl1VXpSrPF6JmtQE9fpvD1zblBPoSOcIKsckDX3t5UFmHMVt
W8swWj7s7QhcIH5vnZDfXqNDt716g1X7h2QUtmbWgBiadVp5UwP2QwYiEYqX
PygxcS3oPwYWmYz33UwEa+pDSGlBG1a2+VeoqBycK8axnnDC1fBslBcqMl7y
9GmIfepAxGoW+JVzq2LkPtZjU1hXwEScklWf/cx668cKW3FTxAxMI8EIaDWy
ePgsQS0AKzuhACfZMRJyKtU9afsh7svY22hfcMi6tWPk284UbJ9bEeskbVB2
9F+d2mPeiKQn+oN+30bfyQ0CKmVClH7Llo7kd1F4YQ8UahJzIUDcNwZGZcWs
4cZMWrM1yDKNb/D6zdEHnrj/t7hdIAC9g+v6PZ17l9CcH6L4MS8LG88Q44J5
4K17rh7wgJpsipiZylnW1JChCXt5CJ77KSvxMX6cF3oUAMv0EpzJpBfg6Quw
UgEDnWnRFZJZl/jnOm3NSHUAzDFRvCJG+f/psVIw6Gw7relzv2z7TsPgZcj6
mZgLqsdxYmXm4mWZ+mIAZlzKyYbk8d5Fv7je65q5AAQbbP9gAcbwZJGzeNJ+
UZK0TVT390xBDN5mWVvRYc8xmbKMfcEl+j9n3x/QDLxGlhYNc5q66lBXOdNR
YeYL4JkMyvjiT2jdp35+31D/Kjub5RAmz4hHSyr8zIGQgornPZ0C5IJA4uV7
t+XM3aJc+P3JrYJy6y6sbAU5KVGs7j7CAffr6NokdJdFnDSVrYWBptERa4TA
3+FFMRCnS/gpVnTOchm01HAzO11l5EwoWltcEjHAoTVIhs01UK+x7UE7pJSa
+/Ha/I6QDPQaicMT/cOpjuK4f5bK5kPMxrjMjFS6sz1ff99wllV2rQ64TgQS
aNRqtuvD2b405nYfQ0qMX0TUCEbL/z5lItfRYDMyZobtwOCC8WOrPx11wYWl
Z2VtXCAL1gEqsSHT4X+zAzjRAcphDEVkGj/om4QSFbl0LwgtbF2CJLmIRTCM
HPb7Qtjjlh/4jdORk8UIbNPJyRbzALCrHNfs8xt+iE7WB6AVnF5JNIZBRPqD
6eykCTXFh+qDbchbn/Qoqs2h3p36bAIPO931emPCjEopZARciJYSfyX/d2Zt
5VvhSeHCM+xCfrfo9Zgqx2VpDQ1LRS7ymsTukAzsWwd53XBW98rBreT54OR3
yzcI31mELsTozWe5sdw5d2RU40d1VNgj2BuKn7Dinu2xBaN/CaVeUNxiidQa
H7XiX2G/NXUbufoH6wNLhqz7Og0vt6fBbaxgWZujmTdaGLXcqVWSMW1T0goh
hVf8FHbpdaSdgSFlGCCi2gtTu8Uy5L7S71xOq9432BXvIHYX+T1Polb83zi8
g5UiNTnDzBnMS7AOMXiQSixWo8XFmq7twjiH4Bs6NkrO4T4+2yMfTcJOCCo1
XyK+thyYxe7X4vR1l5Ux87yCOm/v+S0Es4ZQzKh2xlPj3Vm/enGWyaKjK6lm
6wMqSygxPx15HGeWDzNVIdivPJC2DLoRnwpqkwa4ib+XCcNONo3LSEbB1LNG
fo1IzdOpJNwWDJeyuvmK3td89UEEWLApQGmXL2AkUXN1hP5OtrKkY9A3rxxU
zdOQ5YauPleSnSO7J3dQF+ydXB5j6iJbx/FVCUqc6x1yD8h6Be48wTcZntq4
1mWUozqsTIsM2Iq3AEr7J3noABvaMmd418w3wdSUQ0s9VH1k8WDISrVsNQQS
A1jUjjvuYCX2z7aDh8Bk5/0B7/qSHg4CIifgJqEwY1NYtEim4jGGowDko89Y
2u4omraLH9M8jOmlveMmtA6oaC/z5v98KPSQK1GrODDybUYbMPiqtTM9F4Rj
AVVVTqkjRTiSfz62lAoAXm8kJ5T7L6t9Pz3ZakqENqfs5fW0E94JLUL7zluj
mgbSAMZSRaQXAC0bZT7ClIIZbBLVF8Bx/ssjhXhBLHRywcnDtQGYHyO/8Y+t
AXeyHjUbwE5+zm3M03ODWQacdT6JwrapAt9jjrMTOWlTGpa8eyybKTkkKlV+
JutqHuXBwVKWhGbCxnBF6e4Cr7SpHYOjLWhvynEZqtt1GfFmttcms2rM8Jrl
gd0FT2UUY8KqGrxUKixHOxA+SX1ArSyiaJ0jWHA8jQUSjk62DP4GcsD+vS57
F9dnqhlC+RfyUetN9aDg9QWF3gXzsGoUy0LLX/nM/FiC6bedHdjuK8L6I1no
W+8S20EqBk6OScQajQI2hnFCxbheuEADXVTWULG8ufnIVZ//efEgkjDc5b2F
ut9HuT+FwlVQdGRDjuhjHK6MdcVM47bu+2Ft1qQK0FN7ndRh80ZdpOdZ3wsW
Xa7QCCNFJaboAUl15iQtuuHTp+SWNyzzjuJy8msRvI+lxZ77W8TgbCB3wvVd
mZ6r8KUd9saU/I/Xv2aJW6A8Qqi62A9XnzBkqQ7TivukjMaTiDLVk+OI5x7z
xzyjmG2LRsDyJET0tzoCFDcahZDrc2/Qa8PeqRxMEyCYlTRJB93YrYHZ3Ka6
HrO9AaWMAniAs/pmgC2Xo/093a1enlGgdhtY/b93keBw0mEa16EF59lFp8A+
3eMdkI60yaSY5CuwFeAhS72xdridPtCldEdIBGwMkc6smbxzLF2/Ajh8jFTg
cFqV2Z9ZQwnGL2XlV7xHGsiOcxOkUsIIeAyr9hGmwCGeiwGhpT0Mn+oJjLX3
kurwNUhLBvhnrnmEeYdD/kLf3qL9vu3S/8dao7dZGxwRyojwkm6YuhkgjGvd
xh+tiVxweELVtGFrsCx0eKlG3pzDSrrh83LpBtdrzs5i2aMIUp2gV5SMYQLV
7HGmbeR5MKEjLnLNs6BETNDaSgrFIynVpY4J9D1LGwN34DisJsaxaXDt0O83
iEYsDwhFP38+0V0t4SQr3M8G+ZXmd2C+Uo3Chp6yFV/06YHFXo1p/VE5ftbz
PKjJLc2qUix6EbR+Nc/6idSjbts7cF36LJeFCtjy+nJbVxG2jPXdGWMuFPrz
j6808U4pcjQtJgpM5KhUV7VwknNBw74MOtD5y80rvONw8ptAK4o8QoOEQGp7
U1qWIbdqmlenh/3Fb1LG04xQOlBO+IpiHvuAOsHORIif2qHy58p3kYMwYr2T
CTvPdclKmZoMWYNI/Bknu+zM86T/Zg1jLWLYWF4GJo/Xu/zRsTQNG8bAAvJR
MvCz9apouVa/Ac9/zCVqVL7miE5qhb4XJoT4paxK3dZf6kU2EDPP5yExJiEi
9ZHsw1NJR5RQIiIW7xl80EurIJhj1oMmj4WOtds0pPVbaLkiTP4nOwdICBzX
abOQ8bZumj1hQHnPKtYwAFLgGMNn5pxxdEbmvKS0P8euh43tc1Ye3aotqxvv
8cw37NVs+WPu42TOPTAERWzAm/isWAjAifN87kE7T1iZaIyfK+hmp6rWDHLQ
llH4aBk5jQJe7oQBmGgCJm4Fq219weaVer5pWOtO5SsIsH+yl/Dj6vBVEO7+
oYJDg5LZYTDu0veBAVms0UqJqlDU9lQbVNLMuzXPjlfzpVfYYFZv6W7p++mT
lCOvxzz+cMUbOm0V52CyMvknxShOKmDGQWkMm6Ax2vy0W3cVJMAY4ml3Q64p
zubu1tRh2WPvXOhe2S6nzJ+eaSZ8ypksmi6fQGS++oVwGDKisLSdLTGIQmvo
la/qkDbHK1nQUMYakfrCZcijGvSKFPx8bSNqd2K6BrbTgQQhAFQOi4p54uuD
AoNzG2TDwV4pWFvS2bWiFwTczeHQ8gt2re7G4YE8CoMoSMX7mx0vyEtEhbWf
m+vlEV5Ifnfo48cUSmPeYj5JWWV76TpxKfRgC0lOaktyJ35VHlSgGiYaCR0a
hQxt3wpnBHmZjS/OVVbRFodPO/AlO+MyogifEXzUVMRuKzXTetDeRDKhYNgW
h3Xow52gnaV5riogchXOWeWiCQNFM8pyV9fRIIC25sEoNuM26aZPjS8AM8mU
1KPIeLb8bFu/2heerpIYu5c6TQyrTWZOf1KzILg4AJ6qPpJhVZghA5nZC7o+
cCQAoRS4CLlCNO2zcWJkICXmY2H1WK7Tgnvw8ZTu91dp3LckQA/44E8lkWsp
98mbgFtLhsAObA1Ucbxh3b6VLPF3RJqG0KPZ6al2E7L/lHDaRmE9xqPb5z7Y
PDD4T3Csh8IAJqWq8JFxecp8ObCwjU6diX2rxNZ1Hw0MLXpt8/8dnt7BwIxt
tZ+rRtcflHdpZa9yA8LyjnwRjexJBF6LkJvYSYnKt2zbJHei2YWAsAPe6XMr
cPwU/jO6cpjwopzs2KoYJm9OPhzaq967qtB1Lw3CpbbhXXvV3oTwLzc21b8z
ZjbuQhmgVbIirHUZeINwQBmVZkCWeORm54Btme7uXaQHUXXdnPDiJdpzzkec
kYAODSGkTfKpSpvvRgOi8OOy3GUDwRxqHB21Q8h+JqpiL0V0yniVloSYHNAU
/CnIOzWe/yBv/EP3P9PPf3EGHNTtW/jStq7wHWjyWIznr9zRwZG1dhupgvqA
Gp+2EN8R5YErAXfcolmi9mkhSZKSq0n4rcnxtJ0qVauq6aAnHB9Mq3tcqmo+
R345jiDUI3bV3fg+kexOKx87MsqssZ0K1CS5k5Y4VMLRt6dTCAcfv22vL+JT
86Kvi1a+zj4A/tPrAiw8xj8qhgzbXM7K1vX/cNAcTJLm7I5qIPhAaHBJ0pir
arDt2hSrV6keyHc9Seixd833o6kZkdr1cBTWNSiQnL4uIdFODBRHGeaMvInk
4C3jTK23Cuk4YOY7rThuw0UMdxWJz0zgaltzPz147ac1KVB9kRAUHsnPDcMi
qtGxPITD9HzBcPn0ru1jndawh2E32rnSwSAhuH0yJm0nQJ8eWm1oSI3EK/X2
ImsC21qKhFjaFnRH1n6uXuSdx88hNQ4HgFvTcgwTBWn6DlrR6rq75FrKspZO
2boFXIBIuLp4eMx2ivIwbF/YpEfU+czHkO2yNnGJjuZtwnmcjwiiIMXnyErD
1iEfdyIGRDQThCRym/b1f+G+YzeLBozzMEuyAcGkfN9Aojfi7pyLtgJOLLKu
qjU2Ahq/amGJS4m2VtD7XLqcyWkRJR/4XV7VwBFXodJuIw/g0HmxjHEQ3ino
ivKfiDhwpeu0MuLrwSmqALAIm29mSXGlRwivZTqtw+AD6ubT4ZT4AIdPYkCB
PglZwUN67rtMHSl3NCqp1JYVstfhBYFXova+/d+T5mCOD2YeQZeajJ1t3ee2
QO0UH/zZnljMvK5YyyuJEzuBbnOt0bdixPneaifwWzzFG3Yhj+AbG4lev+aP
eYGBmoVvYLPqk1yAGNT54Jpug0kLxvlGsl0LwVk6FaVYXqSMAgsellx3iyM+
1nc+HXPcbHO8m+J2GnDh7YbGSq8S7Qz7dLosDIs+iW75YAa8Zn/5zfeRaKTp
0Et2SW1Ra5jz+s0d4WDaTMiVQyRpHkEi74fmstUPTxlgc5tDxvtdOgdFhn8f
v5HYDvWz7n+5EEE6GdsfW0RnPcEUAunyCW0ae6+mLIKMFdz9krmlboOPRbEk
YZqk7mVUUnMnUGdlU3TBJ+j/D+1ZK8TBAaq4N08z5XpopCKu+VPBdurbdotN
xLsNvrgjrlVJvc7zaUK6i4AHkqpD57g2dQ2MYqNXP4d8S5ZlUs9Gj9j+95W5
SoetBUSVwbN6ChpPcmSLbBpozQIPnH0ya95LZHRy9nRx7708bqrMfWIUip1v
8bOcF4BXh/0ybgc/myo+VlUwvVSg+bSPCsOd60Qx1f7p6Xg8eVZ2Icj2vizJ
k69drdTUA7Z91hKInSzO1jrTNTZmbK5I2jVsilfdsVlHXp5TYtzmvUrlyLZJ
EweEEuxxkKHHwYbd8UNbdfH3H3AWPHTYKjiuq8qrH2QuauL+s5HFXcU8EIu/
Rx1XDVV48o6Mdqp/9O1Xwtvjw53fEMKx7y/XnxyhsXrjoNH7u4tds28wzfWR
wHSbzplz79DIW+0EG5ihrXiX0WUzkocxxgevqA9tu67VRBuufxPe68jVIWNp
6a+zkczjgkU2SOk33alHrmlbQ2+8WGhFqFeALrAT11x6f1XzLXrf+Ojsy9KA
ddBZaAqNRsLG0bQyB03ZLORXpsQl56eYCFrk3P9PP05sfbofeDd0CoTUcbRD
elJmuOSSaDNTPppa5CXkpwHoSAwqJJL+gaHDSz+elVcrzMGz2Z2ZUqs1Q5vg
Cpdkjf2MeV6JCrRLd/hy0P8mXbsCbokk3OTNjf0fPEmHMHOUMBfa1MYgBY4p
MnP8tNJ2A5+ryYm1vauZ0qEq1aKvVgQ1KwNv/LKe8PqK1L40P77Sdi4dNBIw
pcQpnav2WpITEsNbQETcNaib8/2OQ5mW5ejlUvZwqp79ZAcTmNeDbaYbjELR
MVgTucd9Mr/1eWfqxgKR2p1UZ0oRGc1Lo3mVk4wdSzAU/3nF3L9fbbcydfTb
HO8MReemIkHzNHhrRJuZoQ8CO3M0jEz8DzqkK1362ArYnfnTEeLmvzqDbNXr
nbHspX5RJMQrwrJFVh4fB82WbLH9zoU7HKIh/I/gw7YuvXMGuatYBVrQKlE1
WJtStePzYBPO2++MmDmJ7Ji3Ovk5wwRttn34K4MKhKHPePIvq4PML4fkWvV/
lMPJzssWKRyrIXzBg0DfGJaH0JueCohGAZ88Bcgam8p1oP66+Kr/qiY6SFJX
Qy32TWM39ptpUe7B1Z9OV1IadM6+7qhtc2f/1ZBZP8/Uc8u/vsmyFlYuo1kh
9rPzKqkUK1u0VHhWy1MgD9cg2aAit7wiFFM1HDkFg1Jg4jLzu9IHbXxC8I+q
2EHOy5+Z9I1I8X/lkVa8r+NEhXoz9yVhs2nqB1btfkatBv2ryiMJ5mr+IWM5
QVhUUsxS+Vh+obXrT3+2Tfx8to/lZUOdZzggLzkEAX7CsHQqahp3vZepo21H
/jCHmm9Icb1gMfFfSvsAw46jrwFlP0Awof2lmKvdHp/VgPEpVLfzZXMxxfSW
1m9x+dAl4W7oxIRQcgKxwyc4jDTeP3aKhx/uLbiBLf7brSodwFF5bLNUpzS4
s53w2asA3OAZC2b4W1zSxUDy67oCGDC83XBrJdSV7SS079EkcU2uQorn2aKK
Xihpdg+NFFJ3P0byK8jonyNit6coQphRT3+HziMeGX/SMfDDs9J1lXou7/u7
8ganONmzvYbtzvBvwRlQaermRP7sJOEEKqNO5p2a9p4hWX/kxYRMQyQQkh5n
sP8vgakYtb3DcwKl+AEpC2JRjjUO/duxGkFrpypCSASopgTBEx9V3KfG8xHm
4ksse3vvlo+a01q52BdpeoXXmOMOHCqZPXEyJRXYzpED3oiQ/HLrT0qwd5UL
4wUSPnXGeeI6ikof0xYYcWSx3DoE4YRR0eTQLSUieiardPaqSaKg61m4Ntl+
WTD30sEzGRxTI45BRWy0ZRsaSld/Xo8+/wbymB7iQrpqlAtr2uB87OZLU/+L
64Q8kS9sVNCh0sBUAKzWIjl9l+Wd7HsHxzM8m76VkKe6tKmyolmSk/7639Fu
HQsV4LzJet0Y7UnYhBJU0lJFjD/QS9qNbCA86SaVvZu9L7mk2oqPWD6bCsuo
cCZfGKyHcWKe7Pf0WjXpQS+Gapsr4wjcWA933+oXVKXU5B86G7vsfe+HPTe8
b+Khk54af+5b5JxSeOkIST1W8w4vddWIQeNhGJkzuu2EgLGU4ewhDPMqU4ge
1c4KW1pUC7Zv3mY5DqlnhC7hGPU83OKTbCIImgeZ/YWK8rDWH63xW8jq2Yah
jFIDSLNaxckCzNJhs8116p9baHysUaJ7K1yfO/SozpaukxXtU2AI1F0gFlXG
oXUuZo+H6S6yCTf4oWVlnil+X9lm4ai3dxJHOoCoGw+aQ+KIQFrckRVuUbrW
LP38erIR2DbaKbxLowGF6qljVRg6qrmhqLihi6nFzRLDrdcOKq38FIqD6qDF
2aRwSlUniJK/zrurS8IbdH1g978gHdwXWldueAsoyz4gd3K6XAtA4ygr9bvj
aOFw50967o2wzZYPeuX8cpge5DGz3DVfEuH+LVoiO2NdO8eoPhH1m6aIpOZj
dx249L6xD5+32Ns6T9be0tevRG6N84jTggl81TGYVQ+/UIX9qGb0FJ6x/Ytl
n3Vxhh0NO7J36GaYKMDZajDEQSSVvCu9V7N+j1whgQ3kdFHFPMrAlnvxxMxs
Z0Q5JlzwreTqP27i21nITIKY8FU/uPsyKC5otWYRh2Zc0w+4VaLjlhfmaZm/
OlqXXytdH+NcOXFEmWaWjH1Jfwd0/FjoMA0rbZsyXMhPNTtL28f1Lpn7pyns
faaiQcoB7bpnmq0YcY37IYGUn4RcfrJC9lDt4FLECApjW1ORFsD4J3CKGfan
ix0amXi57sYSsaAabssQ66oXuV5QTRTqxdkbDZvudfmGauMWmz+8DZ4z3uw/
ZN4AoUaZCIMZ9FjWQgJNOnIjsoCS86+qycNIJ+n1M9JkOON3giMQRSs+1sMb
lYrXcsOwoJNEJ7uF3Xpuo0HhDzYQffORkdC9McmdQ08whhxyikQcLeVy2b/C
Jy7bdOoLI82qvKbVjh8j+fFMX3sjUnJpT4BUPPeP2Epc7Uu3o6GtsNS7kSfp
iKDrQZwhmgsV/KPwEWaLppXuPsNBFemeNhGqWDS49YkOlPE5X70hWzqxVD2y
A5vAT92ztD59ZFqFcQPKuGJ1dmQDhaXFn/0smpjAt10J1g4mmEe2rjLDWiVH
yhfBx6BB0MC6sv/njhlIUp2Hnakqv6SlqkXCAoi0MsZmAgZMSKT1xIyF8qM2
5KgEN7VfK7JBOVJdzJzClaW9y6ExPxcO1wdCVqtkMVnHi/eVFP0vaj/gPGZ5
2vHIu2DLJMDfp2Ap6527ZKSWfPqqKekqfKlDRn88c0ew/YEIDGBeFeqB4ock
z9n7DRvvJzxIbQT9mFUbd7ZxqtQSHt5R/6HJR/5NvVdJsInHdnxvsImJSBMb
cM3/fATpDi6qKQyofNHvQpulT+VDBInqqFipHIQ4BCv5CFjHz4jSzmhDZSh1
cXFgkVNWtOx0wfLNhwEQq9EPPySU5mRVDlfwXliiUHOiV3PF3tzlAyx4PWEC
Su+8Jit1j//7ZlJi55F/O0WG08Yhb10JCieT8Z6zG7nBqRqgGJqtHV9B3+V+
OcKnSrRYkTw2iYp/Iuu/0iHSKRFqR4k5qBKaKhjDPa0ByOOJLQ1RrXqLoE3l
iXRocrr6sk39npQjptwg9+ap8ufgMFA+56OjVlTGFWGXWJl0rUuCA6L8iLQu
V+tvdQHzTWpoc32rjY2IFY+2n8LF+EaqhbpsIJSRVWYJnQsUXic5AF4xd41C
UXzJq2LVItUKQagdTm5MRPNN3hH//ibbTMboSSjK3i4eHAwsCWUYLToTkZ3n
Dq5XuKJfOz1TBVlSUeG+W5YLWLbCEwTXaYNDC9T6CfZxDz+hQFJmJhyQho99
/iCbT69seKc9O2XlgQnO4WKRlyUVmE9S4kRiMZbFFga4jozRm7gMsv6ciO1v
9H4ofnx8+XnM2lg0kH+4yLW7J8jRdSQcF3fifFXMZolcEzr4PhDeDOiVJI3Z
DccKZ3WLxHI3PwpI9xX5G26JQvTPCowp7K1CRK777fwtXlSdDtCYI9PWFjWC
aw/fmSlTvrY2rigSz9C3Obd1l9M06E1Dq3oOdUfNaCCU/qNx1COMHsnoUkn6
yZuXC5yIuzSPTeCOI3BeTyHSp4/EI/tyZ6NtCStkhtSFvY4JVvqhHmWNnS6Q
9PMbKzRbdj2XSejVWSXmQ/tX6oKYSo1HasXnS+NzbF0nte5sckjPaLzfQa+p
WN0yX8W09zIjhuNtxaAD5aKqywfyXK8NKQKihVFxj+giwFdjC2qVAsyghVpi
AhJz0PtDMn7GptAu1OvNStvzZILBKN43tbfCcRUBS5tZoXIGndETASrUwkSs
Naka+POEVL5NqY5qbMST83xDC1IFecjIfvafaxBzXDnEjFw3cafLVZOJVfp7
hqgUYuGrzeEaqRLhU9bJAFem33saGJumNCk7kaEYtTzF6Vv7GVBZF/0FxcCM
nfJEJcROO/8nYrU2rqqiZVAqIf2foOJfA6ISGoO5gOfMPpYovt792jbwP/bz
FzJAvX2BgeoemIBEkG7I6D5f0I1pp0ofgymwzgNAqkGR2vfNHDTXl3gY1Z7E
oPGqsQJ+cZT0Iei3XWxAugvxF8f0c/iRb5zqyNJ2q4UXWGCUxN9wEoxLuaZn
ydMHMO18abslSy7QUIetza8qk3qOKaQYJdg+bwtWsw4bB1ndMKoTllAjVmy4
A+irQFxh+lySan1y4wcGmBiVsJlHevsTfuGRR2QXp4PqkSq6JbaYIeXl4cWc
X4ZFU3ARc1ZhVf9wJcJA9JwQ7OipFso8Ge53HmXqMXiyJU/Wi8UfZ83ikyxK
yyFslZM4ndueODE1dcPHh0e7i69YqQ5GNcSylw/9E9/7lGQ5VoHgR4t4Jgcn
la4sQtG+7ZdpdQzCv5cmeLDKKerHPjZlQs+TcCrvNoXl15EndNmoia2bsmaW
bCdgIId81EDPY1pQu3hOdGe9g1O/X2Uu25QUExH6ROSEQiCudevynv78+gal
faWovGWKbY6OOj9YT03hMYoJ++yaLmnpHtppnUqh7X9R73o+0XbBE4PHPbvc
5nJGSTzau1zHIpafkswR+5h86i04aRKKSWCc7nh9Y7zlOuIrJTQkmcWYFahO
15vOygzz4NnZ7jirVZhD4e2euwg5JoEQUFd7Ents+G41tU23HAa+kNsG2B+2
BArYnzm6bfZFayTtL15yU1JJAA4iSHR5nFgiZdKZGog9SmF1iIxpOAHom3et
cGAYK0ukiS9C/Oab/1V3E9C6OKxyfhohuua5liJJF+vw+wvj1dTof+50sbmO
n9pMhEJeK8MTtwj7wkLgrPXB4L9OmCRIbHMQHmSpDjc2PMvD8ido6DeXpNCY
t7tpmIH9UB5uc4tc0CYnMT2NpNQwm8jG/y41d7AX1mxyRlpAU5ifo9PHke68
gT0Jj8rWwzWvyR/2CRt+Lmcfm18Z1LSNsSB36eufC8UmFxdqhHnLDfzFwhEK
rkP4FgKb1wa/vjZM5Nei3xM42fNSgkOMS+gt1Ne9gdlK6KPXWZcrVG+4yl8b
iQ5w8QYYhLwaw13jhpfNNyaZ/ALqPwaAzg9tiqzIhM4e+bHmNet/xeqiw+tO
VQEBfaLEPapIMVrTKYA49sLF7UXkaqQ74CiZzRmt31HrvRfALlthlkxVLg4x
ymBJK6NnMj78iKPfAvTTl6Fd1OxIjI0BA4aH7r6ODjGh8mmkMOufnuGVnOyA
cKijNfLQ5HOJFrgPBRVts1vEmt4ooEDGSpJKuHAAgJXXdxPM30svpM5uFPNE
5rv9WNV/8o26ZqP4k7hSLbebfXz3As4m2iq27+6W2xC7u4xvV8/E50aGLIGa
2hmoSxe5nGReNBN5dYvWyPW46oUKoeikUuumPhjgg0qbcJrLTaGltx0bi1Qc
/5jgS2JgRiUm9Or42GHIdxZ87qtUNU66+3rdIteIht/rEK3lz2cKU5BrlmHA
Snax/9t/r1C4ZVw1c65ZOr0/L7lZIwUZs6aO+U1kd9RMyxJt0wlIm4Dz1E8R
7n3CpwdHLM05FlS+Yt+fL44QK5mm1iEya/jYuZpOJQoom3ULs2KGeBxSMd/m
sxqUmwscEbbZ29cNEr8PzGzXyNL8ePD4wsYve/EhnCrIbR9s0Gfol3RMnz+W
MTIVBJDQF5hSCimqKDft7EsaSfSgIk8UjfCwHXRCwwnh6R0VgONifusJklec
Zn+dNQ/5N9tFS1IewAnaqxEDCC0lIUc41PsXAdwx4qdMZCjxrjyYA8w88QUQ
fjZDI+yp1G3ePzK33d4qiB7/hCk4T6Pj9TZ30rBaRDQjphGCHgPK9yrTHfhL
ApmHNHhu1kbrK62lMVkcS1dL7j+pYyEh+YakyAnfPqtKpmQRdUH5NgMEF9rs
P0rnJsOCio0LgP6b7HegmNmRcws/Y9D4ANCWIbQZDJfeDMG8nL0dwo6gnLOd
lyn4eUylAEXmke3T+EXHVdd6biRnEVP5WU8C3zeQbxU6COwKwdKBcczKrEiE
WK6J5+W8yM/0iaX6530X+Ut5d5DiRDTtB6OQynl/S4965+XY/AOBnbRPijzw
X1g9E3SnlCh9f85ZtZ1WSuwxUTyp+pRO+YVFcMcY4lGV1WtWoPieo225uONr
psibTPHZh/NqzPaiYXmL1WrIGayA78Gf6XNhMH7m6vwhi095kszP9dK3vsSF
NuHPfAG3iBn5ka236zyOIb/GBW22Inwh108w7YsdR2RM3Yl0I1X/12G7RybH
XdH7P0vs3jmcT9iN4GJYMF5IKPoDG5kXO2ZlOXu9nTWdwfsCAzOvW7rKGbve
yk8L4DNnTBnX5YT6lUw3ilxEDriieJuCmFhi9WrcSEKneJpDm0ozMOwM/jbV
w7PUUpPbhGx9jt4n+Ie+urp7z4TwlTSs6tpAok2HT8zuyK9UVYiExI32MXD8
nSuBWKFD0/mE+7BtUMEa6HVSBAI8jyQSwTP2cAGyypsCiQFkBxkI1B7WzbwR
Pu7IqnNn09RCnQP7sLrh5iBgIh9D+yMvImsPDCDqMbtlkW83uqIj6+LEjwRs
I2oYcUtZJsfc7+VBV8uPH+bNeSxCgv99yvUV2Mgq20D4UjiZFJv5iFzKZ6Dt
qkdDA6JUGjJD1MHhoZ+Tvh85hEC4AgvDyk/5c2tCXX8DrEgWcv0+6LU13lAm
txFKkxnrxQuCFY0+j2qIg6KtSprl1UbxtImVx5fcIvqV8dfJsbGmjQT93x1/
tz1Dtaa3EiyxbHLUIMiL5VDQAAwOKP/WQL4MRjVzph4QfBXtZfZ4+Iftxgtg
jWnZOKXZehtiOq1qZEB/fPzwsywaKhpM9K4vkhgW8nn4pqnnwjoRfBQrzvb7
siP8GmB+Nbr15rxzElou9Ao/SirmA9HFoBgs/GZvNy7C7KbIJO4fx2cjUYKP
b9nsX47FZKwcSK/QywCI15MVhSe/ImC5h282klFudezL7VAeRrZpeT3wvAnA
D9SZDlvRWllgosZkwXzmQJU7/d5mzwNV1PLj8GpDbjpIrgKcqCm1ros+gtaY
2S3cJ7Go8Lhdb4dnL/zvG5udajPk6hKDeU+a+4eXacobGtdhIzzFfO6+ElK+
BqNG3jiYYWOlJj+OVcTwLzQ1A5ujKPfm/QhyOAQTPJoQpDr/Mepcf5k6IqkD
b3jkaH4aVDmAl6AW/EpVbTbK5xbHHxdrciqr1yJmagPq2opggUuPQHAIPwCy
E+LzpY7JtpmuDB58LYlyJKbvMSB2/OErkezzX1+mErasVQCcQTor3Q1FKsSu
bBLPFd4bPJBaSuWPcKGKbnS6mYX3bqCSjGvRMe6wbWXb+B019abns9m0jpXV
bc98wp22puUXoCFHb9Et/jyJUTaguKN9tDqgnVnDRgQjBkI9CsSBNg40uRhH
3jh+TjWAomV2FuVnAU79OwzdEA7koCa61q8KJrzArKThDSsjMoipKpSwiBM4
UPZFEdO6UBzVlH1QxV+TUqeslBaWkik9hSTs2y5BrhIih9Fs/+PhW9OqSGeQ
hBgB/HDEqf4x11OTYnNrKHGrG3QtjbO71LScrN2vIlXImkdqVzHrg6ilsvMr
5ikvQXaVsNNtht7QM0QaMI0UGXQZr8nfX/O4UfVCdP6BEH5U2h0nit9mqP5Q
Rym36GhOdLzuaxOoMY+igunauni9IioRcpKKrfZJkXyvtYpRw94yxWrDOnfA
0MV9St9BZWCBly8oEa3gU6xOT8aDOx2KveXZeid8erlO9P4CrvrjxWafzYOu
c0Iy8ff3YnDCca6v3ru17nQBEgM/lFdx//xsj77nOrMypTZWnXJ8DN4msZ/k
57we+4fnJFnLsFde+m5Psd1ht4jxsDEWQxb1hnfkHtVDd7E2c86qftz3f3Fa
u1ctxvKPvs3MxoBrygQ0oLk3mWRlRVGbk9mepnFj8fgKOzEN2bRGuwBB70hG
0vjXDp881/X1Mbi4DGPV/RAN/rDyziNynchO6WCMFTXFphOqpjy7AUy5Kmd1
bo4zqMPXLRUALu3JDwO1F+wy3FDcke8qHQfPHSHm13neOxaupxYbxkrPbb4c
cTlbNQoj0xysRChrvwJooC/R5+m1n5VpT2Y47pGfuK9if7/zhk/NkGQPoOwr
QYkFz7ZBWLK665iI+R/04IZ1VTfMVCtBTQtneBAzHtilmFlldMq+FeoS3g5i
WqugScAcXgtHbbJya7wwa3wFIEc8inWPG/wEwlcqHGTNpCMg/sjv5JgLNIuD
9pAC/+LJBhMxXhClv3nZDP2wj/JRS7nxIqQslt6llvDxu9glphHx+Vi7GNZl
qo3gxhruj/FDPzw2TK/vcka2cGW2PXaqPUExkGZw/QY8+NhxKtbLc0YBjKmG
A+iAPcaNNNHYj2mid8Ru9l7zTaA7BgWNkGELVQfFLxP917HyZR/GJntimVPN
7r/elxpA2JsdOThNfsPwu9HbapUiN/YZmp9FFgPxCEpX9xGv/NEuSwX82xVd
0yKtB2HhjlhHpfKNVyVAMoLjLSU40Igf/kfYryseH2AlFLyEjvwO6CwUgupf
kg0nlE8bC5skyPpbmgP4EHv0fNxuZ+/poYz3svLMlVcRaPaQmHfECyWveV/W
5ThcWbrpET5XzvnBHHtTTS7gHvhROCTKYg0mz8xUR5Py/ge+utV3RXc49Fqs
WEg/I/tRe0h4Xsm9FaUliBudhnGLdCxKS2GdgnOXcn4vlj+WHYRrKAhK+C66
7mdQQIGAjSfnTDqK/TsU+l7cnnPBBosejLJf/9eTJKcjXqbpJzLruzUehnBh
sxvcsuEa/6cmWOXRy3JO8FdjiCr2SYziWX/gX4MweY2xVNejAGo9IQU3U3jL
umDK4O+2DDzU+ZVx53DH2xTyYNvZlr9fmZepRuOa180lkG7BMNBPDme/d8Zz
/SzG9AcORFTaeiD9Rcz61ROxkixHQPoo6UKbfIrIduEUzajOs3whATjFHuUz
s8gjEdkU6+GGgn8CGLpodKYKqSyMU4xhb3+W7bFJliS267EnCsUFXdvn27Y5
mX6jVfoSTifNDOcC/m4YUtjBCvVlKKdeHvvPLGPm5T+/C0qvHjZygE3y29sj
bPUOv+BOA6P7Lfd+/mQucWj7W/nyeltoTczPqciYUBwhC6+bl4NM2U9o9kwM
ojXH/tCBeikrRw4xP52rxzCXUPgnw2VIUDIzAmVj23C9qmnsG/OS2uTjkN0G
8ABKa4AzeYqvaXj3QS6SRkHZj956ooM++6zhicogNqQzxmYiy9WZroMUtP9U
jkkDY5qd8wvz3ua158FlJeMxfJ3M61bFnWEXmvBMhZ65AR01OZxJC/APQoYo
q9xdBOjUVksvZ73xIHowx++1qGjVvRTqvcbwXDSSsCzIFJQikaeDM5DGQDyN
5F+g7v0XJrHnxllSX6hnUpp2E/oIxvQIT7J8Oio7uhQN0ylAeSZ9LzYk6N2i
wm6U8rd1uuY4Az3MUBDPlHcUR4+D7YAXl4+ygUvd7iamlS784T0mb/wp/m61
1Zq0Db3AGrogtOjUGyuVMb+IRKE6ScERdh4bKG5NIuOJ4i0MCnclhZp8AtSp
tcAeBJ/AtMUN7iVQ0y4LU0ftQMlYsWEOQZk8mI05q8mAClLP1b40a9TJ16Ui
eTcV2swkyASg1o/QHZgJZShLkmCBkfV4tt6Nrxt23ln2r5tnHEJk989StTQe
3vblAFMuyHoYwslvFA1f1j/zchgWTmNFWSemHkIaOO0RpaYeYmzgUhM9iFpv
+uFIkTNWIIOoJ9VnvaGSYCzsXbLrn227Sb8Dmk4iNqJRRkXyA9uP+2Shv18l
HedDUKRaS2ITehE0r8xKjEY+Jbxw+Uh3a3To8SivyxDA+xWSLxREtoWrqGKX
PuWSshe2u7HGjsPbsXEC8zgZTFG90aeuQVoLnNL/IMr31BJxX7DEmuod4h9K
QFHofPjDsZ8fNdCMULCno/dgznq8j8KbLJjI7DFaOIZvqpcwZ84IaJz2a69B
rRm8DX2rBT8OLpWolX6ELuCNPSD469/Ar1tQnRHJMQR58N15nupdiMYmamNZ
W8taWpTeir/YJ87NSEKkKynux0z5U6PxeTaRhuBc7035KMs5c4jUkUUQlb1S
kPGnHH9OdbbZGOZQWIyzTb3fHS4egJ5tGMBuwhd1HfpLN6f4L+WHsiQzr22c
S6mW6ENOz9ygrxTJn/FQwvDWMphJQW+zxYq9Npn9LqN7fi+NUftWstPhWQce
9awYt0wleunPsHmRnhIGR2EcAuPYb8D20E/8391qtwWEc2eHqPW3BFc8G7oH
HHMZ/wmxHPnVYUONWZEwg247LKMcfLN/yjaDUAArL7vq/yQxyoWZurmwr8vX
VedwtU+bkZYSXCscQegXufFeyyWK6w8ADdFLkWqWCRhcWbeoQsmSWEQQayGC
xkmNPsudDjHE2aP/tJWQMLzqaN0lrxzIcCwCkJTY2w+wm0brX4SHS/mHDmf7
/AiQszgHlRKn+0+526xXJusXNBz8SL9wQj7a1nPxg238+fl8IioGoE5rhPz+
/KhBEaxVVebXDIH4WIQyVmSneSbMVkkSuIGQ7prnRz5hnfeUbDoOPxY8e4Dj
oZJ5x2iEPb2Gd6Ne7lWrVSWLOSwLdSQxaE0hkGP/cZk3QvaDtonjVtpHO4GW
ccf12RGzvLolKOJKcPHsl9XZbLsotmvIWIfyU3zzQbV0hSvNrU4PR36IEsJW
kcOLB4MNfh6M4fkF4WsC9CahlWpJnaBNiAMsxqY21TnRc3zTu6WmSFC1c4bl
sQTb5QbZSZHp2Txx2GMBri9AuFxyymwdQhubXHrZuOhyVOxCOoop2D4GW//D
nAHui2s772VH2HRG0s4MXH8/Pc3TJo1xEml+6WMJUN02ZkOIKuWD2vtR7TT+
wfINqHZNoTHUQXBC7Dd1dQgGJQTrCwgeVRhyUTH8ptzt/+lbTLIZyn+avXlx
WHPSDYDWAEVHR7E6cm0TTbkLUKxtch/B/WjMcR8iYhLMYvD6MSmYirOxAxf0
sxtOfgatybCRkGYEer5X5+JVqsh8Ofa8S8UYbEbQFmm7OByzOJaKuPvcsYqG
X+BSaLL9rWn91JZhzxHgVW86cebydi2hW7usH/rSEW3KR0l3tnmc4LOm4wyj
l4zETZxgqrHObQnUhUW29jgA+7MHIf8vFv1xbxUKtXT2ivvSF0g21orSy/U1
1FTW3OV/s5Kphupwn996DMtR0HpHNJVM95U6V+pbyR8V7hQM2T9Bpvp2/UCd
SMqyRJ8ubx/7IQb0n//Gd+x8SM12LiQgUponEQcGBDYfFR0tPtd5bCl3zHt5
8fiFtl5jHOCWEWlv8a7IF1b7LLGvs9GAfRHM24HOMYDiQv/icrwuW06N9dah
VLH3t948ZS3bq0xHCmDYCiCNy49IGyWWMzpZyhxKMX2F4tgLdaLOWwZrgg7c
jDfc5mCwEFhT9a5lo4w7pB1wmkoNl4j1GsofXxOA3uFFu7yjmrZDNOqxishI
kvzeaq6UN8g4Fgvc1yjeVS3xRGU7nTeyVkdR8G0KJA53vRdoUJFFu09VEk7L
hOcZRz4qU3Rd8nC5h3ojti5h3/MzUXV8R7EiPwB89L7PBUtWbV+GvqbTWAh/
TnrIZvRArNda/cwcYILzwN64K/BI2L4LHUlLT7fZaOO9MV1qjmaajxOh/oue
ZpxR5saXjadogafM1igNulWo62UuHQpHzIMxs5NAKLXpE2MwTaPA6mwuK6dP
8bUdl3GULQ7/O2BvhogYCpiAC4HQkqkC9aecnmlKrP3EfRtnpf8WGFMHl9bv
VXqwwHLRGu/kiBgVRDiGF1T3UYrKaTwZYtkssnr4HX+VpBIoa2KK0iCAuErC
NBX+iCfyqwBnTDaAxXezGLg5l1q+tH4bsM5sr9Sx6uLS4jwvvbOpcyvmX4I7
D0vP+lBU/psTroUvEU52Fy534OVW1A7NNOHPW1KMxplo7vxfbD3QUUuZKPET
waWsdbag1opATb5bh285iN7YPB9P1MO+JGeyxPhZVKmRy1c96i+1Xl0NhF2+
M15WeOQ1Y+NK1A443FnJdN5AfTgeNJKnZaf1ZNYYN0BPjzghe1jc5IXnJQmo
qbQfBZo1EvNNh54AmJMOePSwepOlEoB/gVh36uaJUcGaGyPCdzj/jVd2LuHN
SEDm4F+y58xq8jZE5f3Lcl2+95AJnbT8+tUj9JgCXj2y1OQC27j+qTvvW5Et
NvEWt7KJVrBhuof5KPpqYmg6/ZW9g3AtoV+GKnGJJqWb4B7Fh4yXB1G5oVTH
Y2MKyZtpgQSmOkkNu4W1oxjqdSHoV4pihj13GLVkFt5wh9TAnYMmBHW0PavL
ZSeZLpjpup6Avjkhw6OcvEf8Ct9PPj43VJF6PS19t+78bjj0dasbQE2DEgdM
G7efBwXw7+OH4cAQqQVi4oCUMmtjM/IYWWD+2TflsBypFXXz4zLMMC6GaWdY
GvXaw/pEJiRDg2Y3XTqTGzo+6TYEJk7d4FN+E322ZOnU1harM7xhzemH0FVx
HnSkAMw/MReA1q4CvTanpa7oyLOP9t93gL710a8LTxL/tih6PStEp54k12xx
R/yAumkNe8ZvFXVDpOnGfTMJS4t/bTz5GujU2NEBwV6GxfwcMfG1hVkHTcOq
vnXi+RNSF/BVK24WwGFGeTCfOLsPO7E8vb5o8XwzUYzoDo68cFCxaYDQk7rP
wP3Ee4gjf5Mn4ZJeUbjY02nrwba0IH9WHh7br71bfJsuq0L7LnvrGc+ay5Jy
jBiXlweWpmzTqUJelWzvKbM2BZZCduPhz0DGvrzU+XUPP8nIbXixLBW/I1W/
CccTTUKRJJgSPKQB+tAbzh/7dN8QvYNsFzNIyw/h74/XXPr9x+jAiHxrLSHm
n1hsTwQwoko5t9cs8TQocavCwJ5T9cNiTSBJMTbDUJ+gOQiCtnQtE4blC9pQ
/QvKmyLv8I4PJGVan0RsACyc4Uix8KQGBah7Jk7aFbp3sVEEUVRnmUBV/Jcz
okeBtxZo/Crg4k0ONkCIj35KgIa0Lcuzme+WKgsg4+KVsTQpECQkPF6Z9Yn1
n2nXj7JfnB2RskVBZodUWwIT7bzhPdWXaTHOVq6vkYkHtTQ676PJhQ10vtNd
YA6tbrHOFnB7tuAe8yYVwbU+Bg3op6GgnwYuxgUdHpMZHN2oDP45oWVLs2mx
ZDIhI1rVAmjQQN5/qxGS8FsjDRrYdC1GlfPVXx9ToZbj+Iz7gSXBS15rfkgc
LD8HAYZ34EHlmlM2bdbqQxZQKgnyNED7y1okWbM7NR4LHP4nW7/ukHIph9vH
7+Y6oKshWsyfaZMCclV3kcdI1McAdNGj5pPAWjJxZ7s0Uw8FKISug0nR89w/
xRNPKUdbO/K7oNbGlejaxJzybQqjbNM+n8JjNyJbLqRKXUpxMeoOaniHA4QO
3yJPLecD1atFPdEwI+FrYpxSRLYWvJh1OGytapPAjbGpKpqDHAKtHztnTY2r
wvNJY7rIohR+wxjDQgixZW+nD4+lfIKPJ3WbjvhIHolc0tV9g2MNe/+lk/Bt
6aGeafBSyEQsLZDRKkJfwi+x49o+AUO3XlUxduu8BETEv4uhu4bt9CyhPAWk
T8EfxXev1ZGzZTYbuydtoS+t/0JbGU+/ocDuKS3OrOBmldBJ9lJLnX0XpO2d
5TXo8WifU7fHGXwuh8klMsN9oDFaHnoK3R71IjDWJDve94dljlMDtCuDFQfA
YjZwQXfTWJYU/05fHwwLQEJw6umWuoqHxTmyU2sC+7GpMKgP53NhxxdskG9e
QCehTsaCm9EQJr8SSFdlJPx9ArwJpxGlxwkIJX+Km5w/Rz2SORfTMrXYg2hK
goZgdZyVfgBkn5DTEcUyxXR/QLOeWcaxWnH3zL6XRD3OWNGa4MADTuDVnkJ7
Oxghzu4ZrZn0xJeuB70TA2D7wbN19g1uIekde1S6aVARGCgqkg8yhaa+uBuu
5gQSXccRCnheNV9ujeTLX0YbAiSX30eP9kXqRqMKfT/OSrAC9X4MbCRMvfb5
CsGYzu+6fi03yV7H9ruNwMQC2dTncT3+CQ9RSKJ75iI+OObHaM7C5K9lTand
uenkt6tdPF33x61mYsIyomO635E3Q2nO2n522kKVmCdwQuupWLMen6aoQpwR
4vsubcuJ5x9HWU+cO2QbmIeZkKqCmvf4qov9m9LEjwufZv6Ho5lKo8mAgTez
Ve9fZi9ub4JYVrr6ochVObEnbAV9VhiwrhjnKkjV6sm7xPce5/okORmWnQ05
XWO46n8HRDsXxlyDCygzbdj/r7y7xZ5OoqNne/K2fMS8T3rUVx17git3F83u
rY+w/BZpsBprpe3lwKeVq2x/2H8JPixRn0C/YPWW7k2GK0PCl022Z+VcsPoh
cyBZVvmK84nVjFZqJPdz7MB/M5xBFPYPIopo39DJ7g/aX43H2SDZm+1ojMF5
8jIpS29BRKs6I2VrvnVRN7fNEH98ace9ss3/eCEiqwsVnMcB4KtyKO9rML9S
kBfmncUIOKDUFMlSzP7C/bP7ueF+FNvxQFesb0+J9jsq4EkvgUn+i67+H1M0
4zms+yvUTT5yqnoxwqUizIUe90qXFW3EejnylHPCDrakfKLGNPw1WEjCsj5I
i6yWqURebmq0seEfsMM4IzkRULBg6xEi0bvfH0346UHRgtmpUicMX4MXkQZl
Pjazw/3CB9Yl+4T0DwOHSDq4FI+SJhfB/c+Rk2r4MyXWzDpHonfEZXqR1BUl
FbnXfrZlZahzarr0z5tjVWFNoxKXocSdPbFIAavuEiosuZwfwWLIPgGqcAtb
n0E8gG0Ot3h0PPh9dR16HbablXuDqhM7O6BbZ9AqvaIIvijjfcUoxtXp2dFJ
d2YAm68lnlMifdE4UFnGZoyy0NoY5WNWIe304T5BB5XLbCAFU30hjbohyfr/
0U6Hjzr//uQ5jU9UaVUO/LCh4ICM4d0JS70vrJK6SjbVlqkK9Ji7udNBF0Tx
+7ta2a6wqlYtWp8XsYeM0ZH7SSBqeE4dj8R65Wom+abbEicwLVqcS5U4sjnI
PpYvmPXrSzKhlyVouvZ4wXPg8aw4EyADHLud1s+vzYMPUcOCe1WZLzRsrk2n
PoT5SIxWpeQRQDk7K2N76DE/C+cXQnwVznqIC42ZqQqkdfkIXGpvswnhC23V
qrS9K1B31yI52hdJNm7MRw5YR6RS+4+XhtEqlkgv4Q5MZKqCrDLrWLK3wRoE
Q7K1K6RvutuMwOEEfKH5lKnS4NWeU5Jxkf9+lkqn0VogmENgCU1ieEIDRfz2
yBltK2FK5TShUTBUtUjei19uluK6eDKQVrCcWnj7rUaFMFCAyPSGWDaeeUxu
RTqTTzA+FpcFeZVWoo6ncSZMHF6iNF1JlHwHJlrAJyFWhbYAWVZL+1tV/Y82
r7ilvEVLrQPo6UP+M8Fb2l0zL3WxxT5PL33KYQRjHoPdz4GQdYcz83pplk6Y
RVlpXGy1wYQwHcdHlj1AWXf8cMfO7W/mHMjo4hz5KFV03/v6OcQgY3ngQBO2
vOyr5MLrZgnF508lZrxIpQtGTjHCVwZp7DdQ1ccnQouqzx84kI0cZHXYEhBl
le89Nclsy0LqGcgYYmswdhNvzub0bKB4l89c8cCb7K9pCya9HgYtGsV6UM8y
pUUHpArkAK4OJDipLFSGNDQ7ZoOZR35mP4IqDPc59oMzvMAo/sRCONyyCZrH
WE+6Gc4rxOnfjPVh7qn4lO289j8BD8KzeTsxkDRjHnNyavoc2RJAfccz4cGs
Rwxhg8nnKztDIho/uob2D6Pjp1mA1ZRXkJbN2m0Ehr9AH68wQxYChcr1xzqW
Yb4YI27UoD2YXbzVj1CEUaP9o/5QeNi1bfMIRF5Iy57+RRVXrY/2zGODFRqF
dyHsBTNg9ohqz0bR5sSVmNZ3rlNV15/ipiuL9GO+TEMR0X7aajm8WAdgn7Q7
UCyezMf8JuPVE1N2+Qp70eXMdkfUmK+7zDA74bp57v+nAUe3gIZjEVSTREEu
y0gDaJGDILbuxUvOyBmrUAC9j1LdPXPDoCvX7qCpp0tcFxzEbmxHCbycsjXB
EHDcmIPwlnDXfE+nhCsm32ztzCk5iMuUTzc08r5CCaGzArLeTKctUXc6C7Zh
lzFYl87aljdX9hBF1rLfpctB1ye8WEIrQAhRdglw0DiD8TxNlHFJilKIAJU1
isrrAmeXo6C/cNtdvKTSe8rljJyt+M+XR51UPzL+omYxYqYKJjA+ZdyS5q88
SF+PHd8X1bzwk+lpkFQ2txCDdApd8CTdfDj7V5TsVdOCWPTudV9wUDpGfD76
pZenYybZuCvYHI8vsGzyoIw88xiR9vLkiq80VNm2JRjNngWmBOsCiVBLCRWJ
is2IyRNVws5MYudB6JN3skFk3XWHlIym9NEfvv0pVcaRDSEgE/LQ+JgYT8cf
2PMm59c3QmSdRXPUnENXRjgJtP4lKUGBRer913XiNKZn8uGKWmlEVthBMXjo
e2Iy8SzuAliXBaF1GbT6wlnFf2aEv5WmZ6ch2z0C5135JWluICZkDsyNsnT+
92hBu0OWVuGhtYmE+zvVn4yHJwnNbvagWO+wugk5kaYn4Mmk8Q2/AFJjZ6Gr
CriMs/2QDM/KgjwPDUkNRe8p1fuSwiLkUx+ItSJWtQC2x8J9Ekr+qw3qAPIy
Jiq/MpTIF5klNP1O8eL6zzxr3zrLvspiyjgAzl3XZl2mTXe3/wN0k4aKrF9q
JamWGMEwSDZtWDQ4XAIhc/xr9sgKMm9mblQmsY+pZsyngoVt9pFHIuB+s8uh
5dO0+/GRuYqfhZrok2t7kEq3S/Kzg6nuUlATlRj1t4UimINASgITm3hdCSi0
Q1lJHoNUBBJPqGL+WdAqPh4+ctsLUhQwKYtn4BE2vHaWoDq5Nso1LAO+6gHe
gUK8IHxAU/KTn3yh9qQePexKWJQd6tvwNSgEondZb56S3ZgPelsZG8h9+HrN
H0pAR3/FHXMgrSaNJLwfhq9sli79EtsVzS7bFy45ECYuFfaLPoLlu1zcjOpl
kSPHXvRzdiOa/hA6O3xuyC3UJQuX57iZwd1kETTuKLpeKCgUw6iS82IzhcuQ
wt33BsGzFVEYOEuGGtVGQ7R+geguFJHqQo0EKDSNXuSfTNYd1cNrZVNGgmhX
Vvy6Xa89LZpuzQZQ8URYR7PO6QpsURPpd3cCw9qvjYqN8rry1Iabf7r6tR/t
3oNyD+xxGzuxWeaSaQLq8hrGYsOzwGeYYjHwfI6IEG1ijYxLF4dF4lu3ocj4
pyYpTs4atwPlUSv1Ba/O59YMjgONP1RxjosXuT1UHCVYLlmTqpdSg4fb0aSd
r+otyAezV3CybPgqjskqZKNuhOV/zZfhltRPGrX0xc3s9M0ME3f4cIMO4mhE
gmE2+vY7K0viBxLq6/ZU+bRpLUOwRxoVkGr3HUxOOQ/0F+In/PW2eGGyKmSl
LXRFisc4G2SYQp7JCYLNf4vKMlMETXe+pM4oj34LL2blg3OrRYsoHBhTMdJB
qeSC+YrbEfiXkn4S1ah8qdaVR2+2U+vP85uPbc8RE0x23Xzgau7LrOXqoY1q
LtvWkFSC6FK7foPBZxw873qF6UM138mCGSnFQniCuLjonKtVT6jJqXEw3Rv2
/HoDsCSTxB9E3Tw+lM5rYuxPfKV13ga+b2VqvgapqdKCBOx69cNQtM7N+TVi
w/lQ4hlmK9+Rgc8dad90w73YmynnPKYdznuKq8tx0IRu7ABLwjrA2cd478jU
LpgZpHdSuOxIE0UA0X1C2Mit2tnOt0nzYazHKmk/yO8q18NaX+ZIN68fccbr
dG9E/GxMMNxTS+61JiJRD/ZOAV2kjMH2Ec1r7m+XQCMaLBUd+UaZqjZLZ3rP
ImUkLEmuxhdYV8cqF6jVuwsEf42RKQXTgu0gDrUOaTLd4/9WoOiK/was0ohF
4TErhNeiujRiKIdszWQ2yEL6mvttojHMIZwKqgEWrEXSbLKUMX0TdvjR+voQ
IssLobgTeePQw00Tg20XMizRDcs7+TYbqbPv3Ut4ecJslUK9l94pdExTNh79
LfWXyNwwPrTDZQ/zSYhW+1HpYTVIpjPiF+v2nQ/lPV1UFui+aO4xqy8uEgDS
Vj6yZMO1tlyNTu92fqgYBcPQCWqyqkrpfXbnxD23paT6bjK8M3YWUQBPo9/K
M6s/98ellPBRzcW1DvVvlY+8i9tuNb2RHTeGO66ght3ypg7WY/6NqekOGrGx
zChBSh5JjLif7CVrjEZKRYxnUXAc3+dPtaCVSB+Wz6mkzd6xuafn7QdKdq0m
HdMnVTZlY0aUSfdCKNscVKXegqWKcugvaqHl2SifLRctESdEJhnJTJ7kRhMB
oMHmkGepFPCUYCCOtwdzY9S/IEKLxXD3UvGCMj3kkgO9QFUBmg5+v/pMVEzw
LDW2j1X2Waujxw6c4TwxORh0L3DOSSyYGGLDt1/tdrgOVOEiqV+OBC20p9fk
KEFKn0XCDPqUFwlPR44VxA++NSejidjRosGtZudNxJ9U0ZTH0jUcBkLiH9gt
9+TFGDp1nsoaOVTWVoK+puLlH5B/8nHvi3OknNrIu8KXt/4jIVWHe8GsFnFR
Auij0TOniYAUGowl2CMaqBs/MJFaY/HFPzlcsz2mCTow0J7cQTIZVv7tXtnC
PPqvkw3eMjvAIxHtOUepgF3cS6p0Cbs/7nXKTf/2AF76Le3xieFHR32qFPW3
0Qc2lCerdXtJ3+3Q5RF14imSO6dLyxWFIubPMTE1WrIwJtZ8beF70KvV0XHz
tFR5JFcA9/yUhpxmbod4LAXqIwtmELwyVdQ16nXj4foYb2roUBvh6n3aF7ou
QKrp+UMLShF5YENzp7BtSTaNz84FOwlbVyxErFnrFcS0KEXlVAka/pi482Lp
AQ5M6ykzw4y3GX8P//pmfJ1cYk3kX9qnD60p/EFoirXTtjkzYu1KqvBPDZIr
h5c9XR4wDQT+yYTrYnQpdJytLnCFo3FLGIEKoINctv+Mw+M/Ezb5Ksy4mGSz
CrbJ4cwuvgvdKGz8IKzGTKfJb1/ElOeLSVP3ld1iEnPAj+wNsgVcKWExFFwE
xMElS78lm8zq1g73IjhSWID9dpmgyqJk2IKQ2SF/kFrNSRPn+I4xQGrtbIOd
jfaWAlNYJ/DwjNjNXEAL0t1cZZVw6ETvo9Pv6pQjxRraYy9cHgP96ur2fZV0
/3HRs7diSc+YMJvhmgZ+QgnUlTO9aosK1YY8oLvFBZP3ZU3aeStuHsgvfEYM
EKdN44Evzj2qRhkm7pU449+C3yjamQQ37xkrNeOumRoLGLYemTaMBt9oYcmq
r4my01IozyR1Ss0RBcUy5ZzWLYv511vwcjF9+DJ1ShY9cSahfu99GVi00YNe
YIVf+ttrMHbGNFTwJfCs5D/qO4z9q8+nKL1AGzpcjqlQAy7KOhwm3Bg8rm78
0xo7BCx/RD6ty3f2973SRGIr/aO0idDCm4p5LhXZqMZq5LHDwhD6GApyRkdg
EmRbsjuxe3OHAu5ws94PAlPITKbpLdmeG4iX1GY3Q5issr2M9oYXOcHq5HW1
LHtYJFdvcfhvRf2okfUh6k8k/0utONaIKUpCzS+Bi+IonpiuG5i6UlQQ6Jwi
tKw1iEQwjPqMJuPnFWW+cj0LG/yBW/NDDO1hxEXgl6MbErGA+X/ZMpWVTXeR
WCnprM8ylQy5Hr8ultv07SDUgxUBJyfH0EkjthrgXgdKfBSengQfpUupcdmm
917fIP0RWcxAXMtLzOMLWDZhVO7o0cd3Av/BN5ZPfkTW6mUfk7FxHEcLMND8
IX0VLRC5PSNhWYhTjHZTXBc1/G+nFJsIqXxOErt1TMCOjMBdogXmWQPOKKAU
fV+8Mch0K4z5OS0zqAik29slGnd3j0scFYoLrki0QLxcoI40KHrz890yxqnw
UPdFfTNC0eg3METdfe8McsMFTc+bSKW4UNygjwLL3NmeNBrCo+iUUrIob0dN
XwXJV8bu+67x9LaeEb/HF1vpy6fKdLeAtW2b0cWPutFhSc6OpR7e2AyIczXM
cVFI86EyiXJufIMcLOCqbgadrK8V5zpKpfw+uZj7guiIBhp2r/gbVn9fhIMl
KqWW4J3kNyB3lDdLpnc2xbidQjZgK081mWBKLuw//c7zgDMgurHBepXSlnsW
AdO1rN7T5ScWAHzwQOCWXAUzyldZgE+C07diNbZsj4pYFTJ7C7ExnrYk7NvS
tXZuDGwq3M7oat0HsMjSZfAy6EWxhQ8U11MEBDkLKkjJ4g8NPyUwb4d3uah/
o1bI2aonj9IaiU99OhiM1M9wVUomUu3N0ocZZwRELZmg0DjlcXzzn8LkGnEr
5QJGFeXnMzfdLS4J+wUDWkbmMdN15rh5ABViD49QNsTkr6o+Xn1c+BPDd0tX
HN4bTNLbzoqEOuffuL2cNfXTFwn2qULWaAxfnhK8or52V0Bb0gaeCcUy1ukU
alg3Ikf+KHgWyc9iyyGEKI1+DkN0h/AYoawdJv4GMcKRnLcY57O+wQH91NlZ
DdS0CIPbBcpFstDqC3ZcnempZ1ikDpRotQt7inn5IVCjiXkaHyrgwFqX9gbE
g53lzX2m/lJV11aT2NTDoYvlTS7odbN/rJwSvD3YSAuXGCgFc3d4t6U+qB3v
UY8aFfQH9oKIMYO+6+IWSXArx8kJO00jAVk2Cxrt4D0HjgA235PIbvoyopJf
6psZiDJUo1nvV/BVfJ6T6K6HBndUH1iYhH1MQqUIrYiDuzYKnyTFzBdwqx0R
sqFAD/EpGoOGUnfVBikDCuLMhyAH8OUxKh/OcdZ+1h2VtdIL2oBmEKUBydiV
pPuI3SWYN3EZXeng+vPGV2PunbvaB0wu6t8Vqnt196MRrNRSj1v20+X8Yi6V
mm586fXcc0D3zPKF1OpF3Nh/urHHedCIFKqjcMoqVxIzOGkhqgo1nuTcjo5y
NgMMeGy+IP497DhDnJX5Ch5Bn5hRT8f9DDx3AHSQM28wQ5FT+ZZBebbjGOn6
a4vgTJGpUgL66wVW43gwgJnhS6GmAjx+ySyGz53+0oiGfSFORJ8yIWOR4Q1M
AkbFmpMP3ZpHZgSSJei1Dd7YgaXNliJ1fSKpXouisXJdFwSLT/S7SL3/ItN8
DeJE7+z0XU7Fe9hp8AQZSqVGXSA8Vbvn4B9SpS/INC7aqREVLm4aFPX9H0Gi
KVSWfsxULIGBAhfmJomwMulRbTt2UIUuh4W6J+61ONHuJ2lfYmC1k52u7Hg9
sXh4geG1Uz0SG+w1e6pqT/+GJoEmjkU782trLPNlHiW2CRKH1VJ4B6hdObWp
jRqhcsZPFhPtjKavmPvobuYPo6toKuswA9aex37wuzXCyWXmphZ4PcVpOke7
vNhyKKTDvqv559fjQQn/eD+C0MWQ+6SYkcLIodKRFjr2aBo2BigCszTf8RBK
9wNud06wR6nc04xUp13krCCmsb+kb0dQA6pQ9XrmtJnlt5h37O6o5EBm4Pww
wWdSx1WnTg4gsPwPBA9vNC84s9QIrdbN0/BnM3xNYk8jDJ0V7G29xQB6RNBl
nCCSwaTeBPB55all0iEM1OdrgOKBopu4HrZGWPuDahc+n56Az0sbQaGld2vq
01tzE37ocLYGamXMwLY3vy96GzkzP/es7izwkz+wMTHyCeacVv1OxBT2hJkR
xg2rbuP42zj3afbJfgENmdPd1+ATc3OTJv/73UgWqCsRpCNdAm20fclM9oYx
5e52eBM5r7ROlbmq2dbfx7XIk+px/bJrMVFDJolRg+nmxJfpmYZe/f1Kr7nY
u8XXRxNGTTwQ5lTPUkbnrt1/zRxvYp2nJPr6DoTHVjsf28ep6aVrGS8qtEp2
l+noWfPEAGs3gmJyFGb1SNQjMO1H32/iiGBDcXNJO1yE7cIT9n1u+ReGt2BZ
7LaxAdkm8raE7jlowDZTg3uGZa8yL5xfVf4AVffQe2yBXVl9tGIUvt2oXQvd
hhstoCQOGrsAIIzOQ8mz8HsVe0n5D+YnbHH/atJkJWnC6jwMQ5BcAOqp4EwL
eK228mVcILZcpQg8bqquGBkL6MNLBCkJFk6P6b6+kU/YJfXkM8HXsr9tN4XH
qkZuyEhvwW5V6iA9BPBN2YVpyNuNsV5N1sbPRR+Zn4vzfL8rek9ghK7RG4RZ
xyXcBE1By37fHuJWZmftjGrOV9DjG5RgY13CBkpEo0DU23uhqJFzatthYlKk
T+brOxg+mSPnTDgwiKhgRuQJYd5FmQPeVR3kHFxJN/0BNqSb5bJFnGH6sbqM
9TVW1UFE6KLGVkvMurvXvjFESOqVLE/mRFo96lqd8mSo+nm72HB0NkNrQy80
QKiKiJ/r3shHyTsSwqRIFXf+edi2x9UUOSKGfjPYf8I8HK3rejIWSg3We/Je
oeMYfwZgD/iyM5xjxdmGg2mM8mPu7f647jmHoPzTp4p6nYi5xl0TIxWRQvMd
zaQho7aw+PFQwFXfwxi7MMGS99GD4SRUyJaC8OI9DRMZGACqQ5gS+E4kOa7j
ZwugM07//Cm8dBYHzVf95zWK20sjGEvcrCCJRlkLHkgL5deKv0R9ldbryHvs
3o+yb/HqgG8s09j0GcLVkagNJB6H9fMn51fHW+wnav5L2vEVscRApxvi5d3d
BDAwp4kNW0MoQE8iwTdm152RctG7bYZy/Bu20+8bAXE4tzluI37ASxp3MLNs
aF/LrDK1rvcn70r8/9W7WX9q1Cfi70ic0ETRxUWBCq8DR9z13iiS9eBU0jlo
dwqfStqiBrz7MyUfBZnPh9TJyKJyrGqQRNeEaVgeGbg5K6VCZ9D/PR4m0q3f
1EPs46Wzux6yub/23NsrwSGjVC3VYu0fbsVLznKkt9639EiNfk6kVUsbG1jV
o6d/Za/VZEibLfynLHZVWszl3nFhiHKrri6J8ht/jOuCXN+krGRcJ45ivAg9
PuvdAlG1M+sfdiNSfym5UhH92R/02g0yniLpTEGCHV6vSGsmpINttYCJ9M9N
mCsVt5kjMSLMXnhH3qjOt/iq97RrAd5VunOV+auMO1OkNHrLT2hLxakQVMDU
h90VLcQwLZdolggOCTzGRZ3VEraOKsgyxPwzF3obpqESXe8Tczfp8G3c1+FK
ZLKmGbBZDBBZQhJ0zuqSXW3UYlad0xCDHso1uVZ7756DasLdpHTO2EdFmRS2
yGkjLeVIUlRWd4+1FXFcTz/UGG88L/NRAgEpiYteJ4Qowymsot2FxUJuHbgO
1xqqkVQ/pZxNP1/oTmjnPQUCNQPtpdJf8MWIAUM5TdeZGOkRvp0jEowcykRl
APXeH+bw/Ij3JBEn7Ft9wOJNV3hh2eiXVOcuFNdfTsfBQ5C7Sz+OfBfpqFUx
dE7N6nk+B4thKRn2FBxQDpTZn1jA+pY2NT/s7NCo37FOP1CcOARRNHviPADx
J41ZpkOZU1AQaq2FN7OZKVcKzP5IF1Z4HHTxX3GBl/i5lxbRBmg2q7O4QHHn
Ij4HZYixC1TSY8L58xqCMUNWhWEWBOGvSXYLG1TyZnx5eYaBWfoTzP4FwY6i
iAHQghDH4GYdYiGt8WNA4iC853/aHLTvNxqEiAZZQ3C132mQsAJjMAKeKKGT
xJ027olFF+IrHJ+g3JkDK4iTSVmPYSSR/Ae//BgDzBHPd0KHIGBCgqXlF68/
rxIdwfD7JEKy/Cf34GDpCOZ2+b7zcHU2323CwkuPaoeh/CkO6J22lg3P8T9W
kR2hbsI/mVrpP2sFRG7l+sgAhgFOLXmdkf9C2SqTu6j9g3apvnyNK2KtMbHN
12bYzd0aJW44rqpIsJ0YXSvIFyBCFg/8i+3cWUwfgez35XAjIZenIiCujjs3
SNBEOkvTh3Qy7vCijDNlibuzAilEfz4VFSqbB37eqUKyo2enItIUYZRWUhDQ
WI3dhtudX1Ybb0kFJa/57a6bXX05KZQCJngAy9Uvr4VPySBSZzbasgTx5Iey
lmhOAEcDBPjgti7jLQJoDYrtNwpohzvU2QtGcuPARxdxQAKYaGq8P0b55PQ2
JNzyBmweD2Da9xTIU3s/yNZf1XwqE4JNFgaxlzS2ozmw5DS+UjfVjKI0wukK
BbQLC4GMM66eMG1903i604+nwaVuCqeKUZ2zJ36K/SFGO7BnsEgo4HqzRhqQ
8G/yF5gLYK7j1prsYyYmtIkLVxj7NAsqGPce8+Cmf5l0GbA6Gport32Cmsgz
1VqzSje+eIPpJcTBX0IH0SCpC+lJkJXl5D7jjOX9nKpEnItZG8IZX31veS1F
F2xal1+5Zxs+OX4VtAMTPuI+gKWzR+pA3ee7lrbDz5ZnQmRkRbg0Ndsp9o5A
PHLwvlGX7Dku9CcGhq6c98v1bJKptxL1mZdtmYJmd5+tYWdAChvc5kWENa+u
Lg37+bSX3bd9P6hiX64cepiriZetdKrVKSVPeKrfCLGkfIgR+ffC8MB3Ld9/
RN9M7NA857usPnkx5HxU3c2tJ9C6GIPLfYNwFShPq2bDT3KzJXbbME/J+P7e
GlRRpRrJ9S5e+iQZUHraA/0XPSvH3p7wGbTdDtWdexGlWnmthpfkb92mnmdh
4miAJeAAQHqvZ+dU19QkM0NEU3XwMr3R434dRccYN9tpC04LvhZFp1m1w+XE
ibfucpD9nuqM83v21zvmwmizHSQXiwd9enCbunWRciixwT/jbRSE/gR91Igj
XxO4JSh4TaLJGjxA85XsEuYkTCLhq+0sZd7p1g3xBu7R3Bh0GWMuldDVWRnc
6qLg+8X4k1LDkKwo87LHg4po8GIRcvETl6A6cX69tVjMOTrNmHGNTX1KeIFg
vBzT6Sf/oXTMw/nQAS69P0eXdGEaDECRespnTnzAq3rMQ0zDXqXAkfJyGSOg
yN0viXhefcpzu9PKI5mwWTftVWtGTpwRuHjZOHBUT93RdrAhpHlrmmZjd5/K
OngCByrMdvMn8G7NQUeLcW4gKYPXBbqV/Sdcb9qe+Fal5g92QXC/ucHGeCt+
zjprMu9YHUZPV/uSektOiDWULbnY3NnZDnpb3Q17u864VFDts6NIfJfhn5YJ
e35ypP6fY2Dw5YB22oBtE2AKQE5ppF1hPjj0dZ4LtSpucaGWtXNKi9aurCF3
7liyGgDNo1eWH60FAGqXgUaP8ihSyzOx1qWMK7qXarQUVRqLEGt+xnAoJWTi
7Jfk9dA7WKX4WzwA1YlcAp2NemPIfyZWF0pk9aulh/D4daBtawQimtK2JPOP
LEYl82qx+q+dbOeCUaGhGRxCNHh8YUFXz4gPxA6cpk+ROPt1+LlW9VKC0SAG
VXAds+9FFPpWf+RZ7+evVeSxjofdqR6udK2bCtWPaIbiNL73V/8NSX5Y7AsV
oEqlOeVVzdC1Hdr8ZeB1610mA9PfAgjg2MZQVgYSjgT+pWygkjZ9lyZn0kl+
BmiuUOyMEnxqO+MowK0g91sZtpGJqjLI6AGVO7iHDwr77LWBfoU7f+GS2RMt
YwdPnses7K7MAo5n5U61boqTPyx3waLFdKpKlKAK/u72gr42+JZoonXyEWO5
ME5btnHrXDOPLlzGeCrhyb2V3NCQkafyGQWxmQe/uClpcMN9XJJxuFSGrzdm
21TLS/6tknJpcnU3DNgbr6qo5Kb5HP4JwSZFjDbu6N9bh1KHlPQxvDqkFbQg
p938eCHtzkKdJ4lORGVo+9eX0Qq5p2GCZ0HBe/NLJGCzhjwOeeA0IUtfBWv3
qPpiCh60Uf+4MKqby5MuUViR9aNhS3Qn7WEmwpwMjdT/IoHQBXReungeRXb0
stZ+9mHDg2GhJbK33rt6DtzJDqNGJxsGNhFxuYCan1upvPKFlN0KBnrvErgJ
R2U0IiSa/sJQ1AluIVMaxSva5FNKi3A0Ez7tcuMa3jAqKn1bmGkEqTOCAwgz
an/WzwsnH5DLnNB7uYZnnxGjfXll6eYfjrvqzl35ELQEm1/eSp4AN3cx2Fw5
jQkDJPUJNzvft1tsb5pb+akqClTyx3MD/cVV4AcVcwmit6O65j1ErvDDNXO7
iRrt+O1A5By7XCk7TF5ScvjWd8GsH/OWnOynUNLKYqHI66H+fUtqL3C/zoYX
yazaWmxf9+okxv5hu7N7doLCmOv0wb0FsmgoL3e4vV3lvB0WzPqQBqaOY06d
al71jSrh9Lq22Xqf28cBkxK45+NN7LxohNqHvizXClOZoB3FzsKOgjaw3d4W
HbH3T8t/Df+cRSsqR5Uy7VlUACKCMzxiaFZVmGSn0BHfzuNga+/HJ1iUgK21
mWrpfksNqYwsFnDWZLtQyQXRyF9AvWiIBWw90Du0YjLAolYY4nnh+n7uPMiA
cRELEolzdRdPMoZTSc5y+bJ34fh6PpRVUp1BStuwppol3AzF5f5N3Hsb8anV
3+PbfUiA0s8HtrLPy+sGb5YtptQpl5fUf+6ywCN9XnVNEUE4GmVZ/6Tl6idP
ZYB/yYw/0fEd+Bi8DFirLNm34dSKCubwKu2qxhYQq/cIORPTi54EcbJErTDt
nbwWafdLr/q8v4ARcNhc8UH9mCddd3lDOFToe5NkVDegz2er4JgmfWO206zx
bS1O7lTTAndno946ptN1mmIYFarHuL7HZ+pGnoaL1cb4usj/wZyvG/ESy9G0
EqeNBS0F7QN7OCWUs2Aepn3NGrdJl5v0LL9mKA4Y5iAbGJbR/tdYcQalxEYL
sz4oc6tKptKV+kXk8LY7C16+NnLO7dwb1G4i9tQymyE92Yc+kOL/4ORCOmKA
N3PbnbjbH1DMxMMRbjurTCRciLmKdggYcwcYMiDmoZKvPpF/2w02I609VlQJ
Ig7lPe75rhG/iHCB4zEDIUIpG+V3RUHSkzrpUAeOmLLKgngCRIp2Ikv4wfHu
FsXZvbIk0afU/5vO/FyPkcS1lwbMbahdilKAlbBregjJHEgIULdrusNmBsWr
iu/ZDpEiefic6Hp3nlFpR+fgBLKCYIidJN7OcSbDiTjxv2PtBnk+iW+X8d5Y
TxWkO5vL2mHiEJes8FMSD7j4WQIm5+HTFzbDdR7sZYuwLqH4kv2tCUSy+z1L
oG5Fzq5bMZ8f5Vb/AcM5syhicjG8XCQ/zgMCWVESZzAPHKWLQ3JcDqxKhIy9
tlT5VPkN4ZnV926h6SVV660clqzV+Ur2LUrfu5iZALMildY5ijwsVu6JOw1D
bAmmMmVK35S2d+r7zSBi6gv7Xzb8l4Bf5r9B69yW5NzKEaVzjPomaWYu9dG/
Quav1vsyip5ycXKujZ2CLNuUaSTbXxcqqrJT38sLw5YhDhLu9VpzR/XpPcDG
q3KKHoxqzMoggtwO7GfUQF/gi+CKRtcyStsEv+meBOjbmDKkmWfqqjI6Zy+Y
SAjEUG/fXP45LpNXtRm0EmGsAJkZDW88t21ObxEwvKATKpXq88rieIfB+YCE
ysNnxKcETXogBt8ABqy06ozqMtlJjKlxt3zRmUt09S2Qjwf2bmpO2LnuHYKF
Rvzc1PGKXvcDT+gAwCHxAQIYFd79hgUpddYa+Bs4SyyWooz1WVCuV/5uo1oz
8XbetE6KwlIg87xC5I1T5cnAqF3lhlK75mn/S3wmYI1nZaBHfIu88ChScp5F
NIAO9hc8oqFkmyaJwUtscw3lgTQ+V1oF73FvrvlFEuw4PDYl1JM1RXAlLb8W
7NOF0CLkhf18t58Hv8X5d80EfVP4Wg3zXFfX92nHRRFWTq3HeTeRjNhHtxC6
xaQR0J24UlWZJyIMrG8WRTqCZtZ1tfti2FV66SKEz23PtR2UrKb6zAh2FL66
4agWMrxWlZa64uWBlIo1tRo7So7T4Ck64c25DbHhYAuwGVaekoEoA4xjKJx9
Tdjmtf++7M0kCfvIvCa27xqu1LJ5yJJgYbqwBglkUvhHSBa9tNR9ZYiAByy6
dYqgJRGxNt02RyRiIzSlMelm57FN1yiAaXmRxN2iDJs/gvObJEZ9c1BHau6A
amacnU9gJqBIsOus48LNMtbfcBU2H+7G3oe4LZpRBIaQLKKLPWhZuDYzB1kd
xj2HcWWzziz1yS9SdBvWxP1LuthNHOq4WTgV2J0Oe5LSU3hVbiG4IH8ElH/O
w1Qecy1WoVe/4RnH/YTMtMIpJFO43NBj5+zUtXsBlaPdK5s/LD3idKp9F2ZA
w2uaThjsH6Ie8PGqj5e7jSF2j98e9sOQsfN/UVM3g6qRZ/vtTXthc/Wk6Jaw
ku6/5b6ieu7PyrTIZeE1sVxLkm4XpKQ3UMTkvtiCJEXCxoIx+WjBaBwzXDRH
B5Ur7F0BGozNOCh6/jy+ig3GilaSodE03UK4UyyXj5ntLxJIBwD8NZA1njbg
ZcSB8fdFXSpgjWyMNtMjxZlqAPM/SZFnRxm1Oz+RVoBU1/TlShCSsX8uh3oi
BMgyWiXQ8lFCntw5YSvQ/1LAsDInsiAv2FJlMFhpyq48vzfbnu9wIsnolZnC
aMZaSxY2hfsaVQGbO/+fFxGQNcz5Pw26stXBf84Pji9ZTOYxm6H9dWaLDtkT
cVps1gdQVBVUs6Ay/dUOk3GNHK9Rs+OC7rSyH53Pk14KPhTj7hGo6iuWyr5Y
J2ZoS2qaXyHQmM3B35xGVSn7mKr1FvRNBTy2b9tr7r8Or7YO+6DkY9tQMcLr
VkVdfYAPONU3sJXd2GhW49JTW3McvCC+KAd+VzW8MvFRMUFKythfv9SeulBa
z3pJgEVJgUUW+tOHW4t+Zq9WxOv3na2mZbQKMSxY1nyx7Z79PtPvbegU10j2
Dr7pUgOuZ2X4UG7LiYlciTuL99oPY4GePlK2jUzYqhQEQ6oOts475q24HFEh
K8K74Z5IGhey5p+u2NsMr5JcQQLD6L5Fet7d278PVNfGVYj4kfK/vB5ow4Ff
QRZXx3rji3mksakR1zZ5kSR7QAnDtkN1Uh9oVGAId8ItejDVhqs62qMb+/0V
yWStJEfrCfpKBQcr55A0/7SybuDJCW4Boe3VNwRV7nVNf+uFxdXUqvktglh0
zFcDb9SSVo8tkgxSCk9+HK2Mxu+dClvQFtX1kqLEImMh1IEiMM3/WYeJSY2N
w9L4i70MtJmKiZYs7kBKXcb8i3gSHFE7E7CzuTTzopYOtIz2KKZtoqB+1cdA
PDnq/gSjKyrczs1YOG7qCN5jjJOCYXihJXTUgBW9idObR16TkMhGaDoEK3Zb
6fw6pstvAvNZbOPIVi+Q97YOUC7G1GgCKdovgPfw9eQpYbnRHZRlcdYS3nMC
O2Dc3e6NBG1H7S/bpnzHqWdkq4twWNHKWTb2NZLnJ6loFYRxexg3GZMlR+7v
v+OcYMdgtn/askyTQhTEB1wuBtpiicv89XdwfNhPCqb1NcVG5nB27cDEh8pY
X1viytQnyTbBiCN9+UelJAOi6e+8CnN91hT5Sg+AFwXyi50cp3qIkDCJRd1u
Lt34t/bFcBjm2bvUFwnDSoDidowTynLpjV0GScC1fka2NXBcmGtfzmarMX/y
MmXv+2PMz9McZQkuXnug2lJu5n50TOx6gK716hXRCcHXTosFO8u+Eetgu3Yn
mL4oFL+EXApkvKGHHfeq2gGHre4gBGvoP5DkHLHVLxuxV1srRDjHDCVkF5Qk
kCBGxhwZFGsahpe260s4sWDdY3bpljYj5qAr8l3Wl5P0AYX8MCdCLgw4cOyZ
dw3DIT0EJLtw+7xaRpgiCwOOeCudnLeOPirpzSGIChbcBa/YnbnIps4GXCd0
FSYiX0QSdVEE5cP1a305CvVSja7hcdOfDz1Am5lZz+m4VQrBYr0id6MvrU3V
oxgla19pvICQwlLkYB9S4GJQ2A840OZBBvG0ul2KsL9WiY0aujrd1XIdn+Ct
izDyovopSmbBrY0H+5hLMLdYriqpULQ8BffYbuQ9yVVw9d4J3Koh1eoYrQr1
WePvwyaKjkEMPDlTLZZERZTEHbev85N7A3gsTTyRdLyRz572lD2YVbrNShBy
tR+rAj/q0e/iZ4wEpQ68Swt/2F76BAEnduDN0XwZ/rOE4q0d49LKGDZ7IKbg
M208gFZkacHxW9gcjsVcwh+5Dnd5xoY3TQbe+BulxtcxCr9QgeD5lCjv+FIe
jG0CPnntNzK5MoyjhwVRWd1hdAC+YNZzDbz/Wo27OLDehccQXwUuybH6/x/v
pjEQoMpx+jZmK3UhRlWrtfQRUupO80t/cWpzgnQLiY6mjiDPLdqYYHJZaoXg
pIENEqeg503uPVbuQjntkxp+tmjWquv7Gq2QD/+BjnvA9aRdPyDn/waFwUdf
64OLiz7eeBAuq+seyxn6v/7AvT3EVvqUV9Q6i5IElxp4nOypMaiNFvzUCoWT
GAojPuXAwQqFrMg9GIzWS3E4xDp85OOLNIDT69bnmFaJ1hEwS82eH+rMXtr3
8G83A2lb4g9H+pqsw0IrxlNVOiX4NdKm/Dq9lfyBE9S9FPZ4D3p4hXrqDxcI
YF43ftFZVBwO6SK1ZstS8Pmefg64Z4ss6T5AWmD+Sl1FCNTOJNBOLVZ3nZYQ
NMKpN+QbMwQQ9/whl/fvxbaT0TN44Mncm+DcmPE9robwJWopdGkesMOZtQAV
BY6uyZJpXx6AKipOmIljEZAab/Ox5tI1Vg9FmYMDv00fjP0V1OQlrMRMBxqk
+ts9P0DQbe69oQqBSou+uKPLaNkuoedvxwKmCPkSr73UQNyV9mYHwXRY9kdW
qd5FL+r5bu2my/s5vG7KHaZcWIl8ATYkqiO+LwQz4cpmk8KfLKD10buqO2gx
utkrGZV2iClmV9gWD/D96NdcI4ZpHShtXXsXIGYtq4GXG6NyjvXQATTn9Eza
zDj88yX/KjYR1f7oQRLn0sjUIH6Rfpm0UESUXZAh5VrNUVfpt0OUnS01+AhN
MU5Phqj6cXOtwR7dEe+s/MvvWw5ZJPaR6Ug+Fcrcf5vj1sJQxvL/YJyhNJBQ
HriY1E/4j0zHczu+BjiFygGSL6+3Tbx/oukfKg7OZWeoy6uTPLT2zxjj7JRz
c9Uh/QZLE00lQNe1lYC+kaCdCmn0fyjPFUFMdbiFQ+Ymr8+wIJ1IZMiP3uGs
0eWIbTGld0aEpekXBrCjtBbg1zY1kaFM/njPLy+PoWwROdeBQ0PYHovgnHe7
m+rTB3FVb1qOAYvCGB/y8YwrXwukRcOOPUz5GP5pIP4Nyse/Rz/D2y6ypWfs
Jdc9ygaEXNvTOggjumBLP5IO4yOaF6XJ5EEX+8SYZixcGhq8b5Csp5d1PAkN
3E0i6jLJrxQ5Va2QGQ8+IKDopNqKg9OJPh4JhxELmTQ+Xa0F7GzxNVqPnaF9
O67eTzVbCldhlOs/twbkoDW7jc+MZRwqfW63UlOYwSvkBi1L58vpyOgEuAwG
qBCC7gg91aZ49N1cLpXN5b8wQvOB2DN/E26cjJe7xBDPkWirdcDz8ApStNiS
SJmBwb3vgmKNZucdNtOIoHIakrBsSseDveMk9giXOptGfXmSZWBn+jNWCLt1
E54iffB7hlTGsOsMsev3LEx00Qh7vrJv46VGmUbdAg6bnSp9NNweiIdScADr
H9x2yvMyGwxfT4bW5nDK5HS+KfmuYgn9OUELIt9ZCPduG9iFIjNSyKWPto8g
/VXHL1M4qpg63QBJpCJBnCIQgl35ahVH/LWvBlzPxOc5uQo6D/7SsOSe42IZ
dU+WvisQF7wH2PGynsWwvhfk9qe7b6uaTLVM85hmeFShy9Z8asvsT5aFrA/A
Yt5K1me9OF/k1JPq0EH50NfPD3be4EFqVwJHsRd6uL5FHmDt1mW7CGIUmza7
cu+JRJ/1mWloJpUZPsS6k9psxMykpmpnrsid3zLSHeIwjBPBAPBuIiW0x4pR
AS/jLZqzlgspjFIq7Gih2sJtjBJhLHpHsK11lqeIdgjQC6DTetgZXrIGn6IQ
XcAFd9D3laK7ZUvVR31VQoJchl7EKFKlVjCImKLpgRNBCtkJpIwve9LB7AGE
NgFoSJOavkxifht6ix9up2OUjh01wbnbn300QgfBdifdSJoMbdLsXGTeOVRU
3ekYLkMfSoMwNxVbgxLKQytxWllBUgdMJuk7ZkUzkPPXqC/z52abrQwITnmq
q2O3Amh/xNo/UaXtq2tv2OaWnVfyJTzzhzEX5QI0i4qqcGg9m7KjXZDuUzhf
TuDdIVjcxIwv04kemGdkJVAOUv+NYwKP+HM2g8otIO3furkh2DVX+JNqs/UF
GF3ANFaLzyHAvQ6idDBHNlsiQHNHFCJHI/t7eTfBpMBMhX7t7fpiQhUeQcvw
+M9nG0ic8un4R81D7O2Pj0wuSizOa03RMG1BpfXxBop8kR/WPEiU+SySbxAW
JiDvYlAEGgrPuXDsc2e6qODCe2yWrUWQUrA58ewS1538LOT3NAocu+AYBElU
URsYEGK0SXVF3FIf3du5ubPmAOQKPezIcDIc4e/nHRXSzDRPtU1Uo8KKphh1
ab61XXNfjIchEqSfMMA3+JzQxq/6PxUimxEtFAqxfiW/7cHUotdTvMFOJ/Qx
2phc6iYDm7D0mVKmBC7Bf8lNvWs/j3GsJlTvUF0pypei02pW5ecEtxfacaw2
FWs+Whlgbt5RqpvaVN1DyzfojdM8mZiG4ZG+cEkKyKUHrCFhRGNSnNRIgi/h
3DQbk9DO6lRDFXqyCxxsCw5nhAHplvuXXPCjxrRMKucMxWi1C61NA0rXef5I
BQzsGsREz/3ZVlbLgYrjR45x0SHk/tOpg3tzKlmhiDClzLhhz7qlFtTc5T4n
8A3uJcYycdS0SIx/0jgR9gAOwLhuK9Wjzhg8N9/y5Ey3UMei29mcG8VHD87O
NMy8jCA2UjwSh4+vnNQdW4GeyiWIbEoEGHjEVSarnTnm25SwR0+3UOOTcHun
lbxZH3e7aDAdPken2XzcaP5ISRAxO4JwLi+soA9Koqbc4PMpXKzZFYoSMVFt
kEwkOqjjHt/LABvJcm7YnNsPDPFxq0zu0J9FCR1Lgx0DkzpQIevqfSW83pBT
U7pH8aKJslcsIWvkDASw+AfHGo8ckyF/ryDAXKxM6jABklrHlxcguRgOGZhf
+Li1FRvG0k4FdCdLdJx83TzNO/Pe6c2cmQzvc5bV8PgJMd7qpaXddqJz6UZF
aAKSfnq/ojWSyd9U2z6C12MpZ+OpvFw9fvZSFr0guJSEUMHtlMDdpQPDan6y
LIeULeNXTioMq47YJK5vKUy6x3QsvojzwbMJbNK2kpAMWaD30sD34gVxiWmN
k1w4ku7jQUL1H98BaSyY9JAEjbjliwwA6xrZbGWCpNBRcd8XSYeOO/qUZbfE
fUwLZIjmbZbqtsrRLHgyUbJRcOr0Uj14KKRqyhrchb2o0chnG1IHjzeN9uZ3
A0AKeh6EI36QL0jf6a/KVl6llYBuAb7qvpoCjXzMa1SS5iMe4e7h82vvZcYv
N+gwhtshuQXlirOk17qIAv4+DWL4Ss3qN6w/Jv+rfF9IDSCQ9MdjrFtkm41I
fE18GGx4ENGI3DJx5oblHdm8Us+TmBY9bpBDAEjl5w93Vm66n8pEDbRxR4Fm
CczRNa0eRwTAHWBdfHfSkzU0syIwJCpV6nhhZ1bZkV3K0AUywDHE9pGIr5yv
ez7+MYTOqtKPC0bTlDWgaHa3IDiNiEaM/Znuv3IT27N3iPmpt0+jCej0xjws
tBabKgKaT+LeEaTaEvX0vnmTid7tHGRrTbIozp76i2oxMgH0DEmSN0IEHJJF
FyB9Mv6eNw6y9qtbtSIEXWx5MpkFXOspwL8dfUCDVE51dyFndsywyxoRlpBY
EiU4rzDMgoN+aRZ05AFBhr8BF5ATA/Ebjgx4lCOeQnxksUuDxoN+or6yD+8c
ay8Z8aLNO7RGHVKpQhVPbCrMBR7YzCdgy94nzD7PdDMiR91J2D1Z2IIYs6AF
xwTdsXKlyMEonPoNa1he54vSMPOeykcSudtCFqZGEtLsqaXprQSaNLRS8G6D
k3XccUFs7sedQMh3XjsFdZ7L65yOmhVBe4EzqSqSEkWCrk8eRN+SQkIi6zdx
BVx7f23jXGouHt+OQTLLyQzA03iZJcE6FwZmyM8zeWoFZ3kR2NvzB3zUMe1t
Vf76toXTFNvr9j6l/9sBgkDJM3PpYHxZXclOFYwkG6YvepWpaNEQFMItECL4
5wKP3LpYrY80xpLqH7m3GnbZWrfiVPjcN+d9K4OZpAQXezTnXxyWDCqGRL3R
j2ITZLrn/jXpqCjIcWrrPMzqhqfAfZJ6rA0awwr739Af+9kyLCGFtvAlqs/e
kI63cXfmGaXeJTPlI18O+wHmKbtae0kZ0oat+l1cD1kHAHyqw/tbt0OISHP3
yf9vjSQLrJzNkCkBSsa5MLWqxpyITP00JpK2iuUl+MsaJOKaqUzgpbSvcx9F
hMJq/CG/0OOaHgu0BhoFs9TjJBzV39onQ9YccA3kZXqNl3RMy4JOLoB1g8vk
YS5brFSPS+wrGOHuVqIgMZYZFOLd4vcvbsF/R3CsysONyHIU3oeugLdTuUVr
TZN6cwQAgKQb7SzjRLUtEP8a3rs2iSWtBZ10xRIboS9sCATNAGLnz0rfhg4M
f1ldzrAy56A9EK3F4PVDLElb1sZnTMdpYh2HhGXbuwyhHYgiAF007bsjwnXZ
6j188JxPX+5ekGk9vpnY2BU5TKvbDZWx0PMcf+iEF2yznof+vc9KYJAMelxC
nY6nzMt2SKAiDh4uC8L4tYtnb+0Q4cw11ahH9CiQlPungSvnYOsw7M9JAMht
r8zl4wej8t/iT863d4ptRWr0YyB3XUYFn9iap4fWyLBIpMdz1QPadChxiJxl
5PrORZIa5gF8q5rHqvydARm1RNLrb3qRmsocbjM5GGgHbZN7MLhHv+UcezuB
NLROTqJM2leloYqzB+PfOGpWI5zSR/cIBXqGzfeyK4WeASO3Wzbe7ltL4Ury
JMxFvxyqlgc2zRDoSew1s9kMeo0RPI9Jbo45zJIsc8zi7ycAMnpAkXuKO5cZ
V9tDn4vPLso1h2zraYMxiw0tX1ChnQtkqdC8MvCC2PLzEHJVZ4yLjsHJDtaW
M3jeB93/8tvY5Lcc8D7u71MDg1zoahqVndpRqBSYHtH1qy3nos5j8ErL80AR
Qt/+ozyLixiRuV2MBzvVGcVy6mORGKxfU06JVg7CUI9G7iaOtRofA/7GgXfZ
mYnVBqHLro8eE36YlejcCKnlG00xmG952AkRcIaOuQRRVpaHaCAQhwWUcsDJ
NjCY2uWxGxOfpWKTU4+4rpUw55epQwkTrsGvmoiyIRZBKn0qUwN9uqzlq3Zd
8kddfkbhvmYWadgnSkVLylEE5t2u3ERzEdrznsvGKrv51hBJtn9NXDhBRQ0k
qVmTylLcYBsyXJds+917KmPi0MmeL9FXqlI6PAVek/ioYEOQTcwARta+ti2l
2IUvCNiQ06axnxEeZFpijX6qolZHjftGQ3y6rKZ8+gMuRyBK6dbV/mvP0/Vt
nFcxp7FjOxh9FZbFeWmXzHhgVrH8iLrm/W1dB8Od2hQe1KkK5sqMugEpBVB+
Lg77FPpcmb3msCDvqM9u8NSkoQQH4FvJ1616ICwkB/mqlhRM6wPDnsA6H5uj
e/eNQrt3ZCVjlckFJGeKh9GFXUV23EtaJP7N27u2Td7zx0DIXx3NW8D6fkg7
WsgAw4D/wbCAJThU4XuVK9AUcYmL0s2iBEBcjO13D3COs9GxbnhNntBlXLn0
AFxt3Ec8/b3dAgfO7pTX8eQN/BBMwWjsMsKtmWYWJOznXW7VEb5q9EnGVKLB
9zczs5UOlZEO53A7I+YB1ZN6/UceBrOOIGPI9gMUU9uAGI6qpexEMHZSOt5Y
R56aYzZiubQsmlRIg7qPJMp9oHaUnV5D9m35mGXXXfAwIHsBfahUtJY3SB1K
KdJFAE6RFuPRu4WUPXXJAClfqjbkYSffTj6OYx1TELqWysmgVMQ1159Nn5+v
89+H5+e80lQW5TO7bnW9pPGlBkjpfj44GjmO5NdebcfaoGYKIAlRrYF5Jtce
4fQZ00GpF1vB5WzkHO/yFBrt4U6UAkXUJlLsm9V603+TveSQL1Zth+mnxkzn
W13EIblH99gQaAKNkHODSCuhhj9OM328JpJrnTIcK1FY+sRl+EQyCYvyCgVS
5irBP7kzuBWUlOpYU8U4CY97WXbu2GX08saxeMIeKHZ/JvdoCApcwC89wQ+2
hpXSDHpSshzYzncXOYQv6kZT/EYYPVtoBaSD6NM01T2WOMX9xWC/1PWGMcK/
aUzSjXdFKKCMRTNosXDOfeuhLHZMkHta2beg2m0hHtKDmF5DG/OlfwOnGYLw
oBtZd1K6UfnuGo8qBgkrO7dpewPG0+QieMdw6EcrhwPDb7XE0vrJH4WVVbQh
hUm0H+7RP8JaHfJbSkc/lcxD7kNNXapPnJFn7A132df9VbvwtEI/3SH5owNk
4wtvVmS2fHoMOqaYIJdAYZyw9fO1nx5ei7nShBXO8+XZpuwHeIMp83X2ZGwX
6vOu6btlT12WYpD1B5qMKUOZlJvgSo20IQtt5V27RoHML5qJGJNJ6V9bZe2j
zOLYLYjeGwrXD1Y1tbL9I9XhyWLX82+RtnfoVm8Wg1JEjm3gwIlC82gtCz9h
BbXHoTWgXROGg+CNTtIEbWgI3VXXk+oA8j1NLRHxXuUNqTbY9j2Lz33yi7sI
wEGUKeEe3f2rfRMoNxdopBQyLp5pWWoUuNHZXodp6Du1aTUOJPrQR49IFuUZ
7alY/gjWr0ZI40IPEb3mB/XqZcXvs9rDsWM09XVVQO045XZSndrQUZLxi5mv
WG8P0HfWwcgKfmXOt5dD7HSp/UYrOVxCwluNcpVgPNfexNWMD3ulw8FAdJpc
UXhEMccD5C+ROLq1cLwiWEMzTCTIZtMpurPVLByZdUghxfdUo90n21oXE+ng
99dYVA9dS7QvJKD4SGJ693n5JNSzpj/qt/QPTUNG9tuhpGjql9NFTD9CqGiX
wcXlsnEIZgdonPL1tjdzvtpjuuIPT/I67Lgl+2EZzerJWLsD5hgx4xBcr9gW
/WvYt/JtGAC6/Mfb+qDY9jZQtg3ZBl8yHCEgsFTzLr50psODbmU2Cis9xQ+F
sTTZfznwG0Y8TNIlKG0XCW+KjUNNJeLju1Sf2r5A49vNA4Dy7gYpaWQsK9hF
NESfWbWoQSneZgAbda5lp5EBHlUXY0P6i4CjvcNF+EFpZC+F7KkqEIjfbZyC
ajmdZ4mWDtpzI1kANvjz6jkEsIlYdpGCcOLmzjKyLaDBfs/jo1l+fva3bjuc
jb0ZrV1ejRDzC8L4v33HrMzo1siXyRM+HiP+PfdQOmX5W+hFksvneXTM3Trq
iQfhKO2OLClxGA7w6EWwFxhGfBA/9C6Qy7NJ0ubwDZzOB9SEdfWoc658QVhM
INhqdH3PGP3NNlS9r43HRjN2jAOYGkYrj7M8OXtk2uMW/aMc7OSlWIVuDzWV
zkdYSljJH6ApiZikg+nG7tlg2kRN3UkVMxM1BfqGG55XFPiwjmC0q2EAQKAG
38Q8T/i8sPDbMilUWvkCGsOri05nxK3X2KOzyM4RP1l+A8JTlRV2PnwYMVrJ
H+g/ouxK3MDDdxdYX/sDxv8esaePt7KytUCdiShnDrG7dIy3mv7dlw+zAyLk
nK1FNZ3XUM9tXAfXdzNg7PmtaqC8eqRRk84oIF759pQRoXxWrVlVibOX94Y+
Bqn32JydWnmmCA/UAlcsDk5xx7t+LeAwpyuCPEtEY+Mob38+CPeq9/8TSPtx
QAHoSb6Wd5kx54ankUNuD0Tn8yEoi9JnfNzSNraTjD0T2OoJ4r22hCmItzPu
hxcJp8CtWm3GyukRn5yHr8J4YIxU0mSZoMlVnoT+FFr/8jWbiLFHtP3WgHKB
cv+iv2vlLUA2jQf/nfWvZz4muW9dTqHaRRghENYVALwcXBQWZogV58hjr6Un
gxdbuSqUNMlNP5qlFe1uvq9Vws3qzs3Hs7Y9Q1/CcUD1QGgw4pibqNBu2vTh
+k6zs2uDB0vkRRo0QNhCWQABr4bJ4BPU8I+Mer1uXxqd/l0qssidUnNRj0Tp
jwz+H6UCl3EeODGvkM42CGSMTFcTlKJzvNv183yZPso/YZEs2rRRO1QFLEAM
yftPRg77sLrnm4Mfl/7V2lzKpTxdzgI3l57dXuOoG4AZg1Xko0NZzwATqb/q
qNmcqgLePjPCxuVjpMEuh3V1oH6Taqb/GngLUo4AAg1PiLVBtIImp/Q4qRl8
Pc+vnfb1K3WPkg5+fHP6o6XmNUC81ExeYwlUlUbDhDaql+fw+Ln4WnWA3UOA
aYrJFMwnE/8ZYGWKB2TubiVKVDxtSwRI0jLMrW0cKg9HpYTkbg4gnWgJT+V+
r1rEKsdTft21JYfP0GG0Rs+l5rcImBUSoaUmf9L9+lPBeGoCkShwVd36YuT+
d2Apm/63d5hYStVv94Jvhw2C4d/XLJdUl9XRmO16JZ/i/mrgb5HxHqSjLEpa
N4QeARRFKxq87OWp7gV/+ABlg/26h58mUFVG3jXZM29irr8DcJYLIZ9Okecl
sw5mEx+EWTzGaZoxF0VuMSjE74Pz93salW5ys3GSXKonSWVGhNox8iBkHMmb
RRRhznHjVEJlOFOC8aioKexgV9rqPOc/TqtsgQWaVBrCOVnBvthFXL/ITOgX
FR3iQR8j6BRaanwW8Esup1vjPjaFrPnxixGeI+Yx7F8TFEp2/44/CmVIIjNP
6BhZY6cs1lmv37cIlQEZbP5+iimblfigKYMYBiFG+n2/gtiAaqidxxhn9njo
TvTFJVmr2ySyehHl5UrG/g1ptDyQvI3ARZcDNBY/KZsoz3lbxY0741NM8N2g
B5a6LS9hv5ss1BMQwtUGGUTLlZrS0BkYNMTvodsnGD8I42F8IDpjswgpLXUv
TtvhW3BR4yVQfv1tBu0LKGdngdNolZ4YqAEQ0sEmCuy5PX3cQIywjizIdZgt
2WrfWxE1VMDWewbyESBzfgZVFmqrpqfQzGG1YawbE9Rvm+ydMZezjBcU4alL
U6nPQ+qkZnZQeBqZaAO+H33Ff9IUi2P1sae7IbkiEmx9HnZL15dKMBAXr5j8
icg0OG2oxf5/C0lNhtlUiMWk/hu3ld8rz6NRDtJKZnVHmDViERj4TVNYOfgn
hTa3FT7sKzorHdzIf1AM/xjL2TDKBzRpQn8fnRzHaqjL8/CspBjJqMoXWQUP
WgOYulryO8j6N4HD8J+wQ22l11CreIGF2BEKhz6bai6uayrLYZpMBj/G905g
eeBgibfbuWxBvmY4s3bgtL2BhFBXOpYJaJvVTl1hnHUhFEd/JGjM+CPOxVhM
CVrRNJdG7qjS5RPFRJf5aHalao+owlBiAy1cNzEDN+mcoLuiobNlfVMwKnTr
v5O0QLeI3Osn9sUN7u3syq/+qmVg0//KFUIC532cZpmlLnSBaxNu4HzppKrc
0JrEEtNJE18+kBq6bJYPt0wXoygEoLNYonrKz8yGI9sRNzr9aXJMXVByv2HS
05NbRnEiScvyI8/ZPE5E+ZwUX48c5VrFQi39CyTSHAxdTgw9Sy1f+ORqVDwc
DC43s33xVe3hSnvJPoZv79n0qbPU0iSfu0yp015GA0R+FsrKh94EPCZJsnOF
rMCfkjqMrXpccx+FCjSkUWbvPO5xg20urcQlWZrQLqz4tRsMXXc11DddbzbA
h7FSs/mE3y5XmAwMaa0ZHPYQ9fF3C5dfJbPFkjf+4jHaww+OoHlD8sGLGjBj
LhnJkdwUtVfF36b7D48tyui3nsbwqMCmrWJ+0qrYIjiX90KHvNJ6J/6n6Oje
NpsCIyuMBpkpaUHONFcw4YcEGWMj7JH9xnCip0+xVA2BYjNQx6jFoCZR6mYi
8wHklx3mYEADaoa6YmRdaW4dxHmC4M985Ptviv+Km/1Tqv7iRFtNYh9iQuC9
+4art34fzZQEioFlm9SAK0VmpU4VsTvqRPx49M93na81qRSNOYczDdtx82bC
wEojkMFC+BzkNAUxcFNh74Bc0jiI9wcCw/jDzZupWYj7w/CUiMsl7lt/K5qq
4xy+NtQbWwUd8rVyDTmiEdVBbR0e/XZKoJ+Icgg+u0ngHTKE29UTQR4m95sZ
982ShZAemMghLdRfLqa9Ybptc+2FIY6+qNtdzowjwiRD3xObwoMtodJ9YOFK
OPbTDOulLYuhN8lddN7liscNYy7ivtToxLMUh3i+/vqzkew+FuWvUb4J7f4E
FikhLg01vk/nhE6/4b/NdTbXoD7H/zR+Sy33rv/tCSWXA/vsQk8bcbxhEN/0
VgU1BIwm+xNhQ3dWAIZ4hM/Tv8JLPsHoMW2jG7LDVb2DcuM8kgr+Agzg1iMo
0oCkY7QfSgj0ExEgiZfIJxDauffihmD0kyLimbdz/r8CAxUTmbDGeDhnHhfx
tVieAcNhxuOdhwTF2vV6c3SJk3SFH4kxVFEul4Ca600owXZYIkD3wnvkPsn3
WSTRuOTmObzcAmxKpfEG7UVo9YnAQaVItIDuVYrU+HaxanF0JquriBDzWyvS
IcKpkhdYon4Qfy9SE68jEBh9hDwvjHstVhT/pzY4FStIhes4k/bZMe5rR3Qa
vfxzMCK6yYO4FZgL7j/3FN1mXvtYNUF854YW/gaf0f5olYXGNjYN96jyhDqG
xCnzSK4F4B/q+zZskIfg5kEHX49YqHaXVq+vw3a9QFH3of4jprD/0vEGIH4p
dtjGvJHTMrWNTuIzzl3mEcT+FB+AnvWePs/r1NrZZBOMtBV/+kh4YWE/nv+t
1SNkWDtiGnI3XyzIxCwd8kwoI+hkPzbBKvM1w/YmdEqpLpUw0//u9vD0A/QT
ksEYMgHbNs3ULmSvrOI5yeFwqK9QAMRMST+LciNpq4t5iyCqg6/+Xp5m/ryN
Gavf2nSKUyFRmNYLbv/wBybGv28Wn6IJ3P0pI5ynNQSZkhZoHlA2+bIF23LZ
GODm14lk7wM7Oj6EWVHXWqqKwm6dE3XYBpTvlwC5QT8kCLvGc5znNSQQm6xD
6G4A1Bk/I8UHVbbTLcgWxYVwDXzZ4Lce9e24sDGxlcSPlyqZe4l7tYhQTcEC
1wWCmz6mgZXKyVapkic8Bb17cP/oQAa+TODMIL6Yetf0pQbolOhHOaPIXaor
Z5S+3K1w+gR6lddKfU/68gNXqqfNOvzQdsiUeM/GShbI/+Nh1HjzsnzvckYi
ZQUsjCX72X0uHaEHAYln0ckM3uktPQWOpaDY0mzKsBqhnAw++FloyI+XY5dO
3YNWly1iaxiA9SLE7zdKxwmJXC9nImrt/t/YvdS7ls8I2oTOXjPWpQummw+Q
QXdNaruJhvAdZPCCzu20P5N2jTT8r4diP5sj4Z0MouN5UmlzRDpevFZKRpr1
/ki8Dg8eJXjIm0A70n6QCn3ZZ94mLDMU9J8FonHCIzLpRSX0c09up2sDev1Y
WggWWD26h3byUX6QNMO5JocbYUVFzzgwbrsCofMdUu5hqRxvRZD2+JT0La2T
AmOhmTe/6s7YWXvvSSaG1bkQ/YO7MwJS2/mjL7D9kjF0P1mnM4k/BMDj+fWV
KN5ZJ/pn6SCugbuB+K+eTZ9uYrbsg9wSMFxiFfNkTYtU38NVLNObHMsh7vmx
TwMfcKjFawAhaoB9SdTYOYbkgEX8WuGA4Ddi8qrBrj7EcbkPNsYfC2DzRz9w
25nt8onx36cUh/UiJPuPzAbog61CB95AfYAc3zn1fib32gj4m0itEP17U/GT
dMIeMi9Qw8NYzjXkTjlfNFAk0z+Oow36tgHepIbMEp2H0JpoSYhEvJVYVi/3
CT0WjxwvOPocuI6r+8Wz5Ku9CSMCtdqaq8P7C5JDrSSBfVyfpmHknfTxbgDI
0QRWuSdRLn39Lmb9tVYfXkxZBzUyLUwIc+0jGDwvGK4vQjYN9M0WuAd5ty/c
8FyqbM55t/YXBq6rQwtjTF/VOCI7o04r7Knd2REVRGI6dBprYZVCLK4y6SpY
2k7Ny2YE5LURvGAhrA2e7s6Ct/Kf2Q5NlZ6MOFSX1qDj/SUtoI+dOiAhQ/PG
1sC06ZiPXC/PAD0Lmxxt2o1kx+h8gms83WpfYO8Ecjd13BXSrx9B8dXtaGQh
7l+9WHkNbuvkxPw5WDKGF58nnRmXLM4KAoje7mXI+W5W4RQoNJ0qr5u9a2Is
Jfi3byFIpfB63ozE1l10QuMYfIyFdw0Oiy1cKXXnZENeJsVNqhgRX1stfJBg
eT+UYKKyDrG2nzN4/29pR0PRD1GGwAG2MhlfAUYGjqiyfSq5HC09J9IrxIgv
nYJM8SghW11Pm8KEdOBLWZogS1TXyYYWe7sSNpm689d6y95RM9eRMAZyTJdO
4z+q6pvYZFqa8KRvkKfoWyihP0RITNhVhbcpcdKWZxIJOLQlrAWxY9LKWSkl
l37mne0ULX7lCXjGmtYgXjlsEERg0DounaS9MER1iflHktwEQJ1ivMYeOJHg
G7vbXgdcQkMinDQroAV1fOj4jmyyR+DqlzSTsFcFXXPzkvUkUKZO3KprrxsZ
Qb7J8fAYJECyYfuCIQQXyL0/gC1F2BKfOFjyu/DQYZbDNUOAdssttmgZmod0
Y7bBf26R9vpGfJJ/D3HYiTI3xOoYyJ+xSPnwJu4jlvX02DF8Pgg/N2p2tnR9
zKD5nReVtpB07hmqUFW7krkZpVOr6TFPs8FBKecrvbiw6Asw97owm/+oZGTD
wvQY44s+meE8iId7pjeiGOUdqgb+EXo/aJ0MUmtsmSZisCenFdDdPtnfVd/o
Cn83Kgnh0Su8UHmoi9iGPjH8RAxlR4cZMi+iKdtH66KvCcLzlvswp4K2D21h
TaLbrQYede40x11KK5DwPpG2D90TZKI/8/u+M0vvjQevYR/bPPCo2UXZ5/Aq
LsCQREwCxLTyTA7T2/rZ/RDKAF78V2qd0JTL1BEWuKsHXzqHCj235VmRs+yT
Cr/8zZ70PmSJl1sV4hoDPm9k1pzWzoW0fcJk0C0BReRO9SvTesfkPne18gbd
fDGQ4xQ4ktSBZp33hLtm8u74iP/ot9LDdLlIFtMPp50gGm4cSU0StbDcCwZb
MaaD7slMDt1+bVxAtaZt1Lt/kQEBFU6pxy/0e395RbFFgywua9TVGeZdCEpr
y5IWmmOk+xbvLAFdIXcqQl+ydKFTb3xUw+Hk1ix3OVEWEMrUatZXVpOqLcQM
espj+w52VIKvrVEaMGjTzI+m7S4J6d/ABolKTL3pdxEKW/5d/8mMcxV5hpQq
Ok1NpZWJGZl48lRVzvFnOaVZ6iyT/z5UVbfevclQPV5UtAl1iLDFXLnQFXoF
G4aSzpl13xOM6U4lfHo3l6pkSgHYTwAUSFNaDGgDPmtB8LhIDSmBQ5XDGUsr
+Bxl9K92RMr7o4U7G16iyJvUSkkRi+4boFWCLWjhYfyAVWNdo+HtgfOZm1cw
kXoTQyqI25VmvUikJC5ytsYzXCOA97mCdsysxFflILVFDp3AobJs2trB9DhG
q/f3k72norABuyChAKafpHEA4pqalcyIpEANKDg4kq/yiVXZc9epT79my1qM
VXWikCr15fViopI4sfUNlKzwevuHSS79z1YGPVz9cVUMrpaqiw4yxl1AIFJh
gYcacLFLRaDy73SbHjh7/hpeiJAJj8ijMTmTe+G/hLG3skmV2uCnUWcLd0Y6
gi2uM6QSv+vZnISWZhj6pxvXQYGd0ghytkI5iddypMRauu0douhKHJ5ye7TN
UPUXrpPp5jb2LrlWMHfQnGWHgaJ/U/sjY4ZFB3SxCsEx1cjI5KBgMDs9CfRk
1yJCX5FHzzMkn9tQbAugwbELMt+f0zwdJX47tVSfB/KoqPjAyTnJI+PDQ6Mm
BdY4abIUJjwmQjzLwAF3ZLDSkgoEgizRWR+1HbeiIKwe7RkwpsMPiBVFz4WP
Mblb62S0iWzqT5wr+TDYO/cY4QyhFny7MpblP+IaaZmxdVmaiCRf1kg7J/5P
Al2bj6FRCJcqzQ6WlKt0F3KYRFdBMH/D9UYIrB1FkenXlFzc7Wy7u6G8rwMz
8aBTqgIU1pWz9rlsB+d3cJbdYPMr53sAtvkTSmpoCLdypuqwL3uNriujMa/e
UPzqxnZI4tF54zGTRaPoZeheqehhxYfo34Du32G5RTkrCgq3s50QX9IThF0s
+7cyYOpeKxytbfZbY/fCTsh4jJqZ06s9gSosu5MFxg9B/i9uONw9CLXx1mhz
aIpgE50JJRgrpnPUkEPYuXCLlcvIKas6MNnzDPdOqlQq8UTAKzV6Usw62pu1
gP5qqDh0EJOE1PmUHLLcbFb/clDAN2TIJFSHDj4ZwoGEgUOsdiKpgD8U7uMB
k0YXGO8Aqr4DBi24GPrATzYLwLGEBL6OCCAsZ/VPSmfeue9nMAcBvrovlBG1
lYvR9Ns9oipLWkKys3rkeVeUa1BRrv2plrdGCLtNjxtuj2a6mGu6tC4I0p97
Mzx9qKm+Xaxa6L/nTAFs2AI6cbYCzCIPP9vur274+ZpPavZivGb9fQj+Gz+E
b73DDcF+mr3j77HUStOyL2FuAtVWc6oCFW1K+0BzJmTtKwNnJenWy/D8Eo3j
tXUemCAGVYHvBTkSDcb8yb4XAUVIbqhbK/EjLjLW8nTGJ1INr/ftXl1z0p4L
hZonI0psfNjPYNdosIAWZ+6itJ5U0x7FrH75JI+1DkUNCxLnrso2HaY59Gwf
P/lwRr9U2b3J4G14XjH/74W5G97OEOkDoWtjmqF94xzyss5XTsWDXDpt73WF
64IOd3IvJXvUrMyPRH/W6J2Z3GjihdQkwA0m7JipuWB5t8Zpv+FSGPq15NDM
fKgAZB0CnjYUQtCPRovefbWCI/HxuZrQIQIvINUP4OBC2AswYRsmRt27ja+1
gR/d2sd/NcJpaHYx+SBFLQIt+kats9MuvJtZyqsSLICCL6O/mbXtn/SQN63I
Tb5Km0NPb5u7qsO4qiCeOiIuWyCYwLPBB6lGK2IGALSDYBzt55Qj/Ykc5Uu4
pRgeedwNu9EWHoxbdveXaq1H1M0pO/XQzIL2lhb/UFkOGkSf3Ynaew3Bovi3
dIBMZeJuFrpvz6tlxTssSMvYFdg3FXBvtSVYiNSfHwt89Oi9mO/2GSM8cukg
jYBDaSoWec3pfdDGvkJsGdTpCrJdN7nOpm5eeZ6kMFz77FVteXazZ8ieGzSz
vcw/jmSgBcOV44JDMg34WUKy9dUYMAhD41fcF7lBp8q1auHevaRHQ3I+re3V
M2wU1sjnJWVzLAW0TGNVALR241BS6UihF8AR48zHE1ueyWZszfs+V+sfA52A
oi9bXUhOKhfH4l3TBN248pfsVA/dK9rT3PVbKJzwZNvV6znu4gG09ZleyqWF
zfHMf/9LddC+uaYBON7abYGFp7uugDiLKWnlk2nNCstRIzrgkq8uFh9nC1H+
ciJdpONMqhHHei9fD2E5zid/l9zqmXCC3PETLCFHFnwGQETIO087dUwlWaBY
esB27ZcBH3cDdZKzbZ+RLX6f78bjERNanCxbulWTH9EVE4kJPnUsusUdI8zF
W/NdUQsh9J4T6Q87mt9O+8R+1rH+qdXjTQcls3Lw+x8K+mnefa+aGLDnVxmO
CT2/cSnCwe+9/RwthOaaGvprYrWlkMfeFvZsVsyzRA9bon/+mg0RrF2FhB2c
WY267n5vyTVpStwzDsr7BYu2TJMipTb818BU/AQCDP4lSU9WZR1ROxeXP8SQ
3stlIoFFH9kH7aYWyZnVCNr/J2EFlkJRklLc9TFmSfxI0C3PbWg9kGJbtE9B
QsFGvGuGqkb5b5qFWrhaVfkTG6turBV9P2pHbVsFlboUJDrcrdAe/tIu55mP
GYH8HQp+C40HrPJerVqdY0mQ0loZmv6Iw23++nDnRmYAROiUVFedrAeybyzM
KPH68QAdhwByofduWebQepvfwnt7Lsa4mWMaQ6c+rfQJaHalrpBCHlJ1au7v
Po7AavL/UWnfes5eG0nPkYGg+uBxjAnTjSwWCs3zlZlJWHk+d66sNRrKWyPm
+ZtVRkMLWIrzD2lo87zQOHQm9gWf4MDjLBFHRjlHCqM2Pl5DfYR9a+dgPf4C
RPVcIpLtObXrY2Z3S+YTMlcuHq5BfakAE9rmO6SgUUsvtgw5h8SCmFtFx5Zx
hWjgBoxS+mzZViXKXoxixKaqtEilwmV6HqGT0V0c8ST7AaWkZGNp7G63oGes
YsiJlVNizxe9p2svmMSxMSHf3ix0glccJ+kNr296FEfYbiR8MycaEtKf1mqe
4OG4qlpxVycFr1nu8tlwRgT8JhQcO4fiqQDCJeaNcTM/NFNasSn+kirtjvNt
6qpCdtVqVgUozr61CeVJV+wiDfrCGluO09u7nN+5VGJxQdJKBUERU0tVnSua
bRucYkxQjRQW2eJlteCH3DZPgDv1LOAwRT4sCzBzIK9kBaoag15wbYtGucVM
ShB6NY3saUzV3G2eO9NnDZ6Iecg3xRMB8tg3j9j8CpVPTJqJnL/8jBBo3Ku+
fPnnoaLOUObe5HaImQQRWIxKDDbS4G90VdIA5qQ3m0G0nK3fEO7C17s8n494
UiHYo0QWLFogKH+8jeLAdn502uJff4SoX7D+zY9Ijm6e5KHL6ilyq4md7jM1
gT1U4C8AESkd4oTY5cqBV97rLTgWhw4XnUDjDYgiAKq8he8a1P07digemE+j
JMiTLOCjb0ZaDFkeSMBvw2ayfNGgoiW1nwmC9wbM0Fz0hWB1Ii8WBMc1kJl7
8rbXG4vchhC/PhhcX0nXrH88MHyIGhXCgUtiC8K6Ed1/LOJXLezZbwQXen2E
ruDA+3BrsCe8r/BYLJlOeIwOMsuc9m5JOpgT8E2nHJqzTX9gSlCtMfwvY5D3
3+yINuEFuYPZHxDmkQHGXScBGpwJF7XhS18GKzODBMpmvCm/JWUjY1e0O1Sm
782aXywIbYrb/hUDQHKbvVfNMgfLdYS93HZFAGJm6DZuOozJdwP6q254gbHO
oxlMsD8Zkf90lOnO0Sf2CAME7Tpo+/gme6xjqaoLeuzF7c7byPVScwrL4Ts7
xyoG+6L4WMnxT6LQcrzGJ7YygoP1w09UNrQT2kRdf7XFhCe//M3vbj5Bkcsv
j+dwqGMNgIJ7vRjENhFZNAj90eqIxaZqKobQE54Kytoxk310cTrQXr6Kl0gt
vKM0vsEjRuX7WWj3R2iDOCWtC6MmeM1+ez4VezKv/L1N4YHbKiNzz93aGfr+
ZK2Sys+u82LKB0imihrCmABtW9qluybzhpQCyo0qThTlcz16/wad7Sr38ExT
kshzEe10gtwu4V6q81eLufWWAKyBQI3QSOCxtaZwyDKt9Guwwbvo4DnK6nYq
0k1d2h2vPrHP5mGdTOlnpIAsfFMqz/5ozsRqpMqwuVLWEKtbMR02FKkyqJ6k
BcDY7LigZzRxYaib6b2dDRV3YlOGOS3/jYSqgqYGN+4DCYE6iSuEh+ggMOC4
0iIh1BpyiZR7/XimfEMxiamHVNuTF1CqXMOLH8syImnfe6FbqwOHrorGP7qa
GmzwMD3qdCRbX4Q9xPiVP570ggSxdzjeq1L9bNOrVrjdW6x3g0zhPkznVqfO
BB9bX3jJ1Yf83aOnnkSKfQvw1YqqU7ECw7aMFKFhz8HVpqIWzoSuV7vhMEzP
rGTX1146jJ7NNM7XP9+aOUynZLVXELcusqBobYuLJxpkBM53Z88LDIlKp6YN
bTJZcI+DJs4TvX30kpS8ixH2vricHjTy+i5CQPSSl1BbMktgj4exB+jSvysz
YONJ3kvp3gImuFffdVoZy8r6IofCWiz4psEXANLTsKrtjEAquC5Du0UdMdZh
HhQFgTrugcj34lvG7H5NdguiTbhMpDSg+FL51dxhagVcQQEyU/cYAlU6JYKS
854YOe//IENMGiylr6nBHEbAGYltW0Co6lXOIq20bi2qPza7amOCenYQyIh3
j4coFP2C+RFCSo2+ZrUf4UP23lItYSyLC07yQTNy/uDWk4DOVjLwoNZ64Z21
sy5mlGGOVu/kWwbz5rs+xF/NkIRpDvV/9XfVWc29pClL96qnztpWM7bdtegG
w0J7nMjhvJ88pkvMEj0sHwz0g2VvTMIXpRLIccZhYg8/lzlKUBWVg3oO2TAP
pvE8xOF7scMUmy9Z3kZWAIEa3N9DGUtNq2n4HSjAdTx35/XPJlWKgpGRlUu1
TZoUxjdzYH+TZ4UI+digzNv7a+953r+7fV9BkvN/qvUwiiT/Apa1n1FoBrZ4
JsSy3z/SIF09n5ck+SVSMnZYzC6i+PIuZ7WrqcfsNa9J02FEMtb8O9AxxxSl
mm189J28JCadLJXUlviTOR+7UWx01ynwqMvdSPBsu6kxTKV71Wn/LZ0ONaUO
LaAkoQpMFC4i8OiDwrDoWvQn3Im6NsURe8v9X0A1JG/Y/15ENgTejJM5yWUc
syGacvAoOLZYziCyc3D4DODxk10/tb1aWJ/5Ne+hogF2dye5PUSHFIO+KSYt
ZZ6zmj2i8e93pWNjoU20vry1fepGdLZUaxL0PP/xfhd5MrxjHSajcdFWE/iu
CQJd8vFQM71CtD9EL1dXX10+mm8JCfa5cYrDK0uwdQzqu9kw6jwLyY7eI4ei
A+ec+zmv408zNG9OJRfp59VAS+wnYqrAWBRaKWruS3n/rRESBUuL08BcRJDd
4KL1vbSyEgp+tCzGwZm0H7SmqeHJXDkCjB/bFHnVIB9PerleEfeJJoiuwNXF
+8zV4BGIkKa/QBmyFpXjFn5mIIKEVvGQQkC2zCq+Yv6xnlgq5tsEXYhk6a9p
f5IvAeJzWK7zSS6hJyKZTBN1APXCp5QC0kzy9ZK2T4TpX+pJzXytIN6T1vlJ
o601o6D6mY4EtcDUfW1Sx+jzCmbmtNm2NrB3IYqNqdYGBQ1Rz0EZEXpUKRq1
+E+QfkAzDRUs9kz0aBBCTnUwDHvMoD/BsUE+EWugBv5qdLhef3C5YtFzeC6X
u3cvEnp+FrIYfCZ209L+Wr7Gzsy8wkwEX7g1GJsxiez8pxkTlGwxE4OEgTDJ
GTBYPdPbjtw+tPHc/6zqwQMMERocsMg4uV+7zWnuKfZkiSrkv7tM4OG9/8zK
NcviHc0hEkQYJ2JEVupTln/G3It68V8SHCPIyJuATpzjd9sxEE1wDGkTtTUE
nL11kUHY3jMJPbysCz2Rog26KOqqUgP5xA9wdF530rerC65rtV+iE9/ITPAK
V410sX9ieVKykqegqZs3ICl82KpSm3ArGpLZ3Hl35ddd014YhOncSlG2c7VN
ppIPw5r3pllpUWmN6ax1X25yOQh8nf5YbIosBg5X6OZes8oV7BWbD+wwlTHO
awIL+E4QQipGj+h+J+ycswjrEqzeADXALSkPpi0feQEDvHid+MQxcuc1/nId
Oacuz9OTqo95X43KuSKQAKPBi42m93LE/hpzrq/1R9pw81l0LEFoooUipRVY
o+AW+OABYfVx2zgqwfmVN2r9CC/+QMYzYMwt199QyHiAkOYJLpotPUjd0p+w
EQQ9sLloKU88hCGn/3IlTodmj7x1GovOU8s9dI0XxF7oKMmD99/MUq1QgZel
tw1//TSzHxGLq12wH3Q20I0uzn1gUIT3pMPHliU8Xd6A4/sUrRb9FbMPyqcZ
ljxOc+lnhTNVGbBUAWSBlp3XrGNoBjR9PFzbJYSxy8S1CQYByOj9Tetj3JMp
zH2s1pQDworqJvZes+VP3mJCHtzYTBvN6xlPDdxTm4Wew6zb3ilhFrvNxsB3
EQxRzwh7NBkW/B5LkdkP7FkL9ifjG8jORSPwqItZ/6wAbXpg4P6GQ5MoGtS3
4oUkyigTzi0ntSLrpOUqU6uu/7PVVdYPkXl95YhsMIWPEf/p6mtkGMNo0kgn
kjqFMFkA363W8kNjnNHnGxfwzBElhQN41B0BjmuTS9B+gMkjaQEIRApJV1dZ
8sYRcehlQLbpRV/pwvEZ0Rlz5b7qZ+rnRXvG/jIh5ra1KTvNad+WDBkU4iVd
4aY0jw+tXqhAm9WRHUN3uJL6zmCWN0UE5vFQUj74xgPfxfHRQCEMweVjOR9h
fbpUYLegx0fjGR+TgjV43IFJ2zu5Xrb/okAwSDGB5b8uzlCK2QzClZ3deu7N
/LSRIJBPrVgXCsQzYedwgSMyKkWUh5pe6PqghYlyS2e3nJDiuAn58Ka8Zzpp
7bH0h61aao8KQF80xt37t8wEvy9xzw+ZJ79TbtTs9s17S5skuJ1kSZKeqzbr
f/hqEjdTZKTum8u3D5qmoDSxw+HagRaYlyIBXodJaS8h1tGSG3Snv4VnHxMF
g9MLCoOC7+f+QvpwEyy34SV6+iQoYgC1er/68f0bLMPnUjhJBdDoWGmTVecz
glZwc5Ucdz83OkLkCVC5ER6zL85lJZUj+VqtqIBKJvyzHsolEAH1mult6Av4
AO/1SJgZHMdptSth0ecWX52xFJmgHdj/iWv6JGl2DS8yTwq/qTW9240jR/he
KQKYNYyhhPg7dkvQJv6tGxdYsjKOG1jQPmg5ni6Ko7BOSssmVgf2Kn8lSymw
xiAEguuVpgfYKAwD0i/1zQkZEN3N7OrVx3/5ZmFoaXzGgaYNNwYBo4XvV0dv
HjNR/DHKQBEm4k9DELZhfDUbAv2u27tp4QNmGgNIv4Mbakra5+2pwuv5vMXH
4p8LpLynrGzZNjK8m0MPsLShWB8A2hpOWar554ancD3MKF3eF9ZMAvh7JVjQ
xVCBMd8khM01MhqcesHPFOIyuAluDz/oRlpNkC1gLVdA3YoT8/wMY4dicvkK
JHyRirIElvAkQKPecYzCd9kbOv3FCfZqu8R6fx4M0Dzk6NcJrFfmBrgNw/2H
J3g3GWye0HXh5LmfQ/Nwc1iviNt2q1R0cD/zekhQZtmLSlNLcK69mtkS9UPI
R+diMDioJvBoHAH2jDSjVM9RNkjpKm0OGfTj4NPYn8DzxC5y7qf0ugdYzXr/
S/hivg/1yPHUYw0YLbfZCiNzJ+XecbV8XCrSpuvufJXsR+FjJTR+9c+cpMbR
7foPo8hc+Cf5kT4LETqWZvtdpIqR7WCSaoLIVFi5V2Ntt/ODp26cH6Oddr80
MVMvp9yfR1zuQoNBOiUbndPBHoTYlScvYmJDv1HWXM8gnvLlXyxYsMDvUVTo
JvqIVejfznQ1c/GYp9K9UfXOJIhS6JMfa8CApuQ7I8cbf1D08A6GCNkzozV7
E5WafSvd/MOhoYQL/AJTt0+lPWPOMEZqMcxUDd6Ik2KhsdNZle0E4Ki2Pmp/
7L5N/Av2R02SlMZadSTem5Uze/+Md/Fp5KVYpBc9EW9MGx8upVPS9wCFu/Dr
ST+bxtHR4PNMSiJ6wLaA0d2CSTpm0Ub6vrXW5hHFDAD+ce17ODVAbxyU8SaA
CHYdZZMNtKwDyX2QSqyJO5iwEb8FxAVbOtsvdzn33Of18VkHKTjZ+fYw494c
fPDIBK6fb+XGIv0v7ogbLr5nsiNVxCDEaljAZNgVciWU7oxzEVzI1IP6IXbe
vYdmym1eDwUZeTZFsvCLJiFUSLilD3A96+uSB+sd7jPnWdYMu2EzEkrRwwAf
KO7KuyvMe9d8vJqgup/WkJy1nu+cMXQuFGcdr6dtnupTqtwnyGZ5JRGOtELs
A7YyRWt2+aNLBhj1pFf8IlF7gnVAJ41avN73p1l0MJx7Pwug3H+EWW/70lra
ZwyWAuv/J8ZQM8+1AWFrFmd68jRqQ7U6EPxfF9hIzSZFlJmaiW/wcmdnE4UK
hJSZnjxkFKvzSseqFwosHGoe1SKApA2GDYS2iLpvsK+F3f3QrJlrK4NdYwxD
bzGhYsNw38qOZbCXdg+58wLs0bJmjy+7LSuZQoDqmhUuzlSW8z80JSW3NcEA
/we1XAeOH0rLHzJGFA9uWmiVNdb4bThepT5KZy6MhXi2jjZbtsfDoNkzVpkn
Np4WnLwEAZVodSLQWWvC2WH5iHepWa3pI69VN6vTWbKiWAncUfWq34tmdAKJ
7NYJJ28R+P/AaajflreUyRTabCuGdFUGxQhFpo1hEVS2qVrYpLS2br1TrGeM
06WGy1ftsSoRlQIu577ncUFoUFcSufxuE94nZoa38lcAS5THt0Zg8OzFbyPt
DcbNTRdIYXzzW1Gwrx3huKqo0dn4xBTA8pro2/PXMNxN3sapgHvAB/W1OrP2
Z7aK7/Z/Jdn1zlAM/3p8MvFsry9p0SI4UtUvYBdtdfmWvCq//6tzt+SRWKKR
Tow1+1CeCjzAYGkV5CdcXs6vMvf3wWv7v2r4RqTySsDxrqMAk03fmrPm7bC2
nesU0QEiHEEF4r7VwO+ygGLRWE+MEPTCPoQJ9hSpVsS4GYAq4C6GwMRB2OCF
/3DFm2zCZokmICLli3JLvKSasTUHSWqlHBrriu77em3S65d+5SPMXxEKMk5c
LPC5dYW7/ChYGyzhncrmFlDx8uJzWlzt2cvmC2qhYE+DuQZT2Psx+lx5VipD
N0+JDvYfFfSsCQtXK3bqpsj91sILwhxSPb/qe9H1MVRljjJc3icSh+PEv9VT
sP0VOPc+3TzdUqT3ROBPthagsfOsPot6CcOhS9ZP62EQLLzfHHLXNDrWLt8u
lCwpDC9RYrkqvkJU5rWbH1QzAZMxWhd5SSlqsuGCUUv7GMoDI3gSwKJoTcU5
5Brq3CU3fK40XFsafGC2Qx6FI0069dSkn8MqhDQE0O4wzwyBRWjy72S7o8LO
ZuF4a+ivrwXdB+9GQwMwnOIZRVBiUBK3dKUXU+nVPOY3bXuruDDkD69egKcc
yfA0uK6ejsZd0iE9XHD3ZI7lQwtb+ocJtMfG7syrlZrro2UGD+JmRot21mY4
kXPr7aB3yhA8RQ9sSaE15Yjco0p9tTpvugdBpgtlaVJryM92QATvemFD9V6M
ZsVZ++LiDwTZYGlm871BxKitjt2E6tSRatxPjsf0wwjqmpfeYnItNfiZh6hP
8A8p1+kzOJVFnxX9QAXqMA98MXTIV+btP9eCYBQjFPBpKMBDKOHoHCXrPqVr
R1EQrDjeWRcI5xVKFLa/IcUvQenIE3fTSiYnjigMoR1tGwyk/bs/B3H5S2YC
4ivxcjSEOgiRiflgwHcgPC/HHCE34xh8NPmOyput8M7FqygtjnglUnQS2l7c
2HBy0YPaDC8ASAzhQzJADzqFqZy7LenY1mntKeRiL6aKDfuaQdSnDVb2H569
pqxB8OTU1K1NfeRUMRIXh44JTJNCAYCrhkLPGb5DEXWg0t8ZCHqwSnHZI+4X
IF5II9ZpRerVI3JtLyf3ZaliXqPVC48iyxlWwr0vZf7gnQtUkTfsGJhNlSox
P0ewF3B4HmWlWCweoshyFAqy7/MGtiWqaKA3C3FPH+evyyowpAtq4x53wBTV
GyGOKuIrOXLxeY1PeuNS0G0577BwCYxeFZFahLZKqAb65PWSJj7nWe6ti4LZ
u011kE3a1zh8xP4MKtNZDF09UaYlYt8M7HoceChivMSWtTxUBYbhsG1a9V5N
Mk1Rk6HdsAucfsshY7BJEuz54OwePbnv5n8UCicHPyvs7kBnyd1LNm34/7IO
9Vp9dPL3aLd1RdsbVRLsMgpiGBhQXrzVgYP0TdS93J1iE2prZfGdbODNmBd6
czF/13PsaKlywQevRsKfBRmT45JQPpxVEpxaaoUH9OMYxQcmjMOoBjrXXWfV
0xQA3oYg0RREZQAov5O/G3oukPR8GyVSUhAvK/Yb+W46G1tAJ0Bg/zwmUZ9M
kzEwWB8iLoDHfOznvr0i5f7F4CPl3mU7iT6F/OofSbGAlnoHZ6yGiQx4L+S/
qKaTUNSPPy0X/FzO106TBm23P8wsXjDu2Ej7GU6aRSTspHB7c6wYEDE9mEYG
GVFsvHjAhZqTIVNXz2IFnphcO43wLtVI592Ge+5jG5WHvBmJRIx8/0lNv4Bc
0VZ3xbNIT/UGIwDkmNmZS9P4suo0vT3Ynzj7eMot7aiqerv8otYYvy+GJ9iY
gdMur1tPTeU8I+gbnvvLyaXJLx5iI5akIW3bGx9M1Q6N2Z8PbOBUexwbOyXi
xXr3f13Ne+fuW/4WoyOtPzaV+zuSTa6N64TNKr7ojX9oZGWJm2jTvIHtznc5
YFWcDRcAa3ZHyomg3Mr3UdRtFkMM1heuNTucfpogsc0+R7ptXDkGLPxA+31C
bVPijt+pJb+/nI9wp3Q9LRjga8iA0H/mxxs6yPmSszaR4h3zgU3SLz+qqkjU
fJreBS8f/cYHElzDHMrP64cOSGgu1UXl0ExTPTQbwjR3dbuqnM9CrzYV4gLK
QSHV+xGppDV5jlNbxaWfnaRN6YXZiJZPJmsgPSKvbEEcDfRj/BUWsBBMwUo4
FuTX3zfi7Nnx0d6emh+fGF1bEB8ICLVC9r5jcHgRv2d/flBS3uY4KUO54NrO
qKUwRkzZDttxulUOAhsGamXD4vqQo0JKaxeMRNlr6LFDlbdK/FcEpDwkms3O
NWNbZpN7x2XKKGtstYyor/AIELnWdBPkzGw7Q/68XoINNdAwWtrrmVxLZVLI
7UmBCxyImhgJr4NfpaXcFvGNGvhilzMCoOX4WS/2BJMCk0R2rfTEIvGymR0K
XS1DyCY2pg4ACsRqfhFFyoVhClvPNZOcNZI21YOrC69Ec795pUfUXwc5qA3y
mZuyrVWfgebZJlfhx5Zp5HOmjFkv2JTqwcu7SRNZSvzlKT3LMfqmbmBFjby3
h9uh2k0/5RQsQpBR+96JiH5dWVGgyQ4UFKh23Jzu566xq8xow+dMJdE5totx
Z5x9onFcqIHUHVcvh5oRrYBeb4h/v/zmOIfH0q0loNfjTwVnFHgcOAYihFoQ
q68sXwwlwglAA0BkOQ66Fcu2MTrTC1QfE4UpIe+w7cROMlMw0G4pBuT5Zuq6
lbskL9DmMidrvci+6IES0OmIoGTNQd8LM3HKV6xgfp6L2wMuFEeKB2WfdXIX
2lZKxqF4POGcgPZUhe7tWIpPr0r/p3ur3XoIb0fWa47aiL5ICcwHN1vOGOGQ
MTH+x0KYSWigYefJv1usTkWtlZK42DrS0nFSQ4CReMCvLNXae8tGi529y8pa
lPdFDsf7z+xa1M3M7iOb3i4DN99C/YOnVnR+T8jHHrExpTbHhsUTUA6wEEcF
noekAEeflrvnJVCF9Vv1tP1KGgkXKkaizpG6EE6JQ+F1iX+8jb2PeaG1e516
C7mVCQ9Wi3vpvplzAu1pPDuFpjA2YU0H0cw0M+7lnDiFFM9SIAnJLPx6/+bh
cy+xX69h59WTp1FaYAchoKOWssv+b2cd+642kWqPZSMWxpAjuf712kNJEY4p
lUsNN4+q2ESgm2SrkKDAnn4hCikbxAgqn5URhf25vrvuSDV1TYosWuBPNvi1
wJN4h1iJ/NhcJPQfgKSHveC2S7dl9belnQNpIPD/hJQHKBNpaN9UhCRlysnX
5vu8xf2DpWuH6kh/g5V4Mni1xesJifmkORAExpo7q8TY1P3ZdWJb8HNPE6DL
TkvdhifXtPhFxE4MIO7WFlFFUDJm0tWgCDBhQtKZF47T5Q9Tq2e2bAwWLZF0
j72wZA7bbRBSEfWHjcs3YZhu5t6DsTLN7pXlVNbQtXpdq5glxPUDnQN555wo
UdzniNaZyh0gBfiG4s+Oep4gsbUfL8a1VsCN2GsD9x79po9/ld5i/x7+/sPp
LHUylppdnkChE1v3Z6cm8QoWNC7vur1U9NYyWEKr2YT76sLuVtcc+RcYGUu/
CVms7cLRV6sQILRW+UUduNRbcLGrRvV4b+jPERV4v81SceJkHgzixj6PoScI
euIjoAioPBlTR8hGzdAIjGlNVhS/uywvSGN4W3fgfw4Y9wtu5sx56TzL3AV6
3O2LxsQD54dYYMVtKEy8TJjrOA7TgtEm3gi0DE+HiuAizzAunh5+MG/v3l1J
tvGhVoOF6ll3pl70F+xSWxCxZ2GPcFmYGjRbC3WA58WVnwh25fSeBI8tnBhm
XM57D9WFPWKUj7qoplg5Iazpd5hkutaEv3N0u9H4FKDr9Ld3CqHgQ+67f3Vg
9SPm6lFGvMhkP4yT85sOqMZUurA9iXxeQ+dEKx0dU1hIkwSbHmJrdCz1UBG5
1qBwJmrUZLvUpZSzrw9DjRQOSD084+VYRZQUgGCZASwH77VmSER65a2jkiGa
tW//w/XvBioiehtrcJdqOC0oxeOLuhhWEVkDM/2oenR6uS/PzcfWvVoaBss4
iYK3TkiVDHu+Y3TWVhvU75+2bWQajDKRffBF695vhJ0D7bImnYdoiEN7/8ML
gDm5ijhzJ9WO35tR5WOC9+J5S2MOImTu5GZI9RH3/GsSE2PGT18ccYO2CZo5
yucRKH25dtqD2INngFgUVS4bRFe/md4zPal7/rF04adDbl6S3g1l+pVBvP59
8IzZhZPIgiEgPh3zexmj5qC1zCabjlmiRW8ttnYntZcY+zEQ8UINDamIhBmk
OOwbzqja+iEZbdPltrRuW9U8HPpamACrZkVrYY5yRBk1J2tl4tDshC0c2uSJ
KddULQlCsgkoxcs+oFuuBWhXPGKRZZz5RVgawTQwtOUDN4Zuar8m1NFui5gt
FS8FLCYZITRODkl8J7xT1pxAnqGt+oiTrw90VjZ0PPjMiL8cMisHNjP400oK
StEy9FV0lpoHjEoVR2w3e+tJrTj1Hxu5X0JdDPceDmb6CI+9UnP29/k4liv5
lGhBW3ocl9KDmSLPi8NzxYMWwlEu0s4wTDs3KJpynd1pmNW+fFFeivp8Ay4p
T0Hq9M6XATnz3K8rGi5J/P7XV4OrircKnBpFZ5fPw/IIX63UTxwody1xJrni
ES+lERfO9tVn4diJHzFKKoxEh1RU6PeWo/ilEB/xhtphV5G11PD03hdrOKwH
2MhGsytkq6mGwlXbmx2mCj66fILQ9vkNb6TxatxtJRPSCAwqsxWTgBFnHgum
iSnbQM7m4M5MhAmnYanr1g2azVLX01mNwwZhDTPEyOZXDTdruJ2Nhoam/xK+
hmVWtX7WUdPZRPRKBmxpA7KTH0TyfSPJgC81JpaiE0h3fUlBZ9EhHjzau9tN
B8TGZpoXOfqAb2H03kR9+RJ5TBwpzVNcXt5FfxZ7hcXgrh5SyUUswKpMNe3P
tJnWVTD9NL6pTlZadOHOq5l81IgyDJl0wJkEyK3Ekf+i/KqSqPZzi0SXIWJE
VGikgBGrFyFhJq/88rr2yABW7Rtxw2yx5+ouHbekKL8VL/F707WhW5rKvW46
lVlI5vgydUGoZxbvueFtL72F82j/fcNwZ7jGBn6rpkTUhsJ1mr6rI6tE1Kk2
HXX2S74AJ/nW7QdSf0z0D9dYTvpNos7pADQkGH+4hQLIyEc10KucBf4IqHuV
XFBSPWhSMD5uVffb2L8GshWE1bj+jLE4MvDMdiNpdJG8uOe0KezS4+nRr3Q2
lhjHi/AtGGSRiboHexDuKqWGeekEKYTgu1GUsa9ThM6UpZ7I7AQuX8Wyvo+M
GaR1x5pXQpHnwHLwlFdNjgcNM7DtQKWigXs2c8Jhk94BBIMto7EMLnDmxG8S
5BKCcG8OkeK52DBWZj2Rv3uSj7MlQxicg/wytORB6Gy2i8sVjvbbUKYV0t7g
nqgY8sqMPCZwP+UuRMkEj+7kGcZPdZKPwz00JGE9Y+qNNng+Q0qhSxgaGtkw
tl2Mk2L10V5cA9bZPr8tGIcznYOyzaRpEcxIDasLIMibqXELjHwty2jLVEth
a8zpPLSxZWkb/SfQmBvsOWKHA8azOxlcvGIN7drw5CqkPDe8JWsDx2T/EUsg
9ibdMVXKBNiSl98IMXJix4/SRM4mJ3L722YPm31ybOtJJKekQGgO2veZWYds
0KFxdihM6JRQSiTo0Qz4VXays8NrqEBfhK4VTtm4Sjkp99pCwNSfADWv6liL
a6mCEyvHkOjNC4NlORp+xkQ0A/rNtktPocoGI/ry9J3SVhOtCgfro864YQ3B
7ePuWUwTuNi07PDSxxIC/T905iHYeUBqrC2Wi/iONHufkiapkjPr+Cg5o0T9
z7WDWlmwezr4h7xVz6h1nvGbxxA+SbPQAxdEjMXACmSKXh/SFY5nOn4vmla2
4HhMk/EiBifXAiWmEeMzbzIqE0Ysl5D8/AVfEdZ8AkXYNJN+ou0O8mAMsS0B
Uv5Bj21tDRuLP6VKuhDECEdNJnS9dyxHZDkKB3Nn3nF9QVvBdHfbi8mk2h7q
0riFcwRoHoJb34UTM5L5RuwVN1Eei3xS868OgAgxuyycXfCfO5Hcyj1hyF5+
BTQJh7Nj58Aj6omwAbu/d30xpAtzuSRDNCAAqRK1Uc38NZLeGAj1WXSbqlLD
3eXlOnZUR1LLRGV1B/LXTMCLGFqWV0byYv8lMAOTCtak60ZT64QFZxxrTcev
VC3EesafL0Vd7w3WJXALT6GYpu3jDjCHYP1mPOCc1CRv5kz3eYGowEroY5aK
lpbD1Pb8WbFCiLctUaopItZQ3B/f6rzWgYjTHSWcDAKlZ0OIgzvdLEGG208t
ICEsvVYtu59RoV0dxI55mOFrUm5QGXm/0RACFLdOjrACCh6OKNJP53YDmPkY
bVcxdKQL7WIbDU6DJtTtaDGqozEimPe/bm8y+iE2WzcZjdrMo86FCUHihVIP
xPufveAHMuLr588Bt64SHTe5mRxB2cBjYOswpXrox407ML+k8HhZkSgC0Acp
kNSozYaAT1uXd3ob+Jj9j7+FjmuEPSWdDRsREx4z/AX/mFINPXCfArD+Otvo
hU4eeL/2/tbYfL2Uq6uLZPBUNdUEaYDH1PR+dr7/qpqeCUdFxrdIVMogjgr2
L1dzeAkdh7AH38f4CJy5XHdk9FljYdlwAgZMVk6E3FzYPqq6mJtLIk6DNFgl
NDlPpWI6y6Leux8Otn5+t/aNBdAaH0dWSQat1mpndM4GvG5C2Wor+kX9rzYH
us0eIUEsZI6IyC2YYoGOMqMSzoixW2L6bTcjzcgtvwxgl98bs9aH2GoF78Wf
gTRyUfYXS/n+JtgsS8+qjmsvSk4l4NhSnl1RYpEFFZsJqzov+jQoW/hwmZlZ
Ymfx+gtVPTaoejuNZA6GJJff0w8/oDdfioiuyOXX1d4ALrIy51pGvGSFMyPZ
Jut7qhBj7uXddUAcp1B2QJlKeJeF+DknYebQQ3UKwOTLQRuhTKnBepoXQ3gQ
ZRqddpNV41lETGh3smN9RzBH/kqXqwQikO5PGG/RgaxgiF99nsbq0BeHvc7g
O6iYd5igmzBdBPAD4r+RYqLwWCEJvhr922NELgfy38BAUuhgkqNpaFvu/e89
woXLpiqcN76Jybkfz+Bzm9XcVRyWrNeOHMH4fDasXeaHEcVAowuBZJym7LoH
ieJ4RRuFqfWXriVSt3GTO48AsGhbkIjdvMEJpcSafY1qGh5c0X/GJ5BQpaF+
wnZkGyFgIJA6h5lZvrq6mhNtd4RvAdohDvEtnhGtJv5By7u9VEvIDiRzkLSw
qeyNUu8aSH4q8LFT7G0tgtKUYFxhXdskHd6CGNgSbv/SJRQXCVNNZ26A8tmV
gRZU2N9EiXGISy9w+m1J+IuR61kvcJKwWQ0V/mShQm99ZofD4ngSbLMJ9f9r
JA71+T9TtxKTb9pKTL0m57hgHTyGwFtrUtIsnpqNR1uTJuj1NgN75hfgmnTc
BhRM2RuESNb0NNfZoQEV739yaW0XD6RNOdyAAXHKl2xBEwzhA4bkjJv7wgwl
MhsyoZJTDXWh4dcbK3dj6VwOGwG4vLaCDZ6tur47v+ihCbwQaUAuYwG7vPym
GbEY29FgQy8C/I52hSWxKWUUp16eQKRwyIaIovcfhJsqWGXt7DOdi4D4W9Ja
fnd2BfN+RL1wD1OMpr6WCsoGObUKUIx/hj1fSCA522EaW5wQxSk+n89h0avo
33RmkCQa4lVn4OHabHKyBJHjAmaK8iYtapFxVR5CUKE4XJS1Dz3c04fe0SI1
bCmhJFgyLkRUk16V55l3HgeVffKRzCKNGK5z8GAeRxudl93YgLf7/9OfMR+m
53Z72SYM3c6tUJ3oJnrbYh8054YkyIGtxFkIlz1vvDRuvEFNXvDFxJOiLzaq
ugzCVgvquN+itzNo0bQKLPXTAzUYt3iAO43wYlcwuvuzvoBqjEC79APOM0Zv
Ffyqp3PlQMECSOA3u4SkIYGYsrHT8pFOsy69XNHPrfAG36tb2R47Y5b8nbpW
9IxLRhsAtgI0JDbbQRnzRhlaXhs8nKGdiOlFLFEyKAdZxhjBf9ZZRLkaptng
yZuNfIWsmiXqF2PPSi5cd7c7eINMGp30axKaxxDxY3we6cN8WURrIPqU829W
d8dKpWkNr3UhOq0srBFLCGuyd+hC18mOibRdrtCVfvvbV/Ndix/9DfJjov6g
O8hKL+ejykqBT13xXxu75x0J7uQXPtL07+gjuCBzDBfZrskr22ICfMQ3X9Gg
oAegbqzamSubnVXgctgwXsIOP+QmAus/voVJ/wSSGdVB0OY+WUrROhSPf61q
6cnYncyxNKfQzV29ygs7pJQnnJgYIhxYflAcULT92lWdnBQIv7bs7X7/wpg/
d6htX9Wq8ZyWuBG1/bXWvI5jOZh8AZz+YCDft8m6u8UEhxHSOG5N/kG0xhK8
Z0Yuko8CD5PlKdX9Ftn5yBO4Cgj5fdzeSS0Dc8zOM8+Nbu+13jl9PqiDvjbn
lzc2PVZki0z+aSWW0wf09gABGvgu4wCXrBouHivzNdFyjp2/2bSxEqYv9wCW
GgUe8N7OW748ljrOcdtMOKzmw8JL9Aja46LX1RB0vXzQLP/ytss+ciKR1b7n
kkcFjWziRtez1bX4Wy4Dg+fIeF0Soie/6peKh+QU0Md716W5OMy9yvoGhUcb
EEB0K58Bunrb+gytvQfkqoqPZKSOaDTyKMufe69rBMtHd4hCydGTzi/aoUuO
Cj+cZ8FR+mWScpN7b102x7CI2LbSlrwVgukmcinoTVjy0hFrwh8QsoHvKDh7
J5R9+7i5/jPa8p+z87l3RljgGkWNcwkxcTXWA5Um75kgQTNNZrjiuoiLC7T1
GEAqg0AwrFVWd5goZyTgSY/VEAwBVV2lZgrwJJ48rbHLxYMa7VYY70bmUBhu
SFpJBmreiiklg+5fE9a9qGAQmA+wRsg/BexGVQ9HSTqeyZy7RuKOqx0pvAp8
gEg6vnAmjRtQlJuK4NSm/WHYG3JiYg3AQxKyw452VgMQUQO2sV/X2OGSyPaJ
EwCu6wY8D3dcfkVJBRTZi86sQR0QGyEmBqAEwI4eE8lyZiqMG8LD3PQvyCeU
grg6FB6lwLF4bqeTZI4o0BuTYGcTK15nZr3uktTQO01IqDyJfrU6PEXZgrdQ
taGrct9nfYBZzsvCAcqFD7xOqK7nDcng/jQpFwHyW0r/T4hGrDwOii7JqmPo
F9aIx/z103xl+RXKFmjSoF7m/+KKF41CLOcbFPPuQ1COJn5ao9z4qFDHdXRv
CqxeLPdYg+U4p0s99MkG0EMgTGUwokZLOf3FwhYB216qkpzO4yX/ASbFHpjx
j4h7cV+XTV2d/pn9ts5JDeR1MShHKuQxLxheabzfK1D6EgB3C0UtWP6dmIVo
W3rlPdSFo70khfD1f3H9jnNZK4hAfGh4GiBNpRCa8AzKukVH2ZBjYrb3GqRL
6g6S8aIX6pZrMacNZWaPlBUPFHAe2LT1xQ6xIxj3JDvPY88rJAgPRvstHvwj
iIInSYZOrycHkJSGnoddPqKd3t+g19/0V+ZguyCHtJ0vaktti5DKpgekq1PZ
a+iSXmz4Gbmu8878Hwhl9EK+sXfuTvVgBdEzp2FMxh7gaAUJi5TsYoq3926E
it4gViadunwk8PynT/8xqQ8bDj1dOi7lhnZHQVnDUTFOQMO8LFhxIHdvTL7P
K4qd2MhL+wSxiTA9aXuhO5rksbGOL4JnpWT+dHD7NSto9sGR3PtwryNw+Q9q
hzpcBhs5J6u1ydxoOrRz1aF7SXnn8poOQQaOg5h05RAwVM7xGcSlf5WyM5C+
4D+dfl9SBqTSv/MobRmMLWxMhdgaCKuy88JWONytIP2+qU+WoI5SmM4fj5v0
EG8TpC4DxgDZTexNFBo8HoZ+uWOGIn05mkSUa86rJkBZv+PR+0JgNB3i4/I4
VH64GRZaQYjm5d1TI+Bxr1jkyq3+PL/P61dQIdiWEK9xr2RWzke/LqMaJoVq
zxW0YezUhm/78HIO2UmTW4vigpVAO8WFNFsOMrbTXSRgSUhAqA6aNTErkncG
mtlOY7dYV0l+PwEISUhdcyR+8ID7DvRoRdKmNdNvQOBJiMtt9lw3B4oJhoQM
67oC6BHdOdcki4CBtg7s40uM0u3LUiXVpSlVJxrO2csiMiXpunW47+nQ6fde
Hg6fCi9z00FcvAp7ViFF5GugRE7h0sUOKcyV98aPfXwZWShMsCuyIhCw8ui0
d9j2L6QPc+hzMF1YNz683uDIDjYQPXXeT4Dwyeq/nl9bZNifX3jfzTaSkgco
eSJ2nhoHQzUGwvCrLCZ/Pec03itbXjrv7bzVI015kcQGSoP0j9YAlVsgigr7
QQjBFcaQtZE7Pry/u/OCSVJLCRUWRc/ezYt47UNd2XleuGvD6NE8TsZktd9c
zuO/Ou/SRE6rRjFkqUvtuvO3zuy3EotChVxlxAjXFYJ+9hU3QMo9sN4bawrq
1tPsAd9jDHxmWV7GAoLLmFoewvCENoNyd9R+qiwpTLOF194y4ymKe6vnKt6O
fkGRm68PHRXz9HksMG2zmsPYt8FNUm8c2E/WTTyeXiFBPUNMHSao7ePtoDMP
59gkuNDcoRSyBm+pym+jUTGPMf/wBS7xsqi/kJeiOjIETKmvTVWVNfiMbccj
PoANv5nNsl0nrs6msn2v8F5uEia44E1jeFBv3CCOhRjD2giIuXyOw9R1Obxw
cx4uefIkr6TG8DMdLh1t/1t7eRRzKrn/Ad0m6KPzbc+QqYysPoNsO9T6tQ43
y/RHLwe7u6Nz96i2QQgjVTa3xbsVJgW3p2euhNX9oPU6kglLZcIinFU/0Z/u
b9zlYxjeJBX9RASYxLMrWmLJt0FRZYpcu+xz28NdtE5uPmaa8MtWqNqeqU/f
z0lO4tEVAio9D7aITDpDBdhSVxYQ3kUh7btfNgAceAisjbyWUaxRugUyZwjq
/0ErQqB1zBx1kPBYoj1ULGnMa0Q4C8y2QDfJIw09+46aQ7dKb0ggn7r+h9W5
tmL3hlS79rN+gAxZut9juem60ehkrpc9auMpyRHR2Bj23W0TQddYdncOfVnU
hAMGjIIYymVvTRHMxZx6WAQV0yJ0T9IrI3639WBNq7zVyFQQ8IWzog9xjxrn
8lRaGlkrWNg9XwBulHJP+8vBbx+kgA1QUZRviyygRE3EWFB393FaGZJT4moM
RD05FQ8O2lEF2vbbQnsYxOb+Avebidqkef781JChujnB2MgUFfLNNJNc4FY0
CkDNPE9xmrKR+ataz2ar5pKC/qu+5/0aJPqPunp2UAIOtvA02Bl04STUBPQp
w+f5hw1Xw4T4nzYgCqxm9nesCsAVZ2bwVIL9DYjgqA2lyIPihJQzJDfQtckL
qE7jR6eOlHIMwNsc5YepphoGagmTR1uekZkCYRpoMoZx1/DMam31XZI8tyzA
Mboa3qGlzC+JGF2kKy/u2i7C+GCiumOZE+gqvWDaHixNPjXzpapYZdCe7AEd
jNH55eKSP5iP6N4tPIdQwRkbCRwvQ8hngo6LVZouxcQ0iS96Gzk9vKzlZ39L
ezM7NdrBQEg/g1NJ6eT/iqj3pu8CJmcPVomBqt7NYCXyrpLv6NejlDjvrWGJ
XC8pQt4sGbD3MWBvEFPR8yG8Zp5IJggf9MaH4f6H6VtRzgqD/DIRyi+yB5Lx
JDY7ZbuwBhzkfT+fvCnGmlVsRA7OsIgQn7drS95OFimVdxu4fEi4c0Yhiib8
hk71Aoip4iNa1YXEf0WhmIGv6cDAhn//jNYuz1AZEMKWviTX3QGTjYbLCAcm
+MNOpzNXveAWT7v+/t9CdQJ7hL2koQTdy8wzqNka4JrPJQvj1piLPGMWsf4H
NwMKUc/mYX8sV7RxJvqzNh41PDJYcRHtNRNnelzjQi1ZsdVn9uJHrHoycOiq
VGWirJBoYF/AAfSa3BHupIlBLlFCK1uZq1tCCHPzw3JF3R5cbyGgo/U/lL6s
69B0vpgrbgHppIIwrRJUXRNtAHKTgMyF1mHA36/wDvvISI0J/vQF29a/qMTE
liQ8dvuc7GP9o5EbPozKMK5k6Jhzsj4MmYtr9XDn4KtYkCW/FkEuH6q3+uYG
dSQcN1wNC6ydTUNOlBsiM7p96n7PzWA28TnUWpwS9/UyRTQP1P9EwN2URey2
2HeKoFKXxnHPlNxiLko5jsXKmuiv43IkYn18h7KFw3045z8ow6PZAlu+kj8I
SuF7zmMJnRRpBHgxv8UPVr08xXHiojIR259ugkx9BwsKTtlc65cmh2aEOqcF
2Qx6cof92WPOIZyCcaRKXRfADKXrrCAZF2h5N0jH1xaznL6nlWT6dW06gcOl
VljNF8q1K6SixW36TxAjHne/7hBH2TjLpS9tGsau+qxJ18+AnKKsdTrwwpgO
nUg9aUTdfY5zU0W+VX3tCRv7AmXK3iJ6V1roGyHNid1uJrrGZ5I1QDWawCVb
dVVPpiq7PLy9QMudpg4G78g26w4ZVTFWk/9b1X+mzhutZQl706FPLIuHsThF
Nsgu51M74UG9tShRCvM0Vv0uxNH23BpDSTFF1AgtrZ+MTVhMKiBJihSYCCdN
Xdu/hIaNXRJGxkAht1Xq6UUjFz670RIwYXGPd1M26Ig5Yfr5z+fXH5GVgIlC
KKJMfnE2WCJGsnzEYEIyw9w39zFezTqR8S/nprIUKq17u6WWshuVPRRbBsbJ
+lxc5yCJYfCkI+cC522cp6u9QTjwEbAhxgs4gGSuojmQ59cbPnnaLCXuynxA
bM7CnpisgQT3mlNxXZ+VSrrTeiTXNvx8F7RVxirNg3QKKzoQX+kP4/LSbuE1
yYFhzYNkoK3VuuL/aWnE2wOkLkxovDoJJ0NasdjYbEvriT8tTN/oTojv6Ft2
wtT7YU/5lkhstUw3EyfTjxXJRn/5+AqHqvEE/2YqWtNMGNclwRApQmfNL5d6
W6DB45YuY3/AR1wbleh68mj1G/XxNWOLP7SePNhxRAi0370NeeyTBt3tUmoa
4gRkL0c76+rYXjtPt61bwhUiFNiTs60VT6Ey3pA6PBdAOAwk2/HpoRDM9Hgs
bBpIr9q3gkIdfGS0J+Q5cyHRpZm9bre+Yradf1Q2qL1ABYR4UCee+tvLP1ZL
9k5u1XMHG7NiEa0oSGkejQKm/oBJxupGQynILWNUoFZBv112VJHclGSjsY4g
6UsC6OuyBybjx5T3kSAExCtsXCaU6SDkTJhaKz8jRISfVV4e5AVvsNUO9n4b
eze5nDqY4C6kibh9a1VUv54eSjKWi9TC3K1WlqHJtqd1FOrjG1CVeRoRRBy2
xBJY6mwSal8+uIS0C7CAUw++z77xA+SwbL/+3ejuPsXtcFvNZoD+fHzWW0Ym
JTfYt1YUilia6xrnct/w2KxjPj+ii9Lbv8hCcYCHQd03cWMbhs2TaKcXgazn
uu/ZUsAk38TVPsZXQ3d1zKI0kY77U5mTqdMW9TiQNXdkDThQ0LIivWkr6Bza
tOEWSKtBvpWCyDwfHBe+SiFEtwug4j0Tlx67+i2Zu8vsA2qdC3JVF1vufUd1
TwxAF1gMT8SY8im02wetH5hF48Acj2+fsT2IfKhTPeGHHliyVABuscbSHtXN
34ZILp2o9e8tUt0S3BHgUs7ixg+rBe7AC7DGfq66jDn/PpIe9LJ3lHxfydr7
8oxOGAwNSx31JUSRAH9X4qDBMVPnH65L4A0zobjHsLZXTp0BdBlnz6XMYCdY
mLOfGErsURh+b3qFpE8ntKbNE/e2/9gn7NlV6dTf1gfbqcyWnS6YljF2O+FO
JnBauDRV5+7CLjLNu+UQ35zGt9pLa81agjongSSHEE2TMsQFWmXcOjBl/+PB
TB49UKQRdJisGMRTYpJtWHCd3bAUPe6DgeK6oN+9FVyl8NnKftOxOvLiUhc1
LhiBmrvFEOlfr6Cegc5lhY++eEFK3pd8mqRKCy9CvZ+4k44Vu9uNVdiPhHjz
sPLJx0XiSkdcxKenT6A7sgGzNflVLQgM4vet/1uvwhHvmdnY5Xgge57m2tms
rqg79/JzJJrv9RR70fgBblekgZuYqNfJU7JQSf0gr3cz+V4Ojetlb4fEhJPG
si2rMM71F31ZDzdhAX+ZvbzM8UQoO0NYWphf4VQyCIJ46ZV+S90e5jhn/rzm
cFjVIdPqKEt32DpOADak0tvfhw7R6HtIcYmfJDi0V51Hm/FHYQ3iKgA35NuC
5NCHuk+6PrHSprgqwBaQljDF/aSopyIKDjSC7Uh0+sEykAV+Lr1tPIt8C2lY
WOef0OmkNsExtM7ZjcuNAdRk02XPr4XKNJo6zGLeuUU5H+FLPgPMbf0/rpKt
VglBSWmvhPxLw0gsNFxGHK3OoG/yahQAzDaqchfTC6Xj/wuJmVcMhX6BKJYK
fR6k+sTVEu6WkO/PByQq+yLmOTqN+jCYXru6N97PDP3a4IzndvMVSF+YA1C4
o5YSnMdH+5gTOYQ0ugQkIlxanYQoG9J/4OMRbzG+RT+TH6eHkblzmecjj8ft
EQjqXiG8eJolzroR8J9D54UiiReadMOkAmo5yMy5L37sNR4HupnffU/3N0NJ
Fe/XE3G8csN0dgRVGjD1FGWj/Qnq8b0tY9OcMx6kf5THAmTjiZ5vWkkZRwet
B+tdXC184ZQrCNZ/N9QkGzFgxBQl9KkojeJRtZvvgpKAsQ7ZrJ4OQkGuE6VX
BJ+g2tfojMU6MeTvTaY/fG797z2TueeLy8OiVO73u2NRXaCRh4xah6fzXier
Z6732mykACFboNXIAu3Yz72AT+rRp/wOUQddpdWl6kV3knyzTHa8+NCJ37gh
5pGKJG6IjvEQMbPciAiXF975Vq5ba0BkS4TGQ+y82KiC8MwrzSsgmSN1veUw
qxj9ctx3KmycWLijZ50bywtv9v/MsA6r6HaaNqLGgY8UIHNy8LHLm3GjhVtt
urVUJ4B95/WV167NgfT0Lc9xOxndGMK1GWiQo5WouQOQbcS7ggTGI/GgIRcK
y2HXYkoYb/DQcUDeGgUs6nvPsTzqToEaHdUeYa4k9UeNWaAvoWuvYJugnARm
+38/QtOkQNPYE2bn3aswpd2hSYFQ4Q7pDWILKa3DHEioXYHWsUJ6Vl7UuSuO
ZKJ+AGEr2bmGVbEBH1kRlPV5CapGYQwdWtj4+omAqTauAWyUDRO9ac1dSfW+
EHlgFCxKJ6SNXJE+hTjLNSGwKduXPSE6P9S8xZ8IAwQXgHpsENnHYsV2gblU
AOZiiynnItPcQJI0lwvN+y2omkG8y3uA0690TMI242yD9bLyzqNQa5K56008
kevYWYiIR7UMO1f9KQ8r/XY36dUMzyPrK6+qXkHdsscFwJ9LsCOuBOTNPV7F
ieAxB/WiQeigAp+PNyIGpF5fGHnN7/FezUs+hZtBCRQTaXxndtaGvC39CDAS
/lCJLcEg/fQVFvxLUbFNUcwK5mFEUkwd9Y7sTAjMOwwbLq/IOR2knySXp3jL
y+nNuMp/YEitA2DtPdVsf5N0zNmbJlKb+jqwig1N7snlW1wh+o36iGE21iV5
mXcVH8h91y6oCI9U/1vhwuby/gEwui1iVClnH9H5PaGeSd+5qAI52qCv0HBL
LasjcxGmE8MXsSWcNwlTG+xM6QAghpIi8eKKd5SRFdkkrSCrrHJK3+V2JhXg
g0o5sjOdKeu3hSY3TUHC433aSinvJYtHMN9fowLly/+1TERgUsvDXkAAk6hf
wRcLuMrAzdenSYa6QjdVkxn3mVkCgYzRJiGTEVDQSQyv+t5f0A4qD60rLLcq
GPtAhF5Bt8huv8iO+sSDmW0muRQquNLHI8uDXOxzbaObfy8/ENHEfgc2Q5Vr
WCWTC0RiZPWeICYu4UYuxwfw3CP9BX8r6SPIQgpFwbQA9MJ7P5ASdnDelSMy
wOJYDPiSpLRFJC7XTrhqlAvBLHLXY4kT7cdRJtIfYffJZcvvgg1HcMfduV09
jalGhVZ+JrqFM+dey4fh63LVqeMpXVQO/c8/V8j+VppmsrmVHy4Jj/3uOGwz
f7oytuWto4A4IFecGxMR9b/rxSIj8/zHZ7LMJv56xokKyrtb3IlIeLm4x1O0
7eTKjIal5ZLZS69lZHndVj52XD1vP8sWRPlPzaGx1CT7HtysvBYbSu+g/cvf
oKN4+dAKGumBdKy2c0vbDBgoGtxVoDtLe/5QrJWn6jcEwEnUU4GN9uwLwwhB
LJiqEj6wlovCnu9UGjnJcbRFn11uy46jgQD2lYlHyiosj78F0+o1ot5JuFMB
4ZIAZBqTuTtGWFVTvzdRyJvmzwvhiHgvNDNpcJKMgBrk8tuzaq09ly238/uD
kvPwAMKCIQht6UPiZV0wpAio/WCUiPJy5OPE7J7g4U+RNYRusozV2ZbuLJId
MIavZpn35sKrfg2rT97EQ8yBjzTc519evRqQwHDneECE1gjbArzCP135hd2h
jzRO8FRh1gCADqCP+/8PXz1a0L6p61XfbT6g3mfagd/o9jUNJH3anNhIihiq
9A83khl+3BddQ5a+iJ16Kniv6+xa8nrOEnQ76nwEuuK44v+9h4l+DC72HafN
93Im5NOZeyscq6fMfPRBfcnCvgyOlVx2AHqfkZpGQjXjuKkvYO71XMvNPiXc
nG9RNcV9klRpWcQJl1CvXo4kFfQiB635uk5oZ69RpmB8j/xRmm1XePOq5K4y
qYignJ0d4VYe7QBObDt4znuh6oVSGylIDR2NdFq1TdybS+fk2L7/L5JwKILn
g4ubpvzBVh7N0zBf3V5cjKbLNU/hJs+sN8yA9g340FkR4mzAfbHZTwms9diG
Rr5MATMhN2Io2eFIaCqmvud6UBYVAH56BQujQVo4nt3LX+M6moCIYa4+j44b
4EeScDel/tss/Ti2eKPRssLN2OIjST6uVBylIjTJltJI7Kp1hMO9WwjGl6lT
oYKTYr6qkgdjYZ8XD90TP+7yfuoKqGNv6/MlikkvX0T2zH/s7QG1vA2ASuvo
86a0VZRrJ570iLhaAb6DpyyDK+xosGU7iWpHbqO8Y6I3SL/pmk7riI7oA3cF
giToHcUjtqF640vRm4uXQX3ZvSzrq7G4ROyFfV3zORPqWG98gIllJnkamlaV
WTw8EdN3tIL3np7F9mnzyu2rM3qf7yNMwD4mdqtDU0uVH/LmAWnf5nJCmqzR
xYJEI4ikvbN4dLG7UDTxb2StGBpmc+b1LeVXzBfB6BBgTXY9F0eL4Fq9ZVVA
gO/4SG4x7XgVdz9GU5FO5dwjaKN5A4kat0iSRNEBTGK96CGOGZyZJUDCtdPJ
DkNvY0LYn+CQSjK2xOsNteXuCycP6uAe+MLcTPKU0maIVUzv/1dLkwPqFlsX
vgEHDnSyx16aaUI88VIEHGEP1pCKGNx+SFw+GQYkxu44LQvpPDbnnz+oL+Qt
a3fM6JGELbA+rH6ouBQkHILov8sSiccEXQMN0AeDnSAFH6/8FwYyxitW6ysO
GotcKOC6/VDRgAuM5UtEvOSLsOz5F2ESJyMXka2bYW+XwWoRGwvrDOPidkqO
CYz4eBl0eARyuDNz08pRgx1l/roKgVa8C/mm1XcAslRudh4uxOQmLe+az0SB
3ikPGCWwqnP9BiTFQI0lbPAVqjrLphKS52C4VxXbXycZqA/OoGzk+4c3R8xA
7kpoRrTmvOPNXthsrEuM1dZuimxDlHr3NfLhnVYxSZ20HpcsffGdJYdlLqYW
Wd+9Nx11DdVedmDVtptI+r23VW6uqM+77J1cdSdtZTOS63K8zjRigtsN2kQY
TJXhkYKV8Q8IeLL4EA2a9gmjyN/b72YHgGC3C5kQgGbF4NkTDAe8f2eo0Cxh
zKabisN6DWxzw3N/MQDAbZapWLe4/WTrCfQs8NpesK+q8j1he0v5p2ModH10
zeX8NS2yBYpJt0LVirjKts1I/zsULStTNcQ6/m+mIOYqMzJSJzCqOLWQVbin
yTzfpyo8TzLeEAhF0o1I6B5I2lqfJsAgLfnKCDmEtKdFMLCgqCPITlb3HqAM
FXNPNxWjkIT4Auj1x1MLI1SNgGJMptPWl92dwTctv1u/Lkb5WtEDvQuGHeL2
w47qtvFbRbdRvi8/bD2ltpeI5ka5qOpE0fUpnzUIgxEcsVEC0NaCD2pWbti6
nthmXbaTAGkiA1Fpvy+PVnVBNgT2NFdDR7I+icjqM49xZ/C6beyzwpLBYwln
Cd5aeIssMtzj/UHyKhMnoyjtWfio5FCGtK1dcKBHNKwtY1KEYc4QVhimT5Zb
fxjPkAn3F1vI/6UK4oWJi/Q3zFkKfk3/vuEgw/XV5dkTd/o3gJSE1Z34D3wy
bSJ92M836/7tFeWv47Zum+hoEsbrQCMUs1oE7pzJk9vLkBTYVOsGEwzqlE0E
eHC9emRjj4tz2QXEvzS1WS7dogNZFJhpmO3A1xtQSgeycYia8BS6GT4Fjcon
ycnULB0cEZnNEUZQSdGKkbHYA6KtKrCOLT+0uEfyNxURahJn5bKX5LhwIa2F
ytgwbawoSddvw8zMRkO3g24hyt8PUeMko/y/hk9sKLdADGsJV3jN17nw8D0a
jswzEQEszX00SviIzERSNxicqJax5aBn5fcaBLEN4mnhZbAMGnR+WBAOk7zW
/SZawYQHc5L9YXKBs4A/74XjZTzgT3s4igKtjAunWeoi4RirwQiYUZZROSkN
qGdHE2ijzmLkxbq1ysAYEJFTT1tPuQyTIBryCNk24CMS0nTy4gBRwT5WYjL0
Lg9U69XweJJRlOi/3FwtisFw5kzR0CblygpkD9ToeNJf/uIhtXx9DADKFW2T
wNUqYMfjBSIdUwTN4KvwMhr505jJcI3RRTsjIgJFWGafFingaId9N2EJyuzS
onQxNNHyt8DV1ApFm9cBRt35Bwew9DxSEcBV9cUO8OVXnz4ET566AGwLUOHd
1+zfuIUvQMwBT0qpNiNWdtnT7vJLcsajvux6P5LJ0zCtvx003f9VbcJQHv2z
DI6i75j6WxEpN4vC2SrBHD5frJKv/pLpobrb9gZ7PR1ldIVQYvm84gIN/X3l
vVNlvH9E06uBQBxhdW20PUYJONin1qyH1GBRlgSavPwijqMmupZ/N4JGsTia
0PFbNDbcXaxqq2crW/Z9N6cNXyNUR8Y9wD6xXuSLmNWQgg1hakW7quoAt5uT
MLo/FUVzRcz4Jnx1UlN2bsipx6U96ydPNx5yhUtMwjrwNdFG12jI2Far5ysc
WgDcWxvVbIZf9DyIH9VLx1aoibTIXaDm83vSH8bZKS5gxNUHIq4pHoMwIA8C
aOek1b9A9T0/4I+y2+qcpT3CHpS3+KNsGqZgQhgbVbz0LZ0Bcf6rh1oBd732
gblh7ou4AmyqzVuIGpLeQM0LgELmI6AY5MvpV5YoRD3Sfd4noAxRUODVIaRr
NMookbab14Z/YRczVc4OibtU5MUWKbtj7AjVwONNGMSdyGTUU9pWivADzZ+M
LeKyZ6q2BmYxpepK9bPnhfoFDH6S/d4ytqNkpi1qV+nAL/x9NpLZEB5WKn0n
UXl/VmhpX4uuzONBYGu8HvW8vooKg3Sf6T1TXgYp9+pkSGySkVPrzgXXnv2O
I3o4rsWvZQ2bMvRyAal1HqSWDwWKCbfCSRKvNto3vTu12Sr/0TSJ/mC8JyL3
jQpE0ODej+tYw8oisyRrOSpvU3QDyOdf8pOhJD6zAU501iYos6T+I7BVewZc
913R1na1bB2kp9LgTxI/mub5Ib8KmeuxsV1IvZgCvzFdMcIElKNTipbwSMjr
BhB0dwi8bjYVcLRP+MJhQVGeGrMchxQwU0ZrLYrFTPekuKW+kHkRCtf3dfaJ
06U/VVYnDKI5Liu6SX5eK3uTdI9b6V7DPmvUiSWahXSgjKGXtE27+n+8a03c
1a7LtzXbT7fJ8ziUURpd/ahawfbylQzTVkajDaSiaYQsyvCDkm8qkIgdOl9r
t+lL+D4Q17sJWS2JupbywqHEGiy35eBHW6mOt1tnomZJZ31mDy+nq7jsGbfL
15qBEssLarwrIvOBVuPeocdODkDM7Zu3LoHXrRSrLwrsQhoNhMmbNT6fAvLP
aptlKCuWw3rDZzcQYYssk3tx2BqSfH2X27NqTFsKJuJmduDz/DFOHTNsnwRw
Ynzsfvbc6tXsTG1Juk98E1T6V1MiZq8ki3n2Mb8vd+fRHmu7ljKvK2ugYDPa
fr0tamNMSrGNjqw8MwWV62Zt+G/lL9fyA5VCbbqQFnUeGi9o5TPfDEDVGBZ2
ZDrywKBGUDEypFTm+B8b2GaRJUBTPe70ik4C76FtFSpvAL+rUNjT+ffnr4Hf
PGpHMViS3UqptMoYnxeGCNQ7nHt+DFg6RdOvj0tGq5HrkygNgy+bjNMAr2uW
YRMXDDpkCk/AndZQIlxXJOmXuKUTjEI+Q/GZNynSlcaZmVJBEnyY301m3hVB
kuyHzko+6dmhgA1gqeKhbRytRACwA3weN6qsBwqkdLWSmKZBF3Dft/Fxq5Yv
N/89MvQG0WTQHrGqFwWXCBmxwyBNHe/n1+P3+gBLKCcRjj7jAyGANrQrVNP/
/qGdrxxxrZTdj10oFsbgiqahfA1KQtSwpop2KVADyESAdk9g5YvgCEHuMRmn
Lle2LdvOu85BVD3w6A4sk0cRuSuOrKqNec/2oEYGnUDvRHnRMyCBU3OcFUph
3twG+hgmDosa925rw99+F4eF6qiYsvYaLFERWGdkJrLfC3c0Ziqb921lNs7j
PHFUhGgDfOeQGkbTCWjaiGwlGXEjPQKvcQrs1Ko18M1UhbtHnL3xwKTAnMW5
t2IekBFzadxGFjzjgKPCsCZTdsHpYI+zzGyb0nhuIHvStRJp1mOLSP3EgRgB
aQbj82xUU8npNGpxHxv+AnEwhhx35F6krZRUJGaLWfnTp26p3ISCHvNcBPiN
lLWNFF1CxG2fidNP5/69KD7ocmyiJtUSxZwfv1SAN4MZjvYbTYaUmmBINUCC
/oCaSqiXntAyxREObqkfuxbmxoyZqMFnRsg2kknTs62QAGUwitmw897CW5xc
yRLQpl66yTFsU2X5QPwg0jRDuIRwME15oiRQ6IPVLldTkMNL4dzdUPv3Q8ab
enTzhoJ2+773bzWqwKMG9EvziklBJ1yStKdXneKU41/ob/larZq8qc1k+IOz
7Xy5d+PJy+vo3xXpE7KKJwJsyqjQoAzthmQ4wTrTIWC/Jpp0dDjeeqixLGQQ
tBOkZkQdd9PLMTBVaP2/dSrB1MkGcEsn4vZQ2smSX2neXgNIKI+7o3KB0erg
82EX1HxKS+Yohard+RI5Et9VaSOgwOOzbQ/hVx3/KXx4G+dfGiioIo9IqINU
vVvNDhlXeslsW8dGMEMr12gCx+gB/y8FF61aoPmO7UHGpdkwNLIz7lAfhKlR
JT1qp0YG98IUOkoVHjR7d1oL7MtlCwUCfUfb8vV4PKWuzW+y3vNYe9MG4u0Z
c/5WIJWEvPHTQq7cP2HI8v9+0sjy9rchEsL7brcAgHbnsUcOxKopFwfmwj8D
pK10lbRBVvE04QPKpqWwOW8kyls743bfVbNj8QFyGPfVUg0pbrz4/KCzGSxF
qKQjCFAXOt+QOjmbkg55VX35cbShUyBlTOJnqyS7QOkGHqT1B9yOxvoi7vlb
5j1Y4abVP2pDzCLK7xH/JNlacW6wO+N5rZbVngdeEc6kwBXhyYhg7NGFh7BS
tJ4duiXtSiS7Nh4ArFgPaKKkEbPne0mtYw5mWo17NYZ4QmTfd/04XEoFfiiK
7uMl31BE8B+kW698c+t8aplTi56N/Z5S4uQjeHE6WAQy85uPSk6raVYwlLfG
1vtLAcipPARS8g7++UBLjoSpv0Qd9XzAznoAB68dVUBss6A1yrgH/AqRtnYO
505QvQP8bE/MUlBwzaqv2cvXYFB+E3oX2KNg5Q6JJQLLSLto2dLFlOUDFJjG
hwu/96tVbcavMj9KmPGKC5t4NoXPFNd3wJPysd2bwW7pq3kOOiXOsSQLukyn
LFGrG3e3ID0Fm8/+amg0/yyN+mat77EFNe982nJoYGuFES4nHCzrbSX2yoSo
DYpM8v2MkI2AFzGmrLYcxdmXWEQExS3/l0r9IPrHM5qylVcX0ZRqntB3gt+c
FmDg/Y86eCWX2AZIyYSF0fSIeiJK19CtVryHP5fLuDEhTKwv2GurS47H32+2
Ypsgdt4wRJEbN4nSh/Y6etNlb2/aC1fK0zUCwOKO5fN2mzCxARiXBj6o1WYW
QIzcyRmOsKoAz+6upqWKEpqDFzM3N3GdW0YT0FNE5X999r1Y+dy3T81HQemf
FHUN2hJ7aIEBrtJrqNk+VglZCdAWpAwMBLzq9sXACtE6aG01fY+k76c9YBjX
4fIQWqG/2aU0HFTsrbkSaFs1tan80lKpb4ZAbB+i0l21WHblbalvMYFiowW1
H4fQX3I4w+S5nm0Ei2FvaFZLVVeRgtMT/58HHl89yCPQDWvF1G5ElrMQ1GYU
M5p+RP1OFcF9xYCZnAYkaMAtXIYtPgCFPbOGbocwo8h7OzlpRX3aBZEBVgpl
ICZ6G1c0gcdbFrMUVJ+PiqZeHqfqvGLOPQGHF632+xnj9uv0xGM8pJfIgAO1
ygEBhKqZ75sFVRzS4FvsfCb8CeP//SP/UpFPJRRjzWV4u9qXIUG80aZHA1eJ
NDpg1XVDmw8yAkz6eflIZMFNypzdvdMdzfZJRlm5FB8QKHE62Ly9kEuNXAWm
HUB09VQZmyKBHExvP/O+jGAYCHQs9gvMYhslYf6Kr+3h8YAHFBvvGChJ0nEj
tOCnZBIggnX+r5b0RZBelvzR/vyOyzzQwYhgwgA+QYcOY7kJxGHmgzTVB6Yi
tqNaMY+Z/lFdiN52lWoY2K8r4m1o0kNkpd7egxbWHNMEIErwm0/egAI17yzb
pHpSH3e+ukrzF3WINbHtUX5YIY6+MXNDiwdmezQDPcEMlRIKOp0VbNnzkACH
4hTHGdG6GJ3KWWlPjB5FzMupqIgtPd+Nv7TFz+0oNGYfwG0+WCPClxyxXnFq
txu6SOeBIdcMvBtegzA65XJkn7u7GjP+K1ZTyLXAoiRvbUnZokHKvEou/B5z
yjXv1MDASXC29IFAjaahIgnpsueIfr1/0uBkDYYoxfpwbuCT6tInsOkqbsk8
dZdQtjJ7bWwuGL9cC+559mizMrQOvYreSoIbfQmvvUfI4oBZlFLzXoVsdFJS
u/PHC6JcIkYUaoVpmaGDaQrRQCjxiMJvW0OhAWkJBxInWtyG4z0KvorKsbKd
y84En7my8xkU2nhlH+v+2PhiXsUEwKDLfr/qookqLras6IDF3JzzkM2Juks/
hjqpAL4l8xZlEW9lVAlrLVc8xF+QhM4w22LI7q/elzRG6hJ/zs5Zcu0HZdpb
dhzW9pRPJrTp/dXn00wRUBLc1/8nscgHKk36tyQOrPp8Ull8StPGFq0J/a0Y
I+XFmNuoPfioMy3KGSxlEY0tR3lWUCheuyYUzK34L1IIN1VNPyee0EhxZy3K
952zWW5SWQC59HXMASyEMvP9Nvs5qIRGjJtRSse2kHs2FkHO1ZQZbCGEOxda
Ci7UsZhCOH8x9p9O7wMGZxEsFQgwpocPQmULDpONa1MwxjpF1acBa2Q3RDCr
bZzgONGng8NGk9jX/1kUuwh1kkuj82nkFBvCrgekKvFEVvn8amvtjT3lpoUM
yRwmgieCAU99DBM4qWu7o8yf8r4O4UwbJjrVWxa8Kqwej1dPBPvwj/NFF4XD
NWRB5wgNUuq3+63/KR+ZksOuizTS1icvA2dyaNU8KlEE/zgNbjhqwHnWKpif
v8T734Ek3OXpRlUbB+Du1BePVAjR8U+p/Evw/UbIo/ZMDu/BETJTAhLpiDug
EUPoUXFMec0Mt4hcsSWz1SFV7FI/fyad/X3sSI5T7PZZjX7NUsaZYNAqmbrm
N7yMpAevQvI+f7u9lCDfEqP+mdgUvfK4IDuY9yJF8MGpvNDh7KAn9oVnYnkS
V13ObzTBtrAcZk+KOy/nchsy3dkvmDSkY7UF+tGshHVXTPa12F98SPPVRV17
q9yYIlWbu103isI7Hi/VL2ejgFQGnhtT2VmyPgUDWb2lJQlwFEIkTNYOWG23
Hpxrat65Fqwjo/9jTs+UF3MBerEcW8ZOKtoIL5FF1U2nW3XsF+5Lr8RPq8xz
jXOlJFNBW0eboPqUsVJiULk0/RBroyj/jS0cSQ0E2/UtP8zRAOvBbQEqQM8b
JvCDc6NlncAAEoQFQDQN0dRWpPxP39NeCrtxytgnB+OzadwwRLi/ZOf9sabL
uG3D4Y7FJeY5djgjmtK0n7z6bqKIT4RqOo1gEzT9Xwps2cYmBcXCJremt8l8
CQ/73HALgNaWCDm2bt5U5M0YqRDpRjYqHlKAsGQogA1DgKqCujr4+VvTUsOY
xRJc8NwnY7EDGji1FwML9BVQvGUlE5zTLAZj61wzXEfqOc0fiTcIt/ZMnzET
P/8xXGMv0MzWNlQM5ojrL62bVexB8qQZNADVq8kbMYy8mlpm+swIRBG9xGaL
077p3cxi7p1Ew8JwzuggJU3CCjfEUEsxJcNa67xKl8PDxnlH9JAjUeGW7k+k
vL6c89ILr0xuCumbS5CPpGn1W7TV1N/VvoiG20hDC828apjjknaZJUSb3v1+
gNlGFDpgsNOFyuI+iIQxZYD9BmLZ8oCzz1CUGQKkmIix/KCK7dDv4rw77Z63
OibEYcSXl8P6XdL3TSM/yIwkim/ZYvAO9XVGzZFuWyFROKx7DN9Bj8uHsf5O
FMDvOGOufMF+QeU2W/fJoDu0c/wo+RYXC3BaUxYaxFDY+AESHjFJ2glpxDd6
gINVPQPAK99toTGJCRyguzytFQYhLc0o55royXmeT5/9aKChVTJYj/yL1I1w
wLYz5ew2s0RdkkfvTFKFk8qY4E1WSBXRedRL8EtPS8TerotEYtsSHPYO3RES
1lnoUloPgXDlXb9uZLn16Mp6LqUZh4uwI/GaUeRvfKYJYOMIIMQGdr+zD4mN
KEZ2FpguYbb9sCl9tqz2EHdr/MFOdGBQzbyhuQK2IV6Y3bR27jIitlq2rEwZ
KMI9nbbhwQ2ER11bcQ8tNwg7/yWlx96m01xqBXsnU6aHmJK0HeLNa6+I8doS
LTASZy02QRa2i1XWfEN/paY5/1bYKC21U5Azj63udEqRMqiD/ZlSh6fMrJ6U
BO3f51FMn2RRJ/3dQDR6XH34WzTEyattK5kSvDcC2IJK9s6VPG4PEG6Z8GB+
hSSxNV/620lRC1tCVkEk5CCn5ILj7vOgk6uJ79gcTqPblhxg74pDYeeO5QgR
jQUrsIX9bEklXHtGsUe74Ip4E+VaobkIWKiZjVhFWrgVSF7G7Kzujtury1h/
BKanAoXosh1Y0TPT8YH0FCqVcByrJIQx69zigUNdHqFrBKmxTVb587BBO+LI
Jehl6NbKaHLD8Kd5ZOZ5EE1/Ge1Z1CF6Qi8vPjlau3n08mIur8Ye4MK6W5IQ
czxtoa3+IofDlMjtCJGWmlxt5XAyZWrSwfKLDsPSfA2/8waHM2LQaCJefwAG
jcP7IZDLNB+MBvgsBullROuTIjZFZqVKKILfwFj47M14uDeCug1bsmaYEM97
2vfgpc20TL96PorcYQxUWrVlmrPeJGo3h/SoGACKtsGYWvlggF1/ilJoYLef
zx8VOnI2RghbDZxmaRjn+l2aXtwvoR5+Eu++H6T9cQZhYpc/B3zZx3D6Dfza
UMInIjKbqrOOhHqSEHV5Z05x9PggWWR4NYJz1QJULrH4hk7HojnoDN+y1b+2
GzkOBpMRfHOeUf/GJbvY94wGJFECefw9LXFpYHDmsbl1lSuN89hl/oPzxE+f
p5uKtPmHFtM/voeBdWNNioWuOxOmhqdLC1YB2I52yEZtFAekn3YK1naOyPop
0BzIlNXEr6bO+lwkGI8f2FM1cT/YQsboyLGW3fyKQv+qbR8rJe1Pc6buRSCU
gdLzML65Idm+ECS/8ZCXVGpWITo8rrP4+Z8fTP0QmRUzrCwyNDFglzpHxTNr
5C5ZHEe5/g4zxJmUFHq6NYCFtRWVvMUBNVlIq67pFxpUIoIElAB0XmXAnDgx
G8oPU75rTBkGpa1BXxZdEMocvc0X97MrswQw7xdSZscL2BoxYQnnRAyMlSow
Y3vvmtfsgPMwPlVk9JtnIPSAD0yAePRlt90nnR2aUzadBlsqz7/0hbpdexmL
ihcfIGKTGt2uTFHjl1ufBL3+ELoLQdADVP3E1fJAVXWhE0oIe8LCR07nSeXT
hEHAOD/mePI7ioDW99rLjwVbx2sZXzXAWZIadu//OYWQX+d5dzqle18jpl4U
tDcbQJsfruObwbVQN/LPkUuBdGK3+9jQ2zJaiao3QgNZivYbtjTcQzLP+tid
9tCET7gtljfFH0Yvd0R4n+evXJJ20SFO2YRW8BW6nULRrbXuF1iWSFCE5UQX
bhDlw2BMzqtT9jgz5qJvdEu7AZOSu4DaVI70hB92Yh1Af4LctPPI3aHL1OGi
CHr2nYxfAbxnn/0R9bpfCfDAiyI/2M0Jko01qGFVeRP6AQWsBngtqB29Tf9e
dCOkvZc4WpiXPYfUPr++drB9Cr4szYYYh5/MWNFVZe26PYYCkDLd/74neKdm
rrcwFbxsWBiTkr2uwDxJUlheaSHFMDngMlOgyK1EAWXmZkaC5Uuvb1tdNoUf
ojQuJt5hu7x66a2ZuwfUyyyjYVbNPo/ZC4COpxL6Rx7mmPICYwH8Xp0y1iKt
+yh/BFGLzXroCvu6SGjb9JXNcwWfxdt/NbGRcXhUNP/g7DXh+tlAx01YDqbg
kEMdOfDYMsBW9hfXIspCkGd2orkRNhMJPJY+bpkzmeCKxMwiobjssCqtuTZq
60imnPbEK3y04aWoqpC5PglvWrWwQDSr3H3dv630KusLIGpBdl5X275WgX9r
AFII0W9u+BsQVAw/OsSTs6y+kV+2S+cHg0r8TAFf1kp/LTD+ERbKuY/aCNnq
hff7CIAutpGwzo3BBC6FpALn/25KIbx/i6m79OZXGe+SNxjcJj233l+nAFkS
8tjGMnG+J9j6zRR5u76XRI1rG/wQ8FrYG1Dl0DLyODbSbOzBbNM0QOQRJDZz
ogNKTujV+Q2T1tjbRm8dc2F+Kb1bGIbxy5BQtDxVApVGQ+PLbOoUIt92b+je
E4ATynl4d+7n06WTddvIrgYD2PJimBoFYNR8ASLN0N6TFR84OhXi02IwIp0s
dMUQmb4vntXtBxoY6mN7kkk12lm8gFGCbsE248IOnLFGF9r1fzzz6BionLFY
8+Rp9IyZqLZ9RXVGH27DdmIRqdk2tjAl/UEg/AHx9AKCxIML8QAzd3chyUdA
dO/tP33igF4dHb6OLjNPJkmg9zuUHb2IucZD9SJEEfoye9VM0CSnaikLZjCM
byd36EWgwajdVYYEkUaCbqUKJQgsWkDml+rlI5gzoJgur2h2ZlxmeqbqcSbJ
mIA1ool5p6576W68DJbfInLFacDBFqUeCoLiqynfhdxePvwmXCAViUwbHBWJ
3c9lBLqKAMOHyJXreelvbpfSLuApQ856/RNou3kl/aF9dKsAJmrKFb6CBWaw
v0QEGl+JufCigbbTL6mhUIllfYWXcGCLOR212xm8Rp7l/7qOZ/3zVTr3iSm+
QXEJ9rX5gKigTls238XVk9hd7S5a2uux/oLOkCDG8q+Zwx2qoehcifrhFlAv
J3dgYPajN5b6GIvGLN0b8CChsUaagFsxGdavhBc1eBGwtd4GWGujGIRo9KoP
NJceFHgRFIXdSP/G4a5LDf8VD3ToHKJ+uM3F8ibWkuwKhHbdCUmHFiHf9VbP
RNQKyj5Cqef2Q2vUcf1LInIWDwRVTJ7Xg/rnjTmPKcRDDNtmT4Syq9P0fK7/
L+3UyGpiNRSMoiq6oB5uKxo27haeKWNW+0qA7MjEtZRKmoFNrEpDLC/mPvh8
dsC/oIBrpi9nOZfaBS93ma3Rh0G5mCCzKAOhIlZabi8gI2/zSPzR9YFoMeXa
AM14hoXbP3pZkph6osXejXjjCK5tY370X2G4Djw4nqjycZ+im25SXPdvT6eF
u0aBsb4eNPcHtCgI8MCu6xldow0TdNFMdYp/cHIv7lgL24MZD3HvQT4eWFME
jlsYfomnpZ39FObffMnbrw6I+PvLgycWGWxytL4F+yYusw7xUXtzRQuEGDTW
7cZ49tejoPQJ3xFiLywZAdktJp6HsgjZ96h+MRgiI2eibMEb02kV4fTEtP1X
iAs6dcXqueicX7VpoVB8ErulZlBTdotQqF3RSTy5hHfFz9lSYxcyQqJCL3QR
LMovMmvpdX4F4lmWSmUoZCbyjMnybBMssWqzSUuLBptiZyownCz5iwTZfe7z
C8BUYnSJKMj0Dh/cpVeGtFoUNdioSLCju2knpcluhCR/Z7x362iMyR7x560+
YQONAF+LjUU93s1kQmWlVpmU6wLxNSgwF3JOW6IzDbGsA/O+ZAYFByowB+cE
PSnNdY/dsNwlvRmmALZiwFcDLVMIqzrOYsCdTqh7tR/GHLrb/AEhuJuYiD8K
zWmsBTuaAJSjZtriKAO3MP1VyS6rNma2BA+JK5++Q0feAKerP4+sZfqwh3Ew
s3+N4Fu3bYbp/IzktakMhmJl/r3if3fHMmgKerKKsrO7cCR5Ta7XXF8p600C
nQWezQKOdLFXZW5+H9Ah97eWkULNyxMlRG66vnWBlundCJw8DIJua95mdYZa
4AnJSBtXp8w5mqgIBbAWzyGY6+0SjsnEuE1pJrM8AQbVzohWiEPOV7Xof2hq
dEcl7HRIL1HDNF9gk9r8upat+x1Edu+/DHDv4Tq46NvY44LZ2bWzMMjn/ufl
hNYlumy1fs6OuEc71ykdVQpJiAamXdCo0CgPhr8q5tgAUdeHdEfpXUPjQw4i
AConP5znGeqrW9xzcDvQj+HlRSY71vNYGX0dOt6VUawv6z9QIEWHsYxa3TiN
ggU9Uw566h9D8Kz8vCm35kn39OXyX2SJS4WId7rWZf7XM3orH/9aW7S18c2w
IXkO9SpcwDPukBjzW7K8NyruQ47QSKSj7rIvKrnCixiV/VVZO4o33zSKrWpv
On+B7F+/7MiHRnSbeEU72K8vmUQ/txEoDFFF04ZFV7k8r+MqbTqta3Gkleqp
EkHnzLwveK/UDVIapgWV7iWRBSOCF1KhxDU/Uly9i098h9esPzuU36HOFmC+
JagyUe06s74f/Bedad9yBIUgBGBpKlve783vxYhksRmpk6omCDkkONjdCOZw
CHbidp2or7Q+kHkcyVftKNZnCHKI55jT+WFJ3bsEl7fKD8LHGAOPbr6yKAem
SkzosdTNQ775+Ccy3bAn1K3C9XzmFd92oXo/V+OuGMWZ+GAarDc8KP4MHW/6
D+PYEp3H3NO72ddz2+ztKyxlL5uXrd2xq3Z/qvKbBv4DOvBDRBB0ZijTuoRt
DM0TZ8wKzOZV1fnebjXux4saeLWHCc9ErDk6SNwJ7URb+9IYRo71T/CN7NmK
lpCddf8rKBPybvhGaSX2f8craBHqpH9lFUMGhQqmDtJiQcX8aTOzH2oRwAGN
1x7/IXSOwC2FCEtH0R3/U7fHtzIbd7DgKULCx7cWOnuEe+R/NLoPf5XXpgXf
8aTlQ13jYuUDEAda/JOoJiMFZ3DOjzSJfQrevWwFPJNkzglXs5/tBvETAbHW
96dEBiEshIRFF1KlQ8svUr0D8xxgxwEdvPLiYL1N/apOXbSwB54iVyJBD7kn
xXAkyQKJZwrPhlkqndtHaHRFIJHU572kACEPGKSw8OKkKNAfTVv5xv+tiGZN
pVOVNb0q/B9iiII8GSbBCbdJZN5wo4Hgd9gwrgG2CU1T5KWNzX0mCKs4OFlR
LKEsIK4rhN1IqSvJQ5L6ZzIjEmVpnvwMPUWd+FmuwgIoDqV55tDBh2beH/O5
v8fc3vk+YkJxG1u51BJT4T4z0TyJeEOg3E66Z4GOOG9wwscFGNfxtXHTp3ao
qlb9pC5eZZWv/HpSpc8V0zgUstYR7orVS0v8yoVX44G9SGnkm32d5T1YaAo2
Y6Vs9Ym4kstU+yLzduZEEGCVcH/6SHZbwzpVA4ZEVQy/6s3HFxSFVd2PvaAm
8x9d37Qvbk1aDwXxZ0fvcbQfk5TmXPxWQOA+JI9UosZ0n7T8JLQu4taoDrhF
ZRUSJ60+UxfxPg6bASLZMWSnFhSZJs8PpQ3aZ9fnys6kFoykhRDldedBFSPd
OvIBVh5UlEtxkfZyjNYOZVB3ei9eEPeLpgDaMAIFN22ClbwrJ+fyX1zwr6HG
O6C9xLNmhIaheN7h3EA2I3vNR3C/PX3RCvjE+Am5yr8ce4n6O5fJ+y42rS+P
nZtbaOLxtJTGM7beSS9+AbkSAv//NzjIYEK3lUtEZzFxrqw/oLWHD/dvjhj7
E/1SMH7Bs5evTPwFJKSHym/O9Eq7VXk52EYH4zDUoatNMXwZzKJcNoDqdXcJ
Ra7qTg373D4vyPC1PUP9IlP0TRXB4tYZf0orUeMnLsGUU3EXE0pB/cS7ZkO0
E4YuUcpnkSY35hvHdCw3OReKnfedpnVwmSZ7WaVYBwz52OOkYQwAwLRPvP5f
9QPuei3uNzMejMQN4rZLNkQxXb8Ecq9UCuh6R5GKBRtbtIVtgC1D13FarhGI
D2+zD3mdp8zIhkkUhqYr9Cu5Kimp+nSu9U/AA75luArmlx6wHXTf19t7qPtL
x5Bsx8/WIbRH2BnEQHwfVp0t0SYD9MNup5l2V9WY2q2lPgw9mQXlRFHW1FYh
7mOLhv7FrlTFddRzlH3X8WuPyw49wubBuB71Alb+lAGyNMLeJZeZdXqY0xI7
8wqayx/NYidm8SxYsrvh3FpvKl4NH4TyafdyFcnMqdGZlPi3vQh8Ez+rZFST
xziYKEbUfXNEBlRrG3e6nQyPHBeEv9HS+dGu4v/ExrEd0Lx1bRvxbX9MNaW3
lM8G4ZYUh8vNd3PE/h+jRoDgXhTxltinqikASh67JjOYqQk6rR5CXI9sDvFw
cAx/tSM2SR2dG4PuYt6SqeVoBWbWOBoQDN1m4o7+1XYLBy38sGc178ZDXuxS
ug6QxR1fbqm4pribEzSKy/ZCXBWF4u/7aIQ/rhy/2BbuLLyUYEwlnmTQW1Ea
KrNrDWEPCFfFkbMROBhDfhjVu42RvUGHpkCT6I/6GJwegmqbIJ6e2mLvYkLd
cCOmxPIXLv+Q50HC+5xESOA+ZN6LbZ4WIXekoQGOZtwR77+Su+UdqTFIDAQd
xuyBO4bqmyCAolCZM+B0iz8ouOcV9I0grKRjWyuAjG7vDFD4LjXqHBiFLoaF
Nc4m7A1FrFjSBAvaoz2kbuJgge25+108O+w0Mc0t9ZDzBksVeGqhpOq3O7l/
pWYQAnXBZyDhelZ0iHez8e1WyP4Vp3+UM/bh8L7eOH0Shx9qkrG8McSW4RgA
1H9LvfkurAui5GC3/uNWZ/l4tAVMgi3ybM2e+V07wGvn3HpBoj9sNE3/FNv+
AUHYQ1Z79UvzRBaNtOUxjDkaJGusMamC8Uc5InBic8cTItR2P5GOLIlPXJhr
EJGOK/5DmYn1Ve5Hkxzh92hcp9w9a1zMeT3iLWFm+WYN/ARrnD2UC2AtZW2I
bUdEZaGZlnyJepQX9ddnve1iiz/1GrpkiRHFkCb2zor1CBKGDuPLw0F5XJ93
Za0XfU+Rs+hWYp0mzTHAeAiD/kYnAnC8DtpXnohp/Rg5p+664HvhPuufpv2D
cxRl+sMsEV+7aH2YRR0qPu4jAWzjstuM9PZz62ZEh2tRPz/E9+u9LGQV8w++
qexwzs3a3cKyYa1WmTMCo/HphuixdSiadRtpF8o1YbeJvMKJi2a0eUtdxwCZ
oIsxGwILp0uC6dW6IifoUAY6G2M7tAHKH436F3NTQK2URg6+C2l3btMfgO7H
IAgMES8knXn68oFZ6eC8Eapw2hD6EMGbVerRNLpLKiKeQ0M4Ig04dXFgEp3c
oBGg9r3/7jyXJDkQN7LyTSlyOxMMxADwEIoT+94C9KciBwtKPNI1nDWH42JV
qfuewqgu8xGQjZqJPbEmQv85fd7QHC6Vou3iKX4NuqeUN9qAznoEsYVt9U84
hcg/C0MhSQqZuHtWo4j/RNeq/vzzLjDcgcu+aclAAfQiGCDgwUq75LzPO36m
ZN6mov4bBV0DjqfeKo3l0dYgma+Zo4FSyv0Y5/2ddropMtJBNJGa1QOQFtMn
Tl0lk1G+Lx7j+gwTdOlYK2ZzSXJ4ZfD+w66TzhKlKmaEMEy1xqVYT7Fi+MrO
8kcMeQRlV5FnGrlUvBP2PH3baD08GVDqA4lKoUEwJ8voGimu0S6/ek9ZkI1e
NhVZSf1htYmUTTRvpKdVlU7yx5oU5gXb61W/iaSyJT3dV0xX9uuAoPPNsVmq
+O50HDT7ZS0oeVakAN/afTITuIdb7CkYlhcnBT9SPTtSRxSaJexqPfB/8tmY
hlsFjTXANFc6Pg8LmmkmFZbRyB2pPdKFBfEW6q/3jsmvb0Yj3zmN/Cxv22XF
Kbu8CGKQwpNsP8NDHCihutztpiv79ojL9Qa/cipceqCpuc0oKqPJZoUBzUbq
RqL67dEGQcK4rDonDeF/HN+LmU3Ey8/zb/ZhT850UnVfr+mEVJOK11I7xfh8
WsEsFFrFWwC7kBFy6XmgCaO3cM4Bq75HhMrf4bYlzqagkAnTcwirKWkNKwOM
ZskuHz3PqaLt+i2l8G+Bw7YdYVySmGZcvCgUCoihwEv9X3lLeZL3yGmvA9+2
AxYzKOeqAON8/jDoRMoDoAxM9kDTrxly4q62I61lf2kI3gwDH/GCPPsluOGO
GMDply65uIOs3j8YJp7tbmqK6xyuWvbtzQQyvLs2T3x7pOh8bIcOO8DR93wP
FUt9YOKOJ5xE+ijxT62M+c0uCoVYHBHWokOldVgweR6afjsQT2xC4S5QECG2
sjEag6TIh88tj7/oHo9OCo5xjbeGCUMw2Tzae9CD9BMPq4uHgQz0HGRwWSqQ
XzCJrhS60aNY89M5e0+oIZt6uE4nzhOacf802vimZ/fiYqiI9pz0TlOJ05hf
gdpgXnUAV7vFC4t9kJa/X91ZNwZUbU+YalC2N5WiEy4pDJ/54RDkTq6lY3gt
KPJyk6ywBKCw7FG8d7OVPu2O7itZka0VnZMuapdtpw7dYPkged+Hhaikd9BK
nVf4YI3UKSTi1Up/SQkeAi8HhXO40rRlNM9smGfNAMhlcBEy9NEmnMT1Kjza
lQFBN4i6rhkYBYftQ9GGlBLGOYlXIjGD1PvglVYJbYKIoaui4T+5I8XRYpOL
iqc6WQEvFCL/DXwXlZhYnbclMNeiQwXQxwQF1kBSTZzVxsZKoIkUM+rgDfZG
DRm/5Y0i4/vKa6edFq0/EA4PzvjvS04zrDdJPapbBknL+HmMRRlcZg+KBhTg
rlvSJDWyVkHEp44syE06qvaiveehtKVaQT539s8IsO6DiGTODnUWqqeXyLpi
5FLpRTWIneelnGpM1tdV0QfVQalkibjtlNlEMCf3tjcqPVH9UjWDUiV9ZSO8
cSjJpFxZQkRFwTkSovsolRBrRIG+mPti4UZmyngZz03btBbRyCcOrhqm0zIJ
iUiAEqkwd/tj+gmcRjMhtxJjqUXnIaZ/npoFhRUwVqC86497smkBeWYbh4Gp
d1LP/CYB5/oQ3APfs6x5JL4D++p9tNAW4fbGLNGnO72SkFdk4J1XzJJ95zQn
LAgWEcEB5ZidcnKiPvgZk3s2f67pw28q+iDPmTiWoZCPN9KXuEDb6OUVcn9g
OGM4rN4LZOBoVnykeZpRLyZ+lpUCEXM+y3sLqjK1mkoMVMUzWhI4HXoDISKN
fpW96Dm4j79k+LYrnS03GMwoxwnNfnSp4/OnbExwWhd+l/nvDWhS0b5RHhHq
+firyLpgEaPkIyIJinfb/XU1s5Rvre/VT6pqjmINEsgRMUdiaiHHRWHmqj9U
2XVfRD4r7jgRXNJjWLZQlYAkVEw3vMhyQFbI4Nqj81lX39ljppeuTz1d3No9
/TFiKdge1Qow4yC5CzkuVwq5weuSeve8huLxyebQJ03XyIOUZAXxh2VJViZD
Zt+cP8fzfog+oJNaR9PADu819qaPIYZN7jRqy9RdVPOvK9dqt0OBQohqAW0a
21WQtBPTg/X85bo1AvK1H442gBf8Itj5RfSqRSJ7gzMG44VIkT9aHGSF1dIo
2RFSxUr9YNi2DsTbEBkr2CeGtGqzBRLuT25mZx/p0lGW6z2MrcTUv9WzpamB
nuubbat8gYpTN5wHOcY4YWF9IfqVlhbNojesum5LjxAJXzaad5Vko24Y6j9v
WtqzLzsRJyHYLjQxZVsad3JJDeJ70540oOoqQr8VwtlQlhMrGAvM8xrqtF4F
YDaoITkBJ4Bt62nMhyLZeuYtQp77m0yc3efrDad7p78boKccsxEpj8iupOxP
ilbZfVEasipO5/b9YrPNXMDGy4RFrEKf8JNeuFPwzLMexIFpdhKkDuoBvbCH
5IMab/lmYK5l1uMF7FEonJkF2JI1q3LPXgevYOPpdjunoplLcQ9uO2ofxfBH
p+HreXRg6eXysxNx5lLQqdGY2+g87VlOX70pqtTMbJ0FFsja2uLBDDCnpWrv
ZJwFRA9B14dcNc2WpjuMX6LiEl8lWyLY272rRP8C9I4dlCTRKPEj0I4CWfpM
CBRMwvm4Vj/dDr6XCh9T8dr3ESXGBQcLMvZ1aAv4kuEDztBqz+hU/+OZwYc8
AgX6Zg/rLD3J2FVHh7r9UsPRXQfeyxAHl1F5iRt77ifXj+ilq7X+j483JbNu
ij0acfDXLOpvl76mn8FHBuygvIPZUPsaRNY+Jgn9mlGk+ZIl8HTBX48gG9Zn
xrfPL4YaCkvandDJOekkP9uVNlHJi0K2NXZQeb0a5o1b5S7gaM9HCF+WjoyB
qxGGpu0Hffq5Zfv1ZOW/EgflbNmV9JGcGSpFyGzK4YqJUU+F0G1oFYVWFAME
v+5UAvwatJaLqAjjtDHqvefrtWCLnRR1zdWJBHQ3gQk1WouttJCTM0HwsE4S
DdYHW8wDxfLUN6suLUCxI0jYnS33mld+4WgHElOTBT6kDEk4LtQwYJM9tnCd
/NN3AwWDEJ5pl3fjKOKEUnKDFS3fpRTm+cet77sGVVy8hjUzY2hP59PdmJhb
kZRf6un4zrjnvHeKcCzvR2zRYjg0MDksD2r2sMq0bzcxZbbk5BW99emDGmHe
sQEKVg9eYeGiOQV9U/kWRVaIjffmM94Hc7bMweBDOlhIATIDEkjgKpLUsqTf
vIkIJhma4rv5E0MLGJ13CR6q9LAqMXoEBxCBRF08GhfZ+W2MlwW07UhBA/R3
0XH/9ITL+b3/2ptHEJJQ/CkE6Hn7RIfk3CaGXWAZlMxkxAhYwbMvrMOtV2bv
51j7Z6GEDDH0X9AJv3QffEG0FqlbBQpw4e5JPH0diLGtpkgk8mGb0PfxdGKf
vjKXH5igh9TTguPMiMNna9aet/TV+4zTmpGlki7q0KSCnERQxtiODH5XQ2Ql
e6tsFbhksscVtvnQGv2sUs7h9xFY9ie9jjm3QzVYEZ4pmWdqFnCxtONi2f2c
5VLQ5uq0L04fmwN2olP4MZuDzpZfTyhSi5UIR1qXk6mW0Dg69mCQZpaGMJBE
qNhp/vQeCp8vA8nmFB1UiDJwHlU+E4T5CRh9iLzHnVBRWFXLvUG72tNoMqBw
hHZeXWDNz+vLsjQXSnhznD3rXP3pt0gihB4z/1iN3b3vw+bUs9f2ihBWdBtr
fMbLiERSFz1n3T/zg1Ip2x9sQJEDWF6h7qZvnnchccGluB46ix4W5TvU0XzL
DS1J/unq+aI8K+oHnSZ8f9OTKXiFWsGpvIS9b/f5CXqcuHqiLxBb2cNypAvL
OH+v14KVE7TE4AbprtU5bmlk9WjoHuSkVG2EEBUPRMD2B9mRseggMlTCZcJC
YHKKh912VvEGbBJCNCy8x1ZlOI6cB+9pyL4BbK8nryEzTFynxTkszwnVE819
nCEu7OVjOwYeL5ulPgeNiOX5QA2F273QSM5yUB/WsDpv5dg/PYUduLggYAYu
jOQFEgxIcL02EU8FZtoVUacW4l12Oscb7xPrBKtxGuptuNFaerffwXMT4Thm
LJmdYfSzHF8YMXet3hSRVbOpZWxaCF8yYcWlaiPVQTDyypqBfb54bJBSfEzF
jKKhJTRZydVFC4uqSUpN4qqJfW1C/i8N5SYy3/eswW8PqnbIIv9+BKROWTOY
WKLi/tc8lA/z65eVx76cNLkmq0ja9dFaATu/GKSuq2ewo0dh/Rd6MX9sVy7n
qKmOtibdVlB4Gqo3qmf3o4TKQHRhHefn6UG5ig6bIRqF0x5u/10GNlaRyfiI
i0jdGZvwX2eA5myUirS83q1MUlglcNiog1xCVItRcm9rQE8RMftVn9SgUxX9
YdJAKkYp7d2dzpbUws74K5Kz1Q1UBJMajERkVfOWa8x0mLNWywA5EYQYXDsd
46ODGrGwyFVaWB3A+Ek3vcp4E92a6S9UTBMmf4kIPAppF0BIqoTlK0dkN3OI
4yPC5H2TfNeUKPt/0S0wF42aEpmntPiyKRWWvPjj9Ngt+Fy/Nq3hjArPTvKR
snKTEQYhObIldluBKdSZZEhKjhos7dgRiYBQqGtdpHkfw2Sg5xEYlu1PX4Hv
xjFt8Zds1yIpBQtHpco9b3aRpVNlDnU8kfE+zGwQ+J0WenWjjrjMxJ4xutdi
lZyyarKmna2WSiwQ+mzG8RugUFJTCkQ7iS9bmGHQ1bdFPcvKyPkWQ1i7xT3B
GYZyRMsjxIlNJxo/85mrKJHUEuDFLJVipeWrQSl7J6GxG+Paq0Vf2zQnn5cA
oC9f+uRhS7jSoC32RD36snVryZZBpsGRFiXAOLu8QIiqAbYxGVf6TPlD8ht4
0IgeaVTD7iDyMHEHdzHSgPOn0bojfjWoJbADZ6KfJFrjdo0OnII4x5aD+noG
xtwYkHUGopRGutYYTA43VIztlJFgnA4j4R9utl0heSACZjl4WSwwMFtGRtCp
hSiTS0wpgYINDOHmonnAwJAgw/s48g4BmP+rwwaBMekyPmCy2M7wkSoMRrAR
n9IizqdXq1OJyIcsRzkcE35Cun+hZHEb5ASJIM7+Hyg9Q6rRpt3efz2xoXOt
PbCpHcGdUCOX4NPq3h6O7yEp/DOb6k2fi4YCJ5LIMA0lTX7y4o6oOgomT7A6
SiC5+H0hcVrF+FCdeOsVpbQpHZ1KHrLHy65xBGt8BJPbVQM7srkPKM6WAxzw
cBhdNCjBWVJIMF4DuT59lXp+OMZz5XhLA2oXI9cab1PRJUiPnXujhCvcUAMT
uef179I3Jgcu+hYCJc1vH0II9IQtZfQmPxz+XYv2Jk5423g6r2E7NIzxSG+n
3f3Vz3bchSw8lBtf1kl3kMFHBfR5d8Y/QwlVWbKG1CBTOendIrZsgGLaT8sd
pO87D+3liMT1xbuiWcOxaWAI7UXC4hAI6V27jiozlD1W6WC6nZvjn6b1W29C
tvNBxhLvuZNuyBXcul6g/AwWIZv33JPipEE/rdeA0azzeCn/DwzO8DX1tyEb
aotPYvHEHfVOBCCdx08tZ1PS9TUHpyHa1RKb+9zV4DikudqXfLhCXm6Lp2xG
WnbkMZOfgoIaPDj7iuW7HumrCeroi1I8YoCZ24SPmSkEwG1Kl+XIVM8BSYEv
YuCLjut9bFYBJILkjCXWHjVMxl2c6EdtWqPyAFpI4jS6oLmQFpmDEcYEhctb
qmcriQPrDmkwHwtbIzBVz2qjTIu8s2sWRZuoivbaVaAMDlnubY/j9XeCEDk+
HvQncvH/hmoHXMArZ69Ni6VL7a9aeTQjY4kBRR52rb1nmhoJoHO2Ik/PNsfO
siD7pj9PjOLqFWbe7ndB+S99QPQ+RPsfp0b8KIzmV7hdBfKOCZhlHDnXaiUH
iO9uIvTL7X4j93sX4z+V3kaeL6GmcGAr5I0Tip0QC4Du32FqPFGQ+jYYEMUb
siGvjtYb9NKyjcgTGYcDkejKoAaLzW3VvkztNsS7fJ60HHhM8D6zMCGp5ZN7
6z2scqqm0uMaTy3iflcGxO5vHX7QH9KtDkeQHmL2p38B4MJBUXPHiGXee+2d
Wnm3EzgSpvmS0nLagDonSDJ4m9OmqmFXP2/pTm+7ALsusFm8bPOiXQjpKNkL
r756Qscxn77zjtxD2ShdmbJ4PBUAa5RYPhTokxyqxv+QCfekeXrZwsF9dwXC
p+52cxNFD/RFAIAU/nHVRhzNoNiNH0TkS1mplYooDFghfk6xNHRGWEl0RcZw
w0drMy72ssVnwjfr1ZxcfD6ajWx+8E38Y9uZb+gMQMFeQbVxq41/+J3d09Fx
yGBcohzjUFl+zgadkXhobRTpmzo6OfAlHRqansYnk9GwbRSG6Upngz/+SeeB
O84UK4YsGaYUM7Cy38cLE3tNbnciQwV3S+QijfPxda1985EbzaPA9KBPmP88
memD9J9o3rjZeR440hJZpLTxreWgTVuPHc+9wTdjaupAZZv7vXC32xrzsIw9
Fa/KNcD63NZ37lxDXNIvgJys0KdezQ2gPJ+5K66+eaX1mMDVJrL1YekD/LI8
YeYmMIycml1Rvx8XhVuShojqzwTtrR2CfLJ/OkNczFbilDeX4qYTIJIwv2ls
AM6GsTtqY0t1RYkeZtX8AXzmOcI5ijcd2Z7Q+iwH5L7woKU3oJzwEpHNJBiS
ErC6d17raJtVKWvRmO5YAMW4TnvTtNE9eHCCstQC+HBFuMBUWHFOEpDxw7pS
p27PK9FxNizWXWvfyIWyJKIduO982acOVe13fqzqJA3qUh7DWb/rlNwYcFaS
fnvl5r6q4IXJAJ0x8L7TjAsBa5GeMZJbF0OhrJ3nLo3Ldb0ncInvxb9ylNUJ
KJT/amH1kxZVeHEQ0BfhEd46CQjR0R+g8vg0uYlYYRV9tHML1ftn/fobMRg3
YHRaTmuqBp6ozDGo79qGDdMHGbYKndlWSOqLyj2FffNiUb0c/qtKjIINE+9V
BsM6mpqhiZGT0DDxY77bnhrCi/5SY7fYW3fGxRipD3LGbHqqVEeLRoShE9+J
vR5PqHI6vmMoY13rWdTyNrzR7jY/pEgXHSQtO60Lp7aL5Tv5Kv/mWyN4Ay0q
s1OreITrJMRS+EDmR1eJY47Rh64MNHqS/TgopdHZqcZ4BbNqX9ERbFAdgli6
U1iBUygufzkLSOHKIE/+C4DIEWlwSeHQpHMJSzk0vUfuegPCb1IsGgk47inN
OrymVjBe2uJEDBLgWZRjjydU9M2UNEgQPQrpu08l9RThD14sEmwSyUBLlV8S
j9fFpMZcY310WadQh6bq+yQyuFIABDwdWuh38W4lYvEeRWFqyBgnKvFtm6+k
ENb1fZT4fzzDrk7ODZHKkSO113xX/xZQWffsiaQVpZ4BBPaI0xi6tmonymnF
DcdDtl400hqh038s65STkE76LjeNTOaD2Rx/IbY9cGaXAoD3Sbi7QoqmMIxg
IoEuogexui2cO+khwwyAZmTAhhKa4hdGfzSh/FSuauWW/dtZFK47I2BTXl7h
aE9D7i+K9q0/eb24/LJLiLOfZ3xrlNhJkJgMBHztXZ1ROqO6fBdydWC+GhjN
MAtP/Q70OjbgUkdXYHsF7kfn1wxOo4wgqKP1CwfP1R7+EPFHvFwpym2jXA6c
5ACglv3wRxtUCwQZP5/3nHQnsP73exTRV6Qb6F0sRl5jYUBlxJVRNvet+5zW
VjJDm3TWavTq/3tYzmuKXF/TmKECE2e4hl/mU4gR+koKLnvGuQygNoqxRZ2S
JTTcNNikzkFOH8RlRTFf5V9rS6x15crciETBQsgJIvdhqRzdzOT6yxlkwqqJ
6MVPkMOridIIL7hEBLhp3rml7TCmWKYSy1jEHNztwJDGG0zvihIkF2XiBIV0
HutjptRyZiZxuSQIj+aA1NHuEjhzSFf1Yhwb1Q9JGJnaNIa7wdEkDeWdV5mo
7u7NOtwRcYCusJJdQ/S6yiAdC3cZWv1V1b5nPqugogwrOO2TapTQCZno2sPa
2+VD0iRgzXouN12cfScIO7iJu8S6yU9PHdGGHtl0xT9mYLHmlpADRLIsWPBe
Sm7V4W84LQMyZ+0IRiBX0PqFs2yAJmV2B9V2tOlWWOrVlr1rQJT1kvBU/tbR
BqBvH0WIVrN9O1vzjAvazn4XiMqyHMiwsZvQ5GFqqWnC/1UUfqou51vGTNR7
VG+z53Ma6Hy2LIzqzYHLGusTQGGi2Orm7IMbC0R82Lvy8CFYmBdXw1v3onhL
qcgIRqvi4gJBNjN/VPC0DPfA6vL8Ruofp6WwEOSvjtlAAf7gec+Etg+ei9KU
H2sg3ZuzsS2p1BO8qmT38e29fmvkC4T0QB9Y4VQ35musMwAjXrRPkFrE5zDg
6c7oiwaONZYL8AYezjaSvSyysDVgVjXDNMFHzv7ZZeYuAbwHDPNumgas6YGI
/jYhK/TAoYFoEx0AE6h8Xh/5ITRUrZNXA4y1KT9MhvP+JAaK4ejg+jJCcq13
FR17hZ7bv0br95w71AmwoL6jxU/alDd8TZiweM0+MJoK8iuCxK1ArESIkwCk
bkaECWXFv3MbgM9JgFaQEatnx0KdI0m3sZ9ISPlL4/ewoWLiHqavqTtmI3yO
640w1AL70hBWFMkBMZTJUVt/44BJ7/5Nm94MYq7pYC1Br55M9SEFVvThZ3ey
sBwO8gwolEjDbksDkHamlK7UJ6upLMwWfpF2tPH9nXfcx5W2sXVQNcRztpzK
x1J0YJvRfVIOCa3PCW0syyi6+wFJ7yUlyIij0Ls3uOHs2G6v39aVzoU9Fbde
Pv083rgP5QcgqTsqrHCFcK/XOHkWysyq+/brl7X0AKmRiFOSmrNt5FlQXB7w
rubzKVnmecs4CmoJlDjiCv3AFzrUQCkQqL8XXqrqoiF9+WxIkK2GRr8NLkkd
GL8t12ynisWfo5+oQkR2BFIUh0pb2i4Q5/ZeqLhwQzSPz/NKpgNTDHF14/pS
vqjxM4ikXnpENiFco+crJDb1QNOJPogo/3mYDLyKcvb7jrvom6xfNJW2hZNH
hhoW9SoyiXjv1SdO/NoaKAvfePoFBvSBoOC1KvlOhB6mKxp74/iFG8nWx0Dk
MADRAxl06D+8Ni11CrYRY8wPfqUAE2EJWHaz1yjbzR+KzUscCWlBJuYZu0m+
aYVpXTNfPNwL1iSx/vsc5PpVdPmuX0FglXmx/qCtGIrTgOSx3pU5cmlpxC73
zcianccw6Rbs2WfPf6dHquUYgiJ4ShjRekfVHXEi0IwMkgc3YXd/K+Rusr4M
K332oF1msgRg2OyR/Q7crqtubMNJfh19Z92TWvd2DMjSSgWosVQCouQXg6SA
O1tV7rVEe70siEmlnyk3/A1HZ/Dn5rk/kzoqGuqiM/+sBsztRPvT8iRoZ3qE
D4f80MUpQlPqFPiT9TjwbKRc8FSqna1dBmBFZDVzVliqquUORH1xJf8mVHSG
FlbdNAr/Jr4oPSeQ7RoDD0l2P2e8XCR8b5anfSxrlMXJWPGHSxK0fWILI2fN
MHzntNnoqrEtqqmCUK4dbuaZcJoQYgLM7yA68kXF2GnCNFTqlu+SUznqUZry
+xYd9TVJO1yES0Q0A/t2YpSibWIqZBrS1z0BEthRaXiABht2J1Xm+nZX8qcw
bMOE4tYmqftMD4cN7K75+cnMWTWza5H6MIfiFTF0PvtRDtyjuXdR/sFC03lR
8XsDmXyOgA9Im2jo2vIn4+ER6vI/Ev3/6wDJR10+KOn6Qmwy6LlutoLnypg+
c1gDhDrhkRfRwXbpdNHLBz+J9P8lHizAbmENykksIpnph2BXY1tFCgvcHpp9
N7kvbslo13Fj/oJJSw1w5NpEnculymIBJNtyxAAL+MyCgVlV7nNygNkqxFk4
5p3soE8ZPPxtMsC++AXs6J0rsoVZuxmpHkR5h9jSLBcWiOUB9oGZxai92ABJ
xbtJHKG9vZGBAJvwz+6Dgt0Zs3vU+Pa9fmrPRU2Qa+Dnachn00ZY7HU5FOH9
WSuibZ49reDG/SdSrL1q4h2ZBt96vVleo4DwSFqhT7c+JNfl7JanKSaDGpvN
y084jAysktdmPnulc1QBE9DUMY197+LhpHJc3ENeI7D07wC2cENqNe9qJ91Q
9uDKuIhekWKmg8+d5aPzt9+yFJqfh6SrCXaRNm0ELENAWuOc5ulGRTL3xxN1
iz9hnICO6Sqd92GbYnK4kj6w6UiI3utk9zcr0KsqZkz6vBUh43zjiyhdwtvX
0ElkV5+QViUC2s/g7Y8RhVimtP3HV2xtuqR2Uy8SGl3nJJ4HowASI4YuKqCQ
Oo8wco9zhcmzIQ16S8xsIlp5sR3XfXQKdayFl6VBthlNIBZEBdjU/dx9lynj
ajIM+h79vm73dyhuneb1NGOjlEapJCsDG/z8B9JKoxLSveSvaKvGfApCeQST
qYXlbMD/aBwcal1g4/Y1YsP6pCMESJ7AGdjKEUeF86E4amOon66lgCjVQM/l
+SXLtQx42Wu60vyHpv+tD6+N3ALrq4/YSquz4CvNkhNUttocRj2YcxuX3Hdw
FpmcjS057X6BCLfFBtJWg+klCkLIpgu5k4v1cr3CSsuF6UhC7jKH7E3u3wNf
FnkFSyt+HRrrtCSR6UrqjzvqffxdvUzlU+YfS1mvZEMOfzAN10H5WslEz+jW
wYNYgB4B8/6q/QuKPFujEP0O13enMnRHzztRbEKX6SYLBS2u4SnO6tAn1gYC
DeKzAtO3KhYbxu0nlutBd8NcpLFz8ZWFjJP73dyDquc2Pj9HUkOBHYviW+e+
HZi5ADHGgF4L5lDmc/Sua0rtPPG8YCWxUXiOioQhP3Jshkv1YvShIs9MousN
/r8xfX6m1PQugh7BzT+3prhlMbLzB7VQwX84VnF7u90w6EE+MGonVj8Bjdc1
qPnLokcKYTCo7le1SeryPjvJL1khCivpN6JKinil0MfotAA5gfGJbddcymVq
MfqA961kpb6DA9T4B3HNG43SsGjdY6PNY/kf9WO8haKb3/zeOaS1z1zxTerq
NBvWAzS650kkllEQ7nRFk5h5Adm0je2btecZZXnXeu4A9ANPgNNdIMc5Ih+O
K2mFdcd1l+OpRlvgbqWYt6A0vcwi+Ryvi/SNKa/K59atEEsvnu0Ww0uvq1J0
kmLIsS9nKsMfyEYg5r9rTruC7SEQPDN4MI45/53+Gjdh2R4BbpXTS58KraHG
1yE63jAPeBvrY5FPq28ox3WqDzgJwzj4cc/63E9yp1Qdy8Dbyfg4fp5hLJVR
QoFOy74plZ9fq/xpXL3Ip8gKCGWBa8c1pRNc8vMihKTZZsZvHBj+/w45V2U0
08Kpto8cd69cUJgw35mWx4tjPjoV7mjcDn+4ZpfWDTN5jmbinYEl9qMj+R2Z
EVlmo5KDd+aQCU9xNi509W18jQLkD41lGsWpm0uXD1RL+foCiouTpOHdFFqo
5k7tjZHR1d63GGdwzMdgrkxVQ1NLTl4thYp8Gf3foHq6XdjFCZ7HRIT1tJ6u
rIXm0QxPCw96PnaOUxA78/KwfRpS8OrYlQDyjueQJrYNma0NZuB8/+/URInk
5DPGiuJOFmzNsLkQWIpR8Fzaqj0X0sPse5roiGmofkgi41+WS2IPYEXp8255
VtzpQ8JEISGXKNw8/LjnlXtRxFTKNQdrJyfDiqsTzOqPq5axPDwmIwq1IJ+h
EgVy9B4pn3HGAKN+e0aWHIihkkayAV5ITS6K61K+bHX4+DyWwxXnrVcceK/j
OxhO4IvQ2hDtcqhE7DzU6pMLr0u/0IwULPzvjtuSKVGGOkTryTn1vFhP7W+y
ctAKlxCfx6h4fbgJlMTBl7qyvbOvlnJk9E3ezUYUkT5IIkT9j+0F7qDKYPQO
gsSLdoaxJQKKvw5eTqsA0XjcYg6Qqo27Za7nwgNo/XlOfc6XDlduzhT0dkWN
i54bzPYzzw4wKlEFZexzmjUkSyKiGFotyXJiOp6/+4qm3yPFGh0Tdmu1QMmT
MPcVHipzp5/iJbyih82pnWI3lLq1LckSKCr2tysKYbidlokCd42QZjEps/Ti
4IFU22YGoqftFMiSju4Q9YSRhLmth/JQRrpxB2zuJX63toT4PgxRw2eaq0cn
VC0ESL35kilXkbjhezLP8a0af/rXF7RF2D/JPo3GTnZJB6/hqH+Likwo6hKK
IiWGk80VPl6L+PWqm/fLWOAfvUvUsEc0AD2vJ+YfGCKyybyW1u861pSyMPc6
EuSyIzA/78WZ3EbFxfMZZ8HR2Y/xocysxEkPlZZEn+I40JNkW5iIVD3vBeuT
eNLIGRXxbGZRayFaYTxcC3YoawjgSszjoiNa/o3YWUbpYsEvDSw16TNeanwP
TK9OPooIZVDYv+ZUnJQgoMAtmh7TBLWlsj2XpbbZ676PGX36t9YfTqmMaL1r
zeQJKImXiOGJcts1quSA8ukIZ54dRmXB7d7wIwQMQhFMGldf3wjt+n2kLa9C
NjENxVA43PfJIP57Erw1EiFGWDVOCkGmduNa/8ETm2qJ6OAGI6DwLkFAxzxk
Mh6rbgZ7M/nWR7z+8D7OSLUfqfdfeo9MTS16U16OqINxGB2hFcdMZufirpL3
xbEKqXw54Pv8GslLwGTUn4HINbjklLA6eF4SgKBWNIMRs9WswA40uKfml4y0
DvvXgTA320yBTSVNZloYNmJw25qfDFldj2TIVGt9bU36w9ZgXDX1tZ7Yrs3x
GAH4p4O8PdRaDZp4lN1y9lYsKAEAXzjKU9UJxoi2QAmSWPjUv6v++//M7/Lq
4qMMBpXMmCOzmjwF6rQnYBH8OFC8HlAiYuIVCLZyioM6WIuqFulNYWoWjyzR
2wF47t4e20xa200PIMcWWiiGJotaMewM8obUQR9H3JjlH2IdJLrEK6lvaXxi
DslEnIXMFpp5ajYZSqXhMc1QajHa+C9SMmBxZJzCMlqNEah0DZzs3UgyzNvC
7lbLbjPk9tURKub0nyk4QWVCy4exH24ZjDxQalq5GHV+QHgyCDcxPiCHcnS5
W9XTC+sh/3swYqiv52ucdavrnQFeoUG7Td2E0a2mKi7kjShq015pnYCGsN9j
tHA03oM7HDsa+g1feTvVfmb2xCenMDBIDL2enSC6m32SuzQDCEqi4AYLEA7S
aIVKgtCNUMSABuA7w7DRK3B8O6+7CYZaZQngzCA4p4Ky5PWVvYsYT+eK36GC
KhTAZd/gnkxb4Y51/Abi+h36zibG18skWplV3C9DiPqwyHqO/oob/bqy1P8v
ZA7UNdPl73H9EQPvF8HqT8w59srR3tJCqa6orjvIUOu2WyPHvkfvoLb/XpfR
CS+skNv2y+ArJ0DFfbCDvyrBR5Rhh5QFyespp6DjDNDDfF5DMEU/fnY8ED+Q
vIE2JhTgAYhzLbgDKP6V8X8hYrEkgCr0s9Su0RYThaN4psqDnuL6cugk5UAW
m1HT4UDcZEip96+G4CvpAqi4mI0nGZZMpoQZkoCHypwIPR+dWoZ496dNzx5M
eMabIR4lYxIrdddfsQR/HSYgOxgsfRGL3qzrhZhJUqP4rPfzr8BMSdmY5h0w
ck4fdDByMd80CJQ3s1veHnu3mDHIiwcPWwCG6kcFBFZWI3nsY+Fvk53hDxuT
10LmcwhQ7E1S1Zv2eZFegi8FnXmjg2sX6uLe+O7j9SC85v7zuzx4vbv4F7qn
efooNtuPuMa08zp40LEZehiaCqw5n+/g07mjwfHl1uQvCXVbP1YjpiAIOBRR
e43FEWIOzGK006XKyIzS8sx6XRD380grtgtQYu2iihMtls+hMtbn935qBzvJ
SVebYpXm9FRpt1PDk5JcoYv7AN47/YnlF+/6OBgksKMM38i+fLQBbq1VtNLx
WsMcgoJZ7xQLX8S/oqhgnWIjg3VttL/iIZ08OAJJqnA203ENM0sA390lHUqi
73P02TVPeXVp8EbLBAHy5toR5WRkaupOmJWBJBVh/5aFhAVsqHCtP9ceYZSO
i8VC0UJq4kq4x3JT81Q4iuxuZAvHFzrSIR0Ljjots7SFgpM7CFnowVwAmXMk
82q5aOG1bIRzBe2L5Q4ObzIy6wObEpUvz4OmYjOUGWt5Ozgti5f9QLXPKLpm
KE8z+nOzqvF68MZw89xH+Xf/7rQeqtkeEZfJ14QgbxJRP0zQkbt7djFwIR/n
hjIbEmwCPAYf5CsB0H/nJ2vePGSxow7XKsY4X17LN9rSA5i07Vo0sOdmyrGU
3/qf/Wa2PH4bmg0NKowTvprgbEpNrJdC2gTWwOcCzlCrGSiywXlZo4n3fOoG
kDolLdfIEgLkp13WHxcuAh3CojPUR1L0+2im0zwScUCn/s9OqqPk8d7D93ax
t/t9zYBqqAJENX56WSsIBRm226BJRGS4F8dGGiez6BUxx2BIQpj9L6NO2gcP
/DXYoGh+dQnekn4ztm6SNsnVRCPpBxe2Mgiupm3H5wEu6xosMS5/X7xuSQ62
aStt7+mufGdFVFVGV3BWLOVruGK4PV2y8MUgqhx8PPfYnjWxlU7rqI7v0vYe
Tud9FQZiVe93MsTInIpy8OHF56Z+UBZOJg3e1ZDBj7La22fMzV+3rOZDIQuf
NxXLqE1Zd7BQtn5kw459ZTvvvQFA98V8eyOpLwOWXTwPh9hwSv3+wxN9o7+G
wwRvjSV5smmmdRloTIzP9Ji0YUlI45FFNzAsAvrZayaIGFJjyM13pMZhcUp5
3vXTO6LkZecyDyEYw7/SREMiGaDPp2jYjtiKC5LLEWsPIYqPxngu//vDQuDO
w0KE3QOoKkM+dLj9KdNBWkVFMlsGIgdFOFOf0IBcQmDZC7fZffoczVn/c1EQ
yTDTq/NjRJwH18w2kNN7oovYA2miqw89nPXTs2FeLBlYYYA4m9ZXNQLoHBkK
ke4L04V0Nk5+mHGYMDql8Z5twbqYSQrAbB/E3u1rjIZ3wlqUUYUFw8pKCbDr
P+dSuLFp2vWYb4c9iyGmVVE/lqo8JJvFFoqi2BnhzSWRzs2MG8sYmLV1fDZt
0nGdwLYVyIN/g2IuFogInC7AJIzuwtZkVbWpNEeEvsT/dmHE8j+qgVReNZzW
JrsoFIORVUTrzq2Alv7BrwfQzGzN8+ePIYSBMl/pZl5JG1NhECynehxJ9xAX
v549d0o+ezeREnRuLOWYRNfVR7LH7NTXf+bzW4jA967fDH+R8YnlTxD1J4jq
gBwoas+1toTrK2wgqeE4/tG+ASuF2pEF/6HqW3QxM0NuPS5B+gDdByDbR8Lq
Q7p9wE8lFVpyjW+jXi20gTZxUNV0A/RnWg7zlo+nW0dBxuN2dzoIHnBl771Q
/cJCWZ1I+ibM/hHHbMONrFbGNxU1mebbQ8GBt4k8JrtpGpz92t141epXDaiw
udxAIs8cbE2FHb+merLztUtRg/3+7cJpP8HBHKLWivIV4deYFvlMq3rdSmd3
1o3CAzy0hO+cQGAIEmEazT7yn2YBDTxMrneM7fjaMqa26NZfwrc5Mp91GamI
eedP5Kgrh6p54MzaisXkeDCh45jxZWS5zepafeMrKhgeisnyXC9+OWFv88ot
+8zaQtrKh4LRtcjvpTE6MjRuRx9L/JoxuxtcUTz0p9wC/hFzWSgiDnOJx6DH
aWR84UCYgLUyE0NGeRviOUXuZVOriiU9Zunco+DcdaZq73k+a+jLeMyRJcTE
HdLfzndLdPiXpyXc/FuIyqcQLcnREt5QMFdUzV8807ld4sL+jiqR4CR7htX1
amUerYNovcjhSTJU2SsphNhiWdgMmN2QFhrXmpzwa17JpqsBTsavDckefxCn
SBwz1mkUKh2W8eV+HoSU+uwQopTAsw9tcJ4OwXF0cKwexvfiFEXiLCmZRRss
4OBA3/UJLAu87reG5RuNZVBTIjQRFUlfPOU3IIHr+AGM9pYS7Bpi5x9FnDkN
SdLfWRnm6diWfl9I7lY7QMs4Cnk8XJziBCLA15wCRDa0cFF22zGofLY/iu4/
EyycWqUuTWOQj2CShdNNAzVJnpJft5LwzdOwzzQL37nb4wi4fUyPCfthjp6o
zdMiSSyb2ScG4D+lpzTKAWTTmHJE3ga55MqTmrBnM+QXPdrBH0PgVEQFYtHC
uDkxEYhqagEddSiA6aCx2GegOoZxeDoejgLID3UEsTsRy6k/KVPwtrwx/EOg
HxkZ0+4BKwwiXmzhMBtvv5lGtzq6MzJBYhDyH74UMFJlJVAgkQIW3bC6uwIj
5iAv81cW/Xbf3hILHARmekLKU7ncvZq5z01Jaqos8lteyoNFBNUZd78ZVQhC
CHY9ENZuOKn1G8iYhDHZG/Lu5A4buncnvcu7pxKz3cVhommTAvK+bp92LJ1y
ltHYiYnREaOvk3Y14kJrlOouaSCp8T4RWSIHnCTqLPtmTFZVGAcgQ2zg4MEj
BYrdoH3qtel9rh3yiE9PF+tHOgXkKkWWf2JY/ee58or8uLhugMUUZ/lQ+NF1
V5DPOjH5oAtNxHpP89yCvlmBv7mUZ74IlJNB6b1Gw/s13iqya9ZMgG2Rw4qJ
n+FXRMgQNzs3yN7MwsbSyVYxgTvcNPb1yZReEb7XV/SNb8Pi1anp/ZaDPCQQ
2WviALetUX85JOMgDCEdBBxtFnB2Q0R7o94W3jeNeJIQDO0JLCLl8d9hKxiE
tytYS/Pzas/umLT4Zoe7dZVHnwB9ZZW8qpN2xyhxVtbDsF2ocMDJ/qOqpafr
LQmgAX+8aLttp7kCJ/DVQ2Sc4yi8rDX2+DTehEWX9pNrkv0QOid5+k1qpHwV
Z77rC03hD2oUdQoBsLEX+AVIP14M84xjAgEquZLbMBhR+koAgsNOYgWZHsnm
cmkgOlrE0ZGGC32dl9O4xNvNySiFjPuI9ih3MRXieroGADq0BSiQIm4pLFcZ
jSqrzrjwZArw2aKdx1X6oUjCDJ7IqNiQyUikshYJypYhlaIhjjwCFZjeVUwS
KZXDY+sRmmLqAYAIE4nVtyRRxgGFooE3wwEdtRbK+nPzmn1ZfWW8c/PCPbNg
thHJYyUXEzYJTeQr10kF4wPobqp3dhhHU5b/5G4RSLMV5pxwNVGeFu9XQV1L
3CUGU0AF8HA4TTOApvsBVNLVy2rF5CJqRDEL6AMmbQ2aOuH9TUC+qidxdCBN
EWiEpO9ThhrggIjuyLCIB60Lu9dZLYUadaQTGIiBTto4ZpWJsVGWymWrdDkT
iUvrVhosLjSWqYehqDez1/SMd8hN14TaM8Pr5qTpTigLqddvzfA/LfvxnYN7
OfcfvMloo8Ltcchdamep4ZSp2g+spNeURkEbTrzn/m4fMIekKZ19XDeoOvp5
Zf8ULQDALxv/FKIV8wuBkpCuseH39QgxM7PD1T+9DGjzM/hqUODOlTGwGEWY
zTPFA1XCX7yQXhh94jJmQcZ7RobPwEHwEMvDowadBMx6d2k19IjSpVQd4NHF
6PSp0JoV4IUf+PSVk42WHQ6sSjfs3iNgHu64hHo5X/3NOfBq00jdtjwXQbbi
1bN9c2nYuZHSH4MVbWV99B56jSjx6Dq71wyyoTRZoil5H+XoNmDaQkdyq+hK
pX0yLOnoXNFQPYBUHY5denAn7mRU5lo8cC8BGC+IFJ4KH8amOxPJ2mlloAju
03wX0lHY6L0FiHdhG2I8rRB9bWao8+ugAhkWm0/B4U1Qj6ay8QABdTdz2e6o
uq080TZWlT+LvCTvT+/LwWHqh48h9Wi4szdYBNP32WmZCDLOfxMK+Y0NKw00
LROariI2h5T6b1zMWU5I5A4L2zhkKj2hitSw3yaN5zOq/8oIk2+z69TCR/pn
CidB0FGAoYqh3RFrV2jUWhVsVx5DfLfRTWFIq4hTijkESTnpg3JunVYSf4ic
dGrKSA5m5h2PBPuS30ImIXm/ykNvGOvInC2nnZ2PgZJ6rcH8yhrZCdQsFbhX
RrZ9FhDsBXgST3Z1sWb53caMetMg6e6pOK2xYW3qBQYlektVzp2n+bw5hJMX
pqxgbRTUgDiAsJ3Y+sZn/Wm2eEnUya1Hc1rNQ2kiwOk5oV1+DmjXSlyqYjB8
usVNZ+5YAtmuak4VwsY6ugTeyqkywx0ETrtXTOcgNbYRMp4J+H46ekUdX9dN
H4vrJvTy/q0Ebr67VNP1Ir3gprmRcqHHf0Zxvnh3yEHHDMx0LufWp0nKCUvH
sMtIGZQSCTYOqQ1YAuiOhjp64YC8qkv/M/Ps5IFbEsTT0mVqCQUDJgJAa3Ks
1sby1UG+TDLPxs+jGcgLOZZDv7VrnT75ogMInVZqXoKZNoqSUhfYM7EaUP6V
HXTbs4xj4FC4iN4FrECnyzPymmjs74tOaOyHynkRVFt7kxUWV/uUeabLVjVV
2oCz6qeYsDedHXE4uhe/u0WIU7OsGRtxnxS7mPh5HOoWUFEXfdXk1GH/Xpfh
VUxBn9aVR1gHler+QXgsCSXurLF0QNFOYGnzsBqRbW7AtkoHd7oGXlOEvS3w
mRLaWoM7rUS3pgQNLPQpmUgJrrF1YmByP3hDk+ABp9e3g4fGiFhmxh6TxvSv
kuYnZVLDSPp6xuz5vzosNAFtg+EsZPk79sfSc6Oq+kzAFk/M+RlInw8gtHEW
fSW0VOBsKtrVpQWm1EzrhGFFl11b4Bha24yMN2ug1Z/6lLK0Rd0THD6YUe79
XY/SuPG0PqrhHMPbt3fvN9G+Bh5AZ92bqu9CeUQJhuQUiLhKXYfqFXhi6JCR
mJr+3xVoEBFX2Vb1SwgbU+tmkuSy2mJfc4S9VdTCju2o+5hmCd+ty9oiZ+CU
FhWE1aLAo2166Je8FGk54cYjfxd449jF2q+aLLK/IfcpepHepUexTw5xOAHE
OJoUcple0Fd6f7Bg9I8FwmAAUMNnqh2XzcCn7kxzn8QAOpv/gK/9Ktq11nLl
EnLlq65qXNDTHQiODTPs3nGdqhOyqKVFNw2yRdHkGw9YNcxlNSxoVaeSoAxo
m1tnfeQJfA3x8Qbkn+alPaf2E/r+gSdhGYnFEUCh/7PUJggQWDfpyYKVNyW8
eitvVunNHX5Lk+C7fDc0GVFy0ryPctcLvtPvSs6zij280ngaGASvNJgdcIK1
jcwyuy14nOYwAV+4ucDyYABgws1+U+G+KJjejqCvCm3u0sQv9ca5sceABZtA
EUZXB3uAu19CuBoyPX3br6cqBo1ayVlwKHmeUBJ5HKs8ZWzyCuZ07n3sULTv
DKAgErAEMkJIkuLWaPodqKcuK+Elc+/sHN/f/OhRiNKpXq49PmS+H9RRiIhz
KHE9/Ikkj+YLZSW0UncdOIetP7AfBps1JYOfXoiSPY2T3rxe8/NYz/X0nLgB
joaXo+WonLKqnmeFdF7X4Qrt7WXtY+rYWDxCa5Q1WHCuSECgeoRjkV/ISCrK
HLjcpg+7OTiR7J/PMI7IWj0AzTECZy5E5/IVhYi5DM0GnXVM+5OFIDBeEtMQ
hbvAh6SQFFGANSMsLYP4NIIa9PDRMciSFzOqM7NjUtCNjQRwRkT6Ywt6bBMR
bcNzLIOD+qnl+DAgDOR+XJ+VKShxp5IK8gQ+XqHWaE7y0WfF8iAjNpQhGrJs
0qFnmtOvOvQPRNXwklglfExxRNHOB4U+Xtrlr8NBNA7WjsmY+pVCcKEAwcXS
JtdnfK5h6IlWxQ7Ew5o/WhZlfqm2DG9VTvbTKQo+OoD9A3avHdmqJcp0aMG8
z535bZlmlHY2hRDb8BbK8ZjwRwrh4RLJ5TLqv3vC9ydZSKG5lVk7JzuKkaw5
eUOOlYUSOLXvDQ8GT4HhsMOis4T5gNnKc28XBKjvl5GMeLqNC/20jfpsWKh8
vUPCDsWtMPOGt+vXenAZb8FwDTPnoe2P+zcJVwMPapPMtTsTY+i8NXP8xX/n
kLzcv3sfivnB4y6Q+DAAdaaKOUfUOnMFvHMEXGIPHPsf7AhmFG6a7FrpjMNU
jdPzVrsm9cP2bNkuX8njqkoqXE/Xh0PRUQB28jRqcGINsJg+MiA0Q4fWWpNU
E11KhbDdf+S4ZqF0NLgWuehxF12+t1ft0nb0I+StVhEb4RkV726a3CPND50y
28Mf8ewpzsqbsJrHS0Zq3m181SMFlmGsLghjPAL+Y/kA25WPZ3zZPOWffY6R
0q8Ms8Sr64pToTUe8QLFLFOJL88qGx+zJWMX01Xar88RPD3/21BvaDsyBN0F
lnyQmbQUtopHfyPbsFGa2KhYrkP59R0Lrs14FRYQPiMPZXoGwWschExp55kG
OLQfKed4YrgoPQ7tyNKq/8CtNpU+YxeMSsUZBMKZWzXj02JnudXZ3zI15cLP
hJuMNZ8U0Sciywx5IQhmiMGp8Iox+y5GebHV51gZK0v5fPJ3RDgh34JNtPs1
3hG0Nwt/JUsuuM+Fqq1TTNj/5yC0ph21TnKycmj45ToKR0JaK1z6KV5q1UeT
4f6mMitG3wTuri9M1BD0rQau8B2pGbvgqx2ZlVHQf1T3yGRXj1I+ojk0vIAG
2aQIHLQSfzaQiDNcwGnByIvfxTJwh0O8DPU/f4p0GTyCaT9Z0boN3emnL6jM
0TmR44tBeYFyfaZQshmRuO8N/APakMkGTDIrvecM1io6rHy5//Ga+nSdZHPo
OWsF81l0ppEGlSF2ehxbUGXq0pLBOeVl5JtyydoBkYpc8Gv6rad/cTUIW1R0
F3naHkod73acRIKNBU9z7fOFrkMrMy66mDrRiOtaVxrbXLfUpcsnBtVp2UNV
d/OdPDPf200v5eeAxHF2R7r65Xbm9owpgHtSS8kguKMY3h+KJ91C/SujY60m
T89xn9QWe+VSn17ah9N6PU4H0vVFN3nkTkNcVUVdi2w730DvooN7gDFj6xPZ
dXOb3qSxOF0VyyMQxtd/EVtqU4tVnS2WCv0WDCjFXI7rR8hFXpYIQDvRK1bX
8zUcG6qr4MfdOFt3zOV43yo+5t6+VKYC0nNaq8okBxdtUjG9rUMqHtPF2y8a
HyX7cpTVMQ4fa6JtWfqOUXyGL4+e6c4S+uYNuTLFiMpsxZ6/d7HiX5+1Q/++
MPJfBxUuUagFgipiGualCipufxqeCdivqJq/++aO8W/fTN/1Q/BXN9Zs5qAw
D2QkyC+BnOTlv3h7zxV81Wbvq9v6Qk9TtGZPK25dYQ0X2v4IjMczUY/gpAsm
q9v+53+TfOQiEOtLrVDxZ6SZLLJM0OxwxgD/2hxDZmiqssw7DwW2BP2VBQB/
ymNPpDcvfVlbXE1S6n0wcECySpX7Kzh8XiZjthdpaVDto+4aXk2T0UVE/isP
kh4eHrzWv5ruE3oxHddVXMj6PY0HlI0xZqGacWOBGqZZ1Y4NjY1G4ZmCCU9q
hfvYFvIwq3m70fqOSq92SKBPwUJ8V3tncKjdZwX0n0OmjuJriWaspDb7PG91
BauC+XOU2SXUN/38x9d0B9TmPNMJDFZVZ6+IDijBZ4PvQGdepmcLCBc8pxHf
J022cW+sx2olpD4uiRGZa2kPOnhwF0QlkcFcIdp5eUXQZ2dmcauG2+pKVU9u
bUISMJD0L+TPXrXh2yxLbT0vhlGZl7u5zFj5rqNqjWTJZmpCc0tY6XQ1SjmL
bGlaZ1gjZ3q2V1X3jVp4f3EjDL7aBHGndtkRC1s2GsfgTnwO9jV00pNYJgOQ
BDY+FsYIvTbDydS/fG3H0zoDpndUN0pKIMo96EquIcO6zAJn9qn5i/S3icBR
iSHIqLSlCViKmCTyEn9mk7UAhGlS/o7oOSv+LpasGRnfs4lvnW/j342N86dn
L2T5V3xth7rSfWupHhN7Jf0U6I+np56AxxzRIkLLR6L4vuXTY7n1pqFQSOdF
Cn5jYNpz6zuf4EuJNsrxnUzIbWsTS1bHaO1LaK+VAhxgyVEGNzbrn9P8I0Nt
4eIyK6qG3422sgejH3h12r+CE/pjl5YXy/sZbfD4t5oxY7+gij2r/tttdoIJ
n+RAy1nN8QFo37gbDjuIUHReE+SS+Z9SlJkp4AxLjBJNMbzhyKX3EqMsbVkU
WNKNul8R7Bu1UcP2XS9vYe/xapmUbCdiRnBKi/C1/7yTiTjwJUYMRIphSKS+
/i27EceN1yOU4xhVrj3alD1mWeMLeWxKtwCu6v7SpqTXr0TnCQNpNsBdOIfP
0CHeh0EI2qCW5inHcvLNMLbtpepInLHObRTL3clABYH0e1WUAsD/CKF9bYZa
3yvPv4obX+/66xyOZ2ps545TKWKNGeV0Xy7+ZzuXhHnPPurYaS80gf3Lom2B
nW5i1ojVXN093qyExUpRz8VYxVu6a0pWRWdbRvI8lqsr32JyWnu9TIxxEoRS
1cm1g+fJhoqd0xyX6KEcOsZoAqz6khNs6bMynsFyS+Ehv4TNeMAYvG+wvIWb
ghcjJj6VenST7KD6+niH+QB7ez7zxpJDNn4G0G+bKCsEShrnEFndOB9FIFRA
vF5NtJznr0sIiZBQCzLfjGGw7+kwAmujL0Igz4dQBs0EFAqukaIqHtlXXDiI
5Qj5JLrokxM0+L1RZtPRGQ6H4IGBzg2T8LVkUCHkZGpX8ec7NnuwAtuAUA8m
IdUQO1Xss/4Kn+L+DjN7u4n8fnyTnXpc9+HMjS6wHjLgFN9mIdMRAynEcx/b
BXXFJJ8fH8h8FQ+xPv3aqLEn8W3jKWRo6aAQjiqhDZBkS7dSsH/rB19BezLP
yWkP8hBVPzMK6geB6Tv+hbTZNPUkOjfGcr5Ds8zKts5/Z1ygIEjFiHyR/Ly7
dL0N6tntK2k96mDoZavJCEYgSu/cVBCy+P9Ms1jlBJekgJXfBSIoNnrIzpei
t7zigD1cd/Z1tUGJbP5e+FBKkNKrSWN6QditinX3rkrPqCtR0ZUrv85erUql
lZgh1H98/hW6pi0W0TdZL/SiYtfrUa3Q22j8ax5ai4hjZmHs8IQerNaQRJ6k
41MQHf4yZkzjr1BhviiqIYTAvIMP3Odazy/wSTd3IZ9Nygi/LL6cttfPzxY8
Hwni6om5q8byKjTTllY4jLRIBMk+U852+wtDrCShHu6ow2K2Tce0+ZEziJcr
E2gY4duFoju2EvO/J2cq2t+RYv/cQsI1q9MX8v7qpxdTbrleikBMOBMa7T+G
zUr5KM39rjb7Tnv7p4BIPWcd1KUFpOzLLPo3BnCvdvNMkJqbBkAGUztqjede
D9cn3DNqz8FJCqr39/fkcp5rleNYvBAg9BhWt0MzOrkJQFrl/Tm8Gkp/l5N8
lYIDrafty2i2UMN2yTmSXnSA+VmRFp4VcML/oj++tC3GWzHWaqIiy5/GERrl
mBwa6HjqGlhNqnX/v6CcMvsd7yrqdTBAcFjBJGk08IAPgj+I/CkQT+BCMbm4
4h7MOLMlzLoVhwqtwmyabllGXv9AzDgwx1qNC/Wf+wDBzZbJ1lXMIvj97nvY
pl565/l8dXowhnCd/zNwOwBCEECOiX48r7/h5lpFb1ewDd4OMGefPgTQqywF
EAWIoNYZwf2rbR3DdoLCxG6RZKNKV6fhyhqM44TlDwkqhBLfsqfpsvFWkhZW
LogSj3CtDvIsCBkh4z1athgav4qM8CIi8G7CcKUzwE9kclsecRhtnUA1k2Wx
mSmAe3dNlY41MnUYaWa+M+TudcjhZ10xQaN6MQdjbUgAGibwvV5tfspGAZfi
Kvkz4OtOFryIHgCov1lTvPBfGp4wSapmLXB4IDe0a7N9hEUinnv1OPLwE3j/
RO1OIXUaxleIOIitR4Hq7Pd8stJSwpKFixpxfc7T3xgqhk5nb2n9tDHGXRB7
99GN4h8JtGNX+gvSF1zcBiY7lwgCrX5mLTAMp85ukjO482HQrYIyQJoWMIoc
uNkoHswkucRnOl0L+7FPalJlhV8A5+Zx9pXHBzknnAKA83QuRAb1qVGGkV+c
1zocf0PpItvHjy8lobP2e1S3ja5kcbaolefNPWTod9PdRRGQTcDvxQhGXcTM
Zb77L50vNo9pGKaEFprKsGJmJ+Wkd6JaGhEpW1HuLjaZ3kgMqXoVr6obwYPX
bMruiVsPE2PLYtP0+Z60fsv+/csWsJHF6j7nNpwNPxconWT7TPwgp+jA0lba
s33gyKkC9Oe5NnavsP5yaJvKlpynZGqyD3k0sAeCfS64/za0w0gaIK+pWHzE
dmt7F9kT8YBgpKuCVturFYvKE9DVyINDUpfYA07MBqBYmY7/AQCI2bKFqsfL
XTXRRO5Xyq+5f2rA6s3PCrzXoykNcuKP4mraQWgq6m9Y2JB78bRmQW8jKdsC
e8Y9JGBMHENXdCQWvnYlDb4yuzTUcf3hqgcvT8NiyOFvMXgurjEZs9cAJASW
8pZ5LFbwq/goAuJWsfJlS1k00HImGKFECYkhwl7eNY2nm0//r2rsdECShtzk
Iu4abGx5klRHS9DG8LAHSWFdtJe9YGUnkLjM+aptjpyeveaLIaRSwG3+BuSA
ALeSapQ3Tc1nnfq1WQum8xbXMbExBkUJsLNh/1eMXQEWad46XS+6nDTV/Lyx
BxvqFQT8ylAr3WE5hSapMeW8eej8ZuTc7MS4/oxY97SOVCUMaUq5hQ2wxNO6
m8q2q/6QX5R5wJR+vE0uFbzz6Y7FBmAz6yVc+F/klQ/5x1l/HjtZ8UYyXFap
HJeX3QeFs1TjWb6CkjcY8OV8A+ZTiH03HLV3nGeeSlOL4SztDQaOwbwlRZqY
lYu1T9Wp4T6UM2XFaBtH5C7Fd0blh3InSkFC5WfxdFNsGe8yYPXvlUpExjF8
KM7SUjPHvSkHKu7l75j3AxVhA/8sRyiQdwQsL7IiFZFvHuWl+KpNzzvKnsfg
K3exBjTexCWOODUqBSZHHtVzOUpkLPxox+cLRZhJm/fdbmN9jGRzo63te6dd
fWz7KZwnAKFHAjyP4hUgk8cVzbLfnI1VDUqOl4FpvpHGedY3foyznd2/TNKo
rD0nLjkPUW1BXA4YEvlq1gEwFoswryrME1jJYF+NlQJ0l+obBR07eoYVP/S6
BDaRpn8JE3f1Xs62Q0PKwPBi9tGSUReJvEwuA+qEkLR2XgdccRfSdkaAdiCZ
yh45fM4bmyACkW/ti1TjvrYBXn4Cv7NH2GC7C4M5Aaio3/8OqIdplHpU2OdX
bUgloZySTXfZnl7WkV7Yc+5ILz6t5EnwxaJZ72x5aLE9wU0Y1EAjDi2XBHko
26fW22kuuF7ExIQqAI3ermf+ndLJP1D3WXOH4SdongQ5c5IUgsHFTmv/i4UD
L4Vv08o2/SFACh4qWYb539kjL/DnS8EWJR0e58wPwqKXGxFlhZ3OQdTR2a/h
9jzJXZtun5fFZEqUA4I6E7SmIkKNC/AB5Rh3UBSL5Mfh73KG8SXREIw/+Q0n
/W9hjQh7LA8j1nArGG2IrbSw7Em/XHz8aLuojXRPSWHjQezqpHrsczBvlbYe
A1gteqm8lo3mTRPnRD1ltKFWAZGeY2BOrH3SjAAAjkwNGyLeAwvDBuy1ibgK
FQ+Pq/4Dschfbh7VoIkJ4vRoBnXt6vpl5yeFugP4ZKDvV+E4BaPGj+izK1mS
l3YZEqxK05VauZ4hJeXmRZrBtXCoPPEd6cdsQx3oT1bK0PmSasC617qj4UIU
X3hV3fphovS2Z57J+4rfeFzcaV0CuFchyaqDUDEjwW3sorX06apM8JqWwK2Q
tZb3VrrWATr4kXuBsp+P0585Jm/rU+kiEI+S1wcxhpo2XWJMUqFiX+npiNaw
qkzm/14vEaZTfrCG8/SLzNAfKRE+E3tZphs78ztmRGkdps/J6P8BbWLYOD0e
zcqbgUQFHWtezPamFr497saD2faa6RPwD4ZchVeSEGRMW9Hn99alwG3jpYQ+
cyUuh6fa1//ecgMmjRCRqMwprxLJLTAWAbqI9fqwI9OqDWRJTEaXO6TWMlTM
e3nop7THNzcoNDj+2kXxEKQsQfRbyMuk17chv7xH2gvBCvGzorxS/lyCF1cO
WhHD4D1l4f+a06hIJmTaj9uLGw5IqPXyod3DaVEtUmVFTZfGpRz6fEdCD0+G
tPwkfWL57q6wk6u1J/M0rp6FREj6jLeAaYqAZbe+RNiuz5+t/tWZyviZYPSY
zyQIZrBNyUeAN4TPlaV00HMiudxZpY6bLfY0/i3eNppvnWXT7JBwJnTrBut6
vXKBkQrbzpsF2BEl1Gk0IFjuxepiMTUbG09VuB8nL9V8wJCBHp/x15wAo3/k
R5eMJY9X8sQpsSYhVUwC/d73Q0K0QzY8Iw8ePN7QWZDD9ZyLyHQoWtdlvz6G
J2bHWzU/n4bRQgvHW5ZbVlQ7tGJLIGECTbWhLHmwk2h/+u1OU6pxL2e9YutD
MQ0o/45aCEcTPOAIaBvHq0tpPMreuBOhANbbUVPT/KMO0a5TzJ+AyBhaYIHt
1t9YbjMED/7XzomkM0ocT80NXKDTJGf3Mqyl3IUBDIw2wdXAYXBZrqO8NdsR
gHJg7PsA1TulC72kGpWvIcXbAolrxJkdnagscs85Emj5yyxc4ZJ6jD3G/Zj1
lp4dGMfwOE3G1FmigjVCEudt3s1G5rGu+8Ai7eYrtJqXxwFy2OHAjbkmyZ3f
ezdu+UFyZAQsmPtWXLALZnTUTMKjs1QDmY7WR1y26G6rY/gc0vqF9gMl3nwQ
nlhRcy36m5gZ3OhkS6DrAxcFCtwoqBq9twk29P5cMjcgCIPvBMu1xujdmuPc
5X7cb/0QHXL29FDBQU3bq7JHQAtVuz4Hph8R0mtOnTX973Ix77yQY0srhK/6
H2orpJ9JzN/JOwz0fjAQ0bcHpq2nX8Bayh+NwczFVhfwWVa9XfoRvblUE9Va
gnh5ihTauyAjOs50G2GZuJVtsnGM2+WBlyJ7cCEoNsrQlI0mxJoTS1cbvFLE
AEnZM5PHDGIyoTi9ciq0aeBJk5/EDhU55ie+cZuk5IhIFtwvK7JTBdQy2VG1
7DOsM1iBKxqRWV0lRRJJVVlsdY7Z/CVXU/xjwwhvpjxzKJnInNtreTQzJjzc
mUJfHfsuvUunnEVhqwa7nHStL9BDTVDKl5dsDOXJyy5XVtb8r/8wt1w8Meny
8Ax29gnQeP0GN0iexnH+mI7qRsNu2BJblCJ9521Wg5uuRA2l/qPHwM0UT9gb
XC6Gcc/uM3eTH1oWsEMLCMRqOiJDa5ltU68WZdOvu4Y34gMuhMvUzaREiwkt
DugEixMC/Qp/1S3mNmKE5SUs90BjPqQkWjOciAwxYqezc01kUKD85WM8qWBq
c/uzAPky9hnELQv4DPYB095+WBPIwVjGQHLZ5fFRJeLmG3xR9NneN3loUGTL
/yEGgR1CmajJJatLGBTJerDd65jBAjfrfiYuIXr5hLJS4YaYRWF5OekiIvww
qdmsA+2qWYtqS82ySGeQ2ooLr0pF9uURZA1xOxU1SXj93wKqWt5UT4HK2dft
oH0ZnpzujU4Rn5JwatD4PVYyCEkBmtsfhVmNNIJ55Ka6jsVaN4DTwMdzS9To
pgzFWumIgOElWd7gxzJgMd67TfR+Uisc6gZmjrwyjtFd7GqIeFnK98+nmPaK
Z7mBK/3DzTWvWAG8Dl9qYm1+eTHOK8KVAaSNXlXOVpehHXUn70jUdhnnYUqd
2QCJJVm9PnLZYQ4r7iHwiQISw/4ZUuaUn91KhtCAMMxFngWZDWIncGiq9/bj
6s/OxQLpAz8vJSvI3Vxk1v95zUIKMB7623y56pcI+iKODKSb3BnNzXNXb8gV
u2X1QKqSLkJmqOoxPSSh6ddRGwkr2soF1PGQv5DfcPiHrAWbC07YazFqNAf+
3E/g8RCRf6+DtUjn6ewl5ljCmX0hdzQdyNGC1aCMBbtqP3uLI/LHNv4LJmue
pe8q2DCqKDqdpVpTPhywGnhEirNBtle9yVZIb8K3yJiJgtqOdpSnLMawNhaU
pFBeAeL2HWePbPaNTw1zHY9TlzKm+hgb9zhZfz6s6ODVPwfntxW2VnHTgAgR
FBLXPdoxJy2/N4gOY+v5BVgnxbbm16yJj4Lnxuu9zj1sU+ugeSrdII4eXxdR
I8/QePQIcXS3ia7fRaUeqXy6mf7LonittkkvTwfcAT74hgS4lyCbxDEQ/wua
HfZzPRVdLubWVtkLooxbfQ+UxqUunmREL8cgEW78q5zL7+guW16PtXW8xF5N
pRRdGUuBXpwvrOKJpnxGj0RpwRoa9iuyY2cNAPCX5tbsrgGDP/wFbm32X9PP
QtYqa6Hlr64QZ+fVyGxT8qLhhIpGIQ49Mj00LCyaDi3ec6yonUuu/04IvMYV
tW4xS01T0W4e0aKeh2DMrrjN6ftEwfkg78gerIpgc/9fg0x5he4VdPsBEjJM
cAtTs5MVTj7Q7d2RaICAu92CURR76kAyZ+CVBSuJh6N+jlSrnw+ahlnYsxwF
2QfaeOVLVZ5K2qAhD3JkBLLEIIKb3xe0m+Vv+RcmFYArmmHHQSPBa46brX3n
f7J2A2SBgOrKDtIegNpLabgkUr5d0jZLXjizPpoCRaHOfKIFRde++ZzgmmxT
QVgXKaXAgWyximgqNrzJfkBGFyAALEkQnwHbbTaR+fTsAfUc0QoRdcKE07sV
7wdkbCtP6gy+YPYtphKjRro/JV+G/gPAsSZIzAn4aqFLlafWZsYHAenfQigk
qlK19/mGbgVdrAFJZMuF97vXxARQD5p45MIsc5VitcqN+ibAh2VLkEB94moI
GTi0gENn1vH4ItT5TiMSgUMeTm487aCR7A+SXTRA7KizczUzBJlfegvl9e0u
OG8ndgndhkJW/LCBinkg/jpvuFkBQTv6Lnl6Ue7wYWjULdF1WRTWJAgqEEbM
/a4PUoaorq6M56xl0BDq/2nClWMlVdIbz4wSgfaodQ/5FgnafL/lfYZ1LLXQ
Iq3keX2DJNX36xz/6wDiBj7pUASw3UEhxZT6wZx+VGc0dzUnJFFsZhTekvNQ
b6wd0T3McdhWGb00yv+URRcfLPWnXrAqOoKekVri0QeZh1492/0F5FpIPlji
UgN0zq6NmZD27SXqq24jwCh3XiLGWJ1f0/gQ/WJDCRzjh6lKI/+ZCTLCwyl4
uBkimd0LeAmGlybWFTXB/xMf37Oj68y+IbCaGmgpGqN7e3IciUIbkBcKUZSs
H+QreqPI5QuyKSndUrNgdDVWZHCk38rTTA9tmYwL/Wia7A36cx0grQYMo4Po
r1patCSlZW3X7NfZ2gu9QzDy9CIjJuKfWctg6aaKjs/W0vQbOIg/qzzwwLJp
TYJabdwiKFZIhMJ8k+A3zYN7LyEqx1mKxxUBD2BKXmQZVwjNhqnWPe3Gdbki
XVmJh8qrNFjCWjaduKAUuAqus2G2UEA183de+oAIjzTp+sxB9VfwqO6RmPhu
2LsFQ5T2Mk0lEjLfkuy0CwV1JobYoVn5iFq7OTKbgMupKx/Kgk69hlMQZJYl
fRQUyPSYA0PHY/+fQc177w1t1ijqF+r1Q3X1G3bvRtrFN7sVt8PTVNJudZuk
Movg3wO9z8CjBzai2z1YyD/nEiMZl0HNvZtruCEjqujQzJRyQmLKDDdbGDup
bZmCnSNDmRywS30chtspz0jiWdr2GmHlzjg108pO8qCkaU83ikZTWQYNbUec
EABYcwrCnmfU6jKtkHpA6bgNGQ80/bXrVUvAH5BJ8LhZ4QqEXzg0I8oH3xim
9lh9wKNwWgXR/Um168a9DoKuhm38SRk8Y8q34VlYxsJt2ky6Szh3748lUjHc
u3OtpzX3gBym9MH1/brVwswFJEHm4l83IHd7XqF/2cYPVB6WhEcXGwU1Jd7s
RcrOzdWz3/pm8x4RxF0EL2o7YXSRgxpnKY4yxnOUUcssBnaa0Ma/cQk/sSIc
1rXqVWHW2qqe2ck5ftIOR3H5JuNBEzixsKznP7lSk5J0UuA1g8BCn0qWDVNJ
yR9XIWrIelAO8eWn3SFnhnuFczvBW3FPH/2LIi1YUt0emYVakyBO1RYEbaF0
vLohd6NQ0Qv9kBxjxyMjYNRZJaJqKJZo5KqfahuDdBFmNfjewJ7Rrf3MCji2
dmd7zqFirX5lWCd7lb01kteYBzxvhbfUSlggWh4+Yz0zt2bAeU6KuOtVThsu
4s8RyuS5OD53BWd5ozQcqWLifFYNcCaN4D5mFuMWtjAuTRK1zohBOQxfZakQ
riJeKF1tRCEVTxCbUR0yBJujWqwwvY9M42CyTS+p2upkokpCv+08WY24SVKS
qru9LOBP0hamVzzDR5KqTfAAeF71bi4Gknz3uZbdoW6VGA8yzJ9uslme9Evn
Jo0cJXSglwA+w1KBlELU6+oA+UzThNoOjXMl3A3ZkoU5NS5KnOVf9fFDq1UT
TeFs0e5b/oPYuI8JnSBiVCitJfSAugoLUOgHH7+rZDfcn4Kyj9WKZYidAgpj
xrUxNWytfGF0Q22lKlnypYI0rE6Afi4evfkJQpCZKGk4KlrcjAlJQPqUtWNr
euMSGBidsdM8yDCTRzXRBa5OceMbJTDmTw9hMEcDq2lBI7AP1de5H8HMtRMu
hVk0VtrPYXMozPTI484zj+gCBpPazENgGWHSQ92mkLYBZeX1G9lrUDG/3lFd
KgLLiaycZosqoPg7ROfuQHuQc9GE2bC2LlvqWSNZhnfkQv5vaCiJf3O9Za38
8dPhBNgK+EToz1sCqJjKO6p261WRUTMqGjv26h2AAsFI41U6xbSK7r0slFwK
jmpyUv4hnPI2dpohAy0g/slZrEo4Ih/0AZuz7yW5r/Oipr+xArYV/o2pPZdc
m8LiwWRgLBGAWkYgrv7gef/WCtn8f/0sHKqYwKHPmwjUrq8zMJl4/Uw9+ugu
RAfq4nsBj36MjppSRz51kvtXNpyk8ZHLLLUXuYrLHnsv0/n166XZK5pZALkZ
wSndS7ZOX15xX7+BsOrerBl6vTFbmxIcUjuCKEvsvYamvgfAcdNzK/butv+0
2vvAccOj1yC/2lM+DeNgG6+A+fP/39aqCQJE/qNTjx3Hi779KOdYJAGLtZI0
Y25rGptnzqCnv+sZfmzm4ZYhiip21sozjrVXror0YAJeQVDZe4hWTEXTGreH
XMnXsrBCkt3AUh8ktj1uZ/WfZcfsDlWKcQ9pdbHzDH0KtEsjAmxHmDsi7n5S
df0H4Rd0J5NDaWuC9Lreo6N/kiGk+bgUWDnRRUe2V6to23lrOpiS98wjFsZo
UieldQoxBLsWYUT/Fvp0Sg7KwNoM93jHj9SHquHAL4KmTxD8qnjr/Udfzb1Y
j9UAcroU5czsbllyis/sl9tqh81yMc0r2K2pvSQXJtGV8A/qE/LJv2Tl/RN+
vCkrT3Y7Yf1ohOMzNWW+8FRBFUk8zypvWluVscTMD/e65WpiGojE+6M1s96A
wIDhNgZ8Nld+MZKtRqVr0IA/SobBs78MGU1FR4clnyFpNNeMxSG5GoE67FV/
FqywJBjFKNSmoonVSvFByysbh6FpCX+N6ywhjXlLlBu/da3xb9pfr2e98B7L
D5J3Ndiz8uXadSYsh+WzzUfhe3NRpxQ/sCC90A5q5yl8oYRLFVILSI7UvzNu
+XGTQgToiSSmuvchoRKrqGFHy6tiybLVslh6IGlwR1jiPq2HitqTyEXm1ftd
8/bNlzAwqQV9QikgjSECvHvLpz8B6cuk1NeKMrxC30YPDBkF1PfI/V39S+fb
jDNJQv3dCMJbjxpc3aqrTmCRv2NpuGKJJefSiFZ8gsXBR5QuDRLtvjTVlpEy
Bdi9pfZLaEEj0OzVGacoWCxSmEVI/6+/0rycr0DivCgPQZXDFWbZiHDmUxtm
VJSr2ROJ7goh4gcIyrEc2Doci9orRMLpdiHBISXcRxNz//FxAiGZj30WavIp
S6ofMlVTfhpNtLDAH1Od5crcYC1JkdZ0NhKFxnHolq9sR7pBP+EOn+d5+HlP
HzPTSdr/fT5fyJYl5m3ZgyBv7Kqcv8IwibeEhnMbFtLqLQgA/RxSp7+Fnyi8
+AxlGKQnrW1pSCice/PLzZpvMyAtAorUNiiq1/B9qmVin1OjhIFA6qKAmDdI
35SOLsDtHOtrtcokQ08RljhLtJ8SrPRRSpoaeCuBG55m3NintmSGBtLJ0tC0
gsk/orXE+CVbyFqg41tFueIDOl2Vnx7sricfNrM+LyhSezdWDE88xyo8X/Tb
6zpG5Lz5xnkQLh9iMuh5HB/NlwIoGwMv3x3aegAu++/IDc+M6bfqp3o+e1Sl
3uFzvdCWP1w04JVNE5gvawVQHCAqj0iK0uc3v73iEqdyiyKGs+hqf989yNl7
mHNz29CJN3o5T6CnMPSHwr6KRekkaF00uyZ+3tEDDC80eaTHASwwW0Tc5GPz
qM7VwVzAdOtvNCOT1hiQC5/R3EWvCTGbDmx0Pr3bTgheJ5Cgki6tqc22Hc6D
AxoWYaO7tczaI0Tb+KO6V2J8clyksVB0vNu4Mc77ekyxTFOIQRn9/sgdBxMl
SGzEElLiXRgMCtXB+/IH8VGfOas9lvd6A27gkHoPStlDCKUlckF4FjPOXTv6
Osc1r+HNvqB9pe6jGKMddndaUSSOEgfx3jLcfihh89eOe4UHwJMzrF+085Ct
m1YBk/J3a3HE2MFuqCToL6iKgmSDcyL2r+Ts9zBurnVHW1+vror5f4KT4DIt
FtzMYpRyFuMfuj9jNNBVNb26a+aom6TWmPTxNCxBWJDpWHeAtfTH+7864sIq
7AbvdQ0Vxdw21hhSjWKCPRchbi4H3QKa9OOF5RcsTiDTJ1iqbBTgGIzS4XJS
PHGRGk7R4nxGlX7rBj1CHFxg/OLy3u7smlDm3gyIIxsF/c4/hFmMDyFdZ5Gw
LYzwAkf1CFfJXw0k2QSyPyf1vB+UMxx/Hmz2HUunIV+gYxZ8lsEMmaW9wXOv
XabTBV1Ooi5U19C7cKK/62NG4AFu6Hi6tg45LS2lfHje1lf+JJ04ldcKrlDL
UVWGtiLk+hNTRP7x3odI64jSRtE9DusbKHBgSEA34QjcM5wr3YzXoucM2+Ad
T0CWNgnGxK1QB4uzEwZJEQTtrAtr5NEtFgyCdWwHz88kvrSciVbQKR56IFQR
ESHvU+L6CZN6W/EgfQzKUxu4hTVqAc/xMIwTVSO3Pto0JR+9YA7CaiBbPLyJ
ONUhRHltVj/XWLajQKKabQJeZXGKpWLbowQXiPhnFo7d4EJX7H+J62pNSRiS
EIUWFbac//Fmw+jQq8mPfxSBJ+cCKZqoIry7RPwEQFpMgZIJbZRo1C4Ub6YH
kx8JbiGxhA5oe/OVZS+1m9Qi6OrdipfGV2bAjn6vT5ikYsTMkWstB6To/iZy
e3taW2tlnoV3syso1fewg471Bu6eLoztxYvx8LCl4b5bXtyaHxDQKD1+3i3N
6PI1LhkUShH19neQztj1fYNl0IHlD6A9OIKRNxBpdvbCXRYSc86ZVvgX2NsX
saNO/VouxIBNDxBm2hc+F2LwRtUJtVQ9jHtXvJXUmyDvUSPaMRKUg1UlQCpA
nu1tHLW/+6LoZ30p6lGMpL2T+jfow5NlpSPbseY3YqLVbhnmiXRSzfl++xPd
RzbO67wI+c57kxwEBWH6jczAQs3+mHKnG09+U92jZ4tKKqLJ0zVRV5oCpwpc
37ltAB0SM5u86bWpnwvIPSnHL0fH5AxslE2MA3VtBaJomI1j72TuDx28BLNt
Wv0ws1A8KCecSkP2UUKoQNfm+HV427E7WQC9IANQmVszRz89OefkM7YcD1Gc
jNjpzoIOPSIIPpijMOiQiSc7PwTHw0ZQHy97Z4bRYWnNCPoPBkAi7XKd6j7R
R2EySZ5M7XYru/BTSWEV8hMDznK7vcnmFHCpWmFdz0Nkczca8tNdDX71qqPe
teav3PlcS9SgYPrmZoKHSks6ai71oIjf5ONM2h3ZfGpzkfIXBD2nQTl0evd6
vbliTeAokB6Cutf0i6thDeMYIvXiCpDMFSO+Wx9Jke3XQp0tLMj8KAq60C0T
9SInQRo9u9JY1ddY+VXvPTrV30fSbVXldV8ubLmYA/vaJyHBT6JH15LQxqRg
XK3i8u+RmebfNSMTJK1x0zBk6dQDzb5z1jLo5sxM6GVjsx4+7dbxY8EpJ1Jl
1vLLIbFCmqLkPz6EBCM7uRUlqSDlbJRYV1FjloRlap16a+WYQel+0VUHqyic
WU5rsVFpGkjxKCXpFVono8TRWsEEbBNx27SGkmy4CCqii4KopsEdiy98Z5hn
gtX0YI9k5zlKgEh0+B7qgI8iLRCddbOG5gClWJDBpZl6s4paUsiJmre9A67O
puDdUqfto17UW4wYGRjA+MqL6UkU6GmNoNlmZdkX0St0ce+9JggVidBOyFbt
qKZqLyt1BTQ3P5OE5RwwHDsi1l4ml2mueyUWlrsVT/AoMMoCbo4V4UCBzQ80
/XjaciALcCwTE+CyMyjJhCW8gtGiOKTnviEROKXcaF/26q751UUIsQ3XTb94
GG26hDznB5vb/ON/Nv0+JSneXI7PcBy+5dFBpe/F0X5N7L+8y+HqqFnCCObZ
N03xMwc0HxAapxtTji/JZ1a4M+r/Tg1u5c/SyJtGzL/Ie7AZ7ML6jj5zmX/3
6Ztt1NUVUiy9nXVRRKzbTWbTsGZusEatP4KX9HOvZX0/XZEx0t8GibhaTkOZ
z0yNWL1T8V6WfDax2M4WoO8oyG0wWKenszCdv3yO6csQiH4BWJxv5jvbyPG9
yWx+b6lILYoLW3VE3ulu3AymtTMvLb6Xv/FMmKCNXgjYICkbCzN72riaHxnF
qokigYEIFmtzhZd221BEfO30ffD/zanO4t2Vklku4YDuBmW/vs3BR/F1WE07
WvxRuiNUceRdYeO5mt5DKJrpp3lc7N7Sh63EgUtNALe4hDWJO+A7CgdV6DD3
ZGZGVu7dNgYk0SwFPD+H3xPOyQQlgcyQJICwl25o/1fG78B2tZJMmWYqbkn4
nde59I/JQ3EP2ekaWw9z89PU3s2nGyDnn2nMOE4lZRERuo3+S7M9bdXJYmMi
U7PZPRFJA3RvC/4sCWDktNDdPqnVZhskIkApbCCsSvlEeBxrdTORgSTITH9N
IX8LJlAv48EDcr9JqVvA9y976S4VVXBw0r7LEosUvi/T99R/Ke3czeDCPdZ+
oWBOnM0mHutWmxXA29RDjUnXFVAYLABQOao5KVNA1dLnBOkjtOXAXX2Gy/fJ
5VvSk1nyQF3AMssX+oxDMlCCjV5hQWVyzSqCEfZyormnXsVaWfUcYWlHVoNS
We+irWA2GtEEVTeAbFbAr+x0iOcVSwvm11H5eq0h5JBGLHSPiNm25v1EVviL
ORZ8gk+4WfXgtOB+1Twh5n0Aq7LJIrWIqrQwIyipqnmTKoqDlvaMFHItrZHU
jUM1wkYOE+KqZMwoCYApZlDNXfae2u3E7w7k8fbD6r9n/zXdWq9WXqpILds9
jFlmCtceWcRkOJ/W1n1Y+6dd52UH75Z4/Njl068W248iCNbUdHSfltuCBDh3
/Y1dgXmjueYdSnGWWNnjSCMKddKrXiRpyCx7QvGdYq5OYUAbssxXDg7Km6BP
44cBdxwRKNI2B5yqWxWKGNAcKvQA99UENrW5te0s1fRigIVJ9v9HVWNMe3uz
Bc8CXZoxPtMQeHPe1oVhDZf5G8v/lT605A6VbX1ZRhtnMM2GcXtfRhHHjJrL
up9VbIktKyEGz8JmgzPac9cfXpE8RrJqvzSOwDtmkW+jyUc4NCKI9qxq+3+w
jg0JJzZfw5ayoxweW87PnpUi7hWfgm2YeD7A9byr0Mq09DAzyK2cKTSmxQlG
fuLaStgUdjPVp39NQtwKuBWCeREvz3sGvVJrgrFBsqVxifPxmEW8mLrZ+pJt
VAKCYED/cWbuKg+GQ0ULtJmuuPiVisoXXRt7venTvZw7Voz0xnbhkUZktUhf
JRx4VPyA+RXFN2W3iCRyD4tktFHLssDcF5I+0AWV/nzQV942CUbV9xzBUXfL
19MkWzAEvbs07sM+46b8dM3DJrXHVTRj5/fnQHVs/a3QEobAW5HVtcwW9+fK
sF0jta2o+po1UsawZ0l2TF7BBG07jT7cT42PQfvXI7q10JXCZBTFa0E43o7J
qP7D6Sm7I9D72LxT02idiB9rl9iEEOYZeerYPSfaRYedjNxzmWuLFPFAkiBq
w8/7fIgLZOJEe6goxqxKQLw/7RbF56mz1KdZE6rRigvCeQ8N3eJYy8an1t+d
wywJbh1szXktN9QVb7v/3WC5Yj+b8P8M1xg+G1R+QMZgt3AUCl3o8i+u6I95
TRB7dtzLzc0KNjZYHMah+eRSzmaqMWbrz1bSFH0W52bZcKtb0RKpXfH5lk22
nSdKQiLYzry3/uJcRh6lurfzXYx12Y0zpjQ/XQRTiPp/nDanCOwB5HD3vAPc
rbaI1eAuqu9Pb8RTQGNKftnaIVm64aJGeu1D4CjEk4Uo75U2QNpF2mraVuQj
JfkHV1XIpkQxmTNzhJhosoXCiFIfZAfJbEXoAHOJQfkT8YAFjKnEPEcN802d
9cgoXI51sQaSItonOIl2xeTr32UWSLnLrY8rzpzwf/2Ugm+dakmx+Rd1WJqL
cyD7cL9ewDak4NjRwsVb3CtIS2wSXTkPuku4iL0uH7S32c6Us+hfwSkJjKIv
gTk52U9k4iBfI7tiOci5TeDucOEhDyjrLqYRFXb30stcdK6+sePpC10XskP9
tLUWBWyrIf4kl09Gd4nmmBNmBfEI6yGn1bgqzlPOgwvJFHe11iDIyIoNQ/8b
IUvdEbnr4S4ykOsHavSpDIDjqD8M/rlPARWD+OSvFixdayUWgO92NIiC0+Av
8w0YB3ZjdsQGpOBi3QYI1yMhcY3eLDAgjF+Z3ofBx1YVg7eikiI6+1ydWpTp
1WTlu5/PoJ06NHauvYqfeY7iFo/Sq2w67D/ZjFrzIo+NcTeV4xXG34IECWJ7
rBorqupDALqHSZEGbcII+XXk41qy0rjEkCNHTvx4gCh28hUD5ee8fBcnZOdh
V+IYImKU0dy++GJMdYwGSyXCNl8SlIlDIewrptdnurrg2ojhVtm7lNhdptH+
7pg6c8OhlFn9Ypk92epVojOE/c1Yu6Mjnf8y2E/rE8jehE5Y3Ssi1ajHt5rP
xUfCno5pPE4UlEe13hTESpRXsQ1PtJXzuutYvPn3j0JP+kRAN62W0cCYFHa2
OI922R/jlZALxZxd/EfN127bHy+gG6fHwvcZFRkOZn8d2IJf+vcCumL6eWiv
f6q65LR+bkME7olWoSKsNXzLqkricYgmIysocZdzdGM9FyjG/uMh++fTtNPY
r0zhQgT77LTI0IXAiTetu7QlGuO0KW2ZoN5znErgJFrOQkvWcVIdOErYxLJk
I2A434joOJ6xqR9sv7+sx0iOvIuR4N9ucWALT8noBUjBqU3IsgHgwCxGQ2L6
20M81ABJMKHaQimXfjczCx5mBDNcUODqVjP1yBl9KTZv6QO71+qHPAwLsSqA
8sMilcxtV+NGEDts+9IPjZ7Ki6cB5vv8wEn45Z0L4vjs7CClJCszRbPQ7pAu
N88r+AvTBxbBVj3E11qnYa2k10rXS5huER65QHpI83m8mkzA4WZ/40Q8Llm6
IQhRUU4+rVd8YuDzgAjvrJwXLsHTIqykCrbFfD9G7om6gOgomRYt0V8tTsCl
+DMv0Ynd+hKjxYSy3I6REbH9IqTg2iKYCJtgANX7yFVhe+c43Pq0zzeMrU0b
pQi+L9ucHj/uW8DdpvvYQQg2YM7Kv2tEaos9t5EKon0Iy7t6mxeKQKkiKNOr
tOiVXwphVc5MpFvHypKAnkhujPlz6a5gRArmXY5PYBOysafZ1bKZd8uGu2+d
m6M5h3JbC6Z0P27lWPsAF1uWTSrLi/W4s5wS0qOek/EoCK4PEAF4EmJy6aI3
kcrG9KnIe9V0uQd76CrF+Liig1kEgu1pBRIFSyci9dtr5RTk0Xeemhs2/+C+
11rSYfS5B2Pjdr1F98aIKrv0tfnkJz+am5kkHDZ1i+bc54f57hCL89wfNWpc
P/HCMbZuI7xWiNe0YAWFRJcmejDJY/TagcPxk39cA96Yn/K1xXP/rxPsZU6y
zad3PlNhpb/LJnNRQV9Y6MJyTPvjohZxRAGJbbAPARxZpqBz9xPKomeB7ELi
TFEEP3zOyleZl0m0AAejKyxUwdg88Hsd0ELmvWzpuRVnGQb9sSOBC6ph+iLA
HW0EHKW5OLGPZ6+qaUJIPaxeoxHvrd3uBXf15UlgkL48VjOECeZcdoaSDCRb
aPAaSQcS3QwsXhfux1bax35N4d3AobuBov2fYJIKNqLDKbtYQojW3D9OlIHV
ASpLqfwIpKLYdud1ApXp5G71Ny/haQ9hvdBYRtt1UXiqCb0pNsxp5mt1qXgD
Ac+w7X7b6k6zQjAuQkXDMIaCIRNlScUekDGJpjmkX6UegX9iPNJaSs/ZqRkZ
SXppxPm+Yk+vwOaFo2BNMZyinwL5NcaSxg+NV0b4rt3QjSkCKX9efoWdSGq3
Q19bJMakXjieezjQxddUKIlSDNiof9IGtq8G44PKxA5cFo19528sAu/vDsIj
9j/AAjcy/YURhub1+sHVvTUGq+tPQsI9pigsSBsK66rM6q/paY249Lj5croB
zRwXm5zrbNgZUBwwa5hPFAgE14+DnqEMIVzAeJfx4XbPg8YQ6ECBdtyHpMFe
kXI9Yxc1bT5cMuOA6pRQChDkkPKZT7WtXUph0w2Y0HBcr2TVR8PRZ8yzYzTc
3Cx5J28S5bfF2zNfiR3wPAVZ4eCkwspiPpfwiCWm91fQMJ0cXD9J9m+4PYOi
DVyTsTwCkVzP6PKVmX/ggp8kjAo/wYEjJBkz8DJC05Qlzy8pyKlSeyce4X46
p19JiB1Zo9A5ON2UzB97CDQ4o+NyRclF+OqCw6tTXBBRTY7AoSa69XbYaUY7
sIy25SxaupMCIe/jG5lXc/VkEXcrF2/upaGmR4ggcrUmn6ErQCF//l2I7LUX
N3+eAUsxtiJSEkhZOFeu7Og4u8IQWjEUxRcOC2jkc6fH5t/nLlXhMBdWOnun
/Z8b4NELm+HuDxxJoFTPIAmjgGtCCO5y6gy/lrPxLidZdXbapjUi7lRTLoIV
4P8JQ+n7esImW0wlk1XHYQVbeU7MSuXPDwgw5R+8G9LqXzM8KAvqFwWic5y3
i6OlMFiVwhQgPVLPefZnd3diOJVx/lV/ZDjFXfvmJl5x0GT3XLMIYibpeRj8
61NiAzMA6vBvKjpm0pm8+ndPC7bn9pIx2E3Az6YvB7C1pbXFthJB67CJDPL0
wcXw9+W8avNalWzAgL66Gc/FXpzHu7XWImaSdXqza6dhccUE7zn1SMQnhMmH
VWmEkRt0ze/Zj7GvcEjW5Bfbp4y4dSoyckT9eYFvYQj1c6lnUROs1nO9GJbU
iNpGOB4sfs+U+TLZE29gpPPz3As07Clpg2sdwfifoeA/KZTgmXjApULpOfTG
S3889fpbzo0RwVIN/zyUj6rjM1cFS9hmGQopjZhZdB6zwsO3bKu2lDfYhDig
YQXDPyyVyrFciyyuncb017Oo2JmHz1hmD0M5COxJL4+V51YWg77WKY8VOaiS
+3HEdvZbazy6ySREP7250aKGXTVkfMw6ya7Sk7+riyuM0fc4esuSlbSjaYDX
q9wOc72hBFvqIpDVI4Swc7d+PF055Ebg1For3u3d0hapkLX0b6FeIEomsFK9
+MzunZz1jjID5X9LATqMOAZ5Q551csg9tmydt6nO6Yk8kjIAb01NDZGkmRoJ
7Ko7wmTlm6RWja1plVq3qPPyhsmY8D4oHRlmpwOEcE0nt8Dz2i7+mGGeacAe
vtsy3wSK6QQOG6DiJC9L70qOmpm9k2tsfyGMV7+JFkAuVQ7rDS1H5Z17hjIb
RsWvbZI9FuvkGC6mpV9jdqPQ1jojQtGkyXM4TUJ+VttFFLLdYidti4ZhXQAj
GWjGkXrWwjHoF2gPWwzQ9hxE4bsXfEJf8wJC1CjnW9NfHSg56dTnAkiLJ25C
8a6kiLMVgNKMyAQhgDKzQFl4itZBsDNmIjHqTuh9LazDNkeNiNF9ykbxFNpN
PAVhFRLgC7hJNkURScOffq5VM0LIKlL0yY3A0KhGI4+2pblbKrbrfFbxu58W
8DRR0YV3Chjt9x+EctbUpbY5iOBFrnBYW9qD657folYDk7umqZamLvS+5xLZ
UV9FdT3QSEsD36EF4Y9wGtalKELUxb8j16Cfo7de+1bFIO+0X7xEvGuZmYpx
bwrB+xrYvFaWckdF0hQHcb5b1vX0I0p5SM5sji/kVD249rFNQw1gWm1W8nUv
U1Hk2n+i007r+DUZ1FPZDCK0cqITaVU7OpGujw5rVx5CnrlVO1z8qc/KBJVz
bzskPdhctx3wgL6t8jHS5vEZCjlQnuM4R5GAkL0p7NjeZB98Gakm6MTHicR6
6XYNX2m+ZDrmGLKRXiw+BEHqttbyzvlQJ0rTxVVhfXeW4iDgIr546GT8qn6w
PHhEcaO1kjj8yEjIfPWYTMeEApztGFLv1jgl6adTMSKg15dycNtbIpKtpi53
2fq3eKBV1pzFHiHzL6pRoTbsbyGYalUqSxMhOE2PX/3xoTaF773sC1xHwukb
Bz1tAbhS2Hzl3j7iElHJ+YJKLzFR7A9pOL2g7u7VF2szeIBAcYVAkK4mnyzr
U7JEWe8mcDpmTRxYfKGn8qxGrWqWP/AzA8TDoDiYKetgjizyKBTIDX1vM+Bu
3P6vnHsi5JPvvIAqA5QNlDNJuqMq/gGIGTZPR/jOoptuEqDx5dkAP7FA/fP8
sdcOAmrTm5mgf4HS32xbScT2Bw9rQFY6wFH/m7O+dLWW4G3iT5fZBojaFqx/
5z71GKV7dVtKOrYgpa2QPu+ax8bbhjf/kv23OCwwl2ZXXOcCQ32QP0igYvLk
+GEvwjCYfS0SCsIevoCSF+rABrsl19TQzc+Rq7/lhSFThKcQRtWDCC/LkFjp
aUtCEm9/1uNLMI8A/4Ei6595ibHjAVTwAm1V3uJqcGNT/YWdH+fagaxwHRsH
RkDSwnBW/6Yqy3APVqczzd8Ut6Dp3TnWbZCNGZFRlQoGzaHCg0H8L7fkIMhL
YbrFTH76TmnEPLlxsT7iUVzjxPw+bcy4i35Pc2XpE/yeXdV+ZVTgzaD/vTwM
hr+bbyv0wxGDpaka5q+Fs9QcJPeyre03/lWXFIfl5pu0zjKWMgz/meuKhWhB
K7eXU+2l1h4aa5EYzWAjhl7/5TnwwGESzkNn3cOikcwDbi3bLKRLSFrunDNq
5WJOPB1dR9DGVwM9+veL9d8IGgjTOSyNodhuuwr5R/T6UBILlcKRXbqXROar
2mPCYpr4Ozi6wDyFf/2PKxcRcZ76z61QQ31A7fL/XBPe9ZtQxn35Pz+/vHdD
OYczvH5aLzzx7846cMJRtELTBGjJ4lTzuinXEuK7WPSUsVR7HM10ygntJwV/
rJKXPYrq9peE53ei+q8OHoYO2Jtr3a3rmdZ5Sb5ZxvFFt/0w5FCgJqH11puM
esaQ0qPrykNPlLaenQdmTO9+8TrW/i3RRXe3XyYR/Z6bUX3i+eiUcTeMbiBy
vHEzcKaCNKDfmCG+7d0NMwV4JmhnCNnEnYwcBGdB63/ktA1x1TznINV6xTfu
BIfalssaYTII4iEZDvd7SDXnO2xdDXuY25M+ppYaweDjSEqNL2mhlsZQ0KGT
TO2529CPdHMdllNwPhgve+xuTOhXBGg2ss7mFKG07lkaZw5qwIdLjcUR9Max
thcBvqtDX0AmPyeB7LRQ6VvgSk+lonXa/iP6leix+kiKCPkMxviZqli4XzTI
mX4SZUFEx5w0RPe4+LVQu/pXad9h9sd2cpKiJ604BoJkEhtOdC48mYYfgZVj
gBhKKP+/Ynz2VEwPcZQA74xKY0qAARyPtlfStogZg9NlUcafRxHsBfgl8OdJ
uNn76qJu3XhDmn5QgN3vl5tO410yhqi9W360fjpM4ECYwxQ1KUwqSxuxxcC/
E3kRttAKHe/o0mpfU4cz2G3lvMMqFqSMkD4G3nU3yhE1Z3Is8e70ZzSuNpGF
mspNiL5eNMgX5ZUTtyKP3Sl1mH+RKYlSVsBBGOm8b6omA0NpmApF0ATH3yYd
B+K9ZrVi75xEZhFB9/Z0HAsvCtfwT8wiC+STuYNar/hYo/2fjRlNGM/MrzHq
3jEIBqcp/wyxoZEAr5FpfX9B5RphVdErGHvnPokLgnFctUa5zzljB2gZ/5QR
oPEbk8gKLqVzI9Ea0JpwvVPPbiA0Bv2n+BQtOl+WvHUsQuP+SQlUupJpRs3M
BfvjtoTr5MTYaCU8NaCzEZSyoELZc5NMmKdug/ZOaZnwfI3ptEflRA5gcwRD
ukJMSSxy1TybkP9iPCEd0GzT+4bOtaMmtOVDzBfc6VKP1DQr6aO0J5W93Rj7
TqlBNJGeB2+NQ6iH1/UtxYzXKkL+G3nzNsg9nUKW6FH0iirn24dXVvuTUE8f
XqZHcb+pqtgfOGqiboNZ0EuhLTrU3fgpAcWZnn/56eXsKQ2TrVb5GY+aEl/R
WaXP5Bp4nESbuPv5qozpFEcwa2H0psh8k+cljuPrq28JIq7wP6vgXRvkvqmK
H66Xr3IOq3Hp01O7ap8cc5b3lCnVL1B4UN59lj270/HC5kuQEOYy+XHS3hig
uwrtaFLwj6Cwv2FPlnIO4YQFnDgu+2DiEXmAC5RhegcRUHPaivo5qa0K+6c+
lYVFEnSNuunzPdtsrK0E2VoxY8WQNMCxue0Qh92QhLV/8FqC4w5DuHSpEISx
NF/7OFWWk/fgVoAwXxxfYKngSPzOYZkV50rkS5uCGmLSCQ/lQtnvHjs2Bj7D
TNG6TtJUR+5cbIKjYlRp9HNli8fIa66QkWpWm1sXeTyIS3y+mP5gX2zJ4EY0
rSY5vlmSziHBU/C6J2XGsiUQWiof7C2+VdiT18hM7S3CQN8riyIAwNpp4y5T
4UFr7lPs4zZ/IV18YNWaf/x5J/rotSEUVn+JJiZNd+H85n9ViNbybcG8LstP
05CU5yKlCYXB0dQZRGToiM5Ae6DN5wuox22+x+pb3bEADwAn5dVq6knDrfwz
dwOlZDeOFD9fwtdYUkcctJiGS8GOTvgQOLl4fRkdDTYI5dvxtgM2ap/q3O3Y
G3U83LXXKWnmhCaSKuV0H2W/Z8pxJkmszr4dMuNawRH29lv5/PGEKhs9ORq1
Zs2kEt8uBe6BMB7KB6gNszfIeYBAZpd8ASdY/8xpPIVpHZ3KH6CAE4auuoMU
Oy5n4s7L/qdI5CwnmrFDHPQSZ2tPXdKW4/cxWqkkhE7Gy1+TcNJscLwhnLXK
dDENcsMv3DWJuTHCFvg+UkJLtn621IWhkB7EKvib6s3MYoUCFXYI5ARk4v/V
nXaehkM1FMvMm4QS32CteWncugVXnsTwFtZwqnQu89Q+UbMNSBaQ9Uz1QJSG
Oqen1YhMSJRbgx34sEuOClgaF1zdOqzUTypBoUn+EXXxUhE1wKgkNhWNkzs0
SYUUr+ChCohXXGx/8MvyuwqhDU4RNVaIuBNYRLRjLcmmVOxeRru01xvBjiSE
QC/uh/sJ6aoxJ5k1/VZfIksdY/vh237Q8gM6cyfQLDBQ558cpMPWxXpOG81F
SkaTevaKP3H6CFJoZ5yBU6m0ZHVrF4avcXUmMtRJTe0lAiO6rGBLKXmX6aKD
YkGmQN7x999aJfcq8f7bUFdclcmthF74A7Yo5j+G7BCuW3aE/3R/UHnN8NwV
kis8FrM1zK0oCD1EAbAMM/1IJSrc5di5iBQPn1rCiZBrbumMKxEz6rH7EBWH
4/uSHCmvbh0TuUrLT1mx7Gf9DpGylVTu2oXvRqIKf7woHlFJGDkjCtfTPEvt
92chtphzgRUd7ihd8H6pXmqn9qXWcz1AkAPHCWD8FM3YdO73o4bNdYTnw9Pi
sfSHKt9se9qH7rjTZPnUWnPbLuJYxTdlltP1A4NdOVtCmi/i1b8j2h5t1Mqb
vspY6prgGBe94VMqrPBlob/sGNUsgO+iwR4B1UaAAcD/w6Aj2xr99mzUfHy/
gpxC/RDwUB7FeV+vyVDRm+1fUlJczpqUzQcVBN0CgP0+JnLUt4RcRrkLYaWZ
8ePPVgtlfjsqGxjLsVsZYPAWEtjIQhVMWTtuM5eKBDXAg8hPr1+X1e1uphH3
RCSZhXRxnZlU7YdCQmZe51G0HiVGgPw4B9ZmJU4WJVVo/YxljtETE8qimehB
E0P01qioAOnuEkYWK/1gv9INmvzmSrwRdJQziUgadA9DxgnEpF1AanLIo2P6
sRLZ3yRk6jy642LUDbla1A4avqotgMmAFRg1qL9UANgeZWeIM17ErYC2l9nx
nLHV5qyz2rgYOFg+XnH383fLmVEMdvykE0SGnC8n8KfgZA5VNp8TZM+qgjE8
vVaougFl/EaTaJ3ymWOrorz7iNWlirK0V7aTBS3itvZeMjRzMdDMGMbvfgRz
mxUYwGamuAqhHN+DnuE0zZO5B/s2WVYpQfuNkN8lO8Qlh5f/tdP2q8+i/k4V
urteQzoaFW62AINgW76EzrPkUOzmhW2TCJFYa+EsSDTd3E4DFTCAYZZx5urS
ohAlfdApSEFe6IDFMZVQZLiGvvTLA9huiLRrMTveaUvgKV74sSYzlI/twNvX
2WIY0CsOZJDfD9rOP836z6iOyY+s3Nhh+e6+YAfByZvDsjI9Ddun1HdBRFJ+
//gvy1SZHeYDrsJkCK4jV7mXBS87DakHfFoHxGf6swSBVM1cCyXWEFQv8VFu
4b1yomxpnlaXfG1/wVFyY+3RGKsKiY2dqA/pTwwT+aEd+pJvjRuw2jXXZmiU
jrIGqiGrrNhu1A41JvN17Q+wcCKBNYTXIjMlMJ7tGUUxNv8ZxO/lhPQpf90Y
xKYjdlDfQLL3ech6S6MudaSlQ/crLgSxjFIdZHN2PrkPZACzS94KeLmT1AE2
2qNEBjtZ2JExBE2jE1Tpc2v8/hpiX6ZHAg828RnWgeA6ndlln7/p/ksEVig/
25TmfWUY7Tus+3hX7ao/KmpvsuJUTctf61177TX/eRT/LrfMk5eMCluhJyZc
W2OZNami2fF1YByPAUEjzRacMdTW3H0Zk9+UKOlmVnno+xZrZEJAAjL4LtVS
m3i7uhryd3zp1mOKip0hpOgMiLuNK0bY7TUo4DBJQLmlQYlUnrbWIMU5RM/E
As6viMBqvJFYm/VypHQ2FXzzCwRHEv//5bJVlNigbpCGBnuYweKx5N7M+7Gc
f1Wg90T5iyKRLpRssbhrr56SY9z1MV8LVLCYlFuJaMCOdhbz4LdixTW8llbI
Dx/UEmnSxJz1EH90YL7f2pp3MK9bsFEDEYbfpasvhEglpq7ev7KlEyBy/9Pn
aOtlBNfkdIILdxEJt5cwTiPnO3p9TzHg6lm0EL27CZvuqzofSiCoGm4r0h5X
s9aDoAJZKXvzUopCR+iu+IHk2RLu6R9xo2CO2fQ64g1UmKHJtfWaB3KVeXQd
s0h4YRXg4KDLskyTxxRrGXT7/wbMBekoIleqntwEXxTR+QXUb9DiC9yA1eBs
Ckn7uPv9Rb9KFbvGN7bWwQux1RaY5ukVUCKLEmD9MrTbCc9NMIkjXqTdAcey
Mmj1J72yvGQydq3b/3QX5QOrGHIDZ7BkaAPgWhyaOxLQhOKaJlHWFlIadGTd
qXu+rO8c6wBGXNg1H7AA6cPa5wF91DvJuLqweJlCn/d3MNHkS2gTq7mq1SV7
ZOGXDhIM8BDlRq070zcPnOmDMQpnHeKLLz2u8KNZx0M3hRZuC5VXwiBlUqYJ
JwYP+W+RJXc0vvguvsz5h+TdyDZXO3soPo056wXlNmzRSaDRVDIRzbFQdp7d
NUNCPzYpRGW3pfazoU4CQPyxkSV5YCS2hUGffPznBZaQw6Mz3KbXCApDDLEk
T9LraHV6r24zEVoC7YA/Dx4DQR7pdnaf8RsHtRHGMjjkmyOeTZ/cIcXfd2Zo
kJu6C8mwX97XYW25n9/Ffg0Z3Ly3ZMBf53m3uLGqNnD+bCo2qG+4BZBHnqun
pKQgPYP+fNE5twuXZA4wQNatC4yMnrd2Xkge81lfX/efQqLtjJhxUEsTR7QM
9EmKq2kcC0WnjEZoEEWSmi57+JXW0z6y7QQICamnqlY/+17So67LUKiYAXpf
NMz1CWMH8WdOglZ9wS1elnrdiWVZQ6SvwCLQKRf27Ecjc7LUTtonuTHPGiiR
qla5n3/xnkwKDugR+K6dRxHj1HWUPspJXFHSVQY1VynOb94okHve+grIDU40
nZqmR5pziy9atlYOF2/8A+aymrFcU3aIA+GYSf3205RQU3gRh21iQftNVNao
BtEKi1+QZ2iskuQTN+YXvMLujUGc98AXY93qrXEs9rDUqXddzu72IfOxpqea
WY3+82NVaMNVh6N5eTPqENkQB+hm0b0+p9pMf/UwzPgd2tblLJjjF+AH1Tz4
FObprDzA3dd5HU+lq9YrZEozom66mj+kJGJgkhDTI1wbxy27mWTanQEMhHq3
tZzwyRLSHI0KayWBpDi4uxdSunxIOGgO5wsuabyugTRwpvKl0ozWTR5Px1pe
kJ/S1S1PRCShoA516zCKgHOgStaDWJdP7WkqI1whC/TGAKMQtsf21zKOLt/d
nVr745xS0/K1or3A1iu5kFayh3CD2oRDmVBBrMSiEyOv6QzTnPSqG7nzC5SU
qp7iZNzEQgMRHXhhbKr28J+EgvlEcslZG+n1JhV26hY9LeRWEZ/QA5eyRkn3
0JIqmwZFjq8bPteFye7SfMkAa2l+Q/rjF85bjIujlW7T1PklzAmKnu7C/5QM
D7/puKUQGGYBQgvSMcmzcbudm7vaLymi6ypeZTTXEpdJgT2yMlxVX1ZCCwuU
yzTzVvlyveIC6WyKv/rpb3plyNu4CWjvz0RBG6PLMRHpbMe4qIu4LenRJm4S
5K1XpMLCLh9I2b8BTofa9LOOI/bv68/+wjeuIcPoNcfweEvQs9jvjiJywuut
MpZlTcCcmJWF/6gmAQS4+rU3Gsa7W2Xb8kuvV3aFOl0HOd/hony0anbCJ2yq
KgyNpzCIJftZQIV9B8LoahWjNSpQaxH4rMYbA3BQROuglOYuO1L4dd5wWkym
gZhiSrQW+KFvQQEsN3NYuQhqyILHq7kYZY43pClNLXU0GjgLJH7deGHBR4Ni
aJJnnVMN+dJSvn8GQICNrq2bgrLN303jirA1Oy9T44kN90egr8OT+zJ1qmQP
2LPP7+eYm87y/f7E249GlCwmAxooAuhXRGc7HuG8q1TNr9AVvaRDd2KTA0cY
z3YOa+a6PuxJSnKPq76wDP5mAJ2Ls0WqKBFUozrX5nivqLvSMhJQ6311k5Ni
uU1QLY5RgVHcp7J7zQY1U1hdVvGPcTZe0fAwbewKj4gorhSsMUiS4URLgP2o
9/Kh8f0/6pRtm7potWuSnCBPfH7qI5IjW8oaKQ5+t2W8UgKPqnQA6VTUPIfD
6blTYqcq9Shzvmcq3MO5Lz1NsIW9Qry3/NaLjF+jZu/lAX68TMNblu4MQuI4
svpAypNznwhzLxuFcsvuNfxpFXednRKLmvA66pubZJhu3xqrIw/bDOIdvCuA
0KEckWKwgh2pjPASsqJtf5cduUrzjX9C2tONvpycrS3ylhNMN50qrAVS4O+p
wNDY5IbtR0l/0YuajgeZPHjmuVUV7EXUdE0tGNCaWsUNC1gDkR/XRysBpDo8
X1BT/Mt4PSE3R7JiaoyU6qzsjgsokwf5ut2kUh5XKuoAbNH+q1YXDlUWIsn4
oeo1Jbs1hxu9TE5JztVdZaVfSPyYWILHJ31+PEKl6JOxoP6nNeYu8b9k0MHY
Yffqh40SraQBbPcIYgI7ZPDt0X48+0Km7Dvufd4eggTIzsMeo6CyFIlujB1X
yZcNsxhqnXRQycS1gQ3XNy88se85Q9i0CgJE5Aj82RO/ZpnB9jFsEqhb7dot
lQMWMGwjWdtrwTNy38eakRenjObEi6jbr8ZDS1wvix4+Ore87iJ61JFsLaRp
Cf9xPI+xPD9t66PUJeKlYTwWhODlu3B2k5nTC99lMKwdpPtTVl2CF6UNSQcC
fEF0/HoRTd4EfWKVJ8fFljdN8MZjBTjGdNkUbT/SoJGeOJbwsBeXqCIz1DJX
Zs3qwJfbmIGLPj/7ljO7Fai8hlDdSw1aznFQqvlcEH6DLA8dyl+PAA6Kk4Mf
l3n8y9IJjgYihMkg4rC3Ail1GLhmxyNehsOPGn9idoIbSgtFRF1n+1OWJ5Vg
4oPjF1A5SIhS7cNaj1VvE5jk/Oj+2pIXjqxrAqqoO5IBwO2lmxVo2jYRNOjD
wHca3YRc/xjp/9uB7/tWg1g0F4bo7Ad1hIYVZUEZJIOA8I3WC/NOvE5Gy9el
tqriyU+lBQXKzeMA6Xjs6OK1FyBDoPJGClM8TDnBz/F5z315WW0h3jKgYHgo
jdszc7u+SVuYVVEPB5LlG8fCwtDdvk9SCD+ZuT39cgAbOR/RHoOvXuPnWLtX
35I41y04G/TQv8od1E1Oe610vhUQmgz6MgECFyFRxc9B7OgWtT4Iga+RuaMI
xgXu9/9Ej+lrbj8K+8NMcUeMPxskryuN/mKXrxWVkX0+ehAX+vTo+TDTxeqf
nLiSJhWemnWZYMR9mI1hciXpfdKfdljPsiQ7kZWuTNIWA+4SDBk9QtAz61fC
AmuD8Y3ARPl1TlYnSmnbDJA6+Yq8prve63iSWyqrOLrUdOecH5TuPz2Opv/q
webaEsvxwD7yi8UAkLCrf9sjSaJuden/0Tfe05aEnmioMX0c9+5miBfG1+D9
0uZS7qcs5A3ZogK91n05SV1NxlZm9F9zudLZUJbjhbq9TNIY3nFRxMez3CdU
VQGftzNWwdInPxxuzVfV1u7/gHF71RBRZJ2duO8IzJBc5UvO7J/7skIiOltr
Z+9SJUx2g6s/ye5Q3lxOmhoom2LYsml37UC8mXH8OQtrjEhLGld3VkYkYn00
f+0/Gi5NEmWXQ3+b39fI5gn6/wRdf+0hNarn01XABE5kdQAHyV+toUItcPyf
owbqn7ro8XpdO6PBc4OGewcOeM2zyupevQC0KonUZrTeURdjbVTYjjIE/htm
6qZ/S/KZuYFh6DrWGeoSbdPV52uMkPkjm9qPSsp1+1cme6vq40tQeZP1VpuY
v42d+kBktou0Rusu4JnW+RFh84UCN6vMW2MQ0km2tRhx3KrXOjxymrXEfupg
ok0iqgRrtCJFo8VDrMsk4ZHPEmXSyBVvqkFX+OhnMYUAqV2/doCXp9mvZIzz
nTO2zuwhFz8NX929GI2z4icmmFMPp1JTum63Bysgqb2XCKpRKP4y8/R1uVag
gvKbbPsX7+ZnS2THygM4azBgib8BaRYUBNqIDZngZWNSW0cZIDdMDDJIfVhp
6QH7ZF/uDrVVvKNLWHbwVfwovbXTOj2XTN5irV3c0lhT4lwqQL3XDa0DaxFz
0V0Df/FG+HELjE6mGdRmDB6H3zpCsslq9vGjx4OM+ns4QqTDw6YiGcfuzybf
wy8//j8Xc3EEId8Og5hWzxE6kyGJaqK0PIQLvB4+whyLGpf/vOQZwpqPjGLj
ZywVVKon6E0lblWcDDH/3AUdXKN+j9Zh/rFaQr8hRwVE8JydyJ7uqp1kihJI
XSyMAWCyF5Vfeyndkg1v5LYlpWEWG5pyllBzEFcvkUwxOgQJCwmWm6iQEaJL
/0OdyXhFmpC7P3xqK/EWN5+jkdt28odkueAxMcoXICjrOH13M7HL1j2wHCay
vnr1w1Nb67lK8SLFM14+2GAZ4Wq07aNXI8p+LYovM6qNVfDHTh/h+RAz0au5
ecAxRFOjVRX+Xri+cLeL9oLIhwIKUV6QoYMZ+kjmm79Zyowf5sAKflfSnCTN
n3Mh9YQ4rZkQEfYuMir2tQ+7YRDmnLNg/evF+X0NN3pPUL8riIMIxyZzzI9S
Uzh39eX2Ut0oPRpktCW5gew191RPS5HcMCsnpVFru5oVzUiGr0Py54wSmozE
iCk7gBHhPk2auebtMnrIY22n9ZaOkebh7b/rpOeQYCnZxHCw17EOvMQKsDCI
iws/uGDraivGxPzhoqsbm8rMAhWcMnlsdZAcQEshdlVOVDsLZhpZsS5ha6Od
5bq73EnOogBA4wJSIa2umNh3+D+GeWQvjdYxF/r6WAhV7drmHT2DDH0a0lDH
QbsNyHn+IQDxJKAMUYEjBqNPtoNC2YMQNRwkDUia2seSkhwfDCicfZRXO97R
s8KT6blUUXFc+P/0+a2XJlJMlfg56Ons6MzuHPLDgo9p2b2E2mw4RClELayl
ip13N7sCAwmlAaWI5TAE8lvkzj0RZsrJF/HGfsjrPU4qNZ2bVbKNw2+pd5Gn
0t4mnPQ6df5zhR5DgSxIYsygWTZnq255wwF8WG+HEC0X77blJg2tFpzMswzW
Q8mAM/918jNMMpmA7Alfhq1j4O2NPDx5vHLFjZe1tbrhXF7L2jA3eD59CnQJ
k6/0arb5qiZ2k/mTfliWl+b1uEB0wKep+H7ptoadaRxo49Pqh5FdA+8TwA3N
CfCj3YPbAXJNW97hZGv7E2kDuEJc8SmX4ZAAtlFCciB4wH62/URqvAGxE+04
0Fx3zOx7ZjuvlEbSbbFIvHU8F0l/r7lGuwZQi14dJo406rGqiilNk2R1R05F
p/yabnVZDuT6z7WwlpQ/ctPpUuz5AH3UAwkAYLvhUtjGaaXvJWG9QChmhhCt
UQRqz2tBj7toWxHf2W1JetFEZzpd/NZ9+oxeGvAytqAKdZk/96OoQ7hQAK9/
ASH95pJP9R6lPXk7C6/4uctuKqJEFwWPoLYMBqhAYFgt6VVgs5IRk0EFAxdA
UnwMAXOHs5tUF2b+ePRUVQfXDde1vOaDkfhgdf+dBNw9MBVWTHsMaA6Dg8Pk
o8LfQ7BvxYnjJrsrOf9Hr/iQ5MwjoyfE5UHKMTwF/WltgmIPTyLBkx0f1QP9
Qp1SnGqdcbf6LI837tWEXiF9L8C7i7ih7QrM5JPwNTaPG43qSJe43XWhB+4E
45KXKQfxyFiIW4e7kpi65Nb7ZOHCR0oEmeLzoIqTFslatmAQp60IHk88tIjS
hPjr90ygdFCfd3YjYhCmXGMQZmUGk+/ah9Qe9ACbnkRF94ifV/g+JHyC9rqm
g93oW0DUI6CvL8056d5OyzDIGu+McwmBHfHKhipM6ABtyMKyzK8JbAPOtZ6V
Hpa8tbmlCjqMHvtytGJNKL7uxkNNvEGYjQGzp+3mG6+aCO9vUWemTd8CcH/A
izE2gAIaSrk+uoiCm8DCOCprztnvK63y9Sa0n83/uPv56AkDBleDthdPYPfx
Pk1eiueH3F0qZiW4mHAJOXf2o/Mr6qQkf+Cty27wB6kywFr11swbP/qL2Kem
EM5zVO0k8rb40r0rjGv13hhhZ6Xc5BFFhp2m/j8XCvNTS8JZLFbwoEcc60vR
o5U29Q6ucqk3moWCbf3sEHof9ZLfpKsC5ZeKB8vRcSjUa6bWNqT+TDnr+H4h
d+M08/4lH9RpjlKF1rJhe5t9Ksas7kUJ2uQ3k+PZznH8AVkbNdIfVQdgeftd
k3q6KBv8DvzsCelTX9yfZoJ1SwKy6UHud6Me0P0zFkjVt6WmXcEW9kviIDlW
kpBRmtXWb+fc9aZFY7YIlZLr+QCertLOqM6QBsQ3smi6ukTCR82vbaCdtcwl
JuObvbdbv3OjjfEk7+Rha4Ej0kiBvP2OmIDeDow9Qzzay7eB7fKAaEgbsnL5
lo5JF3sJrlSmns2BXlhdS4i434uAADLsUbMrKmu8jLMAmVIaeC+tAkAnWDE3
Fi7w823akLh9OzXvI9nsA0W6SeD+d6Yane4132Fu1VrCF7RmsAw2MGOHtYGR
z6VB+g/ahR9VWPwMZzrwwFYo2onsdlFUQVdryLvzNQRQhhCrBhMNwXS0ZNIu
q4Xr57dy5Z/jAYgQ9yy1wg3Msh8PfTSK3bCg+Eb4qfxV+gM7pPfvjoX1FvvX
SH6LmeUG9OWxcQ9QfytWvMxz5rGPKZyfl0YRxxswCrcp343MMy749IQXXjmM
Qqm4XUsRi9AxtGQTvGjfOfhqrPnDCcdcRrCkn+YdCf5MypnwdlUiqJyrjX0b
h/Siu/HQhpMB6g4mFz4pjgD9l0d5kTAi8UuuuBgncgIfZ85yXAuk3W1R9COI
piWo9i6MPz4Gn7FM9ewhih3OdZM/5c2W8VR+oZlPV3Xj2IUNAe+wUoxoRUtw
MM5sRyXBK7j3FvwzYjGBt8FWLATdEuhxYzIaCWE0pPncy8qrorVTYFmlNvfD
jEB/HaIFVhC/igeb+mLp7zjW5SAmNXMGI0yocapbs25n1gF6pj9SfgJn8Yua
sdHjZA6LFLWGKdu5qrnMUjU56VJcoqqVmWIuzQeEs0nFOrXWmcSFCpiG6/7N
XqkZQsh+ChC5i11+Q41IdFQd5ThJFt1/OuK8kGYdVcRAD4gZ9EFp4dRZWJhs
yanFarHWZL2xz2rbhnWGJBq4Fh5eIKFnU7OKwMl+izH1V2R5a681yLRd0PgR
LHESvrMw3CBIPI8nrfDxYzvJ73nXoVeUWxFKsOUNLjnISxZ45nn5pqov4V+B
CSlwGX4u0JdrHJy3t0K8FaB4d4We4KD5TMqK2hkpOuCjpt2mNHuuXNb0LtLU
v7YkE3iHlmyT+miGPvBy/sC0HzHJImRXbZHzNc6X7BfKTLMlFuBYi3AQcjqW
4qSGP0UWlZei9Qpntyw/5yrynT88kT/U3O/ZgERWyNN8Hz5wsRraLdqB3jJ6
/pzRyURT2EeitGEuVShCST03qhsmxEFoCp1NRgrnkmdY1dc1yQMqaxncztzo
DVQ9foyr9P/C2XXvN9eqVDrzi8h3gHzcvT7U5mmxCQd9z2O1zoz9aFG5QWCc
JhSQfrKrTAMTNGi6cgxj7+D/z7tlquucIH16rVkt8wgrArooSsd9PXBGlWyX
Z2q6hWdwNJJnUCBCEVW3GzWgXZjor89igj0beMUTrb243xgZxJixXwN6KR3G
jBClFF+1GvL936wL8BPTd0mP8AfhTPsFi9HFXOCe+vK3TNIWf53a4tngKTbj
qjpbb9g5di2VzPp4I5GI3LqN1trnMPK1dRqsSGSlAT4hnh5SjDsGkI1YJwRR
Ai1yFzDntAei6+sACm+EM7hnX2BIjHRwevkmMHEYPASRN+4R00Rbrzn9guX2
ZFVBsalJFWRTMd3PDGBKpJjbQ+OPp32YcDBtCHOLadtyQQcCP5unBm7M+Ivh
Df/PiOHr1ws5c8cf9It8Fjj3GAv8jaOID/ACHDGYvrUpO9TGxtD9fnghik9G
rPKkHCEgYZOkbT1/VQv0TyMG39p2CyzD1j3Mv6zPxVUKc9CviVquCNdkyp6O
z1cDrtaMbFnIlOjHmzgSOEodyFYZUozyA+sT4VZ5LWRNbWgKuap4vnwu2J+x
appyJTpfTv00M+I8eBUmq5iOF/AZUGfV8Voz6M37auztznr+mX432s7Zp5Po
v/kwN9z/6rt5lZ4VbmVSDlHCv5f4i1KXLhKTc3+cldE/tli4sbrv7+RCjguB
v3APZ2LOTWQnRjOexm9b4VCW6dQcpc+PQqzy+FTmDGEwJU6oB+NOpggsdsuu
QVn2Z+JSBwhnuXhqEa35D77BwMjESCAk6aTadUqKNsICYzUQ6HH62FSOdINr
CaPxm8zpwl8Car8xfbDc4iSx7xeKyc3f5uLIaN3bW4iEBwMRrVyGEt+eobGb
YZlMcPjcN54Cw8gmey8R6tDzWOpcBr1AefOIYaN/FOXmwnWekwogZKJ2r7q/
PA1ZqY0XW4zZaruw5YjLPQ7TTZ0p2pUKRBe6qlIa9WBY9gjO3upz5fOkf3/J
RwLyrKJrSj/hDA8vFw4dsrrHdUODQQWFmQeeU+eCutObB/cNiqqkk6++K5EK
os7K01+OpEJcqqMmt9xq5M02YHFIFad+2Co2eGjsA7amdYZfxPsvHUPplRld
jkyvhtJ45aBaxOhkaGqSP4s1TFv66rvtoOqFo9qafefgYT17pjBXOjAmFXBj
I9fih5nE5lZVHKXCR0MMTon8ad/YxTXzQc6X3YRBKvwb6G24upPyx8by9+Wu
wDi2KXlg8AbzdhD2HBl5AfnFowBEOe/OVIJ5IMZ++i9R6EXA+cXhJFkRnpJ3
1ScUlZ9CV9O7tWA0QoCz3NZsNfKwDYjtQEH5bRb1351I/z9vsw3HpYa87dSy
+aBsAqJzph0JpeaXEqjpW/42IFxye+DSS+DJkN7+GUlbpi/vTE2iuXeYQ4Si
xMBKi7fR3KVhs7/ekrMLMTXyYi6MOz8lNuOZ/evptX8xa5Q0KmvwZ/ofTRrf
KVaTvOY2BlRrPKeJV7pOGCNfqC5XVePrZv98Z51B6YMq8lsjS58AYvLb98Nc
uIRyukNn/phRHIMesbT8nWu2a/88P6pU1TCh/y+5j4tZHsvnAQW6XukGUBXS
j4ytYy6aG9+lABLK/Msd8ce+9F2L5iGQGdnbVgESV7oQcJsMiTlBFuZbqpTF
FrixnQVj66PM0/ccKFuhnZbAmhT1rLpvSY/RrzIjiIPMCrZA1QHVtSMPSiUE
XkIjxK5TeMhTkWVIE8KXPcaxVcaY1fyx2G9qhgMcHqapsKk2BVtmYIIrNtcV
Oqxlgs4vEiCEZ8UB72FNhVciZaQlcj2My061iuzqSp2sTC/sLz5QjpOavyDJ
9FmiWtTf0LtMepSF5AcHjYEu/oWZ0j6q2/cR1I+X6PEBhEGdJCXzfewDUEpK
xAaVKa+5inSZ4EBECirHZ+9lDYiCFR4VM9lY3k1zJ5GYAbLvZALrAfXEKxk5
kQt91no2H94mR2BxKTYJ/unUdRJ5tMBCtr8Jdb7sH+FbmKNJ5ldX2nmboy8L
2cWvqLukXiiTe8lBCzJfhf/YYc5PaaUOz7Wj8y2rt28Qyil5ePT0hjKAA/oJ
l1fdtS3RcOLXBpfx+T6EWazdQKptI8WBYTVCAwE9rFQ/MU0ZRuefOvA5xOi1
9YuEymjiqFjV+HD3NzSatdDSLxkVylboovuVuIyZiDn02RzYjM75PuSott9q
NXsch/Z0egOjQw3tv8pR2K1C20cnLqyuBTa2IBNSlpwFihoylfdK2nyoV8MG
S5arGP2gk2ntIwOG/ljiwM4C6odNhDf52QETpsKWd4ufjFib10x2PgGct+pl
sTnAN3BcL2FC8EOfmli4CE945ldkIXd/2xR10H07xuaeTl/gp8UGVyyXndmg
5CebDOW6EaNP2tEnjcv5F9bmQfKQxu4C9juV1QL/rl/5d53AU1B8Sx++dw9x
fVYcRBZ36bPRi/uZe1GhxT7XWPME5EiboFHs6FkaRMT5vD/Suoz1KkxqTvxV
y2feSMJDk9BpQ4zlsFFMikMSszBC+pmHkiy6SIaOgODOuYCXPXRUn245YNa4
plz0yaZVHq2yRteQi9Yt0NM7JQuY7qrvcEqGQnQVuWJMZMGGNyVEaEHpvOnG
OutCLumSs7j2LeHPRwrXMi3iUcr9WZbuB03Wce2DZv1ObODqQRvimqBcBYM/
iJU05JJ1A3wRhMu/2oDjsgiQ7t7PQchQP4s3wE960ZIqprIe2Ns6lqzBS6cK
FBesBg8maCBw2GLTX/6O3b0fUMIDFl6q7Im1IsiSzw7UbXfGkxu+S8j7IFaS
k1v8l6qnppQQAv2xvff5PVhEJg/94QLxj+04zRQ79T3YTCtlgpyL1KuYhxAr
N4qkPtSf+h4jzFnD5p+KV1omL8fEup5Ac5sIrr3CvUchpp8EyUepHw9C6JO3
pqhXhUeoUPgguXI3HIkNdpIkC/yQcyauYjhFhRBfE3uwS/q40NaGBAblpeqe
TEg2RLhmapx2rTeuH8CiuvM6UB8rGd9Axw9n85gKgfZl+6xTz32X8K7ZnYZL
ajgsbz6LIeV3qbvMH/1eZpRj75xG0erP/s88InouP2KGLH1fDWz8ESs5RALg
dXQtF74ioQ/hZ4TeCH3Az3L1Y761hUcfAiZ7RTiaA90yqL1GbSs82qAfJmzu
cU9l4bptwhWck5lzcmqqe2XHGr8rDMgivaHfXrF2/wSFNOubvL/P5pnSRmOf
v2HR5QfJLdS4Q08Uoy7dV+EOfQRhBwgnO6Eu09r/fZLyig2IfhvkdAAy2DPG
FzOtOaUq7xPCsp2+pb3hyp3MM2F0pyhDTsE/cJxAiPDhlpb9/CgpEJdEORJX
AenaHYVuA52xjDOCLfi3B6JllAATeJDPTOmERXGCPgDFX94mrq9LIxHggVli
+lyJeuF201MH8wzpE5FnVNS2NGHSvZ4M8IwuOxwqocqg2md6rcYpgHdPm6uE
S5K+xRvPTtcjldWi6yfWvMy8EWI75eNKbY8SIbOi7uFkabfUyFtUUqLf+T7W
jWhXuTkCEynSoUxjOQTvEgvqDl0j7mClHtxe/a0Nu6SxBJs4/hoHP4dp469b
0IJxKAIn66C5NKNL/xVqjkwresVGGdM77XdmhpN4YaFfJIcIiGP/vD3RUDfv
nHeARGls1N8YfSq+9xJFxY2fSO68W+b2i45nc3G2xsxd9xv/ygSoD0gjhTyD
pIcYH4jShNoE9SCVGGEoG+BwWX9ZFN5m2wOs5HK9S8Jya/FQ7NL5r2TKngIm
+a0rpSs5zrQ2a4ZOfDHzeZwiyW+R/x8gg4wTgWvoCMIVjBRYqlAEDC70cli9
D4pNGeez7G4VrKxsbjnvW2fy/iUWWxbreD+q4PFv7C9/fn87Qf2B8ZNC3jTU
GO/J1Fr9kmpunwAMFy70hGDwADROQ6pxwNAzE/UTO+okmsoV+mqOX3F6hWOK
Zk4cT4XQxAxsODyo5r+fc0tn+v4CHABvHe0vlTQyZPbw5cAuaecNwtvp3uxM
e/FC1xfBAQDpvonLYAkv84zUpVlL2n1ub90WUnswD731FULKU81ehmFK8BRl
eaPj6lQ5WwgQfeqKixApxY0snJTiyY57JMPqRuvmn0w+/6PqhxedtAPI2ABs
wmNh3Z85a/uDT8DxXjzdTrkAemRC7CFGAjN38kfvESvIfdL/WtAiT8NKOdyB
MFXsK852Oj+pF0wUg7PPMJ16dqme18LmJV7wjCUg+sRpc2gYPvnUNxZoJ7RS
wFqDgsZFzViJW6p41jSqQiRlhoczyvSUDWCx3GOZkIfSopuptPgvTbkQCR1c
6raVXzakK1PlsEMq57OI3MklKkX0/XRQSb6JPfADLKzwAnim6ewOTWrGrnL1
0ch2wKD5VjLVm5Mwdmv2rvEeuD4Jk1aZsgEuyj7QtKV+2wHIwQiWcEaMoVsr
lmAkVgWO7o4poJKltGG1PgSST2DBjrIZ0hDBJtTMY9MuEjM3MZslIPN6lIKW
FmxiWOTCgSSK3gDLH0seOKFUJDjU1BRa7IGWjIA1ZB2VStNZyf3pKZg14LSF
kv+C5oyW1XoKTOQyB53KZfTEWMfZQyL5lNrQvx1JmAHUo5m2c1IEucBZ18Dw
QiTSiFIeQi/exfM7jmsGABvTLa5kSBJhzyLwZz9gphVYocXXglxLF4/jA7ec
mjiUTi+YAVA5bF5vHY2rESzlgmHe0k3TD58FR9FqqH0cAlSXu5l3rCy7tSHJ
kZD7c6YnUcceBPT+XtREa2zF2mFgpb5fTOyfjPxj1tQm26JtDJOqp6RV1vUJ
j27dczvcE+c/VeJwmiPdFrPrzI+zB/ioDUzyAJchV39y7i76uNAhQmMJDJZD
IGwrUjaDlvJ7yIAr60Rtn9ATwHFSYSsrbmaYDY6VJsp9GHi/20pJY0J9nGR3
4q82jV9Yl5YzYGuuN9UyPILa277St4zxAEixSZ62/omyODt1OZo7a+/OurER
FakcqFykOKg5n7cYsp6dnmHVwPN6Y5Fr5jK0TDAhQxRSB0W5xxnTdibAbDvo
mbkvJZ/lrf9TVTQlTKMqA2zecBEMAhkjpNUOQWQTb5OEktabqVEf/nJelg59
0HRkN30XnzLj2rgNpJCzXKNROz9G9Sh3F+TMTZQSAQDM7CYMFmqYLX0svQcI
0JU8FD3cdwy8v67DoyIMjPbcN/T7RQNYRHjklT18T34SbAswogtmy4tg3r+J
BLAAOhi2pqH6vk0KJZ0Tsk7wfX1v3Pon5+oNxeFQlqDDRQ36DTTQSvuQsUU0
edBlAIuprLofZPGDRnBKfKYlg0/reFqwGT3s3cBfQSc6j9rccMLkt+/H1Ow6
iFpZVNj1h4wAWDVjtACDJfpPIHB74h8jKTCfrmMqXAJ6myVMVsjCFS/igV6K
5y+CCQZUdc3esLYfgpqvdi1sNdN82cxlXsyt0l8+Iie5/Cmsa8acWzSgTQYy
/F+eN1vqeiLB7T6dxOfCTaQpY9BVGNTldfwAmNqOpjoxygMqVBa2Y4KsxQst
n+34EifcBOqMHPv0jrxd4uZ48wkXZCCBKkMU4DfofOddYo5GtZ7oFE3I9xGQ
rwx3Qp3TNm6MMRgFgEifgDk0YkrEDJcJCEKS4oQHsnOUBI0K1WKYOfDeNco5
bLrgotNgm7T2w6zZB5GqgfSI4eGyUid8ApJ/zXvXBwmEHNmj7SztDk7mQIQj
22RNup65VhtPjOzv17w8838atrn15qL4samO55rIteJmMTlSgN28meGPfbza
Q3sqQICTQNp9n9yD2xWA43vh3L9Bn0i8BM1FE5CJGGTobZ3GkK5/AonZzams
X8Zbag7D2/GxqT16OyB9XiafiZGEW0eE0pAxr5+h7EwdYGVxXnC/BAR+ymBL
1THf9Ub7FHOtIi5xNQ3sYNEkDqQigW3d3DtbQnp5bm5sip8+PzcD8ipg4hjU
XjGdZ2Zx/Z/1rXpxiyDsccNAmwPbVvryd0ePH0wd8rvqI/cfjzbEYGWKTotG
eXApRyR+CHswVkSRIOc/WXybH1iKMkLWH0sUXmE6dmMNVBHRzUyEkiSQ3gx+
51YlCsQbLtlMi56KVFKYdE3JZUtC0+ja+sGpjqS1V32FIu6IDxz7E9cRyaBf
lZmj+6z8T3JUzT5Gm4/VfBXNWHsadYiRXVcMd7UeuLgwIDFJccpkDo/hvIch
SkAP3J8mombnmMP72XFNeuLxJZEY547Iq5HXXUOJqGaQ997yLmnf/u60NG0/
bfq627NxWQF2YFlnxffms+qNa05b5OW3gmLtDxfsD0BC9rMe2oeYgUgo3mRI
qRAigdZXf4/BlaJBA3Tas0TBDtsu0ti3y1HuEzbICziI4orZekbvZAMFBoEy
04uYN5Va3/81a9+I3Z3zXQxvnEIUuKr/Sdy8oZnSUYv7mz2gH95+iYw9DDKW
tQszuTiATh5cVQJPMgEwe628/jGcjLog1mBdOaeGQhCS6wk/nIZrxw52BUED
JLc9wFvXg7Wsn/jmH8O5u10QhIzI6hmO/ujhMRhR2Hch4qVFO8LQ5PWFW1dN
GN9BERIyt554yJ/FKTBqG09wfixoBNBw5UHV2fag+X7ek3bfxE/fjfxVh/y9
smH/e4mQYbZC0ruPWEBmkNycXh4vvQvkL9leroM+c7CbakcTsJNeenO5GTRc
HoKzCpvelPwdKurL04urwrB3iuveNn8hcZHANGPgc5yTBUg6REdPrZHEW0fh
f9VZbncQhYEMXAPyKta7LAm+v07MevN2A+6AoX6nvk8sFtttXCyxTX1PzVKp
3JxojpwQMLC21+rDjNbUrwmFD4KUOrrGVbcKE+2Gq08MBWQdvzmvF7PsLwLd
bKMxav7sjBY5sf1qmd998WuDKgqktO4cgITcM3rH+U54lDHqxcO9jSb+TfRs
/4/KXElA/dZsukKhh+u5271oooO088m9kEupOpIgVnZThuN8XJq1CrE5ILs5
WdQJTUiB40EkQjKRlJ6C/7POW9Qt0+uleItcKp09NQ46aTrvR4ZAaczezYrD
s4FZNiE1JSxKSFZnJ7+2sb8kA1OTYWhIykE9zyzG3KwiRl9y/DrTJ+W5t0ch
fTMR+eeqtPtQ3fSv77r7ge+LW3GCcFvL9olW/dyIsWcqj23y3nTh/sCQ7/lb
0iwPCVcbWw20cqAWafi9av49/Jjd8XJkmYpYuwd/2YD6Ltbm3Do22LiSkn7Z
lNdi1dbfbzIq0yYXseX4KzCRSXlQmc+wAQmSdHrgH8CNdad0XUSF6WkMyxSp
+PPhdme3bBM9HGhmHlv/cL7kFdgiBpBe/jPOYBb0DM1W4WOtMBasWGaxNUiE
04Z89Dk0EkNHAbFxrQ4pNtXZeskJu4I76HEg3i6He9mMwMuQbcZL769QxSRb
/hRp7LCIMbvGcVy8uQHk8PMjx3Oi0sq+ohUZUGPOT7sVmlxGSiG7R4mUGIpx
P52qGTdD8gI11qxA3Fs+m1Jlhr157FhP/LtbLI9BJ1AkI48Z5B8sZUEQPPY7
3WMPKDcTDCF2lI0lW9pMvEaNV8284CbLrzAI8/NhhvInhdL1FfOVrluAZ08v
96tyXBZKiT2Yie1TG0T4MFru+cF8mZ2gteWpUxnwhPHMkT+ii3KtBxEq27Hd
C/DmmJccbRyvHcR+l4A4gv/qp4P8m2tpTaq5OWloQGVcNkWvTpVN4ENiX1yz
GpjnebRwBhG0GcM1oHay5mOMH/RvJ+UsSBi/o1CiWTuixQDxZXErUC7IPv/X
I9hV8JjG+t1GOpfKBbjy3c2wrR54ag2eP4j7gDU8Z6oUoy/3hiVccMv5Z50o
XHo4/xNxMMlraY9SKNNapQDmOJSiZO+w1TGKL40rVvnZeoccKh3P26h0+rb2
RlCivfSTPswsGmiQ4V3//Qf5HblIlvq39Egdk6PEOLeZKlf77NrKKpAp/zOT
WpqkcJxaJJoFxQXzWki93uubhIrsg253yfQxwHY1+KEkAYvzwbYoOu8ceAqC
BmXfrdw1REY1Xtb5GAlulQ+2RC9E6litkThh7SoLqr/Yl2qY9VEBTPfkps4Z
SXcmLyr3HEox7cNYM4zu9O0tjA0Zfxbb3P3FlnoiQyCHVM3Asrkdy30hHG1q
d42QPV51PXhjQHB4KRVA8BnHT4uiQmnS+8F5emCzb0vR/MPrmfRLgdXpD3sB
C4Q/L+RpSLeywL8w85MVoB9ajoZsJftU8oxs5dd17eNsJdHYCvZ0cANIuJZs
5OfVW3bPNUhUTNHTB7Jtz1hTqVtc4jmye+4eUtBiz+Zogq2ZCalI5GKExVsx
H8Vr0FW20u9Fpgh17tLSiTht7YE7/djBc3V/3rMwN7HammSumdv0a5WF79a3
pfXK3W34ThckZUorss0tImro36a3OZfcNrzaSS/ZbfS4dCe5iIh+csLY9uyS
bwaipLxWisAwPf4zo593/YLLoDBfBIs2ByU82mEyd5hhf2+mQaEjKE5YXtE8
9jY7FdVWICWSBXQkMlNrWwnveeCFA5myHnZI/5Xt0FmmhxtpHUVQQQBzGn9q
HOFSEv8KTL9rSaGocG56dA1fLOk7L0qt6dkjsi+uOTWiagQo85AWrVZhvfHV
eA5jSy4YBu8PEWivhNNy/EgV+aaDGA+eJs2l2pr8Xi8z0m1/ntlflWflDc2p
MGG4ndpncwlp00/Py+m+TB8gCngHHIi50kxu6vQpAlGfcrss3pUcZmyN9RUu
CGL2UQVvGsJy7pM4/e6amT3Tqzs6Ykpp6JxUIcicDzGs/IIhxxcFjJThJzps
p1pOhJn0XDr1wJQzD8M1R1lYpJ9ylVDgDSoQIRTL3CfmQygNXkNCcnnJHd7e
Or6ZMGa9/IAuurZgHATxeGcXqkgvee27rrCW89XN1yBJ2OoCSCOwzL7B0rS6
qkR4oqOE3TBO1gamHlsqupAPKl21llJyS9dhKxn7ZxM/+iJVce/FfCtIo/gv
b3krs6T+CBpgyN8t3KF4s6MsrqW8t8XrkUOaXTzOTqIV/9ajqVles+xMYnng
yKhF+oDji645crv/BZd4GzTujbibrCLin2Dj+DVv37jd9nASRnOWA1TtS+eV
xvHay2k+QLlFvBrmkpsAuirBsRJw8CEp9NQUNn2h/0WBOdZ7QQJgIXJdZr13
8+r8X3RKGcBhRGREdf6+mudF+GrIizKZN0c6EKwSkLGnz5uB8Dx27ig5TAR6
EMokI6wBpgAlw7PfGQGpOBWxnmqH0EkKtfJdP4cq+wls24DRYRo7w7ki1oaq
TrXt5TYejk3rGuC7pcomwG2NUL5Kp22nU8zc/naBo7KTyzStYRCQPHHa0dHM
fTeUW+tng8HkkgZfids1DOUD5aRb5CS6elxdVMxbiOMqLSvjexz/PhJ1H6NU
YvtovurfT2K70dXSOOx/wBTjP6eWE0rWu//VwlQcaztmzfxOOO3L8bR/Wz1M
YB+PFwoXzMPV5y/6KkSkjF4vB/eI4dq3vBvS/IBgFpHf628oTL2xabohrV7M
NSfNmGLev6GVuoWGvMYXOdeBcl8O+Xxhd/LcM5yczh/4xxTB2kSPv8V3Qidc
VLXuJVr3sx7rXbT1WvUDQWqSxbBlG1gFCX3Lu3zSYohoBL6wCDJSkHb/GFWv
OisH+2myVBFNiJzqOJNiQf+BubAdhWaKpoSOm5wV3jB/JRX0kiJydfbktcKi
bMicj90qQsl5fvix/+w9F1g3yh0R+6IdN82HnBq433RxRpBnRORAAjBYG50+
1EgLYDCCQTJDBG9o+RnMBwCiEjw0fpyzig7OQSJD5PnFBJHjTjaHeCLewGPn
ktdaSDnxVzrb9jU0GAMgzPQDZe7LCpq4m+NOci5wyblfMHgAGBuf4PCJOSf9
YBP0uhxRp/FiATl7i8Q9nhMW1yHctz+8PDvvNv8tTlEhdjl9XTDM+ktcH8AX
De3DWp1TbBJENeWQJT7TN0lh33y9M3stozJgk+GDca0387wpMcEXQTNhl1mK
JSCi1cMRoKpYBr2pATmXWxaGoJJt4QI3fmDVUiMhjcsvkJALNmQyR4A1A+gH
ZHnRaFYMwBtpfwgmuvnDHeEq/rdsWh8ov7dONJbwIM6vaFpQs66to3OFWo+t
So2XTMBWh4JWDO7UbibjzZ98SlzdnHlIvsuSHcGsPlfBaNOCO69TKN2jp5fD
q5pojHAzvIlWRv7Y5z08P9iQejvLTbkx0PihoXDGdUdCI48T3CwK1KOxPMhM
MLAfMDFW6q5AAHVqd0Fd1Pp54PHDYW/Uc7+H8jqt7/++LFS53XeFy+o3h7UP
PqOyeVg+Q1TrzQc/pHwWuEQrtHiRVCAze5F2bWacavT4RupRulwK0QYXN/hK
EDVBTaeQHSnZ86BsgiXG5MeULBuV6olXxTg4lXUVhLpltZM5vZnOKhT5XRm7
x8zJwpNZ7Fi8i+H0XU/4el6CX3uYpA0wC6+CH6K1VcPOmiQlgNcgoNnmKxsM
p+9kVLk9ug5DvOsbDNHviTBFJt7v1NnsEa7FYVGYSnZmjIG39VZ0xbWJc8DK
ZOaA4YLon/jL92H7tQSbJTZupw28mXG2RSQEQX0QH8RJqhU3wg4fXZYjBt2u
nQ8O6xLnN8grUaX8vPGQMiWun9woC4d871pRzwLM03S9SK8/KgYxyhWG2mB8
4NFwAiuCb+nMojJwO9BbWaknAJJXU4iiJlHtO1PP43/Sh1ktMUVCutCOpoF1
IXu81k6WUqmTDcK+VmMoPnQbUQuw0KBW6xFTV/CzpeDCnGWjNJi5Ueyxe8oU
UA3ZmjNWx0YlxCDwvfzQstaYPrtR0yS8Qxuqi1zH7b1DxP1Y+YKhqkdry6BW
U9YugPVkVucNS1tfX0MgPgQDUSiprYU4mWoBVzeoEymvJNtcdtOm3qPnAqAq
FbBsxHvgE9I8PaTP+SMCpcv9TFM04KeWW6TAUETs+e0p+pHy6Bs8RMjuhnfQ
Ncd15TxPvGds5p5uyYDGqIoQacJzXQu3YZpZGtryNDtJgdhU0SIEjQ6Ep+bd
WhvUj3FwzW7TZW+7klM5Mbg+QAvaZ5Yj/B6Ug1J4wkp7yvQveSMtVo0aCwuD
V6BD3/ElMj51vUvCqw9eLMAVf+a70/QJgzc+trIir8r9cY2MLHuPGSAOTsRx
w5D7BpUEja27g89XNri0Idnx7Oh3oNxXGoTFpm6BHQ46IAdrAbvgsmiWm/K6
w0Nah0sp5ytzkTbLn39Mxg1KAjxSuieubldMRlyxU7SeR86iTld0yNcKNSR9
JZQlGcgTxH6CbkKGx5+cgmT66EDyjYEI7xhrLQt3HibhaW81pdvG1P13OphD
YrpHIttlnUZLR/rFhdOioNDG4QRTcf1RKrovYdAuYaDWmIRmeVlXs5dwDqTm
fjZBcp5lJg1sbv7yDat6J/jaV0WBx70YuULplncwusl+KlvlsbgbroL6VLA3
k4GbDlM2Oy3D6gHTQ3zA79sxbUT6MH0lsFkWdOTKeEe6fd7IQztD9JyDYW0I
g7RckuR9i5pc+Qg/rlcKo81XzJGC/hj2wC1lDeWq1YL2FMfLKFPiWBxC3ra+
tMU63Nyv890dOiUG145S/6RQjBUHeHZNjCdyMDlPrUMnPIVMWNvtBkCN15ra
OstzYiCgTujEQpQZz32pVVZ30wLtjx/E8qOQnn5++s+nbrJZp9bVHwYHNoI9
ReccTyDnYtw/RT9BirSvGUnQO7ssamyG65clow1AKp+AHYFcPcI/WVcY6wUL
8Wa20mTwiRwa/FTGGBhcByge30gsQmAz1niWCAg6Z25yBxRiEaFNtMfabWNL
LWtyhCu4qkS496iLRSylsu6gXC+/T9MoRaGyZjDbP19cbd9eldQSgc8f/nb3
mIP9C4W+q+grMvT9YbXuX93RUkRKqHIz6Xf5RwQDjtpHxjVz1JXYI5CRRwlK
b2jrzqUuA5SdcP6X/e43dSOdjTsvvw+Xj42BV6Yw3IBPn520I0Ls255u+0Oa
w/N7ogCnLeZcDsHeLo0pp780tQAz9uyIUe7v0oShMIvdedL3sSzfBiZB1DPY
Zl/SIuuS5QE4szuDehWSe/pbwZyqNZin5EHBwc8a4ZPliWD+RZEUY76qU/mH
GnzDDDcUqMTqISMf+5lMHLnSuAeOKyw6big6JsS7/qe3o95U9V9nNrC8Y/Fr
XoH9KlkYqLD3q0nq0suQ4h5E+Ulj7Sa+pi5ezqqbb1Ysv9jfQF6rR3tGqRBT
FGwmWtWQzxanoihda/0Xi+Bl+4bQOjEDwKnTGjo8RpUocFXIf9uKIZsymCb5
URTg9eX23g9Jcg+prbcs//Z1pGKdUo5iiW9JxIuZPPRrx6A/2VRGdJaO7Dgo
3+XDTF3KlJGxG33cAw1Jc5Sg7o6wY3aCyzr+goQOd1pWPC/dKZGmxfPwo8kL
43/YtstK/LAyV6aEp7eHB8fDzx16DZhpJ33QaBR+TltUAmMmXIklEVPFEHMt
p00DOZyhBxBX7Q/2Yy2mTWRz5UaGq55xDrLXKlS1eHnFhQ7M6gRilPnasXtt
2zVNs1O6bir6wH/rLqd7NKdCIxTUGxKFQFCiOLY8K0megN6yafu4R17bEeHC
15F6PMHZ6ij59QDBOCNmPHeM7NK841osqlp8D5mlS/E3lrL8BCNP7dcKgqls
iOZbcXhkH5uQ1UyHB79amritkrLWGFzDpOA1k9WFrh7LdDi72ywC59vtLSqT
E1L8t9ciJuDcEmh7E4rSRGIi1prDA/An3xdpVYBelhpjpX4UILpDm2/zQypJ
4oqoHBecSkZbAefZxEaW4rZA5iTyTQxwxxmHUg86DFlZxjrgVh+P2tuPlZDy
Jt8ng/eIM/MgqqOYzo3I/O3YtG/Xhax94eqTK11iqcnAA/xWZkHLt4g5AAF2
/y3AJ+duqs5tyVkKqDa7Q+ZW5W6e9Z3Y5CYsnoex1RlPhmPOE4+Chx+4cAF4
4nfRSXyTGTE6c8lFgiZLvx43zxPLbI5v7foa6Eau+dkr/j9yWwF9dMeGAtzu
CQV2eQfmZ2mtzzmlECsFyM+a09YLFGSc+mm+ND9dODjPkEJ/5xnj/Ug5fgx5
wAEshHqt3fc+srMrcdRMdXDGtPTA1Tgwficmra0nXpiTxHbnZuclPA9RgQhO
wn50viPRCyFTvnxE7GAsSYfZH80TJFlncXF43OhomMQmYSiwMNC2D83zf0xU
7DSdzy1zLnHQeVDrOvx6AI8Z0axHtGthMKLVyI71FT5A3eC+wnNlK9VENTAQ
7HNjAmQF5eN0GTPVxENIWi4m3htefO/aBlF/SFcsdxuO5L1h0KWSelaJUhJH
QQYuxmQ6s/fFjOs0ubcklhErZOotFzCdsDxbT8T+tkeFRw8CRED35OuVsdQa
W1Iffaw/7LCeBnQhPuvWMnRh4YmrJmAPo+AH2hWZhd+HsCtcs3wkanJHhD95
20vi89qWiICR89vNhFOc1U8uiLPGXk+Mdsmv7vu/ViiSTUniw6reHMWluIfC
wHaqgZByUQdrXmzuvKjiJYYoB/yYQNuIPR3n6KyW+FwTMD7afXk7HdEklJ5R
iroQXR8Cx+iM8ePDGdZLNO/+T5dJ6T3qqOUt62gRRJMYdpKGxjrJyqijwtDe
rhsW2JjWA1af+T8wPB99oMmZGWbfzakdDncJGCSkxpo50kv3EWpYy7s8rkH5
eMAn554aMaZNVLelYpHstqaSgdCHrHV7t+FftHY4Bfcf6cUnq0MiQG08y06Y
1DiqOvtSNoPl5aRU0xmVNps6HlGYajhb8HIJiBDv7QfWI3RMbT7PbHcde2AX
HgOym1wSiu6IJe3DORQCfILPqxxzXYdf2/ALIFoXBGwdGRfRyOjoc7nsWhFl
l9JSX3DaF1EeYzUVDi8uclx0jHK93wF3evr+lbdn/CZ09q/Nrl7D9ct4UpNB
jtu/mUYFl0fon5V/soaqQ5UbSmJIg4pKwzX/LC/Tt12FW8gJVeIOPhazkvo2
py8H7jJsPe8wAFcwBgzRIqB0LsP/A4WSDIrWrmkN5zXvJJb33ED0zkhh5757
Z1kqKgZFM/P1QfH84U4MlWCrIEqEi1lsw4yCzNHXk/9oVFTlkCoQG75Z4eNt
jExGdtz6BsRGkxGsnUnBS2zs+8h3a2hkLwhFo4nkR5x/TaPD0DL3axOIb+uH
b1PTOPsOamEDnuWOVhuSgkl7WIWwzSzPuFZyn8fFo6TwyJw4KRmpj0I6ncWC
4uzuM35v5VcT3zQAj3/cYsiTQbj3Bbw5IRQ2nTzH1m1AZvsRclWFbcMrNedh
60jGt/eW87b8lVhDUx5orBx7Rr89wKUOKgnLVvUwbLntE+lxcrTI4HtK7FXi
zQkFtB0CEWPZf6XtVASadB8Sxqcvs9cescpWj5GN5AveqjweSdYP8uucrlru
MMTUbGjR9GP0k9PGLAq9CnfkfmoEc42JaeS07E7FEKmsgqKrM/D6ba3XSsdU
6kLF00Fs7V/oMNWJQztGqmmHP3c0cTrcBRxP+shDz+RwGmDBQ+ZWyW5xiQBj
E1L7OGHgO4O7j4k5CeD63R7ILuoNdI8gFukxeKOOo1fBpnWJTtIQz+c7yUMd
nxAE3EVv49gxPgts55VwUiGAIO8F29t6+4RkGINrqadrlYDfUpwLJVVxmTQq
xWGQlIXh1CU9iwCitqnwMLS53ajZlp4+JMEq2AcRqduDzT6j+E8inzlPak+u
JnkmICzNnF5+qh3sHJ94vFf7wJmSDw3LE+tf1o5QAEN6y+T23E/xeCyByY7Y
v78Ca340pM+1lFLzJ7LGTgsHEVKjfTFJ2XAyBhq6+BFgmYLKQZQm8cy3lAMx
rJ1mznwMF3vJ31nrayruMbSDGRDRBtDo2EZfsljmy7e6VAODlL8HfARpQc//
qNUk7mvZ/C7Q8apB4RMzpgCUTrOnblF45SPyJLpgOzHAyXBy+dAnKkl0x9fj
HiBnFiAlbrLLHTshQdd+JQXXKdslpYEPjOr1G3PvWyOM9JKgKrbV5+CGf7ol
TwJjhvBpcBpzztVPhwejeuGHvwftbltPU9y2A5lxjhh5K3wgdNN0qzUa8hcR
kh09yH+lKqyfy0MiUYkvKi41PVF3yhzGbuDh6cBIyZQblXQHFF138UroG/na
opeOx3faYYinD0DzQKfaVxvdoPnloMihWbeVxCYv5khyAa2lw/uY/KuPtfge
Ldtp3mfJm2uLy4DcIiA9ez1Z46Jc1U0SKlfnHf0csNvQohmmgqPxsu8oj2pn
dDgdPOVWGl1eJjikEE/VMWLKO3ser/45jJqxKN0j3pWAJH/w3oEOTZhNI10s
rqJoVyqfb7M2u/nO9b5TcL5Rytra32VLzvb2dzs01QciOc+uQ7B+g7b571Xm
fcxU43lYPi3l8D4qIVRtT5qQOp21T7xEwk6g05cAyzNFXm2d5x+yWDnPdMnA
lwSZiHki9AfAyZlP2v6B2S16JwCj6cN5RFtEFLO1sAmAJZY8POVbY14+AGFg
SwmzFVqnR2RRs09lZUCBmna8xDqKqnQPGWcbuk9tBVjD76OIM5iHcRHK9CWs
mjL62DzoqLpWL8ycf8K/rJ7FJJK0MZ1YtCKEjPQ2yDheB1o9MFPZlnq1Hsvd
8bNjqUYJRKGc/riS0aaCEUHdwXwZiEISJng6y3ahVNRaaizZ2LTufvyi8gY2
NU3A3syoim5IdovYkXmT7QuAjQtsC0OcZwtTJ1064fW2VIJgtbhqhA00FfK8
1IxXG2kTeSlf+Vnms5xtPeiqBWQls2GJjRcuKZSCeB+NJzLu8uZ1uFmoipXR
QgcaXHZRDesLcccvbI7QQhEr0aCw4lbXRRw97t2t9UAcu9YxR37wC8Hg5qaU
1corDgpIRf4fcBfhXcs+AHzRyEbYE5eAh8SUSVskZLuo+QEdJFuanwDNqJv/
Bki7ezyZBwpBnnMB3GvOHF1/8K4vn/Toinkjnt/6TNnNuTypCCJzmodrCvpX
gf76wZexrNa5lCyxYI4RdliJ6ZHeoFNWGpB7I4WrsIDP3wXykrnTwzpXGxpx
y7p9SsxvT1FmuR6IpAlmVrnLJEs3tQUXfPx1BTTvdPtr+gtqdqhJO7Ie2ZUy
UM4bVnNUruk2tTuFeBLN4J2RLSCZdjbuGNmubLXYUIOgrXo7velzvIMIrBHg
tP316HqEKrd6AI8JxYj0Xt3hvHWylmlR3DjqqWFp1GmAWPzM8a+vpGx0mMiG
v54ul7uMzExyFBnqTrHPHRMoLY7VStNt4K4KDPYDgm0eJ/ygum7E0RZuqZoL
1VnvoV6ZK80KSYRHs6nAYwCRQFaV2qizSxT0HK0OnHHL7dT76vfxSoK9AI21
M0XHA/PVeTc5ASG2X4rNJwsMFDV1zM5ioTn+OFwgV/m2QS9AOuF6NY9R4eVx
bBExSNd8n6up71i+xdveQuE/khSEsaIfiwkhlRRpnEI4H4Bl+qTdcUNYrZhW
ysXOruQ5fBbKS/73wex1IHVSlP2s+xZJbvY0kXjd4y7seymkLDd2oVfd09qy
T6A3eQSy1PiyqzELqqaLcNU7sDH7AcqOGVthFKhaz0J5IuUJ0Fa0O04UW08S
YErn1s5v1hfPNrnBsVykm2hm2V9ECUSu8WI/JcBRywZkKHZbaTyiaPw+Glam
aDwj5Pbmfy9mty7bKvQo7Sn6ks0JXxvvpFv/Q5DQMGE7r/DwTE52g015dZux
rtk9lUl1TyzWNF4iPisWw0/BTLw8rmkL4hzlBakyyPTN0XSLU7OFBIR5+pOp
ldtBbvPJfK3oINAdKXmD/mQKGP2Cd5KOI/W3eYuMvC6aBsLICzD1biqSMjdX
vrHybLVAG9mFqamWr6LXLdMr2eDH5b5Qhiajmq/+qV0ov7MJ4xD+fODnvXpC
TDpq35VwVewUveeqvozGFtQxI8P35lUvOVG1bnnIQzDFX/FftyCt4HCEQwyF
itTkEKhR+qOxp5N00oP/matOSrR5BM2gkXba+UCOOXBLLgXk30odrlpc2dVO
u5nE2CuUihmM6yReUgen1LyAzTQUgyjUZZS3PYvIVpO0zUYnhEF/EBoZmmK0
aWtqiB+SjP6wkAVLDTALRyhXUV1W10HXoPYx9tKsOgQx/e5GWFZqAMhnBcOP
6Sv+CxeCyGvPEA6wjmvVKxRklK3FN3xNFxE+Er/an+cl/EzLwp99jjKsh58r
XBA3OkRNsdKRdo1IIte5C3IzEDN/msSQnb9WQfRDKYElF3WQpkt0Z1Jtlq4i
p/gpZUIFqIyC0lONrsGZzEGTcwhIfeoCRDvyFYm/Dzov6AHNqmUMtVdG2Nnc
FHOyUuDVZ8g3btIInqCqDg23J/Jm3SKEAPM0Mm57vtyD9xcEcXViUz/4frUU
FFUZzsuHIUjpgtYZ7MXXwc2r4KkhR/IfuELfKVu7iqp6BZtormrGVgaznJzk
S0HwKffjOYCHWtrv251eSsRDxuyd9I3J0LVHoYADFuHkV7PtjkePlPHILNJM
F9McjL1VNZdWC7WOuJFsrWEUHO3QhQ8c0NV8BkU5/PrKdHmSKhLAxN6gmF5O
YTMuTJvxroHg6AkC/hDPKCgvk/0q4xwDVmGGRLgcmCN7zHP3UYGCA5xWvOKM
o9J/efsi+qM/V/uN3NeAByOkBkK5LuDtLExzN6TegPLT+SbkDWQSfMBfebKU
P/o1YtxSxZZaxuGV4LgkSdATk0CCkkQEqr9kA+28XIwuezxGvu3JRWSb2tg/
61uazuPN8+v8cyPoBIPoO83Jk3brAGMFrbStjTyvj7VrXblaqd8o1pK6eVYJ
oKRuU5PsM92hCLhzZSbmmJOYMKWhJtqtlgFuyWRp4xlDcC20SRr90pwwmsYU
7u510u2AskqkiYYnJ9CTPovwth88iQGP1Wq7Tra9JqbNY0O9rlMpqqcsvJcp
ygpOeOaYX5Q/R+wjQwr2NJ1BHktTYtyjmY84B/PRX4SEmxbkx4L7Gno6bmln
htnkrxnioVW7j4xleQnT9glFNx/iPN/4zdUAbiomtaW2eP97Xj8TWfHxK1aX
QlB5CPKeX6MOdX8oC20FkiXQ6puQDBhj0Fx62aj7jktqaSoAkm7a+PMAX9uZ
AL/jBpt2SsOSxV8BIKARy7T8qdNkwa5gnbPIU7PJlXDRf/1jb5Wqkjlql3BU
CEekiqQsd2F2ua+VW3c3dljZaKZRMk6Vnfrg5mBdJrtT4TnRcovQSFeeS5DS
FKXnWdmEDYEdFo5NIF4UaNZy3tlowUA8qgBqEvBIOll9OuiHKEBg6RxlGNtW
PkHq9PZfAz2urUn82bZ/n0wOtamDQYgjpACd2YfhHIXiymHTa6XkBAKRs6fs
m2g6JM+loxuy116VSsWvvYoBZihp1Dqb+0F9TLosb03TvO9KNyEFRjclFA5j
7sbX3Abyc9g6TGl1/xuWPDwAbmmi8hlab/MaHFH7RnMu0p5qfH8H+l9hYxsq
TtZcTI3jCrGejF/y4e8MZFVTGU0qNCEcRLi43GX52mAG6T0o5k95Gz+TBQb3
fAfgHWPkWdKWm/tgGqlaK0XjkgHEZ5uIJiIkyOC/hlbZBgNKisFAv/0Fdl69
78iofFxEiGE2c0UUf++B4em34lwAFTl8iSmEAtqdciP/N+/pt+F4xKNirfMM
d082+GW1x2+G80DcB+xjSjwuMoTbHRKeUb4w8UQP3utbC+b3kOgYv34Po71l
lfCkq7I79FKGJ9bOADX7kGLmdvV2QlwnUysKLBL2cXK7vUmLMRhhAY1fr/E3
omWUN79YsNxUOdqmujJslON7wCf6ssqpBM2Swrirpe7MYrFAh9WiKFjX23L4
HpUh4BaKtTsMubJ6DNkI1FLBq0Nz5mkMGzBw/qJ/ns+oPlcTqKawsDlw/Q8n
4xuqCGAXy+hngHokr0tu4jFGdlNO2eCnGsc2iamJwOKsQ2AFNr9XJ6lZHOXm
aDECQ+13udkLxXwA2MAmG3XMplfv/osoLmOIahyRfZdtzc6opxqgNcpzB2q9
leVejaiV3o4BGrQxaLo2C8MDnDGInoHnBefIC3OS0IKXKY6lmCmtS8/K9a52
7uy/3ku32GJaReYSEyVvCsIdV/kLBESMy+XU88O8Llaz5SOwmkJhNolzU89w
9qIfRyDC2ngkU2eEJKKrS/cvVJ/jt6srQC/8NjLV1gen1FIooulQwLEN3DtX
wv0XpG83gczI0clQtZvLAGB0QHXLY+MWoi/vhYiUAtOW/vQJ92D8l/UGS3a3
FGZsGCatrIliXWw2pNOgKHCWv0y1pjf6Je0HIel6ATx0udCpCwhmm2oHAr5L
W0qRtlGBC1VpbGfKbAHsTiD8PpoVYu+/E8Rhl9Kxfc9BimXE96QebPnRbQAh
axgU2S01Ob7jseJoP0IRXgf08TRPe02wDLj6xaP5hwPSFJDm8B/SGY/M/4Qw
uGBhD3FoYoy4byo+Fk+cFi/XdhaYK6nfV6WEYxSmGNFxiwTJZz7+GHd811O6
Yh0J54qUeTk04oZqkpBWDkd+WXJpfLoEs2r3dd8M8oLkabvnFj11dVu/hm5b
dMjOTTUEHRTtzuJgTgJremQ/ExG6+r524IVbT/W4EB0wMrtjC3J2EKvmn3wF
NUofC1ujmQuMUUFJNe3wxhA5HD8KRQhGcLp4AEEz9vSaSBMzNxF2NnhD7sR2
d7icnet3pwLpYLkMlVCGmJT/r3RuWDJCCveRhNE3vZMZwoVhWEDIwb/X+WJE
wDR6rtyMAxHxP17tn6i89SiXtOLq0nNXIsLDj0klXEcM7KqTgmLah0Oi/GqF
JVPU9rINAerl1Oy4GvOoVA6kCMrzIm66sAuDWIW3NfVIAPG2qVnwx5CqmSct
1BwoXrAdGMAihGwPVsuqb5Ky5NbkzMC5AXvDi9PrIpHYfqmYCPlDwyWFVky8
41IJ1FNacS/R9oMqfImuXGKiTWKCBOgNmVXpYEelLoMdMIoesoevXOjbhzMN
Bh6z2ccxwF/yrgG9wVH0k47+DfR+8kYsv3Vweg870LJI92jBh4+P6tpBnK99
j4PihYBd5ZwFW+up7oQrbQCKU+4kjJzJDOzMb4+luBDobPhpYPY0ktJUoTxu
/zVvhLsrkPOC1EYZOPC1KmQUNrHc27pyvpd11FRKyzzcjx3laGJZboJwNkNn
cGVpfCBLu4Wg8nOi6uan29VgJpx0IrAPg98pzHjtJXjOc9hq9KTsb6BSFcOr
JTwKHrHMCIgJw3be7DQDoMDivBNG+nN/5D6tMcUkUgfAkOvSvBYW+iQLWT2b
rq84lV06jM+52wKBJJjNTXdjMfu61kO8+GI1gzPV7DeIAVgrpFKigFEPA/TF
6ZASL5YESBCZAyG0Y3hn5WfsXHkEMSaqmrSQYoGuGw7BB/uyhxh/4KL8+nWg
mG/QIdaTypuvzyzkR7gxzgMEFJbHcmJtqx3X3fdwqbCcy8+bS55q3VbfNnTO
CJsyBp4QHuHEVeYPBpUQXML3mcZPnXHAkbpUChYidvZpDeOghC1C0wyMVyw6
5OUyYl+tpOzS04Nw811IXhDyuV40jb3kk3+m8eGC/UpeEpjyv4iKtVESWpoc
jxiTgODXKbQy4nIfGsnBJB0/3pJ9y0lYzBRkRsbHEDsPxjHBg4+g+IwzEgdl
FGvvNUixw4zXJb5RzZBCOV1UEKwRSX6ZvGPI3Z4bnkprvfSjTAtuKqQ33y8z
04pYP3I245skCO4tFzqv5YO3WpFDNXYEgkCPoW7ogOsAIPrhe7JR/77DK0Dc
Oyr4bwUjqB4Vqa1yFhWxzUHVS+qqKLJM9orLSWBdO27Hn/9jVzIs0ZqE2YGr
JnSdVDBUWkiJRdntnwmMAj5tEWnV8/uEd7Wqjg+RDC5uo2RfIrvfT+OJ5m+K
oNKpd4CUZLbFKEbPfsriJEVd4S2CmEFgFiN43dCk6cVCnGqxKv5OEc9G2qq+
YLIMoI+H83mNbTD2c5pIoMooJ8Vz9SquZzP5F06f6VhrrZfpAhu9GOjxvuVu
ERTEc9t1PCJ60DBYE3Jof1ifluWpteQX0C+N8AbB+J/EBRy/eZbbPIodFNuK
Lny3lAm71OGZSnKGa13ocwuFr+iP2lXo6rVeHN6TAl87hrH8Iv6sn+FZlx5P
9qg7K1DtF2Q5OdOwG9jnvylEnonxAV1GikwNmSb1rL/naERSJYvjhXiudpqu
Uk84eNcmlXFw9XGxMzM+w8c3XCV5mgwEuEmyVKCbpFzb16yKE51R2epMxrWJ
VJPNwYWp16o9iqGBTbV5jv17oGcd4SRCsAg55O3FB8niYCOweHeQT0WusQLe
3spCihQQSNPsyUMNtcK76XetO4nirCd3aNzkfuRazkjCmQfVfrQeFIvA0MWT
vtoAanN9kwDkVAZ5FhRUCmbaZU1ASoDfElCdEgwZigkmwVlalxJTO65nV99+
cDEJjB72VMkkldpiovhhO9jn2qPM1zlCdtsmDclbdFlySLoVZiTh/Ff7zuY3
PrRlzGmtVdanxEgAa+Q6Adgl85AEpccE9GDQF9PtcGSnppWAg3fQDXuNTN0q
Db8tx/YoYj9pyJcGQn2tlK8172hDeG+X/eZZg4IOdw7ODNwON1w+uidXPgiK
b7hbPS7GZBjvTKmGZSqrwy6sYBpFbJogsN0bMjNI8X3HT0oyRKT4/0GsVzCh
C2Qzhlrrih5L5Ozt6/DS7HiavaWumNrh7F5lsNwYZe8Y1WN6PSOxKXFhnfK3
Qr01iZ9YqcEHM+6S7Z5tO3Q8TrQgbI3qSOBHCOrjzHE51iD2A6QHJPQyx0a/
aSqxOvXgL8ayk0aUuNSjkzKte+7HBzwJukHfWxcUyr9hbdqxIUpnXCzFz9Nw
PHIlAGyvgBITqa6v7yQzn51DmVBrwKuj0wLT3ju9u2IkSIdJTEaVZ2sYK68p
7toqG59gnFnhW7eiiROcJG01j2EtZSRhJiWV3Ej6lqyJX2dxVspQGE/Ptkcy
GEuvNWJAKS7ux9yRYeuPALha6/0bIFfRp9cesgtC3oppnFJi7hE2MK/CvgqE
D/fH9r/4cIG2jgtf7f7d0aFIP9pmed8+zSe8z+xDqucPqWisFUp2oivwgK1E
fvezbvsuRnAnC51vRLUpaUpcPjyWushkxfFSKZXwMtnl32yLV4p7MLCd0I7/
fr3Rj4XaBhv3v1ixqdGCHuV+uT90D1qMr2Kc6hkz6KgXS9tmUDqp56+sxI4j
qO8pyHIlmwIV6TCitcA3r+WzeenqD/mVPOSKApSWoy1cfpZD9Ks0TCKqpZqK
d9zlPB2UcCVD7iBFazNEeqgIWuhRucqrvO4y9G+FqZIrgKWIWP1mlA3/U4KX
eELYNc61JNCaYVbnYWSOdzQAFmJ2lpisnrjhqeWquhZVp/GwyWNs6reFReZd
S4rbWo8se1JCJ+OZAr2qFVYSrW5QpE8Hbr+Vev8Rp4xBU9SLGaGySXr7T0p9
gNa1xt25dum/rYx3wmBBxX1NOieGFf8HsZS9/b0Ep7zVXo7XSGxHn6dQw8Dq
8EFRpQMR7DcrRgFhqg8fkEurRaeahAcagh4gaZRY83yJrFUZ4kbp2V+nr2xY
jLFWnZy3S1k+aTmdTLaFu2pTfz2yw0ssEU/6xpIS45gNG3Kd9EYFpnYNKD5/
5sBvveB9dxbSgIfma3x3HIHWcH/dpvrBHxcWQ4tRx1Mor7Z5WYruvbdaRnyc
/Rew0X2up1pLAPwF+M9YmPPDk1dSelJtPhs0SIum8M77UbB9hnnmjS5k7Zmm
lxV43COXN4E4OBdq9L0eGE+3et1AU2f+NoqmeLtrYHg0vD5MHZQnspERP43L
OZh2KpZ7kpvtXEGyhPXguNIEn6kw0E+U4auDgphwNX+Aar8GhGd7W2GYkbat
V1bFDgwY6WJUEzHl7Z3pSMym3jZPpY0b0OPlIhHG5ATvmKWMgJxS8SGP8L2Y
GE8b8YxCQE4ejFeJ9YWERbGrZ0iMI2CvwLAhGu5QW79DiZrWDmZGLK1EoBus
25d4G2wFGByCxXRuSgrm7WtEtyGak8tGKixABqpX5XNbSbnXT+YyQjRYzlHa
sPYt3b42QLbZikojriAkD1PY6Mdbe28V/Elmp2zE2iF6XOi1htlefBPK0YnN
skfd2ereHVXXFFLtht6tCYPEhlcHrOx2Eb1hojhl323eFObTf6u4sJoFe3t8
GeHSqt/yKZ05pIp1d/SaCfrT6oFnfXdPjJjoAgsojpumiTIGhe8JeI1Fjh70
DrKHNK++khhGVVIcUacqTiA0qUHizMbMwuKo5m3OvRwJC7kGwjCMPckQ9483
qABk1Vsz1O4wZ1sncILVKzTQtdwkbl1Oa2S8fRNv2afZQCKKwCPxsfaAl3ui
XQkrvzJpKpM3+iHj5hyiEhlQUlV09ckBbF2MnIMWVGtPvgc3m1Tez64i6u2T
EtZnWU5v4SM8l5e6D4mROEoP/jbQkTaBz3VCsxtzQO0n5cSitSoXhTGxr3ru
8l49OA0dDxsm4r5lJgTTOYCkPrU/PAGslWMCAh3aFcN+dyWa3RA+ISvfXhhi
YpJz4R+SHh0h3nKQe2sGomWPNShWBwiH/kCvW+ZORgEvJdVJOVl1BXkk9KHX
mP2y9gn6NBFNNeTcS2/YwS+DGEOlpoe4FLvD5P/YXZgmL6yKiTDWoYXG18cY
n18CWMAeFQImX6Ze96I64tTPdD8JA0WDFI6jVdZRt5GSGyqG3OKCk4J2ZidI
us3rg9cvz+OdsG0zcGgHln11Ew7Bae9iqps6KYdA7BDeuP9KPJKI7PaW8Plc
dSBcXN2uJt5lbK13CwL3n2CCYkAEPlugydIHzmLNRM7hxpE0s7xpygHBqabi
K/liYWaGKn+1E+KRZMONjtWPb+fY8l7DpaVV/xLD51yM4cn1owHF/x3ktn7q
bBzFIYElxsGfbJj16PydD9P/wruoUQWuvlMyFpp0l2hdtURKXsx/toGEdvY3
JnbrQS2/PKYfWU8uVfzcnxnNvf5Ejx5MSxinf+BNWcUCWoMW2gJh6sbsHe/d
wTEJh/8mBci5dgaelzwutOfLSB53k4PCMJ+9xdmZZy/sYoaHpOIfYPBgJPtT
i/dzihZAIz+gb2ft8KUTaL/hIrEXblvOsKTS6FzSMJWcIYpdgJHqtOiX6IPJ
U32pmEmiRt1ilIwU9MUMsLhOjyN3WNTZtiyE0Cy25Al0Lq3dMi4p2Lwqz+YX
CdJKKWE+kJJZnfDVFwviVQXKxN1fvXgvihoPPBKFYLp5LwkunlVh4YgM+Wz0
5YJyQF4GIaNFmiZjT6/XtV1oop3450slTjk+pPOFFpJqa4SZIecmFW+KkW3D
MaUI4L4DZKNaCNFA7KIrBMd2pyG0722B0fnssQw0K0Vow3g0DjzX8n0OarqO
N3IOqmNf77MFw5+tPM13dNTz7Ra2eirmQm4o3hYvXChq+9F81Z5OhAnlzi/N
zZtNvnQBwEEbPt+Z1AjKPrPlFeH99zNaJPoKa5BS3DKW5n9OLLfFB18QROOo
2guwUINhdgO0AnwMms7NBkIVvnIUXYF1U8jDjNx81k1/ug0mOlxqYEkJvREj
LjfTJKOEhf494z/h+DytROykR2HaK+SUvmuzJc6RU+syaY43UGC8D2O6jDpH
jxBFT5P+/hBoHM6L4iG28Umo3UiCFGM8fXLW8XwWjO6Olt1yZb2RztP6Aedm
DIbwoU4Wjn6fd5fRPareH1TqYyirgtqaAV7LFPVIBGi5UvGCtz63PAM05pPg
k5uYKAxavPh+ou2dSwoMwTYVIcEgc5deU490+TFrCaozi5u3+ajR5be/5Cii
rs5YI7tISmC+KO8dhncvnJMVAr1QbhOb5BUsBD29k+/pYSgCBs10AUdGnvP+
aw17rFnI5UUSLWEQaBOE+t+6kIN6l0lTg5ygupf7Vzu7o5wLNb62y3AK0qJW
Pv4hQcYX0yis+JhkPEojMuCcfOUxup2RVo/YIhmXljsybVScygBCU82J+bQB
/k7UZMOmRX1jGp3zl7KiX7S/Gtcy9yC3LU4FCsqFcAq0wLz2WnybqnOuqb7y
MsTSM3gQXVTlcW9DhMCSDtUwT7Xt2Ey/HP1UBUkmBXZRTQInZSAevGSS1k7v
s8JGVSmR3c/Jr0HdNwWWVmAkNJJGsadtuXlh/PiZT/9bOyeX4/ifXeHm0RJp
GKvXOCCupHHPj2FwX71k3djnOrfxf7zm1VkhlCvB8ks291HGbN+jFKlH6W15
EmqDcQPxg/GjrobQXQtOhMh2cgn0dnFF18lxa3peM2hDX75EdBlGexmmjgwL
k9gj1lOhn8HhLiLqa75PhZsi0BxYNLX18CyxF8MGszur6Ee0yF47EhHjBwxK
oOqyG3NdiFZ8558g8Knn2ywW4jqbZD73onKqmBvgQ6qRyKUqZUokWuY5Gsr7
0h8Tdz1ZhwVaFIvR6FrZsXaR0f/+96QrZa/DF33AQh1LGBiv+2MQWMkaHeKP
TWWwMUg65zMlI78Jbax343uh1yYOwIJkLm98xbn3VR6iltazxgO8OrA68yzK
/EVxVwIlO5jbQHfpoAcRBShIEFkW76znoseT15lhIpluNlGqXeGr3cieHRzD
jWCprayfHlZ3vMFVniCwttMhZ7GMYTZCa+57nW+KkW3N2IXTfDkptnSsBbh0
IJ6pVux4lxGFXcR1dvDk6OF1ToYHjXNuj1BQsQ/HVdwU4AIYRWBAAQv2ESJw
V+JfL9haWHtmLL79aRFGCtruThyPWClbO/1iFS9+wtuPMtUSJJyVgGui8uyl
Av5gbbBkUO6mLrNJyRlKxqugyCksrdI6ixq+4o2DVeXchWX1AtJlenac8rTu
m88E0UhWVKqa+urFw8ZS1uKc37T/n2vsh1Z7LOSM1SDWRxkT/y4HeK1rE0Jx
rnofSnskkvVMPJGsJTBryKv+dFv/osHVs40D1u+GMVc1yk/PvDXBRfOOgGpx
dQamM16uorFOOc+/mwdMqoibckCOf0QPaKMpR5cOEhSaYZ1tq61JsqXC6uVI
JoQkZlYHTT0R/foynPeHdfzGvowpuHrteS3Tsb3pmyokdiUQzu9yBVut34bQ
4YoDzLhQGs3zmQIPHNhB0d2nUWgxGsIJMr3dviDe/QAk1Gsnc/cyjFGmQREj
XYRaxh4nTQ/uR7krSq5K2GCV3+QhWQbrwYy81aLprcaNFFcD/RQULt4NUFnd
UkbckcLscw5BePHE/Ueu2JsEKiq3t2NL5+A/4x1I7aRfaYHF74s/DWa+WWAP
T+3kuAHXDHbJ7wWkoMpw3/YM8RTnj9t0HfVEwdG/dDllko7kObA7oTGYTZlu
l1YvMWayzXODjQWg9a3AJUDIW8IZPKuV5HvRApFrgxj4dIw+A7xRYYg5YGFE
oXwm06V70W3d71vrKlFAZx3N6t/ixP8UFtNPzYf4zIwxXap66+ZJfMTWp+H+
//a7/CEpA7y5ie8nt76hzwckdzSaASItpg12kUYcHcNze/RnMg6YpIavkoEk
iuqCboE+I49SLWaPYYjdq2HXH7X37ylqJdcAvmOMNF1h0LFa3WgxCMHbN646
TNk33N0sXONyXmcBP6PgC9bzRyF0Yd7BUrUIRfuYYblnyi6xiFEpCqQggis1
Z06OaQtLavaq7SkxLJE33extoBbcM5mWFoLXZRm87FJNN3Meb0n9Yt1BSP+n
ajIdWB1vIDfaCIh/kyJc63XrQP2pwyfu2NZ6y+VAvx2lVVmQyH0CoYd2QxOr
1lMUnIRUbdWUPz+4kwr/grtoyRQd//PGtWHooQJTTC5offk2CGrqMbdTEqZA
21QCoSvR4JifHb4OVL2YAi7cd+I8KhwQWpiZyoyIwbyuSdOlIv58inBU8vyT
jzytYg5L9/so1gAi0CYP7b/6kUNS0RP4HN9UCaXkClHHT+2UfM9B6Ov0hOM9
+NUsgJShRkUglWODyHJQDrQKf+de9e1MKLOA8r5Vo0yFl+RDVDqr8SNzetvH
+tvIl4ZorpGrA1fz31i94sySyFCDZhaz9mMi2JVAatT8KB0qHTbMSBWRun6Y
R/jaMBzjYEtYm6gDDMoMgewH4fy9kiRrWVyyDWqU/xnG0PIngIEEgMtQATNC
1aVGKieYc0Q/yv0m7N6dVCMEfdXWPiUZTsWdmvtkEAOOe0+0N0rAskqrvZwC
InIM9qB3UU9BIBi7TbMlnf563BZbcj1joQIWghVs7WWh2mcYYmhcVlcSTu5W
nvZrpM5+7m0kWnyghGC7khVeUbusAnVEStrC/D1gEl1ujvtSE5NZE4F4XYxo
VbKuhktLQ7CJ4pN42wSo6ttPNVLSqm0cHXdY/I0a1HJLsLpK83zeiRJcfyuH
YvQ3iudqIU/ShQXQr5cQyxm67HPgF3mHFSfxZqUTHnzTcrMz9iS9nsuOpzKV
bUHMZgkbfASmxZQz/Gz26xQOoia40nntH3BWXGiqqdKQhW8Vz60Yj0OQzU1d
OCkghsOAs6LwFkvGluKXJHKwkpKy5Cv1ImJb/F5m4pC6QSJq/XwZhNsiGUT4
iqxp8w4PDYgV6dLJPnpztH/man8FvXIltHhVKQs72Qqs5BU947Sz47WVyyn0
HrOr9gJs2dSsmxDbNgIF27UZF62magZ9OKF5DFNXxUJwxfgQZ1hbSlb6uDJm
2Yelb9Rxek6B8WQZVyA4hrJH2wIXjxxBqh2jt1gm9wN3qubUx4XnkZu9imRp
poFBjSFyFvTGHO+39KX64xGb87vewvgbl0yPeV4at+JlA85xThWpKF9jvGUT
3VmpUz8jUWwNX6W1O4B/4QwHnvLt3B8vel12y5+2ir6YpDDWbramTA+T9lgS
ZNSYlcBSq9spgMv+0K0PtVNwmO+UgoGIFuvTUD8kTF31q39xNoRJJ84B+qCq
ex7Fpor4t86x61dZnt43VPW5d8p/ntfc1tQ7qGlOMiShQlyEM8P//moczRfH
AUghdzLAs84NZVjikvrnwhzqjGyaH0bQikfrgEbWj9MOlHBpS1PoeoZqg76W
tiI0sHLkrkflh62p27NH6P43MEma0M/PVrWlPU19cJByHAkSdtRe0RYfJXkt
EXQAoaxzkoWcR8riRfOgMb2Cm5VcDllSiIUAvRVr+i/PwTb84s+9Sl867kTy
KNe8TpCo/H+Z1YBkkdeueSnjpNpXzm7/k6iwNCYuvnNSnGKQxz4h0/vXIVCX
lOZQsoabY1H9f/rA7tXoyfMyOs6n55Cp/nc5FUIlsjweBuCZ8VpG6JiZiHow
274yUGPykcQZWES7sMptSH8lJpTggv8oAGUoN+/aone2l9ODpqgS/EKgX84q
XYO+nHsRFhK3cJDBvmMSryAU3DUqOKPMr99GsqabxjNXpvbhULU+fz9iqE1i
Esyh5Bua7XaFtZnxpdTgI5FGl05fT55BmJYAIxH9WdCsk6nXbHPcxGyU2paB
0gUrkZv3jEw7hXAiMnmc/+KJaznfNJ55OQgA+wyYHsJSxuqWZakZjtgmk4No
fKTokVJCcH9ue/sOigVfNXTd2A/L9xayim02wsdAtZz88jOXO6PTZSxTE45x
32Zou9bZ9FJCRnDo962/AsgKcZZdXO2EBMiVvESIWfp4silRstyxwvtaBFzP
3Q+6fUUcYxHkHGcXkHM/6LlKUxwlBH72JtZR0xQQUErqBWjly9KPdjhuyMX5
W8ri9EKubaoyMhQZhAk1LGLBKW3lUK0uAb8/jjguimC1Bcb+rjzdt5e7XJ9W
6HDOlOJCRjFVr5/EEOUCu3RABc6W2r8BwM5YfmrAEXythDs0EZFT1cyrMIV0
yPvBO6V77ZFdUo67Wi/YxvRoYg2EsIQWziC36PN+A/pfa7gaAtQVUlUhI2HR
Y0IVX+nXWEvP0JRZ5XkVJJvNHszMdxePrDYzHwj1TJqke8qHeX1Y/584hvdp
gqzNNewB4ylRcOsvzipli6CCnugFaL4ZpG4Go0rMwAbibVIYgpGn57Gf960k
+hNPjMRXLvK5wdE4Ck3tVPh78ypWBl7bfq7jtdx3r3wwZML4CBUqvdLifSJ4
xHstqYt86pb8+EWqwVoqJVdeTPg8vVGp1Oil+n/0jggg8JuKLph3gdKw9ZU1
zZA35GTTgCwkqThsKj5pSI77fginkg9W+Rc+QRKLp4k63cbVVZKluLKoUXJy
wHryapijUdJfbZGo2aA/K0CRl4Ili+CPSI8ghjO6QG38OqeXDW08+hpvpQHe
CZ7x6N4A9sCgYJcP36UbLDx2MV0bIgAPFrOPfi3bGPa1n6h+ztQhygcp1AiK
VYYz9kYEnBF0UekZwtQLlw0hBP/EucIIZfJ+o3YP6cLX8ZkB4OFScm3QQNH1
sIHc0qRTDbAqRZwGsD2VMTHo10rIVyQ+w9ufaOPWucjq0V1I1gENA1Y1fEVf
iiCrcJMdA7S6+VfB1n0L2ZHmw021OZcDrbYdcITx2pmx7tqd9kzH4/dXblB5
Vd/6+QDghKlEu1VVzGWG40oNG0uZJBJdOwE+wb4shaQ4HAw/KBh7XD2D8Gnk
24vVeivzmm3tjmHAQ8n8Z6TJ6ob7p6GDycg5qgEPVJ9f+o/Rek7RbDY+Uf+F
11J0aYIwIOte7bKb4vT3ubS3GUHHr2NhZMlLX+74nK0G9IEMMy3beeLX8yaX
KEZfehgwI01iEp9HMBJD1zwSq0umCYjj6KoEQUi6r0foubzxzabGzie6Ugex
zL2sKKZg2F7LtSnU1z6FfVp3jy7bqJMlpeKm0fPqQ9Yeth1xl5mxfdFN+7DQ
DIXthS1tuVFQPh6ghZnZN+Koy4IOjCq3yJd/6KUS+r8ZVoLGyG7+UG8w8rJo
t7r9bXyLLObK5zz6IsDdDc30ztLNY5lYDxcDArf9aRD4uQrdZsiDTkCB6Z8J
on3vmlUnC6mtVAv5uEDaXZV+6jWOziyGlheg/UuFbytIYNeAlq01zuaqXeE2
KryPSr5bhi1TpntjOtK38AIFF8RUFmp6Sr3Yj67EDA3hLSCHp7/YYG8WeuOf
uE5KVJxUroLiMvVfcq69R52SfDldyE0avk3Pb2kd7zVwrVPe4W+Cd7wiqrlV
kp5fL4RveOxF2S8ndvdtHr8klZwNuIK7lI0qVmqwHTj3hfF6M+XMjyiIIgCN
BD8JMYcedyhteT6ADkJs2thOIzwgM5w0yBnBMT1hE4D2cSQhR9TKyiwmyMTa
z+OZ+qJy/Fbn2dYjby1cQeoyT6cvH0RuWFfm2zx98RwqLIOgdtCUxgaDTx2w
1j39hZJ+C+kFz+y8bL9c3+padwFyD7ANgioVti6GHlDxqiORmDY+mVgAUC80
oXPRoraNuEC6is6JwUzTJvZ+mAtgYiopkpEQJiyi365WswIQuvQltbqBFzYD
2zMjYKD52RPgEw+2DRBfFkwv1uRwWKy4o7Qq/dz2DWwnqjbLLpnnv1fVs96w
kf361pX4seqDRMBiVh6L9Fh+oi3mpDXpIZcA3CtjZdeeb9VC3dEzvAZhjJ4R
m51q2yoezvtyxa6vTBmCw44feuDUvM65y5APRzdAcvdOstHv4kExv1NwlaUC
eq1oqKCZiHE27ac9z4Upkhl67UBqmfWuDRCLmna/bofyah6EJhYZzreujJoW
imTHMEcMRyk31XLCfltioeCnSBrFAfmjzYz1eK6VIjKChUoHfPP0ESa+bobA
FlA+xiCAMc1PxDSt9YL2n4/Gxhaq1/D56snYGlC4IjAiEPM7lxhCpe1FUiQs
Sq19rHnT5JyBrL1UANaBgLR1tYN0i74gJKxQCn3UK6XDJ+VEwem9wta/Xz3P
7uagpXgr98BkZ/eq7CHGTnTqUIcAMErXtTXY3XUFGNAgAJo4ubYRnGhEn3Lz
TpUMdKYDW679h2TAIhkmI6VGP+2S4kzIiZMnpdb0ZiABcSVQvYBrj+bSv8+6
ISrQiDVyaA0CK39bcFvZS6EdP7d41RqmBtneeiDhXCB0yn53Gh4RYni/3x+x
YQZsIXfCJtlyiLhsV7MsFhGKYnRTGKD0+tfziiZ751fbklzFbqn9C/2r1/zT
vHHjXuRffmXvsC8SR5gWF8NktjX9oV/SwZwNLb6oAKZjHCS1609E4IHC6wZQ
EQTP2g/eLDPcCqy0tIIP8SZim1A2BTOwH8uA8r8sC5R4F4yNAE86KIIBCy8z
EQq/A3MTWrQWzLrlcaJwtOFcGsNjxgQyMPNcApl2rAL96ZvNjcYQVUJgiTf6
doboDjA5U4ndG742JhZhZVVxe6v0ssrHN1X4drXk1T2AvVat8wONfUVstops
6oWGnPAJ3C1VA+JoMeZTzFyEvk0IlCKUvMx9NeWOPVy+3hdRkLevVzMoK/Wc
OwqlelHZ6DWlLl/hBSw7/sZuhQvWvd6dOQw58ZtKHrye7W3wh1cTUMUUmKLp
XYw/mMFyRDWd9qd6qgedF3o+jMG804u7Si3KA5g9cN9Po592DU45vAbpyrlo
W6Q6Yy/WYcrPkHpsIrgskLaLDjBPjd6LN9lvoSIBZp4uV9FBpNBi7NDuDfEx
csp6V49ALA3YycpdA+n80DQSH8I6prgKhOvyjfo6rxvo+1Roq+nNed3+0rrl
XdCwVdZm4NZPkbLgrTp+EJZHLB4iGjZ0HgbrV52gxSCp39WyNW9oIwm3bknT
ywmBtxeudGzhSz+x9cgeWBNWg2t1LRBlU2LEAt+Jf0sx647EyJdXb64Tfcfj
KU0VHKRTVJtDnCDeTGReP7RPpSp+AQQBocMpiq+mPkGoVg5eUIFegAZQezPz
HxS8h8NC5M4vPZIEBhM1HwxNCtAHJgrmnmBkvqdhNMxPhZiBv2U2xarHWSvT
YMsMYqCm1ZbolDFiA5PeGOCeWsVx8/TeQypwoUt+FtFtONgYM7ItLQDo/Aat
G3k4L4b8SGAMqIWX7sTi3Eo01Xg7YnAOkbfpSxbi+v0f9CnhV66vZWcDJfI3
CtcetondrakdM4LW2krfOvKQx+rRR29aFw3xSvxsUq+TS406XgOG18+koxth
hslN8LvboNtox61lpQmFcluZvqEeS5NrHY0fH84BsoFAwzgtNmY18+7to2tS
KOaM3f1ORlB0a34khULN8GwnTdvQHZ8Rhsr38zTFzMRw5R7WjkWgaRpyq/bp
pAv6hGz2PSL5ND83RpwkbYuKj3mJQHpoL019VPnvEn/uLwiX62jZmasRwJRn
03JKcCOUeSbCICLQhjzvSc2+neQyD384M25kS0teq6xFT9ZlaOAKncRuyq3G
SoVujzlUEnbuWYqb/V815lu89b1hOEZg8GbBp+o7RvvzJ821bDb5kXpAtmFL
bYNC9rclfjb0gT4Whru3aSXo/qGKvWp80k93lHqwA19r6d82VaQu33kK1WhI
+222hoArN/9UaNVdPJZWo1hVsPmIEdg9VlhEDxXaFUcjb0QwcsIhItoPHsaU
MlFgs1AuoXZ5iC0f0KUqb0T5mivMZGLRexwOcwIMky6+sF5OcPMLE8U9ZOMu
uZMhO5LZPbvJuTcH1hRLn6oSwLHH7dBH4sduetYCxCNrRRYJlgvfykWUixbO
svun6g7CUOrrDsbCN8+YsYvskfkXJq8uJ0OAMCWhBG+OwsRPE35fvZPw3sTu
oLhkhFQRMHL8eHk+SMLfmM/4BpYWfT6iZNZD1E/IpFZ3jdc1ZumYrHeKNJ8Y
Jaz/HLpR1kuhvF3uornN15CVekjmtav8SoSLwi9jmqVrsYiWIF6AT2X6G1sm
gjBEAUxpLGqp1XTOKt91s3rDpKSOhrj7EeDBXFN3Ww9VAe/AEQ1TuJFx3DA3
Qa5Kuvg9RxU9LS3ARJj2eHoE4naYwzmZZSKtFKSpmfuNTXgBYWRZysi8D4lW
3AgUi6bMG3enORshQ/SvvWQrSfoC58sAEpCmGDqSO4g+yYNv5vQjNIfi2j8j
jtq+cQep7bAQBQJleh6yTOn+P86wPJXE3wFPz3OFyoU6AOgLvUisDR1Td7vk
pSQal92umiao/2nVfmXfJ5lp0QOvUZGZMoC3QrRuA7iJ2cBbCn3b3EBYzQyA
npY9HSwJowiNwNN8nkorMglb1xHbd+jph9eosBc6CrqPNYU92H2Yzipu+qoY
PevepSLH0O9hpxySFb/a1tNZIWMyouIu/wEaFla6OdqpcCkT0PkBmaMPOD8x
9teD6AtDRbCjgk3V8HLGFKylws07J1PFOJqJJJDNt8jZ019kMyunGZ/KM/uu
4oBSW6Gbw8W9KvB7GttfVcf6Q8FJ0HZ1biQB7J3vhZXFa17rtzxY/eXQc9Sl
BwFn4M9rVSP3BI6PhuwJXPu6AJ9B7sPUwElbCIw7IWGFRd8Y4kT+oyWERVvy
NP3A+EIsCMwUc1tm/xJ8E9YhDVOE+HtgqKqPJ7UVCBgmLWecPla5Qw+t9oY6
pkVo4DIloWV8vC0SMuvCRqrfkztU+x1GehfQuHotHw235ujp2AF2NAGoXXC/
cg0WqqcyaystvDUKHucMflLl+L6Z0+k8X76sY0FkFeDXD/b3v+o/jbABI+PH
MgYGKe/nJZ3J4E04oHL3vPBBuhCqOPvmEGPcyVoYwxYQpL8dE5R+SV/K/Odu
IIjtbVGAqqKJTPGrjHnYylD6aQTmxxuXXhzL/sarFo05Omynqid14kWgajUd
dzLb7CdxpTgj6mh8zQW+bHEVjFPVcatyj36CMwD1i4K4bjAavQNkZksQloam
NIPKLmoC3qvV+p+iVcHdyQ4bV8ym6SYdl7HtootMewrrhI0hRoVuy8MmcdMh
bLqPiGT8gJhqeqxwEwOMTmAlvKTxXRnsrsuNrLC725NNZN6rlP4+bswQUvGQ
1QuPzGO9AZLNJbTtBYP3J72ibA9j2t9y0rZEp3KxRL46eZEvc/N8PDYX0iX4
8DXyCzO59AhO/fLZUySJu5mB1H7C5G08KlP+8RrZsFAvzkMdhF3bmeWvqJOD
4Z4rBchkeOPIcBeI+Wj4yESOYrI+biLp9kP//pXQiO5b0Mi8JHlLjmUv/Zt1
huEM1LkfTHp1H1/ti6IG0aJuZdx4FlQugaa298dPGnO7lxMzui7pWbUuVF+3
dbzK/2UgZieEF77lGmfiELuCjEhPAuKKNbwR66VmV9YfIElazp8ClPgJ2BMx
3lAxR40k0oeDJV75aezgYQ53uy/U2919Ck9+Q1VgQ4ZjkGPMyKvVsuCoMcmz
q+HFZcuX7QoOWrx5CIJZ9w9rSDn9kvcr6QYUTRzVpdQyMp+KoRev2d2YtKkW
GkAVQMMfNN0WJaBgXYZSzw0Xukc5LjnDvJlhVZ1LLqYeJxezGU+XOrNRPnHJ
zdUVIR5qhwvM/aS1EoKd/t/uTZkXeOZbo5XKD36Q9m/Z/kGpD4J5qf5VT58U
KV6PKGkleQlwhXPbUphRsBtdgJnCcRwSOE9XO4BaGG+ps9BWTUyHrBk1oRpd
2mJVNKMJ/T+LmL7qvhR25+wS33e2WdyVcs6wJTU1FilElXSWWo4/c55nm78o
U2LDv/LjQE7UEERk+AUOK1FI7udt5VFaOPBlZ5oR6QR8aHzS8lPoc7e1vqh9
fP4hxEvNjc79i1kAP7AOHKtgsjlzlmUHg8cy7AoPE5Tger40ss1fPd/5eYGs
bSWXtCbCc1W/lqxcg2xXciiLHFzyTQBAVOm1KWyYfqrO6oTg/r8Wbvf3z5T0
h7gdckyAN7GBfM7ixPh3im7xOcwlXYESrBW7cFsiHoCZK6iTK4zyGhcif6z+
5DYsJZyj5NF708e6puSCX5qDSGZnJ1rMZqPrrUtoPL1ro0y4sOA/kpQxggYt
nE/vUwldXknO9L/J825IUBjNyvikUrOhJZtzrI4Fc7L9NBfZbTNt1RljiNMv
YamiqkME0x/Tlmm6TMTB96C5rQJT6sdV1irExtvIsjGuWk9oAViloOLdKg6V
yDdCvv1JohLhAst/UZ02CBxfjYTsiZtcI3ztN0CXeNDyJW5KKJnGRfPTC6N2
MYpHqFNw3MYBUmAZTqwwXww1H+wubW41FbT3s+Xv2VD7Z/4EoYIaPss2Wehu
mSngZGmBd91hiruoIbwPShmUMlydmS+lbIITm3eKtgnzV1derFHKdVtu4UxK
0PaACYMuKY0/xWzK+d8PQ/daZSU9aPiJB1THxVUFr3WIKkZfI/1ea2+/dW1M
nSO+Fx3qRYSLIKvDZ/bGzEiKFBAk0DRCPD2flBHfK7ypeYEthJDTvJmv+MMM
SkA9m222/07hDJ7R7cGOQ2spUnveq7qCwS9KhWf0mnnbMzSBfiDGxaPMiX93
aN+anap5ruCNea5ps2H0Hb/HotZr41bi8nYOlnN3/WfSVMIYSBD5a+1yyRT1
/xAO8ROgKxQVYuQo3cF9cXI+k4HiYbgt7CYHidGwvm8ZZgCHgmpLCCiQqVR9
GfN28SGKVBc7qtSLBXcIeGy7/B8VnIot2twBzkoVqRHKy43E7HnqOQ3ZoKEw
xx68mzlN6jux8ulxJK6j2uTcEq9W1OIzsFnA6d5EOgzglPsUZvOi6v0rFwPa
NDdkCG42b26OKV/ivLN2GPM1ySH97PDul95Pb0AiKGXAkWoC9anSuZsxYDS7
lpW+ZYx+zlkvgkxRznId7iW4Z+9mfCOXgee/PQBaoiiN2I3Ae8R99LIDAnxt
kpgAEISjUyvVLbTwddp0Hzw61gmdrColpIRI+NoTYYP0HZqJ1ga9G5901AHI
4p2MskvKtryo66ZHetEDBxNaxZ7qfxQYI15wKedrX+v818oRnLMBKqSbSvBe
AVfQs+WYJ2Pi0L0xpvNI95a0joPgnhRq3k3wqbZxguANUpbrxYv0Zcg/c4XT
9qcFNJcgQlThvXv8GTMCHOmz7TfTC7aC7cBLnLAWewK7pxuAlnEXlDQw9d/e
1Mx5tUtE68VJQG4vHfrBMJ46RA8CO3wZBytSw1Kwqz/cpeFKyq+1hR1Bq7Ki
6yK+zl7g9/EgnrAEtrIfYbziJIizTJBogqeTDUN5+r3whyDlIiDLIicaBVPz
Ieaz1zl/NUfr1kiPmdlrYuRWBNuXDzXCe31rLcI9ZI0tR/Gu4CmkiAZxHh5B
UgP6TQCueoxYrCaztmRh2TXa0dKGtX6pWnjUvCeHWloH1FA6Yj21hRORn9c5
VOc8XoaY4UVRHvgcLJGEfAuMG3tuVuyC/kyzZ/c4PjCb/Zt22KSyVWXnmikk
XPYwOkm4tysY1gKIMXRLmTyDFOc1oUaLnb4VBcg1EwXUhFydHXPUxMwC4K+5
5MdZ44Wlt2o6SHMHK1ROgStqjij4Y5otfWRSTUvd029ZoT+OcOjSwcDep4fo
HqN0GtSUP4eTuUqDhuV4OLdHPoCM/Oq/2AibA5dVbMi7p5XJcUoiJkFT3sgj
124MZXIDLQ0JCaT/hdUFw2+GfGjbv7ArorAONncUAB3gSv2ERhHpgALOs/aa
vTDN7hEkRlEQjhwPhXuIGB/E3SzXKKh/JzzHcWr2jtKu2mRjlqwG/3qzqZRj
X1u7A0AIqZCFAbQRUZOaqqa6Dog2jWU7v/ngJlD90te5qyiSIvhlAKFGZ9ub
nRAfmhliSCwCDUis9par3ayRlN69BKBssxtoOma3U1qgbqtrgsH/Wtoc8qiR
QiXO1k4m2A2EJMSF5wnkB9h0i4WwzxI5a9aDZzaX59hZzeSwFvwKPEoQ6iLU
23eCjz/840eYuIEnWGPtUSzcmXzdhLDuKKo63f+H62aZfBhivvgIi1KOBwYF
lvLuhVLw0gCVOWL7y18Bay5ak7S8hCAYMJ+XxxtZemSPSb8Min+Qb/NQXK0V
m90tE+Kd3y222BVmL3JfjC1f2c3/gqEnCNZ3jkXjZrfHGh3jkorKL14am7Pu
1Jlpp1oYyk37J6+dqOgJFopBt45hrRRLVAonwqFrkfFWKXABmKS5a1dmZKob
ZomvegmR8hGUfEVYN0U8VwzNUl6w7aDjGrH9K3YRL4V25NIs66iCHx5JIMxM
+S2vqn+hOIPIB5iWD5CX99pguqoq1osm7k3BokZ/PGYVN5cTW9mljeTuXnQg
+z5GVYaAEw+SWDxEUPQZJLpDtDICsmVAoGEx6Q4DwwcgH+Rp/+JgCdv0AE54
nPJa+wMX22WhqXn6GQSGitK7GYHgM29nJ/xmampeEWerY7oiIi1h/4W/joGe
waJfXqaJL/jR0ZJ7dty3FCav3gA+b0lpWcV7FWuDW5ZSctNXCUl23lmZlMDs
eLqvVWolIn3f/FeglR0Z6As4egU7xtdVR6wvDquIoq5/uVWvLXFLE4031GGQ
mMX5MXkbT1s0fOlpCs5ev6zF4fTyEqCmzK5pfVwx4GtooAilASoMQgB/wwKQ
R8i9e+Zv1laC7G3ZMEmaVsyHJ3YzYUAu2JJae9E6UVbQW1Xu+EkCGSKvdVKZ
c0iIuLohY5FUgfXjItMLnLQGzL0vKNmyXrPc4mKeFgwPpa5eCx6w3JgG9pdc
L8Z+r71Vr7hLwhIzmeTwBAURIX1MWEZvNtIyFHCKVni8yBJMA4gWRuYx+/yn
JpNji7mNxcp/oGDn3EJAhVCPzpPUac0uRwbvW1XGWl1TFSKJrz/8wuE+jiJU
FqR3fbir6T/RELtngxl31YJd3z6hvLXtxK3M/Fmp1Uotlj/WRrbzoTHSMoyF
4sf02iL/ZMMsU/ZHBAjoIM95LFsCFrK3BrL/WRqqtXDZ2Z9ZW8a8UKiiPu6s
VfFEFslVumdsJXuR21vOtvMNKA/KaChAfNm/8Rw3n+ScWLoXRw942LvH/NAZ
dPCvxaXV9LDKej/yj7b6kBip0OGO36q2x/on8JSV7wJmSo9VTbhj01J8eg2f
K5mNS6wirVlSHFSYi2v8E4U5npKAoiazjEc/8fgKzCrwF+gfgz6Y/dpPxZF6
pVcVnSozsNzYQbkiGImuKWoo8OSQ0hjQQYJwtUb3HImLeXYAaiW1E3N3zVGs
LQycev9u9tPsGSsVJztTw1yLKJUCKi3oxn6sdyYENJu17D+3JRehfbzZp92o
XiBKIs9cgkfhS+b2Y0UFLvD/Yql5GYDxoxLiVdJQ3R6r/ZgeTpxO4kx4ragh
/k+Nswi8fr05VPNy00CauNch0XtKSg+Oz/VmR7RXsT1Y8FixJaXW9ANdJLck
JzSkUVkiyLqxN5/EqmsgxxQx19S64tzbriTHg+at8c+n7QKwaRGkh+OsxSIO
FwJDdpYCMftJVbsqHKmAl1lQA8s4vsOchqJaW10NolY5D3UvL0UvZaILEPla
AKpNIN1jJOZ75a5qF+76zx0G5An9xTWGeSQYpQE2rSHwyLqHyN/a0OXgy2VS
4NsMwtggfGKVRyUoW30Wo8vomw9tcW9x5aeY01W4He3gOKLeReCqlKJu7LlZ
2za7ZvIl4VBt51y4JRyIXgdaNgVOXe8RuxL4ogjau40GRRavmvcENFZRcM5O
XpMuWvma6nx0ushnddJMHo24DKDCD+e1YpWO1nELjMYlb7+/842eljLm2M+2
sXy31XWEEYcVYePT91gq63cUoXAIDXTguHQKrJ9UDklvsz+P/63DEHHfwzZ5
taeD+x5YvnULqNZR/EuW16WwAkxUPTZIzznzahHUpabt8W4mbBLrs3hfP44P
BBerufMbHLvRGG6snV/tvvIlAt5iUO5PieRp7+6LcRvEeXqkovsZrReT5j/y
RWQl7iPaSUeSBDQSd9CI5Sy67Mga7FW/sx8W9Bqvfw0crHKTbekZMPYEWoph
LLm7LrYSU9o4VEqLAZHArOwuidWg+wN4CNIS0pEKwPTYVsPd/SYobhcuwl3R
xWLecVPXbT9GJdylNS1UqQCMW1Sua4Jg71N4u/F64hNpBvfQtWamgrV6qWjF
wc8O7SnidKbsOih+fCi69+bzPngCcGRJfptUjhHENog3KB1jYavtrDZedlch
sZJMFbe/98y3smQ6YKUtHJlOjZl4LmjIW5fTj8uTMXuF0Fd7pYkwmveUICcd
/04n77kVQGq0ah1SYd3HA1UHRXm/0ap+0GytmlRFrooBWJmY15hfNh4kA1wU
sQjcEsIbxwkSJUg5a5QbIqpippNgvJ4GwTjEE/5+2HeC5H5LGw22jdemUOK6
ZhxPrNBaUjIqk/wYoAI436HlKJHP1IJ5lYbbd0QpvO9BCW8d4ii7DIDL4y/H
HOtj4u0TeDdd2VcjJMFT+pkdMLlPvdcp9OthNThCJhbNkEo0dYfqZMfK5YCW
zBr+4aiPjL+8wtVTHBeATxO6WRjUs42Lf0ix3Jj49P4EBt0U70uZfIoudizL
qiLbVv8Puj4PI794dtEE/zFt6BVz+mp/8084oosmDJHDW5lq1UrfxaIpAtu4
ihnfbu1gVQ3WOTxoZoi2zJR8ESkmjSZnUq2TC69bXT711GaJ815aPuQYgx2r
DahkmpzPuCOtWm9Q5p4iYC7Z/mAfvk2uX3VJuGhEAcg46/C0Db5en8fw5bS1
pdGSkc/HQZFieigNACZcfT33l+zFdC6g9BBTh/zzfo3I7OTCuGXhH08O5kcJ
FjkzkawncCaVvQJQyxXiEWGur6iZNxt5gN4bv+OukI7q3hg/YFgnwxVZ5DAE
o3iBz6uK2qD/WJAkFboCAatyxm8D6vJqMiJCoHvnxOZbuCuuysQWm0bDV9xd
+hfEM1cM2CzfQxtmaXX7eur4TTsn8IzqNXB3Be/iAX1C0qAvaTIiO/5VhspY
SVDP9XjR3PD6YKn6utoMJSEdhZ/gJzaiNXLV1Tz0dfb0T2aCWsaFuqIRibBX
1UUM8GO8nZlbYjXCr7Wekl2MuSKaYC1uT7d1wIu5IbfeMVQeDqwxlJJeCXeQ
ijP5TnvYvIP1A8QvW200HMv0CobQjrp3J+EMvWx59krDw/mhoRlFE6My04tI
LJ9Xvqm4X5Q35a0I+qRYOE8Q+sN7P82Bh9jyc/Gok4TPJMZcVYkvsLzAy1v2
6psPJJie1TrNP3DeZcMtu8wfBiMKTCFkRpxjo/zg3u4XscMhbNmi7OXtpqqZ
WYWvMhSa2377xTZEXzbds2ep8AS1jb7oeDW5N9uJ5QTTgXrHyUgp8fwgC3GP
gqzoexwrdZegria7dRPEETUqG7Zls+8lU6LrI6Ef2/e9KSerUnwE8yBGG3SP
8BmhKXXB0C3lQ1D+WtvMO30CiIdb9A5oFIFcXUP9iF+89yckyPdw3exLpHqW
Flj7A5yYCNcMeWzMHlN/nThAk9efHp+H3kpCTKcB2P6MPWtBr9WIB6sMWBIo
73aGiyYZlC2HZ4twzd2Q1B5IG8BAzYLBwLVgVd0aYAP+GKTdvqY50/csktnm
o47ahJmlJq++onqS9S1b503wykJhUWq0cZx0dAekRr9i2XpC3V/pIq4Awvmk
r9/7ZNLIFHZ2GOWUJVsJXxq8P15GPfJm/Jqs7ixHIXELLPUOourk437/2UMh
bAcnqDPhMq9rssVjWix65gxM/BZjpVdeszdShbQ4nwArqvX4M+HbHXaYNV/Z
yHaJoG3S9oWZliGUC/z4d2tkP+nMPSGjgWNm/5ZFlNRTT4mQB6v6DI5IE8Tw
G/oKa1QFqyqFi0NUG5SdLUbtsH65pp1wJbMn1khnlKd/gIzm6cehuplr0LWM
aM2Q/AeeNGs3xIux+UPp5o5Vn5JLw9qIbqWHyEmyBo+4UQ+kDGhdRsggYDPb
Z6X3TD9spTvNbCbGKW+YMXGlz/NtmHSY6ub6AjnM+OJHuThG7OrySmTTkIj+
xod+S+RZNrKNJlrlFNT09d5Ptf8pW076a3uuOcTGuMwHeVOZtSe9y2ClnyV/
FcLhT2lx2Vmye8EJjttLzNNbaVF/Pi338yDxaFjg7+LQqg0jnjmW66ILUAM1
1+/MeiDlA9O8xLsc8SMriuBthHXNMdU+MAhVQ9Y/9RpV/nXTwVWXFzV25NW0
eMGJ+xVeyWoQvCJTsfLtwUsCC0kGjLlOK4gvk5Ce6AQSXt/0BDxUe3cOX9/I
BVXaAmr/PfZCaJxL/MvLHzs/EvvYA8LSbrlVU00UwfeM28HQ3BAO69ttTcSb
QwdABEWm70KnXaSWdYk8aR+A+JdyfBDboqrHx1zmyVXWTOkaWZpv41tOUIOH
Ooscw9wsZ7VckdgRaAVRv04C9kGef7S8AuFA40K3WUpIugK3oBSJ7YOK24Sl
nFyWaCHF3SF9hsuwtYdBv0n9hzlqJ8VvE/P2zBXnK/0zjiqIUSxw9jDeboja
PfM8y1F34r6AQGnIqJTgIi7ocpJ2TT7f2Uzoa9JyF38TKSmrA/eBlXkHPA68
e9Z7aHsq3qwG3EediL0Ak8/zqYvMYuOq5OzHi29Bs8o33AZ3etZH/gkE/sFe
6RHSkfiu7QGoEGKdlCcLWdIV7ov72a5dOpR5aC5qkJJtwg9drzpYAE6sumS6
wHyel1wEfEd7EIwkdEJfVtP9dZ49rQCv/7Sxd9j4KQQ6CKSYCKM2LHrnCM7B
lVk+NyB5RzgH1EJo7uEpSR6C2uJsOU3yaQfK07XSEnpB080JTBydx56IZpjY
y4vD7+wH6mnOspQLK1DArQmAIbngNIYo9owcRxkWijdjcaqGm+uC83+WPzCL
jQui1mNX7BI2xvtKnH1J98PoD/r664F4D8+bO4Ynu3OKrz9FQ2TcMqEXlwA5
3LLRwL9umQVLBTJ2i6CEYIwVWM5bznCQAT63zLfAq4lqHVktVcAx7rPsDJ4P
dTFNHkRK/kybhiPWcD/2f0814Wrv/5K1kWDqnWbuVtUH8N2cgSDUaHCf843j
HjhbUq09LRRG7GPfmjRm1FPEMswFPlx4WGFzvkQrODMm0ivyLafmL+qJ8yVQ
uS2Y8SmCKMfOUG+ByHwec7mpB98O+h0Ga3OGmKSmk1PkTpJ6YRyuLkFOK0py
llKM9qOohaAm2WWWFJNFpN7KaOiinMzSpWhSauMJpiUo6HaZwR0/ME+0KX+X
lTY91CxS6b7ITcqeCAKCqV9YsI1wa8TDtzIagMxaOjWaDEKANQM6lCCHpunY
+Ge+gEfmXq5cNcSNHXkIZSAcJCUXQ9de/YqDb7OJsK2gT30jwhpg+dNlWW2w
H9YNxEiuzkruiQGijb9IK5o6xft2rceDXaj9YGpr4NZUbKZfEaig0H/8mBp0
XdXqtz1k67Kc8vvSN+LV8stXz8V7NluK8pmTHi4C09PQkW/O0AYLP/ncp3s6
ZzWn57OCnuDRyREKPpWFiH+ebARgAJi2+nkXrZj8+bzxENF9vnIQrUiC5KlI
+5XXBR3vCdqnUQkyaHVHMUtWwcR3GOE8jUsgzYfyrbzHLbLd0IavmuV4MA+n
VDHjGtQMnHZYIcbq8i/oiZdS7RmJHk0cGz3R0jQzgJSJkSr1Xk0+s91HmZJc
wpSAIFxFF7nMmuuldGH9NUo13Lherw0uCxcQlNO5QF2NSI9BSFXtXSvL4kGv
a+7rCdplHv93SRdcvrfnvxwhGn3cjlmOlYN5DwiLgUO1JY/ZS1cfc+tO5vmd
DTmMj1QjFpsxhkt1/f1bvrl/30WuhlgFAvs32OjMssaA5g7Pfw4QewQ4cOL9
bBwT4Do0FYbQ+OFaxsukC7JnKZRAmNT22uQri3CVOq6MS2fKNbPIDRBAUMRe
/1Gf98ApG6iTvnVwaVqTe0rajP5kvSoE/M/EY1mvTu4fkmzcBhKr1A3Jh5Li
u7qTxFj/UNqxsbABTaaf+zqk0KAv9zVu1ujN5Q7ynxE5P0BNOziakUgsF0Q0
FkVNN5F5zqfpN8tOM9e3Sz3gaUr8B6RtXuM4rrV36K/xPu0uiO2lwTMaWh9h
hfU0Iit98djfxDVBQJCwytfoW1rmAWHWaBVkoZTRcUWbLAXIwOw9tRm+wIGq
Lhi7xuC6xgneGmqFySr47fW/8OG7GNSUMMqANgjC+05ZME0V0GW5kqnEZcYc
GP+KCsBD/BaNjSqikdspNO7joz5P1bUN0GtObbKLU2+T2HCJyHPIW8tpGcLq
WP9H7t2M24dAwPdgn6JCZqJOW2/FZfNL9YETpoaOemmSofvAbVGTkAsHBtsc
UaTMJqzQ2RvvntEVQch3/Z35P3mhMQSCI6ezSFuSXlmOss9Ku9qqXFG/TSdP
ZP/p16aXHdE8lHnfTdJb6CHYTeQBRMv/nvJlhkx4gH50CQJGcNFmiK4R7MhK
ZnrQ6iJhYQxsmN9N5vL+JoYY7c6eoEmalxQjVkloGVfdHojU40wbBydrm1O/
I6998ZUllRRfK6Rx8WaNDHD1u7XbFA0dYI6YaD6z3pkxD9jBQ//jjiS3pyHl
40tnKCDIemWbYtZuaDDRP4ZInYLS5sU7FOcYLghhe0KKUicVqlUMda3m2wzA
0GhcfYQNH0JwfPJt8QJyAhaf9Q7n9yoG4p5HIxHn5BENDfD9U+rpHOCVJ9uQ
B0veU1NZ/pG9LYAdeaM1qBJ9CISaIfIlzzzLor33F6nUUzzisbYyuWSTEHbn
0h0RBmRyg5va3d4Dy0hfgYdKhhi953qKf8xKPFrRn9Yopgeamvp/wPJ27AlM
CojmHpZGkypGkTOoMPRCiI3jYqy/DwlnMoOafmk77av0PJz0ev9U5wdqtGG8
WSAo+aH0Oy7SvwwXPYS4EaWy7WmtyhmPTJR9snAZvjy5uzDEf8NqI9hMVX2F
pCY9esL2Bw2ilkgq7xFhEhAc1XGy9THgCWiHRKicCdtF1kFeR+5XWFdJRxh8
9Rx9I4mgkHq0EvG2yYUI0PWc0xpK5nKz89UJ/f+nUOlBCMRsJDWugQJ164tf
j1xFIZtSGALSXrQa5g9lnMwzN5fvlWj1u0vzTS5cYN94Kdzz7ltPHn9X3is2
MAjm7/8E+I7904t/KOlu576P2VrZmMgHynpr+rGMp9ASiMEStVXORjwQYUML
ASKbeIR1cvcH+H9nSNDdwEQudZjFclvg3xSM6TSzLaksFC3tR7W50x7UmioY
cHGvl+ROrMdwq980L5ZOaq6UXjBmSUMzpNZcyUuKQtiFdemnnwNE0i6iS6zr
ULWtlhEgHOyoOFbadj7B06h1sY/l17VBWML88VIrxNcZJzvF1Mq+ihvAL2gB
KPpU3IrfG2N4SCYigeP3f2rjkuIXEIwjN9BOkAtTCC++Jyvstg8DgvCjhKeG
ZqFKZjbjgws2/l+vDwnkS/XWUKUghSGy0Q+lILsQkK4L3thHSPpRcn+8m067
XY0VIm4iD3anVwJFpzrV1xlg3U1WD5jI1bRSrD4mPG7re2yRyUVt5eFJOZrZ
28MRxVTCfOXNCOVUogb2rfji8EFKmtA6qNRgovzVv/RqCVuVOfk0iqu/0Rh2
GJLtRQf7XxBFuy6Zi0C+Bal2379JDTzCxNGK8useqLFMR/7ZTTKZiYsv4QIs
BPub9VW9GHUrTmtmkiiOYexiHGzHOq9uP7hoSQrXvuw0fAjvG2njGXjpkhyw
W29UNrdyyzr/7K6ySKvT0sYmVAyB2G9AK3hnO3ooZWGu8azmd8pKDJteT+8d
zu4hcWPzN0e4JxL4p09V0pllo/hmQnABmv/lfaX78cxQpoFtVfzves52h/X4
eKCLpHQvMJ0B6S0MMawl7CAVduz8yWguYqFEcVyhqrWdN085IXGhnljtLcYK
lGqicozRIdOQqcuBRfziD78XZEwllun+eoMxMbbJU81wTrh/Cwk3nfsN6BRZ
PkBLZy9ePt0h5Ri4+VVTmi0lXJlgAUAtoUuqxV4Xk7A3WTDHVBtPa6m8SGZf
sG1GDWKgyoUQp63t+LffTAnJlO03/aeueH4nUfTYOR3wbA/K0oEkEVR+Zyg1
d1TeQMIvGUh/tyd8TmTOexT6Dwb/jNimuzsegDn9NZT6HYEFvCyjS+lqbTh1
rt2iUdCa3H71xUQ3bIb3KygyxxbMV2KjXKUq/rna2oB6kwyaktajBL0KRIgD
dqlp1iUYj1StZ3VubOkJRGpXBnFo/wgma9g66jIXvpzu5X+MUyRGtMFTqARp
c03qrrM7KkKVKU8G09y019LqIZd21AdI0nWQeOg4kCWKs+DIABy0BO5KGrFA
JpqG6nYvfq2JUiAPCaEr3oNr3ubGmYNe65sDzMlEHmU6YIsBDD2l5glmiZK/
sDPbVuZ17oruCnBsLZqnyPdH6KRj24MQ+56jkb+s1aumJKKSEztL0/3s+N8e
LQ8IzMFsw04g7GP87JeSgNsqQ5O3ryFmEaV6ss1+Kk5nZBdIwe0svr9YqFZX
ZdNVi8uB7mcoX4G3yQNjqiDJuZUOyoFDqS6STZ9l3wInJG7He/KCtXNBgrKu
eXsuOs/vMGInzpgEA6nYWa3n7j4K+pu78zFD6pvR4Rrv4MCJ21MUiLNRmOT5
FwI9pnXznDC/BjIakTI9vkOpuwQ+aMvVMDnt7dzQkr/jFdNmXZyJNb8bcmcT
0aP0pOQsPaM299A31lQrDNxyvyNnaCSBDS+lYVjcGHOFcM/79zezS5x5F6lF
FVOJRPe/XtclRBBIzIQX5RAFGNFdSiIVeh1MH7Akqu8f0DlyQ4Qa++FDT7wU
oRUsl5NYfBMMQ1cbrdkG9wCZxV90IarlKcELiYrDqecLZ3NNO+ryVJoZwrlO
VUawDllbIKVUWHZ8DyvGX4jw0lEN135jYey/VYy84g/g4Kxvk2glDe1jcxS6
kuEHkzRcymJj6TI9dbJSZsJM6WdVu5qO+8HLI/kPtKoAihxtyU9zFVMR4zzt
ldSJEMrdJjnO/FoSKaILvp86mK+Co+dDNxZXN4nsdU6JsXO1233rqd8PlW+M
66gqtDYU2jU8v3IrVwHTWbQK/CS83qvxYcW7TuA5zIIrvLLfWB3ygklCIBmF
0c0fqTmduk3XDIZ/w0+nE/KMozgcTlrnkw/AgboqNI9vMEKljPefJEom6PFG
73M/V59M5Uqt447D2RHIOvUqFEOS3p8BP4RzD97TWg+mT+YHC1YmpJ5fWHuv
wZnb/t01XmaVJi1gxmAt3UL58HCdv/8iZ7lonaYU8RXRj8t86LyX+aw+RW+g
A/WHL6IKjAMdh18bBfdPtUd9qsLBUpQwOHOvfc0C2UGANGNZRtUTkey2ipQg
i5UYegbuSl0NRcd2as7jOi0Fif8OW4BUwEwE/qmqDkY8etgpYvrOghziKRvi
YhGiHThOvZgQecCqIphQT0wW0znnhS5Xi8SRGm20VnEtNfxaCUbJQyp5qNUJ
3uFwa1+WOCLrTx+Rvwi+qF9mzGFeNi8Bqy7xEg8AotOfaSVrhAv1Va27iBla
Ds+CskALeB5cs0xsknZSeUduzgJevOV3yLkejzVUJtb+n+9hD7H6DVjQXx8n
ASvTYlEvCdBcBaP7txTYDmznAviZkQC70DPEdY2QCKJDiQUOX0uYG0oDNSW7
oMjDRjVMIxtelilbCqkmf7W8xPBwyv9ewO+vSGx2dtPRHn1xiPqDw28Q4lHg
n4iIQm+55u8/86/HZvpTBmwEto/ZIjehNZU18wuNttqsWEGvtEqm5oDYkSP0
JCNXvVc50e2bQDx684rYDGTrnQrkRmsSqofOiMdUf7MZNyolwvQ843FoLONL
ac5sxW1B6yU4MHmXbS1JL6fYxLYGe0l7i5eUCBNfnKNzwYsBdVDg9MfXKI1j
iDOtGmNH7rE10Yz4cDn4f46uUxWQNsfej4GZLqtyzuZlon+somqQit1149xS
H+8fzpnvpqoKYTEqoLVUwyeZH1Qzk4uNMGHDCVNvca2LBTd9bk//r0hJeNg9
AWYPXcDxybIwA97+k9rsjUwCFtbjaDKJThV3KR0oAqhhSJhgOqycWa7QX6kZ
db+Yic3nNHjmdyko7H6NvWF+1ZTbrQCTNRSla2/bpv+iTKB2+iwSkKaTdERi
pL/YSrO7MWd1bKpplI/wERT1wIK5NdoPzf/yIqWO5vI9N/Q4ikX7vWEoCTv8
9/GtcR7IcBPw9esocmLNjSIJYHsYqXwwnZ+YM2hfSj/rXOG1kDqFPCtMjdv+
4ki3rySUVgSapZjktdQvLpVWngsD1XNmZVrNx+yJdffQoeoFDBUbkZOtDCn0
j2nuB7QRIL7iUbhvvC9YGSD+kf8ocFCIfUpxh9ywykSBIO4Q4jDbOTWK2FCV
HWkOsSGzGxcqooV796ZYbUa4K5DDpjK3Ge85xjsXMxix80/fgNh5HuNNL2L0
2F3WykvnbTPNIC8EvV9SNPVnKTfeG0PMnpyJTsS+HnPN/PivlMxyR0DZc74x
Kuw5LAYO5NbuU/h0g84FWo4vO2by9vFuUK8LXjGXGtelVHJy11EYUZ86vtnx
nuW21YwB/HCW3TCPrsBXaDAFyYB5c0hlxF707zuzWDHDNb7hxQxMZ9fqI/1x
BlqYEstlpnWAGFicHW4g6o7gjzVF8SXN2lhfuKIiW06dadSgDRacgrHrcNKq
pzIvVyEWDwyr2rKy2UwT88xGT68aAaDZGj+CDo62/GvVlTjV2t/zXahlbm3o
z7OWevg+lU+mewYPR6PYQVnv2a1bwiSEQVRZerTmXGBFrpkKtwPeGgMPbxnC
6EtvquLluvdXYLdLc+I239rjajzD//UDrWtZzcBgVIcth6dSSlqodzyIoi65
7NOiHsTQEOdR60X93HQ8h3NqxwsJzvqhWPxvV6zDbIOtu65MM4vZtnu1bUNh
z2aL7mW7uIdejKMEz98410kUJtxIab+oqwwURL+PkPzPyfvX3LvTRiWPCQbQ
cJbltIm4IFDHu1SNJ1FFfiw0T/SsauiJpJ4buuHvABWivp78p0YA0QTfRdHa
EvmDI4Qd7vxu6Mxuxue8/LmkgKTh+8ho6c801shzzx4KyCjDIafiQ3zk6m+n
O/hvUji8Hsbml9AHehgZjHwSXvYR2310bahDo6l55PoCCJkasB/EgBW+aVLI
EztNAhJBIq4CII0Ya16AS2ZgGToVa5dQkTPfDqM96+ZBJCBlURtSMUIJpmGH
bxj/9vXpGop4pruDo7dFs3tJMAMw3sn9Wra5yMZjKAzfDOAnYx9Ua4zNH1h0
xkDh9ZQ+nwfOuHnfpNYk/MXz7XMNVFHP0HyhOSAz9gJ/1dTSjTxK1ulsq8c8
aaIm2+gzVfP/9Suww58IA0za5u/hMCdHTsFKM1qDLC3xrMigrMQ1OfcctsVu
PyWTbYdzLQWErsUSRC9D1mlewCM6gFiShSXpy/YUYKbzl0zu07frgs8G3s81
0tTVgnlv2UAFU0JOGxKiNzqRUHpHzpBcPSA7PgtnvZKMkdbneQoo34CTImEZ
LIiOMp2qpx8Ypb6LxwLtE3L6cfDlx3dakaumlI8G4PqJKHLQHqH0RRibDlBc
FlTM67VzwOgpdnkOUEA3qY6zYvOzb+EZUjRT9ZH79AWwTNhGq55zPvvadlVz
e9TZY2fEk+EtK+lRT6xrqCSVAawl8FqbmhQkH1fSHKvQ0es+AGDSznQc0aed
dRM2mL5+FOPDaljDn/qKwfyITryrv6zWksOKuV6IDOb/+JXJwldJuQeZgdXw
5fMy74AmpWGNavGAtj1U3TyvKTiy+lhnLGJFW/W6DFy+OuCCqyPdunRIGv7S
NOmvaUocCilbz5pRYcXsX6yl+iC1JKjJvszkrqvQB/s1HLed0V0QaHIe8QqV
0alAvQJX2qgPftzg5r496G7IIYgg1qzy6OuDp4kOhmw/QCRDE9YyvBoxQzf9
sF86xNAU7pNcLJl9NwwIge9M/ziJP+dSEZZOQKpqJ5FmqBh+ILFYRt2pSRfK
R0kRbadW5TOEka9uvGJlRq1yX/mR0w7NSUzkK4V5aU267TX9iqcOHCbp5In5
a1nsLeI9BHco9FduqhY8YYhFNOgRuKAM0/xM2TAtvZtDEqHp2Ye8AGjhCUYw
N/XnkqxbTcbIrVFVdNpRVY7/D3HDT/lhjvaNMyTXfcTPgnPtIk2pZVsrTw81
qNxt/TPl1AXArjfd0rv8x4PZxdNisLNt4ILVSRWS6ifV4TjP9LjUn2kPpYuW
FQh6N8RuW9DehJUZ5iL9tkE2lplD8JAvPdTjPFLiFtDZul/KX7bPORYMh+Ty
5vhYgvVs4rEs9OYbFxsxjZE4LmRrZmAzVNbRKKWSpdaR3Ll5tz2q8Qe2kozf
W0WBYKsL7kiX9n/eahbgzFCFtaa3WGxLyC805MwB4VnMwMzlZTDwHblhGB5e
Z8zM/NXa5Smd3tFRu0VvrNgEpuAj4HeAzzwmxqcs0ohFl+LPI5s9DqECpJNL
jM0D2ZTG7t8mgQvTJ8xoRQHBQB3SK79/u5xVMnYhSsaZ32FutJywv8lQtpIC
fhN4h4eYMBAzHCU2P+NYS1kjFWJtolq9pm2OcAy2wuJDv9UG/isfIZPi8l/S
GE3BJxf6N7Gmu3WT+NTAHn5MMiA2eQtFnYXCZy/aXLV4X6WLo7UUzUepuR95
4uKuEJC5Iv2WVlG8NRIn0GEQRjLy3jleLeRAbWB+1pHPuRkbDm9XbxbVHQPe
B1mgw4pLnx9I/SN674MIc9PS9oA5o/z2OuTjN/fE/vxCxeZLN7+YDhvgJDdN
BOvaYerTvBTGuGGR6To7r1XGQod4d4HDw+dCAG3C2dv2WRtbeFLB8qX+sYqH
wIeTKH0Dxkp2xshWiXq6TYU7f7EU6/qBOBnAUFxA4FqYFsXTzXhR9KLcRhkU
ul87lS0uDOozE9qMNNnIm1ZDcvtyjBuJHfkYYBTeL3h/JsiQjAo4WK/9KPKx
Q9C0aGtIuuhooBtdD5d/X+V3I70PfTABH+vQGfzvsoUp+b5hva/9XT3WPm6c
MU+Sva2fEVOAbqzvR4B6SQqwMzXV0JFACgi5OKVKd7kCqXptV3ntHPfBzMz6
U/5MfJ+edTCcv5CdbXwD8rGefSLzJEYw9vHvD0m90BwVovVnXoFC5YMI4ZpH
kFM6zR7+Vwqio4xrL58qEDVOVMJNbuH9DSPGHEFFICkEMCbmCYCGKKcv4low
rv7ZsGSHTeDx9Ep/kZRgZynZo6UuCLcEU3FTZ75FGxqGE4wa2gT1YpYiOm1U
MNUeileniMAr9E619A/38MbBeHfciorqUrJ9Ix1Zl1HdLup9zuhUz7oTAEOE
3wrcvutTx5oQhDPZzuixvogILiHLTOvhRxk5Y6IhKLDqGWd8LdVbmArh5Xhc
XOS+yVZPPfOPd1zzhcWIt87f7a/mGOjsExL4fKAAHCzqm/tJ8bc5izSUY9fs
VXZzzPGtsUSn15ohO5ovUFtkkCd75ZRbXru+QVzfJOMdTktRQppXN4Qg7hsB
R9ABmrfprlr3B7/9Vm5NfSalzNjsy62Tt+e/gCvNrVnlDvmA1cuJka2R3fFV
/hth55gWuGORz/DAi3SZVnl5IskimfKCKOgH4gPg/jU4AvIphd8eymyPem8q
/FyDfu4Pbu47j7qJUpxle5DUCXylZtRhoJvGc/dAGgRP8d5UdcqQvgeyjrN3
+qFsj/5tV2KsRxyXHf+nbBPf7iIpZRTirNxqw+ER33qYMHkP73DbdRgpjfLx
v10imweZ4m4+qUDxPBaJfz9OQquYfcGO8xon8sgCpwEd5SP4bPfAN0Es8qye
nNfvx7MWol3iiRkY1KpRURgljSUYnao2uxn4/V78kQ48X88MYG/0Gh9qt3hA
N8OSJPBhnm3PiD8pQgbPX1x3n9eSpul2RN7X+S84ePB2/5igMfiXO2xeqDlF
k5xd639BxtuDkoNlaTYM7HZlWYa6fz4fSrPFBz46JeJwazHsEaTcx8ZeAPyQ
dWt2EH/bNj5tX8FaVtC0dG+NZNE82WdCafmIa9wzLNFXtSmWvA5zEDUiPheG
z799VK6leZK9BOqOlnWhxvWw4gI9ShAR2DMhobA5zBkRvsl/7+ATySsoEzR4
uTNkxyR4ijHKeDMUIHxTqypHoTo8FD+M82yKVk+ZuTrbcO7BZ7jEADNje1Jl
rDJqATOimbSibefmQNEiGy6e18qU7d4PCjyLMcOkezq7YlqPb678X189rfYE
YjD2wnx6bQlecdTExPThLt4NyCSla0dGm6vmIdXYzslms/33zjn7Esz+Wrep
20fUsKu9Bqew+kTnygGpec2+LVx50IEcTuDsKaX6cnsBBgiHMaN4Zg/tnXQk
gfss7/eEcEUNeQ6YedlFgC69zT3P3WVI94TdX2+sw8YDHWTMuOt12Oo45G8t
6DTIo0Xxd4HKVODkb74Sf3aiBRtszE5ieRlLY56ElNM17PXEpoohxzCxBlSy
Hp0Zo3X3lIMJoLVDez423ECtQVn3gp/4IAnv6nmm/DLaYF4dlHz9Kj1cnqJw
Lia7wYxgNF265jGvS1r6x+eJnFPokjV1T+vMm5gx8ib4fhPHmSFKQXzrPb81
jUhwmrdul8vchero3USdbmDpD6rYEK0zmByfkfGB89Gh9ZV1mU5ZuLN2ycqq
MbxqjTkL3zAv+CuQeKSp72uPfjivP9c134By/LetHpcVqYkUildRYZtsPm3C
jfKtQ2NEPRbsk/EF5hOW+dx/RrARg0AgjCKXlS2/YOoBeMzNpu8ztsUdYXPx
GT5tCzNxmjv+C6lH0mRz1Ts4VUVM3XSCRYiJS0g7akSLvAJEQfTyBSI/14To
rgsmLfteWlSuQfvGEAc8Pue1tNm32enZRk9dMu2g+yY+TNxcVKz2TVsjTIIn
8ECx4fqNQFGnjUPOnxjkUDTnZTg4eEPNDruJxnXusUYC2VduKYjrnL2DetgR
CLs1fX4sxNkh7U1900JZ3eCSSIMCruAjs8ZihBXx0lF0OOQ7NJ/Ecc1j30uv
s3h8d5a4zHijzH3sSoDYuhRU3lJiNg+ANpxRXVEHbAvgbt6JHmtxVz0HQt3t
mCJjijChERsjNX0iFInp1e4F8wmy0uaam9+//mlLCfOXCnk5EBaTkJwwbt/j
lp5siLpGNzzfb0T2vJ9fhW3tRGoNgkIaF/LPoZb81mqbfxMtA79WwxeHkGZ/
I1krvspwSPjTRHLEKqvovHCLy03zUWy2xQVg7QDtJBBeYDvne6+RCtUG2ID2
jWEZUFufuYvoc4zGxX67B4kF5jbwCktdH/oMH0VFRqXGIrNwMYak9Q/K+Bm5
DpU/F8Rp40QAbkQBEhlOiIWq4jtMdEuGggRSB4D41Gky46BPcpTZBivzsTfM
V+r0uCEe3ZtVCnFAiZIBPcZ/eOhr4epiCwojtuPrTvY4WbyeOhyllD1pFdDl
sQ4YCBIZzYFIzlV8rHvMAcvKpYuhH640w2eYqyuHghgb3BerWY71GflQTPm2
ug4PUwiCERnp9eusuffC6x+YoArVjxfg54Mue08MyUUuLJp+6Uhe/kdO/y7r
FlsT+mRIgmgIUZ5FXqzOjAxGklpC0I6rl4BuuHQ0BfstQ1QbZsj8Fr3I7c0M
qLXDQrioVnPbacf06txu4CF3TQUTpzaa8qV5LzpoKd9zX8mz1eQEzWPoRwTc
4hCHqDkEHAsdRFHufMFffRT+ZUUGlyKW4oQ5wH8UpY29pkssMpBi6RdlxWLa
HbXyssysk+C7eaTGIVAbyweFkUs26hQfUCDH9XLSqrhlcyULDtKfdei8vY8X
fwFNbB5zNPLSPe7AUj1zxCRSc00ZlKjG9G5kGs6jWXBr3x+NTOPtRjjHyhjf
lisEeSGuZ132KNkeNHGdj6juYybB6KgtoF6C1wN8yv7hTMaJ0AeFqiTBS9Vy
o9UXMUf744VKyc8eUnHmSRNnSld2p3Sb2kVqO/sUONT3wneofyScjaYnkjCt
bqHHXEwUKQvB0Ghp+P7xVR8mFOG587IENBjIRMVRo4YMflFh3FywM1kH6x8z
9MspF33IGDOZXHsFbsh7MEAGu9AQJeVKWq93YshzFx84GZaROwHrfr4yPvqx
0J4oTDrcEqUcQfYPHFMO2sb5YF47ErRuagRk4rIEMlO2Tp0RJP5YzZC/fyUx
DTdMG5cRqMRCtaAq87t80K03/dY6CbDGEh2ZHG19PrBHvVHK/qv6oQt7I0nd
hq/+7FPvo1O2kuf2Sn0ZGXke1FrLZnECWPYP0NfNfTXpiAtwCUw0tTeQjtKl
vAkwbt2YIwq50vazCTh2KUHJeUovu1XmhpCaluMs6suLfJDn8HW4MvLaf3+E
MY4pD6WGV5ZrKZV+eTmhnMnNg052AeKW5hBZLZyFW7OrOteqWquvsabCNM7X
oF4vPi+R9NlOmS7xgPQ+MakrM0GKq0PeaJ5aM1hTJvaazoYgtb+ZK+bIL74s
cRfKO0/OnEp6PxHlxY3m5496s77WyQCKg751ln5KZW6tuCNlYayOXiz/8fId
HcqjGRdx+Q6bs5tGS8D4DEBsXQ9aJI3BDxBKXx+HJzRGmmUY8BpPehBv3EgR
yHf3baMtF4+H9N5Y3VN4XGkOtRgGIbzCNHEPOQxkSkow+ATqQaSuuooPOb7D
NYAT4j2xb/CEWA7ZH4KH4nL6Jpkib8jynAi6YxrQGoNYleJWKF60VJOWiNAa
PDwk8eZF9Ai269p8j9ytzis2dcBHk3QMTf5JHPLpkTsjcs2e5tGA6/y4baP8
XmzYVfFZL+50ovIOoSm8XUCP3b+KH+kp8ZtWRIe3tyUIYLEdYCdDYsP9VVxp
Evq0b3qZOINpGaB6xxnspo6L4nW3FLsEVmVpO1gt88rXKOF6rzhyiULLn5Q7
nvfrrTiJlRg1zmNykO35L99LkOUKtlm+NaS1YC6hFna8ghtYQEZ38TDErKQx
IUilxL64fT3EKPLe5nR8lGU1ZpaNFBREwILt29qdvT4PXcdN2dHuNfQ0/QJu
d12lls19rk7tEZSevIR3lI9QYKTWL9rFnKjqrNIOU6ZoD154bAX9iWcrYaYz
3Pwbls0N0CDblY+NQ/o+Zp2hne4jC5M42J97YuQoWitHVM80xAspDw38P/7i
EEgUpn9a7uf9o+51cs4FVCnsY7De7oJXv1w0FT7f5a8UJSjtC/qc4VmMx5oO
KU2Pa4+2imWQr2q2pGPWFEf/lC0XTibZ0ttn/Kan0rqUKw2WdNjphADrq8C6
vlbLZizS48ofVUdWWR2P0BvTy7PHgFvPM8IA9Zrt6RvU6EwUInVrMGP4u/H3
7gwuYsDcNGa5Kcn6zz/gI/gYN/MHDvVTn8Kgs45zzOVBxbEpLTJ9J/zV2cWC
DkB9N1iTjtUaKjwtt36Y+VeWX0+aVBf+DlcY1i/hWZsysJB/hnvzdDIv1C+x
i8Ff/wqkUzSxsBQH7e2LP4ZH2TLf3cWcJMLxLlrMr9Eth/dCMy3Us8ZLNW1h
KqeoMWti7SEVUu7hXhpS+2Kr/iKWYu5QX0n6Y9EIGRDHW7t9pJfFKp04qZ7r
gpI4eRCQJl2KB8uUY0fJ7MeYGjjktnHbvPZu4I7eV4OUs39wCTO5G9Xk2GE2
+dy1N3HoBPBlcK9qz9/ov1/Nz67UUDqk4as1dFUFjpGWWU8D1+y92Y7FV/Ne
ew5lc6kZUOmM/VHv2teivan0FTLGzbRCWxI8d/mNH+1LyNEdnxNC1f5SnkM3
EbauoKwyozE9sWUTplAp2EML333LLssd5AyG3lffmfHKsqMCLiOzLQG0iFEi
x0T/0cs2vkJysUmKlXuATkNtjKKtzSV/a8ggJe2LydCz40ID35jHbvvdYpbl
zoAtaMTXc+oaK8sUIrVHYg8aaKg7WN/sfNe2ipxWsY0+UDVI4LI/Goh6yndy
TJxZ2O2xi3amh9rjEZHknhx40tR12gCA4ZAyNLFHB+zxfAelSLpToMIf8v5U
npkjZ6/48rzloHigUMPUawHSBF8QWzMhd5IN85T3hgJs/eMOX9igZa0K0eUC
MIjKhVQJtDZT8nn82nF1jCHfWpONYjb+6RwIb3qCmviSS6+yk0hMEe12lo1E
FNOwFRn0yVj3iv6XF056MLw2ZohKUDBG1FHatCFLuu06Njvw+9bSu0TAY2kn
xSEuAUOlwsyI5QFTB4ep/BUpUQhZXoerYoODWq2r6/od2g3OyZptj3nHTQJM
SKUXDXnyox3EvEDRSRzmhr0COnQcCpjqb+lVJ4pRlLWj30fM9K2jATh1YadT
BiBAm035uijgcaLY+ojKviIziQuGjdZQDXPairH5jQ/R2ny2eFfEWZLAAX3O
fh50vcFJDBnQjfDXkQeRmzxm9Sy6xRSTQlUW6of41UBXSX40zMWiVE65YK0R
78gsEcHoiT2sxiGxY2/a8aS0h0aP+IuqGkd12pdh6lthxXzdlvt3qucWNeL9
DujPK6fEqmMjLvpq6wonbpO0y87WhAXgGAR0nZUjqv3qcxe/71OeYtIEkTCf
RFi3b4TJdwXtKh00Fg87Av1DUgWSgd1DJo3Dgmf9p+OOX563JGH+iB1mHN2F
aLBg4QVdeErxWCtWABYk4ANC5gheK4PDwD4fe0G/lhbe5GMTskLStHz++xZe
89R+NWU5rf6MPoJSbjrmjN7YUXIpPyBabGvVoXG49SyZr+0Y2IJR2B62x4el
DzSd0+BieEvl/1FkvLc3x5DbN5yWOH3p4Mrze4k1QOW6bzqBQ71TTFY0X3CH
iYoqOgjK5IUDNGKWaQa/07sC0sDVgoCf62ffkQhnE4S/mhYLjcxGKmjoT0g7
1KlE6p20LaukHNAdQH6aC7dPvX6vauhN+AmbLGdgQIPJkBggnzIw2QD/MK5D
CP0/RdQW0Am9R6ef8Cj2Rxibv9zC8x7FIehQaHuchSFfdbY/TvRZUOtUtZlB
tv2MiN+EcDUe2CatYThVItitJWyb+6mBY/qkcCLvq2U3poBfsbInpudGUtXt
lBVDSVek94t+fQdZbZMhJE4aUOXQd3Pj8MWOgsQrdhPs138jvpk60q95pqPD
gyIeQ5Dp8YWDLv7H1deeYV8QGmssoEVVCf2wm3A5siM869ckOzXhkL/URIqs
6DQg3ATfMMpPIOmeRjj9ioDyctP1hJ+B4mLiL1mDAp7wKsmGotr8DGZdPGry
2doX1cfmbPbfOpiZNjwkrLqBlB+MSbi0klfcCT0jB7uttB7Cot4ZvW5G3CC7
dcyP5R4n8fh4gHK49u+0blQjKqb5rQrYH+S5eAYfVPDJMX3q+wA3ESO8c0Pt
Amgq639bxFNx/SyhM0O6x36Rz4QSqAd6zN6aH16kNuGeYfz+p3TWkiz/am5M
MrZqxuY+0vIkotFxXN2QrjYpZwdQswgNoTxD+vaSRd7Hl+K5X4NvSLjaVDjM
PWaovRm+DXOSMKSVpJouTGpeIVqp7zBoQh3PGVfxRO054gs77X+wvm3aIo26
X+odrtPhlqWwmGLM7R2JRWWvj7q64kGeo15EkCRjndp5ungHeYCC0sAN9YDm
jwXmjzrJyNhrgZxR7QXO1bZ1I4Upvi+6OH11+QY5ur02h52fDsoETyySbCY6
OL2T29+1+XnHdYU1wjT82HTG61B7qifpEENGRmKURCoSxelCcaZg9piAkT7t
US5jBiWT/oMqwJwMs/mv5nnt8wTeKmkgwsvriXwU7Ji0I+tZj7NL/jcRGJuo
FxBV8NOIuyWz1YfyXy6CDhUq0rqTs7C67VW4ym5Bf1h4jyfeQSQQgeP8y/oo
tIkSWxuVSYeOuFUm8toJ/hXCz+KXicMLv90RADDEkapWGEVHJB84uGFBaibX
iT9dMZv1kzZuhCJZmTZcfG569XCKLDEYEAtK7zlze9Jon7E5cCrl5Rqc8YsO
pwL4vYsvrdXY5qnUlx8XiPUXThEiYTuex57uUVlO92IXgi3X+sx0AVUl2J3u
1JJCjuuBQWjFAI8A/rCnjeCIjRUIvIcTRO34uFx5SoO4a4FPZ7l5f5uHqwn7
y2u6sbwbBKWS1yQycyHSGzWshn0NM/ohn+BHXcqM1ZycI1Y+sD7DeoJQ4KfD
tjohp4QgYJFe5ZcYkG6KNOcvymW4xi+OPSoZdBpHRU0iZryAlDkxlsccs7LA
0/ESBESYRleb4dodXXTm2VEhGlmtOl4CZL/nIOt319h6pPTFX4wRXweaJELf
b3cgNKEi55/qmFR4i4bMvdtPFJYERLap24TckrtWUsBxUZ5B2me5t0rm8gih
pgsBdckV2cJNsZtPxj0ONHJ6Kx9lJFJHOq7aI0BqN1UcIxhXUgmh2JDBkQSe
ilYq+LK84G+yFJkNQbzceUazuflb9mAs2qe49qy+lT06zJ6NJ1tYBVSLMxBg
yPMVaDtMQmla2wvwlBv+wxEmQ+hfoxTULvTG0W90huUrCHuG7UZnchqprijK
M4gvxGfKMGtU729KU/ldSrTSftP2jMGxEsWaDcxYDx4YofqiHT0NVosbWDDK
OH4NROkLqAKa4pvURI/PbyCkpErvt4Lj50OLWkRtlAW1Vsook48UFuDGYn9J
+QkgH3KVOVY7YYhALTv2lFQYhZm6G5aS2GQbuAhoAB7zUA9YMl5kodmYMKty
v2z8ujJ25fDdCymXZSu9bEsuxD9fa2opMDv1uyarrmtw2hO77SlGK3xViPJN
V21PckkHd9dr19Yb+V78pHmRENSRh5LEHjrdTHNKmHRP5FQTPs5wSh/UlhHP
EXRwIjbkeCMWC1TIshR6IKrGDEO5sSAggTF2BpHnw6tJSMmpb9TgRwrxkEH7
HcQ9KnQWEm9B+zMkCrYJ9Ip9fEy2o1xc3vWZ2wH7OCtQpxXMSntA4e6fJR5E
OmZuwXTug6pLCFUYLwMmQ0zJ130WiLD8LOsTXdpBLxmAO2ABuoissRSmtkCm
wpKM+f/wnISlQPKIqcPDewQs2YEa1V6tg9r5i+J7c45+86o4G6dizO9XG5Y6
1Te5q88JrY4SlCuKaLrf8Q3e2GmF3Gh5tUQCWBXJB+JtRnbRANeHZQWh/bBK
dWo7xtJHwZDoT8vioSQtSsfIdLpMcFHnUZqWZwd8nm7KYJPy2FvPEScfqtx+
gzlRAGDbfLlzo2g9+7ou71U3llEOY++d2cgO9TLyYhX4i5sAQ91tXdf5D90q
6IGY5EG7z1vtef7WkCn5Td3CPJxNint/LUy3heMNhf/UD64VN6LgjWRmir8r
J7vy/cvxe35hrL4QjV0raWgoUUFzlh5nBGO5FkBIUAr36BWSV+saFPd5WCLe
i9CDtupUms40r42mz77LiZuTKEoyRqoPzwIwb7o8fVxA92naS5gBSRgO1Pmm
jzhHyT871qLdyLSkxVn9gyHSynCL1N4QCt7qg9iZeLT6As06O6TUP99/G5NU
HnZ0+mZ9rakiL6iFpihNO2Hf8105YH/MHwC7N3vvtM1z0fSqwClgJNmh/Jx8
IxoH+QrPFsJi2SDDyKasYnS1DsT2DOVeK4qxKiXiaFZGMIxokxGg0vQ0U50T
guyotBYC2E2jez4taTebVlMB0d/Mm0RxBVsEW0a616mRNyYw0eegwXq1Wsla
WwoWqMsHb2+Bdtv+SnsmJLzMqIklaZduECqR8D/u5gxRPQuwdwj4D/GtAhV6
+KKdtk9/Cd7+cRJmO8bh7YnoQTXt+CsuhGCLP2mroNaEuG7i79d/VIgOmyKY
7CqxMPXGw0Juz8nnmlc2k2IaNimR6iv0X2mPPA8p4xYvQ0bf+DUffIoI+MGP
WEXHZkgYLwanOQRivGz5QJy1ijLMkpJvfGZMNL7d1mB6NGIEoJcuygkejpAr
4S4ZA0R7q2LRIi8a1gxbGxsIzm1rAEtupAuHvxaTe3kNcdeOA1gGPBBr11To
3TeYqp+neFfe78GaRGHjXMqLBHc3ElnJysTgugEIo++Mef3CEonpjjZy63sV
PTQIHMoBH04xqfhyygqqXD2pFYoyPVVfxQaQFcQbqqcztLY13quFNkwjFvNh
B36o+4yuiG8X1LlF88xucP78YJN286G28HWg0fDG/etsW2SdtiV9uLil6sBF
rVE4ZKBC1lLk73zg2q5q8G4PTWrUNgYTfQrg3fcs9ZZyqvuYmwLja3SZmE0A
mO1TiwRT0lKuxvdrP1ZqPkVc8t17l7WJNqlcY+Ks1vrzQIFAmLDrFb0flKxN
DPT4zBOFC+LVBTv2WLHhzh4uyMCCDLdqM6k/STASsj8dghZoIxuoG3d5GbcX
32rs0+rxWb1mdVipFbS5AAkq+WgHhUSDT2dCU636SQcJv4L3AxZHl1zUUYBL
IvSjX0FMltv3VAyMoOs6J/8Dfc9qmIxPgVmDWMuf8sb5oqMuWuh6tU7T6KQg
ot0gRVCniE4GfbHVG36TqNRZ00StAtoLBKxVeIhyTQ7meNMCs2NimsWMbKWh
KAdFbQGZanFsKBsnhce6q/bNJWu82P1yRHiTQv0qtobUs1jmxVMCfKqSx6WL
T1wIg8vexnAWH90v0hSNTAFCld4z1ukZQLK3Zns2bEexqUtvLKJZynl1myOJ
mBggQ4gy+x4ClKI0q3hjtWwwF4eJEzEPwAFDRaSxOXFEX5jj9cExN5lWnGhP
i/cFT5vJG7udCZmpgrJ2j4LqVYJpzA0I0ZuPUtx8PszRrDYU+PZBlQdl8kxQ
NI1gB5ctYwFzL/QsmhPj8jCwZen7S3RVyFicstk/kCVciFL2Q+iTPQL+tIqy
8fYCi/nnGpQaq4ILCRd3kTiG+tOx+F7JO7oy3Wxrg5PdafYiVBK2MCodSCS7
QzOqMmNe4AKWCYkunM6gonVdDxy4FhWNtLbmQ6lzcAvflYLBuY23Uoz6pbia
dcKWvgHIDMIDlNl3+d6aqG6egSHkR1DB5prvIk07BfqDxtTz8PXUL5jFGjic
s41sAnusCDPgDDTlWxDqCGIE1qQYJCK1kx7TfMlIKAACtqs1LdRV29WD1l8y
JKUWpzvCXxgPzExC3Dj8a0V8AW8l2greXWVM5SZtM1jTNvOf6Ugq7Dg7895p
oDv4+LukyfzhaU7OxxkCSgGFA2vBqt8TraVcaQQKCoFPQGk4R9VPSZm2sx7J
0RRK1lYonNQKYt3yEOS8Mq/Bs64IQC4MrgSESofmmEeUwApYdMOOX1BqXUbO
fR6d33Jl/9BsfqI6eWTXMDj2Ea5a2CW2Y2MSQlisUfBXjolLKSBM7+3vBdDa
MV9e9JEfvszOQ7uZCnl52IAKQiBSnPPNL2ZzKLayA9PesUn9B3itK+v5nQVk
n90Rt1bHRJ6/KqmeEUpZmg7CVNpvQixSnmYrV06I6m53zzsH3n2uQRIzUSoA
RKGr+CnAfIMdEjp925x4nzeEupMOKHiC5Jjle+lQdfbuX3Vk1SE4MHJEVLHp
bw2rEx/GiZA4V+DxtnSlu4NoUpbq7SNoTtOMM5pM6PYUp+YU8vI7Dxf3crXl
SnNCz7cibMdLRiHiUXLDIeQ3cas2CEJJRSWQc2nmJT963j3R0z2Pc+4bQZeY
JeVaLF6fYlb4atsNbafajqWn0CDqRi253A+EUSWrOshM7cQqWxv8eylIN5kA
iLIYxUs7Mxhut1Rt1JCihGkKTJzf4dPTlwuAwTem2clDixsyyr+wDwInb16t
8o/kw9gjSgkUJ2qFe96E9ven5O7WGJiMDccr6dJLH3V6DCkgMmIGgN8UgbBC
hwi0ACfdEu8vXO0s9gOZskngByNAV8YHuqLjIZ51xEXrP0fC8kUWvzEE/Krm
lR2hzCMZH+C1HDDcLmao0DfaSuaSyOtRFmTRcTsbmZCMWCVW/Y+2cyov0vG9
/vK8raccIXykFC2cHQ/cdEGi+5wwqLrg0DJ9CNlvf7V0lLMhlhDkkhkhlw48
RsqwbMxU1SHH5QkrVVeBnyRHszvf1FO7mBdFTm0Qau788dM3nsxgc5CgvVdx
qU8EhtNDCLyqwUNeTXefGgSnT5FFpjUxoblHCY5+AvIkk7VBVUXTEuo1UR82
1ADM8622SnA5sF/08vyYXtPWcn++R57g584IBklmfGDOHTO3BaHCSfBTQa8U
lea3ejRs5HVbPoBWejOX42r0Lpi2uzVSvE24uTZ9+NA8rj5j7Ti03oHyMnVf
+5o+uyVxx+U5Hm4vcHm6pnq1Q2QCQCRPc2HUGbbIR1zP+VTE4ff5727TgtSB
MbkdWYbzhvxXlHszepwXsZ/O4628L/g0dynIz940+rHZLkTlTxONPjHR1xx8
zvaOfbANIghubhg+UYwVmHKfzDtScvGUXdUmKQjEWU3yUumUc98FuNIjmboW
iS0vShveYwMiLgNkYcDtzS7lft7S48LH3hFwt4RWGGSmbWyWhnDQv6EaZDsm
eVNEIXVv1wapDUhwoV49WTJOW9JQt3H0O1U6pxlnB7MPtX7CCUN8BWwUNkl0
8yOiTupc03DEPnwbr8ekUUzlNWBxitZwQ84STAhW3dac6XCDVM4/Kduz077J
ydW2oD2sVp0xC1PX/b69RMHPkjmChSl4MX8Xq95m+C8YpYgeUn77kYas9LU4
DdpGVT555a6AcKsaRbobw2zjWr3SD3uu3/RIZIKyeLMBEtWT4EBvjwxE8no7
+5/HR6lk/QOwvMigs2gd1ybNpXPAHLzU37vvTrVQQpj1ffHIC/nQbBOZT4Gr
/ibBlexb68GjnHqFLWpr7ofMO93fpGZgR8pmws5c0MevIeojyTLWspWOVC9K
Hw50aevRsAZJNjpz6GzK5qInRterGMit+P2iH+ULaCMUvC1g9QsFPsjaf6c0
sBsJzlhp4crJcojr5jJ7aIL/qNnaBpcxznSuhZ5vqMhArK3F1zA3qR5JBf3J
4Rnd2Wbl3vJIz0uzJlfMptFt5hCZIAGVfmW/l162dQocusAGBk0UmBTBsQ5G
gWzHOhwrLfZpAnr+fwfoqTBX/e7WqiTb89gBZuvCHt42N/S5gquC0gm8hpdE
nEHcr0fCUhajdW/serM8ik/t7FC1tUxxbNSdTXqBe/z9de+JcehFuSYfH/Zc
g6/7SiPdDYINQxtKNXg6uFhh+EoxtMf70odH0MFBo5kmp7Qg88HQlZ1Nzpa+
9RUHrki+ZBKp23S/y2b9Go9nWLWDf39FB9S3bKF5jd+L20TQAfvtqdxAFV7B
2YFxohVT7hSjy3OyxyzqH+DHhIbHs9q6xIu6qhgMivsrp3rWsuZ3lRzt5ff7
Oj7JpbDBFnPBn2hh6isjDdK+iSHNoDhb/HsrJPDWjMjzahFEKelHxuH/sEYQ
d30+G+O3cYfTJDAGzZP/Um+IsHekgvkHuCq6ZM1xwhLmyRg175wmIvHxt+Zm
UGHjTU1PwzqmVpn1Zc8fSOD7elIwKYPKpijQZ7Zas3++HFqPTstVtDfmwyWI
Xst/zzfYXBMppoj9sGqlqaLiJJxGBGqyW+S0baGQOTV8fE5kyBs6kMkb48GY
O4mSBZyXerpQdAbrhCjSpRFcdcjNT6a6NblXG1SqmHJMjMolykyOhBwLwKwz
cBWchHbr5LKfUNq10jIU8fBXOhk5aKEU6iJyfSERTgALVzG2Fl9vwM6iVZFx
XjNJouAoIw7TCsysgqGBj4krANCNcyXPh7QJlLl+ZiiLji1d4uNEAgXv2vFg
ww9xQ5uJj7MH5MSDnC/Hi8jwKpr2RzcOYkTQMNEmhr/PA6JfEbg5vyX+nE3m
dAZqrUV9b0h4fG59GEP3v84/rxxpzBq97D5DuV7E4h8ulysiEjDau2M2FFpG
ect6bSYbin6EAgU5192pmh1ykHdyifpZijFPnc3Y9eVu9ZSz49UgB1spTlzN
uolUqKG2ICeJ6erUOy/wnpzQL6vHohKEGUtArcIwNoA2H8LL8j666nE26OGG
5/+5gRsNuelj5f3J0kB5NUqMrZ3q+pCiw9ZnPNm6Eahi3uLZqFI0VuqOzXlX
Yer4X5lQuhvCzw4XWlJatqHKEq/eU4e5BHDZteczlwVR1oQrj92bkOslEgcx
dX40Xgqnh5XBUPzJuy5uSiWm2WSwDMQxwDrdTqCG/jAtLCboWovEAc+L6U4P
OD6VqwBtK4W7lE4DmQ28JRTlnGRZqgFjTh9xO1CsM88jrXJfvLmFYNtrQvys
wXILEpJgKvVddMzcYi7p9AMNnNRsI1uF6wpAhDiIyuO8XaqF9GAjdsH9mcWN
QFRTbLLBBEtun3DCedwpw7NbNH0INyoDD4+tWIvVw75udee5xgOabC8lj5gh
oCKEzDQLsNMdO1NbvC2kVKGtMXuZhKCmKHQI3yScwBDmx3UFVpTWprAl1ge0
stPZU2M2SAEixo0aozG5ZYNX8d6MjETafj10WTZwVODVP3C5ijS03B9Lfi8l
MA7S6lGao/5TRPAFFWQoWPoFpTPG+vFYi/cqqRqfv9P6Qar8FfCrXkfSEbJg
rU+eI8M3IcXzAlW49Id2j/nPEGWsee2AgRFN6iEtzFmpmXorpC1pjBLQhuEl
yuVPnBLU76riFPqHUunEzqcdgp7dhLordaD5I/++AoiKtxwHrqgWMM+qwkVd
3qDcIq5/3vt0cFGodMkXOKcijykVDpzxdLS5XWHggb3wKcJjkuEumJyFezzP
/zSBj77rethQ5OgelVFYwKiyEYPYIz7MAtqGOKSViD7WSbKyuWVkOpXDCVhc
gkrZK83WUIGO2o+VjoPTkflpW+iJIxgINk6kmSQ+g0JPRl7s/HizbzpTFnRx
5CheZIJjNastIHF/DPMW73qKHrsVQMSNQjYgewL4ceNutVd6NKZXX7Vdl7Yx
9PbX4vou2cfIR2mMfHCJDwq2sg1Y4zwALeEx+5iOrBtIEpWPiOUkyBa2HAJP
tiXa/RCEyW0vm/Uni7BazazmiTYRPMHkAYcuLtSJaHo6UWXT3CbFKGXzjL2P
kF0ElEXbtyht4l9484Zm9TGL0nraaoJ0crAMWl914F9OynMvGeuMSWRxSHDP
BtWqVyJbnXIc8G80LuuoU+O9QKeYZ6nRR1Auq8qYz9KC5RAdXoOMB+k9svDa
0oGxYAwgJTwC76J3uS7UXLYU1PlxYWTUJ/aP10ULocr+4gf3s/ngi8n3qWii
FqAa9Nvidk5KztPDgxN9RBQiq5g+NQ0WAAzYjvnp7M31/A7ND2HmOPlwhuBx
+zxHfQKJBtLm+bgOAwznpFFG1lilnOFrb+sySdqpvQEn3tXiR1X/mqrsqyFE
GNat35nsetpoamK+eKl3vmShMpbPTKyp6gUFoXDp0Jbb7f5xLaoBIbkUbQbE
jmjFemiMvCpbtRxSPvjQzEFses4Qzv08cQLqlo3VhXwb48Sz71rzDq7gUZxB
2yxZTUTgT5Cl9Fgwv4hT6++DuiyTZx8BFFEmGEXExu+ArpH5Pc6v7vSgN5Lv
38FQpvQQRxFkF4WTRKeoe5YSBEk5Wj/art1GAwF16kSLvDV7Cxm7mhAEXziH
86PmQ0Oh/l6juTMHVZcug7ZusoWT6P0VBeVXuCmcwT6uM6kkuz0G2jmPc5N7
zlzSpusKa1vKlGn8DJqlMwIPDuZUrXmBUtcVADCbQcY9sk5/TFNiwC/aat0/
ipu1fth1kWuph/WV8flJSQXFmhbpTqOYUzvZXXeAEool4VFDTzd85e0izqyJ
r2rmo1Rd9nvx0AMTzWM0c6iZ2Q9ur90aj+Mk3kxUT1c2yZbrJveduzYeZuDh
iXSKH0GGeC3izU6Bk9m1kRu4LNRe7y20YTD6jgBDTdH2D6z+tm0Z22aFJeNg
kT1JqGIBlnh1VtyJCNSit+OmvUI7UeSFRNFDiJL9IXLXNRgjmjLTjPTrqBGr
usvtNlQOxtduffy8bbEWG0Ut0cWV/0qMaestThLgC973FXleCcK8/5p2zsUr
47WWd15ba1oi2a9er77G5gITcKG7DLp1Mm6o8DNaQRwjQmgyg/5Ia9h9/gQu
sPQat0rcTZ0aiA2pbcC6io/JaUiZTV44bZteGsQ1Jhz3ijXsmofP+rfr38hO
iPj5hqS2zH9o+Ne2kefws3Dz/VXkTd7dM0p6CjQCFlH65AjtqOoRmU0dpS9k
wgMpQ9kKziApa+0LrLcBSgZIIPAdV0Dlg+GVmJfm+z8xAP0F0Rd9ZyyEKMDO
L+wXbIZQadSOuO8MREvVqLEH18dTifOGHJUfmSAmAV/9Z0cBfqb4puJ9IcyJ
7cdrT/u/7A9o8MsfwUVq20ict2n4/LPQnlTH/S7vhfMrRexCz2e5Z+f3vccb
2oJ0vS/bJLgjeIk+Dk+Scquejw19fDppkSwK3CLXlFlcFqFiWOiYzBJIrW8h
PshKwOnIXZ0vE13FNrGONMoj5Jgu1IOMcQukqz0qiQLF7ektFPS56LvRjkVi
YlPdkHGlO5wPZaVIcgz5mpE97lMdr+7X2rT+9ORSJmuc1bcQb+ZQFZmeo3kk
F5tMx7F+/ILsKAjh1aA+3uQXJVC6EvzftVZYVzTJhdmfPpznrPKY0dhOySOZ
AzHnlRgiskmAKkRRzAc/uRE61MAg3GhOI2Vmap1wgbgZjfjONHmLyUxHtgyC
gMrSkBUy8owihm87HM6VvpKrCUxvVy8TgXAIA7YQ3E8FWX4RDTcVjX/7y1WS
l5kzY7U5y+luRCgf+GyMpENRQqlp/3oe/wrui/Y1vt1l71AVUYEJa/Jbq/vP
cSCU+Hu/0VFQDL+uMdCLAx8DHqPmpMebNWFtNKcKw5BkI3qEb9sibpu5XIDp
6ZSDr+DV5omxDE3ZdCfOUEbcBzw9nErFU6acNqpJllRR1tPdrIEKotLpEtj/
e2moS2CFRwbJIQg3RjAKOK5dhvCnxCOpbAtojtfQb8UlXiQFUSfV8KjUaqKW
t+jI/cCEYjBFAuhMoOJ/K1v/CTasfjwkHK4VwO6Ep2wSBu/t1ApSC78YkLSd
lCEcWxpjb46jNtjxgDRB6VSFuFtYNUMylaBU936nvMRvbkbMuRx6rkSrf7OK
cuHHoOrSI9gYgRthOM7l0OjOhW5SCKYbj+DKWJneYfXJxb4v05s1akA5YbF/
yJKG8aNeTnShsdMs3UMiF5p0qMG9RXFZ+OIbJm7hkcoCmvWddZQbLEIhjELW
mZ1xt8k7u0nGaSMjUJW9qsQoCG9ZcIOKLNy1qIk7TaoqsCJnXU3npl/HqbN3
JcbfwCzo8p+1mEWOqIK7aR4KIn2Zbu0ppeP8xLvU5kGXnhTd7Tf/3SkE6iwp
kQZm+mVgpqVxq5+V7xfOvBEU/RhEpA4ZAxhxBS6A2XUBvW6pzucXIBXX2dk2
IkELzP3583CLxp4Sh06ZlTOgjQUBvcN7PhzuzL9vgbvHbifT6Nqiwz7dAyAG
pjHlyTV1SLyWkkrCVa2M+1lJdMEffqOyoqdigRNs1TQQ8g+p+D+G31CfCy5z
VZUvOUbjEvWff+Y9rWgMn5C6U5JP11eEcEqW1Fnye/A/7Rtl2LH5xh6KsY/0
BGKFn2cxaTGP0aM8AWSHvGGaL4f/R5fjDyvkS114ZRf5wrRI5QhNvjaIAbiI
n21nCr11MHji53dtcVzeoTeK9jzjITB5suo5SJ0aqHMjJlkQe0dv5ZboTLnf
zv4ksjSt2F7PAE2F8xxJlU5iHvyfLAx0ldiOfuepNbt3gVHkAS6zdxl4WhOn
QXeJfT/S7Wm7m/2X3UmUc4aEAmExDluST/XwPgsXAt6rNctHE9tRhIC6xoRH
Kp6ojxj/xGcJE0xMCdFyN72gWKzdrDX5/XPAPZlx+9ZEot3s5P/N8JAqX6Mi
Fzm4Zce+Xb7WioYweE+QjeJt1H83Mrdc7+DyE+0D1VUl9f+Aq0eWkMAGiArd
i0YVHbB59zwaI87PMPQnP85BVW56GMVI+L8aER/zr7Ppku8Abc5fxk4d+BCh
GzCweEsOa7VglRv6DUD7C4ozttKO1GLModQJuTifx2A1XiaFc14k4BooCq+X
tNoH6e7pjNGhxnlpWSA6DRIpKjxKeGT3r1NCC2dKErBSW53Ivht2Bl6eC5Ng
s2x92BFMbSQcdU+reaFt/ro2OB+1N18Xwks8ivbyFo6wgekmVs6X8Jk+sPZ1
J1Be39ug2/1kZmS6UibQXL9DCUfeJfRgxdTfqzANfxeG++j+oi4u9lUj02pM
vIHL2nJIKXRCnlRCiy5YqCIGLsSMEnfKDmrDcCaWgHRlzLmByaMcDCaJVFPX
AaJ3uYqg7S3OHLkBT+VlxFkuzv3D02nVbeEz0nY6qPMsQnb15ixM0Kiyv4Ij
aHnklWFHlBB1Xwx5zjxmeuqBHqEDxDo0ikqhGs3glNWrdail7+UrC5LJqLwm
S0Eu+ushsMB0bsmTsK07AFVDx0ZqZ+Dzvp2ebTTw2nvXrBSHDIpcaBWrPL8h
lCRrdvtjDF9Z0wbyU7DtQcwbrKAMpo09xMBLXeEPqYkZaFx5VJOz9nEjFy6z
2ZVaA/2Q7OmLQQFO3zg+1squfmQdo1vfEvjD6WaRaiEbnj5NvE36c9QSWHIl
aUnkQCEnf/L3JeJmApY1n7tTNoDbBWSR9JAssbNDoS4pjOE0O+cRzqQv7kpE
WiC6EJIizTwjws3m+7qAHWgubCh7+MGoChv9t+lJEuhAcfMWbUsX3rW8iKAz
8LiyBXJUrNA73EqTsWlm4ecSf/2ggzTsn0QMC7bfCBVMoSax1MF1pl+ruuUv
0qgjO+X4xSn5jiaatVh0kxwMd03CE0CWO+bMQrnDXhiiJJiYbKb8A8lNStHD
UG0DbMNgY90Pzx8JT67y+rRG0qkpmlJnfHzahEVWn/UmIkeZzUzdh/nTBKV9
wcYR4GtpP/RI3PSVWWOrqq6fDfgMBHyY7l87J7k2XAfOPAbpr1kowGbzFx/n
mC6dBbXYJaXjd+GD48P2E/lviXM0l494WhqekoC2GdLGdC7i/mNWGv+MnCUI
lzIpg0ZpX2HIQtSe1PPxW93DmCwrgfwcI873cIgDgVQKbTA2da4FUIYJYnlg
BM/1Bs8vJtJ2vHyKbp/KmM6MpvccAd5dfMyC5LO9M6hICsaorVaxi38dRvyQ
TZ265JqRWLivAEiV6mvaRswjZBBX7g1XbIQzSmSfjK+FSjMFdfBsSFvAkTq9
V6zX2ppwo4kyHVAvxI+/AhqKtj6yvlA3reymWW7+5n05i3NRZxHwMl4E0NdZ
lzyGbLY6DhnN+H1n+5Dj8UpArqts25PDvVYBabh3v/dJX/UOX0ZL+EXUnNW6
4APpWhPxsUZakG4szzB7fO0DL9ofrfwkldq0RyPbNKPJVMdMT8WnglXabe3m
IXDnXdH5/Hzxb0xxlzqcspNg04HIICoGUEMHvYLUhx6tsQGZFAOU3URO/G8M
d4GtrBDca7HpJSNIE6hBvSop6pnOo4l79Tf7QzZkujWuyoPcXDO3XVP5zTKc
oKtj/XGvmRcdSUzYHoRDswLvdiuDiYQtHUm8HGzFvMSihCsaUqoaFv5wvYjg
JB3fAeyDGJDGHmtgavFy71jWvfuySl6W2TS1DsqAjXx0w8RSH1AbzbYGPIG7
qnXl6kuu5vjU4/Vr0ZvOrsRSf8eNmJPiK88Zse4kLG2i4Yby08SisZRGTZ8k
1bKlyhMagLHk2dgVSg2RNv/zO06CxnDxb4neUtkSmy2dzytzr+8sPKUczEeQ
/cz3yHfiVKT+XK69g9M9DNd+s8icIruqGBx2SnlJ8noTBvscVJrmONXnwFoF
tSNVu15GLPevWR4o1zKTOsY02QRFq7LORNZZ3ePmBD2a5nwtjQWBR6aH79fr
/Lj3UWvP62oi/5RGF+zRZ4L3t9V/nEecWSFoksVSM2KS4bpYH8eMT4R2ceJ9
9dLdhqYkDaKd3x389slQL6GJgQtK4GRj3HsyNDCMfbYLfJBQY6mEUMwMshv+
isfIBm9y908tQVI6hhSI//HAyEhRTdNs+oOgWyr283OGWQlgK6y5SWsNmxSt
DysL9WtanbCG4LezPyJjlETsGqTvnqzVDPNvcaFq3WE2N6sCgp2G0+gI3gup
+wUiIN4ujSoG6pmP2cpWC3gzKRUibTxxyB7HnzlcvaFBVFvdZgw0iOByFQtG
BJrL3PpH0W9ncNBLjNJw+rL+TtI6+DSzBqRRK2aOLE8KYfb0U6/a3K71LiWb
U6AhWYMgNISnCslO/4GE2WZJigibRoMX45POjM34lGiOnML4odZMDiEYuv8m
CFnFmMZSiRNFm0JZycTlnM8Jac4IHwyg4Rft8EgTak7ixpo+LDnj5ZAWABdK
ZNkqv+qap1XRy+UshM3cg4CHiKE4RR3BfpYN21fW1bB2Jbm7SCREnRekYpUA
SoIYm+NoeiL2XpvFRKAM51sZEh55fs4h/cCDOpJ6YB8z7hkoAipDA2/VopOE
S/K1Qd8q1QsyBKaSATgqv7Ycanr1EEZ8WWqcTB/JyzbsfE9GrI7Br3wgrowv
dhDBE74dSoCGsfO1Q2oFVtrMUFa6dDhQbTln2mMH8gADnv90wvtJvC62X8AG
bipS5GtU6bhnWtM7Bt28ccMUXVvsTXjDFqbakd00HVzdGwUXCHb1Xh5+Tn7J
XaS8ZiY0kcA94Wv4FIp0YwoH1eRqm24PyRjN4PJgzXNsEbBzqLi/niRPp891
cG27yl5YW3hFFO6glKw4JvMjMZviTPupl62M/SjhHYgrxiFTi/pYej0FWtvX
E4urGLfeCN/oskPlYC7/EbxMvG0VXGJC98dnsQriVwfT+HskSFhJFPxtez1F
DcrxFqy5ZYHZJDd1sECsTsr/enQD0B4W8SW+e3CEZlhSEJKFtFbb41Hx9zqb
OiOPaq1ZskdCISr/Qtw4qA1aeU1Y3eJ5wgTcSAxofZgL1R9s1zFq4vPALHQb
KJqBDHpjVy4AvwkPOqq83dXWwj/dGUqNEB/0Yc6P0A8vYztUxpw52NcHR04A
+sz86iNj9W8l73Ga0rDDUbhGdc+pRyGCIQGCu2QdAi1qONvaR+7TZHvoouUq
0w+HxOldclPfBHQoUBycB7dL0EGL05Y9D+QN8FansZ5x3AQrl3ezPuFRa3wN
RnRaoWiicRkgjmxtpmJt+rpUmpVjPxhq4IamYdE5Q5JhI2nM3r4Mw4FBCpbr
3fgzaDsalrCCBYQyeNqRwDp0AjJn0sDR64Xg2ohkVIEiHd0KQE2XOytE/RwX
Ru+UTNTkSdJ8GCJ2dglyO61aBnf/T7MheR9pHBXEExwxs67FvZ8f15Gm/Rs4
554L49aqduCwcsQEuIqJm7MFlIfP0591tQ2f1JXyM+p8hur/Ki0ZrDGL6lGR
nri76j8L5klUYJzWJxjU1mETEobzQULRjQEfGhSPvW7Zhr1V3FVW19jJvLGj
JamGHhq0e5jfORshkn4eRf20EDqBwpvMhcsxDCZx+qZXpHgUK3EfYE4dqEuR
9XnhLUe3wcbnpEWxxnJVZ06FB1PwL/aKZ+tmyR69nWheJYyVUD/3cxnMnkbh
+lXZCMx2FFiKEysCJO/v+eDNzo3V81FQG+u9ViDipCKKZ0GNEXuWJIdcpTLA
JZmgC6/p2xKg5sZuamRVH27icEGo/BCWHVz1P3IriRzvI9fiS8QL6c8N+imI
51OJ0xbyv+f5EVk0tyXMHYoA1V1grsg9EL9iDq28PVXTtRSbNBuTNoN9IGzB
z7hXvrqjcpptSkxr2CAe5PixzApFHD56osUorc9vf1TFmIZJkeIn5b3hNVaa
iSoriROeE7XI/pJuOwLd1v2KfoSGT3ThtfeSy3XtorJr13UjI6o+iWtugRgQ
Y4aDo69BZZBifq9LGlIPxBuqPmHFDTOc8u813g93dPWxu2cq/XI73akqRKF/
y/+i/+5TJ4ToeOG6rfikgQ0kyRif2oyQasyufsDLATXN8X824oyTNrp++xjF
09hYXc3i0HVBH0kM3AdQZbBrVA6ezZ93f20I9CgTY5H6HW2LBIg5AxdY1Tnf
x0XkwC+jMpAr10c0z3MpZl+u5SIyPWDbVusTlXFcJqCxGZqxGJDgD/UNdp6m
S6beyozQl0RRgNegogwnDWk1rkBxqJaVkwt9/8OF5jW1amJxIWz7zpIn8AgY
dCGgkNb5DvCZN5yGk55buHBwm39mwyd/NyWgfu61aWKd9139csfBKIkCMFDG
2m0/Nw/z0o40o7vmP0m8URru73tC8LlDFN+43ADcEmI1svMZpDmVHO2xOGM6
HdgG02UFOAYyMjc2XH8GWT6QebNf1tj+u1BJzvKP2bhhEey8CyHJHF/wGPUA
9XIV3D8KW1pU8ytyUHKziWn6oS4H1L/Fzt3Qc69g0Jv7lGN6i2kXRtTPfhXc
hjEbGIBwFJ0p0/lcoiSsnXFKQX1LXVJPZBRs/Gy8AVp00EtDOafQYGuXffkR
hF2UQJqSwhrtLK6VHcmj2ciIxK1x7bbN957MMo9OzVQbiOlKj9D99KJIrJpc
SvI3RXOWhXLC6S7MJ05bbusY85ClL98/NEqFQzifsVxHmx6eX9vo01VI7jGj
DU1q4pd9i7kb33yccorpMDlDJyKxGuovYaZfEcjlPxv+6mCAT8vOmQbWQtvi
dbeJg2OvGpjrX/4UUqhhzC4pb58xom+N7XMYdt1OdoPYRkLQgSvzG0+I6hHl
foh/oZ6DMnTYDpeGrt0q45250aknPRrhJ/A1nutMlBGQ4kUN/eNRZ1Zy6tWW
p6f7G7r4LRzD2ogAGgka4+6G9m54kIZZAaokb01S9Ppboh6qPoDnWjdCHgwJ
PihygYehdajk6hvfceMUtQESJvR6VH+4Bz7sVgT4VjGejf7HpQ8XuYYMDhYn
a1WyF8QgT+Vugq0ItYy97ii8eXJbrLSTr5RmG4HigHBLV01+FvQ6niOhuTRX
e+muExnxlXblr8XvhFNOrWFU1d9jKh8y681T4JuPob6bw3/Go37R/1td1EB0
EegQYstDTKD24BjGZ56XfY7Qe8X75atRiSNRgJ2jhy2Bizdy7w3PlRqBVBiR
jETDWFtWNPNwsDPnvY30dI+HAWG8/1bTCLxSNZl8SZJen74H1f9dIOb/WgCX
YUYc040/axUvruQ8ohQk8QbB1VHrMBe8x1hgAUEGaxqXifXD14DgR90yfaEN
H6edC6FWh8t0xTMhcJ+sT/gxR2mmprfUVDT4aXtDURx3hKu134dExhdmPBcc
1ayW71bQM7h2HPn4h73gwdCNHWA1t6DC/wdIlqI5WYH4oPQOTlzzC4looaNe
J+78+cf+gpLUr/gQ58I4zUPUnzuxvEtkLCSC+dWV5kq/B4AN7gLN4klT/YSx
WJspw/Mf7icQ1XKJoXGdOp7YIGbuarfR9JMIO56H5VsjdpZfr3lp+dv6UuBX
MIs/rQ3SX+/CCUs1SSb6AqSODmSY9oTdU2hvUcDPrNekbF8UGFS4mumZdicZ
oXVN3zXBilunf0rNQjX/5g0F9hcYJ6GegmXvoFnqPXAYC3d0s/yvqKHnwIB6
0nu8jsLHwLCGBx4iu3BYETxrYoaPztwSqsyULFO6/YuhHXOEJrfuE6EAbgSc
tN2cPaVK7dCW/JRwvAtr9YqesZyUo4xeCBbDw6Xy4vJezhXfe4YzBc7yW4L4
MtKEZ9/raTprI/0xWTTJ7TFaBpxLOdxp9LBOu6c65ucgHtWweaxogqXSEOBy
kqM6C9LV8XsWKUI9sdKcoeazzEhZvZ6REgjtHtYy94lA36liGjawtt4VYc5N
/It5lBQyq6ADd88OGOWcSXTbdGLuESpIeY3ATUPdkD0SL9zyTZqkgP1ZpxLB
MH+Do5q2uPcqxcMpl3b7LU1Hv0gAzJCjCcnrL1XnMOTK9nmv01EBmz8kGd3u
ZFMvtnfU6gTXx6SkRG83H5Z7OZBT68a5/LgK8RghRYcWPeXNvRbtb0XFPxbb
E5fNSUbexy3S2cSp6kQKk8rNsoBhLQk6k6j8vdGWwW/51ueY49tafhzjpX7B
We0K0+MAFRQT618MSAuRMmBYAmEU+6l5TJRao5jhvZoWWQCdiZTCWw4Ua5aX
W54RemnWQi+ZGeYDTV8ytWOWPhCoqiDPLtW4ssJld/i+W/j3Ns7UuGAk5c+d
7hHZgMOL4EVSQWQCjgKOWmCkcDaP0mx1fm7ejipAgrQCKC/PKG1xNLVMwz/5
kJhchOQSTVKXhb5WHHYWkI81MJj4EeNFDXXeDa3eXpFv5waJFRuVZs3sLbwl
N3iP0HxqNz43Qp710g5+EijcBEB2Nv5NLdGCTYV9Y1iTqXyRTZuvlhU/r6s3
uqCyjROqbzNa88r/M4ardF3qIu11Wg21piOJCOfeGyRxlISuiyPRS7LlEtOF
cDtXY0G+E2cPuW/FoxhqluoR/klwN1bpt3Zz/RbbbhLbWMd4+n/NxqciTXOJ
5NEcYuP/UDUJSYAj7jTgNtHB1+sWjZVC9wUxWEve612eSsMlHkEbIZDOdcL+
fEmwxEAFq0eG5nqmhGHrWTrsyYnqO3Y8a2lgtX3SLW7AUa2H+EzN+ib/+Z9T
gR261xw6WaiGSwwFnCH0Hc2FAtZLo/Pv1cGBQgkWX2r9l6FGsllfCP7o8Und
Xj2ZdB393OoDX02ncgzVEJ0Y/eXcmaLlrjDjnaD3Nef9KpFVlziN+HJASX0N
u7lAqjGK2J+xd4EYmYqsD4IEk5U9xyM8qS9ZkxT4c7SK6nZ7Q5srdDL7HyPl
IZyQvBdCnE6y/teLUR1D3pLd6sETsQD1hS2pu3oHgGx5NS/TS1ieNzkHogL/
IqKt6CFwwUS68f6SKNMEUyC4gYTR3MyCXJgFHVfJ4Cm+zsforZbPHQZO6g08
hhyg049+kV+0oFOsjaHbZqLUHrOyfeojY2B/MRlTkuttQo/ARGPiMEjY58UN
frPqWtPuom/h1azes4iguC93F0x9wduDSialGi+sHvOyrCMikV1IQ1GEi/8r
Zsly4CkybB9wW1jgXPC/bQQ51M4IV5Gr2I9sPxvWGmhwmknb9itFAlhaRrMN
3LY2XszLjlyqYXvUps2vhWMohbzn6YI3nIScypMhtoAPSPgrdGOGshHyk2NA
Rj4fsI/Xay/DO7OVLJPhZKJxtFBZEYYE+5Kdqf7XK+kvFqXpvO6QQ7DDdZ0w
aBrtq5WC7rZVY/df/eKsEOVVn+AX3fy1VVbVYA/cbNYGrVdULlLqNWCjZ+td
nazUgmuM0wTNiNOw1Z3see669d/WGLiaf+YaBQ52XOClvwWAt1HMBwkulCKe
HnBagnaeoZcWfoemUxNepm1M+jeKM3ZIS8qsdPEs3HrUwHQUBzuMmA0WS5Th
tKXuybQynW+wTxkbCJk+LSWHyebkz0eKYL15vKcD5586Xy3jH72D9zJg78jB
dgpWTzwXIF4Q3H1sWep0vLgHCQ/kcBnqF80hXevC2ef6gBZ0xnExCS7+EeOE
sPnr0rdSrqbmZuLt8iAwJ1LLavN9QKyyI3lvN/dHRFiLmOBUPVcUdcbnJN0p
wb6qOYSaH2FqdfcI6JRVf1exIYU3DZrE66GBlO3Hd2Hl6eaG5c7oP2pt/GXR
yzvtjuTO6cdHBWS8EBZslMkpJmpWLKVInfTM4JGRUBCF8bQXru1JwZgV3DWl
QHXJ4cvrm2rnZzQRvkcF5K2+oVITDUdA6FG3kHQLUNGGtxXGfZ5v8NRjPkAY
OUIePcmo50UD9olAHln1opaCSX+CH5HfXxJrxDY5gOXXRKb9vMG6NcDK8bpr
KiV0skghWLHRxwz0d9lkRNpVbotPorQiqLwb3kTPC+zcyIOn539CLqWNHtqv
+fspt1r5Qe4/sWod1RnKjdid+QCG+qixVxZ5zo2pWeznU4mJUgiUe3Tzu7T5
1kKZaagJGDzrjStKMYMoZEV3b/Nu2KNtBpIGaDoXYQuvMikkfrwgd7GcJdkV
B2TWU/Mxo0vQMSGbvGvzhlJ5SQ12XKXMv/SdnA9nbFaMY70APHG8S2drNRso
Eg58nSpq1R6cvcLH7dvtYHeP6g7hx3Zm/S0YPXlfespWIo7RXbN7j7I2NVDt
Kbr516IjwyvYKRxE62PCJqiHl5sXqZYBDe3Dsvhpb5AB+zCrzzcX0ifR/sJ1
30oQaqeS5Z3zVxMOUHSS07TRjRLBqedT8UvLb2LssrWzsVGiN/ihFPBWjoI5
V+9H+ZfZDsZ69nfKthpOyDi938JzVcuBSf9Shpu4Ru4Oycs0+I+vH+luL7na
4RNUooHJavKXVXC1f9QME13P9VzTV3NQYhuOJm6/868NZIhaCtOgwhJFWooJ
x9m4i5tW5yZNwYth1a2PXMfcX6G6R+tWc3E/ulJoK6JSlURTUrLkTjnS5e7P
S/vHEEgIjbsHXTsJz7TpKcfJlLAiQATAEGElyHtILXg5bFWAaYp/lly8ju0J
NOgPVH+YNLfooBCv0taosCDQc6OUyzTn21mAjKAbrS8zIaejXT2di18tIOZ6
T3H1jMKFz/364JRRp3gwRaNWIdrWAVN8lCy3OcgYfyxcCYFJNQekglJBv3NM
atW5T0GiuW+DxoAR3JDLBYHZvBkOU/OvQOkayXtdyzsBsK2+31iaLf8pYD7w
HjWBxY3BRr+ZlhdECLS1H/62LyVqzM/05rgKV0lr8ZRFtgyejAhM0LwM2h3Z
NPdGODvsWnVgyfdN2qRlxCQd6JkxbqQWxND0es2TyDjezczzFXMYq1gyL7aF
a8KJTf/20D229SmLLcuXO7IZrieYHGbGt48ORvl6zzCom3jFV3ItqicxO0iP
og2nq/N3E3j8wSVEgY6s7MTLjwdhgfb6Q0JMAw7vJipagsv1/XBIHq3Pq88f
EQcNmzWJMxMjvxMTK6JCe5sNu1FL+vRINtGtPFO85AhI31em/UOb+QGiuLPb
MOOmlzA2RheZ6fef0OX19fdbcHvcq+04nB/G5ft6Ndq0gusWNqgu1ws9slMz
eW3CFlrxIUaGjpvRnOtgXQWHOg24tT1EDvtHWg5pGZK4HwADl0gZUPVrwB/d
IO6z3axqXxvuGsdfchbGw+2L0CFPNd2WgawOcGN/DH/tgU4DAG3TQOdqr4kD
z7Ss0F5TTC3BXwfICILDDLJMcO7P2WEn0XBnf/EDdSuKwUEf0gXXrF6VmM7l
EKK23vyzvWxlWjl5SQCoT47bC86gQ4N4rQLIz9QscBTxUfW+Qk9R/gY2b60t
DHATHHAnr3fCtM/BF6hZnwjcN2Vs8Y2b2IboYnpY4tRP5GO0lfRi4DaFf/SC
zuNS7sZTbjK3RCfbPuq6n6TnWwMptS1WPtUUaFrNBnJLYRkDuJl4zFkAV27w
yRiR8RZd50013HqXVeqQREQeka84kwvkiMWQ4eDV94tGmIQQchzy1DDKUO6x
69hxyGswJfk6CfLdHn+ENnIPrR3/Dhad5BrWbRBJqfn33YDbIZEEsov28E8e
1uKoMuIhEWjTUKPaYYbuW76CLoWAo6wKIERDT0aYUXorm5zxMe6ivBeyYube
x/SndGr7puYInmuKosXVAGrikxK4csV50xbAJrACN/19p0F9QzCWswjGeXxr
ndQ04LtYJpM/2gOEm/YkDsTJb39Lb81AEnGqPlB5AP7K3b2oePKBnf/csPMu
hG6Gga7h1ldD4Y5FjsALaR1gGMllJSsbQqp19L2VwBNqNGyezZM0CUBKyWQy
IV7y73dnUbEHRM/H/7OtpEuFfBn+rqHCS0Z7juXIExPqjsW5e1HcckcQmhzX
XdXjQTAp46Hu3t+OuhmgcrOYmkUxyzgmkXveYDZ6byiDbuMEqYSVmvsLrbUc
DO6DIWd3Z/bMttx1dd80ECMznweChkbGgvmgBw/ZrinXKaajSvRsNM0Cs6Th
IkcP+F4GTIoQooMg6hjkKHr0Nbyg8Lhq6X0cD4YgZWGfcHCbwAM5BSuUVLv2
Pou/MLUtBzl0LkYjosXMrJgVVlVgHGRqlNkCq3JAki2kCA5yNWl18gWVeTCu
6LxNIXWKJZfYdOjTNw0zzxXZBCYwKvzmTQAyp4ZFonH2DdnEnQWqt2rEs7um
9/myZMKHi2+Sa83jlqAgho5kb9c6gvSYcJ2vTUxE1LB6APT40K9mCPlTj/Mm
uoG8+VRuAo3K1j13bBiWfQmq7wQ6mJ7O3pCzFoz0rh/1B0fLKHAt0Pv8Bf4u
N3zAXSmUUfMEC3w06lpLEkRwmJ9SAz2sdo8zkuJqPCYjAA9S1km2CsgbUQnS
iqL0C4YrpNhzXdf/gTlEZ7zL2SSEo2MUXLmNkKrSS0V/U+WqOuBHz7toXwAt
9XMJ6/EUWbcsqJy5jqaC52weDU1AmfCU5JxJEnyewvZ34pHE9NuHqNtfdSl1
AiVx03M03GjVDMJv6hrLabGOgyzvhbalotk26Kz24pKDKTnpWFQj7s7v1w9a
DIkbiO5ISMIHG+TeysEZMNliUSPdaaVXpP0Jv+pQswp6XvQeV2B+PhIQ0Vyo
aH4E4++98hSyPD07uM8XEV+WIzYFO9ATAGPfqROkGrWelHpGwv7zpw7IOAas
xETZaVFmgKV+h8XF0W3ZGHBYLEQ6XgPBJmATxGH+27j9IJ3toE71gP/E8su/
78fyJdnZJumKLoax203meoSHhCmMVT7lRKOafqkH2yLjEEZYR/LuBgRFczsV
YfMe/d8bLoRx5Q4pe6tP9R3ovHD9YeSMH4cRl+HrAdiPGJWQtImn3Z7xbG8V
diDbxEUjJMPIPvydjuitYk+5iQ26eSiqdvzuV4tyKqnMa9CJhgu6n/eIg1ga
isGPWvsVGDorbX/jjnQMNRH1O1qK2EwVMPN3l/ewaYXZ8gv/opkaicLyudlB
5nkwbe5VpTtI86qAk7g+2ENfH9mmpwJVayq9wW2Pf9yy8YIh1qtYKm4BSauW
AW/1NG9du7snwx33a3Fc89g4pjaE4ABUtGhL9VCybMnKF1bv7yB1RF75Fpgm
Ys4iG7OXjcLhsmBOZUHFWykst+aufHlMsuTHawdRLMy0gHI39dkCZdb9x+ed
T8KCPQfJIp9+jGTmOW2RM85uJOqx2qqQ6P5udQJMZhdEAXP7ABBriNA+DkkH
J2X5UfSJenoPmm5+LH8Op2iHS5EqjxYZGGWc+tectieZu8J1poSoObzTDwTc
WF9XRgGzYfwsAki+6k4T9/gos0hktN7bk+BX07McY1oHT9d3XBvzKigx3Ei7
p1TsU66PELQ5yJlZ73oMFDZhtv0ch3z1ETcbU0EHlIsWWkKivHMq2wXhr4cQ
kIT6WyAxYCk9sxJaSES54+0azsj7eqYeyLZbZrp0uHOf5o6wRqu4F8zF4Iop
TK+pxBwCJ84S3FrR+yl4IpsTcVyUcdZUiEGe1mWHKYqxbmctrFQLvqMDPsk7
2g3THEJd3Y125r+zBJVqlAPNI1m18oI4BdJdSiqiALxB4q74CI1JVssTgXqg
3YEUC3fnu1OIzHCgGGV07Ff7I2t+3VVhNKuQTAXuTtnQX/rjCvIo6i9uYsqd
CndkOaNnbi5yvDndHenXIY2V9dBFejRIoxpbAJ60lzZ6xs32DqIOjJaJYf/4
ANggZq6POSorfjZ+OeoXgTy0orkM0sEqPDhNMeKbZwh6aj0RykUqQKrZQlI0
EEF8ERzzGocRXJbwZ0pRXtH9NZi72oZMyekj2z1m5IaCRahee2aCdC+NWxgG
g6Yftd/2Ywyxp/tDFOwWLPHKYpR5w69mE7LisfRyAQqLTYaMcMWTMUkowppP
eXnlCW8cS8iAkvUY4l1o7uW934mpqgjV29pVbwygr2nFLuGeTvdzdDAOrF37
VST1Qwm+QtiXuS34zXDqOUYbOooOGrWvoEwB1F7lZkmq6tkNXp+UHIaOZ1eR
qPx5VNzY40ai7G3UYJ9JdbT0MLWTyvHDD0NFI72RmwOfOCsBjn4Eie6rUUr5
GOCvmOjzhkUxv7qsnBl4QrEpLv3lnAuWIkDfXcIlj3/oAD3rsC5O9MLxoRZF
ibzAtRSRbD/rCMtalkEzdBcT+y6kz1V0tYsso9V3tGyjsYRhXEY3MTJizO1a
/YjIKbDLOQ37Evpr1RdiFW6DxQd1LHQbRkZwq10Xvex02GhLdtzw1XZzKqc8
VBcmVu1J/1R/KG24LnF/Rcgt5iKXl93YMCAsnopxvlx/coY+1UsSG+JhDCmm
kc6tmtOjFsty9uArf7cl/VCT/pt72souUws7sX3sCaIxt7gQSEGHmPJyBGJP
ieA63eOmY7tGktmgjMeKcIt0Nb/L4cIHqBQzfV3DBWRvpw/z1PZRQOOEkWh0
CzFWXMSvS/JM8dRlmJZyquz72li2Dd1THhdukZOcIeIsPR2lEuxlHNrolVBb
Csw0gGICRGEy1eXceRWZ+TOisLexR2L+VsCQrqhty7zl0xs+qO7vFmHySOIt
h4EDy+C8/490TZ5WrEIgePZ+10Npmqs1yRNnv724+S1rtvHVPzl4xwXpdlyT
Z2vTbzf5n23k+bhwxTsX+ED4USB7znWO+gWiQruDyVvro/R/WeRSZf3oFmpd
9aUG0psaHqDfGNoi3rpqj2jYUEbi6XQkFTmxV0zkw6jQ4HD1v0A7uuE00Wem
fvxay9wnY8m9wbtotYCNpZVccZaUCMYIaCOGnxDQpjJmL/KF3uxhzk8a81of
rnlKV20G93MqTO5OqGLQVYBiB2QP4DfS5xHfGpP0Hv3zThx67FdNqJ3o+2Wp
gOwX5Wec5/H1AQLWbfcve3KXb/PrT8+TfLUFVyrPY0bCiwyOB9p3dJx0PV3U
/MA7Gt6pC8tBgB+RMYdAPqt1gfggkUJWkk4aidFQf0jWtco+iUm0SWKv5FzZ
AAyYOFoLj18alyqElS84tPGDQEDp41SO3Wo6YdGR3tvAfoNo6mJ0xnrSKild
9QAnGBr2FJYr1Fl6OiE89mR/KgvSpBO8onUgOxXHmK9qNscqopYQ6Yge/iqc
1wWv3lAMSzlop6Y/xQ7ATKGAd2ub35i2g4ogcS8cL1XNynDScMGD99ZXNa4o
MJd2pfDQW2c8ySdupijKabg5aLSXGfWNoqhIudk+X22LguEsgLHK4VejpNPR
Wl/UIUNkmDtEtgzyUl7ixC5ZUq39/J6wuamBuociAsau0nHZm4S9XpUf/9T9
c74FiLWjYbgtDrXiNA9JNCOXFpmLcBV9pNb/63ks5JINpQv+B875K85YufDo
FY9vsDyX6kLQH/dobdNDrhsoeQ5POrdoRRmLBsyqTc/XYf4eAAYtA4j2uHHL
Bww4k5vQQihwv/RXexYtFeTpOhNIoKLZHjbksw/n1w25CVhbJjin3b1Zz0pT
fB7qqOj6F458Xk1b23GjMuVxoHWyWVxJc5p7RHTZUZWOPHBHE5N+LR8jWtjB
zycYEofo6kH58U37XBzPgNiey4KYz/X54UqCy+GT9Lm6C6RyEWWe+iPWf3bj
OQvhs81D/jiUmTxD8VYD55r494bhKXUafK/YnLXUva3RsJTNsLsslZmFq8mA
Gzan8rzvZ63dOgava4RBeazLeK4+lfzBXqGuTz3epLZ/QfSay31eaoF0K3GZ
XBCSx8C8FxXN81WS5q+7VV/eHrlMXWbU9ub2dP4qCsZ8+DS/ZSNl0TYcmv3r
QG/B4kcfMvBt9IrX7EhLjl4BvQcoNTqW4J0qdCYrVh8LCEjiwjimsj7M+8Ge
yVfeuIW8kUZ5DdtfuYHarIPuvXnbvyE1JBMmRAcmoWKudysGOvYqhwRUjuHk
hCH//G8+gk5YEZsW95hGo1bG3BOHpFpDkLuY1VfCxP7/o+hqZPG5Wn+y2QIl
k/+z2D2V+cpHh5suIuFNuH0GjApVYb6A0G7jqT4clo772nK3W6Bw9DQugLRp
1oy/6s2f4ptnylGyi0ri9HMMKDfCcAKavukF/pTcoqJP4dqsf0pJ9g2YASHk
NC/g+oaJMDXbKtdmJO9Pc3OlisPOauT2SDo/ZQJi2XPqqkXPO8S0SdO6Afyf
8y1jAujxnOIgb6LUi8nbbuwT5NM3DgGng2dW5r2hqzNnGneVYZ5KXBa0cTB9
ymeYFUz4fJwZUVvKAFcpgOMv8i2xa/ioGow1m8IuOwGiS68CPlLuMTF9xhYY
nAIWvLSsrAJD8r9LgMMTlXSG376EEOnifjI1CRVTPzt6vzvgGgNEelmYBwf1
SKQ0Ahs+RP5Xi0GcJeqI/b1CvASl6gaZI7ZMfwZpA63H2B8sXbHhjWWhTL8C
BcmC5PbGrxIOWl8H8R3nmBRIDNkELjUz5kaJfRcatDXKuUTEazZ2QmylxrqB
kpOUfBgqxZ2Eyka3sJRJb3IjoIOE7zAECqnst3PCKnBXmCNXLB19x8uOkvjN
qC5jmS0syTTpk2PQXCVozTuFjPi1yTBqfkXFLl43Fu850MIOZaX0y20Ficv1
M7dAAl3TeYkmDfYtgKloPbtRmusb09bVO34cqKoym2ma8hyo1ZlHsPW0a7j6
2APskMozDMmJaNsy5QKSPMvpnL7qwXpj200zbLz7nXrSWG6rFXKJQXBpqeox
TyPJzBN1XkNU/sEjCznuibGMfNB0pdd+UBo4vylKO6MDq90L8u4qIL5LYEa6
B9av57f4vGZ2ECdumrnjg6BoB/xy+KctWPhqEjvcmYS4HLG9PX9J9jsnnteJ
5mtwRD53BPFD1Xtpvoorm9g2BAG05i2wero1mj2WyZ9iYtrl8FaTMmixLBUd
unUULBOaTJDd8Fahj69UnVGtJ+Q894MNiZ2yTpPirUbUotr/mjSdSzuuxToL
hsSpdrjmLClRTNFX6arZQ1ahdXXF2JI5QCCIZAt9yAuvnjTIM37qkSXosiWV
/2GndHWp7jVToc4kvzu/RC1TAdnqfxlF8QzlFEtFLyjDVdKzYCVPHwFp6q8V
CaUK/LmPn64LGDqc3CKdCdM1FVVISF5HsO/Ld5Gwc7dJGSHCIPBVCzqPFWFc
5uJ2KxNbRJWhb7gOEgo/uH40hu1qNnoTwTBquFXkq/ynj5joQTQVpPyt3UXX
DHVWrISnMrCN+nrYGxBsYwdfVDDLifcQSqRkiEW3JvksYJGxNW0omy+7C58O
9FHtE7XG7ih/ettiAU8BEmDc9PpYSHn52QovMC6GzchzrwmwcdXEtGiglicu
f4zDhLDpta8PsXdVcUR/6DmArLOjD6Tf20XjWT4uvQfjw3nsiwTnbsXRGbcE
FSgZKMkkIr05gcJb+BPT/9BlNJqdoswzAC2gBR/Hx58ogxrakNCltTpZnFdG
o28wV6EHhhtjrBuXWUIRMqhEOlz1d22v86DMdzJK0jVJdv5glMzjQzhfy3Kv
fiyxB/s4nHjgvlQhrFWGL3r5xflpRg3AyG7lJkilW+5Pg4cnaYtwtbqfVmKt
asbMJFden8p+9+ovlGEsSW9yboWO+MGm3IWu1zxRq2N50YpLkJwW12zzqi3g
nuCUgRDdELfeuSJUKZ5ptQ8WUvqT2GT/RC62RH2To7OQ8cDQ9SdnsvvGuxYG
lszm85ywQ1EQ3/nTxeRoGKUvYZ7VSKjjjwLegsIAJVR9zEI6vSg2eLshe7pr
bzar7n8oFKcm0gjfuKx9k09rLXXSokNj/+sjVymKIGPFGEfDmVU25g9wwlxv
rc/lWPZUUqOsJdLcacqz7rIEaXm1gEVMkYQN2/2HKFPW0ufkb9WK0fXFlFBH
cL8p91n8xOeyf5IuFc3+Rhf0qy2490hrII3Dcul7X3x5/r+o/SgAu94PbahM
9LwSaEf2bp73hE6EvAkU5dnTiL2m0toBt/21A16Y2ViGvk5IEbebN1iDi+Mu
LqmAEky+MdgR16yHTA1dsS/DSwhwmgUZl4NJks2LWfNhLgLv/sNYgh/kig+S
n1hH/0XDq2EegVpsQKSzgflljuSqWfOX0UuTXZDn3myZ7EBu+C/uNCOoNY1f
AeMeKzWJdW2grgK46NJE4fTw2UOK0ewWanCboE8/j2u6fMdRgIUtSfjHCX2i
YmRGleo7BywIFC/dgTtmm4Ji70w5K2GD8ncyFockwx/iw/5JIts6eF5yqf0k
9HQfeTojL0+/6BB9M3B7KFTFo0ePZJRUsSy/w/PTaVPLKogEBAk0D8NLmoVx
nQPYFcPoy9aK6XEau63LDA+6VWp7FFBYXE3glbtnk20/o1jtSoLFhvXOeFKn
FELolx+v5RpQgLxaAgomFYkMjy98XtJhOxZHpHAXxRXB0QLM/0zpV2EOn2/e
+Olt/ytX0ZIYNvSbX2Zg1Y5EsLxIGowQOw5ksJwcIFs0Aai9eENR8yVc12WI
obh7fi06nFHny55COF++tOK/p6caqbBI+Xfv+gZ6UWu8Bot0A5yIEoNFdTPj
nm+DvoxTYcu/gfSIG9XME9rVFGxl20YBbBCgeFb8TGQSPg3aWvMudpNYGgby
N5mE9jmU9AExQauGPp8+0FGprw/WLhp8900iBtE1xjcoJYJdjC+Mlvd00zuM
/T9zrTVVWnj4vGoPewWANgLjLDyV0BfzbTfmZVfLa1GvuZBJFkj/TsZWicK/
KnGj2B3+/KvLn6aSBLf8c797uZ5zvZTrCI4of/tzmux1oIB+FOzuBKZQUSQd
cEZ/7COy9j1usx7ilkxqm9RlmhBGhjVcyz9GiVDSzOjASds0IyX3LTh3i7wf
x8s+MP0OQIlkXNng+wixtQjwcDDE5NiyNKZLLGgDIpVcapDjwxRUMTla1/Ul
flXh/1cw1ELh3yFKLdl2jBHvPfJ9TFW0MVE4q7rc27Myhf8nA7yuGQf4WuVk
7m1o0cVz0Yok4EzXl3svbIErXu73bxN5rMm19oeWLCpY5SctG009SKMT0iNT
CRvogsN2I1XuGes/l8xisuFpgDCsAN32sLsXk+6N7vyiumVnzd9lddbVOZGa
Khy5qwWfiRL/r5hLmnjm6C36jkwDxrai0YyX/WMGugoTVkVUGT0rzEXwDioP
g8IQ4v61HqixEu7bKZ2YycN5iZ3bguOlhT8v19LrBdcbEpSLRx9gQPGtmRpI
q/oPVQQfC1t5N00YmwS3YzngekdCbKzBqSkj7K2Vpy9uVWRxcPnmrQsliYDi
DswSeS7PO8QunPPrJe2u9U7ILr27ox45W2PdETwBfaknmmNST0PbVHYlz483
ApchVQKBxIFDNvcgKOlLOIMm1Ov+N1/gj2tUHtmtyfEyb/giSi0+sM7tXC3p
3OY0UyaoIJsKNC8EZKR+Nht3lDmx8DkuvL3nrArCCdY2e9ZQZAV79HmbN5xo
3oT87x1ptd0/S0wUMdAPBa5J4A9DB8HYbzL2kNhm0ZzbxmacmzModFrQxzUW
Y52B5fwndgAhmgDP+TOXiFdTQrSBee1IpMIW/fq7x2yXajMuI268AVyR6ZHa
bAIpXhzXLGIeOWGddTNOtN2FLunvuQYHs/GJINZokOGVlrytUB/LuNH3gQlE
y0tADQyRR6FhRtWoYciUtnqYzRvb+C1S3tC08di8DP970bQ7dQhPNDA42Y7j
SZqan8hhg8EnLyC68ffqkOo91NTgwwDEU28yXXX62V42n3TpQmCXXlRq8ckN
VhwmkbKlSM5xOqPKAcZok0669B7cFQJEYKI8qBs6DlCEkyX499JVkZ+QoPAY
zFLUMvm9rmKewZ3kXWYvoCA1ygBS3nSMkkhwgJE063qc1PgM7rvuZH6fSRdr
y1xN2+VyT60xE6XqZxtW3rb1fNgDV9tPYRd2+BylWeC8TP3CFXjXzOGK7Uye
jN8RjDdBqu0Sdho9dtvBYXzvlpm2zFuj7DDR1WfcBVZvOYcr0Uvc0w7ZqoZZ
QS+QedmreWhPhRFjPb589GcqFZNIt3bSCveKUAWPofFNyi8tPAHbIIcFxpTR
SbR4F7SOJJA9nyITPf8XxbIrBFZwOZJsJMoe0QUHojugMF74eDAfVImzksbF
Sal1K7cI3Dv23pd4vKxLewjZgQdo7iIwOX9yNhmZsmwlW6XJDo0pgTJWUw2P
jlzprcx+RdAMIJUUcr615COuSRBWxAGBQWvtxuuu8QyslNEL3oMFqdJklB/y
xvo9XjN+TLlxu85tO/VOrl6efE1+CqUOTU43w9rTtzJsYU6NIoTY29D8K1Nv
rBHKc/S1J1LVg1Ln3OkyM7bFcY6EKZsarDC7cRICDWG0PsPl651Bx8Gihnhq
w/yE4XVzKYzR9W7ufEcmnziEpySBKS/MzRfscRtDQK47SNWKUuFuv6u3eNAD
hF1v5rYCzZQiMFSZgjdTYd4KIkK3Qq+NsFX833dK5OpZUr1YlVIQDKoWuk2I
TuyJRF8B/DDo+Mggh6HlTAQu2wyG2fw4IW9ODmFCMKcFm31IarV2TM2oNWk2
iA8SaXihptmZA35cmimMRc1wytZB6DyX/82rfXi6PpZkp5t/uvTM3bYX9sdI
i8Oewy5+g0FieZra29bTif1ElkhXFflMUKCNjPnRIdHhg071bJfsuJaZTA0f
gTW7OnB2f/OilAq80nXYwTHEvBi3ZdAKqzbatvfv4T8NRWTb9bV/wxHthfFs
voLhL3+9M3MzDxehWPUxZ70OEeaTYDK3lSRNB1XFLsDE17o68P/PI7o+gt5N
l/x/POB7gR+8jlEet3eq0oS/nC6S/xmYUIl1hSgNy7vYliwIpLuyhkYBEPQu
ks3wWPwEmIAHNaTFtU7b0W9q7FBAduh+BTuza8Uk7nFUGNVB7uyZI7nfdZIW
xhuuEdOnW+XyzXHuN2LlDjOVHgF9fDeEMCCO8Pk6/3lL0zGYgz2qiPr6dze4
A9pUc5b+FcbLri1B8Hgr1R7ids+TLrpBMyrdINyK9+M3uuk0m5sw32JMgHNB
YlUiOUfpPbAXxec+2E8e83chdqdzfNP9K5fmM/qfKZiAFb7kOAurOYjMg2Ko
rGRseAzgRtxmZExJxZdaQY9ou3a4PwoHUW85+n1CxpYWW8pgbfZp+GiCSFbj
rnNbFfNF7ye8CXk1C5vKj+YD+lxIgtIyZT4UGXhfG2bxLoBw7KFGb4KlHrAY
2DxJ0Bl91DkU86gjZMlCsl3ft5Ccf83ZxzZ7xNOwQr2RArs8A0PJbT+1vskr
TEOQjuPIYunri9CJHHGWA29B4AaGyoJbESoqgTDPOZmdKaLL1mzxK4bAYux4
7JLNmL6aEg5RrHxY6noo6B3f9876zz7b5XNWWYV/Zk91LYEPzdLW+tcmnWWm
yyNczVPCWcFPxQaKPucDc2Y/IdFFO199k7HK0HoFShXtUMMiY/s84pjNrthf
GsU0lhDJRjXgBhSEGKvVgitJQFOl2IMWT9jicMQ9olqazr/GEZrvC5M4Esbj
h3gAbgJalNmBLi45tFWzjY77RK9QHM0zqGzWmjbkBH7nVpKXEidM42F52lRL
Cf2m8P/xv0jOkhj91xN5rKttdfWDZFPMej7mMp6ec4Mesp73sj8gYKOc6gqc
a3fWKs8/YYyhmP9sWg6hSAohrFc8xygG/GIe+mzD+IAjBk8Ln675qbDubmaZ
746E0M2asd9BG54eWJwKIusOEYjf15Cd1uxYpSEtIhKgzQFzH+JeIQ8R4tfT
wVvFyy6bBKcSGtLvxJcoV60nnjpprxutGP3KcAfRfsoNyXpoNgdd6sWiwMzL
1P+2Nx4QPOw09+ofw3vK1OxyoeYxBo/GImaUbvc/3t6iGFJrdkvJxujhx/dF
oESX4KemGyHsgfUOh116+KbRqCnctqdLnfqQZttJIVHkDby8XH5oYcQ/Wjzp
UqpkCsDxvvizvOWQ7Q8DWO7k8lcRqkh4m9XTaxa4W7WhgE+yZkoUKImvlEHU
0kZl8CpULia2SFApmVAM4p6rfsUK05DaGyB66NruZkIFEjWNhhKNCnmb4UA+
iENkFmP4YgRrhos8J+BA893V6YhQVX8rouVj9IaNh1++S3Vu3icr6DYJVtmD
bZ0/Ys+9gt5ekTuCXLM0G4sCBaEWaJLcu2zbK314gO4mwT6rNNcHSldHH7tA
76vG3V8ut8Nd6USLwRqrQHP22zhn61tHOAgp7Nl/HuKO3aFuIxM3p1YZ3SuR
/ETtkKYzakn/gf6fbdYEp+9f2rxjE6i4ZbJoCksw+zD/OgUcsokG3RmqQCvc
7KS9nf32MKiYv4aP5Tway14eEjkRd9oOOzsG4KP4tPSjoG4QtXyZqmnLcCJY
NWQ+HzgW4s1WCrfUrM+oI7UEFtRNbvye70ssC1s33X82QYY8oI3de2ADk9c1
zKugrQFBubLq+/znAp6+/wUbQ+oEooVGsCe5UxYmdQUqZOjhZRX1ZQwB8vzn
JJC4BiLUJBVI/Mj+uAOv3bmf5FQocGKrMKieEO+Dhvpj8IPIMhjBIoYUQ4sw
2uE+92zwyNXXse2vXkS8GyjL79DxaMZT/Mnhu7HOgxiH8ykgVL1W5o6TxpDY
EPrO+8kiRD/tDkfXGDuS/Qt9Zd5qAdFxl9e71IFe9eaRqsHS/mWPxQgI1p7/
6VvOyRX8K7MteWEwA7bDjV0rSTEqkTgeaOY+rJzzTfpWC5q8/v5Dq2s/GO+c
O6ScLgxIxshUDsKg3MwERj2ghx6Po3ZI1CIcZG1Ma82pIFZSCpa+KDQDwjmF
kpNCigSa8il75rnHaSFKBmomrf0b5y5I1sGRThC7IAxCvc0AkQCVxReBuwsH
CeP8i5Bj8qvWhWiq7Wwc4tJJcLhtXPA2QP/FDgRLlg/6mX5cueDnsWd/zRPR
DiJVvDvqPO2gTTtZBiCn/JLCAxzuQbLs2lTwT/UGr8qTGar4Ov5eTY6A7FQ8
h+hveHGmSKhVCCEc8GGcYU8ncgawzRm6a5Hfd9QG1E1CUJG/vtfPpkORKjW5
w1wvXk2ck/ZxtpQuLUxI6/36UH8WBGuPap75f+6UyhtHbHvXRTpwo+eSFK6V
gMaK4jMgd84R7PkirJoxyrZCh/jN8/sCj6/qgRmcXf8YBemNh6UMqzHxqEDK
FiJrcfRra+kZMs/6akpHx6gjnUF56kr3yWgX9SUsyfsRDE3T1cheEOTc015B
73l8RkXgooEtaxB/WZGJNcutSuR1MoZD5QsAReSCHfoatTkGwYJqf6n8o2aE
6Uk1NyvlSL1ZAvH7ZL3KKcL5rdtN1J3144u5wVauQHAehm92Coc6AMonVzhF
INTufjcdFsob/NxFZwkRfSMBMgBdLdVJRVotqt8+/zsi/3eV1+ZR4LwIg5uU
bwjzXyizeKJfheiS9hGIW2TXJE2ARQleMaCQZNY/+n7xNnP+0wc4Hv8vpiv3
WogaFHpZ5tq3/HvKcKFEZWjxe78ce7KDHk7ftfDnD1GgeHtjfrzjOCZFzUEe
OhbR+0UZijuHsQ8r91IyOcUpxRl4ZO9OwsXpqA470QsMFub1TIPZKhRwCzKV
bi37RHc/xiUk9t7ZKEEv4zLyOZxaoyLfd2ZIYhs9eQ9T5tetWkKWP1tk5HdU
kQYX9dS95FDs7eaXi5bE9FPmvww/18bHY0dLdw4lHxiBSm7+IPpFgAtRssbN
18G1JVrEB9b4q4lcfv57mHq0/iKtu7t6ex0HrB/8rTu1b8eC3CgSbX576uPw
Q5F59vHPPImPvWn4pgWiAOJRGTbGgcueg3Ja81sUxg5wHUIxddaZu5CXeXIx
CSkFp9cLoKvp1WMHvSwSnpwA3RR5PBnuvXruqwD8FdLX8aG0FAA7R4MMobNw
vvEi3EsVv/2bBllrwl0PWLDVu7H7vEi4qunGlNH5uUZEfXInYPARCFmHNjXD
5jS7154YsLS0BfexytHg2Rv7Vl4Dn880FjS4Hb9zgoPlslOTuODKVROFhNFK
OPQmG/TJdr/iZicVYv5wpacnJaEkIwA741oorZwP9hhsrmr+pwfArebFThDM
kpXKNuGBkNNSgPc8eKAe+ZVP/zAnLwuMC62W2yldNFJ89B8YklJ8C39mmTM2
MhaP1P2yxr+VnrOEAtLhaao9g/F9eiAa5RQ7QWFt2/mT3DRiCKjTxkwQcxDR
nJCXB56I1FCQeS0sr8kI56ZtbD9yCtwbbHgDlHlG6ApVqpwAgDUNV7hhxjDv
++yXVMZCkUen5CW2u1KUCpgRn/klG5Zv+QxCcWtkKcN8qpcvbks6Kx08YhsF
WigiV6aLNpfBqldQdhO0XDkV8F3kFHPWi7Uvkb93XVnNnRmCkvKpoPImZnFA
JgAt97BFrreHcCN4x3+AAnKQy5wL/CB78KndbA6l6Tx38LeUblqAePQEmX7Q
6IaPZEQ6w66K7x3w0BdVVbmJ1KTjpEpIApOEZWUKksMWWWFmWLB5xt4kJIYu
mOPxMlTc8K86E9Gci8PXOOBcs9itnOG5IrroZo1sXBhZerpjvzM+22cD/Adj
Hw8DZ35Pz9ReHeC0zMTI2y5kKCndGdd1H+U1BHjV2kJQaTUmeSczWATLElsm
WD7kqPKBVqi1qMKbBHauZMKOl2GP5vIyFG3Q2bJvW65pJof2FYy1u1ue2X5D
D5TMPOXKroytN4HXwdM6r2HQ74cYVNRlYZ1Y2xwf0u9DRVn9TkkkKR/uroVg
1s164xb7bP4nHgSNL0mbvKwL0lY20zEVJ/yyQkDmWoFDUGKmrAr5z4umamq0
7zc+nPGwaOvJOWPpB+YrN2fUVGrvXgmtuSUNuQN0DZyckck83J+cA+X5E6z2
B0izkeHjqa+6utn849JFNIs9HRo5+5HXRAAvrSLTvX+xpXSIdykAa/QyICgy
YYik8WnoomA0NsULfsaHVdRyaHSJCJ1NRwcZccqUSCb4CaPLc4GoiPuDVhpv
NcRbdrcsY1bN/NRlijOBheGzrfB4oddUjn2rzBgRqyTDVmrY3yrQ2VJ2HfU9
mqF/YV3u+tqcZ3C/KHfjatlixt9t+yKq4mRzEVDZHR6lz4tVEu0sh9C77NCN
67JfxBgUQJj3hQq2kp5s8K6Rk4FO+xgPUJuvMcDvRpmc0pDcCOvak41wRpjX
fapxPfPduvA155fRcWLfwun8mo4a7l+2DfbWUfWBFaRe4JE6RUdV3jN/PrRa
Mm6R5Zz5iC6sQXLVJilrVtLkvDa/y37Lp5ktgd/Cf4qrhJO2ILYx2klW3O2w
pFdFDsg1Diw/G6Vt1zOOCGKyJH76RuUz2cC9O9uCLDxTvbobGhSY/Db8d59e
qWc+v2F/LLpZA2EGy7wUvhpwhIS7idOSMaHPnCTEiPe9xWHrc6X6/A7aqajj
RFzr/0q6uw/XsHE2swsXiS49S/GHXew8A5EAMvONqzWl8X7R6GC5cR8mPOkx
WJSIKaPUF6N6vQQeIV/L+nmAWtE5MwB/5ReQv0TsSbaUl5U5IrvVU+Y3190u
kjiou5eoqewEqP6YZ/4AmkA1pXV/AIxdbSUyfxIq+4TQkq1hf6rqEp/0sNBJ
nPeikkMO90vM8sGQ0md4BH2lgU1YmAu2cb7qpMHmpGEWS1/NGh9MGzy/vJB1
f/RtzyeKCndkcjV/xr+ynKfGJ4uSbkTSUyomhUN855V0CJWIa1AdTCRIRX/v
sYqayV0E9GZsHuX3+tV/2qaBUx8A9nGktiBwFqKVCNtztjG31b0/FxtWL/Rp
pMLbKsHwnajzuQpepb2ldhCHmMM3W9CMyi4SMh/46SK3rHtNvXUWKNEwhtvq
lAUhzXYhm0dhMQ4r1o1ZQFvK7OT28zCpG6zZSSgvGSTB2GYZ+8z3EDctL0MF
2Sr5kETAUVmzvv9PPd0mgH2XHRiECgI/5cIRmtBbU6sCrQkLjgoV7nXI2jxc
LfYCTUahsAtXGr7HGnbRqcikdWmVo5JGWc/RDlRijuQdbpdBHjDFvDPUm0T/
npAcnUXWk7haQgdKGxjl9NoWzli7To5b994D5Mx8aATmv3JOjVVMAXcmK+LE
SrSQP6D7OW45iHImf/l+cYrhTAjnzSh15/ztbqZA9c+cWy/GVHzi3NKzr8SZ
kLmA80GDf/+9iqOtLbt86G7JOF202IDIdBLD7fiAm6yeNXXkx0DSCyHlvLro
2pBe9ZM1c6Gd+uLJdR3LaceWZWzaXzkdpcpmlXae155vtx4Bxg5xzPitGV8O
v4DHiTb02XeXiLxCdafWnPJEYqbkY66kfzW+jf3kzqJvDayd87vn/+9Vw+NR
iVNE5tczAyrqcBs1E4tBcnjnMn9ETy+Cl6dvS7E00YZdH1JQSlSfnd3H5EX/
fDUhmIwLYiSMPdE7k4W5yddnwrV0JbSx9CUkCtDO+YhCa7AhSeQDVXN6Cq+6
KtzY/Q0W/1j0RLHR7GWKHMop+Q1vWTR37aJlUsQ1hSvIQwv/JuAFHiIA4epU
omMzq1NnTCqc7UaAlBxWZJ4fr7yYwi62ResMKiLFKwiQD4uBgCHijGx96UEf
df+O7Tun6meK2vI976DYeqvInaokXYR929SIHGDUnhgSrTNHYAag+gW1Dn8E
NfrGK4ApL3EJgSKBGAWBYmw3MZyiogrAhSAOOwlCypOCu9P+mP7pARccfezH
yky/Jb5BtM2o/6KaVxJNHi6s+nZe73HIcikUqCg+B9KCGFs1q2V6MYp208Tb
2R34fZlXkCoWPXnPvzTlA+Pdu3XIUyOHH/CycyEJH/wZZH32XDE0IQLBujrj
tm33ngfHtjFE2v2NXH2HT3etoQOw6QWuAlF+m/rvlwWco3aFIHkjgyf2MBwE
7MklQ8gKZq80lFscn7lVoZqE0Z9qztt/H8ORywTb6B1XPYKSpe2Vgr9X48pm
QWRDCGiwsmln8JH8pFfFLybLYRAaXUf/EG/GiIVHJQBCsT8Sn1CengWdrCNi
Js8Xu/t4bqmTHuwlMgiEfBLqdN9Eh/5Mcw1B6yYocoR9+jRMeLE14DtW6/ui
H13bbTI17PJeGZ1JjGZHQpH8GLFUslE9+73U4RLCzdBGyu5zULLbrgpA/SF0
//DenQZycaoGQR0q4BUCIs3mS9bPDb3LCpaWflg/1rJhYRUWzHl4YmMhrckb
RFeENKh710B910gMlA4BeCAOjFTIOO4jYboFfeRyg7c8+jw0F4DcA7aTl3Jy
IarvmzPudvEZCDKaWnGmlEKBtJIXI3jFB5GaZHxavLUZDk3Nafyi5Sp5Jlew
Xb8P28rPTJt8/0IABpoATzn2eFWu7+BrRsc9ufQTilIRnDlGlv4Y/WdfOy/6
lSfMR97/KdPLobtcaYHIiVbw50pSSnKHX8asCpeYNuUIQt6ZWvikSse3d3W6
9GF0D4ptGBKIX37XJ8uuNeVF3lAartHPh8QB0/pkBMmVQfZuxElSs3mMjaHh
cdQdoDrYnYOCzOL0TTnGXDw47wSoQM9jtWxfpEQ2B1aRpQY3M+fkZgoh+TCI
Obvq4m++ARk4i7x8jZE/EWY7nngv9yjaW9fHOAdivlWS8FHg6/oBTbmkgnqg
UPcrO2KaPcf/tzRqW8W9EDrSKzU8iSMzzLJLgvfaoWPGdRO80wg+U5Vl0FBI
VAuBwws/20zP3sWOH5MSpVTfbf4w++SVFwtnfoFVhnmEEQEI8pCoV2bTYthS
8a0b7kJDbOr1qpVb1xuKUHw2M1FpEKnjy4o1yD276of0EaBkDi5Fnz+DJDRa
v2DDnqU13CrlPxdpNlqft6IuIdtLJTE1shMgwFa7R5kTPC/7sZa5iYcVQXb2
8xezVaFIbu0TBEbwf3D8R5ARQcFDhTIf+mBIVvvI7+atpuHT3kneWxdOLt09
nUd2rt3zPmvZRPpzlaEhzpIMOV9XslI3Q31I/qmvdNRi3DyPKISZKhdM2tb0
ppOByPTz/hjbEMKX+NtRmEvv2vkZTILSsOg/0UvhieW/R/ky/SEn8OQ5/EHj
h71My4aGZBHbOVJ6jpp8iqJvFwvfJ2xqLXwLurZ1FuqaryJHseiUeLQR12KC
QoJ/DGU9LPbPCxLdPPYdWO9487Vp2MJjA45ECZ9dXXGSEgYLFHB5HdbtDWPz
DGDCLUtb1gporEBzlYZshj4//1RnVD1mspU7n0v6ialK8ECa4GnN6GqmsT3I
B15MxPDF7khHRMW/BA9Pd9370Md4E//LjoaDcF76oDr/EDIdhjMJQLE50zuc
VL6Sx7t+RFehKfPTJse9thS/qwb7g5pggz8FQo9SXkAQrx970uL8eq6RiTAJ
bfPWiD5ro6mXhobSVa9cefQjIWbU8IzFGt1lpHhI0Yr/RmX0cRYccwl383AS
CDXEfOZemeON7zuqxGoipaFs1nELucu7b2OWSAl8QubdlrAbSe2C0V+Rvgdk
W/O+ap79TcNj4Y0Y2wQIbGm98RQk+78ngcGjkfwhE1hx7pbzfnBAisgkC6cA
L+geQ48Y1/xV489W7CVVWXQ9gRUrLSzMxzWcVITKnuX/2pqwrs8WIMVXgiUk
njZmR1FlL5R22XaRe4n+lG2CaJA2IxSz8QdsYu9dgNU5BvV2n1LX17DcsskV
OQO1UsIkRknO3I5dBQPYZ/1rN8f/Yo3BTIL/uY8fVca/YdeZnA9387Iwx40H
ucDd/Fcc3ewn1JhJQYvZ8R5QzawKQTknRGriNJ7M6F2YwwYe01yUG4udZHQd
nJNiIc9qUbG8e43a0bijocKDNbMWmjnUuJGkQ8sp20xgtu7p84zgh+WSv3r6
Ey2K3mAB+WB8qvptJZGmihSGnOHBrFiYMWyo5RT4/OcIsuNZ2mvpDBrEw77q
0zAcP6Sa4PfNR0usALlOTfrKaGc1eOaVAQpi0Z1pbvQczobymbRz0/toKNFq
pAllLsMMsWhTxnnshGaq2wYtmoA9HYvelaT4/RJ+O3+ehjDPcbch8yQEd5YE
5FJCMk6noNG6t/w5X1U2XSr07AbAfJnU4f3FucO16q58rSFTIKT8Si0HnKXS
BltO548vnxVxDxVRGX2Acr/6DmvfYwI6tUwmy+JixKJxDPJejNOIsv3/in7F
Ze4NPXwDmVxWlXwOFvHm6MuXsJRnsmJbuhf/455PJE4IeGCf9q9yiydcjisV
37QBU2ndbiOZx55+61zS8F3ZBA6oDxxPMQ8IlE1u0op5mH0MBEnXOsc/4MiC
k5K9tssFMkExpEEOTsMp3xlC7jbvXuBK0MNJp2wZujqIo/yJvxSY6OXSVFBL
gIfZGboj0kjSNFjwYvnZeIpPh+3kqf80tsoPzm8tIJeoTY3gcKjanbte/ggY
vTJGZJK1Fl3OqdLPAudtRCAXt2pnpVv6IAvCftzcfKaRlAxuV5XWzpmOB46I
2rdbVHxfYubslz/4HYY+n2HgyI5SJ+Cnx/sUFqSXmvv7g8SI85y9BTFprN4Q
d2FTbyouTSwP7vKn///QzaW2tSFjTqQuq57zttrB9MkEsnTSwiLSl7Yobf7B
GZ46oM9AjKjmZx6fLeCb/DqHyT4jhD4IXvET85Bo/sVN286CEPhGLCZBGQ5s
mBnKRWCnqok2vxH1v1KbSrUrF0BYetg/7zgEDnXurC0Q18mCDUGPQwQBAbZL
fjdz2h68PHtPzTDKo9eStPBBl/8v/LNA+jT1hw/mwgyJXfsfYAIQ3awzlx/g
WLm5daUYXXyTMMn6gn6vSKjjpeCjBCMbwwYpC7hRhGIjF6L8euTkA9Ux3A39
QsuttG9rBfG/VtMEaNGx0uoFga98GDEwgjAThdN0T20JCOOvot72FKHlrgla
19dLZ2doR7TCz9vqz4iOeMHzVVrmwtNv/HAtJzMucpPwARXNMZUGgEnuaJiF
lCmDMDXWEtAQ0BG9UOS5mneyojgBjHX1Axut7jv392H+vOoWWMqLjTXQbMAO
59HzQiC1+u+BAXqyeJgNtjPqZaUY5Laouovw+mBr1dWKiGU/UyAe9OEaDopv
0zp7nEODlY3b0xEAurgzJBybIPl4TJ2YEL2ISfgA+yB1H11Z/WcWd4OoujbL
Y2cvknqEbbkDkwBsFvsUCz0JyKPkKhoTL8r4QEaMYKF7P55Vg15+oUDzfukr
/DPl5JxNOXYAAQ1F7gkN7l9/mr6A9BdVc9lbEqTYFzLpf4fH6AYkUDF1KI0l
48oFGAaBUIamsCkqV/4khoLdwR7xmfBLBCe/cfwjiF/lAG+2UHBnGmEh/snp
P0QRBzjD6aX4brwZqfWgc4PZrlxGVGp7qXlJZQhm8tPmqvfbjOWcRsxzHxr5
Qp04UFatLqOcECHBlWnc7s5sk1yDlVo4AFywooloUjgrBH8ONOCVkT3aXUTs
aRSHS8CothdCzf4rluvdYRNiQr2Y/rmDhsYDYsAtm6yEwpFNs5rZx1p/AA0K
+6pdS/WFZ7JMeiBBSlvhDgPkI7VA9UJlICuFUpJ041DO5bDW+rs78ASnyC8Y
eVlYXdlJy9t+i+X98VthV6/27ItJUPeOTAjQ2K8yd2TsXEqTPEooRFvzeCar
SXaSl26/S9OVFqJdexgNI1YmuzQnrONoGF3mbr7BixLcXwkCirIBdHZrQaoI
IJjPdyjVYUSeZMVrAai7mmWAacm0O7HzkEYuz4UvlDd7RBu4FfPF1XUNJVe1
g9BnEHcU+dikjctXiCW2EacybPZTsTwJ1nRAgHzqwTR+ZKgZUspFyP2lPnC+
vdmcdmWbTXBCgSIEd974vaGvhwPzK4tWg3k0QYlnCjTQKVC94FZUj2vGhTGx
Dof3oc3Fc/rT4kz4UkDhW1jw/F9kxrKGgrSmTL6jl3In16RBWGPb6MNK4rN6
jOKof1aQtu0X/H16RUz45X2SKs7bQg2vAuc3GHmkXM0Drv1NHwF9Q/Gaabgx
JieEeLCkf8mgmUr/7aiUTtP+EMcFFOBhXqUyoUQYimPeIuD0dhPYoT49AsAn
KipHUGa78C8MwpFUdz3lTAEz6ttjtU8EsWmzXsN5DdsT54/uVQQm4IUhH/zY
K1wFKN9XToeI+BiblM+G5sZaDBjyx+isX1E+7N2MhxhjBgXTer2x2kp9WHGk
REDyD5JtHXvX9fGY2YDgEdXPjjoWIXS3Vu3EHSsqAdcsUeXFCblhYxU0Eocf
eGK0m3l/ogy4I4/ykzzIbnMEYicfCueEuCYh835fwtl7dUhp17DL00/l0pdR
nglkAGMm+dflDMXscG9Q5QqX5u7F5qe9fZqW1Z49eyRu1beI3Q63etOL773p
8BCwPRXi7ZrRflEKg+F4UZceyBgVh2fslPX0+gR4NdkVOzFQrEzdbxRx5mWj
yJ9xoTkkhZmHTXVUl6Omea3a6DVGTaeP8aRCRrmaTXdch6vrtqcDyIlAdGM+
qKvNpKG/cZxJQQWUhYIjrsKADxBf+UUZiDMheA9a7mZqWeKL9v5PQW7+W2o1
33Z3IJG+Dib4WiD5Z/a2Rj1B6ATcrR2qCboR/eYO0xa31IqqrqyRQJjNT/q1
DkiafaIosbF5UEP2x60sUQyswRyZkZ8ZWmnZZOGmwZ6XWEY/WOlFPugMZdzg
DdG9G1hwlF/KJepRPFGN8g4sQ4TG1CnI5v3VBnR9RC3FdHMe2IGmkgJUrgTY
RryLnxEcZoaQYqoKpLe5l3fnVvFlT3oe24bADuGu+Zlr4B333bFQPiYKrEMR
EFup9T7vgRT32rrwihcdP4R+WalT+l1reuj+3ITO2uxWF9xYpY8xuCQDKZ6t
FevtDM3wF+0SkvolHYhA9oqpirk8s6p6arREThfbXFY9cBN1tgQiYGix8eSv
WVw3xy734uSuytOYZWRPY7zzCqgJgoXZx6Oboymd1b6TO404X5lYvPpC4nam
nYsp9bWRL/bkzQ61wwcR2NA08s2iZLtMFRwh/EdqpohX7xDtAzHhzqOT5BGd
1/C/vDroBpuKLYHQHOB0lbUwzWPkiiagbYEPM3LZ5RUPQGsrGDaaUgm694Kw
hv6YCUjek5q8KvQYIykC0lm88PQVOf9kFH442FSEBiF/bB/eq8bOgN00nINi
ew4KdKIRuLZS7CH/QOOetWqOUwD8nvdrSIBY7aaQN1EyRZ2GtGIfGO8UO9sI
z3qh7LiKUPpTSivhMrN/je0AuNFt2yllAq/COJ497xa3Ms21E6yUChhFNIZZ
Uggtvrd2OX67OBVG8+gb6nvIZ3LPMtUM1HEs957XUik6a1ywUsutVuOHRf5E
8zr+GO9D/fS4aWmnDWEM7+3tUqt3Qqa2OgszrrHtn1UMJ0sBLs95iVKZqixG
Oe3CF5Ld8pyR6EPnaWVrFPV0Xkg9F8Yxl9z2CY33L909YNQbd6w9PrVzBw2a
SeVpJ4cP7ktILcGMPKIk1oeCcWumUyXkKWCHSC8acohNNkOKPcVbsopYQaD4
kBNXD3InXo2Ysnno2b3HJBNfkBBcEZR0nltVb8mXdJD2j1FFl+y9wg0UsJRB
FQ210sUlzlEkKFIcgdo6QYfnJ5s296F1B35aojY4V89XbSJyyQvXZsgeGPy2
almMqtK91hHfVYSokxMjWpG0kTchRHA3aDFBTPspdmTBgjaAdEqNHtczgkHx
RZo64NhihFtjBH0kVSU8hVOuilIvwlw+4RUHUfOya7V6ss7bkEH6AcERcYGw
DGPtLN00DyeShtjDlyAHOEmfYlQ7KKJdVjOdI6Sb3LT15Dlxes9IfufcE3ZH
hg3Ftowiin/NOwfMK4JkpPYBiqhH3vxUIOV1MVIvxlA1oV5gwIRQqoBQu0bv
Q78dZfyCgvq8pu9jMGOPZZDKhHaz5EU14YXf8+suURG8DOFuzeXnyqXn7JWs
LoWW0N0lXY2fGFcxGQUgOubUhgmqfKneQ3ZF/1RgtBaGL4MV0aHsn+sY9vdg
XuARnC3CbpcSY9pg5ZQO9I18EJNW+CQmNj/svwAdle8oC+2Pj1wDP1jNHKUe
YRe8xTLj+RysQ6n1lODuY1cOA0erxUbCZ8Bg3tzq+spHOXNEeSEaqneoHOon
EQwr1wcy/Yxj3PKhkbH54xfCxXHsG6yQJ39vhf6w1TSoLyXBaLMAPl/Al5mg
C7D9Uu0l1MbxQtSWd1z1GvdF3R8b6RNpwZ1Q8fmjKcIvKPl6teAeU/X2qVHu
ZsYZS7iKZrP4iNImLDEl5DfteklXjerNG3QPCbtBuO4m9sQI92l0wpWQ8ujd
5mA/gZf1+1awKxoKW7NBefyBUGqZaPqUDLJdIuXwnBO9Uh81nDaGSOu689D0
xAXAWY2RrC/F+61R9r9WBpVPsdGHgm5YZhVCEEoKpWvagi05O9OMUWj66R0E
JFjri32/VJY9eRuINCnTf2cmLTCYqqfBinaiBNHzHW1oJ/Ap2t/oD0jozgGQ
zDnyoQZbPlHZ/nKORjY7smC9D9/2jUyKQuNxwPCE6ZITxNlIS8facdWvtsxk
Ifc3NOJwZdVskdsfBmue632++4Cwvs3QELyzWFU8U+pWM7sF7taD0Dap/u9L
Jf5FzrPJzy/Oz4iN2OoH5lhSEZGf5umm09OzEk1rmzRp1wym6jmABQj8aFel
niEpWBoyshXmADdAwyFZFolmdMrl03uRWN9H8GKfT24cEig/6aaREB0+1bzg
rWZFtIANSL+/66euBYhbexkKBDpMjlMENRArl8YhphYy4RXpGhWjjKyy3DLA
06aBqwCWJfoLMNUVdTs+3TEiDadIE7li6Mspz+NFfv/U57b+LC2E0g9XlQEK
pus6h6V3bfGObs0UKu5SDfLaiu1Z3tZT4aSBrx5rvn9Wdv57I93ZHpCPD6kb
zaR6TUjPcUwaDbOUN4cTk2bG2v5jbfZ5ZUF6VcQxKQ3Kuh4XADawo6Zc7VbT
yF6P1KRcGF0UdAyk5wWNu1hV/LCcpSug4aUvWNkXkNBsmdnUbMBcAMfFn3yd
iKZZgc6TiWZvv2khQ2MNunTnm5p2XqPtATeHyBb7klkPyK+PuI/qPXVKVJG9
d37NBaCnnK4Mf4vL6HVuiDVcQql1ppgqw76QndBGLM3hE4bYfDpPitVgyfwv
4xOYnRM+SlnYDDtl5FCXG2xQ3PP6PQJc6Pm8WXvp6lkd6fvxztiGItqly5w7
P57LdVr6JMys2SvVDceyWavrGpaawj08+j+WFBJFJPIRs2tvaNGobtUuwOQ3
rv6jPGxftV0j3znbLDZ6BgsqkiFxvqVIrp9VQNWQJ3m/oW3b7r9Ik3wPVf9F
OXzhurJ6o2j+C8e6z5CUJIPrLi/oZ5fCxAAlmN+j/ZKgLZNqsGDfSGzVUsdJ
CJuZHL3RY4W2NPPXpWrmOlDzmeMgIr25Hc22PCMofgPBzHAn2OZgVP0Gd3UW
uSjo+NFRU3bXwcIaLbyXnK56T58Lpch8x9GA0CQmiTsEfn7TC6vleRyh85HT
WIkUDFeYfwAkmSs+1BHCBVne0Nx6K0LhZSWzejSN2X1pkgpy111BAt3fuR3g
ZhVOIviehV+FUrGcVJB+tARYVYIdKOR8KxLMAe0MFq/mQHKjvb8NgZdGoyPR
MTqL5XLMUH22R2MYlYSQF6ZwJCmhRswP5ZsQDYZB2QYSvpF0NU1bAZ+7uvga
FYUQD0fihMGu89tNVJkb2O8j+2/9X4ksPbEBi8h2YqbGLtc6tbsZQ7CkEL0n
HbcKNeR06RqhJX82RnfWrNCtjUDWa4Hx9Aum59X9nz1XH/nJDq+3MyicnA7G
y5GunTVfI3qh4fTzHCFBDEjryjA993cdMNNMBPDTZkejo5WVYdRmOcAl1fr8
VQ1ySqBYV3BLEkUs9rgac4vYXNrmIo95gfsnUo0qEBr/zVWgnyn7MPG+ACfE
iBhz9gV6lLzkmLRux7yO4lfqgzXP4Zoztl9Ap3pvnMOjaKkILxA7cFQGD9aD
5ic/B+mcUP/ydqPVtUJ7DHpnv/OGOHur4osmS4zQa/Kqkgfc/H5M8qcSYIin
YEN4BA7+AyXiqwjN0gdTsMjs3BYIEjD+PGcikASZikMPvY4yZSI2ujHbQDHJ
77I2h6UnTcjuqz/0l0Fv9HFZGf1kAH1c7KB8U/gBwQx7Qh9jAcivNYHqyvzm
yqdqISYhSnnRJJvNlTSBTME1OaEfUtbkEmtEBjW4MuvoDEySK+RyVXmyJO2S
Si+ndZmEHVqe+NpnaDfF74F47DMW7WrH25KQUuD8LF6GL26ecAJv88uyX93u
3DugyOiAJyqf9TnzvxBf57jippzWkZHg4VKnhfixgNzclrCZDX5xVsgOqfqF
pQbH+uu+qKT9M3Oh5vLV+J+F8B6phyenMcNorqaMUtbm/iV7s0V3VLjc+EhB
sjRlLHANaR42rdQAvaDf1OEtdYkpfchHBOBfIHxfes3I/L3JtfIA0zVjw08e
IDrt8wllcA+PM5CQifedMSljA1yE0zflwcVNvFiMN0RPHvi2gxwhgdTY1uAv
phGiVMw+JYKUL1BINFIeWYhKBDvxO/6kUM3LbN0Lv0BAON3fhFU+ZmDkprjy
8u2Oln6JNYQ0x7TRjnI8Z3+ZiO3Wa0qRXA5bWSUFlyt5U/5Z9konfJartgtg
4eFs29+T+bf7mlS9Dz+kUzuIMq/fRPhWDjJ47kGcmIuY97m1x5WaeHEQ8px3
uumaCCWI8/qsglORC7oTqfTPCcfRoZxtvSmBiTLlFHi2Rph0K2K1jEGpXM2R
PmDzd4gWhZksYctNkMBth7SDTgEUTl1eNaoY/jfBXt+mz0D6PiToTEO8VNpm
jm6R6v/SjGIB/Lz1yQxa7FP7jnMwkCqzfQx4oaeLcemgT5RKaNhENnRdNkTJ
LWiHLZMp293Wjk9FAfm/dwCZ3/dbWlGSx5b4fg17YAqhBKVmgxuc0Dne2gpd
igPAZVlJKJJSVbM+a3lcsEjTqGz1kQFSCxzrNTE9OzSRB7pKbdLSeTl4IPMU
xUJPTj0iy7OQ/YxecFnZyW9EOJr45J8Mihdv/A3vTvKLRxhAdRRDvcywcTbF
nRJVvzrDcQ9ukgOZaspbukTgGZDimjqZnAmH8y2BJsZWlurOfdVMPi37vZJl
axYAQ5eUM5q0GZuHbm7IS8pE1TM43mI8zvoUgNeyXImtK0CNrUdIj9tNvAf+
+PrITeB+zQnhtghFYqCcKxyD7MpmffjT7bN8nb231JatYlvYxr/I9R8bVvys
GqpkbwUMe/ZmaMFjO9aTk2O8xtWDxX/JTbhbPltWj6R/7D6oOoEOwAIVbaAk
lJBZH36g/vx4z+vd9u+fgkeD00cyQlZagh9jW8prGKJwg7DSJpMycxdSQBu2
6cYvmgyi1txy9X5NUyN7bcUGCxWllDkwjtx6StyaMKbLI4i4J9j8LaH5uM98
aQ6nTH94UQ0wPyVpOxUgVPpR6I2QIYe/j7urnqWgDrv+GcXi0fZVJI0Bd40f
p7VaoPr7TgeroQqZq6CcM5BLt8A92YMBEiVnFLh6sNdXUql9UXUvZrlxNV9a
0JA9rgXUr+yTjF7lmi/wYOY/5bkOb/AlYwn5RVhQuJ62jMEZbC/3gjb7crtJ
A0kFuliia3EIz4zcj5+qJVnyHfhyWobk0j9AdQoqk06+8+E5h3ntNKvoHCb7
8OOYxYd/M6tLsuK3EKp1aQYbPSDowWYQ+Khq11u6pCjCqSz17WQ6XAzLuV9U
bANpkO/c1jK4AFhdGbRLBNNUJbxP6zdz/p1cudIQw/6ZQmycityOUJmo2ezn
nBY+qB2HggcggMuFB1AVcQDomkTP2eLrrNKC+5przSxPiSXt9KwB8z73w7Uj
bRD4ZhK6FSDtybk37MM0gWxwYMhT5hZZ+unimdbySWqqhw1RBQJVhkwD9Zde
W0A7c8ZTHi5Vzg+N7NA/oeIf+7VifQt6CgKdm3Hsw8r6RotBBaI/7pnfZfwF
KxsMZjcKMDACjEXqu5hWs2MUBwSByk2Cp5Uazc8tKwqJgPOH6DFD/uFy7Ubq
nd+ieJy07Mfpzf/X0O6ra2bAq2GDFbBhFYFQYwXqr5h3LI8GqKZzOhEBIPUQ
g6Zf+5FlUou8pAfUzJLTDwHEWijFqNGuAfmlJWCPfSdFLzPgM54W33pR5rn5
52fnM+4m99o81CyBU9pF2BLsQ8xyX+jBPusphzwr210htI+kq8bE1r0ZBORK
DU2o9/VQzFuL8qTRlKcYTiU2JZu/LeUzlXNVaH0C/mJ+TSmTh5my85kjPEdJ
ue5WiK4tZRiH6MGnJ3cWkcbaQwVZQhuhnul/nETYsINPptSVV82qWqx7DtXr
Zfk5i23pIEr6hn27MDuah4kgqtV4IO2tG+kJl8PK3to8brtSMap8IB/tHz8t
uNPnCE0UNgH0L51Fv3A1BHWBN6V/3W0dBYqCnT8z+hznKsBhrXkZP4cTjcoB
R6vw73/RhsN3fnaltK2SbgxgNMLUDBiERFZm9B5TSn7WY3KNSA8MtaBLQBaq
R1dk19KyNE/KVoG9kFWlGe5VXX/mrrwKUyj+xYjE+n42YwfK84gP2a4TZYhe
N1khlh+9jFtM+MbxBo0XLRNT6JCz/JrjJBNV7aw/vdALMAQVfxNaid1W11Fx
+QOEY3nWnrYAydPW1C80P+CKhWb2HLdCO8m0VcDEKFQIQq/5x8C4xaiVrPi0
OvTWteqdeo/x6q+esF3ikMI6jhE0g8ji2L0yLkUX1q4wCf2gZ7rv4oTNijea
UeGjlRUYnwZbCXyoBG1iFDZ9P7/XFHqyHsOdsmK9nGyu42yKfwIA9+GHCscY
tdn+BrxNNkaWOZjuJPLFVetyQ5LYnxxiO1IZh/AHOqazGEJVMjTe03mD59dP
8NKj3s8LwARthDLVZlR+tdESew5kSHoSu5SFbYTFAO0Yw4PHU3QgrqVmiSdc
sI4TbJTW77gkq/mCaGluKPnMZdeLmZLGebhAbxjRTkoYeFMUGxrVLFoLdWy5
Ze/46gEP6dm1b9AyzdZth3ZuiX6k0yomfTblEItpG17sTVZubt27VkRHyAPX
KTJ2iBgkI60v2gYmQ216Drsopw69RJT8hwSwERjqvbZF91FepJEQz6G6NH8r
4R/GFORWaGwg5QcnubQHlId7xfJZbFnp1LnqzwAUDh4XYMiiuDYEC4PxCtM4
cn66v0m+b3JvFWLsbNU66G58INkzSypaQY1RdgC7oZeKn18CxxBLRJyypTzO
D3JnwbMi0uahVXD6VXQjgSjSdCk0p7W6rDZuYF5Bi/pCZGTgPiAruZfJ2Tuv
Sol9fUUpgHYIeDfDlUUoi1LeRnuxJwoGmeylHLwbNUvRiFmC/m15TR8+Nhu2
b1OqYI+yB1b5sJ0ziLsB8/wRiAPukG13RFoxsWgSOXWwO2BRoh8/eLomyff+
QMDoweItCJ8xZ9DmLyfBVf9/DBYu6QF88p4Vm0BntQ85rbGPFbEeQvUsLyp9
OgO5yMdCflzV4jYAQGyLgBro8gt+X4CFEvg8/X0tEdJS67Q0m3uArLwrz6oi
O+RJSMN0AZDKvv6YQsa07CrSVoRMpMQymXPn4MyGhqPNo1cNgcjBxfYSkj5a
sxi92RsAahdcZjt+dC5Ij7v3oBoRbv4TimfsghDjAJkY/4CdhIaNL+sRLyCY
WIiKZt6xtTp0RQJ+j15PClMQaMPICjhCYUqeu0YAphF9KZ2Y3YCjJVvsoxR8
GoG2MRpKrvg8SikI2bElj7hzNfwNrJnj08fPEgap6QuCIG2gtScdpY7tkTqO
pDVhLpQj6md/9oIJAuChwCajCCxVLVJ8WGMU0M5P6hw4JnWjONZ+orZWnr7I
uWMsNYjCHP6tpC/DqdIMq+UnH/p5RUbHeyuf3rduymOl6TIDQqS/tFAb2j/A
aBAO6pZ/KZajHUsJGknolBDnPf4nPFNOdqGtScRv28QEC4ViPa5E4WKxciHp
ebgXA3/lQWk2bmwNaEDmwS/2OmGlaB9WhOTzzVHZiqeA5MmbEqUk6VkZWXfq
DPfqnGyvDF1+Da/TnSY9diezguXmEzBMihQYGrtYxx5SuOeI46r4D3jl/Wdg
mPyVMgE/H2XonN6zMC9iewAefvFwgVSB/NeBGHeHjzre6m8C5Joex1oECmOM
SffX2lOWixzSLlT+GYrGwsjW2NkL+1v7pQPA1mREvuJb38k9GmHs0hwzH/U8
dqnAIul3bl8QOteZnDzUcB86meAdmYGUFKP+0gh6zTNGStpEiGRoviF9iC96
ZvBjLZ//wkuBtd2Jl5gjm9B+9EDqdhXiJiqAqObj5c0Etp5Xtjp9qMuoDTKH
j9rJr0CSua9tOq4J5RCmoaIaIbTwi1l/gdO7dZafNS2FNeoGnkRIpjOjgOs7
t2/nsHSDSjjxc1rXki6qb6BaDRjFonDbKxf2kFboGOFrK+uTBjxS3T589KTk
c6DJk8Sa5vGvGpr1K0fQSDGyH2PSd3Aw8wzuPxRmqT58nUNa5/nk3PJe3725
PeodF24dv3QxsEXhhm4o12nF/bkThyVM+i5eQC7ee4RjSwW2UmyiwrUVuoSG
Ae13jpZ3UoXelSa3chVQZyB5YmhOk4TIbhvijI7bBF1XdkWdJJpVVBSsyhJ8
ArIpB2NImdtNUXHaWLrVnj4JaRkkNb+0RWMb+dx2y84JLKRHqjSEWcpSKltK
IIw0hd47DgHzlAdHBTLmF/eVXaoEgQgK+nqikMzYuGFr93Rs2mPpPIMV9AXf
pYiO473BPygBWsoLUH0PJGdei3IVbFATtOfuFiEZ4AExgg/WxcNOXZYQjuPF
ItPPdcWQVY0Zc9/nMPufHMB2Jdd3uCuvV+g91T+mwfZIh4UUdxrei9uPx/N2
wAUJAkL/OqFVu+foOmKvkfyoCmv1No4knA8TrE5VQMlHvcxo51L0yLSAKuX9
RFbR9MXuacqU+z8+BwPAa6ofj8UE3UPkABjpZwxRCPZgGWrQ3rJgcjjfn2E4
fciISUL2MYxEaCcEq73TD+MYxm8UOJfTtQR6cCI33DJZcpv5Q9f+MfcZlVw6
x5qfoWp44BfFtxtkbC7SIJev+DKYI0ZyncMW+goFtMcrfbu4OKnAOpcobfln
2GTeUnyCNW2nl2sMgK54c6pyPXVThaBvsk3cJhMewErail5OknzYGmz/G5R6
k7ZqONLsxSGRr20RaPx6AohxoN9fe7MF4CNJ46FTT6u2j7evtjdvd+I7UKJI
XSHRLl07h+YBNgBDhhCKyTicgpXCAuvrxojUo5i9dk2QVKycV1WOFnwx/F9x
FzPr/jjbVT/I8PrBZwfhOeLgOtW2MoaCmi3+vnXZ1kGhYKtbUsm6Qcya0aoi
lF+FQNbX0HlY4Ewfm5tTOelF+hZe2k6rre5UMCGbpPh1Z0gfS4x19SGi85Oh
GfKRufTIPIP2qT+bxGD0KYpnXTK1StSLkiX3k7e1hVD8UBbWcW1IEE5vRJ9S
Q3L0mcDtOLM307bZswmDDQA49Feu7/Eyd/Iu/P9c85l5ZnmCyIc7CMOt6hgR
GSxoLm287T7iJPbMFYMrrrFKSqzG+/8X7xz0RScdBxtQ6CKOMlVxRK+KbMtu
lWhqmPlkTj20aRCWyMIUsigozX8Kr2PuFLjlVAleIaDd41Jc580WlPEJWx4c
w70VUkWQZU4FAZP1acB+9V5Bi3KNtOVrE5jLsK+L+uNB0uR6XgRBTbpOjRSz
U0lpluPzOSuDVOV33Ci2Bg5LbEFRA1Z1fR9iwMipEis11ohrvHvfQG5VlIjx
v3wmArP1+iUqFqPMTeXf32uX0LGF577GQBVmRFnBNwgA4P9Fpgv6aV/qDnNi
r8th5G2cJEVGWoGLfY1nY3jMC2Hu5/2n4R1zWVdbbXieog5U399G30WhniDU
T1SXtF2pl38zElDpNSuHCpEMWKTo8495xDTbjRHC88XVrjSBi/7mGlK0Gj+m
XIs3n5Il0uiEaxaxhp1jMhmGPQJjKt26eYQOTfYxiU+VrpZPu5zRs3psr8fM
IKVAKoLlZuULx1rG6sbj+js3VE2FlGsSsszRyJTWahqRKJ42sNyASsNl7gIm
yEfuW+ZOBcTBmbwhYbSwGrqBbnJ2m3wZCKrMVvIZn12ELxPgvWVcE9jonZX7
8eDE6hyQnJPR8fNvgnIE1bVIrgQ6lOqWMtZ4bazS2CltUX0hRw57vPpkcTBu
Uu6YMaOLGpuS41QxF139gw9qrPSx6Ep9wnulidxt0VhMQmLT2aHthOnTuEtq
U3iBGAHLSDukbR/s/w2DmU9Jegf0ptjyupNhOU92BeG8p6yKV5AR1CxbVjss
AXiZlqraK69KI6/3+a9kmKHbfnli0QtkUAJV673+W5Jz15H1JV/ECgpWiuNh
uOVri9tQAWfSc7WdfNtxXWySRYMK8voB4/y1nifhPcooXPgvP5KaVae1U/1X
LFzBxa0hwH71ITFu45J6uS4FFy4D9INDOFZfT/PMY8eVvKEkE0vbvAKgx5C8
9VA/WsZnwhjK+N1kyQdIRiqkXmH4EhGyYaKTzrMw6YG6IAs9fQb/UN2C6rSO
W+9AuYUAVIzlntivL5CnlzAk20iXH7UnrY30h65jvy+eWt8Z6b1MW21vl3dd
i26/icb1udbSCdnyZBWoYb1EdW53+bp1sPI2Q4RpXrzDFx/3YAgAhOIH5Bx5
qHo1c+lXa40TUbH3WpGGMXR2vRZWA33SLMba+WzJ3+uvFBky4qBEpLVxdJ3f
8dbjMeqhJfGZn3n2bKGLOu5nACa9EFjO90BLrghCpeUfAkMp8qmr8+IlmG1k
zcwa2OrzoohLmpban/1TJjwkuKlIbmYSgfYH0mLgq5coQzSUXqtrUXDJ7wi0
V6tPZ9sgWf2zUYBGkDtU3GQdDxdLOEPydO34B71WCeP0QxXZc7/hxJtMIqh7
0DXx/X0YviN25aN17MSCRX89qoYGmA0wGvBaVl5zNOqKCkON7Ut245TMoRvC
HBxwMXJjouRhi1Pr4QLAU1dTOIi+AiM2a/j4Kf9mtVKgkG7jWkb0BZzqcG0Z
URFQSZbQZJIEx4DUflOVR83nFOebBKIHu5PF1GNDtbek2AjRZLZW8UFmMthp
BHIki660KAfilPfpKtcU0XSYJc+6pvYRuart5cjPzyTCBmDljbDqH7ay6lCX
0vZZP8AtSJRKOFdSb9n6Ydaju3OPEaiQ4832DAC9yOQ3t8gkVZ+E58iBARHR
8hd2CPpyRji4TCIrKDPGhkk3FZgJTMt+87MsXpGzF9iCDJBlyYfgHcBNvQgs
KxpLe/Znr/TeVf3MbwnsZpf6FsEOj+FRwS9tx0iJuf6L5ldB5fEStZr34CEk
4pbX3d1D9OQME/PcX9YDrxF5Fua2WDoIlIpFH+sWRe/+Xw0qG/BHGtkD3Q4H
IVXW2Oh3rVqY9ZZcMNIV2g8kU0XDfZwVSvtpJKEcGcZp33ymSBMHQ3lx7BXR
5kBT7l2stOKLR0gnpotUwAe2nDuzDHBE1hZmEm8mJ158FIAbCSWQbsEy5BVq
8vVpHCPNrg6UQ9kppFhnt6PJD5QMJQ186khGW1/WUj43yHy8FUNIwJq1rTig
sCpLNWiccpaFoRJpcq1+Eim/fUfLVW1Tds81SDlaVKAEDenlWIuEZ89mZBFS
f8+qg4eFaqjzotPzkh6oi1zklSqkxVkIlSAXcFTKv7Cj+4Wi5DMF7EaYAIXs
gMeHJfG6U/1fn21bC8NW+2MQ+M0XRniNmZImGiTVWTG6JdSbXC9tOUem0yKW
qxlByDK6WPgKcgqIRDhzlACE0uunxMzV/YmiXUJjAbDMGTP/Ri1GmPv0HFUy
n4uA3lmQ/E+e0tyY8gPGoYdAstTrMtF5qTcXWO4NVM6HOvba0hOxMVwlouns
YE8rFfn/Mu0XPu6elzcRtDWZTGZhuvBSzCbSdTiQOtpkiNtO+OdDpfsPaxl0
s7oe1pP2jdpO6DI1ewwXxWoRRUm6fmKuHDoLYeBvdYZgOKfQAFgXW4x9D+N8
OJHFE5GUQnhG3n03OOG0QGhenIvDVN9bbza6peMbaDu39FSFjzqkxCbYch0g
839F3jPrAW9xlVm2sf2yTJw0ArOiX1KORwan7BbUpDojDFR286li1Lk8rhlh
gD2VReHmFEESsCZkQ7D1R7cwyq5wzTJXQvSXibblcRqSZCSyWmt+FTLRTCfK
ODpfrBEKsE9+MCNQ1rFYc5G40vFLxh3HerES8hli9g1Dfh3NtmjhQZo4+gIP
Ui0Ua5wJ80UJfL77C9HleZOAnA480mYbTOu3TlcidASeljfoVAgiKs9RJrVX
XfGSJRc4WwpVQ5Y7vRcy1UiCwLENlZ6iYFZP/Gipl8Zu+V0XSFV6Vr6xHeRO
MRLGawbRgpY7WNJ1jllYx7cC9N6wrKvqTF2Bhb8sNN668EFW1lEoHT6xrGE9
hYos19J3mhWNCuw49exh8PCLZSU3d012hjbCh2fA9LZudQ14QtUQ+HFwiLvH
ssluzqYbOlvhrbiuujoM2l6SMnEIVioZvzWyb0RqTyvT6lGHR98hpf0Qu5RV
RfiKc2JR4GTu0ZSoFK2ckjw14VTMPRoL4HOguvrVt9S+oIP37pPSeL3zGNll
65JV4ZT7Op9fEZLztdHSz1Z1ZD4138Ozw/AWeOHTTAwBeyFza0iKDhzUw0Kv
PfndTjNnBebmNUfS7M5se2r8+5EzZaH/Ow2ta3l2xykbAGVEXRL3gJy55x42
pqLs8T/VGyRXUdiadhEx+K1FA2iVCBXa0KmeA8q8VCVyBpkQ8pc06Ah7qql+
Etu51e1yl+j8W2Z0Iu1GSnQ99ptZICrSEucTuZWUnPa7CIG2jJAdEx2XB603
vbMvEu6h9gDb4pI4jikLRfA5wjghE/vK2VqgvfFoYIM6pSwJWQnccM00Ovm5
VbrREsA2ExKtarDjtWA7p8Xh72l8fjF1atA9zqnrdtktdXwEvEvBzBDrR141
7Hb70/08WrtRoXtSI2DRLGdzlgXxL283IrXP4zA6IV3ke3/cGQKkwH6quh9Q
AohEmpmqoDEfH1NMhrTgn1TGfSH4zEdCuIj753SN44b1e2qqpYm8G1N7GG3A
jPqpAmmx17vBt4PP+x01piUMNBYkPZdbxbvOA431DCOqh/B2Brjdr8dl6Iwr
slJCC9DVf/mifkhzB0wZaBCPKncMNXfkczEuXTOuZYALRUO4zJgO+t+Z+TjR
0dw4CdsvABb2Colq2x6yXd72fh/wnSgZtsrjkhv0uKeoiiqlgZUluUR6vHfR
5WSStE1SDPNPhtNMorCQtYE/7jexUkjrF0Fza8RQhAhuRPaI6JPfQ9xPQQu3
KGIB5wJTNkj+w5gK7oO2HHCVVneO30oxffMAWt0NfamuLPvkJ0iSS+voJG4e
ifvn46mcpKDP0E33i11Lc1ZDyQun98TH1GI6JhqtvEY17LUhhnM0tTZHbR8k
mS505jTa0sFHNCBj5wfOiM51UP/AlNuyyuoeffEZOhhoz0+WG+OV0pOOCgVt
2ivxyIVFCYkfqS87+QjkZrDVYK5r9J1BUcA8kp3Y0GRwWViO2ZwoR3biMVgd
MOpXNDbv20GKqWOkPj5QOOhIkNNA2gGHjT9S4kWpgWeve0TQxqg3VOzHuQOc
TnTATK0gnYqP7gLJD25kYugxmwcy9Ny5k2bz6yzbNu3JVSYjp+Bi5T4ZT9rX
KHm81hBvj0ZOCgUrebVa1sko1Lqxg8mpdFiH+RmyAXh6wygSXbwB5AW8PXHH
+OE/dUWv0F+yhp6hY2s8A6Ha6OjzJN15O9KWeH39yOYuucxHDI1R89EnUGuU
inhjpkAiHLz5gXzIZhmpa+bXO8tlt5Iuka/awFiF/Rge4X+sUn3gUwSffN5X
IlxBvRboGwH/aeS7ICkNAODZpJURbqsjmDBwVy0SCBOR5+/BcWBYMg6+tYqm
cqZK2xqasdHh8mnUGUgRlvR0jIlxPS2d6ri9oHS/Fdc+HKA/yItV5+UfRUgX
ufGIXtxqTEngQsiBpbAUF0cxnYN7AiiNLzCnIbWEF+FTa9mmFyBM8sbboRlG
q8Z3QKpxUKKoOlXRUDHNB7PnycgLsLNdhX4V73fDh3MF26B5J1ZSfxa7MiXn
WH9YX6JYr0Wl03chjurPnCjCohC4BRvQCHofFQf8YulX3Oz+fthkdrt9cxup
p0g3IsTxxFB3isQPjYDC5QaOn7AMPJ3QjY9Hbtp/XDmgZHoEJ1GrpZR6Bb+b
5RncvYXuQR2rXyVRsuWVk34AKN6X3+PfTui1QOd2xw46XiBNpebFB9aXDj2N
jboB23kvptXiiKuuQprlL8LGmhVUjGBlal+y1awPJ1HEOa9G2f7ANXJJ+UTG
OyINUcp1Eh1ta5t8sySrUyivHkdRidLW2tGZUfBILcO5UdbJYUi2dHLyQAtD
EQOBtFeQqQJ0E0godlJ/LCCUwxaERqYNsmL9EI8SntXz8WwAC5dDC1N9E7E6
1bCdj7TcaAX6Eye9FWvT3F4sEa77tT3BYQi8j1E2idcjS6jZqorafly7Lmlb
sOaxecycUEtgMDOv08v/ifDT7TcFVvn928pEbbX+Pbk0knQCuLV0KmEvSo8V
PR76ZNqTQIEIi3WMtJpjG2bsdzckedunQPs1Yc7YaFp0jhq33VATYkGUP1JK
+G04c9XmI/3E1x5ZxNJ9N3mgS9RMlWSwg3zheuY79RLQiL8M4LysaaRmSWqY
XDsNVc0uELEB2xv5nUp3Q4YiLNr58cVPvzedzviqZMWUtsajXLDEp3i2vxOA
UtsnucdUCYupEEaqgcDsnFKMpze0IftVyvYQZQw1MTUIxLrXCoqiHuyvgQLo
FxXUi4NVo//VdPwHSRaGaQrCEBed+Z1plRgQtQO6CWeWll0AcavWQNoWjOZH
5pQuPM2Ria945C69yBiQ+KeavgSiYKWC7mzbt/kozNBhmiM4MueCE0ayQBEc
yaKj6voDMG/YbL/lZyjtK0O1bPEuX1gy7EWIFwvg3E0WGb68im8XUa44ujMx
xMfrptVAcdRwT9jHMrdbtMlqAw0y2HGLRbWQMCeFZMEPAph9/u4O92Penshh
G1PEBtHmOQKVB9n+/GMFjLj+sCGAjrZYm/br+lbq4WnbMlGIGCpHsm52jQIX
/l6N2ioM1DrHI1pKn+QWeXQkPCFLuuo2/HoCjk2fIYO5N6aW2zBM+rSOyxoH
9LeQdQVL+k3jjcDJiZpqwDu173/dcXP6ReezuUa5A4cnvV5FCEyIWWZoyesd
wf1gi92HPBQ4ofYeMWf7t9f26hWpHjFPnwSJ1RLH1HHAJwT10mvkQAEkIhGH
s86q7Y/Mg7LTvNWa/0kgu0I+fPpg5y/waVyReq9IUd1aVWeKxTuFgBzrLSCI
lQfbKYpYirxaZZZvbPrzxRBZtqoWA8ippiuS+PbQeFUyC/019vHfW9d0sxD3
thFUCF5Lcw4GDiprxCYjXJiSFVETeRdFiSqj+ibBddeFnuppoQ9yfJVxVBNh
87NvJSTFzO5DUXmo2xCnGwSkSyzoCo5E2u/42eEjXeQm1Dt3cyEhBLnoQ5cy
7DrFRkSxPB+r7p10IC2adxdkbnkajW1Es3V8/qlnu5EjKRWcHdxtSvarCLSk
2rAL0Iq1OND4YPFZgTV9TeBz5UaYNuynaS8qrR+kMn3v9eimBvHJhfcrJjly
ixIKSxBjwsSYE9ts0l8c010tt7iQRI1H2WZKzmxIITXmvVqnuKW0hr0RteVi
mAGEKQt55PNsGZmQSswH1qtYk+uhi5AxrVufFnB7iIXpd6hj5Ud49h/iLd0Q
xuadt7FuJ17264x/jztMhVxBYkR31pBWwAIdbrP8MLmc918B/X0SHNmw/thf
LIw4Jl2CV81OpDOCe8Gt5VKi1hoa1OTD7pBD66hL0tSo9ArgbaqeLB+A7usA
66Ji9tvRmARcp1yhLKzbHgEMLqTVdF8uB0q54vaIqaWBm/MJBlSJHSfHGmKb
3PzMn0qrIuwLmHv6FOpVAG1XDe8hXmuCCVT8bFw+rNqXN1p4DB/1u4GZ3POi
iRXrcPgcplPINXeRtf9R+NeZO7Nw9yW857JinoVCL8MSKLdQYbeqfaDDZyUR
nFl/QZEh8I2B21P/EprYXF/zdyxblBp8IIGXkuS143jSe9TNY2sjdsAAHE5z
aCUkKSfMTQo77PgSgXTtTIaWAmnhHYcwyi99bBgY9tb73uQlE48lMUNiAkWF
QNOv4XLECxWt9+uaTzrjfKoeI5absqcReeCEQFWiD8uRpPHVCO3bUsKoOS6/
PpHFwQih0V7TW06KqRvzodwQCGsLeDnsId1KVstKUXn4AOt9zrcFIJjP4xjh
6u8nMx8wb6SPlKhUMK6eIJ/IuTtCjGSrJtS+d7TOa0uVvRVyukfkWMU3Rs7w
pgzLWLqFN2CBr3tTfRhARWSdmeCzrOgwD7F7OC+xipBhJgjMOqTKXo7ZDiQ1
AveKOUn/dgqBZWLH9nqicy3A0X5qsYR7mwAowv2jbTzZO/E1oJzW8xO3A0wS
uYh2NuIkiB4k4bQDrUF1lnmU+GpNJn4nTIcgtRnYMA0MiYi6k6OrzDj8kQGu
ZkZodBZJPGAJiPvlsfDf5suin+bjcgPm7gzOySdL0S31ZrxPOJl6l75QyQsJ
lThHTn5CLSHVmUM2i1GcruDadL3LuyTayIPoFxdoVxUsgnXY50ITqwvIHKlx
qjOByMJNaV6Y0UdNNDKEIw2g2HjuB0vY+Jrsz+AZ4dWHxKLcKPKIv+EfiyCV
IrroFeXBJfhp90aBiK+PQaBiIGjWSSlrsfpq8MJiridBmNfpmXAIkrWljXnb
oM9S/w9k6T4JTWiZfQpNOBA1CGxgwmEwno10xXcNRnReriPCnaryQ8LvQ8vn
+Cd6U0vPV1xHJKu4T89iqOmOuTTdXo8mV0OovQfKF7WYToNoLSJnU35y3wpz
guS2jBv2xagOJblskIhIZsmhKJlWWCXT42V5dN/93eKRFCz8ZMbrXJvQED3u
q/sC49YIYdEZJsrM72DNrdTKyyLTTVzmPVxdSLSN1Adt0wySi4NP2F2LPLHa
EHwSqD9kNPS1H4YdAIGcawEn84IliUs49z8n9JZrga1hxQ81ofY9yT9+VNM2
tbXqkSFT9wUd8x/ORinMhPHBi4m+YQEABMrVbxrlok7peqRAgKcRYmAx6i2P
anyDQo2k24DX+x3vSX2P4xb+juqeqlkfxgSyfjG53Hm92d6HcbZB+SacMMOD
6KLciiVolHVVjIZ+4mv3kEjnZOU8yhO8MLUy2dHg1/m8AzurkDYe3PRM/ddb
EhWkwDFBKh4JjX+jPXdsBE+DX9ig61pbHwYn2CUziS/9vpxYqVgkjgy9Cqzi
6sTPxdMScio0N00b8linXO53sr9ZwFWuOuWVzrnJ0V+zSq8i8ziDWhIvVlHn
A88WjtMxdesp5/g2JPmzta3ZvGrtI9TQ9m9G69CRUD563zkBIIJMUTvQrK10
Biyf60Os7e6VbcksA734/PB07Z2qLz/6tNnrAixzg1rz8SynLzKBLNfeA63p
6VYqC+1b8UT2HmrwQNwpu1lcisXDrJ7owyH8XdK3NU/RMYszwUNFfVNOP/GI
B8sXc8oZUfxN36RrssYKDJxadyA1+QoXo+8TFjk3mr/hb4pYY+tuc4g3Iukx
JoF01ndo3VpdPrtelKGzBJuzWasL9ULSZMRGADy+S9Tgy0uuoMYxIMFORdjd
8yzBUXVGU+EnOGgTBjbblqJcSWyAZUuJ5agx20nVGCAAjJY3GQ0fzVnZg89v
TDhpd3j7ZHQ8yIKWmCeZa7K+7fuPLFATRrFKA/Lbge/mWIyWHcqKLGLJGXLp
fL/vTU2raWXCLEoTF8Y3krybzyYw0wHo+YUU3+NdiX4akgTRzNCfA2YLqiMV
//I0yjLnpX7sEIXFkU7IsmEuwWv3FfB1R93JD1+4+y1zvxrFjMdxavLdSu5S
sjhcWLY1bOTu3Gx7npaxbf+61XMeVHo4juo9dhslseLgNIYDRQgkzJ3/cA2v
xci95V1NubYv5F4UhIzg3dBPZLjmBU1lw90xCtqtAL1qCVOPzJb6bAtl+16K
x+GOY+mTWOVIZFgmbmnBdxCM4vE1wIHhL6WYotzVB4j/+jlhEYspz049gWFp
uoVU6PsoDPtFOY4ufi3NRq4976ZBkD4KJJnBrVHqQvJtI0X+iqH59sgBiItM
sromghIdvft+yWGVblkTUY890QVWOFCbCuKGs5sXSROgvorEUcZGDkxQEBTp
1LZQ8p38tvAhWIZ+mvBjt2dyE2u+1W4QssQBPEL3A1IO5H2mR7VjBc4t9dfr
dtRkebngBI5OY83E3yh7XfbJSsONsNrMkMes0wMkTjTcAi6A1NwYvxbvTACn
Wq7bjiHkUbAclxX+Ua5CZeRJO1r0mkgoz+7CnnlliUBSIO3Th2kD7EjzrpkV
3RpVg6w+CAQfTZHuu7Gt/nd6PfzPubfVr0Vl5//XA+7V9ZCF59IT4D+oqmKU
aZOFYfEt75eWNWxPkErqb4uEz5j9ISJidsnb2ikCjH+fs6iTaDAzu2iduOHC
oGHVBQ16pepX9fDqgKzQ9OsCgHwXV0+DZx3vaU2UPJ4/eSzefK/2GTr/EEVc
e82cED/vTxe0e3LtiZBSUo4jWenc5m/cUk2xMtSvfqRrSByQWjBhy0q/Bs23
rLvOcWwvonsOh3cbPGcjj7eQqXhlWZC02lt/xWI6KajR6ZY41WwuU0vc7La7
YorVM5EA9jZLEt8ACFgPadJSGnfFQZa791HGrI5kg2DQv4EtxP49CvBo1MUE
poroeIz3OOKxo3i+0jhAi+ao2YXiQsJYqhUhXVSn48GyqvwFoh6sfY1qRTMB
f0Xwe5WMW5R8yKYbX1qkGvU01YvZR/Fc8X28FOUdTLmDDk4grggLUBgA/y0y
jwY3NI+TqdPwrtIhgdeLSYSZkya15X5pz0JbMvfDW12QHqDj9TFvyY+ZaLMB
drPf94aPMSbkRLFQBQI+/4iJTy4JJORccOHrmVy7ov95McVIPYwkp2DDadXB
o3/BFPlRAUHsItVW/muq+SPOz1TEI+3XhPg7UczC85PABFO21l25juKVtrsb
2XRAF8rm9bRI7rvhYrn53M0QISTGMhW/C1T34EL/NyijxtVZbN4LA7DPmkCE
u7ag8i+P8AJttIzNUxS0RfTQOPpOp/CnbPfVYG47blmULbfpa1ps9Xyth/Jh
ISJ+SovAhh3UQj4vvmDN0BHmoQB0PVqBhC15B1Wap7WhGyV3ugzr20iMkNVq
IjiLghBV0PLZassJh9SJX8gnF6NyENtIfhwRQ2CkvuKU+xu3NaQnxpot8QRY
jkO8wYrbazJuv/sKRd6lpcnyPWZLB+r+79ia6+3qk4EplkHxVQFebLcr99vl
U03CBTOGaB8wtvxkkbh7n15Vp3Ur2u+wfnX9rEQrfNqvNNmYSuHsoXfzRXad
vSI15kCl3t268q+wnGORdHllXfaA8xxAz7vabwqwJYLIBwmy42sH52DMh3BZ
/ZQh5sCAiN7MqHjhk0PWuw0vSzNUxtfAaZrD30uav5SVe4YbUXGRY3NxaEPE
mAHqElNJ2dCisRymsooqtZ6yuIqXX+1s0QHvXWiqiBZgCUxWkH7nwkgINotQ
LKjh40zK+ut/UXoCJUOgf5VToS4FFxMQq0id0Nj0+X3dG4xbDPD8iZwW0ICi
Owp7NbEyf1AJVYXGXGZr03PREJrsbOn/zmTeAQmUmqXSTJjY4pYEcL8MIxpv
u2Z8ChxNt+svQmCGeAkskwDZYm4uEaqlv+yL9lsVWxhvyFIuVu6TmaPH9wiN
ung8BYSmd226TN1hyoDdH6xBlaswYlMOhB8KVS0dsQuXpw1a/gcY0gQeYxJI
C/N1CzTCd1OhrdW4Jj3DppbhFbYTeAW0Wb91wQyEO03KWpp3w8rW6mrTlpZC
5el/naOrmQdtb1IEbMVQ2ZHO64zmjU43Eeu5iTnhUyTm/L6skLh3RWT71DpY
l/e6ej06vIhodVnziM1x92sgFL2Cst21SJ8PNj2Qr/YWqnhUyh2q5wBNHVPw
VL31hkBYQB5FOjZcYi6gczEhu/beDEFABHmX9CO/PqMDl0/vZPPOnvPc2cbN
cJ0v44h00vfiYN0DO6hguWnEpN3/+vjizQwB1I77TAuGJMaxT/ZY3Stv1hc9
DtBfwYpopV8cuOpFKkMdjZwSdZwQoN5sTD9XnHYBMiDcgHusvh14VFqxVHsj
vKHoW3Q+OC3/ZacY12MG7YBncDQV0Bo4d+d89MF/KFhtdMlWfJkxd7JRmjzC
CYD0ymd0YqK/6kE2Pd7W30hCpBIpDnX0jurnae2yFqLIVguIukqGEv+a1oPd
p+P+dH/fepJ+pfbeur0gp3UG3C1gKgETereophkEW/ZlNKWxrxngXAezE7bw
NuBElG5CbPU2Sgc3UfrgFih6yvaFqEwRzqrkfpUTx5m+1NX5JXysjtYkQxm6
5EPCb94qepwuIMsWRhvkdK7eNB1zqN2BWKq3xK+anL+gCQZUVHkvX73GnbgE
hlo0TIeuHHdUk9n3l1uN93y6L5z7qIqoUOzjbXeQE+doQzlOBbXUjTeqhyVn
wbPQGp85kCr2+bdKVTyzVOzr7QS1nGfiAtmJQKXLiedgem8NvlZWMwEp8+Y/
PYtID8qilZfk+Hp+HwLpcJjT4dvV7fp7BUCkEHqbE9zfkJy+2oQe8D4HWe6c
cQGroBu8aI/vaAERGyEBUhJQ7Jqs8X0Qj+jT8F/QJVqwVQH8GJHaXl+9GZSE
+w62DUEVO3Eqi24A17ViEVkQH8XSoK52rFvLgDLqHLF5BoqMWhrv52NVxUPH
4CIFImsHL8rodTGI56/jjow0HGOlOHoehx3jWDOJTtGkChQl2xY1IqDoNm/H
2DjWaYqoKGHmcUuW5KVBP89h7Y6D7PgE4Qd/P4xJ/uCfZARBptAvTmBMX4Ms
lQ8c56lobTEhDVFgMNXVcAgku+NtbyVd79p5harSHMen7+wa/+82IJHzjGV2
xth1EOPKVHnLOhDKXn1jhVr8x72q5b+R/on1asBhdK+6YyLR3T0cs8Tms1we
G20vi5RsGWGmcoEnaFLsuYDE2KL6h/bXnjN30xxxjLYfbwsscYOl7LxuPkZn
r1MrCaBQis2PAlyX8vGEjs5GN8otItNO7ihkaqdaY8Kw7i6Drn6g3Pr/DOEB
meDTaxSj1yNBuh9jBrXR2fRqUjUZWpVqhYjfam45778jJWCISy5msQDQglqx
ODU7tYC6wUwrE/OwYY2AP5LT1/3y6k6fcAdFtcWWoU0ZX6TyLoBN8iYdRYa3
Kt43u9LpeBC9QrudOkv5RDblU98NYNIf6f8561Dp8f3pxTfZpCAz/4eLbfyx
MGjGqYinrFmZ7F/Kp4SI39/cfrXHHAVNDjQMNgfQDCOxUjo/1UtylnC0OEtf
La8xA2cwqX/4o1OSPoXIb3FlFnx05d3jV1ismV2T1LZMQq52wlvYZTGMoVFL
yKBVFTHZlsDlnGqMI2ac4VaZhC9mmkerc59FjdEPr4zYebHF6ZP+1XF3uqv8
gWJ2jPzWeCcYDsrzBeWhjd2g/s7SjLMdd9ob0QWRUkgLRuLAyahxm1DugUOi
+ouW/wX1caL3pcRRIyZ9UAjF3znZKxfVUfjNV6s8R156xLj8AvOzvGrrlS/b
eyjY8gCu0bfTeGVSbfoRPRBbzGH+6zB+z2XI45jIyuWoU8uRb4IvKHN2rYgQ
KLRvQYvzbawbbe779xx6/VfbRb7CqH7Nb8vNtEZyEDmftLI3RBgXdrVDOd1V
ulycxFRFfdEJQ+zLue9AXVuzx3NTqXlijvod+LIA2MxnhoJ+zU8cX1ca5vN0
ZDzYXH5lDj2YBzTRNpWdx0SOQBSKH5LabrfLiqHlGzst3/YaHjbWeOpV/yek
eEnsWClKIXaa0/oAjXMsxfVrrV7TWGWCPeeQKsYwAs6YBuOyMXBIyT0hCweP
YeuqFNR99BuXDKpeXZKe19WhMyNJqlJLRXv8m5Xxz2CN5Cf02LgeSKPSLIU/
P+dAeTeu5imTqXZahmYk5k/MMwOVH49yMJMmWwtfQhdW1aX+RUj8j8Fn95KC
Q8EgptzIaJmB92I0nVU7NfYkeABcpv+lhYVfnztX78cF7UsGnSkvj47ohxTa
/LtZ+WNlfNDYpSJcz0R00pcjThgMH5MB4H80wxCPEWpxVPqbV+Hx0WWk8i1V
dagshZWH/YWmnaZ8AH2ZpnznojuHBLztjSQ1pgTS2J9smXkDevyxsgSqza0q
jlrj3TI1xHcSOkJJ/pBbL5qdATJMZFzIB3DewzwMS3S1Y0/LIkcFuiCvTdJU
GhFCMQzMGmp2aKGJo6ALDG85lhah+uUJDFBGJhB8FOp7Gax43eyAUhEHsFcU
4PdjtFxmZghTNRq0NVWVQSCafJTaatIDXzx53+EMXFpQhl4CCv0z6D1Q4Ss5
xmbJy/4QLLLaALzBNlHQy8Stg79l0/aCN7E9YLMtjRWLsye4+n/uHWHyLjYn
6rsn7oeYaNKvZebX5G7muamGUC/k+iX4O08sr6bGqCtuF/lp135M7I8zGZ3E
h0Nsl/qJvvSpQ/w/xELyOgj8RfyeK0KacgfayDUvf0kkeEHo3mrM7L9jEm+q
PBZos/U+G9lMRFUKay/GYyHLvYr4w/M0jK0lqmwaxbcNHcwuVdHptX+e9pA4
twCeV5BFUC03aUjMyX20y00HFEQh+6Ua4/+pcdwSubVi8G1t6HkWusUbvQxU
k0lBmWCxWJpZX0XjGxNL1vsNA+V8XrOAT+SbFpjGZGSEIaxgjkse8fBNT0sA
71U9eMUbrnlPapoyd6ubfnlTeFJO/jZLksaKFL6mNiZb47HJjZw1YAv6bg0q
m8aRUiXpVptqIOplexdy00gB4QfeRQUxCEkxKZATeNl8QlZk5cKPIdPOW8LT
5xlLQ4zAxeazkXJmAMpDiYWHLkmINMWzMFv1ycE6Ng5l8XiF3Owsh+GkhG9m
BeCXG5JUAESpyDEUo3+QX8ogGKwlaze7GKvTf8wgvcN06GV59Fqx7nvVrrnH
GUDgfYeemlPFDCZ/JMjuc9CS5nCqdn2hQm4r6FzRqBUpKWrMfDmWD7ukg3Qw
DcLsMAkr1BXeiax8B7xjAqNVbT6/cw+BCI7rVH/cSBlSH8Qg9nPPEaeUzlyo
Yw3eneH5JDdRWn0UWZS7CyaUUlsYce+SQZbGPwNB8u0fMsaSDYm5eLfhfmyG
cNXTcgq4jjhp7gLuNeL0ZB35OZx2jYTweJ6i+Z952gNUpaNNPQrXaWitb/vI
Dv0iV1LdWYaigblUg5FjI29T81X7biBO404etajPNPwUu9rjW9/IUVGwdB+L
QEVTso8k3d2Z1keg3PdrgHOn84iK2KD2cPLClbRhQl6YK9TQkz3/IP4dLZGP
vgV+LXGnCDp+8mCtz20iJzu0amG4IEUIaF5bC7931PIp4aLoGaypc8S1ZwFF
9p7YXF0yswgsA2R5QBrRKNprIGlKzB4v5xBB6V6ooWb6L5E0hWa0aT9UBGpN
L1DBe4br66yzrWHLgMFz2x9UL8SUT+HFHpB1YsZBpmcEWAsIH3IDR4ljvXVa
c+m9AoO2iNr2/d6RylrdgaeLH74Y0o/zApG+otZECrVYlCqbuYfB7oCo4hhe
b1q/R2LXrKcy5rmDYQ4P/R+0cA4SlUyKfxmmpD7neYY0x8X+9tgvNc1PZw7b
5uQLO2VfyLuB3jZtRaZcX+MAdeO/rA66kE3iK8UZi70xy0IKRqjL9i8mc8vn
LKp3hQ41+HYiio4az35zVlvcqNS3dF7Pq+gUDZTNW+t00alZhKGPVzw5iAGk
xhh79pIisK0T5LfTYlwLbyEtTALINRQ9nPxAI9rR97EvWnuCp+grCy3h3/Jy
sUlH4xfM7+3VkHQIjKj5CTk63xJUhJ5UPeJ4MOuRxftD6RBBF9W1RtRDzXSm
bVLnMrm/vjuaxptfxmyORPRJ2QCovEM5aLvLW7evWWTRtNVzQLhwdCg5UmW0
ujiQBQLBTnss+JxJhrJyE3ztFbG7Es4z74xKu1mAUWDCw2Uq+nh44QUIq20k
ayZwZkRAZ2K/6EJdLsqizcWwe0AlOv1Rz5KgiYzVM94LwISrHRXEENPPqxnD
WX6FKN8woAQYnfGrooHc6+LhbqEa1IxNHXu9xKic+e4IIWSVSIUFGwKBACuH
sf3LeVYz9c7vROaGWN+k6ZdNVYoBcplYdD6i7RtFlok1iegpzVAnaBm5qqgg
C2ZiC8fFHhQKfy9lxKY8MD4ZSWhvA5W2NGUeYnVd+ZkUY8gP9eBYlS2ZeU6Q
AVzy4yOK2ckXq3ZQ4+iN33ZZlsLeiLLDY0tjv6+KbtOE2hXd5cK8Jor98+7H
kMz18FwEh5jZZusGhJ4L8bJpAu35xIPZE0+1C0InTKDgpEAJBYJcc7+7vdy4
bTTCFLQ4FuyZIl2oYmjx98FYovS2Pk0V/XqMkznTf/Mtzrv0SmWlmiUDphFB
S2yG/UjMOhL89b8TBxE/msBYIy8QVdDQQoYtKhImjjj7GyNZRf4vy5IejLC2
7nTBK3+fcHKoQ82YC99LMTmtgq4IHHIWYzvgSLXda4gqy/Bp/Gx7L9j5HF6q
OJE6Gw+HleFLe4zFULziGxGJshnrgiWN9WyX3dVpCX1fOQUQc1JKkB0cp+hq
liCY9Q5h8PNkQIzkbk2l+NenpEA5y7QXt44XEHWD39zHxsQ3B1RNFjIftoC2
usxfSI1gcouwnoGrGWybadVGnPbiX4xTEY28bpyf/iYNtdOv3ErLUEaRb7bi
xYzlAKCAD3shl07bKHcM3E5W26Nu5xi4TwiOuwaxHEX0PIC6qElOWC2SGGQ9
QCes7Vo51PYdOECTfADq34dm8vbcK5JhOxP60JKCDU8MwXK+i0CfWTiI10QN
09P4wXmM+4ZtwFYzaMm5sMXRIgliRaJUwqkuizg4G5oEA2U9saqYD/7+2ibn
nWTMgMDuum08yU9/CEKTwsNzj5wMHee1ouBoLgPRI90FU8O4sKgeTJBtrpJN
jTHfl+udgi5BrV0Bup+juECFIHGr7DSyolmvSIXIdmHaUeyBj3sMXgFlOOcE
tofsMVgj3s0jqTL1YcEOAK656GsdtS17wKqTnIFyeU0HpgFlw3FfkTcruAgm
D83K4+dnT1bhXWkdhml0Z6cvCZhJu80FYSJ8lXR3CV1rGlaolRxflMxSnQ25
tV22s5qTsUct58ca4gr+Uw1AICmTMc7ML4n5Axmn6s0OTlB8epDeoWgn2CDy
bo91RzHLzvTWK4iuOKkmAN6Ceb4MR8A3n9zuEtbe8OXXfAAD27oLHzAqy+4Y
OuUCAcYwjqfEZEOVpIsnOlmvhGHTG2M1thgLpNs8+Htb3uLY7STCAa7EQQa3
SzFK7vF4i4ehJgUEt5ShP5C9GARng5sihs09ObulQERMHAv0XyDpZ3KOvw1f
0uGDUhtUj//GDkZhaY0TBhQqYTppboOq1HADViF/awdQZRUbJfLS7/3nD0HG
gE84UxzKXJ5dYoEpnF/XdB5RoR5ai5fQyGHGfWsiJIc1q+vWcbS959dlyUS1
NX1WBFIr3gPUuGgjEApMUVobFw3SfoUI+d/u6Q5W4MoMCPenncV0xGcbzZw8
P1No73E8OmGmq6rQtYHWEtpzYVkoYhw7wwOgbZG0sC4dmwKpoHoHk5wMv76n
JoDEK8rkBKEP8t7a5FMYu/WyWZDGnkfol7W+KqrbewYhM8vb4XPH2Ca1s6jA
YvuB+lIJ2xEq2lTl2qac50eYvdLK/yT2pS1gux0IGVRnTIXC6yIsr7CG4l/U
OI5+cx7qEQeMfhBw85LU0gJbk1ATPGiu2R6aOuPytvCYzrmdDGAs48hZ64Q+
3GZNS5JHE2f2aytg6MXPtBkdBuj7Jn8PvmyenL65JFoVIexuRggvG2CgrU8v
syE5zfwkfChJZkmV2IOlQkVrc5hP+t9d8k9saakFdcViAtvypy05gQUGMp05
iyNd0Bn53rccr7vcJX9fJaga4xOYKoTX3ECXqZ/41uV77o/YoRy0sHdSSU3f
nqcbOP7xPKPEDh81ghXenZHBK2raiNKyI6ZZ7SsFKkN08IB5Kqblc08lOL7s
NNO/+H0LnOcclrIu8u+Ut4YbEBSqQwT/n0KuRpAmucBpx4+etj+WH+lUQUh8
6DEZMkDHYwyYJP9qMaiTdQmOWZDhaEeLMPiCRuUkrWu+zPpc8CeM5c6EGQFy
L26WU+9qXVd+i5xRLUUDmqDN9r2hhvFo7WPCJ4scGdO4nPqxL/bfHE31SHNd
vEEinfQXWTiifiFV03sFb7DJHiJLlizuK3Oe7xreBLyl5XEMjwB/U6KgT40m
sjbdPySSYLJBVgvUKAcgKeEgsk3LPq5lQ13xuCL+mP1DLOAosIQ5UIa0IEi8
H4ER9OfTmoUSTuIX+HbQEDbA1dfq+VlXYHQ25/Mx7ZPbyQV0pc9BFKAktIen
hgRRE7bRsxTx6kZQAc25G1RGQcZHVGsBXASr/MS2zu09eHX2pUctOXHqefel
aXFdQHv+79HbQU1bIBs8FrSVDK7t6r4/S8K9JeNVVEiemTbtLu2XZvPLROsn
oXfedeo1Qywk99ZdEacqkv+JE3v5B9nUmi0zqXZ/oJEHAyRlljjzDkhPdrba
JJRybYvQnJ99Z/BrX86wqHBTQDE+uMHxuDo4XiVSbA87z650fnKmpIXul031
zEZ4iWPHOFQ3k6gozlkMNpEuhiuLMoNinXpQ5RY5QiubiG69yv99K1Wpw7aF
omwx9eUYvH8rlmTgOwzNYy+zcVylbOwfcraSvHMcf3zjAbBOOBmGwLbNF9U8
UzuNJEGQLZqur2aY+zbW7Z8TJvUyXYjrS4TVkgmHy8Gqm6guGSlvIcLKVC7q
V9MbhE6DFfEWu2GLxioag5FZUpto9ErP+Udh/a3w4b1zSPMTUAqMMqFzWuDU
gaaxRaVlfLWIC1cFQzJLrr3FB6dKgmkXwKweCwW1fzVIbEqF5wjJo8J4cu1/
7rw5c47JGS4FPXXxuLCaRmnpKcaFiffBrqL085MWOyfUNZ4WO1f/oely3Wld
/+qE0EcmgZ0/M8AtCUWhhGNNPr8YgEahPgFVvsDEzei9ZgWiOUM7fxOUj2+s
xVQ2B6CYVYnfkSF/A6hXN5JhQyMjEyynJjWsRXbN0yw4ApvA/myurBrrolY6
IHtJoFyqT6gtMF79358SDVlc8A87LAlDUgVZwoOemomT5VkXu2Pgi/kyZfK5
bCnZKu2F0Pd7/8c1yW5190CjfAjgFGBYdFWOwuKehRbOitYTZjWwrnPVPAdA
GhfhyTXpvmZ+kAuHnC+9lGXMQhEOy5nj/YGY2X1jK9rCXrmEwbIjFJBSJqse
aQq4Kdr7E8pmjvXyfMP7rl4KT0KoSVWLv4i2jHQNIi9BNCmKvkc2kfB6NKD9
12xnf5cb37IvCwNinlalIyCiqE6DQPG14Pr7ERr+aQGaQjXGDEikIpN+y+3N
s2F0alacIV1TQ6FPDZgCpaVByMu8vjC0DyryEYUmsRkFoh5RswtScvKKAi7y
s7Ri/BI5WPta22aYGahESytWMcoCOEL/YjSWbWZqhNp2R22BxyUHwEcKKm4G
6s1x1KtRGdx9Q3aX8ORa7kXd+wxfoTQM8TOioN0qtIqyF+uBTtbnQOGiEifn
NzBXnuH7jlWoLacIrLFa4QSHsdaunOcy9Xtb2bFGbbVDwysNqe2/3n+jTlk6
rzm1S4oHM1jKI8xRe0p9uE/xwlro5lvOdLbMp6adn+Agyt6AxR6n8spOIgQ+
HOa7aKx4+TZ2I/KjdJGeg1t6CnA6yV1jDX8zOPvhQwr1a4+8rzcwpyT/0xzo
7sOLvK0TId9XBuU/7ltvQ40JSWjZG5M1ylUTlKNcDoglBGbsSWB0lUQUzwsj
DSk8ZNkx/pVRNHJJpn+GStdz+2PudaOYqYngZEAp7JJdC2XYQijLxAoHVOkk
1fH5HK/lZoLQPwSEYOGhUPKxNMm/aqRpkMpo+Nvo0ZjT+psSzMLGyFUm+NnP
N0DA6Wq0gaZ/4/t1yl509PNtTKp2Yj5pq5Fa+m64hIPXfKNNeU/WePKDvjsJ
0+GcgrfuurlBNsS8bvYNMKLaAzGfeuor/2bclABrtfNY1MTWvRz2GWIsWIZq
iA8lFTAsysD06Bhm69ruVOco95F/Ao/S8/mBBAdSzKfoq/IKJRRqOE2bOn1R
VrqUaNKjMTeyVsIjKXHtUS8VkkKaZiGZOwSMoPbkN5BoNd0d2XH1m4eeZ4KA
EeaNZ7uarfj7sbZlSVZJMe1TzLXEZUT6w5lqQFzTxt6Iiu4ALk8aREjeR3ce
ZCNNvy/8QY1OxmHWVexFjmLG3o5EQVoyt2H3Vcp4jgYssUFvFyEuAaqgpYu7
JvXoESJRy2p4w+hUtRmVe9HUppidbjm6tHd/qp7wxO2io9PjkDPUXXfgeRBD
R8P+ZnlguC0nCWo+GeW1vdZu9GvwcMSSsp55+qBnznR4nfDRtzHn09pHRoSv
GhMe8cazsKMeLtkRFW2cM7693gWMK1DNkG+1/HeFKwKDtbUFfhRYDpyu+2V5
nmgFrBZntXf3MZUlznwPTlKC4LFxnvZ/94I551w0q/JqjZ0KYvC0Td67zg42
ruUBuEyBOs6Pya1fXh4Koo5mhbK8nE3Q5XdqbN66dFsjobckfGh2ka/mC2zm
lYtUmnNYWKawlYxR5rjulfbWjGmZxCCVVstGF/46jQ7WevqtHDm2CwVWNM8o
L5w+qpgIxjJCiW9U0tvbEc3g3RznuCP7oC+MOHBR9z8GuCGtUpexh4x4Iqh4
0fwUOfay3sLoHVpn43/VPzpQ5VdI4U64IL25+9iSZlZP+q9+DXiqf1Hku56I
b8MpbNfddrka9BULr5Cmx7h356gBxUtcFl6lkUTvFhDoG5+Zchsm7Sg2zJC+
bfN6A0PQXkarb1gBU5Zf3c76LHddmskyXV8wFx+C5urWnaXB4mGMOnWYLHNi
lk11YF3vn0+En+6qO7m30ZaV2Ke8SLOnQ8jgaAGtxoJSjhPq6H2R6zZarWOh
PVA5H7iKqJ30kKq13grszz4FozeAuylayJ5KOmS/hdxItDXPf/LbTObOmG6q
Jcrk+zTqE6mqHHbsOXS+deEm4ldaWZLaPehuEryQiqlkdDx8AYuqg5F/46+C
eC3BQslhWM06B+sMbqX3GCcbCtMMflF4H0SzPH2xRJ8Qlre/M4KV8vW3xsJK
Cynx7vul5SD61ctx8A65ocmGhZ+toBmQXfltCT9PovAX0kAv+2hFtz3m0EuB
B6Y0z2O6e0jbIzhuRp+eJQKPNQx5d9tzw24MDRvAY1cvVLWKdHQ0gUJtt7vl
R589/Goti48AYz35N2u7rXcf4xZkyQnuQ9D254D51Lr2YIbF5fbnLwjh3VjP
5MqUyz4PRk4WIecskCTMdydAp2UlJGRKYzjwypIxNBB8hM6yMtSGHVs0Stq+
qKnVfjJ2uzOa89AyFe8iBfCE41NuNdnJo+89QRHZqGBP5sdIHq0l3B9/waFH
6PlpNwkyBeuG9JOCmU33TAdYGEH8d49h/EQbA2mBVHWCIghBZKAnWl5s69gr
vji1wQ/y3GeNvgc1wmjLitVHedbddDOcOigkt4kJqeOV93sQYS7BDRDzhNFV
q4BhRJaIxSleVIJMaY/CItb2AjwxT+WtRDcPVrz7edJixhU6HN7PqveZWqFE
K0JczEmsUgKnAi6XAzSaHSqXwsoB/iXUDO/Nqrh9c4C6qGNqhhtHI2fyGhxB
/bUs3Z/EVsRyVrYPC2DlMHsXOHC6PBeaaN0rWIRGAgTEMF11of33Ofb32sLT
FRmiC+Bq2kdSLmXfBbbLZGm15qJopYTVi3T/4MuruVnKndGTcPBpd1qVKjQ/
nbb1kxFuNXGPgIhHyVpwilet211J1nt50C3yLch52I7I1+waF2R8mRzU/3eI
oRTdmYivD0+VV24vn+ohoiKdc+w/b+zHd+vxny0lw4opQmBmdErZzX2UCKD6
ySDmCCU5nKOonIoOTwz5t46FDpS39lKrpsenZmrfHWDX61URsfliETP7S1qt
ULoCjW+dLNHZQP1jMgMrl4DDe/XbInUapfyIP2fARsTNwrb6cXi2eEEt2J0d
rARAm4zrhz4aIEn4VvWfuJfzp9PJxMB3ywNGeAWGEGBm7gATuy7aVSJtEp4Y
9cuV54y4SVcdNOkK6cVUwCq3BczLGwb8D68B4KI6eKDT/C2BNsmCJJ3g9PEW
0i0dFjVl2yxOqQZzDlDJySB+zMjP63wvrHTFFqlddvqIFzi7jcS6st9rJWwP
Z+XCCTCySMk8hU6EQNbdLEjlu2hgzaQZN9FFA2VKu8VxtZiTDHAEgR82+xf0
MeXhcZFL/+BgC8aXnrckDfdW2jgusEbOZ3JWlcSRg4JS3fUeMKMlanYLrSh5
wcW14NTTpk1/b6Cx5iHz7c158xcutTAuFZlB2LrDeQIofTBG7QehAJKcOTWA
fvKpc3Bi3/aDehDMjWYi4gHs6TT6ywxcBXZ9XSRtX4NOkp3vXuKhjC1QLi78
OjFSjKJjU3r8BDeu+ylIkt6bNNnv8rTHQHOqgaReF2m3FyZeYzYQI0o7KLs+
qH2VsZ+QgMjwOCg27aVlspJXqNTMDhl3g2zVykOCRl4ujTbEajhLHY0dS4FL
yF5pv7J5dJxjaFxEBy6PuYMkn2r/ZxfYo2Aw5qC9VWO/fzcFTUQrIge68kxB
oAmHYJSmL1kfvGUwA1cZoEWTHn/1TRZ8LsvLpMnsyz24KjunwiY0rTWybKUg
6Qb8+z8NK6e2kCpRZu0qBfVEXVNEewpKdjQIO7912qxGWSadgW0QdO42SXVk
CY4WZ3bwxTaD9QEmgaiI9xvux5zkZNJHO6oj/8KbsaKLi5s3sV8U282RfTHx
X70B3i5YRtEUMF9YThxr2KRDJcOZ0tiID3PA7cah/L0ADIqj+KaFaLvwsNf4
QjcutTQkacqf7JvFZDzl4bfRxDT2yBAgU7NGfMMqZIA3/V+3CDcBD7YpI81L
H4SezZKUrQ00qyUbVSC3r1CZmR6bEX4Ues1zW1PVJ6Io5Wb6eOPmA76qW+qa
t5uI+jq2uchsBH/8HCMybaae/M+bQNf+5vc7yL+jAq28HsQDle1QE/ml3yQW
w92V+DXYGwq7LKmVaChYTPbuxFeByJYTU+iysvNEBN/7nwydfON+LJCbYGdl
ziL9Th6uLZQaU+IjKQ92lK7xoqj/JbkSLBCPBpHjy8HS513HFTkOOenYUOQb
JM7FKU2L1U590TeVGqxkTBDDnK2LEStCgsjU20doDyocoBBPSELfhYCKo5pQ
miAzTo0zl8xACdzDB7b9rsLGgz/pivvWD7h/5KayKagM/32Q5ZilQzyr6io5
dIIR3ROdge180RGq5Wdaq0jr/As4uCfcg9zZyuFnR1AyKVQSyZIqRWp0ydiT
hh0AFc+MEV/pzlUSuDrzccV3H7XxggVCJw7MU0ORi/uA4OdlXMETbEeYl//F
ypKx/EGMS7qf2X7XvHW16MVUBN+5cvKWThhM61UDFcwliwg35HBeS56O1Sw5
WwZh/o24406O8A0sqp1eTlrZqGFq86dVl4cLgmbRufiNpzA63vsk3rmMRXUn
wYfAC4NcDpbyLGiJS+y5hxzag4zZrOrExFRvd9ZTqKEPq+t8GuKKyAGdGXSV
CV+Xqq91hajleYNc8+fPLIX/1XWoYTpYOMW+WId19jlyy0rFkhCR/lxyb0g2
nRW+NE6J5Aji1BC7CUCD6z79o0RYehaFVi/6P5Oo6p3EfrXGj1GzRlkjXtok
rEhBJgtOjhkGGyzbWAEv+tr6R/JbLFNSiywBCfgIHJAFTEXjt8LEnJToxAx/
9PdCKHKCc8yOH9kBptJaJAi+kChVGF9v8Zaz11YeoPfa788QVW2F4g1JUP/M
epnoVH299BXNKIrPL3lrnmxJX9wSCDUfrEwsjfU89F4L1vV7CeEcFrm72FAV
u4X7J4qTOooUhxWQkWGjGqp4/UJg+NGC+IQdlwyl7QijVrjBLuydQNRUxdYH
R8ZmEwHa31wW1K1o+jOBASM/K/QJuATuD36lSq6vitNdMpVy8q8pbT8szcgi
0uTB/bnniDLH5oPHknZAIK0HVKICVXq4Urw2M7p5J/OQ5HPrMxDjbuWR03k+
MJuHpizQyDiqPY9IO2JXh6z0U9xrJRREsk78ou1MfQ2fhLSJKcuKgDMUakkf
qBw8g5m8vopkCRLhdaXyL4n82ZnfQ0WbHN/TD6i2TRY+PjliaM6FWoaoG3V7
yVVNHaUCGOScptx4BTlL6T+Qu+eGXnhS7BtalRyROd72DR6P8I7CywT485lm
HiaGPLZAw/1TKTxT6wVvzIvhJyrIHCusgzp/EiNAWJrDWzikAFFzVyqQBSAW
9mYipEQdmrHIxfQt0GNbplRwaFEqETCjh4hMyyzEZeJxHz3ior0ZCWJ2EpjO
Yfxvh0GnzMP6KNjU3aDQX1H/k4fdeH5bxWxbWammm95IJKehH6rmLcBjQO6D
pZYmDUjMmRJsmjXObKBHNNkXu5PobEgN6Qz/lmztpATECqLiO3sSm02ow+Ue
7yVF/utRydKWLPcDBpGZ+VjhZI8nUms0XIafKk85elnk2SFLOifchyiR84vq
/Mi1ZjfNoDIS2w9DJdu1ShrLjH/vg6GOxyzO7ipfapspxjRE9h0TQz2osb4I
qEK1qciev3BK4EZETXJXU7BZZFk6o22C9QF5Zy4xt20JXQFzR3AR+Vlk69+J
cIALEAEXdoNeyrFqtiIX0SkBBxgqIino+b4t16GibsS4/IIZIKVo2uDif4jb
2lh9vi2Y7PyUkCfOWtF/rA33RCSkegsc1sjx9XF2jb3dbZ1G8aX6nujUNxpO
5BOojgfmIPLX0eJ63LYcUNn2gK5aW1n6SjaIbQKL9dliOZfIq5YtSfhC0R9X
yRE+8lwdkXEszOH11wKD5xBZwxEeTK8SUTKSGYoZhxk4I1IqF4t65I+MhWEM
fyfi7/plgorOMvb+yABJuRX79wLRNLa7KyJ21+VycqFtvGWCxZafH54OQ7I6
A2e1hFVoxXvuMdFYwWMYpMXiNvXyi2tIAM7E/ZNvsU8eu57CzX+fhqhmQezF
GXUsj7/Dz+j8lOsC8G6tUwmQi/x4vr9mj4g6K7er42UEdiVUYNue/YLW+cg1
RzawT9nCyCvCQ0mbqPT6tlCfjmMb7ZufPYaej0eqHJic/J/WlDKJa9D6C5v+
+94M8cLboVLBdCWkZhLuh7U4LuOfL1adeC7/tPD0EJ8QRsBKCTAiBV3Z0hfx
/coumLo43COKsjUqEgsb0U6iun7PQ7dngd2Spp6RJKC+Izzx6F5vfQJ9vyOq
R5Z/sDN+I7F52TUD3/CMPo67IyFMJN0/hiOAPf+jm54hepKUS87B0UNzUGqR
9DHCVNp5aBcxctBl9R4w9Bz6r8xSQTAU70P4Emya6mchP9JC3/MVEkIt2xTU
b/Eez30rNgPq36s0gbgbIst4mszQKZVRRtRGZj2G+hPqjxDWkj+/65kI2Qf+
c8pwmcvRYjakwLBL0NV68xH5zW5nUmx/Z5DafyJiYQwALvTl+hqO91XOM4UW
B/7TPurC+bElQozcSdTFoUL0vbBqUktOwVbiU3RFhz4JZYCb5gPwVRM4Qe3X
MsXZndWGEa0pp3SDYloShS71uwEyIyZrrd/IjD6qITe4iTBVaQZ++dqDomN9
aiyV7kBeiA5VLtz3ah8WMKJIZOiA59rlFV3brybIWt3a6j8WGuNVLi+9IiZL
BJofSl9aiqSaCR2MaeyK/IAh1jVJIAhRJvUhb0hPKWSD5k5Mmma5i6IfFUwr
S7upOBritz0Wqt/PzEQJwGR3lMS0hzjdI3ofejT0WjcEfYcRMBoyY3pOHMVf
AQALbIA1LlcBSdzFox3sgrSU72N2R4mRBRcfJA0+618rZnjni0g/LAXK4CoF
vRRwK+gBIHr0ajraZpsKjEvbqgT1zp6478qYx9ZHSN04c4jXElkSW1uwt1XX
fueDw2lmVGHW7JLq8eWst6IBb5yO7sK9rprQeIctdAJK1ikIfd2k6nfmzMsh
AnsPp0JHygr1m8T4iMgCoqy3+SYDpQcZrRDkuMA69KtsxgNhpSh7XgqlpWpH
l3Gc2P5hvwpB2QuJ1a/mCZWrqZTbO1AYpZM0bHiq7sEE7XIatoSfT/riw4R1
kOtpKg441aEJ5Tny0pCznCvhqLuqNN2O2C+J3Ndyiy6LhKsYKY5JgIs6ckJS
ANBGfCYS7iqpmU2djwehN3kCm9pC+bFUNlNWnD/L2urN6dXEt02uLde/PZ4V
Xbco8nSB1YSgLmwO2eOo/Bvj6VbAv35WygdZTmf+tL3XBS4dIwVvU7/7wfZe
ym/yLTXVWhZ+elTLpJv5kbtWqfnmKBYxmQm1AL5jS0BY9Q5Y8qc3s0A4lglB
GB7QaTHpX1BHSB+gnZ1mWyZhPF1dEgmVZYGlj50nXk3Iz82wA/kZV+ZqoivA
X3gcXiH3I90S5dN49bMO8nmUB7TVA1oQbtHf57MWko6IaNKeQZyVGXGSUT2w
9VY25j6aJQrQ/RQzCKmlW2eAHXnSaJ+DK202qXDoBaR/fG5EHu9nxtBs1YGh
mxfIXISB72X9T9CX0Le0YXu6SJrUaLXEy9PEGNbdA7+1d+YNrMJ+Tg7wSa9X
RFYh7RQDzH4TASp3jlUf2o/qyrmvgpMpySXWPq9FQv7EIgOXy2a0zRcvkRr/
yVNZzd0tEgC1BNYOaSLJT8AZ3LJCDHTNkfGTiR40+XV2GHGUI09Uf+0S56hw
312WLvCR+kSKnS7RU++2hY9owURQs3s9TdHe4vYLfNBTNCsi2KJJ0saf/bEx
NgBu8R85IOyVyoRatTXKlJXKVPFXtlCjQc1CCHNxP3kaZQtvW8v+TL8zH9zE
DcY9rzs7+QCw6n/pE+DYBOi8wYdZwjgdFOI7wgk/RWXxYor8tcogOE1cHyCx
bdVO9Kxdo7WTFojvK/51pXXLaBPrk1C/Xp6zlY4+0K2bRieS8cfEHhD1QJx/
vG9AEWkCUYgEgWBFti/Ol7l/ba/NkKHdAgX5mWxoEymYSjJuwaub7nhWXQZY
7W4hSiNacoMAniSdSZthc3QKUOLkhbvDbBXxiOdM+apWFlpdt4ZpQUazrQah
CADOBoscV6edeHaoMoOOjrnr6ddKS9BiH7NQVIOBZS/i+awpDTQpQMTRmChS
LIYVmuAquTKq7guDSXrp/YlNPnxNC5e5tRyFeRMaeTlV807wHKn0mhVW1ZIO
qI9MTglVAqOiWhf7vAf4Fo6LxnDFLx2KHsWIS6GORNDAaZ1+P6oYhRe+7/oC
R0ST+vwSEH2zJDTA2RCXX8jUHjBm7a1hnFvlGgt4G/vFCA9Nwmeai8r64Gl9
R7iBMUm/kb4waJXfgmsRypn6axASoiVZc5ERmSDec5/kPe94flcQIX11Pyi7
WR+V3bCEK7Q6aL2lLCPhOIk6X7pzhIWW3+AW+THBscafvyxBie5qtkrTYXY2
SSHKbQ6U6poKFNcK7h5xeio7syFV0DpzBOErLkJn6cdYoa083GhjGpNbiwxk
V72RiON8fGKqwT+oqver3JHdIeFuMBDPQfjbXfK97wQX0wlBGUZWCb1cjlTc
0qtq1vqwvl7QjggQXDF2zh/c2JjR9HptmQIZyAIMPs82c/DAGuC9wPRUjpSb
hcqQOeLDpkM83+xCNrhGyM/MTU3j/0L4q+ilFWFXY4i32EaQFf4WToAm9v9t
D2kYJCbx1N5mM0g4gg6IuhSYxD2qORGWSOizyjbZMU3XdFhHbk2QJBHBNYC6
9uOVnsWvkuI6AZfVUsOPTK4BI3U2oRx3MiyO6dHrc2HPgkQNe6xx9RVQSVc5
PTps2pO7pXLLtuRO9waKDuXyIIJGgG3yWPzegsPYHv1uf/XKfoF5GEeU84hL
bNASwmSUZVhmqIQdxqfACTXP2xnaNj4obY10RH2X+rDBczFAQ31U7Pb0AciE
MVSjBDPt8er4PVotV3JK1Q6CWR4eJijp+0MLBaWJi2iES+WFKkQvWipXpiih
WcgMRuMCFI03ZRhO2LqKtjTqc8RpWRfgPyT/2nOp7ZrnVkV4IADwD3xOg4oG
EkCrvck5Bi1B2vymEp4yvVospo20ocUA3VAWYHhPsh2D57dUW99D7DHh8vet
6iO6pWcpEAJQYS33uithI0Pj3O3BLW1G6nkXVpTfvRlT/Pre80jbMlImCHgT
gW6miv6INmPWSmHspaljSTq3tX7LxXOaCvqSCDNwHmQxMrvT8iXpzW+N/m5S
9v34MDmE8fEU5nKnQ6io4omnSOEl0S220in/P2Nq59zn4+BAc49GjtBwOU9E
X6qmzccdk6sJSrTjUj90arUMZDil+JSY3nZhY2OU/5M+kKEG4IQpUOyJhbne
tkcYc38rk852JeyzT3CDawEWLS2Oezoe3yfsmqzezWZRHbPJDc/iQ834OtZL
bUGyDC/94gw6QHezTvGGlCQH09P+EHig1VI+VywTffjPJRayvxZgoVfVSf+i
Yf6Wy+DoeLbW+dPYtysXmoBk8UunItQucKTlbMmqvV+Pmqm79liiY0ry/W7p
87iTz9oa0r6lhNPqBFpcKL5BdhiOKrbaR7WhzCyh8NCxZrFpRONZQZOTLSke
MjvjJIYOpFS6TiRWhWiSsnxVauIA3k5Nbg9afEJF/dtv8xyBjtcnltowj5hD
2BueQ+cOFl/FfATUlc+6wONXxwZw6lchSJWD5DUB4maE1Bw5Sw6mYPF2SV6T
I9IcnBK0KBg0SnbYEqDjMZiWsSrmPhqIGlmZ/j1lmwbUPEfdQ621WDkOoyS+
Y8kbYDxLL0EMSmiH4wKDOvT0ArYoOeKAjrXxoY8pxyj9gXVeX4jL22RsPy5t
L9Aa1dEY5chfQ/g1TcE9XKQ+nTlRkB4JNOIj/8uy6Qc1tMAkHSE5EaHzLAxb
N4/0fFFbWkvyLM2VVz0IiEq0ncKOLvFOdbgIDJoBD0SsycKAwAUiMRNLD8Bh
i/kCeVppIA/cT74WF5PO2syz/SzDDsEMw7GanyabcYu0/2IcBWlYDAQlqoRe
Etf79NN3qWmkf1P5au+9GDMIxxXJ1cp1OLTf3QuxF7qQSr0RrTajBFHCIHWp
t9oblDabRJZvS0es9Tf2/yFlOlTILJqsXKoyZ2G47re+RdnQrhYKeEkqXXub
6mhKd86y36lVnl+ZpzVGDiMkKM2kCOhUWPtcZajy7C8aJOX6asHZ6eBdy6Hx
YwZK0zQrPXboyUEPExYFjEV+ZOge5ExRhR8gd1VjCH2ygzUt0UgABbFB+Ixv
D+gxWBcii5DWQV8FFKY75hXbOoinjMnEaDAD5baz2hDlmsrrShpg7LFPS8Bl
7OmaMv7JyT8cUJtSrOUyMntpC0B+FpY0F9CLu3m1LWJOPpgOcLaQLzi5CGpz
6pKIRRAfh7O/mE4OM3fPLAGUhMCAv0kK35cYuKqsWASu8W7nIawomZFyUice
lko3IMct4D2D3CNKUtKY2mPPdn2Xonq3i/4BKWu4MHmdB1LJOYPR5qjems06
hBPedwtiECwjIXtf0YNitsPk6d0vi4FftE0tSsoAC7BnLjoq+xwaqgwU/a51
kVdAPzML8J3GKUNfOd8EtL8n8pl3UimNSNBE6EPT3/eJwgcwyCUvcRvYb7jq
y2JiUVNgTCvM9WyG4hjsedsG1IoyppTdpZxEGw6B6WsHvbyArS4CE8bEBtTn
hW2DSocBM2mVm3ljJzsQUTam2nA0oTtD6SJ/So3JrsM4cgx8SqkD7kiHnsBE
yLrz4a6EwkK6a46jJoiwCDr7WslCnzijdak74A4ARhKLTxA0ajRp4R+9egbm
wTEQwSrU/v7ti+SlY9rOmqvxEX0xLfg4wplsoJK/ftL4sH+xqWqj92+rweKo
r0+atAmLuLCeeMdoTELGSjFcGweb9V7IbDAEKHf3HvqSrP4HInkcPjvsG3wa
wIXl/G2sSmOuL+WCf/vDY0pO7a//ckXdEmGrJ2KtSl4mKmkuASYJMVQVL9AN
4lXZz1kIrZf0n5AJ1xUT7oP2ha1m+1efi4yg5kfO47WI3CyqOrRuuiTF78bv
rCBLKtVLSDZAZAMyy+SKJPUkdfSyDF5zWDOLvxkXwOZt7PYJbfML0Vs+A+kU
19ndL2RyszcyxzW/v2gYZ47A33axt4/4DSSlG0Y1jmydWNfkWhztIPHmoy1V
+2i4usuMFaLDYgqh+qug8Fv5i8TMlOQJ2ASVbQ5N3Uih+K+pNX4lmhQDf3YS
bE1XtCKWm1/x22qt5KBLAOp/vbVmZSz/095JcGDeSNL5susFI2vtaOvc+s7G
ao2e4ZlvU4KCRN4UMxBIWKylW9Vwilqo1oRWosUmKZujkAZbh7LOIswhjvwj
WhCSucSE2MS9dpDWE36K+GN+XtFCK6GMOpm1mXJuLRcz7Vp96DRFk+5AQZlF
GMU+LAviKKDf2jf0dipTq/9FUcMz3zUQIA1qW6t4qHGhN2C3VfCCVaqo2M48
CXjK7oMoCffclBKmv8S/kNUm7ljGtcwX+QMalaTWn5LfArgTvPQQYuNhPO72
b/r0T9SYTb1trv5YYoN1UgYx9US+F885micheuO0cRN8EoBM/VvumZtDgwMy
FTVUlV0G7wTU9MU6euAWxW4kEcPQNo4eNXd94djO+AK6HWaiSyaFQtweAKxV
uvWiCDyFoO+3ncQxDy53Atf3Cwn4OahhbN+tLgXWdYYFP4z6jaUh1+VtJItN
QRvxuwfpRzQqModr6unrWs2F6HLe/ZKzjf96fDtTlnxl5eo9cSKpvz/WBwuF
Y0p678SxByUwUHC3NVKpRY2VqKen5Oq+fbeuiSf3yOeShV/yO9OI7VryZyYw
EgC1QVUvu+FtZF7h+Q7IGdWpFlo+LW5apd47wXbSnODDogoRzC8KrNYTOlZm
7MWbSTGEdTSFOXH6B9nEqk9QqotJ4jy25821FeE7fc4dVh9M2jRaKsthj+2J
vnK1AZInyZ18jCVeSCDPMfb9BiP0zQYPdKdAQCbEnf98j7CQDhdIZ4EWaaVB
p+5WrQdojLk7ApjM9s0XrU1I+rHW4dYZI+q+bX7woOswDsvB90izD78GNjPg
LLx/tyYtoW5JM0FYh7eQbx4rLplxzP1pX5N2IdNY/pJr0IrgkJBFFD8KyiW+
yNa7v+EbXMtqGNvGKq8w3HWbMYboZ+I9lo1thGp+72hHpxVZDVKaBa8OhWNF
UEYkfrfOjk6Xn/E8tW8tFEXXoFT3NBclZq8VcaQBsCI4Q84qzNPh/prxSiTS
mmwLuYlRxypxPPTXWk9PH/w4if85EKUj7sUJLFqKbgI+Y10ZCgFtZoSn8orW
0oMjwtm3RnpCYwn7e5H+zIHdU2h4pLYIGkgG+jfOZksOuDyzG/thylC5lKTL
wIVZlGuiu41KlaoVAgLtadYG0X46hlOTHXh+M5smLACVrV38Cotv+G3lqBns
cVq5o3ught61SYgBTIQo+J7jWWo/80SvUgCkl7IgwsCl0JLqKe/fk3dYrODj
KJG1UF9yXtpiCXxs8YclJWYVPjwzWCc72Zr4zdhgYOqOp+Ysbva1jWIpno5B
en/1oueEuR/cmL9u4aQDH8Jm8pdHWRkFrAEdRTdHrN7BVDZoxIQZhk1j8VXU
/8KiEc9GrSm2+zClH7yPxfTYa7YdfE+2vd0QLwkI1zdUafm6okvJqpFLh8sZ
3Pk5+3ePJbyhx1Zc9F0OrXgk5RXr8IUh0edUWv/zPAHJMVh0zb+SS5m/ubzM
A2ZjrLElfce6tqBhGzPUzC5mMAnOpXn6xizhcE86Nldgq8qOXP0TANDir3FM
6zCLhaSrBAebJa312i4RGurGpUY/ubOl988zDmNXSXQX2MV//34nu3/xjYUE
P6UEOMe4KyNp04UU2D/ZJS03O5vNonYtHMPt8t1fBLZ7Jf+OyOl/gGgm+duJ
59d4ku+TXnsM2Q+1N4WiQdwttX/7+xhjjvM60rHRjmM4BU4Fi6RHA94XXgH3
ixC71pKCAoC2gdsldrulslYpgBsSKFoje/skXHm3Ubma6xOFUv1ujSMhyUVz
TcF1gTkvTBGVlcGBV/JTKvHFVtkLLQFP589qlK9vmaUqI/CvlvFMPwRQ9k+z
5iwM9345slYk3KY3un2h+STX9w+yBRzz7lnCyn/T55uCBQUqb8/q3SW8ac5T
ZIIKlSxDpzkhZ7R19jCX1ip6JY+KhrQgzqRuk23eYsx12eLmBr7xjVXQjFwK
COkmTwnMt/IzreFREPh4P5zjVNxwxXU9vHwPEZLkADxm232AnhXeSt4dCIhV
FZwCqeMRskPzegSefqw50Q6MAsxHKOKLYE/HPOZZbazz+VozUP+ETvADjnY/
DVt5UlNbhr+w1k9WsR0EGqsTTA2F9999QZi0NFXhuqoytN9YLqC6p53FR1j/
giWZfkbVAFB5uqx74+oN2XswK0wMiP/okTBiyEjq6SfEBNkMU2I+fvwoIuTd
Bhe/D5XLSP6xcmL4eiJvUFPDaHoRLr3s8ioeXA232gaGN39v6iD7jaNAaB2G
40wDVLuhdDyPqqeZTZjl3IDfmScO+4QGr4PM3nznxDVneBcSxiRY2EubA3WJ
0U3qS+6E49zBKs7EZM4qMTwAg8v/6JFPwTgqiOmGIp2c+X8OuVjpgBOsKCOe
aD0tiDQAiKTKReT1CSQceOIt69TpAT7kWG8QxLiwlQHV+gORjb8BQgWVwh7i
vvIvqz2/EMnSwWeDZRgMiQS9JdRdbw/nyala8qhDBFGgqJ/cJA/Vgt24k1uz
IdhrLXCt/EaxmFAGS4NWkJh0scchMPuWBrXPeEHen6iQlJTlrG+dMKRjTEhr
WZovnDD+I1W2YE8LgfHgu91+Jgx9HefcIKvmOqBx+ivIpmzyuysSLPKeRLTs
KnsGRBNrOaISe6oYC6PGSXuKJ92wWGBsxGffBZGUkzSNhtVovwpd9hbzMbuK
aqyF3K3q0U5IWJtlM+LJV7V0v0tnHrjDqAuA1jufI+iZ3zCelGPiLLbarKef
Y5Bc1GPycayBiAZqPq3caRKY8Vne3Jbu1ZBIcBFmK68suMiO93Xo0+TrhKpH
Ph3ofXBzNkwsMvOQSZLMc5raLwrW0pCW6MKAzGA8ua5++21Sd5K4CMAbN5Uv
9ded4sOPw50xpPE5/Tw0X1FkTSXS+xQesuj/whBel4gzMWOUUsfm0bVTXz8j
14kJrLdIYWoVQI+qI6wGUog9STklnbFnwmNErweDdkvHvCtCPOy2hGAmNKJw
/7PkxSkIeeZSFXRlZDUJ2Yb7qUGnbOUXRXCa5xqKHPhdTYzyWnt+rwqjPbti
bYjL2cTKmHenqiNjJvHUO5XxWchMzMbraDK+dv5So9FTGX0c79XYrrx6WzFL
pc2crUA6V8HcDgxnvm8JCyr5C/Fr0EfN/JIZShHDTE1VM0wemRROLO/KBb3v
Bt3VR++MamqnYWgpIf5GrPEDH7NKICQfGUB/6AEjao8kK0q0IVt1xp686MV3
KFp8dFHlx/aGujhZCyCv2wyAU9DpxsEbp+P0qj9MyCfNNQaAAyTMv8G4OKqh
hBNYZcdhzQ5/ydG+fzSzc8IiQOgXn0fRJNj2OyK0Dkqe3aeueWP3YOGzDgXW
ybmYRAbuhd+VcH2PXkbJLxOF0FIuI5FCtySBVMBJG6HO2fO9LdOJzepK+vAD
VqWMl+WtKkZvqqye/wvfL7YA6+v9OpmHkOss8OIHjTBrW/YBAY1/GXolRH+C
oolrvOooq8xKgOrd0g83M8vxyIYzS5OLHvg+ipyWLWQmScLJXmNBkHarUT8T
Z7cIMv/7tgFZcDkbt+VWkN4Z2ns7aE+D5w2cCxH2Qd+1JkCij1/c7Ah+1p5K
JTWwuD+7NBqhwxWqRIlxqdklf/hfqRSGZUQrr00doULOwXz15qc2WNE9OQrh
snxGbh3Fwp/RLRYkjwrdcrfdTjr7deCY4b6jqIH1JK0NjkDIXWITlQwEBP8F
7ExP+ar70BZ6jQKIpWvInSFGmudHoun0WvWI6Ko5n5DSIB4H4hvnsiyZq7Ai
slip1i/4/xHyoLAsqXviERMPzMxEAC25KbEFzs5PofOGbRosWGRr3ME5BXkc
9wsfiYnN5VjKrdlc4LiOci5/AG3G+z1F9bsx0lLaKbqwmwtSCZNc5DN+PIZT
p9X73Z0lCMQhczj2uQjPIc4oQ4agm0M7mmE4tY0B//Hy1FAbmbRk3MJRb3jN
GX/m6+x71ClhdPPM1LS7D0xCWYQwKP42mh7706zMVt5D1sljqwNCOODwCXl3
5nN9jQs0BcE91zAP1qvPQIyEEBJvORjfEcAQZYcd9NG6AYl3pN/6+n5DE7lF
SK1NLDyXel1KaaEdV2mXAqOEHcG3cT+7wbYbccVAUCd/uOUSs06jjENvaml0
0cOOnCffCAG1vUVBzVIYah3GMvNEVVsPbsqX4KNK3GYz8GlmB6YXM6UBH8cT
DT16X/cnDn/VWljdUs7H0/S3SlqfuRr25QimLcgSMMnHtgyATlrqzbkRaQtY
LkPs5Aac/dD/mlMtqhiKBAdKN9SFIXKHnlHvH9uv7spBxGAzwcIXjmMQZJ5F
UrEpmQqnYP27EKQEa9csj6wy70BddAk/osW+tujIy3RHMssKQbmqmyuodsue
7hqKF5U82jfZSVlzy/4uLJk/RZFMf0142bMSf8mb+bBSiddJlHy2LJ5Gur10
52ATTgQiAqAzWSVdMZh2ZfkYTHwD5xplFoG35vjS46hMwDLBDHIldWuV0lHs
fEeHv3fUOsdl3VR22GPd9dscZFYo71Y7gxHEK/uYRMFNOWM8zutAOCkwN7Dj
aTUpTtCSEbfkJ8wuRuVu3ONcNLEizMmoFT21vkyVSTN5e173/T5nELjO++DL
FH09IJilmJJvOmpHutB/8wQSyiTrFLy300hvF0fwkYWzwFZ/QhGjNO3z9EX5
JotTiTN4h9MgTIrO/QjTBHuWyh9HYqP4EZXa/E4is9CNJB1kM/y9DykZYWch
w2Z8QGqdhPwHEBiSclNsRuSRiXjL8jEDJyWNiMcmrHynC/SYjrFlXRxZEhK0
lqN+Gz/D6UFywd5HdCB6EeZ9Y9LyHigLNvWvspkpODNMrlgIdOW+kq4TjGBT
cSObokb1jkk8MKaqr0P2ZE3qlzSnHBLT1zaaRQ1icHz6NeDQgj8F/pI7lUlP
19df3b5yknUa5+rkc97O+EuE73wG47WFUVRsCMapjvQqfcqjg2m5fOlx+7Bv
KCIE4uOVyri8uTkAU3NxJ0xNvp4gnn1HDs4LMydzxDPAx3obzVDq3ZDaGZwo
yqpTzaz+Px20xXzla0dzmng154lno3rrRnp9cQJj+dhdBaS4ScxSwNnKzCmJ
abs0VWZbAQx/0BkaV5betCTN9NinWWL1dUFsZTThmxJhQeBHh51ne7AWzVkX
w/ZJNWBn2O+MmLrATyr5MT88oCpVp9Ve+e3uSgLnwhUUKAWMme1Y9OVqamH8
YOdiJAgTRqC8KzBdowcPumfr2rduL1Uwr7TQM60fwX9bsEwrhINhDuQeFQ95
jBZR1FLWXGyG8fn7li6FyT+LORuF0z6WwYA+E6WIfyvp5L23DSnumVm/4ae2
4KP5ULDw4CDRcVYYff4TLXMTRIc2tcFohqZd63XY2eTOGNaWm3iLLMNw9z6Y
yWT5c8/JgNV1UfCi23XmYyK7rRl+F9dZcSuY3y0iIsIbvGteuGTNKqbk8ElQ
zB5jUKwTF8fI7cSiWMYhdwgLZF3OmMXnyqIL1FiGl1NoOqBObuDWMDadDwIm
FcBYH8FQ4evRf+SWiyEuHMbHlUvooHN5NjQw4KTyPs1n9fC2GlooW8jWuQYW
lQiqffiNxnfgQDeY6me2oDlkJ6ztRHuQCUu+Xzqgu57u0R1F02WIJRo4JnCR
FnW/C5z2tw5WVRGo+8ITJ1LbZNO9YV+jxsyaKRGVjmus4Uw9xizMH7gE0aEK
vzP3h90mauKPWXH+gudNjDiRFUHAemi/oPG0AaCj3w4L1w0HleAgLc4Dpmk9
9w76Mbg7QT5uOu6eARjghzbo/NP2mPHaMfhaOoWm6GsUSEUoUR6rtEiXKR4W
CFBLJqqeSmNLuPSHHzg4Kg+/oJvg/14qvrzDNhTQcsSubcEQVDo+aS4ehcdT
JAqg1GzEfPhmJltrPx89tnZG2QuOIbRfN64vCBEFEuuXAKUpm83EHDOjYEKK
dCdbKWrElaEJO67NnWfrjNI2FZLqqtl1W5CWV81O+E+dxBxkIzuf2aeiWtK6
zpokyHyFAfhnBkIb/UTAD+DEAtdw2JJ7cO73KUZYZMLnzVhmG6Ijz0VtNLvB
jkwMboafX2EyNjF91pgEbMUnmogE2KeqNbBWkkSeCzqvokLmC2OVjL2ybA0r
LnNQPDRLYkz2xpYYpVdPpdx3PBYuf+4XP/7QcIO6sJ/dMz1M7rEerkRHUBPF
P3vzYivktAa49ec/72/nDYJUZpeQ84B/Ukj67R5ZE0AZ9OXkqr7UDLkskm78
wBKJF5YosShLbBx4/1iNe8P9Yg789j0kfH5yzDDHyiFxicgPdgxzOQ9wxKgH
bfaDkayBj4z5xt79/PoCZ8OS/4IYTgKOQGdfOXxzQ31DbZoHhZDVTM3l6GXt
oNhaXs+6xUIWXYTi3/vCcJX4oVd/xJTm3nYOLwd70LbB06ObdeDDACiIPkSf
FQ9RP5ApHhh7+6SP1Orc9sJOzTjfVrteVdxzK9A1xTi05uiN1ixurYkF2Vjn
+RYqkeHCaOZLKrfY1uAsS3QYTH1PuNwVW2QglPe+fFS6SHNVjLTicdJx3tBb
lOE0CBkLOgp6Oc2V8Ivpi1WiPPCI7mR9ccAgtDG9X7aHLEM91rPLShkRb4Pm
QDQCDPc6Dusb2AjlI3Rpv3r5CbKy+wLpKtq/4Wy/LTbEcbILX0hTft+oZ5KW
xihjdFFB/Wo3gUzDc7rVfwofPveFe7N2jGB3S+5wdnKVnxuLbtmDCNfwCHqA
vgc8SYQKGmwaQVU0xD8tBLDTqEywh8JM2zrIwmt6hDz27Jg9TQ4PQ3D3xnMT
F8HseEHDDPKo3ezsjB84KT6BKpfrXkbTY9QzV4QF+HBYvudL+zpLhqOEL2Om
mmHTkRl5jBeVy8ixEAlYyLXzeAxqhN0ZExs6ABWD5tGcwsKp4S/6oT4I/XOs
cXx1Nn4yVP0sXPM+VX6XxzUHd1MJACyX3ULPZ6rgxp4lmoZU2ihqTdAM34bK
yF8Kj0WgsYhhmelhjv7EO+W7q2Q27MTAfWBKs429zeLEiB2hedv2FiHljp5G
SEfHobg2wvlC4pYaTRAOReUQqcD2z3nSZRiYn1FtJ5vjrivc+MeLYDtHayB5
h/SaFGuyOUB/sejg81NQs6CLnQ/8F80DJWymGtx75nSGaGn3teQzLTUsksDP
RUsAlWg6wOzIPNI6XEgM0oZIqo9PkO9JI1a51zxiATkwDigRdzwNqUJeI67k
ladqNfD5ual5sqzANSyFlVBMVYPvKWy6Mhdz6Ov5JOZ9m+fgf/V0Uj3nRkvr
QitQmBiQ9CdM9sJkltPrdkco3vBtwrrqBTOJwjOAXa5tQmMqbTTO+NS18VDF
ig0EL84MJZ3B3lev3mJFTpKTBNQ58WT6V+/1ZmASjTCOPqWnnq3cKG3NZPzp
kQd1etZfvUN5wP429fQab5abmKOijcD6KVgFctMlP8ptgcwwQg9IhIk6/dhu
4waT30f0HcPFqYhw171kQSSMZSqE7+Fha7TejYTCoL1cBZireQ4IW99/dayc
tZlzN7o/jj9LBYFi4B6kO9UqI7kHhIHM0+P4wyQQ9v7vMjrOhHg45pgiujLV
CSexdbS6rvM9SCx3yDIHirGgAZFXVTXyNrcP+vrUY259SgFi0TPtZF1dOpRe
nL/G5r48nY80hPMlgjtPEn1CkQlyGgyXPg+aiHwDodk7yXKxahcCJ5vtiNRK
nshBsCbjjHsXG51RVIXMcYysCTCectJjucEue/J3K+JSP/pwnDMts2zqzYGf
8Fzb3TY4WMDW3BOvaeUmWtEu+OE1QUSeMtnd+wbri8nLJnxdiKT+reZfIb4U
AOvB70WBWJWX0pCIJFzfVlLgNt06P2bpBcfNSS5ES8VzyARGPtZMFw9hoYeB
4syDqaYLTP80mnjBfrjpqScwNM81cIlWs3XRTVOLXfUPDxsZFjb9+bclQ3/L
dgZVpxsxdfLxipkrYbx1vOWevtnP7ytZWMYib0aZsz+gOiE+61NB9+tzVoIW
AhX7b64+mMGVJ548CSsR4tFYFvLAZS4fFrVGphJYH6n8fFJyOdrCgWHXX+Hz
7RJ2YuI1gsKFIx3+PvIZCUCPdZRM0qIkroNGEn1g0BfLrAP6gI5A7mqWcr5C
LSb3sTqIqoy6Hul47iFAj4WBGYHfdhG0UU5Qbo9quzj731npwKNru9IexTKp
i26lhZBeO9zkDwKIV6FxrRl2zfBl0qziT3nKmcAYXLl0+TN6u45dkhkBWPco
C3lN3ut+6cigur1NiuYOVr1yzfwiWgAd16Grb0D1awdMbWa6L8nhCDYiTngg
EOifaL+5DGJx/h0Kmw8GbyocjFVqNr71eDsriLcnmk/ivezhPJXhCX6y5mUK
CPBQZUaCBPAo7XrG2RgXS2l+eQhh7GL5tVGOyNyMqAn93giwsm8Dt5WP7tS3
XVb4pneL6tatrLP7clAeg7FnpEm3RYapSu9t4vuHjTPKZFZhxPTHQn5bfuSQ
QuxJHSpwF+uMSiGAN8b5iiWyp4kUFLrFTd+yyUFjfdNKIVBqD/HJiGafd7Gb
DfzwyV/qY/m2LUTrkyjn7ZabDFSm4uDUeZ/PbT2QLmbQdgXCCB03hm1zQRec
YbpAYOUTPJJv6DsHW+vb1J/Zqc4jdfwJpXerPMufVdjU97CQsW7/jlYUMT0e
kEJI5r4nv9msqSjoglp7oiVE3+slimS3PUJgD9VYSZ8V0Til3W2vG0BW8PDr
/otyjTxxUwModl+ifrCskH80zHDQ/DvCH2D+9Xcv0syvvlD1v9PUmr2pXKil
s+aCw994FmKTKH4MyrOwXERwXTqn/oHXkL6OnIuRJmnIA5aRab77pILxT+QU
ptklU5GQjSYerSFfJ+ZZ4YIJ6yqtR/Vwectb3lFY05r5nOqtzfmsDvUeNx7y
aBtfB5osIYiwMvK6wTDSROmxFnkzV77Dnd6iDQbMcYKkmZFSVa5nWz9If6Lv
EQS6vKYeJPIEqEtqKQjv/nZ8nhQvf87wc+BhMF9o3h7hF0cncthpARAoaKGp
kro4CmnRepbsHPM58/lXtX+yEh6p/xWGtXPQjo3fbWbHhRhiysF0zwyX0//K
g4AEXmBJOxCxzmVMYClHdsqkNAbiLsGflcI5eMABvZ7nZNDRnOeJS7SozEFZ
UNm5TZb/fL2Iu8Z2jHo1/80EjwM4E7P9Lxqlgu9GpNmnuXj6iCJdohpIL2hC
5lw8DyCH77+qcMgxz9pWQUab58LfF15XkJLvFFcD58EtvwsUr9JiFpg0gy0f
+txiceXvYqOjHD0+cGmnB2Mhnu7VwXYmGvBXjgMfP/KEIOJocFSKvZFJi2/B
i5dDLZ6dOYjejpEELDCElC6GAtaZ5S9/j0pemMILloYs1z8kZ9mDkBmqjHdH
R8R+BIs0s+G28z3OrOsK844emXa/LUmxbzGQ1LU7DysEti/kEVEMHWQvIDUY
gREspmUYn+VlNIZ9LUKcuANthPG1BrRK+xXnZjXw18Uwo5OGm360fE8yBzEJ
9D2R3ALh6OxOck31rmWPGAY+08032eZE8mmXWKGgKun1vtENmqdtTDgmka+O
aL9pHNidPUMYTeHUDw0Z0oS/RpzTZ2+bKArMSxCYrvg9oNGljjXSPT8YJS8K
nstUvAMO27q8eOwZK8LAjjNYNFY6mZxQR/voSDiejxCDl0bUG5F/WQp2lLbX
CNgTy8YvegiXZAVx1WeXVuZTRUWWB2iqBV27uDmWhVU/LHhqMgyVgDcxWefc
h90P32rKDzWTHA+cYHGlykJDHOhqh5Gc7cpnrvd/z6qKfGjA1mtxHvMPmbT/
sjZX+LbYmLYLI1JjIUDhT+HYN5XYwtWDOrEIlnbnBv6+qP+GPkRZNrOQ04cG
OfcgJnahf9UKpDCqccks0uk/OrLTOdhLf3NWJNI9evADi6t3o/afNgONMxjo
MPB3ZgYzcX4gzNS4P8f2QB1JDZZSteOgilMJ7CFFjbcEo12/x8gGP9Ejajkk
IwOsDxPQLl+VphH/wmg8cHUbdf+5MnwJUM9fHrTqAIMIhSO1lAX3oa+LQBWE
fH6Xf40Cz4AcJYO7uoeyfhu5L9uBALEh2zWfLxAjar321xmMwhO7D6d7GCv2
Xie6dvCp5HMSbka/c3N2B014tIKcPxBKoObs+FcutXDYdIAJEbTrO407WyUD
O/B5Cdt3jWWWwYkBw8t0CBe/G6xDnKJoTueJR0gv/D/ck3RmWW+nxBj802Mz
9p+vvVLgrZWQiDfI7VdhQBWsO7YIYVVilvtHhv/wujPQVu52f508PUonChu5
JsX1sjiTszWq5Lzdan17LrFEyHrE7DMZmetONlCRtDpQ751EjfWltKYnV72B
Hv8eDuIsCLj11On2YPTORvOMiyPBrk1xCRCYFRr2BGzQ+0DATcL8dg3Tnwws
JNKKu1eP2sVaVLK/Qk9XtC/taiT6MTB5UujCpjbg1oEvkIAH+Dep3NkS108T
inRoOuw6gVQW5o7Yp3cLvRzJHRCIWwwcN+OfavqTDnScIyk2yGaS/WMjR2ZK
H7XoXhbuQ2QuJlAodt92+gQwxOsGvQgfL2AFGpMUJD7zqnefvoSb+B76Y+7I
ynDrCNJN83DTrMeG20Wq5QrjQJvPzKaE2NvDJeaelbcS1cYxPPodchF4S1GQ
LQIOrtligZ3vM4La+jXVT1l6fxlMXZMaKt0i7jwanKsJOkhHHGn14kVSwPIM
ChsF0Y9pCQ6Yt2VjPi1DCKhjea9b+m8Uo5kePFvKaD40eSg5rvzovB7gxI2q
U6DQEVVv8lG1E3Mzljyb68pTtGK1N3GxbPB1uwFeUO/qGgtsGP8dVZ4UwiPz
wIJG+xa4pGZxvH+1asG1w8I9VVp7ihA3AlKTxffMgQRMk9jC8Tj8xixiP158
5vudD5kb7BPPH1ZbEwdBbXuQ6CxNafrqImfTahUBA4H17UlLtKIyoLSQR9xo
yGzaHHdB+0kONszTcYaynVbL/0kXM3inHkvTOKJA8eKTysrUaFrOmBdHxQWs
yVS8Qk7bkyQRV8UME+eGTarl8ux8P99ptxmOk35uwNbNzy6DWR/KOcro6CQN
5J0qLDGHTe5wl2Y2vP4eaB57TY2AjLXAT+dK4y6gR8Ip0o8NYwb8G/AHJrPx
xGMUuDET0J1lTQHiY+HkHwj5EZYRoUwdIab4U1pEFpUNT4zWu2mPR6n7ra28
qGardfH4QxDPHGqfIe2q6DvglcZh4pB9O8w6mlvIfEemjlUAUizZpDc7ltH/
5qpKij6MKvyCyVjJbSOjJOtRrmmoPnmrhwJrBQag2D4eOhd3JrHxa3WOK2tM
7KtryCnpQUpiwIVgx2zQiWXFnke8c+pIbbyhWqv/xfQgWMZFmucNhXRwtKmG
bQVvLj9l28ut1iIMBsh8iMKuc6MHvPE+odpgX6BTY29rG3YTVm7QWgOKvx1+
YNmdVE4EmdrqxbyQqP/7w6MtIyynWIfSPdBvlAXf1FjLD2b2TH/6iISNx0Ku
hsCsC0HkJvVPbmI7V/YvEuEfeFOGyuy0FKaT6RN5a5mXJFIxvXe9gXkOQaZq
CON9MobEUJm4XZTuyhO8ZcPqv1c8I3ECbb2HL6LotlHalBXCrXWpmWxdnIpl
C525rzMWXxfIk/FkafoGtwuvg5rOh99y/GXCKID4+rY1hV+PFwPEKWRxlpFs
JEi0EFJDLjPKKQpfkqZVYmIC0NcmHQ1HKZpkbxg2iG+3v1k+UrArAtB79U8K
1UUgirCDkM2EoTOFRcvwcxMfreG/b50ZhqCXIHD7PqCugtRMN7BEVm7kOiRV
OCZtD9brQH0YXCUjk05dJtXDj2WE75fTx0jYl5lq2Jb+0I3fIcznhFLcF76J
I0K8OO/dV+uYsQ7wNYTcyQQt9X0/rmc5aNlbM8Yew1gJaEANrrWJdaeAqq5p
4p81MTpgxdg2Ur8Fokp94PQaiNlADI+UnKZdAah6vKPpaUEaNkuOYCjQ8ksD
1OTaTOWKBiHImDchELH1P5cF5BpVI6ygHWvHCfgLn7K6HrtV7Vdc/obuRr8v
qXORyzu2G2TV77i/cX/Nta3h15Qc5Rzni8vg4Nl2Tkqsv5XDQlslBssERINE
xD9LMGBqljQ76ctnYic0SBXjg3UTJJlSsF7tO01Ij5SggUPDe6uDvGqU+Dnf
EXMHK2Nu4KSYz8xkwlVmemT0HWueeWxNT4pN45T81JheHgJbwKRLYJ7p2umu
DDyyDVAAUlMcKoQZF0YQhwuHnsb8SiithTIloxhDYh/qDVZVgNVpAxlSlLDL
JbWYXVjuSK9uXm/T0HVc4E5WExolKsBxmdbJIWmeDhSmbFz13OSsaR8hWYdU
+o4H/LBrJDpNrO5+bVbZbKVOIGb9H0xwCL1wqbAgUvwHBeBRcZKOj8tEHcSr
fJZUFhvQotoIrqELspgkOCElKdYmsS/xO6F57NodJxsCbr8G4451hdq+5ff/
q2NGpGX+uDug9ZdtxlX8H7z+3XODicmofumUH0t41jC8JNbjfuUnSu8oaQ7i
4+gzG4IGeeRpNR2Zek5MYeO+4AIX6gCL4dnLb2xr/c4tkTIXUTTgQaKukDkx
FNi1RbbcpKZM3NzCJaSlogfGEUwH/C/SvOSMvtUs3+6IPIn/+ZybM5mMS3KJ
iXKhLbGV2ZhGtembQ8ODxAsZ1HlLhiyqlPgvxG4zZtN3OQ3yA3/I1P3ztd1N
TVkzE/xNaf6WAy5CSod4oM8FojPrHr+2PUmmHw/S2VFGHaXkp1sLisUUjR0+
t4HhB4YXMw7QcRZrWfTjQXH2C1ZTA8K6RkzwWjgvmspdmTm/Zoe2lcarr23b
5GG8R6d0/4Sbv6EH/UZqgWQrib6AGm0ho3UtzWGfA/o/ZgqCUUUXVPWcIGh0
7+L8VakMX3t8fHxRT57fEHunUhp9rkWgvMz7e9SXGGMOF1C8ZKnlF8LmFUv2
a9c28NAolrGAnb/fAT4bQkYywQZcdW31DLVxReiD0m5EMCazt/HJ5bvaqimL
582X7KjehAktyWgY9Xmy9x+dIrc2CzuwVIUFcqjbiWzZSmGO19gbbrZsYfe2
TmjwYw2v344U/E7dlBaY9j6KUWWe9K9a6PsdZXcbGiRGK1ecZETynMFM2nnV
+7cCVsc8dDpOp3ijQNRld2/kFGu9jw7bYCnDrGLlO06tgkrFeoWXC9DykhSu
/nEsP/fJBDm+x0ancv+xCVcTqpuIv6v1zJ7DkTb3zaMLs1e0ZwYj6meRXcUE
bddmoH44QM/0pLu9X8NmbbXgd7gmrzJP2rxkcxP/4yrnHzfFRic4cR1e7rtG
4C8oXFz4cM+5yp9cUObPVypNbttiakPRveq4yH0f7Q+HXX3l25fVm/i9KrKT
jNNEqb9V1s8K6QZz5MSOs7ZiuwxjCGfGu4A9rCgYxLoSVTwfwIldOuSlH+za
rlPX0OMA0PSNvIhKzyAEiPKptWxl3AcwRTKTsjaHdG0AUYMyZ0iqvTIBWRp8
pfJazcQNaBuqkUg+2P3OQHpeiilNnJalrhfS7WL1OhxWr8jNM6WeHVC+xdZe
Zz2gr/7/cxf1IvZaGtbI2XV484RKyRkj3AsKbHaerEbrbRtIOZ21wV4QUTbT
Zpcu1OJNn5c5Z9BScbtBy+MfNv0ABlqA4goJlC390aJ9GuLx5uBnNPr1X0yU
BGoRhSBS10xGGDB0iDnEIZGBJmMttVDdS9L+519IQRIHzQwq2g0qes04FaJg
P8EW8f4lOfbc6dubDrFJ5yscW2DIIj/NkKsSRcCI18M5r6plR7wPtmyZBaJC
6sJMjlvjGB2ouTFx4HzFNU8LHweU3V5Vwp+pvpryTErlXHjONqVAoeQ+IMdE
DlL84Kvhs5FAd+Jg19sUSpdOrgM8mVsCACAfc6lWCUtfLVcCfVgbC2rAioru
gfd6S2hYXRoY/Xx7NI3PfiETsl0HtkL2YfsSfzLiZdR28u3IVGM8VYzyGBf4
Y2qrVH7EOBpMRkqHiCuN476qoBX5xFkho+2qN23yTasJfzZk3Nk+V0tWoqJW
r8qdNBXVl+3zrkBkZ7odiZXio7/UNTegl49pAzCxiC8N6gh7K/uCe5InX80b
UeyE4WT05w/i68M2KPrba7q0vFXnxwMLn7Jbe8X5s5P9Y9TMUW9b2pBhUigP
XrCWpucZTxzwBkGqTGHdEJaE96DyfYKM3yPm0fFEV/rJryok0HGikUlLwMKB
9fVLbDUMCVwAwcjaAftrPPO7Hq/99y4N1yOJFmz8yRYOV4xhWg7t1EdP0lbT
Vp5bK3UvzCp/G6lALzr36xX7LKo9kguq7H6MHeCJGgFXuSRzLo1Cqrrms3rn
SbxCR2cAr8a8KBj9RveVkaydiPRct2S7SkkVRxvUOtYr34fhm4cZaOGbX0Ee
pNKN2EIEVt39FoPxicj5t6Y/hvsCQloheseG/8rn5dhuTnqjESoKtSM4OsYy
uw9d+a1rPikoJJWti2cwKQRe5bXVuAyUjNzv+yS8/zF0cOk/4LoOIm94gLWA
OKNe6hma1fwFpMmhp92wFj8sY0r2wT0dD4h2AVpmJ3opiQrO6XB/A6ZtOGdO
7GWPehevUgw+veVr60po+hRv0LYBE4dYzBz3apDipKjhBtbwLaQqN7GWOwHo
a8QGp0w+ec5kuSrmDDFyRv56AYwes6Y/9LNO9Ax7EDcQKgYmNcPgv4Q3wFYv
n0KiO1kD7ovUBC9ey46EsxMM4M1AN69EIO2BHP1DN8byrOo1HQYgrXVAQ1Rp
QQwnInPIt0JRFfyYa7jxAKrsxMi3fFfn+RwhsiC1KJXo0ISluKRdnfTSJLbW
NFscFYLebYjMgCLvWf+jVXMGiZORrzfi15erYg0pEga5l9GdJUJslCKY83k6
IOggkFoVUrtT0Y/VHPAInZMejTKxaYXDRiFSbx9+r2qYVgjlA92nyR8eJf3y
bhNvEoUYDj8RD0jnOR0HsczH3PJF/IHf0Vcwl5E9yuZ0gIJKSzDl9hOqDHyf
PEkWltj3m2r9U5t8U4a3OErufqDMyFtr3k53v6r+ZMXC/vbP5kawakkBWhPi
xMIlRMCw/T/t0wgUtfq97T66BviWJCNmWf8lStqsgrfYsrqboNRoSSGj4Lzn
kHeUarDIznjkRQUOf+Bw8iaUtROfBXV14AsHeiMgcWN0fCVMoSzqHWM1lARi
ZitUk0mWS5CYJwokjeOC6KF9y2eHwuQ8CY0nL5uy4y0DBnLbRkxmRIwMGdwb
9xnoDZCFi82o+WiTPXHqiNHcgktI+kr5dipDuElNBRArYiU6IP2BCU3ljQse
38xbTekeKSYPwBzBshILqiPLZF6aMGaC36aOGPai+pd26/dlgwwr9rOrZQEV
DFmOW5RIqtION1JGgJ20Az4hcCXS/O/9+id+Y5KCC8ujta9sP0IZm3Odgoue
zleIm2ixYGQwW/Jk63n5SK9L+9VDKnPkMZzcjEJoRABsI1guBjlsruq6AomB
ugMoiOhBun8+hOOtidwibjJLlIYKyh0re+RY7brNP7k4rjmntlWK3xCCIPc+
N0MvkKjrmB9Y08Y3CxtxVBsMrCx0mA9rWKNJ7l/RywQVYAqKQAnbUB6rnqcZ
cEq5daUvcBh6fq5/BpKjhhA758mHwQek+xDNK+xdqVbGhQQJInMEMYvb0qBv
DwWV4TMkc6/eWBx5MsqCEWJ7EEOjCqnfzngCJZNZp5CDj28C8rrqhB+k/U9W
/x5r/n/Qb/7qcHuoZyplayVmP9/k3oDnPtXyXBiP5Rr8ihULfJcF1jxTNKrK
qM+ySh2ypWc01ar4xnmCVhSVD4pZW0y6AFTI5bJgIKp7HqxE19ffyAfxMCqx
4Zu8tAJDwy+yaz2gIYadT7QRJJ8yXe5kH8agTXDIFFn/06R2WFQSc+Tbhwa5
AEiDAIUDieIgAJ24/oM4bi1exs7DNhno53nxfD+3rfdSRsUYR/38pQSq9RBX
IUEYtTm11zAA40opDNtrxQ/K6XVD0lNNvexYWTM+noh136KlE44pc+5S+agh
5KpJYTro/EHqABEh7AvJqfhLWeykX6YPoyVrjZEzVAV9bim9M6uxIKfY7Vf7
QQlevU1G8DeoFqiIG0auxUs9MJfCfGUU0S10RnM5wBeKrFjkcYFN6Z7zeJUD
nY2qYEIOSquctg004rNZmA9DlRsmxVKcEShMFLofGFBfYrI0c2RTKsPg3FP6
i7QM9xTYPk5ahSKjkCcJRdqfYfIXFr06F72LCMWF/iMqK58Ef7GuSCaMdhn+
Zz+A59BjFAbYWAumQ2sYDn4qdaJgYN47tQpIPOJR/fGeUcILUZZTAD3aRuwE
wuVVdm1DQLuRwJqxWoM9iI1LQcq0wzrpkJVip9LYiPyxMsIm7xkf954/0lz6
eekqL5t20cNkWBuV0EQB7DbSszkkVvMBp7/vmHQqXz1gXJeC0DpsA+weJNgP
xTGrOaZDVUco0N7X/BogzaQbAQGimFHrJuwgFJ13imxP8J9f/pI5+62/qlmp
GhzGvSE4fQyGuCw8h3FaRlKZQgILnX5zBTca0APUls2+LEk4zzFmfEen4Uzh
hfQ43yLQlDJ1+b0z4eYnzlwKo3Uct30M5KeCbsO0uKPV+nM0pKm9jYtB4sA8
0Gp4Zkdp2Gi2vKTjj6objc3TF2Ka185XWB4bjbMjCjWRNE+h6ktISBP6gEBI
Eyj/t/Likawu4MhfO9eM2Sw64F2Bp992GZNgk3RYNtSF+4TO1JNQaCZaki3Z
hQso916UhGfJZM845NPLMIptbVN/32VTrxr3FB/4yw5Vab9bjZVO6/h3VM4+
SSGwYNNX7saF9WQq9yJSuLPuuyw3C++YLMRX2fXgvYRZWHKFgX86GXPaNeL4
RZKfqcUEDdEIpU+giaZfLJpznlvaFF5X5NXWVVzPpeHju2wi+tlhJ2oJ4Rls
HQvRcpXSQMegBi9HvbWHZspsAej0xrb09ZtdWHJe/fi6H8W6fDaBCC0H1NvC
tfGxH6VFHOSJg9VmRw3WsJn82Gb6SUlaKOcwqoKYB2q4QhLikOhP//reYbVf
4Z4AGqAJ0pboMPnRRINiYJo1vL5UQee6nipLuEEzPE4uayPuLH6K0i6Tj/0/
osR42Vq/jlGEoZeMLef6A0Ovc/UKrYhKY1yPg5KUCBXJgzBTdeT7neiZOC9a
E99I/LTH/g8Jj2bJzQkOIWx/3QE5WUnSS+4rnTyemTVgJ0zPW7OSkxZoPpTg
qay2X2phfFyjc9/K/zmf6kgGrxUiYbst9y7ZEExEE4NJtcybgISF4oOHLR1i
Xf3i5tcsI+h7dVNdKQERqWqGiP/VmbxEhv2QjtvYtmjpv5B8j1dHObnjUCRx
rakEs+vH8HA7TC5LXKsfdRE+Zi9Be+LqT2f2sExoZFMhYVkugaca08aYDNv5
rZnXvHNywS6dkAuKdMZCfxOM6W4LuP7iTNSB5smFVhQ+u+grLBcfHfR1SMEE
bhZI/Vc8+ZViN4f8r67eeI9zGLbKI3DFdkfZabdFCJWbP4wyL24VFsjQpR6A
JbNCVNYNWzl1CnwA1SFtUs9H+FPYqSovNXc/DU46bH+VaebtwRucH8cGRtvB
LrwgL6v6mIjRftSD6Y9Jt/GtDiGOQpZvTe2X+kukVHvprwOK56kb8MS5O6LE
gQY+sw6bNT3qibutNz/MjTOZry25gZ4OAsvvPnWQmycaFkj3+msysJ1f+yWA
A4FCyjHB15VF6uWJ28cO3rUAfsnyguDVq6iXf/Ks5pZI2ZTSekGYpgeJ/TP5
7XosNbdvLbIlAMBB2U82KWoI0+ENp0ZPhziu5mtUKiwUqEvzAD4g/qaQIjSl
TO/RxRJTqRiQlbAjVOSQdGKLosTiKtmhInLUsI0qHzzfYibivUoktwfY2PSI
OS232tcNAtd1UqHz/jqgkVHvZyfTgCBxr7vyXhZQ73hx9EGKScV848RcAPOQ
z+zQF6XCpFS4FVv1eQYPtH6eRFoqX7yqEPMPE+pHqQDAn2l+so22H7gexd4c
cwZ4KRwiSoeqShj2IYJkJvwQK9GBVYPIEWh8ek94G/sK0wMUydH9YnofunYn
sWCpEyDrV6SJpeXZvBkk/nbPIVJ8XHsdhWtK7bguEf8fT3OrPcc0H4FO9j+B
cYK2mvJGMJzEhZnIuzqxkpG5N0NlkFI+joroBwTz2sb88WgMu3thh3WIYFJ7
X7TJcJuAjB8XY5BhGP6f2q9qFPgsH4VtxHKgFSio67rULLXsX2UOJo77zBVJ
RBZ8SuSu30e7iIi301sAkuAG8mf5FNOFjCvG8SiRITq6Bdo2nx/qBXBvO9HS
GBGBH2A6w672cxh/nUv54+cKbG5pnPGTZzXLWg3jOhV5DGht7BN8wh2AfP+v
L9L9qdg8HvW5NNP8z7EZJLgwpFLd8gDtQxHz0P3I/1P49K0eWKL4WVmV6BRt
lEw335HOY/6YgU4w99Bg9jQWzqgW++pTmO1s/0UfThnOj7I2UhvV2sVGzjmO
kvyIb/qsWVl6bgNbiac87mZziMmb14wIBLBmDVfznaWsvLERlBLffvOMKFnW
rjvJ/jrgGJvPc7nw2u/Up3dpvESZ5GxF7A3adaRpHj9iLLkjqZASywO6Hjki
rgQ/fqF2ex0HiMvWFjhUjTwEs3oa+ksSWMNQvj/6BipAz/v/Vx08hhM4uGTQ
HLmBFX/Tta4e5OSql+K0FkZKUUjbGHKi7ZUGBYb3KV5C1bG8E9MQCik9Emzn
3Wv6s5B2wHA6cC9lMkIt44+PwWpVay6YN+86Kxutsz+geyj75bdjUCgU4Ie0
ZVxlO1SeQplu7YStOAPOT5qJ3HGiFyZ7Bt+NFgG2BAwj/X9OokHlP23HsoPk
AmO61z1GePdM1O0fbCHnMBCy0Eq4l8TOvR50NLTyIjDvX1KlJkBk2RvgIXro
H5d76zjUe9DL6O6HyDrMjnQSLMTMBk4HUUQAEVWiEJSU9f6NSi88XE7RRJ2w
Ven6BMCSsLyvgGF9G3RI180xJG1N+a4UwcCOl/be0qfKIJl/J4uuldCfNu9A
8wLztDB4HQrunMY7fdRsmU+X0IbPz0GDX/ph1CAkSgEBufQMHYu4Q9Sycg9z
GZyXinjnyefrMU7Gu+scPmWirAGktdDLZ3bu9B+NMQ2Qf2qmXCghJpkmWWEv
0kY8mG8jh5966mVa2DvEaACJV6JInVWeVOjT2ktcEqJZKtoLk1m6dq/BTeV/
XQV52Fn7NGc694xu22xEbLlZYTPv3VYpqCUAds76FkWDeA06eU9UPrkjTRQl
Ws+f2jyAQR0wTsFAMW+beWVMl6IlncFvGtd9sdxpkKp1sfIqnqG4ZcUnVD3S
86nX/kLHdb7tFE/gPgOFc4eoXgJP4x9q0RmSme+CJBPV7/rtfUZ4NCJEUwMP
ky5NWAxJCxUcDdPohgM1A0m9zOHMRCePHY709AAQaKxcR/eefmPPqPus6c97
/TWL6NQ4PyKJpu9d4pXaaSkD2CSjpDK7FGzAhpMJDp14IT0t+FyyWKeF5xUR
i/ymms2g/Mq4S9tqIZElsbfRMWiCd0tziu28SwigdUa5TYHBzueoyl/tuhDT
PyWsJzaFOMdr7LW6b4Rac4g0vZqdpnjvMQCeYADusrWBauoSS/zOD3rkyqTX
WqvpYwC+1PwJ8j8IYV45NFkHOaXqxI0/MU9UXqBqEeRaaqIfzcAKfwRFJZNX
M/mIzYCFw5H35kwAjeCAy19dai35oW1k4lCU8utwHfBVzdTSWEaeCwKYUT2l
p142rTyweCiMvDrj87mPF0N3svXMW0h+JxBx08K/n7Y58CVNeMU/JhM8HHAN
Ip5zz+quG1Wvj+YmjoN5FXc46HZvBKkoVXDQJ9KVFUlXOEpWS0MNCaFpjbhM
B2IlyH/34s5WO/kxXsQtGH+XqGBre0DZ+Ud+edB8Qoa1A0cnOQVbJN4t1Nml
Z7NeW2AeQ3J8AZAFAwkix2Hg/eN6Czua0+Q2SCR/ZtN9Jrefz6Febl6WGnvl
Xtpeh/eJknghG/m2XBbjb0IiFtE44ldxLtW6TgmVvcA98bkJvyEmzAvHLbMn
BYwwjwmtZsFJ475qZG2WJJekoVzc8wFfpobnm8ZvvhNVDSRXPtXd05T5neBe
O4b8LQ/lT3E38UivOUjMwnarNpPl2MiHBiJblo0rOiXHQbH99q3Jy3bQxYhs
KNP4LmZAmtaqDelNyEkd5ZiVHi3kJEdVRFhWC3jH8SRucgWDqaVsU/LMYwCt
35hjnguCY1d0Lk/oy3X1vINGenYTv49LRJzHNwqJC4dkW1tiMrKGZPUe0PFH
ceCrWfC/xcs6AuUFR30YNsV6kwp3Ami7adQCeyxkqlt4igzNOwW1SPwuRP5s
T3rhaEI1+q4fGBz4LrKJYOpc0GFlVyMxzw0JF8KCFqLzXc3X9qblzvk2BiKy
qR79G0i0zK+jaZfO4czED8rOsJV0wla6aebQh/EL8Z+fHr510tXtq8HWVaqN
8BBn6TbLYIAsVU/r8ngICzd4MUspu2el7fOUYq4g8XyFOuPNW6ldztbCGI8t
lTxmYzlcZAIjT1r22OK8KZqYvUEsEPquoNsv/Fs3Vo6kIBEfeDZT/Xe1vlfA
giAb1ySe9j4JD3PhuzsFHjANjd6Us3eY49tYJ/3TtMInoYAMTTK1S6fyvr3I
/dbvOzhISwmrD4dWNMcsGp7ocu8RShF8F/3JExWgLb/PfvMs9sy5UD8D/lpv
vAslj3mrscYdarZORgYw8XcvHxCg/d4984oTA5LWGVGFaordSPlaOuri5Igq
7BrySBl4p5aetAq5uqnJVjsS+VeCLSyVfcrrmsGv5q5gdO1oPBaI+QK3vZQ9
upKGzHjH9iHkBhpM5j3eDVCzeMJaKDitnQ4LxCl0BybVJne2ZmxOIF5CYOND
915VVIFKvcLxjn0nil+Y2FYMC88V3FBkUVu4pstHvXW4v7Jpeh/ApdGff6XJ
Q0KckTRiuXirGXR9gpeLFGYk2INi/UV/ZzQqw2wNfZQ3QBhJE/ENN965vn3w
s5YKcPISVW0WKcoJsWj8H3nh5JpHlomPY6iC1+33bI5iapD22er4oMCmvBVf
FdCHG6NBx6DNl2+MxosWTeuVQyx6Jl7/zTWedkoADUz9ogEeXIPsbuueUPdR
01nE89u9Yc0384l6bhE4gFtRhFnls+Dg6BdezODM2q/dN/+34aFNTPr+DV9R
stG4DRd7A8r52tLc6uGGAch/YMN5e5Q9oztR1F3XGKGikJwhcg+WZ6wF6Hiq
n6yNXXRhjOuI2JWI9K8nIjM0aw6aChktnmxiE37XysR9DwIxQHFIRG+aAWWB
xCQEXSHhbXgDpzH4EU8glBm4WbOtOKDxBdqTc/dHykWCzYYZ7i3kS2oW2iWd
OPij86GLYrZ7D2VhpRmzSmCzix6bGR3vsWGU1/oX+a6Vf0mfoYX0in7cLwGG
2H14DNeHCwmgBiqnBWP8K3wTMLeCmViNliVRnn21bSOLanKZdJRucuy50nSC
VQT9o5bYa7dx7AVyN+mO9J8d1QocrP6rd8zKZJ/MCn+HWGaDBDsySk34rkeN
zpvEGxMthbVHaebsMVkLWsDoRlupif6JSOD4eJh8N8IUIIfV0xV7bz2OvOgR
rUXNKT+zrsf31mJyzljqDdRYeNmCeC853yg43ggkLLOu9E+415dF3IwsymC+
CulQrhki6MsVckdx029tC/gFcYmTY2SfKbNIzYqQ8H3E7ORPzqpHSJ3YEX/A
wNk5wDd3AvDgaNJ98wQARZMGshXdW68Q9zyMRoT7rH99mxq4E3GOpNgGm/4+
MZH8rGuiLznvdL4dYS7o2U9kO98C98HcYdJHY4u/7IOiJ99SSVuZJemToS4q
u6v2npytvTMRqwSgPg7LPA5ybkfBa/6yIxq7KX1ZOMyqYdYtAl0m4WMFjDtl
Fw9GDxMY+VGiJphMhcQ3MCZPCRHvY6ksjWJtYnPbmvbtmBw1rN+AjHGjr+JL
g/bmQyoNh0vGlcBMelrjSoClFXXBqUisC9F3y+Qg+TvzUsUy+to9MKT/HJ+4
ZxyzmIJvpKElqJrUoX0+qhBZQcbzaW4fH1mi+7xE7ja3BlzKPBAdkrMZXU1v
tidvxz2/qWwcodCKkaM3NJi74RFfqU39wnTPz9iJd6n4ZRycWib4cUgJvpC5
c5TU7DXttsWEEB7AC7x6SDMtdP9IV8MkDRQjkYr0nWKfo2hoDeAN9CEGyvNz
60AsZb6gRAxYk9qETEeEcOkHqzimudorszfwkGWSIl3o6JVnUTeY4JX9vKaS
GMfVWUpVhHOOT5Ku4AKkpKb6vjgi0CRYgApOSaMMmC+K7jx9QMyas5Ehb1y6
U6vDYw5BKLX3szqnwnB/VkWuQG+IJM8sbbE9KuIcVbrolgflnBjsffJpg6cX
m23dIWRy/iaasgjSO0PDah5r6cgt2TH21yCe/tCk9CnG5DUnluqo058GuieX
zx8zaAclWlyFRMUoMVuam9Ccq7Tu4D04R35dzslBR6cKCAqhl0epHhslibIa
eJPG0Vx5FezStEfoajaBJtvxNm8GCuFFWY09vjVP1FAkNxDnhTqpk8cbV9x2
u56FyNLxOtzrLhbstuRq/Rhc1RibhDBi2cN0pNkCWXQZa5mzBND+WG+dcsNk
O1J0FGGOJ5g3DXoluMw+NskHwafOUyDDXqdlIdXWkUqrFl/fEwBmCL2D5qxI
HY45xzXNEii9z2dFPMret/z2FdkmjCltoreNgjlHI6GsDl3cu/iUclbWLNlF
1+kP446zxjS+wdV9JTXMLwWemeU3/DZQP+fZ15TDjZIIGf989dhEfmjz8LnN
MzPj8w8ydRvnJvhahvcEJPRXU+QnfCoVrlooqnB4WZH6mkc7N1qaaS0b5cJ5
+iOiJvx/gSHnrG2SXt59QrHSbdDxgApONoswETMbK1MB2HPShsiv0xsTtpWc
WyjrGMtvXUmI1aZvV5kJdcrxCXDmFZwmu6b1RM1jNyiB/n9xG1J4EAkzWZRr
pyn/NM4zIXIoTTADsgcGmDGLH/7eyaEPpbdb9zTsrukY9V3SfvJbMNuH+pR6
zsbpV/l0aC3/C9GuNREcsnbhfsMA+pzQvcBf2YvUTEG0Cv07GGJYBKoqXEOA
+0jInlMjr0iWGDPKwIG2qNsakL+ByqA7H3dOYM5cxU+A1yNUMIX6dXqYNyHD
EgoGP1/XYFGx41Az3Xjt8KyzZ04tSU7YExSbMpETMlIhVZLXQwPrZoQtE2m3
evGJaRexjoXcp3RuQbNPBRBVuUdg4htWfliQT2XDUybE2xxkTed3nbuajLl8
HmJzrq1PPNzSRWLnRn4LNYp8o1+DlUIcyqUYNTmy9y5t1IqiyBZb6iYbt5+j
Inyle3rg238wRFkfZUMt4dD8cOejWnzumQ8YUoEWAX4uDcVOWSqDWBDYBaqo
bL4uMKKZpJH9ltP/cQTrBv+vHzUWWPtDh+fGTIaURGN3fIcDYZQOBa4nfMr/
U+eCxvfNre0Phw/rgDDhksH+hT8vcnQKyxufjEBsHi2ettfInH17B//sfF5U
YM0RyRFP8JRhTy0DmtCzN/zJmd0/x318blM4pi3/oY9TZsKnIQcAoGGRvcMQ
5guzhqtwZAIXZhjgBKap+qCJWNSLBTO/5wf1sSlmt+1fF5VbxEcmMFl42m+E
BWBq6Hl+CCTCfivFxZUrDOrCnLvYuRRS+mZcakD5sWeD6wq2tijBpxHU7A1q
HDcM/ig7a/mJ5rn56T4wxOcgScn3YFneMXY2IgMXwQWhUihZArH4DcyC/e/g
/gG/KiJw/11WQGy/x0XblLMp2Ibr2WQLHyJBsqqkrZVuuHwO6rXweFwzeig7
IUGJBZsknd2NLr7oS/Kr5Q0qbBv5OAoSvqhsh+tgzr6wz1Sz1mUAUhblPByP
eHg5qatLg6d8SSouGAxlGLnDMu0qOXVM7NoVMNyETrkZ6/V0o8PmMyx1mpDX
di7lfoS2fVtQ04O1UWglkXxA4TcrouyFitqllv2+Mp8lGEfhH5DYTVSpu2Dy
+Y9Fcup8HZpRXMl2gFRH7FrIbxzBB/OMuFHAzjYT5SO5ryp1Kc0fYeEDqJqe
Px8iEdDmGJE6KN/2BNwn7M/uBpWt97ZZYzQA20jC1IGNBAMSxXhxhiWoeDzD
z2DegrowvmhRPHKteNFQVwS0vrWPzxcl9M8kMZKTUB0pKvUTLGHIyju4iFZb
G83/Gc7Tq1XlxydzLnIZ3ummAm6c4pqZnyIsGDCV8atmCBpxELmsvCu3RDdA
qipeDjGQWcI0ZOVWnwhMeSfVLBFnOHjhhI3pI0ak/2li7u9rZXmS50PtVJDS
k5Rq+Sw7v6nGCtU1rOgV4Pq12jdxkaGgla6ZSUV3HDDCqcNWljU1dlq6H/De
UEZhaxblgASg+g5ghEMxY2A5pxMCPYngornkza+i65fvzD0wu5UsRWkeVyy5
BH0J34ENgbZRw8S/tw7v5R2XqwMU00aUTFbJYQUslBO9NUKi1B0U8s23dUCH
970tMr1/dv19mrSaZ1HAyiXfaWSukSDPGWPjQxhqgrli7BvX87HP8t5bz+aS
/plO4Q9uh2E5YOWHwbcVjElTvgbtsq2jcLqno/d34Q2o9ur6y12lNUBkf4pd
cCJkpmgfgooP34cdTVNgXJ3xoLev7LY5NyPPLSlQRSSPpnWHEOf8Qo4+u1h9
O9s8geMuxgIsrjhr6/RYPqw2FqZUXuLmTjTBM9eQy62n6QRArVyCEYQWH1rm
bYafMwocC2McuR7FGanBnW4lgXvZc3kNcyPQn0FTo9NaRqkWT3/pXzBHhZrL
AdHhDYGCFUfQx7QehJavUus3J/EcbI1LRVPWGJktaY6vBa9Q6EOpyXBtch0C
j9RqsSuW3OG8+k2RVxB/OdFjsui7Xluyyv6N7D33UgAUo/IikTauCEZDbTof
lknsC3GzGDLRqnJtxhkQxuq79QA7DMQJep2obXGHwMoIwezrA79oPy3eq/Ai
IaeZDbHYkWLunota3t+JIDiGqsMuPvsgqTlmgWZ690Qrh5S99m8XlrDKUcvD
e/YEC/gir1L2lOfL1RVlNb8kWOc6+NV7XunC6qQ0q83Kg/ytA0fXuMvsflfJ
7xHdD/lCmDW14bR6Bz9C2mD622KKohYBc1yemA8lWIhmKIqxuoCnKg+9u/Qp
p2EWl2QgfOL31PB4UvJ6Ed/sZ83qx9RKJEHjGSbkNDudcxSz+cWu+99GK5Kw
N4y/IcUezij8cVMzHcRKWLfP4+bNM+YZvjbNiBCv5JlMjK2FWcG8ng00RTbg
7kW7gKpjM8NlwIry2Z9yTML0LRXX/pG9WxKKnt2hXAuuXy5CyHwMkjJLYJXL
9aXoTEPM0n6vUE17z9vzGGwan2JdF4bYpK6kRrOVER+No5DdPrlWeBVF6yw3
18wGxPIOThFG8xkK22O4rljfZ/fkpYhHEBO6ObSQo7m3WdxrhpZ6YgeLwDpz
hDaawn3/ohaI642cuzVp+CS8t9+kx3fdv4dlYTtHnqQph75AOsYMj4XM2U33
vM7gjRb/dA05JORHfV/4xJDTPs7EVAVgu3c3rB9g5sF4sN7L7ncnBLct5ORr
xhyzTfcM9BSIEhGM3MRrhVk1h3iZ+jWjtQu2rplkpL1AyeQMI1sAYO53wpOM
W1m3CclMxfde6uIpu4txrTgJ1o2cOETJ/gMTR/q3SZNfbDjnN9JTCH2J4EYb
BTQTi3pWo30WUYvK30A2+5aAdaxS4Bca0tga9PFbMmx6UcK7rUgfVx8nz5E6
cnpS1L+PTi5w6NfXYxdq26n8l6WFP8ODp3THJBg3v63/Y/GqhiHzokQfQIRc
p5NpAxg9Q3G9emhFBMk5Rq3vPvPpHEsTDDX4C1sM8xIoeExixEDjxlYi9PSB
rva25IS3yT/S8V9K+LqI41vsS2HvSRfCch7SIhW1tH+krwJL1JqUzDITrOET
a7Dt372VRxS0tesSQx4aeBKUqcEMfgsUi38vo6Abe4HGmrLM1AdCAkf0qbGo
t7Y6tglVplOYCJlcnEZkujaWWNINArEs/2H+m/zPAXFPs1Ko9MihSR/7rUmB
ecdOG0jbeBHbCNK55TdW7Uisa/NLmYa6UVmnJGeLPExaZp65ue+6wqG+KgI0
C/YZBWQANN7FnkSX69bGfejC0cliv1PdmEkjfuO66C1eWXxlE3hrYtwdEdA+
EmEpBVRgMf7JTCTcWi8Q1/F+ULcwa4lTfeKgBQhGhwx0VKOgMz7wd5zOzx8c
ALGPfjlRLeMBgmRJm+vrTGac0ttwKsX1EL/T7y0+9JttAc9QwuroWtYC3CtO
iWv9NItodE0lIvnPf4ThJaMK2OFI0C7NzQSe+XHKylGtEba4OUIeE9SWCkv3
cmlzVbb1XEGTdyb8SQ1JOnBdS/xImwJwuwWtpI4la6/oAyq1K4razwpS+trt
CP6/+GdVqX4HZYi9+/LSpEjj3QY/2K7xyveBRFk3vFnPBksgeBRep3fqlONy
KfEj989/iPcx8spEC+669YySQepZZzhDVbWzGPrj+MWsSFPhpaX1Zo7Qm5Iw
LVgYEuW8vn+4EL86hYWsgOkufLAxFsApRQPK/CgkID/q+bC3Z7UOQBeo1hsF
6q24T92NJHH1S/S8xf+yJ3FpezLHpytk1B1Rb8cyCyH4NKz7TlGtgF3fiKJt
UMJiwrXJ/dhLgrVCTZN4lcwnXH2gjZayN6+/d+W0AUHStyVgw1N9oqoFzZdf
gBUInfLjjDRM/gGOhiNXo5hwDUMyiJmbuVBwlcTp6iZdAxVAaKx3MacCj/Ur
0uUFja5Jjib/ulc4/ARmHv8qTkx3+A4rA0KenD6ugWXPBDcL+klsI1oS/jh8
WkI/2yTbhdbmDzp0q4f0tdoScLN8i/6L1tRxCcK0WCG4IYr7r3IEXARP0Hl5
I9Yq0rGmHl+OH2LKPJjnJQT6X4qF/kuJs6xCvQC7iR2ON7skhoNeG4xV2tsR
MmN1S3AGqapqq9LI41vemjy8A8+0pb7FSJa4C3pWNd7ECEC0MmBE5e/i7Nba
a4fN45mtvGowBZwX9A+m8fWC+3f7G/AOJlVdPteH/y5s12AGkSnsXFTsUPWf
catTQE98YirsaId5VMHEyi4MubYtJgpdIGrNzIPGHT7waGnm0Ce13X54BbLv
wUnNsfTcWKYK9xNLXrIvR0ksg+MeWzAgGXIi9cJRgU+HlO7hMolKC1HKS1Sb
JEd8RI8EZuaCfdYJqym5MKpFgnI9d3PHPGcmqF8Lbpm0I0a9PPi/uH3d/rfp
nqWjs9cK4VZusUz0rk2SNho2tYVK8fqlFAWY3kxsPEzwyidM/XJx0SmObbQU
tHYrfESiVoqXG0JyeKqH0ZBtPYCm7BElTKZGU+JYfHBRAG/tU4shdTaaLPRE
Mh2CD272VnK17P9aBPwBMcvEx/nzq+xjn9KETLzqiLpI+ET8FxDmoiqlcmOa
zvFGKzReiWumDWLyCOYyYLr0/xf9Q5nS6FZtZ83DnqnUUWzkNnuZMDAF57B7
myhBZPQxzOjZmGhkdrfHkfJ1e5nVVFITmaBLMH2WpyW2fOCCwAZCJWTodUvS
EDBH4ZUph2dG7g9chh7smjPT+AQdX7uFI399+odyA8VFFhW9qcQBbA6HFyuA
oNCzK3L1tYUwvz3funiOGFnT7701yacXfQmQ5FGbgj9WN3OykKXV8IqfbK7f
uNFkF7jQD1OgxAwdOLNiVvVLZLt3uEXgyYRs0il3wPVQWi5Pw3PAILyAZon2
VUYgdLlu7ZTOKH9zayCdlIdGf5QMVSoHv6JryTLwynlHvqA0g0hnkneSP3+p
ExZHPyn95On/RnxLUF3umI3iLkJFxdHP0P8SZqQT2b5hByPd4YZ1TibXlXlK
bAXuaVCRi7mWNWrSEh4cLdp2TUBLV9jBezz74jhZ9gLDnhold33A5ecST+8u
wDQQT0Megly0cUZBDTX2rukOMU3TRQhQV3A+43pXySJ9+LBSYZUfSlf65HyJ
ZwDYp2RcM5pzQEay53S4ywBJ4YnTneuhEnaRe2EHrrOK/MsK0H9rX3354mNJ
yzDlvI/+JHb7MVWOW5ruMnVKXGYXV/WHqNg3uAydLdkTB4yBwV8UcHPRaaUQ
d1qeo/YX7LbjUQV6fBDipOZPZ1L1mJGEIzS6siAktDst1k2Hbilnmn74Kguu
GoBDzRnXNTuP9tkzidBbVyCE46t1uUDO6ufIMuubeaMv6bfkNb+5hzI63xud
NcXjTRXJeq9UcLqdRTLDW2BmV7SupeSmakqg7nD5lNxPpZHcmpm6YdYCxl7B
uGI3WFFMrJvRgwQ8Gz7Moi8SyFZY417vDC4PVhEYWjbUm9d5aWX+7DzwnD9O
JyDe5TJj1wUVijyXWKW1VR3m4qazlkZcct6gm6byIJgk8VXeskZjmhPr+ctE
S2mODolfmakglgqwRduAwi8LXQvz/jq5uA9I/GBmbAMNCol22ahIkztBruHL
n0lAFjGtBor4vOHVbZkCf47UmnikbFNCNTzG69yOIeb5EBCM4tXQ6P7HDD58
+uUUyoREW/TbiRD9KcB9Fw9Ks1/CuwMSMzdTsNTkU4VrrxGI6Z2ntwxHmnIX
LLlaN1mMcXrfW8cdB/jMsY2bTfVDNGXCiGHucrlZHsjXnA2GF+Dn4E4UERX1
jNXSvf5FV4qKBzNotYUGT1WY5zo6aN7P9igW4YbBhl81cXMO3KLUCi3m5MeM
t0182yxcexZYhqfQy+3LhHj5ZfiYAK9iI5SXD9/JkSrLXcN5Ssz6QQWi+UIV
FlDheipAz2frbfSJyLeUd2o1eneWlExO6uC7lmfbFKkvTdPvayUu4aG5Vevn
oJ46TzaH+fXBrvve0xCWPzJJf6sBRPq1QO9Jjj59EMbSEksPtkoavL9kMCR4
H/CoduNODN5j+JS5zK4xbYuO3cFemtx6XhaLZB/vEGVqpLZakc+IEqY9vTIq
cjR2slo3kwVNarYVcip8d7f0NQ3VljOjrs2PoctL/OcETK2yZtSUBkEbsFUo
jIvRAWlgRJSvcojHeCAuhzzoXZB5OMWt59WowLSVIfQGb70YPF/TrrebtZjL
SgaihoeY1JXc2Ex1QazC8GvKmAOgyOP+UiN4z9Sz9hSM6XZOjzf8GkM9L9RN
soRpdy844mKhWzEXLkCiLXzIlmgZUeBy4PacTy2qQlijG3vyr1KeAAaqJnTd
3RFoJD0G/knaV9n0MGlFGiQOsfSfp98vMY9+ktQl3DyWRvEcn1faYsEKroGX
CLPLwaAHMFRaj9cUrB0KvtYWw2ooso/bFhIojbwR2vjgKwj3Ha6gjWpr/0VT
mjLzYvjHEAQi6G++Rv4LsDNpWR+8b1Cqd6fQFgjRsg87S4ydUJG0dPQX/rj7
5vg1Yi3CBtw0PuPTXDdXH+Qa/89G1kJ+HLbyzUw9vUPViTf2roZyLzgDsjhA
5PxcxHevLRH1DQcrbMJLykPmr/oM3syD8NsjMaKy4lnLebfUCndKRwXZyOkQ
cAZlLn93BPxRzPWnXlmLrAtqwjKtY7o5H8aVfwobr8GJrXsDQKIm/+ZFJAQR
Ledy5tR+RWrm4IWeKuYlak/DdheUu4hIIqir7LhOlj888Szm1EuPrJiMEaNk
OFq9WnFn+Rk7se9C/VcbT0iWJREZcJdoV+RQhoCk9jyvsQ0RKYCVocOSXobg
JxDZFcPp1V9q1ao/F1Qp9s7nJbZIbeUxdhkEyXEtoW/Ge36nnY4aybERZzyx
abh7ZhIOodVuoA9oKlt4r5hfqKTCiCDQ/PV0OKxsPXL3CLTZbzrNF7NXWSMg
bgNKdZx9L8DZBLRa5dDBzUmkKGjizBWH0Lc6Qv7xANK7OIy1Wp/rxpRxNOXU
e2anoZp4TdTrdOPo8GdibDprKSig32ssttu2m+clIggQdqJkkwtoiFINL2BU
3TXdFNWOxM5q3cVkNlPyvVFofbTcY36Q7vgfcSCL4zxAcTQmZsdzyDcRv60E
CdiQRCLutuS3B604EyCKhIWS9hwPRupQeLmRVvPQ45yrGuALzi9pijyGGLsa
0xu2QfU56w7f0Dv77Ggq9kMO67wU/TMQQQkhlE4gZtXNbKMHMKdZMczQH/Yh
HFbUGP85egTVbjRo6JdFh7TZsw8816K9MWOs7vDDUzuC3mQDrJoKiuMMg/kN
6M1Tm/mek/7zm9N3Dkiz7xuQJoYjkS4VpldstgtgMFn0AANuqOju3rw3UOJ/
uIX0Q1VmsXP3ORc7S5bo9H1vACvZT9DGV/0mNY4+63ESAIUPp+D8MT7byA25
Uzvb5x4j417Jp+vzLwXgiHv7PqFvyemp+tGQm2PR95cPrPbeMfMfls3Llt2e
3dVJ6ULWMRxibsQr0+QFO4+AtcSpGeSQV5LgW6EKMWiFh9Daxkp7qkYpCjQy
vyVMRffX8wAUYiz9m1ZQ7iMaYZaIgFGuuyRanAvKYLpDQTgR1VqtTXwSjj9t
UJHLniUKl4LXCW3xem65M3f8MwtnHThUSTtBj7cre6PEgZGcNUL612dX5K2m
Lm3Ch8ZfIJZx/Xb9PRvf0oQOhEepUw74kSLf3Czb0uDeLO8xZC5+sr9H4oGF
iogcXVTsTNTj8zUJRZrU/79tjD832w7oTICrnzBm3quwkWquplfrkri7aDRB
HBXFOuK4XEpJ1Uo8CSXSvO+QcE9joJDvCPiqn0ScS3wiGe1XRf9I1LLMcuYj
bWDYRPUfkvTcjx9Nf+/eQBykXoX1as6prg9+prmAusrfgr5UZ5l9IWCOlKCN
l5l0lfFjQkQsydeeRttv7qpduPH9e9D3wNNV/gih2+tFOCjxIsagR5WrqMi0
ubP3kUsa9L3UKUdG9LDh4LdsxmOAKaMDtN+I0l9RpClzs42KqHTbUzierb65
Pof8Xd/cJItIAdi4ZrxH7/K+5412nl4Io06zeZC7gz8ko+MrKB3BKy0Cc01z
mCIBxMRmrPyN5MlH2w+KKxmZ3UUCZ2GwFe/yTZlr2tJuQUCRAG06QhQe8Bxc
BkucaOrrfUexY4FpxdIO12dhKqw4R70rP9dyMkoAcEIO51oueIx1zLHsdqzM
Yxp4aGva18YYI/n43+4GzuSbX0AIrV2t0BjRdNRqkur+Jo8+7eiHZQiqpHpR
oBERZEu0cimjhCadBopovraNcQm6W7P1o1ginKaJoggzoxMBaByjuzlQFYon
1UhAj5mic45qsKReTgagGLyeZHffx+HuZNDxU9NXN31T7jMmY1GwL0n5XDfW
Y7CRPE7y0KaJWeb5ecIdlk7Q79PPDSwZ2YfkMPQXPV6drjCHyM9FHrOUZTxN
WUxSlbp9ysZ5kOOOWzQ4Ph9B2+7H/SI8dHIRkSL1HQoEEMXMVB0Uitswwg/u
2TCEZwSI2brr+V9KvVY4foDx6uWLZfBpohuNq6oLj1Cm4Ket14W0sYzfnhaN
b4oIX04tOa5WKVVBsvPsLqpypX/oiRUN/QX8fIrXZ7770dOa3erb2VzjfNuG
2fxK+wSygi2iPAAvI10RITXsk0NZ0kPpuN/pzANmzMPY3Uxbfun9BvIn17jP
TE9EBkb6Pc1rXJ6JhlRuuW5M2/yHFJJ/li7dqF8j6mqLHLOXcxwgeB6klQ6n
fsZ4bL0UVZTF+YXk7hXBGC0z4x1cTOFfni30RBxja3wdLQOu1ahaN3LE08QP
xgZBZHCTaUmDTZErROYe7T7SfXCnmBzKb4O6ZeIdgaRiooIu/7d7Jtnb/6P0
VW9heylEEH/Zku3pcLDeJOcIgHZG8rua3ZYiB2XJB85GFRYRRBcYXm/7FVbK
6hCn05lqdonLai5gvOYUgCCsG4wb8Tl5OLyyGqgt+DWsdcjhOMj4LH5M6HjE
ncyUjqzV2H4cbCIZVMYpoGSyNIWpufKJqkxIsKsobnaID6Jrki8PqIwcBPQ7
9jhZ1yhQXFdIL2pq3oSrvv07FpX637vhTCpizntKVwSDkYTnHjGQ1FRH4Op5
7yVAKEVp7yW72EnxgivX0yiJ+KyiDYjzX/6oH0+exiJBqF9LQRN120EYmK6z
0tcJs7VEXmplOn3QIruRLP0SQCJBA3nfYPw5I3byEuEDcD3Knn4hIbdcRmmN
ZTNdeq6eOU3l3gwnblYUdBvcjeSyLN8Rrr1If3p1gfRilKiZDeIGlTBtf0H7
k7jBkwc5bOjXrurGB8rSh6miR6EED9Nr+ZvmcHBjZ3Dy0YgWq8QvycAtOtp2
6bupLuHov/gDZq65qFkqI6T3JmZSP67JgTUTcGQdStCL0maxfA0ObnNMEysZ
rNqXZGYrybkthIRduV5zKe+ChhtAh6z4Wxu6Q5cXWw5VIgWnjboD/BuaKRJx
wByYy+Os35Es4NPKMGKeQ5cyL2lF22Bp2hMTBDzzZGHlHjGfmrlREL89YJxh
zVdXpAz3mkYoBeI0fLtMs4pJogNsuxu6vb0Z5OevKLSehcsuYLd9K0+W5xc3
PBaiTMPYhP7nJZqtYsJjpBVSkUg6Gz5a0Ywwv7kVnxNrp5Tj3PYCa0itVXbu
KZroVeQpftmK9k/JBWBOxrf7N5L0EsLhKisCC2epBF9df3X708A+iNfR04ZV
ewzigSdQQGM0fGZggPPC4HYtVQcpfkexV22mM6IDXg7uWq22cKwhY9iO6kV6
wCDDVbWxUzyePMnYG2tP1Q3+akOzLwc4zhsNroowvDDaCrRYY+2+51n2ArDv
9cuCE19dy6B9SlC62NUzJG7W9OluFWgyxrHg4NyuO6ItuBpaBCNvrqvGDwei
sboF27IbTGARvivb5UM+IrU9wAxcK50wbJxVHqpyyuko6Iicm9CFq3CWYusx
xnxuF0YL5wa14PVNXpLuzJJNw9/+wFOetgcfvACAQjl34CDJ9vAeKZUNOFfw
8O2pV7LqFGekozI0DKZ/Py4B8secQMj/7PphNTvbVLtjPEYLtSksCgguNSJO
WpTaTbG6e7ql4hed915salYFD8PDP/v9BVp3HQiYYla4Q32B372A04G4EkpJ
rG8xhxSCVXmGUJ7OoDUeE0tVcCeee0+pSD+urTyaELsVQ6jkyBYckBilTssC
L5Bp418V3ISez0jkhufHNvPalpvVRGxIoqt/Q11euroVsS//Xr7v1sBUaBPI
a2DiBqeSThbbTLUFs3Yg0vgzXneUJUfRZEZhmS9wKDjnl+GZOKcvp6qqdd/4
duzWLUHhPOw+8qwuAYRJVLjHNkaqSX2XvZJeQwsouO9HC12DHghTSMA1MF5U
F/IA86ty1uRvPUG7/eoCrOrFHm8ScO40GV5/Ui7uu5iUxMp2vBRLBu9K3uvV
4iB3ua6WpclGQMAdHPTVNzwIfqK74D/0dDhzNN9vGEfWu8C+TnZfG77fwEAX
dCDoriNXBaGQ44irxee4kyVZU+c+BFL+XLH9N4S8q91bDIuTep0ihvXm420Y
74dUavXjWvnwwkfWRT+21MA+4YnTRzvJXoE1e++gEkT4Y90Xf/k01wTUOsVr
E5565oxnfmaf1K5WbamTZjqFMfAuWiclCutbY+4d4sap0ql3ZCntcBJL20Mg
cLCaCKQyD4ORhleykoCfC5rq38juF8KjlEKXcaR38byYxkIIGQWuk0BdCYeh
v7vjcOzf0W0WHM+7Zj6H9ajirubINvRq6eN7c73cn7g/CdF92aHvnBzr1YZE
VVXlgezA+53ALNbhQgVa9MSJxId+oc4/Kxe8Vo0ONPv9pEkmYtIXa9h6CELF
q+Xo+WPEebXvOunz/svUeWniIHMJBT877hTYYU01RLKCVvbE7FoNo+p3OLyc
rIzLWGJ5dIlNq1rEuB8gG0k+3rGnamqfmLA6JJr1uBTfS8xmCDwHDv4RwV3+
xZfSL6+0/L6Hvp5OaqcCNQ5KD6DfBWWjpZg0yJ0gv6T4NknSiBGdQzUiYYUt
cDTY6OoVXeaeTXAbS9ScIGTAdCX33zI96eOSLSHDW5i3U3IkJ+aeEXXBoPnD
msUEW4VYLB/JiCFNxS5/1UkKf0RCm3+ZQcWB/2MPaVIgWY3vCTdEvjZ6mptN
mA+na5qnibp4cJeEYHjobur+Ho37Kuq9QxALCAfIW4GCpQTFBpPkc/6N3R0i
EDuWTXbGdBG3cGAwQef1r8x6271A8XH1R+ndVVDQwku7Pc5r2C6qwEXQE7lQ
JI61CkvCwUl7hPTfzLyLTLRn8nZD21q03vQPiGHdvfmBhJ8/6VRI7CseN9qC
WVJ2ZF7PTa8JnhOrKP1GayoeoLXd2SGObOKLCXJmfiwW2yYu88+G+1y3HOnD
RsTFC6l4X+T/9HWVNJx4tOxJAWgi/D/YoGda25OF0YmyRR51JnFHFsJ9CnYx
fjc2/u7KK45VBw/HFtH5ISkLDU5i8BM1dC9UZt1aNqkuQ5WL8mK1NOY1H1F+
mT1zvqEuun5Nx1GZ6wVpi939PTOMMP9ZO0GE+azOP5pCLDL8clz3prouHqfP
qqHhA48JSGw5KiNlavhUo72mPE6Ide41HkOaqV4n8iwf42i859y5OQt4uKKj
sHC3BQlymUu2S0P6GjZMWae2H0YutzTzp0CaMPGJbuD9hCImwqKQUeHVFTCL
y5+QYXoWXCml/NtJFr3irNuADsqbX1yQ90rn23s+kEUH4UR8Glva/2VepdZo
ZMmi1lEjYPecV/fi+57Sq3gyRUAnsrDdZvKpANwO5xLMhe1EtD72o3M23sTD
o4XKB1s+dSMpP70Z5mC6zZV6KPc4f02080FuWBey6O1TT3vHHMF8i2myZ32t
+gt+RBDUN/BoGBUySYAwutPUfwH/oSKQexFauLpfakEuEIIKnKQLzLiw/oT9
8YF+v4xTGzYS0lOuOPU9l6fXVBnlaKHjN69N0oCUzGMwj0EqSZ+FIllbNnZF
Dbpk45iTIZNDNkDiFqHYiM/6P4DLHTrWn9PxDD059gFH67S1TMUe1eP4j37W
qTbHO836oEnsW7CtpXFKizAFjyc6LuU3KDlM+d27u+LRXg6GWuPukkz3EHcn
bQjEo8FNZ0ba2u3gHH+Wuf1fcQ7VGnDUg5hyEAfQ/0hZzx51Is0gTgE1X4Ev
uFl1m7ID6X6a6LMQrv/9zp4zX+2lvNtXBC42Dh5jYGQn/olm3TIhtPfvAB88
80ZpzWy7sIJ18AXOft9+8Vc/9FFPO/u6gPSo3KAEsO6fk3c+AFf4EWAc06UQ
47VEeVz8poabBEyOdS+Yotnc8bQ2g2v8EUsD48gMGx/1fLxNspt5zIcXGkZL
RJTgwQK9OqlJMbMrcYnpmaAnLXUA18TNkNr13oMj9iByWbP7aTdwmeN7+Yat
7/5bWHixJx5BTdZ2lUQHuxvcgkHRqOTWzFkDjWGM9rgU4oc6qpE1sVAtvtwZ
uGGaugSzYBgCgDPc9aDI11MuWn/ZtYhMMdRraGYO3CzeEpkwksrjLjPO2hHh
tBAsQfGquGMs04J2SBcYiQsSYqdt4+dYmqc8X/cLNJQ5fiVJW5b8pQjbuhSG
Bq2+gDThHWcEDyk/0JQ25uCjQOjKd7u7WJjpXRTEdMOOl1vr7Dw2i8cYbt08
cHR9BRuxqTJgFcIfRwanIBFruQ2dqMVZaRsrZe11uMigFvJ0dtJQcF/6awpG
VtbFkxz1x3W3WrAg0ErNBor/s0u1YimvLFEtHLWmHFK/Wm81eMSGZRtlbfao
fUtLxqayRequEDAOetw9ENCj8Enu/Hrmi8gBAxoltNlasJnLTWPEo8CVXFJA
zYt35KPHOx4RkQLqL/z1jgQM1iFfCCyZMA12+zlGfR3ivl1/bi7RLBnf1l15
qoXvsEL9WXdpYnrf63Cef8NPWkt3Qnib/oBDJDS6gCROdLZaJCKEvwNhqm+j
9pAIWYRJ6oKtksp907GqUDJ0J4uLWEsCyOjuNB53Uy2vDC70fHdSEpPpMb98
mCeqSWjMTjMCcAi0YiiIj//sXDfiqAr0E5obxDMMgs3742LGjA74/omciX1L
VgwouhJShieC1WX8zUK+KAnQXWn3NEW0UUxjqHGWodGn7k2K4lNzhwrLgQ2Z
vLjgT/NBeb8IKDAq9zELA9LN+xFtmsiGbhXmK0cJlrb3SwAD5ct1OJL1Po+M
ZWIY1Pz/ZXaFjquSXkuN6wbXWLhpMhBO2cAh5hbuyhNBhZ9Hn6fLqw2hV6xe
H7I3s0eLqaYKqgVD5Zudckv1/+ru5lM60NjsMMixgfPBjIPqJz8qTcarIZtD
nrBDkXDoAu46i70nNm2dswP1ANzOKcF0SoA4NLbPY2KbCYbAFFrCGS4V9z1w
7K0yGkJCrICkNGbKlLtB0wj9jSjxkPXi9aJ0oOeWirgbnDPpC5Fup3TAeaNV
vQC6x98i1FWDhNH6kEThMD8CCNASCRj3CSTIBOuyzcG+XRqF1rpQSA/CWT5z
DvFS4Vp9813rSQm+s4BGfcBT8alQ4AO8JzCUfKZRrtGYz+caEFTvUyfYW6Eg
xZQKQloCVn6vVjnz1Ryq2ScxfpHP0OxM0AbYXqDrt9CrhZfJg11o1D6f0VXP
bu9no3ck8C2gGj1IZfiGN2QW2diQys5BoZb13jnI5iSDZflH0aHQ2LTn3qyf
X0e0CfMh0uMub/BQSwA0pcbCUoYaE0MxHMJGrJMoco0QIoWT4IA/Knhj6mpV
LCrcBgMJqkgjn6QxExBU4STUW5VBs/I2feP1Sw0OKR1+v3xkt8H27LEXn0CC
BUuhXPxXzN/+2JUAezsU9Dz5o4bEy7ZCTUYGQyTPf/s6LJbSljw5f7JAvSBF
QsrVfeMUMEwj+6TtD8Qb9z4Fe61oHwA72cX+wZLuAoucChpZiMoy3OfZcbK3
xPgCe2Z8Ltsie8bvb8B+enIdCdr3CLT7yRamB187un9rmrmKWxe3fNfrxMD3
tUo/Jav+BQYFPLPhHzumjLwomdUQ63n9dx8j/W6sF8nZPvIGRkoyawj7oRwZ
/fssQspfhpsVcE3d2FLwa16rsvL2WfIc1m7dc+Ld+Hx9Xpqv7650Qb3v4nEs
NJbkfuQ0saCLT4iX/YKPpyYIQ0oqkwT4xQEGLdNERPHvskOg6WwjXXwl4+dq
++syJ1or4u0rvoMvbB5zgFsES3IXFykPFWQbX90M2r1AwlfsiwQTcyYYEzv2
CGDmmECC4SRC3u+qCVb1EGKgkAJ7M/Hl3qLpex20PvqToY5ajdcnPiyn6E9t
pgeZKZkdHGP9Q9SB85GJqBLuElwAFRn85z0wfFGrnIqDn/MN6UmYs9bgdK3U
2N0pM2oM7w2Ku4oleg2w0zxGKElSP1QXWRkUHySLOknAQ4xs08WWwepW2iwR
sx8z8qEUIY6rDMnPkqKFRVBGQfFuEf1OYbqK1EAHUMYko87u/zUAvEYPA7dZ
FfbgsRe7w9PFvfI7qT/nCftOr1pIJVxj+fwNEUpbzD8rDlHzXoTpNZjpl+D9
i4k5DbPc/65I2J/YNoS9AZCVPmRJRLr9DXgDQ4nSx7/m0Wd50noijwDc2LVX
axXPM9w1Oefssh9id0hlI66far8jnAa/yHpIwGnKR2mgV4Kw12y0zG0WcOqc
3aAWXrwqkhzP9UNWwQGf17DnGtvOpJqc5U4mQJZ4qmMFl1QkoTQYOQaGCoTp
apaEqGkpDWOTAuLsC8fCmxLg9ZFS4HoWcgYAGITaO/Vqd0EO2AYDdWPmbKeb
wWBWC/qoQRc9bhfgcQJPYPtQad3BsIcaStPr00tGxoHI49FyJh+MwvmK8YMM
FOJfTcuWGEio24tMgJuwi/5ltAA0hIq6JmLJprHEvQ6RIiw3i35Se4vG0u/E
eF75He/om1HPV0yGV8s/Wn8zhTDR2gf3+eNIBHITR0WU032ZZZm2gF5el2oF
yvZ7Aar32zkZS5BeXQcT40z1wzTgLSRdcOQIQmPniAm8/76cpGKVNI3wfQIC
KsDUVhezuVtCIDiXQ9Z0iWJuAqjDdSFbRyQ0i0rIsDZNa/cM7CVtOsq4+lGt
2vDbYtzcsFv9a27Ljb6LxF5IhRpubWOG3PUq+hp4Hp6mu+u+iy+dlIcKFXDO
rrLPX6D28v034EpMZaNYlIBabvUcGQy1ZPLYEsF8enaXudAhxAw5yMzI9Rhw
xAJ85Xz4GYFXM36z/LSXRnk6VEbLy2qW8wIE+Z9sfi3p2yE7zpx8VdW+9PF/
JGOjebRm76Q31Ntqj6QMPMb6tkdsFAmBTpNYGO+kH6OGwjobIOHnCtThV3v8
imko6qs4SYZFdhfYkaIZIUiIxjv5xgrRWGDl6XAbVNIgSgG7UlJpocxO1yyc
COVNbMQtSpw4WVjiFx4lg+m4wr5dNOfAv1u6Snir6+XZRnIj0FwbvVGR9Vba
3w8P+8lInvQkqtUYqlnXwQXVOIdUnSPL8pPNZWkh5DGH5AI5rwaaYyey9DIC
/3X0gHX6Vc7QWhjaFT5faB3uDJ8/DCVjWpaibv/cLFUIJe2xeRX4KfvXzCnU
6r8nxu+ghfNzhy5BK4kctu16C3S7MHAdF1rFHvz2lHniAgNMboGVrCHGmAtK
D/vs/kHIBQUhx17u2B+1iSoskAjvw1bX/up4cbkKPutfJMAa6oFVtAOzDNPv
hhBgQMvUqc2h65hJJMrnKgfkrDOooouOebWfSSTkXO3ye8FrFdJYoGv5O9vp
73QM6qiXrpXSSq0jgnd7ijy/m+LhWK+SLbyMQq19PqL+2naY7HV5FA02zgyM
QftV1fZJMf9IR9wC3CQHkjRvC53EwYoIjQkqTzWehid1sMjn6W2YQK0dQVhm
7nyKghjPWcgP/yc9zhlxUgpFW4G3FA0SXEekSuMVrKWqIH0x8yt3WYqId+kP
ZNeNUA6c5LKmjs5nQK4TLxFJbCNK5y8DInVu1ddJcwwTLcVbrrn9x35T/n2l
h/Kye3YQjhq8Gq0MYVv3zCiMNhAT0EJuJymMhEuZ8OGXmOdB2ZjMiy+J0opD
Bs6t3Eon9Cq2rIWgG8K/BRiaPE2/7MxMPz4hMlNFOjrMT75sCarRspyg4LAi
ZIT0c/bY7Dy8pGvzbZT9BM2tBqQiVidtGK+C/33Y/McKcAO0D7AsAxvVwRIY
saQhwVaNT7aza8++uShvN2w2UZMP3bB6p8cOcDiwA57ikEQGUXGKmzU5Bu6O
kbjoVtvfQWLUkJvvvXwEUYUfFSgLW3REAwXgLLkZOW++gLbkcpnnm5NMB8tz
/98q22REhow5RnM/MNNwjY74iDKl+a+Oaxqy7YJsahc/kFTZHKU1Z+kGT32C
CQ+H5BqtPRXO0FTsRr/vYo4HIMMVmfJi70DhtanY3GDAEtWcJwwOimyPADYn
1L4Zqj3RPzlBgGBjDyHPKkNBlrAsJ+J2HNhJK7tG9/H9B4njYDx6vzb0xHba
OPPljmGOgUIxgoFKqfE6Kx7/EThApDGb0kDHMl++FWRSMq9Ila3+CV6LoaZV
Ash+7vFqImtd5sPErG8dyo/3ZoZwZXP+hwxzzl1jTq7J6lHDdGVfa13M2OSk
lVr7UbNYgEuc02ZMkCTakT7j3aI1rY9QT+B/vxHAVN32dVBvM3bnA+mTJQKv
bov4HN1Pmoc6Lort8ZrqZPWyDCqIMfSVCYOuPwyMNxZdLtObWRcbZ/YSKeCi
LfX2Fp1sW3Y3GvIOMZG72QxP9/EjdhO/9q7wZXq0WbnzyVIe5EaFN38USm1I
XgxUFIxYmIAzt+1FWWarifEGrIm28u3K116jW+QeDrEezJ2dawtK0mkiSS2h
b8Kc4V2VZg0yyN5HOcjlYc6Ho2sy9/VaRDsGnBkb5hxI0vlGlaZuNaYvIICQ
3D7No19lTko9gGbWi6D6iNRwXxZ/Qa/dxsDRFCoqygv91qWEbGKuPyn0QAs3
rIpHIccQ1T+3ylfngZzdD+ZflkwV1o+CqmnebN1jOOp0qeGhPJq/7zitjbtp
XiKY2Tnzujac6HZdt+XbWzTJSRRaoTgN/KPoo2en5sfosKpo9HlpvHOK0Rhg
WQMnqceV/WUkxEajEo5TatEJbEQjgpf3z9p+ceHwX9jTrBZCAJnYeDEEX7bG
DlNE+Z8FaNyPPACJWSJPfhm/V/TjEwg4HwaHoSbTy+f2dQqf1+jwiTzDZZj5
6fZh2Jz32vL2VrB41UgPVqueK27hTtsrLaiLk0jds2cPTnTN7UuRW0sCziR7
R2kWvf8whNqE5tjT7my9UirrtBgeBju5MBUp+uVXOjYyMB5tnq0Qt0DRh6k+
9Rs9C+uVcWA4sqz0wCE8N89a81nSJBO4Vi8TbjUYY+z6FoiPPMr/bz1eTJCO
s5YR+nD6dmSer/CM4cCkAx56Sop8jMS+VbAGdvq1iwBRHwOU83m9Njn0El21
rMJVms40Tp3fMj1ZZX4KOz9nRGduzKsRKkU1TifeQl2FOp7dBgRa9CwTrhyt
rQu/TzpWTjbtoJuWHNTi8bAYpztInlEwctJ9KsYBP071HUxzr/wdNVB+gdh/
T5uYGvNI5H6q4GVtRqYUXRO6aQ1MzOSMD5PH64FkfeZKQLE6uIVg+1Ta80QB
2iP/ynDJkwPpADMxXHwSo0vI8aMeFpT+THPrA1NNuuAADglkTEzNeWkvzo6L
r0cl2fYh2qgWhUQyN9MTEkk6je3s8mEpIEZTDQcIrNVHx/EdH8Uy4ET8yC5x
m872nE6Wy8QB7Uln86YR+h/JZKnRoaZ1ltcuG5BpMgqpKk+CBdV6HPky2nGI
U2PbNjaq9Jiu6akMGg9N6BgKWVfBt5NNHMlz/ymTi15b5Js8xvcK2IlDGxyT
EKkHVLkpdcVlwQ05GP783nhaEUqo3fi7p+7EssQhQoaEBo+5GVLV51ZPP59z
kSTYNGVvwbQBx4cFnxTONUsignKz2mRtyEsoZmZlZ09ZFJQigK2lzXuH8aDL
dVhEu9J1OsFNp/lNWn861TSO2PHrKzG7HVVXOTwTD2ujQ1+7Jx8iZ3oIb0Um
ksfIEJgREISVkv/YGARnnfFKSqYlU0gDOY5GLotmHkGLv4lpCaTIWbZ8XcrG
60Gsz1WodIu9fUw1QDwT32C/sJLBTUniWmQ2qQCItnX+ACKNwxOyX3CkaWin
VCI6gYRR1UtTVJOTwsNHraMqIQIl2lyMwuObXTG5X3m0e308SxjXB2tFK5pJ
FEqB0azzwujboZw40wN40S/ij20jlzUEh9d7kod0ehN3XiKi+AAm6r07Zu9x
7xfMrVIKKGHjrVuCSAnhUy+T+EochNt9l8XLKJcgJ9eI5U6plPQpFMW53BtK
w7p0ZlKz0EHR3dJUyaPJqeSpL929ai+6xfDldHxvKXHq140+gkVKDhRlLLl/
CFes1CDgVA7hHBiu7Txm87fG2BzX3WBU9Ybx5i36Ugpb3tIMtOgd0luTMPuw
1+7OOQyiQFaKOwZu7FMvwUT4LMcEAa9AeesBYZlRnTUTsrPCH40P82caKRrz
n9NTHKWwYjZ6k+KU7BODwXrMnQaEPWKqjK5eCnPj4iOHtOfgkn4X+ZcjyBT0
l+PGyMwuvUCJMwP7KiVTWKOr0V8rXIqwRCanjc3rfxvVER6Utu0ZGDgNnfEu
JrGYQpd5qFaNa4Gc9naur1wNdRSfBsyR1iF3xEYFfZs2hWzzlGRaY2z/K7oC
5Kw08ImIhxXWrg+jqHCg0BXGu2Ps8lKy/MR56ccoAnK+TLMpB5/i/aIVQfff
jZy7xao/ymKyW0rO9mAabe3qTYjxm1961FJFq2sKZxhIET5tJ/oR5N2QQu9O
R76gHlZNDcF1MPqOnTdT/Fh6AxJBq4oJi6nz4B+k+oJUfZnLgcOvV0mR1AEK
UIMpdB3vdOn4noIOfbpYN/Yn8nrDwZ8p+QogUGWb2ZXVXQoKuhqc4AB3HX49
S8NmJ3LsraCDsf2pH2aTK5vuC7UVGmx6ud7lr/BLt3Jiq66OAPGFXW7kGUre
7gFZ3B7j9OerCToACI0OuLaljrtjOUa7BAs/wxItZYYj+rCRay/1+qsKnWn1
ruds+xucF/XMeuF5VmD1NBVx4vzKKLLWkzuFuvs63EbboeGDsOwL/qHeLvJq
HZFXVkM0g5VARjuYIGZmpRAkFunuAtgV7AqfId9iPNHgMOyEuJ4oqW5fXM/v
l8clQ4qjnp1fZwUHtrGd/oT8FT51Bynss3mhpXmp3kjTQ1o48YD2IBmugqyR
Iqf3yz15YATni6F2rKxHf0sAX/V9kyi1rwwetKT+HF8GE6wXecUx5OPQSMgp
QP0wMTYE1wEKgQGoiZ1CUL3njXmwADzSj7RNnEgYL8a5zajtkKHLTdKC0d+n
cICol38rvL1taBRh8LuJsCRkuZiE43HRJyA8YiT14RYLqztoO1qWwcgru7NH
q/DHNz/Qi1c4rQu1/AfM0oUDmY2ys+SEnRoJZ0xTpCrQI5CGwEVR1SnS5eWO
X+TSRat3LzUfOfJS73wZfvekcqaJi30xTBWaUzVZB+uQW8kqcJFWTxSvYYr4
TOWJpUi0yOUXAW1YoBxGTt+CJHPlYY6ZlXzwaG2SCQwB5sRr+BWpmLGq9hwU
E5Qw28Si3tyLTC/qNRmALWzt/Axlnb/oidoOC5Nb7VGTysTtthQyA/qwWH5K
C5OBQh1vt/NrcsT1hT/7yAmKWjH6PkOKlaCO+nsQBk1ZPZFFmhJAuBEOVipw
cUH/RznHrX8qWPOLofNZCSEatuoEIClqDfjFXI80JI+jAdwsnD6+1BsVBhVJ
kbq7vl1LMBm9P7x3knbEa5lcHtXl6fY8Fx0h30IdGgLk+w3aES7X8JgZgoNb
HSndpp5LIP/tjRU34Bv+mRRqnqdLTSbo+OWvY/0ol8GVWCoj8Jt0c6FxttK+
N3c7SIwwTI7ylEiB40kbk+aSVfLoObCvRuY1RKUBP9j5rDnwimQSTZCaXsPd
hl+/3tMIiJJ6RchB7GWeeJtyGVIkcg/SnQAnIRmMKGAcr8nYK+AIrAKElkB5
9HcGxz9eL6rK/c2D5jo8fvEAZvU0FowmjslvOpoSVx+raLh6CdVn7oa/gktJ
5MXBK/+Wh4mvlcwqpOE7ekHqpxVMIMlBtBFmnivdK//ofMtbkzt9ZYBQWKAw
AkLqw8b+YpQ6xXADb/FM4tUgJEH5Wz5MdBoja+qVkOGC1hM5rs0xM69tTyiI
PjnUBdKpcn1fRD1KGX3D+sWczyIglJMEqK0NW0EfryGPt1DRqmQR+3muyHCW
lSYc9O8i+S62LnioZsM4o1RhPZN3dcC+jKzGDsAz9U/YvdjalFuJyTuQ83KU
+nqNseDCAm68UqLxndVBrKgGz89z5QnPWtbbyFWIk+C9sSsscso0EaFZp+EP
fxeRNUD0qQtsWCbCeifqc6NiYMD7RuV7Zs2hUIlcm6afpFNQAPlBIWThpHFV
CQeV5WB45csJCjyGQOQ5hIm5JWsboJADl1sUdQnM6ep8UVegSLslM7EmLPaj
972sjJFFyUCYUFI3LCLoZC90282ERKJ7ac96CQjFTJkxXA/qMGUraMwIJDjB
96zMautf4lv0L/GK/3rqQZJl2rVUNMB7WL0Us5fbDfpTi8iz1JtpEoM8GsnS
23cB0pPcz/TQhQvZ3nZyAoc5HXovr+EBL8JDBhgyLzjNlJqgGQgM5jZZcjM2
xtC+SF+h3C95lj7A4Xh2Al/tjIkbxc524ChSd1AEqf37SLKF9MvwKkqgoLkp
vOWJubSSxjzgMk+nilXoXjS8UQAqlUiluN8eOEZQOn8HmcAWNnfUc9UTvdRf
hMZTqr8i3bgZ0QJ1hVr7tJkbl0zQZ1RY8PaXTqTxJDAApEU+LpJebolgcCS3
w02aTtJr2ebU+z2WoCDcMvie2GtlhxGiGSHi0cwcNUmwdoNC+TbPYPln0guP
n5lRpzaOIBBv6/DsE41SD066sGpgZ4GFixk9exyURLFEfV7a+jp/dcUdDQ6v
dveffvVrHdcViU5nBl5TgForPrdCVYXtXadG7QLD91QiO3uWxdK2H4+tUDac
aO8WQ2oX7EVzvq7nRTgDzOBnnUPZfHNPD3WT/DskJfvUwLhjsVdf6tFugne6
mI1GGfQiiNkXz81uHnpjECrRx5EEQr+S63Qdl7EOQtCPO5XVSse3iMAJ7wfW
TuUgtx0XE2xGW/Cb2rEYKBtQYz0gV/klceus9DEFktO5Z412xz3OqIjIesGx
8YG16ahFStPbaZaLhT9nt7X/vSv9Ht3xrxD1z2/hP37dA6vDrufL4tKYidW7
tLo8PAHItxR1Hyzyq1ht3YDtUKZpp+MwfHiNc2u0KVYuQu4tRvd+RcbzydJw
pVM++jWOHAg2Am2nHnBC1ES2n/HiAtCVYCIeLH+4qeR8OS1HYvdxQVj1VY+x
GJZs0BHCdS0CFMb6MRoPtLCYQ29TyWaUXKEQpOJ1dBsau8xoKzSPO4Z/3zfN
cOrhtZjyQn4K1UIhBRn9LRYTBhFsN2wqNH1guaYivIdpE1pdKfItprU6LhWN
uSXXnGuLlBNyR3MKL+000JKb9/KnRYy6ihN/MBX1NHBoe7RRBNJgcJvuqlXO
IReTiKdldwF9ioSQIO0PAQOuw3g6eAS18QrV5bkOMNQvniIU04VTjQj9SLF7
2Ze3si03lkuIHrKPSnEfUTyFzKzJ4tq83w3iRW6dnS1FzUNiPD9WACvPIlp5
U7OSB4XVGRtPSvBasxAK1EJVVCvnd7923hKXl99M1X2l2KGhaeSy9p1OY1xt
NW1sUpiJx5r/CQ8aIrUUQlKp7REx6YFKLFjfcPIJndCuAlG1RPaQR+GCuFlH
v7CMfbRc+FuvxupDSB8/wcrqyjYpYiigMbVXIcR8nVQ7rBovpaJgJGKoh21Z
Lef1tsUvNjLc1fXtT4vrYoPjmmZLrs2X3mBwGdCY2ZRpOJWDFOJU64+DI4lX
K7MrHkaVPm4dXQin24pEOQCWkpx5tUx9h5cu0BOg38Q6KxHfvVa/nK2nuW8R
2YV/Yi9ebinz0odsnzDEcUHjWnohFh3N037jqxpeGVE2G4DOC1s9OHjxSNkF
gnjHZQ6I8conzPT/qrav9aSZeJsRpiCMfdjQEebPMRpdSXmeqiB7CMsW9f3B
hXjLp5AkaFuFP0y4ipV53QWNjjuMW74f+hgktVSx1OncTG28+11eP9TNhHnJ
TiViQC00q6tNQd4Z60f3PIr0pI7z9GsvDe4eTyx2fs2gB9/8NpqzjeHtYqz6
NqQsUlewIsmw0lih0Jj1JHrxHnG2RR3/nO8kuYZZ4hq60fjwn717JBQQaMGF
tuWcuK2CWy3e+NPjbxdTdSbMUmGEARU1ureSLy2vjUo9LdaHAIDwfOmalC9Y
JF1CYWA+qygDfqKQD4HEZRvBedl+TWruXibVM7mq/wFeu/UC/yc07TxrFQn6
NpKaJPIlKSVmpmhhnYIRow0BmDG0zkOulxbRu3JTIRvqGKLKj7FmhtVVJosw
dCg68YRQJse7gvTjhaOjKYnCOBedqK1n8FRXgvhinNTk3Rr6vzyxaBzK72rq
ROrGriOFk0p+MpgGpTdHUXLb04dT2kGw19c2HIuWGsIh9zLLfO4PsrytfEX/
McJ+YCqUNHbxuTRoN5SeBTDEx29u1KCwGQ+pdCl9fWZRL/GnDmWDYKiaSLhY
pLFLxzFj4+p9BcljWW9tZCzS3gVI93L5VixX5osa561rnK4wD9hrL3pxWxVg
Z9vV77ytJBLcLL9S4E4p3DWHOyBZjdJIh1l1+PaPRIzpSX1TyndhNRCdgz55
3C5XaEE3T+bhmYFPpJ7/c2kmVadfg4k/hHXSSrfDf57YpoKqAee3IwhzCx5s
uQcbUw4ouvAszkM2sGZ6wkP+meEw5J1YP7m6NozSOf+dG2FZGurF9nQeAzuA
7w9IBQGU27s90VB04fJSuipxb6ZoacLaTsa6d7i3TwccbTobqFN+wD9FNd66
FuOp0miYvfA693ReQ8hxnpv3gTWkoaGxCn/z/ZxvwMRTEdRk3pBbRPgIPPdM
hdGOfIPHM2gPcheShxcVr0SeLsX3548QTBiAVH0rsIhrt21pr2kHec1XlBMm
rFoqC2GTJKIsjZF17XBEUqlfx9KSx8L3YbBq74a2lGcFHFZBBQIKcMRPag2o
TgaYzVUBTMw5214oX9MMxbBfdIJCw/T3xG7ct6BR9kq2XUVyeuIcoUSq4ydh
Nz1uYndbKktzdOyXflzz25FjQ/hsb68SOAe4CkFWxP3xe2FleNWmQLHoeLO6
xfC67lxL9PRPUeAoUevyRrKiJgIZlAp7t5AYshegUm8OJKJEmMJw9qGWW9mY
O51al6eHEB5UV1VEqZG+NoC/U+sfnXuY40v42zElV1EaJt27kFc4b0jKU0bK
fp4lpUnIf2cLicohXcmOgdEO64DEDQuNxm6UilxF9EVVx/hdR1ymauygN/4w
9Lo/YKOFWWWotcyriLaRup385Rmjv28/4r61Toe6PjzWzonAl1nYMA4s21Y6
VkUBfLVCUs5lT3S39EVByoSiWeBajrDwLZauIsF4pCUjQ7mb5mkpITUooyEt
IYScKNuVUbQPP+9r5p/GOvL5NQyi/5myTLme1w1XcsdTCdTYan3XeiAwDdIK
R4T2eDkeaeCtR9ZLK9dcPE/b8YJ7Lp4Vey+Fjzhx4fz8/4ESVdQIgJGIbn9W
FUPUlssX92E3QJfGkFvXAA6erpevhJxpdeL0RwmpiDkU5LtEQGIf5zLUYqNg
3mtERqoV0gLAHm7nhBi7s4H1fvKQ6oVcHkhjNguiB0db8Lv6NdJMlYSaN/pe
9ydf6GzC+L8ES17Xniq1/TxkY7yg5Sg346wdcm1nWjBmHh7gstWKDg3dPcRT
ziuVLgegbbaCAN6h7DFmfXwIiiqGCj7z0icv0xC3QXE+XdLTq1BTN83Jr13I
4rpHISLZL+qzEko0C6Sf9M0HRFvyuTU1aJTcpji1b+69wWbjc9V4UcYhGT25
mYAVjGIeiaVWgLcVSJwkEXVAK6oPkYMfFw8LHWF9yDlQTFPwM1qhWA/p+XGc
889fu7NrokJb0S6oJB178y0AJoGj/qNSStPfwe9ihECWNlB8WDG+h5Fi+Zi3
mQO7a2ZqGSUnPXFsD7FT02iSAF80c5uFlAWhHIwo0q2d+hpanJeKH3YCIwkN
W4LHiCMmo1MTa5ue7bzw1IB01uDaaNfH2g7bPoyhQswgSvKRxviMHCSFImhY
T69ntIKb7VNVtb8aIwKVbZ9dhVb2rf2x983P86dOOfD+LLREMphvFvuZ61WT
EZpP/KpqhJ++Hng0R0YhhNcNOrVdqIF1IBTaQawsW89sRzX0uYpWiDcJ1F0Q
j7RJ6SFPow/jD6+SV96Hr3AgMz9ZxO4JbOHoQ5AZh+hT2pYnCVGH1CoIKNmR
Ktrcikq++MJfrAICnwhcGm+swvuUM13oQKcPU56wgqke8WeJFHo6aCaeZIEV
VK7do/88Q4JEPu3SMcqvaHZCBHXbIu3tldbGv/7oaWFbpRC9jnwt4tiKVIgB
reMKMXHhDXdf3vmgNmIwttDGAoElIoHHlHHWTmiyhnssLK7QDqG7J73AA/Ns
55zuOBl5f9eL80aTtfcW9KqWVqMEYccALvxC/LUtDrnsGgMCz2apJR1HmogQ
Pj5P7rvvTcgRdHDIzmC9Gh3L6nhwytnsVhi4jB7z2LxQ5bkIZiCwMfju3Thb
qwxBCtdGn+ueblRYYYxKhkX5uidRfIam42BbPJ+W8Sr3wwi/pgxmioY9KH5+
DxnUj5VKo66t5iwaZ1sOjOVS7ufjzdSo0OPYcXGATJq1ZNr1m3v7nuQz3OYY
uhFzR4+FolmrudqlgfqchOlNOEd51LXwLwTCKHmkb+XOmr2uhmtsrxENKmjj
/7GthDB0jKr3d0oPncHXu6yv8oFvtSc1zBWFHvBfuAWAGB9PRmbO+50EV5fQ
9ox3K/+t7lgRxO0NZl3Lb3i4NWuhdHlT2+Pyln52bHVobRx9ZQwo6WnWnyXv
rpSUxqolRLWIx4Uq/d4KQKGZARGt608YR+AeHW0plBKPXJKK5JXBwV8+IC14
R+j9xFw7PhOgb8FU2uEWK8pKAtWn7wg+A+PnCTXyse0v09ahOFOm31V5130M
yLFoccEc7EIwxkQjcDxklA200ldhP5Y7xmso+D1FaSqMDhIOveZ6kpxj/A45
lbUqocZ5u8wMpzNymTF+Bxgo/YONnJKkhxAs/a2DmXJZ15itBc+TZG2Gfo8Z
YPKGu2z46wea6BZ/3HysM/Vrd4Wyc7ZK/oQSImIunS1BFOnwSYds3kjQMEWd
kG28bjAh8iqOUmagO4BZ423yOP7+lZ0LEIufwJbYiVNGrvZVBAieevlIrmdo
+UhTVK6WQryhM3ECOIZyjWUAmh6Q7zuL/x3++1bU7d4YgL6hAcGSX90V89tY
wZiMtO74KhNTR7A1DI1Ss9MuSxnUNUqVpNkpHvyHZpdF0r3eTxUZjfWWqyXe
hpgBljlptoEPO3RFsgb5iH/PzNwDQ29sKd+iN/7yNvKXTOpgqznC9CJw4GOA
YzF0e03Gj0nNczni2SIjQu122TMjncvY9QjmMjkIXLj10y78J8bwKGeTrTWN
2GqkcGu74qcY/YTUYPVL/efMVH95dpJIlTGTjsBsgbju5zymCI3KFoQOc0HS
gE3YfRB/PcxLzvxWDnsImd6IqmIeCGTjr9I7J+PiWv3E0Px/QdevnougrDFi
QTSk96LOtbuDx9waDByvrpVNVj/DcZXNesrTzDpxBtd2iegx/b0/aW62iz/J
PsgApSgIfJt/GvEBZAfweAaeiiwYVFtQylJn4c/R2VDaSkJOEYcrONNBg3zH
w2JKSPPv/MztGQ3lv7zSVrQDN7EuHU0ogWlOICdpnPVjXOBDybojbwRSb95o
TtIkaNQpVAJEGzu1xxs8ZJs0OdserObxdtzc9wjwe8MpT2A6xXCX/D/UKcxT
3Ckqbx8FuUwrUozFsgGeCb2rk/R/NKZ2kmP2seaForcuJbmQpkqYNO9QLLPT
O75hnwquMKvESRNoh3DGUyor3RQkqKkl6ClrK4PAc5FFbF9pfUo46X9BWpre
1OiOEw1uUphDJGj/mTXu0Ja5lThd+Hn0KCDaI/x9Qbd+HmAgmFzfkLjZazec
QyRCEG1AVBbz4UQMtfK35am9KvYVl6GuLcLhw79pJy3qqDN6hEAHXY4+lkNJ
3nwoch7VmOJ5g5gPzj5E788sz8M+FabqGiBAqIpgmFPfJjgHmi/QjG2aEE1J
RpGj6d4tpHUqyyuqxk1xXg4o4aHKtRcjXqF4MMOF1jkfEUg0UMER43FtoaPD
OCGGbHkJeoEtiS8DuKEAWrBZVJN0ZUCgdm6EejiYjh9eiVnY9rTWGAp03D0z
zqbFgxOZv+uRlvrIlN7xT8bZ67ZS4yatFL2xKj7XuqLKCgVr7uLFSiOP3IRv
RLuvOSdMG1An1fBeNL4nO9ZTrEWK2tX28s/XCzI9D0OyDjFrzmLhBjoqI0hq
KcfAX6YFC2k4qC6rSw4mcjAl27OyWwaYYEiSQu6Ob86jxkSCQVkIwrrWxdFQ
B/MpDUHrEO800GxZy/sVWg+VmGEfnzrmqNF7QZhQeuXUw9ggiSxrdeMq8mw4
UPHnttp4RlJy2QCD/nHzyqLakix/JoPaRA7Gzj63gkQLFRszOXnISz3+t8lt
c2RMXWFW+ZPIeUEeXBZRPdS9V/f6XvMhrBdIqx93TXVcFTJGJIruSyajr5WC
JClGUsDMaV79o0SvLsOextPWVAsd4u+NTl3hfCj32LfmAhRyo576RGB7xEcy
9/UhNtDt7Ggwz8+OO2zqEYUeuz+HKbsfnSGt2soXLFtm18fdHsBWa/1b1tWF
MfXwOrAJMCKXA08dZxJshDb8x3iQEKux13WfnC6vIpRH2nSHi1N8I4Q1n8Rm
jWC7ucSVuNvUWCqn3503V2S6gMvY8JFkd3yEaQX4FfpWc/ZONTiuru7kOZ7S
8aQ4tGzcS+R4R4fSgGLFqyvq9JLF1jmjthOT22vOWDmCN012Bx8aT7ZqSudF
8m1MlKmg7Eefv7Gb4HNNG7lm98cGsV8X2U37q+R+MAoaQSMuXFMuzglxC2m2
59ZuDOeqLbQYOdXtCOrUgQmuaut8avogJvVx8URNDkuEOtE4O1pkj0esVaha
rulTRNik3IzRTOATgRLY8lBpa/mcVnFyrkmwhNObK70Rq0XSy8ytIDil6Nuy
tGE3LoOu9E6pHmFBJhG/FmQHdDb8UXNBIXRaTWR69e/HeiRltlj6yWX8c1TF
qIAH9DDc3GGTC7IP9bxsn1TsxRDUOOLH/5r6zMIjvOSYN2RZBxAUeniKhn6a
Ieq5DaFEdEDRwRSel8P87Qixyeq0TMTWzsyDxd0EfqXuT7Rt+aaZmyEgfI+Z
jOXu7RSxx7xcPW/hon1bCme5hHvZXOicHUx78fPAlKXE1fP0tF+avqGIC845
fTJ34DDKVYUaEdIamytl7SPNvQMCQSRdKiUhQxpu6Uq/sBoF+/gRARY5VyeN
GB/WjMlRRzYYs54/EAlsJ0PT6eO4x5RtwK0/ph1xOFMAcnNpMGxo0AfPo4HU
qNATTjc97clhJKymah/Hx4bLN9IScTaH630SZ6Y2svBrWdAb1aTYr6g09hjm
Wm9T64yxe7cbCeDT+1YA/O8A/+Mdpioyhv1fS10fIsCCUQPdVLj4CNe8Hv/Z
L/msYtqaEjN7C0lhfeB9g4MnKB65K4rp6RRwY28QT6ci8nWybt1L9jtJpE+p
hqKbTg8vQZGX6ZUtGamoeOOFjfYI7qhY8J5sVKXJzLDvo9kVo8fr/O3MMS/O
4GjXT8NoqjBVI7CQow6OsBxXLL5/N1wRbhm77HZfU/wBXn8AxE08dhjy0Txl
9kNbERUXCCNN8I0PIsTxc2seiv9Vsb9h9lMS8/mPltrVyxDWIL11np1uelGm
wgcA/TnPxJi4crOewyv1nsJRGZPq9HXJymPkz0/vkZk/hCp+/97SgvV9Kd9G
q2bZhdZ6wNm77Cz8oZSPtmFCLpZmy+wx4vttwYxb7RSPJgZhzxJWdnr9fa9+
SNZKXx3jgvtybGz0+gayANpP78x5c2BG8ntAJHuQzydzh+CXP3pHNjv3FPJ7
dB9qkbov0GBrGj4yiKhAqF3eENBabsm1sY34+Pg4aF4eVusi8N92f/CPQ8lW
u01aKz3e4g3hJnVGq4Tsj4/lBW3yg6uBllJUxehWJmv98Bm4DC6L/rwmc5pN
G4aGfV3NRvg/XXEgXm7NtEaZkPYVc60Sd6mQ7omk7Hif4jOAMOY3x8XxuodN
xHjgRwkpdNJptKDG+r5eJu0Ov42CKDOD4r3L69Z+QZYgfb3qnGO60F6DFZSm
LX6rW7FFHZgW9g/zZKgrkYrduNzMo2q4GL6ymF3x8PwRhL91bRLqk65xUwcU
SWA6aX52Rbq58v1qATt22O6gYf3dbNVxDQB3OIuQs3k1UYUPHmiA1fVFWgq4
FhdiRisNdv6mYiShH9JmWnY3UNj2dwZPpnGRvTlHqC6fxTFGOEdqX1CyV2I2
8NTsqMRSO982nYdAzbH9msgggmf67JwOEtqF9yilm4WGFbMtWJyaoYvp4nb5
v8o0U1eDp0jFTpgcoPJkf8ZfPR/CTwHzE4Bf0QJhOIAArnRkq7iwn0JG0qF1
O1qLu7Zuu5fsjMfpJOvSE2XG4z9MNE18bURKPdyHyFybh2GXI31TpwLjYaqz
uJDNv9WBUFhaLUuV/wUNAboxtB+OiD7PzopeNvGaE87F1OzK1QkY2zHJO/eQ
eEuRf8+IcwufTwTUCSpByTBn1CCdIlJByH6HU0AmMYrhSdPmCZ5ZxbdyXHpc
9TPWQWMFN+NpXDgCN5M+VjdBM+dhQtjS2muNJ2AVWx9qVDp8J2oBIHQNwa1r
qaFwxc0Psq+fm4RVHClFr2vmfDJaqzeeG7HaDldpm1rm2Q8MauGx2D9eOIlC
NKZiJOIh5sGpKZbv9s6pMNgYRcA59uofO5Ys7Ol8oraSPwkMq2gluqsScibK
/6DN/yVokjVu7iG6gY/2ljJ7ec3ZYc9XanONZKc0ls1FEtVxg/qwGpg5CRDS
hecPsOW4kKUJST0cPhN+5ZGlfbfBX6z1XzjzLJjhsE5tubtfwdm96jcIJ8xQ
s5OEZARMRdoYgsCcpCa5yz33Bguu9AoKfjXxAiq2EwznHCjerF8atFX+8zHj
Y/7MPtWchU7wg3DWVdKnzwXor62RGOAkDO0IqfxN+AUcIA/9b4O/Uj7SN3aB
zlbgQN3TJoUqdyrvzdiuzoGLTxnCQee2IO/8PZ37JvPSFRB3QR5GGfzuvOrZ
Kn0J+wo/F40OTq7cNxcCMwgQL9sZbcDOQ41xQt+byAjlSTcJmKpBkuw0ZEKR
adMTwlYSzX4XmpDK+wYRxWB0jQXNFc4baIsEj6kQm+b1AvgMVlbOAf/POgVj
U0yZNkUUFxxdozcSrxn9CKlGd/tnEWr7YN0ueU0Y7EAGQs4YUX3RszlBlKaj
fW/HYqZ+Iq7HluKoGXe7bjQRQwhwdMo20Yv2Y8w2h4FGGt5+v0x0uNaqF3Py
Yz6K9gCE3ouynYVyVYuwOYb0MGRi0jNdzD7+lnYZ0bazCIKDAnHjMb+q7So1
wZEptFakIeESEe8MD/tGt359qu//Wl35LR8RWXiVGCPiZgGKbqo9coiwpt6x
8hzhdOWib1rgsLVCfSKMko6ybhhSFruzckucdb4QEyyOVXATNOe/ZZ35NnIg
9rJMhi8xRRBP1vvR5Ry34pSFCKlUM7IKRekLaVzpQPeGk6c+gvVEmN0/YUao
fAaemESY4NtxKGpuE8VuHJVTU4u0uzrxKHD5qKyCG4wcHhc1VO0zLFpGnMWK
GgPM0++hEEitlvywrkIaA7P0V+kGgfQ2ZTj3yGPvKe+BfG3NRbJFXBwIxFOn
UYnSCajKjkcPUFLQ+O/oMRq8/ejRxQDSb4Y6tW/DTnfKYNS31I2chLP/rWW1
3psGEdLSy5iFQc2TXkvWlSfL4atiAqvWrXViTiYHlyas36OZEpm6yhD9TGKP
X5Zwd+CRCEcTNXt/kFYDW4r5Drf+BwoWUTPBECSdK0c1RrzsDyCLoGrdm8I3
9+lLTKuza5q5Y5IF2DLuDwtoILCuDnbZ2sGdEEPdMoq98j3qVVAo6kv9Q/k8
iifQTSbmNVtjGpZBvxULh0wiF1lLiN/b76ipO+cEJYWntAzWpI0D2KKdr0f9
4rPCiqECM+0bfTc0nCIzdaIvMUaNa3R/bIBMZv+vPGN0EHnpunZ/Wl5B6J/A
fNm4dYrQbpBsAPoaEi0ixMpef8QWRlq9IvBXTVSCQ2n+2ILIfQFHsEwC+3KB
hCghqsowBYFIwddlGTuQGGYKg/arM4JWQnfNBpXPY70uT9krtX/spjkujqCP
q3mpvkCuzk/4J15FdqETFUMrW8r/uz1HYLv1TzpzPm9/HLF8Sj1/QwqV4j81
/K+UhpyU9DWD1PBINLHZA/kxURSvkBTQVkgB/fXxzBwUrVDsekeomjRBnkIg
cqOqB0tGhnXGJVV9l+DwpeNOSQNj9ij/CSyEvetKIyy39XWRyxwUVqwCytu5
4AYjxmDNFkSAF6Q+2M1M26mRD9jGLfaXIdeyBryvW7D2uP8lMNBOJSHuww5u
Uk2+yB1InxOz2LGFhZTwwB3S91MbEtEXG3y8BBDU+sRtNpiwdhRuhj3inosB
H3MgYcPyEDuT5apa+Sj8p1YV9jovCbBsyNZlHZ2dGo8wsagKItQxzr+yq+t7
VZwVEjwvpOvAXjK6FYUBk130N9ZPyAJBQAJy21qjlxZ434LZtd4b44MO/NpA
n5dKP/3tFgNa2tSzWJSRsxObjPai/EgmOxRS+AdursDNFvn8vLA66O9UETbI
x0I8zrjOAPXItTMWlS6n7LpCelu8G13H4c8qhZ4oYrh8f9lfsh6xzWhGZdQ8
lo+diFaBwEp2baZZ4URtDxY8IXLH+IIBrmm1P4XYMKslQEMB0i7V9mAHRnrE
gMPpZJGm69Sxm9o2MK7oEn5otns+vTUX+1cdQWx5GpPB+hJ5PLD2Es7RJC9l
iFM7tCBF5BJVZ9bV3bO5bsZl4IBwrGzmTV6CKWm1XD48TZPSNYcWa8snDEqO
HcGm8VeslAkf0qc4BNloRwH8rCLKIyk6RItUKwqesfVV+2heymP4HbAQdGax
p8o/645Qwy4C819TPRGySBzkoH8QSjcBNmE2FoOfebEk0tZ1nWkGYmxAUK7B
q/On7KKH9CK6Y3jwp2vxfl1NrVvcZ/S6BFHJdc/h74Nyi+klHJdjaU64YzVS
hpnhubrRbmMIKiYeSPv1D0l/Itg7cOF/iuq383A9gECRng07O1qbTelyDqel
r7hugJvCH9V1UFPWvXJAvBd9325QrGOIDS2wFY9CfIWV3PdPmDYRfeW+uhg1
UeIYrgTTus3XRkckZ/KdM94QMfaUUl1otratIU4nAVvZabtrtiLLhg5AJYCt
tjs201VZjsgx8ShxyLtAXN772AvgVA17dzuPMMAkZUwiwjZpxAhL2NqD1Hbc
wzVxxJF34khaVtEH/cocQSQAEsPMzGF79OdE2JuOl8FecNjejji9bLABCrlq
V6qFbTAzoXI61tMT/BHQJh+dCGsSC2KBj7l36L5TkRUZQPg8Bqrk5+/WC70y
GafUyf1aKBy+RP+cgJgIYMzkjrWerydW2QZn2TSIIktkqC+QGC7VPhLMcnHm
o6E4dgRIH8KEebZ24JcZho89y6qHLURzZPlrCWYHaab4LZRI5Af/IqdL9dAy
Wlg1saWAXMe0AgkdPT8v+Fld9X6vTGlFBqAwO/1EMbVqew/DtMPjDVxJSAWi
a2FnCEfC1pE+01EW8QlsuaFWbu6MhMiQHRca3qZfKdtBV1kW8Y4SwlKguQs9
SCiH10KWv47irfwpgItMcAii3ug7BnZJmuLQ1agk9luWsyT+gafD9e2Hpu5N
r2ZujcXFHMujPviaxWmMIdjAWt40qOpzn/VunHm1XMuVE/Wj0U1zRsFdLh4/
loVEWcfc4JAg7F4dUj2srkUM6qhqTwZ5gPFjn5J2s2RrqB2Ef6mIzF97ia2c
DteiSBXIkA7AVUR9FWZ+QxlPpg0HUsApMxMNLurKNdfoMQJs7h8aLu5Ffdcv
1erVVRj7nSHvE2+/GYp4+hBCaQrplG4lBo7eJ1nfKw8/RShqIcYslHnDNhu6
WnMqyqxsgWoZNG5SYN2YRxn4hFQTMjuHpGCj1nkbU62lBut3/Meo1UvOBx97
YhAQJHTAFQU8o9WcXAuGKw7Gff1AXTmBsToSXDoG2smPRjZ8HYcZrE72ITDN
dZct+B58PHegqUKvMb46WTEQpy7A8fiOC3hfjdvDj430bOYPRMNG9UXDD9Ag
/bDLhLIaCmtTHYhxLv8MvaEr0wnwACqGysOAdsdDTQZDtlQmVBr1IRHP8yuQ
+06oS+1iKU+EUcE8xG6x64PWce6cmUigwT3GOgwS82y+yqK8VOJQG7voc+RK
Y2I9FQaSVKiZwdGjZV2LWhqUrZLGLEO0n8UPh+KeTgRzIf53S7dUxvccipWy
NbaChRe1uIIpy4bI/UA3G24gNQcstiHQuiJfZQscC4wXd96O4Vcw05/N56zp
fgO6nmJD/2BPMI2zCIk8WeEGfGYBTt6y5TLYtKrrMspBHFv7zQYtct78sd1S
/LVJ0+fs05cJuQMzqfsDsNaRRFYb9mQLNGHY49crRkWnJDIRLUcQ8Z9lCZM0
6iiSwcFpHdwLU6/oHw5vZegsa+vEiGvE01ao6RNpz62aiNj6NsGfbLO7dPKo
8YCu4X5IiodKFacYUxYxms8qHacPFvs0sgcm2tj5Skhukf4peOF27CFSl9ES
f27IGCXtQj8EIDbl0qY7OHlrWKUUv3ghd0dC6cp1GIOHxVZSg32l9UCYZmsd
+RNWXx+onC03qAyAa8DfZudnoP/hfiVPPmwXGiDw2uxwM0bdZE9E6fE7wgGU
Shyy5d1jyY/gcZW2oar4TCtU9ya9aMIxKO2fAe8iKdTPT47Q0uplnNU4sGdU
eoHgpg0KiBLAK8uUfNrzay7QEhAFXFcEycu2Y3+KyiEeB0j5M6kzZYNWUW9a
F+5ferecnFP48sF1DKcjI7QE4i/tOYauHt5Bj4pJkb/63egpcPJI2+aFSLwj
/bt43+2BvhFPUhZNeQE+nLj6HB7zb8JJyneSuYSKbHLcG6m934ZMI7KxQCha
ra6kOR35ECoSVG5hLFnyf1JO+yC3ZDViWt4jbILo+NIeRItG+HNCQ3FqOzKU
XevuTosPHF6ZwKgD9rAh3c0mpZYThWmgF4zZ1f4MfhjLvGPA4s8XfG2ab+Vf
FMaB/jarV2OxIVkSqu0H74fKUgUOPI3C2XqwAzCB2ftwxcRjmwamHvKlb2ve
vouWyA6m0EPX3vLnYVf1Iex2DVUHVURWmW1HZoLqaRdviIJAkLatOb1tkX07
zw9NuWn6TbWUWAp9JLc6EApFMQ1SrnO0cm9Wf0kM0VamV4oCLmJLzrB3+B8F
SlBZBj6sYM33ROrxPAtfOg/Elci7cf6x7wsvcChP2z0oCIW8UshX04Fph355
QTlh2iJC0QW/lOKQW/VOdUCFxO+nAscYH1Q3GglItY/WKatiSfM/NPp+pM01
vH5292buVbotrmxzfV0NVO16O8DJJD0jWAm1i4kP8OQ5uWqa79CVCn9OIj37
8yZahNdK9yaad9A0dBUODiYEDlKfrXegKhdfvWnPb9xJWMA6cl1eL/yCi5yW
GO4ZiFNfXle8dhEYausTkWwhk1CauRPFBd2hqb4qwR0mQh+DVa/4VqtBz//D
xWrpd9gr6qajRQomNoBBeyuIzBKXjO3MSlgqfYtxyiClO1sXcw8vPsNgw/PU
5UtloiWsOPpbtlLDvbV1trcyshGb8yxH+af9ECdB3yBgFeT7jTERlEupV9T/
uuiKt/Vu6/1sZSIwSZ+nGCazmOs5SEzArY82mR5ysK2PTF4JkYYoO9AEipq9
0mRAhsqee4YE0YackIbqdMZ6hlVCUbALJHpoHCwaoWwXQ+F1jccsy0S1Xxn4
hXk9xxSjhC9+Z2HJG0Bz9PmA2KOr0e8fBwBy0unlegVxqW1HSrSXIYA/4N07
kwYOuWb7m3BZ09YKmDtp2f6GgRKlJFuMbG5jzuBP44gMI5ogRuDJKoNkHdZT
JYZPjymyPx311Yc9MmVPIyOEgl/9NeumZGHSou7qT63m7oB0oU8dL2+pBKis
mSZFeXkq4vQ1fDdKSby4drQWDQWWnBQ56JrrFEjKHmjSDIjBsm+liLWVDEdM
DWIWeivl5AMOqZGbm+dHbQuy51SXLott1J8GdiOiavAsx9jdTzdXc4kUHX2j
VzbxEhEbvAtFQq/dDT9OcN9WQoFJiZz+kYSJzjIMBc7e1qccL9OBTLXlbL8a
DtPHSpOvO7RvJ6MGWWwX4c/mznhawDgfALLV6Bjdp/oic4mhZCbiQRCaHJ38
a1Ww4GI3lqB4HLdtrqaSmwfEi/uzYiKGDuJXMPA6MQpRwtGqjQEvD4hyM2X/
nvaj8XViV/NF/0vrcraVBPPaJF3r6rH5tOVXypFXCr+vw60+Ah7ZhukBmeYz
i0IJLx/i6Wx0SysPvyne6R1LqqhigqoVB51FrmUO78WlEP1/8OzwpCKp9t3K
o/fTivQW/qNH6K68VynVgJQP0lTiFoYYO2cVfX/skJqAl9fgUqZ7SSgsv3cN
zxBYdI33gf/+DUxaHWYj8bo0ZcubUxPxPI9fgJ+8hjdv8WDkPqdJNsgc/1Ry
IroGms8MQHgPoq8WVkMhU5QZ67Va7upsJPJtGa7nqeMAqyFA4cqqE4dVIl6x
VpxM4STaqxw2VHkFJxnSX02UZlp73D0bq/zhP4TPD2UbrGxIdvzi/f7gDbTY
8k0KgYMeE8UjJDTdBPhT0bpJGFLBjt5buXAlNhI0YjRR+dvu9lhAb4toWBE1
l86sJ/GbfFPmASl75ZC4VEumH2TfEUMuiBAw75UzAZerrT1ASt1SyddYqmnF
AeSCj/4fdqzYoPxmb4af51f7vHF/Gg6iGfppzxRHFMEL1e3lyg7KUQgokijY
zqRrStv57lGkazTM6OH6vI805bfsOr4IxnmUsiDjXcIBnMRP2RkfYiUfwUN9
yZQtuvnNOKk9L1GNISyPz0SH52LTEctjfpWyiClHi/oUpSJar7noxJ8xQpUf
9JcsMVfhfbvQ3IkpvYkhJ3xd5HRD8PoxWOt252h7Z0lx/KQ9713bwYLLn6Pa
d4QzYRA7hB4Lbm0S+Uo9JsVDoOZSvCLaH6mVsJllqgZspxs4HQks2H4mABd3
vd1/3lJPHRhXCZedFw1Anva5xn84cVaGizKxFC0jvgH0QlyEgSB18i2jr63q
jR2+SUoK+ETvcVxpUDy4uFnI84NUkXJcm9Ui+KZfAxqpDkurkXoZc5aW5Qge
PkoOZ7BK4M9CSyHjFlj3ULhFiwss/ktJNSwzDFz/86TjqpUde1yvTufal/1x
lySeBjL62KoWaDfUjz4cv5qvM2TJjd3sWtggAToqMBkoJ30zGkYHF4WnsRG2
ucfEMZ8bxPBJLZ4mrv+dotl6XcfGwtvd3uFrHi7drgO8KDCUEluLX1T9Su2t
gKqZQM8Whbw0CwGi+xB9eA61OJQCryvL/AHgje+O59WjZ35IxHX8dNjuc3jn
WHJdZ8sakOLzJ3pFIadfkaPbtBDmY5WqtWjTuE2zFMf9wsvqOPrClMduGHKD
ngzjTe7y5GNs1g20gmsjIpf29TDyiGO6Z444VW/fubR1J05dghTINqLZ6K0c
M5U4rpiQ+5MVveLr9SypYPe3EIqTLZhM4UK1dQo8qt6JR093BbBuNfcQKQN0
MK7bQiJ2R7zW/zBI3bG/N6LklAp0WaED49e6YZLOAu6oV0JWhpi6BUtzaDI1
n/0jtDMYz1c/33QwW7SN5ssqyBQryuYzZ+nCmfg74pwqWLl3l/1ZlnKCp7s0
yT9R8DcgB9JqNhACZ0wupjDWS7yT5PtgV5W2Nvc3aPYUQy8X3joEJhTHHMwA
+jnJf0NOXlxN0hZJIPLjgcgyegQLkv5rg3ii33lmGGHkS22sKohgNFOSQrBY
yEc2uDDZsdLXS9UV8OIp2SSFXPCgAGLYZDKyGvEzMh2D9hDNEGJNCbinvvCl
oloylrgjuKJ8OgTkVQndcgByMQ+V8qrT+eazIFb6tPDcwHXY4D26iAzC71y5
QiaVIPLMPH+zaDxn4DjLnJ2EcbvM7AOtPIuUIYldtW9fD9J1HnFDRbzAyN4U
HB5YBbLkhTCzU9aD9LMTDUSPaKks9RUDqmeyWE+xEbIG9kBw1VAU4R+9nYtE
Jh+z48GqpWa4gMDZUs2F989x8puDForRGdnMES3eXFdZQNlbe/OfKzOhO+hM
Va/f+bTSDDnuuPRThewYhANU29AKkL6fIBReTR8zEyvRdmTRWJf6Lgb8u7Xm
lMyaL1elHN9ICofwkWZbVE1IV4faAIrQQAO6qJ9436qERiJudb5fqsVAPeGp
V2X/WS6L1q3XuzXMmUxMpok28KnIjgrG8ip3AbcR8GBQSHJD2NptJZnxPn9X
FQb3y078zYFSHxahhyjFO8zzWlhkb8/P1UdEJvI3cEJVo7ufMjB297Q64o4o
SMYTpIQA6suWBw/6jH3LXNzIMWf+jv1e+8o8xef5kJ8lAMa5beKZh+AiSp+u
XfabQ67tH7dhsW+JyJOtnhlF2POTGvOJ638woKJ+vhzcpBo/RYxb6edvkXQI
aJvlb/SyoMhxNRpyxU6cJAf1tCVjrezg8DC+2HyMIgTvhJ31gXU6o5WtlxpN
oiTudruT40Hz74b/H+5yEtJZd51y3qkPxlZLFZPPUJeRQ610QD/RaDCdx+ae
yrXTSIYAoFN06ltxkD4K0osOTu1i6mhFgQl4CzbdbWo2m7Rhb0txBOk6yDaC
40OdV6EOcv79dm5TBazN7t5gQimXfj2xH/cpefdh4mO6maaj6pem8dP4fS8f
zMYcmHTqQ1ZxVAmWLo9uHIyXceXaTGwsl2G9SYKHdyowZnxgc9NAV/3PTi7h
KYDfP8SuEb0MZTQSdyU0DgJHGqY7uuUfMhg4NcPoi/27cX5IzISh2WYtfhLg
5lP/W1Tx/bgnSZuTYEJzno47oKb1xbYF1fcT3ZKYkxJP6V/axAsux+tAIIqo
xkW6IcxHeo2mGn2XiYhcWYM3oHWwOMz5tirkKMXcOdEf4DGKYMnFIm44tEJ3
vOWSJ8ilyYzTuymjKFIkcykkuHKKWtCWJQj5j3h87E7K/pv+jv9thGA8Z6lw
0S5V54kHu6i93bTA9SUPfNCtrf0PTCgna/qBogaddwjfGtgnjkU9LgdwD1Gn
VIUnlL81XgmO5esH9MSVjZWb1UM4edkwvjNSA/pDNBhxjLTDeyRwFhnBZceu
0dGtjx3k89GBZ1u8KWjseInwkS0dNIQ6mrLfhIhZoN5Q3AFcDufDQ6pbTHLP
y5HFPC2CuMd9kcnPd5Ao+SjgG1j1o/a4oOC+NE8Onh2AizwLOAXe351KI3nn
xiT94YBZAUoOfA26NjWWglWWticdhklXePaTqoalpK873F6JkQ7RVI729oh0
rqohz15L8eanBD5LOvcE/JtUfSvepWIZcSIGRbyiAmcAbPXSEhDhJFLGLyDP
hTe3z/PcUuFWqbXHHKXzln5wOCBXvmbdrV/W4wj3yrBvVpavslT1A8T3RrmJ
QgfK4dbUWe3TJB3ZMMi3OQgrx4Yw5w2v5UNq8z5vXo/4KNqWJgjQ/9eTndDS
XMOhhYzTGipGFFUw2jriuFHMDn4c1V3RCBIPZGxLG7yJRJDQYWPHSA8pOeL0
moxmXR/P2VKMcv+II5VEGs3Xvy0SIMDuODV9ihZ8ycDhjya3fLrdVpBRrK2d
+Ehqx3WDnvVakmxRkIsTlDcpET1itIAnh1eSsQ8xeoruDo8B9ZTJSLZPAOLU
X1xm8s6kTuZEeDvmXbgR386bN3/3Pnwdu+sJTIEnWw5nYe9ktvUfvWK6mdWs
TsZ+9tN8fHXYWio8zvsmkxb9ixXGbYrN+JKHU8iI911bL1S77dF+EoXFZLII
9AhoYPPkpdWP3lv942O1AClSTq3I2+z2MzO+NAMKKiLgk/71youKh+Ez4Czz
W42nFIxrmkBNb3A5l7LWGNwlYp8yhdh9QrBI2X4eqs0Qq+iq0tiJ/BjTIa+g
7DgtxxZZ5bi86rzgGMmA0J6QVw5x20FPd55RbCAxk1FvFMIgEj2HAVdehR/q
qoOnOK7uZpjXOFuj6xBlHWi7j2l+rmWHioTqIk8P6iNBrmKvqWU78qtRU1Yb
jzCR9Q63LteW20cfJzo66Gjr+gjj6FR6CNfyAWSiJVLdlh/x4R6MU/zjk0u3
Sk4Uh2oaHr4QkQQWWsdhVNa27LDEDFKpSNz/pe1E+B1lt+meIIKTOyXDUBFK
vV6qJo07nRr1006hnQfeMPlx2Fqm3fXojvF+u3KXB7fCnxZ1fFFRPx8iFW04
G2Jc5jXg5MwxQCVZH66xbbjpK7q0CfELclw+wugyby0zkQmi20Yb2U2IY77I
/LJ2qUBEbTF+4m7MgPqPUfBXtGKM6N4UISz+vuPcNK/67P+IgDHxFl/f1CWs
XdiH8ZpF2htU2vWqo8Mcc+7GyUogKuVbRQt5Ot/AQVryrSFZR6Mw/mz5O/1d
+S60piJf4viZSnPhf/hZJum/oxy9fYfLpsxi24B4WYM9DR13T6jbobcktFft
jsFcx9UejR5HqoMonO6iE2Ltv5uPjtVKbCJkBDlCovo+eOPh8CN2UYxN8gq5
AGcC4q+YbFfHlWzzt/975XuhbyHqEpSDMs7C2xHEzLMfdktIdWqBXLjnJoRy
jKbHbKwEPQb2nlk+nF1lICcqkQS1Zq06vgsFMsZ5DAwPfWiyd9qkBxEw+ej7
CVV1tCjCbVROwEfmggjfeYBne/HZ7Szv1LsOgZxN+5yCROSKUa62pTIZ0Zvr
WpmD8vmrgq8anuB01wRTVMUrJn4TdJdMWtQNDpKrJEmB1+yBgmg083OjgmPC
Ko2nf8799xEB8s6n71pYAgLNY4VMfxc9Gg2pEF1gBeQ3+DBMs/4pfRj0NX4q
uy/cj/djJ6Pt8DzhvyYf/6t2G3YFSd51bIE4ZPLA5s6qRVh/541wX/sdoi5y
a/Km+snvOoEA1mMCcVfNEt4QpInD0QI/kZ+uZ6w9TzIN6INgLQphPf/L3ujm
ezLdWKBRBpE2lfWPJl0bwaNt7q5lNMq9vWN33X4h0Xmuj0w75Qi41zN1/byK
6cdcA5GX8dGhRWHxuGk5fj9OUo/xef96WVBGlXMcdaBR+JR5I8Zu70olEMMN
fUtSTM1UFU2R20ba1MEY4TLd7GxzybD6pzyfb4c/FmJs18mjEG+BwRQpTpz/
/ZINfnNcqLgwdKGNTKbBG4OSlQk+pXOLqKD8PKfuuH5t+nAbt5lQxSpqlzaC
gs/IYpE+tYvWAcC1OOEf/om2DPFGq2akuaCzrsnmYw66V6D5RDTknzOP+Fbk
tzrr56pKCr2ueKyH/Fsqj73umJDuIFs5DaR3sJS6jBjx0kUEl2U7Lc+ztubJ
8q+MLMDEo2EXzkdGIs+lETUnG3Tp6rpmk+AbneVjRE30Z59ng7h5Uz9GrOkw
TwiHf4v0cDOJCYvMZIM/SxujPJ7lx2+hG1sEFmow0nzDejKySudzEIEScw7W
3bciR19ksljtUpAZhUAPos6OZpqSYdzdvGLJ8XPDYDR70CnP8Hzsj1aj+1f7
BDPVOTqk4ZVvYhue6Nt6dh/8g+MBXOb+BbJa7lr5f6ByyWqdieOcRGVCOKqC
FIys9vwB3OljbTd4k7ZFPz3VluNY+zirdiI5rzAZmqjG19ENy7sjiDC/DE6K
6sNuXgB3ohjR4H+4nTlo4o9FY/G/KnVZzDUvwriV5Wor9lfujCqY2/NPFz4s
7NHn9+TSm2aR78RJuHxo9kfEayZh74Lf/UbmeoHLlsXb5RZhDcDp09kwvkry
9FbshAe9VuiAQGZ0CLimIWNzGAtgXGLzQ7TLfG/zhz/eofG+ZNtKob4vN+iz
Qhuv7KRsyewFK1kRdLqP016Ran8hWOng1pW6EL09Rxz1vsygsf9M6Yz+ORGy
Q4zzEPIcMjSyeF2gUye+bZjIhtG2XCXlFK1ImmxbkuZULj2JvjuuiCAReTak
z6kG3O02g112I4dUjf0CDhu+e9wBzH9ZA1cEFDYjErFsS+kKRgOdmxCUD97E
1bN1Momt6MZGeWXs1JathzhzQtXe2A85VJcJmLK3RdqP3Yn4Li5xKF68Xx9T
YdO94PxSsdaL8XfEDLi3sX/LuPGVR66rh5LKsRqG1+JVN9jYw7DbMpZhyTBo
tPFL/rbeUylJWYmlZWvCWF4dEkqONGeoBhckobpLOApaXfj/kcsHnbORhqSg
Y+T4FJbh6AXpghCs92VzjZKon8l3buimJzlVapQEUQFJBmBT+4IuHksJqoKu
uRSc0nzNG1MjvSwjozXIdxLX/fZ3V5XnIbq8LwMK1YXIITfglKPsBmoNoMiV
lo13bifzUhlKrAlnJ13oQrFDrL5aPJKDRYwLzavOD+9IpgZbIfd6rDkIG2I8
/y9by4raDxktj/sROu/wRnnY+8KaR9E7lwpjNsIS0hkMKloAAfohakr3zJQO
wS9waLY3yoX0nrbFWvcotzOWtbakQYQ5ifBM2SpgJokSGXYOiuwk1UsglQko
E2xwf/RNSRxoKMdEJq91CCYnooefbP2/Fd/Twh5NNaNW3G5ZGDGspLcyaBJm
dEwNAdw67ZtcmGlyUMArewQd39brwkaeJSRe2/9ICkZh6Tu4xW70u8wnrNQ2
Km3p7XeSdTPDBeHTrJrTosY7DaxrGH6efZNeAFdZRbV2yr1NTZMKWO3U1PQt
bc+gHF61hUwdQ8Mh9DYbl0uWLI30U/p0HO6NmSCmAUNzbGXVluXN2nY9icR6
xSgqB8TSpuJrUFQ2whkLhrT5LKRlSFoq10baJ012l7e/PuzK/44+BYy9T9tm
PQWPGuzFIlsO4dYJjeAw6a7uqxbmuKqBL/hXs3XT+OD8JcMhGBMr+jRAFPrM
h61SbnQwuANY7s5/8ivKsdLE04Qh9C22tU+hoS2NfCakIlK756xLvJrkZKfR
HRHs0OeHPEjswGoxP9GHa+4jWhaoHMECwEFSPzPcSJhRuVhPlFHy00c8R0K0
79TqIbJGvlznkItRrcJsmIDq/0UwYJJ/45lMp3dT14jx9v5DZKXsBQ+4Ucs/
tILcUHDifnNa8Xp0AF3ijk+r49sX1HWBFl1V+4jCj67KiFO1dme5Lrg22pgD
THLEVsyhaB/SzIgtRgoHOkwRci2ubogAfyBGnavjkZpAQKAAZZwPAwBnC8/C
7VBA0+la1L9oO+5ed5+HmOMVboy5Jaknma2RGWqaDBtpb8TvcJkIrQFAF+gO
sWvXCxp0IwR2FKPG/iUfHLwB6MW3E0IEwisj+h3I656EmV8xk72JbPN8fxEH
KjgpFJ3BO1kstSjbRfmSwJjgbqkLFzPD3SW0SelCNRsd5fgmuKdkgO9G6VBI
jb3VreCMGipkCdeyGJn71xN6tjKCMj7aSYAXSQcxPPqZtM7/hXQzfRFIVzR7
EPP18SDCFK/nMa76fOx4uAR+mWjHBsUHZv234V27Yq3hwz7oPxEgJaMxKQgw
0WRY9PmiXep6yUZCYUwZTP+BCcqCTXrwV/z0YfSsI5+HCZiYRPXWYvnhQYi/
daflFsFyFdfm+oQ0cCf9zOlBQ+L02UhdCTeGff/uKBpOa6hFEXXTMKn9jFOY
1l77oatbhJzGm6Ns9lmvKXWWRK0xmzSTqkyJsbo9mpB6qscAL0m2ZXnbsD7M
8bX+y5O3jQJ9bCwNRINL6Eo/ajFo79oZMxBV7xONnupqN9cC8j6BhWoRD5ts
QZGOIATGbru6m0fwpAkJEE0VZRB/1omJHqnAjE+vlGQCfkIlmf3iRih7/yLN
2sql67Yo1Qw44o39OGnlKXyag5LMAPHRozYdoC5WRtIaAkM1HZv9Y5NTozr3
wwfbAnDeu39W7/+UFUle/xC2MvOaxiYhJSy6Xz6UdgxnIxY9gLl36plruWvC
mk223EqM4y+GtffMRtYWIcOszNIAo8zgi8WT8QFlRd2fBqv3Y6PJ5Msn+b+m
lAH193fqLu1n6a+QsxAYPoJvhIHAh7Igh6jTEoY6tiHOxH1GBWhcqzCss1i1
zsYaDnSKarxjqQcIzEIUotHbTdC71Ic+jgYcU9pa4coa5lxqld4YBfV4Hq5/
/zF9X+LjooQLrsCWaH1SeqK+GgEa0vsAMAqYVYFMJclS6MTZenKOOYJU4MOf
33j43jKNKXNjHn/RTlYdEhmz8AC1dfgGCtoT77q2xzw93JvsWWNSOKSixmi6
zwi0tbOCbr8WI/Td40tqtO5a/NJi86WhzciNYpFTmIvQiZCGab6JURYoPxcS
+qnOSPJQrOVpLlBGWu1+L8eNXbzReri0QOl1ghdcxpDU+RovrYhNq/3TIqIp
tY4rt1ISdbBXS9SdCDgQGDiN3da1Ln86RJj5dZ50cvmB2NG6x/8kLKRBhdqJ
O5jRnUwZAe62/bY18eFtcMxH/07UGBlBp+6CPRnEUX4t4zKJInvzAzwMEEoV
kl1dL3WFuiYU0H2pjK7WUfJyFbfOsvfvtBIRtxZOuYUyZEsT9mvGcXW8pake
ixIj7j1BpQ7SYqiuSX2FocTzzM5JVBhZT08yLp6fFvWGOFJWoMlNGqZ4d6Sb
z737H0beU91ov3KFe/xDMOTeeHQ9hlXWsP4QfHSVhsi5Za54idVtbG82Xsq/
tZvAm4YwDspHrUvmv/WZ+KxSkjvh1G4lXOV9y8WI+ws7p1N+uslsInnjaTvY
ZNytnAAY2XVHmbguBsQg2MM66B8x087F3sLF2iDygrjLwKHwPkXA/b5Po9+K
DoK8ZXejdhU4G/nptkRhK6ZjA1TWM5TQ76szyFhvVn0ik2THkuwLdTtvYud3
t7Cd2HF3Yos89CMXrI7UTmcSU6BM15EwCJsAPXSngCHRhO/Mc+Dtowd6HuTF
Y2ln+wAjjlc/qLGUBZVhsi67tM43a3arqT370OC1JUQpkVrpWdT+7YXihUs6
uPzM6VyX+jXg/3FqDXfJr2uI2OPH/5/zc9ofqmSEliCnbS8OF3nbfwoNMDrJ
/WpEpWIF3dQvlQVKl/Swlaxvp/x4jPN9olTB2AkykQhzLzeGTbz1MPp4+HUn
srmQReGCHdnTnVPMJTE4V0CCJmr1skzwai47oPL9GKsfgZUYkXWHOCGnIrAA
ZBRbwratIPs2t/klxsOwSyquZ7XQ39zayfvvtnl4KUB85RHIOFG/REQkDRlc
l3ukOw633wXlUTLc7OKHaUF74Oeuwip557fqTo1V2Y3540w/69FEWaQ1gK6S
LgDMIRIWghsGMBPMzqTli3SLMesYRR6nHN6wJZY1b417EXcrUkILZ4PT1Yj8
B6cxk54Rw6sxnRc3/H0U64scgXZYIHS1sXAtEzxKdnEfaqiE8UIkpTfyxZsG
IHoo8ta9ezXtCyBKrHpohYDEB2NZs5gUNZGaNxFCsd+2TUaBQLgNGU0TmRsh
VbwwUOa4cfsb1svq/s1+JGgm85mviMUwXkVSN94rEHLQHFbjRlH9hvEIOBCX
Yv/1ta9ZOTNkWmnSLTQrlcNW9IsSWyXDlV25Ayikz1TivHmHSTQDVN8c9m01
b8/BItqF73mJnNzgeLel63cbsStngkU/muTADiQGxJqxS4mAjVfh73WYAj/i
x3/m4Vz1u8s0OTil8lD7atStstXkoS3e+yn9Z1LfHrNBsdfzxsawrpkaRU1v
ohiosuCKA5mwh8gYKuvgESLij3tOh8mSLG76I7g5C9hyk5ZH4tN1ZozphuIy
L12zJqi1nE3GJ3BJk6mpZR4U0AnRkHGGTricNVs43IdrJEy0To5U96dehVq+
T0J3eNNgJ+GKzGiQRvt2b+s2FG5fWdfUtTCRSJFr+lRrXjCmJYfipePd4rA4
ZeQDELEX6MQ1qKg9zrDOWq+eXLiKrw+bty5FDfgxvIsnmJJ8iGRTGCivyTYF
ZsJTWrglu21OBCqUhx0rPO/CfM2aJxtcnU5Jev8vWt61TefWuJknI1WVXEyu
WEKrFxlmQhj2Vevhl8y1N0jNaol/A14aOoc0sPiRX3I5Jn6T+G9wPtOip8tw
aVGlVEbIV8HGcr/EiKMcbAckKs8ttsnghVnDBoPozgh28PRYN7TqZYGdy7XO
ObgAYBL67ByWM4tOz96nMrKI64P3gQsXI9Hlu6c0uk+U1dZcHVTkxLChkpUh
dUvYgcmSkP9KzRujdvc+U7Rfle7rLZAZ9l/wNRFr9L+KQihzg8KLVBbHKdRb
RhzU6DUJ1bZH31Zi9UmFWpUbYzxvLQOkWxehNAlwTyv4Tff3MWwwOjpbdKZS
/XK6OGFMvif0PbAqGiHM7ewmgck/zzcF53+UAC+ytT22xfoyWdkA3Rf9Y638
G5SxrEB6lTTtQHrJV/Cu/EViWYZapFHa4MKiMt0iYlHD/Czx7gakUCdMf3jz
trZE10/dwOUznu3G+Uikm4Yimey8/i/oPLrXQNSy0NVPzaM6t4wWJyov/zQa
NNh8JCOlVGDT7xNQ9pmPzpnI11VFSHuFqnrkkOe0IlvO+4OA8BLiUAbPkk54
fFkJo91koMELQcb9E86ypN8o1X6pVngVsAFVP8pJ/BDwfRH1i96YjcRwP7Cw
vPpJLrvIZnKriCfpjaYPmqfd7kZGL1MoISpS9V1xazgwJCvLj5ZgJgc+3O7w
dzXYoJvcQCZEiBNfmz8OzMMSbbB/hewtc9AKw65dd81PEptmTQEa6ejB1Dfn
HhLQi+ZyvS6brG/SstrkVFLaslvUKMouErcRtIzhSEiU0CLujqtpP2R6aoRq
iF7U/m3mSpxUuAC4PX4qS7kvnnGCVf2MWnvXZMxpx9lyCYhVZEMtMkK9AXZw
1LfIi4xe04Cpsqm3vFqTHULIoglUdCBMsbJjjf8ehvH1PskTuhIH3Af1juQx
g3SPbiPP+H9j+uD7+ocxj8y/7NF32Gedhtt/E+cWdzwc717F4alKHoCTYjYp
epp6RFlYqBYryYSBwHhr/HPmoPxqi/MsdmpCx3vJRnh40QZmpUWg99+ale3R
xRgCJMZ/yOZNp/RO3/ohShEJgeGGExDlTlr4COj1Dbwu9yg//5XCm6rFmlyQ
SyI0F+7pKJUHsxW0PXAxuO86RQkqGLbdlpvPGlkj+yE4+zDpnXl9Oeia+cdt
BK/loz+PE3Ko9dNMt4MhiI5RDLzAIxmKXJXM/KW9rIxqtTiDLPfRRkQDvW07
BtfjEJdXGz0SiuK1+Y+S72ubqRP1zeu1vLCaKRKjLeQQVKV6/Kmj5wzY+f+S
RPR9xmzN3PvSHcJC+qUkoVqQ2+GRVExfzYPlW3YGMDOR8fgoA6d1a5tWQRSk
EumkM9qTw/4YQt9ffZFea4aw12wzrbpm4ydsZnpA1porFAhxxbTmha5Z+n/3
92TM9+wpFEzYSQBHUCp0/RIwACeL9IkmpMMW/08F9UL+Kv55j2uQGiZN1gXo
fnP/Ti1WWw4AMnUlxiHqEYxmH/xnqS5nc05KjdF/rNU5fMz5OT8JhtIkVmIo
nO+xGEShb38yQrjHEN+64vlzGBmUE3e+mjamq1BXdpVvS7wYGwnxbkqfGCN2
z0tldL/en6ZSjWKsEpFAHMTCSDO0YLl3OJRfcB+zeXMkFdYwtRP+4d5Wjsly
PwIRaEkS2xcAm7zSYfkXUQibIuz+umumYK9ILpDCPbgEhf1KP07UcP66PdII
JA+sNTJjy8Xl8H+Itf8i7sU5rn8FvmLk1OOX7WWODKsPv3onoj/gZ7u6LI0o
9ITSLJ7NMruptfgpH4hS0sSHsCoZgHlvG6vD26HO0sWYxbrR9b+9TTgDYtdU
HhI9OhdmXEkAZNYQx+RKcUNj6E6tyWMhiuE52ttGCBfgoVr7Vx8p0g66IILf
duRg7y7yzpDb2a26uWbpwMjdAcxli3Xuyj9g7Xzg4HVibEyWoY1G+mkmljqJ
oYptsllsIZyBkhAKoUhSAcqB8O04+/8fG9wA4YfXff3U/XIljipUVSYcw+vX
diZOm3PrEGvoT/SUox7pJEEC49O9fZIHa7WWNaKzlET/r+sSxXlYVgeV03Ew
zrvkcwvirJR6xH62xV/PnTu7DtaNOsFVtUqrG5811NDktR10Lsw/fdjLFQk8
fkOdvM2fkNE1vXO9oKpVjXq8+jqvKfcUqpfawEF4E+mdBoSscUKH0Wu1k1An
BXr5STzwGuyU1lZcLIuqiPE+22rmGxR2Y6VYBbJMrDKhj/BRHTDG0XnLSFe2
gYMchoJHi0F2sPH6/4Huqon2jyMbzo69OCLjFcxLVUzb2nFTwwQTTsDMREON
0SF+uXj+ClkTSuwLco9UMBj3Mci6ue6t2nqltoNslxOZg0hPn911IoJt/oMl
TnhDq02tpcm4m8Gvn78qMJL6aA+fDOGmP3qSUMe3cbXeVWxTYg9fR5+VXQbQ
GWTWkPIEmt5K4XazC8WeTSbzaWOFn/EVjFB0m0xIzsyxDVHBK03fLs+DMfXx
GBZsrveu+j+smomBrzPuMBwlYYaoMDNDgvPzbWmy1HWQvob8CLAfuy5xi6ZY
w6xCeLDUlwofOdrNTB1uqTt9+Fx4VCvn77Oov0JHRQUo9oh8NLFF0gNY+6Hl
U1k/u+7WpUB2Sqq1TbynfjXUOn4ogGX8gyftV0/e/WdHdDmNZvk2+fm5+UfU
RbVorKa52oNPt7TM0gyz0JpD7oQbQCw8Krw52eaCMh9aVg+AlBXW4xYnKiV+
BF7N0muImNqlxiQdUGVVCK2bldlmQZyktC5gtsEJsLFQ831DaMlVATkTdIZW
pegZJrpOjU0Wb/rO5muAoZo9gWrzi1I+yR+xJGDp62OYELRONexOys7iDNSf
dKbZ4xQ30IB75ioqKJ13PVjg49w37HBiX05hguSXvKG3LOAKxiwnpYn+bV+b
fXkJgVZ0Lp3cAk8emo3DN1KCoBgYet1KRHyQBW4TgldNWbKn4iQ1oCsP0B6p
O4idkc2ldP6B0dhnU710SkHxkPUQ119+9bI44u9xd7rZGN0xYaBzw9foExxc
Vb2KWHDOHw27h45NcwZe4X8LLP05k+LfqQGjSxNmwxBKDskB0PRL9OaJw5Qe
sJumndlgUyTRclZlSTbcxWylajylYW2Xejs/DxNQTEz+efKY907Y0grQW2aS
E3RFpPkzB4kBRHEH9InCfnugEvndWJaQvyLT34X/qVvg0kJElXKkFR2gdaHP
TjyVVLvmD0hao7UXaEpdsOxdwOTmfsgQotJalb1/xWA+n46t1SnQKS7LwOeF
Y7JT4XixCuKnOXohgJk9Wcf78z8QbJLN9SAS5z/is0RnDTpYEIjDqiZ+JUMn
vxksT6U3UJG7fLNTTuexj536BpAni2tbPrykwf/qfgvCFXo+yv4WXLiC5oFj
39QJg1z4Zs0ghHc2TdEfoDz+T3Ys3ZiriXp3Q6TSUC54LnSCypKfu1jtpCLX
oHoLR8csnT+p6R7olvqP4ojCbyi6i/P2m/hnkThwfAfx6vsdUkjlCsbx4QHN
1XsA9kHIrBK2ZCW/3mn/Ydbbcry3YYOHjcs4/ycel9Qzt/z9587EjISmmGyw
lRNw8ybuCnlcXcOh2WAFixMbBDZTrEMfyQ7wmY2D3sF449+ZDweyq5P/IfRz
KTjB1xWvEtIC7ECK2qOLYBdGJd/k2xd/S9lPG3+o8ysHXKJhTzGAtExJjSEs
suxOhGQx5d1fgBnK8XkMhgr6JiwSIovQlbWZa1j5cIeon0A3boB76f4f+7/E
DtcDXjpfYgvWwNyEzUOtWjakJ6/S8R5DndBfRKSCGAOlgdoL2JlbHNO3LGeC
3bXzuT6/Cr3se8FbrgaXiSSWFGbG8CqkmIN+A6TBaWoOVt9/Sr7CQdootCh/
jdgV/2Zv+VzuCH7vpHHeIz7WETk122fSA+jDddY5ChChvj9xFtgxcMkHl6oh
yZifq59rPA2rXmXWx2v2jCmzLJpHGgoFJeq4OLpfP3c2J3kSBcGfwxXIyYaS
6AENVFifYrDBaUqiLPLa5qvac5bJa1m1XBkdQA028GSs4qbfc+UN+EqVORU0
wn5xjQsYQ/XkdfNxc/bzRlhku/aJ4CYctvS1akJGbuzGI0qxODyXwkJUlmQW
oO0pUchX4ty/Ct2ls2v+kLkjxsaGxIX13xi8EPDuH9UFliU1ryBgyCt0ainH
NZaZlDxH7fofCbJnyEYlL87BMwN65bjAdr3XSU45O4qlp1TaMT1NgYdJpwC+
/XrYJlb82gOblp9bCokYtM20LLURUVxPx/T+RcCgJwKPh/2EsFhz/Uo1cW7p
1nBDDDVNvcABK4iCcL+wDjAe+XF2OmtLdMK1BtrEMDDmTPD0yrGj/O6VkNBx
JK76XT+pDPga4AJBTwJZhJpEWMVrCbr11we2mTwn9P2IF0PaPz0q5G7HozIC
prmUoUosdSOZ521m4nWKqaeGUoGg60rIMU1vmDhd3E69vK6RObgvW7y6CT9i
DsF5cJwMrkQnmkb+qGkF14T6dpsnqU4fpZKrbgIxX5TtdR2sHJTAmGgs3pMN
mw6Y5XIyG8IdOzffPpVBwtUqA1xuwkKX6tcTZg6CfxZk2GTDht6IU89UMKzg
otR0iwqcfFYRc/+RQXQv5UTwl82/uqJN0lzParYQ6wcd+HM8iBOhHiSjtNkG
3rc/E9xs3n+26C0NxHRPJNpmi5UwBfwwyTzcBiJjVYXrE4WNvMIlvOyU4i/L
dYRPb1QIbN50gsCRMREAkl4C59z/HEHwt7TE1ZdF/rCTKauYPvOnkcwz7PL1
LH40tEpMchPFRN/18wX//Jb3+G+XDuJYbpdIV0ALB3Dd7SxW9jKvBkkRM1le
SSZ9aPczd9Hxgx936+rknHQ7YRf6nJi0DPA5Fnhyi1lYYBEpVl9DPpvJsfos
lltF/pV17W/rl4Maie3CQUA/F7xnQZBltUxxN9HtoJsJ6z3px4kI+/6ZmgiC
IbtFykHTidfk4L0GafPuGHwWR5rWpl2hrMYkJ1Iy2668+vKZfwxPXlGt1I1X
OZheqtH2UdvpX4eNTYJ+4uTzCXlNmi5Hmw7xVdAIGHMeYBvt2bOnDYuKS18F
Pq7bro5MHY6d/bLDgyz4MCO82Q2u8nS+39E8KqBeRdM0ZH+xEG2q/nqBlydF
zHEV1LKyEzo4qkfrRm1ePNCgP1MDJ9DSZGBi5/bWU9gI2lD0VVBgHMxxhfo2
+qinFtODUu4urq5uJBofxkjjGXhIXsh6OoL84HQFBV20zrb4NXSdheDA47b0
1iQ0PUZS+czyqBgtjpohwAApxIREeo3B0jlEUrACGV62lSzW27v6Dzs/oA9d
weaSRoro7n0mhXMd+FsGLNY4QvVcCzF+SGEb1Hts+hIyGt8OIEcaa4sgsZ5s
GLmIOIKlF5TbTR8z+jxnc5v86ZORKw7FB/woBT2QdS27o93WvnuuXZFuogtE
UyZEVA37TnPWg1j8ETXHGEFAJOc1yDXOnmC4es2W6gvw0x6cvaiGvvUnw7CM
keDKsUBpna/cYkYeBfRS6WiRAnsjwox7jLId5DeODrp93/aFsfcGODnNNhnx
BRq+SgWKKJUbZi5ihISO3NRrv7EYcMYpwR1HxDbpNV/vZddGrhpoXwz4HQmX
rcsS7s3xs5bjltuM4dylzGy3XHfEGEOB90EityYfqK8y3u+Jd6SUNYxGxEBt
8i4TSMPpKlL+ixeufIN7n+gNzc4CabEmURgmiWqkNN5iwGiXflMhBry2lDFt
G8zNdG/NLK4gpvuWWbfrYe5h1bVb48IYADGOzhR+q96aDK+zcyXUTC50aj5n
qM55TX8v2cFy6ZNd/1fyY7fI+nx4zouLrn1d+kSv7MxPkPqF5V84PExAJnd9
ekykjP/eg2qrkABsy0feqA8Q1jiazd2eYPIxJ+SJTytdLVjEly8NJ1a8qL5s
IdQG7A2+TSl/nEHk8VCB+zAtbuwbxkQaz6Yoxk0xvnQChXosrqIVrDYI0wBW
wjCy0zIbl4xDiIPuFgSwN0TEzg2UGW2g6hPDX1GgOI0K0tv9eSC44F4eWMli
aUvE87H7aNnw+DZW3snndAYN+YwlklnUW3UvjnBGMlTIfvrLFcuN2moOTOR5
1DW/73xDogaLsVrLF9W2i08znXr+O00ZSGmgEjbk2Xn9Ib1XLuQhxzyGStCS
Q/NCwZlgdU1KMswJg//jX61JfhYLPUZgh9GCaYh7yWATqoshAv+szF9m7LqC
0w4wco/0wLVSEK1Z24UCllBzA2nC/ugbR6SCxONsn8CtUSYfRCSomW7s4udr
mx0xevr+Lo0RdGUOiq+TsMaVXDD5zzerQKl6ESyktx6b5mQZXwQFdhgIgJID
TEVLfw1DAX+hrA6mcKA++tlNLLog292svSBPJ79RRSqV5HIYq6J1vdN6Ktq5
fsZIV9JAKcNFovWn89/q4aTSjHwvVtDUebSQMmYcGChdm07SbyjojqwKNpGy
Fo+0bIq26nUWiZqWrO3ElMwOy0XM8X/3A7H7B7zzq4bD8CeAQTu0RuGTktkP
mTizbDkeahdtWFH88Rcut5A1AUnT0UubHs77+x8x4OmbI86Z/2f1jsToqK1/
9K61dvflGoJy0SfrKvsd7eeHGV2pacYmd/wCQT1PX2rU9tfkiNfQk4dzFi+y
GvnKtbax/P8b7K+Hr3Y3NFAAkdyjTjijsmim34nT4M1Cp0AbtQQw+5Khy+aG
/RujuOc1TSuvALH3AdXye3OEm99HUPc+aBDMFcny5r/2GA3+UTuaycf64iTD
0okvpi9jXWKW3TZoxpZecZr4MbQYNO3o1L7XOSx6jlPZqmtvkonxW2WXgvcP
jMzY4UQ5ST0jF4VICBfaZ6mMy+qc6qN4NySEOrdS6pdtrPAv/l60v97ZOZuR
gv4o/+3Xr3nC/3xFMLTPjFIOpsqMzUXTCQSg3UTDttvRgMLhdRdFKp7hICz6
tBOQ3EbP1jF1k2mblMINmsuX3QcCmvZa3mP4GPJU7aFACWE4fa4A05iuO1hl
BN0d+jv8nJiO3cgNWj2o6jiW+eT47GSAjEqz0ZMOd/oOOcXVkpHTFlt0EAcI
oRruZi35TaCCakyXZkbNkl9kqqPpsaxRvCBAK99XnbFiBhvs/yUTd0UzORkl
yCuv0GxAnyD4Ytu6012XtbBC8L+7tZjD9pqYN5GntY/okT99+NJn7MG5TfQM
/AV1tsNQW7b/cYfG11ib8PE9BnOywfe9+N2GL6rGGAOKkFogVUjuaQRN7sGL
jlydZuxyBgENtjLaRAw8aPd+l82xA3Wk/u9aiQbYea7OgX1pZpobwDySc2eY
NqzzQikCu0PEI0lXbboBFZTiEuzXN9+xmzPeEV5kd6BRqze1ANc+vcazboqK
7llwPZ+fAbFAfPAMcIcS3Kz4tjvkuo8S2ApgdXR4MI+TV4/u3fsyhCQGyi6K
rmB9n7zcCGYl7ZoowMbZqu2TDSxsbd9mx090KZhjGj3PXO88zho3yJ9NLq34
zfQMEDsHWLlxIjWaOSDrAC156PFgIiFqM/PHKZ20M0FrJFxjOQwrj8g/PIG+
H1gZqhWknNUmI9hO86dJ0AZDEkwnB7BKBB9C2V0ZMD14ZAqPZykU4eYu923o
fVhdjKIG1s/0VH3JvrnJq05J3zKhmYYdQ9yFkUjsKEaBVHFdAQBZEWoBghFa
ln4gjURCdnWBeH7M8anK6usz1kbQU3ox64qkuUjbebtWX4pAOgvD6MLps7hj
TvY66SKIzYZ4v1Y/vLbvB+Mk2SkHydQh+7OWb9aV1OdBAynljF4r+9f2oZaM
cSbExNB0EMrAMIRjb6MhWQeoeQfnWbuySsdm+AFKg/f+CvwSKYr8W2c55y89
GGcOKTNK5QbU3qG+kw5zliEwR5c1K6sO6x7n6Ta3/RYNSBnq0TCckhazC2QI
YLqrl7iNgbhoToU3zarfPrPv3G/QmIGhq29cSujPifmEIo/TbOeCzYgCWsvQ
0mNK0mT/Purv7Z0jfr3vZMNSUIzIGFSCJp58s/Y6L7CrFXFuUtkr7b/hG9pv
PGf8jNd79udvKWwSSTC4l5m23H7Csxhv/uQcVv7V6W7U3j3O65vXW7jipLiI
TLemI/WriqvAtNBR7XYU1rYrlQVVFiPLnsu+6fjMlLGwySRkbfoTUjhZZG+h
XIedEUAaaHUNUxWC1HwSVIenpWfrZjDkLc0aSCR8Lp9D0Cf8Vg9FmpcaKv0l
n5I99fKLhH6/cvqYzsf7W2cZnT0WJloKbrG8E5k6LvHnGYPl/ZXoSyIYDyNI
vRGGVjMLgvwsgTk6CnIkVbwUJJrTwhaG7e1Y4lbW2AHydHBVW80YFfn8N9ql
9YZ4nGjGOt6k9zto4XbjJAkFiisy3tGgwizo/ZfKRfACWTr9zXTh9XPSq3LI
0CPUe7MNpNlRWtfeNW40tEmDLAtSb2SR6bItfGdIGJEvi0Gw9ncc/96z1vmI
HGg6FFV1n7TzXTC3JMyxXbtpC72jUmZUFrA3LjCdZQsAfq99hrl9bPRxM7fq
6SjXKj9ZijiR/xE3C7vtiyf04fsBjjGuafnnVSU7GqSSTCrZzft7LAFPyK2b
u1nArrkJiiB6LLJ+rWXBLhHWSgq1sPEdAbdspMjtY8MVPgcpiz53GLMNofEu
dtrFM1FcRkQjHXhfjrbHbH1G+lqEEtGPFbbOIAVKfAc9T2eXTuVvYXiY3qMV
LgoBYjDjV33Qax9auEa3ORNbIji+5040LE5t0nl7RBCqGcMjSJqyFtwxRQwq
bcH2vr2g/0FDmdm8z6mXpHBdbccibct5PbDweC/850lqcASkbDXsJu3HQXSQ
OwMXRVT7yHbvrmnCFjBG6uGgX5SRBZh4/QM5b/NR8X6wSwT7vIS7WfWOMPrJ
oiZ/Ot8P4kyaoVPsfcGmpkirmjCNBlYa5VxXzGCPxrYYgGCfqfdpWiHyAIQj
FYODARh265RFVmAnQayp22xnZwC05u7YO3W2GvTEzJgqgDGRX+Y6JtDh/GQu
QEOP37lI2+Lf5Vvm61Uz87m5n2a3zAkhC5WhaeTLtRL1z/AdznQsxqyrjkgq
GvdbjkCg9m4kMH7YrCCdm0Z3kTmab2Tz+U9UAIm2ufme0ao2sOMvy04y2yEa
KQ40NAAbmLZVq/7brcAEDwAFs/2rQyRQyhN2Vq2p3vFhDuROBlJ5QyeinZnI
KV8QA6iZmZvUFCwsVKgMiwplsZzs+HhpeZLmMpD8askXQYw1/AbK7BXkmTYJ
nLLqO23n8+PQuk6LYWYb/CfvsEiM2O/WVuxmnBwl8wDwPLW3VCQPg2W/2tfU
18ebaSQ+D0h7Y3zxKs4h+MloO2kx4x52cZJpsxVYgGjy0KVZrZqA4V71qX84
LP3012/+3zqx28GLjnH6Bg/sMkEpTb3sWhZ8Wm6Jh4IzcR71hvYGB3081if0
kOWPJz5qcnKaZLbzMotowNnqdIUNSULSTRK2qHhlsXotbEtwUmZUDdI0m3m5
U/YYDSxl/ywQjhrTvIbZGwYcqp5XK1yXKh/o4Q0c6Yxy9DsMI1U6Zu9A3u/e
EVvgLPS0DEm9cu3bZBazF2J82d34aphlXBx5g6iGyHS5QbjhJYyjQKzbRNn1
3s8+bpqecmXYAwADT2Uc1XwwIsoJPuWTX6tQXljl906yf2sI0xI8OQL3LG59
3BR4OEXzUQmRNIa4HrALkAh9qPV+zJNbxarT2Zk2bz4C4hL3GlKV9AVz53sC
eIvVECmGxrt8Z+gyO2xQRLVG0apduYzDC9UZ3sV7xJP14LlbipItPpSM8Ade
3+MbfiCu49Ogc8sunbN8YUL/4Ia4v56yeECf3pVoudM8yLqrP/Y5Kidt1ucT
V8GBXvfia04RYd5YzTGbWoc/u8KuyMSZu/vOFOjM/WND6fSa47gBba/BkNHf
u0cYApjZXwAKJph12sTazVSLynoBR0q8PfdBulidKMeAULO+QDnfbYAa/IKG
BF/jlU3zESFXTmvGTZm14MkiZp/gE+/z1lpIpAeBd8FG/9BpTKI9AQBhOR/0
wXtAHxmag/p9aLJ54e4ZGtH6LPwOuuNrV/7JmtdD9nBXaKbkC9mVVlnvslB8
SSxH+wbHTPlVZBowhTO1qcG6woSPV9Ip945/xmdlr9Wk2XV77udFz1g9A1kD
mRTc7h5fvzBqLB404d+GaP9KH+cPgO6sUNOgWwwqurFECEzLEII5fOTQwiHD
PIxa7Qn82WTgBysaOdt8dytMH0AS/2T6fVVOJygCfP8iy/x75+HBLyaGNHRZ
fT01RJ/TkKQcsuL5wP9WtTS98RLdf7Ct5QuPwBhJN1WFfaYiLGfplzPWb/2a
+UjJ4ee0SQoPDCVh+ew/Omh+Wc3Ki+lzvtWw2ko5WQPkkGTp20WFlERyIrZK
bB1+NTD+by7n/ILuB0iW9ZWJ1sBzARgOrA3dc8Dh4apbLhJ2xo8+H8E/rb5F
ooLF4g056MGv+F1WxtESroqS5c45ADGkI7PAxDjN+9iqcSXYMzqhxmLpL9Eh
QxccAkM3B5BjJU5uQMlewjKYKURu7axOhgatvIA2WWQuMcHYgjx0t5VVjU64
2d/b2m6EMDJ1EmxTyl9aY7cTHagDMlc0WvC7V7XBiqIlBGHKeufR8FwxlK/e
Oed2c739VCATuhota7smXYAPrq6C58bEkdhqe0MhdSamdK8nj9sybmr5tDE8
aXHydZREpdzFYNqz9wpPmdT+QfEu/1CxbO78KEikZoggS4Z+tiZdmhWrhPTm
iCttTmk6JoGnU81+KgnJvFR9ohkS+eOB6wHantIc6cDmSTQI7P9mrMI66GB9
TCu7zZkZjAZKxtxfXMOINSP7GQG07a2xOktFQLm9VJt9JQ5U9aaZzF0z/24b
HYudd/n/9sxwQprGdsf4/0Qp/oOzI87VwPkHIowP0GyNXb/0CbKjy2S+jrjW
5brjtt6m7mrqzR2dWnZSMDpG1c2CslE0r99upSvEdUYdDEjaSixinj8pGr9m
vb7YU8t6xrSshI1oqWQIwRyxjVPUvLiGzWUabixPJMTrgxN3YQT64LQnKDjp
5mh+yP5CeOuUAZpaRGPqFvAnXNnzvjlMdK0mCWHvfxcxNFoCZBjagc/VpDXT
gBBuA2essDzAfnSy8jnnuLZU8L3acMqTebsR+ERvg7H9FR/qLTgt37wSTaQl
W+TeFZ0gQFdsdsTb3JUAzO5VTHyiys9K33bxtsaON9/1y6WYFTOE+d8d8NH/
lQFgAFCXsr9Vr6hVZgN7ikm86lp0Zzc3hK+6Q/GdLykE9AF7qDVvSQwYBqLm
7C29ymmmT7hXGJFxbyTAoVwPEGEQ20AHh7T8uXZUjGBwKuY/oUxNeEQQL9jf
0khKreZCIbb9iHDFvKSfV7P6VNmfQ20JyUlbr0YvI8L34oov+SlfDCzA6luS
TTY/m5HuAXuOc4kqS7mIIRfnI0fqIm1DHF4UsZdLI4bbaADNuAVXtgT36ol9
2yoIHfS4KlfVnwZi68ZjS41j7rQ3qFfzROKb9DUQU+YbMXeUARJZSh6sAGPZ
8SBVL1rmizOWyiFrH14YpQNmdbAgQisnBjhLqaO5IftC5yuq1n3bM+XJlt0N
esotspamhSmBHL8gCMIfC4xauubzUyLova3WlM+99/8NFofYB6vVwIIOn3h9
IJZdqIiafC9/5qUZHSK8/C9QZKS/T7FaJE4riLIQhiDVVNZDY2ga/xHahsKt
fGNCB5q+Nv1MvUnzLc9vnNeCOsoHpGeopaDmbbVGy4GQl+I9uSED234HVlaW
l0PyuWt5cghs1ZY0UdV5Jc3p/avhhfP6MtSEt2VI8VdYI1O6D6t+fq1xFkPq
R2uiyZRXlNfjfCHHjPvhlhHvZz7Z2v+ERG6clS2AxT5/RsBviv7btSE0SnZT
s4htdHA4H7mHGFJmhTinZz/KYiTfmPaQNWumQIpxunOUCsS9d7PnKYDd0szR
MbS01CBmwnfGOInQ+Kz5Fy7rOqLD+kbIC5zjc/w2PQLHiCFp4KsNRR2OiVhS
8DJc7RPBUDgtrOPbsW3ECmPtR8eVZA/CAFhyqUgIylw64K4kcqEcRmJXpDKv
m+awdIZ6uRd479U06ZCNKx6T9gDUSJoaZYOgDOUq84FKbaEFrEE1fndaEycm
+afCwdKiSm6iAhA3oD+H8uu3QrD/ELP2Sgr9ePxV4tiaSej6wRiuEwVmaJ88
XXn58l6MhOaPjARItxMAV6olz1huBIY0lTsCUTe9fp3eqBW0j1UX0WnU8EAK
uRxtgN2zCObWeWSslgzdvc3qYz6At1qJmTYDWGohGspENIaWMsHbgUQiLgOb
5ZgDqFkaQsWYt2EVUfG24YrNrpvxk7Sa7cYuG9Lwhz0OQI10N9TJw9s7HMbr
UsUSW1KimkMK47JiU+PzM1/Y9DpkV4mA5gFOR3xL4BPVevvqfSassiAxOYfs
dZrR/rF6LWpk0qwKNaccdwZHkpPYlpmtDYdfMi/qtBvfYQGt6lUxhveSUOID
LvjEFsjbs77uRutaUQrjwdsnsfzxOU5SinyaMizPYfPh4UA2J+mFPfZIXYFU
IKxVkv6N3CorMbQGo4W5cwphVIXt1clwGrr73Ek/ci6UVU2HX5TpZnRuhYkX
XOUNluZcpgrX8f8pSdYPUM/9tn0w1BO6fz70trzbvY6sAp1GNzU6oXkDYSuG
Hj4K1+FiSqoFnsCkTdSdhUIkyF2RlGH1aMq2Zw9kfdjBGSdkwplwVHD9eKDx
FbPh0Pi1gsRKLqSaG9todnamqXx4Fy9n86+0arflPcx2z2CT9JCzS2u6rchY
GJUFG5XOgGaHYS/xLDnflBFRLvw025XxpAp+53Gye4SVbUTWFNduV3lAsFoD
iSh8HrxNbUURQjoiBtJxQaVQ9py9A9JwZ6mm8bvbhET5ohLmhIg5+2QYlg+5
REnXQJRWAp3OrqDzpwY2kirGmXRkolursX+Eiur+nRUuZMuvRctRjzFRQB2b
cPNyLmajoQEofYzCBC9fMoV//9uFvD8LmiBLfrg28EFs8M9tI+tphvHGG16A
yndV8f71J1n10IFvoPjrJvbJzE4YMj4oOpItrS/UMFREDN5L2h8VR9MXSZ2M
brKCRiPqYClDZqztZz+jww9v2fZcQyTi1/YHOwDzW9UY4yZsXqXaEc1RLFFu
d8nOudOGZuFs2uRq2HWtSn2MXEJEK42PjOwVc6W6Wg36iGA9D7mhmO1x8Re2
nocEfFtWsAeFsFk8/ZbddzpuYVWsID98nvCHyfNmwzve5Y8zyzXJbZbg5YeF
MIF7GTurMsGXY0w7VgmX/LTgTkvpOmQK7cEdX+ciBvOFsf8PeWNykeMIYEjr
3Jxt/PgRiO4DT8BvbUr5jbS6PnZ8dPKTobRLlMI/sUmQndspP+zeXzqmdGC6
VpCxlTzizYiLNpxNrGGwlTcQXblVY8OsJOFXWtBtuxBYbEz6vcWJQHgQ7VxY
xVwEl1U0KMqDQagXaHuNUtDDcBErFmGf4y0/HkZtfSCL4BpFXMPj8eVht1V4
SYgFTYAh0nb2CFbin1jBsgYwBO9uP+sDePqurJlGHMjhVPkpshKfkRBBnRzk
fFiLYRdYgNkV8pCZ3W0uHe6HR2FdIiiwONNJpaXwR6jdg5+A30r4xLHYx+r7
/PGP4MTtGIWv5lr/h0JUQGqnH2FkPlO6jx3Vt6xP/mPu55+R4zDoWhicvBOy
8dqJAT9HU06QwJMzBUZiR4I6PkNGAex2PIb69uQkGjubrH/CPJnQ6ko2Xydj
k01cjr74z1CuESfi8777nyG6UVZLDTb0nr14+qDmch0E2iC2eOLxUi8zqS0t
xd/ObA9hsRcTNtD8sabUvqR/Ijr4KPuKhFDF+o3I+vmsczuweUqPKuF/9A52
9zYMlfBfKqFtjZR0kW3aIJw16ApQZCAcnnIhtylGjAoRZQ1VFp8yrXA1n/8v
gw8etVppi8STICveXxvb9zEfxf3dw2du/5h8WSPpbxX9LNsSC6rIRDptwKYi
dx1v5ltkyABnQ9pRXEgAmkLIjeAu4n9DllVgEARkOPwlLV/mpLzEC6rwH8gz
eMRYgqKxbhkd++dWz0qlMdeOZSS8pGXlqCC0NG/kwo9o2qEEkBfJKl9CwZuG
WDqQX3T1NEKLfAtf76TdNBYtR3zGGcalttb8XMFAf7zKiBXfG9caUAY2X2ay
yl6VaIkyhGpM1hJgNxllRF6mUYxnY5CODUORMMqHOtTWA4kfjIFE5Ay+Md5q
heD9/K5XMeD5PCSNxEGOjj54JenPrnglw7L9Ljfhqqs2Xq6Loz4e6atQhPc0
FT+5SEzSAfaiqmm6r1nk902dsMgSLd6/JEoDA944fMCfPUyTVNbJ80JKxonf
3o3+roOCONebl5K0tJjGcwgZFECV86gF1jr+I+a5RBcIV+wRHKXPJ9h+VhoD
PkH9GdclODKskT7UElzVDWsHdBcnH0V6VEpHy02RoCL7nFWuRONp4gCCWua1
V7jBBTg9zq6BVh4NMs/FkLI6nQwCC2YsR53ShFsG9qDrSTYaNdAMYBkGYLCF
FNW2I1Knh4g471Ld0nulmDgQjs2mZRjwfiMIPNdSVb1tF676o2ad0fMlRuhf
f6JAxEdChd+wJa06pMz1cgwcko8jpxbFRnQL8FvzxgwGQnfccgSGMhN4IH9x
Fpqb/NA4TBisrqq7+aZy9aUg8ncecax5NAoXXNIa3iLDoiS0+LUvOe76zQer
7BkZnE8D3dNPrDG0//fIIGHKGdR3+l8zVtTqxXOZpxjDwG3V61HRO5RownTk
xzl10eb8zuIqvjTGQgJI5epv4XjCCilTJ/VQ7fk7Nx53d6evcRauLTW4KBmB
tXWDN9+Z1Mh5910ZJDAr7+nLTv8kj5LYCIBoS0JYM3kJ6lo8Kr0juDjtYthH
pHCDC5rqd9iR8yeJ8Imdii10FFOKDnb/A7p16aeLwaLqygdwDryh9Vlz5cc9
QOQLezlNvYKgQYBvqInbq+9QGY0ugTNX+1vAwqBvbvRj0DEOPOK3LPtcaYHc
RPlU226nrfyoP3FkhVckwsUPjHCNerBig/v1+pMM1ji7HnZzqAif3iGICvxN
lnXjPymKQabBtL62dIuAs2k93WBOV2HVIhkJlOurlZbIfF5Soq2AVa/OMEAn
Gk8Xpk1l/dsozXgpVznIhr1l8VY84pqUrKg8AhdeSvhBMO14rcQsurvrMWTy
t0W9J1pZ3Bw1PxhPwWkN47CwJ4j7uCS3FWqwq1AZe5jDRVlpuK3RSHCpIf+9
P/bUXD/QvOMV0p2kYYg1iTu8y/B3HH9o9aU5UE9+B6a92Dde4rVXD1mkWG8X
jljoTwD785CtH7zUQhtZDhgMxFClMmTUDAnFO6ZzlsXcifGrU44r7n+bMU4n
Pm+NqmCMgWpODyeCHMMczd39TbhBimSGdJiRJeIbXvUALHhSXUK82ozd6tDO
xHHTZM7j0xr8nPEgj2gZHtNlXm5ttapKCyL4ByANxvsHL9TbgC/vTCTk2eHa
pTqRwzktJSxVn/c24Lj+vNjeWlCFLYNUcYbpNUqpTGgHv/2J0A3iT6A02v04
J4SEM5WVN+6bujdvQnuMbWduH3yG9MqGOmoCNqHq0MYJIFFaaGJx6cE56mbj
XpmV1w76hB5F04nlwL1fyBd2Vf7xRoFgCRbd5NuNBMe4S0qAawHnf/drWbUh
1HtWE1+ABlDy0wtLxQHXZE2JuR1MMI3RN98dORb7NWFxEjyaY+1fZpsEIJbL
Eti5YDPQWNJxcEUs1Vm4Rov9PZxgu7B48fROEf+PcUFdV4qwV2FImExBk90n
hHb+UoYVPvW9F7ry90I//lZtQiN18HrI149ngmQ9knlulWZcWtX3cvkn5Zf4
EkqDzKIAjHWygpcqbDZjKQ+a0jQD1C7V0NBvWK9sxgpvihSPxHKL2tg8z1YF
t+J0bUDp10/S8DiyJsOnvjZYXyULGBuQLy159uyDGh0LT3twL6QIyqRvjnJq
o3waQb3oAkK9qFTlt9YR8VK59cUulckG9Iu3EYosJ+1gtRWxwhQih6zO+ZVe
qhyXa8diLMA2rZWjcdvITizbj8doXau7uIwDTul+Re6y/4KY0MSflqsF3ioy
HcegUPE3zHZRZHsGppnfMtAhbShnQJ182JQEc7w2gizxCv+bdx33FplsCiR3
o9qXkvWjvgoooBuCmyWHWOTjrkRdSGydGG/WOVsltIuHuHJav376cleZkhuD
g5QCNNGnqvgKTLyRORJSd9qH6+F1Fh2J80GlgWDkFxwtaicRvcBJJQIsdlW6
0cuUff21pgakipyYJyJ+Vxbkvgc8IWPH5RWhFZfWjPOpOJgnRKwvmDzDGdue
rAwhEtxs1f37SLi/wpquV4RVnxpfj6s1hZzEQYOJKbkZUUrd95DUfDhAvREm
2utwWS2dibMi8IWlZqFQd1dWuhuUTJiF/zck5TmN9ewz1i03srWTYGnS1ZUK
0RoqCMqHOZ8qq+PjkXC2ZOAEycXjPZvEfJLoty7rIxMyF8809NMe2zRfFTfD
RUedpZuc6zDgDWhN5OYHOt6xhHycxmdK9J11GL2tpVc76Pu0NbZNZks/s7BY
Lajx3omZCHaULaBhBk+v99bIZRlP/Vq8qju7uINSeXTjGSvifxQUTZ5r0nWZ
/S4/CwyaSBy1D8EJhK8UwePVh5Z6MFXsbHvQJG42E1Q2W4hF67B1EfYF+2Cn
pM13FgeNuEDExPe0fLcetzmepvXZG/ukOv4WjhEnGYEFIZJ6Cr0Hmopr9yE/
k6JdGpO4aGoop+84sYeVdC/HK7L5ac/UlOUjNxunx1ZgOsqfye9Y2nSGIrEq
lY3TY9TdDhJwdJCvUeVOCdize69XOjrk1Gz24P36FnBpshamoAlGFCLPr6ci
4WEqkF8YfWcbCCvBdx7QbPwuKWQWQWuqhrBmrJoAgrtUaSqdMh1avm+drEUg
cR9cOEP4sANW8sw2KACVYubjqNim0o6bjWKOTPMMOhFX+WY8uqifVAH5hhFI
0UrSki2eAZUQ4ZBckXEDD7jZ2nqgS7OHVchYFrTYqdU81C6d9bQ52us7hjwX
zIUb6oYGJ15oxNKp2tr2WOeEyJG8hNbIaCKOwtl0Y/sMPliIAdOu/TdOfHxJ
VdkHeVdUE3MyUdd957AIXodAhF7oQvBqWjmRrjK0pEkOgCqEtknk7AjSjxvX
anlAjKm8BWlRjfrEHNwhJY/tnJ7s8oTmIY5ktXoBy/UxJ0hO3dH/TnHHQyt3
pTco6kd9osYV929ijQZpe99OljunHVIwZolBYXI5cq5vjbqXlRdoLDRJLRZn
1xxfCOzSrJFK70oONWTmMSdJrgOUpgZ10yxTY+neQWDHP1hG1uPv/pp84Fzy
4BTy9YM9DAVNxTGHcMyBhqDmEWNpKVu2C1ysrHRiddXX56MBrpOL9BiNnU1t
kACuf4mh60jOUU1scIJjQXpVl8h5SnUZsbZEbNPQCU09FBeyxygtMB3muGXn
OS0lP27Oj8jlo3fl6u5Xs+YUwoXxbQ39QjKAK+wYlhfJIEY1wzqWqGjZX5B5
gBQE0TKkZqSX/VEIlcf2DcoPiSjF+Z8IqUs7uFYUgTFHeVEpXYb3GMwuLkb/
TOACgEU1gvqC7DhQnrDxNp7GxpayPtB3ZVl3P0hX22oE194CZ6thk9v+9EOM
eDqwAOMyY9dyKkDqT8oAoeP2ioWJUDaYvb0G/rmH3kayVmfg0d+ZKMeJB1JR
/YiSxd2rKuV0720eClA8gxAvDE7ExVwp/o6vcje4ONYvq7QVQY5CGZcyNCh6
nWwfXibKfN6vKFZHntNmNm1i1iCmkviskdAkeCaDhG+dFUIu3q2SXoIrQrS2
eQhJcVBWAfu70kjCfukVTD8g4DugiKevzPe0o1uTAhNtZgwFJW+Lx1eml77K
KD5Srae1L5FObaQvmJEcXRt2VaqSSHmeWXsj1fpVJ1lB0x+jmBDGUeGV+Agb
m3xiTIsryGj0rPZz3RdvFacYoYx8zHf7x6V5sEzK6Zb3rabhZ81w9ksk2dX0
tcd3vZhdCsNMYFQnRZcO2Lc6Wr6/3qU+Xm2L22vW5XY8DAq/8w567fZHEOPV
LE9+S4J8MK5HN7pQVmObOKvkWDpA95WKhTf+g0myQNDeqwIx9SwTEcRTrpYp
0DbsE7uIRzzXj52IrLL0rQ+fBfhSdCuB8C10zwmYsjFw1mT07cqt+lGTPJeD
4PQUtOLwgXQD9yt8YFtp+ZLb4IpSIWsAVFAUFB6StImbRIheFLKaKOlwCX32
8nfxvwDhLYCae3PLYKroRZZKy1a2fAgqqO8CU1c2JobvCYD2Jcm+vnCO88jQ
2HJJLXCZO6xCc5AodpiOtwtRvYELmtFEZnPLHCPQtir1L4Fm9d9J0KgGaFnE
uL0uBTmi5waP3q438D/Sd0T3arKEBi07JosdIO72cpgVgHe8mTqEhGnOW+4V
RXZm3YKScqtYrWNNgsp34i4ngVWlYa3lrY6vlmidS0Dvn2/hmlO4L9ybIaPA
UumCRNfTnraU40CtJ1nxi4NIoxzEIIXL+qhDmPSijQA/1ju65prXyZDPvGdq
lcXY54DaMFVMZy3JiP7UyR80t8uZ1CHmGTqiPYai0HsCrsmv4uTSOHWF8QFL
uym0qNzagKDS23mMokZPcH2RgNGgS4eWwEzLzcrIQY2pmkNVQcPAtiezJZHW
VWkQXytpS5iRZgFCDvIAW+EoEaFnKhEgzUDp3WcUYfwQ8U4ttl6YhAp57RQz
QVAVQze1VBaFAL5O2vnnmt2Rb7tCoN0m8GjLTb/hpXgXcHAg5q9YQidDzyBr
XtzOzq71v1+1AWAqrWgtR8iDtzhAe60uiyXnSfsnJT1oeKAQWPyR6A+oc0mj
FDGewms4vd8i/n4bTkdSy0lmzSfgmsCSe8QwCwOfT2WBn1NIU/Z+zboaH0gf
rOZ5y8nlBQbS2QRTvOxOyR5bUHQ3AB4KBa2ZUFPxkbN6U9qChHeANhmz0dU2
yxLOzP/37ZcFWL9PPeuwTxXXLgT5TqJBJii3ywiVlRdjBpq23Ktqv30eBqf0
13dmkIWoRvitnxOCTkzokA+ZWlTcx5oAOHl9kOpsXbO7tktYVZwi5puKfVxg
+Ivq8QUoHMnFkBM4nfjfdx+d1KdK0VqAPCVMBVjKw8m984cldfyr1DEKsCT2
wmWZf7zggUvRIwGqIfYS/XI5cQDbKm+7iSnc/lI3BiwdIMhl14EsXSzx+BDB
KDnkQbamjKJDsqsulQE9Dboxgm+z5f/vaChbf8KXaklYWf2z1yEzxpfGbtdZ
Iw1TBNcFTqyBX+wIBe0TUf9PjbqFtFiCNDSpvqhwqfnLWTXHV149hJ+VK/tQ
LEDBZuT8uDF4OuAcsz5d6vO7xq8WLcXQpkNpgh9P6NMdlH40S5LmvyVv3Fbo
2/WFudvagWCDFb89wf/1b9HPuq4Hi1/3CLp7k3rXgwjfXXqm1dN57ePgZSh2
crbi/prTdgc6t1LkDAlRvHXtpDYMmvCatA2Arfu+GHpq+dqiyHbCCbu/RRYE
jfGZyX1yguI4+DofoTkPwcEuB6CT7nwATpKHOkxoZafADwp9vqE5Ys5PrbZF
Bez0j9tVLyHeFeqXG1CcSS8PQkYAMZCXrErP67mAkS8wWgA/r9YVMhvzJz3A
sAFcDcV/6OLvxf2k2/1z0HYkOT6OBNJQi+bYB7DobK9/I3w9zl7Sg8pL4Zsp
iizVrWkSbTC3BXZE7svSSNkvaCAXmDvgCTQifHXWhwiFTBJA/T3/13gX8kyc
VUQv3fGHHBCUQbYo+fzDdx3Z/K9IyhA0VN4g+m2S1gzXUGNnR1O4/YGQhnAn
ng9z+BmGv4hGlNIUI/Q3vbwHYHuxa8A28YEJZ8G8TJxrL5s2zOedVR+oHanp
2pXHz4brgwsQ9RIM+Lcac3ItO0NZUfp+9mVh82GjIlv5CHjzxLRvwR6uW497
G+vmPC6sosKPAeSs9m/bsS3+HvsDUirz5WAe6nRY5QPwml4t6/1FjyoqoGut
vmyswcKASeFV9Mnl72LUR89SJku9PQQRqmnJFe8nzAkpg5CtBS0iytxcqzAV
k0twkhxtLmbB1Lk6IAwUjUFij+oqAOPMJmSsK2BPtmsHf6EtZo75f8i4iCdc
TsdqX5DrNzyeT3iWeKrKKTo9yQ6AMJAfCfpCddaj2nAanir3D2EiOEyPimGv
aYepSsM3VTwRwOjbd56U8oErakk+IppWISTNiosfKEg13t2l6aoM9JAih4KZ
QecYy3yW1ZokUMUTo4Z9vbNVWFeU2QZGoOvCy9wQ521rXHAczTrtafSWnv0x
AaABvxIsG2ZZIpx0ZtSMw88W97JXYSHyRIaaOVGTCOm4cixfdKwzjhS7gYr6
IYS3UNCDkMFQYP6j1I4rskaGA08u2lrWiYZd+f2bEML6Z0MWjX24KrUksGTI
wv/lq+tm/MM8D4YbXHREN8q8B5ZcJ+lcNK6tIMTNzGR8LYjPZcN0foPdqv6D
vCnldLH0LBEBscphQXScXq2opPMd2lP9VxHwMH/5ojA0kSNb62ACdm5Hoal9
91ZWKnYpvaZDa9bidKQoR1HLIaylqkGSkP3+S9uAbzJ4LYO3TkCcnoYlbSST
z8bzt76VpzUAokti/ZbYuTOuztaNzwISZBktdo9Q0C22Z5ni4Q9ldTyhbQVs
XNjfay0V2C130ECj4ke31Q4loR+ooBNToxPWHPfHNfrN0NXxUqX5p7W8AXQm
fdan9EHM4+aOSmVH2TBY5ipy8bU7CrxCHhvSB/2mk8N/CB0I5gVTefmn9Y0A
o0fTuOCe5jT2O1QmGHHvNqiAW497V4lETQ10jJp7A8I3XLDzGNHVX79t/4ai
ONUOSCbsgQwP1iFmRiXaeRcYbUkp0voeMRxXnYASgT3B5dHuB8NXoQmjn+mR
Z5R7hxE9yus3+ni9Gd51fBCdddYds4wrq3QbnjSaUu7Y3jYfWWOOeURBfqUF
qStK3BrnltJERhX6yl86neM/vhhRLGO0gjbnO+DkLbeRNHh2RTCK7qN5/A6/
Do5qKJAeHyP0QNtWzNOpJndxyZ+KRIKEZLmNdCMxKnQK9iHsSVRQbyh5u+os
Xqz8G4mlRM9ryGD3sTFS5ZnVzxBO4Z9WWVVWXDDmK15b9MQ6esn/Wcbd2qBi
O0HcBSZlVYQ3zFY2Y5niNgkROyg/2xcJ9kktrrl33OJedND4h0QkdZ9B+LgZ
mtZns6auf1UA8V3qkTmoDQyFFf5bNz9Q8hNkp9PnnPCuA7K3UqTa6EUidhQo
wBnfaqxZKHK/5jg/cgPtCHRjaV59QuxyXd+kWTSzxBQXuha1oYUCHoNPW0YK
i6CB1NvvvvhKU5EmmPqM+jANyoTNt/BFd2GuPGp9SoCQ8yArmSRc7ptb0RzT
Xx/JvW8U7VQFfAhZPsKlLRGjkyU9K+D4nSpEhNipPd0bmWNQGdCZllNGvRtB
WgIW9Hz24lphPVFYyarHfap1cf0rlfkmk0fIJ9u9I0OVGeGPzfiKOWTYfORo
TUZ3OCr4ZJ4RH2BuBFmvtOniGh45fMvlfsYK20hrfaSbyfMhh+uAEPpdHWHb
rz5q/N1QgXRaoIfrX2Ungpmbphltkvn7xuNDBiVzhff7oQET1XC3bkWXH+I6
c/GejOKq6qOJrkI3yiXnX8GRDNJj4ymAgB3qBuTI+dNdO4kIXiUnqXsYhAKF
xN5KCo2iisUQtaB8Ut7Jv5jZxjNc9D6994SCUnuQdTISjO2LvtnxP23Yym2A
Fv/9HowlbxoUB05Zzv739GEOkdek6aQVAl+JxBTrVq1/pK+Ec+kPLCCm5DEX
88JwMujcaUMLKkc9U+URoTLEiD91Yi8pndQb8ljbLhc2004mch4T7OiGGrKi
hJmkAW7kNTPtfyx0sUOGs38GMBrdrctAcFSK2ULOISMCsGjnFCjaw0tqtoeP
9wLGfdA/iaAcfrRl2QGgSQkg8HE0Hf0d4ZbHPmEZt2uRrNYRNcYheeq7S4qY
lmUGzvB7TIiomf7zpNqG6t6db8/ykL0r+JJuWSDVmXWR6rYpFY0vAhRggw+A
4hQNRmtGvl4pwPP1mFN4MBOETDe0mCVu8eWKM/cWAJZo+pDj9dV/epl+emdL
K/Fwkj63YrFp1UfSb0CCrWgtwo/gZWzklnRh1gFFKdQkZjeJS+jHmNfMu8sw
6bTKgkDwJAu4ZID+aJJSOQ20MeQZE4ASVNpEghCxfNm+x7sx/Ct1X0a0SfGC
wIpUqJnl0i2zOfX+GBTqArH+v034Wns84TlSFflGH0efUIWDO+dB9nCI5Ixi
wN6FkUQY0bdVlKkFLUkg5SjZwKnDx7lLNGfi/Ir5jSE1JA3A5sPoeyxvZ8bX
MX55YFvB3njM+cmKoLuq5gLsrTMImTN/w+vYXzoRHB5zlR5kHNRPYk1enL4r
/4+bkV20zmNXDrjDlCeJJKK3d+iH9NVqtzRmSPP7yVYhUa/aoeAKqFRLOn2Z
75/k2RwFyfpv/6H3AKfBrhM4XjNnk+baVKchnbF3Wgv8THxkGWJgt/II9lqv
6GPU2HTmRrdxaHD+rlFMroPA6XgpH495A9zk55nZWwB6JaKULa8Oq7dKQg5r
mEBaY9CSENvP0adB0uY0tePywaN4LUaLMfcOt5khDMiDSLbGQ9/Mj7rC/l96
bZ0oKK15VqXd6I96NAp7vSh/0y41V4OTcfO9c2URoDdSh0S64hFAeJy76sFz
TcT8ik1RTPR0peA4icBA8E3t4LjH+rIXdBtlViUR83n5pMFJCIYrG6rk3g++
s80WH93pFzA55VJKSudV0PuX2ph+IomMt2jB1bLBnnuz8p15m7fsX0erAuep
M5CyWbUB1Fshu69ZsmAMbjMLtc1dCPF0c+3Uaq4u/HXlD2EHR1r135aOlkFM
fVHSMmRtzxzEsy5J0pu0br2QnMwjXcoiUsCw34CSP47rMFl+4M5arrh5tABI
LAoPROELv7rU09RPjuCFxYlMTdbOwXEU6zShaxPonCgW71PdVYHCu2vCRUv2
SJBw+pHotLUQBALxtacKc4c0C9PguE9285mIbZlR6fe5paCmrHLqCWMAP2EZ
0S/yqsjzRtrL02kBWecUTnufL37T3dyk/bHvd+OJqxPgze4xqI6AARGRd0mO
1bBY3Ig+44oz4A5l3PCB1BArQnLxpj3L8gouicPBa8+xhZLgx/mDu75DU2YB
f8oftPkfBvkMsjWvVLAprAlRHW84gXuHU++kejDrbCYanwWQ8TIEJH6Mi8Yq
xM1Bk/+YQFd7FZk2CSjgsLxLDYJSv1NK2W8WIkZUihBDSquBBIFN8DMzusX6
Dup9wsJ2lFkRboNGfQ1tXXu/KEbFKud/m7sC/OjdR8aluByG8SXQxR2Kejuq
CTq5I5yWsAYvDvtvgkiHI3WvzNNsqHe6B5gns3MG+y430LHfgpK3kOFOodjB
dK9SrHa5TQHBgnP3ONH990ZwJ0/QwTV2aWW4f8Y7UCEg3LjvSD12H+VOjFdm
qn3Chmg/hACOU7vlWcfAfhX4Ri469xGYKx6X1sMka60sRYsRLFe8xXuYzA2o
msTEdZJG088DuSJUfchGzZn2b2bB22Hj4fHegQR9cqyc9PD0poE0qcV9gr8L
n8UNsKia8gq7ptprkRNrc+8nqanP0x8LrLkko2sH86BWLIJNGdeTAXOg2Mvp
q2D33rICdNh0AyN5pIbciQyufXNOy69Mbh5OJth6vJuF7MR3JqYGMzTYMkRC
WYwzn3xOD1imeUHamEkhaN4HYu788n9t5PY6fRsNPAo+QpCiHy0U2dMLYFP5
izOFFlIMzcPAaFzDJT8RbbDlMloERCiv2BljTyQ47azhkFswCm8YezJiONZH
lZNV5t0H6u5ii1SD7SJHrbjB8AZLkTeRr/hrVUlP1y80InNGUJqBuFXQyZus
0rV+4qi/5nDX5JUZyhbNfHtGZ+ze8GWFrDif8Xlzg6ZJRPNuTHcXdCUy5NOF
Kd15eUF28pJ04/k73VzONFjfpGlJaJ7UxalAu9tDQyirh6OPl+tS9/zey1t5
SnGTpeQ2MEGmJ3pvdbzvGVJLm1NhsL6SdB+NJ29I42Vi8SsGdPnZw2tPjnCn
tOQHkUjw0GCxa2dDsDuLZ77lfXj8g4+FNe5ph5R3Z4fKjZgwd6VFmgf9oqdh
fiEkJxPzbum3pY5rQjMJZBZFqQR+k3xrtih3cmgVYouw3y8Zoy442frMA1+6
BwxbNUCibL0ebxwsplRCegleCe2tXpV5Rqj2vVSes7QJgPAU7TH4VVfo8yBg
aen8TEwbkrEQ/ovvLkZS1LosTCQ4VRIzn5YLOASSLkbl+cauRC6Ed/RPUgTQ
CoHlLEDgFSTrTCcl/jxuK9N97kGyQELf5lI1GUyKq8NXCqHpgaEj3VF5zEzf
GCs5n8c2dWo7gqpePM3fatNOnJVS5G5bpVRR+7M2z0MMyo196BKoWuRwTdmr
Rvc580bNis/WbzShQYXHKJt9JAqOaUo196md/Cks+vi0I5QuBU0rjI7HA/sA
ULtG/T4znKJjM/X3iOMkqHwAzoyM+28+Le4Zc+XFHRgv57DI+OQUrosy+JkS
ROkQ2YCIu1c+id6gw0idDaIa4P3GivaJrq0LMD4IM+XK21ELlGxWXo/I0bLH
kc/yrCEuYEUWT/Iwg7e/v1r7yOfHUM78Ki/BBkogVbsawxy6fal6lFqs+wys
CLBhEDStI8dWA53KNrDpW0WGuwW5C63ZI6AxJzdIA5kiCxnv4wp6/6mi0egO
DRqOOfO2J6P1xIZY10yIfGEqA5itNx03qVKepO5KriKWuK7UDW00CwFhFbl4
EqILkTMePyPePTrkZZ/atDMaesAz7LZysubA/VIk7c1LG0eSjNN46XPDNQh5
o5VjMqXluUQKkqTTlbxeh+njU/QTmxbzMB3+yMbUTWm3e0CrQrUSHtV2fM4h
wEteqXJyokKT1TBbuOfv0FA0y17Ushy2hK6U/cIxHNX83MKQxmxLo4TvIFxJ
89auiUvfmaQPda2Lba50JxHkv8SLsKRUdupwtOzYYdGHfz5o6MfBMwwzUWeP
2D81T1tbu+BaApAPWEyIKQf1RkDiefJDFGFIP3RAmDKYandh+liNx5hvkR6V
ez3t2WYT77s/YDwR5Qe7XyqbL1EFwBlN0iVSmYDtZIrmOtQ4kvPVzVHojVcZ
A4KPV0cb/eRH47jOsJpNPQo+Ze2Xj7P1+CSCs4+6QqbJfAsPLlEcdgV0rSw7
RQq5CfVTu2KsWXHHRpbadV9XZR0r/as7syVFgetRs0+1ivxHyFJaBIzW1eIN
C838WhQCaGem40nJoZT7oSmbJEp/LGdKsnoryTxN6jMWvkoLQJuTmGo4jDmD
e2EkdytQJdON1p7rL2VXPVjgcj1kBJiegu627rxQA2/+z3e4UjsTZCfZgf7A
7Vb8BsMWE7UlTZ14nYiq1Jj3zgB7FeZE3kSDdHZtttJcSkFQkvzq/3jjo4g2
QI3+EiEBr47mciuAm82BKdPbZHGS6qs2G+6VoEGKo4tFeh0EbIRq5vtOrR7G
SS0r40hOuC+/9fLWDl/h/BO3hA7rHrGhaS0lTiGegsBbTyXVER3zfqH+FihE
XV4N6kABB/77wsmHIURz8krF0YPbNcrLsQGA1bPqztqEwm9UOWwXaV7jnACI
x7c0J5t7EeqKKpoi1PEPy319k1XrpE4RGEL99HgYqa3rVS+g7qooozeicFfo
iBLx7cW1artRkINC9ElSA/74UUuQkL/wNLjGWU9Vp9vegU0o9pS0Yu2XBVZo
QPvrk0IXkHB4jipXIJsMivw5bLCHlL6LPnukZqnctWNc4fw+SGFYJmxM1KyE
dKdWZQJwTC0TC8B/qwrBVTfLXbboZPaY5EdCGDwfuzugknJ2Z0MEBztTGNZe
MycpjR0i2W+LKTkWqXVobWJu1XNjXTreJWG8ko2bAgFIc9I5wLGZsataZVhK
PLh1wErTgjSKzEZP1w6gXGF3Y/a73l6IqsT/ykIH/7xtBd8E3fQOL4ekX7zf
iqI1WOycQoSEKvrxGiBi42R3lDw8L5lsI8XEVtMpZ76beVfVvkh40RK9/rhF
mKqWruRNkKKgfKlmfEx28DuQICHE1R2yn1np+5RrljO2iWVeZLLdV3TWl0fz
kLDjEX8pHra9WQ8KQhD5uOtJ1HpAQoeBybQ/vqstaJNMoN0sUnrjIsvFnVBs
W9VtIqOZFy1az1qCXNZ/J1UF84BmaAJvS4UYQls5mRJCc0oWZMdFwZ2Jq38o
DPwQFtZD/sphOvRKcXYXMJcloOWmurUocDggMenZDhzFpLhuzlXfISTM388V
l58ZsRxphbnpH5ZCPXgIRGrOpGz4kbcZBJ7SBuGmZyG+b8Zf/6UVN2Z3gRCp
i9vvKz2u0+l8nKW4QAZQ5QplUwJGga0CjMtclyf5/D7pkrhUl3NBPSRIRD13
ElWfHbLWj8iDrM70vvaNqYyAGgTr4hRjyFKEBziw3pn08PdmwLX2xhlhz4R8
JODX7gWad4vriFwNhWRZKoP54aQIDtI0AbErStUHIQ4jxxCqI6jmGEcq4WAC
VRfznSOpkGPWYjPa0rNSCyuAwGQULIUFwbq/3bjmofkzz/bUMkZnYZSKLlMw
Vppf8kt2PBcOALmpbuIJWjN/PO5koerajvI0v88lmovmfQntRQGEDnJCYraU
qa3Mb80yEZB31A5yg8OHGOTROW1UEwKQ8nlLSeJAebxhuE4VS6ITnlwyfgPP
37u/AmgdqGnkfc+p7X4ds+oErjVe0Z7saKK/USXdEptrTk7NJRQyVCOTp97b
bzfWR5V1ITQum3URDh4OVuxoh7VfZAB40pAgCiZsrbjkKwgrz/lF9DMxD/oT
UtVgU3fOTjwzaS261A5az55zbdPKlCR6LU6QDHIbc6yyBTG7RIRrJfovQ3V7
yfXwhkXani5oIM35Z9ZsvSohIpJBE+CCSBsdhTnIA9G3Fne2/9iLZl/Fn0Az
Iej0y0uqzmriJEmguVK+XIIL79DuGnC+mrQqrrGBbatTiAw2npp2tNGEqtSF
rYl+1qq62tO0fASiy6B9icxzrj73l/0oWF5/KvpoR+pHToBIu/JNT/ZAA2HQ
BU+T+KDjORmvA7ogB0Udz/6O/203TqUrmBE4LITG84OP6z1QW64rH7fEA6cL
aqvKAnbj0GR/COq1pqpAJGx49g+xtILTt7xWtP8vH0uRq5Qwq+i1nsPwFqOU
2SdUl3fygE3gEk0t3X3kQClwLb8FAyCNYT7B9uDSYvCFGLXF/lUAkSoZoeiF
6JDMrzkNgzrfMUTG7ExedLJGMMM0AUjlF+ClU8VL0s6YoS6DuKL2G2XibgVN
K7eiFd6w74XBVAuApewdFzZzBs2w2CXKBcVV35EdV/L3oBvgZxKzo+d7znk8
KyA8bLk+3lwlg9URsOyPvZehk6HReEWYEytV/mSj2oBY1et+iyi/Tn4b/lij
Th5TrQu6XZ+epqe/mn8/cKiLVakmzB5z1K1X2tkzZB7v/ce2a8T+Uizl7mud
Y0Quhgs+D5jvOA0pdpq6WCkjg2F7Bya5ubPm8APcz0PnojmT8TxRWPuMh92A
YWRKt7nKVrtyhFrgj43Su1VkKemVdV8Dv+bjXtDb3VGj5TZmqH/p+gSsie+r
monHaD8PIyBjAongR0CRveP8DLsaasx27CwbPzLujpB0h+APnhCwr8NXsuOM
DpHQ+2hycZl5pGU6iH6RscsqLT4vpJjJJl7RQWEIBcRy5pdv+E6AbDECCUfo
4ftau+jTtGw2i0XDtdxTl40fSBElShzZDqHTzW3Q1nMxxuk6/nq2C6P8L0N8
K5MUHdUoQ3OVT12Ji0+6oWZvf1+M7u0kT/Vt3rJdXgFBGA9o6LxP/QJRf6cT
rHQ8mrzE1/mYmikm9S8ks/z9TPbiZFDyVQ0n7ws2uBcae9NCaohSbS6uK7+I
aUPbtKdaxyicmlgWf1X44mrr9NPTNFGFxDjP0DXPw9M4fLKHSsG5ICCdN4Yl
vL87BpR9ZoBuElcqUO2laI3AeGeJAMmlb4nM5fbZK47uKjt56DD90XZWmouu
Ce1Ue/v5Z7nbdDHfMhJxowW23wdzLmiJq8dFdfbUu5rrWi2JLdr2CyeBx8p2
aBH2/9HK7dSL4rCXfovvqZClEptroBWoMZHfvnbpP8ef8n56WL1bOTz5SiD+
nNU8eekAxiI3WrGWgwiomOyQI+R1tA3B3tycyKDy8/l082SWs9axi0lKBK71
kv9e24VX7gqym8i0IyhUOdduqq4Drn9xTv7nFeviHZQSjyHN8LRUNyjkvSNd
8FPUkiNZH2yJvdL+6AvmKKC1vmUepOBF87aS4A0lrK5M+FX/GElr57/dYUKB
jhY7q7L9gbnFk/LpLeMuunrC4YbSufu/Cm3zk0u/Pc9OuV+TplqiyG/JKQNC
2RA/VdLOLN2wtixQLTUcfsY8uegJ5GnNs/T3HRW7D+FJ3l+nltZXfbIhLBXQ
fSaTBr2+Add75QXHsg+Q+xI+9puY2X91p594W8mCTUtjlh23kfMlooZVjxgG
eMow9l4ywn1ALElSqb4ggV9DeGh+j/tWp0v8Igeez71ryz4X7O0vKSCSyNJz
vXdBeRUy9z0Q4xWgu4nOTN9sV5jtM3PvtIWcuqp+LhCtAWCFbhVEUEUOvlQ5
MXw8cDHK9SkVkux5IjngbUdA47VgOyMlwnUMn53OgSUY/B8v6a9DBefB6ILs
lv/9TxrwBBep1W8HHhDpPJ9ugPU/OY2dEyBZllnvOIb4u1VPU4rua6ZFvVO7
BcdQcQUnCeyd7eTycob8fYHNU9OfW3H/etr/hfoEjySWYnwxEzVHC+4UFVi8
0r9tp7RzG/gPdPjKwIHA2dXCboc+oTnIjB2ujmlMbu33xZ4MfazVr1nptSNs
q2C/ajEZYPi76Q3ov8LDOyqyEG3ZyRN0wVGKIP0djLH8yEyFhZ+7vfWWEgdP
uQlGwqdSXJ3E2ZkxCCIpsigSLL9OUTHYrlH2NToFYrVKJczB6XENSWymKsn6
Ig+eXxjcz6LSyViu/SrNVk7T8Cu7jWVW7YrZm1kZDKPzn5sVi9gzLM9IoOk7
7eYubdNuYY9jBmSGpZi4ulVUleOPzU+7pejIY2MXYTDVeijU7XIojRq/8S83
qG4o0FK5oJhvbMDKE3P74A59pM+rj+zPUlVTHvPcfcRPq0x95Yl3Y09duXNv
ibkIUC8zoVRZN5hKapm4fZ7coaQvtemmIYKV8+9h1dnqSqwQGWO/kcB6lAdT
iGPN2+hl0Q2RdJblbH3GP+Aj3L3+PLhwWLgmXK3j5P3yNFO2HdLR8c7r+Xht
x5at3tlw6aPNvJY0p5XC8dcrvF8ZfachcCo4Dq80GTQaohFEQd+pCEO22iiT
edKuLir6WDiXhB1P1luUay4QKpEi+/BbgLpwMPAC/o45c6gtMksAIFo3UyEp
LuvI8fJ9qHnYIV5RCMRELKJQlOHKO/DZa3HfMD20uW8SeJix+C9EevEcANHG
mpwSHmPerY3QzlQ1yU2bD3rERVT3o8ZdjZmXFMVqgr7Gav/Vkcu7hlPBsuwv
jN7onh0m0JS/jctSdrRRNuUBVZrv23k9tYvSH4dYLr3XgFRU3swtjXH+S3jH
UWQbGLxX4wqe6tVFgIbz6rMfYEPc64wFU8gpsSQfBWw8U/45cswuwoVxl63H
oPJexy8umaPrO9k9MbeN/qGl7RSwFTOikuBNQYelwXhy14CXnyWIzMUqKiA/
ntI7gAkurRWY6Jzqsc071QmNv6IYZA2hyCq0b01Q+XJoJvqmH9PH+p57bTuO
M8SUwvNsh5geWwknOFUjARr2dDADJPiRtFYq5lJmPvc39uGLlKX6kSzlaKq+
uXegMn1CouiJGKR4bLS7KSfsT5urHg2qiBypNEQqqg4xyZPCUuQYcn5UbMI4
1FxrWUVZKgtvMU/TE4X7mLMmKUzorf9j3icJDGqXSC5IMZ5pL1ndeZxxQvmo
NdvH14h5XzJ+4zoWQvRA+hDpgowGCuHTjx1+FX39XE3wR6XPWcUaZwq32j6n
MTgv444Yv0EmPQxBwVDaXI8dvtSF1BO8nMBjO2/16Gu28eqrHjtIFa+5pgm/
Ns4imgwtlpZjAuwoNH8k55klOSTFzP5FunnnQ3NiZ4vLD/97IFrUQgrL4uAc
ObgEFGYueBnse74L9TVEUMl6YmlAezoP9t14IscVaQ+XfPftAakcN0oHUby3
OKkH/DjyJGGglHvAjHkZw/OWm49lY8zchEFu90f1BGpcTmBjCgZ2cl2Pd9wI
QjRF5GTcDNg29BtZ9jUIvLGwDI0yrqtsBrewLY9sztOKdvclenXOH+xSelRp
pvb31roIReZMD6RjMwINsyiKq8B80w4ovXVMaBA1CSR/VJAd4+aVPzb8IQGk
+7GneIzIF0p77xYh41lhr1OdeLJOCnhMo+n8YgbBvrnYmY5VxG4bF16F0e88
BdHpXWhfl/sfX8F378h3Wz8QRxkKDj/bUikSZE5GPijehW5yVb0AC4EBkVQc
3k9JC3tvxz4xAoyL28EsArt9GdPmGJ5wxbCU/fP+RIKBtyCA5b/SCmJP5ico
7aLb07HUOXy3d3j3FiQBFqO9kbrSCfUtGcWh8cDmSGUO2vxCtpACKBWRyzFM
hcWDusbgUT/2c6hhjrNbwt/JcavNNnI3u3fwlt+1Kl5bIQTwRlNYM91dxGIF
6+pCBX30j/N8AQN/30CyHSjdQgf/MKFv32Lgqkeb3bYNlztLK/kNTyYDST2L
crkrtxoEkXQiYuNvyTdZ1PVUPqghtOJy/N3a4uB6AGHVqiNLg/d4U+zJbXUm
c2cBFv2YktAD8w06oKnAY1JBJqa772FQDc1LeLadag5DWf6b6HCRKvOcJ11M
qN5bokSuJj0Tm89dMGgXMuEubf46w9jfG5f73DWSpDfja3JYxDhMNHYMddyN
zyLtPJL3hOY577PzlWnPdLgBtRkBBHgBMY3wKF8QxOS5lf5k3V+yRzYh3lEx
XPRA1YFNLLLwBp2hF2youuueBvlgXfMTq0MteqtmM16zNhncdzoHvr/laX9Q
1OrjtQoLIPSlv/sIDGlkbwU75V/+ZnRR+uCWAU7HzO9UbrgtGNCqEwCTnBYP
mWRFpp4rofnYG0BRwQPAe7dMB/mZKoMl1JJinmLUKk9Wdb6UF4s494MLnzln
8sMywNQhERBdZhipMKbSTWVXPc2JI8/dMPXLhiFSKSpsHiBK7qCCoxG+CX5j
nbm9wKOtF6vqSnDXjIgF+RiMp5PI6bSdZVBrGco4f/gXxZ/5u1Mz+W694bee
w6wKiuU6TgVim98OC00ktIKNYS2Fdu9pO6JLqWDBCXgCh+Jd36uTVDmS4P1H
2L2Mm1JLoXUFtokAoqxS5bwa3jSezU1AhRNFeuPFOyrYySvMI3ZQ92Bcu1A+
Gk0pWh9vzDfrFtQnqDOo5snJhFFzNyDYxLX9H0YLc5nRo51MLe1mfL5YIMWh
6nsL871duCFphhA1YTdOwMlzhNX/CkPGy+Nqg0hwnpqnLN2DGqQK/Wm1ft1w
Vk/yY0am6b4OPlQJM4KLzMArIxru54jqxLm4XHqm8AO48rMsoUTBAYctybKO
CA04lLDKBJgoiIq+pts4RJp233Up+sz+nh8oRf4f+BT1CbVmcE1GYnPUAEPV
3FTxe0nPlz9hJID2FvKnt99W9UEHa4915wgeubbDkr2N26ArOzUwGN3ecbQE
I9X33/7jKOckKPfhSkfanKls1nMtEIRIVVXpLqox7j3hkB+KeTQv9ESR8eut
yJLmuQvan7pnM+kKktXX8OXaGLiEJMCaWrdbJdsJBrqZ4B9ww6JTxTTnJzNf
wfobqPVf5NIeIVvrgamIlFsaIIIO9dcemiWrmU1XUnW82SDOAig9ivbyNs9A
B1RRnG/n1zVMDxCNe9xadymg0I5tfrhebCgRpJlA918C0mclWkqD2c3YqNWV
4QRaimhEYGLo8XlflcWcGzy7WSi8WPoThlQZ+6dz7CbstJEBcmDOR+NPN7u1
qb9V1w/1jbpXu7yYUHW5WZmr+nPMwxXn4r6IyKOLXKzTi3Eaj33XEu/SWV8w
eKQSWtxx15a//AnBVBj5R6BVPgXTevEiiluG7ScOqhIYNpzVJoEILZLqO3jc
gl4H+SQ9+52pzWMPaUFpJBT7zC3Mpr7KYogRWEpcL+6AaQ/YVT0mSODmGECB
FmhY1it1iqnWbwD1i5MgcVRal7FJJpxOouwr40zMU/VXTf08+uVOePza8jtC
oU77x2e29USwpAFZ9mbL2iH0ensHc9Wr0I5knIAYTc/IKok4YayrQ6GOcoOx
osPm/qcLcYIUu521I1KNmRFIQFVNPExmY7Nos4TZbAmNEmDiRMnDHd/pt5tv
7mLO6WWv+R8pFhEM5zKQFsA2gZuVWvmNpBhSgjsLEw82O60dbb2mFDvbJv1r
wQKaLv3jgG3qelt2duVT4v10LIWBQXGnZhSmL4T4z57btbcjNz1XY3KiXVTn
VzaW3zHiinfnFaeuoHKBH45rWOD7Pg54Q6iqNMWgQlNIQI/mKCaCYJVJgtme
cc538e5rP0cSsgGp18Nxxe2m75Ux57ikRoQHD05vXuePo75Aj7CTN3XavvWW
BsZl1+ncy+TQN/ndM8x4GJCtG/DiwcDn4brwo7gjtFa8BQZjE0KLl4JcJPxA
l3noUEy6u17qftvDs167OQ3xqQf9OWRHo2LNMUg/mP9xAJ5ZEY6E4x/Qb18V
Gh+++Z+NHzl3c2oj5aAzhp4G6gWk0Yz94M0K/6b64ZRKxzjnAfA6np5M9DQC
ajS6dQdfbvhSCfB1FKlexk0eFX7nY7b3seldxOegEUaB7pFK/quiZUuoR6/v
g1t1w4gT0SAOL5wHk4ovTTmsCRlY0SOIwYTJ6wBl+tvmXyfxNMrCG+L/svZZ
DAe5wTDZ+I8Z7la9WzQVkJnBvjklyYQROap5xfVjbXyA/UlWCC75/8P6f+2N
iZ2DlYtxfoT9ifO9HGqIF3jVYMIAZl//x4nYdxk4WC4DXLy/S2xPrqt6tcDM
80LGyYNNk80Q/abWwaR4Lj5uNO8+6Vj+kYgcISDyWfCEFD7zJc/V1aZC5cfb
Fg73We16kvrs01TSmlEwQy7312Kv764SW3oO2PzqjOf86W5qP2WV1B8M9ugi
Nxk9ei27dFzDREXD/O7lw7C516tDCPS/0UnKiXb4P6fZUrVCUmP7+8WnL2zk
hXiIydi2XdCUX7Ko/Wee3pp/FQYu9uTXI1egWSncxyXjlib+pqiibrPIy4I7
/0OOalEIjqDzwPyKMxqawPAH3e90ajljwJ+IJbew6l6MHXFi4JpVXBesIosK
GFgJo6w03605E8G9yc1AqBu2zXknA1C517DP4xym3JELLRihLDtz38pHgUMK
o++sXmvCtk9QUN3qzf6kaul0DlGFcbLBtgQYMLKZ5UlfY+1D5c1o2cr3kIe9
uMEgZg3snt4QOASCfJrRzDhYi/idLKKdr06tklQaGJnlKo8GrKUXR9mA9erj
jsyU5QihGZ5J2AnVPN8Pq03n74+DUKRe6Fdit7JgK6YyQKXz31HBgHPLBLKC
A0j3HKsvviPhjpqGr5fJ1v6Rd9jrpHURCn1EYbCVmKuj7VDtdsQ9fBtcEnzz
VvGTXUxE256oobkDy8G75gXDwHSYAFbMn4WoW7QXkWW4qPRQD59fnDjzzXrX
6zzr+wG9dKe+7u3ryHswIMy/XUuh1BWu7Jfb6ZFmp5wAPq/iIZ5CXgXcQC89
c+KJfmt6OIniUESi6vU2ysTG5QIPG2dxUQaumE7JVHBBBzvq/Mf+Q4hX2+6d
A9gdzJRFp7SUtEqkD3Y1jzfkDHkr6mvIEv4UompmfDKOzeblE7NPbhaz06AT
dLojYrO8dnSd/lRyIHcn6i1qOYTxgYSrTy1iiGMd8VS2HevIpGWo1NLbizXp
Khb75ChHSScQ4aHcjMs7UHkbw1cUqW73tY2unIJYFuzfgr7nZQ+SGKVbIEah
UD5CjkKkB5XW222kYeYqhf193oDVOlTJkIyLVwaGMUx3dt7E3OO/H4MCFiGb
ACscMqZczdbMvq4ChJWqSA1AS54SCuxAhELVgfac7xo/OI9ev5skzna2AzNz
eRHFQVigzxY0CT2xfwRPK7rg0dug7E1YRBwzKmDEsdGpQC8VaolIrSkApwB6
wSI/J7I82pHnVSAsnByrOd8rqEMwhTLFR8rJhXZrRCmo3OUJ7kiC/Azf0tb9
y78/2l0Mo07vSG6WP8VEX1S9KRA717KWN/AbcuZDJOox458qtIkAq+lmdvXZ
Py/W8D2inVIkI0LXhowAcC4atNRSUmWmIf0AaIaiT+rBT0HXq8yJhikT6Snv
/DQT1l3QCo3aKO9qJjmNX0mAUchCsJ5X6Hq3/gIQ5eQ33UcmKsQbFJfsHLVu
JZMWd5H+ympy0Of624XzDBSJwt7HHYOZb+GWblQZLgyLvV8U0ffix6wfuDXf
s8aX5+7+rgjlnCHeIP6G2vcHSGFFg0u+OHwUKgUEUYnDbFB/4ItqhsB626nU
R6jIB+JuCrDmg8Pp6RM0doXOXpAaC+4RtJpU/dPZN07zQhonNAfAYn3FaJhS
PgnwM2mHbclcGwgIuAm1U3qSQScuU9MeJTRc8YFG8jzK3K2D3he5B+woB6Ve
ilfd41NQBajelt+5jhTXJXa1Mao0BN+pM1CZfGU0rTfkeV8FyADX+akuxLNo
PVyXB5Qk7JTM7FNh9jO4iFy5hHxJ8JbviZJ9gQr+D/nF0B1gI9ffnmUPIn0k
KnNO7ghHdwyUIY3/EBPwmNSF7BliWJw4GtUgcKoM46cdU4B7mWJya+9xjwZW
Q+XNRGF3LK/87VOYD3LAK3bcZIqDsTEgxcFJ4P8x/k9AjABZHsE8ahqtHidi
kYPeO05gIGhZhBVqdaCEGh2H2urE6g222YWP1loCX39yn9cU6NtsCnQdGHOJ
uzIuPsadB887vNFMJKsYSMuf6IRy7wDOl05kffQXlxlfvxxCJDdLCTYP4RQb
7Cd3MLaEe/zA+6+g/NUsQRJ3MF5DhVVgEfQ2fGNE2qEPLL+h2bjfgii0Xibt
pcEs71trJQDL1dQQSfss8781UPJIKR3HcvPlLOpzXdR1LrB5nqKgAAEuX6yB
F4eWpOok1jPoeqZeyJRcXo0rxihhO7MvcgohpIMCW76cyktJvh7GlQ4XwuJV
bgM2Pob0WSuzonwPGfEVXbPGhE4NyGQWxYQKZ+Cea+/BTBYQdIEOrGBc/nC4
Y9Ed4gJD+Y3BOaHwDsM51QLyFlhlMycxJQL2qJeq05Nv3sluI8dY2SaknLLQ
Z00TKvAs5oz25jwjr9kFQGJMUH96nmIjpaP30Hf2CYPD14AAzKgC0uqAGLL2
fQZ1+akYFjXxI1g9u16RpztdxFMjYkcKR1BeF/CaH1xSilwRr3mqgECwYBDx
RVOTqtIb32tqdQen9xIO4uK9y/h0IH3OuaiRKCOimzVPWzHk67kRbW3s2hat
8l7WkbfFISKjf6Iwo72GpyoXNjpTScCK5szwL/lKAb/Diil7M+Xkkhy+z9u1
TGi5MmKI2Elg3XR8WBFCN0mFATUXxXtHu6r64kIgvrCvBw9vwidfIA0NINle
tb8xzZIZTTBOR6R54QLcZ1D0OsJFWpBsdCDA9zm8EK4QaMr8U/ouOGrwbMko
Txknv2KD7nEWsWEkQTuar3EWoqh2NgUgBgXae/kCwmyjG7OpicC7nUDNDnZy
ZjnA+bFI1xhaAbSpsytfuDbfOWHBS/iFH2EadWvPNfNZqPhwesC3o+xJdQy0
FaFyNnEx7Guog/8/fjDGq8vnYV3YDYmgdm0pDo9scfaWDcn7UEqT4cwpZOkB
P8/Cq4Apri2juo4mz88X7wJgSqpDyys7vE4nDVemRxz6Ie2S/BBtdO2VMEw+
q5CbBdrvcan4QDfHsX2XkpIc75IvqRaViwAj5hzDuy2C2srx007HOFRoTcFF
4fCjr7FmLDQGP/zZRZlxK8KEpI3Nq/O6o/dxFbbU4KZRxjmKfhMI+AsEfTlr
1jAI94lJvtcygdON9Kly8bRP73UEADDa07m28AMmhSC70kmDffLXxuF5He2z
5ISOuyDKVVDaNruZAYNXD0HCE9mGNXRDm71HkGcY264NiPhuYX41zSxxMVvA
EDf5fmOdjLRJ4v58NFnPqItkLCzOOYCcSjF2F89ivICkTthqRdUF4383NJd9
AV3N+jKq/5HDXpNxs8aKaCOoOQQucMsNfiigj/C2vr1XXnMpW/KrlWMBUfOG
yPfmuWmwgtqCUJ01EN3ijXCt+oI1LRy2QMYdvnWbT9Yva0RiJTJGL0IHybyu
ag/Bf6w+PxVqhU9RJ43+WSwVtvBTkzaLlz42ydjRnDNN85oOMZowYFIskXOo
4B1d9r0HfzIyaLS1pAgq7ZIuIjzYXqX8uLX8tCzWSX9l8ETMN4JX1o1hdzq4
2KcvP+f4wotbAFGbMh0Qn1ghZr58ypUIBjc6fTciKHYDP1kwiCwT2baPtxvk
k7eSiaKN7wuLJDQVGGgEGBeRwrnR4RPh/MJUqy3luyRer+embhoZr0XOOqWM
RMakruTIP0GiNGKXF1nf+BHe3TDsH4iNA5xMccSC1LlxCRskYoqQw+l7BYTl
fJSHd3yVhDr5DV2Fu6EQHxW6etTx1fgI8Roo8RISc7QIMbdh6v2hSWp1UHmY
Cz0m0Yx7fBAovsB4GEptbuIU92G3mBDNH+Cmt7ak06AJqJPaZmLH5O+w5G46
wZVbOdw3Q4gazu1M9cKbJvZ9yUGMABpzLvZwvVqsJc8BacSWUffmSBh6WcPH
CY8I+PititRWpr+nKiMxUnRf43dFMcrT5Evv9lfnya4LV8HxEoBrINJ/3Lbb
LXRdwI8HafcgJXLL5pmBU+Avt0+mue0rNtcV80X9sW7mlL7y6s8ACERfw5L4
H+SvF5Fpnd1Q173dnCJserNZz0cAVipoRe1M5+LnqNyG8dSzzNJ6qfiDGHHJ
C9zZhRCdSvGDSpod99ICOUS/3w05+XzCzfmT266vLL5827MvMUlAZ/C3J9wv
9QBQJQt6x3WI8KOW3g1E/gbGeiUPQLeZas9w1YIptR6OC2V02XNWj8HQ8F95
/oVU6yYSucrX2byPEztplptqAvC0BjaSauPVjOJkzHeRt9SvngjgYzPRcZ6z
fbtMJb3742TCID9ejB+Wb/X5GNTRf7qeM2u9l9D2v8tfdGkuSV0tFmsO0kg9
StvILvWZCXSq87GhponASJVV1A3y096xKLtjlxR63fqEjU+lYrD50uGqBjaD
Bp3Y+edXtLY4ssMpOkT0im0jm6AfrGurr2wWDQoT0/+eh38R2QRmQy2HtW50
IuEt0bivb1fxPpb2z5fXYnu6/F7TuBuRlv/cx9CvRfzM7XwyyfMv3DuLNN7+
pEIIUYigEKjbmLxypl0aa3LxF6ZEjx1QkV76alZqHGuPdRC31Fm2ttxYcEWD
1xcmlNkUfBXGGSt2sCiTFMFB1a1MykxrAN0eN6Jd411+0/kSaSz9eHRBn1uG
/9fTzT8Pe+RU7V1q4kLeFx0sg5d874hygX/AjsdrJOxOCi/oB10L5fJz6Jt2
B0iPV2ZBgcdRkgGNaM82cRqYNlTBbVrqWI42akSHH9q2JyTnINe0tt/rTEF7
RO9meZg6Yz0qlTwqJGduk//6ZhbB1tojll+RtxWtH7EIdJcPx0EQXBIhocOW
ZR1AKXA1jrMSbmvPSXZHyzO5fe5nGKUktdkCdXo4kdMu7thpjDCuHSM5bn7z
IMQnGPb+jRZ9FVwFNKPDpIjsgFoMrEgpOUk4mOZ2AOBjbhYG9ijdg8mN9JJL
Kn2AYu8/5UWvbEHVjGDxx6gBGnr6eftCy56uTUTbLqLfdvPntLCf/VDJzLJo
edJkSBOZB3cWlX/xYFGfIpkDrDZ3aE1/+DuFmes59IpZlIBepBES7bWu3CWh
aWoXeno0Zzz0Gouavm8DM0nssNm7MLGTbN1gWbk/OT/6HS/eKLAKKmo/W5fB
QFMw2goQnenyR4+8qzg3SjQL+vSsoH5ELKoXHvtTdb+CFuwxwCZAOGUD9HOR
9hJT2aWjHcxiUG5wqGvw4tBW/Kc7mv1T/cJx1WLwAkJxSfgSKM8eQylp62SB
NHTgUZSFxe/I/8X/xXxxl+K/4g6uawR2GaOByZJR0iCGFMqAuz8JHa8ZMcQO
2F5E53NLHO9hVHA38aO0gq8+vraZbUA0zvglsWbNCYRT4CwhFHjh9w/gislY
hL37Wqs/uv0OFzzlzZg+LBKr0m2Wu4y8Aca+YVpeah2dHPnfEdwF98Vj0BIx
Q7fg1xXRUANz5vpryzcs/MevJUEH5GFMT3SJaEJ0r06E9urit6esTEe6Qi1E
aXf5X0Eu64Bidk4syUxNtOyLbbxr/6aQPJrvtM01yZsFTNOdZKaLkp7I0Abd
U+gaKiwvBnkn9W3ZA5F+4Q6GsxgQdM4m9K7BXTic4Kmq65hUXE7yZlacWtzq
SWMRkIHMD5RZ2aMklq87whQcn57UajWu74vdn0dd5gDIh7WnOOUY+1f5cAIZ
1l+9Ot4M51KPGKiIJIM6j4UmoXqQzuRPh1LwXMeIgVmEBLt69c5pBY0CIPnL
CNxyEyhA1630uSFXT3mz9yfCgxvMyPdrPhJua8yJaXPTE3w4EM/tGQZuyr9d
KUleSV1mmMTY8FnGykh90quULMfq+wKc9cmDf5Fa910LzsqG0h7SYW/+yyCA
uuP925H67JZbUcRDK1E49JHAnp4ePfG8DaKAtWBGNT05MUsh2ypxeM84k6Ab
cNeXtQWn731WBB80Oc9STNdeBGHdL78LHiNvQxA6fX73/zlCX01oMNtDxXYv
SvcrH09QPmoGLwcnJQzeouhWEmvmURlIDsvGPY9ggG/FlAFeN1ZtGho/sJPm
LvfsZNs2aSTvYBUoqDXWFxdYgGe7u0dgnzzE6L5gj/DWCsypBytwa/w9K3KF
wgqb6/4bTXn3826BdTf4xqVF93A6jwjlGul++Yjt1VdHDwLDhfJ4lmfEgYGz
8CJ8kjuomOu3GWVl+e8RG2dCO9+mdTF6es8WBMOWqcR90esPU9SFm9WRTSxN
RHiMne+IXTPPjpc0jm/QGkBI93MR7Hjf5sqN+of1+SMyFurukjSRrhJbU0mW
PgfzadlKuaPeZf4RVqAOVGNx6GTObmcOFdkJ9lqjNuF7djpxhF/koJm06hlc
6A19c6QTKMkAwDtWbeQmtVxXgqne9vmT787jOamBTN50WAvtb/pkt1FkTliS
RiNnPaZSnUYlQV4sQrIBafJJQ8o97gwLH1xdw4+yyHG122PH2FWPwQm5C15G
nstOg57Nx/Q7kfiapZQzujCCGhIeTdMr77ouGE0dNvLrlFCn3jGRpLiM9amG
SapWCYB/Gciz6OzhpEIhuT0sEpTlaxMEnRFvjkqbOlHVZdnmtyrwghi4fm3g
tkqR1xv+IYRo8IWbMhdWdDL0DQqzH0YtX6Lh1fFs8MiojJak72uUlenNKcCo
H8Mw0gSZNTIyN9AY4VqHkykr5mkkXkWTSI6yH9j3a+zyjpb4WHiPM/qJsQ7P
r6zy+Y4dcN8pARq2aTzL51XajwWlSaO8VOIrzg0ygLbkaf4rLwDQ8Yj5dlLA
EKO/moUVKX1EWMgEND0x371rd96nhxRyetXFBV6/xd1TOq3iaU1Tjk5gpNQ7
2clwhPhuGfuUsIrY2405pVRPbOA1N72tC7blxfyzOoA098qKe+Fjq9XFhKRm
+t5kowUj5EbOcaZXVv5WBYbO7ka9Cl4Ow9lsuMGfXVGeE4yS7UmQC/OtP9Dy
4VRW7kMGv0RmabR3h9apNvPjqBc4DBjvOm/kAsfb0P1m5IMHUzUB7pLF+UXF
OY6cY8fgc/fKS/ckNjyfJvzAcsTsGaNALCJakkkLnuYGBIhAg8cO1yMm5dB3
jzFs7gehPP/Z8y3F8q6YUAdfk6Gi0L0wsjq2le0gb/ihxf4rHukGdZZlWh83
7hFKQ8kC8Hq0nrVQk4vtKJzeVbN7qG+FFI1KMdTyOPHRDuZfA7h8DKYPaevk
jIVanG0kuBUHPIpxN806vI19u1Wb0EKvA5YnsNBAYRrbVoVqqA7VitG1SouC
CJKIbSG57Xri8ZmlRNUc/2zFtUL+EOpafQx7j5mHIrhMOthbrjs8xP/VGoaL
XSChD1Z8KY/fdxel5Z1++6GTcLz5z60lBJaEwUHm9KF16BiwdfrGtQ5Il7P5
+MAm8QIGQJddCwi2xMBCUdoqhMA73/IOVqEug8FlBHmqT+p57OcLGhklPN3T
l8M41qSxYPHHOG4lOW0Q8GMab5Q15jGoTVD3N3W1yhJ/hyQTYHFtp19OZYNT
UU7G1kiJCbnEKFTtkvRFNRx2xAF1XAnupMGiFMwTvdQPk4R63bU5BXAYVhzk
AmThKFgrO7wD3P9L5V6Dhfbn70rquevFBAmrn65RhatC9pHfB82C2FPNd1WP
P/dcnX4hWNdwNmxHrsK2JwzV0gSF5Tx0QYgF1FRs/rKK3U8Xe4uEu89HvdOZ
sedKmDt5ikg0efmeLy6X6sP0+xICHn+C/HVdb5pqe9E/ryXLKkeFKf7gpq2Y
9cfFfdXn6jl6fBhdb1t4kRjII54aZkLcwGlGybkolAKq5fx73sLvDWBHjNLG
oLuJ42Yx2jkiPFE2QNSOu9gidBxN9cnMhKCDftI7hNx/1LmJDCpQP2hDHxVQ
TzPqhhXY9rKmR+3InWJqZvORqnMr1m+dvQdBwzNLammIyKw5BmR+W53SiYt3
TlqMwEjHA+CyPLLegWSJffnMZi/NC344WS3l2fDlqkmTwFE3hPmdfEdsHFYj
IwMUkfl9RSgIfFQfjB2KXHNCNwFaYdbJb5lu8rrDTruHMEl6fuiT47ToVE6Y
XJsJHEnO+P4yzu3t7AadRpCKtsxG8qOx1Hpt14sStqkqVstkuaC0shBPeEYa
CGRazsxvyiskfVoCjGxRyqRjJqaaWL+PEzKD5TZaZBRCs4T29GjF6ciENhW0
xBQUWo/bBxVOJ9NK7Tl5a0Ona9hIpUs4g5BFMOWWszOGEM99U4kYD1BqK3NN
3KmQbwBImZ980vecB4Bn27/2bYO4SMbMidSc/j32vrris4PqM1YZfZdlBH+E
UqtKeU7KrZDQ7XEZtDYbUVIcyhfwr7lKBbmtkpi2uspmeXNcQm1GRw+Y+1jm
ruhYXifuHGmCa5hfIrHCeT4EmonrBlkZNJD197VyDg7Wymt9roGh+CfdCbZZ
Di+Rrs+TxLsx0E3cVQxKZ8afxPNX3PU3z3NiSEU2C6i5c2E+B9GmxmrHQ7Zs
W+cEHB31YUiYAyIySoIK5J2EdjKKpMefnIzDFisguja/xMj0fgmV+7IHwvOJ
u29uLiVkB5D4Xp0W1xvuKSqFadLo5qepWmp6vcVhM6lBG0xGiG2WVqP6KuRi
+ZuWsMgcs7nY2H7RrqCGtE01+V0hrF46ahMWRRgOyumXwvR2nF1oCgNLuSuk
fcXcxVPAcoBgLkVGSv/L2hpHzknf0YH7RjFshbYG4lACmEEKqHXh2dIFDqE1
DlI4g/qfIAcZWkarYtDiruizgFj559Car/PzeJ0EdrpLvIUX52OOkO+4sm6z
S7fHEWq1GmA5BDJcHOh6FbEDPgPBN+f6QniGikFy+njYJt+7dQOcuoOSRy/w
0tYgXtPSLub3XKlzy3UWNz5UY+BQpb4ZtYb/0yeQ8fFSXwj12gd0toYdAjlm
x0gQwuCfcA3/UoInlrl0kcE1l+dMFP6GMKjIyDsG1XriLAXHmxdkqMrs2wSY
dTDOwpbWSicW7Du1QK6UBd8UfN69+V6Xer/qRnZkkTKspeMKmwL5pF9TEo4b
LPChq9c7WMhZC2/ZrjKKMG7TkW/HKdkcR4sPDtIhe8vfoCLHobtaAemZZmy5
EEV4ix7FvTlliXtVoy16h6Fb3vAI30kGUqj8F4IipO/OzSJo2tdBUi6xhXQM
WNSG0nmMpfRdA1N1kiP34aWmang37NyGxtaWJOHez8k5SkpF5tDPtNbD8k+B
rG+WK9uLCRIqyFC3uX6w4b1BlMkLR6haOllFudeVgIkm/BEI5ZaI1QB4DsI/
HFw4QZ+3uKBaaFcM6ItjfuuIJ9UJFV1RemI5e/wjClrLxmOvrbkxfAIMZbsP
g3Fvqovm2gJYlYu7L44T+E2Byt8evRsy2PxTTdZPeuXySlt9vGkZeyN3l9F4
aVkD/3Y4hd/1wE0jUHMAzTWJdsvC3LXBvGwIBW17vZEC/NXSgSd1sSKAULtm
ANa/VNQQlUDz6fUDyxFtZsuXi3vBnwuMaBRg9hA2q1/3/c1Dlj2AekiD9jSC
GPaMxwwpr8MA54lhh8e1MRGb3kQ9YAW6Zt7RLLPNRqSTwo3hvuQvKu63BcRk
3YUKeXhrMYIzSCv5ms5+jX0PgmjQjQxRSlsOqHZYKZPmhBRHvfGTlnG2jOj2
Ht82ZoTlwi+JZmY5k4YuLQwAE+PzhcZnKrVURY18IK+Zm6JragoaW0Jh8sz9
AqnT36DKjFlEE717K/o+2ZMn9wgoVGalW0o/lfCgl/clZP3Ii5r3e8N2YJkM
qkHyTf8xXfXWKRgvtxZ9ddL/Zrl8a40naHWQoYIcX5mM00zO+NDGZynutbhA
NJgl+TECIvlVPq2L4cb0CEnpwFcWNv7iDXHAjkhGsGJkcJcSSI30PhWj/BFJ
6FCeqBgCldcWYkpNT2E3RNirSgFWQT7HQRpkzpjS2b/29HFakpdlnO3vNrVt
Qr50d3j68I5wCQPRWGPmztG2pVl5VWJEs+J4/0MiUzAcUE9wHycs4TyVG6pL
Xm3m5LF717nrIMhn8XPzzf13cF3RNbhUNtLrOX2gi8v6G4N8MUfEyCnjjZ58
icdBrLW+0JotkNGQk1QZwSkiRq1ItGpQyWv+j+nSW5sxB9Jl4Hw8cWyYaIab
5z6+WMBszls6r1rcF/TLELb1S12z3yW8+hgmSBHCuUxZ+YDbJ4aedHSL80U6
1gMdhKqR5LGXY+Oz1bnlLMBkRB2wWJUjddM5nqOTrIzwu19gOk/GNQqZDTnB
ASSAK+piZhkJgmUj2sWngeVmm8Z1dKBeE3aQw2AKA8kMW7DxBG9+Gr5FxQdH
wME18F0arp+UH827tpJ71IrgSmickp2kqrv7i/UOoQ1w7TBXb6yabxS6ytAc
TXN1jR6IttTeQpT4hBxN6qbAXaiiQV7ENyFHKv97dkd1OnCs479OJpD+FXu4
0Hj9nTxAUn19TGtWCED5CoMT0cqmf/dR0sAT8Vlwo/mJAm+ggeVOrUuJo4XQ
3cEFVfw7LWtyO2J/hVKQLK4mI2KqbEms7OwZWrs0ygB8H/lK6qr9vmxvpDHL
mCsvylvSt6X678u5XMJ6qnG3X4E/BEzIuwdhD3+VNKzCBwI/xDrMxp5M9oya
MoaA40d5FVfNAmrVqYPdQYiSwBHygR0nxWy2XDZ3ZFsmVn8YKKuk/JnUiMf7
ity4uBbwfdOuAtOt1Y8RPzQBzATzEPbMiAsvmK+1AeDHkVj4iIsPP/rs6daV
/yXU8QQ6JrXl8WfFLRZogLjzWaX29uuxcHnUJ+IFyGzcfTaTnwOS0dTeB10W
BKGxHIuMkp4IEJFomVzlPLJ+gcDesL/K9AvoF0w1FUiVcxhBuOPiBiDG7uxg
3S/X74bnDWOvDV+WuH+P/yYSDuOU09BMfC7r/GyLTPlBX8Usq0qGDhQgZfyO
Yo7eFyxcUQElhBjNyhn/XnOTfCvw5w8uVXWjuadWDSlnEjVlnOndzrvq7sT+
FPmU6y67MJJFZqSHJrU1ZRI0NzL+UygqW3JEpoqX2xTtLc3SOdJGpkMufu7Z
u4qBb6s1Xd5otbDE/aCOhK82i8I5P5J7EbvOpBTADFiyi29gInIfPccTvnjq
Z1VLMquEXM4KUboK+JzNSkslwkCMKK8rEDDx5LLo7/3R68f8sKm8iKKhcM6k
JjXTcfe4O6Hyt0iuHBIekHN8CAkoTeHYF594g7jvZeOpOpva9IQL2DaZU8hQ
uiJbq+gCbCVIzZfYnQPrcljtDAWkI1qUvBlR9CAMgEaHZrcr0cd/eOjSSqiM
Ttw2KGFVqeG7OOj1ir/RZneTkaUNzGz+OZyvuS13A7Vlz10C2b4xLFD/9frt
TGx0QnZ0fUWqlZawXYl3wsysX2JFntkjZpFzt2InVJfGsQItZ4ERu+DB3NPt
8lZNWVGnRucsnqpdpUbZztK9WEWM4GcPP6qkQ65GHhqpftpxXl4K5Yy3tDLS
FtIPjwUhFZPIeaWOZvFR+rrIhtkjLNhR8W0Fg4/C4BQluuUnnZbLQae5BDJv
uDuzLWQSDbs4Qafr9MJCszpQWC1W9Ql4ScXPVosMCrEjlQSkKGQkXGHsx58Z
A9SJU12YewaxgMG5zKLbUho2K+slZ39hhSAeehK0oegoMXFGjLTNUawB0E4e
SL9lEcdCB7IS5tlB+RwGc/+23IrkqVRAEc4turKoc12+0cfgfvu289gxN5E4
ndNu9/asjifVFiQYinreYtpi5u5AHCkm2oIagEdLa87d2DrhRw2yaJW8CmAK
BbatVXn2mvyXkP/vBxIEZcpo7kl+55SW+y6jgiDX+87cZ6onNr/iLcRXIw3d
GYcx7Rxh9JPQLnYrN1bSCAiY6kuIKdruJLBWbLeneADatkjiMoxmrscjyYmj
r8rA55AsMEBYYa1iWae/RGcIlHobutKHfIuUnKSqTVIE+4cNNRyxnEBO1bOd
5Z7v0l+d7lMF+KYUhAZJYoG07XTeJtF1GjmZvRihTF5UjuAMAX5rkQWfDXZW
TwkAbOkrzdK/gcB5E+YB/W/H5wdE/Qj5thL9V/qkJKBgWAwkm8UAQQgLLRBp
n70mTQvrU8bVwh8EWaoveOYRRxqJd8C6PdSMrpQoNfIe6BkKewsqn8BUXmUF
DDNe8x4FmjM/0feijqMecx244CSHR2izLXkJU7tyIGPWi4nsA51F0+A7b+0n
t/UP9KjihQh0eL1icJzQIg1uph8ZnlD0Qc8H0Kz2yfHxAcUUBFo9xjCfyZhy
h+MOLityuh/yRy2cUYK34+bBsFDYBkC9Yghxi3+Se4EX/smaVsG9qzPJdmNF
/bdGWDdAFXn/8Vq2gPTznoaSf6LGiGUksOEY67SBm5+Ni/UuJyVs0GkM+v4q
+RZd9GsssJbsZIJKkGb2k9xyUymDjFkHRdYOxhZIjXzAMHcls2t3IPrd2dqj
VxeN2L7JfjBxa0YVeFryTxq6rjeO+58KUpnmKcSkd7c0NH7CcL3+GT4UChgr
xSdqLixIBTI7CIwEM6Sp0qxyOQfcvbZZwUUG28w8Xxjx6g3mCRNyoUgxwLdX
DekjQcP8g7jCrNkhijjuLUe+XPB9jScx1CkWDAk78f7vhkt3WiXAEw69fc5N
f03NvRJy6dJ+WwerT2q6Cw2Nu/7ip7Ea0RQE/yoPXznEKrSAWAAsVlYlUUtH
kkBnsC9ShcJdWzs3qnzrNRQuYGK/CPpyUcW68tFQGX4USSXfQpb3qmJ6AMKl
MYTprapLxmo5ay0u803Hxc344nzH6H8P0aBCtEVTWIbn6cNms3cuaFc1hBSN
dyl3Wzwazg2Gd6CDN2Rijjebe3Jd8rAAtKqmF757YpQNEPA1gYNz25QlbDYk
2TcjAwJMnM2cHjoeZdXKXeDsKCXEtT6wpiGT5bwv+nff5wNeiXCThMl8WRwH
dEUB7CASIxGTxtzH4JoGfzy5nxgM/JHQLoKCl+sH8tMk1D5dtF1OpJPSp6js
TNGyT5GmN46Ivl7veQW/djgOyeIutY/lfjRp1TCHF2oKb26t/Q8TaBToVU5q
3A37bVEpwtXS91Bs69XiH+uqySIG+kLYEoSFxjjgzFg7RqHyiCTCK/sS9xO9
uJithi/l0g8lD2ZBw2s+VGL0+yK6KzJ2gF0LY52Vpf97uFRrS8TO6fbixpLU
hBVeDhdOXgOufvgEBDX5k47x1bAVxgvl1CTnwab2uLmEYxb5J00FO0flByHa
kjzgCMygaCEuZQtBSQDW7y+bjY9CwtPmbFq4VRaHR0cSotwPkuhuBOAeozwG
K718VTOPmR84nS+Y6M1o37vbvlwqFoeW7tYB/Olh14uY8nvPvIiavycMw5Nl
kv6kLpdd+hucjj0ubs9qNct8+Uz0f5XhWNfq7Uig1qryhb4zURnYhME7I88j
OzTBF0Knp0CPw4mwop+U9C3wAUHZ3SLusI0hQbOzCO4vS1uSnH2GdbZrZ+Rz
k7ePyMMRsLy96YbNnqvvkTQWAvJiupEUutsYx9wfAAILQ6M+TKzFvmlzQgyJ
Iu2Xevx8cfKo9v2yUsbOrs7MIq623wmBgN3w2MxeYrD8Jqk0XwTFIAjvLsKZ
4hCa5lXbeEe4cXKmMDYcCk/4NeGnS5FVx42ci/+HxjmldnzHZ6onZAAOlgxy
x3ihtTGPYwBAmUUabqmp31PAuB/I/bCBL663eWquhyMLfQVBXh9kkXrArl+B
+wQm/CdxNDXbRWie9/5bUbl92fk+cnWkbp3MtWEywoxDUQCilsWQNNIo18OF
4CepBDu4YM3G5s1KsCbjSMtaGdnTVyaZVqhMczldmxBHfFORVlrpkSW+3aIC
/f2b7GZVvZDjy6H6iPfrprsDgMQ9xEWVAqcjBL4/ettGo5ECCbZXTTOe5YsE
jXz5jKCWxta9jUZ8u/4R94TWM/0U753+zP/uzeQ15XFQ2XHNr6CYpkw3+x1i
GLdgYpbo6QMBfm7UqS/cxFslItg/5O7L0BI5WnQPbm0f0jqhi7t2LAjZ2xEd
Rs4jBEBOu+CzN/m/Wzc3Simkt4k22K2KYQ9Nd6bXY0B0Np4BUp/Xsf8ZqQiy
XwePx0ctd6gw7vyFqznn3pv8P8ouCiA9aLvroYiXe02RiYXS6WU0j7B3MG42
n9+7fo0OalT3ABqph+Ti6OqbqBDyKXJsSqvgbUDdidAuXs6CelilzAMUy+NA
LLJi6J2DnL9VCnpNCAY+lAUl1Z4zHRxa8TfI5HlfR7zcBnRzFXoz6qrh77Y9
FoBvuFmuf58PLyQHPnZ+mxGGqDq+NXfzCJf6MGQvXjPitxlnaB1OVMUM5o+Z
R2Hpoi2plEq0l2gKxiY9C49lcTR56mk/E1gmhdtRstvkWMuH070nlRRkzUIJ
zARU0sAL8jrhiteLgjBbMuIQFtdmbSvUmxUcMMQafY/GQcVAFk8XUARRDT6a
d6fKRP5s66sXLgSCwLg35PxVUkDkq4UeQ/x4vufmDP8U9WzXX7haew3+M/oQ
JadIIb56vKRzz0HpX772Q8pt2UcxdH3uSlXLQgZ6fiW15BWKeQHkjTQFDhfq
ThxUrP5bpl2QfbJjwAZmSsy0E3nlK3EgYcyJ/7niuNe1lqsNGbJ5xPhvZjGY
/ndxDZ8o1iLzBnp4LaR205AO1JveUmY9V9hYzTm6VqocmNYUyi31KASpJjai
JB7GztTqW0OrFyEGM83I62Xi6tgvdGnCuc3HG3Ob4ZL8wogHWEE42P8TDXG4
LrYS/DECItrk5OhC+om42y+0/9Kc8S04TcNRVocAueBMmhNIQis3OIYXiDvD
jJQ9EtSDCYue0DkpY4BATddt4lnDuU6Chyj0vUXS3YiHD6+dSH4f9g7I/kjU
Jlky6CkRKH2pAGydvFGzh2k4/tH6i7DcbNzU7xBXxzEOWcisAjDiAiCJkevV
xYWpBgRDYSOmgmMTtIBXcd+OMTPGXB10YifGwCIgC54/WTajbDI4C/ApXMzo
41W2y2OJ3oawU36K6k1R62VyU73oy9laHQiqG9BU7VSvGBt44r+DlI6ZqssX
mIlgbWW1LvpDnqSrnT80Jrx8GjNFshzYjeKrj3ZKzKBnOYFqiqM0KFD1n4+s
0ccjIKRmIwrmA4EzlBi9r1hCwcmvy6brTQAW6PJ7hco4NyxhsoWrkqUZAJ1B
LJ8rMWedGOOSUDLBOIMAAlFRHjbS+BZgxMU6W5mabNGnynwchjpgH/TGI72L
JRODkfE0KKse24J7c9MBZJC+BBYHGkYF4vgyuy0ufe3cAamWfrHrf3AJgxHE
9LEGWLUIbhhDzk3kWh4vwHOFabC5dRMsBcsmfQttpitY78iQ/FPdkvSLTK+D
leKASKfem3FQaJ1Vb5KyJl5eVOOxe+q33Nu0fG3RyYFpsdwSuMKogsnaEeTz
g9O1zGKr+8NKqIDj0n9ka0tOd7C728P3rpOgZd8A9yK1Y6gV4+UWWXMdTust
w1ViDVH3TCnJwRCqfZFuUsjivpIhze+RH/QT8GxnuTZCKRt8/nf+bDR/X6QS
3Ch7j0B/80bUmdGiiDvrvniMHBDPV/8AZ2t+SMd8m07tHK3oFZkAVzfa4PL7
DLDbZlP3b6YMbVoVKyOfFhJnwQ51wtfQ2HZdQPufsxZWLcv7XDYAz6+coKvS
bLAVgAcpAYDOKlDzySSjCn7u8k0PYCDfS2w3W+XCdihPomw8RDlHO4IyB8Er
w2ezG8oRlqGjUl8JD5RJTPlse4Yh2RTbni7XFC0BILxlk53brpQfQJioSjkD
CAjKAeosROIL0lTWTidHeAE77kIRfvGTUwl2+Vj09giwEDayVL053gisrEJq
Eun/Dz4TM0ilq5DiJe+UygPzhfB1g/otxwmrbjDHtTkhdQjt4Nwq9ia8G5Vz
E4GckU++YRrMRBPf/QMd0ldwJaFc+0XB8R7ai7Y42urzienAwTBn+JN+fjMk
KZ7J0J7+MxI9CSJJUjc+uppyeaZ32InhqG6Pjsr5vSv0b2XoHwJxcga2KeXp
eBZs0/tOxEmAnYwI6EdZOF6htm0FlM2POHH2EBu5WLMDTZ/M4Ysn9k+3/PmU
TMF3caPT8rk4A0qedTE7k4jhYYZlViVIUy1Vp22wUYlwc/y0ZFdEbJz9e9BA
6lna9SKnixVSj9IyfUT8IqhNC7DYS44rwFeHdhspd7W9nS7dfEa7N4QcJ6Z2
vlLAEFk8d0cpceF8eCpqvfRwbAml885KyHL7qLxre9SpK9EefwRx+RcJcH44
mH+vHv0MXaUSDbDOH4c2Nv72XnI5XfILRGPikwbqpH8VhXLHGVEseT/Qvzx6
8KuN6DyjsdkVxdH+0WBKsMPrb50G1mNIAJfA5K94WMIiwVP6s+A1uL20zSED
QrTkbBbpuvJv2F/h4JIF8s1sqygLy32F41QvRw58EH+Liuwq5qP9KsSM/eCz
/WY2HyE4TTcwNLJg5au7HMfb8VPaHi6uvmJZHZIHIjQViprQlIhL/yanGxmG
DFDTC81k1QnDq9zrlJim1noBHqu2K2ElyF4OrmxzqvBqLuITtABX+RrSPI7U
RAKMIO0tiSbjpBxGpQ41wSpcxKEf28FYUdvIJX6Ow+CIAB8Szn5vvSNXnNrz
2A7yi/tA+V15gwpjGcNM2bNkO+zmk36yLuDPSx4bQKG8ll0KE84viqFD3Zyn
ut1okVXDcrY6tUQz0WrCXByKeUTKSJTY3zTu3RjapX/f5du/XpKU4w3AP1yo
LBotttZGO0rK6D/Atb+idtoIOpyvIDtpyIRl7qR2bWxkOSDHkUuvzwCibW7W
EC9bCbECpd3oNK+akOjVXnxn+MoWJhk6+hXQTIdkl5iio1+WntUG2GkVQDyb
NAmfbDrS19Yu+uErTURk0kXMTaUSqmt4TMC3iixh+yymXZetIjyAIL/lK7+0
t22idX+yonjVcxIgBiMDav7ebMAJpJhxd5Xsd9bHSnHu/5aYusMefMSF25hr
4fAu8cDWBPcAYcPcOOl6+RU2TWc4EM3uVtCqw1YWwyLD6cz2aU3U+LZNRZF0
PtrSarfXUK8qjs51JR/8wbCUfKmlAonljFWuPECdPEHBrn4ddw6ctZqXQfN0
+mP2+2/vMJonKFU7nqXF/MMbXHyGUrkYRAoEgmvJ/ZFJE8nXdVERkBcRBv3S
f3JInw/aiSzjj3HqJLku1dYDmS3l+gMTynFzUgjhdDIfybc5HINAyGn9LCXp
2DgBOJooge8Bc3XRtMiWsQ5imGrdbE8urN+Mlh91ZQiUb3mDm8U657DUWYLz
iAXds5J4SDKrBCoHGHY7TTt6OKdA+oggPvurumnYxOk4wpBP3BfnTNR+d6YV
nBBPwqenyKNyCi1NLVtHvL3xE/qO/rPOWmzfjzYu+ZKDBuTGKgapUEC8HVIN
FTDCmOlDpp8/VgVXNsOhihAsg7l7RRAnzzrmVSThzj8n6R/oIsJzF8c0orOC
aMoas+3jtT//EvLARhZOg0TinxN47DfVGMxhFMi6VG1DbiZdCh+98herzCvf
Atp9avhOySrTIiGg0Tgc7u/UkqUipKRPQQRKwzANlnuwkAszqzSZAtxAyhpf
e0k5b9deckj1mPN6zHRgpdCFmfkIBvYRbpJi74ASO7RZtMyWkbENIVWQiJQT
IUDmJDGZ+X02mSGdCLJ/9C7LzAJRBt8Ke5y2E9t34EZ9qh0OpA5EXArVmcKl
TMMdyFpRRGJN2meWDZaPx2tlcTuFQExQqxfDS0hnmu1TXBsjw6RRr06WVLKR
zo5GyIf7Z0iGRYNUpDjAFtWr3vKjGb79BWorW5NZx+Em3PmFQDUz2WHwdV7Q
QtmdMZb/nGT/XjttBPvtVjdluarcEPL0c2ueNGDIoEoROFaNxsZTwJxrhWCA
WCmrJUNEfHwl5MewB84tAvlGtHbOvwvEVbzq+f1RbVwyjHpvSEYQrQ2PqHDg
Iu3YmOwlA6157/TV8JECDz96Xjx7M1P9nXDL3NNRV5unpcp5qs9Qaxa9w65B
4GUjm/88/arHCRp8GQCEBy/zAreGmv2kgdEU8ZNwwAKtZIzSVmzQAVOpb1ZJ
8A1jpoX+xCVFhXwJDRkLwKhLUSXZB+7hcJlsVMyhFBUgqGBIs8+btfTHP9g4
rMmu1FVwBn2mU80x0lNpczO2SYR1aerHRkeAm15SfHPsTaf3sIBQFFfJT2ea
QVchr2mLhmQ5DaHqP6Fjj/cbe6iXU5C4dIihf+FE/yWXANQv6P5ILGZ23rmZ
M6kiTrD6xEuoKdDrekWcj52ZKzg3cSckyd8powclLFwVBp9Vsed+WTzN5tQV
KkjyzX2NzysLPRKEFksZAA+A5HWHJ7146ZVGBVUvdS61I/kZWPF5gn2XfQBy
Gtu+e6WOAcxOV5WVO1MPaxKV/1rOMnd2mBrWieRLFgbyw7MbJzD9RZN99krH
WqNDi1+yhJ23wGzoFcDgDcvXxYapJ+kTm66DfHmGTbbApQFohynL3K1m/9P+
HwVkCNCywlxpdQD+a+LRYUKywinxDIWpY9ATJm9ukauR/l/6nCWREa1i1Nm1
8AeWjNKUZb0xEX2H8OG3OlEIetiJZATMMv98JIydF/SQRGE2OMJPErnGfVp5
K+k6tpKWY79oYUFhIRuxzkVDNKc7/FfnNYTiN0k3e8w3coMM4MaUTI+854Qt
f4dsYitnQ7OBsN1oG2lwy8dBpGyegJoH8gDhgjme7oOuRFlLFv/QSVRmrhC8
CDlO0Tc+w4gEc25u51WNLxhno86PUzabj708dMGXh+f+zdNX9q/FYwSOZgTY
Oc8j5CRFEevM+VxLB+yobqQmkJDRVLDuodqc+WQOyBmSbZ3adfZpBt88OrHM
cKRWN8rk+dRhUvEXW4KSYqAX8hJzKNSdeFaJjKBw7hjXxEdmxtQIjGOF1fPc
6mVGncKWy70g9UHErfomdZbhKNUlB1oTK2t8xrNDSPKkQ2EFwtFn3RF32PeK
uQ0lAEr2f/aFU0Wo2Gy8OVZXdDWtrXDctErmyEzZFd70cfLPCsSb5+0Lr1F4
+3unVOeRWm5Yb2hG+aMWv1rFjLL2Z5P2ij5AEd1Rg8pzdOL16Wng66wDpHiF
KmC6EA73dpmwvp+5ecttSihk1u5GSjicuwtDSl0msTRKDnvaBz4F2dossK8s
KFihTWS3pC5UielGuT2cNyy8gXEdnZmjQjW9EpjO7Zas47ylbqDS7zLkSa12
Tujl0dff6e6pB8imepDyv3DOAUK6aq82h3IaZeguWyDnnaph5QpCsoF8/dnW
uDyq5nLTGGuLtmVZ87Jc1xpIvoaCjDlTjNc5/Py+IgHCmyPjZK9Gsr2pChAw
c2C1D2ilrUJy3/VZxl+6avceo/LsZn6zkoZ8OcLgK7C1jfQuFJ+znqANI3QB
E2IBGL1AoDEENjGCea2BJoOLVCXnq+XYb6yQC9Z4MLiQZH5rZmpZZ0/EmIsX
Jsi3D+4eorATzrMJR9GJH1E89WiypLjWupNncaxsjqV7FWRI7oHROvJJQG7v
ybfcNrmwhefjXmMEusqSHPK/ZaVBMqgK8eDRBfwKQupy7mwesO5aY0pdYrXX
MHQYxcYlJOeZZr55yVFcDmJNc07Ebys/J4/2p9amEnRmCobmRVVdSiLCSlCl
kjkiOqlru7RdmeND0a9qU2QOEMraC4HCW853gL9eHbtK0Ovy44lFwdM4bVck
E76WS36gxYT7yWHSsqVTxpsI1CpAdV73/4AFw9d64MTyswL3YWTJ/JDQwacc
xabp3r+uk1dWQKq9Ss4Ic0ni+cX9cqhjSeYFM2wPTK9cX2A3kC9/Nw7KTDH3
yfg9Uf/75FXr5unfHuql/XxhgEpDiTeQ4dTmSLk3vX3ErdUVccKBG1k8hygx
M/My8RiJdMeisN85eR5ygq015WWLcG357mG3w6XxZK0pI/p5F/wp4zzxIHqr
kUeoKmBqE1OwIAKtFxclmMDE6yi2GO5HfU7uPkf/WXiAQBcWU+nxp7p9ZVoW
7WUjH4YHtby9GIm4fz4BFwoXjkPWIgO4bFNJ3iYPqb1NCiMfNB1ufF9mklMH
D2bznRLYe996KLxCeVjbUpsl994BUc+67S89Pb/Ce/pD1ytOOaD0aMP6ggmV
cV9mOPcZ5AQTbXWQ2jIZOh1L0PzYkmDzI2HBkrbMWrQTwV+fnnYz5bBaFHF8
iI7KsT2Udum903QqrjSp6SXriTpi5XmXnIEtv8Ceh/tTPrS2xE7kpnmwzmH3
mwiiH20/kJibMGCvrYNQmELMtCgfqvgIi5YcQ/oI17eQrG3TIN4v7f0ni6+L
uiVSAd7mDTEqMgjX/1PAUf72B6kD2N9LQC4G16t2fM96RLO4YlLSHtbb1ZyX
eMgvlejXdgqEY5hCSJnwym/Io5LxAHTjV2poy2rvJA1pCpF/XvNZNmOM0RjO
x+nWGaIbHevEsU1xQnFH38bLFFNWc682/Q20QwdjpR6KILAVGn5SW4oa8UEe
aRnNug66gaup3dJUPNDS6zsC/DQXJaZ/VYHlD0OPccd8NVuFlY5ec4T3zNqH
ndLArGnY/nqzHRV3Bk71aAHpuEZxq2uxhuM4tp5W4rPWN+/OqA0b7jKxW0Lq
+er+Um3joOtMKvELnuUft7jFyU7KYIEEmcQ/3tIkMSbMI3iwCeo4crsKLox/
mnYLdjPHB3kq8weNAfm/3FTpbhpON7p3hm28pS3Z0WvkQ8ea+Bw8dVPtIqqk
hVYFtdH8gSSPOCycytQh4PoDxh5z4c3usyah8KB/UBH1LLPTq0fOG+/DN5pV
0bJJFpxTHrQ8/YlBPWCEr1+RWfFHtgKZuzFmlmDPiKWMfNI7NVKXn5pgtCmA
AohSrC4jOasuzRU1eVEWltEQiiqSXu4K85ek8hDQFi4uhJgPnREv3Z6QEvHn
caPNSQ5TXrcfnk/pug8ggUfUeFZ8iw8g3HEZ9cj+UQ0gYw01fKGr48eQCVJh
Zw2ZM/oc37vXRQi/yO3lHZgtnT9EV+/g8f0mOx7nXqVfx7wDe8kMRKmEQaiF
W6TcWwg7Az8RWtZ7Gwa9MHvrv1vwdCEj2EkM4dpCPcEDFYnQSD60uupsvqO8
m9Wn4w3PxPx7vXc7XlfIHVUZUIENPpHrkUq4CBOClCiN+6UFjc64+Vk1hoPT
0TtxFxyGSqW4sJOB9OSYYqWDY4pE0TLGMwc9C+rXT3zaFsfSWVx/fmXtqs1O
rrqVpiJ6yNFPkGwHfc3vBPg3syWLYH3idJlrgKPdxW+d7Q9O9Jcn/4bdVPS9
edUNhjyY2FK4fjMW++Pm5y1+ftrV++yI+f7nPHmKUV8Wta79XJNvaQCgvKtZ
789VONXgwlZJAKB2Tt1vkzDXC4tErpWT81cM/ems9W7uQj9XMuGzug8RB2DZ
3HP0+FjDOCU9X5/Ydoq9rdOA+FmH5lnazFuPd+Y4uuyo+bmzFlrFWziRuFKa
N0lkEQZuP1zKgOSGb0oC0dmHwSe8N4w7VSQHBE9UDpIpNfPIXd4+YpmCkfto
MpVfcezifqInzk0uUzbPfjbgUIyjmTE5Zm0XY6RRdT4EFqsWdo9Z50gf0glH
o432UqhJ0AadNfnJfH0S4Z2ROuABwsA+d6NXhTs5vPrg4GBSfltacFDcsJok
PpK93/QiZ9kc+m39Xh4sXLReQxztMRoYVFplzopwj1qYMC8Lx9wDVfmN3V48
VdNbU2w4wW71jYZkqNMyo8aExKXBgbMEzB2+eBap9/3q6JMuAiPLEpY1aWuL
XBsGyDCh807HTA3cys4UwS/neJCrNrvsae4qHcQtaI3qdqsBubZIah43U1zk
SL16Lx66+F/Q6gaieKZOtOxwxeIG6smXhAr8KI7hAx3vtdoN90PH/K4WC8/S
XRthRT4KhYU+Rz5fMCJ/GoGNm5f8jCOVLsbu3HmwTNtoFEqtm86PJyNgMsze
6uE3iWx/EHihGZ2MyD9S+Q0W6XiPVvgOgkTllC1CMGg3EQxl45Sb1PEK3ROc
oK5rFVj+AiQuiR/wIs+kpGMV6l1r1elQaWLODCCGq5aaqrfRZg4cSMXCGOXx
juEqZVsLWLCRfBvhAYDIJVCwMmdEGj8pPXAlvUxSSRMwa0NqG+RurLK6uC2r
EwjmRQC5R13cRUxa9ilpOURTijnFn2EwBjOaxpCnJau+4sHGKKXstRetIp34
gD/PmxtpdhkeULkgWmPM9+eeM35AwmgyhtFHYF48z4B0hkKk++hzfAC9pHmw
+L5o9Y9vVM/ezEl1e52mTWg4ePaY1j2kV4I1ObY+zKGlgCfOqnngpE86V/3n
ffaaGCq1401oimKDku4dQs6o8lFAccAB5K0nuC1VSTHdfhlVb6pDsuJkG97F
a8CS2iAW33uZNugPjCU/FQL/KXsyL8Qz8IVHk10g0XohuZ5pwLJqq/Kj8NnG
K0D1R6muhB7C8yMpQIYst+ojXDG9jGSCp9XE3HtYDC5B9O3zjMPMZ25caMyH
5tjl/sYcA48MlVBSNRMZNusHY/eo2z80vWmvtlplxo17m8PzXam2ULJJovEG
OYdZ+UQyxnP3iDiGAh/p5xkI374CbFKC9I9nVFMvAp11w8sr4US7lwtMZIC1
EquFz6yYP3OME3QqWFimvqdOvqwf6pZi8crX5T4Dtw7q4B9arHRhIYi7KJrW
lMqIRx20UzaUgvJse78BxK1ngUK9bmV7pGxkXwCu65D5hstEkp2e0EjbpqQX
tmOSyQmOpvY/QXZtpbcAmRJLGoY/wuAP2rzOuQ0JSGSK7XzinSvmZ9IakeUj
aaEuzzyCzH/xm+iYc2xonFZ0uZbZeKbyKY3pw+d5qVOVe+JNHdJPJLVa8zjP
IB1GzWi6Gw3rSJE0Sti99SdqVqLwr0v5NAWExAteAs9i4nOrFYlplIJ8uPSf
3QOZ0m2Z9CzYhKxPfDltpU7PH0FSio1qNnrUMTpxYeonuvd49puejRzVAOt9
x3BHx+GPkJ+oFL0XmbRxkM/esPOnPAUg4aJPVZNGv7O5653+56Mb5Bu+MIe1
FXWj8TMvsjxQisiS0z2Y5KdrmP3epjupz2Q7um1Izrdsk719I+l77MoLDK5x
qg5i5H2vg7v1QzPBh+g7Pn1MS3uAy+Vq0mDk02B8FLZd5WUWW9lqFamEWl4N
G24weQB4KmavCqzyXCYpFVirevaB4DN2v8J3PAIZqYFqh+YsKcTRRFoo9t8s
3BE7yfeS2Z2s8xRZBoo/O1aLEMbnsfTlZ/Bt63ICEF0wcMBC0CBEopWVA8PE
vmGFlsbh5E37oHKtF7NCb+Ez/hw/TKqmNhMlucID0r8YFLKb2vLcSnFRBpjM
PJdkyRyIlz3EB+s8lAYUOppFyR89HeMFS3UHWuD3fU/zom54ysRNXnAUxjcP
i6vvq2vggHlYgTuZRQ98pmnLEYh725SFhyGZJs8pLgeDDRTPPfCdQ8DQhHMG
N/o0qN9n0auQ9VYcHWKuwvAEVfkaxm/vHEGN5ttKY8uQ0iiMJ7u94Fw0F+pT
/8yNN73potillUM3Gx50+IO6ljVgmgWocteYtSzaLsjsXg3SFVaV7qHa03lT
Cn3V7U4MKPz3X703/r+Eeop1vL2D1+maYZQrUC2MjzN5tTP01iieWcy6aUGT
DQ7ioHs4Mp1ac+LN7frKiu3Aa3g5QKNLCP0FKAnZurrF+MwpbzN9wDY+2v5Q
LYoYYfRZhDASMSCWMH6H7a067lcBqTnM3AHt+3oFUBQayolHBrkWqWdIwQ9j
to1itkfCXfIAundAa4Hiecl1TqirqL+H/MP+SIX1xBLctwaxzjqag/6mcERW
grI4NxlhSjQLxNcNNavBZfeFMxM86NM0LoAoCc2q4sT88hEle68jyVB55yhL
y2k0kPWQuPClO/7i1DOJPhG2psPxa1uIfITbuijh30pdW6erEgJDfD5qfaTw
uNf4VMn3OTlfeHYElc31VwV1MaMV7IgBhC814xkqeAMaO8Bri55+fPIXnjWJ
e1JIbZCZrUpqhJAH9fEvgMBxMIOwq3OPyHwaj1g+1cImAU0k0Ja+d4jM2HQh
plm270MsEEeN/phaOkKtR4kS0NMfg5pcKcULoaYPNCUguJVQlWB9Nsg9SS0z
KMFixnT9kV3oXBeo8+htIkqZQfH1PhrUdbk0bJuydmkrf4m2QvdTYkpnc9ej
7boZe0M0gBtg6M1KcShEMiWv/u84DSxnfiO9Kgwne84gsPRjwoII2WHgJw67
FDfW0aMN/8VkPd9hBFbaBjkEsQ4w3g2OaIvzUwlOUDxgDTdXnWJmNevx5ZMg
yoecEHGE/m8cFg3kHS3oB7QvXJ7YzAqmM9tNi0JJS2ijpE/2OS/E3Rz3+3xD
TBBc6XAdh4C6fXn//DASzjJ+3A5TOB5Iq0GaySN38TwMlcnP7vPBTNNLyX4W
PkmUEaPbJcub4hGN9DmeX7GLA8vsg/t2ntps5KkeeYHFFD5QQdQ5UcztefFR
ZDNmae9jyAmqLcQSO8X9ok7aISwAL6DaS4Tse/GF2bdyEPQU1vf+IUdPqBLB
m2WzFxi8FtWp6VFPc32UtW1V8LBiy6hBpOY4aMgLKDBqu10nmp3tWiQkyMxg
jV9ET+A1E9SZIwrrIeyQxf7BnWAQySnNtb/jtcxWwdpHdTwiD2xRR9Ktj4Mv
k0wRWBsYyPGlvyp472DGjYdobFdhNPWhiQMghzAbib9cMDDgfQ6+Ez/bTz9U
Ml7CWOwmf4IDQr2jBR9fmxDD41TOi59f39yiInECZEer924HRJDf6Y222ND/
nxVoqdNtKBCfQQiJpQJCC4OYXyodZD2GCv2b5zAi/+CY7L5VbA2f4eGocuEv
nkPLcMBE2Zg0zLu8bSRbJf+zsE2gFR8kRHdH9lvR63t1Zng01K5tXpYS0HST
KiM4799+7q3abF2vT+OJUF2Z6XwgOEwFl5tq5vNKJZfwEAsA/kCA8ac2cyy9
5qF8nlrXDhCbm+N3iBFEJPdxayozOmZiJoSyT123QrH4woEhfE3TKyZQEmfN
bcqnaJ+yVRLJZ6N+3GWr3V1fUYfCgJcyPBC8dHEwrOMLu1T1WZDDkXL/BIg7
NJKUPv+X5Zmy1FmhS+QkR/QW4xNjp6co0TM/N0Gash8xrH1gkUgAHr7KiUYa
L8CtuVm07whJlMszvK6GrNnDtbJjSjDHQHcjrupkpfEBT657sqB7PayktRwN
TFr5kYrv7PrZqVHKR6WMNeBqa2FJae3a0vrmkc9s2DLILQ+WSyELzoDrH0lZ
NszjkqRGvYgIeYG+6128nrD3ntEkACJA9iRbV8/Ejk+NKIdKc5Eqc/+5kl+W
DP3jcYriG70aEJM+VEyBHBOtGbxruVTUK0oEoilfBT/lE0t6mMyovjxFo7JK
zOLJ2p9lRQQ1QMMT6nybMDa7ep+pxabFE8msO5uZ9qzAEZ6pxFgAJRATOUkC
nNpuhYL+qt3nsi7Wxmi594iMRFm+ZB9W47CLNZ0yWZp5WarJxYEpxV/lmsgu
Y9ejLz6m+q/iXXm3pTCEBASJ+uZjO47BXs6FfN2071/V7oE0XabF/1fJU4m8
PpIlrbaHDnFDy4T36Lhvz2V8eX/HjvJJxX8jJs2BVe0xwcXN6240EDB0mj9C
uMGUUjJgyXfclkPnmHFJan5upo4MdUhFm4yyg9sWPYHqOhA/7AsOFYzkU5Ha
OxeZB7LYf+uUKfaPnLkCU94nFZDRwSIAGfe6MvpBQrRYVJinST7ky4UPgeSx
IFyqzcARDo8dXetE/m0bqd8ZaqFEDzAcG3YKdEJXuDuUfyRqTAEmV0c0tUNm
Y+o8Ri6zTf2iItSOUDPdecnPHRsT29sluT6NMqg3dX51HTUAj02gLJ4I759z
sAXwrWl7lRcXCOOVuUyDG5m7JUfcwcFqRKF6Urfwm98s/1dsi1Zbc1pYsl6d
S/Uskxcfcbv/LsTIPHxmwTsnUn5blcEcJ2uFP/U8IK90DC8RgCHNAFZISU82
Vbey1mQOynVOP+UTHtrRp9CBnq5DZXDwat/muOv3VDVW+v8eO9coVEUlH/g2
HgbJbvXXBBfMP2EELj4n3/yn8Zg1peO1hC2y6Otl8tXJmPlWVOqUxiFcjZ//
hJmmqgVwu1LDPYzvdX4JFD2grOKlxArVG69wfgm9W01bmy+7WZf/3zomXuYH
IcVocK78kDXump39EAjYjK5Gj9rKJNxkvC0oM/BFJpOWXMaN1nVmPMwtOIgA
WFS4Pwxv1Wbf+RV8uHIX/A8wjwnnMETd5/i7ctZY4+JzoRyjR8gr+NhjSG0e
ipZLqgaPgPVx8vhYfJ5WvtygZ5tX/I2dtXgFx3mpTgQcFQG0m3YkF38XzIXc
LBGb+3ONfdj8/SQTIc0rZQl2hJkqii+dZPRUD/RQbJ+1xOMDw31CvFLf4j3J
fo/aI9bSYH6FFO72NK8A2pa6kCS6eBWvw2gFgCKMhnvP/pc46kCBbN2+rsH9
iZDav6QxXyLNgH5+poitV5wZs0sIYb1rFzs8o1QMPpq+GkDvpM7LoJUD4OV8
dzEzPKoj+eiA7+gUvLYBXtULX4v7MDqWeRLCCvvJYDvxvhauQiu+fcFRskpo
75FMz+GFTV0RTW6//HaMTHL3LXBY7aTVdRiAnuOGoXtcGOJq07aKWLzqdJnC
Fiyydyrrs/j5NeomFDcS4etCKE46Boyh0o4tJM+k8wx/NVSSuhFgZ3AXS84T
ZMvhnTDklzxeGKWV/RmUJpAFr6eeuOC0cW6xJiKQPTJF0n6yJYAiFGNsW1T7
oUvDE/vLJBuiauNnG7v1HiiEnywg9i3a6hCjFf+fuCzmE9nYYPm4+n8L1Ooj
vWDKYb53oRGpBzn7NJNhGlOO9Iqo3GAcXsQfUoq+70xWVrmPCo8+tSPSXyWM
6NVJzPUi0YdP7U8d7pLVQQzbl8EDJFDjuCMOHfNQd1xX6jvVGthAEn5QM1qu
Zh6U1kbaC41eGrU9m+316oM9cRWS5L5pxHapN6x/OK5JgcYhvjpdyJCy9at3
z3yHq+32Wgjnw09VrT1a3qcIjxSghpv3DWnuCbd5KXHp9nuEiJ3d+x38MSQ6
uBvu43inBvlcRRx+yi9/2cZJb82EEtF5Xg4Iu/o1Df5CoTBNb4cAfOsu/VJN
BPk8BjKUj2/TD4WvWD2kJqgxMozyLNH+Pwx9+VDu47vdP7drIOJerpwQurKj
nRAzPcnNPO+xId1tkuLJt7gTvGYGodSWJveUG91oFq/Vg+JELfar0Z7xKlyw
wg64Q1jjK65X+4/7NPQ9FDBXAjlgfvcAlRFTX/+Bo15SnQ5yvHmzudXDif/6
9ByvakGLPlD9y67CIDvv+TZydI8Q8Ez+CvigPA+lo/ZeaCdmIh1JE5+jYhdl
PW34kMe0mgb1l94It4AqKoduG8N5Q/j51iS+yq6kPKabo6fTFv5LNyepTD+O
mdCEijmRFtR1ywCwfBWzIXRdQsAKJsngTPc+OnHqQrTsTeAMdSAHfcuG/9Ov
SpF5/452Tvr3kqOvEg5lpGIS+VkpsUTMTSP2r3K4Jt67GcdPH6mExCK0Lwz6
EBKzkdx10tbcWS70lm4PVMOOFIxUM6BKzosqqWigb7RXxSTvamkDbNbc6R7T
QYitgUpmtZvGb21pAnc8r8kQMPqFLYTMmJbputVIF4P29KiS585MyuEwLmnD
5kxxW8ryLg2td0zMv+DUuTf1m1L80Qm7PYmzhqaPWhulBdt+06/a9/x5YaFF
jcUpQhZ7duMc7D06MFaU0Ascx6+nok6FQorBuArr81vgaReLCvVIvsvuv3/q
f6y96PrGTwTSBVsTlGw4kwAYXdEzZwhG+9l2dDpvsgQ5lB/SG/G7NqjsStly
Shnngm1eCfZIFfiUOc+QSMm2gvZhExUJxBebve+zI+NFiEpGAc4iLEFlLcfV
b2j1XuXTd1B2JlUQda5mFGM+idTrbrh2HYUXNJNPyxIvaw1Ct60VxpKJccVl
uiTyiXI9aSphLbhe3hNV40pyiDcJxPl6WDCGl45c7V0lBFics8B2imae9qDY
xEhRwyqPEXHZo5XJfZm9kW5jEwZPD+0JgH3fSsKxKsJra966MgN2bgJdZ9wf
nw65/mYHvE5Lh64z3W+W0NYoF0PvaUN5ihBDHb0YSY7LD2V2LOVG8DR5yZdW
3eDvht19KuHyU78ZY6uOYf0d7JZSqTW5NZmX2YmfvRJUO0K6pNa1TKDcAmpF
iCI7upAG3EO0j93aGrw/T+Ne23FasF01Qi+pxqp3RFlohsT8YeSqDHeFFV+M
N46LRqRj2ZPKaXg4dAoGngD1FoQXhS0IR0+1X1ARoCeWoyxoFDjYt6YaEg6/
aVzxxQqPVZFT2TStU5N0RjMr+Csnv9B7+mJD02+pFA279gOhni1bSW9t/nTS
6fLwTJcPiZG6i96LcSzAmiDi+CBWocMlwGJt+UC59HLqHCIRmCFI+WMk8u5E
wvRqedQxoOh2BN9dhK+NEQl6IQ5Q2g38+WjVDDaVIfkHwgeOYvmUB+znPtbx
Bp6C7HyQl8ybVheIb7K7JEnQHkrWE9lzu37Q6IWczIV+HyCBJNGi2/ZiVvbO
mlmxa9Q4DNwZSKiYaiaAokrxxzgdjbTh9nhuXBKQ8jvkPsya86p191KFl7FX
9ojN8v5cclJakOZR7uO2jBSn5EbAzAmj0MP5puz7kUPIpj1gBXvokGQDqj4M
uPBvTNim08EBKL27Q/Qn5C//M+Gn44/O05NBlAfRoj4ZoOtPca7qFQgJXT30
JYwPzgsBTDDWcEaO0Uy+ciLvsbpvwIx+5djViEkTNTeEXheIhANKSHfwmfRJ
aPswpm01O0zYDtkWU+xf2JpCACIoXgGb2N7iq6JyZj/dq8O2ogNTR5X5Fo3H
NMdLoMKeaO2M85jthIYD1hxGZtkou+p96wIUcem9YCshBpdrPAjhet6D+vnV
qA1Uy9GvnbxcNulIj5UrQt3UDuMD8SOVLoU2+LMaqZOnQbxHWwdSRuyHPki+
rJVIGAfRq7nvX22jcRhPWPKgTs1pYZLOvOagLFUCei36X/jlpupgFdoV0qgG
lL0qf3aKX1ns1lnafHS7KGC74XdZWwV4c79cQ4gK1kJLABLEDo2jM6fptEn1
XVIT5wz59HpbHTfOlvra4JgaH8r7I3rZAsApRRkBxdnHR5klrGLTPQBq9Fs7
Dfu4IG8v+7GDV2bEvBLiV23oyKe81gUnc6+0IF2a7NsyYqgdSn/bBiwLbrBo
fgI9cDDgkTn5WE6YDwHjko9PIAQJ0caPyfqwsNFkjVP+xUGKSIT54Klp/sh2
Z4Acj1qcQKC9g4Zkpt7LZ3GYWY2ZKIX/QnwMPFLnrjWxeb4GZOQOpiQ/UAwP
WwLloS3E4xRdPPRLQdsrLXSvIuo4typagLwL2XLvrFqOG1eg9U6+nors5oG9
pEW698BtL0NPwCnIBOdThEfUdZR2Ee02C3CLhm0/zr9A75s3CZAILLI7kW1f
NrJcdMhCjvX272teHptGmWgGyz+QZiyEnD880WHuaO+/z1DJdbG70/TWhw3J
ZHBTIF4UUgv4wu6U4NA9FiPoaYmzjbsgvH2v8nmewpxmSiEmDMboQzaBhkGn
wp0lX6INPksZIQuCJMQj+0t6PfgAvkmoGN9LmhM4KxJMf9TcpQ/xXhQoeoYV
CD1ZgMq9TtciTg6xtPnerzGIfM2Nr4zj0bTlk5EpwQdYkn5MYPvykKi0sKUt
UMdK+WV2pWVGfqwSHydTsmmuWomtIHqsi0/OEjiUT2t1AfGvjGoe3WQ4++Ow
kda+ELOur1gKzYe/XRiUHDQDPhClhmBrrYnuwNiJji6qIuYup45QsGhUFrhO
YewhPH2b8lbATVpLe+0F3VgW1cq+Tdh6wg6zpoMgLLcy7RpodCKF83n76Lr9
M97nH5FTEnRYE8nSk6CQAGVh5Fb4tYZuNDSBhDfvt25K2UzBgFOl4ireu3QB
Pxv4hE8PR7wltiDjEIHGoCrxP0xNPpbCKsg9xad8/WbFuOcQgbQn9gvf3AGC
htMeUe2rsKAf4jDqD4IiiEDwme8vu2lt9LYj9nAn/JHB6BVgC3W9JaRxiLVj
KoW/y1gEKG0STZ3H4YRm8c+3zocBh8qb23RuITxc8CD90kd4q6E7nmntcLHi
V+LtqsG1qNkzyQwRQM75+QsKerici13hI24cBnojUKzBBUH6mVk2xX0GfZAB
tZhq1jsfm/Tq0FXL+EBonTC2zFpgePbYHZEsyCMYC/u4LdSiKVz4IaaZYqCP
wbyTHZoxYjKpABQCg4ZLqSQjVak3FY6p0mZQr8bGgVrm9BQN9n5oS9OYEfjs
dMFif1+V3RAdpeENFKkRRg4/piG1CXZ3eXvmzcXLxyAT5kh/D9FZrqHrh7cQ
RQG1zX7P+ydtA5tqu+bRKV9T9Wogv++rsqnuzHyrS5hbFIuulpQY9zpKettx
El6lZ0DERZ5QzLnFxRycc52xpK8hg4Sw8//xuIXHDoA6Lk6OLUD7TmwY8JiR
pnv7KxTdHTPaJL0EtGfT36pn046giWH8H+Gm0C0zpcbc5slf4kg37lK4SbHv
Z1E7HuCl9whhmazXKV3ZUP93K+btD4VsxBP7KX+ultkOv338gdTqO8+YT6sa
I6BrKNQAHXBFulBOz7SIUqUSC6o2tGWL3jltApTm3c+OfotqKMFzmQNjqT3i
oQwDoyLTIPIViVkBCyFNq2BFeouz/tP60jBpsGIdJAv1rYXj1yYET873EWlK
ObMOQCqFfd6QdUr+z9WJFB44HCzUHfodgYgSgRJVOdKENGjU2vZfHskz++vV
iMmVNHyzz31juGjRwuH/O/bj4TE/BYY9GKVAyGHMqlmHRTu4tBig2pONg33r
GoBEaILnjj27DcghPClEmKZC8/051e/1bZHbF6YV8OcMRtAHTzvek5KernHW
DPdKLjmoWYShwl05PXjPN/3PTboQJoixqbDjYPKmqDOg/Z6tS+tP4gXSdY3L
roV/UNY7EWv+etfZhqw++zhSnwU/i6OZR08aR9vk6Ud10xcZVCYX69otSORj
mMZXgu8x5TGU/vK2/PvPJ88Mmk7gkh7i063YGuvBwYGQ21+EnWFsFspV59sh
y2t34uB49Es9hwPKE9o9XCeSy/7yMatgjx46+nKWr4Mv8RBg4LhsXgeSMhjq
2tu1B3xQq6kpyeof9gUaGb5E1v0htserrKnr6bZP1/33phesh2ubDhiKlhem
6La/tLRfW66OlE5ewF6/aofQc9pCDu+bt0odj0qqVjfk39LFWEflx2h9wwub
c9iMZtY4Dys6SjezwqPiGr6kfhzLoY42+VJ5ZCP7UPeJo72cm5DPCWbiOSDm
YEeY3rllIBRv3BYmBdnjOCioNdOoOjJxR2hx/ets5ZsCl5JC3F6LHVg9uZhh
oppWyAHnoao2kQ5VYowaJi2pTNAa7gru2WpKaxGy2DeKzbC8HbQVPLo573MQ
RQ4mculvbmShaUZ6WMmxQiCDj/NFobE5G7oqK6XUsVw1YK4w8bEMPckVyLuc
I3nsDOESHKiMkKY+YGMmZTbQmST7Yg8Qqf8fN9sHttAuWZTZ44T3Nyixx1iF
UFX7ZXCZJ5EXYTFunNz0yjy9sLKQeWoRM+YkDRbcyd81JQzWetRVBY4eV8uv
6a5LUEHHTXmpyrCSjAuEePEUxN6KGyrqFgx79ZZ5015EtSW16R6y+5YYcAne
px4kPPr9mCgV6856n8K/Lffi4WJYn5GjViGgqS+FR1656dROyiEYRhMTYHme
4RrPE/5oOwpawCwDEsS/Q1yK4kfcKrKPrPeQALojwTLCCdtYCebbldk/cp/j
t6Lu4O3qN4zetPuXwD/w8hr+4T/ymh+KkV1OUKEQ0YUTjXrGUYfLLEn+hU/4
uADxLF1HKQZtPBM9VkdHdA/eMwAyIaQUV1ZpTXDIpyq7kfqpGlDpXu2rYZU2
nDfRgTx/nXPOPgr6g1MyUW2WjCJn5HGTthhg90zT92g4N+IFBdd2wiMG2MJ5
ipWNCTyCfYWx5lFNxmtlFuvFSbSws3j0NXlG2+CcuupIpmY9RFUh9K2WTrI+
aJAJKIo9BsEZ6tc8+1AIHnoVjrP5ai1MwkdmJlxp58x/lKDY3y/9WXgAdyOT
SPnwKVvYjh1kXMmsxXrkvDeibV1tTvKUINjvCaJanrgVfaVdvLxRohDqrryT
a4la18fWi2/1MXuI8Px9syiUkaD5mWo5dSC6hIqje1LSAqoOt56U1v2j9tGO
V0oyYbMZV6VMBPI192Phzq8NZKNt2tmW+UU3V/hgq6mjkEx9CWF7ipWERjPg
xUUPJJKcyem6Fm8zlYHugA6zN+81RDBefkDivS3uOOpRsyDK/vG0paZERyII
aS3kQxI6welNblj9Dd7eaScnQFKa92UH76vQ/x/Cgd1a3wOinb3F5ws7Lgaw
+Ln5WdoJuhsRZh7MzaiUwulXOd3RFWnd1bZ3O3DhitWg7h9+XR6gzPSRlt9c
GXF0T2jlAE+8iS8Mxy9RLB3QhE7c8r7+cXzC0JZn3Fcj8OXGvp6I6U19gUVt
et6cCV6AUEzlAmdonWtZpGbI7yAu2JNk+b9DCE1p1apLMAzNGrCyTP8DAX6P
+hc7IXgXDqviyr5w33AS4RxrD8W2BUqZUHsLR4Zx5H3T1HchH7l/M3FDoq+R
W9YVR4H6fWdWbcKnMoZ+XvnVcfjYoDhSKLblFjIwfQLyANDFOUKGsLPQyMPD
Wa4uzH+zYsKDVrKELWVd5NWxVfY9Pqzl7Bd3gIXnwjUIY9CPkUxckTD7eMHC
JQs3xbuttb2R8rhwCOXIMh5+QjZj69k4ssRu4YvxnnSd/GlI8RzxnQBl7Es2
gYPor/75zM7r19XMa5016KjzR0J8e+bB3XnZJDefeSkvN8vUhT0WEQlZAx6N
nozALE4aV46uTcuyAH8poGwy5VsU+6L3gDkR4qmlVQ7aDCQSyTPj3te0zIwQ
/TnVs7l7MEUsuAc48a4BleLp2FS1OMXSJmTMmKRskoqDCOdq9fbjb7832sCx
h3AQpPmuDWUMein07/6j5nIwJKfHe9Y/8DToqznZ22TQUtc1r6OTD+FCyXhA
Ukfa8ejpX5h/DF/6SbLr2bLMX5gDLqPXkbPLVoe/LvOQLJ0yjnv05xYvDYoe
m8JrqcuVCbF62c4tXh4RJAb87KhQJQrvYMXB//wz2AXJ/JL33vt63iWjjv+4
3HR3CaILQnoAuFMFJXLa1ZoWfJUQF4vbJcolqIZzB6M0VL75HNX6MNux9TnX
0Z2gLYTCv0U028Xo9r038kQQIZ2tYxaWboaGsd7AqrRZHH1Vacp+26oyuHyb
cu9V5EodSFJXMajWvBpbJMtpxa92L4HhtkO/6zZSdBL8J4uoJtI52qYmSA0A
aw6/5C20aS/rZ/lSjqxioTbprJJPPxBUVXGTm8mdZYYQQmdtvA84WNcK0zL7
r6pPx2nKad+p64z1h5ZpoK9nWLB0w05tPYinBQq//vqAxkwQi0yxJgpaAD1A
8lgTtjj7V9C2bhnnQxepqY6rmSmaCLYIEP9fSCHWrmlHwUh7Os76JkxAcsZX
P/ht+HALlVjp3bsa8TOWMvUwnDcEZr6+5KsHzm1bxeWXOJuQiO2k3hxsTJby
nQ6xw6bAZElQsOXpc61zlvYPe4is/jbIVmWFDtpt/52+AcbgJuuyVT0zHLFZ
VCI5k7FamZHSzVSYq3lyi0B0Mo7/LOVR84dqzBjeA+Gd+rfoZgf668w6sdQs
dpBqvzuhHKX6xDZojCLkgLGLDbVqHqaovvCHK/UmjCms94cDC0J/OVbRq5wV
RF6qZB+r2XWJEy3Rb2latbKI/Ivk8JTdpFE3U4apzoPfiUSmHlkvZFnsV10v
c0LK4WpdY0MkCP+elHCHRi32jFnU/IRrglhxKyE2mxF+AmE+5DFJrHIKF4jy
uzlkpUPV1tRrGYJKAvmQDm1B4JisJ5+jCCVVB2tLrrcS6JB0jt5GkdllnYVo
hmL4SpStn6mblnDOk9EFjrtpdIPNdqPEhO62c0V1mIk3/zslm9lgKjv5wSAt
pmmsVzuyb9Uv8vsg4P3Nq+JkBiIz4OQHH5tpIRL6BwcP7kBoLlhgYhG7bv7H
7kupwP4EVj7MU1bNh1vb1IaqQMRBLfkHcKX2eunREJpd1W1tHo0NPI/UXHFQ
hmA0m21pNGCbKrrZGf7RBvDXJ14kuTWpW/KRYQWKnjhyYUGSHquEWgmCZcNW
mX6hHoMO2McnBBKSu0z1AEIvKNSyk+Np4GuU/ytbgTE175Uu7S5asdyZb+He
kxokRJzKz9SYlv+R7JO5TUfoVDwcu7pp6bizzY4Nyvr3Fq6I6LYxd4yTrftY
7c28IJDge9+n++wmy+nMreX+/n45nzpavovxXDvFuKT+SJs1af2/orRYCCxn
n7iTtOSTvd9LTIZ1/GlS6V94Ggd7NtkWLL3WTAdQ5Ycs6A2iXFDdWHEXYjVg
axTjXrLRgjWEpsqlVtaD6ZYKOLyMZG6zPNcaW1sIT82ob8pJ1Dzv5biK9z3l
x7nPB+HQ0983WWd1zHXup7kWw7LP/CbaWZNE02lNU2gIFvm9VVfSEaVfsUfq
++TLGGWVD+Cvj/ClMQ9yZQMe5lBJFURNjnHBxi4nVBxEtjdY+Ltbzq0s75RN
QLqoS6k0A/ZXlZT3SG8fHN8kcOwvqpGTPNTbCekxNTFbkcFI0Dn26ls9LCT2
t3zvgXlX2GNpJ4XBrJeM00lREbT80Zw05lbaZ3l0irAW9gj3XtBTl2Rx0VS7
CUe++cF18XQKhnR8HCwQE7ppwPax6kVFF+dp7N1fiG7DNC5Eo3eiTjNXSIhA
dmbuCXzmrri3pRRjSJXLiScRM7jO4N0AYmy3ZF7+wsDRUqg592lnBk1KoIRm
dYXlyYbcDbJbQVLfGqiZXOny4ksfxRJGMlJz1cyjnnoKBxCaaSwnPHzC39k2
xRVC3nUBizHRlero+T+y7FNYWbgVRknM3OTUGucDicCGKok0RLrb2/ugIM8M
BJyxQIF9FCNuCsNCVmPcxYKZ/O4mLowizqO49XcFrgfWEa+O1fu+FpLZ+Xw0
NGahri1mo47G4K52H3K0sqtRK5p26Y/NJ0XIi2fPDPhVnhhD1PgNcbx5Xt6W
CHpkSE8EVfnjxN9V3NfFoG0oIG9NFkkNLxLZgOVsDTF7qZjpEnHDkw9ayiqt
LE3k1uIac3vo4Je3XtaPWMsYEvNe8GAuAFfr3eHZ5P1IB9iGfRXOBFqhq+EW
SyHJoJB/FXL23DaMFHWS3PmCV7mWjEvcsoTd2baEk+7OncmQKIbssi7tfCQG
E0uQVt941IFkXUiD034VQ1SMISuNJ0mZDM8h4/6AA01EAO6q0snrH4NJCsBn
8Ophf0RB66UkLP4a1l4iG2EUEkBVdcfM1L/tDMxhq7JzohCiEA/JIcdI/ViK
AljDK9e5LZygqpQmObs40grIP5ifzWSXH/lsQXicZq7H9brxI1wrQGG050fp
KeZ8h4+RlKNOcHEw0eMYAHSjuginP4Xb/ufWPSCxchlu6ub/XZxCNIZaWjYv
Hw0EBRLi2TnQ6QhzLmW+Z1Hj8ZpAR3tkVvueRzcE0WlbMqJofo28CcyiaQCs
9q3Qisc1qRvegg95l7bahFLyghihUEom6DD5KgpCEPVCxUnZmbiLbF09w3yf
AuPqgUl1jVLU0kZb17ZaHKg4cjhvTK0YuiGOAn4BZ4HDmQpxFFcIP/c0LLPG
JylrZaAmZs3d+vOixCeuL26x0UQY5oGFv0MIKOCg5rBhPZKaYUl2ZsIIY4fO
H1QaR7E0OTXmY8qNqSlXJSqb0xTFZHn+TBGWAO/VZ9jsYUhGLggNYNdlQDpf
t5dXwFs8j9NHvJyF/fcwYHgyQ+bb7SHaKsb/V2DwDe0z5tsRmQY3D0vcYSXl
K1MsbxxxZFtrPJUhBBTor6yf44l1J1244wPYN12J6yFFVMzBQNgy5KdEfg+E
bdRMieTgTh6Q1VuDKEKfGKTfKZuA1wdhbx//1X0E2sBDFXQB2Xy7D46wOV6v
eMqmZVeRs8iF/xaemsHB+F4kXxqypuhPOZq3m8YMStVOV5gM8L9zqqcPKPCa
Fgnl6huhPmrXyGCdI4Vv0XxkK3Jy9pgEqzPE29SNe8kfV7sIt0DF837QPI6J
gZi8dCCm4++yLAcuPYrf2vPhLPjSccnepZ6IntH4CEKeWgSUwIJ+i25+MZuy
AXs+9R3Vn2Md2x5F+ST5tpCBvjUk4AuYmPgmMa3HwvY7WKX/fXS3VNYFjJ+E
IFnQaUBZ53dOZBElnThs2EWkzXlYSJ7l5CH5D0Losy1kDi8XRORoFFJOW6em
21ns39yWVrnKLQ3pk+LPe7hDddnYnz4Dko8aOmCLixyIVLQoy5ncM6l1DSBE
0M6jvZxWL2DfCRhn+Q1KRfbEX26xzZIbfY/Jlt9Ni+NIFiW35N68tqRAJ4fR
TPVB2iW/BQGPuepFnQmKWf6L1PONzaF2egA5s8v03ESOAW47ZyXWI89FpL7V
+NFeL7Ga2rmiAP640txHquU2kRkppmPX8Bs1hsTAPmwjizFVFdFOpfHeAyXC
TWIBFiUhaH3/t7bPu6/ARUrs58E2YJfY9qnukxtM8XFs0HSf6o55QTSZxs4k
szZnvFE6B2RyPhkLcNCIsPhSX7jkbevc8sJYz8Fgs2U+DoXWKkavPVDs5YKr
1ZnYtGQo+xy/OaWoyWLcFOxXr7qs99ikTvylyKEtbw2nci3N9m8fpVpSMXqL
Esrb+F7CULHL/TwClj/Ub10VLGldmcUPFzWcezDGToX/U/jTRGe31T1Wd6vs
AaM76nHBZg8tRTrNJe5Pv7zBc9S/XT6HqgbXh3EyTa0ZfT9slMMi0NZxpqsa
HL2DwxLLXr/QlOpB7Y97a1QJ54FdRJIv0WfTPP33UpWskoIEQZCGumKN+8jQ
wA4rcDKOY2ZyTbyY0kbTjjYzjS497JmAi+cxesi45mDM9xYIhzHlta8FnT7B
yg7uzszGUEDttSU7n3JKf/XFPNfInTTvfmaHslu1xFK35nVFrKuPSxg2vD+2
gYM9Y2YCsW2EcKxNBmADePFoxS+GTmpSFGUly7vK+3uxxqOsFxKAnVA/WG7P
jzuoROHH8PXBapFlT1gagveenyYpKr5QoRN1vQJTtbxbafTT3tONEu7XTwa8
pZDvUk5ZaKsLR1aOWKs2N0EROlA7w9ZoFmqVm9tHZWQo1Lm06smPJOlVF6f0
Bz2BNB3TkEXvbspVTuHtPxgEIdqGgLwKw82m2FRUCEDeUNi8zAn6gB3o4WXq
lOOBi9pxwoEV5BLU6hzA6FRuNtHPgN4CQC48ZSH6PiAiaNRC9X9d2jrpTF4I
76H9wkXGdGrlEggeAunfUwVkRiaCb3ROAKLmdXIWdrBXgQKyrerdOcjfIImn
mbm82f4ntvu2IkM9AhnqlaLAa+MstA158SPbBnidy9b+XO81nNB4jfYKKkXj
jyAhAzpODLBli6jUpcfJiunbogVdbbiaH54fm7+EFuQePPQDdywaDf0SQTwI
DWJ3jjGm+rKDW/90kGhLgBcFE8fVFXusu48zHKhnGZR/p95RtZNedXelW7MB
eC8lv/beXIJPcBiRBAHIO3WY7a1UWoozcnJlFrtEEkkYU/WgyCLvaERRJkKn
4dYrNrFQhoHVJUgTDluortoueGQh3l0gEFpCdboNMvi2s10bL0VMdC+imgQh
AkesCUQM80rbgHMQYN5Bk2/k5a4yFOF5mKrvJozacN+v6zEWKF+aKyaVh5M+
UV8q1XcIDM0JqH/PUP4hi8kXibNBObUc52qc3a1kvurtZ9rluIQ4XiMGU/4v
k3qXI2SuJUJAgmtzr3K7HAqtDewJzkETHckQdqM7UZmxjYiqyaEt/6aXN3Mz
uk8FMPnl8jWgEWucGlCMKb0b2urf4zi3f5lL4AW2Sww8Obx95IQVaDEajC4F
q93ppvF4rKA/GbhGh58F3zJrkg9ZxKFRsrfLVbz4kPPWtRydQ2LoY7WNg0ga
B/VjMC4WHcwmD/NEcWL4IgmS7mWe2/MM+HZFR2WY8fXiBci4ANaM+0b+gY8n
K6Ql3qv2QCwlsjr7CJwP1OTKyWYFnHoIRC2uzLdTm+qY1bDGsunFg0rGjdgt
auxIOtN3dcGjB4NZPXnJygTRQGrN3U7KyNAjFM6ZEMsEZumvTKD9XGjxBCAz
ezhCNaSEw/AiaBqDmmpCixP8MvCyIhNnFZLLLZTwWlruEbyACvjS6xWUchBz
56TSqlfyYXVjhl13mz0tBUiWVlpxVQqAWtws+rVbx4XeUbCykVjY4cwfvqL4
4tZInBMkaOiP5CrTxHXKRJnwws/CZOM7zN8nBcoH59y5D/g5RSrbYkIrQ2d1
FbGC4OMd8oUL0d3rC+Fn5A9L4DoP7c/AnsOHGZf+uTnLhz7bFPwvQeGPU7wQ
vVFsEYtpO/ebpFsEAvuvXMImpo3F/QVdY3cH4UYMmWmNoCo1Y2OspN7v4JUV
a80Omi6w99sDi/XGBDykpoKMWycpCBF8CrO5bmhmWlifjk2utyTy81RyjSZV
MWQ2Ft6tYUiYxH1w9rghsbBbbC5wRzQT7OW21VnusbaGD2PFivZh4K8ovY04
ZKens9RPQmEPEOie+iTAzUvd5RRHysjpZOJlygvpS5ETEpO/Gf/xxlQrXAnc
hhv0wQL/6BLqdnHgcT610z+2hoR/aRW9vWe7zPLyMUJCB7D+3mL2zSMcpQgm
NKUwlHEd/VdXubQ5lV4dWnkoCWdQG84D0MLyc2QGaG79lsnPOCHmdaZfX2+f
LU8QcXfRglYov5ehytZS52iy2PJLZfeE0voWmdZ9wwerJozJvYeyQs6mY0Si
EknVso5cfsaE/aNjeGjqMMcZsJ8hqPEBc62s+QGj1TlHjjtT18L966yhPh3e
IPyFIeu3QZyRlb63/JEUoMVlrue1DR5FL39MMaIUQlXNgULD3ubw8ywT+JaG
BiMn+A6++u9GnejTNhmL4AtCqla3QR+RlSRtp+aDO1AJTKbGjR6PjwmeLdZY
BE8sUWKcBYi/yFgu4Cy2YgU7OM7rY/VWydROYErX/8tA6ZtEJxscQEwmtjpj
FiP+4aIJstlQ6htS4Sd0LsImJzJCcMIKIpplfFNiXGDt2ZOq1GO+cZLcRRfG
MFjQ/7S9z3bzmUvNQVASzYhc941uYiKx4LLG5HnlUJEURdbJkxneikWKCsuT
qpVz4aqS8qnRhQ+xeGbGSjccY68RpNVjK1AKJ3j1SgzgdsJ7CEufJAfCl15p
ehwhG9olhqJjljaLqBgI9uYTlvTc9Kc4SFHbHMWXd9LzhjXr4NU2A2e4BqYm
uh8/VDsfLCJRzIUABjF7KRHDJN2eWnqOO55aeWLgheaZVPUdstl7VIgw07wI
N8I4x0O8x05XVeZ7arxkgKsEm1nk7LeUvo8XkwVnHrF//pHFF1G2wHxCYNbx
yB2dfHOWAk4o8a/PrbuNJqdmKMRPxOeQGIrt3Cndh0nhPUxrf5EXvz26yPFj
JYxAkgvO4au6yRQT7vF32BbreIy0xFVjZRkTjxDFVPKY5HoWVgNusrkQV9bb
Tjn4SnCqkF3mmzAt4C8aPEpEVWI68TdeX+uph3LH+OwWNbNj76p3Wko10zqb
hU8IR1qcq/r6I95esMXJ9wwWZV0cZcIHC5Vc2b4n47d86oJO5eyFV0JER0v1
0YJlEG1fCKGI6ky7t5Kwouq3B6YYwpZ6xYh6Eh1FC5yL3MqAbEuDqdzBYIK9
VjdvxIS91EIa7iju0M5ECmdvzl0ftiuR0rnPX626nF33JzM9784L9G0HkOOi
MgaduYK5GMHiI9MUgJSON9UsmCDiGp46ktuMdMzE0qRDS371pivO1Kn5JN/8
NfJZUNNA3wWXVGlzaVGdzFjMHonFQLhmFWz8BX7BijaEhAVRpoyvmDC6rD+2
MAe2FN4K8xfOlBJ/8f63u/wB/rOQQ2gsqJDMfxUAPezmPoDXP2ED0m7yagFP
E1//aRmLyXRCS3LfzwxS8w35MegOFEofdjL/2XHgoyqu4BXstHjOTMuRt2ln
jzaJNjVbbCiwiC30xxrF3ME03ceXYdkTXUCx5gWN769IIwZFMHusOdfdI7tp
h5nRsnmauw8Zv6Bii3pZdEAEjPUkEJeP49j9EhQf1IYfZ6K+9Lfh951hXraR
nuCLWnNa1j5QhbcbMuX46PX3VVzgXlKUExkN5MQgDXUH6cckZ/AVYUVmXzo7
KDM9rBLj2mr52+KbeY8afDk42p+M078Sf69VNCiIfmPqHb54hPdR1m68ZECl
BVeBCVMgBqVk/yxNQRPRxGWzNQHZSlMjzP2pOXzcPgZrReZlLlsfzkDqQ9K5
MysCtoGKPep470rkzwa3iLrRTmCE4Sm8lyrff8JvxOibbFYmB/E2mXqBdf3P
aMBtNbml1vOoF8Cwkt7wCrggV1HFwKDg6+/YAv5skYG/sPx9NUOd6l9XP7Y2
yvlosylZf7GghknSrU7B/bpNTsw3u1YjT+5NsMw9tntRwUXEyd3HXF5YMkuL
Z+2FGWtevlGANMQSYxW6DdYX//KtabkmFNf9L/jSl8iTatMERx8qNql4mqi1
kfoCyUYu4FJ7TO9+24mzTm/fdexI8I5VpSElZ7VK1aIhhk8YuZARex3INx6L
hy+M7G3i+or37tsbQSNbKFfpl7Wj2rPs0PlZg3Y1noLd93IRUIgkUNhaRovu
J95w92mlew6R/STCTIbLBTf7XzBbcTWGpyxlfuCEj9W42bp2mKKQVOYZIGhg
Zb/VTgGyaQs7Fy36atT0GxCZkeJWEaJatE/gIMrinxO0qVXhctBzwQwsMpse
tJ4BQgovTS7YNAX0E4+8WbfKjD4bAqtaMaoaCxdfB1azSRcjaxhDri6wodMl
hhGano2ir2xeGBrgHZ6lYDrcTwZWXvfIN8UN5nslHuFYt+YL9VQAfUAvSUeB
/DjTBG8bT0GKt5s2EjMKEuSowNDIRKgJ47lQebPGVHd8nsrptEQBAZgjmTtt
c4kW1nVT8PAQjLk+2SBLdqxIANBYRyKlfJ7bp4aO4kFej5PAY3liT4TgLKN9
Z6bElp1aJetFdCeU5gEQXOoU+tho5WmYI592ASdQsOWh4Hz9v6xuGxhLtkTb
ygAzIKnVHExEqc9F0+ripxW7WFBTI6h2TGOnMwNrTUSl2J3OvO/E3Y4/QOPz
hGLKsW5rF8c81MmN6I0dlIWx5pRwcX0E+fmCHaP7bVK4q1UO5DORYhf3zusM
2Rppm5g0nOyRw4tXhGqgrFwcMxb61yQc24vTm5Srj/IWasB/dQRj2fgnyuhr
V/KdazUC7MUBSEA7XrqqiY/UVLfCCKhRRYRSdbmXh0KCSKxxkHS4buNcMWlV
GnF+wUAWDf9pq1I0Xx0ubRXCH518qWuL2b2HAIWCyDYnwHYVm8rMkwK+qn6R
ij+PIxez2MggU1bPaIYBJ+lOwnFzOtDC59pt3F2Ai6QT39ZTJLfOuT8AeuQV
AcKuN66VKtD+BRm6KNCyo1pcC1cHlu2IhpEXJODMwc6A9XIM+jILnHaL1gBg
HDAba3e/eQ9Wd1UD8JvOye5CLeqr5KQSTbTT6RqYRoUMXEQKRgBeuD+I93pm
+ib6+pPrWQcW8K8hnrxKaqILXr7CKLWZaRzfQ41SFjQu6jpofQl+gbtv1Nhe
lPH20VK5LfuaXx9X6YSld4NINni92IBCIQZeKFJVKiK/s72xkj8iXWJ/Dxya
OYmZ007oNJXhf2+bgcmxVvsHsMEet2KM8b3q0Z9b8LY79AMoBIq8bcRr3f7m
mJwdHHbRG1L7zty56P0gZv5qRL672yt+ZWQj5Pm1s/pHNCGIrWmczSrEKWdp
bz1u2NrsV3EuQ7Hk+nwqaK4ZEVYm6fW6RNuWbLUw7blIx8d5ei7KRP2B/T53
BnpFt7tCDQZnd6tY71Io2/+QhjIpq3tRKTzDuTWNtjxlsPNuBj99NuGiR1Rp
PpZ8MFQu1PL0sI9Jk70+FcdfY+rZjsFxgQMPEoWUEC7zJ1xvmMEGTobL7tyC
mAIQQDKTSkOSPsfbeedXjvUSWltQQH+soXvNAcPjk5oUtaDcVeMB2pC5057E
GmMuYCdoAy/IDmEOjVpC/qQyWKWpW/tgzYdY5V6HPG+Jlt8rpvEWNlm1PpYw
wH77attDyyBk1SyuAbIqrZvQLMwaYY25uLMjxGzjJRSHV2LgzKXgHV6OkK8x
CIgv8bkEgUvSGkN3As1z1/ErQ+urshj+zNWweAyJTp5lJ5Hjmuy6fy089khN
M8suUy1uiyyd6KW3grfGvDFiJMGB2Xao1ef1KWo729K9+Yl1JH/37GaDg7jw
8tk581FpmP2N/475mDFYEqqRE03+Scknihbr7SlG3/iv+NQ5JrjSi9OcxclZ
N+YrgD1moEO9MlAaRJSEs87FD9+NeDBF21Yadgd+IP2lHv2vCC+aAqjU92q+
Ii9YZf3eFqR0t5aYaJSE6GLyCue7BOIc9u8YwnC05yUIVHv7Tnb+GJcg21yg
PVxZnF6JCuzpngH2iQgogayirFogcv8zfT7mOUUlakbVJhu38baWEZ+MYyL4
Wv8jqnihUos1ZG4BO6nG72+FubYihMUZSvvCLVxJPG04rIo25DNSLfbkmgNs
4bjl/1FjMBSgpWcL9Fsdj3xS2C3YeWi3eClURCPX8yR98XtrIBuqgkFCIEyM
F7Bkp/Y+vLh3JU1oKfa9y7Lfe7CPTkM2s87OoBQeGf3QV9k57C45ILglH788
zadYKQ1Y6PjL6p/rw58mRjWjsW+dIigLQTyRO2yAEO/Uuq93EmGz90VFRX7N
uh68kY4v8ln/pjBWf+vdtUZt3ohb7oi3DTFHk1PhCGNUgGvokQEtk9XEx0Q6
EfIgH3a3g8j1TU5r7dFEwg7dTSSglZgu3ywSU1C1SUgxY49iscUFKb6JLXL8
I6AXjHOusLca110v1mxMT8azPFLK5Dv3kWOQPa52PtYRFVo2NrcS2JISHbjb
3KMCMEUXpeAiwpQ8pwwcK1swAgxD2Gwe50S6Z124DMEVrAySDKVKp4kj94PO
r1DtE3bSmHJb+oSYNkIw3LsSv1nmAgOKdPCn1GuPpN1V6Xyb7ocbl16VSXu4
KziRRGnXhsJYm1stmdO6xVZoN7NGkX6Su1cFN+MivdcoXoCA1SIukdLQreYk
Qc5H5qD58vF28dUqZTwicvcjRE7wgpeU12X9gLtJAbX7inRkfnZF/TuxuRj1
BvPDPXtA/mwSvXa3KUhW/G/phlqxAoEJmfgkFcR2caglVEDILE5esmzHTZu1
9biq7aUe6RQJrS80O+CqbMgdaH5iqZKsl16X0YRCDLn8bs2nKUT3a3rI0V6w
WAQ7v+rlow+bUHUstcsn0LK9ZfJGvNsGWeP2S9f4e++ssKV135G+7wu5mIcz
1VZhP9EaW9G/N9RGoPA+nWOb0rIz6UwOWKzwUYJ5Vhv/lPkbNlCdATxEdG6/
HE6WdH1GKU7MN2GKK8ksICzzD0DmcRNJDZlngJAaqrs1S/djcG5ceGo78hO/
GB+li2CauC/Xqa4zGTl1E+z3lfiroSvN602SEcag9Da/SI8QhNZup+21y/h+
tb7Py67JRh3bVgTfSP+I6IuHwXzsT2sLa0ohL1p4f7zOdRFy4Kp1NBHy0Nd7
ZRSqGK66LCYuEkF5w8KlPRnJwj1k4l7WS6x8qU9vtN6dIzda3AmY6Calu5Ta
6TkDyxoSwuJ+XtILvTma630CDpra6NPrV2ZuSswUsWfDlt95DD2ckwLq/33J
Vk5Fm5+V+4/ZlapqHEN/CqagNkn0Ld47pIh6vDIiibTFxY1yZU2Cm7Du7HvT
ZO08396i8E2AMu1c+8pK1GgpLoN6vry5G5T8vz+MSL7Kbog0/nivHyYObaNs
JyjErujwzCaG/548OikMTbZ+iICqTVPdiUQlZT2dERimqjpIPJoGdNqt3+jK
Gpbaq+tadd/sOf/2GuGtQMgfjEPqGZuAu/gBdDyXm8xK/T1Cdr4b5cyMfbhb
szkwGJ867rAJ13CO/Clgztxiv8ue0MIOVb4dJNDEL33aEw0gR06JMVZc/4Y3
ASC196C6B1hTvA+JptyQqINWcn1O0bXRshXz8cUz1c49J9onafVsAjxspt0I
2BEoglsVp8p2qiNlkisyZiOidAiuqWAcrZ7zLW6zVV8Jum3+rFJyOlsAGzeJ
X+6+n7BfePFlxfbBp5m7IaKiyCJqNwmbTUD5G8j6ETqsi9pS00nfmN2PVdD3
80cETfCmp3oOwWUkn/MYJ00/mgPBglNP/qQewmO8dAF9J5/COdTopGmfHx5t
kGf0r1SSHSy9lf1YozpsS2y6iwUkPGqytx2kwxygEKBYn0l7fGB+yb0+NEDV
r0+DxP1jp1bOcpIXWeeQmUXTr+40CTNEfkekuxup1u0qCVUTsI5LhwJx7GUB
iXFTUR8JWy4zVm2AY+xF8nRMX4rBnnF4ztofvJCKrz+XPzQ8IY4/3IDypmw4
eKDbmOmXmSeRZQWrPViSQE/QrScwyYuew/KdLmgz2YLwpHWi4WJVbLWqApDh
YWjIUquMD/dR3gxlR4TwUNPdG9FdHdL9ulftw4ywFMmAchdQ7ieGhLQAZlCb
nFOgUq34M/h3Bh0uEiJuE+y1954Gc+FlyM7tq34UWyJhxpC5RvKlgyzxz/ym
qhXqxgUaznVgpRwytSiui+VxR8lCJozrVfxdkuXTV75pfRG7BMCLztdSwfqs
IfyuOAdiupdtw2gZlXFisY2dh+k7jwUnB2BYWUCfFh3sm9skuJoboaUz921B
RoeoyHZ630MlbBL6WTu6sVF5rKiGuJhaz+Gg3vwDZIDcIXBDh9vFst+w23cH
ryU+65jeVUyzy6enSgB1jpBmf7OBT0X0XtyAg9BETARI0zFI8QlQUesAG8TH
84UBpzGi9o06/N78tjuafXBko5HZnWfUuaKMzdeVZYIlXnD4KOM4+LJUOi6n
q6XlIHCrCQPu125ro3OZRUrejr1jXVGlWMhEHLCC+M0i5aifkj/UkJzrOqtm
MvfG7WnuAMGkaxMcKuSMhzAphGXEsvPR9rxLf5vmHldM5NmXtyUbEt57iFaV
L+4IoSmIFyBbP7gjmHLjrtgCae1ZbklMBjN+UghyKR67LjxLjrdb/OSkynzQ
T0VzvFN99ZaavHNT7mgZMQUyTvbftivoxpbcPbs/PdiHtyHDkKhasfkEnxkm
i3JM/zBNE5zFh+bg6VXynVp7w3YBO3U2zt81u2M6zsVaYEWXTMqBkIxHnh7/
p4NfMNlrXpe93ZwhG+ywfR499004eGqT1PjaL/hfyot9/YrJ+/TE8FSYknln
3NTi7n+JMvcZpbLqMRD/vMrcc7+GtYbmUeUsO5uP1WBSbQ6v8RQs2sauXSUt
Gxr8LTCetJsJZt8QrMnnpLtc0/8enF5iibuPzBnWFzXIxhrOT57q+waS0kZ/
//lxtU+ZI3EHBhmNRX590V/XhT+ke7Y7XpqLiBHMr1/xaFo99r0LBTW0iTO2
phM8TsqRezlUA2cLzzpT16UVnrXvyco3wIR5PKulcjCfKs+qYDVSyI0h52AG
THpM/ml4e59UW80gA5lGvvisVpAz91XLdmfjypgnrLLcfh1NBkPE1ATb93rD
RcyNxcWIfNpTMrBuoskZJ0ey2zv5TXocRzNF28uZwOSBoLHZ4GFpzfh89nOH
T4rUsHOk+mCwejPFHJXR62kNlL3uFJ38wZ2PPiwt3fHq0rHWXtFbaQW5rD6X
EN+IRBd052Odp/yVXgFTesktqqqIHzKZnkAk0AECWbLDpiwrZjcI2yHyYAN3
7ih3/F+WNCVmnpZRuxqFEfCBVNYBLBHYYVZvQvXwpUBsYFUfbfJcd3kABg+n
q5tXrP6VGrYeh2gUmMzCfEFLY45G2wTVScS8VMClK2t1Pg6N8ScYmdYiGY6L
1BsY+diwbNx4XFSPMeHrHUEeI25L5Gq1aJ+24Hrl+P8wsroyUW7JNmMFbhyu
QBlqo4DT4FxSzOZoiRhs1r77fko44lxEwh8Uv0hK0hrIuM1q4k1E8zIImOy2
W/MtT44vgdP/svfg94E/9pzQltA8kIBFBAR6F1pbEE37p4oMw+dpI1M2Gdhi
mEkPfG+hksaKrv8rBdplxsiQz6NYaRWGu42uB3tz6Yln9ImciaeiNpqGCt2j
HN6jDxlXFBgQL/9BAvSKZIK1WtoiRb9oqPOkob0uYQ6c+OMTJ8l365VU/qvw
XEz83yPNtrZMAsfYKEVzHyqpNi35RJZzQr+L9SNBg8dVqal14u5kEfvVXFwO
Q3zz5QWFRXFX16SZ9sW52a+f8kmnB/g7Wf+FV9pD24S+W9XPJLKe8+sn3IwY
7LdM5GmteVTRInaPD0xH417q3DJ+OjwB0/VjEWD5hIKIvRAOPRGjQgyZ5HNq
iZwSUE4gLC5360QVbAy0Zb1sC3mmwOxh8a6l8B/LuniWPz19QY/F3sKJX6q6
lcJG3bPPg7CA8cbTl8mv+3XHbLqccTBf9YAHTUEMqZa9M5vCpRPU9McTU905
k1UmdDVbUpvI6pC09CQ471AP8j90/09+UcZ0LRkhby0LPtflRXHxXTKXUAaG
0jHZ/GpVQ1TzfEGNjgQDE4xB9jNo0lOgdDDdRnrjWdZA/v/PAoQGB1DkDJ0O
xfLMqzKQ1IacVXzhD5FVuOZGGg5bukpDfv4/jkuhCB5Mph0UkAQ7JtBZi0wp
rAzY0fSQvrHPzZcQ6y8y6SGbj3kbFxtms7vMe8hKjIQUO08XVgQ9FhntdrV/
9RjVydetWoMp4IjYLcQrH59Ag407lS5yvVMTE6skBoTSjtVlsdRFDXK49VG5
KfzAajZiSyKa0TDg4z/SxieXfvDOMGbugo1Gt1GVXfujnpqYbg8XhhGjBDcC
q58e2kE9PUVwGc3/P3DxgQEG9LP5415nTyoWbEOWLkJqC9q/NpkTR9iyBoUO
O/JR0m72rH7d0aoFq3rzLOUmoKtoX44Yb5mBAGvI7W7Z9bdKzSKDU+dO3/Ow
OvdgaXF8eY80IoGUrU2zB15+LfLZyuunWJw2Wc+k8XK6XseSEZGgfUTZ2N7V
JOiV3mO2lziYuwcgK4ookGkgY0orENvknj+w6Mce1Aji2OUQf2YD0x2Xkn3r
9rO2kEcKTHGwtZ1TPRbFxyRIE8yuWxCMexBC9pg2D7TLoyxbgsc4OOylJvRv
P4Jcjqyjabv1B41aqImU7VXVaqbHyIXkH2V/EhjPvnYL2XZSN5RU+P/nK39A
vAMz2DUTvMOABTlDNdIwvMiczmlt2VtBpFOUzL8aqgayaQDbsEh1t/Iblhsp
FiBfFECBXl90TipVYcRXug2dbwLtozS93A0mt+GRX03dj/dcpoUVMfvBvsB/
hhylu/JUMJoM26BHGAGuL4DjieO9fQZ5M15+DjZ6hjagnIXFjm3wMd3FnLta
faHQ3kvZi8abwLPEF7/f5XV+3nKHPX1K3NIKFjDim+BpvyVgmrDEEBp6YvKg
N0+q+48vPigOCVU5SFSTkqeDUw7zJsF01WSQuP7CeGz8QLQUSIJWmvUbP2o2
0uFSrdUwF6cY/zCsyhk8XXkOpU8HjUD4w2wtSkwF+4x41zGXvqBmdeH9yukH
BZ/az2ENnvMBIfS6pUc7vh/1TYhECRz+VvuU7Lv8/KBGkKKDVWjjH7ScQDzz
84CIstsl++LvZgYnTwGzm0i3RjIlhRFNJUh/stmtbdil//gWklcdO+L7P42N
GK+WR2qJ3AuNAPiSa1z6thEz9CJ+u4gT2R1GOG/pWPoZps8FXydYH4Z2yqNa
cF09P/fDd3uLZOit6kJBMIbn7jnXk5JUG0mBb4+2ny9xbliMX0leJvo4d9uN
u+/b9bAPv7eZ3v3HBUrJU6IuwgELiP0q5vyp6x409x65TeX4e/etrnS58Vj+
MDha+2iYRPzFDhyeLaXMIeV8uCPEjTy+ymNHjWq/RjreG31t/pVIyVhgEHCh
ZWCyD6DXrrJtKCZUjE6QYiBAJ70JektqAAgmOByIAwoSL3kLxlOlLgo3btul
nEKsWmJcbTKnJxvR2kFcssbv7KJoR62vfFOZhGgc36JJWBh+yyMFcTLild8T
Y2+sHncXRnUfMIX3tcODMUggc+aBY0Gs2ZiHVvGEUUP1E3Kc74HZGSDrTLqW
IIbpjL166mt4iuA6hQcTnC8HfrbF/83xI9sQKMVR19inBVfHc81MQR8gE/V9
PxIVDs3ataHwBOMhm2TPrNfynmYF4aLAgZQ8FlIAvlWAlWkSLAh+iBgPPZkR
Yn8KguSwqp+JcepJdNzA+A6NN4d6sK3KHYmv4Uth0C5HAPIdZI/Yc4lV/YXL
hMQ5QuQaEK61eloZbAvL+10K081dYG0g5b4mBTeVQGzT7auUslQEPXcgSjED
uMGu7S/CXpQBWcu+GE7qzzAyOsEdipPOQQjOMXnNXZ3o5ZKKVsEZhszqztco
Z8HlmT0ly35fjlNzfxnZNxVkByydzEVWGjEnNXQ5mXLvxdA66YnrtOKZQM79
xj4T5tb4outdN2/JVI8jEvTRGsvI/wIIOb8UCvoq1uXQb78zESb/qqt6FFbv
4sohPlJhFoX+QMFABT1Q9JnZ0+EEOXuaAzXJwnoA7OIOzuweSmwByhy49tU5
irEZ+Wgq+s19cxIv3lciTFq0Jmsj6QXrcG4zwOtz9lrB1140SPzZAFwfyNcL
fiPK+gVGJhuC6/Dr9NP+72y2eYNxxIuHdheccoE0laAEmcLoBAc6b8XQeHSK
nnx4TTLIA9GX4HZo/xCGRMxMagFPAw4neiSwMJFo0dFmcnpcCl5GKChxYMnc
h7ausFwcocy8lxi90z7sTGs4p83QALUYOYjMyovmRzGAOOva5HyRPqjNZ61L
0AexCzLpdkHnvdAHBYY7aGKnoi4F+IibS7H9fR/3yZ9GrsM5yD7G4xQaKDHB
kNX7l/ZgX6h8WfIYnCWL0/lDhraH+fpQTdR5TAGS/G7pTbEZp8ALt4ooesSF
QMysTbGdmVeifvMdmtugKtciC1R1XEORWCJrHCuh0p7RV5LLWA9l7REzIEyJ
hf03A3S+6kYW83nMyM0bwYAaXWmTlRrJMO53/iBJ0b0ax3lA20i7y7XboweN
55/xJJsfIC1ja9RtrRhazfM08PtCUAUw+qG3R96ePPahXA8K2tGcH2CpGjE8
i/K9HWTdMv9z9sQz8E/yTsTZ0PXt3gAHTSPf9yVtgylen5aHW4C6KWaCVdZ7
Bmt3LJi5AykfRhJuONMCscKX8Oj90ZPOM3/0muoOIN62egfV5Zzmuihs+WPY
h4HWFBSHJVkzeGEuC+F1B/xa+iZ+S1CzntchCZT+3H1ffTe0EdeD/6pcvDz9
QAadsGt537NmC8H9PS7LWBnnn9BkyoajnC10tOddQUwSr8xIQdph8egwKte+
eozlm4txWqFcXkWNJlfq47M9PaF5hxxRAe3DukL8fZFfULgZmZatNdKcZys9
2c490NHBSJ1WK/JMfmltL6STl5AMBJPWFQmS1yqVSBOqwpA3bF8oYJ9epvp+
fPfsXaGV82OI1R960r4UU8jaC1rmDgNcgxb4ocF6da94tM00oDbj19T4ptm7
Quoypk6uG24IjIqA1QwPy1sO5BbJOVlLlwEGD02fTlnQjDj6clyRFZy44eQl
VXywoc7vQ/JnDtUuIyNdWaPomS3F9bbb+dtQuy0pcyMOX24jod2O1cDdXk+P
ym2K9vtyzewv/BLImWlqWVDxzNpLLyJ7AKJzr4MK4oL1C6TEWLeuqUjHwJzz
UK9yPN4HHri4uGbxykyiz6Tf0l7yDzqrDIm5V41NGY5F4tazx0s8q2cflL9l
6sY1M/D0nT968A11vqX105DqYHhAwPGClMCdIPa602gjZKRZLc32cz6Z19jW
xmB1gid9b5f1KkWljdwnydCPRwOiH0aJnMsbx+1tA7NUGMQUUatG0W4/T3vI
1+nELq59MavHysAZtzOfxObYvtepe4TnylWV1L1rEcPzeMwe7wMTIZdKK2Bv
wFB+H6fyL9HvFGRJWxeNGdlbOFUmwhrH+p+8Dax/TR1+ZQdyiAxYpbOPvcRJ
8m8SUf1zQjwHPxbmwPgHc/4cmWvbHXD32vt4oLCWxDDMwfiKiU6npKRWLVOa
Ys3FCN0w+PsbOwfIutyhTvZ4Lt0TmX+7rwZILUxHVOjfdyOcoUzYu8T1MxsO
LdE1DdNeYds9dCaggIjHp92xJ3jus4ctKhLN8vqinCx0pIPg1iG5rEfE5i1u
6GDb85dNz7Cl1GtmicavrlDcesF3jHEknJnHHzniYn46DmYXIdo9nml/bfQN
x8Q8io4no7wZlIa2VZq43ELe72Nt+weQlDbXdm2FuSKMgpW9SPBQtIisI2UU
hsyHBe+z1B40UakfHyb/A17mLTD6aZx5lFMmQf4uuAbPI4UlYWWYJ8+gJQwC
n3kFH6oJKyxmTu8ufuDWV8caSHOohnoD2SDfbBwJnCVKWF0ApNXMTu19BM4T
lQ3okupiN14WXaNsw1v7q+ZxizhNN0x7qFrrKCdo95KuzSYq18I+p9BzWdXg
0mPz626Z4eOGEdicfnWiyV9EEIx4G5HomQySnHAz4+La9QeuP9NKPhrbGMl9
EHjBOQlWxhJpgM9unrFkNIGFyxbh+tL2X8b/6O/3WXUpxJqrsSOkFHNEXuHr
x0K/WevL/L1++far3mejOvuU1DvpcbSuYOJ5T6UrhOCFMPIqGLO8Zl8ijYVK
IWsYF3YRumCAPLR+C/zPVMLBUSgtqcBb0p45OkcJ2a1YQyyLlXV4ZSdQekiO
LujJ6BnqPVRlR0ferozVBF59JZ+RwKverP1TMemSpKCRRi6baSgpt2GcwDEE
P2+7k9PplfjvngzVLk4p6AAjuovlHLAnDhnS8U4q1t9NYx/3ul7wIhbUdfSd
GIT0nit4oXnl6pnZu/OfPjJHsvAgcxLmdAe1uHLVcdHwd1oMSNL/waPGA0o4
1VN+17x3svvNjBWIJBaanbpoiSDzhZ5XiaLXxRcivZUO7Z73QnSKQFD3QOXT
bUe4dcdU2H2SbmGnfqy7lUH0Ys3BHWZn6N+mHCuoQuVeqmBSeUpvMlN/2Woh
ZxHVUtKuv94mA8LsuHsnWHzjqWvWF30dIm16YikpwZU3CBF14D+Ys66cJB67
ka9UV47fxZlMekSsmqu0n62xxMApAIB82JTjBzHo6blCmNPh/Ey7w4CuWEtJ
4vR4qKAk8MOO8ThEMwIDTABxk731UNKa12MhFQENtWfPZ+h/4ucpdQq8hJ1g
zBmxnrIYn8bYqqsVTk3aLPXfRAMRLGBnAyBKY8BoPRtCIEV7l8Oh+7VnytUA
V5I3mApsArZMylRQ16x7lTPfwg7fnL4VcFSUQZT4Gb/yTfN8n2yEvrT8gSoz
dRr8AXQlcPJXk75pNElMY6IcjhtizCLMFW8LTGuXuH3qbmBGIW7fJlxNz9at
t0l9t5xXAZ9WOnRD5EgXeHndwlRGcPTtMtchwf8WOX39oDa4bZ6Kb7XVs2mw
3ApfNfpVtO2Cfh9ddCzv0m8x8E4I2kk3adbJ0YlJKvVjFyr+J93BLRn6XJwo
W6n2nckpE5Zo3zHdoxTtNxJpDm02gpi5qfCkCfPHN6gp61tsR0gBJHrRvttp
DTlV9gRcwTsuaXBliPLxTkck+k7CXyb2Djpd9ihrkgaxrLGNKzqvGJLiRHI9
TkjJR4s/sY3fIMGiG3eyAZOPMzfyv2ln4RJdOldP8AnV7PQShN82+m4NAsyF
w/itlez7ztwiOqcxrN1dD9EPODrdjd6WRw3TqmA6bNSq7xzc1xk5qS3xrX0+
nczC5N4f0pE/IlWJdejYRP6xXNvNMGqAtI3+XGS0sULajh7nI2bE66iXaT0U
5XGUUOI5hylHbEhbNDGl75/JFWsfNudGVBS3b7hRcfVqb86ak7W4X8/34dnc
3Ees05bdLKTSOOl/esZeFeQnhUn97mBnpOFt7eQ1i29G06m3d/PromZ+RUJc
PWdQ/fHSr3fh+G8nhYDf35eK8OmDKQyp8B3q6S6x6EhELq8qJS/RhaGIFEdC
SPX+eA+Je1TU2acjGxZBdkzr/8Iuegq247R17vI3O431nMhHkzjXWt8fy1IY
8UEpqrijJHvayIy0iAzsTPfdKmkAsxi7jlDhDdCQdGj71Kn60q0gTT78g6fy
Fpo34zChOgfplVBupLqBf7DAaom1GoNGvXPPs3ZLW1q2Ufbp0lJkfT62qZtw
u437EL4Qm8SEjhi7VVlp07CZ/YJcj7hvRnQ7v5dbmoDERWNpEiZxRq6G+HX8
AJ3BKWCOCvav/PxQ1+dOhMS9cCsNFCJlX1qkeGGMBSEHyPItdpcEuDqCiSb1
1yr5HUm+M5ekGDI49uPrGklWHu8MjbqT60QjFG6vqp8jIEN2GoxxKyGmC1j7
kQY9I1+5NSi6xL527Twv+oSJ02RQd161BKvFGCfZ4OfpfExsl3fIWO40Z8ow
kjtC80CXqGdR765PR7b/NdKXxlfnSSmh3Wv3uVmw05+Cs4z7MUJ22JehzKFw
MlRWTWsOzy7ZxTiVdO//r9aWcDs8qJ6q4xn7guQEcaDAM2qsrMzAEd8y6cfp
bOpx040qQf1USEZjhwR2//EqK8GDBdR/lB8WFo5NZoM4OFvsc4sdOqMFS7KI
dHQHUQqETxEVOO5R02K/0r5gU9F+2C6O1BqOc0ttP4VNTF0MN9QvgGJGaBxk
SacRNKycXbkNoQ7HnYwGZNZ57Vdlo4JXySI8/YejqSzD7ky9UdPHi2TT1+FT
EJsma+EolRufwvMkqI9Zya1RdLlqNJnPA2rzJmmKyA4zoFaltllupb/Xbx5e
R5ktc+IiHHWKJTeF8gGTQz01WCWI98ZstaY7C5oMxlaKOwK0uEFlfsd9NgdU
PMzZGEIGTUMV4WCwVKgLw5+AruIZrMuunjcnPvUupg6qh92viCzbRrnmenqS
aLsSMdCT0Mb2zW83leX0gxDdN3Z9mDJtKPayBM5SFPej+D2rtou2nmDnxl6F
OcIXJaR5KJE21c+Jwh2EsqADmYQlsankWMreVT2OI5/Nphg6KogHD6+7WmzA
R+m1q2ZoZDJPO5NJP1eNGE4eLTRMIvnKlIHMG+IizSEw5f8bDtVisaoVirh6
lPjTJJjNWBjQPL3bpbHotNEZpP6UGRijTk/4qFFIEtlcs0AIYT7upO0z+MpT
fi0M07GAaZugo/BzWSdlEDeDmv6GXiTNJxPKkk+2de92Ijl4YEbAswO1XoDO
IwB4OpcfRuXZymTswKcHAYCeZG1hIeThyHcAKWL16OfK0fPsY2OFvM4dsgWj
G4SmvMfkXLOYLCWjFCQ99Gz0PfycFojFJceVdtULgDpf3HW2fRJ+Rgl2cGU/
IuExaKjZwVb88o4U5WmJ9s2bUKw0ysyfFKiT7VCkNBa36tGoHQl89qzYz1RT
d5nuSBkJ1hhFnDax3nNIqw1Xnb49HsGGVkWp0RKvrijtS0LJF/SzptqX7SGb
cuiooCb3BwAOEP1wLGr8D9jG/KOilVtW39zjiE56Wr5eSpa6Um0Mu7cRwV4i
Ot/ZZ8NrlBA5/bduCguQrGYAl+lU4KKxVSDTd95kPxnN8NDz7eduqv9T8OCu
TPaw+QgzH2YxFjQSuGFV+BQWz+D43OYTF2hMq+5RDoKeAypifJyxb01PxvuW
xujK6MJ4dRAYezoBYeSsgJUPLnOHl9NbXv4IAqJS5ivI1FCO7oFiIEJZscJP
gYHdh1m+idkn50MXsVTnLj3pE62FIpirj+inMZeE+1KwAUxclxEBNrZ78bfr
Kal+H2ianvxz80iEYR5fV9vx7/K4tXja3N6ZGw2ebZklI6cjYMsQ9gUQdVIy
wpPPqbAXdrZ40yjRX6cucsaXxB07g+rBdhazWlZldSJ1v0Hir4y1phdMw4Z7
v/LVT0F5qAAjTBvMTLKOeIpEHVmEVWqtNeM3o2St9SR4RCd9TyBYP10oGtU2
B+Oau2eOG3Rt5JKjctShLRjI3w/cVOYUYg3yiNfyeApzyqs7a+PkfOeKPpEk
yOtis0HXwzS6BnxyXYQT6gp+D7W6efUqDD0nfw/iadUGQYG0zIQUxgKzBn9I
Y/64bs9EYLDxIWYhobOt3pbxoGUeS/06HImuxr8pg0EybSmGhCjYQx5Y4FuU
OeFONrWaZYVYgEG+5Kd93snGc3E4E2LzZlb2nYPOucRyVtEUg5pICrgnSbwB
zFbxU7/XO/Che807urzDWSwJouniBJZNATxn97wFM/B8KWfkhBGA+1jZBLv0
AjuBeMm+fqLhO1yk0/9bxBQgTwfO/JLsI82ekmphvSMus12V5B3zjarxvd9K
2jV0NGeJD5qGTfh5HBYEjHsippD560uH1S5vcAnveoUKPYDwG3CjmoPAt96A
yebRXFwacQjGXNw6PedDgST06MGIaYVVEjR7Tb/dOkFjmejjuX6zg/i8GQ8s
RjDuy/lsbl31vGlRy8xSWLHhkSl/YUzFo2zF/VtccdXltRrT01f7MBEP0gFl
+nJ+9NDiy5USIXgXtFgV31KT0LryyIorNOlGrJFbgePjCOB8MR560fpkn0rT
3o6adQa/7HuQcaNR7BG2ULrRpX80qpcvcKerAqajf9XhlKVXaz704KEXK0pG
0jJcfPhb4efwtqywH+WSnaTD2oZ8aC2+NFtuXaRDaESgTYY4AOIfqSWBDOzu
pcYVy1q3+JjPs9jTNb9eGIZ5BrgOLfSgaSnC4aNA8gXHqON5BBUsdrx8u/R7
Zxo/IBZftGJW7MOB2j42aBlRaCwfNCjDoVd1vSdWPma76H4uE51j2q7N9QTM
LKdlLx6NkLqey/fU5Q2hg4kni9/8GnrE9dc6892pg7az0tuE/76SamYfaqK4
WajdHkWuEW7EfgJbXaygPLtxdpkpp3f3vVG3tH8WQRZPn59WK0EkVJMTM1Mf
RNHvKx2TyfHmKQsH7N69wE0DjD2S3kLNyNQaCr/s+t3V6PXA1YlDiZFgr4o0
B5LR2rXNhNGdartG+w+OY3o/3/qoRhyjB0rK9C438ShiX0OvSLnWCk/2uN1E
tX29vsJkNtnTNaErrfVhoHLDlgYUneAauD/nXlRdlpDlhciFO8a5y09RiQhp
Q0Lw0iWh7OKs0ifeFako6mmdz84G7gbCknjnL2NO7PhOIeKKrDHL/O7GNrfC
3N+AU57uMBt8rHhMqXkCV8p2XKdnaiFIPY4zY9c8jSq29szbkJA1hR77GnQw
UhxQ8pQ8SZOzgIQI2HPotX4b/dapSzDsSsdggo6xjSAPZxYfZ9JPFe0Ur7AQ
k5njT6cPZecLdfDy0M0NCskvfzo8QspfOUBUoN1zONHtRg36p9/ACuYR73H+
tqHCq4SN2UF0vpUJsrdwRn6XLHF3FvkGTmZ75jpE+N8JDb+b9YghsPrBI7xu
xIVRhty7gJm+6N3+65KQz4njHjcw+c+119vBS7R2MBkG9+sn/jo/C7OvQIvm
8Kmp6SVF1IQ0SDDWnvKhv+gTOSmyTI5zpqEq0moTxsJ2W3PSqYeLz3XVtH5f
xxAcoG1gquG5McdgIbXRynV+M6wywav5fxKVspqvnnJaCu5OSkv3QgVqHxTi
AWtpKYjgkIP+oZjDzwn5hTelMgUYzCVu4yLZkTz0XX3p68fbipUtfGR+cRO6
/DGak++simXPwCeCt2J9A80lrfGgvpTaJBECjMIb/jvbGrhvjk66OF8sj9BZ
r6PCo3KrLoP8OeClurrBcYDdBq6uKmk67LsN4f0gJ5X0S7uiToYSZQPixUQr
Dk42VYtppGtPrRwIehyKyNvtTb8zyW4kILzAHAxHODWqjf0ftPWHkPAyQv/X
KNTybK8cW38NyWmH8/0paG/3ZXMSz4ca/ZSXQmmn3812oKzgkhORwrlwARJ3
QmyH04XVP4v1OiBo8eztUERRyAD8nlNTBU7T+SV5jlbUTgsWTm3fumWGutC0
wQbkWFfQnAmRCFoSgEO7GqPhVRIc4fHf/YlJqpBs5uPcHwabYSgKpUbydx9R
Aw6uB9r13q1iy+YBQrjwDeHIeoglypXI5paY7id4Wa0e9knMkk+hyQMRmSSJ
nnKugUTSbUrF/ENvMw9yR0PqH3AACEPPoGjnZ0IipKt9q3T216UYQsEGekPl
J99EHP9zeuM5NfLPgcQJu21E9BCcasnjA8Q9ARPCYQOhXM568cXN9AElrCT/
W5L8Srv0wSCmeo3B1AH5URmjINgHJQRuiFTmTdeMJyRlTGrKdIJZvbuDP8TO
+kq0VUtWlIcAZVSAEUOnKHsCuUrgocxYX/NiatQ0ap66Bcq/xKni5p8R6R+E
Ht5TwaRrjkVWQd8hwo6iTpi1M5NMQva1CroWQwqPIMKs+kU+FRsjVpurYROp
F024mJIOvL8ZXP9bcNeJbZiAxtfCnO5Ll4gDM603Bk4PyUH1JBfehyl86BTZ
VczFeXKSk80cOc5EPAdd5KaczGsyfK4GNIUcfcgcXo6qT3FWC51hEyAJGLeL
4SP6w+diK/XNDid1lxyJnEljIP4Is9a+oTSIvoCsnvzjm7P6xwu+Dk5xyJCn
v8B+9po6lKu+2mnluGnAcK63EUVc6SSev1sJssgoEPslNIDY7J8iUm76FpPG
givfloEfhsEbaBiqjW86T6fNOAe0Jf8y21jsyR0IScIdd24+cM1qJcnM8KUV
PouSwWrIum5/arYFvJP4EG0ccnseZ6lr2jtZ6X/0Ra7f8qq2lh7BzMGgIYy1
O1iTp9mDohsTUWgTswkmAnhdk5dZdS0cFdQQSb2Q7bB2mjAFyFNYMgqJxOqw
P1zk9qGeynXM/ILPMMlonflI8KhoXMni9YoXlUpInV2czI0cXC287tnqVkAc
J28Mi+zeacLuYEmk26r+hiKq9ENk8uMVO6RbagjK2NRBmULN6O1vP+1Hu0OY
gCn7xAViMSey86I/b8yhSfpEqVG9EneVK329Nrqa9TN/TrZafOJ/UQkJZKYO
RRM/o9KKqzrxKd7sxCwEiajWMLwYgaSimdGMK0GlXcuHhStuSlxGMpOQg6cV
tH5JcvL/KkXSXS6BiOWFLNn5cakXpOnRbTuKsqWt6X7GJTn85c8QKwLTo/+T
JrbdqM4Vg1d22ri/PjWnyRvi+i/pIPWds/MYohij2AbwEo7E6wzSfRlQ3svu
X9QOdkn9ivwJdMnwFdOE3xM5Hi/61R5xir+VGcXnaR08oZ+3VvgVi1EtCAiU
t1WAoT5GqeQTj/fxsRcpZDBNWgwzR+FHdvn4fG38s9NlEEHSCLSEkvNYPzCT
kMe5rLA8xI9AsvyzVAfhq5UZXt0BXRiaK92yoCWwf2bacvqYGdiVD+meKCkK
8sxFOQaCxHXkqkMlVyKuKWtpXuObkVt5XHC2oFpJa3ZJ3lMEMqN2I12eb+fx
mHhKhKj5zSF5/YI6U82B4Ux685MpUGhwAl1ppsWbDcPrGWYsFCfJK/rAHYno
t2gda33fuQs8+tJAEsp+WTWA8XVIxlZV1rkJmDPA4pnAkNZpiQd31h0kYIUc
Nei/nzzDyb4yYljP7cSYOUcdbtO64IIsBWerXV7K7FilqmFI9lP3Tm44R3nr
sI4ss7VuXr+R/RqQIVDPqzJsc+q4tPJQkCDBMsN2gxPQg4fBWMselo+xbk/A
uEJCpr734bAnV3Bx/ST7DXLBksz0+mHQyD+//ZS7KC96FuzdCWdnSsJqaHgg
SZElomFaVrE0VKU5Qnu6ujIGkJeMDNM+bhwFwyUvdWyhhUbI1qO8F367OC+z
xHvXM2AhFQGu5ctpR/RW2jRjeZxanQxwWKVg7Y4EyYDnlJSp0UH33wABG+G7
qbn/VFMMrgAsMz0Uanq5rXJ37JbybVby16ddxm09Uc5NIEJ8cTAumlsGm+m2
/hfiKP7Pk5eAt0JdlXfEtQbXsx5ICt5X/3dMh0NwydT6IEAWgpVfOhO0pl5x
saYqIwdBg3ScEw+8iRpxBBOpFO9GkhDK3FG2kKlgLXLFmun7QOCR4sYoFt2F
dqzX5TXDyKhJab8cNXPo40rYJSqK89SNOmjY/7dDYtuL1gNz+mfw7UBNAJlo
9lPcmQEYfc8fpwqhkMcjChmv5W15W+rzxvVdn75sG5iu3gDHEpr4luhWLwVF
I+aiJFTaUQh2c7vHg7D8pTvDv8eszRN3g43mMpni76dV5OFnrSB+xDEu7dBG
9zynsgg6Im6V0cDJ3po26yX9mDOzQ2L9OwA8Ncon2z09q77NGfaIFw3uxgMS
BxmLbAsrz/3A8gDxdstwMOoWEH0r44XL3HCqbX5QdZSYIbFonwmnXUCNG20b
KlAm5CRNrWtS9mtCg+Eso30KEdT4orpi2Hl6SjYQhDTuGv6kFTGHBC65Be7d
Fsd3gqIAzu3Bf8CrP+GYjNROx/6Bk4MJ0k2QVIHp7x+tdEJXuvISPDLApCUw
JeGxQOcGtrWLTU7qAUr/ayhDI8NyGR4sIJjGbFS5N8FtH14MXylDGofMOW+h
meUiB0/98Z6H4DNujCu0h3C4AiJ9y6Lcdn4IOTPUgRb6I7cuuY9MgdFb4/XA
xPE3ETcgj13awKoGt6IfD/09cc4hZPEBWA/GvwxXdjRFvWBNnz9TvQGLYfVf
Q3KZSS/vhJK2DNTqSbI4e3ESowcY1aoG9ENmHj1ffld7v1SJRmMm0qcE0xr6
T+LausINW2qt7Gz5GhkneZtHTMUyDSJH0gCq6sLoaQBzor9MEqWOLQo8hBtn
DCaXEUmQhF21xqpNudtuGJmUNTBUpX3HW0DKIl+ZUMEgxVLciaqYJOrLxNNY
uQm8oUMp2VaRMFCitoMOOximEcLqAgvLh2Vr5IOLc6etRvHyTS7qjOyG5DnN
DMalWk4TETjmqxQke+gjEt7s4InU5OQ/OgjCGc1hIXBF4tZY65eVZuf3NW4J
7Sq4DW//vNfe+SQGSqrsNIw/rLzQZM8pheiB+ooh0DEJzSUW99j8asdryzAQ
7gea5aFh1c3nFTajxxucqZR7DBaoDmAmArUbbSzHFlVswwcrK2aAuMeINWmz
EMZPq1dWYudm6FHWW0F+VxdQMyE7exrLXoWKqnx6hiQVZamWdRqpzg04THdU
Ke/nu5myoEFh7omExq73D4CHmQ0xOZ5lGyLpFb6Gwq6A2zZXhmKKgyjesJPi
c96IpSw7WohfeZJfeIlGRn+zwP6NN6GemLjde9+YUWkaPdasbxFy3EtFcimp
tam/caDjuj0J4CIsF6Bm7d0cvbJXqzpqTE/7BXbuE2Id2KdXkFjYhBdXvedL
g9Soa8PrZhl+n4sMLxwpANYPxNob3rPgGU+RsnmrWy+WyNflmSe1F3OCdYnO
JOrjy+dogVara2T3Co6jYIBGFAgAYgYXVg28zZmBcDwYSg2tEVndNkiXqLJP
GqGIBaDUH8vavmvaxKgLyuZQeAzfeOzabvpakICO5sFBc4pOtp8uS+nP/80f
Ma4C0BByudaki2ujs2TTzCA9fvFoEBKDMm8Y/8FKzZH3pd3Iyazq13gzjBYS
RWkCplm4LazvBM4Ei+JARgEFy8A9M0AJjjdJOUr433iu8wsuyDFdTfCXSy8K
9rKIHAX5DoenNEtp+iu6Ts/U7KyBfAOElOQR1aTmOKEmvAfliFKn6aZ7vb+F
6nhB9MyFPi5gwH4b11wp6n/PwB6PtMBlCY5FcHmcWIvjrCNPPuV4E3ogPdd8
eIF8VN3zcwudFSfgWXLOiAFMUyRTINYJrxuuBouCOvch2cMYgFzInxQz6yYi
WfBwcPHoTyNl0lwTpNXyPmLBJcrqPGJuOxpBKhQ69Tk6zMlPiXdWw1kC3Uqj
hmKTC2dPod8lyfxqDsWMkLTtxIaNKu8CKeOfnre/rRQUOhTYUyVhjkur/lJX
0ZgtqNmzhybjTeTTCrNVbrDGvyeD5bcltMBLvhmiKM3pqGqljzXD3ycE9BvL
yS7VDXVb3O58jjxAqZ5oZ7M4kisRMZxU+Mm4sLWX+3/8LKC1+ku0Hys10e4H
KVzp6hOW8qSEOVt4x14fDyhqhn09teCkdxyi6H5qIq8girnwJW4XdT93Ty42
Vupw4vRNmkSFGZEPTFpqhTs7DWtenJ0gw5KtSbqgzFZRje6XNGGGoe/AXFWI
kb7jG0ppxvcHKFofsjHhpIpcoG8uV5ZfI6LQu1cv23ya5EnftyhO0G6+E/q9
fixGwpS1wuw76MI77gnqT8xcJIG9HRNxGAugQQnxH+72YH5i21Dg4T9mD5VR
l2MtEU/vRlWQmaCPa3cAW+PP1vRnZVt9uiC6SRGsulus7+Fihv1d2t14Ju7e
jL7wfRgfep+D83ykVYkG3pFxfgZTIjbjvbr0gw2+TtEs0cXUMJwiBDGxYklx
51hwrA3vBXfHSamau5sh9xEssHJu/xTFEnRU633LikGatCxrFQGFTKzo4xxX
99IllWf63WxrfKJ9qPpD55yhVMjxPxJ+cq0t+1sEWGudtz1HwVnpf0ukhhv1
Di+N6xnnZ+kMF+DeNPXKmHo8t01/ngtk23RpICM4SuuXDoc/N9QA0AwTvhec
ooQz+82OL1WYfg2leQ24ZHSf0QkYy6L8/XNHSwK02TY9zheCUAdwtCnfIP/g
JZS0rCpZdlL397ALSugjChRJtTix44Me+1RhecInr34vMESKDAEm9ObvvVfL
+cSZZlOU78NGeaxQQHQ6y4WOMmUYIqB84N9dc9uyrq4HpjXNqHlUQi+xVnBm
2GuJFGWVh8Cq+EHlewcaF5eCDCS6VyXvpqn90dEhmF50CjTsFLeaECIOHjP7
poy7G+e9NBBwod6AwkbaQ1iNuw/EOhpCGrGxj6GJVPcLB61DKEh4uAYeUPqk
RsYvV0Q/lAxl21TaLz8hpOnaEgOmcY0JFgfAYk2TtRMsqrihFCRRx1SFfM5A
sxGkCKfqG+VkzY0gYZ5JKQq1DNJRLu/2dxn9HScPR/gP/lLzQ5Srr/KzYnAj
MbWAKIcQ3uerXiD3I8TgyhU9QvV38YZGXJqRn6nMXQH1Pq6kWbpNa9ZHNm6k
chaqF26JOEtIBegEmjKQnaybjJSamc3B3N2x6EeXUoiUizLJcHx6oFYdzbGQ
8D1MH9q2vPv6J+kYo2d5iOtzK07obPzsxnWcTUEDNRWpMPwD1NjNB1LPuEKr
reN1PXx7Fz9IjSfGHKvR/RtQUy/S1bAGsrhtIA9PqoEMpaNT1v05AxRKp16S
q0RKh4EtVzVo95yHJRePz4ayIwn5JTUoEVvEwhqtnKZjnGH0BA+oI4oM8lVF
t5gh+d6sTxs/lFESbCgGdxxChHJJkvDJDo5tZMMBMzgk+y+WnaIjVeiZRxVM
fu6xlhihAfupXoARmUMj5igxIKhmEYcV1Rz4RfDPBqP7Kf4POdkfIrYIdqlW
knpX4hub0jeT3D0veGVBI2EIHSdiGwJHExgUr1i+It3cEoFleRH4gkug6xwB
yBDjbIhaGhHMhtF7nnJYiwrS3bDd3+bAy+Sxnbt02+2230bKZwICnShHcrg9
U78zfIqXEgbESKvByHDYU3vTT0/nEUl3yc7TsgvttcP/I4JnRvFh61D+0Nzy
VRHuHU+85wGXYv59rGclmreTIs4ceJVmFGkDuAeqsUZVGlJe1Q8IJfHet5U3
ZeK1b6pQJZ055FivAGmnxHv25FccaM/0aq9EbTR7JWsfhukzcrGsmEf+9wQu
TorVRmr1AWNPJbWtH+O3giY+hxTvx0CuxnSGMNPNmPgRS0ITghaTvIRFTYdK
nrAxHGjEgbqhyLln7SKEGVEk1Nzx+eGIuSk64RlEqVBccDCwtai70omXRx93
WScSjQjTZ0J3eiqUVaxZ6h5ya15c5yuaVVAUY1pXShs9jkK8h5SkNDsgKDby
UWBKdo0Hg9Ykunb/Ztdxmq058wGQiZm94AEwuA9bt7nDfBifn/HfEkwviACC
RxyoyODIHAsjOp5M1CPQvzfkowehX53hN05t82LdZWT2JY972LG0oD3dJZJE
+Zqs/Mohvfx680rp6XUuHK8dzx5zyFkNYurHQtQ4hRRIfHIapT3FdfJ5crJy
r47x2pqE75CQ7nWwZkaTmaR4PcBzbPWOhvGKOTPoR5F4VlnLFjeHYGb2kr3k
VNv7x7d3IbKxACSlPhwcHjRF9yD/uG/W9ZNSIBDcy/kqiyFSotetUub08H6Q
asPb0O6Sk76oG+2ph7/9LnSI0kvw+2lGZLmjhZGKfuADmRA2CZMgN8N1Ys3R
dF3amNdJ15QE4e78fwaRhGflrsxeoeNoc8w7Ya6HAC00YJ/+QqnFcXJz5UrP
iu/pYzYBbFo3coIAh/PHi6t1A7pTmOyKLIPPYYTD8GRpJ1ApCs4gSTHSLmYP
Qx5GtkecyTXpyAtY71bIlDzXEXoCD8QNA7oIeRe2SMhS/L+jVuP6yVM9ojgI
mhrt3rtRHoMzWtyJFJWr9CsUcD4JtjwkPUT4kZlsVZ4UnOpDtBlzJCg1AzRn
/xUbKXHOGIG+9FjRSe7fOgwbBV55NBmHzdywoLdFmroLG25RjTmFCBeHdgAR
AMUxIx4btsuWnm/5HW2X4CaVObNGK+hNLE0w2lCDgZyC+FDnelu24RskYIAV
oo9rGSxds8x8n1l+FKle1t7Q3jWmTMf0iQYu8uZroIIk9WKkTHPVVK7XIP0i
BSgIZgkQmK/d8SwZqK3Ek2a2RWiJpWgyR7qPACEFrcaIkOtZwd/QPpzPncE5
ZmUmghqX/aoCo54mTgaw1TLrUZrF8SC7ukOXJvAlTaHvBNLPZW6C7XEEBL2l
CzXCWu7VczuBWDob6qDUnl8BBihCFPUyiHPX/ffKuIUoF5iXfxzoMeQxkK6W
p/TCi+WvHz9fTppynzZPWD+6kGzoK5WxCMB+nMWbEaaAq+H/n18azZR1wkOG
RnyFXL4NK7Qa+TJK8jKOJ89a5CjtSTlFKfrdmCjgCt4v15RTVAPB7THbdjVB
OeFjmI8cDP1Vg6aCL3oX3o1m5fJNDUs7N3wDHdpHFo6A+dA1madSmTS1LWzE
xyd1hfmynRShRl6sz9r9ZNsqafOmsAGUYGTY0oscKzx2mjHaA7w1FQoxBwGb
3tLMP0R0RThHIA0LWlJ7tpO4Dcf+RDCDhQMp2rEGGszHNGNMb+eqL3aY2ClS
oCyM72Gvpkwl1ARVoI+qtBoVBx6lhWWTLduh6r1XOdbYK8TjOhZbO2aZlCzw
Nb1jez+gPQ6mb0sSMpy1rh0SZm+9nzxgDG7+lVc6UOEb85NjeFf5WHQT768d
XpVSq3LwrJYZO6JnWFbibFkh79R7hvcZ8GU1y5RCzNDZRhmk1Fe2ENra5Tev
MpSkGieM7VOOrlmr4+AnpsfiY0cxd0Lev1chIX64Dd10UELuahHYI8iCBjv0
PDXBUf2T/BMLbMtaz4BRiqTR4gUbgilV4E05EZjczck8m0h6RNO/bgM6yMNx
v6/vnZs6QqBrt4+tIlS59g5J/+dq4PwBJREC357I7BPwRu+TyDEzg4LuPYN/
1IinMycVSWfbErOqZv3wHIdH9SxyuTypuJovY5saO8f9bgWAKLr9nAUa+ttX
r3qwN3Y6W5aciCfxy/oCBsXnSsCGOC7rn8qyfa/Yv2ZwbCOLOUfrCcPrNYki
XfEm7YJeTkR+P0ecaF1biQMsnFPHUb/p2QvuUJpKrw2R90m6umeeK57GKIBF
hJUGlgdWC3HRT7H1cmAGXbFvMv315K97Cg3PUlOxgKLoYX880WgThH+FSChD
Nr0dyUglIWq8UfjJ2eb8D5BoFNfwpf5zJvWVZZ1XHr6NVoZE9HkG4Y9fHR9H
1d1CaeaKHwAvMSqgWmF764Wa8a895HkbUkLLOb/yehG7+65dbHzSB1tNFvCe
NmTUfETVMUtjBH3jTDMiiT/FVcrgC5J6yUj98D5evtnANkJHVQYUQjl3xbT0
H/Qv0PpSLcNh2hYbY9TpIlbIMNpppLhXzK9n1g39R0jAwr6BEKyGMS2JgQUq
tow6XTmb27FT3DeEdm4Uo0T4ptSl+ms7aUQRMwfCt2TmRQaKgvlVyHShEwCu
FDzXY8/lCTYGnGoiE2oGEseYfQbzSN3iaoviL/R/ug7uGvdvMFbzmK4KA3pd
BpHmV8j0vRBPDcoV5/Phmgod3wgJJcANfgwwbJp2ICDvFEbDIBnnCQsyWJ5Y
vuCw7dZwca/7GRcT1aaDZDZ9VvEp7qFmEH89tqFrzAGQzyEUyOc04LhE+dfw
to8mVtzq/iyZnYYkyFlxqk9MCFNHW8j4jqN3PaBkJ4YOnTJP/dkwlBl4LKsd
MSTECUr6qBmmHXTtsgO+4rNv1/wIv5W4xX54vxv8CdR0O+JBQlZSA2ZNMQet
WuNUUuPeSvT2ks29WHAWMeGi600G6ByZ0scEVWqsJV/h9phHgQXPNDZOnPiW
FHNkq10fnTk/1ccu+wR5KQY86x6Z1NJAwCOlgsIN3BqSaRAETmeHC4h96NtX
o0PprYTH7mPRrgfviy1u3ljFUrJQfJPDdLXb6L+fq+QcZzT05ExwvWQqtX/V
8TCrLgUaeEoAs8nepH220oparWTpmQRN716OQx0FqvDCaf9r5ZNJzKLjfv9C
tsYgtYgmcf79admoF1UBehOELU7AqySe0TSAc9yqRfxkq/bFqfWdJkVORPVQ
rAgEsJWkk6CHQvBpwVONR997NJZF/wkZo/cU4qMIKy66sRYZ9GAB5EYoa8EW
5e+sCCl+lhOl1m2ObhiyWUC3RrMC6WZ1OSGRUZorrNTJMzer8KfwL9ccJbXW
8qJ5+GLrqsjbaJehPb3R27ruASkWetCAVkBPXYBS0dg3tm7SDzk1feD1hnY/
Qiw58RlVuDShppmzNwHQep1fvnLpBM3C7QsPzBjfzksxhe87BK2mG9k4LCVT
14ZfDxgVaLYjywSezDUHVVq5pC7/jUMm1XJ1nLlgivbnIuWp5fXPW87+taWk
BMoaVF6p/di2ClZ9mRGhbHX9/n/ZdfdL/ugB9WMw4jfoLtXvQ+VWSyGooVZh
TzCMdpLoT8MM+XmD3kvL4iLkx9Ms18B0a+QAaPi2+1WpXvgvSHZeBFh36Hw9
8lWOZWBew+mQI8APEBGL3Wfcr03xOClx/Q40fbjYBxEriMa+6Q8FUXvmw6GO
BlnYMIuhzSY+I2vQaJLAKRK++jurddMCpHgUxMZvWi4Xh9U/GA7twcdOkQA2
Xl4VpFKTONnpCEvKJE4XdtkqxwBmU/Llpeo0BdnUQJKtBa8ks7kDQWsZk5Bc
ScLtSxEU3yfM4D0szxZD3k41ySHoiwKTKXc9OgaZGrGNLcfeoykmIU34rS2y
7nkBucZMseuKVDJNbinlBGGi3Hfz1WKr6AOYYnszCILNgpOg+k4nrnulWrh5
xF7BJR4/lObMka1XVpJ77VxwOPuq7mdyfqfw8sDi2DANMg5Jootu3SGjdySt
ZYO01Uj2AR2we4kq7lkK8OLKrbkaa5sNyMyvLdSCE8sNwq5vX/cN/WTKpdbf
TkWEKwqsQBYgB42YdMmFgFbvVMOAYhTypmlvR11c0iXAWEd+W5BgTN9F87Cj
mRsdIV7fBQDzILtRkLfTV0KUaH5h5xOL2RfdJLZdEtKlD22CnXKbG8fZdlM6
HoPua2qC8GOqL6mwN/M5CIQC7G1qFrWWGJ9OzXMpJy6E241QhAzZyQRIzw3Z
Fm29Q0QJM+9fEiwj0hqWQuLXhabUvSZpxzX0Tj33S4yFx9Ap+cEzp6gqIbRY
+5C65g/o2keM8uhmdTwerA48FIqM68V2CtTZPgf+rXWooAyzDVqVgURfn2jT
am+e+unT5YcQoNc0a2Khdj1P7M36ddp7GA56gfSxWSuVwOZinpbjDBYND++1
Zr7cP2jGbU/beD0kIdH32My3lpqpbnm7EbJMuKIk5i8xxkkTVpeEnUKJ4/Of
ip6fRv9QmsV/Fwf0cFrxGk7WIJXAp/7lD+V1yEw4Rwru+lPRzbyvG7aDcW4q
KMK3jgE1b/TIvWKHqkKy0yb2S+Lc/u0JGy59Wc8EcP0AbhCp0gagWrTSN8va
Cw3YySWC5tuYmj8NsQk7Kw3qbtXa7vAAefqiFvaSa6uMc2ddZnR2OsClu+YH
TciJxHHTLn/OH/P4APtjD+csBmxN8ppoFz9ErLm+V2MRQzIdNYIozLD7gFVn
XS2oIJ4LTRWq/LZjiTkiNvh5W/URhKegxaIP3OqNtyaTPBAk0J3N/tC1AqOi
wPsMr6jl4cgC7xuNzPrugveQC6ImGdo8m7NDIxaAWsPv5rvcvg3NljJHFDr6
fyUsgcYh41pvI5mEM4m69tXFGs+6lCHWO8rtnOgKNiGINIHRwvyxesUy4yf+
PVUcA26Xas03c1UFBIOtsllklhSX6kfL4mIsHDdVXFeBv15YAsZ+yr6d8uoG
vroCSoqmjt8ujUmUdKRrBSihQ4bSm5SXH9GVz2UQ0ykrhHuoPDYabokiR+9Y
92IFwRhLmWBWNI6NA0r00P2T7RnwnwFiuEU89e3RFloIK6xPGQcWWlcstgLa
10GigAMyP6oRKFL7L5YKtGQgpZQRn5Yuv9eO0+83AMkKptXEAm34xmE9MAMG
hTZQD/Y5Wjx3KZqbV3jEzuc0kuj6F6cRoTKY9r/D3Dl7vH3AFN5jOkprbWEP
/RZrfd+1HxcfN3Bazt5yWtyIOnqk7sYru2tOzr3u+jxPECDMFA03nh9Tmqiw
tAxeBBpC7HG3YSOBe1FYDlCWSblTvjXQxM7zAeLfZbTiNL56Y6sPeF5O4jBT
MIwl3eXw3WVmrd54F9VUk6qkOPrzQfB13UKIqH9qjCyHl2EtKs1W9JxD18yS
HhiX3ksRHEk6TmmrnjyL33yUBzcw0EHpXc3a4bJnWgYZnvIm5RzOYwPTw//a
IoZ9zaTbhoeyQjCQXGcyfbKmyj3iLt13DAJR4KRbhStXIwoU7b+WH7JPvUVy
q3Rk5LPzEApWZyiP8pFQqMuzqEMTtvsoomLk1uJM3Zhu2SgDNSkPlY7xtdCV
iwewwQ5Lng3eWYGaunvBMq968+x3uf7IQ5t+C31FFI88wuW9k/aCHGMH5ETP
EZi7egyGZ4mnPXcqgv0BtRylt7ZeANtFsSmxzPruGj32L4Er8rz9udy/DFAM
lHllTNicnlPyuRtaI4J/gnnagx7yuZ/X+28GpdI6GSL1mhl4YnSoU+klVzYw
xAP9L5zvPVxqNvxxNsW+c+64sxPxq0SdTIpjzZX1oMXETnvFvn3k9cb4rRud
UPU/FOZXb8Q6SFAZ39deCV3FajCtit7NuEn9+NoDpZQ9MKzZ1lqvarxwZyUX
veJSVpAP/KU3cQlVM3kUH9yz+lYSQBKovmC3s6Us9MAvzBZJoxGwfHfcx7bT
jnPUvLi5yc4KeXGAt8PIB/G/Zp0B157gq4NY5tgt9x/+57BWz+hYdtFWN78d
N+kC8zSVvGWMwOz8TzxZVrfHtHNWnpgDhI3EkCZAJfm4uZrFsT/0qtl09tyq
4JfcImmW+eHaaHXaVd/2/kUg8BlEVrZvb9wSZx8EEVNJvi6C3+unJA4vLkdq
B4RQ+yd2EiwIFLKn+mr86zYiFDWY4C0HaTvsJ3/+J+drRzyBw+7WMJTZ1nWQ
tNovl9nQpju3aNKNk1iwMLLj49Pxs0gNnd68O8eTJ4I0L8GwGRivRTkf2p/L
G3oedfawWwzSWAtjHYVQSeH/5itaFGtf6oDYCuBTtvOUHyNmrzMTdAqHGnn1
uoIOg3Y1yOg0t2OavgaEukDK1UjEb4rEvgV+V/9A3nt80VhBKN79cCWQwd5d
LwjQAmvRfnN+MlH/PYlA7+30IRWxhxw5AvTJ6B91FlwyU5J//34Gg7Kh9d9P
iJ4UaWQoMms+xtpX21i/mfhPyq6nq8UQEBoTil6/F+mQKonoJRUNrUVi5LLl
w7OEZIAMyHVIva21qpjXfOvCmNoaPLixSDe2uhXkY6Ba3uVHagIwZno4c8xc
mAeUUB+OFFT48Hy398PaehU6Uk1d/hTFaI4bQb77QQqOFVLsApfVO1p35dLc
r7KLNiwTJu6oqqwfEC6cAiy0lOF9SNpRqs8vhZY/ItV/yPGDIfnPpouedAZ4
nLJ+GYI2RBoppjuvO6+UTxJikQAQkBUhLUsyyIE1LaQVuqBJzUBH6euxMMu9
G5uy2RaiUvYH+BaKaYDvw0J9W83bRPLa3s6kRraEZSBEt2n70RgtQ5mdM3+h
GIEbTZgr552D5mcI/FIh0ajvGI+B2X+E2n8DuxYcg8wYvv07VGpB2MgvO3b/
1vgfkRIjJ3t8PrrajuKBwl9V5HzwsL+t2yVMU3OlX9vzcK+rLRq3nLFmxlJZ
in8xm1r35aBt9xAfMwvb5Sv++KlvFid8ddDAzJojaPpClhN0MUUGY5PHEX5A
X+UwaVt26FxxRhkp4JHwNsAPrSIPdqWIYu7QAfBAvs2/gcwQT6RClx/HdbVC
zEKBuV5oby2++lOB2USjO9w76Vbaf9WULAiFR+agGrHnS8wIrCq6yh+PFfcu
M+BNiTzGFV7aZBpXexonT6y7NF5fCE3IRwdmLIkeQfBiLPYcTS8hsookiqLQ
Gfw4Is3V/idZ/tPX32MiaxD3STWck5uDAX8LkAVuUF5hb/uxVRB3NSXKW0be
2Cf2xIjMcQW0ghErnGX0iZoXMhORREAiDOf0bWTCMNifEqsqW5nvod+ErZQD
UxOE7fNIUcDx1QUQsu5j86CR/FzNr2/DVOO9tNLdBuznqlcGq+PK/GMIWQvs
8b34paGyz5YDl5Q2aqZ7/N7WDvKINPp0PYy1WCpIk/HNXqmJ5FiQ16MKuQB+
coCaXFbU22ip8nuFslcymzGL8SM1UnH/n+jF2756c94AM7SXx0LrOcRdLm7y
u4WZlPSD0fzZfMa8wSWJK90lgZYMoR5mHe0H/3FEE/xtY5uw14W7HSKIj+4N
+WPFjeqqvDTL1CfG34nK3FZuNSdwBo8CZ3GNi+PTQcXmjx6XuuttbdcZD0gl
MmQYNVNrRGko2z6cKnqpsfWdPPmSw1fFawU19WVFZeznzclBrJeKD3ErHlan
bT8TohPDGNuwEzXV/yePDMulVIIW3G6oLuzog3SIMHbxXPnqVzIv5CfZti8r
dHaqqvMjdEzec84duwLROPBaXEIk61PKcNEv99JBzFyc5TXP68e0PILrDj0d
kSQzrRDdlaP01rSUgZ7oT1JsvVTIDQwrqgjqMzMOMZa/fi2Htqm9bT7H4t+4
ZIsCf4qARSs3LnmbgjXgPJj/2Q17/JFdLsv8i9lg88ytJ48Dh78zDpz49Bcg
Wp8dxn0vDj6ZmPPlmhzRxO5TLHmU/wgYHI1aRt7WBPPkaaBE8pwYSCc9gsnt
FOQVRrEcDXMCcK71GPRsGYoln0d0oUTU6qCD8auyhZJwxGvOGE4fkGLw92nm
gJwhLkCaRlU53VTZS+EsS9JtjHj1BJxBKgtOoDN3a1Igd2M+RKr1gfiog0vS
yinr+es2kosyb2wuRJAcykGC9hraaZ2oAs0tKZsYhWeiZMrbVEgzueDXu8Im
aoW1r04oZCgYmCFE5lgTQnpKc/nr+w4E8C9Td2eNJ8SUSKyOd4sw8UWj2dUP
P+F2CCFYhpW+lCjjU2G/R8jiLhsDkAU49jpE8CR5+rQyOZx6NB71pz26cw68
f1MvCGdFB1691K5Clbzsw/1fsMKMWCwNqMjSRokSO8ivdPyZxGBzy6OJhBfc
k+B3CAEqQlovgQN7HyZG0EvTW7CvgBtoTKneWIs1guyy4QcDOw+HH3CFe+2D
j6mWVHQsFe7TcejmhhZ+YI4qMwcG4wRLDonnhGbCgro3LRKlXq2xJ/bB5ZSm
fVBdJItFVBJJXJspOuEow/sOLdk1VUw8DLNXEkOACAnCRDbS9TAEM8bKb5ge
UTSwyjx6qjMlD/3oWtSUAkjkwDySw4PYpjgWIDmPB3YftyEatbcFIvgZ9NAS
zVnFjbGM55CWAE03L2YHsSomtVxhMWhxk/HubYg5C66SyAIRPM1UnJIQrqF9
VN4qHTiBHkZvfOF5G3f6KajZTTT2aa0Fo9TWE3o/ZTJb+di1w6zxVklKxSRK
+5jZe6QCx79hu0OE0/tgsGkzmb9tjED+DLlFj07a7UmRNd6uFeP20ZYiqLMU
aQHb2jbmkmOH1D/s2TyjCPxZacuZ0qBUnAxXYSjvLWSPrGeWrR9agF94JXqS
MOE90PAacegsuyhCm8Lg0nZRp6n6INcJkOsP9TL/LmEy6giPowEJrJ4NsNrq
narhLYMH+3TG1WVT2hx3QULR7S5PncTRXsR1xYXQHsYWy/AmPpnRUzgj8D0U
k8nDoe7gRC+Lh518IGSraps7tgSFWHKcJCQtpQkchm7+tWIdfuY43PJ6zOvG
2+UPFqNbc/lIRizXFuNCxsi8nlAUIdK9fo3dEnLzfNBRJC1M8xXgcBtcAXx4
jf908bzvXRSQjSe/wPDtGB3MUJksQvGCkJi5Eg7rq1NMj6TZe0d1I7LXPBic
A+e9HNv0MIFiu1kJTTeoF5R+GsVal63P6kc4HsYvkSGCu47qIlFLTI0UFqJ7
vGDbDFfSoD6tyAksFNkcy6erdOR4Q4NURnt1XMgTdxJgIT245r5FkEH+/uiG
UPf4zOK1n3M87q6Psj+15kLgoroK2yDV5ZNsOE1yCVUEbsoBuL6di+lVpZOR
AutQTF5RVjvHXKefvCLWKB2b+okaCSA+ASFYeABGl/0jaJN99AONyQBcecV+
iR46ZmjnqCKCWm/rIzRGvjpm0D09LYWVa3jTnHWZf0wnOQBt5eEBeRpo/9iu
lqhvfF+KniFnVw6C7XqGucBQU11m67Pd2z7abeHlcl0gyE0abTza9RQFoW1n
tNzvPXkLqhW1YWVYuNxm54BX/k8SgZEVicdTjAY3r7h/B7mVEarYtgZCDjQT
i09Emjj0Cjg5Ye7hD/nkKjWYwFHC3avZCyz1rGFKBAKeQqO6UoOTsBA/ZUwJ
sDPTEFlm/h+Prm6bgQYrwwuU6Jzijy3Cx1RvvhdC+4G4v5B1GF5ip/b0oxND
k7dobdyYrcqxPBtHawjOki8kZMCiqLtNZDz29fGH+kTV3QBnVKQRXHyFPmp+
ZWfFRXpeP8v4DkdHgvYSJExqkSCojx2bG51zFdH6pxdMPnQF5wm1GLakdXSu
r5ONhU8UvVFMOzKYfR/J3OyvlTeaWRTTOBn5v7+E31Z4s3IoCCBrtMF0uuvp
WuSf4sIEjv+cb6+kTikOcL3TALZHWTtl/AfgMhkMY9P/5j3OG/RrZ197QJrh
PBNQ0S9qrWlUuwGD52ET9spx1TB+Jm7RubueDWKGSyoxAqw7TjAlpl6KfE6v
3Mg0V3+WjwH45qC/M+stEsYTSduNKI5n0LRZXQNh7t6PXhWbAqqvwqIz+iij
nwqeO2imgSyosXrkWWWisyfRjq2HiM9GEDpZbxddK8BlJWXVdUlNM+Hy7lKl
HLR6tPEoI2LwZiQoWCGwBv74bXMl/baHijuNegzrvNn/NFRiKiuKTQCCbC9A
W3/fYlHIR8c1SZdK0lX10hd1wYUckkScaEPkfp8NtNEFebgPAPUbKvNruz5J
7oy9Il1Fw3L8pX5bGL6mgSqAWlb937xs7Uv5SuinwjMIG4QOBrihw35/MtYq
n1sr6rrs8RXqhP4mmIrO9Zrs6sRLeZbhZnh91uJmG7RrCbdajtvPjQgXQzvt
jxVMt3P1aSgGYnnb1hpp4w9Ja1eD7tNBy8z+JeKVeDKsKH/ts6k3UouEzxey
2nvOf2RU2XS5j6DwjmbGRUuWzbgA+KSaesrYtdeM5ArVzh/Ei+Uw6LXiF0E4
mMVCOb4s0l82aV1fuCKVpeBDbPOn9ixV2h0voTi/ecTySjAdSa6x1GVZxFzm
1nBxp5wzMgYzZPaUtpfkRXeX46uXKmCVjjdp1nNYq81hr2Ol1mBV/WG7DaKV
Tw58ac/UJnycGhXwKbLcA2XbeK3cHEgyn31aUmOSnoad9eFeHlvzT3XVCyyP
G1n+lHAr/osatAzulVRcGLEMiMIs2WpQ/Pt+kpexqlgkl8gtEk16wNedErvc
rEOdm2XNz0LTU/u8XFF28NxGmzwptUommM81Wy32pPxUhonz54nUDyPs5JRx
O5QmuQrIjpzThr4kgyddQB+WefCIfYnqeFcg8C8gtQ+8PYrJ+m4H1/UyJ2pH
CngviRbvhdMdG8TXsWDNHhnCS2J2qsM0FaUNpzCaYwml9LP8ly8bHHlZAozt
rRC12NqqY48wJnm8DKAXAfapf61+n6VdaSp26Krl1P9r84vE+yfX0ehmhwSA
YEDJ/cRPW2i76ReU1TCe2qtr/J4JO4OiDcLPcg/shx/wUkaxByc45fKQpC3D
9h6VQb8EtTShYAbeWglLyr6FLqsurPxYVOM7uasiJEeJmTsZptCNrGv/mYFm
cL+BJCHn1jgIXyrw19Sau4SYSC2klUhb/WqucGRuPM2RSkgVZfy+i1IKPhAA
7WZVPVK2API/PhyXWcBkpRyLLp9f6TI5YtREmV/GQ1NK+SesDPz54g9xdCC+
Vgy9A/dAZmSk2sx7jOhIxvdYAC7xvGDRvG6Srpjkz6kxcBiUtPyqhdReOJo/
GX565ai/dckn0R4y3BJeV6FeDo8kkyCl9sWWeuM1tPZhoE0KO0gH+qMbcEzZ
RpfoHI5UvrLRhlksaefaWDlksrzF/LfpuyJw3D0BrrP79HBYHxbbKFgyGqMo
UAcuwO8PI0cLY5HNdJKEchLuoQdJld1V/fi/MVc4GNDXPync3zl2zeBKGvpR
nrxDY8gfWnlu/VuS+Pgsp+1udcTbdnOZ2o/kRKl/H3Q6/UgQb/3Vf9pLB4fA
C4wIovb4PuLVBd/piTFbpy9bJ/Nx7YBSNiHX0N/XjqVxc+roko6MOzSq6rdq
lSze+jrj8NTM4hqzXLOmjh/38I1NCAuf7uHS80GtyTC8j+qc3Bwl4qeSBASH
1uoU+FXo/JPCBPio5/vFra3Rw1pH5gU5sao9Y8cKD0G4vcloe6othmyKUyin
FMy3Sc/lUBxaFTuohfgk6wX15lv9Or9qLdsUFAFpXOuMYgS0aCV/rWvqio/7
9vHtx+l1zcjECqyoJE+rpWgh9KxqnGhEgvfqDH5NM/XmFuEvc86g5zCtB16Q
QeOJ0zptBGatfRrDWQ0tHAXOO9JnwTYHi9QUoNpvcubXz3Nv3FiDHi2sWSf6
s4ZaFym1y1vNHklqI2PZH0CFmupI8OLTMVy5vkjtysDvT7fRnfocURnKMi8J
sAVi2qHf+Xa3s/uTb5cCPVXW8h5m3yQZZRwbTpSEoX/rwnQcZg6+458PaoKD
l3XkxbpWv4LUoIeMNjEqOts/iezlrCS/qe5VAgb8UG04ApKtVOHu9VAiTK4b
CYhIj1sRNuU4Oo+c/0b73h5yp+Quve0q+3jdDlRhZcRcL+4uqWzy+aQ8IFba
A1rVkr0s6or/s+Z5peTGea6chTraEAXJsHSBsu6YHSxwdQP+2+3NfZspQvqD
JCBAGmuNqNN7QvwtQKS7cnEi4+uF31LqBLqCRB1EoG4G29v7ffHAg9kvdg6c
BzBcXEB4teJBB4QblkniMccNym4/42/XRJiimmhdsIX/fNkmTqtUzjAZ1ZvQ
QZrebbIXnOFNgkwNliRQZJQTGMaQY5dL2NDf0870n3CfKCTan0rJOd8f6vuu
saU0leCV0svkm0z42UO+liEi2NKzEWJzzDFO45wOVvdtEjRN8JaHKQtRivEw
rfvmdKbpc8drC9RxVPRcQTLOYZdSXzNsz7ga27vBCgzAuq1kpR1rcscUuiNF
172ly5JM64eH1nGy0Pu5VSiYhCxSRs2qGV9ftycazWgO/32CPoTJWgVVFd7y
CEjVXUqWASiFfV75VD0yPGmMtLVXV3OevPl9fLZjEGUeGAm/y2Xy80Onl1S7
mBbi1xp6YvMZBTqEb1AP78BCpT2/zP2LGUWiiCoL875sRtKSjHNPqRA3GZhm
8t8Ea4+E2fpatKCVkurQuJ3tmd8Q4uuuFlcTm6c0KjnSg3Ztd1l4yqrBKDUA
nvjBnjJOdkVNg89jZrl4Mz0+bRMonEIIODmBitJMuHPpRSTQMxrWlzWOht4X
IH1TXKNKF7gw30sicMtA4ICrqqckDG6n8cqm6YLDyghRtY45+g1WLTeeie8o
NHylseQM9VFIS8VnIMjJDYS+YNS4xj8YuTAOzvwpqpl1oqGo1WznpuFNkx3s
2o9GLVzHWhB1/5uEJy7B7uU0grxqCMLgk7Vs9UEySbF3PuoLPfMi9KEdSOG6
i1g75pEUmWDdh5ugxHwLyPNv/G1zFiGtOUK8lvHNip6fD4J+TVnw0ma5niV4
Z+5JaqGPq6RZXX5VzhmKjF+ujhrpjK5+p+qOvwK7hEN+N3gmR/sKtuW9Lk1z
PVIzaN6YlYYLTVSlwNIBGaa2YbIutbqLbkvaIOucCqNfSNTaVCAwZsIQwITO
hMNFRY4X2aazhFp8Qpb7SDRL9vn+79PoPMHsheOKp7khHPzakb7uzopULywp
iZPdEbZnqVMpHVPTI4F1ah7R5qwgF9zAGva7pYyoFoRH66h2CIkXmwa6y1pt
CJ2igS+zQ8J8oCeT9UUT83uuqQ3oCXvUF5i22u/J61DrAL4RhlUETAdwwJH1
kc3b085WECFv5g6+vSZr7aK3qggSGrUXx0Hh6d714g6y0RhL5cPTDIAd6uV7
rQf7Q41R/1RBhyhjQryGItcSZ0G1t3IB1mC7B6SOmSCp7P4z1qXJFUgN6AuH
VJn4YRc/OGH/HWF25NOAVLJ32/JBkERm6bzPUufjdu05Pv8SWTxfSeQbhvT7
DzppOTSg5ul9acVimyrtvJvyON3J4/lrZn/qR2Bda54A798WcoMy1dpq0GcK
w9zvssRlPsc+7ed+NNTBqg/uFHYNFckpZMn/CtYqiWj2Xo/O2sUVNfQ4O/nJ
94vt6VKOqfiUIei4dXyywKZakTh8YlOcAyTxgsZrSTdUIh4SnZVC2oCBotPo
nBpofo3I02bnsBknsCxTe1NQvRgoVFWjJeuS4lIQPl2r39TaM9PyIb3MD8iR
Hkz2QU+sOLPck/h4EJQj39t9QD/jV80h8Qhc5B+yFBfxGNs6C8/45SuDBXyi
u9ijCy2EeY7ZqWDI/XghJUEQXFYpoRmBAbWMlCKR005turKjjeyiPXWFWKRG
BmwQghPph8r7/qgKRQh4eZNEq/PEBwdTrbEL6UR0AevsY7yWKcqw1PJQWiEP
dRoQZq9AutdyBzH9ZzP78xuElaG9Rlg1UlZpRWwJaewlnd7y87/BlcSyzKcq
SsX0iWO7rrEEUP2E87gWWMbBCR+VWfsZkViwJlt4F8W0COR03c4Y1HbU26mN
pwWK/PxR7TQLs+aTas+ER2xkSeCl7IDaY6IvsNjGmWKC62+GHPKSBjI26sep
bgMehxTaUnqx3i3Zb2FtTmfpz5f9IT/XHbnPCDKKE2Zqjnvl40lznL/yy/UM
w60Tzw+x/FmLCJ6MaXX8nQygDyXPyMLAGbLXoyPUuLANYOo7gvZmvoFIlk/Z
1auL1W9nYqxubq6yaJ1+bevlFXSderiAeWJvre9vfMeNtvYgFPNgqPkTlQBb
odd4eZgIQaobzMVvkMIlmTWYFQibOijtLMyFy8rOvsQd7dETHZ1432IiGREk
CXvJbGjSkfcfgeromuhFDMy9KPsNJtMhWIWsx+H5bUB03NDck8e5Fl/wKwGk
FFK/81JWqfGeLgELZPTZ7Ipo1fiOJVX0RJrzkZHHI/DpeNCw/RbvU6qnI3uK
mBRAMvl6zriK+AZRINKoKx2yf9If0lviCW+DVUe4r9cYRj5l7rSNz1ZBfKQg
cZJl9jVSqkzow4AKVA28+WzoKSDNjd6N7zwG8CrbRPzhlj1KzmHOQc5T7rJ5
FTDWBxhTl4I7jGF6Xv62y+aC2A9Ufhsozg6exXj2xxMsRf9MR5tyxL/myS3H
hvtHkW4vaPDCBDVWfyMMaw1kG8XWuie+rDpw2l/0VzfOZn/ad8HHt30MeWF6
qWR//6qxeuvEuefPx8/xAVJEW6JzdrbafcgbnHEvmSbjdrtq/OTP2cTROV4y
ZVeYbHqNE7npgOeJotgXemTWAppk1X0tlyoEIfSMOAvBvZb107gZadXCiLXF
ADMfdEe9GaAiEZFmiH5DpW4puSIXwP1ir0fPGRA/FFbNN0haHnVzuIw5w91m
jQYVrbxYTzcPIvpX/uwWnGmCS/O8XeFRnYvzT1m9/0S3ilGLTZTpt88WZsAd
9Ypmub9oSE0Clsxi+B3s/u897H57FmrEZDj7fh6iN5cC3vyK5VjRqzMj0Csu
czrTAme+2RBqSMIzWCm6xkrGU0NBF2gXPnbI3m7wCDNQVboYV9/ZHaoZn5GS
yQkk3V4qDfa2H4OC6TBBvML7N8sZb8P/6V0z0Q+NC1mVyUrllzh03naXJgdd
0kVNr7cPaQy1B3QPYm8s5Q7oPNpi9DH+N6GN9+jNa2ncnf4rKTYougKa3zSq
SJw78X/Ny38Xkh9SdVW0CGNivVwp7aph84zxT31m6EsTUM2ZWZG73WdqrRCh
5n9lsEqFodnSh2BYquEy+jFulk1FA0eT/6xB5VEjVzUhFL3zhJLPSw6HrP4w
bG8vUhG6U38q/b9xNFG5lxnFVWCxTgEfEeLc9HFaTWZwOGqNWiXucBPmH1VX
LEKWHKE9DXT1Tya5IndCANMIWJCU0IEoowrsZvlaJYJIlp/oHnPcIET+NflM
GSQ81IqWawXZ0BfICfH1NZ7WwlXUtlvLh6HsiKt6KXSj0qJlSlyJnKC5VwE3
7IRYxzrvGJyRm94/JiQSIuFwJb3hsMVyfigOGySBStSyoaDhMbqrT/m14hX0
sUodk027fo5nAzvwNF2TEvKfLCRZRDHWR/hpPYwBxcHlAzQHg8jGxCiIAnSc
GRuTsJO2On001yYw1qYuuR8Rrm4JlULznrq/G8zf9uexM2fAGIbBZUqjExvd
X+JAnE7cY67ULeat7OjRUxdM0oNxIPvPqrn2l/x3LMGLV3kfZn2MQqQatjY9
LugvKfJT/GwzskFka8XNe+ScauUpvwaSkyMaaBMIrq/DVWdolHmUSc3T7HHj
YPOEFe3zMGumhVDmSbL2i1Ksm3VljodXK+AC4xgEUFSrtQz6OSSTzN4pHtx1
jeGdI7IHS/yNKnS5ZjQWaETTMvCbP4V9hzV6nO7PncxIyxroETZNq4ydTwlt
zvejmJFOBkNlQcjcfFEYuYT3Hp3ggUYuiycpDNxwFa8YtO6qrZsoo6IlX0Lk
lzd4oDTEffL/iNu++EOXgMWSFX8PSezuzlLvBDnuEhFtW9dG2dT2MwZ7Nvha
h23hs2et5+lpNRT+Vl6gZmE+sy64tiso6oJXGjRIHTtEATki6EDR1VVhWQza
sC4Yq0eXwaER3RAKcFzMD0MS2vW+jRyuqdmDLyjARaWSKSZYRDeUQLudW2kz
A2RgoRi+ET23fi5g3lTnZsTVows34EtoT7Zsg/FMRpPa5WTXJL6cSVRHAyXR
FvtYd9EKt39bYxdvElGr8qHoipiGO2ZtnV4IrxuV6lahJpJP3tHmmGEikGEM
tPE3yk/SBP+om1dLX7mny/U0DRGkjNhABV+lZBbHcCDKOpKxiClUIzPjT/1u
MtKJr+JVcZO4ahPnnLaESz8Hq4A4qVh2odeMFtjl48whKsE7l46r4aUph2Cm
xe1jrfRci7v71hfLeSh2B47qrxPtWmnKFyFxnYy9C3vGp2t4l76hkGee4MwQ
yy0gYQAFxp2+WW5ZZmpykRMcxVYe5+B1/eGtiCC2ADm7tVGjXiehjdWaoQ8M
cyPdjP4bbzONHewqMzCVfagyIqGProS5Os4fj8+u+hi9BDV87T1jyIZ0trV0
uf0v8pjPTsLUtLpT9SH8q9cZFLOElA1Wl3AbVhrTh+eSl3FtqIXKys98MDLi
wB1Ovuv9H9HgauLMRmqj+gdU5WMnsQ8J+uM1qSHvgsssVlAOy/EiLedascq7
+jdgg6OpRqfLgnQFHJTMfjoPEfKRbrJPvQ/JYx+CoGV9PwlmmTn9B8RvLJGS
eG2hp0vRFIWdPjxmBY9ulWmLIgUTL+BiqcmqRfV9jVMNYnxXjJGqGOZywu5G
qGwbcq6xn07de50PcMduyqQ9DX88LTAf0L97VWZi1Rf00XB+Cs4vy73zhCon
xXre/Vgh9C2xA+ZwbeV/8tWe4M3xYzH/mLUOeA/ii+ne+VRCT/HqkjYL2C02
CVVMbc7EsKiiCAn6ukTyuET0149vUx5wmxV998n7U8elEELuicwIyK9qNXql
jAskwV8y44ZVdaI1wSVoSr1PyQjhLDeO40DjAQ17V93JjqB95Pcxj067T9wR
eYK86kB1a9VbrvbHsFHL/gVZxJJg58oW/lwDUjcwKK3Zol+A4OG5a36vCFbc
t8oR08jQvd9WJwVRkVfPqgzzFcUBYYz1scYcnrqJuX14/H55ISr7Ii0LGxPh
ttm0CN9mU/9vc7LeyLNdoAhUGtXO8NJSKqq21ffF7Gbmo9fx02yEH8tG30Oi
575IxWxeqi/mYawPKbsnRhYahq7W67GVGgc+FlCRkFUNLCmngBF48tT6dK8V
vRarvTnQw9tkMT3Lf5/D6mml78Eqt1IklJyMKwmptmMdQxX7PRC8UqeBzRIE
nps15w1b1zs3stqPh67DAiLCX+kPffk573Rr8hJaG41OienpUFpLLpCE4udH
iDWEUoRyY0ySXEqTW0ekTQKAtH+UnsGafXQyOXc4KGNdauYWrDGOgSaXqC9q
T+O4vMKSf6ywFEpHppnaeZwJOPCiJGZq9O75Qxwcq8JLKr4vI6+WwdKlEMYt
+rKVRwpbpfFVT3y0WogofDQfXsJ5idAFQMf0vAnAL1494wwatR8JnOcQjvXx
AYqx339qT4YeWkyTR1j4FQAQm0bBPMws3xJI9RD1wyj8HLi0xnEHNZ+bj4Oy
ESURqZaaQ9nE/PvELMC9zhlhVWbEufwJ4+nw6P5vZO39WLZ0s2u6988JZtHQ
bClOGAr0b3wX7KY6ki/BAe/3uN+2JsAKHIkS1kaYHStYYTICBL6Ib/v+vh5y
eV5f2MvhMkm8UIl7oypSKx8X/n+8H7iGzKVxg0+4yj1iH6yYtJPymJpOzZKC
wWtpn9zCxf/E6veCeUSIQTWmE3WYTVtSkRrgHYRnQrf3xSJ2BKE6tY0Z2OP+
dew7smiXofMTTYbM4Q20rqbSd14mHH+UFOOqvd8tZ+KD0Pi5qqt3zQ18Stim
g0zHbjFyeuQyG/kFDh4+cQMgK1ffvJCoLzC7tuaq9H/1YE1/tZKFQ2t4twTx
uXKu5j8w7eUXtzdVnI/tvJwQHe52TbWBzY+BKMjArNLRO1H7EMtpgYvqbmiT
CY5NuNg+bTfKNCzJVCmbv12nc3A3ruQs33E544Bi3tB0uuY4gpFLY69sMZE2
DGTxWF7V5Yspjs43oSF7eED2p1H0rUlTjROF7ckeXvxI9TGpgHmIoXVLDDqb
zgC558MwjPS7F4yZoU9LnVXpm1B9b4G3PehK6DlgXhbgoj6prqHku3qz7r1z
B5qpa4q/W6fjNcr7B182xvEmKjpNwCVJDHPMaQpQ73O4aDrOHeORSq3aRtl7
lhU8RXejjTwwa2bxVCOttmEq83C6kFB/jqQtdmCj0s97o0kgcWdp+njGZ4Mn
gY3vlwvPwxVMv2lZQCI7owXvomVFwAYP4AH99Jip5a2MtmRqzaISvAF6bccw
3uqrcTTtUaeNFVhv/HU2Eh4j6yLH7Im2UrEsOVhrVw58vE8zz7mCqf4ovBDn
nypkk/TeA0i5BIXBYfH9XKD+9eM8/qH4hjW/pU60f7otqN0Yt3r2Yo0uOXUK
nLAo7YyTUQVEG13nenxXKV5ZS/SS6EiyYiwzO6EmVfiejzlJ45uNL1gmlJV8
P/fHrs3S2Bm+2/EFHTi/BmfntbO0/ZkfjlU8Cekp7y6b8Q8RiTUdlhoka9Hj
OP1KrP8QqNOZh0XhfHYmW0tKgAiW1ws9kz1JcEDTFFrWc8xisER5j5Os88gc
FB0l7ST9+oFqIT4Jrsq/KTaIQ7ooCMA/REkUqUs/McFI6s+bshpYY6XoVcbD
aNXb38MYbZFhLVVQQSLC/LNcNuRpFmOkwmVipOCF7bBIDifrtGSyheLkdKk0
1V3nklF5Cf/KmxeD4UoDNFA1DzU5SlewDxg98McCsVuiuxeYySZ1G/tJ7Qzy
lXrYJ44IluR+c6q49NLiqzZwjc51jXSKcjdMJM0BYfReO54xiQsLReyekjKO
WS6OQswr4aBxjbX3U2+QhbATv/wgyxc+51aRSJsXAvURoFkHF1Ek1kfDlsrs
wnOQEXm/lYsHq/h7U/lRA6OQiUetJpmnSylBFINDjvvgRIv9jyflo32VntWs
HVE3SUoupCxg91ZSkgH52nbGWifLCE2ueSUBJ9Yw5r8vmxG1BeHgtOMY7XZc
LNHhVehVTBrONS263BkfliK1ybATkW6LUkpS3d5hm3BhPs3JQmXFzvm9v5Bg
+zRtolODg+rabgH7Y1E3pejuUdjPE1JMJoQJlv4o4m6h2DIQaq2wYeWDhNcn
iBNOT+9vTd40XxY7jYJfizuagkaH9zJKnfC27G6j+/FTnz8sRiOnzB5B7RWX
wChlSfiu9CC1lMV74ol/sQqmnJGLp56/V0hPjisSj+KHNz/A3ChdxsGqJ4Mm
nE6DQWKGDSHBvZMghQNYPsfqN87Y3sIDZlG0lHFDTB2Szc493O57WAbYuXkF
3tUKV9bQEd1onliWIzr2+dQdfeEaJ72oA8vbj30V7HTI8fu5pKjztsiqY6Om
N0Bce3uFGe8fgiFiIsSwsEUfXWQJ0VKBz74ij1eJg/keZHxjUNj+Q10YcbVa
6ZZMFOFJTD1eSonidmWRywwlxz3jv2RnDXKAmRDwX9CWn/DjY3P80KBJRdHn
w2DSTV+VQ7ieteVsL1rPzh4h2cOEKOuAo3mZ5ZnwK5ukhtGy7Ug12ZrqNW83
Jardm8y4ArbBSlvogDMpyESKYXCg1b2PAO8yVEYeJ/fjAOZipUwXXcX4OABK
coyqqzrur4bnimqakbMFo5sHuMlaUhJaSmeRHyjEze1Njzg/Xycx/LHhROF0
diY342ayVPPuNe7rW1uCA0t+g0CEnXiApW4iANAUm6+nNKLxMdYou95DPSf1
jlHoK/cGSp0GrdUd2wK8C6LUNrKVSJz8QmFEt5p29rsfQ4fIPzA+V17nHyO4
VY2hYz4MwL20yNLJgaT71Cupn4MMKPS+hW02SlIg4trUYRHQnDDoX71A0us7
M6xgVo7mRk5kSakDt1YZ42lCj8k7PAQT2LKRx6tmtejB5FjIjm/WD+rg47ln
aUMxwgzM3AG4qRzzzF+guKdIHdEpJup5eKkShlYaiug0BNLjb/JT2YedIucH
sJbbeiDuK2vaGGkKQYXBMA+NWTmST+4ACsMk/39mCIenW/yPEyyptsP88TY8
Cqv4glgzIXMz+C3SkSDaPWSlVTC1b6JDGbI0kZ9AV2HDxjXMOLrAmU0mlcec
ZGN8TcdLSedHqdt58uXU0ZyCbtDE7CAIQ1nutJxjszu5wNVuR40MPc5w/CjP
p0DZtPmdxy1otYxHNqZT2IuXPWWbs8q1DIfkDOe5J0HrvAKYUUiR4S8rSClG
mjlCgSsq+yWxL/AUZQeXd34IY+wfxbt409fp3FROZ4hAPZnJ91AysHqyiRLb
ZI9d+JSPw9Bd4LphI5DcWxm0FqVFW2B1iBsYrfoW2y0lvvlC1cqZkAqMzT88
/B01Vuw1KiaNu76B7DOriLCCXS5XolSJVGa3Zkkh54BlLCcwrFRrEbvEYReG
tnzon5fWWunPF3ewXS9m37WmO39BYqoU2LbtNzFtScvOFWSaot5A4e5pACEq
wntfziutZqyMQgd9RYNpky3tUgzNxwBP9zlx2VbiavT+cLl9TI9cYa/W7MQg
i+4OH5alopbWnArZr8c7tXr3Lbti2JNI9Vv6lIee+RUq1maEupeufilhZTpd
FiPFWgv0o3ncvD1qS7L/pcW8mVKgiQFrPXU0NFIXIoMDM5GuntEG++ZEVqRt
NvdWahKYDBEh0bGNchH8KUSCKjZCRAiig1Fp3fRWOOZwiYo4COXTpZnreiGC
R73AtLJGsONZjpcNzJe/zg4Tttc+07m/PkGLhca70pXNp4gJWRZIe9CTG5oG
P19bq4vlccWkUvREFeRYwswQJBH7TrqAw6lxTG0ZVeQXMxl3g/XlRZhaYKXa
IY/94kpeQ4Y+VjIlKUZm8EjVyVctVZn9J4R2+4CFnbD0Ggtjf5I4aZRKej4O
z9Kqp/5Vn9LVDuVzu3OGMSCs82j+UOJXKE7VqOjb3u4iGDuqjyeDUwMsG1bA
4/n0bFCyQRtj/BgPFD9pDrPAJTPMK+X8SrV0Rk+epeuyhydpFsab4dLk0tQ/
EbTJiaseirBsQtJHnG8Sde9kNKva+HhCwsdFTkX/U7D7RwyEU652gDHAj0Ys
vlHj+r7qqsm/ycM8B61y7DhnOiY4l4+s7ox+wtrhKrPYyc/bhnNhmlblsZL/
DFq19jHzVtRoxx66O2bojt0I4SSMV9dm06k3ekalvKvxC3nMjjCft81p00VT
ENcqTn9j2jxVPXmI2YITUUX5goAF86BT5brlWNqjtHfXpsfBfy4B3+I+qM+S
OPw4LnpYcAAl4nTQislFqAbQzizLYeAbl2yeXNxEeKb5HMmSo+NTDm0lZVgG
2VVindDFYyEglw5iN6NonH9kWtiqQRs62OOkxtZDo6BrWlEftOijHjwCTlvF
UCVjyNS3+HlagW/yKUO5BcGedfNaX0oezr9Akg1UuQopKzflkx5Fk4bRDrNg
zaz2Mvu/AVrCLlL9LdwK0577cPtpygsv9XOthn9lRajnL1p5V3zFmq1RyMBJ
zsC6QwSQtuF5toMat05U8GSA18ngRNNqwlavEUXvwb0ya4Oz0o1Mj3eivwlb
nmIydhy7S8QZm0yrVMeQEbTq3aCQtgq3jVUbknQkif8jkHW8C/pgd/CjcieF
0mfNu3SwqmswDYbqmqIEPbyvmk5mk5rRrR/+hrmrUDnDicnbhiyed4sUo+L5
ZYIa+Nqfa69JuQMsK27XrADadFw1vMRL5U45WsbDlS737GZHmb6zQJ7KjhBT
/9iECX4A/FG7zhEopFX6GztImQ8mRvCs0nPgoyaAznzXDnPF2S9QCqPWZsBi
CE0ixKnqI/2Pk9fLx2zSImKFOx8169UAU30x+ZlTPArJC3f885xj9OHniHDY
maBtEEH639+soS1WAj8oSt826zA5xa8JvpODkxFEAySYvr/Ab3bYZm5Fj58F
YCCmj4ItZXOFux/Bl/4Y/5wYL60E0boqtn0yzpAKS39amacHfUdvVFMWf/Hm
K3gEA/WAInH6y+FVY3J7PYCSt/utHjdtFbDJEE9WlMmKl0Fbw3eifdFJbVLi
vQ/cBT5+LCnwA/7xW5rx76NL6vUJjmUrfJesT6QPpZsbcr64svDATajQOcBE
2ss+Ff5JC0wsphMUuOhgam1VlX0yc9ieA5kdGFV/CFhe+qh195BkQZTW69TT
VhfKZTe9SC/+mF8iOl9NK7q/16S389TskiFR7UE3Ii4KnV1Qv1sA2SSc9gaJ
4cxWNJG50LsviZjLLHrST74Z58vcQe43tuDlFH+x7MkO1TaM+dRBk9EnvOYn
8AJCXrk7ggio1Luf2VjfEIwO5HuEo4rAIwBC63kAdBIVLc6FR8ZJeAjtVVAv
43u8mW8TREcjR8cFLTi9C4zqLafaSbf+8klE7Aw2r8xPLaZGSNzsLpn/yuXm
9XJxgjCOWFLT9RLwgDFcDdt7QqIFtOyIUiUhMyNkzJ3WBd53Y0ZCVl2jekyC
7bWkQK/LEyi9inCFNoucSHfAV5VjthnrNvJWNFntmKpHIlGvSly5fJu/fma+
PcH2tdlptjX65k+ZD0ta3Z3DLBy8H92TQpEOlx+eDzNQ4zssXLuircdX2JK5
+FPWNVpyiYqs2CfVZzvVdv42g02+tNBQETtCtrmR94rv2p0wXEM0e9xbxg6P
PHIdE4PaeShEKj9Vl1ocPt+kFAhkLOwPm0joBVw/qCHNbx5haGO2qnKbYePj
tLNQRgcwyeHEHdUo3LQk2LMab5CxeUm0wVtHSSG/p7X+tbVXrGerdG9Kwbdv
u7MdwW5LLX3xEg59E8yNJ1Kr7cXj/dhYPG52NMWfinpnmpkw1vzfrMD/n0/m
pT+p/jKLeGXSSk2tJpFjDnM7rpA+DVJy7HleO16COEqDhbQOuKNQKl9dWxiH
9YDBzI1d+K63JrJpqT5cG7jljsMFk8mkMibtiNbcv+bZ6rmgO4+QieDCxx+b
DMvQpRCcZQ5eWipSLC9jlcEkqIeOSiKgmtkE7TFHfwKg2tMH3XBkfzGqIOdc
1BiqNlaFicFQ6RYanYLhWeo1Bt09eR46RlBaU5rjQcszout4RfZQ7h2PLA2u
Nn3QXF2fWxeeHq54RYJVYW/89oELSKk/94GMzLrX+fBS5VQDzY1gyfVThJLP
go6NxNTRuoSGHYJaJ7eZFGuqCgV7HGaIdkPWKpfDRLI4hSJNRVHug40Tcm2v
9Yzs47rMyCQsYUfb3nyuUIhhmIBCW9H2Au4Ru5c072a5FoHWvh57HukVFjiP
vDpCaMuRRXhC2ukD1UAjytM+bwnJTyrHari727/vR+dUbXRSYBXN//O2Fwlc
W0PDwHR0Uhs8KMel6iNIv8LYB0hZK/trj2swYoQfAPYIUzmCbP+CMMVIZFOm
V1mCFCvkWgGJoTlcCj9lrsFXInXl+9Rj2SN2Klb9ayA9WT+5XTrTkUWhDUah
GKf+gutF/qOOYbIETiiJraGdq37YOI8qSL5h28fQhi4JT6m+hTgYc/I8Xotb
idwEj27uP2CrLfFWGYT2j/pZxWgSYTtjR8bEK2kxr51Xw+Yam5IVbDsG69xd
ayoTq9AvUA+GVONgBTqE4dkOXDe0/O1lDXG2spGOAfwAvCW6V2kt+WX5OqYU
fCWxb98xluoquwNH36500irvoEayQby26/DhNEVZdg4LwM0E++0S7nA1n1qv
ZkFNhXdcriqW+acFXJ99ifx3wN3rgbSWfcD51mKEpNSBj28VT8tGzcMgwUkd
8EKUVoPW1z+zienGWTBlHZT/l1O7Jm6BznRmi2cXBtJSM+TUauVtnwavUAs7
Yizaqa3T7fLa5Np/uiab8yPk3RYqQyKD9DrzFqhEg9jOeubXpdb0JJeZVT/P
zm7Yabw0hMyFSdhP+tPCWHDiGyvN6VWkakaPN75sinLKaXfRSEq8E9ARnvNc
vGkZRQW874XJBzqI2d5c1qxenGkMHoWKt5MSq/uUVwhPpuso4usi30fpGB3l
/oQbQjQFfX2T0pSlkhvz0MH2dLrcikCOwVpFA6mRA5TVZ2sUOqYsil/Tt5qr
XgsuQkH47TBZNQpoDRri59aQrE0D4talrDUB/NMaLkUq8sU3KUMkunsuqPeR
aHOUjS5pAIvDqirW5QdTE+PWBCVVLD+UOiG/zMdSmj5xqtdLrAf5q4E6lMvq
pq6PCLFryxfEgzm0Nbbwz2deR1ER3CVzmnJSqRVdlVaFZCab7dF1GlHiOuHo
eCAsJcGnd/RXpAovn7lBLrrj5T9V5bFQKCRUcEQY+s5E+AmxjBrSrkN7JaX9
vPRC4W/a6UYEjlEltTQ7QytbgeLxRaB+2dNeyrX7vWUW6caObc5g/oOMJCx+
YR6nPuWNuCztR2We8f+gaYfueQO4vh7C9wOQ61MtoVKgMvpePbICES867f57
rAw5YLMgsV+XTpYG6iuRMvtPGvq9Kk+m9dfhXJRKwCkoJiRGYQPppYpUJ2uI
MmRBwKleE8D9hR9awOcodX6ESW/xMSzsUW5peKf5sKQzoKSlJm7kPzJP/B71
vblVKZbcknB4onhrfo4hdy3fqct3OfUFeoqFfeALTJuatxFdXw2brZM4cBar
AbdxejT+PXdpWkoXsbw3R9tBZOPBXDA5IjnWaFVBoek1OUMcPGamacf/0eu9
VNmajUYHBL+qp4/4eF3wyteRNDyVutDJ3YtjU56jh1P1rzk8SKAqtYV8O1g/
GCIqbY/D9arYvdiJXqcWqC9FPoyrlvT138hEZns0N/124gniX+tEnLzHIziX
k7nZcAI/Mj1VolPQBYUAl42JJQ+8y6rw8D0USHJB+W+Vu4wrBazTD/yyqUH8
vPgBD/S2IPqD1qNdXpqam0tQRcmRDeXBhT/I7wpEq1JIn5wAgVOK+l/3xUkN
nRfq0lQoKHXSLGRHEuLB+G4tzV3g2c9IgDfTyc1dPbsUcPCIzu/jBg40Kk/u
o5wEmODxB5YJnKUpii5MlQHDQVuEjPKysNFJr26FW3UeuYyOtj+qNHTaWleA
UirR5U9h4Fo9y+SVk8cHpuBR3S49TPUAiG0aJiinjj4UQy9NHbmHFJBcDocG
CxyA43aGqCyyo1Zuu1TEX984aDW04G9zqAv0PPR0AvlcPkoAYElduM2RSNUx
qaTbRl/hBz1CbR/M7ldsx8LQg/CTzIW6eu0kEFPdfIIcWUbDfn0mjNZk73kO
bLd8FhdJ38DDr6U6lpWQIlzuN82xVY+XW7VSd3wxLS+rdlyNWSuRLoo77N0D
qAtpwp7xvApYKz0W6v3WQm13AXYXDnRtvB2wuSQINc2UHZG2tJIe0tT/U3/d
CT3dWfp3pcy2wIUgXntuC3vYImjpxWSlmImvflyH6aIXjGmO6R70RCiHeCcg
6/EWM1sGZTWZ45FRYGzDR/DxLE+MVzfHY2rGQUJhSHwxA5cpqUJnWxu0tQDh
Fgpkass+rWTTCXrGwbpS+3xaJt2/MdlWCf0iRTxSjuM1yAmdWNsOhL9K8sdF
sVEiklNuvffMY+TeDYaP5r2gfXKMJ03Pg3CjBM+X96Au0smSb57mbB+Afko2
5dKOoS38Bv+dKVD0yy7RVizwYdtUQIQVTvw56mt6QdZnVXURRa6EnbEAgr8m
Sh98nXKVbEUSx+bWSMZ0S1CO4R9twmZ2LD29v9OLqP9e5NUHq4WtgH5b0GQw
8LUpHz+MFhk+FkdqzK31X3rKMqfKQUFVjjYtZyXay4cI5TC5kEOu1k9pnxnz
ATUsu2a6TbxTPcZMJ9Ralx/98hqzYpFQkqK/UKd9eGsnRZz16zXz6sfxzlXk
SHx72qEagC8qaQB+vWZLYtkzcKOrieJDXyH1HQcfY3MzvekueP83Iy2WsMxy
XA+F5FU2u+jEqlQc+7JUJJFJV3HXTzigheh5zNoAWT6eIhbtUQKsINF3lr4x
DX63H6BKqyD5gOxg+UuTUL1kozO8F5HpFaXQ1Ez9DxE7OCbKYQv5CasQwiZl
CpQfTF72Dcg5rkYu2gox3Lr+F4MLXILqG6GOuQiGUALMyEE5ZG/YNdYqhhy8
4kv0Pv874OdmDg312HB0zebbydJDyrhHd0CHn8PxswN1iBPZv/O9CkS1gdEm
ar+q4KqbJsgIALLLkb8aTxbAmkprhRoTiUXVQvVrvOGZ0a8x0AKFxJ8z8c/l
AT/FR9/W08jabAgNQxjdoKCmrRTv7zHomAT+JxxUvodtNZufQD/QfdT+oja0
jNQTWjIdJ6LdIFmidQa5zp2UE+fhq3HI3PfY77BiApq39IxIJ7JU2G3z74Oi
xbLonNoW4oKzbdr6eIxIyTyMU/3ncHASJBAaotviL4wxaV0tmjoMnV19eErH
Mk0HvyCN4RHw6ivTvOp9vizz3nd1U7phgmZ42Rgz2ODfFzwpou36TgkwdxS5
9Brfd5TddD1OcWqVDfxglriPWo+NcULOz4w9a/8Jgj0UyF4Us+5wZFCbdNq/
KcOGkT/HLxGkgT9kG51OW7rkezWXHAQMyUUChft8T6twCYx8NHUwA5rgfP4L
csIVgFyS+seXnv1PtZYPpOfACFisoByfl68AwoNNXCa9JXEBHxyMOeoDFd0d
XC/D9Bp0d/jW1mHvydSPQ6mPcdhB5Ldy2IiQFPKrdfYGamxqtEKSfnsgj3VP
fyAEK2UnsGQSFFozjoroMuj5fI52QoB6mogPnlWs0wyI25EbFEb0OE5EsoTs
6zS5ZNKbtv8xWWfCXQnT8ku9cHQdWCXWx0Of3JCtRj8hlN9orokTs+jsznMh
L8zJoPx1vv9eZpg6jS0bn4/blOZN0uDaSvYIZr7QqFjcjQOnT3V6yxTtT+a2
iiUydsASSt5a/IKuy+TmjIgZUmATS+8hZtmI+d/7kSyfDYNOD0+6iQV7RVKQ
QGKKVoXvwvfAZV5fKIP20yygetvsJ1+yrOGLji+h1h/XSqWzqmZtI8HgzrQa
PGfR84rou93tfG0ojRWqEAXN2W+u0IQ4DUGEsljYV2qRj8YTxP8khGf9eRJX
Mf1AGtEqxAH4qP9Nj2OkCZU08PwvDjdZ7MVMoPT37xCu01GCxASbN81j4ych
OMHpZKxLR0NNKCMM0mBmmpKXlMYZdbb7UmOmuyQ0D3GamnReuH6FJaBrGxRC
+RLJNtt2JW+dWiLfSP8pNN+qqhUGh9F+JG7w09qKbHr3sZ2G1opWltZG8fnk
N/hF7cw4EMqh2x1s2uuHURnb71TtMUyd6YSIXpwRC3zQAve6Zd/+p1FKI5Ox
gZFu445zmbahyTY8mmkA62Nm8zh5D/kvZoPEEROVcaOCUjOQP0a5yTXYHdD4
ZZLS8tlXTQBODEqQy0X/dBtHrFrV3cEQHKGH46c+64d8cmxU/eUufHrqZ6T7
XHBTja2JwVWy9kf0u3cd/O/85Mft/O/2Hk5x8ofoN7N9Fzi4ME1EcM98gc/1
40mGfA+nlmLvkVWg7F9mHaHnP1wjswSPa9TzuVQFdh4UD+o9tC/HoKsYmHZ6
gwCba0KED+WbIggEBuqPrZur0ZwjdPGMPdcJRuJTSXxl1KjEb0iersDwLS/2
rCU8a2G/040CGnf5wh8A2OESMyVaP6ezr2b3ja1xL2cGvlkaB4oSfgDPrIY+
RnJAhRQWM8NoWArWzf74uiT3iZ77GM9+/3Ed8i6dY9y2JCFUlXyKaIwTl/8u
iOKcWBiyWEAT2d54vgB8C1y/I2vwDBhIFfwH4P1eLK3HnQDNJReBdHga0o6x
Mxc6pWbX0qLxpZbqQEEIC556OankN+pU3I3bwhy7oWuYXJ21gTlufbjyW5HH
d/L2g0bov6lwbu63g3VaQaFuDKtRdObd97pX6hLiI6fNKPfa4+NT7g4SfEGG
Jrjfllqoss5AKgcn5Qaf7c5q0LBM0msm2so7/J8VBsua8glhdpIhEHNzjZJO
0jEs7/kkKsQU+gLd8cTOrN17mgfgoYcTkYIJx76SeCjxH2PvopoTQktE4Kma
sU/rcztXL0iVtf0u61GVZzLk+PBN+m9+f8KQstnEm01ZEGWZ8HzTnc8ulT1v
7vSpE8fobQbmZ6BtRq4V0X9enedYEEIYVxLPpo1x152E7CzD9fTlsP9/0Z35
w/NoSRWlwNec/gPBqX7OCnjt+4DZlIL+kpDQZVq6FevsZZqvEoAkYyKO7oke
fRW1BNmxtY9p+aaaGdoGluWk7MmMcEc7MAdJAt8du71YtIXoBi/u16Gv6W9T
CAgiRzcT69702wR66T/+Z28u8D1XypCul7bXXkg3UYZgUqHf1nxxQWR95Q+8
lmazb/OrT7y20K1fC1qgD2uDEBwnxyQcrg6JrcEInq/umk+hiEniZdUtxY5d
KRrQfn8hY1hdvACI0n2Jf+DI8jhgRMNJmmFFAjG3AK7/Ah0cla5OszoA+Yaj
CeecuEuJrC1PLSLU2Z8Znbt3spdFZED1OmI5MKBm6W3c+wot7oq99BUoTFZT
DPQ74EKbrbA+AJrtGJbp4NEBIdO/X39zTl6Gf8Cx3yrbkxvbyfErWR0VCf5g
ATumXmSD7SQ3cboqdutuj+bw1I/YLeWOewnUpFWa6YSviKITAhZUOFEEjGPB
Ck03kb9AHRY5WrhDhQbNpqyP8nUF6ncdcyhNEV73XYp4n5rNjgA3NgYsEykL
6nMVvt9JfHPD6UWkm4PhZxxfAj110sXSr60V1jnaIbgkWX+mGRk2Z648iOWh
zbHqVmjCe/Ttv+sBjGCzPyOjINrTc1aYTmZv0DRrCikd9oiTPebGvIRSXznW
tAXius+fO7EOOqCfFlyfyRGcRGQTS1VmtNCD4CG5PvFJIeB/T+MQkTHtJKKg
Xm90n8pRjUtfHiZpBgwzFXIswQwgAxNsUGUWoaou9DRSouQOagWJZiI2SnfU
5Y6Lcq2bwp4pdUGGbOu7M2GXRLeE67CCwAun/SS0ZFEx3+qiOybnllwMFsD+
Bcwlc9dHjA6tU+VFutxs9akqieeaWLx44WLA92OUnVJ1xeBeygMDXgecQM3x
8U1MtUSyw2hDVAGLWAL/gygNlzeihsnSpHz4tPPEe+q6JIej0A8Zi5SEewjz
GAJ3IF+9vJ6Zx8paHmJZ2fUl/6HtfvoNNGBmjlyAlW5esk5hcPRS7wfuf9as
CcJKgHm5HMAihsHFayoaypl4ilDpsXsnHuB9utaEVTvZ2QW2MMjbe7M+6X79
l5FRDde42+Fpj+I+RINmF4Qy6xmTn6iR6qA01fs4wIvm8WFrQO88NT9aIF+r
alYJNLEeNetBxnpBBMwztNdDuVWwiSlQ0RMkI308rs3dyiGVab4iXnZpRD8T
fscfaqJt3FS7KdNsN6egyBE9mh07qeWwTMxAvCLYuNp6INoEGaJMShOoXGXa
ZSddm5f1Fx+ta6RY+na5iq/UvZMlhOpb5ddiiYWIBP3g233RI34T0WEKr86W
/oPIagMOwkRTIO0J0LFdBVDF2nRFcN/OxazEVYzGZX2rYpUsfT2mTLNQhUvu
OMH+hxoERr/++m32k1S3X7eug1pMURsBC09Jg5fmWe5WdjKJRbUPFTi/vSjZ
QP45cEraiZnzf0arq9k0YS31gDWWb8Yq9HANsgNGNFbrucuIQdiMx5nj/WM/
gRXiWEJFda+rcMgNg84EddYvaRTaeU9v14G1Mhezx8PX09p39CXRi1AmQJBG
Fo+Bf2fWvwY45lFz40kbi+cTlSZXTqjxCTgUetL5OyBmtmYdpWu/7O7jrAW2
jzTMBd/RmGmemUrjil9ZFpqGLA+rJH4q1FiQMv0gVVLq5QsZuI3g+w5MLQr0
yYCNRdXfdmjSDocbKKBN1dEnYmNcHOQbjXbbowRrGTFig7BhHm9gCvJahREl
D7pjPtkgUeV/QIbUr37eymoXAwLyttGMLo2/isAZukB1VrF6veCwy+IUJm0U
y8EMIxdVWw5j0vPo72VNqyr+ytZ6BjxKTSGi7Rub7FSWdr0FbXCdUecuyzty
W8IivJUkrWV/bWzGWFXKQhY743im1JmYfsLNDnNJKP5qfEcJoOXr6SZMrblt
Cits5ID8V4elfAT499GuRn77Vnn2EprdaL6JzJEkELHrJoZ+EW8WBZod5RkR
2WTYZhz9++IMR6260roGJwpUIUEX6A6qKlRUT/fQkiw3nB9PU7IDT5OdIbAd
tPxZZVduLbeVhXV/+1qpAujHR+b6WSvKKD7RW1DPCtQmvH+AEFjcQhOt9KUX
d3mKkslRyYP9VMIEI3ZqtEzlBrpOIUc+ouiLqONumC0GlnkuCNGKJoFfhB3j
yZrTSwmXyHWPJlX6iMYZ9UBvF4rqP76WnbK54X2ArsTyX+9u4ms07+y3137w
Ejj/MaehyTnEdP10GGNlXQyfUSOvKyikzWbvFyDe6tfNMA7cPAOu4EOnWWgD
92m63v8VGlyW4t3bDMVDXuYHnuq6JLZY+IYZoJsM3qtIbrxJT8LbR2fomIxT
0scr4yWyLjET2O8dNNKP58oOFlere7cTIHMQfBGsA5mIfPYmupKTX1kjVriA
459ueJ7RT5DPnOFFU1EpG+ZBaUh6ms10AKs0XTSyQJ+7eAzKkgF+KipC6ud1
lFn4Sjj39JBtfxIb+TgC2A8WPdvsc1y5vZwnV7LVe/bCs8bClIafUcJjsOB5
YoZcjguZJjI66CAGYnElyVd8vO9ew8GhoVDE7zGlPCo9XET01H/wt2fU95mw
xZWrBp0ILc1oxocELE92AZFvBpFiemU1+uqzTGiH3GPVH9umbrwRcwAJN/7w
VlfXA0tB8i0BPnqdN/OnsuR5BoeCGnhLO+UAyIfqs0S4IGEnOCpmt3IjZtsC
afGRrsNbkLAcTb5LK7am2MozYeMxYxzineLn8MW3YrQi2BmA7sPmkE0Uo1/7
B1QAb4OXwYN8UvY4ynGDdc/0/NjJp7fyz1cJJcmOxFxSIopiXD/B0/pCH9Cr
yuFvN3EST3YUnEnOxsmjYiUwrS5gjSQW0e0V8fcqOI2IiuatTSRXEfu3bb4A
hKA//bviCORBNzc93GmpSWFRJ47GBHL2BwTLwCeuaoR2nj5M/wJrdNnwOYgQ
NSxPK4TvqAZZWeS+ASzz/6aCcd0JQ+C8Un++5lQbe4sS9rKWlDjZBGdv/R5d
+1JB0UJU5KNLdiUvKz2Lnm6sxcXzXttSB4ofn5mfFavG1+zJfZUw/jX2QFyP
+ytrI+KLDhZyv+M2If4/eYwo1kwypw2Fkr8l9ybRpUXOCY4ufhxYdsv/sxti
7gFK8ZkRRn0MWPjbF7RjLUzXm5MtFBbRXFqekmfC0g9I4TJ6O/1mS+2CmqKx
f8sKCJ+/revnFy7vViW52BTrkmCM7jhgYuvkrkdpDS4N4wuwigQ7ISva6SSw
/92J9UC9rIanGqsFk6sbYcAv8YD2TkwBrNdeIiv6mQ2cuPRXmsZayAXG+eCp
ZDzFgUeupb9smK9/doAQ387r4dlkI1z+Icpj4Rl9kfEPofWO6cmLxawAH4A4
QR9oER71zwlisOsg+xETnnJxy1sykDjfAgmueYs4h3QQlp6Yv+m7Ipi6+BVY
IU3Tfpg48vbKKnOScNmHrfqzYtzH+DM1UIP/9seYKK7FZXB0tSpvELbtYPmp
cKe8YOMXxqJDIrF7VlXv/mJ2Ef0vbjiru6teychkoVuksDM86xsEh0kZ3+VM
3QF7UGTp+H8h1kLirZXI/qUgf2WlgqL6aZkSBLRn3OZcQpPm+NR1kdT11DE8
+tG8BKN4mjFF5HEks6PZW2nZAwgu6nyUZrKCHTgfUGxUk0Vnv+EU5NgUwFTc
FCcdRfRKhT4DRnyCBt1uopjtBctgncYn9cnY5xsANiSnigw8/pzY20t456Bw
3n+UIx5sDiWzW2jKAlIWjL6mcfN42gbdxPEqd85k+ZIMW/N9bsURjepI6n5P
xasoDg5aNWtkbRessLm2H9uuNUr+aPGLPgT1/8aus2AzI1UXrIakzHaG8YZA
5rOnZd36ZF3zXv1wO8XO6s6L7tHBkbLkZPEqvQbtDF4KnjTRH3ZE0Py4wvYn
H1qe3dqnw88/2cIWfNSD0kJjHxjqwci2v84mWmX26VKTVJ8Yz1sctzxPaqKd
VZLgpEidNW0++exT2HHtAAHS5+07oA4Qb8vvnShT0Kw8ZFIqQeNN73cXOO2B
rIu778A1jsSnzdSVbdKawvb9N1Yi3mWBl9Ke7+Ps1pAmUMANnIaPsFhpWeZc
600tvEByEjTpfyoNKSaKXJkzMFd/HAwtM8tvUmgreaIBJ8df7S7E9E3HvRpk
I3zlIEoIXxoI/6RVEzKERLNUjk5EIyWfhhYboudU2f5nSwTvM0iH6tJPl1en
+q4dSUeDt4T1UHAcjpSWc7PmpDu1pqu41A1wuQ5hFpGC5Fjv0MFvOYwMlZ5l
gkv0+dDNAB0J2N3pmNOyqwU+2iEuJSe9mSiCQKPxrTa0eODiwtOHRfmbHVC1
J3FGXvP6vQTmlApAjNj3W/AwAq+ieXHit/edmef6PUGq2BXPeROVXcnnpgwO
lIVvh06C4fk6WHiCJd0YxOTRwgCX6KxhEswN+89uLweQeoHACfPG9d+qprc5
zu/BgO9b0iAGn0iKyEC13DkSjpsPl9d/KkdkyLIOtyKXttzzBYFfh+f6WZMb
HTseSIVUdl63RfTLQhuRvO3v5FdrQW8BgGLoPCX4su6yB5sUthEJmQmu7E+i
ngqK8OeVDLYq5XISIywb0uCp8nkbEFNhyraueBEPNpyKMWaQfKF5yUU1VCqJ
6zPEFBCvydNdj5zLiPChPiaTPvOwQyz28Izr82GMcubtMJUFPVv7ACnhCBx4
Tv7Yu2h3ZkeYmH+Fv15YiI5DYYUU8DogppoT28pGs2rVu5oZ+uutxisNGqyU
nNF1HVqCyRULUSaSzBltIdQdaW//erFVDkgkXbgle3kamQM7++RJSLaoQ4tf
HrF943RbecSHdXCXeQFK1m1IuWjDD4htLpkUZushroKjDozCHp2UByk8vxVN
BvMD1dZOsQMfdT8yKAyqMhSDLHieN5D5aTI1lFg9RhZt6uPGMxKXbNmkQoZi
SxE68VLQkmVPtIEMeOkv7fw+Im8ENFeiALFNJvKSDkwsi6HDoDZJpWTdkr58
s3cllIy37fYOxprCWIWObvUDuc1OGXGTwd1JtESK7B0zHYTSfoOyyEmy2LXq
CxeEZxFLSWGs5NiBxYty52QlwmX4YoeQuQ3S51jxm5tqYXTSarvZdn6qNsu4
vGxiWKf3WvMGPPWT/48u8oq6BY+b/0fZNXysf/dOY6A9nMFYRYVBuvd03CIi
AYYQpBQC0YtsMbeyttD4V6sBLK365fb8DaPt1ldUq029RaMkdKcnr2cRl6pH
9Uwe6h4es8LV3ypv/NVh13vAprCvJLf/dqy9JJ7L1opbUzIzUzAKPs6wvEKQ
BbQZ0zmkfvZvmVyInjjl20Ams2SGAkAnHIEllUAhaZ3EUdessMmsa6D2KsQR
Ya9HWtiRlWCrX2YAaSV2Q4x1MNZQwl+VYZ+lT4S9MGJrK7P9cBTqx2w39ndy
aofvvdrj3rUs/UbuAS8Se2GB1IQglAGkh471RjiScGQTqcHzPEedXg55McQn
zX/nsaowYwfFVVIlorMbtLZmD0oD4C1fl0/xl24MU6To2x/6MndKPJVVz59e
OmSRQ+ginWcLs8GF+e7FCTW7imA0JryEAsfYRTH+5pLx++zxcJ7BIQi2AzcL
xdZSzq4lM11+/NijDKjvJ6HAC7zSrHzleL8bvny5cOAS94GoryqqllV+SKxZ
vLOQwcjbYJLR3ZhPVdzxrEU5Z8Qd8UxHMQ95Xfwer2K8LHt1gmgg9RJh/bZB
ugclhI+4Ou6z1ncPkO/ZM+WpeyO8q47rrRlXDnz/DNUiDxyKDUeGVt5lHipg
FThfQaLmSl4xKy1TRY8Cwuwzkyw0zVtWvLsX3V3PhfoTBCOlMVvitkaR0lDp
jMMnBb3NaL1ibNGeI4IKnPx51Ordo9YlPE8nTNKw5orhA3vzAa2pPlj77T8p
Rv8qYKdESo1Bf+H+WLCnVB9GFSPw4rMuSdY69imgqs3/Jii5Cld749uT2r6x
vH3b2S4HaHkdXkhCV+5xrO9cLTfWtswrTDWgqYWtw9Tdq2qHRgv1pDVbtpQ3
7zQJqCG9isvX6H8eRYqlQh2sP0Hvn3ncddXBIE3S5tmAw6Jq/1fKOeYnDQQN
79YPeBCCvalNDt1IZWY7h2mpsJBnxPeklWbL3On8aJWKz3B2fhPW4l0rsp8l
7+SYyLS/vacxij7xJk+1Hw1EUD6va+EK/TYvbHP8egOZuyF90s1HVAorGARV
d/5xCZXQ9KyDtGbQB9tUBI50BFX+geqbEBMSqYlFBgXXCKxlrbwNdNdSeYo4
6McTyu8J35xXhFvgFd/AMEj5/wQ6UPb/dPdApgDkHx40q5XztSRNdOU/0wXz
Et37hW7MJqLWb5xgrm2a/9zLKeymfLwKqZQHwgGDL78u9GZ/fQBXw0kxIdT7
gDOj+d6gVmjyth5yVQNEo4v9sfIwWHeY8W/52bwt9/J19gnFlDrIQI1O2FBD
WRa/Ajk6EanemJuVwqiMOR6/O06YtGTOsxLp2xVlPXqAOLbFXWw5LBwpnUFZ
g28WiyJDbAsh2xwo3bcyq05I07ycQBjvjK7636fbctfix/vOslFNpxRhczaZ
JIYUhl5VFQoA3W1B+ghLYpx/iTZ+Dq8UC51dvYqvZ5yhEwu//EJltLXH5bxP
Pd/UivOLsz2PlvOASqI9bqwsareT5kOxoxhvnz8sJTramiV9dTLotNIU1o4c
4lHiiConjxGpV6WIKIxTpTvRSMqfuB1KB/+2xYrbUj6+LxSLpQw9RKd+3RJJ
alyFLYPnhg/QtO5D4JYDUqJTDn5r79VEJwIkJtbmZvsabMhAd8ypPwmx7ft3
7do9Ny/G13fW440G7JXD9ttiTADN4a94rAlLsmytsGVbFvu2PuVblR1x4ruj
WjGX+lFV077eloO7fuSu3k+pfJdqm4EIL1ZkboiWGE0CL+NuQm8F9PPs0kJP
uVwMO0La/LVJ6RTvP3oJqknpyIZW571e5n/AcZH+3Ipuyk5y1J6vjol2M+Jz
95PXdu8EVNOvWVG44L1NJClE06tCkdOl7te1bxbqaoXDgAhYuCMXWJOCJYqa
cyqorWcPQPcL8LDQWXWNlbElWxCEtdF87csOCRedzLRilTgnn3frpq3N0h3P
9KgvVHKGRTwC/aESRzq3KWtOKKaXi7nR+9uoI0Ir0WVII+7YlAFjqNQIolr8
I1LZW0GLmIRKPAn552s5JyTljmjHRdIAbOjq9hAh5HQW8h6ZsoeR8m8HYlcu
yXUBVcEF7IyuKmAwNnMmHUFkkFiJb6P4X+qIHI8qhhtYu2A4Fo9dP6iGjw47
tbD2j8pDQajfWdcuV5AO/IpL3b7ilZuAmo8QmLpR65f+ZwpcEohmrYGHk1te
9OcMfgM8TYT2IIjqBAehixsOT3V2/Mod4NEg351x5+YbyZqb2oJ2ou9eDl+t
xgPQf+ZGK84pYBg8+eWX93MScwYQTJ3RommXTPFtRLEj9jyTJtuZ50H2KDAU
6phFMdtApV6wQJaeynm9SaG+MLfleVM2wg2DLvqf0t6PnwpVBUkANGnKRYJ8
vXaqSZnD2ToGB2E2ILzF1IS4VqTOgvnRyCEb6DO5+jp7Jim+fdgvkz+6tAPz
Ve9YCgf4H8fCDNiCw7A5pMEHJB4zxFxbTeZAJOX1FbsXBo0yOTr4DhzBOCC+
eIsB5LXR88WLddcSsRI53AU5ea3zO4TCajlKcBBnVXoUOUnl0LmTUEamQorU
yAwuCAlnaRgnj6jTqv/NUuS5xcZvs+tYSBHPVzUuBV8+4ADwYD4/aXLboRO8
NyAVKr5i6YoDiaXIOxhTMH3pGWW7wZ4/Yol1dpkfck2T5ILzQTzMlt0lgQjC
Dhy/NV+2D5XOGT/VDeJx2KYFeBC5bC05zmvldlMsGjGzNzpJ/eEDkwTTTVWa
E9wV2HCi6Y8Q5mykS5n/hkqqxwdZmEU1peVh+ZrxeR1JEGaUFX8BeMSZMUYs
MmBEKzYxHoRtjEwzU0Qlr/KvAkewTAB7+FeyGHm1MyV65JSm3aroay1DxSwY
buiHB6KUaOVPNlkSFKFXoHuf7ET5IiOE/LLmAy7ndPJ9gbAXHSp/jkeltbwC
hzLWzw6PX5l5z6//IMI3R5ky+iVld9jOmOb0MBVuVm7LtZ6RiruS3Ms/s/Uy
Jsehn9QPGmiqHI7y975ogANyWNhns8p0X9ZCLN/RAOlA+wsoYRLzdA74HBjn
U4XzYS26yOJ77SZgMD1sckHS1dr65zuW85jJ8fhqCJyRFQNFwNKq1WCqmUq6
RmQU/d03kMeKbUypSzfbL1vsMwP6nsntkc7NySil4ZPcGuEh5gGi26qX7ICy
aPrzYewKZEBZqOBj8+7RCYsP/7o3s4x227iatuN48km7EWBhmFJ+e43M+MCl
6+w4RKR3W3pLxd5ycW68O7axJcteVfk50MpOlF/6dMTJ+9yfOlmoTE9yvKPi
m2YgZ6tPha5c2wpFno1PsqdY8MMWPIQV3NKUcG7026ttdHHv2Au341oUN0T3
SphZubVjIyNYF+S+mso2/c9IeBqoO5zp2x4kReB35gYPo4P1bBsgNjgC1/0N
WwjYF01Djk9RbN3BsghpP1Y/QghWLgI/otQyQvIkdVYOdhFJPYjHmu6LUmNH
O6zgUr3IrKMPhZaWEZXxam337aVCyuFb42Byslv5sK1N4C/5HZArcaIg5J0R
UTT9AqkR8mU5klQYVm1XijtfGVI1kbxGq+T6YaqdpAWcSSySMyGj9fGOEhnd
ilrqT80551yMLdZX7qP6IJpHNTWQhbI+aGXRo6Z6YyXHb0pzKhT1aa8/jTT3
lVUy4X+OA2MlRxZONU2jZp3Basu8K8uq6a7GtXBFbyZrmMlb+XxGytdzaoLy
lWFP/sPnejTrAI687YiQ6VDAFfh+DIVZhiB3Rj7srmganS3P36NZo/viYNJM
VXKQaBEvXAwBbJeNXglgqZYpVhRCsn3Pw7Xgmh4clH3bGOm++m+6D0nWmEzW
xETh1e4ha2TJCarfuTMTvO9MsBskUT1xSQ9cYy7SAuphWlc5790wQFeca2t9
m4rvMKdE2FVX5cJcE+KoaE1qfONtD29Foa9j9bYAeqgLvYIUQPHwqoIqIKwB
4U9cCO+qRJCc28KbYQ96M3cCGKYHOVwd9B7BYyat77Asd7giMrEc2t7x2vSd
uSrzIa9xrLC+OSwRg1KauQ/pL/pczPey5E4QQIw0u/lSjs8zg9H/OWpUx1gy
NBBrGjb70b0oXkb1Pssrxbfb/YvW+QXUV3TdGO29AHteFXMpTL+vxYmIQqqO
FdO+whuGYCFakNO+PyOW/ovKPQ4FcvUmWBwoA2jiGz6AMOPOEnrhqKM2gIIt
YibCJKPNrkCS3xxFYvsLNlqucVsA35JPjRS4I9JbdoOa1GyngqtgUUgK17UC
mIcoPSVigapT6t4ZELBIE7IZTkuiutiJ6oEC6w8ypLY9ZXDT8vr8NYWSI1fT
CVjbqeP4ahDKhel6SOBs/JehFhA8yZzXnjCHYd14mRiAhRioWuxTbsUdv8LP
N0XmICrFaEIRVrGEFJfttRrPjBKKxX3EjUCy2UdcZCip55SklBfw7SMALdh9
ek+1+FY5IMeefYafH4fdmgjWRkCvXwMnQs5vFaZCnLXvLnQNiEBs9u36VxNx
KR/LcH6jLLESRAbwaOmG67da+Glud8yRUgyrf/pv+K9gRQ8EkfiaNJsZXfHM
uVdzeIYkmPB09lYGDhLCeCGWcC2Y+U72NAQAUH5YgStI2IJS80NF9aYtLxct
M4qreFnjk6rwgSOuSPWlfNlfz6XPKN0FR/ND7JH2Xq+qfpUirdmRostQe91B
Dt05aVHUeH+elAJ3FkvxuWa1pnz0QRpHAB+KQvK5pDsP0L7veW0QJabkNnhn
Wpmle+b82v3jw9vneD/gHZYcRe2w25I0IHEr9NXB+rDGvpLwd/S5TRypCEIx
qQHFzAGUrxJ95laJJKXnkSEZXkYAzIKXIejLv9JZGJ3st/mFdXYHVOuVlynq
8epgAQLxOeq3EBVsFCG2/YvaCfIvfvHl3xM3pKECc61lmKg7sbVWxVww6jah
qTS/ni+IJHlyR9MD6EJmqmQ8b3uwl4Dpv/HyuKY26wUCcM1TXNAxrRq5v6YE
4RVqi2dVigmMabJv0AtvhfQSu5z+fIxgiWnGMirD2mPPd5ByZWagkSJqQCSC
Kdw2msmGCXY9LoWYw+BFQT/Ne8O8wU2bSpuD+ZYfmk7oRAOlgP++rCApSUn9
BtanFQYz2uFNxi8SUaeKwWKOjDUdRdAcv5CNbKfaGnd9AR5M2Z/oYYr9KAgl
hJUSTlH8Gc563ywUdplMw21uiYJ0D24aySckpxvPRcEcX0vn5kXsvmPYPDKj
0bEdJ43jL8B0oybOuOTqFvbRnLphgkOj0EMKinUGErK/1PARMCUQzmdv40tv
sL2mvxwbw6uMbJz7z5wW7V5r04Zi1y96449EwxOi1PAJcRxEzBK0F560SnHA
5lmffvY4C2GjtZcF2UMn9dH4veTfbr1sdyTKU9TkuMSdPHwC/CZ6yr2E7H5K
gaXB6Jv1MMlBUghIwqeTL+naDhwdf3V+/sYCt5kF4HBTiFnrWwJpz1neW2IP
WXgKjlTIP3x/oADJS3xUb3f4gonNvQmCpRJetZCls3QlzUilesxBmuSW6QGr
gxs8xY8zIAUtJSpxPnNrCmip7XzJGaK+X1xUBLaWQQB2eMeQIsRw6QoDB8iu
KQtWEIioBu0w4yfu57OdATxM+LrTPFy7lpsClOjlxJIu5nQGA6Wkch9gIxEZ
7yeQPl/imnb2xWUmNIUMQIqiHRRDbbmbHxmW7RFvGHFDlHZOvbEOmJxcP4eF
fm+Nmp/KYufyVXU653KLMgb32OWBrAi5rUCZN8g3N9rsyUnpxq4Y+LLCyKZC
DTvrkD6K3q3XmgDlY3TM82VpFfKZPt08YBcOnB9cINl2FEYXCkoGCNKFoQAV
/vbUww2yNWo+TvDpGYDhy51dFaPTsvRa8gHFW9F16Mbkbuc3/VRP/DP30x18
dGUY5vR+kEwfiS0Co+7JZ4ezhAuYaLLRwzyyHLvD/m/5WyqCoBjb7BYektAQ
O+9fRkoMWbjINCR8lSrWoIygX6VT54s2Mefe/QT/mh95xpCFgVod/C/zi4P3
d2Yfyq2WBfTrpuSR462ttxD1bxAfI3L2qneYSOGtSNKqYxlMeTSf2/Hp3r/e
vtPwXpt4dNknHId1AxwyRnGMNd92VDkHK+vgc+aafI7J402PSrwh0t1GkeQ5
EBqw35szoqWr7ENvBh90mOi8aV4bqX3BwgdA8CruUxdsonDzhxExUC58QjSz
+0sIgUlZHdx/b7qOiCfYNRKjBJLXeEVx02ZZ+IB5b+jBHYc+Clw2DS4MUvPU
1rOLFdQGVYtnsc/latF95unE9gWE2UA+5BJsrDCE8NcKFrZcfClfi4Xr/Xee
K/I5SZ75GbjAjL5WESAvJbwVu2/aps37G4CI+kTk3fR1YEDN/f290YfTiQ1L
nKn0oJzBYfX8Bxvkzc+gEkk8s0MzREPO9gvYUMttq8cpwBKQ4izFcwsdYGdV
7q6ydqlw4XqrLTQusW+GKUEEwrt0cPS7C7MZdzgjAkuLAtZ51QV9ssZj6awu
KQG1u5jO9HY8yLZqrdsKcFTGcBLvcJTiRwu3OFdZk4cQ7Amm0/xDrp6T+N02
i64hwjDcBTnHQZ0to508HEaFO/q66wwwwFMoJ/ReIgvjHArG3ugrS2aU7ulB
ZKPJxIR94HeiSFT2YgDZLSET348RZ/914xIWeTPuvUSGKJxqyJ0XqvGpufSx
R20ZFIzEB5ivBBqKJnm+CpOSMI54tVcgGLHlp4v/70+qBU98eaDMCsocT075
DfD55Q0S0GWxAJsKR7ltp32cP7O01MiRk1cvvTiWhITE/rczqPtzM401dwVn
eUdq/6NVPQD+ZNGtQ2NYp6JYTYXA46v+9maadPNd7iNN1H4SIXd8Jo9XW6yC
WyIX6G8dmph7O3a0XshYWmN6gjp25Nd0ppF+tEKlSjbAxkHLO/vy6JjzTvRX
9mPDsS2DxSq3cicxQhIiufbx70JvdZWPzUuONwxhwpPKvGsmITfqP5Ha1T+H
nElENMO5Zjid2lVCYKbxabNe32Qp0zsPXu6QsVxPkyV/U/Gfsw6Kvq3VfjSf
qkH5W/uA+FeZpBf+x7ufjfhF15ID5KsvnTbSmBeXmujQBzzxt6SxNt/Q/AAm
hTJdG8KRhy/23X10z1rwu01bDE1JoPEX6492GhM77NTGBL7Z6rlOV7+EmC+D
PeYNe/tNb6H6I2vgjKrEiFAvUQTHD2oGRDm8hS22hexQcgM5JnZ+hINWp5iQ
3f/09q5BhBD//HWpWAxvIsf+DuaARG2y0xIlnEm/B6R4UTg9fSf59ItK9D+Z
qeXGgZOk736KMGYT1SLwogD8h/gqRsvyLsv5MjEP4pKgDmVZcGquuy/e9TdU
JxnOGXX5Kv2UZDPuSXbwFOZL11EIpR4GyaO107jXjdDFWrlJx6ciMYlEAr4U
PUo0TBUlj5JHr7ScpigSlpWaLvIIU00uTbpCQvmq4pRGi4m4XFMTpYMOr5fJ
xib0igDRhbUrgCVkZ5t48etXkoh3knICuxIoK3mg/wyZ6BpQeQ5W6BI7ahak
GBNHhyk+3mQiIz+Qj4qlNEpEI6rjwPfYfaLJhhUFoRTnAv5YBo/2TUg86TCe
YnJPCwHXW5RTVtnAQ6O2MO/PJD08x+G2jd0dpOKzyqbeJsBEEGx2TDUNdSuU
U3MT3HgjtL5ZEJRi7MWIj6yFNgqSnp5Vnwe/h1DoNgy2LhYz1I9QnyCp8tz5
KtHhXN/KJ3vxucg3KEZt76AITzdbfe74N4vDShsWh6yn0G8YNKu5ePYzbPL4
evC5GYYUqfv2JhETxd8aBhW4Uhj0E3fjrYBn6J1YVCJKMBV1Q8IL3u6FW2RL
YUpR8GIOeVEahLgNcoa+0okeAC39Yx6ZlzuvqNI2S9LYey9F7wSCKTNhZY1b
9DQtRcly4aprN6Y4/PoxhlvcgHdbTosQ43M+Og1sa0a5/b5kuBdvaLUOt5la
KvKDgfFqMyEiPvOfpUwBY6N974YRvtZuQfTupBqI2yk+G3fCxsD0v7vms9my
Zc74ilNiGufGfyC5b7ScU2jAA9fAIbS4uH+PogChiAWH/hgKLkZnn3ZB7xqB
sR2SI4b2tBjCKEoilSwUpK+1+ZNYj87gxz7aZlWa2cNZBCdg57+bAjrjNx+t
HNBYVkt1vcZ5l3S6xbO3g5qP1gEzb6R678QxeY4hGQ7SPEGtEOtWbLXt/QSy
7y6uEQzA4XKd34IA38bdfzhtM0JGqZmIecZGRmUF+nOZJGbnMLNIvox3+/jo
0prD6V1i/tsBbInIEKJLjElcTqMLwQmCBhXKow0rKwAkwsexGi41e3QsHiR0
WSrrIecLzvy45uyR7mV04Nof1W+Kuw1qosP/NzBG+IRSqLFUmRZaaptvwzyR
tAYXsCqi3YPeMbMQFbd3Tf6ymkJ62YhGxkRqmZMgVVVfCCMNjKt2RlHqR0r6
9JG1USsQXnc5RmUJ93UgWQgYYYsXmfpX0NPRXfo8UUEvuvhCeEIEb8S1+5Su
HFODXTkxKssnXJ/XJo+asrxPMaEfB/ZrtpgYwsZrj1GfElCkzkMnKS5OrCy3
IQivgong1DcXmNHOMXVUd7ncNclW6lS5yTe1XhVuqYN51mC08RSqlLYVq0tK
M4Nx/JeOcznxk9ziWvIrQCV5iQIu16BZqezadxzqvknk7JCzVPhIFvIyIauH
kU5nSYzU8LXbRZdYm7f4eah7r013nVIDu+3BT1t9+icf6HgcULyQJxwbNh12
c2aKfGIVQkdt/31jhwVi00+e/wOscPKDSif/OCJfFhiT4angkIM6Y6EMlczb
megk0vWfsnUwZ21vU4eq1qTm8nYJHkokVD0CF2/zz3idpFaNgLuj+vzCDmpp
xoeUTl0n+8Ab95fz38eupC5ZxupydRX7JZT1bde2SJgwklpzdRod7PdBurnc
HOkjIAZm5Wy/1zudZUWPgA3P9sTdIzwqJpCyDu/qmB+wqKhrqFk5lB5/lhif
t3GKqQydEhBZEh2Bgtdtg/A0SXQ1GdlghgzdThlzXPdWBidM1V56vzdEOT3G
pMdKwwD6eQxskOEwU17y5I7ssOuZX6HC5H7gS/6HUkNs7iddEL/c1IqctxRu
uwqIAoIWLdm5HfLWt5HTbeZth8ZtGWE4sxUeDYLNcgwBPcztv0NfgRY5QYky
L+Ao0r+qg7C4o1S449SwpClUre2jO97BckOYaurcwAwPucMrAuFgHNzuW+Ow
vC0yjhB2vC1bEjOTjXzg7vAk28Cd79xYKT6JKbe7vinGenzoEUSIwc5dKS8y
09CFzeMuWDiwp7XNS6Tccf27BkBkzCc4jWV+kZhE1nWU/WnWH2tUDU/fgeXG
F+BS8t89408XpyTVZ2hE/yg/tAQUyqMU68xFV3Bma4ACKyXn92cx+/JuZw93
oy4lA1DSRw9Th+5W4a76Ck+dg0F45UeiEmJNH/5OMZVwDM29buY8l4QaNZPR
TnLOgj+pLPcbZw3s4kHmz0djZT38seo/Xi2ok1hTPLsHMCCwPV18HH12HbIz
tLeeIyKu7YBmZM8cv+QlR3errNTZKieWuGb0BZy7YvTn0G6pWTxBGwvmkLJb
8nMVmIG44qIxNGcNsD9SfKXcuiCXTPDDrWQ1NwzQbz9d/Af80/kmNtdglA38
/kVWiuM/zyVRpgLHcRMdXREr3DU0AR52ykRrOZiuqMJiGDI+wYiAAp5/qq1E
+85HNUE5qKPGbCjFNo6kpesDMJz1+rMHgg7ZSLF29WFYHmZIjviFLfWhYvnP
E51a+A6m0O05XDxpsNsoCU9dm1SqT7DvEY/VvVoOMH7f//ATqyVHqO/4yqM0
YHGCXOzzhKwLRFO3XAow4FMCg/MBjdwsrC77CnXY4Zo8h5KQFtt+th5Ny1Iz
OrA3hoi3taVS3MaEy4TjXXuBtd8bE8LfP++GwjQe2bl4wsTA1VTew8ofCnIg
TRPr/jnRDVlWz025dc28e0GwLPjYmwaqfcCd7znoXhxTml8PXVPfNkyPXRru
CKpdCogldzcmlUY0LrJP79CL0V+be5VQCqsX5ThL77aEibTkd9c83fD5W6Ok
UcuVwe/Vb4dTXhwavMmFA6n0SI128AGwj1KFk4uL7RXHJT+oCtBOYvXC0MB9
sC3vsSxeiMf9brJc06gpJREFx0jp9TRByBz+NSwh2RY+Q8v+CQaloeotLGSr
rjjMrUvbX9A4qm3Z7OBWsZRjdG8erT4sVq4c6W2CizXcCwFAkISZpyTmPlRA
eDLlx90+HRZGCUQKnMjXJApG2mcDiVakK8GFeCUCt9u4jDpLOO/WruA7mLAm
8jpBfAR3dus9Z2w2JSNmFPzkSkbdio+WhCaO3RvnD9catDRx5FnI5gff4dO5
mZV69dmZ9W5zGciJy6n2j9tO+cvfrzyGCwE5dxdDQVJLcCgXesF/43iRAm6M
UaRAefzVmRtxQFMp9B+DDBmNefyGS8VyQzsm+ibgdIr6ZL1X5x0Ou2CmpDA4
v2xaZj5DeAlCdZAnaksIVtlF+qVuc1YmdN2I3bahDp+TA4jieTwf8BUIfRqo
PCwMGF5zMNB3FLsQqSqVWoNLrKgBFEIWMsQds7w2r0kF+9f1PdIJqK1ng1AN
bPT9VU1uXA9/VIPs0eggZ7Av0Hu0Hkd9XnHpWaXVpFuzELt+Jf/5FGnj1/9a
ha4LqUZ2fNsaUmlJFPmikQxjdoE2ExNEKXei8M4B1CThlER4UMGdoEilPCDY
h4Pi596GaOoMHVFXF/ThEQ2F6FZxL8M5yr3F2FBFg7x9NG64kfYJid6CjnkF
JCJXKlOfVYwe9a2lw/+LIP3KQkey1cGYwU8PXA7gJoAO85kC2BhIuC+8XbJh
EPtCp9nKVqdVVJ+oaZ+YmsjrS1ZVIIcweRv67rUNcKi1SDvVs8nNGJsE+oyu
bntwxoKXKIQE8Id7oeszWVc8TdVvbtDfNU2HuZdpSgYdd7BteFp8nH8mtt6k
gcb1Mi9qVvCBLmzMWJTM3gnLYkkuMbP+dXZTwwdboj2XfPL7HiIZy2n+nok6
JkxiMBUzNUY7kUFSuCZgs8BhEgOXqToLwA/eAtVysTCqOWEKKtaHS7RKN26J
+i53R6pTrwHcpc/BW3jGLZ1KTtfdR29rHDk3w8eblgM5sIooF5CklWlCIbXe
7fDDQZ4lyGSbOndhzppdc2SlbU6AS0v5dxdRDbE/HLTFr3ZADeICP0aAFZPN
i8jHylhYwY96EmA34zgVkVl/SICfdAoAc4Usn4gs1xV1S00JZihIjRYqeMsY
ne/PMOypiJAtbwU0RvfuKcbntbQ8ALMTbEFq/uLo2D2Grg47gccPouxHNMHv
oXCfHmWbFwTXhVE+JZDEsONVZ8Y++qgltGw1oEiavhr2hAWJxRnZJH9ihkcu
UxzEcGueo8jknko2QuSeUthj+1C8ImmFwzZ4JnK7ejl5TObrtjxzDMjJ2L8v
dzSVOIJX6ZdJnTwJHfRSzKiZKZimsu4mMh+nLs7LQvB8+WT79tnNdAa7HAnH
K3YnvtyZRHKpIF3mjzoH9pA/z6Y4K0WsddcAHuL0xbRLvd4h0LI+UC8H6R/0
wDW10g02ex0OeuvsgqaN5IpdN7L6sjMZKDIOxkEIjBmF6OIWH5k1Wb2syBdI
s1aPWHiZWe+loClXWpUlmhDlQRYUSOOyoy++w414F4jau3pshWe0n07F7+t6
bwdnF7l6mq16s5ybgQVjXX4JYR8YrlPXLjKvS9EaW5tkDYZZ6RA7er7PlNcX
TU4kS95aSe0wMmULyxaMxrhu8qxVVeYcNqzqQTtJbQFwhWCt0wkTpL7DE218
3FcyWWH4AkxSDt0J8uVVNCdkq9sSYY7DLgCQxj0s/m8TIlLNvN6K5/fG2zRC
OaBaU/+uWuLzqGGgwQuu6Pbtn+BP6HP4aQeCZq/BhmsTp31OVv32WLerTLNT
serVrVGyUck6qYxotPVnitm1ciMFwMqFN/YpXKPzLQcRMK4GyRGaHJvvIPX1
VjBF4ZxY8TRFVE7/sHjPaPAloyMRXO/3BemHqw1hYc7PqPv+jBuUeIzgozEm
kVYP+RlnPofe8AL1b6BGcFiOZJIOQF0EA2ltAyxOZFwJj5HEm0P+W01jfnbi
a4qXKKx2UyJjm+6Tkp20jmsJNANS5/E3Quu97ZYFl3qfd74gcYP7VmVP0HeL
pzE8iCggO5mBJs931ArhyfZYK4AP26Qe02WV4PYxOFnqPAEN6iFvZog9Duev
O3TV5vk2CS5GBRKk3JbbK0OBdxIqtxael3D0rjF5pRlumS3NdH4GkXynuV70
QfJOp6wlqVKW7qwUVaK+bYEypTNZ2ReZMwIz10kRcWLsru37JP3SLjuR8pxJ
OlXDTZJ64XKOsWJgy4nsjy6wbYMnAmcIolP01oY7Ciz+cio1RCRxDYVV7pDU
mQNY94BGClZV6XbNfCMNdL4b1DxGzZBLj70YRm9YM5s6e1yX1wCJgRrUJ07Y
RMIgQP0Px7z41e+sihFTpWdbhfwEOAuT6OY7VB4sYOydtySsISi3s1Tlsl00
b6Ig7exNo5T/u38tUu3wrDvV2OIHzST7OhgrUhpn+R30G7n0WJjxbiNZzynI
/sGxZ6tKT9+p/408c9I/noFX5TH9nlbqyT/9aqChYeqH17tbreV+8BFW2u0J
GkrzrbeeNYFeVJxFmRe/URRQcQMwSHVFkRNBJQlGOlzCAw2XsXXS0aSlaIrf
5bqtN3FNXjQuilIMc2nPxllTnZu2wKdPyeLtefrpMMziGM9UrVkR4pV1qzc5
ptGNk7cULlAXHBSJlfUArMfYcY7wjy5EWOOYiiLD3Thy+BWQMU50IH67UNUz
C091tnhMSSxHUjKWBMOvtaivj+y0h9QeVqRzk6KkBCTi9/xfX4TqhHkpWQWT
Hyzoo4O8PcCck4STeBlZm3gfRZjSrJBTgei5eDAWGXFAO57COvRga4xMGYFn
5Ky4yROHXUaUKaxFwTsOwT3dwm6evjkvKVuEpjLHEQzbhZEcPWm0zDDk9SEf
7/JaGi70QoVe4c2oTU60qtKduER+nREvYOGLc6J5Zj5D0Z3ApvuMWb0cLlS2
hw6WhxrNBih6bFqIXYoFVa3vlnKugo9TSzADkspjtAa06IanhcZKcCzaDo5B
2E+6CXkdia2du0FlGxY3h7BMyhGNTuAlCi3Eo2vrIuE2ZlOsI+nPavoa8oFb
54o9k4XlEYBu7HewqODFcyTSygy1mQC0rU74nrg3jGtYT1Yf+emimGp+WoPR
sVQjBkIo3ET4d9UOWhiO89Zr/eYt9UtgtmPsqhqNymv3xX6w9aPXCEjLYM68
VxnBHB6QA0Th4A4gFn135EaiFIf4BTHZvghzGkcbB+g3JSOWqsM3MmbG8kDH
1k5GU3cg2V40JIGfE0vc8iaVchmmApRB26iHnpreouo9oF67EQUIKS24R1p6
2dP4L0FZXFER870d2nBhxLV+ikNbly4yXm+FuRuzlOQXgdaJOkaTYq04hyh5
W6NQTeY7CN98m2PWSKL9wuOcMeVFD2AxBMzX7ADNLSbsZEhruW0e/h6PAU2s
StJtMuv4KIkzY/haFPwabBBV4ICMS40CgE0BPcB0GU0Ni1XdsD4Dgtnd82Es
2lujoSON19ApKVOLvOdG4KM2R+Xqqi5CB2z1ozaFKjuokVg8MqRZ6sYDwauQ
h12HXrCCXXX5PJ879ai33N/iRwjFE85hZ324cycNyvAyhDYjpLsYNRK3Ho3c
RwMD2BVPMKDPzLMc2YJlpaf9OoEv3jnJDG9U1B7+YHXZ1YNf37INFOyKixeU
+rwY1jRzPZYDtdVmpVG8EjbNWzMilomxkGSr6EnH8s5WEumwpozOSyay3GmH
v6pcnMtoqRYnAyzLnHghr4lrGWgP47zU885ZaId2B4QwxXzUunqTp8t/HQvV
nfJQ5HaEc5w5eeqptTmCNLxgUyP5+9uYcD2i8d7A/ECUQzZPcUo0gwduex+G
NTerYXlPcc9bzeG6KwzDIKleTn8TD7sXeDodeVk9RE+g8skeCri3B4g6vzHy
G5b/bxflY4K6RNnLhXxwQsLt3a6U1fbeKd+pp60qx3RBaZ1zY6LJgsvnLLJv
jYP8f+fqxpO/+7D9sy/GBnPcsc/dMjKxokSpiZMyjK1vSfGFuzAu+lNhrBPP
ujZiiFc7wHphgi/N1ObNT9AXw+uYw6g6F2tG1ePT/PBxTbpJNXi5v80EBy1Y
GPdJVPJypSwxtkPw2coejOeD/hbS8w7BL8VO5CbojTMJt0oOyrfMdg0OPZhR
juhYJhXTUFZbUYcWJvDTXjoS8og4bj+QquPPrSJmlk1Z+l1XHtR8gYP0Tv5H
wMqVuu5Zz6XHyzIbgWqTx21mR3/ItzQ+TYjpdFzLhitdvK7VRCgI0d7fd6t2
lxMOjObDdyxpKO/I9ZfCoJZIgJ8Wp68z06AnIcuWDCUruWC+E1/AdlJPmpAL
hmJHTY5eUm0e6l+c1jvk8H0KP+eS4zkfDfC6xegMmZAvW9U4OB/+BdlZpW1Z
Jle5tTFZiNRMZnBDA8b2b3yw/Xu7Ow5WVO7t5ztXrwLZshvfuGsu/jZKMTuT
jO3JoHLJFwjKstABybaMR+7PmeGVHNGOLDZiQ5P442F6hcFTJCh06xn2GCc4
24Hz6SLuEQvdF1vV7iCzHTPu0rzILSVKLIHKRv0aRtnQFwCyw9y0JMx0LSuH
wguGT+yjm7jK21TH91p+6il0R21GlXdYLhsgAIK2sU9jGTHhaWFASf+muXvK
Xs5j8G5kBbaElRKQT4NnuZA8OQnLCzdjVEEeOP2lyUgG/mIBqX0p+Z2JrC6T
oxHopVyk+7BOnC904uqbb055DprIGQiADjkn/mVHcki4n/A4h2kkbCBiR0Sg
s+UOsKA2dwsZzs51lP902VM16/dAN/U3MGppwEZ8CTDl2mf7WhGGDBXB2cEl
Juh3zqTzYVOzXAB3nBI2IBlIihtYV62QGZ9XDT6wXW3XyDY977vIuMZhH3z5
F3YcB6ZJwuFt2H2a97Ta8sci9ytKH0CYDA957xuYsCk2nuNqwjt9CZUzUidd
sNgS72kKZmGHAtOsYmNlnNtTFLiBXolesCd6tLQU1VITBYnYdEsVpKI0yJCs
qNrMz3sZsK6ZcSwdaalku8twT5GUJ9C9S/55UMYZFSmlHb7wfI/vHKxMZriH
n75ClyOyjkXbUa2fagRG+NfxpeO5SnA8KEo6nxIBMVWHvCxterz385UaMqgT
S6Bu3Tv2hRq6lFaBSF7PKXRdtzq6gRRFgbQd1nQyNg+vFiMPTmKuDcejeaJT
fQn8PRD1Y42DJnicx2f7svpqO1wpbLy1qzEtm2DzfjWxgbUuoBi/HsfR9HiI
FYvrE8INob+Q8Mwb7vxwKLlfMaa75WyiLhPhbo+iqOmAniJQlUcRUzBvzMVU
YYJcK5oDnMHVFtF/eqYEu7hmVUCybbDH5o0IevxIzGrCZY9KrlAeL2EiG6IO
xyls/UHJ3S1QTfR7sRytZNitXs8JCLE7wp8kdsfhTyDO9HAiWmkeMhg19i29
ggJ09y4EGw2hOuS2pIq4bXzk7BhK1AdrwZm9ffLfxe9l+/glzbdcOEL6JrA/
YLe36Q8jkBOZvqUnh0cegPcJCrx90wwVFg1wALa5aUO1SaBEXCp382T8VDMs
ljhiZg8WBo0LcNhSdPh9XBLr3vGcc3g4VCBccbIWLNmuOJZ2Ow702CVXVfSg
iH0PCI4inwwXkYOLSV10iH+0qmJB8/K1XDY+bkhWunosAdsBTOsd88Ak3kQf
NbgGI86UNCAYMujNtH+OPCcOL7i6tfkgJlAU7RyIpKFwcFYcfg85c2mkUcbB
Ipnw8ohK7ExKdTxPdWURtpU08myadltRTCoD43cHyuin/ptq5QRrYQutBsE2
jZ9NjcrjtzHBwxKr+Xrt85z4YL5O6kYxHWFBrz5alTqABqUl/2qwkIIlQ8Mb
cANlvwuhWnJOTH2lTYl+4DFy8AFZzjqR/hW9sAyJprhlk0YVKclekIwT+1Zk
trxzABJyMqYft6BewLoWPL9Agk/6AHsEOtRqAaM43OHvBJjXts1JeHHzIB/Q
xuktJmyufuY9kr3jv0RF1F0QQ15eMtoLx3T+XxYdyXiZWQMi8qtPRqeEJlt0
GGvV+f4asHQ8RKC6e7VsawgDiZ6KAjJ5z6KONhJfQLng+9g/BvKtZiT4gwdC
o/iyeXeBZ2pL9Ft+5c+PWhqpnnvdyNgoaQSwlmtk17OHAOnszdL6MDP6cC7z
AwKmbHkOaNZJdb8FtGdKRxi3S6C68uQHxFY4ndoGalUv5bvlYNhTGswkYUGG
/Fm97qcIOPiVOvbqsN/q0xkBWeUN7JIVLFL/5GWN5jvhnL9fkVjLGRecK2CM
YJGrTZI27nLHaF8mesVt8Fy/U0dv7PCIyylyHA9+V8iNFrpDgdf2QX8xC3tc
S579bUa73iF7iKtenmkwM85n0N0QWXaCaAkWaOW1tCrhySdBTfAvBxZY3Ygl
u+1DWN3ndh1OysevM/tpiCji2yntq4InLFdVGYwlffyDn0I0md3rTO7TfyMW
yFsp5sQSQf2CKbas+SL5h2XIirw7tJr56Bt9GVQ0/s6wxwx0C4gc279GO6Rw
lNO6TOKTxz5OlauG5gzM1Sbz2iBtV4UNYa1RxNGvHys5/Ik0rlENhhHM081g
5E/ik1dMqAsRtjUGnyhR9ixtVocPKWhjqxkJHuSN8F8XsFqLccW1AVzdlAgp
u+XB+EFlHkrJ7h+VKfOvIYky0et+U4JuIYyF59wYx/qT5PiBP0xnainH6Zsp
QIF3B8GA1S/PxSYaxjU910+5FW4weT7HppqQcbPUBWos/obZ6AeR4epHYeB0
gk4SUqmPSku9Szg3y3UNFCKCTZeFgwdEbNvXo/aB0PXDKj/jchklkwrxhuPv
ccTiwxIzIyqLfcPTZw2E/V2iEwkGpzLxVFEH/2BRWSkERBl/z6RcJ+ra1IWi
qrf/1VYWkVYzuiOi6YOcOwke+IN/H/hn7U4XkTb5JKguE1L6CDxewD6mdmx8
FozlicPF3WkL2j11NuKy1x+jdEB3BG856xDY9vEqL1HKHWqJ6AkdOlSz5HP4
NQb2tc3DpDIiOABz8ZFwMcVbyYRe5ueCkwxF6FMrI6W87Ewu4ufe0ui3ivzR
PKc4WFRjxj9aj1kuHbDrhkwzuT+y2hDrHWDdlFZe+U3rby/Oa5KvpoFFHYma
k/c+6P0DotXyjaleeE5Amk/XToYh1cEFi+eBi5Wd2gO9lE/1uUazx24fefGH
XT3v2t+SFvRs4OuTQt2yh3KPqNoAdH86e2sEjetp+6qfQmSFoe8HR6U2TIRS
xYaEXm7wfAqJ/6ogUXjZP9BV1UGuSJoHK4/HX67rnzzj4XKgj8rHoBXfGITm
DqtYGlceRcjk/Amn7Ql2qvqn/+uMAQbI4yESbk3i949cbx4lH8Otj0FoUup0
9LNRzfh9AoIhX53OhBddMN8UmPwFIAsF2Y+4ObSVQY/29d5UqWlwW88oP5eZ
aij6pRk0P8xYsdfU7E9VojLqa4BEq+U8/2AYNzhhP+0UKkuYtHAf9o3lPxGz
OcrLAymOOl/3bowZgzlcASraQIIwg6LS0P5WMBYKFcbWNTckJDrjcw4njgvB
yjSGl9AgZ6oFdhzdYNJM04QBxph7oS83xTxVkjc2U8XecZi2U7J1Wco8LLmc
Q8yRKBRU9S+SSFHDB8Q/NwwiqTWUtOPDxeris3zoUj1/C+TmpCcs7OavHpz3
7ZitgEqR5jDHXj7QnVJiqxK9IQwwfrMJk27n8EGwkOOmBTqMlr1/JtoJSPHJ
8pQLdlNHMAnF2Wke0LqQBavs/piU6ti+imPH8YySHbO7k24XxbZ5NS26vVMr
aVWtL2xS7Q+xAyurodJZ65+1DP8/TuKdPSZi2smbwYvlpb29JyO9k1osku+B
DNzorsiDigIH8MxffKWiWjtswpGpjKwFla9JPYjmGwuKMo8jo/gEuI395M0R
PLSo0df1onP7YQDwOyxjB2USuxj7Un01rGWEsOxBlrxoT/zu76n/oq9CKQxz
8o95OedaarPYuoF80c11q8bVPhS4aB9kDzbOx1M0DjRg37ahEjZi/LzGKmR+
yub4Gs5AQWz7nUJ7Mxk4FQuhvbuOLPQrymkdSa314G9M4It5z1+mV2EgDVcb
ST2oY6nA/caxyKYfohSTTvTD6ndnaVeXg+Qe9dpRODUZqXsFRsp3JAXuoAkT
6ClDYwp6Ve8o9Ha+limxZ5t9kuR3SxUwuYoKDjI5H1ozwDGseYPFU94MP5Q3
byNhpUIBzeBj7f/YGp7cGUb351xqlpGClOmyxQhaskk+367wbdbhcu2agwv6
k6XUapGobRM/GYvT5qFJl26XirPAqiiXAoMTUNmmFhTg/YC0efxpeK/RCce7
4tyg32sRy5nrHpMHJUx0dujSjtbauhMKlWMWngIkDOMoXzTk+YM9E4v5PsK0
HHHl+kEIM+Q9L1xUyB73LK+zkANLABPjudKDRR0wssxeiLYHbNjPlYXyze1E
CanFqHMNH1t9zfXjxNGD/kNKNbd5Jquvhms2F7GuYpHhIn+Vvu0Paik+QI/n
fSMPsFszLatCsCjpCr0xOGjpLv2XnkYLh4PMe89782aNEnkh7p0ud8rehaVo
Ei8gcVJy2RTynmaNmaNI5+Qom64t3PfEiniFO704SS/sYJaWxOvOMyJOZN7g
wTJjmByP8JqtwSdaj/T1aoqKMNAcWhIBqvYu/mwop/tgwfST14pztR9Qnqnh
6LUCC5sJbwKcte8+PfKx3PrF2xcvzr2Wy/6QSpKuL2H/K62L6SLW7o58LolT
TecQah8bUUgxx78UtMqNXKm9O8FvxTtWBM0p4RCTGWIWCvGO0PTdE6zsNYuZ
4pgl8YxEyp0p8Wfggz8dzmt/aXwp/LS6jr8mTc9ljlVed4xPTSecaGsZuPH7
m9C06qSVPrLyjTQNU4P2waumm172XuR/gmUJ30mqVZjfWs08x3is8tmnHDJC
oRxtXEFazHmzehhch1CnTMOqsd3ZvbZtpqDHyAl7Lrek5FqZoLRPlZ4slQ1s
KJqJX2XKFhUT5dwJGCPdaFrFj04WFE7F/tFsd/cT4vJs3kmO8HI07KoN3RPM
5nhq1lXJL/VBKKu+nktMaFatxNL9dQEpBREZSkYWnGJJwqr5N5R4NjqH+sYO
9yaZJlRqhAICJf1gH8dxkic6w1nymMF4CrNHfdVQ4AGliJRMNXYr7qOm4Dy4
KxNp3XXZGwnFzIZQQSkRILb6RpMWbd7N/U6JKldCDewmAILprBDmc5CAU03d
49g1LlXs3k7iyAnDXMVlh9wqynwG3WAr42VBQTslOLkS172w1A8p6xuvTgYu
r1B8j4nKtoNCw8CWsL/R2GyAxTsc1xOImPqubzYooa6MBiwlG4+tE1PZkxOA
mfOT1Z9gV3loaJ8VCrvWHWNmzULUdtUYBJKDwYc++jJyKfLdvZJlqzubqqeg
Fb8VN658EgHRPN7gHeaix2LQwB4vAPPlnt/KH1lMLrmiVOuS7822Zf2xtMTb
j32N/O4pNwMXWx+tZtviJ2hnsxKWrZdDDbOQMxS397H4CiZyvM+DiWYCKRW7
kd6uBhoxTbSfTUKqJAB5Xd/CM4Z3aHWWnIPYcMNbZVm+S1z60F2rc7JvwIFu
JtCsNl6CeS9c3Wbr30URtJtSJ6AKgHv/dPhJJGpmndUjmpofATank1Kd9tte
aMoaZrQT7nvQIyMKLjL/pgVZL/flM+j0EAaP0nXjyMwF2m/uF86Xi08AwFp3
uVtGh95SlJmnPJau0w/u4PYdm+4ajlKDB6Nvg5pbjKfei3C4DRSXfKEURJMG
hsKd8iuQYCiRuviQ8Xdt07hHrHVxwJct8uu6IygmAMgDi7OaWhNrY7kh4Y3P
lyOgVXbngC3pB6PTJ+AW2yVaFuESCOnJTdWo4/qcNjEWHKwDQP7aqtbrmA2F
gf07EU55wRu/Xcg2YrBELYC6fsr3DdDwd7nxbwLjumemaVVdQpYWe0iYn1Xw
9T+uV++02MCJP1Wjjm/0ZgtKAs4Rh69IBfd6bma0ayMycXMr7UbQp5EYoG62
uxymEh74KhmwXBpZY2xNdHsQO28Yfl4uNggupiEVv+4LZZkn6gKl5mB+pj2m
amJMUfX5rvvsoziS4tV7lHocfyjSW9yBSnSZK4gl0++vHa7MUo+38ymMdgp+
Hd1azMYUpbaKxd7PK91xcwGNZKjq+wObGVhLBvHtius0XkFAzdoCopV95cb8
n/28NachZAlenwHs2flFEa9fDjMo9WBai7yTHrx03V5/sM58Xsx2GWLddiZ7
1qwIWoCEG0t55ujFZ93/OzMQQ4NVuWIngr9QIxNQOd0L/s8n+69imd3iumwd
anjhRt3RITKJDg/MFchF4q/IkrUq18KcBN65VeamwjIELror5LulyEzRIvzN
S532M4RnvwETx5VyayRSkBm+konOQ9knaalxr/KQptKFy1UMK8Use4NDfLlN
YdamOo0IdGmIJRYYcNcDn0I2LFrM/LQVET+m8c49/euDJmgQzFnLNHKFvHtk
nBXsHOpi7oQZmtNMISNSEqnJ+7GXWufmt07PEU8uxFeCDNBmSaVFB1HtYhVu
qXedj8ebmNPfyub6jAKwQbhscoqeEM8cekvHEA5jSHGoz/HUtdyxMYr75tN+
8LS6NtP+D4xx4l8QoxKGzJbHri9+QOkJtfv21dbpxyk6cIN+THJzJsG33maw
oAnfKDLnhxDuemcKAtlIjUaUMGkn7TU4DQpkJUsOMb5qrHtMHrbq96iQy1d/
FuyPv8EpYOZjL3koWk8zZ5J1jJtylqsxD3RRHUme5eF1GD+VVZYtefkvLnXm
/Ul0cAV/uyQXAeqBauqnLc9kT756ZoooEIEoCw7SHh9CaqK9jnywBE7674Nf
iThxeDi3WfLJY6I7S4UnHb6I5pjQ8M/leEiLDZNEInc35hSDOuhJ3Zj/cIbq
Bn+HI0+u9oxd8pPP/MyGK04MVfBFgVYrCa82yfeXUP1xcxfGoFJJ7UK1kIUT
/Z6m9f1DfsddsFGb8urGPn4jZkgbHL58ZFaoN/NnGPL4CGXqZnu9wEWTt23+
hZmgGmTGKMdbYGxyqUu46LTjQde//H1sNsON0ZCDjC6Bk+DCxpaYIAXjfZ1S
o0sQCMQ9NBbYX1HMEnyxxZSp9HDm9ZZuyYLgFk9EhSthlBKtC2tVHEVWdW2o
YTJrhKVyIe2I5gEbEZJIyHGTi7OMnjEUtxJPBhEGekf4UWeyuP/VeGm7k7QW
vgxsD8TmK7BfiisdClJwz1ouA3+yVRJPn4JRninW0elajljkUjVoj8iPCISm
CkbXSzKQy/7SgwBkdgtQV9Qo7ddxtrzyZgVcMy6/S9D2qtlcwfKe/dAMGEdF
Ukh0kEqfs4kOKmjuNSpc6CfDXCwfzyFaYKA1Ak4ymrJhYGNyRwyiB2x3bEzI
WwBBmhXA8CNhj7PblA9Sw0lRZq+ggeoSiO5A6RTlQWOSbv+vGrdiFygC+tJQ
ENbCKQtjubvX9Rqt5h7v4ReOY4Egs1b0sToVedJxykwXju0TEUGVY0tzcOR1
jQQSrue4mYDycNqwRQLiWQJuoXqEPSfTZ2cSUPoBe69Hsm8JHw/cHvI48Whe
n14eAcU4v2AITd+kTYSGJg4tjm7ubFucTJtY/sKKfD5C9nQwn8gsWu91DAJW
JfydXyYNHEUhU1ks7qtsOkO8lJBXQPBytkE5AEoVEH6iDAwiHM5p++jbZGK6
FZW3fnfY6Pz0GHEavT0hgIkTC7OeRM8XuLtWB35fUn/2AtDuk3HpNjjz/jZC
5UuCV9RiEjssfPn4x42/Hbd1uhvPXZc+nzWUHI2SDy74p1LCoXV2tbEmSUsu
M/WOPgy9UNxB/IC0WDX6IQiyD0okavZ7D3tStjloWfaP/q1YSabPNUIxiXux
6k0Ke+0rEZQLChY7q3Cfx62cW7Ayf78y89wlrznzJd7X5PTtu0NMtgBczoVg
FOW8f3xpwEKtPR1gAgCtDVl7M96fFtyh+bBE1b+4WMlY1BKvWztuNXyhXOU3
uLfSq23aUxkkyljt9Bpbwf6pIAQvqXmnUuB0NXM7v2meXqa6fwst3q/NS6sv
sBYofo5PrDbz/I7rBh2IS8Fi2q7wOsI29qESHE0st3CuKnEqN3p5ZKwN2+io
T12NkNcrjdHGvAh2Tonp5sGJdbtyohR+51KqMXjXxuop/oyMNeIgTD33mtTb
hsDMZCiEjT+Fk3XjRJZiUH3vnLDJagtkg7+jml3vy2qy2DZDnglEvzwO2jZa
w3GlDkwh6NMbRE8NvP4Bw1f6/11uKgq4z3vuVc/Dp2hnd1YTZYE3UdTlNhpD
rYsZOLnInm9c9WOebpKN8UUcPXQbrUuQS1tlNKk/aJsZvsPxIvOjDngLqQPj
8Jb1priCmte1Rcf3q5PcwN3eN9YXonvVXVWuLxP+JOukOU6uAW1W9NZ8vARy
sXwJRDe7Ls2ShLbtur4oOVjfpGmXZ3zDdOnYn+oyNxzaSVKAV3KyT+4b5787
ZrvLBP3KOkttI+1yzR3c7XuHrj4vuIKrE4TZWWYRnrkI6dvhm8Ih+/1Ng4+Q
lSSNOTyJIQbCQFti4eWx6MexvxPYkg8tg/MDKqg0lucdbLaqwilwGh2h668F
2wwC3UtsixWsE44Xddia0yUREmBJOTrO2xygRA1dqfr2SrBlnnTBVhLtACrV
AURuk1fX8JD1eMvQfxC8drRSHktaqXyaWvO+vb7FGhDd2+aMprLXHTaDWiRc
DuCzo6MuonfQkXjDPUI5yBWdkXKkxWYzXayGguZzSIJb0SGZBdJOoGGPS29+
XLMegFDFC+yv82zqScdTl9Uo1cATDmgtUQrop/cVOaH5YONHlmdEWDGEaYmx
LQ24+7tQWeUGcXzi+fkvH9WZXkEPfMqbIc+tei/KvPZzJhNZcbfnMojdVULy
zW8RCmhZjP4SrgOE9fd0aotonXcmlyaQdGivZ9LtLpnpw1VbAwk5piOnPUFz
AxHZiGLvpKTloc366Z5w1M7YRjtRJFq4TtCcVq9o87zCdMm/nyIJ+0c9ufUm
sSbfVDbuLHc+hxqOT7aGa6pZActolUCiYS/nB1+8aVs645e/2UBuomWvXZ6B
mJOH48PMnzdDRZciwDOQ7iJ0cpOtapUz4CBae0gtEGowBcwWN643x2VZX0CT
k1ABLIn++O+czdI/JougiPJ5hV3+fXnbOoti3HXUC3jJydDxi4Jkbz9CDRoq
4sX9TypeShFFoEfs0y9O0mhT4TWxVHnksca8KP8BLBmwCkQPce2TRn60hIMq
8v8OuNLfzy/QfhpdeB+4SW7fsLARLghpJd7J1dwQ+yoR9ZPQOuoeU0r3Dayc
IlEBHfDgfh41BlfP9SMPQZnA75939Vk1jIZxHbBIFNMjCbOeAVt4XflotzaW
Rv/nljUNJWOebvXtiSOm35RkjzDTqyYK3n9IxTynTFc4n0LQUxv0yEdq70yq
FmaoEf7rWZpTZOmyURWeUJKQVEwGoZJvPp6NmjUlLiuwNujqQAa0XzZMeFR/
PB06CiabliJk4S0X7llkxygvo9dnG05uG6j6BHapI5XTURH0Q3AznjF+FTnv
aC0qaGFUwMHyy3jaTbpbANo3lrWpBaXi3rSiYBKjafXqCdobro2hAADrCNjE
JENp72omGfjdZqDKL9jjXoQKXHMy9q/kCumg+qn9H1DB4Tnn6uHZoelp43IM
jF5A82cOoE7+W/VaIvLyYsoI07nCVo29P7i01ayrX1d3wQMIIm3XWOzVNNYk
I6RmwbrZJ1KUtcxmoZXq4DiPhpUTWJWSV4mgtIG4wplJrDcLomnLPE6Klfwa
JWHTtYgrvhEcTHL55q9/YCtJRhCSqtXni9wa1tnyATLXx+ZjHvUAIHRbwlpF
f/f6IFlaod2t4S+OHGr8zYLC2vrjlp3vTumLYquYF+PUuBmq+7lAy+JG69uA
k1TBrH4ZsIU2lvELG0XONTuag9I+aD1B8PY9oICmjc2KqMQ3WsNvMnNWrXhz
6wyWlDnGjawhkcp3GWeqZJLf3CyPetoolv+kqOwaakCO1ShIL4+nSkEFaztr
vo8AtEMCSf6+or98f5N7k3dX4jT0Z6AxgGrlk2U2FIdMnMCApusWUgyShg4+
8j/Yufgs3u6los0femSA5cgtzKrpRZEz2tr1QCI8aAGEOUI410M/Zq779TCW
lisBFLkR+hHUc2kXw9WBGQo9q63cGMWwCGT80YvPMpg84ITG6bC8yBJBj91F
8+RYD4pwYHnDacg9FSBsYPeyrYU2Y2u0HQH0Yl8e5JZf7n54DeTzvUP4GzCL
hiK6C5DgSdDGs55C315U15p+hWE+r9ALJiuR7qEzq8PcDorSGoFvh/vw5ZGw
BtP6pCxQQ89JmXaAS/VW8CKAfPtdYUrE5+Bjox6ns9XYgSEXWmZdmM2h0HRc
UxKfE0gHlmA4v76IEgQ0IJh/N39KZVpaQJa7SThvhmog6Iem75tqYdarkpF+
A+FzzpBXdevXr9MGFL+bElPDHKJPIyBn0rY7grFrr5WmtxxFnxDMv/fdSdJw
LwgFGHsXCb7HWa1FD7yrgpFMC6G8h9ZWQ0wZd55o2oh35Fe9uou0xP44OhHz
64KvremLJwf1QZeJBGiP2t753OWbEHkpflXJRv3ze58QOyzVGiApI5OT8lkx
0z+rcReoriKAKXXZK2hPd9bE6Ws4kBy5M3zCR31S8+g2KhGKAiK9NcvbQ0bC
LWb61PYYgSkgdcDYzuP8FDsNXyfGlSGyCdoFDdPOBUyvK9kp2CRfZiJ0XAhP
qSabyPsj9NF08yFZdErR0OyOfw5BZzLq8w4S3ahcgTzZ4ckc7+AhK17fcDD7
0o62EDTEkF7U8C5xV6rj2yXd7z9IPN5/T6xibmJEbkxRp5IikGvPtnAExBws
kgfOTF1b8H2ADWHqNVAUTflhs4JATUDoR0Cikvje4LfqsHasDZ0Ch7YLUvTJ
+qki3yRi3BWf0bS3OG2gXBWZccOqIQSRqPD0jKHOqNj/C/fSmko61cVOyHz3
Edtl+wW/Yi/1l2TOK9PwKFXONEjsr66drffPAyE+bgO5L3bG/hMrwCL2xEXL
kV4gIsEuwZ2Z3ommMygJtDqHIjv2j0q+L1gp8C/XyaTaIC/lmPMpogwoid/L
gaGo4ihx4j/7l0fKKZy6VWYFpONzN9rDPfFKh8AxjV1ujJw8JNUHlLLykn80
PrPLwKceaLCMBx09DqVKZGWV43hFSNKAyiwWsSbKIGAmOFD7NZeNy2a2Yzuu
F1U1QervC5Ht5WBdqb54Qg0bInj4ZbS809B+RTNSdH+eq7JXNqPtbM0ubIic
PEjO8bXFFfn8YesHLw1BQ4BnPvaj8S/oOq/MD7FzPFhbKi+XvZrdMDhy3rRz
zUhhnXlFmZ1mTIRrCYH5k72c+R8AwvKuOjZqaf8dufgNOF2tphCh4FpBmvpP
Tp0OxwrEDXwIAwWSslxyW521CUTZxw5TkWXyCC9wub/JA8G09znyg9N5IY2U
VcoLvXKNyTEM/JpCa3qcSl9ZWNKmFxwdF1Gv7P6lod/9ZydrxHwidFMJ62lZ
7sgEjqdAzOUwtrI2FAT42o9LeZOPCwTHFz6ZJ1InDiR7zbY9e/szcmlxXL5O
J0pjy+U5RPV3M/Yl8wkl+XX2hCVriyd7xmbqFFbkhlx7Art5HfpPhpw7CPJb
fe1MxCEE+jKYs6CROA0eULhaWEgnHMCHyy/zYABJlRNUTz+BO7LAq9kVuHee
x+4pgug14ejHmum684iVTAb1OXZkhC6S7M8TzQ35vvkdKksgFHVlPds1wP4l
gfqyEXWJ0rl3BV0w0gq3YV0y5aLBiKcFV/vREFjLv4CSr1wV9inkRAwZzs1s
AeLT/NCHcw/12Dq5umFP6mFS2lDC/KwbVFM5ouTNo+2XAzVwZCyYSutA5n8b
LnLQ73tfMtod0zunWcFEeSElDPPxjPqc4B9dN2Idr/CbbCBBReNzfHP5GSu9
doTvvzsQicsx0quRBbho+qfYIIy9gpSER5pSGdw9HJDUcOPfqGSwd7SYvby3
4ZypLaNQ/m+CL5ttawzZshS0bUX7IST5ddHPIoMO31hVr57voOmlBPa8MMPD
2qeyqOF+i6iZ+Yb7jx8kkgylIhwWsCB56E8HeVcMGoMEeRQQ8hQ+dNDK5wm7
5ITQUb3DRwQGCAGHmS2ZnzuqcmcBlVAo4fWfit9wPYhauSRN4mqnr8OfAPjE
m3dsomdZmG8zJVVYSspo6yB3Z+AnsmJ+G5pjwj7F2ri6m0jt81njpp2V2Uyw
5qlr86ei8eOXTSvTl/kT0/CL/8kE7SqrKJ2elbiEbSeKZr3zv+ccF2bWK3Dh
JtafQIq8wWLvR6GA/gI696SUD3GqoSMfxhF9UKCKJOP4Gfe7lYadhO6GZnJo
2np1Ur+TlV7jNz2aaj7sNSPNcG3dvazORRzgSxltPA/1WszD5udoU9T7hExX
YIDKVAt4Af8fA98MVjq5isu+Ifl+1s15ondeAjGtOS+WsrI4YrdqLyjAFXSU
Flsjpn7FTTV40Uu2FxB7ZJNO7H85z2srUFui1qt56xQCPpB3G2erroLzVGeA
LB1dK9XOXliFMgBWSV6mmJw1t5mz/pobUVS6h7Rln4qFGPi3Ab/7eVRG8OU5
VNzCEFbnAYulPQ1a0bqPGWvpIbFsY2gcBXh5MV9PswDaRYlDM3sjKWjwR7kv
cZBQfIcUc2ZKzkJ9yFJ23+pgUptmwqeJCSeqya7sm0674Mf1tYQfo3BJarRZ
Q3rA8HgbTa8YInM844GWZY/YOBHmIaFlh4AHLWCXskeJvkkOTHulXefIeKSf
1XdhmGTl+faL/O7uWtU4gAT/VA10ZvU9KzGsaRunHIcwgX4Qbu9/o82x52rP
3Cg5B5Vugaxd/TqrsWqBpzjw5tCdf5LP/4KNc0Fd6sFhOQJOR9oi76N7Xhgl
0L7P1FrjXmZ9y6F1OCresONa+1v6fGvwmavYlys9382HIT1Svz3ZsVPB4HHc
pfkf+dc7ZK8lwu6HCvtVd0p3KQp0cqVaqGrCmP0nThpt8Pexe8tJ3bTpz24n
EkCUtBKEtVcEaF8bgN8UOy3VXCDi7oEjy+C6/aHQzQ2mT/9rwAQy2kWs+Od4
l4+hx1EzNyNwZmMZOVBRCjf8S7RCBjw/Buowr4hxwybFWOUtkrFUWemkybMV
2ASx6YkdG45MgUBTMagki7nWkxSUUj0udtLMBGN4krFmuiY1o6CNlbj7Fx6/
QaT5Yc2lPQaJTA5FWeUnyuZ6o3r+8A2jf/qqZHrMXqEEAZGkHjkTcJ3h15cH
SFHe+wb23Nl21p1dI+Uie4bCQxvOZZcPFjuqEmJmfKC+4XjMjr7AhLLbEOE7
Vl8Ye9AFy+5FdbKPjH8rq3Z+82arRj6zz51UsXnVgM/BYaCledRcfRaNvru4
Mi96ukjTwijObPCpi2EDrv2rGGWM8NFWT8wqDHWtDQukxvLiN/gG00QZfHDp
rpAAWZa21gq9Tfux+WmhejWR0ghuT8DKz0yPrPVjNDG5/jpP2Asaet0UAN7h
xzaDz0X6Nfm+CQJe4F5p1eI/MeIKY2cjch8siFBgLgXaSvh5aqIZAykTyaLV
ri6kOOUVtzTvz0RkqnuPyN/rQp600vcZBISOva8L6fqNRbri3Qg0GVl+sM1f
QiuS3rpbaVv+AEuEhpWe9PlFWLwIcWck9+hHNKnHgb4g8hjlz8NoB0XzD9Du
oEj/ZTazDELPrK0KOyb4ra43xiKru6DbCD7Lg2AOxwHiK3pC6lljLsqrvicv
VmJhJilvl0dAxPHYIaTkJSLQ9CDwkYA08xP0xAQHa/vVZAGd88X9KiBBV1lZ
VOTfhpKRsjfbZZbQXeu17DEeEHr+/yujZfCc339UGo7wbIhE+tPDmxuoV98Z
4NNRbr3g24Y0jxTUWAqGPElX6IWkJSGDCV31MdQmNwgFXwnaEYuqfG0q8D5u
0Ld1PfAEEoeeyEa8FUh5J8fCq6GZrAWsMHRzIg+GjMFVogvTib4oMolPhB6X
r9LvoxCnWgvqDTqVw1Dl/Hkk/sc6teU8hpKwQwe4GNlduoSe52vDl0bUXcQP
Jry9KHVP34PZUIJJ+g+f8SyXPGFQY0/t13s4bGj0my3tePyPtHzdsb4M8a5q
zItRrNJZ8/p55cvfzqenIacbNkESjS/HA2X31bLsfvA1A92oOCsGaHAIXFol
0poF8VfGMmKcoMHhlkiqNckKmQBeQUOCUFNKoQY0GrDHs4bzCBGjYMgoK4qn
JqhOjEUJCh0sDkASFvTB1VaplGzberkJuQdqamkKxiRACtbkc/MGtqLCYbAi
PSpTqKSUn/F/j6fSNwgfTnDOGRyFQEbcU0k4hl2iYHz95mEg+OhYPeFO5QUX
pmNfPAp2/38zEseBeXrg1Ru+KQL8JVO2qDgRiV31Vefug+z5hZG4Y6uWy7hc
zJY28PlRzC6cPWEKekgDdheSg8ThU0ADbFDYbAF1N9I6SPFlTvN69bcP8sTJ
/6+hgvBXx57GN8FiDFvv1MqquvV40UhSoT9qrAW0I13g80cD1Zh3DLkx3vLu
6XLy1krXUpMIMaeOWrazljpxFpg8I1vvEs4IfxFDzu50JgwmRkBT3S1/HOeq
2vi1+b0OatyS3vNYxR2qtpHHklwQmfluFqh6msoGI9l5Gs99ZLgGYQLzrujx
T7jBeD7ex8wHIJQpm1bOGAPW5BXrTBUJkYaBcfl8WhDiNYxPaXAmfEk2A/C6
+5YXZS8lqLqn9DVNd2vuvCDi6LaiexlULxZhKUdkIBw/24fFxYsfkfOiG5WE
qPpyYvYW+i4GAp8ipTkIX2Iwv7lJyH+Mr1JA596Px140q5oENuOIYowNY36p
YcvgMvSEFUVKi6eQeGCy7Rbs9WYVEeqt4S4B7XlOmv7uq1y12MZhH29swmuR
Ski+EgzDmMgfvjZ44iWevZJDZ4BZxwGgJ7jgpkLPKKL82ZpKDZYu+edHE71M
QjSBnCo4prqMfjSdJpi717JYEJijf25GqHVKOaKHTJE+wqhVpjH9YZnxZFvP
MendCnzWuW8KmDDkKJN/9crSBkOaN2txTxz0amdWLEl7bT4Uqx0IsxWeNOid
NwQHV6GoQkueSwWQMmEoVR5dfhriLydTNtYcMq3McwtMPDoGzAN+ATqrn2X7
9U6nBEF4Shlm0omdEjyEIb3CFG1TFZtclI3oFR9d5oYN5HwgyEZretzyx4xk
o7GDeOIyqy6/aHY5CNUlbTuE7BR2X4UfYGoxqMH14iBZnOphahYez1gptbca
03bplvBORkfmypDwUbXedeKu3zilJAG1YjkjpPkOXSRajWYEx/1wZ56Gxm2R
3/zk9ZTYB184t8KdJe817mAYqg9HYKdau+S7yHQ1VZAczG53cbkq/Qztt5Hp
CU6+cBGRouo8IdJy9YqDuMwjBm+l2BZHzBME6n+l7UJawcGoV2FMD7rcPtv+
Qje9TE6dWYJ8NRb/ijhNW+4fSa9QbVvI0wpGnjq214gDckrSH0vny2bayJ7N
6dNNeKoS4+QhjtJ92VajsMi7x3Vjo35vQ8J3I8+33NeQPKwSgIykpRJ6ykgr
UXbkx92WOIiKkle+J8a79K2HQwgtRm1EJJRgIN9wTI5UJ308JGOg/bhpm0AW
hDHScUhWonY2HDEnArp3iIKPGKt/vv2G5ETXpDKxd5YWcGdnJvv0P+uDR2XR
t4xhkH4Ozk7++Ho3ZiyFlVBxzyrvYcIURYEcBAeHK7KdHhyzOj/HfZqZOtww
YoX6c62A3Vxd2UsdfhJrYlaMnKidZhqJfjz0Crb5mYZmc1zcuTiaW6TMz6kc
VsANNre3azpPRL0PT9en1YzvxPAhbhNb7uz1zes/cW9uRe2L3cIM4RKPNXse
HySBhiBKOjqG/6xlRIbvXUEL39DCSOS9D9ZM2V1pPiIBswScbHZvxxnTNTK3
qK5GorGAwRaogN3Vbrhg1ptlHV5zUbAKO0EZtAKktDsxm/Hud5bZOcWSXhVb
pKK71xN9Hv5FTix6H0hAsvB3FIHOgsUOrRNmVLyPo0733Tt0WvNIlj7LyAc2
PTGiA3MgIFzRYvYfigryi7WQTFGmYlp+BgQHDbfdy9nuls1A/RxjI9hkMByC
bEhXZoFmJLeRWdc44dijWDomkafFzhe2FW8Ns/YSqCiBxEGNX6D3n/8fRvpc
U0l5YmS2A1A37G4ut0+DZo4377/wCbbevQD1WG06k65sy9Sdhd5mRAmT46wc
hJ+NvEb3Qdgxt3kJpyAeZ1eCYiz5c+buWUfqRlU6PqF8YTqcCgrb/4mH6m09
ZhcpbOQu/CuVGHTwR54VzkOFBANu54+HHVUdcagL7WHgxnGvXzUQtwOmJFiJ
cJeM1AcqkypkRFWtewiGCfQDAaE2yQK5C2p2wv/zcoI1WjZlxsRVl8L318W4
zQMhMzuQVAJMQp4T3Sqgx/SUDIXRkJjOZVSUwNgVUNyG8gmv2XEV51RApjIQ
jb1XhnQlsvYVqlkYP+vbmwDfsFCGwkjqrsgSEe4846gkXtsBG54yqkGGJpSu
+Zn+uA7uYEOVjxthGY3KLfbMe8B7Yo56q5hiQkt/uWQk2xUEflpk/VCDcQiz
IGypuneHwj//WNr0Ztb0HV8RDmsnZnCDDDHkfszWtMWmLuCC5zRRFqQNoDQQ
D2pN4MYHBYhB3k9E8AAE71xDhinuXlAReJHH7SO44RX0C3VTg9Dd0tzsabpv
VaWAtxKjIlVYavKIP5MT7BNn5nRMreW9WidTydwEhZB1deT/NjQ090lkovpH
FLhoMDSbQzNWLmVwXj2Syt9XQ4Xylq6Sm7OCwsa2mu2jFboV7XKCXS/7tYP7
nidZ4b2tB6x1AYjRPsuBexy/jrVP9gzL4tD59wWvBn/Z8Of8JE59tirsQJEg
6v77U917bJttIyB1SPF2NRJgCQfLkzlHk1zYnrBMntiLrGJsx0MW9rrfPqVB
MNwhVrEj+I3MI/69OA647kmwm8A3OaevdBzGehiKjVrUCPEWi/ujOUnw0QDe
f3ly0JSK8Ytl+8XNa2jvUC/mwiHM9/d5nrPsRBKfbiiMydvHcGABWBCdZEWa
hm14fz4B8wG1xl3zzIxem4fD+p/38JztsE6VrcaLF8ifOhFwuFOBEy4nZTF/
57RHM8hgwfhzYKOuDnTVIkRMUjmxsPfUg5piaLCcv20XEzbt+sPB0+goro6h
hNkKdlonh2N04zclAsExMoSVn1zPBf4OwBxnBOGI+G003mN+TpAKAgLRoVVJ
8XxeF8FOxzGWsQJ8KZXDogdV+BI23Zy0n4ZI4256QgsPpy3eajh7DdAQTTwr
N3VX6MnAuldcr8O359JEzJcr+8uytqXJIni4sXdz5fbw94NVyTA57u/xSgRT
bZlvHGaclRkG0NelZ95MkFj0PTvTxTNnc8ZcxmNtFyXJGw18bIR9ac7guxzF
AhIxi18LY6H6P6AIPtGn71kj0ZrtnqI0S11x9gTiwqdwXARQdGOlUvVUZwtA
9sRH3/XYZT3Djq4xR36Og8v/kUqydlaAyd8xBrgNpJMQMcjA9z5SwnnH01K1
EnX9c5a6r5yMJzOWjWIO353UrqRBAz2rtGzvgQTiSyrYaNJJ9SRpnTiO+x7c
9ZueOC4lSTUyNKTV4aGsj+yUzxo6kCgLi8kSxPzXJA83LDGnHNmLJnicFotX
4HJWHlKc1KuNDWU8RKPwpiJOO6sCD1/IYN08TU8Lih/PNQ8Kz+gBmXmWKt7D
uA9ShGyckGxaA4tcpavET4kBJzv0VhG9ohJz0b2kVYdnu4mmjqvF82ryMvv/
gaeJqOrVz2Pavd6XFhX5nse+D7MUcxltw+esZ/Tvg7ji9uuwikFwb1PohebE
V0sbByR2WFz98R1lsrrg7KgAVXKLfMpw/3Chf/4lidzh35kjzsfVx29K9kW3
j1l6k38Ufpoftk8CbvQNvAhPBFpcB6I6HODZ5zNDIbC50T/5v7FR3V8tc7qk
hbZpO5OFrTitqAA3CdgML972zuFeyp62Esb5H7GGJRShMYyZtlCpPcfhpBBv
vZ8iBIh0gKdjrERgroyik5l+EnyI3QWSN/8fcf2rCkcArFNhrzgEzzIUu0fT
F/3xF8uqGTJGofThtjwn7spVD2ZDBkHuxilX/LMhDUJpiGhU0Ft/OShP/Ufz
mMe4udg6ySmb1Xzs4SmsqfKY00hhb+YRJCLVuAgLJYkAav991Dao9Oj0KcPa
/dW3hc5G6JDvx2zbFVUXVrmcaCwMbW+NnHVwfsjmo10IKMVRQF3/1ds6EPfb
Nr5bJHLZzYMwCdmIABQS4JYTegMCiFHCwudY6DhpN862TCd7SZckBy9o1x23
VAlrutflMdVN8g0kWuEqeh3Pig3IPIDeGZgJ/OZFNQImLAxLGZPFR9uo12W/
PPLwNsx2CXiNCeMr2n5bQe2yN8ZnzlXZpWgdBJAHzsFgEKr/heRNA0b6d3FD
qrSe4nqVdYYFIf2U/O++mAvkmVg1zjg5P8+u6+xNjmKUHWfxm02SS5Vz0IL6
tOekDUE8PE6bXhDtY8njMa84AKi+/5/JOgmYiH9FIvvEZKQ44CqxFB7q7GWB
auDTxi4CaFQhdbBrmndTF7a1QZffyJea9Ff9CC86BbSx68tAN0XzpiiXKorT
Qb2UUh36MNRHlZ8qtIY7V+MBq4W9/AEMmDc+/4pIJD2/n4aMkhEbn/o6m4zd
L8MknFTowoZPCtHgFPuUJiLqKlrJ/A+T5tK/+AifU1J2WUjYRg7FU8Zsp2Vh
HWTOz88PTXvmmfqVkauP+rUWm/ljF+PbI8sVJ/rpQHWHNK2HV7Byq/9PrD0y
b/ZamV63lPQ9CeyWL3n6cBIzTRa483fAdh4y0ig/WOD3W7vQW8UlFRyKsUyS
DysuDOmyvdP+66bMY8JNYs8uQJx+2L+xmbdl4zfILdiPDQnFEppFuna50dLT
iS49PUj7oXjrnh+wOa/OqU488EU/iFEHww1dvO73zzzVVuq0OSGbRg0O5FYc
5ntb8F3LGUMwH6fFBcoOQM2++5kjyyMwz3x8C/Qxumar0Mb/gDT5Ig+opB3H
3/cbqyO4UN66h//Pe5k5CYUfZFbh2L8lt4dZQ1bIIEcEcdcGFSLvXEMGqdOn
AitTsRrXKKi0YyuPjBOpAf7DU6onmyyLVlqaGRznu8kDiOzGJdSzCTzgSZVI
1VfPvK7LLiP1H+bONryEzu8FW2MC+wrpZCSdzKhunDqXBoMsa35HjRhTD3yN
24wBXcNyu6SmqBwyZA7LLEvAmeWzUfTdlryolEwLF+pYj8kHtKZXLnCX/Ov5
1S0DrY4J8YF2X5txYEaXI/jBCxcigTU81en4CRcpG+ffyGgtatfHwzAOaci7
ZoTv9rPa26IB/+vA/nMoYrvfFZYcl1Nlz7iGT06Ldis3Tc3j3SuB+0Gmmz19
4PYz/YUNMaRufii9jXZYaCLSqF2/7OyAIO4XlRilmD80trMTPVI9vHfwqq1N
oF2WECuy5kLF4CJhV2g1+NP3LUxa7lHa43Fkoop6v0tnTIRrhLT9bgCW7tT8
vDSSX3+8krYoIz6TqgTLPctGtp2tzP1PlBpdwwfqUMVt45HLxD85sJcrbCQe
rCJxUtTCPYlUtj81i6+GKIysX8C/yqRATAkkxlAg3XoMGErc7E3guYl/sEdP
+j0/KbgylxCPqhnYKEUNxy0nLkKVz7Q5mFRGxNXBa/TCeg0/tRIkZ5OmpqPa
Koh2zWXEO08JdlnvzmialAZoz5ToG90GtUaKewGVfqk8RwtGrWpDj0jEqp9G
UC5H6Hv9zJ6yxXGLUmJVQyrhKX8kSVkvHhohV/2Ot/BGFELPNoKtykjVIoe9
JHiWg8yUPACFPYMG+CNRQAiQ91V8UyQSeYl4NCOOv1/vE2J7DF3ceoLsGZ32
xVsFnTwb/Y0Rj3rMPgu4VBBypoGJ+GYDkuo51iOHSm/EUp4xG7aGN7IYjjpI
Cw9hZ1N5ZdX+/g6an7CJw4ZfWjLZDcgrPoW5gThW1dPOUy8kV9uhbGtjihgn
l41Wg4csyygnzVETVo1f8RvWsyX83ZSzdG+TasJVVqb/9QDdUumCjot084LZ
HZsaugfqxWAko2pYPFGYugt5MuIAgx6fED81palZvm1AA3hcZA+737eipoUp
Xk+k6clm8/yz+PsCpV7cRGxNGIrgSKZ62MeXEcBkOqhn8XflX/x3IX44Inbw
SP5Ezye6A6UjXIVa72eMS5ZU2tVZCTaV3tv96Ty1glJ0dgZCj+IRXVtkp/Zr
pd23RuMzPVVnwK0vIfc/03+jZuqICjmYo7ndaURHZzsBfV+Ekh+N05VvhNSn
dNsBnEPPk7nsd6y/NnItU/lV/uj9RsVhz+1ZHX37YkxrmRbZA2/lmufgqZHH
HZEfszirKzAw3zTT5mdHy2j3hg4HKHgmHPwpvWGuTxfd2H2KNEEvGYxq0nVF
UmP47u6hPHg/v8TEKHnmF2ndlrulQrNptjdYOtPQ6W6bh+NQuVUqPfcwgfRT
z1tIucQNg3xymsJz1l4Mmv5en2BJ3Xu8oHxMWO/Vo9lyki2TNX8kX8LNSm0r
t3eWyc9CD3YPDg/25EMqNjfC5XwvCVA5PM0eGatC8zxfHC2q5JGXQA4eBhBM
ssBH+iy+L9HN1aUw1h2YbPbutkk2qBsqlt2qDUHkNIxYgzUdu+FbNg23Gduw
QiXBFHoq803BbhaIBu6vmgogYFH/aROPgbSvloj9d8b9PBUqKB+WX9etsscl
zYEOD7Z4i1dKMFpmE3KSw3vZoqcXJxj1sYads4x84c0QsFMT/O/SAj5daGE6
/L1wiLub16AM/8cshlUvffjwrH2Z24SbSRw7AOjtG8rlIXBXNyDCKIhkRZxN
130St9Z1Mba0BQZCUpXJ1MUeBo4GMEWJ35/g7dQDFGiSUTx+LIz4mIFixyn7
T/f+G4W7+Sb4VlZHoMA7cSY+ugMOk+KAACrxs5IB2BC6S23vgGdGrzDx7FrG
BZ4LkhnPRtcWswNuwKVf0dYvarjO6pAg6iQWFbsLFScQmZytvwbOvsCMKWaQ
R57GRaZ+KtQEwvc58GJoGot2cnoZ/gYvuv90swbiz8FHRA5VC3Fojd+Mauuh
wDn+Eid/pOrzH4+OVR3N/RPiBgUGA+mftH9XA77kDa583ifQJ/XLWPDU6Eqx
4e567U0ZCnLiNXF7Jd93aWvDQ3if5FqdDW4sgofMla6/dQVY4CerfEKENJyP
KtV6+aBGwpDg2IT3zeFaTzzf9qgYyPzNe3sLHCGk04kZkkwwLdTfa9VAeXkI
FboEalqxmzNW1tbLAQT5SuF9li2Ia1vfpHfiii30ILpmIpdD4h1qfRDTjz/3
9+zecChCZekoJa65PiCOo38rNjLLvIHb09u5ag/ZwKTDTbbFdFPKbV3JXFCR
Z3Q/rFJzILX0fa+uT4Rnn3NVZSv62b6cBi3ehMD+I/r+aYAo1/mp6ewVb2xm
/QczI0QQenP9ShZwqSuImESsXL8aFqhpDX+jV0zBxY3bN5+Ufc0jKxLTLjE+
KjWKRFvG78teguttcgsuQTedHOBhFvvCdtcdniVaJStbgdfDxaPoHIDTtBUJ
Zd1dAKcM4NaWWI2aMZpstHNAuXdax+zGYEvMQ3iFDCXc5PhQBDdq/hr2RyLC
5Q3Tc7S5J/GDxfjuTGkwWHnaGn8X5j0ojsTRYtQMC0wo/brpvOhZGLI1yPD9
Mb68SSkGvNzmLPunSejvvl3zNFezFfm9ck6pLQt+zdymibDYKPvTMozrWBso
0zjRc0cHiTKyyW5dYvG12vC/XkLVQJNF/0EA5bveBurdTWdZ7Qhm3F2yltXZ
otvbgzGJTldbPO23xYhym/3VyL6B6JuXpnZSUD/8PbnTAIfi7FOn+zE9Bbpi
VMWYCDQJfq1E7FsJmuJscxu/E9Lgh1WGvfchk36SoDL7iO6RFf5CeyRH3iDU
aSiGSVPA46F76x8Z/YIRyuGRYdrOIQcJ/dpmX/DTsqhYsKrSnt2Dppv9yC9p
zig4didx4Lc9LGmf5gJi0lqN36lr0k7RKV6+XXM7cxxV/B5IK/wKOrmHxi9J
VJ58I3J0HRL15ZYCuw7FH2mNXf3qTFL3AviZB5wbwceZCPGYg85qZeOv7bMG
5YD6FaQX/pop1vnjqBtqfqcaaKKtpACsR/28tA/REdLxIYfdG9Mg4tCuWPvB
Cis2wgSkq6EfPAOA5BBtDciKYhruSkYElPMGQe93pqSXDg34jFWrQUBxHMO/
n5FALUwXMBIGB4vNvW7AtMWiW00cFf4cegrM4zzpRnipMC39XSn+3e+HIa7s
lL/0Fy+OFSwNA9oZn86f5hCScwSBCOp0J/MimUvF3r7KBS/1MQJXcK0K1Uz7
Ubh/WFwLHzNRm3TJRkoLsYU55wkF/Soq4mBEDeyYY01YHupymIZ0OkcQxVpE
KE/k5KQ5aaNtOYjiO5DJgVcdbBbJontdk0rYe29B7/QgHSO1BUHZPWbuuuly
e9fDUhBby4SWR5iO8oFAFnkQ3GY8PFd9gVfd56A797UrlQFehjmDS/MbogoP
1EK1GEP6lJehAZQXLumhv+VN0DBrx4R/wKK8Yl8iQf+gdcz/rK8V+1lWC0sK
tD146R6/tBGfQbW7SLXxl3TGuVBMVgKssb27QoVfWbd0h6+/bTk546hqjTjV
ncSVFxgJyNelPSSveyZjCtRcmbwQcaU7toEoKKkvuYKatQAjUZIz9sx4GSV8
5AtIoHmO805j0cxItMpHIPa3BG6Llmh3+dROWMR6YzmPYMrl8E/FGOcVlngV
VCOoqKxI01Dq+G+AqzhcuHzxGibrqOuO2t0iRSH72qqpJEdwZChVCaed5F5C
tmvbwH/Tp/hqTftiBeN44VK0DYM9EJTDVwB1NonX1IlS7bwFQjHrzZsmLHy6
10RG+RoYRCiiOpcq6mVXXMBU/6syT1oD4zDQbj7gjgobmpxcXrjqnWH+Ef0K
QPVRoB1MbrNXyu8HFKK0f+eyqw6f8O22RlfEFTvCWoL3B5rHIZWeL4nOOeJ1
+bs9a5NEl//PlaaJL6trd2k7JhLbKuDWABKAEBNU52oYMIGxna9YJulFEorj
OmXRUWcxG+InZf/dUINRipXTt2rtBBBfiDcnMl2CdqsDGiSC6jU2CboO5/uu
fuydN8HJ7JsYbK6NWtIxVe+GCrkaE+Aa+4TDPSfEZN5tRhiRVhqJzi5zh/qz
ZmvC7x2eFBK+EWdl0HZKY65R/lDmfIoOOqec8RgfNeOCbiXrbmvzQLukIZp4
crj65fKx93SEJQws6M+pQMKkrKVFTNdTIriP0myzWowUk5AiMIN1KREZmxrn
q8YHM6PEy5nlNxmNrBCxjp9j8ofQppjEV/tLIZwzbFaS8Bur45q7RMbsayCX
SN5xEXWfMdIDQPG19r0hGMbSgGV7NqcX3O6dDF7RcISqCdq8tJRMgWqThm1E
4iutviloUxoT1C+p2g4bQK+W1XZ3cUmHdaihLTWPKKff4RGik4o5Cw4pYhzD
B/Ka3uVgKh8IDyovtpUL6tlJa0o5iDYgdi9x/sc5p4VWzi5qHKnKqWqKQDkF
sojlRp7GgIDgBcC8da2nF4MUPO2fkuWG/lcYQsNxe3OHPEmtSyxPLLKuzIwC
jY8b/p5cc2EfJjQoht8SaO7b10+sqkqWSA8El565G9osKGG5nuZTJLc8PsWb
89uXSHZk4Ir9cl9xMpFii0EnYEJo4fPpUc3Ug89O+o7l3GSK6muSvWK+MfpN
BFGqH88BlNpotjBOw2pnecDR8dlrUBWz/ewAZ7rw9sHm1YT0F7yKA2kimcYr
Xg1BKFWI6uZiu4QIBWdhkl/Nnhd5cE5ooVEV6qRi0u7/Vy5y+vFdGaSvxJOG
OL0RVZ78EMgGeK18P3XJnvs1i8ol79jSmNqj9Jr6uTs+prQo+dZ0/yEqO00p
4+8X3pRZpNE7Dt+Ipayj7I7fbXAPodcEOYEifDHoLWQ1l5s07WeH6uCaSqh4
AyuXxIr7+mU+X6MRve7tyccjGe5crliUgz6UH+7ezvb+ho+GUJl1dAdlT5IO
VJSsmm4X0ZeWsTqW1iAXO+GWF4dCk/0iofO0/jhbApCcEyqKubuxpq30k4kX
YcYXc/Bg2XFNtR0xvPV+VJtQU0OjqHN42ik8Uj25PipgjRT+YjlS3NCnWC27
zPj3dZoZOkawWQmblaS3tb6mAKZeteJIx0iuCHXL+kAQxs49F4reAFQVBdwn
KEpi6aKNIs1M2aJl+LeOoNFT8R0hLsrhB2Sre3StmaOx6aFxynnL5agEaGWq
VqGWQXjdrjXibGViLHVMm5GPa0q0BtvMWK2tNEak6DaywJWr4gxcv4jkCPBv
FKuRcNzP5n5FaMk3birZpUIVyBhoxRSB5U7OqP4t4Yz6V9ywxdBT2QoocgmN
+4Ez74YeO+8N0OOT1LlZS/ufaSm3YdO1HYVTzXWPI7KcEOq1dTSPVVkeDRmK
zElHBohGdAG+x77IrDhLm73fIqtWHGJUXgMHEWd60gNCjyENrmmoXJX8pqNs
BnAoAYQBu5TFKAkOZt8KDj045VtyAZkUbb0JNzFlxGtw8nw0D1AXo9mpFoks
MCTAuGvNwit8qhUVKlZS1uT0e6ddAaGx0Ny1UeGlLPZM22Cxr8m8c2CgSK8i
OADF27/gB8vEMGYXqDrWE9yJHzp8z8KVH3Wy13FWzZDnoUuvhk+W/MsdySqs
Sbg9CY8BCXhb7vau33nSrZu9Q62lcAQeE7zlFKxlz0IOynA0Wm3+qNjeFL3z
pSkJn8PrmEOAKTHDZA6QUSOdIA9UIIxxYNKww2LyMt6wSDig8oyTdCGhSXoO
i+Y4h1vwruyGaKm0ILT/6v0Pn3Wlvr91Gw0URp5czkCdKmFBR3MM2hCNYMhT
LA2lNuD4PjhDDH1yC3RzZeqUnVsc/A9kZnWQF/kTydExpZGpUdOsqk/JZX65
N6bdqhsfXxh3iuKj3+nFnBRI9jel0ljl3neAdqB4C4RXzrYxKJcycSymekQI
4Khm43S5CNgV8Coy6dxAlh1d1x5CckHxdDE3aAnNY4na3YV7eq9wAsrCysqu
uCJLZCwVTlWargurce4Z0hGJrh4GhF2iqWgO2GQaf+lYQY5qUURW6iqJIra1
5iRgjrXPeTjH51J8jnTC8SLNSUI1Qe+uFZ+gRu7fnOAGPgRhjYxVOpDBE4b0
JHs7Us+evQvUd47RnCgltizwue0/bcR0xX76N+NSc1I/7GPgQ3IltZTr3Vtc
YZTTMZkiOlim3BGT1csxaWSZeB/xGbvgcF0xECed2gP3DbnBgckePDI/fjQ4
eKc10PWn8fd9dl/XxBmXBmvyD+wvWHNWFfmlDNJhhaivbqHksL5WzbOpxBUO
YSOLS9OY/O8FU9COQgIivEDQPXxifnm3obiywGGDHDBSHOiCSl5K/u1oevmz
6Se2LTUc/wi6aEz9sKPK+fLgE5ulzxLH2vAX/Fgv391u5ACAa78hx32XeS3u
31Pb/m0oJBpp+NZPKIeLAca8x4v8FWqKufyFwLAoQf+M93dptsYGF4jOwOdk
nczfgPxjRjE8Eg/XWJNrPsPZZVhpBytVwnuKanDyZiiJFWfSj+/EF7byYrmZ
UKoobBTFap6NCcxkSelb5aMyZK+GuD0PYBgUrFFOL6Gzsv7dLNg98t6anEom
RN7H+tIgZ18PCooRidLzpekVPMyozBwuTE5fp75YAQsxSukqhFy2WZE2Tzx7
ulKjN6BqHU3c0JkuEyqTycf23GaEjFhveRPg/nkbHFiag/b6lDObZImRe/VA
vCCSANeaqknGGr7PjaDu1EqnfuYmBp7cbXNzWwBfsUBW6eLzDdV4dpeY2sea
k4OfgY6ZYqwBHty2jsqm+aZ3TJHY1GGW86D/9VMuCS3Qjshw9eGucJeYloBK
0MhsOf2niaUJFVQh3GWatCEfuMPs+lgcjnV1FXVK4R252x7vG10q0MxKyS7C
2Nx5PB3932DCy7NzJkwsf08iuw0BN9oAFJRCThDfQgHegloos641CpAYHpAM
O7cgklWln//i3gz1sv6mwgKrDwAYTXeSPfR4LQKHDrTkJYb2wwLaeMAJf4NE
Y0Pr1FvGgsCVuEq0TY00VZBiwISb67N+eTwL9g0tWtE1+rs8zYAOzzgzgE/D
/g68dqcfeBaYfaUPfcss6DPVxwtvXZF6Hhv+IL53pmNO9Y/l74uhlDCpWfrC
PPQzR7bXicBO5nFUFqqrebF2o5d4WrZlbeG3soDc1fCOq1C5X8j7XURSI0Ve
HvJHZ798PTmaoCawTemUHQumhJo9f2cT33XBXmqqc7NgulKy8chhBneAr/OU
Q9CTtoWbUYTPmyD3SyB1PTlEsfE8Wy8Hzlqdsk5fr+EBY8GBflSPPUlU4qgA
20qHZiA2oisn1e77nFjJhGW09SVmgBndmxX+cmLkbaCdcg+xEF2TVa+Wyqy7
737TwtVOHZ8IYjzCpaNWZrMEtYihbMvP6QD1a6L8NYjRJOoXtwLy01ENAkFv
wnS1BQmZTrDuZ0Uk2wzO+uO0YQwItaOqtwooo2zQlfciafytuzjOAcu96wQd
01iUJnY++nk4ifP4L3kN6EkNiC/drWJiu/TTdjDRjJ/Ffttki3xj/YyITyVB
drEzaheWbP4bO10+briV0y7uefG11H7idu6NfHMeW/12NMfNDtk+KLD2UtPW
r8/5UTcxFDMtSPK4IW2jiGbyrSk1grylApo/MXZJL1dd5DEx99oEbm0a+lyj
UBH8VjLvEA5IF5q3rD+gGQrthkoVhvJVe42zWLnc0/Mm5TAnk5CNUFyLfbdT
K3RW1NN6hDuq7Q3bV4SDVzf7K3bOG5osWqwK3nBW/c0gR1JoKitAE8hIN2MF
UA/FelN+ZPV+MAv9/mISsXCNM5W5jjpFCx/A9X2TVDXTwG20T3bD5nlUwZNt
qaWwDWXcjuSLmYg/xNyrrubwJrAsa6jOYILXg5L7DBUaIEAFPuYgZ9yOmov6
RDiLjgGa7RQEQwxPWegwBFyLAHSE8GYatp2ByOAKoSi2sblGSAR6A8by+7qh
WGsywU9yCAuUEC3+CzKstuw2qDW9B3y9HzUSvyJoYIQA9sx8UHS9k8iZdAVZ
0YnfE7QuZunH8ulkeK0OrnvL4zlNRe4jkzdDzbll5YE3O2Mls/5QqIa75gQy
vh9Xs9ZAZ2RRIr6MyqqLMx5MOTQ4VOHzKwZ/O8M0rY/uEH0rDqV5v5H6bzOV
ZS7L2tFVXgG/VLTI6N2uOqZT+HK9S5/d9qZgBeIyC5zFjZGIggdeRg7HS1Rx
xre6InJlooPJ99GVzdWnnI5yQV2rRkuyHHkjHAHYtFso2p7UVlmcetJtbVhN
VaakWv1kq+SLNFhaZv0o+/DcOy9rxXw6HQ5seCfn5kwfkePK7W6BVeny4usr
6ZD+vezvOaAlBOywZkf9RCh20SCH1hLd/7ZxAWtM2YdMtw6C+9TWHlAwYOOb
B5uRyN6ti/PEclofTSBa2fUFS5BqCXpG6XoIGnEL2ZRWJH7+zBEWfX4MdA7Z
82feZM+obqjvLC0hN0T7igu23uFePD2GWjANJiS7S1oF9ivrhY5qa31V4i5Y
jhAyFbEGcohsENqzgNCIz38A2IXalFG9fp9oTghwwqslBr4WcW5jC0+azJFW
FcP3y2WjxmHNCmlNuZ5ivQKQmTM+TV1+BfrznP8O8lPhfFhcsBH2CBQMT90q
BMMcwI18ejlbJOVBhI9B2pmo3v0aIK98Tc0feO5mtAVeaDyImL1JLq0iaIv/
5AolRM2ENyBS9q+QdRLLIgCym++RR63dO2C5X+D7BbMjnOOsSEpwh5KK3itN
wfF5oK+bjXpoMANwmksCHsHoILCz0QBLj6ht1Hd6jft71Iy+w2m6jEuVmqdn
LZnfJIADwdrQTrYqtlBqsRIEsSnuJ7dTJ5g/OAXpCUOY4ydnJw1Eew/IMJHN
8yDeG9Km15ouMTYRbBQjwRO0Hb9e1iJGrxXe0Fuh+B5wmgFmmn3BSQ+W4LXL
nE67nPIO5wx0Bwip6fwwZgK7CBLsZbIO5KbcZ7uK6G2fV+zrENQOiwx1g+h0
kAYYWFmSxZKfXAGiqeXmpAp9wBCnBGTEjQmRM2mSo2c6bvL6SZafXdIzMkOD
qmhL63wpsw35MlLMylQA3Et7zLkMEXT0uuxz+cLPR0sM5o3X2m3Jav51dboE
fTCRr6xmaFxWt4x6FTn0Y/Q8FjTVBlsYXwdFJc9lBkulESFo7yWSUVE6hbBE
EQ6q3ng9aW+iT5tOD7TdLN+M34k+tcvvTfsB8rzwHed8OfUpHEHYoE/RIHNm
8F/uJBOLQyAqpVwkDBDTlXxXCkVX4Ffa59/ASjydE1CdMWC9oEws4vdpmIX1
AAfXglAoPO4597ML01Yh2eBMb4xuCXXE1PaDW61RQ4SA5GQAs6qxyZFqRZtQ
1bsem7C8gIAO/Pn2uTXrsJ9XAUlC2HBQa8TrSIO3/SfJMj92IiRUqcRfTQZx
6WREGUalw4OqLvRwtIaNNOKbEEgB2+Z8ZRZIMWxfTYshLBteLH4jC00snaxx
wU7c6ywMUgQM67QateiKCVGsBCOkDwGz1QjXkf08R3yZYHCZ4fCgR3D4cCLG
Uoir6d4R9uVOAtpZSS2yaM2JWngsZAAcoWKmg1i9tvaCt8gwDfFA2ahrfLQH
zjy25T/1L8U/qpHSXiXxUjR1W3cq3caVqlL64wFLcHlHZKthnXcPUOCxKjor
+E4lEAmJ6V48GPrz8diBQcw1lLKpZGv5E4ljD1WvEz1i7/mjb4hewhSpItSG
ZiROnDZg0qeUcGufF6e6u/Ttx3NF/fpag5maeJ/fZzaPj/Phv2Dl9Hw5yHr5
gXOeBZ4xCV5kmLI8eOKV3v1Fs/FlsvoTkR+4iHj+n/V0EWsvvwWU0We/Jkrh
1EJiF7kY8dtjL2DGN7fThsfzd1TMDAsfS6xB4aBWEKZPN8S/0tyDhYfl4+6X
2F1lOho/kQU6g9DmkBXyXQF4GxleDjVtG4OioSyfU9oZU8Zvl1cs8m+p3q2s
eqECUAz3Sn5Fa8mBKotXOpgg6yXQsMIfCZc0+GU1IWtji2El/Abxqkmcyybr
LkAqYZglPqS9RR1PdBO49jFD99hZYjYuwxsrPKAWOcnd8I5WiISnIrd6X1xE
X2Y9bQTGuEOzROBnJw1VXCBXVPC2n+kZ7PjPBr5IcpeflwDVwa1EIJ5Gj18L
2o7EZwRwpRQsO2EYiYwnXd9mIVsNDcOH/p63rPh95y5uwwhpYGpDtT6ZC0tW
Lzsb8C809I+Cd4ueWRzg3C0T5RhtBkNaGZp9d0Y3JBrKgTWZ1+j4RC+jtJeW
7Vz/HXM/HkfGznQVxUmBLn6oqQlEfJhytYv+cIRQv+Et3ZeHhRzt5PT6nEJ5
mstRG677kwuy6Ushy96crfpUXmH1L6zKVwrbT2/6IeDH4EYNE2Oo+HdEBCwR
c6uQXLKR8RwcoyHSeMy7W12BfQBWr3Hu070XHng/NRiW1UBTRGwnkyJqeofu
1mcDQvUIm3dfAHOa1LOmK0eKM23YA+hN9HdAEtt5IaUPrX4ze7uRzpizYvmS
HPrTKlDivDIQG+5QIigYXb39f7dm1TEKTXy20RoUUSMaztgBaQ176TM+aNbc
T2+3AsUmkrmYFEbyzdwyaP9CfxXaYmGOAHw8CzQ5i4uqWERcNHObSzSzc7/l
FJyYePQl3JNmTjWF9j+XH20NjExWq9r3Il1efmqhSMJVs7yVXQ3bwGybX2Ap
EOQH72kaX6M0o1YiCxJd9qG4C9hCw4ktkYFwGjo05sy4SFRM/Xqa2ClzgcIb
m6noQ2+i5/Wgn0YELMGijZ6nvVdoXREBye1L1N2nxVVA6iiRiIIucmp51LBT
2CctPmtBvPKiEdlg7g3+SC3NQQ9aA6KsiAwEaKKQIQ/lsIRdSTtL+RlQfcbH
SY7dHzEGiqUhW59U48johocE2aZXEF+wItB/cuW2DjNf/Gt4vsoF8pxjlQIu
YZ3SDCAFppSmHCjYFXI6w+AX/TWQ9tO/bHUx1UjJ7Abwst+5fge52ES8e+EU
UCV1THR722zNf/E/dP92mL3NOY7ELZDVAIKsUaGOFAGXpub737ZjHeNArzuR
PXEoKUauJLqHqf6P2qFJg5AUMtYF4Hk7VQrykmGpp28PFkF9stw6NgUKqsjm
e+FQaD4Maa/CloGdOZqsm805eSziq3wPfvQUurIIXgt51G7ZmqhRYiTQjiJo
SFRN3Lu1plf8YyMSB4mtxhbBMxrvO+g3BYq19r3KdJZR88EDXzkMUXwZR0Uh
vS4PBIfj/ibsWBGIWSLIbdmkFBVQyZVfGoiKvr+jw9xB8TPHHHRF7S/qSUWc
d3I6fgdo/BHAGJ3F6VYqTZhz8U3zRpSfj5/Ei7yd9N+E7Q0VAEiOPkDzZ9yG
+FUqRGN5YdW8tK1QXHkKB3lVpRKu4n8KXCSgqe99DrmyY+WuLIjejk2QM6Dm
e2/XWLgwHGUcH8nroF70t6PSnsnZOsTvvRxAEplPcD3gSWeZlGBT7SUB3GBc
RcPDznqfbAKAWrs2KMxYcxwTNZW/gLlPIPNpbpwFDoQDnjKQSw0GZmYRhc3E
Kjn/ihGEq7Kpt5D1t2AcksD2wSihqornDzQduV1rC6t1kZvh8KD7UnKU/JSE
dOGWxXG0pyINKMKDyIVVWdToVMqJ9tHFneD1GmuNZu7ShoS9a9gVR3sJmLUb
DNHVpatdx/Mr1JFVdJEHop54TWQ30bQ/HPynXC8PkY/CzojrBMSybtPWkd8b
BZCw8PweOR9CHOjkbn/bT+FFvtwk80D4RnrJ8CI7R4aBVEkQFZV7y4soFbgC
X40xaKE5PJHEKQa3LFYaykEGkTn5VJa2sfgVAq/CV8iIKbA3kl7O3Q8S6EJD
P7zLLwUIQ46g4BBpg+dQtjAb+ByiYMQ6bS4yd0g1UVjdKKmZSxlc3R60KIlW
dJK45mtE4SlvsMiBu/IU4lbanDbkPlyjWQn5dt4QO3ovcmyI4hQxH2pQpzf9
+U61zFD51+SzcDEquAhCt4hljhmedHuXEXA3o9s5P26jcnAa0c9mLhzt3V/R
lGQTT3bExQXxkeGHVNBHuIniMdSpOd5/30/MAHOTnhXMfl2iSqU5UCMh+P24
bE9kUmBe3CpR1FIZQ9dXbgKk9DonZwvpoWPRhWcTJxNCysYk2fCibMol9r47
iCmjR6u0oCKldNDHaZZVdg+F3eJBEfOKOBnIF+wK3ilb5W6FejIoWnSktTrq
RDfKUUIVg8FaqrZRc9Lb8iN5M1A8248Hp8r/2ZNFyj4tB1+kFBDrKRfZcsWU
oz/BtjrqrblJn1/gbUZ4/BWQ4NqDkuyyjsu0L43sT9djNyTvRlPOLOoqsh9x
UAJMbARktXGnD/VYgK6wYlXdUU0OfIje/MAZDxrVOns2ojLshqg0HaaAIj5g
xkwOIRKFPWdqHubQ36RQgPcQkO3lKUpVShaTE2UcnH9JS281HZJkLfKWQbul
DDDXHhoeQCJdjS1o3r+amFaYbh/BC9lEURvQSaomMikbZjQpO3Lv8sONHwEv
YAzai/qHAeU4iD4y/PqkhxSfeKPI4xulRwX5yds/CyKnWQyaE4aS/TIRku0Y
AQ07ui6bvf0W6CvJKERIjIY3keEmx8M3LegvO9nJ3yjO3H3H1J7fouH5Sfpc
+I+aP+brW3+0z7/xOYn4B9KWYvxxJ182VYipha1L0J8MVj5WfPGQUZvohGiC
2IbNNj4FiNOg1XxDEXls/fwZqPANGHLOLag71uJp+hfOabrLG48RgdWQoTxm
mopI3XahNu+55tC1tR016Z3hx4QEQl7FEXHEksonyhYF8BLDZRI6d6wmOfgl
JpT0eA28y0iC4LZdNbEOvy1PDYK3jDoY8/yqaorDbARZ/ZIXjIq8ahfvIT7x
VzNenYd6Gy1I0V8/413L1jEsTBEH7doWM3q8GCVJ/38SQeCGoIYUH6wVcdld
OLo9p0NtGYURpQ3UNH6Pnj21Z5Zx15ey6+cbiVx57zlSetALfmbiUTxvLASu
qEvbW5osrW5Z8VOQ6loHQZeiaM64IMMWTA7RZpYEHp1COiJWYnYqb2f9qvVF
conAxzlD0fz8kwVQIBXx2WZXMqpJooCaoHuNSHGmEd+W8YR8QoaOb/9v54dt
8OYvFXVB7HjhKjH79caln2tTiuN3hOmPVVXGyc0cFlb/7k56fG6D5c89J2lE
ZCXMx8y6Rm4bDWt9QudS3eY3piLFUXts6F4ncyCfyL6fWKP9MyX2USMTisYp
wWJMG8yiEyLbx88QnEOZaFzAS4V1dTBU+2qJcr49o3NbUx7ntm5ViBJcmWEL
19NXcmXALOAms9pQZAqM22ntM5MDNAEnaryDW9TrbD90ut1DkMD/DVM0+0M1
xAXZ3nSdkXBURee4gJYW8tm2lVODf4n5bIuFQDA1QWzXuikvC66HInrF2WvQ
t4ygy1fuXMTP2x0crHmrMsxCJdo1jUec9z38NHwTaqx7H2ZefTePnF4a+olz
7L7mSxyURTFdTxzbuiihriQ2s7K/QZ5ayeWpE52iMJl03v4QIr9oMBc+kzQ7
sziKVZic6sc92cbYhOgHR20mfmOlUwr9xZUMBrjDjAmmvJS67WQH2/IjO84S
lAfp1Enu4EBkniAUR1SM7flKETMGIm94t6RuI+nRsces9vEcI1L0Jw9T/fKA
4U0kvIVDBz+kUDhSR2WXSqA6UTJHQ5iSTq9/IoyrKOralvyEjkI/mMAQd2n1
ePKB2F2epY+0TFIs+cfHYm0JPjPe6Gr5/MZTs/NEjkrqatpODLBBaKwZVqhO
9pZ1dIJ/M+bAis/SI5RFWBehqDH4JBRrQKGksQjwo4AyvrnF3Qcwi8054BDy
4daCI9yXnZI1WSPSYPNX48hwyYc8OyaL8YU2rdASkNPiXcY1Xdu8rWJWQ8Yc
QbYst5PpTWIGg3A684rHCn5NFMT3SBXRX+Noo1aBywX9vqY3xksva2+X7PEi
P1/HR20ghS6N7G0j03s+J3hUl1pMAM1jAcLMjaDCSsTd/0U+/sLbycdZqP3v
dsbDd/tFFOeNJnoc0nvHq+XDrzzvss0WoxlyvwQxUBCYnshenyOuIXFyeu+R
N7vBLoJ1q9fumPhiAJh72fVLq7vX8zRFtwvEjkk6/PY20SkeAk+C0ycgEieL
EhXxixJoqzajZkRWEhpgeGTa4TwSDqR3YXbT9GEEW++iLPmMulD5Hzy+Q9Zg
poEECcpvvNFfaTvtmV6uDOJOa30JUgbloSp6yeXVsiDyrM0/NRKF9ECt4ZyG
7aZBiw5qdFq4FAqkl3hLv6G/C4h8QYsIgZJ2pN5wT7/4l4ZgFcA/mvkg2l9q
a3yQ0XIpv+F35pWbictB5zsxKRgdMdU8LawVMdh+/67ltbbln4m2fvq8rKD9
ofNETrJVzHIJP8V6SPMWwhsSkn8DZGzjqwVTCqoATR/7kudZ5m4ZNEU64tac
z8a1f7rRpeJuHmMdkzNLNuBrt3KPs3x7qpj8BJcsf8t7pvKQZShx8qNJwXO9
VEB6a1U5CMwqXngJsKMg7r9EFSxQIWI6kzNLTlzFcLZAHS1QEcTBmvteScB7
Vv4EQjMNsN32Joy6SeEuoOSqvKDrpVe4UpU7/GzoHpvnI9/Hbp9VwekGL4XK
y8eYWGhyif+VBd9gS/eFzdOSL9ge9D9rcyEsFETmgj+Xr5Q6hPxiSNF+0BIY
GGo+Qa+aHg83i59asYXG83VBqegBWjYLfud6XXN/AoVtpNnOaHJfGqmuLA35
b0f9vbJ1wB4eA0mYi4rW0cop9xAyaheyxwR/XXJ7HlX1k0rn8bZbN7HLzBQk
1IyrOp7q/y/XGaQbxhUbdAEJPOerbNS4lvtcSQ4pPgpmfYsCRy6hkztX82Fo
GmkkjO2UhLG9U8wr3bxE1k+zfmhE6D5ExMMdtkbzAlttdmigRzffAiECAb4I
sqgtK/LIIvo9Rk4FieC2nTUlWnEooiV4GCS+ZBx+SraAIZ5hjgvp0l+vEKUq
AR4bQokFOfKqejcz/HFCzkLijNtZ+gtwFTtW/LngbRZl90+9undQt1ewhUA5
SJ0JZmumCLOX4l4IP9gqNB3KZDFg822Gvt8crgtpXEzNdJ7Vog8B6LULfYMj
1vGTTUnxwVAuW6Ka2abWCn0B742c8+7s6BFLxYdk+KrLhfi+tyKXxwFUDc3U
EQraxSkgHvKUyvc7rBAy+NfBpLjhJDyQGPpnKImDm+IjnLGhFxlG0rF0v00G
zPKAiYnjvFH9FUJbnfzQUDiYe8hVHzG/BpPh1Kao9C6bnApITZW+70xCvytF
ybuX8L6TYI2bXZcikkZb2Lm8rPMusB9sl/lZY6G3IKu+lwk9dqqQ7b9XfR0i
4YuhWwR77IMZkDgIRaTJXZKivQC+Dxs/YDZIo2s/SlzDqrO9yMEcC7jkBEE+
14vO7qhHYhG8BDvlKzTa3Yqt9a6dNUdOLxbe969CRU0G3CVTnjoLUNCHHltS
Ev3EA+3CUIanDgKd/WMfG5clGelokknFdz8T9pZog6O5D2GhQ7wId6n51/jE
+WiYBgoX0vtfWE0MuYMs5zODumdoOV2F7UA2W9uZteA3fJuAZRn5Vip/w0kM
kcp4cVWjaYrRfSsek4W+XqyiWHF1BvQPabsO6RUXAfIH8/lnHZqhH/XDlCK4
4kLVfzBqZDXiDK/7yZGBAY6oJptVMzBtGS/jFaz0pKqWXZKMlL7csCSFrRdF
ST7YbnaUdQ8obSV6Xjw0TMuRWJFScPo41OMoULTbkmhBdEfAuMOgzruTfEES
QQCDBHWxcG/kYQR5eTr0Jch2MaKubjaw9c9faGssaeOku2bD22GN8xyu6zL4
OQZu0uktEx+lPWewY4FmV/S5qKC57t8GWumiJqrqCWbE5kvtBqvgtbHFiYF9
fruZgHSGl/onAmMv0pSpX4b5Vy9gWmHwBEVsjAo6/btgG6Vl6zpq+SwRJdyT
rJpnSh5jp4kiNAfna3CBUIaoB47f7zvl140GP6AfNubQTAYHgoQmugOWal+T
fAj3WYMckX3XB4BKox9MB+gJtF9Jy2lAWLFmMDM6nGGeISbLBrNJtWCPXQd2
lOaMjrX74kh2VL9ZQInFJLsUgeCUICjutOwqEy7KA/55JlGEM0EQ1W69bgXv
wEYqNVXMojQ9PWMxpLR1VPSaeOnroVQ33b8RZHkXTHJiPUJN8KN+2p/QmM0h
V9RpVvZaITnMaaRInO9Bx2/lhOfbUX9tzkiVwjTMVp3hVrZy6JXiOeoPN2QW
26U45pZ/tpDLaDq5sl93AhlwRh1LwyyHb6ZXqAmDuI8CjCjYTXolqMm7PgN/
HHhFdxKgMzqiHRGcb8LGT6kAmJ+NEkd2tBDX7iNRC6z1lXtY7iLwYBctZ2Tl
bw7Trgu0FZ8/EUZyssHhLNeUqKXf7TnkG1gGLMZclPj7vI7zJGvD4xYCskSq
mvy1NZWub3do9CigDR9ODfBcu4Gjj2l+UInQ4MHHdETlC6L5SXGCT82qawyW
cZU4OX28hz2QPMLiY5c5FFxR7kXHEYJ+0rxKVFnTFMYpc2eU94oMlbxERRT7
7uEeTH0Biz68y5nooBUrheOC8DsEDyk3kpScGm8Y5jVFgKRthsFIgfvVz/Ek
wi/daxfHzsNnrenIcudKIgY89AWSRQ8gHsRZHd/JEp+sNbICAmBFLM0CU1Bn
IyLTSMQe+ZsbbuvEgtIOEUcf+4HTmZb/6DmnDUpPOo3AjZRsBLEmPPN2V3jm
mXBZakEgSKa+w2pc6QFKTLAHoFi1DTadLRB5rAA7P8/6/UBr+4OZ3d302D5C
cnJsBQEZTH8BtpEL45BAVic6dcQ1v0kdC9VqZqrhD74AeBIUL/h8ZCOK4Z08
/Wl+KeB8IK+2uu1Q+zRZ7BuCM2WlV+AWJduV3e6CZ/qTgHGSjXjScOHe9d+7
DWkluBkGrvEe6nI+ieBupfvjAZdfa9sso1TFsvdzZ1+U60iLOvHk6+cVCRV1
rOMEwdBl/Ple6zpV3AEL2xT8MFtTOMo60EXO00Sx5/1NCWFPUnVJSrx5JqLn
XbdN68J4GVTH+ou2lAmWED+CDp0tPGPzYB3pjgUYFd0mBgMbju4fnBVYjTIP
74mqn+UfzGHTMLPqTtfgQB9qirPiWqEnjMFEVZlMMn5Vn6wIChIn0Bo+Rxtc
K+N4wCOMmakKkeqsnx8jrMBHV93M9H8zBLd9x7ex1wtN/+kOAawZjQVPnX7C
MwMze1YJqzhxXCs4djJjZvRezSVo4aMwmqXrtXCbfBsV6GIZ1aYrp4ats7Yr
xdE/LFjuxSUc7bAdAz+AvFNYK22opZZdZg5c3uHo+xvEmeEh6l+n1YWCT3T/
Fbfga7AAM4VTDCPomqo+blHATmwNYXqut1zVRpE4v5R5JDqJ3xneJBrCkX5h
C6fjn8c7qifqo0k5tsZxpqjaBQzR/P2REXbQzm+68+EvZkQdSoWBTn3RV/Kg
gmWaanzY+1Ha8cr7Dau3HkyY5qOZkBRP1e4R/67xD22uIVfOOxcY2jrSR8WC
Y97Cm12APjPbDwCDX8/x6I2MWlZ/662mMOdUxhXYHgBgFACRk1c3zVYPW86T
Xvy9I+XDTLy2Vh+mDs6BrXF5+eOHCSpZ0uMreqHXwu2SaafOix7vyjYOBToF
GxvCRIZkgTuOZVD5prCaqfz1juusMIZ7XJKwDe/6Wj74n1upCZC/s1O79xAJ
tT2I7XhOPoRduSxBTA0+HBIXYI5w3pRrJ9ZGSoeQPlyNsn2YdH0SOtgedaud
hNiglcrAa+XElQKM414OF6gTZQHrTOU8EcQe70ur2WxyLG7ngp42CuLtZhSQ
uZeu5dBmzrxgIRMG+VU5lOl6LJAi9FPII2P7tj60mbjXTJp8l1ypfSXbVPiB
TaQl1eTz33eFsxTQxQcjBglw8vvHxiFu1WHrYtwg19H2VcDXAKMfeqDMeZX6
JCDBkAz7qey8F4q2nsyTQWUeJjUv6N97eTlXodZjqvDDQ1nmO1Y4d2Ua5V/P
LwqX0CQcACo6CAxMWLQDBvidYIauAXTPGvIxAFzP+6SsBT0y2iK15r5q5e7d
mdLBzIo4WwC5uGoe6gx+lhinzLyGJAoq2U7IpPvwJBgKkg0pb0OXUty2P3WC
dByFXp2dBeB3GvbkD0pSW1yC693pUk5HibCNIPtnNT7EzikcM471UePREWGA
S7aBbpx6tFr6IERvX8a6dxbEdy56vlKlsNDRt/aj5JteehUTMIgVIIFHe/Xc
HjFAC5Vr8JhunrP0HWMk4T/AvTvnvPAezL/k8iUhfZpkBBNeKOscPs/n7jnr
eY5R4XV/73Zr8B2HABXtFBigy2743LQ9EkPVC+rKiWUMIlSMFcid0JR6D7jy
I3HqsMBD2NgF46L/WGXLSbFSI4zav8XYicuF6/q//dZhRLzh/zrWNzzzrDn9
PGtBtBN0KfTEHEKIM8U/8wxfu5Gfd7UlNYFfKx+9uxWwR4wm1E1t215Iqv9d
LPEE6vEQ9JFBY/gPHgI8VdK5y3UMm1FwpdGoo5ffzrEoFX2AxqtL4BKEdivT
vCpYygUm1mHSYGKdLhCzXn+3O/nWKf/dg7/gY7y1yKsuLzZj3WbUbSzr2IAB
EdKrFF1xDn4G6lIom/6KidbJtXXuO6zCHvqZUJMP4jY7o/SFhrkmxAvF244e
q6fvDi8zRJsM452dvWQWfuO97QYF1y7eyhH/5XTHNZm0LJzfMLNS3kTz4lRP
bCqjTln2P0kAxco6qZJKZeLwRDB2tkFasapC1yUVTf9qsxpY2ZRf/cravzzP
IGXigQ5RFTdl4uLVlefetGVnMEXGtOpEkFkXcynZjqC1cpJezolNYpeyk4lE
DW3Fz6TpB5lUyxpU5Im00plte1+nXGvx1fxkN5H/20FiL5Mru3HcpHrkt984
5fwIRL+5yZuwm0LkZ5/cGxO5r98tWkArQiI6MP4UQC8MmuhYVtvn2ghhkqD9
BvabEih9vPL1UbWD7XaQHaGQbkO7Op9QHBSjT03H2zwlxquJ+HS07UYrEM4N
ulVXY/6JIQSDzoc0ljg0rcd9IRwsagYv6VC/JBwwAffGbFMRe1h/MdjEzRMD
9XGMOwpedRh1nk4hJEjsSUtDvV+P5vBz2wcfgiP1nZJJfhQj6Mx8zaGcHvkZ
JAcRIkk6TYW/6q5685MZ0aZDD2u2sMqdIV2kqIjXq0x/Mt8GDaS76WZOw3H2
QJDzVTcnZF3ImKPVYBzLzqHTvJlSnzFzLjuIF4pQWaFi/CJ+ySVhWZEQDNQK
4bum+vPLPcN+iQ0isuy6GuTEc695RzVeC+DSiWXsVksfr9eRjV9h9nMl7x34
9wbU3Pv2UgVLzUmd4rw96nPhAgiwpdH9GCnLCkolQ7Iu0z7FlfJ5iMl99Pb8
tgOD9BjiZjjj2NH/SmdaeS7lfwiSTkRj2klRP66kb0B3VLGZKARxVvaWH76q
TUcp8GtMZis0z/kykpN7i3LtNJE9G0KtY0t4ecTbNnNe49rXgrN42tGzKM31
w46UN4rJSm61KTBjtE4k+sa3JXszqpr49uRqVfKQvvrWWxjd3ittin4bZRw7
7WaVlevOVllzHo1pC3LkK0csc5bqTaKR+wn8q+3R2/ab+41Lrg15ATnrsdek
5JRHAMCFQpFeUPS4cOXg5UlmkrBBUA3XPEORC6X8AYBFu2RBMiOcbd8xAkf0
K6OvNeD3WtPxYfikqtWRgArf36cdf/Ag4/Vck88Eeyh0KXjuzMlLsRgwXy3q
u5h/tftrsNGfJ7PTBk9hObMffWpk+gDu/k9LTzdFhERAENsRdG+EqPvs6m3L
jRlaLFiOF0E97LDMORJy3OhLoXxlIPCIcyNG2ylqJWiIXICqrrOA7Cgk1hJA
gHV/dDIDR/nqDNdQwFrrcD09CqW/zxSGnvjh+x0rzsj6vzaknPX/jvqDXt8H
rXCTPsV0zb5ptucXupGwHkh1QCcOeItHEL1N54vYq3v6qs8E/MEOw4k8vuHJ
0v0U55Zzz5bJ0zV+P2P6rPzSSp75es7PhKnDiOzLa2Cje2l4r16LeVfE6J+e
eRtES7vDQN57ppTX1+Rsw2eHSegZqeEG9fxi21fZLB9Q2IQs/quURzH7qzFn
wAMms0rKbmslA/snxXc2gK92x7bztuEFgTjVJjVBW9sJwU/MHWvCyIM9vCCC
94Wx86Ni3PstPYeuBBSWJBNz2+7GPoO0OJPeWxPT3PvJFvX6SfxHJWaA42a1
+aTyK8pOEKFlCdxk5Q9eoZkCD3xg13tAaxoEX8N9D+EjLmJycQogyaOZqCxa
AJWSH502lHH1V1kvDyYM6qUaU25hZ6V4h9CTz3EIO37KJEQlm+TygNPqtSGn
9zVtXtkn1PHoQPtbBSmyS5sTc0YYx8GJisrr2GQaQropU9bcSI+ef+46rxOw
GQgHIb82gM2CasqKlOpgpNhotIc7utlqwtFpwPsOruhwZmKrrV52K39HTVV4
NKH85RCq4JGFxt0JnvLMA+7cXOwOhHOkAq8TSGpJgQ5QPB2rvCWwdIDwSaSv
kKjf9zbXTdS74Qg+fPKJauTXLOvsmaQsVFZkBMSOlI9pEg8b3LjV745nTRIb
Yc+KtT8ypKhgWNxwN+eUTL/ixqs0FBomP37OeSaXV1AYg/wYgf4Yp0WcD1f5
HmcvSXc5WKzQUVSqPYlOpfZKi8bFbEyxrAgNcWKvhBGlXjIgjo0FQbpJ1VuI
7cKlOVMCTbqdtlb9PxwOdo/u29v/DRGbPLs3Jm8qdok2EVlrPZO+TyH19vCr
v5jH+83V/USGsM2y1EeOYRhEh5cegWvok1iTVxixLo129hKrUsJCcP9Xku/K
1cDfHKL+oPd9vE43+sbP+NSH+tj8AA60qckh+/XEXLpUBDScPoooL+2TY5up
9uy2BgvnX519hzoOfEu67LN92ZHuYidgZxZWDGQ3erPzEI3ZwuiqhBMLCubO
alwkYEJSjazwKqx7Mg3aBTu0XDrrENpzAriDkrKajWKfw69g6R/psyCVFAmw
e0Xgx22nQ7AW1G0OWIaCMGJSTHcvxfpBQcNApO7zhHbWQH4hIJdb/lgVaREl
Jvb+TYOWoYJzH7YKNUrnhYMDhlYOkJEkFlUFfWIWd32mbjxsKmG7tGn4tI1C
z1ejX6MbSISbOMWEVNs9kJcJLd5m7vWXMsicbPTuaGzyCLqu4bVLy4+38iXd
faPINuVDpWDInMPte2c2K8iJASN3K42r9MnPLU9GyCrhJpvG4i/y0UNiX9D6
hd/cev5rs2OhYqgMGN0w7QdNXhJK2xc7EAkQCU8kP6dvRBgkIIDouGB0urb/
ATv3xU2eUi3n4/4/0HGqR+C6Jf44cUMCbwcORXcveuWAAZ3eCDF7a4nTH+Zu
3ynGAbXvVAIuXsfkzAoSB9sJT23OZzh+GXAdpt/y5RnB5bJ4cckKW1H8bS9P
vYLWV9AXKRGaz963w2z8ITdfTQ07f6VjFzXTDgTtx39CbrxDGRXK0edxVUZX
7jt+pFkPoryDpt/Mof56PF1pI0BwCYBcQtieArBUsLUgRnsMMKJCSSRaJzYh
BnvdXapJe7p5g8SbHS8VvjIn9ihItTXcQ+/JaXYalRdw6VoV105pvVpXcA82
9CwA1QSJ2eSU4I3US++K8BYz7c2Yifxu3c4NGs+sezw3GFNXtpY/oVYkuL0+
jTC1zwVNP4GIfQuZ1Y1EWC7Ncr3zuJOiWZfV/OCKdYa6UJQS+7+PW1YYpuSK
krFIOyV3ZV7UhgNS0gd4XPYHQXfNeG3jNc3omJhQspbacviHHkIA9+JV6Bju
eCo91GbHCLCNXB5qaRF0QJ4jdjp+ZKOUWbAnkc5BMOJVl8c/PJOm/3qGQdEl
hQtK/4XPcDGJHMnNggpzIa9/DtnvawBden8TLBt2L+14GAW3eXc39hH1GT+x
ZqBuIZjV3o/zV/1FeCw/18zi5GJmrXUpfVwR7EcADYjMA0AHkrwHP3VS7PQX
dKH1TpRMroq681CsROu1uhm9fcYPBAlTxZneiNcZ069SI355fdUP9pZG4Imj
2O41Vaitk7DHRVizVrtTT0D+DEoCLPHMNYkqCCXob7wCyDMdyVA9CNlxmKgh
db3a13S8D9MSqU4JaT4yW1XCW672JzLEHF1VZ+Pi3fAGKV34Pu6YrNFQbk1t
jfGuchlPyqfsDdq1hCu/HfKBDesurMnnbs3e9al1je1TTA5pk4i8abPXGYRb
2QWIjR7Yz5NP0hMA2LclxwNjS5iufNg0IjHXj6sz3SQ00cYxlg0ZJOLL5vaj
nCKYAz2WfXifZ0Ubb4QrnC9z9ktKodwJ0DZbYEE0OnBG3gJOmA2OQo4w7Mtg
I7Ysk8JIkXd4FJmsI3VRKXp6p4ubp5OZ/d6uxi/cN8aSdM/L9ddQbuxf5rQC
8ByoIENkZ7eR2opLvpR917vP/LmPy0nBJoowTcoMYY0Pd9wAIKQ+BIg+LwEQ
4QJll8a2pSLw7B/Qb/hA7LtNPtFFaE6PoIg8tFFh8bAhLz64gp+G44jvUtC3
E9Nnkqql1M+tivVoVclng0JJ6dr0+XN1wF0YheRKA1asKnKMkQT6PBjvJAgI
/PM/PvPjh8xZ7qBBCYyE7RsS0rZSI8W6j4zVp99im6csFWtodlxtviqdg9gY
CzNs/NlbDyyY2MGuSeAmI0WRQIBEDdwYg4WvjHT1Gpev1vPc2vQNcWLWAhyY
+fKQmoRmwv3bBqokPslaORmqDtDFsAtXd8s1nER8qg4TO5XEuHFTM8NKnXfY
ML+8WfENgSi9ajXpee2Z8KsNiS984vdCveRyQt0FujTi4DrF5u829aHihCfo
smMypVbskEvFBrjenkYO1O+5FMmfssp8BorkPD7H3FWhIwOI4k4LenC2zQoS
OPA7qk+Ck6Y3phsEh90iO5oZCDIqUXkj9awI2KMnwjE4K8+z7vbtKi9zaX6B
sF0v6HgQKnyYGEW7ztW9S6OuH3BuMVhHb2dsjrlmtMUM82GHJrZCOfjPgo2r
yCw2lVXBSGHNwjFn6yBARd++tEGGCxytTYL0d9dXxwoHxg/ORKD4uQF5UmRo
2VD5XCD/sklimnlpiZig9dRvF8vCgq/e5bnHEN6nFL2be+ARhi/WBR4EVHXq
V16FcaNd10qZQ2RQxUspScEZDHjFTrb85tD56IqOkFhRMe7i872duo3AZklS
P5ViR+mabEYI09fw3YpVWd0evPRkLPZ3ZI2b8I5y8m2ZiGIup4J/OHYoyT7l
Ewiut8sV0YMiQFy+YOnx5Oa7OrQKGJyheNy60yH2K8S6JivbNVq6s3+ZydpV
mAKEw8GH7JUUTpAMuP9SorN3wcRzAh5C5v+q1yhoJYqqtXpqid2fbSNRhIJu
R7AHwCUeOf+YvVpp0o1VLB1LYniwjTjk3n1zd9aL6MTxwgvZeWUXxPg/DFEQ
DjAm/Kqm+c6Hdp8nW3uuzaWDVsgSTjfHWQjBsOO2IE1NCwaR80B4ndcsrq2M
4Jchh7oo8pKfn5xfD2IcXqg/DCNqPnWSoF8O0NBxWhh8mhqcrmeeseSfOny7
teUbZDoHPAtdjemp0maXHB4W9XXU8XA+8jM+3PLlgZ6nWrlQOA05rQAVDgu4
FChrcV/DoapvKcTgPcOT3oSKCgca1SjyQphUPPIkkrqK1CBn1327ObsWL79e
YN8bSNTRVvWcaQ51jTzmEbDGWmp0NNWgLoTBdawj6cUg9N8c9K+PcQcOKm3E
Xlnp7n1xDCWbVeKl/4DplKiLwiIRRbr8hWqawse07TlhE2sLFZ6NetL1odlM
onDHrTkODSnj/NWanGcMbAnamdh0K+zA4aPxq9PGGJyq0lccAFZoYtZzlXEG
sZPKaze4jWjS8FA6QfGPDNQlePnHc4RuluxuKUTOwVlwuZOdWN8LPwF/fIh0
Li9j/M2VHDMitELO4e+QesWay1LpyRm1lCecd05KXyCnliI4mg8HZ2flOdDc
HYxmTU2VT2g5atNe4G/zexPCl1X6INT2xfAYuYe6h0DfEy8rkXRsq5H/ZYrJ
9oMSxzwI5qhouCqngSv6VAOUpMjXSPlb/ymfPr4tQ8J+XAnKU8HCIOnBQtPd
a1/5UwnJ3BV8/yKJG74h9k+wNb/OybfPaePzFBT6GafH7OFq1GLvlkebzx0r
GAIwUKox7/e+WCs4QBgDN6rHADfKgjCv8Q4UYk23U/td4r8M3svIGgV2mSo0
GttP6W0VFOJ7UMSxVuFv1Tw+8eGjbyEvaAwAaY2bnyU3rbrqw+oKT0sKu2iE
boI3RzFZPM76hEpxXac4leV82rVDDqlhPNzM+a+t9vO0FnjEx8BA10lkqaeo
O/qPd9Ql2+osFiMNEKbqvu2H0siGdg6ZI/sVYlRXza/mSjRwegxvS1HgVJws
PgM/QNyNU6ZnfHPnUwiQliepCcT/3QEpaIJiUqfFmaLcgbGHkOUVYcRphrqi
jXclqgE9mwJkE8ZAFleFogYRIGc4UhGd+pn+QiV/sTV52kYPniEfTiw7WttD
eaTAWi2S0u2PzPkJkDtlu2nugLjep5YUoIWcZOMsbY5lPWAFaBwqpnXpfkZS
stltfrHy+n6SRjqlETRHtfFx569Ll+Y3IMuEYPTcD8tYnzqn5tDLZdN3oHBQ
a3MWQqcDBhLd0Abj06HbbU2CaauxuzepaIXryCnnKYpCbYPjjTjO/+auV/yf
ZiaoatLCwjme5gMiRGRrkZjZhmIVKOgDpkz/rzzPxpxkhVxMXHBFkvg7UfX3
+vQLVQ/AZFYtz5zkpnWFxLDnwGTm0vIL6Bzmh2dyCcY/iCCnePY9TlCbhLxR
YWMWdnDjo24SnjawylZwg350CNq2TRJPyh6GsH6JwxJV9GuPReOAu28POW3L
ja3RXgG+n7BhC0OLFL7bbCzzTmdeJmXbSKJq7aQDv4oQIOsoa/4Uvi4xnPTi
lyZEpPulZNJuo/z3NNOXzun7n8QwEIDaxPbiCnrMPBjcS7N2zF/NUEm5sEK0
rTaSGJ3iV09XkqJSf2XotJ77c0Msemi3O08o9vC1B/DL8ZmX6vj7XcBW7C4Z
Oa4n2k4VehFP3y0F0kWtrcIicZTZTWy9T8Ng5oe8iUSKJk6x8+DFKpE/BiJP
ZNQr2TWbNewkdhEG+3dIyL/csu4RrgWJcxF6uZXClxHtedu466YzBFovau/2
Yh20eXhxgYKNe+8bVtzzvEBQh461xN++WCSPEpBjZ3GEahTjn3Lxl2Xvu9sX
YW5bdH6GdibDSFCzMnwMIytYrJwZVlAIIAH8Fs+pg4BY+vrpWlYMpRDCnovI
VjtUoNUxgFJzTpZcWBeZQXZ4WDSxf48qkKqbUHRiKvcD72R77zABLIL9M2jG
5FT+aM8vaTmKWcNA+N+kHi2r6S1SD2ZP+2W5YbY/doO/0Q+rePVvM0+e+hk9
0UyIX1ARAvyAyRVTiYTlrYl/RLPmIgSS80vpBi2k6wL1k1asQjMX1czdhYWn
bFFOzWAbBsV6OyegAlIZgC2OLPD14gMSXu8xvqYPizUamA8S/Ihvav3h1/CW
H02yaK+RQlL9Kl4QNBAYw+zU+t1mNIyVj+JPv2faRnTr5l0r361yPHrbWCZm
8PUu5s5dKyFf30cbYi6E02wrsjmeLxINk6vnosD6TMkZmcale/jsBdjRCISK
icTKccA03ynMONKVEqASXRNgTKnU2kgHm+SeQb0koa0ZMG3o+02xdzN84iot
HDsvzWOc92sZPvJTF/ha0Z5FN6Y7aSrQZINtUgUssvDxdTl+XsG4t3vNntlm
3TgbOSYl7aXLyfbvvH/1n+n7I4jEMUWj5GO91jw6SBD8AENeGcLBRvMYkc5y
nmpKaZlJ7RVbWCmaCU3MQDQ4TJFrjn9LTqfMHv9ObW/v5XWYNLeSYVOy5/U7
bfixgv9UkaRufYnRwUml5duz8YdiI4j5M3yqnrwNBVlIRu7D8ys0YtlMa4us
JhImieMWMal6w47ZsDaz5/j2GqznrzTOluT7VAY6bNdTwMFL0gLe/CSXshLo
RKyt4CUx5rYxxTothniUBN3rbp9jXcuJVsBDnkNJJaaUtKyjJctMcG0+iyz0
weJ09QEgA5RiwGWYyZcpXth0VuB2Mf7m/Q9Jxy6hNC06tZx92KN4pn8m1E9X
rD9KMXa0Ui6v+hpLrsqgpMJxwPVDYduPHjjAcj8UAvxz2MN91Xzv1wipDXvB
PO9/e093OK77l7LOnJBdNv96uucpjiW4trjUXgwMV+CvLZmFUfRra9NMCd6r
86ejmqeeBDB+ajwYW5/pnMrKsgoc/ZYM/ZXhq+x5UP7voQ4evy1UZFM8ydTJ
gnE9dJOWaNVqIEvWIb/EykBEX3Jqt4MQLNJrUqAfD3Gkx1qmeNDbVUi4de33
yqH1G62aDImFo+fRK8ss3sbI0j8+ukhRF2DTxLcSign3gyxRzaMCTb5vj17v
D9yleJbLkmhZH7iGLNLxB4Q61mD0yM/Ajf4ZCfyPDDYyFZLYSTZa9N6UAv8T
2Ts1NvVWJMLci3P/+GdWBn6Wy9D1n6KYIcp4R12y9WgWca4K4H/szJ0rzkkt
tp1yFPEUqjWw1EeWCmDdjrFVWhdQFrDCP+U2AKUdtSMaryxoyVjDyXcXGb8U
+foMuv4mR8+9ALNJmInJFZB10Q7jXpDBQ6EQDuzF4taQlR4v9AHlfGH7xk9N
N3foDpbC40yVroFtsjXVJjFXv23ZmAMcAmygQxts43jhtygCA2y3n/hA9N7r
0B7BmmhrgFKtCbGQhBzOYkvUTMjHvaHOPhiU7/v+jmkYI5krhUKF/+aFnVDs
DZvDX6GrN6ykN8NcsG4H7QwVJmpK9aWDm5Afp6sQQJ2Ceg+v4eBLlKs3rYb5
uqyf2NiW9o4Rlku/a6xdEri2TWdiryAleKwyojAuP074fLB9LMB6WxXu1exz
dWLsk19SRwohkK3zgi6QLQdWoJIdlS3vxhFDU/KfwDyHq01ctpcXow3Gy7c+
y1R94D+drHTwdKqf6jp7RIGvKhDG+LzWwaU6627Yk5t6kVWS/+TRY1TiSF77
3TtoVmAMQJeAnqFP+3uGKqAShXBzDUYBKNH7ACkKvWYvnUfUeeb7icPvSqv1
kxjp9OF1yq1g5L3iBGFNQqyavGIkdiHH+ILzHP5GMTEmUhgHe8lXH/SKV4iO
XSw/46htUHmW3/omb69M/qyWlzdZR9qI3TW3xfL0XqdhwVXuR9b9M/Z7hnaV
A72BEOFlPTcBdTuQtaCUvh2Mo4EwQjkW5CedIiTd/8JW815EgpR+8T1l61cd
DHaJmRWuR+xxwY1VBVtLYOIgiB1qeC3/dev1n7bAVyZgYcKKN7wKMpHbQJwe
vFPYoNeCWC8sdOiKWQ4FRndi9thDZtTef+Wv7a4V6cWnUuVIbbean6Sv5Hlc
MjVWH0YlierqqgbmKDWcQEbrWTSnwOZ9oC/TKyEeQp25qD3YXUePkkZLr1yr
RcTbuvrwAgWqGx8xEEX/TqxVyMneUvJzCilMPmZg/dn1BWOLN4knR8b3Bx//
xNjF5UbqDOufXePcLshke6HRgLxgpS4F3mndebKTrTgWgbUM/oZ/33tdycND
csV+9cMQWhev3IafgN+sR5mkEctLz+qWrpg6Qk6BRHaQvZgerF+t3IrV6jks
B4js3aXG5Oyi25V7RAgHSAm4v0f/IhhSannWOrP1ebXaPYPiG/CU0qDsr6fA
pxp2eE0Gv6no0ZuJpZI5EzeuQ+d5iFx9XcepVw2WjAXBkYzs/Cga76nX5oq3
ta99XCfMEBJbsN4iVMGfLIdGpAML2XrWwNhTW+UX6UCimNVXvDjfgOxhGFvH
YAAeZNTCOWihLSz0lt4G5bZYiwLD1mmlvM5NBaFvnqhbuV7jqrfJvUbxbJhU
TzS55rXv5t5dMWo/Y0bex2RLH/bgawSrA+s1YeLIi896qwa9wXXnc+NQK2Qy
WD10TUqz4ziuxE7varUPJ6ZuAJqjzHmGK2SWsivvUqKf+74JnRZBQZNa81Nv
OkxxRgPZKW/hnqYELOW00N8S/olklFba1ynvXkvEMBe7m/FK4b3enTPy7gCr
8gIvnw9A1ADRMfTA6OOsojU06dGnfoJ/rpfSiRgA2SzfsPgFGmkch5E1UISQ
Y9PPch3wY8bx5PKEauXp7iW05n38aGf6Au+5hdySJxiqzeDnepBGFrq5hnlp
rG7jURuwaRCzqagVMcbA+DeaAOFdTUgZu1bLejqgn7W5K95Qdosq5ar/nHKl
RS05ZpvmAAyTbA7KZN6EyF4gfAQdaY1PKd0wI0fe+dMAUivToebm2JTqgRzm
o7Q7ww1e9y+fk7l3JByyxqesWN7aXqf8x00BjqW6kT9FWFEcBKVQdqKrFbr0
TOiJ/x+5IjQr6R63w/A+34OuO5D1yAeuk4tNjQEMinRixJA80yEauluRhMjH
lCHTUcXwre4bBIRDb4ChRnVF5GUpd+XpHSyNeDx+oOqgAgtjk8cQ/V2Ppyin
ibHVNGlh+rhdZqSM1igummkAT/FrGIbIzBJy4JCzJOqrFCpk6OjvpqTVqRDg
192EG2DTVV5WvT91Ehd6SYg9N5zgRcd1Yksyuw0rqoleu1BcOh6bwQYFyFgv
VoqO6uaU+EWJg4AqgzDZGVgtX+obkjHQY0Hbf5ulB5zBxJXaVHLjnafa3rZH
D7h+qyj5MuEx27Ju6yexMFqP8CrWYX9psltEIekVsEj6cYRf60GvmBqk51PY
lQXa3a7SVkl1tD+X+NqMrhikqEKxxkbtMLe79JyVtZdkpIcXN0SUflRSmGXi
H3qVuKJkBwSCa7yWfNAg9woYnMlf7VtS+Rsu8XY4n7Vv9Jj4RG3jjGBgl/dU
u1bzkpExgyjDMpHg6wpE/ca1/QYi8IgIdwL0hsJ/xu+vAYQn1s1jhGCp917B
7ZCciDM//2lUThYsHXN+ocjLvCIo3cfj+cU5MRURRLJUh++xGqtv+fCXVhWe
KjcIjd7dudmy3N9cj/wWBrQmU/0tp8LZciP7SzP3BNWjn78dmO4XHQaOm7aQ
d7yIwHT0ETe5ZAXepAPEvCDhLto2CQqjsGnF03p+XjVLIuhHx38EzlBtksdh
/4I4FrEadQpPJczMUir1q+cq7aBsYGMgtG731FnVuQDD7FWg85b00Y8J0jip
VO4VWtuvOnhlhuBQtr01vzEmakPAVtpBNESHVS8Jn1E7M14lyrPoQUQpDY1m
/Gw9OVdpFs0QTLMRacIbZeY4ZPqeqs8O4xaJraS8xv1qa/JmRjBCHLgFOgwh
xtkK9IO+QnAn4CdzLYpSwALyDG+xZOMVj01Fj1can6UU1AlcIZ8YA15BPV72
X91pnZF+/6yZBIsLwKaIvvyt3Txy/JVExjUVF9LcwdrMz1hvf79cAPjAMzKk
njgyh6FjE0yxh85OZKC/+RcdaMjAvXwfaI9KeRcr+MbJmit07DtOMTymDgQe
mTwK+eHBhrj5Sfex1kyFycianmFDqyh5N2o1hIyJBELLc7cXEI31+pgC3sGy
AFwjKntI/YpgdRBDPGdcpS7ZV7Xd7lrYQg97qB+JnKLSHQHMZPUbwncR6Cid
sCPcv/p9J1EPHtPB9RPYWvUyeeiPm02Qa6wf3JW5wbre40t0MLqnHT6QzGG8
lM0/7GLNBm8XcY8g7aJk9k8tM1MGAqKy1bBC1vq0xMXo1jhjArWc6wtoFWnb
FWYUSU4ikL2a5bEJE26jRfbBNgchqH7hoGJ7QpKxwnmbrNjUn3UfT4gaPn8K
bD4L4USi/smeum1pmSi6qNFpKhSZFug28wC/9ELlIBNm2Iv9iP2Cco1ulKuU
fsU7z8evNgqlx52TVdu1vBwXj0hZqFItoaWX95O8PFSPcPE2ullVTixVxwPG
EMu76XmpV+9nszpUv674jYnOihDY1ubCMNIxvrNqBs9PkQ4RuZcfAlIJo1hK
2G4LZZRNcqwVZRMT0qNI5itvmvFUyxuqYX8fA0Sx0ixlaxxv3LAOXf6Qtqly
JN9I4D0899X1IQ/MbEJuuOcEIGKbAshu4VH6OiC+WIlXA0VzON32P0pMR6g8
PbEt974znGSOrxvGY0nsE6nY2HqLaRVCEsW5kA+LO+qkAMDaIL4Kr3STXnie
Jy5St6/Q+RZXa6OW/wQrNca83JN0RWRknRqaN6r4EenRGshuevJhJVAIaG1X
1GWoUmwMYoEmjSI0zCJ70Iye5C05mkGbYgEwsx/Yk79d8S3IXaDpidP3uMXa
y/jqC9HVNVfqDU5Qg57yBokWL8f29p5+FKGYT05MTQzsO81SvAnz/KaPgfH2
KdjrVJEwQ+DoEQCW348SxQC134WoO/WwvRMiB3vMCU2NumjndVkAGJA9cIWJ
EHWWhopkRjWYruDG0UWPVfy/fHrzMy0VyOnXNQgYxp2H+acOSyWwCTfqcLoJ
1YHnQk4MX6k5k6VUqkFjUsFun7dMtK+ChsLgkNA+KJ9Dt4Pexu7B+icQGmHX
UoTWWVYGg9JFNbQ4BOKEDgHcqzfxRi+ddBbRQ7CmiqgOjQYsKFST7XLNwIK+
HDxa7UhcQj8RdbF40hjmJNs8o5iPkO4P/LjAdi+9gIS8C9vyS+EPxtzpm56o
MgA01WHOWG/eGh30Ue5EYI0Su+eDkZZkHRC0BvT/rUrRn+vlBNL6S1gkXVsx
uQj+pzl//snIp46QHb3q4zhcT3PQCg3uEUst490Y9TS2jTUKhuVoBU0MLA+s
8hOf3HymGr1EXBj73+wRrVobbk+bVQCgraeyoi3PrbIowGqTlPOfIJLWw9ol
mrduXs74hZoV7eA2HSLg8bOeqf1/Ej5EVuaQkH38eg838LyeHJ9Tiaokuof8
/73UHrw/6EWKlfk8Nw7i0cAHwwsvyISU1XP+r5WmztzR0055ckI+yAnBu2xm
DwjttsW5gt4/mHGmVgqm+dCCyRiiOm9FygY118BH6TAurbXr7dK2xhFoHHWa
sfQiCqzMuPnCQLO3Fr4jam+KpFpx2ZzVrQ9X/vlt3NvKiY20cUZauI1hFTcw
MiAErtjGfnnFWY/wuidLmlckh8Lnrn2mQ9moTL3gEscaJ1Mv8OEtmETwYHVK
LjlY+QAEpDb7+6xS11KYs9k8QpJ/IjUJbA0lSD6OBIFzKwpDSMIZmJ7+9MkZ
IYUyHPT95HoFS8jfD89jvIu7/NUL/dDa3AZq7YGs97t9rcvO/xaCv6sQtN1E
EDvZJrRpV5/TGjoICQ1Y8HF5nRWqencdfwupliPiwDo4rxdzVG2hsUKduAFc
czsDpYdbA6spq6y+7GHEftcE2UV1vfdQNVkCMoha97DC52Aw27ttEaS/ycFF
L/pz2F4lboG5B4MxHG5fZyJW45/1ut64bZXMbVSQnyHeU3VYetveTiacZXgb
WZFQLthsXVwLJSEoZ29Oimr1TvXGARU/mou82MvLYp+n2/uTLiifGXDxjFYE
7yppvlZs8+5yknPHjBMiYa0tH6RMOWwZpajatMwyorWXShunnd4U/sY3VXJV
JZNRszzEDTOrXEun71YVtUz9XQ74k+uV1ZThnhcIfg5QG0yP+vof6ZWhCQj9
XX+UEDIQAIX9EJFjAd/yere8vvC+snOko81dvpC/nth8reCnA1NhnRUTOrk1
l5eFLFrYCsw+jHHpASdZ8zk4ldzu+e9x0TyLDr+YxlUVx8tPTzPxW8GtDZc9
z4pO5QoumNGjxtzH3AxLVuUaKHYqp7+078f45/ad4hvB/d6a23VhqX6u/kF9
5oTnP/LfG8aLUGp728CH8I6iAVHoIhncz7BzSy1dDY59Xe48zLxdfcIcKOQV
1tKttaPP4b/7AETEwsen9mvbPvP/MuKFW848Ra6/zzp1VYn7PrXyamcM69dn
AzMVOZoZcZ5GORFmH0D19D86saKqDjQiLCEpM90llEJPpWN7Hl8G906UmceR
+lt3pDHMz6ILh1WHSnJfx5OxPgZMXpLhFM9L6hf3XQGdX+0lzq/AX/PPstdo
cEi4Y4d1UtC6KjchRhRz5LBivuMJa9CevePmKLK30e3S5DTgbtHGAO4Vmpki
qev1tImPI6wyWOVlonsZXtGRBp3yinTpZuk18iFSFuWdLpbxpnJp7i12fS4M
kBo6wMshUZ6e6qhTaKHOCcmLZWh7PgCgt2c/0aZA8O4MeNaBfF8yxPIAgXen
HzH/zmBx0nOFZCbzKgf169a05ZIOo1fwdxXHkxuFP9ipHawKs1PDVGCmRyyv
TSdXFoGT1+CFWioAjUEFwF6oUKT6htXz8FkyEhuMynKb9ehCMYb4nYs4m5K1
Tay8By87Z9QarxYr48CmNs/gzz5oS6ogTLouZjMwy8WguMW0hoIR5wI1Sgyr
LRu3So/hidlAHv9gVnX5ITD5KOTuwF7AiAWkBWecZ9Edivp40j/1JTEIBxWT
805IGApSOBJV110gQk0TbfHiQ1ug2xDHoIMS2XN1gAj6iNPSc9KJXBy4QabY
AR61lBVbzjSXGp0fKSIedmgiWsm1Xjho7DlwIHiSj1LIEsozVAoNQFpphxDR
l7BDNshIlMvW1FtY2/LVFiNUDS7q1PYwWZxV/jbenx0OXPYK0BY6X9nuiJJa
FxIw8j99AbOKQ7I/nbOoVamWlAIfxpzwjDn+mDxW7ZtmA7Tk//35gTW9hErQ
6yTLOTS3vvYLaiy8ufJWKSLnS/k06Nvj9QzD4YeEHMAPpTTWQKLgQS4oPjNr
JKUdUA8XUJqPJvS55JTLp+fwAPHuaUzUITZVY4AAV85iA0xeajoMnhTQQKuz
k9nON8rrBncDJ1m09wSBHhfiKhfYei6eGMecEWpe/4dm6IVhDUcXI5dmeg16
REDlCivzLP0H2BCOWcAj01cyRY0H71+7X+qEqNGlqmu7mcHfR0o9NaqwGN/H
RlsDGrlxj1Sv0rSdWkuzAd4dLdpUbsS30sU3FfpS3DK6Zz27HI3EVfRA8FJy
9yNyzVhzE29kdMEU9QR4V/WitVbLP0+6CgCc1kuoilGryuBJhhseD6jXXJzI
pK+xAsSKFEeKi7q/HwKvYTp20cDkV4vpxV3PmTIExydyqqzQ6EDEq1iSn7Fz
Om2bZN887kYxc79hyZnwTwgCZ8/WZFNnODuLBn2g4CJFth2zAKg8lHD8Isi7
1C2w7K4qLMRVjWJepU28q88nGG5nyRu7bsD21VX2SGKPeFp4DzEgxvx2p3x3
+EqqKCUtTguKNkCXok5/KnQLBm7ydQRGKJeZzr74rIuEqJ/sKhBxLIkYsdf1
ZqYfrMnt5IcO/hkrC0Rdj8jvvayEOxDk5z0DWKCHaRqetvGuTMEqqkG9mH61
gnihUTBdlBkky1m2Zg/W2TDectiFWK5CphTvg2m/kd7n57Ng4Ww0QIcVL/xB
LUdkC+XlpX63SqePzg02SD89siAMHrVee0SvxddOI/6hU5OGmzFMkFQHOZmO
xD9a9H69WMOKzsveMKLQHBvSz+lF382gA47OhKeBR15mh5JX2ig5oRvYT7wZ
QJ+kqKanp3hcW1xdyQghQFHIhnf8QA/W3K/Pzny73+8IHGKoR055p6whG2dh
803nbB2qlsiI19CxW8GXro35q6bYz3K2h1gjfRDnFteOL3RZtt+Jr5ll//QV
pvR7PcnDF0HuFwkkyI4PNIlccNgS3EG1DmBZV7Kv8fHPsQseLQ13/9DLlagm
Ig5/U6acIGrXyr2My4Sr2YKLLeFZhoRfo0b9QxmWlQk6ZnzRJmEh9OspcQ2g
96CEplo3uRF+M1Xdn1OiD0vqVgnVW0/8JMujX9bBskCkljfgSJJXSYoH9UQy
VXvE7di8Qse2QCjlpHflOPXX+vGr5JehoOYr/6ILKKGr2wCZH+wZ0pmVG3Zn
BGbK1KxFpbINMygpnCLVLDviEXnNDRWRJx7Jfz1yWfQ31eSXJnQsXEFLNKsC
EaUUY5YtzKmAJoiMx54Bl2A4VpK6PYX/HtZBxSx67yWwMm1zxgMMQ7efTQQt
y/Gbl58N6fuyCZfbeAHjO7pZ084GrRq3WlEyjNWrHnB2aWzjW2h/HluBU8Ug
RcskP/1hltlEma5Ky8EdhhI3eA3lemRFjdkG/VRVTFoNMwkqoBWZ3K0BYMZE
pNyyQFfFZNPJuhKfVwrlcbv5yOAmoRogj+fl35HaqoIGIAE55/roq7o3M29X
knhKwUv0OaAHmOxy/ELq4uRIcyetG5hBuriIWrf1fzK70lNFTKoCpus/dIu/
/PpfT8bzuaTmIsCS1jiUkSANfseL8ucmPovC6AeQlYzBpF8SGbXHUXuEkVl3
9qOuS4pL5mS2n+jVkj+lBd5ncp/zF6tVNWdWsUmbe0iUIGrESu/Nx097LcpC
xUYPZ04SCt5qMcqJaq0QrEf+IO4XexjLl+5o5+nsIEqNei4moRtuj/lvavE3
FbLaQKXA6QfeultHcyfONdCVVPbNhU6mQJqGl17I96HK2762jkRkaV17Vk8c
dCO7FJIO2QsG0qV+K1Q9+6nzkzakrndzZOFuaMpJZ5A9xdDeb0Oed/hULrai
9Q4JTZUcSLXWDDIxUDJJFnQ1mC1INhqhiKFdtw+60Y2FAGEYmSzFcU6u2Is4
xJVrAQwcjjg7xbL6oRYRZ0B2WPKgDdLgSS/P59PeLYdy/liUJP93VmHpCcQq
fOPhTAeNFxNUVaohLRcvHqBrttVi34pUwhCHNOBDSKp9Z3QuWMoJ6RaGHps0
VWfsn2wFz29u+cYbK1jjw5VPqBynfCJdDha3MDFFNRpNzZqwZe+d0sRyoY6k
eqa12oZO+31l5gf9PKTO4gXVOoXWGuTCofnVEBbXfTCDo6nSEa38z1V7jRAC
rFX8+md93Sh7lZDohccGn8R6yuB6TWzeD+8WwpdwBJUWNWhtkNhvQhD6O+R+
vN3Bm5vTGLRSmsHa5Nq6TXICBmAoNsr2aJItUd7QeiPzQOpvWixxDx5MKTQl
fo5uL4LwSJMgieUp/tVh1e+/o+IBERnYXbU7ntCOUDLNrFGAvDvmiU6JjIc9
7sGpnEAD6hSVzztfpBt5f0jYh/o5LazjU+jEaGntxfe9FSiSDrg7Qr8XgWfZ
KrcBl+JLHgdnJdObWjkxoOO4bH3nWp6fJiFNA1alx5P04aYor1NsW5LbZdGh
S3stuB7giXo+CgNYWhSQKsUW5qFw+BH52XR1/tbciJOHAvo//NUWmlJslXgh
daBFONkbCeFy0Qg+OtMVGwqScN9gZ3NHjKSo7wvMOcMkEtdNuo/zg9lG5sTG
kxzgEgD5s6NwEPpBxOxQbgRYeFRy8esSAygktrxwEOzA5zkB5rtNaLDVTyeg
jxGlwMli/+SPK9QkgsH0y/uklRZbOFxQPQPQzzhKrUEzYZ6T8Ufl8Ye5sbvm
vuDlYpqWLioIJLyjS76JFM/6MPHYjO5xDeYOCFmjO2zWKZ1+jIcmuqUDxYvs
9qMPmL3kdWQHVkT7FbJcZZRrYWdeADOoQ1Hwd9ABx7D/LwNdkRY4+34BZwcz
3mnTKVtzr27DJokBY1OjXdQxZtIt658oEIiLjp9jOjfrWhXeRngmcmWxTB+T
KEz0jwnbNoTq4YJiDHMCzAtahiw0wQxnxGNtKHlxlhmrSCN5v3U9btbYs6tI
60MwCOKgTflmaYUJGNzqe2JdAvND5px3Afs6Y+H1MDdXENwtdfkv91jA2U1K
hwujSW2yVU/B3Jq6hOXKfZbHcPknPR10uc9F41SstHL8KJlxObXTRZ2fPKFq
HAQXoJYYKtojeS6Ss0A0pk0CbDtimSQJ9/WafRYSoEtcsUqH3B4YA+Af7j/b
4RaYCm1lz4BJNBUiii7XPqYTN8AOYL2suYkHQYL69lS0YBjCvpl94lTs9KtT
Pc0LarmmBguf5iu530jJro37P+uBqYmCyqRvW4gQxDiViZ7jgaWoAa1kVP9Z
KaAduK5BinbqOrDKS3M4D9xWIGXsyMgrzVvoTSvCfETlx1As7DXgHnoeJVBb
wXMvdhNBPEFX+tEpttsKa5uLD1tyunikKzyQIfOzCW92SEu9iF2Ap00qs3Bo
GmiJnSH8cZELeJNBfPjeFA4HX9q9nSU4l8imw1042fRpNii5Daroi9zcqJn7
pLr8DkW1QST9ZXgoWBJG4XDwoIzCgMSUxy1GwDEvpcekvAYetWZtMx4HaTsr
enlSHCzpS6ZJe9u0u27MWT13CsV2NUY4V5u8LP4InEaEAzrqiy4B+w+wmsxL
flGf2CmKdt166hSJvoDNShuvzzRPPdtlOvWMU5TcuGp56yW0ufG/QtG/XIlz
u+nmHZ2RBuDs4JOQs12OFheBH9QKbt5efL5m8xa7d3gpF3NqEqKaviPRfN28
WTTDa/KWI1d3qatusz8xltqZU0LozF4AgWORlxPchU9lgwhjKvOrew1trimr
qXrQjHyxnGyX3bVRo7SZC15z9Z/URJUagwPqHsvdRz1MqXLnRImdVapcHTfC
yXTqpDm9jtPu6Jk5BMQ4YGeR+coxMl2HlW0A7E6h3/gDnI9kC5CIcI4xmJ/H
0pZmjCLdUt7/ahS15ARp+hCIWVy1eOQeMMltgk0roA/rYX0h2mtbYF42BbNI
Zi6EeEKOIZ+fGFTFA5541KSTMptzbkF53HE6H0ElIZ90lwy9AEghvDwpk+Ij
pPEH7ducYXyW2uWjPiOeUbjDJP9jr0EnxJ1UgtX2FMS66UBVPXbT9JNXzA3o
zegpUs2Kdk6VThO2F6VYGVHTPd5tJGl6ZKby6LojK74AvmBFqMvqUnbADKLx
WdHBUaVO9YR135Jk2spBnYvbKeJwVScTr2UKECKiJhymoFLqbPrxnWs/1gNg
GhbqDOHtDPG2fjZqfTTLcHKoP0J/c8QAPGj6fwrbooPij6Nt6fZQ6UEwoGCX
g54T36w8OCX5Jm8C2P0maIrXM38UrvcGzzzaVSFCYUKzcLCQ5ucrLmzqHLEk
vrH1xK9YyYYYAj6eLswrm5eL2YWIBxM8/RKIWRZmI0uAnFkCmopy3ZNixsAM
43W11+f7gm2O4TG3+/N/ufoahbUmCEiykioTz1U6fkwTBsp3z9irYh9/0pA1
cK5ENKhB2Hae7hXeSzPMMHFurOZam59owgkMdzRZwPO/AFLaPy2gX9drbdMt
3xNGH4+f3xT1YHB7+wejeml5MlQ9mhEvn0E95iVao8T66C5w09B6k5LE7ze7
MNMiUIlHLNGzKHFNxR/AKxh/sRQ+NmjwCrlBNJupNnYodsg59CKROkidGxHr
0ZhzJ/w4LM7g8Xreix8Efys0FhpnecfPoD+Egq+J3XdFi3m7xgwWrb55oMCO
GhmPdHA4SJs8svc9vlQPUlK5NFdTLkxHLbmKp5MoLfUaJLSd9Ni+eyKUhdmB
B5YIMfZARUUDoYkNbmQqkwCiEohtep51/ByPOCfxt7fL1oUT33E1c96l2ejd
EjtXi+71U3BdR7PJNyoG3gqilVCzkUtcqyAljF3jjupcbQ+Js//Lt+/QXazH
2NwEEMGCnwx0j5CU4kiHBITsHpJJ+uOphUIQjyzauOvG9h+45Q+FcyIIvIwv
bPODoyMM+7lNpSJr7pXGO0l1RZ2J6kwRgi+K6GdhlNKN1PY9sRUDCYGuNGLf
RRiGDhqf9S28FP7y7lCUoR6VU9qA3XvBH+xxZux4qTY55XKRXrRFK2lzsS/v
Et0AheyKeDOzB4djAXT3PYsY9RBSe1NDvYgpxKDbhSq/IznGsL3OOwvgOPht
wHsn3sLKWBHUmfNNnotd1ZIBsJtkxrjCbF/HULVRns5sd3hINaNJI9rWoGGK
1FcmOcA3l3HISbr4Ood2LepcyYRVkLlAxnAAMMpzunIXZqoVOWc5O3jjHqmC
+jYRaHktmCXwdVF6H6e6FAkTyBwB4D+fusyRX6qaFPAEa68hT/xoVIRhEb/8
IgcEkoZ2p9VvCj3jVm2eZvMo4Hl1n08No0hD+53uBNw4urPqzAW57s3F9vFO
Vl/TnMANMB3uaJq0d/azK7GsmcFtQJAwjWAUK9upTCF9HfkDpEbYQTbU0SBa
WYEsezYLok/GsZwIn44UhmEohjTm2eQibflmRhaBuYaB3PJ3mWFOF1LkPTSt
mnyiPVStXGFpIzCqjHO0OxmNO94N/E9rbna6xkUekKv6msjSIsQOEATeyKoL
HBkz+sTZQ4wcgZLWm5W0qCzlMVBRZfsoGAriwypSPpCBZ5BrXM5HYdOcJdcp
Q3WS+zwhQ30vak5nEOrvHvwEyLmArBLhlxNDSvjnspLyTipnaCrWGnk0LTZf
aKPXEaSJR66uWgjiqUcskFtNqIKGq9oNOYB4W2ulCdHyCH/9OcjeTALch3XB
0OAZMkhgBF3W1bV8eQb+Aef5ecHkpXp4Bb4WiSPG5YaZA9S7NryDQrupNdCy
obW7ynU5xCuBslp0peRi903IbuAsRREgv9hBOzNKCJ1hobNr0m5DYz1EZ2V/
IdboAtD78NozzOWlMFFSERXlIfBWB6iQkSURDFjll9BPK50jH4u0GB5SAjf0
tQfPqtDBYroBeAH/4z43MubZH+DUeEuQdXMtGgebWSBv3dIRWqkjJrD6P9W5
rpunl2nIU12t1hdZlzcJeSCCW6N1lUn+ITZkI9iy22hxItWSYpwkYfGOqhzj
XEfrXOgfVyD1lq4GJuO5D6g0j1YA6LjZ+wLYgQAwmuNlHhlkmrMBeJIPgrjH
Kelw+6Fv8YE2QZYmaqMpadI4KZm4pbrBEyccIfxU6QMa1lr4VTWvDz2DqsTi
hYcbYJ6F9HtTFDZnaBvBTz7FnjZiWmpYuxB/tfAQ3MTBYxR+RveQNRuekAyK
25lyQm5ZJ0pAzkWJU40ioVEl8iExy0683wGGljSxW3EFqJIOYeREIubYZ4GF
tN/rXtYzP3pUQHHKBtt7BAr6SsBoQ8mcrS0hDAfF6aj4C3e68xn/5iSl9j10
I87xh/dxToTBz1Brv5YysIX2xUiHz2xkJKz9x8laRi9u4CSywiVLiDAI7eIT
xRF7a3aLk+YJQPiA9Z83jtTvLQRvIhKSWprbaSxCS5sZDajrOk0DPonlWTWR
KwyjONpC4VNy1fe0ul6kVOhGS4/LjbXDAD3AhP0AHUZ0d64euQixoHACsDVe
NrFNoeIqEBkaI1s3Q0HuzA1F/lh9AAeEK70m0HjHgV4mfYFTy5DlipJZcUg6
wZnUzfyT5eiGU+mIieHcEsW7p8dpZ29hAiNfoUq+v45dHUyxM8hOrBL2XXEN
Y/fwIrhxs3BpO3dmoqSqeSzwctaajCNGOYuhBkbmlE4vc+x+UkHHX+RAZ+am
qEAVnb9mBIefDltfS/vFh5euz9OAvGppDtOPC9fkZj936rYgDmlVypzaFTS3
7gfAb3X8BXdMIqq9l64EMcSkZ5iBDZsoeJDG5MpHKW+FeRk3lV1PH1HbOcCw
Qs5dDmn4JLYtsRvEbvkcv+D+G1KxgQaZ0slWLZCAgJ7NLPwH1npwQSzKWT5q
MVJ0UAftdi3KDRZSAMa99Q3gXKUC3EYy/ExJzLmGLRuJlvy1qFq6Snyj8wwz
sPtl//WqjvFtsF8TY5BMgy0ngDi1gRR8UKzECESYLMAOvaivAW4lGj0OCAKf
tU1klrmqEs879ZtfUXhWPoPSxZAGWTHAlYUrYthhu7bsZrrY2Ia9YQht9iLc
CBEvticVeHEcjyY7UaofFkPks0RC5oQfW2hdG3dQWPiW+9sHJVgWrHYWjq3W
Gd2XpkFnvk4dap6BZ3WGcbCkXdSDc4J6l9XJCrnzylruQf+OJlJVLpL8V8m6
t8n5agDuINFX/kFGzy4ERep6Ar11ZBZOLUY1SdrVLLdg+x6RDpduP3dmQ+Jo
418+4LQRXyPYfkJoHQeImHZU74yLyaGoXX1GtHLugUObZpO4ACYkRsMg+iOu
ck0SRxTgp6RO+YE0DwhEKkYewRvPy7ReW7mC1dom/UwBb3td5nXkdSkx802O
H0YjSgj4w7W6LDLUcLKajwdhJENuvX0O3czKafgdtG8WZ80Ay/jmSIr/Ps3F
uhjARKYZMSaRv6h+zNO+miUtNEhsVObcMzPqQecTSvEj3IQVV8fHC8RUQe4Y
9bDsFyp4gFNDQVwFHO0vFJPX8l6X+ME4Y3jlVVP0gWSlitfnHXkBRcpEQrsp
kXbAztyJyX0YXAIiIcwT2jxdSRLYUHGxNLkZ+Y04zKyLuEnSAB4HgvINY0Md
M2USf2nmaC6XahY0dvTxar/PHNs2Re9u3Cw1nYlWgL9RcNQO7G9hsRSrAdHq
NcY3DTkBKtqxSJDLX0vSESBDEKi8mvZcyi9oGTHMOMyKvd70hG2pZeuY40IV
aGXgHcheiiotVlRMGU6glBo5FyaEETWvT2kVLy/aDe7Gm0DIpk9q9GYfRfm3
U/8PMU+ziZHfCkdJIiTMi8VOSXQwoKJc8OJ2rxWUERX4pThkfHfmakHH235W
3BV/QdjHU2N0dQJQv+jMaDpHS4ax/rHl2AwFYCKL3FWaIcX4B8JxSHPniURr
299V3R8UjgJP1Bw/9Bnl6k8OlxxojN9WRjJrcyP40DwDtrFuK9X2C4l82pud
tKtnthJefEMPUWNZ0ZvflOfqL0XhMPzRqpbxonNWZYsBbsfNF1IWnsnkmNFP
jxb8Du5OMxtxGv3CwyNFOfHzUwR/3HK4Ffo2aqVWDWPGcMxy1ZbvhRcVbGVG
w18nVlnZ73kVeTZX+cJgZLbPPFGTByuMTRQzPHQK1h17nv0m7gR7FrTJOUB+
Xs5/QYIdq9FWFOA8m/TGmy2DS3PPmiaDvC95M0ChnxoboujjguIUBItW0Z99
vRKJhtqdb6Xs8BqZp0dz3Oh7AMujGvc0zYRGJbDYzWOexLa+LbgQeidP0tio
M4s3CGAxLXXi5U2jxpsgMmS76xhACg7abnYi765MTu3pTIz5PmHXtmGEgh/x
sTuebep0naraYPmQ0BZdBxlb9XcwfIK1ikVIaMu3ktjhXYLLsnIkvqqQ4VLb
Ap++zyAJ4euX8g6ASr1+242OvLwW9qV//WVsmZzJR48xlkrhhcua9etxIwoc
NY0TX3eI1Rsm5eFef5gVwv4mFkwYLvYkL01vEBmCsfjKFylaTbErTpVvASDn
XSzuz4ZUDOhKi9rJJVtZ+3juVgFrusM8ORCWy5s7LuuWcv3aBjDcPr45LsGX
+K2ldu57V/6fP68KWdM50Nbwnyu7cCVWlKvODaOKkLdk83EFi1MIHJh4Agr+
4WfQDF5aXmUwTCN/XhV6tQMBJahHQ5NmmWXnQMAfnSBOTnsa+cvrTjvraox0
Lnca0fREiOyhs/xS8gjyRCXSfcYA4W/PFxLSsx1lGzdnzmelA+XO6AesnV16
TirqTKNl1hcJLJmX3uHzHrlmgrUK/61iAiG7g6Tn1GxHZwIVI5tF2YJpuJXn
z5/nrqIEPrv5APynwQHw5VJ4iohcqaFpnZJxugTDSkjR/ozZNLQRacS7PrX7
xAJ44anx+kBwDHXKIwZIsROlBrRpOvwUio/W7VlOJ1Nohhb1KHmiXyEyVGZW
Miwb58W+mqNzmLr/cs24MLEIQ78bKIMVHLxl2N484+ZR2bpNcMp8fzc9XCVW
v1rm7v+7hMABPAlMHAQhH/QbEaLdkgjTpmM/LqIU8J9H2IyXS4TNA/6SBsLP
OeKgFqZQjGkcKr0RaM7dFxJPdl2FigKzA/HqQGpdVFZV6V6sajeN0rdqpNq7
GsoklCGX2EZbKKtPiFp8HfnHNPo73wu7KsSZU4IHeRB+jP+EMenl74PCqPgt
LMv/Isk47ngqFkQbj5avzR/QvkBp37VsJf2p+GzrqDwpuZ5Z3UxUbOVeFjmt
mVsslJvg2UqPhxL8g9YPTzm23eEspiiTIAjusXC62E8ZwXi6QJJOoYxSGLTl
2Cv/6aVXAdyRbCH59HN4783wHOS5mxlAKL7JWw6a9y/1buNxKCmi9apwdQN8
mkxMqQckYlS7jKOxfxmlDm/cRhizkilmH2XgcrqZJ6RplKKMLip0IMwvcNjF
ZBCExIWXXnijbJiHouk5EbBciuuvLsA8eYs56E6ropqeYkanpxFks+cn4BGT
MfKbxSXvM6+WeNVdquaJu5STim/D3LWzjxHKW9REXJBwwT4iTdFMvPjLQl2u
nNJCrwKgd/lNsB37YjbG8WjST6H0sljB/XrQ+tF4JoiECd0GYP+gVRZKUfnL
tFKBb8wFIl9Y6tACL4zjt6vjHt2A48uOrZzRGaSVvwd1T1IVpVwfJ4WDE//4
+VoO0HzqQk5buDbnizBYhCNf+iOfdjXaXb8rGNpENwbAOdGvePnsD5C3dlej
j+4nGpFYHeQvFgIwfB4GmoiuNJzENPvjafVsdxL7jNQ3A2ZquYzvlEoMtfWp
YTwPCHfU9lf/IeYFtv5cQibUuIfiBUFRUZfIrIKujypM4dMZkI1c+B9w7G8P
4v7JQpCDuXWo1Fubz8y3fYV142qe4y/YUJim4ovaOxtZydUhaVdZClCIucrE
IRi92g5eBSJP17lJNDo+wXwLlGFopbPvF/CQtVxvV+43LJ/3DV8QCUVaZKdB
igBv8vW7gcmvyHlhTrMVKikKFTXIZl+23r0wQX0TmQzPrMyD73aDYJks9+1b
bczW7NAdyi9a8EHMFPN1mAw/enBhAkg3V6JBslTOQbDXZIYRS+OkjYCPnNqq
jf892a3a7OWb9ra0NiLo04vIFg7rLeapTuTe+HTXcbBeuh/c7hhe8mTtux9n
AHSDncTPhe2rV4qxmA5WxBqUKvrwMrrCblPsu9wiZN0xJWUz8v6hkIYhjk8v
DXhIkY5cHG50UYi2WFPbRaOH0p/2IfMvPFAqMIyqT4ayWtBGPvnvVcIsRYUq
Cy7PqhCLmYHZzim267yT2OJZ8C83W71Y4PnwySS6/mnGD36/5XQX3T/MP3a2
NlJCAViVC/O6nT4VQiocQj5KHveoKldgxW1iiTIY8wZ8yio7OfNWHS0kf5hD
JfGwoWfJybpXnSHSC2rrNGouc9XWeeD7M4Voc7XTzA0wdTL8d5LmNdDvQBcx
RMsl8vyE6TQNt2r6VqbTiDRrtdvsQUJL4GCLEf75C0qwVYh2y1n/Qnxfe25V
40Nm1DDkb8S1lMumjjzWoI9YH6gMdg1Sj1Eb3EGQ4MTDSf3ckCgmNwIOBGlo
h0VMrldqCyAyZn2doScFJbG7QNCAzvfmcQAAoB+gE7u34kTvDUBUCEuWf2e6
ayowgeYm7Nv11zr97cc4ivqbrPosHTgMSxOqOljk45cx143+NMwvj6mpNZCB
Mz5F6srUDzstOijLDDfVfpF5O1kZuu1ysXQ/Jau4eht3BKYAo9eSwh0Lk+Lb
SuA+X11HgDoE6+x283rlQFqrTrKZGh2k7eaEqA0OBTP5pQ4tzi+Di1b0yFyO
srHI1Hxu+gXuNXCTgeOkJQ7ty+F9Kix9XU1xISxP17KnE55LHRGR+JTkrVV1
aAmDWBk0rM+8gomUUi5KCDsoLqNwWujUcg9pK6bD5/2PhUJrkr8S0y8dokKw
yXXymjWXnxTFvsmjbIQNMGWT9INd0mCgsEjpLDagUOjD5pVUj7MfqlQ2gI5k
il7NCAgY9//+Kb58RO9pGfsF1rK5EVEESRm45mI4CtUBsXxiLKAwUoziK95P
CkoSPpRkNzFivpuoqhK3RamjpvXm1xJicLomIhEAEjzL6i2PbKR1Py9btQzw
6Z9/9YV5MYSh7JbZ98HSm945HZ5OhNP/A49FoCumumAjjg5cBK9Fd99LgfTM
XBeRaug8n50gmekpGp7YcR6dGPEqkQohK7TLpHqiG67UHhgtBok2/zQKS6SC
VqM87RCZskjKIX3Kyv4WkRCx3UjatSu/AJFcusjgIejvaJjqnmR1a1vc3QOS
EfgtX/OPWXZfFUf8hYS/N/EkY4MgcpfdBvuF2G0kIPjInD5tu1aqnQ/5QOTV
QXkc97hPE0p9yN2srDlBH0hPQk1/J7U1zuOHeFeaoU11HI/DyV+ixauAzso2
EygkujgOZfikWYMEfWxgNZfgIlQmi5KGmV4AM7VlovHDoc1AAKWcpdqWm5Z6
qIaQldQq5DuT+w/Vy6CGam6Mv+fbVQT8WiTN2BCFtva/pwJl/bb5RmuwKrPs
ORo5rHPSjaz2rX8zh0n0OrYYgJiEJR6SP3XqNrX6JI4hmXr5kjJg7AghbeEX
Gfz7KM76oORji33SAHXdOm6qWqiTb/Rp6gl62nfO0pgUf7+1/I/Rb0Ujzzmc
uRXpA/rYU2lkxq9y4r/xepCdqsw6rFW9ObX8iQt0FOsxdxn5pTB5P5gmbKHe
0W/0KD8a1xIWdTRwgwym8D0NdGgNg4n/G9bh/5LPSbFRAFYKNT4H3qsHdueD
iNoR5cOjjm8zwpGnZ6X/WNyLfiyTJ23fqSskvCI4hwO94p84jAh3HW9eSdOl
zjo78h85T1N8IF/Jq1sr1Ex8LFvXm6+37e8RjkQiDuETSkZ0ISgivnk8uFp5
AIt+e4li4IMEC27ydBrUw9nf1NZ9SGCCO6osOVMtqLyZn5Yb3NUeYMIvg7mf
h0Clm/E/YoCRt6V4j7/XzPGEc35HzW15MVtSgRdrqx9k38xy0xqE4/f8aCd4
fiE4FEaiHxhJUCW0zHWg3z9pcVCR6heD1eepw0cxSu+5ZbPI8svAxXQK15yB
CIbFD9IzPUkh1x2tMYSjgPXlIdD0WBQ5T/jEaH+m46Xqgk+LeMtNlIR1uqe/
3+F+b4SrNV/pQV+zGmuE9WSIridzgT07MRI/wZ/JBLarLI6zSomuvhWHG5a+
k1LEpI8h4eCmqg8pHMHcisMEPtylTYBg30wfzXPv9WR1a5ZwlMn5rPuUfoM0
ZNPuLWiRgcyOvHGHN5pw15u1tFrihjjD1RWpmupaaQZuauyYVsx8CTIIFVPr
x8ue038px0OjqJQUW/mu5cSqLNeYz0w5mD6PJiWnvIqPzUYg1ndN7FCqSd4O
tpT7v2R3A5J/FMqYI9oYGGRcRRiHkV69V0xzwHbds3RmSbWJsfCWJa2b46Ov
qBpfKbl9ye8/+zjVLM5kY9EN+1bPqWcEljPGqzLJttCKBXrLUcH1EcYwjhz+
hz3GNpLV9h6wfxgcuN1srI2hZq0Evr4um5htb0svnGNIIsTF2/yYFR8LTITR
/BDStgjPtErlR60TuSNmqlxpCuA8PT4OlmSrj0eRVyktrSxLd4GiphYcd9ql
9PZqOUHFMURmFAO5IhK5bHK1842IMsMqWidYs7aZrpNJi7EL7Z8+BjpoMR9q
JmumqQKECztuBjvdWbG7JxPS85/PWbvP5HNF0ht4LJwu6Lw45vM7j5Xvo/0n
xzPwivWet21Nzu1ZIykVX7KdEciFBJCM59KypvG0Q64ygh7WTCVasDCAUzSX
11Ugig17XFMXuC+CLdi6yFjgkp8GC1tsmq4+c19vbkgP02W2ys5vYbdolo2r
Pre3yUVd9AdjCb/t6R8r0wDzlv+jX0JrSTihlyYIWaOwOCqg7YkW7NX4q5iT
TADrHoALDmijL3YSH+xqc5p7UiYiQA13bCz/tQ0jiE2YVPfqA/Xw23wwc0xw
Y0mGvgbVBkpNsh/RTcAv7WyZybezAD7Ag5snzmYYnQ7mnCCAfXXG/odOqYH2
udo4MU4etyrfkmSqdu8jZJSx87LLIDeh8d5YCT2VTIEK9HnlxnG5ODMD8r2L
mcwu0GxKRagiXf+neNC4apK+SFCj2Hub9d4ud7Y+jX3M04sIV+54mD/UlCcy
/DlPdUn46YMTk3FlYUZbnE6MYYLkh/022AI6DJE/vNEyyPNG7pxI8ek+tOpj
iiIUhx1PAI+imWpoyphxHdXXDFaBiCpJkZ2y/UcU9N/ezviDZe3IzRuRW80u
VQdIoK0G9/9GreLyqQslwM+HqZ6zALZz7d1memj1lUlU5I5m5Tsk+gAPMSro
5LghYsYfQfKA/HbFMup3dkuemcglGmMHWg6LAfyJPY/eS9JU1r/PM4CCHuke
KSS0UZ8fxauXuQd2ucJWBMBQ2Dm62SS7ohOtcHjYqP5MZY89y3Ye7ONW/a2k
w2pUqVeYOHH/xqW192NKliQcvglSBTGyF5/dTCCmrb5mWNR74ARFmnmoiBNS
brx9/2sUPF6Osz2YV0RO2Np7mM7Q3mske2CKVBVO0OdnEpTAJvWBRNJC6Bsy
+qkMrAJjUVhy7Q6zgi7lx9re3it5tBSsFcTuiL/viaHdwuNaPo+2GwgttLrH
xGdjwmwWCw6u7A1qGOUp98dBT6jeY0xB1DQ+I7S60vc3oQ1gSHw2pEfH0Vc9
iAhjfowOrtI1rLce+vuhlNKFCp2JPuKsnjvn9CKJ1XdIvrPhJcHuz/2LA38u
MbqN8n7qvBOOWZeYJmL4UhQ3SGhQ33Fea8NPwcBLvwyooKvsjNtYrBr+uVnW
O+HOI1DO/k6ADSUUu735OPe24GXHeJf2BKyZ4DkypqSOy7knlUHWgIqhYG3H
FQRl+ZDgpWM3146/iuRxIBUS5XjFrjoPFA8LQSPABcYHarl5z4B2LbLzoDWj
ReYP4TiP4K1GnwoxRQJs20yMB/fc8zjoZzcogTy7hPkCRVu1gcgjnH9mMcCg
Hd5dSd6OQ/5E2sgT+U7XS3bhOmMaPXWCihvp41uzfjKEpzOLffOqRocl7pha
y0AaLKSvhjOnvXeeM4sFdpMjDurLCHG3abYPSsxOGPwltOstVMlfxYyy/1RH
+/1LqtxC6yPJ5iI0SDzsQskY5huaL4ugpmWgO+1i0MrdhssYRMaFVtB0RY64
B+VgXVx+0t3uV1gw2s4+v1H1f/GBWxByWgKvUcqDy36T0N953k2JD2IIXsLW
6NRwEjzmpRPsXcih1LxUGoypubpajLI+1IkKw6BoLusz6ucZh5zk7C1kNflH
vmBgac57zRq3SPw6j1G0w/SLC6Hh6NGMj274XvxOfWedqE31Y2W3UaFGbOc+
DZKC8OxCjz+VlJbSYzW7Jy54+QVRcRk6AR8SAEoM+3w4zWSEVqJu5XdRMgft
ntT6QIZMfdUUfXGHo6jVKwwfV8sFvphwoYWxon0UO+9o0juxqPz6UopuxiMR
en6bSCgzyyuEsux83CBWIOv+rqSn2pFApzGrLwOjM8RLNcVPvvUIwlNGFY1J
JpX0qnJx4oaF6qktpEkWOKQMfncxVJjjCjwEg54NeK4dyVu/HI90lZr2OmK1
vdWZGJyB5QOyIs2BGnyCkDBIa4+dw7Fh5i49SxiQNLHe+3K5mkqV2NaofWvp
tNEipnznE0sfqXy2ZzGGgi011XWL94w0nPNHGDKe4AgQo02uJy03KbA6x0LV
5CM1r4TEbci6FxmKBRfNXlR/+xiWz/XRkPztdqzKIyQgEtj5lR4H60+q1QEh
t+Tjk82e62JVJjIsOebaqWWaAgQ7pE6/WUETcAsCxBIV4pxrdFZyjTCe9QVD
CAp5T2xTZFEyQOE7sOzRK+fbQQiexHPBTzf2goeMXGEfG2GFEcmlYALwYq3r
7m1HEedoVrPuGe9bXgwhnk4lPMMlKAKimrNs5KvEAJgKOtYqGPOo31QgtmD8
auY2fJ35zFVLvS6xLrNSWgwVFedLZJ1OhwEAycu6hDeB+S7wfHz89lyr9UXq
mFVzoQVjsb7/HBHy7UxZaeiUBVDWCNxcspBOQjfqktEB13Sujy1pm6jN5hzQ
QNZbc+pLs8TV1J1d2qqSe7dFZU8rg9kPH38kA+waQq8JPh5yP8RGKIiXLFCB
9mEsPYkWLfFNLYbOw+hnj/mQhyhBU/e2rPPfLyNSJKtBxrAqNryZuXRdK/Jr
OpRIeZQQpjK/xo766dTbRy+HD+YABNprShbv7CeNjIoTec4l20ROqgvp8od9
lS+qewFL3Ev989KPs8k7xZ34yEguH/jZiza3Ia+yoPq6PxomE6OtGMYF6Xk7
3EDMEsbwhLJ/8iaRBRwD8Vd7Vwa2NS+HjtoOQEkeQFsf4mEvhzzw7p9sBaNP
vp2DiqIwfMzbjtbaTlFp3Uu3bNqvyW3hwk75rq6UhYJuptiZg54f2vsMbrzR
gkBA41pXz73vxjJ4W/rjk1PaZc0MiGQK4J0aw6Xnl1JXrHpZv5cMdGsbtHpU
0sol+u7zExTX+VDoF437SfdPuHIhR63/pRGQM9pfg5L4Y0Aelmo9LzpakTgP
F4tn9zTwC3CA0CcUTr8Xq5qJzR6TBYmk7LV6eFu3JnlNogJFhKLpIOJWM60y
R27wCqqdDPcOMkip4aw5ICmwrFV+kKZwnTyEPbxW8EKifquKrONGCP9+yDyz
to50qU9T4z9TVkCKFKIJrcNOTvjDkBvJlR11v4YDUqU4B/t4HP0XU1P8Phcd
34CjQIOhjuyWSFVIQHhK5tq/g9kld6YgO5b+j97f4kkA8qRLYsBhY+LHdVRZ
RL9NeeJRnIWEv1pe3xneithTFvcuSb6jgkLjcbXvz0+JVEHcP6dfcLHROU7Q
WuY6Mbww3KG3mWwAZeAvgag/Oy6tVnk6ksPYkTqqkiXgY0AAqbyGCEn04/GV
QJ6GyxKU5hBwNNswMmuV+7UbTJ0VkJJIzzAXm+YQuytP4ZXxJ573BJTAYDZ2
F/cktDOgwe6xC8HvfQ/5yiT0Lqw0VOpUhconO0Ucuz28QyxmD4TH3Y0SMMk8
rftMhwOV9Al67mDI/Fl+3yvJB2PKD/O8Ai7m++n2LOpnzSCUR/CYDBwlD8wo
qhmh4L8+sSJRui4/L4tCVwGkiJuonGL2IzzrWPiiFGFRqBAEhx/UvyZiYC9Y
5MKjNq1izBUrLAD4nWTIL1H3lrBC9gZp2bHJchSYWzfLG2CQtHuO36ojzIZl
5fxUYZ59eAccFcb4l+vMKwom1FTkJHZBCPALCppu6Gr0+o5g7MVJRg9uQkk5
jJYx3vxCjw2D7jgRD9dTmZsGE/rtrhAuok9pCHtR6n6iBElqn4PLl0o97uRe
gK0UFWzK9EYeLBhEnz0/ndXE91S+6At3e/ZN8/YfYDFSKAKyiajH+3RYFBd4
vyxJVzrkv5FPi0L2LhTPBfI8lVqgmu0kIp4QjXyeWRmB19Ipdk6hZWqgzm+H
iAQXYQWnrS2AnWdOCahIvsg5ef6odScG3qJL20V7aj4EJMaMOw2GrZzJ0VM0
B36FdGX/9JSE4NcQvQ87mWEo2BlwI+uyHJQhqpvY6rfXWHhaVh0ij6uXVSPM
9qhxo56ppHrMOfZ5ElFNeew9f4HNe7HtM68giTgdkrL88Ph6DcYQFJAXyH2b
sDlsYx26CdffK0TpuYqzNYofTaLl8HevlEBwtqxFXt2B/JPVRLsxO+LqDR0O
Xi43RQ/BQuC6EyJIjXTzI2uzNBXT2pW+D3SxiiMQBRp1ao4MfZuOFBG6lIA+
SI0adbSW5EXOr3rVHWYpfT6q9T6CqDoR0upJX+azsrRK3RYMbTl+5z9+5ur4
afXfGogEAaala8ogLlAm6UhdB3vozXqG8irYPXzTpqqFkimbtpc7R5Jc9wYS
v6o5EDlubvOLA96/vISgtH/C2bdrEXuACgkzrgqvgyDA7BnrMvIt9eYz4P5c
3DkV2GD5YhHLdiZZoxNPF6CWSpF81XA2kAzZUczk3WrOmBf58Oyt62M/ZLI7
ofcTskdehPotvYO0xs2dmDnrPQGmlvbJ1QHPu8kqhOQMYxbDwT8cwJYQ+ESM
ZD5jz427XWBQs8nt280u1TxpQfDbpRYtCyD7SJNNwUpHso9TVKYvyBYUx0d4
WINcZE5dBlsihKKZiBhEdzdoyySRHyFAI4ZYDJVa4e221uYTpkB3vlAxZ/cn
EYrqqCb74VMVks4VO0YpiCBXrjW6ibbAUrS29LzyhKXAW9f9/Kf0q6n4C+Cm
uZl0DlaEMXd0xuzLsSLM0grNEexiCVYaQArQtF+MR93b+px01J473NAvndaR
DxebQR3eAsZ5JZNi3hYfimzcObRX6qHhbKeqrY5SxsZYPdo352xH+Z2dBP8a
5Kfcsc1vlUfVlBoOIqLb1PmAvFkl4XIhWVBKPFnv72Oq9lR3FMBd0m7dGH39
rHzJWgijBkChJB+rJ6BAG/zrCR1/a7neJHndCRmzpR+agKYTGc4fp/4fF0+2
oWbSkJNUzYGNORS6Sf18HTl2iZ/PcFd9mFYazlEXbqcJkdJKBTCX4XbA57A3
4meNsWzhkDV/uAQXsXmq6k3KdmnKKM9zlLN9nhx+Jj/+V6kS34aXL/uGchbu
qo9DTwZJoekiezc37BWGp0ywn/IpPQLYTpR/IdXcOkR06ZUXQ9arByQWHWGW
8YmkTWBLsWKNYUlW2Oy2/MEskQobNY5Wcy5UE+LPzkPF4Lc90fsEa/3VcFe4
3zYn68VSimtl/0ydy2d9AKn5UFhrI2LrET/UXQNyf2KVbUisxdwouYUYrQ3K
lAx1etdEVD4f6zMzAD1Pp/t2TPRt/UERPXSPR7YIgStznIymHIeKz1x2ZWN4
LDSUSDE5XnkIfhwaxsLDZYtADRf9g74B+8541S66EKwFcDtpC1Kn57IqXtUQ
yFAwHbw4WLKp6WU2BvOjWJk+nRhD0SbvwOVfl/kzJ4uO1fLoWxd1Ek89Z4mc
vlqdSKJ0APbp5L12nzF3XaQVQWTJs31UT8X7DJeMD9KSnGU+K5iyHagQHDLn
lMLfUI1o5zvIDavHOHDp9vZoBO87QBUVn+mBQNIFf3R+/J4HW56yOwu28vYJ
Q/02X2yU6YHnDPOsjk7IBhkjd8F76PGGOdaBR5/39+9txQB3IpZfKBY84INq
Cjsj8Qvc5kFCunaSUeJCkKKjcij37n860aIiSa8CLdBi4K6HgVA/RPZ65NHU
gaZMUWtFE1St6Rcx2u8QR1an4slB79OARLbNsaAdaB2haAFnZrfo3/ukJGuo
3QiNJkOG/ytsQD5qllmkDgt4EDU6UwbAAV0CZVNuWFsc6WMILrl0MQEODl0w
7oRJS3sqoth/zUUNHApb4b+rk5Sox9Kj7a+QMp/NyQKdyyHoOXbVy7UHQ8XU
DIYb/wbUhGsuhTblbwBdf7RVXlK2ajnjrzzzSaAnBrnOWseM5mLM9GNPAahm
tOrGJo1thEpJkeIzVXfbbqwazdUUQmZmSAOv/sJZzJE2TanO/2G619SdhOYO
LOzyssKw7mtQT2UTrElk6QuDOb3t/UL/RGXOhOAQ0bJDNt8bk5We2nAmcBTb
5V+8ptblDAQTDuOMZMr+jevmFplce6rGzdrg3VvBTJIfy6nr1WP18ptEQOc1
YzkoQzwoFlM8L5AGh4kiP+yBEcW8naXhdFnSAbpOk6cuzWVLxCTNJeZfJF/p
wQFHmgwxqtt5hkeABA/R6yigD2uK79bKqXWURrtj9vJTeL+aB+82q5GUvJ/O
kXwWy3hYZAJ/BtPiC8hBaXCUGuEOjzcTMqQnxAKh/+dkMPhXuAmf/npGJaUK
hHrE31vZCWPZFy7oNdpq+RFMeWMKrcEDf5dFwnrnWeZ3rFEDDr61Ua70ZoYD
SJhRf0QZ0uRsqaBcDIYhUzZeG6kJGR+f7K5x9iV3PpOP03RScJH0VdAPuQER
ImCNDP4+Hgi4ciQrt97RGCk1kLjUxJ+QB+Wl73ZTEl9ysAwegKAKU2pYLBF3
AQ6aulCIKUXq5B47qIjg04qtfVIOdvyGlLpyF0/IsFwGWfguWwqUIOhsbCyZ
Znkgr0gfXsgj1vubBwTvTdvt9do7MBfOGIsoPyLmhhYvg8lhj43EDtC2xUbN
hdQrSqPC/Q2P8XSKiORR90HWqMqw6i5SZZgIAwXIm7XAEGzXin9ILCk14dcB
g2+D0n2F3oompfEb6xsW5Py+BHup1s7lR4jUOMO/em19+kWIbI+eqDC4cC5j
bj9OtJMaVwMbt2mAn6oRkrTNcerwFZff2LQuQ64S6bRDuyPKZBSRRXAUWNUZ
nMfxXrQrlQn+LjGDw4Ce4eh71J7xBjY7YXwmWx0HPJd2D87xZmJ7NcJ4xcE4
fNqc3D9A68EA8x2Xwm5qTDaeZU2Bynz72uIxMJRaV0Qb63++ZN5waqDCkgb7
774OUmG0lCu8z3C8GqUdXdO4wHMsfs9YDATD5vNhhWpShemHy/SNFmxAtrmO
AXL558YsKMoSHrrx9eSTkjb2+1+KJ4rH7rB4gO7ILftYRrFoWDK1SFfIoCMd
6ZfqrhYjjiIa79do91UyGPQQB1NWow1wg28m+4wx4CtjYvbZeg6tdokdGSvF
XrKc8FLoetc7jiZUG/ocEyfFHic/6R8Kr1e+52icgJrh7Wcc8RXiyM3Yh2Gl
r9Ri7alyZ+hRqfXABxDTOE1Vu2syJ4Ae4I04av7pd1eIO9Kj8gNDUp9Rl3a8
Ru/RPR6sYVDSL32x3dIep64eqmH5wTini8BpPrqjeOOSqrXxBxw+iX3xnPek
5asO+k1vUmdZrs5blJYcQdkO8vMstMQxxowKD8dU1XKOg8OYDI8UyH2drJ92
dC+H9MEA1/obuOT/OHPK/i9WhFxmGOVYg5z15QplM9m+Ac40G0K0mb0ViSSy
Jz1xYnobvNGZzDSHE1282HZc+Ozc7SWlAfW0DuF9G/nvAgQU/4lQrEuYquOr
Xg8hpVABmaqJ8cL/wIEPhWrn6UYCl05iLd0WAYB1yvLEFEwtLxW6xykTxRLC
oiCtS1EFy6DxuufpqaPmXA/noG1Ufg9LdWevfDlnD17DxOcVXJGL/Cl7rtjF
pURexA077AnGMcnBtLsvQGCkt/gW7BEsG3TPqEbE0d6p+GwtfTdgHaYBhk9B
DjjSlI7ryACMnYiV/4+99d7a/QXtTyAYQCV7wHUupoNnc7jSJVSR1T4Hq1K1
9e0drStBBg6cWgP1XhtOK7mb4BzRSJgFjQLwI114tCpuAL6PCRYwOmP3jFZ3
dlfHSLAxZUXEkird/t6u1K5Q+/8/FVzJ7xJlluoE/lMlKp6IPCFf2ZK6/aVo
bmdo8OaX+mtkO1IbZOJ7X8jLp8rPN9A7cQG0uHg2KyEj11rZ+a4BrXVPpC8L
9C9eutAjRywm2ZW5saztRor7QmgKJBejzdB1p4qOBkUcmPVku7G/I1qXkUvb
yEoENx1qZXPzjSJzj+MSGeJAySr+PmO0KAiIQaQ5SOdQdM9ejQ196ColL6F1
Jro8wwbusWIVNpc78IuE0cAXXufu++aWNAZV9mgfPUlY2id3J8s2/COQL4PF
NZvwm+vYHi1VPku78zuIJylz3eACU9loIKSG59Fbn1vjDKe+vcD79InW6/gb
KXWUJS/i4DDB0weAiLT+HvO2lat+OzZKko+WoTOl3xoiY/i+HrZK9rY/fa+a
XR5BzIqPw0CPwMw8OWcWN6KZdnD71kZY83epxXPb2Kfi6KYhwUu77o4iTnA2
vUp/Hk66o+lQfnKi/uqKmTA7GF1gctSwCoa/Oun0pNf0oIa3pWahW9AvBXV9
A9c+PjpLzl54EZkHVYP/UFk4jXZLLjdEucm3c3m7PE9/qCfCEZiARFf7/UBu
GrrYFPmSrsWY1RSqy9sh5/3vmVbFow8a2FOLigCm9ZB9UiMZbnWois7p+8Hu
FNmAJcPWF4xecHyVDf03V5UlQRJGBqht4GxJfvuW2CPG2F//ela6Ssj3KlaZ
SHPXX3Gejv4MS36ZuPa4Wrrasnr1IntRmLwBAAIfVGFrh7wIfXU00xgoNLSN
KKjb9Gli5IZUXezuBGGhXVUIzp7X8k3q7MZIrTIdD8rB7Z5RrORf0yx/R0ln
1T77KHX6zT4uiRUYW3Q07x6ACtYsb2dn1/M+YEB8p3dwzjzgMsBiCLzL7dg6
Kfu5u8m0WK0wu6jLQvNKH6YtGCha2QdpwEHQZi+SzKzHugOUP8YvgOZdLtT8
/TEkUOoLLkQsgdyof4T8JdRphDvtthU7VNWhTwwLiNZNiyi1RNOEpjljgLiw
m7NMgXe89GZa1bzQgnH7F8xmdoNmmdMetRXOkFnZVUxDYS5WC3fbbW7BZ2eV
cpJLEyQsLSs+JlQxtXznatX/1zeNNd6VDhc9AhIzEJfLQ8xA9hmPIom6tLGS
rk7StH3ugJcgY7kYgE8jJoZHWpNj/7m4HV04TtlXhuIwq8rrO5GrB94KUKir
A9jHSUy4EQkF7SmRiZgQBM8O9Ecr3PStIZvOWA63hVNHiHTIZs+xujMazhJU
JcChuZvnCpJmGMrESgu+/YkwJYMDBy572qC78DCgcuRberrZhhBqSSdpTGYb
O6mDPIkRH4a3lsTq+ZLMIKwA6gBE9U63doEqXJiTmNk/xfIoWg/b0kwu2HvK
/xiTl40msiPD7MuI2VXeb2u4WTnOAJNNd6P68xZVzszlXvyHLZwSSGe1kYyy
ZpQakqrhto92NWUOkWMtf1wpVqenJUvxHaLOP1eP1VkNJuUFOZ2H8oQKIxuv
efBZ4Ys+AcErV1Me/iQTP+1V3MQmoC/KDK4xfRMgEkaxtu9qkwCIh1Ydbcrs
BFp2GWKmP18d1c1Ld73kUaCMi5rGRDzAMa21iHrtxhRg1NAbRsnwvxmVr2bv
eC3VjhgHfRD0GLdlVFyshUWYSm4/8fPBfp8wjTOV4d7JrLe0tvGAMDnPZgrh
HvBYdTF6vV2CDDuiJsr7AV7HB/V3aD67G08SwZma4tOsjhpgXKlKhRdZCmHn
IFARai9J5G699QDh636N2LEy5Ttv2L4VBf8ezVIZIVCoFHTRfTtEyGGfDMWC
J8tXWUSmsIXNSFt6aFaYYaA/z6fKK41QNGv+zxQ0IQ6GdCe7IXTMCAwk29ys
KpWplRzhUbOcOFOqj4i5EbiV1fu3DVAX6M3eCz0x3EuqJOp5RZGQzYaP4dqw
N1GtX4Xu8u0K7S7nlhI/L0SLRbL2U7wteCKYnSokq1Gmr39CoKCw3JmOT009
Mvanzcz0oJmjTNfLuBK8Cgx3BqnKwh+QYCJVOV1dsI2cET8t3LX627DPr46T
OSa9L0iTeYxELsYavErbVrny+Up2d+pFocOug9tN+MFrpzYqy50bk2o792P9
6s6GpgXM+XdJDHURI4vrgIcFiVkaA7W+v89uuduEf4ImXRpzHeWWp0spQoYg
KJN+vZbKAEBazOaDfIoI141Hg/Lg9BUrQR8nMlDVrvBLG+cuDF4kLJZojhCQ
AROqJMoKIgNpGcuzwKSfzWdG+yUrv1faLdPSu9JBJYkXcykYyIWFpBaystGO
q1KqBpChXKR06KmK9I77n4fXjbhz6yPGrRfBjIPrLApzOKpvrK4n5sDRl7p6
3kxvgTL4GRuC4C5gzmKXS6xBKDMewPnmwdz9AYKLLMxQUoMgycFGvg9oLsW5
uiv3b7qMINLOFmexoO4ZzJSxjQ4DdhxPp+3jhYuy297c6PZVs35fLsJND8ge
w1Qo4hUr3Joep7A5Yz/T+H23vJEbOWS7zpbNpFzucwZDzvjL4WT42Npw2jkY
PJxk+qhLD1kzzkMAIHLeYRmriWps9uzR9w8wcuWdxC9dhT9RQIpDTWJvlyon
WySAJB6/MxXBfPU9fAa8msBf537zNyfb6/PwqRNJuSkkbLJ3TlREPqhvAtFP
LGKp7OH8jEGxEpOWc7btxw1gPRWjWtuxLPLzTbpbdlyyyyB2b/UTGp82IO6C
wB4jFZigJ5oGvy441Mn2Xs0qHrJs7Q1qBp6bwe7u4l8DJ74ONxskxJKOoKo4
Ex/54HzScsNlY3XIjEZdAab7JbUGKdDFhnrfv0oBsJhvh1R5ZmLffFaLpchX
BE6pN3bOyd5wuxnuTMrhcTXNKr4uQRJblKZ+F2ps0+GGwnV/SizgvCNR2vx+
k2UoS2voQqMy36acDvQ6uRD6mJXEZdhqScdMjSwwnucA8KzG1nDIMEYc1mqk
gq3kOoIri3Es4Ek+/IdI6KBP+sD1E8u+LvfWsxKT7fgp6Ntren2WT7SPifnr
/fzLe/Imx9WNSxJIg1whTBbIugjnAQfgMLXaOMYk4i9zSy/fZPCOOVDUIpJK
wo3mMySKRbv4/oWMm2p+qX0BiDyM+Eo5m6dxKgzcfvMPcOCN226PMl2HqZuw
OeM4IMiS5u3jx+flur66MhOU5ZyikkaayzfBLy2i7uQBhCN0nmKW5sy4oxPY
aC49VeTltzGgTZH7BEZ95XPqUea358E3D/kMJfnXVP87/VYvuIF0FPQ1nA1U
vCgxdJ92ZaB7gfyfQSLxewGSippxeGdCzfYYtLdq+Wu9L33puOC4frVW0hBq
2HmwbvJz+u4SMRHSh1vdyenXdo1K2uGJs0J2F7zi50RRGRJfuB2a+/IW06Dy
4BwOPN4Les1Dp5Q4q6JQ3wqRegNqTaAQ8EMbY0fLBfY9+7fJ3edC9kO6YTFs
DdsTjCgjzJgPS93T68kdhk/fdOs5P1C4p3YdIFxU/XPNKmVOuEAyL744yKLA
3bZfuk24cnLi/duS3Eaj2urr1jY7/G0gv6uxSxA5BM6RCUI1Vi0rKCBkrkij
VQqF5PyA2hh8ZC/23IqOpYBTFUeoTGdOSWA0bRedZEBvbEG96bY1RljgIaPe
pOCBaf/zdR59l8gTBZ338FNjD9C9xZHmyGh2rzw708zr/dE115JbBFGLDnN7
u211pUxfdYPSU8xSdtuYfYo3vcpGdQmRLYaMCXKEJFZWE24KygYFE92iZlm8
9OVlOeGnFjsj6ugrFH1Zai5SY/jqTYa/H9dESBjI3bw4VVTMu1KxpIICM/fN
waKgV2IsIZHZgGbIx2ahMmRtGncMKZfabQIbSL9l9a9mVszaVnsnFj3oAhJ5
XTXy/yPhB6NDOFxO1HWPnIrEngHPrOBwHdlzWauM34sCWhWzv8ml4GVVmWL6
B6eI3LbgcS/JxBeiIdVFhX9Nzx4fKoyz6sCQiI9MQtafWJiklIjVKjatJQAv
Ptu42sjjg9WKUNsIFV5QXEg8sL1nQRQapey8aMDGtxOukuKDyXuMWZrUQLIT
obkhs9aTFrignFIbhECxSprjBuXFZ553kU/UzM+d0wjpdAUwxiE96EQURGYW
FthKcHnsHN9M55CC4xUZLSfBWtLQTZ5fVmXUD1WJUO8FtwTORE6ag+NbL3ke
qTG7HVmcgpBfmVMwOEcB2MA3L05xXMnTAgtATkbcNRb8Ohlm3q+asv6L+qXw
1shbnaSRPD/7l1WRJHyqKDUA7JdMz9Vgfmf2T3C4d9Jn24iBVCLD8DIoc8Ji
SCkih/XEA0IhrrMFKJ0qoqTQ3FKya21MSB1bdN+oEE9vD75rp/mTf38SBOMN
eAWuXVcyPtqlanMH+dIDFRGYw3AEgsG3h+uMzRPS25dALr+1x31c0Xdd0LKg
dNU5uwzhzDnystaKViq3KX7bseamEnuRSECz7dHLCuW70PwkDJnpmAWZDlSJ
VdUfGer4VVjxccuAjITaaBgD3dPtyObP6PaFMt+aVjA/ECCzjcoXejSwta62
bByg8vgJ5LkTBt2A+1WCRNJhcgciC5jlUnzj46zn+84J0LpAX7ONJ3aEpi9L
Hvwodf97TusOd3NSG9QT+1o52TBt7v5Zn9gElUESLZQksKPykwqbhHYrmZ4F
cpEOoXzPl8K4rNllg3IN1E2z2tVY9zUta4wW/6o8wKwJnymt9+KUpVH7nXeO
t6wZesDrOEZKwH0piEaHob9lCJG7MZauP2ATRqEqHN8i8c0SNbcE4xPRiKvj
HJS1HmeNsaIR8BKN7ERgpuZgrU9Uhe46Krn/1RIF4PUPHL+k2OiJWpmvU29j
3ZP+nvTSvqzmKZ2s3prbI94xFv8hw9BkmsnE9xmpUWY1/TksU3jSvmqI7wuJ
y/Zm0Yi3eQmiheIIBGodtqcYzeSrEZevYp0Lzct1+crq4Mm+uNgd/2zKLNng
rQ0kbRfxKYLD0XAC4nHecfFJ6GSVkexQkj7oKKZIsZPVeITgl99ed46lK7oZ
3GTSiO4taPJlcC7m2cRgwAMt4CTRwOHMnE7/d82AYfp9lbSdbQz+X9wkVQO+
dxqYy/CtcntWx4QnsJiFszzdG8pxLZTmioiD+qyHFGoVa3c0cbxQOb0RwTOT
j9rQpA3ulce7ipFmo8FSmh5CYdfdvdBHJJZdrd95s7ahISUwWglDb5OMCHQM
N0vPerRZ4qa+fxinjX1t/Aw1zaxf208yRfiro29LcG4Q317Bui8Pq8++ewAj
z4wJ1Jeo1/+LiPakcP2Bd9D56+GL8cISvrE4EC2LkcP6HwA4iJdnYVbxnkyk
+5a11kaSYr3fLfIA00x58SUExYAyw0LYy9UwhYcOsYryqV2M/GDTMeFJCxf/
+nnQ4wmF+jlvRDx99pKTCMW2/V97bymZYrc+qjSX6tE06/WGqHpe91oisaPI
UHaL8FGLI41t995/MMeqJ2hoMyhbv4nK8uxQzdjBfqNlWHAyIZQM3BL3JmJi
6FXY2x30ELf9DTXeaaas8TjhLOtuEcJa41ydLHhVr3SoBXGmlwl6IFZlaoMw
wVYtTejCB9cPFVjkmFD0V7A6+X1WSOU2mif1dh2TobftzAbZ8MgfqC1UlU0y
y+lliv5gzphB87i4Ao7kuSYeObNsxABp+QR5c6LkDWzXy4jnao0HKirDXSTX
ecuBr1TAH6T/9hFu7iPiY414XaUlwHa6QuVbJl0vR9f7rv5s+8NUs8WxTSnV
B8GgopIvld+rsIvXAxYdnBok6mEMEUx0EkLkECNESUzxhWJfvH9v5Qs50C57
ZFKdtWW0/uWzt0eRSG0aLB6wSXeBq+uUF8gWD7CR+SuxghEj4O2Tq10hXQY6
JP+GLVMeRcuygFg+Zgszook9W4+lh8Yk/XpJE5MI9VInvMkdfsFGu0DjuzkX
uCJfweO714TxVnQaAwtnF+zvG2hQZ/tW+XTrJlZVw+2VQz6SA9Y6zCafG/Zo
gvfS1I39bAdc45Y7uClZF1A/yNNP+W1bYcz6iGGifyEKikdeBqfWYVQwhceS
geXLxLTgBquQkIMIF2qUdm+MkZ3cJorXxLVaTlT/7iMKIdGw4ND+s+Ny8lgh
cRpegyn+4W6MObstxySdNakYMLbiu4g22hlxZVFhft8DosRRerPGblbev8A8
puzwwH/AoUrtlP2myuZADStmX6GBK32ZPx76DO1JuQlPH0BlPHULy2lXgZgP
IpBfjDd76xA33xpHhie2HlLP43tnDCfkctz+IVmJcQ8Ml4mHlFCppUgp9qaT
mmuHOfIw60SRiIJ7lSAQG0dVEhJ0242ASvO8AbdtoPQfIKyQu0shtlAcNadg
JnwEpbrRFCKNbclXMTvQa6igs4vgXtGBC19lIhoR+oxiQetl7hbOjTdiRwtL
RuYurPSfPnMWfzdWKzPMVjrU+R6pqzymuhxZ7rvj4iY4KHZ3K/biDTKqS1Ni
gxo+czhPmnJb6ScmDDKSYl0cZ1dPsiJVc4/8B/rCZGC0DoPgaYMfQ3N8xxKY
qC5yJMpKLxu0t2jv0NjoCjnyc9zHFLiWYqxPaNYJ4lUECOEUxmjNNH5eauYX
TJp8S1R8qmJVbKFA69VC2GK7flLVHCZvQ3s5POQMxNnRiDxNccdq5qLlRA6h
Gs+GSPFqKZG65SZLHLD51WEUQzwaS40pjGChJs7j8uGkRGAka4zdh1YEY2he
j4K9dgFwWG/6/CihSeGSwqO/twcyPGmja5ELFFDJWgY6k+8CVdWLSc9f2h/I
6SAUAWmNCnjcEX4sQZVSZPGpCUMwSlNt9xUcMD9Yl6aDGOkPxObSW0owwX6M
WurKB0pg+xiPk+eRvEUYxK78t9llcSXblrpfbrQ3BWOoGt2Hq+Dbg8AWREGZ
LN+4HYoV8bTKKrg4HDNWmJU+V/CxCYH4RUT/wmhh4I7QQ0VQgS90BSXSDtZK
IiuQcKOa7fJmCb879fBNGT+n4sAEfybr2TqQOfpNRKRrVaFA88ferXCeccKZ
kXmsMYEI+aoVbTK2Md6gbDyDoigC358KFw0TTibsvcK6+CHt4n6grV1yTS/T
kiSGwsFa66FbxR2mpfp7vxn/J/TzaFuT8bVOlJoGlkXfF4f7fcGwxJqYSqkk
Qc1e2s1JGQT3i+i7zmKlzzg+uonu2z9nEykmk4kEOhJnIo3K+uOIlVPj74lY
/QZ8zLdLQnhe4z3k2GdJDAqseQ5VpFCBm48j3iXHdZ4GLhLiNeURSuEcvbJD
v7rV/3E4aAY1+TFC5zGaEIr/IbOCQw+HLMhNOF3K9ObfjjqbuFDoHhKiJ5JC
b25ltt/rXw4gJz/JlcSzxZITL3Wb5AeboMxMLpznAtbY9KTDdZRBiUJB4Gk/
7sjbcAIwsaJ/Esdh8ldDeS9Lzpu7Q4ZKLuF0MnRS0wjgPmhIKKVlVrXH1oJw
6bdC582mPU851CflOdvVGr/RfOMrGZuDrON9tMYJX00XX1DJ8fd+AEk/R93K
DMepHVnO2P068aw2yU82qGDvxRY96FjRK6ShySAaBoEYi8eFqLbtYCJIAlAI
RVPjgX3+UZduAYyHiUy50OKCA+zOVOACyuhZ80nrwzjUpjx75zGs6yaK79GY
l4c1vfBqkS6UHKblNskMafldPXMo9PaTLiPsOrq5NLBGySZAsOn0IxWIlde3
U0ZWNcEj310jH8IAGkEl/NSbTl5CsXEXteW2LtvoLnxPyqt/qvxzPfCqQtia
RLr1cZwd8kXPsLZPMVADAESOLI0CxMJ1HgzW4aN9e0coxQeCJdpeIN3mXRPG
e9cHKLtS6eMGmqI6nXq5uwIq5t5Kd0SdH6FESeoOb2EQhHvnIRpGGG2C2VUX
fu8VqAY23rjQ9hRGCHu+D3bzScaGCxCYD37z9PysamOG3ESSexEGVlqx/pts
afWXC2WXhr63E2sVr/DCKqivjs5xmTlLgODcDcPJvHY1D53Fp3BGFV6sT9w6
0qL5j/85YF7QEaHGawXt7zQx4xzICObt/PZmfLuF42OAaIODLoP1OAnpp5LS
W/UagT7NF+QBfbTqNO8gA3ml/7xg8H+L2cUb/vml2g1HzpmMfK+sd29NoHK2
yq9gknAmqaYivKzkUIcWwrh5STWrFUcOvSEqS2QD1LYAj+qToC3JwoI7VUYD
TZaKlvsR6NenCeh9GgsS2zwawQ2kwJCPabIQLi1/BUN7scOR5XqcMKYHbO5a
evnhhI2KKD7bw17dca9pDhtv8hyPsrFG3onWYNeULOUXq+b3Pu4zrU2GOZSr
aas+4y2OEQt4esxo2caHwOPX0fLBsb4XpI3lTdG9APsPnHcQTsCVeQHRZwka
rBTuHIFAk1Kpujn15JWpYn4YObuvB+WGt87An0yR/DP6Feao6dfk6SlyiZX4
KK1IHCLjBy33fx96zLxZhGk76X7oVuJcTXAPmg2FIDk7Tl0BmLfK1fOKq5ac
oScdaMbHSYRHOupNJ5v4xhii2kn15dQagGLQ6XJ1BjD0VTI1z+ZpChNVgiBa
HuAy0ceJbqGes0DnHAIVEPDWhDoGr8OjpdXWO730Bn7ReiA3fmDjB8FnNtgd
aW58RUQe4HRPRGcmN8XM4CA1TpTXl31F2QRjdRA//iJdlPCdVuqguYM0kczj
06yLo7DOSawMTLryV2oCCpucs4iw7Fbfg+a4MqEUJwe4DDBvPhxnS2SpZ+6C
e6upGHS8qEHWvrakaJ+94UgFsxCl0QCAUyoCR7OJmz+0W4JP5q1LiV4QCYe0
NL/Bc3Yx2UeD6BpYCeNI5p8B7ajlSLdt/QTmlpw6P5m882AJIV8/ma9Sjmk4
pHjLT6ZvgG4TPSOSKUmGy15Q/AMtye9/csFqtsSBpDRI7TZNCjVpHnpvY7Bk
d+4BX1tNPjGhBGCoEIY/GWqKnonHIpUrWyzlo+hShuf2t+xp2wXl5BzFnBEP
FNEKT462kCker8PnPvyP+i/ihbbETz6UStRaJV5ghnYLdFKL1nbUc0LvvoNW
WC271FUAGJpFuke50aXbBPE5KdIULrcgW8mJS9krBzeglwYdrP8x1rHUFHKU
Iy2tWLg2MVritn5aUH4eCg92E+91cnfFWVgw2vslw+M5uCXpJ//S7NXHSqAy
WqsoARx0lmFsHSfUoHeAUqJZPZaxhQM/5J0y+NcjipcAPaMx1GXDVGeFx7nm
8cCkmkNuF6ux5gz7CpqxQrFOJ3DJ5dXkQ5Zj1BcTkqf/q8CsBhQfEWcupDtz
wtXqqbSTN4GruddhuSZ02978ogLn9HjcMVFLyF5gHttU8upfWaW1FQ8bdt1b
5jZZVH0UOsHHM2R0GOA+PYg0fOXsQMBjx+Bl0Usqfth7M7RKz3OCywyAr2mN
R/hQrQpxztLhJnZ1enFIfB3r19FAapsWcaLiC9Wp7uS1dsPvKgTQl7rYPStb
WGoNRLEVCTSZ7LABg6XOyLe+ON7vhwTzAbVQagsSiQm8xhjRnBBqC1VQta5X
GMzu2EEgZr3OlL6nOtoT3WA//c/lzrVRgAPXj61kYi+cNSaVCxwRSS/+S0N4
luzDrTXURwm+8h8TPwAV4HI5RIbLs9aMHXYtEaGz5zXpQvHFN+zI2JTocMFy
QI9ULGiHpcn9UYmUGvSK7yuKqtXAI9fFqzB+P3ojAHiNWy7XQnyiHh7qeugb
4s4Z2/jtDY4icLXoK9dS0sDtjf9/gGTjMh/IRqUDHfTjxStWHUGdc2eJPG9L
o//pvWAUeZNCTAZdPsyoBVksZl6onYbw6t0e78jHveShz06Y8vshe7kbKPuE
REw4ifvWZnK2mxRebv0b8y27wQ35zOpR4ZdoNioicXxU9DeksltnpLaSYcVV
vq7Q58euHb2WQsbD8K+IXVdNclQgGatTlr1KDRexOUoi1uMPQJLx2AKG/20V
aXSJ1i+TYP/0TOQnHhxE3PAkfZSgsNvgIdup+k0gPNsBUyMrR4J9JR4bmV0/
umC/UhOMVNMwzT8+owJSDhkzxvYb4n8ntTOjZXcLAtzhaFZF6G7oID/NTe/u
cVvjybRk8zU1Xu26gbOjjgcd9V/j36t7O8ATHmFvg1MP+VfiRbvhJo8odhg+
mRsoP9MgeS0cVlxegclMLHA3jFFTQKMSKRJrH6wlg/smwKXG+iQ6woHInBPE
qT+0zTa2H4S7JOq5ef70jwu+ahUq1VM9AYPX6NIOErT8m2OHI+ylNBudu8yS
2z4/w/xe2Yyb3BTr0eyrA2TAnORo2RPdmtRge9yb03TeP7rNI+syvWXiosuT
s+jR8RmLYKMvohTOXGImVXd88+MsJtcoLeQVApo0SQAldPHhbpnfY/Izht7A
pSlPq1JzOTaXp+lq4oZ+bvpa+Jh1ETkGnr1fe8uy0V8jPQ09OujDGga2IbCw
3e4LjEvyTbfvCV+cJnsKFM4VeOaXeSocd5XgW+Fif+CUyZ/7211aVBaRoJ0r
eX1IMEAXPOHUeDKVYSQEKQ5HEOicXLShjC6xg6Rbtj7H/hyao4c0qBk8FCwc
SnnLGGBsPHshxYqPJNnxeRSAMPO3GPtJYswCxb/SrZvjLiLO77Ay28uBN1XV
dRSHynJREXgPI9L6JAOIf4EsVEAWVdbnjsHSFI3b9ZHzpaLgvC+1Q/JpteCg
XWgienh6ws3CjIMwXueeR2Tk4Okq0grpwGtlgIFdMW2oPcOedg1C+1o9atai
DCJefmWQf468CalKHhFMS4WuuB2/v77CLhibe5VaHpHn73yeurN+K+7uACLG
O6DGnpRsnQWcjmPiCsGJ9tWFza+rMVEyyd/qPdsB3RWA2v986wcEYmyfxZGa
KmpHD76XMBvW8xxJ8MILAcmbMpDvPEWIvNRUSFiQNnobJ3+/MP4XRSfbMXFf
6BtEzFRkptXZZ8s0wsi94ewacjTF2XPgYgwRIyuooyg9Dbh8jhzDETNCCtPV
W6lKsktZHlArjQCUJD9bBEjSOt1EKFZtJFbGWj8+aTS8mYDfwVVc6JpM7zVY
qDydieEfRU5w3GEr5v1hhT+1xRpKcgRhsyaPaNFBbprn5hrCahT43sudsYcq
9simdmNJP4e0OSZgsS4zZ6R+nwofoPv0XFWipFXPYN77dTbaL7QOffM7JPk/
HvWxJ8FC1dd6gQIkzvrAuoP4D2w2jaEwQq5DN9kMjg4cC7IvlEYVnKsN1xTw
ywXoXU9wcE1RQn9AnffJoxoRb8diQYA4JOZ28PXRMqc1krgpWd9LLkyUNRZp
832nur5Ne1Dkr4HUO2bPTSFPMf6t/JCJUU/v+zmmOG9BUFkE4Dxm4rbZyfMi
QiwIewI3RpVdrJIW/tHJlPNe4BbSR+p/vidnLkU5YVOO9mAm9Yy/cKjHLpmw
KjeIOhkkAUioysRGmq1fCfTqr4OzeyMUMVwR2ea3NqTqH1Pee3j+vprO58E7
OY6TAgsCfG5kL5nQwLHKaGhVQo1zcdXfqAhHl6rs2TeGjwWRHWuvg8OaSzRV
NBR/OR53xG9Vu1mFRaZ3jjGgcS7NI8A4OmTPrjFkDj8Hz9Y++jjoLhJRMqLD
3WuLXBJA6tc8EzOmV6+20d6vm76jvgp0kQTvAUCkBTOOEy/q9Tu8aVURnzPb
57lv/vHCqEYW7e9P+Qu9F12j1o9yM1FGSS6bjFFcXwChYrNsdDPvgTRaXLPZ
oCsaqm9pSDCpDpovz0OgdjetUqJHD2Bwd+te193lSR/RZRV5miSgEMXz5/jH
mDKBV0BFtZ05DyjSZulPu99f1OM9261NeAKUBwajpB4CjeBFCjeXVX4RN6jK
W00N+n65CIIslUomXF5tJ1T95BqKVjEN3dV5+K2QFpqUhm4MSpEdNyfrvtB1
QXklKRxoMEpDzvz3/K5ofUxZwRaNZjtulrSLKOM9HSGVPLKEErQ4tu8apHhZ
5hzoWQcHsd0CwO/yY9QK5V1/j8cP/+O3v0dZnacLQA16G+pNEKb4EWL5+R2t
W7zg9wJHdr3jQyoMDTLuctQ4nz+Qm4sY5bwTyvQSqvhLeVVEHe1EdRtZEl9O
xluqlfWC9Y+jVT/56x/EuT+6uHiuW5cv/QebriFPh8y/rSbOtoIKzRM1Gx8v
zXmZSQ0z49HQUB07RuRtvj/NdZtGwydjro4hxNVQGI6e7OZbTfVOkMhzz1ef
UQVff1CpAznTSlACH9NgSVVamBt9t9UDzNyRlMzeG3ibsKLkYF6Vu7w5X1LW
H7FiIne1ztGHLB/SRnHw/rixzF4I+PO6xkuI3eaQQWhN2DgX/1XE8Ui+Jeml
yxLFJtfSkAQ7cuxgQCtFZ2YW1XEo5KVm29jgu3kJVLBMebwZwhUILABNKYVB
rwM2x/wAtYGaJ2WtDj11dKuDf/9XhmvanVTQAyIy7iTQtBF1HUOvzNRabFDh
Uz+Z9OlHEHG+BhRe9oajnLzu3oq2CC+RyUXJpu19mb8oCTAsC9+vyuomMlQZ
kC/eJW6MCkrhP8YRnt3x8b7wbAiVnH0xIEKULoV6JExEnH52irqVQ60WauOy
mdxtCd00sTCpAr1zp3u0f0fU64IEfPyC+v3/5JYD8Ua5T0asyZ8BkiBXSFbz
5elM2G7FokwkslEcI+8k7clKktPDU8RWkn1YxZgQwLb4XAYNpP73WAG39ngq
+rgEPoTtgJfEpGAQ3tI2P+LX/aR91s7NgFvi+hl0RWCe6y+EKoAIWO5HNALc
Zl4NcHB3WmSuw2duxoZ0gX8kJScmilczmFVnsyy4RsDbhJoQd40Fn3Kbpf3f
caat8Pv6chWHTa9TZQ4KV401msCLba0MnUDZc65kfg3CsLNvDJ7tVfrQRql0
RwFqXwFEahnRWinljZonNpgotMXf7Ox79dKIZoorRqHpIDT8vmlZKRD78aFF
JslfGMIDhgx24ask1y5PvxmizN4ZKxHx3mAxomUtXejc6GhXJf7hEB+bU/TJ
bcd+/cTJkIDHFYhlCyOw0qYzuPm95if+cckHi9wtFuDjLhANYm0INWXkM53i
XsOe7gJGCIkOYsrwI8SQGqIzSiOnyLLysrwNntG7cwlXhQ2YCxgN9a53AXek
bqIPOvL+D3PB1Yi6YFDTZy91EcQNGLASsYezEoumHJASpDDC+DIn68YAmPat
dJKCzhqIJ8zn9g2Xi+ExBmvH81auPvjagL/Hv+zEyRZMHuVD9XND6OeJQ7A2
KnIikEwYAO4CL8qFymFyuAwtQuOvqG39ubmrxmdpQZfekqU2y4MH29PE9wwW
G0BZFRDNscnDSPEgF6i8PB8Zmigt5VkwLuil0wFzjGZ3F/OkMD+y1lyiuddL
qckTjlaH02qbFCh6tTOlDVb1IG1ur3LmwbDslYfviqYFed+pYFtckUDaJgWd
732NI4Z1svQcLgcn2xEU+6cI4UzNjIkixNxgqrJjOu3YEVwZBvfiW8La4pMr
jwLssAtzHtF6Fd/cLAtjF60+gtoVCOQ+wf2uHnHBELwWxSQHB7yqIt3Wx8bE
nUT1pEaLCNpODhN4WtT2orrSqAxF0XyRhH4OZlLgWwoaudZgZJN096F31Y1Z
LGkOHJj657UKw48OyFzEx2pklDtSP1KTOFc4sk5zXQfkRQLSnGfYMfoOMGbY
jsw49pzJ/e2mOW3TeMdwRZYihigrJT4cSo61hIYDFMSQbsLkg9y0StB13ijD
2s5/X9TsZDBVIAzXShU5RIkysESIt3RcbYSJpT0+o/elAMkhQLl3ezgLkOZa
1rVOBntENABozuhPRRS103bRrJlWkn0ALFF6a5t0pYuEfjccCYbbBMT6iOrp
FUbp8yiRBUTUDU3nlhDkxTUnVwJfnubwCL4mGkHY5XPIr3rfYw2Bk7RxcP3K
PKxHIWhYzTqpTRCIoPgF8e39UcFXfU1QrxXLjtyAS/GrVlusA1rNXAwwzOvG
LSU64x8qV0CCwtvUNabxFNTjQRBrHY3k5WYcYD3/SrR7+aP3evacFoD+I20C
2stpJlSLlzSJWwHIGvu15dvQ/nQQToLMVGYvZ/EaeoBn4U2xQKUrg6+k9S0i
zhSvDYsSoSaGgqjpl3bTdUIYcZzu49rNvdAeiVhKxPbSAEZNSU2KXwyX6Gws
gxo4qd8z4PU2TidpumvEaFbTyQmZozma1v6kZ5axu94N/r/Yqda0u5K7h3++
QBRVNEKwyTM4aBFlvpTnPtV1jri4/4UWmeufNbl4pA5Q0vN103NQU2K6TUGJ
t0Sq0lRxG7AyzCS8Lz+SBLUp1Pt+oSWhteZRQ57eFKnKFGKXA1PiptdfNve9
yNJQJ0LStgen+S30sIVWO4GPdRUSCkGjPAbjvVEdR6BCIWseif196wrtQsvj
R6TGCMyeFX4ifKzduZDYx8X8y8CP/VOxsVIxUUyekL+8en+83ANOr2sbGQOs
KWx+XzpDG2Fq+gGZMqvppVMqDW5AHK1+HISIwM1Jqe2muQIZhDSG3X8CDTUj
KnTx6YysJAbc5sHzBINLrgK7hF8Pt1ksxSEIud49/n60sWbdLJxGkd2+uRYA
8eFIF3C92GZIlZ4Xwc0qLWKm+EJ0ik11LUooNxO3TFA96NV1Re+XiS8nGjgW
FTC/oZ/WWTi9OoxbHC/uuk924wpzhCwYeI9bE5Y3FAgHfDZxaqpWfqNDFRun
LqbYkLlsE13YqetlfWqhTJ5hrwVOZdRT+0mXpbmXqxXGxeuG/R5jvKMnHPLn
vhoWX2kcIzTrsRP23jt65mnHZLCDOjtxTRiZOnDm398jq/dwvPyCCEzgLFzy
QqDVXrOV6HmOodMqwhRktZN9oZeJ8ShTIioZaEiYycFmEPEsPftDBTGTGIGl
68uIEy3BwCRn3ZJArUNwApSmQdprwh8J+kry1o1RiuK6Y3jEygNPzGxEoCPH
Q7j6O5UkbgV8pQnD0iyJMUWihNyiCuIZYAxrM2ys8sqY51luVPoBNxqILuHJ
jLuk3bXnL7x/UJzQTS4TlOMuxCgQtgz2I9tnxXL6UWZvV8LEluCg6leItCFf
GjV3ixlNzsrdUjhMKAsGnoIeGnh5i8p2fVFSuBA/TbCuIMO47SNPwFwyjkAl
2tYW7HBW3844uAxDHF9V1/FeAUZKO4s4un18w+XPMP9kQDBgtPMIYVYaQfTT
o6TAs6uytRg59XdSNG8xFEs+hyujbys5Mm0zD0pUhbTPXxyNzyOOXiRaea6y
IUfoKZlgEt9f9HvGl/6hp6rmsbFPFrZ44Jx7ve5vJt7KjxyWqkHk8QyAPlDG
HVZrR0R1by9ospHZeOClS9EC1oodh3tEIdOfrpIz6sB9cH6wEJhYVDie7l41
+xJ6xGMMnchBEtxusLe1MImBzAPjFIsehjh4l8Dv/m90wRvLoKC7Ie5U285E
BUyyafB3uVUXXqSDjIsiGjLtyV9IA2OAYNU0RxiAA4kqz41Q/zdsQNVyfn5B
loHskyqn0p3QSHedSnnSH4PCt9KHEHTohY8P3w+985/9pNZAjF11GbSthcz/
AvCnnpr92otkwrTtz8+FG6GVq5MsBFblNNFxnr1io3eY1BnE1c2+PXGLMvvQ
W1XAjS6/tKxk6z7tTqX3t/14YnfJ2Rcpp/T+d0qwjxaC8Y4uJSv+uflvIXu4
3oHPbdBdrlKGMr2rPKCrHnA0HEfFWlhzrJLu2VLTa+sBwS/b00SeFf7XtM93
ZgfMGOcDyqcK+uhYXPAfabQMST1wl+jAvGCxqpIMTiSYdFYctTPvqa+GIEsh
eLzru+znjfBv127s1tAGdE/k0zt98FJnTkUUO9NgxG3C1NAPbVzfoBHdnfg3
liIgcKdtl37+JhJ0BBnvaamD0/VHH1tTbFwGIBFt2ie4JOkoB+SMcMKGfC7I
yXwNsg9K7fXAdfkhnIBdIt8JuHXg+Y86zkOzwlJlFY7jZ3hYnIDT20Y/hr2y
WofTSWLXelTP2EvEOKaVjeEVbeDbtaicGR8HF8kn+edJdyEoBSw6uPPkpR22
Kky72l+FGebFn/SGG05cmaERYABJ3WSqEp79ufckxeYHmbVOLoEZjfHyqzf3
PwxDqTA203Vzz+CVfRjH78g2PNR22Ob9Cycu5oynT8/6a+4LoVtLoELGqdS8
Xji18hkvoTHXmTMdyOhGUauwnrvEscMVEZbMFcmkR/EO448SwYP941wrLjSh
PKiIRKf431AbnGWtjnXv/SQl/xef5sWenB6moPiwVbr3Jo8CjEvG9kc6MSzR
Nu2N7h3nrWll9GCqhfDeQGdeAeI3b6aXlow2X/nuPeoyESHcp0dn11k97T78
WoH9XQyBxjfKJmV0XvWaD3rUvgblRKP5htFxCRGN7i1TnUPSeNnR7UAnIEg6
Gk1ZPo6B4WW94tKqH1xipuwMY73GT6Yd46Co4HLhG2bpqxYKf0Yd3TE3bm54
JpVeDCM4Mix1YjBLwiazy93PMbqEG/iZk2VV7sS+73QRDo4LWEVCyIlLEwrj
7plKVrzjU4yzsag3AkUXW3IjNjBxPdjYzs3pig4OCPhYgMlnDn2Z28ReVTv8
2H4HT2VokCThzQwUU8dxBSA8AbnQyaZuIkisGzVqYP41GfgPSsJFIu1wFsc8
DAZJU9JhA6zcoj2s+TNfFX5/31dqOcrIL/TWEG+nehWYyRFUaWTyCx2RjC1O
3z73nyZ1Cv8Sj1Skd9PrI+gxFKEVuyjd8wIPu3ZJQZ0WkMO1/PaivfuWxJpl
D5xXyj53IGulK5tQm45G+QY4M0NzUTGAXx7G46xEmMZGXuJbafXdxMoUjFy0
2qvpzvG8i8V//xUhNfIKu9I+a36MnMFVND8Ua10KhnCKSSp2RW28omlGocyH
DQQYJEpptLAl5b+ND1Rw5k8vBd+vrW1GvOu2Ua0satJJ1gvO/0TEzP6nuNv8
lkOUFCVw4zk9OaETbLaeQNwDzb7F7ZLX1Up5yhYtqn0t21kT/sN/pT1hLCqJ
oOy4IRHTtzfbvrrzjgayjaf5X8E0HrXaU8HbvHb0FKhC7FbKl1YCbttMv3t+
GYLWTu3a2o/KcuXWZvOTBeKwk5p76Gu9ry9oqCMy+ukvO0PXagBMQIhD+VCc
uWCCs7142zz2fQ18hKiUlGrJsq8GOQhiuTnrOu1TYM7g3bElw7heXSeUS9RV
nM2ZxAhDBpnvMPclPulnHWVzOeaWoSG9gEWL76QvMv32bi/t0KPOZN1Gjo21
ivkYfiVVwc5EWuEK/LtMAbIMHHm7/Spqg4wOY2ToxjAfmUUjfu33ESU59Nas
Ix1gVID1KyUDrV3GhHy1m2m5FdlXTbwCYJrq/o6YLnTGZPKL9zZ0k699xXeA
xcJhYJS9h7hIvIpdKkz4RA4o47vEy6t1gw8rQZBgSuV3N1y7NZRVgjSFXnoU
Fc71MmjgBFYZ+KJfHXGtwwmIZrhZ+e5xKIsC0S+Mi381YavbCceTfXR/QdqB
RnxRVp/rvhayJP9kDuX2RpnL2N+8V6/H3yuZeLsAa+UXOv0DxOnKVe9XFsbA
SOVP65/jX8pQOag35WtB3l00V87JyzIXcRR7LVsg8axdthAHUCxTV1ClIGCW
ZkhlXcNUSb5e5sIVixCNFYy7ti1N/YtIYoelzlKZmHB8iR2t7fzE0X4VoAFG
lI5OEvrLi6HmyJtKBh9OIya8WwfgFDFIJkPXDzI23WJGsP/j9vreEMcK5h6I
uvecI1I9hVQelGCrj3LHlBJhF5RAIIe3eYxKQP4HoHkEEBiCTMgMQa0BGKgt
+KRCntr2aBC7zd356xNlOQJNv4b1Zfv7X3QQfCeivG8ZacJYNBaifaQ9UjEb
9iclzrN7GYvIUkwww8E7P0hroWdC4cLeRhUtyzSDKHBiP2zWAAax3Up7lORq
DdaY1WYeTCdPFPSFdYWso/iiS4syYMav0LuhJ+dIZfTblJ6YuOaFA6p/ZbCJ
VCjEFOHE/13J/eaMnw+ae759NX41l4kZVdlnsFjVpcx/JSQ2jI9JNMRurci0
CaIfCGXg9L9kugI5rL4d68ToYLNGrKqxBkAKqe6eUSz/EwWSE8iRyzj3rYdc
QZxtn0+hEmJRkexd7N7+wriR8ImNRXOLVhIWlybbBKvMclpMAzfLB+O2ZD/H
rE22erhNptYTHcSzKUbSUt+U2taY+G9AxLtt3qQNEZN+p8dD3UySdJkK7v/g
sDwjGcb/oYuUzUVMzvJxWVMB653obLz62U7jNmTW1SuRoxo5Y8DWA6kBMGKg
hTYlVRP7jHJvEVY6jk0EIzqBJlmXjqj99Fsu5TZku8mG+zZBpEBmb+mwxcsQ
ssKNlp4I1W4i1+Tr6K/jQIdQGiDss5uI7YDqUQ9OsvLqe7qSWxMmPhwFBLL6
xtJrS4iJZxmkUey8OhTfgNfgZKIh0p4eGOzmSwuaDtbqVLRQyQSIX6Oxc0kW
zS9fBNhJiR2PPQaS5RvYWjYK7pSTwNNr7qNgIB0wrMBxlqSOtSWu5xh6sYSV
pBHgZCs7eRtbuhyrTHtKcP9f3t2QeXVKEftvaDs1GRlSH/Z0OnSy9+S9gKqt
JWu7H+dlu9VzPSxs28R5jGdRxfUE01k9nAphNTFHYNtETmFypLn0tVmWpHsA
8RuypWw5BhdWIxbL5kbcmSoQosB1426YGMMjXwvq9OLSosn4GLbKiIb11du+
zH/8tJfBNBjF9SaunEEfPXCYMgvl0JM494VxtPvd0KggtQ+3eqlnjdoco+Zn
lZCBiCROkevDagPAFdUmQi5/O64ExEaeo6HxUNFMbc30OtfZ7AOEfheADjJT
KVHxSrH9lPoAukNESbDBtiiDel1bK8O0rWpQ1XJe17wCtsChWhN2lGtPISnL
sLbrdgPoqPE0FymAd/okOHB14i2UfdLHQCf5YvwxK1jnriBgj+VykB8WM4Ed
Hc0QTHnXMvWVx1QTCYTVxB0rBL94LYUSCVY5pwPxjD/J/DWF6gFeEzQ8eoBn
RkACYUMjA2MDaNKEoMs1znDt4FWhTwfQb9KVE0I+GBt65vdgx0jAxO5Ncp5c
YpDfko6U6hJzViHeRpBkVa+B7bZmwpLnxdE7hPzFcmwnfH+utSTWzO6omRp8
jsA37BjacItW0dHsjhIL72uEBl/Ibk4VXKTans3pGnj6vD5o3xnyUJQFzOi0
xHvMM7hs4q6cT1e7QnWi+lCqTMXzvfxf+AYJYCP3/0TcCSMbj1yccRp6kdxf
XAh1gG6MukbfItO3PFH05AQlpy8cWmyv5vGwia3MtmJF5Ypx/Jr5wUYyjhOT
LtpggH+QXGZmuJyKr2eu/5yOayvaUWVWWYuexslROp+VTc57uPMoXA9p5J8A
ywCQweep8uOdEPrbdyCoJHrEEW2k1MRUICgWc8OXhaeCa+4RbBsuJRADt4r3
mhAJD0BOp0yKPp+qoZOC1GtVQpK5AXVCPgx92/ry+FGg6B7omZxGIj5RZ+Ls
e2qmHmjOmo8DBdEW8v2/vRZLbkFSUg0FgViBy97gMhNnF2SCzXyL8RxIW03k
g5JEAyM2TSOmbrv0DPjAR/of884BfD6uZ0Q2XjXLYSIrMTNKuFYcM4WSNcgB
yQpYtV1COFLg+xmfyWUdfRbp/iZ0jDXFAqVlrei0BtVSn3Vx/j0ytme+Y+tN
eoaWc3HOB6ud9BVornvJTScdao8/Ki2SL02DP25oSDu3GzKsC69Ng+fAQN9K
X7oL4+ejmieMK0tdsEyFfR90Bxe7oQicVQa9WbmS6Ogi2zEGUuzXIoXvE0aq
N0qXO/5DVdDqg+PqLww9XG5njIPiCGiXQSiZa9BRqciQPAIYU0+A58ScK/q6
6ISDc0gT45JXtauPngMK895u4yNoXDCkcRapm5Ize4O0acS6rsRw0RhOByJJ
dSRTvJiH5YTHGuAnL1OhMg68NQLdjTAZ22BRcK2fTfcJzzzoPGjv2K7Luvn2
RHJM6QSHf0I6DKMI0qbuqcuwrKGsMtNVROKiLX790WJs5bXDEna4wnQ0I3TL
61o5k4btdaAgEkwYIQ50DynUuK1fskn6+W9VlDfPIOG2cFl/qJgkPGSk3uaR
gpq8TnT6v4dc/LizXje8OeHvOK3mXYamaCREOEJ/MY3FxMrecfVXgFqKSxFg
jwCvHSGaaZwxmHn6+5rEjS9Z3dnuEfrTA5CXZoCM1ZCO2l+bPgA0ymEi6Lsd
n6CXHwFZyULUYmZ/agnW0uI2wH3lLM0sshlKOu5lZfIrG89wgkIJ+OzOym1j
ExHoW00XD3AoMuuUW+fAqp0v/NpzQm2BsoTI3YGpbsKg5quUiCtk69Q+icap
6lvsNbCsgDJJSo4otSl4xvqG5Q+b6qtxDaj2vtbzj0Uea0tVazR/MSmpWZrY
sKmo3xEuveUzprTvA6ind6PAzykjenxnloPxuC+LnJo0mJb5lQ2n1V/nO4l8
ix2Fj06a/H0lmAemUFmNyCInVblf6Iy6oYv4kLD7LHDQXoRhle1YCCDqqtM+
56eZBMCDihXNTojYjZZ1edcGzMSbb0gSNcTwb3j5WQzpxfjlsFMDtuZLgTJx
uxjFMRR4N+00itMdml7YRoMjG7Pa+/Cu7omEBvsOnFqCUUhoT0XR0jrSdyiV
FB9/CS8z2ZsTp1hs3gDrtPiUK09DlT7erH33OfjKEYfKc0kLHlEFJzUVJ12F
tcPFfUAxBakPVPFGCCE99v+LroN1W8zWCWHM7I97O9bxlSYyFf9oAGgKr3rf
RR4/GSDd4t0DFXlNwmCY76RICGsQ5FI/6qJTiqHLsBzLC+M8NWYmsTmCY2HM
IZhMYwPiYihm2DMo8EcxPu9zPnTB+8o1ZGPE09PSIK/iu4u6wPhheZeHW7NH
hs9K6R4R6XKXnJdnGwIRMHKGQMS5AGeiHsWSfbzfz8tkieZZKvvd4j0s1//E
rgDy8yx4XRIrt8pFSyf172mzTKjk/7VVvH3WVUSJgXQr6zxJ3mhmcpOoQH92
8OUEb0SVoGhsTOXMDxEl5ZbzlpVWQh2syZhOgNulnCURSWcHPOZSW2e+qU0f
RdBDD3Z0BsOYDMDKXQkALVQ0MIvkClupP9X+//f0lNGjdUL5GLBC1gQ80gTj
So4Gaw2EbdoQiHGUqMrxyR0+vFAdqGpq/za1a0SW7kyNEOdh4W+HE1CjYgk5
v9Aye0QXArKHLEofHsKqIkx1H0Iq8fcvrEPMpfeJvIfkkGYucmORM/dFgrDw
n2/ttLYg62oDHFefbijdsfmzzQHvFBxzlBPB4EnPRq9z4XXg6peBjrwT7oWU
dCjB/iz4v3nHYx3NDqc7Uoi1iP0HnA1q4X03bkYlrwlvjZx+5ZjXLC3aayIa
/hbskSrJgf7KtdfPr/YPWPuE0aCeGFtwHhmzBp/S6M3cyyXeEdB7qFYZGqp7
kviL6pt5iWBAbTkKKMidzpM/G2MQB8eyYhzJSv7y1riwt+qgeEaG0TntvQ1e
UGjPT1raq8PBZqdv1HctGU++/FocfZV2/A/WcVeXrm8otr05TpxE+UmDn2Am
C8kjNoBAZPqjYsYf8FO+ANWtpKWVLY8UJTpCwds71egME0iMEzaKULHXW2xW
UhA9aSo9wYujsVh2nY6f97Eiwe4nF3BGT9svn7bXYLlAoRUsn+B8iX8smk3w
xDYqqie5sR9EtMN7KZ+t9naPf5lRgJBcQEuXS4jKjsZ5lUlHCsoIaV4Rpkqn
QR7m8RJhTsbweifalqGIuCc99aqayxi//fdgQPJrpIdtgUNDFfjdxYp0Lxzi
xxc7GnXl8bJHooiZKicM9KspqS6JxhOly117alfKHxAtPYKY+Lz3XO44Dr3m
/8M+P2/WyRn+WEYYbQ1uChEQ4y40gSRp6vocXxOz4+0Dij+Zokso4ieFoEth
jFiYl1onVPG/E6hsPnnrCU7on/w5VyIPMhB2aOlS24XRVvgorGS72hyZUOxf
J49Kklr2WKUcw0zlz657GK0TSIp1LyWcsnQtNozYAE0/ZmuE8K2qu5DksCIU
6emeHirf/QdpU74mooBXneXqY1LPTH7Fjs2xHUs6KhzgznqVPyoRgSSQJ63R
0ODrts5PlFfikMI07AlBHMIRD/Uibxfnl2fPxgtc6VYXahdLQuOVGp/n8tSy
wp/lHrfyecTpYA7mjeSv/1y9VziEVVrr90GceMSuQuHAo8TK4IVM1EeXp7ru
06S1PRsO/IUL7MVDdhV1qaKcmEEoOLD/kPHdRoo/R00G8DbCPgKX3Z5b5qWu
Uu5bsE2ARw53wSVfoe3zJqyCR4iHcDnCJ2plj/604IBZ6Bsqn3LQadotfNwP
H04ocPamrMJCuA0N1gCAzb+Z+LebvrhAUvwWRHKBg7iHHenxZWX91RVySTPQ
Zmy8jD8YcTfRFZ6VCV/Xl4N1S+gMKq5//kI/fDz6OL35CTT5DwgsC2/o4O8A
zwR6vttQhAxHWl6I+zLh2cxiZnw77Kg3BMHfbYVzy93BtFtSOkvPPevx03kH
VAr+XWIM7y3dfulfzAnXzSa2/rpeuc19SHIwkUkULwfO3nthSsJJRAMz1jU2
TfVou5gRze9OzqsbLiVHf4WJj/E2ebL/HAoV3UCDyi8623WH1nvg/+CK/S/5
I9lqyiNM6MmfirOPlkUxD3P3Sd/O/USVMENfxrfd3xiQyMS6MMcUMfMZZtR7
hTHQcJD6asuHvSCqaat3EsiF/tk9gj7+WRK/Xump3Bk0kNzWHJQLDJqrTnxT
3rXxNm3e8l/Xm/j44Y7jTOXrfESdBxtMXIm+9ehniCvLQfvxjwah+mdYt0aM
0aBpZkvcDLhIjJBvjx+L2jOqbLMBFlZmSdnxkZUYfIUpsXMMTjYLdxV3smiK
RWItK/NJHzNcAwNwPpkwi94DQcSxjLHkquhKwCEsh9rWigH7pj5B65YcxH8S
wkOVHOM3/LvAftCadOaDMsNvS+iKy+k/5vEglvgxgqP9+59PmO1Cw69R9dqA
ps5b3uzbB6kqC9rW6XxOJr6a6LXzPikmF24gzpIRLQJlC04EJTJoJ/eT7lrv
s8fDBxADM6eNFYqsCi6rI9XZr33miVj0UcO8n01viUE6AIT7Hr8I48NO90eD
ms3oKxvLGXKyZvWntEJD4w4eXXyF8SSj34NJqbVpE/31Z/MkhQv8f7N2P2u/
JXzDVOMzE5bT0gjMdohbJvoMB7PPHAsDWtXha1Zrej/zjp9pv26xHFqqA6Bo
9rkbVUTSCYioiZN3IgQd3UgElrVT+r6eNt2p5zKxI5becWq2jPPOZUoE8VB8
s82eZpP8OCKD0C0pdZKN48h4X7d4pvcmIVWOjLKbf5f3/YSCNmwT59xcOO05
oVU6/tQoBE+cCD1gwPQ/IQhThwRo3VkA3NxnGXPJYPdz9MD4j2K/mufsH/XA
RsB5MEaHroArN7abIpaXfUE/V9qSGVcqc4VfiACzWEXDuq6oTdcslixaydW+
pJsCSIFGMCLKjUba6wraH3jGjeROjJmYcAQoim7jHEKREsJJDqE8FsUjM0Ob
PtlwQPWocvh3bpp/Nt5ysITZAKOtQA1Xp+luxLZCm7v0NQD/kBmJ8m92GHsu
sOdAKsSutFKI7GY2duamhKdeAqPbzE/OJtYHE11Xnx+k0FtQEmFf8ixFErAq
4t1XENVq5IjqYzLW8p0+0FInSZ0XZgY9OCYY9p+JLW1Bp6N2UqSRbN7WTJCq
kYAift1nZkepnAzBxGPdBUN2bpTB23p6146SuRQ4WDOfhX6tjnPubYFq3O/Q
Z9irQPyIoOlvjqxPtud7mUaN+mlu5e5DqZiVGekqGQ/zN5B+wgGaLdwpd4s/
80IMeKOSZ5GHb80T7SlS+oT2gbMadaTQ3rx5JyJrFxzYlPD9i7abAIkflDF0
+b32qCFnUGyEY9XiUAHMsgL24OK4z3Kdry5cINR776o3jHyMDOFYpdsutmzS
VMUCySYNDa8dW+t0+ihQHC/Qzq1Ub1purrdevwYaBxJTVq/DhI/JW53j4s4j
VS8dQ3/WqATMyAAVocMvy94RoMcfhWyCa4rtHiSa1FNthIoB3axQnsv1I2nv
ZkneF4F6bBw+vq8Sfz/dKsNREieiigNcf71P2C7FWUXp4W46uIVbazAdUZYe
0Tn/tQuPBfU0mNjgxDodpR+K+2Ir8cOYEiQzf+nRsvuq0p7ur89Bz78cHyjU
u1amv/neywgm1Kx7nXIyvu1hCI2PyEM6xZ50QfVOZABBXtOo2XZnC9o2UWU+
FAVFzOrEmlzj9/70lWtZrP9/1TBqODhZJmo/np9AJuggkIs7HD+s1nK/WEgG
pbjLuD5v8/ZFGWsno4EFkAKkk4/qT+u01Gl2dTmGljSB4LAWVe/ZRWv/s7MI
QpsTV+e3Prb0lQ5u/teXH769KmILEvHwc31pA/w/JLPARnYfg20NndD37iLu
WazjlKqMGj8pnhzK2xqIG8jftoCTcVG2OptzEhTYbRVwy+0A2hH8e0S5HdSX
DLwAMGDNJu4lTMnJ0Xnomsy2X1IMsO3e/AU43DLgEQX/nfjmAWwRND/yApBf
tBR1sXO8aPCemBacApEzwfqm39NegJbmPUfJXtLWkxft8F8NcHte25NTGTUR
ufG2rPy1WYvESUe0E6gfWrZHdQfOHp58wDFx5SOpNUp/9/tQqiFlGCuYObDM
foVCf1RVUWs12p84iF1+NvXLVRMA+TwUYVlytWaWbYR6XlEmCvHGulYFwotv
eQEU4TIwO7MByagKjYElqSq/1fpgckiTVz9r4hBXNJ6+DxElInyklr5z1ypF
A6LoaIt2Uh/wrLppAeqT7/O7sEkY2Kuk5BQ9fWAV74X+l4x6zaquSgrG2YSm
Flm2JeWqeBRKieXWidQKrxhaFSpdenJ9FEF01d4LsNtP9Ib3SrWrbDFZAH1P
U3n47l7KqpPeSbslfyb4EXunpyh4yZDvb8B4hnkmnG7gqFqaMKvZ8bTcV3l3
s+V+5oSiCUwcsh3k7oH3HGuqFQkRVfM3bW+J8QtsuBLeu5DmAFtuOpRpYeQl
xNbsV3Ia8J5KMPIU7kR0MdLbsOW9tB9jBOBYmQDHpX+Ark0xYtZ+yTED0881
6X7IXYgnfbtVaC7wz3+am+afJSi0RoU0EBLVk431FaCRCmY3LFBPoBAaeqoP
7galQ7chjqDRo4lJma35vwZmsG5tsCubKiU83YYI0pZ4IE99+z3UAqXp+hZy
75WaTa7qDabFok2l9AvqSY04M02KK0sVhVV3oT1ZlTsJ4dKeZaM4JjZMV/yY
NELrWe6EIZiNuhsWbdYX5cjVPoq48+cGi1thMcwKPtJgdqlPzGb5xdonLMRW
0kpwcXmJp4dTJYALo8RUd1mZ807OY/WMUT/3GFYXdC+jfoEZcgO/PqjiMYhu
LEqqykU5hGey834OFPgm+PlwLJlsHLA7bUNKgy4QCZxBT1FYYlPV6aouAc2T
0UiEXnzKzRh+193+mvkzuApUg0gyIIJzwjof1+m79hJV97kh2Q+MGctv+JoQ
rzTt2G13zxfIrJ2zHIMxJATkJaaEQewpPAqtBQ2VnmN8ggjtyhz0MV7TzEDw
8eKcgtrlLd6B7sEFkt/mDLtL8eCvRpgTzpnUpi/0YPvMissWXug1J5GQXMKd
SqmztyNEqSr2PzxlLSxSQcEsd+FtpPPo7JRYKynkgDR2FZrAk+IaTpuBpqk/
9/bFxHuKb4HaxshKLQXzRA0sCgo4d/zCDGJl4s3AJ1MK7lIRuajJhBpPi24t
VFqgMkOlh9uh/ZjxmEzqiHCd8mdWq5UlK49f1uPDkrP1ECAfsQqZ0K6B4/1n
edrTp+d4LhV1f815ZekDaMz03AHf7jDi0nh/0UXqMoNBt/Ldo4Qui0e8kY/J
WVDubNtTa0i3PbLonCXYpQFJqSkRZvihuwyf0EsSLaRUi8B5p8SMZGF6dGSi
0LwnMtnddHhWQ/J/Cn9ebWKAYiK9U1xXkEfEFkCgDhQnL7p0liYmy3/cKFBV
Up0r6PcY48kLX+LazQiqnf/1d/7NZ8pQCs8g4apgp6rK896mGMCH0AdQPGAB
d9lTQM4cvzGGiRR0jEBq3+FI6/jMRIbn6BOdMzqQemkgJSypHiVKd2NRsAIR
P/iHIydZSpeTbdfKi0yYmiDZiYs76ORFSf0ueQOUNdh5I5RJX1//Ao7By1yZ
ntkF2pvzwJf8uIuY8B8ajiFtlk4dI+c2jKduNdgHPJgkSwHWZurrThaTQTVF
TMV8qxI2YoZSLgP7GOHzqKuOm9k+Gg8GbmQNz/Xs6pxEqk8T4UOVmFPaYkmb
WK6vCjecE3kI5MNnRFc3CXrshbpQm3ibC87SsPFZE2fYubLgik0bnbZ45T2a
n322dYnrFWdhgGwQRX6x1Ytg9mNjcf0K4C4RMAGaoGH7C88TXdecuX2Tk15f
1vvB0p2t4/FJnjP89c+EFcla7qG0TSqOIusqWLRLbV0+F3xbI+jOPLWqlbmE
sLEFihmUgrqXvR15iKgD4oIPxulMFC8yZKzoIijoZCPwq8beW0Re6DQFKo09
Pzzn5XzkWuGwArqKhz0itZ5KLIz/EC6nvmwUE3ExMN+vTY6GMoXyY/aJVtul
0Kho7IoZpoOoE28YWifNDqwdwqAHKpKnjVRusM0TS9Cw56qUpkmq1lTpSPcE
xlDFBEEZSqByXX7WbvB54mTHEuqhdlZddI9Rh6/2VQcWAuBKvHhfT69CpgTo
NKjEZFn/P6kR5lpmxtAU51w6ICUKezh2PANWzOrE1GHwh/MjB77KjORhpbZC
aAZonkcifiqoKo896rPcqM1yfVaCfWVJDGwqiNUeAczfTtqJZJuAOiNg1yqZ
2bkyyu25HbH03oEVHZUQdpjIEjPBzN3FLBKYW2bm1H6vDmI5rjO5akZ5eT72
zss7XpwzPEom80iEQGm4biTZpF4Oz3BlAIV0la9Eq2X258032zXVOTFr1YW/
uYD6SgvGgTalX0SCjRqUuNSR1XbM6cNyJ8iqotC6J8y2HYFkqap2pvgGjaEI
+VrS+IHdncIqkhSxhg/7bTl9uOLNnaXvhEgjXtJ7L1c5dObEgGcF/DRkfjQz
L/PBKdfLcoAqrK4rBtkazNv8IQWk7O9wUMbup5bEW6OLopVebWzlh156h4HT
xAI8p9IuUXwjsFnFHEjgZUjsADlSfPMkd/E8AQDGTVVkqcff5kWEDjQbLuZA
kTJFVBApfhO5dqThywSuGkzJubfOvLvATpxEb3xtlZuFdvydOPJIdpT5QlDN
OR0LdQOah3hJLibaEPzTXQVxkZzZS7K67PFSQIzGJR0wfvw+jJiQPlt891zF
hZNg8SsEd6zjPyE1DZpQJzL7jQYP94WevOGJLo/v9q5gvR1I9yyXPhH94FTK
yC+Ge5jYNiXTECEyNwbDVyXrRUEh8HYrCK/b9AEzpZ7Bnz/SGF0K9Xp+RxFY
eD4sxxTvs42hXKVv2gcZSyrxcgO9wYe6U6ITMNRm/XU+eD3OCZmuDJ/fB6Rk
qZ7WdKIYGPbTGduVT3FgrS6gDNchX4sHYp8CnWfYVbNq4NfmoB+juljHQKTH
wK2fg3PeTAQQaFQcjcZiSmf8tS4poRLwCnEYxwILa+k1U/I8sRJPJG8pqLOu
GxbWVCosNS94M0GJ7JwD8yrZ2b3AgriUZFdoCOcPSOeCgYybg2apPZaoEgXc
Vp+jQhHCg65QjhT9peoxe/YS33AqjPjerXm9km2Z8rHW/9xvvibK6RrbgJ//
47IHp/yBAt/2IPpxc68LQqPRFFkCyJ+KqM4ni0sTTeifPtppllaUq92cjyjx
8aOWvapvlZsglGy/DVzVSyVkRvepBp3sVZ0iiGFC1qi2ED138K6amD1cSOPe
tA5aKhQPVWoK0j/KRbbo4EWJYtZ9Jt+Ub12Tne6DvHzo0OEkxCA5qBUeod9r
3dtqUdGPgC7yJPGVcP7eW+iILNd8FYHp100Mnk1TVGg4I6mD4EZIW3+eyLUJ
WPpuZsJkdmbDpT9o1gcfwiH96b2s6f78hsw1jzk0r2ZxMSkZ9r4u5yPv5XXN
GSX49ppfbZuJtOzLuBWwblR3NliY4IdcXgm0lV9iy/cCIXWwSE0HLKoxnI69
/ZT8sfdiwZeOd8fzKSGqf1kgo5g7fSdfCD+1apQr5A3VN0qmxgQBv/Oohc+r
anFDBvK94e6KvQci+tN7MhLHaH3yFN43hmFwgBX6Io/v1KBLo78D0DGs0b4n
ICCzi5pcqNwLFpmoMEuE89upFZW4vBNNSKc2v0nDTb8I48SnlG9TXnA2QiPq
lWQAlplP3o2JbigpghU9z7VvBuzAQBJjqj5cqfxf3ilteflZX/iG24mUj2sg
ZP3BgCnJLgIYmq+9JsgwEWsR65EGRkc6qBHVYOvHzfB3SDgcd/OGnbub3vi/
9O8wjB9VLizG039D4YOZTzrqweMN76bB4w/j4sGAFDixuezJ4p4LnVJq8LMe
jPsLAbuU+LYUufYYePPCuvrqQ2x9eVj/SIXeepowmnLv6zppO+rQb56MNfgb
2XrROGfkjUp2u2C4XX+sCOQYviCAHWgsgxz+ROOUxN74zqrF2ay1ZTGqVxsc
s0qk8V1TZLbQwPt4nF5NVQhaAcLwOqS7qRI5P10ipG+2chgkQi6U2CJqIz2c
g0kyKVTZ/Q51Uvidt4QGgDYs5ozzG5lnl79vcQ3vFDSEU6+Squ3e2IuvdZSK
+6wN/psQyz5YY79TfyOXcHDVr2MAm0EJ7ilwXzOA+jGxsPmf9yjruJDiGSZG
lw4hzcQefnRi+BAX5GE5QRCSrsM9iscyzqY1XDrjIKKkoXpdBeSQhB+Yen2Q
8JWAwLHjcvTYl0TQQ0MHkdINLm8/p5xV7OxX6IPi5EQumtTsUMruFrB07BOD
+q6iaEm+CW1L9GL4VEsC3Ai9dpq/Z1jLQKWwcNLfEAkuwSmv2+ah1z+eWH3h
X5rdTVKFMcabo/avaXvKX/4br8pU6U1DCwv5j4CMzHIvcPNLxrYGHJqBoL7e
DirEwyIJoin/AQr8Jb0sVNKHQFVak2KymBhroGd1vTxxkK5gfm7NEzr6SJuk
fWZtGKtNmNbhp2wfLgBysHPKQW52S/tGTqVoR9+MSNFbMYw098n+AcxAuOdO
iklxOoe/xywpuZk3SRgcMa2OkuY30DizzAFrO6XEjVsnp+aRYhWyn/j43/qS
dukJFt9Jv3ZzAwexFtOsUd5vXXSJQt96X/H8nQeB3zMSgkMm+GWtsrZ7cEOW
buPqdX1KNL3hx39g1tezORlsPTz1ccyG2Ir6mZqOSVRlWT3cj0uST7kfk7la
hEEqlkyo3r22d3K4iFGJWksgrYIPg2dq6gj9qGrBkXA2hHq7y6YvsYpU4H0P
kGlBkbg1nUBhutw5vAlB+omFs0iTJtxor3BDs1kkUMkriBqrTCMF0fXBn12G
4AAL9Hf5hnMf1SLL8q3POySb6Ig/8ZtyORoDIiX1H82vapb+16BSpHpxolc4
WR6/gLjAau1lJraVmclgr3FEgB1x5h95Mfd329yd4q73qEIifha/6ZOzPpqq
v9fBOEpgSAzFAJXqN1S0P40ySD87D3PAdineGldDvqUfELsrNSm0EMN7tGUX
KfZ0qB1M1LUX2U1JaW7tu4sRETLBcqCF82SrLqgiRzEOezFVqew8zfh7ID03
6q3n5IQ3RQzajinLRgQVqNQrYjVO/gmT1MqTtpJ0j99osla6CHrXMpR7+dt9
iRYNi3esTP5Gp7k1/NvugPkbw0IMvF96K1H5Z7rLyAiHA9U9gPU91RjpRYJR
DarvuIaigO5BkuHCENWQQFqoBlBwfBDxSQlzkLX2EECcfrJckA3zwP+eyOpq
MNXE/FifHK8VQZ0XeRsh30J7HxEEet5IbsX8smvyHljVS0xo2LCk14N7YxVE
9gS9yDOoizsfMAL3effuhLQr8repYtUwVkSj0oBx5dt1evvOSaOv7pFZI73k
bpCgd2+65TpiVHOTXAvXH+nuZW9ZZROvvSoEIncYs86HAYiodVi/qNm+ms5R
a43nJPtIBp9OaEAXb9yAEaD9GJRx0h0PDWm4/NZxW8rVsSfI9I9w9b8YdPR1
OfgBaCT6PHdBxGPD1L3DM9hjdxD8Q5nnO3UexMbb9giEepivk7TKb3ss+Rhs
w2v7jFoeuIn6vInRGVdczI+YxY5H8CxToMFqLzUxP/WFDAqP1XmakAn7SLOV
qXBxYA+WUQzQpiXfF0OrmgYP/EzD6d+3DkARusnvuJ2mTnHiAzceg/JxYRgC
Z3spjbi9rh8cjZFa0iTBDE8YPEF8UVKTGuwS5I0ljLnrqmfMP4AFlGh4BI9o
Ta3+7+i59mqXJ+DvOmLV4hQHAXZF3zCvdkUWcoCLT3X0EAt9jp5hXz3CwjaD
H0zL7Xi6D+TKz2aemE92kEKkpITIwXtA4fNkk1CrqQwu2uDVBU8tABdhFte+
5VVA4fHSDOe2nEMPZPgFGPr7MbTA8l8A/2m43wCFboxAj9TfnoySZVcq10+k
I7oG48pbrNrK6Bfmf8Fuu2ii6di55pxyU7IUA8hjzqUnqqsZVfZQrN5+Rso1
5kXjpVWS2bs7+F8PFNGpUtWX3y8+0vGKMHSvWLfv4p1RIctmiWcQ+oj8aBBi
nDvQNBFWimuzVrxbOryBaDrGqMMDIZIByMgb4GpL2UAckc9dbltp0UWRVnaH
Wzv4j5/Ve94ScDK6s/SoJyoobT6Gx1A9gjYY//Ye9+Ik3ySiVTB2NVVISqH0
mYOeahkB0pTMTDb9ZkGqC2AWPyGIlqyoH+T3pSI8DhWw17HG2+ovWbChJp+I
I8N5u9AUhqBNoHWvpvgFuw89fVeZWtR7A6NyCnesnEsVLUudiojInWDkNLYd
wAy7bpWWJEQIS3Qayf7Zp30kIzOY2HFDwuNsM5X5AovxFe4nx88wOoPX1QVT
Rig9CBfyH3KXroNqGJUH58ovI5O/tKbs0W/nVQpRaWc1FDmyv9hpaevV7d7d
kLgWkIq/wcp83No64td2PN4uCjVf8s90kb6eB/yZ4dq2z7TUBjXi6pcBaWWU
RzBF0QrVGhaWxWVHWSxQ5FAiLdbkmir8YOPHopU55Ql4sVTrnr0PWt5racpn
DjuVjzjLb6hcwkcFVhCBkzfl2qDBtTF7TqoKQDjvj/0ow/NfZJaxL/Itaevl
3T52T8H3wiV74N/riY9dgr7i0u8CbcgKaJ9rgOeia3IB9pIwQRXoKcKJyqA6
qnNPoTOzTfKGH28q3dk88IRF/93eqklipLwD6LYseg9K0BIh+b9uYldbCQGm
nt9jf9yOyLO31ziK/9+hylPcxMV/xs26qnAVpYnDBYhLRN0zjZU85Y838LaA
/1CamGvr+267y/50qh+EyThnSZg9y7NkfwZQPYhepLR05CwdnYlywdrdonMJ
4joPWNRyFGfSUS+TAvbYlM9+e/YhA9iLl5sJhlcGUB6lcIt/xvrarSdZqQQg
/qV00yANKmjWWUTK0DGwyOnoRMIfDvGGle/1xuf4HdUfFqD1R9YBr3TZ9EHH
GnuZQO6NXVIsr6onIuYrM2YSoyHzn4RGkcesq1hixbyAzv6cj7n9JN4z1z2F
twopOWGNlPYCgHBdkhw2A5bGFxZDwaSx0wRddz2o5zGvvvYaFmAkEQLu4lyI
s25G+8JP1oMBaMJAqGNvNHtUfPDTtnDQPGnu/HvDH5XpGl8bTHaZ96grMfNY
290gWLryQHRHnLDqT0ky6u6zVT3j81fuaeORRSfddSQ7GskMpEoVz1tW8Wny
p2KKLgb7ivHFMpqpqibW18TG2K5YsRff6TuajEpYcXIkQqCeCiHxJaZDyDZg
BblYJgTSpXZXvwgRbYfx5ocuut0s0iyZ3m8IurX3I2v/anc21mYFF3D2ZylS
S1Wtj7cnz3hL8HQtzaQaemqJ2DIwnFZeWdYJ7Jld8TgBI3Ejd9loPz+ZtPII
iZwZONcqgmRzBOeZ7GN9Imi68DS1d8QqOtnUGxcVy2jraRTzZBaUMFlq9GJ8
NlQPBLl7b52up7+bus4R3fEhZLtIPvs+0tfpYtKXpT0yiHwVXxTP0edY4cCu
JiYDaoSgGsHRGFHqo7UIn8EEl/S5DpddoiEKcCC7SpjfFnBa05LzISz4LWF/
Ao0qaEHfQ/7JApURY1VJwYzxOlUfzmwrR7XqNVw/ePTf7rp6UGOgMUQ5iFVa
7g2Tr4/Qv3daVz7k/X/ITPXUntCG1y7N9gT12UPdSFTj94u+QpWWtubt2JkH
fZ+2XOCyjq6NlDwS39ZRdDPJ+vWYjAt3v7ke8kI0koRZ851uZtRNAVj2CSn/
KN/OOCEYdWYljkQiFoLe5BGjrPaSKpv5QCWhWNYlaP2J2nWhirs5umodP6ir
q9OmVT6tq0j1T3uUDtT+l2q1O57HSPg4koUNTvW9E8ZncmtzTGGXbpV4ucAr
OzipnwXvrAplu9uE5GNZQvsRhWyLcVQ5Atv7tp706mRxCBL5MMdAQ/1RCngJ
0GQtprpFMffSzZny8Psl+WxRyfPkTlnGbG+41U33MgSaCX6MY78rVfXeOz2/
XOXO4yNvxWz+RZzo6YiXKDvFMi8xcqyjheNYWqDuzvZ84jDSa8bxgBI8Li7S
jQCNV0ZMBT4SN673VEiR1QZ9TlprQPo7mcRQsHsQ6kQ2SyeM8tZOCkq4XR+Z
oeYYHVpQDuJOd1g2pC0oOO+ky4+rZSnpwlf+S1tuiUn2CMxpeiNbGQ8AwWM3
gtJ0+NU9VgYJSd6sZUWdbop4Lz9NdO1Z38pGgMN3e/yUesC3AtC2JSKGw2oh
KpplTdpPg1G2/pC2Ey6N2Z9/M0FPdpZ/q2/YehQKbfRjWFuRM3q3hG/aBOUF
2MHM2iY040/gDHpdy3BL3+u0GDLZyYaXIbTbtrHKxUNlhokHFM1VeRFmZuRj
a/58ZPK3sdcZ8NHPBPIfcw/SRMkKUZtSGHS1pML9mjbi7cKHz06qarPRHYmK
cu8Z6aICZ348BkhuEBZro/o9pXCl/pIrNzBHpcv4nfyMyurBXg1d9Tdv900N
iRU3pMBuDjeDUgiYGauodANB5gC2yW1CgvWN8xcaVTaKnX4QRSdNbBgGBp3S
EXyniJgBHihhB6lOUe5JrCGReO3UDVsYIKe95roJ66s/RtyKw8tUfCkkQ46V
PU1OEn+z1Pf0rvu0RUaPMsXrnejUy12pvPHjJi/wapCQ0JFzJ6FbksXDb9Qi
STfTyX0OurXE/FZlJwpC6WRjJu+HWqnzoO8W30A2MnS/K7MTilx+vp6ViP4w
qY5v1Z9Kp+yz56kcCenNY3N7WVj3UsMwOeM045pBwPS6oNznqkr5kJqXdoK/
ik5mvgYeHVFjRd2gr72QZwlb3m/kiP0VnGoI9OwaVVhtxSS4SAHURLcUxCNF
Kq43nNw3wgbmM/cZZ9jwQN4juh4UuoWOg+ZR1zA0IE3Tz+VQH1pv8rI5cuWY
luH1TW/73EVZuP7OY6PzQ6BT7B5xpU0fapWfEcSiPiId9vgi1OFyEW64LI9g
YifGGqsDZxi0oCR56+C7ir7R/J2niGdCL5cFfISe6B3UtXhVlREgLnX+a9O/
EWpnqi8Urd9t2JaWZ4h/kdOEQJDxhcNlSmAURimq+q/aUk5d3TzxmX/pGdBy
Ezlt0cniDnXrq8P04r8DLtFRR3hVe0SUvB7wPZSzz0SDt8XN3Kx4eJNyoQKT
3JTenQRS4Opsw5/Qt5LP8S6unXBseLVRPEVq0MUAE6U07aDyU1zcEIPOuhmG
ZB+crj+M71XhctOXC7yZbhuhZf1h/yWEXXIZXTGocAEgiM/RUV8Fzs0PyD05
PsU+oTJxFrAI0+3UHO/+DVf9GYHz3TxjWOP90aS7WXuSn4R0/Un+oItCLKB8
/NrXv+OAD0Ni+KYuUpLsoLmp9r8eUrzmlyMREHqjUWwQktFL0MkUmjjfPHbW
MhMjuUfPLYRJrKVipgwR8JIOBlJlgoDcwmyZW3r/uvvRwxG1nCfHNtnr5Lv7
pu+qVVtOO9Phuz2wj1keXIiUKThG3f1ymjshm/XwMfXa33pqckCFGZMv85lF
0HGzC2qHhn4D6wa6lL2QT5tgQtS+vedMPgs7dIdU6WTJc7RhytUwy4o1CFPu
iTGZY/ppAjvIYwKoMlF4o/H5UVRo0CF5Apx6yJJc9+zmX8HUVJNLQXVvRwWE
BR7FEVRZVLZ6aNNyK/Qex6xCB62D0qSSDqVGJoZ6Spsd/nSBHuZp0MGmjT3a
soloofMr3N6LUFHOaFqykCWaJ0WeT/NCZa/MoQGeEJtlrCHs8nS0dNmuKnbn
HVVPzGkrbDwPg1ByTBWBdkbeRqcqgzUiwHRCm1iHUwszKwXEeGRkJE3S9T3M
uRf6HX3rKmBFbMIalfzCOOSR1yIHRIhiGMWTuE+Ou/7/3n3+FfmGG6gziJv+
MxNNELMSgO5ZSYk0Q+YvPsehosgByRDPkjjzurD+PcNy6Xf1uSCnK/2vl7Sk
R5ChhnhOojdAggKlacKSGBZTg9M4jy05C3Yy7wEwIfYLqrt0X9QDF4PubV3+
X1KRq+T3gD7P2yjluBPPT/3rD35VnekShHTmnepKtn1+S/HbHN9eiKCoKpfs
1IYuuwImQw+aMMbk5LFog94m/O1WqLXamIfcZ4Nmqf7dRUXgtGnS106iHHZe
VRt3OI+tcrTPua0e0lkPLZnERlSUlp9ow4h6mpL0ExHYWCVSvGdFqptqxSUd
loeK0A350YgCOVcSBBFOcxe25txqbORdue6UF/8uS2350yohQsz1JQmmHBf7
2tvAJHkj3GgLtjqXI2SqXxXq0SG9/HhK0kKs33EFlBobManwQK49g9h980rb
qaEAICeeWPu4wTrl3sVlVCDJDaPOhpcg6rDU/+3VP1lgSw1XYTLibDTdCe+N
02l/ZU8B6YkOJzg9spKN/flRlP1U83Zb+LDrDyLuEXGS3wTMRsm0PzRCXlNV
u6XIJ/QUnhqiX+UHBEJTPj5ETmGLUiseTmxVCqRucAcuZ+nKBIhkRBVv49sx
GN84NDl9crlnHVQ+LjLBR1w07adWIsGgT2xVplbMpnNOpb5A7X47IPdHKCiR
VWkAGwfSIRl2SvpmbWV0PcCS+rSQ/AHaZN5otn55C6Kj/LCWdFXBAW1YEdYx
tnthkszWGE9rmjuj9WhRGA48/XVF7knqBzFdTMJ7lj+1D9ybB1fsyagTxm3m
Tpi/XMdeSFX4df9xSEXB/e+7ZwL3Daw1eoiCt7xKj8WpPavDOlpNzNQ2yKXr
wd4d5nxlHQn7ZSHuBflcLuARf/5SrGlVFGT8SZ3Fs4tY/yudhd95A4ydpuk7
pwxuZoMNHvsVhdrUUh4V+h+mNoJKx8uzxyfYN4unIGx+vIai3CrL+DF03FUq
8mr3KayflbVmAh2nd71bhrYS/XVEJgk7WpX2+iymw5AkYNUUmL6OHVhcGpUr
EgHT38CleBfAR0c3rBDZLb2HImbYPCQ7XH4mCWzWnUlN7eI1pCZls13OmDnq
VbTtAliMVhp6PFWaaa9jbj2KZBdhugy6UB327nLl0XKZ2l4syYM6S1vjsi/j
sFS7giV79oVQrfEzDv44YTi8bgP8P88KD/KNvKobWb5l2Fs1bCKlIp5naf2e
SAXkfDxUlXbM0Y2hPCGqwBI8wpQDoL1ve5TqLbqZ8Xuc0hSSimOeT7q6UB2Y
c4IWMO82UBXkkQFtmRMY7mB01kN6dWeLJ2GOGMWygL7o+ARUjPs2uO7dw56h
KUDkvT4giGBSZbyd/ryPJ3UmfMUP8+DaKi56orp+lFk8cM4hwoPjx0KTTlzv
LEBdKiPAqZjoi+ewfnbQ2suIk2TFB6KHAN8CWRyDwHGw3uYR9XINiLmO+QJE
5fOPmBU+sM652xgdWq0Cd6VvraGiTtmWGZwAw5uOfBidNZjSHQH6ObCXdpyT
i1/sB+W7sS1rCPCcHpAfrcQrJKzjo537i5PogydMNyVQolRLG2PNst6kpjbZ
Bb//ePoQDqX4XdF7r6g79Q9KHLp6vOfBlsz0Ne7HhiAR/rXbgaE/LHY21jyo
eORPX7PyT1JBpoyBNGmOfs3wqIMSRXx+bYQ8SnDcw8tCoxdAfpzOg2teu5q7
tEWuS95TapTYRTs2xwXGERl1H/a4QCMPX8KyohJI0CnW//LzcdM9aWQ/jDZ5
qXV2Vlj4LHhMa3YWvyV7gQSfrE+li7b+dxeZ5hkwKwqNXINgjJJ7Y42R2Y6A
Y0pKC76XoxwU6z0N5ywKXb0I6VRs7tc/E108ppebkc1LhIutbOAy28kJLxSh
LQbWdNKwr9REVv4IQk5Jlq6XXjcd7mG3sUiu2/jWPayDzAxLsNVErSVjb3R6
6cmp4JoXYE0Ho4Z8A5T+Z0aY19giwbLFOR8N0L3kYuN2hXNIMB9PJVN6ChaX
g2s3JG/7PuczhoCfOq0cl4ZOvlvqxVZS0y8WloZiuf4C6i/mjX9o2Fq7N0zY
Bo6ECjmjehkOvbiR15So82jKtu7W1SWUsaYeUg0AYk8hIMWWzQC1vQNE+GSK
8qSD3qsLJePEzuxHGZUlebq1MFBkkk0Qn1rB7ofxRLGpuP+G/xMhV59SHVI2
SbaE6qw2na/a3uIDvjj/IwEjKndJkCPcMPmoufF5y4rX3g7OkOjHUvfIFhAx
thqwv1qv+HyVjdShcsdKUtBEqWpG59o4aH6OUAs1f3GbNZjFDWD3Q8Y18oE8
Ntt/ff+kjhA0RkOgj1Zrl1fEyQ34neYhC+zxTCsEJgo4od+F3GPsSAlaaRar
HFEXdsfF7z0jTbQJpT+n2sEMTuXWGbufIOWPgPZHk8kGBkoMJ2FC4fqeO2h2
DZreuWToaiKCeH28nmyvJFGRQJ1qabiZY7b5VlrLK15kncMmmbiwI828cYvv
epEix+FKGYBgQetq8RdFKFC79DJ8VB+qU8Jm7PLrRbhfzeieIHIQF/kIAHHs
u8bTznCs3LlfOq/Yw0Io4eXGprlM7JMoiYbuF9xth12nWmc+HZtIkUGzhPE5
jFw3zk8tY+4MII1PDm3aiBLP/qwD+f1SjeR9NOl0TyFLfUBQZhHxHbA8j1Dz
ExJYtAvNYOzUAYr1I2gW/07RKWI0V+YFk9VyYRWrU86h4JgPwueYti7HQTpm
qGC09McODZ+fmNJAbwYSymljyc4r8dDot5ySAaPi0sSWNjUBDZCb7F2JGKa4
78y0RJELYdLPvDjkJ0GTtXaFdczJ82zvuoFXb/09i7F6gtBvNBQo/Bx5bbwj
8gxQTp9rc7voUScrxwHUaSCic0G42R2mToowh/l2gFgC0M58oPf12TyzI6qz
Jv9HAM4OosA/f9h+V7S/meKUAVA0/KA8eoGsiFPW3hO+s+3c0ZGB7BKAnMz0
1bZ/5LLF6C4lWu0yurgAB5nKc8Ble0q+FuuZRs6xNmHvkVxq/tuiCreaVEyi
9JFd0HkFaMcRK0o9N71sL+0HvAAT3GdBXtI8HRDwCln3xVFtIUUfZngksaf7
BPZ/m9EGYbVLjEGiGcJ7TP7Uu1hZey/t+DpSwaNEzMfmCAV8oafYb9e/8TLk
+HspHaUNOd6pkGTvCXT5Gw1GYgERrPa8XGdcg4rNBI804YjExVLmBOoQZjRm
bae63iaDymovOHii/F+eO3cVSg60GMY+lzad/bGY9aHUa6c8vVTo+hgcsHvV
gBZQDsQXSMyHzvQ41GUTJYdNNvXlMNeL8hxyI27eH8FYJEp6gfs1uiyO8id9
mHYhYtxiu7VtBIHj7Tan106pMlefbCn45a7dtrcB7nmSSQiPwzXFOlFSSPf1
ECEltVR/Qpf0Gp/AJN2C4oN633cUch+ysXScK7YixiRv0Uc8Sp5eaG1kw3bl
eDD0ozK2bh8JMLK76GneoAk2IFYyNztaKtLqcirTVoGB8R54EEPQbDJuaeHD
yCEZxEgaebVMkjmVyDGlcJpvxHDKgRFBg24J7XvUgal4BJdBGW5qdKfDJE6P
/253RK3yj/8L332+fXnknLSWoYzN+bHhBGlMkf0jDjUGkJ2qnCQVqoIC/wHf
P1z9jpNeM2XG5fc34rSVVX9WNamKPtUz8N4f/0SGn3p8IbeDGRvFGed8VTDW
+ifGYbGHbVvUaHdqnyEzFkgfuBPtf7j4l4LcyGwotVEFOp3dAfGMaQJbD7kl
KHZrGf+1PTK8tLCUIXENpXUQAQDESRMqvG9p5lH/QWteaBXxXyz9t4ruNAka
WcEtkB4S4gYjwwHPhnUQNRYa4qD2m9CAJ6Vpv6b8gnY0SWShsd6mpcaMhYAz
I6QcBmt7+Q8wjtGmKRF7KlwbaaztjXF7W4ybee/M+TZnSPWqfRZ7pIhoLb0n
61kf8d6iaP2p0UpbB1/9DHau3lXIHJWt/hhWqAO3/hFFxFVZ5UGFq9aT8dby
BXOCtWfP4AtmpAEphpWkhlG5eMZnPHaZ1P3fQjcFzNQoPbr2q4tpPlnkXM1J
goSOhX4Nk08ld9fx9KAhi5ZKBLt+lZjbOlqPwEh8mfFPet/yArm7vt2LAz4K
2/6ykNphsLiP/jrxZM2Kf6K0HQ72s8D1UpKnORUVT5tssKGaDrU+MD4js7aX
CTEyoGeqX22eZ1/dSIEYjTEO42Ybo386WmdUw2lHXY5kX/qqd117BWodikr7
ZZK8VDbSrjwrS9dOd+YQXKGiwaMEVNJ+hyoDzCi3NeEMcVButCfb4Bk/XB2E
QwF0hFUd6zo9nm3eK9Nqco+pTzAE+LOlWgFFCg7jxq1HjoNuxAzW68JLzRHg
8byWxD902MY07uYjjzyLY++Cs1fjQrl4r8jSRWxPuCofKN5AtRaOoPI1c1Zm
8xXRjokT/Lm3NexpatPgcFz4EfN6/WqzjAYGUd54kzrwEQ58WBbJSSGfi8ql
EL95gb428QU5F/e6OmRyVs91MKhzT7zLG+ctclgYDjVYnlySmMM62+bHfaSN
M1Y3VwK4YDGRo1unb9rApy6hZCfG6Acx1O3ncaDlvlWwtBjhpBkPrJ0ZS7xq
sW/84VB5sv+pGChq2eb+P/pZKnu20DpXJMI6pnGhSRNldvcxp28xjPC5gsx4
yhaGKh0qGY9aLKzeysZaFRGQpt9S0KcwkCaUI8ODuMabnC6hTQlTs8OMw28U
BrlvYoELhB9duCMRy1lOIf1Eo+MfhvoZEvmB+bIcHgHE0ptA52nj8Y9P4RfZ
d0ULQUac/KdvUhUUCD4Q5a1RrXyJ3cL5Kg8cJqHW1qxlYK960I92hwB9OFjI
otCoIhhzcfsiQVfHfIjm5EaGyKoDL0RIdUNxkMrFJ3gMciixLwbCBFH33Lds
mgTZBPFmBIboHgpTgLPZDiusD4CB9LnGVqoOmKyzOBK+Z/wiPZyfPO5FxWXD
VkWIOAi74k+N4HAV7zpabrPKYNishOavtyVFKUMyFjwwcJ15GOKzTwm0FPLQ
MXyK9UikJkmqSHRhtpb8CVF0ryB6iN3wb8QcYKUJIWGVRRo2LDqwoe7tJCXV
/1btwbtjqFdVKSVTvZJMGR+iT8anFbtNs8gDCrVNDGY+wolUwo4qAvqBc0u8
Hk+ayIdVogRxotV9q/UkTt9DXp44RuLHN0lDcpl/qQ9tIR3GO6k/73KSzjPp
26UGK2MLG0jQKP75Vk23KCgk6wyblSio7NKaLAoBhLcDMKF52ei8JKXWQ9eB
72laP6bLc9o+VIdgL9ek93XDhkhE1VE/ypn8HCUqVD1fiqZT7lFyJbK5Jrv8
fQ/zvL8W3HCPkiJ2PIHlxEsm4shlzjvRCtbELzPxLkOhlfeZfiLJJ7qePCYV
18avPQ8KDW7b/mOlb64ahk4DxrcI8/9r0VMNoykK+XQ2yV3CW3OyIeQK0Awu
u34VOBO5J7NR8iXF9Llf82TpmQn5j29TvcLliABwkWFBBC/YN+l7rKgblGkx
9DXIW85fq5O0llbG+qmqh0+dGjpUlYFgeKKebYD97m2OJ0NxG/pOqfoCYHTH
pCEblCDOitO55Wom9tJcbi4hHimjMZ6W+/F/wKzvbNurX6/F/WQ19t2MVCvb
Q837E67tjugfGRpJ3u1sxFaZwjnhkT/gukcwuPE5+wBDPHrhmDe9W9RfllpN
ReZSNFpttqswa5wUNxOalJ/7P/D9nZuitIdkkKKL/vNSE7vhmgrXsA6Cuq6E
H+lnPldTZkl2ZV2TOOYCY9F4NOOOsimU0CYwC5AzZWWnxl453l1/rEI66odZ
I+lZGzdq38ytSWvjW1bVPtkbRByOw1qkTWC4QbvmCqU7STJs8p5GlsQtVHDH
ilXDUOyDgGovGxUdV73SpQy5fAYH8hY3+O10a6AsPC0ori0vB3mIrNaa8sAq
Q+mL7EDQjUtv2cRYEuncz5PSkYL3Q0wymKn8FFlsIGgoIpGuUmjeUyqTcuB+
iaxb0oaDLVvtdK1+3inBXZLjQ3STZmEkFHDmFIjsYR3cx3WzxXNy8cNOAmsz
qAdaIQkPC7z4Nw+QXHsQAC1AvDEC1gLYMhUxeH6bjNhw3J9S2nHAWAJtU1Tz
QqA94P66QNrKD9frjXNLOCre9Y+j9rLXz6z+cQigzJUYa/Sg9NSkQnkimMn4
ITw4WVeNAn6Dp7C7FQqvynRGWkL/jyFDHVbKl1q5hbgsN1d/EknbUkaub/R/
hRnzcA+jptvXgJSjrJi85+EVhXQozZioQ/OTaC4Wzz/dIIfirI8KJIYSTOg3
qR4OjdzMcI33bVYEC5/EE5w8RTG0VFSFO4t2WPI51dWrbbqkvO3Z8w80pqpW
g2ytzuxrh9p1LpwVqNH1MkA/ZyLNY2VNlqDPQrfe15LNiXvrA3zj1ypVTPyU
cAXVaKsXGnt0Tc0wwXN6nroeBRJ8tGWgaloQPP77NH2zyAVEWPmJunOsRhwg
/Vf+CNj1asVIlRYQnEFdjqaP3/BcBaMvkzf3lceIHrKuYc8ngjAWE0QgYWRT
MzgzGel0OQjbzpC74sYthNo3gz2xepDunGBD93e6J+C47xfVRbqNbJ+kAmLE
n/8BJlrtB/1+aflmzjvRrKZVYx2Svsx+FkJa7gR1qN2pb31TAy6k0cjQzxi6
6UZZjPFYmUbZ6QEpw8dExnXylcW8OiGNTzYzn+7cx0VI6Um4gGJP3aP6sLfJ
SEFb3Bc2myHa+cC3q+IpZ9HdwAgtq/lX3AxUPTJSNLJg8l22DHXG0M3Y4/t3
7dfEidskPjYZDH/2k3VYs8HQZLfek+W0p6hMxYmGOE6Fw2abUpaEXFTWPL0a
lbADlMYFs5DqTqIn0Lp3ntmTF6MBYuOhjEetK6aa/voemd/7fiIYvqXu9fOB
58xL6UxqoG+rdW5Z34k2WlEW/sC5z2ufmd8fb24VICc8G8ffC76vavlZEUPm
ZhqaSTNK1Swwy0f/m78HV6Q78YfFxK9Ly1BVRNR8NdObcqpDlQZQNBVgxGsb
lU/WjUlONLb1tYaR+qYWPqfaOC2qvExoUE4s4KM1mYtXMqCFany3arW5AMrh
2Y3o0xULEh9RstsqKeD7XJdGhaZFrztcg+TNqtI8qMOc1KWB2a44icLP4oS8
SiR8qUHjRLIBWlSBJSXqWT1PtgSOwzed9jbBwTeaCeMq5+hna5vi1rpPUEbr
vj6kWYsMJwvsaSD+4x7Fen2loF26EUmnF7c618G/MkpfvTdFBJ0h0s3yXyAg
jwmli5vlIfErRh+AfR6KANiXWdKFL4eMNiUlim8BWX5g5ADMnJ45vnHjwRC6
dVbV9lmoSVifSNTkWESbX3yqMpz36hpCoA/7Y1TIbnNHPli7LNWNiZjuQf8x
jZWaff3UCN4cJIZjELdkRv2tu3n42pAVT031m6n3i+0v+s46LANFsZtx5g9p
OPbcojOen5/mn++aPWF3XXYJt8RHghzVXfeaLUSrAdSX1BKFASEuuLU3Onea
9niARM35nip/LOWXKlKpoubGSvCREGYqPv2ZgzL75CNA4mC7nqAQ8iF7olmR
kbBm46/cHZwzukXjR/rd1CmNpyPXiMDRTNMzGaNCHl0IZRoKIJuBATmb+Clv
n3Lo/m9Act2huBDvlT1UueybZIqnB7f7bScr+fWUf1ihr6WQwVJVuXFXlmve
NjRZnnUyf+dhTzE1l16CTYoMVBVWFG/jJzfgITExhnvmYwNwQr1DNBW2sKZl
Rp9lsCl228t2mIWwODyDtTMDFOnrloPaxa2GO9hg3EK0TC2Jshxc/Bw4UaaB
OIN+5E8PJaK5Syf1Y769Iz2qSqL7Kv5fkSWps3Ddg//IJhTEuuPKLnQWDH4U
3vRyfUNPTYLu8okifk2TKDgpj4ikB6S8MqGL73WzWzTQ/hvyw5GYufNX/4dy
Q4rD2DFL9rhoHYznxyHM6sLs9o3Wa966lryFWvW3sE3zlZo909L10UBurP2V
CxFOpXB4p+f0e9TUFijqWDp7t+2P/XGi0QB0CIr4TjoUIBmnfRbkUX41cFvb
4PMscLjscMgd1kLdr/YwVGKu5QGzPdR0XzfcW5oXgYazAUdWTxDcaCSCkDgu
rbh/W/86JkHZEB72IhM6LUNZTC9VR/lY1qVfCbfOcyJritEjRq6zGWZplLek
ilBgfFL5Av2HhcATfPWFfd3kRQBSImE5m6BuHITPhTdfPstj89pN2fyTFLBi
50yG7FMpah6PwLgnIAhD+4ufKpzjwFWHgv0gD+wJVStCtP+KIKqlx29bN6n8
Fb+qd81z3dcDoimpozfM0E9FbD3TPvFT3NWONPuyAicmvEAJs6/I86tevby8
YsjPdYUibmDG+ZXaXQNVhHjjDrhhX3cE1/GhlG6Ob5H+o4sc/X/BvtS7LrqE
RDx5n/wnO/rVHKDLWczWCphz93vwcsTBA4aHpDS5egqN1DbO+eWlYoEE45gi
BJj+zr6+IrUdXqRgdk6DHSsYWLt2QjO211ZMToLcVB0eFKuv5YiyF7nnMFoZ
oOH+KNaTfCvPkzvr717uD2PKn2iwnZIupfYG00Kad9V0aRZVCmxy3Df6Y0+z
CCpTKPImnsIvsa1buXFKCjYf+mCOqDcmFBOcYNqAptDN4BP7JZa00RAe1ASA
MGFR6We+QDFCf1cu9j+2FPUs+GenYkC6HNFWUgI0jGzL9Htx2iL0ngbtEBfz
HPCx/PxjAnNdb1alJMQQrujuCgNHyjY3gftJ66iKTeY39maUQ0K8JF8phCLC
eY0ler3wom6wWn5IYQTviOFUxis7Z3NqPrDD5HAq8P2rIh2D+jQRPsygs70w
6RqDX5+NN3YP4HC2EXmRHmDkl90QiV9fOvSbqfh5ebkb+nbWi/cLPXpRkGk6
4RMdisoG6AsbAMvaTdR/B8auIBPSwCW5rqxhLkPQhoWzH2opuo1gN/m2NA3E
2Sj69Eb2Vf6f9TmucAxkImuBMS0MCcRuGpeBotvzIBHZB1h424GPNZVK0iL5
0sFbl7fuFyBgqVKOFIQm2v6gQWr963b/B2gMcHUjO++p6iT+Na2vyonMqxjg
dYjwnmcx1sRtio5qfjjhY1w8YhMvWoTiYjFTvC4DI+b9lI+EVUuOa7fOdWwx
jyr+uC7aQ09HfVBDGCL9CODFwgHAXWddh0FHDQZdfRHLRWf1CTK0z9GOu+ql
0yehTogElfgxbDjkCtcuEuL7A6RuLTQQYW6GqVBcChkKSmWPnP1KHPdWf3vF
Nkd3fyRgE5Se5qCfjaL8RTkLxqy79Lkm71zT+Ay4kNa57wT//Ab9T9mjAEYK
JCQXBggzG5AXrzDTQ+ul58q+A97tOnwDGDsmqFLidjn2RMWxJtCMRbSOEevv
o7PeZcXltrw1EEbnd4U0qPi8DEp8g3wlUhCWaxYitVWLjMZfth2iH9vDkCyv
UZsCR/CjLa44xmYiwTwb58v2x3zLN5tRfGcw28dvDrqBQP7payI/fhkFKs84
hgY/uvqCe/CO/piTBcB/bbwH7LhJ9UxjOz9ocXlRAdeQJP47GnkoBFJ46u2u
GjTDx9CSePoRcyzFE8mvcZQbYMppewv7rSDwOc3z3u0he2/6ydG/wWSCi8rM
vVMLpJ/jJx5NYCvpB0eQwzxFhiANW0utjipyBJgUPSm85IWD2zX7btWA8lJZ
ghvQRpZ1ZUUfllDf8BLJJc+Sp2KG7aIeJwGitI1xhXWRQTJ2suL7dUjprHZB
YuntiM5upL81b354Se5yllIURQXCXhgUcNTSYA/V73tFzMmZ8ypf92+0F1lf
f5j/Gp7eqvVCzK61HIgUW7+5tGuFMCqi9HI5MtEj2B8tILoTciJ9qZqmh/bM
LzwrGbenuw2QIHL9oTzmp9dr6fiFXnruw/Lb/wYktuJPW0JiHtkyoJz1MaFd
f4OTPbTVqCzPBXOMmNIbiBaLdfG5sGcqfLl0QaTH2jzC3kgtJ+kIo4/2v4OM
4hEh/YRTN0r1/YA3AeR/p3NDRN+zI5Aprw3DDgJmxi2CTqdPyNGP3YCeaLCM
k9NPKnBHYOoAXoMbtIYF6X9hA7AfTPyUWkjNbrFL8p+DCHHGgwK2Yx/MoBnG
8n9aMtA6ESMRKkxTq8Iz4dgIUV8ZvOfV0oabmUf5g/WIVbKxy/kfCYhyTuoD
8HxLqBB3QW0CEId1O4c7MpYq3p4ABr8FjHRr/IfxnEkXqkZ5AJg+pKACZe85
vAMfgJGYt/MxlFu2tnj6F46S7uF53qNc4xpzeZLGlMdCLMZYrdBTZBe2Ubl1
O9rv3ZwCrrimpXnkqwf4DXd1BFECeOaBdXCFjBC7jqg9wWRK6NsL9llIuq6f
Om8CI49OmhR05FUqw7pM3XmJQApgieLDX3kotFtesrbGX7KXUkfm9fzXzQ9c
4K/2bO9LgDmnoIWrS8NfJjwVRKINvmBjnnNnEsRxXNxdYgWTCbJt1prQOSqe
SugE1Ka4Zqiac+x6b0WQsHMU2hgRgr0+4jA5y2miymisjPeyArXXOm8YfJVo
XKNEkDt7kHz8QxIc1HTcsP96PL1PkHH/dHI09xVV7X5NHWU60EYe75Qqv+TU
y/krl6wuhv5Ao9hbuhWL8UWoxzedixUg/ZrLjtkpVDYC02pVIoExsBJFgXpR
jqlnbsUaQoX1e56/zQh2ZuCJd9AaqOSEoMd49TathLANo+wXu6ca/ukRgpDk
Ws0qYJnoqffeAmdEtbN2Dy5fKdBZqHQ/LVsjljvP0hPw3spuFMxXAM3dPPBy
7coVchoMckeK7qHjQkbTB8Kk3roLwKw4kbAJlk3/WWq1TNxzUEstvZMAbhtF
axl732g0v7cbg+ACjNqsEJCSsoHnVEkfJscdaH4amK6nfHKXdfrqGE+FCObx
f5JrXs6vevdjYH0k9sYgShNxx0Ihmi4lTKvwpYuHdkkiMtRRfi8iDmlgqu84
XjT7QPJwUVBJqFO5Us/UsdaV0SZaq53IZfQ4xdzeeECgcpBi6ZdzYwg3lstR
N/juYWDZTZMdqfiSfa64YXmrdvbzXAyCHQCHicjdlp9iXMV5p4Z22mvIebMW
ZOIdnBtwVB5q8O6v6mfoJ3sJCL+XOOcIZYgqXI940sX+qZGXKD+YxKTKhYjL
O8/4BNjJK6SzuoZAe7k8jc1APYblwE9q507gTV5tIDd9JhXNB6TLtMD2T05g
+uUKxm2TAzJJhdRYfw75+IyvXd6BZloEKRRM/5Ut/JseAAJZGBS/qKsqr0xE
OQ1/UbdDDPMf415Nr/u2FDuIR6NDQvGnnRsQVI9f+jA9Etrk/45M5n8oPJ7v
mgWBJpQDc01yFwCAnB78FZwfi6YOKbAnZqtNSPi+Ct2UnVFTC7p9xj7uxAWq
GNw2OJu56IW63AOrTWd+olOjYWmzbrW3NgMqwiErF1uldOcq1zqAe42LCrZI
kIVoaVEAh4VFPfig9G5gji7vqaYnE3PWuWGe6jXxj8AymKpqDPgCu/gANt3r
IWDl42teh6FxvEJBmLrfG5iFGqhKddFbv93B+7Chh2ufjxqFjITDVoNrmpmW
h8Th3Ez4wwI0fMfagdkLrRfnrxir4srJ2Hs1femoBuoNpoEuhs7XdyXVjvqf
8JaMSDg7kn1Nzr8TOej9c/ouPfVMY24nYNxynY9nDo9fl9dDtvXyS9Ubjz9Y
jTCPsiGbwq6Y8q+cVCpmBGU6GCpqUtVyAjU7DPtojEOzzmZNfXEDuVptDnof
AM2dj5KBfJ7MJ55BiuoJxCCnzIbjVUPfKR9BhwRDYiboUe1WpNMd87zvOohz
xS6oiHVMzmd2Vo52TcbRsobVuEJDdTCRFZG9+gxThPybIpMOJN5KwSSPpWmo
AXQg4bp/9SZ9TJNlfjFfYolD8g80r+VMAdSmTZpUrTmVLokS4g0IkwDiCh89
zQzDWzw6NgYLEZT+HWdLOKSsAk4nHzh+WPHJCdMNLXWORLSXkGVNkbc8v/k/
aTgmA/S/Jb0LhtTDYjp8Gf7SbMkagxyVFfCsVPIGN5a9LFOR/YbJSZZNjbfH
ICziaF0fsBIJDuBNy8kX3yXMPPttBvnHOzznLAE4m4o12cALolVtu+nu+9Iw
jvo06iQ0hLKOjJp57TkSYd6/SyKQhTzOfsRS9vEVmF++7UZQXQJ+ROoSQgRm
C7KMf2408+mnEZbyg+ICOhvHmg8dB74LL1uuL+gfBBFir7jI+3QhegFOqWgh
LlT3nGY89JZs6riXxdAt0zUPLNoES72NzfaaW99NK8e8JZG4XdAKz9GJIrjh
ugkYL5nm34xpLh2zAc5r1u6Dv8t2SLDAxl6itJq2KsTSIJq2tt92cIx+3tFd
/Lslq1y6E4AKZa8Kbb6yWWv+y9WfgpBJnw6FDko9SCuml3dm+yGrqDcR6e5n
G+yvZFAowDPG1jB6csilEFIMeunTEnB6nuXyjORMfwbNvPG5lh+uvO7shoLN
ZnOFGeAhzWYJXh47acG0UMRdRkCyArR9zz/dgWQzksdoseqGS/NQxbLQKW5b
gePBsruzmN0hPeIfNJ0NferZUarD2bMlPl6vI5uWmBdVwk2AGBhmV4N3eU6w
sSLAi9+kidknu7I/02eCiO2y6WnFy+DqA4jfhqANrisdhKTHLn+7UFEe3qYC
5vas5LVrVHY+YxG+XBd/jR0pmIPX20FxTlCivOl2aNUT+QnnnEdSsi8dGzJa
3h+fnRoK5aO6mniSAnxblCG7vxnumlzJh3AUomccY0j4aFtipSLtj3dfpDmp
9sXnJM4x8pMdw+nN1u2wRiwIv3vLXI69qCTi5+6WcXE4nJlh44Xk+yXaiZRT
gwbRZgjhI2SHBvzLSpevr2OyTMujU/1gsw/AHULNoGwIKebgDQAkT/3S/X0Z
3aZTyvj6OQNOfq/gjMGrnk55tT0H3BVWi4e1lz7JMWvaLpefa0SQ1CrvQmAa
Of/FCpd1M8ylJlIKi/Fmq9GqUU31MUB+AEF/5HeAu/qXlHgF6fSZ1wur7INb
rvCI3pFtaNOW3Ofszzz/0AZDbvbTkSPX+UlbUNv24kwqkIACZP77bBdRcHo9
XTUm85JSQqZK7subqWRMkEOcIjuqom1kfgDIeduWcptDACztgzKCzn6PSXJ4
SGAztuopo6yobCytQj/Xq23WXqt1sQfEGVe7GPhzCSTCyWxTcYHXAvh3gFX7
rYuFaFzNntYFZYGPjF+xlIkkWwvAIhC/P5fTQfa+c/QxZTire0vuOfoL4j+1
r43m8Lh8y3mLOHUtRNMzLNR1Qapu40cdMXg2dIYodeA9wgXwQSUOIDcgyF9h
ierN8RI2OQD6RWycnuQInDihwWfLnGtI9JXQkyyR19QDBXlp6mVXo5ySKnzn
ZTq8rG8B3gfX/KRLhGRRtnaYpfOCrHzaUGNKxpukaV1V88T8EVFF2syMCzkN
CLpKkf6inRGm4BKtyPGDc5h8Xn38XE8jQ3VkhUNqVa01hHs9dhTX4rDEqEhG
MLYJCy8tDDrK1uRxFYJCe0/YB7PpYOBExYi985iUayz3yNpskXirxDGSg15J
UGkYawfrqQxEp/L+NAP18Fggnas9BpuP++Jn0IUuQLaxFBd0iKy2ESEfholv
KhHCliG/0yI+HLbbiMvxIGA0dQFnhuLQSv/4nrgVqk+i92HpLfBaGdshMp6q
JnGH0WZeiYUddR3GWJSt/xDF/2BCCyygHNB7TKwApLXcIciAe46q2+UXOC9C
8YaqJmCu/1cAzjesVyElTgpqGw/7NjD19A7w89TFSlSlQm2n9mcBmb2vVVPJ
wqvJvGSUK97kHm1T7mfW7cy/IkJyNeDrJewoseHm9CbkINnBX+kmAf5wM09O
ygGXrFZtjIFNCSETIKgj06N6bBPBEmIjYztjLcYLuerUgLR7pqFc5WEwluhI
FnTwP2WZDEjK1o+HTUda5mhjZRamXziyZHkedAvTqFJgByE2uJV193lTYQlt
immoGCEKRaKz97MfLEYtKJgLQoOt1LFLYahsBTp7E0GG4SU31h+u9Yd1ev60
cA90b8diienDe7jd0f9xSrD1s7ABvvEvzUBnbpFDQ/3ysENc7qW4Hl0gXyO4
0jHcvqkk1yhwLiIjr/qAGGTMMj009Ptgac1nTynkZ0lAlRwnpLRLViNKZpgk
Z8mSjT/Nv3vOHAP4FG6cfSbz/vEOtktbyOi1D+I3n2SXtvyWOhtsZItEYeqR
oy9n19Af19e0H+MxBC9BPWu9DwPquy4Yejxpza0dNk8mKKcspWuHng2qGt29
JQMie2wwsWSiH8wrH/OOKW8gTbVmvgR8sYvqda/iNt3JaaoM8MMVlDYC5lqR
aka3ezjmvrUBpR4U4CPVhuKatTxBeByLWJPeC7gBv+e3ZHUc2fv19oKPariF
cmYaT2+k9cZZhNCMhnawrAqzwRabHJcE+IXxiIm62EY/evqA3b/w8yPZGSoH
pTyZJ+xJalDSTwvjotFR+6uBjIqNkjaKAkueOSXWiLUxHUsVrcgZGA6jHoDX
ooX6/ViNiwZt+MLdkqx9LYMGD0c3KU19bJIAvrazi0m4b/KxiQZ4VZ9yAb1S
QDtPf3yMIPZt0q7qqb2DSORjoGZKZSk0zZYayjxmrCDtWweQ7ou3FvjLoPVK
LyCckz9HynnckCYnh8oiTA/PsYclHPfc0wvYklL5RNaFiPRGiK7DNXTOWB6/
oRuSyGmXpfbFFcQ9eBVLyPRaNUW3NuwblKaiyfuF9qZq47nuXNqWumzQbv6Z
qyKC3XhhA1sws5t7C4K93offUmXIFKT9+MmHFpq6ioEiPJCzXsGkIWNVlP5O
1MnO/ALhn12OKRf1gbOcPKIqtaqTnWwMwf5hOX744cqLzyjiMlri4HOf2397
ztZQ7av/0xea2tDFtZsmI81gOo0HkRJ2WBkrPpo83dg6omOWZIP6ZfKLOlLL
6e3nGpin/ZWVBl45Pk08a2/OPO8EufnDa8cKXGEDWzwX+KX310b3zPC91rgp
ZGbpzHHsJz7BHykvrMeMHMqpG1ie6sxo+wbltmkGpzG4qFh/bRA03KZfKPlr
ldwQsnA+vHRtxkbWWDZPeuf+CU+scIgQVXDqxTxf6glY2rFCtLKDZOgMubVC
eVTnIRdITDA9kZnFOIxuR5VAPrdM9ZxLvXfqUdZm7v+vAj+1utFSvMKOXO4c
T9Im6hXqriGF9763dtpGO4cz6P8whJ7bi/gBqbPnZ7ULD+jMX9re0MSg4pCM
MMcS/YtWETjMi/kMwveoK5n8tuEuW5gsGXFmgAKSwlUYk76JAlZ8PB5RDDSN
tpfwlBrs732JAvcKCDHUeJwIEjAL+BCa/xSVZ6jFEJvoF+VJwOirKFazaPP0
sX76s2A86eYVa5U61tpddQruGIYJy8RjZTnkZ564Wy1Qyr9oiu0tLj8r/yLd
hJWuYRSJawD5C2jb1eWFt2fzMsj7GcOaHNgER6YGDwqtZVAb1nljofhb/SeR
AQ7JlBnIOWcJg4AK/alZ7yGaKKUiU7I5kEMreKIPtS4dBVmVmV3g4IrLHYJu
hgtsIhdvj53+cFF3A74GzhFxbcCvJy28OUX485aCpcNZJJ6t1t9xBSPwskjd
S5FFbT/x9rJ4E48GbdL78ic8itb+kMbeXauo8ZuNGomOHBXRufSt9NQrwvyM
NcEGfEoZcNYJ7isxTy2Xs1t38JQp+nS4t5fEHG5oP9vChYpWio/FTms6qTbW
oTBMTk+tYLR0vesNObRHoqdw2A9Qbcj9i6Ilydc0DDy1EbW8AXTDtkxay9V6
i0XPfvyECF6zvMPVLzqCJmhqxFItKk0Lm/3gXZlDY5ciS2GY1dJ1JyrxjR+x
y5Wy7Tdn56GQsPQxpZ1ET0jC9nqLDAfNbiT3/yer20TrtsSYexZV+YsO/uay
ed3iyc7m8kV1xMIVPyl7YfGYTaA/HvEbVt6UN2ls7PM28LfUR7m103gLDuXh
Ln+Agg5vSSKq0lMZFGhHXVF2aoHZI8+eaOKVF2I0YPI23N+2BM1ZZisWxYl+
3aPwykqX4oqtkSV9BTvdNctCqQOOi8Ak+y3Gw41fZbT3DMgek1agPawW7l03
jkkfmDmNnVM1XaPb//tFXz7eRItkWZfaecCqptW3UF1jxB5dp3gtwNBUcEju
e7UaOvubA7afPueE1W0IyuYlgT4SwH9G3JsfPDbRjjK+3mKYKJTF81Ll7i/7
vFAnHq6gFABozLSdFsdpsNMUfr0kgWOh+vKRfQ3mSMHexgAgYYthDxnevg3D
KpdmkeBb4DpJ6lO6Y5veKgvT8zgwPnunnDicuxcLHBzzdd0n+EWmmB04Xj92
d2upsldCgXDIQbkuoMgVsuiong0gB/gLlLDEuyHaodNf5TAfpmwv6KUUDje/
IEYZDbgNq464njnke27g3MIxh7KIhn1QdrsRQDByNvtN2fOCn/uE5A5jSExv
ykdwuSHrZrYkGOeQhCDhKk1Dkea28D0XpVfCwexaLPkooSxIJvjiuR7wx2D3
jdUoplkzftwGo5X+Hi/jRUUiSRjCx6OZ+3eEt0bxf7NV/ztUWWWnS1pjhod/
sY/scsBbRaJxYzqnoXbBHdFmWxSW+iy5IfNV3Lrof4TOThVYoWvELGSjLAbf
g1uhcMMKQO+2l3khjnyOkchNTLp0EC0TvOZURRogBlLpBCFPGuISiGZybx5U
1nXjfLX2GJECkxVm4Gp0RC6OI5uZ/kW2hsI+cgVOMTqRMEQH83HidUzKfiVU
m97eF+QjVBfcB+63KzjprqLf+UuYUNTHMeplgeiE4IgqzemxDeDvg1NJIRA9
Iu1o3aho/GEYO3tw3LLwqn8ri2bmA7PhE7nvGI8mMEo/Tfk1hClQ9Ngwwjr5
1ovLZwCRA1LdhZrrVGr8JQgPfeNjGmznNbGH+pv0s7lVJFf6SCrfWNdlcR5q
M/pOplF5RGs89AjuCmzkecr19rKgdeW6ZWgcGLVBVySMktliBl9+2iPtP+ch
+NETzLylxgfwiRrE12jLggPdCykl8Fls4femcW2DVxZA90ze6uFgW0zu5SKo
o/1j2v73IZJLZQ1FoU/S0U3AJNiZLd11mf/LCs2Zf1IUx06lAH27Y8/apxp7
ZrKUUda1gXgZWV2V9dzFzr1hLofrk8f5uzCYuR+MK+DRJ/QgS3+/hsL2uCoW
2OqoYizfgyuScpFK5J02hmZQczEtMbpxh5DSSFmj7bmA1Zg4oR1DImvPOl5V
NuL7jcBmqWMWjoiptYllQZGk7TtRT45iD3AAYByhbjnI817Pq0mUYjAcNmf6
AhPvMY9Y6u8a16BCVyyx/CkoxfN7/S9t3mppd+lhqo6j1s+eeuPBhATlUTJN
bUhE8cz2KXrs3Oen4/RMq0ZInNeXQQILCgny6D31lLlvqRDreOcULUl8BenS
0eLh5IlA+hIkGlbz/GW1YHJme9pqHRL3jUCoJDAw3DNTKLE28JgJST7GEpCo
2124DQHXPRA8J1hAoNFIkG5SbNW0YTrnRRiUTtrb/lwVqSiwXOWorNQ/5cjf
N8eRLR6OEL63Q7zJE4lvEPxqr4NBtTI90OnwwpFavBFvKyZUYqIKCuVWzBGA
A3/SPE/EDijZPWDcz0bTwRYPCcDYdMC76XS0Txox+1EBPtg63TQb1QKssLPb
iSxfy0X19UME1s3qf1MkNBVEm4kHlihDPLL1MmbfFqilLnMXMvgodg0y/Z1o
x3LNE6jOepcMHhlMNrMu3pw87hCTVky8ftyHRR+GnwZjROH2P37z/5UqreOr
CA8sQNnK/DiyCi1FxANJ0RiD5X1+vkSTrhXgrOe/4zQDxTo5sMRjE3o/S5aB
1n8vT7OkaTglmWEye+pPB25JoOGmzBYYTBkV8SBkIUwmYw23fmevONVSCFmu
PH28ZBOmpZHBs2nz6SrQZ2PzgsCgvFyCyhYyjU9zavN+JW9PuJ56HpbwVAE5
4SIhTgm9RMK3NT8EqPECkSwQbj/ilTm43bK0s3M0QMIalu8qMEJRpEA4pflT
101ax9sz749An89UHlRnf0G1IExXbXU/QvF+vf5HQgA8HJdLxTHnlnt7yK3t
+PyUR1Yw4EpfvUhDgFlnIw9pdlIovlxcdrH6tNcq5cs1I1FcUcu0jJgZguB9
q04FyfeZb63wETSFfTSBwuZLwJ4ttP/bUJLRp9MPBMXFTpKq9yvabE4YXWX0
TkCnt1p0+CefGZ2D+p1+0nEW2CVRX8glwl08F2m3rAkDVjPJuJAXIeGdZpOn
vyV4x1p2lqfJYdH0r/BQxt7yw5FMjHyBxSvByYgZJ9BY2nhDQzLDb5Wi+hXW
kfdWy+5kFnm5cEwtpJZ0uR2msxWa17S4k19eT4DfEs1Z/cS5JWbTVm6bEugy
Ow9vS/tC0z0f1JMHi4OWERuOTX2+/cruDIJs8OW8U57pFuyvP52rh+ZRHcb6
3T32UMmm0NQHb27yzwh0T6NEepAxuTA44tFLM6ls0DaTtqIJ2z2hEOQg7C0j
oOBBUJvIir9r/vojlJOYVsPiCZVQ6/uR2IYci0fCpOI58RH3HqrTZJQZTLp6
A0BArAmIAftwamCIUHwWfydMYh7MaZwTLwTk69YgXf8cY/Kty2zdMlNcEllE
pUL69nJgAn/2e8dzght8+JmtkOHInlTgCB7rXESFjCmCXfkCXc2/x6d03HMb
MnPhSXp4alBq8YLbs9+UuQFsXO62QOXsn+3ZbjW7ULSmuRyGvmGU/OpMTmxN
TepRVUhS14PBIoVaROyMLdWu0Qvj4lCmBBv86xi5TDuQnbqjDwAGnR5N5GGG
+giVrkYYDrkziZtsjA7tVdN948Q39r94YsEzhUXkqoPW6ths3egVqp7xnufR
PttmNB/VqHKraMXig20sITkCkxt2vuDOBzuSAmoDwzR12vf19zd64LenopzG
nbf86LTtCAUPhxywAqadzze5h7CtwUD17KVKOF1XvxoBV4xByZ667aqkK55I
xjL6JE5D805o0zKcvXShdRG89Z7JlIzuwAdXvqhdS5O4807XaA1TPTVM4/2b
Z330ayrAscQc+DW5VfxEbQ4VJcfOyZ2smJW8fy6mi8kRVuFy8QMaRxgin3n8
ShqGi3Y4FDZJ2cwfqKU2zTb0PJdyLemQwvjr3WthRcf4MaoVTphVjjDD4Jag
df60SRKM2Iz90Aih62hJqf+qksCkMNNlE8HIOwzGQ9wNWx72q3GX6jl6/F9O
YpTEK2Fe5ZB7AqAVnqANVwDarOXKiQpihftb4c2ixnZLtLiZCb/GXvcIEQub
2iBXHMZxsvxuCp4UbpUN14/Op8xYVxGM+otG7DVT2QX+x6C50e/aI7ZLgMjk
4tlmXVqd0k91kGaOAWO9H8aKlaisFIU0AA+uNP24Fn8/w3NpB3WWnizpO7Z3
D39TnQF/H251CNB2q1Pw7sJesqg0JLZqvZQRZ3NCTCm0PaWjo35zXLpxd5gT
gC7NnaIuc0nds+hATy9nhWdzU7s4IUV7HGzJ/2tKqdDIiOwFvDi7786j9ckE
eRJjsaLHaPDw1oXGS3QDR/UqwtVJPDOrBLaHsu+fKh3eVanSQaspPxCE4HpN
bCky6+TzfIA/8BnyZkkVqtSOTJKTwV0ZKCZORT8BmkDPvaoY7sVptmh4mab4
t8DZEMk37ccyJe1XYbaQDU6oE79v3Yfp7XL7dsY1V9pHGdWfu6MLafqP6H4j
LKw4OeV+b5XEWXh7X7HXBqUY/HROqoiPmIoqOI2y5RtGZxsDs0rrUof+nIgW
ixC2UogXT6lnKxZ08IK3bWxiKYjiS8hYZI0TBszEi/4cuXeDjZqaDuJUmVJJ
6Bx2fCfATdcNYTLYVYJH4hmxbouYnN6rt+HRPXsWTyd/fufZtMiUhUz4jl/z
yXU4a0Dni6rdJIXmxZKIzpL5zTLgHqoXRd45kHm1aiZS/y9rX2S0hLZkGdBU
DO6yFKlt6gkqbAjcvBcoW5yN2mLmfHrUmxejcUe7KZRx8h3BM5rlcpp0JUhL
iC5iEukMMFC7RCt/ex/WFD7mhTVRQv4uuCX667GBpR4BKzf+cYQJRt6/WK1K
fin/h5m663qm77ZQn+Qv4R1PWLZ+MS7pzPyQz+zErFWfaCxr1n+QV0ElPv/4
ZjCwCfGvuwAHEH8YB4w1VJY1KBh7KlyAG/kdPmCjnxCs7p40eHvhv+4p0hOa
KmBAaw27RfleMyRbVzlQgJofXbVJ89+WQjVtSPtvHbqjgBStttVWZuNOqMG7
k90AibleuOU/Buzpmyaot177Vc1kc3Rkf3f6i1QajjOKIyzgYVVRbVL+uQwl
B5NXIAy5ovylZzmZmf4F0SKYF+sGui72Nfin9+o1Iu1MvXN5kQie8gfYQly/
t6ZKQBMJM9R3TjYUfOH6n+mREQPfW1pvlERbZxsmHeoRuje6p/WoMEFSxUAR
TmquQs51U4OMROA2CLe9UnDSi9ZB1WjWOtPtQCLvmTSd7caEna66SQ1R0vll
egDd9gbKHUt7t4boIIW5I3Q2L3cXlcEtpvZ9AxEJKExHLaTR69+t0+6jL3pA
oBVvpSMoRYm8ItMaEGlWSzMNMJ/0zPHft7yKgd5Yj9xbgMxvXxiU+7HDV7Ev
hxpP1YipQgk8Oc8PRv+uF0mKN6pZblt5jbzzq1hPim11bHAPa1GhZ/fF7tlY
UIm+SMsEG/febq0qB/3lerfsopDV3J95/dkazIg6zNRaYnSi6SfxnLauuCuh
RZoLiK8ay8d57hauDYhRvtn9vmFb3Y43i2nrJOJ1NRGoGwe++oAD4onw4Spq
oeHIwTkC3o58gGk4u5h1ecdI1SubglmRv8UTKnyBVTyueS3LZ9OZPEZsjvJ/
P16buv5LT7zZDhze+gKJHpDF8sYFFTyxyjASVOQNY//CDFw9LRIKMh2tSwV4
m+aRzLyLSaKTaJHR4ZJtwECoT6CcHZbzNXKhUUGRIe8BJOu9/4xuAfo4+yrm
UTt+pnxpcnYi0swFmAFwdqYC91Jkb5yUXwmE6uJu0JZn7g5hqcSs9uQ2DUd5
BdRn1LOnLjTWae2oAaBv6awU3Rsu8L0N7HZKqXCjRCdNwUhfGn2xeDeOoarn
KYIxbsQ7ckLpwXlHKEv7j9wHAe/0bu0ToMIPLMs4As8+zwfvvcRill9xzN2t
J41uuNyu0wv/QI4WHOGLOfGKS1a7b/1Sp05r55HKTLLCKjKX3UdOyLGVtAKz
ykVjwcMufcq5xgwKC6P8Y94zlIFJk2P7hlzbctEco3n7QSf1O5Q3SgU1q6Du
8KIux6MM49+5CA/Ofz9WhISUi0XpaGOA8lLRt085TbZC3XqPLltt4rNjbL/y
XAfGeR60mVvdeRE0OEW3kujzfjSDLBO/kr+VAgde4ldBjTMDIMixDX9l2jXX
bzWh9fFL9mvLYGWJV3cCY0no+TCyS8q7sdHZ2XkaEEsOId8fY8C8gQsh+p5i
3zK87gVoSIbjEURGLg7GiLh1unArepEvkVTpJxAR2GZmba3bM1OWYweGClpt
UW5NQlXn00UqhVPTHFnVD0WbjAtke50UFmjjXQxajsyVxhjnFqDbAE/vsnod
Z/btS4yrMNzxj/ppDbhBXbOwaNIJoL5yg78gQhMNMAy+AylhhuBRNErYovB/
Eo53Y07uGMQ7/sUP+0zqDpnKNiSR9JVbphrFT4j8L8ZJ7sUfQLurJtNJ5jZn
OlKmSoAMp7pZ2APu7BJArOnHu6nNvgSOo44RCmYRrMuHSkgJix5+s0lC5Mml
jxWffsVHUX77v/JJtCWzN8JHIYF+qe4f4j75jcz43a/RAJPUtdU7xpeZ2r27
Sm2xB+Uy6S7dfVOKIZTfYedhkK4sz7S1W0DLFrKkmYceU29AmRn34jBbBW+g
9YmZFBI+t6H4d3g2MU8A1FnnW7NPWdfnSev58u7zfPB3q9Fx3FKAAFVxbF+b
daWuPGHu7OyFla4O148HHJ/WYhrE7ILFR9v6HoZBhwr2nJNMp01g4VYJFDcY
ZVQZMqAnqn/l8HCYc+1RKT0Z7e5JhNbcepIasZJVXEg689zSk5mlmoVg99Ve
uRAd83/SADKiSDUZcp8aDYcPwfRCc7ccUMwdN6nhn6hPGloY/M8781LKEjBN
KpAW+YaWRmqAqZjvSj/dvQGGoGAyHA4NONqe4q3niMHGg7HjcbgW1+YIIJc6
T9wGf+T1iw5YNHXnNmlh8AjtmaJ2ddpyKlvBId7led/+6425IjRchvvtVg1C
oH7e2ZsScxcTewOLiTWqYbZKHZ8AfHUL9+8SL+5T8OtlqAXnjzB2lYqtnJjw
tI9Y0QrRTidAveYolIwWu1Q1eyJRQtOYR0qP7ajQcAe8NcUCNsetVFZ7lplD
q5Y0kvPxYXlm1n8Jj65xzqZQOyKrHJr45ODV/55IBE++k1BQ/Aq39U2aSvQJ
2XgE6wzay3/XWwFSpyM5unoGYB3FaG2zO+lUtQcQ11FK8uBQ74G4Nei16cQh
SWTeX1Z5mWfHgSDM+6RAtt04rRmP8nrGnF0A+feprj2toAS79LxmIWsJpet0
CPp3jxF1BzdajXPKV6uucs6QVCjRXeE1/8/TGJ0sqk3KqjOM5G78ZS3QAoMt
suTrkg+1z0cF1piQQss3C1/Q73WE4xb1sEfcbLivq+HnqwbgnCZ2IunOrIsK
l7JECvXfFf5EKLzNX0Pd5jB9hi1LB0nJ1EwYWsiDpycJdpgtRIck5WEqehjD
tgQ3kEbTHYs1ydpHEktjziYXQWHNOYnqi71OrOJPv1ZGhkjDvz619XQbYr/J
jJZjkxRcRcM20CqvMTjUF61+lbQBcpDEKGZ6YHUEsRAMeAwGtaXtd9Q2oCOP
nYb54UjZuI30rPh4kwdURsiqxbenAkoJ6bMy64/pHx5ow40GoovUg9yoGxqW
loAhBilS0XTkS1GiX2DG9u+zWHXINBivjuTNePQNGk7ULSzo+4paZovIATje
paYHultQ1T/fiqImOIFj0aBuViDUfN2vQTt3LZuEuZc+8Otv6UG0fhUVEQJz
8TCiTZcDoG5T5TFNMXph4fXXyu3HLEjhV018fAzclx9jiH2H+0va05gJ/Yfp
RB0YRL2sQQmW6pZR/mJX5u8WabPlU/y9Ki4C7WNdUgQT3t2Z1Vdb94KB8T7m
vt6clDUgN1mv/B/H1WIKXmecmcTuFl4/OSXh1l9Gg4rh/ezdVN2wS7+T4yeg
TaxL/1WfL7hqZ5iHzhQuK/Km2aygm8MFonmh9ZKbgF6Bpt7KO4cMk0/T/y7C
0Cwa89maXnEpbuyNylyULUJZ2sCl3dZt41Tp2aK0HURwrXWHh5DvRpIwQkR6
LZT2D6LpKBicjq6cy20Bonc9r1xie8kgeViw95/v4LEaKwyk/13D7OAAT/IL
SuI/KE3CoCTjXGMhba+/lS3zQ/wdO/rY4tngwA2VMBRoWq8S1rRRoJy3C1yM
XhdoPDCmhortqkgkyyy71tombpYXqSwMNzetMfsjEQBf9dF+qKSwJyHpydov
OL2eJQxlpODWqdr+uPqb5IlXokv5n4b2FIGRXgfl4K5f9WOmGVrQhMYbMSly
TRxlnWAcJ3RkNhO+czy0CwlfAbA7ag70LCMw3A12l3kVkfasZSu23bOyqHk5
a+jpRtbLZrhqfhkvyUzWZRecWoFpEAoM8HNmI6QbVXJl3huaC9GKHBP+9wKA
Uau07vOjPg+hsn5c1klpDhZ7wlfSmXPg9ThsRsVBQZ8A3GdX2u2Ccd0EXISm
Hn/gYO0I1T+qzHcxHxHDpsYyUT41KMLnGsrnx2Y5/ordcgyhHfI7CLGw/A/7
MrB2TtPjiS5b/a4PsGQXHd3ENmChzd47aRH1OT87XGm0xym8V3FUkI9Oi8G+
bW3Vt9Y3tPj3GJ0rmujEiq5BLxHFUFEC5ZiyYooAmQEK74ppvpXa9N6jveZP
nbKvhQmdei8cZPBrWeyOfJWLx77cNptBqMToIyvtANsKrUa4dQ92BNNUMd8v
QxyNeU+ex/LCd6nMjCM8nUMUqUuRxtL6ysSHifbER28YWn2PHZ6zaaaqn+6c
48+WOludT4iZPqSsHYEtbvJqx60X+Z8/E3Pe1HkewSAaar7GryIyeMRYaz78
wYhdSlnoFI7w4ddZPQcszhnZ8xnB7iHYN5oaOFPOFLApXOTdhoFhJmDMfTZn
0OA8WZ2FwjL8BrZ45bUotlZnvegi1csyqruz+iDaWJMeU2Xpb5JWRbenSpsS
vOht+5rGndm6qBPSAzY8KWKU2/c1I9QZuZ5vS80cYBz67SaSleymjiS+sUVl
i9gOoqUgmtGPjYkKbZTTbPo5kZNcB3Oe5S6rl3aFholcb5FsfMLQ8gtuXE7M
gTppa4jemYBqWVw1lY18F81wlXBikpYNGDrLQcUCLypxILtt2fZPm+OmdoyC
NItaXNBLLI8tuFBFn3Hxe8c037sdpQ+2mXH5vI4AQ4QuBA5dJMBphzWHVEsd
qi8kPEMLQLhbsUmfTUvRCLVMZ0JPiqiXe9kciYxuvY8Zhqb4VQuNUdCCAac6
KhaQw2XrzLOmMG2dO4wYtYC8mFWAKWNAuARdjXwjrNWsiQdvk7T4U+jdrj3M
QLETa3dE0D7+KNR6Jgmel2lojuugNWkBuLQQdiboE7D4RC6itaP7rE0mfWUg
mrFWi4KJWWHdF56Fdyt7S9NPTNaql//NBKLIC1Bc1bOP7HJUJEiezehQ9QZ4
OHL+3+lpwzd2cPuseYrrx/dttIJ8C3wlBxx7eyJn1qLqcDSr04AgZkR1G4Vs
E9qd2aeYrHIxzFCb5OSMmu++zkZ7a/qESAxTnWAwkM4hYk24IH9rtorD5mk4
CmWU6HwqR49oK/20VOKW/StrBqvB0UJGFc62MmyIab5PMEDxUqtKYl7CtGUU
gHb5InMrIwEAyKFxc89X0W5DMCxunA4FK+MWOAKEhKDgmO3do82Tmav2lG6i
1q17jzNwFr+MUhFwabGCUPvvizDYXkltdQW1w2+Y7rpYFH+B+b6lppidXhZ0
kt6KYgB0HN2JcDZpPXRmSlNV9AS0tQ7WBjW3dU6HsWXmkpTiEzio209dasz7
yW51jW5cZSnOKgIPYkk7dAO11zRgHa1A8hWND+aXVU0cG7z8f+EK8oDW8LQp
zLUAOH/cG8P7brxIeub5r8nVXuAH8St1OwTIKgGSDsf2vJ1qezMkDyKIeIyV
7ozu9p07/0LuJHDzlZl2b1IHalQ3wPq88WibhyqACUiYbJWCkvPylpAxnN9c
5MCASEcl1cJJ8yJzbS3954TfKEOr8zFUfjor6Ey0s7F20F9hH02JduR9XFeA
IA3tNdEJZxSnM3/KDKE5J9j6bX0SzMddExTPAOYMATXQPrQolHg1b2tYjk95
uXZ5/aFpac/SNHmVRhOYp3nV3UJKU3IlT43vJuh2XZKWGk6U7796cxWqg7kH
nQ5RO2T/Jbhp0XKwt2rr0VNlQ5bh9B3z5SuY0TnuWqr0+cSGmGx/BtJJD9bo
XHq3i/D0e1H7SnKdpziUhRfgm0xQgAZ3pZEXweFAKclqkvzqJu6MRDj30CR6
elcHrh5TXvJRpBgku97aJR3pz9voxCgCmxF1z/Xv5iBRcH5OEzkzFj0X6Smf
H8sDm+4VALdmYJvDr9RL7nAs1TqzY8XX1/0dMHSnlR2iXs78jfb5SNn3HUk9
bBONfZckGwJE+IJ4iWxjKgnBTx6L0Tr4QDhJqa8xkUKS3N0ep4Biggw0hsTo
d5ILIctBxK07JASXrJrByVCuiT+OVbAWJlW/ozCZy0hvYRECalIbLWxFac23
9rF5ywVULls0eKJ1hIPILrzzGA2esjAVYiEnuqP/MyNVbzWtUQYwS+APWWBm
E9ZlnscMcAOE491DeFqwEeBW5jJDe6sp4gJg5C1qnyr3U0u9jsnplWTLZUu1
LTC+GqIA6p3IwT0RCUw20Cv+EjE3rN5AgttLGOTd/65o43aAIpDgnK1aJW2F
fLLaeAbulwrWvHTyKtfv5NJaGGzX9a7JnG+5SYkDcd1GWV7ZSVlgwqFUUfwJ
g+HnwFTD10523YM/6jhsEyyOWerWS++wNvbgF+qWMX39joI1xTDu7OPeiqqS
inr480dUnYd3ZiGNtE2g/O3OTJgEq8d82JA9kgvYDWNzLL0yPIRZjWeZDXXr
b1L2H/pvdGawQp9zva8W92nxIYXCsXM7/BdZEAqUt7a9FPm9CE2fbWJZxbgP
GpNkKtc2Iv6WCV8Pip5+ZTn7V64O8tnchcp0PNt/kYRyaNVEku3F0odjfLf+
9NUKfXZSvS6XTnBeftqKX+tnue+cc4z54/QegmQjjerAw0/ihx2CrydO3+TY
cixNjbj0ef5Z7cCrgwLKTOREkktcGiI+6zpuCzwk/7BOjtr93oTy5/kM6dVe
7bnIPdABLFQ39roqGiErthUYT4D/LFT30Vb56ekfGxU6CSpQ0JZuftZmTqwl
qhyVmeNNUreSnZJbaIgX3cW/OmNFl6kdz2Yb7RC5U0d+oou0+L9Yjip0qGVy
Isr4QzyT9kF7o/F0eOi/kJZZZGR/tsAKwtgc6zj47pedJhdU05mbIvsb7WIn
pp20a+kCTeYb673dVNp5WsJjYbBShCngZWh7sf5wemuxg7G5rfx84yiRm8W7
/eaTwBW3vc+r9AsmocIEbiWpKlqLx1yIu7adWzy0/5idfrw1z+Qa3SRXlit/
EbDmmc0Ke3XEvDP88ESmOosvACN83XRzZByfctHqKNs+CxYPH6gJTI8oMiUO
MBxDOWAKkSvMyRbZTY/Uk4kxHCsBzvxZah/yOccvwP1G9Hods1Fupt+M8AgY
6AWMXI1r6SnhwSIfk9jMkM1TSQuAZN54aSXGIGR2AMeGAIss8VcHCC3MTP3i
a00X2UvIpQ3oinLehL7RsFV0GxQz/2XClQii/pyvREuAOZQb4bMSGIF+Liqc
hZjW0mF37Q3GY994TfT55NlW4JPIQQbJV/YNYVXbWHQLoqdS+8hSOOxXEG4C
IKiOhuCq8lgz3IwZ6ombKcg6XNPadnDXTU/om8ECyPiAuf2k84qjzpVKkF01
MqFfQzQ/bG3aELs3xOAseP0vBDkYtZx3skrlF7BMlZYVwNoD5ATMvTC8Uc0/
9ujfFxlb9y1nW6jxdVTw92yNij3yc4ivCzRHPSHHP7/NG3aatAtRVpRrJg9J
EX0WLzB3NRfp9aU57eEiQ5cauQzU6w7h6sbW1Y8TfXzSem2wn/aZseiE6u71
CcXgap74+cMWxmkAv1PM8COed8vg3TO1NmKMB2Wr2exK0e0mIEA5l6/duwtr
UbZPhZaFzF+Re9DOBnTJdlS47IviEvrGkarmtXGDsus6mDGJnnprAVnAJJsu
RlBCXUsatW9/BHPraYenmxw1y0QvXgxZ3/NaP0H/Jvojm0r7VJba3Hwdkmta
eml4pKzn5SAl4B0gUlCM5vWFUSEF6WiDYfE0GI1eSfFntbKEVWc6F9ukYRFo
Na3p2BTgzI4by0/9Cpjz+qHb7LlZwzNAe2r/vMuGQVt11LjB5C2Zf8AI/ryT
DGc7jJ9isrcRtua4xxpLDW0JbpOQMZ2tP4hv9ZQhWJbBFfwCVfPCUHTvL69v
vXFzO1K5pgV6IREbIB+Dn7OI7ioZ+GZlip6vnHV+6Nc2FQ4BSyEU5cT7+Xx6
Lg1o02yBJlEsPZBNWiaWzGAZ6qAdrMpYIfXRg3pjb9aEEiqsH0oS5fkWjMnm
hgQuhSM0vJMBnNQhrfDygWcPOoZHgsFZhrAfLsNu9AU35i7Aa6F+X+LVxutw
F6WOy/cEUZNBJ9FUffZsWozAt4lBFTky2zRmwfBWR6CQmpcZeG/zoFwA3Iqr
8Etzq98cqpgAK9ut2cilCtVZlYM7l5/3jlCNKslvzsGoocZPyLKCz0DwU6Hn
7Ffd1VT2P3clEFVNtLs6qd29fqisjeMNmkB0gMzzEXrQftqoMymZpzau1vMt
GiHFruf/C5Vi407/FNT5KpNAKKd09EHZE+PpXd7L/qSjvhZNeTaH73yAw0sQ
v0X4Y66oc4jq2NsVkJ7ODc8m1wJ0ztv4D/T+6yYOgWhvQb4hgiQQ4Qr6kzrp
ruJS89A4vWMWkJxNfgPQh9evPLlppTRBiAalLxUz5UikU2j4v79kJxA+Rs+N
FdCDV2Sm/i9mmkHolyEPROZ+ICOk5OKnSpxteiCHjRoCSn9+CI+qFkIN6nxm
2hefzHkcTKWxTZ8EaPphHUypNP++n0Xti1QgEnizw6ILyFoyawDUmDBBMc2E
j8L82wvn90QPzNlJy+T7xjGRzzl9fcSGrScm5kRg/n9/DYuBzrBRLOTMt2Cb
CjYQN110PWI/uuFOpejXW/hSrsU3uKwX2XZA6vAxssaCWRTCOVpsx/KBqg3M
4a0cX2nv53OOLoqx5kstH1WGFXVDU3iSLwhqOOKRveLQEjVppSa36Z7SOjbt
LC3Osholb2jq5UzRU4GaOdVQT5Cni9rbt8iSadkwnDgT2ntr1lyK+4zIeBGf
TVc3N/ZUF5uukCuB6f4bhajRepu23Fq/UO0NMJ4vGHN70m43/9vHCvKHxh6X
g1NL/Iwee4JAX5Et+LC6OlT5f8PZNXs28+7QQIbKTprHWJ6OMFBx2h9ipP6L
J0r2x9S9/ONz1B9YZY3zIydhDbIHDvf8NVloS4myM8TocjP5HESxmWRUsOA7
Ne8qH3EngvqYW6E9qCPs0S/X0v0drTUiyaURI0JfGne0K5SbQXRnG/TmExLi
GLVlGrX+vmCjg0buWdfwkKRTLA/yOscdbEszmH1RFrt6xCeTG2tO8dkeuNbx
vP0jpcZ3B4zYdIwdGCSdXVQ8b7g1mM8EDx5xmkPeY2UZxDWy+wvF4fanxoot
kPGdtsdswtY+rOKy4Db1NGzmLuvGpiuVKl2TVlWATufjJjFpsYn1YP9WA75n
ZbzlmpF1J7MeuEW50InqxkEKtBI7FJ6KezYlXsoUXVQ3AsUy59wpYIOao/9q
Wnu8D8nPN7NwN31TLTb5YZahelJh7Sk8BPXkqcqkzZQJ7cJvCHBL2gfZnkdX
QozbwEc6YM/Wv9f7HJKgjmupDyotQKUai+cmy9AdFSdW/xMYT24lMSBG+MY5
+ZkEhITGsS3PO9ZUMPhd75piJblfOXHaAnceOB4o/pjjpq1dhE5unbB1Y7bp
BD2NHTeLvQVYEP3toIEbODuEwik4ScC5Q7RlDA4mkS5Z6mX85/t1YL27/xBm
VZ0rmNth42SY/1u/2wPKzh74KuITkj0WEV0GP+V4iaHEm0Q6AFfX1grOdyyV
etqkH+s+tz8EqcTMGMyKI1sp6H3CLZ51bbhgw1SOwc5++FYGCfCBm+wsHsdy
V2NiK8dPq3vBOz/xJVvRyUFoCfjUQ65bxFKrFEwnzkb3ouVAWqtPby+JyjIO
jS4q+NXA8hlTWudIB/X/FJdTus1BFQJnBboIhCNsz3fA3rPwmrqC3OV4C8pc
u7V1saMVRBppRhwLDYPUm1L/nY9qpPcNgNMpcTaw0ub/E5Z7O756LL+DZtuH
AsZW62Zk8hyHVdYRJ9J6uaD+fAaCQe89Tg/z9F7y4riLF+vAWvebO4B5xKJn
UFvABOn3AsKZAsLbwgmeMZpJMKf3+kRvpgTJsQ4fF+PWWkGAH69mj41Koq+u
JwQZih+aje4KhjHKSUKceCSE7wDEBQhZfnA5+v+q2poLvTIS9T+mAOHNwFIF
o2e78KfTNPsodOlqYVbheaOGMcHbUZdS41nQ1vs/qjeXBUJVvr5UUqpAriaP
0RKI9GN3PkiyNh62Sh9Tfi2iDDlMEIvChTppmEw55+FObqqTDEdKsERRvgka
S6Y6WOqsxcLse1XABvdEnF60v9B3GckZYHYV4cj08NHU22sM5zDKaFmAYLU5
LyY1/Fv9EuxZUiON+l+hXxSggbPVq2XC95U7M/VmIHMl4PqW/GcHVHWewplQ
KbdDdNETuiHKSouOI6Rydz6Jtb51KP68bZjxi9PshBqGaylP4nS2yEl04QRz
xrbmNAw75Lcrco0Pw/ZIUkhvXIxI1Bfj9tmGP13xrlUs8Ij50lIE5p+NSdTS
EwafsPAnJwksCuKdFVdgLqC08OE4PqOURqwH3XUPpafzaXSfn4Hr55duvWRq
p8FFp1gsC6pJyiAuNR1oMiZNWQgPS+jRQ5JG0gbPchXYI7sjDTzIwA94qe7u
saFMmZwPPufF3Rn3czyv+LfB0L+bk18BFA8myRHCdGgEEkM45mGCDESbZGOp
VszhUoCxiLylI0O4JB/BveOwcpolIsAbJKbWX6BzCTp1gzQQh0evJCGORN0P
XOnWLNgCnSN7DciMOfE9rf2m+h/ffxqJVQ//PdV1eqEIcyCP+jYPMnLxiddn
DbhqlUcxzdSv84LIOxCO049gUkgZOyjKzICFNHPQZLEla2EYuL3CBSFhZ+yO
F3DntEx/DO1IPf+QLIdBGWVE3X/7XXCFJuPrn9wxgm1nI35EcSb0zR2R6ttN
AuGq1TGrxSlCd4HKkOcdw/JFPePX6DILp8kCwqow/FbZybOMN5GnG69nDZw1
2DN6FFhDkUmWUkVd4nAm0NaxFs+Y9lEFDRPkQcid133EWsVR9XYniQvuRNV6
UU0zN+rKTSCzt4ctlGHYAh88sD5SOKjf/tYlAVQChWvQ3fx0XeQx+8KGBiVF
2pDxEA/TJFO9wKvm1kGNmH/ecqVgz8a9e26X1xW3ZJFRWzH8Ua4OHk4Ghk2v
FTxoudk2WX2DwdvwQfLFiHyoCNljEFnepeE7jPonaVjxIsGWQkP2b/YWoZju
t3KWLqlf0QXP9EgmCzsmIl/4HyMjdf798sc/Q88osSYZ9QLBaUOGnxVNwUNn
nGnMBdYNjl0juX5Fu/GsxiUaIPKRbQ2OYt1Mv9ll5LF9nzUWanic7vSEfU2Z
1qTJaNv9Ho8na+Sr8NdzLk1f+SnWuQxtGqC2ZEOtbPqHwOfX31t7o7xjuFJT
+zRMV/EN4S73udqCfjYVEcVgl4fC5qqKkKYXsKMG/wDfXpkde0Ige0JThvbb
Cy3ON2CESHhPWi4KJyDIeXvH2QlZ+Z6ykpFCjQnEWqUUnSBb7dRusQjEXF1e
Pwwvgfz0kRHUyry9xeGAlXmdUL9CsQqv0jBm4nzqxRD+dQzcOitv49H3bHpG
KM89KWX5YnWKZqhWY5nHMHOe5xQTyMNHaok8KMJ5BUcjcWqRShCzm+8l37AC
HjBONiZw1knBHnnCrr4z04giQyRH2AaUmuT+E9dx6O+ki6g+sjmZT8omS0EU
1cCQuBeba8uRJhHqFPHyplhXvjj5uFvuFXW24m9GSsrFp1V7/qi5B+xRzEva
0XdysEdb0IHpW4Xdq/WkUTkJud92dtBETqzgUwew05vKKdvhws6PLoeEi6dH
Wsw7jTJAvyKKpZpc2MYYFMv2brKLbRpfDuE90xm5evucTZMNLRcJ65UrnQ8O
ZZcEiUNvd/cpvE8egy7+C9oyMAoc3vpWqZGuu7ay7VVpRc5VLzCI+iTUlk/k
OWeitE2iJW8bhsUVN7Q1C0KxrlQJ3ZwfB4p5cjzFeNvvc99X7IlksKiijJU+
MKoF50lf0YrkRyAMNlTWmwJVr704YOebqVIWOevw5L+vaNgZ1aq6sNJLyzf2
0uZ2U63R6rtqQ+8a/sPfj8lemlBxl2dHU8RbYj0gE5ytEJS7+Hkh20LeXQCh
N0a+ewiPSQqrvjTfev606v7aB4u1/dymr8S1Dim4ZRQZVjYDNRL1SXqhxeXH
V4Yk2e9kwWuOQT6yytUTCv8wPxGVlFZsY8zTU154SN6nebdfzGIGCCT6/SRG
bNUPLaWh9/8r24gOeY51vP3MfSHbAEQRk0LovGUWDo9wc/hseWCT99nUn17r
WW9IpC2qSCBGbaWFibjdGtIl7xmiSx4yN8ulqSEX7DdrB5UOSZs6qFwY91Tv
BP8vI10nyuJoZyw1jjwFnvRjVPJ28Bx+FvD9ioJg9kwrlV0ONBljKUY2bJzD
0RuzKYwNrjBT2kj9oyWPsX6tBNyWq5vt3Xdf40veuH0c8lDI1kW42hf4U+PJ
qY5RkGInSlps5zZQ00ol98rIFh8jZDYOyGNjwPtPnByjeq4QTVQTeEIBPaYG
eQxjBHAAfZ3ZCqwFhjuyVVf1fCybPDoZP2jeFOax7r+CWt4a/Ivr9HG/V8mX
CTs7A6dpQdASVUxd0c409LqHlPuCOtRtUZmeC6FhoYIMAP5V1/giVWN2nR6d
DUZrALJxMkjVe58Rya0BcCk0VrGk3M9V9UhfVSEl3w5XNcsM3k4FyhHpNnID
Zh9yGnM3V6R1cGXsJS8ZiYP06AdJVZwfzKcZvv8RHZVylUkVkVo67p/6mWjA
/qasczwklkzW0ApNcignPY37Uwp68X4OL+Tu67hAAPot7WemG30Eyw6WnGYQ
bAcTuROgZlP5DOyk0EQ4mSAlmr2AbUtIoZK79dWfxHP9xsCk8NjAJ9yR84bN
Tr5+KU+MtJdIUnn+29qOMP2IGSJIR/OLQQCbb1cJiC2lD6L+z/pyeGybOy/V
MNaKquh+mJjpcE2jse6LZHBRzqqwX9wdznYv+/TGbtV1tY+JqtQ1Bk0/NcX1
Wl5GWiWTxsxEtNqZYlr5VE9Qs441rsJjymFxGMvzZlaHoExu2c9VffefpRgc
o9e3iCog5iw1Re/1uicZg2YqSu0IJFCeZPpXdCw357N7rvArchUEUISYdB5m
vNPfrR12DdkYmacYd2wmI1sSm8njbS58YYD7WT2/CZySUFju917kucM1rUQw
jCCi0Zt6Lp1C4HM5C+uCBcw8BFVMuNYo0w6UDY0NW4oVQaIaZL0bidpxzlKH
3MTFwvTLzr61JwIr1/xn7b7YE6nQVjequUmsvnbsND70nPyEhJcQMCByUH7I
nv9nGeZRtczsnAtkR2lf3WqM0Uuc5FXRTqR4eLvnuRfCw9kEUXYNxJE8LFDV
OX+q66jfw/erT5IdUibQghZIrmYZqA28ZINSMNA6uya2ZsA1kVvqm7XudbNi
esbMIRTxt18FS76s9p+za2Iodl8QJtxsgavDC5hBPRGblCM5ukh5TEvkl2+C
a3aZHcYiN5LLxNE9cSgKYAnhRa2sNFCmJQz9Q90kN0zLXtFl8VrS0dTlgrap
UP0bA1SDWxCt2IpXklsI7GSB0NaO8BABSWcIgbNZtRvRlSuahCC4PlAhm3dB
EQCIAIPo+UYDWUfqkRf4rTo54dBuI/xkx1N0q8a624B3hFm/HcTWU3hPNZx1
kUZUiUKgX/WNsLTGSYukE5qToQHqruUs3u5xgA64FVBhzjEllkDtPOSD2Ga8
mVIOI+5xpzdHr4Wu+Oylylx8+ds8sDj6yy2wiU+bQaRAfUFuizkhjw5bQjL6
RCfvv5+xokjx0nJEpyP9mcUqB9ZQw21za+68nbAqT8Nl4D93DGFoykUWNbnv
z6f7QlARVRJHCW/NmuBEX0XnY7wUA/RIGEsvc6dLI9W7rINSgFyGPxlk2iUt
fJ4LBNIeCn1OD4ZVCB1d7KzAHu/NmgBPTxtxuxUW2wIhKR7FxJpDLYzH7QOl
OcMLVyqw/r+9DAgLIvMZlTCO8MwBRm5euXStScIoytBcu+Rs4WwEx/fxukMF
v6kvBG2Kg+HUBYtW/L9qi1Xret7tzNBwzTmc1NXhQiDKDIC0Wyv1sIZHG55u
i48OIMqTE1Pgg2xhQ5azgpddvlJ6rYlU80MXI5UBtiuf97DACmNh1PvF1vJu
jjD3EyLiJCzs8U/4It3bfM/xGlrRoIo9bj5Q19l0XKLV9Tdc9wiSLSL6ZQWe
GhylgQ2CsCvdyzSJq4DIThTtPGwF/nq2MnKnNEaeBzka3DYuOfphPMbunVeK
djPRFCPQQG6zf87CKn+x4ye44z63mT683WkcUIqefHzX2KtkDNkSn5p33+6N
1uqchZQVvkOcYWQpRReDXnF5v8z+2TDh+l0WPtCeIc1sA0ab8aRQJgcmCeyP
d76MdS82hVQrLiZyfIrK1ZlSaypcpbQtA/+jG5p/XcYaRvW46i9yVW7LsPcb
UrZGZYyhjrbS1kt3cF7+8ZXBe1RijdEJIRO+WPo7zUl/9mZUlC6ukX2DEzY7
LRE15hqFrq/aZAGhKf735BYG8ME++cqkHbHkvKCNzzxOhU1+kLyCEqZvuDrw
3NmVUJxSyIdvemJNZAQD3qbAbke+mXYw7x5GB3QAyxBo1O+NMxb1goikYL/k
f9FJlL9nPRVWqkeQkFvCA38hQpqxd3hOviYviONaJM9m9DsWah5JmKpvH5S8
a8PIo3u1Lqu+18U7MT3WKxgJDBcJQdmj/vm7iTVg7UXY7xqavgqKc0rZSyyz
ZzbZ2oZA2F1T1KnxJmj9uYJT/o4A/84VaZLOtA92usCAkMS41xuZrKf+4guN
sJxpfTKMHOS+9cH1233C/kacjPEAqkfKgiSQVPYsmaTGWaGnsDk3q8Hehv5i
JOnVWM7+MtrdHwN/mEOnpi9XWTMfmyzEt+tJDi+KNNi6nq+DuP4m1AWORFev
gpq8iI73AhB9eShlv4LjnenZjFUyhkYL1kNf+/BHG9qKFiHEo9fFuPGrM58W
U8JqCOIGEPFjvwRYJzgEoAPS6J4e5XXhdMyBZK9WdHJZMBUwaIPxDsI9vxR3
imTgBVjulDi63cp8I8ScW6qiypjjcdf/iON7mWfsM8IxDh7Z19hntHi3KgUb
uuP6oFTgTpeQ+3aGLL59Xt2kIzQdEMKB4kwHySe+yC+tqNXmzq1GbOuw7ynJ
dqqHdhTyDwSqgqXaJSk0vesUz5QzlRy899qBKTPsAzbrKv63HuXQxXE44YRb
g4z9KmRdkABYD5a6/xhOEnZ0+JpBFaDWFSUH7pgKWAWNqffxeq91NXfCt44f
QHzIw+27P9vLhIp8FRaeefc75RgQYLegWfCUCRfmIhCfnYRmnOsV3uzRXV/6
FC9Ux2k8QzCGNsblewAqOcBoEb2RZUO/t1DOA/9ZhMFG6dD3wvztmHAvppYn
wknsCnlauJa+AgM/3UCbeUJxFLLsyhxB0ZzYUGYH15Aq7ZDbSIG2cGVkHxXu
KGSMorE98R/W/8dbnTITQVvwdMVYqg4j0fu2Cf+0TEXvqGjruDQ7p05VSD73
u/4lYYWpz5kmV9e2t+PSl4/RKTOC8mU8+jyVkc9pbc41fXjJpm9op+lmLi49
l8Gl8FHU95gOn02JVlTB5Cc1LmNs9f46QP9tndtpysuFY8mMw1NIEnDIdwKv
QM7774qYSPuFrT5X9LtBdKwu+dlajEt0NyTFA45Sm0vkcxIFSoVEPUPogpEJ
/SfjDmxyTeGF4OaWDSGc0bl6Z7fyr27yFGdmAhauzZKS8iCeS5wGDaQsGDwj
3v636gElMH3Ofe0iVpOOdsIl5/crAerejqz5gSqDjqN3IINIf79QeCjzRWhz
DSRNQLePnftQh2DjYrIAbtyZjQv6BtkhkU0JS4r2/5lOoMY4Y12SW+UMn/Xt
Kg8Vzgl1xfjeDd3HyGxhwR7SMmm8Xdv7GLuQd/EXCRIuYCjqshMC/JIZbJkH
gSUWlucvNDx5U8+t21oljswttyHWm8DmcwlGVptH0JzC1cMddmUSa6EZB1oM
lrS24Jc62la5DM+F7BchRDRrZQGGMk0tVlInKqZs/775Ppc3Axw9EE8v84Oe
yEi2zEYkeUqIUhUAYXD6q/HBFCbWatWFBscUVBFFntmJVtkimQgpnzWCrGER
XVVknvBbRhP9bvvbj5kCzZDQlNe0LvntbK7Woyn6tIERQi3F9QyB2nUc19P5
a7vNGMt9QzbgB79j+VDkvmO67JA1BU1xovu8tAYaq77MZh1K7jKQc8NeOj5N
FMldjw8J+tNoj5EER7enRzX06kjVmi/Xmi1OR57DA3uCTbnpygcqaNp9V783
WDuV41IeiPFklYP0U7TCOuC7IvlFU8ArX5WRN8Hwj58V+5B3Ohss5KgAiDuZ
c+UwUlopAlFI2VftX667lke6kw97brjrub6lwpzKBkD7L++M9KGZe9uPKN9F
jmcMDeTbCT3tZ6yT//U7EhJ4qnJ67gRzQ3rP4OHLKAQ9LsF5/QpUVTUg5hDI
vJL7seMLiqhl/rApoI66U4T7mf3nKEoHVj5ogAuIcXGUVRsgQbKj1YNA/XV1
bLPTFDnOTQ5KPgLGfK9S6VNgMAp4qBovuyA612GrnbIS4eKTLnY+UiEwB8y4
TRmniOgGiDIZZ61D8LKcsz358ghEDnc6ZTBqXdLjSUPFDS9Y/OpMzKhsfCFh
VhcKMp3sX/WlO7smNEVj6/Kkh4t0x7qr9bwRSjoubjlIgkfjt5pGaqGURZkh
Qh/3vh/uES1rpD7E9vOiLr7r4VQS3D/D3VvHtqBAciQoYpGIBUJ2Oa/JuQ+S
POy7kR9AdaFx3/UepgCzRMaG1ODA9v9hm3qk4HcoNIC1YyMtw1UOZOxn+3TP
qmbd77KFXJcuVNL2pfM0vSuYTmS/1m/As/PGvkiiFizudTIemqHj4cp+H3xM
mmDTmakqAxXBqhs1KMAwnwwSTDfp/FY9eaS2CqWY3m0GpOS6FEzjlMP9zdbY
ggugpDfbXqX+xP97V4UaUDpJrY0XGU05r64GaLnD4oVMh3kB+B5fsuSZx+mE
ATqUZqjoMpSnU4PcJKlDn+eFZ1oJB1tqvW70WdDDw/41GVtmopkXg4YX10Og
r3I1+F6jkfNVjMAn2o/We4A2thFnG9fdNHoOqD3ZG2MEfbmPDUqvnzIcjnKY
h9gh5RZZ1RbbODrVYKn71tIOt1nc4FYfheFaqN7VonxUwrOgDNfXEnxq9iJ8
GnMd9IABpDvMBKvT5mWjrELCdG51yeioy8K3h5G7s5is0xcJGOzsh5w1oJ47
a86r5J4dqCeN9bwlC9/E6T+nL6EhOMRHX+nJ39T9ticNtZt/ACEmHlQVBNG5
fXzqI1adajnlIc5d1JyY2ivgQTsjdSccWUcE4/x2oQL5DlNMh2wtsnjaIh39
9Eb8xmNtl09zZF35DIeQigTP9QB/8vSbERam9mGSLEkPrwfMDKJGbidu+7MK
15lLGGa4LnhxTbsfbVt0SfrZBErIHosGURFC8xGlKlKIB91UFgg/C2qSY9Z1
RHoTaZszW4fixcej8dq609aItYu4qRqU8UhKcNNz98djFcm5MGfDWa/F1iD+
kfHFKi8ucYDcIfxBLawNanqY74WzVw8754p3SgzJcgrFQjf3xPec6pCZ0Fbr
NcFPkcgkqYOWD1FjW8ltSleUUvZoFHm3khbFTaE4y+zjzhdkMBHmNZjC8vet
oC+BIyH6KrdeqdlK0ZKfC6t/SC6agAThpfC7tCWpKPREbAxYbUQ09Mi8H/Bx
SPvyHehUnAOtPxq4PQzHpY+QGV4Z/n+vhT9A+I44X+g9kSiyiNeDKUM3GRjR
4JUR/V3Y+znPWC8KG+Tj5C10JmtV5qASPWh6v2XzC2NZLw89G/bEzPMU44j8
rs5G/i0XVvSeqL7mgtXR+9yOSUNacdYnJwL6cxM5/MkTYEu9QHkn/gOwdeZt
k71NdNbBkIDBneIBcuMZu3ClO5r5A2liSAGd3vPefPP0UCbxCcWw1Oe9BL05
+G2XAxKMajTvTf+xq5QkG4OE+SeN1W5d0cHiKS0JuzkqBRbhQNM5vPJVhYpq
fphm2II5WEVAkdSXJT8XnXCZbK44SAb8Y4CqqJh4MTmO8j7hU6ikoQWcTeYx
7e763WJUVJPiQbsmMNeseMEF/LLZTCTEB2ceNl5KFs9uMDcDO0kg7zAwGdyZ
t1t2QPjZXLF/vVkrs8lhs12qfXY3H8jfesvrJXpdYssgHoE2ZgzPa4mpKMBk
Hs9PtLD3QPseL4Bec8BVgK2Zf0U/gw4zWPtmD4/J4J8rXq0HkpH6Gl+yfY3/
oMAFf+ePQEZCSa4Z7PBMoiodNzPPscTrGfDM7W0RKL+mwKf5P9BDB796psDS
Rr5GcwZrKmalLNzoO2sdyY4roFsMknELoHNF33Gf/ThuRaIr2gpA70Ecgkyd
t9FlSoWmNOos1EDyOewnx1JUXv5XieRQhygHEQDZD3fV8caJr5cGw5FWM8fb
qjTFG9qI6IW4MKUH0/4nMO4hwE0cinybI61Mm9NB/4TrgO3U9wAVd7cfmNFX
zW9dSZTK1TyZtMYUj36t5K0HhYSpQ3G772U/6Lg4/TI6Uy7PRLAlsFJZLvhY
Hz8e3zJ6gglQlKv3Oe/2GkSrq6a+2Th/lpccXf3yPezXJ7y6szNt+/CuO+Dt
w76H+5yaxEttGvNCZhyyhuiQX8vvajIQHgAc/zlaJMjvHoy62hUirjv7RnPi
kSvV6yiAyqi6mbK0AFwfx4eA8DjLvAxQZDbsw+eh8tLyJm6/p/jSzQzRYrRN
iDEc/rs9e0HJwOYKANX9JQstQ9//DZBD+jxYFhcc594fQpEayFJwB3l37dAu
BTmvoKApmsidBZg+tB0doMIIXPyWNa7oYAq0Q5aVpdbeFsFZuSZwbkOze0uX
qo7ek09YKUgLVCZ4B74XNjw0CrhUkVE76ZSgeSsUrZU8uLpJKYZDXiKoXgNt
4aJ54Vv4ac6XRAJLaeQEyJ/WU8kKmg2JmDA8uaGQ36CkdSLY/J3Pos9DvXnI
vf20oASqeVBWwimu5e6I95qLvjkYAAqFQQWXTE4YPwCPNAJMJxm3Blg6h9Ux
Y+2zN/Vynd4iLKGphpXgUq4UIFAJuK1tTEndrbzqW/KjcTAtHgVD2P5ECjNl
zROco1/0LbVmMYd4XFj8RuLTc6Bl5gXuoltE+IYGgfHalVBxsKkf792DXU1v
rQP9YMbePx9Q34hbVo/mtU7UJlaJPw9b7fZJS732bomw9g7M0V/JVKbDrep5
eVcgQ5JeHrmuOXb7ub8NG3O+d+f1CgKdFzpOrtj5L4zZF2QB3+iBZ4iGriWn
x8dfJq2nlmUvgqwgTYY6f/21hwfQNfgDyp1VpQKOHrHUT9wVG8AsV+0ptAwm
sgDBZr9d1n2+0BLfB1/9Ul5Hb/MzyudKW395++IvBqE2n5OLg6RDlxiBsLFU
ra/NOOq0FI0Y1RdkjDup+Ki1ZNNKutf/SYNlCqiunK3gGZ0c9qftxohQKvPL
pxz/yEDzwn4b8NgMFsFhZD/hHgktpR6l3Fibbvi9itGdKg4r+sWC9WxxtFcD
qsxBprjdGCc4s3kFUPRF+VaE1qWbZs3ggTk6ODmFA5VNFrDn8k7MsCLm8TnM
WDp6zbVmvx01jVYWpohBxAqsYHrHc5DGJzEEkipsWe8XBAfrvMGnrckMmMJF
SBowUhz2CCKI2XzCQEGYe4+ZuGj+0zRbyK67VSVZ+mNGUNQz7b950uYPGjIv
MB08kSB6suAKbCt0PvtHvD6kPFyk/bmA77H9JJdf7hB/a/YzBtIrWAL+50O+
KtszXlMA46cZVoQuv+m0VoAFz+GtVt5bI/hjR3FgQPH/joduprBpLTf5VoqB
r+aTzMKconwlUAZDQrlAe5nqSls9HsaTLZViAMIPILuIObnmCGN1mkIpqa8d
tDqM4RuM9hiv/FwzWLjA37HfnFI44Js+/IgvBGI3TprzZZMLiIcnf8b10Xj8
LuqbZtefvD58LNAbLAXmiOW74iLemhSDX0W2Jp19kkjt+nN0wdH3qlFDyNZM
vevIRNx5mCI0p9aLMQafcUt7nBOrcB46vZ2tIxXZLy8qbJ+o/MYmhLx6mAm+
rygeBIph6Oj5JVSsOEj2GBvBAP36TRoLS47zFPk6pnjvt++IwE41Ei8Hm0BV
Tu6oSz+//o3CjpqBWehvQ25mb8qkAUtgSUh145nGT5OwGoGpTrm8+yQT1eaT
uVKm2B7q5k2bZkS5Av3L4RtuvgccN9UCfpJQmX0gpoUe19QjglmHGXcbZ3Z3
Akw1NVatYcxfmJ+9JJ36xYtsc/ixtimgx+V36frkfAdzrLCt6EmpGeEtV/Yt
wj5IKK9Ef3pJtId3pHA9GpJV6e6oPH4ofD3fIb5aQYXijMMd/LHonlYIq5PP
twjgK8RE1mtTo/aTm4DjNe7+N6Du2TDyC3crURU7C15d98zSxPUA9hvv127O
oDiqTIIJkyQoGtZcncPab/gFIfzqUklpTTr7yS8Bki3UYRgT9jYQYQsGy2pe
9BxL8GQCh3vTsViMsYqusUxy+wQHc+dzOyHrweIsUhmkNIY+bGq4CKX4kFk0
i4rhVEz6GIMXyoGMHgx58ZO+RkjkRaWOf9sj8rNqD+8htZTvg24IrxEhqy1o
oC4UNSYgDqprCbA7sDNTt8mcIddwOZTG4kXvgYSAIYrbQ41+bmebf8McATrM
PcxOLwY6vMAiasvQS4Y7cr2kRKZvtEJSs37QTktT/erRSXVtVXmsvef9B3ra
gXv1PGGeph9zfYeipoXPQ1znvCcCN+J7o4hGM55RCZuNunuUTEfuKfdy0UTj
+mlrJ7oHvN5OmmzcNSAhL3n33VmmeFFau7Bq5caNWwV3kZlkKQOz2f+Ri2gj
vQv4u//7VeDY1utirYsz/A6kwwOZvQscX5WHMr1VInGXrv75fvRZQ4D8zb2D
wb4Fx75s1Yxmnu151hZJDhvx6hqxK2jBU2Emkef3dtTzAjJd47bktaRXWh1f
4qo8LO03ou7bEj6KurOS52VwZsyBI5XXYYcvyhJh7FRHzr+ZWZK1w9KDT7Q7
mpK30REGkJjLYH9Aim6rgoLXsRAYxaGy8AelmhkNZtYLlCs7DJl9mmDviPb4
ZPdXELzApppZ+TN/GSb5dWZ/Kh1fYj47awYgvpRTUyNEbgkSHEW3nCyUlUkI
jzSdKG7fKfiH7432pqnz3jkSHTUY7YEFSTMYokJtHTZ2Jg54DC1t+NGHLdjj
1cvIIECvT0+owHZyWubsgSQFy+5fhlOnN56+LSCUD/fyh4kDHDn8GuWijqUD
d77+yRoMlVI4Mg0/K169NrJw0Wbv5CZor3KRFunpz4z6au29PImitA44orOG
dr0oFTmKnP0aC+IqMGNmWw6AADgNm8M6zhhRLty5RM0+WgRiqM45JGU1OwwF
fP/cIFZbomwkRkCSz/31+zAUaUQjfHg0m+fereqFtY/uSL/MfmDAgPz/XmRb
at/rvmHhFFYrAKITLUwWo9Xl7Z419971RxNAdNtElY5rMuixG2JbOWC7PGb2
snEr2dwq/ymeZV9vey78SZtuz29MHJWw+mrypiTTIdms69nFwMqVmgWxR/hv
lC9/5O5zuEagfjVgSRMGRiBiPjJfq3x47usaALsuT+R8fy4lPOrRoyAhjR8o
K+NsHcHuI6nrHGPbTvI8QJxKBlbJt+kG1ZQnlDOZYkixI1RYZsPAF8r/lxND
QXD6XufDroU0amHUUTQWXijgasqAldFe+C1j7kFnRgo9KaLbUWfeI68HM+l3
+voLVmMmt91asot/LSrvukAfkq/1SmgirUOkn7xfeOWz3P6I21Id9SwxBk8x
MBoguNWZiOOoluQ+LJyasnDrsH6k0UCZ28xtR9XzvwliyawKzOahB0TbXBPK
wKHpSPSAu4xwncSxzeKTCGJfHren6pZ8v5482mA3Uju2PC4/C6BzPN9C62u4
egqvH7w7nxXnyWrtID6WSLV3H0VqboUttpFrQ3VkFFc6bMQPjQMQqjvDL+si
o4L00jWW6oGI7t2dM1weRRZGDJVpSNW3U/4Y8jjlQqIJSwU12MJPfGkPLKjC
jk+ofl61HdCLlIYip5gWwbEzWplYVYfi63X9tuTUlUmL3AX1QOtk2csPcH+r
DJE+NnZkgTC2q12btcSUeMe/krbXfEj2AkRanAJuDTrWhI7mtJVBfB5mEsZI
nzIEGZVaP4GB5S3RifyRC73tfOsgxRJQYioddBJopKgu5TqNUXiadrj7UvNU
kROW4OT8sCmksTMqH2B01jWFy1SGprhn1bIGCX1Rp2xjaIBxAOFesLNhuH4f
OiYuuNdZd6bveSRNcwmWP7nG0zq7WgGvL9J9O7dfhFN2edUUbh78fftWJxjX
J8em7prmB5aibSfu2+YyLQoMdguQ6YFHCBC6f3KMp8V5lNRIeTVyRY9kAzuY
4DVDCb18DIx0Uv5rRn/+ER/j4x2Rnbodz12Q5mcXhfivAxKADI2ZN1Gp79qe
cMlOudajX2eu0yD3faqJgGFHEpT99w5JrcJOc2FtjGGAN9gzx8wUe53smzJb
eL9QAlhaHAKuXCqiXaOR+vMiTROOOz6+H08/Us85PBBpqtI0+IlEbzsummML
Q+d86+N+Ix+yXfKMWrw0RfHuKjD6dt6NqLLlGa1ILHjyhmAwhdCZcEqDuJr6
yx7O3ktjMGO5fQX1ZbFeaohU48/YoQT4K1YBrQQlWOig7ERjf8Rn5/rP7/Lm
isrN3l0NbkAHIRyUAnHQgizDR3yESsGHkT+uVTWma2L885P6DZ4e+4yZ82xG
ZeZHn1f1WCnsJjBIpLZxNU4oX4teAQZbXJRMh4yK05akBskXmjpuF6COmEWE
2uod4qAfiW8mKDsza5blyA+3JJlBZT0nx5twbE0m7n+2pZgknZ/3iaTOglGF
CTHNL7UcvsSMMlOphfQLhosRkxdAupi2pdTpL+V1ax7ZAX/t70mzntAydMz9
t0K6H6SVbutk/BS0tQYLNPJ01Fzm5RaSmAp0lYggQM01JzLpyoAmREGncxM/
THAPHqNlG8aYmuihiJ/IWFzGkpkXsfDsk4rBKEWQJQANtk5wUaYBtGYK/I7W
1TGzm8OeVGOJnRLTLZCKgW/O1C1BAxiwE4rYfaBMvpUGANeoHM1Bi8qc0/tN
RTbYRi82hcVYtWMOTVFAlFgBpBnG3TEmZycFxQ1Zrd40AoZNAmh7qppjtcsh
0JHV/ffgN76tpLL6fUK6F1ivvjqUgKXU/T9Rtn+FDfPkIhMl3hI5jLF8vIJx
vM07AaDGmDu2M+rYnDwsnhNqE2cikEddkeSNsYSPSj7Yhfw+TqfJXyt1BssK
Y8/Z/UdmnFClPqWug3SGN7K6WX72Ll1TzVtxOXr0Mu8H/YA2xp3pqQ64IIaa
TVyzj1NGGCUY/91oHyXCKO3DqpitsonGXeH8+4Q35NLd5kbldRc0N4wHLexh
HgWlzDDOKcwU+KNkRWCr9RflDdFDDeLr/Z96YAAlXjWL1e9Svfc3/2n5Vu9a
J11pV5nlwKpIub8M8ESmH2BXIqP+X6Fz+/0cX4mlR/kv67+gR9usnjXDq2/Y
2goWMJokrLn3D79giNCUkJJ0v5/bKn0V74KD+5uTNw9N09OsvnfFgtT2QdVV
EVaYD2A3OmbCOODbWqHq97d81aqeU0wyF8m77MPM5IpLZP03/xXDE8lS06lj
HAZva4iDvc6UobRaFP9RKm7V2V7JwEeza9eyBi7Rcu1xY8yhUQvnSCPFhBts
LmpUT4CNji0MD9/uBF3C21ovbzIEZZAu383wvxBla9bRtvxMZqlUTvNpeygh
cnVtUwsBBYGWOncgLfYIbWRqeAh7BNW6i6nJ5+7uzQ068UQdOskBaQ1vQEiv
PIe4IOp/AHmpbuKrocHtdwDwiA3Jg1vNspH/Ad8TWINH8nzLzf+9GWKuUuFz
V5i9tncrEpb5Brd+bLsso88Z8BMO8CNr9vhjedFeOKwqR6iuBZTJbah/bOk4
ze/0wRW0Rt+eUmqOw1NAICfdfit9TPWkgcFMTQmExzDRVyA7xuNic9sGsZ1x
fiznp0mXxzDZo98TwqbE+e/C3Vw+eTFAvSLVkT5olRZaIPYcqBTqh4jcALcQ
C+1yknag9Wp2aNofQ/YGJ3P7L0zSdFXiB8jWVfU2TGoWL54XcJtjFJdKtIiT
5/zb7PgCp4Sxwxs5zuRgAo5JQa9snTWp/HItHlniMKEw9offTdPLjbyPgTIl
wKSDJT0KddwgkrdNnHrtbbhWB7KXg3cNR50pkD0D137qb9R7blEfHzOXoKW/
aAMruWaLTVBvu4w4s7Bny7UpeqrEX5m/eEOzp1u718NiGpz2Ms3exbAPJHcF
Kf0XOB4GjUQhkYTwhcMx2MOLjGyXjyUeip6pwAVFRIjqw6GTmqEK2VnV5qyV
iWZ/oYqsv/ESRfxhGyjt31gpxIB+/m8RC+Pw+YW4d71gac0mdws347UfuGA6
DLnK7uDgDKgRFcVMbp0pdWlbkDb4mJ72PT82I/CNzubMutlW5omNKWlFETnW
nmz7T/urXSFZyJV1Jk9cnVkup44m1VP9PPpNPH54yUGXe5LWKZjJM3QdaSrL
DRILCufF1CmKUYJpmUamrJuaBfmUAYDg/JIHYbYppStNfd+854Y8N8ZZa6CH
uoWs6/1thfXwhYFD6CwSn1abYP4j1zO4WZspJerf5wC+KgIBvuI03lFhI8eS
V2JyVPD6bkhMiPUtWw+OAuTHq+fde9sqGDRmRuLJf1mtod89nPo2S/N2iXCS
uMeIl+LJhi2Fsh4tZ+QR43NAh4tWpPSUh5V1O8SCvc4H5BTdGyHLMk9zjq3R
NoMEKTTY4Nqsx6wJNVzeEHoqQ3q5F7S3KjNzzB9yKUrNTtUDCa06SzgWJRSj
PnqV1Z7ZThjILIlittlX53MaOOawDnA9Dbyk9ulZ/PWumL3BNfTyhsxr8Nec
n0dSIp4Dv72xREDMhntbvCuB0uChJ7CnAJilR3dfGCF8jDBone4H7QypzesZ
rgIFkstT7N1vxT8l0nNRpUfBAIXM3aDujJU4gTtkYYAbdzyV/nIahUrU3nQ2
nI4xhaiya4R88K8m0465KPTj78IjB6jHHUYbAWi+XnnjLi0hMJd+S2v/colT
8eQVtTU2ZEqYfcp5V6FtmuiDMRpDuCVg7bHcKqgjq+bTrMgHxNksdfjxuJ6n
xwbCc7ICAgj8LEuqTLr6fSifoUYmg3qWPiBCf+crjWl9AjEegtYQgfjfGoVS
An/xBh2RdACPuzDhbp94Lx3tAftArcUg65MBInN4q9irkxsQraM73/KPywiM
fvBVdP1wgM8mMxbYFshQ2hW97asbv7v39T70fzgDjogCCQTkhCg331nsmLoD
HfBIyFxitSIuEDzJdKLEZbKMvfwFo5zbNtasCXPPUx8/7cZDll/38efeMVUr
EB/qZEBMU3auJdFU8wr4T4+IfItrjKFsWpXNbFRON5kyx5oxNzJJPQI0ZhnF
HWAy/trp6cubFxd8z3SDZlmNJEBSIHiFqe/WoBrWeDnP8Im4T3AGikzLFiZe
860T1OKE3VVAXDjldCGP93fCpL6htds/yg1SnrS85S7whecLJQJxVpmcHbdU
LlTTkdP1Q4BT4bnAl9EGVq5msEHuS0Nm7t3M3Gwwp4XNPvN7u/GwTzxnnLXy
JMHOb5S4vfNDGIa50PD18x0SFVVVIagcyKYc/XdevLRUqpyHVe766iTh6RiM
gD5GuR2tLW3Mr6q2jmvUmeu9DEZlTb0rplZtSbezF6DAbZF/0PcmWLtg67sx
tWENYTQJFCvPc4D4z1h/VR4N4dV/w3jkqX2MNzUGMotpq4agB94tfln1uT1L
6CzYLM2uTfNMXw6XROaQLr2k1H2szhEuJnq63V21I/wfvOjvmB7t643DVgvQ
IYREQ1B14oVmijkcLj3sIaK/PyzJlo+qJ02Y3u8uU3to14YfqsZ48Bfm7cq2
+9bj4cTg0T54RgFbwT1hUB68gUUuPRe+TSKqWJK1mwErrB2YkSGaQ2sIVz0l
jBUReQR8t+fGg0RbQYQyaWBEk48u2uBEgvYsbYYGXHLaJv6N+Y1A/BuQb9lU
VWUDXw8/DcMSTdo98CPRbq8+qLzpdQVH6cqkPdVm8r4eRtBXWFzpcsmulInX
GboIgtOOeRWDUstnDZMt1IVIDsF57KHUtPEAfwcsvA7KBbp2unRoQX2x/Oyy
nztaqIBmA0q3/A9HWF/AGfxnnc4qHkbHp7KQFMs2Oe9j4X503HEA58psCIv3
+6h5DUd8dhOVPy+g2gyG4wIw9zkDKOnxaYrnUVaQUAsecQyRDKvTubnrcFLr
fGgabXgjPreVZba8QstzDK9pB/GL/7FQoyJt2JTaWoqO8C9J7fUpPhfbfjgN
Ff7H5RMD7LVYTOvfvyS8DhyrwDR2qvY41iZ4quDlAfrFTUFh5VvbzALIPe9S
GGzfjoKt92XOF8YC6jqL2MWbXRtXBPS2evF127rUqxy/gLwqHdNxehnWHRXr
vmjXEtDICrcda2ctFUuuGLDxXqLsqS6yP+pjjqIpNcSLr4aLObUHIFZnjBQ/
//susRQ4YMAPQrS164dUo+TI9c+HM5UWefb/x4I2CniBMV7J6XlG5jySxCzk
WQuZW/4qQTI5123EJKCRrCdQXHxnQ3bgbnTWPY5JHl4xsXsfSqP5BGujOQq6
Ln7k+hvpCuvLiMd8biD2+ptzNpPHGwWtw9Ej3+nrgRERrbsoA8rpzQl9leke
enLRg0DtCpmTTEChFXF7QStKfqIiwWAEPpySYzyi9JIeV4hVI2+hdCPxD/Ab
aqNfBgp2hgcJtldeS/iIrMJXkgNt1rpCYQTJLmPfeNQoH+tT6mClk/Ty6oDu
H8MF9UkYdVhG4nPlyAf6cyAiQ3oBPfq2DCER5OopupGXVDf6tPgaT9pdS6A8
ihsL4Y/G45xzx7s/WlYXMAa2iyjEQ1aBzSgnRFZ1sbnD+ZXvg09RfxXufpbG
W1qzm8e7LOvU1HgXeQmL/MKgkAT37hrTBaIR+it6pEiopq/7wVwtY9jtZWe1
9F4g265FYg/OIhB9C1RTxI80a8WHYZngjKy9P031ucuHRjyY2aKyUaLs+zPa
t+2EZWkCfviYQTGLZNjD2M/QyOe0bH2RvImC92MzM66YTNkxgeYsyYGWKY7j
3zvUoPH2Yy2rmLLZFatcCfV7YZ5Wsexgdm1924/G3xokiN6CadxGP4bzn1JV
08g4xaA8yHaJnmzqE4+Il/0aKe8cJvMgTGV1+19xfYJs8MX4Eg6781dcrMOL
1SYX+z0vltBFFH1vNKS9owYA00TI0NjTElaaQo/ovySoV4ejjiHsRwozO4Ak
KHxU2SkYeAsd5KyATmWEoPafPGgwlNehGZuy7rK4smBMVRFzlvFNfAGlVyvR
vPx6NqovrMVA/UBLCfV0GEB0stAGUw0gHMgDDayjeB/l2YR85wkDW599gJC8
ktyPnd3dPZYrF6jBdAuzRv/nXBfCRkFc7OPL/Dk0QSeey695iQ1babjvhhyk
PFApd6/6qMFhfwnOhlGZbtj0z/uNGEHE8d2lycl7OuuWfxDzn/+zEU8Sj7Q0
0BX2e4gdnTAyW7TXsscvWgu/T6d25UqHkb07568a2CozEYsGvooyMGhW3q40
z0TimnNEOeqHbHWHMKd5mf402uXgOKHE2zCdopAe1/BGMKkCxF9G+JUrieqm
ujP27ZW4r2AFwQJGoZ2WQMu1oV0s2ud3lphMRHhaBEvGzvl/2fzzPVfIxUuB
bsgjcAX1iwe2VlwhNxEmON+QzBVAZ7b5lFtPHxF6ONwqqLkPfZKTAy67Vevi
lu4EAQqwbnaR7VceHDMZ20Y6Yags6asVI97OPY80pc3hlQjBVXIuiEXJMeIb
6cJYyKKhetbb0N5ipsTgaPPi5iv+sFxF79LlApG4lzrSubPG3lSWzE56PMgz
o4GKzI7gvTqIFMK01vCmdWpJ3q8f9+l5CXFlnQJHWntwq21VHod3nMRG1ivu
YnV4NLAggOq0flzJQabcnFZFO5SFdq0JNKdjCZYb2Kgpp0KjotrqrEq3ER2h
r89mnIV/5d2h51vb0ngmHivDp1k8ujMFewodCFRG9xT0xQFJk/v3pZ4pvpvS
sp+G8bywPuoS1X61HJiTcg56bKhNRsfioseMTFtRZzQtCIF7k2LUraq/RBLu
zzsyz9qoFotqTwgt5OWyTj0ok3V8OpJGKd18qidCGKlTt1Nhj0EMpJUqsp8U
9z4sa+T/0+YM0pknVTv2fNozBSbmxVZTykWCkiDbZl3QXE9dI0vUt79KrosT
cUlD/5IHBWqw8/+8bBE52P1evWZaL5ilsMtM41Q9wrOPTzbL0BbMmawjoNap
hy/K/hYlngae7xA3QqTNrzJ4vBTVc43aq3NUY3OkGeBXZO+Yi7LhBpYGZ4Fp
vuLrQEpEWaZmU/T7opt7nKFc5eHWwAx4vjBlzJDk1hCVz6cqXSQWy6KFDT9S
rORQGRyZ2ahmw+rY5foIN6Xrhh3WKoRbqd0w9Teqyu5VUObQQTZOYH9gdKfV
/ZD0OjisjkflyteZvr+P4SnLQ4q66IF8PQO8twHsU9Iw8bwDfoOvF9xaO3si
6QUFpvXIdKak31Bufp4uC2s3+QlWJM50LYSROIEHaGTJfj620i0ircIj9FBU
+mwvUBs1umONujD25M7zAZ8KKb+U07V2HsLWGKfXqLesT25vujzFoU6amCYK
A8bjmsmmPHo6c8PSNuY4Yo0zgoBKlrsFbe6yuMXps8vmOAffaRVYjK3XEbgA
CbQ7bD/cZdUXxt6vSYg8FrNETX5Oo0Qul/PhXb2XU81m1qkekOEN6tcME7qZ
vbt8CyFy7hOIjoF25MHp4Xa9OSrQSEpBhs0h/fszjGgyJFcioTLjgsLuP+mq
XBrnlKndFcp6Mnzb55Jbmozj/kTYhHiNE/y4bUKKqTNSg6lqWVZoEYrO4tV8
WJ+xpZ5reaMOuGB7/oGJ5WHGdsQj9ChkLY1vvg8ahzJCaa+3bdStFu+Ww1dk
5yXz9Xb+mTDmzqMQ5Cy13k19fwEW0AoXYWZfhCyFjUgUILixsUYWYXBaL/YN
WPJGTRiNtRQIQS+Drz3gLIYnr/0XjlltgF+z5TTBipXTDVkcvWJ4qtSuECeF
vzp2O2lwna5p2ZE8J4NQ/pIEdkBEOcqWsDXx8Wz4GM8OerkzDhx7VAWtS9wz
rWvOFvSIuDr/VhHoc8XOM6cmIRluQlpdhipsPL7RZhpCqHxfO1DVzzc3avv/
xa45iuLATc/AI5YZ0STIxPeK9LIq1nMpppajCgdEQvyNQgF1cCc1nDLUlVfx
1Ath8VPf0Vch0p95WFxlHObBjds+a7xVKQ7vSK0VfN2Nt5QkJuyRUoJSWWd2
TxJSuK6bnfonF4BJR/MUu9J7Tu8CBISDEUPqtWanngY0Q1aVkC2a8Uo623zk
d1Fr70e3oGSyxgBGfkePzo5BSIJV9EhTTOFANhRrTNHKxxRrfO9KHAcrjXvX
UelUJ0uORRFBw0uIaUpPUFI2HDrGKEGdSmGk6TWiFUmSBQhycFW6kIPv21ud
qwSFcDdEVDDFf0oBgc6D/sY66CNSwLozJR0NCFYJXebs6YfYQMH93i6WtlTc
daBpeToY9/027TwDR3HykeRfuuMbrzQOBCb11cnadB46YOGNzK5iW138Y+WF
gaLwKOT1T5kIW3FoG34G9bJfLj3G+gggcdLQfcEdCNN3WSWel8Rr7eyoRaQi
cdVFNvy+QHd0AtEFGlQqOkPqQ0EpkRqvVkznC6hj+685yxf0KrNlK2gnHnSi
ENRPPiBrq668hUdG0sSCNKWlJirb5a+a2Njn8lL879RL30HnLz/rQZUOmPhN
zsCIOZ1AEuYVOJWk8SOBZtog+37UJ5vs7BZxR/iO0KtAPiDCp/j6oS6k9R2A
ImrqWtJ+wpwGqKe5NHT8xsBmQwFsnFSiQCZv56c1ukipUZDl2l7CHp4gGHnq
62OBwWCY1OsBu/n86fZ+Bt8dFHQCb+mzhoFQwbbJChz9bQD+/hpsQArmqh+P
OLFSRPXMvgtxIsFDE44O2htdY75nmzOK0w0x+ErNGxyWhECHqzWlAOE+4x+P
NZ9cSoc+U0GybcJN8fMeUnoisaQh0MMSQW89jOwI6ybTX9hrRgsV1225Yy/6
daChZF6Cx3m2am1miEt28qr9q16B5MyQL5+xFgqOlvjSnFjAxGhpuBokf3kp
jUilNB4NIHHCO29BOBmvQdViO6jWiz4UZ3W0NkK6EfpnTvzMbcK1y4A9CQ8f
ZOOdtVIgsrVKwM4P4O0NxN7i3Z+KHq0uz7qz/CJrT/4kPfSGD3/rBTHP7E6Q
C//0NITUlXphZRb/ZerSoy93N36YIKwoRAwjXJiVEjZnWsieFBTzwOWmpOFo
upL6UWIJknkRUVN/A6d8OfJZAl0T7HeOvWPLrF+DZSwKfnSQc6EoVA0VXncx
OX6DZeBlp1pBRWx1iyzduxH0M/9Qb2KR/o+G6svpZLwAE0h2zkEZJxinOJCH
i6w3NvzPHUUvqB9fYO1HAYZA2KepLzyeQEzo+2re4gnNmcoUxk36heqcrVlx
zsVFSisBsRUsdwxFz41UWsFESA17IirdL9F0Fx/6OgCv6NXWVbuZlHp9nsMY
ry83Ur60QGNGnEu0hcunOjyVZNUIZ5W3F+cVCks8JGodlqZAzhoURvQmnPjA
xqaafxzWiuKAk6cXyeWHkqOBlwDpjJrnZ6jlZugHt95RNSm3RBEwY7YmkeD8
CrglNDGVLxQCif8BUuTZ4JA5PJ6QBqgLNFDH59VyMYA6neA3V1VWtAEONKpv
xucoGDzuLy5rPBK0oBaFBY3Ev9uKbtuJrS+sj4EzFLTJAM+hHXhtVl8CZds0
lldWodnB0F/UtjsuRyC7LVkDcr4TVylPD8VZdJ0rsr9R056WImQ0SrSKKG8i
iwCtHguNhjnifEbfSzpplhGcj5bQ3eNOEj/LSKJB34uMFtLGvO/cntubvs17
VCzUlNDTNCPXmEQj6Nkj9S7y8A+ECjD+6zWWbW4LQzkIYoxydIRKO662NvAS
cdbDJm24BUA0uE87mYV+jeLthV8kel0Th3gdtJaB7l7PkhxOPSQW3dm2Vnqs
y+6/5e89EzFchlkkKWW9vPAMoUDBBnGekWFwls2mWZCUQPn2WG4eGgpUDT+8
/y/tTy49amBJPrW0paJx/PmqCYrhPN4+maRSoIZX5ntb9CCrq4xeq5K+Ww53
xrWkBIdcowzj25jX5Vcn9YGAKkUdgPeCnv6BAs7ScbF2CU0pWhB8yLPpQ7tU
tV8rs71/JD7XS5e0hp5Djy/sp0aQBbS1bPTtQgFQ2Hz9f6H7Bobh06Z+uzky
ELZqaG/kwqD69SQbZVh0xZarelSQ48OkEDTa8c9XOVqnyHiVlyU3nYE6bbSA
4KvoVmKRUHIrMPUo7n476hTWnDHvCezfejxJsu6N4TpoumHfqZb2dZenkBg0
ZVO4VjHe15yOGyTbSsDeKaAMGmB+oZwu/EubR/i23ImvuJf+msCu6ThypiTO
04RgL5RuEca/zwIFWLdkYSxgm7esqkjdwm3bbsWRa+Dksdde/552x76qHE6p
Lt60EwGIa1jJY7UkfmivPFURd0G0snxaZtXBXZbT5WTxtB67hGcsastpcnUb
yn+YOaHn5F88FUdulgBiAWJYEoffAOC6/YhWIHBYynbZHuB4Lf5infZnpwUp
evhioRqSNtYGRGxCqPXa0sWDB6h6JEOuxBYqFamh28TXjpcMGuIJVnWcIH08
cFPwomi5LIa4xq3Eh1Ekzg7OSMXw22euRnK9tSSSSZzTE9aZPhVpIZLHgmMh
hbxM5yH3Adn7szgEjSzhokgcuLPgIKAln73bmbLpy76KIJNvrYCwB7GUnaic
eXcDXqz4nLuDulscg0DXmUDgGgR7HNDNexRd046QMk/CMI2Z8katOg8mvgfo
iFoogNcf5I7aH6gFT9aA67icjQqD1KnawkKDGfh2TZXaiYmcuFTG5tFIIQmm
5hckYuqFjRrdOOj7vn3M680NEkG6mespSk/3iXlw9JU41FQQeW19RQ/jsGbG
/QrUepdLWWHFteZC45s33r47JDDSQrPQVSrZPG60AbveVCANXjy33xU2zWJn
ns5o4tt/LjQ1/9zQevtvGn/EP07snn2vFnIpgBwaxPydyb2Q1NLsbj/ePOgS
cK2qBBUEe+O90wOrWRxhd5KVJ5UZIbDh70lnU62nCgixOt78F8iSCeKQ9r6m
yeooQNj8vjgVGsGQXzC9/tPRv7SpL1Z/Pq3G906xZywU9XP9U4lObifFlCTR
2p2L3tM4e/zJjgcGIMXizy/1wDWQfeq04ThRr2q5i/jmdciFdpDnGHAkaQzm
IQfO11XfVy3du1iCU35LKTU+MD3UPm+vVGaRFNKU3ieSIZDd+tZW746I3gk0
x04yocH9f0h3w9TNSX2TSM3YK7FBF7GY8A/1yXrDlB/0IThUqECinJ84AhLG
MTturtnVCBTIr/PkKzSLS1MmYS34Gk8CW6TVSFoYDDTHRpawjtAhzwmGEg/J
uX26dT/MwlpO7sKFrrHZmO3LqQ8Q8qfN3UL84sOfP9ACuDKqphlu1vradX/b
i6cgHX7yRdGw43tmHOQj5FVfxYIzZh1wrkjjRB+IafnTULRpVm8vPssYjYRD
MqyawjD/382Zxqqz6SdHdQMKZQdJbEJHSt8HyiijNQZzUknZM4Gs2egEnVv5
X3cPyEsVYndMc25nQVZ/5C4z224IwpoA7zTCqmCGzQQtF/5aTwjpZlhQOEi4
oUQOcqScRnUcEI4pgrf/ko/Nn2tFPXhopIMFi4SmUbJ8nzLkOTw5DLzri3kB
Lh7o+zbx+wbE576epwIkK+yJknX0D4vp0cwJ0SpVQ0jJYTvxj3ROBQUEFK26
G+mso08IEBNHrcOaAerdR00aulqxHfsNaiMieuU2v32wcwXu800igdslqjv3
67iw2+VOgPakN4daLJrZRjrMvYeEbHNPQFKbDwixufEqO5uFF7r+Fsc8v8UE
5VmvpDfCTFhjs1Yrhgr6lOOl5i1wv+6ilXkpU1PEzaiwHtahF8v1Evzr2u+L
p+0Xq7WL5ewFojM1ekFVw9roHmU2NyQs95CV2Sg6lgkvbJ2di8rY2p3yVJEY
jpt+SXdaROZyJOWWE6+CQ/GemCPNuafudGlWAzhYuEh029QfrtX//ceACbEZ
sSlAy7w4QpHxRnYwhxCRsete/ZDKS4R3+v70YYxEL1TSQTVYh3ArNz0PFYon
v/BRCfqhOvpBSAuOAlGuzffD8Nz5uze08TjvXkwjJq950MHNl+0U1ccyfC+8
YXcHMCO0sdhypHREWRrgS/z4pJ+ebPCmSfFpPim6owR6f/0e8OelGH3ZimY+
ZfXg+ESHobCWPQhpxcGwQxtC+zpNl4z3BSFjuXgjm/TvuIoSASdRMzYt+2lA
bmZ3WMH7jMLydMXai/srBm8PcbB4swFX/3AsiaUB6IxA8oEaob7cstFSBNnq
kgfdDXl1YzErbhn7IMTp8xZa7ivJ9QIgKa8Z3x3mfxWawd2PD5rbebF6M/0l
nYagonp8cjfuTbRcxQIRi0GfcYPB6knvzLprx2xT5tlUFwvZTyxq/tG1gYPt
LFZeJck50wWZzTN6VcTle8a0V683EXVCF9aqVg6xH+FJOnH9UBd/t1ScCrkz
6JJaRyY2XMRraLmfsLtCEN7UTadIKEAsaDMFdS4QZxc81aGdg8+LTEbgeEnn
gYRmSe8luWZ2CcSBeFmpRcHCousBGgpb3DrjlimdwKUCCyz086iJnTIsdcGF
2GmpKYk5W3AUdcbFZPjq55RUlKz26xljL3QQkPOb5XqiQWr5gOd5Vfzipjar
xC1e5XrxDCxgITS7kwXDctoVarOVlx33WhG/Hii5qBMsVK9PgsOle5yXwFxn
NJ95e2Ib2Bq+lH92MxLZMj2FaoLi6tQ2gd5z/edY73dHYbhemHZtyL/J9hdC
gvcpjnG/6+bjuiaSxzQET4ouTgkngaYmDDJSEYBQh8RB74f/HqpE51HX8DJz
XVo1rc5YMF5x2CNWUc/wLIzxr9msluQ5ACbx9k3+jZtSQCB5k0cIT3DjrrC+
nRkjuJaEP8eSjz99fhZUvdZB8u6Y+3Mtm7bC+PNpuy2tgjdixGeMrEfYooyk
0Wo++NYVsF3SvuSVxR5YtX0uyZN6syQXTqxltBtQ4wN2JYeXnF/WoO6eaWG4
4XcNve0+C1OPIUmdWfyiOI59ddmfcFzOc+tZxHL34eONJJCKe/OMyELheIVu
u5eAMn2CnxMUPJFmg5a2IdMVjTQzUpbmETw5DJ7ee7E1gTx8HHNI2H4OMW8u
EWcfbfVMhpzKdrfe0bI1uSKP9VQ85KjirymaWOiP3jox4jz4kXid+3u4S7uZ
rt7xSLEAT6myFKRQPRkolc5bnro4x9nxxvtg7KFVZxd4DfTcz1S2KXRVcxiX
hBSA8tA8J+ZuiI24SP73J9B13JTIMP4rYUKK/Mp2PVMasUg/rAn8KI/qqzym
JVh7UK3nAN+HGJlAPq2x7Ogjw/hU9P9aCJ11+lD2D37XfvIBj2m2lwbuaZYE
FOya7iR2zLglXFL4EP9KWeClRlqrW7R5v48N1oyPIFEXO/YOO+DeW0DBQHnf
wDoDA2RJTpM5/ktnyP01Wjnm+jkzT5xUQ2h7ev44KLt3W0DmStWeS41CaqNO
eAuQRi3MthZiRI6b8uLs3O8ZDDxcYODy3gjc5CyX9ry9vbMWW2+CrgJRRkw3
q/D0TQXE5zlix60ACLCi19Pv+MNcxgPI/UZjJzc5BGukAyOjY/3970VJTTS2
c1bWwV72RsYCDzGFe8lzNP0xioaYEJlcM6XSEjy1QdVqiZHoi03bfI6xHDWa
anh+qW6UCEetB71UFgmQu5+g59/SESf5h77k7/R5vqGm3p6F2jP64I3E7qRT
Xg5IJ65e2H+rdRmsAhzCMw++IWFYwigM2JxQGtO/4oCeru9w3yJOQvcahXn0
Z585FuO0At6MXDHxWMMQ1Qn2G1Yl0K6RvWZQo0VTHbCx0DKOlgy9IhMc/AnY
2fA45ELhAPCr9/J3erEZF4gKi/oZGRmPf+Sx+aGmUC0Nqm44j7Ks6cu/nkwZ
TokgDWqVOs+/M+VEtADOPIL4YNubFAuRlI0Pyhoz0fsyOqSsLjp2X0BjcUok
VnhqIrgMTDcp1mzJYj3PNmXdopRr5rspg0YjS9k3V4YCJb6cMXVxRByyRpCf
PdCF8yhcpAlFKFvpDGE0SuHh1h5+1/Hg5SqAoIUG1c1BD7D1KU8bj7Lc/KT2
fvyjY8E2i2r/mxV46A8tktxOiRW3eoeNo12MoSj1XvwEg8gkfN3lwEs+DgiP
VEFBQ2BfMRol6xLna8klCqE3uNGL+IaMEXbDxz418alnl5fLfsqL8pYK9u61
YbkQE0FSIDaSchXfUaYfjKxAQSsZfTepjSGiUByVOuYIH4XxGBH+uDJuL2qK
f+Tf+Jq5hTlNc9YPd85PMjrl1ukHytbQFM9FyZlyegc81iU3l0G6zhtVBrlL
BOTDBNPyw4ZoDPglRtNfPbVJXSsIfqLBnTdgKBQ8i9KCLeJUIdCGwhLNrJNr
PjmTI7GKeyJSnxJYL3ysF2NvSLJXPysFJMsywNiO772TWI8M3YcJ+b/LYKAZ
0TLmkkWZ0LtpwVCQyXunGX0w8X8S98x2tCH4+3XS82vtwQ7aBrICclix6dn0
sae0iRWTqdSO0OT+AHik4B5m8ywtMAHas1dxlym7NILTxMC+PRjtxskzJzyc
LNXlhsjFXFtOcrs/nf8lu7oFCxwbvLL5cgY4Ix83aq8NpzBrxw1SN6pcJsK6
ud/RHCjZ0Ld3HSS3DXh4AyQapJVZCo+ZSGjurGefHjdD1i6IjQUZVT8S5Lxr
7hO0qbWlPTe73b8pb36WwleuVEPmdelz0tdGWBFZmkxDWlCdEaR3IqCUlQpA
pB2Gj0Vc4Z2IZgFb9RteMpDCftcbSoitpbEkwoNVqidkIUsma11aSustr0BD
pDY7CMZQQbBj7tNzhRECIirgNjRMzUWb/5Wp72nmD8gXWurr0KV/UMSZnaV5
gZURv4eSuqM0rZ2k6B4Dpo7JnyWM8A622hlNdH+JA9KIG98zIssK/553POZw
nKuqoct10cnEi0VyuthT6asReYVtKnVcl+/QeeVBw04Y/OMWEvg0LYKAsR//
+7xI9rIG6FO+FBZhqJc0UcqGwm88oJ/737jitGoA8F/acoXNDQTk/cTIABaW
6Q6CYAf4NSPs5hS92GWU86ILkL8jF/EHlY8Fq/LfGUN4XqDh+dVyGgdCnRUQ
IBA1YYB9392zF8FfoVVAD6ZYvgx+fud7HXMmmDUOQSAUeYseXcf86Dsq8MFX
gxxM1sPaYKhJvSgQmM5T4QVnj8d1/QupOxa+kbyLfDQqak/Kz+FMD2gF1luc
mw7+OqRsKhDV4BkcAu6bkK/rP08Dule7MsLsdkC3W8eUMeZGNuvbMxTg6w7R
pXE3SqyS92Sz59YdSd83TpCffzahwV4LOw34ZTKZ0suc53UPiAHff99My48b
LZ9QCiJOFYpIQYJ6yku57O2qoloSIBzLcEuCbZc7S6FqFKS5pKa1Ta7mYVN2
VdeRA6jzYHDIjxZF8YUNi3Um+7oSCwUt9it+S+GBoqFs9q1+gl1QTYwvXSUW
hSbRJhVqdFkJNCqBQfx90mpRoQ2SPfG0PhLkSODWGg69aJbYhi7otyxqOxwz
x9LQSpw04bGaVufpdqXUsXf9k79JhHGg5E+r9boPFjc2O++NJyL83oxwIVgU
W0VMbbPj/TwoUtVuJgGUC0jGN2phWAVyYt8uGS4J4DjwFadTv99AWA/MjJkj
rccfZmTkWDqulf7M6uKJ2lUYJQGXXSOw595gZnCa3houVSFivLqeRKXWiYSn
ovw3yuKsVScmicm/giHn3q3uBARKXunZIOl8+OekOlEHc8hebE08JgJSwHpI
eSVqaDL5SH5o+eWoVbggC/fDtwDHUdawXNR2eSDsoNNvVnx1tN0tAVzT1Ocj
SFBk1jjL/hnB9g4EJnXrLMaxMGFqZyPRG95Evb5XkwLLEw2PkMUjgqBuvk5Y
MHMJ1bVv4/bMtI2VUuhAeIPbNbyX3b4YB8tB/s/xUkZQyHHfDzG2agwS6MW2
fQFB9nSBck18swIv/4mpDAcs2rfVl2cj1y2Zg2Z233pEyvd33iwJ88LybFNn
3FXRsRUbnN9R/0vmQ0iH+ekBxNNDEoocJa9Uv4jovtGv4HMCJvsvoneb9TPV
JkyTFlV/KqiBlYwdiNe/4OJtcSEGoOZM6zceytS27sfQWOUpuraMC37Aq5Rt
J0qjc8b4pgQxwwiwM+/49X9e4gNSec/tNswl6E19RJqGbFRdXJEJ6/orcPNj
S3lnBuE8XTP0rdlH2kD6aIojka0VQVSz8cSeiEJkd4V+V5D9+rbHHctBPbzi
zH2vVM65GWiYNGeE6wZ6+KItU7y79oz/AXl3y5vmMC6oyDbHUkRkS3vskVyh
rhlypJkIHwlYujFI7n3/v1UUehbvy+bjN24RdK/Q25cWPSp9hyD2s6Jw0wYp
iO8Dn779hAtChLbPCKXRZWt2r0YpSywWregBrftuJd3ZpZ1NnHGxCN+EfO7p
kzltxv4t2R9eTdwUgWj+P4PiQC6N+mfAZ+N5BKaRKtpR52MNVXrt95dvWg0m
LLyML1SR0hcz5cOHmtSm66HUAKKtCAvxNHw4eHStPYG1qdPXkLFNShJ6DLXy
woNt1r7SWpxAkCxGxcZZhJV0TK53aDCvSvhYK8OdWQ9ifFdWxklqHPwQU5Cd
ujL8dpY9ZIbj565XW9/Pgy3U9ttq2i/BmOPabb40k0IB1TgmH/oZBtLdwdJW
XjclXVfq//dV4n6yIMdgR4W4FBoBvCJbmZEVNWoXEQK8TdMcxneF2Q/NHsTQ
B2UNs04sQHOnNmn5hUk5upWAnZpgC5tJXuX+ERRbHqbZX1+cWMXa32Y3M5LU
Y3zAfYvQzZxya2c735sVnOHzDOY4AnYCrIGV3BudJhfX+nxIxpBQoB1B+bWN
a3iH10gaTXOsUHUBun0OMVSBQesA3rf6i3n2kJMRBxRJHfDIR82mpNmvFT+C
YUE6JgGwHWS6XEeRqoo8VTMdolshh5dQQk5Gux3zkVsMl+qQp1/kjP6q12q4
HmPEx21zDJEpPd9jTeV6AHBxQGM0TSzJLjUatfRPEFC6glQd8K4bGkf8BZ1V
03pi7ohU0fucHsjjReQ+bIqatzXL+WLP1W9gdMYOURh4q9yKtKd1KIDUxmFV
3j3d3LZzWnydLmBsX2LjNVN922j/8nnWUTLV6D3BZEOANcKOM7Vt1Kapajo9
cBlNH4h6PCLOVr22HdWPDfp4p2qea6fI7JqMYlksCrqEVLJNfemjWquSvHlJ
pz2x4C2H4SjvdRmsrZR7JtiWkh68v6OudQMKNNA49h6tdex5S+whAr1uh/+f
Nzmg7UPjpd+FAH/bO7VCxUMBKwB/ePyiv9GF8Cn6+0/klk2aFMyg5GZs8q8b
B+Gay/ZSvLGFDbHiW52y/0G1j3AMllWx1EhtAXPnV99odTgJR8l9JuMvpdjS
HeYDl1hXNDj4aNOD1Y7uDLG1XSo5I+GGwsZ5uAhfEUs697j5G/7s75zzaFec
lZ07jVRZntzopI9YG1Eb09izAkKLfIB4gIuA/dJHtY8yqBT2I0Moqvz006SZ
9S2qUiEvDvlEmTd7pSR6qUY/ou6GMrZYDqV+WoPUnfqpz+OKBSMJGSXYaWaC
eIP6jnLPtkk0NY5NAXjxWzUIkzf6vWPDy/l4OhrZVHnhMVJxNoM0QtsZIe1U
ZBBWOkU3T8boVHGIr+LhSFiQj3GoYQ3cGpqmEcJ3zfafco3PaW94IL43xKwP
kxRSPwHB9AyeblZMF+WbBFkCrYGELg/AA7qevDShAEt6MFlkyRacobrqD+jB
JD+HmNeEhYqQxWR+XQ6DZ7lb8dM8amIGXa1+GwC1I2vJWpGgohTrtl02X4H4
k3i8VFnV8gssg36zmdxUobORz2K7tr+/lQSgJfGDvJ65FakeXD3WOTplw9ni
fzhQte34tMSPayZw/wPTtgWSedmch/CU+aZ0pl46ya6vrVFcuLcY0AxGbOxn
DSTWK9u071Tx41fkKEZu5Fe3e8bN9q8Ar9fB2mM62Fwr9Xc+1M1weRQ7fMyH
oX9AxQnPS8p36KL+eA9iI3aWOT+0d3N5Khfctv+D2iX1BmDysr2ZU54fMGUh
Cv1k0+hi5N/efo6gCDC219CJ9nE1lbT31bYEXPRaFk8DsP03X35L8YURcPoe
m5cE82ry4T31wPi+h6Vkg3dlIlahx5Ytogcg+uXFwGeDmnzOJPg+sOTQO1dP
824evJzvs8xKLp039V9nf5oPp670Mo3ztr/XnrmhjuYfhZ0J+eU5ciJ7sSmn
q2WMM6KhbSOpBge+Q5FK0KxtBKWiPhi0bRB8Fq9bgn+hgGmrAHstIBrPzBzu
XuzGOMbc6CHhLmlszHbpCrgLMLyRzUdom9fWJUwXx+DbnHWWNAb1dQXkPYEv
7sovGYChU6jblkm6+sxiKPEm9o7E0mE67ErvK617aG/NKj1NTTp4KY19KPVk
nRkGyj7/SfROA6wmseW7IX46ZP+VqLR5iQn7T1LY/WCsXc620YOF5kakV/je
u+pHt73mISSYUExwz5fje9173Wq/yqqPdLPdES2kk2sYxjtl2tR1pdpTU8v/
+Oq6Z+Ju4KXBaGiAC5nqqMSoCa+eG7r6GnEU18degmPvIrcdl+4vWzwXK9O7
4ufRQaFHhwsXgHyEITZ3GZ4GZEP6rcT9yEkqC6meou9K8TvqevblXsInO+MM
/Vx7TUbZTgeCq2g1oj3l425vRCyFsfjoxxbE+tAfnTXNzys6A+PxaHgnICGg
mWTDy8d92RG7cgBwC6A9J4vEIOGEwLOn98o2nkYF+v3T3OWDLfMqgg/J+J2R
tXwF+OoSmwcpEGMM+qHjn1ZlZrQMGKWN3accFRWIEt49roDsvvAqtweHIt4v
pZopH0GFvcKAjYZhiQrQs32OJ6OLwkI7230If+Iv4b9S01YB/zjSn+85raF9
U7wSV7WKd70j516t4MBuIvfDjr9oWCvp0dh8vs0D8DFrPDymricEMU4dBTyM
5aJISDFm1mUfJ23Ma3VilotAmOIvDvGOaNmFxAOouK00J+tv9OkMh6I0wqd+
Pl5RSN3MKD3g7qGt8xCj2nEs17ZvlF+s1t8xJc28KxdWU6pQDqg3ks2FrtTP
IsOMtXY94ZVSme3iEG7KNp4n+T6anI9ZTPFBOzA3IIP0FGf1BfLwYRogbSGE
kIZY/tDfPHuNm00n0+BvFx3Ac182AE8dhJaZRlPsnlLxWGuxdx34m+Of14dS
GhW7EPy0I2yNPgH4GE0lA1t80bQf6Dh34+LxTxrU3pHkbfW6AXMT7nX6DSZt
+VD0mq2oQ35hty2UV0p/85LybBMvgycbdzI16VoeBdq028yU3rM8QOFPBIFo
ge1HJxmwKvcKMu8cK/5+18gMYdILnUKWrWQlwOzBQZ/Uj+8aJ4Z16d/8NedQ
J3U18BjMCuX3f6669r55rUu2BvSmoFi7sfeFTX04IjhsdRULKE/RAgv0xaoF
KwP1c1zQWMWwbgKYoexuC+OG+kN8PFr0ayhO8GKDrdWwOxSt3DM86FeDOdY2
kAyjh31NgzAgYYUtOEjxM4q2GvakLlkhYJLyCKAEd8UZDyJDlm1gyGNBkf8D
reX6r+VR4rMauqFSVTg5ehlSxUSYQt5RXFmLyMQdGan1/jrWc3fMJ3RTfT50
A7xtExtgWIna757jSV25GBEK0roP4EHhbqFyPz09xR5LcJ5twPC79ZLJd7MS
agQZbPfaLHXKk7LEtrcq2mMpZ1DzbXJjlF3IIfvCFzeW67CLEQs7pKD2SMGl
/nSj/1+Rqp8Xnnh6Arv7UgLwPT5+udjhfAejBX+8g645FSU0JescImlaDK7D
PGYytyx0E55KBmy2OJvCFee1mKA2qYTJ6YBBht0eUM/y830Smz5njQ8BLUDj
5rRv3YLpwNetJmRkGGA1ZAVCRG0WGjodnoXRID2HTwxyM8fN3xrCKVrHJ4It
5nXwZPFYRzPSDk2tVeD1NbgCk5HpOb+lv3KPp33jeqg3zDyHUbeJTAz1Mgmb
9upxSE+NngdumqMX1jVISBiPmB9TeOBXb/EIoVhlPSxZMNVXG1fWIyk4XGK/
O2u9+VWyyJ9yHo5OJMK2B9GMo8eaPuqNhCyqNOI4SvqMAc4bFiFngJMV8DMM
HLL2iBilXr2FGIa43FqUF51EudOF8IP24pT8EP3mwU9OIZH8mt1DrhL+WZpx
DpGqeltNBJIX3/h7X8X0iuxuQiVObHosMokYFs5tVkmAP+YGnzi3KuDrYRMi
Da2mhTab/V74JuawVbNCmArvI5Hngl7s2CtEz2cFX1D3u89Rwc0WgWI2p5tG
JJj/UOjwvYCIFgv/+Fd6uNE9nSt27e0jloQzRlH9EA0eyH9Hy18bMFxTsEMu
+4slSwGZsm1M49M+5lcpnmCzPKdmfFKEJceOD/cfMzLtd1zRHYEYd1a25VzP
k/Ver2Pp/PoiWGJ7ORLdMTM0uuAQui1bCrpHqFX89QdW+svw9wqdkhuF87gt
0PRQFe2X8K40OxFcxk09grkGWwoRgS6T7JH4XwjaHZpB0qm11uMl1oinK8oQ
nK8VwnHJ4ksVicuxCgqPNWEwIm1iZSEGnl4pOB1pbYTsZDNhLF64YZOxh8Lb
IwUsoQgSXazyXRRFSofG6fZQNv7Ru33jBz/JTubeYIINa05vvsHu08HEr6BH
7Qhbgali232B0zDV7YdVULvYE2LEqThpUDF9bte3NIh6p+XpYi9jxoqyrvqW
qTzPuoannwJmi28tlw9RgTMA+YxcYNtreNLFKLQee5RsthkfvPtCpuBAFGem
g4KQxtcju70zqHCUkQfg4EodaFOZZohnW+09ookZTYmT/6MMqJF+ZQrfwKqu
A/2m+d41DRezYUTHjlvEJkD1ECIZTG/0XDIr0524Zr8zCGbazizsFdDcH4Af
Hcglyp0gENjq6eOJkOygF1ZDGM5SrXQpmxKKLAjFib5rdrDqW03maLKCzBcf
wcG13coG8gfMrDizkf56KyntDmprK27yjxI5h3wPUWUrSss2SvB2rMvnamvQ
QbxAck93BvUE7Qn2H92cjLA0d0Hhxk9G33DprqWWL+6XIBUQkSKWIHLXov1P
SJwAgUVTWLFt1gSvDUCrs4+gJqWkmsM5ZlvJQrFnXosslnkL6hJ41UAkLopJ
LDhTecEsz/LUBXfSXp7hMuOlsWr3GXngHTzriOt4WoDqwe6rFYCV455F10CM
U3TAFPsZ+UBfA5Ru15UEwW7i0+0j6z7sYpvymTske02mG6UFlULktoKPQUN4
HZ5Cer3Lom1kwCHgnlQ/l54BCzNcnRayNrpmM5wccIEBYYlz0nlgQJmsk8Hf
f2gbffS8ta8bwp2SjM2MCMxq/z2eYzNsKxn4tPc037MIXvSCick+A1nXpaEJ
2DdubHgiT/cIUu/9/Z8KW2vzqeKO4izbxzGLuA8GCfhhxZB1oxsiPSa3Ua/b
rNVxprDtlhRSzKChrqdmF584VTwBr/HbEaL8sJc+DMtysdZqhvCW1BlfhoMz
UN0+wom7bh68tsCPlEYDSZA5Ifj6He3gJHM2qtt3BQ7kpen+5Z1gS1wOwKxQ
f3VYfSG8ITlaQdX3X7vrJE0TUvgHtX78rN/YTumAxRW6ywgtIWkskSZ5C/yf
7jVTvxzZV4YgIl8ydbqQZRvhFyFDIobgKHe5t2W+drf0cjw7DZxlcKp/IFyh
rpSDabcI/0STq6/yfCr2qP0UVLouh0Kp95UALeiad7m9H2huIFlPcOR+LrEW
1E/mDIHhFRTvf0WWpqYqQ1IUrLzJLoenR6sGk2kVwm+ZId2QZWCU3WAT9Dx7
cUk10UsE/tk5ikip42agXFBwOyYlSlCJL40Y/Gci7xf2Hqy6Hg4xY7FbAdaS
2wXht8RlsyIQjM/GLNWpDOrvLlnxY8DXmZwnbDwnso0TNb91dTx6EG23UuJG
zPlgzk4DfKxuTX6LbP+xoTpKLi4qSmyMsm53KGoiZ2OsF9qXSTNsOcMWYu7e
BEEk3eUT6l4EX2TkexgElIVopzWEsp+q3IbFxoInCk89iFUqt5mPYfW3Wils
6o+M6ONoJjlvOK3PAhXHmQ9vPZGToT5hAHMn4Xtvdwmm7N5Tz/+m44YfY6XD
jUirfm0J10b6KwcxbuRdDXF5Kma3EqE1H/r1IvWsR7k2FpoxLMtUL9Ms+7Kf
yKZXQkHwmRIw8/vThg0nj6DOaqGKym9x/nCTK4FjJbJgEVwS2M65cC3FJMNK
4m9RwGRCW7MoFEgCEgmpWCF9/Hsb9gULgg6I/R4Xh8BrFcaAxLkdcofil54o
UuCIvmyo5N13Zvwb3OO7o3C7cNzaKaauQNwO0EkqLV9VD9D/Sufuo62ljUOJ
WLPtSyiEiqZ+QR01S6sjsP4aETQVlPzrtHQ3r37UYk9o/CNbErU1gxc864xM
gS9ciKr8epvzqfjxx/Sl38Ea1aVuZMzNTzzqqskgNXQk2JwJRiINSlToWJ8x
GP0nOENqNrDvpcOCn4aAF1ZYoAfHVT5P8K83e5SkMK0+9erzLnq+EbBhPvBp
PJGk3zAK/nDyh1SZ0OiWiM0gTXlnh17XhHBnL1ewP397i9sID2DlfmcAtPJh
EmCmtFORLIWa9MJIqD+geAvSQOsebE43KX4Gx+59L2OLrTVk1IKgAbZuGnSb
E7+ekZVCkOrpue3Df/gyFrbuO9TJkeS1BygxChsbnpMiK4EzoiRMOVEOnKE4
KyJuAHiF6Q/U90PbgGIONF5NbkHyEYZ83qEbQ7XCCm41kNHZrn5AzY7TTNCM
X2wUJl/OyFtzp7dzFNaRqBLoXKekAKqvvYcwxIuZKmT/qTKA9W1ojZu/WZgF
lNFCiOP6iwBbjuoB8/uJSSHrOXRdPvLUg4eP9Nc83AoKocVjcflu7HDGFwJ+
akwz4rjChiX6AJc3kqoZEJAW7RMaFhGInkj5QI/iJB/AjjwmYAKBGUmVQ/GK
AF5GIgJi3tchmQeeEjDCXiXniUcr1zD7EdBBBsjdm6v5Lw35TKe1E/mwWNgO
+xVII0ENinIR+vj0dielNvOTd7PAbdf1tGtcgP3LewuI6njaUWurWoXyvOgt
oYAqZwFyd5G+1xjwNNwqbDVJlQ07cE7QKkvU+3Cw27SAWOP0tanjC1Bc440b
qN6IWhWzkhTJ+f2NzPK1dSuTwf8J/OYdX8KBp2SzB0MhUGV3awRyjAjEDxL+
Zw0BzxTFdMUm58PoxaMJw0EXYWuALxLzy2byOhbmsMq/sncKyc9xxT8AMTX6
cAsJrex1JqHaq1tzoVGGxM1DcbFrmRoqz1zgAx6To5gg8kLRGqApOV/IbSu0
tq0rbYyXbdh5HdFxTHWIrAQMq+pCPEFsXSAfNbv3FI15iNTR7xW2Y4ai8JBL
LLX6OVoF0s2IoOnrWv1MwmcYx9iCh7Wa/jWzLWivA/riKK8umjxRYI+X9RB1
d8B1uZoKrYppAvGKLyVrQJfgD1gJW7SF1Cuq+9OPADXCZi1iCL0Qg9dCKSd0
EJLd+rkSZGdhd67xWOiA83XLg9DLKsF39oYoml4EvIylohyfMFRT3zgyVzbp
Czy0oKKx+xYsfqmBC9rjjan+NKTVhkKf+vwLGkvzdu+MDGrHpul1XVY5pCBp
tL50sK8pBzRiUswv/x3yNp9nyKoefSZ0kDwz3jtWOlPqjWaE5jjoO6vCYnIK
2ajndHMwV0D1NkRzZAbKI5pn+FdEgoyg6PJcDZVIY4zcMBVp5UCsr/zWDrX5
JS5K1ymoTETpEaEeIf7J7SiYpu/5FuC1YJ2dVsE1DYEqFL7JtMYlrUQKgt3Y
IvM7by79LE6yswL2euVN8ZIa81uWFl1sV3Yddq50zhnVUNG7uKYeRDvjTUbI
9KiqpYD5RRvPTqgygu85kaPs5CE0tPKhbGJzhOu48PlGTKItSekMri5afOp/
+E8CPMr35Wh9GjTMm5qPNfTTqblLPr+dbGtNmPH8h8IdYTiClPyjsRc/dU5Y
mZ4WRuQW4S5kYhiKYU9IAMV3lA968QmHFyubXoUuLRSuLM1kfg8IFP/MRwK2
vbhTC5wydeB2YKQMpNpUqOeF6kMKDsgYPk1VN/oxL8SsVJXSHVDhclsoh7PL
BU6PyuSRtHq0h31GYnX3Q5P9ueiixtsf30bZpk8KxMVZEWXFN87irbCSF6QU
Ymhmwy8FKwnurDA9GViMh9iCZbKVc/4NNeAyk3Kq4eJw6Gl9lZjuKA9zEC11
BRYpeHUJdw/aVU+CHABe3BnnlP5LQMxDvrwxsCrJoDs1mJSsq0GbO7I1/X9n
LzaPiovFUVHCVp7ON+pcfBFa3BANMcMbL57Oc8XrTrdL5dpR1d5vewxLBXx9
YcNLd5T2Qr+d+mKEWS1m+XfEH0UoU4ij6gENSH70zz9eRySMehEYh1XzoFhS
pluO/U4wYOml4VRTvueoew+YERfujobarDeDnmu/772el/vEwoQHMOW4im6A
pSSRjM5HWiGMX07tEudEikyn5rqhtPRD4TppppzQW7t6v1k8CVlXSQsNHIK3
Tg9HmC3ormnVPAYbnFguZFdX/oGACuE4eZXmjS76FbfrNiHRB+xhc4vD2zI8
ejm1B/dnDbh0fRD3fma/UKIq/L0wbvSgX/FD7yx/H6yCDkGjLOvOcB8Y+uNQ
XUTr8z+WgE62yzlzXtNAAczIVNDe7w8QOyyE4DDvs55cEtue3xPF+NQoDmHP
kTOCW/qHGxnFIwf7+eSKOJE9wiQiaH+XLegmiOGe8fhWiY9pM55+IkGf8AU9
AayThKvXF8VrooUSRG0+ZnT58wQrfsXgDiqD6Us4lMqEO9PBvWhBQOVjMzLs
ZtY+MVXuPSZx1ef/OIa0WMqlxOTiFW6cRLjrIYXtxAF20Kyl0KeooiDPK+GC
4XdpJzYBA3sfGc8eofLjdJa/BRYh+g9OwfnSTnDm6jh14qZK9lOcjZjw00ms
c1CXA/7P3lc+EHAEImLUVNTuuNybLz5JFiv5wB6OOk58uS6G2Hda9S49HiK1
FMvRsagK5A05lxp+t4fbYRB+iPLU3B5uXlmBqqWCT27adPqg3EeOoUZwVd8K
TfMxrFXY0veSzxkqTIdJIgcEf8emebuo7XPk+GPMGaPhNZO3vMNMgpmkA2Oq
Fzl5KHKaRyV+7iqlygJ3AZRXI1sEpVaYvpEF9FT+UTW/3UowzPD0x4dmoE34
xGNO0N6pXDFsIKG9+9oNywK/fLLJWeM+Nq5meXu76ziyRRPXqs3Epy0JxPvA
NbZxhVUMkSlkJLUx/J1FcmhIuQ+qEYC6heDRRnQWnRQxUVg8e7SLTfJtW9Fx
XDIbYa2XEXYe2pdZpBmLdvHYmclXG1rMzJyQkRE+wUFw2bOgNpYwC25HfVPP
k9mBueyFcA6NgoxeQ9rViE5dYdRfmeWlrvblUvLRHYUtmAa4fA7qi7swsBCj
+Su9mh6E2ES4RyGtHJ82u1yUIC0B2X5tV6MfaEtU9BZ/f46SfVy5uwYjoMCm
Ol4Gw6Amcr4CFNP8M0GRU+5BErGIteAbiwMV80io6k62lXInh+TnPBT6W/7F
3guO9HiU0LqgPA5IR8E7p+RP+l8xH5Yt+v4Z8zrx6KaBcz7C9KZIaEIkVAGE
yQobHHXvhuyw6Wjjp+bX9C7BX6t6YJIBzIT7MYS5yOtylGe6VuJl1ug4j9r7
mVphvn+6tCL+AypWYe6xvnUIFnUBh7gWwlfDIvimpUtdtR8sOmwcNfVoxnYO
0KIYgIxh5fdgPy2qTTVjDK7Awc9TzD10NOO/M5vzuvLcvWrCFWpm4HCbgw5Q
+w7g7SyGPN+BXxpcSGWjLdueKczKguH/3W8D7CkgTc+BIfK3Mcg1dvDKdGsF
ICYuJINLlNHdJ/9Sy0jHbgV6pRuYL9QqU+mCu7eVGnpedBEhk4sI6WO+6hJV
PloDd5eJlzUWWuE9K3y0ZTtlY6TuK7X6nHgONddmnscpdwRT+TmiVJ5Cq39H
3TSKdt4hI+oIIgAwp4iQPD9PZLXNwEuGSwtPei5MnzsVw8Jpigi1Oiifn7aM
E6YwSddbE6pjYnfDCq5EHOadNAcBYLcMFKUNUn+VFInPBS8fLLQ2GCk2kCxF
q9nViSNe/jbXkjQB0JWHCmwRpahP0V29sUiBvUfW2QHS5odc1UJ0jxTxixPe
gdP86nfeueo0JPwqAWzE4I9dSZAOukBz/23cJ0614czi3U6331GI42+0ncrw
s7i3gwVs05w7Vl8sc6OuPrpbcde+z6AmQjR7W1cm+e/GLP4fmhdx+2b0L6S0
R+g/BntvEWKmQsqKpNhOk6naWbkzLUGw9Bua4L2OBM3EKHFb6lWUqdzyLx9E
V0fbY0kTRE1XVFrwKT23Tbx7wfYA1tB5xrRaf6JjEjrUKkzHBXA5OEYibBfi
AsV+hnp7zCzDkaRe1jk0OmPjTUxwh4p9BBtWMgXSLrarYNGa2P1gS2/tmGkU
USffvNOlkyuuXkZN+sDcv09uBOnjBtBawTYcHn5O8s60cBvci7ez3+c6UwV4
IN76Rw5z+v5lYVl36Lg0GSHK9tleT7NZwpbg4Wx3BtqErkJ/q8SJEc4Wfa5s
r96WkK9mBGkyXbQ9FBKeN7N799jvAZ8RecdnKwtkdOTVt+b2EBt4vRyRWkPn
MiL6+Rrx+OYuDYjBVdAcSakDl8abc6bXiLFyGZcZ7DR13w4CxMlj7Ii9JpG5
o5NZ2Qo9elKyouDCDFnkOGw7zeFCaXgYLWpOBr7PT43sbqkt+SsgcoIhTMNJ
rz3PyCBQRC1FXhHN2VQhox9tVLkdHBa87HiQXGeHJgQQnkFhDKYbgRSO7TsT
p/tyLLoRdl7WqC2zbh9ZSRBgzvjOC/5D4q59MvUMRLl49V29qOgawyTXkbQQ
OyrYjWFCQnwVw9AVO5LPYlOmT+PA+LwjTSp2szEkmu0HihrGFAeR/OjxoeOL
II0nLlx3hym3r3N+Zd6Ze4R4NM+bpHk7Zytd6rYDHdkIiKk+1hkg+IgH5sQ5
CG5cUFr9dQGtghdiG1IFi7F1tzCx3eX4MrUFywRE3scJ4GcLjuz+jkGaT2sZ
GLPiOWPqDeFLFPvLxcsGVOk2gr924kTb6IDpTrd0XE17o/hwStQYg8dtpI5T
4uZON6Jtnco+FGy+EmPDgMHQjquJZat4ugDZ2n6AIbCff6wHbM/xDpqITUWr
o/noP1ofNuRYUFAVCcfgelG8PWMGgvriz6/04ECw9Yc5zjUFgMKt4uYwu0ay
50G7PMJGhR8dr9NrElJ0ZA5lOWfWJ78gOg5e59nWlsfe/q3rHZqxwuGBWAL5
bQIdRx3StCN+m+bNbGHwWnNw6Hg45Xvry8RpKVtFw4O4gO4OeKtj3GEsy8x8
AOeENf1O4Tz5zzFQkwQw5BjPVcbrxFhfUyVrDC86ke/5VzBbNoIWzbUhkIwI
xjH6O+cklS8feEhFPL+kqTEoQ+o1e9wq6h/sZF1U+Mt9aqrKe2JM15i+GKXn
+B+3M+GEfLTKxu/gTlxs0+B8VmL3GnrF4KZRn/A/Bfe76KJvluSpaJguqpEM
T0ht895sVhq6rDct/BFvLl9RftxZbSMvNxth9IEThdW1PZwuqtp+iklknY5i
6FM9amxncl6aQb7K+ZARX5fiXiuQeAYkd2pLu5E/rKNe+V4ZJ3GApRhiIXhv
05RdgmcBXdBXlSY/ZsPCCHaHS1csL3TgQ/wii0b/nnE9LI9ZaTsWFBxWpS2k
98ALKq+VScQDjFeL0bMvWQvGmymQNi6tGwQtS/0R+jNjC6/UT69e+3MeFbsG
XW31HYCyPvuDDM0q9kr0ZNAObIIysc5fBpvx43R3Md6sk33FjQCCt0jgvZLJ
KIs6JnIXuT2aP7l7vv66X/pi0FqfyQcc2yxlZIMNtcik3DeJNwMylIMVRMMP
FfkeoLKRjsH6dsK0KV/C8URyx4hiViHANspeI22gE+4zQgUAoTQPqF0Ysu7k
yLZcaY5O8mphNXRyMnQ1Gv/TQJldrybLANrN1L0a9HdLf0EEpFlkPGCYnpRy
BJIn6f3ajuwshhqZAuP9rptlJmmSEAvGvmVUzTVpOFM+4veeXcDQJaIQjNju
l4lSJMmcW4Se2lxNJxNe/1CqfzIv30HovBhJjKNQPCLaWG0XInoPkYTixEi8
S2cS7o4INjNWsCEgDy1Z+sptlsHDRrbQYKfh8etYAVlELVy3V4vSUTDKftZG
PKR5I9FR2x1JTrzoqQZRSwGbXlL+cNz6q/110nxo5xJ/A3fmYESxCTTn3vm2
oVwRq3KfnKfXdahlHmpjxM8GE/7aXu2M6u7H3w7KequJmxH/7ie6AF71756m
pkVIK4w2XqFz0WfXWP37tZcKbMaKOaJ+4qbPlYKSS7eAvO/AqfcPp+ZV3wYF
A2lmEHVQrqUpjkgGTjvboyW2go2CNCBXHLtVMUG0MpID4NI34/QDwH7JPMcD
4bpHLOV+LYWfL0mLoE4x3jvaxx67OU2EF82dbCOTnw+T/cJjsIT2vgQSdHJu
hiAglfZqZnyBGUabD6RhoQO4eiEWk3UcbUU8w43GHh6zsfMPu16TtDgPAxrJ
+835asyEGd7jZGDBMzvfsg/jWTpsBBPl/lEIvdpnED77QC5Y2imXSccue+/T
aHj1tbyUF+aWcrI6nsybXzFAqUSAJ1j2WCWlpvyYwPsnsUuX4SHigMQkCICG
ZHj72yLGjqCxcRYVttUWR8E5lnk5EkCLP5GCcHuViSntkaXLWX3ZrledyDXh
sUhudzwN9mYVwfjKBdMKxhmJtvIeNIJeuapLad1nTZi+JBHnKaa888RG1RK3
3V8Q9gRuUvXDWD0gIfkFXMA5Bx9WqccydM2xxoRoIz4q86/au15BuaQ4tAa5
0gxaNOj7WGbSVcAzWRrWP3yMANfcFW89ZtnxIz7VTfigbRFHWAnSaeZrDiHb
GVb+zHK+SLzOZrTl8523m5qRCWCvVzYSqHLhzv0bnLpUnfwFSsx6qvFjxF+p
7mq8e49WfECdafWy3BVZjH6dP7M8YpQBzMnFOpxJoCp2uWpOhSIbatqBsla9
X/09iJ8Ytp0Zmeommva6GnefLgfXMRqylFheNIDxJ5dRw68aILxxwu4RHPq+
6t4B05UVnL95rt0w+EAUGAq3wOwGfeLv+gbsDGsaF80I85pv7UAN/jMxzZ7g
oRaGonG1IZ3mdsT45vBpOvXqv0pZAHKhOjy9OjRbKItjsgjLRqoIjmEG44wr
HwlQnlGKImY0LnghZ9ICNPlcdlQZ1r57k7CIPmC3F/WFubkQYJx+9gX3UHT8
GvVIc8xx5JwyZfZZsKl9FsyKuzJwJ0TXSQKvpLflF7IumLxOtUC91+t8f1ys
WQ4ICSuXIcg496gTdWxl9GgXcISzj1i8jBZ1GdwA1qin2CALxaUTg/lQEPgD
QLqDsYtZ3YBmgO61TMututb7KRz5fDfSL3zgmtoUfjTPbaj0FNEjP+jNdJek
FkTo62PNa9LuvlY5Fpzpgws+hdEpqB1eORnbYungXnWXtPPfKJWF1aWEb6bt
z3s3Ccc0h1zTbOM1oqrZIE3f8ru0enO+1e6k+rWlqE+xsd/kYLpWzGWziNMe
AAjeSEd1FZWj/DVs5p6VFNidrFO0bW+rMnSlztBgyeNRFXFLVlyknXaieEWR
ENVythXS7dYANlgCIGhhhmHH0/M1Ie9wEeP6ppbdurghVJhQBgPNoN2XTvbu
o4OO40V6zDMBZJzCAhNvY9FDlne5MGXaXTrRL5DizsbfMznGbzt6iBRQzAPo
A8g6XohHyt3MpwtaVW3PjDSQ+7GTWI9Eb1SNu33tzo6Vd2BaOov7eNzUswb8
dtP9Li/CdW00iRepMNteCScF1mObrD3npbQ4KEsrKOxFkJcABldo66/2TMpr
D88j6He/Rv37Fwf2oEk0Qldw6jRhpw5Tudd+ivkC5juHC3+u3r81yiyhbvQk
fVhZ0/f3wT9QRe6CnWg6HXHg2+j43tFGAlBZx84lpDRkZ0D/9uXKxUp/V4Ai
K0LHGTuP0dJlTqb/xrO4kyIbPausm3j1AiSpMsdYm1YzL/U+KDC/vXBLY/k8
ygQq+5s3pyrqj0VLUohZHSMzg5JKyFNHB4osW8hH8HvyZjUXIh6h92GeRk/9
Da3jq/9uThfxypIYDD4Xks1EdfCCHdx1HaMwyLWqUtwP4q+XhwxDnsafFlCp
64fZiM+C7ueu5H2IdDEbeC8tjUcimO3lTvz/qOjCVAegpbI5AR2e3Y01fdLt
fzx+BRtHE/nx8uBAiphcw4vdoyqsJ8ZGMs5296OeEk0JXFCLSGrHkE3oqqfU
g30Nq6zq+WMbPy+rYMe/yNyR/jD/V5THnqFYiLaLcRUDpJ9HxRCHEJ/Nqdzi
3po1usJryrJRfMmGhvIRXZ42ImKQeAeeX85eEnRc23Uzco7Q0Ax9H0piACpf
6B4R9stnQVUpoiulDKrd/5K/6EhWMbNxIflTa1wTZKHCwK6G/R7GPifpg8Ay
Viu/O4m5b7GbW09f8ngI+22nRh1n76Um9dlIlMQf6PLgiuMrXpGPJAGPGWXX
LilfahnU4sIn1uiUbkoSOtg01xI7v4naUhZ+ZpzyEbEJW6QgUdwlLisvbFoJ
M/Cw2syqzbt8rS9aEm3JgcEUazuMrKqFo1g8cw6jMYh1xVajNcF10haLVKBf
vzhVKUxzLClsXL1USCSWDnnq4lB1hs3g3VZlTQk+ZTV8qesRwZWleMxfSS79
wNsdMTgSN6FhCH0165s8KlA/4+JY0JEafEDhR7xOgGMKheU04uJfk0Xz5rVU
Q9o4ETrIGcjTos8qWZg1wPySerIRX3cjh/hMH3b5lxQ2LLYPJjb+z+jbRsqN
kg5S70dGS2xctLQmYa7eHXcYxL6HjI2ioOhhxwYlte7YiD9pOwPQo3l3Jv9j
m6HE1vzUG+VQYl46KGQZKo5r474CUeKB/ZJJyQIi4WNTRqeygFVNpSU2qXuO
0muY1a5xZnDTN5qGVqKHWZWSHobEcPOYxP56oleJyw0MZwZOAbgZ8o8gZoTu
7Y7hwjyqc1ewzF/p0TeX83OO9eZmuc4S+bQffUQUZJ4XCFj+JOr2BEkaO5G4
p6aWjqYH38kO7UU/UcZq+g/I4TvUACAF7ceNv6+ySAiotPW9Ks8xZwrC+ndT
L9CB4t90wtDvY91yIIVEWaA87nFj12zRl8wuNcXmKaMrtJh0MyXznsDVAt8C
zjIydaGZ4aANJqJTBw5H4oof8yC5TFUQS4HiSqH7D5WsUPKTs1Qz1m/SeXFX
i/EglwgWWNCFzV1oIcIwQd2pUMwhlLfAFekZAHOUt7DnZlpWgn+5oZY4XyOS
dZ9HJfYIsF98Y7J804elVUushrHKJIjqdj5bPw5xUf/hwjYyt+/EMBPTkVAl
Q21yR4vyEpKdsPs8gE/5RSv3Z+2qEICJ8i3gVkO0ZQRp+yt8df5MhAUU3W/0
ieg6rkzk4ybtMHfZ8Z8jRiyFbPLAtokiL/q8rxp1F1KSccvKJBFEXD/uOZcc
c9EOBBTuPRWmMDhs33DfaVrm1Hpsbe/hY0KHlmaRjBi8SFacAk151yOY0mgk
c/XjGb1X50+vajLGYMzQmxm77KCxZzMcCOR8JnhIkr+UGE+jit8+jW+QIdHs
9QH+Yp/M6tT/uZu89MVJCfFD0iIeDiCVvQfthFEAmGz/V4Wzwmdqw/24m/jZ
70B3WuiuXZaylneybcQJcNQNHNVaylJ9QVY11/HSiejbBtYJPCWPJp3IwZw2
dBKGkzce6A2vcAblY/EzcFcIR3O48Cj/PCVI7NtsSpUP+eCcySxxBQ2G39Q3
1WFSkg0trVqAZ3AkooctjzeXsskJHKIl9wlWu0the96wyzF7PS4XLuXYCFHx
/bMZwc3UBHT0mmBnDI9M90adklrZ5pri6CnjcerZcwQnu5xWDMJ1/a7Y8lEJ
nedSdFAx4cKCPh6cTQODwP8vbMCWUM2NRG8Mv2Gv+ZlXe8k/RVS7KJo8F9Da
Hr7OLQ+3O46mBu0Fjk6e1L8dXizERZ+SOfZz1BvQIRQjdgZyuIQ19NAbqfrc
NhqGeQISV8Hw15OTCnpEZ2pHBzBjBEiiRd6M+XGJDDxXG5x07VR72QW0cUs5
Lteklfp+2PpPT/7+yq/9Z3Ihj79FHVO0Dvx7tjkWMiHhVy5BCuD5BlqFKf0W
IPHFlQBC5plgz3KpAsIfOXHZDdIopfPmQ2IPqcjcyofXyxgsEZWis30YFrmM
fKhxxtMChGB8jWp5GUZ+fmsOeocxFdQDnm7WqdntA1rWs54tEdF4dy9AV61z
ofid5GaZhnAF9iicbm2Fbq9IBmhU3Z+vLvAqG7QZmOVYqCeoxY99oq8zdm9S
NPkWJRuYlYUuIEpkkFjSaSdItxtp62fyp1N3VH2EW/dof38upPlDzL3klX6T
Onumu/cGTZfSz3kl0JpMcBSg7Q2q9CDAk4U4QZivMBRDwALFrZgaMclEIdKH
SqOgh038PGY+uKUWxfua3bqw5wkKqxrzf3pTojWW6k3089CcPyNpAyPnmOVz
iY612XqXGm4kSoTERGGtLi6sBQMdy3jiYE1n9qnfWDhrZy4+A3gOqwTOqxM5
bevRbeE/LR268tIm2BxYcNqdI79zRwCCdsU0MeN93EOyq9sqXLa3c7uDc7TS
JSj/AIMzEXLuRxbiSaYQTI2zBvy3e6aC/L7kQad0FOjGo4EbUoUyU5EFAXHH
Vp0j7mOHDhAVfjJ8C2WOUl5RzUcJTW8LKPi++DRjo6Ran8zWqBP+1fWHFwUi
JnNEBRXaX+ARVaascJLNbgm5MVed2GEUHzgfW5XQt305io71kUIj2bZYVAiY
8wQgZxTW8h6qJtVzv9BIh7/aUs9+ojadsjLflsaPqJ8f0lHVXsnBYMiiGTsq
YQrcAVAfc35M+59GYtQyzLsTZD+aQ3HpzmTiJJKF1VBGt5US+dpXORT58mkV
+dm+tOzgonyUQwM/pDPGqUNhM9MTKFyOKPdmJtkgRG+ia31uUGv2SyCjzB8m
QqCF7EkmamoO1CspvCucU0d6WzHrtI8keBeWUo9g/wXn81juSj8VPQWmzGwK
6RYX/zRTYUDQ4OU5jOajnsdED5ZE/2S95XQamTYSX1VU5hAPBzhA3A96M18C
mCPho2+xg96Qh2amgI3W5oQg8QDOpjtSvaU1ZuvICQRQG5mlfgNeZbVC/SkI
uIzeyL832T+8fipVTsU4RoEDd5EW8CAMC0kBtKyt+asnuTlYLjXdu4mlxeOS
CzXzBM/wREDYtupLpWmaMpkBfYKhLgmTScwUMVzwScJ7eEipUZ23qwyXIqeA
+A7b4bnBZfqS47mRhEhPoBsdecp6bvg6xVMyQPxr1SXd/Lczrlx7Hh2R/aCk
ihW1AKcmclA2+KwBJhqM5nxymiZFs21TT9xzSTHZ8Y2BqFouh+7G7kFrTo5E
UnUEQbKIBJdiEqLkPpye0kSnJxW5vibBHiPEFri/s35V6mZmdTzqBFUHmQCs
+DdyyzbGPtxo3ujQ8nyaZsEWZU1Ljabj2f8kiY6uZzV0oSfcOpbiiYORbN+b
wPsQ13/A//IVlwBd6Ts4+Amjf7GxQJl/5bymVb2AXfam/oR/LCoEoNYoEp1A
YBzEK/YvmPpTy3x0gcsCa+nLukeM1NLgHuQBSJwWCrBGbgEV+s/eW0qRVRlt
2WEWjO7fFSycoc3cEo4jMdGnyNS742S+k8iewMS3IzTc6F/TSuMbKKXjR08R
iUJNrNS4UTEV+lu34Bp1r/jlpwdqXnzpnVJXu3Y85iRwQizgThPNQOXzLG0F
DgQSQPNYQqHBI7r0sEzZjsgHPU4mUdrbfMEI0cZkzFRL+3J0WM0SazsuOMqr
9Xk3te6QZY8umwnikqVUfHiPHJvhcl5InbhzDnySvfD+wM6h+MX923v7e+m8
CXPid/bwykAa5+rXX0jADzsxadCewMTAk4vIYHYWhvkk7pMHPxpap7KybBaF
9B0709CqST15e55ZDKYp8TXUXJhQRWYCxdypMvD7jYJ7TYP81ZIkaREivjFm
mbYjO2k0dExvzEr2uZbXIAkWzvLL5kqawZXV2/TlTTx37Mnij5k+yYWd+xaX
jzMoY6N56X1Mbj8nXidx5HATUUtGDiVQdt9IwjnjvbNYT0AHbjct4IPa1Ut9
+B3ieQ0+ER5EnggzzUuSo5fsfXsEh42Qq4TvJsLX4fDd3qlu5HjWVodv8uMv
jnrUhVAP28Smml4jSxj5CrxTA52IeYq06D9cZuFGel1bTSoKLQ9FvLhJqcjN
Un0N7eNtOaN7uNwJKsHPHhWdM68tW0vGlvjfmYsyLYmSkIg7ghdM6+4L9YzU
ew9rRYmjNJhiEpfquIl8iqWNUDnTT+8h2F0PFvxMdiRYQbcXi9LE3C50FTop
jzbod2E+szxky3PVUUxuw8N8Ag4ILfCA3hLVV/iyxyDWEFYsCtGrY6B+Mijy
3nGqGAMoNe5LwdjQvL5xptkbgxUVXyVvBi0t8/T4YWuFKrKt7L6JsQhGmU+f
S5MFwl9HNjIYS6wmTX/Hm9Z9VFjykQy4BXeRGHPgDqr242tby/7k0Oy0TQkV
r3DSGDOYl0G5wY4Rhjw1Z13y6jftdjJPHEKwsQiLUtDbMP13sF32B3t3IUrO
1VUBZZf2TdPWuk0qoNx4j/PWb21bbupFv86On2bCsaGcqSfSDSjWVdHb58um
ZTChdkuPDrt3V2Xep8NQo/ex4567IUYYKkoLzfhi1ixI9OIQ+GegcBpI5VJF
uZG92bQSkKb6ZvPkiLCDISgSgU6UlY9bWCy8T/TSfGI8L53H/5n0ykP3CaPK
7RZqDzcn/jxHvy3e0a945SpJRhJrle21NcQ9CeI1ZL3MxeNP3bsO6yPAAqDA
I4amB+TOv6GGQchLu+6sNHMUf5MePmyTNWJZHcQ29dXBntzOf3x3mr4qwRLx
fdUuvoG+Kc68rAQXecbsoX6GQn7IW4wOb0QPk5FrQkFnGCphdg+tkeSuKw1D
mRrTbc08VSQiP1QHhiyvxFYCBjolIjGvc3pSu65KMcWYmnqtcz5Jh0NWL1TY
NaAO0eLGK2zJUP/csBCHQElDbn7McOk066agJ59Qr6kWM2pkoCLOUFwJVgTR
U6tv0wid4P1tQDIPbdumq/64FGn9JY8jnzgY+51xz1jUvDkxxWrf41mFqhju
piPew9OpzH0ogAKv1IgGZENCxROrdGdtmmv3WBZaBanb1KzqY5Hyzk5KgoIx
I7ntSu+rp7IhVAsnSgHq0ofZ02P1UyUaJ5/5PzQGKS9fRcuQG7Z3GP5n4Z8f
e+sN2j9OsnFdDuATe5qQXvwyQzQc2jJ54C7s3FQdbqdolj5COIulvj1XQ8SN
FuvDqV5HKDeti0XJsHdYoHDgSHl9FZac4ie0KhCC4k1S5DbE42MMm0ORBRw+
IeJ8qafswqGj1YMc1J9d3IZmpycpa07rM/tOZhAlmablB+Pml5k8w+GWzeVO
1+Sxqh91HeqIFfF8ADQlRpJQpWH6JkFKXbFg6BoVn5AP8xHMglQm/jqpXZ9l
CIlKJZ+1pn7W6RJ2trZlIOrSQXJolZfcG4+hK8fPBDONsHG3sKc6Dm86Ei0H
+l1+2rnZ9k9tWgsNZ6tK/7ahlv3+Ex9ilXhcB7/KARuey5pUh8DtNocgtgLm
9O5/9m9w2bKH/nHiqn6eWCKJdawHgheBp2WJGptP2MbUXUkeKJN4AcJY+vKd
shKQHhTlDFAksecsGhplYKt1XXni83wpktTE583t6Gja091GZ62Df1Ud6AuE
vB3xQGz1WmDZfH0qlMrz5QmwvqcFT0J8Y1fEeNcIlLGVhyAkKgZuNwNQtjBq
aRybHF2HxjyaGvqnkAkCK41PXf5n//lWx97HwkdXPIvtI77qpQ145BwsVBy3
ETXoIy1EDz59q9tHjyh2WL0AIrNamDllZfhkjwpZYiuXIYwqL/zoARynfxoO
E79jlQ5+87p6x3voce0kjcdCpAeABvACNMmhOIIQ4ZfmhqX6/8J75IurztV/
rt1LrOqZkzrXCGJgz38tHwi1VykrYLm6rpHgH/ra0qxQjBxM3rtsPsZRbrWL
5RlC0RD0IP3qmIiAqFRUxKYG1cULDHLOoehj4/sbBvdVI0MXg8wiYd3yW2p/
MNUvLWDLxUa8PiQH05hGKdE3GYGmCZlFJwNnRqO5gGurPHeckDUOCw2ExQN0
uj29Dd+/hrwD3I8bHarUzWU6u0pffh5STBV/N7rLjPGuMdg/EwGqTN7b2KP8
ythb4YT9a/5BN3cKvmz/VKTr02ZJQbqxj/9jvPGJjjl7VQmngjPfzctE8kD9
TZgcjuC0f43lqGChbUjY2inu5FRkXQYoxz4Eh32FpHjSkoAEt0ZRhk6ujkPx
vElioOoOtkPMfp9qbpv3GennFiOMGYYOrdaQnswSYCp2sdWyKN0wcFyeorcE
6psuYgghlOfQYWyv6ZmEAtNtxN5UieobUL3m88tZ1Ncf0VwKSSyQry3rS1fF
8nDHIsFkNprca9OaYQ5bYiksq/tRTsEPIBHakARZ9QYyVaRhRewDjpoPthP1
9Hh1CLlb4gQtDIuj+/I60NTCsNRnzBld4SiyTqldTPn6XXhgxxIiQwVm/f2w
JInQ1AxSDeUYGhBQEije87xMOBHo2L0ID3VYnhiBFpncEfMhRKoBj1XftTGK
RUrKySKXXoZ7Je45CVhdSgonho5LPEFN9IXRSDw2lR1E2nbekvt9FWDQMEE8
NQ08UzH5mEPr2xhoNMIIhIgGk64Fuc6BqK34A2kGh/zJoHzRcgiX5/LDnMZE
omNJEWPAXSCFwAmg+ehqgOsSzCAjGd337koGxNLfGP6O5OHvY4vP34KRLFKZ
hbypLUSUBkEQw7E9yLlEHLxHKiwnt5kDqXTcGW58GvWc2ilO3GXKUDYkrorg
4a+F4FBpgW6bgtqyGnHI5JJ6s6f2BpdLYwgK4znOYtC2SZkfnTO816p3vWql
kMNFsjmV9xX9NaUAzd04JawCD9YQhQOYSsbmuvqJVjsWZZIGzTVE8OyYs3Dg
RsHEjQbGtE/hu0v7QfbFnbC/I0WTaA8EgZWJUEvuuFFpANHxYHt+09689hqL
JJroEccE50D3D8hw4tpsLD1FFV7QY9zu1/Q1maGKV/5EmeA7Vl/hJG1p6yu8
NHWsjSTpdVMLk36gdD3claD2SSc82P6GSc0qR36Z+pCv8wgTzdiAvfy8Oo9W
53DPSuyEZdWn9eGRLIxRBtw3asVDQPoTNVrPrhR+qZiVD4i7nFP32q++CnWu
+CUTrRnT4pqWYR6hlnWKWVFKx3dZ5yYFJv7l2AfSnYteWf7e9cOThvUBglYn
6TluSsM5MOCQh46iX9ySj2UkRhMzh9SifUVDDeB60uInXYqSYodQPQb9S81Z
IplU7QfR7iUjcQjf+xaeA4tfctjcKUB5/rWC5YE0xjSAvWcXYmGBNWbyyAHP
co/apzWLbV1vY1N2VQn9MUwVPLfdU0zfi9XmhBFXnMuU/JYXNplYJXTNPCjI
s1rjsT5Q1knlSnEXwOHaw6mW2Zs8OAgkJDy7ILM2nVSb5mhoUkKjzo1KMlIa
XzhoznuXtYASs5XGxvtXXzQbQPvFwFdPjWrrWHvyuESEbNoAnLZsAKxhRzW2
MD3uo+vBdvTX88KlovU2cPsn6d8G3ZuHU8yJtNqKNBhGoGBfODiUweRCd12R
yOctYAUOdA5TnjmvqRecVP42e7C8/rjUhyvmczSFGtOBDaDXv/E1uEPdyL1X
ZEJAebFNsutsuOnur7y7VOJbXkNaz5B0fXp5YygI9PWXB+GSQkL2QxAm0/tb
xryyZMcahqsZnA3mcC0PYhGUFqg/qtR4b+/BZdMv0eGC0lTvSzvgZxHoSQUV
Hybs/ajWfMI/ByTmoLdzOJKHNak6lJjP0xNXpyTZqPGcU54a/94JJQiWrRSB
Plmmdmp9DO5XmbkGY3bmamWYjD435KhVxwggB4EK6CpvqMwO/2S3ilhlMuKf
hTEKQ+zIwCCjdx0q2iCL4IBlM7ZAAkTdcvX+HzJRB4B0RzLgVWACxsSnz4lV
YULDV7DEN2wpO2GgQdx5ffpHObNYB8/qk6l9OKhHTfK8tUfZ8HraHDQkOCmh
IDPk2Jb+qLvQzERBFhKD6M0HOrCxJNUnask6CO0U/tDHEL0BlyjIw7j6zok0
y6GzuL5xmLEWrUe9dmFWSyoQhp+pBm27DMkP5iNkIwAmsrdTCMjyUiPB7Xjw
Nj0dwgmKIXfczIbYSMOijLRhJqfrzh3Ke1o4ikDUQnUgupCOtJdQjvivHdUN
nqw3IP3W225u6625qf4gMb5Rxlpz1hj9ByLk6sRfCQZDOojw7AKwyMFXhjSf
dsv3WvpYyZ9F8maspE3cntKOpkjyqWEL2ImlEJVdblW2ROHDGI/5N7JMeYZg
g5osKiE6fnhJJStmokgo6k6ysfoVN2c4sglNImyafR/WhIQBeFYzdEq+hIdu
4ee9TlvKveINZzRuTTk0dh/pxrzFaE3jvPESm96uoy1edxR7HkFkgX71Y/lL
/elcC2T2qAWWFRuxSfC1qT/K/KTDQgdLeSibnbosOIL76psu3TcXtHR6nem3
kMY3s6UvXLH5KT+/KVK8+Du8zGSF5mHwcCZmvP/dMYBCAPB86otJ6SGQQgJc
EqabHmbELR2eww9Lo+O9zEuoq6VLYIowAI1lpOajJv1oLs7ekyiIRh5/P/xY
p8Om44on90oDviGtRbkcPv05j/rxgR616taoj77Sq261rUZtGZJblia3P1X+
sex69v5pKa6Lg3Aldm1reZMTw+6i0marv/hnZj2cQB+3cDSjA+o4K26BYMCE
/pYcWkGkTH9lSlSDx0UjB4YfTrZYtmd7MuY1bNWbCvRazE/AftaxCaxPhNql
wGZsjIbCALTjnfqrgIA0xhCsQA8hTbKjVIikUfq/WExzcYdF3PwdwWRvl4Yb
sfR7IxPwm1v0xalpjP7O8n1QwBhIYcLzW6101hNxF2q/znLngYwSnT7tXrQk
tVeu9ymWSVTbl5zPMG+GGKZItNDxYbSEbsSINQuDr6ZGOnLeAK1a9oV8RD7U
bU8jP24dBzOhqj5hT5gZxgEKf/oBGKJCzzFvOIujRpxubCdIKEdPtvGNumuk
GbishpILsGOHA8eANi/U4NYAn8ZcyvCQ0upb0RQLMkWA+cOooqcrUKUiXRJh
yrg1ohLflE9HCx9IrFoYxHHsSujViTn4q0OeBewl79z8lrV7jyPcCWh71NZ6
+9CP4JzIV6VVyZy038I8bERdR+Bbc9Z0HEMCCADtAZnEleDUpJYCxgABydZG
neEa/h1y5H+nPcSYfMceFK8OFM4Dh8/f/4DbBQcNZm8q17OrjGkSjpwzB0+4
yCOyDTv0SXVRVqq5adSFwmvpAXNPN3ITwVfi1PKbioyWoCJ+Fr/JLc8FJga4
FUL6nwdYgakxI+o9f2cSTU401v2rQ8EQ/3XkxagqqaJjmfT4yql3XiONde4P
keERHBiDCmVLYQAi9edb4HfUFHDI3MOSwbrGVjFK8EVl9wxhRC3Eb53Z80XX
DI1Bkupn/xqGmbTPL3fwZZqIUs0nxDvvfk/OkQdhgja4w00IbH/G2F5TQAr8
CD0t0CXgAHMdqewcELPxRH50btmM0zF5lTpCt4gLfJwlFtv39Pc76j0u/Ki7
l5px0UeO1wtUSgTsRWa5nQ2yzKyGA4Wyt1R9z1NpVChDftPyMSms3KYzrndj
to10/YJwL/ttdERfXHp8cLigocqW/DZXO5DLkuOI3MUc2OBbIgjRJXgedoHR
QiQVRWmhFoSK+HCb8KNKyGO0mEXEa37ac30WkB9a9VCzbSzWXghL5JfEULTA
QmOVLsE1IqjX09RIWmjxvlBPVA0r55CQFIAcvJmc7iQ0N/QafcH3rZ4SNWyL
rjFlDSundUQ+bv4/BD3GEk/AiiMfayTQDteLF8cOkCLw7qkv9ApQj3ijPoT9
w6Z8zEdjQXYJMVk5ptEd08qPol6el8958nulo5SA6HgumQjFpWdUUDlK9lVA
ibFPOa6PAUGWDw1tjBgiViigvp5JPVYo5JrL1USkEcbAHBpSaZv15gait3jc
6gPdrQr1JKHz6xG5CdWv+343g/We0poNNKark6sHf5CzbZj3bRdnsvF8p3uH
j5dzUzkkmG46c31XnAbnieVzBXABDddGSq3ifKTHa/KmEPcPJb/LNpeONFVD
rbHsTo3Vq8ZL9qf/2UfWthpp6WAw47UvfLdJSKdBvL1T7ewg45H3Vw+bLRSD
I4/JH9OwlDBZxiWJu2CtiCTHYWXDSoEuolV27B+dw24/N7B2MILIlSx5+2FK
MYor8GvPDcjMPUtjViQ1qX/AcyKvFyHp+gWtBHh2qMIZY1H/1gyyZ0++OsrI
HozZF3CWIOmja2qiA9bFkNi+ZBkcyHu/oCQ3Luy+SGWggK3mHffBrseTbPMJ
2GQnP7ID63f7X1GlC1TsaO6MtTEyEqVSuQtgDqkf6U0T+Uh+nXpsYQlW2w0P
O9z/6SrZvOBK9SFLkLIFHYyC4WJVEczpuEve0A5nkB0z7cm1IJK8SwY7gSwb
oOrVgkSV24i+0o/kk1rNzlvDZMr8dhQWxA4+l4F3Dk7btMHyAqHd+5ogeuee
rlTCEs6+/Hmm85bVUuJqxfeE0WBfMZUfgRAmKsWlemJ+N4eDB92ONTd7LdCZ
Y43z9x6tNgialFzaygGJ7ou2se0cVd6lBcJk/G5IjPEoEr+iUAGarxebZxEa
HfCzyWB6nlrAdPPd1eNAD2Rofztq7V8G1/nrXoVnkmnd9nhP7CyAB1sR4Tpz
AcsXRs/mG0OTNGIX4Ezw11hFhlOK0i4pFzEynwusTfRfU/HdhGlPEmj/vTMc
D7Ce194IgV9T2xxQ6ILj/G3fzzUiOIzl3/lX88++CAwHAL05mXoJX5Hu8saM
zqkbe6ZJJIPTyfdEpYO/cMHM8HZb9Uep5hEQgXGNZ94S/AvrDevMuynHAIgw
6tSeYgdoQrmN3dDn8Tg6WTyu1qT6VCxwF/OHRpSpgaA5yisRPuZHbWb41c3+
bCYUb1zs6Ey10P2+KoT3OgjNGtL5tQTP773yYzW1fECtmRpEwYm77dDKU2BG
SkCk5BSOAgOUZ2HuUPa8D/LO/IJ3tScLTqre5bRzfyJrVL0cd0+vJnkqGXmD
jEjp8bVCNr76kIQT9u4Zts316CgCaiqXPw7ZWBFJ/ScJPUBvy+fp56XdC4mJ
vgvDNzIj0soLiRlIKVdW7qDgwAjHTNDaeZbr83HVyRhHDAcOaq5PY5iSCizD
A+7mijAY6FbooPQ7M+iv/k9N5ZrJFx3rpND3YZYhEqEhOadVRo6A4mjKC9dc
jvQbnwv/m+LnVHmC5uiHFMaz1CCnUaw8ERnOar4CgMjiVh/iYY/+9wf9CgXG
3GpLYI0pF5baiYQRXRa/0nXcqLhLTYTglwvgtltjtv0nyZh4I+OTUjH918Zc
WKkR+gU3B9j03aU+DrQzumvviAr3oX7d0AywTHSEZkutB1HV7621an+6e2cw
lex0YHizRHDzp5FIHDiBFIexzhTqeHpGfWjTDE8eM3WMv+yUuYWfpFw07Rnl
6+04b+3dAvTlG2xSwSy+wUBNcs05X++vIodsvYck0ZqAgVwevqo0XDPiwPNE
zl6+yniLfomEKVajdTBz10Uw7RRePWolSUKUm6LSjg+MR8ZE7wuHCcG0oDfm
L+cBhVa7A/pctEFduq5ZoQgjfOKFd9Z0/iI0HC8kEqdJJth9Zh9+X+S71PdS
VAzRBFVRSBahgv/YFiHiQgwfQBUMUo+gZ8psZ0CjnM2oNRQzK8LLu74fpkqI
Dp5qjL1G4A93NZLd+O9MXSSdHCx2IaadOPiuoEVZik0t20ZLzLAUyfyWevUR
Ipa9vMFNN/COAEfQW2vZldYccAuXPeEjG+vltOZjH9NERBswqkgjsZp3h3WY
eNQeWWluPuVxelKYhBkrsHhYS/EAxYm/PW1B2/HFfVBF0Itz83JrAV+vXXgB
VfRHBE++WFiTPfdMBlFiRzZ2Om424UiTAjy4KQZIbYAAiD8ttIx6Xe9RW82t
A49ktkZfxaRLPxaqtQsjfplEt6uqOZgBDfalQPASw524q+H+zj6t/ByEgVif
3RmZwq8vrQDHfdg99EbjHKxjBkGJ2LdwlCoFuSCXj4Z6EUbry7h5C0lhd7xg
CO7GpCg48IT1cr6PbSXmiXxhv9lyyCiDcd4GyD9gCEYJKx08eVNA1DHkAUP1
ASSM/i2/0RZnxEtdoC9kddQ2MEOLErX9TH78jQsH4VwM0cfY+MPbXc45ucp9
cQueJ7p0x88+IoVYitIFDDU1LBodsRNCarT/WcoWKoVcOdRxXFvxPmm/zE+P
S5ILv/58iRU6CA5VFPkmG/ljk1C1Fwkc8WYGKjP7FIOKTRr4YUDNfpmy7CYm
NudUPM91CHk791bF3prvrCenZBeTd8cXk30CR1vJ5g+XuhKND+0ELT3wG2oR
S/Wke2VK/sM60CXQ8/Kq+pH5U6wePWA2keD0dVN623rpgJqZecoBFp3N6uPB
GABOreRioMgxwqZrSp8y3dt0T+qK52SxK0MEWY7I4FMZTGbSoqJLvgKkB9af
25xxcd2wA4xtDt+mB+PL6QzSvZRBpDp4J/PHCmlNtM5XOmqw0ign0+D31S4G
ZQ/EBP4/D1Q2vgMnASP8dnkeObT+p+WltgXeBckMgSyQKK64Y0qBRD6YUAR2
7Jej1klqp8Fv4YicpYIhNnB8NvjwY354xwQzzet9PzfD+7EBtW2edfh9PTDj
luB3fBiQBd+9tQCGIiTfjr8oYltHfYLXxxiLFib3gFsVt1VIHIg03KVowKOB
EyWaWrfZzesq77NGiw/5/kiL4qHfpxyuQJeS2zN/7IfuqZ8PUf9MXbdgJPDz
0qMvGhpdyrsY1IOSEQfXMXHO3F5ZEsD3O6jC12IWIthALHFS6kn7Vt0TpYsq
XEj5WHpCdifL4AROCV7xCLLtczqGhWoK82s9OkBJ+HfltrXJvT71p2z400g+
NILXRT2nkO9a9LBXfNXsCTOWqDAZMG8vBRb0KAY3y49tR6Zcv+HoWtUFytyD
GeZulIt++wSSRONvyklt3ZKfYEMMwVHyxowpOIwYu1Mr/eHEQOHKMNu7mBqv
b8NwoAmC2WNPk4Ma1Lhw4K2ZVfi5FEXs8b47B/5AeAmI9tHZ5U4kHzb6FQRh
KmGaM7Dl9f36dDRdytaXUBPlco5Iogjv77kOq65HE9kgokeBwqnDGnuS+JHo
RdhC1Y4Gs02wTXb0o5naTqvJSR9hfkIFdtrnrpiMilugR23iKk1VLMdApNrL
CipfQLS3d2H4ws9ltVHM1oQBhs6LcbJoRtQxJe33waU11sHCq1eeTX63AMYR
GXzfOJvIbTgppyMtXszweH5WVN0BzY/DgUUfgL+bRXKEXHGHBcJYOJ5+bIqC
AcupR2/RY4o1cMZJclkl57gkPh0G/zkzmou3y6jnWYSYz75MC1WcPg2LusXx
GyaX+TNQU+WHKvKy8yUNZEPichaqjG0k+AxgLPlQjL0i15zcgFQG48kniEmI
uCG3RCWpnlFlPn6Qs1mrlMqVNQkx6D+rD9af5mI5E6zXWLFB0j8flJ8iLwMR
WxkkR1RhOb6BKGnCzNSu/n1XrXXe0dKGvRIViHjqmWXTUU4pDoZyRfbCesA/
CW0C3YMW0i5K2XuQv2Lae+ijTM4oik7wZ8lEknCt5RLR97PP97qeBE7DQSnn
XSV+4uYscWJ4CxFmAByjAd2L8K4VomeepnTUI8EW2uUrYucSVIdArMXYJnxS
xOBh3LnOgVMk4WWJO7zy2a87VAlSKa7Dkn3L4u5qa+kkV0TNmCITY6Vi0SCl
hwSc0yS9mNbHmBCY27DCIUkNA7tjKFBrmusg1ijVGKawFKyz3Bh72/EFR9Ld
fUNDJ7kzLDplmoC55AvfvkERCIEbLvJ5JPt8IM/tK9C6UMxXdQYoHUH91gdA
YUOITI/MlzMW5C7+AakGvVLpzuboEXP0VUgvKhYWCni8QecDCXYP95ofNWeJ
c8ECUdSQVejepwjitziXFs5V7fPhttDjH1nXjhrOusJEpxIbrOkN74kA+gUm
pzpKGZu7GVU8HNFTvoIfsdbfwGX6KVkaPDyc+d8KRQMOogsAR7cRDDMYxTwf
g12tdUd9DotVPldTq3IXxNj3qr2g1593tqx/fFev+H9e/rr77GM7wCqZw3HF
tozjjQN/e+XdZJawJJZm5JwTQvMXW8bjGepIFqztixvWlczWpuDGydkshOZa
4ZCmFCtG+VcDLYk95RJILtklmb08OqHbt0LK27njcAzCw/YcIsh5pQDk7RwS
IlqZLCNzPq75NwkXLnc0bqTFv0r73Ilwb/gSzZmCgUXp8jARz3Le28U9PCr+
iChzVFB4xxs/ktwqHmEnYivw2X6L8Un2ZkiwQlDDPX5Mz5+Rr/fIxv0U0S/l
XxfZrUQdxHZwJLLV2+93o8pFdBKVy45S2Dn+l3Fq2Fzt/UNpNya7lMlRJKtk
ciYPpgccJlkTsNjvX1m5flqJ0mRXGwE2J8zWkkK4493NbxMcqbe6nM5oMXaZ
IhpUwj2r0EDrmKTLvnzP00JM6eB19PVzysy70RwkA5YY+S0rzZmZ3m3TdNee
XrWY+Ol+BwctIa7tVk8p5HUCTwzsiEjp7y/AM6uxIHBjRH53JEy22HCWGOVv
9wrqwOLFXU7uCqkEHFxRyHOFP1dl2r0pLTAnQsfLVCPGtzPuZggsr6jz1f3B
rAJE0gnTK8dIkhNqa/hylkWAsOzqjPu5v/eZe7VVinmbiCOuZdDj7mG7ZY8Z
eGfx+7qjy0x/NoFb59EqDzdl9l2Ih6BU9HROwodTVBfGmXIWCJBED1FeHVGE
M4uTsqQf5FnmSF6JdwnZLXmAePTuP7dbAp6qNimokhO6aZKh4i6yxsWLmSju
XqMvA+IJvxMUfVO0qiht0FL9URQe+H/w0OofoN70HneTDf0eraRG8JJXz4jt
BoEmTARjF2ZXMdwoVfPPsKdRujhPYX84GExHIu3LfexRMPPOk/1pB9URXi+G
5rFXtzcFXirZhxwuLF4vWUYLWedJZuIkJdtOXu3ZCDBx5DsfRLHbsnDke0tP
R9mwTPXx6xwGryQPC3dmN3LtF6cHbnvBwEqDi9PM8RihQA/8ON7pLWsgiBNj
K2abuZ1U9zsp7jg/c3oIJh9e31qKNMPYnndYD2JgTZTceNpNRdI/Yvor2sHv
g3H1idJ9toSC5ib5ilMVs0EdB7tc/qI6Xcyye1EYfsr+Epk4G5wDaaaJiplQ
9/5XJovGehwigYKJw6bHV4nGJxEb61k8yLzVb9LAZ7xGC10EQrBUQLV4uQhJ
JKmTx33SO1dD9HDlNKqGM1Vi0xfj8l36bKQoGz8rHfmtDq5jKle2W4r+LxFh
DF4wkJMdyrDH9KqoYwLdY7QILJa9mdpIG3ulYsRaLpHRm2auwpg+xbp/eOks
XDrR75hHyYfkr1C1w9F9UUpcvMnEU+eqPjxBHrUqIzxkeo3sEXStZdVh32fF
FyXKOuX/R6UtLEap8/IoaMScOHZose0HdOXdyImsUsy32lyF8RhzESbfU/Tu
zIUymnvB+PEOyOGT6/O8d7yYWk3VDEbZ3bXdLlRaPFu9Xru0Ct/bRl7YSmS8
numGbLi6xcP1NkDwwWRIHWQMud2YeTTqVj/7GkUbCkGTZMPU71XxpkexYxQ7
S9Ldd2Juv8+oBN0OgkIbpKUY1pojIg4mp2i6CE1yWQ/JDgIMxFTX4RGG4A2t
ml8tsSCNCx8S4AmoJvMmH6zjwBE02+4WrOs8f79lrKbXdoCYCPyp4fKzyIYB
jKlEdeJVre+gMge7Fj6ahrsyc8Xi20bjyb85mIyUcLE+dCXXQLJ/XSyInBuU
f/xZrg2G+bDlB+q46ggJGU83yy5vxDJPsN5AmaHu8A0QGdm7qFIwm6Ph4ofW
R/U+nPlku2kZjVwQgBjOXilxPDoCaAXQajncYKPXpzzEQL/FwNqs0ofXqBFw
z9VJPS2ivrXDQwlsvfppBujjEVr3018Ikim4cU5Cab7DwH7V+cMHyfaSrBj/
H8lKbDouqOoJ/r69F0IJ+K0QMeDUJwfZZAAwDj9MopwaM3If+b5BF1XfVzCR
8GCtB2eNFshSaNURclXA4CfB1yyGoGyz6x7x1aYFQ6KbO3QqjB8Ce/YZRxse
B1LIUyij6gSBDjKP4P5ftfh0ehRwRHVcbqbyd1T016CDKhHzytlzLJgVQQ/r
bqmv7gUoEPWzlIOs10OWk15hjO9abjCS7xu/MIs8SN6rs300RrMTVjKsr3QV
55Ut0leMpw5ypyH827XW5QlJ4RTh9XWQMr64u69gqUnx+yeJqjXeqhfm4kYY
qyDjJO+TzIITku/WBr5cVCqnjX9T9qIMNehWwcsJOoKlpe/i14B+dJbiY3H+
/NPHXTo/4ReGBhEjkwre+bt8IMLkFTQ2w2DseMPOiwkcGKLqY7PXWhn7ff9U
1BrjtoSZ9fiSEg+T7sSbEXqGOYfyqxkTZeXyErns4CS7Uzamw6/whEDtwFyG
a+xco77UhOq3IbRHM5ShLdj5TZbdgDVBs5a7Tdc841Mp+b2EJRJEm50dJ7XU
FuiJYfd5PPqddLGyO02Bp9flLcMOUwwbz1mzAgCDAOECzcmatBPdbA5ySXF3
Mcn3KOiPgTHIVUk3RGPgYgBBg8ceCgBJlgP9cX25M2beVrTeFx2p+yRYzW0J
rrmcOrwP+u2719kUxhN6nVNMyCwThTPXr6gx+2uAHqMLIE0mcrELo+WBMAng
kmUEWKIBWFqshW9PLiUhuJsqmE/EjMHv9GkstKJdjoR7xCBKVlEn74Gl1PBR
R7RXqQFj4zYak4Lo9EZAfjpAcAAMz6FmtkSg10rNVexLS0vtymneYmsLZMLk
zjigJ38dcoHILd7xvFIf4ekXss/aTH9+am9ktXHkKoWcHKH6tojQtrMQTCD+
HtiFH1JcUl2AChQPqcxf4LdD2KMr/jnvjytxJni1qBo2yGd1OlMJaPjG0J1n
V/G0s+VWlNYbIbt4v58ykhfOGWxjYS3cByRDqYi31+bgIX0teBYciY7UjIgm
2uIK44rZOGF9mBQ9wxWv+6+5nBVvewyFY/Zoya2oeafHOF3Md0LVYytWbGHb
QRkW2YK6YRxB/DXsRFPlbZ1oRnuv0hG1T8mqNd2DsLE3nAxVwLEPy0IJSjdl
9QYEBnho1bFDm11zMfYY+5OV6YvQPFLsj3poaN6F+cDokCPA8qv+lMCuXjVk
mwO6cUQAnH7fHbi3chF6ZmguX3NfefuTBNCjmcvZ78qkCaf7m9pCesFd17dS
SN7xvlP+9h/n0edAtsmqY82nuVc53y4F0Vxh5+AXbOgRHokciqM+d/Cus2JM
ZTbbRkU7+F2OIP4JyyNw4wnyU7xTzUMJKxL/hVSpmrWt1RDmVAp83s5WakR1
FOj+YzJ3Ni6zaQOu4xPHJRygWCvpZzO0BxX6C2/dkC3DxAxMSAh9Y708Pqey
OKeYOel0o39U2VK2uWOYdNehKETlbSt1pNo7wezAPejzfz7Bf4wZve1lStpe
EsX/uMen0LMnNL4zYDUIfl3q34Ri5aQZmPQnaJj1fj/uHw2XMlsm735AXdjf
9v4g4dQ+ngu6OnnDPF/dO2v4aSLWFOl95pmyxYBhUBO5K51UlrvxGs4hdYUJ
webKWyXDpT/QdkaRh2an6PAhihMjnTOci1PYXfY+hTn2XKdtyOaYEvbvOa5Q
F3/7AZtiN8SdDyPJjQijefG6GkbxNA8WZlZV3UHg3a6CKZUNQ2Kio7Tx+6kH
lzCFOmiWryEYzZKFDGEyX+vLCa6NqOEQlh62MTd0qYJTatE5rLV1qW7kX6T8
cwpO4n+1nMcRY3zf9aczQAHdrk1dORKKIq+dtXU0ZJsKz4YOmKqV4Qvq1EYL
nUxTze2WBDSv+ZQI7i3bKabc9yP9fVJkJPQmJwx+N4yPp+9SS1HXTLmPfU0a
n11dLQQH74YMPIS0+KQ3DZUr8s/xUq602VxTt3I/qkPjcK5eQ9Lb634QFIYL
CMROaujKUFv4Vof6AeTArQjJ8k1YUFOWeU8GETRgvJhUAlfDIYd+HBlvfwzq
qbAIyAbtiRFRIENCwh202whqasmbCHlyySU8xi3ZkOn2RRA7iOTLyEOL8EWf
QeJAlT7KdMf264S0GGVgHu7ZpWI+XECmn7HNSB45ljod5b9pDT+z9mu8JVNl
tpqTMQr2lk6cwWTogjTvSlsar+SrF8YbKh69SRAQDtNYFItskvPgqgZ4lZkY
6czx6bHdFKxyHscXj6JHTGWzbMn/U9rI5N7/+7ZFeoALKOPFI9zL9liLgg1V
GAhfrnqhncnIwxALg6HV7xFfUKy8wWstgvP+6RgGnTCYjFOI/oNruD8cMy5U
/z60g1rFBO/eJ2ewFUDGo8BvznPGugHhCIZSBtIWkfprN7tDK9tdj1Vk0q5Q
ubL5Mnu20HBKVOKP+2uzH8p6jBnUpyGQnI1GK8ZzPS5HNfy+4bbvsr6qHERE
wuiJsRJhje0ljJ8ipo7JNv1LWJ48YqnexdtYBgLBl6ec/bTe+0UPxbN8iCVF
2oW2/nn6SM/PLP146hTlpy+3mcKVasAzTOtlt95PmB1lzHVSx+wwe2VnazSs
Nvs/mrLC8g7oXdqRn116JLZAdIjRaKMyy4W8QBy89q3OGUe2KhjcOlKx5VSD
6yvLG3dcj8AE041heQv6Sy0VYpNqY/Bdhq7sEpFCbKlcKDqwrP8n/zYAxJTE
cZx1bJQw6VwjcVu4FAcrvtE492iMhGU4UNy+PEU2xrxoi7Dw11xj8YxCH+/u
04kZU3kfjJTvs9sOHa9KKAHXJKDhSbumwKKYMBZWk+q+SdwHVCkwZ8hmU+gV
usmNd55IvK1G6mmlHuBI0jmtmkhgBCyxKOUMfsE9kcl1rem4H29a/Vv8LsH7
5h3UQJFPQKBUSl01ERyUJyJsUcjdf+jHC60b7oW6jjNqbMvpcEiiohnQUTIk
f+DpJVvbfvxMm4k6iyG62k1nnLWFOSVrVeXpuzCfzPLimW344+nrZmCmjTi9
JVl0qdLr11thIckCwGynFTLYmSfIfxxEjAlxd6ZqREPXtFCWdQMxdruM+fNE
SGWyxrEiTr6h61FJGE7uvHXcSpXNAu5kj9F/gh5kWN2XicxQ0PiF6wvScjBE
Ve5edTXbxiYnUMKkQ99GnOymnqzs5lUhGMU2l2GYuqRb57kzTXebRG0yZln2
27EJqVMtEduIaB+YBuqXp8ZHARRkA/Y3rk2u8grJ4n9G8JDXShLoVAQYEeQ6
dJzTegplGC+9jgNwm7G5ZBlssOL/UStrjjIWc+4eOwjSmnIEIU1lU5u2+rF5
2tIESL01Py9dT7Hyb/hcETwSBquddIsD7TMFZ+xKbTViyAfScwfMNuiFclj6
9QsQZex6MD4Q0x36UWfuXJBheyRqZX6FLFANcZffXGiald/MRFmjiBbIrtwv
qfPdLxnrrFu+kVrpVwgdnoM/3RAdBNMY0KVgsckvrLt4xjl3jzaOYSYjEEFZ
/QW9zpuc6XZ1FHQAv6B4ueZHz3TUAvROwbemlySpDjH0VEDLNOthhQGUIn6z
m4oEtS/L6pGDG+WAeO7+2dlXbIGykwIi+s6V8Fauid/pe4NCKvJA0zQ4xnLq
ftRYXQbwQQFTpbbRTBIiA0Pop1oHHIpYef9cLKzHiiYOEMNkgPDhyMGIbnW7
GCmW4AmENdfITy11Gazf4o/9c+ELLAhV145z3CLejGyZrvzvbDB1J1EGuCIi
IZn/SBEued5ogbNTFhI4rqLXn8un3yuMe/FvCREpSr0oNOTbQtRLdHmLrN1u
gZqoC8HWjYeYZ7KgaYmvbrZuTfi3qLD5XusyBFraQPrO3cAli5Mgi2bMtspw
6MzISlnzTjpPbzJBgnY8B4kfyujF1VXDKjGD417+TmKkhinZmzu9unx6xb11
yiPkN2CQWsiFTuf4us7inMsTaRqMjKeksawH8d6c0Dw2os4CPgodEmWrFh2z
8NVz/K1UP6eyDhUE5osImrEJ+g75VnxG3B5LKUe41Ho/0Z+CWR9+7EgzA83b
L/Uk7ixjty1d2ZP+0LB+Zr9jMTFm+LKGBVONT+dGfG/D+hWz6qGBCpdoCQJ/
KzlnNXL4adMIwKLZwG8MPPYVBgqgFspwwwR1qVHzNnjITqbBnPKXvdXOzvO0
Sj3bgdKdYbqQQmZ8jaeXsKDynfSqI1ns7l7nHgyuF5AjKMjfpBtUwl3IhGt0
nAODxtfzrejWrEcRVsfrikHInNBuSyasAr35FA1HBvDPCm2Ty63sYEwpVK+E
+7Hug/RgmacG78rporvKguWfi0c+knpHmysAwZaFxQ70NaDqFaEzd5KAVmip
OskCjvqdmWoKyT0wBnWROgSWgxpSC8cFzN37eXRdCHJStGwVNiCS4EcWO8Eq
lPHkr3n/Z3n6VCT/EXJkV4ApFwq5WatNGsX+irJv+t+JPgV8Hf2RdjKguGAU
kaihKdv2n0ln115Tyc7DSVTa+tdV08DEF7L/ufbxk99hCCuJuS0Tsp+KExuE
md/ddtGPRjiqt0FbWdetCeLQ58MpdyGhfBSqoGERu3dIo9YDoMROsXAg314l
XSRzBf2EhITyTeNuR7p9hbSFKfM5WYK5ygyKQUnqYKlO5Mi+bXx8zS2W1RSR
RkL4uwVwDsQju86M/Y7Iop7MJbWvp5T/nRsj/CCKlT8WpPIYY99h+9mQy/FJ
2O5NHXkXp2cMLaa/RIUGdiV46dJZ02Yoaf8Xz7tRm//sgf7zL4h6sMRIm8gx
YaD7jyA/TkrPfPk629+1gTWneamASqOWx68dHD3MJ/0iDGDbFRXc7+L5/d1Y
UICtsmaV09OCX57fdSf7XQGKs9cZ1yJCDhZbT9S8h47I/EbVyqduylQJhS+G
MKwzqJySfMdLzyrXM3OACg8neludvzKMbHpjpsDcBdAfmVNPacFKyts8g9XN
RaFLttUi36oYHCW6LFZbMo7C5YD8o6SktScr2MoiWeeu2jXW/VMNI3g6jQCx
Bavi6hum1QoMnzp6v8WXb2cJwF7D69mrQTllaZ5Mcri1AA0fQaQK3zQ52Qlc
1fgGwD0eQvLCkQi1oa5YlygLxzUVFyt8/ZnG3LPFllBGcni7jSam5trQaWba
TS8ZhxexkZ96QvFs2ZvheiAo+mxqBR8Cwwg4UK+LGflrhPEsoNeqWGwAxFQm
bcK4P4Q7sfRTgq9w7iG+CSzpMty7/x+vjAK1i91IDNZq9bU+ywL96VSSeoPB
6e4oMCNjtaqAgmrBahhzERQvdoPKwRzy02lVSmsDD6TQTtEiKkAVqxmojmwt
2G/ant9KUhfcHeviV9gdwfY/0TLKbD0gmIUHj6wTU3bv8FGU2aaS5CQhxS2+
XCuEHcwwmqiOLiuRpYZe2u3N2lNNPMBlRcTdP0gAu238x+zn8lrX+/EIVlsZ
1c6ueptb5KFsd5v5XmUN6L+li7R0yWQ9S3rLOy/mkRrh2H08fFlHUgcbqu7E
gxeor0zeiESnOnM8PXTnvMN0jV5lLTE2rTmX8eITSEjZpMlYTamvLiTgo9At
39XUcIFsXNXd7EGdEJHiB6x3eioTVhULoprYq8s19VuzExHW6vmdyWmtU14J
c1AZCPjio4Nt74OF5nGC4jMyQCkAe/EvIZ+2OicnGXhS8lFnZX0oGun3Ac4q
0Anpw7Y3y1rkWEacH6pG2mWeIEtEgbM1shTT5JqREDgIoBV9ASt2S9wH/z/V
wUold8cB4UurpZ7fWg0Y4ljjzePfCPC2VlhFw9KCJ7PBZOZTEUfEChB8d1PX
Z41toeH0tXiS6kd6fkPaUuIBuq4gJEHaa+fX1nZncnEiPJ82l1WoNW1FKMrE
wr22DT1daRVJLXIWw2aY5ZIImkBJKQUwwV2n/euOxJP+4X+zErx13wxMXcxf
jvLrQtqB2wTRhRsxvRw9QDLT8NPE115NcSoTDe6Vm3c6aHwrtL3M9/sPJZxV
Fwcep1csnCzmF+V8S4ROrodiNXQcDYaVHK3EVwkqOETo/3DCAK2VOzaTKbH6
SlYtggQhNkwulZSNmPTVQgUwWaVivw+6mI6hNsWT53H0S2Ahkpl1I6I3XFmr
jvudN4UBvXyt9jKYm9Mkl6w91KJAQplZDjy6i9oMQ+gdrrX2AWHY4V7w8SXf
iy/6rJgLCfTKfHIIwI4UntP+txmLQVd19n/u7jm6gIkWDCaH6GQJIBvvCRF/
P6xHZBdUH8OCWDAG4s97aknCYT+SdwEBTo993BnqYmdmGRkztMiau0hzRH+j
yoxRoRx+4Ex5Kbl45jqwZYOTRRcdSAgMtETtK5C3mXeNpnoHm//tAa4jr1j3
mPN+VqPGAqhrpPK1fsAtgF8ivlIHNYWMWCfk6wb5H9eUs7PSR6S6i4HONiY3
zpfkSFj9Qx+gmLk+lwH7qkY6rwPpDqP1VuN7pwPX0Q6Vb6eAnWQSBZlM3c2K
Y0JmoAccAVHgp7eoffns49ryRmL5QXVjJZiiL7/dgHWYTv3Fk5O+KEJvHPN2
J5fWN9Y//qysEKOcrUeGMZoxcDla26o684vjdHt0tW8gYiOl/4oyVksEcH4u
8g79JOAJn/CnGKAaI/4OUz3CUe6y6308MjIRqIKzshL9uA6am02az6YGC4vw
sXfgGd7RTLiPo+ZCpCXBEq3Qz/YrOeeAaO0bb+KA1R2yfsHWHtad7izyssup
rBlhzlIIZJ95ubjwS/0xfsERtFSbpScq7cTu8y4lwISr5PG2SClYOj2SsMge
Kpuhqnm5657NnMDO2HgCh/f6awTlTLpgDE2jnyavEOvH04v8R2ByMfEr233N
pb99DwQQzL5VJXGjZ2Ve4hJY7aWCShQUnRFptMTaU3cnF5sB1S5PU42DumVo
pH7ubmlkO+IxpnrAh03hsWcUENziL+yR/RXyhs3tYcGvwPMNATaBPrtFks0y
+hOeBLyxCiBJqd7HGC/WjlENgx0B0HtWW3Jrs8+iecBAR+u7dceXUtXjYFk7
NN/COfb2c93t2kMHt/RpUq69Lo4ndzYd/+hs2+4AuuhcFJAFGIbpKcG1UHR0
TN/2bKg6nu+oyufmqIjfMGxsZG6C0urJYrd5b0f6hQ7LrF8Zgx6y8jhVgia8
ZyHJ6JxVlhobb2k4pgvBjwxBla0pZixd/DTI5B4cTZJWPJ+EFfunDi8yc1Zt
RTgqPBqR6S5lf4tgh729sNA2NRW+LFtxymqbzMY/FCaeqVefT32AO82Zty6G
nkYAZ7AZi2+jXxpwiXdx9k/YQtn4bqEMBgU7wQRXy6Xj90mX4iBpaFyQxykI
IoEWtMTNk3Zu0JFbiEPIoyzf33CAVF08x14xCVdc5HtndHwuoOYWfBwkqD+g
eXTDvYHxXxOK01qePvRUgQieV0IFJ0KrHoo8GrgsTyBSwQ4JsYx0TjrpPSlA
hhKl49GYASI/bLopQujAR6+wnCQLPDPOMDSh5auVLqOP0yKPVHq8TWKEgmI6
VbG2lLthi1avhwkbONW8iO6tnbA9+RTx+A9XIpK2PH1VIGjWlgnPfecM6SrZ
leNFgrl/eyxMgjMY4JxvW2u4t5Ngfnj5Pp9hW5phWkjkwtGKBD169to5zVRS
wGECH07XCgSvWGEah6e4TC5djcS5SlrNdyTG+OxJjuZvT16cxFH0t6UKorf0
nlf1Z/ZYxRd7ppT4CxtdtdTquAoFvyYe96m1gBp6zdZ7Y0OlOCBKFntL++Zp
We9KAA3RuqR2jA5MU73PVrRGF898BEx/KDyg4SJjk/q5YQUmzUtTL8ZsNetc
Eiyr5q8VaNSqjnvdOI6dAbqzFyQKo6VR55q4ma9+/oDSPBpp9Vw6fDVOxvcZ
2WEB9TUHtlnYQE5bM5fpKAd9UJumUHQg3XZDgxi8vcBizCd2E+czXYik/eQL
+nEJPfL3kxJFUWL4I4xwLa4lusdXJbbQgCsZX2sPtU9fIqInQQBz0yY6aTEg
R31YK7KTQPeGpKGxuIWgotDCen/gPz3CssZ+rcqXUGUHBs+RSbUM1bf3jAyB
PJLglM6kb1ThzMTr4Ejxsv7s9sYGCpVxIfXOQolvYMfff6aK2FTtnkYn/JyQ
H1h5z5IMbU9fL1DKY1Qeka1gO8c0jm7vYWJfi5z+AEOV0CHioSvtaYCT7uHj
Fyu4AyrobgJGQ7dVGhBYKG/Rtyq3af6um66pHISqUB7UMtV8pBOR1R0mNh5n
LJVrWYswWZhgfVGviaAvEcSH1QlYf99SVZykowujymPW3yVYWFbpI8yTpkQ9
vnj4DMpixjRsgnwEUkLIs76+mcRFcsgkqd4H6wNOwNxT/9Pz6BGnslaCF2FX
tjhgNKUtPplEdoearwQ9TxHhHLJeJY/xSVrXm+elWJfrYRF/3XHVOZNAul2I
siEcgdHiCpbiR1X7GqQPbasanGy6Gs7uSQwnIoojGpRDDbhSf0Ha7Xpp9Ld9
q4BR1xfeuivuBp4hD6UQc5ZUkk850F1iBkPjGz72SJAtQ8oB8oM0UdXs9EcH
cV1zk5Df7wFgmqjwA+UE7SebgxTm3E7gL4xzMzVIePMrm8iw9hy9lXTGQLvt
jHcL8D9G4L6VgdChGYJqqbtgq4Bm4aJO0j8EG0ULoIgZvjXYB3igRLh/SC6L
IcW0ARBWi40YZqRlp+G2OLyVJnibEZBIei6dNqvnqaeenWNL1SKT89mCMUlF
r8D49GvbQdA1RmQCHaAICgo5IJLyIp2Z+B7S8nnkQrxIX1Mb9mEtIRsHvuzB
ujTUOfsfzse2sE8CLeSBhfBeR8NEP3IunuGOnnjpHhwkGzs1fTt2p7IKXm4d
x5Jge50lz4Ir53jmHOn1FFjA5yg5n91ynNo49N/HdcjApEkFQQWFRilbk6wJ
+JM7QQBZSow/PtlabAt4yD8cykM2cfQTWovUrSuSWx9eLNIcBCXqUyWFIPQ3
p+QZDQS1FE7X//1vxBsw/wru14tl0r6F4ij53hPrE0mwfflPY+xN7C9SS0Qk
QHhpl1PP7qx1bDXz3q3aAcqKep76IlQIbmzNjzubOSqYL+boyb/u9/mN7k9x
RSMNEO6MjUa88VypvZmLjLUKkQPPXRwrVjXE+jj0MfXIQv00j4V6pRFx1Gfh
Z1u6HyDYogzoXB6UB15uGWZxMxXBhiZkh9HgZ3PQbaGYtx12pPcFxr5BQUiW
qYvou/m1HPTivudPoBjy2UFhN13xHfoyiJ6PskN0E956la9pw5gEnAattt6a
NCmpgrEZtuKUoV12s03K0BxDIFlx8QgRi2SsZkqpzmVhrsQ+iU//SoHpU6yT
3yNLGzq4R8WY6EmKPPHUUv+DxE37E/rppICXZHQD8a0NZ4vQKPMmH1VJfu5D
2Sf2sOtxniWGVpfsYsLd3d6ySzvoxdcIzFjcWI+8B2UYZObgJ0sVU5Nph6Gk
Bnv9sdgBy8gm1xeTBq5K7QSYsvRmfcLrhp2Pgd3mhysz2EdKWmSAPsH4zNzU
S+uBOxfR9//zCcIZIjmAFIeLchn2PMGDVVt7xZ14Coh5TU2LrYlLi9QJq96W
1LMPtg9nEZ+wjXJA/YYAN121oxu6OKxR9jq1/pmfoagfyvyDehMGKy7WVDVd
nP11B/HtFQX7dwDLRNFKtAbczwA1hi4w3QRpna1EBjOmFfED1DdmTTEL8VkY
7HOEiKWMG4pR4k0C5wSk45b+02GVbQKexCCMKg1fijYzy85J62wGIKs6CdvL
qk8+tjyq3EyCbZ739aAQAmAPvTWJXkmbVpyoVl76eV2PQVrNCxSs5M03sYWy
OBHtrOslKl/iMIz/i17wrqHwA2pMltoB8NvlDMn3aEE1gRmCeLeTYAtFFrds
oJdGi65wjSGZogte33qIwo6kqNAY8zW1dsEV/uURc6fK7GelrvZye13E3qnj
bYtd3R8YbA0AS2AmJCWhnOkMbrOY7tjQi/yOAnv2QIuEHDk6IYG9bU5c/uK/
4CSLskqzugxSbo71Z7Z1CBJ8iVSkHedJSJyj5CIzkITNSJw8yrV2VBKbtmqW
nV6gRiDZcL9SIY3/BKN8D5rFXyPYV3SK982UeKbFLXPBBfcmIXuhua0JUqrm
HnyizMHl1/gvpyOOT0NVK0ayQbPLpaVHdLW1tpw8Men95TLGuPH1LgAI037I
8DgB0duP5mU77hGu6ldc5HEAKnpw7eNC58XJXWG3xB/BWE5wudYr0cBBwAfg
t9cQkecFfOu7Uz5UjO7DK/K9S5ErqtClOmy5ghOena48OneDWG6PA2cj13Hv
pXS+IPx6SmiUfTyZ9O4J3BA0A3t1AIvgAfZqcGkdMPpsb3KILhnVqDivvmgq
3z/ZQht3J7BuV3NaRWacXQgDmWxj6pqAf8MpOgoG/JemCEYLaLaJi5axkBmt
RBkCtKYGCQ1uYpVwXcarvWzvrsXp2IrNaaboCS6+32c1yXJGVTSor4CZ9lxL
1ovsKvBkXLNUDKLnKABNG7VT6rV096ZV0L37uyuocdrWap+J79OlSrnF24p7
wTS8knv/LaCZYBUEkSJ/Li4plbSHoNTLqrsXHlvHFge3Da1r6SFRqTe6WSLF
NdO1d1TMdb9wrWFJhAs3qMPWQZkIgfZs/TtbAl9K9oJa78speKxlEcY2qcEw
+I8Btir0N5fKNuZetv9Hi6UGfP2beCO2h5vFVsfsf7d90gxhkGsuTdA1bPuf
EUgwpgwyxIZouBE6Ekw85tOmqew3HjzbYJ83EOUp+d2ujg+RUxlEksRdunrg
CzHv9kp/71KXOI6iu2yn24ivdecVQID5KP1JA9SGDvqzGW6b7lapaP73eUYl
gwpBAVsTDtDc4Jy6uN6l3kiArU1ag7op1Vr7neoHnc5Rf/BeLlZYogqgvUIZ
jQ9fvI4lBj2xL8iPc/4h30benm8up6W6p/FrvPW0oJFiuxveYcQLng5ugv7R
g5RTQOSCp4Vr/clYjF9Sb59ACYOxdkUkCUTVwenVLcBnD2Ikl8EV+TdcSdYT
kDlFRYHtnqATkKFciRuO14Qs5Vp9nKnIa4oyT6XjijYuIUBeBJ3DiFCJw2z5
ZWbRqVQsLxp6ROm7FqbavufEu49ipPrFft82iJcVuu6+PcsAZEz7npUnISZD
+B8sRMv3kwmIA3EYXgp4T1FzUtR6X1q+TczAFkl7cEKRKhqEwlK8yv3Nda+r
QvlA+b+JF+B48Hw/rP5dAZWhdg3nAYBIQ+KrQP5YnRM+s+n0fXx+OFpQmpRM
zE28FYYD3/NnqVooWfeHZkkLT7bKPZMA8ikH6d64omhEfb1XEjGHBbZD1C88
3zzIrtS7ZGKvEQ5EPK0lfcslzlu5k4OgY+vjUQ/a4SIMUJBT1EALurMKBYC/
GCo0OVIO+hxKLz9azpHxjJdOAjqcOhe0/36BseDMjNOB2B7Ejbf2o6+G7Cl1
boNFOMkxgJx/hfeofKaGPXf3fmOzVPm0iffrvDn3i6+AtkElS5euKUa2UuaT
MkdNBUvM6HmRDqzdlJ3/MmXGZl8VH57blC5WjT8yXPCHLOe2qp7Uja0+fsr0
KmlajDsLzoi9vVZ465bgA4crzz3BXi6QmNhpcKcSiAuxWLDK0Fo4IfZ6QA1n
V5H+Wy5rTzn4L3w5hFCvBkEydJzySNtu/K1yGOUY9nEuQMWIbiizT/EjSQsF
QzEXjTo8xGW/K/GWyNnsD67DDm3YyyVjbKMfbjYIAJQOdA9Rzrnjo4qnqeEe
+Cue4q1jE34o0aJym7mn6QV5UccVhKvyzrAzbXlh/fQNVr5/pSQsmLxV02tk
Oz89f9GtQZDsscSHjaSdraVzLnC35k+U6oVGepcKKC1SHxCtP5iuaYRPztbL
hXr2u5aVB5qV+mYVEwU8GumnYm9RXs4x1lvSEwRiMc2D4f9iejFNf5YYo8cN
1E45/mQkfSa7vHRYs9QceancGoaXH79JSAEzD2MemEghSOrcW0aDS/z4qlQB
atUJ9dbA4U4BDvWexEMoqyEsPgVm6oIeeSFuyhC0m7UAVGXjirVfJOtOjoL/
ZKPYFahaMbHhM6VVKzZOakwP3sfuOjzG1oFHppYe5Novk0t3z+XF1b3ZaIG6
L8l4Ms9lc44YKkPMisMhYKXlHsriurKW+A4eN18ruXPsGdOd5PpRUBHzxh7y
wtjCgm0kC/uDAB+YHuMUatunEUvC9r9OPP8CeWlmwktuwuZMvr5RaViROY5o
RD4+kTkiMkoGX1+LEbMEEpZWzIVvq8+0QdNnqrEUNIJmRRS67rSq14x2xc8J
doNiYtTbvBLI8c3IRywo9KvOPehkHO/dR5BlanKNqeGX1EemWkxh8ACFSGGC
fibEL4cqGdm6j8znU1CEF2s4loRqR/IDUALgyu1k+emEy1qPcrnxLikiZcQF
q8DjQ9F+eJMqUy7Zkzz2jWk0y+YfoClaw636/uee7rUEOv/u+8hlbBserCBV
OOzhE43P+j14iaZ3dLdaEnUaiVDKf+WF4vj3+RCLs3e1hNKThnxxl9epN/HO
K29WrpyuAOEowsfNCCUN23eiRSRaBdH89+Hq76EKMApS6FJ2avhqotOI3kZF
E5DkQEc53f5lC9B0XYKTzlNnbARupCe6DtaG0tSyhuLyWsXzZ0iyOhTyP0bg
jPW3lOOo/7HBr2L8O1g+6wQA6oIyO6DUWPt6INwPTEBg+P2TF7dexOJShwM/
rdeN5dBa2yjV2dn8Q+3b99WnGA3Kpz+EriwUm2D9g5KDQCaIMOaUMyE/qcjp
vwG5cdLHG3g+xfM2M4VXwF+/obgIqYI8s2cQpg0sURjiMfvb8xBsQ3aziIdX
Lcm3i5VmIT+QA/nirPImzZnG/O05ySFe1+vu5Mb4YY1uT0HvgwuJ1FD8IK4D
JxcUeJVKVH9EXEw7vRSK5llrBZlRFbJvD3Ntn53bvt6WaVcUgwT3kgqj1PDc
cE+JMsLqRD7grsmbTesTvB1K0ul8iNQZFGjo3E8RvpCcROFAP60Q15booV3k
74oE8zSXjvkugS68CQ1UY6kM812wj8ZmDnFXnf30J1FX2KwJ7Ye4kUF61Gxy
wGmImOWKma47po5oyabDw9mrZzAJL0PAYFpsbAciId91PEwkxsFz4KwIwsMs
hK1jvLmv5xo/qc9SYo+R2RwTO1sDPtLgbiOpw3WgHSFBkUTge6jyB3hJ0bSy
JIVxEalffpkHJtTDe2wLeAthFw+lnLkM3gID0OBF7fy9x3dVpwyfpZBkmAH4
1O5uOOICAhw5V+p6HaWpyRe/k0wtjeAKL77km1smrx+Zl2X8J5XcpsFyWzvO
f6ch2pVm9W6PHjXNsyvmz1HzOYthPvm51VHdwauc9bcY3hnSva+zwi3WTsi8
K0rQ4ePxe3tlIvGdGWxwx9/EmFG6DUmFpyeEFmbuwaDhcw749zkZ8ei5qlbM
92nhUDM77rJZT3Ro1tea+gifgBVkpNwzO6/IEhd/4w6jRRNsM2TcYzc8jGAV
h9KL9pjU36cMScbcuM3oLHD1JStPMgMbhAIWIAIHBaMWIkdk9vLESv0sqHYF
K1/ikelJ6Av47zPTmvEqtGDW/hWkKjefqaqmGSeIaJ3FxQ43rZsMohSi/KBn
HcMk3Z5DGPScMaij8IXqlVs6wg5LFH4NFAXwRZ7Qf60A3gisCH+Qzbnigskx
SxQtSa2cFV3w4QJrdwBzr81QdtmhJqxE301RYG9x/oLRo16/EsfPyPTkuZUx
+lpXB+fOPDe5X8DO+dZ3KHzst8zXYIcLQGmM1+J/Gvi3gw1nPWSLgnFnrO8k
TT7BvNrQuQ8t/Btk/FzkaOksK/sSwaZmMs9goZyY1mtgnxzn44d7aSb8C/w/
YKjf4R6tWW+WpN8mlD3yabGJriakooIZVxK3YT05nSnCo2yykdDbiwRpIQte
R+PFsYmVDaxYUqNhk3PLXkuRhA9jGbn69JyeGMZsY2QU6S3aNXYXY8eWsLu5
SNaKhLhulDIVLFTikhqBGXkjGOc511dTALtULDqRHvJQFLG0t3pVKgVvbZMj
xAeiBNMmOIO96KfpGB+Zl33Hj2lh1pKB7Z0U2gFHpci04pChfuqawSRwIO+b
afg9mhZRTG4wplIhFC+dqWSMVcukWoisdj8U5IuAXQhHTGCvdRddXRue8f7T
8pzN06rrhcS/utbZ+dJwIgN6+ivjbZlEHW0ZsMPR/HtQ2d5zfBRA5G88i/Tu
jvPD63NCUAsFCq4P9F7rySzppR5XfTIXRiXz0qpxP9W7dku4/kVActMOo/pN
IMlLwHfZZ6CFX2MoQHR1q1Mh4rly2FfjC5GoAUP6lGZYM3pIY+mfpFgTO/ec
ZO7AL4542/ZM0x0h2D44/6iz0vYDAVgmcV/geERHSYHrUKPV8NoD75N72Clu
6vszPXKPdJUlxmQ9EwPrbtFKsTpYgSyvM3Gui5hUTQi/FsOU0tHkOCT6djgm
QFYjynIMMY1VBQSKrxRUYwyMl6F6IXU+pENBlNlQk07Ian6zGRVM3Og8UP5K
hotT5dM6RsHhW7JluRGni1iMwyS5Hd+awzCdabp8utcQrj2lEQj7tgfJcr4I
oJraqZSnAiP7IEs8tNFzFLJje8/Xyl3SLxMvyIOfgh7ZOBsb+mR7b1P5M1fW
aGxfSO6LSiW1f4TlYaCcByKPFj0GaAKXIQY8ppP1NMQgIokpYeifDVefVY1F
A/teaHxGS3zomYg7DgZS0FrthXVHwuMI1cXjSSw/100qT8axHzZjkLIMZ+sp
qw/8QymCEwYfOTJl2z6U5PucocmdFBIR2odR82NJccmi8p3t06HuAqLOEsmD
jI9kmf6/pdTJyTz4WbbUTDZ8w7hAr/A+YUrpTRkINs3BuwvoWSauXvCTTc2I
kj/WVLvrBC+45mvlBS6H4/KsOwq90qRaaSNxB05Z6rLCsbRWvV9I3JWJ5Q3Y
kQ6nmBMliqxkN81B4ga5RXsqWLBQVMk2rEzBE+dCjo2Fc1LrF6keOoWQnT1P
Ij2s0UYyEXo3rxr/mqAWiRNsAv6cNLe13orsuLElfQeRNmZXi6zLg8bxqv4J
WWNYWSFybT3ZFqJ98i3W2f0YSd0uUFodD7x/Xnc98EE7V776BP3+j0uZJ6p9
A926sssDwtvZdFu8i3cooyRF7p8i2wgEP1qgMNi7F0B5GW+1ZThq2w/RW5fb
JaVn64jTKByMK2kVUwI4ZAlvDPPYE6K3iiXdkIEm9StUYiEBCTJY5OC5ogt9
7IOiEpz4jfLpFAWP3OZrD+0VV48FBw3W/+idQYfxocZgyA19OTG6zZbw7SFo
NaktRN0CtB5Fphb2OFO8JNy0QkpW9xNrOkBGqvjXLl6AfCmPRw2Q/DBx2U+U
/zGLRD3Xo8Q3ot0rest+SLmJxXePCBXszVA02GuW5WoOv0MKCeJ2kU00GB9F
CFX8Kl2DfgDJ+1t6GvhQo7Xx5W411/eOL1HQa3lTzWlbWXQnz/9rvHDpx83u
R2MYZg+qFbLJ+OWtTOyUgfTnWL9KuJXeJ6Kgf4EJ1XgOzTMpMV9E9ko5k167
6OX92XNHQ5O2vf6169RV3k3d+bguk0REcl7PFCV85e1htc5gPUceuFXsDAA+
xy499ZqYRUOTOrjDKb+jCyoZAvNEcNmqvjWfNsyuNuyu76oDa4wi3Cu74K45
4S4T5CvJGrZQdR0yBmDL6B91yJvB5RMX4FaLkod7J9fr1g3186y7PLAUWVO4
z5hnj/yilQxyO2bPijhIRmynVDTysoijM9mXU8p7lzUjm3CECM3jK6vTqWAk
xANy1bGo7vJWQ2Dadzu1v4JsNmTBomydyHWGjHYhWUthuVUVhO/5RecVYNHk
gx8Zeguk6jIc1+FXfrZE1yjo2+sZ6JB12OSGmy2y2EGBYhxeOMeNKoK+BbCI
6tGapo0vsv6MoFWyui60aKc3rB3a/7xsrdJEXlPp4LnPqH9lG/eBZ0HCUXkh
psqyTgnMswyE7R/KJVB77oIBon5dBD5Belcw1ks7Iq15Z/+uCXrIQwfqoMzn
S3nluPuLF0JZOkb9RJvPqVjHfQ0/1V6o5au5yLehK1obfbfg3tiuA/eFmqpM
RU+Ud/ihuMKyjS5cW7mk7t8iJWvK9WipEoNwmuNsN1Z4XN+uGiPCw2Eu2ZW7
tatzeaYPuyiu0xMI3Jf8uEyCPFdqbJB5fKGC0DL9s3pp8a4/xTV9AxhCaqtH
3+ClPBUPybI3eV3pNWDXvRN5PbywXt1Ml9BLu66n7oxN+7r37KGlZG+ACL4E
eKqi7wCWj358qC5O8adQKQLejyh9Vavzi1KE33MuX1CF9Fkp1mHTBGCXMyRH
npMN4IjxHFc5syc0hCpEjrYnJlZYt8P0igWxy5eEFTzzSeUnd/F/pG8dCd6m
Ytl9pPXpDqVz130PHxg/ymFLor2rJfAcOBGt8BhzmA9clGBXqfnxnGM44ivB
dHPuTKU4kl1xV+Xq1R3UyOGHwyq99/FJRmHdHhei85q7UJ/iNj/Rypnw17Sg
d73YdLy0BLTdSMPZWV3NkidrvTFE0zq2IZz7YLdcMhoV+YOnYrTu0l8f5pDs
eFxic4C/3m5UPgWJQ/8GEG3wcBr17PCkj6YEsn0rjKxat7orRQWsBPL+a3C8
8HUDBnmFf6b86ciYHJw7XZ2T4ThQXXVCybKHJ5cidiqtuuQeJ0uHzhaL5XKW
5OPb3Nu0kKdVJikVhok87HIH0K+ZEws0zWydyJA+gZpnTZoxXq3oEOrD+JQ6
Kc3Tzdwwelm7gsLmxK0n5/fvt3uir9NUXCIOyN6MGCNkeBJ/VWl5pjwje2yh
bOOEm3ab6Bf3beFxbNhg9o8s6ppq/EG5vcmU932YU42exgsccn7+iBfCmJmh
W6CyKmCJUVsqQ75MBOksNGWVGHFo/ReKpNzfhHkNm4ySlHaurSM9CaLQxvvy
G3zG28HWcClAHILuQLTyPkFzO0hBsvUZleJkGwLy5kAPGmelp8Yiaj0inD7f
wKU4lXro4IdWvF+MniqAS4YzRIwwbKg9tHob2VWRA4R+OfI28y/MSzAXEwda
giE53KnE0YSjmfsMYJ5PyvBYIYLwgZ1+/1hm6WLeD1x0iHAxKsq9wVqmkSo9
NPnt5rORjYA9mtCdWpbrumSuvGbRPYrXALIbbhelZd/J67SGEj5UF4Wizx4H
Epal9ASDMl4F4RvGomcVO3D63vMl9IPukT+WVz2paB3f5ZwUtPz9wBen9hSL
ypuQS3hwp/2Dzf+KTwALe3ZuaDV/m3fN4NGxjJYFlkbPHtEjBsFit4mmARIw
VGedI7/+l7gDSpQIdQkBpoxhNxnebedxpAOSovyrQEsWPg8cIraO615rRFQ6
HZQBTuITBPGT4CloxM/a1E6Qa+1XEqdIEN2xB2Jx2YipUjlvcQDxuBTKTkgG
bf9azvliJ5U+OQ+yS6pCrdgxILA+TeacUu+s21DVLfqFBxOLBhMrrgxBOThQ
7NIMCnCZcdQtgtR0/adELDMC+gUlipRHsh/hEzXMjiP63l6oj3KUiotgqm8d
1r9AdXIPQh+5MZMmDDdNkVWC4FgGeWKZQN0XVxB7Pf3UUmCku5pplBytZ0+M
F8EfwGthRVLUGSY33o51U5p0vKlO4A91i3k1G5KFMgNCFX++zrfYswzqFJBg
/3SS/3Ocg2Q3hMn92WRh8X7A6sM4zTCFPdONxeuRp/pnhIbwCb0WN6D1XWTs
tw3qNBRTQwd4HaFel9NplJb2X2TUBzx/t1sMOh+aFpNp9lxBWQGRIhuzdMJO
pP8dMAm2ESwOfOmPoHJqfEPBZ4uvpM9lzvg+uI4/ITOyxEW2B6Ia7tm80Xme
xgdnJ1SSSFAGer5HeV9V5zV2pJbPSKDEgmyejw+vghOOnyGK8lynjN57ZKWf
Ebc8tvDWJI1qYpNf0SedRRhGcF4Xm86iHulV0ABXCFpb/wREcI1BczAU6aVP
kpXR2Md/2dX4QxugK1TssiOHY1VIyRYSBJwacL3qAK6GBEmFA71QdBNMezSO
y9yiEUG9i4lBchaCBPsTrO6eEJMCHLiHMwGxvetk/tJan6k8BPIyrgdCXdqq
gFTE+EODRhOS7cZZVguBZxD4EFG4sa/lDiulAQxf+3ZePdC0MeyzNFmyr9jb
2nW/V8qv9YiMZrPkiUq2Coq7rH4EpUE1fYvTD1GnjnB1h/8cApmE4jVLKL3+
Y8pEU1cOIDwGEJD8Eeka5bSRJyj4qHFqIMYqXAvf/h+AdzO5wPGkE25agA7n
N4jGzqDCQet3szoaYDya83tXvCWIHbd6x3U7la3O1DbqMdey9qRZbw0BaqQR
a8VElqKt4Nqm0swfFk8M3c1NT78F9c7o1p1D1Rdv60+tGcHD5fOiPoiNKzGp
dPWIcn342IJGQKi26daPya7AAI2pfh917+oZqKpG1trlXpZ+ZV2oEQtUNGKI
iuFd/Mip+SJSCSarZcz3GhlmCiQDVsWQocG9iF/vsaj41II/IOaJ0zu9/Jbl
wL4dXEZ8WjbyiZpEKXc5D0nytp+/nTe+l2YMjydRpFtje0/NL8dE/mE8oc2J
3j1wztA5VOKE+KEtC7Ke9iKFeDPbzAsBaFuu0U655eVHVjOE7wpbhhFeqADf
3c9kC/smQUzjfB6GPumBNxjPzrOz6Dv8Mx2QCQTo00a3Nh7IrNDKGI8KleFz
jv7wkAqmS2/r1L6yo9COs3Hm/byGy+1Iz/mbMThBOdv4ugDC341Ly8sfDjAf
d/T6z/3wEVca01jxu9+WlftUUtDGqVR2Dx42bE+u9LzlaHxOjJxPpy0ee641
9wH9spq4eEB17tS5tIIig8d6I5ehpBHcYqmzZuiYzDyirPlJeuRynrENMALE
EhcUS6hipmLNIKfbAwiCftaafnlKB05HXhOqy1id4qM9ii08zzmcAQBTmbJw
d9Idv94CTixGBi2HqZaKyo+TGgt9j3RZldBwX/upEEQBF4nA/8ZgO3QketJC
3012ATlA+hKs5m0VkKy0cfzyiSeqBOx2XHRnKJCMPgDy39sUJt5MYf1tjTFM
P11JETLeeMcLvea6pvW3yDaME6DNe+RKJvbJsW23YtrO62UiwgzGAjzc2Xey
ASh8X987VCEXU77JdpUVF/OrGMSAkNbv3MN1HbcTQV/bwZI5kysmdX6zeT//
NJx2Lcw+HXK+1VhgzYr1QWtbJDp6Wz2VXBNN++8ygOcDiJeBINwt27PfCctQ
Tj76RblWbODAffScksrMBQspmezdPVQFlGzKt2Xo8YSnhVXWZM2f87ZIMXjS
WQTXsEtM/UMMmcj/Rbmyuxprv3vKqESf3zeo0A3axiFEW7TDOPaO6ttnEBMj
M3aQkNpRfkCrjiH+qSS6zmL+k3H6fFa14k4A/FsVfHYILryXSS6fjd7tb+z3
zq/nK73US6kSW2EADLtr1dc1DXwKYDGGL5tRh4Tg1KO/BW9Glbn8IGP/HSZm
d1IbwnnWtnnGQBLrHnOOw8zAPMMj4C3tZD3ecUsTsno3kev72ZkWOvZ0wbP3
r1nebPVWRnaURL2MdYIT1eWMsu8BsROOjh2qC5pstfYWo0ziOMlYfxsRMMuf
zSjukG7uXz2lniG5xoo0Y9IaIdHz1Md9HHlInbOWdPrsc9a2nJTPCn1oPbJB
5CjMIMtPGvrUCvUzcOoFCCaExigt+5JPy0HPrAx1zHYF2aQ/bo33WMz6LYoT
xpBEf2Y2JOEFDQrb4cJPZRw6TKGOVK8upBSlYAwz0ua6SIIeCguJtan/GMIL
XA0w6TEInfuIsaiG7vYiXRqw8NIlW4rVwF+EDO5IAAlEJCGI52qIMXiZkenz
1ji5GK2OBYPH+76gvHF40tudZwXTw5f8Ln/GK84OufS5cOaYZu5inRO1ZgJa
OADINZr+W4HCSoebKyggbki3VbYdeNAWHvKHK44n4ddpt9B6BGVXQ7QyFqm6
0BvgnQaibVkSR2M6x9q+p6urSxlSMCf3v6AGpRa4IW0ak71vcZgCLoi8Lk4m
4njHcKAOTgDjINvhl5yMxgPKgbsTgjDkqYZFQCmrCnddOxg/SRtIJZkFMF+f
hrvgdUkKNX+M+Dhc35poN42MaDtVau3cQBHJv38lrf7PjYVKz9qR2rsQgl3r
+tV2vWOSZs64WZSGGW9TBt3MpuR6MxUnXtjVR9v5nfXDmR3J4Bg8ARJ7bS/t
UuNzYPnH6o7zm2ktcQ/h9WrIDl9JDkMWOokHaB7YkPmdfJJbh7aizEKrJIqn
yOJMa2JidgWW0NtWyzIfxq+8Vfr2g1zqyRQfArmJ/7hwxixBnaf3YjsJv3Yg
YC14b/pdLYF0WGVbq2F3H1CMm8c2v86Jq8OsKLwu4ftu4833MJQDeGjTU1tY
GQ+4ptfjul4NcDS9KI1mwsbqy7iAiU4L7e4EbuxBkp1Cbi+I6tIFrvpnHaW4
pYO0v1zv61Zbb8r/a2DhJWNae+IEL8p2oJz1CC0rObisabt/RB1EjApkFDJE
VFZ4NmI2LAtQTnIqqn9wn7yxpHKx9pPYocwE+tcNuGYaZ7Pbahp7Iig5y06X
Z0bhP4LgyA7lh0GfpLcO3ouHvhU2PqFDxDARvQKMmcLPWznYvtITM5q7q7M7
mkUUubZOXAo6oQjgs3xRxP1Pec6pgwWWvtUr3u4wS5RjGXq63WUyrMvtKvhM
ALHcxH6JvBvUGh+KCt8R4bSkYeYOeU3yicS0J0z5S8LdM61lUB2BNXgtl2B9
9Sbg3uvfw0eb5BTD49zrzzTu/ZiOgPzNjc5L7hqrxT3U7sGhgsfBzrWMLpsO
UxN1mInJqDtBGLX1q3ArTJGug9Cp9Rhfe85/CL/TRo/UKUAKMgtHAUVf1up+
nC/48KKuEdbfYFICtEKi1mrI7tpHocIzarG+XidnQhDcxj7W/Aa7S3THZ2ZX
gM06c/GK5c1jwtAImftSviIC751UAPxbUrOUSL8sN2RfLuNhXAMBCX3BS1df
Fkk5/jDfXto8PPz2h4ClYyhhTZv1WYHgmH5y+NMRiEZI5r07AL2zk8UT397+
VMisxFPdfInhPwPbE1+I0dubJn0PEuGPkgmImLVdI6lAU/fZQuE8ps8GorrC
VRSbRrID/s+ZFNYQP92Qqe5VBRaPd8XOnBsuF6VtI3se1XiPMGHv4nk+oarY
WuDSVqYoayu3TFrcj6eGqK05xloIjRBaKtVSjdO2uOPUgXm22bfH1qgdv0lu
6HfpdvxKlCWdfhVD94yHSN53Guv0vw0jpYEUh/Thpi1sfLPwrg5TIG6ff2Sa
pd/R2zlSIOmSRBDRXEbuFERCjvrge8rlBKAhZ8BZ88LBgsC96xvSjv7l6D5V
2Trb2MBlLXsFua1SzvXoGVyKYgj1z+VEAyjfqom6XbiiwTQ6BB7mA8G+VWRC
zw9YbfN4NlaNQHDI3FhTgJwzk8wkKKnxpFZvY1mTn8GVS1AxxEhiZN9w++0Q
vSa1T+AGrTnY6WVMlWLmW0UM08DyyB9trp9XbCvmrt9zETV7YmWaMOm01ZWA
/lZrSqzJcaIdH0VwpyN3IZSZqm0H8AAsJEqilIaNMw1GyRfaSmPepdys9ElW
Oph5QwZayuRJg+7V/CEaFuXggnTUnib9q99CD+2zoI43cfBLngPZXCd7hfmq
cmmNpCnAdnJEj5QX/5cuZUly93lbHLWwcqzZ1Zua43BLBI23609h2Rnvkurj
kTarnJXbx953AND26K9ivpyTJWlXMkPrNqF5lAzjiHv5WfiVFYBTbZ/luCbS
pfhJ3K//AEUvRfZeFWYg25kuu7taVJeV94wDgtd+bqw9IVsV6OpJ/aK0fNod
eePLFokgBoLZ9aJUcJgRvlaD5nSlAlQ8VPdy+dGyQwp5fbHE8CXrwu++os8x
1azO1WFpRPJ+1VYVOjxJiOJSegHUrEnsogblpcG9JalM6L2Fir5mrl4VXDte
VeKC9vvIjAOW1xOFTq9jJ/wwLTM+2OmaTJWAfCRiqW/86N5qsTdlHaPyeNKA
XrdNFfHdITRTFlv9N2/llK1Jv/gGzv4jiXhmo/wMoMkS8K7WXsfMXuq3rWe8
MooRFIjXwU+k6TgHn0MAOIuhV3HW0eOt0dzUGxnmUqLAFV2ycMob0GgSuJOv
IWnjbF/d/o1yD+6W79qQPkl+i5F8OOMYAMyQzRsem70FwQ6jfTY4OdptrXHw
QXYak+lgFTXEnCU4NvFrduJznul3cEdJ3Zn+pa8CC/oqoIEeVJ8AtuDETEAd
29BuWgkABHAJgI1Ayat+LZt6atKP8KsEdYmBV6yeBO0bkDfbUXwO4+8ml/qF
tV4KfPsb/z01GB0Vldqh/ujVls829ZzAUNGa5cIKyWTLQC4YzsgZXFJsYCL+
FGMoGzKrsAgtusRHyMDFMxZLOMiFGKc7tQZtocOLOHEisXLWSLd+qL8/hBpP
E8PxSJsNJuW8itkCyfPMF1Xrk1x9dQ7iZviDP2BotUzHKgsqsplUm/FFT5qn
kAwtB5DQH6xaN1ZG0aVvB3wG9k9G+/RvFx8KkFckmSY81+5m99IwfScT1OOj
ZfN2ANlAgJxwBKtiKu9hDif6/HRMQ1TkkgO7k159aCJYLiv1TQ/lk24Mfegy
YFthsDqSebPt/fxr7ziNaJZlOe9PnX8BdOycgJD/uJAyQ9yw7Wc8bWbw7VgR
LGEjtOac+frdn65SpIeyrW1y8tuXimVWvAHYdqc4Ng5VYgVuoh/zkjZbALA8
l4OH6rE7z7EgD16HORjazz5oUQ56kUdNwjC5SXZhwP3Vw+Ui9xbOZc1heF93
Wawbqq8ORfEL0j1xDxkKNXavIY2BjTPQkWdCqTWKSUGxx9bO0KhAztU3YY91
eIB9SkK4EVVMZW44qCHyexD8QQCLuhIYN3aIPgIa4lfOx5n2su8ZlVSVyfD4
6mCHJZeqz6mVkk89TkAwLGI8ANuOroO0Ay0AruvSdHYcky1jjebJGLKQ+Xt8
vYCw2gpWxE2q6uxndUvjWW6vKPonoGP6Szm0IsVvli/bXfoXhHWR2k/+VW8Z
0CdnkR4jaaIfrWl/pSzMSCCoauvEV4awe1y2tEQe/l7O5duRw9LpSZWtBu9g
TnwaXreYKVvCUOf1fvNJGFY1BbenzwDy13e5Wz1Pwr0drGtJVyP41YcDxpKA
RrpRaoXAl3on29zRAlGNfUtSSLQf11a66VHavXZ5F4FnwG9WNvvH9DhqKpMC
4WOUBOFshx0BnSCy+mIHXXGltTgr/NeNe8z6aCEgTw+VJoOEv/R9YZ9DDXjM
P4ifrpyZ4ctULRW7k0CfNJCN+AWNiNgRnvM43fyojX9QejgwlgUOJLsONM1x
Rc8oDKd24A5Z7+NYgPzobANDvoF2nsfnIcvJtnDni4PdZ2RgKLIgtIfLKL84
ZvpEXk1yw9fWo6KVTw5n7ONuZLgtR5evyWNVGbL0V5sUC1awTNRGvu7R2Ybw
TohqlqcUVDIpS/fkSivKqXsYvgLzJ6RnqKimh0t26cOEVEbwI26D26vrZCIX
Pl4SfrlXEnbJFRwa/QCAn072Q7P+zdo9J+PxumvpcDPvkkjTEcEb9gvF69Ul
HZh4+rmssqbnVFyjWG/5SINVA2G5N58cn/3ouR8Dk1l+3+Tn1/lZWLwuyMBO
Mw6FiGmzWHhNLYUONyqdN6x3C7wun0ig1UMBJg0DnEVLofNELHNKbSA3htvM
gTJrD8TRjORYuF9QWdutus2hisRdak7IEVVNyX9X8K0paMnueHM/YN278Fl6
K5J4pnC/tmbKXdEskvZLejJAjgg8s2s/8kXdnEadmIZwg2YwZ2rA43fZcS3j
XCqhuKuIUE4wJRs3YA1G2fHmyy2QPAQF0wUd5GVe/fFS5z0beRUY+ewf3mOF
HEWHTmvACfoLoZIaytwauUMg6aP2HIdgoUUzasnkZqx4uO3k2+/XIV7Jou26
DJ9LgqxdFvdEpJtFBP0m6lFZxrzLlm3RbuNGc5AtHpQBm0xsqhEgF942VdQF
88c/jUp1TJ75HHqJc7uS6982hNlM9t4e9grIuIYcaJgeYwwNKqXNmEuvsLcX
g6g1VoUxAp88NGtHxNnyyIdz2XJHW8uoQrxp7ImTtZWKp8RnKJk2ZmoR6K7w
TxgzQK1lLrdmWaWK1XILrCiMYI3qCryu+WQD/ZKy/sFh/zg4Luq8xI2xWN88
fjVzdKJyc30ECUYYUWUmLSjO+ycof56pFhRIXnA1LXg2oStIzHcTtHgCWdNs
01wGVsNgmlJ/P4iM/l9OjcVLyw396sPoO2OznGhR7IpUjLrpbLF18rgmXWhW
34ZzAfLwl7zYPpbZTQTPx2pK8s+Tr2YDAR2CKipYTaqZ2b1TFFmaznGruU1P
8CL/cxYwtNhfn7CUlsEJZRPHi2PEaSkiHNimhp9FsOzYnKm+5V6vfO0hNtx6
xnTEPqTCczSl7Bv5zve+ZmsXP4OiSNukL9HxYlzp3NPybYjdQbB5QYjw+yJb
MQcRneaq3VNGQZwmBxj3FGZAgSWPAh1V0PFYyrz2wlLilBVRpDtXHii0zl/T
7Q7DXcBgQEnDVOeSI9ySU7znvg/FTl2OzwsEj6EN/BVpHLz0r1MwQEOkijWj
sQBQX1+s+eCXiRPUeTg4gvntYp6fC8yJC1DJT8N/5rzM8p6xMYGHtnNzBOy0
CsFpaUmvgwi67tHW5fiGxOh80Wb4jNcETlC6Lg82C22xm91KXayfhXQx6Mul
OBP49UsubCrKeCw7oGmzuWfyFGeDof3ldFgn+7oUtd0Zo448TBZH1WcpNVhc
ak5XN9cnPoNsd/ByYJSHYBLyChbMVyezaGXkQA/opaf3RgQh0TMrmEBXv4JH
MFrvQnsbB+GLBeBizoGj1mwGf6BgFu7Z0YTsouXTpCtdFDbY2bCfBWsWAu1J
H1RKAPz2hf/MzYyPij15KbIKwYgNyXjS/UvJ7t6aHBJa9a46v7VHsA08Ibed
9iUb8wYjTGTTaqxFLpDeElZzckGiUg2F5gpMsFdAPsMyOlfAPx9qS+5U81iX
RhRRXSxsyRx5PXt2A1Z1MWbGuTn+yrlR6u8KWxV6ZZe3Af941N8yqzA3oAyF
UbsmmIowzIJwykI/ePqUimjCmerrYKNJDsWJJbfKRIOgqopqnJz+1WjXU2Wm
BDASyXeVbMFUSEl1JmGNSA1ozz/BtDnjwl1H4P65OntCxsg33k0v5I1mQ3+Z
MJGE7A9sA19lbL/hf9t4Od05SyVb1m/fCFM3viyiWyVx6zAuR7+fg66kgF2j
dF1/3nFq0tqbfyJbbT0IdekYqxMSpQLvnN6p0YKAGW7S5VjXJzsZYvxi9m2+
NIQkNltdDSw077/KU8jgwfdV1U8UtKoQVr+/4ncT9j6+pYuQ5WisO1eFTxyL
NIPo3m32DaXTJMP/4cfKvHpPJYZ/T4JuHvGmd4vILUO2Xm9wTkwHczJuu/pt
OZvuTja+llWeh1xBY4gHX0J7w+Ypuxx7oLcpZ8Wvib8NPHcq45LRWT8NrJUL
8LxoLFiJPWWfs3dHRYkLHge3kci0I0iZqRljBsbvKoeuefPh/c8+fh2JYhRE
REHmjZfdN2Tk7F56x118UE9yRpIT7XRzRchTI76/iHBjpfUl9lr3CFUqhW0E
epjQ7OYiacju75MsBrVywOYOw169X3iDNRt8k7ivccmI6BGUuW7KjGcBeYFo
i/6Dmksca06lDAQsQajmGrFAjH7gtIOuK9cP9Sn5y1k5KPaDRNlMGark3CIC
aIPNJLV1CCdOytBpIHWujTKbYTMu2CKC7Xs8MZBS7sRph3cenhyEivMiSiQ8
AeOL3SVKTs3pfusMCXWP+ioicCKfFlpB/RExopUw0yUqFmfxS8I6MvXSdG/F
SQBreGkoNJScb+6K8xQTITUA+4VudI9RnMSEfLMXlk90+am93/N+KJ9gJwDj
IxUb2UkXut4V6VAIQwgFx1w1Hl/COdv5B058NrjAMZmVP+UDPHCbk884Ov5l
nQ/f78hxaWd+9wiPiDu3V4ll6niSognVONxf8OAhX6iFUtksbNpv9diY5Lzl
A8AjgDH5bMyKB5HyYCU06Jvb/CeKMegVk72W8sbdz2tuY5OOiCWSDZ8PmzBM
bbjQ5TvLc+TkyEnPPucXO7bdR3MoQ6fFgxjvq8bzzrqGRCpiCdh77/oyucXR
phUT6eJqomffPfLIvNNvjsB0m6PJWU2ehsOJHPtfXanZrpIzG0LQsVVrgpPn
9LtAWwJuqBu+SmK74Wjs84+e8iH9Ht1puvvDaeR6+X9hs6tizpD2agBXF319
KgbcWgECCgNsc1c8hNva5rFY80r4DFe+23tNALGARrp5Yt072r0qxuYtFhZQ
kyGrDld99Bqp9Y0AH75cWAmJ4CCxDgcsnQBd0xul2aD94agaG3QhBsQbU2zZ
b2X+kIVkJwjEEAnxvP8ZcxIIstPG3plb6mw6w5ZZl0ElXroUY7c7sNHoOgje
9r5vbLijiDqNQjgh5SEtBkIpjtDOAWSVNoX3trOn27rbqgZ4u5ytYDSDudVK
XR1ngtFyn32lon0L+0hSWSoyeku9P7e4QikLMk2V3+7LCgtlXC9FQYRsMXp1
kNL+p6kqqIMKTLYWZS6txJIjRASQgW+fxiMQw0hcU0DL1b/HIpdlCGE70jFg
2sZW+KkTAosV+vqhJvCDRAQdhuqknPQ+x3Sg94NcSPCnOvX5d//Xl908oD+g
89zqkLyGu0ipKB495QUlNMM2PsWZLV/hq9n5GOYSLB8UpT2YvHO5XefqWWfy
Iw0K5Ml/PzATmyoIDS89VVEEfBXfpPjkFsgnn6pVNhfAtdTIjs5CfaaxNS5p
QXcu6bKlt9n8I1WoB5IXAreHZFwFMb+MY3yWHBR44BKEW4AVn0grPZfvKJ7E
xMRH7XZzMkaiee89cVH0qE9Suoi/yqEcD4hFy0rDJ1TSJVXu9L7W1MTCvNAs
Y9Z556Fw7Ni78ML1Q/ggUK89xYxLkQ4bWOgisR/4SXabiFFIg+TLmiedT29J
9Xnl0DPuEBJCThUqk1wWwMM9X6GN2ysnG5T66/+W5PDbSSSIgVZcILw1p/mK
nLKeiGcJBnbuv0U2ZFfQkt/jlJtvpGOxk7AsV859N7L+eWAkZWrbtDTcFtHW
NXSylZBbX8NaVwvB+2nXO/+/77ByRsJyVggCEsNssJ8M9PG793hEyuMgjIwl
n5wspWrdGCpEVqwMlzISHdDYi0Ptff+KSHp3w44cHcjr58Xotr0Pw/TZBds8
V4CU9UnTWu+k2JIwRbtD7LWwnbEFhV09WZZifAftslq5z7RxrNHPSU0dWh+n
yy85L5bVr1t3r8nYNCYCGH9HIVIoTBjxBosv6PkTRYsBMIoH/KJG+7NJ9LJw
rq3+lyKWTrdQ+DVVYwePPdhqWi9eVfFWk53K5zrDf85ji54VbjcU9BTtgMWx
o9YTsGtMpjTyRLeTpNoi1Xa67DE4zFpv7IdZvEqQJK17XpLuWtbAO6tSl6jb
+yO9551ZBU2jWmw6mtY8katEIH23ZZOTrtbH7IxCPctXIYJ6V9Sw6XxvxLQX
THpUpafZh8mQnrOreAexEfmAvphCaXXeHA2ZeyMZL8pKTwyj5eiOM1uss+S1
pKLssTrsXNabJjECXQFx7/E+VMyGKRYsiQUqN1lXwPncm7tTp7inLhVmBSh6
QrwZ+lNghqesVIlCqi+Pz6mw8+2i6dVfsYk0QrkHFaf42qAJqXazDQ9EckbK
sdkT/EUznmFLUe6rLI4qByBe3RqvRHiVdfa5HFX7OEV3CiSh3H2bmsU8qMPd
USkhFXT3VlGmHKsRp6rEBH0ewyxeBeFzgvb2PiOHPOQPWkqByexAHN92sYtR
w4K/hA+VMLp46Ow/7KBce/E9VHOsAK6reNjCof64HGf5CmVSlFVccZEh9Oip
XwpTtAVNqnxs98AP1PPYqkxAnMA5dse5XRQkuFJ6vRu3EFFbYOLR6fn7uVTt
MrMkg7yfvfVGZZ7o2iFh0NeRgnYh8n/NST/wzDS2g75f8NRi6RFWS6xtVsGp
6ArmLa97wooFtoAXJ0PtBH6n09hxnSuOr0smhINmDv1u2TVVXMRnD/ld2btN
glLmL/5s9kuOj2hX/BwVw/VkVeebiES7K8LUwpzKNJ3DCUnZjd0hMjggaLti
tb27oGTUhzKkYljlFSIK8lu5cKKaTrgBr1HaXOQgFetJkP4P6h5dL5To7/wi
eqkn1jEb7EXMEzFZxDJ64SECPgW3/GAfsXBsu1o0yE1cF1Ct4l36UIflYg77
1y9t2JZLYfm7NFU+6t4SIq5tjqsrcX6l0MwZxgB7HHvKmx96ZZpDj5uaU2jL
FOYsz0ngDCOK29KPDl4v77yBnqXsglI53QGgXk1VUsC8vBdZwu09eGZZ5xhS
X/LkLdEAGjG4CNVfGoeu7Z59uBHSmxUlft1inA6YBe65RyRdz9GBhlEnKiLT
9UoFv9PLBK39Q3IDrenuv0xDjLh/dDVxMO9Ywg1ej1FcP97RMsWzqcpqz8RR
62g8pDmL/XmbZ427x9xgbYDZrwu57a/+Eb9qDMFCXPphHV2CDxMOObkTMnYb
BPR+UXAyD2ciEHm/WOYI80CHkj6g0RdVlDP3mhHTmE0Fwlm2JZsYuIzA/LPo
LCs7iUJCAxGrlIDLKaJ0NKA/tCa4ytbWjC7IyEJz05a4cCqGBiA2z08JrW1G
018XeXSJN18hawp2TVjTAtnBEul0C1QgOvqTeiEAVJaDNSb0RoMNwFiKHvHF
wRxk96kLtIuLtsd27LQk95U8i4e3XXJwpJbpZb8xxUUSUPf/yP7TPd33/1Vc
NgzWWOfLwi1two3tFQ8dDp4JhNXVYo6kSZoZA/iih3k43Vt1GTv5uYf2LD17
HvXata+/oDbtwsON3HuM2q4lP9bpLT3w1fkDzd1Z5XpEhHP9WHXQKkDHRG04
atnScxzXeZYyzGNxbgGWzCqqg9IZz5CXyfx5rwRWT6qQZflXU1q/Je6qB4CE
gc/5k8fd/3I3QlOY4L1123w53zHwKXMGOfiimENQ9YYgkGUnO7MvVIXU2SjT
cfbVFBN9ZbxovdmL9EFaZKqdrpQ1TMml0mhjRFyQSP07afLMbC03FmjIVMZ1
QCixht3WGao3D6WAOkuFUvlMt5Hbxi+qa/+/hgZ9j9lNQBbf9XQ6pCl/axTU
UOZLVj6m3jIjmGxP94/fIADl/xZSP9EKbHEw3fftIpTSmClby5zQuaA1yRne
+GKfwHnScIY+oXRFcStP3ebf72NN98GqgDtsbyjThSJV8KLTMnZqPuLeD2Df
HR001xXjo9F4z8Al9anzJ/jdtcgAk+zPfo1RBvutZH1TFirnqr2+Zi342ECx
PixHEX93vJ47MN0ebh7yFwwx87j1WgiJIIIRCi1yvar8gfuifAQaCDCmlciN
QxX7bIqBf4j5tnaRVVo4voJ/IoLSuoL13U7hv1oFT0MAjcZCALzhDfIhN+un
/c2bCKwIgMCrGYgkbRUjXi9D4St2kx1Oo+USuwFnXvfMPjC73IZaxg4VGo6B
oj+z83q8z/sNDFzpkG7LGnmODlFdssRZH3++eNU1HKD3Yl0ybRl5dXfEAVMv
AR44sS2cOcFMKqvX2O2qN07FpKj6jlZi0aWv98Tn07PuqXPBmG5LdkSiYb4h
H8tmgsvSDOaE9RmhIIULaYSUUJZNjO9gi6ngJ+KGaH19GDzmFDHBrkBIE2FG
LXPoM66bJTege44Y36AiFypsD3OX/xYJO9PfpVgR9e10da6Bb4YBcqDwjuzH
AKuFw8p+hjsR8b9Q8zdTu2wDjiwdqJ6yOIcudLCcew/WlbUsMMO9qHg9oVrw
2WMSpqbmaBcaWrWutSgHUiKkRiEu7sIB+Fb4DILD1yUVvea9WAZDKjtXRDNM
Jf3lbDwf3uprT1Y/EgvaqO085h+gERcXZTtZr7p321Mq+WRgF1h/nRHowfUO
3tfgAONOtBK50AGvTTXQZ2k4xPsDs9XH5b1Q31HC+3ifRSi4BJ/Pug50yizr
bBh32UR55f2r52RhXUpEXHrUWXoDeV+WWFxgeQYPoVL+z+xePnBHZv9lEtDh
4G+qk0mDb2Ixo/1WwTqCR/5EvdKiysNV2MvcTHKN9ZynNNexFbNUFlayUybG
Qi5I6kAItqMndbpt0R3uGeaRQOaYGvesn+0bXg2lcBmSn1j2R+anUTIaZgYO
6aay7HBSsxkGuFkuZcAc6Fn9E3W7gv3DBdZyucXXGPh6DdUdc9xKV4ZXHckh
x7/ygVCw9sOjktPmoH8l9hmffos+ssXIG7YUMksflLDSleznjt++g0gkhTmG
3V0Uql4HbTqlDft3vg/817CY6Szgy6hsjotB5H0CMn9l3sr8VouidkJcHmWo
FE1Wq5p4YUzg5gpID8IPG1K1sVTdA8WC2Mcd/h9+L9do8U+Q5r9Gwj3Pa5p3
X44Y7STcyE5H5ZlzrfEa7F/zTK5n/wHyklNzBK9vpSnuOkw8xUO4O4pFP1r3
91iAlXmtnqqCOC1yWYLyxvda03D7OvizCb9K9NXi5ssW9aDqRHj3eFzOFHwD
rOAsYj3N6xpl7Cl5Pd7sgOwX+kEE8EagElx/0gaW3dzBN+7ytHgeDCtdJ8+4
BuYe+Iqw7XABvb1AurpcT4ZwWN8FT7S3YMxouvuMJSd4YrDsquFmcSaA72RO
+Zn/qmLNNzgsnfnHuStsPCaC0jFjuhxQ50+W4JW4+ZDarpX73/yCudWivr+U
MP6fHzdPnVUgRl6GBnWaYFrei4LcncR2oydmD6TGnZvjp5cDtcx2QQYjubYI
9xANOWBFqOZf96wveLFqtlfyILfoLLFIBgciSrvIEewyWnKXqlX1mHjSGLc7
rcNv+WJJXbEqrmmNRc7No0D2SZbPD7QzSIKM1+e8P721Ot+b/Iqze6VbEXz7
ir85IdrMC7BDkLGqTy0X2CFfOWJ2in/Kdaz5enWcKfAm5Me7LQrZWbeaIdHu
IhuL/Z9IiE20Vlral3DCTecqPgLFH4DucTMZ6AOd6tcED9EK6iG5lwT3vf9V
iu0ddfDOK6iFcdHRJaJI1aM35eKJ6zTFnymuELI4nj7UVPsuwYYFTV2zJ2Im
aHGur8mwonrW0WXZW0zZ/yGoBv8dltZev6ewe4w73uDmb2M5uc3bTIbz5Rnc
rru1hIQGaeEX6BEI9r8SnqP2dCJcE7wCfVpGGJN3QrMhj6M4GFDc9ItfZ/H4
Ls+uUCX8aquLXCzwmmdk2dek8RhUC1Xl/2H1E61iQDc0TrV1zFjSity5DCHi
/KvnXygluThxHicFqyyLnfHOe9JOmvz2tQdhuZW3I4G+DxQ0FsWLIxCnMZUQ
k7l6nS/FhYqalzaDuQtxSv7/7O89z3FZ23R5SQcUqSLdBGibnAZqxIVGgoWs
BYpQs79N5qp7J1Tm45e4ZjhDNB1sGtZq0g8UgQZhVNdibvW69fhRKKgST5wr
YX0uoQi68OToUVcUJpQsslBwsTupYi/QtcKXHa+4ODl3/x2xBbMHjB3d7YAF
B7eKRy8Y3V0ARlgq4whEyUOG3CHgJbKmEk3NZAzKkbJjX1r18+FbNON08qiS
jqBHMfplH9qluaXcsWFDyxSXeUKBdoiOl7aTY7VjdRaMTSosENRkGtWwEQ30
6Tkrmja9KpGPew13zdeN/v6/RPRCMlsoeKKPrSSmU8HwWceevnYP21Y6KMJP
lqb31oWrpXS3bKQfXWuDEpNCYk59S4ZsrUHA1SikCHllGMPXAj5f7TrqTIiX
94+5mjU45CbKfGrEp4PYiEi6KW3ksp/rA7Wa4WbyUJyFhtnN8sRal39zG8mo
7YkilylxjW6UjyuVkTseDjRs/SaXr5ebqtwpshzUuQGYGxdRzpyJ71eIFEVP
xazRhT3NydNwBVJr+VGd5ykDLPNW+XPnL9yJSSVZhyhQB0Jw9eXMWJeoiMbj
i0dT/QhriodbU4uIckB0uMWVw/Co4beB1iDPMv7DPXWN7kzNki/pnDk4rM1r
199ulX7ht3VvJDhc1b1Ka2/N/Skb0+nv4zSnGlb/RcmH6Hg48vzehO2ps0vR
cZ3e6JPHGaP83m6Y7ltL4ZiMLgWHndzZaSpfOHY90KdO/8+RIJOjtItAjKiY
rwLCjnb/XFX127Kpl3JXg07+Xp5Yeoh/OWJCU5NskAqYsdnb23VwVT/Xd+fY
DcnKGxvzf1MZKSs+QCjj+Ac7XE5Dje7ODLkAL8AH8I2hEpUUdo6kk7WNfgWS
DvafMuftfpcfQ0xXIV34va3Bao12Fm2/7FnDqcH2uUma6lBkFSoL4pM+IBC1
I+WMBqFqIl4E8/f39d9B2d8OP/f758189zo2bou7Bz8hnTsL6snrokz8ukBD
Z5Lw73byjOeX+rL5TPjaKCApWD25xY+S8qy8LOxEjClb239hsCksSwN4KzaU
S/F/03EpfQmU38Ucg5gtI2q0WprNSMFCEGP311+GCYqtFFoWQ26cFPXAeIbP
9JEQUjSWTVib5n7c8Yq3eVEf0shHQ7WnekW32gMvSBH5cMFSUMeBHSIu7cuM
vFUsVhWIGude2LJoqS/JLm3rjDCDQvGiInPHL+BGM+qoT2vTVY1BVmjZMCNh
b3lTepNCsQ4SZ6WfeCy9QDzpCSC6r4y2/OG8yVKKBAhfBnqZsY5W48/M8Gzd
ZGIeaeUkOp6Yzsi+THz9EzWNKSy7AUQ5pWC1W88VParlDCXjO+a3vzJj+J6i
6soVdfwj3hFG4Ps+JaYKlR+zQZ6IG6A4pRbcETvPQU02A8PM+v19ABxzYMwn
raLpJrf3RjDfAYcwkhVGNDR7fOaHOl2G31uHM7UycSLFFFG71zGpDuofNVhj
nIwmon7XqU17qQMQrULF7sozFKKqTGq6+dzUATlxDVybRb+/PsoK+414LhKC
BGuwK19wZxG2SZ/NEX7PQo+5y1O70LE1saiVrE6at/md1oM/8C3tKK/RkYSW
ddC8DQRw4Fykz2ycYiHOV1s/TY0ZKQ3QdnquZzu2Dj43EBeu5Qg3J2uGmLY9
YmH45130fBBmMdoCGuVrxfRyOdoJAYk4lDDm5SqQFPlFL+seEKPweowNAVhr
5/LpoWD8GC+Ri+V56lIQs+nFpnuDZsX9ChMYeNLeivLp8K8w2uY2wyB2mpz4
zWAANiC+xcy+2Es2r4RM1PH6PdPG1+dUaMEZ2YElXCeTLYQ3HzAJXFaHTvzE
QFDTAUDdixC8LwA/eO0BMgatqflH0S7xLEGltUckmZ2K9I4eQRMfAXiQOaBv
k5r0bcI7GOek8qaOwZGKEYUgQSQVUWsxwRjoLHvGp75RMcJnkKCj4ogvX1Cd
yQtkazBMazJzoPQhBc6k4r0m1qALEoP0tBW/vm/Qp+G1yQ/hJ6cN5Szv8DKL
vKyrhLfOlTamG/RROgLMVH4NK1yLVd1ian2UxG15vplBXfZUxGOYyT10Nuct
PnOXK1waIIXTcAd3GHHh8oNHqExi0XL9qbZe2tI2r6QRTowuMAuTEIeuaZds
BNi0+UP6WaIYSs2ScTMqtXUS0nbwE80brCZA6mCAQA1O9pGlJs2Gqmc8qAx0
7mUrEHwqLNcnF6xxzYxmH5nPOVo33QZpD9gU6b6LJyWfb4RYTx3kiKJqWDIn
Nq1E33Sk6qFKm4prpASemGVr3dQ9uwzQSUDILyTRvLrz9aXMsEA+UFSe6whR
IiPVDiF3lNXd4JbdFYrO6IsKqWdMLB8zVrZbl56ytYAP7OvsOhKYG7OEYsP2
c83NJ3bN0qJ3XZz0MGQIx9eQt4rGJu/qMsNWgqOy8wTHB8+xKW3akifLqzeE
tVtS501l1SNrN9qNANX29u8oVj8IZFOBSMG0D5XuIQMKu+6CrHNYGZMTBdja
clhnFmD0JepXqodhWMwcESIhMn27zZxoaNvuZRG9mWr37zmgHOomLWpD9Ssk
Jb5snJ3LyP8ygQOJsIm4y2+XikD/jfQcrFv2m/vBjw4nzFjdLX8ys7ukm9eS
TBXT49O/PU1AIlUykti0ImxTDlu6PcbnWHM7yDQ5LOWeIqBkqaPP+td96ZeJ
zpkfxikL+tylOOds0LXvavfbFliYPulFuAdxmSyo9jSaWEJND9f7y2YsY7gU
I3IKJ/gEqPlgUhJfc/WgsOL+Z/c+tqHd+i37z6fvDvlraSmE6KOsmSkj9Ba2
XhA6XdyylqUjQfo9WINJnYHJUAEgY29xZdFGUnIfCk9bFx3BscWt3fZRm39v
c3l1d9XhaiQaYm9xCWwyLyZzwq5yjsLpmc1nzYzaJ6v8PBYB8juWzbrE9R1h
X2EYt1sZImMi4uUh1x1Zjs7b8CxqmJMeQFjf68vLZOa+XaDeFLUZQzxKhhd2
pOjpl137y6SZ+bcYw1U+8KjJ7UQH6jE7Ov6qCrEVThcnTxIYucx4cQPz1gjO
QLWkiTTEYYeHrRMOVUVZwJ7/lk3jikNQjN2A50XGDgku5VrCjo0RmzYjemPw
Q7X+Yrm5aoNpVWZF6PWwwRVCdqZk3I9MW+zTcF/PCXQqR58F3K4J2CXSvRVs
jGTcI4yIl5W4fQSElpQw7qWtzKFQels67U3lYR39PazCdb/NajdtqUt54rwx
aN2J+ZiXtVLYrxgko//2M4x2o+prq0krugsSy7SLTp981DuV9WCd/WUvCv93
iCrHiydxwxDtADiwy/BQbUXX7EC5CFX/th/sj1AzsO47PKvJUtVKdSmGyS01
8vY3eMV0uU0srtexqB7GRkKDzRCpeW4m+SmT1D1K0hVLK/mCBVOygZf6ozwx
NJGpq0gQQcHZWG/8BLyxmi2Tdot0CD6JydorpYYGVToDDZU16s5yfGESZBdR
T60DDe23+WDexTf/JvZPgEK6hKM1QOXkkSSXJBw+PyFxdmb5Pt8pw1dJ493h
sWqSpTijuAJdaiGU3r6f6+zNgSm7gZveS6ixCZZfsR+lVKsExqfnSjaBrH35
nQujLHZBrHG8jMx/zuYKXbSU5CC2HkRIBWz9PiHoqTNYwX57aNWIrkUX9CMd
mI5xfimW3uNExlO1DlM+fYtt2/v9gS0b5aFqeYwYNrLU0n2BuRsh+CJavxfb
+M8oxIj6MwA/4CH3q8ipxhKaWoytBZEFtu6MiIu6h8byv9ZjQ0Uc6K7yd0zI
fXBs5HBs9cnlvT18x4Q5OMafWh+Np6CkwXfQlFG67KgGnjvyEWwP3xaZsLYm
KokGVo2DZ2rWd0NPRFVddsrymNsPbvydbw01UbUITXL9GB6+k/iitEXfemnN
aWMr6b5V4ocIOe2cskPMgy0ihBoEAjsHI2JgJnmQrjcRjVXF+6N33IQ2dyqt
yCLNPXqXsrMn78P5y+qBVQs5OU2KLzB6+GopBddhkeDIb0LjZyvI3Z+SkzH+
PEftt+s8yNrRCfpvuOol58+kgZiXUgYUFD8UL8NZo4VALNl3fxCrzm9HcCDM
bc4qis9gxQk9YxBYorH316vQWLrCtdJQ/lxqw2sxI+4NbrCLSg/G8O7r8KH6
P3XGcuy/KVT6XvBkCF320jFb2b/qe5mtottFA0uPKRLDWtgDU8dRLZb5lUMc
rvLI21EsaVrVcN1oWGJUnOIGnllOFIVNcwl33D3LmscZcDi3xxHhdDmnqGaq
mOEViNAa75ynpft99EqtUGShlWaBVZ6+rvaSgFUbSno1wPzlUJEzIujQMn28
3Gw9PP92hUzqvGDZjtAleEaks3n9/wsouNddQcovOLYkc/0X28eBPhMXcUow
XwPcF0ikk5y1w7JIu2xb3huABn+nkSUO1ge16SZf8KdACammWPIavULzmoa6
C/xMrX8WS4g+sEtRy1P+uNubD9QRuRJv9KS1cGPjXEMhXDbG/WFPiVboCWVy
Awv+cypZBwaDRQvHJ2CMIRm9rXPkPaWc1gxAu1qLcECBDm0cNjlQRryDz57s
lDbesfdzhujE0arCpWp5YQOsdyFSvw4T0EjkizIt1yrhMnQb59Kv4JBxe8wj
FA5PYMzxU72EQTPesvyatMWfEfgrl8t5QuoVRHLrrUqWpf+C9hROb1lDL1dp
B0w8x84wfnurVHaH2Akq4plUMN7zDypKXDuleo18HdHTWohhv5QO5QHwMRZS
O2/IyKasljSY5+Xic7wGCJVK0VMtCJRZ5GOE94VAm9+V41Iby02AoCex2fec
PU7S5sdQyYHJmX3hNX2Z2kdOIH/kWDf3G3nK7nNgYlVQK1czYbzU4546PXo1
7M/Ed3Ktot6P+vsWp6vZP+NoH79328EWfshAAKqzkZc8y2lkS4LqRdgFAnCk
EabNkh+2o8lQFr5ax5rn/zeE7NlqlVSELuYf9nT1vcwokALt1teqolSjcYWf
HOGhxUDKeeH9jekiwNLSlbXHfQbkHNDwgO/uCQXofk+/Ah4Qy5DwZYwbjWlv
KfBLSv6TTyrrbKBK/PrMGyfoxa5FZaBTfNXS7tGvZcQoh2lttsNSFSVsS4oZ
OsMB4pn4Cae5Owy2MclL2AU9NXMTn+mHAFKz2XdGpiVbY3PwWTwHrn8vb5hg
4P6O/YYym7G6f5H7pwRUJiitS8G0OZV2ktjQJK1MFQmEZeLLJDGHN+OHWgzC
aQhDI5mpOaYkkzuoNJXwLHXIwDSsxi2nh4md0bBrPReZbNn/HhqUt9aE30Xx
ukaRiSmaniJ4x3Rkh8H7TVowTN2U/ofDZb1SWNFNZOfO8jirk45kg3352r7q
8lvXcvYM05BF3LiTKCXoc2guNZl3jBPutr/5/99t7uyaccR176cmkFuvvGut
yC+/kW8qrJiQzBBuvU+NMwvIDkb8wSMs1dbXzNlKD/JvJJ9ugrURHjOofZaD
AWefTJEE7DjVGurmSdn/eAdcxjNag0BVjvz817zNhBGzNu9Zu/qKQpeYpEQJ
Hm4KtFmxNuDOQ4yisNhq8f5IQwrT50x6nHDjU9PVQjGq9xYbEa/m4/o0X4Uk
rN4OdiLYi48WNc1Mhw1L3KIJsa0nfDjHqrdcKaMBjAIKoE/XEFPdI1Xp4chG
N7CyiRd9kT6JS45kNZx8AcIyd5lEV4pecc/vNWLN00HNfZtK/fsGZkVuuub7
ROy6TRsfYvPiSWe3N9m9J3MXUZ8vcdGPudPrNnjJqix9ZTXoxNqoKjfYzcfe
pwDUIv+vEn/DGY6HteSA7NyctjIucZ1hdgvvjI8YkSE05yehFXn6V3PYb9nU
Z2xirJiIBux6xCo8W8cWaktYOoXJK35NBJQWjbZRwtwZZWmcSlqtqGLAPdLu
dG6YTIuV8uyXJ3sHWGXfGqdvAXBF52wIdz2KvZbO/Rb48jQxKlD0BRzaeasr
41lbCfxgznWPzEbWLB0DJAL2+R/pThrt0wNGhzHUJzoFSpYW2Zx+YNLyGG22
r0AGxGCZBbbVPiE5kqHaEmLWQUnD5UK8mO/o3w1VxPLygMS6XYGkSl8oS4yc
FQ3PZZOFjBbCwVtVl0cPLOnGn0MC0pRWcyBDr6lqJxuPLGjse6q/Yzc2rvX3
xPHeO5+j8NXR4qoU68rzm3jbdBggxypl1kX7dFfXamQ6eKKbvN/xXD+o13cV
9O7zHsR4ldm3YteNbfKCJz0JXZSLOUDCB8mEGWJ9kQNT4to/yKoRdaNtRDhe
ofP8cAGqme7M9Ganr6ciONbTYVbGHNK/TypwhCeoVEsWR594cP2l0m5Beq7q
RaYFauBKDP+JVTRhRwyxWFome0Oh5Jwfc8feMlnMtSfXurYYm0+jR0N4cht6
iK3v48nOGZUgCKfXiCIB/dgCaDOcipLtwoy13jSnhztekxHgVNjQhb/pkZum
Qqj7z0UgBu8OWWaBIKe3TvxwhngT2JSbjrukJi5XyDw+bleGVbsTBxXXCSOf
dr9leKms6w7b4k7ZcTyTp2hhI/DMq7ha7uTqDGjvUhAWUETkRxXyT2tyq1FE
Z4Zq8Pk6wnkEJTIKvu9+c1q/PVx/ckRlJKVaiILbxegCUgOP8ZVYg95YeVYi
sp8o7SkIHlfDMJ9C9SPzUHsKelTL2g3w7FmrsOKzVVtxznhg80xXXS8/LXTF
6BXqeFIcSB7v3B1Haslzn/Nma1sPMYNldJKf+e96Q4JPb48MQqlKbDr62lG1
GxtapVIgJfwbelSqFBR5WDGWWkcToC83Rqkh8+/UMcXLsN7YHybhAv3rIs66
xrkHV1F/BOJSghSIl0qB8TCF8ohIUmY5Pn4zxQEI675336c4tQxev54/ewdv
RihphxZeeCeOr0YbPCb5PwC/cJedRMk3bdZ4+MncsypKweRPG/Brnleev7rc
0knvCc7wjb3VSBxnIJ6AtDzcgdF0hgw+qVDEgdQQ9+cVw3Se+3G/e7acebDA
nDeJbQLk2gbjXLSBbgMVjsvuJf05nJ6NeomvwRV44ngsxsb7lxOtzmsUYRKp
nHadBVpKNEf2yoZ8DeC0pQHrJHKLcIkQZifJKCHo7GWyBrxeKM+C45CLErFu
iu3FX8HbY4zlP7Kd9+o+G63jvRRYJvdzro9zoX/e39R/LKnnX9bTDwZ9E8hK
tE1QWXXa5l8maQZYhJBx4suhTeSi158lXYtnauqj3VazaLzuV2c2WeJ2qrTk
CwiDRIsxqM7sLF5zEl29Fe8Q7l1s9YO9yF1jr9QY7CfDyPKz/kEVlSNYnppq
Txwu4iTev5i7mxJ+IfXqgGNBJp37cbvlEkrhWBOwnPgNfiVrc6gG5FioyeML
7Xj5Bkn8Lesi3LnOwVkkY3ClCOiI2ZYn+VLz/3JGGYTqN87kRVPWpUOqJLlj
deyGBAMrOrFjCFRP1qTO1xlvov61flc4Q6NKRhBBSamN1vHwX0P35FRnCnjC
GnEHFczKSjmkotRa1xsN5V8N9ov2QMB+MjQgJMYdH/0Nz8Hoi4hRbImsDzxg
/7eZO+9WwRb23HXqrxwxUiIF6ePr3aCx/L/SKKElBmnkkh60tUZR3nMHP5UI
w99XnNXqjQqawmdytUzl7Ltlwp751pkMje0luYA+XTH1UESnbWlYceyH5iUA
YQBeGBw9bQJfUltm9KTuqUFO4FxtLNoksnWdZitR0vcsitkvsVDD86d8Dr9I
VVoECTOvEeqopM3ljDnFINmGAHmXbXn/2p36PZ5cypOCmmjkh8FzY6u2PwhD
OFhxJJSQu3QOZIllGUo8vX9DrggMYTevQQBHzqmNMzGSJl+a0CcYctyChbcs
iJZNO8AtoRiF9XO67CVEtI5NvTBrPmIGhn3KopDHB3aSk6TbHh4ZgqBPaCzh
Xk+Miu/bM6TrT4IOhCACq2RCgrfIYH7myeoTBRfmpFQpUEji4Y13qtbhoc9G
2+dTkAb+IoqBFBJuTn+GsPzwlino0h/0QUGr9OYiH+2GcLfaHps5abu9cXtD
Lm201Hth73jOmWHs4VLU6vIp9UMsaueUO8NKMnwnTHdiCjAbUwqm7lbvQTrQ
KYuUucVpQ/+gj6pCBL7T1nFQT8Mkq3v0UPQZXBRAzqEhff+ZcETHDXgjafwG
8Cmax1I9fqhgrNCDdvPPDzgiF14X9vxlGNF7YBM3L5u5Zt01KTFjMT4y0PvZ
ZaepSEazy+Rz+IQE2V9/UcWgZhmP0nK3iL4HqxTJyubP0KbJUU99npp//lAm
wrvl4ZloyxyqtEGfbhEQmP/MdRg9bwZ9BqrLI6I+199Op1PzWhH/1R7Nuq4J
t28mREUt4efOmJF6uO6h9CM17fG6qrhBLi+gbk/3FegFMgLPPPuKbKrQxcFA
UPcWk7IpPwg1fKyJbgrdjs2F+6BqnB8TcuCkPC7onK8tTgeMkr7RYtW7RXzP
rcTB/pY1er7KztGRsuR5US2G3UviyPR97VzKFpyt8xhNA5sd0sF1I/uVZE2D
Qumfv1M83gkYZz/8WiLFZxzQllVTJ/ACA0T/juBTuYmfIWwHSD61zb7a/hwU
eJUKcxlCBwEtPQO9vP58Vt2v52edcSr8k1NwcCoD7VgkRlqp81D+Lb9O62HI
GSUPGgZx94Bc1ALpLBcROdCpfyiE1f9WyhAXobUfzB+M3mhz8BJEReskx0NH
RRad0SsrWJtc0Xow0mJjnj+Q+VBTCaPQy2O1kpDx3ey1B3QefDid0BcVJhsu
xyo0LQTxzxP+VLsKm9KQUAoBm5V1cjscgd6SmB2r3Xfwo1u2w7qrvfzDrn7F
m3EdSom9YDYR3qK+1jy4h/yYx/bu6bWJ6ON8VcfTPdrJ1sFreS/9E56RDdBb
vA1EGFJrxaMx4I06VGlNsLQrzkxDIzX7HPhKbQJozpr/Lije/0gmO8K6X6uY
dFXJPOTzbyP77pY4FiikBrpMMxXP7f5lhjCZMWB5Q7sFJJPgbprWKBijj+14
gJ+0D1gsZY11a6QS4axsbsoxm6s64EeM081w1vFDLeAVM1L6DDCbZXMQG/sQ
VfAvDxrJ8eQMr2M1pz5p6kRb+GFNa5+9F4ISu3G8wawjorQmuSREb2PN2FEy
3WtRuyfTVIVru9u+RPMJtMowrz3jhBpbK5J2GvlTplX4maKzynwxgKZqF7MN
rKdEVV+nHYf/6tsXPfTtOb+j6gsqxyxjwxL808sqM+Sc3P/Ae5Gj1DZqoO/W
vQ1Z1jIxgWLA21jHDxk4NozRsEPUgy8/BFx4BLWuB6AXuOvwfzXyBvDniKCc
n9iAe9ABhvqq7Bz7DSrt0CbS2OS06a9bLmHT0yIZXbWvB4/bN1r93MTeLgq3
ghF0Y0yIkpJgHzhEZOaVVQqBGH88A/o549hyxAmKJVhrM1WMPsHAQC1zIBCY
HOiOfGVBJ2gCEHPHtNa7kV0ZdEhkKERy/gOKdJ/2Q79OAv12jq/3OR+rDS/A
LnNgGmQhNzy/d/z5BLLWPHseCYho/othm47uiZUeM0bx0tc77T+AG920luRM
D/FxbxDIBlarZsWU1bZAi6R2kFAAZG0Tx4WG/MonY8IoPMR5Rr0dZdvV3461
gpwKrbOhR+tqRr+2L8HW7Beo3tYTqHBEGsEMJMSUqlc3bzN7L7zgLKx094D2
vgGc+DaTY1ESUC8lxYy+TEY3A4BrsseyP75X/3KnrsjV9dFxwNcPN7V5PUII
Vfx3VT9W64dT2mgEs6dsUGVMKtbc1SicsVwZ/GL+6wav1G+63LVbieKCVSUJ
q+eVdDWEPpnn3GAajtSvPTc16FwoLRFxQE27+YgpXpedtiFOgSRaPbBQ7YUR
zZ3h177TpGZUbD+53IQfaVGgf4zGAZd0RMN7msoA6236QQpeStawl+ETp3Gt
uLd7a76+COE8TonKsQhSGkDNmhZmnyxlJrKXE2Itlc7cNASuukW83rckE7I1
X71KTrFzL6A4z1eCPhLXs1q4iY8wiOLIQsAVoC2GE6K2WSf1/zp5bnvct1nj
tIqdpKrxxk8rJ18lGJ1IfmIrV5S6n1p8FLuJV6gvTutFDaWWV94gQ9ySVoAc
5v+JtfcdoN9ByZV72hrFa911xapTKXcZypml2lUPb8uwu2udxDMXdiEeaIch
5MQOCBPr1N9tkOVd5no1qPlwT21C5lAUxojmNXsclcMZvzpSxThw+fadkwGL
rdUWWWuOThUi+GTEmbHGBNEwOwSeI0K73VrTZi51eUG8ew53yMx/BNyO6noI
vln73/Pq8tTQyvlwbEx3sA/Lr0n+BPZ7lUaDpcC7OXzzeKShniQmD14sJRz6
CVpP0wyuiE/0WMw1vI55eBlZvnvcjKJXO0piNIPWGdBRngIu8w5NWtHBUjMZ
LKmhlejDhCi78QHRAf7fPPgrQF1EtDYjN4VzDZYe3CVNMI3h8gcsoaybjYtH
StbSERmoarxWR6ZsbsGuYQ90Q2FRP7MpU/bGvjOe0K80w65k1lgSluk2xunc
QmpRD0zDXt5T/RuGfB9r8L1pBgxSJBSCf9xgedTe2lstsGhSr0kr5V7W+Gh7
YWA6nFppfBtruOZ82jWprISfM0d5ylLQprausvySjFUbhQKOWfA+eMyzCRho
QiO6x9rDyXLhyKGMm9vuTbEIw3LZww+ptcP8hmFFc+URAI3QkHG5cENSKoXV
QaBKjeowZyWQFhCXSEIRmLhMuNLG2YhlElXL1PvRWqfkf6wJdYhznc7gwkvx
TeqEcCX1p/1o+sy3IJ7P6qCX18n3fok9SauOLgzFlrGWvX+SRJq69dEKM3Fj
xHQ0mOvSjjUvOIDhSeT3F7t1N2Tv9mfdc1B+aarffoHV3253ff2GF23mE113
lVwgBSPhkkGCD/GMVBf4vyAGSdJBAOOT9FXEdEfnV/zqeub7J9ZL82NoQcvr
3pZWXb94OgiVhWAd1+qW3f4s+NQYFew/LRqkxF0oNaZdWqwCUezW2cv6jjUI
1WY3OAxoyiBIJSqjWJypZGf8+D4j4UiB34IHoftsqLB7vMkWYXW69h8OZpgC
hZehgIckgUD/gGNqo8v1YM/kPChkrpgXD7oI1YNZmBI2NEhGZkaMeszx6IO2
l0A/M61u725w3e9J6rqI0Nuwi69kSLx0vxLdXSknv5I8KHZGI/QZznXhJfcm
G/SHzSuJWo7Fz1m4jxfGx3tdiBxZPxXY+ZVxdhN+6uxO7CpNHy/qeMX98xWb
Hm8+EMQMi4MelvZSPmyLSVK5Y1xB89YJuSvoVQhpOppHRhaB8qSFmUX6R8dS
qCUm5WBfHp4Q955maK6By5MB6T7lyIIbshgdIpxfaO/rwDiettv8AH3TETzF
hAsfpRmeLa0xsup1vq6j+U5wBx9GaAPTGOB3SmyB+LFYePAjrLzqml0KNT6m
ktgIQw+91W94LxyuJb7LpyqyRhiWJHtIkE7R2btX1HJLBjtZClUu/0MxrWwT
KGmK6X0Bfkom3B7boRoQFFb6TSJ89oEaKUm2XCenGNGdcW4IxZJaQPUpe3Ed
OUXN81dbAY/K6wd4lcEzc1ldc5kKSEHx9S6xlCrUV25yuDSthqHu8GHsZZX0
tCWho7HGHK5tP6kCXq4xuHZzOpN9QmdsDMOIoXuymXxTOCLy3GKkwwKP8xyn
z/q4ELrK0diOyoop223whCu4UE6TYazyByladi7UxCM4AX28/AeJuCCWyuj0
aRT3lG1xGLLmGSWsRbrIWEbrXictbqTYs3OOhCUoJNuLQ1ZBgnkhLJZXq6aZ
u6UwC603d92cjAJEfxHmSazEYnP15zsvDW6L9K0BcED8+akTrop86otGHzOI
jOCh6ae65utB00RsCPU692N1z7me/U9KKq5n4+JZXm9cMcf/6ySByecNuaUd
bMSTZxPqArWmZtwg4DMAnPRuJoz0hseSBbzep4E2enDcsXP6MoGq+ODo6wMs
B0WhBtuOOJoQjXlk9nw1DroTXOd6qzzC5APj+U5qsTCsF5lORvdmJF2MooyC
811D/dA/mc6bZbA+jSVi/uZmZLpZ2u13GRg18Z56TT9Wq1pD3iDmxBZIPLj0
6khAOJEV5oPmxTla9+YRYRpLlAkUEZVW410qs1DT6jD/oJ1zMnM+KIO4xeyZ
8Dj9EuBhLUw5EMuI74vadz/blH7r/onBVKn1K6qbj44NGKnbztFTR/ETDu5p
tq2UW0Lh/1SkXJ73nuL4X6prOL2GvKlLHLVqqPzzBIXkPSijUsdcPx6vk1mC
IN6RmixzGtt+f7NpTMwkMjTqp9BT2vYvTG+xvZtszT3o7g5gknArNKiKjfIX
CJknNnFm7nHf4naXYh4BB4PhOo7nt9Ggy6IB2s2q5y4z70IFzgzWbwiHzEfl
kjBO098gk0xnfRsUhz/tskr8LwrxTeoJy434F1ULX0s/ajbVJITsx3Ed4J8h
D60Mh4BDk0fIudygSafti/n1++d3xzjuNLCMgXUKl5swscCjO0TgqJjLQFuT
xc5il6t4CQf++QVqV3cK4QtkS8NFLMLhsERyX8TO2PioorQuCWp843bPMGXY
EUQKlJY41CsEJO4quVhw5aQdFmFHYckp4YPWKjA48vwKmDLkAPWHCpoFNCFy
ScGnHoWOjdJGRZPLxPn2JZjN83v/ycnhyE+EtiNdSf1+tDsBRc6OjXzgJ1yg
lYAfttxmB2E8PMOf5nvTgFfzzFOZUZ60+zY5IenBL47NbfAwkoz1jn8xe7H9
tARLMqHzH0UVr3c+e8zqxOpHsLL1Aq0McB0bnZ98WoEfWO6WMTy0YiGFpwct
sI8VmeOtgIrsZVFqEBkrOuBXT8fW4NQWmNfsHItdutkn3cKhxLVpTpfcIXPP
blg2Wk13JVBrsNWRsm52ptljp/a/Xz4W+m/uP6745h23QD5KncjN7dr3Dh+c
w2itCZJoI5DIDCdoWHe5sZ1fLL6olurHPUHpO7Z+2yzrdGqxNxMRlNv7wfL8
EKv1nXEyfytjA4+PsR1+e3TaJe29tYqyti15mNYRzUXlz8zeQmmqype/Sp3d
BCTqbUaXtN/5xUGb+smSpNIbTKJ/IGKb2yXJfqQqkvurFCsEK6CGVQ7BnKOI
+BEgrfwGhg4d0jvvZXI5Ak3vXAFZFHuXhzOWFPth1Sy+K3LykBjZGCKbOnV6
l8E43EdvDSb1vR9Qe2xKNU8RU6u1lP2ZDNH1mIIfP6srzg4nnBnkzR3CXT/r
pt4yX8PKXqWX0LHCdU52aWFICRF2BPiUs6JVDSVyaCOOXK5Z9EeN8nC3pFQ2
sI6GuFjFW+ysf6mpslJdp+ZvM4Wp6jWLkM2iscmBBZD6ehgi2msebqH+dLCO
4Rg18qpcL8Fud0I2/Q7Myut4fRlog7YC9PXH3kvHfSS71pvRro9G7OnTxAMh
kX4F1xvz8hi1UmERK+Z3FSWqKGbW++kP5ApYVGXh8qtjtbAj3Gh9qZ3Dka0i
cchgShqM2WDx7xKinnbSDfb5cVRrrJbuNwCvEGb6jjqqCcstS1LXESHV87Cn
oDKtn006toPbx2NFnsYbDNiHOSRzQtxCVqsM6MdUc2VquspINmiFEvVSdY6M
XfmvwcwoIrFKJydIO+oZwerQQIOxKKnDQrsQqkNI0RLpmppNHfHXq4UdOfxp
S7Wk3yKt58IXchC4h5osLBAP6B3y+q6YVmVFEGlbr9BZvcnVGYlpYE3KuwGq
I6YbMpjt85xycHLCk9NZ5l5cpKgLRf/qM1PpHM+76ltj9sZQ7IUdqSW0iZdD
9MSyvwXYhr87DVIVhvYV9iLNz1ZEgiUFxf/XFvM0xAmFYLBMwSB0HGDVScX6
k7l4dNuemwKom+ZW2SVFyhJd4kmTauPgmnS7O9KFVHLeEi8AA8+F3axyw3CP
glWp/8nKF8ZAWbyUJLu1t+Fz517QEVkOtaBdO8I9fG4hsYwAIFuEOq33R/E5
4XHfPTInfX81hHM/bdlSI2Ns1s1xk5k3fj+pbxBQn/v/sxgxpDGCpPvEoPuP
BczHlkM1wGCYzBIyfs3/0hTka3b3uznusej59Z+ub2knvFkjUzFdUG+qm5XJ
nX2NrdEMVhR7sfYOYbqVypilNMrV3G8BtqHoabWQkK3HGB4p2nYszP++TIlf
pOeOUx9dq+E94J/HH6pw4U/WPs2603/LV9fDPsF8ris/TQY9jO0GxeUWf2f9
8EszM6SJjzKabdniLaqdkv9QY9rLT4YMNsMaG9FMfduGsylZ9D3nft8zyQmI
ey6eeiERQrRQyRUxDmtYb5ApaV5F3Qn6g4MZsi1/pyKGvbY+cfc8ew/mshq7
t1mczSXxsy9f/PaG0merVRoGZIpLIcNzjobO9p47nJuWYU1fTRJoDEv+8MZq
Di/qKoBFWP1+Rv7TqVyRHBg8ElM5ldA5E2gnBz72Q4JJx9U/a+H07kft2JKM
5SOY46Bbxw8vUKpQURRXw3OJtGFAwzfEaPL3Lj1vMKgjVM3TXUohPoVv1PfR
ckpk7z5FBcrtBSkfguOQVYx2l9MO0fMH/+nvFW/L+MLauwg9LF0lddxUnclm
Vz8CRJF97Gc27feG+r3bVwmmRnuqhaxzjtV0zOo0yX7O+oF+dBwRNrF8sZaG
AIXunpb/F/2T7hMJdE+uIoH9VzRcLLKNYNFcuMT6xBd2M06D+98+qGK2r+mK
zZnWe8ExpIVCx1fyNiwx87i1O8rk0rindMoacECjMgTGdjJQL+mMKGoY78Xt
w33kgrU/Qljc1TnQglS/k+zsLL7DpYRRlB5mT3epNOqDrr7+ZPxYyefSJ2yF
ge8Q4j0Ic4NPDk0LZiXi8XRnGi78xFCjOGSOaNCSFx4H6JJ1feHnUFMjz+Xn
QrWSemuZQ4MCBs5qaJFQyKNWyTyLQpN+OUPqMBpzjPmuWVfjcNgbfDjIcIHW
TnFxKVRUm9vrXPNI9PSY7iV1WWRlHhFSCjg+EGz1iTnttg4Oi95llrg5/8p8
S4TjYAsvwteq7rW7qCbNrq5NFGZYWqdb7/NHhoMycRVxSFy4Q/AFmEMBPBIX
/V1MOe1pOJLInlK4EEbrEHS4YfirfvOn1bnJX1rS/vKK0u6+69zaqVUUsBeC
WtcQLoQ+3hZlX+p69A5sbzD/g+JLFTVCQboB115nF0UhT1tNQ/7L9Tkx2FmS
LniJnmC5EFKKVenh8gqPSn3KRJsYFg4uT07EwpdRqdRGn4v4Yf9yLKRCd+Qc
b7WPDwHXphlj331P5stGpQvWxWb497ddIAQwbX4QXcMgzhgVu/KUjspl8mYW
duuP2z7YsroF2ETJan3sXMrpF9r1W+QUadYOWKE/2LPHqSM1lOan1uH+ruA8
L4OI1xWEd5slKvPE12RXDxt3JZSc5Lixleb/NEKLELQtdOEMR5bsef7+CBbg
aqxmp5h+ddf2SqwyYPsHyjvo/6wumJGbJvg0Xep2D/tul76vH+cRb4Ev0uNe
hgrjg45EyiiNCDj9aRKdrEN9gWuqSej3Byyds8SoSBVys2uy8z7naFHobCGn
34RZXexGPP3ozvHGhNqzIvcd+jDuWrqWF9GSacOrJ9Td7YSRHHmFgSc91jpx
phy4z6d36ADQrIcCcgHsTeDlDLlaJcBlwCpW0IHpHqEMyV3M4YGnUJa+VeOl
tYOF3HeV8aKgggF3D4uAHhLUusRs3ees5B7FVL7seIOMaYkHLX5OZ7vv3eAn
SSlRn6y05LHJUIkMRk+RvHB3mmyP958IcPU01zK3x70tipRzDfQkmmBx/N4R
EcC+Sl7CYqDYWGJ2czuj3Nhs4KsZVyMN8e8HRyaifDOyU7bCpk3WfZMFC8NO
zw1E9r5fvNChmwtQlwZQzxRFUISy5gkfxtUEXCc2ok94MgluEHk8CGxbCeYC
X8XRlAm3eNYJmtz2aYnFglH3PxK4kEgJLKzeiRlqYBTFi4sla4g3KC3Tn2ga
zmpQq64S4kZoMWQljOtwdhinPvwRuzyBKyshsgm5Q0XjRxip49TIERzwmwor
PK9eY0jy2b/P+exEwXMu2aXvDXjpkJO8QhQor9WX0sPYxpKQg7eTUiiNudTB
3wIK/kyh9sAcqPqnCFd/FTAUTLAV+9bwHWkTT/veM4DLKLbtVDQ6hOcnAOL4
ctgrlaKuENudMe1thiAvETsgNCh4iDWzFY9xFMfvEtwyiQv30xGFStxM9v4A
ZNHHK6GJCAf+ywj+KSxS247h+UW6Kb464vXvO+wlIDkUeVlTBNHOahNShg6Y
XkKFEOIiZd0qscvC7iyGEIVtkFPEDoni4Zu9+2KDUkSCZS2YuKylYEiezARI
e/eGxCVf7V8PU6wzwQpd2Y1XtisDCDWZv/47NOkB8+P1qa7M1dJ0/fsZu/+A
wKW5jiKNZoq1e+KlHeHYeWCmOQVzJ+M5q5nJmuyaVDDILrqUwpjGEQRhliqS
Ta7I8dfyvGkIvchon/jSCdAqHabA2OoD1ue9HqKsY7IJ0DUAarebFgfycGTb
Y2ZhRQppVxUBm0XzYWCjN50w7R0PJxFCClriIlS/6Uqi1KYe7tMmF3mvw7f9
ACCEsTzvu5slASgcBvB/bYFbiJzc5WIfGy5XmeiBQjDR9jDwHf0qcvo6OyiY
Qhp3APPNegMEAOTWF637I0D0p1WRH1UVZCCpfiMX+C5BqaS/jpo4hp6taELQ
Z8vQxeAfQZ6/XRb2nnprmGGoLUcdGYBevN1+YGqa4bHJgeLRNaS48TlPPBZ0
fqh4PqInVMv2AVWaKuzGKl/9xiJORZccAwbzeTaE4+u18GsoG7KJoZh8FxJm
Htz4UkgmuVdmh924auG3Yk8y4If9ACa80uNo3C7YBExBt1VAnTXu3Vw0fjxV
q+3S62HV1qmKcMOoW8mU8OU/6+Gnjxfv22zg5MNJWQ/YcG7cbVNhZ1NFoWNx
QcvHE/wNNiwXEhkNcsNRBam4l9Jc0+r2/b84V1Q8BYUEVHHWP7i6u+X/VY0M
mpW8cSIubft9ejz0oTmiyhFvnszOJ9/rWLwROWj5LLpeZ9KiSa27HQSqMKeI
8hXAGTw7dl//2uljJpkoEUCNlUZq+nGvoSwg32CXM05YOCl0cX/ty110kmuu
isoWOpgI9NaLyuNLSfxGRzZPbcThpqWWObPXxRl1XeiX9us5CijhEWDR0hLq
eM4cYXNZ6KK1GJw2OzsNeVYNxy0jSqb+pCa19T3NGW4P92gyP4i5apYeL4D0
mK9UY5Wi0OpMRojQ52YYRU3Gb1ukMIY/Vi4zrEJchPfcOV16qOaXgOm8IfO2
yHX9LO51JmKPfbTz5Kmw7/6Qvb0JDNhxyMnc/BLG46L1IRECOa8h9n8sGkzL
gbNvo6JuuFKKts1iEIXW/MCJgxIxKgsGCVgFenC0tcHW4DDR0MWCscpOlV7Q
NguH52h/qoarSRfu9bO8F2Fa5cAWsFO3RGUz68PqNdm6dSQumQv/WVF3qVQW
3Kh/EUpAapBUSajWEm2khTanPjOmEfmKMASUaBr41KhNAKfdlHq31Xvowjmu
3qLd9W7rgdtZ9dOASxS9oteJ2eATmTldNpKSkO5Mj/DFEwFcy2PfE5Vul71Z
epwyIkRRAD5oLiu1sMfbvOQ4wghMkKIqOCypJQ3hr2er64Jnb5s+n55mVYuM
rvo+JEGhvMUc+2tn3ioDNPgKtBiYN5Mbuu/lg4/mkvQiOP3cMq47J/FXg29a
vKcshm11Z9ReCN+NqrTwMCYQAvZFHlA9wr+jK/jvk2SsYO818ApyixZJGeRt
PbtjNWV8ZU2XeK8CnOKlpbrrtXJNsytV6uavN/mbuOmj8aru/KnQTt09nEOT
LRmzorgkqU5I9lHLRjehfIsAFt9jMHHzBbBfs5xZTyCeTbr2Awd0gob1MUwV
xChAMz2EgDDOvDAVlDZ+TQYZvIVzrYrq3F4qiihMeZsrjwX6pJGLEMiy3904
aFjvsjepJ7O7Y5sVfHW1xYn6VxkJ7++Ly1n+LG4ZNIvqMdshQE8QBwKpGBK6
BR/G9DW7MHSvHHm1f3EGDwHHesfmGbU+m1Hgpg9GcE48TTEa126lWJnDCOzo
nhkDtE+PEKeqWAA97wXE+K3SsDKQCh5Wha9WbqDFuOAEsDAbECQtWsYKslvG
EJqpy0FmWQyaNuVrsioEj5a6t+sIFz4EHXxI0SYE2g6CsLp0/5T1QQjgbqfB
O1Uwo3cfMIW+6flZba+hHLn1tMAxCuOOLCuHvPKMENj2vKyeYvZttnMTMI57
W1pAiM9QYnPWTNNgmsG0qzOUrihrZ2znHimM4aeNf4QDvkFGsaBZdoG6ISpy
mQnmm/1SoQbHyfxZxJhivNyoUxwepPKqJ4MSpDxEJXLVm80VnQaAQGbI8J0y
YwY7yFUbYBfR6nTMvA7yoTzyU5GG/UlDakJtYDOBloLl+IloXAG6NeGmRni6
U4n7SpIFswN+sHjaFIN8VCJBpb4lfZZn4nUzBcTOUcuIjNAhGezf/qbk3A3V
zgb5YEQ+nV0ruV7TP8X4EtgJpvu53K5xSoyrZ2JHunrkO93178YcuvvNkO5Y
JUk+s+opgHjJ5ntaCBzJ40EnOubEpqqoFLbRdOxgH0qMMvP1bm6DLuhy4IU4
oyriIpUTPmv/IT6h6/T/jqY7qQU8s3IsjWgtCPmHxhh6HN24EYZoGEBvwGNS
QS1jeXryQ5RdTbSc3ONWB1PtzwbYRk+dKXQBJJymfKoOLZlWjAW8xEuyf2gD
gyFhsiqD1b2HmqnufjeHjuPadZqiWxh57Nl9zp+LF/3AAtcNwsIZMGF9Y/NF
HYvW0oKp64AXT+XbM2/ynVyfaQyATYZQeklapTfA8VVPrEQj5v5bTXytWHsf
tV8Ioo5DJyDK2iX/SsX/n6Kf1T7onAYVFY1D1AmyEe7IZsTYoTIjrly3rT7Y
8gj00AO49iIP/C1EbFL34W/DT+vL9MMvHXx3LNFs+wrVFXBlmPNk97dJXA/t
jLUz2jz3D7BwEO/vMw6S1/0skPxsCctcydRF68DkeY3XNctqLWDz9N6L+PA9
V94pLHbqpj5yPT3ptWeCsYuL4huayi3XjKDUZfrM4hnRTrKDv8uDTMhr5M5s
IJ345XySZIX0nVgxiuIa9MHPqaCY3iIy3sK4zCcrPVffizfC8jrxPC9myg9E
02dymYhPb/bztt4B0hDwN6asFZF61g8ohv6Y3u+Lq+FVxo53X8JIpSdWpUu7
+HacjGw3gcm8xhJuyrv4iLPpw2SSv/AhH7XV+ueV4FRw9jWEAA7Z4SrwPXAK
Jd7Q41TfXHeRJWqDlXhNWoux06d7BCLbgkMBvzqTA3mLjq8Ku7sTiBkn1lel
UJG7ysgoQtuP5iMjIV5ZvGPJN97vpZLXHKnBxk0P5RR/PxCfd5SvAT6nw8E0
TDU7C43oNK65bmrHC1NRPfX65wk/6g9abB16imAmu/Mbqv8aA0MIpW63UbXV
zgVtiSaUKtir1KbuJfQq4GrJQhjpDIeqp+xS0yYs4UmHKyLMzUYbX7eAiS5j
n4umsqYM5V/Pe3SN+9clEUZCClrPOruo9W6nljh4W3gGYrG2ubMJJ1fGq8QR
STq1Os6MpgLE+04FP/pAB/9kZ9elCVeHY2YtN4xCBVSp34S9315kofthCYni
JC2Lda6r6nGNQxuAfaFqo6k5KjbgPXwat5MqRqIhvRTYbWBXPWh7Sqt8a442
iMQSNjqmvRgX99OLBYRI0YKt88Mp12AjQNu1i4ITzlqXHd4juY7nEzn56Qdh
euerpOi7nVf6uxF/M9FtnQv6/54oCJkQ9YXpv5Yp2xNiTwvvMzboeukDCOR+
ywkPixXgeu88qToM7lbfQ0qHqwaux8splTUxv+mbBX7onp1aKTdBWjsuvKar
qTizXmMBlhN6MyymD5KKNb850X+81iQkaeGaLeRl6cX64hjyckhzIOUXGQ85
jNhvWC4ES7HmEMxxj0a/RhN0pEt8KztKw7uNwlyigaYtnQJk0mi8EpoDxt5b
hAFh+wRPOgDbduTyg1CS/zPIIivqfEK6ZIoRgK0iyGoA2dlApa7pj1/210e0
bYsLyBExdbEWxZTzyiW7ixn6WlDsXTyEzswfPBkiDwXXbuLw0+UERLbeicfM
jT9WNEONqbcZEtTCHTfwNaqS14YOkhycZghASwZFk82NZXZgqNDG0orNcNKI
qOymjnegYq28Kv2XAvzvz4FkcC2CzTNElTkWx9yWlitKbcmVXCk7Oj/tHCVI
DhHVk0vAnPm36N2LGSvmyJmwF9zqQM9PuRjljN0WY1h0aLDJxplrqHX/3pVL
jPJdY0chhMquRIcM0IUkRd75qO55+DbE0PvTwneEavJdQn9aSLiG+9O4RTyM
y+jRVI8Cid3Cr36LmF4Xfoe8pw2trgk91/MBNrbQ2ZgZN0q+OiSKHE0ENoe6
HkFdfTEZtLFv+tEKEnzFGbMH/qBNwydhd0fOlH6UFkSoJuFd/hAB7xPt4Oo3
vXMjOWPXIAZqcFG9eZ3N8HaCdVF3rGi5n5ppoC8Y/CoqQxg0PlrW2PMKM+VJ
8k8UMRcm2hXpx0FXxkPR8xH8kQDAhRaKFZSVUMFd5LjugZJF1O/scENNBytm
OKItS8Q7ygZQNyUE6+Jn3DlDPvEzVbvwaq0PhMc7ailM/LoU9YDOppqFpFUd
fn4iYTNzSgsLz/PI64Hg9F5q+//mQY6h2jh58TqZNQaAKJSb4HsFR/v7jgFx
cA3KCkkGteLQOBQELfTXsV7o9NQSAcSpxYqVfCFRVVPp7MaxDwwWhMm17pPu
NuaM28PMKFRwr13LZ2MwS2rPC3/6JxsH37I1FoxvzbyDGjdzh0of7dIGrhtg
2ePM4Uo5cA97aYNak11pMMcpFsfH8yNtRu1L5FapKXUQo4Mn8DOK5m8eRzX7
NdQdHBc3/RdIYgnRFUOag+KjL/qf1obB9UUIjNkpPEWrZT+av6qfghf6kxi1
zE9+d0TT61eIG+N/wrX7FwZzYSZe3MIP34ym4mCejNTlhTFTYvM9BYeNOa/O
Ltp7AZBjwDf0e4HVG87Uehzy+liPpCy7JV03jNyq/7kas/N1EQIJgnmnahV6
Jd8kJkNKTrNW5oDRRhY6zVwYPmQcCKs2XLaqhknY4Ma5CohR8stH6ZnfBCpa
/6Dl17GCIGBvwoe9MWBl1hROJyDFD4D6FBS8L/cHZWMLirobftCXjavZRToA
E5nuuwP1PDrBNNOH79AfaUjY6yJkMs/S6/bY3fKXn8lPeTm7V8bI+nYFO/bW
QwfKYCbtlf31TthedXxAVTyQ1DWtVj9BkPZAtWkrFQIHg7zt0R2EeXv9/psF
buHPh8/ekBLBOEODOfr61HXrW7OgA3zy6HfEZaYSXu4P1YWXtH1vsSveBKgz
hVV26MZazUSofRGNBa0Y77TGBoz/IDEq371Ve2xeRn3lmu7ftNxVPYiBrjQO
6iz4Xpdw1uJwvxuELVgo8EQAZzAraL2en7QSxes8ZZk06WYkEdTCOhc9SRA9
+lOQbqM4N7MN89xFrSfmChooSeSI+LOtd28fUuvAHowzz3zChVplxnKvBEMy
+nolQ3iSgv7ESJa4kSTjTWZbW8nzAAIk99VwHs4gAy5YaBEBRVZW0rAyKy7q
NMY/WagllEuGheIgVk6ERTfv3JWqGGSNEBrgDjgC1Le0K6C9BMwz++YjK2++
3W/MqMhfIWgfDBu32s2RSc71ZJVeB4Ku35L1vTEBCa1G6gXg90Dr/wCkn2B/
99z0ppzlBBI584am/OlEmo5pMCHdnj1Gtplye9fupaN6PMvdNTiOeXGQTbM3
f+ZoS2z6HS89vLNxNwmE5vbA+X2doDwyzytvvrH2b/YUVB2L9pd1YIp18KCU
bISg8CdAN7JOrGNuHwAyza5BZxkc4az3ozlXGBQZnYGgVgQioMhocxFyXrgr
H6TGxJ7cnDnAYCPFMcx9fdIWcNVAsP4EQqneFpx0vOknOQ+UxOcrpWYZebUR
3sYcW7zYYI+kiEs3XbiMedkEuuw8SJ377Z/qP9VrohwTSn0UTVQd7BVcOcLG
CUsmZcADrjna7gjmSwCy/q8zYYNgbTU1BLALUpyXfV6WW/EHe5AhHvE2KLmD
LtIO2I/2g9IcLfU6JOOU+w/I0RbT7pAyB35V9LWXvCbwQdk2S6Uyk7F30KsD
2ldXOV5p1Dnk5EIH9ZDJQhCvlR2fE7hcWwbqNb0hzTzVDHTMbpdd9pr71++x
5nW4PvgPFZq4AhdEdLVL1x2caNVa8veljqUr/LE/i1hiIQL87Ixc8bmu7EZK
guwLVv74hMfh5mZelyKa2qAsK447QcT4jd8AiP4+8f6ZyWnsKkQhpD9Wyr0R
Ko7GGo4l+8l3HH3vJAJdYCCybVN4YibjSgJu61reR8nSzQ1uJoub42SjaTfa
lwgwh1wkW2eRUVdABnnPDVaUdiJwk3ZowI0ol/I/xx+aYAB1p5NRCq2LYUQV
96fn2OtewN4XyRm8avPjOkDASH7ixbU5yXYKIqSDXbBlUi+BquB4GB1/jAu2
TIT/kr/8TPv9GZvO2LtJ0FEtBxUtJmTiqE53DmUJ3JZeuGTPtIvfV7cnLttf
qLDnIZ8mFEFadC9VRgY5C3G0LCbGUhFRmKt+R1H5IvKBOmencHI7uwOtXXmG
S9CcgQHWIWAjBzpRVTI8FKAXGLqI9EkacI0CoeloZOupaElzKXxXmkry+YEV
QoByWzpw1RVxKgbdSe+XBwSBgfQVm/ogdq0rCQo8f8cIguKVm4bLw+Wb5DDK
ETAfKkbHfbL8ZohGvFY/caEmZ52d/RngXN55q7s+IiEiouWw8OPZPrAgIEB6
W8+ahZHY9IloCzdWDQbfsQZa4RsTUKsdkwwngakCxmPWxWXwCbCr+mw2o+4F
rP6PNsk8RQn1booH1IqJ7gZtBLe3JwEpNT8FVmMgv3HQBrGJ1+2Nv/T/mSji
MlZFZLD4C4vSHIXRGrUQA5ddt23krFu6jLVsuCl0MgpDCLo1bsxYRlakU4He
cvibsQpGjYYBcZx7HiYlWioyMJsnCha4u7z7QxnDs53/8ZkL7JQegCPRDhee
ZU6e6RwCksWHzjRs6d8XDyHxaV7uK+KmCerpUZJxev+LxNHHROfAQOk/I9Bc
VZnV2AlRXdUl0+CyZ1N9hfcooQHKxRb8rd57A4ovAFy9Pf+nlBNYa3pKI/JR
aWJLrCAIHjLDsL2tXDqBSvlZz2PvJTsPP25fXChka53N8AqjfnW1ttbbPqtf
y0jNcg4KU+6algXkBcisJVVPpjAgoMvpVoCy26fh1ZmBmsA6Q5O+04C/Ddnd
w2s0U5tUDjc6aMT+VS4ESvPpSh+Yvh7sg9LNxGj2YHH5E4Pb8tl7wEee0XPn
HFFKStVkrZf5dJO+uslkJVjuaWEhtePxLJFpLjvUX71ROcDsUMjpo6b5/wlE
YB7WIV0tJqO8g4znFLt39Agxw3BhwlvLGWHQru1E1ZqeuW+kNTWd6nLpSXeR
KQQN2VZtFcPrFEC7I3EHvnwgXbVNINSq1ocUgDdlNoJ0bwiaK3KsVwE+SLxJ
G6uWUB5vlBOqylMjzs0iGgq1a2nLHWkoDPx/ia4gqMVhENS3LTTVg2TxcUDN
yK/DPXA0KalDFokTmnVyk7n8tsfspohE/yte8OE22sYPeh58SjnhcbEGRNkh
6cLdd7CA8NlsK8b3Ajh4epatIbd452zrEglUbWLTrSm3z3v3hiFkfnFCmXQw
yAnEEfcOD6edo0Pi+MjQn1Xnlv9/xaMkFcng92X9NgaFyom0TPtCLrccY/ZH
r1k1jS3KowUjwWsVlaOt1KcZUITCke8jjlPbJqohTaWLDDgaiYgotIoAkcJD
di7xx1MswaktgOkoTw6SfC1JYz9uW+xuFS2YiioqwTUFSvscfzrKXTm6i7gx
O19HWBD8lYHqWPd7Ylhr6Y/B413L4NwBi85iO30Kz+gbqxWjxgKD7+OBAogm
1mfw5owBTxdXV5WRA9mlc/Wg75WGmqBOFZb+rov0vopdb715IMDpa5zf1Kio
DaRbo2uHKSWlIW0anGoKbAujfvyt9mUilWkGrm8Iih21sC3Q6yQzrxaKj7UW
a9lkRwfc/BzcsoVV1W/Qyg7kgeA7vtgCusTxVzXrxoJ22MkXUgL0Xfb46Gsg
qJ4A9dyw/jrdxHFyO6EqRbugswroyPePJKAEK5ulKTklna0adBFstwN1t+XS
hS+2MJPp37XrTh8lrQA3T5vmpbvPXbmTMx6+Ta3vqtNqmdvNnV39WVIubHV2
SB2jQJvnCgogX0gcrTvqcIvLWhYOPlJwgPQNoBvY/Z/VWN+8npxOLMiRzy0y
wHpTee8HqmdrZD6/Kasmw+c5pqyYeYDsmnXmfUeofld47i/V1wijaByXGhNM
R6s9Ei4g4SA7sW089lmSmRFmKveBFwRuDW9BvM9/FsDRzbrH6Oxp+sOx5kMY
GmzHqpmFVv8t3CQfSmhnf+pswr8nIoZ7hsvK0UfEA0oQiMatcm4f+1Dr2wUX
2HFunA0QCg+S4xFwk4IKikg+2GDdeOBeoEia1Qc0w0SEgFK263CNr5SlxvxT
ze7q5yceE22mNE7JviZW6s91wV1Y4vjM4+WyHCbJhL6pQssyKnNhcvmUU2Rn
KQfb3ombhCquKVwEUCu3NrTaevR4COGatsvJlk/cB9fPI/OPB/edFUkYRcQQ
bRctI+tOOkwFEaZXtQ4W1KeF6Fp871XI++dV6FQU/eZmMjCHacxQ8BcWrV9B
gc5GX/B5jMLoJ31ciManRng2HFKGT6UUZUUXGe0bvsVzMnJ0cuiREhitlpWt
TyimxZeQdscIXLxYgFwHvm7nyMFwe9luUbBcLuhBIXfi1Ed2wLqW14XrkqMM
yNf9l33pyT1nDROng41kkOP4RivOttvt1rXRAE9YqsvSdXMYcxDTgnocC6F1
ikp4BrKCYewvu4y4ZPM3s1y5Bbc9AecSRGUaP3Q+DYLMRxk9rRaHT1Qu8L2j
hRN8tlTWn5Qf80zCX2OoAxmHG0GjE7jEUH7WUymyKVNUNtiz8nQgsZaDaQad
eDPmEffGjBjyqDdfW04qodi8ByQUrlXg4gLzt5tmnyA07YTlqo+xp1OVlXL6
hMyo0ehVl0mmRZ1g5RVV/XZjoD7w5CA8hx5ugMiF9PJHf0HiY9Sma3tG1bdY
6caeIZFMH2Yg2If436AjKfgYEIrnHzGItBLHYlt0K3eyZSn7Agx2BR/UuSCa
5QdU6z4som5GT/IdYqjxCIkrMG1v53Zv3rsRFx4VmkzagRQyr/blYjdHacDS
Y8wz7HdqSxHBvPj9jXx0AQZI7NQ6Sv8KLzArqkjLWFD6rdZ4U7fvGuzeo3SR
JNxGh62V4WOWglL1hSxAj8euUBiJXBbUJ3mk73Dyauxy31uftMnh7ZqkkyKU
+k+PziLW/icSgOol0KlnKC7fw0ijnx1A0j7LPWodrQLk9cEnBWJvjwTE+XZe
4PERm66SfjOv9iBECjizoFHKdjfdVGPHAnIxmWJuWElxI+Xzs22qZJlxgZmN
ZhvMhQPBvC6q/hLFlWBkJH76RTtbZHOv3XqBPf+UMz0/b7zlQejcrjZSZoj7
Piiaw4oBBSPGtb/kl/I08HW3WenSbWf2dpkx907uMsYEuf6Jrl9XdZv74JFQ
MNgKBFyeUEtvLKRXxSouKYDCSRnLWBVQPfVTwcZYtdmZGoXH4eCF84j+XYlg
rIZeNBa26cJ3yH0MI+eHat6Lv3upvNpauEJG3D9lnrRl5UlnW/YScPHb8ggC
qRSjrPuWwfhKc8egqx5tPZ1YE7vUGoOv8l2lResIXF7WrSZrch2l7VknfoTV
f+w19szNmCiaLeiqyGguP+mjW8V9D+t0zM5kRFh/uYIC/SvT7IgCmbqNTAr6
PMVF+/S3MO1cs7asTg+xE5iXAifHP/1jsqs1adqMn6ZWnZvjLwMFAQP7bOW0
O0w1lXufE2ulKvyY8DJpsri3yhxBAVLNhHOnErINhOaAAA6G2tSe7kGgzFaM
YlQvzHo4q9C6U39yqqZOuDj9XnqeUztZrb84V4YOCc+6NY6/mXGwUBHM/Fxm
raq22R10K9Iqs3xygrIDIqbPHFXPv+1beaZ2l4J75YcB80zBbRCOV2plDneI
yBG9IHb2CLFTXdnoGrZvg7QJDIlj3DflYzVi0xGVdqcRNaPdb5/zpvbGtNOW
2Csfs88qyeIZj2qTiNiGJB2ds+dNmIf+VVEEKr5Jep/9vhtKKW3D+cc2a/Zw
QVkgAw51MMCdxOhTSm3qeuZIqmthXVF7FWCL7y5gwMcHJiQh833J26/eUlBP
jkSE1gZrVnLMg5n/2Hynuyb0UKr/rSBZVxT33uaNjJB4lNDv0J6IXoQ9E2Y7
VL3FOmwxtIhk0sbt1vq03bwz1PDi8PierWLO5GoT4sly1D0rtTZCwAmT7oKr
Xef9VNScmqKFMOKP5BKV+4k2LHEDUC5POGYygfYuh7P9z50WPGlD2Pn5YzCk
mjHTHe4ROYJe7DBdyebyQRuSUb/Eg/2/MMU5PWLhvFP/30lnkstOO2YC6zpS
UFzHgBl+yKiysB2ERucIGGnoIo6Lp5giSdqJd768gnC9G8qeIXlzzGqNs2V/
R+NhzcAK8d7x750d6ciyuMmI5LZA4RsRla+QTq1QCdpYY+zLwAoJJPzxbAba
sQdsyKe+68rLgCREbFRM6buwdqrR62xiHfbf7CxBotLHyajzJ+sMEfMaf2rL
BqxRuFEI60uOUa0SSKGvqyEtFxD5OTOKC2kcyxYJhyhseuQrKDkPiWULtQYY
iPTL/HC0KgVDujE+yyK7p5SP80WBTIfl/AqOs/bnQ6K1hgCdTBbLmJ+o+oGb
dSgm3qJEf3hH7ZtaP3oOFTUgkordmZvpi2psBDDxUBPwURS7Sa3KZV3fnN5Q
WegNZtTii5ywyBJHrQp4Wm2aK2BhiPYz+l2BFmGzEXd41DRPPXACI0TrWqea
1eAl5AJPVdldueCsRiiBrF0I3VEoNbk58vbW+ZR5IxikilwfZc3QgHJFmC+Y
WRHoq0jNS6qAQzGTXIDoj4jJ1eFRovF7K+24rvRT2yvZUKNSA5jiu3177B2N
Ux3k0BT8m4MakBwSO0TAvGtrNdMd1YFnJEy9v404qJdRy/cSyVcb6HMMrzVL
cZLjsEPpxQRTP++PlBIkzjWF+ZHUqFXhswLfML2sxQQdIAQZXfxC91CjM1ep
ka1Xj+BsTVs/pn6/tM/AJrpi1XDVJMMk1LN3Rf1JX3iJom6WYMa6qb7ounDI
oXfmOAiSvAQuvVCGDMupt+BIj1sud3odKm61xJe4pKC2WibKqqxfM87j5m6L
D3we2/gul8CEHw9utv2X9Bv2iHKyCvIPJ8ag8K2Kft+wJ6HureY2tR3rFa0j
KG7EKvPaOIClNM7OETsXIFAjObbQ6jA7sz6TF/jpcZUB7Q73Sh8iSSu8U7Wk
690oYO/+oRt+9GhJzssTKAN8jc0Lzb9epPWrvFXOhk5Bp/l7lXfONwHqnna1
aPZ5IHwJjZDSRt9z1wLRP9oLAF/qe/ub3vu7fn2X2gvru0TmD93d3SzCS6Ai
H7Do6a5e8a0/hjqPHc1v+szS+sfDdMFk1gJHfOMvofPRabfW64n0ETwr/rUY
UXnAGDysQIzTACgq8g8DCJsOdc4pIkmqNw1+t3LASBrc+o2MAHTFIMeFCPMp
JigShM4SFoBLazTwfrLk9abiyWkv8RbbSJlKjkz5dMN9+2MU+fSTokieIC9D
QkFTVYeCQF9RMQWQpYCyg3YR8Vs79O6TM1DI8Q9P2u88WITJ0RTEkAbS9mwx
/2GbBI1lIfYHKrMkHFDmqKQDxI0FiP6NSGzQP9LXadFk5KxCBbOx84klS0dv
CASclPqvYKJ+zfqQ8dyGCclAz2YDgv5nEtwupdClwd8a8C8iKUxzv8+Z9+3K
VhPoEZ5OuNVLYlbgi+4l4zEPMsYnyCDcZqvDmmwRMPyFss0zmGjwIVG0KTyN
hLjn8JTJLTukRaFoHH/cdWD2FMgcA7OiJFEELXxU8ZChh+yH9ThiI9tToeVI
AFPExUH0DWXOFraYWrK50GLxDZHkQpDKavt83o1EdddGyOOUt6I4uniTuIuA
iYamIQSEQnvGKZmwM0HO4YATHZEMwIEj2pjKCM/5PPIA/copHaikmEK9v2eF
KP3Z2rDKasloXD24dcwNRn1Gv2bjU8/fwzN43OyQOF84QNjgubuLTx8scGpZ
dtPGCB5nw+hbWnMSvt2ILWuEWWNncF3P8gjJjC1VhzYLL5embptcdiCGRt3R
94UrxgMRuWUakDY/pHbl+9cyjlfYB4ycIXPAcNb4bcIEiggr3kArONhEMLyc
8zbV7DJTdXt7itD6oNttMhTTMfKl7/L63RHAaROslS2MRTjIOXXB+mGMC4QC
ZYSemyXLDlFMm9JcYz+cD1YngqcftpTEuhJpfxiiNy6PpeD1YFbgjwRD74ri
QR0P4Z5oEwilFnQtqR8j3HYz+Ml3neCqejzQF1GOFF7tLKAotiWJSPA1Di3l
PIMMGdTJQ0d68C0kgoymvVr0qf9K9AEToP6giPRHBCTXywGPXT7ByGcfDa36
Qys3czip0zR8hJ2ut3bLzPPhMd9IJHiK2fXzHZvZZSYBMUliLg4seXvr4zeM
zjtrTijIu728X9fjjfRkE3wCSYa9OCuYJVlQ/iTAnbK15EtSHaTUVD9BaRAU
f4EdQJXCMJf9liIrd87mJj63M9JfHugVSuTmSjm6qOC9W6J/45c41+ujO0EI
ElSnR0uLYhOqYp2LJY0hyVGP7MoJJO8hIVTiDLpAyq15K5KTfr6vyjLMIwQM
hhqc/aQK92xVnLNNUyCVWNsZrC+I/93s3jPvz8wA1LCJFKsFnMnQOXawEfSn
gKslHBzgbTr/bj/XQaMd2cHT9ClKVmMYexuecSEQyyyumpkvlINaAr4BouDC
7CqWRBP16lVyNc+P08W1gnW8lmWFJ9DZ6o2+F+BT8bXp3gdvGzWrl9ftnnbi
mmSmYZ9qoC6tLs8dCxYfNVEmYHHp0hdm880Lu9hMpD3W6+zLUuiDvyDVviER
wS44kE/kT1IVWBUAOWiEB8uObj0gk+AG5iw188DVbhqBPeBwHolDF2xchOmx
vTrvhRvv52iKck5DjyobumINZ8aEkBeZ/UtH2oC+Wb+8fURKex2zbEKQjRFn
y8M9mmv4laYOWTi5DKQ5klJpX4w6LaFYhTjvNFqnhF1VFXkTJGG+ihIiI3cV
RqAWs30Dko+naD6rl7HOeFMZhnAuSyhqFC0sdNpF3ipr+oqRxPv0pQ48Q5pd
MADW7Ooi9w0d/SFcDUfQnhb/3Ht3FvOMwGc9eL55oz6owOKoSt5TDiqHW5Lb
4fVnymVy+KctRFXMHJrFoZXobwyhccg3iXU1rS+0cr6LugzDnhr20FDOoAfZ
d+ncSKrOBe81aQx0SaUKHikT2nAYccl7ACPjs2+dGO50JAuLM5qnECAgS74W
l5oxq2j3qhq1ngJ4tUK0kJsu3HXXNkDKCVkI8NgC4WV/Ge1S9gOd5KebxM3e
JpvjjSS4MRMX3O5B662PUGK9qQcqVGKI5BEH6Y3spjWfsVgaTzq077hF/X4d
a0IKyOfp4wCWrg/LXaGLS45PWkiFv2+1/I5cWQE25JoBwvjUHyAK6vnJC+Jk
iu0JltScIHL3vZnB5NVBvGMmDFST2TpNvM/lmbVUOjqFSMJTMX0q55lBMYKz
SdmjsPjBQ1Evm5JbQvxsMdm2cxoUZ6TAUODvnv4dIPYi0mSkIXJcR5uXwuRZ
/8as0xu50ZyUYzwFq7+Ov2F1hOloskOXPCR2362wJ+6IQrw7zd9Y1VXxxgFO
fnTzGdpzcJahz1gCzwvBjLgwxObWxrmJSmtsyiYpji65Yar5J5SNltfP1d3p
Zykwv+QJ3otaDxRCoSSufwIWyxfdYf8TERWPoY5iU7BN8BCXbRt+kq+KLKDu
iqSQY5PnkiSbouEfjhPv+IWgWwsLfFP0AnMxz1ebFLhUjmliy/6rHdyGdqX+
zS81myhjKTfuvA2HE8RonWxDV6Sqis8jHQEL/RO93GStVH7FPPKCUOr65JSm
B1pqDpb1bwrmezq/NduMu/hZ4/sI7QN8oorJ/EwYpSEUonb2zVWiQPFL6zDw
sBAGgyTJBxhQkmqG3oXY11hYDuKCEW6WZacyE80+ko9yLtJdF7ga74CcaCAm
Jbv/a9Erp+hVIeXDsL9TEYeYFllPXqH5H/xMPh5+l3F0zi2xypfOONIfbddn
rW3CUUfRXeatcoHR7KlazYaze3OCN6j2OnuwK2VSnVJhx4nwABWSeLEG+ukz
aGRRnv9DkhbKhaHN2ffJtZtpp+kzMqAr66Qtx270u5YQEP+oO6Z8JcCoboid
GzIDB3uChPvLsBYsyOi5t0Lg8V8KebgFckjY4fA/FePTsBwXTT4mJG19qm0u
Va0KGrI50sDT30IHE+vL0VPKKkGfn0r/otvWqllv4KVJyTkFkbdFYksJlXCW
m5H+tBNK/EuIWKUkisWwr9vcpy/26BEhevNYkXNkO/w/S89hYpJmljD/ok0v
2IXz+UCXf/F4ZD/XJsV5/hOC533ZXFtvSHMsWdvNm3lAdO10lS2YoX17E4nT
J3vcB4HAMLOSiaXWGlNCLqNu5XirniWxqUyRyde+W9Rn+dd8umZXmeRb1N4/
tizRF2+ae7fwZttMF/ZPrPndHoUD/Z0wnxAo5Az5TM9mD2NkrgVKPZiDFf7I
IDZomUEbzhSAgN5CCCrdrZwImgp3HGyEy0GCIwh0zJDZn/s2zNZdCoDoRZP4
Xdiui2AlbVXPBx8Tbw/z80CFrCG4+oI7kU24Lft4+2dvZ4VkTHyjn4VpiK0W
AyaFfgbZrGBKclvkyDLvsJNJlYwTL1FMG3s6y0fQc5ZPufH9Zhz/gMrp/wyz
mL0b2gWVh3+Xh0ShWB8wPbeysRh6lCtR7fssB4De221nwmAd27UcDskpdNE8
CgxHEqLII6B0To06uwtx+CFCQrUSCeYmAd189nf1BN9rcxOGDA2lVgJfvpFd
0coEFcU19zmIFzsddEZNT/AuvDYq9Mxr9JTTtV+N8f7vuw+rf3X63rKSPrZk
lQuQ2d/AVnB6/GeMfTxnYvEX7ii6q37nXfWPM4qevkirlWrcMUT2yxtMxE0t
0Ty5r/0wDymb8qJnEZr1pdk2sLnLTf3kxw8qKp0yl/Zunpqn4bcBxysX1Nsl
PlnCRoo2xTJIPeDJMeNzDevNyk/cvJnj/rwiijpFNeaBXmh9cQ7tFA6ZVtyP
pFmZiTlANEye8t/WvbEf/mLoDDlBT5UDaZsF7DGNFwv24JOdqoUV0ZIkqFVy
KkgwgLvHdi3XUqrIAWNiieCyYpgcMnOODRx47LS5ajZtiVYiiIcTS8w8IuZ2
D45d1P2roi4okKR+y8g7xBlAw9dpIpQayPTwlkhrRP3d+P5SeHuW1xkKdud7
Jds5rec0vD1RwzKYHyQ1EO4c0A5vh9Ax/PY/aIZeUJmB3OvYtwXOLcePGbLm
UsjL04FbfipLoXb6bFHdOAMYB00uGRJssI+sRKvt8FcbNYiD67fOYmdr1KfG
NOZXceznNZFXJkRVMRhoIW7wf8/J4vXu1d/FguFPej4bkXGPQS6YiEtQhDvd
kqzQE5JR+uklZ2k3Rx9VhzfYDDQFGRVXPVXE4xprghlBpEFYBJOZn3tHs2CX
id4NxyxWOaNcJhox2HLc7LTV+Ja7CvlKavUG1HxN2hXwKEN3FaoBKWSVzZWs
SGNyCMFAXtyecrYkamuYSiTirIDzOiOFjkgjMYCrwkP544D78PeY5R45nofR
7hgA4b02bDdSx8JLTGwYj40TtXE+1vRJi7yR/z3E17MusuWEgs1DMNUhnXqO
ykvcu+5Jq4q1EoMEsRLfS1DZpbfR6bTMZIq+d70pBKe670ntSobKXvV6/Y/d
yaAmKAykLQafpuNDFWGt38rKWP1NxeArnCH98KHfeUoAB5JHh9yklkctS/iB
j2Ua33s9RvDjp63O9Amu1utWH9k5LEZ0CjEC6vHRRm2KE1VfSyWlgZyoJfSp
z26g74JaCdKl04UW4+P9wqdnbFeCwdCROqH3uQdK2lAoEi8ZjcbYc2fTEJHU
dk4pNMUp/HFihIoko8zxZaXWFmEBloCJ5E9yW7wlI8jYw+ZVNttzyxOKaFEE
PmZ2wcKRLI6L/UyeXNl6u664KOx47o+cVxMIzSgWBgymnV+FhJaeNlQvl705
f7+uYaGZkECBHosMZmYDo3estpe9jv/nwbGc+3O5io9LtbSE/nFHWZ8vYjzJ
PUdfW3cpkYPabV43fE3uiBu6A/apDq8v7WXfYKHNd+JYF4fKARG30vfdfz9P
zS/VavDQRwLCgcpTmsnks4X3herWnl2misOssWN9Fe2oN6IkoUGbtudJTkA4
5cM+UlbxEiKO5UUKaTomPsHxrMH2v4qU8kWAdYKoqrOJh8Asz0yIBSLzNgQp
WsLHfTI+2XgDmXwrf7Pz83X96C5U59wYLSz0tjA3mPmgXIkyDzpfzweOlnlO
IWVaBDu0FjSJJ1SYLeqELRq0o6NYcPPkLccRBg/1CL37dI9o4Z9qNpUGvKOS
ZQW5A+o6eh45PJ3kuMPExJmp0EXPc0gQDSIYsIe2EyS7B5aFj7mgGvSw/BRK
E1/qT2paVA7QOINLUeAJGSyHrPg3519PVsXe0bWeF2j7m/UYCDigiFyPyCSv
xhRt+kGTSdzRU76LXYWvM0AnBVTqpOiNtx/6/ksSuZkrHb4knVesm7ca3pcP
QIqqQ4pVTkhOtpVw2hVSQBZSWm20k5xbs+brgM8YSpg7aOS8YXuPWjJkUHRU
RFpHUj7ye5xh6jeIb5S9Ugzkr+PRwDOuk7uFJh6wQ//tFnIbWXCGxmc+KzrT
5jYAM/45eCoxcE87Z5e2/qpjCECsfOGm1EBkCrtAyKu2WqkSGeZFZUFdlILH
+R6lBzRNzZQimRkDiC/31YifywHU0YrA/KHAxtwrWjCN/DNGXpc2yOxzTe9x
GVsBQGHC8JNdb6hIgQByI61EQ04NkCNJKmPRO1Ug6h1z9Th35bL20KTdhefY
x9YYjvSaO+fq5xeD1Qo7PPE172cuW5lMfAk/djFrXYAhT1hGXmbYSSkXj2oH
L2c5ahyN5nKEyziHX+C4m+KBI7H78nRKF6ZM3t1o3uigQZ56Yfv10jX6Tc9O
G1AqGUPMd7qFZvcnPxV0fODXSDQ1MPs8YoLaZvnHFLSFUrZ+QGwBIT66nvoD
4RHv5HNn7NVBSIUPB9Q4kRwgB2NKOKvJB2z46HEfM0H+jXZQHsR5BZNfjuyI
BBIu7cGaKzIzCG2pbtiJvV13m5nWUE+XilRcQZ9M8HrCY9AKEb4KixWP7nck
GwTkzbAKya2tJTD2O/nYsYJnbCrVmbpKq7DJfr05Mpqu07/L5muI2MhFE1xX
9lD3u/9UyMzZMoCKF9esm3TuAq8tsuPb9SJJvqKBCCvsK+cA2v9OhkrrCq4O
nmO2XZSxpYnKeRZ1xJTG5yeeSmAXJdxIjeiVdwePzASWEW+GkCl9nJ71GGay
E98EXgvfZDd/QO5X6Uk2cDoQJfR2w+m7EGB2ZtUCQNVMNlg9fMvHiRfooS0H
/55R+r4fH1s9VohR2dgr/OpWEY4L1CL4MKwd6/MYPd8Bc2B08biO5tmKcTXP
WwFchJjCPgxFFAKt3i5kUXHaQEfIhTpxfwzwVkUkUD9QkzUxnDM6+jPEtyAE
BWnlG7jjIQlnh4YENtPxiT13tq/Oxk1OdpH5LKZMrexFGwGzNb0kJ4prbne/
4w+VjAne7156fiTm8NMJ1MRfd7qog2oNIxsyt0Jo6aY0efIYw9BXyWhkA1kz
ysUwdG4WcHsIFdO6eSuGyYV/2+da8bBiOspz2MrLbk4CKW4+0fy0lkOaq/IR
OVhD2f17Y+KniPQSTHh55k64NX/6WaF4/hXYNDzqi0a1db7ymr7pvsG2+xqL
b/nmiwjwcbOCoQYyOQE7Sszfn436AM/I+HMLkx5oqiEibDNoIFyAU3xBsg14
64ixONkK1b+2dqeRVVa4ji2XdO75PQa4GC86TMy9gBYtuxj3l4T7P4OyU6T8
OnMtPS/ow55/8ihckZRoqR5WoYSIDMsNWYXWDdRZOhVqoT3s19vmzc/5vzht
U2uQIXtUgq4z85k9lQBKZUcUGqcpHmEmSlTV5dTLsPahOxnYFbArW6pMhN9x
+6e5DISniLQM0udnOFGGzLxKPsWHOSZRXdzvoNlylQTaV5Nx6lhQ2rQ90F6z
WkIJKpdPrj7UmgkhE5Anzu1V+GmtMSnnttOmwLsp3nH58rQ1EB02UBYZy/T8
qSoGQeisqdJKRP6+zjoQVJgesW2A1zSPj6Ruovpe6N958WAP0FPJXLiIB3gZ
YSxkneKMKeKmiMFkHnXuo5L1NA34v6Jm+75dfkMu0Jxp0FNA74OO0WOs54Le
9/G+cyWiamzWDl5SpcxxV/k2jys48nRZB0KubNCPwBZdGOHQsvNv3rrxsbPO
Fp3nFzyCV8YsYZR2nlz4hOiEziQ4rFTVKlOykOU+4Ip/fGEMa1gKkaDCu3Ki
DQBufqgfQyYRDa9aGLFqMZjIGSwWSl1v2o9MqmLOOOlrJWnXWzedk214ux7Z
hBr2yGR0bH45jj6q87svatE6e/KvY/0e3M9O/2bg8sQaBL1UFHwSPcsZ4oQX
QeaVVkEKx2nlxlRLYC7S1s0rVD/n9kU9jEGTllo9wzS064IFQdk3q9ESiXCT
SR/hAvmLiRJ9W6AaZ9fvY1jRBCUfTxEg2Wp6Ny5noD0VVcvDPlJ4PbkvS8OC
v4IZ/+XvBbQ2tbRe8FJuSEBEqblUfrJF5llGrx24F+4ZBNXJNdJTVGXj4CDs
co/wP21O6K48l/J+dsm2ZPJVh+JMSo2fdJ4tvn63I+VNbO8bhxbCuP6Kps+h
62WKEi7EieBH0gmkWgh21P71KJ5MrKifE9Kt64x244GIGGKBYBarFjeCXV2c
fKKf4UEq2zSwlft8V5w85LSa/8i+iqemhOcDQM96cANTKd3WSAoiqWvetGf1
Y3QOlr8Db+M7rSm8SIGu/QinWnvXsOfUPl98IvfdxQNNSzUYOt7AddoSWjS8
oNOmLua/1F5PQGGygC1MB71aDm+8vE3Q3ccH4joUrlWvN1sdHT3XUlsOIYMG
YgVJB+mKQF2BkOstCb6Tkh8aqocQ6p093Jrc5KJuvKqQNu7gOJnJYwAwp8Tf
1Hit1iZEJ8qp9w0BmSGUs5kKtLOaUwFs5rseLToxJ3kC4BqALs487fGabh4Z
F9/iXlmtgCi87r7dJTpuXeS7VN1uPbg5jfo/UObO7A2rOIuQGNU4zyE7OEIQ
FAv5LGLHWNFQcMLybReEumgIwysaIFIRZhhFNU2N0nKUEhSXiPrOUxnIF9Rx
kRkCvDncB3TNuCRAwc8MXwPhKSaNEcIxoi9mUrtBoGOI+WScG7u5JWv18QX2
bqzEstVHprSNJ214dpWppH7PnH+aG1wmey/TndQzr0pgA5xc6FgoMJBb9RDQ
wg/WwC04TGAm3ujAogPcjm0YSaGpYLs0J5E143yfcG+ZDit8amj/V59uunX3
pi+PhLObTp8xbBL0PL4yag+vojwiksmZje1RmS6iMeP1D0P7miC555pnbsx/
56WUM8znzUHNxXT8qzDG4THdCWJ7FbyWMvklxvEdKyemBiU2AHR61sWrFA+h
nfrKWTTKMjEPimRYe061ViPFZS8Sh4soU7wtSCS/d6yvM00dfZWxaK3aNd97
/CUnbORfiaEthvc0F0R9qSZl0uu2UCcXM0XqmdPcjptl+O80ccqsX49AdCNx
FEogvs/Zn1NzKB+yA6snStFWpE3Mhr6CHKmqLhxACPOGn7Xxz1E8EBhkW08l
fg6gMNHGm4Cu63YgClE/2D5wa40QCFLlvybDLzsYwhuAHVJORUCXAMoealx+
pyztqfUJRzqXpyldZDZHPUR2W0+oDRCo6YbtO2yevpWXj/UvdW0fK5E3bDR5
w2UA1rDiJBBfFdjP4nj1V0/65ztvPDkCtxX2VJyTlAwkq6Ppid9wibIfCB7h
vwMcnvFmwU3hrnGuC7CrN8nufcX/oIKlpYUk092n+vRd1uNykh9l98TuQ8vJ
z+tJ5+nm/u4NjITmyRcj/eOOuj5HFMg5xnfC0gZqh5VxI5m2+HOM8Pz6duJM
PxpmNYa2Alf9mX5f5o38GJ32oWcKBToBC8njf+y1RPclhjgXTSWlJ8p6fB9h
Gf07s2//ogz7RaLSHX8X0OP+JhzzZZV2S4RnfpWrywe5teQl2ORJvmhWKqT3
q7TYulydOjRpygCI8ryey2XwKOkaHPWbu6TGy0ETX8T7T78zaXYUmpl7RNkm
eh52Qvcf+quVCd3H1IKuywCEjpllePSaTqM1E7xEqiwSb2/mxaHIzfD6qQe8
x3LVaJIIKeKKls7fxlASVosYMtc7A0XAH/kfepyUR8ewd00w9ducrP1M2ERb
zGWHKAkbcqxD422vZJ/uayNDrqiag2HuCMoZeMVKpjR6s9pU+XXn/H0gYQle
YsLvCUVC3DvHjruiNW9PX8P8YHHCID7ZsgFddBVacePJypfZBMED5ovevpJ4
0CRwpa/z9p3I1+msV8VD8skhJBq1sW2fdfxHsVy2CpoTC6Zb/XUtuSoy8WgM
PvwS416GIZ5hkkKpAQT5qKQnpgYarpWz93IlMMUHcfiqSkLXrB+lmd922s9W
CpPDNOa9OshcK31iSU2/tgOGKtUZL1Dgc6wsq7Jb+2lM6z3fGB0cGjJAQ81I
Du9LxKyWZw8nR+7Eiv39K+sVHPa2v7gikFDf4SV4rx1DYJEDbMIUBc+WCYoo
w3cYzQEWT6HOEbEDPk3vdj2NCkXJV0kbRbOWEtqpT8nYO+RaK/G4EixcNURY
7mj40AObpqCkzWjaj2EavIoJ1p4i29YggQUeOFvebVc2WqQye0krFOzqMch+
eB70sW+vnLr1v7lAjaMpm3hfFVsRhSVE8o3EWw0cuFxxqx6MjspKzuWf3VvP
ismaZvlYYe/NAqK5bzw8GWCSAS3eCtuAvQ3rljB+UbRRQVTb6GIjXeBXdWsY
DbQKQqV/RJLulpUiRPWrurwMvfSqwXpeOjd2/wWwpI9RL0yM2TOtBzgxhsHw
SZqYqzGfME9BwP15U7fCYLd+BbLjvUfMwj9yaeBNA7+THTxA+kDyp4NQDc4w
XpHdqOEdGkw6kO8wxZfVCSddmLmZtyYezyDmwpLd6129nc2AspsxT6i0Nxgs
42FKLjVde54ov24pSZjjBbXYwGobHDnKVomwgLFjCH8FL2OglmuVpAYboGEC
gTUH2NOSAToF2gBDQZEWTs+tiBBkNu6O2epwczVrjLL1HcF1GVouzR7nmeNE
Oj+CcfPKbJXXNVl2UkS3qBoHoKvlYFgKOfZ4kzMzzB35Xvu3FUpyBFTlGm4k
3iVZE1+/VFTlGsIfmDIxiwZ1nQcEVMepCQA9sw/y/Jcr8OSPKYWip+RADqGm
AXtrjvxzqWBCrJB5wQzCE0qqTsvmpYQWOg6sFv2No4hHq8wxcdI0b8bZGAcj
JJPorLOEWWeKEP8cdtD3i/aGwJFdIOA3nL5f/UAczm+Lo+BbLKedUXUrFIM3
oP25W7dzWSMaKykcOpP5Bh6bIea8Ms5SuBppQdy4wlDcLjRbcDhFSGehPaGh
JX88fg0yBJK3cqsehwcZHD1OhwEJwAksv/EKPMzpTvXfL/S+49rsCtiNLzil
c0Q1/G/PUWOGucudoX2XxNMm97BSFpNMwuiv5adjQ2KdLpH75T0wxP3zzXMJ
HBkvRxflSUua6pom48Wtxt2xrQmG6Ph9TckoTKo0GgykMk767JW5vrZCilYF
XyH1HoUBmrQ0oLgqdFtICP4eSoyQIZnaehNKayBxZucFEifdj+2pbjCWn7Y3
S45OdDBfHdz78K0iUtiBaLyGsY0BdGjie5B0UhzYJDaPADY7NVcb5rOhXMrf
fJJP6y1UI34axOlrqOyPfwSgD1aVfuN5DCM56/49Q5400kL+gHxKsf5XifaN
62LhPqFmfd4AvQ6oxh7VQoBf1cT/h+rIa8oIm5G9yjnVPt5OQnReg2+i2ltK
96QizG2SoEJrcG2Uh9nm7KA2Kzd7Eh0lIZD0zYGZnvZhfx92Pqwgv1/auM5g
3StBa0DsCRtr5y1w8t5s3VL0XZhclNxukAkzPuxluwwEScKJQ6iRwrY5pfQx
hQsLbbp3PbbsS8tu4pnrWjLX4hqd1KPn484gUbmzMaUfGvJqCb1vfZnvNMiv
hJIUxJzHPueJrYvUh+fAjsF3COVMreuQgGYwaHfWsHGAYGX+mgMUMJNkFyjV
JDJ+lPh5nou/+h9SiB0gLSUUukvZajUlVsL6OEMX36TYcHaQ7P+iNZ6hBL5n
eXlYkRP6tOt/nbBkQnJ3tcJyRlrjTnU+ufqhW6Hlw8xjgoDSMo3ceDnqJZKD
RUxeVgF4omS5wROZ3t8YhfeoZj7cQkPEOvXnu4YJ2IVzDwrAFBxQgbStWMXq
X/6h6kWT7poN3WZnNaCDDzwtQzAWJs9jWMKY6LzCExTtHXYZ9Ze56BN+bibD
EYGQ905cgwwJT9ey8M7U47LrzXRmxazNQHvwabuFAVU2bb5MAEIDR9KOv6AP
xGhi6yLUYV1nk4FKMJMcEK6I2X4sGpOB4dT0OQIvoqwmthC8f6n/2UlhccQS
nV8j7MUMRoczPTVUtjZ/OGcuBMlrDMGuqjW8bvGeJqI9qrdmtuUMVuImXRK5
xRdBGmfhYFviljCApgH4F1P1xeU5aozJuodA9mMwnNKGu9CP99TOLGs2GXcH
TL0u0h/D49WiIvOdmGM7OCtWnWJuLJtlGrMPxL26YTvc0mUB0U+M0Gg+wE5y
/bSGqCDLTUZie/bgTz/Incx7nXJmxOzLoRl5wix3O4+pxyK/Nm/aAsItntxc
fbzfH8KrtO/Jb4Bx2t5qVNyTzTp+bJYK4+0CaiuhFq3efm/PeGebNfyIQUbS
hDp+pOjLu4qYuOBgOwjY4qk9/yApabXbQz/HEri2qx2speaTDEwfg901jeT2
Gnzz+QDSyzLqQnnDMn+85StPeBDQQJmBjiKMYo+oDV6t4Ea1jbG6i4dUxgv0
VHTJdUlpwWZvk82eG1dJ9QMp9jcOjVD1JK63DlO+5o48RaqwMRciUajyo5cp
KJ7hgNLLYL/mJu99AyzT+DHVpZej1gOCWzAc03+5GVHDtDl2yK/99DQRnmbz
2JTRYPUD43Vasl8dK6x1XRNsGVVaq/7cjHTN/Gg1er52GumQWQQ5rF9gU1dH
QATZ3xVN8pctcGAaZsnHlwzgMJMoG2NB5mBoAr9s8M9kVmigK0VSs68TxUsh
QBMZPkj+818lpbJpL3ktKAei50Z+wpFUhly1MVeQCWjDCkmLM59A6IaYZT8m
X0Iaf6uldCICwX5DHmYYAZ3x+ITmm2hlftfHJ4KCHdwIIkIp0ESsoXH7u8DC
AbKPBnxWLW9N3PlVqGpId07zS7HWQjGi4vF4EYtKRptnDwrvBAy27PHOzHSy
fiwQhbaTpvSYvvWPUXAgLRpuRYQDLWmvXT0cBqvfFgpTuARBW+j5IeatQEcJ
lZkBLw4Ot4oIosorMMPq6/lIDD3rguhkR4Oh77y6338sUX/ikQKdD7EPV9of
/aCL0OUVXFWossOW9MfOtn5TetR4wgTZ28tL3O/WXWGhvkJu1EmiYUGFZzKT
YYxO3GeakmKu4CjIkr/ZMYl37tSR2zAm2vk1A8ymOsgHP/Yd5gnfx403N4W/
AwJt1MXZmi+uDqudE2AasPrwdhzC5w5OdDmnrH987ZsPleYt+obIToxrGA9A
d2Cf2qb6zhVbsh8dfdR/roIEso6bHcw7dRAH/R+NsDCUzds1QDC6/B98DiKr
3A1Twb1Ovn/GzxAG2lsvgTytEjbauCGMB09ucqBBFrBidfdw75It1mY5s2z4
ZhDoDwAf4hoOKdAp+zzkJL/sIykjHLw18e8PWKC4cQLkRbJNEBAhxP4heKtU
Uv7L9STqpS9vdp4WgnhPwq68Gt4VZi9vTZAmuFoYljeXS7a4leJvBl6AD46j
Ix4e/Za1uQqtmRH5EU8YXFKEJU3QeimtUDWoZmeyqghKQ9DcC9mj0EtFDBeN
LwRkM3aSSMRq9qF4t92x+wlAbHQS2Ro3xNusS7F6/TD5fkGH31C0pzEUrm0q
mFRWfE/kWGo4mVIWs7aUZos7LimnLqOX82e8aftvUvgdkUO2QSOdbc1MtQCU
xK2F6rRetam9WHBBImZ6/mdsecOSSzewg22U27Yt1wXFWMAbRQASaOpFqEoW
qJXBO4BQqjJDCBMg5o532G7zvcVxy00sfIhCsbNTjJorRuros+IxExZoRIyY
AwfcgywvOhRZHmZVsD3ZwEnpI6Emxvbo+ERw+9sHHyLAlLdoU5e+u1EVXgwt
Sd66TcyiEEZW5C7JCPX8H9IPgABwdZhlWQwnklzdAKxrxz6VeGtN9dSURsac
75gQkkcbKI9yU/PsqhnzUxeukpZwYBdaNWKEjz9CqpK/FX+NZkzjfHyX7PkZ
k1el4BfyucHiO5n8jt+FlKZwlzBheJT+MfWrJ3eJ1PQKSE2Y7NR1sXlC5V+6
bFg0L53yn3HO4zR76RK+n6iTmVys+zznKpoukh3LK0um+Q0zgKX1gnGXrEDA
+jbcSaDCBrF+GyIeanqPa5Uj6xAuE4ggmzuzP3eyh+XO2c9hEi1FpFuTu8Jq
Yb3SLQIESQiHEOJ65pdheTPto+QZhzk9Q0ktVs1qWKe4RJuO2FZSDvt82U/E
qiH8/2dg9BTRugPb8YIuXOWRWEkhMYdahcgkCDI7eQJvaCurO4bE+0BxrGSR
ThWcO9P1dssHifO1FaBIG9n/QCmeXA/eJLtIphSnY8GRpXYimGjsQXrYSj+k
K8yGs8WwtLbeALe3155gFA5y5KJDYlygZ5B5SNn6ClHQ/dPszbskSs74YsXz
Jdoct6wRvlI1dElpyh9LVrw1hyMqR8cwEgjrQQfg4M3Suycc4cm+0/EVnXwk
XlzNHq2w7StbeINKsdEbPoCJFOhR26pweYIDgqDUfBFB3apY9DUFHDzmL0kz
nlcEntE/w49k+oZ2YS+s68b1wbF4D2fopMzAYqU/YLoir7VQNhL0HzZm0a7F
C162XCuRIEHFrZLz04W/n78GJvDDDu1BaNOopA45/YkmDb+VTV7B87h9kQnC
iB3wKaAzSHnlUGRFqPQ4xExMgRb/vqk0ZZupdVldkQF3Pz0Bkt5F1bQCkwsl
BADzqS+LJ3mxjcJ29xvJT/eNvPrwym5yOVIdR+ecP7oDHLs3kr0GFYHT3buQ
cNg4RQ8c/4VkeLx0zd4z91nm5pzxyX8fBdoGCx2Y9+RJKz+gU6wKlEpkPjgk
xST5Ig++1XZJV95XKHB4/BOmD6qlKo1sQDrAfIpCaDeLVU4N5NHLknhpM0qt
6XopFul2t3G7xUX+eGSZtcXYuyeF65UukX/kmHqgkI1dgJDdKacQrX46pTF/
Zvc8mUxWNIoOGzyyect7N+CGHQNtBKD1aH1J9ty4+qK0ZpQSnEifc43kMosB
Wk1c9VqrUhzPBi+gY0DBSYvB5YtL9wl8VYC9HZOBHcDmS6YL+opKqk678FEd
VkVr5uxDUa7qivArZOHmAVxK/4yLf8DcNM8Xhh4He+bCbl/DtfWCIBq/fDfb
oxGIom4OztSCcqjvqyW/khOdaREuaa3xS2hBC+1Q34fLAdV++wXemRZ5KABS
CJfWdQE2kT4MTnRfiF93SJbK/pkPSDkfCthR9M0dlIMfC+jyGX4BqIPw/2t5
3PnjVj7C1x1pIX11Gd1LHz0yqH/tInLbg5BfSZthEf15PYlNC1qpycDzEqGm
Ob73Yp7rZOcXy9Sgi7hr26+P6J92P1zIxuHtChEiwEC1BrU8z2+kzj+o+cUx
BMSMQcfxtnUer9WJp93pWfBJeDRDcM/hfkYXp888aASDPiVbduzTaNmfH8Ab
n22K8JoPI035Rhoe1/cZhoUPVeA5RJz5q2fUw+4tYjaNTfR8IukLVHt+Eh7v
vXZbFK/0Hv3AFyArseLx/Eg4yLUmpphnLdlLl0bm2twp093DfINEnDjWQmXP
Po7r+EQq03R4jjSYMqIDBOrooWuqRIGADLlqAG74cM6pCETFtTIvQX9akB1l
8c5RoPlDpcQbQpL4Bry43Ta0062CIRA4LFvQel4zwC94e8xSe0QhtekaLREV
mDxEzLe8ZtCIg2lFlqm4E8Foo/McK7cg9A6hSNlVXf90+jfa7tBeOeV6blyX
kHiUjeT0gURTE/OqEZ1uyyyaBIfMGSKJYISPL7cv9qOkMs2nnPASA9DXVcbs
4Qpeao6DYMUblLRENUWo0AG7UsM6RK0XfAykp0dk87UqmtDNoUZ36UsGdDD9
g7H79g14EzPZMI5nHOYRwhnF8vdBCIzNxw4Fh7o2udYfBYig/0RPQCmtqyI+
U+E+OpusS57RgNbGQ+tzXY2pHpXlFYbgKA5TWKMnoBKZ6JuUhYOf4Sf+HAgy
VPBNsQpF1vIdl4V1KDX5f5+RYH8T6YvsDv6F++46ExWPhdWBO3yrNQyPeOg8
gyj2axdhUn1h5BaevQIGk23QA7O/uhYeI7rtIcmgYR7u7mROhFmsT6+ODRWL
hUuTyaMGIG5ThzZY2qU4A0LnZ+m8DssZ5Om6jJHnX96ur/Y9vgfaJz1uJMs0
A2Hc24aDw0AMk0pm2Bve0M5MCicxBBdDlVY0syEgQ9qJXdRiFoMkepd0PDt2
D2lklPgTGu7YJMBmYyOWE98OH649RnxVOIlNlrOEefHNg8MnLQzxe9RpZxod
7xl/nOoLAmObF71waBUp1L+4E7u5mLj/4PVVfBMns93aMV2jZg7vwe/89gfw
pq8+I+zh+h/sLN8p9FPWTIM7M5pzTSVtyAZD2BZfTNcJetPEFFZPmp2bOCF3
EFF74zZmI5jJW6YSIrWnoWVKK4deFAtP4vn3o+8FAgwFlSd3Dq/3iN8rObAh
GmZ1OKACCz+s2koEkimJl1q3aTIzsRCpjqpD8aAdM8Udt1SEOj0N5eL/AJjQ
ToQdKKB5sh8mP9DR3OQGTkRxZh8DAm4lqoaWeYU7U5jYnEdk9gcUJEPl+onD
adCC3AUVWuDqnoMFyrvyWXv57FiKMoV95orKZFLeMq2W/8RV/KQwhhYedJHM
/84dsRhmtdwnINTPDJiINN3UQFQgEizY09AzYneb8z2MxSoWYGFaqAahnxnr
+RyMYbJR9+4QUCx1OmD3lfzTKyHJF/Qe8OBZn5CC1R9MaBJKCJZ2ti4ZowbP
3eSJBPUCu9xKJbAAcBjU7DbQqdIn0AqDIlk1MU0S6SxKhI53ZSAQOy2p7itS
agOCicGNdtyKVI8ZP+galVYWx4M1DxSPP7ua0fDPjv8SEyREisSkU7gIKCtt
a4WrD7Da93RacxKoLN1OCFRFBszkDpK9jRSmLFC7BZWvXTF/MGwCrusBTYYs
cROqXlCgVEaAwb9lQP6tmv3KCdp6aivDuZllBUkXcgF4fn1nhruwlZ6BpyiV
2H+MsAPRhg0rQKgokeJzHpu8nLvJyQiDMTJrdRvaywnIZOPpx+ZFFXs0yozv
lCDbSy+KeEpH4o7x0r6hDc8oHtBqgyJygL4bqlJoeTLuwuNk+dyyeoRGVhcH
G6+eZjPZSUgn0qUfYujmXF2w71NVPCzhGsO0DrehrWScNFF3lwG/8PU9eBUw
vWszF6dGc5Oeersg+KjOpWrFLc05zgmS4DDKDbrRzJqzE88lM90Ydjh2aH1h
mjmka/Y76lB3FOa2JekX6V7ri7y4EONIqnAo4RIv7hnPHc6qip5BHmUr8AOZ
fs2JjzJI4JqlpLDFTRfJ9bH2zR9r2/82Z143Ivke7QgZ+XvvYZip2kMoOZ+S
Kd1m7kMKKgTozJW46Eh3izYvLkplRXr/b+AWa+QzXfKu8dGQiV0n4l604SNE
jPdAUbVhZqDUz+RccVDTcI1iqlq/M2Hso2B56IfFDX/9RvM/iYvU/wJawu3q
UsU7Cs2s2r60rLzS7wrbDXP+9zM49iOmdylzUElS7qJJvKtDd8iuXexVdLGX
13zHqTdJWvEgKU3aJx/ziAr36HgLqevKfK4oTEbpX0iEizM8XQ5/1yaM/a16
I7uMvDIYOEkWOpANh9fxK6YeiWwpZT+qq/hGOJJi4wOgN64Uga8Owmi6O0yZ
jPwmJ3QebjQG5a+3TmfJASdpJDA5tYmhvJLzaci/r2HZiIVnHPDHF0g3PpoP
S07V3T7xXQwAQpMZm7xDoD6b8jxs9B31V98yUDDYkSdurB+IERjmVGAZAY4x
sVqdyHmDwCH7PDqK6wDzP/PSQsrp35PzRgUQh3tW04kr4N8+fJwfi/ZCi4lI
39BlDh00yyjPsmGiFLqsbMTDK99mhQ9LaJK5x9PJn8df1dsdLOdu/HguIbTV
m71/WUgS3WShcKS/NjYJ9B4FhNbOmHNQPRLy+aQ/rgKsWc66r/NoOGVIMVey
WmdnjCZCVrtX7EAoPRNmWeMesKF0kxcoxcqY2X5bt2tw/q8efxNEELhgdfA6
uy1FSGEVlRykRVNaMjpSdmVgcG0U04kl5j27a0QdZtvldLvP8pwprBXanIxG
fIYRLBde+GZj3Abkgq9hqLJapkmCzhqLA/AWwFUPKVED6lFg+qhf7tULGGnt
562Nsazpcm2BoRNGp/qmGHMHINn0KxjXlRfEhrEn3bI32UkIwwaxS+NgZT1X
qPrvBuR7JGt+10SnsL6DmjAxu+9exR6gk7S2cScz6+GHi+lur0KIGIiVNtDO
a5V9ofQGNQNX04AIGaTRE5xkYXydHC1V3ZSl2+SgFvUCARCpZ12+N9VVBbyI
KaiyHpUDsuNbiUQ8+4s/H3SJHYd5rDc+Udh4oFV7ZCAXZWroU3gaFAo/4n6g
RuJsBVn8uFV8MIHJEIdQycB/jIkB0ydDEtH2NU6e/KAl9qpi6rLj9sOX2ao4
Yt3LN5Jc8Urxcb/t3jePjumEafuhErN5uGBnnlWfmsdQmNv1W26R6KFUdauv
lkzAnrqhTJb/1R4o8CaXg3iM4I4zAr6385LRVi1TmUGIxVvhQ+DmbyqhqkcU
nvOtkMDJst4ca7csZ7Mqr1P983v9jRjPP9tk9d8ueZ4GTwBQd1YAioQp/+op
CbDS4GNHqRCyku2UkHJCv9LH4t4KfRd5+QxXby8FPMEtkHSlkxdPCKZKxPy7
ZEMAQvJ/YPpZOohft3YO8N2fA7fsXYo2+hcfYQYTV9db4A4oGLDNmTy3HSCE
nit+6l5ZwO1gWw0DFDLvyKpt4B1fGNkdfACIdOK6M/JGH8KoKBGkyjWuJ+UA
xXPD6rAedIattQZuypZUoJu1OrcsWTsCHA9xi+4Whogq78XLjeErTGXfbRhN
M6zLB4GZoVXgsViidPpr+lM3rlEd6bCDAyLgv2m5zwAyaZ7cEnbvr6E9zAbB
HAGrFci1khMiefeklhchM9YeqymBhJ3Okgh7C3Ple/f7MQ8Brq78kkMr4qs7
FBBnjnRCyLd8KQ+1sEim51RN5v2+V5LkE8nWUbb8PwqIAT4lLSDdwdSRPkCL
5q8/ZSFt3nXS7fH3uRZEklfGR0mz2RxsXMoeWhTri9PXX+LScZC5YTCdgfSE
czHiL01Ueiv+z3sJLrYGjgk0jI8EprpYHXzj7bpDcFEMQjUwzRvngEBhHT6B
COByCoUrV1RCooZHL/2lRoBP/TDDUYAMtjBe85HzfHimEBNTkrhuV/4Z9SJg
lir/uWjCPqo/Hji+x+lzeatDAA+NCm5X4oDaPsovING0xMZS68RK/HosTPS2
Rn+tRmVT7bi+62Bk5o0X0lXgdCM9bVYC2NLaYVi9/7izVcaG2AgcZxjtCvpT
1GhGjOcR7qpaZl8WbcX5JFYwq0ORMTnXpgUk9p82i/I/YP1zIISEBPF8yesJ
2YJ57kOfHu89IIMR+yiCWAv8mYeCH788omqE2aNmhieLL/ygsYXKpI4UX3zO
IbcjBJDe+jvNdri4dLR6pcbkXiZzJmMgxKyvALPkUqNG2PJwVpdNFBa4uB94
F5sjjVrR+NIIhwQFyfotc9tZgiB+6SmRbkUMMVZOkeplZKMDaeXEYrbA8juQ
Whbibl+yee7DHS/2oD3zxzh4z9bDjJdbg3gILOdpt+5PWktDlggzbGjnOnuK
uPRSmtxieMQi2VJJEXtU76uxDsQc2nv9l/6mADpTw3Lk15IX9fbIBwaE3Uox
S8Ij6RTwkQixddmhngvPh8Ex7fybG5Mr/r/pxTIg1WADeOTREqnnIg3kCxrl
QVo31XLhAX0oYZC9bAhJmvbXx8mIe9HFt1uSoKBdv4V0uhJwvtrPo8miX8z3
+qhlP5Mksbi2WEFyLYbfMy0+068LnWauoPWFwU1XgnyYF0r2NzBL3xHavNXi
qBblYB2X65/DbaH4Z5B5aEk1CRlG9nYxquCbSpQ+kZHulrQcuUrLqur4sFYe
N0S0GkhSCRfnEEpNLIhPHMN4Xf+omeSuKG5yd2up8GhNj2spGQJ1teuWslPV
fr9VHyhAlm4MRUYkRS05tjMA3PpCDS7lP+0Jrs1kD+Nz4HLATMBQc7gyT+QW
326Nzz2w7Fi54ZFnFekjSvOZ+Q7lLXqia49gRvESilyFIn9D+J8JoFI2HH1T
d+S96wT4xMMrMHSkexOP7UMM3HPIYr4Yv853gF6rRI8u7JsOaM6uf1OhuOl8
JQSLd7qjnV8PHDiCg8KJ96kwDjM6xRen6W1eATdk/pEzEDkxlPpCxTJRX4Zi
kATN+Y4/9mho1EN7Zs10rfksxQBgsPZ8Ur0ee8FU4k5W2WH8TQGNBBxVnVNO
S7QKj6KnrFMAejDYw0F+XxTaNHA04DgfyNiGAhcUJ5V7s6KMMXoe0VJ96M26
jFSs2iohdbbM4JFymEvVJuD1jiMA4T2BKc8uLuk+PMY4j4xluYNNWR9tFZm+
VOK8R5e9hg9RQHWmfS9oU9jBxgGaeqNclGJoXNo2CBSCDIry0Z2ulG3aTII+
N1/bb3F3pRf621xb1tbiAkoejVjssqLNNKSkqSqtxFH+iL6rHPANQSQ1tOjU
0UIuEo/d60cdvIejQ/6OE5WA/aIWn2WweQjDYkg8W/odF/m7uNEdFlgmG00q
vsL17f9yKHhMPymI69Jgr/sHHgLJTrWvXAxs8MX1ONzFYh9uBIxUnshSMCSx
mDxnYguMkYCWA1nWnANnjSativy474+Vjv4GFycGS7uApVLD1KP/0xPqEkMe
kYm1i0UttP30VJh+zOnJn0P76O+zsRonIXZsPdksFwQYoGqSfGQSIwOnoxMA
IK8ju5/XXXiQrIbM80++s3N0G6HyZ7ILqMIJoJlYWxJfgNc5PfetL4W5f4WF
eWWcOUXIvveaDoEcIZYLFOSzSof2II2GttC+li3cEecEyxEbrHgc6xCeWDXo
+RoWSRFP7Uu6BtiWsWBLDpEmEqiPJbYf/yPBbHZVKX7Pg+QNruH4wn2XTUiG
hyY8oRygSXvScM0M4WT5xs7dZlQCvNj3c2NorC5i3pPquG1h0+jthe+d2vVZ
fb6vqpXWcUr9VTH2R60ugDYrk6lPioJxkcNtSsKPn1ImrXwqtTgWkvUhwoLi
BM8anHAJi9CyK/Gi0RfkYWrHCB283MiNoMna2DymhRqYQIlfzoc7jID9l7we
aJKHtyQ3zmBB9fdu9/66x5PZULBwRFHP6971jfyw+JEEWx6/xRwBHYWW00Iv
y9FSwCsAqNPAC9sB5ygutItlAy2N26J0VQVFm5IW5O+kVQ9b3WyBHKD9gybJ
wGCrfwuv812O1dz7tj37uXZTzZ92GmbH4r1FRwEaxr4/M9tJN/U7sAkYIWeQ
aiGgKAMYyHUly83nPfizkAgAmiT3GHWPQaKTlXunqpn5TSVpEvm58NkoB1Ea
befkJ69NHccvayeIdlUPXJJ7oYKxy0gFhXj2VL0Yznae5jmMVAIMquNmUShk
B4x6TwC+uStStWQfo5id6akZGhwSauFlkN9/5gyC5GKzAo7NtDsbGitWMe6M
/H8TElslNbmou2ERZcjtI+T1ELrpVl5hqNJknh6+A9/aW0RIav1JA8p/vNu5
mO4UjJfdNEPnJWKM/jNlNVOZ5Z0PkZcf13sez1LQxvVAphfAItZr0R7Uobjd
EIZhgKLcH7PDdc1v8UFK9G5CDIR/5XrlIGSMu+tFUcw0KuwxIrASQrGzHu40
SH1A6DIsUcd1zHIOR/r8VzMw9jtvGOBGGkm3ZYNyOUMnGgmBp7lpJQj8aFlz
fmjondAPfhLBYPgbbunNzjY39nkJT6C/o9R2HQWg+9SbBlsCN4xqt3V1em8b
hptVs6FL9X2vQ/bpYWMhqn6jO5M5eTvaAfqo0o6dM0+ONKCgjbweSHliT2OA
6W581Mi96eZPAQO8qoZEO5Kj57P80p+0Nq7L7bFXM3thgK0YN/TiriPyri18
/GPV+N6CfERkBoQIsjFlw6J7kxeK4myYMek2VEMOSlUsGWEV5wA4vXR5HO4G
FKsA8pmnZJQgI6S6v0dAuLun4+z8gSB5dT3eWFZUmu9rzEoq1Wm1dpeG076t
iU7nUmgDWyE/CCEfeCIU+U3ORsMIlDfjNNmnn+5mbJ44jpmHb4nQAAJqw5NY
WPtKaZRdhBTt5hGTeNAiyPhumc8+PwjDlpXGg4LfSUQQzgKMggLJxSa6mUZa
dRCmzujMoIA4SAdQpTgDRUlxQXbF9chsVNGT36omsKfaUs5kzSW9qIOp9UJ+
rWLj32QJZpwoIeQJo2H/keYCRIVe0p0lrnrFt8rqhrTiFESyZq+DXg6PkbG9
VjPZgkmvZHWZpjYLiq4ysNvn/MveHismPTrZvLwmk0hQ5ig7oYNjjF5k03rD
v7cSYarbhgwoTBoJ8EGngzhDP5RFCXE5LKd4EhoHDk7A6aCBoXt6rtLjfQwp
xysbV/JN66Tga/iK+7KGSIqLq9IJH+PKcRxdC3bL2LGMUlHd+SL3R+AN8DNt
sGNNLg/epoOyv7BaWatG+DS1qiunClFSH8THUtVn7d7tdxrOZh11b26PRuy9
nbn3aWG2058AMwj/rO7uX+hNxULUu9OFHgTiv5Z4W6eWc7l9toIgkqDNu6WY
O/cTK+xhdKMUDcUqEX4vXeByFSugwhFeC9ERcpRpGWWlnVSzhvvHwPYHJs8/
DcIFpDq3eXTjd3dW2aYW6Mbp7L/BjbEnt8+fn6zX5iBqzJxmzMKhqgK9VeFB
2WMjyGIakivKlVVeZRJnFYjzMvudqXAszMt/wMULwBk9NHsuupJD7T8n48DE
9LUJodCE3PwRKeNtQiNwWiVrF7r4/ZW7kooLlxPHFqEOCoLOQj3uJFhJaH9H
/9tSivmBElvy0HMPF63runWCGp8LDqFb9/k6tzCm3cAqjcLTDhJ1QkQwjHGq
ppIoxzTaExjnlATUvNVGSV4mPbJpZmLMBvJbBhBmeP4HGDEEwF8vuC0DTFTU
PHT8iO5uIAoHwOhBzlEYKnisq0hz6YBuELI9C0w7S2AOlcu1c/VKJoLbrU8n
vLmQPz4whLb2+bgoYnfzHgnoJUofsbeO2csf+4HpMuiJ6fxtd72AML4QHrEP
Z8XxmPIGIHHV9/iMwqu2Wbe1x6piBE9nl9Gg0avIQsYDieTyZZIwqhfD0Der
RRtIITPW5eWShsWEyEsKRkQ7G5mOmNoEAVWptb57/V6KBUP/YzhnRKQLdSeP
id4a30/OIIm/AHS7tKCJ6LJb5Gk9cOcevIpPVQi3gHBLCkUzYM71XN84eO57
3KkJTsbOeuu0yel+OuxCv4T5CXgIflucP4izfgntWUsRdEQtJzmIxAuX9cCv
tJ2+zNGLYfTIgjQyQRSCDHxqOC/4C/0tWdkI06d1B27403dQ4l+QY6ug0O3g
0z47Dl6klFtMDsfuVR67zDQG54QwTpJC+crUjd+tCUSfZJYb5DtnTzuRD+v1
Xc38YMwT5avDbmv73usxJGtXKwZawjo0JENlLDOtrHuK4aMSAORniCiRi7wk
FNOfNK9Ix2o/O4XWIzOshirTfrrw2M+sRlIQyoMfHn9jCrA5FvOYBaSmobZI
0svsAOg2byx3baHqo+FZteGFDkopctTmi4lgiddMb7kfGOIWWNanHikKvzmA
8SYUBgSkljpFvuDe4e5/lSdkLb+Fv0seJy16d7HAMVKZWEBoq6pBrhXGDeNQ
iHF5BlcXjLtVbDyijjOdZDnScr7fCXEvW/2ExdsRrWDDHe4qL4Xsj2jn2jz+
iDl9TkswYptruhRheEzY4DmmSY7L2m37IsUtYVwQnE2lzSS8tv/aiCZDLGVG
HUURyUBvlSu1GGAhgR3QjpYthnAxXuMfNJpWPe4yzqdAsEY5rOoFURGPiGeQ
IGnIsenzm75c5UKfaaMNpWfWwwlwHnZYvmTwKJ7i0szIALelR6LLB6tsCGhJ
McgUlabcAUaaEr/cMMZsC8UWbyfeklx3EMwE/B/TpacHmVkDVXWqfBTR7rLO
sDsa+GEUQU5qmSi5CKXqhhLe5xOVSC8sjcicKyRxPjYnRPl9RMfD8UvTFPOA
SDtTUiKp+X8iTCsZry0wB+y/J8bk+3uGO/sIsCwXQMEwpMZr1zl1Jzx9bQVB
MJ05Oc6AJd4tPwNFd5NkO1KFdHloyspwRR+bs3JniOpIiQGMdiAMdieIHO3a
mlfmdSKGM2orvjjSoiWCnWpHo1j04GSPvp3/tUgV+R5+MsNwbUzkqi1rWo+F
+aTUHoAnYUwXwaQCz9qkSw8HRlasN7kRIqz1OiXWz8Ugcl6XkRiPGNbm6qtV
+9PHF9WCP8UE9vUHkZEt+9NVP1l/4qaJ5LXnK0vx490TL7KzFZ6rKiYZJv/B
pU4MF2pJh4wmeGWET2y/uOBM0UxdaNmiBR297QPL/hAxanI7k3Qpjym/fKsu
SLe8a3+lEm6q31FJ/eOkcmWOSguTJl7AjCJWRI10DV453bmsq2y8FPDC7j75
xaZTkVn620m+xWHSKUjMUb5jKFc5daEScYYRGuRN2n2nui8QzM62zwL7KUsK
1CPZBbaq7SMp7VqW4QFBQlHlK8L7FS9dvFOTkGmbxzlEh4CNUkcTKcOkf9h0
SYEVOKSB1/PzsrkJssys2bjQ+593ist6HCmBDNUud1GpNPi82MIWK++Bt4X3
AbrY94iP6MsHAeUWUf2MVTB4v6uF0cf/cITILCTTDXiTuvRWRN/P67pWdZ++
d4Qc4UnIAIW68UyOiqBJHAXTSKEuGAakuCNeEQ/uL6PkHBkdTYUnDxax0B9p
fo3S7Tzh5wgklanGHtgxRw0Z2/kZTtH+9lgGKu9Dk0cLoK437U8QBv+377b/
/JqZcY111oeb2a73FUZO7l2yM+0IFzmkautvFDShLxs5oHYA3shpSsUE3rdi
/QdME3k9slDrUl0SnB2lgBBdRzP0jcNGQmsJj/oxmX6J5YSiyoWSAZxDpveZ
rct4uEZw+VzTg/MMoAkASArIjb0Wy+JwBRZRVLh4HZnE6nX2JIe0h78Vpvfm
85n0wYDH9Z5rL/tBPT5ZCWLHWP48/pS11dDJJIjQxXqN5hJq+LE1mZeHOd7o
l8yf93/THVLL2CE2RWpL0Sy38g6+PkOc6UEnLJ7OCEPX9rlLWgOH6PDQHZ1J
13HsSllPJ2ilZrhH9kXjQU78P90oPwqr0lKZT7UAjdIf66pbuRKFCKdUhS4n
6A+hQ38pUpGEA8DF6v826vMKU9cId2AkVc1lJDcqBh+y1YU+BvHGwrzskbSp
83wh5OWJFhpdMJlf9e5gA8WitxYKw3eBFV1df3oOzGuOxbVOkhxOdcz+UWTZ
28BNPeP5uNjCXyzC4A7WtUZhTB0xnLyFNNWKWKgEJ0nOpd+AR9VUFiMoIeXT
6E4pxH/Rs3dK9m2slV3N+9g+aduoCmxLsQ6N1XCAFu/f0ilLroLXTjG1mUlu
97g5VUTmYGsZJULrHhdNACvhoHDDUjBPPiAtJrP/oXzXTBnlBB7dhUs9MaUh
HyTMOHQBFggnZdzDY49BHWCoLsSPwsXl25n9RNKR6Mb4H0daMId0+Uhrr43b
4cHxeJF9jkR9vx/NvLSRNwA2xUrQ+pLacssEbhnlSI1LL/ElXYAt0mJOBs64
Cw3/olh6d9ear9vXiXFBPqwdG4v0hlAIg4kQ0QQMkykde7Dfiq0L4uErhLGO
/sugFMjGe6wygSDWBmr8Ai/mFV8PSFk672/qo8nJzKTVESuBtS8wrE3yLgvI
N7vOTRhPDEd18S4MJ0n4t+UBXmXWUSY4qR6x2cHIfd48Fr1ylij9L2bqUjBj
npbIKIQC76T0PhOS3GpfYltqdT36rtUiEyjA3qt0ktZO8vBt17okPKp00w0Y
g5hUpB2Jc9t6haZDMVhqk0La1ATEvdr4UDVs+4WptpsVwXgT80UMqNoqpCc0
dmheqmXAiA57jDUtIGlYdK8c4wE7DffagW/S7iYGkRxbDjWhiHlvsCNFHIi6
uTU5sfyb9DkD/Qz79NAJF/GtpxU4AcvPr+XSqNFuQaPBfybWFiYdVXcgiRP8
Omi2/i1waEpcCjsmdtKDxtyhpqOL+ig2tXAlnjRYQIpzUtCqvTITk4v06KYL
cbCqvInFkOQ6Yuj+LJ0XPts5hkelUTYlfqlEbP0qnQxYCwis+9xJOxERbNT6
r3B+0dkPHMUccMaLO2JO24BHN3BhdMKbnOrORi/lOEnMjinNCmjXoRVOIB/d
fQCis2qb6pgXq9ArRQVrLEQDsjzb+9lhiCydV5vBGS9WXhI/+8DuDQFBVoC5
p3Fm+eEFDltA8h1sWsUH9+bWyvKYcWp5OKhftOTiBwlvp9ym5d+FBz1ox16a
srsGXA1zt6F/IR1EwyGHo3wnlHxOdCS7ZWkTtH0UAJGs6GWU+8EGTBJJF0yS
acLI6DiQTnHiTUG2xEKgIiyKj3PDwq1nIOFXT9luCeF7gz1EGeqRRjVpaV1z
5Ew7iWIablWaZXHTZrWsYOa66Vc0Ul82CZdf0xYdPZtLfXMorZKOR8uVPUJD
w4fp0HVZFTCmgxSX5+nY/n8RSgCzhdk2win8f7BK11ly8OSNx+AlJTT2drd7
HP44FJGs6wcT2Lh4HhwSQL3qAK8cHj3Cv/SSNCgF2zr4tWewS4CzRavM53n1
jN6AmFUOMbKwJnvu2cU7cYpLIQKS2TKgiuyJ8ZAHLj6pyIGZtFXG/HGGD2JZ
KxvLYD0et6n7jJZq2h5i3SSnj7FMdBiiCR5PGNicDJXY1vWG5bDXzKN28P+b
3Qa+GjjAbZhCkJjwX2J49Tw7udgaOfe3WnKRiMz5SsuGp2tGeitUO5e8eeeE
qu75ColbYDooho+d9jShcsLPg58zzCVOHbwQnvGqmsrkEwKC3xeMDjcXtZTT
eNaPGDyQazWKj7NOKRCdjHaXVHd+RkNVvkpVxdvb0b4e6zNbUc9YmP2i7sK4
b/IDo+bluX6IC9BqIpJPK56QiFIq7YSDzSMTLAWY0Mm0S9k6EAKyOg2d7Z43
Lh2iDv1BdlXyBaE9YXwjPxKPEE5tXZRRpmZe9uz7z7dfr5ieym3UOPP6U3Iu
GG/6Z9GK7jXcODbr9acK/AY+d/ujyFXJoUMj8+pGeAsRnPnSWEenQq/WerHb
nDE0BxMRpmOMRzqjlsgX3ye+U3q8CmMvczy6EUjwZgINrEqv0w8vRIaWJRoZ
0Iiw5z96TaKEHzY2UBVzNZWb+/27FJvHZzK2DE4QDCvM/qIo5c0lx0xMX7am
QHKDuBW/q0bv1uKNNLg40jwCMYIgF1TgIGmZiORSh684AnoXJHihwqJFyKxq
zm5l9a7uXQc++g1Y0+bcybzEJae/Jy3VV9NCeXHVATWqUioNlQSusBN3Ddo3
6VwC9oTXAHMnvcjcZX8FwTWPVOujJS/KCc+zP0Z5LI3P2xRR2mzA6wfAnzbJ
E8oQYcHN5fOP5bX3EDsSW4vXtEZBTPtwmKAOc9NZnwwhLBnnwXml/gMiNvaM
dGESrCpEKqgQUuguIKG3BIgcCl7oYsipwH067L8EVhh1O7mWBeSOjpXb1v1y
vGug7pJPVk9CSEq7F0yZOqNoWdlxWzmW8XRO0Cw2laBUieKWxspv52lN0mRV
LvgQvl4PUweN1hJRg/XNYBEXSPpvqxkNQsPu28xkOoyNnQ5WBxF3s9Kj031X
suGVXEEugDw+Ckf1soHcHr3eDlXP8q0LFp8qfDD7klN5fySrenf3d+7Hi6kf
ntI9YVDZnnw2c6Xq0x2xO4b141QhEGDCqbpxAT6vI4FyqHZawR6/Ds0wCApY
U6Hra5nAZYr6tsgXmP7pTTuHDt8OtZ9rKrBjm9/m2Q6usMWkQaq/RSjFKaeu
VQAVqYlNLfyVXrcKzy5FcGHRn1xqQoJ6pGU0txSsJi2H8jAi4+aS1TnGypwX
ifUVhwtuGwu/EmYhGIododInLMMgIqJHZlOtsv51jDK8L8L/SPpi7o2lDUB9
GgRcd965FlJ9xcfPIUjVGjHpj1hYi/Tr5VBUqUNYY1QD9HpGssoJPAxYYNiD
CdTT4PLLi2+3A9Pi1ywNH+4P8BxEN58memaXnFmoi42dsWuULtDTrWZK9K7Q
CWqZRN00ayWyFn84Qdfi8gcghrTsOfazW0FJ0HZ0ufw9W8iBaqynd70Psz6Q
GBP1vAzgvkHXVStusPFylD4ZlKFyoX8HgZPRiRBFRE0Stke2KRG9sUaWS6QB
sKZ/o7B4IHoHsi17WswUduvOzxWVsW2eKUlrb9xdz8+kGUdbThNw8Ddzqy+K
1gfd84BdmoDm5N6ZsgDbNtxXxJv7TBzHKDN36e90muD8J2oOupQy9GbDdFes
NaiEmtJeUcCmFcOTM9Dt4FLBfPoM894WLzuK9WhSNmUf/vDAi1ajnpkyuxMP
+s3hPRzD4xtRt/N5iw9RadR8xmbSYlHX0c5aaMCc4XlpkRRTGlJAW1MNXq2v
UHi2KhJFrWFwnTEVR/JKoEQxZYT8aB8HIQuoNic5LnxMw/3ct0JzQNvl0/dX
QhFJMvavgAa7Uz60ZRn/221BoK6PXL4h1ejyVCSf6K6F2C3HUUXL+d86g7Kd
W3gjP1YqQfG+uqymP/32sd8bT64FlB35k5RJuz1MjWtKhnh1CeuILXwsnTaI
GssHiWQ27bwJSOppdoUBG+iXWyw7BIrnAjkycnVpa6bhD0tEYyAx1eO8+W86
KgcdhVfbCh4Ku37JRwt4HVc6KvomJ8ZPQHQy54xWmgCfcAwW4nok818TyK8S
jwc9Yls8qVEHZUUCAUtq/qU+PSb9SdTxku1Zhv/eGHmS6FVGZ7o4QnreYyOF
vhLHztmJDK/eeVy65dB61ljZrUFJlA94s+ZsuXKWzwIC4gTsMBmFzRiwrega
uXdnByXzEK9/VVmSM7P8OHb9GE2lS9eJXo6S9LLS97YdzRKyP2zAiSqGejc1
lcGHAearBYJu4KmwJIfudFsO0WYIFkDLOkErhoSFbhHFZ9ERaay7JU27V3xX
8pGVIiz00g1ZqCWHPQI+Zn7Jpj70sw/Mu9+iBvgiWprHGTXhKYOjDmtssG7L
vYGj2SIHaA7c0ROIaE67CHJAfPulg6npx/rJlTrYSV11YB4sfYT+2lgRU7p/
Rasqxcm3W1nWaUceaVegOpU9z+8e2/hVi1s58oRJR9/UJjR1WH+7RcFCRPcl
/ytzhGwDm7/I4OJJ0c+PFJfuVip0naxAbBObsHZbWRRo5rtLwtCn5TR6Ja3n
b9lUIjIYJRh9+CL2Ix1HlwMNsjFqE9dC7xv9k91SE3uO2RCwFPZHSDJayJ3I
L+33rBWEro5myFIthHw4Gmm5SbcrYWQUNI/7/5hqdNfb30LubuNwX9zGHkBn
cZI1QRFEoa20WpKf2l5NMa90fuWTTnmN3YinmRg+VBq4EmOA50ZjOn9jlAdS
BpnYngOMWBwdeYQ8D1/AZ84fzjXz03HFbLqLe/66zTN4QE9V988oFNyr6Hnq
MC7MMFnKaMwwjKc0Cqm8lPHDCWUdY9Lmtwenvh9RRHE55Vtr7BA2x8hVnkzM
hVYC1JXFjx5AvUUP1tB6SvilMgEfx1sL+IufdmpYx9i14sTfvOC4dPbZI520
7h8uX+pMbInpi2vUyyTMbiRLzxDmMQLcCnmxbCd0y59i7SRRk9KSyN31oJ4g
oAN/k/Lj8vlobiwOZ6MJwweKOxnC0FYzHKtH2WdQ8n/HRm05WLzwnE18mzZJ
5AXE03h2BMu0rJmA64oyvuBi66ZYWjHi/yrm5sLjCYSfuaj14jZVLVTNbl3q
4jEreotvaOSUJzTmCKmd9mCEt1fiRiw2UwWcvJB75uRXW2qrPmNBWntSgCDI
xjdeI2V9AVC9T8sK1Rr2PHFdos+8VMi82SNf0TXRAir46DacqQR5UWPdJMJ6
6PVL6f+PIRUEznAstlX/Kguhn5sL48WzOYTDlHJivgfWJkuNrZ95JUK+MQnJ
amldKFZu9xTYYbq16ZzO8y012JiLwqVjPNypBExLAGcCA1y0rXto1gfkeFGK
F9He4LKGwaaFXTVBobRlbb7u0Ub4sfDwWHvj1QlOZCSq1m8NXyZSDFNNaVOO
sZvu7GGQdAEC3ceo3vGtQ8pxRYA7HtzRXVpha3PhplishvOAe6tWTQa9QD4e
Wxwb917KR23UmfAIlefZC1TbO2bVJFelwu/fvEDTEdbHA6nZBbitf2tT3ueY
oxlBmGakQ5gIIXtmOpX3DgXLEVyl9MvGqIx7O7gzI4Ni32vJMUamB6GtlLst
SSzMEFLTJsvvX3wafk9mL8q1QQbHDGymjrxv2mp4H5u7pta3vyYp0JSa44Q5
LA8AutgvAV2SVBPw3UvFwx/cOsGIztLoLcnCImsjJ/UKbOh+jY4EAmShaUfH
uVdBZNQ8IFJzcUr4DeQ6q9lyn9S7Rc4U/JdljN2BTG60+bin9GODTDo+hKR+
d/utw178NpdHdMf/1syzkGiDtZ/B3sW6VOyM9Wo0lDamregcp4EcldDoEA+J
eJ+V/UdEX9jkL2fSWjHY+BztHVb9+g0eMaUzjYLVFTysnKebilIqLvkZfVLQ
vltvIWChDZ7ue7lbTDHhYbsNv8nn2ujWnHMobPvcERgWZdfeYHJ1JGOLIG/g
LhA3xUd0g6x2QKLEcn1NMvpKze8+fEjLpHpR1bxfmsBKl8N4ELNM089R5NHR
b/adkXPFfPvVekNE7M8ZB9XxtpF5Nt8ogkySOeYuSJQIu/QEllm8s0FCa43a
o64QCYB5m2FxajVQcdgj7GWtNADWpnTYi/+6mj+Nyi+AWDdO9v7DEXw5r+3+
enbIC3Ealr07+iIv7H46mc0eI6gHjSifKAj7Q32xRtLrhWZfPuQYnmzgZ7rp
EX7XeydIcqOZoiVb2pzBMzbYqrQI1ImsgoNV0ANkrUcrm1RFCdk+1cjnnXby
QpuxYCl9hilYtksLfaBlhh4rRQecaZDzMd7FGySmCSQsc8WPhYkVaFxhYAY3
CmNAFmH1sL7uxh7vaGVM4lqA+0iSzBYMs697FzPpL+S7UY7Ezm4iJLtjSXho
nWT7ruuGi0BDcu6q5sg75fVKNCDk1SfgMfmaEYF7GIrDIaW3n4GrBAk+8eUJ
LzFdQiWvU0QC+nfbscIjF+9IYOGcZ/ZuaIKo9OC0kmD3XtlhA1QBVIoBg1Ll
hIL+o/ly80wy8euCVy2tyf9gxnn2z/c8aRK3dqHIzTvmhMbeXN/Y7ZaR7i6b
BLh0Pc/8x9LAzn/Cz9Zlt4cSEbewkAqXkDLssk2orkpGf8aiyAdEONo42YfO
36b11KkYeZTIlfCDVkFjGJo/R8gQsNdrnscYryXrXe9IW23dQlWBPZvEHetP
IP4xzJl1dBIMx2t5FlLF8u1BhjS6HHvy0gsDsZvZmezq1aIWrPQ0GT0c99J4
1C1xTesG7KEZfhMINcxCvCbr4SyABSr/Im9YHMHQAipuiZl14/6lPBj19YEs
PKlKxirzrkuS5ZLfkxatYOCEt/OcMvyHTTjFYiVk2TpZ6I5B0Ud+Rs8iKTw+
w4KegCb+OW1d8E3DSHegTCalVlGu/LH/mY9waAtJ57dWjgFHAeu5+eJ28ZDI
L1V7rtAQDjWlNupofzBiopKwYpXtQR8aIvTJ848Em2x/xEWR8hgCh/OYTEvv
TFETA2zstdm+NBCO5Jqu84maq82XQTU3A7vUIkZwFBo6uN0Niq609K6P2Aem
pOgeLeowmcBLG46DtUFDgkaQZeb2KHbBJN9siZ9QwPwfIif0CBLrZv2H+2G1
VnzmtNmhBAryY61NsNjuNXLx0uxQtGnM3fmvrRhwZDYFRFCVYAMus+gE4L7m
kWhKMmykbcR2xxRzplVGhRUiRYU2LpH2Mya2RHIoo3QU7bgEmqQDrR7UVe3E
kbJuIKwSAJU1LtoFdCXtVaUL+Kk6TE9aCeRMnT2cRl7eBPex0jaIXrdseEOg
/NaxXFNA7Yv6yMqQV713S7Zwp75+44qEFV7dV36qb5thXPjh5JAbeeTgcLeJ
JSmHker9SeRR6oY1PygbSQEMXvm5jDljrs/N18PzZmXp6YU3L8Jop2x9Wl0l
7VZLPyF5CZlTaRoohH6H/9nM8pREQdHlMSRS6E9zYam7govbuC+yfO7cUKZK
sg4ooJN+H7My3rVZ9x/ihuSfiEtziU4gjaALfJWTFXsEX6x4gg58zX67t2wc
Y+a+fcOIbpYRxATsZHNs0SynLJmoKOlw4rk/WLsPmMbnpAaR1XgBI+mLnA1E
/WEuug4fbYBTF7PDt4PGLgfRh2A971b3Ckwoqzj5XWvOCQRPrgIsczXOw5iW
13fmp7GmBaqvDhbqAJh9rXrck3ulSZv2p57n3sijKkSDoSUei0ako68k5o6b
Wezs0RyALyzK5KwzGbJb5Umkv55L4J+sLD6Brfsq1xp6cdw6zLGihvMOLz2r
DzBumkA3YA5bmxVFiOYjRZrES5fPVkYE+ZQbA5G8ZP7alMukCCnovmIAVWc2
cVE1+lgwl+l1SQMAT08kQuRv30u63g/YTkIbXs+eRPmIBO5h9f5VgprZhfq6
shSjhjJ8FA9OJglluiid5cKWy8gxpvzY5ov8jQqnwYJ16wjY6u2nJ8wMNm8t
ZKFqsy1wy73xklHSp7SHgIZkhbNiD+qtVOnuKD4ya0aeydiUW9LgQRnlUK7e
5ywy6A+ikurJ/ewY4u/rZ9rCwwkoUA9iPsqy9ZC7qEWHkwId+nyM2l3kps/K
uorl2DI9hNhLSJwEnv2Y0GtgbSjJrIIeTfFM0jrAlo4746pJeMTpFBJeisKV
EKPfGl341HEDMsLy03Mh7+xgSHnisB7xUP59kRGtPN35fnvq2nxvAna/Bkdh
+GJrLODCLr7blZyzlQ3BUuobysfr3MMUWKxtSJ127NCAbJrxTvzKOR6YDjS0
XNvAN2JipDsRnOGajGCsoYFvnL9F6EyOa5gd9McQbFDALpTqPdDMHxfF1ZzK
Snqus8F3zklPM3c5oQjaFIBTo3rMiUyNhFMxj2XhDSh1zTpelGE1cbETugY9
VOcSlqzYtWsGHGmgERCMalqg2VgKfgVlUcGb/j/mEk4J8Frpf4yS/ZPiM+zk
mFloFnHxMp2mU0Rwh1nGrdrDKB/aQvNtJ2jqfi/bz/HhX10wO+sK4Y9ElVaV
6B7+tq3T7jzfefSN71fi5nTgX6SBrzRGOiiHB6YE2cqnkgEpwjM6Wf8HyHtU
988IM6kfdFlhABlBfTCZWiFYfQpYI67Z+isVaScZcP3F+k0uNJRuINHVWbWJ
SGHdQ7Jz6U3HB2w76FesYEnXiIzGCQ+l2M9lnQ159IfEABsAmDgsZSqpzS52
nZMe7fZlu/Z/gkD4L0BWl3zFrhLPlOFfm4tG+6cY3Q/8WT3mxaHGsbA7w5MH
SkPGfMVmBnmuEEvS7pvCbd98CGUwDDhEjTsc3shUJPj8jwH49jtnRpKeAGc6
D1ccpIY1UyMXGdJqMyFlf7ggkqwVeuxRLMgq3w+J7obcEmtZ+VBVeKTIYNcQ
hTQ5Yvb2eVKMm+RtCsnaop/2c3OLvIOcSh2OlHjcZgoR5v19tW310fI7CzZd
cn9lky+4cc62BLuBkYPKH8EMmNpwZyMtt6cwFxS4AIE/xHgfjVDm0GIgSprO
j/lIUb67QviOEo8FdkQs+xB21MJCo+HDTm5ake+35dfZuUyiaBwDgwhFB2vC
GPAFVBApzvycire9JNSq2haYCi/ZjYVvAVauAGd+Or9ZgT56ZIAVqQZ/sIKQ
/Lgju9WvqWeV6knzv7SkYKVG76mrABw2MqritLDt0EFku5Cgds7QVsKlG9ed
3zuHjewUbsQaJnr2AfLSNRVveisSsUGjqf03qbYUPntyspWbF/BQ/7aeJQbb
F1P70qNGGU/ZCEhrOqA1B7bPnCLrhU8u78BIF9tjU5DvcbLw5MZdrHYbKf4N
uEL51LdWcSrTuDVwMdu7TYiCdAXPrM3E1NnWEPNVbyDomJzrDRuX6uxh+dRU
Fp4czzIv6Jxi9SMfI85VhR6qnc74faxKu0yDlXf0ndd4ChJmYFnXivxJGhsp
sdhTGpJt853LljME+a/VVKmkkFu3oT3uz1TYWmHETLsbCJ0W7MnF/+Dt+mb2
BLvbAQggxrR34nAhrDDjySH7vvzn6bw7oftAe0AQ/lJlZ6VyH97eTFmj2ihL
Gdj56aNJYrrqZ5cXuGUfMFzoqPPOFsxo+7BZgNjHxgriI7duxkJY65FhSinc
T8Kl5meltpZ8W+lbuaRp7SXI8bEw+2d4QPWnhdY7+qNtlXZWbXq+E4nxvlEe
TvVL7VSETtIf9waiGfnKhrRneAbEwmHYs9lr8jAoBO79dnMSdTJnwPuuBgDM
maWIaa1elkiRWrErLOeHUOrooBBo3yQo4P9uHU02yf0ZlD4IiUAlnKcVjqmq
STXd7Gf6+c56QvBdreWNN9NSY/GHK3P4Gb//r0LUg24UrWskPccYksQ5sDu7
ki31cj4EeFWmGwPwPLv4JOt6Iv7bRr5yxLsVoEdUef55MKSqG4h+izukQSBx
F13GTPsCUKGXaW1Nt6SESCAzWmT1vBMCkn3TP2iGHc395Q8eslMSakLXVoY1
7KYt2QNadXBLZ++Je8AGD7Zhd6EpI2OrTLhmzwHS2pr1rCfvmMt/fO9iqzai
QGwxtnRBh4xhythXr2Q0teipbHShapc3UnB3ndZJSNvAOTXibqunPg60RqAj
xc1OxmWxqRC785fQRJjCtJeN2c8lfayJ7r/HTQMfidr1Qes6UOYeolYSiZq2
wnOwJ4CGaLSm4+qWqJAQOejulc+eqBTEwYaYNzsQoOAFYIzDOD6+U6A9lRoG
WtfRdW326yGn36QzILL5V4kCyKf2dxrz2jwfth4TCPaYsM6gHdkMRrSQZcnb
b0RABx49YbL51WN/nL19+/TNvVTfdwgIdoMWuho4wlJg+voGvNy+7lmp9zhm
Pe+Hoy3pKmfYRQFvez8UMZb44bazjec+LNpgVKkAgqDzR9Kb/uON56IKiZ0w
7DggcpMk8LQLwpISIsxTgJklgyuvnpp2AVmk53QP8jf5F8H55VbHmbCz7ZU9
ElNN51Y/MWxe+W+5EywFSKdYH7ZxJF5IgGicP6GdvtuhwANg6VtjHUPnwxTd
8W93Q/Vs2mAiqvEYmZfp32XbN29fp1j8lPCTTyt6yFBBSsXB/kdlLFYcHygF
2Qxk/6r0yUzya5Se1TQA80EkD6uon1XBsS9cbn8jO9sEm607S8ap9/jjIcql
Cps0jj3FNAoduTs/GdycVheEWYyScRE++Nr6YIEI/9v2Q800yWsMM65qOMTD
XbX2sDbrKMl/h5CfFg+W16UQ4Xube4L2Rk8E+hARt/2zg6D1iYvGZnjEhwnu
IeaUnbkMXOzYINsd0rZmhgNgnhAE7TyJUXt2HDXg0gD+p4rib26xaCNXdEBX
BA2cKKMmsdvKXBhubRaoxCnTLWQERqER2ds94gq6zsq9dmJoKbR+eoCKl//4
48HydBTXCY2wQTR4VJq672PKF/CWAgnepwVl3rQWPFuOSpoOa9/3DSu5YlVU
nfXXlIJeAwIEc9GeWvYWP0o5BkQLtWjIg8TGsOoOOlC4Me7U69AjyTFUAyIm
/7vxynG0oaHpkHzQZwK9RdYkOpYmJiMcJ96xWoCNE54JzmV56mkmmkKddC8V
aNpKl9VwcRjxSxQruD3L5LCZXrhGKN2hmATde/9ug+CQdUGPugrvE430VNYI
83Iw+Mn03JMg7qH5pdlmfm/UR7GWBGzEckYSzZWvWQe38ZqCkmJrUMi5AbrN
qgWvSZsJEUJWAuXtHaVfVnPH9vDRJkZ51QJCS0QIIPEpFZ3rbTt4+LuGHwc+
meVNVQ0XCTqzJQQJxqzi1lNTw2IgQxjzfmRxdEblK9nMehOyHl6rXCDt3A0y
noVTRueeWhOAWuBC2B6nYCiX7KJKe/3hEPVuyLG4SCYa1hOzFQf1BMyRb1h9
yPb682bbufLMoixn+S8n3yVVwKIZ8AHkp17ngTSgAiHDisuBOAVDdLWYGhKX
Rxuey9CFhSz9iZb7dvnrIiBkZG/e2H7cxioJh/vPSSj+Xk+102DICaSglIdS
EYttYwKdGqlN7WgmRARVsDpW21fqKBXng86m3c5sIJXB1NP124/TpgxpnKN0
75c5XRzgQwKscmaJOFqOq2k0AevAQ1zETZRYhsRrUobrvoB5tn98Ag/a7iVv
bRgq/IRQ8/gE8s8mIuYEsqYGrUDAN/M0OkGYQ8WzUiOhszfFz8+jZFcJ7k1n
9pX1OcXL8IwZbhkJ2ADXTiclDLH5aR66PJKROv1Mn3qlqWDGNfR8Br1HTQRX
xEcglCAyp1F0syTCER2OLrhUaJxyLBMkzdEr3JoGik/3V350OngMGXPfeqX/
FsPoANBpsAycHx5Cyc17njgnN9A+sOpmImD7oUTpIxwHFqTQ0WnJ+mdid0wE
+4K18HG+2H8aN79XD+t266ysb6wijKmLhoV6xb8JFOPLGQ/OOFaPLRM7gEzb
8VxiWPAS6rFugJG1Jr6yNUR8PcDZffTPeTOdLOuuY02AiziF2oVx8e/ze7qB
CbgJCMfqdEVfXW6uitCrWE9BR8H1GZHti52qRbT57+ckKjnfyC5UhmOCzTBp
FACziwFZXY9lvpxn3Bx8ohwMM/jeCfVr2DsqCVmdKsr8gHD1Fgpv4Ai450Jp
W6bOqFUhC8kawp/k2SP8a5G+8qr0l6kaP2RjIaiL2yHk9bRB/U60iixludNr
g3P3+b3+z5C551ZPYWBcbLf8EIG5E20dqkIwOzX+1byGXhVOIYYFJPNiITXx
6KSBz3gDKpFPY5nrPPEmrlKgIAvTm7bvStovQ0GoFBzZewBNV60leI8sX/25
Eb4a+37hAiimYZWV4j9X6xfcTGm0clKdgknMNfHLrTPafbbb1yZ5D00N09ZC
oL1DSlG1STBDE9te2VZMZIer2drP0+n7G+0plQJFQguAqdbarhXQJVUoK7SB
rHoDfjw56XJhV/QZcWnGT+Y+He5Y0AKGztrrGETffYmCFSY31JVAK97Xi6Ni
VesHITSoB2muIFe04TJamnXeCo9nwgUkucMJCw31DhXXRRkIr9XCmTUwhs+V
7CHM2nNE0NbniIDsr/Bs1CAIAB0Io7tni4txdiKyGaYE78ldWa4eFvl6E/TA
VnnINcDe6aYxV5rOVdV3QyEkSdZ0F2E8uCa9Eg22AVQ60SVPjCbrZAY/p7dc
eIiuppfmwBmgeyamhI5IONj7d9qmcxZZwHCj+SFJmC5BAY5ezHb0+/zRg/rv
39O/+RtUXGjcojs97Bw5hTOpHVQ5z9gcuLAHqhOD8XbPFqCXxnkLEgV0sE2e
65EyZyA5kmxGw5a7YxhTZm0alZEONHMQeQazw/+ASeXihTx0jdC20rMDHL3d
KGjiR9SeEvT898MAugP6FmoOm05wUjFctPitzVWVu7f7XrU7OILh+T2O8UQR
UO7EqbY7n6fSIsDJJL3qWKA6jZj8zFdBxjKAeg4MpHlH0o+SyshwBoULTFH2
7SIk4NbpEPOCUlpoUCXP1Ut6dZT/gGo+d7yF2h+8tLDU+7Cs4+bNtc4/Dglz
1QTFapZjRAg/zOEJUq7bIBPrkD3ayAQAUO64ZERSOL5wGS7O1o3WC67+FMdY
nHrPBC+xSMRVn6JYBMj4k1c3VSWcAL8xs3KWgdpLBa3MfGLSNFnAu0ibrO8X
z5wChPz4zzPWiY+FM3hzFPEwRGu2n8clAEXzqrDbzexkYJNHjPJLyDSd3Bxe
sRIZCrkvfmqAyf0jMgXzyW6tkagZ9nbgNkOBtcZLwKTtguf6CykdztlOu1Fv
a8cCWhEnDrBO+wv7ifFCXY/QaXasfBbgOGNJu35lGzOdLFpA572BtfwYZPxU
JlkVztRW5zben1Zffgi+1+x3/Hfok4H/Zm/JKo923Ewx+kf0AxU1Q7CPD3bz
GzmASMjNXalJqSKStGhc8zHKwrzBVcTI2Vje5QKQeVChq10y4uLOziVBBVNV
yb2CwMV3cmZwc6whUbSBbEUZnCAMCqFc9bCLU6xT321fBCS7hC3kSZkqNlDS
XLPVMOPjxlAVT6RedRlC41v/JDTNQys9ZjBMGUu1px13kQ7rZYJ/PCuPJ6xy
rs5u7SWyVb2nfXyKGsbeSqVOEgfb9P/SPKI+nNxed78lWRVP4ZEF7/LhCRD1
xLkdUhMhOxaiW11dVOu7cYQejzxjZw3VulVIUFFMk8fzMXajQ3tyvHeIES77
2jtlMdqxfcuSFcNqDbAHKX1YYFrq9ZARYO1yWkKOz2233jirtXWW897WZdiC
vESRRvmFB4wtMZNCkbXoOgUp9FAxOJ5DX7ZvboCoT1Iyz2NK41qk0d5Zxp2d
0vL12PzUzd5SWp2DrmsFEcY3z/udsjkIPvFvVTJhw5tUyUPDlx9xat/+RfnF
d/WTIjmhFfro+l0G4QbzkBOsy7avyGVDfiXWGhb1JvR0HvKPhly9s6t6XNBd
aaamsuo+LDarMwR8nsIJoLfhL8HQ02lKyR8PnHdrce2OgB9gIQQBLC6ZWi8I
7gtRjtg44zl65Ci6uB57c7Wx9jOU57wWXy/MGCw7LTEE+m54cBkmXK1XqHbR
09sik9d8Jp0bsXrCNWK7VTRNDYZ47ObS+KZD2Lw5zf/JxkYHJ9dZcfdWFpt4
RCc5VvCJsufBDEDeo8U6FbwTrKzRtgfOHK6NbhHnL5WzV1VN+xMORKn/GcW9
GxB6UkSL4XVUEgeAhkYnGZMBnEjxDXyzHqa93ie6QlyiEdzvCYJc7m5Gyh6/
YUFawoxY9jzOEshCyQeYwPlsppdOG6kzNvdOSi1jzI6goT1WFm2dISYIePRF
8Mp8KW1Gk8HvjFLel6YbYVAlV8gmNnr+O222gJ+PWOZ8O60HzNB5zrqvADCH
WgldguqPJm/CHWWqNDHtKPrVR37wQgdq9oXFvHzRuMLojC/KYpY5UTQ7zOXQ
kI0+P5S99+orBnsNeEJP8a8tbCFSSLZrDxuRgpjYRufnmzgpxtXdIUGgmS9j
Ii1wq9V6liVoewmARMg+go8dKfImol7N1qC2diBge1oJ28/gppEv+rjOeMMi
48lxnAbhi7qXZ0Aba1GIfrTGURFSLLHBqF6OK3UsVhh5irpR1ex9F9aHCuQ6
+K4TiRtfTu5SPzDUg7CIprd0JyoyNa9Qy0dwoxXrhlikOoVBhuIRclERqKBu
bo/GE1nccgmQtgel+QLkuNQQnJiq6xS6SqcV+WylRjaKZKbPSTIhHxitMWl9
OfiFsCHsXKxSynv9o+jc4kZ1kxzNPMarphvfqCH5bSfXkepTA0qmwM7Cv6mr
PsIFewRI2wNuhTNbobW/nM/2tSM9ZBnUbkycB29HV1YHpPmFmHbvj+/zfapo
XSAR9FNd2hPVlORYG/dZd9I4Zv02nybyPbLzzx6KG3rmZ9lgMAIgtufZA/W4
kSW380uRSb3cimgpky31W4uOK0xL3jKdGF4ibgmrBVezmm2elIRI+TOQeji8
KysccPl0fUtN3/dDsXz9z4RwO/T7eUujN1dzzCj7nknXI19S6K7pWhL4Kcyd
m9xfahKJRpZYdS/MHWBTZidJ6zrN9N1VCwwZuTAh/ZudyCjBClkCshVtxC6f
KFryLhZQl2CvWxDljnFn4IZ31C8Y2/lN9BD1zJgpi9FaOOPgKsLkONWYSkyj
8tGi+mvrIoGOFPBHhRfBo43BVb9xKc6Eazv7+20zaNtVgFVI/2cUNXBHjLAG
cPSlOeNtLJ2rwPUv7fDzE/BkimgyhfHryzeBSBBOAfvaW95B1VMNAT9wmFOK
MyWBk+ywgRFnPYSpj52kPTg7EDX2dijclLO1Usmm4kzaTnjW7OYmr858NrN5
AMJ2e3DEOvqT9AmbgOktaHiO/MeZzCSgC/7NyryrQCvWGfj1zb0U5xkpMAI2
uJSZFfMmfr+8aA4n/R/afLz/d4yOMuQRc7sPWiy+vC3QzZVG1GcW5NZUGNU1
eaihXhFYWe3dcwBD6MUXOtuMmT7pVBb8rKc3vuAV9D8M7Wc5XBRoxZBoAL0z
o8Lsj2x5bt/bRG6RNdifpIrBjcWuXPfI5+pmQNTmqPU9dYBVXxNP4ZDFdlXu
RWJud635mNgVVxAa3Wjc3mniDercT0yZ9OUjcDZmKmM0WE3jaLdLeaK3YTdN
N/lIyY+Xt3N1W+6Q2sX98evXaq3cs882gQZGyn+a6A/JIvg5d0ZoQ7DJUeEZ
j6fWVQrenNyZa/Q+oiuEPNOCjcKrYvS7PurxCz2vxqUCgnILzeyrFpuySoh/
lhFJaBb+yegpiBLM3gmGxTGN6coO6luzRbLxCO4D3I3PvVjx7VkZioVidQ3y
K6oY3nO/CcaM2GlGcGm9y7Ehv3iJ/lFKgervx0bUcA4Tbmi+v43a3o8m68b4
5qUqoOWuFQeDSbcpn47nN+29jSrLisgSalc0hk5hO5tIWJXGSXnW3nOU9qUN
inZ6+Yw8QXhSS3dodfwlCXfwMrlGkXMCVbKqUMug+GmU7HdrPh6cnKSOKEZl
2mbKGb3kEQ6rfM7Cs57hYxSe339Awx7u7JL+gezuBbmvmdT7Sm/Itz9IvGYB
Y2Z1mSbNmPasG2pImiXDaBz0Vtu6Cqe0MhH0dArBYIjzzjX4cxrif1kxBBvm
2YPDPvBK9q7/TJjStZ2SkxDP4XyGM6Ky4FDOzqE19djuYFqi6erZ3YLVTiVg
02j2+Uq+EI6E3cxeRjxdVyrkgr3gzxN3B8MidCzW6PeNtBW3VNeMyybFJzAh
Gyjojq1ejS3C61mv4YbNFYC4zyJ3EFbWToVqrxMk5z4DhTMSyozwcyhAEStj
gLGNkOEX9A8p/yXf3CHfOPK7qXdEAJM0OaZZglR6/NT2fe+OxvUFDgnZX4Ro
jB5ytL/rEV+X+HJOOgWRgKT2TqZ/EyquaqXaBV7uACEgQvFxlMFdOPIsWl0y
qKkiHsYyjnbJj3HbLtlB6mcMWm6pdG4J3MURmQUj8HLp/5FbIwRnMtRMZ58C
i1lbapMDVfbRXUjHmjP4WZdaKMv9vWx/VsBLw8oqIjsbiVB7sCLtOUrcN7kh
lizrR5joUMo45rCjHlY/qd8CZEhvAJjo4lqV4mtBUEN3IaFYfaQhlFeoLE1M
AjHOiTOlYS57DyYN4h7EbSZ/b8KdSEk7qXX6Y04+U5WJu46ueWzkRDDxdQy0
mpD1SbI72uAfeOkJYS91eEjpBroSTJT7jzO3Yk2BobfvW3tBztoXABy5LoUG
FHc8kj/L4IQNt5Vb6MABhlL88H1ct63jOg1CyhBNRIRSCDyS1NmUqYmlYofs
lNlAVI7wxXBiEcvKgluPmeceuDYnM69vOBBRpArK66ak3Wo3z8kbWdcg9eE4
2e+W5LC+1b8aXv42YvC7bIW2oa5H2RqEF5c23yU1pcZ4U7Y+2hkoyJfnieJN
EeTYVgGPGo1v+7f1/SdZlzL3uou8aHQM8X6G5N/eMKrXg476vy4UvuiJxdx/
q8xMZTwewBUZTtxkMQPqSWY14Q/CgU1CW5VJk85H7Tvzx50W+1mLuyImfXbd
L2mPfqc6/gJkj14IZZ1rAGOhw/6rtMU2413cM+TWvJTL0SPtHgc9Mxq4RZpD
ogfjLxat1Y92boI/A9C/pOZvXdBHsG+6DSzUO+i6w3VzC537YVCSx4LORxEZ
d3lnn+D+pY2GdVRXZxDbxJENKLgIYokIIxderWrtxpLL+gFQYp/L8hYIO7OR
tJg3r28MtTjYL8Ein697geh/+3cECN5K8G2U0iRKRnVrdNUEDoN5zvZNzq4w
Tm2s5JJ12+yZHoRR1KY0c46VYMkwxosmPvqa1TwJv1fKaly3t/nb1L7bGVHP
IwvdsymWkpsSnlSuSlEbFJabHBjDH+yLEBLW5UZVnN34IiiHRm6Q+AzdflUK
bnZ0pQWbSJ8Xqq796kN+GjTleMaWMU90Ty/LeTn/aFzP7aF+eo5dOELHG2wv
8zOIMV4lTzBM5446YK78+gS4ZKDfsFnj9PinD+7XVj9dHa18Fxu1UqgTLBC4
5bNpZl/SSloZ6Hf5urVywhEOYFO4HahO9XUBAgm2vrRHu7yn8xB3f217WkMM
n0Tc3CA1PMnyawrxfYlrZtNYLmXsg75s2/KMSgiwpQIwo2enzsycWBwW25dH
CG76fpgOqISnoEs2m77sLYSyuHzMXPDjH2zFtCR4AWDApIF5ecPv5uehsjy6
0qCZCXV2YrcI3V2ywAj1qg6G1Jlfaxw9eJZXYrVDhfSAvMVwKC3QHCxQdwu7
i54taLEEPiXunniuIy7Q1kDpt382rbqmY586PpW8Zi2t3zxVTUsh+t6jtGCh
gT0IzdTH1u5F1W588sx3d218a412YP0xjBd5qFUTfOkqmuewn0YX0vgFOFWq
IKsJzugdatAR/psNyTcfDeFfM9s6f/3yZNl5AzN4qBYwJLjMn+cCXo6pTD5u
GuqK8Pz5YFOrT1jsrNc/E2wSoShOFkwKMw65b+VW5EEGSXjz5b9Oo/V6WhgO
sN124rlMSuMD6cVocGHRJMFQMPrnvubPNju1/eagya/jhfPHQuHDMtZQjlVZ
8K0PfZm5HMfeYdrr4ykAixRzGyvd/lEirQRmDu2aSGOGPDTmv3qzdKS0h9kn
jJ7A4hS32+jufBd0QHWymKXiTf/XOcFoWRDbDYhbnn15N/qM0oDkJxhkNCzu
SRH7Kc7IM5OfvkRuTcCQahoxYKgZ3fLJXhicQJZsHT+CScpKqMq18jYTvNSB
Mjtx618U+6R/RQWgMG5Fye2KtIkeRnHjbsP4qNVO6dQnRHBgrZ1LdX5Kc7lN
Ql8DjU4eZher0Mdb+JN3Fc+NCoF1oKj24ekkY3YbJCQA0U2iYGpJumUJQnlg
y29KAzldmkUa2A/EUcytr6kkxzg6MSHOxpvZxDKUev/W6mtACrIB/a118M38
7lEpfJQ3BxzgAQuXF0FY8sYArQeqykym0DZrBg9FazOH4aM0+8ojLUi/kQ3k
w47nFviIcGk57DpAjlUz4jVcKtilarGtCriClgEkljeymITXe8UiIIazl9hh
CDcmJJZW6ZEZeZhIMnhq6VfqqwqVogUSZnPDX6IhkDNKHKJvE2E+6rzP4+br
3l2Q4L5CACYk2PfHHsnK5/SRsT4s3eWSyf/Amh8aBbwfFONjj0NibIQ0o2oT
WpDwm8/Gl2pEPcGArT4RPco2mJzQZOG0t7pZsM97d1IaDfg/BZYHGhTKdwld
9spaL/3v1rVj5hWQQ9rwSglcFKr1Y0IrP8RL3lsrrc4rdN++PI2pOaYRe81M
0RXHr17dyHsyBhH5frIu6edYCdicHwm7UpJeMQsJe62kOy8C3kzWLbV+qFRp
N5zJDhOIRS+/SDZVFB97ZvqxG2i2gNATbPHso9DiBCMwFOOktDxsbdkHpPLc
l6QgYgHrz7GlqvNxwuz8+tRtHzEciM91kHj9OuYn3IfAeltoa6xTkPQXqw9k
kKVLWyXAUapa2cuXq+liV7xcnBs8XAvu+a1Dh4vLOfJ58trBFi6yzPhxd7CG
/8eMwqJzUGqoYlrLj/uDYV2bMW45K3UQ1pItCYpxNfx9yasrX7QDHIctpAxb
HEJ3QioC67u73CfVGl1vWMmxjuw2WpDkWBxKKCtBrVqovZTNWZfqxXlwUTjZ
fMGBRbj0w0f5IMWEVveMG2ocVKasoOOk1gU6yODAJKO2FuEYzTcPB16Cr7gG
oe0FLp9bdCKhURBH0p96vC9aFA+6khpKmj7jmQ+ot8ExLhCjo5SGE7KQ2xjB
MLicbAxXxqCIHsSzLgEkLbYD7lKumk301lcBRqb9jNNBlJ4ct4c7ZLNEKrrV
aU6lGYooaXRG0b78CAIVcs00oU50XAK6OELdthQ6atX42nMzKsFjlXPoZG6S
BE2yY1DNOkaBr0d2f4EepCwOkGKjMR8Avs7IOOdtDAa6ayiGeaqKXaJqU13e
2NNDFyY7WVoOR/yPM+jRpNN89uS1/Ac0PZoAYjWXOjpY1u/+nbXCaiUbyKx2
X7x/aOFFX130zLQLnn19VqRneGrvOgKB0bq/KJoY0RXLkiA0FHwv+8KU+ZMJ
pIYaI8rNAg2bSnyGDXo9OxGY2T1dPR/DauhlN/VLu69fml+9Fxn8oTC7wWtN
zgDLS7UAZYJycEOFR5i8YwTb04Lc05Xo2PEtxJkyNblufqlBr+xltUtCDE1a
DSsqk/124hgWIb6LabJUnPfGawapmPY9OhSI8y6K7qPCv6w9cnC4PwFDZD3d
Ik2h/GlWy9hHoyf68FKRs46gF92+E07P9oETlGTtPoIPCeCHE2TkKCFr54PB
MCzCMrVL/y5emUvziu8csMvCoGsisNbGcNRuQTQKjf3BlfIUTnt9Gs03dQvD
uw1VuC7aKD/tX1QYxaU0U8UWuvj1qNdPMBYoK1+9eCF75SDSbpmhMPkwkCr1
jtiPoGwkeTGCoomhHF1nOv4BiNacqZ2J4A4oKZ8YT+e93e2z3Kh/oHflZbik
6PpG/E/1bmkeNvlPPkEorEfFnk+W6rTq9FeU7l8gxQTKq9jCXm0H0j+glTOn
cSdmFJNPyFLz96A3zn4sHjb8M8hmo2PC8Bznjjft2G1XW/5Vs7ddTm3wVLZ0
odxhcN15xcq2WT06dCTozI3RCa2sclAHL854Xrguzmv+VFUx1i4Z1+AE5few
dshbkmCVeEHJ+EL0BV5wEFzz+CrxwORuqx0WydjmjzVjpa5RohXUm9z3yDhc
EhIY+D3irAxaOELbnncq+MXFM+5LGa2RRCEXvDIY0JaU82S0izaOoiptTtAz
b2qIXoE2BAKd3DCDN5AppFyYPCwkiYm+gAYaR4RG5jy33HhRM6muDbMEH2Y4
MSLKOeZVVeYYke2F3auv7DMTSj2qf1ONeILjCjaW4eCYWiIO2cyXc818YrDK
HXaNJactHwMJrvk3m4d6tReYVLzlaJXEmHGuxgmrha8LoGokXk9nua1GdVO1
yyYA8mq8XJVOGFwa1pV4GoYtsGN+UqHM9WH72M/p+3UizZ4zaZLvCyW5u5em
FV6hP5XYMk7dEwuQB1qTpXcDxMrVM/b+tsaPbfiCLLHuWY4H6TnAFdnyzpU7
qfhEvDIIh7Ma4JerVR824wbCuoRGHJC+lwf5VTWgFDh4nuQKPxbuUtmKd55c
LkDHR+3dRgA2WCG3NEKcDSi77DSvh2+ai0N7jw0dTCYD3p/8e95HbCw/5pSP
NFgc9ayBVx3MZkvV2ZmhViKoJwmZnHgPd00tFNW+XEj7K2ql9FnGYtSqacUr
LTyB5KcuAmB/IzyEjGV0oTZVaSQxOYkBDoBwSP/0gWJgkUYw28htSEV9iugo
koAhI2b1YQEPUPddwdHbWzH1FW9dxokpA0T8mehNNG7OImJ/ZPcK4FFeN+lk
cSzAw+spSTYCqMk4mGm4962NYd14bB0doZjjY4Z3NCSzmScvYwet8KJwx91W
GyxMY0DXoe+jPvcH9TSme1rrSXeaXqexqDp8ss0zACIGIuxEMZNvvt4yPvbM
3yXbMILTBM8iSsa990V+pLS3KeHfdWRFAXoHLcRX15+Vx2DhOUC/1QJk0SWl
l/7ouYe7BdXIrmHNzjaKFVcRsqlQUOCw1+oBX97epGMrWJB1bDDg9wFNRtcx
Ca7Wu+FX/UaDWHfeNFg7JIskqd+gTLqMhzCYUUwfTDTqLZ08c/DoN00ml9AJ
34et/jT3hKUrbYNznT3l17EoMWD6I3tJ3UzhgVRTwaeN/Au3dKRl1o0t0wzd
zoKrxvbKXCan6eGegU/+pGtyGkgjWW55PlDtfZJpJLkUnMQyRJ+RZi9qZwaW
WyZ0ZI/Uo6mTHMYkPqSSMLuo1+3N5YO/phG+7JPNRqoK4oglRhv+dYdFf6qT
TDbZWxd5W9whsRY4YPWEpqF4NYQHCsIhy6H2ASfK9TLzj6MqXTGi8zDHcprr
n+zFDIcjLm2Hik4maA+pnJIFbtnjCNlC7ZMfid0/YAxSgUfA6J+yidyl63MA
oLk2qxVb29g07c17oIMIBxy9KlYt0OcxwcjsQt8keEnNABeXPdDDZQKByxEt
Loccj/FtO+IW9KVoieWb/QtGAqjm0GsbifJDPhg/RXY9QXuaMtj0AWQ+1rv8
AyKARcEAvX2UCkIM49uzZQsiKhiV8GS7HxCRkcrMgc/SRGbdL8Roz73heuIo
5cndRVp2Gdvrwrn4sr5vAuj9TujAPdrY9+/09dYzhDHZ69Z2Yq0Z330c5zTT
eA/UCNksfJTzGccwn0NPGVYiKDp96zI3UMViG3Cl4FIBNhqbqvjhjkfKDYi9
RRK/OCRVFaH84Nfexoi1WqJFTDR7k+CVa1n4ztCIzwJ54FgNZvIYIkv6mAL6
2VkAaDwo63lenu/wUi5CI74XUQq2cr6iAcKOsKNycGM4mm+Vu9a9OZwH7J8T
KYQNz7ZNAG4c7NuxgCI7IrzXdqt99MAQZ+fFpRDEUGnUjD+uvb1NLq62qWoh
K3nTWbmBEkOJkp/d0cUPc6wBo4bCNYCXNvXnzifA9ywv2zyd38AqoMGKVzBq
3e//nZ+/7rRjQbLQWe1QqBpZDbkZ3wXv7HHjJCaxdhiLAScFeh274D+Jc+bj
m6A/UewDGb92ywo4DHPrhKL4ICqFNY1DjX/oS2KgASx1na2prlRyydOPrUPg
hZ2Z13T1OxGPkaJKbR2ql3lXqGWfQpN8mqHCg3csiLGmXpBh/Sr/6CAxNw1h
spMtsgPjIoQ3mOQLIos590dmEJ7+BOWVM+giR9sUpOgULPDa+X7pPAmPvH68
BpLG+oArEAGHu3X2jnBwBHc6LijWZ3DB8zOtxOhEJa+2BmRlv2o4hhv6ges2
lErIQq3b2ipGdQFz+mAwLfOHpZKnT5siK4cM6djUzYV3otQzqx3aOamLZLEK
Rb8ogpeKZwtHesjh4NpkstDavS+X9UfQsaGP/UeS1fuKaoxzavmGztQG3Zwc
2+IjNzT7T+7H/7QLMnn6GMNw+ePVFVj2O7oiiBk/zbV4uOeeV86cz0ZuV0cL
NcJNGgHfOKqMPssUZ8cXjC4u/xfwpzeaROn1Do98z5L7ooecZ9EU5ZDYpUEF
K1uGJkTgVFgMd4iM7a2OjGJwwhhuroOpVpnXdavfo/1RwxAmvcQGrfmyoZ5R
ObgzHgIitivL3MDbdVGSqsan4iDS9dSL1jqZtGVzIAfuxlMBmW/WZY2WsTii
YegRE87wLvXX4CwgHdDCNz2qLDgljWBElXOP4IE+FKipRDyXb5HDvlL+9W5y
0MW2/a1UYJaYyTtUxvaecHhiBOkT/Ux2bBz2glqNy4p1Pu3UZvtIAAtRFud8
pBpVyWQQcJSsR6mt+EdW3DDtJVuRt5zo3tOBt8g0VToZItrSNNfj44rKJVXo
O7zwQgxAqAkWBmLfOmeM3MS0Af5k8cYVcEIHuZQWjICTxdlB9vwCZskpsMvX
KpX7GkLHoE/QJZWNeUI/MipJ87SaxKwN4y/cwL5KGFi/1gULsN1chskTfOxd
GtYZKRK2zBWd9cj285HRncHb6poWeyj7lBfcuZCtdhGSkbqpsoY/5Xa6gMAp
Qw66Q869IZRAdEYHjbTfkmmIQZhQvb9j4OVCqCL2JyfZk1yv8X1Mtm6gLMkn
g9gg4xqLhb36B7B64MNM1sYSyRuoo7WmZcnyhkZ6kelj4LqBZ/gj5/KgPRxV
Da9PRPjvb3h9ecXGwvq8HEsI1Nd57lIbNfise+r/Sljelt65PLlg34GCk8LY
qtQ7I3km4EU6Jh+20QuscG26UuUoxjiVY2CzWqF3rBjbPTzFulEDFHi9ICXg
28WN4wwUKr3azOKUiTb49NM5F8ncLMsaODcpyf1P5NcbzPzCoT5y43Xyl6VU
+M2z2KI/K94+j912lvkNrmBFyuPM3QDsq6cyBSBuPP+QA2t1EXwpDxmKwILK
JoYzrmRsOYzcV6c6ILo5LZmcskk8uI7txl+mURSaF0MRr0dvMUvKtkoL3ymi
17UlyK168qDZGP3q+cJGiE1FDrhaUJrAHBrz10bVUGPJ68pNXXxUZ9GkmzTc
7bU2NW+RVQ10wF67FX5L7gDKxbV4NaTmKFuNOV8FYYSFfPcqeoXStgGZHHcT
NjYV4/pTjZwJtopkV6b9KLj4zYTNqgyWyRAPNXjPTSuXt23Bef5Qqrr43ikf
BDUt0m+qIsF+Dz0gvCkrELSNQQQXnfF2Z1SaiNAi8IjCHzTVtBi3uJXgKbP+
V4X4Rgqkoh96+FRGflYs97PrNPeibO9JArrRwjcRBsmwJPPAmXZrCanX8bUa
lriE2BVdB+BiMHYWcNMaXhDbJlzTXmmvFn9PSF5sUuxjMS/R0I+MWbDQnGPv
UL8rpz0HeEA3bSHMc7uJNnVcVfInv8XVSLHKtEzpxLZo6v9452C5ecCBdhdt
qoG55a1JmGzqAgavzAsMXAPEhzGP/p6YGrQOdnFwpjMDubf/d6gby6T9dm0I
Y09C9JrJz3M73y6BIyoBHUS3SzoTxCGcCHQXv3MDPWbWOrd2yJabDDtMd9H/
SI4Uko6JZvBT5lsblMaNyiJtwzDU/sSbe9+uXXOFtZCjKe7+5qhpQJp+AhdO
Lk3XMezQftGe6esEswfYHCWK1B9UK68gZal7AdYyMxfLKFXX8joSaoeg3nkF
bfYuPb0JBexlZ4jlOz0Hre7sV4sQS+MnI23j9ZlvKpyYzqbkwHzIyoBI8DEC
Jvvpi8clWBznbQbjC6/5p1IqIOHzoioSr4qZJmoeRMppNVJvSfItG8uaNBfP
sVvJJjdkIAArud1/mFEO9SrZ2aSh1NRstmThdtgJgMIxztdzzvh0kBLSkkIR
/ph/eKMH3NOyjBETQgTDqUwToGtDF2tdLym9/PmgNb8dGlSnYDy+An+az/pd
kyD96gLl3Fuck/eGTICMckGjU6YipW6rUpKHHwBARju3JJtE8LZoKyxRqYle
7uDIkTS1bzAnCvquDpgOXQ6Eda15jPVzozy8CqKnBNFAIcsXVeaFNHze2GqC
snc13xfUTc+GaxrxaJWRh30c1gpyKxq8wrd0kSRX9HsQ8jUU6WHbeXsHVdpA
z1M34aR5bDEFefzZ4Zj3nzcG9UlY36dd4aUuJ9PNdtaVXnVMI8t4abO+qqh2
r/VuIzfZH5Ec6VqLMRQK0dZF08wcQc/IyFZNT9YH4j2AgazDpmuJFnRopUCA
JhmAVaxGRmzj+xyXh7PisxN4odgq3hblWSSvOgXZstXvlQAAhHYNpigjEFX5
Ea08Bp7iPYXJEQQb7in/37w2rVSLDGzbyqVl3tpGM897HuaXudkNH4Ha4LpB
lMBpDWSqIgaLL61hfUCTo191UVE/PkhQdSZ6a7OG5jd5vuPhIlHT/9Ou2fq6
yWfrCjJnx6f34Uulm0Tn9W4FwV71jI9iKNFIJA3nUUsc8YSAB/GIW6+ytqFd
PfrU3WeEeumFZ6DzMOgwabQ9WCRVXDGirtagCkofKAkk2lhqAQJnWNXdGw6N
RdmYtMOJbmzwyIy2f725OeqkfODV7vQAZJFA6KSP1z4wmPr0wjVLtOrpImp9
k0aNivLJcD22kwYDHi4h5oSXahY/Ytu0Av9DHNEy3tTtuxJ/95SXIQF+Poso
lltwSnMTL5fSilIrduHwqzB8wxvbuMuR8Gvh68JRNy4x30piGZoXJRo76ofy
7mQ9f8ulAaw4P44/AxUWymgFcRXOGwbTuyZ7/y/PSIDYDd4J7aHNoariLpwI
0Rcj/YUjYCKTbW/BsAynpzLUd6P2JeX6LdOhmdo8Sypt6yR3Zi3GBwIF9eKU
SWL95OINmct5HyVIqKm4kdoKQ92cdWFWnmN1wwNUZa8FtsE4IDYUJyVFzINj
zPDr2U69AV2pCwOFHmyJaF9ZjaCASO1zf/CSL1/OC62jkPquH1S2LCkEgr61
02M2gDf7Xawb/Ih6haNwo7EjYOpaLayGS2Xs/umZq7PJfK8LaX98oyW5lDNW
5hrFijR4izpBodN6PkBnlfPWqK3CGhkUjhASJFgHob18IsPYDZgfQg9eRE5x
Knu3A7zuJl/Pg9joQvITcxpix5rw1o+S9JTN7x2OLDwoTd5EhTUE1cEeuhta
N6XTxqLzkw32BCS84iIkkCQnn72vfX8Y5HMVVeNgNCTtGZNC52g0QD9Tefug
GrSleZxhn/pIS/F24DXp2qFfQHkTcuGJMCRJVNqLR0h6CZmwCrdlffmHSn3J
U4gVfVfutsh51PFalBbiFV8GgcNxETUB3/nWF+9Z4b7crdQXAbKOhTatV49e
SlC8tSJLyRswJvch/slAwJngJX1YIbjD+l0f8PcBONnm11e02orUnS7GdtUv
2jOi21eP5l6ToFWN53GjlznfXezMcrH9kGBEVkZjdqmfOqSWkcojFiv4V/7p
tjPDKoeRgf5/FkdyUXUjOSpT0x9M3INmOHm/V2YDgZ9tRZGs9azrUp0vwKzG
XRjbzqKwnsc6yvcE8g8LVjheBsAHPBx/YW4OXifwtzEzLDlfrYuPJP2IoAsT
jIeGk+i/lA6rifjLL1HyKNtxtDQI4TLwV6I9LJQpkm1E9HSpZLO+0zK7z00L
mUIYlIYk8S0LjUU4dQ7SvqF2ZE3XIWABKxQR6q3zrnRIQEPKlG7TYI9KP2ar
gKbBliZP1xGh1vI0qJrcNs/4LWmzw7sSbUC/vN31L2GSXOr05PWVHu/f9q4d
App9Es1QQxcCtlaO0IUVc7BtuuheJl+jgBA2FO1d9WXyGoDFKyXlhdyd9bsI
O+b+Ler/tdSmhs0wRkaXHOjxA4Sw9g3Zu5CDtbLKRQ2xPre0Zx3nPEHujIGW
d9AfYRg8SffEQsLD8bcqU0zWf8cw7Hn/sjfehFUqjXcaXNFfrd0InSC+6BkG
S7n6nvxRQw0eP0ycMrcAAfxqSwYn+O/0IeZgBfE/SsVkGQqdAg/h5L0sw4ML
xUpGGS2gb33bbT2UlkTUQhelu0/91J7LhUosl4wiRquX6ferfp0kU0QYiZye
ayAFdwrCfXvXSz6JNCUFYhawGd21BccvGSfu/4LhycK5EMfDCxvJJnIVzbsw
btaZG4blV2EEopaXhdB64apcaUH5/6IuQVMOLbqiJ8bvYhY1ShMIsVFT0cA9
m1+he+ddrRTOvwWK5R8oYcYKfwIvAcANtFeR90Y1HDCog/5Kui9yQgUsvsTn
dGC3Au52irPmykZvUx6R1cS0CZm/XS3JMJT6SprCiOFboThMNBOXDBEC8bcp
gSPrZEpWgWsHBl2lMFrUOzLEQNgKvacPB80bTVu4AUVUcBAm/UyhaejVQue7
inD0UGqJihmYy4n88hhE6k0FoHdfDCeEcSj8cSpbeUGBBKXXES+U/LudxcCK
QTk1mq3hZZnh/FAl0wPJ1+wcAjFi0lpMvuvyGxwaD8NOA7ewExys0Sm/TDx7
S0yu3AsM5eLEgalbTOix8j3HYSw3zjnTqyizXHB3An2OBcqIsVNZ4UCfMhFi
J31AWEY4pLsbngiH1ZZxTP5bCGQCDZxtRapMFNvk7ct1xwiGRLdxWn//Fioj
n7RrhAQpftDlXcc0cV3H7QufufEO7JCJiRKQa68B7HBj2wEWRAzVxkzrtuUF
vZB/eFZWdNCBD73LMzsuXjYdSdluzKBJdqu2HoNYvjidjWrzGX/Iob6lpbpr
guYwRdAkOMxZDnaSQNl/GdFuw9LqChTIQuFBL1iZGKV14w8lWQe4hXxYtr8Z
3a0/spzlb2UeV/NkPzX2WGucFHPGKIvIqrBw7ody1MX5c3h2bgVTwnyUpHvR
1ciCWLCbUtwZjzOp5UZKqjcr0QEAJZ+qiHxe52AAkKcxYiY9fnnLW6vEIFiU
/Welgt9kinku5XNhNdw5yqsVmuRJHrSJUzp3Xg0G4arz75LIjZ7ons2epXy0
TMKhA5Rf41UUqGRksnlQ+pN/7loO+jgslYy8F3mypMjylU1R5Pdg31GIIWuk
WrLKdAMqx32jlXV7gqKo+B+Bo1KbWVblOiKp0D/oPNow+/mdbc55rnujonE/
vgvxYTTdWa0jipmRdCeDY1WFnKXGvbr85BoDcSfFUmEgeDHPOejU/IdFyvwp
KAoT8engwYaM8NW3w/JMyyGF/SPZirflKvTiE0om+3QQQ1noeHKAcQ+y+Trn
PHgyOFGWL9ixA1ThIZmf7ciG6Gl8lBrAN981hmccf6oby5wvGmc9qIfwwebb
1zoD0crF++pOsYmeNAo4oCTJKu533N61hLiO1wUEs5e30RjgEL+sB0Zs1iMh
IzuqSqbbkNherFfXteeq3tvWYRh5C27jN8pmZqAEhlYZWVj9VmDKt25X28sX
NqXRm9EXCKNMBuWZfI1s9B6ZZQmIlkIqX7lh/safHFUhTQ6hYG8jTOZTtmA9
KS3k2KznkFgDs7Myvs3iLGiCVQBl81sIPC/OTCpo19tAmzBZz30YZC67WZ8C
+oyqRz5Y6GUWXGCtwBCww3gTeRmKAnwCyLRYfem1j3zG5Lwgy7g7sEFNNV5/
4g/hWjG/tzTu8uwkFdJ7Qr/yw7foCr9EMyi51yLixczgXiKwgV3r9irEVIfK
iBB5xpWbxwvigEqm79prOKmK48RGvd6tykcQ8eGKzbtMCBWXlDRdttkei79Y
wPojYqp65a4kZxPD0alaTpVRfTTzfBnf+xHLirUivUB/9ugUWiPXVOQWWbBu
X/2cYGHlTVkf5gy+Co9uzKBoB3HzhHmDhzEYh2ql4MwqhlgOfDWaRwt0xgO9
tsjP7r0BnTTXu/1Th5S6mLwkQHgBwk4Rh2EdZjvbTn2TUIT1u5eWeGijeWXt
wFqZASbGnbzzB9nE4DUbWCRJrkaPZ38szg+FeuNfxdBFNzpUhMpd2tADXj+7
RGlMoMcxCklEwCMpNCcgsB2/ki55yGr1IjHgzgzCay9Xb3K+ptXOc0qu1C4D
B1YZ+Dny7WOdc51xmXixg0znZ9hGXXGv/AMYs7WX4jCuPvpcdZINqOqtmhlb
rtW2iRzwI/vxXuY4RxcjeIV9mOlgYuDU6bLeM3HrFRY2J8zEXaS2fL8whRLS
ePPdsMdvCvIJNN5lQdFonEQbZj1bLnfGFh9c9AoFa+1m7iwPs7GNUhMe2zLg
bj+ZDDdnQYBlBgBqBBUmuqg93PFxA+l+7+hwFiBXW4HkmaaOzqJDSVIyLq6G
azQD0iPM74GzC2+TSA+xN1C2MoXeegF8XabjAeaTphFXyCFVGBgPnyexqIZj
fGKAH8gJjWhtP0g/UcphLdFJPD+/A6HO6JuRvQG206InpeXQHNLTk9hSa+Gc
B/LzzwllZ1P5/XaDoScBF32KtvUm6K/2VfcOVG2mcz6Epfa1/mZIlNmJjCpD
+wnp8WcVQKlWiFq/OR0J4uZRP6jbaXsyeHTTKoe5F7FO2iHySb7NskWWzW1B
8JCQeWBqreGPFtE+OqBD2ZcPuoOH8dZ5sFouzvrPpUg9cP4du8dsXsK4y0GZ
xFRRiVJgY+U9dScYKdg0sLreiR0NoAnacHWFetXz2oFc6PzBZ9szQvjEmXde
wxTZB3QbRKGEGDoPhaa+72zKkX3oD7S1rsQcSjzX0iRPkgMa6wzu1Lo6N4sf
epZZEFEy2wMtSy9bQF/KCC6ir9NV8t1M6dgQUrvxdYp7WlLM4sSA2MPJO+W/
os85FgFzDABm3zIM7OK09DJZfrkIEXOZBOkc4uxI5Q1KkUCk4RuPta60sxU/
HO1v5RcIhnTkzqnQZq/X2Goc49d/Z0zcZ3ELi0F+lmYIN6FHRNiVBqgAyz3D
suCwmktXqzApGXFoOsG2ObvXpa/1dNeOzLQPEiPGJ7szl2NHdVKntx3kPHTe
81nwnLj+vt8IqniE6YQWmpzyHLsztnijKrDhl22rfc64CBMWALlscbP9YLJc
TbQYwNpNgQ3N71xkX+PbQGABo1gvdvbMe1G5O+bssDwQKxPf0RoIfizRHzGS
9KA0LElwhpRW5zEZBCnlMMRNavwtYOYP3oT786KTyh+AoTIJNp4vYrkHpOOD
IWoe3wXlwmmhONGGoy3dp8ZeHfNOXfZnpuMqraLpv6EifY1yy2l12QS4jiv/
2Uv64GD3ngrVUHTZzmr789W04ACUr34blZ5B9cdHz0H7aI5obkO6iOiR8iPd
OwngNXlvR02dnT3RrhK6PDEx7X7JnnIPF9JywfY58qwbrhEaSmxp9Gy90hLx
GaP2wML9U6uEtq+m5OJsLg6CFG2zWVbFQA9QxY1NRGQrPe8CgsOxrUqgJuvH
WJ4mcfc6z30K9zaDcC0Nfa2SFzQENmgD2KxkL3wk7dCDx7+wt1vnM1CCknSG
JE8hn8XmXFzc/tkKm7Hl9OgBeXNOBbHnUGlF0miKfszdjT4aE8KShRh00wA/
8Hi8uVzwsOrtykZ7Q7JxqPvcnj8kZjc8YjjYhBCW6wByoa2KxaFhMvq6DlSJ
R+8UR2XoJBHkxVorbaEOdAarAwrCJvSpuu0oXcaWSFCviIzA41JWOZcRhecG
pAngEuLoe2rEH4LEyddCGQe0j2P6yTL4I9B0/omHL7dpc4cnmMtDHW6dzAO+
zlgNHPdG/yHwAo+Ba1mjMw418Sbw1J9+TAdYvx1CwNfgls3iRzrQJ3j0tsI0
Z3k70pVpho8XmAAHfCrHLcV/r96OFWEV+noao+nuzc4vfZ3jvIbj+2arx45u
17QwizLPpPntmuVtji9b/khXmwrcRD4jUQ7AlFf8UP9lS9tWHQQccOjeljqo
soEbIJO6Dm2CHNa/gt9R7ZZnJ2uZ4wH9T5FKc3R1T+anxWs1ai6/Onz7iA8Z
s5Nst17LHe0Bn2IbUI3wCopOG4Z/vlmfBAl6nLbhkpw0iEpW7BcQ5HfuvNz+
G5y7+PetGd3VMQv4oX6bYHHw24PKqtxC/ecyzD3vqnZFGh7jmsL0gwuQBZpl
JVPKSdH77CUMlDorvkvNRUp1KGNBurnzxTCepYcGQiIqMftrxQ7kK9wfK2+e
eojHBSFFgomu5AZfXiWckcOkzaP4O5UzAb04+sSfDj4yjd3r+2ccxRao2DrT
AbZD8QlmpVT/CLy8sQaEBdx42uvgwMiK6fZIbB/kh10H6WP+kUhxJHBxRMF3
Lrp0qw6QsXulpL0RAEq12xYJDnldlE2cf6huL0LKFV9+UlJ0NoNizDoQgxMb
V8k7GcXlwPL4yrG5zicJ110ciiBn/loPaV8N7JXcIivyKIlPgTKMj0P7w0mD
1aoLlm5E43w7d1nxC/8suaeoKpLzVHeysd3CduwqhNl4KDL4LePNDQ1TphA1
HikalSuxmf89Bxt/zEE52fR+VtY8JG8/euACb5k0OaOxbBCs6Kmg9A5TYr/n
LwYhDnBImL+15cr1DQSs+F04MoosaRVBz3aCicLGfbc9jkcxU+m9i3YRTwLW
PtfOdQ8Fo3nYz97kUniJBuoi7om5J29RNUMWbETyZHf0kfU+csZvx4izTcF+
ZPRFgUq32L1p4HzkjDteTHqSvg0k+RYqEgYEIDFOCBEmu0WBlccQW0l0ng/g
D0wqNVLnJDy7NavNyPuW1bnJLjC0rlvLORB++CZlhTCaLQwD1/HzoEHSGGUr
BK0zGwXpKqedCRcbXnQTvgcm4UssnU4J5bmbCljkAzwexJiGsxy1ja75uBKu
sdHX0HV61hT8rMIB+OzUDjhlFPv1wp1FaBvMYcAI286lx4/EnmCD0nDPqggP
CrSIO8D4IQT6xs8dB9BjEbWQfhogKvV+e0EraKvxYiNNfUsBiO/qGEGM01J0
Hr69pJDcVlQdVNKJxf3kUiMmqgmrzKBcHunDaj/XL6YnX0yWOYJ4BdtD8cxi
Y9nhQDf0Xe/82W73CgAcfGKqSIkfJEl5blQWx7S4I/1c2qxgF7i7XMGQ+TVg
NhRH6IeVTtl9FrXauXE85EOOxG+hMhtkPLM6inuoQGmLAukYhjWuIJuhNWAZ
U4VOWTcWeSCRMrBm7pFR9Et1uZ8FTQ4TVaSKUI4id0YeDKeAQfPSN6dw/v1L
pZuW/JX1DxxP//QwHX4/FhLu1LMesdbI6RgHcMMnpufBTy5ctDDmMxzUSOsv
tgO4zPE/TFEb6huapTCkjzgrGzgxMn0eKjclqVXhufa0GnCJyzkziu6Z8wQZ
oZQPvynArY71i6iPWLMnrH5x6rhlgGitMlskxYMmRW37BWBqpVt9xHBbpTkE
eFT5LB7f5bisypMlnRYzYrkaGcQ3KQaZ3hQUmqixUlRBlc8hDBJ2bulyPSHg
h+usflo25b8UZ3o5Ikkb2UM5zNyNHcDZIlLbRzVjWZ4Ngqld3UAkiNp1qF2A
ATzbPlyZL4zj66T8C0SjeefIclX8bmqLipWJF/5BPyQvToVB9puXt4VRYCpQ
22c8PqNugHRKaDTQgRCEam/qqOAWBK278/m9QTOVz1RJrKV75PDyhdBZiECM
Xn5SjWVCDsWvh/CjgylgsBUpJVsL3sXOMibAEiHAnxmrO0mq8pzuofJF+OJE
7oDMYAavnlN2Or6Gdd1OekixAGogjNIlD575UA86YDO94nxkqy5u+3zufU/f
+yQTVlVU1TPIvNtwbEPSHYFq/13jp3dKFIocHd1MLFgbboUYmblNC2xWcZM8
OBrCUb9HiQteik0AhYG3mwPXC7gcYqNrwDAaoYF6Igod3JzbCG7BTveTPPxv
8ceZrs+FGX/GKndhb75OMkzYBez5AFdeeGbfwHNmOH+y3Bz8/Qb4CNp4sci7
W/Kl2tKmpoeTJ+kNDDjb7t53x/26/lOJ5jwjnEY6Vlq1V1G5DbgcDQ27/hmZ
/Dg4oeH9gqAPFcwYEoE3Xx/CMzBTQT+X67BOJJACLMM9q5rWzFkUuiOhoYST
Y61jMszmiKSidERcjklKWlkx+upt8ARVRKYETZ3YgBseKBbpqfflnOaa85T9
Z8wAg4gc4xj+3MKXWC6/TAnpISJhq++YwAOMp906U6mzkR9uKoKAhVsV7bkQ
9eB8otXLFexLcH8rurEd0czUL20IVqXTjhIzUAx8YhJOXRosY9HZQf0Xt8Hi
v/YuSZxLHH0Ctv6pkBmkqggNPiBF5mZjzDTlECZgfeKlJInqNL54do2pOVSf
Q9zIXkbNttTaHd16anoWqDah1ARPcb+8hHBI981GmDUL+/9QimLMVpYb2qBK
gmbzaR47SgcaLrNus3+/T1C7nYk2+zlhGYsbdBKYmXlq/eAplK7SLQBJSSnz
mFi2s+xdr5neUpVe12uQWzKCQqdqwNRaWlm74LGC4Xn5xlGUaH6zBrmVoGoU
oRnrgcNhQfPkvMOj1dsWO/KzpTz7vCSuImoQCljCjvaA33dhPf/9T0wPxWz5
6dxPNQ8Wg4tNF2/SSKkmzsnFF4cC2xMJISWHYpwtpn2UI/2ucl001rpGIHLn
2BZJ4wBZpv+GbLrJoQCZmdJ9cMli1LK3WBmprDMrhTglaVC9ASl8u5xcL9do
gfl08/F0tPDscy2ncfTQPJvxaAQDRY+n2tY5ARTzCJNrlglQmINYnb/8556o
7uVZ4HNzWRhRgE5JmAn4NnJwKRF2rEltV59ML2UUZkz0wKs8sGbPp06hRu/9
CY23icPIjRxpPl9foBZB4y5VYm8uuvmfAYcQGHhkZekOsTvIuwd3ilYGkhOS
xownUweAbvZL7Jt6QH0AafMkgCluZG4IFEmQgbLr2/EF3fz/qM/6QTJABrfN
fieRjRx6OJNiJBX2IZb9wKO8g3nbGY3pbA+iU1QiRQUI/TMg2XSsa0b6qmQ6
G8RvFmhVg/IFrtpjRtlwycaXDN0Jox8187ufHeeL6MmJ8RdEIfVP3vk6mjt3
solkPA9cbv6bxLwWFHCWAyplaSuvihG9EKc0iocizTak4B1J0Pgu69/Vmbi1
yK1CuM61nmHm4up2xGCm+mgj5UaythrBh2WaBaA/nwDy1ytyjzaKlDYzrKBy
o8zx75DDK0Kubn4hn6mFbq/50RejrFESIo85O5PZ5SnoFln6YExCJvqP1Lsn
nlqLGarES2i+f1GRZQdiUnkzEZ/qZlOXWL5ed7lhKmV6nt3reUwekL4niYnK
mbJSoG0mqsWm3/sTgr7lws54eRMsTW9Vw6dTDBiKsRteSrw59jdXTV7mMd8S
nvuGAQICnfSx5hYexQpILcFkQKCUNQuBPfRYb4kpSzIlG8FEWJwHqsW+99Ow
K8iCjxASfUP0fDqHVqo4FUYZa7PojfXd7RGrQpyLDIpCiZctq5evLhSMO62k
KLl+cuzYlFwEHOp0+k8+u+b9dAXNMJUkzxyw3UfOPGe+GVxJHMcG3aXlOO2E
VCuhOJ/mU9InxxhNAmU/2x3k5McIgOXFJ385VDVUwPW25ByWYteYHqg7E/bi
n0Gq9YGuw0mmyYy8v/yeFoJCR2dCnk3zBIUrgZ3S+XI9VnHf9xdzte4G91oX
Pvw+Au6Zao83DtXAC7KwV0wgupqEjULaAsSzw40MVPAqJD4GHnUUxaUaoyCI
rxWbF3fBwANdezAp9LTmBMyqHitP/WCWGWwudWIqTDRljn/ocR0EB9p9T2tZ
EhojxlsheY4igCAbjrr43F5HWSCAkindl21lwRhMvGhZYtXH9EtrbqtgS32H
19V1FxV06s7lHtqfD66xjUe74MHoxC/McI4DCx0ggor8AVqnSXjO3E1FCOht
7dsRVdaCodSZupLs71VGQ31Ru2My1av9jahpquUtfJsF9nUteNgKcKgXCVDl
TZmM88OP3B1Lrt9xfB0LXcp0RveYtjGWyqQZBcmKjxMJavKwE36gquFtn7hA
H0s9KmH03fMZV0xh5hWrtJ1RWwrlhT4Kz9NPqeBCt6bmD9v0z3DY9aqWYZ+w
b36Uho5CRNxxfIzf5PZk8BquWFtQuIz9zyfiUTXblkXxZRpctTz9U+9hwbuA
+aHrxIemyO9KN+bdl3KyhPN0nEBonWcfLLHxkaCv7kXXHGMPQV3WkfDtV7Bi
0daUv1G4+7JJjRGC/UrfeblPgOeGjiyOuRbCoW2kCu1jCHlt2OdTE3tzcbqY
JicSlFNB0ZXCOI4ssu87UeqZmOdPPIG1gxx/Hmst4lfSPEX8tFtfYEvy2IoR
+Gof/hQ8GyMXilwEXIjHt+CXNjvqLabmGH8x503Q1qfkZjiVpy1Wc+45nBru
cPM9CnhofzpVD1arfF6ju9mJSETjhMpOR3FDMJTpkcnQiJbhETYbrrt71nlE
chU0i35yIE/XAUmKBehrdHSzSFvmV9NVsx9Z69QD+C/oCf4Ix7GjLe8B9rgc
jT1k1gpNzLT8nZxUi69JI45tWNO6N8LRvkWn3NLBJ8Kfu178BWc4c0nCeK0x
t5KqXcE4fliYWBNsLQ9SZkM3mu2gU4D2tpsor6RpxVhRfYTPKssCPdpzjkWt
h0EoydwnUy4v7Gy+mtlWKUpIdwf4o8U3SO99hm0KS2VagWGiIh7UdBXuHGhs
Ggo+eEL4lQS6haqveOeFO/LYl4ihGsS2qHirgAsJ7QdOoeFLIt4WMFwI7i1j
bBW+Z2PMCpiX5EYAyqghtEuxlJrSHrfKIvcWxOJraVGaYgHEkI4AQp/fmWtU
ayFLl+4V3//sSlOnmTwzgya60jVg8kzyfjRsCNowiQsNbyI4PReupdYhUc4v
Xp3nO3xmGt41LW0LIauFUED4SW+udwvJP4HahsfcVGEHoycGs7izdVjBJBGh
Kx6HICLULIfFq9ywEgETM3EmLIqcOPo38GSZsXTFDDaPwdzuMGgX1E+OMQ0O
mfV+HIi3O5mWXM74zUvl05YOIkJZYUgIpA9/NCDMnYfkubmRmXKO7DANpoa0
4PY0yfaTUeYvYOBCnMNv5wayx2AsoxRwRmo8lAPA8qxSsXzBQTWPAH4FNsQd
4/oGOaHAKmhOArlzLMOsffKFcZN1kVGzZuwW5FyuLJZKrsCW4GsgXlkYiOT5
00qGSGQnzasBse9IUHMwdKNTLiIxFlqz6vC9Qo8kyakNDyu/o0zIo/WAgbYl
+Hw0sGdaVIwkiSMdEzRgK7NOhPeScLO7DReY80wpTmyeikx7NBcTWAH45HxV
HIV4ZtsIlKBdVcghzSqEe7QMVyIUBzdYa96+R8mJI16M7sBDPVqj3BYQVkSa
hSjcfE+vDXYQebIXUJYSdFV2uvYA276FchyOxtMWGtjeDIV6fgEZtAXxJz/r
PUU3vGn6bPR8JYZmdi0P8lUoiDj7SeygkNCUmlDaZ6p6/IchnjqGdnCUgsRI
z4Pg46oRHmxCtT+eDfd3Sai9Nv116CuaickrkCqY73PXy3NzvQH3JYwPVEKv
tnEI8oafeYnWoS+g65gurqKNptyhn76mWdS67OhWvqZbdwj9kzgCCOe4GHKn
gXK5WaYP+1EUNKD9OaaHuaCcCeTotKpgCgeGKFfGdY1rFcXHCmzZDxKgSlkV
/fQDb5RuAtlFanpPnGsegdTyA92AeRylJjRbN9tfM92ZASlrqKoJCkfbzRVr
fXilpZL+jxhRGQSpBtVOSYm3kG1t+qHk1ELma5vkrDxhKVcY1wQe74JHhTrg
e7RCMtO3QYJk92zQHPBpl/T5zZdH6wCV1aJ20oJ1agug81IyY2jbm/+lq405
h0DTLq8Q4hOlqzL2WlidONLZXYKgpFyKQuOX+n4Tfwhp3JIVuXXDOBxEPB0T
ubYch8bT+n3R2QpV+ASbAJdsViay7fcSDhM3rn6IK8U7q7LLoRQYa/Y3c1na
q7WgAIBsBuQLThaQt2gaQMUQQB7VYZt21tyOgHiftMsVgN8gbtyroagcJihQ
iowJWu+C95bq9JBQhBiY1jQFvhrhIyTDQujVlZAGMFE6qSMWa4c6VKIDKZH1
OD+wdI2201bonUBIuJstP+oeF8wq3KvOGFT9D4FGmLuKl05VFxFvktZtGxL4
kDt/MfN1XfPXKQQjLQ3lL9laQFiuCK2h8Bf6zMEcUvieyhpL8XhQ+NODLm3f
GKaZxB2AKEKDiTVmwntHEcfBofJ0T5AdpCoeistQd92afP6/1wUapi/uaUtx
nMGBKDbqFbRGje2zdtSdVcKE+YHx21K/mjPaDMJAhYLCsY4vlIi1J0qLU728
3AzvrmNRnsqoA4bFQNLyOH0tVIU9jha4dZ0+ggf9ufgtd5oCdPEZiXk9oeeB
c7XJbhW5GpE1AHmJ+deyMXFH2GORSHqFnl+8KTuyaZfHKk/0fEQukhZVMbm0
n/lwy0bzRNw2SJvmQ+YbGcWaadZLa1X8xHYKHTHXDtL1tYq8iIql8NeQpwbf
ty35ik4y4kl+Bmwkcj2EIOeSiEvUDwc5O6H9I6zw/2/IU/vx9NiwnLMhspEH
LTDzP4W6koe74UDTt7IKzL+marnoP+jeXGZiaYF3dpFUUNpjiPmZ31EQ9fh1
hZMxFGJoNFtVKo1B4niwYgh+VavYuoLRZg1CrpnX4v+hXj27TnBtj/JorkUS
0HmqG22kU0xwFDgJRt1W7ItZhGlV5YXK+wpNVh8dDG0J+aVHmqxZJt7iIiSI
w89p8Aawm4ll6YuGIIGo0nrp4ltHDb1mfCJeEmzVh4kWnoAptuG6PwrHrE2U
EjgxFImVVjplfQ2jHejvwxCz/PAqZIIDnUI1C7EC+xFFqTN6ji+285sIL6C7
fpWNnjPzlc/+C+qCnhMAH+I0R4Lf+37KAoievanYkP+f3KvPE33kpdbXO7uW
8+RSqpM7NX6z4mZwdhOvatzewnS04BIsvX/85fjCHl+FnU+cNiDFBkMpLr7E
kAAWny/rJ/zTwBGovaRFChkDSFccWgeMwERA+ulpFqxDZMhTMLLSxBawW77+
gDoGBxBgsCAg6nEpWRJuyfWHd+EOI0elJqK5DkpkbzT1d83KH5z1GHUnSWPr
iwRnZbGm2ArlTPpVMZvqudfP83UN+M1c3CH0qeGyF0TkyAGY7+WJkbEUJmZu
21AYW4C6xj4YprZJ5+16tLAvAELLuMt6uWfpVfVPnPBea4MLxLv2hDGxEqWF
mSugm1SiANIyz79+UKTXQdY97P3ne9GIFAQEEaqeqKrGRfYzLbpnS/vOn1h3
dVEBURcF5NnJEuREXmpp/qDKWCfd3NrX+kVocT60fQKARBdJ7r4Vmqt82em8
qy4ce7Bt63zAgtPHr/mVBVjTPJvhcjcihbjTuLHw13UcknrQjmGO7fuW029c
5GiOVDl3472+p/DszzGosO1Lw4QBURkeb+HEYBYY4F4BFdUkzt6SWL48C/4g
q90jCQrCBK8V8daYcvgyh1Jn8LJUX1cFl0ZMKK0TQj9fM9cnkWNzsGtM7V0H
BkxFlp/rXLccalf6Aui5DKpsWPk98+gG89aJCQlksmT0JApuV0fSs9llCzbo
cgwe3cbxTSXGdI1rdgJUtDEXtyvjPnUiJAPubEKh5xFfyHtVnVKsSi3CJN0N
x/dGQzhWcpfaEAKMMW3heQ++V3yJzs1GiJjoU1gS0nRYlvjaOaw/G3wDnyBO
CvnVvTPBk++fKXzEGvcf5/RZ2/UzBfuAF1JUyL19u703n2RgTh8Kb6+89xY2
NSffeKHBwxJqTDV0sSGGXN9q2fDY+zJUB/Iy7bCSpGRkmn3nNONfU/NmWAps
+UGsSGuH5Fx3L5c3NSfZKmzFC8WVViEReO0dRZGLVbNK9qlaoJeF8R4viTyz
ze7eAB8n37/1IM7AiRIghZwXjgmOcixWKxXERCFsqWaOOzCY7uSVfpuzXPr6
DrXUI8YTMnO6C4Z8ZgDxRz8JO7fA+ATxpEfLo0ZsT/TMENDlSqWEjf/+EoJ4
rpChfrl6T+NJ+jre8UjdxbPAIJlrEypuPxK4lZpfnpk9CaCg89eLi/AzJYiC
n0kS+IMEAngTO2/0VnEulqTRTpG7Hla1wXfqeRfwJ3QlV6hzDBodJvq+Nd8L
UE/w/GwGTNmaDqGLkUul3c+wQW/E2+tdVriCpFTLcxlWlI1z2svYTT+df4vC
OGRixOQcVtKtYytf0uMBdfaiPxQIRQz7b7n52SA6TVq1e75RSvVPhRZ/IXNR
JHFIk8CfCCjFTBw0krWvoG7kE4hqb8BbV+XxebZ3zcJMBf5xEcZoZPi5ilai
3w17s2rDpRgvjmm+eayTn+l2r/di7NbUlryY14N5ufry563VSYV7Xa16nmTm
uS0lvpy0sHpryheJGby+PzgCTlCsa7233UD12GnYYTgAYwHpPE0ruUVG9iiI
8zft8y3jfKQK2WjfYEq66JbWOdbQ6Oh845VcACpv9dOCZYXfX0TWHCzkOLbb
it551eTOK51RhJ3F06rENJbMz/puZPrqeOkBs9bB+A9Fe+hs0QMcA6qIXkyh
VqcrpxVEuaUG5/aoYbp2KL8CwZH8a3yknEoJq1J/UpkdkkSpCdL6YBZXneuC
dtzF/JN67slz718upO2eEmZRi7zFQ8yLTh8itYtSC8yF2m7KNOutvnEQSG6r
aiTJYLDz9AqiWgweHUMZEvtSXImoTa9xVQPeDFcgvIDKii1TIy60eG1mszT9
TRxKRd+0WEspyYjZkLWW1qctkGjZ5ddjbB8Ed7GESod0SprB17/2WcsQUcC9
vanZMtNBb8mVQU/yaKah1z0f1OMvuO/oRhSssEFKGq2KS8x+vsNJY/0B4e+g
FJHfgx6VY2dSYGZOlc+6qY9woaxqqEedYPOct8p1xsZj4Zek5bUKeHnZiNtp
lOHYpsl7lh5izr39NOj1i5W38XpGPYZ7f7iE9tM1941/wyNbI9k+kQ/oPto/
HYs26SrkdFhhFOrf34ecoTZTeq0to4VGYOFarrSJdGLKHThjwuFDoA01OXB/
O4pJg3mbKD75NuQUdqybTH4VmnXUUrNhZco0SyFFmvMSi8f8AtuVbj9MPpMh
dOsCjyBmpNrrDwFRu46hKcLbLgLPpKkRy7Zx8TcdxvjU9nw9LxwW2h+ZU7mW
jp/Nlb7bC1snBQFxPeMiCW2z4HF1FHSolw9aw+nY8QZrSq+3Df1FisnhNWE+
2H8OHPGD8V+kccF5qABhOqq6ex6zzfO5cr7EBPWHx9G+9Snj+NlypXYQJ/mE
PM60wOsoYBM7GsVy5IMEsa2O4DCXuteB4LlwYcU6WDvcC+B58VYef/VrTE+W
qrZqAH+yS+dbyBNkt2B2A1rjJ3VvVouC99NqqX4DrHxelTvmHhr6mi+Therp
ZAvChffJIA8ygZwhfPTYQRDD4jVcqnX8VTIZ4iylut62e9Tvj0qq2Jpo6tvv
puMuVRQ9uMOVltz0UbbYbyn6XyA8wGBSnxiVPb39VrR+7USl+iGSg347/dyh
rIRIz5JAlwIoMJySHwGN9Q19l4brs2LgRxn+CfWZSoQ5vX0+qsRPzuJ/9Vz5
7H/XOU+uB02E5yGjkI4a7fP/o/ZNnaOhh7fp3lMF+boOmsR3RD8s9F++TaZC
kcSVnD5D+q3yKtA4G+VUnfXybMz5cYaxSyob/JyIkH/KwOky4GbEMsb+5tlM
HlSQcYzamG4c9MFiv2DXObT6zEbfARqCRJKwEDpGiHdm86pqBbNJzbJU1M9D
gSbbz4Vic3PoVtxDh6bscCTdePlgXWhdIJ/9Z0vdJM7M2CLfMroM8//fIrzE
aAji7Bg0NlQ+ZmWSieqkyF74Ifj+Oqb4xMuUd1NZ4St0B1JbKXAyKH/cywBs
txJB8K6n407S/44Kkh478gIyovsAePzRpG3c6ymyZehNHmUWqgEGHMYCQMQp
QF5rofPgjsxinHM9bouzMtfZ3X91DjnB41o8FxzltonHVQac4mA0Q6sMQz0k
92tYaIHD0ybDl2S/ZT9hprVvUkH+lNUdRxcirJPqZssLpuEW73wrZSEf3DgX
L6OlXCDn+jSy+1Ckw58zUJxEk/oZKxq5EMe1JD1sBz0sR5WJAZKOr1lbr30Y
1rB6MtMlDLZP0vXnLu5Uu/BWzkPl1pIDzF/fZ0FHri0jXMdw8TfdKeIvOjLS
QCPzgFRcvhgRmBAqmwhiF3Fo+twf+YwoGMEUQr6ykepfBc6mhtMmPIh1MDgL
+56dgZvs+4If/WQhRvIAys/Kkx3IQeHttOZGrq6uo93uOOGmC2/nNRw8c8Lx
T9ozdKU8KLTuq49uaRCMy56AL0LayGZb0ciJcsEb5328s/rydkLTKyaGKIRL
DpijtzCZ+ABo5qozasrPZRdE8iKwdrJoC0aaPhIg7g8I8QGEsvJTM3HO3ADH
fJks9AdhKHElQT3WYv6CQPIe/CZc3BuRncvjaLzbdSHz+KGzyKvB2qqNj42+
/W3g99A/q1nRP2W8X8NYL3QhRuk47vYZyRrJQPhN3WasdRSg/qX6dV/WWi9d
YEiXOeOGVhdPi4gYowsZ2Dmi3YzxSVNmvY6B7u9f77QaEKoeUgN1unQukeV0
CQ4X5CJ5M5pFxx0gJY2tlObYNG7lRWNlNL+e3hOR+PkeeEkxamye5zHaY7SX
apHAJzW7BTkfK7QbwMpBTs0QKj0+Bwa0LFAofR7XX2ynm15FTJJt9bS2EKZK
/taZ7OSY7mHpv8JjS5lRsQX3RWmAVGpkZGaprLFmGBUrtWnCPaoy+HnGVq0n
Xcrvv3UL28TS1AUOtbs0JYgVX7it4LdnHl703YSROSLan6vS3N1alS3HENyp
l1YHWDEL+rwjThbu7sJ7WgGNQXIT9Vm4hPBKNysA1FpvOt/0G4FBa3zcAdos
JWSrO0bSS0nw9747BRy3DfeCLfOSAjYyLo8LwJRqJZYz+XUWGWi2XGR83cdG
ETZ/HQF9y5mMlNkRLPZ7S2S1pwwB4g4GQ1V5ddB5QJ0Z/i+p07rHOgX1ATj8
3HVezkNyrlthFPISqVSize7SNwLdqLXwh8xHYVY+bgw/EaV5etcRf8bjKRJH
jd85nK6wCtr/yCkXsGJ5B/kDTV0UhY4Gtd7AVeogv9bvNpWiJ1UtFdvHezxr
v4gM0Fg5rXUzHhZcZoMoM8fsuq010GNSdoEP9Ok002GJxoyQrPjI4lZ6KMHH
K/LUcFOxnasVwQWh72EKIfSBLhy8Nq9uUk+YdDTjJzkGPdlr+tM4Lyp6FtCk
Ozfl/0YuaKVQFo08Dk49x+4cAFiqD/uHgQOEXDPSQxbzBCDTHrSDhVMNIbnk
gFKjWTHOMCEOXx4LMFCnVKQavLG4r6cWEDcNBLIKCCwfqqdxGztuEIUz1iyA
6Lo15FwywAluWbuCMVRnWhUmNSj3vAO4f2WQ4hA6miC7UhyGoAzQQVmKvqwd
S9on6F9ehoHstgnrF8BA/l0STYTTJUzNEUD1f8poTB/M8bmO1mU+CCFpO6RM
mdZ72llzTRbG8Kr00yWD23ZTvmc4Dv2WJWZevpH92v+yGnzc8jD97c9Y3GmO
RuORk+Op4ylStlq9SkKvFas3ukS2zjAoObbOuwfblRgxH/6SL+IDYjgIbQ9h
bkzXuIXKOoyYz43ndu5/mkjdEHUb/DR7bLesL4geTOInbhTzNpeW0DAwke5T
SeWCRrjT2D6TxgsnAdthnz8NmgU4666JCpR7LTPUEHIEIsUy9sSInIqB/qXD
Ec3k3173Me37rvLEpUc0dgsBLhBmixjfy3iebWN8NLGNw5uzjpxAgV5J9L1D
9aM8NXEwXOJ/jV5AHtZZbuQmuQASkG8geqx+iauuXw4v7QU6Vv6NtvoKB/4m
/07D5nty5DuEPK8EUVdOlPUngiVQ4IDEwN34padw4WBsVpkMwCIWb/Lb9q+H
tSG74wzJDaB8pI0XwdOGVewhuHDZiMEpW13MjTHxYLMdVtopdcGkcfhzvj4j
cJsF6xtRjaUf8k7ZmAiyOmMH5o4g+ZcR2gwReFh+e81UKkjJYCV9kUoz+4K+
ROadWLmEDLttuElwbpt443NkABG8PIrnhGcIyqIwgjbFv6Ph0lPeDwdLXCQ7
tlYqjUuMIce6UP9/bAaYP0uXpclx6TmXtDiUwQnK7SYyEKFf9OV4rx0ynnxk
fnJBYRZ9mYnTutlt14goLXAry2bIAnRJKwR7m2qMXN9WTVEpTKmafc8LiAlj
bhsD45hJk1qkECdj1vFRRNf/OhCAAqpJO0fYj7ZJ1VDTZRD/U2ipvRWZkZJf
Vvs2dsU0Lz52ZGu2qKpDrzi1M53gf6x+ctjf1PIAeos8+AGs+SdFXob7Bi77
BUiUFysH+Rs7APhkd1smwGRKv0fjuZ9mrp4oZ8JM0nuudsmF8ZU/MhraHrns
h4s3v3zJYWEFy+oeVhuYZ4WJvjm8S64E9NRojm2fJ8jJvoMwFy2LAYjJMSY7
wyY1YwTdvb6hWnxIfZNm99O/HYy2SkMXZLuosuRyevPqdkLYZGODQ0Y9Z+r8
asED1oHs+W6wCamdJzulKFPZ4vCZp7NgVFXMZ4YLC3b5BZijUMexfc7AVN9B
F/DUIVXXcAOrcRZBt7yT9iFuJFE9hVmBxvTyDMQ+K0sBJCnBzzqipeTclCjd
3alaC8ttItFBCdIS8gVV50crxuPZJociJwxiJSkQWJq0xA8nJZApDd02GUmr
3H6x7xk1RdAb6i/ggPkeqdPmaSITpT0Ifz3eWV0eB0bkfVDQ+SNBg1SXnVjd
pMSfPvb1Du8qfQVV2WXkpArMnQo6iWnpTU+Y41H0SXrH2mxKKYz/VkxwafdA
xJFlEGdi8B7bGYwlEgPuT0WxaDC3EegZcniiAgCU/59flsm/AGotP62X+os4
k3G0pbALnA2OZICG9S/Sxmr4hXQP/ABDcOU8RAv2ADWvQvl2kZc/iPySx7hk
Bsb07MD1xRJfGs0CCx/Anz/3W8Cb+GxA+MI9uwn+ic3dhgYPEc1jzbudKmLB
yjUlKEZ9oa7airHaK4yb0I/+k2qVeswRkq5j6Tc9Qj8j9Ic9P866tkLuMxjB
QewrmgpIa5lF2+IPu3E7XGNeeffUsvN7qoSJ22gfYER+2Z7bzbTS876+i3LI
72f2JtMkDi0j1NWcEuZfS/f7hLFdwQLgjtQqS9m5DzAqdPlGibhL37ACAjyf
JFWkSYenhvJo+Qweme/xF0PRXiWt+RtT/U47woJoxpjCdk8einyTc0NIpivm
9HD7pCTz06lqnW5pzj4VQVJLqDPoarlPlWlksAMlHZL47MlmOb0WRmlMvtvp
NqTNOwd74PlxyjLZQ7/pUiQnwCJPiwbRuWWc5qu9asSUYW9RhmXi1HYN6giY
P4Q6hPINq4h0M7JOj9hDQJfSA23ruJV7eoSavvUdYxSGZQQRMUSSKkM6QEnJ
Oxj42jQ9cmWibzJdn6qlAv10sbdZ+iZVwrSbcqn7m+fUwuZ7oFJthrZexeeN
PWqaE/UuGYeGu09wHtDo1EyIeoI2/u3ejEtpEv3rs62haMCtB65quEUmF0ol
aXBrP4JoFNdJfhB4jMrT/1bnaAT8BepM2UHoxVHLMQR7NT9+4xgQRxUnSYTR
dkZf+HFll+q2GKZQ2488ctiIHrb/dRGnaeWRzIIDhI22UgeP3BZZdYv9i+Bp
Ru8pof2y/y5N/MQPPw3uctzrB6trRitMdWZGO8XnSlgMulpqiELs2gUzdWRr
VJVxBGQ+KKf/KjSfDZlyJhU1NNF9W4953hSLMKvI9vroRdS3uXYPz5tM19J9
xDmP4qNkNJvm1UyFO+dmCLNSlHlieb2KDtvgcRdJSqRp1Na22KoND71Ynt6j
O13ivi8oMxOXHk2zUvNvv/tx5+GG+OWSFo3RGw5eQdNaICBEfy03atJYG3N+
IhvT3KWs7jsmh3boR3zTmuZDRPuISA7ASZ+6qLNoxAK9rlXRy5Tz/XtfkZt6
xFKH98imX/K3GF/WPhe2OSMqCjmpOk9JKOJ7pqVZhH/p2NNn3Zd0wA+zr+qB
50RZHZWNMeGGFxnSJfvw9wK49iqZ6uw4U0RIWn6nx9fvl+MnUg845gzc2XzF
EptzMxtNp4AM6u+NEMfRYsi9td0k3EhtWbCMAljA5/ANGn3jYkojqKRk0osX
E3kMeYIJWltoQgSiwepdWZR+TgboOfruhac1zuIrS6uvfMuxlluHWfmi8ex0
qE8vW4WNu72e1aVyZ4FB3a/qa+f0GfJgc1QjWWttnLauos8Esn6J7xWIwC9I
ecz57i/JGuNDo5a+B0KmSoqOx138PnDSM4R07DwJsMRzLyLtksXd02z6LgIA
2Iw29pGm8YY7RAeyA0FH/2uwA/1cFHqmjaZ5q9V8FQwNFYsV90ykKxxzhtqL
35XA14ctrFyvzBq77BQldNPlW/7WpfTZemkpt/rkORKP06Xg94Ffgx/kFAfJ
+ql9axXcXdkUh4O+J02yxpeEORoMaPnAMICY4zzRN+o/QkH7tXG/GpUoUVR3
k5KjXk0K7RUKJ/DQb+/Rog9jlAQsBenN7liEJDxA5ooD/AJLUgalvT8A8MGC
uAFesrTDYacm0+YPj+Zb/U7OD3T2hc93e96kxONgbZu6CWrOOGLOc5P0QdxB
jQ6ZxaTjg+mzCxWCt96vuqmjvhyIOpsdfc9OcmleS/6sWx9D195vqZ9kfZbV
uIZniBkSWyK1GJKsu/T/NNcoPhuswiQj9hBhdBF0TEEFLtyFOQ/kLo9KiF0k
209aMxgz4f3gtDTt2McA+xTAIO+LvrzM7vSr/VHsi2dKTqVfPcv+Z1Vg9G3G
kCXeuGPr7fyBOeqfUu110VA/eXcM4BmVgh0XZBO3RbY2zMWGDZQH9k50zhwS
S+Afm8KaKjaGWZEU7kCo4vhsvT6YZm0sbwligiNDZdha5FGWHVtQ/auOIazS
KPzamsYS2gJqU0yRSePv23EAHPeZew2lJrw+/hn0jWpWydWMlUwBGMaE897H
hgK8cTggC7NHAkkAITeekjC4NuayDtkkz0IgSls0j3Ukl5aZ7S40L9eunKfK
MTGHw9hBT6bBSRFiTRRPUsBrVZharLKb93JebQcSXWgTwf3RRPOZG0FjyVim
Xn2+4tiBc/IkUmxJpFn2zEC6auVJtRZrx6h/hywSTdq6kgLDxpJFAFVhucNa
tOQBF3p6LyWeA7OwR1KtU+2lOVyP3nIeHOcfTZfaCL7M1armVp9yZiwBZ2kc
L6nCB3k2nGlD628f3vIE4z/UYmkyupeUmuPUw2Txiu2DoYUWs2DIE5+ISEoM
9NGJx4hlmlILxLo5vEGrsoTDJSI53X+/xabV5FybuiI2jzklCo5KcJz5IRdS
9W0e8Dz2uHUaKLIWroAzgZxgvz2BIWhPaiIsG6VzjNRc9m8dYHhFK+8/NZ/I
BFIBQEDY6qbba7vk4fKQg/RDSctiSqZhATmMv1E+NfD6zE/fbI+87qojLJXC
21dduGuebsChPtNeBuUWoRecynaVL/N8g3zjIYOhxGQ2cZiWtKH9YCZ+hOwb
JavlqyVv4Pw/ykeaisHzNmhNPXfvNhT/rmkAb29LgfVgFEB9RhffxaJY+PZJ
pX+v3fmVxe//79WwuCr0jPFYk/lsjuKCGJKD7syxnvgEoHty46s+ERtGL/yE
fbxAn4jLUhi8OrgTKTQHtE0GHJjUyMgraYBnK/4eju+5VZOcu0sq4RH4tmXk
LYsjujmcVvjx/fn6Wt0+EzE2TilmJkDQODmUcoeYYKA5/WUfzYRO9UapDdGn
FGl5ml+HZwNJz6GPVOTWcfGdSviPE1rZKCPf0p6H9mou07d9oN2tP7hf/GaW
hzhXBicR2vHXk+pkRewbpT2eghDO0sOXDe/mAFsVkMrsoafrlqDHA88hD7Ba
pJ38zXvWTOqvBB0Jd3Ausq3dVIOD8tEtSuK+pJj5d+l4QDPrsE/ghwZ2lFUH
GMkxh4nCeTtNTzEV3kReAOZgrotOfdvN4J7R8PJji7C38CNLTFoIXwqtL473
XM21vA0U+Y7eWWITL3ibAsBaXJ6KNxctv8MPhCGSZCHQ+vhB77GeUVAJAl2y
yTQZSqT9IUG4yXDNGSZNp0nfY482o9ekNS4fyzM/kvC6GyrzY+a2YTEfQ21b
PcgLYOsuLSDf5b6azKJ45ogyln6qJD4YOiGBTOFfOyRAGbVh4YXQXeW3EBUU
7fk1YEepUveMsPUa/V3vzbD088N/0GWwtk2m2qAEQ1YSX4fshys7cUcjbQYc
AL/fM+FQNm7bFxlh8mYOhP1pAA5RTvnkyt6/I+O6wDxarzMatDTx82Tr+y34
Ef2q6QRa7zyZy94CMY/I60NGoxZuEJNHoA5yY7A8LTOHvAkAhZsZRHf5wRSS
u8TQgybsgy7EKtH8LJ/wQBCKQXfAdS1l8D94qW9MlGFBRhpKPwpLylynJ+PC
Ci07UQ+U5OcwTO4EUsq70IAn+MBVF4ZdA/JjBP2swJRedjUc7/00MXoYB4pw
jakEr4kGfHVHiSEV7f3I0z3CArWaUmlPouZLo+4l9Xxw63rU3M/mzN8adtDO
P6TYwbM1HpNwRXNCU/xw4uTBON+f9gL6luzirt41yt1tvzM2NDMxrzOLdlpz
OYM5ti/jlyMXeQ9frsYkof3W+fkyUgEIKTi2I3U08ra/efkqNGPDoXCNByhY
4lLHGZY5J2xaaUsZSKNeTfuqMiBgLF3uNcsRoogLagiK/3xEcMS5ShsDhv0O
qMVfiQK0wmmflSLpQY/ZNgefwLuBCHSKjcTKfZgTsxA7aJpGas+3e+O9ph66
AJAKjes+Gqaq9ettg4xK9J45wX/d/Id0Lzssjo1IrfcKte3wX79MvriwQMzS
seSJjHlLeM8EMlrOqdFKMQwnrwAVwouPWAR0SWPAYh1ME8io4yDTZpWp4T/L
m7sqKaMUsfuBIt0+4PT9HJoFUkGlNX141LPQjLr9OK02itCgHAnfZia2SLih
LFxCGb0QqrbTpAJSUG5ZkiO4q3iop2H5JO0EgMP3CkwtZF4YWdVgwxxWS8vq
85Jhay8vH0hpWAcjP3HX0VjrTLej5ys/RqMy52u+B+9sKcaS/O2qDiww+4XT
PrKxpeTOLyxInwtoErz38bY435qXUravJqIHhL+LR3FReGKT403410+WZe0x
m2p3Zmr7uCMzBPH6GaDQZndTAS2XKZjqI1bdvDw7SebU9EY/YXajmCYgP6Dl
yjIcV0NX9U+7qmtIf9zuGld5IdDvQPLA7foiPlJ31hSYDQexW0cSc/Sd5APx
WOUHqhcp4LqUylSIerm9c1fZNuionh0Vt5q52XjX8ulHDtmYiw1onXtpCk5P
o1iB0KhW4Qt3o4qq2HGZqzvQWFQ7vO3Cy9G+yv7pSQYQbDNV8yyOaYJe6ngi
Mh7cVVWD0iY9LofT22Rprpl+rxgvDU7WoXRqZ98t4jUVZ7ryuac1hHBpyXjp
wFVwHL8xYiG7VJArn3Trid3oWxMryVXzh8YMjVA18QIKtL5aCfjjRp2kWWrd
4WqGB+ISeHFmlqswAmHAQBvYmjLBHarsy/+mS5TuBF3i4U65B57l+R6BYBUb
dC9VgaaDhRmftIpwBhxoVltgf3SQqYQyS2MlxBl9nd0Lm+BUsH50x/WiUcFN
MQ1YRqfbc/sD0VmcVXdsUtQcXHS4Mj7mGxaFLDXjjpNY1McAN0LuvnhSPi45
rPgFiRyL9enLC3pnxbNqZHgoTliH1uEI/UIlB0SnNzVnyZpwBnI/Zpjqmw7p
GjgE7R8yfoTPUtKB/kK65UNkRzNqsXOZxbH9ygYQkcCna4VZtdIoODjseqCR
b2uCMkUbhLpgtc0B/op4/81r/5AF2GGY74YuNLGEXLf6pm8sPjsW7ZKbkPkU
5iEICiLuziZAj9/xrGXKQZPSUEvoMnUs65XlgE9kvPW2INxe2AhI3uO7dvar
bu39FR0wp5xEfnLWIV5krin4+kDzPcDETf4qVPp67zJE1W6NcS+g1HGnuxfx
xk4pAVISA8jZoZmgKEfbUunzS7FKYOVFvdX6GmIaVeTX61fzZm269RZ5UCFj
wt9JuAKZ6bMW1z9wvmpFXEjMsSKRuYSg0DeNUKOY+E5RwxA1f+1H1P/tl+xw
HrV211kHv3oJvgBQTcDVqdpcarkLVzkSGLjZR4v5hy3ZW7tgVdNjzscXU6SJ
NgHJApExST1LXWymnW8ep7Sq8V8MIarU0Q7OtQgzLMCtBNuu+M7WTNTHmOLM
8AptMk+jvV0teqhoTRd0XLd/HGertJY03FHdl3DSHhmOus+jque78xDnLMvV
Kdxd/Dl5P8VsNtGPMQ5fHuFF2L9GUs7LNNL0Y6X1S0c0uyvls3H2bO09d07+
0gqPQjdyuDynHTJOyhf1tIwFg9ZNj5OUSPyjGdTGq/Ar6AC1cMCuFXWhNK+B
iIhKut9iXqhzxTbU6ypy/Ly1i+AFnVO9Y1PAOTRHnO/Ja2uSexjFkH3QyE3g
v/xmBeD5ij/U4/UHSgIGUHGP8s0VdYS79+nkFgIUfMIrr7Ot4UdT4tlIsaMZ
wxCqqV+TBE0WppSx5GeyQfUfMv1cuz9g9+HEfmy8lJtCZ7201+DpgiX579RG
3nEEZXUJMaVwepSbpw73UGWqh4AfSYGXgPSm9mfOyNk4HZ9Mw9VJi/5hG0yk
0Dh81CmGMSty+/MkmGPUn5afaAzjnhm8wahIffDfRLHEBc0pFTsBj7SoLAsC
48zXUaKwz4lsXgAeyCDfrAbD9lusPOm5dKi2RrHRb0l+2mZ8826b1GR7GNWi
NJdJ33e71Qvjj2Mr7rAfrIkg/s+FrG0Mzz5hElw2K+X47CdGX2qt23j9AIIM
lg81NXbx1m34hHbgRipE3mNhxWdsBrs9qgUGebERMhwXCeU7g69RKIOyVEQC
l0jaRoKz8Xb7hQd1MJfj5DO98FXSoBRJ/fjTgtx5jDB4oV2JPW0AGr78wnpW
t92epRc7AbH69mIqv7HIFUZcCxUEfHmXiYLhXOV2jmsx2VobMNPaY04K3/BE
kvRrkGgGeXV1m+EJuLzt+tAUeW05aiJOyC2Cakbv7F+tbDPyymVabR+0bKcU
hUV/TZKyB3D74lg/YRQjIoTB8IVcJxpNeZy6gxLCbdTGoxZah8jyR6ZY1ZcH
Z+KhBOmg+m4/yG6RRyu5RFM3YKVIvknvKK35nJgSuH7l+AmsNTrK+/F0gzLb
k5FlczXOO/JRhPq0STKmmVJYABQEqwzfmmL/zD4Ncn5VsgXa3+cRUJhdcZjf
EkQxCdUVNIkVMDifS+kF/o1A/6Gi/VixcnD24MdzxZZhUkax/TNmCsnZrQ6a
VUTpIpquXv9IpwEcSXKMcjsQaguwGC+rXnvAcfwvhg5tczsqn8s/+7Eq66/D
su7D9P5mmWjwbeqdHGDKbjnI7MkxnMNqdmUCzOMea18yfc96ZOAPuYoMOEG2
Rjgk8+Iymw1r2etyB0/gpHC4Mqq81eyfgVuBnKeg7aZA+5Uekg1f89FoieLh
eiqVZQnxL2fKcoleys8nGs8aq9l5zipKButUwQbOV6GYdqNsRAF6boyB2JW3
nwLv9bI/qPzVnuQmUY0fdcmFFSPtLsMZfMZr7c9CamY2xq6A1nAluqtufSJY
VfezSlZpDnJKe+f/rBImKX+lyXuHN3JVnIrnhinUlBSywPahEB3L82SnqUF0
Ttoygfz/Mi5fwJMnkxJnRgSmfx6FUj9ONp1h/kAY2hDza6lTsMApECPXdqFq
60AXJxM/+onxMrB3H1e2RTvpYFEJNvvjj8ZbwEXl+Z8d5n0R7SlACPQz3r8v
6SbJ04sLY6cYLiLWY7UKw6bfmahz6frmgb+Ftiq7/qmUkdslaeMUCclnyoz/
Uf6OMh8SKw/w7ZfWgjzQvER3OWJTG/RUOLzL+gtkcclu1Qqsp5TC0tx/KR8b
TqZGsDm80yAJ64nOXpJ18IcMiIbYtYzEVDbwRkDxiFPoHFvTgQ4HNVeGYzSF
XyJ0mf3oiZuUWJpyRFvJCl5OeLDwpwJbhMJVfGfmsAOB2/F45eqWiHvLD6Q0
mRpYzsk+27yzNVPBcil7eSElIiB3j3EYdD3m9Xpr7M+Wjzv1ae4op0Z71FLz
tCspJk+3YvNjrYEwn2Vnve44pbdnn36b/w7HxPNWdKeUV1yJl8WWBn3rvQ8y
KqgJgcY4ACVpbIHlhuEaA5EWqLL3LJPb+KAv0gQaXjGNl718ZxmaOL7+BcHK
J7MPmglYj9TYD1o+JL9D2Ydm4N52pMdcWFo+MfCwjW8OzOdr4JgadHGbV94Z
0wSvyOsT1LGZeNUhIZp2IOXWXMaCI6YeLKM2JUJKy2zwSdMLzLvM9B0hlTWa
InVDet2xEO/17gpj9kA96X/wLlwFNpuFmqBI0dVDjDBbAIsjxgUHNKehBNmv
prSEThTu8b8KDI0Ay+ybRGML/dtWNXciMnJTnRCbO01wo7rNPWA58TgZD/RL
FmSHsAlmPAUwctFjardr6ebvT1kMRf8y+dHbtsxLnQXJEmc+7DdJGwyvC+Ch
7F2FiFa7qZtKd2zaVZq2J9CyIn10FfBuXZ0dAS2hSYF3Tkpo6z6ffq0SMhdE
GqTtMmrKbe+NTBE9Am+Kh66H3QgequRWJZLBY6vZR6IZo8VaAZr8Cjn0E7X1
rLjCYgNkxcLSNUoPNZz0MIRbDEEQ2UT1wozBTLf2IEDty1xzQXL4L2PpujxY
udpvb8op8+DVVpc46SiZv//LPoRDY7hxYKXd4/a0LB0fNiIF6/5puFuQ7SK0
NEsWKhFJJPmBO5MOSUmSUEAPTkplhodFA+XMOFspAe+QOOs9w/M+UDcH2Bw0
0Y9oXOAgobxkEKdTajbRrEejoQmMbA4RWu3k3QaiW3aWhbvBCCqTlfEaqf0P
DOxbEQ/GnYbwD9lVtQAXK6QoM44KJp3w1ELzL0mjoNthTPWZ4/XGNXS4WgWo
kUBUrff7/F0f10UkEasdTxA4i2nbe2/0O5GsUB0w155pSEH9dLuuk0n2Uq9N
/MK10mLL/m3DQRVEYMZWlJfGj6xItgYw/JRbsIA7eYuvPFhUEEePpQ9gDpWd
GYaMqJ2oJyyCAHKO5AaW8dO1wJok6578TjUFPzZb2fE9N6lDEIvbrKS/MD+Z
O0xZR/5Qi5gDzZKJ3/hwbQMHlOw230eYJx0Oc37GXB5wC9x5cda+UIwYKw0X
G0PQKKwytOwBbqq1nPqd6UgnWjDR34mdVytyxcRdUkE+IQ1ApmYDUdtcb+cy
WWjJqniLeURH76cJ+lel2dSaiHV+kvqW8tUYB//XN+U1YjnBTL/Di2CtRfrC
GG5QGo5OOg6cSJCQyw8YOwqGG77RVUZw6ZStP3JJ+9RrvIvbFK5RtEMFsxfz
FZY2gwO/A9B4jaiN+4lSKIoDSTXmAC6YW/lS93Pbcl0lTXrlX4yIJRLZF+jJ
ZTEwnR5rEarMi2Q3QzpXL1LPKNjUatDraIqIEPjj6QsKKCmJxAZjYwGzLzGr
pzMaRUJeA4BUAFuZAHZFhRQ+m4rjvvIF6QNdlRyGoN9o4JI/Dogz1IyZg6vA
WgtlYQoXHej7LeQ+lVcFWa0yrQjV43a2Df5fUV8ij5c1NsNLH0FybD43YTuC
J4VgDvlB2U3ezqfbh9OsB6WKC2PfHCFA8Roqfy+4kCHipvbFSbAenu14LvHV
BgFVO+6tguiPXI1b/Zi+NjAbiFb/GUnFzySBFMO7xnCG2V9uNE2wn4SyvoU9
O0Y7EbEpL8H9ffhnygMIQjvw1RZ9/xRC9RtsedhhEAXBbHP5utkoWJcl2lne
FvYgRM1hnpOCbv5tNZn5XKJDM8G8slNUATqh1kRwcOIMyrbc1LGSNFkcgCNN
ub+jEp2lWbZ/7EaP68uuSa6XslVlmoRJQu4Fq78mtn1aAkZ6NXjXt3zenQph
n67LaVzTRrX+RBC8WCp2CfmdrB5tVzGB/KXFm4Vbm6JeuMucRjZc5T6vUvYY
cgcGcztmc0wCaEj3Z5hgHef57r5IpHT9r1wKmNsABQZXR0v7eDk/HdbSh+yJ
fuZ5qXpL19vtQg1MxoJJSH/+ujAOiPh2qagGe2L0fVKU+8WZmHySAAFmWXcm
b4/US0zZd8d6qG31lRxyG2hC7QxlDERiicJLcGtYsdNC1nXvR5nU2O1GuEvm
Bvw5qK0C1pbdGNLMTkdcPfmQKU+9gv1C4oCA79Khsi16NLN1GV24YImv0nYg
toH2AIubQGR08gvfnEcEt57l0U6tiOcVuFqUPkcPD9r7O0tKR+u2qxeMQJ2o
QernCQ6o7CoYIWs3Bq6z2Bw5PMLJ5qJRFUZJMAAPfRXAS0OotocsYEoQPkCZ
OcJqKB8YaLgOxc6s541y1DwQJEjGYzmlUCwnfPileR1qR4W0xW8DCi7IHz3v
1Jc94G5dSiYm5MRuN/GqPyguZkTkQ4LFm8zEOnPfaqzDsk/2bbXbwjHkXZ+I
vbc+rzTQ67otJGGVj//Sr7csmUHIWRr/ri0ZDWQTSmbaBmPxivFvE80JGY2Y
gymCiBSS1QUoF7EmE54uTGS3+NGAns9UZJQCHO+xtByuwx34F2X8aQinn6Kb
hCHs/Lkh9vCKGdVY5HSJxYOHJ+dt3O/LEYu6tI7IHWE7Mqmj2J+V7UL6nek3
ZnqawQEf6pwP/MbKC+Lhj+HemlUdXoVk/bageXMJKlskGcOAJq/hqPkWeCny
HOKLPNmeprihWJ/TAso1mNUU3+VChNV36KDWgFvVO1YXr5nCBZBZpaSR8meQ
vIl1kdvbnas7xG1luIRptP2rrQW9D5Wft8LyvLZa6gjbtB0Epc5dh6uFNPvk
z+RfdsfLxZrijZfv6+nxPtlbtlKde8U5pH1k+jIwiYak18FvCwPeHpp1zSul
Z/WirFYYsxjAVPGTiCeKnFXxPRcnTOdbFe8gUPOe9Jb6M1zG0vtkO4zpo3M4
JHz40ew/3Ii1Klij6gw3BDKj/NMDF/bGZ5k8JvadxJ0lDCGfYlrLEzyu4E/P
CNVGAyqNuqgJYgELbIKC7yiYufRKOHymwqt0RvQ4dW8dz9585I5Zk/td1SHJ
R6nF5C6JadRypVOW1rg+QldmlnHD/Fo1g4cEL6PT6uZNMkHibdS/5pB1HZGX
035KRzka+2Tk1/BxqQaKFnl++SA8dOxmABzeQLhVgwBU0DzpgbYvaOGgJeh4
VFSCSwEuw4cDCejQ0K6pBwrZhK6hFkQCcubRFr+eGUsmYWiPLs8LzddtZnjf
K7fMLMw1I5aRj697xwgTR0nIQoxvr7tLPAglBzpvPPtoeU7WzvSak7qw7x+q
7V+jD23YbVfe4mq7pd5a7Z5ntKhkFVwNzpRoo5XDstG3IklI6vXXRpSXwPQM
Wcv1rJT/qYwHVf993QomKwDa+41pvLBXHAi/m5mqJfM1CyRmBUQ81wKbohEe
yVXa6Den3Oye1RABc5bSDgMocXA8OVjjWyBX7JGmcknaI516C8q9Cwvf2Eim
Cb6uG0XFFUoDqZP+9f4PNVOw9NtcO3UyhQVbJnoR0b7a6QXX4LP70LhGKbaJ
UJ5Q4YTyFI15ykrzlxLGV2hOAM/OCYvRecTO80GcEIXWQhm5tv+lCdLJ1I36
j4nxNDCL8ectyX8aAdvNdnyx/kbtLl210sRDkOUQlabSR+HPIL+juasw740c
5FToj0m2zOknZ8lCnmm4VPFn439CaTB/uIQTIuufib8TeRWi2xPTis7d7bjV
xLQ8LjzeWpzXFmLdSg/18lh0giRTbn5ex/K4a9WtHsJw72KWtjDyQqq8TT8C
IodGPgfHqoGOe1TI3I75sNc+33bp4JoEY36T/+vK2iQzyUM+sS9Fkzy8v/gE
6WvRqcZILHGLYZXCDtYsRqh41lxw03G5BUG+znHxQxjCa3nwo/pTozNjl8Kn
BB3GZ+DPcwBWNKxSF6LZjgHlWxrnv31ZCtOp1E2KcTq/v3ZY2x6lvCmQm0q0
p9bPPoWQOECDdfs56DohVsP0NdTbS4LySeLoxWZM5mx8tzUL8kZrAjxag9ag
lJQuqUQFgtsJh33jODT2+eElsz2XNFD6SSI7QO87TehKVNQ7tZZBZwAskvfh
BL2giyXAsUfAsVIg9yl5vLBy5D7m8khATk3fDoXNQGsgLCkrRDGcudHNH2oQ
R2mRnaN3NhdiDlItWPhfSuBNTxQgCUb0nLAfrfL1E9XH9U3DcG2m0NfyrN9w
TB+/Opc4y+Trm2D3dfFfMPh0A9mUdxOcTn9t7WQQgUmXehkVZdaZ48SUODLo
EhKo+tmYcn23dfMjLDX5whj0zifHRtoXL1X9R+PyOabp8NwsPMzMoWDra6nN
bAylQk1HnvUuZF93ECBLzsIaM7a0bv6A0vohNIIdOVuaQ/nGPS5mrPANq55C
ULFg6qWZOJgtI46DzixKRX3SuSpbPM1bhT+ZrjupnYP5ErJFvGaTaMFpLOXY
4SsbLlTsnTvgzpLDNGZs2oTrZvjjS5XE5WsPmOanCQKowRIr6LOrjCD7S1CN
wpmhJj2GuYQLLEqOMzdcmYsF1x1/RmZx1rX3EBN+VSkUBvRPVYZ5vMdsH5pa
L1PIA+icp7lDqyq6qEC533C7MgSY5Oo5GZ/SvPv3WMC+d0Qi2Dy9B7FfoZS+
IxPl59FaIG4AhrvjSK1Xerq1ntezQlL2s34q0Yecjh3nIGym2DAhY272Vyau
5qGngn9s4bUk8qFHOyhEZkyH0uQE/73VjccyftIUlAm000CJUrpyamHrgHce
1pc36FHrXuAXIagFDzd8SlLV5QiGKlEWGZyW0nz/qLXywXhAlx1sPBATfnzG
U+dAkyB34Dzzgp7xiAli2oZoVZKAVErs01YgsbNjeW7KUOW7Cfso09aDPbiy
lXDKhjSm/7uMv8jYEkPPVhafi/JfvBJetT+bU5MjHHY/4FTzUAex2SvqUZvx
mtVodkMYdb9q486ymjqzqcY3w6XieJ7oxjxnE7XKLqBMpO1zwL1TEVdRoFzk
3pb284bXFwb6+sjKFg8BBp+d7yyG0O6pZEFZUhVbyraBck5lGKZZEyysZ9XN
o0fTIZJhA+5wfAhZiVS9wJvvEX3BFCRzYlY/9fPDgeYS2NSr9G9IFpJg6fY4
+LDcIdNC9s9qGM2fI7RrGZFC2Nk4oSj76TXVPiAcg6E2aoJ2NA9nBSbFdOkU
lWMUtt5Q31fLfwXfGmUHpMAD1LPBLUNdlJ3b+HKkJiBZici8hbTCvE3GZkhZ
7o+9cxM0ROOYGJtQNnly/r1UJ9dclEleBjJO4fH/q74O3BRy81jGCLNIZ/W2
gg98iM7zSRK0R3c7IEe8qk478CKqu1wuZT7MslD25WEpgGyz1NGVlumGyi6x
3eA2Lhx30l5Gapt87T2BwO0oR4EBL6AKA9i1GnXprzcMCJQReVf5yIsWKlUt
SwIMI4RUo3uopHh/ERhdw8Xolz3KeP3qLPvDHX2oqwIqwLwRi7Np0xwVOcqa
dVdFZZqYCPG7qYyFmMDa4DXkWLZJv/oLp+iYcjQAMhcfS7FYHwO7BNjSoxyX
V4O6zFuEZx256B3X7MkCEe5clP2vx8+1UkzpHlAe53MnX34rRsqt4wJQ51q3
rmmBTANUfYAfB9mSNx2Viq2368zi0OSIwaycWrJwZ9mJb6vDpmLDjJgnzTyr
tt93/e5WX8PaLFQqvAk1Zheg7JJ8L//AT/+yVQVzT6tT3Lrmb8Ny0aDjhV/A
vM8U8b5Lizq4SLp+1CaKNX+SrUHVX299YtgotNNPJ7x6b7GQZbk6wgrrROwH
gglhCWAsvQ2bFxn8pKdAwQiho44RfGHTfu9PBu4Wmds0q3zghxGKuR6rQLKP
pXb+Kk1wz6/eT0UKhq27xTadVtPFIqeEsJ58oNpd+2CeYB5hXf4ePCJCf9fU
V3Rp1zn2/OBw6/6mWkq66fFbV/ZH8400xON8C3QenJm81i2C/PSeI0qvn3sS
JXlxoT1o8D3FIauWaXtSePCSJj+A07ZTH4Y+D7SsfgkY32aa3SuN4hMXh5zG
sfkY+uONjltQVNZWsnEyTu4LQpUCyMN0KxjfJC63OSXxeAoTMUVEcUtf55R4
Sz2NZaDjRyBcAt6xXR68T/7QgumilX3R0qdSY7sdaVlQhnE/wpcnG21uETo9
+ktFN5QoLvrmL5ZGiMYjWFKgm9h2ZMYgCUv1AWSToo+Q3PBpHCdWfaX8H0H1
uOpuJAxE2pkAE+zygbTY39XSn6wEUSE7D59zYaOfHVYP7XIaMD7ZHiiigYUE
3zC2Qz0er19owQWCWCRqvrer0g4GoiZTyPkfHv5k4HNveWhRfTwyuhEfK9Ia
esD9Z9EiBSLLk1flrW1q1uXMgP+z11cA5FG5PThuYUIQaISdljOkItIXQ/Qq
k/583vt+GOLsvIp5obAJr8GefavMGomdn3G0AKhWvMmlf2ZVhk7Rr+OtQ1IF
saT4d9U56HjoKiEbK6KMivd9jN3ZoTqNKKpu6x6mQ9hf8PXCFK6LzjkSGDJq
sxG0KHQ5/bYVPBgBX0b2AjXmwxU2g74vdgwjb++lOPPZHPfvMLtLQ3KKoki4
s8/R7GkBC0uWpA5MDvCrtsVsvYwfIOF+UNFvHAXy3gGmsxf8xkqW9RsRGB/T
9NeM2KCOEagFTtDK058MxuYHWxLA3U1owG2/DNKHwjLO3YIaj8VjpyLSdMk7
Egi/I3WPOksGQqV8Z8i/A10d1ANQGO5BW0TByVRIO4j4Ntw8Y2mupC5n5QR1
ViPSHQ4B9mpdh0wJym4HsFYfQIr2XP7YEqiih1LWIa1TStYsjJaDkr+wz8Y5
XBNIHWcUuwUfkZpGbDyPxcOyEo+J7Ww3nsYQ3N/XT5tfm1zAPzRhvM9tlsos
6QcleF745Ft8OEvzPOsDjEjqBQaRY7vULFM4W0Goo7MG92ZvVk1J8eLOjXN+
XteW4WtTiJZAGeEYQ5wN5LuNvgzeTmQ4GwLJzTpMHYYabVaFVU2CVUP+Dq8B
LWn2gy3MBLo2CvZi3FDFW06AnjL7nG57gTbielU0BsNKzmHyWQ9MytxHWSw5
+y+qbA2fSvl8cdauzG2UZU2pKoffG9/U9769rRuadoqvW8eeXFZo5jCHAdyM
/rjBtrH/2KnmelHpGhDeWcwI9cGQQIMWmDYME6Wvdcc5yyRkaLNskp1vk3MW
fEplrLiow9mI9kB/9nlDiIqTN7zj7WsM1I7fYlCqx2vGfNBTOSNcqK8xXrOy
Mz+5La4M5gzN1biTcg6UG349OdHq9WqAVmkWuSpxQlKheZAlfWk12/s6gd1z
lRQG+woQhb14xOm4h/x+4+rsJdjdeuA/SBZOzg53B2sCbKUePrXSmkBx5zfN
e4i4DhieXfjv0rno9uIbKpStAsVRrBJjlwI06BwXFt5eUo+r3g6MYJDrCxOX
uflPmJ9uPEhbkpoRYywMs1rCe70nEJneEGFSRBNJtaGlE/VsRY1KCbVyb7HF
Tx0m7AFsV8+u2t+toSiqMrOoH1xxMN//5qrz87r6oiAw8f6VIdSDUEijegc0
EMhoFmvTdfZRlWNBV91u2eEmMkXzVee2/E1otvceXu7oqZXBE0rUsXYMneSy
eLEAQoXCU4pPkGZVC54LkjgXDcvs1sWb1I6kwe6cJyU857+ZoOa3WjmPidwt
0CEvKIUtyD9RSRfvco3EpQD/65qH28zK1vA7QcjgLFvyYduhF/ldn2yFfM0C
vx/+35a33ThW9evphv/a4xEDLhtsMNtRyFJSE2rimUdJ1qL3iGioiO97PIbE
hZrzvrbLg5cFy7Gv7NiC3peBGzGNfjx+e+32PgOx0edG8mv4WYSk8yZEjav1
kSjD0pon9FZ41GDaOjQJ+Mv+UC5RefnUDaBhjLxs9AVWBCf8GuoplpkL2AbZ
MeCrLIqtrbq/qZydArtzKVs+DiSTv5vXI/55Kfmj+OfRPiVBpCMSJ0HX46nR
HfkRi2hbpDthfYSWkuyv2P3KpNKifaGysZ3xRUhc5SGYh0r9W1kbFrNeYxAy
jiV8kg9aHvuPVaflN6PAQJ/qP54WwfkKz+73rn8o0InqiBDtaJtQCJNXPDCP
sAJHtvzem8zONIcxrjcLcxnYbHz+KQ1hCYcQRK4Pfx7LxGQqGUmzJk1cwTyt
iOphfAgLIy5aN0X7wkwDlbHJiPVcB35ujPeMHzPVUdVPNcrBdM+vMINK99bc
qf2yXgPD1JAn0qqSA6EDoYr69goqXagsc/XHQexdFCLEzXqjKpjiu3e1Hl5J
/EBKgCVbLxvlr3bWoPYLvg5UwYvQ3UM7M9cTY4ESj/dDO7f7AM0LB/Pn20Sf
tsc1ieYbLMdm2VvUWv1o78KfvHcmHvEdT7nrp8OJqC0RPG17NVIvWt75hkDL
KM/sebz1JFjjVzPd3yVxM1VpqJhVy1yLHeFsahnZAVudLVAGrF/3KCc2iz1D
qjZoeWkfjGOd5gvfbXj8sd9Bv3gXdDyoNWqFKfBc9fVYqsBfvigLVrMOJBNX
yifWL5ca7UNlEf7cBha5oY/4XwxvMRVJjPrSlW+YRiSwnoNXPbOOTwHUkAEZ
oMrL12c40rzjBpfHk6o8mbrQjRE9oWYoP4seu6AKc5VrZ9EY81FzeclpUomI
IR2722PRMjFZvUZg76N2CGhLYaNvxPeaEZdNWCR5EqykgSFs2J2ejRW7R4kI
j0uPUfA0YpdQvv40svL6fHEfT8P6MRhzMCMtSXtfejCPaYxlEANZoOERXY+Y
VTNUnBlKtInx5As4CO/lWWlAGRrb76lqgEaLxY4VM8J87yMHG4aD7+pjhEKG
xYkrk5Kq9XI3CsJ/Wy4Rrb8AWNEPq3vbQP0AbMeKEmxOGVkXTl+fpJAgqic1
4KjW7nBglV4eObbqvBMpR2SKQUm0XMJcq8hPrwvnWu0J/xiwasXz5Upe1vT2
A8gh8oQMxWuw/5cyl6e5G73jkH+4YxVAGxHdhBMYiaDB0EoRuGI8zOiB9rsO
enXK5xNkmVwaKqnOrB79rO5WyjXxF+LGaYENDpz2DzwUDDoYKaEG1NHpIckO
T2QFI/ixmLZ7rdEzScZ6yc9iby48ITxXhONIFM3Wnl2W8yhKgrSVQYS2cspA
K15NAQJw1/G0PMyvE17eEHl363VnCCO8fow/V7wBSA/xqjdMSPd9FPz7/wVc
zWaEJakQNTR9rgYQTzFm1cHvZzkb2ETanSdpoA3TH88UvBEWnuZirg85nfNa
yXoGfWv4s11hSeYjKIaYnJLhmDcsWV9mmp7TXenCQDE49eJbMqXQrbFRkXmf
w0QUV5djY4fT1x7/19R0Qp8i/7wit3gjgmnRYA0O8vj5RKyTTtTuNExV2x4l
e9eLAXGKCQRhAW5V2u4Ax6mUAd3kvDepPfpCbN5xWeEG2gNYEQHSnHJKFq3S
F6Kj7i9+46l1fgm2N7J/YKrvHOmLqS8jeDcpDbTn7p8ET7ME8LFOwmQfgLqF
pvdpB7OyuM7lBU1TpA/M9xGXu3DbsZgCYYtaUC1UDpXv4s9wkTN2NjD0A9xM
NYsPpnUguISsgJcY5DpFamzL8WrTGQDbpnC/9oUVzowoY9rDmhTGLeaZJG7k
9wKteVy7WivrsHbFMYUZXVhqOgtvgSYEUcZkT/0dZ+ZCpAxRPOhQYCkCsWL/
MuHiwtiHanNVV/NwRaw+D7K5rq/lxFHwnX+pbuDF52vy6Tk2TKbbkPQmqOZb
RY3M86frfihxpp3fTLzPxPe1PZVEgN0vHIrGJ9mkKO/mv+Ba0uEgZ0S++Wr1
XnDNf46LnzO705ODARznsrmrcQQixFifVUitJNALlcQUncO9vHC/7tBPTiwF
3C0kLel71ylmNMvQnpmJgx76HiFZaY/WJX4c/ldWFYYJSU1LQa907i27yM3K
vqFELCdfpEzT3ndE3ENBAlsc68DN60SZo7JCYZPTRmTwxqspzO2a0UuAYQt0
thLrWhX6eDDHd5xMtQw+aZIWFT/RTL4rY2/x/K1tYNgxUiTxmPaqdS6dTQx5
PAMHoFsmbgAXJAG4UuD7drdpoNetJY6om19BV+pA2EVJxkg8WKQHNOX/ns4q
whxg6NydG7U4SQ4bn+bjVWQ9KaM11zJMIDzauL6sDPZ+pLZNqnyj89D7n+b5
M/2F1FZOGmH80WIGdFUg3EWfVbCJ0m11NTHDrLyrokxAjEnLPiKVpTUyRfQc
3EDFBhIc92r3KbVr3cbB0HvPzJi99WjPEsm3yUoKYjFS2rGZrxY3wx2mtmfJ
i3yYRG3CqUldfw2n25m5X979Gwh3F242i5qhpGTjFsw+DUlfIfyqLgUjXufw
dtbVyCU6zmU1EuqtCIT4kBBmlXNH/I3IWLfQK5Ej08S36ImudpiqODghqXwS
mzRwf/U+mMOoZCMGp+EbAzINASjB4r/BSMfU2uc8WYMn8YHUTEuNbRxmEm3y
P1izwwb9MfO3WGh952meLnyEGkYw8jVM7vNYXZXGHw4rk6QMFtRrLacerwEy
AWWf74qg70JE8ejDR2YbPcTwMpYFon5efegxFKR03Y5umBJlf4SoZo7eDbOS
K6tLD8R4Db/2KjxMuNFR4q85Y+V72zfaU4tyAswK+ihA4iw06JkqCxe6L11h
qr+F6DX4ovTV6TKfP2ceUd68RHeedh6Y7R8bzUVKSgBmSqdl5et0wWTq4dVo
ryMJEt+0zC9D1RvCWHgk1pQgohEtNYzzo4mNPEc5Zf2qwB79dSLI4fctQjFs
Jll5j3kZUgHjfNp6Om3r+F/daX1zyJNMOFD+XahWCGW5stN/bV8d1yD67ycs
7Wk+y6V6drHHnfE0LQ//yvZNNq2liOckxFz1EYLGodPde69cJsRkZCaHfSK3
gztWfBkf6HrofxTiM6aIaINWKmi8MfkaVqbmLAcFA2jBm0U2Kjz+eM0NnhiO
2gSRRj8Vsp8c6Q2v9caPiteKS+aSMBszGn7gRUGhMgZTc96YOXUZL5z6ZOjE
IXLpoHiXkdkWjScq4ihclU1WpQh2rD+65q6zhFm/EyWzqUij1Y8OBskct4hX
PtnjCFSXL8y4aFhBJk6hCdCiEzZee0YVNGFsGiU3iF26aRLX29ze8bxv+B3M
F664eU0PXFGT6FN10f1Dba1ao17noONan/TAUz7WwEDuI+kaij2KrgIMXLw+
hcjRqGzvS4VJgeXHc5BPnja1eJaHe2435ttzOIHhgUPt+QWuWCLLnxHS3CZH
8OBaYrnyFDetL1zWBejjg2nXS+FevdnxFqTOvzOSn/U9dZo6Deebk4iZR37o
5CipZdlAGskesgV5mLIEQhfh5/WLX1tjZkLQGn5g4+Bi13dNfuTZBLdi/mXT
uOaylqh3+8MvSNmN6w4e0yOj/MTeXr0pRjKG4U/KxV7zR8fqOS0QdBnnul5O
WYYoCkaGdZD6otSjCMRWdQyHmnO3mOVK4SgZ/iTvpPGsOwFWrsqt1Kps/AIF
70sQpHo8Msg8ePr36/MiqqVB7+SmkO+I0P5tg0Qc2H6+zdd8hLtJKlXzc7z2
3ZWwjK726WaqGecyLV9vSv28tTOiOiNPNmBBPdfo+/qdbx1HZcFgWmO3cYCX
k2f5kK/AF1eJCmYUATYRKSSs5Fl3WimN4vWTGxP8PGjwtON3vexfKoOYywnf
1Tas5ytCwfzulW9K+f+MetfJ8kSZeKFy/VHYwMAFB9Ah4a7e4CaPWZ/MtG2d
NKThdGR5eFFt6aJX+t+uou0O+740ncbOKl3S2AW9LFUT2V9PHTY9NqBq9MM5
Y6mPmFZLU2ivrZXchlPZ9z38nK0cXwHhuLRczBVYDg2IMkUHrQ6fjZivtSaX
kOHIxvuDLg8z6NfxL4UrB9JDDoVMe2jUz7B9XtKoLLllqY2euzJ7jBj96knM
s/8aDOiVzn9Bq777dtgbG8jq+qEavswMuQspBV5E/64t8p8Yi71MgZRhl2bT
Xu7gzt8samA9/VoiuW+eTuPbxdoHVJImaWSMBvekvx+9YleNyyVEgg/APTOK
2pXEp1APv1bdS4pOZfN8NgEZiOXWrPRtnwpomddphhI4DVYh9DIOgSr9HV2S
2WGMk1TR7EzeJ7HbeIImfpNR8hjViSRu9l/3aY/OCothCckUc2IUXc0oEPpD
WgPiK1QbIGoDs457JsIF55o/tsolT2vdW8HrudeW2w4utQ6nseqSl0KNVm37
XA8sRASCVt69TvREsDZ5UULbqz95wMQoU2VHBxDmW83S1jPzLFxII4ZZQLL/
ryxZxMVfSUuthgdOu1JWm1Ds1/Gtw/XIFjQLT+s+QB9x028aRtpfmzZNzVOF
Q/g0gwV7Ui6NXHPksDV4KeGmH92wBJeKLXDlpELnvsGE+ky+uTNay+HGCYv2
gStxvg+5rzog7TQN1Jev6wq12TMx7G1J36mS97f+i7IeUAdA2wc0s0NpBBiO
96+JV1/pGjB/hQnGGpNU8j1a3SVNxA/gWCeVztgIF0D+aVQ8aY4Cc0crspOV
BXrv8LeXR4weqmYpBwjUpet/D3q30i5+Iht2s31P5Yt8YPPusmxBPfAPjuuo
hrmxdIOpGMGF23Ig31M0aa/jhPmrAuK77TomIQTgM57k4Cde9DIGSH39Zd2x
+RBZzU9zTLR+vWjCoupC0/IEjJheBEpPx/UqLYOuOj8c7lPGdtJT5fye7b+l
hh/qTteJUtY1K2yd4Ej6RCvq+Rau/InWScxCnr2cflqFSzBtlBsJ4XkDRY9R
oFSzUvF/TTxkJv+wSECcA404wmOh6FQbeoTH1JoNPgLB0dRp8AjGKJd0n/2R
INgkWGfkpzhkS3pFq8RXUNvAC0YSGr1GOWcPGUyzdS666xrwjTtaiHnhxyOm
mbPIin8xjc3Xp2z1DxVlqK/i+sbdPk7G0gQ6t+LhA5k7qMU5fUoZXVEdSIJ8
anI3j9wgPIyn9S/2IWQVx2K5PkT3Lv4mHFhiemUY/NJpbI3SS6oPcGVyUynN
cAYqg3MpeJq3FWp16j+5KLBNdXJWMMH1z45blW0MYMzLqEwOF1sc3biKvZWa
UddSiiY549ahZkMAHtIh0RtBkyCfIhIN8IfUwPRiGfzoju4WcG0CKRIhpSQZ
5J5uYjz8NJDQB6P4fV3PCI0YL8gHKGYOA2Nsj4MN62Wop0zYJGQq2Ar0MnU5
7RR5Y8hhMcikQdk67Xy/EXgzHL9qnye55cwfoC7qKM+pQHnqz5NcaWcgEXSu
c+KgCj8BFpqTob00SMlCcwBSC+GX+oh2bW8PIQGroZLsBEG2GkgQe8mfIM7k
V0McGD577EM/+bwD8h6GK9LEGGP3VbToWswtdHACIATv4MyRVTZHzFHK4muL
k77ZDWTHNu0G0Yzwb1h32QGm/Iw3fzO2gLRG26904bhNBjZsk5RxxJKWqYrc
QmUAND2ZquGTwP4BPnCogCLKmyXkcJnqyyhN0W4cvuFi4YUlGrTmJm5HMRhP
Ouwtl+un8BStC4Ybat2RcwL3GY0u1kuqBo+VUUvjn7M1oXvQqQu/f/AL4SCX
C0UPfDh9RyXQvysnx04hE0ZRXRj9pXiTTBgneV0MvUVVnZcNNV/hIHeb/qco
OXT78plS+u+jBVDjesDRleI7LEVii/kdX0B2iH4eFQbDDsVsWkNdjvEjf2a8
DFrSi41M3AcBdUaUpIpKRHUFjRUeUTsQ+j2pIO8cnwBk9kkH3t0Z0lRmqOCq
+wEbfyWTVrLBFxrper/PI2b2HwjoTbh2qkLWxOfDRoxfGAwiFCXkfseJNQ6V
wFaMvikvJcn1SN048/2VYDJHi33a88K8ON4YqnJFi9JD/UYE2unwf/4emPH2
UmgNmiBUgUqKOdIEdYBfmb7Bq3UziTDZ/jRYfMDZAcpV+ra19Q6EDvh0aexP
zGwJRRKwG+dVHXur6wB4xGkM+kAHoTb93tPJ70CuR6x7jPmt12RUGLq8xzEJ
CLXBe2PqojBKbInc1dSJ9qfDjv1uLQDXviHNH+Qe2zASct+R647Sw6FMOojy
xUPJN/KaqMMGpXRC9smmbiwmJ5LiKw6iVMfeezkHsZ8PkX4lABc/AcsZt2Mw
IjWynHrGnyidFBdNtm1ZFem21nuHpThHGC1/jRudBMYT8d6hGU0OAC7ILawb
JH9i43n1e55jX2CFfIUr9YLVEWUiP7uOwTgRcxfRidqZMD+Uz1IYsofGERCD
C+81ZFyWotxzQfJUIl/k7x9puzXriud4T394uQ3mKutlXF8ycf9Ymw5nmdF1
eGyf60yHCtAhkrLcKTqGokDbxJCTjLoRvgoSrBUknLlX62PD6ek2WQrUqkSs
TGmGjP1kqY08DyEvBYVGTY0AZOTuTfq8Md232WGM98PO05MhTYdioMFWAK9K
k0rfZjKNVbKdA8k58ahL+T0/6o7Vnn7PZCq81Zueo32reYFkyzwwBGdM54L3
YUQW4bSusfzu66cR23jJeGnw503S1RpF16n/ESctF+wg20PFzbspnHB0iRhb
cdAT/tOCVG7sWWicGjliNen+pWc0oMoeT/e3oqiAuf20i0Dw7PX5Pr1LvTwv
S8cvWMPQdiCg5Jein7yJgxsscujXupycZ5zkkgl+UtQVDYAVJWtWwru0M4Q7
C+6FA8bt3GwsCXlZhlBzV29GlrQhL3wooebO4259k9c6yotO6g5rMrIogS2w
n74Cy1w8nAqlGWyIJa5n3VBdmwY1YVkfD96vw/yMD8VDOCdImD/PCxnLkTOk
Gad2Cv80n1JQa2VqjQboga5QrRgYgIK0BcFO1lZuT3Qdd9Cugx+hBu8D+zUb
5FqP0FiIZ27SNg1pQeEBXc46Xo24c5cFHzGvpHKBbu8LBiL/DKOITyZXPLIk
AxtLF1zYIQc3Ybdk+RrvPyO/H6Qbamh9dDoSNu7dmEqZ1vumY6WKjMsyE6Zt
zNXYrB26pfDHhez4FOTkjXrRlTN9zhHZqs+HgGGf0ve3DtPJT2neowS/lEsI
cIyPbT9yfsM2TgSC7cLFmSXux4x5Mtp87lKao8L6KhtDXefjIfAPILKit9ev
tZUoHq4hCXfKdjCLHRuItGJeIXBGQ4rDO8p8i+BkA2IIyODns2kYOCRCqjkx
iv8eDoFfcOziOu/eROABr5fn/r9k6Ho6iZz2Wt7gore04qApHxcU+uN7swUc
fsfMWGLZlWzdN5bn/4IsjSC2Gs9FYOe/2ioQO+unmTQjJBN92lnj/B7MRXWm
HpOsxOyN3cKD532mSxG+RhefhpDzQvcP5T9AoQrNIoqoK0CzU/5K0meaMAmM
rHXdek3J4Wl5u7v97NS3CGZmGW1GwqhdJKkrnoMiLrKnz+B4DCothS70d3AW
+nN1lE0Onwm/KCOAFCwe2mvxkNqNpMicw57ME7xys6yn/6cPMtu6lwxh6dUx
MDEYdykSVV+gYpTsPjWS/9wDnehzrdBDAjhzeWebi8fGbE/f+XS3yLLGxfNk
A5ynO73zgaUTmSiwmvwCbYVfo9tVWCRCoB3+7JOzj76Uchob/6nI53NbG9RO
RHm6xe7/wLE39GrvX5Tnq2OBTQNMz5ngt1pWv7/sWrDejJ0vBhFk+5A4U3az
12wtoFclJA+JBBqt87xY4BVJ+dO6GfYV24OUWRD87vENj+7DyxN1UQ5DQ8hi
5IJ+f4/eP5tmGG/cxdOMOZN/vceFZUeXXZvavEyHENSBbcmCoYsN4oNTGwUI
Ag5vKEJB/z4J4wjxMIEvbtjvVvKAgASm5/8pKttMDWIfVAwcuYzV9y+NNO3v
kdn620+ypV8jT6FE40jmfZkDDA3NCqq0FsXndcdvOMf3CkS6gBGaApvuYvJu
vo3X7iwrwPlolVpi1LHqk5zUBHG446NK2HxefzSCZeTBLN53NcIYLD7Iw0X4
2J6Y2Ou9lC8f0Wkq41IOrAfknbuvdzFQt7cJac962E0QjLeUuOFOj7DVmBfx
Rxpvv6Pi3wIwIBljZPuCdOeeVY8TZtLtydS/GwG3S7FAsoaFnkIwAfjT0GEF
FGZgOdSppPE4Wcbiy4YklzuxK7dcjjQdmNNpG/2YbkZTwkfCnKeFRx5XieRX
rjn7o0E/0aFmR3+pTPPLpwgxqBFWIs3EW07XM4gUVBAqBe3nI9Vks9MXUmjj
FdB6el0D6ElOdbkPMFaoGJCDXtUe8cnQEy3cPolrm+hYdAdVpJWMlr2lkAei
v9Rx3mEwiHUDVAhOyYSNqnyzuYKawKlMfJXaz5QgWquNKvzlhPHua220B7fF
MjjipzUM/Yfr6fwj2czaeLuVe3aYDkdqBv2TL6vefi06TKO3pelXsIRB25xU
J4iREuh8AelZXVJgVzZxeTevcsHAnIlZnm0eCsFF7Rd7RxXN64FmrDia5dLq
MygfqBM6hCHk8OLP1mFa2DXeummEuMCFyCGKxA6tkE29YMCzUZlhpcsDqU4f
fOgbGnodmz81bN9Tm7FCcM8br3EVcStt066RAs3zEEyV8rxxc9jkIz13r3Be
8gC4tSYN2BsDGTHja6LUJna7L6bylm+gJdeCz4L+nFF7YmBSydF70Dz8/k6Z
3fXJXSBISnLwGiG2ibVRN/aFqO9UVcgGm0vx76+ai/d/wZT7+njAYgoQC0za
47ak9BGbGPSAvdlmf9MvVEyiwk+ULYk27GfHnstXIy35xpSdbGFev3bJ5HZt
BLDkVW4DGHqDwB8bmclM/2OPQ/QS5igAUDGILswkMtV28y+omkUrISN9aKwB
Ko75xgfqGC9jXsdMb5GrAYj0GvhL2AJh6KtJ3FUWkoDmfOJLDLDy5COxGWS+
6hnn56Y3+BKaG4vqp+BmiJVE7ED7V5e5YJ/uIK9zU2xVVETk6nh5mrQ1Op2p
S1cEkmUq967alGCrnyiZE6hZI7yXoPERggMKCzFozpue/1IqGzkf4tw0IQCO
q6v237qz/kPEnSA23phFwjf6sAA5fWO2J8jb+vboC9SEENDnBYYSQNfEX4J3
K8iVG9euSIyTbjj+J1lz59/y7I3nLUvgJbkb4v99Q0Ha8C8zl0Ex9myaRyw+
7w/G3NBz/w2ij4X/TBCjM5AHDhZGQaJ6mOArCzDDP3z9GK6tFR16oPo45GHR
uZ4iCW9XzYGVHdcHyaLdELaOHeFFBvbiklPrBhHHcDKwsnM12mVhzc3SSWXm
aZTrDbgGV7m8PL6lyquSyJXKbmychbakk/0PVKbs6LvD2GRBRxSw+nV2fEkN
IYT2xiNkcKiXwKZYl8qypTDg/LWZbGTuv4W53CQJNwUpJyLl5Z84yKIpivkQ
bGQhWDY6eWB23U4LLPtKylpGl4XBzZ1kxOZhbEIde16myTe5eRJCw77uWZga
LCeDEV9GO9sMWsS7KIaC9G9Npmc8UvfoNKHKOID1w4XkpqGdVm6vV35T28bg
qfocUd1RIuRpk4irCcaWE/HMMrF06oBzvl48lfj8zLF7e9v9pvFI8Jgh1Fq5
LmV5+7+32COzTTzA3FRuKOjnKZiJazyJf8jcC+NQtWRLqKRm7ZbcBQl5EzIA
1oEHK3s5CZ1yvrFV3dv/60q4KZHkB7KWDiCc7wF3YxjJgcircZHruLtPsTpf
kvEOKlBI1Q4X8vvD+46OgLEp8dXY0pPTXHnCKsB1NN0mbE1pulVXRLJfCM4r
fCAyQiU8g4cq56tWJngp0Rb89n4GNqqlJh5qKKaw8tbJ92zIJyoIsK6qepy8
NhxP/64Bjah5Y1qbyOuBe3xhzqw7yWqiQr7sBIidL5IeIn9//xpEj6nXGEUD
r7qNRXA1kOKdWbtOwduqau6G1q1lIyl5I7mC5lPdug7tb1Q3SPdciZzNVvDo
bchNEDRRaK0etj0NTPWqYbOegWl7NQLJSoYLs4O4rIFwHjYPjR6Js3Flbt2F
PbkMrmv21UzZ+dhgLWOuDoWFDYsa9igRz2UZp+oiUP39MPF6Ad6dyOgGf77k
XlVyJUKj2V27oxpfmbxuPHV5HySAnfjCXOuOMugtXixhWWzJKHP31zd5Zt05
zMkf5DjYoQu7eOB9FiYPkm+XBWZjBRdt0XSgcsr3uIjWInc5sp4p98jrcCbM
k5RHSGme7C7SfGcz/kWc+K82UL1lfUsuvMiM8MPJgyKnoE1zGjSY+joMpqig
MSnLSeUnxGJsZHU838e4xrMgK9syBId8jdSv3TkHwQfT9IlAaxFO6BftmPO3
LXM70tozXeSV1SXsyfm6kNaWnRouvtT98SYA+K/yPGIZdRyBzFb0LSMQ6x/O
vYa5NEc3IYWHfjBcRtJafbi5AuMkdv1tZYL0XCQDMhfh3y1GB9TgexzhB1Pg
ZgJWQv4kWS+4GqkdEdYDbV5Zcpn2mmzohXL0PTKW6v6C+uHackjn4KgLAEDy
XouWmFQ2xndrIuevqygDA4CRdOOL5iziSz3XoFvQn+XeLCCpJopk7HeWzDRx
AcGHq39k17Dl/86EoIJnLDjIxxFgwzGwXGtndrFwmNw8RfoXBZksUGLlVf91
OwmX/EjBCjLotyBl5qKOQFSna+byhFKbsHyggqW1mj0LzcvLxhAyqBKXp/H5
VrDN4J8Ckyus0whh4qWsCr3jOAP/JtmOrlCmC0u5S776NTEJx2cCyTDvAiQ1
Vgl40RK2E0KqJjR2pnvRz9A+ipujxnA0uOpEl3oxFhMorv/wC8eLtU8l5Lff
PqudbQoB+WjTng635uwIN+fstRlOtH1s58vtt2N+U8QjNef2Hi7tsY5JRM/D
0qEPqq+k395iP5dhNHkQayWybT3/rEs2LhV6acSIJ9quaS96Z9h46ujPFS+M
WFoUOeATM3vgDFAez7SgCijRmR8g5Rkmn57PCICQfjhe0vOW+RC5CX2hsBuj
14h50YMhEHM6PitU1bpN069JpmbqiLSW/fd3ZuAifFsKSFgGQOa1ZHG29NrL
008CcdMgeoElr9U9El6pg2X/okgDnTNxII0uVQkVNVJtbODJfMOBZ+elevmT
smTjf2rd7VQma1aOBqi0Qw8FXWGBFDzR58CuXnA0gU7VfZ3aKhurTWebWr+U
szsG8QW6E3SJBEfgXxRfCHCGfR9EELq8gNDub6TX/p/rR9TxaIOGlZ3d/b5r
iO//1B99dZiwjozBrnKqv3UNK9BlrZG5narEzJDRtgrxyhpxn65RLcjScRI6
rHa5bFUrlANTZCi1QLr9wvsvyZ6W9S32CBoB3jThrgKzw6N1Ww6/fI/kMxmm
RTG/NJ7dBxOY5yUZ6k6gdX4CcEu7wSDiavlDEJm7v9J7JZ0FfFivtnYtMqkl
lZVbsFxHO4zhrU5BqlwWLFbzGhnMmpx3Pt2zHi0+sYQqrFx9xLLh9pQd/zW9
llUtykZ3Lbd2T+JKKM5YATP+2Iu/3OuuD5GVm1dxme6eJNusy6kox3FjGKJE
H7ozmvnkWF334z9O5r9tSYBQ0mB346+SQgxE3VxeejBJ7C06eeRFmWHg4/uh
nTmwM2O/Bqmw5WIj5GPt/tuX0Hl6OBnfEVMJqof0PX5BfeCAdsYs1Z/qXYFE
gfyp+VJ+6EEsY4q55v1ib3XHNcI9sCyutj4N/gggK3A8DHYcdRVSWFHhV8af
3ZpwV6Ft6JgoCnzzq2b3Lzs1K+osbhP9RZkLoNU4aM0W7IVs5zMeL2VmZ80J
9cjmmy49Dch5nBu/B1LTY4ckYT1Tc+a1N9XoI9gVuOuuCufoleyukAJ4hdzY
zQXLV6DNGR3YVb2oIv1ka7GSBEY8pRd/GENjcwOeOUpDGfGcEs/9MeFL55+k
Y7mx1lLcQMhR+x7/fsVU2QdxRzoapo+YMlyhyXLzu6l3sdNFEzRypTQ9EqA0
YA2bQa9iiziPMTbPFT1/HrUM5Uko/ScnPK1L6MKnkRDwZspEu2niHu6u1tWc
kEBqTcCgs+/qvpM2W0ZtFfSThj3gTS3ehV4cUpYVD/ae2ldMuJBoBdsvA6Wz
U6yc4bTyDNsyDml+v97J1k8B9K/kbjv/bY4pEv3kZm4gddTaPcJ/CZhIQZ9A
9XKn/fB4gtnG0kDHVYkHCLrhsZQqK9HhrpYPTd+2JlucoWF2rkJoKFq1AHIZ
UkVIj5CAe/DIZGjpyGa3GDwYJus+1C0/PGc+sJXWluPnQyaRqEiJvC8YJTF2
BDuAt5Dn48kjwDuis7lyCQfH43S0w69oXOn49k7UL4iTCZf0Zcr83TQxVCaJ
opO2H2wnszppdtXq/B/SQxWM/ezh6XFOk2WpgjgOftzgK6qowEg53zmlOp11
BoVZbhEcxYVp6GFipHecKT1kT3tX7B/ycTIG80F4zfQ7UZFA/JupBUasYXBz
BYA3Zg5FwsLMmXd5Cgv9cPoBx34jV/gVJvKoNzDk+GxFwjyGSfPsii1S+/Fz
CfYdKJJ8/6j0SDfJubNAALIJKYwQy9rkorCjyA4zCWVXKETACZJ5qe4oN6C/
jl5yqU0Pfq4CMNHy0lXAHlnlkPYYoTXKigVu3rqsbv3Zh0B2+Vis59jMY2YQ
LcRAcn7wy6yzeqecsjjQ1nNwV/KK7zeZlkGLZ3jrncyPBvG0ibSZExY/FVsO
pRmppV18X/BUTLajzTJMPElwpj0k2h/yTpx9CGgf/fUBuoz75Osh+GX1Mr5F
CKkjrYF6cxAIG/iPe+OocoiiqRRTuxP95aSF5Jzdy4wZAcs7uiYc4R92JGIc
JbntdlJvMon+BxkFCv9vKzSEoJBYP1badeZOLXvGvbdYVxTsyGChKwuZ4ziS
mHkbhceduTxKMwwZo5/IwchfjWdmP1Ad9K3KsrQtridcpphq876tNJa87pEl
2jhL4JUoeTbQhJnUo0VXwlB8EbL6LyzoFqfWsunv7sMtUH6jLF54VtuUDgxw
SDSvbBIbvvmdnR8NVJgKTbAANItlt3mK9laAe9wFGVKpL3quXQ/DggeSRpob
SiVXqhiBOS8pWCOXq3XHDoPVMMVTuqrCeii+59fuX4BU8hviNQj5Q7/Lxtfr
aGrzXlACujTABQQ5ebpPLjR0nCLrW4fzBoAe49+py4f9ag64R8QVXKovBPHr
RQ1XSBFYMMO6RRQ5L1ZcvD9atIz/2h9zgVui+PKJZUa2g3JJJXpVGqs2vUpi
hc0yu2aV2wpancMr9LiWJ4qKxS0oK6uuiLf3xBbT0bYr5mKgGTAU2FXFNdzv
a4dZ6sNh9OJhbODq1SqBboYTK/lgmba16dQlPa/YcrVPQ3Gvr2qFhppmj/qi
sBNnrOSbF31Tpj+KLPXuouLPqWhkM9ye7F8VQIpsDmDPJNgQisP2pskD03a4
mMbnkNfvb/5C1VIfNfK6k2E+R1YXOUjpCeS4Ww+coeV3X1B7lkTJKCFfvHlF
ME6wYe6neWimocmM+bWfGa6L+CcD/avTJNOtNBs90CqeTWWMmdA8rNXw4XH1
rWr0EMUiCbehDIe4scTmnZ85bJJ+oie9vYVeNId9WOD/58MXVFV/mccdDJ/6
IbZnkLfDl0/RPEezEoTcK/74QI+kWWC6Gc/To9yOeHERgfA3QVsswBm/n3rT
8J4x5tttS4sIIZ0lOMPTE78d7AZ0nI9/+yMZSgTBlT4tEBNw/Jxr3vFaWNql
uPdwRj/JeOG6dGRtmc/h6wcKoGBnQ7kAJe5KG6R7bWDHoTcEgdShoBBIJXLH
nUM9/XbHl+5jL5kr4fkY4FwPAxF/fShW2dpxp/ZW6GTnPR1C0K6RRZC5an3l
cO6woQqtoITpfiV3UDfnxYePC6dwdFErMELspKIqwe3fstM8pErhFg41dcgl
PaGtWKNrprh8gRFMKiKhaVY2GxLjwI4W07mUIb4uldlD/Khy1c4OxvxroL/h
DW38/IxgrdSlMOqrQOsXP4HmHVo+HvJMkzpyQQEj7uJxutYMSlsVCgc2M7rH
jTkH6ZGhfGLRuF8f4uO5mNxSQdMr9SvbwP2uKX5FWBx4iIYba0xO+5nS3Z1J
y4g3qbyj8dU178rLIKuho+evWNuK/GgeHXmtoNf1xKI/rHNhMCfxX2hBzFFo
dX1tBXJ/HpuymASJUvqLoySDrgblwULIpf4D4IkV/tK1+qbQM9hvD2UNjW/3
aV06ByIBNVzdG/XQIBo0g7VnppTpz5NAAt8wOqLPkhNLdYSeuUzU4SvlOirn
MDu3eUxLdi32mWMoLiCx3sXTwVh5jDImoNICD8H1ny8BHakAZaYFzVnL0xuw
bvsXnyTkcsbt6QKEdGJGi/WFVPxwDnA4datLIHseGpVTOyA7mG9YOt0xOrF8
FYIECAzYlwk1LJkRZ7AE+8A9puSRm6YSDG3KcMmZjjUOkiZYJ7cWzfL7CyvE
+3a//r3OuwI6EtTYvc+r+yWbaQ2NnaxbzbraauBeYO1oRoacZVN5xORvg0qT
JtmLo37Qcx/Qayj7YDy/3DMOrYakEBUfB3JXHvzhrlPTonKnXJiYKHU1/xM6
P6REg5GniT6ers6BsJ+SUC7sAnz0yqAgHKHVVK6EZiBLk45j5tjKQBZt9Key
tEPQYEl3X1U1ShvHeNnIai0McVIqqg6iWPWB5iTiivx+hwDTiPo5ack6gIr6
1HzSZm4QmdBZVVGqgHSGlXTf6mbk6UspXRMsO1+OfwIWWAeEp9/yZPyK540p
u/Z+sB2ho8qGuAMHdOF9TTJKhABjxYTPMQuI9VKu/aJMKe85yQMXHiMu4UpG
CyojGmSuITwkhF9CmrDoHmF4y/j2cCQdZmf+zlubkBogx2ZEKjFjTJM1S4Ah
oaE8fLr1mjV5+huHWTkvHAaoNhTYKBKSFj75WUArz/zGnezZx+0Y/4AfQK7W
5PNw/D0v4TnzLewDY8k1YvF0F0iUNxEaiFrloUwvphwgktRuUhSDKbcsM5OX
asqojq/H/5lhZni6OgsJ02b1qaQ7V9TftC7QQtWV5jah3xVje3+He70zoSgj
oyfebko8wtx2evDVuqbT9UsLDl/enLybhsdEKMGI9+PWvZtVFn9ZiztanjCA
FOIXrgIu/+RqwmXe4fCqbawDuYK6dN3kJk2hQWqP1XFYe4kOYwLn/Bv2TRhj
n/aERuIryZT3lkp96aA0cMLJJYjOArENWcDPW+Bez/u882SQNq8QvsT84J+2
F5G3clTxeeZwJ2kjyHDbKKJOSgm6tMCbIACRjBMf2GpIJzNcoJiEoYp0NY4V
klZIms9QEucMmQjwD4xcQwL2Ju2WiNplb0XU2//n2A1KAuvMt/HALATJLift
nXXGl4rxhB63mNTGu8u7/BUnj1drRMGNOjXaexXtfgKkyyDZjxFuDNRSrJLB
7j0zjsMR6b0aw2EN7f/OLhwLmbFvaKC1SphKkXH3uTZAZSx7yQWqxT2GNT2L
lJfBkWRtF00VESrukjLbJiECtbH+Nry7Fk+rbp9CRjCpAwH3F/2+wyT3aYyJ
oY+WKoLK+Yo1AI6NQXnd1dceVAopazlJEu1fBtM2gE7f17PI28FBMEsle5g5
t5TD5EPmvcEPQZTDI5rYG4WDVUPAihu+rEctXf4d5dren4zk5RUH85CJajA+
1jtG4xvkGevKLHKnNM6uaPoAojQRcuceEUrzaHCnBUNFK42IOujiH722plDk
TVqbEL6OpBg/2Ojs+WVkbYXCyC/oOsr91d+GEoWne1DFs9McaFQAcEzIo5iR
zMQWUoIM7DfwJZ8LdouSCfKIBEXwsE+K335Hh42TzYr1Lf5NJkjETwCGXzHL
KUjtLQxwa6Iklz0m+0C38hYcE8IlWH3clQ9X27a9NIucVCVWwXxZyOU0H5Dd
IKZUBSucU9K1fEdwJ8NA+y/Nttg4B3V4LkSBlfWbWGEpigUMbGieEdlqw7yY
8dgbOusmYwnoQLFVfClGYp2dZkWYWwxLoyotpXyioGiaHj09KtH4GxXeLkwo
kzmUm76tmdOwxwT7dawA3NE4vClaWxhtGFNMUU2Zfk3HwnnZbyN+IjE8NXZ4
AC8lfkTcSYeKvayPbMxDEIBijXY6q965CjsHJ0YJh54uaEJycMycQfnBzOyQ
WcwCvbWYFhkdfD0c0Z5c15xjVu4m7dwYeN11YohQRm/B+UqXcTT+L7fLsF2P
rSa7YUcyBoGcuCR+nk8ojKk+OMoOXSzFUTblz9ZPS6MrWyl6a/seKJWmFW2R
SwHhxtVcwdceI+Pw75Ml/BAMLpxMEMm6SsMfhCx8PF2PK5XupR5ifY/AWGLH
jY6E5jD/aSGsyhvv5ghSF2JTUC/sNEJfWEpFMkV21YYRRcTjx7XkVNwh0ykD
9QIl99Mmd+ZIXvoT5VXlTxmsl4hhgNEA5KZN/XhUQGx1fMxIzN4vWWqKAfQp
bIJlmC8tXYuow09k0FlAoK5ClKWKCAa+U+OX+b/5ddugDCUTCRD2Wy/rKvNz
kvKS1uByqJVaiU9WfEpIKSl1D4NbewfyVFV2PVOXIJ4qhpUDjKpuMkeKuY3a
90VAzStbCSIaXmkJwOoUEXJj6TbqW8j8etGTTc0u+CRrRjFPw5oKV6JDdebC
49RUMCJJBrEgcbKDb8veuDVuYhIcQQYEs5TDO3QWGDj8oKsT2gU6IrgQq5gB
RN6iF2oS6jykfcY3BjC8x7naI/V5bcgmijC+AKHWGpe5eLP45ifVIbSK6ktm
WuEP6Y8lelY13+4zy6+fLvYgmh9gfCBhxMWbKv3ZCswT/WJV7Z5Sp//7Z6kY
0IbzRMI/4KAjK+X06i51OGJwclXtOD7Kp+i9CqSBbB0cp6MO4w4sioom2JvC
Bl3P1xA4FTmjX6U3m/Jun2UYA3XHrJWhpE6ol/Dic8y+7rT6lggaaPTk52v9
YbJpulBFLqXek2zQowFZtjOXo2v1tI15zK7mmtXwOQeum61Ww4wKsIUOOSKG
IfW7qBSSlQDmquzzRcf3EoUU33tLHObRo3uQVCpKVZTCWWGrSQ0vevTJ7i9m
j8klxx+E67jJWIptA4S3y2SJIVVbu0f9tfDinVM9vON14kTevmiMf/GTt8w5
uW6uUCn4TjyJJ9QM5TiRjR9KIxkzcZNSoDUoECn2ctcU5E/D9wf/6F6WtgY6
eab6QgbG8bSm8v0TXptTspHY/o2lfqiv+s3NeNCtNd7td97x4YGcHdpZOo59
pgMcihnxEpp0Annc3QUtNdefJHb320oq0/u6JomIGLpViq81/nalJ3BMjOzG
J+2O746fbzjJ1AF/NUgJjOR0zwOMsg9eB/tkHZbi2DHfi/NVf6+AlRgg02c2
h0QobvKy9Rj5dhRC4hap719NuCsrRXyFDHTc6jDhwezcmGvj8FfVLWJGPNaH
KgsXALahmQoGKwIJgZtU6vf1fHi/ItRESgSQZPSwjx17Vkytlx0UadpiN7lc
FPXs6AZ3PbiOhagae17VO37LOfrMaBxFsI1SER0wYYXOT7OsTbVV1W58eHTZ
wTUzyv9LvXcDwX2lbpoRCTdSzz8k5CkN3Ysd0qncUlka7bLZFe+v0kVyqaBC
kGgj0Cr5iwuKg3Fbwcfy853wyyPrwBmfSg3jE3coMxuhZSxb2pdkzoZhE86X
qNWmP/Jjbio4gVu8MwWWVG+1Fmz5IqiMraashcFXnl6PD5Smo63r95ExWxas
Rn/yiI3vSHlLNGxKiW3Tqy/gql5Tok4t3jmienveYBEfc108nhv/MopuQmYx
mu4JXer8ZKwoglcSbgXkT/neC+kRSqmwXPp90HNS3dR1JtryaGKcPnts1AD5
d3z0RYVyTg+8nC5ynfhBaYjFWnvGWPrqg19ZeRHKpAFCzzNEnzGBxuNrQYEd
LVoKcgZY/Fqb0SHUj3/wBXyMIRLUO8bgFeoZIx3Uoe1GxRSQmz+n34cQGW8D
4KTnwOCKQ2AurfNFnwM3cCb5Y94J1KS3iuWwkDY+znVeKBsiry/KJu3AP93f
/dUb2oKkehd/FphjePvDi0o/0GMQcuY+coaFFpwdZcycjUC5QWizF/9BJ8fH
pOaLs4xGMsJJ98oXcilUbHWLkNzcOoBeqta0vKf5JAIhDo8pZM884IuIY8a6
fsvEUn2G/jUPf1YLuL4VgGdXd935cmLB2ViQTuyRKw/GY1DUMZnQOnod5DHH
dlzePLJy/0B4GPgQWs7xzCmfeGat1cVawiysQPRioZgWdIQl57uOdHMOGBH9
hK5gStYKd+WkY0h+FSRRTZgWNfkj47DXWJPPUe6WLiRIIMU4uHE+/72W3kiQ
SOYgrBeEmHF0Jdcf20c6UZZo0dmp7QcpBKqYT8jvN7xv4VCKfGIAhffJ7/dN
dLweIlm9wp6wY8mnllwMLBlo1F5xfXIY77iK+8PcfSsRoM0MqiWTmG2Efivz
L3KL4a4YRRuQIvK76EGqQA6VqcQlQYy63XBGx2lZIYswNuv6PR9FOeiRAwxU
5aSCnRsYe2zc1v2S+BjtBkD/8DFJ6ieMCA0E8PcBi91/xT1AYGqyc0R88pvb
TbRdTJhWp1iimzwwtNFNIeICCDdNwYSCiduCkejdFjOF1h4cHDtX5eAFaIIg
XuNP3vKuVEZh713Xr8PMDdxTLAvfgyMBTGo83r/W8cS5O4+5JZWGn4lgD0P5
0xSyQliSxkSOhblEo7YpUkm2QEf+HBXJvHM9ba72Y5/bDkzF020Rs0DmQxW3
CRWwQTO9Hpcn+JMpl1FERHp2QVU2Z39aKwy6qxnoey9lZenSkEMIh2xaWHNF
ZO2JtAKlmRixHnWG2+hO3cKts7b80bSS92zDVAjJB9Qm9kUCzoRYpDmqVU8D
4Kgz0EaVH/7AFxhoiij3+EbZ/wZAQHbsHZAx884RXB8tYaNFb3dxgUFR8lpZ
4Lo2U7dHThekFR0IKshw2P5pt9etgrL1S3w620O9dH1P4lLGwYm5cpcZL7UX
5J9UWG22CSeeobWliZaIMv3p+q3Kz4dFhjH0KNiZ9O21l6M8GORisupvKPBE
t+knU0WSArjmA2mHLFw6gY8DK3inxMeyNf9kKNpme04OXM9EYdMHyzNJ/pIr
G4yW8BCiCD08HZSknzVwyVFKM2SfcpwIz7FDiAfqflbvRPxK16bQ0ipJfp77
lhCqI0/VY0ZgebIPp01dcKjZtd20c8hc12EoJM/sQ3foH41oocSBPf4hf/1/
21Ji47ATW5LXGdfs/dQ04WYU4nzyL1XMtNQz9iehIM36ZkVb3wmz6VoHSZ8X
dEIJO4WMvHP+rUJNBXkN/pRthMtKntB7p5wRG65RDCeDVekbTPZl1aZnPDQ9
aTdcPiKBJ2agSnRq1+48FcjSdRMjS5bRcjStClcvIlFXZJcPtvwUpChShS/j
dGPfBIQcZPmdp2BjY2oRLBrXr/Jgn1Wz+6iYAxo1EGFlNsvAM5KciUTY593n
Oa8SetEHg/kH4J6kkuUFnoFVbq3XGf5y334VoLGYxgVVXohc4BpcE8i1Ix/0
dDrenH/Tzthy22PNUkrTn8IqH91SxQ/5UejYeVekidXWiL4Wif4hJPGxuNqp
szCrIcWY7MTEUUF4ZEL/4ZIUvtFyCHfYnCtfBE4uA0GzECn0PIS+0QpZtlTx
UbglBiL/C0kDzwA6rkh90oxiSdVHOmK1mmNGtHtIhOg7jlD8jnYs6L4gayFW
1k/kduRjYu+sFRLXTR6bFipMiwDtG0W4FEvbn8fmCgLmynl9tCqdzNDcHIiQ
QjLspYO+V3bJGad6FxAOwMltff7DdJlvhQPuGu1fSAH/P9rxaQlqXjkrzW2q
nUljWz230GszdWO/oPXP1BPOirOg413FkZUSHntIBOFUyNmm+6cbU+mTicls
OXUZcjeW2wXDV5QFJCGSCTvHGcGi9HypGAUEOeMSSv5m93us7i46sOjr8gir
nyuH3iaa0/67EGQtrDi50/moWuafYwckK5WbD2tU6ck4NqwjrFva/LqfGVYx
vbXdEELZP8XHiJpLaSpUHdKJYe1gTxA+fCnqExamD4g0pch5PeMMCvstDqrb
qWxQQc/6lF9ya0o2rbLcQZpuoTUJizi20/GANMez3YuZBa5K3npQKkeSxylB
ySRzuH/TPb24IzlPpihb4i6ECS7OSdSnol/9Urpwm5B+S9PLK0NPPFnlHhI9
UdMpUE4dTxhjUljQoHPgoI+Cq6Mirkwa8MeWG0S6DVvVtP7jUWPAddronyt/
a8tAszlleCuDZYpiyKDFLirsHS1aAY/T9XsfANm3sN0ufNwO3rPZqnMdku8l
kwomN478w9ISKrdaer44saP9Jv/+PFJxYpxs6ZaqkWDV7ia4mWW/UyXW7ual
MT+7GI/hy6N1I1wjjdn3CX0BydR8p9wdb99JzkAB3v6XmJezKSp58Ay8/WNa
mpoaOShffVY3t11xgV7TOk0H0ZoJnUI+oBQz12cQ6DS39w+UmjBq9WGo0mTz
aolJS43WA3j98B/XRQnzJzcOkX5UNB3IKb1HwE1GiV9XafP0pVC2bdRCJ2Ch
p6jH4hglV/IJXos+/Crsnxw2t7MrcsNaB9Tbn2uIOdjiDMaY5hX9V/ybMVPr
s/YNa7NNpD0oTMZmwR0eyt1WEMMk11CGKm2m10+cktzuPudPyuhWYNfsh6kz
Onw62V3EwR/M3oSjvGIWIu/Bb9w/ZH3cOjs1kgfzA0zKjaGh3mXebU0k4p5K
/r7X730XkJjyI64v0fUgS0juMv31+nlZct+kpxx93y6y9lVjwtos8hC6QI7f
fBYrp90Fh6Uc1qUTsQtGt/+kKRDd6oAfJwiBmeiPBnM4MXyXkk0S0j8fv7Lx
77d/n2yhTnf8lHDWtH3Cb6vTVYgYQvwfWhKN9F3+cQIekgRXdL/IlDPxbvvg
+zm3dQr9KxBIstbWUeBUDMb9z3rqPLcXtty8zXrTu/k48/QqJ+FaqqHN0G/9
9HUZnKIEaqFsqNvLC7RILuH+HUFU6cFk70/sZULApY/sgXcF29Y297Dq6Izs
7BICamdZ0jP4bGA8baRUIKuHxfedYnkhNFqDvvBvidTMN0ur/mL4dPEFvq0o
vLDrZ6AXSKLeZnCo4xw+ZUsQ9SfFqs7PCzIFdUmvpwc721JaMTSq+skObplj
8ue5FGdLwgVrldjTuIvZamWUcS1KUd7jhXUTUr3M7BOL3fJ0WEdrysGx231P
tIw55BDWwBYKkuoqLsO/fRNNR17reme9C1fCnFF7lLJWUAU8R3u6T7CVHeta
554ZU/C18nD8iEnYy2kQW6TxihgbRnvDOJhuegku/sEU3qg9rh0cWPVnYiia
8mP010w71IX+jl408L9p79BG9X8CnuqNb2+Tkmbig0aKBQ9NyKxSegtP9X9h
mMaZCK+loAeQ9tUmTp6wSew+HV776AFa+Zd6o3V/2lyxkj/54IcWM8/LPVBJ
7MI3i//BEnMtgODL8r6W8AqPs0YKU3omgRrx+G2tzVY8NaFIzSI83Ps52/ny
Aw2vh7+W8LcSbu0m+tSDd/mTKIn0aBLjfcCkngsufq3h3jUvyaETz6jmskZN
Yb1bkN6THSYKvf/HRhioJs8Do1Udc5dzFV6XUCJRkmUKF/yVNYqoNI14B+57
L0taoz3gaiKRvSaPqLri6zQSt8C6sTF6TZg4h7rm1z1LRlIkOtqwvbu2+lb/
vY4NW01QpFDrudLw5OU3WLlj/eEPU772XJ/Eq8t5E3trXRl/ZU6bsdpnQ0TJ
TQJ8vDkAlJiTPQULt/r8TMzUwAn66SOefbWWIWcXTaNdXvKg9kkn4qzbK+Oi
+kJBuvsdRpxmCS1MC1z2vf4qPpPhxjfayTdtWdkCUQ+hPCMNoQWdkmygF/dm
dynhmx1HyApw25zzc+n1utdVs3n8yB7qO1JZg16C62xGdNTSP9pzCHJg74Q+
WNVPiJD/e7fSYqsaX4ToA2fN5ci0jkBxgbkkqEakbujnxrGT5/a3tFEsP14F
455CVWLT9bHVOdQKb6AQ3RgWjiz5JwUwDnrqXjhHnZNQ2Xy4B8jV/kSRqzCx
9ogGyNcG+yxxJvuLPAl0wYukMe9xm6bmgmEJpXWwZby85ObVuY4W96vFJW3z
p85RJe4FWeQGTsofuIXS9Az4D3Tixn8Mkb3727NyliRgl8gqtSBDRQH3uWr2
cljzKe02tH0wErCM63lFdf7v1I/xbOpazN6DYJwdkmlv+hXl7am1qbKuAmqn
A5Y463J9FkGRgavgAhjwWvf8/wcDHM88ZbYy4J4/sGxK19dgST5iOzAh3m+j
4Mf7pCQ4x4BroBpmAcFuwZyl4wy1k7khCiRkZeD27+1sJLkBSTCG+l1QDjLy
eio6XHMBYqq47BvGM42nMOXezZj4EoNwVBCxMeDTEqv1Tnam7LKyXCQi/BB+
aHzHbbpLNmNGn8ZZWlD0U8CWVhIvslWjwRKaGlvz1Zq4ZaV2FooyjaPBo+9q
8rNyhF4h/1TBZ5D4xdxc9oV9CLFDJgl0iJvHciNUiHB/WkL7VkgVLgDQDYVT
4QD4Y1psf7uQ1z+nII+zINmb8XRfTuxIDsa/qTTqWk7uDaJ1cWakWj8gcoCY
pqOoiEp7BMvS6x2lmBuZX8SG73HqQfH4X+il5tH2I2x267uYEkhJeHM9j7Sq
kZuJPljSpRJiaZa4kefAIcCaHDBPQUJghHTyY528Q7gzrz12rjQHphwlqh+t
dgUVPUWjO9jDrpplq/r/Qsv5CE2SQirBI6d3k5IwQyDnJWvux1nYX3LvzQ7K
3hEs5du3XCijO9PfU7CKViqNsmOUBvFdDwJGO/PdZtanPvWFUjuQWPSO+aVh
LAih5wM9p90N1rnYDMLZSlYACNPHqOr7TMYzF08AUhK8gSBIqoGKgAyhTJtS
LrWoBEKxTi3dAZ3kwaOTm/Wo5qmBnfCNfeKTdntdq8YmWn/0XPmYATUEnnDb
iGuuRqdclSrsrDpRJi4c12Db3gS4KC/O5am8DsL57s0Xg0NkzdNpVVAyhNB2
q6nKLGD+b+sOLkZBaXSowixB6WvSKrcGh9CB/mq1VyCwavfKet3b0hsbejbO
V60F80DO1n2gpG8Lkng+hQyRssiHBwqplJg0eDAbsDllGNTmjB47freP3onu
4jynDPrTwGIkImJg2KDk7jl8dXGOxDySrlImMrIoM6sd3PO1NsKgiRclu9+U
T9FF5MfhtviYkk0kp4qAFHm4+wjNDbf9Oq98i3NC73c4qKxmXjvNzznLrriG
dHYkUDtyNlCr/NnToKakxf2C6nvPRZ1HS79o/70RXnCSqGCFjC/4TfKfZ3ZE
NIqFjz+uDWL6YP/PI91eV044M7Wg1KV2vNxV3TrlQi7lo/v0UYl7RvVgw1wZ
Uo5FU2ko9yGLQW6WhON7Kfs2MHZyCqkar1HOPzijDZbWmiy51PXNxwjtCCXC
9xJ+j5/tr48iGbH8pmTdRnG8+O5ZINo8o4BZbnNJ5aYS3v8PVcRTSWF9Ii0z
8+P67wzdMM2uXVdVURXKuiEeO3GY/jDw+UN3AtSQgphFWP9BMmYsLFZHDVT5
NEpf4tm8/VZRtS0VFCial1qLhRDx2HY8KyEcjOfyH72tEcN7GNdOFwW5NUaw
X4Mov8D6+Zhfp8JSqipm3xMKjuKDT5seDx6WDB09goQJ1vW7yRkXtIUfZ/nr
RYYIZ0G9ae0DHzXyf1OCw1ruTq2bcD3nZ2IZYmLbm6Tui96BWZAwUgXdIWPG
/8dYcegjI4+tEm6kCdbyR3LFEe1Au3hZJ6utihHzCL9m/i1RBfs1n53ktAaw
UphjC7GTnkEXvfz+lsInf6DwrAJxwxPtFjrLXhoZ+DU7qPChPGCi1DBRl5E/
6sFaix1/ff/SQcjhDylnWlCVFdRYlcLBmjdyJurzQef3i319VOy3/t+QgGsQ
ofWRgJHnINCdb248Imq7qcEnlB6Ltq64JCNpc6p3p/z35SKbaqDoM7QhDI1b
yYqA2HUKptmcCtgk7+RMsrq9fwVIIW/E7FsVY65rNGoW0P9m0yLAbGf+VTR7
hjDAZmm2B/U3T4inhImqlMeSp/nE6JlErnQ/Ga5Rlzx9Gs1nzWchZBs9WnwZ
QU0WVUASIWMJRL3EXGHwslBu6Yxlxd9E6zf7kKX1BWYYEkEtmF5+SNEQncob
RU5tVR4q4IW1IDtUyoGTt7CcltLOizRgbtUmp1ULxGcc2k67xQiB2KByBLaW
xEIhaaMUD0GJ/kIKyFm3Zffp/dDIqDw4h7LbacwTT3UJTjo1hjgChekRuv7i
k87cOuYyBjdj/Hq0q++AqGiwpN+7+J9sgGo4tRQExCxRm5hXdSu79oh1ea95
mY3udqPQ6ATh3SuJUY+xCY83pSrYChQmCABoS0QGnHuTUWdv2ohsjXyeEjmX
ueTXd1+E+aO3qSOca9e+WXgNj7wVc5c++o77cd/M4v2F4Ut0mzFGpp1d0qnw
OjjflhNhtMcvssg2hkuQzM/UAGEQrKNCx61WkbWv52cQ40ZYmseq047OYsWU
YvfY7ounKUHG/VFueQxHrpz8MY4KatgG8SDsAHEwlwaNSjo/MAKWIXTMCLpR
x9u0hmijlnnC+y3IkIsPtlPTuiD5QQOsRRgqs8kjg7m1ioztAqvbEUodha/y
f1CgIFLVgpKTxPsPgvsX0F/xvo1szaBqreqkB31LIeVsYTvsbrFFhlbcuWyG
QX+fuMnXT+9QWMWlBaN/CEiRuW/nftUvnvwTCCfKennEr8y7PrrsvruUx3YA
XY5EO0gOjrRoT7dI2o8m3EFFrYctxfajvFpeOj08zUI8D1ErP187bKll382b
iKzNk5/LYOBYnSOcdqHIcV9Ve2n2PxS/gtyowCoHpeKs4MQEAPRb26Gucg/r
EkJpomYf4Lr/4gtDX30tUwNyK7VaTB9Zkg+oKltoRVf6Pq14d4+7UTFiZYE1
Xx7SetFdXhI1kAREHm8qXRoDt9v0j/ca7dTKnE13YqdSO3WvDnhh8m90rVNx
yf2OgB3JLWx2NgINhp/29wTRVwyiTW35TOacbdWgr1upoO9FAFAdAyek+VrO
J6fUgxUtU6L43mQwnnrSSMs6QpOLRKDoyMNTSU48P5zeaJHw3NrXksldSWQC
ZZahsBtPQeTeD/o2xYqiXkcZGStgJG8qBrP5DrCYKYuzzD7Rx1DagIPfVC9G
b+MH1atHWE+Ai5bpEQn2KfwhVj1zEYphnvluXuLb6vXdP9dtmcnz3HJSjieh
A0srzDbUUwoaxSuqpqNrAO7jz/fA/79ymXyjAngV1odRnViV8GkihBaC5mXA
oP/NT4Ygw/ihK2HddyTCcQMACpxT9dR6AGkmI1gU+ZLissqMW2iHxfDDQxTI
6sR9oUV7QHvnZ8/XNxgZWT2BG8BMhDsftKYWyoWR84+Qkb4LnMiMVzL5gGIC
9QxA9VLx0w58yEeXxz/CRAVA1Dxn8g7xMB9/wUyyVutHTGpmEQkkN2YYGyoa
m9zCKX43HHWtNTVpJZjgoIzTMz1ubKyuJusI+oOC2HLDRlmt/jIh/b28sszo
xEYpXxQw40+goY1qsVL8SLTc+TAsfB6zCQGylKuJ60HdFFjKf/DLzytwGKrY
vbo4vs3YnQ78NOKj7SejfrptoRnzHCWGSA6n5Lncn/gNGfcuioGdJYULC7e+
qrorZqU/xrdrB1mxyAwHXqKD7Bdd4GiK3gv0dECRNaWtDyBQbk9H/iGRbm5x
nCQoQ3AKhTOE9cvkfdVV76udEM9vKdPSUk/JZIXrnFdvEmfhVYso5wMtKkDE
uCIQ6+yudPC0dOS29EPzB6HcBsNSshMSpgnM/hCc3zxjXEd3i1OxSYL2YUHH
gfto2Ohe/kURkuCwqdoJ5IupU6JMys3cg17CCC+NvYliEc+WpCdjb+F+wf2N
CEGzZ5pYSJigSe5918YEgmD0jqix492x8S19zMffKmyojsZ6Wh9z3Y/43w6i
jKm9BUB5rSwl4nx8QD4RWOdOk3kyqU02vTG3N5/GBok9SxDyexDBVnMCU8e2
ZHJgflmJhvoeScHNPf4jPC2EQ2JJFP+LWvJVP8s/QAXwo3veJUP8eVOeG4kh
ZCD87bjRWJCFPwPtuUr8UoWrwwCaCHiSUW2BQqKvQVh33I0bykNIWnJ+1Y72
sy5QU0SwQAWzEM+30HWsPdE4uubCFgJE/1VvTCbeeTQ19q9HVEgco67DB2ST
GJXYrEwx3IjdgxUEAgUYZdLwKL9OV0biwo6x7bdfQEvKA2cDcEgl2P116vwp
rgAe+Vh27CTdycb9NiJp5ZNTFaoYcRPHOJ9MjweLoYwcq3LnifBsSZnNpBCy
B47xbwEDtsUpxAADPdmujlks/isP2bDg144Sq8MIFfXfUuSJlB5jyZuaNjSa
9+akLVn/4AyVopy6c7Fw3CfHlorIjZVxev1bscNuef4YFW6Uz1sMPcHU6S1w
3NtJp4AOpqyxjtOhJ+7orXzoabtYxIdcgV/C4JanKMGpar29ziKsZcaU6RiK
FAhd5Nn/1zffcMNsJ5k9RB4K1umV/mEjxS6y67piKjU+pLGOrUbfi/gg+vQa
JB5aLKZvrexuo/YJmhHlpw8XfN3zmiFdaqcKFqFtqwDW+hOAV2M1+SQGrnQt
oQFL5f7mqb+DWoG34kooEdMLir74paPlXlYB5L0EQQ2ryUFl7jcMa4CQewq3
5DCbmgxRGotB+gx7+pikTKL1TYi9UZCIxoKCpFQp1Z6+F5CcXe9Hosz3vKLE
gzh5nsN+RSHogap++su2cnVhivTe9f42t26noZClWlDtF5hFGuE0qFax0gV3
iB9L/33Hipeqv3KKEJnd1gQ1wB7da5bCT4PZYiFt8KI+E7T0W9ioyGJ4fdTt
ypFbhhh4KuUBz7JU/eQupSH5IY9nyfk3owwllvv8EwwJYNlZoZesu9S19PgB
9x8yiNogtrqnSf99359Ep2xI4M4HGlPPcI2FbEnuweds+TQQ5dH9PcU8pNda
RbMky+cucBb3yTjq/zws4X+PAswGUCZMBoR7moHi4zYBeJKqW8vfHIuE9arB
1BrQ6C/1qnN72mTgFe89sRsvPbDi0PKQ6grFb8DDGzOyGD5zXCeKttDlMux1
lTvXUwDdD2Zr3KQUnSdvnvr9+xAclk0b7nZq3b60o2Spx4yvy1HPaeXLx3r2
aFuPSYcPRn3yTxnwdbd9Ih1P1aiRVcmux/DWu45J+YE/EfEL5AXgDxCsxFd/
cn5R1FdljM3QJHftRCbiETL/qPEPuWrOiYTOX4dsIFKS/ZXV+rxVNYjtJZn7
PLmC+QDqVzM0Y2oSbVcl1EEQgsZscNdudRsZKV01bekE7riDpnLHbOTu1aeY
m1hCgWvOw0ygLOIUdcQ6M8kmtlzfYeYjKXGEmAVpV2neLdHt3sXyrfHgqOri
GKR90gFCbPje39BleJvJUUtxbB6M03xldY4pIEOnAJNryIQn0XqDMqiFmh0N
SYZ7ErblcvFcLPjOUq6ikGmgwnCSOakJT5KCicqLhInQ5lUeQ6W3lkwcRirA
IjSiiCphEFruUwK0Y2V1HrYnGjwrX/Wg3kibimqkMGTMlJ9+F9rAQoT4Jzx9
oMwsCX+fp/jGDKuxvEDzc+YJ7NeiLI3d+YmuOmzVH9rLN36QhWbyly399gqU
vrH25KO6DFhR1Gy2oFsBxtv0/m5W3HB7JqYK43Pbcmh3NwH/cUKs/8DCjqVd
MvA/0xBNlNY3fBDfN970ECZCHZMr0jQ80RU3lYHb83daYOmUww7445dzPZSO
tWJxzowuvpnY9bvOlXTU7NWSSxKH3TO1ZvKT7bnnrqTdKd3AkCIB3v4NToww
B/YwHSVBXBlopvftH6ILlemaZqvqQFz12N/FYOEsog5WlrxbZi2F06rmG+8t
2X8fFQM0hbdEYWOWRbkfiSro0ca7us4IJ5HA9bV3VtZOV6cOsSorg0FQ/qv0
rOEryCfwq+udU7AFDlhB6NF92u7cN12Ug6FBxXxWQIRtl2EJcQDR39uFjYD4
kV1TI/m0pVKAmTHJZ/6mCnve9xJFl/x9DfOwmUWKPIc+I+kNb/px3cJxNEqV
uCe/8BfPbpgm8bGLh72nH4lOZOxYq+gGKD4paZjllUdpqz0TZfAqWqeVANlm
TQssu+R6VgxaR1xmNjxpdoW6l2fRSesOoK3fXJwfA6lqtNuwqsvPzL1bp2aE
FJ7bM8eocv7qYH2maPyIZ1iGd5VLSd9/tEJ/gTNPoApxhtHdLCMM7JQLtHTP
SW274EccFxOIxDysj+ZYAB3iusIKfcTgZuM9xYtVpPJ+imvt5dh1D3ZwPE3U
zbBhIiG09nygC1F/vM/WYUnu6zkPJ4MdShLlJL2sS1mCaqyt//VlY5nq61Nz
1YuzKkQh6brrqWGmYWzcw71dFjzKMNRpg6ldyGoksaWy44VNGHXQzb/KY2PZ
StpEgCqZky/Qyt5CuOrTsMW4YU9qF/axQiVVxlq937JgWwJa1uhx+wXfx+fQ
QDtQr6x6ZcZsEpyVIoyudX5lF2ED9ZV2MusFgK5b8zFFBfjgn+IVb+EICBML
UbJbUWRriNsKKgCAgKG/GlJHNiDuCZIOPUBDsqi7HxiLPM28a6Z71Evs1wd6
Km6OA6omSbE9mbhurFYHARvfnRU6eATm7jfvVAKdm9gDEKTHcU0XoGERK7LJ
JwIxZWkpTquj2OqbW2M/y54Iw71FNbAgNPvQpEApMadWFf1v7HcBNThEgrCM
Wii8uzBr1TtofmSpkDwxvcrtBRrKoYXfn+WdSY5tS8iCSA8FcMD1WNd4nTpY
EjOr2anuBxuww7whxUTXWEOubm72le/OiffsjCU2l2czAjWT2WR5EJZHYCDx
uWtz1MYo2NbkA/o0HD/DjnX/wcWt/HjW+6GLwddjwA6O7z6XXcHVW4COFrw4
gFeGsw61KUA1Lkm0xRchek/PF0ifIHhSZE17i3k+YdKZKt/83W5WFXvkMhgm
hjWHBxDta0HsDAgoSjdHEw7pVh6K5UzWH9TA5rQm3lmQ6Oz6h7EBB2mKsguF
FfDXKDB9p5SypKSPq1MS7Dw7cgCS/zQRGgK65yvGrduSskMybbOB9brtqMQ+
zBMgC8rZdfec4kcZNzKs0KVh+gK3diH1yX4FutGjSFSsG6PvZYUpKf533Ogu
WRsSsZrEJ4uY7jvFLXjcb9eUBfRDv7w9UFu2jKbpVMwTjE2fc/F7x0zemY9E
JWwTeDzTpbjM7NytwUM2s9MCrRJHP3sXd9A1XBTc0BoXb4U0EZa83cCdRyk0
xTMl63Zu9dER/MoiYuhF7YqSVLMlk/ywHceMJ6W+Sa8TMbDoQ0pDCUxNlIoV
P3l8w/1/bd230sHn5LOwscF6T0uDhIbWtQK+N8hFp/UEzHpNe5dwuzIFwVqH
r76WRNRs7bgcrEyVelI6LyiTyzbbaoyFZhEIqc6Qa5Omsjrg0bMd6DWsQNCM
/zIDmLReCiXXRbLdL1Krjqta/MwCs+XaoWfd2vcl0o1u4ASFY6VZOqzHpg/9
mRwiVA1ZiwL3wUeTYrnYOEsKaEtFu3+p4xwpMn2DMjThi1/MBrWQbIS4oBUj
yvcohP/y9CBVhMyI1yOMGON7DZj5OyTDvl0pWKPwivvA/bvEImUCZ/rR5DDo
tPll1LlvO1HSd82iaOG2IDAh98J4vIOV5rciwL1WHnYEZjHW/2ez7bwLtHrj
KXwi8P1fYmzFBJs+yZn5EYuE4tbhCmyN/G5C4s6AH38pxUfjLs2ptETCjtcd
RVEZKQ/1GVL5RWhdQFiEiM7iHo31RskL7ZwuLsEizmpZFI46tuHBt0emD5zg
7Nzi21FHgeGandodlpXatmZ4qb0V7RQiRgXBVF0K46CTLnKrJL3PCbG/A8S4
djywDF+yTQE4QnVgH79rxeEXM2kFz2uDR3p3cwr3/1fBpGQjWPxaS8cNPZkN
XAHHLY5YKpT7UG87q8NOpLF7DVwf2yPBxDJ0SN3rTcjqlz/gM8VZ097lgEGH
UjtVJO1clIZcfAOSxfzN95eTSzdX0TTgb2vXK7nc3KEFiUCeacewy+AI+GRU
DxT1dwqHmt6gFxdmA2irjP9yNBjT5WFxab3KqoIJypYAvvMu+5TLAmQM7fkJ
xfox5jkhZgQ5CY0pnRMD+ucoqgecK2S1E1IOXCFKDOH3lAUmxCEaBjH7GhSg
bWBFhIF9ypLNhzm7d+8QpdIbw0cwTby302/QCGrn5o7010zqhb6fT/vNL+a4
RApmcnIy8wX2j9BPbWnmyvfB2gUQrNS0Uzko8tUc5dRqy3dKDUCgx4yMAB0J
24XfE5JV4fDlylwZ3LRMWpkrh+O+ReEMz3m86SFifU5BK4KdgdomPS0r188f
aBsQD6jliSKiOfyg7p5y9klg5RWnAQY3jHYCWwMjiFTm+VDEOQfJWnpAtY0s
dAbFFJRlFFoKdnbgKjfab6gHdbTvxkUMoSrEMsadaZgVx4e6kQbtC+4IM2vP
2RYqx+jtZcwAaNgxqtV0Rg7NJp06JbltTBEJu8TVn3sWsynxzewWceCa6xgy
WdlYW+gZy/9qkeqAZAO1Y8AuvqMSRxVZjw7QLQzM5cLm5cHnNgtvB8zIHs/u
7XQx7Bq5/Gg0L2axt+wsLeR44g8/mHlGmrEpJYKObRuwHiMp7jMmyvWA2b+g
FdZKA8zDZDDnwpkZAccuAn5y2BINsnCBN/muZ1rZWK8scvEuikGp91keGPSa
+KHjU/ZMe2rrzpA3dPgXTPvTr6DbQlGf6TqsMUcdjTXBnhnkPkVO8+kdtIWK
/tN20hv4LRmUK9pvwAtlG1490G1LlbYDfo0G6xSdPPMzdIgdVJaRlYPlrwXm
yU0iifv13bDogM2nQ18Rpr7KG7Ji8BxxLVupvS7Yk3nYpssiyFfF89K+puTJ
CS06hNyYn0xa0p6Zi+CWjHrBCyWgRlJCyhF587mIdqrUJPWLiMgH+IqtdLmT
Mab9SmkC6J4RtXxr/d6fJCoL+YERif0cboSqe7imcstgGmifctFZe7Rw7KKD
s28fc4XcElKph9Ux8TC8RQDVWAlSQQe29Lmmy0pm55RUWwTjcO3B0SfEbYpg
VzBPl0yt8U+t3vTXDvBifpOVERrzOcqCJvwsoJU1ul0n0yP2WCAUo7Z11WZW
T0kKs9LcdXyRCYl0HjGVFjwdsVGVfDtdDWJXMcjBpiSVGxZlGV8Wh3FufgQT
2E9S8C4VDA2wv3E70yDOwF9TRDoqn9yCBZrkeaTV8NSXiEbWFpyessPSjL9f
5eZkBktRoqv/iTPO7P8ocQXu2nWVqFpLo802KRyDdPQmGpYkZK4jjed5yc3M
+Fy41QwBDQFVBjXBppP6b4ewvCS/gjhq4iY3OY7EkdBSsXfV6IAPwfkOspQB
e3BxrFBVQInqO9ZaEpYJaN5kUzVSWp8YgvEnSeYOIExnSfH68CdE60cKCtQz
lrcU0WUd9MaN9Y3jTy4WD246/eGc10J//34X7gw5FJ23S6VPFjFGcjNiYM8+
Oa0rz7t5AJViVacF7Z7fHLdsZJodeeIHJPrQUh029ySaWDV7lyV3DARUq1lt
xyyi1VlN1aLlg8ljyan6Lgj3L+UF48ew4Tve/o8pihe8bL6brhOmGcQToi61
kdxG+9XgieOwQvnbzqoswZrmyd9OZpB2gefFa/nq5Hl8SjWVqpjRd+gQTI28
9Gj4YI8Mdi3whXlq+lfhATn3uAjpPvs/21CvyonOwCoM13zrw6bjTZsLACPB
PLXIJufc2SW8i/nyYUjA7zLN7n9TjVSWmxKLRMmIx2JeitXt5txg/RdBKi2X
xaAgQI1bD7IH2ncxJg9mUEoTLwJayGxJHzSFd//Oju9FjPtdl8ELs0sIOXY6
onUvSTvs9/RP8ygt3trYCRH+fCaah5/mYUHCV4X9rdL8QFlQbyO8xSJdo4wE
POHi7Duv+YahnYW3Q990qhrxjAOKhGejVhQilQBbYPby8Uw0u+lxYdtr7WI4
uZ7XDWKg1m0X2OAd/8WJ81nuTqSflnNnI7C7n1/eHksMPdl9fzJ6vfJomTXy
weh/fCXobnYM951yuaUzaK8Usqjj1AxXs22thVvX0Wr0QDP81zaTMme5BIGD
n7y+7JntYnzBkfLgN6bZE/wTj256TRknvA3Iw34GSg/FuuNi0/5EXM0sMng3
nX2o5F6D48VQk2vHbxI/q+LX8XzrjkR83xm+/GgLp3B0CvY0GT+DgvDeC7VL
FuX11tLSRo5m7QNHJpN4CEuQn4tZibHJXFavsYA8g7/yKZa7BdCGlXCBIBj2
sg4hdOEfgn1wfy4Y00ZSHMb9ZOOZ2q6OmgfwVBPWwH01QuLu8+l+fxemnuNf
SfoWkMndxEPiuHWsxJBMlXvvu9ud7QeZpwq1ObMp+ZXd+Z2fO3GJ+C7hzxZw
D61wusQ0t9/mbQiqnhEV/TNSVG9ehu4T78jE2BvJXZ3YGbGvq73oCATMi2E7
q6ms8hVuGghTOAOOq8WBxYe7Vo6/5A9CrJ9Se8lyNKcxwH6OEE0BgvVkQmwn
+f53m+/riKvjkGqV8ZNyjhULyRkrMbyBpMtDUjx3xTJwUuLWVFUO0m/v5ds+
9VlQkVN/cCwOuXhl978FYiPtdQXJVRa2h5Aos2dzkkU4MzgzPBt+BJwvRRre
QXlFNs2aG1pqKQMwWFr0vVUy9hJxD0rzb/QaQXYgiuDSmepbxws7HFssLekV
tBwVBzcDeYB2YpYR8QJmmHU7JvOwxA2oDoQ98VX/UIv4xG1iwUFEg26GhRn+
ZyylCsUWu3DTbqJF4y9f8D+pn74bJ+0BkrZUy/6kFyrYOu69jCl8tZJR8UnE
4v6bz3ujF9KIS0MkmwGh0Fm855WW06ZLvsyXdarMwfXnG1PVmH1mlYtFCAVz
eVYi/fVq7r6c5zQzoLk9iDYeqDuo1DnImhKzMbHHnw3OEwwVOaCXs8Ru0vsK
X0kCB8saWkMcNZJAB3VrYwac2n6G/qnmK32xFi4UEgXZDE5DZKMmXpfcpaOT
nLRvblFq8JnZDdTyBg8NlOUhI4LEhCcgR/alhDWmi72w/XoslHUs8kCZn4Rv
2t8on8816yCiURPckv2yABX/TrlNhccHXqBK/7d0sS7Ps1gR7hIrCIu3ezJf
8YBPBbWoIKjl/mVT/5KrTA1GwTiIwwv1JfFMOmYmL9HNC72vwLIPxbD4dS1g
AQfaMEZBYzmBXoN51xDvJQSn00L95NPO4jmKbXzoFeTq2Qr9Gg4cFWR/+gd5
KlN6yoMp5rnMe+lyI86N2fSv86HgHlEOrNcn4jmlIsw8sfCB8aHIq/RnUoDq
R6kB+Fu8lzP6OqKpemm3rp0UGwaZGZnKvCv5qu3ay6YEuV+N9XllPUp6trjL
m2SzRkOANZiO2wJzOEnXXOwVKrwOLtstZrN4UOlmrepyz3Yw0kXtlcY1axnk
b+OYDvHatK5I8LcaghydNY5d1jAVJQcZIuX0Mh38WVvYACHNTysCh69gJuki
/bInogvRX4RMO5EiRpxSCUDb7HxbslXxipCERzNpiWdWTBDe9ti8jmdfdppA
vEjOMZr1uqMIO+pfL8AC7d7PzqEaa04BzFDLe4S7JzE3dFGnTtCidPTRzKIE
QeFUdg1HyTVYXbLdshgFrj+eyKihssrN6aiTsd4v+LEGQASDvXVK9tq48WH5
E77FabeTBptwLANcIgeRmHaTFMf4Yr8rQEsKM7M+ZRGZ0kl2DptvWqCPl2rk
ee18W57R1lMbEtVZ2MdGAqiRNVXzbk5w9/VPLjI7Z4KMvRUDThsK+OR/9R1D
SjI9IOCnXa97IU2a/UQuk3KcNSxnk5W+7fClN3EUkil7X51ynw7s/DkKyvpu
K7ak/meLoDs+1Qs4rUZTaagZzAOtJSJ/SglARRpd5TsCPocvObotij7aQLPm
J6lbC8P7yzD56M3/zYh6mzechq3GDiZklFUMsprlRS1Thsz3Z5Fp82HViihz
x18BqjieyjEG2qzX+mVlapM/kkpShTUqu5mDEPRWdiuU5iyiHIW3YTlEt+o9
Dr7BcTTyguU8vWVsM3Sjx1E9vpG7vGKNS7hNnyfpvpOdJEJ1xKdN19pkke1v
PvbUY75FVzCdwSqXEPmNQnxxMaOCcTNZ6hqy8AIMKAr8W9J/8aEM0ngIk5t0
o9xEVhm2cWXGKer71137bQdtaJJyIgVlo/VsnPK66WFUjP+A8mnhCT5FL4YP
R9PDXZBdKozbGXZjiCvVec97YHx5kys/eN6+pLT+D2ap3isdTGu1tsGDjtoz
+IcWOW7O0r2pIU0bI0PXRFM/YWYIfkZTnaWop5CIVHpgvSH/Gd978/Gc+xF8
aWuG3s65KuIPHN5wMpa64abgm7c31FEVRT8ZTTQmu/qqHI8vZFDkRvTOWRKj
JWgtsOLxXpMjMX3u/ZbIU3Aw7FWJ9oxYsRXCn0aOeErhUTSbNsJma637AtI7
r3cCUIfgxETSTJazOR5n9eMbDMgmB4bifhta+N2u5loS383V6yGpBUAZin4Q
I+jiRigHYV672MG7mKtKoLzWwOEZxnSTc9z1U1fYYcMsA4uU6jooLIwkGQfx
xF2GgRjYpa98K/Z5yzdSu6gnitHF/1w/J7nOm0wZBWXB3n9l+ZpfGHc+5Ld0
NFIIVsVn5ZxogQauYtlZ6yiEwKqP2pUUDik7tUTbg9SgpMp5SMW2zV3zo/sN
Hf08risyXXOrsiD2ql4rwAcMFkqnPNaEVjKc39sNILYEKlDb1CV18i9Kf9DX
U8i54AsrBX0CEYOScTSPVBq0X5gOIG0f7gXtVHTrZElrU66fcpmdU1ZKvFhQ
lgmAeUBFhxcwIVfqOtPLbcJpq7ZNTPxtg4stecNDdZyImH92OvOMWpAUkMD3
+mcvZo/wmgz5bsVF1//VDp/4/hLJjzicPfuQrxRJjACld/oP6LpF+HiyDL03
OO7NelNcmLQIoTaUXH36QWagB7af1QHy3mkTJpb1UamnCikJcwnBbn/n5oYC
cUh5tt0qdrFwOqTuOhN6Ms04Q1uVk9JKjC2higp3A3d4x5LTuhub5HCc/UX8
9E5wjxqzo6xwEdGaSDYoY2yLC+uSAmpq0lRpaWVZ0QU7F2Ds9H/+2AWUURk4
QHKDfmZV7m40zjiz8AjHi4wE7AhK7gATjNYmVy0+3dnPQ69n9iVnEsVVt8S1
KzQbY9h5u/GNT+VMyY2sa/pXM8x9d1l2Z4c2rvyi8OYWbthMG4PVCLM5vNIR
Q9pLiJhiCKSCm9rICYY4XY8I5ikVTwbmVPWpz9VSsA2l/9KsC6aS85zhIqau
UFNbaQjdQUbIJscBzYqOdLfJxhempO3/d1DiThMEY6p7SpDvFCyu4spg3Lc1
6tzbQUg2V/TMhPX+hNyL9t4jj5e/wRK+J7ckH3Mg++mNtk3vicrRp05fgl3t
RuKYWFUc+AHNdpvu+LcNgE3SEy3kDegurgm93jxXpnQdwlc1JeqjaNscDWue
pAxSJ2aaRY3VCfD2NZPpukfBAel1kqmFTDZ22MpusVx08Lo6dTksq7IZWKL5
euQb+1HVnO2ABLhex2pAFG+Ukb0e3Yz4JAky8u/+xbVdL9gnJqM8p6wxp6ga
LHoBvQ641WqZWqDO5qzeCWvLPcD6QAf9vZUnvV2igyE4IbBvCvx0ek08qOKO
JMzTk3gBNKAjMtdacsMZFKIu7b4q5qz7KVQpzS+Hf/SYBp9AJ6rQJXfYX83h
2qHlwcdrIGj5ZXWABGLwUroQoyBdis2zpVBs3eVcnBXRhhJO9q7AYV1/Oem+
2O6dAneQ3fNMFFMiWGKHx5XOH1K3llsVyyxg1QwI0F7p/VgoZ5FO2VTP3TP0
y8g+cqI2nLwlNz2QBuXiNbUWP+iZqW7PT2k5rm1tq1+E5q0L48K1ELFgSLWA
Xtq4BBidR5Y8ZsdA8FwS5a3LYl8crgdLTJOMo07eygiTfZo4hioPojO2L2FI
7b19APJYrD6o3lchbJoQ8MTfOttE2IyLiTuKJHYDb0jYnYGtcFbXVRKA2eZI
LNZFiSAPGM+vaGNF/+ooD+szAdS4B+kJqNYN8oRxzGkbgUmAz9BKsgFDDstc
uKbPj/FhtyJNCH39BMjHniee3/JbfHhqlrg50EfawV8wsOlwvLVhJY2YebUo
dI1a/W74jV4I3HlAxFrhVLZpZR63P+AcMLRJE12SBlgny50OZPQMFOvknwO+
ScZGyozo4PvDIOTEGZz9gvwnNfnbyHGIhVoCFDl39h9+7WiWX/5AlFOFLmA5
/hMChAwcVjIT13ezdndZQISfCerS4YPXu/Mz0oyTcyVZc4jmxJ5zsWhXL7JF
m/qYkVeA4q2M2tl/5LYPJK3t1A09I/k/1sSiFr2UyJ9arEe7ewC/5ZN6UcSW
5oazyFfZjhzCLOIm4ZAuuz69UlGg0Lt1GNjMR1OuxGU/SuiJCPmIVvMo7cMs
5Hdl08sMsZ2WPPy+XBkCk8eHGLqfGcq7sAl1Xywknj4/GuD3edUdOT62lGdf
51KnKuRMF+KOOYsEDIjwz+pv1pWyIXmuGlhtM6LArBCL40pKxEGE2tAv9KHY
EU6i9+w3ff3KRmY3J5fP+xqrsV+n7bEk1eqIWrDBvtQReGBfTuqIIDlRlqNr
1aXAaCS2dXadFxyMjAVanBW1N1Ntt/lLMwn3CVhnFy7YpQ02GCHH4etWsCTL
dpQvc3XnmtYobkBHiRxJANzrktsculhsKeRrL46BT+uA4Kv0PLw4ATanjbdP
IJAsUtU//uYggIAhqVbB4zf5cUQd8hT4MerQ3G9kvSy9uOtA6aA8fEGR+3EQ
SFXefgUEDXFC52nYLSxhk1guJVKkHgb+OjCeIEPXKZzWnP291//qrcDsgSrQ
BuSLmXwIzoiqUhlzkBsFAApQZchMVgv00CmSZRxdg99hT3N8oqrUuI52ykdV
Pq/Lsm1qiieJz3ocrf51P5KJcevNhZidN3zT5jcuErxEpWhdtUJkIK8BfM1O
E0bCcqvDQy/ZMcPRbBjKj+riISB6ZFC3TC8CZ/7s85V1wN8aOn6WJPzEMXOn
2XNx/3hEfXA/FnbRGMTNbxcKYVk0GEd7xcZCo3aDq1AS+/0U9KADgLCyKPyP
ws1r+EJwwnJdofSiXXnRRci6qzf2F5lvtOrT/HUcHZMiMHFOWdPzmnLfF/5b
GP9jYDDZlDPRsdnUfMk/Ejb+TJrSSwlSM+VFOo+Ut7JC3/3bvPGW/e36Hb2J
+htIhOy7CjnXDKz9pPFq94DMZlvf7GcgBC0cv61wm7uDPMk+oVtu0+o1TeCW
1HGkUc+jzySmVOHCaKpaCiqGnzpdMiKHvyZZJErvvpiaCKVHR8gUCQCABKst
OxP+nxDtmvpouU0SS8BIIwhxzTBW0LvmVBGTN8qV50YQL1Sizc8dzUc2xPN4
9SQ3glglJ6eld4ZtlalRjKPWvajNOG9Ywpbld4YdRscZWySD7tGckFZTDV33
CoWlYwC/y/fnGwtoWfr3NLb3K0uU8/xFLBL9atsTi+1rAGC523+2tFqhnj5/
GFj1bd0AoWurQtLvvO7vmsi4psfCkqmRKnJ5VJmLmqbOLzLtqxcLN0XW+Uy2
1CGU1Y/YhpqJs+EOJnj0yMbJtBLatPFfFWN7qQPNHusPWmskqgAgfZ5O7wZd
gp5Yj8aQxUJ4++nS8eQWaaEd/8HMC2xtQ91qRof5phuwGys/2nL9QF0HN0oQ
ti6NxllCf/wOLTC7WK+xGN/srdNq+qfDXAU13O/jV2FvZraVl9dZ+E79Kcp0
oIydFmgWjtErVJjWc1Fs1rtngyuM/egkiJGaGmLC06n/A+KOmX63Kt+ZIYq0
bSfEmExXrwiKOr8pPC8YoPCI0FEWPmRpQs5iIz3LGOLjBv0Net8bbOYzDUdG
LT43fKLxmdnKkcDjvY0PynAG9gS3mwmQ9521RvCxmwbrtxN80+AO1ewGUGJB
NvUnlpQBTi1O3bgkBq4GRuUAvFz2uhEqfEPOD1xgmmIWFtbmG6kP8xON6rPo
zZJgsVTKnVFdG2Fwehp9qWepMXW0DOBkHHc7A6t+UN/VY/OYf0ThIK27axIX
pQqZr4SOtI29z7Prq/Bi3K1J1uI1EIIolyMKvZtN/crJIXCw4MZkI3DEJumq
LzRJANTkJUiB31HSI1B/nL1yPoY1/i63QyWx5L6dfmiLe4q8MQA+s6m0YF9x
cd0tCFkp538SVYM6hWHYfshWjA+BAj7FBRH0Pp7/HLWJi9lxeVTXva+b80xt
XLnuSj6w/FK1sI+Ovw2odRcjKBoF4bGM/0bygcyf6R8i2gKbfFZHvANHUlPx
y0Kme4aR10+QExRSTiMwceXY64Bq6fSNO2SoBcbawnMzfhjVYEQonGjz2e2o
6kaUlMJegREqVVnzWK9bEOaywF/5UQ+2tFIHCwHVbl2yBeLZy7He0xgkS2M+
IVcA2M/dj86gGWXTvAif5WCGZ0iWIXmTrvA8CEYlOGdeYbUfz+w3PqTpl4fd
6ggE4jz0fsviz3ETP00Qs9YZTbK9RZ7Blmw0yF4lBb/u9T8xFUxdZgh7Q9gD
nZsnqAeWBrdlSqkCqfYMVfVZR6Hyna50MGvNBfKqfqzVP38QXpph1zLaELk5
nRhPZM/70mHqdE6SrPyZil5vsv9WBHTtgb7oUSjjbVHmrApuYXoxpcXjcO/3
Z0ZGZ3qTGGTtYL8XGOiKcFeuAmZGGlFbs5r2RX7EXy8a942WBbJJsjIWrsur
QaK7xKY0I+LbLV5fc9rV7yFNfRiCP/0oms+E/sJLMLJrWTaYEq17YeBLaUTD
SpqTj4tlPhWSwlaFKJEM4SKmDLb2ajZ7/nO+ao0nxplG5K07uarLI11UExSQ
1DjqeIwvop2YnDVUlM+uI+zeKh2Sibrq2UnOSnyvFKLMnOxSXOi+Q0WCSzQi
DR+wjQuf/5OuTxlVTrvNKV8nXNP520eX9TaPJc0LYmb/MhXW0v++ED9pJrnH
jhO9d9DkEIS+UtoQHG37I+tb8+45w+3x6gm3exQ+6Rr4AbUDkEH09di87ol8
jlWM0SEHWU7Y5UEJTm5z82KODLFIbz1k6iSokTr2KWuPJSpHuzgunVTNixNz
ZCnd/+EIJwBP9ttYznBFhUb42vSKuTZdVufGgVF/GiWKkyHhxuJSNhZEYYp9
C0jOHZMjscWoqqytvcY4TwUikcAJrSjkmX1OQZZfm49XJaDnlEBG3u3C8lJ1
0sed2Fx8iu9F2WsoIg2D+/RgcVKUXVzFj9Xb9BkYpWQaBlIU0J5+8Ze3ReMZ
LKXF1Ivh922vVYZfgEybitKjowIEaTWU5QeCjaM/OPoCykzhNWFdPJPXaMvL
VVIZzhDeTb2Lki8XYyadNW395TcI0yvk67TCDNkD4LTAGfDin9xnIx1ENrGH
tBhh354B0viV6gsPdmvHBYD9EXoG9fRKhFOjksUuC6isBmYFy/5M3wtegOyD
ZhSCs/aCUllr0aNqaNu0KlZ1wPyOAnn2j/Loe0f1sCU3zFJyv18koifZCdUZ
L/OLEsshqZS2RxGW77ryv5/vH2VsNfAPQzFx4ipFJ9PkI3/+qiKuIzMc5130
30nI2U1ihBrEDORiSkM3kpg9GafzOUmZA/3mnuwgBwq3D6gct9gNPSARkg5C
sfVnH+M6QM8lpxE/zsAxmuIAx08cCUwa000rFkFygj2Tll0ipG+NkpofF8Xo
iyyMwxViFSrhc1KYgHyPiBl0VSmh1PY0mPhjXKwM7YstlpmeIttHPzzAVpAE
Qs6or1ijZTfBW5Ub2ELdW6y2kPcpMj8tbrBl5DpplWR1w0fBHp7xVZf5/Bhw
zzRKVMdrjSwF3SYVk3oTiedr+A3q5gsaadi9lpfF07pPQa0BkQY1TRZ9l2Pv
/gPk+kpl5a25utTxbCd591gZzM+6UaCpAWtdBEKcBvemUVQpFdPwKuFIZ17L
4oN50VRXE5Irm9CeN39Fidke1UVXlm4ivEwEuOCv4XD5b2Vd2LWzYNjTGR7m
kFHJqctH7ci4vharN3f46lnM8L27+fzhax1T6euG2Np5nLa+NlY/TpZIy8rr
kfjnDCjcsuCEVa2X/kqrGPhyc6rvBsiHPCiZfBV6R0zBePCGTnKRcGVWRi+a
IwdpbSy/NT5jRCCkVfiw1O6F/n/6nNwAVo8jT/Tie3+D0ZLILicCegUBJ9Y+
qA/h8ty88tf1kgxMlCbGLniCGU9XoXMGrpId7iaOwCO3XIyY80h0g1aROPoD
sKanGs8sYhIRUrnkdlrETef6PL6OFHqEWnTrSRDgsxYu42heGAbn/Fx7v/iU
ugNoto0ULjzwbhhNKavPsjimw4oe5cXD6dBQCe3V/QQ6YKM68I7zobpVKGEs
7L6nqe0B6Wx1GWcDe54vyJaNMEqJXEz0D/14pIGUW1ebYTObFPtBoPopzxtb
Bo+wLqRvqY3aI7HqiyuATQ3UMI0kvSD7rZRUBUJfWvDKTZNdEI5cWXwLSdmf
5l0r4oE5CssBeH/QD4DsDv5fiN3D/z1orfntQU0DIkdFNcw3idOoAmxGuu9i
rFOf4XT4MSo9S/bLGxEqzRHNm6N4ayTAwUrD0kMZuTyP5JJv9VSCzDMXNI9u
kCcPl2Qe/6sWXfj//KspDHCm78rG7aw6Ohs32N4h/R8YTOQePn0MUNtDJbMX
333wMYteL7wmM7AhIFKt50rRVAOPRc7iRyVPv7jpT1S7pu5fQoq8KPW8CmAF
6nhJLcot+pK1ZHD/50tH/x0v4hHDowlc9NDcsB+MAJn+r6wCObuCF4P6Wox2
CM9mfUVRPXtDLfmeCz01bBu0ynrleigaR09lw5ErkgM4CMY7kegmmDHjjeSf
d18vZaasPq8kDJU1eX9OfznE/ZQc2ErrC/cqL2Kxx3XsXAh1QFXnGmNs3i2E
986+mS77DEVzEAeSbo+wT17F90/xsTGOVV7dyLz+I3T9VS9z4jNHxwhajjFS
9Us4WAFHPiqfLlsBzfX+EVYGBZ1FZed+JaiwNE6wJgsawfuvuCDr43NqTWo2
+QqguOjKrith7WN5C9v+n+PPV71gqScoXdq9RSrkNe4IF3zjzSv49fIX3pAB
+cxqOJpn7pg3Oycvb6SUgynypcdYGhInDBtDdZ7hf2QQyY71EyTczQxSumUw
ML8wAvljZnrSnULS1AoytlGDZjRARCK6iZ8shppnn0yyFgx4fS+FmRjWhFcT
phm/q0LcloOjRK7VP+X0+/fdaFXLsJ53Rk5crdyotwR8PJ53saXc/fz0ZZyr
RxXkFEjz4t73CTJ35Xj8HL1obyVfoSpIlEO762+4F6dVQBxb58L1vpmNRMf5
r215b+gNg2qfsKNLp7BKVTzhDKPrnArhvdN0M0BCHpKyeyXcFkvnaPllI8DT
af2AC6iuawf2q/aAkliaLsABmyxs2Nk/kDMrCWSjWm3JAg9s+AgMxxXle1sM
nXZrUFK0tpy4iY63zA991wN1ALawK5C6nKRAB7LKZacdgrNKfyD0FYHdpFOr
dnw8odimH6HfCG+WKatEEpDU3yw29Kd0t++62ss7EGqoPd0C+Jg3nsbpdq9K
ik+dtPOWNHCvC2w/GqA3yOyCEvYYXYPmgtwIOHkAqzCitKAzt2lQV6aJxHfz
3VJ2dtrLwMO/kswyZbxyYwqPLFWYPmJJupVINvYIhCmfWr9h5wxYSrTz6KXy
Tx3kG8Z9odXigcWwRab3vAjEcf2aJZmjZTI5vY2xdvO/Mh38tvBeTBXRZMkr
9gxGVtScNDnzq+Fy5bJFBWLddI3GgXZZUYeYa6f+yRSv23ESkKkpZ4HVBeoP
PIN4YAJCCdwhzz1IAO44A7ruxygvhpV5+q8zAr9aem8mUxlbHXQccZomhnpE
mZeEiBldoGJeNfDTiGyU54iwuHHsE+W3qjDJhgIOQwtWEYzwgw/wRcxWMt4N
qtG9xjCfryjyWViH5g//uY2ZKQ3UB19JzdP2AecxFhHmFoS89ig+K/uKMtm7
NJNe68vpYiqCp8BwtgPDL2uvhu9Zb598EeX6PUnMWni/oKjraly8y1njmGuS
6K3jsSjCm1aXO1dBIwcNf7DQdmWCyJJeNTYl3WAOlwKOznKJ/OQ3+7O2D5sl
mhOepqRboKn1z67L0AaUuu3kgyq5Hi4hPTGzYKheFPR5CtATOQasMj429DH0
eV78a/znclB7gid+VoTvTUYgrnmPjiQSdPuHITzJ9RJmo00nU/E07US31LBm
PZOGY86kTBUUxUwOzoxs/LmIAhQnBt65oZQwoqe4HYDE8lQgd3y+w1PtXZx6
HQtqI80LVG8bH9obZcZul06Y+vPP/mzt4FW9FMQhEfyHOjzL6LxqCKv0m7/M
yq/mkfCWcCuzAuCD8Nr7DsYpyxJnZhpOx1TvqZlW4uzfdXnCzHR0Wyf/4QJ3
3pMJiuxzH5c5if3CE6LSLUmhDDtOSKAV8Gj7MDU4juPVNdfZ+K6nS94Jk4+n
Q146dnveVo+fwoBD7z+miLwV8qvODikI2mOGAaH8oWvPmch3/Mlg3/15amU7
FtmbGm+BeeI5DA/1dhXLfWp4Ia8ZhXYWrg0u6qktcPpJOK4pdM6+RdAof8EH
nTr6pKD2NM62p8dkebE/R91yftrxMG2tyLOUfyF5RMeZi0+RFPIeKJkt7IPT
nRW09u5A7ggOEZdvy5DKMVhrWKwghjdldgJHqTiR8Di28HJ4OFZG2aXzn93B
9+KbJEu8waZWD8kfqcnKnc2XB8W1lhjfCZbkpk8GwZE1TXW1bRKR63zKjBAq
IiDi0M97eYPl6OOEdbt0lmUgbUVuBgnXA8UEW0X6b0HGKAgilzaVoyYnBy7P
D/wlnI79wrDQnalNApp8rvsLueO7TsYo4CI0vatY57vZ95A+CZyuhbltgZUf
vp/jj3HlKzXOmK20mBRKrHM5XknboOKhD+5IgFfXYL+8GJaVttoLWH8Txy84
VH1QkHYXoqW15a3uiHi7tSAGojkqZNNoMBuL+qvgfEEtnJP+QdaZLzYtzMsb
7p1Me1U+BFEAlksrf+4sNR4QkGEBPSHrju5yF0O50TAJ90zh3uOzxI65jeWD
8ls8sHLZgMPjCdS8wWxCRszeXZtUHvJz8emmtGe4NOKTimlsSEZP/HwnPuxd
bEYSeSV4WZ+Cf9/eZnKLnJtFOXBM/r4qDIjSeHpX6R/dmvNX/8IAeZJO5zdG
ypQcvaLU/0X1v4dxgFCmPNm/YmU+PFrioGeylQ1SukbCWigmMDDFbfj5pYhK
+fgTM6ymXvg//RkOybVso5EQ8uk5NVRG1BA7pfoU3TcN5YpY6GigLHUTEWNM
mwIBcKwYcCvOgmlIAfWe4luwPI7V52anOwSuYLuvRRl2glTABxffJcdoxIJ8
piMpbTN3jLfO0e5TIOJM+Y5h0wSVC16EBgxotgzDoi2K1Ocazxh6nbvnJzy1
p53UchwyLrGBASuGpXPDtOKSW6Z9RuQ58m2aLmoqv+qO/XTxs2yrPkjcfO+p
1nJoxLJQrOxVlaEBqDRqOvsi242dVDuKyIxzY5Ru+SNAVU9cmUcly1hCGxdf
eStwNK5Fqtat0JTMG9rnBCBL2i6fotw5PVlQIpG5cQo8ulZFKR5PM3xlIpY3
Ti3MYwLKrdIRY4on+Echn3BcqJkKZHd24b3adywNFkZLPpKrZFsKT+uz/TmR
GuSmE+lhcYOS0FmYb/3k71xaJX/a2R1Dmj2qXrpwgeSqnw6kqQIfsUd7wqiH
I4U9Yc1iAubOzI8rWhezJKT/oxwlOj6Ed/WPKftZ+I8tMhZ7l5AeXebpIkKK
JCKuzFm5OPram2kOA2kfTwBBEyT7bLYrGOTj5bhDaTBguw4mMCoSrPiSVvxL
FQsB6m90xZwpqvOjwWfVdVuW2iIyJ/WvI7wSwdt01psBPnR+g6CyuCO9gOfN
1Lsto/83HgkbQf9ZSuL6LHXchKSqWpo4s7qqzBfVVtkBnBTWqZflE1ka/3SQ
Gfn96K6MbH2Gwe98XOBax4/k4dKyjbWTTpqfGNL0wW9PgrpaOrWcqHskBd36
Yv2n+fAJfHDIzS+Y3l7DkznBTVPGPCZbtYgOl4L3s7xEg0Y7B5fF62yx4oC8
ukq+KxziqFGnr0ttKqAnNP1M6/isZ2riY0VmEuiW8+1sMsTbuBTiQ8R7PJGV
7kiZKIMUtf6nrr17I6ZOb4VqxKwOLiOghliLQRv3rZTEzJNbmLkNFgX71p2J
WLwSXSUY0m2frUxXc04BQi92pwy4vwLyG+CUjLJuQLPpTvvmziDv7UkU3+O2
t8ev8jgJhI6ABm9lYjAj2zKdaYRwqsuq51DhXcTFQPV2Q7UJhDgwX8Ow8Xzd
CLzle+sqwJLN4/z4ZdzfAicgy1vibfrMmk5abffPUEmtfdBEXF6Rb+udiAeV
ZoVqcaKHrqhg/YLgzLIVhxDYHavpKVQVZ5K33vevbSRTLek/2ZG2kO7OINHa
DLgqyr6NfHpND24xkMZWd/K8zaFhOK6LwGxrCIvA0qfIvP1p3v5od48hKJE0
KjQBB3pk+7YjOhTKekVJvB7K2/yB4p7t83l5V5UBn1moo66vpmzgyLhB4ddS
IceDHAzztucuIIolb5bizcf8fdmYyc6Md3X/x/bb+D9JKcj2Oz/jUdacPSrR
aMPL2+vRzatojxaUELQkShTZrAdm11w5NwVq76QFUzhjGGKh9NZUmxWZFksl
XikDu4o3WAeNh0s01+FXueV9ccnxGMKXH0yddN+ZfAptVQ0FGgNPvraNJfTw
57xtWUbueyvw/Jey0oWJ7s3IcYXMJp+XyxZDZwdALAiYc4a7+4VnPD/qbNXu
Ibj+q+s8cly9OQ4Wl7AHUkeYkMugsQf0Pp/G4whWDEdPydseAkFMXx4YHwrV
NE04b83oV5IQwskZ9bNzwEx8EClmyazA8JfLOnh0ZvBJdJ9Io/vP5C+MY47r
xkwTxDzZb7wxbe+wPHq5B1tznz6oztBR8kbc7CLR/KEuItU1hO1f5tcBwsrL
NjHlcnPEORX+QFYN41pTKXVDyVpYjqGIWJBWJZ3+v0reh3A2lnqdE9jsTtyf
M/BsL5VvHj21GkcK96bv79fXjy7QLutI4ol8sg85LPKgQDW1MUXVTrD5lhoo
KnJlL+lSlX/LYGyS2NQzgzTpu+Tx8sYp0n/qRJD6hbww2smGpSYOR98aHqYf
+jiHixZCCqGtMJT0AClSmn1jiB94rXhFqCov2tJQL63e8Tzo1ND9iI/uF2Ei
pgDnnnA4QM3WDAdLx0ptmWgO/sOHAK/MfbQNDuoftRgl5I3mf6lTPYTKZaml
bR9QoTAJjc2/RBDj9kkNGLDrLwtpohbAVksMoJPWltUs5mZ35bUr2xHrA5Dy
omfnWV+dKUew3UsC2bDut9w14mBLA+WITaqPr1dSa131aLIFw/JJHeirKmKl
4Vv3qT32IFaIFej3RADbCoSg5SVop5je7aLIfj7uKI2q2z9iWfM8SiX/bfbz
2qvJNn32J96qQENTlJT2RUQd7XODmHGGzSlgOf7sw8CnING1L6smwbcH/cED
EUEOlicJ0xQa7x4qL944UrWm+d7fjn/djt6sjRYp9MJeQp03uCokH6gxRdsh
qVoazS87Nzv0fA62VN2aKxh4HnDEcG9Lvr7P+dvjzpMNNI/zh2V9p07Uc5JB
G2ZRRa3HF/TIjlmislkb4iMR+tghKUOe6IS4ar6RkWGDf98A/pITQROWxpTz
JgfqcUEbPOrSALrJyRZNYvgOct6fI1lR5TPC7XSIcN2uQAWkcwNdWopXiRTX
FKYVL/EeGAKY88v+jJHPv8B33nCvjSLkm3Nc8qoDnlFUvuENizWGwUQHvtl6
S/kf41JszBY+8fQmf0Qd+6ueDaZcM53cWJv18qxBk453j1v+DnyJ6SGMZDeR
UQ8gSQxv8ksAAnOsptZ+FkwuaYDAz7Csj8yElKXWWuN6JMFa7S+oTuqhCQ1n
hbYeYOf7EUte+DC27YYyBTk6ySpeHdVPGdOO/hR1EusLxC5FKEqFb/lUhLgo
KeDCWLCM/atzFrMTfN2wXqOAVOfxmdDTEHTOODjW7Cu5iYpHmdp/C7VWMlCv
lYepcz/HrS1fHK/p3eEOf2zStfetOHhvVO5ahBlfcq6NGo6Yn2XdmUwum8to
H+yRWTkAIABjNkzZG2uJ/v7p0kFZwRds7Jd1mAgbtKtUXtEl5LHJouRYwXI3
5Yj7lh9mhIoZ0VfRUIS+/OxEIYx7dzWhKTPt559kwTWzy6ioNMcKmlhHj230
1W9rXj61x0bIompYuEg6aJaPEAKPunhJMUhaqvbQH4SW1SBr1xa9b/2Ga2Iz
uwPqMHZtvfAgo7aP+YXtvI5YS4l5tyP/WJ0GzXg6zoqRaJqthkVxUTf7s/Nt
quI+Zk72/SmRDjAG/kW0KnI7nMx1zvHvFjBTk8qiGFcOJfT4LNuK1zVhCWQb
9JIrpKRBZzu2EqKzq4Whgd8RiWfjNWCQhJHfVuzmmhiCSXTew8/ay4dyVUvD
vg4rpEpB8ZBGhU33hmGYssbxL2RfN+GePhuC5+RNw821dAxRTs/XTKALBgSi
qCY+j3Q6yYZZg6OfGXWUoLCbj2Ij2+2pIul1oPprBTitPIkM35SGDs6W2/nv
qNENACNELiG0Hzhoa29hRB9SJoq+NA0EFYnMf9asbNw9GgSnjKlySD+Bsf4R
QCC2zWsdNmVDpjZ6CrdxQYnIid9FV9LGkmbMypCfeMWjyz2nV8PoGwPq7eam
uQgQnuIqML3ke8RrYXFaPiVeYxLVFChDXlCyjnb7mzHf0Zs7AKCShGuzZw39
vTbcu4Ep2cRtcGz4jSQqeX8Px6jlExMw0ZPQvRxPsQgpouiszvaiLCjMN0MA
9BdacZVMdGPgnwzQK8mNmHPv9NIMKYcNrzRDCtRIdthM6N9ONchS2DbqYCo2
QDdUy6s6Q/jo8/6p1lZNFORqYKuOyS5Un4oSx9yWspwbZX9PkCrUQTEKM5Wj
md9rXpr3pXxSPWY6zx1dxKOVAkXUkjlcF/eNmUrlojhhMlAtk/roubObGWef
watPMOAC7qGCnXwwLdobeTwEyr8scLUY3tiANwjso19WxCo1nZLubfmJR7AG
qscObNAkDg3kBlxsGuIhRag+pMVaPhPPgKvrjQDSNE7o+ptQQQRnPW02pxdl
ZRYlbNb/N+Lkt0VYq7iQMJPLUoIb/R+6Dm245R8KZjJ4+LnMmvrmTV0G/gjz
Tm0X7m/0bptF6vbCC4GDLeGInR+vuaI14601v8MTvNxu40lDgAFWCppsO6aQ
Cw0CVmX5ixeog4/SaBzHhZtdzpllXkgFbV+q61Sf3NSYUcob8Pq1pUXtcmwj
FfCWrlF9sbOtkaB9hRERrmRnanFdlDsNL5wlswJG8MB25JLgW6im3hnPotPC
hmwUl6/5Y1foJkeUAXuNxvB88qeG+LQEc4bmG4jeZj9RA4sX3/DuAKeNHQIm
C29xfBJNh9s8JfDQrHrUr9s7bKAApaYz8ew2+G25qgbev3Ctpo7X8wK/9itQ
WHIeCJ/olyW3e50Bk5IpRAHhHS5IJMS37Jo9iNLT/aEBY8p8D1QNcGHGMxem
Q76WCE10zQIlhUZ/NooCUVzEq0DCOSKe0LboDpaCGweG6LJiGg+5z/wrTqFc
raItbSZfuXZ1/QdjD5yqWN4j2+rxyqAIpXnzR91hC1u34HWlDK39ij7e26BD
h6JTwGu/wIIiTRovW7RoCmUWpeE+4UlC7ZBvdmX0Gss43hZtet/rWSdfNEHF
MgRpCay9IEO773Pl0m0M3Fm9wWMai09lFw5KKG0HzzcHWrBGqEvpU4JKef1Q
UjZUyNhpQ9ujNzRf1ZoS/x++n2TtR4khOqjxTt90FDO0WtJ4md+XIneG9PfH
VPc5bC4q+1OQClmn+O5RLfHSqpzMxeLGUWS4vAczqEhaWbXlZX6Rz0nipsnL
Go1jsbnUOJJu666YeajvEnpQkqLx26ZYfm4jonymHga/Lk9lPCs3Dn20E6Ox
X6aJc4Xt8Vr8Rtfb2SW1IVgXObdvSLAX41izcjb2Sra/2CpMBVcB8h5Z+gjK
3RMp62QDZlskBrHZbO0duZzbDNYRHGwkpR66syXQhb9LT4RohbM4gEEQtNJG
oFLB+JtZDC9mc52Ki2hepdAvKOGJLTo8qzgQ1mQ7GbP5liKc8zKx8uCpNDqe
Qp8P5O+9DnhtMNV6nU/bxUWIdZTzx/iFymqz8uVmlM9kysO3CK82NqVlEY2N
KG3x3x97qqU3nnPCe9nUygKSQKICWkSzsJuNGM7eYqMpDHA0w1wmEy9jywd4
XiAo6DJNrSE+Y2cfrbNYaobrjlPZRZwZmUASM4EjwqvIf7SZBKrkiDhqCwKK
eM3UW9kL6dsVtRnZrag1fcIhKUyFcj63iuDOfvV1AvYhw4Yn4hMJcMpZ4hI2
uMbcTULkzlOX0Ul16oI/MZTfsmXhHN3zDLeE0juVAbJQQDdPtI70xq/IIrUw
plZ/kSuc/1JVmIuCZlUJWIjmkTAU5f9zvvstthu5sYIVlRBAKCU30eXlRib9
ifZxlB3YyiF/peXYJuMPypElR2R/Drrgv4zrLy788g5ZsQ1vgaZXBESmXott
dAM+Gmo37JJ2r0AQASaSCyPCu0Sj88Jllz/KdN0D99+VbgJiafVmvZkxVFvu
Qz9VnHfN3gjcR8dOpvQO0Atmoqa9aKnm96+4rlbCx9Zdu8hvSNk7ezX7/VT0
AptAGOGK+YoM+57J3LhNp5q39nHu2xkoZWP8OVdIvZLZY8qsGpaywHTzN6/q
AGxFT3ZrZHHbKnPyNC/SfaODJkXIPg10uP1mZsmo8Uev2JVh1/uSqZfn7GTj
gqOw3YMoRvtvO52iiF/zVaMLS6G2LVI4c356kRcRSpXf8/paJsrw7VAfO4CD
lMmxmCjLcmGVHMijpDUvvHfkk4wRyej6rqRNsE0hwDXNoUIBimFropMWzjgp
FF22qujX52F9NkOrVGvPA5hBJwVpIEiB70MUlYuwItz6Ws2/QfTXJWNId+P5
jnDntjv7Kxsd1XcEcC2AiyTSzrOkBoqgPpUfTi8YmKl6RyPOqns5+tVQKKYY
zTfi5BoIwASmykcdFlSuuRn2O0IX9eVRoiEY8GxwJouuz6efy+ujJyRwzQWS
V0HT6euK4hOFmRk3crGgEZOg6LkezeV28CH4TxNBWNmMNPy0RtaCr5lVQv01
fkCBfdVbjIgc4tLRJfYhSVBl17VJFegdtqoDZsS4Ka/wyBhwVNts4C+AFGqC
hAAw359yEytmP3Kp0zURfS7nQoTjx+P60dwtZfV0KHz8IvJbcrS1GhHkq4ek
GP6fOe1uwYR1NktnZhNBK4jNlM2hx2XJERzuPf0esyXgNpVKqSGGqCCVq2pN
GatJo3G0Xnd1bY/fBSsIik5oWa2Ood1Z4s0gBZO+Ad1ZquBsogriXW75jkSy
LMEbkEDfIsU+g0uHPZnCMAJsWKueJ7QPGouGPPyoR3KA2tevk1deOPGXLKu4
Y6onaUuBtUy3epgIyjHZu/3g+me8/gMMZDSTE6Pm5O5YrTRYRxg2Chuvtvbc
zVr3Qscm1wyV7nqP0KDJhATg6cpGYU/9kPY5KNPzfitRIUdKDo3cMP9p6IWF
E7VcwdUMu4B5xI6H/+afjSYcKOMDYsuHzn/TO8qVyOpOT9YlojNS5cNOwV9i
OwNIwTYICoLQ4+r9WH3seSO6vP/ftawbiiEq6xs2gWzwwfNrqGZXd40qAe+g
elh0elJn3xQbS27vPQ8oTEhCo4KGr8+tJUp8/6vMraR8cL0dPvlIdm9+qYN8
YO11DUG4pWv4jFI/AMytzH9HeX6gfplkoOBwGZGznOFbsmKSpZprmbBE2r59
OLqXsR/hIIBPPvHRgc/EAnXHoWhkXfbfCh8XI+9o3RHH+fWvUtY8yTb865PA
Tc1y+KLUQ6JkmFUPezurN1oRjlk3A6qEDflYrh0W0p+h/ngQw9UnFcVQvrwG
gspZKDmgbTweb1hHbsD9CYtiPEHeQtHYyvrr3W1IlxI1HHsCR/untjEFPoAY
5BKCmBcMBuVM6kXh2nS8p1+Fhp13GDYhTmCVvWp5YokfSIVBetjLpvAQ20LF
ayNXhl0jbJEvTXCJZql2R45Hs0lzLKSV93sUvqwIVGjUr95KGUgirfOzwR8s
fmdeLOAYq26rMQJT4DM6Ah7UOLcLaKdoCpCoLdAD0s+J7dvp7pMdwU1Fcr8N
wuxC7EfGgQxFspUyUDB7NO7dveE4wLtSFa+rrCyYSyaWfzkF0oJ/9+SMbEtm
SdSWA41It+j3ej0p90wVvJ6x/jnixmEPIL90vf9477ZC31HsNgRVezzAFeb1
0KxfEymKZu3BxEeU0yjRwCJbXGKLml6CstsVgCnAvziKGeGJOSQ6XQoSgGFl
FbpII+O36hZjOwp+u64KSLbzJALX7AJzWOwOJVF3TRkTFLNou0hDjNofXqiR
Etq1gRNwx6k+kmiPy0tJems4YYqPv5co/ZX/Jjt6ZkRJF4TiGGwHNS84/5EF
t9hU7Ol1OEEF7U96ubzXm7m1hD5XY69YmlsCwOh7yS1bFf4vQ+37qtkYmys7
MECDe+Who82U9+OkGLJ6jiZcKCVB5HVv5y+cd55ETm0jCKztTISHzg2p5f8P
aKWFxUWyUwa0t5mdjC58+PVp7XHKbl8TMKuK2n4llT30mfdV1nSqjUXS6GF5
JFiscUlxwOfa3gobriU0bPcLPSh0+smvAHwwC4YoMMCapbIpoc4h6xofn52B
Sjd1sRdQIrcPq5UZEBaaeQhHdD7+YhTzOL0702cfJGWeNFiMAYo0jz11YuC/
mcHIlhpsNVicBAR1hY1V52NnUaSEicW7GFtaOglnGpJlNO68F56VQtN64cKZ
pAH2GSLm0R986+RixiiMtyUfQ8LoONgx/co2Q8GngJUZpC9/QLIofX2oLQcb
tKJ0A5UVgPr7Be/ni02vJNGnQO+i2yZFkzukafceegAIMNfNCmaGMbXIxvDS
C7O5dJgB2G/2dqwCigIb4wF/xL77Mb5/l48b9+qSKMPbxrFeP/sGbcFW/bbD
wMaIGW8FTPnsa/lW7IiATKpGtdEwSY5XZbAgrbIKD/Mz8hkItC82D6jgT0px
3AZNkykkQv92mO2XCmlFP95bdQPqKAgUqN7VIq0UD50WtNE0R7kPNxYKDE3G
aKQQ7+/fqOtDCXBwydBpSmpbBaQqCPOAcYp97yEn7VcDE6Pn1DUCEIueDqu6
jZ3t2pb0sshkQm8Bs0g5rego0ch2NahKWGZ7k68pzJ1es++2eN8DTRwB5Zo0
waqchRMArQ0B7iYcKMG8B6Xf9T446vo5rOjKYPdvrsgiuMn+2PKlbrLlQkG+
zs2tcbWy55wJw9KpyBLlCnkh1qHchuZZ5dsRKUo5/dYyF6qVGOtgy1fjl4bJ
BrjdqC2HjN4pYrJCk3e7er5IEkqAcLPXvxxAYGPTIR5VEwi5FdA95WIfygqO
0lpJMiv0GtcxDacZx/Zmeb7tWBvukoR2f4szBvHLGrseL4H17YbHqBrWx+mV
/Xa3mVb87D1aZ2Ooxc6I/qpvEu2qr6IwunZoow1mWasXg3FbsYLAPBoCfLvY
H9JCehtVQaK6Dg7Y76VfGRPvrmwUNQ7vSFAWxoOsjWfhfWhAzSiJlcIC74Qa
Wm9Fyh50zzuSJfTXg5jwIIABH/cZgFcKHPQk9hBvxMEY64hEwEX+KerqNPfE
MxLtj89Gb32j4ygjNcRssbD+w9u0m1KvTBtvi0apJ12symwborjTBSeCYdlF
jyL/aRnIqEUVBEWBETCNE5OCGQMaj3YV2hI4yVwYBHTjcBCVdJl0S6/GFVYn
mCdMOj8tqjFRP1psOuTqHR3lMT1bXmW3SLdd1cI3t22Fmmkp2lq2BZhdSm7R
NopAVuvsaTaezJm+rcD069dfZ7Pt6yGSEf5F39a9hU7lIcnx0BtnmesekI4y
7wjgWlIt+MNtJ/IDfWkDRQcghW+i7fbhPnq+TkrIznPiONWQMVzQUriRrI+2
zTQU+Cs5fL0dz11i71q1iWvCvGg4liTNBxn6B9aof9feFsv/SrDBzCXxwtcY
q4gOF/6PQeuyiEFOVLrRo0TXK9kO/soztJhzQkd+Sg/heCNZZBDbGFiTBb15
z2MrqU1bUjDjm+feui20T+wnXrM/2+laBf3OhK6h4O2m+32xfbnTlAGxpDKS
lQ+40ZjbbCf/ssVExmw9OEeDPIFT25Zoyay17XadckLQE3rKSRP0IQFmk4VW
e7iw3wrno07WE3wrM1wb3NtzV80oGeRYz/Oc1oSvljDe7nCk1IWD4P4XT79a
SICjoaiOXE7lOqGV+bQp6L/mrnjlW7nEn7SmwTEpsCp0OiPXonWGPMUc5x6d
snixcy+uQV3uf6hJOjs4wI3fLduqI7IATX5ba4iFFMho4WNSHjolFd1IzB4+
5A+6ze6XYuY6hUQH/wcDCNI3H2tQV6ealhHTF938U/DBVggNU/f+bjQlJxLQ
x3wwF9ImIjjqmLBMKedYH5OlYnAcLSraVKtELHN+3CFzo2bNi4sGasmNPx2T
Ji5i+4Orkxe6oEcw/BOqx4R4rsPJNSTHmPyo0GqhugrWWepixrCRaD/Xl70s
bwLnpruvofFkhVcaNQMVzWptOJJimOi8sbWUgPD/3fs8ZuPFYrvMQvD6/9+Z
rGlF/d/dVhdsSnF1bkBuHjuvF7ei/FKKBHpfOOV4t0CKE3I3HOSMA6dswSJb
c9PIpAR3bs75RCGh/IDe2WWQeNPtZ7r239EFSy+mzYpBgJ+YGDcfYLTE26bh
xgDzYQkD0KupbADILwAs7k+rj/OvSg1A+K0hSoROhp278S5Lhx4o24mDKrcP
AfNCzgkVdYVouopHq/83oOzriSEUfIC/Z9cP7weg41kYpsdo2T4iCdM4d1kT
7ClgKoVwLts6BCmSt3N2FtMB/icmsTk7fB56NL1HmwSQJFBQAY3hqbnb5slr
YUHozU8urxKSrSiIcPsVz9Gx8ZevHpKoW9N3lgLpHTEb5OXs7yaXg1sGtdZX
uLoEj3TYpPiFMIMPa8PXYtmhA0Gj0JBNdR49nXvaU8i9MYOcECpuYOIj3dgy
C73v/XXntHROqA3abWXpPCGQ/H/XZm7nChsTikDJIZzAn429p99jCz4KoU8W
zIfeaRrCv6AvjxTf5Im1ysMJ3HdSHDBw/2PX8nPgYxadeVBmnvhXvyy/KXm4
Bi1vWAzzbzdwX5Nok+xrcBmtSMvMG5IAN62f1t25665CcO3BruANv8ZlMYNk
TioiBWKgDzcjZEy1v5RmDgkDn3tVI61bkXTPNH6JvwNhp+mMAuDrzGIC4Ie5
GzZfdaZ8Dg5nxWvQRhUVVIJjTP9Bz9vNV8BfZZFvIyE33qF5q4jda5Cd6eH0
PXkwbYh7Er7wDj4gkPnomHDfg9MJI0UI0YUOwtmsfenDrLjdf/pkODLNnPFn
PAinrIFmpQhJ1sgG9ooep7tAPgd7M0IJ0B/cKtJajit3WjcC84JeINJBudq7
nw/F6CEdOLVW/oQaO4NbZZLvFXqAdUm5in9P2tsKgBVSX2tqh107QT9K0yeP
2ynBnmzbYnDeT7Ho2eYLO2tEPaloNKuzdhsRY0Yh8CBwn+pHfWwoTTzHcitq
jUYM2Hnm8BnNOpnfT/ahX6VOT4wGALY4mOJbNEZsQHGPpBx6AaaYHUngfNaH
aV9wrQeL065YS5eRoLfjsIiVvD4QS3XT4uKr8feu35ujNtoYEPvKKlv2zuU3
Lv3YCYS+EEK4R8h5Qj0diP8GfkDLuFQFVoIAOQo4/s1KVlLIjWSd/VU6s/Lf
yYQBoBtNF4MWd3ATYka8scbdPfC8ZQWRvlm/dMr42f0pIPp3cd8LWYg0rrr7
k8IS6X4NyQrqVTtDfisVzmFzrY/deGHI1aisexYAyQdAeciFckLbYmhNEhwd
KB/D6tItz8YofwrkF3sSAyLEgkcTOMKTcDaBiN+NoVchjBKnTQWdS/V3kApI
MzA1Kn+wc0JrMF3AKgeME2bP2qFETF6jBiCi5O0zdeOI2fackzsZjLZolnXM
0T/s+6puRZPqoET8p7ycRHvbsY+sPvs1nvmdfd0d73DKX45gRMkpmtk+euaW
s8oC8bIcqSwkj1i7wpsyICFKasF9hdA1A/+yVUsdtE4QrYZri5ogBzyZBQMS
kRekGPlVKsh4JaE5XTGPekFOc0ouBzXTeHI02ivBi6VrtoQssJLA2FLEOsFw
kWTsx5W8TTMHOC09HjtlBdysV1E+Ljx9rC9QdN6Quvk+Wl6Ld06ARY9NNMX/
N8YVUcJ4csmtAWiBSc1Ge9erwinYlGbvPu+SMVzMZF+pGBGEUVuBKsWywdlW
D6fpkwkNBaPOsvQ/WsK4I0F1uSqIc4A7anw8zlXi/iB1QYXot0QHEmf7wMn9
DgQUDavFl6afTuvLxQM75+4LKX7ILVeAhjK63tHfvaKzbgFwBBMTdPMIPDqT
t2QoPOP4c3JEB8XOKBc3+aT9tz9hNTnMqbF1PpgAFafjbvqrueE1ybQtL7wq
/9/oIwRnnVarbMAR7+hKm9AfV60aJ+T98eePHcvptyy8oBqCazqJ+Pz/touD
4reiIQZNe2dwWRUkdTLl6UBxfDYB3Ftkqs0I8JdZMDDioGygwM+40eTOBWk4
SyADq+ks4mO0n+CjjpLdpd3JtETP7mVr1xi3Bm3gQZgPBXu2Lkpw6nZRnGnh
FHrTNlOwnGXWHjPMkvS5VvuN4LqSRt/1epGQzCnvsBZ0xMXvd7fBjP0a2gs/
eF7zFwxE7ICXXu3/+nR4LItU6PUHfrAyYpu3ykm3dn2oqS76oTYqx9u4d9Th
l/UZSWYHGILAjIVXAREJQdaIncvpKcuM/+xAWrabccNYX+UorW26jr7aJOg2
DUuNFhFabpba9coUCJCEYRYUPviB0Etj+NoM9Q8oU2m4vTEsL1nsCtbpq8zq
Xbefm8PkVU84w6tqAENXZZ0HSMYfzYRYafquj4QfdiVAWXK444bxBipBu7rn
jS9Qlp5gGelglQBUcip4OUzh4HrunDQzl0mJ586wwgpiOK52/T1YuTa9PomD
ZpOUwaqDEpyNmpzbCG95W6fR9LNyT5JcNpaPS51fnKr0KVbL0RDjvwzcaCKy
gU54n/kRixsPYEfx/tk8p+nWY6/Ov2p8NX+EYZ2vlMPMYqviEtPI92z+LPbi
jwiCbwA6F/58r9Ra9A8Mu5dCB9hlDAFcEWZn62M9t0hldnxaXhfmL7cbgS2L
hURud10qSTLc41KZw03Hc2b0m6yurNOQNBFNAEoopkHQiOuGPWl0CSspmIoc
pigwmJ/hFF5y0hU8FXZ+dQAZV4uGEEjFSOvRSL5zsIMZSs4/dOEphX4k6/Pa
LCrO/k6G0oV1Q9Hcp+Zykgyz3u10bxZsAVfz0Q5LiJKXOYlXhpRD1bizgVe4
bHXDDB4lXojNXOuA5JWJ9dcFjb8XlLZrsx+rpRY7xdoFRLy9Si0T4PzJZOJa
Q9lvjoNXps5sqjqjOuPAF8oZQS2KXoYLJe99NXNkFYEu82Ydiihd9ApmX/TE
LuV5kyDLoHyUU81OR9jrlHeN3yaLFbvaZBdlY5ENu81pBY5NOarZbdMWpwOV
itNnl1wbf8LIqqwNtTaUMGvOiIEmdOlMtVEJXGDkTgCodS6eXPc5XsVpfGHK
PNpOOC1sqIf45t5G2ZydtIJcx4uvzqezaPs18gYoSsuUmTYwvbj2JDvzeaWm
8Z0tNTk+q4bOOefo/58K4TQnOsbRLy2y+6znBzo7G8UFhC+HbmpxA4Aqya3v
6RBPEEuuHPW709LSW66Sv+o5Z6A+E6EFML0+ndhL+KXlrNappKKN6sulXTCi
yHPyKR4b/MPNcWie+vTe0nHoYwA0eeeVDIlWh1HMeRBBrpUHxenXiiRwts/X
qsWRUO7+yQy5j9mVG+UBkyFOb5QkIikz+jvsPK7z1lDdcNAWpgG37rP76oFt
D9wnPkuVFwKsGaswGRx/Yd04pxFmwnQcSSaFHU0y2ztkhfTASVWMirJJNj7m
LanKO5n6rE1R4Qa1JZ4+FOiEeG1NTdlWiXXmw557xZBHD1T+P0kcvJ7+8sYn
2p9cMAIDeZTWp+HJaSf4I/NSrWbJ6Cp3DRaIqaIylT/bs0+t+Lzp2m6w5dwB
2VSN/aia+s55NWJdoxnSWmPB4C0NVIJXuaXbogIxsyK88QX0Ym8w+cpiGJ1K
PGVOS57EwMyjvsBBwQczcp7CGmxflW8FDfZr2u3fbaZVBVUhsWKrMnGXCIJh
KSsmF1xTzBjsbfCDTC6PtOAiv4RIVdiBUtLJ4tkyZBs5Q1RBVsVjtoeAUtyZ
TPyxid5VimDx6AKkBT7Jx0e5LIsldlFAmbb8QDlQ/iydMUA3SVHpyyG07iLN
PYWItZD56X/Qbe5JWWBAxrAd6Bjj3y8QechxKaYi3ugsHO+liSmjW7E8558x
WuwovSS0YkzdTLSZqQQMIcBk4QCEvDpCrLS2WesGzRE22k/hrWKkA1OGWQw1
sqMtt4UKnSjVSTdQ+OxPRp0UuspmsW1ftRhfJGqJqNDdsJ6Jk+fsOQ1sGTAu
tKoHPGQ6yrbN2uoiN2WqRLkjES4fmlnpaSCi44axsI1/fDh5uqSVg0RRic/p
NUF2w5qBpTyBiGgb31zX5QzUj0Jpz7kY++DNVU4pPr1BiNPZ5ZzwD+EDzkLw
qo3ELn0VDr/asnXpSZmzKpumfnj26h7iGDBmDwbDc8ZjdBbY+91PbMGf4iib
KQpszr9E1DhJLc3Wnwk9KcUOk/7X4KdTi7w6hHU7wgIwXts1OFgbyEbtvVwn
2JE3N45R6nO7dtkVjElaI1iy2ZX8txCfRmsssEhn40IFUAVQ6QxBi0wviFh+
lJPo0ri1l9zbE1Ax/LgCfxPMArT5CT3UiCQeWSmllwSU2YqVa1iv3c2PjW8n
ElOJbh6KlQlfbKmZzKKdQ3yG7Z8Bz3JtcXFOYKiedYmNpGjdlskZZ5yqBAJV
apND3T47h1Hvy3eAMUJvY7IHlUtQkm1Y33e14QHhZMO6gRNUwT2l+m8tUU8J
RZwpmF8ESJMVVvoWVcpXd28agPKueEOptGrYdmLILBFDJVQNIb63eh6F4sQp
0MXXCYin/F1yXO3PQ28J70uXpFNYbgspwEwxECZu4RdnLTJnEyuqUqIbMVJ/
fdx045A0GeiwJK+TnlXbsKO71BNTgOgzu0k88knpyGe3ets0g0Cn1aVufebP
RwHXcdiitGyi+9pPgin2bGhyhlQdCDBH/RkKZU2A0eJVfmb6Sb3cUD4ITxM3
ICwCvjUM8Du1k97fMlL7ALlDM7b6LmTLCEjBdM1DzbqcvHFUdC4j5ma8TnwI
ojLpgyJcK8mJ4C4410TIFQApQZYp0aY24tkkYnH7hWw0leQvmC0OW0LMP5tc
h9ZsnoNmAs+LgfaHIbi+mvvS03nOrKnf9bw5hcDV1UInJzXCWbql0v5p8huS
vmoKZ0+AkrCgWGywlR3wZBPIZJ1GQXjN1IFVDsXtLnNwZAKeoAssp4OB7kr2
D79jJ614EfMF3ncaimFFxijPuZOWzpAGNG/7tucpDaBicERsdSXOdjsPLnIb
u6qayRhSo7D20mFzJZBBc8kKXGDvi8UtdE51UgTPLb3MLlHaAjZW4ZAWQRrM
p39PhimsVFI6SJZtwAxiKsXYgQ9ChPx66pAuDoc8yDEKlE6QPAdagZ5s1RnW
PPmysT0HvJ2rwt5GfNdLJc4EtTvxE/v8KZ0hbd6W7uWqQjSAH/CQ0+pB2d7C
Rq7CkbvcdZb7tHnajafqh4XQ84CXtvrth86CtmEl4LNFe5JbOiV4s4Mu1nan
jVwflbxMsvP1CPusosXMwrocqOKc0BnGnTlijYkOgEemWERHRbSfbhHLZaNQ
spv7zqPop1FCSYDryZGtjtzXCyqExvG8KMYurK0WVILLpIfu+6+T8ACUVVzd
Xfo5ICPTlgNELgVGE1vLu7tzQIVmINLcSsBao5kvysmT853sFyoYamw2pJ7g
fyMDAIh5Ns7gsHaWhrvajS+CdlZR2qw/0mTPmIrGa/bKjPichmHnoST1WnZp
jnkdFISB3MyG4HQGJ0P8tVX+o+uLS3fDjkKUhfzn+NTPYq4q+D67vdF9jD3I
aKAMrYT+Nh8EhOUnTFHN4aLpP6HOh5XNYLAF39mQzWhC6gS6YS6p/Od7FRXy
dUHJSzqwDJSLVWTJ0tuh81NCPG0bVXk9z7uTDmm1PBPrzbQmzO/Zk/nKlirY
cblyMMi40WxnIo0KehUm7cpuhWJZAFXTI/dGSwkfFmp2jmZVBCYuBWOBiX4h
eWbEcmpO1DJ+xnEtbeHKjwFVbbJL40Paf7f+PC5S5e9XYi4ya5BG8lqUarwi
frjKHM/oLU8nqdGa1mh2GIH9gInA4E6iZsF7Zmz+ZqbWKIm6LhA9ZPuWDQg9
jha5UgYTPugK5+9ZPaYhRZVLwpIK4iFEAiByAIFQcI4iYSOxpHA5YZC549lQ
lCH3jTHbRY5yhsR3sPrAXzMX0TW8uIeWb2xqWo99CRMdjmNs3ZH89QQ9z1G7
RioulnkoY1qo307dtkNVP5Wfy28xM7KpBBs0fF9OssYl10P8JYvNZZKyyHS0
+4JdNxNpp3MZTdYA+FW3epxurq46GQagYVTaAE+/3GTpsjOjs0m7AdWvIsXz
sXVOa7FbbXSE6RvWIiVqgfNgbyUKQN2T7DsdUnQWgMgfMl64S1drO99O3xbS
+A/PxpQyc2OahlUj4SszmBabo53xgtaJnh73aCO/OK5TeoGD4lNMKFpB9LKz
mxU78KQ22UAqIQ0QYE3tiz/MGNZdkDZ63GBVcEAstcg9rLTcDNUkU6HyXybb
cHzrV6a2OVkKUWBHGved4MiX2H3AqtCuSLxtciaHhtfxwJysJ8GkOt/0NM91
DBVgDMXPjGza4WBC6xgob4S0CNhiur+gRvS/r5gNVgQx+4y9jlyzo/cPZBMb
ZvFXQ1pcm4x3F+eVUHCuV5YW3drLY2UTumDSKtASh2/SLAril3UG9QBJBxts
wty/P6i6TpKdh2iG4iIBzUHyRXyWgAbY7Do5Cqp4a0jo1HJdErsDyjjfNcrL
wjS283LdT6R7LzJepTeylu1vs1iR0xybQecJoCH38xlXkYhjiK7rxJ4mKR0j
zaKtJiQuKQvNJnL+w/RFx6gqGRMoB+zQpMGQa4gF3TFccWs2XafRxz9UZPxX
E1xoiaV9scQSx8bba7YkEv5F8/gl1KgAGXc6h3uRfeMuPq5rFLmvPvzmHCPr
qPHEfd8MIeVYF6BmUy67StldPe4o25p9Bk69jzJxxjaD7RV4/osz0Pze3b9J
KBXvRuAvEiE2eeJMVRzhOl27fkRbHnBl6DSUJIJOx69tKsWUnm/uysrwez0M
bCzv4ovcu9ijNIN73giSYsrzhOGk+Shh+GmKCpf/XkgX0G5wcxeZ5bJhtnrH
sClkjHcXo+PS/+R1oS2wwEYsVRyDJfspytaoIT55WPlhFBbX99FbIEQ3FxSi
F7yKA4RJKzw8x45tsSqWcRWP5v7Nl55BNv3Qfonvl2UbjfZ4FKOH+MA/Nkgb
G5il85o3K2M1t3bPyH+GFj67e1bM5ZZEqXPo728J57J1R8yEBjWGUPqAAxVo
5czYtB4BJemGvCFej5fRljRhLuqQbNrMaJRuj5EblyLnKdu3d6u0MUjIr626
Lf71dx57VsFEBRSdl1vqMxwkmgwp2ErX5/RhzL6vLoVgiu8IT4NidSTfjh4W
wQZcSJWOXNgtj6rdm7lR9Qwx+Sm4fotca7rvXtAbjiRTOVDOc0x6gGj82tnJ
RhmBvcYkxmo3o+6CnQx7/zmlroJwqml/7vDeVQut8DaYq1ijU7X9/+5Cqz0C
T9/FK3VfwySZvW/svU+ynTM/MxPhYJxSe+lO7VqwGfafO/DmvyjubmgoAm35
vI+6XVkwXfOE03jG/4BHQdpe1wW+j7WaogqK8IaxD0tGyP7vQZ8hhWDdn5MI
wjA3CpvbzpHZQQ6gZjG77FbWONkzJVr102euP1Oy6VrnI7RSpCyJ6E13xJGf
l7Aan0lF0W4VMUxHrvneVUyEJ/6++ueXKXrqvEBTgjpEG8nVI+AgdKBiIGJw
0I3fjJi+7LdiLzEBJ/o+P789DjrhOWSK6qpI/tPq3qWoaEO22oGxpPIULueM
PLIWnnJwgsV/2Y3WaMqK5Ovwd3T++NPNQWeUbcuKB9+aUf8ezLoJ7vS7nERK
d8pbn1Xnw6yQIWHQbNAXtIlgQs6Nh258+YQQbVNyboqRCdCMMbDDvKyo4rze
nE2M33HtfWoCLUZ08KPP1ek8j0ynvMuzldpfX5F+46u36tO6TqBPYwMlNnXw
FF+IOe5MEJwJ7R+EwkFt05NNgPNTt/Py/dEBpvM8HY9p8tYff0DNHjuSx38w
Xs6b9Up3OnCReRDtaiZZzAxvsYFYrb/nZT9g7SsG8jY7fAmCyhfuW46nkHEo
XZ8Xfl11PanB8+eCwFYb8XOsltCppEfbFNMBJhPILbL9Yvi8dwVWDUQ+Gzf8
jTeDCkT9lxnTUks9iMHzLsbVIAumZLoAmY2bB4dB9LvyKrrKsay7yPHW1MUL
giEfHMKe17JsLMlBveJzMjcJi+kZDYaauKHdSYbVeopGWUmhGAt8Fyvfq6nm
5+F159JTZPITK00hAZ9GIzdEHLQnuxwNrsUi3I9shJV7xUbzpeA0E0dUUZL9
dRy8KHy+ILjOxegX/Nn3D3C2TBCvrLerkmnR8m8fV3sYAwO7TCqAgWUsJi7T
21qtqLPxoN2EB8QZySlGtFNTWCLHttRIqmxk2LJCALWZuRQVa9msFAbUgaOe
Gp9cO4ZOJL9AMeKKVGzIAcgivGoTMum4adUg/W3+y1I1CTMKlVDMIF0SnR7V
eQtHgKFyGScmwOz82J7vHKz2RG8kF2jk2la3apTrqKdCb+okQZuYKMbJSTcn
AcBT6gQZ4jV26nEE8CJS0TV76m6dWst0pKtpMS0u5uWKACXCR8qIou0PC1Ir
6VmfLS0xHAvq958Tr6pmWlkO9JJT9Q6SOwYpOHBHzEG77bUIlQOszFMlgT7t
dyRerYQ5Wj9iWscRkPcDoV5i/4HZKgySZriMnZehMqxynEJWDUL7tTVJgiPX
njnNvtiXF62eT57bHKhDHXMmBcxkphyj59h35Eujw8j8CLkdH7zGs29Dm91n
0WE8j4ha9mojVU7FPY1ELIaUw3mZj3xLQweYqrznUUBCmQciPJrbwTl9Sowr
VvtD1yQIouWks3Ax4PuEabuy9GmGthrBfuzq/dxkO9DPCADRRpCnhznp28Mk
OR6LmLSKJQO9QYDQWWK/qCa7y78YC2Ozsl/3FhFraBhYD+fQsRam41VmOlcJ
T7EZP16co0cJdH98ADkRttL3aUG+2i02IDWjcpIkr92VGrZhS+uhhpABjfif
vS/pM0gUrCi0/K0pAr6q4ZI1muKXvXAqxFlqdAvR9AwwGXBee+KLvsPNFTtA
Y/1lpEYYFgCamVnCFYd4CtvL6WcQVxPBrSJkGTlbo20hZ9NY5YNMAnPddK3Y
BSD124RJSa/wjukdsHuj/s+ZR55/PsKSPDu7BQMhXqzSC5VKdL5u6qTsGJSN
E8VnQA6bUrBoCWrx078RHCgh8s3TVhhd2qat1q9h7REwGw0Xmimf8Qx63sQO
f5QiAYD2X8k2YBC1BgRYcA1yVlK/oEfHicViiYLkxrTRi2gceZgQWn92zIJY
OjMP4XSCVyIImktboNBykBDKKYevyCkqjik3XoTC4jHWcZL4yyM0gqFWrGKN
wbuN0k3bqo3E7n9hKEAk5cyB8nx1igKQsp8zSmRq/dEHkOd8kMp+JKS0J3ga
8UnU6DXUxj6MODdk8mNg3/bDSkS+m4UHxWbDmGE4MTAk6yPTJ8Rg1h4lhGXP
9XiIC8MAjYubHPbHamLroL5pf7tv19jDIftwGIUfSaSuVhMplEAYxODa39j3
25ujt7IpfrDbn1Q3HmEj8g5Q7dthtr3Zx1RTQcnTOQ4zg/usn2Ikqq/XPvcV
qxwk+ogrXlH4mJAAZDp7T/r4k8StLPrbYO2VKKSi6Uhtt8AtH7/U0n1Y2m8u
CLSqplDdNFp+ifXZyGmtQ7lrqtwZT3SjfQIkKWP6eu7nb7CsSB0HvnlfDXT/
E4ZAjmyZRvTohwu4uG/Hup+uAdkUVitod5v1+vTOu2tYcfDfgNcteroJMeth
Ev3gbu/RIaLHFYAN/uVRASE1kK3q/GkhuyHA7DJXcpn/ECKWRexb06x+Xn8z
8OGhGmmRg+6xYVcKmBDuB6Q8DhbVrvbzSmGDb6o86rNPtvf+9yzfy5NkEt4c
rIibbkBIyfR1WWu0PUOnYm+eLTJvB9dHydBWTj/GUDXbRZY2Co5jzLAT/Fl1
f73OHghOwA6PfZ9m0pc+vobBSxi6ogMsJhaiYMdrPUfBAnguMPk+qSkdR5ig
O7H6cpdOorS9DW3DxYEbXfFt82iKPldE3Qd4e3iTMYfb9SWa9wQcR1pGzyTA
dO1T13yIwM5N7yv3RSoypu8edXQO5uS2Ypele5OFArp/owNL1ySJVZXM7Sod
FcfJ6O6uiX2dRBCUbxdOe6koAsy5bSSZlfeOzVgXRoUsmggl8gNDCaeUZ13D
9x58tDVCacc7JmcnDRLIqY1C6MW7rZ6xEPo+uWIdKJKk7Za63Y/8hnDxaKe0
RbiV1kvzQbA3b4cmjwUtXm07PqkX0+pS+uTrRYlyFUDUmiTFHBQJ6ne6Vmtq
D311NE2NIsyhorxcGiKljBT60ixoKimdpnQm4Pc6qrIU5qrwOu94cZgGsE6i
tdaKUoFPhRGnxJZyopqEoBhrG8z/auPzN4FxOJ+ltCFyDvLECahfNxls/W2/
fdD9OOyNjfHSjUaIovqs5SJeWl2sh3/NQZvWqyKK9wZBQTwYYn7TWDES4lPw
ngLNNJhSq+zYXclDl1Zshh5s+AKulZNLSO82mOUtl2SqyKyNxapSRLoPo4u8
LswYTaxk8VmtE5+Q+DyNcwrQwkFsk1bMMhtZ8qhBPdcPM/elf2mFzl7dCI1Z
vIdaggpZ4I4Joy73VWaEQbDpsaLcFmnrr82Hai9UQEUUpPIZwi6teoVkoeLa
6GNQDSAi5y84uxj3dSXm/hNGNvB3Zti1fajiRCvOppMjcF0EoQCDGK8uZhQm
z6kmNqQva1atd/WMLOW/S4FFWd+prejFU1DkWe+K1n5kxviK+7YAsCPukWve
ILUW3vUPGkd2v4N73budnABCSdHaQruylpmkwFFf5ySJdtfEbUQcKB1l8leZ
a4UmqU0YA4VoWr5jdPQxzvjONtpZ9OdvLoQWEoVNj/gYyYeSOmvpDw3jKb3f
Kxcq/PlmWV1lJEW3kueIfYqKL2d88PczeVdNqW8PT15qE92oP6WDKoxytNdo
LdZf3DKoEk6dQYjcsbNlN2msIq4iyCQxBtQEeO697nkMf9i7ovTLVYvCXaI+
776JoFOk3J0PJq8qt3OSrUq2g+KyCJ0Je/4+vjSr2LBoYGkM9ZD/LsU+aIpS
cT43smR5Mw6RbqeywK0222s3dB0ymer78j0xse5rtb4jm76xWJRyXMMDtPlH
J0SuZmSqXPIgkBhAVDOIGJZjRZmPK6SGpJucdcHS7C3gt3Y+McdimpJ1M+ao
9uc+JfZa8WP8j9+uQUkaSz16DmHX1i1X4mfoKOPTjPKxQPlH2MKKqzcgv4SQ
XfxTe6i+3OhujGNZ6bc1mmhWyrlirDxMyJul4OHWzBsiJq4R6dYSOq/FNWr4
kSpUg/KRiISXgmu1V8FjGR8/eTqcsqVk4NQi1LaueUpJb+k4XoPlCOPxVmyD
Ue2y540xV+dM84aTjqGaPtTzbdYusAcelIbIN8ShpU0nsSlbffHg35fvzBpn
Hr52rllcYB14qd8UMifHZfVCE3zQvI74amcJjaZeFGCNcXI8sxpJPTwTkpiR
7ttVmiNtz28tehe0gneZn7wiG+KLqMpIFVhqtY1wn4c1hvsMcVm9qeher+yO
bDR1GvNLUJyl18kqko3vERug3hvTnYcSblWzezTxxWy8SnpR5336hIjhGLpc
cqYfDCWnxUCYA4i2u+u8emQb2ikd/CrzEsxoIa0Iaw+jueCbcas00EBEymDS
hMJCoXPF92XTW3exRzjkxwBLEJwxsbSQLg1tK5PqLOZwimFy4AAqhMBTto5Y
8j0z5uZ1or60cqoZZdDOetgmBA7+zMbT0abwpO6et6twZhqF2jgVsGv+zQg+
Rp9n+Gt6bt7RcgsrHNheCfs+5Da8hSjSPkte4+fwGTq3S3FpcKX7xOipKP2t
MaPIqoqSbIZ3p0RaeuXIsp18HSjRqjq5rm/R5luFkMnx+1F8VvkY5LHUoQPs
IKWT8w3zDYa2rZxO07MavyipPyxEIAUnS9DZAew2LGA7HIhX8P5KJcYfUjoe
SAx77pBG95jk7gwQgGgYhhS8l1Y/QTBM6BUUWYnusyYYHJZiT0rJyLRr9BRs
UFUbBMUAXtZbwWWPWVhXty4CJfa2lsZXSHduPaIHjJif28nzfOgRrMS2YB/K
8sHwdfueNCt55g1TG88DNv7ZYDZm0E5S9/sKG5QSmoBQJFn8HBoWrWKNuoga
EKCjMm42fK7HvCnP8qttTbG+a1Zmoy0CVgHpmDkk2SseUiILaQWER+Q9WwCm
Yw5wH6Um5UJ4SJT2vi08RKaMjMy3twIfRlhMeEdIbBNQuhpJ6NzZWvbQz/bN
Py6Fgcs/NEtfUhrORVgEDmx477AoQ5DQ9Lnp746sbRuHautUTDyisjI6/dBZ
bytFhV20L0m2iTJB/x4/oZyHRmoA/OJc1RoxusQib5yBiER7tSHJ9ZC7cBSf
WO8ITsKeSeP0fLL9cI8bZAjYmYduMCCfeSSDpiHun/fV9XR64tG4TBephpNl
x4iPRBg8UJyoNquSJM6q2qbxES8My0nOFblPyrc2DHWtUyjofRJbOiQA0AnJ
FW11+Q05rhjrOEhz9FA0WywO5Y+37Hnv3z9CoiJhR9Utro+ln0undB4nA6wo
GtrUnRSfMYkAN6Qzqgs3BrrkccCT4Izvpcs2Jtj9bk6gLjdkSFwBOjly4+12
qxHPts5bxgROQom1bCRwUBDdWVPD3DUyM0dOIC3qWOPuMhCszkn9LyMFUBnU
0ke+9LHD8M6ExCX52e/V7Uo/CXL4NE0NOZ3hoHgUEq9l9mgjAcivADWMxumz
OR1a4MVifGaHjjs0Z1DVA+f9/2BU9vQNwTy3nvOf9KZwju2YmYVkTZmTo/EG
9dS0rVMpcaJ4RyMHNuC04n15iRCirn67kRUt03pIxQtUbyGjW6fDKqzKod42
U2MlBtTfjfXBqS60LbgL0t4tV3+FgvEfK4HI1ALOcmjVnJPIrjQiV+EDEYaX
gwwZpnmANXt45OYTQTkZ+Rm+9oCnbcQySd2mfEfvpvczhYTiAenE+B/zZP7V
Iwy2QknqjocVK5M7UIAoU94e5LOakXTPuTjuvA6/4a53wCKnt7baHeHVLsqA
x7YKoUkSe2sqWvnAP1HTk3gGxh5Xe8KrNovcLhMOZ9GPZTJcdUZnakIdLGtw
fXP74Sbvl+PHQ2E6YCPWWXRh8U3N+hlOD0cK5V/caoePppsJMUuhFblOX12T
E38uat2ec9foF2l3azRYmENcfQSawXCINuV2/Xx6PypEHAT5UQJ1jFaXAv0r
6K6d3UG9dq/n5opcLU3ZQ9nUiFcycc4qhMxkmPkkeYCJaC6S1c/c4unB8Sfz
fBkNwBS03NA3XLn3EAiBkxN3SETG7kp2hOvyitKKVy7JloKU4WQ0I0NeElkd
eYcKMXwhjEkz6o/efUJ8EePxPNJP9/YD0OtITU2sGq8S1+MAmtvUhhuC+Bpu
Le0cuRHbhqNPV6syEOVn8JR4XPdkuDEr3odGxkVV6Yw2ifZp1YSFyX67r0RA
r+AWAECyZ+xQSE6nXEaHXji1k6vrAgG2VO42L2kEPubgAMwySpPUnnZC8vy3
KBfGziKY7+vEQVci7dXpayYJ6R59eTCL2t7rKZaK3MHZXPCYRnGOTA3d0ztn
+ri6/IQJaH2klcWRiZo8/FzXJZ3pijhqlfCpVjbt5/5dj/oNzM26msYFXPhy
wU9jcArpUtjs1yBhIgtPRVnNoxWbv1R25idxvLiAskzj8FjwR3NQ5Mch2SDG
4qGM8MS9Kqi6GjRqUteY4sGxxNP20DAgD/42OraId6kBDeI2RNa+kAs9i7vW
+lKjouj/cHCorkQL4sTsweSxqI1UDGlSAejV3URCm3N2yXB0MYE6Nryf7Fvw
+9+/P9NRkdvsbr69zObMhtjoJQ9Cwb1xZCPa8tMLNDPOaOYZdTOa3ggPyRwN
Yf8T/5AmKKktrBl6skKtTGxA8R5n5U4YRreW62qLTCIwSv86QZK4TT8v0JUo
pQ4Iy/h/vDrBy44UG8GzJycRK5pObIxe7bn5+yZQhUcVlAsx4vxBrzZu20WA
JyF+BzkitV7KiKP8GKuqgdZLs8/lHum2YfMrpbcTP5MC4w+KPHdUxkcmJtLT
6aJBGyyxISWIlZ1bNWUd6CqwnHpXL/HaGWE3qTY+ZgpJaNW3W4EzsK0QEXjW
b7KMMxFpw23kQ/EiA8LQe0ZIgsMI7EDlU2C36K1oqD30GxkRcskrEhePgjk3
wx6w3faVp83U/xXePaeGe0JydopebI5Yp1+9h9Bjs7Zdst4aKIpLFoR6Fj2U
K10E8BpGldr3KlLXfannpXRl3/mG0PGb3kJpYOpcQUUdQOm6bw5O+FPeEiHA
aAuhJ9/64UVfRWlHoX1qLPaRN8dWj+XJrbALUreHlmsWExdvYknSST7ZVCyB
cFfXeqwW6ZUOtSYhVL9dmZlZTUiFCdFehdcvzW9U0iVhfjoAeblseDqKpc4G
OchGrS7rZJ+XFa74fxP691MFQR3NNIu58UY/oz+YIruON2rSTsELDZQSnPqg
QCATF2Q4UrKQix8+O0SP1vA0E6Zg9wJkZbKWjHoOsKz2HPRsunOG4GyFr7Bn
krwabgcmZb6NUFPbHaTn7gilnOx2rmK1SKe/if/wyMN9BUkhAEp7+o+CnIzP
9jSvfHzsyydDAEtzARhW9D8Wv7ELxOJWjVhvoImigGpjgQPKVNBlw8d7VpUF
u/TJQDf/8WJQj5I3Ct+CSVZgIfqMHYi+HFlqJkE9f5f9mfDkOj5c5xPB+6XV
VwI/4OhkDmcmjg7KjNYZ7y1BJjZO71zPrQTkCYBy+PIqsqkPR5VaJI2C3ijx
1jLpBMC12/TWcdwZ6NKkU2a9d+6mVgq/3EqkcWOccxo9d2ktPlSrpfzQFhPy
5UQcETX1CWmdYF1FKqJVp9XwVV95jl2kSeUMISc2gP5erNhm0221OKiVBkSH
YnhN3wpXQ8EYUiA4mn7ZZS2l77t4EoH2IiHSWVrg89jo6/WYvp7hB2jVeRU1
GvF6zNnDMZpm8yue4yw0+QAZ+qJZGpH7hLrSezhJzXmV4A4BMsGadjkDmois
2h47ptXltPOL+vLlR4G4zhhowfbSXALsIDgmH9D+kXz5Xoe4pOzgZjENjfwv
6P/6+AVJCNDNVtb8wmxOmdfstut2QYD+fh4ZdflKq0AFFcZGxa3JZKHTUZF2
Pc9rk82P88NbDAdERRdYWJNVmQ+N7EqPNvro1DbnV1wuklRo7f/SaO5j2pYt
vSyWs+BJeLztUzbrYEoMYiFqUuZhnSfMxVZOL8qWFsBC+xaDj8BbreLH8LTS
1mYXYNKfWdvBtJADJDidNHPg/djPYQikRLJ0bup2/Bg/LG36NKaPsqC0ZfI1
CM9dRz/hYqKCHa2ZDqueRmVSq+u0h0xi6AYVXnlM+jyXfdj/jozEXGfuXf2v
6xtqzzjf7hFYsZ1H9BhLZu5oduN5OVZYhjMdFf+3UaplvM1/U7AKv78EcL1r
AYPmxqTVdZuecKOr7h5GOsjW7Qk6tA45qFHxxzyYqPbEhpPyQ1fo5+i1xoLA
/W5jc+h6n0hbaIOpc22K6FkZXwvlN3NHHpc72JZnvX9fbwg+BPupFd6pGVdl
h++YBJ097++0jOA3pDy2v0CrnMNw6G9hTPFgibUbo/1t7/9ozGXGjuKM85Uj
+Fhzj1U0kRviU2LbG58aUQ94nebGxTrDUR16VfvI0sA4I7hrJqqDFa2EaeMt
+yeUeyiTB9jXycJLzb2dlc/mubzEBgbHVzlsPqN7RV9eKFPCj2zdIN6H6ciq
/+xQHateUaN65QsfIqjJUXMexhUCkQoFIkXIfKSW3Q920FkivUuh0oGwQuBb
JGhTIkYG+elrjDxGcljUgM75Cq3l4jTwJ1AeAEOeR1xkuVV4VHcJ2FT/6KGz
nRUB7ErmwQLEAxoFx6qVY83R2YnX/bzlBU9aY/4ppcoBYKiihwZi27bp4Xvf
xPYqQ3roXKg6VYt5uDSmu/FxYrOcMdUGAPBYGePGprm98SX0UEA/1A/2w3uJ
Uz5KLN1YhP/6XrOYgaS7Ae1Vb5YHuo4qvtNirZ45xpGxLH8Xfy0Qj90Ri1qr
0xKGR0flOgWAiOpd3ytFKflH4aBgkAdEIr7ajNbzoIGRHiwJPZChvKdQ0Q2M
Hnn0GKiFMV1udeufJDW4RKvxwJXHd087JLkTCEA81SkO9OQi1C337W8TvUi7
OMLSwo5FOwbPZocxdKsNNf5W2PRQvBbFvoZEVUi/3/2/SSWjIm0Pkytw1SmF
I8+G1gqJ7vL2jqn2FeZzWMdn/OMoyy2aGJcB+bG/D6A3VX0K10Kgg5ra7Rrp
blBY+qvjsVjPCFjYhXlUphnVQ7+IJi345JVqJuma4ENzBwfOAteop5mGiWCx
G/72qT5CPBwC7Zs4xfolgUR3+qJlCgYZZf1pr+9k8rO53WBeVs4lrRsMO1Ul
AojDHCBVKawi43deosqc0sPtgqkGg/GQT2F88vY5t2Qlj5XDndTn9kZ6B5D9
DFcJwP558T8Yxwizc7ZNrFMGmJs8cwWU1nYMCW8HwnqSmO1R3Q5v/dHga0IV
7QWpdreOQQQ/jjK1ba+VvkmFvzqqFHq4krbpGnv/ZMoaqNqWulL6UeXQ69Wr
rxUMG2PCQFH3UDGRcMjbnx+TJc758jG7Rrc4Qpz3qqtQKmwrVW8SEDoqROsj
MnlGrcMCIbc/1SmoEwvcwYOHUn6DlFS/XGJdSUyAlAxP8wVtA6ay80r1YNO/
POeGZeHH8+OSrx3HSST+E+GnE43YZ2urEAupqsgW4iXCIvAEsUgXopoBCE7X
orX3Ea3sq7GcdlowdVmMQBOXXaYANV26VfvzTaE3vjyHKnFiOgmiFqCwhxdR
bGHf9aDWkybT5fdG+LY2oEuuM3uOWW+sCD0QNzxB+pYGc4sBTyI9YBbVfj0f
Z99J2pxuY0seayG+mlXL5GXUvYgO/ThGE/7DvCEafvik1aI50FLeNz1KRe3R
oi9YKEtx+7pRrClgNmAAN7sCWLOaMMuZWux7Tm7Ee1o8aRd2woMiqlsxALfn
jDsvSRr74MCs8qMHFSJNZ2psYegTvBhmtbrjrhBQIj/Z/TbE4aUmZxVAqSAr
1SGpoj4f3XLGzVzbEzFGpJ3LNufFZC36bLL2H4ZKfbNW3zT4UW0R59egajXR
qW/Loldz/xf/SYd1cKCVjBeih5DcrbFSPPFGCPA6+1DeepsAYiN3Pj0pLOzo
0jhwNhH57nC0uaa2uu0i5PJPjdqpRZFHBa/BF0epmWPRrVLKvG1s9+wgYYnO
LjYCzuz4aUK9K+YM9VC6GZPfa6ItGqrK0HldmsCSl+O3nW5IPcDy8BDJW8ld
tnq5BM09BRSWIez2Xdv7zXV80fVip7lCkb4BtFwVSgEoom1CCqcy26BQu4c9
APBa4XH26yrJpTBQPtaIeXtdbxvRdLWs/USrgKsx+FIzFrN0bI0iVF+t1GbY
66jY0vCtmIyCXDQ/K1wX2euFC7h6lznG5oF0y5RAF+TbtV7vS+JhTpr3uRV9
PpOjFow59oU7jt2OYz3A+DBcRIN6RfcSB1G9VQ4XgTpZs9eqjM7m7HNp4WI5
OMRrhFtt+3MKWYCxIaR+ZHjb4fxaWxZnu4XLdZEZn2G9uDo/jnF8f8hJMWVl
fC0n13OJEr6gPxf22tNQ6bzsqWneaYCftBKJYLW6aSG7RAy60IAWgC53I9Ug
OSYBOAypEZs7gssPu4Mbytc970TqggnCmtYPzQ7fEOlpKrljHgrz2WiSD80v
5CsGQSmuqaUOxx9l98XyRrDqV1oGUkC7akxmwfj8WVn3ixTVnRMrKaj7gYbU
uzX0oKFocTDd6omCxlJMOKGWkLKFLF40oUxsV71Kj42zjErSbcVyz8j8HQWn
EKXZrrPpPG4twBSd4HBsB48JDxKCMF+9GzOoalAVrIpTUSsOg4XI2do6RBf7
8YGSbgPWzM4/LSkoSE75s49IU3RyU4BsCULsojQWjj8EqSnLzQmeOlPuC2Dl
VJq9B6r7WuGVlm/sB6rb2HsSMK1IHMpQ2n4rL4DKrbusXCIS7SnQMOIDK8QF
AhLCc/x9VGkZmPSEsrdxSwsXOaFjnmBtxPoT9mFDsJ2orfheVnkEZc3q645l
VbH3xLbKjX1A0eMG+zawft++lOosIo+4iNjoQK6BumW/JdCIdOErPlwtsRbo
Ne9uuklZRowPZv1JYS9wnAyuCl9JEog9s+SBUCyHbvTO/PFXxmwO4ctqTERZ
vBCkZa7Ig1Ikg0FdU2RsbCJYeIDvJt1UQ/vQGh8pbACjETvyvRuiokLG9ZB6
MrILfj7ubEiFRMPyWcMmAYR+ylMXQ0VU3Bnii6RN8/dhGJftb9rAqRRPpqsr
KXvmX9ntMMvbHcPFgzuy3Q+N9Kib9hwxKGqj+FRVib9k7lGbID0A94vpuE0e
Cfb0QqZ4NZBvvjx3p0hIKf9zZmaRDoCCTGHixFxpPI5GtkI1R2dRHysUUWbz
ZI/BAE9Ob+kthn7+i/0fmjhJ+f5t2UPsquYS3KhLAvTl0Tq6zFLj3oNO+dOb
G1NhTybTLCyIpDeFrPBjlA6wQcXl+pjgwDV0wWLcfBYUTsQhrPn9hi0ulm2h
CrzSx0OFfd80ums71XRD2catKugQ3ZUKoEM5rvBVmADbTBWkeZYzJrVbEosB
fJcJuTOFFfCVsYT6qrgkFL5t7hye5Jo9nMqdCRZMEfMkm9kGKThey+yiHjJM
3dN2We0bd2q14y6ditJVdnlgAKOv3T1f2CmehZuFf6gS5ZbdTaHlXJ561sdQ
AMibFG9G9ibXMvI02OtqQJNiXlMJzzozPmJev5bzBhTKiK7oPC9g2H6m6Ajt
EHv88CBfohzr2uPhEJH5MIv2um+r9B9JwtA5KaePZZNW5Jekfbd/CmkgXDm3
LVTRnzz5Xu9Jqj/rEE0qUGYyT1UsMFqAx6yAR4EtPkKudThXOK4L6XgqQcRl
2HTx3XKH5lDAeKChiH/sZbgmNkzL4eHf79f27T9FsY+uURi2OsaO1fsiOsMU
aKFAC+i6MYjCvUxPasy7pbEMiLkfwMKiGZFWFBtV7tHFwSFEz9mhTX5673AS
XV0BxTn7qOp3Yv+lk4ULyrKFQheX/Gyk6DX+0+ymghbeqmb5iL1sMmSZVHSS
7iQq7OZSsN8cz3u9iPHz6TnFQZT1PvrFt49I4hYfFCFRaWg97brSk03YGa+I
gZiPlLD9cb0+OU2eSToFPmtBeZymsn6Yk3whKjhi0qFPB8+bFRAwGIJ180e8
qL9pUMrA1of/2ToT30QotgTekFouQ2p9L248FWXLQrIJKYtM2jLup45AdAgQ
8qomAfbjHWYiujpZ79FNkto6xFZIgcFbKoR3OQHo8IiCsjsAE8i4YlwwJKsN
JswlNEXz83pGi6OX41FE+jfo08lVnCC6PkzxZ9enKmxhmQB5gJ/DGSI2oEbO
s2IUCm4zOGRu43iIfA53aT6Krc/TlNXpURr7eEl/phVLHf69er0tLXA8DiYY
rBlaPRMSzr7UbtG+NWcViV8TZXnnsBd5eV80rMkvhgzlzR6iCciJL3rm+ZI6
cU2yyK70fOC0gnvpMom+dpnErAfYK/37JZUnJtWBS1am0I2bgLpgRpkVAVLq
HSKGafs/rqrgBz+DL7EUPP9Tje3UeNYlP5HIsrz6T2JPQQTn/omWWqqejaYI
EZZ6CQY80JQbvYKsmMwnDsIllTwWI0pdcokyVYvYa3xEj0I60H6Rc1eaKSsQ
9NxwpZys0tqwQcO5MbUo7llCAVWfRc4uNOvGSkrIcs1eo7hrNPlApxZt5Hog
bY0y/doOsKZ/BpGlw0OTdOfeMHS+OcFhJRO2dfv+NSLDOq0LWyZHEdK+Lu2u
xyuoeeM2QjhyLlPuJRHK99TXD2i4ZiYG6h+951fJ3kASnYY6t78GG2sNyCAW
+6Rd6wQxOmfQ6UdLY9s9ltxmphEoRabzY5X2BXfy5QxpRvED7dRQD6IWfA+Z
ZLXXgWgkPFzrrZrdIlhp20wFZqvtAHN1JxFb//kQLm3xk+UVJnodHDUfd1Il
cPeeCSITq3YACruxhA83Ae8bT2gy/AembHq0PArA5jKe3NyP8flVjSBil0uo
pTClgDEGQ86WwKKvXNXcQmlfKD8kBz/5l6RUZgWmGzMYy7yhS+AG1ZZ4vdCm
GtlEZ7zKdCA2s2KhRrY0eUbDhRK6IchS0rSyP1+ehBq6XRgCWTsDgpxMhmo3
/YwHhSJdUJA8+fR40Jtb8tedcvyvMhERlvTsfjOSBVsuKJMY9GptGiMEOEb/
8pW/UQau5I/XLeWO4i5TEmNqBULMifnzsZHbwxWnW8P0Dkp/PHJAj/pwZKnF
7+TG9nnVdYKio4S8egN7KqgTshCnQF4wF74cCGOSi5pTo7YzetXJpZQqiAbt
gab/NriZ2tBI+0mawECuEMEINY/EHg+p6SZXY9o/MuJHtXOtR4wmGhopZ69/
ZriECCnL6mLNP3OUMXn8z+10esjlFdoZCdXuUf4QwpxvMJYhX18/Gab3Ijqg
8uId/4UGPtWMoHuxkjKvfNopy2tmm0pG1ACIIv7CBxy82P2hiNyWtXMmaGLx
2Z1D2Dy0QNIk4VGcgkX3/YHbqFOkbo2h7Bvo6tl1mXZ767LCsVJ3EKpQKz35
oxMc40H8ne/BSgfsMuR9zhOa4MHs6DSnXv9o7SZQ9jwt4W0Gw/ixhs6CrZoE
SR1dmWl2lfNtHLunK9TTDHLbMZmgzUCmJfyS9ryDih5zR4AUsEYzD9b3T/45
Gpr3+FSaOZl8Ne/YAuVCAlFGh7Nz1BHlgoHnS2WDHl1BiVuRg6jYZPIP8nqr
8avDeYVpNyYjqbORjOv/oJwNF+4lyMl5r46pAS6HfO/QHM2lOFnTGVySIsAl
6EwFCxRk7ldrb3meKk8AAYxS+WkPweVoMkVthe7s4CE5wSk752l/bJEc/s7U
JDEw6qzRV4hs03eTeS+7fAvgA2YY0i6BmEV+RyomDUnGziTdcibuZz3Oe4vR
XQhL53EbGeuUlLdWDdOVSxHJAVSu7zYTaPYiadRUTt18lBuT8XZLdzSzUbyY
gjw/dde9lHopmOEx1/xPtiL+6z2sEoYUXdnPUF9G4ip7wE1bqqBxysuPXSVd
NXFsQKQWJTu+l4wQ8k8DjsDr+MGj+n/RgW4mQMhdi7ltSg/EGWrq+M8YcA3w
eNitLHtg9VoANjyIOe9PvQrbA7FW9avEQpPqBuPlNU4kd+UiCw2V5om/UbbW
d0yjkdoVlCgbPloMEEGD9LBkVwY8M4goTYLctjDLk8ZpPGTA3CeUYP1yKe8y
FlQin2xteQJssGBgbxRemCY6lcKeCmBvRMZ6tipRE78LR7TA5FVWSbAySQ9L
HHKyryUO0AkDFRghj/u4NWd4iNURs8jsVM9+xLcd35ueGM/qeGv3lSfnbeXb
kg57UPHVBVramsFJ76tewJCMzbBSWGbxttJ7A62SnxgDrsrcmOoRQa1GjY9K
BHxbww+G9lS7DmfI+Q3f0mtcqYfEjlE5dHxhS4b9AYVNMX+NE6W+J+iBz5nN
wSZvd/jioJctHPbYMNuZMRXGfUrKFFCpog00wILewnnsKx/97D2MDgZ6sBHs
fM2KzZ8Rfb6rInT6NuJBUZUeZp/30qzBvccrg1L4T2n1iV0e3sFCAybkhn8l
5qtRO8T3DimBAdk0h1aZwQt1L/RSqXbwfSOv3LLI47mDX90Eps/s41vZR/8D
bY1SM2sDE3Eg3zHsVEZyFyhqLwQSpVdApm7PtXD/acqVOd4951PHuNjvn74p
DDEAGvMPjMmWlw0WaimUXBqGe31qAvZ+a62Y7tWS4uPUUf9a9BNMnn3VB6or
d+BV4x//srhpOz/7BOGn65MIxu/hsrlEEB0TdoP6DUZem3ZMxnUuew61xBJz
9A9w/WA84K2VuBUlpndfzvX4HdCg05zEQACcBaXHSpq7QgfJGo7pKUv8RbV0
Nd2oiMzE+G3WSeX/4LDWMkxSjiGhjMAZnwM/BGFMmXZMzZVOEcWcubcO6Mmr
B1sw14PmgtfkzlLKY7jaYM/KGrJYT4to63vhRgyrNOhyELUDbzGT4yVpjfth
DaojnFZFanlEuY6OjZcjcSDb71Re4yFbx9agV5+wYq3VUo07SKFWNmLlXXOL
2eiXXBPFPr7WUudoVK9ALgE3iaRBHLXpSODRPdwGC7aFIijr+nAPwpHSDKpo
EW8kfUVvnkbK+tOCA/blrZ8hSyIJoDMCtChVKEBcwHmAwRQjc/kLeo6af7sr
qzzqL7m+kGmqcbv+ebeEgJc2rEgmj/aElOAJA+2alDzjFda176auBmCIr8qO
Hfx3Yb8WEnHd2xppnztAYIbRJtrjnJqgLBIKeRx92py0RtBHTS1K6pNA5jSD
WTocg80smjV0n4FW3JPhiUBk3eiSe4hNMi3NRJwnsvqoCube0TIhHvpZhiYj
A7vH/WkHSuYSaF6Yn8l+IYaJv///Y0xqmx6YzUEnp5zM8GEiXIUBeaT8x3xw
sIy5/u/bVFn2X6zeFlnd2pI2xXUX0HD8ZW6F7kATE9Ya4aES1Wm7o2J66qZ+
GLUSDKdNqHkhCPCNzbGWeWtftUgNDLcCBiWQ0hRIKZbapP7UYveKTo9r0tiz
ijJN6tRQKMwLdfGhPZDsawI8taY+44+MN4TnHFb9zdaqUrfM+/J7Imvlh8dT
01ZR2eObJJQSR7onwZ27iG+Ut+z9qnH75n4zYvP2e6/du6yeZlGaQJMssd/w
dLm95KtV2izz+qJk+WYB0NAOrgPY4rGElCIUJ3poKVbRZDe+Xf8s1B/N1XZG
NCGrm/fnZh7SDtGswuDTuKZJVGYYbVnFavyPpG+E+UM5E2x78H/2PLm+DQX7
rxKoe9jzrg5ZA0eZL2BjVF3bPc6nBUUGVvHqjIdSmPKaxgihJVUP08rBbksW
fUTvfS9yHMgE73AKFibN+d6uYpG/9Yy/59GUWvSWZPkvoyn5DuPkED+6duOl
gTvCMIJyn+prH4VyiL3Vd/FhIYH8zUQF1uj+HpLMNF6YG1gqjF1oLthbself
K/bkK4bwGcw3vghUX+3aOV+cJ2cv/2MWde2uIBf9wOwqr6VPxOQwNL7AwE3b
+2OTpfSLP1DsryIbF7kQrXEuBAoBJE9//WvGQBth4S9yEf6zJ9V7E7h5ab3C
c+0osLUAin+2Ngh5lDB7JPKbbABHC+tLV7rZo4S3vqtWkBjVN5acbA+MlXcf
/xURrlM5REEdS/EM+N6NSlc2crUbxdUTFAFoirUDf6pT/XDihgrauOVs80S2
w2NiIRiV6eP32tUhfg6AFYZxjICeikmhzZf7jpyafCk4dQKtUo++mu8YSWOS
XoVMvzJ5jViMgAeuJ44U+qoF9j6YItOusfCHcL32X2cAo4MJ7R8ksBQlWZ2H
sOiRn05T1dXpTwicibMATRjgW/t5TH5byM/yKpjfFDPbKgo+S1+CFjUzXAgc
nXHdNoUZ7R2YXGEGGMYqB/WIJ2oKo2WCmmT/KmgI2ok9V9AlR7t0jCiktghD
yvTeqIagLen/hXuz+XFMyzcR8Cnv1Ulo6D8jPLy4wtHPJ5OU4UjxlfoRWSbm
8KBr/Mf6zy4iYMGnE5HWlL4M9IHqkCj9A0rm9WPtuRYY3bnm6n9Awl7pn7Te
A97blYo3RgKUDd1vsat9JUUDlzK4SkNZXDbCH7fQOWfToVdQNbu65Wts1hoF
SMIqd1Hsv2EzWNO5ay73b9DuCLrkzlBDKvtvQ5bnq69SbtLZnVQF9yBApB9K
TlaBX8ZTIwFsxhS7GPBvA9bn3g3fpauGwMn1tG8zeSPFZrQtHMGyGsODkAsj
CLuJNagXwLDbyt/jdGPSNk1wUGMKu0ELB9QDMtKRtnVz9rmwKnpAxseuNZQm
go+JBbAs1Jdr6rspOVZuoZOSdp8S29OchFnUwqT4GmuLpkFqZfjiNqI2orhD
QRDBi3KC3+WsFZ9qXAOFe0em37kIrYpLEbT0bTHDREyPcJ0h7HNVUimmC5cE
rGMn6i72o239tvPr6CsA9Y8hopMNOaR61m7t2Aweg+DMs3Ja/1xxEyHZUcNP
aGAknqXadSAucfOIeV+r6H8tiVAVr/0A6d5LWdwDktFXkPqPXiVl2FfRz6Qz
mtPY0aoOAOBLVJsq/A3WjwR+2ffMbegGOf3ua/XrPUfiihjrMm/a0cuM1gc0
KHj2Omg/U+vLvOVATY1tmQe+6yM0el5zgcgeyE2aSZR4nGNs+cXUMGzNmIkO
5Sr4qk9/webiOM9mIOljPI24l4zIgIZTbLhyetj3Qo9BYe+imLxVgFKI6uii
hKYdycXjpM3GHO5LSJWwsO5dAjzTjvr5zwY8+QHxwhw5qSuhNuAme2HQZEm9
E4IlUq8+R1YlbkfxXWAvwP5hFW4LhkJDutS1+Ufi0xDyXjBUJnJ7HLk+JcY0
NdQS463UDAM+IM08ZldNXeRUCatipXSPNlgxVpOW6h5tBjoCJVpdwo93rNNS
UJvYILTEA4P1oAHDSfGYoeMMN+q0KiHD4WqjQADxS/RsBg/r2tMNr3eH6RLh
iZaDL8X6xIJwpgaDzHrLtDLrEdQ2HETesL6N5h7deTJSSElsL7jwOQswU//6
lW8MwXycZSz66vh+CdKlRmTS5j1GKtxWcRWEFvIpPndwzQNgUEvrKc/Pdic3
dzYCzDPRANWjteIb0SM7TRapdmifrtimsWA4PnHOG1oPXXFN8uhx9A9H7mUA
daqgm/DllRCo3e9pcDLlNOH7REhZXSrMAD9aiccftWLyLztgm23nihHHsL8T
OkBvtSMRyi7l3v8sa6nQuR+xB1IvM+k/8rZKKLBSQxgCoAH5R3jT40JumwBH
dLU+/JfEyXMYR9kLz0WGCKYoInwK0vf4I+W8GZn904A250t9xTtjNH4pwalM
MFny67EXrVQulEwNONCsB/65YASCilbWPzRm9egJe291KT2LBC7f4tvjWUax
p9oUJ6Gu3io1PB5eML454pyZNq9fGmXAlOzWtthAWH2uAwpUiSqWiRWzGO6u
JTn+G58EJ9C+p+uI4hYCteXt0lxExCR67j2GJpV1s1zQTzy+JLt1b3y56dpn
gYYM5vfbEtC4T1cw4ipCLJPBVg5pruOGQ+RBwixQFxvldFRkZ4SZVn7TPaUI
Ayd9zR7QJiZjcWskCGOGwilTgPYMTZMaqx4HqWN7Z1WEK7X1SjIN/MxK+8tv
NRvpf2BMaIEKMDepiu0YuFsCWFJltWNtzQvyMNeTFevLzIkL7V9d0mmnoCIU
iPs9RE1NX7RgYILx38cQVz5aBu/TvDlCGJM6J6Li5PuYRAnkeGbxa6VLs+zf
uQrEkAI8jvGiA6gSaWzPtYmZwWtsigmfzjiMkekYdLrwzCioM50JszSeAEic
A29t6kS6/zp0pf9XkMBaj+IlfSfLWDFw0TjbfhimTGhs0Mp5CS23qO5xYN2L
FnjZtl6zXR4jqrO9nGQzME7uRQJq9n1uyJy9zOrmw8o+UcZQq3DIafyX7jNR
CPi3tJoU5CFlp//P5tSd895EzP9DG1KX7XR6/J//qDfVeRBi4IpUU8IaOdHe
fiz6FKK8+H1D/uC1Y9kkHdU0PcxKYS81BtI0MzAQJ0O8PuFCPVEla9Ecs6Mc
Cj77Or7efMCnSsLEB+aDSeW2roGDZpvQNwWWyFweP4H1P1saCkiKRqRjzPms
is+Gk8GdLuahUdlNiUaFXeazTloQiwS2B+qcFUu9gVYVfzkAbz/9Qbzw8m2m
osiEZAY/RlBFTXNBj/wpLBFdJ6nwIPyNHJd/Rbt1wSfi9G4FhR7aOf/nHRao
6D/GBAbFgznMD9UPLWkuNygmW8moJr7LljULOVioIzisJOH6Jjd0vc+6fcMg
Mz1qu6nKM6fi3Doyqi/yqyIaEXuTfvzyuZeme5bHsrFTlZZ/yDTfoo6Flo6S
enp9/GXP/UvZ/PI+S9N6MeYHuOcaqIZcxczdCTO6Da9OK4ljyT2CGCEWrqf6
prsOOa/OTbkk/fdrSI4+T7gHSdawuNg9AEA2OxmBmirYzyvuKTRFdy6hfd9x
XtMgjJGQX3xmbVTKUsxt+E3nh42Z9DyywDbjx22qMsBM4rW42lq9YqWeHmtu
5K9g2ggRKcvQs2mo1VP04LZlngSppbOkzh2hin0FCIvTHbXrGgYxCKW1ANPn
A6C84TbFSr83qVkmSA0ttUNs6jPCJkDnVP8L75dUQQeu6d750iT+TtNaCiRN
IQdhh4GDx9Evpnn725wgnl8mjEEfTWhCyTohdatnR97XAwAGYL48uNs3m12u
+1EjAKtwzy52wg+UlR+NNWYJy34pfY0a41yGMFuBOiZNoM6PflfNrzjv1Sj5
QdjD2zctb/onVMhVtgibtvhSnfkXjfiBQ63vV2D9EGXg3dTnJZLn9fBLQvVu
NxEnlepQzHbgFfNaTU4f+K+PH37S19zQSEx5jepjCY70O/SymCvsRFfmcEzW
hW4e6Jgshe2J3ZC4w63Jifry0tfMxsMc+EA9ZbyltMFloZJJkIdzpUMrQCuF
rWycc9nfUOBHFr/Nu+WJn4ec0akkXemrHrE1PS80rR85G6BvGwBtwRq3kmy3
X0K3gYcyyZSKAJdTGj7vufyUn7SIlRM2qsqElySY9kk3xfRnSHVWOq/BztTT
nWPWJQHExT7xhMB7t7zJVUphCmYvrKJk02djF+z0pnTr29rt6FpvP2fSzTJn
JleDBkfSZaCJp5UHPJGDK1R/1pdAiin+1UuLPYZfr1Djs0QmdUYbW67Klf6t
8TzvndsQfLOiiGJds4q9Zvp+A4YV8s8T+mGsENHnn5tVCLLqU1cScQJDhhn4
ExaBw+BXDM1/90xPTl/mhP/EfzV7NG2KVAQF9pIC4ke+2shdPXOisNoyaS3h
PTUkXSjspnCZ/ww/wZTV+0eqtCNn+Daent9y4WrFYW1+TnJN4wrJ5HWqnpS5
AfBPAl0maGqxR8X72CN6taKFek2jK03EcabtKysYn67uXUh76eY/5ynzEPpF
+2iFkdACqPR6YFL5Ie0YFmYJfuFCecKng+aEMkx0NJrY9W2K2dgDvsxsL3KV
v3ZxPkDciuW8n2RD+k6mVXKGY7sFD/wE3YvFQS5rI9xSGXzgxjpkARgdwWLX
rlw9Ky81i4CpoP/Flia6zUj+CxgSBTVBwtneuykRDKUXxfLiLoK+iYT4pkdU
Zpr9FQN26QFipGDcqe30NTyiIEkdw/8AFSejWxewJuh6fYgeFAA3o/HVZcBF
Vm4DFFit5r0NNO7QovQiX9G4VIQs9QecKDrEY5ehJn8CoxI80AxYQN3OVxRL
uK1j/5q0qZv1pIW0v+bOQ+snBp4sdVUqc6JKxck1mTcLygrNuysIZ9UTXvA5
gqNdz9f5KdyoWkcJ1r6n3tAQikjQoV1K/0xVUE8ggvnvDCqqpy8RWYGTSXVe
YHmU7A8uACpwKF6rKQzV3KWaWSQoHn8VVby6T0/tFyr2BooeqYtLrBjfxDKn
HAWG6rkySEf0eQ5XM6tDoR7uEq87ocNpeDP3YYMgWW2xPS+Sn1RSfifE50xO
bitfgVeaZlLvDmpt9EWrSB2APLbv6HQPvJSdyflMjtAM9bSeLO0v1+ERGtNZ
keObTz1CODe027dDaJF9fUdPeK3KhSaN4gFpkUVjsoLE4XK9dHNlq61CksFn
sdELCVBuDZuvPW4IxigYU5/I+ylPw9Hlblx2n1gdB/9hK5iG/BQWLzoCVGHQ
4t5USo7FpGYwdgR1jye4jT11E6RJ2al9/k+d0P2U9IRih/2ZstMr0sHfKxY1
0gasixehBFjyYjGd3lW7xBfyVJHCxqes0tCk4wpVKDeFbpWVcGVDMbUA4jjf
RCiXTjn0zyMhAxijJgV9P8U2Gcv1ccs1C1ZXk83H9A7qfDFEjJCrLokyN37r
hff80lmJa2fkzTh4pFgPyD4fkgZB+jHmUvico5mO/Dy05cZhFoqStjLAD+1g
UODlgyXjQBxOazA0I9QZ8VWh7r2WT1+3g7j/dxDbSCrkgPnpXqfux/aDNPkb
/LI30bx7lOkq24zslsi7CMInQ2WR/PWvrkbknOpJacQr2ziVMN36ygsMfKMA
suZMkzcLYTvHMm8FHaG2rXSPdw3hfe2c9Mvxiz9C2N64GG6w3cAEBa3JclCz
Jy7u3InCUtzXEMskmUbY8RRFVt4N4WO/vaNvXPnT5SFuzedIT/pH7tob5No5
2RLyQOB+g4kJNGRnmlFgmCDlG+CfaCRjK6Iie/rlQPFO0M1OcFHiYJ7MgjGf
oQP46JWvJSEMoNEyYmloUs3N+Z6eEOutv460fHfQh7hVebnYAdWWnRwp67AJ
tWA3/dxdzuJ1cuv1rev4NpbGyzc216atnvplj0EfseWijhJ40Xp0VY9KHH6M
Ot/xzeJqXhRnCjPXSVL2gdJZuqz3eVu/Fx9lJ26dvqYNdIFO8Xi5ZrHsR0zT
+MGCgtT8UPav4NUyb/jQbnhkNbXUvpjaUZYO5oQ1Lmtrx93n006pcuHNFRQm
kcNRTSVkTWdaqSLTf0Qc5LaQcV9MxuJwBlo6Cs20NGbn2MQWeY2KsSwZ3Qeu
FGbVlu4jhHELKaAQ05YngoRVrBXxJ10tcUZmp4p7DOBOf2c04zbtY1evu+r/
PKuq5/pnHaRdS6aaYPqayTV7yHpxjnahYnKVs6MAxUhy5PgJggwcawD/6uWm
qkA7PBTPBl4fpQV4FRvA1vBk3o4M4B77RkWMwAcVrPn7ys5EoC+3oPGawsl3
CAMWWm8qShDEVgjRexqgwpbUzvbhSkQgke40W/eL7ki1ir3s//qa51uoVZNO
PeCPL1ljxEFDY3VYcPN4om1BdFDhmr4tDk/uOfX1YcntAkBEIPidLaiUfVi4
qzj6D0hgaRx5SeZ39VTw7DdSMHQwJwJku7CAEUq4/c4/fDSRj+5yjaSLMUMi
K2yiQ2ajjwtwkYy/ZbsnXQ0LJjuze0zV70xmWOFdwKZTCikX7z3AllEM96ry
6GPqRV7FLaDxaI/v21QKdxxs93AFeXrA80aoMa8HhqMHD9mvuz1ZY30MUJOk
OJ+oJkVbnD+p+s1SFyTGh32c2EghkhkzGKF5Z7HYWjNPsHxQAWWgIKxmivHd
ONIeBVvVfLpo+etj9HbJdA76G2Y6AbF4NHQ2gFbQu4kbk3BobFx5hPvFddFp
sRe54fOcAcv2yDQ1tZn4tEP6G01Xt4eAmr99v6M6dOAfq2rxba1V6Cb6xgZZ
7gPuPAT9wE9blGCbhIIiXhANHEm39a2Rfp8Ui6TlfL/TcCRIeT6jv6gdVWRn
bPMS/5WSjlSm+b8TWDXDg3xW6TA1Mu1eEjqvCygv4CzSyjK8M0UYk2flCBOG
0SWPDQ1P+m50i22RkVVd2yeiraOFf/N+NWT4H5amy/TU4PZlMH0rE5Fz8G+M
K+iwNdYa4l7GsuLxg6ND01/HbmH1WyBSy0XcBpzxt9XXNCxtCFeSsEO8LLLd
7s+Nu+eLmgAd1DR9UHgKcfHcqUACSGXA1d2rxvIc/eEvhjFkCE6+e7EJm+uU
gexriQE6I2/AbiA3ZbSTY3+Zi46XDlnNXkWDcGcY8AX6LMvek7Jd0AKWZD6X
O/zwKUozja1UW9o2EMvMnJYmv7uiAc5jMWwDMDemON+TXocyofg+TBKe7lMc
c5+V3p2zmAfaKmbrUI5fzvslqiKCfgM6GWOJrBI1E+wYcsjk6LxL7mxuxPHZ
EgTMqoGR/F++nPeKdy4fIXq1EfXkO6RpGjBQn9zKSepUc16iIrnwAywm6TlU
JZ9n0w0yl+pPLE9WPSQPmCu8uABIFsKOGGjKmQKgF+txRuqRtajDcdlZXkWR
IaWXKSWZHdfmxroBA5SAHMaBmVE3qZdAQL0zvfSmUxlbr3J9ob2BRqLRRKEo
bVPnDHyxVy/UKr0nlL1YHSLXHKw2feR3RMNCOPsFwQyc5wh7SHqg1auE00T2
7R/D30kQHeYYNrYoG3rI6GD2Xql/HysUwy59v+WlR7XucmMI6mYj+IdPfaG+
KUBv8dGpgMLX1ScRrTC6rpj059s50FY16sBmNflhCVAOQfkMm+Xr3sHXOpXy
O5Xcz91+UXiRhi4IMD7/cLKbiwLYqJ1I7c35rMPw0m/RBNTLRrMaDXfFbGXT
JU+SpDTFYUpGWgYDChSPJvvqWDHamktAeA3CA7szwEYs7mPnr6g6hAdCY/gh
yVFH4asKVjM6FcNJyUCnA0OBqM3bnX2qr2Ylw9aUpRhVPsdUPSpAfDBcPhKp
mRJsEU5CYJlVb9pDemiEQwV/uIsZjH7MduO/aB0FELpmQ1os2Ws5tcafrvZv
Y7+T1sWmfeDx7fUHSb4aIRK3FACdu91erz7OJ6fT4Mz7K3j3smaY9K609wQ+
2ACzZjMgskCqVSHo6byZw4+dfu5w0NeUaAzv1a2rdkiLNtWEO/88S0bq7W2J
Vi58Bxv9fbeonLNM2WjH8cOp5dGsu9WyDABmP29upRGWqrEBiBovgfnnqwNk
aVomrMNgUSMRE1lL8C1Gz4Quir33+UjZF2wJqcWHkOmH1CG4Kp/zvHTv2qDA
AYiPzWH5gFgEtm9Qq7jaXeT4JuHmDEQYB0+4zH93pkGrkIt/4PrSffz/6t8z
65hz4QKVFISxSN2EJScj7TJlb6AxVBBGMMiSslW2rcy8vG6S4UQCETucj7BW
+vLDalLp0n3OsjQAffW/JFdkkbz2fjoTKqm+5BkTu2KqVsskU4PuDDYJSaUf
9/lg58z+aHsGTYDqSyuJGk0/lakSJcfMgmegqXIOwtXUSIVjPZku8p5xHlmu
hgj2P31cHcTL8h+2wOueRLYeAvDiTp97EXkGzQbbfJLt5MZszLHIxWOC5cf7
WAOowXXsbD7By1j5JWf5sJf/Jbz672IAdciiuAhL13kr3tO4jESSeqS6uPgT
zaKwustlBTfJ5o6/IeR99/JmfxEF2trV7X2qFShr768I4Sws0pZv/nIPigxa
VN3P0QM6ys3vWPvRHLDkUTbkkks6aSnSUgpTQQdLjtIDmO3fXIWgyvFqs53h
1TA3f5590pCJ3YyjIcKNJzITvA84pdAKuQNuuLdtiYG7Qv5sX+sYbVGx74LI
hJ750NuLyir5kXz9vuJnKVB7qXpMF9DwRCssfiaK+hna3PSAUYe8+M0FSZRo
OeHJCAK7PRfdoXGOPcQb51IHzoHOjZkMxviWlBcWdnBJ0/SsCKxxoKCnRcWj
Mj8J3mcgUt1VMwH+RbGUgBBB3vdVDxKIooG//ST61FT78f1SHDrozI+0ZYrE
PklYo8EUQBrXkhwu5Y8wztyyiqqMyuCD4SLnH1LlTKYmx2t7UhvhH8azkeLp
xFWvyPy8dQtyg75fYBG/GsxtgW44/N/Ke+mI4YHCtFUXh7sU1fVNlXbhUnXb
HC8Ydi4pIqj0k13068TCsr3tuR+q47z/bPRYpcKgs0sFZ81zSO6G6T56JuYY
FOX4SSBzxh6ngeBgi4Xy8FgXKlttk6dCY3bf8olmiifjIgAFPk9QNlrkDDmS
KogkNe8Nz2a4YcF0o9BSsHoeu5Lbh8WkoJHCtnmCLMc3nGixsELMiwPAulg0
zH2uEbiAhtBsugkYjGNxIUPN4u4P9fGe+XGEHcfk1IVH5cbjv0hKEWGFWyMb
92BgXZWHAmGPjYBH5BrmN0jiOt5xL/DtkhoN6eptWSbYXeMCy4OWVDH3UNMu
KF+k5F60i6nAiaTddWvZORVwxFQhLVJCTHYWwr8FK9t74nku+ZbAWTbeuS8v
9M3Vpu8wbWMEQH50qF8aCrMcMi5QLhzKvlLq6o2DDGdhcYcxuGqKjuKrnSXj
052UKoug+zeZrcT07HMst3Ho59KbtyXXeY30UpYUEWY1sQOiqEi1CBIsIM82
GXEZ2ri0qNqQN22BekQHxxhUsHHdPKAM9AFWkYwpjqpHzKxeF1nkRTAXcy88
muv6U2PLbg8uae5SCTobN9N86rVLHBpmoP0i/lBLr15I9XIY6bMUUEXr8Q/8
1jkn8hp27CvFjnDzYz1UdGfWvCEXjCpG/2qcUCvM061ZSl2UARaaRtYG8gZN
vkLacSOayst8Fs2UcSucGRgNYKZ6ugxG3j+VAapNpTZFrgXwk97jtj+U9wEJ
IvH/LQ98OpRYjHC5N9PdDppWmVNgJf5nIoY8aPjn9N8NpYiVB+v5nRcGTt2f
TEayei+P0YL0ArAcP821klHnmw7n3lrGsqHhBwehQ7X9cG+dDBjabzmvBrEu
yJZu4UhybeAfIAt/MEEYVjTlVlAbePlPCi/9+wC/2yA66V/2FCOsvbaqAgOk
yLXEi+ipWdnvY3HZgJViakv+5UOUPqIY6NLl2qlvb11U1FdsHgMqQWLDQBWB
Wa7VqnZYUjQh07IEaJqFxzUv2b6JrelaRTlB+FJROgvXycmokq3ssIIh5q1Y
4cOyzv15VWJxDw3VPfUoh6jTyOllbcT1enpp704XN+M+FZZbSfTkbGBE5pHm
cepHa1v36sup4psEsbRL5ZgrIiJCYWIr2iFPP7dMOeIgjO0c3+XOxlxtgEv/
Fo8PdXBTnnWT+joHV7Tl+o1G8TTAFa3CheL5mtBhkQqkQoq+hm3l+C5mi/h7
vNCvULzDWuo4Tisfq3v5DjV4Jdqrc/szMp2vfXi6evoEWVxW1qYvgV3+4IPD
OrqumtHZMd/gZ+zygruAxpLF6E1i92A2Gc0bNtVLB8lP0nObM4X0QOVVNrKx
CsedbMvTMnpaHR5eRdWE8CLvpe6fY8ypTWm+8TB8+cL5LxZxRQ8SD8kYBs7x
P8Yx9nQktRPR0fthkNWzBaPc4V00F65rLLPE5MT86nJzmi5/DDrvQDU6Ezi2
gwIwEyZN0KkUY+lIsJFVQtghjk3jHEKAB6m4uLZOOwvg50QKjKGSUiVBnVwq
hsnDdU8wH3dVmZyN1UZt20DtStQNeHt2OvvIdz/q9m9hpal4ymIq0q/KalR6
hWSLD5aWIdS8gSEkBBFNbiihajBioSunBlpM/pJqRzihXT0w/6JxYA8UlK1Z
+zsyoGX89ftcb6/PoA7gHDfyMe4pdBG/GtCYlNWfRdwpSDAhRk/Th1QeU9vQ
Qpv59fT/m6j6FJfjWQvXp7bty/n3bsOV5kHTfSMFVDBhBeoDw8Q+ZBmA1oN2
bl/zXga1XDfhOcr/SWize7jxG53FalbvqR2N98tEAhwf8ITeVsb3onhdVYV+
hjegjxlEYB+W0NxRiEOvvfhZYnY1zI974NRORkQ6TJ4b2xk4HGn/jcRGnf3T
5GB9y/Yr1IxIneQ4n08z5KfvNMc1p9rAOqhd1IboNfkfI0YJ8+LZs/9kJnnY
Hl7Hkvtd4eGit+dQa0ZTZl3HaWG1kKTECMs8rHl0ga/5aN3jxMce+y6e2Bf/
+H2C5J+2QBj/vBizD9Etp0pK9EP8H52dx9PEiORK6x2Hho/UtF3PfT7u5vvW
ZEeSFQSRzubaOkno6bC7254T6aB8jTxQYtzO34naznZ0N3uOzZsfzq8gXY0A
5auppIMS87W9AzsfCHGDg8qzRzvdnDliDFFWjvs2TKas6XcfVpmfuElmcL+V
LG4tWUJL4OXtYt4KxK1w56wIY4W4Sjuozxqke/1i5lrJPc+Jy8MATmBZRE2Q
IgwSFRcvrILAGeV/3RmmE0vLLETtK1dPR97i5+JPbkh4LIHBHOgQ5wfXAPUU
LhWieFh1W/TkkC8svivxGcNhIBNvqmF2j9uip2632tmTpa7+oqww0c9660ST
B06p4mSmKfNGmAucruxZJo+HsDkYN2e9o6flguVeLcp9QBCKq4YycFHBLDth
/ZwDIoT9mF9lNSmfm1tSd9aijNXoiSovAZVXbqGh3ITsUZG0hMyy+lmeyC4Z
6hsQs6d/fwCNCxqXun7IdgUI22ElWVzF1YA1pJZA+JjuH7SkXQocIPSAPZvv
lVRt5VG5hJLiMqbBepmNHoizTGYoJLWzP/OwDwQHvm64lT3j3Im9NvZzueIo
EoBw5+ZeSATmHviNujRkGlXdKBCBG5CAHTOF8ecxIBhUB669DyGLiQ7Hh+l+
ZOZhjdiOPWLY3a8CSLp2X1e1MjllfHLFe4HWpOswQ4lrCXFTHkMsdP8m+O5k
omrhst3WAeEZUFU2IKb+Ft02zsjcuR8YNaoq2TznVJ4KQWg/gj4W6zo0nONj
lENJ5DpviLOh0UpdsAwkO/1qazZxh2yNzHOKpSONzEwl1y1cCkSCCRIGGmUX
eXT1qGJaJfZOwMj1mb5Krbb+SNFCtFhVSJKPj9uBv0dZ4/haflUTz+I3WY8N
j9hL/GNXfO+OR4VlJAXIZzBhuDBX1/PORvAIMvafpKDxtEEe29osKV3evTJ6
96E72yAnV2s/83kmJkfxmWpHEUjy1UCcrYXgt0rrZcjzQ90qbwiBpNKojfl9
LUu6A/ZJNbW72c8aN5l9vmWv74MuaCreE3oLo4FU/LN6ss2/D/2Ti4lpxl3Q
/2TFxG2D8iJMcWsi9993WLspsEKYjThss47qdXV4E81uW/QF/plJ0ivhJnwD
Ype6QdW79oi+UGMUsatkcplNzyYADZsWmtvYo17OE4Y3QLZK/Dn9FFdqlHUH
MzDee5aFb58UpuVDOzpRDYG12/kktC5CF75/ae8wVGDOLPmZNRLrfSd5PFMR
RSHGtdZiK0WE+pneJ3l2jUjpW3oBj5xKpBy1jKWnfI6SHEMfSRNmzhKdStX7
jiYpE/9Ye+CLhEV3FEidwwM+LPnnZIQeCchTujPYzFMR14eprspuvyDtI2s3
/dipNIKtrbULxa+TzSllRPVxVHh16ZUsrDS2PYdIUL2YEhq85mpsQGZV34mP
iCSbCnbKc5aMtROHjB93TWC9oOWdShARDGWrXFsUMOtnlg30PpRLLLjnJvaA
UVOy80YVwck0OUpsL1EiuC4f9lfugV6GKZ893Oo1M5gEiQ3X6qu1xnrDOHNX
+jdFqZtwk3duwEK1fzUH8/0q0wEJwYfBXoTYxB+A015lKZAWBX6UW+SizRAU
jgAf9qUn2TSm51wIi53NH7yPc20NBVeVvbd1z/B1pIZdM1R11wSrdWVc5IsP
pegVHVo2Kiua+vZN7zmlpoBmanN9Y3lRHUauxLov1uzOLI1yOrUYtrx/R+cb
P3LuhVqp38Lzpdbk550c9IuiVah5pS2JL5Ws7Yl+f9HalRkC1Bwl0nJClpLw
21MGsdw+TcxZF3gMvIzLN5VWzu3vG5QEgf6UB/VDSjMdAt2IkJXbWOrtHxnX
JO5HvT6CgYiJ8Ms+dE5G3+dsUDsQoJdkTI9Mn3FHMU2hn++Zk4nAYQMyBSC7
5lspCjS+UbZqWQrFTiR58/tjXGJ4OQs3DFFse4kkd59FzLa6e1pv4noNyjK8
aTeHxCc2N3tR8bgVkE36G0ILYLVLBxLIvpXPCZ4wQnOSBTzPIKlb7VutNlM/
61JFioPTE7k0b6ojKkL0JL4Z5LPaq//LDkOzh12dGIgfNjfCAINzYdmr20dF
pKdHDcY8csq79DW0Pb1VQncoj3Gr9bduad/CMgZTv2IZk6gVbTQuO+EUgOte
QsnDUoZc/M4BcGHqI2xGMx0KnqviYn0paK4Q8UezcGZbMNwuJZDGYJY9vT6e
m1G321yvl34p6+6okSqqwOJVHCCyH+WBBiqlbQpUjTgFmshFr0SMxk8hC9J5
c7asM8XiiXcn9o9CLxJdhe1ArmjIICDSUtO3TwD96DDrwNLnHeahuX9eD4OI
gZkWfsscL81q71qTida0szdSAyikFP9A6y6WGXA0SLYOKtzTX+y5q4LLss7x
0+Rk9ISJG6gpYNci3bHb9CA3KB+xwlU0rLbl1bRkx5m5kevemthmHiAO+73I
1kpuoGI1/kqjxXtNwC/5Lio367+zP3JtAF0urIR73SIZ3Pw1MOvOhu6fOyqB
g9ha8LVn6voYcH83tAZ7EwaBWJ2A/ayOimYIQCquSKpC5XpDWy08InNi0Nde
w+p6qYv2JcydEFn/zmrk3rTtEmcFwbsrwvLtP+XXOEjMHFEAASjbZx5tRqnO
ffJ1RgcgNuMIy+5usVCpS617WZsTUkJ4q7ne6cQn0x3rxENVDozNypfgnOSx
rqcS77CjtIqt2P7l0tDf0keMKeTwj5ptp2Qh/oqtzpPNJhiworF8bTPBSjju
nYMNTtqtZ+EOjrxkGIW2j/lCfWQ3zjdhgKBz0xNimo0akF1pKuisJAHDPVKE
flILo8Qt5RFsS1ZXuDAlPrzCA9NetH8HXBMHFs5FkxU/HYMf2pozLHCDZKTn
+BOMhQOJwJKfDAovoL0+wj7RxtQ0LLlhrLrm+Dw3T42O02wLKuuF8Wcu3wCG
9VidaMFkHXWFfz4HY+1BmLQcBaJmXMqYAe5uFlUyCnVrivWeuNJ87g5VSKUM
/HHJnin6+GzCzPmB0DP8y1PLgIVq4WGapBZP4W2ypOT+JcCWQ1t+J5dJNDMu
QIto5yqB3Rtl6VXxr0ZrImsxoE9ObHWrpfKYw/cjkguuI1PveHl955JU93rN
KFwfDOBPR58SX+4QBglH8Uksm7L+sRawMqDcDXMWt4OMDu4bKDSZcFKF9hsD
lKUiartoIQaxlEhMh6/A9yir7+beRbTJI6D5MuR44IKSvNRva6wb7DfyemwS
nI0qXeRd9LEiLzz2PcJCTaQ0s6dkN+GJnSRwdXW+8FtW8UAvIGGxlaDkSeb6
1XQytfEEFT0Hks1ZOCtJ3sAlvaOES0xzlQdrKkB1wl3o4GdLLKkbvlqZg8h3
r9FEjvYCGab5f3BoxDvdAWd4PcLILE3s7HpjMuWLqwn7w0MXU8SJ8l1mrkrJ
FxX6k0ISosSsE/xWOZ4/02jA0Oc6UUDGrToxy7ezD8XmMaX2jWeO0u93FtTi
Y6mXwRp/fHYBC2tjdHxJBeiwrA4j/lnc83zghAVn84+NSeEFQEqFyTxhYkbf
iQLK6vVXzQzVrzFHsMBV2Y3BNaNlhmDmj5nY0nhSY97oPRr1AfcsVdAtTZ1F
NGHr18x43dQIcOozZKBk1p1L7fqGa+CoexYKLS0xlQqhADfI44FaoiGmk0mj
DiDhPyV/0STNMhIlPQmnNtE85ZU+E1o0EoHPKG6kFf6Zf5jL1sZjwXTF5dXU
Wfd3kJxb8G7nqWXL1J1OLXSu16uRuhVH4cT1LVUueLvr6fHsDP0w/fUD11BY
8Fe2pw/Ckb70zfyOFP9bziserVvwavjHFuW9y6d3cg4W5zWMAJKQxn6AzMlW
DhrKJ4ekv0CtSwXYVTKZ3Pv+a/LbV9zPh7sD1rrtq20BJQyewi4vt6Fnpf5v
VQrcCh5LxaeaGBUd2dP7qD+Rrj8u6dk40tL5aKMCItpT9yHcKH7RbRGPGSVN
kJ7M7DbDpVKpTm+/bGim3l7U4QvCN9mxY+O5qZuCZH8W76bvs0pOYQxZAmkg
wvgMt0WULi4ob0lL8SNcpIbULt+SzeLEWuChSt3Od9ZGfFaULvRJ/d11pN9H
A0JbTsIAQHvYvKWFHVmGPWi9rRn5a1t8JImuhvy3p2sRh+6+vKvXlmRQhmTL
RHokynmDJj/Gzu7MlrheAZIPlAWhHGWpUXxWntB3kbI8/47oCF2akfsdUId0
XpFTHjgJ+HLHfggyuXUEzhp9q2dboGdzwhB/T8GjP37QQnI+J/RptBG92L6u
ltlDaVd5dr4F77Mnp7SZbcT7RGEtAauMlrHle5P5bm68sBvmLYVdEzo8xaUx
A9e58SHabArLqXLxYcVKPo4eCqpGZqIYh7YKS2kidVbzPVWrW0DtxNCTajQP
Apq884b+HvziiePjX+V0b0eKH2ckQv9ueldn1xbsRhDP5fV32lOU7D1U/BXr
o5qoU9cG7+b8Nn+Ym/vHXOg/LU/XdoTZBFGPk+yz1J4VpwM2nNjLKMgKhE4M
SYQjaEr6wybetfXqKlo4U3qDq/tO54MMdz1hEQl0lOaswFCaKGaZehwm3s6/
VX8I0DXKV4nfcXpGvGL9Fw2h3I6SKqzaau12QC33H7DT7Oyy80P+zLXHHIOy
nPUQbphnnj3fnSM3l18fIFbtHQpOIFUMtmYgK1DqN7BMTJs7O1X+Ss5H31Gz
u4ar0rJI6P/YDl1fjuXpM6/gC/fglzUKmE5GFxss8AXwNBiI+iICD1b80D9W
BHqObWRgGHNzg/Vk3PSmw06Lh7do2/2KHmYpmCy6p17IbpRhqxrGjRWr+4Ei
vH39umhhc1CrF2NEgRzdKMbu5+v50ostycjGG9sjVUDOH+NprtgP85jJKtIT
r27X4DJNcNeaUcwiruMYFdodv/9UNTntE75L9bxwH956ZhKZ5sX/bC15/Z1u
odhc5WtlN9ayM2fkKp4g8+llRNf6udPaivnFzY9F71SbHBVRYE+zLY3kvZJ9
GsGUM/3hgx781U4j8EUJOKJ5egxdXMNHpFe9cm8xvyAvxNjfVdMyP+OmCEVK
vZH2h6UyteYYHH1MgS7OQf/0zuU3bdbRZRcEIVpclIL0FdE1aaBpJWkTRbh6
+P63x5lSLnOEY+Jae4xp/fhR3QdIIeOnw2f9kvMniHw6e0ayhftg4jocPg72
oBCTtGmNysGlb1a/hCES1QftrJPAiNFxJTSafuSsDSKsN3gfOpaATtavzrEb
cLPpYDuRxQQGgTQGqI3w3c/d0cVlSmB5TZbigU8eX0RdItZ6qRw6HjFZIdn/
pNLpebTV+F+SNZqa7xqu3gEENzL1GFZoaXiLblek2v4h2jXwypAAX8RYtb/X
7neFHBIH/WJlUcfw/0HCwd0rqZZXI2CzlXJo3dPjRoeKOAHrhuA8Ejtioto7
wdJcXAEx5jDqp1CCodgehBV5UtuzodHPvpMCqTE5yicVSHPJaDP0c1H+KuTQ
8A65J+CuWK5U82ZW4YDFnq/7+9Om2PxRoHy0nfJyuwAeZ7CCdmv2xdIcLvCF
ctMzu/JDR7n1ViO93CnemW5nOhgXKTx/KuguqrJ6t/ROtnh5YPQiXykoRVPm
baKsRmfig2CsJL5UxRK4iQF0kRmx/b0Qe4+pHf8AD40a9vCdglTyVxMyzHBM
P5+ijHNVpHn+d2woUPBTU6Tajp13DxfcFiaswTSZ6i7v8LTmbWNAP/ZU9Q4d
DUzAQPuM9t/AZgJwv7UbqC4GaP4ZLQ6tra52osWC5xpV3x/z3g7VNsDwGcfB
iLmWG+rBY1WJQYgtIShSn6Z9t2FIXeTvdwNUgqRTGgag56FIwJlAQ1+0Oe/X
a5SgAs3zYKcJzgNME2t5IOkY74IdQ77JR6hDMAqWPo0TS3ZeWi2TrFDhFPAH
XgYf8UGWc5lFe0vi7n0MH7O1GeprUmGAcM+7QnvStoNvpyvBLM3b8aEkMLGs
ph44h9F0VKe6KCbzFOmHDaTjHDEf3EH0B+2br5Lb7aGDlT4AWGLbWF8Wkf2S
x0IoXiOF4G8rNDDqFkYg7963DMg476iQynN0kCmff1QBq7zZqWHOSyCMjNWM
6bGe5De1opaHAVW2rmxh5Qj+Ez9G/FyTTa38gLKLlezP/8jwGdPDKzE1QvYU
qU8bZFOfnxQGGoDEF7vS6os/sXoFJZQXMb6/SKsRwLSHPRPNXO5eoGGvlaHu
M0y83DcoYgUKtmD8KSnvSYhtfk4HKypZuLc4YdWS0a786wtvTpOe2y1F4e3s
RCcpOmJiZNW6TSGIHpo/kmvB7Li4MR3nl+9FVSKJsFMwppxcKFVYI7Qo4ufE
Eojr41OBAkh/tIiljTnofFF+2skWeeMsCiJqiGM0/5rQjX3ZW4OEMT3FXBo7
XiiwL/+zjqAto61qjHMwPq5K0cisZMIXgBipMRNEip7yJmpYFbmkv8ldNfqS
JC3Quxbgzp5+EBR6+0D4YPB+CcT7nPsZK8HZkcNw5fW7PNtsehnse4ppV315
RE8fq5NFAeGIc29OinMukYhT3biq9xjL3pSLl+5R3x+o9lz/8gX4O+XmDeZx
jwwN88mq+y7ZQvTOQDRKje67ex1sIeCmGBkArgC0OEUBQnNRaL1HbF1JFH/f
KIOxxrbSOr13XZTcKDkL3tPX6NIqAM02WPCWZ/8EiaJ95k8KJp/I7nRVOTFE
3fJyz83Qfg9huwT2joyS2YQJQdhDEx2T7YiLUnuUzWk5KLe9fstI8TTnn3qw
1SPaaZc/cn5o5IiLc2EmkWxXr07dEe6oMtIO6G3AxqXkqeBSJq9AwWBZShPe
MGuCGjUYcpJi8NcTjsTBaWCytNu7t5NMgEgjNT1DPycERJmVkvxaWmwFR3HY
oLlp0MS74WEmfgShvWQTEv3GcF8E60m3Oxg58XF1L9jC6fPf7IutTufHv91a
2KvGVl/7eabH1Xt28lWfEG5JPjTJoEi3dzwwe3pA3/+uN1VWM55Y2/+T8yWZ
ZyRNxIkwWSRgKu6C/6bdUSNgBh4b+khTn97qVJdw5BiFEz/TgHWzaHWMucEH
Qvv/U05wkMJfLf3mwrB9iucnE5D1WluvlQ6ZWOiUmE5tEx+hA2jUBWALgRT6
1ySoz5FXwTfsgEH1Hh5fXAXb/2d7VXl0DxonJlK4S/8GvHzu78H+zx1G6hFV
r5bHpY8QM9DnjNyGvnQ0GcGXF/SRHrFLGPe1eqQfRF6S+jUwYucHRmcakGF5
p8ZnEpPClnNP6fWMa4PKGHXlWts3VOtPlA1VTkEocjTxJeYd3vZkakJIAayO
Daii/EUbBEdsFlI8uu9iakcer9L81HE3v9H4qIcDs1S+tk9GTmFzVeSKyCL6
7EDZXNm3V/T1och/sOzGk8z7r7dW69L+4x0v9vtY7h7oUZ7bpEzvGQRSROGe
RsQgGfNjF6IGd9jRqmfQHN6z1Li3rmDZG/lnd9AMDV8YXnigIaKjRCmNTPBn
sq2K5LgROtjCrHBF/Kx7Bq2PTzSXJyUG6ojkXZ9vCu/rcCB10A7SXesUQfpC
XA4+8PxD/SJXVqnnBBS3925/q+w/DGVX9iBaPwbLBzcT4Gt4qmUIJFsveGJ2
oJU+dFsMHkM8vbaziOPJEvbo4S/ru2+G9xsJFabYFxJnyBVWVzAE8sCx7HaJ
CZBKdD3XnWWkyqx4aLuikokwVRp7D3B1igJhn49Q66JQn0uTMi8cHS5OYwF3
rsQetOywVcrdLtNWJWrV+TO1a9tGWnFC40wwA/23ajbo3vWeQQiuwtcdUj9r
0AKxx8LOXp/Gq5QhPQZZ+s6acngUu8I4nWxmZ+/RedDC3GjM0A8ndQersqZH
rmDYgEqPvPaPhH1TO2wombRqOk1VwcdxY8xeKcoQ1nsW4Mhh/i2vcvPUEhGW
QiplqUSbLLhK68ncXYYlsy1tWN+CREt75d9rEL9gwARVj/3VyuhdnAJG3y9U
wmCTrjAoZpZ5Q0oPBfZMq84x7M/B0b0XTjZcMsuK4BpXFOE4Yy2/Yed0rvea
d625RqFZ456q/sK/JWhGScdgDoXSB2XdYjXbkcUtCpVDJiHsH1PqqW0+51VV
cii/LpT1tcyZqeOsRr8JGzEdMEpgYa3KccecSaWbjXtyvcuKshMAODCyA/Tl
i7FPtBnbLFMKiDf1G1wReD1/VgLEvPevyvFgunMoRkVsZoe1/tewu+AkqHOh
wQZ5P3tw/cpUHkzQk6dLsVDLzwFexJCPm0ZEQ8w0gwLIlg1CmMMfx2R+0hZW
azcjr/8cU+oqYCzKVmJfh+OK+beqpk1/IAFcG2j1vEzWOhkJBv9yy65fiR0q
i5xwrdaLHFfQdYz6jsWMDENpMRchEdjE4sEu08t3TczIQMi0c8FULVF88EZ7
515uDfgXiqh00guhr8uK0MNnlb3eX5xdkn5bk8xMAhCCPN/XChiVWR6hpKBw
6/dwEE1Cn0ElKT/FZj/sx6I06a6Bl8MXh0xSChFsBT9vYZVBepipo4Je9ir9
CNed6l5G2RBP7M5eseI2UPYJEwExNhRT5duZMULrqkf0wcwJimpEWHg8yLjW
VIjZhlspbySRtNYCOCbfMEKlKuEAjeec+iS72+KYDRit1epa7p79NsIWoFJe
GH+2/BcD2yHw6zmrQlx8ukoQDLb6qP+xvbQbLLmmu3eKO7zb+KJPU64LaGFq
JV//5uReWdNXwaAdhXac5CLrkofC0y5wHlgTqtRFKXR9+8e+LZBheypK6Tzw
ISn6G80ZzVZibTSan79vRiEmNMwy597WOK4DUT6lI2wWwpKTA/dbd0U9iLkp
VtBDzan5tliZnXgjIOmP73iFK3N1xmaOK2tCad4L2Ix1GC3kIxY+HeK+Jtw4
C54UpC7JSzgbi7Y2zzV0bdJWMHjYF8Vry0PZca8orog1wFWAHpF/unJ7MoH3
aOuqGy3oBNcMv27Ys+SXXUY5/mdTkwpffnZ5uwkHq2Td3HpTp6hFudI04mJ2
O7G2mFVTxS72lNPtScRh1/nZEmRL49lxeCiWJKA9qk/Tn8KjUsSQUq38ibUr
9IWeetQE+qAlXad1GqANVXH9879sO+O5tIgycYYIWwFy/t2s2YLZil8UTj2Y
nVOlf8WXQjzvl4djPQ3iRfxsBS1G5JQyzx3sGm2sucAwT7S+GDcM3ofdkt9G
h5lt3vfPYoFQXfBgXkUpETK5MVUoszhDiHtHGvJkiGXENN7qS+s/Rv2bvKAg
/JkyfQ5Li53L4vEVroa+7TotVA==

`pragma protect end_protected
