// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Ok2Zd004gL5BEWagj0yYDblOO7a6uwC+ez83Mjze+GLnitUAONXGNHR8/YxDwSPZ
TT8pRynfKU8tctEvVlihOVx9bJTHZSNRxsENuB1fD+NzE7DlI2HLcNT701CCN5YF
yrGHy/wfDy+B3cVs04VHPrc0UVgx62VzYJZ9owzL0XE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10288 )
`pragma protect data_block
itAJcBpTKQZDmSiHGjQQkSyYPXaduTIMdxO/srFp9sQyg6gnp2kf7UdheQF9tsXw
n6OdwZ8qVJqPqVfHGbr0l0Vx6U5VfuoS9I3b2zLRpLWOUaote8G81yUv77q2d9vV
yVi5rctW59V87bb1vrNM5V10ydBpe5Bsb+c1RTwy5TdsP2TjK5YcZUkRGPX7/U8N
f4DJikgM9idAtww8YL5OXF1YL93UX5KApfgeYTDl111OUwd9Whb98Rvy2nT+jlda
3X0DfNLV1lA9E+8NNneU1bF3S0Zw51DCrm6XPSUgrsq7UQQoSTQDtwZmqKsnyhIY
wUHm7eMz6hwr+El8pWAg77E9RFqWZmZzJs1+5HOICoxgbsR+T6A7PQZXh5tcVBVx
KIn9vhBr8EZ5ADrFZGSO8BoUYa+Hi51ZN6c4bcSLwqklXf4WqcfphWYOrEZU0dR+
aw4EDGv2KdZu3VVk5Zipppii6olOh+q6UMEqqM6vL3JfnUct6Gxsq6aloeGeOESE
bXeR5W9HdBeNY9e4njpKrgGkJ+8qJ12AtmCayw8IWte2jGR+EWmWoheGAHVqVV9A
64fOlOU+EIv3gtDWTjWSVuD3hbw8U3rlkxEo8jjj+vuE2qmMgO5oy972VeXCGIM2
VBf7l7w8LxcdHPumZjxh6xDWQ+TpX7Gb8CjJgUnSjWV7XF8Bkr9KQDA/EPhLMIkh
0NhuTib9reu/hbnoReovEwkEu3zE4WzaMY4EN4u5C4biktG1ycEfdqtrN5aTL+dX
HqEOFY6zFPzaDvUTihGpGg5qv9nek9avovitzkz30i7JELoO4c7BYFgHZRXZdqoH
9PPCcq6v+o9LlimrN7sVmBovD7ksYk0L+aEI4dks7WYKGOmFWocwJtx8MIZoPUnM
Jx266EYle4GIqGqG6Z2+tHvVYTamEgkNT3gSknVGlljgPhOoqR4xJX5sIKui9KOa
2GFh+PCqP6GrCqiqEGf7FXdGOFM7Rjo4qE5mna47JoNa//lk8+Yq5y7oeQFuJ+xy
iOwL/roCpFu+tCa8+bswoph+ny7UevXyeg25asz7kRkGRiJ7RlJ1N8bPUyE+PtqK
PDJ+X/IhqCTsAwl7kOUOcTKojLRpfiRlmITkMpWNGovPbHBqksd6V0PmOSnLUz8e
sHdnTbAFFglwJRuBe+CjxT0J2dJ0eWj/GLyWQMPC8fjPvQe7Nav3b/0CRGR4Hcgs
UnzlCouECpyBk8vKd1QGHiQZ4R6cW2ssESQ57kU7wGZn9NGJnpj4qbDPbri1JVKL
YCbWuJ0x1wRfLJaB6wKxpEu8G4H1IEzb5/fpZ1HkTKI8qPGp4Mru6d3aO5mZbHkv
1k+zX1DtI2m47iPGAl/ZvbBijqpphPI/oVGJkthnEDORWmm1sIGhNOZarGOeETO7
ODJNb19T720qfIYudM3tau8D6iFUoKAxKlaHRvoifvxiIGXRve2+9spTuG7KDCQx
7zinN2Ea7FnQGn9ITW17gTibgj6jnztsZ6y/eX5NDdPR/JbCsZTy/AVHdTEXZ1yj
bMVgx1F9xzjHmBxj2bRBGcBAWTebPB68BUG9hMVrxW77iDL/s/ZgpdMM+hQhsvMH
r5GV6p2JTnct5UDjSKNO2dHXcVabDEyTKsjQWflKAopS6WI1ZDbmwM15hYi97uNq
vf6mgNgdBkgeECfmjXTxVkd2UvXnbSMug6jQzZVkEEtgywddOkxh47nwrdstjbbi
tPBknn2XG7edL0kNRWZsY7NzfPu6SS60zuEHsVR4jvNRqdD/Bn4jhfbST5T4rTuY
ks4sYJwySuaznng8ad7VC2+eeptmntrsfczfpe69eDiDLh8jEf8fdrjUOb5xeD5i
yQkisSHBRaPtkyeoZ2p7S6dgR5J3Xc5W66V7vocueCzS1X617XRX1QXgnHP3XMq7
hB+HUSnacRM++OJr2vrR03HRt65xj84Z5JWux/WrjCw3timITWSzifxnmo3+ssRv
2kjYHx8jKfo4sHG8HeKf7rVAyZP4BkuxdgV8Aq+n6rP6KM3yy4llgZXbKGi+vFqn
lalwJwgPqp+01dgdt6cx59TaLoHVDllCtZRgqPtDWrs1Vu9vlNecMQwIca6/Kwve
p8IOuLYtYdXnDNZ31abZrFyRK7SnwKHkKUmm3eVtFTpDV/UdbRhY6A92H5YHn3tG
TBGvhQ9Bh8XXq1tLIetSgatgUGLel1UFMJ8i/fDQVvBOj26k5NZKxTXTdkavOCFt
eTMCMCr6djMKLaZpBSu3E9TMOtiaZSZs2NDURir+KLcBxBAvFbxmOUd0SbRdmhi6
Q/YSbC/TJKY//ZMf6wsJ0g95P1vity1sVYVufx24VjpM0CfxK6W35LOnNz0kTdpu
UPE2evlmD5rDbZTc5pkC8Hak22MdapoIdMa7TH/wW0j1YlSXR9mIkKs+T2z0K/4g
4Uy4buJmAFxnorNhGkgm3C2pXd8DkV9myws0HfNlY3gZRGHTcTI1ybiyAyJgpOjm
/wyE2D6PXVIvfODXtrcT1yl4Xcdr6JYSxKKtUsaQa8dVdnom64Tqy5zTlE9cRLuG
IQqZv5/2hbcna6wWviSI/kP8p+l8i5JVVwc4QJj+F+EyCR7PjU/7B6+yCcOLv4Tw
lkeFQ3U5r8q94j2aFfCLfOwIMLoj0EF+AtcuPmH5yS4QkoPl+zCPhIq7m2vr1Zyn
fkeZEMXJKMSvdIfWGf6G6kRPFmA0xvVsbusekPuDTpxv4gfO0tm65wvA+qehaQVo
ZMaSpuASjRg3PJudS/gMS4IQikdsgYbD3qPMo0zOALjtZRg29fEQrjtqlsUyVV50
L1ETZC6JgxUb7EXMwHv/lKmu+pFmxB6cPjkLOlMiY3iHYUlp8jAJxOljjIwTeLXO
v+VLwsLwJk9uzwT7dCcpvHCHEjWngYXGUNfELzJi7THbwqsDBh8WeW0HnT79x2/Y
QvSAFm8Gb6w0Iv0ufoRHW8Hqf6YvhvB7dK9RkXcb3t6jhD9MW6t04Cz5Dsq4ylwT
Mm6AjmdzIn1FsVbbEey7FoCLwnInyR5Whc9t4I1SijW3UE6gxbTkh8BVXNs9g0eb
JAu3zuqIie9+xLg5fXx4ZXlzEYq/MXc6NuRwAslXJZ6ZOKQWG1FCtl5JPCssFIpu
2ytf0lBHxRftycjhB5A8cNBL40vWZUSeQZ4UcHabQD+HeFrus5Z/6jdN1eQ+z5/3
gFGqmWbHobLw3ZCH3mfDmQg7DJp4J9ks7ZylQCHGF0vZSlFuWLtlPq0a7tXuTj9I
8X2WM74Rgf0mfZTCbWHfXlOu8FwgOYW7xhwJ6mFQICMz+00gFIkHuP1JGmtIaIMh
fE31vuspenTAwrNKqjVh/J8W/zaxsI56IGYgE+381D3Sv3OjklJ1/pYhxRBoXu+M
c6li0AZWyjbWWaMQ9HbsWfYJtUOzjrXQHYGRfto+7GYwrnDzQowA5EYofKMJbdse
nQWrjP7uBor2iQj6XvHRMShrAtN5YMr3tDtBtG3ABocoCaDJX50X4eBMBUAJFKVq
DdJuAQ72/49nsbDusj0sw5tNATepSz8i3gkZQokUun1cR8VhU3EGPn4EObEeqmgQ
4uPcCYvwNGHZx48366c5zeWWfL9718BEAzAtYZyS88s33IdF6Aoghbgzt883V3Z5
oEqVFuZbzYfxMlW8kbOECOKRGaekMi/tqEtqmlatvU6hz2tRMwE3s+o3d79xdjH8
FfgsHtNW80nfWoIk8+u2QxSAXzVf+nV7egkxAE8V1aT9FgNQPuCA1xpKEtqxpg1w
uy4GTgR6solAPb6OOx69vC85XN6tY+8qBc2qO39aguXJUC3G5lrMfBPAHRaI9Xxu
TBLEF0Q/i/rOjgJm2P3U47ZRRp+i6IVIKbSmUH27o9Ln2bMnQC0J+5gxqRVlo3ut
6HbQixsLlfyTN28ZaTnfO8EdmDQDv4rHrhYGAD+cIbC82/NTl3dp9NvMGR8pJ6AX
JbQf+2rEZaRtin+xIzEEQuTKcASX/9vMjZ4GeZcYJTo54thczJkB0p/XyT07Okzh
2uM3X/lIS8x2zHH7ZroX/e0XCRPcATez2SVti3x7QvzYC8/Qh4KvB7JgkE4aZql8
AVRi+tZOleus2wM0fuWZACBckYiYG6rQcjEcfpruVqN174wAfPFngHkszFnpU2CL
Oa4b6OyrnFPJfuneQt+pEFZSxN4ePiatBD9w13Yv7XtSDI9R2QYvQXkUzFXaxF5a
niQFp+GGzAJRWxLKgh5PrCpevy8fFeInUcg9hSqP8sY+UMlEIC1zoSy4CJ/hLGYu
S4bVQe5vNNiw/iibR+G7x6/eC+OCXQSVqKfv65wGIqdJ2/G2BstgDIXG6N1hnVB7
exyeT9xJ/C5uo3h0JjzTxTj+Cip6QhnlfEJcqYal8RUjrWd0tC0+6Is8xWszfV8R
Ne6AfPRtKFoU10ldaDDUWV7fgkVGsNVsvHL+ewIPqkI3147X9kxZF3n52po/NnjY
l/vKNdL0Jatws70coZ6zxxOlEBFRsA7XnmP5q8W3litCetYlJ/D7o2SbCkHU0hoz
XyhIiqFL+/ZWOpQTdWwBYRt5j910jDqyZBIDhSFLfhzT2lzbit54QyZccsm5D+HR
F0mMX490Lr3piZyauC8mLtK8YBHiB1ZQxIuZvCdcPHEQiGMgJYDNTgv5QVBuBRP+
ouW1zF73PBdKvTcDNoLvbinacsVLa+DjFgqKJ4qsqtVHW75hO65QY66lLdFaFTHp
WciogPt1N9YahIyDEtKKVom5BMd/se1OA9CN8wTvPurQP33lk+eO6958sd9LmuUp
oUzG4mqb7iEQfrMkFSBlE4FtF/LRiqgtsltDLS8ATPEAxGyR6784Nt7jQWaZ31M4
DCHRnP3wi5EqRSEoXNurLeIxLZvH001xOasxW7a4kJMfc2/O00jQTDcXdvNGzX2g
2EuHjl23WuGRVfJk/Jwjp2nvrxaEqMN2ZQSLwB1cOzrMt5T9XAHNntpjmYevXAwd
VMT9/Ogwqb9oIXdTeRu2rGREw3pHpg3cFiXg1GCNsBynFeZwYeCkFeZu0UE9mDcQ
71W9X9imye+QopFjfbdjj5ycoUsDKa9HiJJNv37rYKmHhJkvwGpMnY38t7RWBQIC
ltHhBWVD05TefwgzGpWkTslqucjWIvtztxw/IoUswNFUQ7eYsIciBd29hnEElUQi
AHnKWwuL50h69qA9Y2JGiewzjPwULcwG9+2REMtjmu/ywhXUGRP0qFWWvk0hgwmK
Ic00OICte0l3Z495v2+CcO1YYc5X0f6wt7zdzpl886eDzSZmsnxvZnCPTNBH9E4t
uupqDv6XymXD6aKnZ6NWhnAT06ycypC5aaDAHChftbLiFp2DCehq2hmwIkzt2y9q
lzu0Vx20pq6t3xi8FDFLrjHd4b8YSv2sfvIuEiUecJFtVcY0cRvjCEMB25fGE7Yv
oTXrVcSCIJm/7ydgUFc7isUGL1YACj/Rq57BCnnUoTLVOyb4xIvfE5UmNaBw35bx
65aM+zrhuPhK6srT+oHY/+sAMvNmws9yLhvUKZNrrBCwe756TmGxQ6Hbex/KvkhN
LFPaR752trh8JcW/Tz/1JOg0H32loA+2y+twm8Xi+gLmOz6NetTkg+9m2tff0Ije
8vRnFszrobFT0jR+FGnimMyeg7IX2glCxfgg3ZBBtAA3gd8y72CqnnKP0pSyL9jV
qLKyc9kR0r6b8OjDyKbV14qRG6BFvWf2LaojLoZ5YBeOlnTg7r7V4KzRBdULPjI+
AwXpe0gtvQSfgZ/caKmqlMItLijkyJSYtu+0fS0FmNYQBd7Ct6RdBCd7iUeWzmQF
U6214a0S24fKwyWWBVljxwsqkUoTz9mqWSmD0jbfjlafn1jIc/IHILx098paKFma
PymE1cuY+swiYW3qPLy46HqpWImLmmE33S8ovHU41Vgpdhmvk023b2MoUGZcT4CF
KCsb8kmqWghYRQOTr+TYubGomUn54DUJ2Gq4CVFdMV/9U0UEbOVZcs+Nfc0IglYJ
abQx8ChbO7vM5puv0odkciPiJq/4maETdwaWqVFkq5wprO9zoQakLI0uENigv7Nz
82//gjUzzVZXFcVZ04oIQR0YpyKlPOIy6milKr3Wp2rf/lG8lIafB68WwjOuCcSy
RvZfT/wHETpwIBiQO9VkKYtNV4Bl/MrnkUApiGMUyNL8hFvOFnEf1sKcpcQXQ1g1
OxduMZqvq78ZZKWL0tqPA9WisAjG2YW+9fO8dbPv8H2aefyrOv/SLv+46FBcBnO7
FcGPlDJ6G7laeAQTtiKX4vZ1/AQN3b+2p+z6A88DdssZJB0qMknqYHbDYSp0vBnq
0Jo6ZajnUiu29sCbOGwkRIRUNHBvEce/OQjwQAT79ufQs3kjidWR3fOBkAY0TErH
4avyN49vN2zMKyaxAabTK7HcNQ89RmTree4Cemwfnm4tBab38lS07NWQt55c4Hop
Ia4X5ZUnQpuQ0X0YU1zH/aquDxS/+L0yW+C6zcfXd3iCmeisnNxzDwn1u4dwIXo1
IsSGruRwZriJ21LV/q6Y018FWO1RGVN+SmJgtTPNh1gBZ/NxbJWY2j0LV3tpj2Jz
d1zG2Y6eJzoo6+OPR2Uh7LBJZMK81ttmkY+6k6rEDBL1d8hvyt2+5k53snIUqS9V
rSv6AnC75VK87c1wQOIcWuBzI9Bfs3ER8Wu7SMinpLG3CMgVe6TYxf81aSxc0w2r
8UH/2UOb2h2fBvCEME3uYbjUUJWRMVHxeldcZyaFnofSmLVlwwRF3t7dr02VBFEx
vtzhONpbo3zE6nfcPWhXV9qrqnqQj2hsTd1i78x3Hp5fdPzxVkyDTwKQcG84Qrlc
Yxbxmw+m6TuMSzoVmPH2lEl8x+UOOYKG8cgVJhkqmjG2KugXVWGpzswFJqmaTlCi
HYurI6OoQ2Hu9KCzou9Wsow59CWqY0reHgvJxsnOs1mC5Rl174cpySwK8crZS2fg
dv6Wzte72FE4iTtVRx39VjWkqFxsNDCHdbR4p+ZovyZVpYg+OMj6uBbkJk/lS9lz
Wx4KCiIqxiX/QLUChAV1sfARVqI6jNfJHHnUdfQRiQAXdS+sEoSH1U7xQwj+IibF
eDjK0SL+ZIgHW2P3VpEoxrsziO90bwyVWu9y0MAFW5ZiqoLCnYrgCb61Svy4f5CD
R8d0Mja37FWIQzpPH+ySvYHED7f/BvlxR9ScjfEQCOrZl4mblNcL7/vxxJaoKrN8
znCep+yvL5G9GwPfs0+rfhHjUv0lxSlweicp9GW1Hxi+wV9sQfqOx6yjNZOQ6g0Z
UMsJ+vSw6sqpTF7MF4otovR9TqJV/g4lftPMQZ+MqwSlqfe2uW7qYbG7NS83xHC9
4BWeTmzvk/1dWlgfdaaW+3dcjgSf8cB5lvZbn0QyjcD/pew825uzF13qbJdvWqkd
zjJq0yYO6Twp2Ar8QubBiMzA8NAdxwiH455DYi3ABLH90CGoiGQlp+uF2jBHsq6A
Z7a1A3HmeUOO9/KlPE99+BnpEi+Mh6RIDgvfS/I+cDeZgqKl0ZFUkvwoIbx/l7Eu
DOLzY0RJ7gUCMHJvj+PXhIBcaJZ9+wLICLcI289X2BbxIGXH/JOuTvyunM8YMEEc
puH0N9FrV22kFkoFk8G09LLzS29UgL3IjQrQPcDnuKN0AGyCny7uCJRVMTYNlZ+m
Oj4sMWL+4pnFm4RiWjDeqzBgSOiTixghD4tQ7OcYL7YyOFzTp1CX9JBEVp+5WGRM
f91JXUZ9du4qQvkHso2Pzb10/BZa9zgC3UkNAnkMUjeiJ8styybKwF+2Go5FSeyR
fH3I5GeWhzEADmSw6Ry/CKdv5/x2Vd0attiGGwihzIZ2YiI+ecuAeXqg1oPvUx93
GLep+F3NZwLf5pLtsi6VZL81sFErdCkVJRtNrVj1/G+AKyk0hWNDf+gsp39YLTFS
xYiJLokusKQ43RAVDeyigjNZLwF4ZUzAReHxTMW0pBViCbBVPoCIyM94BUiGS6El
KgCa0yumeALvKwE2uRSNMcj1b09lJp6D18sX0xIkQ3oZ76QpIEZDKMDHJYqMjGnx
SgXAKmkCRzrkx8tE6dajj2HTK0l5/YcWY0riGJaIIVW7nnN0W+a+BbTmrARZLyc8
yueWxnNTKudlSctTN1jE86lzSqWvyQ5Ib/NH1gDnFR7n8HR9xqk1M6iZBO6bz5BR
aDNBesKGMPOtDWY8zSryL7keowLUCod3uAG7Mz4xjKqosP4453VLkHEmAgzkuyZO
tgfoIsu7mgdgV0ZEVzWybE31XnRMsMw8CsGbD+Z/MfjQRvgvCTLBxKPviRBghRRJ
GSz8p+TCNgUvYwis3zF+qcwLlv91bV+TpxXGAYGx+B+1cHofgQgMIK2NskNxJR66
2O+xDhS+TZ0MmnNsxj+KspecXA6invH2XXp8Aug4AtiU1gwY7YmI6Pp82yjV1z1p
If8D3dRVpgZrWQJwEsc6/1Dw7Zj3mqqIGvd/v0hTvej80+ngZ6h+Q1Ua9tzIwZtR
ZDeI7jfXUrv76pZAvmELXncqSYztXeOZoSsAOO5eunQfQYt0syrUBm8fi5wtYIYm
egmn3Vpw+j8iGeDDZ0FolS9E2tyd9PYjB6oPcqZQHZQGNIon1mPgdJM9MlgFx9Ar
RHWCAbkcg4hGigxndgAAd8MuHD4SFBZ8kYC9hn1pI/jRwZJ9M3QdJ90Wp0Wen09d
xRWGslrrsnpGbeovEIhQHk0qLiXJYMWTXw+n62FYeU0tOIOFFWk4HxIdWfI641la
CyjARAsOihqEyHx5629wLDUl2RZOjtlSNbb0oRqtfHax2k9XfI3IRElMlHT6DkDX
h04GNsTfxECxS1zvtrmjvLUqaGSmeOz2sCn3IG56LU5dklnhByksaKOuVgcH6s2O
kXRYvQ1CteF0esCX3UweSLQCPvl32yhqfXXk3ZSTyu8buSPU1mZdVjMkAAHCmq/G
Ho2yn6kaQ70MgKJ25JzsBMUFRCmiq92w1nN27lGif82ejjWOwEg8+cj2wdQ0iVgA
VaGm7+YVTcpnuxYYy4zdPa6KgZBMG5Uhr2bGftqMlES7twUrUsY//vUGSaEScqwV
ZyDC0aHLyIrLBKQ3a5wEK4mi9HCTkSb/ForY+Y6d/VcE5qDEIv2E5twkvb1+0T8D
7Hf/+F0VdbdqDr3WHT6Shwj/jDKE2sBwxM+Rs8yozBBPhFCsulXCpZSRy1vLsuG3
s8EOmlxuEm/Gy98lBSN5Xcv6qh7Dw8xXrK8u/h66Uv+zmDupliCquo3xit9nqoHj
VDXur0fhN1x4WmltIGpWumOLuvJuR7NTnKL+OoDxnHsg5f6chGU6Iwrq12RRLf56
lTPVRAChAxA7axBo019/yXF+YLU85q58kiDqpjXSAbVGB+3v9Ge8Zktbk/0RSf63
lYO9U2XYCbc2uAv2Ow6wF+T47BtviBoevURJtFdiOB1zQrTBu5kZwaDIqf6dQdLo
Qlp0aXHwhD0bnqAn8JUWho+OMtYz73czyM8xP7d2CEE8mUo2qDbN9qTJxrLtUyqm
+CcBH+e7O8E99hoHs3g0Y69FxvGmjHNvt88qCQgaigq7Zz+AZP9+5v+yQyL8+YYS
iVLKQmOZhnVXw7ymFk4GgJJbSVv3mDTyyyUVbIerMcXu7rH9XJEdbJEDZWA9caTU
mJEriScWUqGKyP0yr+rymOgOEYOiN6jp7A9HsXwaM8DAHYxp736zY8Il4ZcuM9n+
+ZAr1fky3OeeWsyHuPykrn9aYUSOF9EP4wrmGPFzLTmav4fWlI+UtLUOxbhksTcs
8e57dspAk1ImQuHkzuabRWaUWqyntwoCxiJ4pUkOkOyIY0cg06c7liwx/Kna64Us
dYgC0WpVEGar/15rB09wWnMC7zxEdyFeBBX/I1PIouzr3Fvo1rEMKX8yb23sFQIp
tBVr+t3NpJ0t5n7aFv0J0pKt58WNCY5kM/N/8Yo1TRZ0ysTs4B+qFk4GMP436dul
DF0cczUOTvoWXMuKej96XZUWzejEx5JqP4SvUJR2cLyZk4hER7bGgWOwATez5jC8
sC2KTTzP2SejL1YjWJfZ7Gt6rdFOGCZjBixLIdpKuOA1oozReaHZQIoCVC4ER8dM
5dE7Ieqa0o2442+u8Ssfej65Qmhsvoxr6lokihpF6tACCQlEnTLUReHkrRid9d9m
WhamfzIkxNzDQNE+eeHY3EqVqROXbcmSNHYJl83SC8R43rqdacJV+De2XBMqrzSn
OElbGjwqqljMQ3C1epIm7vshQAhLyTiB9Wnl7K6OJnq68LHQnxUpOl2aqAVPLNu6
f4ChLFXApmgxveai+wsqlj8VaBZWT84baj5HILVLWtkHE49gLfsHsmVFFnXlsnOM
HQX5E73U1zJRELUlfR9p4t7iyX6CcdOl+98bhwNFDbz/gRm7oftwwA4ML3xR5PwH
XAZ6c5NDeXlDytI+7A+X5OhegqwpfO9IDpYA/8i5gw9oi9X1NOHr9oeQTXEhPLyj
uhetkAColX0YVe8Rn2lf8nVTzvMBuyPn35udU4HTUX2fY+mqclIzx7hku24Ci8zw
Onj3ZLrXTC63qDvSLfQNpPhzgRUk2cbfnF97rPs6IfFsjYOPMQxxLTh197EKM/Q9
A5QdFUPFIkpCwFFiwUWE1bXyuj7ZXChsb6fzMR5fkdmBRt+NE8wC4oPftaYH9Z5S
79fILmP7vJ0Qgjx0T/Yu7FbaXDf+pBDEg6WuCjzwoE0ABbpSL9QvFDWn8rmBmcot
pgLQ9oTMXErpbTRM4/MF22kFlDUX3VYLAlSNQmjd1nc5TnsSN5LoWTIPeAgejcY2
yFppJhwBkYPQp6ykZR7h9eNeXuFfLaaM3J0dQxXoLze/YNa7DmsKIAu0q3pdtzmS
1zhwYMEOZ+6qoakQEgbZx3c+LBurLG72cITzgXD4IFEAxJq991G9QV7H821s/P7k
Xf2/xsjU5FqrYVBAdBtzjPY5HfLNxszp87WKTCtEGxE233bD3+mZ7z9hPaRadvvl
LcIU++htqjK7mt8zgtAqpPgtDD/5r5NfVB0G5qT57535uvdc2Nm6QQ7QLullFwoz
5hHw1/tXC+qSek4t4SJqKG6gO5SwMSy73Q6qEhZSG2ZFkK4H91dcGhpkNUZj4Trc
tbSF8VgRlSbkSZXNkxw2kU9AaZu+R3X0PEfkH68Dzor57mo7sUz6Zfhbw4R/D/32
I+3W00juLGaKfh7HWj2y0MTDPfVpSyS0JYS/2K8dDqKUzCQ10t7vXu2TljwEJDct
oXN1A09jQbcay44S3lVfDm3SDEo/7pZq6+JqeuQz0eYS018yiXbWIN5QI9v1Nwsi
w92AVNGgR+Jggd5AeQW/4IRr7ND7oHEum55WkWTBDSXYqVJhfFqaDCI9EXvrk/7p
APqIP/DVOC5kx7QPTwinfzuftcOz74ddR0qnAktKA0QoQYYnr8OuoY+BXdhSY9zw
1QExH56xsPob3r9Xh2LXsBGPmNGDl14HYr30UlSCfM1HMpWWil6UF6Mpb94zf2l3
1jfW3IzZVMW+1kkpiYOH+Ccvbgyu8LOv8G8uj8K+yxT2lwacUp/5S6JZI44+Zqyn
BXg3qCf9vBL/PAECt00nAQF0JtRhcgf6Bw4Gp8W8+kR1XTsPaCyWyYkmJujgwwj0
2JkOtThCEAY93CTz9VyN0zgv827np+tYUx+ZYZhl+vTdJQl/XgTx7QSjtEP7LVpF
TQoOg75pWckte+w+5Gp8OsCDNFTgPpkids8noWxAIKtnubaKqG/OtGiZJOlba7FQ
oACZ2oWhqdTYqFdQBu9uhSeWO/+pSVRwI13Ry/PF03PHz0cY1jhJe6MT+9txK9Z+
Hq5vresIFzGMjEDQ/uS+pLh0UAvMORJbVM9VPFNp/qzao9ZPXnE4CfUIjfiXNec+
JOLbNPthymJOIX2CTolNkPXsyUim2YFkBjhzJfS3VLjoBtabEahAqmkFNZMIpoPI
WblwJE5LpH+0tMepTH2wF/sZ3ukXwGkLuBRhWSqbasiU6s3Pm9OV72YUrwUBZD+8
so1Sk4BzDvw56cP20IOfekPAh5atku454P3D3GIdfgcv53wcPfExEWA4K2K259Ce
PGPeWvHO1rtFdN7JSYibd9Z6rI6btMcrJ6340GoL0AzRQYJKg+4KQVn/rOpFIi+E
cxSrYjpuwxYa+Fd7GKXdWRzly5BELzusa/LAdN+xOQxCa8T+J/9I6JT6iT+eyBCf
cfU03vKwTnH9pWatHugwVIwzqQmKjlbEn6n/fg5w3N7JbxUskcA6pTXhuGI3NaB6
M3ySAflDpH7+fGZwjpTOSzGklwdR7Jhvs3Ec2nFdk9SfeB60amNkDfgS1zROEB6p
5N9lMpZ1fT8CehEqP2BL6RWQubGnO7UxGly7iicW1GE759gwYqVy4A0/ZlBopoj4
6PwpQs5xrVpaus90rEEXXNsv/S+Ec9jhTsbWAH5j/oqcBQT+vTVtCo1moIZTa6PT
o9I7i0kodieJnA8cGKipJjjnu191G8DrQ++L4eCT9DUoAgE/KlJEIpbOyu1rSTlv
V2H4h+x6jwvyHMBb7pVHDupkR/SJOIsyLzETm7DWkjw+Q/q5MjHl/MPNj1e65CRS
5jCUDxGJqorCBZhJSYbXToBQ85xp+ZKQkPwq8lroUgVEIjKFyvoVaGihTdFfLJmw
nrVaqsqrwDC/36IrIcgiB6PcrdoxZOSfMwlktjgIgSQzSurOmDw5OV/PusvTwBps
tD8//Sjxh3h8LAPuxNUt0x//bYeTqjW/Kp6ZHB2x5XRw6QyTiX2hPwxuHGipun0J
KZiGRqK/awpqq72oGhiWywELBovyJa0E0uIjK2+ekc7do+/bs1iGuYH/gF6Z8wP7
T+l48VQt9WyQNUm18E+6elz6wlRf9Nepp89f+MxSOr3iV0StW4aHZhKaTIkWJjYf
gKySLAgfnttFFYBSCjMXCkU9hMUnjew3/pyWpyNm15IdPHlj91tAmgDWzk39Uk6+
GvNM8Wr46wt8UrWXcBwhgIsGLfr7A5YHzb3PubujydYgLx4nqxojB7NAdtI/TiRH
AcJZFnaPioN54z7b09PLB8Ofn1d3KsvkvSj7hJJn3Lg1tfUv31IvcyQdbG8ZPm4C
EAGiFwpbec1j7qEUF1m1ldaISt8VBw7eHTTnSgRoRFwybq4Zi7/CWQB3bHZ9BGAC
ENgfHS22jT3r0aMQ5pJMzo5+56pTZyKrWKdbSdi0s5FCW6x52jIsrZljzj2ioiUx
I9Dj1U+V62DMNUsaOJpSBJbFzgpOD5Yr9opaCf1JLFIgOxFLae8ifEO/V5gpoIm3
3c90a41nx3XBoEMLv5qAtymXgglJ8iQ1m66hcATijBis/qb9kDaQLAAffAF1hqpm
j6b7j+SwnFbKSgRBHfoCEME1YdcBCPU0I7wdLIRUsU3mipgX3yV3g+uz12XZTqjz
tdtkVmmyVbtb4FtPbrggcSPvovKZ3VfvWqoBF5c0OqCPRbGTe1vXQzDb+ZDp9Vmf
oDnhEusUj4tFhbzHzd6yPnjxjzlcKMu/VHrL6d8STa5R4wKD5L0e2x1DYX9VSdCw
Y/oGRKpVtjzwRPZuf1EqACYdyBw1X6SMNL3eZV2lzFxUgqrXd3K/4eWCBv6k5B6v
nEudm3y+ATiyzDwGMEGhb522A/GOQcsbFSv6TrhghGrXZcwDYWMkEnXXuw95H4WB
vLIXoL6qXcRcMv1/jDxv5g==

`pragma protect end_protected
