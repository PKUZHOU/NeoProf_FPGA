// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
zYkj0R93kpM8mFG57xWGLRCYTfCkJlwHAnmmq8YqtfKBMmzEe7rup4vZ8OOn
mUkeSriIxAmWs8spsn8n5Thnb5UV2Or2z6x8+jz/EmmFg00HEjFDTDXk2sL1
gQKbYkCDMCjp5yAGNRSWYC8eyTgGmQr7XAu+CRXZX28FP07yonaAhGifmKNZ
fvk9qSiWfw4IGAj+kT8d5rA/XI3at0infMPHWtXwe3qHrBxN+XsLCljFj00L
dvLC/sXx3OEnvFuCby/ueVe7+lBWi2jsxKM0LauENA7gG+imBGNaYmY3qwIQ
1Az2o4s8wVz6aRUPSWgUbJhgxd/LT76Pd/SilHkEVg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FN7A2Wgv8lDsi/2oGIwLcN5KeYW4epVeyJZIJ38KSlnONdBtPB8grraBwbZo
SR8sL+wv99E+5/XgSV4c2QofK180vjarSmM+8RDx85RoOxlfkspz2xepO9CB
WhIPQtuydDXMTfTHALw4N3KqqmClopu8/jJEAUXQx4+G2cTaCip7dj63GGKg
v6YixoC+WY7mDB/CXnjm7SsB3bqWm8wOZZRY8Fb9fdgXwwlopdX6XbopwA1G
7SgKCmPtPWzxdhTzKMzyts0xEG29rFhq+VDZRIqZ2rK9Asj+qFgcVfHjyq7s
j6cPPNupwWVnKrfC2Pp+xhfocEIOm2cfu5B+d8PttA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S+l5iSpvn5fXe4NDx4ioOhbrGPBPw9fkbf+uYK3mhdOISVca+34nf/eloMxc
2TI54L2qgMRD7Z4TsrU35ed/MX8hsC71Y3PfDniW86/B7YOzCaTnd/zsJ3lh
DejaA6ykQqF9MqfKwHjnfex/vgup7ncTJr/WyGzCwdzNb1n21prKn7vJKuk3
vHR1NWX1kA/twcruktfweuXXnDJYlM6QbnxeZ89HJsmbbt3r0RhLrqi9776b
UD5o02riW2HbGdpOCsn8iHIDAvHvgMmbJoNvFO7UuqvCIId94odWLthcwPQL
T8M3CUSPfj33lQtCRQpOt4e+dj1lCYsxaZ4JhY+jkA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RiwpuWg2zkNnch0om2gXCBZ1Z/Md4N+wzEpuQ+WeZ6bvr/XUU/8/B6nfTb+s
+CFahymm5MFxgtBd541YcpwhKwJxu/yc9jz5EdFp40apXkcfXGTz+O0nOcHU
LBx8XZEueOlv0pvb80B65KHd4rKd+FWMtooUC+/6/skEsLdYlyY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
wCuoRPKMwC6hWfH2PWHVWVizCYxwKeIG2HP/hiwSXIG5YKbROpVg7A0L9jun
Dr+rlGvO6gQgo+KGKPaB7qtj7ANapqWTZO+pwPPInaOZdIxU4iVUcnsvEHor
cZ2XIyIHUXfRL17wU79pjqBnofjNZ1X+k6m9hpNpd2fxjAqJVR5bOeMvMrWn
pL7i92kO7mPPC9+YwHpRIGLDaqhD90od+1jXVmnWnvLJPzEbu5TGU0ZjvH72
pW7NrGql69GnJRL/XQYJu2WByGW6LFwP9GdIy5wL6XmVDKthBUY+5ygkRQD0
LmO+h5y0Efs9HIdBuZDWRpS9uWU0x6TfFK3GZdfRklt9O0mpqfTvQGelJA0Y
cRpPztjEm8VDdGK0b0IYQF30FnsobYmyNmpvPjHH1AYKjLbtGKXKKkM9gKz1
7IkIUhLmQfwV31PUGzKbMUqY+0iVtK1wT98neDEvpmggg/Hum/NU9yXxGYsv
Q7QsZcwvAVIqkdm3kdEP8L4Aj+kuPH2Q


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Uz2uhG07Dr7VnCoQWl1Y2YdautPfskB4V6ZqNBQzAh0Mr6SAQc6Zwgrh+s73
W2Te/i7DRFBPgxobXxwrv2eNXxViNa8+lLsyVgHPqMA7dXbsWybsPwvWkxvE
ZVlXwPy8t5dwBdBRcn8XdnAB0G6eHsLyAqRJVEcJs59YrP87Hig=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ab8uKN4ckghDXYpd1JjbY01oDOP5n1JLvEge+K3hqd9w2Zos1YFxq/LORM5O
r3UTQrYw4lZPx0sV+ob4k4kmBrXsOt3E4skSjbrXaEYu/PPkMQShMb5QHdsL
hMNI+cxMM/J0xKdAEXsIjtZytq8zG8/wfL5lXVAEPPj2F/FpVvA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12272)
`pragma protect data_block
ecC5lB0IMrKKju60ck3CnzywmxckMOkgZtkcRgpdKTKPCUTn3UrBGsSmlp06
f1zUJ6whPoN2XObDS/ZAOCyGfxHsrwlxk549c8SkgeZm+NAG7N4FGQoToM8g
dWJ0VvNYS9CEnY/35rfc4WZaiMW8Hhwt6Yhupi7stuku2BQetQ/qtoWLVqPF
JJqYBbG6mB4+SgXFTLC9ahBInfpCGrFx1ndAJgR2ay1kvRsDvmOZNGGuZY2M
bzwKUwzsIAH5FuYAbV/FsvAUmqYULoMGGpjGOIPer7h0mUMeS6z3jZPDjcib
d7BNWN8acGA0hUMMWre6CKR5MDZuOBh/ZEGE+YZ9q97qax67fNCyVic6rz6v
Cr1YZEmqnJqtvgYmn7EwDV2PoEHc2u5nCyrRPtfjaJPzhStdZOLN/fx20GUJ
WTzXymn9faWnA9gz7RZGcZ5uAEa2xF2aC6AGKHtaX3Nfxcjt3sYt2pPQuc0G
6r8XhuF6+oj+vyMD305YIz+p8qwbMQL77NusgdUCUD7WYuwTW+xBlhSfbDYx
NOTkhkBDGZNj5kB3rRfNx4XnQJCYs2d5aMEXm7m4AfJRtjJHZ7UH+htYApvi
XVgLAiGk+jAWzxyx+CUjgWjKLE6kTe1DXu8Z3pzkChXGETDJ/0EMD6O2edw5
sxAI9UvoguS/DY8Ig2iBFvKCFXgRmY2MwCSsAz18vkGylCHJpQesTbvyba0O
XZtKb/nwIOsaAfVqXNXN/M/ulfg1p8vx3Wr4bunTsSekkHrv0khAnEnJdyun
3oeviQs/JfLxnUzXjWodKKq8IEbkBW8x0//aLh2q7gC91xHSGJfEh09yFzlv
4gzv1r4+rc/Y1VDg63YC76v8WCc08Xis9EhZCq+up33hqZaw/nTPb34b1lHG
y6Gj2micZu9y9vmXew1cNTlVS9NtP9QZ8NeRNcW4oTk0ozrYBOBrrIw0qa7a
NLZrjHBvA5MJN4nF1BjNduW/kF+LFDjFlE9iBAcfk81CpGpP0TbjeYOHdTxs
3//DD6pJOiLqSNE5sqM7jTiErfpiU2/ELG0OsO8o7gaDP6yU99ATx18jYT1Y
aaKkT9uuYM2uM5MrlAmAzXFuLfMpA9B5v7qsP4iuBw1PbGq+y9/oSa60y1NB
EuR9y7pI1uDFPRwyM234FGQrp38ODs5vzcNUbbc3ELs81KMJL7pt11YnGRev
8GWwWADt63xR84uNKCNZ1jL8gXL4/JOrE8lW7XdzFb1dlcFdn7hRTwY6noh2
FlKeSwjEN0kt/KycVnD0uQZV+GRcatfXyTarGlwPIoyRNJbddpRvqRtXF9br
4BnzBKz25BSd4t+UizaDM4XG33M5+tYH+FhcH1y6vkIjgAOB7qlRZqKLWH+w
M5EOqsjuao9f9NV7cizd1nf2IISc4ZMFz9TeK7TFlQd9mXGYk0X/fpDhHDH4
b7LI78KCqfsi4XZCuYHU8B7dtPGQHILyoyxKz+h42YBrneoGCa77HY2nqkCW
eeFVmMBqcMGhqtmJYMxAk9YWkGKb5KOESsvnx8oEgh8IgKdWfAeBmVVMKqXU
xySwdLM8fblG6uWgZVyck/Db46cVy0S6TwHFjN4goph/5XACVuuIXyVcC4B3
wQilKJflxl8Tv1zB5MOkfcAp3bWqQI/uzPPMsUGNF02w+BUzvB3h4u6F2ZuQ
R35uN4cHGX5l8WLIvAWH6uviDB5sxFYepf+bGiIFK1LVus6cfwgzXC5vcHLm
FcbKeggGuNHmfbCUXyVOu75HdEXUwQxXpiLvhILMiOmcr9ykUhMZHxLddxTA
/CM202Re1EpK9FGo3BRfuoiAGr0BYXq/WHzVVymoacs92oUSLaGmXJoECL/V
vd/6MtCt7potoiSmwO6M6MqW8FU7bDSjz+ls7Bwlc+tbm0FqdTuYtMU1jHrk
FZ5Mez1TVgEoD8tSr0jZjEbSj2ocZJx5qiyikRBYmYAdFFN/0LB7sY5p8oHM
eG3DkrBRWsIW/e0T4puRNq4aqG2uKkB+OV3Xv48ikHBZRaJi8+bgxhEdM4wG
p6epvZ0JAP/Dfj92hy88f14eYWq0k9QNGTQ2/ciTA8l12du6ol87gwKvm10s
LAC7JXgxLx3VdBlXDNTGbhCJMjqRFq6XJDdgKwH4lYksBvbdzFg+4pTQLy6B
tmnGEwYmr8M3cOaKhHdbayFm/mEuJl/09McsGRmRoDePEuom4S9JDnwAtxXa
zeTthaw69H98HBVl9FBr+AeFGDAx0xX/+9HzxZNo+SjVPNeWG52wBI6OlKF4
20VtddZdc4K+8mHHHLiIK111qdDjJc4r2d/2QPNKkjkoxz5WAeHoXdpmcIjs
fSH6JBzA+M+kVXUQdiRNtemXjBKrB2fMYDeyd3nPT/20LEZVleEmUZMDzKKD
+isfXkpe4LZepTlGxIoR37m/2o8ayNF1egi1PHMvpzbT6RFvHQUhGJp27U2K
BXoWD9+JInURwNfOzS9JY7wpph1p24QB0wqYdjeiq89Idgzsub/cVcREcV1g
7Ysczb2+yKA3u9X2UgJJzl+IyAu+U7WamWeavHTP0ZCZbHYrigKTiZtnLwNK
/HAD85fv2h67VtzwYv2FVW5HCCWpiH+vHWJOaG4jGuPY4lKyJtzNoyInYwOJ
L05knBrm3B/vp5PlmqYojFvP7q69SMXUZISqqJrZ8RdyXpNa8dATOgH1TvLs
hlR7yW78R/Gvqw3csu6ReziAvomNTkeuoOmpajoHfx3M2pxn02SvMQKr+qvv
rHV9L0B67j/po9wYn4HvmXByINciUyE53p9/WNITEucrb0TRZqh4HyCjlcnG
3XUOVy2UNn5dqXOG/SKYH/caUd9MtP4iqlM/cp+fC4RbfCoCfGdencH7p1+z
cvzRrEn2nKZ27gx/7TNuXMy/jBjzX+ynWq2udffL+y+VkHXhivdXbPO7e+fv
cG9GIrQROyu3LHsH1o3dBHGmt2mG/XQPBTsb3m3p7cnJgKA4jJ/OwMasm1zX
guGQfSysfJQL8Y3qtMYLNXtQoWHNG3RpdVhmQD9IcmFe2/O/Y0bibV9sFFrU
8CVluwoBzBt2qwXpXhoP3fSt2pbzCFl06bDlm4toT8W/3EywVyPD+pGcyM9X
S5rtwT7qBJY5/Dg+A7WCJC2AyEzPFfVE7Ii8VpOSaoM2PI6COdiOmuzMtbnG
yFh21l9J+2GyYyGHgXc9VwK3DijqdbQO7oZEvGE/49P6rF0nMEvm1XpOIonw
9t+5PJPPmX/uXZXvNg9bdcDhRqQhYoWWZ+9KTITdJnFTloJnQyRRgPJ7R/A2
ZxHp/JFnruopqXyYxjoYTou3N0f0u+qUwol/AM2QksXXWlr2DhUpuCUPXpLM
m5vBc134Ley2KlUpmIN6N1mp9W6ruR6J811a65zi8vfMvMvW90g23lhqkis9
0zk16uhT6vQPtChbeKkRxPg5CKf1szNUvUU/WxKvaDsFwo5BbDLUbewA560I
CXRgxrAFiTOb4sRa+8CxJrGCPfa8ZiUuDeEJefQawJY2jpPxolBy+UmkQHf4
QtMbJD8QE9ExzYgF3o6T4rgV6+8qhuw0R6yyrVkDVWXoPSdxSUdyzgVwG4ZM
3Z1YczEhH6SFh6Wnm9cwTlaP84evYJdFZB7vZI/HgMvMoWYohLL7/v5Hbq5p
TpqwEHHtZncyxBi+deioeDxhnNkoAn0kY74zhfbnjyZyP1ELmSphDJDGe1oR
wz4/1BbsxXSe07iNYSlkeqqkzv2Hp9x/TZPWJhVKebdhWw+DxEIqExNpm4mS
Sj42QdnoZ4YsVZK966OPSEvFWBozd/NDbW3Cxv5X5yfe7yHXTTGqPqKqSL9g
3XMN1dbuOxbRjaZT0UFb49DispxlsOjuCHuuIeugDmC6bnWC4s2Hl4MQ5QTd
b72xWnb1A/TWjs9vkLlwQcaYDwpMCnNDIdDO+cnx4HSdVEeydzjAkzS4RMvC
o6+TcotbndXeKBKv2qs/6EGN045UvG2yJcALodB5hmvgWRv51ymHJ6k/pHJL
N4ETkF+xXXlGD+eCIXzt/NKyiUmy/jZm/pe9P84mST3YWIWy8/zdw2cqROoR
cRX3Don3MTwdADyhBt29p+5zlkBIsLNBMBvK3qQ+5wtEo9rqth+Aui5OJLxf
JE40mKzYtsbDZtozfYHe/gZleOWivLbKc/hclL43iFwufC2SFLHOhNp0kT//
MauXfoY801v3mKwQnfGjXhNX6twbYN2JilmwEiEec1V1kY7daVg8O1dI5TxD
QrnYcMAYoZ3h18cB1kJy5+e7UB1VUj8BOCgIwZ8Gp+9OxIFSbQJq0urzb1id
dJKg4Fefrp2ofxROASmkDqin+LBx0853BvoYTh0Nk7kf8NW26dCSy2ItWGbP
K3jG3gS1HA1PeQZINfxQEhCcXSZdZPjRG3k+lOsZbx9bMN3nwURNQibntZSh
TubZzzdUFv3Cb2skR8Y9maEY9N9jsRR/InZ8sqYM9RXGaS4WQvo4Jd3jmDq3
Jctmf70P281mPjhX3Bcm4mW9yhqYdIeTRWeuJQQBpOyQYkMCU17K7LcXX70i
ABgmoAOJe51VLJb5WXBm7Hhb/fhCR2i5hp0M5fqzPouXR7JCNm9HCklMZnfb
BoGy+90PfMBBrzdDCsCO1651J5VznhQXAnIyci/3m5gsWw2Y3NnXxTxLN7x5
N4xZ5uRj1RalmMt1BPwvhh7Bz8OY20YlXPJIDPVyEiu6euiqrhIv/1X14v+I
pjZlKzWVGJH0feaUw2jWzN2sFVh1Ua+r5y1t+lavHqAwImOP5AjDT81yUA57
LUAxw1P260YrS0vUR48pXh0ags1CthHhzdZynA84eA+SOsd70FwW2D0sXhl+
+x28dtWCo4h27xwWvjs2N7fhUoOQmX6POmXsS0rWoCf6EvKJCukSZo0IhWGn
eQ7ZlG5yGGa2JFq4vMm+Opw3fJL5evkuh4Ghyk9t4TIAZcGM2H/y5e3G92Ls
DQFsXa4lSXBihW6gO/3z3Zim6lJckikc44BzUoiWDvI08NJMxBOe2r6wRAvS
jk0ScGJPQ76P7YvY4CaODLgUnjCM8R5TylUs1Q8Mz/B3goW76323UYLWjM1M
UfSAHVUJ6P3Od1jKeUYrUYFxWXecumDdmIoaNa690G4339yth3U+UaZA/OAb
iU3MDMIJV4PR0EAZmGujSGksn2ZWsC2JjsQ2xWfB9h0YuS51w+vAOybEQvHF
jPAf28t2XVO/rRrOpWsNCicXJoirwx+RHjMqfXnulqF29eqP5qrltrksnUOB
PzXarQ17Zb2bikMoAJ1Fq1++trm/u+69V/rgrg2guMxG5Jz4tJMRjhsTfFfO
jP1p0/wm6tqZKcIa2yohGcH2j1Q2ZYbNbtcatMgWm3mJzthk6g/9ZH1TYN3I
b5sSoE5pY+bp4AL83e+yNuiccv4LnA9ofXeSj1L2WCOTA1yuqQeI5tQHOtQL
qiUDbrLFqcMEKAUObglCZZ4PrkMizjbxgRiGTKPFp76TmPH6ozu7fpsXcEDZ
WztwEhowCEhdvUtaF+v/Qj09xFD9vyu2v0ug4GoPcEZNTRRP5jHkHAbIQX+l
e6DU1u7F91X2Mm66So2P1Kl8X0sjje2PmknGHOLRVKK3r9dA7qAm7hoYLLnL
XL/L2Rtw1MT7MNi6VHfj7id3kc0n15qC5w1fD0dUFMIZvnP8gcnYbmcvnjvM
C4Fvh5HPNkd9quMQiOgAofVEfe6L05eeh4jMuywvVJN3BtU5umhhJcV/fw7d
dGMMeL+1VJub28aaPA/r1aecy+94cQ8y1kpR2C6zrERoC64YfT3kZNE/CF+u
/VAR98ZAM/8jhcaRajOuHKxL5hG32XWerPFa1C67ayasra14601+fTRpt0rA
VPnIkNLNtNw39yo3h4OGqaEJebYLMU0gaNh4yucxLqf7eG+PKUKo79LNE+ft
pEXzWfQx6ViWV8G/ufRcPTgkNGTVAmkIs0zsLFb4cUS/RBf/uuyo0DNWbbRz
aWxmNyYNKuzcUUxNxVb4JyZzFtnEogPHLzTsfX0lVawUilsy+vkCdkh8qKu4
/zvijMyLCP9fahd5FNGloqHGpEWcnanVJ+SRK7CSezyOwgAw+xPGThRRQGFO
Abh53IGGGZekuDGaCXH09McWSJw/8xbdqCR1umHSJEUye6XfaiZWUpav2pqu
SbkawRY4zrOCtvxUdRLWEwk/bYLA+ND2zSGIQPZG8Mu/EinC/y0PyzRCbstw
1NDd929i4OMc0QWLOY9UuZ+fedtea9Hw2PjzeYqU9I1Y7GVN8gez32JX27q9
31esNo64n55eNPOaOq+9weeYilJhL9rnM4qfiYaPrEwRCsspezkU9nRtnWcF
NeEz/DBQiI9smboqxDXcPCcycU1HNJ73wy42FUnU2mbmfa9Wx9WtoFYeNhHi
m4/9wceoI9KFt3m/zrjgU3ydk0fW+EIU56ZqBUhmRTWWHNAQsXAaq3ObJ0WM
UBSa73X2xKjPCF+aYPaJN69yvXQkzTod4os77N9gPrKW44VETImk2FSQvdE1
mRuAdbkfRTioThxo4geTbmjTiC+dCiGEgPh8u5YkqMYI5PecaMXe86IUvOsl
te8xFZgaLms7ReiCDy0Z9erzbWWG1SNtewTt+dYFg+S+26VBj90MVNWW1qV7
dw+t2V192JGc7PxOav/zS+y0Opi6oklb2R6qLrYSPwNb0HUfywCbeOK1jn69
brsVUQPuxX78VY2ol2vPt9K2IqgGoyvLWQ1J6XaKYYSZvzhlpxUXHLRqzjfq
OwzSCED2217XHTIKamJ4I4wIzAHKstfkgGSypEXM28CKMSaS7bvMBJRIyyxB
5Oqp/lFYLDhmz/5vHzb9vBKT4PRwYuUrsz30M22P/LMuBpxYeSMGR2F3WWTt
EwYz3NePNBXV+C2+GcCCF3an+C0Apg2gq4irPWjdQPOKkYE6yzKUYyRMPaCI
eKwk+Ufz6ylY+5ifSLSYPfnFdNvhsf00D/QMJh8Cs/8QIb14Dn0IUkrjOykb
7mPx/UdfP/sAvfwYujMBcVVpc8cdRcOGKqV5qiIF6gcR5o2LYiIpgjtIaJZG
of1liCZUIaZsnPV5iRwCu8+m6H5GLzIpBkecTvjvccIcdFZ+P/qMD+yBEcvN
8p2VwN4DFTwtISDDRD3S/fU4L1cips/8Hos9JJoe9XDeOXR5BV7khdQ3fats
jk98I/iKZpehcGC2YlMeSKSS+51mkLkoN+WEjxM5X10zO8ttleU/ofYMwRw5
SUy/hK77XrS6AIR5IS8fqpj8LDkHYSKPd6/wZQMK/r34jiEiyCbHQkUUegqu
pw99GLyp0M6QLb377gEMfOl9KfPZAZjWGJw3R3vDmU4eKQyaabMbMWQUacNP
mEI708dBa7nbd5sGnmvAJp61hrJsIkV4YzKR2DF5140BpCFj/4tA73+E912X
GN7BEHmh9SMMzfGSMkfexWNcZqyVL5XuVloxPZRziaAPovc5w1qD0SS/oONE
f6a8GqRiy0xUHrcrZuKaFjMAnbPQQlg4RHa1kRrzKbb5T57KYAxEmjfYIP5o
i1IFCriSpMsZNmKS01CAi0y2kuSSJMWY3ykM/tnPYFyRXD9rnb311m1tGO2V
kjxoYssyC5uk3oofG6nAYAIAXcXnXmVJ9hMyRJzyZpw3WXn2h9RVEyZN3YUl
HJ/Wz5aotrHtrY4mt2h0u/xZsLrlgxaobMlV2caG5VcZJKL4oIJzdIGdBYrr
i407XzgqK1IyTTsrIHP/AUCqISX7mXuUlm1zQPOVK5mzjpDjjQVmXmAlo+YN
ey9h2fui5nv8h2XcoLu93Dn43nN/0uK4Rj6LXWi7DMS6y0/sZqmMTopfxviZ
xGpSj1Qr5NS6vQHkMYRfi5XfDJPOg/Z9vyJi0yTv34bbgdaDcWsk/RBnTGHT
+INz55b/JlHwq/exjYa/kJUgG6NFsOh5O7sET11Fd3YFUH+1jrMa6imBkcdW
aS0Lr359gvRmGlqIte/ANBRrcgR2ynG0VTyS/IdN1QF4jMfFhD3HegqYw9Vf
wbxzkCBSj2NijN1kWJFlJm09kGJGDJdb5jEsO5EyIg2tUcBUiLa8c2LAFXxK
pnGDNrhJGapqNzkJ8Qv7JAxG1K5YVkDK0OTeypARMJ0gNVbaainM9dfhvnRz
WEWwQFlwPxZ+hD4ey2rqTp9ZdgNXMtgfIINk0GTFgFKKcsiUzKOaSGM7SDbU
1I20PCg0uR/nOjZBQiKJ2kiHvIkGyfRVFFIjspLvmOPNQ/0KY/A+7+NQx801
oXdXahuF5VkGxj9U1IrsEOeE1I4KiaC5Qs1Wx92HSZaMTzR5mZb10Q20TaCX
0p63x8Qhc/Gqy6gcdn19U46tJbGg7KGzlXFnVGWymp2FWVJMa4DKttGUmWCD
W7eqc7TnY8DSyvCROMNIhU8fgE/EeHTKelxiQGEtPr4LPGMKKhTVBveUxwl+
OvIXMcgUoSUSx4qBQRKKzHxxZXtbt2B6VFU/LXc3tmgmwpRVc0AXva6fd5/N
OuoufhUJsh3BD6DVXBbqiRGKoA9iG6g8f47L1n3syWvdDQF6rnZIGs1mBH4y
rKNAfF8wwbe28BFjPWCY2aeQfLVOaCO58CwiSO8O7ID0Hv4syNZ6DAlLwVJ7
k6YjKsDejZycRhEAw04uqbHZv5RL7pi0sQ3YjYBa0VvdxgjU6i0ysciF62SL
XfaYhYAh/KsAKpqYUD44jzjyRtP0nMXzqcjqUbhrgGyRr5+mdWJHDyDduk4U
/wrAlWLFaS9rpsttuU840ebnXQu2sUFGodLyrMd6KbVAWHcAQbMrj6NXDpkB
Ys3bxm/pTyIOJhxlLRzeEtTH36jvNrTnOPezvYGTZZPJJjnn6FRrxslNhaYu
7kDymJL1Z4G63k4Pq0BWIoNtrTqtvqwMe24+ki3JZSDuaKCNoxtuQhpamO7R
gUIDbu+PgnT9jQuD+INqRaAALO+QhpAuH4IkFQzqKXVYMycab+tbAvBJypDE
41jglkGdfnEjeY+TL/zTaIeTAH0pD/GfuQGInTTeGKAoIkFR7r2IBLF+PDzk
NZlS4NfOY5hIKp9tfcqxSlJLllGUR5PDFnxi0yCSqFBi3JHLe8TxuuVgHZos
Y0krRAY8Hxal/MUpbfn8Ob3/NDAQF2jFaMuXKnqbykgp52TQPy+3Pkjzzs06
dkzO0QOrDXFGys/WwIglJ5GIeuTQuF7tMqlrkcZUYAntbQDjI4UK+SJG8EUm
YFQVHXrwyZkYbGik9fVOJOPUueHY5rjmL/Mxi7Jy5WGFP0FZFNpa/F9Pl4Rg
1ZJg2EfVWc8PPK9vDEGzyZFOUfybSw4PI26TuEDBPycfVPybeiG0iG+o+Ctx
kgTc8dzlylDuM2gk4dheYRnGsmBum4NIP5VB9iYIqpPz7DBNX76qX8EdD8kl
orl47HHOuEokmKL48T112X1BQ7YdDG+FEA6K0ZXZY/5AIShD85Z+nZN7bVys
qV2v9cf2qA3QOJQSXGzHX5oquhXffLHOu5Q6tr+lvDUmv902YsdCP1JNUheQ
aPL8s2jz6s8KV0/D/iWHuSacIzWEZrmPSWtVf5PWlthNiNadhEr/Dyw5lnb6
JS25oH8ywgpka2ZGvy7VEly73yTz/ohxie+/oHEx71IA2Jr/ZxQewNKts+4j
PndnDXtB2GP0Fe2BwLzbZFNffEMyJII4LkRqVmCDFSyUoiTfWpLqfl2ilOm7
zlW1G1Oo8x5TwrWD+ql1XMdQYgNOMHIyryXXVcfwFGx2gqkN9zUTi2iXaNio
3j4z2ojIqSf7sXjNc5l9EWUGtikrgeLX1AxHRymA8lNO2r5DHXmIRdrqYswY
k11JqDkERkRSweV9Bz4hHGP6nu/hXbzix6vmQNNE5IwJEAzJGKmnwgk6vKCS
jj/ibyrkCkSNq8c1YkWCiIMANtqYUWi4lCl9FxqTBvCt4DWbrIso6W2sK6ru
JPK+5fZKMEd9PBcCHYK7nzBddrIqwKtNZXlg67fI9Oc7fk5+BLY0nsKTpyFc
u1mPxEkp0nQhB7m5fWyrenwPLaMqVLsbW1FQg7lTkYCbvmct9/h3m7M/4uJu
Yp4uWjcEw7U8QKN2RFnD47KnHPoysU9TUJ9rsCz+uy6W8R8cza8JkXT2e06w
ceI5TT+A9rctl/Su/oWtV7TlEZlKPlRcd0MViJ/XEUhmI73Wpf1xpuButWz8
61xKKI6ArE7uyRTT0e6r47XKDl9/za2yQUEs1ltklLbrdoLReUk0dbHvHhhm
+/EO0fyYJa3NkV/wtogfqPhALYhK/ApJAu+UY/rftrW1U9sk9eFKvJkoTlnu
QGV7Rbn5xBR4/wl89+DZLaX9qv/jjSSOoWLqBe20g2VXIEHPXsg/vsvgxnOZ
OS3i3akGbDuUf4DvqDQZvX0Vp96Fg/CIUgcBxwY89fBuf1eF4GGLeCJ7OwcQ
dbrEt83PL5BuME+tPXG3WdwqrfD66sFYglfjyexCs8qY6eq9Rx/THdp3mBHp
Lzrg65gsno/PNu9AExJg/xmq9KsRzj2PGeldZtmk7My0fQ1Ew1mvCBwFgZIR
8LgbbhXhxeewByyWE0g5KfLSBn93TQLPKpl/LUZL5LymVHGPjVnfuEs1R0KI
dB0QMBkkqSMj7Cl0N1toF9NPI9RZBG71+woNmUfIb5reCupAwFIE0a75NGzC
VZKSsXPh488kJf23oHN0onbV5dt1QyP1kTz+bpfmF1JN57/1M7qv9O7M8cJ0
d/zk83XSEi7vGEv0gIChkLT9CbYt6MgjW/w9M/FJZvwefw8BFYJARfTOkDrf
8OEo/yK/9B6RgVrrOCRKjrtxIgsN6FrU9TaXxWP5tbKsTnnKG2tXNemfEdx0
jGgD6QP/laipPFQ9vRwk2229Y51NDseAZREvjbj3YYrFjJSYOI0BCjRTnB7I
FD+ofVFJU9YnjM5eH2EBSyS/41aoveKWHbmhqWEZOEjH7paZhohpE5NdEDeY
J1wa9Z0FJylT5yGk6YXD90RLc9sW1+oNgBCl3UGKy38m55jrEyQlQF0/a5AZ
cgUjkEWsP4a7Z3kJ+q57rYzMl5Nhr3yPUC5jyBAefDIo0SJANMhg2ay6Ndmf
DBLNRNKsv9PgGvpPrtaKk2mxnpdtOC5K9atYxRFtHci0goKomk8A1fhWy1Mp
kDGQ5OOCIbQqwqJM4ass12aswENPKqZPyjB4YEqZe4nUZ2fXczbYV3Dfi7lm
+xIrJy0Qq8xZ82W75t073BLZHK15qf/61e47v9mQZfRvwxQWZsgRdmi/iAtV
fFqpveY/erodQI/sW2ERaCnEzKj6FYS3NX9ddjrzk27X7AULKSH0GfnpTgcW
F77KS+v/vzOn8EKK6pE03ga4iijvYcXQINhlN2720oQJVIwQRT8kSrguergY
EtVP7tUuMM1JFsUjkFduX3f3Kla2/apyCO0JGGMVKypF9BoOQraWFUGkz+1C
aa36tqrCUiHXuTYLHXBQPlyvHDq5GvjkEFcZbc4yLLSqyEfNdlaYdUvD06Jm
j9AUsgyTApoJZbc/OvCUqL783jbRu+EzcBt+9f5A23Z3GsqnYRAdyouLFUxd
RgLiCbjKC5Slloji5QNsllxNq9fzLJL9enJnYHstIcuxjwHuN2tcAZZEQjvw
bjasKjhyUv8wLC2tpb/8QIoNkMqPzuXcVTFeXARTyK2n9jvkYAHH1wtyiSe9
Fq+bjrc59ZRrxRz3uFdIndFSNueXcgCRMp6j9MXcWfIPJuKuiy6ZWIBsKwaa
BtzqiqRg8XmjJ1FLAERHvtqiTa1OERGPGFiHaA6A5WUr7JWUNoPbFlJkdqw0
sfVYu1dEe402ktMoxsTybow6pezrhGTCZtByGSA52DDGkdQWN+lEMBvP4Voq
N2TiSGBURgNOXIX4zm1dGox2804N1CGbJFimYbxdc0h+mu5YigANXIjMNzMm
VIXcJlVThOmwt7s/nFL2ujPnu/VirXng4GPvf5rMg2TyPLdiEqbCQqz63frK
8okpJRLfazMtJTV5DIvCCyWyapUliG7QRkP9yeBtxRbEaBSYom1cMpXF+FoS
R2oXQYbIcAOTsQE+9Vq8gEgR/IvcSuuGPnM+dRrvJUiWNooKo/wXfvy73LZ6
0JF6tBejVk1NZtcw7sWtN3wtvRQIapDbzNqvFiA+200DnDn1vM4nrn/z3JKd
qY13/AyUHw5TL76eGPvFz6RpzZgagwEqlhHdDuWVmN1zUxyk/3fMgHYqMzDi
EeOQ2bOlpU2cFOguNIy+39Nd0Lparg57TijRmvfknSF0G4DYu0SW5xhjHXHW
Bz7PAngj8ewvrnBSaC5ApiAL6TsJepUDorlhx9BPYTaT+JW4R/MnXyjBD0rs
vgJJuUnekjGR17PslePl8SR5KBCO9ePv8xhUDajBUu2qSG44387KpFGgxEuh
eY91BvAaJuUjVEurlyTNUNUzhczBBc0jT8FIoPxVa+WMNEC54IymFPCjl0mk
3yFhQDUhGIw8ohbef0fWXTF+pcZ4PY2acWCAYJq/Tefu6EcHpWksrLrTfPl9
IyAkAbBLfgFdtwT52ww4jSsCtgsdOVg9+lmGn8UTJz+dbICusBs63pUoqypu
FXAzgzg9lQ8nEowRy1mOT9evSIsdaEOUiC9MNWDMdQpF3vCFoHI4SVqMaJGh
r1UJZ2nYBeFlikEJzhsVbFTfX/IuJkMbPNUenxoYE4ZJcupu06zuBTRTdig3
SfLSptBA6645T8YCl+/pjpa03LI7YWrO5h1I/llaOc3+uOJHolPerUig32sc
+BhvvaQ2W3AQZxwHTw93wPcKQvEJdMAOSBXJ/X/V22SL6QIW9EPcf5FQKvcn
7hLDan7h/l7eAVSRFDdgLxKiozR9im92WAGUi+ZmVwedlQT0FxVzQfW4jQWq
EyDN1dnwRGinrmajotVml7pTQ4QjHw+zb4lS6hddgO/8kQbowfQWUSiiy+4b
f8/ykoKuKBRXzbPUmSSlz9sdigG4Jur05Is8bydr0R7q4nMt8tp0nJBLBM8P
WACZHWC2zlveobsJR/7tFrg6SYSuTdqFbeoCLUM+0V6cIZWeUcbzAx0JwHZG
DMkz91Q7FExWh3VlSxhd1hVy2k1cu6SeTXkwKcC3cGXJxwT4p2AznygkSxlp
nadXEXjydKFjVY3LT+SCCoUQLlCdg54/yEzQbIBoWR5lO8Xo1KHGSWfJRrcI
3b4K0nx8CBsa/jreJ1aMmFyVXPR1F1UsSVOOX6JMufUXTf/GIewHbK3FURZS
nLcSsej8D91aJJQHRYwnN/8ZAc4VCaybdfkymPI5/m54bX/sjvHC7ZK427fh
6PXl+WwMMPcJk0I2O0BgZd7pyUA8kyGImDK5vNrAF1KHVsWPG+tPJKD7t9a/
rTPcB09sMGYwMy9/ThOFFY0UC6R+HnDH4cmn/RkE5sLXUr4P4XyxTkAlbq7t
0ykvy3uqOuO4ft6zWtvy/M4kaj8GYTyaNkSYBaUOv6ifofSH56nRC+Gi+s+s
CvVzabb4wHOnM0Jk6iLcxafLOhkvEujQBYY2WyZSUh+ppoQKqZDs+9YOQziT
/+hnQlLw+dGQtCbXQ1DWgNMi5NOiI2d76QDe3URJmgL/a27oJKaKoZORCJu8
DipWSDnuxJrIBf5YfSp7cyHJOxE1cf5csm6E7Tf4WrR6PnQGoVA3/CobcjyY
QNAVKQPdYM79CfTvj5GDp7SMoS2o/oGpv747RS/VSaYW05L6N2hKwEre3+nt
8OtMgggGOY2MCpvRhDwgu8qnWp5AlnbJxZV2Wr5EgkGS0Od6wr9U2ENbG1xH
ZOw+fxM5fBHf9FpByOQ3TPIUxrIvOu0B8DxM1/nR7DGb1KPQSMZxBcbPNZ2P
d60tC0jWn+r2gy1WoMnts1lpSR+RsjPxPQbOBVwYcnSe2fvB0j+PLNX6McLm
NRdgixFWsaUdxerhOKgxruB+51BUEcoI5lrW/HiL5iIfBcDmenmRMdB243AJ
FwxGryThHtYrBAtmyYHZORzShDUacBDXQG7pcMu9PucUIGyOZ4x/WjO1IMSA
UbuMAqlmUKszt4j3KSwNJPYkZWGfmaoa2++dzMcQBYLRlt5genWcSbh2FERi
aHNzt4D/H/uFp8hsF/5VvdjHJzlgTxDSRUAArwe8f9FmdIYZCzg63N6nwA7J
rWTWHXRSt7pdHQ0Cs2DCazGlke5y4qP+9k49EJxSp/q1D8aN4UIKKrtPYiCC
HZ1auHbzBgCGxzX2KSBThhcoNQ7Mva+6rdX/SV4DOgO9z5VtgFv70Kara+pn
TJwLyrkgIWIYsus6rTi/0ZqVosSLZF0bNO0ygWLfDypmwOTEi9W40EuPvB5b
B5Fi82w4VKsTCjAKmYg1Rg4knPTt7GKfhK7ueukdsOxPQWXNpab/BfveJVNJ
nB0nZijbf5cF4iaWTh/QneGKIHR6buA4XmI/97YzeUh3ST6VWTLrBEhILF14
j5LdMV+7ToRpxQZq8LsmTxdEQJN73fyDfa14MHbRC1SsQiE54lyZaRnPP2p/
zIqvvWl6CO8uN2dpgr9LhMwgfpw4skDsqDPojFxG6zqjMcijrwmTGBrWzdCI
erRx8ukXRjxx1KH7WmeVdKqvsBJspr8ReNtxqnHVYMSY19QSzDFmRqU4dk1O
C3Otm6pO1d4ltO1mSqE1WthP7d7C7qdqcOwzxOzbuNoHe0c1hOoZMv33yfTE
qvoCSHQOirTh6lqvCNqvdmwrArN2o7pd8wPXdoBQrwi/qQaxFymB3u42iFMB
4+wyLpVJCFVv7mDwPc++zWfvAgLJUH9eLbKQ2pfUqBIcgg1IUEszLwKcu8Jl
3mrkNIQF4CycD+gGeIjmSUIWUHPVevIiaPogLk/j4Nvd5PmfhItl2EFTN2Mr
dX0HmpEEgJ+4mMRKJ9NQRgqm6fdY4EaweOok62bd3yjgHvNgGiWM6PxFI3ha
snbhEhxWo0G8YlHI4AO9fdtYIO2pV+LlUsQ+MjRBWvMxoviO6LFc1dYX7mS7
lIfa6aYEuHhr+6PBS3HK6xTlbbjysg+VKmlPlUgKVe2YtDiW6mdUlH/25Zd7
kfw5MQHKCgiTFS8WwXK1jMe0lCO1TH6bSh8uTE9rSWEIA5mJNTNQs7YLN+ts
CRMS6CZKwZSjM7bSZsn1irO1Bx8UwMM+r8O6UN5mMdZmKs6Pd1h/2mJI1/TL
VvAMQadTzCgzudX/4+qKM8pJqAwB6l3dNt6jqvpXRZ3E6Q3oofihZ+LRe5tY
kkfI0XDtTnK18xsvHAWWRhJdYJvcvI5hORd0+5fDn2BFdPs64Mi2pbedxWSV
9EguZR/OgLMTT0GK01FDuDUtgAGW47YHJAFLsoUB5UaRb4rRL0ke2w/3/New
/cdBMxPyRzBq/fuoVdAkt9zW4aQF8iXOF8Jq51ZxqLZVBQGlzWc2EpuloPf6
BooPGPaLcPCPUVIbss87mRoSuYOtNgbF5OUGbLsyUJfTfNCh/eUaZHd0ReK+
9Y190haonO28rCKNkFwyn3Ams7Xuq0QGyDVW5pDmg0xSA9QD5/DaEBu6qq5z
vGvj+lr3WXO6vCa3x9I+5d3MFU61x+e9XVopbOO4ViouzVyjSeqDNIQ8pxS5
rS7qJt/kMqUvGynyg1Qp1klqGmFVrFvxpfHGuaKAIk6dv/afPhIGoZrY3CFY
/TphsTqAlemCwawsGJzvXfQJB8tMZ/8btw97mEIcelee+5CEcnxzt6nHeFod
0NMdwnSvGIOmdkbAhzerWOM+bAWAn3zxuLO1LnGFIgeZgPSY4r+rZTGtOhwi
MAKZCc2KjkVpgcu4D1RgNZxZ6vt2mUxZ/0NO2g9V1rL9TeMYLVlngyqqrj/8
1Fmjy2N8mok/g3Ss42aDqFJzKVVxqlgUGzwvvDAYjqZoB0ctMxo1Q/v1cf+k
YyN0OEcWO7QR4vXN2foC0UYLBNELVqtA41CvDze7E8RP4vmwpjNI9EOVohgc
uLPtRZSriFOe9uNCsSdw/m/XKm2Eg+h8zRwPBq6S4eM+1Mhlj4QbZPwdYriL
idskhuFhCLOl0SNVTTNvW3FC9NpSln+AI26fegwLuRXH7NlC5dH1EnDRrxC1
aTHBi/WbXCrXROTnemh3LB1+CjkIrksh9pNFqVV7u9kSFmtpxjaptpOdOGNO
ncwfK91ckQSRpZvWi+WVTBUpr46TWIYidZVQESEw5V50aSlq6A1yEVbWM4tt
8hAaevvzqUTE792z1RoKYi2A+PVAv7ygKEm25R81nZtuQDFOGMUAzalVXJbb
6d9M09fMwI6eN/EntIq//vFkCAEh82elK1B9rN/fRNyn6TYsw0STvUDe5B7q
vQ5b4ClbC7hmesTqovy4gBI9WKoZIW1OlyaiXHFFLN8=

`pragma protect end_protected
