// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TsjWB+fBINaD5eWEYSZuiryrBayrsUnGoQOffms9IEv3uF/QWBU20vncwmL/
MnhEf7KE7Niv7VrQj9h+q1fkEXygcanqEj3g+jCsITvdF1trEzpb6eU+g9aj
xMO6pgttxkY8WgKvheDx+3gbic/Kpp9WrQS7sAvUmUxsJbkZBrXi6OEuVVpa
Akqu9kOvbIw9bLhutkUOgitcbPsqviyARPpYXsAmfahz1xGpGCd5iKVMtfpY
8E9a2q87nyKxRbl0Q8ZTychZTr0tRaVMyayAhXVx/NV/WSNMOKECz+/xbEFS
9TiKA1NraS67h3Rf3GCdNVhJ3b2IZnFChTC64wzSHA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mlrrO5VOiSJXHlDe7SqBxoaH1Q2J/jTOGgZAU/Y0o7iZjcq83pD9F6j1BD88
B9ANV042fYEb0PoHIuZ+kEf1A21BvKDLWqzFYe0a/VvEd2RxD8VIei+D36Eu
Hwix+UVDeq3+dm/9wXUP9McKwfTmvllxTp308Dn+8Tmt9lMlt1bCvCoXPrGy
cU2sTmkeZMDgEs0rcxLhJx/NMhN9ASS0Q0INfsZTgPz4w8Pe9w/os56hz+SP
Br8ZkldZvmQJ/jc7v/FfofXsbISDyVUqj35kfkrmgCiGMzdpP6B7S+JVPnXo
N0ZkZVlqgD1batYZ1qhvTHHW3iT4nzEhqbyD5H2MYg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XiQgCYUhZS/It7X4bn1cFAtdAE3GucPQAIiDHiIMVrzc6d4GojHdgZjywsI+
RBpKhVHjOy+Wj6hE7Hbrd4gy6mlzusmpnMjZiefpwXochNWwb+9StcFcoYWX
lj74iPOfMOSOR9EIW1QX5CW5VEPF4hHDivqFTfbD+VA2iSxiY+l+3V5IDXt3
PlY61meAatr5xTR/j8HhGLd8sNLCqjDf+iQ0USbHQGnjeOSwngww6r/Ob/Vk
aNz7lC5DN3LlJXR2lwULeEeqVmjwHGFVh/9uJ1QzPClDHXHQYI4nIPbHK0jW
SUlvorMg5CJSAUCef2K31oGQ2Cdjo0wR0kTOW0D5Kw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lDt+fR9yFHx2V/XEEx0OsVbedrsUsgI7DrDSO9EuCV/4/oniLTOcEc1d7Zks
S8xrhwmfl0NEAYuo24nMR/KJMiXqqDxApD1Nm3KVOk0OiUga0mihP5yBJl38
SYQWW2+RXxGRnT6g8MMrkuf0WQe6l07duzENlj+4MX1fVFl/NTw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VJAA/3lNjNqIFtyHSXFiMUdl4HIstNXfgPWSgc/zD5P+e6n4Itvp9f3Er4Lv
VkhIZuNEzvoBdhULIf0TT2dqp9otpvnW53tkIYFmGS1dzbeo/rjICF4QsHSZ
nxNZgKnn+KqcMqGbqRpYLDW7JP4VTP4hje4oGP71sld90EjwkSy2VzmuhKcb
wwcu8MJ1myuLA11Ip2S4q0/3NOaFtMjtpQ/k6fhAATWk+10tOkBbkr8jYpAa
uPHjrbuaFu6ZTFJnWdptr8RC1C4nvhN9ofREWpGj1KRt/Der0O1kW0uUhllw
1CYJM3zYmlOyu7i0dO1iCtwYZSVqkYr+AWF1MJZo8ZOTAGa7fOl+H3q5TSOD
IdTUalM7Q4gjxskKJ8kTHEoORjYsxgvZAlZ0RY0BRV4xLpG657pvelgKezWe
3W0Lh7DVCBrB6DlxHI8IdV5nB2daCUCprzfNUSdNhNdja52mvDQT39Jez5dV
B8Y1phcdT5o165qCoWEXWOFWu1OUSO8P


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sX7nZZsO/x1THpSY+5i5wsjS85KmOS33bExV7aG9JVJPkPtCJkACzjNjApQR
/DfuMcjtv6+yPFedP6fRE+1OJFIMWQTJ91H7XNdlIpzLd0xIIDVVGudPAsGN
NOPYCIHK4ip8hkW/Bx91oVB7d+jqWRWJ6kgKQe12JQLUNnB4Nko=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
q/qtCYBAKa4PIGzmb322agKQ8c/Rp5os3dGy5nxjVkGa57YLYnhJPYIMr79X
AGTKjs+2dEQJZzg9kRB7hppgL51jdjHQU0TSeNrHQVx1XgKVKu5ZoCbs1xSx
PAot62RZwJ24+0RR+qgNdIB4pVGPxtlNL219YlsDimjTqVkd/jY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 23664)
`pragma protect data_block
4ZMCceKuupXHVTuHO0+WyCWt3xypoLF+qLo/vVpRP9AydiVzCn2Shs45gAid
8H1rcBkBmBLseDhWIQAqXSHt28biuj1iL/2PhlqtQw1N0+VCnEIVjwtgfK6T
DMaEMjJ10WUhhujTUpY+zVo9hTOBXrqtIxHkIDUtl35FmVbRrjP+0c6NN2ET
uuCp8OCjrExf+VdhBoMOeVIJnhEs1g92LmpQXBhCs+owd7ZSQGHpj5iyQ8Ko
fNJi2QHI3pIn/IGvpP93l/0cOkmbzRW5ydmHQ5kDmRXXsdzN/7en28Lfwh5t
ICtw1vXcoc+6Skr8c/mFbX5+qu1pQ2vll8fPieLkvrGXqqqEerAYFNTlZSo8
otLL/H1hVsrckFT/UDmgAMsWi20OS2ge8uxYoAW0muOMTcydz+TOOXIgVFaU
xq9BD+4aK+lIA4NAVysbW9gRuGuOcTJwsxp4BXr+dRv579e6ib5kx6kxtpzI
bRR/a8kvmH6hWIJJ3gOP07EW4gAi8dkP5j1qnFYZhggVQq0ZMIcYls4JVJ32
hssA8EPMgKMGuaMXvbmjRx2z6Dwq57Ugzeu+VQgcU8X243fdhthnoVYQcrBI
P3ABKMon9cFxm1a02zfIs/qxBtYNwaBk9hVItFR9wrBsiNRkmSoF6pCSugts
gXyHJec1D2k+g83Ji2kOoQdIFdiSkEu/n946ihTFNXpvr/ncmNL+8KHc3gk6
1GqF+cPZa5QA+IBZO1sFYekpy68Z40rlfCPh+gfUAOhDRCYy8YbxWnRm6kcf
NRbFQdIRNoSXzV3BQC4hlhRwxs3o76aB6tXyKE8J13ve9Wx0STXrJk0BQsjj
rG5XvTx1LrNtnaAwVl8d4duIP306LA/8bZzwJAUT9YDMv5pEhZMmU6JVVc46
TYkf/ncISPkdsTSEo9OfLiY8uLQHPLfmXiM2nHsFFxJZe7rfiieQuyo2ZpxT
YZFboBPtvttegI8iTfhXtbdJ3NzHkUX+H1hEO0cnlW1qw3ljbaN+/Oc4YrjU
VHsV/3dPyTOaUlG2/4aRlXg+fNL3Ur5krhAzhuv2wR1ezz42wALUOcokKXsA
p2sK8alF5T/evxxID0Y2Yfip06EbrA/GW07+O4gz/lQ1+CKKSHqvIUV0G5WC
xrL72vCPiNk6DoGZwSRw3DyT+RUzpHt0Tlowi/RJihewkTcFfEkrvcGGWmGy
vhDqN/KqPpCqYQMknDaQ9FDsK56P7fKMgu39NYSe6Nf6/jhrIx3Fup+ttr/p
nqbLBhcgnu/Bj8RdAaSG83gRP0NPZOthJRuhZKJZyQXXDCV+fhzNZPpvLFjV
kKB8smVq1I6rag7qAflhm7W3TVx2dPMeblUw0wKt6w3sBJZNOr1BL4bwBfFV
gA7vx5/RRG0lTweD0N0n5Paf1tVLngcU62/bLTE+aeQVwlHj8D6Dfm26dbDf
f+Q9Uc6ekNh/JtCR8AjKq/vMLa7KGTKsJMQjMEH7GePEMHFQEURUM17aTk8W
FtadmqwZ9WPvDk+9EfQfvAFbkYiRdV0Aff9Vl0blSm+mBGxeGTOHUWefTOlb
zD7x+cWTG+z8eF6tEs1RKwYeor/3qwRoLJZO1IRA2wFRtkswT/MuQtQH5NAI
KcT9mGKg+P/4qJufAjgdhr12nBdsmz7fxXqjHhEbL+/0RWAXyUyMdO1JqUEK
VMS0Aj+8VqzXnKZg8svgd9YtH8DgxQbixfYCChOd0JmRA1M7q4nJzLEArLaz
76fX8BfKycFxYQwYlA4er1OYWxYws/JZBF29PEp0LaOevdTohLySMtF0Arpz
vVtKwqX/6C/xDM4Er3wulEsihgjxdxzrG3q7A0CTu93LnP7oGVMY3UovaV4Q
laaT0zbJeWJ2vPMgvSrLjSE1kmOTKFXBYRW4i0fCIQtOxM5wpEaZf35z9Otb
jmj30xEG61DKWNt21pqquscGMPLX0Ws/6PNDbJadM1o5gscc+EX59HpAglYC
pxGXPpJ7jt9qWg3zEWtDhpDlhujV2IlYCwjrCp4Sld3Nmqd+h/ZKlxxvecyU
/dBQswuPn7agxEwir8HighvZEJ4QSnj1ln7goTMgzDv93nGMvM85Kq/9xKYE
h7Y8pt6DxH8Ur84tNxVo3SJy5YMq45UzSsZJvSs/tMAhCZwX7JqIHzRcyQ7f
apG/UaseBrNScbkWROY0oNhjl47HcRQrkfcH3ReU1wswj3LxDz7EMyRYlWoF
80dPSIb5m0OwvRQh1uPXAs67yAxMwDq7gJgYFSVTbYPi0rLMXSklVrzptLOs
GAfZPxpYFu1DYGHOL9fKRiDTs7BmptqIoLbe7V34werWh5k6XZwBXxWJe26L
rJCKTY/tuCU+yUnSOEerdPMVgDWWFDe4mJnpOO50a20DZxohJ6Uys0tuCavd
hTRQmJkGfRHxIcImCWHE1lCamrCkHMjbkUYrwRzthW9/quZUl9MC3ggXQl1M
oDktVj9AjSiraD2tkXCZpGFsUe/ZzIL0b4WD94yxapsPiWRWRNNBJrn8RiR8
/wqByGgz1LG4Ss4jx9MAeVGe+YcIeCLNJybtvgvcHm2FGruoQQpjqfzBvjJZ
rvmChMqYyNMxGvfdFV5AA+4I07Qkyphr3xofGLSnt0wcxJIov4QDPJNVyGFl
N3nHbAZ0BVnZyf915DH0DQPtCzEIrHHlBSZLfRwOUq2sEqZ24+m1qc+8PG9A
xDF5X3LIAHByToZ5s5wBoxsJIE1sWiCia25c0yC3s836UR86fUpTZ4ntcEgy
TTq3UYfRK9J0Jr/9mzHFMJ2IpHZAAk4yrQmjhGZ3PrInbSXcea2OmcpHNJeU
9rHRq0cOUWJjVhPtnHHdxYFdLqxRH1U5O4/QfWjMrW1FPb3DkOLctIYGc+e4
TvrZxerzeZtuAijiCFtkn83R+bba5ZgnO5IgYRFe3aYdArZAvcEHqQ2FWNjL
EdUMXr/HmlOnm1b+z5EIrUintexLTwchg9g3KiyxLgzYK4gPRxY7wdLsVYyk
1I4FtoTLQf/CS0qs0DpxhYjEYFTSRds2y4EYCv9NAvJ98eE/zWa3I6TzjYvq
AZWj16KYGMKs1o9oC5/OqwdgFVpDY6FvEzxVmODAaYn0lHlzDkmooLmvLe2Q
lA6Jod7lIPOiTC/frISwHtvgLqelUzQQuyAif85BgHsh9Iq/VuYCKivAFTvx
YeYShg5PZBpPGvPJMTWAmHonQLBnvXYV5CmKiImtSIb8ZFXgA2F17RM9CI2p
hCRIV/Dm8q6+TtUiXnb5n4vYXCJ+B6GEZvMqrGh7+QHoJM5RDBP2xjC1Jt4h
sPjnOrRP4pxIAynDWwFh599L8Hn070Po/AAJrylO/+kwqbh+m6H1mToPOPcn
1FaHkySEJU+prTP++DvNJVAwzcHQNhJ0vio1PVvHEgpw9Z9yavXmEnUILBkB
gT8yQGnAVX149a9rlILS6RWlucWUvNpMVzjTcNNfGGpOBzB4kHrbl0KWirh5
a/kMbTiBQozqXK+aSk37bqB50VEts5GJq8Mlmocb5iUOQZWAawTWCv78JrSe
QDqAzHulpd7F6cLzPrzwaC4C0wUP2TDuc67qIgmKU6aWYazSS27tR9uRJc5V
JQVjoL50x9z+RG2/+LbseWoDNQPVRUqHcZA2jKpHOcdYW+5A5pjcVoW3Flqw
fCaaSQ8onyFtmBTOHI2qQ+jyA+MsgUbP/NdT6/q4TaMFuqhhryXXlboKudra
/5aM+Lawu47VhqDGlsTi2i/lR9My3y9mYw7q9yY6DrvH0rHEMVWvaMYAiN1a
6Jb5ikwX4pF0VsK/8NQzvGweJvWLJB/TsDYgMoP2sBKa+X3cJv2v/OQevmN+
DCXCx5wXoJyeIWvKbt4mYEGcfJaP2jbwSTM7WLdhura9GXFF++FWonaMBz55
xncE6n+xEPjbJ05/BW0yBZQX+r/wpxZ9gBARUCf2orlIP8FHRRQkg0sqikLV
mv69doZsz8GGttfmXbTQwkLFvDp/ftT245iBIk8EQWt79I6dvBg6Z6Mb8fGf
HfA+YAvySkRylTJd347lOUxgVc0Z8A1kJDvsxenk8g4HQH1MjiYVeCQs7BbF
HErSEwgaxAljIsMHaSOH33FD7yZRb9F56nZh7VVgz3zmPW0bEXFPzXmpfWLp
iSgibERuGOx31/lSOjjefAQAV9JbDUv/v1iqS0XjnEX9ZMSZmWsYBwujuEoY
XublJYEbhz8cnC70s/ZbZ5d0B2XHR+ci4Ce4L4o1094KLdj9oyGSttlkQw8u
mZ6p8S4oOsEGwfbkZL1+XpkU2fpQG3vcw2lAnw0+Q1FEsXZ87KZt8vmZqw0H
Um2N05QkEes+IoI6RrWzkQAbo9/AiQGlot09G9nWQIesMBJ8nvGLq93Ny31o
2rDzVUZTfWb9DO0D273ApN/tV0JmU4jvYsXCpiShRZsjkRirukHhQpgRGAF1
eWM+wTG0wJXfGsUD9eFOF2Vfm3j0UScWqB44MWt9S3LMh64yGznUbmOsianm
GeAVSMzjaIhLH6OCUDYVczRq1ipx0rclAc9jzBEPLgjdsTFb6x66n5rOymby
zR1AOCfd7nPxA8Wz1npvOaIwcKUDDV7diN/jJwRAvfnVocsDpwLGvDAdrowH
fitnDOVmprurV8214ENWUQsV6NT+4QGuT1R4ubCjMIMrPuMHLqvs7OVtJ+aU
oTskiCCFez3Al5eXUJgE46Wdy7RdTFpnSaCyVjRMDC2/36c+edQquD3nDTXY
qbA0q0HLb4XNorwFR0P9Y96YR1miKMoicWAzYvGmw/BX/BvR6wpB4LeolFPs
aNIp/NP8ky9tP6hCe+nKBXRP5JqcyccNWvSMHqkefseO58qwGcXj71zGRwoS
DrJbyj3nLMZNpQ5eOFZnFe9x67plQDyTLVPmY8ZlhpWi4L1zLUZjL2ArAinK
+3CMLVlceZm8R/GEUOufd0BejRreaLHWBD6L6FPmbWYiuGxFKDZSXvRZww1N
AKuvwUbZvRr2KwAk9UesWq/LE/wbrP3GICxWkJ8NxJ0rqzRbDK9fydmsI/In
g3hy4fx9TeVr+Y8c6T3BaL80p+7pWC9TUnsojFrJQncDgQs2iU8/fAdJbIR/
IHqhcCgxsZIuWnkXcUFVjxe7mNTFyy2dc7Hq5ntWZW5g83Tzwjw1SsU/NIbj
6bZAAxYePo9UwoHtA8SbK5YF3WaoWZUTzjnaN381z8CJFs0f3NvJPwz4Amv6
s8joJAqGc8RLFAmHGsaT2ayxyR+8l2XFwC3SP7/lGgBU7Y5HswPzwAsE27Jw
1fzEw2Zy1h8OQP6sf4DODNSpRPD3fEBgedPVutAQhWiRAiOZ+UZXxHU1eOhX
PHt7uM3t4wVqQ9n2Egpotl+nTAScXqBgESUHxhfFoy/xsZSKbNq1t66sg+Ez
Y4GHtH0+tuX8HxLpS5W7JQ9v9Ud6XaFsdTlnHwEi5F6M0hDaPO7C3XpE+8g8
0GL7NpYB00VIGnhynV/guEDTd4pmuivVL5gll2Tr/isnoOIzZb/W6b3QIQZ6
CC+mhhI92Sdik4u7sbmyJq9j70SkmuO/9Zz9s/aa9KJPwXPPPStoehrASdqU
9yUFgjXbx2MqycAmVWRh/Vga9Ro6r0qRCqlNzPSLpM0h6QdZE+lGMUha997b
FpK2XhLD2OAySz2lzQUqoum7mMOjoJ6VdRxjpM45jrPaxXEdnkSsb1M694Tr
v7LmspDirR2imR3cvkd9uZSQleG2xB3RzfuyDlV2qzPeHBhpNDYDwoo3pZdJ
1qzdzaCBz7Q7d/meBL+i0YiLFPTKerVNIYDkx7pGbnYUy/oy99vzTfkast2S
A/HGoqw/oTGgCsKPhx8yxBISOVXZgcRaSdcVSD1Ey1jgU/WyXgv5yZLkVbM5
gmnIjglrwpSFPZR8C2e0xF1E2wxtzn8AbX/Yd33IxziEuWnIiCf9TjuP5EQL
3w5NyYhe5QGARvDR3GIK6t9vFFQ1nqXAOzdt0Nk3OQYOHBMMzpoQ1/mG4sLW
t1SAe/4AAmUvJ51lJJju3WG8ThZWNISyL4ovf3uHGYjl559J5gnFUDfAdPtY
wKW+eHGwZTLkHEt69c1fnzqx9BsphkW1/mIuowitCbGvlCWmgp2TNTOsG/KH
p44x3bz6tWVre+AiLs/SbFTbhiyz3IbrLajsmm898AJDill1cFKEQ5Vz2baQ
ALCded1uHCLW7pRM6/aWdlhX8u47fqGT3ccqOdrTxLmkv/zQmSBAsdYYD4o4
i2fNV2sTGMfsqVh5DQcpCGwATflp+e7WZnov2y1biDdum/0ooXVbAg0hxpdk
cmYt5jBLz3I8vYfgUTm5mcUzBgZkyY4SGwPuYq9hkJz8ZOQZl/i1oum97MCq
A+O+MmwHSUZS9ojUjx45tuWVqFYdULDldfwO7MO6ARZT/okYNiqlw4eHZKiv
khn6MP2B3SCEi+ZorGIXi5EF8nUiTJHkVunsny0MhviViN4f1esmkC6bbPRl
2czXH1fa6uoC+y6H+31Xw8KjCowhYPyjOg0UNMVsuJb0SENRz5Nk0SD2esKl
ShUvWF13BZJn7qD0ySTFtWRwM8IG6MtFFkLhR7pW5GRI3q16AEAo/h1xXQXH
jQZkbXA33IIyRNMEgG0rFBBPb1D+COJgBXb7u5HywZfTAqKuBv68O2lu3b4N
9RZf1HV4A9kKVs6lFa5nMIMCdzjl75F/HbddKxyXZUPrTfKCavHaCbub0gHZ
30I+tjsOfIK9OmOeDGPBCfrJGFM/hS4cVhmQzxG6HSVff9Sl+S3pvawgLGYs
3SWM/QPMKeTpwKQkuQ3LwGh4ezh2v6z9H5mVWQl+tWyOnCxKGHNSnyohpe0S
OuA6Rs7+N6bHf5hsbVL9T0Yy4EMwArH308IxtUt0XqsCHD11CTRrpVELjwmU
jmbcgsLmNglJP7HKJHFcYIJXJDze9DmFQgUymuejAOOlmfMcW20Xxf9+6QRj
qj6pdZnm6HQq/v0B1oLtnQq2ADRoULiATX3tT98YUlRCumsH1m6R24bKHL/r
fxzU7/tPzCHsR3KFFwr0jAeD3jDTc6cJf99y0uBnW6M0G6/opZhx0q9c8fDK
5HLDaZsGLjSwYr2QZeXeWWyFcWJ3vH6wgcu6OWyCKJ55s0a0ENoNFZRffTD7
ThOzDVf3y5JcqiJXonULbFOEumfXzi8atNXF5wgKpqQSxw8pBj+sswWMwwyJ
xvMnr6wGvm1+/Uaf0nlXSpNVygkJFo4ZNZkFnMezVELrTJXpUwXxNudcFlHl
34EWB3xAKYG9pWgXN5H0I9HYDxIZOliHH/fCI8Ez6bPwzjyzG3NysOhXdbDY
4/5Qdeni/nKKK9lAwFKM494LRnH61PtV0H8rw4F5X5nCidFmIy9yPmNPvASB
7zu/hTHBmMSWpFreytYHp9mtRarOP7xVdkg/93S8PIw9350pDMel04stdrca
9jXrhhRSrgyvyh/Oc4tTpsRq+TnLgRGuK0dhReOwQZt0vkvwaFV0thapTtVn
oMN3qUHUI40ea+9mRCGDCerRlc4kT/WWdTBeG2tCfSXdrIUen0Ln2alWLe7T
5Fu0NGequvgClYbrQtd9aEMtWoqgXN91baYbP/xZwf/2W/voGaROtBrpzE1t
pf3tzDc9gSyBzTWD4WyfDWB5T2R3TIjpbX0zdBzITF2PEKxpiS1LA7f3/CdU
z9FpMMe2KHPnxYLnUICPTZsJ0QyYCZjr6SjXpsLINoNbI46D1q3MVN/Y2hE+
hL243FmUsblf6HmLU9z7+YseCwI/0mTNFeP3WfCBM6jb3zYg6OIm32a01FTN
0hVXzsNKN5/IKi0ESvQJw+bI3u7q/V5dFGGhWSmEnTKKSD5kSHyJTxDe07WP
dZEXlhd+a1G0Js2nwGClpL5r2/sSNBunErvwn5jeus04l8tdAj6tDDKm1Eo9
lUYVhiC9l7Obk8y3nHULry8oo7F6n0+rFshHxXHwiolCONv4F7Bt6Aoj6HaH
P5BOPW55A+GY6KCLlgBNhJqK51rlAkELFR6hizPqiDb3dcHFfobBm7AAaEkF
oFZhg5DgPisSrFDMLJjGnsON2Jk98BM+0foai4h0ZjcEN0V3UHFhrDeKtkHq
kid589s8iSEImnU1dlzxo1bhMqOojUkpn+BG6Ual11VjOWmwNckJwsRcgVwm
6M/1CQYCX57pEzb51kY0Lraf0W3Pq2BP/1mhnUX1VuO1v9p0mEVwEJg2MeaG
Zd2lgrCnc+BS4v55GkQY+uOZ3GHSgjMiV0xPZoeX4Ua2ZDMFj9MWSSI2sf9q
FjbWZ0KjsMP5+GmMnBd1IOisCmlOTyIIgHTTxVEAOnxjVihye5tv8cjym3iy
Z5wZqi3jGT2wEN5SXLLQIPKfTRzXz6P5GRpC5C8/15dm2H/J8HHS4oIBvxMU
g7IVz6EWvA7NbidIqgaHvevgJ2bZkt/BoYisbPO+Ou2BeyupIOxrvcslHaRv
ZFfSNOZtNEHH0x8QPbDh3NCKneguFIX5+wGofCWk4LxM4L18i++qh5jBlpiq
zqFhy55ha0ezNKThf1bXG7lYKqk59DEiniYCIhaG5jGS2+5ilYVosq7EJ33i
MM2vLJ6WR3StVLQiL6E92GUr0hwJNZ5Gk5DuXfVHhSV1CI2i/XIfObg8POop
KV+SKwFQBN5lo2YIxmG/oYftpI40+0QOl4Q7Oh1DzBi5CzJX8Wy/+kr8qhTv
yhHxB5NuTekQu15uIk9maeX99FL5mhYp2P7ZLpV2aLEvnIsX495B+ZvE4GnY
INzjA+YJv1LYiM1Ipr5vaDrOlhXYw9DIl0kcmbJvZVkxlbLCHSZmcmdIbPVP
3LFrBMm7IhFkHXMQB3dV9696S6qMvmk/brUnzWT5e6qxahvWB4wcqbLbjWBd
KBN8zOhSHSYkYh4H8q7cfYkljZWP5Exsx5PBYkeQqrvHNfBffrfGSKlSJRxS
c4EgfK8K1oaoyGOIzjwh1Wwtrl1ycvL5w+Sw/7oXG/hkThxBIrscZF0duVki
EUCLKHT7W50WGLqKKjNIICCurgU0ET55Vr7jLG/63sbRilJdLGYvr34UtztT
JZL/nFTUeq3RrePMruHINCBgdQPi8+2Z8KuvA/sM7SVFJYxts2Uxufw+186J
mXJncr6vm4PpJIF95xL4c0KF3zzf3vTbrGe6sh1fMu0hMm5vwSA9oOW99ZfV
X+PRyw68KG4Ak93dOYVW+HlPzUhvaV8r+2eR2kBkuqINLLbMEiq/fnCUX6mw
wPIOFl5f9x+IMyymYJvZ8/EpNCqNMBQFUuP46+Sede/9sxXUrKu5wT6icNCd
xIhh6WyeWxaviQWcrnqlS2MvKY7scD/iLQI5w1ih1uEA0q3TG9lB75wcZ/SZ
mz5KQWLRJ/QmhpHjx5Meqa9KeKN+kUsDEIHEogMWLAOEU1IEuISkPOdBvIB3
zFssOzApUin18sueC7AfsvWZqXaqaWloVHOc8hZXUB0qpkwVyxgcF4k7t6eF
arTWj0tAgT/YMrL/VEqrjg4EzDQDVYamaeP7Dn58RKUwUgLsPNqnddy6lgGO
32rKzEGkn1F7yv0SgZs/ED15lhDN0aONoCfAKA5NHRTRUahQlzPkWfYby0iQ
HBaFQC9F0TJjHQ6jZMWa596rVNyPGfo+Ohvl78Yd71gCBy/PyHEh1bvTCcIe
nH24yq35NhRFuKILW3BCfbgfpd/7xUumb7r73Qf1hweHVyJW8dizhePcx7o5
UCmhfVoBbSF2ZO/gGb7UHqiy68cFMQzap9EJ/CYjd/VSLk2wfDp09d4jV6Ed
1zj9V/FPc3z4aKVzuUA+tYF+p2cUTMYHi0VtzuMAvkPQ9ouw/mW2MuTh86Aw
+6MnQw/bXFUDR6pmfd5BgQpYfIDF9MMMTBXpk+bO9maw0WSo4XXTEF5yhIAP
ooAdRw6v3tdya0t53/mwmuJgwkevCGvsTrDiRr+OIQDnYhH8rZ8fqArwdgPw
xu7bVEMveK+axfIZoODDL6kDYuMBRE5id7m8C1V4k2H/XPX699104wwZ6odp
GtPUF1kBy9rPoltR70lOybjM/LgF5vjyD2Bq3ZLmNBfg/A1ZzqNMG6FdLGvF
eB9yMIpnlOtasS8Z7h1fvokZO2mWRuy6V8W+dL4uImF1zEAfHjD3lFHZPlGj
payGBDwAJEKT074RQs/xJmPjurfm8OHtoaf8MSCeFxo5OorvoPjHazz7VS80
lhpczhKJbtVlE/JNvIxJUoTiW0UenK0jxoms5VD1x9JNo2QaZzju5ezuGnrS
cb1oNZjAqrXQ5xDGSGmDusI4u3jkM3z/erN3CXjF1/1vDcCqwQmOwu9DDh6/
T/fkJSh8Ad0tnDcL35+Kgqdkrl7i0yVJFvBEnkZQbv5CfxsZECSSAfTbusrU
envTt7FCxhcwft+gT4/87ZULv8tR01Uxt/q/hecaMrO/uK7XAr+acZvhvP0V
bIZJm2TZbRyns15lKCm6rifcXfaZi3CIFvbPXaBQgcbOezNDE3sna6i84rCy
HFCTrG0MMufnINDRllc5h2nalMutQPq1wYvtrZQFxkHY3CDxEm8RBxDq38+A
4HrSg7cdY3F28hHIkTfgM8kFJ+Uk+hvN4B8CQcuSRE4oHg2TuCboo5q54AaJ
acDPjFhOGLPZnvz218LW2EcLmhbs0sM0HUzOppjRAOdpujpJQlsg4jhaxeNP
+QSOmooPp45r5C1DKkDgrawaIa8dsaxllnXHNLwxEUspLsRVa5EEu0A3v/Xz
0iTAICyqn2+sY8QWL0gtoDdMQWNs8uIkJryKP+lC5yXbNbhjWMjHfZqrSVXB
LkOBalG+3HCAU9yHjdQ9KFCSC04nbPtyXK0pW4bsCl8AP6Tr2lxmmoEwQSGo
sC9MxfHilmph2oy16gAreNsf2m+71L7QXZATYoAplq3eptNlLCkVcyF4fzKM
Tla55CAihj5Q5kOikrXw9HurzF3peoBCYv6+WJW7rK76G6nX29GOUC8mYSSx
rMs06nO1HQdYRT6TDC5JnXS/vNLwlez6rZ9Ol/fDoAV7THGxdxt/DrGW1LJU
QbkVFwegoahe9Qp7MkkV8Yxcqy8FhRjcNePXsiT4aB44WGUb+WJ/XeW65yun
bDJphTcgz01U8cmuA+4pXqYbgIelJIjvdUjWKZj2Vos84ZCnOFH5GBMLqTIn
rT9fka1jq2pNi0kFqvgZ/+jRUshrUHCKvy+71gCpt3q5ES0L2s73Y/1FucP4
IKcJ7gXGZM7+bF3Mh529J2vTbJhIjElGY/Di3O/DhO9bRFsGyu/x5/in1C8A
AzBP5/qi4bk7a3J7nu5P+F9JfrTj77ix/3Z3uKSOmO5AkcvvKVAYxpCfUcx9
Om4vl+Hl18nD4/tC70zOmYxOQ2rIZQd9fworSAF/U+Nl1fE7l+GpwenT3Cuh
5EZfOEOrSzzVety/0dVOQ89TSbpkUbth35Z67K6+s7s+yD5+8OwzQM4xdLi2
07LHelrpzfESZttNhfPH7k/lmrqsjNW5V94e5NczKuDHeIUwJ2q0j4wHFJQp
p+lIDGqzeUFilqwo9OcKRXpW3dfgOUOzdAMRS+6fzd5smsoshL7H962y5h0V
IlC8+tbn72pXqlJ9eAOWDTB0pmu3PQwL6fJYUFsgt8TsGPGFYwnCc8xfekru
psQ5QocEWP+zT6VwJKoKHAgFutMv+kR6ldbcQsF4B4mLWn7OZ+WzOu+C9mc5
WwJ4mGNjTXj4s1oEw75hD9AYaEaKZP/wVbd7/BO3zqN7ixu5ki08YbYS1i43
AQLO8r+pRw0SFmola2yh24JdjdQ+ChUfYALWWnJJVDmzh7ZcnAyvx3ruFWxX
3sBWbv8qOSa1Qk24paBpI6b8B8dJLJxZgsxzUQyZmEk97J1t9jy819za4HD9
RWeoAuYKGj85QPWQK3CdAdCFVkQ4btzwsj8ZGXSx+zPu7cLDfI/ViSx1ts7l
+IriUmnal2u9GsjySyATUvmxkz8q27W+3Jtvz3SB+G0aq8SGaIjJarR2oWOC
0A0jg5SpPybpmpF97bwYlnjmuUI0Ln7hTifbuq2ameb0Bmo0rxhqZB9ZFF+i
q0h/QkU6nhE6SPt4ZAi3lgUSXh/idZ2es2HsZMSEIOFmUUdZ3I9PKcL2kUhs
AEPN+DYrrV7NpnLi8DtyzqfNuZtsh0dIP+wRamTReXOii2h3Uvgcnt4msttY
v6fDPqOqgg7DRaQB0KC6FwHZILpi0LTJ76ZT5n92mW5WjPx0qZOPPhjSNhGd
cMbRiY0EYuiCPvb78p6k7rTarYvkfAc0l0pwvgdaT9DiUlzj/3A/9uknMmSY
qK6MoYLCCjnAVvFPFz5g6Z7sHOtt8LnqxeKtedTSA91vn5TXWE52qUsXaIv5
zSQice/x+3QNFCxrgPXEVWWb5MbNzWp4oiCw8D6feAj8EAtk9sySyfV5ZVI6
Ziun/XAlCDUr0aFvJsFB1iHpPL2yfcx2QI53i+cO/xCxtwdxD9zj7PW4kAdy
0JNejWovkEM1dxUOIXaNrKV5HDKj8MxvOz2RH+Ls8IENcWzbIWhdllm4nJO5
zNzbhN/thiRIFXrEKwoLhKAZjL33Swbgq7oIJCjSyYHaueCX9J10DROGSgTn
6bfAxX4UlOgOAVoy3LB/H/VIa/93nOpbFhHW+/flaJAROtyIjkgYCmDJhoOy
aO328MDHCchtNslKb9GxZ4g8OD9FefPXbDr8oHykEoPx7yCqibjuY2qDIdGL
kxMyqkID4NCmyqyavLmTHun9nGp/Zm+VZqDubNFoJ6xg9f9uffqXgtJEHTGC
8FspAFqWO99DSX97kegrhP1REhOYILOSt58iW7LwONH8BSjIEAf05HnqGjjq
TNrwCbFuxQc1NNArVjtfefcuOldGs7f2og788MV5ZJ8sAu154jBvi1kX4O/Q
QyXj7qjVNivv5AwxsiuHqjl99FpQKzxojxei0bLpAm4YcHpO3ikeaGhDe0bs
oHIEkGV54cH49Yat1vQWF0DZ78Pj0lvUSG2ZfwDofPdCBXyjE6uYhzfaVt92
p67Oq80DvdYrAktskwMMeoKN0qvVRYXkokYjJC2fWgwkCZGeaMNWdHULlzsp
64D8lxlnoV1OrJH9eZqLePzHCQd4qMTjwMKCYplOsuJO7UGSF54vKI4O9E5+
mGeyYXgDnxEdKo3fS/EVKp9Gbz8np7Ux7Fs3TduePiZB0pYSkdU0EE9fgONi
rpdlfFvxrbtCSi0pQplrjxEXrmVrYrg4D4Gx3KZVd9moOxQRbTmO00Fu+/HG
kpqhV9KEafYDJ94wU6THk0iopTiBj192Y/Hx90jKU7cQtT5FiIos8POq5Nae
xI16peF992EYzKH0/jgasiXoOWMVy2GQjJf3E2uee+IhrZojCsWeVpvG03IZ
Rbo668vtZAbbZHNdPwqIpYRZwkEEVuC3aV1XIlZH8eQX1rNu7pkhb7R3iPjl
mB7WpUSYlGQ/0gxCpjvrde4HDURDyi2u4NsIj+BiZ7+i0C5/ef4Q3V9W4fwJ
TQRVKga2ypfO+h91usoPrEP5rrdCJGLxLJw5DBns/sa0QVAxy69dDewVsFaZ
G5kVIMDkuO5UZ2YUsPGouzXAA7bqcmSfYO8osJjqW6IygX7oL2Z9cxpMhwZI
OFpF2EN4IFw/3EsH+dwYuQatvor6Gfh0vgQ9PWFXDU/M+mNDku8fdlDFKnTV
xQMudp23q7YJGCkGJslEf+8zSEr+FSjLYbpOflQOtNqypNTNzI6/GJwfsUSz
zCqip+rnTpjHg6yBdCjtkOZh/wUljlv4nEHLWb7d6rvj+7ZfPbOB3lGdqldn
WJkcQCl6tBL6KqWt7fOT79Jr40BHqjHnsJY4BQjN28IWxBDAgd1T4LM2bcW5
1JS7aix8jx5to0N3weanTdDhJIdPFM2FIIqGTrD48GP/HeJBgldb2Fsfx/FH
ie15KiRvvHlD6AB9qLSUnZx2qcDymc0naOK2NzEvduqqYCYGlvpXQ1l3UJ6w
YrBjSmXYWtkqj+h2tTHFXa8b5cs7gZq6ZpzeYHm7CofMJ+/ItPzBpOgpD6qX
KeikQ6G+V6vOBMoEwF6J/XYHHvtV2UXUYk25/SjNcceP0/0VtrPjJf6xIe8v
U93QBDG1RUsssQdFvA0xoc9wVPCKy4sR0uUqRfX/kQnKjsQdVWCtIJqe0NKK
qpRDXS5Qfpy0VoQeaE29LdRkKR1SDEW+kuu5Q8St9r/qc9snh8gzMKZeVqBk
FTcgeXjLlelKPHVu2wvfOAegrdCup7URia9aWoNcSvoL7AhVlrK1hB1p5EBp
8SsTXdAMErIoTBjUlKQ5/+uXY/OJhloVjhTm8qfUICufsEt/ex84TG0gOnf3
Sn3lhcb6Ta9WEdQeq38XDTT4yn5ulOHut45ABrhOMQ4rgfwzJANI8nmuJuIe
n1mML2vYLTbXsJyNmP14aMWddEkipOhnO1vqvyWdmEAGhOyKcDX2W+GTMJDV
NtQfWeSndAJfs1pCsImOLb7GK2JIYMMFNqnZDWwNSvROapk/3GVPYOQBY2Yk
Nk9E0PidvVXqar8mbWdSfSZ6OgLsJswhl1st78gGThTLuJTPuy9a1SQYb85A
pbNgH9TEFduQxZSrYd03VrxvNs6AqYGUVN/D8c8GAjOSuypv27uAJiva0jmF
CFC5rBGT58hgKB2L13RSdOAGQT549xuQJBurGRqkGTet4vzueSQ6bpRiaoKB
mXN4KMY5aUvo1E8fmlSl5I1s2LnKVYgD798sHv56MJ/XxzB/kppgLq0KkfYW
hOykQokiSqCCa3KAPpWoalbfUM/JiQ7zYI4rtlHIrMDkb7hzuVt/JZPmT0c6
7oNGVY7T5pv+2h6kt4xRBJuoZXWvYrkOG82NF3oqam5dX7eecKzhGgHiNY8K
yqvgdfDnmvtT2Jbs34Hg9ulziQS6T7/sjVdurFXOGV70BHNXnfQXaZridF/R
UrstGW5HkfqohepgkFXpKaAZxaooOZl83BMFTltiXix3tZ/IlaZJB/H5US/g
NfEqXvrkpxq8qiQSfp61tNc34kPd8WF46xFhWbEhwr6GsW+3KbNHt9/qFIkJ
pV8tPg4VYOrnZX3ayVTwnDCBq1zxU1w8ONuFjGzxPG/hX4W6Sym7VUfB5Tcf
j9sCJ5cT9sA74depuPrsXKlLsBcBQPf9BfpWMv/JKlVqw0TgECqbiMn/0yDi
aZ/+YOQgzyuXhQF7u6x/op+vZ8oBDTxOK7axYJFzw2memEMRb3CL2xeps8dh
1qLiWP4+t8Dpcv4Z7LC5bh11NoX0NdDPJMpdeU6js0mwwWvxO4Gi2CS8xDtW
UnbqObB9JUM6c+OsRmqs/28tfbl3KgcLhX5hIobdFsuqqfRuxLqELwJRrjNP
1uri4AkYqimvq+bT/gGZVs/D0y1GwNlXVTcD0YHF3tsF6xa4abOMqIq9Ueav
p2VAwsBhTeLpWhWp3xIfq5R/ouj53VH4AAM1xkvKiNChN6v90p9vqP/PfuLA
KRw6+C6luNld0mA7YvI7k0WN46v3M5IoGDZTYwkPEjjk8+FU7WThKY98dMKE
vkscDWlqrasmejii7j9955RTsObaF8XlEP4RmSQi+u8O3xJYQk7rrkkxmYYQ
foGRNO9LiGq077ZKRuXf7rtA3akpFfl3fxt8ha4r+qd8FOoTP97X+g1JjYat
ISJmus5z8zdUFXJQh4pZ23byXlaL+FVrzqSZOsSmMiHRacsUd2IJfNp8BbQ3
7jmTU5R8LF5OcOingpXSmQS+xRUzpRM2pdlyNXiaIfxf3XnSTqSmuXD2WMS2
p1bDhN8jB1A/QTS9J7bF5UztKT1eD5vYKDv/D0SCwCJiimt1ddq7L1NAP+wY
Mw9vxL79/QRxqkR+3RLXwiu2iyO2sMRmOyYWfTXp9zcdy2Bpx3zOIDIYIpPf
mdyWEQLyNX9GiKb5BNgOZXJy8/J3NSD67QulIul5Oypuvv9IiArN1IELZGbO
DnTPQmZxr7javkea9wjbVsxnwn89Sd8md3HmhR3VM37jafVfCPq3Z0UxaBXb
0c0hI7tPzGABaiVUVoyWQDhb7rzCMkhpD8AtWNvZv1svZfOA9NKar4XO0TdW
QJSFXDMwptJJmemys6SeHJBPsY362ESSUOpRSKJWDPodLtfMowlSf3MrKRaL
o0aawwTwEqOxUCZrgx2rMaKtNRV9Xal+B6vQzbneL8Lo4qLXREiLby9dv52h
HS8a9kzUEbx+6iXnJKMwk4yWBtlhKY/dUyTrfUELjLuDnIcsWOSQn8V4IYk0
FoAX3qOrba8fu/3yG4tr6LQUBtIWQZaGTYep9qdSPHizR+4pejrC7SYxM+8P
mPlLJJ7OXvtxFcsFaUlyz1aJb3mPYdwr28w0cfky+FJ+rPVgroNU09jhSSJu
CNgGYkQL7+BDuMrcCRVrQVfBzWCIsLg8+OMJk5fvpLI80L93SB/Vt644WsHv
vfDsHzW0kIKNCzEHHbrJjxswTN7FhLINlrjG15nfzeevZh0XVQJiBikzINEm
ahfhNjO0v76dynbVNOzmOGH+QUF81OcYuP+G6YJCSQb7czxipKoh748qi0mz
oEmKWiFFyXtoIp4HoAnk4ybftgPv2Yy1HGRR0NkcsZ625HWEJr+KUjD9NgRT
DBMp7w/zPHDRNYl+uXRD5ZRUKHEOzpOxA+i2xqosAMSEn5wYQupjzURTexvs
wJxHcAWu0wZ5v09rp8g4R9m0+/tK04HixfK7PqC39o1zTjj45f71Gl/7X6nT
cyTPriY93FOFMRnPHvklKLyd8hPNjVvJ0EkJbWlanQK9wMrtwF4vxprVuoCo
nWOsD2h65szf0H86VBR7UrTeW54EeokuzoYCSkxamtmUqtNvi9AhCV4lGC39
VUVuXnFq0v8MpK3mDTLd64CI/vvVN3RW+9JNwqtevV96s+JGmOaHuJLrAyVF
4ofbTt8ZWyS5Of/ILgvKTMqDez9YrMjB5hiXxG9YKDkk3TPTMIBFa86yRyD1
/g4H42Ij5aEXjiyUjK5GObX/NiWlwNTQUZzS38nQqwL8Y/oJn3Ozdyt8XxGx
pjAdWxbSJ0R+oDGVaM3YnnXGhh1mTUNQirK++ZIyRJylobxIYwHSslMZrXqY
DCGHCmW9u7ClQFtJtAxaCYD+uxC6Jk73pLV7B88DdMdbsf7i0d4JZOxAdEhs
3d9Vv4zbAF9EaQEhIr9Acy6gVeHZnwGt3XR8Pi/JpUob4eizh/6SzByMXmEK
J9TUVICnv2ifp7BM1vHsRAC+BtUegRlZVBzODnW8TfO0NCEZbHeASQ3XoVNO
/o+frCDgBiykd+hYeWFEcFzGKvIjKGMwvomVqVf3fLd6611aWHoH5OVFJyAd
Kwdc0Sg8QqGPB9HoLx0EqrY4dkEGbuXEodSycVYvfmYTqFnJVEwTX5sFnqda
A4k/O0IGkwGtkFeNyLH/1xAiC9OlFHmM3Ga6sMMdTFcbV7NhuTpkEeewjI9Y
DPKXGaAVUrJ5a6QQs93ffx+qX0I18Si8/gHQpBGENVeh8BIDfjRmUYuPTWQ0
y/EX2WO/1MsRBpLfER5p4sQ3lXdjAflSzfq423mTF2emgtuaTc0xL+XaJTi1
PwDUtoIPnoU/twNvSoOjFHnq/HSpw6mZiij8I0ehNoUAYLJHMWttOyIUils/
MBAZlG90LztcFzl5SFJTkZgqA5Ab1Xe0K5WDqpIykNClxx+6JXeq+vWfWJDJ
Lp87dvPHg01BdrpluKuFoVyoyzgZPyWoduY5knKSPsKdQe8cA8BKma6Y6l2l
5Eb9ltUzp+qwAH4xa0T3EfVUtZ6+gxJWemMVmjtSe4z0YsYqVa/LfAK2U06m
R/YKQUnjeW3PClNQVjS47hJL4sCPi+Ws78Hh9tSKjmalBf3FKBKyS+tsbLwD
Gk2l2D13oiTgcQ4lwDGT4rpsG8v0UzxljTzbgJrfXOnGqzVdkcoNj9KRyIgc
gxgFLGONhUAb6IyzFdkIj5ULPdEJxwN9yLm+A9MZX1LogVovZiuMMD52DtOz
rUxNgciW7fAiK5ICiaxyjtKtZjWPsBtbi8TW6NFStoJflp2nnXedwce/8AwX
EpPCvVgvDUpzzcZ1RuZaxWhHooZQs5IIma4LMvBrmeBsbirc6BHRK2pHQsxK
gFL2wlmk29+JjX17/WSdqZj82Y24FBiAOhWXcZEre9kwJKMIPbKZMG+BPG5N
fH8+TM94j7OL5lcMnHCi0t/u3rAdHR/ssaFsGwfjOmPP74941D1ojeX1Stqf
Atp9QOdMN0roB8JEVM0QjhdwBW/rvMYXJdNKLF34LP99JO5aFffy2CFgi0nF
yaT7ZJi179kgGUmaPlKP1n2Ec+JRvBesjug8hWI6XCTT8N0KNCadKd515vn0
Bk3O9AMVJnP3Zi7ozPGT5G4cqCHMBCHrjeAaRhrIDY/gupQ/owOHBYYtU7uY
sbUQuoIH2q+0JJavO3caIZsb2kFcojBqLVSTDPBiyiNMiD4q1/wmqaPRRGLo
xarwVi3WnR6i8tIQ2688SuHxyeQZqSf8oAuYvs+r8fMJe7iguf2nXYGMKyrh
t7CRGZzOXWHxMi/hFmf6X5dEG9nSt1w1J0aSjZurKQA7/TdMG62zduSFQabB
y9ky40TV17iJCi5kOibtsB1kSnQJKE+Qs4HQijlGDh8Am24Ycsbc01ZUQ2bT
YRedvDBs/HKN1VeFkkJoBEFbunLLllENiMi4MdeggWkIYuBrjyCCq61lclZ1
0vGLH1qhawQURBdxWI71w/J2xEbN8yuD2iQtO4zFW/SUIg/dw4FFoc0I20D0
6+MTW6qtZlSfDdxL39Gqm3rZELV2AMtVX6r2SJSZ+XNOnlc2JLtCifPY2IUr
VRYFFSlO8uaDfUjocyn9JbMCOyRvFfOnncdT+kP3dN7+8gf3uooBp1WICS0b
MHUGWCriicTOgz46dT8sF3R48ID7pnZJwhxWWQzzW/yPtFvD6KdMJtXZKME+
YFEiUEPhj2hpShapR8z3J0ZnWwP1SO3T/NLQivqj5ho9lElmlsr7btLqPsgP
siv+KT4s+wZ9sMFbyE42+YLkGciEn5MkzVWcXbFy9G8gWd3o1yMXr3Th30md
2axQ80mEAFLf0+oOVyyOVuS3J3iHeYo6RqjwTrKVyY/VbbAJWUtuu1aq/Ker
wawxQCP5KP0e5wYGOnaGYE/jF/TCNCi18LIfPpO5uaDrcUicAxgGkZdtI/cX
HdYgCNGyb4Q5AwduoGxclNEN1CuF4mc0uiQsW3OVQYowzOM5af5AH33OHEsQ
JEwx05yyM9zVS0eX3s9hGE7OES60nfr9tDRe9QQAYLRZBhnehJ4eViDhQm9O
pRH3+e8B4HIAH7zG5jul8CiGWcZdTnCASsBCTs9PSY8cOnafEG8k4Q/9YXoD
JXHDrZwv8GllNjkmErcy6mZAD1Pb815LkWBoLyS+2cDrR2JbnA7+NUK8ybXa
aKi4n0L39J8sJvDXJ7JBdo5YWW8/VTgI31h+8cBnODLAinBf3uOxbyDganT1
wLj/96ZqOe4+8CFh+9GFFGJfWtH2ykmmpPB6XU0A5Qo65C24HTDGhSDp1qB7
hRWbGo0jxm71tfm8mmV2w5Fngip8jqA/hKAhK8lpGNMJn4IwfkyHWQh+UICD
bah9aQEOeSq0XBLkurFJhX5gjBxZF8rdgEsaIQM6m7TAWjylOuglQKWc8DrZ
iKIRi3IDOxLVWKW7b42KoGjyUHy75TjJwAM2jV6qHklhTqSKQZh59nwAXKvZ
k/lpjIanKDBO3I0HeOR5LFg6HaW6iujAtQvshCD2+guIwf4yRg1R0757zl5B
ABFEBWTE5msZLc3XgUwIOLPTGK5hphUVKCu7+NGRGf18TppAZq4+GYbsRiv1
trkAX81PXr5faRLsOFBIwBZiDrH7Q5fwzMF0Ql7z4PXSRNiaXL+Oy1OCBKMV
/gP0Sd9W/0g89hpHTkjOvQypJjHrpqtnXRXPBehV0JBL5U7i0iQbNHXmMpTV
OdptxSpv6wgm6nfZ56AUj4tToJxM0mcLz4xqd2eI/p+KRbcd1D0iTqGzqC2N
4tMuvuMjvozeVVfzWsPMg8alrFHaRUmMaUukZmYeF6EYe2cqBVLR9D/awQQp
GUj9SWH7prBJjYPUseWYuLXPp3D7R2v4jhPV4gBrWYeawrr3YYfNBdvgVypA
29J9jwGpE0o5pLafLGcb/POxzqr68jaABi+WUZbtkI5Z31Y3OsuwOx6QrSge
RZc1ji4AbMdoKTYW0if0Sxsbt+dIDusV1G8oIB6YMNaEEvCMLzOrnArjmw+9
sjRiN4IapOlSBiT9a3FCz7b8Xfk+xTQwqCK6ZKU8QRFvfC0HNv1kGUVb2pQ4
E+DwmogLDRh/tE2ao8fUM3qf/8iA6t71TKMnPSaJ7uCc+XiIBgoCb58w0BOt
HTXxtgI0FH8rkx0rzxYg5N/B3MQ/6Z5YXP6REVnSPqJh6fli/pFosRi/pqB/
qSspzS50b6j9Bf9gYSrPICCQc3AeTk3TkWOf9EeP2FK+nAvoockl+6UlEf2b
79Xh9tX8laReYrhOOByFQJ0DS6Z6cWE0LZQid3OZNwetQDIO5n/EkEaaHF0Z
+FMJY3jICF0Umc9RDGJY0vBQ5UlzxjvHBsGt8NMpOmHrH8mTqn6p89KCmBeM
EB2a9G5N0q/CQZO6xc7rBtealLALXxC6I1YDxcHfLzKp5MQACl9iG2/FlUJt
M7JWfGCl+y53asm2MNBuz1VMtEX7VYBGOqMSMYgS0xow9akYXz8jEOT/ru2u
dth+htuHGE+BAcfgNwaZKKxIpzn8BCfrN0w+w7oKXh2xN97ED67oHyB8N6sw
zwFPEXWFil20sP5pRlU1yNEpOkyGbvjwYXNv15REnGcSgisD+9EbMm8oikBK
TTR92901TT27gj6W2sugBlRt5nE1SaLThzgYv4pnhiTfUQq9V7J2abeNWKNM
33+lhDKhToRsGfvdhdTgsrRWqYyiuB0YhZJJWMyD3JP93uPmm9B79hcJ+8N0
U+Xkx0nv8s9sxA2VefSDHiy3SZNOT4vZFtDqRreREjTOcLWe4IUwltAtfx6R
1vyOPk26XYDdtJjX4WuSgJl+OydQONlBEurC+GXZzVVFev8Aw/wVPSwJjIG4
50qC7RP5BdyHDXV9ATADJqxVKl5xLrnrrMzyurhpBwjZXRtTCxfu6at0FQ2n
WNzHAiiJPDdV2TVg1kJiQVayHsykFMc9pIsmo4IOSRsUq403UwoekmQT0A3i
N3zWvjAn2if3z4O9K0nF3hFeJZbmg14YRpkbGwgf6QgBaZLNCeuXEehG+gO6
B3x0wFiU1OtNCMWP/2tni/TjXRWOwtQIbl4/rapyfuEfdIB/1/0IA0jctcUf
KdOFMdVZZ574UFHon/sQ1g+SWMbil1ZoMxfAk1t2zGBLg4nZSjFraSKSGC0V
2SUQg9pcDZHjKxAX4SDk/c0GM8I0jvJPb2ZGc+v03pHLhPFbWlLHNLcSWJq+
es0YHKyphULv3dOLUBWHXRmZYOVCpGgVqtjNRtswSfQWomZZwIzz4JiiEwXm
FSjs22EkMMBRUBaxkIGqsTFzZ79hhGf3sq6yj9tuf0kVGc7VTZf5/EPVeg5U
2/AlWPODQyBPtyQCHXE/Gk7FXWFz6WzlBrmySfDb6PGLDwG5EXEmjOCahQDq
ZKM5ffsuKDl5HqPMUYs9OEC1cLOgq/9/7pZqmTSpEgLjPso2x74E+W8YCXJS
KFMU2IX0Epuge/HbL+bhYw/fTYfPkjRi9AEyZ+UOvEx99P2dM7FHAcYAEC60
8aqlK9ke2ymPfNfJXKmqjCqRh8nYTRjCd8QpFr0nMcpFU/7ZrxHk+KbRI+9m
djW7OeprNCMYtFMK/LoqrtNLB4BkJ/Zc/IM+Vp6N58+7Q79rYkKFcnkmbuTG
w8pN1m8GFb8nsfBdsX9sFKVACGGIeJjDIfL5nKa/nD0UDXzy4vtMJnq4v9jB
3AByUbqXkGq7ozW5xQCtd3lCherjp+xFpW0qbzKFghAxpadt1f8qdF4+5URc
70qnGvycjZ1ZPrv5U/zJz2ZQ1FhrCDYjp30TBqlFkV1CWto9FW25FPQ4xikr
XuD0QMQATzwXZVTkNNoa5LgDaI47CTVWHtp16E50Act3cMgROrZwLwMQ4lQ0
IukzZ4VdqjuVeMkqYJP72fUrWqA0pB5Oq+u+F5b0ZJO0vjx6ewD6srgCD3yX
q3b6BUIumodL+L+OE1zrWAnb9ZYp3sNFdSWMLoDV1J+ano4rtj4rVF03wvCl
bSeRHwhnqoDlwhhOc3/3/stR9bw5ubhSUVswcxPH32VnSKlq1xBY1fG/HZ+l
s5gT8QSOo8kLotGIBj1rVnyO+wlr23O4/XpLJ30jKKYlvH3wPo900adeY6IC
1584LS+QcjD0O7KsU+vYat245zjIqGeB9T+/hdCSUpV8jJLV5xn/uJa2tUrt
flY3rxliiT6zmbUzNVJ9iqIgZh3yPbOlGLBRxmABUgUSmH95v905Ab1iNpJG
dhDp4MZtA1avQM8JQXH7UF5/OEviYl7zO/8vYR8X6WEIeMM9brvf99xWNWjq
iKudedm4MHT8Tpr7OBUKGpRBf9wpDUgIFkvjoDiIYh7tF4IF6FG+33Pgiohs
Em938OaXc1Lt0tiv2kF9cAHM+/uF4W0lk1gJn0vVPpxNeW/3OcVezM/YxJyF
i9hkPUmbL3HgFrBPAkNwCubjhVw8P3PHHWJaNAMxAxYdXNw9y5LMxQdyqfXP
P/u4Y/DUOxWsglh1ouYL43m9fDPUtXx1sSQKpo9vd6C3pcTO2JVy5hyH1jG8
JPdaxBOQDjAy6tNqIQt/LXdneR6f4iwQLO2OCMYQKzb5Q++fErLDNvU38hMq
v127kdKRGzZrmmRcU1Ciw/hJZBC8iOVQXXc9rjp0bS+AjLbQX95sPjJxMXiM
hzb/LeI+zcaBUpN9qHx63F8rABCybtagmV9SwClABRBweozUmBZ3r+U5jkQd
R+eyrpAdzH0OXHdWR2eks5LW8Ha7H2BvL/kohsVa+KFp+tx1y0Ys1Im6dTe9
Nmv1kmEdcFGu+yVdcPdsK0VVwvD7f8LnUnQBvKKjWtZJFAdf7BdeKiIDAWMX
Up6xpNql2QnvUyqYRMLToD3Qqzg572BWQhR1VN/h5m3PVqDbedbDObjGqj3W
Ch1oJGf5iEDY2EdB3jq9fpoYwlj8DVL0VAdRzVcJQtPIjUXsNftSexSI9qZl
1eIDyehG1YAjYgxRmhnlU/0M5Wum6B2UgDEdIhmRKDTJzcbmliyRl53uIqQn
+AWKNGgAbEl5rE9Kn1sSgyTPEfPDmQCR/NGJSQ4X1SffySBJ/wWncJ/PtUkK
tS2OSVmm9C2wxLDU9iICPGkYsMYiE8MAV/E2bK8qGqBx6PIwjF9IhBYr1qdh
+FfB9qHuLdSO4lpE2yFOj32k2QjNktT+3pv/GIq2xsvCKf7f5WfNrZ4wh30E
t0CV4WgQTEr+cz2B54CG1yR1nt5YZ5NQ3aOAR3H2kmAqsXajJ9p3uPy537Ns
OdX2XuffLUHU4JXvAenIBRI61LobOoc8Em4iOHOqB3k+dKuYZaX86TDrHvi0
97YuBBLK37HVNKF79sNMkQ48Eq0eOyQP102smpqEVFdsHhvwwfnesm8L76U6
mtCLEhgzCz4tMbOS1D8jaSolMl8P59mmIOh23PRmTncOXVBM4oLDonGO607N
BoDQNOoj5a7tLqA6p5XGznNwBeg1OcK/pLffFR+hVlwLTgJPMkwPSElk5yNG
LAzqVxgSw4JCJV4lGrGmhV4apHq1hdLDWd4l91sK+jsrIDIUHr8DzHgPBvOd
ayxWtJVuG9G/17mEqPzVgv9yJUklhPtvQ40Yg1akU1R8HhiwdpgoTTAocseq
1zSU29QSNnbEdrG+V7eG+GPFZuXT0BgBankJr0LTvXays7kdYp9QGhPYt/IQ
VveeM7uQd3Z0TfrAaU9ffybou8Tq3E0H4Ro9L/WV2KH0ybU/xZ6dUfxi5evD
M/7nfdTkGXLSL/qJpYe5PFZ57vKBDRDeTz+QFTu0bqYj7vS8QxpZ/q051oC7
oAKiupCIgXy2XG9d3ykDnLjmIOI9q1ArzgBfglMR35V4+xf7UwzZmGc1hHPc
XoPH8UbR8tP/vqs1oOaNY5a3Zt23VLcoROErRemC5tyoKmt/kF6mQ5TcTeYH
2PMCj/ZKOexliwtXwh6W5L7JJBYf1+JDW1A85w68diuQFwR9OcTMzy8hC6os
qXNyZA6PmP50htQM0xknEv/jvOfRw/CKgjX/tJVdSPToyVw7ayRrF8oZJZLt
l44by7z3k9PBqN4+kWHoYNF02cPzfGc4pru1iyXTYeWik9UcvE3HXCMIp9AB
S8v1VMdfvLn1iiWO8Qqs8YrmFFrB8qC82SQNH7KjyKvfE+5z3l+85iUw4FGu
0o90br7yznl3UCRi5/41B7SZmHtZk2ACquOh6hcJosoNrQjooT4w+LagqTsf
eeW562goURozNj4ABM3mFzeFfxEclhfSTtFHpwi39fnes/AO9BXyeTlVYnM3
ND3b4weDwVIq6Sqz540CgqpLgHCPcT/nwos6visXNsT3BbIyGUYxYJZi+lSV
aQUO6XLGkcyVcOR6OLrZZZHr249x+fo4ghB2eHeS/MVOfqpoMHjgg8Q3n9Ku
BPilLsO9I+arzBApfdXDQ8lOYgy4zA8RmjcrqXFVOZ+1arhYGUgELMcYudF1
ffB0GrQxmZwanHW0iKyKko1tVhdZrOkvb0CKxKtXEO6sO8zyHdpd7o7hHt5M
kX/sXC33YPke77xjSSnjO7YbjUydedOkSkpu6Z7gMByaOoAK9KMKkDTDt7f8
Rgx0VdM4vUHaSzoDr9+OfK30L/XL5gXOp+s7lmTjRI9/wVnyQwIBjd2NjXqf
WYfV8HHCiznWhxoQKsJ1PJXxLnuIMlEcHxxvwO6VpxiDrk9X6htkYSe6jN7p
Zy/yXgk3v9fAak9yGWuKrsLPng2O4ujmurUfSUZwaUNpZe79qCG4+jmNUGSB
TLjvtLNaX/JTmgAQtUvGTBuasN8TtovL5MC6wQy2UTM/XMb/n5+ZDtsK0De4
W32qTifh16UNKgBuk4n0Ds04IWYklGPdUESTtFukYR+0ytt3PkkUL+KLCFtV
ingo2Uy3xhCjFxF4V9zH0CoGyyf5ot/usXfA3+SF8rI0TgafudSCsXREbHfb
cp7riwab/jjJPyBaX7LP2IMOP4MQX8nMpGcDMxMwFGZ2fXeNaWaLdBGs7Ri5
ihY5ALvFzbxMGqXMnemOSounR/Kn21MV7ca35Iy9+ks7FF9UuZxO0Iz5BWFM
gs/HRZLqtt3aWLzqgOFOXLLxXBdO8PQKiT86WRwpHvU99CaNbjtDGx7tSaNK
LCIQjvRpfYOgRCnyC8f8JdUFQHF1i19xDvaXxZ2hkW8QRo/IcBu6hgCX4v5J
GNYOASBMsHXd/kH7g53FrrSZkCnH/N7ZfExuWUdzVCwIOh9giFyCkWKxjUGu
CTxJnOQvBIXVSGS6sTXKvMnlcu/E06zVYbV5WJML37YCnzdio07U6LFFPkKV
b6lQnubMAj+dIrW9WMmjmUiEuW3xV47F/S3Xg919rsIhxujfckqwbGnCdzRo
Env6ViLpPRGjP5sWLoRQi+cHUYwn3aiOC6kj4gG77REqBkSwdQdbv5mqE/gT
KLz+1QNCsRsOWJxPjtaX0tIkgsB/40JHF3RRI/1C7N9OaZneHBxrbGRkYIpi
olUGqfW6VFi0EzIZsQWTfUDsSrRE18j8H5JxULFDNL8H8JwMNMWp69JCi8s3
FlLkO50xlp0K5O+DtruUGkRqv5pCIDseB3bT4GKI6sWhk4rvtVQeSUOoZrG5
rEMJrOgYicBEi/14WKbSKAklAyozdgfGFfzsDZTuREAT2eiuyaOyVC4wa/R4
ZHkDvknYbVZT8eHcZfGlrOaTTlHr+aT/FxiL11zzG3yBi2r/A8g28G8IVYZS
JNzsvi4CG7ifOQrFyta+I5FbmSa2J9wG+Vxoz5RODIk4DnRAfHRqALgXdYSn
TbWvYoNoKarTWBhr2q3Tx8dvyAAEnMSOS5kCfWt1bh36wtQcyfTc/ddIh9U0
gcACuLPn3bxpF08dz8r5IDkmA+bbwyLlK72j1WmbW8Dm1vBwb2Na2tFfHlSf
xm19KKPY+KXAz+uHA2GfLtULujHzajBiyFjqP4oyGrK0t7WFuAYRjqwJa/IO
eKkdMiy6nam7joDSWWa0laouFuEDdz/bnaxmvxh5waM2ckJeXLB3h+HiJaSo
PQKyACBuUEXQ7MZSAx+CFTg8yVwmcpHFJYLUfbTmP0DNfy9e9fJw2JLJhn5f
0YS7tsHqjq9mBDrEMFeODNIof1eaKSJyGEFr9cpBDr0pvpXJbk+6rSO5h9Jv
eYq67wHMqWwJiUy23jrNXxU1KGyVeJdiz8DjSt/KyyibpAiOZvJVePnh3F3V
hgwWNB+1IMw5vxauPXvbxwUXUA3aKMfIrBS2D+OI6nnBzbpeMpKWta/17S2x
4eG81hicyLxP/HP0CAEeL+EhHBMyI16mIPSpKTfSZ54JtliNR4HKdoP3dB5I
qooUnKgZMcpFmHoGUoDwT7PvD6dWTOEgPbeuiIVWiWD4P+7q3lMEfGrg1PmS
OTgP/Hue4EZrVJDqjJfI5SxehZ+EOBRWeUEo5xf44gNp8k3HrrfBpQsbWbNO
MehccMohy+dpvqW8b7iiNC+SpQOvyQ4fw/tnD8dmprR+Ltr0eQjqS6pO4cCf
0SLsjXIE2UEpJeVhbNjoJY3c2Dpjot7s74slMeX77RDKmUpkuwiKEVsUtkhq
3KsMWsQ0Rc0UT6Y3uax6nziV+e8IWH66fl4J7rtzoj1V7hJYlNQwCRrZD7DI
Tt3s8QzWt0wFmuDOcKN13lZJ8E7NAfRPGslZHAPJzNSfFbHIsyZZDh1p8TO0
E0CB9Vx/WI7iKzh8Fe4ufi/X3Bqil+Li6eNicC/nyvQ6QH/wQnvEXXXWk1mL
BsB4CvgK7hs5Y5sNHuTXNV9Pp37lmsO5ylJ+OAfFpzJi+cwYMsOM7R3ywxuC
FnQyu9sYIjKeG6ZNsHkkwO/Qlo1Q4j08xKXb/m9/4NUPNy6DASfVQ5Z3i/LC
rnSghDbA26kNy5XgAQInmQRiwAfOShvo/0pR6SuGvHpAqmyJSEbxGKcVUMOT
OFBa5d+vFtH2lJr/mvTWkmIqK6enIcjqkZaDuSCvHIotWyeB+78uVy48W41k
wksWjJyBQAUfJLO22NoD4NlDmYUe8aAn/30D9f1gbIA2twuZFgio7bvZKJcV
I28CRNrIN3o7ZjkvFlT3f8ytpKzBT8FmaEUeQerVzGdBCHi1NTux3XfmmSvo
mwf8asWkhhWV5A5IT/3H2TZ8OumbB+wkVPeEgzCkCKV09cb8zHYWYsUjFhz3
VYAMJVglqIqE5DZlZHvkG31n2duLGMXjgLDd7hEoxa31rP9dVIdX3bWEWqo+
BXWvJOHaeoobi+Ag5FT9jDkvAc4xh29hZG71QhEtjs9kWm3ZJB/U9CLRAeKK
clhmbta54knVYhnp35dtmwBZ9p8MIp18UtWZgkV+rtd8ic0dRxajyhnbifa+
A7M+7wWSLM+GI6u/ZJbPxLNYG+6JORM5u+8CBnm5E6TOrePDlN++wybp5BIE
j0bfJ1hK6OcD03QzE9ovZCpvC73jhQUbhsCVsz5xyQjLoqt89+Vir7/L9Lwj
IaZrvcHWbJsvaKPEJAoyQ70oAxOebpIrig9SdiZfFbWlEqortbA5HJ6CAJAH
5c8TR5fRhCehGC93LbYNo/1uGOxylrz0hMrQZFHmrzcMO014BAPzYkhlYZOO
8UokOGKYrHirjWKdbSrGaJsCFfLXr1RIHxRVxSdW0eIDUJ8JiS/b8ziiOlMq
t8y5G0Ih8muyWmxLLy2vx4yH+Ot3hfo8SQ1XiwXdxrjmPL65lI0vVSTqyfd1
mTWJFT1xBKXk8xIjD2hJP1uqFDKIMuyFHeFoOVzzRObbrdmL+w7700B4t4DR
tBwAXnKeaO2qGbs+P96wvK3fqbUlH+lIcGZ6HKVaWSRlx3CBe4WJWoTyp8q6
/ZNARXvakVbL6E1QpeFa1PoZJGEbwE87QyHpsRlOxLQUe0eeMwWXC1qMUGJI
6SBfbLIVO7O6byKULTgN1PpQJjsAouHzjiiFtRIsoXcnkD9ofVuFLWvYbM8P
g8bLYugrtAIMSrrO0si87pYqkjS1B4/fWT0RYknSNND47OcL81regJnAbuqF
PHiTbewBUZPDtu/NkZ3QnjecEwNG8fjXt2eFzAOi/fQ/ZQflmwVgU9zmtnKy
5RMxkj+JOth3+OzJTrRq63OdmhOOgDI5oB0vskIk+aeggThUr92bugjl5qoh
HMJbX74lJ5xCjJvJS2pQt3RNHyOvOaR/c6zD82lKrYkQTO1YHKBpYZYlE+Mm
u8JFglOLX9TSK7p2cHgmDn8Nm5Ls9dFbJpBrp3Q4AAldH8YPTbez/aJNwRWg
PS6CemB1Fpw/AsmMXPVnTLI3UKISuX1DxBHx6rDE9qn7yJs2E2COwpXKhZEF
Q2mE2G27jpjpbAaqmfsihi87VT7apcDSRs6MaaeavsGv5QN5+K884lkdlqoG
0+YZDy0gDxpgckRtSa2Yb5vbBpFBfjx+Cne07AOtcMzWyZ7I5kMf2iS8h6A1
k3LHeP6KZdOoMrxVz9Bx71cGhlRzcpck44KhgGuL6KQQS0RzTA+SsrwLPFre
bI/WhiJJZT5IMkrIi3ToETMmxCpRGcmSkc/qysUlmjWD9U2VU8S0lFf+M6R/
Vx/k008sajq/aLCo7sOGkoMc7lC6VwK+Jv+wA3zlv4KIIahSVz5/8RzksKuL
/Ig19OPZxqcA4h5C85Ujh+Cz6AWqTHg9gcotyxSWMRlIClxRiI/EHlkmE5Fs
RRBInM4JWy2edd07tVwjcfjWAb2eCiJiRlUGSys3IneoLiM41xWaoRx32LEj
UfuIp0RkKRyxs2tR1fZ0FxXQYIMal0pD0A126dNAVSmQLfFhz8PlH6pbUAzJ
8vfuejIiTLT4GFBmQEdnw9LjR1T7tG1yd3Qzlf57YiqTzoomiv/Epe5GV7BC
xoY2X1ephRQF6nr1ULkh+ogGmKoX1OEfdvg/uyOMntVYnMuE9eInLLnRQw2S
KkRIhE0WCeyEwmeDXRlzhynv+1FG0umOkwQ1fU4DYI9VdFD0NbdK6tlMcYbP
KT0z0VL6L608HPjjzXKpqF3MeNOXNzrnmKEB1Mct+sGucNeegOBk2+1+ZmQ3
wpVGM3FohnH6PldL79CaoEyj6M9U8tR9F/tFOVGJxWs3RxgLQJRG9oCv3WOd
lGL3b5z4NFvdzHvYpNjbzxtuubG1sJGVBXElSSihfLAZ3VScq465vIcSoeTL
NzZUTsvwJBQM+Cz+/UmPBQeYDze1LN8qJggEnzQk1KDvH4wyIAbgDek4v5Es
7IGIrZYOEgxFWmC1zavpfEZ8cJNH/7NZJwMkXI0pKx65KC3X4AixGhZ2WLP8
6eAwnSreggy+ckDil4UWPZ/egdwJHvq8tYQaG3FjIVK4pTITRqW/RzGw/r0C
dQ8TUZLhkmCpDukGN84lU226zblxaCP7Z2IST/iKvfwO8vS7rDz51lcD6/mK
cu48bSOYyXk/8JE8oFofjnFuBAHdIBsnWkeSEAdQvKdAB3WwnoNEXbYvtZLo
MkfD+Ie02Q4toR7hyH5hltybD0rtVZ5Rc7nKdgAU6TL9wb1Arp8R0D67SIqU
Eiov2JSSSlUiuT4csCUyP+hkI2UdfOPYtkeZFz/roLZFV9TfQOznv0yjH/Q7
K0P9KLiKN4dAmXPx20F6EPKjvafbaO7CgObIPOOylwNgkd92zZpSm6JdJl8A
OsYvPPBsdFAATkrvavXRMSzGnClXeyN4D0cC6nlhh8+kBj5DZa9Ww+jsY8CT
CpVtf524wWPcJ0yPQciSKxFZDADHv3xVKaOw/k9gv4Vvl4UmTL0vqq+s33Z2
HpQKtj+kuVnQxILozZ41W2mU0TXVWxpvYbjJpZ8qiulS70QT2DYKZhyxlnTP
5LJKXgOcuEqxyQV3Ldbg83wxEe9wZHRIB7Ofb2Fibz8AZLAghjUia2chebob
QCEdlBsPyORF6J4cTOE8x5z+mJ2+FicvZkdO0KcMYaMqugQMV75kw/fk12wq
MXjLS+vreRFJK1MltsJEQNnPu58lJwGQgw1LVpTSonBCOfCKKYWcrjydITiz
QXnuvTNwD+4sTOkGQZUr1rTycuUsdV7z6hRLh28gbqnV1NuoZgVwmVMq88m8
YdMprf6siBD0NpZTdRA+CK4fylewW8V4PMFwvb5c4F2u5OhOKWSBYule1Ikt
bAqvIIAespkKugcSDcwnkMWcJFhvQj/NMCzbKoS+QeD8NPXN5cciEfBp4zcM
K6k+171XFoFiVW0ad99bOryuj7YJ6eJWkGoU7Sain+bYei/O0UnBekQNHiTb
xP9I9b1fpChiV6NARfaCQ9sQYY6rHCQEvCfXznWVe4IjHHf86dJoeIp41SK3
hVtGcAAFyUKgHjlOcLP2cI8OpIZnf8pd35QHuI+9t/S9PBQuLNopTous7b2d
JyUk0UjmMTlrP3yIpRugGu4JKis5jczZz0DWXST9nMLVHciOY25CC63/+avL
m8Pp2B8QdLuJGjBmC9J2XX2oLCQupMolP8VIpUcR/8R9uSVZFvmn94N6J5iZ
gsBIpPOD9mMVH3d2r3nGSt+3lJ/1xn6o7o4t0VBjcIOoLC1e24lJ7tXw83Wo
5nB4e946/WKkQH27wD1gfQy+jgpiPJGdO4ubPf8xzMdntaSLEdrOSWYAsMXd
JWDjOnNRySeBMvJJ7UMb8vLyRDZjJLZZOPgOBkIzZlwFxdWQr9PuBb8mEnFx
kF5hvzbXY8ESI3Bz7vmHjqllGixsL+yYNiGizTftckFjen9U8N2ZIhicIO3p
UiqaS03hhSiP+9o/B1WtuV3HWQKUxcTWShz3WfDR31EvTNjKMy4U2TLXNpyQ
C2XpB8E5D1WYm65KJicQnIyy0xdCmmQnROuU4XMpT6Y5djxLvB7zWEQm5t68
8cOynAR75w/DpZJnJ7AXxD8xG6SQlM299ClLDCQw3swq6Lnhxa8jsmnO3e7a
8jK6aCTaAaKMQOexeccG5n9Hb0FVVJHxcXqxsCTLflhHAvYjh+c9y833923P
bMZihs0YrPti2DBWkX/2RnUZQnbD+ygSFbwKkHQjkVKt0jTcF7YvjZa9fwPH
1E5+sQYwhEJBJAuxzMxqXY6kB7puZEcG0kdIxkJu5wRIEsVzu8jlv7Qvaege
jfs8ZMdLcx6ieUCW4wCCInXyiM6bZZEN3nomFW6QDNAnUE/L4bz/MAK0mPb+
3/dfDa9HazsVjFclOWxHUTLh9ZQ1YEvNBAI32QgW2HB0+RPyC6u08sf0F4YW
Gy3k62sh0Iv/Larvb2Nxf/X0nUxQitbAOOflRFHfNKuD0MRTleQd6Pa2gzcZ
2gAv91nsLyqQJuFJ4378wF4dyGNBdVZBKYHso9K+kEzKSXnhBpLR

`pragma protect end_protected
