// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
GfTvyKSHN1xApsAzm4wpJFW4M+OpucnWeM4kplNylOOmFyEfCf+L5v6tLae10qnw
ME4is0TlNO2pkvDwZqIeJjCRb4H41z4/L0utSSDcAgU10r90wfcm1UHm2w/hgDGY
DTki7RVuWdTDVSZ+vQ7B9koJXpNzfI0e+feC0slFEHU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 81456 )
`pragma protect data_block
T8emsR6RFNJ7av09Mr/VDv7XeykR3gHSzMKBM9ynolg6Y+f7jz7WZDFUP5DFEYoT
mB2MFzQU7EzqUGcoyyqNzCs2IPVg3GNNTn5U9UoDScIP38ZbO0QVEhE2VFA5QcI7
WLCzO+QOkuhFmkpplnWW3g8WJXnbnTp0ChK6/AAY/pHySJjq9dy/vKItdT9U3/8U
wBvdSS0xF6aFyBuEJRNuG9wjXY3fzOL+am540cVJ0riVhvzJ8POIfkniDgnpnYZP
k6RTODi8OLA+jO4qS0Ntec9gst5uPLhOhyNoV0Dww0Ems7GRzRQPNkvLi8jm5L13
BZ7vddHWDCHfpJX1CE1u5dOlrAojfpYcVJEMKGpchDeP6cFd3hgMRUNCfPy+J7fa
FSYikzBrv9qNDbT8q1wD8PZWI/+SANRY/iFr2OBgrxcGsSAFCHueA8XoKxf0zrF/
Oe3cOb7qxKQQcmx038q15n3k/HBOszGECS4wZABWKCAZnv0l/hj6fpp6+w0nIzuM
/aL5O8CDqepCC4tc2Sz9YQs19QFNVuYBA3trykYzRGnhlVWkIt5o949SjvG1wOFk
A/kwP+3Msr6Rnq6TkcUvMBn9v36H35Bmw292B9WiXKTc4krEGpTGlWD/WavG4t5y
vRkx2sI4mOseRhgVgq2Z1hKRompGVgaB0DgLNaLw31dHph6Bz/enGh1bqywLvmui
KInfBN46lBuwx9yifPHwtE+UWBDHck17+uxbdxJj2TYtYGeZnAUBEbyALKm1fIz5
TYsIF0aoSv57fwAIzVOHaLD/Es9+sg7STpXgcqr4+uHjvBRPHA9XaTZYii1O7m6s
FVaKGVqsmnl/QhxrA3V0ZLwEsnyx2z8kx4qgB0RYZaho2kZIwrsva0w5i3tQHZVB
YoFSQ+WOpZploMuYzjjiRcjK8CylvuoG+rqR+4bMmQPFSANGvqM18XgNGm6sayJj
1Mv3ufZ+3DnUudh49TElzFb8VtINAAaatbBzcXGphh87tX22nrSxWv73Bmn4TS4I
fsh9ZGrBZQ7bTjFXK/mNlYbkcIe2SdofIpGD5t/fU2KXSQY5UKtNSxMHaWleQ2be
Sf5mqphjuVcdnpOHuEh3wH2GSlIm+u0VzW+w+VDe+UkwwTru/UkgXg9y3bHElUU2
Mod4QS5eINNB9qGdYz+a4KZdYSpWx6Mn9WA7H4CfG+QAK17iQmjFhX8BHDIdvV5Q
BmDXF6eoQL06VHHA2quNSPuPdlnyawui6US1OtE5OvgZWT2U8wwUadnuQZfxF3lA
e4yf7hC42IY2Kq7VlhcUupG8faYrKShtOKNBaifYCMXtVZN7ZJIJrdRVhV9rlbGY
Z0l158aPob4vnksXe3N9c4TiFqcQlNZBa2IkMEmAOsN4oVM38vCSGZCOc4JHAt5g
XOkIdswmTB5eOeLbR31Ulsqt77ZBG3AKntbAi/4Uo2nmBtlU/W9h4dQLTRK4AGYF
vacS23qKeVSMf67kDny8QGZcrRG30fwUlAV+dSBgBJxDaTUJdSIjVWumUtQFtf+4
NZH5MfAWltXU9sZfvdAnRUjSPBXyXNVQPR7zxdV4e++FTW+LJItkrDmm0hmvJeAA
2S/TLnWNotStwhW/6BJOTHLdv2f+AXmzVef+j8RQVSrRbLaL51zzOVcuUzdq3/xF
JTmhCo/Z6tQmhD9nF5lQ3jSuhVSdDkIrpcG7ekztYYQUCKmjz5s0B/4ohAZcjGUN
tMuM0Nm+tdVO6lAsjJYaSEVcDkScLtgwWA628p0cXE73YbHqHO9YuClxxeBf86qY
QzZrTUnD3y0iVdvooHKHPKY32wYttcOI23vDoT4lvaW7CQr8EkUaoi9YClMCfZW0
Y7Dn68oeLtkotKlauWjB5uVZ3f+p7bdpWqzJnlXSi6eEQm4bn51b1pZR2f7/NYb1
3i2JLRehUlxN7zHgc+nCdkdyFHFiLXoH/xz0TNgaBFlYizk8bs58XDvKTNA3CXFH
hDjsSat3qyagdfBgkfUXsAYLaeu60NXqGyUPYASnMIxX/1dUlX3gv/fb6A+90sxi
y3ePKsbeTyDvDYP5QebrU9fqlOOEgAwSwDucz5cLtKfK6iJ7B+3i4Y7ddgIBCU56
k/6DxEWVkTegLxtl/oRm0M/rokuFH3y8INdqRrPC7KUFHZUfLUWArFye+FvXw+EO
JCKM2032AyeRjthp8Jyr+EuKA8pKI7Axw0GqjduB5iFV3gcdva+LIyrbDCuZJfQm
tUHKZCJDmzv2I23JH7HFCBfmaw4aQkz9i3CGCbvg5MV9jitzpYvhN2f2aBlMxnVg
a4dL5KcKpb1/v2qvIbsADReSSIz2uc5i2Z0zmHZO2ZcXQ4lAy1gRhXcl/jpIw168
cdOCWjiyZK/H5OI6tbAEPTEE31SBYVBr/pChX9jovvUsVfCLN1PXAPFu/zMeWKlx
crjkGdiPfX/GTS5ZlBrlqbCvhYIl1LkhQ127xUD6c1+optzwvTzPXtqGhznsmC2T
eBBcBBrcyKZopevLdTZuTI6YtfOkLtOsTdgshnAUyXHu7Do6IDIwjxypdKNZMJ9f
9Jrl2HogfDrL1lnBRYc9sqZg0PsfVTZyR01kvUE9bOyd1NdNNejwkVhYTcWkP5QC
4pyoSrORFGV34+3q+FBY34UHAoXxy/d4y96foUYByVGT8CkHoMHMF12T+zCBlMFO
z0nRMEz9y9GKIMD2+WOuVyDhOZYNkbchCOzyxhCMLmSe2mM9iZpbcjUy2TTppKuX
rhjwF1PusD5Cq5EPYvLNFpt+g/p4g/I/MpkvrYARUNPR7yFHzshFwrqZ0qNn79vK
gPSfEVGYiktHQUrV3fXhUTnjrNgo5ssgNMm3DuZoaBDAqcllc1NAu6P4FS2B5AZN
IFZ8BBz6Md8rj7AT6sOADiZu5lNFJAcwP2gQ6eeR6E4Qeh6FvdKWjxZtZ4feQHqq
4t/8hFiacqCjXUranBPp02tjKVE4jr71nTTXDX1ER+bb4DWBDWHdezVQ/W001MwV
SBUesMgOh+k/90GtHxwrbHUYia/AYC2AF6oU4mwcrVzMZIyRzVWBdZL7Cwh4VwFK
89MeXwudegtOtfL4BEGcncs1CEkDHWLWJJeK/5yH0aFVEwBStcjBl2j7a1FlYfVr
T5QuVCge7Fq4KUOH1IZgvlSMDADfBD49clHHZtG1SkFz7CpyR1h5TfluXu6hUlv1
krbf42KkuVB8NoPu7PdhsM2iYef0wP7qoewRHNtVK+qwaQ0/bx4Eq+DsXD4QJJGk
l2nSVb7hPwh2wLhYX+HYqayezjBMc2InVM9vLQxN1NAtBtBQY+DGQR1adgFA+UJO
BkeZ8g0PRP1TsY4ZoXdGkcHBWrcijKNB8KTlH2SSPBjK9rJA9s/3wzowhMamv1Kp
Lx2O+edw96EelVvRu+C8CsAQ2G7/tkq3p+uLC+D+ZBzbTwaqzAzwpqyhqmca/2mT
7t/FsQjczVb80j60YI9ApBqMH0SFhvvp3ZK9Cn/p/1OthXGdheRSsbm/wmru3H+7
oPa+3439FQb+xwSh2BSIPqcaQbH6vrBBc86WwJlbB5Bd/AWyYg1bkyg09nDVtrJB
1CK2h+Nr6ZzzoErg9q/maW3eIzkBE2v+n9WWAhxWsg1F4Q2KWF4OQvdWXp902WAv
m9Ru7DVAvC69gs+fJor+iW5A2peILJhtaBae024yuNFEmTgucCjy4JtnUlTUSZCI
cE1HuKNtffA9h3M/gImTj2pY/xaCa5FPddyI6QNENYXbkSl+VbWY9Gsxur7ohKsp
mxB1dfI5oH1KImZ1UC6IEPXCqdn8P/7Ap/Y6nGlNOBMbpUCDYpnw7LVCTUmZofy9
Yal52ecyiAxW+O+UsUQTO5+a8QQgpSp4WHQ66cCqlE8NwbjEmonrzvPnWL+NPFvr
q7HGRriNCemsIybbct1X5nkWlMO1D7ZzjOT3F2K05/pqNEs/bB7PsaZihksffHwg
yPqHnkSk8s79zI+1wWBnlfBMb6ywnM+jyqv99aYCZh5rXpeX69jf7VKUEuXfPnM/
Gc5zqpPQouSDf9vOv9SEG6/6CGHtcA0wswV8WAIAYnHv9Zzdydkp4BxOKNKjeg2+
I4ESD0DCeEct5BBThFxZ+gUao+dhe0fyKyq+c6f6QK6v0RKnsMI7Xff29gkITYiF
nHjCBGIRZCkJv8JjFDMKC1BLox+w8dc+KKnSpTRBROl9BU8WCnQnvMIvBNT6qUxI
rzn5lWknS23pW0I9JDBRGP+k8k+5ir/jVn/NmVPLcm8ULmnkhoTDeb77V646kcIC
b5R8ypQFHplX72iY2+hJpEWUs6aLF6dgG2xNaFr2fR8IGJlDvwdLe7+RsyMeF3Yr
q0QnN3lC9eQBTPLPgE6bMFyI8xwbphgm+IwNlV7fyS7crn+90bzUDAP9poO2/us7
Clrq6LlxW6rirosbyNQv27VJAoYu5621g6+hSD1EOaUD1eKzcVmgTW2FbQGy8wlU
QJ+Vo0d/D964tXrO7nudy4JoqtvQQ58plRBa8OIGiIY7mv1DkfOKygH9VfLpqTJR
y/eF9km1SpUw4NT62RQlbflL4TxFac+oNxKN+aGIME+AXOft92z8CgYlquJmLSRg
YqIAdVPg65qEa0HgVWqXIvKvIbxcGdzyiineLUM4QilRyZmjbZ/22lpjBpxbeaLM
tAfcghPrZ/vsnWGJUl4dYZ4svbzUkmV5jhWL05CVAbzq4IsgOJlh6CMLslyUJz8M
qJcuDidkEHjcO9IEG5xnU9fRWpIicyavEdkeDTEYl9XLLGhUre59RGqCdtw+gA4m
ebt+4MxSBo/Tna3kar+yd9/ngde6DXXatHxI5L8ze3iy8Cvp8wLLfot5z1BDeqm6
RkpBpYuqH7CfBOKJ4OJwf0DIfvrGQSyZAS0/MVX2TQGJAIDQYkQ6X4jL/smuQyA9
cpqVWhQfoTFPZXQBnbLxRiCZ8bqxpx/y7wceBdlHB8GtW8RkPNn44vG8zhWrieFw
1Q+MlfPrYdBjlVuiQER0j9xeeRQiwuY/+Bck8jpH0mttFrhFGRUxo/UuSQwsfBhm
/FI1UfH9cGpKm+g4eM7Znlx5VPUJi6gcQV2+yvjoT5TwiIPhWyWRVWSpKPiCVykw
Jm6zPxKnD6z7iVzQ7uBpqO/cn6+x8E+lSKdzka35WXhbUCv3ywnRgRpvkxkM6Ico
TXHif4o8pemCOFiMs/zgCj/7v6idvXktw0BksCBARHYxyCvOy+yKmi6G3I7nTOeK
iuLy/aJbY9HKqfaxlbGnHkrBnU82Ltcuo9dC5NR874lglidj4DlQ/jme4FvGsqjn
ViuRWGc/zkjqmzeep10pFi5NGzltM29NH9OjdZqv0KSlb/1Ibg1yr5NbWVt8Vn8E
XPkLgAmWHII0bphpbPSiDvY40UEOI0pKcyPBragtlsHF6ixMf60FE6d30YayEvwX
Jib/Xgr64UiVpxiPc4S2Yef6nmK3vztwFlAfLehtC+88fhnA4qvHaSfVwjgjTsKv
7ZcNLJGMpBnQEkcKzc/MLxhn3NiDM1sSCxPni8ZrHyGo4Ydm1ij8+EhNggZOvLwb
tWJvoAkSMNk4G5UhUpkD33cNgnV9xQ4+MWdt0iLrvKlraxn18Uou0m/NdsYFAU7T
wjXVBwO9xvTJaH/Qtd9S/pNcT2soMJqGY2CrG6aews3Eq8rvvkMFkeT4ORUnqsYK
RDZ8wIGmZYx1CBQFo9nkYcc7NVz05Am269zsxVYOGrUu3G9bB9EebeBx2BM10hB+
O8qy7s9+zNerZyL22FOGYDM9MtBfNm/pctQkDcFKJhJL7G91oi5N0U9TziN0ZWHE
LKRtMKmSI64FZTPwczm74suIr8zfvGSI6tD3lQmZ7N/sqA1vggAeWgTdSAEgFhHe
OCZ7MCNXKpXP19b4QCH5ylFtITt9SBWT2i857odoLaWhYDvS6iKlNPs032CeCZ3e
s3/8IidCUA+iUH8KL9YmvtYbqJIFUgbfcEipx2ZfR+KnBDtrYFTEGCoI88Jft/eZ
2d4LkUo4fbq1tns0nDdEfRN0QwU5dCOMhK83dKRSlcYjO7OuKD3RqAQ7dSWUU4T4
YObsK8HSp/GG6vx+8KiLuVhqv6x1K/DV8kYWc+U2QObhHCMCSp4+uhoXuDbEoUvR
Sl6Okdq3Ct/N2cQwvcS3Lc2ldhnvaRe4PuBIQXyARUwfi5MdxkeiAooeqKvGkhRK
NrAPqGC6Z6TPbUocTTKHk1AZ8ODSXBp1uYi0l92XOXYaccXwY48XW2hY6pOXBbpG
ONQkJ2i/rcfY/NJCAoLPfX5bh7OmXzL1Vjup3PDf8oopC4XPp06UqEb/mCloEtVf
mVC/R9OrLoebV4KM/xewDUUfYyLkN701+UeSe8xgu1TkqdDfPlMllQJilNno8yRu
jT8u4AvHj2jTVnsLaG1RTOB+00kXH4ThVcuH8DmRmbTwCLcNSqO3I9G8t9n+Dir3
zWMq9CJj2fTjWf1u8k0odCMIJJUC7uNVTG310E0ug6AU1QD7Ub7HZK/GXJwaoBJl
XbPQZmz59hZFRM01wQU/VArudn0QdUmcbtEx+8rIueA7/vVZuuGcXgE5xqUg7GMg
auCvUjGN3tFIFcBJ/xJbsRl2Rd0ACl/YGSFaoHZ2TI2O8o9MjUpWoXOXHf/YZHOl
LhuSM/AZRFll6vpDNgZTjw5n4vtxEUkg4KsMwb/iR/c8Jej8kIqqcRP6tDE7qC9v
PtEy3IsTcuSByuEW4sBqHGdqVZyuRv4ZLnyp/jOoX0l0xuC/t4MznI2OVxpXccgy
0T8bzqDpkRs72jq+bpMMSMDzw6z3GkQqJzuIV7QDiOqnlPUa8nUZw4oXeQMpYMoD
suoFIWym6c//y+8VCQz3d5JYHq8r3o5QBrx5RnJA+PqKoXlu7XbtfHBOYsNsXg9q
sysro2DFLWjbDOVMPiIbJOR5NaZCzDym6SBhE1T5vLG9OBN3t4OT9JqDnWW/Om9X
od8KHygeUapj8RZ0mUz+nbucvhxUVHUayB2z2VbsVxBgIslJ/fTPn27iGnCb4/4+
Avsb6WZuqqVcfRnmPmwVF+5GNY7cJmsK38yLY3Q5OmPjU+9zKZAimNu0wAeRtP1z
QX6B4h8DCb4xHgeCdX+pHiwhbBlvX6dkdC66GUaGj2N/H9WH5HTBr0xZgvTkWqB/
RdurJwykZFUWZNUuiZ4KYm8j8Sn8ihXJylnpsj5tbaskMVX6Vu0a0tdFffhoBmUE
JX8enkvntFAte00BZifym5yJoPzfH1p9ZvWFmTqNqP6i5ZUO8+ytwkIb2YHVnMyz
mYkYif/985NYRZ5zL1Tm6ZZc0YggoH7JYiUeU1F0JIaJIH+jXf8/4+64VvfEa5NT
Ezpm1aRpjaeUKbCYQ2PyDkzO2fmiVh9SfBdrHeKmbUonTFsVr4dilFLiOITlrosX
C7z051VsbfYOH7npB47a4dwI3oAfPfRezQlWyPbKK0G5eg7MmO5glyFFhxK7YbEC
yCAfum7Du0ulrqrUnIWKmcuWHC+p57NMy0nyL3mLOEjJee0/vGldceLPkdSroBTe
6/HIhmmv0Sb3OXGnaJZrXb7oQ+rpKYeTGves7OB7OdwrhUtGbo2WwwVszuZmbnR2
7NhSO3v4ZUoeFdh8PmQ9Ba4jpXPOE19AnNzMl4EV1Mpp8Rzt9pWLMvAADwkfOUa4
fmnOEoKIjQx9av66dpnCKik3qLG3TMz91yRNJpciibVkWPheCLM+sgQX77XBGoyU
CU3YP7kcrtVB4Z22k87yNeJaWkeK6CBd+pMc5PnG8Bu/ivTfAEbNIMX8eYV1AeYf
1bvJ/3rqki9EdiFpup4156D9rM7/6TY0VWuyVHZML0fL2hIMHWzagNFO2GvSpUd6
N9ZdiunhTaaihJXQJ5XiXAJhb0uMm+VBV4CPwi323cN06//4St/QAmu2/1ZUYNpL
f4Qk/d2H8CIy4hU7GKQI1V02qnhSlCXS7IA2fPWUqPzFmCXu6WuNTNXiuG4f9/2r
Dlrq5/O6eM0UhAoa/X4GjaxryPnuph3ZG7WFRZe0sGhZd3xw96jCY77UpY6ASUke
rxDFT8U+sO4lXJdBGarzZhSfNm2uB219AvTnqtFKVAtP/+npAsbORUKu53WYjMZI
Ydo+lXFPhNjXuIcHvTHDScgLhqLfHsqCbfTbp4yAsy9sXU3/BvkoiEKR25kD8X0I
CKQ+ZyleduqxLJ3KXRqZJZ96rHXC25vgRI99f2UfSf1rfe6v1xhxtVJxrW4aU+wa
JOzZgCT10otXXECKs2RVN13fXgp/qLv+rP68+dNjv6yzcHXtflfpOF26E4ncAgP8
QK6f5rjYPT4/TFFtj3yQAohfwR86A6bpOvt+FeIZLSZlqefgOp7w7ViACnt9YwAa
Jn4dvpG1IhXz/sAJq28KIaxI3jzYlnDekzAjbeKywVTD9EbRKRwaxsEgzO/gqMms
8BA3SxurKWINYmNo4DNyMZRkpw0hKfO71KgH56v3jKpp021YgSGATBo6AusHBVv6
4hP4jdr5Cfi2KbxUIw2bvOxu3dsppCCgHFUPMvDBBoxD4i/0qAiL58mFAumh2e72
4xvLPcQvklbTBJS+dBA7EKGTCcEb9aqrg8psfhy4eVNlbqrENUTqLSURx/wZ9AUG
Hc/akFzUzYnWzfDMcK0yiTADqYgjQdqYAsm2j4kG0TVehiYGUZtd2K1BBsQPEm0d
oTTYARwnhGKxAHeUC7JVQTAil2UUJAIbp5msAKFnMYq1nS46AvxN4VQlcnc2ehj/
qUyY57cnV7ndFL0h2UGIWkdz6LoOM5HHkf7dYfAXlZzKtuithS8j0nSj6uPOzpu+
K1uNz236kkiqmQHnTCGjt8yjAPbEbWPFT/G0l2CTX8P0MTiTaI4F2D/VXcvKToyw
LnNqje9HAKylbnT+/mJ09mXT65B0LbnDB1Ec/H1V/wuAwqBSYSsDI5z1ABSVwm+B
qeZUy6EDZ8TJ4oGU2B671+Ww75DWrBEJ6Ytkeai3VT+zcApBUVO0DSVDA0wKsDBu
0zWaL6zBD6zORp1doKyRat9gofSni7j3NI0FCdY7pPlYRYzQrqbgpLUAzP+QCc+l
3QAS4ARTERxZG2YdeeZ+XbmfwLMPDL3nioeodltKBXnbV0/TUX91406eH4vHtWDB
cwSm82Zpr00sMC615RIVL6P+Y4UU0pb1VD9YQk6gCsi5YYNbgNlkUfsLz6EQ7s21
Qlcu7dWoKABOK7en5nGcpwifBHRMxgJ35ZiepaoLVjU2FpvFSt82OsVZijj6pXip
o46JL9u3dUSZf7UBKx0xgxy0foZYiKwnIIPPipfiJ+Ht3M+sT2/zJWgx71ii7Efa
FGbU0+dP/dfEJxKe3Ey7VjrAq77H0WSIBvyJT8496bCtiFrEUOyjfv++FYs0BuHh
MOkr03wccrSnv7dT7qZV7yj0q1uSFIrqIPCMbNeKENRrPgHTVR/UAU4TTVL90YI7
o6+Dc49TPBiCoB5VJvi1Sk+lXQkqMe48PkxaqUt0+CjhTH+0GHkd7WIS2/OkHLUv
fHDgZTvAtKHfSXkUPF5+cBx78dMadCmDPbRPeJqJxAML+Id6auqKdu++Kayjk0ZA
HFrLeGr9DXLePiO4KBKsb9f9Y53qTuX815ptFv/KfBx4ohfICWEVOjAYVTMYPcpu
LuP7fxWe2jZL4/Sjv5jo+n96gPQk7aNcfzZMQNDxISMsLEiMnZ7nQWUXr24Gapsq
HN+ieN8RBorfDu2SAEqtkN8ZnOGggWXZzXuoOs1xFKoufBBulAK0fgUNfxJEllx9
SFMnWi55SiWUuNF9HBoh3VHE88HeFUzI9qbYXZmCW+OpvouhC6CcQJpNph00C8tB
ena4RlrvGXXeZdxX2EEM5uV59USwFpIzw6+qYvWFglD0EdZOgoqiTO+tnoHNsyx+
s4NHD7ihcUWiTG7Qm17X5vSa1IDmu6gK0ffQFWnyRSEVSJGpb4IEJtqtHtjrCwEe
LqnxCHXlCtXyX26wH5zbFpwIoH7WnJVslfDk36+Ad8MdXz2sOekk2DnwMLq9Anpq
gQAa4DNAixtUKoXO2l5UFS2omiybrLktkUJrR6mlStReN9YE3LaoI4cOmxRacsM7
py5B8b5SEUxVXMDycno1gk3kcNA7lRxEhbLdnV4H77/rDrMMzN1RfLiLCeNIuyTI
F1V/k42gWy4kdZ+NroqcYotHVAhGlxJvN1uU1r6cBilxcklCASm8Djk2N9W+RsbR
LvRMXdbAZBX1ATUyPrnCkXJ+whEZaEYdPeOoJ3tDzjG3tG0AJjzC37HtlP43oY5D
QxCwQtG+Z//cVCRJrE8mwzrwkDV1SSNg2QDM9fSrtL4BKMfImgUvL01XEhGWsDr7
/m0h9TSxp9SLLGey2pH3dcJ4VfTG2a0czvKZvPXUjewMF4pAYJd/JrhKscA2oGc3
IveFuDEC+MbEihKmRkPp3UMkTj4JwYiVM5lV4LFsJxQswkHLCCmoMbfI18ij/M4k
twWS0TJEiAYTHMivMhNc9/k3iVmmSXLbCeNU/uGKXQjpB05kTqSpekXPHRRcIhc+
yUMRTX+ZWMM6GPPqDqJYNIUvEUP9ePyI0nLSBEkz87l364XJLQLtqNkSQ6bY0uGE
7vmrwAXT5agim2oehaP56oO/0GY5qrqIVAOWQdFcLjwWA141E20DEYODddA/lOVV
rknwBS/7ppaZKr06RCJiqNxS25toedi0cu+GIgQhZwz5ADIIdbofDWLZI6SXN5oL
U4++Ke3nK2t7E5Jtrkdcl3LPjd9pIJJqV5HWAw5g389vR/K+m06QTHldM0c/4LOB
4sQOX0mr4l80QO57bptuHwX9cV9fPWHIIG3MbWaOxSNRqQ4kS8vEuamaP0g5urvZ
zxj2KadlmsCMLL1ptGQN4+2yqRCKEDsrFxooNCxXqSwihfEfepNdp5Ncd/NISr1j
fR4nx7Q4fJoPkneG+CYW6jdG3+o4rq2u0YAg84N3NV4AQRhZniKUzhhYNJ27OK1I
Dy4n5OKyIUa+t5u8smDyWB2qfN0AUCrYATR3srt7uMbKTJdzP/aC+r8pUPjRtaHM
BLYYMckFeN+St1X9lfDBiIxZsnFKdwKmxgAcfrM9r1ul/GcJnNK8VB8Ga89WVKte
OBuDQnbCkP7z2kYmfXeJxs51iBOZfTCJ9DDcXmBCjn3sY/rSMDe1jH5d/yQlPO2m
xiZfyOInYG1J0KTi45zD03Dz8hYPEcCh+uzNrBEmvU99FAUxr2dGM5BXfQa/15hO
ErZTtHamG4Cj8frLpHvtrTvhBciPiB/oDb1tdJNnIF1cKep5iRKWKIbg1DcJjnd9
8uR5oH3ONSqbLNCAQBtqq/Tg5ByRg2Yg194zvwjbdnO5yiNIy5S6hKq3RfiDQHdB
Soahh/QpXq6/d6PZ3WGgZhZfYFfzhaNHnJYOZTAqIek+TYd5qc784TUE1UADCwjd
B+NdQ8XZE330374rGYR4xGySuvplbdcgrWNK/he6M2Yk3G6TVKoqFJThTCH5Hu+Q
3uMIz4YZfXXyVeMSFIe8NGcURZMchIYu2RUd1fOhvIR5GGgeqB2H3phhiWDQO9eF
jQzZwvQp2QqUcITUSw1oQnJSUNiCYszbTiOOAwKqDIRNTGV0fnI+dRX9CIbFupWw
2ZMFTWNFgL1SBbJ5Qy8hkUgzEboGFFc0FKPFFLij1PGv7zsJRCmkklk8ZKzJeAW9
lggXf9tC3dCMFxu7x6pSsMaASjTVPLByhvDhPwvEMNizUO+yAcFkHQCA97CVJfa9
GdScF2q3sfv9HycLJGVTsV1uN8A8qIyTerJzP8sqNKRwPkWUZgRQsgzPbsXhoSc8
Seyn4iIJhm2M9laXbVinxCdiQBfYxUQ2fMUQAWen7J89rD68CRDRJA3fzILNFPwr
d1ZQuK2bBjVyGF3Ad+phkF6EzOWCSfXCpDT0pDu+YvLB3CM279U4X+x87/H3QnoL
t/TSQ/uh5hVtFepAlr/SxmXMQPQjjATyCsI1fElXA3+uzHsjK4SqVwMobR17+h57
CwjR8CJRtOC5tXMWYzKIrOOTTaH7gji0J9tYV42r/kezPZ9IRp+jvGayA86ro9SO
PYf7jmcJucfb6KQSISfqb0e6Y5TMjfPoOyM7vqjBiRFt+Wjb2CCuks67CdgAxswD
nLeEWOtCDzvmokYJ4W6bbIaGnZcInuoBxR9TZ2H6XqeMdrOEdjzFm7imOPEuFuJx
EelYtrg07GpR9EZ09PHDk2XUsF7Ozc5aJG7HSqb3XJwQhNJTnblnbk+LClR5GiiV
tkald+X606N+2wvdf6Mq5tICUD+yOZVLn3kNaVWx05eiOZas4SzAv7URNTgjHkPA
zqGDsk6A8H6p8v3jk38C27ZdWYneiBCfC+0g5P7sRfkng40SKpQg4EJubb/TUd5s
ajW3vvN0G2ChVlqJchemelKZ2IXwO+fB6Fq7TIiaWAjcF1p50tgyUjRrVDcH8C/2
okm1U6qTHu13whoN5hbZfCYqAN699kBtjqe64nC4s/Y9M92hlLTx1Pbdc13OOs6z
QvV6Fc3H+Kzs40QBaBh8F9COwtXFwcS9Z1FRn006+KYScw+3PNaM1F54A4sDO6HX
pIemTvBZpMwiTPUW3MDz1P7Tm7gvdp78BMRvudV9KRNPPLvtsQiMZ4DiJxtSkxXE
V17+6QeFu5cSENnpQe/IImNwFNFbBd7IyLmgHgdT9g65pOl8a4C9o2z6CCdnMKMh
WO+DF448CVfs7sfdnwSEIZBsNvFay6xbSi2sHUGJdiq+2oVNDbSYiz8Ojxwr7J9i
bIeEw+G2/ddONNuDt7IYmmip7uw1ca2ujWvnhAttv//JlW8bjaxtESRgw66Ubb89
y5+Hr2iOHlyrkPUTIfC6r+gBcUT5I7kPw1ivfYl4GS2Ee2KD2IzowTv7iSDtxxTe
Az4zfbZU9I0S1ImHtLA3MlaNW8b+mWGrvi3MZh62rS4mn4p7JNsXZKHkQGZBkwLd
viHdzSiVV2cu3C9AmfGtvdkd7qiUzOUMtdHLY4OoNrRAr4rF+pzDHrPGWHb73TEm
px8JymlB+rZPusAso0gI3eQqGZ3HwGkokVe0BuDj8AL9dRVLUOBcPEl1xai37Z9g
VmcFONuo86HbUPNTYOf6cSaGexiZGwU9aP2FyN/PbFcKZ5i7hyItDU9JCOO0DY54
PiSmhNj/76pDMFx1uNiduN0dsREDfIGrYOByBxZ9oZDZK5h4sAuGCY6jhAioIvhj
I3QQ4vAVurYZ361DMwieU0NUVeauoPuQ/IOTxVMF+4NJs3U827hLPTQT0Ry+lPCM
Fjq3EbPEbgxCslMTA58A+3j0B5YaRVB5r3wQbPK6iOEd0axklmb/JZ38YUUmrn/f
tXUorOFisFQ2Qj+NT5xKyofRWMzYIM1ozR8I3zL9UZNwrHUQCotKaow7u+L99MyD
F0LUKFLGCfQiykujR3+8jQrs5RkEruYkxj4SMw/nOz/SlGSb+c6sbK5Dk3+/WvNK
qZLfd4KjSyWzraotjJmOolyyHudfYwGoy5yQv+TAnIlLjnf1xXg39h9jEKENRn/J
0qs2qFudCZ7kwpvHWrwrk6THqGMLJT90pFX7NuavMDqdjhn6zkXIx8R2BksejH2h
3Ua56dREW6TG4SKdtZhigNQV8XoM4qetY8CBcXWc4HjMVn6MMmf9RcCnf/0LVytl
E3oeQJKlECbeb5p+QRMs8L+otZbj0+unDlpZjeVbo5YdpRdTcPO3Iyipif/07U18
UXPt8sFjRUQFcRqOx1dG3VatKKkbY/XSKxEtGK4Ktz/MDIWr47VSHZFiF8tJX920
ZPNnAVZG0CmPLwc2mUTXpf17X8NT9iMK+URPi3Cw63DtJEZTK337AchxyjbRNMr1
tEhKzH5lN7av4DxJkP+jXcL7/RU/5R4rbHWrkckAuwyVZKGptmmCgGtZC3dmlArl
yh1kW5K4S+elN50rg8af4S3Wu9JSWNvlP9r8wdyQ5KfObyMeFEJtXgyQM6T80wh6
1qU1BthW0zs0myHgdP3ZyiZzPw6MlX6/kwtox3QzNufp3kus4/cmedhy5XOYKzJ/
O3ZziPApHRLTsnrN/Ys1btm0BVgqthZaO+72fTZkM7LY+jCaQV2/GqHqbOogzJAt
Lkk/kYvJxFE1JBHyRzUxUbxMxaEAtJuFJMlwWM22zJWylJwdRwMaRuSRCCx1tKzt
90zvVM9QImfKUS+QuxL5/8Z+b5YXtJIwrSPeViDKrxb14niZ/hYNKWbrGwMtoLRT
yXP08yEsGxuGH7LNboiKkbLluedfbVWgZKa6ibd6FZOs7/PzIWqSxmXFpFEqucw+
qdqSPsVp+5tagnKRlCa3+jNcERmMDki65WbCBvxmb34rzxobdWR7/FVjA73D8cBT
0C6AdGgpCbxtyddc2c29reAWQFM1OXAg5qOANxn6h+UfRhP1KpFJfEY9eqK2lgmG
PIC7dyzim0klpPDviXAulwbNY2aSxcGdwG4jmt6j5YOAPpcal46L+mFHXJID4hyx
ANfbyTyYlEpaYqpzeNYLHPT7XGc7PAVbHpSQY/pPxcLChDUpiZdM6x+AXQ/O9ede
SPXeEaDqdypQ466olXYb08e6VmS7kVWQErCLWh3hgn+2Q0TYAd1wJZsj7M1CMB2a
ha5q91mLeL9nbj19VZWmXL2TNmSnCl0D0QEnfhXRZHjhpdNf2qdyDd5OfFx2ApB+
lpVZezAdau2myqQQIexggP70LPlMLzOsXwJk1JbOnyCWeE53jNqqAly2L00FLPvJ
AukCopg73+VDOaQzspigZ5/7Kw0Vz+q1NP/wAwE0LpUDGAD5RyYKKpzxtQA2WMD3
iDOzNp4yaeK6gZSZ56BmVCOyq9G4Bv1cna60IeBVL2208hgy/5MPqQeRVinHVKBI
7+ytyZSW52uuTASP4ZWqOgaKEuig2CRtAV08yVZO2yAL+M4nW4DSbY624DLDkrKg
25Z4h30v5yTs5QTHzWZK2yyYSqCnKRynv6zxytsUaBAZCNCKV8KyiN9Rl7J9dXPS
a13CuqSJpCMQvyp//o7xbVKgEufh6N2nfBj2Zt7RlIx/VbA6yPCkceO+IBn3fOFE
j8uNWFT90ObbSjMN7ZpF6XINzfVVd9qnwVcjbxEiM79Vo2TkW5inSXO1pLMVXUej
/2lYUMd4j3W1ajYc50VeDoT7ARDOtnU3JlSdKYew13V1qoiHqpuxA3yBcI+4IO+I
JKl26weCxoStzJSpAKHBtAXZXr79JgVJcPsowZTVJbfdYJK9osjDzmurshDaztW5
CZvIcH1PIX4mFckF/y3WFrds5P0PWQ48OiIDBTbCGUnUBCedZKdQVZ1DkUXQtqG0
QG11v74vRrOYIz4s05AX4YSRYWyOBTLLnt04Qu2G+Ddj4Go+j3d35SaZeptPCvqq
a+w9uC4tLo4aKjdsaUKx4CuED3wZBDQkOxNK3NToI3okS5Kw93wssobOxf1ORuY/
nHe6tRIazAwLga+I+xZ6/HVucYadVeE8lF/RQUhhz7cBFWMsWcenXmd1PWqFzTwq
kEDbW7BKvjQWgq7BH0WHfrtklpBBNbSMJyo4EyBk8AFYxCsNCvMMmKuyQanH+Ahq
gFxF3nJEFGdE/yQGOSaPoi5VeTs3P0ew5OmcMNEj+AXOMHLmta1ezyjBIUA5zpFa
j/Pti2qzvR4pstWADZiEODDDDqXYPW2QpggiSOvGh9KiJNKEtXQfvzBGxwaIp3kQ
yt1f/ZRx4JXARUn4aSaYlM4JYtNSG4rTt4BA+ickjw7U4hHPuAvRIJobU4czHOY2
UuCa/cjuyGa6f/AIy2iQOnRgWqOEsMLZenH2PVjHg2KNMbCFMY4D7XiKxL0iHBUi
dzX3c8igOvhmo85wWshCgSm3cgHzLE6KH39TOCdG619QZVzq3XFcefnbz9IRRDA4
FOTCjIsWRZTsKd0mbCLYdxka8GXzCExqEGUq/0VtOHuPu4vQ4VgI4WsD6lNOMHUi
9xmx5NCHPW1Use47JkJS4cjS/YiRJ/LtXyI7VgvrOyteL2Br8bKlakVPOgmEzmO+
1rt7mTxEnOt07uSVBXgbnIFoLhZzj+Xz7Nqt+FTQjZQZJOrLBpKStdaYMBBb5RvU
DsgHySY0VikUgpYksnAXKNeRq3FbHESaK29lVObmzCb1TvhPx+loWqfz9W1+Y+HO
nOdNKymN8NjnVasERLECdPDeMqAdbQjfo9yd8YOLTenFHDf6z8VgI0Xm177TQZ92
+SjClch5BdsrVNNRZz+blBPT5G3TZhgpiyMewCusAeirFMjhCyXaP9leg/MtJ4Ww
Yml6prWCXr0+bKEGFHbvFGZtnhu+92Fw+cYHiB30kdhdA35ICUURP+TQosgT0qvY
Zk5Ys3g9WpfHedzjUqx0WQEpq2dAlfR/8jxe0cUIw6Pp4AF7kdiD30tWhPYDp/WC
el9cxfCyEAEwSAUFOsWeVLTzbFpGypxOmZLJQJVCivBo5WGIc9Jf1acg3DFEPRiZ
Qr7wFqcqcyIZus4d5RdfuUoE6j5/vuFV4L3lykMrkQEWmHqNpZzoSVFc2kYEXgxj
pjdOArza8OoRVHiAq99VAqh4PDf5+/S8PKM3qaPaWaAI9ie7SyrO/lo3z2ldTTu+
R1jNz0PZe13XcyYR4/f2y04ANw/7p5+zKDJeP5R2ejiefxmQb+3nCPxVlJWwcUeh
TM063oVdzr+Y+8a3gRhQ/xnwZrh8quk2ZfQ32tTi29ibJlXKuvXtZI+hKP3+5inN
IkA0MO2a6/hlLlSDYqoVDB8WF+x3HGjId43zSXlMRUMgkgCLiP6eClJ0OoYNlSkJ
Pzs/L0zQlYLzyR4jZh+roky+ZzFwdJXmfhwLbPc4t/QMY3HKL6LFRYiTuWSGCBue
j4yQbOq7a5M+DT7U9GB6jOBVmBxwOaXlyRfT+GcHyUOpMBJEZ7X0P53L4BzRZVQi
sQpAttIZyRBWdFbLN4nLtylnT8tY+7GY7A1KnV3keUx12PL7LpaQ9Zzk9yIb45DB
YbkviUpmkXCE8H0G4I5f9Vk2DIahmIzainig/trDh7b7a2lcWnPuP00jQ8Yhw58D
ybxWtcLlacAAVIJwlxHHSoNjlhLmj1f7lncy77kvgUAazks5UNPJCN48rYji5rLi
C7ZqLmpq+H9dCMA62GtX0utBKrl4tkFGHI0jW77TYLo5tutL+TDyWbDy5HTNJ07p
WtkRHeUq33pImif0Ld0Z7hZwi+DA8LNz+qrYMxqmfw1kXW2XhE2SZcDaC6WxE2FP
Raxax1rbSq3AhcfGgEcNq6P6ZYYqbYTme/88l32z+ZSat/oBqy1qld6hLP3FQP1q
vXBuNgsIGBi1TB7Y0tTBSwNG5FllQ+BqAkxEjqYkeCaDqYCCDMVsXPmS4eSySUNL
NgIeXjt7GekLhQBe9J9mnV5EaCEIgRujwo4+7AZzRpDSzxYU3ClfWbGSMg3f52BS
0nz/kHrC8Ki4TH12HskkFZjV8BYOY11bdHP3fMafqDY6XWnpQ7IJ5ihurfJSccZx
pCZwVBBZ2ZUyIgCtAlLg7Z5y/mcG6A4cXygW4Rnsc26rRgV7guN+DmUSuQo19MBN
pKKfig+3j3l2G1G/15aI+Sm6RmpOcxTleTOb7Ab/MWv8Ecp32TO2t36u+ovVPyu3
tUPnZR51DcFRPR0vYnj07cHMXKnimVJqnucqNlplCU/uB+3URK8c5ChXgYLHFOhl
UgbmOJlolG/V4zv5FXjYELd5fQqQ6PoZNNFLYBxv7oM4AVm4KwoHSr2ioU6Qqp9P
uyGrys1PcCGnzXPZc+VE34VKaLo4PdVT2m66kAMdyaA22yrXBTH/2ilrDEJjKNs5
qg/oxfWvFh5JyrhqiMqnWNJH8yYv3pXbg/fabVQ/OtHwFvGay7G2VX8NHLYGWQSu
fa6BADwJ83eo7CqlFd3IGMrBVLujdCdvH879u4x99JA+zdTg+Xne8fxUz+EKEjxd
DZP5N+bFEsAB1BUKt8ffmSJ6BAUGXJEn7+K/g4haeibxC5JZwWv6Ak3VUypJhoFl
qprhl8zebZK+HkRsJOuRHJJal1GPSZrDSsNtNofQw2ecIgJLuogWmjKteEY8X5sI
zMUM6WpR+PF/qEHMhXn+4XNRhGFTo+ziLboj8SPEzqUn6MigKJczwxBN9Rncesvk
DA9fRYl2a7SsTrgi+Hm6tNrV++LdifBsithJGYK8CK7CouQ28vb9KvEs/cxEQl1i
WDivbNV5gQax6O7LnI9PZOjbdiS2u9yXC8SQ5wWZ031OGKaUqUFPoAi7fshvMp5J
d+O+NrAWVBVFksd5JtyRpEcIF8sypRmzU3/jCQoJTzEQ8I6BoVtxZcY62DFaAuke
Im3qgb9Bk6NnHlzpRX9DGQ3xBljsyhHWFIcQulGMiuV19fvpoEi0vo3EiAsvsFm5
wy+ZTecvsvtUlFME0uGlYuV4MR1qvc2M712Ji30ZRVkEeSgEKsz+Q9s920SsPFqg
1+xwP+I9dTNGdw/BLqmtaDvihCuHhYaszUiKXtYCaj2FxPmVfOqH/tVrPXHYJCp8
jkOh7v9tXbk8DBnoJUg8aTnBu8Vu8mAWs8mEn1msgaOc0XLHrRQBf9uGFHDQ5gfe
22yyDRTDjkpLilSsJEUJd93wQKjB51qTaCnLAnLiqwP20YmTWSYqD7uF/aeETfsJ
yVbb9STWhrWagAbkzrGisJG8RxYdbBYEGEXhBS+yKsS9wkqy/Yp4W7KcI+nJPxlA
lFJ/cUnUH2FQZKZcpLksCAaAE6ZeM4k4IhHvGr5EXRkxWQxcpNaCLzKRF5jDUghE
H0gGu3B0+k7EZ0YAKJNcSxTFTZbTE+UR7u/hRQurlse6/6AFspWmKaEkVk3vNVx4
N83Bx0EeqboFj7Tmqnrl0cf8WaM1rEO4VivNADleXuOvFD1SShc/nItHU/IU2qhC
mIntzFXiWZgWDAgZeHnUrMCO4pv9mShqMsRK2gzeOeTqGDMyQynjejtJKIker4Za
7D7J2KcDnJS7lBlZE5T3QQXJbR4EJYk6KA8CERz6GOUuTJcCYc/CHs1DSAl6jwXT
cuk2+wLKqjAaTvWolAEvM01aoaekBoONLP/XyVqGqmfwTSs9QEVggOT/6xbWhtKH
ijQrUbIHMwYEZ7ZdkOhUf8Eg4WGryOMvOOpRVbPo27kisZUdPtujKYzk/aE5udyp
M9QZo1Ee3AMvzDUBnaAt6ND7SJ5gaFkh1BaPC1Mez9/IydpBshIZ0pyMn8452PlQ
IraT+f41Ywh4V1P8qVjIiOBSvKLTvaW3LI2B/QcF7UJ2HhUZELo00Is8Qxuq/RLs
mPyv4W0/k7voD86FBQdG+UTj5SQUsvwKJDlKVH9eSjYZxK5Ip7FKR+YR4FwKigCL
jiIHv1kTcH2FagvQXEBuE5eZsq80QBCXCPf/c8/TqvB0z+JmLgt6OmhC7xaCXqrc
8/KKbzw3bZUfH6ZR6WB8bCELUN9mTi4DrMSdYECrqSMh16IqYJVaBmunjpSY1msu
63fDf9g7c8+J+Ifsyef0gFgXZA50pP04zpWpdG0xcHrHru2EQs88oxJWyIg14Eco
apbFJrkF0FOwgC1rvjgm4FIEbf4G+3iB+AU+/tl+ToRcb0eUNyDlNGpzWIwAc+44
WoBZkecMd7fX3ffi0IM+yleYczw2LJ756Kc96w+xRp9YYwtSCPQ4l13MrYfmytLt
41KMtqxAOwZfzM/WosNnoFLCHggb9I1JtJQpG6ibY+F6tgwZJcRw3F/0Ng0Q9E1v
ORB6X28w+VNQ9WqqJ2VEz99ZGWX9LwoqYEqh2DxcVYoOWtg0K9h5Oo0bJjefGt3J
ISODhSpI1MnQr6CzGLPEfntuypkXLDJe8mQeqndA7agUNstV/tMd5BqWsFWQZ9HT
/32eEAnekCtyxCV7QleZDrThYeOKH0pZEOPhwHzQG1y7dRCRsQqfo//v4VYnRZZy
Mwv9DSMIeFRs55XeQk2tih8LgMop8vOXPzi7IgUyrceikQAkQOL0V5PoGAvFlnky
yUUn8PSXdEqfI4UySmNLd3tbrJVI2IUIW7g2iH07tb7vKF/kx1ZhvvsBey+d/C26
0yA8q6sl0vZv2F3FmdcfTlYdk9NXvfCE4BzWIIWgqA1oyB4DWBc98Yq4gLC+EuRO
CInXV7So/JAEXw15zA1avUntHJRV3kkYOInIy63ZMTRaNEcTiL2su1m/LKBrsWNg
PVh/kOiCzk2uu3WDOxJW1Hs5+v6Th39BA/l56s0tE0MoUY/7ZZFJTq+SwjADVwPt
sFwQ7BSq0CPzLYV+39AJBgkkN0WmI0Oy1SIftBb0kQa+uI3vlGG2lflew+ZZN4gZ
zOhcA0Ed1CCc0NJ4uAMEXGX+NIfItMVZgyoI34zU4NCcXQFQoTWo/yJxY5tbQEKI
2hvTR/ARMzY980IZBvgL9nFDe8hi8zQTn0CW60B7kn8x89fSIIBPV5yifPiX28+S
5nxOX0TA3CLHHYFBXvyiTd+gm+tDvuGIk3N8E6pl1n8dkDmBLqBgaD50iUhD4Eqb
TEdyF/ktFVfAxkJoouFMg84Wrg+1rDInMlRuvn81QL+7/Kg/fzsrDjxAVGvV4IZL
BRy5LGRGHebsR3+y1k9V8b6ckTHpPIoWl38veqIFBkRE0TooAIwZ7WYeMhW83OwM
kc8T4+RaTHEdALaQ/v5WxotjUaxeJRTumhE9K7zjFGpHt5JirzvbrwwXADXnb6y7
eB2lxpasR60+Z4G2rfMU1fKw3lCMKKU9DfwSK/Z5e+r0sFeaDOhakH9wgmDs5Afg
T3kxjJjdpNKmAMFfvvF795D8z3p7/h8trWZJAOPLmExaHDoobQYVqZQnFfFnQlcS
1FejOWdnPuY7gwdLPlIohxA3dHPRau9G45RbK4qx/z15xNC1Pz017LK6jmbCNPLe
wNXWKQK+m7edYnI1GZc/2neOlzmpCX8hYlBJvh7TyskflfAHoNOJuOY3Q5oJQT8t
M7v2/ipru7BHM1aZVqD84clCZE/fOC17BlVzNUvFaAnsl4QDPziPfFycSbdDosV2
QldoAs7orBlkvU9dArhj+X3gP+jJTIaeIGbkgx5WLWB8RLeFcMmUn6RviPCuNsNQ
szS5ObNbeddsp6wVplpzPNPyLdARRaupbaeM+AsbYVt8Ma4/8INhVfc8ofvuCGsS
kN4bA0HgKEqpbDok+P8JhXGPE1nlAsVieZBF3SGgmmM5q9Xa5ZCK9uqQKeO/99pK
1AU+soPuFQ6AD+FVtT2lU+LRwq40dWUqqBet/1viLjQdob+aX5oYUEHC5ASXX6Kt
qRVOL1VDnxhNemspYVLaOKl8ZXGeuKl2bKALZUFCdieMKga+UpxSS/HGoP9rcBNF
3B7iCTZW+4JOxuzF07HHD/gOidfb/H4eYWnZqXdexUCubIXLG0KvX9gXWbF/iaYA
Rv0wi+qwWy3lDcz7lHT3DXcdZuSyc9z+l+Uk/IWjOJqlrQX1gsrh+psviGfA58kQ
s6P9wu8LSlBjoeggPmUa+j4t7HzHveUyMTCcoVogaEklpbiW+Mmled/5v5QKwpOk
N7wR7tDwWcjfXjUiqPPa7Zm4McM7D7ZGDrOhbOwyR6rynM/hDeSAwKqQmUWiE4Tt
ARO+OFYaApwhmNjHipJH7iNxlrWdBI/JpmnkqVAlhQnewW0m0eczsT6PkAjri5Oi
PV+9Iha8Uft0Gdwbs7XQXVMRmfylFnXtQhYqADhsagV+JGU/OebwkVsoWh7TkONn
g5/Edr/TSQfbMFDz5x9IvAyEjhSdso7oBjGteodmnyPknR75RkEGMBUZBHDRxUVo
R1MGIa6mqV3Bgb1z+09SMIKkywo+nGekvXa74MkkdZQ63oDEn1ZIQzOgV2KWImFz
ldC1yPzC4t+jQbI7XcxhZFdE2Ii0Y5mm1LqY2oi/yX/to4XiL3vQJWU/oLeLZR28
x8+wQI5mHTzmdPX/Urlgq56nxaKUXTsYQQBO7VBIojzOW4oWNlKtiJ0sg3KPGRDn
k3Tc2R/BSqfOys9Q7W6WqX+M2PVi3grM/aCPiMxarA8e2Klg5niZGjwutKZGhAFn
bEy58prlPezSfgBWx+59YrimPNM5j7T7m36vjycWreRhc4Q+rwjdUz3bagy6gHG1
tUx/k0p74Qj1VbSR2FKjRUcXurYhTanmE//8upH1kMGav7MzYr6tS1V/Lk3Fgksa
j8/e4+S1tVY3HaFkaDev3JKHOgyu619PMMj7XhHz6RWRtbd9KR2yzTAXeNFnU4B/
rLNYX+ggV8EE3law8PPw2knAaOYIjGzd6fNWpsFPdkDc7qDp3oURuAdcYF+WrACt
IPo+NfFdv0oTaX/0WVGMMER9qzjhT9eh7BmCcRCDJ1DUF466xgP3u/vLfhEzggWR
So/0rc7vv1u5T9jtX+jPHfPoUabWpdMCX+/wprsWbd8fC7/Do0Aa+A5OYgWqDZgq
W4n8nIm5fKRZSwvyyoptQhGPnzqdCdHKGhLyhFG5VEyX6zpaOFsLN8YKSiuRwfh6
sFEpGNpqa5C2MlfUxD3EGFNNrjKhbd+AxEdUGe+MN6HAmJQeXn3szc9NjGE3t7mJ
Sfl7Y2N6uiDcSRdl+C5h9n+kOu+4FuAp91BKr9M4h2HjjtfO+WqqujubCWA42g2G
k69jY5iYxLKvVynEoaZ5gq7nZXv4BqfQH8dRm1Hdm5GUAEWfHvA0KjdKlSL7AEWf
cetU0p+sbaySo+vyc3wy+3UjuB2FacBfRkBjtMXgmqCi604TZVHgsDN4Rrf9TDBO
pNFLeoo4ZNIVAJ4y++m/tKJX4xrdCFWdgHMTjPRvaw2ZWhlmCMtskJCrvunGdHfy
KpLkhaglTZyrsqrpiCJVk38NY77/M+v190u74Cn0I+V8IuAwXeL1Q7eKlukj9skz
W0zl0Ee26Q/WnCMGRnwWRhjEBJlRU/x+2GN3ol3EelCZHJLn91CubdX0ejbzZALB
AAaS3/xKYfS/x/CwEe2dCpWb9G50l+ifH11XY9D0cUqV+3SoThJp6GY3T8ennA+p
RX2J+Xs4IhjKrGcIyNxV2MKzb8CKm3ASOa9Gk0owyme7IOxaMrQhQHh26oHe7nno
tifZr7D9F1w/lDUeXRg/hTG97oNOQCPr2EnvJjqhQQV7y6iCZ2DwII7dQcoHuVJh
ekjBr5hI+ORTJof9Tr76NWEZcm0rcnP6l8Ka6AtoV9VAVDmt56P859w9tweBheFl
TKWlii/+51T8/eNpgREdpP4SZkxjVTWbgrxuOFuNCZnUJVL0TpJPU9uGyo8puvqK
27uSbXkIV8bl1RuC2CiBcqtQNsZ/M2Hg/aEcmlDyONP3q4e3Fs+OEtbjT9s33QDs
Knpo9ap4yvbTTLOItOPMrds1s5eIMPLOre4bBQ9GRjPhmkwfBri1XXKmRI2fnj3Z
ACTlYzKIotuKFNWkpk89zc7OPURPhuF/LUgk9Q7igxKYzBLFvC5v7mjcDDDfCMSH
P54klZ47m6E5h9gT8j5QZXB3KlSGSEqHNeSHHJVkh+OAIFyFMRexSeo7vJtj3PQX
X+PQGnWOSYzZUmEbFbQNCDxgG+y6k/WinFzh7LHiQ2gYkWUUCHUJ6Mw1OOVMvXWw
0xtu8QZN3yr2qo00+3i/obHv7CU7BynoDpJ6jXpNFR26wjWuhwPYjFBQix54E/WK
7HaE20Yk8G0xCam1XogAt7AOi5x6zl1qaUGVm5aK3WBTrZJlYa81LIXrYtlymLHo
My21FN7esYgCn/OkyZ5WoJePOjeWKSPwqaaLM597K78g7WwmzxNjppxhYCFIRXIU
iMu5Lpb4o8RTk0sDAj5am9tiIBVNTQZQXBxd/JRjN/slZ+HK7RsDBcIFAagCg/KZ
Tq6EW0Q5XQcxZj3ncwFVvNFwl0hhx03Qb/DHxifeDqED4CRfcU3cx+gHZhlVS6xk
XLoSvYkUk8qXw+5PUt/cTCAFOO8n11WVgKnrSztzB3ghAcik3lfNZx7fWEznZYXS
D7IQra89ZnBy1nEfN2DJd9Chk+z3yPzGF4pJtiQ/8h7a/FA/QJV4wgf3ZEgH3bcA
ebe0lVEmB2IE6iV4TDUcKaO19BJk1Z0EOwm1IZ054+Z/eTZzWXkjJ3zZ3QT5GZLQ
KGSSLvBBOqXTG+0h2c9ltoWchwJIFV9Kzy5M0ckVdShil5i1rH2fQqVBvzsgGiWM
4VQZMtD7ZTgdTaLj+fcyay8YwFPF/rqHdhDt2h+rfxAT6rKGBDfb4NqJrgbSWq+A
BE4E8P0RRnRkDxc/J5AVEu8Q8AVSEAYxv3X/r2gMINkfkVWxgyXPiJHrFe8nAlfs
VZLRfLdpzfZ75dV919cbEYgiri+DholxlPEivqLKxVci6TMhBKTL1U+JyS38FjZu
o8SHeHq7VqimlqQjftlVYtqH2UjbIhS+wFouI+aVLXGi8QuprkKQibEZxISITClc
gAVGsumWoLCQvEvMIjnovRiCrQEd+h7gVyBzmHSjXQ38rcvJHl9NSpGY4POp10B1
ZuKsdXvbRZmN4n9GlA3OrvpWXU9DJe8mbYKytIxmuluaICwWAF8VfiHXkDtRlIoU
d7QgzgMRJZsYfRpYP9VON5kxeaHgsa3l1l+hgPVPVQ3SZjOaPYN/B4wjs/vBJNg5
olkUCaitqPyjflT1NYB4tcfcNA6234A91cdp/Y48zTCQs8DUgPfVE5B4dVYhztlx
rSj4SXDAiz5G25jg3Ng6m6WkWGG3+GZVT+DMNilT8gg0f2cq/6uXOqjg2IBPn1Nd
keoKBq4qMPzsgTFWiZh2P7bJXHuuyFNXSOi1iM9ZTjJ4An+e2QvPIV+JFQ+QHUVk
8C4dflb8YQAcZqCl2GpXT98bWvjtPUmmGqfFoXjESvUV/Ln8FoPxzzYuyZ3KLlaD
cYFPj3DE63OPN8Tb1DLcngAoQe07vNzIT3DyGjpMim6ICKiS0uzYgaFg0rUehNu2
Mk20/2ZC1x7wy7jiZWChVT9k9k8WTux64onbDtv+X3XTqgfQSpcITNi8+/t6ki94
l//tbR7bFW87G8rNpjfYmEj20u5OzT/vaUzxpZOYvX5UH4LIOAYYjbR1H4Qpv/90
lsK/aZVxBts/SjGMBe7BCs4NFtHxt1jj7S3/X60R513xrNlT4dybeadHVI26wtVX
fUz41v1kjcxBw3s4kzDc/QzbOAFMsNb9lR18CL7rgC0ZLH70qYtbmz6+dw49IPU6
GkY/vDcYKQfkotY8SfavVVYNBf6eGRqi0cN8d4HAJfm+ruBPeYrHF9w7e7EAlW50
miCfplFjI9qnROEBSdlY3C0g0lYHyJezmKOSPYKq2WMEHmr3LTaL7iYewNnGPJQg
jjS+E6E9iJ+9zxl2DDmMVwPCPRVb5incPQ6CyZY6Qi6Df/MlvjI3zDIhmPxSl04u
66e2LSWoESBmoGEXgTpnXD82gwEcuHNYZmut7IxeUbZPSh4dVyG9PE6AzKvnbHYp
E9vrTady0YRso2TERXpizoS0o/ULhXshbX/Lm5J5YO6UyUYzFK5bsqnxV3C9sot+
/dYiiWl8kWY/EnsxmCMhWOvwWrcMeE3Fc4oNyoZvxKUzCmFDHI7BUkUQQ/yfYlB+
RXo7ZXhda40pKORX0NF8gh5pA89Dv/cZAtux/CEgAZL1fTcz3/7m0tJYGA1YSQ24
HoTp9L5nP7SmA7X4tnIQ5u4rPloZ2enUd32lrDCFsP4eMSnKD91Cncx2k3WQ0QYl
P1LFRgXuxD3T0gGuAWEJg2mBDBCqzYCJ4lsX94NKa3KeqhNwFNVQrjiRoSPsutcD
p0M1CJ/i6vNsiF2+aQKvayBreHTjBnGhoBuxdlUFMszRBjQqdsn1vhvwBJFTqIes
Th8IcOPI+QiywqaQ5q2/71npkaVu10vADemzg0soOWiyU6g3sihPzHUbviOWZpey
nOsgjPqrKkriGqyb4ee9H4lWpy3c17Xn6tVNeMRdUNKKOQPoSK2PNBvo8prGuWrw
910FvIen/+sTQ9MQYygv1gYX5dPPJcl/+QDugHWKeJDlzH9EJOcZC5zgNRS8vPNZ
5LPouVmHMRlI3/9HLDZLoQlDBf94lLqBCB0AT5IwmqtqEuhSi8qIZlsixKLXpXFl
qM28hIZNNH6CYqUfSCpbX+EiGKdGc5VWkhSUsqVWQ1H/7Whf2D2uH0fz8bJdKwoN
plL4IA05Pp47WYDrX2k2Y99Dqc3xUi2dWV5qasaqRQHc5Wf1z7waDlo7QprRmJMS
68ObfB19Rt8LUfpAkePruis4xzXQvF7I6Yz/fp1CAVo3PhK9Ym6xitqtrnK97IIk
w/EiJblVgxrESbOeKofI5rUDzUI5Ln09yQloiGUqvwK2yCZQfISEbNe7LHBM1am+
iZqVtxmlJL/OlAFa6rxrsKTi5GOmZsMAPK8soR+3UncbYmZZSg2Dg4KvO64uf80D
Hd14dmYYj9OU6Np+E0Ki3ZXw+81PWdKCI72yOTMT1JFs62R7Z/5pOa4kxjkYIrCm
HVC07rXWM107qFGcLv5S41gggvTb92NMO8sUEd4QW2DO0BTEAaOV8Vj9aw+F7mfT
6xsMGLk2+iWDYq6fiMyOl3jIOpXd2+iZvKbVAvq+zpi77RfuMJBBY6C1VIldc6e6
tY+zAPzLww3mJCrkO1e+FWk57ZOjfynWaPH+1fWCU67W+G660yW9JTGLMPrFmHva
aDgCB6ye+9SALw1KIdqpXVuylufCJIhFJdh+XMs49WUXO/2TqHB0NkgRMWzx5ND9
5pZUbStTdc4VDmtqwHpzpPUxGBV9Nmp89OVFs0EKWMKs30chXDLx53jy/Tlq/vXF
xbHI5K9dfEqagRsnTKV6lTXbGl/MrFKCoo+Q76LXZayo1LGM6OMX9wCm2HBKsUXt
crIIFpsV+mBNzBgKh7c5YRDyvzILPOfLlk3BB/VbN7TsSXA5OnpZmllv60NyyY3f
yeaRlFIkAnSFyPSDNoENFQmdwlfqXYbm/OOJX7rO3NeQTyKdIhe/UH6pDxZv33Tv
Gp+5gh/92uzCYaNrgzlLmDsgODBnxdXEalYF27EpTJrllBBgBjWr+HY+GnF+ISgX
phU5NekHg4O3xr9F4vQ05aEweZHRV8Xo4dHqH6KMm7lN3jCC4CL69FDvMSBIfVFj
qFp3sch7IzUITDRH0JW9C3OrQQgNKCkXPq14MA2vvyY1HmQvQ5q0fWrWGwsipscT
S5LDxHhj4GlhI0dpi8t4xiLw458sY7DooJiHrJ0Z9hF1zIxIY4f1aUt0rYCTT+JZ
jYUe/Lf3X7ZQOJ21BLSxQaS15wrxVOhZCHHERqK75cZ8AqTtgsWZ66+O/x8/EY5B
YMcYK6u+wi56+QX/MT2dsp0YvTTBk55nY3uJ4IhT1bfvTFKrt/H70BkQS+BaaQMk
j7hEO2rMg4RklcJYP+MyKVtvCq3RzeX4fGIdR4efB/58BG44okl7WnykE0hcEBBB
VV/OljjI3KZgwire4p7IEh94/go7Y0om9n10GLAMAECeGCX8ShfCh7U2RkozyUx/
X7A8s9fAuS8PetK9jzvvMlgIY85HPfk58kt3+Qfoh7yvUiuU+QQb8aeXjwUAVEcw
t0NVECzPV9/+utJSY60A7iAj/S3+/6IK3dbvHzjhIDnwgIouXqrMEVV1YisiTD3D
FWZ2kEM/JUhlX70iDNpPu/fqoRgce3xS9ka8vTV+YIhty0DkbFqqpI3LsgNz12Tc
1vYa/VvYWD9Uuzet0xgYL/U8MDuFfA5Rddh/PYLUiWY7Qp2aJwYbDzreTp9hiGVL
+sw2bc8th9c+72NVwol9DuVNMuSVqZpgA1+zjFWluVA9HbKaIkeBDVmQM0YXYmnb
AwefPVjr1ZA+cBLMgsO257IqTEv6Yly7HSfJaaTglcnpPNgfenzyRL9Dmz0jds4a
+VK8DZvrbh06nd1+PyUziH5oxizcCK8qQ2hKGWEQJvu5zfhdFEe+jNzGM71xa58/
q9+lsGPl+RTTB1+VpkNoPjoIFXKUJbd+dD9YjhbmQ13505PBXmgJn9GhSUpPcD7Z
KxkKB9KYwWpA5k2AqOZCYwXT3BS7ISOWhVLftzXLnNUyDUD+Yaa7cayTmThtxGWs
3pPF+TLPZSiajyFQgmktWoABaMqTtgplxaGUp6Q78eAtIY6o8E2vmsbJ18nNlmjR
EPkWwJ1picX1nFJu1Drd4Ha05iuw65UcOFg/lkmiSlcOcmL6lZC6jDhMd0Wm7K+g
n0QVqljIxGnoXHCx254gEOHKnNJS2cQKsyJ7kI+1t6ty0ua7S8AHHQSOT0zx928R
+yFxrB907IHY/XsB+FPi8msp0yok2QbrpFLUNeqr/bprBkfxqrKGlRNEJY7jpRiV
9oMGGo9tPZtQh94AGyBPeoSG7773udAqd5eW+G2+197hUypzrZ9YdGBE/ooZbCUB
YYLE4ppnaHwQfQPkSZiF7moRjUpHls8gX88ANivpamm45UZPznXGRFy0wTxKUfMv
8fjGRN4FDB+mFoXnkkBFmyznkzUvGMioEYecry+NE282gHlbYI8FA96lmCcG8zj9
ccaAPhXmjh4ptDCzoHY1jTvy9lwGfKYuVaFvr06t567jPbucUWFGAcrNYNKw04bq
vjy7jcpCX0Bt5g4Irst8k3IsajISI6Dp+mjuja9Y/oT6hNH9gCbMzWlNzyUvl2kO
emeGP2gk6d4qoKNpxw0P2wn2BbDIYh6b8lws0Ul1dkpK3ZWyD5zCx4aAecIdR7Vn
PgnMT4TC2cZd5DjDt3Sv+dpz7uJQwX20iykJtAL+0g2ysMDIviHxL9TVIPEANgdj
KVOcDVHeRuRRz1JnO8hucYaMfv67CaeykCohlHzwHxQZxYnjGH02/E19HfEP18xN
u/DccWG2a9qboM2YdgJf0X0ewFCaWdP/7U32BRHfHH96TZZ0vpkvqKHytaYHSc7g
g7mp9iqDpc6xmQw9Xle4KNOxQopZCZ6GirpvZeV70STJdNmIlD0lsJAjyVSbEU86
19sbtxIxpJ3J8X5ykYrxMlK0HoYQeHLR06whSaV0CdyIvw+myedTyO7NZOZsCHY0
tMgxSiLTCFQ/zQu8/Z57Ez/Rgn77rwUIgkMIMCxiiQ2kJU2JCIWpgMM/7k8scy9l
gWN2yuPW9h/UquhfHOwL/CoXagDoeAiTZhyHplEw0KQ+DDCblyz0RFDcMPgK4CHJ
RemHe7jAFoLiiBmQW+OY1bHm7qTOl+PjksHIQojb1YeiwoDtUfFvODnRN5sXelgi
QMjxUxlka+ii8Sxr+yadxGiI0bYEzben+g3mP0cAPfIz9aSiZwuNSTe/PVBteQUa
zVvXQ/1irt+OEqlvkedaYtWOvtikoQ3Oe2MQw9V90ID+eOi5lNJFK23N64KCxEm+
tCj+g13fwaUlXwfGX4dgjiOxzFhb+iPw5ZkzrCxST2QrGrCZvmMp9VNk/lGBeHJ2
0Q8gpXf5pYKt0meUKaZ8ZEFIVdP+q3vkU5koOtuKz9yn59C+L3rAcl8/nI6I2DK0
hnUVzc2HpK7GMCKCwRJPtFbanP0QutcmVizr/aCC8E3BqwLTZhdD4x71F5W0Eon9
ZbcEj4TuqDcIlidF/lbcy96MEhy+6YhmXM9joRIQ2y3NA3nfy/odCrhW8+3mbSRk
AwvSONINJG1vJzXqCtm3p9syVDeNyvksK/b9ZT+ite3Uvg1KBAXFCHy+bqlxtdEm
ve8RzdnXdjr45MwIwZbsPQy4BLBPjPGJbC165HpoTLTEZ9XERRnjBLM+FW3Ecm41
7pE+1VSNvxg6veZK0tzDG9JHiQ+fK4DkVQRQdWQiRUU9A+yD2TLDdJ/koo5B7JLa
Zdj/xp+xkEBQHKHR3mRWyjhaVWjoGBHxoql7NFkzSym8rNBiBaOrxyX71VCnLlGx
StlFP4O4fnH/zq72q4+KAT/B3JB/rqUXl37dxlchALut6hvFgiZHTJDkbpyv0EFY
TGlWukduc+kP8EE4m1QrzIFw+8Ri7EhCPJuud+1F4BfbzXAnOPIdXCHaaZzVjhmB
lOMeEz+YzQYID8Cxhi9UoDgW70OSz6nQFC7SesXm+ecXsBt10RrPqfOXO/YQM4o/
nAeRMGSbACVwV6OHQp8zy6SeBIxSrnsUBxzMhDpN7MKFKYA9/PtEL6b+5vde6DG4
FXAlNszG/mhvdaVlENIOh/g0YKf73JzhHdaYl80jmQwd1jwbJB0ofP/giJgrEK3u
u5nmA6v1Wo2qNJ5JFdI3a8qfYBFgeBmxBmMwe2GzxUI0V0Rvo7yotsiob4pscHM+
/6YNYZL0pN5aer2u8lzntCnngP7stKzwA/oC3iHiui/BSbFi5+PXNg/OU5rx7+OD
FQIRxBSwTwkVaaKbc5XPAZEmPe2dmDjC2VteFFj4uunAKGUjxnj6VJIYjD0f33br
AVE9q8xHtoVSrK0yd1Fjc49HmRXZEfw/hRI9t6Q8JkYa5SvMXqqcc9MXZyEmIRLM
t/DzJqxX9sq6iGbuuospGhlMFr8SSYHIdE9x8vhygz/FZOR3zijgVau2iad7DQik
uitD3MMUZoP4JI9LKCfdXWEgcML7f2TvPE+DoUUkOAZV0xVHAz4D2h0nCn97Jq60
v6oafhkejlxTSURwjDtmLGe9fBSHVDoJ/tzAFe1xvZ+xTC/NHAJslD+sBVkRlPt+
T5Ns+dOwZEmR2mwzKadIgD0FNGnKPLRj+mnUcPd1IvCvROGEkVp/dhZ6trK+DY4T
BUYgL4KLVEliFIfpmJzn00pe4B4p80qMQEKEBvsFfy3CuHIFvOP68B40ACZdwsKN
2p18MuYV5iWRlM0tFssUJ5OrxKVfAe/fmHC+b30uhBM4fQyqMXR540HQH2LMWcFO
e/HMn/h1131JGSXlaQf66yowHBRdtyW0+RuqCVCJ3O6tGLZzTiLfnWuBQkaUfLS5
nOBJIabLjqAdfuACc7ztCbJz360ayhkYtAQ3TtNv6iKfMfhQIWe4QuJCAyJvZ9aT
fdQOjKkvBakdcRNSuKT3C376yQJdvoIl3JfK7vI0HzbczhUj5Cw4ojaDWUyu1SOq
+vNKLa2nlUqkIfaVBPYTLPclXhmebrAEW73VAdAWWFaXqsGUtmP+xoAhiOVAK7F+
L0XN/tCAc+vbrk7XtFG5QBeAnjxLuGMXTSsK0nDvxkJ89B1eDKLt/xwHq6vlN98z
Mmly57LIRpcPcRfXBFZwCc2RGJhQcCXG84sGiO4IsABoEJmMi50WZNQGKKh35Ral
e3Npyo8rLDY3QrJb6MtWZVzUE8dQQroRSPbUbEwiYB50Pdm6kIiQLsVnhhtp9UXS
YqaZlXex1ANsilGEX4wB4rDISoNJ0EuH0n0Sm1tXTOPrjm/cuIoQigJTdu+a/ao+
FV6/aRV2JHzdhv8yN0uFYI3Cttx2LZw3praaCDiDgQl+EFr3wh2/aOc37ZmeXBVK
FOcbETszGe4QCX8uunaiuqvm13quBOIy3buy9nOxCtedrPqN9SUoItmiijLSAJbc
+Xzug8PfSlJEIL7a7wMbHb4xGE99pn/lKYzUVBx2l1TfsJEgh2FEs+EzJkmyiI11
W6mz57o5XfG6wjWT2+M9L3nJTzYhA8SqJ/Hn8YAEbs51cMEg3nCiklnqWBDFuqpD
GXNclq32TVpoWdmpi3rcVKyRZafvv/TAluD0fYcS+cEOCUzuUJfCgMHu6IH6+34g
6w52Gw5v98K5w8j8fqDh7HSd6Tw9KD69zLCubbeP8zGd+TWFXmEuEV6M+WxbpVJQ
1nBGLLgqi4aArVgJiB4Iv5a9IXfsYjpaw0CJAkartUogtBY2br7RZk6uNIDAySNL
syuPXqijD28uN7GtI5bpaI0XhlxLZAUcYB+xZBKYVOR5bweoyX04PaiT3uppUvmH
flZnYi4ii35NsiuWdHRULxB5w54w5Of4DnWuz+w6m+5eI1pNDuaDG6t/JilOlp3K
g6hyHwVw+uPznNqxzG0LYASSmcU/L+y5+nWa9nAMsVjKWbpIAIbd+rFqWyo4rDb5
IsXoATHHmtSzPtwYR1jOKktmrXFaCgE/fFrNX1JdQNuQ90IAGVvk+Dqu3aymwWvl
vyF+clASMoQHSBucQpzP/RGnn3xctkhFhK8MabiA1xVMEeyoQkJ/EgKqLbwoeO5G
pmmF3XXNErie5Jyc3Mn9DKbavK2Hz/Y45OC3aUdN+WcagOa6+8snGJK5buWq5FcN
uQY7gbXrO8WwRRmpCHvwt9qexG+lgkcZaK/yRPGr6rPF7EuFWxNVpgQ8+9RDaKBc
i4u76edlTmpszJFXXX+NoQu0B+cicyGEHuhJteNt4SO3Oai6bPL33Xek8xb+9Kxh
eUfpXTRgTInT9QMkednKKBuX2TsoGD2uZ7auzue6eTMBZN2gayahbKfVandXXiT1
gYBieIeNAkOdicb1yuxS14IpxFtb99Gm3yf7eOJ5Becod6B1UvXKHNh/4TESqKKi
TbkIU9Hk03BU7Uu+jM43Rzvt29g9R/KdMkL9ZLUxhzPVpTG9EfXXmUy+yy2K6GnU
nnmC5ykRCw0lAeNu/JdIeGQFfbsX4ys/kzH081LlkjXrwiKzQAoMGnwgcyTaxl4u
5CvFo92AodhugjKtbb0vnSb3OYXUWA1i1Yblv+zuorcmY13LepFCXYx8bXJOTm2K
lncfrkZD3eCwo1DeX1jJ0ZlNsiLWhZYxwWGsM+fzBSwNnR0TH3xzaYF31j6Tgsm5
BCr6Y0bs2r3+TXVhU5tDj4W/LtH4vmJmOc7hwvpl+b/N9ZXGIgOiDUNZkeukVzwB
pC6lSZBWlEl0zxW/bat+8cnrsyOXmsEIiNG8hzvrq3S85c5FLvAtKn4pwfVxvf8H
7XveltcRvfMQe3nIJqYv/kvKgKKOL+lUVLBmBUN293EJMAhpPhO6WonEHPlB6ucS
Ja1jxVyJ/r4BjkCYrSYgUW+6TAN539vPriFWCUS2TWftd770sqLAk8ag03PQ484Z
S0yp44dv57+n2MuW5D/iq81Lb/hVrKnmMkdMRcYMnwf7w7kWeBr2y940uyNIWB7S
vQI+TLmCTN7F/YB1pCAhm43+XuinKkuDHV/tH0KhS8LPe8+vmPN8KjvOb3fdRqsp
hcoI+M+KrnC0pdJDoBFUvrNzOue5Ts7v2EgJyDAkIk/PXU8EPfoalLnMn42LXwqC
uXsEEjwo3I22wh/QRM3QuKIaCz8PLSTFJ7+xHdf197tnmc01QtqUfxfAAkByi0vI
gwig9l8rtFVKTsB0vq43SZs+TrP+SBgO6ja0wdO/vuipY8KmbclyiF3LUQl6+5Za
MxKQnXtPieCwatixOgSCO4XhXF72PWbFWLUXLgzJOm4dwKyDNJFsHpsvyLpa3gQu
mN6xwHkhKC65eyggE7Lpi6tSEvbC0krHVOaS+SoVZIxL6KBMLTYSYtYkeCd7EYtq
wpoixhuon4XfTNxMrsvYSNXAI9Bhf2fMrIOYMFKNM9u6uHkg59q+4Es3mwNzUVtM
kyv9UnVI50TJQeMjbVu71xpxKuFHeu+y5bgO79QcWqHXRGqx6FlUkBJY8ei0hNBP
OItjAldc0oDFk7F/nZCDe5m++WoRGtAeoxM4y4u60nTflEKhUzDVFvO10+iENLYA
73JNyIFhb5NFJWBl02lzOLCS9FFQ/cL1QH2Jj7R0joQ+0ojgj/Od6MYun5L43zAr
hrsGweSf94PYQLDFGrgWcCi5CBo0eSHbf9K7dGFxeXwgNKKHy1ZECNdGYGnYVmhF
Orkf2VZYQCscaNxcSqRzqEx/1JDcj5Uwm2Bi2QoqGv5i3dMbhxPbL7v6DMWVUgWi
LLGHkK+qJQrgZ22sMA1gm4/7hqxgWi6Z4JhnZhzJuc18X9C2CJcrJIL7T8OneNGI
kEArAi/tgk8NVOtnm/AlV77EqwvKxd6brQUmbAA3c1njLlzMxjUJRYlULGJz8IYd
M9ALjBAlGHRQLotpFHGdCdIvaWKT8fW4oQCXw7ss/CFsFZwUgKRonKVET747ZRcz
nz+dJqs2vCD470ODXjWrw9QTclJCpPivubPcSHUb+55NOl2dRTAQOCoY4biAyYEg
0GD45afaSeYhWh5p9k4b5TeWNOOCQ0Q55zTbxXss8CDlPP4Qvzf/2lrNY6icB50C
3LZKaGyku9p9UpnBK+Q2Fb8J9HLARXfGGYo9wT8t4FCx+WoJ38YO1ltf/2mOxJwx
kuuqCQgv1a1XC0lmJmjnIty5Na1VeisqWYtMniSoIi+BrlGQc3vsxBboAUitHGI5
P4BXBgjfJ4fxZujnvdevqGA7Adj/YSUpFc5Td12b4S7F9PkPxsj3LN1hfsCawMjO
f5YV7pMCe/GiK8KWqVHhF2BIm2l+4B20EUrgUeqDojel1lkV+ndc2Ix1IpHoPKLL
RCmpMzJZx2g8ToqtFmPu0flpknLQDUNXySpra52BBl+5xRIdZxkKTqmWVcnSl6vD
4hBuI+eNNffAFjVdofREvPhxL9uMo1tch/NHPMZYxMVWy137ZjdM/oJFnKCGVnqv
jrFmka5vZWSUphakcWNkveg2SDrAVJ7IyxZ54/R1Q1trbKGvmZrj8ygONhJrQ9yY
xUcBU4QoulIF+EUpDdXSYh2wm95pUEGzbMcv+icW72zyomd4HOjg2zgQvgQjz3jw
i05iFhpblHb1de43L96ugK8mhmAkfRGIU2zEh099MaGslbrabFEzXfmI67c3wAC1
Z0UJ05OJyFXjYtzCeqZjrCBjy2bzLkfL9IEe/NXoc5Fj8oUlt188bn5DmXOe4rLI
B4rkQSo6EVkrv1iSiLOHDuq9TygVHHBNO0CXsvfBC8zqDoxMr4vBGidH+ojAsWxt
we559lcXJfeJxGswZfP5qGpOvptp9AlJFeVQCQwgfsgDnXwtoVFKVToCkjBQ2uGt
f9s7pi4dmQTyL1WoKcBoJrcLSMwhz34lVp4RPL6CnNqn+UfiMm68IDvPHFZrPkTz
0L5bif8MVFPcUBWeaqgWUBB5YyjysEaSeM9cu1WAMSNNuCBYPAZ2G9pwbglaAAHG
5L5HPplSDDWuXp35QiUk+/FwZ14vQizSutOk3X1iFGhcJeFKyoUtI35zhmMEOz2M
/UnKeKmrKeZ2vhXP7a2RAEpxIYtreRqPPY9tdsqrQsFs6hmxBx1Iokmr5RDP1/4C
yTZGotwvbt35U+AvROFdIQ/7Pres5BAyN5odTdaKhpoWJA0UM/X7JE0Z+0ky6aHy
V0Idu7wO+mR0G6eKgfefeh0CjDeBLGONkSbmh35g4eyJgKqtuY5WrEbJhfGZYVQ+
aCqWRTpuUCEY+1t/M9KKL/94Dv/wp1/7/U95wNH2Exhf9JvGKOReU1fbzMm6kyZU
lUqmgmbI8/HC8rsjq7bYvrronxDXC9k0g3aI9U0cejmSJzdnOPB9UvcLKVMgzmt3
Kbq38WKvirkwMWAHWzF6r+EMMX4ll+wy+KVxTcucQtv8nyzFO0lmLgPv2OUmz+MM
ppadkdFiNfj4n9nK5MaL0lkm31fGtX1t64t4wD0jli0WIQx17AbfkG3UvUKrx1YU
0rgAZNrDFNU6Buw6f8V8P0D7QL7Rx9nLKHgIlTQCHIU5Pmq9wsO7c6/1VpGL3zvA
435Ye0gzu7pby+0FMbvk+F/CKm1TXMt4GwxdshkQopt9ymaaoVe+9uezNiQgaQvM
f4z0GjnX/mT1QT4cSAIufXc4v8e7mPhjR3jUB/Fo8M5DMsHxpnBqg/s/kwLYOr6U
Cqv//Dabm/rqXuswCuVsyTInTW/2iSL/U/kC9YkrkitakJx/p6ZgqMNHSg6XK28r
9djhK/QDJSqdNYSilbf8K1AWio/fh9QgppuB0yp1BEXHLm1CbGKar9ONeiWshB5Y
jZp2mRw5FhUt4xSvVTjn221B69zSpbYy+eH8UDUjT77tgqRNWBd0reGBPliOSch3
gwzBP2bbd0etk3pLVBgTVR8YdmiQJdbaex10bI27RADdIGO9B46/jftICvmg3S8G
6zYrMng6gH9n9o7p+QdHav+j475er8Gq/ODv43fvjg3N0JFmcOu9emxLqPVHkAJn
WjX/+8Cc2CHLLoNCsFa+njLtpKiFuAIK7HURcISKSrs+VcbO2OtBh054/1IvM1vs
tDWfNEB7UvGLk+1JonZTr0+J/jQprFUfiHBa6O45wx9KSVG/nURe6QP+YsDqm1w3
gh4FxuBIywxBxWyvlRvutqRqYFSX2GT9XFxzH7S4C260b7Wx53kXPKck/FxrB0yp
zmw26hWKT7YXlPbo0ugs9wbmgNx3612Pb3p2878B8Ovji9S2sk6HpwLEZbsudy3I
FWU4Pd/NcQlP5z4Fi0gEmO03PQJOim/Dh9pnp+DKNpmNH6OBqC4tEA43GE8wv3Dq
C5VVk/RPlQNbkBN6vBzUBA7qt7BgRZaNyBFcMi2IH9K08nUZISwu0F7p4qoCpw2p
sNKjOs4aCG2hN3rcNX7tRfLTilrczf1+KGUmUjAU2DK0eQVfygyVjl6CzHz6eM9j
oWFToy+hYbYo8y4/AoySqlLrtQbhauJzjCBcBT0xSFs76f6Ny7pVOSV6eeMkG6xj
c01FVPqrgSIBL0CeJXj3SVnY6Q5ctuRyH8eJJm5OD3Sk0CnvZySOsITDdRjS7wGx
XFnF4uVOsMCzGfS0Yqu1JJ7kacxhoowGLiCBHIsuVpRn16+zG5EJe5amkOq4uMYX
1rAAApTGlqQkzf9ZZh7kHCTe/tq6Do1BI/iUTl4JP9mFJbfJgxdg4MJkRTVDShrF
XIzctSE7YOkFiRAEwV8MUgUPKtFK8Zlx5EurQH1lJ1MoAi6U7xSJsYgzGF74ADvU
s33Q/+KPDDdMAZOvMpXUCWZNe2qTflF1qA1DLY2aUiIpHkPkmCzsDJpuBKYIfr5y
CIeN+mQ8bXske3d5FRZQHfmApNqpudCZtHjfoMuU+a5exKVy5u+oH+oCoHm/IaHy
8l75OEOPKk8a4i4uaFDpQ8Tt7/tavWQt4DGTRb7xyTfAglu7eCywhoe4SHyBdl+j
UhT1F11Szf1YZDKiwHt6azCexxy/hhYQvf/1wf5ijGfwjOfzyN8mhrEQXwhsRngt
bCi5HZGStKc9Yj+aFgG4GyNnENMZ3PvSA355YbQ0O/cw1MFwvnU4XIr16x74Rau2
u6fyXbFeAWwrilXtKubAjYDAeVOzljbwuswmn+zK/i2Kpv0CWvdTxA2Fnf/XSgp/
zyf9IqtfzZ1AV2yGH3jteXmN1D7Xy9tkxzADyFjxz788at/KHqOkCWJ2lWwqmNls
NJmgyDzYiU5R5YhEvCcK6BnsSklVM4BHTK64Yz/975nX3xtuJlf7Qp0qBO7thH+b
sHcZeZhX/XeMrW2u7dZCKclKWbQqdC7RpGR4H6m8gv2idJ7ongQhfphzQaTOrUeP
eFbxVMSKPN4l8frQWPdDApYrHCaaRT+ZHcAPiVJsRBOWv92SXi0ebQUJPKxzAzo6
DNKc8xaNhPE9PRjvodPUz8bMtRr+AyCG86lcYDzQgn4xYLX3uiYK/6sYZR9pU6yZ
NPJ9TifVjkGqJPS0yTCEmSe7nc1E+25ZK79pt/oJtlnhJ7QGDWB0vAX+nEPS6+AN
lVah3msIILF6VO9M2dtN3zVgktkC1hHBOP2KkBatJrZBxqSxnmA4Gwef8tIMsY3G
yAiJM+8fVr9REpt0enKvJ/gEem+o1sbc8wA+Iw2o+xH7Ey+pip3dAt1ZEXpuswRb
PXRL8rTqhstnPHSiICmnzdZfiny8XxEdxSX7wlV13C6vAx2Z9edBMjLir6SxmJaJ
zVExmyJ+mtH0HFh0u6i4EI/Rth70axMx1mFJ2Q54rVva2jXQ65qROOgfBJUD+eol
c2h9HtxTzK9nFN0uXW7hL2r5+e9b7mlhfNEFqrdw1i4Op5900riZQ4WeOa+//r+F
kroYbdKr83UruwMR63SWGyRVFfhklEBNgH0NSIB7OQII4+tECVuABjh01idSghQy
dkTpLRIQFwvwxB49nyHIlmQNeYoWHbdsE/7oTjMzukvBa/Qo+SfyxDq56lhdntIu
eiYLykRLbZrDGBZ3vh2M3bfSiQzIJ6s6b0uD+BuVqVngnTdYs40pz/oj/jZeVByT
R+ODUWcW56ftStSmcqUasMO9r0yT9wPIfNqrs582EwQiovCSF/A2kSsseBS1GQk4
ufCiw2U1TLHHdvnnlxIj7ULGWGmAp6gIkywfwFeakvy7IsrV7FT/gCbGkgf68YZ7
rnADF6+XBUyiQjm3dQCeP4fPsNc9OPVBl4XIKW2ypOb5LTzLFJkydywk9fKplHjm
frPJ5tSs6qiXFenTBHjK9p8I0ZGsHmOXqmzH5UyZqAAogEC6Q6uin7kK0Tdu4roQ
whCk2ATFoTNfK79Zdm/0DkDtvZYHPB0PO0p2gDQV3vDu5MT2UvFw4MQeZqXdVLqe
ELdvRuBohNNmeDlpVIO95ZatMKrFFF08FHYqCJa/QI7yMbpj18jYbQDKqiagJKb/
e2hxGa09/5iKWz9wpCgi30oLxqH5TEz2e8k42w+kbVDYaKSRhCR5DCppMFEIMM6f
cOiW+WEXYoHRP8FsjSBZO5sUd1rh/Pd2hB6vw0L7lgw5McyoIEJ8TDi78BwUVQaF
EV37gAQl77xSV41Wuh2wbgbGlfFK1zIDh6V4hD7ztieEdDLNJ9sGAJom4xP/bdaw
eBkpoztILh8wzn1hP75ru8Z5hbbfaObZy4hl/XfAUR3smV0rY0iQMkVJXq7Sur+r
lrIike4yzguZq7u7VE6tJQGywfmmtF7pueiXNKUpbeEgXdY9ap6LRuj9ngjins5Y
LA5MTTx20CxEoO4IXIBzcVXwfQzJoXtBI45+m+g0rgAV2lRu0TdYOOMpIfDZGKsM
LG3zO/sqI+IFE2ReA/3nxk+7bQSa9XJIYxrf1eBcuc5HS24MZW1ZV72kxbuC8y+l
SfKs/H0ssDPWhziLS5Jo2/0bP6rz6hbvGkkhqh04kFXrzIaOCDyG9zPNS8ZxmLhc
SGvbE31CRPBWjMoY8anmfBsp4wUCWNHD3KBJ3eA1u+pP4f6fY5HIwVAS2jBnkVt+
2kfo/ZGxTBVxZNo8r7c5CLlGr+/8tqMX7heZKNgDzUVBHJ2Sl9NeeZBdmH+cxUvA
pJgXKMKdQ6oFb2R113qTJnlbPLwT+DaIIBLSqPFqwD+WumfPZJmo56+l8qXXrVzo
tLvJlQKvqsqu350b1ZqSyeu56xaYrsiJpcghUmpmVeOdOwALMucA95kJNtnvwytv
0QEuA4nHX8L7Q/j/Woy095Tz01BLG5jUc+O1RTNHvEBo4p1irGkmjJCvyapsYCmg
cP4pmO6cjETH66FpfiUheQmelI5E0tljH9NakNjRAKOnUMOZg3gZJyT6OZGywzYx
pH66BHenZjEQMccbfHFfF8wmUx46hRHkTs2z/ycXRTHJ/2nTN16PIHjYKOQJKIcY
B5+3wx0ghLh0XtpsDwCfbojN9wfdR4nkHCL9tFpdhJZA9X2UgiaTl9l80s/b7Mib
f8YyUwz73icAkIuuemfHsgAebnwI6IpQUmAqa/bjhmkpFAFYH02Sszg1Z0Agc0GF
3EZUGXQbMq+R1DdwiGuumYv7rtstHlT/SRxgFtGMZhjZufXTqFHLNOgwwXyzC2tP
UsnzmZcRwYF9xANjIMYrvs5uHOHFlcT2neNtleI1tKQN/fOF+y2iJUR+2BVw+jf6
UNA1J/S/ePvj8NVS1KcYo2kDcKzok+wiXxdefKihlHG+NLYljP/O3dxxYoD3K2Af
np5BYORGTLR9I8xVLKxNhfAFAIGrClvOInD1XO72JUqaPTZFLxKRWjJZ7FaV12Z7
UShNMaLNi0mXnLaDlHGgNzn6AtsgjkKa8YYtadsW0YWRISfaW4uGFeKNJAFwhPXs
ZWbC7HrVWTc0g+yVpBpGTWC2qN0z0bOrfFGHmnOCqENoB2uSgNE+nl/sQi9cm22l
inWkYVVtf/xm/uZS+lNSOEp8fzZ4wOAdrWWg0d+GH/Bh6fyebGoqS71Jfeum1Fwf
eME0gWg2BLg456Zpw8qvehPcnLy6q5zyty4U5QarPXt4+KtY1kl038u9edPM8mR8
1ztIC7Lnt/VJIIWNZ2NbXWLt1RVPuxRYYbEbrx1Oh1cLvi0awxENs8KNfke1uTTf
7Sol9yPgRhVrcPaSNjG5CF0YIxoUFr/fNmYynHHkX2jFKQOIVGXh0WbFmlzNvUXI
RVIOL1yvffClN7gt2KtQ74x1WRLOe6hin4H4Z3rU+q1thzKvSvUwB9qTkaa7oGfS
QFmEZ2WXcBb9+HhuBYGMG/EJ8EcfMDgjjjLSISntOsqTacoogwbSITLg5Dcc7r4e
reBjmcZyyD9XBtt2I7sXnOI5T63oRTyKX+/kfHCishvXSHfD1C80VrDRmkIMXt7u
k89YJ/ZcSR0Il7fgGoBqqVkRGMKiFBxMaWtmFFFmVj/om/otTVxyC/LgPndmnWFD
wLwfHa3RmYp28Rn/g5Y9RVp7mnxrsG9JJE8o/8PX+Ax2o92M3qySoUdsGj1txZCo
Jo6K+WRDU8I/1TGzBnC/NsmPlPRuSp0frFhjyi1rS48XCGiQimz3Vqc1V0nagcE6
Nfsn2bvyAkwK1aa4zSoJG3Ndb/425lAttVgjSPIoq9DDMYqOp48LQ6r4CFu4zEsf
h7AtVSjzyMFVcqRVUcf+GeGMuRl7vdGii8vnDR/DKhzSWWxKt2868xHO1yheiWQN
J82t04hwhr4xWUE2hoiMA6niEsSzYPOku+pw/8VEE0B2KadluB4BMaC7SGRdf8ws
NKDB0l6tFY8XPodIMc6smg/RiUB2vj4ZUyDMwGuvb7I/Iuoke2+bB//1jKvvzs3x
N4LiaAkVFnuWpyq4sF/VZUaj9LL7grT8ac4kNL6CEc1xn5P8unTggld+sU/Fq60S
Oxyk4nU9Fyq7yWWRcub/gD/28x7Ej2/Y4tNC4vnMn3jWtVhvofVKlg8uMXpElrvG
ymMFHXNNt31CAhw1ejrSTBRNbhXPFQ9QmPWwAe/pVySf2EgthIrpGNVESFPP96Yy
JTOTso1sqnXRjvvuW402cBqTO+J2DCf1DLvWV1sAuuTwB4T512LOmtzYTNR380ej
jbWoCsEsPO4To2To/uWgtngXQIHFdFOs7BO8t8N0p5riZPpbJddh7GjVPO4Gf12o
ZcM90W9npyEvl649fta2JO6PV0RzQSAZyQ2eNRHhTbBVoV0ig6HkRgY72kalQtaa
5K5li3Lwc/vJ/6SGFMSPWBK9zFfL5bJbHmo3qn1E+XT/gd4M1TU/4K2XH7+ZBV1P
vj+oC6uRSGki0uTsavJmop6M8d/tEGmgH9xNVOROaFkQyXAEfFfWbK25PP38xu7V
78corqb3xfPVgw3KZ4QWS1I7LrSdaFF6fAnOTu97YSt6nBpccHi053GeA+YqP6Jg
uoiWrHviiMYD8U366FDAnaTr0ajgUgHe8V3F4QAaStCICTsJ+aMo2+LeIaF/JDdZ
QDaTESjEOno6aOwM0LX/uAce25frtuOnzaHNsgTdg5gn5fGY7pLmO5b1EXNP6vOQ
GylK0J7S0mRxkxZbL3IgGD75xHtf8RYDn2y7i9CUo2lSr1KasylHJYfoi/+1/0Ag
joDnewF3CTGUvmOC9OojH/r1uPQsd3vP50D8ooeXvjC1hyU0nveMGjo0qHjerVvd
juuUZLURzJnLMrIW6ovVp8GXd3ERz84teMXhjRxBIAqz41C6AXz5goHXv8fp0SRT
wSZ9fryfJw9md9lzOaCxJuXtl54orjE3hyUF5lYgfFiOahrPgyNRmrbwc0w527XD
rpxqSvpnQ48epSw1PHUqRdfQAgCjKXwJd85WtIb61ehGAO4vVcy9CBQGmV2sltZM
2GQpVkBYTQVrb+5NZ6CyRd9gOTSiTriGcyGLssvUTeOaL31QqAvghDWWZQsevg8v
aOFb/FDq9Ah7uiLWcH8YC48FBs43+iS/uOik46OHKSFP1Ay420ggmIRQbAW7Ky46
hyZE1PUiuhZzXSFWe093J4vr3stJKnDZFzDRVKIZnU+5nYj1UPr6onOeTwSDrKhS
79T/Y5+2NP3pWLeBqmbzfrk4VEEEu/ELQZ/j8ca0GjmKxMLf+geInktsyNwgSjS9
7zSIcAJ2dSuPZ9Pkp7g4ABxXxi1vuM5a9ylHZFUiyQk2BaDCg3WOq23Hm01QMKQG
ISamryetQeLuEJorB/nfaaVQUo8aMnLbeyS+p2t3/USSDoeMzbFxrztMRKfRCwwq
q8BCHbkP1UZYj09Ww6wVqWL7mYTwijPmtCq/0gTWqKeytZZ29RA70vOYDSAA+veM
QVtbUVjrnUtYa/hNwJy5MlEg9olfSoDlA1JEntOGKevj1a7M0GPRS4yaFoww3ztp
VM1oI7nxxxUz/+3GvooxyFb0mfDtYisFZ3bVNITGHH0PH3+0K4XgmYXzNIdCgjQ1
DqKl81Kehczaw1vvHIWWnca0MZjrLddFeBwXQMR11zrB7rwv7LDBGNK6nNc0qMwa
wfEeKjV2rIVA8BVhW2JozGZEN4/b94lgtWEPjrEwTFsdFRnjhCmHJzeNm6pVjsqF
NzMRohAEecL/XI3A1LpJKPdfAdpOTeME7x3GeQ0IIbp24VYX7DLG8u8SLLxb9ujh
93ziNrROSbhSOGjlkRiyDcbd2UVE2KERvVH3qebcoo6nxD6eEEp32vg1kWiFfeUG
mluvNo3Ieg0ecI1jgtyOJgyWMcBaZ7sey7OVj5zJgNTEFguL6vG4z7udglpf71Av
alhRtbTaNOBU3/kc/Raf1Fe21aPhwGhMMzttTnmd+duNWziwRYENKpOBCJri70cL
Oesas1YO+7FZhocqO8xFqDACcJP4feiayKX1crJ/QZaK2C6ZvL2ncUHz4G0p64rL
7hmu4xe48PV9KcmOd9w8f0WnsISWFWqDNWSNJ68uqXjddqiJnybVDKRb5etqJep+
AA3QwiP2LB9iXN8yo5gVQCyyfaOWo4l722KLW5hxE6lbEt/jMCp4I3ZBUXfFzNsX
GTZ31kt3avHDNAplyUe9iEm++cnNKu+qBu7hMl5ffkIefYpKjlSfBW8K10HxBpis
HbN798iBadhmweG4dq0HW4t2orcd0/WRE/N3Qb/gCAs5gQSwTdE3nHJ8/B6OtOxr
2GEDAPiTOiLDYlFeiSnIDyMOxnnnVqeWGo3T42uUZ0esafoo12mRpwMozw7wh6+I
e2iRVZuJHiGsYhSkiEL9q4MizlxGSVAaNpQDPwZTFcDiiBETYiG9H8P0Wa8lLpaK
FDdw93mZkD+vlrPl0LYIyFHAinCh+tciXGNebb3CYXcYjhfKmwLH5KABSLWTMBko
/ctTADBZrAe7e0pUH5xv4P5pDcfCC87xnTdvtrxIedZpIzZKKNlcdSJAL2bGEIto
oitSxcj+NEWMH1seXxQeUMZsVL9ypdo3+4ZCc8y+SXnzDUj/24lQgORwqyIWxW1B
sWhvYTXtRwz25+vDnCR5XFo+3fxqZBgxa9Yaeu4w9sOkFnr40dtAx761yH6LviLO
jxP51rH5jILTlAg8BtbxndF3HGsa4mBWqkfRBPbIV9xPOPAWChSP8L4b8YEbG3oO
XV4eDHfV1f1hJkrpT9BKCxwRQUp5GB8U65hdFC/V6JHNtgLfcAYl8opm3hlzJm59
csgX11Xw1OTPg38vHzNtzfiFH4bOpKQu8a1hheVi/quE2eY3T/ms/1Enjos9gvVL
r08VikG+RGdsfbLPWakGGJyMleSQURUhlREEbJKZDuhDtHNNy0GzRxjej1P1NtGB
J021IyQUz9i/roNWr/942RE4ZtGVUatUjhSGljyY9jM2IgtN0vE8L4znwQAyYOEi
Sa1xjSZAJ4St9bgMUN7DA2AMPvgwlZUWmRDb+1x28pyKaYRJWxyg+1AWSFj+IvU7
bWxaEEI3eDYNKBdmCg88l1m2YR7SrkhVbaeM8jGO63jky7bI0gnkIUDW1RjQKGKY
bIZ+EHDh7w3/6OlAKeagT16gu284oBjvyBo0voiiBfZz0d+SSbw/D+Lh2EMWZB1R
t5BES2Fl8gg+NJlRPn4zx+JmlctXFecq7f79gFGGAmWocOVMVWy9tTtNGzlMpyMM
ICTDv+yTW95KsSfQCrZ6RP6rCr8L3DsxowlY6Lk699ECFYHqz8KeZSbNBAKWyIxU
EJmr3m+/2qRsJXBYWTY1+bJtCa52JZrUMbYquG4j9bR11TYLil9lNpb64KVfqy7z
R2CAKn4eOdr9VB82j9MWVR9E/DgMFzztpzSWxq2yIblYWtCqVhweNakF0K1AhwFU
iE6mUKZpxpqm53Ti5w5Q61jpu0XiynyVXVlj/I4/TKjKGJK1cKXK7gRXBL7U9fGk
jukYGsPUz9+uZ7qgwlB8Unuy4WG2i8J4CP/IGdJDsPYYLgSEpdIK4ZEHyH8+n9dc
TEHAYXOEAwOiGRRNe1i/ivshHqrH1onYzvYc5ZeI5lsXVuzGVGNq87TvJEGzeICh
66aO04DuE/GxViq049klqP4ujbLxdtwRdzsz356/2ZsCs2PvdAP1iew+EiuHC6Es
DB0P+g+rxEWp2cqxNUc9HK9efFLvxB5LgcXjlbIcvKglfdc+qETQ41xP78dVJugL
6EocqqBJRJDycygnpLArf3/cLalvH0bRngOCTiGVXAykTqw8Hjy7bGL8W+86dX1i
4GcwobtT43KNDGSy6Fcuxp0uN5EquHT7QUoPZPVmtgLEth71xEAGjuSIx7zFILJA
xHnoEoAWJHBdiQwX6EpSuI6zjv51slWnNTojAoaxawj8mKrZ9tpGLEOl6HcY0HjR
SP2+WsrQsoWzBiELp0hKX4kG4lOzdyBjx34qPfVy2AmnAUOPw+KHIpqNurLRDBsy
qvdDDCV3BZka2Aqf0QNfpUB2PlYm31KQNV1QmIBNtRpGNHbjrN8VGjrwciCTgK2f
QJyUhUM0UgLt24mV4465UzcR94NcQToMOdHH7tWlFr9rsMkDj8THbEi2ai0oWkhW
ZcArXQz/UNFEIfEmYkBjbbGcdXH4+bJNMOIR/vR/7zXJXnqp3Nf/iawyNyceqR6P
1LoG5irJx+8Kv+TiNA8rI6juSn13YkktX/8wW3OQEzvVzUiAQD+L1bpiMIK+BDe4
oL6/dVXEQ/aDe/dOaE5GSL4xFahKYhQVrddf/Lu7iU6pP4+vNagWfJGZnXsZdOq1
fIoNDKlG2JueN7EXZ7wNgfjybZ331VGbybbbueHQOOs09RGGyi2SSJT6QVSNsn8P
WYedCRJqsiUBECIrdpAocyJgYN1+XfET80I2/x9wU4z33WlaJskK8gVePBOJ9hOW
NZNn9jpbs1cjqgfRMmcTYGPxOF01h1/ATn6XnnAdXZfZsfWhVAXtpK3htv9/WSY+
NzHSy+viBvpqgKMgeF/fh5b7O5XzF9c/LpaNzbBMtz/FB/06szztLLB7o/YciePu
1LK5EzueSgPzj964UIsnPAgBe/nC1GNQeX1XiYi5yQPiL02oKN1MB0c6hWOrEaYO
NwHkSX7LmumBUM2jyaRPxglXkujD6WK4t51q1aaABLOiGJzUTeSMv/h6mnp24pzG
8x6BbwObRgfRWUE5CrsobgTtBAYbf+jKYSn8lnJqY9evJwX0KQY1ZgdmDeMD3Ws/
3LYa2QSBRs0ZwWUUsrqczWDxZjWe8ZgX9cfuj4hSj59W9scTsFyK9AutuuJacJb0
cP/I3j8DK5KwTfOfqwoiz2DZ12a7UmlFjhliehvqVPYerqSrriIn9g2TbhVF6RCd
BPQQ1pHx3AW9v/W6WtVedVC/PFY7gCIPuAn2xL8LzxVfq7CckzNfcBi//vQeEHnP
21h621qOZ0QUT+XMXUj6GQLahEgW4+oSzI4JIYGzPXhl6CltMhkP+pmnH3CeiB2g
xUSpkTQuKGCPlTZB+Q+32fCNwpwq/3NpzX9GvD1zpmkkRp0dP1y3P29f9LYCWVGf
muNkCq8QYYI30m9G2Grk9H6pVeiMmQgw/pmzWoikbLyPaVUBEHZFQjLPBeEi1bHs
JEMM9gvlFlJS4jRI1SOdHH0tfii/9slYI9HEJsx/5eTkNPuIqxJepzAXTROc+JxA
EhYpqgqHF7Ic6kN+fHnVHKqe0ri1bdSVYPP90x1AtDrr65B8TU1ByCrkD6azNQEB
7BrD0MjKBv0IzZ9Dvljk7qdu1kYII7wyiFt4FPdyalk2PaLYmXScphu1OO9Zr50P
2+VJM2MKLO8XPxeyBSBx6KRbMkhE9nN34d7izfiRAwS7FCfDrOFr9cy1vKFy0Dj9
veKy2Hw0BApnITxun55LN2UPu+QXtUKCZWX3qW6QEMUxhyqZ7Wh5fz79XiHH24rV
pvlpWU486JJMfemscqaoV4qHq+7nZayfC2QhF9Y8ZvAFGiYmkpIKKjbruOWQVWo+
xVblWdExwE25vmcLd15tGBIJFgzX73l1WXz+SaGG9bJxoD0EmiMtXJtVGus6xOuA
BDSQthuEN86YhlRX5mtR2rUylE/fNh4wmFh+CcmLYSR2zNJIf4Z/+CLcUJIeH3eg
PGGesD/czwnNiN2NENYE1HGvpOR4QDwO+9POxNCJFDsGJG2WvLyENx5ZIzaTiXNN
kFw0f2Im5x7ZhXDqbOxMa4LjWOQ8b3lN9/u1ls22sv3hALnhm6vpYqWXxz3QT1CH
HU5UPZxks+vIMz7Uz+fai3FNbJuQe9TOQKyz9EqKZFeLLVOQu3nLONpPzZ1LJIWW
fJLsHTFnR/y/8kCXzrxy4VeahlvzEqukV1O1rnNNN+TmxZPrgyg9wn2TlRqimoO9
zUfAXvg3hFVjfjD/YtcJ4rqMUlKzyASroT8/EO5z8la66Q+9eNTTi5loETr++4p8
AMeTI9M7dnrRkuk+q4psHoiskZw5fmFYJl4Zbk+9VYciPhE52alfZgbJvo3qfiZK
/HP2rRYJKGn/S9Y0++3XTgn4MSCMx0e3U1XEqZ/SG0sofm35JViAa/oUnqMp/t4C
08J07T5OLbzpI4wF7M3S8Z/OD8EOtj9FbpReyPpt0MSwMWAkn7nIMg9F40L0qCNG
Fz9tFHVr7Vf+N8J7mt4S+wqbp52THFX3U951LGIo+AQWcrvXOl3aRYGcrt6WZjjj
2lM0tWIsSBFI9NFg+nwP+/WE5CcSSJEndPxll37IpZlVggJHnax26Zrqfsc+MWXk
gpuo3L5TNQomxw6CnfsfO0WJc+U65jy6K6b4JDrJCrHgC0CSStESCXidTTImGsda
EXpadgUfK8OHciAvJlz5cp03e44k0i+jC97ZNLYGwqO62bzeM6mFKNvFnrINBesb
pL2ittgPlze9JhlW2pwF7O72RWFseCcnun15F4/9+cPC+x2qAmEIkxEILxo5uFhT
eIzyDxZZPZYdBuGz/EzoA1h484Il9CCT65KeD+1BqJJmiXmBKLbEM7VYdms0svkR
3lleZj2a+LsjHg6C/NnEL9DcQ+K4q+CY6KHY9htY6WXnK6eEaQ5HtiRLKw6kACMa
rz41adrrcqt3tn72VUvZP5rLDfTIYEafjpz0ur+/PVdAb3OE2GVHbhnrt6ELT68y
2fII+iL6a244dxDy4H8gGwz+eswIn8JQHsWldynQEK1Yer7cN7PXbxQY+qbsvRdi
f25opDC1Oy7wpX+UwNsqeAUJJgvC3yijoF5kiN/qjNKmKGwswLCtLZCRtksEX1b7
FtrfLbadXvBeaRjil/lBRfnXxPZvwGqONgIWudQSg/V+mJ4BXuiWQCo73FXQDz7g
lyeI/JVe0bDKHiekFCQhlAPTLhVix5hlWWGv9/hNu+f0dro9sAaWV5+R36OJ9xCz
v2uDq0uVNmsPhBvKh1wsIDjV+cOI5WU0oGlv8jFmH3fkyERH7DpQC+X/Tc61NcUW
9qcC2fk30SRcnuzsVhzI/RpOJ17+VMxlBaLuRlQWJv8yLZSryljLd9bgo3C8usBG
d+Pf1knazBA4JuakbJb6d/0POT6b8rgEMzgip/FPvEFaiqCQ9ho6b+gTRAdY1UKm
oU+rTEsLzXo3FcL+p34Re1QQvLfs+sN7wLXEvGkL5nf7IThoUglhuydiQ2YM0WzD
qlveGlYLCl3gRNG3TDGvZre0H7NUlorylDFEHpcnYxkRO54lPq/Q8CfMqsHaU4Uu
3gUpd8CEBwFtfUlHvXybSQ9U1FPkBQ1B4Z0DQ6OWl29IfYsXuTXi94qT8dMt47Dr
FefbaIf7HF87x5ZWqToadcsrgaM8WIItDF/OvoAaBFyvW/bqczNRvWiE4SulogL2
zHhoEzUqEynIGTjIY7bKptwXw/TNuLjb9lFMB4HitT6hTJDARXprLFvNUM5Q0/u1
Y+4QEDZzRv2xgfbQjQy610ox+nidXdunx8XnF3oqLRKVpWftWIoVk7uQyHlGkIH1
Cae2Jk3AjfVASAG3w0ZSJPoJ2YE2aM4EvwLKqREYT9itNIvpJFEh42lUNBFrSBJg
ybMq7HqaciVdB+thJOozXQXB0t0t4776/9p562avrfh2Py3ucPjwRZDVzkU+PBQ/
5us9erfNeIKNFg6icY7CdOuEF8pfzADQMNDqRV2E3wiNFmp1scssJhNm4VaA2l/w
D47dRet0HxXjFWE/dCHBfAExyL+9l6aIJzVNaBpOoxID4ozDTdd4JnjLrJeiC2wy
q4JDEoPK1BeWqAAFENI9/qmhQzpUE7uK32uev3pjpchqlO2Qq3Dev8JuVL/G7FU3
3PkdFoSClOlR+hqZBJc8Mp0fY7zBGmxQHiUNr9gwXeHClA5V0bMrihiW+lTyVjH9
RSiPKgGvUxWaDKxP62I6V/Opix1MbSD8gF8vStk/v50GoN6KoxD9O/HHFNYlgHJ+
dVnFJ4CJncAjj80AZtoEAChdIUrnVO7n9raJxzpHvAKFqju8BCxAC8ynVoCvhMU2
Ln9BmqyK6BgSmehZJM3dwUStYj7YJ7oozrOEIUcUh/CGh83P426p6fHR0TBPxDhL
OkJT+LGnd9REnDtAvv/3qMH+9q6AFsdk4WmTFjQRiJR8b/JaZQlWIX/QMCZhgXuq
GLRNAR8xVWiyQZmYADXdOZsUcN95YVTSET21SmArroqFQa+RLHhrLPKUdyq5H2fj
Px0BUEFHF/vIjnWZ2blC0naovY5uVAfFwuOwBx0uOZ1rLosGKAVPTlo+NR2ooAmE
7R2z+Z29c/YA/pG9exEiIuqzUw/aRwmDfr8Q4imw5I89ZIh1B2Sz0F4RGp23ywbY
1Jy98i3SD5rxG9ehFAafZ7qwMWlXo31fPrFSvQA7kISvrPQhw2FF2PCTIGBwL4wN
w7EG8hny0dD68ea8ftADFLzSME1d/2UBzCb1YWm86yBcikUiKX+tBbvgY6wSmlWV
Q+osYDAm/CGmerUAwpArWbX4m8DwyZh0nW7alK1gfXYFv2Zl7rahZvfzk/WIEZm7
1B363Bzh4afw9Y88USZCGB6v3R3dU3eTWjtBM+Wm8zCNDjI1yBODPW4IpZB+PSds
FNZyvNJen96hCfz2Oli2Q8caa1Bq/H9xGyGY6AOm4+kxThKGPUDqEVvnYudB25nk
QP97e/ElspykNm/x64Q46CGtTUi83ZDNng8sMNqArHHbWflq6g4K2vb38I2PkY6M
0yzV1f8qnEXduf+OsXz9BKdaUddzI6hWemD/B/7qSlCjJov3SqlaibAvgRwH52cD
3DsbAD15CjHvdwTABjSec1JOxlBq6r/E4udnpPBkSTQ33IlNp6W6o35ujoW0QXGn
EPl5bkp85jQQe01SV4xQYeV2POQ3o5chOi2GwDvZG1zlqoiWJQQUHQ3R0nrRrPPL
WTrb5QGBgPt9NskPpIPF0u1AvFvQNGjO2qskGkTei4TCIWJpPQq8epLnBUr7bG8I
4NmOY8bbBwDYdFdew11KkUHafj5/MPKCUqrGQZfNNY5R5UOjzQ+SFAVbcO8N+UVN
SPW9pO/+WfqaYQ6vOFk//g5V/acv2WWXilErJ4QtKeLlx2qQkq1FvnNEujaEFHS6
hBEs8dKDZwwL3m07dADciKdcPm4i1qUWu855NwujlKR/YNg+ioJiLqoL1OMkBhJ2
2KNSVZ09AzOc/FXBLQf1pyetbfGjzgGexO/ViTjjQrCQS1KeIyOC/5CLXhe6vRjk
cFYyiDz4a8FPlEepAFMZ/CB9sLRH+CZeGkE7Sz+VGCG3hKl+kUVtE1H5NV3PBUye
cXT4B7dwxVY8l0v4+e7FLyUkaqmw5b814bzJwATN3ksz0XmHlx4Sqi0DPZ98AeG6
O392/Iv6Lw7+jqpiMdyM6pU2XqhZJIDSp+D/r6mY5XGuhR1bonEgr6I5hZv7fcVx
lwELKVF5Gz57hezRI3WeoJQeJPcoLGfxjT5NueCr9jLPyZ/QwgdUnY2dfLU7FLNm
jBZkVwZsSDgmNS4RV7M5Pcs1N9C6FxNUt2ftMB5i+xiD0eQOryyIeoLxysWvDYbg
bx0PY1T07D/rR2WXbAWEg4YN6LnyJlYo7SJiw2i+U196iO6wOrx8J+89o74x8xsM
L3XFM/IV4h1OOVQPivAGjsDwnZKCRtkqColQ+8uS2ZzR5+hI8cspI6EA3o2hOpV8
Bmoy52BHlGG7uQ1RtkNsmMxRN9tlSmc58MLbYYvdiPj3B3WHT2OICjXThsS3p4eA
mvGuvGSgAqPRYRh8RVLBsxO5dQjwttLmsSU5kY4CuZEWqaf7UOUYagqz/82b/chK
vIhN4w5bCP5iFdDSfTV1MxbfsIm3JeLzYjvcnGF4XBPFP0AQOAyUPmJzsNv/vyHe
N82acSfXx2cHu5uHg0fhsHoj1px7eJyMcfC8zhVc8wMEoUMt4molt4PEONpd+Q3q
f2GqcszKfwC05PBbxrvaL5m9tM4r61q0dafA9FiJcR/zvNR4Y50bVSPcHOI7Hul9
MXoWFiFNcJVTjb0IvPzhacjPKyy4klnz6KgLxghocqiMTUDYgfci0az5d6S6MGhg
UBN8rZ/dDZTwE527sHlaxWUZmliRh11Fb+2n81j/IbdCkQbhtt4iQZ33b+wPt5bp
DuIDt2hmplqoQ9boHnfjxUEZMN3kIwvj2DgGSGflvy66V/DsDNspI7TEH2z7UxW9
5KMHmQj+kpzERtaWw8+Im6wAxxue3waIFzL7FrFDWvMlCkpfgGLt99AbSanp07d1
bQweFKz8hTmR3tbmfDEYEIA+QCHBkkWN/OraqcC78QaWKTfUsVJbkQzEqp54G7wc
LIL6iDGhV9NKGrQVdtefmRHS2JQkLI6C/PMYsTA4tg3gAhr6ZQpAUceF6p8OssYj
KEJ6ypbJmjYRs6Xnub5/tO5/crqVmQpQT2NJGpC7RMlSeRMTm3CDQ8omRi2HvWUA
5xwM0Rk4AwzaOag4OZgkegfMdGMaljV8gsQWq4/1e/nmsaBxest7jybVu96par3e
DpkdUpWx064rW+xW2zVh9yAOt9OTjD/LZTTiauyyCuLoLku5DezU09YVsrV7+nSo
8ZXkRGuPVp/9/PbRJXGIbTAXGEKMKsG528stwKvT2nMbPrR7mJv9wpGCRi0GGIGi
zi3Kzjl/9lm2LbTKsvbMAsdDFe3/Ygv9F1Yx990KNfuRG/70asJWXhQ35wGJfq+i
c+AY2IS2TkJTfn2XkCizCsRHXKSEEd8jc1T/Jevna/3raDrb86UsY2gs4ZIEKwYC
ku96WIR9fH1HqQijSPlTWuWZcD3t4qQ8a7+B46/8zkFgMBzCanyUm3R+aQlLB1Ax
NHK0A2E5JaweaPHgGtrHtHoIEWYHBEj1eGOQvNOm2FM9XR/D0soxuYCbUwCd9fRR
v8XcWddmkAoRQgm4HfWsjZkYvU+Mp3Vt3cwpTsqA2QJnskojGEdpLLya8EHVzQKb
tLfRsHAtEuvtlITCjoj5PRaNZNvKA4YG8AUZ21GAd9Qh7FZryeZXcgpBJEzvooZG
KjLJxE8f8pI8r8KXkTHS7sYG6YDHNqpuwiE1EuAcSzyEJioRMcFzaJ2+YgCqLwBA
+w7Hel46m+r/ygXz7yYd6BEEhui15eX+YMw3eT0UaZA3//EwVJK200PM8GkdOKvN
2EVYYx2p9TgoWo+O5M+UyQPutO2uxKvzHEopbfWLPQZR1BMtI136i7PRcUeQzZcG
jI1q4c99Ywqf1CodRf+j6qhLfwRtD1VCnGqqff84COIBtmStELW+I3ZQ76unUAW0
0JDEeKIxCMFeW837hBkL22VUHIpnnOaiS/aGI3f4r2YBT0MvFA8qkUJIccC5M+rH
sFoUQJs1Ype+8KVXmodLjHS+k/ZiwNExJ8nukJuIY0riHxVIhGt5oyWv8t2UaeVa
H/ew0ploKwO3h37/bqPRTeD+mrDBhuxN7VyD8mLglQCGshLr9yyY2wCf/B7rVA+l
SRPl4Luqd9iV6NkLe8XLtorYHwtd5Y+CrpIY+bT7JhvLJ9zfjJZkglDpEoVPF6/0
dj5smVdNFJbOq3qLNXBk7f8Aqb+DqudJ7xtR7IDHYEKF9Cigzkvmb+d5/vNLS53Q
qYE6mjskNYxULeeWRJyxPjOedBAgjlj1My4xxJcflgw58FfGQf+lVrCLSTHfeh3d
DbWxnLSaerEHwzLG8fbt6mkDuOd1nkGc7zKs12CQAP1K0mTZBjL7uqlCSF22Qr2R
88x/ivGALE2rhcMAEIb2fPqMWqtTyB6lltbUJPhrzM5EDeS8ejgOG07Oj9E21M/E
aouFLGqMGqhptq75gZZvirzieriFz+LTglR/sfFQ9gWazhpWYO/8lYc2ij7tzFem
wTrgTYlrMWtZ3xVIbPxChm0GnafpVG9k5hJNQ9Vle3086GnN7eqwbdLBhyL+lMev
K+nAaO7MPGqjUNZVRDRPT22SglAIa1DogHMcnkLLawcYvC94aVY1f2MWMZqKXfYx
8V5wztt5zHWrrUSLht4eDDlAjgqsX0VQbM1lpgu8k/XEtBVU6zTtDJnTWjVSLvwz
HnCo8LE2JDOkOfoviI9FTVYuYW2igGE49FsIZInJYUeMpwA4PWXpmhPJ4or4V5ak
n/rNM/r5y9c+vGv5R3rA7LUgK2LeMqJZNkh/cTTBhOxO0Wu0/UuN5UTqNNEWWoFv
M1TPACTgcVnx6VzsBaShHR2KznzWDm6uMMyHvrqytM06jLJtbtzJynPQ5w5Sf+MA
+Q53mOkP1djNHUn3MSBAQfuX27V6QSYafc4cgavPI40Xgh1e27OdWyWPhVYziW/C
cIs4BMNpeMsrVq4L+f1ugnQ0VH5+h3zWscRMzhu7hHDtpjWZUh7DpEsFvDkRUE9V
PF4GXD+mmu9d8c7kb6At7zgQBpOcapDHgHpSRaab4EZfD/j+S/MeX7gY+5oZ9el0
j36LNL/6ZyiyNlSxyggv0J6hvs57MtR3n9JFBPT7N775ry/kR9kUS3aFBXnV1JrM
Sc3T1kHigcRxhAkr5nju1HDAwS/GkHju0tQKY6gEH2uaG9Tk3a+I9xCQwvBztGxr
0h6ms+etwu6Xc7Vg/CMHGW3sqO69YGg7BUr3labiiHM081BZwMlQqtaZdZNC1o+Q
oBBTyfDwELSOOfikBlLTE13bMB2HC5ETqLrja6KzRPRikcuSL4jv6Z60FKeND37e
Ky13BkqGt+fKAGyY4Lew0q/KHPK043ztGOFENqR/PTuE6h15+LQH6Dlzybu3Fi4+
fAWEIa1JcDNFcoLUIZiDRHGEOAa284/d4RnarX6e8g1WzRNVGoCNm34yWOgQ0k/Q
w3gBhmIIeu9tsAJ7E3OM2UPC38+HZtcLasSgdyT4Uwk6s6D+REUNOvlkzgPH5/c/
3s3cAKVPYmEJ0BmLpc6Dw49uXN24nYQXBeswUla6uacKkKB11zHavRTpY9bf98VM
xU1xXPYxqoRWdDE1rWXo/vWNeXNiQ/JzNYbUYj/xDcg4jO1ltxKhK+KQHwIGYzb3
pouHG8Fp0dHafJiVRd6sdwAN/PavB5OhH0koIRdecfajgx+NCVPIZphW/YXinyl/
tbXKDC8FkJ8uqmiYtMUUVMyYqtqeupnVBPQxDO7JEs+FM7/7dDQNrIeWa7EAv18h
w8qpAN2gPhSrQso+BT+P1lGYdV4xQOkYtVqCYTITq8o9vKsuPsc7npBo2Y7DB6K2
a6q+nnvhfp9a4f1aFOrlVk9yJf1jyLgFyZ2RJFo0qHDM+wtY0pEaH19+wdmhcZR2
36y+H9WTQ0joJOJbUcHfz1gPbXNSanpdmuqybP/TP0O05hG0Lmp/N+x0Iv4MarNV
6Sf7hSQxYEpvjhT2eacc0aP/z46g9pGOfQkHXr+92ZIqPqCmnb0YDi76F6A4Z22q
avyUYClhWv1hTdTd2TTFSX3g2QaBRjJ4en7vVHAVmrUkks56dPu1NXHlsFfLPiLS
VNkTvQFeuCxz4gG3ETLvXJFbIZp4kCSz540SgPHYk9MYFfcq/d+CxRbplh0+kkCy
QUY4CsEC4HpbldNtcVnTJ1jdzYWQOgHK+mpqLpM01GhyUIev5n62COBjUkj7NiUD
EJTJL1oopl/kOSmB+Miwx4EYcXku/5EyJuhGx5x/hau2upTEEByvPqFIuLFzlPr4
xt+hdHB6QFNCXfiUTyoN2MBzU7nphzrDgYdBHfWJlgABq8s3VtJuf03Cxk6iM4BV
P7IW6Yz1lyxaNSoNbTkURemqnhIdJD555i4K2bdnNJg5/BKT2t91qYdkyi+flzhB
ordEb6DEL9p3hZ1BxPrMBDJVZKUE13EIwvb5682+vA/ZCR6XcycVNoVQAw7JdzEY
QtcmH6SCwVOP8GSPlm64XOS1BOdXGtopW2zalj7H9onGz7dd9kKjSiPLshV0sUyj
R1X5/vlGxHjcpzO4AXMvhP+DaE70w1IxKW7gyN2DUG7jvv6ZsUkHPtopxSFH0eIr
qpcV+jIp5Ik9HfLnGYbVm0DCOJy2/FpJm6VgIl8kYo0K0FEhE0jQs+uh5EEdRV2I
bQAk4i8ZmqqW3Vn6yCBK+xK6SgF4GxG7Of1Xnz6YQPhw52tNdD5pozwedKXDNLXm
d26RO2PCBou4PNlMuRjAlSNlacrffEiKVyDpgXVKZVmjmTrUr128mc1cyfM7Avm4
JYhcv0hLMEPC7G6arJE9HGbxKs/5aelXDu35faVzQX8MCJ91adeKGkEEasa3u3HJ
Xr1ngLRTDYzbdmX1GvRURuXA/cygVTZunNR/enamkANAeFXjyCCiZIzuTnc4aLiK
3IBQVEqujRfhbCpwSbfDJRu5P5yhtR8q8VHL9K67b2EibqG1N246kFcchDQlhTCh
0abpNG6Ijl1Mj3cfyVNgIbC5myByipenmtVdB5PwNcmWvr9BikL4diZ1uner6NGU
kDui54W1raGNUN/8/lrWdE0dxephQ5vN868ebPDwRVZKYR79ZFTtvuoebC+TSvvc
lOVsXsrYcjCdRZPn+bcHVJUmHnYFasuRtM4Cun8APNhIjKpDrhAK9bUlHg/vFrje
q6AEz7EQQtM076EW+FN4pqtdiRnP4/mq1pXvOPtPT4O/C/+ENHM1Ao+cSeLc9Mvt
XPDgC/pEBzUREpsmy4VDMwciKDr7gPhvCvGbNdseOxDT/uHAESEUg1P0s2be7WiS
lzI2rLneQcX2e9zTtza4VGY63/P3/jIDhOaRfDw698AccsQGFTuM7Xx+7byvsYPt
P9DYH2kkCrH3efZVaQN4VWMhDW/r9vGlyN1WTF4x+dFdMX99mHA2/dLvJPM0115W
nG4Xh4TjSNNld2rAnJ7RVqVCRToAy6N/u5wD+QO6SvXNTbHVgD7gneze0Yqfvuyn
2gpg6Xu1lZhjDcjVo1Jk4dJxv/3P/9HpA3sHaxuEqYm3bxMQ0PtmLzundF5xGk2T
6Kn3xONL4g0iH3uvcO74o95neX5i5HXGrUqaI6rhmv/J+MVQrA0w+XWBbjXSjNRe
NnOUdRwDvy//YCBAqb6K1wKz1N6Vnp6tbh7Z1YxOhvZ7QJZIijVGTSOijW9c0bqB
q+ytkc9Zz0w6TfRNMl8jjaN5xJdnvzdZ3kFk3NbhkV2RMTQ7iWV4thaXb8URgdYM
8PjT9rak54rHRxY8blYZ0yLsIINXyiSOMxcHi+85iVt0D08+aRXRv8ZhVOQvteEx
PH9Ab1CCflhDuYut7TX7PRIlxmK39W0kS8gZFX/Rcij/X69y1W6bu9n7gmefjEyf
Q4QKIyspVv8U7N93GpdTyJLPupacPDA38RvQKUNHWpGZF5Lv1lLBbitHopZnAlUX
+FtKtglg0r0a+kgo+oa7t5NhF0rmgocgNuEgwSoYbrwyV4/C2sDuSH4pHQEqpMld
pY846COX9v1kXxc780e6dWErrhzJu4uyI0kJBGkNSmtrF4DiLQKjPpYpF5heXK+m
a3a9u3ADX+R6QSVwt6W/1Qu/aznfW3ETQQiXD6mM2bATk6NBLARLIRgmQfN1wl65
nm0FQZuj1qGrqB1Iszm0SS6udh/cPrCrv1SZ0T1U7onjBOR4V41NtDuC3jUQgFZx
GfRMLHa9n6FBBFmSpkFTbvTKEU5/E180t5aC+Y7FJO7fAAAqi3vVA3WLk4w86IHO
0yIiSdGXPcVbyUnYil17aUfZsXx0Przugj4bAooZ6oZ86qHjfC+tassHRc9d6K3i
26m/+HTbzcyZlk+fbmPkvywh7IZnK62szCqDOdlOAgm62B3Y36xv1oxvFCVW4eXc
xzcAmd7xMqJiYNN0PnmGnevKBIex9SpLB3M/myjS2hvjYSsY0jk6pmSL6ADdHfGi
PR53vBhVz2565EKzq5lWdF15oSfLemVZOHs0xvdbQB3JfbqmQROsFjyWbhlcV35G
tj6zYAxWImQWLTSavrEIGGSRMoqSj2ffgao22xWeoBHDfEpX378/dejYUik9Nc51
2wKBYlxrkCR5lmKOgLtPrt1fLfrWc7gqJBFHniUP7Crt/zQVT18i6X0OFkaAdymv
XjPmTGASWueRRXajN6++T4MFEFRQ3WCW7Sgs/p6tOIgPIvUbZOxVgfZ40paDWgvH
JJHQ/d0sNJzRIRG37R+ipCjFJbPnFAl1EFKbFYekks5i7454+nPPEbjZ2RXUGzIb
QLT3RDEHaJAY302dl65Y8Ld9HTVa5ceSYp8o1XKUYimxWstXxXO95+xDMxK3g/QJ
q18ZO/rUjgVjMEHUzf41VBjOAuNdcgXX5zUhPkiRK/dk7GmuaR9nZ+pk7zQr3ajj
z2HpNGoSGvtwNpBoW6/5zJ9SN7PpUl9x+EUog97FcXAphKM0L1pxeCHKaET55FmZ
q5VGtbgHA/kBk7O6P9K3f7JPfKqXTZC2HDhvRa4lk7b0x3ACVDhztLXEQ47d7hxh
yyshx2YE0SiO1PmdVdxFYnU/ySmybxh/ZgEOnoE5vzED9w+1VPcVMCVBgW8FAHzt
hua6S9vLhVKLBjkTLW+lXGkWdh0qGOCGocbpJ52YCuSLQWsJ6X/wP9mGMwDK48qP
IkL38BshJDbFmZ63EdUVZYcGp98AkLwnC4LvVu8qiTVjiC0Hmhlt1b8kh2BswFP3
sHd289oLMArL2IsbFOHecGq3fbzYpbhFH4bwSh9x1nJ8R6sEcQ8+6rBRnHQLIOlq
UrPwTyAugIOIafxKqTERKcrNBpt9OxdBoeTOdQB8G1iVWlJ+giTrwMs9hjl9iZgJ
szFiep6uQHIuKxp+Hm+MaEcI2lYRJe9gP0FrLVaCKJWW4ZpODBtYraMksH60VkiJ
VJU+NM6bq4NWR4SkcmimAISILw2SdvJNyOwCdZ6roLcl2ujp4XcTgnaX2HVrzL2T
2qO2bP6Go40kvOzpLTWyUQDle+k68zEGlQYkABvNr6LYXyxZ208WmZdMkmvEWQhZ
YRqBdsZnFaey0IAgrR7wsklwNsM8md25q+JhxpXxI+TjZfPlJaKOXWBIfScN4uNx
IaCs9atyd/Kv5YDmXojlE7sXaRykwPm3IBAPtuw92UcfyxxVl7IvV0vXAu3/5om2
ewqF4qhWBW9l+namAB/+D4TknciLk4En52cNrQgS1gnMSCz72cy46yQN+ybX91YW
Qp/pG+0xppknNURqwmFz6Uf/aq0sYE30TsZUctoKkQZALU6pQ/SZmvXW7yS17D+l
u5A29vpXWPktR7FbmDDZ18FRhQoX8rz5b/x+Y4HFC18YQIfG5Y2eZWYuCyy/aGkh
3uS8tHKq4bytfSCtEnoy4/g8YsXtRJBHK44/LanOkLjo+N7hB6UyTnEvcG+FM/ha
zA1SiM0ZN2mteptIIJY5cftvXL8D0Pu9vZ+irbpB2I9d0tC4JZNknX+R6l0rngUI
frDvk9/JsvJAnnZ9KnjO58ePQQFPwcDS+yUO0uGKgVr9KtUBZYjmLIKAxwZV3fMR
0qwj4lV0QCOPBPwxotKQYFCMmsn8oe7FOU8q58VDHSKx7nf6TIqFOKnrA+o+xFZn
BAh5kDXeW/4GrGup6dA2D5/nX8LtFGA3t5yaY/dop4+BfRTFt6l3EtuyxgXIbxFZ
//9ErGvurRdrFyEMRMXQi+8AwGETn/G9+TL+7+VMCFwzlIuOS8/EHb/yYsZ6aT5e
rGO7yKMaZ82CetcQKNZiJtiNrVRR02xyMY0ZXcGmfy0GsQdzVHdhYzeRd371kpUC
CFjTmRNxPp7ErBqIEobBmmtOKg6ZedJqDxq/ivfF2KkUL9Sa7Ns4heNUAAy9rwOt
iVWRz1sEY3uLY4DK/VmyA4p/J1/AdwNoGX84rpkxjFwGp9S1MnJ6G2eBPHq8YurU
HSomDcVGjLoj0lF8gDl4BAbo0zV4gi9bJyX13koLQivCP4rCQpXjgsWbmQpQhOEQ
rNg9yMUvh7rOGov4z/ivtbZznHkqYHsXZslnugPzeYATsev44YIJGZXvs5XqQkY4
ljTBATnppW/nWN0yZ3q4suXFhO1mVXgJKoIH6BrM+F+pX7IN8sxOQ33YgX/J5Eiu
FkevIqavD+md2u1Df/VQD71+iwqxXMGyn0lstGN+WEEnH1PcSv2oGimAxOpPCd0D
3CZRW8Oyta/TTo99M5Ddxap6HeHgUI8bAb/xORsea/dPmOIP7HFqvdOFuYjaPSsQ
BazQxcpPumw1Yavw1xkoWUbUyyXcibaNmle9NK+gEKPfMpBmLEMxahYrv4UC+LLD
5ZR8aDGUVm0GlndOdLpm6PMxrQz52mfTshuz5hbXmEkXC6OK7LW3/4h34cVParem
A5RcjYA/01RsF+biti0dIWPFFuKm5dvcq6loCveov2mc7DfEFQAol0HWMF4mDo8d
SSdXY15BbUBsSzDC5F4Q32SWS4kSKAv0iHkiKSHOiOUNSCdIUZCqI9QxSh+qGZWK
6Pm2VMg8n/NNQ+57LG69u7sO5JHcftWQXM89NaS94ZXHffOcY7zhUxiofZpjdbfF
QDabv93UDdq0T9AEiqU6ahE1C2KYBd25htqNuMCeceEs+Q7OZjF1jHOcbCUOLW2S
rMRlr7dTJGhxXN/NQsWNxOwIxYgvV6fHyr2ESSDQJ8fbB7g7I5Ddga+FxP+6TlSA
wokrW8+h2E4ztdHhaMx2TLxjXE4rsy61XY1h8GhTHZ6yMMGeEyMOpHgVUni/9vec
QcaP81AJmOgERM+FE5O1PviuKeEgHUQi6z+DtNB71KfKBFbWyQ/mTalB3oTFmQg6
Q65B5zJbf5qiOysPIyr1ojpfAMmRtBjz90jXyJjwBfSdBf1PGOy9VNKZYiDMN4Mj
dixCiD+Ls6XOXSsk0GGF9kED+C7uI61nzxMZAObQ12MJxdtW7lsmJYtVURuEZksa
+0LbB1tPRcdX7278v8BEO/T5nhNPVMGllFTPL6O3i4iBPKsvZqxq5dc4H0YKxIbr
k97DFl8V7WPQ+z94Dx5PdwyxUliRTc5kQTDaO6nmlSZbEhuXhFUNk0LsbHFzQY3t
kmpWFMgVSPSW5KYY7YScb6ofhgc0oz8oRRzDC0/EGHNeWlACbDz59C6elyOl8HCD
KKC4+CsVlU6eoKw8xQf/P2424pPwo6FW262j+m9I45ISIMWjt4nKtW+MJ88cK29D
rCNXm5vHBDmZJm1F2bL8rcBwA2i25qjReKqzKGNnfJsNczCZ0sdNd1zDPmJBqhlw
eq+14lHkjcS1fRfPuoLa1TpI1BCIuFcjnq95xrR18RIOwEEY5QT2AlbOagv/swi+
spOujVmIMFzzcjhyFO5drpfgQ+LxWA5F6m4AeNIVMxo5MMnxHQ0ys55CiGkPu0LI
KRXWmN5Nq1Kx326VsDzRvQpuAhG+86aErFLgl+zZIoVYE0Q3W2rsIM/c4jO6KJku
IY1bJt6W3uyp4K0yUNN91mIxiKg+diJTnk3zcUOZNQLUe2252jHmlQoxYVCN1Xt3
AfSiuQ2J94L14hcAvQAZtOB7bpoD2htp6BvTlukS721dbeVFKCnx/1t6bgN65BtN
mxOxx7CnCKE0ve/rs07zVyjRm/8OqH6D/udr0ZmL7qWhC7LweoVUR1DqkuSu6llx
9OqbkiIE3J+oO3H934pFBI47K33SwDOI+L87+viiKXOZdIPQXryEBqJkKUGkDQL9
UdOFlS6vy/NWOfLmgMHrzJMhD8tORtcODXeW/ANQ8CyMULA36EspS5PVt1JLhdzd
Xv8TVdC/FFnFVTSiNnV2g3lIJfUHGLbt+9QobDP6oKuYmv+moKaMLy1jGgmayhtv
lcQhkDjyxIRxZt51PvhdavQzKSCi+BKea/GCjziApEw6JDQwzPZBWHXVVwdTEDc5
Li72D4NTnd7WDWqeXBeD0P3KnHzBsDWl9BOlu9Hq0UL424brfys8kvNcN05T14G3
xcUm/6OvscN8r5NHhdGP8AuYGIudhsZld5UgN8O1vOZxUQKEg2562mpeXX1Eerbi
ShGDv5q+AUwxx31veUbKC/LjpukG97MN2QwckoqlO0mcnG6AupWsp3feJR8FIIUL
+4XdXzQDyOURP4ffVe1XWlsAUdtfqn5zOgmT+hUK7/8BF37G2+mrMRZ0bDktQifD
K25QRfG4B5alsr28Nnhe19uM7tTqQqnzhCTkBEtiz9Nw1+A0lW1bp5pkNiAo50F1
Sb4PBVtaleNbDrrLszHB5x3E/PXEgpSK9vqU0RL3d1LWEkYLDSh+DYHtTwNnq1oA
R15zJKA6hvh8QU0uNmgnD/DdJN1X7eg0FVZcxW6B3ptnXtr5MYn7YVuejI9tYQv6
NIgBxQaOYB0d5prdBXoZB7/JxzT5/cSFykz87L0SaTe3GN9QxIZ9q7m2lGGbkHva
U6pYYyff6+uUnEpim2NqT3jDkGfnShqxCdH6MX+3Za3G7JEQP2ywRL7gUsWODFzS
HVfLRl7uao9If2oVU+5lC6uT3t/wEXL55uuIyWubjkkYXNPcGZ537DkSquHLXEU2
6oiFFywIXNFB1O9BvDEV0zVOrNAqxxZW+xtCxtpgmZtTUSbLEI+sG5/24VWUN/Qu
xKFWTVW3xsWlZY7q3TC6dX3YakGkCtczHvbd2YFng+lWIprXJ/7w9kOAEF2CRblS
t7elWhqUjgHU2+t5uvS0xmfyL+Coa+QUGJ59SZWw3OuwyC1ZTv+YiRXHapIzsgNf
A9884zZhNb4o7nrUWgVz1D6iS0Wse228L0yMFn+8Sukulxw3ufthJ/tg1Vj3i+W9
t0pg9YN9efJxVzheqr1BHy7Sa0z0Wzu4MCp9Snz62LonUXcjtCxSkghuh3/QNiQv
2UbcJqT1VdAUKiAHJtVu8Q7kq1yuapyRukmAtYOod7sWqzGj2QvhG8Vggc98+23t
Yo0nLwavkpdDa3nZSfM+3Ax4jeYp8Qh7f+VMziyTZG3MjWLsSLnSufEnR9u7qEWX
v+IxQEVfapRXs/WffNQ7/LxQpM8q6U64T6Sv9CDTl8Sij7Uy/tjCNsutgoq63PKJ
fga6lbPtmF+gkpJUhdz92LugO7Dh+Ikak7WgdsJ76nd7dYNPQYOPCH7T+NMH6J8j
PftSe32tk/AzwSKjMJmy1dXGAG7qI8LjMXqF9lbwqEuhXgLvZb9JsTZdgyAjhJ4z
XgWTC6LA4UsWnEcyZGn7DvC8IDGuMsPq1VsvpIwQhN+SRE7RiOoX2lkfN2dA5jT+
gkPBsQzFh/qZPPS43XakgAigjVWO36KWmfOLywqyr/Q9hBwf41XhLpVCXJwHsgbJ
ER0Ic4yVfftVP9WpH2bmIj/lu1Q1X2dQjCInrLNe/8NmVQq5tFf8h1YPe18AOjXi
wVLfeYeh1Kcg5VMI5BpinuI42qxf+0mV59LWVcmQ0k+oV8djJPgOxXA4xFiNzUxv
QwWMyJmHtKu9QKN8/awzg6mmx0tJO2wtTyEFAJHywwDNkl/IcmCWe5kwMYKitCvl
9tyoQCLGPhNj/0kaqocUqfOFvbu5cys7pOaPQ0QvPrtNoSSyPyBP3YsjrXdzzkM8
QFR1HL4rGG9zpp6vnAXtolkNzB3BYZAec/qZXvZkGWkl+w7JBuWvqyVrnIhZKxvu
uuyoOzxj+kDpPxHxz3cp6YMiMhpgnWVx5duZyepMWMNMzRpufIlAzNk7HFyMFChD
UcxNtfhIaWZKCRjujmLEqs6wL35PvD4HVVjYzM850oqHTVaS+xidl0M2D3QJXi7c
h8mGwycX35jlERuBFs6kBrmB7Y9FH0CWkMQAkzSfjqAx2VeOaxSCc917QamyJ7LD
bjZ9DoIlnQyeHlfcg7tCvUX/jEnnKNqs8CYO9/XXXjUYn8kTi8vlfZK2h7xW+CIy
y0Rp27gTjw8VHZ6A3NAMQ4JnpGQUCEIp6L7cV76F7LUgeYpe0yPVk6TgRQBdZMAo
ONP4hkigekN2lVUd8bRhU4fPmKD+M3WZP5pGtOnnyCkFtA1GvA9XR82BvXjfFqFU
pBe3Oart12us4bCXbU9/9eYB3LTDWXdbD+bhNEAaSYrBZUr7/Wl7cNXQ1+Zq3E6g
bnkOl7hHSbYX3/DtMNH1LUonCCB+sypq1JKYfQSlsp934E71YQPtM2DNQm6W2DZH
johJiGejQjW8Ji2oXNtMc2Rj+ifRiimBinRoN/b1mbl++QLzVlraArfhOENc30Vz
piPCcz5Tpf/6DQiJRO3kPBIwuTDfl0molZuNHluBviAEp2OFhufTZPjy8kWTpe8t
XII2se7WZQip3hzwC7qaT/+F/4RZVowId8mnzeBmUGe82ySJVm1KsxuQW/2q/Iz9
Yeok3Uob1fB6LmAbJzkA6AhmNhvkF88BCuoYVCamtXyZNjc0gmsFEugvMiYRaynQ
clkk9FsqNvwcXvdm4GqfkozCoX65VqbImqZELBjgw3fWdavHhEKzDonNEj7AROD1
7g0uHXc+2k/ewxfk66NNcZNJ16iAI7eKSE6pY3FJIAw5+TAHE7Q+nvoSByDo+wn+
9YgvLogXAxolVut0XX6LUiaCdi7SICH7TRkhmIOsC4yjggBWgzRQ0rdvBWK10GeR
da/Wf1SQnSe5DGaKTg9uvGKiAin7consKNp2LP9owN/5x0mkcuLEngnG2rRHchVP
hdYI5l1Xojgna9fg7RzEQ7AV9yMOVkRutQeBXZbYDidLtU5v0pGyOhOWRPydS40E
jbQlHhbDbphJC4zOPnFRotyeGjo6QIpK4ufCbKHYo5DaxCC3UsIR/GKZ6meEkvPk
1kC70Ged1BW1+zON5O66h2jCmgsOE8Cai6exL1s9yok1Wgl3gP+Lh4d3/+E9pt5W
mH6PBrCsFCzufv6x2K3ukaD46Z5mAqpZ/lg0e1uwlwl0Y1O3hwNkKBMEzrrt+C5e
d5BJbGqPxEiadNgs7ajSyO2xubICpfZ+aqqhyMsszk1LbwiqSnQwx0IXR9CQHikx
1xdntSJ2Vd8fyyVlSUhzi6f+aT3gkLz9JArl7nxORVSjfqpkJEdfC8+E1t8yOJUb
aOqspV48LGFIJO6mweGrBuaWsp/GlS28kElDYBxo4cMzAzOGRJeDCraQKqVTjdjU
tb3PdTRgX5i5HWwcho1ycxH0TAR2kqeNK48aFRXTeLcttLiMYBuZFuxOtsfwNX56
s2HQ+bJ8Uuyo/8MA/FdwERqOBLuMNoC0pbGOZOkGLNBCcqOZdQ+0UyiG+LOwwsrV
k+KUqyqonomZo3uyuVF+rOqtaS908euJpR6bTEGcDF2HF8zhGpAF8YVF1cNONzB0
lImmzuaT36yxKe8JBdBQOvio1ViC4UvUh/6OE+oXb7C0n5FUVgQk6BPwDmdigskG
AjG4WYBfXx4p1eqmmJRJP6A7QMFRoQekpwtW2LJ/MCiHiZRi58mKeztL7ssELZRD
MsfEqv8Yu7P3Y6HoAuu5nVraUP7G27lzUHrGqn134IgBHl5I+XgYAmXiJUbSGhng
O6advZ5+rAiEK5dk28ZYuEFfTUdYatdrWFTJPtrIiPyZEeUTZNR9ZPLteMu7ccU+
xrg5mHJsBzcEhGgI3J01vmvNSa9xdBp+9o29t1VjKpWnC/BR/o9oQOgxe0vI4+HT
+MOCvJvO8FXxxQSqR8e6m0A8iZro6epCA6x+ctQZykLcdTC+dJ2erKPxNIY9GlBK
438O7uedgALvPmiv5336dfX5BZr/kWfo8CWo/TJbFN31UpTqq9ajrqTrIzh/A2dd
jjr6YuK/DP3GgSqPGP28vLdE4AQa4PFppoAkebCmJcOxXAmfob2dpKmlEmZ1vJ0k
UUgJLe1mLWwnZULRZ4IeEKpysn0ksiLq49s38/YWSF0hANj1Fq3z6lrOVVtpytOf
X5t+vKMGTNIj/ggzPYfCh74pcgPNMF0Qsk2sgNeobT9bUwOcuDbHkrHPfVj2j4lK
1KOkAEX60zXLVeDt2vUPSJ0U2OHvsYjVbKz3sY4gSXbfdERutgbsHkKynMDgXWBK
Nzz9BCHNs97nteIvwLzsQnEtoxg/rfzFmifg9GRZUWK6qcMqaGdjeQKFUQ7Lk1Q/
mLyhIShRbr2QsIvw/9USndF5SEE65+nwO8G3V96rd14BrJVl9kfHg0lIIX6VDnCO
WXiruuNeIgCm+5b8Ajhs2eHKH+KD/B2ih7jZCVLBCoBOqddhtm+HCowwNskgsQs+
Xfizew9wbF54/oV2yDBgrqGGeJwnqJCQljxUWO6spA09ozKFIUKtwwBuAiJmIc6+
WBmTMGajZxgjtC8ozwxavPBev2E3i3PNI7QZ/DrO84uJ1qqZtO85lLqW3Gbsuu7P
neT4NtQqxj/tgwOZkmykh58YE3zWBFHg5ObaAGmNkYYpNtP+GDoDZBW7o769kEKZ
B4hv6raN25vmSb0iTVvWP4IjoH9qXt/dN8+gKaGQVeZaXue5rffvsuvWFkHZ63Cg
fxMbIWBtY5NkJavxlcoFGvYuKOrY5gVtmg0on6HLvFxQWqAk7lBArHzFvB6a0KC6
CuAzNBAs7nKaAciG1Wn0yz/YkUGN/vrxr2RcgH7BqSHGEIDEbK7z0xs15a4yxgd8
eukaY4Wje8KuXpZ3PKkd/seCdcx3C9ZwDijb+bcfzVsX1LEhL8plE1+Dx11qGZWg
cU/nj7EyPigtKJKT+3U1xwccbqz4snFsTtY/HiFMw5IGBd1EKmLrUhwEOYugc8Wq
Bh20MfVwFSihwBIVCowDlzo2C8eZgZDd7IpE1a8JsPdfxRZqwJ975Z8xqelBJmt2
HidO12yi0pDR12COnY/5z1hf7X+sZJaVGx5pPwWu/uA0cNyhkJh6Vcvce4YiTb3y
jFV4ajysliA3jAecySTaDag+75CylnBL1B39fI6CBTOiJVY5Q9YCFGzkyEk6Q+8b
N8X11NmAltl7gjGMO4Obrpf5+KJysRSu+e9ZmCu9/1PFam14yNiaVRpbksqzM5U2
aQZ2J7Vx6N9eECZKQZ5COLe5opbSDolbseFkzRo9ZnFTgjOcVnEG5NEKmpF7cHKa
rKwHlZhpcwaxi+Ay4YkwRTJC7gzjdMX2UJI3DFk3AcFYR1doR1ZjhqLIR8KuLqy7
DuwxnQltEjIyH3uWmkGEh/IO2zquYV8W/iQeG8fOS4wsoR3nzSViFRtrh+N87R4G
K5h3zdo6vRySHLdz+qL9AKxoxLlCDBE7i8hgVzvWYg1t+cJjkn5Jo3T+LY+qP/JE
2l9E6BSTi8uXOLO2PfimBuekzzU/a+YDmImz+m6WCtpMBGQW+6IEp7QJZMLwNMdf
DC6AN5AE0PeHbGJjXzuidiEKw2FQvjd0kffB6GWTJ0dzv22dQVtOiW39ltQMW+5r
Pcc+2nJGz0BEoRO6Sx5wfW5fSVLsvxlj7a4ML1qnSqqDfYWp2+3XRitzPzoVWDXj
kIjnVJhgdqdeFpngt4Z2e+ofQHOfidyNcL5JEXiIuE3dTDP96FpS2kRfUTBVkIqV
+S0gZFJMjsGroCBF9cFJeF59eKYTmPDJuNqY/5CVf7z4wFCL+PhnuMxLB5pIPM4F
67X27JgYlbuHp+Amq3Zz8ec13OfGx2bUAeGYSuCEwaVZUGmmbJZv9Pntt/yNtL3p
A5692rZ5ike4uGgEVvqlcYjYlFsITp6wGsS1VOTb/YtNvKRVye/EvWkqx1Q+yCMN
gSPGj8Fo4OZwZRtC8aNCXk48v7mlQAUmDpOfyXSn/S9OfDfGHl2mLrpRf96jWAyM
tJZcNRN9TWClnvaqjR/pye/Ztq6vqzK0ur2wDMpKTo3CKHwv7L1pdj2rrhQt5cYB
Hwb07hE37KW7SXEeIwGL6bB1v9quH+mOU0CEqdBm0GevzzFZMaZMA+trv9Ey4Gbg
qjg2zesxxitu5PY6audOPG8OeKSpDTfy/vmo1FSuwFrZ6ceowHhk+JkQbcFAXJte
AIrzRdhqi6XW/LXQO2l4m63qW1E4V9ZBKdtmu4gdecxk33ltzUtJ53zchbD9P42T
sdwSh3SdyYq82GVoofcSj3iResl4LYSbj4vwjx9riUjbcnkL9AJWwLZBii2//4f0
mkHmCIwo84wc7cqrkTGz4GuPt+QorNFRYPOawXed9pRcXv9SWR9EVlyUQtgYbV4Q
Q9XGQMRCB6xeGJdOBLUsTE1uNy1qUiCnYKF4AzpE/2j0PHBbtrblbk73sYQqWjEA
JoOiPWrh9cksfpGa4TjZlpbKkLD1egctwm5Qw1f1aFwsE9peq9wV327eHcXGLOsQ
T9XKEhHbDvopuGjj7BwldHP8HuUo6Ox90uk5kdBrEbEDHrvDTZ1DXF0+Z5PyGAwF
pBdQJtq3tqnG3033rvQOSHDyeRGR54E58OWj6HqSxGp4NKM4CVJhT7bhsYiWw4YB
mQqRoyfwR1X75a7vy4Jq/KGZ2HE2zHPMNjuVsbpzXONRfl6xg3rGPCRS00PXkJ1O
cvl/1xbzOTtsruE7mCleeZYBGdJu2V4ybDehJRqHrvvNMLn+7uGZsJWwicvEro2E
jpJqhwhobzDyzIwoKoKC9u220fI/OLlV1hMtmtgSJH0BQ4RyRP0CgRHnv+KC/0hc
TYAPcLbSV559WOT7JCNhtS1QcCUaUHNfn1SsxBfrK55+mZu0VbFMWoiOmHFDk21f
0pUVjj9RxagaiRcqVUsR2ENpEIGkKtU3i2l95qqWX9QvFJvGuDzrBGTvHUE+LRNZ
44gipLGjn2g6k7d4Dj0T452OPUKfgFy12j1iJBmiylbELVDi6HiCTyVJV0xGNvo6
xJqNU1mlRiU2irvgAeeHo8SABifzIPFAA90E90Cz2GtDreKilqmEaO7IexE6qnDa
weICJPYVe169RUNiMz9gUd7R+gm1ZXIlC+F0Y2HgoIU0k0cRlOoMygRgNdW9gNrE
FEVsm/pkmQ93YDL3snI1pTzCKuNBtjm/KWEe5VGseXKQn3awXGaWn09ri6kMGH6s
HkKMEGO1KVWs+Y9YLsT+l3NAc/kzhoobJYiiHbghqoORt5FrRV7ageJU9QniGbEo
lXyfEKjYO9iZGI89xA9uYO5+1cL40SAf7mtCtY31lFgKXomIU2AS5JykU14ybpSq
U1HuZ7/iTPeoCCZpW+8WVSt+9hmI79RmBOe0PK40IMKinCO4BaO73QITwtiK7bLR
/+0+h+DBV34lhERvK3gW+IeCxzTOF5XicWfXMBkt+zih3mp0rIUqBLE3btK+v0P6
xkCbML2copdk/scwolgvrpVDwC2+DZh2oRrcfnBdENL6K4NVlxnmlnRnTWbCkIhd
mSIUE/qvnWVXiOl1zMsTXEzWsmW9KZf70qLeLlqZ2Dtzt90ejJlXyR2lGDNdOhWl
hb2CVOMJ9xi4tUg5fC6QGzU7y/60wy5GVR+JFwUOypgjBld75IxPRAhAjqVknnii
KyM1EOft2zbTTl8gxCTSU8+AzbQKV6oR3z272SLN3ESoveCmSDNoRtdRyy+pBFM7
FcOUGFXnW08ii8HaUpoIbZp/S1bNkmduFOxs5bcQbcXKc6mNXY3eK4Bf7eGMvWge
3oL9IUsu7ca31GXwiw6MJaZdZ/4UuBU1MyeHS029Zy4wOGFnfvL0eCwAtgka719G
Tf9yRsbaslpOREIBLum0eW0bO92Y8kPFmF3fhb5dINEJbJs6RfJ8q1SJuZF3j563
4MQ19ny+agcvhJMcK4k5G8sa7yyLUQVGVzxKiS9oRoDB/dkBnqEgv0XdUT65iSil
X+p6Gbqwx4a1fBXqK9af73bG73LI4DAl4dBDTXPgh32pXGtzkrV31RpB9MzRfY4Y
3d48rNuHKMYaIgWy7MT+1JNlhhhpoei3QCK4xLb3Efss9t8uPYr4riH0zHXm2dIz
iH3etebtPIhPI1TWmVSsgxCogTryKaPn18HtfpCesQWcL1FPtAGJ4WUgf8gFWppg
BrtlnEv4YbyYwGwOI8sWrmfLBjbEbtLZrFmjf/awpYmAvsgqrDwy0KqANU6WPNr5
00o7bh+qoSpr1Pv3lnhPqLEKdJUSqFGQjLhFxxAmv9T9euvnkfkpYBegGpA/b7nW
c+GgoYkkm1KqUaWB9YR9M/fD/iTdEjdgZv89HmLQ4w4kex9M+G3fwMZOM0N3UY8t
eAS+czmdpPj67hKULnc2giA6wn9/lNTH61bXcPSTnUXaVNDnrY/4lU98MS5gSQbf
8W4BSFghd3fos+/h5zBSwOT9s0oi92df4uQYk5zDpmhcRqtBVbcosGrPpYrWv0Cm
YGhD5SOOQwrza5pzX5NPKXdSHDB1YmP9UjHpdxzzbKyrJz+llk1BSt+OmRTQSxs7
lcafQH6T//AgUeyMbRLaBIdzs+y7it2sKfyHmRW8iQIyIpsrVgcSlMGaHRqYZAjB
zy3vtWRu7AGVABm7/w69XFCl6jrqSuUb3AGHeRQMlpYk9bF0LBdhrsYdPjiaWFGZ
V+aZGxk9MVQh9v+NQb9ScLuiIkmr5HkaVoxBqfigOeFrQPAzyUdSPgWTzfU37PcH
ULAlLu++jHR/Vvr3H/vicz0hJcwIAO+YwTJ0Gw3qgODN4wTSbwoVLfWAJuj65ae9
oFWaIBsBivQbvPStEBR/RWrdTC34OvpD+C5cY86XkTsHI9KM6Th8EaZqmZsEH11/
X6iRqiMXQ898dk6a1Yvi2PwPNLXnJBFD5hG2EG4emibKM5HsR5gu7aXkjCab/uTn
XS04vFkrhahDT1KIngQzj9MOuxHwj/RkS3m3hjzxLYiA2JSlZxu/uZvFO9/+TSjd
98s9oPqsiGKhR5jOQBh6LDT5CG8ZBl5qSSzFXo3gNpeDpfCG01Bjqw7lIMQWmmI8
WhnwsBGxdBrCrHzm3MHHK0nc2WqBdk0o463nCyzp54wuiHgTYvdPrU+bakScRCdY
hPb8O7t/LWtJ3acSFUmgVqZpHeFkBPir/YqUCYONd//mdKPMqtndMtxqnxNOfb5E
JQP+18BpgMhYV1rW95TglvcsZ3f8VXsu6kN9XGpr7P7QRsuFZaJe/Ogxn/zpYyL9
d4i3qec36IXXAj+FWEMdht8piuw3Q+QtGHEMCTUrkfmFtOWCgKPNr41OTWMXlP44
meqOu/CzWqWac1cw5eaO1DCx38sii7FkFIzLVImQ/Jz2PWlxZT4dLZZS5OMFQpMt
9YeVHN0jm2OsFAKIYRqiyYCGhX6Sp4m1weBYHtNDszq6gZq9QctwX5891PmbZjxk
IrrgxRdhUjOqlSez/EvJrELWDfjkSzzb3Fwp8h7XZbKtEAtcpbWyd0tEuWS5etOi
570Kw/uC69x1JsDTLedUPKMk2llQfrQR4I4fsX9krrqcC6kKphJ5yBEBnDgAOs4a
C6Cj275T97P1ZhZPRS9JcYCCgUUkNJxO55KjSWKGjvlELJnCPYXZm93wsLgwHFI+
sydRQrHDj4o9NI/XNobw/V3Fcgs31gKk6ES5/WgeiVwUTIGGscokx8mBJzfFaBXj
OKVbYjW4AvfEwhTYRvs9ZRGp5sFgs5tsc87vorRGt6egzkvoMKVLuP2y9o5Fpd9O
4+LBrcyciEQyJTIB9Mjfp6ByHrlplpa5Ntxuopo6060C7wxZf1aj6Z0CMKc/9NqB
hS8PXthVHIrrzoajgpFpUc9Sr1eFlFgym2dlh8xbJfdZjXzK3G7ZbZuK4loux/rA
pDG4Cq5jM0S1lewbclnBa1frimcH4dLbkTFeClClFdA+55P91WWYKSkqcLEKswwP
1JI0C5irwDsZdFl5vVVFMS/++GyWKSHb+XG43caZ15j76H78dwuPZL2HrjEU6OLZ
kDQrTaiOJrIvOkLAzcXrTMOFTbvKqmba7RBAXT9f+QV+82hYDGKYG/dgtKw8E/uB
UmuYPmSMwFN57B58pBb2JbDAoYkFXwSQJ1E7zrprm9Ys4giyIlUqLRKNJ5b0CAGT
8SiOS8CelewGeDBiSHZSMBNzrWxxsxfV6XmLF4fBH3sr5UUGNEISfwOw/BbCfR4P
2KVwpbCiEVtkiXksQAHhEwzSRsdZOEeyOKrw6T9W+tnFIFkrXG52BgUaSFPfkP7F
Tg7UrlAYCPNbzqvin6judVYqig8ABPc7WCTvRFBZF8W3OK/AsIHZnJkqQeQ71uCQ
lfBu5S6bHuLQI+DpcM0bzQ459+33SAC7KKjvoa36wuYfiGVZq9em3HE0Kp7MXsNi
K0kQqoaFUQEfpn6Aih6ExCKY9DC2p8XUF8fuGo5tG6hX26DImsOLaWl6ofgMymTA
iMI5KWTWMZv8wQl4ohAcHB48T0oaJtIZfJBfv2oIBBsLD4j9l3nhMNdiqoRsCtnZ
LfOKjxI9H2A39yJNZPN+8sCGM5eYUufnQ3yQoIhUPZnMenDf/kvGaLotl8BnXAKI
a0/LJv8ofarbD87j/FIriWzN8lDHgLkSHiS9bTNsvRXC+MrIkwpnNMZCmEJZYDTQ
X9eIHPjFcu/n8bEGyVXCq8OS5O8w9dAcTDPVXGod0Iip5+ni4kxlzaIWWK+6vnj9
13V/iXHjjLLWPi9oEG84/LYuLD+SIwj5RRr+7IMp68vhOmNPqk077qqu9gAi0090
U2j1g5sFjQlHDZDVxCgVTBoq/biIf2SNNhx/hRyaWfxCT/bNF9pn0ugEOhlPRy0s
MDjRXn5p3oDd/mRL0egV2tXEvoxWa00fX5eEYPqBculhQ6YmtlnaAp9YyLk+UDD3
zADn3ZHEPbwbjMctu7HS+4JTFG8dWfiFwbFawG1vytQAp1HDAfNlo0Ry+n8Wt0uE
UAOZqNDot2hbPQU6Tu92nV0rYxQoP0FyHzxLVSnzpV4IuFBUlMGrjVZU/n2DhvBC
qTQJ2djvtKlF2AUQqWEZENGsyKTuTuRo79ZYmeAS3ygNMaTzU66gD0v39DjbGJHC
sYCzViu8/YIFenuNZs4xq5Oh4PgUctCvbpMrYbs6wOYffk79FMEW3psYtHETdowQ
n0qY1PrM0wbGgbRJMy1PRolbetJm66YFMawMpghtNGx5hOTg0sNCjyYaUcyzeMIA
/qPPnCLRNjs3utaMpQNOXtUTURrHOq6+GqtTdzaZp/lgJXpCyfsuODDgAQYxculW
9iZOdv25E5F4+W3pnnDHu3IDXKloUTFVyjipkmDDQrSGceuLpv433lCYeVI1a/A+
ucL1WQeKRSxBmQooAguaWAD8G20ZUR3fVWGlZTLQrb7LMdbKdSf0jSUQfKGoxQ04
D4S/AoT0XjZOq76lb1Rk1Ep7TWZLUFSPeYv3r3wNNuW/reLWtEPJ94vr9WmDwnR0
3/nSFr3CHcoaw6nGdRLnW4NivmxCAqahEFZccWopTrFvjdcdbkj9AOwc+8Jk2e10
rtS7gtA0hVVSuxTXWdDv2RmUMLiDvGhOZH01Gt1Kf8OeKuMQZYl3S103sk9Kjkxd
MCAxMaJN4jfODvX9pBf4xxNWtSGBBLi5Tvk9re7SY2qHoal+drikXXyyP2mho00i
Urx1Ddf5zmuSQEuMb+EWOzsGKffHG7xg6q0K3nWlIlJE+qhqqT2bwtifn65Gl1Rd
vLD8IkkzuHf0nfwKZkAt/iGXQNgjWQ/c31jVeaPrD8HSWOtsHC9P6F1SeJVfGx5q
ABWKYzLBrFiM4tFLk+NZVW7TKNVLg61gAqv0pvpK6kvoCh9dv8V5blg5VnsEPChI
Zv2QXqWKO7KqE1V/yIm+kozgz9nV89PimxuT9dLaWtomXwuoDEC/aOCvAeeOGqnj
1MTAqomEliZVhQ+kqFiqMGHCMphs00moBBm/ihVE5zSUvRvUUGuCnC3zbJXeDl9y
G88E4mjSqOE87e57viTonrgq1KkA0nhu0Ylwv4EVRCpSy8wd1QWy2+VmNA6ux/OA
L/ArA/2XRH/bsSJuUn3Of3Ql7WkMlxkIduSvKQ9QLIxdJoqQ+HDKTQeBtNd/w8so
+MgIUl8n5jH1e4g+og+B1Q3F/fbMU3jnO8LLkDMAw3t/28qqgHvnlU5Y7RU4sM1W
YrpX6sMV7ZZ1QjTididNN1Ki+x/GVWRoTmMM8eLKBXW/1TTrzPohV2oVIykh1jnB
XeQhuDDCc/ybMczHkESVz35cnQXdSK2R75GUhFp2/UMrWhEfK8pwhhJuwFQT/lOz
nhXCL0tRHBYXMG9KtE/EjdtoImh4c4Ixe/NWHuO8RoybGQoDeBaG8dZVD9LU3UrQ
O6/3D5CJTLYrZhsnOrA8543NyFXdWxuwAm7zTsMA2jLr1d8/8mvZOKS1qmDhfEt9
TgVC/n7UFrrMO9KDDD9Pa57JDxXKMhqc5lfQ18SihSqXBNfzjDMRr1dg4sgHptd1
DStbzDoulTiLeISk7gx9IDoruk0yw7SNY7exUzF1Az0+dlzT4A15x7Q5HH1QRlEc
nHY8bkWOdVQlCZ3wA2wlKkzwfRdwXp5dAVVZbDK53WPdQiiWLE2AkT0FiEBO3Xnj
bVG0zAtD1VOIGJvTVbkqDrE9JRNcsPPabYRD1FpVu5CuD9RP294VP7kBUqlY9L5X
1ciLJj7EAuT88tvjjoEWD9n/SwEgjnL0O07901qfNvZ8ySUCngPd3PyhJTUv56bh
rP2TkJY20UN7FGrM/KhXe7NGhMsPw3UhsOLgCQoq9LBW6EZw6EDAO1G7OVeXTnOT
N0jCH8uqNvCFgZg6IPR9UCOmv1bpR9g6QOxw5uE52kLot3kzYjKjtpMqKvZ6y6p8
pAGJSVt4+LUPRPplIUrSXMWMnhjNB3AMEDRgCMz4s+eoOBjK3fNkSOWypHR4Vdb6
Cyk+9V8Klx09v+rYt7Fbp2g4s0ZlmOGapsnF2dLsXIA6odAoYos/gdkDlNlv3X6p
UUoRC625eHOYkkVXzxWVd3g5o7MJ7fMLGYMCUaI/6c4L3hcAUHUDhbVfQxc9TDGi
xrhPN1uzu8FxldWalGMpHYu+oMXz2Y1V5o2gEcvm55w26fqSjsRGb9px+IfUb/1I
8O89M5ap6cIh/QtzLvwo4I+LZ+StozirRe2Si3Lpjnwdr2YTPPQfhHnr15Z2QSu9
4dArMjJsXwRrwHB8cqbUEdnrQe0aEPrdVZa3MLF7ylvb5wezA7+Pt1EqrfwECy3Y
BX6X/w1VmQkp0DMb66+OH3iod5dr0jl0QfLFYONVkXowoKU9vMlzfKfsHVNzVOJl
gmIZFdzeURcAutyZS8JIA9O0cTzHadn9x//bbFD6Z7xEJxNUtE6tkGLu0vfGckgh
2FBqAUKy6ypdQ23exswqBMD6KNRPC0BwXLK/Jqtq4du8JIxVuMAgUAr6iha0Eitq
Jeoc1hxm4CQoithrWoWxJX0FPGx7N2CObKRJeWxWvvJ906iXSzAL7urSpKMHFbln
Jav8mBDV0PuzkSinczDI2dHDFoM0lpL1dFXYxUbQ2W5lSSfpNuH9YGavHll5qvNC
AE/2EX19WlTi6hGSq3XZHq2lTN/JOEGcafUxmjBlD49aOvTpV4cfJrft0u2js73t
QJEFOf4YlzXqu/yDdaJTm/C9SVAv0AfoYGPXkxr73azh9J1qGWVidxGYKH58VIFE
+R3/GEvvL1rW+Iqsq+WKBwOIJuhI/rXRY5uPKE3Guvk4KcIs/xTs3uo1BSoCkdDc
T005pK3rfHidYeQsfubn8DSIG/d/RVSX2OtvrWg1r3Um0Ab0hLJTAMD0fiMSg+C8
1s7rC1UpNlXb6pzzCry0Frem0x71nvuqJstDTFNTJReVh5ejSGtvig+UVVm3c0gO
eKdSpew+frOg8TJJtSg6WV5WAAw1wFQc4ipZ1R0EE3yPheMpcjK7WuZLGo0Y1yxF
4VSoRrw0y2Bu2h32lhUckSddPzn6XZX7nMhwf9Pnn4C/1dW1KHqqNpg8m1ym1pBg
mPwirv6/us01gwmSch53HJyysjm3xh146lCn4KOnm8lLTpCgYsyC6+pNIwhmuHgG
nP4lTnM1af5MbKtPVoje/yc5SxHRGKZ1VJMYg+3jklxCkz6XtqRAnh60z80giOPo
x1EIHag+XMVNdikt2ZgfjpJX27hHZY5PAzuWz0PLOPvrIOfCyFbfbzU+37hW/zsd
HCKGaNhA6NcGNMWsWwWARUcvmsrQzpuOjWam2weJ+oSgzqc9+SlF4drV9W75wibt
fWGjTXPmr9If/7bzadixlNXAmrBUCTDI0kh6o5c3w1C/zalIFTIshw7TIJK0/Sro
UkYEftA44JClcdmQMRPUK++kDNNUqTlfAkYJVrOSifw5gZ0IherdXmK01CMd2wtj
wPY3aC93zXI+5DzIVozw99oQVRKQ0MyNO+G9NFTcsbif6o7NJ5Nbz8/5M+08Xqa8
8g6BHNIHeRetfCvf52q6mRb0geUwPnDStgO/Kr8ZVZVmXhRNM8rpO4vhXhwDNHt7
TVgswvXKc4vncZnQbxqnSz6o8yMlutyWNFyk10NbljfvfYRVtb77jWRRUx+bTNMb
PCcMk6VI/L+hW1FUNEOUFqnTYpu6r8e5MRKidSSjCBS8Cg6ph2zvi6Q5nBD0k5DO
e1VAXLp6KT+GR3M+RHvb3Cxa1x/gBHR7LR98AO41rzTbTMDGi37GlivyTjTjETgJ
s6vTALCxY2ObbBeOjCNiykmsmEU1h8C2+JoqDdbY7y3V4/8oBneXD0hO6lF3RHic
CcvwY2gwlKi47+WbWBaNSmnpvkX8f0jKeeP/9ywW1tjNyQH8rRWxRZkYLrJN8j9c
vm5q9hte6q++AF8zQtIx90uxwieQYqRo8pyd9EHZNaHIIfAXxSwwuc/d3ENT+/TN
jRyvT78o0E65b6uZBGR6ggi2/IxUmcSbTsnq/5iqukQpSjGEnM2SaIEPlTwu1aR9
3wtUGcBo8b5Y/KyTaBm2iT9QxpYrASrDvAyz36QdfteNLJ4OVd/LDScdWUIbMP6o
pW3AyIxqNeDoUjDuMvPpwQLb8BANLNzRqDFgkcKoTVudWyBX4YsAtBM9wSJHoLuV
i/Rg/Cq9H+nWOMqptLieopu1UNC01QwUA5DdlWndHlSW0LUVEu+19YEoDMlRNfKk
fLuyVJkDhljLXMi0aHmH+VRyP5IWLqpEbQBrLCKX/gNksnEzzevHI2ZLNRH1Dy75
MG+owUYdBXzkbhMeK6OWdS3tH1gVO7WR6ol2bbjEVXTEDAGNVAD1ENeqS+8jF8YT
YLC8RUaDumDbCfTLzVj7Zg3LnI5/HTzP1fWYEBTKuUcJ+qKbfMcBn1RUlV1EwDhu
w+Ind4bTtU3iPN4q2cKX5c+k0Mfx23Yzzcmzu/DfA2Cp4WINntNWjAuxF6YrdZxp
uRD6qexC2pg2m4EBpXkrt6GlxEJ9kuSQhVqFG/JK1dlMTDQs1gskCr0AM7kld6F4
nGwlGdLVgTLe+eopzbENrVHtfZl1/bzFKMLF29NA9xwnGxqkSNuQh96K3WaIRJ5+
Pdg2l1L2njAQCLiYCh05Q6/W3sksCIeNQ2rrslNKhUuleoMo9T51pAIc5krGwngj
tg5KHn5tmPBlPRQDHBxpJomwnRlU1JiSroauJXp/w8HUX9AuP6SuAki+L0iAamhQ
xa/yGb97z0WMEZGyEk1yWeEUY5qRqBsaqsOmIwTJCH8Dh4iLJWu89bL5qo8SZk/Z
hfsVJYIPTw7691MWnFgsGXpJOJzZawwEHbKDC7XqhrvRVsK4VjMDZ4RLMOKxIYHa
bLJFkJ3I+hTtEYk8m9Dw71Jt+apOD9N1f4jWtivZzG4vMuTJbFeOeG+ZplNQvs3V
yjSDFPrbImMQ2XWF5SyWrbLTEoszxq9mg74hFCbyXWV37ovw4iWWSzWTTbbjt+a5
iTOFqMkZCLf3Tn4bMOV4DPd8mDBd5QJ/zQk0k7iP2iiPdZcixyZ4AnDcSnm+sKTf
Eyf/c8wABFej3YC/qthGq6NANtA+PSNnMDsw9nEWvHwTWIcMlwwZxWhUBri06cpm
bkuVoFn9txHpAQmY/DWuzrCO5RewpXquDI3iPxsEkqZIvkSFL4ynFX0AvB2cKysU
XTd0akv+g/NbajCf6UGqU9I8ITA0CP2Hd0nfYG2h5Xj5+u1KQRIYFb86uN3BqoPe
OqEluJJdYITyVd5vRNsPsr3tX9/K+JfOjY0UMr1DCRuED24pRzRk2U/HHSKnznoR
ejNT0SbgB5ArfuTQyLpm4FiEUmTPHx3f9N2i2nznyi+5swg3rZN8lhtpG6TPzMKh
XHTGv1JT3aPdiJLtAWPh1w276TyD74hTKLYQLxEfTE0E+gLWgzYCAetBIDxgv2Y/
zV+8mCz2VY7hJ0kYjwS8hXYa23P2eqIwLZiJ5wF0/7eSmRAtCjH3Tz6EvN0FEdjz
DMCzIwOySf3bGKZFqZTBIUBwYeqaM/f3c8ddgUODd96XNUCbSlTAB1BWmSQSZEFR
FpohBXQULkdO/wt/7nCE4BXbEP8n1aBx67y058+6w5avph9ivnlj/6NhhQCbqpLJ
kls88QKi9eCAoAfmosafzhXZOCuq5Rizc6mJsR4wBxMhm0BQIWernyTzjrNFduML
hBU4HB4s94KpKlQmd9VwYXNHv744SyOqc8469moYqeBWaOZPa/d7ZGDIvO+4sOvv
0NcmkTfW+NwJe/6RwalUEDabe2txlVfuFgH5T1/lfQD9sasp0aoPvW09uHtFi/po
1c/uLg6+CJ4fK2MJAmuTSirAv2VydUN8QCsrmiDyE0W8JxwOXKwoYWWorA5a6ZcR
QeFikEC09n5R64sTqkw4r5MClN5d3WskzZucYCRFQOCCKA21b57j6gDFcI3QDH8/
d1AMnzVHMaQ74YLDrROo9ZqpEinYOT3ndZrOsTpKw8tw+TE+e2HaXU2jQO230+PX
nkGLqJ/FjnAMf6wWUA5+Fu0UZ2kAsQFvYbhbu9t6YUC9zVQCK6DZfPSoC/3+lMLa
w/w+a7WZMtTVJ8TcJouWx7dJ50h4VBnRmErGzFO4vmg6LVYbGwvWUFUNHFXOQD73
I5C9PJos10vGBQRGsZ8QBNPgRN7C5eePFZSCrng5i1NFzaIsTP/yYCs0S4Yw5HYh
ejI11dT7ZRVfuENWliW3vQYO7OtbiXJpLEo3TtZiQPAOSWFEm1u7oiO27I1tqTzM
WOLXxedQqA4lSkepmhHTuVfaJPGQyYFVX7VI3VALlI2FSBuBuSWb2Yhu72S291kG
RxdoMreLOLlIRgR4JxI43Qy3ap5VJneBsZJZ3MGFJGMCtugkneowlVlJY9hKY3XY
j0MQO6sr96/bDPEFiJa6MGsjC58KS+3XxnH03n6t+K7XYfKyZSzkc5LfajZyxp6y
eFOkGZW++GoWmaFfZM2IRa/9/5N1OU2B/N4kU3VDv8n2M75ZUx0DZ0LxU107lKGK
BkgW4ajV51aH/pCxmJaYWhY8WPzVOfyW4G4AGcuCfc8OcI0sEzy9pTVhvbTGI/1K
SmHotxNCAYyrSmSFH+EfXXPqdIgXqrO5wsLO6uzZbyi0UWE30GWb2k7mN0rQZkVe
WwIyIn92LgCeyC029u4boVQsMleM/64UDeTSC6CaYVmbGNvs5AeGGwyXlx2RUqhO
s270uwnKQ3MORWSMuDKac1bVnW+vDmr7eagvFwy0YN3LojmmE5DoVQ+Q1oDMdeFw
CWFgb0eBP/Qli5wA86CoDABgSjEg4IV9UAc7ulBsgdoIGKQKXe32DdHfJPyPuVif
+1ABMLrvjioVIOORGhOUJJ3r05SBJh7F8jPEEMHQkXCzzhXEWD3Qr7DtZ9jn/9Td
cE2TwbA90LmyHXQ6GwtnLD7p/V9qUEZPvMQxZlBsSpDogMwb63vul55rYvdFGVPH
WbpyRhBGeZWkA4578bSI4cH+dcWaRShtZUR1lTV1dTwxI4LGhzV8G2KXB/icZWvo
lpGJBgxOKbTIXZipXWpdiXB4bXjhTrJigeltSAi3u/wRwsfrv4yj06xTia25HXKh
VbumpcxOw2qywTFgd9bDAQbSfJmrjZB8dvZM3niyUzQBxHUxSespzW5RLMCzlw3M
5EnV7bOTztL1qeZe4UnzILKnInkd4eehshi3WN3NfG5z3+OVW0eLpK6IaYxvFoCx
3BOmoUFGfBH6u1QiMmxOusoO5uMaaPIDOq+Hwj6hT3wX/9CvzybAd/U0mk1B3Il1
PZyR4OQC+//t1OPc6b0zRxWKLqZuu0sWSDDdgYX7kuVpEXLMAuNdrohtuEEraSKZ
TpsVkUi6qPJKKDo3EkEzcbrlxL/0JimJT5a+1g/TJ2DXumVjVEt79kMkoRUBnP8s
Vj11T+EOdp8BOyoZ0vtkepk3ieAXd5HqsWuqESSqkBB95bCEC5UemG06981cv1nE
KQsT7nOKkqrHy7grsGfia3mJodAjl4WqhUSFWRsWnCsuRwmPDOk++JnXYBAnhFnd
mGZTioK4IkzhPbcB3dCCGRzng0sy2uTE49r0LTix2C3BbAdOTXHD0eCs1RUrpKMD
SA7CIincae8oblpTvAKTDpHYOOM4bIUJbxTw3gE4uGvwqt+XbXgtXhhLdlOD+z7g
qAhBDzHEximuiOGu0+QcSit2/XnNLRxZwidV6/1LFhLe/F8dLcUViWDlDDLe4jKB
tABgX2ZbPjY20hYRYvRzBoPN9FooGoxFSJ1bUr0NZ7spg3PJKVG7qtMlfXypYwTU
WYTgPgI0K595oTexUcRG5Aqux9HNVYuBKuejfxIgRBWWrqCf/a5rkeyXiDQef9ja
mWLmbG71mBnrljKWvR/vTRMYM8Y3oeEI4Ctu/Cmndu6DxBJorPV7NbseKQpMhi7U
OWVZJdhTGRsxfD+Qqh4Jurs7SuhPdSIzr5clGnJdFxyMWLoXAERZQqQ9yvc3G1Ek
rdPp/2AUJJlX1imYE6arWyVPduNaUl3Th3yA/Kkh/e4c4a0TE6Ve9Ty0Rcr0Qopw
uL4m7IRBd/ag4roWkxWyx4EYTDiqiX8mLavY294/ubUoiRnAk9vFf74R0NFqacHe
PBM3YSM4GwO+HOpqr+xSNaWBc/UXwDppmPYM1Ac0GPJFQ1Mv4moPzWWqyPDYZS7G
q8cFN2Z/nPd3yk3XYQnDasNlXbdca16uWrNXGxvGKbMNipX4xqjO60Qi2reo4oEC
Q0caKsxYuQK2RRL2U8wU0u2wyCV6Xko/9bot+VdKPyS4boaRSWj1XCWYrNw3DnOY
jsfOaA69rrudKLdAK80Mv+ESYDGDDfs7E/DOLxCoOtkwvBQeDCyB6PT5hTkOgKgf
lSuGhG0oB22F1ftyY7uY0yKPuCn4BFNNVM/F0pW0FamuwO/aWTE+0+0gt9lGJgC4
+WGWzDxpCr9/APhIoEGtDjdt2Jue1OsuOChqpJycXUa1VMlkc8kJcv7BQFz2FAUM
YijI/wGusaGOvvs4vJKjwGyBQIj86XWmuIAbBGd3yHj2sRHEr0BofYO7dLjFOBe9
sghiZD/lw2H0gxRpR9Yej9K980c4B+DZ6rVOg/iUh9sto/NcHGyp9KTQSjMAKzQm
nnqqMa2CclGNt1QpEmevC5Tb7cTbhJ8ZREzqCATKcgMW5MbLQHOGKERBGMT/PdjS
t84HWeIuyeQ2De1BIZN6ArdbagnEcMM2Ew3rET11YjCPWAlsXqxrQGY1UT9NPN40
bhaTeqq9zfj8Fe1TATzVBPH20Rv2gz+ZWJCgqZRkCDwHf6LixyCBvDq3YskkKxeE
Cmj8w8M9hlQtEbh5ObYW6HMKX5I+90xGYsjhtbU8f2sCRqVdCD8r09Q2qWU8u1bZ
T+eFQbFwHz+6U58VtvSTRX2saa5LKF0Z6+eM41HTYt+FyVEdxDuBHw9IV5t+rXXn
bcO/yVmmwRNA3T/tV2rAFllvOJDBvEnNH8MCms1GQ35hS9ZTzn1u28wof/lYvAr8
Rur7hgbZzQCDeRATwWrFS4xTOPR42iVDHdAqTVdZUkYgJcyUeeJ4LzxKhadEfECS
o9SmBYY6OwYBIe6zn4TtFVxMcx9mFU1sYTsv+FCH0BwNgbDmY4LtiKKgO9NJWb/N
eurluORgPJ1HKkZ3x5UavtJz+2vbjX/4EDR/I+gJmUs/u374RzWHopwmgdrB3IyW
n0xhkiLoTPYvPYbc7PwHNkMj2ixtlGomrvOYWmHC9O7aerZuWVbdy6tSy3MpyYpN
Mb3kPfrBhuT9w1w95HDeYqTs0XoBr97/4ZMEp3VwV54IKJi13u8gzaPS5MNt1MQK
+eZvbyLK2u7ZVtjVQY4e+vLcdtfYwKoFtwvKjRLh46zMsDmsgOagkiZ6FPbKUmKr
kuC9+xZ+TC8ZRibelODFXhzWbfBafOQQGO7a7w2t05hb7ZYvm3+9CMJWBVegCgsi
UtnsNsViT5zB7gEnkrhmZyxxYk8wNDKdn3vrHUqp3xdAiHOF0A1dtN60Q1u8Yhwn
ZxAk5hdyit1t2+66CEksp+EPSu1jEkY6i4yCaCn1dyLRaUW3phu3QayN5Ap5X2sr
ghQuk/FsnUiwQP101Eupy+hxNR4dQSYSOoE2UstTrFsfQqw7EXmZKSvny1xUMGOK
5YQf6OUUVDOr15n3UxLfU3cnti0bnSWTIiHN9D/yzZGisG7sCx8peSGprwy+oZLm
wVjqUzQEWZ7GFdJcc1IpPHTjwGCoLRR5WjM5DumxTgejOH+80l7PDUjB7ApY+OOt
JppfehR03Ln/0T/0HDv4JAWN4JWRog5mPnYQ6KSZv+tErcLCJZp3BOAZlmj9G8l0
KxwjAjhNyrZOHd3jw+tAu/XgKq2R9+lUEAnRK8vjc+BcrKWTmRBEF76DXlNLr7T5
k5zFQdk1bq/xmwfQyKgNKf3QTUf8hr05ydh9XUF8Fv5h0oAN/zkphbAqlGE/VwFN
Ot8W22RhofxpA9xIOFJpgypui5DxwwTAHmkU767iFeKovrHy76UVO4Vy/4LO5tNb
9hW0lXkZs5A4VrCeePXsQLkjff3oVkHVkcnaYZPQZGUlxVr8aoF3Cl1VnHjktMAQ
3hvj3UREW45GZEkobiIAMYiPEZL9EXqx9XpwiQGBql/sC5bEVqw1+b4ymkKS2mF/
LLxr8ZnhMOQHklT4476fCRWdpOMxq5WdeDPxyNlIpRhiS6CGuNjBw/zrpzubVT0F
yC9rnUXLL5bLa/1LWoW9TOSV55VvxoWHVe82xxV2pcfecD6L9w77tvuUM4eJgfqq
XEdgpC++mjyqB+RStp7MNlg53tDK7XmkCjIGd6Iv0UH5CuEPBPoxzeWoDhTLNnry
t+9qdkw94i/tZoB43Tu6CgJq0GTjhq8SHTPbIIU9N3+ZZugABvW+NR4WyezNWR17
SdDXD+2SUEkJvSoHXVDI8qk/fMY3rSAg8a27BN3AtpWA6SpFfYvGLPTxD5u+tb5B
6brbY2Hm5m95imm05bwweO+Go5+xFNWZcH6UzwGDjP8HTaHGV7h/qTEbE+gZi13Z
NrqTVYFgPl8SLC9F9IUBrT0/Il8zqt2gomhbFbxZ6dz6UJC7ZTxSP46Yof5p/7tU
MVO9XLirWLlflB8YX7xIE6rUhV1QvfFYUZ3rRMGiqKpnG3TkJzm3SQ01EMPPAWhx
whKHkFWDLdSo0OFFqJcM2+FJThQS+ZHahLCdmP3ffu89mO1oi9AxhjANnR8PqZlG
geSj2CRf0eXyOySX3vlPmrjm0Q5az00bJkCedMJtiQzuBdwOXzA8cC8cXp1qmbxy
MkkxD91FJsyAy7lJK9ZUb3JK+UIdKNSdAUdpD5qkrH1UEIRc/gqFvKby/kpwm5HZ
Fo3GJgoOWRT4F6L1R96h9YcQtjWqetroQDqJxkU3PVDxFMu3NpDFCZ5ThUTncx2Z
WNYnA3OyIDSgJFeeMv5kjcMoG8goutTDMdrBa1K+ZNm+QSeF3LLawSYdiv64CNWv
NEHj1UPVzZ4SQtdCZuWech5osvr9DPzv60H0SFLxdd0h9NQv57o5dwJLTOMFnmPW
gs30w6ec5vnUE7sjMo0TFW2F6yBa1y9rSbiEXAthaHVCMMB52ssvpP1HHAJpZiTw
IQm7et/fxm9S2wwjVof3cCnvQb1G5DR1kgBacrL3AIfzXbsFYZWNMVCcVlVlM/i6
RSp+PH4iIFy9RefX5PDBlIBFF/obcloaOKNptB/V/96UvlZI8BpNsC6FWo5ebhC8
KtVXlbUAqtkxCzgf3xEmTJAw2/ixO5K0VJC8F7dcNTw5Vopva0wA8KxwIYJieaq1
GW+JryhqY2+gQdJWivVxfnq6ixrEnGsU7n/NrtRU8mkpwewABJErvhuadTa9o2ta
xxW3DpO8ddA/EoZBQktREFAckiFQjx6q5OrbU6bbr1q/Iz0z8NHtKL+UJ1ytlGZs
mXqrD+xRXe2Axow490a1xfI83qYQeuv62PiS3t75WCbsncxPQ0onXEgU2/AOOLml
yCmVQS607ZV3w7q/xu38ZHzJOSO7p2+hghNd7u7aCWs49mPtZaaQJwKKrh5ItrYW
Xvyr9vieTcevox1mlruvyuLniGsaR5bXPpUtcQ7K1abCsCDXFzErMkrCtUrD2u9X
UQA4lixpq1eANB3zSycesHDaH+b+Os2kvVyeVkUheEVBYM8/0WL4A3VWnIvyzBYo
exV3lKAEZ4fj59/1j5l7Vg9I74+4+Q5CVgJcDkeuQuE8HO8sj3xJwrZUY3/16pRT
GocOUG9QzxvbNvEbNa1XL4S5CZMPA74zSFRdwKURUETLCE3gUTeQHiJOBEwMIqbX
PtjIJCd3gYzMx+y53bUD046vGSO2DsI53JPWKovjR61crI6PwEEu6LoQKGpQBuF9
9ciu0bUUrYBMKM4xmlfzCA/7sktAw8LM+9yOhqV47+QSdQcunkqPe3xBuMFIIIgz
e9PJUJRhJB8Hde6NOBOpUYvBuO+RuBweH0//niavqHkBoTcb2LbEQ7lMNvUCx8Da
TJY8Tq7ocFOAFDOQUOIMopy0vw0M/FT9HgGvl9hBWa3d1XdaCb9dt3DKAfdAUj63
zIAZr4VaTzRRr0AgKbm5ziqALuH1jJkKVZHZg8Av5Y3GzEiXYYGJDSKUqlWdTYU2
v0Joa308BuP0YUeOFNCqJ3V4Q2mZJ5Tpb0dByzKKWp+TxsrGqyz+Tqor2XGAfGCo
o0YvabarfcgcpNZCI6DZoYjPbtAtlvzNqtJv/rNYtmM9I9ajrkrRE4Vsk05cnG0O
uFl4oP8w5WSYhWsm4RaBa8Q3s3P0eG0tY7lKNiskyRGj+Np56AlbeGTXpSxD/2Vc
TblRzFYbD0koV65GKGcVV7JdeVpxxUUhPLmiyy76nv5Wm5isRMGxH+g8ONJZ5ZTT
4zYslM0QIepEStiQ76wKp3ArF3FkL9prqBdGdEIYPkvk5Zw0Nf+rkNJaDgG8Ycu4
OccrLZ0PoI4B3NEBQlxbJjodt1Pna2qgMWV4WwzU41/F4SBA+mSO5cVdnyus1XNQ
LszpaxUQZqEX6QMFj0dhxOAe4Fv12g/jsDaPb1hKUpYUcjW+f6Xlq/F+Sh+2seh4
A66OPhSAXbrhK8vzYJ7BIit52hddEK9hyQMzMH2JBf/M4bYzCIl2U/MVZZy5rsbu
aAURZkvg2MiVz+73ns2ZjbFQf5ro8ZlGAb6PYAlAmAqkuXD6wdelsm8trnKzfbfY
omHq108U2UIqOOczPAssaLaAlQIEKVd+bUQGcy58EF6sJ3kMys7xchpfTtanE58m
ez1cRhUoLbCv9B4hHDgOjf7FAIQ1srniLgZ+7C0XJ2sQjegSmwFrBqHduF/V8Qd1
93P4PsyAycBxhypZ9uA1+V8bMj3SVgdeG7Pdt+kOAPdNoI8mQMco52RGVNGXAz22
WnCnd3B/TCcXxZRrQmaXJPjqlVCvLcusRa8g0lMKZWV1E3txqVaAZeHHxSmNMMkz
fKudfLDkKX3Y5H9iPnqcig7e2Mo1ULHXkxUeh2Mf4G/plxgPYoCSg7SIjuQNQKD+
HpET20jqq2+Z9+2HC4BrZ3DXj0XwAgadVYv+L2Gdi4M6wCIOW5l8qhdX1K9fdQLr
GArUWSyceNRGeULwZaul9nPVNLD+S8mx8CkiSc7ruOc28ACDtmw2Krxs1FARIwak
uWhauZ7as/XgXSStynPglp6irdlKFLzeq/yQqykC20H5/6d0sS24VgN4+ZmHeyZK
b7NpsHLCFj//UbkY3p8V+45F040e1f/yLLG9OIGu+DJztElDmaxdXps/pBJ8bEmC
eDHckzM5IRJlSYADEo9JL4tME9pzF+ebYPU5g+tklvT/aN9DISlBaHxS/ifi4mev
gEdnSwq3CzbpMKqU28+9rMAN/3cz9VyzJ+Fj2qqQpMC+kV3vUkfo+K7UYekdzSBK
L15zVktxdCjWSoxF8MkSlsZZRgiVyTg79R8WkTVNH54vg8aF7XK9YpohqJylnoxy
wscpqFVG6ByiBNOohNIj8Ts37CTa00oO4KRngMy7xzPCvxhwIovBkI8IjkTi/+jT
LmZpdJQfa2PkajaXxm5gRxX/umiAblrD2alF6U6YjYhDT4UCI3IZFY8yO/DNQo0o
1ek6ekvPUkwGnZ4J6u537A/r7SUZWE8e8JHOIuIyf1RUsmicGq3qerr/Ho3f71d7
xCwWH5tVDM94oswLB8TAcYvW3FdLoJeb1597TEoi65FSdtHKuC8dOugTeovsChVc
TEkJ3AvEyI4z7QoWwzcqMxZdUs5i1xDexrVuRsd/784Iumm7L6om6ODfpVtQQIVU
M9/JDuUMcq3BOye9jZsiaxu7+O1j3oplxH9f5eagDsf6ZJihGeI1AF3oh5VL2sPQ
0GuF/fGqxK/lFJvWn3Wf9jOKUSK96uctsrXOOvo51EgcnkzxFK2xtohO6/UHg6Je
1/tfw+eltOgze4JT6xQnBTMPstG3EdLlq9l/CQWZ3POljJpwWmfQnAgwxN/hEO+1
1wKfk6ANP+bRzkeFTUAcVir1w0oYAEhofGajwd9wAEtsWZjLPhRaKW4RMCUGYRau
6YHqBByoyYBF5KN6T/Ga3AohlTZGq178mlbLr94W/aCBiyNjxVTKhNEoDIFHHAQ0
swkcBdoH22lK6pdNrxUUGIwf3ibEqfTB+YRNOT5CsFzoCnIkuYHndl6Rgnn3q7J7
V/K5060xRSos8JYpKkpftkkXmApJfVupd2UTLP+ozn+q5kk6mFat1GAEP3iHhDWR
SnDThDCYzOWsSL57s1ZKSZ/S+yANmcMBGtC7huTjHB8gCF3VWGIpo5fC0o+ad8As
rOTuTf2NQ5T0OxPW8rXPRV6brnaIl78bMRrY1E8BtzSXXkr9TEwyO4eeUmlCuk+H
7JmztaCO2Iuauf9Dsz9lNMDdYVgg0UcRPyffs+z3VfafVa3jPpovPyf2GvL5Q64s
CvjUNjHG5//QU/Km6Ym2LMQhufdLea+PsdpT/oclt62FmggakhNCN15RaXdyr0TZ
le38YgpwaGmNtexS8j3mkASinx7lErPRSjQKbcV4vYxCRg3gjEkIxedGVOcFi8pA
XyV8GERIitwlHZuXuCfCImXHaeL4s1vFTEa3rRGwCWQywD4wB48L9d/QB/aK7/Lb
S311E8KxymxQlzPvARuwMo08VTEDhHsGzfGQsgcQMHhty/glexCbg96HpZO1D1Wr
Rv3mY+K2/tONVzyBE6q/jwVlLuXGc/sQHn1UWs+bxc+XOwn2yRD817tvG/F6i3cO
R3Ml26Qk0JetBilXumBblYfJqSSl909JQFKgqZ+VsCudmvi+EijJBmK819+Cbbze
ZqtTK0/uc1QJJT1YhDWfUoWpIlJtT6krofeOEfaRjvrJOXOcvRchtWWCYd7ZSsKK
MCrvL/bQi9pwx4tYpf71noTAx+lf+GNyxiduFgBHdOzICl5mKuETR2I/B3lZuw8N
IlkTCqesJ/WGzGQS4F1hrY17SMhqXrxLGrpLcZV37t8qIwx57pSPtdVtd641wEIL
BDQX5WF2M2H9SDcvE5cYdXMZsE5Fsm83hnDOWHxE+gXVza7SbUDxMZiCkXIgvJV7
1seCbgo9yivcipu/Vp1IUaQQ+JQle1SPongJ45Suz6tddPJA1dOGr3Qdxthx31xn
+SR6fDmWjfPyLieGDI6jBTPOzvYxhuC/Nro5EXd6ZTOi/a34798nXXtgFbO9FspC
e5v/8PWx4JATv4+Q0z9kuTALXFa2aZ52YSlPXAwhnSd54fuss/3kTpwuTWw0f5cy
z/ApGybrg7P+OrG2BebunZ/3xtGJWcwlnC8IyHKETgqKrRdTjOaMywUS62bwsKVX
BQPEl1RetlSwQJmPz+QFlxv2xMqobcpgz1l6qOE/QKOuMSpK4CJyaQ1/JnQ3amBW
wY3EJLUICGx2o0nlQ3DNXFHdzzZIEkbfpxGIXAQDhz4GsBlH0aNFqmxyE1vlpIyt
N4lPmMIErcgJVD+M3AJnGe6k6kgGM4UVJi05jOQ0YjQlF5oIC3KHF808jOKX7YCM
aUY7Cz22y2ayKOTZG3zpZZaueOiOcGxDD8YB7yQDWysDGlxHzy4SddR66I1lnElP
mS63zLx2J09c80hUj3SsDuk5XZq9V+uo02XyymeKbCxGlZWZIYoZncd67q6e+IoK
G17RH+yss3iUkRNBL+EjbBMZIkjtWpAHYUqakuzd+PGFcYE0fVFe5qvefrh7jGoy
qqa5QGRggiUgasSynND8Pg1Ig4o/JlR1gh7UkdQcfTSdlr8285BHxYM9WzYRclhy
eOC8izgC7iPS3x4wUHUvEQ6v5E2VBCdKL15umD14lqTjoFFz152lsO6XzBCunyJ2
sylAMul9vTetOx+lJzmM8sUSoguIJjVwf66yqmDNBa8K9jTtssZ8gDzcP6iYcb5o
VGV3l7/3SrKJvXvkY78ODG+lz0kY9rd1dettEv+yjvJQWtJtEjN59fLmwu0WfYtL
5pKfuNWcWeWCg20s9KVERQo6PaAcwj51fNE2p/4mbXmc9TVxy1JxF4zvuuRNwJW6
2jO/fufW1hBbr895jqMUd5SANpuLxKIbxW1ItoAioEezda4Xd+hzHnx4ruAVsAr+
AmuLVIPQC0W2cQKEB8wfzOhtEye6aTevAiwr9oLgHr6blK4OXUrblXOkTdHrjyEw
I9+Iccw0JBKMCyhEk5Obxix6vLtbivgXuNU5HwAPQ++ZBjAYB5E7hyS29X01wBih
rPtUXr6K7CnpWm+gMFuq9l/oINoMXKRgVZBuc/QNwcGYlWvNVWgJehpteE8hkrxA
Sc25sbPdXr8XdP0DwLKBPG8gpXPVHxFnKzfEXAy3Pw49zVzXp7GvkkBnHC+2ZM0n
LHXRLmi50xVLrQIaqgVay9RDO3mN4cIiZW6jxcDyDo6jjv0S/jX3g0EuHnGfmyx8
Qtc32ypwLxea8WJhze4IYfApuhbye+bb9h0ck52ZFC8QkgrtLkI86QCGivcfeVBX
52++pqe2trFWVyY9fbt3+irrS/PVhxmDQVey8BNYouaOpPicnMmgavaqnD6gaJHO
klw2p7OfEamC5ZA8xZPoeWvTT3Sdc+IAVOAOx0u0Vx7JRhMuPRAAxwkFdHAJFE/l
QWfCw85+up4IpyoteRkIq0SDq+5NiIylns3Ome7az36HqBt05Inat9LVzhohDmMV
kSrJwIWyBxyZ8LdZj8MMruO1l6PLDqkLtke+2pJ+r4GoROANozwpJk47m35O7SbO
zuRt0gRjSxE3RefqeD+I7iYEqjG+mNyutrVYwi4m2RXPzxzuB0ddMUIwl4RkVrF7
ch22yqRwv4mCgL3aaS3E434j9QmUCZpdZ0Ba7ow9/Mj4h+iRAoDf+m8dtqJO8r/d
TbGYT+2n8qeZAAfHenzNQQGfkkVlw2wbgz5xqViVfUksfhziNMUK2HOFh0f8qfec
QW6LR84W/GmFzAFIBnytfDe/2VY6HUZ2HutxREfU0Iu80M1a49L719eryQyuXLSL
mchHugqoBDZ3VS442sGCsQULGAa0MpiyvRaa5xtWB8Q3mKfE5D8BeLNJu+R8pfMI
8ObsBx1PwHjEfWhFTNLEoGNsuknmL8q/TdR3UyGvG103xxbwchyqri2kUvlu5XLJ
g8rlfv/vHFyEsN1pvTnghBTzyxTt0cjBqheLN0utB+k7Dz8CBD8EHt4PXVSYZQtG
PaABxzzBUjjGuaHYF1nBTTygRypCDY5Laqoy5GGBlc60LJCq3kGNoF1ie99jT+GS
TnZeLOcsKQU44/BAKYOi6EX4lHhQdk6LFMW4N+4rs1l1m5xe0nwYjU7ZXKSQqp7i
VW4d7jJLayZarlNBpSH6i03+43h2XVFJzIsaP0odvizRrYbZzkBdhLCBKPNtLsE+
8bGHMgwviRDud9pbaRRDm4V+kHCNz0hnwcrcCPPP3s1B0QMo6pbaElhuD8fOPEiz
vIm12I4mFnE49q/CZqPaCJIxM1mqx80gKot7A2RKCZWu8TZp+BnLu7JlddeLWmv9
fKh6PgrtAyGbCFKcSFwn2eM32XBSTllTU8PFIREtNX8h5BdxN/4BskB9Gcakg08l
/C2i9umYXSJF3eXjgIA/CgTJVedIZCpNqPUTMmnGeDxc8wJKA+hBC7ARRaYcHE0L
91L39BTXScVHQbuUkDqmmYAyhy7Axzwfjb5ExdjW47HyUYagd5jTdSRV36osQEnq
sVlCp5CEaifrjX7woV736wIZuu6x95t3Ixf38TVrh/aSNVU8NQ2IyU8dEePR1wBY
fsQ7FG0SzKn8tA5iBEgiT3nQTSIOCmFqhDS/sFHMW56J4NroCj6Onl5tGmJrHv6E
gNSYnN+gDFcr9kSoyxBMhf09VIpVT0FaaQyQDtHZUd0qILck7xp91vIzQS12MCWq
FyCH26r3PqWNR957Qnf2sMtqPzhXP5VQ80uUnDDVsHuOHbMWe+d8ioEEZtG9BVO7
SdKEKEyBfglxrlxpireq4DWi0nuXnpIvtntUJvjOeRdoGvxzZxu3GrQkI7wL3B82
USBmN+LbcrHv9MuVFXWXUU+SAK36n8isBo6FnmNb2h2QEAsBOz4DBIq/lwUjYTmF
fAJTP8O9Md+8DVht+ercyQIs3e6pqFB7Vo1E9JNDLdVQuDwP6PSi1mHiM1Ipkzi7
T/a3lyqAamoGsjEtV1KfuxgpHlbolOzgj9fUa2MXDMadf8X9xBfWZxBUvh9gP4Na
2Ob17jHRAYadtrGckC4oRpfbJeiXIH/UmcYesWsxvUSix9dGj5Xv9A64our9+FDA
jU3+RuJtsKTz7ijHMOSmFUG5RHvKAI/iB9/Q5vCVi+W+O8ziC3grHLqvCTjTpD4c
1ZNegbeN/UCqaOzRz/yWZzGa5Ac6Klv7/eeBHo89eO67cDXQiN7/FqC7CNswK7w0
SJDAPFH/qTyDb7qOklLsHZw+lWYtuE1WGQaKiIs+fFN7hYA1bXEzDmcMIG9K3jKM
gDmKfDZanpcpEADJwFndhDmKkiGcy/897mgxUOplIzn7sgLlLv2+s52oJFmHlWiO
ejL9ail3tezYDbB1FAKCFoXTr2LZcETR7ozHGrhq42TV+6BE6csNBi0+w5XKZzF+
kJc1GPezed0Kyy7i3gWu35MPlNu57iWZYxykBg5paeLfMdcjQ8uN51R48Slhqx50
RbtJgJifJ/PeEqsy7NW0/nJy3j2Yr/CeE72+YBV10+aXEJImh2hBdfi9kjcOjIV2
p6ISFMV8lCv8jEB6dk19/1vDIcACVyObSqftuqaVEtNDMV/laAjaqBCQrCY8zzQB
rPTjegrS9p77mJ6NyEDzSGSzXfLor/s0OHeqykCHEUwOZnFO4+M3GwQd5Fd54gW9
7MSjhN0FNbG7HD2Cn0SmcjLklylr62xGr9M86IeDOxSDheBEqmWnitq0HTCNnqUw
NRkn4KuZoAe47WWJpHC7Cm1bk145m086/XrXGuk50XHeI70JUYvWakGj5IYf/G0d
ueMuUrOPanV8Zon5sU6KQ0fEXebb+WOXEsnoozo6b2xQZrnpKkDfXxxObuW51T6f
Q8yhxDn/rtl70SFToCpXeAs0SUrKJIV2N0/5aBUhC7qs/W99Zahj40+8D8BovIxC
VMgh/TZUzi/D09bStLhQQEh/+FdcndTde1wg2DccnKHMJqviN+WUNwPC89IP2Ov4
VyrsB3jKEQW2tEr6vhBTo8WrwwAvsG5BFpumUqK1YXf7ZwkQv6+lxlVQ7bf/IAEx
6PE4OVuEAxuHW9CWpOF+uAuPGrLv7QwgVuu5x8Tgs7dweU2cMRs9t9IxqG2dzn9n
ECd7khaGwv2L4sb6Gee5ruN5EAluQyhlusZvIm5NpU3drCXbeaPzXe7iHOcnf1oU
EVWWNh/2aDBYLjlLAZyGpjDVARMj+eLjxyD46io2MOf89W6ZgBxQrgJT0yxE5U2F
gGaZxZJfEiO+6ZZXezsWMhZU32MnicPz5J3xJKI3yS7Qu4PL8p/uGt8wZZSm5Vf8
TH8fRcjuzqrzeTePOMMujNZKqRTjyKUNPpTGgSHjUuT9znVxGToROHUUHP/urOrQ
jBPnt5q7Bz7xboq6Zw9Z2KupJvfgxugM7kRMxmMPaXKbfywjMIk4tAuwn/u/qjoc
BmAklzcRytH12Ocx6U/vt7gR2hMS+7HoGy7Iu2glCRjOIhOrcu3SIkTWpndK3An4
qkWZCcfgT73LE3E2EoNAkuXoftpunD5J5v5Bt7PFm/iMPd6wSSLLJ4DCW9QEyzdK
N6boT42bYk3ZriKtFnNq/LBqcR9lSVDU18i8Ljps5ZoNnvxG6P8dPpLTPstkPxpf
hyle/zauyBrbqLMJmOuVA8cAdReV4OglEIj/qCjRs7GiuTVc2NICakQohPxW/rvM
Mg9OqwDM5PxlTx853avX7Fi1Ts5gVTAvHKMPLWiSt2+oCBMNv8vfCIjVDxHhnUwB
g/unmc0gVg23sZkt1kEMZ/6hUfD9ImrE7YPe38ojc5+iyr0e2qyP+p7+OzRfF378
sGBjJc7FBdYQKK8fvWVY1OOMXlZgv0FI7BSEWJPzSk82eo/TFkmYmlfuSPemo7aO
ozom4V83egSH56+LzlktnIXmrFWKGlHq7h6MdjD2NyUt1/STD9msiLuEKV0nnKal
qNAlU7bAyvIeDPDOy61I0wBXMkRq27txuxrl8tVqolLQwgth18wEX5fZ6x1b3Exa
fpbz/EfahGg6CGkcOM9vvTZ0hUs8Glei62o2usj0T6SSAq3hiAL/Eo2c80sHYbWo
QJiO22O8D6gy4ihHDV4RWrDZwNut6CgMttIgySp/gYeKHQAcgODlpHi4xnNYCbja
VTLTVa2VieM/4xAa/GG+gm7qlP4X/dAR6eG2vFqD9kLX3mXtNnllcGBs0xE5bajU
0RrnHHBjgmdYFjnRM96wurNCmsCwweAlTEFAIfWJcthnX4jrJXHNCnRG4i43nc2X
eMRFXnyLD3gX+WWUnR4vUU8C/iiQb508MtFgDUniE60eQO130zVg78RLhGAm0NLu
wi+CQxuj4shkN0J27ucUTx2Q7O2rZotuLNhYsGIn3S0VQF9NLIyHdbuwzgjxIgTk
iEDIFsIWayjDOU9mogVPwUwbFCma074Ft1wgJA8QhzC8tBIVfqubYWmI+jo7KB67
uWpWr7wmn0ZaX6rJOMt84lYLjPPJkMTk2mvQO57oCVSPPyVWuMm4H76vuHvl/Ejm
PE9EHLtp2/kBmfincunJTod/fRtluXst3lGGUCx//gCophvyxF28ogtFGtXO5657
4T5hbtbaRXGUcNLGRV0b0G9A/wj2OGvig8uS4f6nlTmmfv9sKXso5LqW234a/owl
yzOiSxYW4cDQ6ZxRZpZTNQkY4VasM+ZRq1No8YEJcoXJHSRdo0BGu4nj1ct++QbO
8FwtizEux7bZnUAStFfBYrXBsWBUqVMCiEZuV1c9ffgR+ZMnkO5KyMPb0cg6NofN
Vnj7zUgpBonKKmlANovsfUnTEDjpVEEfh5UBWtNL7JAc5lFrUFmd4nKLqmj2NmFi
tVIS6NO93UpeNIueG4wS11PpBECklyTxB6rU0cJR4DijBv8pSe8Oi2DIA1LwusYI
qOK63rokZzRZ9Af19ppwqdqgQKY0zuOv2Xw39nbXHMEHlskJxl6JAwdbkNkY/u9p
PfnGrWtfy7Ljm6eZW057thFGINIIJngFwLtSLSa+OSeFbyDX6e51fSO3m7VPFal5
3BAbGFEZa2KfKvvLaQZW28ReY0nGz5YXX0AwtZPvCjUAiPOwCDRmKGipnOxIj7D2
3zM+Xrfnyq3ESa7YwdspZJ9klo+UC6gJ2MsIRNxuZoyuI/0nqZB9tCAdsUQQZeOb
Oq8xGiC7HdW7qj65/YD3YoOSRvr8gA56cW5LeAdyDxOK+DsR38ZZFTJmS0yiq3Ro
njLRTriUGikV2F9oh95zW98+e8vKoRCvMsy1i8M4Y/7+h4XSqGRRxgZ+OrBbxKlV
mjKQ/qqGhjP9Vmt9/HdVNIJNbt5lKWbY8IrAwT3W8QC23rdimiKsANW8dkUcKhtX
f2PkYCIcSYMfD7gLf18PqpndERuyTpgQB31ZNtikMVC//8EJGLOAdMyXig/79SKC
LXZUsQlHei7xKmQ46Zq0SSLylplYKzTi89mdHEbk4qUoAFH8MJD3ln4VMQYelIJl
LinzsFEVFVF8TZz7hoJsGzZHBfQAXFs34DfCt2PtV2rcAcrcSakx84FQ1LBO5XmB
8QuAUcux3Lzy0icZ8aF+3dfpcO7FDd+Uko1k10tgzwSkArbiFiuHznk+ZDs7XlUJ
bsC5k6x8sQUlcfcflcuziZS584W3fMPxvHhjnLas7yeXANuwWQyoU9d4W6/whxPX
UtpEjQQ4mJgobLRSoHObakj7VXkPgnMKOmiAsCfv0VBDtbwv2V0UIm36ZjxPh0kF
yBX+UUo9x4KZD6Tc1YnyC2/Shvgfb1qS1YZ1EsmWPwjAdRplSS/6fKzFdTOlo4wb
hkqDPPntBrwqJynRwPg//0c/XGbeIFJlii+22r6mlHE0BnS+Ouete25GJvw7xP2d
2cwK2Hpsu7+8f+qeeDmtAt+ICOBmMM20RyN0Zc6tw7feP3ShUgLbDHjAit1H9UA7
xQaE/ts7oGtb+TuxgCT4qLXQAq0zZ1lSZkwVUhUKDPCuIsmDMdtcDgAOZoDMuwPR
t9umzuK6FScTCK3KUEX8DvofzAuI8GgnlPIhyavFkTQZEEefWYzV0ADj3I+UAT/n
Uaj8Xt9cm4ixZ/CMFA4fkvhoYhJQkbPA6NGAoZ2GvS1f0ruN7TbaJVJMx6hn/Dtc
ncH1mX0QRWNc2F//Xx3z7U65LHm03DlLq+JdVSdb6GnPWFsn4QBRHBjo7/O/k27+
fdHHKC/wWbbxS8Qbkr+A0tCwkGa5HStWwBDZTE1Qx9Lp23HlmiMaCTaCJjvo6HE+
amcuAvBrd4HIorODkesaSMwfApYhlCBC710Od9yMideI+O2bNxrN7BkYRrnY9apU
W4ayCXz2LP6XzzNWRPNSRrIMkCnuyjjWZCTfFTLQ6jmvLtD8ECf9j63IeaGA7acn
gayrBohW7BAKY0UQfTPs9GIjMQCnspN8kwmNiBMcFDXGzzxeBvmvZBaJ5dVZzLSN
3tLv4YOhDGsuKlYO9Kof2q5NMY186MSepgrmTcS/V9dqSLm4jEGcgklbrMdN1dMT
FINJ/qazAKuKiatvN3fBcjArm9fptykwCa6oHYd3h+eGW1QC5Ai10633SBjjiHBs
n6nvIacwHw+ahkaSIus4VROffYV23ra5sF5XBGKI+3Owkfq/jFkoh1eASVioU/MI
AAmZqtYz+pocuhHrc3qkoZkuALwuSPFC6wRVzGMFJyMLBe4RyEVD0RGsYbTR5GeL
835L0kRASzERYDmBgMPWuKBcW+ofg+w12h5N45vNLZYZDM+S+1ceyro7AzR4QJIV
0n20GzR7q/Yy0oRNR4yv3x2iXKuQ91a8Zt15a5QXCmWfTaIFmVMff2GkGuGI1ZMF
eOEYNQygnxqChAQtXHWmHDtdIwynmAAuIbadaq0aP14Pm5fm/HM1QVm/60Pe85G+
D4bUuQWpoIIdci7Nd3Y5rSaCzs/60+bM3EkrWlLK/1cxUhUVeg5Vxsd48SoP3IZB
q61Nj1rrQjShSEUqaPZO+eEfjEpZ8sbfVYPlt+PltW9xwUnWaeH2g+PDUKqCmEZM
1BucHQXayRNndRTwLIRqn3zHGbOuNuku7vjHBmqBeGzWF7pGehh3Pyh5F8BNor1F
J6o3M3DHlW66mE2NeNR8BPpqE2Qoc+0Yg6DigZcig0aVLutPwZdCSKPhARvLtTNY
WIDvN43MF3BWOp4yH0kpbknolyNjifLS3IGSX+zVhncXAxPoxN3bVAE0q+zlKPIP
g++FvGXukX4WFW5CxzSnFe8IpF1tfRHJWQzOmVQL+kfqHcuztDCIyZu5vf7Mh708
S8lc0gVxlH8GhATYO70zNi8c97qHCH+YaPJoyV5v7DhMsrXg8kPTIDoziaZnvRk9
6d9qb6UZ1QdoyzX2p6pDz4rMhcvW03ygUYH7QvprTdBL4r2/Lo+W4xCUHimKOC7W
diY3I7LWjEEVAk2D8XNGlTb2wQaNlgO2zigsuPJld0R0qH/Cumd3vy/QWlHB5qYo
nNL8nSZbrx/MH6JYVG4AOS1YOs9pI61mu4hZ/ed2+TlQtJtBqRuBjw5kbqdLo/B7
67RAsEevZ/Ru7kMBbd8mdVjybD1Oa4FU+UljdpLFhwBVpJxf/+4HChVF7gzUAEzr
HzN8g50AEvKgmMBhn5NTalnGNcPEoznioMkATv8iBfHuLpswz9QUDZPKyVq11gYX
LiaVQE7UMYQDPpv5eFCh2Qgnbsash0kcawhe9uRZjrawsiihUqpcS3bjAGlQy5wQ
2OqGyOpqGNuqQjx//+vAjd5B3jQ590bN1vN+pOB7xEcKD/q9kmd//WmYjeTJPS37
yBRVo/QsPknPl/N6GCeb9/KLYGFxJf8gzH2D3lZxQQLSgejDi1//6BK9T9Y+kGrk
FT5NsXQQOYBqc/f1nPsApjYlJ9vtHr0LFApetfne6acn+ZhMnriUOf4UBckqcgW/
sjc2IPoarY5Y4Z6ktIVwqVTAFAGBY8HxZJck+HHjZKx2EdBLAJmeN+PtRHS/Ui/1
yZ6d/FHnomPao308+CcDsgkazsXX6gkM3Na1Wz/LV0gE89NOgZtB/a6EIC4yPjOh
feJTXCNiYH3LdBhXmPhTbPXbjo0UWef8cSUXp3Umid1v8Wzx7854nVLm6egHu8cO
4AoiRxcGknm+wHhjyXqIYbHtNAGQhqcUCmg0re8SpPiDsf7x8UgosKGJRezbDbtM
nEPkbxLIfKWuL0AU6DmcIZix5I28HA3EHXEP0QahJbBQvYeLkvjmp7oYX4P0Oi1Q
jh+DNLkbkNUKGXkPZ7hh6T3UYGWNYHx4NhFbRUYMWpnkk7gaPx6V2CUedlTO5lfp
9/RuArH9kMBF8jJfoCCJ2sh3/fyPIrVtVD6PTRu4UIUoqiTAwVj5Ffr+B6M7DVyD
qiyTuC91eunG+V0jDTD5GxykA4yFwcNUd7RUQoNNNPYV6mYjmI/1B7qT4ZiA44ZK
vLVpyIClG4zXS/G4ZA1rZXFWOQCzi2Q6lF0orw49sEsGX/K6HKo2vf1+PpxJs5lU
zqFKZbhkB/wPBM/HVZzdeUo3bTyRimuqAHWxNg5wOqmP9sv3lGm7P2XcxxBnfFoF
SB76dRm6xE6Ldbi7seUIf1wXIhJQSRmx20q4zMYqzzV/aJynwTHdNjPTJ/0T4CrC
oHV4/1YYygWMLZrFMK1afp/wknMvs3YbBBftE5/3dvro3tFZrabu0YtI2rTPv7ET
RrkQiwzpPHqYetV/7KAogGNoglfkNg1iRucHK6/ux1labg9pGsS+l3TXUASIV2uV
CzuYkefQM3KIaLskw8nq8mldVLWe+apCq1QtTeoKzgWGfxQlxDk+aUkT4SnwegHn
s36DwlzZSdgdDe5BQXxS/glCHAH4N38udyr3wzJ3VQyF6cEFD3cOhp6pNd0NK0I7
6suznTui90CfXmSBhi3jyQ3xt2TwYh/+59I1CH41+hXdYN+pB9/zRttwYMAzk1V8
wAcr+ARYtxyQEHP/mZe9unnGJkJmX2P7/J8mEKtG3CU+fphAlyM1qIwZ+pK4zN3R
5uD1xs7E/CaJGIeX1YfAWj2dRyQrrJHgT5BmWqg0lmWPJ1VN5crrqETomlymPb05
hltRmM08fgGOgJrxyHR9KL2vBtqMOn5Wm2iopq4NiXdGWvpttsPFpUmWo78qIibU
sNa9GmCeCquFg3whHU1JunhZ6/XxZhp+0eH1cV4gaOd0mQnIDX774NqzNvuA5Yuh
E28gIhFcXlsPKRjfsBxF6+uPK36M5k/vlEPwi3cAH9WLEGOBvcZHMKqilU1TNpjT
636mQxGq61rWjJwE6UBk+TRRno7rNxmB5X0ybV67khTr2VlF2+mYekRue36P0prs
uz/Eo/MWpPLmPjNL2xI1yQdPyXmUu9Rgz7prds4ZjuI0CdrJ6dX3GAlUxgqGI1uY
xeKkEjHu00L78dP2MigUld0ZcocbH7+OiMuFesxiODZH2/3QY3VOafu7tv7XhK/U
4z/2+6/zBksTTAbdvUoQOW0D9dx4CfX5l3T9H7oE2e7LclOk6VWHSWRKXvBj20Jy
bFQ2avARn0lgeRlpq6/6NBIJDusz4Af6dYXTJApgTlhJoGlzf2MKd1ZJ32AMsAQZ
28MA8Q8+zl5vyT+aEBtV3kOiFtwwpeKQCV/RluVyYzxeZmnmUz2/jOyYWzn5Wm9Q
5feYu0cxY7/MSkmYsYNhrIRdzEyBM81b20RN3yY8GC028+/GyPouKCrE7BxYlW2G
ZYEb9nx6Kv6534IB7dalmNSJ3/HZK6O+aneeUE12XFIDql959qsv63yTfww3Y+53
0iCfT454whmsEkrV/gvcgUyjI7nWKKdAwdQFSi3DWWXgYIDnWyhc/qP+gmzRJlC8
2hTbzX5sg6vX6cqcmPVeCpI1940fjC4HXo/fLCgxThv9mk2wOm8eA0H8H7k49q8x
UI1+J20s5eIrC9mVHTAf1FSciTIvoIEnaJNvRnmwrSZgrnncILo8A3/hHl2TgCFR
P6wdZbTDaNa5isITeDDxHOuF6I9KGDMiBB0Osn1Ul+8xnl3xcswRMNCv37Rf3Bht
iMvp6LNdGQ942SZuHepwvAySdAt3Kg5oDTV2sw7GqNmkvFYwe0vrHJIvBVF/8mIs
mchOKjtjrMEqa6xRnslUR9dy9HGkeOUKUbUxnrvZpe2uY8a+93BeK+H0btKxXDgn
MPcTiOM2vtA2ofkWXBZRii7xMIP2Wck0Avbq+/KwkRxrm9dUm/yyUSuc/De0EcBT
KeJlrUY8e8oLt6Juk5k1wJxzDAYh852YrQ0TZFJ1UzZgbf1qa0TrDgThZ3Zbj0tS
MgShtjsrAGxr21m8BngyCFeiMGJEWVysvlMTCmX7yV4AMJQ4NwZJyBXNjzaV4JCg
YWA9FPFQxVa5iRIgC9BYM08QyEgkH0RkHrMIw6ixqhySibsUKBT0mOXCZYM9M52J
Tb1qt5PxMeW8yxmlCgvkBKsb0Y+esXmwwso/GcmMyJOXhCxCj4yWRNcAuC97p8+8
LG1WJ8BLCm2vXX5wewpR0vJ0M6C+y/2zxtDwzwPkeodQRexx14IBe/lepSF26UOV
URdZaRWqBZGYyTutkIlm/vb/lUShX2hJsZp0/XCu1cWJibfYyL14tV6vaFFzFJMd
w0Dix3z92ae2+BkLO3+B/tL8o2JzzNCcgOSgwzHi2tkXMHJjVfRWoeMgHo+Qji3x
lceNapMQABhGO46UtpTMdHRqRYHratkTcitmVt531srOpBHSmRfikaanezuhO5wC
Uai1wrKxevnsfbUgqPl7m07YVX12w9xkCmyJxW26UH+wU7lmDUJY1Zb5vQRIsCwy
cCuLHkULWSnVsY/bein3BML64fO6iu2rGFIPQ/Uerpv57hB7OJsBI7rXWtG5aDk8
31EtQ/QG/7Kk2Illmq/UrMuG2Y1V6arquDBv5Ojj5XuARc5DYLkLZ6QPmTTm8NCA
baSoBtZhGmxWu79jSY2OkQGpFBH+uhMmUu+n42/mKImQ7FTJs3WTJCGPGhgxZxyC
d/S7WNpfWjTorfu5OJvUopOmKap5hKnIbTqbx4lDB0x5Dz/7MU5m3iu3sxm8qI7O
vwJ+3uKDoRy3jwg/PqhmMupnDkMqlqTKojW2QKOVYqFaaA2bTnDTCwy1Ytpxsfc/
HvLgZhQYHAKrS1CXtd7N3IHntvhcRXQ5sire+ug4TsOc2iFsrLB1tWfQl8zXI7jA
ZPWgtbvIvQ3t1Bo6Ks+hDi6zF6JCeLrz1Ykj0YToZR1jReBQcZLHfcd+17d1qD62
ET0Yxu8kuk0htWOYSVPC09eBil5zxVXwPZ0YDtnOFTvAD5euxnv0GYhJ0w3YAtGI
tmOB1WI/BxOb9H/2/NY+miLN0lSrkohNUZkLMYedPlpEhV8yZX+CZtCEHCuzV0+h
jlDZec8s3QFb5Qoq06/kjeJfT3LLtbfTusZ/dzdVTHvUV7UpdqFH6jLF1BP2ykMt
VVJut/o7pNnQy0GnYuzs0sV4zKC3CzMdKx5FsdLbBrQNELjiuaVBrBOxOUTkOi9l
1YatrQQOm+qYsg/nfEhzUpDUbz03eSBsDMW5GwTMJFJ/L5iCsfI3y7A7fLWXvF89
+aFaW92ZkoGhvBqxBnYvRrt8yKjwHs9fnS7AQvdQXd+zIZc1qvuhs/ebWinPV7BK
17WkezEqr1xAzd/U2sucL3Ai6PLwzYjxM1E2r0QHO6zGzxxAn2uMhE1nqDuUCf6F
1WkjNOezZenYltyB3I6XjTzcP/P4uld4WOJ6co0qf04uiztzqJdQ+5e83poocGvX
1m4GaV1k4d/zVf4jj05kQRD9TfAtsQB+E4/IVr//IzrFV1EE7UJuVq/+MGUx2ygt
3aB5yeBxEvLEViuTKxSeryCCH1TpBH0F+7eBdCR6lQm7xBp3pnCDczv0Vm/1LKLs
xoznj5Weh8MShnIieO8LgvLW0GgyFLLGxm5uVfvPgMKG3WvS6gCPgc7SU1Xt0dU5
OpL5GoNYw1ipw16vTgm7WiqoCjIqtewQ2GY6F3MPagcH5IqumgMxuAcPzxtf4p2x
bNflpzi++43C5M/h9o7EUWTWp6f+G+2p7LTTT9BUzhCZmO0IdlBxt9c3cD4CWNOP
UmWgU7CuKvwKI6+FLIOAF4SaYihO8cKzsWqE5yx+W1gZe6eJa5eJ23uT6YGc44xq
J8X2mIwGfvW/M6gaelTDCzzLDelFdT6Dy/Ig4a44wlncqBcHkxY3KyVpOV2cd0DK
JRbI8KUBLmeFD05wUfd1QKGxNQZYD5CtptRoMcj2j7B2kMbhPiS0HCrUuR5kRKNl
nnW5E3f+Gqw+MGe9pKZ3uaBb3c4pAXEGN/J/LLNE+en1Eei3OY+fImTw4Ph9tz/m
vqekrYaUgMBV/jBAJ8+xzr2DJzySJmIf6SzwS5IfDslCO8No0Ia2jFqwS1T9w2WN
CZb+sWxiIDirWGBe0nhAAtGn0ya5EAy8zdOqjwjV1Zn35Reu1HISeMZoR4y7xaIp
haHNerGnrhA+17xSsR4dlZWCa3iAhEeOb+8ad+9PlSYrbB1wnfT5cyovZA9lE0Nj
1DRIWXkenbHDwnTMVMqlL6n52sA7tiAJNtJoaMJHERwjSRlYYLmRSMICC6x+MUcU
lMHy4YEX+KVnaYOjh5UJEHlHwyauzqUFlp4TqJS+fZRTJ7h7aTEX1RWMjSrkVepJ
jyfIz/OIJszXqZ1d+kQ+qgqDjJA6CBT5nhO5oLFxnKVp9wDWq0UJbofkdIt5nuyP
BnKJYf+D0Dv+oUrgm+x9yR7mSw9pqF9iFgPX/8FbWsLtMuZIGc1nQHF5yeiNty40
3R5RgmwxVvu6UNypNEDk1AMIubIPDQb4YrXV7anCBbVBPX4s3MWuWCqLUROtAL/v
yMziy5LfLsfBdDMaJ6tHgrv2m0TH2HJf8cgznup0GWhZ8OtM/FoA5PcrL4qKe3R8
mx2sdRxVRJejthsf/z8iMt5M4gyODcreDmKcA1YHUvp3ZzuUnM8R7MUM4fhjeD80
R6Xotx0OIrEIZPMvnHLfmM8FhCXFuS9mO6WuyOR2Vj6AUT5FD3aKqkBjTQuecBdO
iOHlMRyxSl1knZVFHPAoB1hgVM66sRT1ksnqpglFZb39KZHpDICN14BsKnuQeC97
3ANx9dWwalIZWM6NqxXGoHnA+V8+oxHybOzL+WRiI7fwGDp41BT+R9ihtIvNz798
DEJ8f9URegUiUEVsCVrGYwGyXWGPfj7i8McD1YwY1bV8R7IfQ3h8wbr8HHGfRdbD
DxOP+Zv+dfDgEh8WfzK0LCxkM9hTwWisdS/EeC6RPCryIV3bW1uwCqINRCjjcV5o
ZTt45+oPJn8pM5kLb77qgGF4+x9WQUTJTfza5lKLSrm6ALyZTAHSi6Agtm3c1w9D
e8vNEDNNjV3U6WE6HcKqpuw8SmSkoA/LDx3Vmp3aqRvBDXFLc91KV6nfSI4EQZif
DPWCrNItbh3cvnMiQjVe0mDMyo2ElJJcGnSo4GhVGBLBklbTR2vBnJxtwn7WFWKK
Vh05m7eT5ynrJ+B/4ySRTRCTuZOpNU11GMhBNKvV+9/6VixGGKOs0iSyBx+ksTs6
YzJm3ofE5y4gKkLs8vk9SPVyAJ+3CBtXJBfvTXwPiYjTwiV6CaAzMFDwFmXAwkMZ
k/g9ZSQfDpoboqm8NOdPUR8Y3TB5DxnEIbn9pvruQI4d2UrZj38o6QM/rJnSr370
YQ4Gz6aUGz6aySOE/Bl4lUx2A0h42DsBEQaEq4UjrZ4Kn7OJBsMq9fsQl1mlacQ8
vxsttP+0iZl/ElTLPCGNyvRRdmZ2lORvT6su4cR8VWVusAl3Bs/TwX9IMg8AJI/S
u4mnYodSYs3lJkkO/7EixAfc6S88kPIQqAgHU3UwUWQZbDo5C0UBFsxLfPyXFxog
lAT79gyJNWORWkKvBtXII99ji/kwZtXy29vndn7RZuoh9+cYwbY+/0fsITWev59e
cSx0D15y0z+QXGm3Cc3Hmvbg3xNm1mX96ixPPMaIGsqgH1151tqqZsE+vjBFlZTK
3r+Msrb8aeZV7N1s2hJOabcm0h1+OLNjjaKo8tklflv/yUSNOXOvTr6Bzpe0q/zq
RiA0k2lJlB4Rhrhj7NiHY56QXw5SaYlWoUUEL3K1wdod8Nv5/TiTfZwapJSY4kwW
idX2LIfh0IBpxSOCDZ2qNct+zqVd5IFgl695wLsR340cnRpjSqgdKfyxfnv/b4S9
2t2MVn8O56mqpbzyxKRd/mJtCS4KXohz6IdJH99UWqxbjRVxL2qALSsgo/BiVl/h
XHM+u5J4svIsPZLcUja11DIPMi3DKbxNATBIDW2U+NMOVt2PUyIs2keGaNJYeAP1
5/GF7JXtNzTugSiZ7mXrs+Si1eg+Sc51gQ9cVYl8usjUk7C71F2s+/NrGqppf/KE
/fe1hJwkAXel28G023y3zDMlBmI3sPyvclTTIr+v7h55ZMmmNNm961PeJ1Cf+d1H
q1VZbps0DSMvwDoqM4zLr2IVe0Kq5fQK5dPuzxMJq1URbJLWT5Xpi35jAPcOG/5H
w1mcshbMlV45BS2fSryso51C1HQj63lR+b0n02rzQTA72Beg02vRxqqj0Xxl9yF1
DFNYwXQ81TMpSW9lNH4958gjTwpODtvfDKy6/+tbUdTflaWIsByLsXbk7xoqR/0C
Ys2jqh+8OJI9B6TkWs2v4Kpjd4XiSF00/ejvzbzHtND+bFrf9slrP1Uuwx5lubIN
QOGcJnOoOfRDMX8THKBAMaDC1GVmq8fGExHyeGAgwnXSPzD3XO/mWa4JhbQv1QzB
yDMd2nQp62raGxyR7ANEszT0CNregMh5oo7HiOjkbX5qRWJ6lA+74fdrqiqaSiRS
FYHchZeldGK0zA5BWPsI7mnq34WnAewpRryJ05CTGY2ZmOI0CoYABqicItjs4mTj
qklGnVdOwZ/VnlXZ0/+llQHGS0aEmMBw3UxScm+0MwFvDY7Vk2NULeFP7Ocgc+0N
mMWcj1tigWc9sLT98ZEnAm0o/r/aUULcR7I/LCU5r5tcbwTGKfWKDgzDvBqy9oRI
2Jp9CttXLiAfCP4LYqAG03/XjYZsfwRtWZft4NbJRB6YJ79Dmj9bL9Qjr9oFP5i9
NnVzgeWgDvakmLXHnApK8IYn7wDL7njmfBNFSJUiGYP6Zrv+i0hAY5u7qr3sv2oN
U4NdCbNfGOLWs3u5dN9lGvf7DBN7W6n48N/YvKsk+Mg0pyu61O8PqDg7k8n6QCk/
gt8A2U6gFF/i4eBMnXFESjzizsHIaroOefxiiyc7ipvGL6XFgoRsRB3W4vf/Qid3
TL/DdNI7Zh2gJkkPz1QlgIak22AXj7aZhMriNof2f7MVxs2lgKwcU2wCqG37gxs0
weuMFPJpHI3HWnaN4fm/8l8Sj+NtJN612R6gEVs+PyJ0ifhzxgOHhMdB9jy94JNa
fN/qTNRuw55qmvLyqE58Qn7YWZJbDjtMuh4iqQ3UkdHXnmH8J+peCGMXOrBa2XIc
wPH2GRqw/38C8R3ardp1vCUti0hUesid3Oj0i+emtJWYVLJryp7+XSPy8NMPg6ba
RHTZQ0e1qmqrcAXuo5uswVWYOfJyKV40QD/0VVK7plNlj7YxJ7ra3UMUvvtQDRBa
8MCQJb/BA27s2ytsWQiSe9HfBGp4W+8Lst9eQGB5WWKTPc5XEiTNaFePU0y5sJU7
RWwgbevSk8a6mpk3dX2cOjFgCUJbJJbanjVlS6QhmBU7glYppntYZ5y+aKbO2RWv
EikrTW6F767eJy1a/0jED4TR7dURzRsxTXvQ7veUSVJP7cOGgZcOR4XU2/w9r06f
iO7O4N+ge19aPMCSHghL6nJaKZzijbb/+eslHWH2ToQzDXlCP38qBxgw+ddvOeRV
9C00C2BcF8CHddc2/sDxLxntyRKfUs3LltG0GG4PU+PpUug2V4sdJvlswKs1RR0E
WIXh7i0RcUYc8WbQl4/fx/4Q6ByqkOMl25/vAQSCKiRFpPx2RoVLgOI/qCsZZ4bg
B+sFihQ8dyULYaJI20fG7FFL5vgurbSGOzdz6Mxe/u+x0/GyzHXYztBSlZI5das9
3kfWVnRwtfVnxiCiclzXEHg4Vf95MOT9Zxu6yRAveszwGqEcc1jwQicAeFXzCKAa
QBfI63ScVL598HTnhvMoNOMtzKNrRX+AFqUI4uR5wNSmpDq2RRPZVKLmp6GSU6fF
fEolCpITc0/2MFbbTK/X00XIINxfR/odrKl2v/aUS5UX+bu8izfBtSpoDSQmHdWx
vJ/dRt+29LOaKCNXidvMAQCxY6sL42CaAxonptcpXnN3H3j/1UOh+Ad4ZC012Khm
HPQm0UvoOUOBpRpYpuiplSDJKRYae3wgB9W8PM3PfTDmKBKGP32UbDal3XIgY3Ck
iLADSepdN21inC6GVCZhf4W5lujuSnqmaNYMVs7ScJie6C9CmFyvNTJwGvejbjxH
OOv5s4TJqZ4wegzhkS1HuhB6XVOt+xmmACWQcULRPR+VuCSx+nAnI24iVbIfPR7u
gJ7bG1VATTcHnTQDye2sZHdwmSuoSB4f+m3v5gLBlYMJV69Zbj9NJX355Vo7zYH/
LIBUy9mBx04t4ZmU/Jlqt4iuSTzCDR/0mqQveK/mq/QHPC+bIN04Y1ljZpyaX8uH
MxEm3I2jjbTs1/QdlACNg4IG+7c73h/1vBD4TDqe5G0PoFyDchv5YYw+vac8tWLA
QL5CbyssOsy9hdvLrEXcEP/T7tt+dF6HUc8GipFl3Nh1dkR/jL4YA0/EFAOMtlb8
xGv0AZ7uf0hZNEyVceVpDnrR/Qg3YgWGEtq1Ys2ZhS2s+tln9r5SfnnS/A2b3Mbo
CHh9mYtgeRGUnIwiET8yn/fDrsM9rdBwiCFoaT6Rekf9LR03+A/e1sm/ddC4miXl
B9tyD9SVZLZzNOWbI+QYCROS9nIvcI/ZPuVgE6MLwjwOljjeeHUIerV2v1mM5wbO
ucXYx8PbXUrrMFSqtAwMKrDxIMxl7JAfqphyDDV8Nu5NN1Vcvsi8005kOzD1Wb/h
TmtkuSxQHuCxJplCYf5xX6L+cUhkrcUrfzx3v2Usdw65JOEZyRRLgh57d4vdQuoI
VRmM+BMkMIUvyic5rDRPi4DeoxBzIMFTjVM5tIHzSfy+malFmJPLVuc5Xg+Ispgk
BxFLfgbytYOgYImFdsmnZih1LxbTW4AYtRUyHZUa/aBtA2iaydM6lbxStEm47VML
uWhJjCyreUY8Ss2p9belit2iytUAZg3Ew8R7qgCtLr5d1SQG/NPmYqcctGDFY0xs
PhG1Y3YK7avuJHaOtSBl4VohZxByVSN3pwDlvDL4VPmxTNyrBVW0SfLRmX8z7uNP
CPLpXoCgDk1f1+at8RxwQ+mYOXYtbsT8BCmDnp396CDX5FEcnurbMAQEm/965bWV
ayulp4Gr/IZ0MV1H4wzFxLnqdHnbHEnceVVWYiOFZ8aMG4h8ruHXc2p4m3QV9xXE
tOmOoft3BfwRg/MBgrYCWLjoGai7vnXacV+kbJ/Ud+fxrgjWwuuWd7ixwne0qSNh
VGHOI75UMUW8LIEEMop7rNNKAOl2AQ3O2kpniMTAhtWtst0HGmNFNCurERLaRST5
nfXoW/7eR/gPORFpqUzynaCdnc/SmixQiYwwS+H45CiImjQPB81EypdLdrI0Sv3d
Mf8iCeAMA5LORbpaE/NEtE1htOJr4kEpRycYZU9LZPzNzv9iv7iQ9ECXuYqbzLyT
UE4bhxuSkCWiJHX85D8/r6bXwz63uACrQAgy77o8kJZKT91oeUu4w+64xeIYS7DK
pK1iQ3rxupYnBsKUoadGuWIv/niifPkq+bPvAm2Vvq0U3nXVoPodBmb0ArnW4feL
LTPxR3yt2L9a7rO2/v+CyOFYr8/BmwsjqCheyOX0ajeFsftARyvEpLvGYIYw8RLB
O6zdvyBMEoUcqDxrs/BHfyIqTYQtkVYOFLBRgF3CWJQHXAbRk4bDD9+vR6t9U/W3
yXZSCdCS0F8fKB4entI06+hRMuq85lrx3F6QLCqkoc99a9oSZ0RnjvlgItK9QB9Q
lXjCGmhQ4Dxyld8GETTME1YTUNvGnnhhQk6qMEXIntsJQluJ490/bFt/0AOjGu/J
xyoxE/U8qDURPFaOzo0Hp8w/D6GCnDPdOjPHoXFgpjKAa8FYsDrATP3mlZ8Fwr+j
YbaB49lM5fi9NhuwfX2UBY5/9RrjOMbYPYB5UF16Boyo3wOt5Lvo25JvVkYOm62y
ei2G73yr8m9480B7sEU4AiWlkiUAvbPrB+4LbdMwkAyOZy5nUvUUqNNvH2PktHU2
tGHuIucwJPVrAh2NF39z7bxRoA1tYx+t7dKuKb60EYE4fxF0vLtZtXb1Xkf1/dVp
YwCkzlhDGwh0TQV365n/Ma75sNGtTiAou3oVgo/d7Z87ea70/SZgQsysUwBHbsPR
wxnDb3JoxG3uy4B/FdkurbzwRjjhHPFr7O8bBvqceNTDEloSg9FTWPIl4sT7vuUW
t8oEqv9sOT5wKmuTM0mvqo4/3NVpEXbckoMxCIGgq8tgUebyGuEGY7Y0lvFB7Bw1
JwMUMEzHrE/J804vdmzTElnQCI/YAKRHrsylOsVzO4OOVomE4Io1d8Je15mI4bSh
gF+v/b1juIVLMR/MaTuvV5HDOClpt4m1ziXIQxW8ip0pmSVxBbEKdaSR3ayE/2IA
fr8m9ArUg6SNhQSAHeRtV+MzsqESVJoa01Y6ugCrwgb4daFB6nr7oy3t5ufxso6U
hv4pzQ/ULndgkAdgAva9FcXIqaP91UNPhMtJr4FsiYXTQd4kU7mY1OG2HIi+T579
68Hl947rX0OFrb08dY0zwChonHemU2gk1Mdrir8Fbzuoxk64/2a5K5QBikVFo0nw
0Tz4QRtLvH08DhcOfAflnt/d2ccrlhIYePPxla/21OYGRl4Qd7yeSh7SM1cIaaKu
7WHlwXR2lDovMAYuX2wbZ10XuhNcgOryH/DFq0P8RPoTuCZNXdBLNi4jfSCWPD1B
uiJCAYKKQn8Olr5Ov/Shw9U+tVaEN8hx97ROBcePf2SP0Em5l7FxEpRhIvesGhEN
PVrRz4Ghi9R5sbC4L5iMHM8IVXpJE1OLMPMxfXxV92UDVqTM+nauiK3YViNprfva
0iYDNEGb4c+2JFVR1qVbWizAur2nV69iSsTK+cTgFDBpAORWlBViXeFWGrG03Yfc
9HfZKmoJjh96zDzGlKYB3R/TcWBeR8DtKnEs1dxkAO2VYUYU6SOB5VobUDZpmv/+
sogxEBGUmVIiGg2kw8mHyZCFuI8BdxI68ABHNgW/uUkdHTABKBCwVXHYqewYYBTG
spMVd+JuNfU8opfd2fiYgSiW6dT0fXNmIyZ9q+xWvQ/q9oeFxITooqj+y8otO0hM
GLLDn74tjkrfn9ftJpoGaEUUCXPzgxLmq6+1NVsiRwCQdwBBoJf8l1mE41bPjGzW
ADEhzcImMKaQIdn4kgli8wCJBo9V2MOLNOAVSe3OUai+9YZfVvJLWlBgQ901QEyC
n83NHXwpqzPduR0d2apjlEMami/Cke5gZYlCBa6APOWHk625E8GEuTRMerYKemdC
uv6R3fX7aTES3yJrQKgkgSU8kZZRLNWkuFtdE+EpRSifYqOSh6HD+o7COsq0ih4F
ciae1A1BZwb7aHsOJFQmhKw95ehScshngaQZbZcx7ZAS1OMZ9rrWtHpDjTBMuuXt
PK6+Nk4vt1bM5sQtAwIU5o6J0EY9fYTpmRY1fBG+rsuezNTYIEQb9PSBGZylLrJH
kKIw/CqOe3zs0B0LNFHQ+/HxUbXoRCuNLHr6mAbZ8kWqgcXFqBp/MvyrgserJvjb
1nEPwume7nyyLr3FYR/Th84FfXrB1tl6wQ0RvtkyMst3McZ4biLyllg2+iZ+N9NK
fL/otdUrxah1A/1D/PPXhun1BHoopofLk0wvBefS6BkrdcYnvBUpTH5WwiBWS7le
VViecZGJx9ikegQnhwoqe+uN2+p9K4MCvRE6yZUnopgxBQgwNflMFljYl4mnZo/E
0BQnYu61UUo3Jfhlyvb0jxzmQnSoK7Y4PqJRrrrjWj1YjBtH1WHmimPIVFdvbEJ+
vpHKrSenwm1QJgjfCFZsTwiUc7ThZ/S+DTqccJM56b2hK+QXYojoQVsaWA63JZcI
v/98UzfOWqo+Ja2UtwOFmPu5v9QMIpCtlQgj2I4FVsTRSUM3/KzUQ/IDxULYiMxs
N1wjeJ+rUCEBna18sFp0TsXserIPFCr7gGbVJcU+87AG/1TvAoi3gh3HrPHdUiu5
dSN6CY4Xbym3xjdd9uSNVtxokSp6k1C0SgYRrX0n218K96ExFn0QBcJHkZNphAfe
GXf5O4KBMR3U0oiBz4Kt1iPnJPQc0z77cAibhZ278wY80EEIV0Qz/Yy+d76d1uUU
4YHtSyBv3xbA6cMqC0cjfFiTXwx46breG8Xt39hNgE1k8QD5F9EyFhbRME8zPkq+
RuwYgBZUc/F5xCJ+rcBoLdGwuNlg4ExkDn7L0ykYCHo3wKAg9SZOlzWqV1icLA9E
Y3MyjCp85iuETJqXLoYURbvXyClyasCA11PduD9sSz+ku40IqCErvhUa1U9CGuuJ
eH1hXd2ivE2TrOC8+qxQU+GH8yCZZ1TE5C6u+bj2Th1SS6KkR/jOHrN1orel77c3
nbBeL+F7uNErDFBR9renBmYwFhgQAvrqCAIAytdyWU8+AFn1/ohDBS/8a7O5ziER
dAltWeQnuWxdSw1fPoadholCNlKj1kmQJwtlDGJdBS4/wVG9Dh4QblXHg05kCsG9
REqZ3KKbKciOfQ5S3wIdep+SLAC5MFkhFbqTJnY/xBZTF8vCz7nlp+g/ykkj7qYb
Waju9ePfIGS+UMx4eOtVKIlWcedYYIN13J5BNqBL76FTRHhGA1kbGl7CtaNy0T6j

`pragma protect end_protected
