`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
aVMzNFjrjMp01lTHfCbLGVXFye0ap2/Q7hequWqi7Ir8AheXmcdtNjtnm7d6OOXX
vutjEzcR6V4nKrDUhgM5vGMMXswLZKty4yNz52HY/XgU2YdSSrnHEzQzWU5eSIGA
JSS51zTNXxURGAUaXQ5osryiY4whouy2q+EXmJYLk4o=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2352), data_block
p/iop0rQQVnUZRKPdXjPjIVbvvCqHDuD9ygc/4Sn2cGhw9wWXMDrVODnMSIH5ZE1
nJfinvvhTt343Mv1SGkNRbFywSYixLxesdjlyvY5YAmcIZ7Z3w623jILp4yIQ+a4
wTA4ONxzIzhKABEVgh5D/5kpcEDVWXxgDV82GlZAiZW0xWoAe/wzxx9d9cI44mFH
dUWcBw0iRsZ3nnnlkx7DsbMVnuvsMsFqdVX7EBqI3U4jMm9bGIiuj4FUMZ+eIPL6
YyV/+6hPRaFejZ/37V2/GlULQYyBAfS049mvUS7EIhuBUTCMRQeznQaxdOLCFWkC
Hku7156AVioJCYx9bQgXA45XrJD2M0wUyZiZiRAbTPXAdrCZXSNug07+CeLJrTgI
BwIqTcRd2LeT0WpotB6G0yvuJfcHUPeZURKhRS2ks1mTyEXMPyxJmLnj1pB7TacD
EB+YT6jC1myDpi53OkicjxcsMqfXdvEyjiDzubNDGthQehaZlITk51YtwjzS0U9f
atNiA+C0rzVlBHPKfr+Smqf0/6FsBNIh4iPP9N1bYNcF0mRo3L4X9AFNIlFtTALy
vfdsp/2SoE1xkz3N5z9nPJ/QhvVi3xXg0MtiINAyU6Q2ddWnGcIAK9+Rg7VjTziB
7qtgMOxo6Xl4vEbfWURKJTVQjC/zMn6TX3Pz6vf3q4mSsyZorlf/LOvX4m+UVHb6
PDe805381wbs5mjWCfWAajv4uW7pSTu0Sj4wTDt3nE87jo15p4pmawQ9j9Xkfkkm
0eIK1tW+ekO8MWHCMDObFNYGKWY+ddMypsGPC7Asdq0wP+GUs7pVbogzbiUUoaDq
4VlfPEo1oFtFKZLHnu+oYUZjoHJCIpv08NoBZcLVKVlxdla07I+slclxG3JEjpLk
SMvU1llp9iqqGDZz84CvwRL/f2FWL6gwh+hmDCJTamUA49WQueeqYpvidFOTDFWS
nyWPqs7D+yg04+8JI3MkWRvhwQeF4d+wsQWIwg8qkZ0GDZsOR9N8CWxKymHKJPuc
1zIUJCXT/JgrZYTL0hTx9nHyIJIpvJ78nncl+yBQxAgR9zWMxq9Mb3QA7MCj3SPm
FoowgCGPcnFq4hyF865VY/aeM1ZNIzG4GtEW+876Um7mS2+D+AZbmWc3SprQqPw3
0abHD7mw7TWjLtyDeSTVMpOYYG6BMTVzluQ2WHmoxTHXdri/1LbOQB2UzgYAe0zl
cfVoLZ4PMo/3RGzCOJNMNNWM8AxnGuVzwYb5v+q/qEMy+eK6ST7FhheXiOS9/asB
5u6CdPh280vZW5qFlvddozw1gvEpxVqHMep0Vpx6jYRNmcn7t5lmcvWyK+v356Rj
1waPEaFktdU2H2zNl+gLABeNLctuFqTfEXE3McTQ2LNXhPB4onHqhx7KdTr+DC7N
jFmreTtgVr8CtXm6SxpEQEo2NA1AC73GqiEEjdyiSeUSjPHEoXyiymjURjoJf6z8
2OwP0EzMoM53Vuddl7CiWjMM4JdO3XVAE1OnljynYCLooTIPxQDipVnoHNFMYyXW
SjkJwu+qpiuKi39CW+f7hpBV+F4idRow5OOmHPgPI6QHZo69jmVPErEcnDltIxe1
GQjG01tbNbVx6bhGDebKLw+UKFfzSq9tk2BFp1u1pqkvg6M0wkw786SMYZGfQHTz
T1so3pke/R2h6tQ60E63op9fgEW8EvE5xHhWbR34UIF5Bs2d54KJOin2gbhO2aNT
cPDmxvyyeiBVPAptKHnUO/+OVbO/gkzjERrx/8fPDUqT3ag/oC4KJpAZ7QS7Oexj
JvcqKHMaaydIZHrYZLSnHoB6T7wAKnOg2JE1ZEMIhSMP43ypE1rwHrPk5Llmmohm
UeY7MFG3nBxjrdNnTg/D1Z/1mBxyFrGLV8WvwKnLpdaUF5WW40xnK1AyTNeqdstX
D6akWAJgvruQYuUGo1BYLwUhzbL86ljtBlYT4hjmoRHmf7Mgr0Tqe7p54ojw+Yuu
vADvaoZ4/LTjRrydsZaqTAPV73u44PkPI/wRsEDSoWl7wR8cTXPQmtg/zXpn9hMv
P4U7pYcZJcLuHGOMlG6kDWmalWIpxyobCFF2Zmqeh2Iw/2IAyWDJmy1am7SO/bOQ
XZvgX9h8e1WUims0BSF6c9zRCMdzZQanVTFOybpOzSONIGILzMJpgvP0mcXav8YB
IK7hz/MVLyeNnBBUNtxNAuzaZWG9gZKXGfKmP6sM4W7P7XjktfH9T4GSEFXd9bTE
ZScsWwRFoDj5AoVqQnyEfREa/yQz0XJ1VjgRffd24QgZUvctJx9CyzlBElmc0ni1
JE9LOLbL4c93nfdRhHYXYg1UPHDRLmV1Ai17j1ZxfYoj7rjJCUCPcTVmJ5wI7OQw
nYHBu+R/LvOxtrAFoUSKOsk8+xWQFExCGBSQskrLQS8UhD9Ns8EZhqJDCBEimllp
E78ELneq91i9wRUdZIQH/MdXHdFFegxP2FC3h4SiJy8GpY61NickN//i9yK5Q3Zy
Z1Blsv9yfh/RT/xRwyDoS4gavjAGY1k0Jfx+QaO7nXDltgRYpQesX6y1mUIbWSNK
OsbyaWxyZsssQ0zMeq72LSJMMJZSpmSrNMLCb4qku82Z2NNb7S9/LCRZrTZ6sYkj
CDRqXAgCeoRyIY9m9LaeyXRznu9a8dJMYRWibvKD8Kf/cINRZaRpxA+wBshNh5pH
SrU1g27q1sFC/T8WxCqqWeGvX1I4jcCzE/ZTHTlrhN2HMA/k04wtzkDbdY+koTXW
t+3SskSq9VEcHgsNm90910tFHYm3kC1eotL+sI9s25Ul8Pk5oZcXJ10BJwPYyw02
/WmoLua1wkJIqAJYBUbRBZTjhq0xcXTvOiAURgzDgepC8Kq0CsE3i+xKDfDYoYLs
ny+8RZORlkt7ceoCrIzzaGGJAsuJcK+c65Tdc7IhxPYlyZicLr5wLiTjxktLXAAD
7FkziV4ARH4pYfYFf++9qgx5Bo9AXSetrAZFhKrsqtdZb/lr7n941rIIlbt8AWjm
e3qJt4do2aBRZDNzTWZt9N1doycBraViVJQdv0V527/3IlAj82D/A+BzpEZBeFhN
QQDUwoxtxKWPJipA7MHTb7DpoZg+rMQpdWQoYirLa8l6R9u4LTXn3LAPCWXLilZd
`pragma protect end_protected
