// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
t28DyKriUSORGVWhlAzOVW1mYHN9a00vvemQCob+JLIj01b2kFKM/H5leRCNJvac93ObF+7hp0tM
ouKER0kwdysjzNwXrVwUYmwSdDVtmfpm7dAr38lpZkYRRECrWnZs3+HIr7Skjp6lZoOF0kBkUwHb
Qy9d+PgqpurR3UIEKvJKss+UtlfM81Lf6/LcYtxeS9El6yC3i2LT/pKM1Fjm2+6GOkpbNmTnhNpL
eKTELjwUSt/hKfwv3xhnmLB0OLS1dsm9yi1vHyZh48d7aKqFmvf5ZYqQV4tlAerjelJj75I9aHoM
BkgVwgFe3i+8SiK95AiXHtspoZunLrQkiTXWWQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4736)
Qh6FfAuUZZqne0bqYOy9V9IDUIE/trwsAUKSF/UIpRTG5turYEKRvnxDBB9DJ2v8YNj/J6MLkhon
xvUVugNnPhtOwRF3c2u5k0XcdLoXgmnWLoY4qzBX7LeKw0FpID6FV/vjNl+Z+j8L8E0NoasNx+MC
WIdajJr13Cje+QJDjILCKGdV8+uvXaT+a/a1HYKZ/uJ/VG8lgjVGVYXJrQdUW/W5KvwbkB5MRD9q
mPSpGpo0Ew84NWcmjXkhSiSbEjpqboli46chl6uhoQMrFMRrn3p2AO3uqrp8ZKd69MgukJd/xeim
lpxIO12S1nlCB2mCHWso2u9KQ/WWMma+xm4Xp2Egwx1km/C3s85Rrzc9m1qGBQ9E1T7m1ve1NeQ7
6JkeJCGwm0v+XgMeYnItGWkTYt66M8dEkxfa8oOM3eMzt0x6vTaCB0DkTSWAEQ4Jvk2CraYBOA5l
CRYMkMLSZTZruwtAsv8asP9puNkXmW91uSy2s/OFdWCpyrTOZ1JcIgLgeQ592v1mSsPqGMeMeRGv
eQBrY8AedaeqdhxVWoLYH6B1ItXlz5/T40cObUfz77Ch6zFqvnLB8elqaPxJmSMMkogxEHT+7arY
j6EWiZW7RLbYbw0/SeLvis4pCb6oBkrRWBS9j4I0u0wCFu94Mj7RNjk3Un7g1wFCGmWpgXDv0akx
NlbpB83GBvGkA8yqjOwSia8uSAHZjSgpPRD4hpUHGMxXRs4T5A0Sb2y9QR+tYzVfV6vKlGJgc5Gw
eFwXSm4zg7JBVzKoW1NrKPyXgjyp5jhu3U3YoLh7O451fOanOs9Wjj4NiDLFTyS6dVxVvV+R+l2H
FE3Bpuk87+zNC4/qEwXs1geBDNmiJBPGy6zKHvK84nPoxoDfiLXYDqoXsicBsu6Ppz0Xj1SGKSl2
bDf/8G/xm3mNBXJRSXWi4wh403WU1uuOnUFCvS2rwx9aUHTIZ133Xp6tBq3kDWr4UmXsH9U6whx5
kzTOi7rvlnB1kLiFY7W5X6jFCfoOjVnbw74/zPSF1ZGG0hrHTgkGjB6SgZA3chFmQGLVzA9RWBqi
Lvo4qkv4oxveD0escF53nmMDK9Lh7EXG8iJHLXQ/O+ECxFkClOykRjUL85IuWOaShcfZE6QrXNSv
D4tYPf2ZMFRRLS1+nvco5eJzPjgzs+hfHWhAyFzRMI98kldcPxsx/i9GtoizUKHMCWY0xK44MrXm
kyAX+JIXvVb9YkX58zHUU6uDYhwuO9t+wZJucr4OxKCf0UVLSfdkEXWRzyHy0LP/gCQlRHOSZWAr
59aiX6E6fb/6Lzw6Wll8AaspGQRKlCwOS6X941b+a+IxvQImUTLTwM1cQMraeKtl40cm0yP7xCgd
kV3qdNZTeOdoownirQYlybSdAYWKBje+t86/y77kLq9mLlwKFodTpj0+ucD4pMNwyq+dqK88+ek2
BTobCAaqn10S25bmWUD/Ae5FgWoIiLBCViOaCn+XHp08B8zOGZpDrfEPg17Uj/NcXahVV5NJf9C1
md3mWJhYwoVoZDb7XU2Pf9jlQ21K7OkIX/eu5idgHh85/epvpPEmh47TVVZfGRPftcs/gVgVyv6s
cQ+PauNQZQxUNxbYMkCMtxy58JwOr/ik93sePxTRmuQzQ8lM9CSELt9nHyXed0H2GhlnXw2z5kel
8AkzfPJBr4CGhxespaBqMbZkpc95ARmdFKg4XwAH8oNsrZtS705dV/g7bzHdgZ8xkzXCiSRF8qcB
vHLUPq8eP1pctJ+JMPyDxQOees/oHIQfz/dUeronujNYioGVlCtkyjspXcU9zcv2lTzVZel0T58M
NK9gv+SOdCcj0nHWjRFPEyu0zNfnnkOOnhryCWtWmDsBfTZukEWpJRSzwrZ3tYJ1VCo1KariVlmC
UwT6SGoFvbl8+/pQ2Uiuqjp/Ujw0HzaYlvG1tODkXq7jMg9YKa7F/M8NRNuVnTYGxKUEelPSIhDz
MnZ3Vt7QTD0hKqWgsBY5uEq/WZRBA+PC+Eu8irwR/WhW2yPUtgQBviEAD5Lk1N/TSdDrGIoINbcV
bjru09E0bSBZe25caAa/1aimRueUfZ+hDubCde24WdIqKvluwsKjLazVTC0dBSgXWjtSw8ErfZWQ
pXqIG8y0Gt8P1/MaSUSGFb2XDSHZZmv4/pBTRH4IKs+8VdvftjwnDYG3aYBqH5Y97MVwINxRFREj
CX/AvWxpLzO2Rp9w2Rl/qhyGiftst4jpzNT+IDSiNLqwlZAVzldFeFFG3s+yVp1y+xEy1d4v/yl3
P0j5koc+MphK4KIssgVo5KlInQFWgUS5wu0gIDL9I17gANid+W2l7xwU6JEfP6EL2GVI3vKeyCui
tow9rAL2e8tmXPt93UZ37YDus8JgXbdOeYMBbylDWQ+p8HNu+wEi3XqO/UJYexC6+abAZfotcO2k
zrdR05D+ypU+w+fbFue+8vb8e2sTCw3dZPAbpGbiPEGr2VR0HXk0D3ZCpj4UzTOQgXd74axS4edl
mOUzfa8vfw5LWDayMKDhRQBoAQXFC/o1JfS3mQgyofwkoOWfPjFy8h65CSSphk2f1k6nELDOqKLp
uplcQ/Ij08pECcNcB56CFJhLm4kWQF/h6S1mKdYBqnDAmLFZ2l/NcO7OwO9tRnLAqOIanUNjVRSl
Pz3l5ZF3k/aEMt1bpo7tkxP6hSWNzyAB+iKQ/P1wO//T7tdrA1OpdjTVnRlP/oYiNWZrbSoSY8rC
gFsGgrVR5nmKcMExiDcsbNCkdeS/As26uM8DUerzCL78GsxsVNmd3asngbb/0IbyJ1XbGj+ItUTj
Sg8cmk3aqjr/+i1ZQ8YuDlvo578l1K2h+Gxk6lm2UHP+8V6dchdp3l7pWSAc3r17W4Ydc+WUHRwv
Y9IJEMQ8kOK4KBg1Db9usUUDY/ed4SYHvc8ds+ykqfZt+1KOhQmdVxAiWiZEOk6YT523XBo/wXqf
gjxFOVb7siR1SDGm/cem5ymSP1OBY3/Qbcp+4jz2j2rT7CQdVTVwuWWrk4VWDDoEidNyidRMy+Ys
GUXF/2JrhHex2O3UTMgIWa+Unv0nGeZzpF/8J1Ln8F9ijqq7iwVrSIeSSxyF95kgrYgR8iWA1Vyy
SYbkBen8g6lzVaIxSGXy1YuGL/o5r80Dg2Dge3gRLbA3I55K+MowkZRlaYxb4SpDdlzyOomEBe70
XRmKRrwnJIxhGhF7d5tapKalagGUcxqJsL3FsG0rK6cuezMCuw1dAeQmI77I7iMGTSApMeTStSCv
/fgvmz0PTaRUk/r/846Z6T/3FAn5T4kEEzfAA3iMe+GURlyNqEgN+BB7txXV5q8ObYAuUmMDheNy
jWU82fP2jLlsRlEkxNzbH0c8pI1hcx4o1rL3aIwysZzeLLl9rZv9RllMa1tMQTXbZwydNRMsq0sg
ib7FIv9BI6vSoPF2JKjyTIkbl/kS19eunsrTMvWUq473aDaZ6Td3M3tN5E1onyv5A3r9Y6BrKVsm
1PnN0fQa3yDxYLBF+t5iP5BWKTlHucfsWvRMG9bPEfggCFP96m2itnfyF8eA/M/2Mtk6oH7JAcA2
hJOCCMSgakhX1/R+FSYt6jPKbNDxB4gapMTKkYlNlmE8cowtVibUzgiuvLff2oQIEv33WK2uw/yX
s+1gzHwukGQO5rWka24xcQck5vvGxGTBVEjLV3j3Ja45U7l3TzPtAZ259pvKGXghFMQnLZpjekwP
C5+VKSSr/rHKfnXGbq2koT1evn+hroWlZ4t/Blm/EXagne02uBfVZfPpyrY5A0ekYiAB0hKv0VNG
7+IodGE1ztV6ghG4yi8c+qefbT6KLyqbmdO+Kx9Mci44s0JZTSbyf3KNKSzjYTdPNuVQBlbEUtzG
4nPTE1ZaMUWkJT4BdOrf4UhyYNR5I3qFH/py+TjBJst3h5pdpmjkbCG5xhyQCPb+aPFIDhb/yDEN
xs77E6N2+m5YedFIlEQDVet44tNv9LxyISYNZT442f3oXaObqShq07qZA7QQvCP7/KIhVL4yhjUo
586/WJHSlIjDkYQub9zcfILlDAb84vp+5Gcls9mNgpA+js3mEGEpzWjRNygBHzLjuz5+GgspyXKK
0sYoskZbdwPVcmMsZi7fsTlyW3iMikuI7ot/gEIx2n/yYik2uinIlWdRwM+JiS8rmk9ButQjTd8q
Lf5YxZJAfuH1HkBW3BF8/1lQ+AY6OaCMBo1hYTDNahWvqrBjbTqnzRNPhZlbIcvrAbhi8wDvhYoM
sYUk3ihzEUgw59RVO27M+cXX4CeZLcpndtUeX/frsekHF1MzwR7c7y9EcDy5tITTPqqtA99TvQg7
nxoRECigWnRUoBNA990etVOT0Srw2ZRgN9dzlG+1OwJeES1ybrvb/9XmP31/lU6ZUQb178iTFNKo
eIv1aCQk/4vlp/kY9VVyUQ+p3r3a5swdGudiL10r1FWLsI5WiJT1Rg+FqMyLVqv0boU2arXKMuE0
ij/fMgnSAOO9kLztGosrks7DGMVscjL4IOTY1b+ZfemArq32A6v8ihVL5T8t/cYluDKFbPindCj/
S23Nb+0chydn0X8WtrmLoJE88rgkZuaIwKSI11n5awM1UZe7ZlaGvxmHY+8c3CvGiul0NmYJJoi9
g/HIV8SaVTj5DSdaqHf1aR2ijJOYPUMZ4Uwh4+0GgWZKyuaYMkJDj1KkNBQ8gwN4PmjowVIjlehy
2rPP56q92LFgwC5KqTABc/dNOEmztnaGp7BlCPiofP/rzpPX7pZCGsUKiHyMuJkd0F8O5qkRewOT
Xq6Ix/0z8d1d1u9EOrvtcIXTwTJXQhyjZiBKyNfxJv6Gzl+0cLeOiYXcKtrh92Rq7KhNayI/8byU
woT44aAxjKENZbBEmZ3nUJ1hwEkYQ8CLIy0TV1HP5MM66/xFS0KRc8j5w++aV4Usnx3cOybdsFWT
Zq4pYc1J5cVqRxMnw9nObCYUX/HGhrY+epgfjI5O9vgsDta+PB0HZ9ssoPuUAKO8SI7vKLO8Lusq
d+Gp7ZJZ6bY2mb2mLGI2r6gRsKkME0R/CY3JzRjpdMxEj5wpN4LoFBt83FR0rlj5nWAqA+WE3DiB
etNJoHxEHWushJVCjJrUI/gTwAEFAPPGD7HKuaaTl2VAhrpfPw1CrDbuJEOonwhjtK4JjVEYwFCh
e6TopjnvDZjfAR0JHXQ6ECAkLexhjWFRMomQMN5pjMlY8QN8AvQzgs7RE7YCcX8q5nPEdyWYGmFU
kCAQDlZt9sC/gD15Ik94Is3Ohch6w6CIRzTqxcwqIQAhdceEoKDwBHpNox75+IFX/htp1puxow31
Wn1RYYzulGJHoyzKQXlSzoJepYyRApp6Uru3qvFmSjOdieqwaNFUghu4JT+rGStcYxsbJUIUAC+M
zCzItNC2AT5opitKoIBQwISYHU9aANabyCi5IGe2nbByYCWA/uQdlCnZu7Kwyolgm1XaH7HRL3wC
ckJJ9SmyNrJ6ZhAjBZlcifyEWwlqtqd45P3lts2kEgdFYDyOJK3i3ISLIVAvtcMhms03CIPuJSGM
v+DzJEPe/kCNnJo4Vpwwm88bMRbCLAkx4TJc+1OLJhsgLyNucyGl41GmpNXlKEB0miDEypKnRoee
/iX3XYifpuNcv5YJXV9oUA2X3I+vZsL0kFPQS8reyq9GS9WKwMpI8Y9WTnNOcfXVsLr+KxvrWTf8
nUbqBnhDYZheKhmE1hvGBea4c68TgFoY7kdXn9QtugtWCZrR/KJ4kQAPUAFpYOxQoFsX+Tonektq
EJsqeWIcKZa9P0+e8ZFn/UHhJgIU2ijPAJFRkyR5nRXH5B+aSKMCRz5cgMtvz+YW4l/jrSyA9quB
KRmhU4atNil5sJlWzQtJVqfWei3BeeDNJEpruaM4DeegZr3TInW0X7QpGLDP+VJ4aSnvEhZGGCl2
3OZNHXhe0Gjv7v2yNN0CfP2PHWw6/DEQ+eAA7lrxTfJNJf2RC0YpR5juH7tcPSMG0buJ+vyWrVBD
V0NwSGyEGJMs3v8WjxmOhWB5upUUXE9W1BQ6cggAWyJZZcrnu7MaVRqvbRq6Xf862cdkTnAZ/TOi
NRwtMftvwhiako8/gzbdPuCJ6J7XVpClbO6tg2sHnvydGpdm3K5syRjE1Pl/c/6pnSWYKWiR5K1T
EPUIWbGUQAtsH58/ZvobBO1EC+PQWD+JdlMdFrVuqAozbf3cxVCC9Alw/FpD+ihlCjrGGnAdutNS
PELA/sEgejyXPFAk8KgPEogcNmFfzTxZ54hfpmsiPi95Ckv3P7mVQINkA9b/j6/tKzYp8CBdkYeg
eyRMqSw=
`pragma protect end_protected
