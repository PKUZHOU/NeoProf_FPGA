// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OarmJt1qLZDDvPVEvx1XgWYycmnHr4DeguUbCAFetXH1jXq/anlNuZtGJnAx
hszxQ3mKmEEWfe2QY3WLgvIqMpNY/8v0kQTyM8/Ekoh8dXrXtldNqjJoVUop
noeCrd4csIZxzRN7q6k1fLwzjto6vJ9cW/i/fTmYYj0grkduZYceegI7StPT
on82hHKC3N7Eln9D+4f10ifNiqOHXznoVVuHLKxZk2U9jcktq6bOGAA7exb7
h/NQaNGztXBzal6jdWNNID3Q+CF3KGrYwQXgdVpGXREvOipvs7vSE/eHjhGb
Tkr84Yic2R1FJBm5VZa94o3Q1j8lOeQvoZc98cvdhA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Yhgkoxs97hFkJ6Gzs7PUGXA2Ven/qNOQvVinoGgWvvCWhpF5NWw1IL4RRBPF
e8BgKwgXovke00/Ll2W+EXCtENJis0q2PGtUKAxR1BrtJEQ871BN5AN5Lr9f
CET+Z3ODymquWKFI7Mi5L2I2kZnQi+yDtNVzVIYBS9zxl9PEMgy724R+70E2
wnW1ONaQjtpklNoTR25zcrnDvkARi3Ri44NLxoeQOFqnRFcdBlTmvHi+em/s
kyi1C730gjpzQGaqPfZvxm5KYiZMtHjNdCiREXvntmw4B+MF1BiN9fZhkH/V
Sy6mV237yplSJeZhj4uCpPCkLjYYSwIBr/JjZSeBxA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VC2oAObqLPXxDem6drmuzJaLHE1qPR5szzxHhwiTgvwOcI0zfdhTTSOIu1rL
w3bKX7mXpN/LWFWxKYNwaoSG6XbV/sJklEn/yY22sXGhzQ/5TbclLL5QKxKn
qEJMlls2JcJoFkYNzssJnmS/0uNpyvNXMFhwkwbJpSwDDInzH+k6AdKhcwfV
7MJ1VAD2vA2hoQIjAm2MBOGXvrOOTtlG9zm2S5WUsp5n6HzWbNkIGO+tBoOx
8vhkdaG7l0NlvCO4vbVFnnlVw3Rkq/oRvCRBi8A20d+wEPEDHkCguQCeN786
UmPdSXbYbFAp8PSPF1357TYXxTbfb+uQzZ0lrs99Kw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lLZNqFsP0dgmeVdlyyPc/FoQj4yuVsX6aIMiUSEB/jPwEs2uTgmFsq+SZ5Wa
nsPOyMkkQ4Mcbz0CSxA2E7bmcJPwfat3y2xmQvH+ogsYGlsOOXPyT3khyfMX
dOJ3SeQPqE9eVI6/49q0JKZkoGwyPa8QbP+KANVu44Ae9pyEk2Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VQf/6HHIhpKVh8A0m+iv5gJ5c+gEAcGCP3XAIRderopZoPJq3xltwp1Umpes
gIQ7DzU+MlJ/BKZq2f4Dze8PhniqRHbYAk80wOKsTUsnyE6pnYY2ifY4PoHU
p3yQG/r6hHI6cDJMTz+C/fvdh+SmrdF80lcNY8/AszC6xye7ocUxJ0Y+gk7N
Gm/Qy/WbbbWYmTzV8iti4aVynm47ZTfLfZrcUx9e6dyPtAXqcg0qYzsZmc1t
6v7HfKIAFRDy1xQJuAcGrdQHyuSpwIekTPlUpgMwyxx1I1MWkrYyeBpsLY8L
BT6ovQm0brJTpS0skWIFspX5hWz/V/SF+lP2qk1b38cfk6PECwTclZJ3jclH
6PoM+AVW4rx6wG0pAxkEAJYsmiVrrFvphTrVDrO87Lf5vkSpBbhqpIDCuRrc
vDyCy5wx7xRPiZ6yr2NSO2LFMHuIIe/CNYdDXX2ENYZEG7r3Q3ejsgGS/ESG
ebj7wrEvaLEDQVSWCtSBkTc/mzkNs0t4


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
e0w+oWH+25JXdFBmWAucRhaeVQeOJoAqCuuUPpoFJ2tYRiwFKTRKFFZwDMbV
ArFw4NJj9r1fjR0Y+HfJRuiVc4LTEb3PNKmyUFzSaj+6ivXLJY3tfu7oC0/z
2u8uMI4zA/kNp8hM0MJXpDRGW5y/s4bwbi/OD5ZfA+d8dyocaj0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ys1aNFxrZ318cdOjrnC+4YYPP++uTBnMIixdjGHU2mPWaUPo2K23BZgdPOLP
rFKqxEERr+owIt2e4j/xBJLGgFbwO+V3JA9sASiD67q/Ar0WzYpX7AnCxNju
5Sbip2afq662sH3ibPeZ3oy1NsUWmI3VQ+BXgpZYOVHjyG3+F38=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 49536)
`pragma protect data_block
DskxT4STCvwEAcWVFERLwDYLv7vCrOu2nrW9lMulW3/YGX5a6RSdfmfFFVPb
UzIs+ZbZBJoYmBSBordupfRpXDem9jlIz0DgWaLDykkvtKSDKo3aXw0wXAZs
ED0Wrjh0m7p/mc4zUSHsCacrmbdaEjDCJzwrYxp9Qna+JNZBP0c1bJ/IKO1r
4Fql1V9iue9Mx94z3XSkWq9KKO9ofS+bzn7M9Ay2Qh8UHVUGVFkGAzBEIlfp
5YYR2mWIrwjoA4eBtnO/M6tKHwUI1wP9kiNaAKU1IoWWl1kyArWbCE4pKvTS
DjvrZZZJimIXawTcHDk9Gp2Rps4h1NdsajauyvTcejVgdILBCSdOq9e/Qtg4
5rfiJkw26YrH2vf7LvUepyWigBZw2hMttdpm+O2cKyS5FnbWqfiH2SSYbyoc
gVS9tGMlGHtSyw22lQqMA2XJ0mwF6xbMa6CT1yISCNDMGadD+lniUdH2GIMo
6v1GTExzC0Z1ZDpMEtkiipwV+u6Yps6S23oODpKErEkzvIAzaJ0B6gldIIBK
kzJU77wBZCU7ktlc0cAeChos8++IvLzdqeNsSApL0JanfmVeNYh2vNSB5mjC
zy2y2vVittBqzIHhPBFKBM9t/8GOnAvw/sh2EnBFxpnyk8VnLS/ZQl0AiJ/1
iu4JzcVBbpjgDY4h1I5InzlESDPrD1RCZhV2K1rAWUWoZ48aZmtk9ftnBPwK
2S/q4tPRECD8QE9azjyjp8TMiq9wk06BQurKSdSJwa9tMqZKIrl2jemla7G4
DDAr1W4KS6Y9OPDrp2EWkJxMoJr5JG79EY8AwtqBI7cUu2kxXPXCrtRPvexq
9exOVXUzVvsUBtQPhUVqAMi8gTZ1aKUZ3ZvFsz237xERaEnbWV2CmJcvSN7W
t4PqCMAgPHewUYVc8Pm1FL0ZFOhCjvs7wzCvVbTpMs33umTEWhT3S5JdvRdt
cwBHYwSKGLZE5++5OzNHK0C3iD5lNrfyQkgyskYfIjIowW4p6F2VNKNFGPfl
HJp7QBLcMsFyKf4R8StixoHfR4kbfRtVuFtqSsqs+Qy2SD255jOxGRxp2UuL
pMW+4EvFSK/pAc4y+r6NBoejQsXbe7lJorgIZRnAxnV9GZOSfQe6DHtb0QC/
RLOma9CaZQt9UtYJpxaNKj8o3qQtOK1G+h0/qgFcYMsIlm70h5zFPjz8p48D
Yqzl2AlPNwNaBdvt461nmhICsCtRc99WieK4DQJTSJ2q1Ew9m2sfkk2Bl7rK
SBXTZdbqpp0K0JoFpTCfvEhKK+fdPyoiJpjxqxF2HgwD6BKepTLpElMQ8ukT
Z0nok2Xm9FWMIQVBANgXPVefYa75H52YOGy/2nEfvkp4xrByvIYqv25LF98p
W5I/wzVb97vPSPNfFgNX9lJb1r57wdxv7bSUe42BgMegSbAFeFUYlQqsRoD1
YnB3DaPU96Mr/uW4GotaC4Vyu86vAmkm7bgxx0hefMJeaXsI6XFetq1xgfHs
yBiaLg/YM3m36bn3p+O+bZvRb6fZmiZ6jdAtmiLtn1nKO5Lnb9ZQxi4Gwppz
cgVgpo9vlK7xfYNWMjcRNlXi+WEk+Pt8cXJGC0Lrqmp3K+Whr5JTf6fA7bnc
P04gU7K2vR7Vgj1hgcCi25SF9DZO4v/ClkQE5EmCfItdWIFIhKfK4CDfmKa0
AkUEWvwCd0Ezbgc78PPNDBg89GpuvxOMPfTGfQJZKHyhlzw+XKjzo8eRMaS+
+34PuLPd4d/u/wK4Cy3WpyNlDUl0DJJ0MTQLkf0ZqLsLgFfMB1XPgY0duPIv
cLcZuOOSsJXQspvXwwXk41rwLFHPE/LPP0Rdo4DbsLPwqmzoriO7z2M1jnzQ
TMect3VxiwoIP3efa3G4DaLTGeyqlPBgbo+TWrsnBAAMktW1AGAFdpjIf5J+
+e/9A8s2vfKeop8TYywHRZKQcXkje5RDiwB3Y5oqCyPA+ltpU03D/7Fo9pKh
mu8eWt01uDvl0Gq0PCXFsNZONHMO1kgKWQoFkQI/UI/SS6LcmusJZ6vT3o7j
1E4kOdnhif1+DyLKQKovbNxfkbuq1oF/H72ZLKxnwxn/lYN+qNwFa0BT8KNe
6d2cJD4eacNyNeUrpvA3IRyUh+0LBd5mC41NiT0oUtFG0sv4mVLHRUPgnNSj
wsZ1Pl6MiRUzxKpIIVPrt5DGXzZehUR7/pZEsKe3dAYusv0YePlgGRqZmzXI
lSdyf1mmN1FyZJFa5UnmJ1iw9BN+rAnqNvuzCanRcFf5rxQbCOtsZuoX7vow
NlgCAwgHqd0rhRJHRaWdMoMETxucOdaVgotESAeqo8eI0oeCzu3zGWkjrfle
94W8brnFDYhGmBRrh6TvIkcBay3brAcMaB+rsj3bwWmmLP4+wuKij5t5YRCu
vstIiLHdnHl6noV5DBFgzfQvfBxieMbY8EiF7S3pegUmesMTpKtPUE4/E3o5
iIbSC9nLWVvqY2NwxpAtuc6hJk/SBy27x2r95TroMxFOZ+obMe3hZXDQP9yN
/hJApklmNYDnuUa4QJ8zoJzABjxfSs1iOLbxf+VLrO2cnqjEkSeuebe6o2JK
Jcj49UF8t6d7OITIjXqQ5MnEmZqmYSbtKbSirRH2tX1JCDEBstsAOWOTIe4+
7HUuIKE9EJWOZDRq92eVKN+lrNm1pKrFgIy1rxEt8JmyJMPXq5uFjMBz8ISB
BOGpcUbTYOpHz9fHFjVK3JPD1PaWjBG51ll6MhRz7hyUYyNkGKkOB2ob/q8o
0Lk5AZs0xjkjGHYzsdypv7qoZ98PWTbHgVz1BxzjEzWg9cEInCaIF/fZckO2
llA6k1BWapms3LS+Qqs5mjWsMIdJ72eo6w8qU0DBgI+Fjr6+F2gv906utb9O
qX+XyYZ7z8i8FDea/xdK9Gfz88JMkxOzNYH7qoDNy6exTeUkwNyg6aW+/38g
BRPD4GV7lxopeoYZTINkpW4syWsjxnU8kgHrJi57i0PZu1j7qgAW8AqaCO77
kj4NOIllQaqV5K+ZdIO1rj17spOGL82+RZDS0s+AmsxuFCtVZaqBwe/KkEfX
lC7f2HonOrU3X6MJXYLiJRv4C48wcOyFmHbSWr+hRQahnB1rO8P24qqzbhCB
lBH8BiV5mOStyzAAtxUd9R6x6O5PndGJQShAPw2/iPnaiPG3iEnsTauTQE/l
10NAdgvqep9RMTwzmE8M+potdAmvMCPJTSxdfd1Mnpsy9Gznwu762GcytiMh
At59SviiiWfZ0rVi07OR4V6KW7TGZeMsC/bcI6ZVVDlSpPrFHxuiDu/a7SOs
4dfkCQ1YNDvsy2VGKBqfs4cPKQeP7CdYUcp1DZeghTLdvndbyAxXsftpRJDL
fn8/0BMTWGPK46lptFQTEvdxv+WNG/pSx/SqmvHJdRb/LoUYTlfchRAh3mM2
MvA2sAd2fbd0qnas8yY/4iyvhA0WCy2qxy6z2rHA/U9RXUcWXcySR9C0De/U
QDAi7nykyQRdKYY65Q8T6AX+3GewNk9u1m5CpoBjyQ/qQcpvtP0X5Na6WzBL
yWc21xsfgidWUp6acUst/6mjFgF6XZmdom2VN9nkdh4kAjtckapsoiAByrFK
OruAgEucvI6TF2mjnqhn2YSUJgbCFbdgkd5d/XD9hf8rBDNDcMjXMaR0A6+e
3i/obD6RZZrDCkfHbhYMKJwD4SztiZOZZ9lEoGsfKIsvMSLtH4NDHjFtotYH
n1rb8VjjwXnRcwuIgIzUA7kyBYKeavcLxMT+4nxdSfwJ8Ronr8BVXRH3/PMY
3lplQymsxcQ9J9tmIa9MH7iiIxriLYxN8k6mP0rlgpIsdoOeGV6+ITCSGLaI
Wo3YmScHIsdX0nfiUmVVXPGZ/UN+8uHt6MH0l4DUUbRYSy/qmO6hsEk+kR9/
KRb7XR/I3BXBce5x5kIXlypkdgPmPLanSllzq3YqInN2V1gK8znEO60SlxhV
hM6QmyVv7qrpNYmcrIgg38b0p/aBTQucujISYfYkU2OlXYb5C4ust2E6QGSz
pLlhIcwMBI6YwXO1tyfrj8sPquNpTHEU24WMUZUPmH0SVxpGFURb5p6IMlJB
LKbLV0z4OAaJDQezf5bwJc7jdvJ5zsclvPWOwK1CGhMDbVj/2l9ELYbO+wdd
Cv7Cs6+bBdVw2d5THd/fo+2CqtgyUJkANU1t5CbY/IjEMQBUPOz8vI2/z1UV
kcV9FHS4dtN/45DuhpSpdbVehjBT2ZLX3Av4MIDxxKra0bcmN+saalqS87PH
nlsV5+hRI9InhnpjmuQjwnivNY48jF/1d0gCgWYro1LCz8/c6agHegCNh2Ja
0m7GvvHOPZe7qGWY7scj4KhXnUsbQnBY61DP/KZl5OdqlqDauXCJjhjVpzv1
iCO/YYYRJYOQ9fo/cKP4wrGBmBgHa6HSawLTTy5XIHNfsIp1bRPHkGXrotFK
2dLYzj+kG4x8T6NlsD5G/gp9Nc2E03jtnVV+tEdQ/xcyZ96wPCIq5xPa2bmF
lQK6izrMjamV86xNSfaxOdkaRp5nusNr/Y5HZiJc0z9T9IasZgquR4ufEU1F
E1m109E5ZlSunubR3VAlYVWsrmuyXj9t5LnOwgYoQ9/RE+i9zQjde0k7TmdM
J/8N+Ydpn7S4a5wOsUWSNUprA5fv+oofZqXemaqfGRJeJqy1O2QgMVZIHOd/
kUpSp//bzZD+ucaGiXZwbwIGRKlEjjNiOQNq3jVYQ5KdHIrP0N+LElf09nqP
qGhFHqVfGMvvwqK4uxH3s6yi/NwYxs6loYrk54vZJ8P1d7bb75NzYaoh3rQj
pj8r4mdZrzb7ZUT4FpvXWMaM7Q6/hrWEfACDQaBape5od5fujRHbgGTshd//
xYHEkdQrEtuMYDmSe9UYIETeZTiTHrDizIZcxhZ6gM0I2sbCSo1rgDv1pEb8
IkWbUTfsNo8I6gWn+oTWHKcvhczgHKo1jatFiWeRaHCnPrH4E+d56dzjQTUq
pzsLvNO/Cm6w/tnzy/nDr8H2PeJzdQ5jaWnrdbM/aGyg0VYAIcwIITFbsVAC
xSWq1QgJbFvlrTpNwVCDAEMj/C19lncRakAk1GXIVXT2N8q7vGeM6dSmTvUU
ngEjZbsfkKuO/1kk9jLFilpvDKg+V1M3vzcY7W5Il627CHQCanuHY+0iOqKA
44IYNIJGNorahhjDSyYF4w6YT/4Wcvx3YQBWkxVQyej35CVE5Fl9nobtYipy
EaRyogLt2/q0vHUdI2Uvz9tC09CC+co3CO/tmG7oxE8KMYXVrChw32wGPFZt
87Dy4zhEonVXjleErZn9Qyh4lnd4PsR/aXw/dLbVJbDcJ8HFMTL7bXPalypN
oR9Cf/Lvw2iCExa/RAqIPLZz8CZQB04HQSUpNUB5WvzHXtNb9l/9ehKBkOaP
P8QiXXWCSEL0sOgjqsZtohkLGtwxq71zZEqJLTjThNRxt8y65ngOZaiKuCfc
w13/gfcNRuvRT+xh8tdnRxiW0cF7fdslYYekcElr5/DmMFCmr077ucdmMpJU
QmGLb/jeV979A1ye9uI9Z8JkGurhe9FpTbB3wJTO8HODnNuAubVKj3LpM6G8
sT9/lmsqtDg/5PA1FlK7std6ZvpPbf9aCYc85Vvz9m9H0np3SvHESwCqz5DU
AabJFw+XHgC4Q9jl7IzeBzQkgQ1wjzzdpSXn8e1sAwR5mzBxzH8uTfhrHoS3
hFxkUup85r5x0vxLipJ4V7hox1lcRyjA6Dg/YQVYHPNeyiv+vnTSVjR5IqpJ
hLVhpaskbaXPA7LZ5IbUhibcLXWYx0gONRYUtWe5JHgAIa2XJEw5kfFilQig
eo45oGQJfKC/Rl7ge/SIMCKlPEOEnYxQMxIsU0tcs2buViq8/NWwSaTywbPP
d8vMDMXoNWlzS0IhEVDNPt2jX0t1fRXyZjb8mEijrPJJ0oJIppKvnLiSHWfD
ElV3MCZp1gOx1hWsaeFAKjEJG7UGkBWG+qCiD1+X0C5mwUONZ546wky1BrBD
xl2+bcjBTCLvoZXsWevzLBnBByuoFsHCCwQAEA9o3HjxhjEczByoqq6acTgl
p7QKHcO+f+qdKGN1JrQ5/ee2fJYJnA2MZUfWizvE8NqM3vyuJYXCaTww7Do4
UmvWLlajIoXm+WFHOo2bHIfK5cRihWDVfH/CT4Nw+NltBy+2i6ywVx1nxaPt
bBDKA+AMo3qdLrr7XfIa7p2NirMviSddhFrhtQgEGaAWEM7KpzbAz2ecMj6k
QNKbzSinXViru+CE9KSNOc9w6JHtV5C5flcyYyvdRRh/PJ46Qhk9H2VfSr3I
EbSgIu7WM/4XeSS4bjGvON2yGf7VY+NrlwJtlAvhrNjpZXModsXEDad54u4l
0t+XWfCUin0sb4sJ8OwUEAR7/CCjlwxYGX9uTpFTKzWAFOHcUAnHJt8cS74M
Nbuf9B7ygTASKTex7MUDUZbqwNVlLqyU5COcQB1XDi1MMlImSvZRx5yA0r5i
4JzKlPFfNE1m03FJSutUshz2m9jOqlsMRuBXX5GllNR1F+CSfCaIZTfPHFEB
vtMjRR0VC/VGlItwYHd9fkiFYPgW4Mmkcs2OA09BLchj1udjXoOuhaLnhjRi
EKqdKkvCwuHYgOYqzCVplRnV7xJOw0v8Z/esbwBu/RYBUZvAl1cNOKLfiWxl
tmPuUM9pSBhc/tvazL60OOZCbCgo/TOTJS+LWesD+MiwIsyMljbiwU69x409
zIiXVynYRgTvbeR/BUe6vLeYPGggHNtpr43m4G/geofIRXVNoPSkSwIlsZtv
vkz/tZu+iYzo6v+rc4J+WZe81Q7jqyejslggZjgyZ8cL9ZuF1kcKZneQAaLR
aItVkg/98XZftpsmoF7up+efOdXKoipgb+sPWl3zpROptRbKHWmqSSAIhL1x
7QHXihbhPXBVOuvSWrBxbIxOTeMQwF5uqzGb91+6YlTURQ2KakaSULLNJfZy
wvXDVEkCDjxiAvn6rwTrND4bbejTeu3UtSnIarqSj6Eonk4xu7+gHXVb0mLj
swaoc+Y9QenIizSsZQN9NSOcd4n45EVXEmrOENEsJEa0MPPtQevyTl0GWyGg
BMMk2C7nOlte5gLYgzgArfl2RDymAsuf8F3CPrWcjK5647Hfo+cpr0hD1s3T
bjR787OmqCN3J5N7yFpMT5Zja5TVUI4KlfYswvhouSDmKJY2+iWAGIpRX7Mx
DFuwnNFSgTHytC5tB9Nd+zh4UnxP/RhCBUxLIYJOW0QHrN5kAy5kVXlEuVGX
8nDN9Q4jGjt1lQ69aPNcjSibOr12DMnS6Oc1VJKnd6CLi/BD10wLmM8PJlz8
jbKlgbkLFCSl84uKhnRgdu0c3FJXccZUL9ntaCdHwmhNj0/Ywx2WnAhl+tDR
V0qUwDnvR6cWxj8Cc7/so4ISwxiMTx469rujX4o5GfakYZbxjdTS6NrFioH1
pMR+z7Ol1s57sEdP0DXYWzXahfEQAvlUA50mU+/F2RcRpArUMCViGoKyVp1S
LgfhrlPqwwi37lK+gaeMyBheLOmwrwSJkYVAqzJThGgZCIELLfS/IWfXvN4c
VH6ioxoI5cwuHXzGGNEu9gXUd+Pb4eFqFm8cqNsjctctwEyeUw/SjEE8E/tn
B0hqoHJi3XTSBAft4OjQGGgr+8rzIEiC1UxjDmd4XSeNPQlEcJL4Pc7qkd37
nJ8/wMkAq32AwXVFYh4w5gCzD709/fLRxFwWjNXgGWdhwDm5EstMHYIXdbR4
2MsIMUvHGpERcGxWBwhoCOTNCmqzhgqjNe0sbcJg/JD516tsjg76ozHGpcSp
KsXyeVOtipFRdhmXfOVSxKdHMKBaRevejqJuiU2E+QMCCzBIyH6tcUYpKI93
UXvxij+WKRZGyyOZKZEvwuZtlbJoc/LhnZvNeS74m7m+bg6lYgtOv/kWDO9o
1wzOeGc8LC8+xq8WizM+dZiwTaXbDtHmOVhDxBUYEQO8JGV5zGj2WblIF6ly
s3tRd1lzSJIETbdcZRj/ifrsekfKCxkU3za4xxfSgSEV47nBhqBiIF1o6jwk
NKGXMoLUXpAC6fexKXvqlbt3S9WIbJiURCO3cQPSFI3zNPprzWUfYeaR1pqx
M2CdEEPmwBkan85zJDsKUCR01mucncG6+Q6kFKE4FBGBgULkgt/dLyvqzTLg
WqOuCBiHu/xjMVapkWhYD1wu0UaWyaTcsQkxLiznFBqFiZ97Ol9ZJTTNuudM
e+eTDF8jAPkJ6bB8FXBtesvXQ9F/2SRHkCFt2aI99PvgyGNQPScYJIB6Czrl
ZdPAwtayr/avNYdLWj6ND8a1WzYE0x2reUKsfsg89dPxVZJqxbR+6NmayzzR
su/Ivpjr2iz0mlFpnAWRbwR3vwDMM62agGq+5+7h8Bernnn2UC9zM+33tADW
zsRDGkPBOziFnIkuyRvGehwjNGTV44NPutxnYDuvKvhoUM/yxvxC5bjXfN8S
snZT4ZCdP1qiYWoTnrqZc7X55vi2fqD6GIx2kFdyLiQDDwwol9zrDJl3xnnw
/v+42XdQN3lPCTdwyDBEpVV3gb0su0BcYUn7lkocumLRjy179Lm1cortzdAf
uUvgLGRdEoWJBFqek1c7hXzb8mAriBRsOwgLfEX0Jv3xOAMtkCoJDtv7Bkfc
ZrWwYYrHl3my3N4xGQfbWjzZliSYhnzWEyfk2QIyMioPaLILMrlD2kUXf+F2
y13NzgBF34Ql9XBBmrXxFdEHIwONeciZHgymG+Fg7whGxAG8s3lxXHSF87n2
00ZEhDTndNiS0eJDWFOLeP9mg9SMR/mEHZ3KQccMbihQKdL9/aRLbheZiskI
DWI/5lvTOyaKmOczWkkPkGAG2boKXWLMvQwWeAWGkCxTr0WqJfCBOtb1QKvS
xrwyasOEd+TuQnKxrpXoH68qJSfEyqWhc3QretakV8AUPN4yVlR0fCWCitlG
GKa4x51cTcNvFm/flZroVvAGH2QQFFp1Y74xto/zeBVYyDNlRE0ldibku12Z
gjzrfySszN21IM+cqb+SXrBQ7ZLCIgwfqdJ0/HlS/2G50EN0mWXOoK7HKq/5
rkHPsHiF/aJc8P9f5q8RrJ+16PQ5aOE6nphDrtKZFJJ6K/g2h/CVoTrMGXZV
3Dz7NyrzpDWqJckpzRW4aMee/Re5mQARKqfHrZkoIGFW7cxasyCiLsnbcc4c
W+F1tdzuKrfJVQWK1MKgKoWc8DJO61lcKoVozIXxEB3dXOCQ0+xbZMgYGpgE
bbn2v5fnCfQYxfj/46d3ftAl9gJFJiFV2qUYxzZmnnYMtWKpY9IlDMwTPeTz
Dk2aW7DJcp8HTkZ7kvZTcTPxLQlcwcC3cAg7WWKlAGHvY28H+oeJPu3SGuZz
snh4gpi3HrqI2pugUlBPwHAIro8YRZL3v/EakrOWKYKjeHyqo8nFhckbJ8pZ
uTVN9RsMHAv8xWB03FAkIgGuFpSAi2WIdXlToYf4vN7IOWcq1z5f2M5EmPuG
gjka3PJD4K6GUUKTnOmzoTKYHGM5XoNHzmYthzZCiEYS9jnjLA2keIAJqJxv
x2ste6Cl5YcgIlps7d+EO10FHK757gizozrHWP23EpA7zFZibTsXFAIVurp6
J4oBDpEQm94VxBXMp+AhhrATKasWmcLo468S1TQt0rfRUOUQGzT77dRXGZW3
9JdDcokhChcaNiVldgUL+CPFCGFT5WfRz5SEuqrZYb+UcT/BfmCF8GbPI5xD
347egsvN94tu0v7XoMZLdsy4GWOpuoFemSui+x1myG118jJ3GKg/crZAgQYd
wpWrepZE8YAG6GJOFXDUt+lleXlZG1aIOhO+WTiPi7j5wonZuvAGO5Ja2uQ0
/+p4Ts6e8CnnTFh3ON0ULCKBSVWD1I2F/WznhYnv6Ttf6++BkrdKWhbTpEPp
Q2rvhzWJOr9AJt0JVGkhDAx1XvFJVPx9bFuq9H1o5k5flZatAlhzUHzkv+5Q
FC2ApL+oK45hK3A5MjWl+m+9cxkNMXp+ZioxDSQQ/aMUHtELbCCTg+LCEPKy
m8vRMdKwt6Ftdmrq0xyWkI8+6Yxru8bFtBnAyhMDCzuVtwZ3FWbiTlx5MFh4
elsYHD98SRPKC/hGj6JV0wYWOkY27DDUSMpQbGo411IrlMoalIfwbaFBAkhq
SvDbkIK/s+vPgwOQXIuMgKxixoOgn3T1kRFfEMr1gZ/QdrPv9cpDHSPUWxV3
W41Ns4UDP5J32LmahWPz0chsd5CDNeM8UUu3iYAdTzg/BoCb8e3oZOHBOcpy
KWU/rEuUJGmy+pxshSy/l1OoX0qq7TUk7LgUTScUtnSAQtwpIiU5CWsu/SUi
N0Vz6YZo+FXv+MXFEJyMSQcHw5cZOS0v+4WayZCILgB50sgwpqrNXe0A4trR
RFkhbY7+TemT72J7TbvriCH3IRJ4i96rDB8kWVwOYCWXEU9e9JfrxvWX/QS9
udx8D0YoW95owa9Bt9Qh/lr1+rT9JKIJvp0hCnHwU82/4lZFroyLX6MdjnRQ
T5mY5GmrPyAKv2bhDvV3toGm6dlBoylxqKN6ajn4BgiLxPrdWdIWs+AxZ9Ko
cXE9Yh22V9I6QGuT4IkA1yIFVfbM9j7I7me0NPaFTarykDA1bb7je/0mDgXD
Y22jwCXYENghvxrw6FQ0bc4AUqGZuhIATYs4LfnyX2OURwwTlT0Ku48Cj1uH
jojtQ45xsTLwhRu4UsWVUgnhrLBH5ncmm26FNs/vliGNppT+qmSQvx2dwgsZ
hklTsktbgD4jBoeMmWp4xsnLl9xeYrQYjwAX8hjHrst5kD4va55VuJFMkp2R
KIDQjN0kMiJs16e0wf6CuGut3pPPS6d48lZHT2mqX9bzsphrQt6SG6or+UHv
5HrY6iO7ur1NLi5RKUdgyePyErCcjn+5ADyUu548tscvlpeP4QWNPfrpw7pm
iiIOPlEvtYCQ9FfPNyt1p/VMhhZsd+fHcnxkkBnGQ0CpW7Jdtp1a5Ev0Q86g
K8iZLxvFMH64V0U0UJsH0zTVkf5WI9tC8/0kmlPhWlVghpWcNES4WogHEiSY
41P1f3Srn09iLR1FvqCA6FimkTKxtDbF2wfH2abd5mVJUiTY+XRkcU/FSEdh
KnC09DySAvhzYijZVbxj6B5nVjFLmqc/GVtEzKux66CxAmuaY7HzojVPlZ8Q
9B6Q8T9iQemUnhXmXj9hGUA/oVAddma3rcPDx9ZiPpuh/NChYcHy+/BUj3TD
Meg5TcY6vXR5sKwo8yIm2KKhiKr37ekxcP85MgOAAmevur3cyGAmROuUrjpl
ej5Jcc92EJiysWuIlk31R/dWZrRtjVyo6xSbrPnEpqL1T7RAd6DwyilmPvO1
aUpMER1pK8SO+/q9Hm0iJlCvLWM43WIflfksvPA5ZleAq3dxZjiRq6mAnN6x
/edFuPcqFDQUSYbmCxea2CCU0gbH2OI7Ye+1HrOu5GxPWywZnpliU9Yrv4eE
6kZRx5ToDomRL/yqQEFLUNR23FCOwWGUvq8zokK9BuSFGrvqqwyWMtRHirmc
QANFofEkZlsF/1Wt0yDgznHVkYfm76DD5bRXUrIFzT7VIg2sk0ymPTLnlDwu
xVCmJaLmOi/9mK+BJ76IbOkLIVSsvM7znQq0PkXbVMDsrfR+zmdpSBtSMtlu
tpymrPwLKByGBbLi+jkrXb0hvc6OT1V2Fn0rMTC0mnoCfGWSzisHdNN3A4Q1
LbLsZryCZ2cT6n7UT9sV6D/7O28QPpfI6i2Lb3+J8lhzokGNa0+aSyNZYJOD
6xfy5c8KgA1yWTtXW6+/0Q6Y/p3QjZ+X2MJCREbCap55i6a7kNJ4b+KtW3J+
VewbzhlVYWVDj4h7huoitLjJwehs5c9oTgc2Q+RdzKUDqdLq0AD9ld9CFP16
BvaBeEjYMqNwHcpeH+h3mDMNc285oZP9UnaytDJYN1jEbR1/NwdfjZaYKyo+
wTCL1LhQBqHaTi+4lKABUWJ9We8D3yElnrY5JcAV5XWlNV//7f+gC9VsYht4
bex9kIzKtd0BFUY+DxtzYNKsiDZxUSipIzrx4I5Vg0t9/R6sgcbssmaBs6RD
J8W0pd+eNCaz/yAdZaBaIzZH5zZnpU1KtWGG4a+rL16V/U1ej0keYgRDCRsf
iI2krPTyvLOEkldgNUAtd/Z8yTu/rsf0p0Va/6oEyLtSkwj3gWO7HwMoNnu9
V6Aos+LF6ZF+fPcZCrwt4J6zZQmOE1Ex4Nqt4x9dpjEFbShp1vxilAsiWe7F
aIIX6wRgunsRWkOJritDtGNmkZJOk3MMRAYLIVlCBnYY2UArsnbHrXG3MffD
XkA1nljws6e9mHCR+Pu3aufvbAzHsQBnS9yIigvEYY/R65JoLRk0r7n3H8Du
qZ4AM212fETOS/o9VVYyQIUqLxhnG9B+PITuKB78k3JyOll+e7P8iVxVeZ07
vru0NOc9UeS3gvrStNooTB+JsMvU+dATn/Zx0VKFDOuG+IYhk/K4WH5QLIRA
kmuuL2BanWE9AdTcem5n0RFmv9ySaaVd0x2LAwsZbZoSgrNpsGkvgtc0XK3t
fqgWUGrHbaQcDGGGlSbCZW6SFTcrdEp9fIgF2Dlj5IhflGjuGQ64iMz2/C9B
38szDk4hMeqEXMhdS4ZD5nRHGSRs/6CSjUzQ969vwMfy9GpN3o7rlrYWZUza
bZK7oyOIVUDuRn7b/R7hWdC3R9cYZasyrz1895P9Mdgi3AjxLSXDKiXzTXXe
676u5HTcyywctU95gS4yLOXksNwsBtbbyfoBr5AXbf5ZJ9axI9L+2nzIZtqu
w8FsJbaqEy9yxUq9QY6JPhczn/yEIbViOWmV16n3OfhNtjwU/pAR6xVbnyeg
T5i08BM0u0ZCIx0+j9LbAI0OAKSgs9rOzOtmtZP+Z0BhaKK2AStTMiEuD9ao
mB2GSm+L/qQ4yUTR3OJClPLx5JcYIhMRTgr2UUto0SCBv3irQwuYZtpPLro+
eZT6VdqziJhUueVpDm/rkKqU6AkG/qp2ekmDFHanJ7PxBkyepxm7YZc5POuR
7SBl81omI0jNr2hhCLpbtC/aFqN0fevN7jk71/zCEmUj3izH/jQOVj6DWLGw
SJKzIRM1MNU0313DM4QvLjENZgU1MsF3Vrv7/UC4I5vSc7xl3fnqXWFEIPib
6JT5bfxBp6CPLyHI/PDJ23ag733/erkPNjNC0fceyOfZpky7VVWOpqBG+ZXI
06PUpANOcgEh8NdqaQGUEyVHRFXfchc61mCrYsjOYmU0mDbFSbnBwzLqOY7f
AW0/GZhxRrtX/r3iYCCV2iwr07igXLYVUAneyF7YtpkqNZ8Y/Gd1fWk4P+2K
zRp6SvHahUYGQ3DZsC2EJUd7dIpLClR+TOXqxQ2Ld7NNjfK7vJ8Vpoq+bhqP
4+T12ql/CgaEWbpXIhSiaDSFqxo4zhf6zNBizU2+N6ePvcitfbhC8ytNfQZ0
7GRrw4aphybFqRZECm5CFSYZW7ku3X29Smv7RRdttsBOAuolnA5+J5896I1P
HHisQ38QC9EjlSidtsycLHTzty4h/OweH8sWuJscKk3bJA7wxfHrXYG0e6uz
RRnKTHkkI+ewkF8WNaYAx06Xj/TCpoBCXrr9QqKb2mcsSn05crBnQ4zt8daO
sxIjofhJnN9FqzUAt+7mvYTVPHWwQJRTNggc3XCUwayR51yH1ZAdKw3w57GV
NKWa74VHqHHmz38Et6Crs4slthSqjpY7CY0t+sLPskUdt5eUZwzIcuBWtCr1
psWcOMvFrSgCAKtp8h9Qa7Ul75G1VaCEzP9NAsFq/hA57x7ChfsRmpkdhrgq
nrmidmF4cWLPzy2JmAIuXe2ia5BjtA5oHdSkj6/k9950pIoA9/Kibbu3QpA2
Khs5a94RssiOKrLm9M/4bjnBbnUJAT1PkLFTIUWYmQweNIEOIX0fb5cB+slC
3MQ+Onlm7ABdi0TpEVoOji1MbOra5DKfUN3gxZMh2A+8nnFEpKT5F9ggSrpL
/jmrnWAdZ0G4CASwjfk/YaKW6uazZVkoTduci0F/df+bhETUgvLmpd4T9vDP
fQ/3WW9LKNRomROjuL6dQi5cdyIbks8JBcJi9J1JkIpSTrKajt6Duobh8UvP
5ok+1XT893PDqDhA9aq/tPQqPtK0omVjXh7H5/jh46otQV8pw2tNf+DSc1I4
FJ4sD1WHU7JAntoARaTeKXkUcq2JTDOWPlBuNKnofJWGYHjxeAgteCjav9s3
7QW9nnHknn/TU5ZRwZ6VeD/6sTOc7fzoSydYBHklYbbvlrlMsus5tO2D3Mfd
jog0UHjDAO2Kf1Yp6OQT7yflirUZOCU3VGnqLzitAPCGjyySwlFN3Ma9bTNU
sMpfdWya1RfY0wEDm+hw6aT7yy5w1S2lbMZZ+OjbBDKckg1ftY/Z/e/4dzHn
Hl8GnchA1e+5plmg1cRn2ol11vEzqZUsezIZYEhbWBviuCVCh4i4FnS3aZd3
dPf8tDHKbPtcD1JLPlP9W1UB3IYsyxCZJKQi2z50vBtZZGq8hwf688EokHxV
PNcwjzoDAOa1v0Svjp/TEdawUevCDymJq0wIxVvq+Skyini1tc4PuG/VkvPH
/ay5blKwC/8yaO0wJgmrJHfbNlUK3ecbVQTpqMUcaeOVRmIct9p7VdOO2Fwq
c4H5HduqhAT9o6BFQjrVrd94/uplc8jRi3mHy22XzSaKxW4DtExtvXbzMc/j
uBbaOQaSB/awSpM9uRqft4FGY94uVHsR9JLiQQH1xl9ckRTnRF6XUGrSFPEF
DxlvTTWzPitnbhXtnhfrpc00El5x0yOAqMc5P5tQcFiq2a1Q3GIvUFDiCSRt
O7DLsi15g2iEzKxPY4acS0Pv8ZUNiFqfpHQsh7tP9Jj90Q0IXhFL+TzjvI3d
hMnA1vqvKmb3GvRh43RWmzs4Ufw55qEMTsRtZ2wk2SSUYeodE/QWv3hKjDl8
WViAUJmqLwE7d7ZMJ3hI6TQtBwZwsIfpFTRaz2aK3prna/xNIg6e8zYaRetx
6crvrGlE7UPiolHqdztBUc+6lReJRRfZuP870ezjV4k6F2aU0YGZVUzpAQFs
alwqEfQDfGcWAgWWiCyYRsu36ro7lYivQK35/29Y6r3WnBCutHKPSTTsQWCi
qC6gnlFWg0Z+sJ1+FIbykf2ogWsldODeJMZmwOBfgd5sfEtDd+ZmMO/otagK
jteh3aVJticw1QvCghomx+SqJzBaDwWbbvvqJeXOtoLi1WxjWFaKomaFOaOY
yM2rOkSONaFy9mcnf+hH0ajVzsDagiza5raFhspN09ippxMutWCUIEeBqHt0
qkZDgkN+7g+fipsi4CXGAw0HHCVAELGMaUopx67Ay/+7kR0Z7MenZBJHC4UT
j/cmrrjXMJGxXf5FLZRl3O2Cf8Wwv3jxp4NvyTMP5Vt7X0JWW8Wnx4s52Dww
KAUTKin3+ei1ZSUdJBcZUOMrSpyyPyBQw7yYGbtSq41K1bUFzTUb3BdpdGHa
RVM1/UROhGZ6nFmDE6eb5Fu58oAV1n5rhke4eOXY32a4mmM06/nKcPUPF2pL
sIkV9kXCFKxIDxxhvyKOCNBP9iYX5KIQ8Zsk+2ZhuqccOV5BQNHV+vXD4Wvn
iKTEuNldk1kk0a9Z1vQ4vgw/xUrqgRWZS7sx8dkSsJp9Ah5EF9erZWmyzZzp
6WervC7I6g68htqW3DRa/Gk7JpUp/b1ZMEr0nkg/ziBSBoOYKvZ5NsG8u1Ei
/E8RgIyouzQinwZzHhzmfrOh42e51gbB7vaANGh96vnymaLQGJw59V3BgHGY
b+A7a29vZgX8d1YWVdWlT9ctP4ywogAyL5TXq46UX8cj9QfEB/6yv37yhGng
z1jdpUi5Yhl5u/TBxwssZ4Ks4gB6+nzcU3EnUx7X+r4tqeu1DDHCaQ99nkj9
bS56tOyF6ks4UGuETHebBa/GgxscGg8idv0Bn52zSIV7E6xNXTdQ8eo3Z0e1
6zC1AIK7wPMSxOAIsGzoxpfh1/Tqr6Oz0z/v/cCHm+WN1fuubdrCoKwBDqK/
Rdq9TaJ6PMMPlzMHsclpqqHyA6x/LPMWV9dM5VMskvSEf+H4l8uEqCORME0+
1S/YFZxx34rQSmqSD8DLcZtvrrV/nZ2eRXbBAcHpwywP8O4Msj5tELSVj3TV
gJSByAIlXzu3FWTqhuwLnDAIxCOdvIK5wQU3Le1pnyUUDrNpqxRK4c1+Yb75
tZVkMShY4Am/e4oU/NUF3T+O6oSrCW4Eydcuo5wJ52nPCwNz68H5IzNKZlR5
+4UtxUWCbYh9Z+PL8yHyZ7xRgGrMVZethRTWIikx3EIWWstXjK7cW4FZjO1k
xYK0xvE4O+RpUcOgreGChe/6HW2G0BYBam7i90M6wv1xN+TuyHpW388fAwTl
SIXJVk/NyvancquU+uIv9kADeDn7FE5Dv74dBWewiNmFd4/eWqjtW0ARaaht
aPReCxKkDDIUJR/uhNogX0JbMyJGFMY+YPcfb5IGGgKmOJ2Ij2Wyxb2uNnrK
Gq/MtKaw4ZkgDFYw23o7HYxiyRcoPrY3cWEQBrV3CiQ3Z5BmgIxVJGKwxM9T
AZGhuy1KQW1cgRKUOETRPtCHfWLn1PDdMDLvBuWWIkPNkywukvIuApI8+w9+
e+t1JosBrrRYOMcFALt9u2kCp/Sa/G/UawYrN6QCFZS5FavII52XVYF70LXY
gR8+vSCbvBd8FiFjpgWPRZETtxY+tu78WSG4XrdgreB5hXeqB5H92Ay09RoN
1VJFtgW0Q+OYwu4CwsSoKRRRXizykrUhcyTHJlovIIQY9FCPNPV/gJVu9BDF
covtpXKUJ9UZI8lbud2JYVyAKXbcZWYMMJKgHLrDQwnBGjpmuQdcCMxcvilO
V7okTcA4hl/Mqbqx+9XCYcepWFHPjcvMJLY7HNRuiuYoKxAFTpwR20MxuPA4
ShR+mRoi9eug/ZnR+5sfb4FcP3p+uHnhti9pq5HQExZ25ap5eTVrB97Jaaul
1eopPu8JydAcNzFv34N+bwknlM5BNaS1NbQMRMrAdOj7CatwNt1GQFXb6wjo
oRRSpwgwVLrSdzqZaQxcewNY+DrGLCIYDO5V/dPWk/3fo/+Lz3fQb2oAOeCb
pRPJna0aVMPUiNYeyc/VAiSgLvUXCciJBi4EaCkFxpCfdPmz+pIlKFNh6txo
wSjQc4mJYLrvfH/oIfHPWcap+ZMsUdxN0YFbymuBeRGhu+J2E45xt3qNDp4+
Cfd69ZslMLb86D/qFstTnLDJEmGO77eVwYnA4smKksdQtMKIdxHRCAr9quTc
PgW2jmgyRZTwFFuv5w9fzscXzaZGWIR1tp9vRnaHdxlB8bsWwqqkj3DAZ4wX
3MEnY1Blp7D0aKOH2zynJHA1hlTG6B3Q4wpOjD0C61BmP4zpSjjPps7zUY4V
OkcwJXuervkE/wmOWa7JLq5rritNyx7tBpaWa3nkMU5H/z5D5C0UHf4hi9x3
fRC2OCLijMrGuxhLe2yYqmUpaAL8qByAl/qQPpb9XRDwpOzRGmR6ZXlvNYiI
mlHh+eCdmqvgXwfc7Nz8KzwHSi1rxGdEXDWppgsK8CFn079pVkkyFG6QEla9
oXkUGTp1DIB07xhlwUIiADmYJcsz1LTJkG2UzDI6HtC7o6MlxOOEErc8Xamo
+fP+vqLEoQoR4ED2DdAqgdwxQYiDEKQ39goBjDOzT+cefUQLINBXqDEgVjVK
nKjHLNq5ifDSYjg9SLv+qzOjwYxRJpd11CG+73EC1LGCOnnpT+X88IvagKke
l+G3r169/VUbZLWDUqsi4pX1HiDvsIdXg1vCpcpEcuy9b7ZSzvr07EezoYi0
JPJLpZQxMPC2qIzPML2Z4OB9iwFu7gDbnxRYqXXxhhUVS2+fXaKQauAtwqDK
WE+LBgnh72oE6bMOsswzQVamj0ABTNj9T3p1vW0IEx3XHDcIVBNW13doqgT/
+V72wEn0smDQKWi4PiEM0SNiTNWyvdb+cAnZ/xzdFFXFpzZwbSyoNZx2R5sH
tR1w7122AWJt3T8ymAyvL7QG8hgryWSqNOMqQd6+3yY1G0KFtueTT91qS60x
BMbhWAz69AKbdLwNMbZckUgUcXa47Ce1Ut8ThOBq03/amU+DxKMpOD8ccAEs
TIZja5fiuZjEIPtaYGy7naR/hzJ2ZD1br2Tbko4dH32Ca0AfBuDj9B5OSFiZ
FflOVso/m28hqWz62IO83Ns9CVQ7E7yNcYcEfpI9ctFkMsysGLdeltO0DdxU
dSKEDa1RwzgQxPYTJ54zwPElEZsRnjvzQkLQljgBiz6QJMPqNuZfUEEKOI/A
qsTRF/ZVokm0JN3BuZaWJ/P1ul0XBWpBCy1GuC55AtCySEaDDxdPn0hki0Kl
smOk/T8dmNHZphVU25VZYwm2fJTZJcShFaY+SDONHTC3emTu0ISYa0biPQps
YfoJrgtUL0V9ZGW9Z7klAw45kNbKSIqs/Fhyiv+aJeR1DsGXE6MvCKKqF1x8
EWPXFLRL5Yfeov8XpkFknuAzSaQN7X6MqElEjt9nWE5ll21FIpG6tRHjBca9
rfEQ7Mxth57rGjdx3YfhLGAtTBEFTuLQbLcuCOW2UODOfTjNIL9+w+VZXYeI
+J3qbwHdkw0O6oNmFOEpM56yNiP4nbKECOuzhOwumpdtzbMTuN3Nmve4SKjg
Dg4mzGKHTZGzzkjgP7mWKqC7Z3A0WTlJD6zb0e7Wqn0hgJ/cw0Httxl43rrX
Idi70PLBKVz3tLDMfWXN6Bv9EC7T9DUSY+XP5+pk8OXFgEIfj1lUsrc9019X
N61crEckB47h0emOUz+1JCKba5t2AlcPejLHCXrrMExDZk1Im2h14L+FJcqb
w1Sj18yJagrTrDx2FYksO9zPeJPmzwO8Zoud0YnyoWxryLfmPhCfVA7qEOl2
Td5gS6htXLsFUyGic007BY8hdit3rGu7aH4jrrmmr/KVc3GIBfwG1LTVjHAt
muu17bfoIz1pNcZ0zEMW2nQRiDKyOQ4+5+F63wAIjLf9MHQykWj9O46bXv5K
XSq33ZiBjVR0yYin5BaHWrdQQ4OXmld8K6vQ45ntEwFXz/IGvuCOksoNSIo7
ZP+YX7ZnPGdDpzoSQm2FdqxLH6NcUldcV5pze3TMNrTqrc0F7sAWPz5dytdf
gac3sgJlK395FlEZfNkp5Ba48P+KwVVYE3T7Q8+tJitN5L6cE7dMNiLwpsfF
rb8s3NZVFKT8Wa+1+ddFOt39fNk5882LLst6mYZqP9y/RxEubPTRnaBJ4m5t
1d1FBFkDBd76ApiiY/MEiQHE2uN+NmjgstWCNRQ9DkPDTYRO+yQFJR3OzBKc
03Wj47U4Io0s3Nigbe3YqCYnIFh4AHOfJ+RKzAEyy8kfLBBYWqVBhcwKyLkO
/RvZjUpJwABah1+JzOA26XB3HP6nddtmf1r8xH2FVMPZlwONTXVkRkvpzIzr
epq2pNV2mxbJRZl0LcID6kX8YJAMpcqwuDmFYUsa8u/9xrOvGbwY6RVAh7rC
YN99OPThHGSgWU/+zpJ/M0KJIysRF/AuMreCGY6Psdlyxl2CQ8Z+FEEWkv3U
LFn/wQIuyo7h/Bgm70QcbFW4hbMU/8gkqb831SG47IrCS5ZYEoX6JIQWD3+4
0k9TI1+maaF7CgJs+nz/yUniHj0FF3LLyxUwsCJ26D722hFQu6p2kkSpxZL5
eGswillGUwRPGh4YaEbpi/Ar65TBRWWYDcXmn1iF8ULvq6xCWo8cxr2YFhrr
AoKbQexeWNaJxVxwlWdq/fLFuv8J9T57xwp90j4VIVjYkF9Ih9CFY4Bxv6Qq
mfnjqTX5PFuXzKGefU7jHKNHBGIW9KaeUg6NDBpBcZ933fsxJxNhvhGBWTYc
h6McEKaETBZDh3iXcepog2EQjMlR6TiQE+m6yE3167uo4SAYDSu5S+nxN/L4
Un6FUlYihVRaaQl8kaCK0oRQf4RvtSDAl0hgoY/rgUIOofFsj++7m1ReFlk6
JSAVGqp2eSZHyHUE4IaamNJLMMG5ZiBv1whiynG/R6rXrsd3EUwQrt1q28v9
shCqjQI22CgeMMkvQ5QWsrkR6a7SvMXObr8Sgld0ugQZBMKcLAB6nHpwmIfd
DxyUADiR4R8/M8Y1v1xqB3wzXpGAlgi56B3hCJBeGd8ZLKZwA3ZbtL6Y+ert
QsQWG/ujmz9FOfX5lY33ENioG0V9SkeJUpW3u5kp9sqTAZk3weEfEIGZKYHC
phSdxxWWeDenUAxPyyA8F1zZwyQMBKr3E9byDH3yV0xdNnejyJs6X7PCqIgl
8YvfOBt9+7AymKK95U0Og/lC3hdcvZuLptWfHEmCqXxrN8yOpRiBfNEpQvTA
OwyAhaS7jCztYKvK3kbyXrpCJ5JvMe2hP43qKzksuGUi1KhpIIv8q1DZYMh3
pxR7qmpklwEft9rqxeac8ab3IoP/C90A6eHJVadVkBkUIppq9CT/QxHtukgI
zhOgkGzqnhiEXIiT8kv32tSfgJ/RRjGZW347C2ZOvlBoRxlvUtDlg16IDt8B
61quf2m7ciXHJqioaN8PD5VXGGpeoKhmt0wzSm7zLnzYP5gwb/UtiEM9TeEz
R7e9O2HjJNW5qf5gR5wqDc/nhtfjLxp82gX+7Fblukke40f2l5G36my6CC65
vyV9mHM0mJmcDp1rmmVYbSjEAKx4aDwTnl94QXx/jeBVd1mTik2HE8v6q7hm
LRXS7axNHuF7CJKNVDKf5Rb0Acmjlp+qiST56S8tpkS6jJqOavWZMC6+17zJ
+J4H1al7I01E1Am1Fbh92aTLqIgUuPXMLsQU+P4GiyMqvDvgiJOEIYEp1bzI
Wc13oUA27E6J7GBiA6czNejBOnB4paeHbIfcQOenQV4my43PYRjHuGpNwEPK
EFqY+YerFoWWV6eMRQ38tmVgEgi7OcKPkZTO7NRQPqmMRInuj1fbqsejdrlq
QGtE2uQSF6tJmvn+cOgwhOV5iQIR705Zy88oWkv0ZrNwCjINdrE57DDF6u33
Mou6bq+FU8OKJ3n5LAnH8X2tNf8ywv736Phz7MWRWtjHYa86EydZuZSy680L
MCFCT7MyvEGRl4c4Pk8mTnSrUu2BNKk0t22SL54CXCZ8Wd/vV7x8/onPDBQR
vCdzuRok6ZcpL+krD6LvlYb8Q188PiPISF6njju9E/i/OrVYLp0ImJlj+5Id
LNLiK/8hL0X+OAiLuLyCAEDk6vl/wVHq4AGwbluedjswXpOJ3fUhaeJqdzwV
XyE1k1FfDTJ8XRAwJX1k9q/p3ErpqlGPg5+EFmlRmUuYVeMsvb0UPM1vlEtb
/ktAByCxd4jKYmc9bv3cQ9PgFkZBj+FcxfToKunzPQLu4Rh9RIgAvM3xK3gS
Ph8N88R5nX20XDlo/ZNIQKlmkyPMZFQXrm5Dn6M4wr92TLhlByC3D3wIsWMC
7ehA8SO73yP8yd5SnSPEKpDK2wf1AYh7fgOsbJNU28835L85NxTgTUWKKKHm
cXSxrIXForo4Y1oK2sHG5MbWQKwdxBUF1dbw/deKZTEt+3fsXela5fiQ6Upk
u1tqScSm8rGqA1jhnWBl9OzerHTdveF33JhFY2YsqLr8hzE5ItQTSaN7zjYI
mAGgKL02s9sl7HQgMqUhwH10M0NpsYfUpa2KRgemLT06dPR5lYxeaw5iYGvY
m3bPEZhIK1NSZCUNWwfWP1AWCFEdPb/vIWeGhaWWgVbStTjMvt4PJmLd8qKb
H75W+JH2R0X3UEjJrRVVO/qeYMQf3Itxfj+26OYdz5sUEmTIpIk5o36BxsZ2
U3s18UbpVL0Xh2ZfKs3XVaVXSyQjpcvDyP7n//+LTIF1vjWVKxPmZc91YnV1
Wzex3CTnF/+skSERhE+hijAke0yczCs/3hGvwNkE+RQrRulK5in6FCUDNvTs
z7kaJocVDNuq21Mg/G+nNkUC8bBZvPPKxucLe807cya13JYTONjrzcyOaSU4
H3BK5v75BGQSZo1oka2IvLSbDzz4m5TSM3TlGPkxex0t98yXwme47FgZx0AT
vwQTq6bQLUeYBx31peaCaNl0eGH3GrPxdFZsdZ0UUpoaGxhzTbVuMwU30zJa
W19d3h1wWNC42G0IwAyLhaJ1sti7ZZJWe8GRt5YTKriRGrvaNx67yi2nE6Cc
olzjrWWVl18r06gHnoVa2ts6VbjUF4Luk0aUUbkout+FqFjJEnJiaCGDhbxP
jd+m8WN9tdkqOVLVd8n0xzxQ4Oea5M8hSF5+FwvikEb8+Vub2B+Ro5naZfcF
fObgA806yROQo13SxOjDeyYXlwkTfHCTrKyKmXNvLpK4dXxPZa9zNBwIFchg
1o/A7LUzGXiOnJikQRLV8qKuJaSEIPiVGA08MS86upL4W0HU4y1gncbLf0FS
YIh3BSUVuyrn/2sTfeg5KLODtC7t+QhTYJaja1sgH/9pSyXb1Tp6Z19vGTyl
0JluNqx8g0R1+TlwW11LQMRyegXuXx5GNLoXml1qTsWuwr3E7Of+m7ha4GdP
Rcd5GbeKtBYSRzAprMV1rn1akGq6lcwKeay65iEs33LlmoG4o2j/X2xWBTQl
cXlCD12rUp9r950uCQFYMHkQs7qu81tY2JOv2IoKowOD2R32h/A//PY/+n6s
n9mvPIr+ALrvfZkcSsp6cb4LxU7NDP13bq1nCCq6mD4MlWsMigGjjKboi/BU
EyvJlZGQ0ohRZ+SHxSkhBEhv0D6kRsT868vz7RuUWF+w5UgH9bwODuldbP+z
WFjyO4sZatHtt6Xot0IdoJZWqSTwiC0laejGNwcRMWCqEz0ETvitpWBjgE7b
WLKuyy48Qviyt59MHHA9lwxq75uVikNknK6Aja8ojbOjyLr8xUoo98tXYfpv
IIMmbAUgOXu2GG9pPDnyDFa5Vv5XeFsmOzmnVrksJt5GmXBssSBlIlSAF9f0
c/mVNhDr7FR7CwCBfoE9laJM7Gzl/5g5iOBFGODIEfjCJ7zPbrdyQDbC4w/n
x+gHoKKwtfKVoNXu/FL1BioejSgK2tbAv3J8Vf4rqqo8uu6Q0Z45YztbX2xW
1od59CQd5fSvBBMt+V23wkSkJ0MNL1YTHeOaY/KvEom++AwdrBhvRiaEdaoP
/gDr4KPdSdmJKZwq4XQzaIAqdC/bO90J5aDbMwWVq3/JstIe95x4O8SbUyy8
l8B5GqVrYIeQ1TLDU3YfBoVAe0ZgN9UgkTPI26zb9f08VoJk2eCTIDnIOIh+
q9gtfNhlePm3KU2hJg0Cql/gcoUrl5y0kVV5ZMoy7DdcyIgSEPayLaE3p+6a
cPLYK5DLnCKLmggzFB87o7Ig+ZEAfS0Xb7qLJhDA42jjsD5Nquxnb/LEhWE5
XME5+CJGw0TTB0wYk7IpYP/RhVIBCiTm9aY6HIv4SyeZFSLhK3jFvms5U6io
BOYkzopQzydxqxgRPJQqMZMCb1qyLOAvs8avfPjk7W5TXxw/Ks4svbVAWMFb
dJq+XYqUP1HmELQD7Nl6cFZaNujYh9Zp1l6qgj6meJO4TZhBKoa/2/71PZ62
/skeMNnIgdQcSN++C/jVXbNNjPkfgTvhy7Bsg9mk8RKYaBapDespfbeKPK9s
cd4DYpLg/mvKUmBIk1sx0Y2CR1jkxiEAjzMqfsR551/U/Fzc2QdxOnyfwXlq
w0yZYuHC8tRkcKTk/3e902YvRT33gMXHlIEWYD2C3UW149vXkBT5AHWFZIPw
eyz+73tsBLZNozReaHVuqB9HUVGu4vpCJZI/ZOhloilpiNND0YBufucF1F4l
nGygzguicBvDYRTeVgvSe0ZZtnkvdCIylFbL0B9rRiqsthqXjruyQmKds74I
oRpuyF+PClCiF+SDsjuMdhGb5K9RYIg4PfH7ZHXAGw69PNO8BHSapjT4K6zh
mY54yU2IRAmoaul8Qv1HVOXCiUN99LfEhPLkEAJLqOmHu5vusJuuT750PyqR
p2V63AGRLKZATjUHv4mofUmYlSICpopTDRJu1AaRXGbxfcj78TbdgcpGRZcV
IlwPEdel9raq0lENmGEM+jX4pXDP4Q8eEIWdlxGi38+loLOqdJk9VpFnoRUG
mrPr49AhrqB5rknLRsL7Cf0s27TAItIx6ajmFGmY9XTur4y7zMbWMh/V3kln
0uMVP8E5aJWbkoOph/3naAbhrZQAw/BCtqjX5D5QEMmN20nww118Z0xMjtXh
+fRxo5hcsP9MnkpPUuKVaGYcsaonqNwDqIzmPkRThN7b5lxIljjWNUT8Cqd9
yRjnzfSLUY2Vez06xPrLGXXHuqvkOAWWK8iG5bzuWDsCf3X0M47I0UBt8toP
Vg6qfT6MYWFJtPIZ14kMpqe8Z9rGBtOa6HGTOaJA6Srn3jWV7ufRFEyzf9/e
whtDWBQszIO236qqOHTz7L0TcIP2n315GUfNn+0xvSLdOmhxWjKwCbUsRk0a
waht6u/eMBZRZjr2FCjIed/cwypcmhGS0QzpRnaJx7gB4hhdAICo8rmLXoft
WRVkLyefeR4fwM/JgurT+KBzNqZVUC1yRLFp/ZaavwydWpYDyW4PuTa/NdYD
eQtvW36Bu+fxPkBmYUJZP0vi4DcZgRkUqdN1tfZxW+uUFwMcwvVGAdrx0gLF
FUTnLlewIlWybbX75mVgVFapguX/0VMQn2RCJHEtwHNYb3jjZy3tHP9DnF0P
TmOeu1gkwvLgHLgr+glo2QJb4vZDo3FtQh8jot7y9g6i2WUznDb6rGWEorJY
Y3Wly0rbKraa1YDtqEvCMjTAp7Eo30xCCwJmYQrWLzKQl7Ga21jl52GDx2j0
Z5n7ObskajwCf/UV/Le8y8c9VLrQJgNTz7dxZlMNzwjdFSkUo3EMKXuexMUV
qUqu05f/4YfWSe0B1n5xzoSCRUaB+H9a60dnIr2HXKPFmBh2+zNo6WtqX6rE
PNN5BgfEagP1zMKln0rR2xrJC55DfDwoxKXg4DaGb12zJFHIOvEuV+zEZBjP
0ZcvBsWTATE1Jaup49P0no5ZvpHIoD6GhrbW7ZorrlJecG1wlfDznJ/wDIgK
RzZa1n0jyG2CxHI/NEp+dvjmQTi7g/IGcQfIMnHC2TmzblTZ83OxV9ZjJsT4
TKxpOAcyycKep1h/RqBOimWbHhBfON05rx46GfxeHEqUvxmDUYGKRpH/jbFn
WvZLuYr1BWzwbSkxXBiymSe5l2nQqbm7PvYz1esdGnl0RhHInBsJmgarFZmR
MbM0MD3cYsSvbhubq52FNIeocJMDeVoOhB/SY8Z9mvui+4OnOy2n2WP0/Zky
uOQVNmYqE71E6e10SllqxQ2pNRoUREWJBgyC2As92iU0Irlv/KwyP8yKjk9z
VCZWaetvZnwQxbh1s8pSOr8r6g4NS6N7e6AyHz+Fy1/dW9YHfyoGFTBsJ7Za
tXF9OOFSaJlOyE2yCZxWfuHio/JSxFBBlJ4opUE9O1QL22hCWykhyY64/PKI
3aWlL0K2O8hDJ0nynNElYYHfSJhKmcRd59Glav6AXybAfVzClwYqWhTwouQk
n/aMBGqhJAcj0MEEs5M9ZNYHvXR9jEjmASQuTBP9f8RyTeMGci44IvY9Svfh
m0yHSu/h1yduGdJGgkNTbCYyWIBN86sKwceHFDTdMr2QImjAfZDiWeqQWagE
ktY0J78Zu5sr2guS+9GD6hcAhpvVcW03TEtpVLasR4XyJ1VemVUOfE3mQFt+
ONJdRjc0nKc3a+YPxaXNBJ8YnNOLITM14mOqB169mXcPZX0aApMfI1u8pKB1
a97I9xddgStOE//Iuu57Ub9+c7OvReaAL+kkf0Njia9GFevwrkuvMKHbaXZg
D215mvdqHMqS4636iIEM1Zs1MeFv5jcEPx+rn8hk/NX/tZxdwvpmkRjGimtP
lKdzzarUX+1YTiPAzb1ubOzrJwNv7NEfHd+gSBTF/s3W6s4G4lA+L5xCM7bc
eGTM5BQzmLCJUxYoj60Vf3nOuZDVqbeRNLpmtNCyWbIYLSezhz1d9RQZoN2k
pzfH+CEUrzb3PcewAd4wtAk6AyibzEGVeGR/M9cYvPgXvUgvDOVi7y9CnWr9
NCG9dYUXfMj1oWMuKqcOnfsketEyb4y/haBcE2D9teWwAvUjzKtIdmOKC0oE
LGSpU8p1xc0snF6IG9eLk2uLKbwfEFxRJBUQC1VS9u5uXVhanOLJrwK0jkF0
rx/DhazWSBe0H8Zf0M/+D5gNSTYOBTxKLswD9F8wXX908M4Fn8UqWFF+AYOJ
hjfEeEPYHaXf3ETVXdm/9oy0DaTUCKWKtuNkv0OoODXRqOYVXruSJ3uRI2uZ
tQLcw1Agz3E9u1yjwLQ2k7QURkv/EeARqo7ByqI7KWdBczGVds6Sx1Vo3yZf
BG4vQ5qLnXDbLAN0lLzRoOPQj/mewz6Ob7JVoPAE6jZJeA0q/Rv3PUuQiR42
5UfkmLMFHODpXhN8i05XVgfORe/jsIlCpwGdtv9zjDF9E1VOXOIxVkaW8H4Q
H02TxxlQcpH5qUzrqv3UaQ2vNsRE+wRAd5id89my5NzrYjG/SxrhpPZ/xbq0
gWJKeYpRmYLS0LPNSHhm24ORXijEBn2J7V7aijok77WnIRtFtRvd4i0Ay90x
BuIAGcs/1auN//CQWRrd1ajeDnAW958uRnlJDzjjPe0rgzAKJEZ9oHtJjeDa
4flTudIHdotbxtujYGE7IxsJLTdybliZZUcEGjDIjWQgnltquqGsCPsciI/p
/JyIYEjYG+MJIcIyy+M11yKapk4+ByL+ltEsWPGUNJecFAZXm+NotKwSivXG
0SLdcPrtaYCUMdRPllCqbghbIx8vAez7TO78CdZEov9BXZ8OoXFgPMyL4XYK
B4dlDaIrli2RDkNmYKEtaTrOTCro8T5kX+O5HXTHDJOyk2IVql+xkkiMEuGI
1vFpS2vJkooazvHMiM5p7d3P5q+zdb6E79rGU/+fei1ue1hAXLcZkzpeIo2k
E92+66W+Ms9muw7u7roax6zJj+/aaJtFKEj9JyJ9KpCwmQX2K7dj7VA5e/Pa
OKpzfQPYy3hGpty9NXuufppKUXkAzIWe/EMNPoV12mmyRdAFUanYHjwNJD23
RzsVTY9lnhc/QlH97EBli0x4CsoOIR8SBjNk8r85ww6ITCgtQHgseUf0a6UO
asfbgT/odGYYvc15rRoRs/W3qfL2DktIz29u7SkPDm1259fEq/Wt1EzjHSUe
om3Lm+qnNqYjvYAFeu9hG/ylCFINYwKCYl3shc4e55Fdi4kj0dQCAY4zRhLl
WCqUwnB4uZEpJ/b/xAljRXNo4pNHhfjbglc5OE5TRJ1lJbABWsFhiBAk0tEe
64tg5R3hb1IZqlmgB6EGyLWs2GsvENHlRsJyp7+212Kifvkzp+MU8uwLWNZ7
T5eHEziedjzOff0lpzuAScQX0sYOWIWre8IlGlTbll2tTmCj8ccLgVvqOGXE
J7RHawPfyK6H/55gJU9jfHIuWbJnBHk9/MMsBCaJueNGfi2ppv4uEBAC+JWN
NOL3XniAJA265jkqRaSC/3gdGTy1j5DMDl7KtuhrzUN0uyyK0p+/7HoLKzHj
BoTCR1RTSN4apIQ7ULp3ddYuPVMGdjWU6TyR+nje5OJxSoPA5dmrqV7OOuCU
/ijdvEwSkNxJdHupHuTP2XAMV3M6hCodFF/rj91dFMYb2xSJ3dsVl47+m/01
J25QYTNmxqCiddLhNEpmeW49q4FhhxvAaGIaWsUvT5WWqe0adUaAo97xSkuw
ZYH7AhFvpVce0mL2qT3S9i1m8Nxqvn5mUeXZQXW2nfeEHKQBOPWSozjobtK2
MpgOozvgh1aEuYesEe9+3WDo4aAnIoCn2MVWI8ZFDHtHsS7WOuQNLTG5KRUO
X21TMmX80su4vqzp+td8ilFnDjxO6QSh75YlG6202hnS+xcNe3HYmAN5MGxZ
ygSbr/uzeXfKAS6Q7hKNsrh0jEkuIOdUfycXgD74vQO+p25rQlR9rAJ8KDcc
QkP/AL6HJs3Xi2r1azB3wjLPpEjHorTmiPXZ0nO8d0CkTsBNRkP9oXRpo5cB
PVOmgnzIMiw84RBmCCb7kYCt73Nb/xpqXbZ3/dsjg1D7dDJUvvm3Yjsn0U6N
MA0iOPgIUliNgWtzOcZ58nCXC57WDrg9xNewdqHLVlHsh9ay7zaswrYe6QRz
TZNIhnmIatytcBKj5G7ijy7c6g6skK0bR32pk2TzJ4jbdbMc/YiGzN7k56SK
MTrm4mTdFPoEjdYXHbmt/Eu4xiuf0ES8tOsqmU2X3wxFbSPwMk5euG5w7Sgq
YkFYc1EGeOrLpBlPy7TfFznodhaNMdDS5z6Gm9hXXTTnCeUyXY/Ini5RMBZA
QUViTf1mP9Bb3oJyldNVqGcPGuXBa/n10T4A0v4cajo/B8V8XDIN+YsUrnP2
qW5fo+LmIaBSD1DnhZa/ubf63mZNK6auxHavPwY9HBm/DcnIp6DYE3CDKNM/
ZxQoOIMnK8dVlHiVh7TQSaag0Zv9Paagz6S/JYkj0It9wywNqcxFYZCXfwOl
QrTv6VLzqXS0ifH7K8Yx6395wnMwrTFNRF6eBeryWoz/rRNHHuL5EbtG541S
8/CUBM37fEEOFMKjOIa95JVw8KVUNGLKpINZFN7R9vcFmkxq6SFHOzf8TruJ
QNwaDNu9Dn2oOaS2Ur1lInHeyJqktO8Oog1TdVKAgIFduKDc/1JQBz4wSsmo
yoWtKasoOKksJu1NJ2Abc0wLoLRoElNjCsBwzVee74VGzV/qCbXIo07A13wP
TL9WR7Xub8JDtUWVIjZyf8ISMwoeUaIfB5HwySTRbT/Asdl9Q5hNqcAsguEI
ysi8ZpnhT+p4eoPWSi/7WFVaNZaLtAzbfEEYcEAKhRd1NroWWxuak7Qx5sCe
XKOrEvmYvN5mLNsTT+9MMC8NI7MXRtFPHgfwdZf6ZKlMh0XLqypL5qpvRuId
wPO7i5i5aUEdJ8BVxLpy6BakxdkuXkYDnSllzS6CeKk2jQKUK6hboT1Xxy8K
THF1vp9hxJVEC/fpzLTrQ0cW6Q9d15BUv93ipYYnAqqPxLyBrGDUb7uRXBJ9
KPpGomvlsaBCHoD3SkKcbMTnqBF+qTnsnZ2tX5Z9fAzrlKfmOhOYf5IPHkFt
mKzAb1ltV/m9wsp+wb/vCxhdcgSiNBM66nrNcZXPYKYyytxju5O9oVi26sXQ
1564YjvbTLwMbGooK4JTXRehXYr3eMr4Xwc9P62BUXYQBellRczgn1GrYcFa
XnSq7VwNw1L9pWV2dCanpIc1Cz/KdsbyIAbVyJMq+bVan74UUY5N1OGRql7O
5ZQO35vlPKkMeyiQYUEHBtxJ9kBAB6YHIe8DLIT0pJS/BmiiVKlLxic3nYAH
wysuQdYl2vP6lx/nbBrj0HoGW78ZKKJ00fAeZqZ7Zp0NQOa2RDWS2LV3gNU2
o5P+KNK24qS4ZeOd4FqBCKPaKxouBOBGqPKWEgrVWvDayHuzFqV2RklJotV/
6s9+2V62PWYpCUF34XDs9PxMKbKyQPY1QOioZrUurFIYgFlC57w9LwXJ41a1
lfBJXb5Mz5jlaO9+RRB5ItlQIHcy6CbYCB7UQQvurUAjKT2ERr3ib5PUPv1j
eFsJnz2OBcqaQl8OCkxzaYfSBG9s6Sr+9yWubAEVglaNScuKCdnb5dTUd0v+
pm0b/Xyo5ULnoibJeyfYY6mGUQHIWF3pUT+2qzOPZX5Uu56axTM29gw1GjiK
LGqpcj0p3fPhmts51RE+XiwzIlQno20MtObjwFKxIi1SFpxmU5gWafg5P3Zx
N7zaGdvn/9EXJrALTmVdGWEa1BoCU8GR5+NDaLDsbr1ALyxT1N2nSx1V5ylW
WV3UNGyTmWwC8aGdf3juOcjXzdkDwSHefvi9euNMf3f14PCuiOXFQozdUmbs
VrvNENz+N4AeYvqXb4j5Mb4ug0oDGaIBhC9myYn58FmLQVJ6yvsiRdARo3kb
C0DIpCbpNG6tUQIPj+FK8Hw0c32zFveMegCwQF5E6vDy8IbIiWTh2e0sD7hZ
E/38QC2TLQei27j9ZJuOF1BFtRBQ0LCzRnQCx+JpZy3HmSnutuINp6Euu/nU
80V8RJwmOx5FcwItylcQ+IP/fAGbNiKf7UxPTc0a9InujcB9Aa+1Uth4P1Zs
K4AsqlpQWYlqV+W+cpOLnLef0oRGBGTtoF4Re5tjHUCL5g+Age4Ochr6jaGD
BaMvLJF4tvBw+UQYxoT1t2Axl3uc0DZ0YUum+ex5JsTA35h3iEMsFl5iXGrk
y7Nt8SzMFj+XZUUR7dhVsurRkJb3Ynw3hW3O++r2ctZAY2Ae+RYenL+igxGp
HavRHeZ8hFLn5ea1DUy1NH3ZLpD5q26HkzlAaOi7yfCYcWZGIJXbhShtzfNC
lsHAFajcuUnlbt2JLg8EEM322W+5qqAqbO0nVMuaAaqiM3KvJWJruSuMZnY1
1ypcK5tPWEKhgRrUXSitUfyuRtOIFNSP+j6H/CQEWmHHq/2+pHSigc/kzXNC
QPdZD3FnNmaVVMGEEGEITB1yeOvIbDZyRcYv6po6QJyisgR6hohjErSSZ2pr
FNrlypUS/ZharMSI3bgayGFOrRslWeLEVhbbFHQrjz+3f6ut8wm9VgGVrFlH
ZwoHXonD5fmW07SnlpUrw9hv7m34IywBVM2SsO+92KvBb57XRdkxHjlwkU43
WniUaxiN/cjW9rlD4eFqYvl7e7TNocYFLoo1oZciqJPNhhYdUVaVHfMaZC0a
KZtLSgo6Nj4s0ItwRkqTgiKb2coocSnJQNoI9SMb3QpuUeO4rnZvOU4MY1eG
3g3wESY/XzHNIj4H19qDscl0/E8KlUl+QRDHxT2jgF6qooOYvuN6qIAN3yDP
JXVFdW/0IbZWQptqdkSFHUE3zVTC1qG8XJx+Z5hn+jbdvQUUHv1tUyi9GZtg
rSF4Ms4RJ0I1Z7tvUdX5BbbVj9wYjAotd1aBTjfdvnw8qnIGJ/7Nilf7+Tsx
J7WPEOcUV5JOU2Rb1N46Wzt/1jm1vVREUR/DeVj7H27fVMs/4/c/TC29bGLx
ZuvbzcQx6PQa/lR4EvG5A85+bggdilkCgecHDCZTzL1W44CzsLCfVxLzSgAT
ZsWiMg+LS9hcmFie08EugSMkjP+C9YNqeEYEjhfpqqnzOBeA2D8M2N95weKc
KCDcqFm6eAA/aPC7o4SEKQC7YR7Jf2NK7ni0BZ+QZk0djizYz/Y2uv0+gGkR
Mi5DK/0L95P3w3EWBIsHEs/xlf01SIkeIaYvrUb4+XisC2qvShufYotlQC57
GjGK0Aqnelm3kWKAXHInbRFy66yxNf4naHv6E6ug4Tp3GRyqeeB8QC+bu3cH
Kr9pzgEb8XC4Ppkg4A1+GOqwa17kn2m/oJetFTaPY/M+cNqlmTd/juoroXK6
5Ozg5iIR+2ZjdNqyFV3vMU3r3kbLFmx2qg8D7qIogqGEyLo9FafIqA6JhxpN
U8CYdNT02gRDrTeJLWsA1bEYKEfosDodnhmhV+gDH5QjKpsLjflWgXofAntS
YdhlS2WJT9IsfV/VhxCxVeYbzt5CwM5JFRBcLeiknW6F0U9KEJsBnkxJz8Wq
5H95gOUVuRYj3Nz4wryVB2z2vKdvDoF5nXiFP/WHhDUx7GYRDRurVTl6Ji7u
gBg6d0avEDuzgzgrT6zjQW110PMs7efJGdoeAoeSGZPKFPVYR3m8Pyk4+L1K
E1mrW/y+zpiylPDyT7tuA05JxwAd171OKPdddm60peBuK2XDsnHOnYIN4hHY
851ZagYVnkOzZLZGrZxAG3AmkvDda9goNLXomIW9LfAvX9BKuLz1PhrHga8z
RGYXBoy+sTjI4SYbhCB6oHR1cUkXEWI9t3FTvAZOtF+08E3JBVvJNHUvQKSg
7dY5JkY7tqXrP0vdDF81JenT/FvmtlWjG6QPQ79nMavALRiBUJaidN/c5iMC
rpze3FZppi9tr+lJakUTyOUx/78FJ1J4i8kR3vn+yaJBIKwi2ZepvqijD2N2
tP7t8EmrDlykhsZbPVlDUfnBgqIs0f9FstRq4v1GBvWQj0mJkNYZazPci9wI
M4dhWuHmDWmIoVbkWsMpPXb6JYvEiYTrGa5SbWNZWZHgGDT0NaFRHeBioKjb
s8uPSc8dS9jpSaoQHJnNobUn3ha5oWkUobf0cGRFgwrjpm7XmMfbHfHFw3nQ
k3kfDQfFnOPwSJxwJPGRUEKKukP0fVKK0pAF3MtWNYDFxtSyxEJaQ6QYf5xz
R62l2dGUAxQiWJOqUBNQwL9bFIAkISI2XEn1t92/qiBJ0qneCdT77sdxgPsN
xghOKU9KeMojQW0HAbgJK2np+dfYiCCKgnUlcMJwuZZUOtNUefg0zBtG71Dy
Acjo9/hFIhBacn908GyA82/jJu5/tdfwmazAKja8eZ4axSWMk8Qbjwm7Nw83
5BmwCzuyQentH0kEog7WCL1ZL9HlbTWa1en2hK8QR2pUyW5Fo/cSn7UKyn3G
GXwHQwg1pJwIZAXFDNnau3BPF+tf1ccm0m3MjebWJj8bGTzVnYU8Y7g1ryat
6hanFVCICW1xrharTCFptqA/cUVaUK/nkan+h1Z1ZqSpVk6XQSTQXn2CRIp/
xI1SnLLvgIQEi+MQXXafAXvcwVI1teMy/prB70Ylkij/EsfplEeN6O6DlfN7
IcXHpmy98TVYlnL0s9NQSsh4aD4NYlejhsjS/4Uc3Y2IngQ2amsbdCliEhpw
6WaYr5F5y6BZ0ddwC2AF275RvUJ6EPzaExy49fRBA8GuefnasvD6ttVYKpgQ
3OZH+Pu/3mwGNfXyhXGJ4aSUPC9RTikJpTfYilIhzRRxgHM2O/cO3sqPPGSt
AyuTOs7w3Fd54dy9ESKlt84c/RTtSlNUFw6Sf+8aFL46gGsHfzkD2oQkxnVr
uOkJLhQVk3ZY6nqza6Su6CHX70lCCdaX4C17OarjcrRbDIE2blzx1t9Sx8u0
ZRy4RXWE2INxL0HRmsC7PZ0ymHztyqVkdM7NOc4fWi/nVCzvknsWuc7WsNXt
18esdRNckRUYbZPv/ORcSUIcvP+/LoCkpX1D6vCj3PMD1LnqnlFC5h8kCq0+
tGpAIgb4oxsz8yz3QmCWglJXkMKq6xxWh1MR3dDS8Lkmf+cee1riVDwluSxy
0yz5DS9hCTv+jYyT8mubPMboeHGkKbqNVvkuRGq69i7ipwi54HNA2KhdYDx3
bWuQjwoJQLIP0rKoA3bDoaM2rB7LaKsmil1aEuXqJvSZpl+qneTrgOebDFrE
YY7CY+a+H+/TQkO+rWP0hDyMudKqmTf5W8wXenyF5TMTh0TvqenccN+iHh0E
irgWqnBmeKxP/zZDY3L7jsC/Q5oV7i+xzcmDGockcuI+HF0vn2zV3ZqKp0Z9
9zxTlC5sdzMgNtQOO+DH1uL1H87vm/vSMjr0Ez9bVq9itQsswhc6Cx0a61M9
DBviGofnNA39hnsPLMHtt/N4fjctAEDCeyG4DF0cLLxpLkXh94ChjxZPx100
9IC+gjI2Oxdk/1kD8wBDDQWuaGqufZlC6DRxLRKh9huLpsR8dkLBr+jvXjoX
RO/pUP/OTBiMB7L7tkdbnwWUUSQhU4SU0wg3oihF7vzoTxzt8I36TdQSyLEh
/nN+ls11fik/ghe0OHFWfqjbUhN+wwOX0/QnWNJ9m0+EewQIxeYK3g+F8uIB
ipridSP0eAubz5y6+l8/V21RSDpq6Dhfhk1CV/z9V7P4ROGm67a0p0cg4K9r
13sU7hROD1t7+NMkSA9xwWyBoN8MW4RtCDPVnVZOz7xIG4mUdsjfci/q3gGh
Aw1gTeutMIDngEbmPbbnYV9Wwu4edKSg4s0JgaY1QA0o2iwcd/QKRZkb6upi
3cJ3opyySRQJ1xxPAvgug/XMEH3hI8/yaY/rAHeg/QB877nRnFN57lkXHxD6
1oNJ9+aQgsMos+HZIaqLZgmBnyYTXEPJQMyw5/rfmge2bIfWfPWDDw0YNn0I
0pXaiboK28OKWdNwt40Nog0X6c4/7ViUvByXaXMUigFCKanfho3iXNh51l0k
3FMPmb11NINdKqiIZb6yRDEGv7GNZq91ZnltyYBwkkWjY7G8ByZGfKWUTBXh
ZAKZMS+NkcnwRcnOnoN5rP4A57VCSsP73jdFOLr89/aaYlWckw3IQ3WHCj93
ST0NdN6VhUAuf2wUo9BZgOhpYDfLHXiy7lqzBl/Ktc49UYJCbkhQARktJIbW
e5CEfQXQ81Ddtvt6MJXdRPli5BfE6GrZcxK8QHgH3OAmjy8urWHafvfg2Sc7
W3Zy+X4ZnL6kJWicQvrWeR73OWw8kyTZTVJmCjNt7YxIMGes+iGf6esmzCQe
UMHsyAlfr7iBp8gSf+mhGoj8iG/j3/VReLIvxcMeyRAepTfdbEyTr2qTxZYa
Nv3vrI3Dq048LK/On28bI0x98eneP91ri5ql+eVWo/03XUmEqeJyOEu+pSWi
9tHHZN/j36eu5fnGgBLBgJuRcLGu0BDGVXY+yfnzHof77tmJ474TcjdPVO17
ixbYmYDHGS9JtX5ITjasPRHQKrIY9L/AVKNIGRYdQ5DrG8Nc/iCIf06Lk1qi
vKjeBtkIOxqdwr9QZgh5CP9BAhrK2Z2h7NyxfXiI9ZX3Q4WJWgqnISphk1ME
tAJqQO3ZJInXmdghi+MndIsstBZYkubcS7hoHZet0rpVbAV0fqnbkr3Ki016
Zk3itnluS3+3CbiInw2LWoFUMzMDQ/Eru5qIol8Y/BdRKa32KJCtFwBtuIHy
LLUbsTsgNj5l69wajx1wvZBgqVPyVqQAm+spQViKChmO1SyNdPew5OoScmkO
k13pUjSxo5a/L1rPMTZyzAL+cNLOJKboDoJvEADiK1jP/lEcMasrvCdcvZQz
Sm/IBx3QGKlm8g+EVvATOXRPjEebcDQ2f6znn6VT4naPwyROfI0dWXNWs9UT
4Q/yzvIbNDEnTHCS8b1gwRfupjjTUeiW7taqGMHZCRknEfAwlP2UG8/ZlKSz
iZ6SJmujenVjuWgInhg/fns+jntZPT5R/XJ5J2XBXv4C5IZkXWCxN8RFmTqp
K+TYeaUzRt9chK7K3pUExrpQQSPsAoLLiYKsmKcTNK7LtHfegsMuJhGYRNIv
7l1ZiAz0ceOuXGqLG/ISx05PacSW6CHYTLms5nJ5rK5FHqD7S+GTzw23io9k
ACaUbTT2ouCz/+P2fBscHaMe9urguXGBvHTGgmSixBFkCWLXCjtTnltf+SBy
mWIIYVlj8WFQZEenxqZg6s4GTp0KSd2oFg1yp2lR1SVX5aWPspNXOFJXpqIx
NKhdzAvNbmZvnif+F6PPXlq04HKBA1iXgBPdCNLncOQnXphUNjWfcyoOXElR
BCKfUqeuBzaMBTLJakyRUzWATnztuKecwtOyNLlzDxDrzDZUbh1hUz7CyYs/
a38Hdv8j0oKcxqylvDIfHP0FAUPBg59aFnl68BEQeJb5Ph7lrzgSt47an8l5
HjN6klowD8w1MdKNKmlkA2XoLU9MRB9kmJHassRQ0sHJ4pUPS3C0vSQGtoGT
dkhu8kpRJMtglDitauCwAyZYBhtqQhZwZDF1s7rAf6nnoAcnNzl1GPibPnWf
v1C90WAajarXlPuCxjVwpjpUILUfd1rY1bufbpux2v4Pl25qVQJ5PD2ZQiT7
q2266Ptm/dwpq8lLomVel6aB8f7yoTgZRxi4VzyNN9P2GFUZe/Us+Kpgc7Yh
MadKnvrXEWs8ZqGiUarO7Ab2669lG6Kf2/XTtUfFYohe5qkWA5Y2PY45dU/0
txnviR5J0HUxIFUpPBp49eBHP1nTNSAULxQ7KUfcPn1ulrp/J/hv3l8MTkAX
Pl/IB0MpJE4YdGhTKtjpja3y9XMrm1faHtVf31iBABiOAJWgq0ZbKpZytBX3
B9gfAHV3eRcgkhUBkjv85o7geE7Buypzp6skzVHVD+bQ9XMkq8z/jbtZ8WoI
Et8Sk/UKJ77EbbA0m2hw2dTFgS5KPcZo/+XVoFeTn/AyEOiLXndBpvFsw8Xa
ldmO4aRFrAIWX7+JJUFpfJaNds4IMk0oj/MXxpR5Md1yt0aw93iVp6O/8J0f
/0bv5szUSpAoKvFd2dKvWN71W9lRID+jpLJ/znmbhh68dHWBUCY9ZywSDO0a
eAZpZ+m5VOEcYvhZxjhZP6zoPNUfXlFtolcVCK+ecxClUMY/fzSmKnTlUESQ
z4UrbAcydFFI7eiTYvvVwh4Erz2xhbJcMP60c1JIjbPjvvArEFjL9T75Sx7n
VPqU7MD6P5w3QytaXzt743C32oOvMrQpwrKX6HzJiSk/fpvTXuYg8RVXE8Pj
KaS7F3TeBNqFQHA0DcPgcBicqw6gaxMi9PDdewxilXJG4VrhYYldbT3v+9mi
SAoGc341HD5SSGoe1Y/Mh4mrSs1gsG0tpxxWAmK3h7S2G7uI+DoN2cDVSyGR
JbOXdQnLRREk2KdLF/8nrqYuwz6hQiYKqVviIdvxF8i/fTPgw9p9LH8B6czA
N+9mx4zQ3i2zTm1VJeSU7E+nFvgWMjoFs/GxHcQEjX7UUMrcSya9A5TKKN0+
aeP68UpXvwAe52rDSxrIlIIS9dqVnEaT0EGn4vtvDDYoqMtJ08wWvdhFERTD
LmlNH+I63Vs2AxGz+lBhrFWnrqBMuhHbds72mIUcTKCjU61/1FHd8tCkl1N3
JXfnsmbIu0uGRURmG76wVgtucyMQy8jRiDrTIyzSSQrBJyIpbJ1v3OuC66xW
4fkjXMYToBnLR6lkZsZYUm88koNXJjIx964Vxl+DFgTLJGtYONevZMEYwJVb
T9EYobKDA94/GHlartX907JMFruaV98xANraO2R31TC6H4UZdL0rLmKBR2iI
kBgm1TXjw7RIZGOTi4hxlBGv4hFqpzyMHQxxQysVrZ4rsdOFUgEVbI3Fpw0B
AMfi8b1UK3zm6+9OMPmLLUWoqPoU2FXsxADThiJYl76qx0DUisgUBBCqaYlV
y1KfphKqlyh2MvawnE3Xe0i7i2i3DKGf2e4YhLD6VJcwRThUyCgXSl2tT499
4pCpgTWp/luQjSBU9IRpXydTYUNNNeNjuG4s7J1GpZ/GslCJa7W2Z9wZxvsF
XmEUPOdx2FS+SCj45BYzGvD0PAltNvIKqDCzxPd0OCMSwzOlpx3Jo6pc0qjB
vQVlwM1qCOohVmvavew4zQQvk2qjAaYU+/aBJ3WrBJ2IlTQAKbrttG1ae7Ig
OOFcEpJRWdxIRiJdJOrAAez8ryJ9tVpUp1/QIcJHhOmyYFXE+rR7zXj+tyYZ
alA0kbba89ognBLkH6hUhyFlWzJV4TQyFKSR9jHPdvmWdX+JNUdPS8ZLOj6g
ScH+1m2ACf7qguNmeHvsBV5xRlRhehWUIxrTa33mR02/mzVr4AJuQNYds5iT
/3zG8qco8m5LxmdOsJv9rzCWZWkazoFY43x7MhSA71fOhkS8tjQx3eF6Nhfb
6hJ23EKIBmmP4aLjCpdPiCNg/cKCXZegQz99DlZZEmy0+AinImFgY24qzOU0
GCsLFSaQWksti39QEj43+GZOVDsdGzGtyy9PZ8aXLoCrFaPSWv9aBTNEXSD2
mrgB+0TuCHxRh+5YBM5u4P54OYNzZaxnq1GQ4gfkPLFbZ/R5mtd5mSoROATK
tbfcqyUcwIV2LIngyzAPx9NePIw6dHSUtSev3scF8xk5aoI+/AvutGlhGCqI
ag5kXkD1tlZuJynJTHy0W3dvGTCpJRt/qL9i4y6ai0hVKjGuGC3M2rvp1y7V
Kc3S0rj6kVBiDNRfSfstr9P3+RPPXIGfm1GQgc4xHJ2RyXCr3H+fYe8tHuEQ
w2nfs1hPuMq3y32RSgMOSjWFi0YNWy9hPwXalM/PFXMKcts2Ai0GT257PG5l
tGmODonAOUh684h8JRRtCIzYXk1o5K+fBwpIFUK8is1yV8NLhVe6+B8+fZWe
9ylRxiDukb7D+JA1dcQpBTII+SjAMR1NLP6TNqAOISWg2ZNKo7Tw/wVmFvdD
eYAh1BtOPgeNf+rEsM9ilZ+oNvfftgJ5Vc0dE7eK1XGIUW+V3tirZN7Qqeov
2wCf7eLNLsQTCKlMWcBvhZzeSSYVrr/1Es6Lf2Nc4GYPgGQUbbnOCaSOE9bv
zl6v4wXDYuNsfGozS8ed9W2kULPEuIDRWqoJSdyH+tQrW1X06MJaw6HhuV3H
VOLkNEbkyJb23/Yn0SrCm0kNohBxb5/XRWKW2DymmaUBPoBvZg+J6PtXxTkw
I7eN1IP9RJ8YVxvYzZ66zX7JG6bErgJACk1hzihA64BHHKEdNW/8QDikkjy9
MQWFbd1UIvp4eFtOD8o5FMpzLPFyqblCg+xf1RP6KuTqew9ttDjHxPmYykqe
rF87+GICgQBDnOfl4wr7iXU4icgEZuxZbz9PJcUERdvBreLPTli1CenVUVkF
mey5/DDE8H3YN7W5W6w0wNFpfldI+YPGBoFmzvRrMezhGPZJMQbt3HsBxG3N
u7YLshGPLGyPZJeuyp5JV1PA+NTm9npBNyTsz+NcDwIwRSawjppgozbOXmlI
pU4H80U/gavsrAKLVvSZmJVkYlk13jO5N8ZGUcWTqr49DXJdXi4MCc9ziPVH
tJlDxqHtxc+w/9y5HqmMJPLYeCdUcAL+f9U/uJVRibKxmkd7qOz62OOQ24Ho
P6nPRbEJqHYaXDJW29MvOlBIGBKy0TRjbKkkWZqlnKnXmGnkGFCjElocFh7D
S21J0GD5EV0gGJm6vp6QOflV9Iac2GJXwN94CNhl/+68pIopiYsALxLft3pn
nQrM2N8DKptnC+HElcpwOpkLH/VlDaTlCg6IXr/Uf1WGRYuamOHDaifuunk3
400MV47ugIbHASDd00UOdpzC0pJcTWlPvNO+Af1uK8crKl49QKNyABuWEUmL
UW4a8IPccAfHb5z+txe18WO9V+9MrXwUNHcWrVFQ8MLRmYADyVDv/Co4kp4F
cJpJ+Aa4EMG1DgSPvffx1599DrwGzh8W360XUjtrTDO9Z1BOb0brXcqkgCDy
U1nyAVldvarzbiV2slP1RQjSRsv44O+S9ELYYZ+pwIwyq5Guuq4kkh8A1UIq
r14CdlXc+pMeYpxmQXmXCSqlvVjCbjE2jhYuqRLcCpTwSaiZ4dpMOO6q9s66
NQmZhw5xqIJOi4MMiMSe0gyrLScZLWJu77MDBbsKyEZBPqjxsWyv13bt5mJs
3UOggT49S1M15YEfUBJdhJNTU1+AppGCDHjO7SgSSMamHZYxOORKp6OIzcge
3A0lxMmLTbW/e/J7KJeS7SIerCoVy0FKtGea1utNjsXbb2e3RYPq5/4MlzOw
iOwMhu2tE69gEVHtZjFNPkdImsVJ3SIo28Na+qyxeAWZ7igRyJiJyPnbMHEc
sxbnPLE3QPC7prXnSQh4Re6cWiY/J2az3u+v0/oj7aXm1yB/8niyDP9iEc1a
HGGBz/Wa1o39+H/7RTMp/05+hWnT/a8yK0Q7SZ91Jo2gpN9NREH+dbpnNCEW
SVyEBcTeDkW+X7ISx/mvEzjusnaAlH+eX6YtFVQ0kDGV1svwtOf5Mbh40AFW
bWrYn+EMdgA7chL/vw/sfRH/EDuw/57JXFX7yWSeYxAPOGUeFtizKJGgOEy7
F3cp0ZpP5UllJwe6W4enG/n6LdQ3Fjlhc0dg1oyRKJiuaAQCE/npYSAzB5FH
19gNIegX8roMZ8KfLStGiAhnfkm9AzI9QuGizPuYgqUpBR3Deig9/mP17heV
jXYmcE0u0NJOCutJkmolUxasqnY8fyhQ2yBe83QSr/EkY4KJtSriGQbLELhL
MP31ZlShILl6/fxR6ite4kdl5f7uGJjJsDtNPKLQnnUGW0P7F6YIQZTNKj5e
xBENEznOKsDTfLFOenMldLX30Ic0/geSmAIvCMFLDZLvdqhXNkdSYu0XWB4W
ik9oKzFQ3uEvqYtAJTb8o4+U28I3CyRyUDHc1rYd25Yie4PnDWOu2Z1OmGKL
ekYl+9vMJoPdI0tRdFBQh4kz3qusRO3AzVXVyualKucN4buXQTEW4VB9fNE1
3T1OK/YyHwgknTvNa7afhpPvnD6VI/8PFUmDEWLdHzVF2YJxx4HTXW+zRPru
+LZLt5NV+zu8lWF5j1jGav0mdgfQeU4aF6sJJzawLSimZwvBYtcr+KsdkK86
uV+1oDVJMuDfyiblS9uNbz4Z3bHS/I8o81iypzJURty0hQRDryt77Ytj54ex
8EdJ1hKUd2l+stH0Vjrrlu+kCTojs0dsWlaEGrD7DAT+EPOgDWu8T1opGHCE
zDlfPFjds+fZkmEFY1OvbX8uQL2rOcFQ3BFXXkYc84NjpPtNmhK2jt6kVtn3
J8fbtNr6YnT6MgvQHtdl6jRAYrLMXDAX90H7yDoc4u2XJWwsDsIKDjH/32xP
LEG+C+mBP/hhOoq+J3gOZQiZ/2WcQ3k2RS8ih674r/rc9ShSYJuOvIIHUSQj
R3p2tH3NzVOxJdKFq6mmjFovlRsAVAUYNpssuiMoxnpB1xlo6PKUCgfXj7Mi
QHPeM1XtDofKf7LC30ScZ7cyJUdI2gFX06cUY7tz7apBiAKEzemLUg8bmtkf
zbujTCAlYAZ+N67aSPrUzS+zeGOrhcimF10oKV3IDYn1mZmI4VElJ8TNWlTv
+djDb5F/bRXSd2oiNe9/8sipKW/bZNJk+0uTz7vSQxrGE2Gm9uuKkXFPAy9j
SPfIQQNEkbs2RwObmDI9kBAqqOPLevKhXwNfNaDJ1rxftHeYn3xV+GdAFb9F
c+CpoikRhAePvVp98cU0CCAjOMZFRLQzO+phmRyap1MtWkkFQeYEvz2wWIrA
C4Z9klbx4jlcQWxPPkBtFOsrZ+nh7cUEK0zan8Sm5akMN1HzZGf2si9vK4Dy
LXrya1YaBfdWun4eE4X22J15oBXjPQqM/YQ4Zr2ygTRXJc3e2u+R6hZHV00W
kY9WexmSAYyJG5RadHqC9qL+OQsrIU3X0Gfe+XVcTr3D/3y3PkuXeI2SAQ2l
QdU565TkAF/53Mteq1Pl5XVCpadOs9QFTtMW9aPm22/+lLKYISXZlf0ryKcz
6mtn7qrY+z3074ixaD//nQ+qBSIkfLAZLbldefO050NkDjDjC9lXtjbhCCDc
S0u+bGUqEm2nHvgX04x0T2S4qGteP0vhCNmgCm5rOV0NIctapQTeTcXoAfCl
J5iiyEYNnky9PwBr4FOpi8af6XoIByY1OxEYVPs3AHG2CD/gGfg3Kgk4XlFw
aUimZn7PtY4ivVBDIcF1Smn/x+GRfBZTtYZy9L01+qmnlUQMXcV52bs/WVMx
KfMneBz3Xg0VmvNTDmyw94nwgkYAIwfVwshOS6HOf09+EuUxK2hPUqsa42ZE
KnNp/V00Oio3SqvCc0FEdJENmwfcrKPfiG3UGG++BwFdK3p7nEpVMewL+ppQ
sX7VkiFApStf/fE202remU868R8RwVHxZotJx9TjfwSl1swPqUrYW+SmP9Ks
pZuDbYaC5jAIo+qbaLxr252cRdqhnnVP2LMLhsXon369DxHq7C47CNrkk2hs
V0AHOGgBU5CasMH7ENaYdhwAJV+OCCxWasjHxKJIfqU4bDTsvQPu+BulGrYg
rBuU4PrDeHGULDBV+RF3+gcUFO9DsBeofdN7jlzIh+qPfQnoePum3vgGcSxi
a+3HcOZXGrN5gxs23mDTICtm+dc3xBI061JKNxK+1EUvZMpO/deu56XXfOpI
9hlJ3TC3Qhfmdn/ozAN7COyxA0SZnRHcj2yjnAL5ChZDlTCk0ZGPMEz0wPCz
r1RLRllTIp9IBEWcdypIMyFrKF2fLw6OkJig9XIWY5hi37ID0c+PDgKCXBvb
CXZ4bvQp9LsuPf77d0VZHNyPx/A3ey2ZvovSt8Y0I+vi+NUGjS88U9K1w57C
7W/FXNtxNIl2EHsx3xMUzbn4RvNRHsp3ZnOA1FD4xe+lB1LCSXyCsuVCcfqd
1V4T92yc4Cu1Ja4+Leuou1aXxIIZ12AwBAU+043/AemlYxkq26nrBaHFfnZ/
NFDSonnTMBFCDLFWmig3iJkuz5zO42Om7SrZ77lrirLX8K3niM5w5b1HyAaI
aMacbvZdTWb4Yi1leOwd2uxGafdj4aPUPrDk2qVRdbg29juBDgW+qzdtnKr5
p2xJvAel30mgbI++/whHZERIRDa3j5ATce51IxHMDOS7PO3C8h4hAj3XXZ4M
L5muTYs4n1kiFmuWjpCaaM92KD236s2VLJVLyAoUgW/lfBAPymRp36BYiqMv
TEIg8aFP9YYHKvfJFoeq4Aeb9rAhBhnALjIJ37rOTEn7e0BvQopycatzv3ZK
/UEGpPxoOV8QU/BmZlNKXJHBIwBEyAj59qqLLXB1jtJaH0YdbP0P7YXxChZv
HzSevwfMObKl9DjraNUoj3hDWcyi/3RTBEXYE0LEBmZumtQBlGC2zthFNZhG
7CoLhDQ+rNuzBnovMmvwN56TDxe3gxyObmwYlZ2NIw+gnjPUZZDHgi2giith
G1h7eDa/nxhlPKojx8xuEuoZ3EgwY1Gqxdd3VR6SyQrsug9iBUvEZdxAwhXm
GjcLHY7fnbMiCoUIAQItLLdbZ5jeDJDPHDqu3mJ0e65vhI1nR+KS1xcPpm6R
qFfldawxuqQGU0NS52/XPpZ8dqdDGXqchackmAyAteb0b6fXQoqVG4ub3euQ
50VzAjcL8PF6V11LOusbFKoOtjsZum243l7mxN+zkJyfnQqdQQcdi2zSO/0U
nKOdFkInoD2Fhs+A6nwSAEm9YTI8gjkexkrXCpNm6S4D2GA8tkxqcKoXYNfT
1jwuKFjC73xu7Uu5MKZ/cEAdq2shwojUB0oXHqGMtd3R5qVu2kZvZP6UpQUN
AbiqQeFk1gGgu7cTorl2iIimjQoyC6GC+1XZuYeDgWDvOXA37hx/Dxem4i65
iAQ2GtLFTakO9gT/iQRsJ5WXFLfaIqxxEF42EhgF/M/ooAw16A9cRsBjl2ox
U9+GZBcUyokZFuuknFx2ojx/XYaWckMrNn4WkZxjZoi61AKM15Rwh9dU1PP+
Mz9uX1KYdp7Kk/gan0zdugvLun5+SrsVvYiV8/cmE1lz6hrSG1dcynf9wyP+
kIScxIvh5rdrfJaToA0YejknBGuE1wv8UMpHIabnQ3sTQAxHoMh5d+Qdbq17
BZcajtNJ5gsQ5+7SwG+BnkdrNvROFDtB366TB7n2a+Oa3thHjwgU8t+zJ1dr
89LoEOZ7HfrmhCa1LcNGEsBrY0JyibtP0AVwtp+/GGXTtPCruIONgQfCIhYP
QGntJw09G7UPXhM/XYFdIuVw6iaQ/ygl7I9YN7BMQqp7ncxAACp6awnQCr0P
gBwKYliRCxR4PFNbv5UcLHSSgQAOHJgVJlWGg4kbON2xsfPS1/OSl6lw8GRN
ayA/HMU2uI18snTDkI4pGAu0+QGfKopgs3PTohRC6DnOZ8PrttI02JlVbfuf
l952tE0hvAzHxMA3E9pLLjb8T2q5z5W3NjckKYSqnnxremHfvzZCNzw5LD/Y
eXJbwxoyCHT91uV9EGm6H99/buBLzR7GWs/Z9dpgOiSXzEMsGf6toB5UjkjE
PFf0Fz7iSM0XFPtwM7WsZHdSFWVZxQvLMlAgin/DN40znJ38mHGuzGZ4GDj2
qsSuFSnHktgFlhMPKlnHwam//FO/+4demGF6djBvf3ZvHWxirin71pqtvbu5
X3AZR+e3DocV2majm0htNyxZQZTloKDUDsBddD3diKgk+OYeVy5VCOs64TKq
o2lhsYKmrULG4pbreOMO6uI4tEjTSst+v1vWwpPoXUe8bxXY/pv4kXiHVKIY
BMk3X/ORCymHRdAhs4BDmium2Xx1J6A+ZlCXXTpFkUDwfxghUzKluetiPAUy
DY7sYCDNLU6bNyHLX4jlrGQeItVJUdGkbAUyypsf1uSdTweUkNPk/9Y3gr+o
BCKuihd6TLgU6mdxPKzOurFrGMcskmNyvPKo10qfgeDl1E0nMVORQTXR5MSb
gBPVoiVetVhRNDEase6yoH7lUSwan9I9UNnWZYaBarqowt6FWabG1PH3GrD2
BxQKs7+CzmrWo3GW9p+shjP4Qt5tdWnKXIYk2IjsLm7tB+mPgOaToYYtlB5p
U9lvnfv2CWPne+g7Ogpop1nBbaJ0+1XUWegJeeU7IZEGItiPFKazEyhTQBtE
OpKsQ/ZDKlhD8aGdz26sKg7wXc7xsZgbnPPrwob8Ci9pnrLpNHN5rB8a9Uzf
fdmwiPkFA7jN0hJyswM2YAKOkYdbGaOkivWCdrEHpXqAQzOQX8674+ehwI1+
ZQ4eTlM6sf/b9EImlEq2mu+2vdpC2zhCLuowszpAwZV0GIF46W/DioTul/x8
CbHOtzGHfs6JRltuJ6qf2ZNXUEupxC9O9gQjc9xlbuHViy8b+UjOPgisWrlZ
/FX08bDcho86QF2Q0TuJmYjxrTaNCu+sp2ZzvXZWWJWXzADW0ETVT38GV3TN
TwiLJgHWEcNqMnJCwqYD3LWJ8I/Cx9qNEKA+H9w2wOk6GpIrFqMb474od7Tv
O988hp0FtVNbHVqsVYjf8P+Pl+HUuE0zr/B+fpfghJ+Jbpshq6ZbMJqpCQbx
0PTP+8tb+zcPlyZ0NrKILncOldlSMP5WZ52LRp7/k+yAIn5p6Pjo3dPrwmYR
QaEIHfD4RnfNyS6Cr8y02KO6QkHJ/uclVit5mUMq5STVsQ6ziycLoJSOlg1r
7Pu5FzA9m1cSFtDrTkx8oS1OX38yWZg8ikjnNRk0FNz1/6K3GIdPsyDnSGB7
nGVtjQxjk7BHcK4BAz/5Uq6OObtmoVynrr0a0zQiLHuHjgE/ui88mK8M/3eI
qLKB7tvRH+JhPDBcUNqr8DL8pBOVp3qxJiUk6FNJS+KCEgn5nrlG91QtPtzh
2bfXx4pFGu/BoZ3c5ZRkgCtljdWG0fO6uR8V7SJivt0w/OjN0DY/RZlfrnm9
usAy03qEgrM9iBnAcNhwqqt9P9ggjayTpwOQ2OQyYYii5CDwM+2VkmyAoiHA
ZzzxeXez+377kBV9OefhQBhYumOgq0ol1DzUpXbj6PCrhObBeiernmbUt8Nc
kIVbSGOQAFspxE6Z78h00nOGxaxO771Hh196tbYZ/nlCzmdqAmLh5a9yDnY/
PMT0Z7r2F8ZbsQwDzFdu32wD/SCmsjqiFBpnrtkvJcmST3votRsVpXwnIcnW
bZ1Qj4spbRUtOBPU58d9OUI35PEUrDH2o28bh0Rqz2wbXNIBz4MZnmlxcKw9
TInVoMA8hUM9EhlNddKvcc7JT9VR025Unt51a3XPHmO6msu4umjxcvkx04V2
B6xJOqzUK5oN4JyGH4RTzj+YWT/81ZSRdfRM12WG9r8H2tyADVTalHFgx2Xg
kjJUv5kTvzSY0275A1RutC4eBez4jHnOKyq0O2hHgqaqOz1dM9sgY2xW6X7A
3vPzKmwMQamanxL+JeLWfpyLA1YPo93trcMbc3h3jJJdGgVfrjcPppUnfB2n
Uzhjps/hHg+msvjD1GRsTjf4d1zUjk+0ZcRorI5WbZhFOUZDPgjezVPmBmsd
T4J9u1tgdjXYOLHzpvDC0qB6wN9vz3bTqvHvafkqxhI/sjfnE0xqzJ6WPAbT
ZzCmmXfyB5HLbxZmGozzOIVeaRvZlfpTMc/b5NBGGQKsgDk70kxYZxSrc5VK
aFMSztSg0cSbb+DzhcnfQk1gZU0U2c+BavO6CxxMj7oNGBYj7GKXZi50ILT1
MtLSmRS2Nh+MMYxC0BIv+Eid6HgNqe0O3MMnKlaw+xqdUA3Epja46HCnpjK0
dwb8qYIyvgbStIzODO+5y4qqtAJ0vHkCpem63c/p214QfjyJU1F30l0noUWF
vrTJRWz+mBg9lW98StMCL84MtdB5XumlL8W74ja0XDLorD+VShfsDJ9bRvrc
i3rwXEszI/qaSexaUkZ1I5UX/f56F4vA2qtrRmua4j75Vk2slvgl5qOdGar6
bypzbCktI9P8D/7PYwXyLS3jbjjQm1VMDCkjIvJTXJOcTYfQZ/WlHne+RTvJ
zYlPfGizYOnt7yMO2sYE4rDtf0pxybs0q6DApiHtKEm1NcLMyiYZg/ohXUIH
ZedMC2NKXhR1e774bf/BPIuW52yWIb2SSdva9qCvXfFVyVoP2dUYnM4iVhqw
lRsyHL/HOFBIbQyAi1MQlQcT7prFSW3lbiAd5D24NBtcjE5W2p0aTHfzI4Y2
01LvFIhc9giOVnpOYLODqaG97nI9tGPsIIHUinfkbAJ5yzeXcmWm2GAm9TyD
jXNxjcnW5wANH2s7YYSdbBVjPFjeNP1b5TzqLb/7OnQS9TNJuaczoPOd5f7g
5U3lyYOUAvq8tKhDS/XGWoojiOZM70aMddHVxMaXvise7OXDhvfFAtvTRbuh
rEwNbZxYqzN7oyYo7rhHb6NMlXjGeiq9MkSXpP5e2xyH7p5wcZXtlZQbSnL+
LuOaRsdEuZihx6h2phfRw478Q+IJGPCQD0u87Hm51KMRtqadSSJoWDS7pAut
quvZYphJI3+nJ5brXDjKOKlOHVYPWCkjrZd5nR1qGwVsXdyE6zM5ZRZB9Dku
FB0kDaVvn0a8ZbzvCTLnEAiIBGYe31B8SpLhjyhPYV8CRu24lykgGPQMHMoj
+uuSuW2J8xPtPI9ejsJbhSXfz614RFzuiiBnkHaS2s44+inx35f+XjYDaBDP
hmExFTroNJkgYZjm9t5iz9Z6Vjsi4qYxqv8h/WuIfh/xrUmU7fwsi2ogswHy
71Ba2/U9u3CHTEESqa5Z+5vxzZf6mUDOgLoSjiyQE+3Ocg9zaO5Vs3T4qWLk
Ij5Ot65p7xOerKwfgMGkLPtkqRFR2s8T79jpTNjYIx8drw92kArKRCIaGuF8
3T0iVpshs6+rYHSOk11q9OTJ/m5WjSErpgmOD71wfsx146l8rT8toRBeEN8N
ZnC0dzcBgJ7/y61/YGu5B18I0PUYHpHqT8MMYhP1oElcl1uXjJY2QWFXOIaT
lsSAGLBnvSqcgh3blS3iQIqB+8HJknlNxGFFR/YN60ypWz1Sn7BCKB/MXTJU
AY/RSuw1b6GAatymRxcggxAGeH5qwxUUOeL2yEBgxjml3hOzfy9alaNDlCcC
7YGb3iUd2dyIAqFEbTmAby/N8u5f/Uf1L9Q749CYmdPkea3z0OdYjBTdsQpa
YNoaRpn0cka3I6WAf7yTR6pW937F2lfpRSlLyE4jBi/1EFG5tlmZhv5EGi50
9jVFC34i7sWpWC3/Gfm8uobGrVrGd7CT7RYP4M5mSAKxPp2GMoTiWOBdWs4a
9G8nuladdRaR44jFIxxr6KOXcwjGMvCOuZmDinUGn60SoaCch09fUSiSz3uC
CuLZHIEIt08lKm1tb+ER8dlWJdyW1AjB2T0ACne2yCr+9w97Os9Pqsz4gHmR
1n0XRjQmiBLN42qknSsu9zmD/wqFisY2x5ZVN5GNiQioTIVuP9dNah3/pDZ3
fgb5To6Q357yLtJmg8BmUuhCJqIyr4pBCMXPrNdvAp0eNKDfUxHT214eM0r4
8wPEsw5nDzzsyyQJJD3gOd4uNMJ6d0UGPSxi1C8QC+T+An79hGfsm9FHtNkz
36Rx6h5W0xU9YqnSMedPDcbIGFYcioL5GY1IBO1EwSF786WUZq4Dax/FdCqO
tFQcrx9qgZq2vUIJacwmuN21LA3QQAJkz4eL/NX1COO1OZ5C1DcxTPKAQf+1
csbI0U7Td4kHNyRQeWgT5ORnltwGcyxE2w5vioPtm/kG5ENlsgBOLXUEIOIO
kkEXR+LCm4AX96jrdWNB6KSGSL2X+lRO/PzbKqvhF1wOaJG/M+nU3YYdrfn2
5FceezGMIBkGswh26Jm8uqa+0Hbun35rVHvc5g9bxZmFONIH6iD/cmEeYALn
ENG5R17aOO5VSqt4pFHmhNbRESAPsy42irNM1EHuQLrGTyYLQpzR/aB2sKPS
L5oI2nQuCcbeiWJ9ewgKIGCPtxKEC1F5IhgP4WhzJSNFlroeJ/uNG50NgNFB
Pv2o0h8Rl6Dhas6iZGn7L6b6o68+4z1eya1Fz0RmGplVuIZmDrawC6GhgFuB
VYREEwkEuzm9iqsIXOiGPCU+3WSINCXfoghrBWEONHPsi5bscFEh74uchIPd
mBIFJKFdKxtduZlXsYBkhFuQZvIEdIpH4W518vPiaZbRaG9Bd14kh2i1Usdy
R85eE1TFf3xwbdtaKzE2tqtvUhRtKAI+8fzoB43+pe5Sai27i07vS/hsN8oM
qxomE2P1xWadAbMrAUtknaJFFT8Whqp86WcnhlQe+0DD5yrxcPB2iAJgui5E
Iz51N22EcxIifaxNdnl6FmBE5gsUR4D6ZItE8rITkNqyGpA9rKN7ejZBv4rR
6JXJN0QF0CUpP1jaMA5u+JE8beTbqH+z1jJm9MPov5yVWCUvG/VR0MQxsCkd
pk83xhrnM7Xi1Zcw2wcGHdafKqUxa34U6duqstOcsUSavJ6FfSLfDn90s7Aw
hRZ/MZT8nG3CFzGR2EB2CMIjT2nj2cWbKGdXSczCpdR1JvfjgWJJ8fB/SrbJ
l+uh8WTYJkAUnBzW/JXokBH6QPHx1+W7q9UtgKnDYbcvoX+lkrFvSXfUuxwJ
850aImBgFlMWUmajS41FVhY/lrLwhbmVK8VtR6Xdl9IeotAjEO+WBbL/N0oT
i261E3TcRt6zUJOyS3v3nynyEx4ldUU57Zi5EFBwxxh6sYRHKqCTy4ax3dPb
aYwASrt8IXYMFj7OvXnDcM4EGNjDEuduHDnyHdn5y21aOniKBLzlh2WhVQw+
tTrl4hdlETNfTXs/ERrXahxZbhRLvLT+9CYc87c6981/56g7AjgEZ1C+aR8q
m8YUe2NesQ8h44zoDW+Bh6bA1VM/ceQH02FQLCjNMk1gnAP8MSBl8yClc5wK
S5C3Js6VlITsmuzpxm0e9qnC3CYH2WRLEIt+0H6pfE7m/MiqnSusQ4F1blBN
znNnTekD5G0GT01flujAWAqgt1MC3/PDZvFlyg6X+tRz0occXExoKG6Y/Xwa
qWw9GWn14dyZICVBwCiMZLGtQWNWFl4J2KvBZtFvmmCi9zj9im6mN4OC5UDE
zqIv0/sW8y23qyYsW8YtbXETaUhmSrekaSKghzeAA63pPQFbtaEXIerXLjF9
Xbn+x+IO3ORm3jQgXW/lHyHczrwqKfVXnHRrWpPsE9aR2L4j9Ahn8NlDQTOP
4Z1Fr9Oz5UUtF8Gkaaa8neDmmj0Q/9QjwTTcg8Ky27SMLVUf+TP2YjOAsir+
t7lddURJxz4sfeTvv0OLgLsfSq33rDGLACm7Czli0rKLcjxEabdwU+oksvu8
ZuFEzSOoMNF2f7qbEgzjwAbF0qmn96+6xDNW0i3QXFCqMSctucZuiyCoXvl4
D8NT2CmvlaDFepI1WlB5uPv4SckIFqh69R0Zteg/6ocJSYdtfDPA/SC5TRnj
xMBwhyWHOXPgEdk7DKPJ+kwV0xKDXlJ4brTkcPP8NIovNXnQaA3a2Sqrvdvb
iMUlYg2wEvrVlRO/QSCM2oklBZPWZg5kjmTnVXoESnRLk2sMz0sW9sUU+F23
yvGlC3iYG03hEJ7ncZn4u/vsj98SXKbudPGmf52EpGc220a8cr78g9iySgqe
V3j1UqPva0qG73dWhP8V3VjPCD+Rmy42ds8AItzAiwByPyAfeaue6oBid9mX
MMNgUgNG64kPlJ3UFTeC0UinC8aXG/qizP3Tiwy4h1D/qICYTgBD7fmSoLZt
p+0ost5Kkk6P6+OrFpIH2kzUdk/3f5oQ3EJyzwYRgWTmpVSHJaPkYVzuEda/
7d/NuglA33cSBHio5FIIzUn7LvZczOPKQESqXjAawzR4Yo3ZMw4y5OeLSZ5m
tZh2iWfqrGiuKIEEwe6oPS3L9AV2RWBO/MV2vjbcBlbwdrXQyH60ajLECSHL
kHgD63w9js2zSHkmQ4e6Ac+Sg7gvujSvf2A1nKDtBtYV7vgoN54YEFVZ/rZR
NmXDZZmqcx/UVoyHjcZ0QRSSsBv6j/Xe/fcVDNJWgWJ131R+OdvE4+QIAvsq
WAAJ177I5TAom8JtbC92gtKTv53kzg/mR/3zO86i8DVLeux2J9HHYApGMTig
RzWMhz8TiiPxllzDBKOYEw1IF4EfoqL1ShB9ZvDdsJLgVhoyGUIexahcbWlY
EJv/yNU1vRdIH3aaIAjBfSnpo0QM+ab74Fu55AV/nAPeOrLB4CqNPAlvO6oX
lWp63H06U3NDAq35ql5jRy0Xniv9cqcKL00X7870C3YdjmlMeXMTdxSkLi6C
J41eJtM+NH8OaR6m7Box2O20rNCo+SR/wRqrBs254cZ2JIPsHllbp8M/IC2j
vrYBeUr8ZwMna494a5h6TrL2Gy5KrhoZWrtkZltYq4d14vq8apOQIg2scMjw
ANoWdnl169xrzjS7ArMW2lVcUBZstb+2oPFbs9B2lcdz/A0emkwijqWqmWWQ
m5LDMkoT7C77qYp1OxaRv6VifdDEDSRr+p/BrUiM3qXFMCHpZJaQFafB5oFK
FPz7hAl71Aw7o2RIM+RFg73mVj5Dh73IGoeNNrYhj3uw9X0XawgXVmwb2wXA
foCMMMvdPc9D4lxket32Y4rXnbIYMA1Tqfkc8SXZymKD3MFT+ajoBOSOKRlq
CE/2eKimBe7el7fLAS32O+tXnMi+iVtuzCRBfUMNfSwn/YLaY4ztQD5rB9s9
tUs6AKr9ZgdxfH8IR4MBNXQlcmO9AbrsSObtrSlcgAP3MtuZySuK1GfD0dzf
0rzX2SGXS5gTZi9wMYWOmwtXaZEJSMcanzx5I5vkwqZ7NKxFFBSVibYxFYjd
8xbdhXmEyr0MaqwgMeK3/0qPTvlUhC7sACI/npII/ahyNjR1IbnXG0u6Etsk
rPramYx4tyD0Cra6pMKitl5RMKm++/idj9PMB0Gh1uDMWe8avS1Woba+U7o7
tyot7Ys9YJPXON+PSGHQJa2hfHoFdRtph8+h4OMpng7epxKnrW8mJHjgj9FZ
My+DDE/TFwApAVkmlxQLqiD6hQdS5BljDwSdUgjCw+cXY1eK4azFxbCPUIZ0
T5wI0hGtbUxG/R6T7iRVDAPYZnqO76Rpb/4ZtCyNvMsgTl4cgRL9+QfL/EoC
1aso977dXhArx+ZyiNTkuRS53FMPyrNiAY+zqjhAe+3EmtzcQUA7ygUOm7zg
raeB0tFNtbOYNRnf3NmSpwaASsYAnda1YaH0Rdf/H667lhqFg8ZlG5HQUT9Q
8N4SL6nsJCvQmDDYaB4rCza3cM0Wztqrll7FlzJf8s0YZ97GHn0M6OWyZXdt
Lp1FM2LPGa0u9DTaXX1Ri25JtXVgwxEO5Y3f15VvQ9abugZfM7DSfsqc2qxe
3VjGEuE/GoAfqPtjExBZHR/2tK6GrUsiAuIaKB9D/x6eIn5bmLqdUEkhoojF
XUH279W9IUdizO1P7i01VBuiyt1FDi/iuGwOFK/X/B8SmPEOOsHevd7LbgbK
FTjxBooRWujHI0Kkn53mPayoeOsjZDZsKWaKPFJhE32hdxrkWF7aDhR8uh24
N8cHbbtjp6z5LDMcP0Y64EVNxOfRV2/HZeWgqrHG18LDJtqct7yY6c1vOECR
GJwT7TGCWQ/hNCCjkah7oR+i/lJvTT7aN7jS8onrkvzQNAqKEJmX54mupLW+
9KGvGrl2IFrj21Bw96PDstyasOeFtPpGtJ4EnhadpZA0/wXjyBAv8gZClSSr
HyQzr3YXTvRYI5McSgH7r+KDjdYQbjnJriyQBJ5q6cPB2f+9KrV2zntO04NM
5niu4H9A8/iu7LdQPDQVmUy5JgLwLhOxJL6pxhNb0+XH3RGBKWBzlL+Ri/Vk
UrPsnhIoTCtygWZQjv8tk7/RjjsQPN38U1qxWzRVTBzV75yRnyN6S9wRz8C2
8TyNTcMmmd4o+gHA3IwWnT5H6pZcw6rzWXkSk1QNnz+0EpQrtlhPjLZNOy3i
0qRkv5AkglLJBzYSWtQtUA/uv7RKwYEiv71MvfA+jIABPMD6y9tfCQ67B4D9
OAN5xc4MrisCwpanQs+aSxeEZiozptG2kKjt6NbptwGQjSvg5hWLrrk8J2F+
yeYGxWLLep87MIvkq9Ojjg9Z3F3hwfeFHrLdHW0Zyg1Hq70Yjd1KuTVvER2H
f0g3qVSprWFrl0FdBfxUeeigI3/wC0Yp5Afsc6Gdy6ZgiHdY61dosyxqownx
HqmFMKb+OqqXJ/FybGQPf9RXC8bgeaMnqgQ7cyur+u/h+LatA7TqKGUQ4KVj
MYfRehazkbmtN00Fos3wzrGeRSJsFefn2mbZzhlkhGC0TeMtBEIIGWhxab7V
kAFZ7iIIFOJT02WYokKy5gJ2kBcUldbqrcVHTGYcPqPXHNjq6p2ltN9EPSDc
76p2wZi7Y0WYfAgfZgiFfIsVe7JMDDZ6OMNGH5VfJv/CQDISABL09b223dF8
DdBjJHg+9+tWBLUuaE9cvvodB4m7nJDSOYYj0zTTUupDpvRtOGbFzoLShD9A
GtgOt8pNNUaWrL4WtYxfHvEv+FwL+Te2+4E/MbQxhpxY6idF8lCJcluXQnBY
GDDwTZQVxgj8LvlKivh6D6RWyk3+0Ac8HZvLICw2S/bveIk5Hies5zS0xBaD
whzN3X7MiHa7PTl5o99WbOj/HT70ktliDwcnBzSqjBd5jqlw59T1x6EdfN/6
bn/y9+Vs28E1/ljUxMH6LTESzunMMu88jMJ3sLg8NBEVIwuNFx0nmT2AtfRk
yvG1nYhRHHshj8ipJiP9j3RTqKV2xnOZvETdqrLB1ze//icPzSwg1ZqAGpEW
jPDPVVw1LjJOyuX4XgMLcQPmNudY8w0p2FhegFHFEpeNafF65a+7TtBErkA2
gUXdGFyG0mmbr+SG7/WcAVRD2WTaz1L0ikd4R+x1i+VsCb+cBxCWUPrgs7Jl
a0+ntcf2uNDm7+MQTeFL9wd7603O1bGBAEVil9GIbv1tH9Ry3AqTzn3994N1
OR5rsJNU0CDCXaioD9XwTcwR1YvHWCdbO+LVrQzW2wQMokL+5dOXy7MXUQtQ
JZikTio2LUQoLwrH59Os/Jgh0jDvcCvdgLsJ2LFpoLDl6QjqWsavjz6mIxLU
bnSeMMqrqxIDyyR1lM1KevWwG2dGg1chks0A0BGS+SnbRRxJN2Vy1XdyHq+/
3hIxT0kS8akyZpIfnKZCHa3jtYkyAzvzAerXqTvhcJdI1kZ7nf8TD0qedXM7
GfHSVVIadIZlaDGrqwMJVHXU6RmauQtv13g7Ez7mDkQRfnarMwC/8t1HdSTK
Is2n++EMo9JPMqtN/IlYYLv2+QrqzQhxl4ietW5lYFSjlNhzprlutDt6hqJx
bKc2XagOPTOcnzqtuf5dBkx67eo5rstwfCqx9IGujcepXEmIoiSX/3qtV3Ei
hu/YT0a4mhqJf3OkJ6nXhxGnOOXErIkrcDz9ZSSfOonkRai3AoKrp2qlfj/O
GFF1MfE3p85GT7EXZkpInHEKZt19C8G0ubWqq40tMTKlad8zRGULXKdJ767v
gCT39bp6PX0XZOZ9RAGd2URnW+5LY6ZG3qVCLCWFtL9ArwqbwODAEu6ezl0+
N+cuQc5cnnF0HSlRv/FWMx5sl+epautC71YrzmPNmE2j0J6J8AUk22CqJOYw
7cOsOeHlnc7Wav3aDMmzKP6eMqT8cchkyM63F1YD2AR3vkZExZwO5O45SUdJ
dRlrFaNiuwp8dEuJckPMYuhydfYHPYVFU2JbuX+nAYncYHDE50teKoxXmncu
6SPbYaZ0QOdnQ79jd3UCbM3HR63nkIxUWJHQQfP3WrTyldJKcT4rSRGnYNrx
wp0mabStZZi+2Dv0z01NMbuVQGIwsrDxjq+5aalBJ1EehK5XF7nD1Q9NbzI+
8p2iaM7m0l6FjpShXY9L3GRt+RGZUHIQQ8MzTkriFJtY6e6431M3hh5nJFfR
khgMO9E3j1TttEAZyB9KMcVUh8D95o3dueaAvMG/nSAgwywukOpkwL81KgIv
63t+N5MMBZPJyUZSUG2tXf3WtbeauVFdFLMUnvQgVaQ0uX4Gy/5D3QpNPw3R
RCA1WnBDqmiUrY1qCOTwBpaR7jjUSGVCPfikbw5MlsRwnZveWKlETbp2Tq0n
GUjgIGMIJHc110O55c6EELNtYXUGVh6kmJ4FuqqMCq/lE0yCkEog4H/q7Qdb
vLoDWwckjBq2ZYlACnUiQayY47yyJho36L+5yijsSUmUKsjEkzXxzCrsSVaL
a8tNCTf0hYwPxNTmm0pcctWp4gGRPJ0h69UHiPnLQN3EMegiSLQ5RJbXwzLo
sAJbYEpi+ThEK3jNm6fKmGZNqejWoWqB9vveC4QNmHdNbE2ZqRiT4mae1xKf
qn8rGcj0tSt1XG+JpTHtgbqob17ofar3UwvBkjHNbTMkLonQ4uyAMojxfAud
wyaeJrggkMSq52iz2dftbDjgyA6bNY6z/8CD4SkY2g0Mk9YwBysrD2WZsM8K
YDs8tVi0t4PLvT1cpBEA5X8YLYXqedRD/qFd+tVFD3IkkX5WxUXgF/6j13ac
g3nkYWsOSp4nuYlGCxATdUXx2QGPAmk1wdOEw3vQjVSfuI9MQt+FezAD8GrO
lpP25ly0Tz2uePXiEDIn6cJBcDD0YDhgkWUSufWzDZegjw/a9jjaSvQ76yMA
QypQiw0E7uihnAYKWLoMMfTgypCLGvqdakTgX4e3V7VuXbpHNLVHoYnIjfe7
GspYnWFP0SSGJGMf+3GjrbAvV5hyxX2mrwjTr0md7HXhonb6DKnrECz6ok48
I++MU76YQwgsJWecUpGmqsYuWZWHGwLVu0E6C7ylBgmsSB79z6ixZh5jeoUC
2sfyKmhGZoLSdJIFY9qnpLTOoNbYU9ljWAtoVPl0LHiGsq9wAIR4ZsDQ4oKA
yT4S2i8pAuWsNAGnTuykik0nY5IvFGvK/A9/ckhxjvI7VxoHiyNTS4pJEjMm
a3ciPVYq6Nb+zyb44UrgCfR5abZK2pS+E7nYRCg36cx6PTV/9wzjpmXGnV63
2jbtGcKQnvy+CzTXgTzFtznLinT58MPEH0S4eoNKPNv/huNQDqE81D46+5U1
Rj14M8819DJp7IG8EuF+HEyCpqV2YYw+D9ShO/0N27rTwnPPlB60Hp26fWKo
pHfJ+tE/Ea6hayJ07iVWvInL3mTRh0bEZpsaVRuwjWLRn4pFTVwvrAja4MUg
asJb/nzkIPm54vefrGSPgfYVw9jT4+kcLpZOloA+WSfmtuefF8UkMKX0HXXR
+b0aHEn45FbeOaTIgEoSFG2JoVJ7xW7cFIY6AqX/M+rJyCJsoHfFYL6whdhg
NeuxSb+l/HKyR4fjskccS2AW9iNrf/J2fmR2DCy31Emsh7MGGqyzE/P27ec7
5+lkkhcuUBpBVPp0KJaF0Y9Jxe+ts9pIQODn+4/2jw4KyjeaYsqPDJw3j3Dd
Fly2c8JWxns27YIjSZNQl4GHm7rbJ7DzUv9gxV7VqY/FfGLl3pH+fJ8eY3F+
G6/cGy4AUnTIZOD/oFGidRrhMuiT15YIC8wrDFpbeO/A2aWJbDlg2xSDBlHu
8w7Xvb2LBqkLK8qzkSFm8R48GNK1CuPWHn2JCywQIE4WGP/XSyBdyYYPuchU
gxuHV8QFxuJICkNOyXysgrIgicqWiInpA3X87M4giDxeNLWlcbXVHhjEVGZ1
FRGhcKkJE2IT5Dxfo2xRrCx3R6mwJNp8lDjLyAuc8lLS7UrOs65G2HPsQCgb
gZkYGRPpat+Z8Lo4ihQaNsJFBiy0EyA7IN1oMKYW6UOQDyu2nj/oMgAkK1MU
1TD1Za4GSWAf42P4L0Rb0eS20nfYNSoFkjQZSI73ZbES0uAj8UOSESW+Rj89
i7JCfZWH6tGUx1sS9257AueH6a/k8fwD3BPwRNJsI/6iN6LupEY/BRSszUBq
zTOet8CM6X0ywwyv8DinenZi3A2ezAjKY4aKWo/RFHAl0G6S+nQM9TASGyei
MF/SFFtBjEEsq6L475PeubQhi2HrbfkuosoOd4UbRUrLPfgu7HgtiAHq0iC/
dcMwZz4Zq8PUHH5r/eCh4sFkv5YwCWrI6SLjGDpWbiaPkPbRfWu99VFMhN2w
SPeIg+u4df9at7ofDyk9UcZdk0Sfm6Exqey4fBS6R7wVnCoZxF4HVeO/j8SP
20YOnAg5bHU1v8u4SA3chOu7iYdkigG9YayhABgHUe6CpJh9Kem5+WKbd++C
c2K0wyOvQ/6zIz17ohcsVAt7NYhDuXWwBmWrZFieYJ9zSuf0b2wNY+4RfeuG
ZceHAEhSZ7i17toF9FZrP9SL0+r1ADDsl7RMxpYifO8URNTw8lbFOffiuJOr
ROgo1zouH1RfR71zDn7067eqGwMKiyd+D+dng1eLBQxkPL/7aTQ+F3mnKHtR
cQo2e3CvpeQYvSO2c02TrhnFn0Xf8nXZ0vOaoSk+YyNZ67NGMPiySTui7+RJ
rmRJQK2R00C3upS02+Ed+BFYvtCRUbCanBZgaL+bMRVB/zkKFbhdIfQW2++3
N/ZL3Unajod7JMBGMBJNuVNuIruDLInJabnrMLTACR1I1nzM21X7YmPKFss/
yi+Hl2u4ApELCeuykKNkC8WukT7nnMvyPkzIi0Hvl6QC5LSDJ3sE5PKhzItO
OULLuE65FQYh6r8LnsP0Kr6DbnoqVI6hXsC6rrHgJWnpXpRP5jRLb+7Ft2re
GA6hJL3SpBjLkAhEAEMo49iQEO0nUmmV5nL8n/afmNiRuZShaG6r9a+8apsV
DopeqFUi9VM2UyvncoplwFogcVkS5av+X1JYp+akGmyoAxeZBVJw8upMBhM/
PsMRlUPeGT33uj34psUrmB1gcqOTdziJtLs/r178uUXczNrZffF8yzxPwi/F
ZquLrAYcTXYLxqRr/W8avj1G2cfN0fIZXa/XhbjTfHC5+rJmL5vVd0SOFlAh
v0KSkGuLuST1l74inKT50iSPU4FN+VnSCdE2Nhq+QdwFKfHjJbWKBrU3anEq
rOYALsWx8nLIrKi1zZ0A1ICduv8uPvGevxVdZ+n8s3chj5Jn3kD9H83T8vf8
pBGRo8COFGGj9E3XaQNeBCzf5yQpJLW5Endp6Rjgn0YRVzmXkyu8AMMhjXKa
CoPHUdZ4KDgROnpWbVg4frr3qpQpoa0Qv0J7sYVYKz+J5P3wbjgEG6MllxbF
877VFqIWKj1wBh2tBo18nGa3rBbfjvmGIumPKnG1tJ4oYoOVyXaocUG5Vu1c
yZkyFrA9kM2i/8Bc/CPTu3PXc6g+EGvNEVpYp+cyt00w/v336D+W1q3bFvdR
bb2ogcHFDNu+gAQaAZOSP3b4N3sbEs0qJRWjuRiW1gb3iiFn766lJEbCCNBF
r5j57o72nx7y0Qrwh7qlu3lRD9783mGKX7JejbZoBGVUWVKzvaAymm2toiKm
0nvUS+1Z0RW7UJtDe4hJz7xZzsSHKnKFmTRlCJXmKMjm02p6/JIjm0aPj4d+
+UEkmwhUEW+VC/T7WCOk+05pjSFOmgveBySmZZcPBU8g6aWw+VLgF4TDula5
aTFWL3ZG6bDN/JhurB0Q21wuSpOeyQE+OK1TYKv6tudirUW5XQU8euFc4rWy
+BhVdwvW326Cr2aS/wg2rqn9JkAUTdMk6VxUQj450TSgzNzPe8+E77g3hrlt
jA7T5AOw/qGobvwRfq/QwJdoOkBm/Ft3GcvtVN2Hs+5dN35SGFuJdXtOa1Fs
A4c8Zkgb7fBXukOULp7CWR2Uobtmup2IT/ngIONTtkXjz93SWcbzmG8GSmU7
ReirR97dr2jfl6eaQXmnKgYPsQ2DtWBDupUZmGskJaQYCD1rGNi17K5/J5sl
qMsSEqyIDUXCLUKms3/Q2aLAKCRPRSMktTdZZuHgvaPS+axXD8shFs05E87t
60GXg67Dd5fgs1F7f3c7e56YwveQSPHjpM5wGuFIhCUslorhrM6oXQJH5y4q
PF25LsrAknzNWg2nCjh0j30Gg8dxPNBIbfiHP13tTo3MOFsAz3DM94X0yA58
qE6n3N39sDc811+LdzmVVhgyqlxAudAsmnqxU5vm1UKnvjWr+GXLvijW6qzc
+LDrc32LxPhi8LWRN5lDfgn5RU20FokyDOBczjGAH/zU82DDcN7Bf9kk1syh
mrC03AIInMusqwntYL9Inuj8/I+z5c7z2T4c/Z2umyZ/dSN6YOxZXFXm7FX9
TAohv6cdsf2UcAu43QknIsO2KAy/ye7vsVCLH4WpaWtalke5acHgXSE7texM
3QcOizbHnVeiQT2CyMfvAYZkH4Oj3lcPU2bdhykDtCPhvLqL7AMbB6ogXfXc
nF9rg5EX0l16OBTvhG5ZqUbXC9k/jsEc4OncxLTISBeaA1Y0nFoBWQr+MBcu
/j5oY9uH8iKDR45fALHgWUvT6d8LhL/eCJwOlcHnBFOopNsALcJpS0rIY3UP
j8IYcQHkuFOdDRT5dlTD8wpvEWuLFjocX3HAnIw1Avg70fT15Kh5N9z2kScu
tegYFOb8vSHBOv0GLnMKAkZXk5BxlixGzqOQISIH4JwAGPH4HSSTb06YFrpJ
5IelksCjbE+DQDsQKYsCnulYYfqcAgNgzGigVIj3FMLtoWkKBkMaaEToco1V
fD6k8xzrVqXikhpAbCVJ13/9PIkqrKusCamHk/Rq/dueF/EdnMl+dxmBQtvR
RsYc9VKiiPdKCXjtNLE3ErPTEnhFSTcVHN98hMKdBcQ0Butb5b/7Ryd5Rog3
w9oHPdqMujHPcyKh7QwTdm7/TQpPswxyAtnN/kGgPRQkgE8evo7XIJERSgXd
EZKPe34sZ31X5iVTLItU9R9ADmgVnPA1vfVynkiVEOXxaABAQPwJib4ZugdF
DqFbBKQUwjFqqe4C+jlSD506As6C2u6oEx5WtxIJmyoxzQIaVHF3Y3ycY/IZ
xWvpVENHDqKbAIwIyUY2HU8o4jPXX36yCLyZ0Zf+1HXHV/c2wZukhlEyaczM
g8vtfqQlUXKx6HOoSWefM6BCz/DljvzfftZEBBbTssOOVRxT370h+SamNZOr
/s0fo1ok1MXetk0gZqPsnKcmhaPwrmW27EBS+tN/HxgARwWHJuxdeHMryzZ5
Rere54nV6nimwml+umE5t0MzhOrYSQOf3pSmO+FXu77xkpQlYv8abo6i62c/
/Z70N+Iv0T8EO8Y5BI9sKNTAS1/aUONW5EdTMEwEaFcnehpFB2n3o1/h+K6c
k+4yGAPOg8087mik88bQ7UaADNk2dMES0LDzljOeW5IUAxnOoXlpShC0A9Qt
d8P7MWYtE5IFotG6QA1gDJSALdtGLHhZpSSrTs84LFM6QqH17JXO0uFYgVpC
XGlxGZ+CJGE6QuKsVVX9sYJTCV//qSLi+9hBNwL4CxsydADZ8uyrbv5ImGS8
tSeMSArXabSuUWPVNLHbV2KHoa7EfxNfDHhr8YW5RRxV326cs/XX0jeBqxFT
3Q+2gbwQwHMLiVXdizK9cCe9zmR0xMH/bcL33eZ3G9fzK7YdDVdTZNFVYY1B
H6VhKSNcBIWfhn0/TAZPacXC6WRhGME4KS8LXa/xYKNURvkquTIyLzjqtcZB
EfV2q/Z0CRiqYtYsbb248o4BjzKIk1SoPUOtUqCVlfDFRzpOwCU9B2SUayMU
2FTxQINhV1OsQLnGdGoA2m8795KiofLDGYeqgRg20bNJg9y/QVo4sJSJIwFA
kn0fMwfX0bo+v8XgCaT+JMYxHgKwbCWqLSFz/DTnS2OrfnOj2ntizZHKdohq
rhUOewCBAQuvF0mWFpBW4jxsLUmCKNhni/Kw9K0PpLu9hc8UGxhPHtbiNdt8
a0XJ0/UlE7PfOV0rc3dwdIAx9gZ2JHH7STF8oSoJSukUxpXNBkV9ZFI980rj
YMLoc7k1B7iGzCi0wAbcHGTyRwjEaBGC2G3aVzvyG7ZljgUS/7qgYhaFDBtR
FxzX7mLH4pFZ7fjJLk400CMadlB3ZLPfxwBrBiAnJzxMChVzlIDc7Lz9zvoo
1flucZvM8qaKLOmt+IwGu4JpyOTApN2bZijAw8gxbFt1W1lsjlz7HfssF1DC
HiRYqjNXaMX/g2S95c84Lxarar3CtMlT/UmF6/xM+fZqgBAbzSQETT0dYRIC
48Rlw0Q2OvLL3K/iuUbabVtIpbenkSD9h4OljSOLPnwoyYTCWOdnPykXRV+7
8T3fc7+gsbjNzgBgIN6lVuOwZOVHJ7TDld6YrjKeO0P2da9xJu7w9NdRd6wP
griW4ov+W+0TRN9i95IMDo3dqCLr9+nKrvi6Y5sqHlZYnT9sW66uPk4IGDil
6clTG0RtZ6fUSPc+M0cHS+8h3//nvWlPpnV/Ol35wVoy4tzc2T77USq4AG6e
rZUiVeG1roDQenyMPQXVJapzMhV0ILSAd2exsEcVbXhCQ+DJpsORrUR62Ye+
gna5ESxeobTMN9NTXQnlsYCPqmyMyOd2CIWiSCaNXqUpTJYTW8HT/tvdeKpC
AOgrQjZJJ1mvr8TQyTdO/lE7DAhEmvfzRC6YGEyvWHCRTyR0efN3jD4eAsS+
3AZPUJAZglTfpf3ZkO2yjsv0VNYCMAcr+ySPrIbYWAKCXi22bmAsF0BEUFJF
fxkLsT/z3m0Uda/vRTSwr3BuPvH4KbBQuSxGRqM2FLcNjcZ+3uG7wWwQULkj
RZYN5v3Dayxhhrksz6p7ua6lNiiOrEH+LujU7fi8za08UCPr+jFDpjCJMBdE
moWhs4RjC/IIRoJjxZSjLM5n+2US/TqBRfl1JIn9vcIerf91BK4bD2EmMV3Q
ZHVziW+AhvACOWoXHQ7VRoG2ZZGI6ZeJHJdBsmNqlN70P+kZl7xkMlpKS8Js
pnyYPr3qq3hhGu92BSl9MbcjLiUSdZdk/mMRhC7Fi7O553f+kw3W+76856Mi
p55vcIKCG5vYOmdLUYaNBOK/YQC/UXkBPUhlDfRzcw3CP298dJ1fhXO538wo
eANXmgq+npJsjC63YsLciZ/oDBvD3lhzsJTsYesyPH81n36JCIGP3ojnQh06
g4Puf00/lJvgk7j/PB9bBqifAlxkChTeP5c7GezI82rPKu1SSTEAe1rNwz/h
gDXWUoYHJJT58tZI8eqA2UR2QBaqB+wGMnkOVy0bg/dxZzI28shFSZh4lfQ/
5B+k+aXPR0j/Pi5i0CpOLL0jQCnmI1yzzzf6D7AGiaSNSmMeTPy/lYYld/Il
HWwcALMsVSeuUTFifjvylk2sGJbt+7QI7cQk5O6F1R7cMYAp7cQpdFtZyuRq
G8nItrCsg/FXTQUN8gyhEUvXAt7jmdwNng5Fb2slgJjsEw6YX0ShWmLwdkVM
W8UqiDiaVa5ysarK4MOOxcUXH9yTT+Bgqi5x1L+zUWdAul8DYFU2ZSrNwzId
lo6Mu81CxE4nCJh+O7QbroLMTKtxHNnsr0hBON+jNjkejkaH6IAGc7ceVwrI
F49y7bDM97eShwuREDwGEoSOiTF6TV6ID4yRAo0dVHJ8+Z/LFBLWdGshXxS9
GtdGDAdgYEEEbnfIGykYgeAiRoBrJ16R+53teZq+Vck9Ah4mXEae1nOGCWgH
q74NJAiHytoFtYJ/WROCYmg+Yyu9xyPwavJFu/8Nn+wT2e1pLFsFZCiNGrjY
w3XHfcSn+hcCJCR6u/RcdrBJBsxvud1oGLbb3AdJlz5Oi1Z0Azv5cqAKlBps
RuTOGPb8wkFo2+d9r2X4J/6i/9TeVWpieRSAH1vtsDlk9/etyHeQU9qDgYeE
FpvUtzg1Y7eBRv6DQq6G8RP5/Mnq/YI9X16GeLLWiYafynckIHC72rqbv6ok
ctUzG0DjvjjjV9um1PvF8RRVKUTnino3+D4BAP278EMOSg15BRNdhn5AxM3p
Hk64L8eagsxs6PHFbmu4S5yZOinXBiVCh57fozAO7+ug8Z/LAD267yuthdkQ
xdr8BvJB+FfEwF5pjbiC4tSoqQW3SHpH4AG4E7PSPuKz9TT01bJLwMhbahHt
ppOLiBvgs2dQ9kXg7JtRgcyua31m0v8+n2VWWOTIvUmW5qHC5SBKcqR9PEe+
g+b9iDbnpYZflIPhKWbywopwKtTjtZ4YWBRNLfBHaCho4kDhNlF8ioHtBZzJ
YdP0aoaiELdVFNicIRJ0woBuVVw33q7aqLG7E14edoY+1gSfE5FuEOFltB11
FLR+1bcdcor7UHALpE5HTlitYsNN1ZOPCKVR5X0HZn1OHAB454rK0qXGvuoT
dxbPkDi9fA4LdgoKt6iM7UK5aE602c8bNuncTTCO6vOE4JaaYZcPM1ecSmcv
FVi3oPaKL8PKBjB9a6hqF3Ub0ZedgwRLXask4ueHLr3H6kSTbbL1xceBB6/p
Of29yet/3xcfO5pLjR8q9MXuI9P+9D89/JjSZg2BgKbIyIB3X4LQcbD3Hf36
YlX5mazV6RCHR4hyft7XshOnRrvqXs8lH8zbUXj2SZUz7ZBQHqp2Bn+BjGnc
OCOj/OJjItVdG20QzrMl/2ckWaP0rlP1jSamTBAvQKCVuIQXqaXIOynJIOhL
ZJP8pJZYKgRGFKtSq6xf1VNm3T0oISpgZJMWv8c8BdmFn0wRax9vUtgu15l/
Sb+nawe8qs837o6q7rxPJknVHAcbtiVGyMG8gRv3GtuVWLhVRJmwqpBBJ3Ee
I5Kw0xYqr3BbXwUAglcGoNN6LqhDQN1kce4PvP8h1gQCOsdjlIDMjgtSieyt
ijwzKNOtF71ucvqtUpQN5fJXUsLwp/OAF4s3MO4OT/5kpvGNbg9VQcbUDnKa
kKepAcOdRJnuXThvfOVgKQGHlFfO2tmcd52+CmDk6jc3PTBvYBOksqNxSFJV
WGgnh3QVmTDa/6FoiYX+Rqzk/hGSoDamFgWOAsn4K7e0w4kScCFgdo5QTvyj
akzof1JHJlnT841VVwkgcE4rNJmhvxdDs2j3PSG+ldcW741e6HQ//TP+wXJr
OlWYa1DRtHkjATUUcI23GtKaVRC8zz6t5CmKYeRiXauj0ITL1w03Z2fw8Mkq
Bw1cwaiRjesG8N93KUG2kwR2BxerRBcw3SZQOl6RNyqNoJd+vpC8BPAkolXH
2R4WJnTC8M8e1rd9GfX3zx9B3Vyo0zVJnrx3stwwu0hjfUTlLuCmmF09037F
B+BVoqnooM5kPx9N/sTFpZOuWSIKPjrhj8x3q2PXdn8bcfMJDmpCoh+Xd2oW
qaunap6OrcE2z2HajJFj3rnOsSH7IWIRyQZBnkdjtMBanW6tf0+h91aHwlbQ
OqvZBqPzbq3BGmEQLriYiNpJQ/YG6Zvt1Ln+5MffBtCLztrMOCvGU63yGnUR
qgDtufJQ9IelVwNSCjgVPmTgThlMOlD5hdX3brK+bAelxda+I9qC4nGSX5qR
wP3NZStaP+sy/d8OHKW6NOEJRA0WAXm8V9zKlOqQhcfBkPvE7Kb/qhh4kBWN
CNOjBZdR8mYQEzy2kdQN/qSWHMGIEfEtxliC/jiWHH2Mn0FphwFJ5nFityDY
YmhuP5ljqG43YcDiN9efyq6OpW/QocaR03mDa4Dw10fEcbvRXQ88FZbbJQiH
CDs1JcWuJnxo0gpx+M3+ni3Ui9q2nGd+mdBMA4C9j30FbXP7vLZXBVIararJ
lS8oD+b5u25/oZKKWbewZ2LbhX3+iaRn6dV5ympAqwVv8nnL+hA6m7HcNzBY
gMwN+QKkvC5mp7qOuwkTXl92uun8xzNUHsccEao+qy7r79BiftXGkbJ6qR2p
WjuuW8paI8yFsInsYzyzu6aGEWeXbCKf3l5Db1JSQJhkmzWdbYcyyaHAo6UU
OVhp3LvkW0CyFJvBH7OOHJlhylgr+SMmcpmb7q6wS/NukGXhtM2OAW67efd8
nhu6SdSL8lZUye3Af3HP5HEdRHP6/55ZWlYV1p/Api7EAUFshBTaYImUTAxW
nLlt2mJh0u4dAKx6zwQzYN605NT8Ca+HVUZPbilcCENN0gxOYwC7Wh4x57eg
R3Mq+P/Pzjn8qDmzftcwLSrrokIMiSRt/BkrUYqEkberpVaUHq++a5vVwTbr
8U87MVxBOXaxNRdjSUXg38RsHLlXnnk+/RZt67H97SJeK1wb8JefiSB3TOPk
GegjRmHIISTfTpmIfUMDr4zdvTp9wKOpjG3lr2mhkiH/uCAeXsKIatzxzgHV
Pmy9P+bR9RvTwra02wsAS264Ehnud6kqPu0/bcxv6KdoK5QwY7WmlOXp6sM5
yiljAWVgn8dqX59AkaLtDMb9Nfk4dt/NIltqOmeqoNN0eIK3N93D7j2+uQJx
vZhkJLjOireP9VwoX87tO2RZ3SftX9+Jy7thnWfQNzoQhXU8MFgN6Jcrfkjq
2WXYhPujIhifBhlEQyAWVo1Y36d8xab0PUPfVucYTdaTPjpDWZvPrxfk2thc
b4JpUQLRulLgLJ3B03DtOx359UuZOYjVtUcZ1YcsL0+GATDz5qXZHSr3dNir
iIzYBkoEaVXoVFeNe1TApPjCvVMgJJLi6IdLcUJGTXX1Y4OKEMZkur/J0JKf
CU1keHUbUkZj86nZ81HKlDem+5dBRtuXjb0jjGR8jpSGd7fAQ8y9d5knhg4s
ed1PUwDVuKzbDUPUZ9eFWFzgrRYdZjsIjyneGj6jvwHN/Y3pdU6dHlXM91ZB
zCeBDLZFkIttMWWqBxZuUloo7h4D53i0XILzM7Va/ZnMCWHzTAWIQ5bh1Kdv
XfgGG7ogp/bdQZPZ6KzHNg3wO+pqB12oPUwc6JmcxWkQkPP2JlIGcJDvKpyQ
DY0u20EyxotuqVUIEFL+zfnvWnGYPdHqInbPoHdRI5Bs97zS2W5H2mWJ8W5A
R5AiOzwYIavbmjcAsf8miaps2+xUrv0vsgnzpiy68ClTIZ1dnfk+m4HSXAtd
vlB6GQ4EPNYHy5W1pDcJ2j2ORdaXdfYP+zzFz5FhOF+FJoseGLG/Q3DsV0zh
ljmSei/rTnchhILV3c2GomWjQUOFuKMNvcprn1ZgMv0I30chAQZ6W7VeJsYF
E3lWKAfM34yZdG/8ZRRp24HPnjLmlWRnvSYqLgk0Iq3YZStHKiwaehfjYggV
GbcxmSpF30EgF/d/2nlOzlpPzi9JkB3YXx+pSB9SCBBKl0Tfu1ZEW/EArrJ1
cey/3nqS0GEQ47OPbGOFRE6w8MPjeX4dRzpbTOfYbtpxPGG9++C+ygSsFo6F
bW3Paq161Cimzs16kOPQ1O2lm3k9zunZacRCmGQSUqCu0zWzOB3t+iI2xELR
4fmhjDDJBLgGv3aAYmMx0xrdI3+eNPeRrrXrkoqXL+5Ia1fORC2qksgkah0k
2wv2E0twNK4wV9JZKPP7iFnMjL+++Qhr6/1/zgRrF4M5anVmw3M8pLL9bUvG
WMln+dMdBbVzEOxCZrbjpm4yRde9FHUVlOGzC1UU/lWVPRqPPzT8B+catLGq
5xTzgJNCWvHG5POb8zdr7ek2ueUDTXgw+YpcNnSUMhugQqt2VE4bNQmlv7U+
+lc5JsKsOLa9MvHX3H5rEmJxzIC94bXU7FI6cHF77fnUptYsK2+yErGeEqFy
oXt9Ml+wkYjueWXtT7AZQ1Hs5/Fxw5cuNVWzPH6awT6y9E+2q1IHn4nmayzp
RwgH4tjlWMGmwx1xusdoT8k4DQpptendZXZPa9E8AaRadiH8Tg+TTktzYS4k
DlLx0UPngl6eJe1gJb564TfKCGYg6n/dMy8JA1bOzQgQ2FozC7QMG4kMJMnl
qreSSnva1GSoazY2zpbs1MK0y6H4wYt+rA38+mCZolC1kSJA66DJdBzwAIfg
IIaPJ+LzCbjEDeSam00kFDShHKCv0DA5obtgPxhU2Ab5mQxbuJauILY2PNee
pFdujdKSz00Em1H8E0z4fKkXCm/Vg0ChdYMrLxi9ufb6MUeGNerpwuPPKBJq
arYKG9rPA3nYcGK+1yuzBPmFG3tTrS67gmqFFeqQwprRiKydds4OUxbbIGyP
jaJrLPWE9RBFjosFiL5dTAN/HSINa/2jtxu3zbC56e1LiJsSJssLfj+5xNK8
xHF16dfvOcKSGH4hhmZI98ye1Re5kpx0MAPiUR6eYrdZjcvj

`pragma protect end_protected
