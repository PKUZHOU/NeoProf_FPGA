// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
0TDDSrvb91883v4WGrRfV7CQb791VQECsScWfMv8MuchjIliZ65btzy2j7Ky1vA5
cu77J+JYdYjAPnKxjyi/jiRycf726Lh15cJe7ALReQzInpi9eq+OGusQt+b47S4C
ryVNsiJ6gjKmSu9jWysKglV44+2QiRgi9N+qW8Twznk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 3792 )
`pragma protect data_block
Q7MMGqIucJzBIerLxrKJoxIiH9kel7p2wVverqeeyAnXbNask0BQ8uCtocQSakUa
tDTj3zVi3Lwxh+R8Eakx1hIFDClaw4DPGf4VnIFj4YFNdmIY0zzEDmdDB75rmwTa
jxZV2TKhy3G7Qw2EXS2sUiQvXMiS9hau+BnLkt1ioWreX+PvwwBvVg40Uqn2kr1F
KuyCsKeY8HLLes1izTdSxmiOoJfmldKh236IJ1BBG83Xak9sHADhncqsl/mIifAe
r0k8ihqjqbncEb3gJdAZ5msj1FPUH6ZVpf4v1dbczZH31qr08s/v/V/vpae9Dzj7
EsDczovOqS59IzLQdlkzrArDtgV78SCRXDtdEETedWNbpHtf8C+8BbEjG+jeTgOr
WY4klWdqsage2yRvYJIGMOzQH3xSolt2WeRKjHFuaRUgO6nk9f8fNf9NLVqVMyso
4cOBcTOWkQa/0Pi2a3EuZ3JlTeT9ZB0DO6b2o2i/rTui6qdFqidNrgHuD+foKZMW
yHLsGbcN2EBpd0SzPRX5Y59O8mkc55kGb5yYqgDrF5WiR/U9GZoUcQIn4fR0OUC/
hE46q+Se+ZdNmfIjV6TwK635yQtMTAQCY0Ft8mV5/OQm06kpy2gvPkTJwNLN5qN/
k3QELRBQX2XTtxw2hmbd9F04CTlGVu5LsGXFkiKUrkfV0Vy8JpX4GI6E8Fs/ETsv
mvHPX2nFycMlqeFXNwnMYa2oJu+4IXnvmInyI+wBQMrpv6pLCogOm5R4sRyr6b7a
G0if5loQEkGebLG1dhye+zUicpRclBJxyb4ejqwX3zzXGioIZofHwPRP0dPRdSQ4
7oZOq5TE2f1HbG0hpv/uZAvIUm8liSspcfOkcMukdFs38GJ20sPrdPtTJl+zWzLc
Rij7aHrwz0DTJwqAE4t1A5zfSS7jcrk5DzKx0ebYjTxalgI7+KCO6s1z/WmqzW3q
S5BP0H9rX8gDICHZds4PHiyGNKOLHwH81z7oFHFR37Sbm6fwQsAEKbUCWv10SQS0
rvl+q5+RoNFQlcvbYowlgT9Kp/xJd0U9Wdk0twxrW1zXniHyXKCtC9+XwrDyDc/z
ZHbP4hOl6JvgpHhhwdqhEPr5E2WJH96AHFiAj174U3ifHsweiGdFnZ0pw5We+K/W
8068MTINVlj1J7x0VaJdVLfKj7QphiFiXltyD+TORfH8UCPvqxJI/M01ex2Gvt9X
HkQ66SVhs2kYyAi8nG22yzN2HoGKMnii1LuyHdCj+E832ToJjHc9b/pvmQwHae3B
AQZtn2uKv2FsYghVygnKoAT3OyUZQgirf+hupToyH1udvsXMJ9l1QM4nhjJ4zp1N
7VQx1LJYfqoF7leQ4abER0jS7YMkOg264pLxsPG8MjU3L4RgBUuTFpkhKeSxeZFr
3kkzEApEQvFOK8GT3mP9Bj55mCoTHxeN92AusaqhNYUnLYaNym1xfsjY8hLvGXqO
5UpJV+mHlyB81voUTYJ3x0TrPN70reCM/J6GRmdoLuImDMPXisD3XmIStHh5YvGT
tVPHGOhB/jML3uivnepgJkcxJqgdf/D+js8NWK9FKCFEErYC/kWnDii5CZepQoF7
kkiDhxx5M+b8vkoNfu7bd6JkpM/x2TGbgg8fFOs1bBeIBz+aopbp0/OPNXX6EdW2
TNaXq7WVDm9SWLv2cTowfdzBnSYZFxVsQLHGstdDCV/xPZOwpE0zAc9oj9tCtQYG
2XB+Dh5kbImKVVMMAn9TVt0tRcD19EijYkOI8tg/Fu4GJFV3y3Kf++CGwhbklU2o
7yfYS+RpSPzOazhJkUagtxpZ1NZiDNX8x5EJv1JKEqywGm5qI3F5GIW6nApITUR7
/59CzHNJ/CvyDycQheQebDQZGzwONl2VfMW0XSI4gTYgHFANWIC/tp86xKfHA0bp
mYvQ1DZofuiOcn2sW/3bmp2tGLQ37RFoLzxfXuDLK2N6sVK7bK8rdGqHPu6fkpqI
BbXLK02WKqEYOKPbDY0JsxZYdsyduYy1YJET1ZI6nZ7KVlNv7Qkz458fBFbQr0SB
SYoLDhZ15U1mmRsLwdogJ/vcwH/KkZ56vpYa+DQnScsoon/d+nsH+VFIXEI0hq9E
WpsA2Ny5PE9muRcbJsoem6jHw8Ns6l5FbS6CdgTjD+GEHiK50uR8SwGvZxGfw1TI
T2czK/I4oTR0FKlrSzk+I2PJJw3l4GmVH3PtrGKyjkxnqiNtBLJ6/Zr90t/wbbzi
R4lBPdPoP6dHXW+tpHu9hYub9xymMxPv6EPtwRzgmRJCQy011oNdCGFuovijiKLk
evScdUPeP2u9qzCO7xq3EM69CEeUdlKx5JOhiDOTfXsKRVMnvHTwS8dcHDuSl6Ox
aPqHgNK6A/XsV0HQ/LM3NoO6LT1gOEUI23FmqOj8LSmKtU4OTOa0kjRET/U96kWM
iKzlFzs7/ba+icfllUCtb9xub2ygPw2Jl9CgpOS2jXTD+huugm7XKeNq6JbkvFQ8
5lnOEOxnqpf/Z/8p2WQw2+eAkqDy37wWA6Q343xYAgbbzEGqsrd/KqXPUAmpXfor
XvXWywNi2phFeYpppAJviEIxbz693osxMRRb7tJ0/bVqJI0fu7sNNKnUF9x192P0
NPlB17NQSl61e09pPMgSlkHSSu6MXOVsl796Ju34doKeO4J2Hcu11IjA7E2qfAXr
qu0m2R3ALpO55JbFqWZW98T0yVw1sB/Mfe8W4cgmp4UZYv3DfiaFO/G3ZGoz2E9Q
DUAlJAtkQmkpFEkVLRiFaxMFqCc0lwnX3pYA9ErmYdOzGZkFtAunCZXGi0+8E5Qj
xneeuBGu6n/SYtPli0371VKXElPk5aGjjMlS2Zs0OY8H6GGzL/wgzYSjrFUI08sj
PFL06XkSSgZkQBNK2h+scrdXKCq3FIFJ6d7MHCdW+R3ucvQ8bwQzQ7dZVnqSAR1E
WsYe4kvVcYI7+p0QXb0UrrdeZAgd9BDb5YinkerGzI8cdAtpSr13dYn11nTsdriK
MYlRAc+wjOBDkoW/9AgLfRKg5voNM0ledKoZU7rg2C2y4pce/5SYBA7G9tStHCWB
hRvKzK1X+YSrU+/F5bH/1YhAJ+HSOwj8eosOAl188sPEsuO2KxbSGXf7qySrdF9U
7R6pn4BjQHt5U0kcuoqtc8c9B+nJ1MN4uVQvgfT4F+TnWjwuHly0Zzs7DpHqzlqK
M5GbVlHuSb87FflmahYbbaaYU2XazAU5979aLFPC6IU2ak4ehUIVj/3EyvwejsuK
SqB53pzujmCuute0tN779bIpLOoz/Pr0FjyJaAYcWFILITRvodKwolr42ARo0oNW
lbG+NWj3vZQjbQqlrsggf8kOb91/G2184Ed10yy4AsZ1QrLUqj5ceUCtH34gZpTs
MhoHyYzsMBe0iqCBLrWxCsh+oaVPoK36RejUtvonqvfPqI5JtKIYV60e2IQAoDxF
kd3Jx5K+mFLiJftMmM8kINSJzb61THjJwYI6Msotvltp/UpvY9dljHf9M7ImWHm/
MrdHxJJ8gyGSErYBcCQ0RdABbxfXtBlQhjmvbOuqMuuR55b+HkMhYcP4JdyRwq5X
+N46nbxyJ2dr7ZBRjuQCYUCdznKZ3c2XXAAciuBJBTX2vATFHnVInLh8psIyZuhI
gOJYT6VLpHzscwLdcAfaG3rspc8GvXbT4I4W+DW1hUyYwm5SyoUnjxhg37cB7qZV
ZRTwOwtWVHGRZNvxD62KXdzJ33dBaVqQK0/nY6wamSj2MwnJPECWjV21kBPmdQUq
NGq1sWD4PiWx6qUMrutFyrEmxbQsOKg/Sg+MFYmoXbzkBq76N3o8p2WIBDjrUWXe
X5ES9VG9iz1LmXuDQFdlMl32lEJDudwkzRWXTPoN1alW+JbBfxXyUD420O9SsS8p
rUMquG9/ouCFv83IFYOhmlWqxGNTud2eH9ZBqt8XbAPg6ugCuhd3Iv0QPQbAf9vh
5wRoObZHCGrU8fgCkh6uV8e8Y/VzFk7Dlg3iBnS7jAJKGVYuoRku+BP+vx4rCE2D
y9ZJtQRwXOfRUqWQ+QhSRs2tHLmA/uxMY6gHxyd9jdyq5tyRtZbUIjGQojoRAcVU
hGJAXJM7tEImNvbx8v26RnBXsbmm9/FXb7sUzaVM7WXmY62Th+wih32IU0uGY4vY
11L3eQNxKGURviSPwyXIwfLwO6QweZ4+JYfwzwN3NCBUyGHuTK7pMl9ob0pthGb/
h1LlSEz+ZQR6tvY3pODn0JHUeaT8bqKXgeWRFFkwKf/MViSJwxHN2fjEFyS8BCTG
hp6ydbGA0zGQ6CHjkvZ2gH3XjYA/EdBbfjb68pOtL0jQwLprFYU5VU38RDvOFzvi
CMDqLnCGYFEgq3fgHLuCooS7+yZSu1HjgkXHYtzM091Ug7vowsAc9A0+HIFOF4ly
dFUolE5AVNMboHzm5100myBRramS80UKvj1MW3lCze7X+xVYNunXLcZFH+fTZVKh
F+pUwmv7Kr7Btw1JLxRbmR9T7cNgFGx4cHaRSQdiQz6Sxxl/aQMco9VKpsPtd4/+
YSGxK0P/9wf5wiXJqw+qYGBnmJMUs2+a7TMNptqF1nxP03jsnGvxSzUfdXbb0cdu
qaGkmr5r90dM3TKs1yOeheYlWQbpAvvaaNNtnbvZifhjL7N0mrsGwhm1d95XRUfJ
Jp35C6TVtnujrgTLQe3ILnCG0UuVEbmKa5iIlACVclDIjDawIjGY5eM21Sa0oB6n
SvKff+Bkm6H7syrtidCTZuU/Eb0NNG9JmP9FviVAfSSnH0NZJ6s4fRCM6ju60O7I
hZ1XxH7jlzg93kD/corJpeOR/wBFVoKyg0gXj7iWUduFkdhNqcqZ3V0ipewrxT5b
QL4Y0d0lFlUCfAdBpHOaRBB4JDDwGDaV9JqmX90AQbpZQaY8+tXt5zjey1sQUI2A
Xczl2UKXSnNIinRavUPP/tYK8PI+AQXlEgyLpkHNjGoMxlEdiVS3/eZAVGOYr+oZ
0HuEr2M9HevSIHsTBSGuIVkhh+pSkm698Y076JE2v68cV3W15xXHoPxEP/D897XH

`pragma protect end_protected
