// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
BWlngHMMF/rRxsaR9wiC/aft0/TzrPF65hApCz4oMEB57ztrDiBVemjBufyhW92zAWwrVUFbDhzg
/+uSHII+66U6Jk4exkaLIhs1ZEKjheEF464ydx5Qqmdr+D74K2BGQdrEFRMNXQJ57o1+RXZmJtjZ
PznwtZxMtTmCTF0xljrP2SC5EWR2nKY1lAbI/+Cmnn/oZ0NjGkgZCP21wQNMCusJ11yZXNfMpvKV
nJP8G2hmORcA12vDsyeT9GztNY1wQ/GwUF04O5vU9A4hDy15QYxkngTptofugZ75QFHf6g7ms9Rh
0cuc4kA8+3kXOIHkNI/UivQhHjJM8NE3WmUftA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6896)
SmHbXrOYA0XdMVfLn8m2m+wjvT+43+qn0wlaRSCpNBhDALxhc/2sV3T+okKWDbuVhXVFwrtFEsPl
qWG3Cu9ihTlO1cQHX+2MJp8GrS207gpMgff+r59K7L1GExBY33hhd+O7LelMuhkF/dVyQjOK1WH+
ikbCQIUFfvPRkXElFd980SBAxOOuLoIq2aGPz0aPTptg/Ecjt2RLIyQq9neRrEBiUSfgH7+l/kyc
m6g5pPN1p7apaw0RKaz97BOt2NjiDTME1TVKKVQ+JGB7wZq5EAp3aqT3NDZjkMT5aCrD4f5ADZFl
GM94xjtPPWyyHEij3B9xPK/+aPc4oJ9EMnjSFvAvTHDV2/cSyPXc41vuKadeTr1UXlqVmQUf1oGt
RR1BBeXsTuG6U4/KQ/O6HbEN00f/FABQJbWFQLjPZvaJDT4SJXbp/NBDyaOhFg4P8MyHTbFKhGFZ
qsPDQ5WXmchVVcjN0bBJ/VxqSP211YOqQxK5RDanKDdWL7qkFZs6rZzuIhlUhAw3tb+hJ3vR1Xlf
9d05OZ2iS/hrpCSQWKHCDrbMWef78GZ3iJiLyIvyDASiZ9JpzSJxTacuErdB2oJIFxQ8OPIl3TAF
IEQ3j2o4p4t+S539P6GFytvFDvx/c6mSVmcPrGT5IPgo00BoTD4lxhyIje0DvPtpbPiaKZyMA9XA
/RQcQt03djjylzi2PAJtI/zyIhpW6ScF7CRkhFEGGW7gIZk/peavWhKhI0+vNLFIDfIYPvSCko79
1U+K9ceK11nh+QBt6tzVVm04TtLOXwqQ5AV4pGNmZltBdejCJ0f4g5o9b5ZWx3BSUITjGbWM8K0V
2cPNe/URiwpb8JfWoIsXE/oTyogt1USEDGPKYbb7EMtDRZLyjJHo0HdvduMRYsifxsHr0t/Z0xzI
Y7vBzwrd8xV8UyWKhgL8jxGIhnOp4k2981wFseOcg2f5f789unzd2Nf3uWlHa61tR4v4+10NlMel
5o+MwN+gJ50lOSbqlewUrgU30JWO/tDO8R+gfYQ8NAVK39jnr4r4oJXwwgzifx4I3vwAVeKrJBSE
madxao7ymqwv4Yj1dIrME9FgSGf7s7UCSrXr9bL61E+1mFrcETqhB/z7EUSlp19nYL5FXF+reaxx
l/EtgPoTRBgFjdZ9q1OSSoudZwLMlNgFjlsMw20D3pWM7ZwLN+4bbNpC/+dLSRajvmAfzbGqKTst
4eY2ZoxKspJbxYZla8jOjrVoSX/ARSAoF1ZGAz5ixJUQNQfjs5nJ9j2awHvMKm9vWypDHvHiKoSE
onVljQ0SKk8LHMK6c1RvTzCYdYik+X0Vla8/YpQS52R1TlqBaxgBf8t41oTkTOfkefV0Qo9kWhC5
lMErt+e8oo2uNt8beO//353hMXHylKSHQYPu1XtlaPVOgtmy2V3FLKYPMOV11J1bMynWxOwTuAsS
N7SkS6s+dwJRhr1AfW89XKeUNiV8zmFTu2QLddM7fbSsaQyz02h6dZCCuGveUFcYosKai2a32JnX
jK0NLHlYh8DLAwR3abOBaxv65gC9eCV5b0E1g+5lrJLa4DX+1eoIeUsZpzdljXfJmUq+J7K94dSH
6Pogmc7cqJP4h1GvRuxjbtyPY+yo/7fJcLSeqeoaHxYjjjBs2nLF0Z1UaM+VaG+deMBLiXxnhbX+
/QfLSb+oGQjMWIIELPsS/G+hyYJPyGT40xjrcyRi1kPzwPS/GPaGMW71X6Dmsh6K6dhB9ke0Jt1g
lcgCoNFWvEA7fpTvH0G72LFcrd1tP4BVZcPWV6+viNwZpcGvdRzcpy5Kc7YnvZfoMQ3PyK8MxK0/
K7+KXp6kFTazyYe5sFnrK9ulfTecPjBnmzynq0fLIUB0y+8EQn0GvysSJGNZyhAqB578fgqULp1r
9xRI3dV2GE9gd5aigVRIxWAsrAYYP4PvNT7Zm5qEvhg20jsrEP5bmxtDT0eqHyLvYpHV9UlKwTox
RVdKYw2O/HpH1o6VHH5WZwZ1bHC4SBr0PRkgrUK13gJ39z5CbAjDBeosZD6oN+qsuKtazoKA2U3q
hQg9AvnUT+Hwwxa0WPPs5eQ9WRrl5jmTasd/DkWG5+DKEzm8BvdxB48xnq2PapTgc2q17VZQZCw+
UNTvm+yny0pyeQYZIsfGZNih5c2BtxfW+py264EgjNpmrDSUWzCcZi6X4SzYn/XmPSmScTCH+Frq
pQiIh1AZPXMqul+W2QxV3gvRYwRNcUktg8j9uC0wzdt7VV/yuJyo04alq0JVwjHzfs3U/bXIJ27L
Z1m0X009ZwVHciZZg5kJQFPqlK1/2GXpypMJnPpjfRBNKZrBJirrfO7SfsSLiLj5h1PApVmwmzE6
bNCiQGwzfs09JYgTAM3yh6bBFFIjq2eH0bBlSjlrR7bYKkcf17/nTBz+GMLYNZFAcvzFVvHbkCM3
FX1rBoi01kQF3zIxqXG80Jr+zkUIcsUqZj2IPgaUtE+1e3vyIECAbu1I77wgEpxxGG8s38hVwWSh
1HTkUMFY6RogO0kMltJOYNnjpT84OroJ5KaPVm7NEXGFVDtLR4W3Q+KncBg/VP0CIuVoV1ZYBz9G
28BHcWHlVpBB38q9Y6jZ2QxsfR79VWJbKuyIUTlbua/+VAdbeCuzx9CzvPwJj9fk3ChYmW2YCl0d
gIibg6BrodfEaTXovaVntZGGXGR4PLDLEs9le8u+vu+OsY2aaGQBNWmd8Yp8idY10DqIgnmPKSQm
WFEGGPUr9x83QGBDPmiycSM3eNiCuC4rhRkBb1zNC+9KQm7EFCPsipkFXDeqN2lNi4dncDhd38A5
PqbC2CMD3VHB76VJUojn4k/Z3habLnrlPjUlSA6j4v4i85n9ygHAm2BF7ayWaZ8gye7CoBC3uzoh
o4CcTavzdZjBleD6fVRJbwZOcbPpFYheWrVWlbQL6GhzperSHi6cR+ql8DVFbD8jLbKLQM7xm7Zc
6PjvjYmYSY4nlVQVNaXnl+g+S7m9yrKhUGghfozPmzo51dyZRjj90jITfR7UthbVGASXm5nnm4d4
/4krBVpjiU9/UPMdFUYhWJf9Y/t3AXr6FWefv8ObFTG4xZn6udorVamrPGQ6wH3Fcobg2fZ3aeQ8
EAdlg6VHG9k47WIC5Ftq4vvvWRyCRDvYo474FE9jpr8Bzx+4FhcR7BfxrSszMeB7XNlJ7ueoESJP
4CJJAF6+iEJVkfVtVkDXDZAbDvsLiUUXNX6lt7xtMTOc65OgqXFiawDw3OXTvq0BiUou54epwlfe
T1wpIFxsEVqclk+yfYkJYnFaKyt4BIpKuWREFCZ+QA0JnHZI6sxPDXydg1uMyE8SuH5/5PF+UH3N
Ir3Y62XENqIdQXxpAtlZciefZ/VCzMKKqtyTFZ7Fgc4l2G25CgmOCav8+Frls5sS+DhglCcYnyp5
Q67gNL3yWfzfhfYj0n6LDfujwOy8qLW7VXYWO2Rep1uPJhcSRIrDvbhT8XsFTFpxpzm4S2IVjbqT
B/gkYSbBZHeqLAiEJCMRhGcC/6Ghb2VECgdM3eUaPStWyqfaUbJnPsRnZ2jrMqKWKl05EspYd8Ah
T47ac6wzvuOTqlwSnCqFK8TMorxinF29ldbTEQhDgckUSiMzXSj+BZK1DYuLUwJDMqwGGfkCkWCE
ehGkN+1Jh5KcUPVyYYrBECAbd2ick7qz/k3o43HUjhMxyrf/ojZusaO8tPlqw4pYQcNEXlII5DHj
T0OdVyrPv1PGhWBSW/fn3z4C7Kghzrwypvk+W6uh18r5AwwuiV9QG6p7191ubdw0pQpHntWgh2E/
goXByeZqZ3BJjwYpHERvwFYh4L8ikpKws6UK+wjOQXtQJS0KmsBSIja0qwBUproxSXhZlYGm63WE
LMz/wf1N0HI+u9kKDv2S+XcuznGzHBLOu5uiDjz1MkDHjSNu3fBbIN1Mte0DkxXOeTKO1VSrihtj
S/glbF0yvjK0moePd43tlVnlRuHbcXBnpwP41pxsyNw4WrpEUAYc/pSyzFvdCDk5raKZpFkvIb3R
YVRumcJTkfLWCuN1fAxkoMciGkUDNBJ8XmDGQIRdjaTPK0JbjFLYqa81WrUSpG/xbVMLKSqOwggi
VdhAZxZDJ252TAASloFG5sbfJN1Gt57mvp9J9heVi3vMaLZhajWOF+MeKwZCVUivL9QoweS7Bi7u
HEHfYPId11wIvmZIDy5GvEpmht/ng68HT/GTZ42yzAbGHtJfwimahxuR2j/J+jtapi/q0314EVic
WEkdc0fS9Q+pbCXD7DioKlHFuryQ4rtksG0ehY2bRbtRp6+1EeoOgAP9TQ7IMcdvOhK3qXqZee4p
8ofZQSunSBb+vTgkilY/GcJhNz2j1YVEiT1Jte6670Wnc9lD/kKpDx5CoUxZP7ZaMx+qQ5qJhCRa
xrUZoZEy3VEdqrGdTXXL/594hGWxzoq3mMgbyYDpruU2x6ORlr/0P1Nn+VTZG4sksYg8HsCLD3+d
jkwTHySF8JQ+dIfOvoljpZvmvYoL1k5JGCygjOi3K+X6aPJ+Ex9+g54d1GHIqYNpiZZxGaEgdwoS
lUaNjXnDoyeKDfbRqzPQOzGeA9jVoVGZqSCv2G1SRwT8+C/m0wrtVlyNMayA0hCYhmiHnvFSqGJl
MRFGppPEGlODkJ/lRmtbOn6FMaqCFX7uvarJvq2l4sVgznFq9VjK1hAV8JMdz9Rv4AsUxPjGHbhk
/xZquHEgDJqGfPGtEoq1pBmMUtMnAY4P+d7d03LalyCgJ7e5ZHjPpENa7ucgiLAdN3Wr1pLm1fHn
yHjfLRK/9CSuI6KkijLO0AgvYWNezWDFKbicJ1wnv81a6bvljcFmPoSSTyhoWLzkM9tdzVf0QdBj
4t1TthbMqIkPC6YGUUECwUn0eNb8skiL15o9gas7f4Y2x1fA/2d4nc0nunbjN3SpwPQkUjdXw/2d
//MLM2RTGlLTNFclWzzVIzp9A1g7m41b9z1Tv5zdqWraHg9bQb2Mtm5aQKzjrpct9dGyIvyKPvA7
AaoIvBAw5qqu6BznBSyooWnlSbm6q7PzNh3lYe+28FWaA9bI8Hg6bMq4sr+knAwNuXutfpemJzO5
zacJV7A19Tcn6q/NwFKCPsiXK+/j2nzmxXqLYLH9Wh8/AYV0QdiC3OTrfJ3nVKF9uCyWrbfy7Oyq
pfcKfmQWqNHMC9fzWd2W+MDru01Sas+9caDXUaYcs1HdEn0eO2uwr2EiWfvdgJpZpg2EDWyztzx9
kMzQs6VlMFmmwYVEXtI9+wgzhanNuVyDaDurUTe8YfD85xWqtRJjRmQdunDmzVMp02BbppY/35GI
X+euUJqo4tdfbRLWtc1JurMnUCPS9z43iPXuESXG2dZVcw4fENzFdA3HH36RnFPJYlsfHyqYFfyr
rhMAcR7yL5NCzmvd41br5NE5rqOSrg16mswX1TtniCbETYnKJs+lk0sB3pwzaVA2kMQqHJRoa1MW
GDITAySqaBXvG5SQlQoBSBNdRjg4A5OGuPL8hEMHLZMOuL+eH0UdeoJvWmQRMdC8vl05ff8p1zLy
k06+NpUyXg2m7nQCZKBLXN1mPREyDsu16P4XL0BqRzR1Et7Gt7cU1pdfVRuT+sJSGGHM6aYyqkiS
xl0iYpbHD6GTKqfgZMcAODmG9jCEjJPJKvZSm6xMTk0SnzmCWDliwVFGxWcmGQVxCeYx4VZLc6HR
jCGiwbXO1JGYvrbJgPNbIJGNthuBh1bTl0oCC/dGmVLodWq+PUlo53cCRkpsJEgbbwfGFo31+wHo
VxIy3GE+2iNNWxQibohQGohscCYqJn+bUzz0WLu68TzJ2s3IcMQgoGedXMbsbfnF1kSfwrl34VRB
eSz6/Pbcs6/mUq0ImKDFb9V2910XyPjwSubsP8ftNjPwDN68VC2f5rsODSJXoijNVQ5bkQvv6m/c
1L/xOwuzeW3wS7eGezqTNhI4OPvjc9rdZNS+4Nc478PygYnWQi7i3zwdUQJZ+o7Qlog63g2NQV7u
ZhX5220lNVqQM1IcP0/8iMwOKbK2r1qKCZzM0CQ/yhuXbguIRdo6ndaKrUdVwuREdNB5YUulgDYb
h//IjOc+1cZ9J1FK14nCtOwaHKLzMAv9aYeUmeCREADQlQI7FXb5gWIx0j89ckhWdbRov2TTuQed
NIqXx9LB15CQE0edQ5UofFoZO2VZmOpsjLxTFXYajsZlirzNLsTYDRj+iQftREAKDIlXiU1dvj2v
uA9Wif4zbliQEVPzoUuYijp0p1EjcbRZJ37nIxpgQGvSAEz9qwj83mDaw8jpwqyZ2wiafQZcnLy8
LFrKlwHW1BV6tbQMNqAxgdK8qwMCfDV9BWCivX2ZPYZWXS1fRE0FtRFCgqCkegYTSqKBvskW9qYW
JQvm5+Rd75LUuJHVXisJOK+7zgJprvp6mZsjAhv1h1yt8kSIi68o8aKI4IOkZ1wdnTsYTTZafP2/
d+5qxdQ5I/JMehQDAWjuA5gRR/lNG6sGKL3gsd3MqWnZIdJO1ld1bmOChBMfhwEhIvuoLw4v2Yhq
hwFNlR7DVVGD8WWALXlEVX5wG6XW0WeRzU2COyqb0SrKHPIiPeLo1RiFoV/pXApx41kXFMAlH8at
NvAlpoheqFGGQZcZ6d3RiNoU/ok9+mVt6Djw7yC/Gr0EJqeO//0S5TW4mtjWWMjuiXM8sNsg9nCK
iHKgqHV0Nf8Y6LSEstCXDfFggnt31q/MSi7gZ5vVywjVG16j+w/Z6pIa3xE2rEtrkXUBvptGybn/
lhb9jorJUifKm6DHp7lyw6F+qY9eEpSUgUinU1ahariOVeEfEn7Z7JD4UMe4oP+0oULYt7TnRdsz
W+fDUdMewsZ5DEWsJMzyERB6WM8TdKXzgNbyJkNMS05tDYUpqur6JG7ycPHbHdDQBilBYfE5MnmQ
4VqBfgR+rVCik2QMb3eF8QRgErhZe169yexLFwVTI9emM7WdoxGHMFIwGO+y34iLVrYIzikSNDjd
x8o5ZnW6e8Rg9SSQUbrpmJAo7Zm5cdVJU1KnlBWnQp62X5u40C0Z85U+WiTObnp4kqN8XgH0lVFM
9ug5j63lRAat9y1IWX4gYV3ZktsBCknjFJ4qZnAbLcfBWyomMp7/tbCmdp8taK6QWo+lex8F5Lck
ga5v6NLQ1AMpnD7ER5QVwVqyq8ChhiWEuo4UQ35YDDYlXQL3XekKI8ERFWURP6coI6OmDdqPsfxr
bzeUz6AfcNBXX+FUpwbxVburwGxKgTHGxHo+yqH+smNGQIKEloVUJY/PsHodr9iE/hAy+aTYAb4X
akiNQY0afa6eikNREHVCSPIglsLJnfY4fjea074WZ2VyUV4OoCW6dVIdPthZr/hBx2/JjxOZolWC
OHFRxij/qkr7GBB7whaZFDT9377CeHrfunj4XUnGiS0cnm11ZdTw5Ec1Egub3v8lSjPEyQe87z8g
An3vfIJJWH1HXRV3LCXAaDrAfSw7aJbr2+hVChU3ijpgPoUpE5YVyz3OpCHOF+m7FBZPu7ZgMwRM
kG9lOfOPHCDnoM9LhAmoIsBkPKBiLz3+h3kKBrDb5/JrPsZ8x2EUbiilYnBC5ESwXPaEtwbYdj/b
hwZ6CsJHfpvQjDft8c0kuwOQB/zphy6D4KT8RLo/FVsjEhTNELs7A73ty/hEW91pk+AAxry0WOFY
pm70rDMgZsJ3sXuG79qlR2Iqd61URY2HxkgMWzMdzt0zHbv+PAiXUUULA1Zx6Lcv2UcjyCxLkZLQ
C+AN4WtlVm+d5M1doewaxcxK4oJpYp6pr+mFn69+8QjUouUqAb1Xo0XcCgSYE1wMUve9S//t+97x
U3foK5QkC65GfOAAhk8q+plEcBtD7Zaw/SSLpz6np4v0fW1uhlk1sj/suahQbm29Dep6FuSw8rrZ
5D5VJ8zd4qbXVbQSIiBkDyeGZzTRDS2nszUOjC3avSo+1tBHKKWZh6Y4TO7WIduVv47JegPtQUeU
wTuAgekoNbm6f076iY7+mnDpT3nWkZQCyyjOpfJrnAUdONqKXboFYVTCxZ2yspytqbDO7Okztn+v
TobizxbCOWtvbXGd3aCwJ1GlmjoIxAJFD6W/tJmqlBQZSD8hoDzYM9JrIdBksN+PlrcrUNtBom6U
WS0eSpMgpoECAAFX0apfHotCCvxby0PEXL+4W/DJxvk5yIVl+a6YvKYxbL5/ufAg8iHmrRrVFU1s
HLp+CTG4IZ6gRyI1IVuNY7FsF95MTN8dm9bs8rR1Kn2XdFk8KzO7g4EHQhPErk7bOvk//CyxYcbk
FPVu8rAd0d+5nfW3SSMt2PMkdpRP51cp/d9Wht3LjneVAppq41VGoCXmLLaTOS49IjN7jEIyrNMx
rnjB296urGuutcwfgP3oXs1ObC3pE/cWiiOBeFDyTe8podJnVbxop0ZKOCMWXGsUo/PkYVmlHGmd
v8++FDuM0UIafpiljLVLy7Dub3u0vbvHPtgt6IT45QI4RqQwdtf0lvDOLRILLcn8jGXqZ2IYoR6w
NxykttlWp1YK2yodhpFVIsDu3dJEJ2XWWLNHFyDbvG8S0asAoVVoZQANN6d2Y14lj6hVbex20F4W
FYk+t88T3MDQY4nftP93GYwkdiaDno7QVU424/1bXoPH6YQwS4FKD1/WmMJD6jvop9VXUoctzXek
ubTu3Qn/X8FkflCXSQ4xwBJY2FU04rrM6uL3egS/uasTVBEsXW0jYwJFzsZ0heP/HQI5fXWruLvd
EO9UyCBjMQJ6mUZjOOnFmuDAKIlCAEUxDxSUQuO38a/DwdiZuwP5g+vF2f6WT6LNhgrJ4pbALLXK
QO9MjM8OV9AgZfOSKocF/FhYSb1ERIGrtqT1H7HduDcrYF5+iSouAror871JlXNgj+atrGq4CjCH
/x+pkD6ataRCD7GwZrWYdp415jfkJ/zNedyCxd+b2ReodQ9Ep/hSACtngckGMCSwV1G1Vtsf+kA8
VLRT93Vhb9kVzhwWKVT2yUtRDjCvYr95iyzCWVS87Ew/1DJAdcSviue7h/Hvw5uuxowUomYMCHTz
hIKov4x5pSWgC53n6QnU1UbPbGjxkrWxci0HYAAtVmRLyE8XN5efxiWvFEyQ79e4Fgk3ZGS7p1dD
qEPR02n2jn3HfOvEdGvLoCm419K74dEiVZRovYH9XGac2/wgz4l3F+AidSvY/toX/M7MqIF1948=
`pragma protect end_protected
