// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
1f9LwBmEt8Kn0VUcGnQ0Su9hrQeY20K5la0fPtPZ17NsMwhiILbB2+3h3BLTdGDM
dJpDmIHRICo+C6sRVG4rIHQVsWxBeoFRKNsPw9s+GqBnBs3yVqS5fqtxOkiHaWG9
kmH8j9YjkUf4E98g+TnOHwK715X/LrRefU0UduscFos=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 3120 )
`pragma protect data_block
O3MOZf5xNe44oktmKM5YY5YpT9nuph9yEKJhf8B6WtPkF9QtuJkGpEQhvFQ4OpZg
fY+rnMSCJ4yemoIEK6YvhUMDR+EGaHbb3I18LE1tX0XVmD8zWXGENRdDap4Z3UVL
28f/3b1WE8GD8XhE+BkxFDxnZYpsdSKsNM5aVoG4Ybfm/Gtgu83sG7zspQKFAPj2
8Evw1SO7NRgzmT/xntsxaWqp0ziQb6ULEH5yZhtmkSCdVWy93Oj8UGQo+1iCC8O+
YeImF92QbeW2PFYUJOIVJuozMfT3Mw+0Ds8ssAI5Q4tQimagXCy9ZP9Bz/GnbdQu
UykMDvkZQIxuW/DZqnaX/2Q0m/P0rD9CyD61P6be5ZNqs25ZnJP0o4FXYOT5ZCw1
9d2yw5tIjAGw0E9Fu30uiqu5ofbuivM6rb+kKIk4fkZNiKSPNhf8jMBigjuTfLks
Kuj7uwdcjgb3HpLapun35NY85m8ggADoAOW/0TFL4R1gBQXt+N44gABppos1u8t7
DerPy8RMsHjMRiLWsfXbYpGgotkbLsBWFicY5wAxOsLj2nkENshS2G5GW8r9VkFP
xsbl+Wq7LovdZH2lFDerWZ82iRZGOhGuGqPhGy3jHckTS3kPB9/eWpbfxRsNRPiQ
Fq+Y2qZbCCJzMF1o+a3t7EFVT6pF6EvOTCC0CI6vSEgFyAQzKvHZD0myaZcNGDJ0
+qN4wF4Zstq40JgzxnD9rOWUTNX5cPVZIz4reywFMsbjG3L3MsD1FBoB1jTDBz0H
1D7slqNs8sZft9BZM5H5pzzdtVR3mqMYXBMuOOKuhQGtftAJe8RKPr0yUtHaY0fy
Wx/4VTvf78Ww2CVYjf7ftrTr3I+2fLUpRaeGuGxMX2bM2Wlocz1LpZL4fwDnmKnH
ri8wG0mMyToyOS9PWRvm9xhG71QFuSuUfSBXRGdxFumBc/IGKsI+09tesruuZC8h
DAc7TfzNRT4yeVjzlM/f++rIbZlzniWKF+cw8RbZHkeTgCFRIstORk3BjD6BIH00
pl0eNbTuz80a0WIhACSG1ZvGKVds6tIKCoMtMp7XMi8C9ERFqIJR9Jvoqxx2C+h4
nUvPx9C5RhTGbdVeCOdYmpsl4MMERXwt9yPeD5EUfaHqwbaIwKCMijMCyvP+oMGC
3KOtZLS33HhkXEPG0DkmLqHigAYEJdfrdC3O9nmIYj2NuiS85fMJd68aCWCs0wqT
Wq7LInT8Ey0cqtbSbmjMZQZdhv/LOI5o2Y2Xtwqyi0dxNO45wCptGL2sk4G9IsRk
xPCfG5HkEHHroua4N6rCsdUt3UAO+24kW+eN1lpt/b5EyBpUQtaVhBemj+X9Atpu
l+J2xW7eAPgaFbUU5+xxYasXGhJXB4RN3gzi7qOlCO/04x0ghWPZgHxAYIH/qTY5
fcpVrUlz2izo/T2iR2wJosKi2PK5ygKZCUh2aKE+jdkuCw3YX1MuoR9etUYDcBUV
LxRLJ66w5NHfCPfbEREAtSPIG/EzkVkR4zUQYjVXJmHtGyJTPJNGWZeU6rDts9tS
qF41kMc7CLTrq87tlkD/gYhFj8aCNp02vQPqE46tjmX5iMKZoAi3rgqZGRvKRcJ7
14mqAEvG87U5iIU/tRAsc8T3eQf7e5ZQThmw0LpCvp9MBQRqX0qfchgUpA/fCus3
GeGL55WbVoygO00lNWXGVr2KC0e0IjfgR0DflD6ug/RjhPTK0tCGtdlou4wHhWlm
RhEQV0qAJhgUD0QaqFcQ54sBykgbn+jsdfujkNs2RSftTsB2Xp2m6kn09frqorT8
RaXKmLhEAkadSNxJtUfoUHAt+64hvw5M/W4Img98wtcq+MU3ORSnnsO3rWEqCi2u
rhnMHtNQJPWyaJUezz7fkkDMJgE0CTEZxSNZZGajYQf/1bz7rpjXdcoBZdeaDKBO
UkunzY35/U+OZN+Te8fMbbiFbwQ6gDdRc6sWzetot5I0DvGey7qmv2uUUT5zLz9W
VeXF/3DC7NCXPddJUYbMLEY1CCKZmiVP5NrEygQZXjdYKI9wXEj3nXWhcpzqkMPK
uMp39fnR9BD9esaebohgGmHx+2cl9ZRoaDEAahygOsMb9Kz0SpBS4v7pGOfXdZWV
Djk6I7DY2Y0Emz8+zRLq8JFeXSxY5+eVCabvOcLodTFJTi3FND17jGd5QgmKGTv0
6ulSbwOZflPE5hFiO6XAdIBCMNEjTjiLFr/n6Ez/2dHlU5qew5yeIYyMEWBQ5p3T
CBmvNpQ8Q8EW+rNrPJtL10fSGwuZF0EqXT+//qlGsCfde3uoxCNIdB92MMGodagq
Fsz5IKzMMr7YzeFYC65QMjB5A09jEgFNBTAGkgSoLocCtfTh8TnYkM1TVt450y9c
ROp4J62cp8LZMCkrhDHtgbzJ7tlfoI0NboOYtFSLSl/E3iM43P1byjkyFEeIIshn
oBPCbXf+dlcMKeZn18SexnyzuAw9TvajdbnlzcBNGJhL/lsh/IRv+tBj8AYiv8cX
b7Rg/WuclwG+CZ/N/BRYNjPFoRWNtuA+/8GIZcnjeAIFGwNzq+2Z+KD666FzEwH0
0n+rb+zYkNYxoDPvqJwxTw+nnAeK1Q2OnCMmHIVEVWs02AQmnuALhkJeud2SaKuF
pjgvCWn3WzE+v6bQGtD6yF3x3DMvASXnTFi0Ur6K3XThpLg8aP0nUhIRVAwZ6ytg
cFtiv8DR7z3P10I2v9Xta9WQRwLlmNRLZDHJYiyP4GjUBe5dQB+1qVKbqbYKQphy
4ozAAWiGOdX3+8kvvD5RZQzHyKswW3hp+yD8UhOFDqIGuLLcIde46memb3KA2kdW
HDoM1MQKzFqXdl3Bs3VwR30cWLvbVq7/z8TTW5jQ0eZzbdMVwKlthDD7b+TlTSU2
xCuZdw7vT9omLr2bbnyYMRsf7Z2pyuQrTILdq7MCC3pmxCrH7wtR6kgpcLEWE8XN
g7bpJum7MBJDmcLTMYW/DSEaS+tYyCR7NiZBXPGR+E/tUAcmLb4ObJfOyZYSPfJj
en5gNmWEqcQWFBZVsWWMnTaWr4BTViTCmi591xrobP3FWv6kBjClDAKuk611CRlk
JZjLUDUsDuA6o986BLJfXSo4JhA06xxriXeeo2PSDFffmqKiTOFHjUPc9ABPvRhN
SiPpB9K6gaL/htkJRict8pGs//5uLm5ycEee0YpNq4197DhmA8TZ4/vggeU2zuXV
6W8+kKy5J3onAXu9uwAOp/LlyaNSaixOZ8s7Xip+t7UBvGbhlBZBdjcYll0nFkl8
VdG6BuuniNY7YkJwRQD+tSEnVMmJH9eICE0RO6zH+BmP7q+C+4j/y8wXbQon1o2d
xAyWBfKh5VOAI0RX1AsH2WNYvXii5Tm+weJTooiiluD//NSa3Egy/wHcyYqkfvrp
c+0Wt1HCcKylBdTrjYTAuONE52WGRFMWvKUDwhxL/S3GgFOIM6Tsl18j9l99J1ZX
nv+xU+zsFwb8g1nojf6LIF07P8XrP81XxjSvR+VAwVTgb7aguiE228ov8b6ymJNM
QD1keMB2wLS1SEGzUkCYHWfmyRtOF0/G5DiDNy3rt2P53h1CzqxY2XHA92mRhat+
+i/XrgNMdYb9JQlat2luzfE6gKsaZ6N7OTzAz8kpydpjnd9E/sv6rhbbYTjRMcdg
K34I/yZG1dVylv+vCU5Ux6V7ceI2Nmz2x5A0fkjvTOev+W0XeXfYt1WIQvr4M5QW
Lmj3cHuvLAC/31QWrrdxe8LbZUuoqsspky4C1GQePnKqVDXxGE7bc5pG8vBzcOKd
IvlOiJNd9Iey9Hrm7M6sI1GyETikYJQXEaBK67oe8EaJJG8N8PGyczVq4LEUSBFm
+8/fckO0nZDMCfXG+mc3i3v4Qm6VYX0Mya8jYm7y92XRQSq1Wm+d6YHtz9usxMje
LvqBJIy9KONgUc9yIZqPgpKClOhhWa6F9laf3iF3vIe3L+Jxlrb9ZRDm/1H8iIYI
byx+z5WO5q4PtF5fjHe0xVROxfeYPVDQ+d1OyyVDQjSjmD5bhMl2JjuvH547fyn4
/UC9ZtheoPA3o2TPuSjSGaVsNgR0kizlmH7r8q9QbyUD5NWN4DGsG/cFVW/BVB8d
jUCmJnC2C1jIJidH7xULaOEabk4ro54Y4RwXwIBcrI1k6lP7vuR25vWn4ZusTo1s

`pragma protect end_protected
