// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
xaO4E5gvI5KvVZVJHa1n0HF6F1tK7Ikg16hG0nP9qYLNjFM/zqfvsGzNGybD
ehG5WNYa3lPpiLyRPZn1+71DfaplTpo7WjbYQj8k+vKmMB8D212tc4F3xrRN
56aYDBGGQq7jCCowxuZbCXstT8Y6NVSnp2wc6K3SBlfXLo4ep/CHARMwvexC
RF+uXd3oqWE+djbZ+H91uoKQIM/Rr2kMZOYPkJy0QPLM32CC/l27cgSXnRbF
elYRfRR05EbYKK/biGZs66VtOc76Qq9DpQWY6sekJhFCqtZQybwU1Fl5yU1u
k1TCsBB3PdDaXIk0Wf7MV2/ujfBmK75sH77P8jsnNg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Wuh+iVSWp053I0eCqXUCgxp7VQn/Vf3PlhXSLTEZjMsdGfs/wo5uP5sO0hLL
zT/vv3tSpJf6G1EFYTTRxdYrxjHOO8lEfOUC0RF4tNsybfqV6HY66boP66OE
tDVLYlHFIyp3j4F8Q9QJpJ3oLpQTiFlZR9l7PNUAe6uB8AG6Gi4HYrsl91gy
1ezKm4vkOlDOfGw7w7/o/GF3UZC0f6O2WOKp7apZ1HB79oeOom1KrL/MT2zJ
zIJTnGjLK4cBnBqYP9RNDY9aqrrVFZbT8wfbIJWh/faAdP/APxe0ZGuSAiEH
5wUp76k7s5IZ+Kwd03K8QLDTFgqgoacBVkwYB20eKA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bq3fDdOVE4aK4evvqtlovNlijEKu9w9HN+h/KSYgPMFm8xN9XZ41LgfXUf0a
u+DSx5a0uIzEWEKHVpZ6sgeiKXxSJ09GK3e+7yJOwTI8KehqCFXeOGAXNNlH
bYi3eixEwOccJqvZVgSEaxk8BQtRUxoF4fpsBMdzzYU3ySscCls1juBwoObd
YtsaPlTUURJZkyhuRSC3pX0o0kLNr6T7Rrd1ZRBOcvJcjWGr68iKbpvGtS4P
Z3HUkJaGf6Z8rVLuSfsuYWzGdsYXlv0VnUEL80Xb0QYPWLkaQh/2K9NrYlmx
XZdENRu17Mk709n9shtkeM+61gNPC0JGj6fhEksBZg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PR9t3tck12ZfwVu5twnx6NRy3g0LlCtI0YUsLoTbxDNRkXrqAFksxqy9+R+S
ntBZxPuqgRcpZfNS+tQPzMwhk7eBTvg4iv/WbdPrMxOU86prv6X2WzIjILsU
yy1jPlag6IMAoJVlWZHTRDbCHrZvw3tg2sqc0sH7jIfhdVPkQME=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Mq3qBJkMfotYcHY5glbzmaMIR7fWw1H8ATUUN3ixzVzKYkZJpF5Cqsxh9I/q
6NQcuKFSgo4yaJU6LFsRMDkXlSWBuXILJX1Mh24V1VcGAbzGB2dlFOPIpxIZ
aL3/JADXtMoR6H+AfBtS5rQUWKP5w6yHzZ5lpZcHIN58u/jrjI96RtfLd+6g
MIHzcluYE4jHX+IM92jG65DLfpv6XbqHNVwhpnW4ZiDWzvAiwNz+N5BN2joF
kWUG82ehBwS01h6WYYE8KKwZDoRU5weQQwuq3qeIUZWwrejyDNco1MOluVpb
mPBAbJFjHmKxSpvs3x8bsXHzYnK/Lh2zaVTHkA4XQO0YTraWeimCSgWO8UAk
ySRPraqK1xW+16bNxRmIHPlOAPOCPbn9EJf9FTZ+ASThkjOHpCXFgM533FSX
Kcvri50b0y31tOnl7sjLl7KS9PJJHf0Cuiqr8KNoS5eIK8EWwEDwccYd4d8/
ogNl/YfwsUSCLaVp5nrmem/uvpOAC7TH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
E9rRpbPgkOP/fLWEmNi6iVUzjr1HQ0gf7ngOdpzF2cFaE8eSKEiRXeTy5bFD
nY1P6yLdy6hRc38eaRgmh36c1eBSaqZhcK1vp9XUThAbtypylEkijsNl3RAG
+cGZUyabD3Mg0xsisO5icm9dHHS5xLIHg3m9xbaDu7pR/YfLPiE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
reezXqSTLBlvmOyezeDzwjN2oIDCqchDZzTGKfXpUTmpF/vGCvyhE6FHKbim
iSOcjjI7GmJeM3eFlh+aX85SJh3ST8GshAhFsTVt6LJ4P9n2UOddNE7jrvJR
XeMnbETh7VTezpNPgujOAWt9Gu9RARPcpwGCpVokjqty32pBR3M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2784)
`pragma protect data_block
tqzYkgIMWzYB7luDY7FbFUkqsw2egS22+upj2+UqG7fsgPaswqm1sM5KwXFQ
u51TdoZlpSTRIvHh5abpYKR0jifguGv8JEsjeEA1oW9gJW51aWIF8nISyGAP
pJcvAOEV0ujYCssmAAyQJkyxIePvEQxEVGnFCMWGy6znglw+TacswFErYvpx
W9z5VTpDavtXkvH8dLW/HnYSPKjlUz+zd0nvR0Pp3c2CJrbqavWzy3JiYBs/
+/60rlW1MvooQO0G/R2pX/qsfvPSjcnUmd+jXdmphRRTQ7PC5BelbXIz1AQX
+8LKH4Ra95ZVa4D0MjTJ7rO12V5NEFpmkP65LbDYhuQ3UbiEzfC1khEb1O1S
Hk06RLqkcARI4zFyY4z8bxW/bklXdncWHMQ6biFaIwoAMoPWoxb+LDxanzV1
Vk4UHkLZwgc+Dg3E3xPLQcWgITI7om4EA043xjYwT/bEZHQAaumtzgNgplcu
NaGL375GxUABWe/DEKRE1R3kA+73gTcp9PxywCwlTthrtJRGTJxl+08za0jh
IwW5k5QcWhqrt61m1g3nDL/R5YZBLsGETtpaV0tfzSEXaOXlSrTs+7PP3CBa
NNFk9DaAY103OsVECJxlYiQulM6Q928grk8s28Nvq7cuXFConQ4TT01OUl6j
INEMnB15ZY+/mOZwPOISV9+E7WuguFDtVhdgz8m/gN0doeBrcZYxrWDkhTUb
LUh/k9jkW8DLkcotbSo0QE4WGV2pM3wEW8rI/xEmE+XA4tQdhkMip+xd9HTb
LWI96UkmrTBQZrRUstNgAceRj+JjNOmPuSuEUquYTzxTHAlO9Q9snwujuyPb
NOobnUdRz8q8u5PdEzAYuRVeXasy/CvxXRlrbCzWADudwEBGgWAUg76jx2gw
TievH+7tKKUclUV8rxpA4Y3MsWyzRbwYhLxz04KpPgnG71/q72uz/T9VvVVh
ej0Y0nnhITz0J4wZ4d5Q+3JzMW3UZ9hB85A2nD4G34pjE71Q8asoXs/S5r3p
PdCSUdeS+kj/VEZqrHPgbWCeonhMmNKfmDsRD4WOuyfS3vRiD5DogJFfdyAd
yXrufCo13Vd//nLTITzDdTaAcZTH6ksAfSzOECdkZw90LsF3GomzqRa0U/JT
3pQuGhFKULE/jpJIMdujp6Fee6NmEeHmeskub6fz3ZbHZHSDPFjoXb2PXmXs
yTOquuk4PK74CML3IrrXC9vEW2kb3NpZUm+1U7eXeAsDBTMMSpqCnYefezLK
fV3w/0FYIhFBvH+othU9LeKiZ9FZWU10m5me0z0ox8MLZ7EiG1h1jZFnlU81
1O/vmuSq3Zt8mTyuBVIQJF1mbzbOJ5QP3Uo2Qlhi/TrryF4FALr45rZwVj+V
MX79IgWiRlEBtYkPY9Wy0UoJVBXb4g9M/oEo3X0l3fRqwK8YhsqP7V/y4sEE
sLTKJcNdSC2fNUQObRPBowST+Os2XX4VXX9XJIa2VVhIzNzR9zHeFUzOb2g+
a3pHQSAym7nr1s8EF4q5xuesvUshBLHU7KDA4VQMFubVHdBvtjVQYJQ0PHrR
Mis0W+jPGnwCKswAZ/qMEPszW6woZmkPFB/2Jcby5XRJpWrX9fD0YuUcw7QR
w9l2Ox0UDOidTH8YPvkLolZYyXTE0S2NaKHZbU4HbtUJoiacDY0HMp5AzK2O
RV8N40nBLeguFPFg2kXFC3ypWvFVzB9pSbl+7squvd4akzKoCPvfMhtIqK0X
1z1FN598/4Q7Q7uboxyK78ACueV8MWA9SmPj6vmhJSVWga6RivxXSXcJdJhx
H1loZdr9/AT6EkLtnOsDvYpVz4DxhCHPEGvpeamb9QhaPKB4sjx2L1CCxhl1
ucTjWVizIX7+64PCkkP0i6Ay9LY6up8FNIH+kdbdG6aHGnEPI9PUeSKMQWlH
zpY3PUiLZE268MoN6f7w2pxz9p3inyedSQnvIOzJ7qaSuGNTOR+xG78Kj4Jc
TCURYuuUV1wudbaVRj/lqljp3ch7wv5rkmuLsey7BnOG5try1DQ8pUf6sqJX
dI0lyh3Ui+KEk3Rxlsxwdf64ICeuZv1kG0WHMKMvbjXAyR4rkKevVqPzQ+Aw
5zgoLSjpyAouekd19izEkv4P/gDdNE8biKO94kcPCnFPTBquzcnjtL9dqnjv
Ry19Ts5PPbGf0IriJcIXvODG/mSiPc2i41awYshYYXfJVnWOVe5mqfQPW9y7
LNcCU9MxrHZ+T88hAjyRLYwGWXtADyRnDyadj9HA7ifvBs8y0kYsX0q0oiii
HSY4qVgls5fllzRq8KvSjSmgxNFSlEOToCwdxD7sqGKA2t183PMc/A3HtNOX
6xKEato7kxjtMun+Rgv9VDfTQZS4bUcMocw204ikAEonluyUxohu9AVLFXwZ
aDdpEcgkIjucZegfULDupYmuxac+XmYR4bWB5qUwm9gIjmylLXnsLmHvnLw9
eKeAULa4zlVE8l8vBiFF7dwNqxTUscJz9EL6xFD5jouDXdp/j3l+KluqbDBA
TNFI95j7t3S3ztxPQOUMAcfFrypnoRmnIddbGeqOlOdiR163e2IujyhfsUMJ
VolxC6fMt3x1QiwDkMI64QEbiDnEZ1LQiGcRE7QKMNDG+TqM5w5i9OtTUF0H
camrUzadvNRE36k+OR8RKDlLzT9UNAqsA/v2jb+MPtNT4h2r9zELfccu6xP4
BhpbQwZUXrtuH0EWnTrMH4ANEg/dkAl1eLBP3JyBtHPXsRBfZhpeEymaJFt9
wh8Vgp8hwFEdF7YcE3BOkzLW4lDtHpoODcygANC0ZpdxPcOlDV1/qaP5M3D9
8U5TgHQSYV0sUO8YX/5f2bdj1Z8GMAXul1U+/vQ5Op/np7myTT3BHL0hUA1X
aTH6ZrXr4b94ptJ0ofTXejPSlxrPufWD3jwbvc8+CdixK8SdsYWGR6o/Rbk5
rZ4eeQ4iabc3csQ5xLPQg8b2DGi6x1JHJH7+AJ3rHvGY8CchbVBRYcKoVWKk
VZpuxX+Y3sT22t5ZZdoWkfyLQmxo9/QM9ChvUSh1As6Yv/Nz3X9/RiiohZji
zK52N67ZzThNJw3ghjqXXmftVOwOqU1umiBKCLorUqARsMZ0CQPk7OJvBGGy
l8Bgjb9Vou9Mn7cqkzkYbZpyh1TFoEZonSEF2t80kcpn4UYST9TYiWGLy4Op
Q78tvMFiHbkQkSz+5Y4/tlCIhPttA9HYFWlm0mD8DSETXQ1UsVKB4FFPHi7y
tAbX26lAhC3KaO4o4O7lQXZV4P1eTa1MnXlVP3AIwvv5jCJZ1A1kvp0ZFifi
Y62/jRaV5EN0MRJGjSLjjeVeL4oUTUvfFKA8UvYb0cblxje1IdWNCBaAF6sa
ix6vWc+wpBCru5TQz3Lx+WoEIFRYhEd4J+fUSja3rFOf+2Jm1PCC3bkqdt0q
ptg6lDpAj7y97eQGDXKJbziHezYLCLkpYOenTYWfkkRXX7ideR2W/YCEY+/n
DGBgnMlZWsiLkdmA/pGFDcdIxzQ/WX1W523RHThSXCvPvF6rFnfdFhhb/mGF
TIVchR2Olom2Vnyo297tZboXpjj2p4zyD45QgJ6g1TO58SCEj2/jpcUhtnUW
7iPypc6T85PL4t1BDrVK7gOYGZMvu3GR9hNGmUeqbkZ1vpBa04EP0nu2ZfXh
xesck8QVfZB5A73ayvui+SdkMmXkG82kKtE2zU5bulgO1HYcXD1X

`pragma protect end_protected
