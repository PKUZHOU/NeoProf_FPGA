// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
dfDCdRoH+wEqfvKAS+cJ/miMsqJqvQUrfBrGX6uN0sWQ4CftaKADPSIN5DzmmAoz
RkhTHE+LcePYcEB6zarBqV1SbdTplHnuYpfcDkiDgOgsR83ysM4MpekXXaafWWad
ZQpzhMw78v7zq4MFVhPk14OaQV0aWrX+Bc7RZf1tD3nxkNqRT1ny+g==
//pragma protect end_key_block
//pragma protect digest_block
gCwUCeLr+7g5dZZXI0QM247RSsI=
//pragma protect end_digest_block
//pragma protect data_block
Bgz4VUCmdWAT2tKMywR8s9REABUDCSxJPWpBgcV+rlEVIKBVzfCbJ7ru6y/KZEJq
DuAHjitz5FM9Xp+GCA81Pzod7qe0MAupdJu6qUjeKMYZNBH2vETXMr3Nwj1bWbWN
8nvfyzlFwYXxIbe/4x4kYEB/T1PZDNL5SHCXEYksChGmYTpmqcPubvbbp3Y9DBwy
CGwXfv3u+gcp2LUvGQoKjnLG+Ktk+7PU+oW4hiajsZAXtRQDZxxAcX9qUQlcCQhn
s87syvynU/iAsSIeu6fdvZ+0yMVXBOnvoKsO50yqaABoMBKYpuJMNXUEueQvMWc5
fdxTmyH1UIX+zVfk9XXPrhijo/InSDljjLBph3tbi+XaV/BJqlRrmDChlojZ7fFF
o9h3J+SL9fQMqUT3Fbj7o88WIOrxo/G24cPRs2hoaetLNHkbzP/KS+wBMmxKZQY3
KzflQazk7bO+qagmjoolWMsmgonUfvxSXeug34XO+E/YloIFxXAghdzr3ltSntEu
lwRRLxfZrpa+up1IbjNPhgVaZWC8Me4yopwPq3vJFK2gzl1/XUVoHJb5CIkcIPHk
Nzj88qHSxhqMO/9WtBOJDDqKU872EmspNZH0LQrRpvC0yIkhVFVAyADXytzD2Fag
IgP/BMIWW0YWphDu9i3cCtGuC2ftUEiizvLJTt5zo97itX2j2GDRYZi/FMNkM8To
VDJOGDgOb3eNekZf3K1gi6ajB7qD8Vx7eVcOqKr9IBTUG443npRvuqxrfbrTcYbK
RIVeZ0WPsNsDLGVUW//+wOPy4Vigm0nC3uVviWjgltCuyjLq4qF8ZOktqZwTZzMu
+zPYXCQ2SlRIfL4prxjPIV9Y9yycjcFXgPSWeFN/s3V5vKKlytFMtHdqJJOdi4pa
IbrXr06DrRHNDo6YDqq1FHA1HnxDHByZcsRQAAM1Q73GGPLz4B398kTdOaZiVPjU
9HrMk8UZbduwVS2PWPhBBM/RbOgIwE72kK/8+5k4Iab1cVTlja1Q7OrTxcL58x7a
fZAsVb6DHb7e2/YaYL1YxNoXrin6clX6E5/v+ql8YxlzwqCeH8E+bKuR1xvpYJmL
DKO70ZXWO8/YLqVcIyhMNYhd6vmVy/zuaT+8U4qhe64rE3qYDXE4ukLBXZR26p0I
h88cEg4GMy7zHHIPXY2NAplti3IHN2kDCbN2kXIsZ1+wdMHuJl51tRTxAybXGxm2
MfkH9FJYzlGYl+jmr8lodpC2mkdW0tb3u9FaJ5nYlAnTE4w/zLCsYynwbJx/m4XV
AKJGk6p0v/yVRhQeoyBwzw/GqGOWUThqwSRl92PiuyVYmClpoFmxoCSQGZUhkOjd
FboTZPdgMdCk/Bn2JAHMwSzymQO1ed+m3YXu89c81lXJznEJFrWKZxwqFUFpe8UD
3cie1+x2HQaZ4yIUnQZfyAQeVBe85ZZJwdJzFS3MYyrq4kj+/UnYw1abv/fO9dAr
/rCQmL1Alq/soSS3gqRySgb3LL1jgi711joacSc4ZLR+0fb+fvNzBDEaBCWRPQsQ
RdldDD7ta3Vx88ASXYH01aPyb3mx6VQlovmL5OVzV9FJaGfb4YmtAwHNyVGVgouo
O1DtZcak6ihtHrFN4KEtxE150AYqQa+y9Zb7jG/eKVWfdLR73wwSuLTULMGRa3Jz
a5qwKmxXVqyY2IXOKGQzGT/8ml7dpd0ra44qv9Itsf5MhJqRDRTXNEPJId5rgjzv
Uxt7YnXigjv4J4g3NlUWYN/CfLnyEmqCCmR4qTL4olqBimruCQSPMlQAIE47Oiux
NGzIea9PgyG2gLJ1hpkH+pn9MH96ScOXtRlicImSsRBxLTQybebCf516V8DXL8cH
AKQc1V9mwywJKoxEruC4qMJcEghIOF+8Q5/f8x15tn+YbfULggCoAJ/kHYyhtfjC
xDlNqQQ8T/1Y8Ew/Q6iweXpu7/mEgOeyOZY07C3EzNeAMRmhepsmMYyl1m7cwHYp
F3Vkd6e2ZokWf4ii24lvJsJ8twR7CzdRrPFbWbbRif1HfszdXMbFqBRACA0NDYQG
BlY2X5iA5VIGYWdgDh2YQGzJO+Iz8Nla6h1wKjeXS3l7lpN9upqWc0O/jFvBhKit
+hr4zpe17vza4k6WbGGqdmFhnvNTWKWGO9kAr9FzYxWaisK/LBcaXn/ud7ODPMsH
RB+2JHc0tRzqux5fjNfG3Sx09466pteAaMQ9LE/P58bM+KqAMkWLO1g+qjNzeYw9
dqLEB51YrdON/YDnubHbQddw/PiS5ZvOauRoZv8cuRHl+SRcRQbugPG7EIhIzp2U
A2ZZjqDgB+CDVu/KT1vCUiKdNl7r0N/YGdXGcr8yF0GKuwpVkLM27LmqvedNIwb7
LUpil8Pk+wvHboJLCDRUvLE6AFiaikm/XwSeZoTfn7nv/SH/DYB1y2HGM1xcbLlf
Xo9stpQJCbvzPvtnw3ijV74ver6KKmMFtNm/a9hlU+jSd/C+v23uLn6FuVsNY7RS
QYAI2IuvFZ4lygTrZybAN+odjwd3CBbRUYQHW30URRU1x5IvGLJMO6tKQNtZ8WwW
i4DT7LW+QzFRUxqWMOHNrOa95NparQ04I5FSonjQolYg15R6QbncZDmqzpjj2Hia
naCdVznW5SvySHTZiKxBWRJAwWXGA5YDwcQVPIHlj7Y32IkKWy6WM22Hu0zauRsA
2OSHARCzDnrmIpQ8UOZgpuKXXM7gx5784rzgxHF6YPmYFR3Vfcr2ydVKB659kOep
zqVuAowZE/xlqmOzYDfFon+P6ogj4JYIiBoLW0yVMAP2pWPbf9s5kLyTqitO7mv9
92PQD8qeaiSyXG0Ahf5ehXyX4V1pRk7ju2KzDZm2ADQPBQRmyUwmlZBWa2UeQb8+
4VUqtU2ThgJID70eXqlFsPcXU02NPfHroF4sZGI8iEQCWKo7JQ5my/mbgwtePd8w
TZ2I6ohGbnYxrzPBeR5wXoVXogBr7H2i2NIMO0o6GYsfO5kxLmDyUQ3q53mniDoD
PDFhOcRHz55VTuJsPD2THe4jII4UtF0JyI/vNiKm4y1VEb8i4J2xbXboUzEjRVDu
IcDZMOIKmDq5+y23U84dKVx3+c9TUWf3oUqN/W717cN7Haa3deemVQF++3iGoMPU
UwKQIfqnHcj+bF8V9/JPQs58XrZVsaTmdvIiSmLpw2OA5IvFo1QyOkXAyqDtXRxB
7Ay6IZ/irA7NqQL9L6ne2J66+ztLQCkFulCjxoafJk+4Q+4ZQ61zuwaLRfnZrY07
DPDI/h3gHKZhKBMQIYCNXwi+qm4Vn/3N1sXT62ggkkMct9ixivgjuZ0fOZFOzEQL
JD7wEW8iI0CRLH6UE+h1klSZwsXSqLmj5VfYaS+zfMlNza5AgzMdnn6d8A5esyvj
sFmGBCyLLmqyY2H8uG2C404bXHjJIx/QmQlBGafw/HyGYrMAWox+dTFYehp0tVDP
F/SSvu9pn5l/zIeugQOh6UqUa0xpW+Cy6VyjJEcTGQ2aOjedE1BRLXtswy1YK7Er
Vi/GseDinUJ+zH5vIVnDvKM4CfOTBxZA5rZZHae76PAT5ygfzexjvJApYM51zRlz
2m350izalnGN8sCrixh0K+2inwiXt5AYlTEI395qjcMpFqtte1qZ6RcMbdeZ/ass
BxHQREBuFPRLpllY00dELn9oPRepOhQ6MnZcdnltudqkg7ubyPsBKIiHHKhuaooN
d73XMnUojmEAxaIJ0K9nLFepFr1gWYPazuWW1ZGtuSADUcu7pn2ILLeXvIkdgV4a
d6q1Jh+3gPCRba3c5gqHvU8xEgoppwO2jDHre98mfFOiy1/BbAT10OdDKTtTDReo
XrYXVuMXOa1RbFweHNLamVXy9eG1NeGl8gR1pT6Ki0ix6r0dncuv/mTyntywcIbJ
StJIvSKYdDvM6hX02fWOP5+8MvJybxLrYH7k3hbAGfqIBz8eNObYgsfTUtEI/3n8
mY180XyLBhim6MR+qTJhg0kmA5yN8Sx4VwxV4OtLsz3ESZpFFhpnI94S1WkAP97D
aeznVB/DOGbhiIDN3QFoiuDJa0IOTliNB+qNLOwOb5tOl45TRtikku5ZQ3VS3lwr
kEzl23rHZH3f9T4K5Cu4NYpCC3T7gREyjAR18nSE79pRQwYrF86jLtidMgSK61dt
C+CXAly2QBgG1pDBQm/YNULuIR22fYe+7oL95qLhuXyfoJkk4AyxrdguA/K+5WKN
bDtc7/CerQLJc8Uxo5MxGGVrd8KFJD/SbXYHtxI+/guezNrZl5vQcAebfUuIW2xe
FviZcVlLIXxCtH+4XnjEyuijCA8q9QRGIfVJkZVZvnqNBTugVf9kiG4ttFzyKLXs
WaMZKc9qORnfjRH06ljSrp+Ds3JF6nAYssFg805FBKgbDQScAP4ZYbDZcUqm6Qgi
SMXq/LxbZUmc6t6LRV9V4vRmyT5DwUu/c0qPiEQQr7T7/KbbO6DGyQjb4AeizBrF
1NOb/bbfs+V+0nipfQAoE6vMVq2zbfDquYBSPprpmV3YYbxDxW+mlNOV8IEhEd0k
yyexVKunAbD+05xpy6DoLSvUSMYbb4aV8xX1GBkGSx7HH7Z7UAviG/NUQigczK+I
kuVdBzoj60Qg3cEKDyOSzWqSGleNqRi1adj6JMEGRk7XWc19Pk1ntoBRXp5tvsE5
OhF/q3quQimxIl52jhYybnoTLhNZfz5NN3IS/vS4D+7nfL5k6TnnLf38j8u7hCZk
DfWAOqClx9Bz7X5ls22sRzBuRJH4V6fxGnDUxYGEmhhyf7WEO84T1QH6Zfkoe73w
v3Fgtda4YtXadiIP+imo5ISVVS6kn/e8L7o3fqRWKOLZrwUpVXuzl0S17htA5bPd
dsh3W2l0srv3RrClsnBA9b+SnLLwVSu07pqlqKfVCe/Zo+PP6dX4Bx6eszMCq/dh
9VbAUtsccTygYka594OgkZf5oGncjkKLERZF+eI84EUiV6+3HxIkJudH//5qeQ5s
tdn8DL5SlpNa2auYaw9OVJvhjwQcjTLmHxpWHgL7kUEafGXNQlX9qtR0IonQnAR4
xmDsc+wO67nU0LVzXxuFXk3BG5LYe0ubIVKqEOPI7ikyuH3hePbU5JTVYZhCVpET
1Aql6kdgc3COIs8SFOAwx1ocviGb/NiqFWF+KymVrn+eUtv1N8IZqf0yeRJ9R/zi
h2xlmyO886t/PnKhIQnKKxqVjr3W44eYM0aopKRaEpVyHDhVkO950O8RvYEVkz+o
7V+pQQgsNk94SWJ7ybDP4dsUqi0x3GfpKERBaTVsAlu5el0qDge6djqbPjvY+39g
KXy9W+khVOj5I7UzEjJ9l/X2y1wOYbgTjcZhd68/niuk6nM9OjrG8DUXAYM1c9s+
Kjsz1pYvp/p61aQWllbDBhGQK9PM3sCwXqBwqcveXwM1s/3xBZUh2DMvB1S1qLiM
GQf0Q4Pxmab9mqnHSKg5/QjveRlePhGo4fXH0qyc6aVf9JxUUSAdHLKJa9nIUuT6
DGmgkoat6GxDcUu4Hw5DCzqp06JKuIuhi1F/DwAJazj7v609lggL6tqwh894OJ2i
h97E0hLSmKB25DslMHHhCrsTauUNPP+y+r1ERcahd97x/6u1aHYcLTxeCM21edJ7
QxfMLD0jSgiMPRkdSmIsoX+RnPzrWw5XO3lQmj8EVliQHfksyI6cBlc0/q24R45P
Z9Jwdq3brd8SYtOsr1Czw8470beLHJX6IHCqmtgM1Kslt+fa6VE0Ob+ePolz2arG
nHqApRJtEA7BRtOYAL4eqoZjIc3yfPgOwj6/996I1EhcU3G5IK6Z0Yx8J01gRmp+
GrnD5TcPQUSLnCB1SVAYjTmzZEqlY6iHz7XBIwqcI28R98Wijzt76FkiDiSspFvL
aoAwdko9TnK2jHWjtNJx13SMu0Uj8sqd96lS0dqwmI1ySbPk5yQmRgi/YcmwTKcb
qS5MYkUWoKrE2XjI5HXC9I9BVfblJZCvRhB8q52b7a4K2b2M4vvJGbXmp4rFhDnz
DRrt1UAcOj77E/wDbpuusyL+BypaUwWGNBsQW+NxOqy0E+ixN+5nc0R0g4FlmhGA
kNzuEdVXcHknxpdI5OCb6YmtFSjUPKyMxxIef//ykzM5H0wt7589OJQWQEo+JQXJ
TIEN0rIdO5qUGrUIGUjoRCVeKcECJ8ed9cAQShhlhypO0/vbFovrZmhKLtk6u0Zf
6x7x22u9sOHN+T11gazolBnuxbl9tMl7gWVns3/4eBESE3g81sAFpz4NEFGi30wb
Abub/sSf4xnrYU0GqLEK5E3k9i/JoNWRdjUPLOp9iO6Vq6uOvCrzLbY5vjmPLxPI
PNUryz6gk/Y/uP6Wxv9nK03D3xDZ9OiP0VVYCbLdgI97L5rBMEAKStws1z4NWt1o
dFusDJWz4vUnczTnPrRg2XdktwY7JJBMYKdeWb+r4p2emEH9wA91cnkGZHqRZ6qd
KORx9bBTfkQ4w9dFWRO2poA8j6kNF/c4i8BnOP8WYhpFJlwdOCXe5cS7jgzsUli4
DBTnZDOlr3pqtZkn98m942AkLZVcDT3XcuNtwOwbIrUKEt98mCA8ZHSphc7ZmOY9
kqI0hJXOMjbZSrq/Lr8FFDYGkjCkoWUn5YwbmRRHscayDstyTitztWPClAaOq8Aq
ArjxVHxD24b/qak6asMw5C8r+nuwbWsiVe1hXUk4q1wk6oq9k5dcqg5PvROnUPPY
va9/kCWJeSgnOac/CREzrdnAxie6VLA4w50sjYbXfMcBGmG70Mne4P5yNsluChpT
O796q5SjE9H9bCGKq/fnFWUy3tW8iTN7fbDldQBW8/vdsMDaEM0sozy5DC2fS9OA
b4L+EBXZwpir90F+GkPNV6CWwBRFUiEWs+Fxl+/Oil6znPz3Ec7e/L3bOt+bSx7K
+OQrQ5vF3Xy9kKIsm28aK+Wi11w19AskV+ybNspo7xNrnVvx3IhRvbgkgGHVokw7
3v873nZSg89hTxrTqRdYNPKm+owmITDhHbEeO7cY8Tr/xEy1yVYhQQ2Pam9Rnf0D
ZwMFd24XZRrRW9sCddVMK0Ac16eI9BqKHgzV0jHFxUUl1F/HN/oIuuvbjk+Jy850
osRwgS12NL2HKXoftrkN6KAjQ7sqEAyBCi+mBNKo8CTq1zxO3bJYcMPMesgkwnRK
nAMjw3shclYPOaq2/c8MFRPGr2IX8XWTRWcKFb8tJQon+f0m85nfjsNKp08I0uA8
aDgr4sUWZT7ZUtp5IgEDBkZcenutfQj77WQBsrI2iXDu4U72J3h3tCFrN8rfXLt/
i+B9jalsEJbFM4YaS67LP/DVv02e0ftl5Y7eSBQfwgquDqmRJVC3u4VAE98E1IlO
GEbMJyqjaxM3eHS4tAHTKBsTsCNKYxLlkOiOrg/rdJHSffKAyxCSXBeoHTnXVWWy
QdDgkPUEIn8Y+EN2ygWHyG1qgWJJ3P5+COjhZ6yC9OViEpzf2xJMfKuJIhTG6SPh
5gRMOaZHb11OgoXayvyHT6ixSt/vPRtswYX70yMgVvIm6k8Y8XeSBXbQBK7kQHj9
gd4WoNgMTGiTs4v6WS1gORz0vgUSFJBAb/3QT580vOxAHRcCYqCgbEOxZiSTnE0a
ngyPkdtSpLg6pQJC47HhjStojH/PyOR9/I31qzUBaI+eXlcEn/HFM8jIyaOi15Hv
+00jnQqAxmdkpXdTSyyGYk/Mts46MLUWbhX6j7MHLBvT9IWieddczqhrSedj8wjT
GBHG+mDhRROZwDD8rH0WZP27j2P9hL7lwikd8uE7E9O+PZ9/qq5joXlDiVc5CYYG
+wqtvJJWgP6x/DlqD8h3b0K0ofgaaKenKVLw8OuvIsQW81g7hf06jO8Jvn889mUl
ZSW/C+vBBEvo1dnEvVl3J3pe5EPRyPVFPTcX0zLzM4vENvhh7peLV0VMZIzOWMkv
UY3U/2RqZuzSZRMNwtbNh3p0KE9HM4WUgindcCRVkH4WMTmtsDQCp/1ggKGIDSf7
mKSDZbytXxwEnXkw0EXJPJElB6A76X8iktzOKvxYGneY6pYXBRKJqv94rol8haZr
mrmrck828KzDjs3/Srg+dScKtRt7EWcNyDzTw8m37LHk6wRkbKV3N4x86p0BKJdM
/LyBgFfyTPrqWCu+f73wpvxul5U9gp5L/QuhHgZqvwbztrJiorGDiygekP/0I46x
HTPocbhTw2sJd/m2kRsNnnEk8Vw9cr1kSl/whXHYrIGci78PxbyBgxSac1p7llA8
nwODJ879jkXeUEG86wpfMSD/3XD0X/2n9Da3ZQ3vuAx4lZmuc45xI/y0KVhuh6f2
f4a8a3s4v33GIXUXGNQv52+t6+zUmB9y/vDVQYdtVKOJ9r/RDQa3ZF2GQLRjhnR5
YxQ0q6mFYZtN6ha6Bs9rEb9gqRiaUhe+8vbFk+ABbmENz2Ft+C6MXhnmVAzyZwSG
HxA0bhvNS+qo3boQzEs5gOZxZSyId3LK35v4EN4EjGdepo+RGbA/ue/ko5jAF+iX
l3XxvFQEUY6VdpnM0nXL/MxPvsDcrh4HgOW/niksPfS8yot2sN0J7dGpquxM7V6W
VkGdf5QRo7RM0GqgY5ZpA7OZvzMdSMfBNHUD1envdgifDI4q6QIdECzv4S2lQSel
zyLaN8NOVotlmY7s4HmtJy0W/Dirx+bRnZO42sKn49OHY++JhJjeIT05uZ/gBssj
0moUFCjnIwFkwGlr5Q7jtNkexFfx0VY5CPi05CBIi1SiiHAGMb8MDVjwZI8LLHDz
AqejupnNkVccMSWUnsxI6rCHZmuutfZE3RJ2LH0VClKt2g/okZXwk3T+HnArrjn6
jG/RCJLZ8Qu56u/y6IkaF+13CSO/WOXsxMmGrOFKdsWZkesOu+XMy5jbgAc6TzwL
KX66btuGMr1C+nnNBfp101ObghAwN9N9U8LCUwtg4oMY/P42dnhE7p7iy0RF+XrS
vlRR8CHhEHZzr1cIGvu54XomLBGw/DF3qnRLGxJE2731BT06cZezR/8c3dFb153x
yw62EgGjQ2F07GcwCw0yywHZ5uq2TeeXIqH+qxWxetIensOVF9E8ibnyZsiaH8tD
DkSNn9LRq7PNsxjFa+sMHyfdIpbNoR+RaTi6dS8YdiVufdf7f2Kbc9kqI0DSJaz+
hG8vVICPZ849R7tAIpY9C558LdstJGkJoVusidGnqWMWs60r4xYrfulpH2jocefV
aclwzQtck8IQGRnbpmnplKIYR2kI8SH0vvCGNPGiWi+ER03jkNSWBLEy359h19r5
YEDw/LQn+3489o2tJtnPlKgoL6B7HDJYpZogwC+hUvY6FlgjG4XVfg3aRCRsSI2O
WyXzCmL2rWYDooBDKgcO2uonckxIfOFoiyTsHq7a0nzr2pR8Riu7YABndCdQslSZ
bhXQc3uGexfqqxJp5unE5ekKjx41cDEs2fmFU10N3xut8Dehe1RahI0XTcKJPk+L
AGML3HHbPC91dtP+9Epm+d11fyG12X7Lwg++g84Y+0Y1jzVcNkqO7R2yGVI338Jx
0zBkDGyQ2xZmHacafQcshQCtYGnGNgIo9t/suPVlGVbrsUmdMDnDkFTdJLqO7dYJ
aM3Vg0ZoiSA++U86o5/9Qxbf4AWeWAUTkQSx+CJuKoQKNTKnbsrnWkSSjfy4SdZv
RyANLOPgtLgo6yKytfOJ1AnmqdIUi/o7opEtSBifuw38y8ial31JeadtqHEPWMCw
Zyz+qnjthSEgxtVtNWai29UuNOgoPBq8ILg3JL+TVSI/NzaX1sxwy7D6fLb067hB
wvh1bLnJwNgynOX1b0/93BWHqmHfJqCkjcg5sOHC4tgx1n9HTupNykJ9/ciNdRAo
/xszxqmKYV8Zj//FEGdh7gdcT5QirnoN/a+/GeYGC0MwX+Mv6TqzTdz24w3RzFR5
ZktoTjLC4+WxNVwXFxKdTrz/AVp2XrR438JNfr10NsGVzeLZiFM9fBKaYqFLCvMR
PHX1L7U35DID6smQD5ZprtFK52z/zCKQXtvxGndJ+hIMCR4i6+tWSyJ/ZLtYaTmI
NP0z5+4GISFi6p28P0g1Lkm/47Vxrxq4i2p1ebjCX1ydsZxew5qkuAuJK6owavAf
0bxNRhcUNT3p9rahds0d+iRWSBoshJ4ybVDlFui90U3qB7KFplGTpqpJl2E13uEP
rSPgbIMTrFpkCoZQBiW85huwTQyIP/IkXdIWcMGEuCfx9LGybT/Q8EzOP+pP45Pq
MKRymC4znPncOtK/BQyyEmrW1+7AMts/yQZ1S0tsfoW342/uL33lSpQtUMAlpS8U
nkf9XkwX4h1UmspgJthfCFP7pw4Lwp6VLRfRJy2rRm1Jur9i9VAogpT7G/kmywxH
FCr0vaBi0QhBt5a9hclqNa0L9TJxjZZ19sC9vD10gK449QzTyVLO19X5W1BHKLp6
04w1RhwRfryuqVsqtEqjHJiQbJwsCPuxqohbDUbDALztXFZyKvMJAbdBVRmu8BqF
KHSx8MwhOy9xzcxy2uCh5YSiK6CUWEulwE2Rd5hgPa7wJPyQye3UDZVsbOWA8npX
ng+7bY1xEIplCjKk7WHHiIltwuiz2Gk0pLZyGnH3FVmsNMbrAFs6UOuKzRHQIDDD
1dpXnek2A3tIiLvH+d/hMOIo2jlyPOnkyhMN8zRo4ykT1CTkuRt+l9+wMD32Ye4G
EsFbMIzz/3CDuj/eQasOHRio947PQQB6rQhurgaCzg0fvbN0X9eBW/3+yM0ar0kr
hW/K6MWPI+FEXd1Vabh+lQHB/rCE+0rh4kYH3I2NAE1k9IWu9ZI6axR+dcDzXnzf
DeRBvKcE6Vwq3iBmTRnUhtVclVbd/PXi2NTY+AstnPzBW9Y1Xf7SaG94zDQiKazF
9Yy/9WSkdPoA48mf/GHa5fU1hS3Skmw9LUO8v0Q2+LKI/xNy/fJ4TRz7ZANuFz02
smcFXUnTDfGzsOhFIBbwbzybP/qkqfvXtav1LC7ZMyBmCqiVQcKH1t0gyC5gPsU4
fy5nzgdZbMa2domfSDeBQLAonG+6naB45zOIcrHXUhKI1e84etbpc2pbYT0CSAVa
mBNGN7VoigwjabTtYQ91CxxGsvOriIX2lf6j231f3XNXaO2iiR7/wkDmF/f3/RFr
JYEEtprqQy6/ERMyAxH4ZzQsHiJ5UdsTrv86Z3J2gfy7ab3lT+lfXR03IUmFfVQL
QVHeMrv4POsGyf72GHmPHVhcIeJUhz7S80MuFmP11MQ1fRRNOrx4IVIKzqPwKHj2
BLVPoDMp7u9bs6Vyp1GnouvJbucoWrBScTPV9prys9XOFBRP1WcaCJoxZbyG5VOz
2uOPpomOnoYw8ixuV/rrwH8DYu+0rldZFFF51/H3Mv7IEA7Qu1a/pGg+tFitxSwe
RCWm09bCniqxtF2wXHuGwZPZ4caNEMrpDu5s6UQi8xlZfMp2HA8s1QMehpuPJlqv
25Y6HsXMC7f7BK3qQdZrgx+xWKOyiwCfvcgke5yuYhIZdVIKEXm9VVjlcvkKOuIL
u+Uw64HACwdoj4laHuxp3VXiQHHAtTIMA+akLcPGxqaV5gVXGtNCiKJppvOdzuPI
TP1fyCgmIbGmNvGF5p2Nw9guzskTAP+PaaC0bf/Y93EM22ZiDwlMt2iHGqtikble
e4YCmpaRr8FKYwEgZZBtooFQpdGw7vD2/ePmgIFQiB4SCkHkttagTsB0nHf0/CKz
H1WMQj/b/iLFACalZ9f+Y7ZlUynF6v5KZmkG8S95KJ0AM+vlBbY08pPSIABQzAFx
xDJJHzqJ+q121aa9VdAkrBCsBDNHGHZzR0tzhDxoJyvdon1qtuA+7NkZWFP/Ak0S
9JPhII4QxexoumjGsDhrlRiSVbGmtFt99uVRY/sFu4TQ/AMlfvi7UwNiABTOeUtx
pc23xvA35yYPJ8UzehmAXLfTIotE73B4lcGtmTZR/dRJLzjgTRRAVu37Ft5+qkRw
kmXQ8iw6VmeejH5U4N/qig==
//pragma protect end_data_block
//pragma protect digest_block
Y+sW76ndF9IO+y9sxAf7XX7cOvg=
//pragma protect end_digest_block
//pragma protect end_protected
