// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qgo4/GWjCHPBizEKdOKUo1nEEyxdlhQtcB+NRrAduYDTNj29+ux+Wm+P/SjUP1OvvtUdhyRDfw/Z
/eJI8p9NjF2IEF1M3hWeVH4hOuDRu8FRtFT9BmDaeJMegG+uqhw9mNgpZPeoV77KfsxDvLzL3mFe
yaznF17Soa79kPF2ilHi8hdew1tGbb4t3O8BGV9XQBhzSFV7xDlGJyQPO3Fe3r/I6EozkWnfRS9s
hIIuu1ZQvdS3zjAhiXyM+XAka5CMm1RjFRTHZFQSMDuR6YH3+OVk6bbKPje15661FVBVvNOK6kzM
r1WhYhVF9vBhwCMb7ZAKhEM9JrwxBakS+zkWow==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10656)
wpdIJnnjM5sRVvfInVDlwh4lmip9dMgZk3FGgnXAFAm3sKLQyNxH1cGWtxcs5UB562G1FflFasty
N8WeBSDRclxeRtrwOhl0mWFm4QCOrSRyKV0WpSch1zaNex+hy99oREFhOfszPAQ4cuUiYIcTtDYt
t8X3ubcgongEwI42AVwIkwfkrtfhK8PcdMsJ0fb9spcHmKH2jBbki98Hx0GbBuc30Oc/NdKImstE
CQlkGy/ZFxgqV9HZiRAPopyrOwJubBCGmCdOrurEIuylHcsjNyxVtbxKmxpKMQeTqgBUgKnP9HrZ
S+urmBg86EyD8Qw7u3LXxtrNCY6vF7MRP90LUQLkXUzG4RtkKPTuoOL7xvMh3vrlDx2xSs2ZCMKS
KEHeTObO1CNBmqh/arIByQoy2k68e6dZKz9+/tj4iXDdAC+NvR4MRAlEsR09TeWUyZ3wP6wcj74L
7GR7tRfjQf1EneV4uKMb8OYktoFrkgaZUg8e7Wks6C+rXqGCEi9kz5Xw/m8zM5OLvahwke00/R2d
e/6Y8l38FLECsKqzZLKKwGQ35MGQtWXA02UCY+p7pQlCTn0n5fYpaxfC/c/qkWC5EHRIPnmZtsBq
JjcjCkwRhhevoYSAEC8PadT382zrdU7NwIMI2JP/te1M/DySiAbNAr6AtJOeb/dKArcSmZH9xQUk
KvvcMpbKyztERxF6LmNeBwMo2zUKM5GUgz9F7EPg1PTuIP1s9rY603qEdD70ErqrSoDfo4rmfqaM
2EGsxE1gq/PaQ3F4Nfp4WwTL9MmUFDy158gMc4B2bGXd9eVhEN154wfFaVAs6PykfwgKoA6qQL6r
mwVVniCvGmt9Vdz2NTEKEDvIr9KS65MjxciBybJFIo9+sVo03t7GSLsuLhUYkrpjf1O9/P814M0w
8djZYzf5KQePjd+bXDoy58QNu7Mxfre57FV5V45lRDixVNJrS9PEqWwSySif7bjTipWdD8F0LSrL
AOWOaM4hZOcAvFI+9Na93/FUmSBdEN6aO6xnaNXxwwgc5Z6feYOFuxqKJGZrgtTBZw7kjohz08pf
Ob9sN6Vs2vFfl4dx6XrxvgxrtoKDyTIXpW32C8O8kHiCDr1RG2YVsDUyw5guOni89QwopN/teLP+
ZxGSIMpcdSiC+IumL0AU3EwFj2My6WYXWnFU0CUwzVad64CqcuS3Z/u9uzs17SXhEPPYYOWPB9QX
bcjEFWsw6LLL8F+llhAQx1N7Isy3pkn5lYynP5DWHP5JqfCrp4cpWb/Wseozshax1rOOD7oYCAGY
PPj56uqZoCWmmigK6IQ8zBNoizvLGMDA9tWkB9VfjwOYvk6A6YlUpDfq86KO1DGxTfalc39d9Ze/
qsjVuA+Mp9okqqeIBqDwVhrR6BXiXSREAyujBUZWcFW4kWL03o9DJEPJ+zUN9L3zFk/b4PP7m0/R
B2vqYF8N2QpTtxp8vB8H77pLvGqhATFhd7Ea9WvqUbDf2ZZBgA5Fwc2LUABO/wMnWHERic14FbVJ
DBvXd2xgYMDfjUZ26MkkixI1AbaZHaS1Ih1Z5Rxx7NxA2zOePiOE8+rdqDdydRcSPUf2VWQ2HEuk
dP/ZxPdNIDvVxPt1kepI+o8jMCl9koBjhTd+5YdGNfboiQEvjv9MPF283CT3sXFz3JBaq53laMQf
kgShfrfNOCmZQ5hXNmLyFveWdp9PoSaSl1DKUR3p4/leKcu1BsHD7qIAOg++pS+4OyfopIDrybFm
q1uNCyfjns3wBFWETpZ/xCWYxMpg8U9FM9n/UbXlbAouoGgP5UZRT6iw4AU4FR9xhWfIhLpl/oTG
2xNCHiMdhYciB8vfQD9qPDyIBJPiVS7y2pEZq73f9jNlz4g++0Mi8xYmUXmgnzBgLhBN7HV4zW0E
eE2IbZBGCBTvVEEVgC0pDhwnMkHsgyNs4U8DqGLDJQoLGW1KBz4QTld56VpjtkosT3czc6xGkukq
faxyH7Miyj9740qz0DlIAVHxfFk9FnDySbJX4XGNjCWfm8XdyLwvtaann26e+HotVGQ30DI4u2ir
t+TWqunb0VUuyx4W525tZRRPWjAhtikSOwX2jvAwlugWL+UJHgVSCkEImMoMH6h+R9b/0fnGlOIn
+JTzrF9W7B5AA8n1XWNvrlTMcZ/AQdzoHkn3+vpDOhcNeYj0OEtDbil/M+IfLsbIKfeJzqL+BEoZ
Dk950IEb+FTV4JG8hw4tLvgAoSkNpWHAD+3CY4C91SXTtARIKzrVi3H7l6kH0GiijzBhVvY+/lFX
svlzAnedN8VY/lBmn9ra3bVQ0QX6rCjX97YYh3v7k6ZSpGb+SIYdelQZybdT8HZXcsyDNU8syMQT
e4zsytPX2ucC1BpKzzbp2kOoug6FXind9rPy8d7avGAo9SwpA5CLjiroGaebma+SXu/YG7BpUDZK
jgYGh1x1cQvlE5YUzDg+dNQqfV7QtC44k5LaCZcNHLDpkUD9WOnvpDBC70T1HnjvFLVX9LeT6vHt
thA9T+ZdnY0pjLP/1B+6QAI912RPJc8EM4ZyDtk0wN+27hzrhZInHXaZakKamjjMOGMu0iVQaF23
lQo1NHSAcL8J5dM65yaszEq3nlryEypNYyNlr7YajGx1yg70LE647mipGBV5uAYetIpHrmbb4BSG
hYHGmQrbbi442Rrd9ZdhoRyhaI9yPTm68L/QkYvsKa7H1XdRGYjSeZLF/VVFrz7VMB3/YMXAZiEh
ybpAUkc9uitCqMfS17BGIhSaiBR7G9dXgGKCZ4VyWBjf0Fkqmcd8q7KBGhwCEZX5VnY3ZpQfALM6
RiZBWeIL/MigLakZRxVmgFFxDsJ31Frq0AunM7lw0gwewcbvFvy2DtSvUG8eDO5EHQEU+62ghQl7
O02JNd1aN/Uc/du+Q0yRE4dB/6kdB1xOV6LHrlbn8N0RbXCbZ+274DeGWDj35MjmDDcgoqpy7hwX
DncRmvHaB28zB7tuvDOCruwSVXBtZA+UJlVaxGmzo/v4xMz/QDwXoeWo+B/aHPrjNkNvtqOxIe9T
wycoz2q0l5X0uBANQ7W6juhpLUQxtpao+9VePWE1JUMc4Ys1PrigrGe7RBiDfh1aqyoP1EmyUo4l
jng7r05c8edNMJCf7pUVudJlk3n2++pilMXdt/IpLsfgBIHFhesylfSFHdNz5IJVOUoKfk3sfmVx
tt5x96s08QG+ouiotMUo185czG6CO8KasVpVE1HBSVCdAm7MJqgIB6GT3UFSMsTO3vl+JRH4FWyk
j5TzS5MEe0iSzfrfL2v6myTCI4BiOa7vFCPbBMlscOra49gxqygEKM3hRucCZ3LjvLk0tb6Ormxl
mqPc0kgBA16gFrCyocGO/qRJsxCP8GDnq6+c2VZZ2FXMOiRfum3Po4GxLbD70waHOKAef1UiOqU1
e6KtEWb7WQrdNaZ3IcTvPm6J+FLt1Nh3hIcQOENBHV48FsOZQ75sdCXgzOPDarffp9FwHO/B7cLs
qbdZJUCGy6gXzkiiLL/x3oFLDLWl08t1b2WOI6FYqEkAwL30AQ89hrgkbVp8pSDpF+hhBr46nWvv
j+te7KVuv42rCkiM3Xg+JNMFyk7vp7Yi2aImymbtDqVSSiHurSbnW7ZIGzmJE73/euTtbSM1G7Zq
h4QlR48W/opJRw/Xa7XbS/D2ns9gcIkCinRqQ7p50FsQf7wSYnA596xN9GvkjlqX5L/kTC9FMKL5
wSaIh4eY3LcLigfJvluXBylBtiUwHdIu1GK3nXevhroM8Sl2pofBqSnUqD29/fXHhnVkR3H6GqwG
BlvZbOPrCvfwEySm3GrG9uM1N2eewzCa/bHvjY8/rcdmniJZW8YYO6OgbFoCB6ou9Vrb+gyLZdXu
/9CrufWfleQ4pUCKiDxwHngsTHW8zf47Kbczd0EGmJ0syhPuohXIUjoq/GkJFLIq4TSeZB4GGXkq
u4jFIG0mI01t0ACRDYVvORhBzlOc6bys6pWm8Y3347Bbh/ZZ0a16nMYGyZnvTeczpwf+JDSvouCH
DPng/u1Wim4gQGMSmFDtfDyTVRR3BeJEatec+c1iwXkSsN/iCiNYczcLUn4s/1RUwgBIJe6GMKcu
WmyT0Q5dPwcep2YuHE6LNMTVLBls1h9ijCz+pbJw9EMOhTNAbyZ8XtroSLbfYYyZIQsAMLRqdNvo
ZF0w79ai8AfRBvf5MUu9OtiOYQ6cPZut5jlDB3v4J/Nzhwc9kpuPZf5QMS78DXhfVfVPM2OLuMC5
xFtCEnLC5YJIRUZo/7sCH8+qNnXYJwwtOzEk8niTOthRgEoflDmLUWjsGRV0NzvVCKdXJMfWbDgM
/tYVzhWSyDHDeXhcRi7WuLe65nMGgoyKwEAiirYubQRpZV5JNwyYQvbs100NOIOtTrz4i1f9ej0u
N2ZyVqI5t1/oe8gjQ+Z6wn3NbvIa/A5gYLJH4cQWv8FfrIXfPu0wq7K5ll0pVvQDDW2/qZejbAuX
EeysOPrgtGIw7UfCLilt5XobyjZ8CTtVcRiEf1m+NzDUwAUVe0TDwiDjvTiLt0L/JZF7d+JG1s4G
y8l8OlnCJ783iqcGPQ70zO/KXI25XX+RfIWHqU6kcJjU9dIaV2mp1t1g1l823nG7V44bh038mwEA
khkoBajmbAbSwGSbkFDt/7KR4GsRFMgYEqCZ95xgURMWm6fe9CJ3cG809llkOkLehuW+8HFZZtGZ
CYjW4fWBjA2+WNQ6y7XRkQ9hqDcY7i7I3u5/yrgRicGi98BRrfA5DSB3QxS8ObyOhmN1UzErLZ0x
zYFEZnUD7vyZU/NCxYbZn4hv0F3rgvXRS6UHJzvpL54RKQZNbt/NZGUffF1/iRycX2PTPMI4GHJp
Hh8nEVuWU02qrGDk2H6ovcds9f8WdfY+rzWuGXmW2U3Cw2ozmsHCke+LnQY4Sg8ldXDYj1VlXLEy
kIY4MNKnJ8dL8e+kJp+81ARZAjtH4c2V6kpB++/1TpJP2h+OnuSOWUa3A4ZkAJxOOwdyDWRAsze6
Fm03uM+Y7yGO0H2AFF5XPxElXuGUijqzZDylH1fu5VvMjgxFha22vs0JMMu+0f1KKyavpJ+P0DjY
f4WFQoa6cZPEbzBC5NlGQe4dltidDLHCCn3yq4/iggF9XqybqEPCZM7s+nR8c3YLhAX3UpeG3Q4h
+8IKX3NPQR+ydNUecOM2wcfXBw0JqDmCYcqPYzdJG6YpWM2Wr8SH1IAA0HAKsAL5U1g7gH8g42AJ
yCMx7FWIrX82XgQegyz6lD2l7oBqcddsUEaCv8sRE+89JaGCLU1914HrLuDtMCMOdx++XLJKJ40i
d4RzWCax1POZC/7wBrnT0cKHv2sCv3jrXsbE9Uce9vynEh0ftoxMo4nouLrpVtm5u8e9/lbv/pHi
IJgaLUWpsnw36imaRrO97aW5hAbIgZaKWZQrHCDusDoq4W+DrmysOyGXyf0RsOmmZXBemVNtVssG
Dc3YcjmtizWCagAiA1/+vzK7ZfvgUm3pQq9bBCy0SR/PeafReiU6ZjhFSTqIfrnjuCdm1kGxaY1a
kBN492ERNwyHvROi0l4mCysq3dKJSnL+4W2g+MQObGfi6nk+ULkBIA27BJ+DHw6G5Kmfz3A39rU6
nmMsnkfTC6e+dq23btF+vH0CRUdQumtdSSSVPFbc4nOlvoTPnGJp2hG9g7OwsScOm226Q6ZpS+n9
duzMyXhLbmwtI4HwoTEDYyo7jAN1zdlLaz5Bzvt04W9fSoDbO+7Gm/7aW5v4fXnPTb3nb7t7KuAa
6IHWuaEH3qNbxQBpQocpk6NbF5JWz6jJBT2QC9I7FyPbrFT5w8cQNIiGUJwylzxLeBXe7EIrJTC4
GcZarejUUTOCcDPZerWPL8xSug/TOqWRby9k5USAtyCwpJVvtL6bd7ARFijkzKzQVoUxKLGMr47K
qsj028c/YEXZmjgnVf5oPle9m5ErniA/GTRYat+8z2KLIRLPyVQuSW9BSjPB6fJw0d5PoMx7ATxb
ihN/MPPao/yLYPSBi8wKzDiv48DQCqE9bkKuVZGYJy6+a4z4ZIlrEJmYDb6oPNKoESmPpIFY1a9E
CK+e7r2p/xoWfMpU1Mhjtlazv8EI1SZ+E1oRG0u/D0Km8mYcxsEIHQZ3gWsrhIAwYwnm6ApwN5fR
SGTH2UBqxFPzzOpRAfr7Q0hh2sMIkYfkEQPCt8sS9VCWMKwaWJXwj6pwpK+3aCAmE6fYUxFLnV16
Np2ZoUkXHzpsTLof83NcbYRvUWRitds5Rg7aP+VGOfxmyPEzIempMC8y07RhNqi5Bav9SNje8x8a
+8t2SLKUs13AY/Sga+qmMx4TGyPalOFYo52kBrZcTqBh2r+i+JKSxdyz3PpEeRyJmHdn1FBXJRxW
EwB2fNt0d6XGL/iK9ObIRRyejH2GC9Xcg95tzJf54J5UyjmwouLnf9Qo0CaxXJgLpVr5jFwWmt0G
baxInXWojVv3qGLro+GcoaOxtL3BZhvkuxMf2rvSgxhgcdJ0lvm8v2XRXYUw24fc4RjOIL8ULm4J
8PDW7xITaz4kOxiivr1Gm1iHIXXnBMdGwJgNotXMDPT1yDhDYAAEZ03ZOFXi3Tz3tJ/7M5P+YsuF
3A9CEdOIdF9d7xn1gBgRlyAnqDzXdcmg4IWpJxjQpNKt3XxaAT8HpH005OVyt3CAIsL4bhU0h5XS
okv8XY8AR9T+cFU0ML8ali+taNkugadsfxOLB3H84iJHYpiNCNP5bniPzEtrn/W6kVlHIvCIaWtO
KJIi+hK8M2dtFO+0FJE3NWFkVXIPly6q8/BkoPn63LL9NpreCWheuoB7Z1Htwx2iqfddEgMtFEVj
HlRePqb/eLFGDVpyNdykWmBjDC0Ue9JVuO4Ush/cuiMoKpGaM2ern1wduoZ+YigQYj9Ts2BOjy7I
54fXMrkR/S5QtrsLP+rY8uFC1RaAqiSzPZ/qInx++S44RHPf1/HAKkpUQVt0kKMUyNrGP8/qdTf7
vRcakZs+sNU013dNYWMMprWIxMpGYrp3mBUuIMQMUFsaHnnF2HczUmw7nDeX7Q8VfxJXni09y9jk
o3hF+9PTRdybBMVTLrTbtp9wKWyG/LRMajzI0/t3AGg4nLwLZR+VpJmyzlzn6rNztUzF6yuRdQ9Y
mxEAkRook4UT3wykCdEUrhUvKZlSyC4fXkxDaPKOEeO4Nz0x4HuNe7reZNRrwqTJ69UCqCJB/Tos
TF3JwsDWavbjxtmonNk/J0DarRYnfVFwZEmc38BaXxhhYS6UHaB0MozhDl2OdY6iLiRWDStWOUs0
pP5Kgc7jUInRYC6zXiVD7pLfJx4vmp6HSLoFMDGLuFqTKGTCNpBkb9DxC+2OhEiOe+MDG+s/G/xx
YthtEdIKTJhXlHPvjbP582twSI5fVdDM0L4VpOLsv6Ws4NEWQRUOB9BuodCo8HF/GCK0rpNuZ9wG
DjGdVEDZ4ptWDGWtHw9L4f+cXN4H7cLjo6agLY91Av4Rjvw2P9BRaTm66k4MEMo94A3XK+AwN7ot
Dl8IA4yOJ9aVKF7XQLW3jAXR2yCMSNTxQ7k0HQbJPhrhgWRovszk49Ezk06J8CC3z122Npt3IiMK
0nKwqHPoF8f+neMS+6h1h0+nj/5rI+rNPuWo0xFMLycZ6QkPt8N/169tvHkGmitaszXO8oUdMvLX
fw64ct72Ekix8xQ8HQDzSI16aaf1XoP5YEMgrvaWAtb0jmfBJgkYKEKDI0qZ+m0BXOd2chRl896A
Cw1rF4zsGdd+97Ciryzt7Vi1kBpmk6AFIwKCitxrQdU6p9iCN7GL9PtitJAXjrR3xla8lQlVF2zO
hu7K+w9Ujzid1dhrdgpb8Cpzv20wxSdh7ZulzMJMN3qSvvUs/g5VT/+yYaLqE1wPfh8NBCKnq5hy
veqAbIVrsaBrFZhCsoP6j0pjf8ZQUAcNS2CnWOlG37WD/ZKoAogDuEKo9KEyUSE6mmTw8ZNUonhw
kLGuVRSRhLjNpwyGcBh13bHT8rQXta6PBM64z/OMTbw/uWzZkTcyQRKs4pddCqzFUMQVFogHA3fI
ctvcwqaFzjypO8lkTnpAM6vyy/dhjHRxLzpS0t1dNfVCxx7Tihck5vEwc58zsewVXeVGuGGn0PCs
pn2Bqb5ZNuk2OmyE+l3joTTBj5gUQ6bwbOton8M2m2UDbu9s9nw5oG2rMO/2n/jfLotymGRENmNJ
iQAMSc6bNupsnkLrNsm2MGy6AZwsAFDO4CSBGUR50zMXQzI27FTp1CPJIxkYO/j9ml15ahkXytg7
6YCKDwTd8eUgH5BMuiJgA3du9QPbQzuut6OuTFYB3GScHTWOlT2SloxzmFvqJk1+kMSdUbzIUkaa
EfQqW5PM2VPIr5NG8ytd8Yt6yLbQQR3/GabO6kOsTiUrulnIQ91mlsfWnobIVqIh2bz78aPz2UU2
/2KiHs0cDcvfqF0o6EOF0muXKxqQhUGMmyGfzyhKiJ4v9O6l6IwTZgPtV7MJLMRxm4saE7aU4R9o
SRL90v7fitq3FF9TnV0mwmzoaAc2++WVpA1KA4O0NraJ+39Bj98Zfo2/cEQ+aJ3/j7cPrpb+LaPy
kkQH19pnPFMRm5v+NBR/uDbKvMavdLyhUU8THz2+Pq76EQd3TDVal1IwME/wGdjYh5e3YcHOwtyJ
c7kbEsGev7+/UbysjgxZ3LahrEqq03L8tjGlXntCrBL1hJIhgsUp203ifrFISKttjMyZVVeR6wB7
CpOJdVoztUW1Ns//cVP+VMTJVkzW7ZznteYAXYC+XxQhepFTl5TsxxqckB/7S5XR7cEoi41w+NTY
EKu7NjfzlYtu+H6BM2V9899Pvbe2EUFGR+XA3DvbbcOhpJsuiSwJx6vACuHcLvv2FUBXD/non9h5
ycgQec4OE7yerJ/RbLcmiQaGairq4hI6MfM4lUzXH8X7FVhBsU4O6baWSfxm012luvxS/CY0kAXs
g+wlG87UfElEccLXs/dT0HDZYCrVuJxla8cs/PSmgOxtLRea2++w41PCOFoU7lAmC/b5MRouti1M
KTlkMLTwHCnFPCezL5Tj0CxzubhfKBSGmADxePWvsM1G33vF3BYCw4OcpWe+FJX5KS6dq5K86LAw
typWs2eCHwFgS7XvPFZWaiyW2NK3VxzuMuET+Fpdt+wq4EZMUakCbK69OzTZetGDMA+vEGwmXdWy
PiYLVU12o3BqnS7fI/X2NERk8p1/3pKzQBXmO2fAi/rFS84TbDpn42tbriZTEraOJDQIsY/Wd0p/
FnawLU6QxOKz/P3Jw5NSkMerkd74QrIJxGAsdADCvIJoCMFjGKT01FdvQZRnvY+O+l6FlLgXNDGS
fYmMrpqQlJmNj5EqyGb4geNy0y8ltEPwmRY0933Vlec8RApWvTRr78oIISe3N0eKFbDKSFbusB3Z
9mHq4W3xEEHLi+Op8tqU3f9MXSfguTbdyYYZPjS1ZKaLoTZfM6WslmXeww4D6F2SLdTNcr1TICTk
3GYWBHG/KuXFCJ5k1CC5RtzTPexbzvLEE2yXi2A03TzN7vsWjNPQA3Tifcj9sOl0O80b/XhdkfDO
dlVn5uAAZXLEtDGGQeU3S8EIwLTYgQG6oUlHcDCQDvmtciUt98TlejDeHqnJoZ4EGD/wgDhW3hOk
6twHQtV/vjfbn9SyF781TleYEahpIfo0gAjgW+NNo9U/0EjBin1WxTzsa3PUI4lopkFI/necSW2b
4uwq5xNKJ4DFhU5eFDbjDFRdbxQ2rmhD+fYXEfo8GEUgsu5R07SZRGy5P5lvaWrXtsfEQJgP+1Br
U7vvPWouhYuKMFaCMzcSS0jR779fdm5JJYEeHfW5FphhjdunAvDx4nisae5EIYa94BdR7QrcWpR9
tQxvOWSN20xrBQQy7wfKY5tJDMPD6E1z73g9gDYGh/tyLdNqyjaQsNlPotKb2DR8OEM73oD+fWPs
Y9mZEs7Dzf63rY3rVc+NAoN89kD2GG3I0j8SfFrp8hkUbPiJjqwAGQ2RXYl+tKIrxmDP1jtzG0VG
tvdX/gsCkQPeGLm9Hys1lUWBywDVCFcmiy5LaRdizlo5E2bnztpBTQ/wFmTp0CtHrxHXLjxnRxcD
3a+hDW/ztdojW6PHkbkLUQHJnLK+uuAmF2pmhr9SskGb/WGpq/PQcbXwTjQ91ra/bcmphl1olFcb
iVEuUXrgoMgOTGBqOaLjVOiIErcESj6HdfLb+vTO5u51X99nOE+rHrCxRaPBlg+85DgxvbMDUKrw
W8FN7GJtqM3c+3qEZ5iDrEC59YyC/zr9pcKuxtRFRgM3jwJHfbUX7Hv9qVw0MhbIugmCTRqE6oPW
ATg3kCkRIVixtTkHDoGFOGYHIkbPWHUJQ8ITKkvMkEiryLsdruyPEZanCJQs9JToOO+JQwHpe9xD
8XbRkLzJuDp7UAMteCHCTe8F4fUK1el3bEf3iovevsZu3uWaxMcuSVaguvCLcPeg0eigoufwF0q+
4VQnZkiGpP3K9qS4oyu501hesrdVQ8zOiR1MeDIM7Ntosvg1zGvL/pvj9Dzf43BC/DOl2m41ggmP
x+j6NOkQPL4RxhIGPvLZ5vJl+o80mVFkcwUCuCKKnOlaaHTjLJkeVgV4HcR5zsfeFvgR6GePBxPF
MQiRbD4wYsumw4y700DA9/5O2voOe+vJMVgC8ddwfd9rnE9XO3dWDzzcuqM7fYuA1HbY9+7R6Qkm
PJ46Y7zKxY70Yv6MXOzgK9kL7GJmjTwvUkPbibcMpZxI+TYRpowM4x0P+9BCfdouw2CQJ59J1ISv
6bmSFvKqwHikzwQS4qyAq0PQbO7RbVk5pTE6O9V6+jS/skqHhuigXhHxNXmqq9sWeyyRE6xX1rPr
R1RRtfOqn2+GmC0tN9aV8Gh4ULBdpmQ1iMigorD3KnHLa+b1HpOUYYc1fSFEK3M9XqRnSov6gKcr
ADIJxAy1M3UQi4tp+haCVH+l9OKhD3aK3Q4BQTH2rmB6o5QJj6WhcQksElAkPMTUM3YT99h5g8v2
0B0+GKoiaF23etqkzUNwHQa2UtjuOOTxdPYgeJ+oADN/iyqMl1H9WKA6fPXhAJ/VMMe2TkgfBmub
1CHMcWcUB6X6XO1va56cVtqdxLLF9gALovzGb0LnT9TB9rXr8SoAEiCiIC6/P+KPV/xwZQkxfzlm
DC+Pqyvo5aQD0TQ/9PccKMVmKL9Vw27hCXFkFV0pwmNWDqrOo08V/XRlQ3eNiZ2srYWvS7QS8esB
9cbU0O42fkn4Bnm630XqL6spITqC+AxkE94kOoDEZ295SkrdHDAr5X9Ab8CEHY7n3H5hoX68uXBJ
/iCsCa9tDhD7rawEl1UyPgYtdEB1GlCXR8cTv9GdCw/zd3lWvfz0ddKwUaa1MUNDjQtZCOOxpqhO
Fvm8x6FAJC5ohhWtJtCLRoSY49m7x9cMXoDj4QoLEEEwpeqY/YpjkOoZLuaKvg9f/r45wHj9OvE4
4a9ofMVLSYXckTCle5UlEZpyfJ9BYhUsINQ5y7QtFSb/1VR7SzYA00F9hvDzVHqszAetqjlg55ly
OsKM02X8Af3BSsytTjkKzHYlB9Cb9nUaxkuRR5RbmfXqNT3pP0bZiAzIVNymQ2gCyTePtalvyjcY
qjUeF6a/oWuaf7lYWg1/vitZS02x2xYW2WRzmH8oC0sh75DdEFgaHKdicWuhlUFWG7uOioaUOAaI
SIL8uLfcHipb0zKjb9Pq13X4c+hFbH9NVdk0FzfS+P8b4O5+/sEJiVsQJ6h74wVBP4lr0IavRMKl
JnUIDbhFwO1nprzMLCN64muIvRvXV1wN+FYPP3w2rEeG2QPHryAclOZzWZFD9jQ8FALRBGMXqhwA
WKIy5QzUXrZZAHNBwaPfC/3Kwo9tpzEhAw8ACkyz6WMXQDZohwNtpVgmQz7g8CVkpB51mtboQgbL
IUx/jSi8BKq+OGPINKmTSc7Jpw6V2q4TYBfcohHW9h7dOPeFCkA16pdtZgwOe45YQAk2OjZscZxR
+MHSDL8vIY2r9WoOywHqjR7opx9zsM58QDX3LPC2FRXG9WqzDBQ11nUbVF54EQ/WapNE6itG4Z3P
1aTXDygqLxZtz/xO5WiBnlw1eoQDAW0TBAO75/ujCHf7um0Djs+mMr3iuODZZ4OkKbie6UKnek6t
X/IpgEyjZdwspHjrrm2ho21DYUi/I6LGUaH9uj+wr0c2OdcdAu4KaVQ4fVwHSpY4WbMGixAbpvhs
1uuiMorUl9bl0V2ywCz0OqtZZhENL6wUJe+Qv31jQw/4iAe/+lA2Aw4n6RB5K7CJFC1yBO+vmVfq
0OAJRY1jScIc/810VhGyhTlJaW0hwamNm+xIBfei79ePNvsgz7AZ3KOEtL76AIs3qDXDXG0Eq43z
I123NUslSE11hSvqHEwDwXO/zmw07en+M5VvhSxZJCgsCmHoth9WBR7T9ZxPCUdPZ0dVG5NAqXxS
/pv7sI1Cq4a7ED0GmJIO8TucFEESVy+3zyVpoI8/qBjynP0uZx3aNfNNWgS+T/GrGCO1xcWiu2sz
vcVXQQBDevQwzGkt/j3kLMOvlZt3MFSaiFs3K7ZXAUjkZA4MiRKuymDi9ymXUs9zmcYncWDu1Ppx
vJNk+4Nh40pFBeG/sF46EnLPPUVS281YeVYzdzB0/WKXf9DjlOddp/dz4Uwypfu1iWGD9xytKwPN
+hinLBTFJA9SYXoJBQLz6SxKvUR2rRgOtOAnqcSwiH5/3WolGlqtJFm4dPYcOCqiFPGiQKN66R2f
VWTIRFyWEMEvRxc7FnFGejiwkR74mrRDUtUGPs8iOjJWigeI72UdH/5GBoCu/FYSJM5cCAPF7rbS
pUptglawXdt9puYUIUu2AAXjLRgS48IOF4V1puj9Aqwuct/jOLCcm+IpG9BBHbtrvml1d485yqL8
79UlWsO3BkQoHX+13zB+nqL/bSwWmj0NPWipfcSUzjulf0sYPOl/WF45DkaBt5Au1JI+ZRnuTcc2
goWY+9C9b/MuRc2pgUD1XlAgRVeYfqMN5iVqaeSTYc8+/lAT2ZguVhkMB/V571vH3r8+KaNjiS1N
kKdoqT6+B1yBqabMTZhLSd+YMbu3l/jKfg251oD9Kh0vMKgmJu2YRw7SLSRxLMDM1vZYoZ71zapm
LTgqj8NzmJob+WFPl7Gzd+y/BPmtWVNeyIo8LppYLaTfTyqxnzudZV0sydMb/iosQHkHd8iffq+7
98xi3Vku10dIxhdyi7iKjSIgj6c/qVsFbT+Ya4dP6XVT4UQWfl4M7DEGEPq1DznD01sVMPSDIHD+
PLN5+5CGnwJV2acCtKMu33Fx7WNFkSq1sr6qLnr+qCAt3oBXjhYaOOu55kVCetjj1cgQM9ZWKZgR
YZfTv0gMDBRvRUWZrjg/Fv+oi76G+4VxbsRnMCknfqtxmmBxG1eDtEgsZKi3+csvCtsXtKyeXuE6
8QzYQXMyOB4how0y1MjCJvqjvd15kSF4FmtmT91ko9za3lPIixw5UNAY/T3chznuM5NfsdrURtuX
BVx2Y0BV7S4h5INJ39n2Jmpow2pbsZdeVqV7irEPG+DTaY5sv8RQQ8iv1ru8mrxQyy2pXh/kdoKT
5s64KMRL3DTDK27P53aNDtGZ1fhcvWXQ8TBbQviSm+NdL9GyAOltXvWLIhKMF0gXz4HL8792STBG
GBOSTbxbCG+LVLj63uzSqv2qnvy6GRL+8rcO6ouqWlbL3IGyWvlT26CRWVZ8cFT1YtVhPVpVMZxZ
Zpw803tfCou5FFYjJty0d61N652bCS7C0jMapZlnJvSopdJVI63k1UKGwOHE5XrTLCi6F0XXBfyY
XUHOwh+pseDx+PIKCBw042dAC7wKSQ+sPJS5p9nltv1BxXci3jhUcKobhXbkJH3A15e1m12LVKij
sLFOnItzg2uMI6t2lK6veGsanNL2N5jWmaHJhdOdSiazPixcf988dS6Gj9bmBxp7x7/7zS8OFx32
fAkvoKteAw5N5zVwFkLRVOcKNPwFp9fVMyLTHuL/l3j5fWTT5xePzlDpXCBIGBLpta03/fVQHqZc
Jp2He6T/ENPw/Lg1YPxIVpQvvWY+vwrRWluz+Q+awHV15DcfBTxxu5WbQj1o9nJ9vGjY+fYHoq1A
E7+zDHGudiylQnUIiDD4oPnoPCAcEeSsw/f6xLbYgvtXyfsNEjtxU9Arhzp+BKUfWKAsLdAd
`pragma protect end_protected
