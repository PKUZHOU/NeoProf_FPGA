// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uACd0UFBOxTJI/kluKwDI+fsdxR/YUH1VBqYoar/CcC/dRAMTE4aM0+SnyX/
ngMZ7E3eS9sUfADNCfB+T0vm3tcPfLXvYa6vXxEFVGN6Srgar+ge5EmmQlh/
mgVwN6I3sG1bR/tYMqmm2wP8rVHRNcLA3LypbYEJPZ0kYG+1e/yA+ZB8pCTp
5LxA4BzlmYKj4qS7NTXlfVGHnX7Fh4a/pj4FMdnOEPLsH3vpC5SR53CigWYN
FePL2yE3HaXjpIUs9xUqT0cEQkPRdYLyBmCzWSiBL8iOmNZFGALHYklSz3yu
4Xki4m/pGLW60joaP7rJm21uFBj/3kKimMVBunrGEg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EWMGSQCLAtLDbiCRCV0365p8cwfShB1oX2Jn8zkh2bGNfWX9zTxhMaZ7hwkN
4FvdZrV0/GiJUU8TeWIZzJ9Nhbh4tTwoQ+3+vKA137gqks/30nDJGiu589cH
Zjlct8CXY1AtluDYwS9JJE1TlekHMTaBIvBExvvMTAcHIbN0/FdL8L89rUTO
mUqYG3JEbTML3HTlo6s97AW7s213oT5G+D0mSq3vbxKSwKmUMXTnT+2e5v1s
xgMD1IYySAbvMX8ulWJUxDnueL3biMNIT1voK36MNjpmWbKQpVjufSI+dVDs
2isFk3ahnmFXgJpXRhZiOYcnur6XBdw3SMIjD8JQEQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
G37Qn83pL09dHRfaVGsyLeZzCl1Gz5S5rqSA2BhbfU8baeIeEICh5rCLOwSg
FSJ8pXJbzW63B+mZCw6DiP6eAAjeR1urKZDvoWrhCbCicKWyvJ8oySsNjKB/
8excaOXzFxqZVnuQ60ON+yLAuLUpK3z0fqROY+Jxx+kLZAoEb83bCyaV11Z6
GqZ19f/jlsdTOPSJamduQBbg66n9fSQ21+qzWb/SmWllU3WDw3agcYlOcjud
uiviKkMq0p+vf5FTF03bn8hL365rJCye5ze3zmB5L8nRFSiIjnIVcJPvWrLV
xhI3Wn9h0uxA4k3GyiUcLRN7u03QKo6Dp0UPalw9yg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
faDkFUCVWoMbKYd1rcixymHUEEb/LfGakaHDe/ihrjevJ9Pv+wJibz2PLqzC
NaXHLxpXL4kStisis4k3HxL9WGRDAdnPSNgAvv3podd8Yg2EAyOVdxelVWdD
EIXcvbsbpgJcy+EGyiJRDNCIJF6nlpl/V/Oy8GEcMEAGVj9Mvrg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
EUyoNV1Q2UbkTjr2EDz3JiNTfOVrtsmTnOPjdmtTtQs2T+jsy42d9Xn96Ti2
0Zzf0fPQY0ik9Pi6u8ZV4RZb75E2Gk6MBmNv+JhL9Sw2ybbwDp7z608ghrah
dlx2YsI22aMuiTblehEY62uZx/AjAUoKZUZN2p4KpVG4swIGMSdnDk372SJq
/udVDQNHyTyxHpL3intg2Cpuus5rH8gCupzNvI7YdDqiYMMpVgbWHuOwrDj4
zhEnMgOyLrQQLQHUrCeKyQbFOGvlOfR7wc/oU+P/R9q/ceo59TQi2uBd74/4
iBTZXySji+boiDm4ocugUDTqHF8zS9Ctsi0I8kVtajBYfd2+TvvmtbbAHdaJ
3UjYu8FBqBK58vQuNJe7qOqlMcEk54yOEbTIcS+YCCZvuKXaWwZNp/nZyffk
gGZdHRR8Wgu3w+3kWNRK4SJZ5UkJPa+ddPLqGHnuH4HJgjAWI5pdgam29yLP
2eqPLA+r97ktPdUDCemJIiW75JdIFMnA


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qVQ0N6t57upN67OFprSMka+GI++OcGQXC2ph9sqkFMysdikoCexdFIhZ/+3x
EZml6l+bkV/MLy5guChxscrGmVCCBs3hrR5pYnPe9Sj4XFi/rrfrlyXmSSL6
V3Z4hPO7+HtLp1Ky9HF0jnNzB15v4Vb0gPQBHaaVFimmQxNvXRs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ReMwCbSkUSqCxvjhbMSRvCF/XPU4cICoQF4CWzOth10NyiHuyu2ZXTFQ22vp
PW+IEcr0c1HjysUJFTYgDq6dG2Z7uat6kA2c4Jxhkyn/gOlYd1U01wIR0t3w
nXwj5coDBw0Dp9RCroyAHUsr/kDgctlTm6SwW79RZ9eerAPzHWw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 28352)
`pragma protect data_block
wzf5JTRHHFNzKLTwevOMG+0MxrJQsU2NF0S4461SAtaBRbKKYqS7eZEq0paU
0jk186K4hWQtteg2sN+q8kqXObn0HgRoSI+HlKbIX6D82zYmlqFMhiAlQyIs
xdRl/oecpW7YKyAvqsdJdtHH3GceDJBcHQUKQGI5IvjJ3ta8AXNg3nc2V6Mp
giC4JJNtFhqEBxeK8YW+6ngMITfRLkDUdFpZ+Ojd0uIkrhda8Pt2gQASoOkU
EajeYin3CoLbg2i1J/ydgenIwPCYCSxdFl86J914PkmRRD3u29j9jL7Hgd9z
3Vikab8g0GlS9zcKb27GZ9fOeYVX/+CvkiO5LC2PT6wmvlBEM+6/NDHEyvoP
Mc5z2dxclm0GNdRo5xyr4HPwrTR3ZuxleUO5vBqFijut+yup1X8I5ZeQurLD
fpqoJMU7hINNV9OdY0U3x8YnaXAaKrRvqwxSUEY38p5X6QYpMbJ7whWaK4cb
F81ltcVzFXeNZsBrwUmMvOXl1o/FdWSAwLDgljPqUP7XliCm2DBXrP/Yn7UD
aHf0ymIM37ZuDMC6BUOw4S1NEUFhosbvYANaWQ3eoeHWWZrvfRftFz4fpIk2
QsuAnOyFqO/5rwjFhMh4A/dUJnD7beQ86fAQ1rcOSeWhPo0NXJZfDG+EB18m
AKSOaT0s6fqNznhRRsuQUcjrdu28oEuse32Kkb9caxleGk9SbDDGSSsoj6pX
brmmj31trp7gnt/n+VmNbRM/NUeXHyPL8CBV600W9bJaXAagooRh4dkEiO5U
LzYihDRvbKk5jHgaFCWjm+K4EE376kMrWyg5QM+r5IvSu/ZTsXLu0g/eIuT6
f3t5qEIK0iooJEl+udWzPzyIYnlEoEC0eftCVxmRt/022gmvtMAavmPvPEkx
V95MVPDbD5QiUbs+Y28QYafPFfbrqHDlxCiefOeMNmFXMowvoBAvDFsBSG+g
m0cEjdTYlBN2/BRU6CiWCW2boq4dYmc0eArmHsJtlnZrfsi8IcAoNAdbBZkK
DCiFV1IFIaiLrcYX0k8D+RyR4xEFOHQksG5RzIqlhbNBdFvwibAwAB7HhTd4
zIiCGM5han9QSew2kfsyfUJBZQqPULbQ/a8OWLJRpD5Cz2N+kaH+qSzRMQEf
AHvX5VIJfGjhk8Vr9jJnu8OEwk/x0pWO5q03sfgu3a5UThuDGx06mLXbUnoR
Rwz0SGpx/ryTR1/YJu+fPROxycrxmVY/v7FJg8A/MAlAoXFkWIPy7NFsSMdD
1yfTU/FcbueXa4D7uhW2CIYWKcVRirfUAV6A0BWMKmXS9pdYWZx4cz+UWKDM
Nzli6lcFhAmXFQaM+FMTZh4e47tnLa88MXcRi2w8S+3AeYQ6O/tEDd7Vu7ap
yFezthTRJlm0J6rpcRTIA1/agUnog/3uuapi/xZJG5al+OrECe+suftYP4lr
sMPN1CCXzLdA4OzmmU8NC+fN20U4+MnxFgzBOBvYGLJq6wZYcSYmQcTHfK57
fqA9qh8eno2cN18LOSeoKhxuHel+JDzt3XOX0BlAeI9x83ateBy3OGm5Gk3i
zZqoFW+KgziBHw2biCK4UVqpn1cRm/TNm8W4X5N4od3zgvHdO2A4oWD78t6A
gxfKx6f/C0O2O+wbYuRd/X9fDXOduuWFIfgDF1RuA6/vu9vGtD/skfAF8YuV
qQtkpiJ8U0mH9B1MFb3LNc64DoqOY1qK1SdlmaoAZCgM/H0R/2OndKVHFT4W
tZkclnb5DONGJ7IzXLBvF/hqP1hSbvarxAmZu0C+HHSrd69q/WkafGI50zhH
FhMa2gmd7HNSfUrwXb9kkVAzRz9UY1GwIev9YSYXUNFeH6WdiVck5Jf8vPtb
bwsvIdBWOBXRvO4xBuQfjmVQF7NZqWx0Et0d/+qOUzhyRMOsZMNNxWQupFHZ
VO8gjOOeqnjxdTPPTKIUJVa1KdJHI9U07JhGooUL0DO8OqK/Nqmg8D+JZ/CS
Wi2+J4zXRDplriEdQysl6AelUXsL+JOjFCnJzrbGDe4wloSQmdhXaGL7G/sb
5sPmEvqAOkUD3pdwFgcLBAtMbm/Tyq62bwL57wFmi12gAkvp5E/OSk7nDd/q
ioqkPH21HcPYqsS05BmTFJ4e6BFPz/yXUYzfB4ce9q+KR43ApI72ql57/U8k
Wtgts0EQurRkMJMYYTIeBhB2f1CFGz4VLSWkj8++1+F/eve1dzgClG163RDA
ttxR6+3gPQAWhSS1P8HL5gfDQxF961WZGX808zf69dAYzHxv5aFtpxWyXJps
z0yFQsY5n59pUfHervuI7IIK7j0HJAmz1rkVpcLPr8b4Ystwp69M9kViPW/G
1qqi1PDCDnn5NkxCQbiAy9glKdH4PqPpI+d0AJa/JWWRiqsRdSSgf1tVzAB7
rgW3eCcx2BHI+47RuobkliTfZlviEkwyJvscctrUQ2A6kWjEowj2h2GLSAvU
dMdGCq8oD1QjswjRk5nbem46nlNz3SPrFhBUD/C9adTESpZqFSN6IFulBain
c8ghvidDl2nhk+GDCs0eSdV+j3FURmT1v1EsVLJ7D5+5bN4lfmTDLAAx8BCR
/Q38w9pA8jAmsGYqkaPfISuIsljlsvnqyWhBOkY9srsEaxv8GuripPDkvaYC
ZCObMP1tCQoRW5CsMDRSdxnWTcwcSwqBnkiZivQilQVCWXrGWXOnhz+F0ZD1
FoA8/qRh3dV4gw3uVjF1SwwAHbosqzyqkVEhdtkz+PQOzHCqrpM0Gq71e34V
N27uCDxvPB2VHNKFr35+wgj0t/A/e5qc74+exaEeuQJfsmRf5ZxsMxIOfuJ0
Cl6KajPpm1Mk84rmcGRiddfOI5jPOna8E7F/Qa0Ig5zRXu/LNwPgL2kQG8vR
EdBkW/ueXPwpLMnqQU6krc8CpZKnecT2M7DOL5tLUs3iSUa/37QOotF7AbTB
RuqZ16ilaRpVbvpKMsqDUDYcaf7uP/AyAiQDMItO+NY6x51ROgIUcx+uf4BJ
TN7JnsGIYPuayMxTtsWyOCqwUzir1LHVUoCKuTZd6RI3KsUSCXvBWkBUJudD
zZuRW1JfF5NxdEpz6L+jo8XNEWRJAhi/UXRJVZqrgEdNAKCDupnyIeNskyoU
HSFaaVDL9TfG1fcLk5QSxKVNSnG+2WhwRYK/heu5vDPbZIAyeV3NxX/dEnZc
jEUWLqj2UcOvIFssiLEh9CmhXATsXhGHs6RpDP12sx78aVpQljMDMc4Y2Jne
FulqqoLeqeAod0s41VYjaTsbw7iUYQU4wdwOuef3bnRG0uHPWqz/w15hXAX7
XxCqAdU/MBvBCMoBu4pO61qOJBmeS/NemdyOmH8R+4xsTpMwtpIq3sTgObXZ
M5Mjz4Ai/pBIXOXvjBjaZUGieYyWY/jmwK9Kg6qhGsopyYxm4Zr4fqBaZSgr
utPacKx6Y264oKg4Hi+q/d11SaQEo3ZdMxy6rPIbO4QGaMmnjmc3yIC4onB3
rkVdB1sb7Qbr0zjjbuJW/a+VqjvKX48R53k9QgUcK85Z1JxIUFZr+0PrwfOU
G1hSlwwNJUxbgfRumHBlBmWxb9opRe+9pfRuHX7U5z6Ph7nTMeZ15oHJjjX/
7Tz6HnwqkpRzilS5cgdeSJI+CvB1CGsBsj+kIvwmoimZ8tw7+EV9ulmV9PZ+
ZWDw9o7DYHkOoqfflMGbQsU/5OT8ngXM32Lazxr3jAcHphzBZj/qNv4SDxRw
YuPmq9aq7rOqQamAoiN0dGI8f3KY2CBDQE/rlWYP0TRO74Vlrw7P5zPoX6QF
t1oKKKHgUNHWgXxI+E0AA5rdC+J8HbFQTSW3+QOiPLB54J2GwT/xo+ZLhDpw
NqNIDu9kKrQZ/FQwKc1bbF7pSG6Pz3QQ3MtV3+sDlP7JyeYDkqTivOQ3zxuX
Qtd3JfOtOp+YR12gHa3MpGXhC3P4lGn5ND2iS7qFl1ycxWWIvMLhmvRdRBu8
jdeS3RdpnPff2zwf6/wbMyNf3y8wTFU2EMJ2Hs3HQmC5OgA59aBCtAjqHR0B
VXNbMdGF21UoDBxTVj4Aj0pru+iogiFa0cHGjS0QSJM+JHKrl+i9TRJMNcBB
tfwm4R2tGyC88KRtZgOC0qiG7ZiLFcZjjvQNSIZPi75FTvrcXY+dnYt+wQXT
cNAcyt8ekOY+wWoMl5kkDmpQho6NKhZEzs5QFgdfIo8tx8D1KxNofnzghr1r
YK8USXO7bz/fBHh9szmEOk7t3zA+WNexXsr+Zom2DjsM+UaAS/2dekSXSCyH
6gbQYZ1QItBdc3QbpDmeY/O043+Drjhg+x9mNqDeomxxs7sh9DuFsDE6Oj7J
d0aPu0GsHJkBbxb0K23LDX32zAct7oW1VLMqrjbBJtacuZdx6TU/riluRMZx
Aioxci2KfuMUc1OqUfzK9OCcti0gIcOjNGd0FZne6mlVuz+lxv88tOLqZIHS
QREspus1M1BZt0U8RsOsPJE/pVs9aUyawvOGQrXEf0+uzaQda0Y05fBV4IYV
upquwg5tx8LKoFjh7UiTD+uEm+VePP2GofIty9ZRoICupAXVicUMtsWmhBob
URXY/Xj8ChrDxJ9QD8MvsEw0JmaIOuAX9iPmuuIHlyT4Vh4WKxxaoNotUdqb
bnHEDNcVppHNlXUo2JDLfadXfDmptNFQtGKTvtdujdJHymbYmTHyvvC0v9uh
C3sutyuamy0aT09MtmK9y415CKaf6kaWTLOgLz45fAWcM646mJn+lH0bQUOa
/MjgM3rxdKRt7CGfqYP7ywwGR0DTFTse+BqELtEHWBOXsX1XcchsaEPpCp2W
GNgY3SICKn1ot+fEDaFY1n/RYt6cV7RMujpnDE2qbY3yX7kOemTAZvsDnzhz
rk1yzhpL0FWahg7Cww/+aAVe+M7MGTVjbrYvXDqKCpffiPrgaXYvZnSuq5ze
fjzQnt3zRPSH4tEQHBfkie1GdkeGglPB96/GKlb4np2ohXSZOJvO3PYDz1RT
oTdapYgty51YYLG6T7ZuB1mGuaErC+XS9B/eddhuOwiCxMpnPwtLWESA20Fl
85+SKoB9FMX+kIrBCT0z92v79ELVIIwS8y2RX+LiNUti/X3TzW0bN/0fxgAt
0Ggua8pVzTRVVrrsR+Lzcj3EO0YQAxyNj0p49NczpMjAAEu+9/0A/3C6S2Lx
k3vgNQIfER5s8Hpma1bwU9omzM3kqzdXf1yV2XsDeibPu7UGr22M3XMLmkqB
OFunt/I2krfHp4g9E2y7sviL6NVmNDxmpMNTTpu2dQe67g0kp5BeeazGuqBH
nNdcOJAlTpXiBpxQAdLM+7l3Am21tiOAqUZcXx4uVilXLUaaSPRReShhZpD1
jy3/p/4B1xxBCBHsmk9fcJBfFAnFF696CGhPGl5jOCHl3DuDwF0m3H1WpM0Q
cxaT0pF/2EGX1Q2kxF2d5bE9ZDPHktlc22EGLeVJvml/oyUSpDr85EOJAkBd
N1dClF2pLv21sZ8zUsWqcNdZ6u0BNwlUMYzcH3KDYExXT2JZz/w6SqKG0rK2
lRsq/BPY6OTpAk6T2iTRuFQVlypvfwXlx+lOmq1D6aHGTCRkpp2oeDlzoGdL
IbjZuCewg84wB+pG3D0Uji/1BShFnvQMR5THYShsHdA4IMlOft8wnJNb2yxx
Gebc+agIuUnO64p9tyPFVptGQmlYZKDgcrPwXzHOVUBk4ctTX1mnpdAUoiGh
Jh2IKIiH6kteQ0hgyiD73VQuYtpYnoczgqfiC5TtC9/lzj0bgnt1vEPTRjWX
8UVOWmCc4vLoxMVnwzGkqqH93hCsOT6CrHbTJ//OMT0a4DO8u6AjYUMMCqyk
gBVBYLVcSgJ447N+xrvzv1UFyltrvq7VAFgsNiaXBwELyAJM/9c8IAdu2JUk
wWwWrvTEv3SA8e0+Jzyfc+H7Lrc/UfisjaLE1hegcCIR76k9dCXX8f5ZLK0c
OAhMeRHL9+oHVTRhp+9CLYLGpGxkwjSHGazC/HBvFMxt/EiGuo1jjer75pud
8DqITgOMZDRhl5baaa3zBiK83cTTYeWTsqvr/UTyuPEBxwMxKUt514Xj1rYF
Zulq46/hzSysi1TeMi64KyYg145OZvkr4nF28hTVvTe3uAPeUHS2Z5pV0qMy
bUqYklu87y4DW464XwrCpcdLheBM+CVDcfYm7kvGcjoyZ6opeYE1f2dx8gEF
+ALMlqqvwux9+oYDPuH3Lq76ZfGQFa9+i9C5auhnQYFOxFvhwq/DYU97bE6Z
W2qnfsrN5uYJPEB/WxzlkMMEpKVoqgbCTK7+Q/kD9r1HFhvplaxy15Heh48o
eMO87yQDnPzVFOeR0py3OUiACgE0wDgxCA1q0vTOa4VQGBhsO0s+JlXynPaF
pcqDagAIZm+XdQF9HmCRYDyh66Nib9PZwxNg0QkbWwAeXiNUul9l2WbuwRwS
vccFBhYINKNh4T3+p3NTj+gWMjwNhgXP4ERFG60mwHRsh2QdabTwYXpmuDxo
2wXFQxvijdwI8R66vkqYjiBLp6V04gYhm6HxZCe0QSb2anCfMYox324ZBomk
DPeSSGHRIYmp1FZvsKRFakWdFb/sq/g4kOwxaoAYnef/RXozXRX4RMdNsRtT
9HLKSvjixJCiUVevE9Hhmt/8gkjtmfHx91LX82V/8OZkP0z00nfP8NHr82D9
xxcT/RuGIkoORZ4Liuql+uN7UFei1RzSNkxQzDpwYB4SQN3hN1UkfQV0Nae6
3E55Ggl26YdnNPnBSvPuOQd0wzCwAHNcm3XWfAiAQaOWXw3ucVptCJ2trQ+9
qewvTah/U6liKYvF4OpdWK9hJNRujbZbyqk8JGDPdNJnTIsgZ1I66uLwZD1W
UrEJrYWnsld02U4FtoWNWs6yev0EYAjOhumBirN1wcqbMEoTQltk5qJ48P15
HYxFSuBEqJxdhpPVyKhvAF6rbExGjlrclO27wu3KEsZwdE1cl9Fyhf15HrWg
ygfeKcn+W1NTABY9WMl+5MdK35bTwz6OImCvI0lMaTZZEzckUsVckFNu9axj
RKkQnmQea3o5nW6nWNyF1hcO0PNK+GwIzf3B1URepYrMAeqRGFzL/g8eKWWG
wRgHiFm+Q7gkcDrPtQIR5+APnZc2xJboJXmMoA8lfj2bkxwpsz8YFDCHVatn
WMKFYN3mz7lJ7C4Pj+tP7r3q7x2zVDmmPYoOnin9wxrRWnqcnpKHR/LZo0XY
aqMFo70FCWxiewx9trgfnp+4zuc9/PRE0WrxrPp85LVWnHUXBBtCUvkmtBNR
ok4CqEQ+W6s+BO7IU6R2ip8Wa0IO6vbS/aO5xX6CPH/UcwY7dte8cQW54RLS
+bvgQYHR2Bt1M3PbG/NK4h3+7pVh35959SIj5oiuTTRP9CH6jqRCrJVRzpge
EoZE/PvYPaPgUCnyFHVcFnJuDoFmdTdRmBigZPkgZyOndQem7zDtx0P8FJwW
NMzvPJYo1/jdFFY2W+JmJxh/7+jZLPC4ctw/PxQzZRAauZFYhRqKtG+vfDxo
ZGLKZkszgdOO0cxo5c+mfZStP2VeG2FpQW64Of3ysatvBapJP1TAHw47gwRj
zsgWEWdClJQFgW/DEV4dXaAppX8+s2Hij2Zy5z32E5d6f5KFVrMop1HfpB/J
C4nKBy6jKXj7IXBOBEe4+X9Ys/K6lEJ1I1O9HB2U9Bgmlnkgbv61TA9e1IxF
t90pgzkO4Z6i7kUpxg/BcvO2iC29xmM7OYCuNQ9xKTos0k8HYaOSUcmoZ4gw
PPwJgCttJdFDekLssX/AcJsxp3gvZJTI9zN6ADGK15LnTz9OLO17q7tCl/U5
rrThynaDLUhSSn4f6e8UKks7tBosU/rnwl8NF4o1fqbeMAI0Vrx7/0crBMfz
gzM+eR1LoVgZHoNepNJqaDqPG2AwBylufj/J/3tiPSHKjRrJDwr29ETk3R+Z
oq1rbLe/cd+erERKoZw11OO1Y5uDj4MpliSITh2gJtvoRUXH6IEBbt4LZUY3
BMK+JmqamuFKi7DTFXQnf5HXWRPSOeogFmuSzAoxTysbPEMtrLI2lqudif1G
IOib+AuM4A/65ttcN4UKtg6cc2uGAM5nWwXCPSojIdShFbFwF24if4EQBKhd
fTPcU30uzPoxiV9TvTpdwd6JoSvfIBza+/kQAMPpKqkbOrR9JsVhQLZx5OHs
SuJu0u9ktjjG7BK2uXTp+ScfoKHu9oLtRdmDec9E5RkxpRnRGp7NgNTEA5vi
b4sDVtUjbZhx1Br5/skC2Ni22HVyukm4kObJ/brych/+v4tXry0iiVzZLOpd
jWQ9OsWMjTWVFAuNcDvfeDX1ltC8DX2bZvOww5hLNv8A+M78YMA1tlkRejCE
zBBo2A+Z2D//pqmrY24VhsnHSRmZg4G0290wqyM1xAEygxeBe041xl+rDCZT
JNuUv1f5llRZncnJAf7fbEabqHPjErDC978QAnHon9AWJGr7JdLGEVvBEuGN
ur28mWOHh/SDhLWs/150iQAcYC2AVk3YBa1n1MpZgFyKQ6qLXcKIVZMiAoxW
EzV5QHQ48YXLd8KZbEjpSAst7dbnKcqFsbkuuL6uZNZBryT+EP8AexdnESKm
rDwMZi+FNMm5isL9+DDqC66d7US/GpCykc1mTToQ+ITommVu1WNIa0B3NXZH
XUyXFKr8LHha0zefGQB97N251Qtc3lAwMSwD7GJV+GVmnjD6dOWVAcG/gaK2
BXCSrYZu56N44cPDAUa/SCAGZoIs/rlv9jWKYIegDheFalDTVmDrujIyyl4W
t3xY3sV85netjqEa3NddPVrLjr8dcUt6Ey5GPCGKxx5UbrcdLrhjRWT2uttJ
twIDMvUlq/gXT8En639ClLMjjwx/Qyr51cLSLAaB4lXF+Bqz60YTTvz34+YM
wxf97Lsnn5cH5hdxzbauz2Bw4Qm+wdu1Fyv3FWovgkHAAzEQ8TDgKw2OqUt/
MLnK+cAbnC4oD4qjAtHo+8sqoKGL91ZWN3rQsSJuh2Z5dWxP+01Wci6lkbN/
z4gt7XaC6bmrNkNSC1vgBM7ZfIpcMCqNBYkBMwbm4mDZHjQQYyiLY3Avz63j
FWqvtHhaCZRkxcaYINNIQyX/KLj3rA54NgC4ZdArkZS3Hc5SjkzWck3HetPV
9hfxKnMV4p+/ZOaWnYjl2yGrBL8iRXIyIT65khAfkUQo6wIGM3Ey1UN/Jyan
rHSphq46YBHcz6w+xCgkknBhK9PzbxoQLANYUGlg/sl76yQNImLp0EZvvzd9
wwI1Bd3XTzMFbzitEEtTUlUygTaUep7qFGFB8F/oJxtB0syQUBI0u0aAL85d
kSoBiw9nIk14cdIG1+3BkR836prvYaIq/aaHdU3uUbER/6HTzepQJVKKzCB5
CbxEqXACT1addDdGaFF2jvmwPMpzHbA3rgfXLR5qy9JT+s3IopocFdQXJZb1
jykCcmC5jtZPOak8xkQPzMS7d5FlClQOwkXQiAZPkrNabNKinV9IgAtIIYbQ
7SX/1lLKogUNylUCMrOSSpSMBjXaicwxwDYCjBD3Q8/TyUgEMlfK/evaJOcb
2Yyu/e6Ov1kNyGLstX5kDnERTpifaNyJgHQPKxN0hH7H3jtePnPAufRbdcda
7d8Gm0rylAZL9PCBt8BNL6eiZxK9UcbRVgwRcnYZxzJGpQFH6SwnJi8fKaxH
QGySzT2XyXbhlFfylp0cjcIj9RU1Cg+OLb8EGrerMudzF+1Y3I/1qbBcd5aw
whWf3dLkfdnN/kaaTk+q3mLvpVU1BzduTe+EhED4iHFJQPn4tkd9EkWD/rWA
41FVAfvH+nEKPZkL6hTGZZv+fKiRhklCVKM0cuXWgE67La1gz7wLIc4a0lwe
LwmEh2wlR7oE/zLxW2u3wS5IJtBOXFJ9+ERPdWlezspV2cnkobwxMSWP+Jdq
tTXso630sQLZY9hcrLjmSAgD/89sI5KbGvccJR4doL66Z26Wsy6f5zDrdTfD
+/CoIqVUpbuYZZ3qcdumbzhVk7LYHqPhBQEtMXZO9ifLzNxPrEV3PJZaWPoo
7rkxobfAuOMnDSfe8HRs2MPQB4aSWqQjz5EGiMNfYU00LBfO4mFzbn/N52Si
7Ig0hLS2/V3ehV2zTID7fta95sSVAZYmLfjaDZ1GqVjw3pZ7St2DrFbAbcn1
K2gRH/raQGaOv6xxdBiREEIDuLLWDGc3gfaHalGRNSg+/ZkyjMZpQ0APq3+8
60Ap9vNUPoCD13MPP9ig3LxO3H5p+Ntq8NBfpi7PMJMO2gya4kpaDSek4z+9
AdN1uL6wflOxkEWIObWatnFs/5vRX2nCx29o4ePyaAci3Wwm43+HhjKDo7A9
3hSY/XwvGJJc5Ybojq5V5G2TDvhrQ1nf53B3xvD6a2Y7H5pNKuua8j4B4y+W
kh/Uy4PsqHel4vOg2OktZton8fbxGx1QmTVFWuCoCHTG8+7iZnRyhtcT7A1X
MRRyd4Q5j1jFYDM/Q5oJseXsV7YnO/3RFJ4rO/TAcI5MpETRLJt1pJzpoLyl
TeX3yf3rhz8bTZnQTJo9pGYL4B4fRghgb+b3mmUeUjdH9+ENuYM66uTIKT85
xPw5GJ+8q2/ni52pP4Zrqcq9tOj10AizON4LywZpYQ8ja1zzHpByWzR65U6K
4A9Xpe3HYotmN88o7xyoltWe93wIx2Ew6SdKz2jhlVUjOMB6gG0Axq14L7Sd
oaMhJsV3SapUo1m9Ao0ChWCIYPxYe2yJn2jEAKiEGtzt4YEhnAUopEwy3DE2
R0/6erLDHQzbVE/ceG6pQZ57L5BivNjgq5t/qLeH0xdlGPZFKQ9HanFehXsf
kL+OtDxN4rhN4HuMWXVYUSxJyhV9hANr49uFnj6EmQZ9g0PokawCqBFUY5P9
lgXkEBcc4Htlll013NUAMlWl7QXncI29WLt58K7zAiZQLTcCKznsgymiUn0j
TdcDoc8XKUmFTH3UfpQu2uMzaeUriHP92Yw3kqNwEsINS1jdKnBRxthQZhA5
fqE+NA4lNxJpTqaTbCrlYHYROMnjN7lQXr/zzCztbqBAgZGTcLjfMrE8XWnH
u1zzwdjdu06VFLMNKt2RsAvaXpzNjNHGiNM3V/tAaNuoUeL6gLzbXVPTx56R
QJFdrjT/CJ1RsaYrPJlniZeaRJjY6idObCR1rH1c6f9xN3cvrKaMp47jw78t
kh8cn7gK3JW3tOXlYlWm4/EzWGeaTbdSCJg4RWFaZogzAn9seqYPK290xqZG
5CTzzkQeJnxdaFH/Q4PWR/NHJy725SlmIWuszySogs9TYr9FQgOcGR4t8pYl
78kJV8baSxwVjXdTyOVP9+SM91IFf11f1spykwCgPOVatkylKCBOqlo5KocC
EF7ON5cOxgQLlNavPs7ZACj1pTCEillHwlYh2cqkji0o+mKAt5Y8s0d+gu/u
GMSOZi3Cd0aIx139EEuH1jwzS01rur7ubddth+1jPxVyTlvTpp8zu/SJqeFL
i0xiDStVjQxwp691qNmGBDp2E8LD17aypmAn3rP8vzHsDH5EXc4dTc95z2lR
c6+wE/CFcQhtuk/jtlPfRaCOFkhfJCrKo4TapTQ6eLmQilotfJLHPjoaYe66
uRWIn4tlzd4QVjxiD1mobOHIlPN5BrAYrCOjAVCKyqULFPLtbacH7RMwbLSl
oCW1eqWJh3WxSgdzJGxvHNOIwjbxjDomkeIv89HAbp7V3tFQSBWkX27bENI3
5FHQ3Q3TSj1cyW7KQbba+Y26lC9NbcqMQDwmUDp3vXnlX3bstwOmqE4b1h49
d6y/8U7Xo0TZ4cWjuGf4yLn0ihQJ5pkHpYithV/A8BPXtjFRbpJMgTvSFrPH
PN6FCF4NDFcj6qBqnu0cJENRb+iWSyFi47wyWCu8ZYojHmXTPv/IVyVK/lDv
sg/HcHpPZAXZdrXW7uc+SNPA4oQM6zOHrCd+7P25LkLGeCkr0oJ5XcvWvQA5
kMH0CDSXQXdknB/DFwju1dXdgmpQ5M1tTms1LuSMJvHpvwpaEewhKmyl7aWn
5xybU66Vdrzhb5EARqF/BeHBJCxd2ykjRuFEaLC5ngLGfjlXeR2i22i67wQl
bUvLF4e/5M6C+TaC+o7gJHj2Ku7BP0dytGqJPWmOsbmva1k33+mf5um6G5+l
RnAzOtexowxcj/NWjNsIll3guKUmwH8wPn0VCLbUNJOl8IXPK6YNuo2UR8Nr
V2VQ29ROGn1TzOzrx/NTlLIiPmIFE6rYkahdXl27HqE3hj8HKH6ic1UcUmnI
NluMOYbwzss7KOox5beZiaqhjVLqNIdMWDu2I5I+I5SIqDEyi1ieA6dnMy/p
t6b36PjDHAqYPatDrs8au23T9XO0Y/RYYGpeMS77WUEIWw4B99eddwNCZKOk
toK3djlgjVcjZ94AUCAkiY/3iXkYBb4aC4NpdZv/Lo6q4C6iMDdCFTdUF7bq
E+cGctIUJYgrIN4/+1hj4MsT/Hwwu6RAjAa1y7mclQPcZgk6hik7uwz4MgYZ
M9Ps0AR4kjnOKL9psNBPQHhy6ejwDVegSHzc96UuTEVs7uLmXXugM2WV0787
Mv8fgpLwXyx5RubXqxrfLMs8jJDPOMbLlMz3069ij9Jb9cb/sPjVF3ahGY+L
2HGw4Dtk16EDu3Txuk7LEAv3IXsrA2hiTzKMn3KgnFIXQf3MuOatg1xgMEhb
9mpkYR6OB/369efFOuoa+EIgpHSQJYGExdFnq+9/BWp36/+ozYud2IvY97C+
egSx1nW5Rr7O1SI79knV0J3BZVfDdi4/Qh7rtdbcWMv/atbwaPW68OZZObg3
iBYiZjz599KKYYTbWXwHwjWN/3U7k6LDxAZPoDy7hMjtrb19jcqrfxtUuVIX
O8H54gn9ynzUi4jZoFKGZz/vFgiYIACgoCV54tpFDMIBLbKQgL9k+kjboOO/
QhY3rR6baDCFpJyC9xTxuPLOOMAQeLrHUhexU504q0kSin5LV5Ul1EVXE8ac
VpWSFLWn0KbCKpIKEUpE/b77wJ7g9jHjTS17XM2QrgQQcTNd+T/QAgh/mNTc
tLZ+j3EfELZMd1vhRKaVgfsKfNDs3asf0+niik/cz7oC+ew8h03oMqvA5Q9Y
s8zTALydT2O5GFf+gxPARtZSXr2XFK4R0UFKHDMrNxWa6PXjCvzNsTU1LMm4
Xel3srtxe7LXZWOvKLwjN4qrEwbO26wpLCTnX55Z/1iAsZDOfegpMGNhInfh
0GT4lWCY9k2nMn19O5sb2kUawi8JkGQvAXiqhiNebXdL84ilk+e6f+2O+EZw
hjFbBjNHwVqevfnuhRO37h+NzdBDe7dKeiQvywGfHdniDHrsn2P63KBLAAQR
lnKxV+sL8A0c+JCtlHpjjsHRt8+SW/+cXvgz0wpHgg85nGOHiO6KFQvFhji/
4JZ5BVteaQmN8i9CIO4bsn3oSFodBoxEiowOmkUBqwa00ThwjBYmTCJSG8LE
U8UEkeyKHeTGL07ny0+SBG7W/nam8FfT7YBUALRI/TIq84QHQp5zNn54NfJn
xU2ERjcBwpHJIdtoh+yRcSnIYZQXPQLXoXQStwEFJYPgdizKQJ2lFXSXBh+t
P+4AqZvmMfcGkdykXAp4cmx9ae8/+CX1qDtTmRGpKqc7PwzTRZycRHZDto4s
4WAlgZdl4rd+y+O1Gxyds3Om+0OTZC98I748DY15Evx5tDjyxfMqw9G0HsJz
MsJhewxj/huWg9TgXAumRvhSofAK0D81FIxpixZgOEDlZMqGdXw6A4qV0pYg
lLKYaF/LahSU9aHqTyWKQFA/wDzhuSeGS5CGkUXjSWfdSv5c9r8aFP/rAFD0
EqGW3GZXYtl9rvKVXINhXZLl5BAAQB3yz9PeLNQoXqQN8lQqdCrXYMcQ0nKU
W9iDgX+u7t58X72wVPoLBaTr+4U3JOk0BXiV+tdl7d8N/cIaCno3Vb8/tAzo
0LSYmjgVWBoIM9Xj8zwUr6XHgbGAJ12r26Po94CIHkS6830cP/iCKJOKjURN
M5VtmTrh5npk2Mw+rrSxpVmgdqyNXMbAmxUcWubCNdV1ku+wBWDbXUGLVE27
Z7acdUblWYDaoQ1P5gHFyq2ScrvqE9Sayn/gCQtU5pC9Px761UTsp8UuMJKO
4iOd6EKKl8bIqPa3O6zjLB6Q8s+z5C03SFSHFPISEs5unr568q2wF3KvVGz6
TlqmiyWPNIpAHEDIbe3JLFYegx6KvgNkRiTLSOv4Q/9t99xugI6Bsa8OLw8E
NStTxuXL1Qp8249MK5HZIv2ah2jjscv6pESYnBxCtUBhEXwo7gHeneymit0D
MFmsuFEwA7NhSIQKFz4wuwXUW6bv0IyrMUZJ1a2Y2Se144Er/oJlQzEveIdy
pqh9I83Mq4JDRCLO+NNz+eYAzpRIzYucD4tYNqAuH0XGd4h01DgIAA5iD1nH
gpYc4AAZc25eIHbiIU64V1xnPeUInps8wdENsNx7PSAPtP61IbYXlcJ7yCSl
NX3cVTpzalCyduOGPO2RR5ZdtizaDmKH9OhqCIo3c9A28rH6fgkmL1WoBdwq
Ta5ZOXa67F6DJqIuvgRmIJ4NZ9VWIVA08MB4of0TPXHI3/ZBaw43S2guuhlg
UUEbjT3mbFGbqHZRi5moTl9yGPZge0+NLrjsvLfPfq3/JD6+619p+RvYnHkx
gPathRzBzlSeIbH+y25YFvjUdVvCtSm2Yq3zC+yH/gpMLaz/wdc2oFeo4DCT
FWB/bim7Lj7uFw8xt4y75/ownYhtM217r5kwL0KHlEG+pYLV3WidpO/Szv0V
8REmFWk2EjALvErb59K0wBcrENTlRyKsLKbkgxouy7jRfBBrcRncVc9saHQ0
0Lw+xcBMFqtX7ORy+WHaFv2IIoTfXpfAk0b/WUNQl+E43E3s4GUYRXy9V8eI
aTiocHswwwEKTFi5dV5KWf7K/bVpcPyIdApEE4wJEUlLeFFnt3ln68dAAbF0
urHr9PdQtRKRfxH+zTOQAa0Kh/Vq+f/W3A40GLX/NMob64ED/xkA8xHGEAl0
tjeOB9DRqApm1n7ikHKNejK04DqHEneL/WCgHz1gSx6o9WzWslX52G1slN/F
KtEnIa+SS6RMDLRo0q4dxV8YK2dlz9qLy3VGKT3EfdEYscdIoM6TKxNgEDVs
O2YLvlwA1y2pAI7hK6hEzDCpu51KbG6lJTwHTygcuwKqxiSUzELsDgw/iOeI
flfjm/4E7AQgchD+aAYafCmsTlfqozdIKpepAQYpcimP4jg/Pb6wlSfcC+O0
WTt8ZzgooWZ6tYX+INH3DwyqGLGIQANcEaXDHh+rU221muA2yIS8Z9sru0ID
WZbaRSO3dXy9mn50nug8HsvLVResVo/D3ZnX1FkVJALeV6aaLlpsJU78WYm+
W+v+VXxVUveCd9TlAgjLC09I8LnWqaKCfGDyDXZwO/4ZXNoP9xASnJgZL1/C
uXk3rZ8W6UGL58Mvx1d5neXXAUM1t0390Lw/pugrD5bulP7SZz86IMRBXGh4
gjBzLwK9FdDpDq2WtxndqSXRSDjZiAolG8PORh4wIpTd0JIdV4S9awkBsWks
sl8bTCgrxlbyRuNCRWVXzpaxfbhtDR9eKifwZJGSQEefLVOd6jTj0t/VvWLM
8UiwphD7TObWu6DZ51sWe1M1bwRGxNTxDrsAFwH5M+RiyfuNHY8Dmo0rbHMs
vAGQVH2lFC4kGYJU0LP+4qYGQFrNBv7fwwjF+6hseqC+UuAa8YN+oJdkz71r
0Mh5wNov5SiFZnFiGlFgbGuw68/CuiqomeMm5jCiLWRBGdS++vXKvs+HAix+
YpqQnoqk/ZeUvgwVXhv+zzmPwh4Lb6OyIiw2PR2kjCBqcqTuYqOTkFa0kzy7
henTNwgsbejKQxFDWHD1wyEirABKTbR86e1cg9zBjjkmiWvU5NsadSnVYWQe
Nfo49HoOlQqIajiDJ5mzVLvZxugTHOoIAaJ3pNu5Z4kcUqHFzGNfu/FIoxio
BQYHoWe18zRbfgiB3CSDCJuyK3TNjdAqTV9okU0IrkAx8NrgF8l0nthA/An7
pW+148PjstLTmORhfkBwf6cHobXGj2VlNSKnfoHFcb9o6V3lQuMsemt/yq8d
Ube0xLR+KC1REWpFFuTY9Ng+ztxXeol1rdprG91bs3OHu1o0M2B6EvWYnCwx
5hhnbmBakwEBc/lV/6Zc6HjKQMBxXXBxe03MmhaPZuIglraXmq7VxOU5Q5RZ
FcYeU52PYnMgZtxLK8L7v0QeDJtHgCDeoisXoX+HJKjVCapO3KijTgBiu/u2
1uMQOVYek7D7Z+t+Eg8uoRUU98K/irqzcivFhLOMcZpAUIhxl5wJKiUQn7kU
EMzID7bsh4Mj55Ec+ji8+XfHif85109QFUCvCj4QjdEI/sdTT1XD77oJj9BT
iqCNpEv79nPiolulPX3AMDcrQXwC0OnVUwjpYXtxtSvWOYK3e8zLhrLvIuHa
Eu61ULW97Xi+YlI53AZ/poOMUWVC6iFk3SVWgOtWbJ+LyZcEfQKKgohpmjUL
5Jnv9LmO4jINf1f5ZpeJKc7/mn3RU179ptCRV4M35Eao/YL8i2TPLpX28uvy
2nsYqaFh9dP2Fg5zx7oIIW5Nv91sMUpqz8fSCokcFqBR+AwdRa+AJKZ90y0I
rrbN8hfGsl5BYi4JR8an7VyuHOQtTFItiYHHOEMeloxVhNusSfHrBGSaBCfn
nPESdRHfqxBv67t0wYRPJGwPlDuok/1gp2yWasU8Js+LtqKwhRI2Yxfqnatw
fkHYWWYiVbReigwkTCZiQfaHXGtKCGHbSNQAWISCQ7FuLQuQZqlpxSRAF0Wp
xHPkwwlxywmtFu/5XDEbGGVw0r8FrbdVS8r5yftvos0rv4pBmfoMVLjgR3Ax
e5PEWYB6CgD2jCFAJFC7UXv2tmTRC9nH7/pQlIploaCnMbLCT8IepQn2Shnu
xCeI5pfFjvb5bgCvDgVOmJYcvG1cvTsKZmUlpH/q78URrhYcySqHaRc40i1O
p+VXKh+3W8BlhBnCo4intX4lJis6IRzSZ0z+J+vzyP8iUi7Ssp2L22HjKmrK
LCxqO1Cm+sQOsN14ulyLe0CXiN+J7KYzXmoMlLAr+GYi3PRvsbwJ2YYcXJ68
PbS83wo8kuJdDjTe7mCBZm9dCkPAvtIit/6FDY/mFeTTabnQz3RL4CHIlTZI
83jkk9z8dcnE56tX74x5ASB+qE6y1GTMd0m3ZGi1eDBACSQfbBMfoR9PQHR/
5Ej7nh+sYIknEoidEsCFo/Xz09WfZW8rd4f9qEYEYG/wqocJQNrPWtWRQ7LH
RRianqZNuPRS3YH9fELxs25EyDpMkHvUdSHvwjbRejCXHEa6eCtTRl7icOfO
Gyh2tN57LIIzPt3kc+DZ3ytZWZoKrK0Hfw0owL4aTzGZvHdfg/148UPihC9B
Tszow3ZKckwou/M+N9MND700ZFmUeHZVAkL3jdIkCgcqcoo5252firENsbqH
125JFlJGtZ62K/uP5AfaY9HADSzqB8JZcP8Bj1lw9a6kgHCfRihcNiW+wb3s
toPgcfvn3Hh7qJpgxHVojKz6PhcVKOubphVFhu1Ppy5U/n87yUu20Zcb/jTk
gDP9Lza0AMxQ6mo6onLEz3nijeZbHbRebLJ9FcJlo5IvJaykIEUf1GYFL4qt
UJE6s+hsgw2YcjI5efYrSbuMouLIqJ750ZG1VDdOdnD4yg7qSX7pV4ZneCZH
k2iU2e4zcA2MlCa7H5b7Vxyha671b2e9trXFqPv/87RSzYRwusGlowAw16+s
C4OuQOP3/ymeYs9GvVqJCrUUVc/pw+XasnXOGodeFJJqYudm0qzvya7dHIH4
ut22RkYUk2QkLw+MbjgMyoFzJ1S9Q3tyF23ygGdYe3AFU55gnsAJwIw/REwD
KFuVUcq9rxvbPZALDO7C+zl1fWm9DHOVqIjh91cis0Pl9YVOM2BgZgNnLuca
i+SBIj80L9VSJd99H4TDdDrG3MrLhObbLEtzQtjUnS5ywsak12wGrrJo5ePq
PEo+jYp+1YILjVlzrynxJDqdt48djDz8d9M3mJv7pt/Yk0E7oXwj3V8UDdTu
omZ4i10ghRSwrnfFQXlTnJNytAzGo4LMHSr+2K9UQwD/Q640sRqB7btXZYMO
H3SRneitBL3/yvRl8BHZZAiXnxTtjRmcjXA7PR1D0829YQC0y5SoXNtlXB1g
hW7wIZic53F18h3b2T33SOhmK9WmFbfKfxQqhkwpJzdvd3M4Vpvj8XlInI1K
7GhAz/zouD6jbMoNGXp55V9Bt7s6zZjc2OuB7rVWZezZFO5QP3KdFswf0lWw
uRqewABfbeSx30j3NF98L1pue8eanXYQbnOUoURKXb5vR8xG+f/tWSfBMi3f
8rwCbDczcKXCi94XK5erYe2/blKepJbCaadbPrQ8eTN+K09Q/8vjLT4yPvT4
So1CJvm8Ipkmo15TsiyDK2kCyzSefgLz6uixtmkMbQFWp+51bFR3d+64Etgg
tl0SHfFqPwXZilapr/p/KGfwzcxB3HGyzQOt0em8AlMDv/Spm7tW6uilotwb
b83kKL8bZi/Jc9JOUpeQQ4RxPKhZsUAYr1Noztj9b15qzx1XA7omZluwgNpr
EzWJclg/+lY5hqvfrnR7yE5cGQqTHX2Z/ZaVTWmvKO+FXf6LcUmc+3MQWUGp
RrQVOsvCrijh22/zj4XtqYmGVXXnatDHSYjHWmyPQGneEcimfyjexIzjZtbE
ff38pk1qaLJM85S12Isy2tY2HJ0Wsa6IZL6hXjVTAetSS3QVP4uAlQ4hJqa7
BRDCiFZu4qt49eRuk7+r7oc4RgRfjtzGrolARIU3zWnlR3jXWomHcEH9zu2C
cSt9MGDV653kORh8af2Rpmg0EkdS/n2IjEH9sly1cAlTt3FmTUQSLXIagq3N
/Aca4OI7a0ejaUulITjDmdMns00NncIK8yBdQT1HQFD4S3cV0iCA536a974j
2bEq9EaHVwSx317ASNq1IQQZMiWd0r+27VFNZAAmrH/7wNOYfuJj6s9Uztlz
MN7tJEPizSX6YQORl9IU4Ypxqw+yM3T7JTcPWckDEQEInP4/XlKvYCwOhUS0
xWI6EAfxhKBIwRz0Phuv/3C/cWCI5yuTIPsouHQYa/S1CZ49x8y/AiYxIftA
21qVux5iOgd2y5QeG/rsayO++nFwtNZiniAEyhbXEJRMeiepb35VJvziFibd
mXMwznqXNLR+3edeKiEMlyQkekZP2E5qaBPptTe612RBGcW5PNHH1TwEn4+G
z8+1+SidiobW5OgpoGCRtEtQKMBldNvVEM6/m2KLVozzmMpxULDRYI8yDYzp
gtFlRn4rsHpmM+MgXNe+Hcqe1t+FswdEZLZAgXZSV8Fa0Vpnii0xSJhwIdg0
9JNkdX5/Uq1hO9Uok+Rx43ufm1RNH4k+dhChlAlGsvUPwN6nApJ/bJDiQAd0
W0aydHtQv8fLELZLG0XDwA9TaPUB4ziR8i4rtA9YjH4zXJgVj+q8exHUBlh3
xV4+5qsT3iJA3ZRNJEgKJCN04iURUOTPilzW3fZ4VvCpqgCYKfgboc3wQ/Vq
aXr+ml+Aut9Z9GknS+rTL5GZZM0ENUALB2xhbyaEXmTllj7aztHpCGKmKzyq
BDLt3kFyGRuWzMcRD2W+ntbuDaxR4Zgen48Z3/0JUfWmsXmGcslve17NpwXu
dBCXvbuFmzQqcSAvGf3QsV2sEfT7ENMVdpzPTtspjz+Vp502QNjOfwzNgAIN
hTpG+WzQGmF1YZ4CKrZs/EjBpzBk/Li36PdlfYU0zr1gCsLJgmg7YlWr7wmp
SMfjcoMHSay00Anu/pb3d/PmTtUl12fQDfC9GFQ/4fwKQsUPb6Va0fsvYPd7
0/PO7Lt3XWwQGKB4xDw6UOAYe4LoJ5iEiMLhc4jQNi8utXbkNzBROmSU0IqM
ip1N+uXLLd80BHZWjqvXsiq3h3TmaErwoIQlbkJ33g2pzUhsaqYbjvLMss/v
d4Aj+10bOyrUvpkYZ7u9bdCNKSEErLdY4WLa7O/MveDJNppHEl9DLiE52JO/
rbL0nSmB/V/LG3i6ZXWKA9F5uJMsh0eMwbqE4GpQSe1XfaT78kPzaKVarJCk
tqvIt2Arw94yGBBg0CN7yDPZjChC2XrgDm9WAhE3whMtQ6Kkn1IKPllEv7mH
1svbZ05L2DDfENP+1S0Ob5eQ79bO3BYaEVhIipELYNGBisTxost1pU4gbyk4
DyWCsdLOzMcJTUcg82MMra+rMeL7eWTY75Hd443QA1j3Abbv9zAizGM1RhNH
6H1q7V+RW2wmVfTcqRaXogcSwXqrTi3kg1ff7c2LnJE3PxNchqFGALUH6gSh
WFg4ZVPLcP5RyNsdXZaw7QoCm0P0eNCvqX6cWkMIqLa5/CALuJxE4ipkKueR
WcuWwpDRBXUuNKyBqBJlxQygwM3CYRY3mwllbsPeNzlsrjmduGvELg0J3K2h
EnpmYQsgL/bF9jVZ4vnr2TYhdHfcEz+7T2lVmgzlPwqoNX18NFJLLhF7uUWk
MuSP4ifcvbg4d914++GrDd4V89JSLJZaG4bBTqZigFxuMvzKjV28pL8HpgsM
95ju+gMqY71IugPQsh0Om8165pqo+FxMOZSSYhzl2Cdr4fLa3b4hgAzLQ97/
Mz65l7u4VpQfyieIAorHhJgQOEmQweKyckS4ye3Vw7kClL+Uw2SuxzIV9qiC
RrBx6yiSERhuA2PoFhmgro921PQVyH8oWNxbF0ktnGi/2Vk4rknvgoJZJJEn
N7XyUBd/0iJg27hsWbul1PrDI0pRvEg7eTUdiYbwllccAiUrAa2s3kGJsyxI
nr2LBM1bwPJRkPY0fxlvXlibe+g7QCaA3qfl7+bX1VqmwaseKGoAfMKCPggm
8Tn5NpT2PZkRUz63EFD2ylrWd8WFiE3OCOBfpILChP5fUdvL6JSNyKbO9nnL
C6WDWYFQAq2U7+DJgU/ls/OSa7vgOzbBPW8OjIYy/w4VU3ZgDezEzopbb2ay
7pzsO0NWgbn7g86mfenY4uYwrVIfT/Toiygzdpo1uGisJ7fPdwjc8MmZq/O4
8Gqy/5IUngoF4Bk+fHq3ObFxdvT032on7OkJdssOU0pGFkE5CwYarWEbVIod
cTy9yqFEbKd2QcGVlEG4QYJo2I2EyekeNx3vuPxnQt299Yp7nPD/rgRGkyss
DC8gyIZorZrZ9r5q0aQaKYYGV7Y/VvOeA3bP3CLS/PsmEIBQZMHHfmizvwBB
siR2x44qRv80pnL3Pxbhbwp6sSergznrTlAZa19ysp+LjcNtLp3JwEuA2C8j
md87r68ODF5Y9HhnaJOcmunW8Jqcrge03qOvPQ6UfsqMiJz/tspD7W/XPs/B
Fj9xgyy/5+qW3+yAVJF/DSai7jf0O27l8l5zF/48kZzsOdN1flJe4h+9voQO
1/dAuiyEGxmDdrWnRFjL8CSOo5lE/Nxcnaw3bCaKmaMj3nmcRpqgb+oij5mP
/2Ml6OV63f1f5M9zx5iK24Xi1VJhBB/uXP5fgThcUW/ITYHu6kF3HaNloY0n
zc16jMlD20RMT6I7MKcVbunOBo+C4C8h/naCM+U9RkcwudPCxDy1gB0nlhv5
Zxe280kDT01Zhi37ESgVFCtdfjKYmOH0aj6JbUFVa19quZ0/JmZFxwNdqCP2
PcsVTEgEIMqAOjtFatONMpIf/ws5QMnY7NP7bKqw4ukmjqI4DZJpzyGHH7yq
NvD5gxqS3Asl7SzujrWi8QzDWgELqdRMFBwnNzh6g38bfYWCqp6c/7MOWlbW
A/Dao+zEDfVUtcBAQa7wv53EoKDg2rto4P6p+DMFA/SaLmOAY4bmyvyD6s2E
Da6h+CEcLrR1GXjXRpzUr42iBMsAx4BjiBGQw/WYMNJW4ghdoA2AjEiouz7+
Z5LPaQ4u/amtgfyUrk0YkGAcEZgnZcj3ZxwCYY8tpd4XrFNePXn4vXU6H57A
tCJB1QZysTnKZ27Uer9mQhEu/qV5xu6e+u3jAZOf/T8xcLd/7rAi9H9GwTOa
FhAzdB8G/exi+Jxu+CUNyLzkEOeNKu7fWvtwaha9tRg0wU9NasNgmX2t42en
DKLJDad5quXMklpOR20jXY5zr7CgeIyAN1TW/xdfl5i48fD86gldwh2S7unB
Q6L3kAoNoO7RZxIo56HUnAdCPfABzL4ny52PcRGKajvYKheR4pQ7UKxEgsk3
ZjjWTyF9EjgaUK1Gs127M5fUHIeISKZhF/F4K2azPqOARse6/h5xn5ggT2+E
lhAa31I41urRNkHRb4W9YUtj0Uj/0bPcezIAtoUEnEQfpBfcQDI1NS4RseoD
8qcMIlK+MmNdB0GNUiEwsG5uPQKj/CqZmqHrK3Oy7vce7CUqaItQ3sf709oi
TxpdJDprFzW1w50m3g4rQYONWvr3b2ceJB0c95NvY6PnwVJcCOjuQi+SDNMx
NjM0/4tJ170lGbAd0XhLe23Y7FDeK+4KKjnRQ8W7oDYQO5/rBUEnVHqs7ovf
pdFvVrTCOUosyocywJN8F24CJgj4WxGQnzSwpNzUj3pi13+NaNQsQilStGon
5pyFiOd0lO9nwxVZHfyIYdKdmtZNwRVFi99bAYe1Wy2IoXGCNIAieIfKnsh9
ohWkCvlMhM7RUAuSPLB4OFsYMFyT83d8YBDjGg0j753KmEEa3bHEPmUl8Qv2
pEsEJjIImUAj9hHaU36ANKw408m/22/jhgQDW6mpvZDF4bZpCW0ZfGW8sH2C
0HhTXuBWrMlDcWud+1LlNd5OUoP57av+71BlQJMvwMffYcKJ14p0UrjWMWiM
DFqZfOmjbRHpZa8aBE6RCSprd/pjeQ6XSeCOW66PXK5D15NoJYdaGryPOwSP
2Vxg5zxfXs1RwrPGIuFPmmPSpVj/gdDEjiC9JxfLHdPGLGPexd7UKUxOEX68
RG9ASSb0Z0MD1f2MXgE10CuCr8K56CjBa2LVMOH3T+OJawG0lfChQUk9TPNv
/FFxomBq7VBJGv9ud19qcvSQJGNlCiMCptvROL57ZAd1jw+taXMqWAU82XDv
3rFb8J8Ty/NAiS+HwLCYo1bVjCiHc20GolvZ5vqqTJEuWIfYB9qoCpzFFXgh
5ugCTQM417LoZWYCYIm/ch5u3Rh5PVC5rWZEDiuQMSTq8zkds11St/UqWW1/
hJ72xVau1TGQthL07/aF0Q47BN+0DQUlvJUFYm/GuxbJDxeL4/zgT91FBeiC
ggO5gMwk8C2tZsBSOABXd9uM/2kQWdUGCd0gSbmrdaINnceh5rrGhJQ52Rwh
uhwRqWy9t8fyiaLWKARnexCgxp/FK/3p9+uAhewPGSb2pFTr1Wp8NIBNBXcl
vjV84QTzN1xdJdWs8hrel/XjxVHqID4cgRxsU9pczaW+gtnEkb6tq3PkxEsl
+YOSs04ZK0mS+Dic6FB+2ZdwxlwRFSuQTg8x7QdN8kK0DLWFFwq635GGp/Ff
FEmZ42Gzg91iaQJU5maEoayPTJKzdj8E86krxITdj81IT3+oqWqRQcVvi/RM
pU7Ja3uj5LZ3rtvt5H+4mOxZTJuQjKtejcKl67Uaq6FudCjv4+H+C7MFdc7K
/Gvi5otODXmlXjm5HLJwibNch87Xa+xEZ3PXi8eGwg1JzTUN8mSczMKHcQ6x
TRLn0fpUlDP4FKEPuk+w5apNE1B87vve48ccB9SZymbTWYA6fW0nJBRyV38F
ZcOePo1U2o8HGrqB/Y5jZM2R1fSWt+O9x07aDxEDb/I6eNWeSDWk+xOmpN1c
J7cKp2X68g4PqHepfIYkvp78I3AfRRxaMCzVYuCh2NA4zdmrgURIlMUvszKq
6o9crV9itlb/Ott8qElw3hH2qcYsHKeMhe6VnDr0lJIjbOSbsadxIbQ+Vblf
6HJnorI9y+UaOgU6xqZ47upiSUAHeH5mrE+8ob9ubeHo75sbLswbq1XjFxqE
hypcu0p45LZUkfBCLYxt4rrrXPtWZiwITUVqktjt6FVPRtr7nxryWTiUOolB
jPoBDHOUfY1Fm6xjD3hNTDyvGdLCzQOJ/4R8VzPHY6H90gGql0Y7qupKJQ4R
7pGTfgLhkAaEmD+09toCoK7A/ymuAarYCJ2WDcdvq4RV6sSQLo3mS39xNA2O
bHlcDhaOs0IY0GM3IZjpyMnS1eR6jpFshWSSH+GU6hlBW061a4nE+4wf8BBw
6vQYzXINEFLSfi+Ge2RcbB2rxUWIi77E5tI+0w9KVUqzRxyu1XqxfoGKbAFD
P3xt80AefJ+5tmt2oQrQwt0xKY3+T4nqAGkJ2OmeAo4wdbLzjGARdAL9yZ8y
/H5P+UsQ5Wu1f6OwN0Ko2xzH8bbP9/DwVy7zv+8hZ0WJwRSMZLCKO044KTRi
n3v0bKXXdXDGFXcCoBzaDHqX5bXTZrY9xG5bWSoCG4gKrnCQWLR/of6eRapv
gpn6ebdPavjjnPOHUTexdwCd7V6709fjGconkXXGIYToVo2mB/N5pMHLogRB
F/4fALt6APYgoaeW1tNRRIEQqd4sOlQyBWL3sdXPaoM8h6vfvgT/axig3Uti
eQfh30LFQ7rJMMbvyTadppKVsIxAiJ63Iu8NpGvESjqxBTe29TQAJs8goTOL
7BmN4Dhi4c8qgx7L7dYqf0jz+SNmHZ6EaWnyHiprchgXqKmf7yKtOOnCwBrj
RvntikFMvmaA9rJ9iP9+yVu+/7znrQVKCPJMwqWEExsX7pinexDoFZcrQAD9
a+XPjEPskx3ePrUNPEMmA8m7tQapVgszTlRmnmA1Gk7Tup40CY0nLoC0sEAi
FGqsTX1pKswXoyUWex2WlJ+VmIkOa8EovFjGZ5HbEUlm5BtDcBkuO7USM5b3
7Uyyam2jquZTgwdGrU7xqtizmddg3f2RymetCBq8mQTd727YmAOSos8SR8sR
d7b44rPU4NPyHyxpqXMSl8+jOX9Vso2e3WMXcS3fpAE6bF1fzjjjyxH86WpV
rkSTnKmc/7n0Oc4QWQSdtWerCOhbcwyOeTTHaweZLKFIiGuSb2A2qKtJgmb4
WAQzT32liJ4JhFwKft7jJGr30N1Yzoe7/+likbBThFFb5JpCdYJE+RPrUC4M
ikYLSoTERMdhPozdae+uZ/I3JCtDKgjAsqbU1b4O5Q+CPnKt6jA+ehsUNOvr
7MJdC/PUaXmed8idrrIrqc4kkthN3PEQKvYvi8Nz3V3K612MMnUD4ue3539q
3y9JXCyETqhs7tdbiVYU4ydJy43UjgTsYLr8djFdZW4lVcANhbJlztcF412t
jP60hEk6f9SIW0mGHZXECfWhFIMW7DWtrEPW+rr3zFQ+9taqqVE7e1FtEH11
3+TkWG66ZLGR9GZiDiA0VeP6lgEnG6pI02VOlJeFVbPEcRlHt7gEzLmBfomS
6gUBOa9V8qiVDwonc+Jh80DJh/reFN0tquhjaY8pTWz5FeBIHDQEBRfpx9AE
9oLTt8Q1fBBQXij1Y4/7KQ+cIM3hj2aF6d4+jwuvBoF/GcFY+y3LySmZzZIE
NgQZ6T20jLxy7PdGQTUnHQJ4E4sy/CfB9r5GDBH4wy4Q2yQf2ciceFtqdS0h
4oEsIe4JkkPzHJBnO0U6zCOxzVOHJvMMLnFhWO22A4yMe1HG04XbLBEcgkTe
M+Pm87fe8yN5+IgdE0IOKXzQscHA+SKBJtbstBxf/IuAelDhg5uKSHQ9SXP6
+gS48fLMuGzGHCV40YMomQU0BlzST3UVJisddC/qV2kDg1k3N78bw61QUxtk
76aWPJUpW+c3gARr9RPLnl35BHHEt6kNLFOpC/ywyhc4vcjym7WM2ccfv7xz
IZkiMP1vkD0Mf4tQ7ipYKlJ9goCb791mS4GVDYN5T+YoRd4o+nx6MdPGJnSx
+T4ASJx6ykdE3MEen7ZPuunLbdJFnS4fzxu/ysEY2SHx1f3BEDCzb2vEphYw
cmu5GD4+L9JyK+Yv8LGty14dJ3hwN71tBTAforCL+g1qZnxQb2qV9m3JAWac
jD2AC1A/CIcXcf7uca/NbmgQUnsiKR2G6dAV921kADdfAC3IkhnjVGYZo5ls
XDvp2tuk/OBuZX7L87e8umw9oNwmPd8lGj6KpPQpQ+BHgxhg6++8Dy26ZkEV
BuD7Pz1+hDnvP3/KM31Ct2YVqmUU1/L1uspC3AyzAWR8avrTPECyXFIWrLWe
8l6eNpI/J9CR9OTn4xaRt4LUYZTuN3OTjTgigJPCS3PV5k6sCjfulZCMdf7T
CTPDyYZ7Glam1+nPFNv9q/mLs9wXKCrZ4FOsRANYnMT/KVyfh/Ow7QL4fGKQ
Xq2+2m5w+2P4SO99DKsWAufGUmlJknCNNiV57L8fEWtsrcXtYYm5nNTUP4Fd
KUn/mtqOosyN8IQ3ypBOMMkjjXpjSkqRy0GlLE1dO00FQEKxUPRvuRc0gan9
jH6mpvWrIXg1s8fE+zjwKxG/O1/B5+PQ0UmakEpGa32thI0Tcv4aQ0ho70eP
5BwkprQtIc1ysOenpIRpwmftppRtas6RFV5/b7K0qPz9MdI8ANPnd7keIo4X
1RvtKJhI7492ydaB+8Wx/R9EbnEOWjrIU8oCzin+M3FAzJE3af0s9VDD9pUD
XzX71DqiR+9c9Rky1DHfQPFbzAJ4UIOWliQLNVrGIXY9l3Lom5766nvF4vDa
2chausXcKeiZenYOYulVxDuSE3Ufuge1tjQIpJETG8a67ZTazd1HBLZo2LbY
Q92gzGVqJs3BRU8+PqufCI1QmMKdRGbS/1+tuCsb9wrUcR4tae9KNq3NO1gM
cFlAp/l6BEUguFpGczci7QIoGoj1TTmlLGr14HFx6ah3NgwioXXQDjLPWYq1
DFzI04JjTojS6LvUWqveZkntYtbJfTZt/R7hGOrAxNXWuzagiMUq+WpxVshj
2Ku+zJ9syhN2LErAyDYP8rYzozciRuqS2n42qPyyiQDJ3OLqzy1YMojGEk/0
36WuXyXYx0rWkjYXYlCJLD5zwPx7U/QP+NmB13S2ZTQOfWPpwKPd5tfeq2wL
S5/29fR6We/skma1VD8ZzB7A97mJJRrUHKdUDZcaW1BotfqDz+VkeHYGvtJg
VGvIHye11nlsJGKC3OMDGuUPXEzxrTg9XQR8RpuhaHkNcaH1F2wF4iDHwHJr
4U3/YrlP9hvvlp8CvG9+5xnmoM/m3LyjbRdXc9swlqxaFEhZA2oABrPophMZ
U9Mp2ZqjZvrOBOj/jdrm08sG4JIyzrVCZ/FZijnlFOKuc4AQwcrVKSrlb0TZ
qj5UCS61OFv5VuhZ3BnBCI6cauXqFzelu3equ1yKQr+yj2WOAYznKbXA8xZg
XPq9zB9AiBtDVttoB4LyWbRkA49rZxBgTg+H8ezSdm2Hf7pQ996ZmRe2RSob
Git44PIebwBnqMRs8Tj6eSsfy+R5/aOsuWzxueLgPrFHKOifHtrxqU4KplhH
dakWM95nHuHxxjBxZCJ0Y5oBUHOjRTLORUMqmzsO8ifxypgGhOPVBbU1Tug1
/UduK3FD9+v0I4vRpGq3gfAqP0AeU8YxFL4ll192rV5dmEokyoe1XGHbVaHH
KXWZueL8vVrPe9ixwqYeLt2EzA0UILbbulZNUTyHRXBDib0XHFNHdxfcTXxM
HQYV2gYjJ8HRd9eqd0tHxua6V9pEA/bl1TOtWu4tZNajki/oGqjh6+BRxK0z
vXCJdX2wt9Uf/tznXY3eKsbeEJTsUwuX0yIYxc/kkLoTNwSU4v/AGUXEUWnG
I1ihEmAMUgOS5wmtjaPzmRzvaqs3Eno0qshWlU/c1z0wHuHVKUlHPDLvyal5
n75VbAncZmM9k0/jY8Jj0tKNF478S22StCVvsLycMEoPRCocADkmQwSSZoLe
t+MyZ5C9sWoEL59grkUT3+C62nCpAwAwmBP9FWPrS/lWWcHgN7hQzDZhSK0d
EhQzjmmXMQda3O38luUOM9BCse7sffcg/VMkE7Di4XhRrHT8VTFpXsiqLuI6
mVCjjDLEOplWOhxxABXmQQgR0VzMM/y9igV0PHsCnuPN1zmRovxf1gTVhBZ0
X8ln4DXfZXUXJkiKLZeKB6kiCC9cMCBzzvfzcKQSFMi8uul7VRsef6x82g9F
QbJMcls2O3SRkCVJRGgeliERf5AIPXUfT/dH91cJrfpU0/uWvcMjeL/x+OmB
X33HKdSHerVBjiqatNMe8ozUmjC/Q6/GALxlAwZeJBtze4EsHDKxr3kLn5On
XaCddqLChpXpXXKSC1EWMOemlQ4lHSkB4VtPS96lsrtyA/lOLlQrhVzina8g
ZWrbNR82XFvLTT/qliMAaeIbFCNLsNg5blz/YM5nf/f+DhQAyBaFZONlRpgb
nUA5K788qcZGNfk1yQVtG8Pyy1OdKI5Irv7BJ/gNb2tiwS/KIK6WS3Z6Wkrc
f6vjBfKjrlyVs+ln/WCZ9ncLdCu9UcPdN2UQZSSJzhObYaafxf9qcNjomsxa
ZxoKAbY7U8G9veKob33Qvou/fVql3pGF1t6tESQSQn1LMg4Od89aKJDsC0JS
LJexxCcZOIMpb3IKAIXztrE0Fzh0RBGPTDnmEnq5hKC3OaMpUZchaTwr5dr1
g0+5MB/xUAZFuN+Xb5FAiyFgwHLZxa4fPEHr3oGYN+xHsxoqHDghm54Tzo1S
8ugGvAsfRYNkP9kQ5VU9mqb+kqupb/ooOkBJoXw49zEyEW2c4lbTlB5SYnoF
5aF1M0gnmGZ1ReTVPMmVJIgY1FRdl8z3RMAwtft81TE3F2BBKWD/Jt2kSVsk
iI9DLou/QjJZYKBusTfsNWyI83g5Em88NsqBb4+NVgrcMOOX438aFeZvTa5V
alaIgM20tPdA/Onlrt0yx2jPgdNQdceLlrlVmK9+rOv26lGQkzFHEeyEgcol
4+uLUm30BPw/1CvRtjK8/Xxr6fyTrKH8ykO8jG+dmmbZIk4bzxP390EJXhed
8VZvvsnNbwSKElEMcvPnAQceY4DwScT3LliS14UTVKsVQ9wz2wN9LYsFl8+k
s0acK4r9p7r0ilpYM9jE75Q+zPSW+zYRkaB5JbLP7hhqcPQCZKPusBGgEt2J
B8sZ3uvuEx19hhqIAb8wVB+a2bUyRXxSvALOTGvZ6TikEBzKbbemcepX5Ltp
ozQhX7cLdoC4WDX55CUWLmhwLQfFrLBL9uyTg0+Gr1I5vOYklV8waM4+4O7z
to3hcF8hnBh6SdAyVg/dVWpEiUVlLSGKH0iH0cLa13W5ahI64kQ4mC7Wlc2n
KCN1ntHXnvvVMbscdGT7tfTnDjTOvxxeKd0MUfTLm/zun9K4yw6gW8LUSU4V
vYd1Xv/Mejy+3IpTt6PLnlFI3nMLeiTFMkcGe5XR3/VhiaBUI3BAKds1KZTj
a9+UuosSaDKmDjAZmGIYVayEGiD7STx0r6zA8P9Sio2jaG0GYfazxJmJ0l2A
ajdrGCI3dqZIfRWHw2m45e9Nk/FrzsYM/9m0cQ3UKHrW/9H+jG6erQBhDEbK
6CiGnbA8XR+xsa/AwoM6KNqTJLe5Jz1Qk3n2HrwGMXE5Be/NQhUoZZDhb2Gw
OOrU4sglCYek0PbPGqHxL4u/I7CxRC51Y4gOBu4ka9L+g9/mrHcfFy+cJ6y/
jRVyNnQkCWJJMtaUAQWgTHTzFRMG6IKzcc5kOMDuM7ru26AWx1xwIcbhrDl2
NBLD5vgGLfr3bi1tlZmLMXql/eicJBZRvijAPmk0nOlOGr2k+MC+JqHspDmM
OqtoCmKgYqgZZHgcfWVliG+W9J+WQ2S/8T1LUZJSTqPe9HDufTiAeY2ydXb8
f/k0oGNwsw6N0gxCZ1d/KsXg7Lf8woU9a5ycvHo3FngmLfUryQC8CUNRy0LV
cWs4fVqgt6HlDdyg91q1CS9giFVlDq5fCiFFEBgO4CM4WbBkBoca26mccTGY
x1Jt5fejTp6q5ciOdvKJndVKjoEGEhGDdMWO4sbOvIWNi4Dk5uqItDt8DrLn
r6r+mV0mkSKM5oibADeVliPcLEiKR87pw1rxuWwBNrpKRItWUjdFtJIAvqt/
VAXr+5MJrD03JaCfZeQd/9HYynfwekpa3KoyopE2iDv8y4v2QkgDAwZhNVlR
KtFFYfIFD+j56I4zedLN8gZ+mNQ/AGpcrCFp1nl0X/L0YKSdLw0IIzMn8qMn
o86LIgawTVcm49PuVt0nBDKmk8PYb9aYhrmpD6pZmhDZ3VUEjAMhjrF5sP7+
gOhTXwuwHA13JzifSjoFPPoZzuFuN9dto8QcZcZNI9nTff3Zs+H31HkcOCD1
qVelbg4X+ozXHY2PMA4eRLCIW+n2LPUj6hfWMjSLGJzmkDapEQ37RXEl9nYJ
a0Gxz68NB2Ok1X4OnvVPKfgaLN/sIENElRQasONk/oEVPFveJZP8DbZaTn+y
1vcS8CG2bA/CGuMel189xBkwrrLV1XNfB9bwrFQB+iGHcVpn9SoHWbyGpxUi
j3YhwSvmeFiqiJ4mprQeZcGqtyLpmEdHFC+RbG8LJWQ2Mv3ECNrodZofBNDX
SaMbc6f2/2Eck26lTQsBE0g165vaK6rt2acILs+Uc6ATmcDWbOl0PCWx1OAS
XHeqPZuKUuZ2Rkwzxhyj04speNXBl+tvSLWvbgjz/Ot59N5217H/VocmEjpp
yAwaIjM/vlBo1Kdu12aGxtTXmFrUonQtVwqd3ybEohPx4g5dPcDeZ5//+5jd
vMWfqs4WiNiFCyMFhrNjVgr4JzsKi9NLIKdFWXEZnOugLsIbrg+a6kn7Hk+2
SDpzRbYL+j4Js8WVfGRG8lpJvk7aiqxu+g0j45VWYukgJ2uYAqWRd5J5xd77
EJ9yXOl3tsLwfWijv6ntr5UbYijYDZzqG8GxIUJtDql3npE56SQmyco7eqh5
oyaXjaDpSog5IeOwyFI5bprE+udFEY0FffJabtRQTZWZciIWdVoUFK644vlY
0cKfxFyogRnd6ccifjzClzndwCPGeR/6OXf9xrpcNng+ZOkpsVo4IKOEL8Ll
oKjm3N0oqz1sefyEo1CF4sjnQ/Hb/EBC8lUvJTs6QE8bsgfWj+Pq2lAjnMkx
treevgM2PRTKdYrn5RyFJ90i24BubU1eV14jk6dFwBn+N5LO7UQG5xcdXQiQ
0iYM5cpcmZPTXwQN+a9lGixaST0/HgVECjXQcuvxMD0e74/1xxBStcTx3NvG
kYYKrxYEJNwUJwVLrx6Z8/0cZIrw2ADTW1ox+Iwd9VD+nX9/RnlqukF+dixR
+isg55+0CJ3QQg2keYx+eKsGoXmmhg9SECP5ZxSL01oNpQUcPIXwFTV3yVtt
W5xbQhCKhubm9mJwkGqo9UChqkWEgc6FforWDlkwb1waAUAMjx5lkDoKT8o6
gQCrT4jCKs1VE4mBTdJ45VlOw5gHuHdfdGyds7DqQJ3/51i8GsK7B58kFead
h6CaqsH2YA4NuXGyR59nccgKvPCgaLUVPJ6wgr580Cr53ZEN8JXc0mFO2gvL
Sm5G49Q7y3vWXhlGYZqgD9OJWbueKg+KXkBsZ7e7BOxSJtsZ4yjDDG4UBHCP
+ygEgCrvWGKx0VZe7iM0MmihW6ewiEQiTsBoXb1g5uC9jKdFW4f1TZDikWRE
C4QUNA+kAcf+lq+wAca+ICDPR5IysKfTwYNiBhAwGtzxdDp22EJ6kWSe5YU/
EhAqKLqRBc0bZIsdAbWMs0TyvsMa/GpftIPNMIOL8iqM5XrZ0bafz8xmlaHU
l/0bJpb0USwVLptRu7GGXXkwRxGdOuiXp3TCgqqOUQ3s5PSgMdeTcb/Nuspn
jX0M4UZjj7/g7u2eLY0eMNEn115dXCwI3SxyhMGWi0ON4zhAJm+34jISGv3N
s6sY64ZzQII/OZcMQ2npKb5VsZyuHysoF7hCZfDGxVCFWg96Zym+vYcgnYB8
ziwG9bW8M+QKxIFPn3RViiJdMmHuLK4/WHFzXqKNEhgIuKmop7EJkTZXgGI2
/lPz/oP4+4GKHfTzgiET267Ty7GAIZycgmXbdisiihKaObwkOHHI0DEqKShd
XZAXwkqbsgbdSFVLu6COuxTxUzEH+VoMqbV0tox8jA54Cl0AFPyRTkI9mOiq
a0V66R3jy2qn2vOlytI12AIUE9NirEnRpjewV3TdLFT0gtN1cIfH8NAHwnLJ
UpkIxH5eO2ZIBbx1qtHYLuaazFz8rFjSoQNgfmDTLqqYb9cIsMGNYJWuzmvw
2GASpT/MY0IdkA+pMybpFuwkJxSbVxPxSYG5MvLGRGEyz7wdHWpNnPldb6it
fGwDun5N4RpqLkap0LXUaPctVWLd3VbUncb6dtTUnAyzmKaGkfl0w0L5rXGt
HTmUsGOAhE2q8Ox88brdG2cJ+lsW/FTdsE0xgVyhQSawyHgSyKMiojT11+v2
pmhAT3IjJBznIWqZKaNzLIYLmoz4HOQAqJTrx1rbZSMWOFKCrlj30p2psPK2
TNmXUBPxcbd1qak6ixW70ChbOSHVVHHmKVYn9F2STOYcxZEmRohYVR+PNxpp
Z+QGmasQLipHCihfV+SEb1NdraSqG0cIOtCqWoMwnCxGLg72ZXEex/+rv5Tr
24tVSMjHuKU6EYQPhxh8uCsIcDIxNc7+k58aY3tNJrygFhuSRgmZiah2WSTF
G3dfhcl3M8VSKOhf/m0nNCn95+zaBaJwi9Yglqk7RBU1p6OubgMS2z2Ias07
LBLMNttZw7j2371RwrgfuNK5o8YSSL5ods5OUN2cKvczf333nPGzrcK4cC1w
DgiZf2e8EIO4SLp8qmRxmktnrnX4h+kCpNIdeHbVrLjB5AdNptGOEMcbwCcP
CYmsRZ7kkIaRCN9BjC2h9HAWQz0pqIDtJ8shh/KUYO4sOqFhAG9kLd+7iGDc
L3cCdw4WXqg0Fku4fxksf+COMCxreoipo+ejr0q4m/ZvwBD/XqafgStc3vxr
VhXz7YLHsrqT5Boq5MCj1nlVokZ5XR552TNv7Y9DjdOeSmr4ngeAEnGw+LQN
nEqkxaJn6j5g8VX+ZBk95ytFqb5R0kWLOOMjYppR76zYlrwv8v53xk/Hq3P4
n2wGcKIddBXZccgSqaWMs/TGSYjGwkV+dGZdr4PwJiK1GplUkQBmfgh07uCU
mk7iJIIQDlyDlq+JZJtbI+ExlVcU6wXDep6JXQSg2xtkE4wwZLdunkmpyXPy
CsHQa7pl1wOY8Vjn3QcIgbATpYu2E+S3GDqZk7pxgu4MKW38sW5bFvh/JmHa
1I+f/pM9NSKKNF56lnGhT9VHdXaxCVwzkJWrh0mKnaFimHhQap23le9Atdq/
xBdlP1fbGZgP98OsPE+rg55UpOEaOjtmgNseuxALhLJsptUri+R97RTfdYSk
zcUedEt/i7YEO1MzjbxTcoWJXpzPezqrXsuN258rgrbLRybDeKxSiDxE0/Jr
JZN64A3Q5bTf9OkZJIDQm1FdID7HrmLx7dca/Tp0l97M7ssVsa7qBC/ye+VB
Owo/kTGGDWHZqbvR07xOLjN88jxEDpq76emPxjonZoTQ+ntQFA9XBzyIVei6
4XsHsr41jfTbqMWQzAhXbrTE7aaH59wT5qkm+CRs/qQipXYTsSJak+4C/zbM
bbUbg9jfkvpTAz/hzD/5OmKAWfimfDhuT5fZAzGGHPJW99qwPNqKeu7AHk+M
oprdnfuJSjAGTQS7sW46AwmclXtss9haf0E7bXUuljNw0PQ/0Ah0pnzNt0yi
QmixcxQ+GB+7lg6hu5vf5RawZUD588HfrXxX5Z1uOtTkPSknYpK55UFEisQq
YG0obTG3S9ZzP/YEY0VhXTCnhF1FXgZkcuedM0neoxeWwAacUh3sYugGLRNm
f5BO9OYzlDu7uepv8PDk6HejEKjHDlQqS6QNs29NkAhkah/VyLPg8eocw79s
DnNz/PdKMli9/ON/o5vdNUbd6G/9GCAnXiyfWbbzCgyihRtXgJwD+n9q5F1V
+btjdlp1eEK8s1LdEq6HaBLwmsY2dFJTbO1Xi+aGmz4hGNVtguSM/8Almat5
h1Mt50fvMIzhWUVrZwAPCcsJ2GOtfWd94mhqpwxJDFYrGCdFf2ngaoRC7l22
R5R5SEebJzvPeTdTcZF0QT6QLFxsa7AlS5MIYW8B4ZgGZz+zuUdSfRuT4La+
1iHf0sbOaQhMczThs4VPmW/y3cVS8LV75Nz6Ilpyk+v8ImKScBxvXTelDjrt
NEVGnWJm/mMXhTB3gOdE42+EeeWRjrBxzuBGpL/syR+y3o3pbpNWl7jnTVpU
kdDhJubVtH/A/LKpDTC07o5qlmh7hC41iNQELGVCIL44HNys94i0ntkHhX0t
dufICc5xh5IZMe56uFOsXnfFcblHb3YbFBm8hUELNl2AY3DLoQqXDcfeiqKH
KEteofvXiq8U9pqIpLIzE02x9Na/k3Svvg6FVEAKWAZdCGPdrmu/K05DdnR+
qjCJGL2MWpDyBU6LSsl/tn+qLy/4Ir+dQgjme0hn2D4/UehVleNiQHY0J+9x
MEjTXAzba7Wvbj9umvEmzoAVFaYewb6EwgNkgBE+20LyNucMi6bcG2JPDguL
mGdjmqs+u7VHZvDmHAJkB8/NC1m6/Xi7eKCu3AHb6WddK5CxH7hysqMaG9CB
DkVc7dslOKWfgMf1YuNqywPB5kKd6yoIA190kuqDjOtBYHix6Jgh39D+cSzk
43nbQFHH2if5pT0TeK++xWckOuAjZvpFOOwc/yR+g8MBvlNMnUz9H6zziKzK
1BfMMX5Iwym05lvZe2pR8f8jq92Xb2QWzVBDdqNP/FLsDbQ2Q1Kl9Vn9oS9+
zlFe/ms5SmPgV8DjIuVXTbvSbClgLx4X22MOX1kanQsh/exlOdgoirACqYGJ
axoosCJiH3w6+mGgKFmZ66qSFd2sCqyI4IuvvgWN7m6GeZeHRque4ZQJl5o6
ATEVdo0iBHqfRbBUhHje+33uZpEYIjF5Vr/pJlcgrekF2rheZ4P+gn4meKm/
UWZIkNTo1wMCYI80LoYlGoLGrmEDr2QGqt01F+XFmNhmE0f9K+NE+npIwd//
he4COfVfA2zEfXUff8afr6M0+o2zrI0ZnQRlySJGcSZSPmjwTOw5XV4stUOH
A1ui+37PtMLqa1cXwNUi7LDVt2UgZIp/kjgJQLI26IOR7Y12Ko2lRWGlfKhE
AtAqJQdf3V60mGYi3MPzxE4or2Vdl0C4xXGC6OLE51tmFYMAeOEOsKcKUhzk
OnPni0aNuc7x8BVppeWjGuLsuZYL+WXWgonrcqgZnN+JpTfdLZ9auAO7sNKX
AshdEUc7SOQgGerrSxsBOuskGkQjrQ585rym/EoAJ/p9ymCHFl5f60tqDGS8
KDF4VLb/oPC02rsq15v05UgJ+v5SdShDNBQUajiE5XmwLkr98/AoLDxFxk1v
ox4v31/AS2DPU4im7BHBmWcEc5hmFGXT1gcxnxEmNtq+3k2sicIyuOWH56/E
TYWaz8u9Oq+MavtKEmGjVIqUQhhKqVQfa2J/ljEzAbm702D9cLfHgmgTsfhA
nVm+irLGCyADhAUmz4MtISeXV5cchRDKwcn5RoHT+Pu7kO5JbFIpDwM2lBKi
xPL2pNhdHN/3vJHPy/G7lltZmVlET7BovI6qdaLDpJiQUFTO6vWyGWAlMzfB
ttBOojxvJcnSkXIMRcgNOB1Kmn965+DOnQxLbzXmbKz1rCW8Fp3C17tFbmrG
TzUta+DFKjKNHxmmW+s/l/JlYVIVKsu6CefjyUvZzITCBYsb16swfMie4Vu/
UTsvRLU4fSctP+/jLaY7yGxBKGyBPfYr06tyMGtPuqlSwkDFJMI+3/Hu9zkJ
Efppxp++UoY/sjvzdf3/Og3kCmFCgqTNoH4l+f7FYZFSuC6u7UG1GHzWWUOi
En3v/8wifDb++UzqWDlYxk3WWfZj/O/vqbgKiOkW3WFzBQV/OUZJ3GmZzfzw
7TJ3eRme7GETWzadIxKMQO+TCkbiX8kMLfs0fTLhPAVfiM67SWYFfMsEEn+S
2GpF5EZc5MlXVxZlbkqxjd2q+gr0Z53Rj6MuGP1oZLnrkBdFXxoSHgNKi0Iv
VvWCEND+XIvef2GlyLSuvgU3vfATc5AbbwKp/uO2e9haWQAiUIEzuMsq7k9t
JStS0eC6JVVEqB8KuH+Ufw6hon+4PPDR3hQdiU7yoauyvdpe5+obbew1DuAt
+ed4NQszysgFRbBTZS3bk1QbJt52/tqB5vABY1B/Q0RW12byhfV6o7xQvv7J
CY0lOo04HdKAcI9jptI8AS8bCkwoioay6amfubk1jNe3+3PE0F7d39NNhOAF
QFEyyx6WWDlTOR152oPQFycALA6XHhQeb+TRa9v1X5/EpExoLBQHQvEzMgSn
vijcKGMeBcofn9Ao6jaWs3Sj8opDC+zpiF3jRyBo9k0EACNF56JP1libdpn2
u2foPRyv7GBjQUmOAFmsjJiyDugmethhPHBuAUaUbhbVm02VeE4Fo0BwiHBL
EUc/48k5OEsPRt/92IdIlCtBW0AmUOeITieOKtJ+8+FpCnZfXhjFZxlTrtoq
6IqrWhhVCEgNqo1bFmriFnCRMpPay+2jKuMI1fryUGH4Sm0crxC7QqzrvM9f
SfSxH6l5tky62LsoSNlPvkrlaRY3uzkaYnjiJeywBXpEz4CBvCzd7/XSHPC/
XDD+MOiAPldEw+oOC4HiaSbhJuxBPv2Z6HyBWu5C4Dbc9FPmeROX2iYm9NwA
t2DNVTNkhgvBvNGQeNnZlJFgSrRqbOF5bePBLAKL2j/X6fCTG3opGk7RjAGd
nIu8lpeS/pfd//kq2YtnbNCN5fs8r4ElemPcuqBCnoMTPS7K8YVSErZ0WlsS
KDvwIL9rWoOGOquY3NmN3mNuY1KlwxFjCMteISvxiROTU4eUI2GleqKc/yv7
bQIuaTxAwXoZfXIsLx4fBy9CLdJFdxLZSB/BJ/J+9T3s4V4w0gvoazvAeND+
MmNVDOTZrvgtkaWKMA9ZnmwJ6RjpygtzOwcOzsIw8BtMw8UMdz+mB4msVyeF
AcygM8Nm1L0tTekiaGhhTPx0y5E6jsX2l4MoyAGMdW1AittgRHxu+zs3X9Z6
MJuJwEPTIYUGyTLVBBWr426YmTVBbIWUet9nBLtQtHZbWuZ2MsDfal4AIe87
55a7Ov5YYiSGo0kCeYCxAX4BNpk+OCtKrPhE7WMV08vBop2dWSjtkMDXQPd+
leXP6/Zi/Z0bHp4EcUwL+bg2zJH9RUh8JKhN1KtIyP/OxHPH6O+l81ecMHWK
ST+qrZL1HBrBWgXIuYVnleEGSGbCgSPUgakYiltzlixHR3yIH6MYA6YRjdY6
17nap7B6JUdjJDa0HuYQ8VnI+p1mLmdjKoJWQi79+ymVce54l0OkuET/Z4BK
XMLe0BlP4jSEN+ghwE75eYkyl5/E0JjH8f7RCOhm4doaJowNfXNeemgFFiBT
6cufWARKR2hdz83Ld6jLXKDRNElS0Wx6TmO4QmDnwDyDXuKKh33QdCHsacNs
wvLTNbLU26gnwFV//icpiJIbj//xYgpfpdeJM5dV+5sRl1AmJllnqQoGoVdH
2ZQgQesIFPhjBmeHIQ/ilSEwNfVVQMisoJVG1TeWm27WeyEuvfR8QABj5auC
2BCfQJSZW9CQlgsK8Wv9azuidENvHkJEZ374hbpcHmbxYCBYWjnSUBfndXPs
3QprrkXhuh35/WuVi1vIdz1bj20MKmEd+UfA1sh5TK0BBbpfxuJ2sO6hbp4A
NyWUaSCyw0QpYiqOEEDo4e88Xxft4aKShAy46YvVghnrSvlHKAjuGGtCb0l2
H1FocZU/9rhg96TbMm7+VckE1YZvxswug+2ladei2ktoikV/TTX8ve+qIL5n
ysI=

`pragma protect end_protected
