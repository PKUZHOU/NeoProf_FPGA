// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
RsxDDDA24DhlpsvYE2j/eVnOR/+slgnK1MamfB+Wvspczygsip4XI8iZhmE4wZ7s
zjlOnSL6U1udsibazdXDfaLubQwFvnLb10EhI5muNkQ3HLIBX3tsMptS9HprKyfK
KJvfsBnLzaB+LNVS32/2qHrFUzljl4QQRxwLwArgysqJsM7Ct3i6ug==
//pragma protect end_key_block
//pragma protect digest_block
zhHCIEKiPO5/cfs4P8EJl4Jfbyo=
//pragma protect end_digest_block
//pragma protect data_block
Gz+IjqIq2cxHQvTbHnbir6H3zgFxi5hLn0YSWKgFRnZrhAST/H7SlHBnib0SMWp6
I9/LA91usrEe4HCn2cemfQ0Q7InNvPW0uZ66Z1yv1LE7DxZJdp4urNjk4cL4NGw0
8xBRcumqFNYqR+KLNHlEhOE/CGLUysRQlg5S908F7Va7KU2UoJjWb5xNczN8F6Yo
GLLumtlcnc9QTJTZKYr1O4OW20JVrASmtvuzkay7xzn46X9i1zgrfpZU1PkxDAly
KiCIpSm5kdMdVx/rM2xYnaVay61zbgyUqPbHM9Hu2ma9GBpUdKsq+riqCmXfrZBe
nxFslpJHQQH/OJpHn4wDu77KX8D9r5+K+Ew8gtcwZRbofkbIwcYHhl3VG9+5uOvm
SWxPu9O/jlihk3nIoNGqPApX/30lQeVsxlFqYuhPTnVburHkxuPExfQUmSE5pQII
VacIgbm6GXO6YG8WzVaS7Po4/aC1WcB/orgQ7Ki4RqkHqwrKBwRv/oBW/69vGn4T
B63zAXw2POxR8lGaUQqJ+M7CP1ZzsC/NX2ef8Y1ar5l45X8IYt1dl0TCKHTQUW+P
XUKZP2m00rQh7sD3G6dMdyzXderzeiNMLRnDkKAYD5+EubPxqai386d1Cax4klQn
Ea4C8WUBPhVoakiR/mEfH7HOGPYEaiENBQb1P4MawRWWb5yN4OD5HCCLFvfitXvq
W02AFdB9YBq07jMSK+57cSAwzQ13qlpRDRNQCtul4M8hlVFNx0gRxZUsr9KGKUqX
gibNzbqwcXltMKWxgxSuYnWApw0HxJCrMelnQ9oM1GByWXw/AGfwY+J6Xh37UUCl
5z7UJnzZBHjzx3DALF451uGk8yPKQnH0XZhK7o3RBHG5Cufx/NbB3adGoEdvcyKD
CgHfDGOHwqACzTsjBxmYvRq+4zsVQrTk7VRCId/UISrROu8HVsQZMFtJ4E62/2my
CltELuo3jVKqkeSaV6MLcWAbhUKYjLm5Vqd9YzfxHQBnXbCbGqMAV/vJi6Pv9u+u
mSubuBp6gjhbcx6D/0Y7j5MhnTomKSPJpaZ7Rpnfeqln6cVmXUXlmLwmtsVlE0zz
rbU82iW60rspyJpZxl2S9B8hiA9Km192yuxDXFn1HPAL32sArAwEWTqzeS1ARLpZ
Jzr11fq/HjQV58YAqaVi7ai24fnOd+JoJIdj/PmUsI/QtxChuDTs3JSsUqSuflfk
Mb7UoBMLrJdydc7Q7ZhfIXflUqe1fHcKjsT5zd/u0HCBIoVLf455dW0PpLHZXAkt
srkddNHdmEv8f9CiY2X19l+3A5cnXOP/DHPu6uPUhs1HZW+kBe0iHOdFBnQfyVLa
bvPKU/chtvPJeAOXRcpQEWDpmS4ZHE9K0dvdduviDiU3Q/cHPqJx467zNEH2Fztg
8e5khgefy4z8mSYqnS87/YrBQoSBQynbaLdr6iF8IV5GD8DAhN/59/52tsXhYzxs
8EqzQzjqEVoIdaK3wRLozr+CYD+DuwLLA6uKsQeLMMDEskwmUtfOl1A9JM/xGATS
pBPThWFSGkytEPEIfhkxUbTj5dAWJLasquSzwE63twqoony4yLn5p+F7GVge17KN
T2ZkANqEtF4jcKP2sUTLvN97HitNEq0gGo2HNyYFIWnnCZj4tSmutRR8lqagUvaZ
FNMSltIEOWfWsc2MrvAfO++RVPCz3Hm0XxiaWri3xavzeCA5CAXldFEJm6FIWg8E
OJl/BduOsgOHZjjx0cWHfcHx0EpdIQ4yyMX84ggNNnsfY8l75iW932CgqLm+c4hB
Kz15aX5SBPskFYr3Zv1cPpuIAAPgDTcWeuCGP6Hp6ZzEJq4iowd6fZnO3+E9Txat
eqlKohmfZ382IOa6SrOCtVIkatisBIEU8A/5yvKzlHFG7TzEkKZ9bGjlf0aaRNlk
GKbUtns+u5JMeHS5OsBd3ORh1d/dAZXhFQsCVZJdbgfk5PhoWoaMakjEaTinLhfo
ZFKIqYl4BIUFnpM3D+YbpXyvxrLqxzhdsKbGlfdyR10LaD7nllymZpO+UCQNZY5S
n4czYleRPZOf0PbyqTXLU5NDq+QWZJAXLPY889XWFrWZ0i5bryAsIELWmjVjf/TQ
+UpswKc0omENIDvKROCrkphzYkJMcseCOYcdFoiATB5y1Rm+8GCnTfXRIBgz4RLG
K5HhuDq8rcGeKMKXqIIwuDz6jiRmm8G2Tl26aD0rl1IdCMzWNFnix8DrXOGFcUI/
VFClqWiDsS7g0PJPv9X161BY9NZNpvyiRCyaRDxieLOmLpYz99UOt+XNwu7Uc8Vj
W1C91UtRfBkZ+uREAjhkQK5c8ZpjBZlJvLpAKL78OKKQawJc5uKWtnRPd6A/gUEM
COTnKQ7kz4jxgVWnoV8Zynzj7X6dLBWr+Ur0XImo6ATGWydBtDWsqk6VgNypkAA/
r55hAHXYK0cvHw8mArxPo6pw+2HwY6WAmIytbHl+8oBgdmTajQa2xEJm4SZK3ajq
6kuSX4wI6xFSb9MZjkzLqRwIXfUB2K1E1CD26vlpZJU6gR8cGfknD6DPPzydtAKQ
hOweeLVNsyJupapyXA1tEIRZ1Ip/Ce/SVjE+mNNWHBCK/qWTY41vRi0dC9ahaqq0
8KoUoqtOcSmYHahFScij6ZpB+kg9f/myqffsXg31RemR8U+fA4kDnA4eV5wiCEes
38vPBo77bhZm0OqmCVS5XC9qePFXhk2U8ozSHA46nXPAZJDk3Lu4BUgMy9Hs75d2
DoQIfzXe+EnfOHFIO63yOdeOOCfCpcHwNnP4k46F78FnhI4aEUT6VfZr1PJhhpHX
8oeUNGJ7u2EVTmE2aHJgPIgeC8AbTPdVRo2FUszQO0aPlg4JRwx0usjGeh2g1db/
tdjgwBHy+F48E6gHeudoJ9DKOUoJYv/hN1zuswYtbmXgyDQ5xMO92BECGbXE/Rnw
02sU76oLS0vYCfpotT8UJaaSD4HMUA0VxkVlWdtLX0Vi5/tVwQZVo9PVb57jRxhD
uvS8HbaHsvo8hqwtRHDiOPNRF5ln7JEIKZmeGa7mM7PtL5n2xt62IfV0Lf/nUHVy
5P6bso290vncFdFRzZU/hI9yIgHeg+Re/glpzEC+jXm1LOjtSzutyHByozEnER4h
3Rwk9cJ8XHFgSMvL0QERGf377u0m23k3V6vw7ct5wjx4iqF6yYVvEXNtxfYWfrA/
7uz3TA1yWPoOkZ0HcAQIs3t9SEtA+X1QDlfdRrOmEfTRJDp9rA457ix5Ee+SCx5e
ikf1gMKyhWfz2PuZ8tMbzbkgFPuIL3QFYa8eV0uTINO9UBp49c/PT2t29rmAsgLE
0jEiZ9z4yrGq8a+2rEhCPIaFLR0C1re8q1UOkhzf7r220LHRjLx/FVWUt16gDkkR
Wu0HdQeoNk/JfNg+sE8/Ll3+DMNlVzdigoR1R9hNkKzcfzELgHxnUiBoLW1/r5xp
r5kWGPnnd7QjnUPUQYI7YF5UImfxWg60AtQ3XrxmEZEkD5NWHnIu6jzoJ0BGTQ70
AxHwBfHCu4lbICyMkl3nbik6wR4zr3XIgwI9atjYcxaMO9wSqP8bfvDMaGpL85yZ
Kb74GadbRQGlUW+SHWlLbgd8A9iFCyMpzkx/3cnl69Qin6rMK27befw9FESkGKvA
gMDCwAgYPYVAP8lJeGxkPw03d3wZ1GkC1b1Aa8LOAWjNCDh4Y3xmnSGTDKM3VyLn
x2n4/jyWPvon5b/sEWSag1XIVB0MqmRyJnwGvpU2Wm2YU4oFtoQu8FlHjq5IgeYL
+Zwur3g6RQ76tr6IdBI4Mj/VdOG2eEu4EW1sBOpfCIR+RwXffRffktLJm1NfbKmi
Sda2YlSwGf8TXciy8dbYgo9b8uSmPuKsS9VU76+vb/Js9p/0dbTh57BGApXPJEBZ
RDcFX7p5CKXDQs4ahd+KiLuY6T+f3jEI2IZvNFSHN7OLbzbXZCsSnuqWbw3ohF4/
1otZLXE4W/+fwyBcQzFCUTSq/WX7xvPQYYuxeO1SHnb6s9RyX2UwxqWESbSFgDSD
0SbNbdWOTMQ7HYeAv/jD45UPDwsIxfjq7or1Arhlc9KEStaD0wTGxmzoRC8k1EeU
90Xo/VdgQIiBhklriVBWr9vI2mHBkPSq+TeEVsNhmLKbt08A0AUTIAld4w0MbdNk
9uLApK53y5tQ5IKE5JiW4Wa1NwCwFtPZPOj9LvKZ+itZXajUOAbAq5fCdpgXeB92
3On1jabAmxVmGdxoCA3ENwV2QUOT3Jk7ch3V5SaSRtKB6eJa/McjnNJVz2/uwKjq
580A0w02Bte6J39S0iZBUakjrLc3aovnW9OV2OpUnc4O9ibxUweuwsYEaKRihsKB
JDLRy86O+HI8yDPsoTutiYXIpCOgI51WQj6rjSsGCob9di3KkxMKdOMoTYMgwtis
kKqmPAyqcIYgkAY4XSn4OM0BxWli4EUTe1N9YAXID09FT56EBkPEMj6T3FGVTF7w
yCMToHhyH+K6heTYDWZg3c08r9OeD8rL4g3qbjmVyTuJ2GvDhdL2r4R5ja2jVCPx
3/PHMy6V9bkBox7zlKBGuOUojktgdBYFFcdocWltKJqMrfAY0hhLRmNemF86YkBX
HRFmtWpIKfmxAJT3hSLaHRdgomMrR3AZy4drYJTZo+aCgar/fzQImr/mgVKDJBls
6tjHJnZaHqlrmHgQokQPiFioittjrPXoohfGylyBVLgh/j7uHgwMAqzJKd4PL+f7
QdlRnTjcjUYsMuXjaW+XQd3ZHGvE83VPwKvtw61Smz6pgdSs/fSOl78AsxtnGaDa
BD/P56cQAX25OaG2m55Tld/gI+e4S69i2nDXVVjMt3ncpzTi/0/NO4IKSlwZUHrF
8ghhycX/lbMBDx2ozheOjWfZ7Rh24DrV+XlPaA4CDoiZ7Ct6nLi8ObXSLc3rZXru
HpQwuRgu2j0/VWaPcjP3n0T6LVzVL9V16vycu5Q4wm736yONasGiETto4iJHR+vQ
Vg8qaZ5e+1CKKIqsRWkCR0WK1V6CLhMvIsFgsgZ0/917RUj+YxyCjBrlsJ6aFFic
NJSxE4uHRyEyvaFmhwvmwSqKxPE6C83HkZsQ0byBrASqqJqUBYbS4qsM3QvU5JKR
D08bfD487ArJV7w7ZU+kezcvrqr+3r/JbyqPN+XRefXtK0AskwIAGF3YWkHGGHka
O01ySOjxbJyMp2r/68USk4PQ7IblceZr4ABgYwAZBrN6leRopZ8Uap7k/foA+b9F
9qWa/Yk/bXTGc+Xt/QN8e83eV9GqTvbaFVR44a5JzzhqaIGneptHwBjj5S2g/X0p
QI4FuXdo6sx2acf+pmnxtZub2mDyjaYUaXXt0viFMNqy0FJd4sJvAhZTTdnpgeCZ
SlPiV9nrrV2T0OGtFYiZXR6vqXr0SF1/JvDggh3W9EXQEs+4yRa0JOYohtuTTldS
md7ULWelTIq49ftNrahIpxGMEKwIdfb5+1DcYpxfYF0QkqRIUMhQIUjGESjAwdst
x0DqnuPM5lLg2cL4PB3o+D3D3whQIXH3vBif0BbgTwLmd3mVbdhnf2MTYQ+pbz+z
lf5i4o1xKHSPLDoLn8HCry2WujYu7sB3Q6MvdQEWvVCeZGEyO9iA1lj/4JEKKJUo
UpQ2o5fOhGNoGhemw+Rm6g30KsIFFng+PMG3ltQqzoEUBEVbAhgMeK55O/txWxvZ
2AST9WqNWpZ2KKZN/3lG4ZKUNZeuAYlyyIwS7SiNLbdlePgxSXGLDG/pVD093vef
NkbzRQQNxFcdKd6nT8puYi+7PcdMBXOF6MwpZnPXL99Yq4MAjIL7sxdAVfsZabvx
0uq3+nhNWRTJaBCf+e00H7fOfj5V5CVlfdtdJTs6o6EjPVU2LCkTa92sEiiwABF1
FyDquiaiaKqJRkPLKQZZFgknwDcKExMPvVcJe8KsoLU4nvdDiakfrtV6DG4UG+e4
dhnAh37oX/Raz8aThdWQpCLOMfi2dAHSyWkDkGXeGNA+f1bSuagkJzPfWe4B+lFP
lKKqZRVpxululywtWuJS4KbUj0BNG7pw3SdxnH6sVu9CznIPNH8uLZdD1dp+mpMi
rtb4pSWc+J/jg1vNvgnB5x3SVJDaAqRTQSBNScxPI4Ic4YkkNeAqk2SwLyujk/H2
Xf0A0Rf3TM0iEkc5RLMO7vknWQKbg8ddsU78mt0t+43BmqsbJKtd48nCZNx3Sgyn
3b0gTdpYp/TlGa2IiBB4nn1wazAGAuzI+B6H96Y3AGHVc5OXRejduG7YeQ7Gaw5S
m/7NZTYjHqAKkPBh/LwGKIhVqDSYVC4zI6WYzmLaLWn/fl4KidmE+mUapl9W/ff2
d26cqbP+M1paV9h3T62io+CrU2tURWsgOWPtzLIgGL4ytxHncdZBsMzPRA6gUCxA
1pye3JI3sLT2/E+wTuYXNM04N2qPmTcCWnFGQYonjH4f3lT0kVDGJwl8c7orMXXK
+alKyEjzc+1DqPlh9YalOcdGihJ+bULFHwb930c7EuMnyYN8U6Gm2tb/SYx4ngQZ
SjBFtH8ZhUsqj1CePctAJkFgJqpzUQSJQcyvPQiG8Ec/TFlmKETe7WZSDoR19ezz
RVJ7Kh3gFSlU7bvkZwrg1JUPwHjPPc5HSy99n0aqDt4SU4bRX+Q83EHPVSi5++uX
rvhjlwz8c4Ser7p/S65MIY00ONk3p1AiSKRKl1qoJ02ph0jp+0aoPLvzoVUjKk1+
aM2z6LgzlxdtrUW4UPz52OwZ1/w9Mqch57DYQIdMrqQ10Yl6Ti35iqQTpXaziwc1
Cy4j7emPcoFPp37ALeSaWejADgcpEXGqtlq9Cgl2xQ4k3ytelAmz3n/TD68UuCXL
AtNZT7+xXCZLTwHc9/5i1ZMMFxjuE+Rw2F2fUwYdZRyXl203Qs8d1+g0OMLeCYdD
tbc7D1S6pA1UF2HLq3jT8nH5jzYDHtHPitE1BY+Rh28G14r20jZ8Pxt5lyVj5G8U
Siq5u9xMk2nBWyDvXCm4YluRJlk+52PPm2Bd79sHtKwlh6baUwupBr+6jSgxGK87
hCqmPKKd576Gi9opZfDv7M0is1pDDWkvTrLEfCV0xPcwL3QpL0aBZtfZ9bF5QCrn
h5TnQTZBySKtO2IHxGCTXCPVovJc3Z8y4gIec+tUpP0Hg5XUzv7IZ7DK/X/yRpN/
FKAWlp8zfnV6HR2a5mCvjGtpytrmZlQNd6LeW0/cwiZ3DdbBnyrrD0vP8Oz0R0O5
mXMsC1E4IgqyrUVEWrPS+clNno4VphTMmc31B6zGAKHO39RJ90D8lDqVyFQ2XvBz
qo+WJPPabM7pv8Iil3qLht24DsunkmzB1ZMRUi+AXQHocvnyOy8LRImkVEKAM+MD
F+uyGFqa8Qjl0unEDySO4ZCuLKIrFlk6zBCxKkLncGftJf1+q0G9zw6IrWjI8TtT
5NUe8yThXNKvqJXimivhvTaW3byR49Pm70DhBawJm+S6CEmS3n1W+3ujPhYK+Qox
jXLJZ9H6E8SBKfWJ+FEYlIRGa4uZejtLOQX50/kFsjgssHad9tODqjXz6DUZ753J
LdP5dbconvLZBOOfQg/ZoZSHrpe7SChb5f2/m40W008rMznc9Vj0Ebk+9h4APAVh
OKdIm5q+iP4en/sgZJl3QGar+l2mwL3eK/p15ROUnDj8XIsAo+/lX4AZHoGfAA59
7ikxjFzpx/sZMuB079+pTJKMgFHtOuJ9xU6RjsLT7Zj/DlG1L6OYu/XLv7haALU+
3iIheQE/p2WE5r72TcMTJ4HbTn2Jik5y/TK8TQsikViqo5tC/yISsgN+0YtxvAtV
loO5Kzi0iDBAcevY+d54tP4UynfL2XHQFpgOA56DoQuKEYmo8GZmnDvEEUF956O3
vDJedbt5ZqSuYZqrlFxKctrXAVVQ+qJK0ZVeobuu6AqKkIY3XFzkaE3PC+0EGSHB
NMokY60L4oEJkGsbq1u4G23pmw+NYenrsCqbpu+1StLaHyO/TT06jv7pmPYhxkTJ
tbYXyZUr6uS18kyEo+/FI7Ex3el/ouR00T8sL+psFm2R6ArRNugjgGWZ4rMRLckW
+miRGO4TP/fNz3eGptnIGOvBFXFItQhRc+kyK6L2MU58+YOPTpoCKMsxJlnhF8Oy
7DbbBr6+zIMGkWBIyCc/8WI4iagc8xY+vhp8FAPIqYeq0w9WzetpISMFV1u+gP9F
MSC0ngqBZRLXtV/mDBUtz3rx3gI4jFfP+eyrOpzB1RlrQ0Yi4teho6ZizoulO4UK
0HdtkwMRD/YGuEXlbnja0W5Nm50y/LGhjvPJTfLdEscw4jVkT+R9Wr5lQRZRbB5d
tgF25wK1J5gxyobkxShThtR/s0FhcVZBVbxMzTTiMVcPC/zlUU2tfIiSt/yIkeUq
O3W0KwfMxnjIca9HbKjMbFVPxzW2iWTI6jys+/OvaAf4mASdnS1Dah+y2aeecP/E
VyKPTyFFaoqvOdbvViUym4KLtTfMkby3t2IVWQXVAlZTaa/vUAWo0dRHYeXOWfuc
dSMO1F3aPd0DnesAqe1ZW51UKS/CGUo2M2vJw4izaX+9joktgSxCKOBgm7rjJTBy
4Ip8usSRvwaR5Jp+JmwXGW63IF5P2UCwf8fe6YcGGnIq7PZUgUaY3OnT2r+sS6Ds
WCuqlCPUaW9u+LC2lAyqSWQLqnifAfJC8eZUzXW/5iv9dRsGqgOWm5UX4OAI2I7s
IKAEujrImzwzWVgCA0uKSTxYOaO0eIaUNDXTaISv6M+h3pqrTo3fIYhBCWt2aFRD
XhJPg+q2KGw/1fdF9ddzfKiFr3hZmChTaEllQZF73zkvJR11dz8+OkpYGj4wyU/v
8c+HgVDkfg7ZebqNnYVV1fFyoV/RhqkgnjZbDXFldDlxCV37XxK2luXTBA3O6xfN
cGpc51CzoVRq5hBRAiXfg2zYLc5BvCrgr4H1Vkuddfl++PODH5NnWcJk0aKI1brK
D97+MYRqdiE6d3XyCFKlhYPbia0GyjEFaJl4iG3xuZp5lpei6sTlgvLp8l8EpSwU
Ts7mMwRFSP2ptMokIy9O8IYfu0G04tgX0i7l8AXn16eUEp3gl116MSXdbaab+SGY
WYiFDWUsH1Hb24uvd1odOndgEY/PyefBFXVJK7o8ymAvzALejLpVcPtkl4TkKOGF
1T3qHbNBuYUmUOjAX0ojSFJDW1qXbzXAMntpWwvgvOOlu42k1jItg8Vi3Vbc7iSa
R2zgj4PYCpGONWG2ce+DIwzLziRC91XQo2JCjq3f+qYqPzpgPJOs+XcbaR6CVPnu
1Gg1AwJ+bFB4oXZkz5icEi4rwdR7juWt1h72kxxMkGCS/Zk28HXJCelvfdMgj8qy
70mgXJUJyzFBrHpeWHLQ8ppp8xqt5zMO3FbNt6LBg7qGRZmGJmTXNoxoVD59Un2m
z9Zb81JM9XZNxqj9E4gmNDZsO4mD+FRLz6afdwoQlth9uHoS3w60CmnN9mriAISn
TEbWAatwkDB2nPv28+uXuMzg8oRzECNLu1xTSlgulGpD0WmtHs/bMYghkBF65g5V
oAku9Umh6924Z69V282/AFuqaZ/6YAIkhLRYYGrMd2HoPmiYnDI/3NXu+uBgeUrD
xzNlxA0pvpD4dtNqzkc9zogUlZ8CBgXShpUhzCsh7PIX7VDifM8pi/HXNtcY+poV
RupHvwrScUl6pjhBBQCGzVc+aFAodG8zcbJ/jYLdo+CDuRx8p6R70EtagXNbgUz3
iLeXYUoEST5ws44I73EevEaVMvi6WrmG0iACoo4OUr16CLx8wQXKFZBtmhfXF3wF
DrmH1bS1yJL887WCeoVjjSHDOkDP3H/GZsyjF8xLqgA8d8rxArWWxsCrjXNjf0uI
DDPsiJ980YM21F4y1gaHKk9IUTdzaCOEIgwJbqCWAQPeCvAvHFyF7SpNJJXxHsdu
KuurNAkdECxgO5CaOq2gshjq8pMHCfldqlWJTclOiSkR3OcyQ0FX4ZyErnmPlACu
H4Lx+Sv8f7ncRexomK+9f8YmLs00PMHM1TMlvFZoEbd7/NypDd6hsSnSfR/7EFHh
LNMiG0LPEXmly88zurgoSlrmQqWuQ+I5BwrHlQM2A0QrKmOzKJQK3ynsS8MmCDGG
GXzeyzwq5cI26tB2T7U0/FY7CQzvDGfriGUcbGAlJcxzB5xEVTKfRLBGWN6KxrMh
RqE7CB7T0eBH2eK/sictYwr3Gvvb+hxSX/QSd6wVnDCDRjNEMYruEAUBs8rq0GBR
SmD8DDyTW0voMbLd9IR/NWDKioxEa/9aR/OLd+6Rq3AKhpJ5+EuoIv2dEPHE7nbb
bSw3E1CwVVQ5IEE+kT787F81eUOluxLOjmHL7JT28vA4uWw0WWNwKQMvWCYsPUCv
8kjAF54T6tAD7eJLOxrplug4alaM7jcLdguEyzE+uTAQL39I52kmLJv15mtIPgdw
7/mL1TubRcjAV8peEpxt9oa7bk3iUmQSqSpEm4nOKEmIUAnuQuprzOllejvaibWA
2mhiHzGDs6sgYmRH3xHTLsPsKY0J2Op7kOfRs7o2T8Tt5mzcIGbEGaUGX81Fg5Np
aG7HCgkIexNQ8n/fROWvOTbe77MdxDQdUDOCiqbn/emvJyLm8t1EEIWiptPo+daX
xXYkD6X0HwDlQKsO9SaO/RgH1NHZ+9HGYii07e+8cZZ3gb4t35j9qNQfUBVvnheq
v5uL1I4RhXF+Hu/hyRmY1V4qClUS3C+EZ8smxTsqCSYcQH8I8Ctr3Wn2gOMkTt9l
op4jWwxP+TbgtUjA/BMtfXABzkKdEbW8SJ/nEm8x5WfoN4RqPu2KDAKYJAV+k9xc
vdo47818epR02MHkjGbQgvXqqMv1XdFNCDHnVdwsvDrh42bP3wKaMninHAw1owRv
iOIUbKTA+REs+kvQ1CtoIOU7xYq4qg6D0DMkDCTgjCLcfD8oZYUUk95bH+4qayWh
eTWAaJP3AnvBSiLaIHx7G26ea3VGUb1smzc/UzDEdJ4xPRhVPVFrVPTY7hi/bZSX
8Ddh20CrnPgl6esMkJtK1//Ehw53cvQDtp/yMZnPzFVygUdoRrSoZEg5XZsjk7Mn
kB7JHKFXZ3vDd4psySHqfNdtNjipUJ3vl5PdCaY47XSDGLulAMykRTj0RFn2c1MY
pp0wfz6VzIxzwwtdzUimwAvV8mMnKGlBsS3568ATeU/mbzQawIb9ZhUBx+PRWZy+
1pCuJTWxjYeJJjSmtGa3gO212hr2pDPTXITerB8/Q4gtqibqHZz4z19lzYe0Gdyd
vk1v7PhnVsYDo+e0rr5FAtcwa9ouS+ibMJG2I9f2GHl08oLmP9RaveiqzPbUZcMF
oaWCI9Qe67pshDGzr9ygZK5OKfrYYpwP3GZ0TQlobbBHP9XYTnrJfgTLhbt3t7Ru
/Y+DZNroTga+l1y82KujNWFQJddGm8DYQm343Im6t6JnJPPZhQWkTN6pFS+Qx4LA
hLQ1PcNxCNpmjuGlsc6dXMpjNWRlcN4YVBrjG2E7socuUT31I2m8aAH7ic1f9/Jx
uX+i31XBSRTR/z85WvhOadHF9D+Ty0EmSjTl2HXrnDT8OmZik0S1/Zfv3DddEXVk

//pragma protect end_data_block
//pragma protect digest_block
wG0hfWN7rB4yaFhzI0dCupg8pAQ=
//pragma protect end_digest_block
//pragma protect end_protected
