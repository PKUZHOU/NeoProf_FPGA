// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
fnk4Z1ZvrxDJIl7hi/VK+tmeyz8RMGosFtUJqhyxxZfJVMwu6S40UYWFmxeXawbGOXUg/iGOr8L3
X/OP7AZYUTRjv9TnAFfRxvn+ieCjBk4mHJV1VK3rzJcL4JAYlYdwipOTYvlXLtSvoHTDQmM0UIi/
ZNlgFk7egUiz3gp+zJf8HJY/2El9rfRMwpYForfmi5bI3GeYUaXOs+jGDBGN1a8RUXbOzu8lbiqx
VwKpHY9F0J2+czkQnCeOr8ux06hRmcB2z26hZcYMXXXyUHI37QlkPYOw6myxVJiGptZe+X77qT4x
hC4icsocCzygFAxA+Ujfv1vsgJdU/GERM2Qfww==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8496)
CFxVDCzm92yMz+N0gDqcI+YJXqPN93m1keYN79+XlgCs0iUOjjQAhCVnYRCfFmQXozqjhEp0fGQv
zuYs+FDZCRDpGTvqYd2r79TwvV5xQQEtbafK+SDFMHPrm92DrJZ7Td2EXImwp0fb+EAg79t2X2sS
W+m1imY1UTPHo5BMnbMjQ4mhpkJuTTkhBFIw6u+HFR2Kyx7FZGISplBJfj9brhgA0Ziv2mEP7ryl
/2Lb4wKIZW1UiSWJhjbd0VDqnrZyKgf23Z9SGkogAk+rQiEUH7vjzxqO4Aikj9ttKvLUeG4gRvlP
dpnuqdFGVvC40RgvEK0g4VsxT4Ypalaj4/eSLRu/8bfs1xXEgW90Dm1f9U+XusyaOvT5nYLINgSe
9QJ9NHkjNjjX3jSAjf+pV3zYi5pTVOhm2BwKQ35CwARfpK5sXpIxFZp0YGHtA+BHTdpU8Q5kdxcq
dGBlhxoOl9tuSKUuusN2v5XzoOhJB1tewJjP0XQTQTMAmrbtB69LhydGyaY2a2BZ8GJoM2MttVzW
18YfoAJo5Oy+56zbjs9g76k0uzgDOpDFP57QkTC0fi3PJUoUgoB5585rPWx8m586SoYIANAeI4W1
eRHu463DXbFOqt8LdfvRMQx3gGaGalli96quGMqvX+OJLy3gbKss8Mr+kzVEqGrek+pS4oRczzHT
Rif/4E9U3x45sWH2vDlCtfJWthEtpPA75G/4icCmOtzrdbMl5RVosy7kgs+JWn27DWnya+C6+izZ
sike/k4sOjilsDp/yOJVxhZD5BIQ1dSNux7YaI+VJLPC9qKPtUatBznzHQF2K+ZVG80VVU88TCsD
ZDgRkLA9+pJ93qUz+jXztnLlZgpfpCD7wE3sVOhyoyzlwxIgs2+6T1muygW2ehBjD/g94mot6193
qCqB9AWzhOWW95EfWj6cgLVZs4XI/SG2ILoxw7rXAsZ6BdkO8zLU55LCyeocfoojyMBNuGIcVIG+
7sz/3FG9IDjmUkKCL/kH7UgTaqpLO2zzL2qwTlhhMrkZYGXDxv/AHBA1dB4aK5eGAvZFgXu0jrBU
RbF4UY7mwVESiKbzvV4Za6Uj4dueAz0RcHDsvypnUaztTpK+vcqRaPrd3/Wp0m/33Cq1/MblL0MC
Lfgioke4ecBbi+bRLFIuu3ZiXe5Y+310aS36xC1x4jA9+cbXLnIRHcLYl061V0WI8xlGdVjZyaG8
wsd1aKTDiFsmgUPW8lHgyODia2P40TWpL7tHyoaxTvgl/YZ5ldGgq0KfCvrOoreqecCdkpq9Z/Jc
JDdQRUfBYvgKD1Joscz4NrrysNRc6KqLWYBV/tqPeSkc3razeSZn5HWrUGS1kdUqpTtj2oNo5csd
ZsXYlGnUIk7iI8N4q2I/F0BpAumPJzqePWygBlzJ1fgTccoPgBBiKUsqfLIAldrqz8GQmHb0jxDF
sQARqrYGFhpILNkRrRqCfcIvfzCQYHxtd71ve8GZuU0U80/tVvPNElruGOuzwoOZjsm9E67JkDka
bGgEFc2VJJvi+fefYgSgSVmum8dDmUW1kBtARaBQP8rvlNHCTamDgIUNYvwSAaxuujXFAlFaItb+
Xdo+yhh+us9j3tCkF16TvqbQ6KTMmKqTclnP+wSDRrXmp4rldOsKIIIJDRPdy35Xzh8YiDungX3L
jvG3bYdKY+kTDDKyyvpIh5hKmVQdJrihbWPCJPmAEhAgQ763eWAXGmdRtAD/e/mngO7c3/5HTuLa
jN61aWhgAs3DefOPNjlGOZ4pG8VQIfV6lh1YHtpSSyrriPjixYf7FVXmN42VKzXdHwUUoKleOpUU
RXNznv/qU7CDjqMcGJx2daUxycDpEmgyepaS3HOX5rcCZWeAtGP2HQb8ssAzqsJ3AwBxhV+UNR7K
nrDGWiCrFHQTZlQcon3Vk/dfLmH2trZXWj5cMJfBBRJfjSJQhjmWDuBS11uawxC6rWHIXAoiwYgb
zG9+qipRjO8LLpqPF05JyYwReQ2O0i65HIGTSogIuzJf7esy/EcL5f/aIyufOcxJ0YlKv5hKI03k
rCNg8O4ofiZr+b6vXcFcWnb4MP5+817C1zykeWu1UgjeqBH5cWMjXkzmEEqFreusUcyYT2WkAIA/
eYUrh26bm7nWuE1TtRh1D12QjMzYoFYRxDexRBHBHo75KORRgZ2vVB5c0jjHsl5jY55kR7kFCrCf
cf+qUouGvo8gg82kv53pcNbYEC206qbDpWEXwQ++SQds+fEcNRoq8rLBNm3wCdeG7KsFDtsC8n4f
cv40TRyVUFkhFQXMTkGBhb5BwxplFsAlkD/VDfc9LznFabjKIdat43zA5YV/TWU+7ExwnTpOQmsq
DcyefQHa2tEIYbGZSgj6MU7mtbg4A1FOWIQ2F6bTm/Cdw0jDAlH5US720yTU7gU2ySpCrPEb+g8+
+IIyqW4tSG1weu3FjUN5T5f3C1WlMCN35flC8GcOELvy/3Ij6iS0d8n57Cmj7cIf6QZQ2dOpvpnG
XfZLqEm9EaVgny+f6vM8PknQTxP1umwy1aZSicPRCs146QJxK1ZNsifjC6WAK1iwiaDuxmbsNdun
aAU1HPfXR/Ox2J2p9uHdGn1JsSQ2TsidrT9G8z1ipTxLinVeIfDMKZaZ/pnXP+QyzQOMvcKy++ky
CkOHN7fVuhCPS3x4Mww+hTUQR5gPMg9JUtCyFGTVsGShBl+XzPlU9uhAk2yLHITytgXSL0ynfhaC
Ywg45Hc5T+cp5kRiypbk7m/n1IPAX72uL7yeuJWzz/O3cleb/3j/fORlaBksPycbpCkgndo4sCi/
iQSEroMvGSA9CAprHjX/8mJaIu9FZwll4XH9bLPhRPgc+DeVbTnXaVcUoXCwsArsRNPeLO+SjwbA
rS/2DMF3TxeTpzANf2g/lH53xNfPd/NvMi+y7GB92vsRn9RPnc0ncIdxGh+Ofm6dB+tJmdJHIjnC
EVnD+so4StHxh8QwK0k5kSqeMY415ILEjo+pSlUxK63t+keLKScxS3tLCrvBs+Xub0YtdK68f9KL
LUyP4YYr08i1G3iLUVnS2yE5SeKbTcbIk8oYejOEyP7ijEOjU616NjtpI5XSiy3XQ8tMXsfcgTBE
fjpOjq/Mc+n3Oc1UAUQ/dPjYN+ndcF1rjPx2xhTGpW9rqOQlyQcb6SMLr/6sVeYXopnNnpQYRfrY
hGtm+374LGbOk7np1QL1M3bdIL2PVVGC9a1qtb9wvIzRAI8JvOY9TRa7xNWFTetpPXu4eewvw8CA
ot9+4ERGwa3/gGsQPvKMU9NmqHXTpFad9dpmwWJVcdgm64Psz48Bb7kB77nJlWPZ3VAR7L439mjm
k84wIrd5o1MunfUVZ1X3Yoam5QpeKBhZTt1eB+8WFKRYYFDDAnG9Me+MPW1CoL/Y2lhjtDjuyn5x
QdI2Wksk6/I/tjB8VtIfi3MsJNgB6K7yQjng7LULpcgeEEbHmN3JxGRBS5z79Oe9vpQ9BEiG1LlR
WejQfHJPjm8uZOtdYTt5hsfzfl9K5jsglWhvB507jMqVBqE94BYImG2Lj+hkW3HjmIgFHhXwY/UJ
c/G9S9ck66q0HGCXwA8ycLY0aRAZ9kEjd+OW6t4e/Zytify4si4KlSN12L13DU7vCnCq1nt9vuXg
cQIWvYY02PyCHrq5dRyrTBgNju9nacnDtUVgFanMx2X9Evuh02OwHq8AeKsx3uXtNvQgWuleDHX6
sE8SjtWcNQBgEnDUjkO/FEMuIemaPFCUwXtQasP+FjQeP7szNjjjjREeTd5ptiFC9IEhZ5wzSzMD
bwokMCaZu22sOhDr/JIytaXPjCOmfVphm++mWQXRe+HUGLrsaIBdrdO0md7pl9H/QWJkICQ2ol+p
lw+YMhnTcJva9Q1VMls6WxR9JLuog78ZcEGIJ6Td6foo0JonZKTUIi/uI6ZKXFD3R8sJNhOuSFu5
aulFh7Fi9NHIVSBFUyKpwJ2qPHF33X+WezunwiOKKX+yzwiYdcz/hCc/IT7PIiiOVf+eCblppIQy
Ze/vvjHL1Po1n51IiCB21Ppv3E0/1cUisvyM2sZ2C8O0k1VPk14j5SaVFgilsL0E4n7BWPCrwjUw
ho0nuHoOcKZ92+eOL8WR2EjUs4gbHMpGuayyq8nsqEaCIMp4nqAO7FLxhNP9wOihzB3d+wwWDgCB
6HYQI8VRzOyA5olZG4Met5wNaRUC+ITAejg0VUD7z7QicrMbYp+aLDGF/j9QBPmzjaidIfr4q1Pi
UogsM3RyI/BmTGUikOolhbe2oek2TOXO+Et3Ov5vDStJDPoVNdzeum9T7BubfM5N0svSPJPOBQfz
iolJH834+umdlqgihawK9ctemgXVs1K+AJMdoIf+EEGarWiNN1LNx1IUIeMJADzCHZ9kW6aQQ3Zi
FnIs6uFFMk6uNGxAMuP3UoCS1mzacuPFhbwBBud+AQmEB/wbirDpErAJ1S6zNy+nRELdfoAe7djW
YePktJ1sP0v64E+U2v8F8NS6Y5TiVRHu0PhlwFriMNei2aaIozDwArdaO3fZg4htjNB2GdA+CS3f
eJis8coAw28PnYDHw7t2Er5eJ4DR1ydFDJ70QeIhNuNIEFZqVWPJBZStGv1owuL3MBOroOmdQ+4E
z87uo4uFqQHZvVvYR08QcjbCF/znMQN/A2eCI9ihnE3UqPTGMJ+lhWlgiLvOcAXC0rTgd3/4pSej
cgdW+RvQuhS4PuTQei+uHxFZPE+yTMpoxJ05ILtL6bm0GMSmZKj3sTuil37Qx5ZPADHjUMB1IcRX
E3Bmu7+YNRU0clRAvSjt08IdVZigzAi/iKWTlILVULfIgwxhaY1qSaCn4G6K95stacx9JYAKkRe6
S9i297Yaai0drjIxgsOaZSJ/QdDYB+yZxd88wxOJe1cK8r+pRiEJNV2aj5ni8wP2SVK+B5qYFaSZ
69LVioNMTq0ymzAPjqjdtEr7St/8fvqRzejA0nYpR19LWJTLKnkbFHbb4mBg6dZQscu6g218C2oY
6dDbm6F6k9bG8J4w8SCygMDlNOzY5crjMfqywYNBe2tCMiash6+DQt6u4Nh5MsCt8mjXuTGPpN//
J9Vc200kLxPboBXqx/2vNXbzIbcBJPRR56XyB+vl/lKVtRZV5UJgN7wu+6V+XPq0outpkSeczADY
OdRJSG8nLgIjpbEp8kadXtZvHXIhKT8VnXdXQVpv/N/pJ5NPdpo/eS1UekYsGYBajo5R5Grjfyfj
aSgSszL1xxRRmZN3li9iwu9WKzrELYD9vAPd9J8rKep7G/eNxYfsd9ap2AyjfVB20Sbi8x/ox+Ht
zk2wqJBawx2lz4Fr1h0GPhUFYbZNqwHHQRRIRghUylY1v/irCPuXCvwTWr6OP2v/u3uhNa1qTkk8
20waPcRrJhW7wrYpZ0ag+LfmGim1Oxeppb2w/l42lwglvXAOG1P7XqXfhzQJbCrgegpYWTubM0p2
9kqsO3n0bVHAkANWluxNN7AQ1sa6JDPo9ivCxlOoJzXDWj5YRvfjAOk1djBDo2XwuDFEvmJh8P1S
8Amo7aET7amna+93WqW/new39VI2SdklCU8LZ92qqINdWGCxmMW/Ab/EsCl0BuvpW0sYt7BYXGAT
lcEsjAKJQgF5lDr8XKb3x/F8fmwGelz2Tfn8hbsQAbfYhSi79idAAsFnYQ7I0xkCJrhOUhE3Yqrd
j9c1Nkq2rn4gvWHS60nOz/Jiw5tYdiL560U0r67e5ZyGjPj9lbFjEqdiZHkprwxoNu4gOAyyc6ee
RJXb7H5gaLQjIzDUswGGe2oUQi5n3Usb7bQPRMXryG8jMYOl6Rly1+yxy1cZmKX7uchjZ3dYd1a9
8QMKvWUxWrYa6ctbRypggIct69F/RQD35a9Hr8WDp9GpbSdKrNtbgm/9SCaSh+juydeK8hfnFdqQ
UDGWPbfLfeYMPkAOC1Pv6jhsKD3ZRNlRmNgtVF7Gibau92j5mgB9csom52BrqLpYQUQNxkBFYCsa
Lwq0XUeWe26xGFH2uNt/UpWAYm/TcdyP0J1fnzOw1E/XM8opC4OZ6L0rAc8+eJcAK7UvH7HgwlY4
4IOWc6tndxWicsi07lJxzNzCGbxGR3YhRnRy3IpHuTjtBLSYkTbQXQF6iObV9mm9wbLo3FKjOypS
gLdqNkpyyFU7MzVs0Xgcdeenf1WUlLSsveYNtEsy1D0tlEfalw2SGdrVf4kGFZkrge86WSvKKOKx
9/ExEQ4w5BHg3PPtr7Ld8TpJjO1FYneK0f0aFcNduAXxYc/WnB89ZeN+wT8bwlYgVBJFdaBGJVXB
01P3rjhyGGXCuyjIOmQoSt6nV4qMsn+U2dLIthX7oovRq809f55CFbK0hA8MWLnh+5sHZmS192Ca
dGxJyZu2yArXQ2M8T7sblNqOG50sv/9xpKGImGgbbBLixRJ56Z7M+294opA9GHw0tBaUlqcCHjSH
LjlS5R/gmYjQ1wByrsQcl06F7S4V7JfY2ppP9jU8t8zEb9qhyyB+2r01wFEDVFR0ARJItp0Prgli
oe0AfNdK4hW8p2vcH+JpvlKG3os+xFnLGJ2/fSFq9gjQobdqhFUND8lDOUMUKwzoIVF8cS6QKQZc
I7i8Q33simOIRk81y322iK6NShE/+lkzcPTdjpIn4CbaA+4tbij+lCU6Cffe/Dinq68rw2GZsL/i
jum6qqPgzFeJe50fX3tD9QEBZ+ZVrHGY6aSbzTT54tHmnSatDSBsiQedkGeAfq679jaCqrZL/5oD
keWF0RjvyyCjBCMc2+Em1ThDcjK4NGGWFSgs4Ic89dplkCR1YXVO3Mqt/pN7/+nNBdxpAS7e7Xxg
tmBFwDfuqdsu5WkMQ1fBpNyEw+DiDjUUk43vgYzklkGI15XSJWPBvnATauRsm6AVy5kacSRxbJTU
tS5wpHkD/vWDs3GaRJSq5tglBPpXL5i3zfdcSf3Sxmoc2dSEl8UxnELeR+J1+GdWJWf8liuGQfbT
auE7PWaRoi6k++/ZdVCSGevAoA1lRPv2kKdXUSh264SrxGenswoEWABvALU9Pw8xNqiGENZthSQ3
sPJ6ahRhj3lrKftdMRMQc1tHhRL7KEBIIAy8rVYes8Excz1Z+CMFDPiTLI1Sa36thnhPvg6di73t
qF9rz94+eltZhT5VUbKMzow43WRUw7zrbl7HX0sg3X2RKhL0t8V313XGnjNCZVEWkart6VmH7ifu
gy8lIwlZ5T4VH8sq4Mg/k6m3ZkV4wjvq6B5kKwDJjVVeYGjZMozEjsim0GZ9/qM6RBPHwurIQfNZ
5J2O3/w0tpZ1Lzwgfr3nadTm+p2I9Pq81VjprPbHyQB+gWbuIUA2mGdNJDgIA+SB3u3hLjmr5ESV
UPS57Ikb0v0TMCq3Z5dwj7D7DV8cAnYMboB3/8AurSwFqBmouEkMsjgdZWYV+wQDvM+q1y5TvoM0
E1JQp++j5dc8v4u8ZMpMQNPdtyTHBquc3DHElVOoBq6KFjLOpeM6BX2mjNvRjdeTtSh3VIfuee1c
L3EG7UC/UAlbW817s2bwc2IsKJ1gdxGOW38C/i3kfFF8tJU5kSfWu//FZtCF9oacq/PnSOxE3N0T
x8v0VBdzZWoH1j0BqugxnzPY7R4XIivrV+u75PBuzmLFZ5Xd9PPK08pIp6HSLZjqTfoTtZV3la0C
5YGO/jOA8In3QPSj7DEn7QiteOm9FzQFK95tnDOex6ltygD6H4f88XCmqGipuzTOnXpbApW96vAi
vE/rK0b1PdWAu0hRnxx/NvkmlYdWmFXjCH8jothz0j+WiFuTGqg5sdF9L36cRn0ZxlI9benuMp4Z
FGGb+nkKSheaDdnv2IPnb+/vHfE7ApSVhASRor+cXXjxcDogWgVMqrzp0FLAc+7rNAgnQ0M5nNjs
KLDIfSWQKvibGr0tkWDLipyPW9hQus0H4BjIbH11bWC67Pyn1g2288zQeH7kM32UuecZTtOuyWsw
MI4fig1QpqoAf8dl72eCBKw0zknVmWdkDzfT/5cVZaPxVwVNiFmUqMVc6iLYdzT/DN1WJIkrxpxz
uMwnmtUs6rhmckz9iRQtycavBh7o9zLJ5LZ4UHQ4jQWql98/q7+Kd5FN3cbiSCDWafe73g91zvgI
WSP3myh/P6+tREULAqt+qhk7w1cvxjVkE4uIvsZp3RqJhQJhNGcGP9LNqK3LyvAgpjv1uC2/yoKB
TENaC+fouwukqgKCBF7RnuK7FRj+hnjjUClxNTPXJ6pW1a8AASUfbEwgcTUwqBELUV6St8md2ZCc
/AklqJemIclFZm1MtIlipQCgZhElRSjtRcQv/dou2pwMk40PF0nN6IYKFXzlRxgiBMQjT+LMoFEu
ADx68h3n58vlL9xMkungxFP3z/L+r6cp1xF6O5vcW0hzMncwO8c/cW8ctnANMnnV2178YR8UK5q7
ilsIJWRUoGpXuXzQEsjWdUtg7mXNKI/8piO8miKtrkWUW1V+ejUuyXMGiASs08aPSHsQdWp2zdbU
5Lez4cztNxGOgty0NWta6cu2rBQE6CyVxDYEu+HvPp+1OeJmedr+V+Vd0t2DoWARzZgCpAGFn1wC
/MeLCu+DDQvMNlWqOW1+P1gt62ZBU+ZUTwUz8Sqy6F339eWmzpIF/675FTwKL5Fq0aMRoOQSD4bM
GEPznITFiOkbKdlce2TA4n2Ppn0Vjpl8MDkU4Eenq78jgPLc1jkZPL4toXASj3jKg0S0RSSQKbrp
PLs0Hy9We2wWmw97R5Lz+pCfjf7S3diuEzdkOlY6QcT8u47bIRU9EgWpIw9tbczPY6CIclv3dvC8
Wy7q6y+0Idm08k4wjx8w0JxLmiph7iBmnLNiLEyWegh/ACNEJ7+m6b1MVmkdL92eW8HkM0D4mY+h
OzDIZNDsYJTYgEpfgNFLFwTorAmZLRGcx2swVaUTknX2ptJg0N1XmMBQ8uS+8mgX5VyRBYZh5DXE
U2F+7HNNAY8c/F6IT8B0Xcmjz/ksk8FQFeKLDrIuM0UJUyzNDSswEHjktGFReNs2MrQ2Rgu6IwNv
wpTfDhTpFgXkdKSn0giL0eRb4nYmgv1kMV9p6CvU+GMTQajLASui7Zk/cMimjXlcfb5QemPiCg4U
vAl+1Pr+agh6pOEVvEbRNat19BK/taa1wRk+Q/qCOOjKXFDpj9LNMXT4qsy2tmnGuoF4NwMyBhcY
sbU2oM8pPHq+ZSOvqQmAzKV87EG7Gl/R1eJuHSi7nGtqzsUfKf4W3ke9OpysvDa4deOhGcSCYCLT
PRuMF/BYopBGYGijzC6tQzCcwsRFzFyweHqxid9fcFfCzMJfcW65aUBKu5Fs+eIpGFgIYN7fVK+F
L9Dw//afbrxrgrhstjs5/UEtkVptSR5jNIbCAC8qW/U7VeLFzxWWhyDyQS8XIUK+MwR+nfBWsexf
InVLQPHRyF/WqS3qXPqFHxZa2omu9g2gesp3VxZ2VEViEJ8P4qrA9dWxvgHOtitaq//JljE+hGYI
cTbccqZkXTp4Cn2f+6hivTlLL1uanmTOi/8ZbiDRSLFnoM4AP51uxMdhseBy6NfCaFhx7w6RZa+Y
n46ggKmTxVRBMvCT/tuR5O23D9nHmoJCJ1umKch7/Rf7KXKH6zKTyktYqRyLu6XvsZ5SzKoEhIBq
YHIjLION7owioGdTWnbE37kBqGWIdNYgfDoH9KnTGhYvI94sbDH70+ZrqaFAhihIZifJJQMJx8js
bc4RxcG6c/a4hULiVCl5nJJ7m4CcpKDgyPlazyBCVdkH6TWR0pEoCffjxbB2IGF7EjIClCVem+69
+3TdvQ4ZTxIpED9S5VHUmIRFiJK24K/5L2djaZmJRqgIMMZMozxfGeAoiDuhwc5pWvPtsEGpJtox
Fxg6OqhzvNqmh8B6cZ/VWW3MDT8b6yX1rizbIv/o6MkfWMow0zlRJ0fYaOdXtYc2qMr38zZnmtJ6
1+liTXII2ASvtayoW8c4GgSZLI1SlphkCYCLgCdIbHNFqNIHRyLWLJPT75jgxYOLV9x9UZ1IW/TC
5qWjWlI1vX6LVAu0OBSAcuAhixo6LCi7ZAfHnS1+OytSOfhs8fjB+66FewZvWEnc+9nKjk1FYUpN
F6inMD79pvgaQNOdswnObcVqsrGv33OM4uPhNa/yf/dZB7PGa7XxyBvqfrmIGVlINzhEATwfZCUI
6oVZ+cFXzj+jod/RUIOBXfTwfeelvq1VV4B2DIrPVQJNFE8sWOZp0hNGpzN8J5u2vOZ49GntLdM+
4JmynjqJsycU+HU9GxAlznneK0OZJ3fRNnjLFJUZBNnpgs1PEz8BLHU/75vyKQ6abA1Jtk2Dms3T
dUaHvwSSpNH9mXFOZMudn3YimqUuMoJFpELV3NJskwkfxh/uQP0H9kTQFpRC5jkIQKINN3LZMPIA
Aw4EJendHeWoKjrqkIY4OS7Vy1EsHM8Ew8xz6iz+UfoC46RR85oqY1Z9KtgZiziUR5bne/0HFT3x
dT98QYT2SMcaT23wfCjLTigQcnWzyIrIKHmyPxTVUAvbut/DeXYYCKCIXhduLZNaqiOBiwaQ4v7f
4DsUmXEYcS41As72OTuQSJVz8PbzTr7BTcUhOLY021Iwf3OuD9f8iDbKbvIg/KClmMtBWsWvDGHj
7ZKQNGd6z8thbxzYCiKpWDl1DmJNEutTAD6m5r9sQJXClBhpto8ouhZohngUTbAqaosl7Qwby7cC
A1VHid4jyGX3dCufvxtbmvnpT/IfSl2J9cN6VR6nPQNiUQFIkD/n3YRJYvVA/2fLa7J0ZwNHT+mQ
akb79iEB/0EOFb+Jj5vuRmr6e/TJLs19J9A1+5QBNDANG6MP9zhzihM6TZ/vVVOFkW7txbSJu+xo
gqEGhzuQAMkwpg3oJSPEs3T8d1k788ywpK9mNN4I0FUbNZEBBrD5H9nCcfNJLuv5FDqNg0FvCpGy
CEncB1AudAT1I+DCXRCuQ9Wp3uCmNJRG1Hqy286sjffmDo1Qsde6XhWONscS+TOujWDsqRC17URX
Lu6UTMUTGxMJdwCuzUPMF5Juf1jg7uL635BdhZVfI0wPPNhHR1MWxBuMOkVJc70gtPcJ230cHZuh
NicA9Xa5ZGUaXvGGmDPYvVjX1+RXHnG2oU242zEcXqZl8oCNHtt7PSDP1UpInQ6vkrHhBjOJj5og
tSw6RbwjZbWf0lyx8FJxppZ6sVaGXbs5Aer8g1uPdBucO2Ajmew/bY4iflgu4lm+F40pkXjJbAGO
krgUhdmEsOQ0fbXORW48JFfqa21yZvsUwYd0tMw4MJnrVKPT6W1w65Fx1Ux9Mb9kPfA03Kes8K6z
IrxN
`pragma protect end_protected
