// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
j9tJ3j5w2u6HySzvYI6wDyj8WDQzrD+9txM0yiGDaK1s/qHOiiPAmiuIV1lwKmk3
XKsv0W2Xn9qr5zMGsf5o6C8MvApI9ugrB4HanZOEUp3AsFuQ0YFdqAlEOkpUENIi
yFMjzvUeqYBpcR8k9UcaYaLXn296YqHD1aSL9LWzVpqVQz7Cy8ks6g==
//pragma protect end_key_block
//pragma protect digest_block
xpnuYicUz26O903/Xv6f7t0o6o4=
//pragma protect end_digest_block
//pragma protect data_block
NxxgpO9pX963HSNLbQrDCLPHV6wk4T3jNmKDGH+ujb4oC7RH0jd6xyHjK0uecK6C
0q+e9sUU028DF6T56mMfHdPxzDPdeVhPWckpcSlxcIDvgeNcyi8x4ZNrupsrT0OY
ZjsCDk5tIRezqEJTM02aeBfWWI3yZtOJZNKDYElmq4egC/CsI7sCKj9wwQnquAbY
Qt5v2ZqU2uyqpin9fcxc54hTFFRCHEbkF5hSnM8UCQ3BnMhUx5N/ZFY9vDAwe957
qhcmVYPp1zDnbk4cZ7qI6dW1aq77JVB3SoQF/NxSR5kdhu/ldX9yEdvCn1No5Ghg
KStzB5iy9g4kz0/nA/4eHOw0Zv81ua4nTk3r2QaloXJGNtW5tG+Ju+mQv+X8F7eu
frdYWlEzMkwMEHS0K99ZmOhXOSUETYwMU6snpcH4N7TbtgooOYKBZU1KTzGqbsxY
2kie4jJZ2+fSghX9nwPcS9kg9mdgjMop0qxl1mRgyhh8EfWnrDtkU2RJdb0Z0DEm
fkEOEFWR9Umht83544J1fMyqTbKBBe80Ua20CxuXyLdofWmkEWez+hP1uPm8FwS/
bprwmGbSQo0IWz03kpP0HUq1EU3G2kNl/okizQUj/CQtNlsdRtYIVnP3mU4UckAL
5jKPDu8H9SGXhB8XzV5KEnBQ63mCETRPaH9NkPFfgosgzLgBaD9NsCX5te1yuQIi
HZ8JDKkuf4vi6egNRQ3XRCbSEUTHqhgphFStbYG/ooFwquKOTwMSXpMbNjVrG8VP
Jy/APEzp132UL092fJ0LnIgzNp5ln4DRn6g/exQoEN2ZyL7LfKuitok0CC5HqTmc
AVp4PUB1nk9qv3SaRoxHAXr7sv1I5rQfbe7Ve7sfCSIxMZbhsdTZFMUsUWhvuD+D
s7PT9HD5IrrPtfjMjTOYPNXaj2a1Y2J6MQlgX93XVQVm3bWRu1ZDvn08fLw2xX7p
5O/7PQ58oIIe473sjOxHTLEjhkwBmwqySuBup2tBUAqLIgj5m5M7n/VQNYaD4GU+
jvvNsZVivCZmzSJBT6IumdceNiYqvQ4c2GWimjCtbcXnZ0gxnxCYx8yxshqfmjjY
d9ca1CWcUVZCjEfllHi51M+aXMbIWnbw3YbcG4dhQUMuVzQJfJoAOMm39wEzxBVr
Q9xOf6/LZWC3sfR1OxjJCaRpJfUL+0Z2Kx/bV2ziGxEM7InPx9kqUg3NeRL1WXVx
n8bmSJUCPQlafgDSFaz1CaytNIOFmejhqYsGqBqiJtV7uH1hH5m+SqpwfCrrlfyi
PqYiqeK7IhqII9pS23RkyMGs0DS0DB/Vz6aGBl7fMT/pCbaDCS/B7jsYVNMYmLea
6VAJUhFYLzmKyxTacoGpGfXckrI8+zoX7r51oeAXSYPjPbxbs8hyPmQabyHOcd7Y
UBzYUiqc5H6zntbJAInN8CJ3XFSJorR5JF3rXUX9i9b3U9lbx6Kibd3gUZQ6HDyI
tq2tjX9yl2n19TotZFT3SSK3UnU0F7cVma0Rq2Dg3rF5ORHtVNZR+rB4GFLMycSm
NLjPduRfwvzP5qw9zKAByq7AHWIc7OGyqLvbQ6IFlErLTULDFHAb48qTbHEvKjzp
DNmeUaK8LCNa/a9UBo/KA/t1zMUsZ+Dg0mXFbQVOuo1gboJucuTLq4S0ku+sqTWR
ORTg6nfYg6XnAzdcgywp/FNqo3uGEqJ0bY+ZpJmXUeTR5VLw9/7OkruGIWjUROTv
Spc+BU7hwkwO3tPmAsDJqaYuIwRqDmS4IMHsGP7BNKOKBR85ZvGqkHq9j9yIXyW5
ey7vqM0tU6Vzva2RHszpjUpNlUx2ETWRXKoVF+cV1O9nPaRzeLOUCkY17kjVcWJU
K4vuxYctmsAo951Mtc27Cn3oYUQrKwiLCwqQ9tfs43NIH1a8d5+qDCIHDCYTwmDJ
j+g42ugY9H2FJiAOih8P74b8c1C6AnhxEWPj1Orv1ygAO2JLvsTiZ8tXql2lvbD1
uaJaLUkiYvlFG8Bxr/CXxW7+KTdSpMJycN6fhNnE4OvMG3xz6dDznH4Wm0QmZ+2e
5AePWq2oAoBydGMnWO099PR0Xcu3MDPoyAEgQjfYNkTra+pA7QApW5ugnOSZStEo
IGo07GJLDwZkj/PPSiA7StrlV+1WtsswqNqbYaIY9JOOASjyom2FNFz7jQsLFZaj
/1ilhDy8mJcWcq7SfqzZ+FHcsnY8bG6TAfB/jocRRVrb+TjIajNB9iwq2Z/OMeA8
xhwGv5959Q6/aH9zbRGHtbzKBbIfjb9xJo2lFJjyaULjdrbafXcNsEQL4xczCF4F
KfSORfDknxwI4vbKp0n8Sd1Sk3v3/LtXhrzsS9a+xJkeRHTWMolFkrX07I7SL15o
ANEmRNRNHp5xZ9iXnFpHqAg563GNP+mktHhHkvRgq3FvAd96tfTc/tRV7lXpNlNq
TDoNQQU1+8iyV6mvu85MdWDeI/TebOG2hpvB7kEt2I6RaseY3oZCP9idUIKT6hXp
sYA6vtNRi2tSzeros90LlDneiUxTK66boosuyFsvKlKpbC1v9w+mVbp8YJZtrYxq
xNnYFuYrdGAnjq2xeaGnMu5tPGPQ4amHoGm4eqwiUwpgLE3yIECjdg4sRt5pfJEA
GibPhT0DLuyF/HW4VElzOne7MWMIvG62GAZhyWPQ9sIzF6XJO4bcBnHOEmqPPa0c
hwr4iU6AmnyKtb1o9QeviF4pPAvI2+ghNU9depx7WIvRfI9WpGSIABJ5E0TF0avQ
jG07R6WJ57Soqk4u0YT+eSrlDLO8PNZtc/L24/u6bw2BFCq+fD6xUCYQcGgZQlzG
KSUM7EMH6QlwR6otd9wPx/xpcmQdlK5JEwU06L0ErWWdE0xqA4fCzZKSrPz7OhPF
coNuLPstUClzwTHFmC3Ufk7mEYgolpOuc27Yfx2gXxnIm2QAfjGKLvOo4Bu8UePQ
+cy1HPYbCiQZgPAHn1Eik48FP4u0DpB1oy0HYneC2sG8Rof71bnu7RzDgCYYhXMz
cWiDLZ30TnD3/mZJLbpyL8xftnZzI8xUFjqvkdZ5G2GIjJ8cputd0+lkzh6CKeC9
Shgss1f8f+VvAA8AYVwOe8IsHt39a+PVkG5OO8XCBxGUkH+7XggKCFlKTQ0vxkE9
XtrDX2zs8kjCrx2x5y5Q8YJtAGGOUJADjHEOJVDfmTFnxxz7dzQaVbjsiPIdbTu3
tUXjrCfHq3dairq77nWaL6k8jLjKQMu2IFzP7L20f9D9wzpjpGLcqQQoYW08Ruef
SEcH79VYQoZJHtCoDCJmvRk7pmWecLsmQodpjyWlef85ljCds7tPasrKTW1pUY1i
KCccsvHlxfP95G/QArHe1YHLLyF/sDjaTnKyMkXO6keHtft6cdU7tvMilaxhrN6/
wWd2thUok/caskGYDLGZCe4WK425ZjwZff2bACL0zITmajqFx0iey3wCFSJ7DNTZ
9e/Bq7hG4N5iAE/s/FI3SA5ZGqibyxvJiwTjCYtxfztc2Vlt4MKdq2Vf3eLRMxto
nfpNymVqhWJOGjFZSrNHPdROlYrhH2LJ4VUOmdinwmhLMAvePtVc5UKDVHhGf5zi
Hw4TThnLzirAjq/QvwcMVmxCwMLRfNCPCdy3Xdo6QsAuwdaYDf2dZ5DxnypnG9bJ
XdWoKZC43O4jKrTvrmMAWLHM6eqmlj+z5S1WdAW1syswUaSy7nnubw5C5mMkdjjE
z30CKbUsnOrPD6sizyyeKT8eN52/l5mqY3CsQ0pvmhWUdqxVKVlVnjGeLTIATVbX
BC/B3/5tGfrNMMM3AWuxfzUXPGtFs7zlFwSky0KFEBmQvShhTrPMQWMAFouEP3gQ
hMFrKuExHW0V1zVbEilqQs48KAv56UYNhzlqKaB1ABoMM4RDWSW/aEzX1dGKzAqm
Tad08tufcvIIbsIswtbMbTwdFeeoSxBwjET7mjwOpPdKhetqBNv+sdj4P7N72H5k
NJMiYv6NZUPdvILiWti3i0xuusQKjxTGRbCMJk1uW3b8T5Rya8dbqJHSj46ItzOY
ojtNc3wa5DEZ3+RzV5eCl9nLbzpcuE/TYOIfDwlndBF9TAyLzdkCopUptAufZV14
MG2VmxMyqzmG5jZgUnjtzcEE2q1V0j/Rtub5UFnKMdO8xcIEUzoKm220sAzj61uq
2VdFifEwZ8S+bCqsS/4sKxXqWxJi4GUw2JSJ45Zg2vnUYKo71AyeQcKBoba/JwBA
qFJYNQR27VKwZ1fByy7AX3XdGl+N6HTizOzvrdeF+9fexqPdyWVAKHa3NSSQQAyj
1vTuG3whxzFurxadfDUgi3iAgY5A3hIqEnHVHO4PsFGEzIVGXZtdnWmZ97EvqJP6
mp+icQvMhbcwU323vHl+XFCoZ99HI1eMAjj6p90tNoPftgt4H+ipSbPOlBx0mRue
NY/6vQxEceXoBLhtfrQM32/NPGGSvngpY0qCYjdyI8c=
//pragma protect end_data_block
//pragma protect digest_block
Pc+xNcqv+jP6b0sg6mHLuL50MP8=
//pragma protect end_digest_block
//pragma protect end_protected
