// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
ehv7bq2I27e25WVgEExxH+Ws32W0QOx9NHqJ3szRGx1Ws+6KNoHG/gjVpXKh+D7O
HnpXQ2TsvFAL1ERLICe0afOHpTpCYYrmHMtTVDXS0zhGzRtQh7Csd4wDZyl51yfj
k5kHZygP3rv2EDQFr2i59NRz0x4BWSfKCDyNVg2a3Zc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 22736 )
`pragma protect data_block
CGaohrLqSxdCNEc37DiAGllkWZYy3ycGV8mILJ7y0lNvKI0x0wQko6R5kcUDRj0i
pdOrnFc3hoAP9G20Q3GQh/PhJzMqg8q38Lf0+YBxS5i5lOh7A31NOiYizzJl7ffR
4YhUvBlVZiKlyoHbH5P96GjHsW4jAOF/eqc3jmsNupCzppb8iCcgavM3KZByfuwn
mYAACRB/TGNUU4M9W4+0jGP8FohDcdI9FWlWCsRe8kfgq0hQb1QR7UhvyCHRhEe+
ywK7Svn34EJ5yMMhusUzQLiAbX2m73lscKbQfsUKXd6vfJIEhAfyTzinQHtvvbkf
oGRlEnW9KZmTr10nDfCUBUHmNDHyywMQ+d69LLv/ihrv9dBoG01VmHy5/x9shEz1
P6CU1x+mVXRC9TzeeyZqEpJZjpxVH71uGXZsi/d7yEzlP4UXGhPIGOIojCvxR5Jq
hR+CwBTQA60Hc8wc3518YRv0+7ANmTddtth7xJds1/9U3pdz/5564xuxPpaVOgzI
FU+i/4nv8fC8edrhqqHxOb1VtWKivKDcZkKX/5kyHf57LmBU+u5jGpjq+gb7ZTdw
IvNj5Ci4t204A8OOf4M5nvHGly7jEWyYNyPEQD6KuJSkraa1Yuk4BGR6+EsO3p+Q
BNc4K6XhDi2YX7rI8xBEj6+3i6XcvRpb1oEOUnTXv1RFbdAfZ/pW9HRiDJEOqM2w
oJTpSXcq3nNN3xWlx0fq8wMY1LnyGA6yF9ZOKwMmkxRwr1ky8xJV3/W8toOCtdZP
cw4ekN+Udy2fv2/TovudgdpXxgbkK8TJh8QJOps4pwQZxYT7PcsRU8fLIMyYVcvK
SXklByoyWzdA05qx5XRFT1DJMQrVBZZxbG15tOndI4Rhd6UB3OIFcqJ6PukcOeaV
JPtqxsyZwzXIMQ+ghnkLfcNqm25kpEqiw8uYUpqJ6HYFbb8JB6A3V6g/2qUKfMD2
ZwVWMgPljyU+mhpvmry3CpgH5JjsKx97/iKmsF7AW++Sn8TfFbAhLPcSQzGwBRLg
AGIPrsFP2So7KgcvE3fWCX2gOu4Rei9IfyYZP6PxGv9r6VqUqjBk5EnLoeQfBC3e
ni6K2Thpi2bBXhPHK05Egxg1jUJ6aaAU4FhsaxMETZ2TTUdTnL2t8NoL8gMuZlQX
YnE7MqDpg54pZNZOjl74s4asBRtaE6eb0cmYFUNSIrvml6Ye65NRUzePvfi6Udvi
jJUtpVIuziNr3QC+sX7Ynu0U23nx6vTN3KzhPSkTe+jdvflol6qpBJJilw02hf8B
RKkvuPGCxPDR/MfstcIB+xkXnKNWwVlwccA1jGzwW8pC1nhaAwAY1A5M/+kExsFa
fFp3w9wTvJXA8jx7WAfaq4GRpGXg/02926nnnGZhLTMI1stwZMrOL46rJA3IwLZi
pGbuNDsyi7zl4qclNCpjjzDybNJpuL4I4CLModkGBeBgsWAfwyiEY7CToEI9Rvep
YPkmmi6jYllkfgHVlSscdQoSMJUCpKlaevzMYwFyQADc3E/KXwM9clmeoCal1qa2
PJj6zTFY5T0wOtnHjLCatsnQO7weKpduGfk1t/Y/tcYXNNZB22t7R2JAsdH6Nbr+
JzdD0kdvFp/Akpr88DEZPIjMFNn8bjEynejv3HJPKPMAVHHXAIVY5oN+694yD50J
/tOWCU1Zkr3dlnRjvh/w2bZKLmBm41LDlj9B0FM1JfTbUIylncU1n2HqYngvIGsg
QwjGRgDMSL1nFOfeNFs+j0aekHU9GioUmcjsL6DFmPCjHxL4MrCE3aEsQYBae9rC
oktGYYO3lLa/nYd8qw5W1ZNomDtWQ4OgFt+FXol17n7Bv3id9fW0y/3fP9uDKYeg
iw3sRsq0cY5QeHlkaoiqm3APfu4gAaAdlM5f17fHi0+ziFndWMNTV/1/hQzMEeq7
XteMLg5YoJvOlVrywwvKZcy9Hyi3tVfULB8lBuxDMPgGbfzzb34oYt1TmhUWq5Tl
fim0GaHIFmhK5AZIcQkcdKgW7rOfyWZFAHECgmbQ642kg0b2feIzP8gQ4AXvil03
tnC2MYBv1+KphOaOpVKhcxcbpumfOy7Cj7L2HqxlaixupS6d79vLsjr853EgJLma
Kp7sVnvavCOPAL5EyEI6YbL6J1EjDeFa2aXx8zCLdFk5G/Q47tVZbXOVMAP/lHSc
vgTN76LKjGxgWsxJY6td5YN1LjKkrd/LWvH/E5Do0t+7+gdB8CvqTjJ96ignY7K9
ZPlLyBhgtEEUv2sPNZJRp2PeoIOA6H4N0r6X6yOaas80ZUDwkYAKZxLfqKZSzM20
JASWTuasvwIlf1L3NpHGuV93V5vit0kDt4VaYa4jfhpMcje5RZQSFSwelHUBw7lo
jmBe5W7weHgjsVoza3qrXlci0udDufQqMANwMfBJFxK8eGm2k4dzekwXvry762At
eqJA0J9lr8Mxq3SaRdnjId/URIJYfNlI23ymCEwRiNJPg9ErvriFj6gBDPp8boq4
BjunQapV8sqnkyqzWTGNF7KXarCf5Y8H5g2LrAp8kzdlbl5+d/fVHxSf9ZiBHtsF
hTDKb02gifMQ1D+gDZjAEx0V9kS6PW7YvyN606ZD7ic7y2SKWYVorPA33ZLXhgCT
auHihNBNQFMuPHumwhFsWHK535rboW0xXG7r+4PiLTwfh597xIQxsM5qqh1KvttT
GyXPvVK9iix46M98Ma9848QwiNzn07Ekj5vadnTlhxOzitl0qA/WSs8MWU8R3riw
EIVm4lRBQ3/JYTnGZzwXHJPJWhTt1D4q5AjqpcKwuF4TIm9jceR5FNfb4o67+7A1
+SKNbVH/E98crY54pGaDkuLLiqTD62vCfCj18s44JXtzY3BdSN+Gvp0o3jW4RRNs
DgHVoDPTCnUTQnr6c5tYrGam5F27KsyX8SfBkIC97gd7sV3mjeoZrycqwx4+uvpS
hz+NAKuEOxNt+LLUFP4Dtv/p1coF8IbDnL7hwPh1JZQSEBR/SRxtDpQYDADrB1KU
LAaYs23jNu5mzYFmnQkYztDFCUHMmgFxulXFefhdLIAl4ME0nTL7AaixufW5y4u1
aML5IgKBr0jE02Udu9heUH2lazn214mrEg9OZ57/mfpVFpHcEeNolGfCkqVSnzvd
8IiHpAJb+zmlnS88vpWvyt5NzTm5AWAlUc282m/rl4xK3HzFKC8vHgJRvoBHtnX2
Bccyll4Gb5GEKRx1komfJZiNebcYIvx8U1l7GKI6qwrBWrgUQM3pNR0ycb8HMF5D
eFcxCYkE1fSLI4QGiOfa6Hj2casCIqkaBt2507ZTaJ0MZfQpBPxRRbYGu3eJQKEw
W8E0WLvOlqpoUAL0S74NVSTKvyRThLEmwIvLFO21LnjhJsGu9+g0SAVjl5hHgen0
Ji7DJbb1l6o9MZKC11dZYx5J/G0KkNYuFzMzksVVOYu3wDdarXKM2WQ2H7AIs8Aa
sVQSDh0x5pYlWuFQEt8rZztzLzBjm6vGWGLsVpxLbRzMxQ+O4gVGSpYmo2B10ruM
Q0ZqHWx42dIAaTQ2fURpwQJsjdYW+v1de2sBh+QTEOmF6omS40C2xBJfN+pK15oT
vreewLqbk9yUkljvXa2Dgv5kXAxyc8rwhMc9BnjrRXq7abbdemO0idp0+Mtt6Ao0
8u4zh34GWBnPWman4F9zrUMDt94bQZF4RL73Wpr189AHvVp+KIex2JQUcwYvqHk3
DOdlGEkOJbqXyhCYIDz0/0l953KADasGAa80JRQ0RYPLMS23w4eNGOZuIEw/FROD
fdDX1hs2GgpQmwSSfQxHhfzkbnfxFfBITdNNxq9i6iL4hH5/JngzzqZEnPzO4JuU
8+1qUgXAkhDO2cq8F8trua/PrpV3VVKQJ+D3Gbw/IE10U6HLvXhoxYTpX2M2hYnc
0YKbdIFeDiJJRNHUaE5bSisQYSFVZV5zDcbFs2wwl/G5HX+Aj/DyiYeHwjWV6VVf
UCuLLU7dJmKOetMvg9JyjR5pgy3onJM5HvILIYa+vT66KseJbp36xnYfWQ4hYe/J
KA1TMvlly7sXf7x47hZsF8BrRZWHIjd6ODX21ZJrObrwoznMGeKpPNJbKcv+EKva
S4GrJVe93jasGtfblhGDLKTSDwKH4T7GK5pLVL6xjXq0IqPjLeBjYx2ap27wonEM
18O/+BX7PppRUtSEE0X/k//mGWqwPcfvBZrIJ0Tj2dNFMf2i2m6QrJm18XO1Olna
nYhzacEUp3wX1xfbpynEfICaI8AttJkVKaZmv5qsqdFWs7FBT0FIf99mufj4lbMw
5UAnR4LfyXdtbG/rRPJ7NkWJTC0ZMLzG6d0OjEaD9q1Tx/GJb1Kp4jxNW5h9I1Jx
LIVz/vNKSMUIsGAKhg/Z0JKBgjfSHlccJaj36iwTVB0L9WKAS3NWcL6KEdjf+s+U
qmhnlEa07MtKiqsY5NgW8/R3OT4pj+5apdpJy67/86ymgo0AaMHHQPImVe8RTa2p
fDi5JZ05fusKcFVr2OtGyv57BCzo4SjEtiPdtb8p7RONvj3JfhEXNamgjqRWqJ/U
V+pwmg9UfQa+6xn6HMu9DoYErZ0hligk56FCvtj0kJLqlQ5f1410KSPMtwpVnHm+
hT+8ZlOKMV3UCHZzFn9LixSBHQ7W2+ob+5xQPuAjMHKPiV+Mh7+QW1MlnYUpYTua
Fu/Q3gfV7ZKtqha43BLYsM+Q7+qdiAyaqDhoFi85uk+GKf3/IHQk+B18zQSEkDNi
JEHlPxKYgo4QfxlgY133/SdHg0joLqyqKkMfJdAVI5HF+ujpf3eXDukvU/wNA0f6
0PivtWUiHo11vFjW2/eDjRK0GZ6T/n7BJEiqvp4cur693mvck+7eEewpxyKw8ZIr
8IaAeVbChYuFk1Xg1Q3iiwV8mV8P+ig1dC/0vj/t0E7hfUV3xgWuFUISNH9h5pWJ
rUSzIKo91O+F6wv38KgM54Ttfyt3SD5I7YrLHwhTWf3FZCBu/b6akfYL5pYvlnvm
rRhhaye5hsKh8Q6iPp8kVDAGsiW90McqhSuNJ8pCIGZXchI++hLIG/qMfcZ1MHnz
IS9dR2t294uy/7UXZWa9zcrtYHZaN+5soReidXu2pFLCKvMVmB+dDfVH6T/kDmIp
2zAcf9li4h3W7dn5sdj9AzxVWmeDWZGUeR8s6kaxft96qjLTD3f/Ty9N+yS9RhcH
TJoqs4KP1/I15kwsVU32fnWIUQZzfmZFxGRwKNdX5H6Rk9zyYaSRtm2756cm+nm4
x8GRtSXO2mfJcXJIsBOEr+hJV3x33X9AzcsnSI6nveyxnZfq88121bm/A0SOZToo
YDTsHYVcG5OmGnxGt1XcF44SWNyu0GNFghne90ZP+4GYxkfWUe93cS8rRAz2U4cG
D5Hfil4a6snhjvQWq+Yk35Aa5U9O/FQ3fThE69JE4ghCI4v2sd9aIml1mCqkkL7P
QK6Z5e9z4FqjoevrzU1vUI1RhtgT2GryeXPqH0V0GQRT3IVME/7GEiGu7X4YMWG0
f6o6LDH/4PTsN0r6Vpm8wzLIfHTgNBO1zZajW5XgEICkfygwhpq+CTTjj+m2JW+m
71IXXWY8hLmDNTAvg1Ry0uSXsus+Igv3WXu+NvxuoFqHhBd8KjymWtsdihrCDLil
aa429ShYSlg53Ydt9AVF1w1WxH2r0LZ6Imj89qHdIFOEKjHbdKBFT2XT1CJBFPsY
ZhjAjdANx3dt0QR9OdReGA9l7b+WUyn37Gzt6lTBs3pZumKx5sV4vNViuqFPpd9U
YEyoyPDKEzDHQCj36Rv+ZJYzsp6f3sQIqAQfjlLityEwjXYJkDludMdBpN3O+jV8
jbxxnX+8W6U5Lv6Yg6m+MoPLPnCJkNGA9nLAfff9Gcbp9v/fDGp7qBNFH30W8Xvm
6eYgf5qM7IYVAyC1tBVE3cqlsk9nINLOX6TzBnLXOw7SKLz1TT3JejrJCRhGocag
v9fw10lmE+hygFQ2oE44igM5Mplj8quc9gKz5CeDwv8r/6mUzNnpnBQyuTDoYhqF
I/hl3+fM7DbQVp20s7ko1Y6q2Dl5kJWSwyKKrv1CELAFUiNaX4PjifBxe2NPuw8l
xgbAoreJj2ZWaK/8tqJhU66lXK0LvxOxek537DfxYFjMxn5c7EBR1ff/YZaOQeoD
139bIXVWr4TYrjV5Y+3pIP9I3++Fdqx/gfm/pzZj2rh3vaYYGYHgxnfx1CTEJ76R
XDczxwxPWReanK0+QwS8ftrUA/sMJR3JgzZBOtQInCU7M1n/PJhz2GMeqcO0gxKF
8KTep8TO2GC7yRLKQmDYJ3OgpjQRSu3tsKRacMMrpy5fWtykLSQs/Jkc6oMM3yn2
f09VKCPWeyvy6JZhUoehFDBDuE664XqyiGDr7JYNFhaJVwau6YGCR8D+jZfE/LG2
wIhcjE49jyydLuaV2irvOBEVzyj4ZuAu8yd8ny995mT/rgb48PXZLrbJpHK/LpBE
w+23KjnyUoTNT/+cI1a0hQsV9YdJo8YOTiYIZIZGfKE3ga+xCQk6ovTUcWZpNPId
I6+BQWObMUS9gEWUytntq4V13X6LtKD+CGcGM27bmYMaKiUg1c4PtO9oRU4zAp7T
mpYXyRqANKfRJe1+Zy0HIRYW7PjNkYEPpbwt/OcTcE3654XvStSl3YuqNrStp6Qa
VJ3NSmEAhHWOo9bn1wz681a30qhkSsePD6u9xf0d/WWnx+o2eAniNB2Wt0GRayEg
hsQ0776wUKl1Ib3QDVUasicMVf+OqvJ1VNb6CbZueKagg5MLcyKQjesAiDAMKlc4
U9QbUA6dvipxs7s6EaaNlTsxO2kzOvjo3B/ZOrbOxnZKEB1R+hNzSlCJQr4KyDCT
OIehkpW+Ank0ZpjdrKO8z+1I2qkP4pttnYlrk7Sh8tNaIlRyAFZuEPdALeoNzbvb
AYBI7gvnsrhFdKW9Mh0DBKdbYrAz64hewFIwRHgFJXMqMdLIs3jG/5YEvnWdlmWB
sUUXm5xVFLrgLKUk/iHiWQSmQS/bUXe4mFUdBeX4DDqqV6RMptObQToXfORjVLYx
G1RIXynswi2X22NY4KHBqGHigu1QVdrPuorNnSML9E0g36q7ncT33pG6GKZmYZJ/
F3YOIj1OBo3XY/qYRpHPxfdIigexVAU85Fm6xlVh8kbXB9tsul7CcWSOsgWCz/zV
h0sE8RkkqaOOaDu8x6e5Kp1/q9/cepBUh8zuZfq10Al4XswNgKd/Sm+qTI898Dxc
pG/cg5esk6PCJBOz9RCx4y4uGTH0KNGBtBfWG3Cxz9l4PKZ17dMDBo1SblSQOCQ2
XQA8gi4iOknh/czB86UB5z+h5W8POzQwcsuXV/0ZQmtl9RQoSlDY62jtmBPD43DH
nWY2fgzzWLnTlqTftURk0UbIvtIJQdOQkBDzqX/rAVx1AdOUSSy5iuFVf9I1egpV
vc1eVdzGClI2tXOB9whwQmkOnX5NVRbQcvIsFK3ucCDlojWpIvXIDRTmUqTJKbHP
6cOQJZTZtYSltG4Qgh/UiMcL0SDiKHNcpyvSqYwh/Jt4Sg726QdviMcmHjIYWO9l
D+LRjKliYxu85hiFQbOUYt8NAm6BMT7EPZooZgiGTBLkqH2YpNfCTEs+/c0Gb9Ey
h3ex3t7/MD4unh9VgxbuiyiBmhtXFY5vbRwIsMfGwlKeyAZQvAgIvO2MdtuJrI5n
45vsvbGfIkwrE0bSjdf9bpa+HYFAY5I5vLkRrkDAJIYag8cix0RcGpcwK7T1FsTk
WHPCi84OHbOSMJgVvrkpf7zGKpNZW3FkUjRcba/clb0tv7Rl6jjD/St6uA3/d0//
ZxPdqlFtAG31OehHd6X2F9pJjsof7HP3LtqPduq+V1/qBd3LqUhOoZiKsWyNK/ZS
s3xo7JmSDAQD9ISGJQ886V4n9OW/Nu+6l7k/X9DUL6rXZHdSI/Kn/RqWXgK00roK
3JGhpv4oQTgkS8cmZYPBQ5c4p1aOcX5YFihuxb+slgZ+p9TgglG8gBaQRYZr7qPa
8MgO5xlrfoSvloQuFQfE4xER+KIG7lFBCZLUwc5i5XuOAmjCbMWd63kXFQXPHgKL
mIN8CD96Gr7nzfVGNVDboK8YGioZ3AHqW34QOlZJVy/TEUvmEH/SZqLiFlgZE52k
tBogUEp1XYKrKavMQ36G2VdZg3SdGzEqOXSaFldat5ZP7zIIxWpuji0KeLo8J6xr
8Mb89ZVKEC3Gnqxjvf09lC6SF7z3RTmNz2uAhzgrzd3ZvAdT9iU2isKuKGWYMI3q
UAP6JD9ZJ4hDRPNqDqvvqNNCjocLpa3ulemykfZEYegwj+7vTQbrbKKhFs5wEXyu
W4hWKDKaLIUD0olhSnB4po26jj6JoeaedzN62zBZczE+FsYqLLiS8/Y/Jn5/3BZn
AWePdAzKaGsTu8XCPosymOXLBFgsSirP31hfyRS03axLjoGumANhPSWX70uM344u
aSxQJkLJMS9q36NC0J2bdclsVVgL5PZEWTYDTMATGugNq0jLMgo0mx69mZmgM2EU
cF6rRyHAEtltTnY5imtYJ5eKtw62WtoZOqwqhR7XQMEkM7yV1m651Zp4XiXOB0Wb
k3TCk485RM/PkBI1hPf7I2hdr34aQHtcU+Uv4o5KSoIAbCDdIK9m1VimgfEPoB5e
END/Aj8/SiFVy2XUICk50YIdUo4yPNzOREqwTu6tKZzn1NCTjw1pxgbZCn6BJfRA
kkDmgMPUPPOp9jU//8dvupM5mON+q2trjaGTnY8ciyUrw9XQlSnnRIrGSKQpPCo2
epbL5heqtcqJQMIm0PcDCivUsnqbHLVyrSlNkguGTOj+Jg8FFjKoQNQrLeF+kp5m
gEQ7LwClcnGWpSN3Au7z3UaXpaECjEzW/SyHV1upPDFEG+yjniWXQQXTvk+Zh1dv
8HLGSpE1qorpEKH3H2ReNZRkusdbNX25X9HqGkaEcoeK6+aJoj9XC/rJ+7wrLaDm
vOyDv3CRX90XJkkEPC0tarNJyzYUCckQVS/LseBuLuAmu6HWav7PWLD2HFDCx1b3
Nh7FcVM54hIDd5UKPv4ECgA38r9i18tNqIm3JzzdtqcM8ytimd3NIHQHV9yI89Nk
EX+930UPHNi6zFBBWZe+6SQRbr0JprOHQ23kDFxH4KQEwflD3Nk3uNkUjlG09gb7
UGW0Ul6kqmHts5w8ZK6sSneLEn6zFf0H2mb4ac9234b4xecrPhaBxvvOtFRwM90G
r3rFyKhK4FoQ9Le4wADjq9uW1mqYVDh9V/NJHrrB2GcR6WLlRAm+B78FPRWwYSxA
SnuE/7cNgeOPilHsXENuGZbyqGpFHE13z0d2Xks4ZGO88d8VMj2xJUmLdsBGTM7U
bsnv0gOQ2WpSmrEWs0gTkudydEEFmw6ZACeOn7c7gmisIbk+UFN37YTdsg9Etasg
NY2bqAQTYlN5w4nkes7RU5itfKIN+9d0OzNfK9rJhcQiIIVPkIbEpSC/Xj4eH0Ae
OPv5X0F5N1GghRVm/UQMIALVVuhMvGmdb8fuF5xkvjJtXe4l0BJELSnIM6gCdvXn
+cOjS09vJQ4u5f+kHocS2P7+Qwfl4DFzxt1bvam9AY9ImTVV+1l3fADPOc+57UWu
osQ59FoUNLGZRbuhfPXI41K4X4rlzOchCk6HM011bNLIzYAs4kXNLPUBE6d2gsEg
G28rZfuiTg6RyToJCk8Y44cZf4Qsjs4LiHmLRcknpUYdkklu5HhmCT5QLJpVp/Zg
P4Pho5nFn9y2Kr1XUb2yK8j74/eKCOEjRlx3N6lkd/89wemo+ozc8ddiC7NnA3Ad
VI8YGnDipjj1ql/jukkeXpzDdXc9iYJLu9d0ofG79RTwwkm0xg91tSTzdJbkrANc
SCnzBkjigmiuOeZblkKCETxC2FBR6GZvuVvTNcaGgwl4AwFlaOnW2vOZ52LapNkM
Q4YqmLBy9hNBaWTvL+cDjhyKKKgFjWKuOmBWvHrDQihqAkmaJNDBXQGCoKwklFkv
MpL7JnG10Bk9S061Ec4CvZUHU++3CuSAm3wrEVoqjOmB9s+ymEnwU0UO2vY6XQue
YWUp89Gd5shrnFILWnHwZTexSo+Ke4tSq7TCnQYyELQBjif2KHDonoIQsq8RqFHp
hw6PfjMmIGH5i+YlnKSb2RKS7BrAYYJaVfkZIFXCD6CO22OS6Pl0Bvu7sKzs+iZs
OV6HuSKCxoHsw0NJqq1igdjOOly3OURo2883yBL66C20DtaGqfJKtcP1PMb2Pqdc
jt7OVLVvEvcQImxD0jpRM9uM5ZniJ9Mu7nuC66q36Nilv7BqdPQ1XkUEXS09xKYM
rVAje8iHE1JJA7Tl94d+4w6+jyjAKRjUYtrJweEVM22KGkAZnQZ/1YI597SFgFBH
+1Vr+kSHoPPPRN5qn6x8ocXxO6cnAiqZ4NaHyYRPsU0vfbOjKWVz0wCbtyAjNVBa
XXiFZOvqMrQcl8A8tQoPcAyDrqMG8u8NC29l9oGYajX1uAZUC+EM+K3L7jq3pg63
SZSsuNLgDj1zumFFmfk3f//iNfiOx1XUyU3k7Xn1nW4PPifPsAzCA74b4vJvk5a4
U5jz2S2pFwPORoEJyv4SimQWf51suMEMRf9c80Du3YYKL3DKCAk5UEFfP/8prT6D
K9INzi1G/VxtpXCJBIiNEb0bgyEJdYgCr6h8+pvbSEnW6AGs0+rwNdVhPjftzZDv
qBG4xMXwVkGNE52pzn2PIfKQsyv6zgz0wKM0iekIojOAxeXgcQdyirF/kr1rgGGs
BDxs4cfeI5kLzxdsO+ezRTIzDLKNq52cHeu9EYEP4Bdi8/09Xt3kEPcaKoD2t8+z
KjsE2NhrDjQghqr8GouCgGcbMS2d+eFRrT8i+vM2pSy7/EF1sVQ21C3Pw7tzxlIe
tArshmPUVsEVbourdwYWpokjm7WdoKAs4Tol2zdz6Nx76u2QAnYHFSPbFPbFUOEU
7Il/Jy3FQQYMywjdK7Ie2NRM69k1NV6Wk3lNubheVdyFZkYg0y8izNvkT2gQAR5Q
SOnod0nIU5PhVD1k1mUBFZqYJbLl4XmY6yUA4NNtHmQgRwAzZKZtSe7N29ptl33U
JrEl1IvEH/UuOhxs0LOmrU9/tIgi/VS7b1lv4zsn4Lyt2ooYDl1WKmUZcnO0p8bX
kGBY6Zw2Uz+ytuMiTsL3YcnWMEqVvpJwSnPxm3AIj0WCl1T7+D9JRQ3Sv+5Ur5OG
CH7IdVyHXl2qE/VqMJq0yMeXHIdYd78E/krV8wrdkahQ8oE0+qtYgmCm3sSEO+ch
OYeWt1bTxwNjSBdNfTyT9BkW1sPQvto0hni7lrtRB+1FdFFnqRXGXQwRFKKstrgh
EYNuvc4d+x/wVOKXQSvU4YlMCK2IUldIxYBF0ZcL8YgGLnIAK4tB4TVaEOEgNxjV
h0HyBC+Gz4Wai3nDIaUkHr6UuPnxoOvCWtxDlQmI8nnHoiXMQgPRHhal3aSLz65I
RefaSPH7pHGAw7Hu1I3M0XiHAGHbmPxx/qe99OWtG8qhmJmkO2PXu2RwCE7jOAbc
cHTyhQ2WP/7O1om6H0vxJ7HHDbdlM5ZvAe/QPytsJz27iEacb4Tcni1zLnhPe6uD
Bp6OMtP0PveIncAvmoLq5qMUv8gvfE4QE7T1tb2mvf9vtsXs0QrUs4b9vPlczqQ4
niEHSgXjizbykMv84R7suC0w6WlQSgwkUAiHOsZfePGuJDgLD1DHpzpWmtCame5T
FifZOl/OILQm7QP9wYHTcG8ATyV4hWuRm3AI0FbIpppojHdntps75YOtxzUsEXRh
UdXMWWaGfwrhVbZGlJYkN//DrPpWHG4Sm0Shrw5yzmOr3rxMOfbz1g8QXw9EZtcM
Mz5FjmhAcwkekulBZ3EtUAySEEFzRxAg10kuvep09sGzqRlxwfxGazoeL0VvY7ul
Xb46SD9ZJDFXcmS5/ocN6WGoNleuin4IFeR6Sf1MNfL/jNm8HqQeA/RwMAWF6Wlc
aS/J6FfW731GnimRlz5AOqIiFXIL31rxUu+sPCA3VMJLrDwUGP0latPHTzajCYgP
eZvxBOXXAyqOX5AppFVea0+D/Wr1nYfEZp3uX4gA2nAMP2U+6+9mr7jGF7p0iEpK
6LhfPN9K+J9yJyfVAiXe7NexEOvTtWbDYWDCHO7K6VKufZiKZtt26r7FOOGCQV/l
PeoiusJ4nsSh+gDnk7jSVsDXeTIJ3+Ck8ckmZPlPd62F6hm3fCZ42b1TCe/ApgL9
Mtidqk+YGIngHsGuc4UMtMhFT3Wz8NobX++SDpTB98yETua6IhI9FbaYbECpicHO
f/9zeq30xIlm82nGbd9BrMEEMdVqv9IAOY0RRIHzLa+wXGaBHEjkwAm/t9Cqm2Yw
CVj89Agr0XMzjyBgicVkLZiSCnd7QQ2eyKchrSrsY3znXZXO9WWeNxieSkta/Bel
axNd6AiE/c6Zhm1CJ6hja3HuR2zkqCRYHsrjl8FuBhA94nS+9u8OVJYJtDB/dvzu
NLMPRK8cjE4rEs81s8lZLFDt2hf4esomaTCc2hb/QscaASIryGDPZkzu254bG6HQ
3RyiFTqnx+oosBmXKi788zzSrR3ogtBjfopgDxPxx7uEcVCRN3ruawGh46qLH66C
HxPjTLAu3m6hlTfC/VfsSrWJcAbp9r33s/pBTOBvG/LdXXTtVxEgB5YUpz2ENt+F
N3LGRtjo/StdJDqDAYffBvDNmXbDOl9C78lQolC/PIO8mYr8YCMldBeLBx8Btb9Z
F9Sz8dJtkyMIZkWJHHcp2TCJUdYuDYhkhUe/b+CxuHG1p3epYBJqpgPcPfY4JxHd
tms159qtJdqc/mcsbaR9XljLlpjhPZ7OU2907Vc8zXsxe9XXnnBNT27OlmcOtMn7
RpJVrrBhbWgaQFh7mYgxbnuFxhERiQ1EcaxI8Oh3t5CDNO0s6/3vtf1WjgMPyWKf
qxzGZvbE2f4mbxZF28dqn6lUTNYcQwtilp3BmY+Y9ubx7WfWQ5ON3smFU2mvQ959
66Ti3+o9SzYi7gKxPQYlbGBc3pEhRzJqx6FVLv8g4wODmAJbILG6NGfRmenAlwzn
ReRyz4IesSO8nh01zupJAi/ueW5/thKpDvltapTTYLIreT251XxNaR1ERJbvq6n5
aYpcpWU0nJHBpmhnDUG9QhzI/xL+/nbB0mQcg0y/5UsDHKCPLijLlkz94Q+iL19R
GtujEB8SewTJcvuaZpg8N2WBoTHsstnvO10pC7O2jsTtFqz9+GU7LuOB9O0hC84s
cGa1nwkD5E1tvIitDYSR9O0TbrVIV11edjkfwsnDgYIxYT8SMe0rbKnM0nGW0E7O
Vev56iONfOKxOyePRIO/qLMp+hkbB/knLM4zAwi8XD0LN7GsnEeR3bS0nXm1W36t
juyV2APuncwCLWm6rcFrREFHZYTY9RZj/RirOKxa0VuAJSZ0uqlxbPs3Lj3HY+fW
Y/4I7kfvCWEQo4vIRVX3CLheFXSuBB9sgkXi0lgDvT3g54ywF4/gwsTJNtqg+cEh
l5cE4rGM/k1ZgZEeEc8I44LZtbLgHDpV9av0/omRszwKMRhmA+BYAvGdijO5jxEl
QISgbj3UXPOIAiFi8RKg3dpaWaoI63oNsykeakTedf5F31dY+3WPvpJrF86X93xB
OBL/9+MGTxm+BTAPbJhiz4LE1ysL9u4w84ciGcjTFfLA/ymd7pSHHYyRQ/1pN9gS
eZCcrH+XCWAwqRo7AYxc3a45uYTrtzOYCf6Pkg4TQC1l9KlarMM68EuGuhsQKr1g
LHZu7EN1QbiBM6815eyKdUwC/sSgJ94sFwCm4RzJeAlSIBKAOnqIDzz6yA9R1Kap
LK+lcVe2sFxM/4APuzAPeDxu4CQagBG0s0hgs+Ai4nLJm2EottTkVX4lmRSPh1iW
Lt5a4IM+GIN5YBS4Vf8dnVcuIXbXSzpq/QasvX4G8NiqvVnKTOMF0pWbkPiSIqVQ
yS7WwJEh3GJurG1SQQLc5qhiuwimTS1eEoaOjuXN5GRs8v/Z/X0EQ/tDIHm2XWK4
R89PEY0MpZ70wVOGhrmzmFqqREE+w27bo2yz+l2ah4CM2bqUFMqWZ5Ctl40XnnQs
ojXy4QfmT7OPOLswvM7Zv2aEfljeKTatXdzUh/wG1ro5AkG1lbhL2DdxiRTHusi5
6IvQsWMqQxDWdMk3VpBXOQi+VQFxtz18oYu9glxSr+BTkrugpDPtOrFy7YNeYZXF
LML5f46pvjOme0BK3aiIEp5ZbM7M4VKbNPzD/8QoZ1V88r72zhECog7xBWW4q2HH
M/nWt0hbRp1n4VIA7JEbtxWyr2dmxumtLoNoT4LKZw7f6n+Btpt7Q0DL3MNIolIp
frEofqiFQ+dzaB8lHm6cUzIPKRSNZKkG9aM1kc3DbyGlDwOdGEI8mPgKPpfwQne6
AWxPw47nKcMcxvxqo3BAVm7sUO2JVHHU6FFIH8TPSWN/AipN5uccwHedZ9Xqz525
WTZocKhvymwEgfJDeVOBEAW5SNlrL6/wj1Qa6T78WWyPeNLqJKTmXjE2lqvzhLX3
Oiqk76yxtcECpqaFxfOTP6UZfl2+W6aMKTmohnQG26Je9AcNKVjFillkfBNS44V5
MGl/GtMVIGpFq7OWGDFumAc8awNyI6ga6bFVKW9CDF+uWK+ihyGZBp7kAw1vHrXB
2lh9r37DVFZuBgCiSE9SaESsPfcJERT6Vu/ETxSAwojLJ4snwX5lukhlzRjSS/TH
HnVYVn5DX/uOteEOM7WRzdRnd79G+/CoVShCBnBpCoQGc3PjCu2JNEIP+eEEu8Mp
QYzP0CYoSgPO5csXx5oxuCUxLRNTtthSDPz3sWfjd5AMk4erVabKRQwbEgh0cP6I
i+IKJ8rk7JizNGA9V0SsU1QkkIBBaNYAdf3JxJ6JsWUIpKRQbkO45vdrMhvSh6ri
WLy0RsoFo5Ah1TKgo7io+oszcjnwlJdz+t1toFZV+reDWtVWV0zsU9x4N/6Fn5Nd
rxvCpMHkH0PQ0y0lKb1AOSe2If6vATvASft2Rndo+FBx+zI/orN+e7zjfPm3SNBO
IHoR3zulgeAwlp80s3MU4GNoYUL9gVEN4G5Vno5EEANYVuV5w+2rC12knwhSgR4F
5kheXOCnYnIwwosSN0AIBZa2ALEQ2v+0bVUrBx15DYAwQRNLNHrX5aYGfw4J7zQ1
Gm6muRdxvpd1b++C0uOMhRmchDmCOy3d9WRev5wipGM6KZk7Y/1YRpUccRK1/Nh4
8PrM+67y4Ov/LnkSmEiyBk+YWw44vi+7QNXlz3b3MglR3zcyfKlATl6z18NlYccq
jlywbbsEU8kH6SPT5YPFPUonzqNb6EaF0nhDFDxhVHBimzv27+ygDahCAy7gPoYr
fHfw/ExiQDW5dqX/m+SGP6wmljp2I67mqFj92WkAg82ji/txM2BJRQ0gtPPh1f2L
0ykf0Velyy4hvZMAUxrzBJUaXSjdDmj2YGK7u7QCel8pfVzHGTwZ5lVgNyEyhU1j
l7KrYkizQJpScN6SALrwCecrHB+XAHIHLcLrKOQR+aGKxjc+PpGaJoQ3Aa/fu7y+
ODQKppxxOQiNPppuXxHJgJyAb6kuC704n4ApkBnUht62G3PlnEW2Et0CqtLD2elZ
jjABB30jX8amf0PxsctAY+dcfmehetB30nrDaVakYjt4LSU9+7cKA9bj6Lfmlwnr
0Bh3Yh/XrjLoBxUHTNL8UGzKQwxIABg9rhTzKmje0H7b3CLdjngZe/okXfQym1T7
1PcPgTb0PebZ1btpnZfoBzvYBNgUiwwP1srLLhDxDfeLIyY1twFpjQExv0kiSEY/
FoioRIsVYwKrBB8IY/S7H0pwgvPd7CKyF1DuPkpatKfabPj8wU6h4LOpKMKNXOKt
8awC0ufTNzz1am+jg+z5T6zUbxIEygasj7m4WLy4V7FXyBrxnZKqCXJUVkjNKaLc
aH2Rw5E4p31Oa7OAIMHvm/IJo5w2H029SfzTForC7rZsTxbLFMmZTta0dT5c8754
UFipGN8b9PSJ6dIsWPPXfIy546IIowcB0dxskzdN77C/vJCf2YdJiwVTm2UrRKGw
bIW2bB06jMKy03nPCbdeoJHQ/bCl9RM5Js9o7Qn4NVp8XIPeAC3ndMVL/7t2nAqk
46T744lGgo/XWmiDiBpU1LJNuUfBtybkN6je8FtBoN3+B8JCa0AwDINKJQhFyHYX
1BWITlgDU646QgubnaaBDdRVdnGAFPoT6MIjQIACTFvj5dZUUhtnTgFrmQWxjgEl
J6W3vtZE0VxiP4a0nb9VXvsSGfoju571m8mFM3LMFnPUxD6ukCKWvoHfT7pYbHZD
HV7g5uduO19F8EJ0v8ZwJ36C/mBkVEG1ZF20nmTDg9fxPqFpcBM43d527NQ3p1Md
+w16Vht1unvCOTLZOAXfJ/S+faXxKU5nyhmIVskPS18i7WYKeNXS44h7dpMWNaQV
Oi6mjEt6jS3Ku55MECTpaFvjr4JSWuF8yMhDGVYPzlgtN6daS2epUgnLIANkszO6
U3xJA7btBpYIvNd2oSoGBDRjNT5a5D3yYUJodLwWeFU4QZoni4EIFUTIXuUQ8DBz
39nHXc2jYNy4ATOuSZb0abF5hWqV4PLSm3fd1Y4HOOIrbzoyAGXZBl6QmIqgzruB
VOA85Fa2YDXvJVOwFQV6l4i8w8FH2kCFETInXbNongMoz572UvjQcrgA5ZFcmbxA
4VVo/8hTWzqtRM6Jb7EKmdH14pKY8mIv+ujhXggZsHjVtLjXWla3gciHZAajRgpV
2chT4ffahr0XDzAyXZtDVo2+eThSi3cEbZHukC0LjTvb55H6vdtHM5Q+GuA9MKNE
F4ICFRsJlhVtlrDXGkNkbgb9Fl5cMVD82NYg5h09Ix3YYCASlRz1vkinIYOWHbfX
heOO5Y8XoheOskQz/2c0uYsi/POqPV98aKh7in2nMC4pEasW4IgblFGMnyVnBQGF
Bv0+8Z3hsl/wIBDYTtQGH0QyQg6Fbmyr1zxDYYqRqTzp6PeblwcBWgRONsNEYjVi
1N60CUbWkXVypIR/Ubcev0leSo77LBybcvPUwlJcfayHmm5jT1Rkt6t7vBQzCmc3
+slL7PK1EnZ9dXCbLVSe6RZC533TqvRMa+qB4pBR2Ha6nb+glWJpaR4RJ140B64y
2fqluTub+tUeSVOpOq/e4+SxUJ+q7My9XDbiBfelSi5A95pEJTv85CMjXWihstSS
ISSl6YKRNXBVVIpxJQQmOUJR9e9c1WP7RGMD932EmD95B/PPo+igLXg5b6b5zHah
6Ie4y4ux+cxdMjvKaJM1w2pMg1p+buJPhsh3YmEp5gpbOVTBZDNO+nbEnmQIu6hI
qJWfVN5NmlDoHmiNOdc9vLxc/b15PUHRs6+XTCGU5FjAc+vql/nj04Z51GlwRLyB
2NqgI3JhFvzKtc7PgNqLZFW2rENzGjonMpn6EhoQ/UN/zSPRClKw3Pw2C+7tjAro
KJ7jG0HE0apyZJNAJDNE5QMDjGT1Nn4H6Ma3frviruuVri4ioKjqCQPsL8xoZIZo
YOtw7McmJJ7i1gZHL+kkHMNVUftStcyPWtGXM+EFhO4NlT7q/JUe/gXHfdVXE5zV
WDKUdBIqMSMck+KP7YHYyG9lXEQAf+deTu4gOIXaPW5tKTD5AFDzS7F8YonWLpI+
vEWJdo6Cs8LBCemB/AfVJaAbY/+jZkFDcTq/inqVYL1yX7KLamb/h04tkk8Qj1Et
MryprrJEZBiz8mI3+2vYtnBp3h6znQ+H/E4scbdSGO+Qznl9eABmQRS2vjcE5i0L
haHfzovPCMKkllScW3kiFBY6kxnAKQS84vS5mJmmNwwLsVrAmMss5d1YO8WTh5Ao
qg+AaQ0bUvMDx1jVW3wIMstT1Fk1EjZO76GKT8XUy5oa30NID0zHZeKbcvFAjlcI
6Fvvoeszcdarg9fTftO6HvEx/Pd0SuzHdl/ifJEl+NhOm0gPsEXSToqvhJ9rf2o+
HBgAbzoId9Qr+FHn8DYSp3CrwX01gesKuLqbFrf0k1IKLOl/6iSpkU437IADQH8Y
4WrDlZlnNNgGjryuJFSwfcxtXy68Qy6mcNMHqgXQxzZoxxaufnQ6pQnwkh1A/QPl
MmPOfbX8njjkLa7C55rtjsa2JZqT2KllOiG4tS1mCSVUzSR3S8+04X57lPfNU679
9OJ8/hv7oTJ+xdme8HynumdPH3dFSAKwwk9dYsDvhBXxXs4JAoz1p59ETDquccTm
ZS54nC9AxtQ/rhvdRMsP/qxcnQ6PlCipIrd6iQ8+PFib0KJt9+AizPGcMQ13l8Ot
AEncEEuC/jpXwx8sMBSHcoj7B3MYX8fpbQzTySqfnGjsunG5DOSzrnU10VVEnTFB
LqWiV53toa+dKwzaNUBdLbeYLuD6O6gipE2iar3bP2LALg6DAc4lFughU97oKXBh
2ThjEdINF6WtJG9IzoH9/MCcX1/T2xPsTA0v09wl0OxkGwDZhBEzH8RRTZj4/ueq
Z25sbzZzyTHHHesh1m4SbBz1rBNOwF2dq7ADdsyELcGUDPDD1UJq6dhOVAnSilzl
c+DMLk+E1NQ+WNzU5+gb+CKmtynElHmMid/JGZZ6FCvX2ePzXGZiDDjQcQBlSE/W
qzofSZowpT8n17l5Yn9/wFJGkZzXJIZAPuNkPHPZdVkyiXjRNKU7NkNs2JxIkiap
su/Om52IXenAGmdUAHJKcsDeeTr9NeVLnRvQ3y4o30K6c/CIlaVDhAUcxv9n5waS
9G6EppIxfbFheTOGtLwG0HD1LLaNBCeIflbl7xuBp7iV3ezgiCIIc+VAf8YZTyVr
oAHTO7gdQgwb3o/KWfyAwdD4UmFT+Gg+VbJnLlRzWX6+iGxBCDUu8nZCr9ijcczl
lAYlPNvWDX9wIvh7Maf1iF5RN03OEBQmcINFx63zx9VCa4HqiN/2DtYAm9EtZ/k2
BQMjAeN2yu/QyojLJ4yUhZ3IOA59OG5lBtQsYWL0tu7DU0vHeGd89evC96xQD97V
bOZ2Typ2DUkNy5vJxKr3Y3sOn85JyBxN97V7/w5JbF9IYFr4WOMC23RUogKd5exC
EwrkF6eNjbQXQyX1p7hQcpn5HNdz34kPQH+herHIoKNeo6SBvzcpBiSlIb9QhfLn
1WYFbvecObzwehaT94VKb7Y+Qev9ubwJ2RAHTObAImjVTvdN0ZXxItQG/rZALJvP
iCnXi1tN+nHBk4vXorxcSg6k/6JLAtpXBdfufTJHlud/4wBuJnIxeyoL9sn6ONiz
Ft0H9DZbLc9ikTsg9RWCSYU87kFyZP/M0ZZS6hEP1zzzY0l3E0eBEf2aGNESE8/J
aOXiOSyjA29TuOZWtlLZa/zIJ6N/r14C9z4aUY7TJcCY9Q7z7gf9FZCT5Q7/gXSh
oxz3mpi9w4/kuOjfXb0P1m8NHZjelV1UBeimeBl2c1pBCBdbUktkB9GLLcOy/nSI
uQ+mRLBDOzdGKDNyxJ4v1zlu5w5iZZde+XkghUJD4iKz+GabZTfYDuF/CveaamYH
2anKmByEyXsF9ZkVqtShBidfJIRovJI4zsCDUqaVY3a7LezZb7W3h+gTZrVWUH1c
eVEBYmYr5E8viN76UIITxUMEIGFHKJ32fCS///R5pyGT13iCOLc7cgSoXDOfhlJU
zC8Mz/S8L0iaASXql07CjDYePNI7jRF0ELn9aDslZjbJHLay1v10JJpj/WZFYABW
GJXad5InGMpcEomozDHU9cf/s7Ua4Hg/+EK+8jdZ9ZJJif+mXXeLM/dO7H0aCFdw
lOX3Xk8kFFzSs94c663pLcgBx01yKPTeCkiAUVsOTRrrrxihLm6P0bsE9vUyfDWC
oj7cQxfqr0XSlXaLE6u9U6alQ9jgl7wAqjkHIQMiXrJD07LPeM6WYJ1XShqMQ9lT
Ga9LImfVKUdhPJWBU6aX+NmqXZG0v8fqWwcd3aW5rZwkN6tzxuYSm2PfW0wH/Cnj
r5F3OOUQIYKgeBx8Cbpdaa27r5fKUAV/p5kjm9VDLDcY107613244UWifvNJeoWx
I4irAU8OTQSMBorKt668v5z7oS7ylTyIFzOwWpLRgP6yksdNb1BsrJb1OPnO9Bb2
vlyv5OyoZzBDCm3uSeNquKrNVK0zxwG8hScABJjT3+xSxFWOc4tXYGYm+X5f03zy
kU1IDFKYlFm09sZn7zivqqWZdUuvAWHaOjcVWWs4YciO+7W/oQABQ6ho4buTMWhp
7VpZq8y+ck3W2oRLZdhDXLSqAbXxRm9LqIm69n5tL5PX4t0xkmYMupB++XeM/BSP
A91HieSEo6Nk+rY4s1sBJ68y2o7/u/0a1oqtxjfq1AOXEhp24i488D8wSA8Ttg+o
qaUVstGY7cE0GJ2q3HaG5ibIGU3FP7PnzfrSSaUR9ll3Ekxwnr9bG28Kyz36tsnV
9bI+pfR0bIhuZ15mKHJMfkxH+3jn8FttV1a21YO30UkcghaK4rz+SXkodub09TwJ
XIJW9r84JJNciUjcbpsmbyDyDdKLAcdA3v1Qy1F231r7Lb7pgKT6xVcgHWH1+ktR
Gff06q1b6uoZh8nczoDVMGMRgaqginhn09+drTOqmEstaAnt/fnbyJLRMG7Nk0bM
RJSsZ0Jbt8+ZMNkTD7UWBwfFALx6MyYBkgtgyQXtnbQv7PFYaq1IL0+2NL7vQVsp
vfZSTvnro+TRHlTAlvwG2ac0r4E5FkLwu/paqbyBqzrscRkqgxXLFVnOF8+jC/8J
E+Gm0Q+z5jM5fGeDZX/xiPxlxg7oPdSRFZoztlbjhKWkVLE0PcxOIjsyVapHybB1
X+eK8sWYKEWs8DIDUZD0dNLLUZq9z4MCWJvb0k16HlpHlCE34c7Zst43KntjOaKx
WIQ5s3QVTXlq7VNV/6gwWKlmzglGFR/4oIttiUtQ1qD5iMU+BL/5LsMXPPmVQtRH
DZIuzroBh7bPkjh7SduHJO7GK5t2qmekVQIgtoPAiIgeszSWOTbvx0WGQUJ6ww9f
AkwABVeOoAlKB/jYYqJpp2euMtKDZ4209n9ji5+nsqzLzJKeiB6sA1jcxdIxcMKM
7v5rCRU91oyJRYofdGlrztbaWRDB8yYswYg9m8FB4IzPHCkUoDOEDss+sQAWj3Kb
7zoMOLiOUyE5b+WFaz0S2XX/np5Kk7BrVBKbEvDvr1ZgwYsiaWxsl4ckoc3xe23I
+ad+Y1kksmwysdJ1rccRpKMaFE0akzf1BFoYeCTnQYqz3Yfo02dKPitVJ/TLcdxS
6P/mHivxBTAlPtznnZkyJRVWQUDwK2JQS67DUoC/BecAZITucFkagF056ObklGPs
0JEhIZVZmbvTq5NKPn4/+xze/w/UZzWuU7veX8Oc5QTWbbWOH2LTX25ksm/vxanW
JJ042AjExwEPCG76uWvsix/KPcjZ3a3kowOXlhgXt7aWQOrFAky32zNB2yJ3GpaC
u+IQjf+k+fiNAk7xeRpXN2EtzOHaM33EbbOR9gfUYPZz0e+gZvxzYFTrCGWP067/
FNcZkyoqC/QnI409Z59Xp4dWdDXWQVRJj+CPzYTeyCeveSgrbrfa6zUbZ8uhmHdp
/es2XW8HnMO1oJnE3uRzjXrDOhVgTp8lgJTBUWVKftGNs631aeOq4aRIhuNZrdUp
7mYASQKcXeMO/OLppQ3kGIVQVIjPt1jEqY9tbXzAx+Z+naW2Af0cXOgeph0f5uo0
3wEBtye9hIKXVB2HohhQmlsQjp8rQCEKfsHRTmzq/2Lp6uLifZ+JsLnsFOLk2TsJ
irf3vWuE/hQrWm/OUrzi0tUWo9nw1kHgNCdw89S5vTogfC53qVrwu4iH+gi6IEo+
StlYyuziN+loOUFsReqmytkSBGDxoaCumZ9Lpw1ZE/5n1SniDgIlebBsAkxyv+a8
RcKR1fn7aXIU1e01Z12nYH+7rQ5nuryO+hKp+FK43NVHC9K1sX6nUEqECLl13bTl
PKrM4EThbLiWkdAK04KM7z4preoTCxK5beoSmq1tDX9BaYzkW5QLsrv/xtvG0rVF
KezBVnQ8xnLj2oJ8nBmKrAJczSyBtutZjFJhVjkvLDInZdGwb/3nbTIq9MsImEbN
HHEl4t1WRV23w4x1bS8pnsXfEVtIqDsWjdMqJfQApawgiYz1YJho8BSArgzHYN4l
j3u2ZTIbxU6JmSafaYwQnuOolPMxGUb1n5RNLOwPh7wb+DXuaqxN1/TtkeD5R8mm
ND6GK/rIbsc8CGImgrDGw1+yI2zKffR1NKPQwDW89gfN/m5ZL1+Uh6JbND43GIKZ
WJFbBCufLgJRK9Pjk1duYyfuQ10fgIiJCWT0iGljW5TqaWsTekwHxUlqTtRa/qsL
hYGZYgEOg7RCiOUDo47yaswT9mIWlcy175agBs2bZaX5uKYoltwoCA5/4HRC/mgR
4zZUVVWLv//JyidNk03mRWDn/C9d237OA/vL5T93GZvyKn7AnACphg0H3ZXFONQI
VqO2OUJIY1QHLh9wCNu7Tk5LgW/jJp8OMklKHkcAOsEytZZuHJgSr/e/3b6ssQfW
X8OqcEWyrq9froVDXBL/xhyV4xU4/q43p9tkVa4hzIzRPx2kU9F0KFF+dGNblHpV
mLgj5OhU1Y468wTGwKDdhqTflSP1Mwh+03JQC1eSNaFiwcembHHpDWbiyXNdWoYU
0Lc4qAibC/h9LFT/jJUp5gm59p8cBRJWzsGFcNU/PBQOCXcy1ItYzVvk222xvPK5
5zNbVewijOWPRo8ZHe+szRMltQ+JInrk0mvU4oPC1cLSR51JFMCib4FoqhpyFVVS
2tjgiRhnO32foPSsBc+1AJQpZeLz1tlcxz1Vkcb8SWqNRSVMcX1dCSH4oOomG/DR
d2G7tUzl7uTaGUJMxaVBNr31r1TYB/W+OXQYP8NMk/gvtjy3w0UUCjMOgZ2Ic4Vh
WP/8AoxZvwBd/nrie+oczgLIBHVf33HhtFkzjJXgGj5TJPYRB1A/ZQNi/afNNRdF
6xjkQMVck9XUSjj6vLmOCQttNODHqiGjxoQnVt1NlRjcep2l74QYh52R5+Bnum6b
hOirSnIMhPAUl32YvnUdPjDDx4rAmu8pcy6pXeeYMNUjkUfayXK7fp7YJoasZYWr
BvWPK6EQB9QScLSlMdHtPNFPsxpyCzydTa8IWOpIOGG/xjgVBtnOlSNg1+NArAVz
gYMpxRpZboMwuBKKxGcC4cbR1Z8NTAqwKUOIMCObqq7dqbMgFtL9YWYQ+uR8DcLU
QpCcvX+JOZlxYR3qZGa/iMA2wQlUf2CHYJL+ToK8e8/V9Jc96sCSppGDu+OoiNnR
RblcOGCnGLXTKlV5Fe1li3ZbeajmutWJrfLlY6xH0RU+NMgyVnuIJSza8DCc5c2V
O7R71tqsfApFWBEI0cjmnL+oIAB6HtGs7H6FqGnlLHMxbikVJ82zi+b6pZFClgym
Tah5Tg62JZnGWPcCZ4T4Sn+YMExnGORwhDeKAypK7Q4gKlV91Y86s2EhOQ5B5qpC
l/dz4SqPeKoGrUTFJQBMZ6rdv3LzMt9E3fU1wzhR8noPvOhAtkaWogp+raAdQRtv
esFS08EfjLRHjy9aWwawNLLA2GyiRBAUcubNd5uelRzWDensLzp14PFGSNJCm+9E
JI3M0KJljuHITzkFegib4Z/ftcvIl7zquVVvD2TzD4ISGid+t30e2BOcapWWm0ax
kvsN1FwbVnTbhwtJVJu58ttniSyxQKI/+D/Y3BCxEdcs/wOUuhd94Ri9ki7veELl
4LJI6aBe3Xhphpaa1QyORYQ6WIQ6WtwouY40oWeVXPtKbxQ2FN/4HXQREssqs8rd
Esl8mfgogkCu8elX4Xv1ig7Z4cfYnv63XA+Z1tnBjQQxou8R+mkTViOd4hI9Y6Mw
wCgRd4YzwX0pU3nDoHkWesfI0cxNKg/3SdrZWLgatWBj7mvePw4oLlHSuP9udi4j
0SDeO2vWRASAzuiXjSSUabc2LZ9Z6Gq0xCFyjWavYp3OcZyYtOJRG8t0XEkaVXqx
xOw4JXm4q3Hv9C698GY++Mwmcf9hmimp6lidGVYcpwZ6LgVppZ4YrIqTzPeJSZsI
i2FURaMvbbdjIboBB8DJgo4KRMXREPPv7evGCa3DlvN+eFEqvVn+/5U1oOp/W/iD
bdZ6yT+oVtqCwxvH0i+BbvC1g0q2a6dz9zKvan5t2VNIumZ0qv2K7OAjS+dlFmmT
U6nZiUsiI312IJtaEi2CzdHMe94TrJB0OPUcJn/oU7yF+FOwL5utFGwhXSCPVNrp
3mkbAnTPhqb8wB+MSETC2Bc0DlAl9AvHD784Z+02WWVM5NAhnnL7n9zqu5xFpU7Z
c8xpbwo674/1V7Wf7DrriF7hJN4qzdzBq1DLTfR5JBL0FDyzeXyLa6BTdiIzsbF7
KoNZCIJH1xJGC7UFiFolpDHXv01zVmv0z3PZeoNDPP+YyDWPAaUk8nreRQIc9P+F
zSAW7xfgcf7SkocXLAxZFsmELzBP2EpnOwnCXtIof9tDjPfH0sZQh4lJmabLvLLx
qbPCJrxfSpJ5u9lsu6jFlKTtsPhjpF2SckZdd+5vjKzh+KkuYqpfdfF70kOdW1w+
qXkscZd39wZ4MFQU93RB46f/Do/nyYJR5878dDlFroXqAwO2VLkVGmiVESDJ2sIY
EhyPL6kQIyWntrzctN3VmXiE0XqZodXoEhRoc+POAiFr/hFBPSRTb0en1BVQG9mT
fQCaDI2YTMbtCHBVFpEpkocnT1mC83MU1S8vTXaQs+l6IlYSx2VckqYhF4Fji8GO
Wo8oO3DtyZTuM/sGEKm91zCJYUc1F/UY/9Tvc/Ef3LfFRadQLcWCVZHqf5HudBp0
DPzxHSKifa/Wjm3LPE85YaXGGvDCFalsFjnTYYGKxL5MWw5QE/J1jynMgrc739xl
JjDbrCAO3DMdW/ZZbGgGG9vGXo0GdEifjefhod6V2WuVOuj+kqs+xvWsOeY9qIqh
3sx+eFYCKWEMAwqCXhCDFcydc3u+PfrHmPo/4yGlQwD4husPOSpZVwX0Dbr/F1GW
z/sOuONUZ/PIg736fQj/1TlH/9siKWjBPlKyG7aojFyxFHAX63dqJNyVTZT67JKO
aQaPkt3a3NSZIOIDvwkYRrh1KeB5Ns2LVmCw+gFv5TfSeVzCP7ydPoE6/hVG/86P
RNw+znwJ2kLBJ96ojuqtFrtavAEfNOQ2RJ584XSD6TAjlgo3LHgpDYhCj+vtA9Yp
FMFqnH6izBecKDYBTnr71nCM8HSvMdbNWeshg85kqW2LEqzxczts1Sb1T7NOIX3p
x0uWCH+2PeahmI0r7GoV0Kr92nlhEeMo+/zktoQQxj9h1OewawcNXT3Y+R5GBNAz
NVrG9I6oSIXcYeJvn05sGWCvBC3F2G7GKJJGjx45+BssRUiTeRqLXb+ODB/hThUu
idVmjyfqYomFZcEWQ0XaueiW8ydQWe1M7cpcwvkDgVZ1EUhPHHHf251eMCuQylNP
6BjVbxBl17N2Is8Wk5vDhUHxyir6VbAKpIINOhmSpeffqdYKqRzevHkN+NhB5OHu
0UzdG5d0EYiubzV33pvaRcJSXvX6AgH/r5Ao6CzIe7+pP1cLRX5sBu2xWZluv2bR
olu7xhSDgjMATqElmS02f4vi7WMuSLqJunL1x/aH6Ze5RV9CHNoZ6x19GNLsUQ6s
iF67awXAyId4R0/Ztlf3hl7FbhJEUOhNxRQPuwobTt0N6QT84T1mFX69h8ZWI2d2
LUNw+fj19aHb2jdgpZDtRIR4cvXF/LbCFf4LDDBIV2VB4QuOYdCOBKD4BeUNVJxu
eOOLSCEr6AGEX1viRe9l4F4C7v95ZOAWaBhxSQJh8bjGFzSkWaK+tjoFIFDP5crA
zHQ+9USGCw/jHcxyDAcxgbunOSPMfuJ6PEchT509+UdOL/tsOOL+P5wueraV2eb+
p6F+oKJLkGxcteKvaAR2OkP6y9WuHiJxq0PyvTDqrqBGrVX5VFJd6qKz7xeTYcV9
3sARDLvStJomnEC5NQ1ut7mo5OobXPcPLWYjZIXebNh2+40qOSDTs/Tvhr/dAhDZ
k+2nNU1Sx/EfRLcd0MA8DpEjuADSzdyFvzxkipog10Bcs45FwRvbNYzmqqZujicq
oPHOtT1ONv1kbRT7KSptVfxtLfuhGeKjtACobTF/nntcAiIUyyxoC0eRuYJbfaoI
nc4fuznSRyRdU6JzxWWdZ347AXoPJ6bL13OFnmKPyCre6kfW2BXEM3QrhoRWE6F0
HIMvoadqGOSUolzVCuQlcz6jkE0xdtHCMOVby6dmhmIqhK8a08OWHGh9/g+I7u17
z0i9LsVwQDG0wMrMZplo8OrcOa9idp8DiXPeo2qRdXqIuguHY0bq+zFUJi0GueMg
Xzihh+najjhZF+IJey1jEPcn7DBdN+8e/a0PJBtEQnVyZGQwtqBtoSDxQh5dxh3y
ZLsvsePCmXz4XHZjIxfSOwOBCrFNYidXS0Dx/93qLWaVJZE5QdqDEpYX2GEI8jE2
oetc5gZzMjYq9L6RQ+4WNf9HNNBCMv3cT/b1pSKH9UIfjK6p4m4hK2DYpt7ibH+0
ddj0Mwh2IKgph+41mFQO8nvDJV0L0Je5XOggwgMxjQwcvLT5+0eESfDMnIUyo4PT
OJrmhkKd0JA/u5uJiCBBLyH1cYMZtefuq7DBFGuc4PRFCPl1OjSKIKf2qXGnHCsQ
Wk9FUiPvw7RpTCMUGkd9M0b+/OnaVV9XqUlR+Bao4HO23EQ7aMiIQnI5ECEMco49
jxWdr/vc9rW7s71hHAyVAwNmDFErNppUzmFEEopcKsT2X13d431yEQ3hK/gI6jGv
MYivF1u9yiXKlF544mO3x3rEm/edM52jDRSVen0BjLtg9f9BV6pyI1VyrqfpKN4Q
YWTPMyybZsg5xAp6MCQPJhbC9I/Vq4FKOotaZeQC0w/uzVRdT0Pd6PWQ+GncUSoB
ZFCTZBP+svTzgODquPccg8IwGlm81lr1RxN2uT+rehq/iyKwvqomnxFO2Z4T8M2J
vL8RV15/tO7hOkSctl20zXZquslSke3d5ArkRhV+k9BHmUo1UOhGbee5AYBDcZZ/
KHKM/EPVtxHS2f9eDhpuxOmQWCzuKtJMr/xtfjfzHgFJlTHoUksIvhQZl9RxmCdm
adHPqhRXDbpXV9QnHoPqMR8tma6z7tZvc1MSukZYv0vjFRU1N5R5P1jy8nfB7aWn
uzFt2pZ7tBrL04VsON5e7HAoPnluUcfeNTow0cCuUHrqm7uwgFbXTkMfonM3r9K4
WpnmY6W92NXU1G8HaeAuHww/M1jRuTdIn1TDkXaemS8OkVm0n4Pl7a6TUjr4qnW7
sKrMwxzmsPKKYK4I3J7o37W0gYjJAngSV8nocLDmn+d0BXxTwOBAxcLeZsJAtHUW
mapP3EdafiJjSlPO6y+ea9jVAXNCSenZqbhwNzmOBlqJUZEyH5lq5X2nGMGRYh1S
xkhuvmPZ1C3BhD/HyZMPZVuPu49ka1ECrjDwEm0fRlXczf2CyWrKUh7Cb7zjatzB
A/g7P04PpBm/c6LCKZKLJTLvEIRjEC8niRxWezBWa0Xdltwk72ZEpl40f0a+hOKS
b/lz4UZ0vdmxreGkrxgySn0qMXNgXkzORgCRYWG9ZkKxJ6QEVKykFA0ZGB5hF6a0
H6AlYNjCAR67fiSjuy8qJgN6tNAM8qfjHy1ayep2V7xV3YnS8MY2xqt+fukqrBEo
xdrozIVSLp8RdydpdoU474WQCbm9nBTLk0TV32N+z+g91gNm0cWdZSWIgKp688jZ
+eqORF8ZgNfFOIrUXti3MFScdHfwzhOKy1lV/63JCAkkRTUtuZJidIlJc4isVjKG
I0JD6/ry9R+6XcBlpLv6wbR6s3kMBSZ5VxU3DDqNPQS/VbMkejR8ixTDtvB+T6nQ
ZGBaheOb6icnAGprMnR3epk6FqtfPEW6DPi8wzaEjWHclRoOLT+aY2gn8EH6859l
v7sYgmxaHpAmle6TbvWQ4SsrRzAn3nTyVbRJlDr0cCRcVGiQaXNuKKne8++77+/a
5oZ/2zDxUB5zfD2VHIRuANAQcMWewC0Zp8scCo6EVUf7GepQ0XCi4bnHl6nRFEob
GLbLrvv5JmaQgkix2/sw56EV0aMKBdbMUdVvosHOqkSj8jvOVRevx13NL5fOOLIr
i1Ze6gyVjHGOyMLv6tZW/WkpJwfV8oF6RQ+2xfsx0k3wkCJJ261H+H/NPH2qIfI3
hbDHhgoxu/T5xVCmH2hEC5x9GM47MWwZ6TFEMsZT7nsebUUPmQQ5nTwtl3gVFmKT
P8C1PoMDl3xuyZS8ZQ5Yp/ymca7qaesqTDARXYvXplg/+6VINKMNynVUwbS+ZtTQ
9myxR60hQLNAGeQ6/DMuhkpJqjEZETMlA1NsOLheJqhqobQSRZSHvlbZLN24gRC6
BQIJdZHYsK1gJdyX6qY2T0d/D4SDn9HLy8An5varIyiSDLu/ycYUf81TaHS41iew
j+2QI3Lia6bd4jBe0oVKrDMvAodg/pVwFLe0/zpf/xYTPGZ5CRITKn77axqhuDrg
l9WmOGvs76jcFhQbunogfQgNKFwIV4c5gBOl5mBcMIQ/YboAlitGXoxIn4NxJfOF
J+rf0xT4FB1NsejFobSbDpRw0yFZqaFBTe8TUlzYsy1k3G/bNvdaMB9Cvu/Pt/uK
m53CLTi6Mp9tnMNkEaERsNgLhC8ptvZRZ5dh1NiDhpZHFXpFfOcOi821d5FG7ywJ
b5SGGIZG5uHvwF3jBmr8JQggm8+5joh+SBWpe+J3zmy1CJrZsB/mifoI5b6gPnL2
aHLjXLTOpu9qDRz22IOc6dxot4UO2BBUdHOiScVatIngbfRIp/HO8Ewd2vZWU085
Nhw/vKMwCIzWrp3/opiJQ60wqLAIB0YQ4FlIthiHYeeg1DqG7qtmephFQ8+F/9yd
QIyCTtxJ1qvN6OOHDXtWdfIHmNV7mYKyw34rCUEIPt2t/U7AjF2wvvJchCQYO37p
gLk4Ah0PKx+kAL8/rENJ/0SRkUpihSMjiWYL77sEW4eYsU6o3ROtVnwI6YShOIii
G/5FSVnWfqQn+TomlXSVPHdUL9YJ9pF+inOluMbAVVGVozlif5EoyydUiKF2o4Mx
YjSrXzCegtsGylKt94WTm28sVGDwjg27Ikgrav14W0ey67rRTd7z2tVCQyKmPuPT
kqvioWYb/nVYXqg84Pw587GQ2W27rMciZwZO6qMMGX5DBt+RI4I3GvOV/b95SU5x
mDQ86ng9SNuCB+qfu1+x7/WtQ1KIQ0hp1dzO0h8D4My8BI9udAgs1Mpek3VjgvZ6
8rzw4/Wm9D7K1eeWagD+7ZJ1PF3YtcbqebDBnCZdMmrJIspy7BmAWrLVu7zJqP6D
J98cnwyFL4UgEXmHdg4XEd6D+GXdizalykh8JcM7pQZ7E7CzlEfJvHetQgDGh1tt
OTfBDPPR3Uvllp397oO6bdu2DKuzulmme8Fy63wUGu+V3gBf0ePkcGUsw3EW/Y+1
AVLgMO3JkqMqfrutqh1Fuf1SgEp5OYI+pbVr4SN4/RoTZDh0m5HBq0zzMCsBSTXo
Zd/uD6/te/5IDGzONj7md3NUX57DUVcLevodRVyGnblkblA2uoyHG5REYRyH8RZi
Ui30HTVDOxl10cQHosb2g8r1qkfN9LgiuWxodipV4+slv0RC3sM594d3Lz+b2x1a
QS4EGUtRbrUX8G8RUVUDcJH9jwOO+4GhAkFPQrgTb1iImiMsAkm/LijVljlL+Nvl
n7MD+rmNuP8oAh5pWeJMfPiIvkD9r3d09pzOK0Yqt40hM2vCeUEWs5b1zVMPpuAS
0aY7EI5+lCzuk1+YfM0idm2k68GtuNBfPnI1lLZ88OcfTD4lmrR2Nmy7pI1Q2F6R
pkSjHWbnjM19g1PbMdpsM2EoDs0cHEmQPWG8dQGrpCb6QBZgqaLyXfrU04oB6IIs
gX8r+WZuK2YOx1rMhMLZWdxexULlA6dezzb2yJsC2ZqJ310gRH5k0rGWpNShFxr9
+ZEtV2Ks9T7Jll3lfCoMfbv6dqV+5+ndmu3qBpcZp97exyy5bjhOeYw+huH64PdL
/FG2gkT/ip2ywqXOQ/cmh+5yGQyb5OA49jDcvdQ7B9OTf0L+XzBWaO1Sy8LVgCwB
vmcGWGGLXSmcbz5W9RBmftH/1VdIZqnztVMI4WDIrXChQ6zEp1ItK9/CKnSsYf5l
xE5MoMhOCBMUvPubFbnn8CvCiJbTxrB/ybZY5sL8FKQcwJXjQ+z0RF9oYgenCsf4
WCCsR52YyiTbqPAu6VNYWSG41xIL30m2PWUjv6qPbCo=

`pragma protect end_protected
