`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
EjK1mnWB3u0nBvBLwj5ZUAnLbBNKYGLtnyqg43kHJWyRqotLhKxJb1/+SQpgnq/s
FTYXY4RGKtJ1hFaEjPobiXrSs9UuIBEeEBdV64433cWBj6J19tDIS4HZ1PKm4T6s
h4TS2nyUqItMnPllpFZmjdGLstNjedrYXP0y2V3cA6M=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 1248), data_block
NfgfjiA1vCnZiZMYj2Frv5/RTw+Cpc+1J5hrmxiaTj7hMm27be7DWr+IRlsqpZFb
jwaEdNj7aIMr2U30vaF4V3JASATwIzB1K1wqylV95uqCDBk1/DsGFtujCjZStUgv
o2DwnidAJvYYYknhqxw6vVGMR57bJ4ZksdMv0fSljdLsTAJwjE922e76ESC3/E5r
2jUk0yKufogttttyEj1vwqBlxfVM991+/okoxCvY90lSJPZZfzXT8/nK3eqfACK2
1aoRhPsid71aOvS9x6iuZeUUchTZPDpAnyqw4rZEO3kpQQ6s8KhyjFUUbolbUu45
rvFR99QYTwwqDqipBmFKEIGBw9/lm7RsF18hQF2//2z9shgPY4f581VtNqYlloYR
GcEZ7swqtnIkjHAlD9wc2EuBY6dCteM6VdV3w2pJwOSKgoFVhajqV3AzLAQIEjh5
ctYKZKw8iYclZoWlDrz2+RkcZZI8N7CeJzqlUJlhKI7oI0+p+1ov3WkFOM9TCgWM
n7iy0NfryDXQ4CeY+TNjPhUDiNB6AisTQUX7I1AbOgrcZLVU2UjHQHeYSlW92+k5
7ZtnQMooiHYi1ngiNZlz+8Ss8pVK0c4DH2B/5AGGn5U3ecbgIy83eauQkrVcqfJo
SCXas7SQwp9kkyh3Vl4Z7OJNIIzWiKlFl0Pi219C3PmEG/5u/w1NIYgp3OwAQy4Z
37aU0a/1AeCx99F2pBd6Z6Y4+EgbipZVK5eJ5Up68GlohHbarIdlCRXkFYTM3Io3
P6qWupb3m6mf1k+sPjEMztRys2vi+ybK0aNXgAiy0DH9qNQdVkp7NXvWlEGvWTJ+
MeD1yCDo6MdMs7QbJF+HAo3HEcBkzZo0CxhQ4xkPmF+xYS9Xo26BOLyRSRSVkNU1
fo67u+nO2+Iomv2oQKHm3Ze2IvlEvhA/ZARMYYwvP/XQznsj6lmoahmLIwlz2f91
KLbaosqTJLA0KBRifo3Mt9SpiVS3pgUMsSKasySAzmxlueDrGhTwTMw+nlaDXp1X
lrNwM6pBmgwtoZZhUmVw6H5oTWUBVx7Nb3Ek+dI5hvqwG7n1RzC3pLpRLY9GeMRB
aG1ubL0TKhKNJjHs/Bl5Rj6oVFXPO8b8ULzfBnn5uatZMi36VaFbEBwTZBjYcm1X
BCGHptYRlpF/+vp/wX69iZ8f976aNObPB/ULznlXFWSd1t8EVSANWrK9PiScGFTV
5wYNt+rVSDRzVHi31k1GBZJLaMoPWMgCWbnJ1EVXvV8nUu0vvHchjRqEnbPGSqmd
m1ZsnfVUHR58obKVv+6GpOsI/D+YYcR4/HaJMZjhhyVJho0vA7Xfw5QtMumL5OvU
8HKUWaYxTaMabbsjJLoVpvbXjyud1QavTs9O+uQeghNE37bN8YLFAxPnB0coBZpr
C0bOCeSoJnlojhKkdOFhAiwvzt0AV3eWDX4kt7QIka96rLOMJQ+g1bI4J/c5nt6q
oCi/SQaE9ttDKew+SfuyqIcPN9hUfk8MWPAiDrk8itWDfijMyXulmQA1ACvHbkbk
i11ocPsvAkiLraDmEEW0NBX8fE45ECFCsh7khHdfi0bAxh8lgmONNPZdVseq/CjW
17jwvk1hjXHpqOSYvmeAXDdNMuJ6vm9Dls+q0xts5qkGkWQvbxG7ZQq6ObQJ6iWJ
`pragma protect end_protected
