`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
jFGJ29h96S/uwBkaI6xp8CruciTq5bLw2bkLi33KAMwcbnsZDrLpRJua7Ctx5cTN
GU6TmziVriWZPYIO9XcTq3QcJOusr/zfSVjSGE45RfLRn+BJJaSP62y1eYFskvWP
gGpmFTzepVEYmgejINhYYns+W0dsYva2kB49PMD5WBo=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 29440), data_block
xDn3mSwAWHRIzgxWOYBuTSjpvVh/0+8MEoNGxSvlj3MIvkuyHatt9XB7+szvEuhW
CXUiRkxRVtDaDpKNh2zYYg0O1GBOX8MfIcwWxlZUK+AiJwBc58+stoZNnEat31VM
/9u66hGbPrdT0aCfwtNbiJ7kga6hMI0V2A+wSS3ycgW46LCxxpH1wmehDK96Njih
YZEM/IqY47JL5ua96MpvRR0VdeBFdEPT96EFtM1Ov492FwSTVaN71Ny5r9hp2FhJ
kcYWRzvWlOommeWTtJMQcYusszP06UobW0iWIav8Vt3sc4cDOSadNcMiQboy8Ym6
1JZwB/pdejt+fc6I/CPKsyvwnGnba0FmJsUW7JQ/0oIiTWVS37Q5hmlmaUGcGqDi
Eb4GKXEvAvIbZOivgmuq+aesmd7qabSS6lS+iW02Ub3w2YHSqM6ZalWsN50ZuE4o
WE2VcQ1PzhgjmQWoGbWgPCwOtC6+zKKgHe/G6Uqc10C468Wc14qYOWOyN9NWDFB6
m7eTGioEr5zLSxlSftq2oiyA7a6n1HXmhnr85QXT0+DDhdN4LE5URvyFSLqCaqtX
TAZP0nEpOE84mKR2N+5sWTV8G5nsDEmZRScZmSR9k1HASYrZT5KSN25aZesDzcD1
nltMs6yOjja8mvEWGaolzT8cOAVQntRIIXmCwmTh1bMWqYKYn7L9jQZamu9ywew+
7In6MVXo02SB+yMlVG1LUkngLafupt2AkZjaNxgjPsIB8SKUR/5OCGt/Ydydh16r
i+1ALm2YhmefHcOevptvRZxx1PzP0Dk7Lhe4B5HUHxH7qJ5xeCLE4k0cF1VKE013
HLtnE36UFKK8fmz3f97+/gBDyAVCOrdOj5TbwuoLC1yI4tYaSnYUfNV1C1gw2x45
nRGi8W/mn92myBu8FvIfkZFZFn8YNP4u3f9TIrYwtQzt5bQs4OATCctq3UDfBN2y
Tdmetk9K4orulvf6D9aUkQAqtSyPTBTfrUDgcWPNDOZATtDonuInzHVJngaU+drp
vK1YhnA1BgbgGiyx4Z9/KVRpg0Mqmoa8+YkPIuohqYklz0EsjfWalt/CAFZ4AXLP
+dVVaddipn/V1GvXsJH1dVzK5n36lGk/i1M4Uye4IuViqm+31/IWECtYcIfRa7fU
ZVHlBtSU+MZNzxz6FZxat5Onz/Twrz3O/CD7I6d652oyE/uXvli+2zFRJdPR0MJZ
DLD66byCSG1YwDPTa4e/6B5e9EnCQ2/IyCmZ/R0pUcvcIFvlYGR6rDReGnEQV0/k
9Bw92TApJ/Y+PMpFxt/PeQ+bRRSO4CD30cWh7WOe2gUa5I2by18cdwvLipx/IKAk
5n7xsAc9fAxrlU1uxhRsMb+jQmaCMFahBGsLp9Z41byntb1Sn2NUd0tGzaApyv9n
j9JPvtDLQdWbYcf+5vT1tFdwnRzqrLBiU7jy8J1Lcy5T6iuZ3bQHqUr596bCBhGI
iSfcLZIatJfKjPFnVrrJ6h2Omq3uFR2JEyOH/E1wZZkYVdYB7Erd16BACVhWabRo
s20bRQMPeGomUPrcHqAgQXnxpV8ZLsZOMwlDG4Rn5rCiTYxqg5AONinAGZ/yMM7a
X8Nfu4PdrVrSM1LD5Ep/rXoLqRz4cKSd2QELStiZ8y+tQHiceMpGalVHt/BNd3e5
WxXk1x97bqUlwrS0/DMl+Xp7tS2JV36qMSF+b4tWCNU+xvJcgu85b7kPATXgJ07j
7LhQaaatbNKZraoQR9s99xdzyovmaVMuIH1RP3vSMx8qjifFHQ82webnFvD2SKNp
ymkkNqd8dW1+vsMQ5zBUfMuquwhXWJGNjB//XsktbaqZobcq62Uo3KfWspArRrRT
7w6IQjvVbQsKmaMxfc1p2DI2sYmahftRkJJvWdk1WynJ0/VX0gGZu+VEeuBrUsyf
RtY2rFdrh7BcMxzIIMg02xYSZvaKH0rhcxNci2nSpiprNv+fuUycGpZ51lpcazMO
gFsd4DNpUvfO1dKZhORi5F/kBrRnW5i4FPauySroAKv9nvqLDRlgQfAfhHVgSGu2
8PrgRg9f51xJbe3Yw0G7NfIzIlJA7uqygypNIzCPF+YPuCNAren2Pf6B4tY6VoPC
3eIYHUqQmVia9uxnb/nfR1KB7PXmAKc+CBtVXotQiPe4QuP0+3D6jumAXPom2Exy
5pxmuT4p8swUcIHeD7jpXiLu9ZY9GE6XDjqNF8SvUpWbat5VnBoUJxXRNZ6lux/P
7CKpxmu2zQJ32l+IlSeO6tBAZWWneScci8ch+Fg9FyDWJbysoxnavDPgDJj8dYzx
WlB0xqNZcis36AhrgMTEiLayB1QYyd4WKwlaq4A++PJhpFSV50FT1V/WdmwTQzvm
Iw7WtIqu0K0k6XN0wAQLJ6kINtTcpOJ7JwxrZ0T1e0O69+xBmHFHd0r7UQhgmbzS
YH4kd5ZeOmHUMTEWFxQDsLeLJ/ICP/Xo+zkbjtbbp2RhYugehY+fS2X8UOOJ0+LH
DDFv5usT9gN5/zHoQsxb6X399bLLdzPftLRocGjMXYT4uqhNdJMHmYJtza1zX21+
8wrbOeRmKCoNQp2ZcxbUt8X94ZqYACmDll7TIXm2LC8rHmH4pj3xMOVRdlchoo1j
rr9tQnCFtT+xcVYq7vEicYh7hGa1hIiGP4U2KCyH0VC/grzVha0b2fqlanD3eL2r
pHCovILDEffpmUHt5oOIR86FBBQoEUI+N4ZnlZSFwfVogEC6l/lPR+opmttIGn1M
H1Ny9zaGcrGVOTtdsDFCemE1ZBIPIM6EQHGgL2OXOEVAKE8MiftXun00BqO1r0S0
0MOP0Eo0NEb/eapTQV8MrXkE0CNlG0Vuhf4/9BnwqIaJ9ZP+8rofbGm5OELweq6N
LWDLvV4J8CDQ4CgQkCNQJie+LdcY/Ti2fvRmJv1ttAZSa7G3eBO11Nc7UEltKf/D
6QO9qe2pKQCtPYp9AJqsmnmpk5folQGPx4RC/0dxfBJUDLyfDPXs55UX8nEjGIH4
Bxd6LApCEpCjyq40a+McOS/2tDS0NSXzcrFaOYIPRWB+NHxjPRURUYcl1TUshC2Y
mVLT3jzwliScEikfMXTksbO4ZfjATu4s3HWacF+B9UPhdRasbUv2+0u0PDIQEVSg
WeEHQtB3bz1UBWCU7hTHDtoRkl1ijEFuOXU+C9OyHu0V9Xb3CIeKdP0Q+w6ibsyv
vH6NOfidAotiiK8E0ESmFzbNYFmYpXwgOlETKfMjZemFuhxNbjJjqCRGDpdJtVhZ
V15xFtqG4EbyZuDZaoR4t++qs5Y96jb7Q0Hr9zm7fvu5LLqTCJDyOXVaPDoYQK6q
M1hHHyr3iLLIbVmG6iSis+2Q8bpOarHrPc1SPGpsmJQlbhOvi6aQma6yCtNW6/b3
5m0Dd7o1Jkxw0GD2bMOiMUEmMeloFIhVhGvnUMCXlorZwN09cTYA3+slK6qXxbjg
Uk/de9d8E31pZoGUsJgGcuc0dCHdQ5CuS4atWx7jTltn6k1scbyIJLPFHAtO0Ci1
6Sj2kM5rPtTs4PMAOqBqKM4MaV1iQUkOdaeM9SMRLzifM2znRELurJo+TpA7tUsD
8iY/XzXQZ45AywAP50WE/whhT/iZaIKKQvzVwFU7/ajialRBKOi5O15m44DKttW8
CH0OG8V+qQax8ZSQY2Gbk8ekcT1hr+fx1zmWmrOUcbin8oD3qH7bG2gxuvoqfgrn
xEsHMcqh4t5ZlwDvC+SNkk52C7z+K6FXAOdxYThEeUJZZLV3YfaAQ19ozNIEP8rI
PhMnyBxw/HEpACygZ7W5Io9j7fwdk3/LGJoykbJUiQG/kgpo5QHS9UXKl5xLa4mU
dfNp0COmvT+54mqDIqWr+fO0PPJ9CAT7qr/LR1BWvVNKPLP7tHhs2wE8CcNYdo1f
ncSmvdrqrzLj/HUyrYDQlNxIq5Suo51YsPR1qlZmvuqniLXHhcm8cKmzLHCm8IM1
3uu69IdYwEtslGDC/W7/ML5JpdIh/ytIeVdxbhJJFN34YdKyhmIC+c1QIAH25q8t
R8P6rRq8lfcUqomlly9ons/x6eBGNjz5pUEfwrk1y41wd9GH5GgDuvzJRPZcE8jJ
mmfpM3FBvZKMv/GLOvQ5RPz7BJwFbmjmSb5MPRbIV4MiRZ4f5fIrBDIay7NmogDU
XO3qKjdaz8+eecnWHci7/Su7/UbD9BnFW7JTZqS2Q4tjiQnlKQ2kSi1eJBFfSH/L
1U1NGEAAe5V7Jj2rtRJ0W0K8T1MSDg+PQTEbcB9utChKD9pvZbPFG94eR6k8UDE3
fuLO1pmlUFJGR3TMwLU08XR8QKmw0sBug58RBGc/EeIpTrMoVeikqaiXb73gN/bC
x1qShFIXuDyY53hMd0qxwh0zhztzp414jD4kT9M0s3ejlxarPXGwd4dkAuz/OVxF
5BksnWDHlu9Hg2Xo3WYBHXPd541a2vBlKmeAFrv0Yr7nGKf23hE7nJ4t0cnaTtQz
Ksqd8CyhvFtump1Tmxd8mNXKYdEvaTUFNl4V6+QPAGaA4PVimo7yNE/glv0P/5Gl
6FYweQoUFJI3+c76mQJNLnN0wIfpbw8ytVSlIWXQ/VjHNCUbNCVEP5GxFjWOXnWG
gw9wRAMJ9JNvdynywc3HxYk7fRFf6nGX7wfPEGwv8+RmhjnkZxCCKE2caczV2nr8
j8SUogwpmUPwYw7W8+OHgbaTrU9KUBqnppaFtlULaDFiiKEsU3NXCFfg3XgosVer
qwPOIEsUwgprkmWhMUIXbWuordgLHxqePfJlUxMHq1BC5xWx+iQlSDo9RPThbVI9
svV+BZ8H1pfItokHBtq7yBpYBn+gN84GgE68YYaxgHKh0eLZ2OlDkWbo/6gyov7A
YnS8ycWgWo6lFs7Lm1dusw9fLS6sFTgjae+Jqh1UC7O5AEcLPUilh+u0+WCpK50B
H7rrKW3pjBbQbo59DMoPUq89YxsFDv37PvDs4PJhF4+Qwg0wHGnt2BfXIBki+OGD
zzgGq83/VcHWmP/8t9rtsY3dLzFZJFInqZF8l/dooWZbdnez62SdATSF7oXov/Ak
VJAoIgFlJ1jbdWmdEPFRmo5kNmPSGcJIVnyV/iJDUN+/119D5eIRoTVTa9qZISN5
Xx4Buaa+Rd8Nd08s7vgquXBvcD8KGZsGBU2+xmFswggdB6sYelvsjJsAckXkaW26
omOeTLGHCB3+5bF3Spz2PV+nUX5EklUubGWLF796LD/STsgq7vjy4odA6qrS8Axw
jgyAtnbeGH8uMh2c4nz3zJY0mL4aNwnOgkXQg0xF0wfd8v3oSDr1td0R6yz29Y4S
viAnTPOhiVKnPlZzGrW50D6nzu8rCrNZmXz2QOuo5QvvEr3Rfd9hML4Ka98JNmU6
8oap52p9wo/oIO7lGojiC9CQfVOYRocdx5AiVOLKG+yJnEKSP/BrDI5RGrTnttMP
x1RBKJynVaIVwAMhFmda2IZv0G/lieI2RuAs6FblkViODOMrbZWxH66pBOshFfDW
Sl0ERXavttMHO0TnejCzC2P8zm24NI3tjQKg1B5f7dDa672YPEoFY3FovLo1Ag+R
Hs85SX0GRH6G9hohs98CZLxpixloXhcMxCf5swP45U6nTqbeVkuRfgbEP/f8K8v8
qjos8R668kksjObdwIE309pPrGQ5/SjuHRpZb1brVJYmotUjC67M9jgLIzj4woRa
dFgM+swhfaJNyeIR6kEvOhIYdLScKmRPePwOaWoDX3gax1XaceaFwNTmTI5y0YJX
WYurLfaYuIIsKu6zsdqemfMMqWTYty+9omeVhmZjEfE0eyk6HsEUJ5RCOZUk3pLo
W8U7csif/HxUcgtmisHIepDGQoGUOfpVOVOg0e1IedXjlspAm/W8k0mxGhrTUCFd
05QwyVoJ15wcuG0xP1ThbPvMgPkts68mkHfBHLmMWE29aW9ecW9CKqtGPc2yrbUA
xYaBdgk0Pxww5FFKMQizCnfhnWHbxZd6ru2NZ10FhcogSnq6wBPIirNrAyOsCyI8
XRVaqa+isjo8tidR0H9fzQEIVm9hpykx9nPqAnhIh/1umS+752YJjPvt8zBPsVSn
rJALXs3COla1SKumMPshvsxXzIkBPZv5VNmzm8r2h3jnYMaMG/3RNDAAIqTNJsh9
WL3WMK1cQDiyDURhcyZpIy8j41oU1kGIMw2E3llm5n4vvsioiJZRu8Y9Lhfn5nG1
Ar+CuV6eik8NUdeAaubvL+zMvmK7q07PpljHbNtSrjHuTxwhNwtfoHMzHtE66E4z
lILIUOWxKBSx56rmvavJDfo7vH7uKtGWNq63NZkAYw94JDm78TAFCcLO3IDu+q3O
uAL3FSwOf7GblwKL71PneOSo3peRWw+yrwc7m4Nuo0vIst+q02UMZdYJqiVhROLW
XQNMcXEyrDiZ/+0WgVF7PR2TPvN1VZa5/D1tss5MjEJ3HTamQITkFU9MW/v+L9yb
lClMPCRYFGikn8hYMpknCg8P8dS/s9E9QUuU/hErwPhroyyD7icRkqec/grawM1R
MdAnNbCmgRrISWatAlqe8Gi/ivSPEB0k0RwaO9y8affOXCpcdIOLoY6fCiPfpZ+w
IvOt7I6L00xDuyGeI6qrQOjSv5wKdplhZBmdaVyufmsrDFE0PSd6Pv0d4o6CRhyf
s7VLjM73AcxAYtcLY3BjST/5PuH3QIXFr0Gm5PLWzl5cx/6wfqJKhEipKoZkHNsX
n2xrISBrBbtqDtaWsliSU2+iZl777mT/9Oc+bGGyjS1jCUhEVkCUpFgx6Zr/S8Jg
U8u/WDk8xpo21ZlmeDW2ZXxW2ukZuHbwmt7PhowSzCAJ5CuS9VjcFdt6qnCw+tKr
qnLBUrW+59qlai9w8Cpp5uY+129UPQBCwb04DLvIdIThMDekUw2p2o0eUks8n2q7
oddj3k4bJETgw9djYD3vch5Zv2gJcJdJ5XO6VghhRRn8o+IV2mpO2qaztem2qIqU
X0/MEl7n6BaQGZv9BRGr6B3smn1fd71x0PsFF2C5SGxbFFWFRoYbysx7qatMMsO6
SLNBID2oRsmGdBmzEp14CcxUCKdzc9oE/AkfH/s7/enUSy1jUkapJMM49/fdrFBJ
ZQ0choktx5nGhHVO9oZF+5j+rgoIIXflxJ+DO4y6ZF4luG9VGTVohkykoUWgAfwZ
zrCh/e1LG2Gu4hyeoliTXKUnehkHcA8PMdeojRdMQRH3hvFLFGyuf9fmXQG+PvSE
DBo+uxGtWPtfp04RdnYGTLupI2DCrLQ8NjzQ16u/BuESTomyTkKmuQ633O8L0DTD
USM2nF5phMELi3abd1eM52y7e1MBtKTzcqJDDfy8dGdse1fGbtjx24pAAzNl43Ip
R3i01c0wY+OmBOrJAgyJtZO/IlzAXq6GxEOVwiTmhbxaumAkzFHjj7yCbydpCp8E
mIjoonYRycWlDl4ohC1FPxsi+RkWrlFzHDlFiCXZSByUQRTRMAEbQQik0LB5YeLn
uzePdv3/G67udlUUAZAI/LGlAgYt7v1YvPPFuRL9nMQJ2P9tP9WsxsB0ve+21DD/
SfHs/UbTI7XCv71Vx7X6fd0BHE8FyQHNFCLX4Gqm55NjDFtw4lNAhXBV+E8Ef8xr
DFFSbV11XHpAcaxChRowdjcIdGCkuHf5WQiyDlH9kw3zupnt2ZtoNYdAmK6aXCCL
kGTp5hZobYGnieoqSQy0XW8mvrBRmXya2MAgAIIQ2Y92WblSCJCpJIU9r+mkst1g
0xzr+8y3epOAcQLNKfHnEO0Ih9AOw99fOrUo843UVdhFo5IvGNKDpXBJtvflBviF
7oe7ZbUu+tP8CNxpI9Yi9VpyYI8bpw+vLGPGHxQTDzjE15UaU0n08e6U19hN4xm8
ESAFx8nvvaiMIrOCWGA+am3pqlMMs+LBgCoxgvVOwMRtwBMoGpSZBiEgmlYOTu1v
RB1CRHOZaEjXueiARsFXj6RJ4xUM6X8KM2zCZRtkcNimJPuAXKcKaBDbZ4FLR6L9
MOwdLVwkQa0Mui3ubajATpUktOKk1WxTWhj8inpzQX3aJJ361BRtOWzokGDudqMH
K6BylrvFKSW2vDA37qDR4wSubseX5UZmPDMRwkyn2REco4Sb1vtC2roxACyAIn3L
UjzKVPF8VsnNNl1Z45ciUBpyvkLUuOWQ20h/7JtI5nCwDWSWIi2CKvploykB7hIw
69wGeD+sY/eG2mbYvkpfEjs7kpuKnITP7dN5vOS7+CgUCN8I0dI/TI96EZHT4bh/
sGAzjcrnzax8dZgza6npyHzgZFryj5K+FdvN/J3pwkOTRG6dqs0tVRvcPrqtl4GB
hGK9iRmtEOD24gOwZbVHmK03vNUtmSnfolOAS8MahK75Ox8oBv+HHSRMU93VBcBi
C9R1J9MftUdF4feNvq7kMJ6yKll9Jf/Ie5Ifn/GCQnKBPTI7lTRgfFB1w5heqcTW
rDcQfwmU5jgo8nzPm11md/duxV8HwhOLU14PESR5m5JyZQUe8dqZ0AVC19NiZfS7
Zsznj7kC18QY1UBi8j/r2ExfNAS9qyhPuFVkc51eGqfrJo4et8v/sfHlHu0l5CUq
2bbudYJDinHZ6iGNypc4CcMP9Cf3wW6hgkl1ENpQ0u5L9tEid37nhGZ2jou+OhR3
7FmChqIZ35olCM5gY3hYvqjJ/VleefyGIEk1dIJ9IlcV9Mx3CV2kVX+6Fr9M16XM
fnQBD/8uHTni3aLLe4GD9LRZ9Pl+wlPVblbpV0sGBKWnAxOsXgF+2xCVfTGKX/Bv
/Fuzwp1tEszcg8v11MjHT6h5k5RAxcDidGcY4Ts5/6EOKfKSn/EQ3bgqUlWaVNCB
gw/PFQjyZYjANlHq4CwjJjmszDMe6BGRoKgZzHoFLbJSoO/GtU3szbTCAHZUkJMB
kSwpBNt36Z7VWXPPi/cNzsqIinYgI9wiOI80AbkwTnARWrSvBSMO4t82Nv7MJhBH
COT7iKi4gsv8j9IGk2t2+lX2EJopv8i2S9n/giAhMRriszqqg1eHWE0PLL+tPT5V
c6xMmHH3hPm0BCh3Av012n0lRZL1qdIHTNEgEM7y3sDQLwKLvMCdNHC4LoZQSlws
l2u62aLFC6ejsgZwWmh8u57jr+/uPHILiWVwWvq2pOoFa2bkU0LbiQSmeVCd8JPF
ZoBtWImtvvabUSUytzbl6hzV0679JAPU3yDID0NnMnmYyQn0dZwQmlqyhHNGc+m4
RVQVhLwkI5WSstAW/12ex2fAlRAEX2YEoeL6zZYJzo+betNvRSADhb3C1ZR8T81X
YYQKY0TVDKmVPFUnrsDi/Xh88YDFK7F7uYFRt0EcHcE0DputE94ffFvf7vIKayam
XpmPUmF6XCjPQ/lXON8gmpvvp+8M1bTfsNFT6YDpfEDK2jF34n1ybUgVkvlmqcVt
OlKenpeOUWXwbdLEhEajksNXmQZI31TUN+YCaREZSTe7sI8PMHM2SeDggHeRV0tn
hEGYH6FBBsPpKoecevR7ysbqTpbxcHhVVLmWKQhLgbrDSx75Fg7hSRh1rT+FfwVk
wv97Mg5HLJ4U+gt05IUijWerqEAuc220+flP6c7Mn3WcS2dQ/srhC/amwb++4eoG
DxI2Ki2fgn74IQTm/M033K4ExD1MRmNUi4JyuxoGvnNzXLJHgs58X56K8AVOZrg4
Uy8txm7OELgSGvgO4AnO1CTRYgS37mjOlxMWk95ntv4UT4QHsm58GPBBAOsMIMjW
y6tI4U/OgeOt3TACQyg+RARtXBI0cvx8L+gFY2IARRGZclKcyo4eMxciNu+W+aA6
hNeVG6nA/WUnKKlwJx1KnXCPRtxUtu9IQYP+Je0tv1Q8NXINi1rbv2d/uxcw7jfQ
AInvjThO+Bud8CflvBsFig7mXfxHwJVmoyWjvM0NcMSR0JIl+dFzZb7V+u90W7yC
cyz9zXtlR2M41JAIBP4h5NOjdJzWSpF3KZHRZM0eIZF/OBwvCW4WJSPyJt5zsRKp
A9qeqHoHS7nKbb/JG2K0rrF+AbIta31orDpovyyCcmA7de/7hI8gH8ny47Tu7WRH
1e55L5/A9UJQc+15SxvL3jEkN6phmJGGs9+x2mrIhR1vJnBSMMCsttVlQFxpm0y4
kiQjlk0pxMHZussusIHqdZDD82Ct/wJOxd5WuZfXQAiUD7z+U4S3VDrdmn99LBPw
pdECvc4eIrhaG+BjIRRkXAGAd81WHsj2nAKkBoOC2F5ReovvQ3WWoOM2q8qV7eXf
hR1a1BofnmJTzSGuQkQWQHOtKpt1FEsniTEZexwWiYnxMGPdRFEksObiJKhfgCf2
JrOU3kiAStEZ4t5EKx2t7b3q9Vb6VTrnR51CGQo6INIt1HA+5+BMuvhr9k+LPFOI
0ihhIMupZW48f8Tr9HBL51BjTn61oIYx7EuvwK//fs3gg9jKp8343f6+xrm3ls0m
efi4hvXaMPqwRUDv2eLf5OihCK7KXkV2666vRrJa1TRPiM4mE0XFfm6AVK6luX0d
wEsOjzfozFoXGDh8THTsd3UC5HtVx6BYKmbRkj9HyP1qq6xBI1Ieiah1CBh7t/wq
Is9uzuqd1XFBfmHCdoAvuWiqI7FUCnhPvga8AszPhbm+r1+svMe8b9dVQPX0M8SB
j/eE+NPOv57IIVr2zaFDT2W8MyCIvm1AQ6MYPYllAveHVf1rVtsAbwRNoOe7WAAp
5m4hNE75CfSwfrB09Tn6OaFfDgwYj95QHW8Rajbhn+GSg7WQi3DtwkLnsSFBNJf3
Y5qW9tytdmMJ4m0kjhUH0tuYvQl8B9fs5NRcO4dFSDToAMoEL0pCb5zEOuJow7Q8
T/3utczJ37cM/jJZHO2q6kgtm4J3/gtMq3JD0YC1pK7e/px03iD0ESS8Io9pBkZe
dkt2HUXZIDGjAfmkuEjZevGtCBGpHutIi3V908sokcxJIoCHU161QR2FPVGS9eLp
BWjrhokkDUyVKZ2euVHgDBQHUzGv2DHcPe7qDHUS235qPflrGsYwgRDsWiir71OR
F2jNdZHH6Gfdn9KXwY0ICSqB2cCLEYcBWpoktinKVkoc+G/fUkeDFXsPSiyIVZzx
v8Gc7Qj/8dhkUakUI1YFgD0y6mwova9aTyEnsH4go/AGwVWZ2bA8sgSRv3rMds0B
s370pHlrkHH6LkySsJXnIvJUUjDE28ItrzT9Oulup7b5JKqI5sjgE8L1MvIJt+/C
8r1ig5lICS/2eHp/YI4562dxPbfsOaZH4QkQQbol05B2xNGg3AIuYSD2b4xYEVa3
9qeM23r+gMDDtGkTQGXrp7tECmSvzehK/4Dp1Fx5wRtfHJYGv5/4XszqIMHtcqZM
SZFhgX33PGocoAFldzKhiV4qp4ofboO+RfcfHfZBMbUre5n+oaK4Hb+TF7lGJd7j
ZNohVhla+aHLOlJYe6njALakFqJpp2l9WWjb15oo/hCAX5HYU/4GPUcgI/NX8Wes
tu+cWKxWS8Rp3kJ10zqk1KWFm4yTOqErlpOZONggZGCurwgrNos7rcm0y15vOmBZ
CmgFUwSh2Ea9hVdPElHVNqgIYkC2AlO+J+s+VGDdlIXDRhJurRloG8SzBo/P7c/l
6bdqgtf0mrhAQNTn3yF7VUYQWqZR2VruRoWhnvCglLh+5b5mDvYsWVe1ettSr6Ab
oniEFmXniw4O7iou+/gmKYcsr+17eEMDCPX3rWa1vpO2E5SjZbRmvrbe425nkhUm
0DmMY1nxet295OelC5/czPqiiUkw8UpqWxADIKfWqFxTWO1isvvOd/iRZdFHPjGX
iMXmGQPJBGruv8zleTHxZx9hlLpmH8fGIWjwVH/TrVxpDEHUFL5uBsJR74PK1u5E
Z4yT35bArAQhdg2xgXUGdkJaP5TH0blzo6LLe1z1Cv8Oit9MxzsrNFK8f9Oiy3Uh
meOF3EMtc3pTa2lDl9+14G5KGyRyKVV5vbUO0dALksKsGcloM5cm+b9xmIKP8J7J
GMuRn3j6vWi2QPXH29LzaE+oWT/1OAYyfBoQVx82tMu8vVYMzcQRb6o56DDlzD94
k6lXArPigLj+gUE2KAvTs63C00hJlBkJByt8FU0HEJESMhFvrYUWJeSDbS309jw0
iiDAp6aeTqkqJtYha+f6TlG4D6OLDyJolyfDeiYxmZ5XkLmueKqG/EKP2GxFn082
W+Uc927J/yXskvPCzg783zRWwJnB0m5EYkJbtkTedjJYLmVJiq4fPL4T+aQNjhGh
JZ6xzyElJYcykmnHwP6Tsm1oXhjiY2FoksbpvTg+ZCZ/l7Xc+RlRhD6cbWMTEjcN
sNZjR7z+IJzxtXC/WNHuc+r9bXcfmhACAR8C2pU4ukmwOABNtuBJ8CBdKS5GlFev
7M7zlJdK7wCowTXtDZaotgkN6pJKPEBfAV5CZSeSwtGknjZGyjapdc0Z+wGGyJX8
aWq1Nsj8GhAToSk+43ba4C2JMb7D+e4bKt+DVfTK3U0zOtZaOIWgXUlvQUWRdu24
gm6Mz6XGIc0hlepsCmHB+lVxieAsThwTZZ0WWTom7AoCqNspimyHibA/EMhj/hg2
8h4gmbRGqe+qgPRbPGdFA3C25vU+rKQTVVSamOxNPZqzQW6MwsJdWXs9wKKqrWJ9
TBoJaWENpvzyKsT1JjpXyi0zQgFz454wizcU+95E18FdPhHSy8x2Dk/OHCNYiivi
s85i2bTHZK/vJ54tp6mXCILhECQH5hlSbb8836ZWWs7Zh+HKWkQRvn/49Hy/1xPj
T/0Put6d22EO2L4QT86p2tKp3OhKiQ9slomLL3PYTa7Vj03289VOiaW+iqxXOk70
HVPXj+Eoq+mZaEAhbYnlztFVTjyF+nVSqhX8TSDYLOz93+XSDza+Rg5OU9dxZPSZ
Bto4CKKR8yMk9JrwIl6HTQslrHpD3pw4YKsaV20xivmPXVHysHuT8azK+4iEIBpG
6UMjb0ly9oa8rLIoSH6OSHB1tQcK/TC61BAOyIRQ8GzIInPhzJtfSKScoWTBuknH
YAOF6ym2/bdZA/hw3X0ODPrvZQTjnSCCtv7osLpIVZw9b9RhgXnmN5meXsPr3Udj
1aOD3/tX9vz1No2QmdEfibwlp19fWQ73JnTVva1p7k8W1NgJS2LOgW0WhXl45E4a
wOkQlvbXn6xh4MPFxXkqdHYdGSBOUaXjqSq0MnimMdIIcK7tx4BwiauGmOFA7WmL
qC38m+DW/pL329WGZo1NNHYl3UrCefaGAsNiZhyt2+jBPkjTTwA7hxyzHTAl42/O
7nLb8CYlFZMSXMEBdgm2hkDSyyDotdgXMjyIrkQbOW29rnyCuhEkqrJz1y+wyVIq
JumvSJl4ZHZ7AnCBMUNsJNKXCLwsZNynx4WwQ0DqQxNEsObLoIykLa++5J5br6l1
vKlhMgKRb71u3tvgn5mrB40wfCaSGEhpQbe96boRaXPXkOwfHcg60Mg58AKDugty
80ywtpNEZB5Sm6PWXcWi8BfoazXWp5ExtN6oBSY0efAoHi2VJzozJ/MbD+sjbUsN
9IqE5dLiYnUGmOxXpJz3Z/3HdSGD5SQAu6Z6YrPPEt8xAFOFKkQq5qJpCDdKUe77
G4kvbIIPV7VVdZ6XVxTru8SwimlKCNeHplR0wSV5sQEiCNB5+5mvvQ0Za++gupfc
7eFNSaKw/xdrXJWNWGw1KfQEZ5NrvxyyA6AN/0DeP0jUufz2+M4Bp/e77LQqPbgK
rc6ojhi2+WR49ofK27rRwhRx16YvoCAM1Id4dZIQCam5cfEtGG1uiJp18GirClZX
3QVWQ9zp4apMtlaG3UuzbSxbg2L7GSy7wcYO/QCEzq8IQOZoVBEQRfuSz/cUaT3U
o/s8SH+W85pWhWrk3eHkNszXSAbaUxkOQr1Enf6k8MEHpjsFGki+R7xH5uhafy9D
JiijD58mI3X6mifD+nJgQ6XXLVbK/Iv1oZ70/59pvIw47P/Vw1bpWJMbB6dMHQri
Bsi6JIrhlCqOs9N+l3Ea8KEWWn882gXaA6zGOfkGKBZrroElkp9p8VYPt1S6IVUs
v2ozB0IreBp4EfM1lnUTcMKC2aJXqxVxXkjzW++lU3Yy0lgYfGXu6RU4W1VefQtZ
fWRiecNuw45QU9mITgnqVJpjePJ/255S63a3hn80n3m9fOWqMTGrmsjU9URs+ARY
qonS436peFQI86NRd3uR6J6GVOr4HCcxrNr+/VOGfjQJ20vwTmg8nHVhUK0AltMO
EVUCeGI/InCJvl47EbkB12VQsx5sDcj8TKGMIwzrEU9QGuUwBX6JsDsRER4pRLja
WnENuqpFqCvRaZ/JdkwYexwj9t3Qx1Zckj4sfHLVE9fG+J69DjBlTv3pXHpxNb3i
tmfN79IaGF2blDs5FzrR9ZJnOLmqCp2IJcQMQh5au1xljxttSrBIn7Y+LaijX344
MlXP3jgHle6dq6QWJywU5BkD3IEalyRQh+rKiH0IkiCcYiLUrhApQlC0js7yiu70
rrn6Elhh+fSYBaRk6ZIaSDhb//F1hHBDPCNNJD0SeRXtfBd7wKeDfR7vtr7F1Zxz
x3l+/BMviA73A4oHZyU/fom2yBHc1zf/t9kd+FoB2SzLMIKc0qdd8pZOKzy6sCSl
IZ4+GvwWRGl7Vw8laUiYYxo98EKN+UVGIeQtGPgFgIGyp/3AQv1TkwLZshIQUrKc
GrhbvXP7sv23xM2dKV907rxwKG5UKaM4h6jObnB6Qlfy6rdNL/CZXM/Kzjo2QAjU
Cr4xAedDW8xw5CRreeeOvqi7ZMxZuULJMm9bNfUjX3juFA8H5jyTX7vc6aTlpTjB
pauL2uoSG054HPdVm+uV8dIUDkb0gphV2KgeFneGUA98HbMub4RTZOba1sjGE48v
Lc0LVYqeKJ5Gvz3JDmlRGf3VsA0saL0ofCwxnnT5TqqGpcRTXbLSYim9xPPH+LJS
VO+eYqHVXoVcSKcYrC8FH91vN9G6j5NCvoqyt1R2SvAMej8znpr4jPfvZnVUxS9j
/OLL7Aq1vJ4fy2cI0M6IoTGMu8+qr4RX0bEwa3cgty1HqowcRmBE6LtVPStJo+kQ
hm0YaXS2HZnhUHCBbpddStUAR4/IOLaWwpKHKAAWxntGMwaddNmyotafzdabKmeQ
yEMGaequXvfkEoOdnEvxi6crfEsKxi+EPZ5TkxVyoW5SmXK5DxNqeTxJsieFHTJJ
Bfewo3/bWtCXvkQUh9q8oPZ373YLsgLfLBVvbsrY02qW3zkzsP4DKjiStMt4X/ei
FyMJkFXFy3zk6J8WJodIIP8srNYhG07n7VtFt0BAAFlN9vHmhGg+/VqSDwZD9T8D
ZCq47mHfkRisYuRpymQRVc7Plsb/YdIRC6VrJSaNWrsqvYTs56KAYkH7i9MECXBa
VPyF1C/1bGenswudXN4U17ABYjpUjwmRhK9obOr2lvYeHTddsjoFS2fhmHFucYhu
tab09lKzZALFPYPzwK9iBq08Y/uUuQYRIDAQlqjphuTs5QVKtu1pXP0k2EGNFUdl
c2Mly/MCZlAumxKlgOnlCOB/DXY+zqOTXJg4Q2hw+mV5sv415CFYbI4Tw9+6pt3G
QFqAx/1SWy53UQLM72vIggQcotA+bFOyi3srVV+ttNB9qrPG+pyrKFJCbaalkt+d
sl92c2NFLNQaEFHfvg93zNZ4wqToPJVpdYebvv+eGvNSX3m4oll/vrSybZxXSeok
VucdqFdwKU3J6uD3NmpcrYQkK5oSB5g6eULFffbsOo9rXzjmB4WwTHBt3Nbv0C0g
awZ0MACwB51Y5rCmvPm8QPsteSKNJ2/xWuQW2We+o0YHg04Z31dQI7Fjr8IqrWaj
oz+EEU/tcOTnMHv+dpJqWNOvnDg+gv6nfBPxYCoSimg0RmGQv1n5cTyj2Wah8qT4
Udtb92/AYMXIvUG1WCcs3VZ6CCfc+FTmbbB1wvdD8hBI7nfrQNaBsaC+RYwR++m2
qlMhM7FqGJtBBxDDhoaBauyZCg6mIELavTwn5+U/Bo2Jsn4BQFnZHOKyHAU43LSJ
o3xRcGMXgVoxHzbw2ckoItwNdOMMHdC+qP0aIQedTLaACfJFjh8v/xH4p3U+rM0U
yonSECCxHRQL64JLcTVpzcEuZv06KikAOQApuTxin6+YlshnVvLkLcrMTYDRiYd5
Cp6zIWaeD5rJf7aXgpcoAMHYESp17cuC7PYpLZfUF+bQzklTrdX9jobslcvFtLtW
C7ftilvvDeAsOOd78eOyaqi5ld/dCC/bi2b8Kd81KTX5aF7VSsILntX5JwPbnvAa
YHBi8nhVA022o51PREbehAUuAEl1eGnORW8nwVPNPcaCxi5EduOEUUKg2FrOF5Cr
6F6Tt6PGreAxEuURGd30mcL9mbc+hiJY3X5Jw4VKQLisxFBzkY5DSMGIWpSuBx1p
fgt+PsCN8HrbJAsMbMWdjZMeabWPl6zgROSGHOKqidpohnGTzgsJEs7uv2FkzLEY
1vcxoFKA0ayWAdaaOTKE1F+fyr+76U9mio9hIuLfGFsk5q+RudsNc51b5NrFPftc
QpJmeG5x7iUHSER+72kZRPVZ6F0xXd7BDSzghAu1oM4sqoixnTDfSp3atBudA17Q
OD7gHfW6uit7SI1CRk6RHG54LPFaScT3GN7XqX77bDpeCpZVZkPCj6pT9S9kupAk
fKhQeBpmf6f7gBXN+Pa4l4qUCrqlYgTzRAYG35san76ybst2WEN2VSN8aXSTeB5k
24OdXTYG/PH7viBlrwGQEi+zsMjJa6olx+rh/8swEQabPwEU1lyQl0+TWSTauQ1m
/16MDe5q3RY/tt8bzt9nBkzCqrwNfsvIkAQKu0soqZ9vrKkP1wMsx2MdIa1hi9Dg
iVIRozLQdOZFzH/050p0lp1IuVj+8Goj8v+PQGf3m+NXLtqB9FtMlDGLLB9C+pOF
C0hIDyFYa+aWl21yshjQdiQJsR3v7EoXfqGkUrHY1YEIL03opw3+PiGKOMjpe4qH
3qRMau2ngixMfAwBGsAdN1ORAPOzgWKHJP6FZs9ADtVx4AFhi8kaoha/Xz0itNVD
K9/bNK/IOEKjVlTEp96fMjC3iF5199qYWWWEynXLZeFDTtkhEg4aS3jvYluqOH18
PRz07a9e+10NpMSGCnsTVy1ITZ3H0sVBCKClu+VZf6fcTwH4oLtiCKzL19H0e9Vs
/X6zctkJzCF4SqLyZizZ3CQ+gvBvKaJhbxArHaA8nH7b3h/NClRJYx1FOov5DitP
fEI6E8eeCuuHu2PlthDdOxl+ivQNtRPuD6yCjpDRs9MeXtsPXrBtEd4Q9cts6pqL
6cE3RKMSSooAva367qkyqn9IeD5D/lcdxuYhmsd1KGQi0khfXGZx71vz4QNeAZOV
touTGvNBpSYhg7ZxdjgVy7fnZcNDISPpW5uzxJ3ujfwZxxfFY0i0YkuCw6kg98W/
qODPFvCwvj/UyQ83zLkkvdawOAzhA9bwus54ZJ6d4NlJo5vAI47tOQHru/vBgF5f
wLRRcIgcQ7U82Ncx5ETDbYvx5V7LjSO2Y6qRmNtu7uMwvSA4wmHs2fYty8EZtQa/
2sEIslotavMrnX9B4iMML+HCsYjH47L2fwB4KFShYCdvUWuSRx+wEMO9wLhqEGWp
hWVCXvrgfckrAg5AMlioqACdui3AlOqIoPYOd2p+S6wNVY6qxGQZcu8YLToUaoK7
eKIfHAYXlzE26bw0wwCGDt8/YLGF/G7Eib2kgPcMv8ofTbXDGAH1+VVQaCg4kX5F
WLrul4f6sk1EihtZCaTgcX/Hwiz9Wm/uzChQpUe3Av0FusCuLl16Cks6MrF18gv/
5jabkMS+sfnMHXQHx5LxiwwJGPRo6kqXFbDuXX1lD+brB2VP4OPsMXQyTTWYxVZX
0/d2dQ+cW8caxB8NEQgyPneIbs4FnF0L/ZDkfes5+UbaelBH25tCUI4e0kTjzTxw
bMz37n6BW6O+sYlyWgTmzThOgvOMnf6GLkmJm6bi+bC+SVvsxsMTmYsSrsVQI5CP
Uqzgx9LcDtnC3D8fjj1PsuFEufW2OjwWhrsA+ptAtEtnrb5FMqOBTuGDHk8ogUtR
rdY/ztXo6hwzfqibkJAgsZQEUNLOyx7htrw8rsVHM0+G/wK7iJdbB+jFRppFLhJV
D+QNReLQMw30qistPZ740mGA3rFo/dA7sW8ACQ0CfS9hwQBSR7yfrkpeZHM2hvu/
BhcHdygpjykW23wUl0FMiV73irBqu9Qct8Owah/BCSc3355mxJcgUrwpezYJHpqr
Pyu6lJQ4EG1Af32SYeyNsdlwBK9WuRXY4JcnvpKMPb9rKAnlHjplmA+xYy3JgvMk
XypiXP3jT3scFSKj97z53F5ZEif47ffvLLpSlhkbFxsW6oFzDwS4nlC4d8h3/fzi
ah8owBz6hzY/N1mtbtYosLNlVcYRlxXLjQTDlgAu7uFmN182cK3f0u3K3CHIBFuR
hRX3pnntLAL4LHpFKlrq1W4waQFnYAtAq+fDpj5Hwxfg/mhMWcCcg1DDehyWKcyc
3tQHyKwaivFqSh4R4OH+AT087bmp0V9NJLm1A9cWna1UUUQjb80+8HPUYCb2FnKE
qgPow95XQrIF4fVEBU8JqeJz0lb+YDEZdLZipSDaldVvZENtmun7fO1qz6Ysh6qf
+8XqKj4v5l8AJLCORdcdXD4/avbq6H408QwqwArXCIcEKTWCOL5HSgw6jdUi/ncw
4eUHjDNt7S9nA5C7GhZbRQVjCHw0nrMqbNvsQ3zKLGIxUoMRmn9qhsGNW0UsVwE7
x/ELv5y2O/iT0ZBX+akIZbA0sH6padE7B1J/rzN93sXUhn/pTUZFaqq0wFrxTqVo
HKl8tkGADh23UNAnFbn8t8MBjCFIWK7E65nTnDKkuyiyhr5SA7Jpdjw61nKNOEtj
oIYaH7Un2+VP/xkLndrnaZavfale7hTtUmrOMKMbmxyR7u1zdNRDKXgbQ71pr6cM
f+2/LiDLph/8a6khk1Npe+GW4YpReBjMHuHntJ8I4eAAxb7UaPOhdovcQF4z4Wyj
GwSvuPDIyPSXjc95J45POhpFOhE5ZpYA8dYRJF0wazgvwbHGfOYZPxxrKEtw6E4M
w25RqKuFODdoWNRXBCB0qw/ZgJqgQ9SgtTbIrWwwqyDDWVsSp04ngGpZUeGOE/gf
AoPLDIMUPcQsKaLVR9L1R6muq47lmLti3/SGTtL8LJ3QcrGbUhXMjEuCx5OLSixe
iPXMTotzg25n1o6aRKtRWjVF5BXVlPrafi7/X/VgHY2kKbSrDyjFFRpcJ3uqo6rc
mEeWP+TlgxCg0ZL+ceD5ZtxHuYcx2boyq7YLwVWpgFtkZAR8iirL4JpMqoIScUjH
wftlL8RumHialrAEUczxJW/pk6QFaQpwJg3jjiObXB5B40bQrv/XSU1NM7NhJz4E
UTvUSYGguF15wgqTSXH0EkGwoD6uYuX90lJnZk1GgOnbJ4YrPNOB2e60TGLax5/V
hd0j1Aa6AO2UktcjzxcVPR3MbqAqXNLltjqxv2Jk7YKz6qASrJR27Q2LtcNfQ+04
+rEGuQ2ARLc6BSz4I17WxjYUnWUgbeKqsg7O8S5hCj5tae5z/l7UqKvZt+R0/O1k
RVQ8jPDnRL7V5vOGdb8n3BCP92tTLLal/hmyJ/xLHYI3Z0kH/nIweLFAl+VYzoze
Z4m5YPQh5BWxRT2oWakjPO/W0HNc7WE6KfHlwhTjGJ/Mc/u6yGWfhZm5mu/9q42S
eX8HnLyLRI4d+KFaxMHn/23sCLkTGhqgB1AzGkZiBYOMa/ChTQBw2u33ie6t/RLP
0GIilOxp09U5qqcMN5cE9zRoJaNTuhyG9Qc+kP/0wuN2gNqwWZWzroC6dSceqWAI
D5A0Jl44RAxefrLRTPXGy6sO2vI3ORh6BLuwS5r6JWtU8p4+1yGmBPha+vD0Yam1
X3/h4awAtKPkq/ir1/mau9ONVVFgGyAkaXGPZ9Pr/5N5uwbaC7s64tEdWK2DrJkx
wxNNpm/bcck3mhFtPfYf89ugHJvWTinaoClJdcIfKIMKhHo3m7FR6Nnm9plK7FDf
awiiPFA7YxAs97A1DDJngnL5lhRgzpEfpdrsO8/XWakUXgfIN63lsdIpJal6t58C
CUpph30FTMmwATh/HY7wT4O9Kmi4uxBn7wJ3FZvriSg4rpS1N23lLEKAVjV3gvPt
q1bLyyXBS5dLzoT0Y3c+wvD/YEpJXvWXoQLUij5VQ9dnnAKTuq33eqOuXC9ODmKE
C3KL1FFcdoI4VSIdXowxBueG30sR+soM7K5nqro+KVcfEEQaWigQgCsK7H4XPyPG
NGlZ7I8PMc1okJmRBht//Q7fohdmVwG+qLMqz8xQUtmKiFemK1UHtj068IrQNTZi
2Ub5PsM2zr74VCk73JGpuoqP/T+ZpGTU4VcZo2e+vkVsXfq6SKzfTjTCxd1OY4Yx
8lSuSLLwXpBmGfFHXwwDOhXss8Q0Cqz9YJ/BdvEhYlTmfkE6s/LmTw1cCPo+khvn
MLZbBTe7jPrU6b9g4m1qWpE0VVVMJ1UlcYUoV5/Ov45Bn8ug/m1e2hdXoAWJ3HfZ
yP58fqHz99WYskMmUPNbAcXkEQ9FXdwu8tcIP+56yeID+2JJb5QVPF0uYjBuHJge
0n4cQX5dVzupk+oNEk0KTkHK3nVqIc+nQhX0c1mzv/yYc3lBeBcu9qWiWEUdW7Mf
CCsBrEogQb8uGbLnN7EzisNuQgEZv2srfOLtsKNJhfAr4mKQtDDZ7xa2KnmHvTin
FuakGqkoHakdOQwgcZZdB1XQ4r0Uq/SBN5iW+ze8tLa1RZYHp7Wlutc5aESsj1Qa
QSZwmfZkXTkHjr09S3GaUJFnPZlK4suwtZpAKF3CGp0ZmOvQrJMbNdDFeDeZMjn3
fXKDGBIgMlahojxp6tpPAsqRtCuoQSFFNHjv6oVqqciketWNjOtovfuG/kLUC2qu
gE0TdKAXT3pywK+XSfB6rxQDEImBlpZonCIwleCsaiddrxuwYXAwxjh0LW1i51Z1
v78ayW7dlJ5VBktRnq5o6JEY2Yd9V7ZzfagjYhgzxtzXcSZHB3l65096X/GD/ou9
qoAPt7gHskwKxsFuRUV3B8UsBLPeyUTQt1JK7ygauYe8trkXKlwDRqTegNt1hVmo
cglHF3tEh6nZDqNZRUgseSWoCpzJwHBXmmnbaR2bRnPhR2XE+GW5n+dqNuz4x41F
i9/84G9/yJBBhE0rxxGneO/+UF3EvYffoANCL4QeRiAPwAExwY8r2jhY4txoq2cu
xcp7NJ7Xe7016/UeznVo1eHjs757/nb5Df+3OeDB6oLf5Xo/Ba6ix7Jyf+2jyNIi
zNcig4Dm1jYNb7Bt2BlP0v7jVmX5OHvttpcZ+0iNODbQ2qgR8/3dTKSzmrfmwmlE
Tf8hXmOkjGR/91KlM2B2z5sREq5+0nJBk7cB+wL/6ZvM6HCu9r5BDzrzXVis9Dgw
qp8c+3pbyeMfphrdSUVzEfhyCFidQs41o3/+bCi7Kt0wLMWBnGkBrizSdZBHQTIK
hyBZulzMMBVDK5GeePsYQVVrxMRFBPcpxymJmNFRnlV9xdLx0giPgVnQ52utEIyy
kKwFIdCX2hanbLXEqoOH7Z+oUeEP0vnm+/GFMyX4nb/FD82YA80nkFmfHNPVTKg9
voW5idkbGRY+Zwdk48uPP4ixTCr/24A8Ya/OAUsTx5qECrY1gZPLXHKtiuXzTkh9
V1B9tEIpNRuBujCHlluBaEZEY79exd35Apu/ss3pp9BqbXAtJj54qzVx/IyRVF43
XueJFxPxaFv4HAf8+myEUbBkPrhyS9cEnOpHCD8LI90RTiTW09qt52eOa1oXs8Ya
Vd3RuNSyYZLAKA887C5d6gO5T/1eDkkTYJT4xRb7PfDykuSB0oKWkxEs4MldXUt/
jlumLaUH2XtvYOZvAD6fzNpI18xPfzA2o1crX7v09DPACPFRgm7PNAWPrakTJnq/
2sAhP81Tfp9fX341rodjnIqZgTJM1q2pnqtgvZQtWkr7UecB72KmyKT+G9mRV7C+
BU18/EYlO9fE7//WeOM8zz1Zc6mS59wTAkiqCu2kKgpaG1QjKcdM5obmN2d1BdW6
lWba3386qWxSyCkkm/ICkp3wAI9hmeowkCHNs1NdoCzm51z2SfK8jywP/ZpiazMc
fTGo2pFK2htjuKE5+hvYEs4ZwJYgfyDu84752FZexBFSN/+jKztO3RYeV6Wu47sQ
zQHWWaic65EAESO+La5hXfe6swcv7DGXvAW/LnX2ZjXE5nnXvzhRgyOIwV6KzXFf
MfT4s2uK7T3BrfVW33PBqlcmhsPaE7ZIXPdHFOnHPwzb743f+bqHjnxoje9jS6WZ
C/64+Ixr/a1TQYITjNvZ9tYlsFZX2SMHB15L2K2hv9D9sjUzUyv6Gp6LH1XA96b1
U+6CZn8fDl9q4i1+/+5dBOlrR61i8iNHjbzWcn7gQNuqwFTm9MnFzE7hdnQ7VtYT
doApCbhMOLCDC1JjMMjraaT3PSbQmFDO866hu9OMvP/aZK7i7O2hBjUV+99U9Glw
Od9KwFfNfq9JHiFydRX8zMj/CdDIwBUPy/dKDknxH+K1oXytLCj7KEZwPM4uxUdt
6AAtD7tDYxLoKJVwkOnLhbx0JwJZplAsgNFaB4rH1IxOVJDV+iZAD0Z7t7VY+DxZ
gbTr1X2GBwVRQuWvNDAQ+6JBj5JxwnweJIJE03/cY/2lEN8KlvvZdSo+vJfzfghj
EWHA2Njr6f8CK1J374X6WyltvMa9KjTUqQ5+QZgkjeJh8rXr7OMxBiJSDOc/Zggz
dyIvSsdZFSEzDDWTyVRRsmUZSxTyHtqX1X9fpx4F8yGoMdrvLp0j3JRFhpARWoTF
9/2qghZRgUr8/dt3VQmOPirCBH4U41OBa40i2DD7/y9LK1Ui4Qddwjc9NzMZ0qJV
uClHa9S8axNuojGlb3yMTtOU/9xQGKCRdiaWk5wBduuArpdUWIIdjewJQI4iyCvU
PfJqp0yZ31cAj6feLsz+FT8hlfgz6sbj8BhzeYMNHtq//e4hSWy3Wi5GFl2f014K
crKp4Uk8P3BZnsfF+CtXLwvr6wzRAbUZM1/4F5TMglcgaQMXynwn9yx0j9ByY6j2
szTzmUk7BaGJEJ5IkjtLe0V24qcQFs/ey6QcKdSQUF2OyUrrPSk+k+atX2cOPZDN
buviodW7TPixwQAF1TvOF+lztdmCeDOMCi53uIh1M+3yY5PSH9EYbAw1TFKPvBl8
bGV65USC8S7bI2RBZ/DTeYh0Caf20LiwamutsL4ME/ow+k6Eac5Rt9Y6Rwt9qxEw
cCL777DUW+wLUWBAIdJby7tQA+gWU3obkymEOTIE8fIRabZXCAIxDT+EX+XHqdAu
B+6J2Lp1gX5h1QIKULj9qS68Vn4Rhgq1T/rKAoY3/fmHPE9SIipSPEfOvdvsHPtH
Tu8nZB9o8DsT9L/L7ehIl6jtWeZedUj1qeP4lvd7djnsLnR0QX1he3EPaRtHx3Pg
Zk67zxNzO0BkMe3EzCkAbIUPFXRFMporCs3IpFzkuVA/XCzlKLHCdlwRYwcJfVbi
3fupW5uWwGwc4i7PMCldCDvmz2zybW1wIoKZGcZ4K3hBJC8b2xzZMJmQpIkbpjW9
2k4TPW0xfWJn7CKeETUgmfrTGc7AmUPiC69oe/XTdS96fphmGY/igWC86YK+0CVB
ZuGuf0lMHJ2kpnihY/rhbYkLTN/PTEEGBgfDlMj7cQAEQ7q4wUba59qAcciymTQI
DyLcyVZm+hN3jyhxL8ZRp2rCifclBulrfOvta+JDS+ikZvaecrvK1ihQWc10gYpc
Sa4UrWc+alezdbaRvoHw6nPW99I5+0Q/wQFzO0qSh6XLjGA9qF8chi+wkidutRFe
5c1WVJ8m4EgxXG+ORSaeG5s2aHKJCsIPj8Wblzx7yM8IpNCyTLS2LVDZGUL3d149
lYfY8bmGUlhUd8xsABGXGREQhPu1db9bYwQ0awQH5pf8aqfVkaOxVBzJedQKjxtN
zTSafb0LTMme/ZlHaVv5GcNNHt9+MY1uYKkMefZdhN/U4mD0LM3AzHk7c1ExuIiq
j3ho0gCSl8slqoY7/NFCzTwR6P223gEWwwsFBX2MYQN2A0hr3y8dEmrCQcNERDyz
vVSKuq/5SX9oi9jvo2vRbNo5FRz44U6wyp4qZAzv3S5tHXzW2r9SRcc/rCkm/C0u
xg/D1KimiUmED3jua4y6DTX5Mq2RuMTOJSVFCZDjRcURwPkDgpgiZncPvDADq+HS
UZbKT4KMsmZCs58QZpKVCxpBDicogO54PPWNs2egi7PKyKWGFNF747k+yfEe6rHy
slWgtYHr/Kc6/Ouve5/7j/coWLB5Mz05OIWK90LikqW3jnW+MbsTTNBrH6Nl5yY8
dNLM2mDWCGGykOxhGiFhOIAkNFUvISi7UtuL16uZYTO9tte01nPOea0Nr7Pnt1FT
ucKgcknpwajZCdUvzZf/HKwnA7xfViC4qjaAkNR41Qya7aBwQkYjRS+Vyfvsvjbf
w2iGom3xVGftFD2w+JtdJZ6FCf2MS+cekSt9h7iXvVAvwbUlinfrvZ45a4bBGiR9
c+Gi+qCA9PNBdjAueu5qgCfEy6lGpgQNkzX5LdUz6ElwRtF2w9ULNlsbab/+UT9l
0UXJztZo3Yl4HcdCCFHOJZEolk8c+/MJSnQXl2ILTM1SnbvOVQJWR1aEcu519gyp
Ljkg0jSg0Nk9Rx3thC/YuPe8tdVKUmTQauFrFYZuh0robpYNRm2p2v8Oi71b32YO
bSMdtN0e8HFLuwzzP+e3sK9JAGIZ3pYTEraE1mC7YlqOedvPuWjRZeZvfnTJxVNM
N0JfQxCKPKKwdYNEm+s4TE6QyRlnynUlX4uFJaiyy37NPgKoBcsDPhWDXn8NJDlH
NZURcNCyfLFPjCxG6hK3MFXteVznpVHFpFzWYiqLOfVVXUSXOVWq+nnDCzT1qW7j
RXrFJ/fML2V9rdWU4e4Y4yEZ3in/jnhdpmkz8G+R+8iu7zVIvHPO3moizFxtHffM
shmqcGIFD1ulVIKGFyijgySQUegmrETixQgfXQCO8DnxHUn7DoYCOlQ/HSDCw/NE
n2Vn2v79yE4EtygMgSXnn9I2WweiYyj9dgKbklEz1scBIch3XIYGklvX3odA1NHl
jt/q6+SZ/reykg7qs3XkJIQMo6AVMKvTmt2WoK7WNSYMKImGbSN9y7Ofo6YSMzvq
a31h1P6LJjWN0lGTZYTaX6C0OKrpGAkX+nSdKVegReYvj7zVbomDf3pLE6MWNg1j
pQNGujaMxghGF7tEU3XPS1vpjZo6SevCcnKP8BjKtY0xeVP1KLzP2lFYssJhmc6O
Fwj4xI7idgW0WrrXTKDAbZ1a4w2S+E1W4OT/FtBqr/GiSbzbreZeum+s2mDqkE2x
zasN9SQNl7pgx2PY36XhaTN2ML9V3Wsw4sqYsIJj7K5F/VfZm3Rdq6YOhoMYV1uA
DOENcuiDU2NNLMk08ziRyraTVRJmYAhvFgfiZ6yaOUFLt7Kn+ItPnz6Uh3MH0n5C
rntVu7u5Wu9z+Ul4A/xYuCDA6MbOIw/BfscjDzB0dlB1Lu0HBSkBoxQmJm4hZSAs
Obnqk3+54lYI03ChRMdNXrH9bonboYvliS14QKDBWcjVJ+jI+CSenvkish67G3cH
ENAEBJ0KTIULoHzMZ/xb+FbhVZiZNihGVFH0qxXF9yeHAOCqb21Y7RXNl6eMlDlJ
vfhOP/L9RfLGttBS3UW1AgTIGFZU3z0aDR+LoRbfZt/8tUOt7m6U4NmGWGO/QjZk
P6OlL6ANfvUas9/HNaiZAEXuAgrPXvoC+6TviXLgcxxzuk5TFywfuJJ8+DqxLmxC
x81FPsK7kCiH5/Ww50zecvFEvf43MlItP+QKp9CS7Elbd11HxBqv7bE2AJKFuqKT
wHzkhewpLmbUNC8VeEaLRVlSmnEwZP8h2MuFRbzgZcmnDhg9jXkhRoNtiQMcpgmE
gfQYucnAD7OPkoHAg7rW29CQ8LeYtn7AXT/uAby2gnpuKruL6WnyUaKyu/8Liuxd
vxt6BZe79CD5I87k5Dg8qicfjoQgISm5QBokRn/xXaloc2Ny04jNbjb3SVsqntpr
78blSItsAxu93s0bRaAMAf3PiewAWUvu+qkUEVqN84b+fPxncKBmrBwzB+FEi1uQ
agdbEWR5F9e8TKf6gAu51rNAy7lZZfrbxcYkAW9KRcwAASkBEye5fjk7yG+qlJMW
zMB7Nf11aeqxyoPniCjuftnZ+79ha5FQ4m19i9vFzQp0iKUPJKzr/zvs4Hlbdl2I
zjDeqkW8shPmBxH22BizSN0SxSCV/iy3PK2UU+MTf0oiqUfVFiZPeVReuYtFQ1/9
/sOx6T0+ooPFLSZfFhr3dEUih6eHWQ+puqa09j1SWFl1Irg4M69JXUl/7RDk11Gw
8IB04/wHLHxFcEjGVpzlNtgAlfL5OD8gKvNR2qb9ixEQSVYB8Z1g8qlihFiX4bfS
XmWPagOWc0mxEsIIcZIkr+dSHeY4sPqeJvISjQoFz2QG0SSBSCJoakpV/KCOM8SA
XxDEHkN9r48MNLpIyWu8M9Vdb15MyPye/aEz9vOW14Mvp5VbUM8I8ajVYbqTlvsd
QhbxWA9viFQu3nWJdKvY5Aygj8N1tOblC9TDimZB2XtosBVun8hJbp+OEkfTbGel
fzOR5tJv+GKPDRn+iVCq3qSUI3AEhRdopj3tA4c3Wp9RAoZWId/hrHQZ84ikxAAs
Fk/F3ngK6idOdhtku1EjmbCpR3Q3t152M47ZnZIRdLp4TU5LzWhq/woKpBT+zJb5
4JYc5CrYF1FDI4dDDOF+hXmSpzcyfe/JNuBgNDlXu85qVhJ3KaIt/W2ejGXgypny
ebJ3DOYguelRly86nKUFnqd9dmNp7vkRALORzDcp26E0RCXJzOpfSHee0kHYWD0e
nIPE1RF2yOzPNjT8/qdpPQG8FJC5G4dbx0JeAQ//2TQ9V1NSGGcRP4yOAmRPyiNX
M/OI6x7+0HCVf6+HqQUQa3Fq23WCdMEecB1qGj2Hh9GDrDgRjc0Hs9f5gilVG+2J
3LXEb5gqcRD3MwZMhdySowPG5oqtMrDgoTZulHyvDqdIgo4DPaM09oLKDAIsJesw
RIzCQjqTLIgqdU2E2hIwXkKWBaC8HYPffOBSrmmcCjMEFWg0mS1lWY1ebqwxhcV7
T48hZ0RPlin162ZafkDKqfBIz1SnOfZxb4hkNEUzu6CEUFRmUyqsQtJXbHrY4oTU
cM9ZcSdJM7AXGIt5AmyDLuwwKsn+85pcDxeBd2Oj4QtCQox5U3fJK9V4etfX9wsO
7JrFqzRUp87wPRAoeLrd7arQQ/dm+LYG7iN5BZBAJqhWuyxvL/tIKS5ltfz59brW
t7CySAyj2yR0aKoq7EfqeBcfogVWDnweQ46EOMc1GBgdKyHbcV+IhIDf6MWDXeoJ
rI9a3YS2cXhx4JS9uxaMbZsH89eyrWXSsJURxEyKiiAFzJlLuD/jmmCFYFU/rzfs
Gsv8um97gtNpD0v4gH2Zks1W7N6CeiBd/hEv4ChYpG6utgcm39bLPDOrrX1tBFWe
GFtMZQktMil+LDf/y2PPjK8+RF2+MCWiX0/3m4BjjV5ovG4vRJ+pU1AmDdfrzSgx
7bOklKsa2iWIoUBghmyqUjWApjRem6xV9nQtxzY1U0FZreazRS1ZWu3WzFv5z2VG
YQgzOyp75b0hFa3z0MZGYgF6+pmaYOt3j4/+LUTjNXP8bn64h5xq1OJ6ijN6gcji
8RctFTjjl+USANrikMFsG9RLqQfZa0R875U0mbwuv84VPUs91sdxiM2XSNMR2ndD
mrQm70Rp1hYTRGNn4dV13tIcxiEWhu5rigsAPEapOZ6pgIoUDZ81cdKhAu6/nNWM
3U/Bg58z8RGijNxTf2YPv+cQWhFx+bsbAPIjcTkN81AEqqugK/dWFf+Dw2jqYZXr
vW8aBGQpn2gr9486r61wLqtNyPmwmBUXBIiKPfH2l+OpOuviCUhh0Zyp60GEiKpF
7aeb1ZXldIkYI9WmkKktaBq2KIGu2CpdK1qw9jhtXH8JbwX8WmdeeJj9/fnT1uN+
9Dl6pMr583MFoLSa9JPhUSFz60khHggWFdejkfJ6Gc24RudkiF/00DVmvcU6kc2R
xK2Cb4b+w+3rH2Kx+LMArQPDzIDAEQghS1dVsQhxLow+tN73H5vpBW+48YmUkOfh
kM2dKIhCd7cDJRfaA7Bi216qw4BM4n8pGk1UGp7SMRvoyvfIk9artcnf73i/lZ2E
+LDxNIPG1huP4ErTUkOnAF+SYwO8PH5RIxhQ1HMf1BryOcsMfnGn9Sme+XmQi1Sq
pAESKIiM2cx9d58W6bPa6da9bsAfQb0mJmhCtfacz/2ryzHogY66Ay7Sk65/rbu2
57UUVZP1EgOqYtbdKRFl1epf+5SjoFHKttrL8VW5Sc4yrQRlofq8xVBuD76/T/zm
YiWObpbKQLKateeJEzrIQMxGX8XwnAy04CN1/7K+OukwxLqxkuDmIilOFs0XXka/
NGWCf1l6Ne/wwOGpQtq83dNmi0bTkvabFvrIPfiQZIIldXB03qpdzFe+v5oUU46b
WR0oVkcpkFMUJaxmBDruWn97xUF/sCASPl4+asB4JLNmlMC5YDcfDeyEzCfjiluH
nFeCrsPMfbkEBcPN2C+swPchjtowCeaVrDbTJ7aZTLtvr9uGb7Ix2QChQH904zWl
0ZOyrEpXEJzEkPOKuEyROf5bow0JyQEOykkLlU6nq5nHCuJZ1zNMsz7XsNh6gW1x
RrD15RZeYON8Ms8KwqNp9tIUR5sTVwGXvappugISjcS6DT76bLRtJSQBZ2/4kNrg
EurlbRdjLiBc8SjDWNKJERIvojcyfhTcDrmqxlxc+9dyDFtpy8LNKRSVrDLr5j0n
d1P3JL9G3wgtbnNNqpHSTzYf7ekn0zC3EzNGJE2XOMXo8W7pOwIKa3HbjLz3iuQn
C60x9ujcEwn5WuIlgpKtckpQ9sW/TFitpf/uBfi/w9uHoiexxWl/tsPFjXQkNiP2
aaEgdI9X90bfXq/82zurF49vjbdqrJgQaCs5CaCjfg+CRLaCJc3BqyL/kyCO830Z
Mn/5g6btXURPcjSNsPbRgYHB17i5B2W2dp7Mh2xBr+h5gFeOwNOCWWlGjUXmaa9N
D/GZ21tsSoqdxrka+tRSsdZVysY6BzFmAg51JizubF4mzC/cl1IzY+q3MUUiLMhd
s/vb/Tx+PamqY7Qzwb5LkK5Mozdton6uzS0Jofk7FnIX3E2uvD7Si5OilfVMNsCy
JKHhrG2KLiw9qauI++gsbRbkxD10qWHR4KGJhpr84M4xpVv+yxepHoCwc7wFCZxF
aQ0RvuuI9juWw5+uwMvlkOsVr/ttwSup6L0w92dJsPatCd/aO9omXhOUwg3pJoe5
DxLEz0uixPPVCN2PUhy7WbADir3MTaf+crMSk1C4PW9SQlX8m0pebxHFxSPeGUOL
U5LVTTkwLFVFx6dFXNAeWfs495eHH6mU9fe3OxVYptE+PbJ6xaGlcHoEEK2Do5Ou
y7QDBtDrZBUZbI+/wcDlBxxcAM19VgVYDYJO9fBVGrM9j7AuLZQ4jpbW+ITw/qzW
FmqiZktjIpyIrNaKCxXOoT7dNcAyAFWfasLGSYInns+0jktsTtlbMTmi0ENchp/G
liVSby9OnfTO0aWoYi8NUsxjhDxaIKfKk+3AlRecvRDG25vhfuVsLL8/nPSdggwC
IO6OlCxsRzPKjDBEwfYlj12Eg7XLic70ZOg4SPWqo26SnhzuIQDqvttI84TtxKc9
+16Xz6YPTUxg7XKQvZ32Lg3cDiFbOdEeORl3oGo6vPOT/of974pw2ob5QihcMGFh
jO38URZNIttBIgIBwl+07tNnoH5cA5dsj+ZbOfllJNHCLsBAOR+tkj3RDZm5Y/t5
ISrpoeyFVGY7oodweXLoxLAif+DVU7Iy0XtJf/SSuAcmcDYSRqimijuaN4s3sTjw
M7mBIP+R5zjQM0xDrbMzA0pvgNN6ld1gr3DKhDXCCnS4c1GpsTkRe8W3emSLVG+H
cpvEwLaT/D5S+goRxmXi2OlUiyVwMUIlRq8Hik9NsWulc5MuacRbh1gN/PdTazCn
SK7FjeriAGJ/Mx+pP8gz9SlzgBAWgwwokrBqxAvrH9Z02GKL3/IqO9QfcitXmKik
RVcqe+d3QEElHtzevYSt6Tj6lxRzysF7CsryNq7u8IMD/l4XrcSrWt7v1rauT+RU
Jem30Vc6H0qI8/uhBX4zgGGc0RNI9K0y0UuvxnK5cWixkmpyvBF9/ObHDTgwQSmC
kuWIIFbOZE5IIZ/0Y8MXdXV12Yxh0TmrvQQP6OveNQm9K3HOEv2qVcn2KlUbwteU
u3/vTkZMPe9xaU25Kf0F1e0WPwssh5TADS25QEC81XWWKnH6ifODYE81WKBeqvGv
3w9udkkxbhiefZRjPD76K6jn3FXySOOZp8yLkqHuZh0iciq1zFk075J0PAnpi0DI
1GJzv6JNaXFcUq19ITckoQQfxsZQAlv9YvvtqmfnBqcfhjWgwFiNRbzsiL8DcpQG
2pScKR0FmF7U6x5BJm8EDE+jdA0ekKLIam60mOhQ8j2g2FNxJwHe2FPtrvtC+Bki
SwDxN8a9NBPFeZAdjERwDoHjnKzEGajrcwETLyOkXe4Gf7nvABUYZp9av4r4P0/S
MT5kJMp1TyUD7tBE0QmBBAjtCGl+tVUlrK28ZNEkAFvf441r8pU0LRXoY4if7mdj
HO2UeVdVn6Spk7nVlA5/2MO40/z5xM5p4h98tpI3vRyv2GM3lxmzhnitDMSWgz3s
rXf7MKoqf907DJKaR5ZOp9VEBa1Yx0vpkBnaDrnegiqpbtvZn/1AoTF1vEAc9rmp
zPrxsuZStFKSjdwVcZxdM9kgd8yK7bbBXp7F4fNkudpqgh5cZNzz0vR8BfiIj2Xr
D8eQFD3rr8ftkr2ioWYNUX00BSxTseEQSgk/5Vc3deF2lXcHpd9DGkXMFjklas5m
7ErIXJOhsEizJJl37xvjvlI8BxZWmuvaJ5E8w5Oup0PSJi8fHuPbVdxtKfqcLw15
J9Vsu5WlZ3GvVg/bTLn8GxToBfn+OrCaHuRDv0xEg65isX8wUVbbOO+hWKZRP9NR
Awxxmt8BKX0SX/UUbx9ZDj3oaB1exsym4663QdHUHP+1zBuIeA224HBmsMIMiqMd
uyZtA0oLOdpq5sw1ist3ipdWAn0nIgWbgKdl0FhfZaJv6T5ydA17Jyz+CxUQt5jq
V7C6E6+sjS4XWuVzMuJ5uXt4HnJLWO2Lg+nh5/WooSq9JmJOISay4hCTiae7qLIY
W81xhdNOyMY8nWA0u8amaLVFrCyba74MwngHvIxTr4MK7TPYmofCCc4UsZt06mEB
T9ybmC7ADUQ+QKAWUspxEzTATTNdJl+oGD4dkNT+wgmO7rxSdsAUB/mvKNz3CHOw
UbvPdbffUb6giwa9/ODCX30UDeZMJ4gfDMW+J9g1eXWtK8PKO9Ya+Y96/3wBMs/V
MJuo/Q+57XK1FqpFFNvPVGP8NUd+SmlTVzcxV8GwyfOf8clS6xRWtjIbhZDPPW+t
b2fEwUzkVosZ/kz9WurUPHzoPQBlwc2dMtOqgB94A5aPKY3Ffd92MNTeWN2BthVh
AtIGjTzn+Q4gRSmyJ3Kwn20MIoPDaY8XYMGgCG8yoE+MGEpsGmc/9EeA3BTiL7/w
xp58S41XSoTRJI7XaYqQm3ejKpO2W1TMFpUwhmqPQdQtjaf4bcODsoEsYs6Hqvyd
cJxFAEeNHLeI3ABYYI+1hrqYx8CNuJgML4gFMGia+ukMwPqwS/qZY/AAjnl1DGoP
OYck7ksmFR7ld9wf08sEtTOnzKXJY/A2X+tbsIrTVR4GxtvSdcnB7qqRgvytGN3x
RSVrMkATlqiUE4FuDARGBbZv1NWaXSk1hcZik4ybmaK0SgkaPCxRvsOiovZCSqLm
JEVad3YmzqyQxEijoZfhA/6ASAIrYUAroiOn+KOpZHGZ4NeltaGMfpUrg9NZriKo
mvsHKMVLpj8rC1IUuDvPdB7RSWcdAIGMYscz+H68tLhOBzfmZm2Fxblr7eGotgmZ
582/CurWo9YOE5CWtp0g1+2emtJo/yJJgyWQ7SICOusfLl9hHTZ64DenGAY1nDrF
bsMxBLUClzzENIpBIL6zTF+3GESonqDVTy2Jm2oy3RWSOhq/2ThVFk4q1XTHo9u0
liLvG4lHqsVJQEQZufOZChSjm8wZZNEKrztIUG5BURnrFqw/zaCGIb1oIt1a9irm
XmKTjLiqupuKM02yGzRV8y4isPBopFh+Sz8buiZr7G9s0ZyQbvlLUZvomi+l6HCt
S4a1heBVmw5t2Lfx2WTfmoDTEsplxSw1P3JXBiBZDcLN9y+stS2Tru0waHeMaW5z
3u+/+5vZlXIUxVYH+LoRbsizzMK+WY3t+z9WJ/VjBQV6xAotBVw9kFm4tnFEwBqh
9M9LxInM6OzhMY5JGHLqEIXa0eLPnS36SUMWrXB8z9Bh7FyY/KTyRPcUnPP3z3jV
w4GvdCwud5LgL/EPA5WYaHvenTzpllBcPat7/Am8pzAhxbMLVKFTxizofB9R1Et3
h7CSRZio5KwrqXg+eNwgjf8GdwMg1UUgynq+7MBlQeIfIjQEJ2qbaHWcBRSEtlWa
H7eShQmuQ6/Vdc7T10BYFxdBX59WN5HuojWp+fPOZlSq5gL3E2m/Y0mbF+hfKP57
dhPK6jMh+xG84V3nBBLEw7TPk/sTMuea5A9qslaVH8Rx78Q8KyouUYeGQ4V2ZLee
heslwVDWI713hswgETLIBUxjvBlJlcO8GHWp1+aanaF+1wnQ+CR2aVZ0gEsuEO1R
yVVfSvlFrjIxuma/TnAcWo1BkVDdCULkS3JatNP3XLqx2bvteqGhM2jHZWYzGraB
syB+MQRGGvYzXpAmyDDYrdB/PgY9kaJZ8v0nnzRK4T3iYMcEzRGZomgIU9qEhhV9
UnGeggG0N6nxHp1O+b0895KB84g+wQIGR2+luq3jcAN+e/28AbCe77nmaX/0qgXz
xXDlBdi351De/NR3rVP2i4IA2GO/nIG4j+blel9REOqu4ECZOAkHKtPdqvmBxdkW
htx4utY/U27pELJAPQNg+CwqkOIW8txaIzXHIuM456DabVloRuURWUUR685zNOAa
Cn8Et6/VUPO46W40pY7RVsl1Aqp9zNtrfgPEaxYuQ0/12eYvF3iXTQljQq0g1Ic0
BE2yxhmgV4p72Yq6caiT3GUWfaY0C4PeQ7xniDzmZGvUV6B99k1y/5TmvL48HRkD
4/jhIkQt8iJXjbI6YjvGlQzIMCK/s5C3StqgLNFgj4TMUluHKhW5dXGSwrjPb10m
Ee3OVI2p4ur4eRT/+bKJ9otfITrnmPf/2L8Oh3HfFnPwUhfw29PxDFWZHgeGCUmY
xMFYsTwIuPT1JSCODrVTYiqUvV7UAsvgUY7TfnR887iIgLhX+duuNK19VCdAvfrs
79R+fOh1Tombz15cHf9syrw21lSR0kbtUUAcwEZrocHRkli/6s5eSVS+KoJWy67k
bkARpqDWrcfZF82/p6lmQ/o56Kdfb7g264TridPeO3x3TNloq+tDju2s79J4rDd+
kt9JQElhlL/vQOnfQxob7V+NdlT4HWCYUjUKQjrasXtcVCV8tdNXu5/rHC8rGpRE
Mmvmjh7wSrs8PjhbbCEv6saNy5KRQ67AK6swwb1s4J8kYrPQJgdGTUpmBB9oefqt
JPVCgXa0mJcV+ORGaNalwVcjkjrNH7Op2I3s8SV7qgqxTblq1GdVIek0+EO0Iy3z
Khfp0szGOc/z6jtK4WHLZnal036hKA7cSy5Y/2xiGz6L2JLfm86qz7OX/Zhe+Nek
42QW0CcWkWaCDGc1gYr84acB+Lw0uZdg9/oW6hi8Via7qy/VAptjoeeARk4pPrsW
lD52xHZmmVkVCVs9wmfMedrP8qVWUoA8MaSrmFDo4yt018nDgEpzFJFWhF7tCn+s
r9m/6pWCX29LLVKvyWuWjFZXOk99aYIMEa4uIlw/ao+YWQQ5+vsVunG5vbAQsMJr
0BcWBt7iH9OjWMfmK447pwP7YHEnm53ks4dp8/80fBJzIVcwYVMaXoWFJh44rqKj
zLI89qcYg+AygmADRsYvQZ11Z9aqveXmK7kkIsWTaB3xdi3Qzm786Si0MgO+aQmY
DLrItNCGnO6U+dAilFbOKQ6rbGyN/rvREzkaMTaC7+xE4hHDIfxXVl4muECWJSBv
D6hZV2hU9vRfm/7XJElNvRl8kw8ZCKQSQOjbUaf3V6YUa+YT782JKfGsBiCC5k4/
SKYmibnIXiZFM4a9eNN/vMlQSIpv2esm5V8i4+zkFv/7Ydhixld2xI5C7Q95imKc
1TEUi++l/Ds4HvLfMdCN77b/54xG13VVP6A5WutXoNDR8fDUSFIEs5/9lvshL5t6
4mo7fod29hIB10CzqrB6Tcv+Pv2oF2cI7etF7xvRvUozdeyX/cUzll4D537rPPnd
B9MB8R3RWU5hevajE0JVS5TtKT05dk91i0CyCglFMJ3ZrXxAimUT7cbg3ugsjqJT
zdHXTIt6ggp9APlb2/N4dn6LQx46EWR50aTw9/zq80r2RFo5SqHrL29jiyxbdwZm
N58wby1DbQysAs6AIErAE8wJ4EaIaoQxsggCnli74Co+YOnRdUFC5TwmdYJfG1z7
DQufiZMZT/ak+sgoxFbMrjfkmsQeOrPRWDkMeQQadwphD8DkJiIqFzsfjEpWg8K6
HTTk1pr2WCWdA4yXqcdwo5Fhkfm3h3TBW4unt/ZuBNJBfvNJttHGzXf6tYCevqVK
N04m7YupiF2pC2OadCzT+58FbNNcnMV5niexfygrQhPQhK6axZOdFaWrp/HALr6T
9Lp06Mf2khDwj+rUyktpF7/upNF4jQ7Za67vGfzrAnxSIWmBP7maHH4YePd+NgX6
aPD+wHl072k+X5oF1Z0cwQuXW7wji+xwaqZdq3kcjMPsUl/LOvF5kttTcIJjBRt6
6gVqIm7ShnI/Pumos2CxLGFqum9qiW6E5gjCRCXJGy9yGXVRhNW+A+45A+T17cxU
0iliIpiVagHmoGRGJ+hgDw0+iycE1uzp5NIHOen3gUAkWXLlwMwNnA7LROlT2viS
NycHkumSV7fs81559Z0AktZ5zgKo4SKTP9PpAfHGnh17QY566qChFBQPbLiWFM27
iOa+Nh5XON8IObXFaLTC1KRGd69gvRRxjkzpWu610ZvlDVe3lYNA/ppRpaI3KgvO
6pD0fpxrOaP/4mXV8EB5GJJ2YP5j6T90EPcMMSYWmCJMtqD+JRC5Wrm2Xn+w4g+D
Y+Vn019UiU3lg60oevCsxKIWvyAx1jVYN/RXpsF9IvWpJCIieuWh+yBmsYD05eFD
99IZBv1qRktKqZ/5XLZ+UTJGpDKFxkLZBETm61se1deIeQFX8t+GM27MsZeiqnvZ
dmrX5ZLGRztXEYwFMaAwbTZghYILInO2LWw4DKZ71gSlLsXf8rzzUzWFmL7Y8/mp
5eVYcqflkGts3DF5Wz/ZOvxjAX5hpKqs1N6r1OPVJP3qYPJxdg/vnHgsOsDduigG
B2kChY0PyAbK3vfpp8ppas+p0zfxzPClOPxFCBldnqGXVPFBV+o3jc9vNQldxv10
UNVISbDtdu1hsVJwHAWQhNiRMVKLdMmTJE9t3+OTxkrV/fH/LiUFqJxmyuKhOZ7N
n6yVBdnMU4GZKqNW8NiAvqKBiXwX1uRaNQPRDA+VOeE2k6KdJWQ0dbqkoiceL6FC
fKOTBAqQTKJXp6PzymoL7bEZ7tMRn6X3rgrSd+SWxBpnVKHl0tWtsUcKBPq7kf4L
qzxI1uxWnQN08XQuw2bDM/Npg6KgQcfOjTZ68ZZf7FpnxnUpTgR+/4MWrZmfLbLY
CIQ5Bwm5z/nDi5bEyhheP032smKR0ZT0/xcrjOlUyb3dD41fQU3pStnyPXU5G95m
vUE8460+FQe5PZ3rfOO3KbDqkfImMQsQfuEvMycB7s3O0rJl1C9l4TWETx2QSi8r
UdUUJBfJOQwfUbcvF5Dq5rRR71f91ZHflkPWF+XLINkMGdA13X2DVLhnG1RHrQsX
XbcfBKp0d6htNwr7TF3fprEeVd4cOXebvE7NgVqsh1rXc2YhvaiOIc22m+uB1HbX
H2hi0ejkROTzHr51HXWxyWehKTW9cB+BzQpAsKhWaRQtcB7B+dSkgaNaa5/zyXL6
NUUwtVPVNsBNKrKPDK/rAy0mp1w/BAL32Z5u4W+INXDaUJz5Kx2drasU5lYxV+y6
a39CocWMrJb0J9Ok2J5JGsu3oJr9HwtVahOhJyVmeeZss+sBc31XLEykb/HFF9XT
2MwtT/M9YO0ddRwipLkkgRX9lrgxqXYsEILu+PDjdKPXyosTb4mXNvHhImeM6V+Y
gXzvx8gBppRl+4W3TBZaFeefksSSl++GZZs17KH0JJuMntzY1kiTI4hYNopxpxkC
sYOt4LrToGBkVYweZYpHmxi1lq/Fk6vphJYeyclQ0ixAehuD8krVm3RTDiZUbg92
KeDZmG2ZsMDYxEQB+IoY/5bsIHHx59SxitcXTcBTxdRO7hjJMZNxKHixJ1zfEMRX
RheLlgogUT6qI1MHGsZ8YdxLIhN2R/CExn0LMH9Vjr3mOng/AYNmC5HZUt9EnXIY
Tf3kJKdkypRQBeIygJxcHYP+0Li4l864gsAPnZPsCSI1pAv4WXuHAizW4sfOsH4k
2uxv1nJ00YqZlOsYaXaY0/QGL9KMtg6kM4dLV7oMFTxv4h9xa+H6qkxf+DISc+0O
o+Z8HXFwvmf2EKgtaMz9fFDx7h20HYNAtmNDkA0qFpTfCoIll8sEUBjJFhmd78iv
fO5N5AWgTkyBXN4oo6Fx6isJ5BRpIbasYdumyzv9YNbTTEjL8w3Zeirjo1407DPj
vqyFJChapMjzlTLRxGodi9JbqC7cd+OYZxyRoVBJlGRMUkENo9NBa/ntNggLjCUl
JU4HGcgppkUWCwJeA0+L7DDHRmvJ+jNv+HGeEAY+jJiuLNVl/5hfqEtvfYrkG3AN
2hVKcoeCa+kxpvJJyfmj/EkWQoUjpz6dNzzpUIUbeQs/dOCspzy8X/nDvlU81c+1
nJJGYBnXc3ayftQob/yBP/lN+6NGzqf5YdR/Ja9sNDGxgorY2DA6dPYjmST2TrjK
Oa3zx+iYmp/M0MGOGerTqDvjtYLB7738PC7TE6MxnmGf4XWCHm1JfRnqBFmQ+GBu
rJqvsYFnWcOwmUC4ci+hwhuYdtleYuqD6kUoCIWLW3ZK91XBjqOmLhKnHpfdTZo0
K+fmcpAioAAYYpZiRhj2Ur7K+sPJxBAlRrvw6fo3u1unt9zN7eiDj3iY6ZHF6j7y
ar3k95aaB6v1aBQV6uCJB20Osy/NCOI8Zb9QEyKVEZVuvBIJjy9bglq9jCLPEJIZ
nr+4ceRG6VrUtBLOvCV4d4Cp6pjHWggMn//cmZbd5fTgxff66SeXRG0KX1Um5zoQ
DUIuFh3PVujIMlqqp0vdl2z3PHepg+iPnowf5+WsRJzZSvTnaxFHzg/Ut7gLYHIG
j4XtegVPfWPFMU3Mqk5SvvLO3exBD9KdEDM3OBLKtwlONihiAV9dU8L/Iu1lkh7m
iaUhObbMcQGILNgVOlewnNtq1J3hjfOmIwjDQQG+KoIGUpD9j1eYE5q3u12pydi/
JMPQEG5uOBJN9pCVYCcEr75q80pq+6ejX5YUM3O8csk+A1oxLJBED8qmjKFuL6EV
aFdkA7p794AkZJbvnZ6qDmBNNelBB76TLqnkVSNhOsln5mTQJhUOcUZs3UWIiUV5
8S0SY0JegmToP0RnmARGNBRS/Z3jK/10miW6Nrwdfcio4kiXD02X8oSyVZavipcb
4calHR4Bym2tfiVpo1GEncPi5GmMTfL8XABtZSbo3dyTTU+/gU5D/jD0+P6+v4oU
QYG92gGtYgb1Da2+pKWBAh49pD9kIRhUZ5jABhWzXN+t0RIDZFBaJO+Iy66w1b0i
p2dkJYLtIZh8Te74eVMYMNojt9uXHCWYaA+zaV/nB0z3CVvZ6D3EfeKNAonK4LEx
gV34dz7FCBlp266KKK0+rNC9uw+xXMmcGIAn/nIy7vcToUGKbqqVLNktdpaYMvtm
U44ySUZOrOC5SZ+8i/lZzfhJsrMZ820y521KlMd45r6XotGupTKy4KaCU+ghY+TX
oyklUH80bEdk0CgiueXTd9w1k0RUCSa0THgJJ3IeTbRMwOTPE86ry7QmTg2oLR58
AZpcWnf6FvpFEGOrMPTgAfcbVYPG7KSEmXQMzF5xWduTRbguVLo77NOjGfuNF7Ui
eS5QiNshMQ2A+4I3mp1dRfgR7CGjMIWbc2bTdWHJ0Ee+88O4FJ4vjmP0olZjfUot
0Smadv2v2Eky2jhr9yTTmguzf8fOShZgEGty0/RdmwRG/+nqhPNjuaGDqBrGhXM2
YlSXDHsCvKV/R4yQYQNEMDeosi8cP0Wk6EyOD70k0/xyhEN7Y1RrycoSWrfbv6oY
JvKKHsUdX2Y3aIRAZoGOtZsyJ5dz/Gka/9kF1mvN9IV48+zIQBtyqJEzXULKPDuq
d786HUK3UroeYYYQ57UQUcxOaXS472JNftuBbTIIHmfXkmEgG32pR02/faRmOlET
Eyx914r8m3OQxv6CI5DUNwRZO8s0Yfpcf242W88rG9YIQcip0dSGv+OoXJCKEXkH
qQPsNllYFxMrkepPmjd2ZwFsv23iLp0xcGSQ60Da0QOmD+Xu4WatFt36gdrN2vbT
Gg5SUk8qoTfnlFQmU9q4ovaohUybjK0GwsLnL7TDTz4zlwm8qjd3pwDxFAW2T/dB
w9OHz7xdmzneFf6WIKZRhM8hRMJI3zzEAsUOx8wGMBYnZRmkcJvcr8JGubX7FAWY
EhGQgje4O6HHeZH3XExft1tpTliMwJ9UDHr1L3ggEV0myl7QQEXhrXZijVBSvNti
3nwV4TZQSQdx6FdkKhWf9rK2I9Vc/P/h92ptcajk0wVqHm5oCUVZVNvXBREEVTR3
6ALYML01JuTVNM+jr9wXgKGvmxUmfpfHxamQdPYFL8YzOUUiMdIyR0nc5Yk1GN8Q
NEV+Dwgn5gKmDTGRYm1feEK8S8XPWTtRj0IzCyZQ8h6/DatQ13/CEZm9tBLu5dlz
sXBDsmWHI9K4DaVjjZvKzw==
`pragma protect end_protected
