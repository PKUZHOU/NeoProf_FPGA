// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dDmCnjSc9cJjfvgRm05WPsTb2msTLBzz7iXG7Ew1ufEQwn31Utrlu5lpcVZe
qufuykW0pWjGed2oK34JUvWcQOUT2b/GvU1XGrJ6I+GGEUXhW9qzFGBGlGJ7
KvHBqBCpEIPDWWCejhqQNRrE02Fa+2zMPOjrXdDJR8cWt+x6Wo8AwwuSUXVI
6z6ykIGMDa3EYCWFMR0r+4OGjwFpz4Y7GdWwGx+eBCqNvA1rYHR40j72H0fb
GuRB28QsU2S/GmlGJeAE+qxVcMPm5ZIyWmE9ENfGjPUbqU+wZIytnzJNq9UB
Si3TXMEagsd6hNO2fXycHioZuqBu+1p/fEjmF56vcg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FAiQ8Ag7TZzeb+eFrCpJi6N5mWyNHPBMEuZNYj7FyvCGESw4ZqaJegy92R5G
FeYkwqB0C5dP7UYl3HViPqVl8evyfTjvw2lYsohJP4e7xF4jebfm7dKvrAuc
nn14Qzy0FDawKR/nFQDPRTSJfXYL4oq5MhZHT77B7GV0I1OhoGUs1SU/8rFq
ciOschPuWwoSHG88t/APa06mRvi8byGC+XC4/EaKnlATPgJuHF8EdIkrSkAM
t8Wwk43USo27doHDi7RNGjFVcH5gZ22jqBCcqRKpRVEM+Wk8ijhMDCYwvXAt
b+vvzhvMeQsG1GAnl9TaacjSHfoFebXqfPWyxpO4Jw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qhtSsl5RTvTZJ26qXI9RF1qvGwAqi40Sh7+NVVXIMZGZPQch/DJMgOjVgJR2
5TAAqIT7lAy3ZPwQjIDVVp9zeLWG1MhFB0Zn4+9RAINDcwkuZv/q2w3kD4+o
oBTmW0b6xLOe0qHhj00JtFntrf9JvCIrqCApWz+45+Jpvh3zPtHi9sBI+qka
yMkNd95m7BdzHoidWNSJaXWv4j4nPDwr5iOPMQGSkGh0VF0r47gOvAR5dfZ5
YOWvn+Jdm/1ai+wB+E4rA9NzMI4s4GHRWpFojYcu7+SMOD/KzGtwDMbSo4SK
NaEBtorzHerk2l4zs+ISK69BWYz06mP4iJXHIwDAqQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pvuqLMtM6/e5A4i8+hDrzaLyWnpvtRNy9FlpG0YNBP7m1cv7fY+Sw1uDjEYL
umyHkrqOAf4yTozuBV/4u1CglvR/12wj82oRqYi1dSZe5fafQhJh52R4Pylb
7ruZqep7LKSd958GRWEzTqmjpZW6lIdcE6QSSRFySW82SLXk41w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
KuBuvjIvQgrteuLhiuR7EOHb0dJUtSIpEa2SYL5QO5dxXWNykoVUvdtUGtLd
D+szdCZ9ko/p9QJR95nIVSiHZKeb9KE/J9K8ctryVtS6+4kKGnrvgGECXKKT
Fh6ygzBcziD/OJlnIjapiJsTbbJm9iMs3SLT1o+ZpY0vjM4P1PyCh8ZFJKkf
9R/zsDSQ2U5FZZbfH1CxihWL0GlD/Qi3tJzAiMUu/VcG0tgo6gi6C+o0T0zW
H+mKwVmuhn96YnxsedlHxVqJ9+f1lPiQ0qTX6bM12JliXI/DODXpRfuRPaiX
8DzZSej7oBfcWBRHGceqgb03H4eyGogy0FfidhZ3lyjA6b9gtaQH9ZHcc3p4
jxjAmJJy4PkLl9lkbjK2q33d5RPFbcSyUGMYLKb6LSXN4d8yYyZ0DJb6+4Ua
qCsjZ6qXp1MoPKzvExru+bOgbsTX71PKdCwYDf7Ou4fOTrlLGao5UITxm/oG
8Ati13drhRjbnHh9fzgjT+xHqSDDUKV0


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KTMyAU5Bl+YuoeXrcaSMiML3fUsk2aPdbSgTQ2zURi2o+zyoFSIKU1PLt1Tf
7sFlfbaQEvQ6X10Y4nD/pHR3gqrfn7Ep9+NXNnVt0VcAg0Ygm/Jyt+RG5XGp
sJWZqcUZYkNJh4Hh8HQ6IEz6sv+T3OjICPQs02EqYvZe3Ku9BTo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XXEbqm46+XUrVF+Tkoq3tb5YHJkPipOB6UNSao4lyyFxcJFHMpOL1Q44yITB
9GYYtp4QoutJZSU1Baef+1+Srj2sEEm/usoCXCuuopGqtWJG9dfP6snpC1pF
hbZtKf4/x6Fyto8pSBcq1a4zEwHSjZUOuoUIKPKOn0tCA/rzRUI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 59952)
`pragma protect data_block
F3UwG3phm2fx30/RLRDKeKLRRFqw1VmrQtIMfWDCGPPszG0Y3HFUYGkZbWWL
hL0vREaLdur5g+/A+lO0qZilycjVTpCC1raWl/Lce46LoEo49UDkCTnH9VyB
z7r/5hbM/JuQczu4AH150oChdlwg1B+Hhj6JOB4DHpO2lm3m6+rFSc9Faz9k
CR4qprg70/2gjqzTH3YyF7qVWFj5PoEsQsHaXEdudrzOk/p4S9RBHI//LQGX
Q+7Csqzj49sev+N/PlJ+RQyFDly3f9zaYUy5BQpADESvgQqcZbRCpY9Wx7FH
aY2w2V4TnTDTO5lGlv1+zBZdIAzjXSmoFnEal9OUX0zypuYDpIPxqOB23xkE
q74TAsHRoTpD6cfYOkrtUxDccukKPOPcNrDm/6Wz6Yrm2ITovMy7NZ2zFmrJ
g6Gmn4eKXrWO/UDGTi3o2hxlSyXVJR5pkCoVoA78DfXMP0TjkiWrKWr/uUWA
nZEIEsh2iVwgrC3eSwUv09duPC2t7Cqk+amxdkXeg1jK7uk89FzBPly6yiVy
r02ISiXjrFCMuGjwMInfw2S83+zdQBwMk+8VmfU+5go5D6yehVu7N9DhhY5t
lRALThvmOnmV0n4VTUITOqhQediYHfzdnu+39zs1AZ6nseUJzm1Gz/esvnvB
d7ymlCbMgQ7PfLDEyQoPP+/c3ayAzpLzOpBk5yUtE8K4skXcqIwZr9XKPOs+
AkzB/eSMvrA/Ou44I8sgO+NXLfktYfawfkMFf+HUCpNjsiGFrcZNtJTm/21E
oINY33olh1S0qcf7hwJsY671d7A5kmFU+UyIHeiUiyODyXDDsEUgssYZx5Cp
CgU8CDtnabLghoGjhzKeRs+JGfiXW3/8WyVkxQLKagUIcqRlsMyy8YkPRodG
PI3r4EesDiXZNLJFRh2UXyTWLf+/klEE1ctGbIc38ByPvLGTa+EMeUBNVYC6
k70RCODbPBlkjdFT2jYAgFD2Okf7R1MvxFv24+KuHtiU3T0BmDBX1vGxXxzZ
JWbx3YZ8exaTQFRt/P2Y6kq0KIieae6YaXvboLA0H8UfuTlQDTdCtfMyEVJO
yn1W3vdT7JUJmCUq/SIs+SufeDuXpcrMvw6snJPEUeG3oh8HTKtN+8LMtQUy
jnVHknfPjRDAR7ttBoI8IuIVTfW+Ji2wFNn+4uwzj5beTafcmeoaODJS+fIb
zXU4aPEm+ALacu5fDo3MyFSo+vIZ6A3MqKj6Ht4idTJ0bzrQfJHqmlHoAOlH
QJMnJVs5H/EVwL/vijTfwRG8rwWxWuVBvVIm4TvH7pVrc3XA5pl7IoyfXr6o
WB2ay8SWsUb+cvXrzAFihNJ1kqs7pit4tKJKPvmxdIijcyTlvt9igvrFo2ar
6SFJLiZR5K31CyecjogOCNNkpTAXypJIm/dLzo486/EihGvwMpToiKLVDgyO
qXZgsh2QvQBM9iGc7Ns9OfM9mOrbUYqjzOFWL6V721XMsVJShvUamJ6HhvYI
JrTN5m2WSQKOkppw176UG0FZ76ED1q8oZn6F5jWeOulbNOAc1qgqHcjtPe37
AMvF1sA3W4Ef+YfKJ99QyaCiroJb1Fi6/H3ZWq95imyphzChuUYXceukSNHB
NFVQ3De1CDsEYnnOCDnk/9mj9haAKUT1lIjPqtKWgvpoaitwpgX4pj0F+yk+
T+A3iAGx4XJECeXcipsg4zPWd9YGvTW3QlIVcHjSnSkkO001hKSezzPhhrNX
B2XF6sYCqSmemKz6QP1ksZgc5u2RudTa52OQWR9GJBIqizQtLmldN1oPL8kM
qfogLRvD/kPu5Ciy93bSy13jCoFX0ohs5wCARgsvr/th8OeFAt4KZpwF7Jz6
JNNrK9t+6K0uS5tSHomfpviT+C99BH6AFguU/j5rMuJPev3RPXATG3Qmcn4O
bJu5eRZmDqqfcSqPruYj03N/psGPrqM/4kGrcatDVdg82OHfxx2MRcoHJ5Ov
DusoZeO4IfYW4db63t9EWNym7TUZiRYq3ioQ+mTeBDAi8IRrVZXoADQ5NZPH
IiUGbdTqC+4Dr8V5F61LtJ1qMb+hkEjY5uGOFshH58QyyIrywGDixtlJQPtU
WsbjxSTuq9WQiCpbKWVzrVuh9NdOE6hVl+X4kUfkZNyidCYDqzGunH3O4qp6
JJa6oC8IBprXbuE7zgkq2911hk+iZUF8KFge8Ih5p1JAV2ik0342xxTab0Ne
4ewiNs+roiNtcGo/Ts/Bpy73b3gYEY24HmC1zGuam2pVav4GtCybkbHmgq+M
cGnrFKc+Txr/SHZ1/Lm8/pjhogskeXVXt1sQW+srmK6AJhpqkCcFL5m5G77K
wQvbJ9vA9gt0P2RdD8w3plAEFI3C3vU8jVpdgWegh48Fv68HNMRcC+qC5ysD
0gMWeBTkBNA05SG+hoTFOCnXZyIyrkyPmiYoU5EYzWQW950niaDVg0OyXE9O
UhDq4XDg0XRY1lMlqNqbFtPPsTFFrWACDGxxDt2t35h9/qZY9c7i+gUx2SKY
Bi1hk81t5E856CuNTRlP3li7fkCQSfVMX27uuw9md6kFwsf4H+GCx6U9J2cj
woFhSRfDdRr1oPKNq8/r7Mw4yqZ4uBhrD/0PzKYUGcv/OE/n8jHztE9yalQA
Be/kk5lkCKVeFwTl0dB44lwBAFmbYvQlIZiUdkdmPNr4ftv2/V7l/EOWRob/
Ty85nkkyu48tVBl0XWX+bufoLuZz2BOPwSVRZ6Nx1So90bv8EOp/cd8zMXyO
YuO9JflN3KaAMR0F9e2ucXz8unXzbhS+8wjk7juNdUVGuuiy6wKwzx3exXdH
vC2r2+L0Y+GWkHUGg0LEJADBbS2duFLBEaO8VlDnJ00MeUh+U9HvmdmDL+8j
Bj0D2NOOUBvbUxt3X0JGQexioakj9IRL2D3ycOr3TvYbCE+dq75Pv3OvQF0t
Dn2D2yQ/e29PDJY/q+5i4mJ+TK58RPxL6VkVHH6OoLYRIyVxd3urbq7wj/JS
0GHOYorgZD/Cyruxc3IjO9wx55fVW4kO/TBzRGoPMoMdcdqwA8TzLZFTele4
bNa5nj5ccpjFHtIo0+kSJMfrqflySh3LOgmMwLc9gfmXZ6gCJFpmj5dARjlK
amzz1PmZiLR4b8yz/XqtVttXMHE5NVTx3sqVMbiv8KbKcgS7PQa7IyGB5NpD
w3lwGFeNvNgKhFH5JsTsa10mz7+EDuGT7xZir2U0E/KCg8z710SREsUcRkqV
IXuEgGMI/42mFSgCgTYJ6jhFUtI/U+0p8xmjssAgjLUnO3Wr7je+RY4g9t7H
HliN1wPypj3sc0lDoAIdHrta8a0+LpnZUCSWaJkPuwRUlxdZ0/qJg2BLDy3k
CviNtmLKfMNT79TTzYk46anBHMnWhjlyQ8lIHGF7yM+ImqA+kcW8ldHbQHcY
QuwoAdT//Uu/RyTcl8gRIlE1uAE30XnICAfLVOWrZ2KqZ2jnpH8adWpPRYjJ
xxJdFwaB6uUMOW3hJCzClCUZGYY4o7xLXD+U9OowqPcCv0nQt7xf8l9lYcc3
nRiAxcCkGfbLazX86k9xpUUg0rr+Z0px6ndJtPayO2w9xEjibbr8jYSTDAzo
pHDDY+wTODQ/SlXak2kC4cWluJcHxyI3QdNxCISplVv8jBkC/FMSHITbAXaY
RPeglAmHNvPNpEYaImgX5+ca0Jbe7kqJxW40i3Nsk+DDEaxCK4LUd1A92t99
G/wqsL//DQDyu/EHm5wYIaMMSvHZ1YfHM3YZONHmRITWGZal4P7XTGCvybp0
6J5pNsFnRntR5FMHfR152hlAnsUi0QG9naWI/0lPYYMETmK9/wuM8J31LtWu
wxDWA5uQv2Cojj0xDMV2Rn8snoA0mqEVE1+hTiA0J24MMXaEns6vP1+Cxmb4
sJQXCLvZmLsouRd/bbGh//IA62n0bIaJkpP4/bJE3c0mtORO1QFSnaSbJSHx
iI5ZqAl8cz79t+wS2IyrEkrKr7kpXU3d3OGC2mHpun1g8bSGak+ySN67Chbw
9XPxAcrXMbUW2uXREcSmQrBSJRfGdyFjsrr0ezx8wbWvvuWOt+KzB2RhftY2
dUjiwCXIR0tQcDGnvLwYWmp3/d3ac4SpwBoz87ipkWuhi3zk/HkbEmea3bvL
z1kYNoTDzfbZrQT7aNvz8okNk7lrH09qZXanQywIz7OYPpJh9iPP7j+ui7d/
fbzc0chHqT3Eo20i2yxen/bBY5ZwRcV7wTYVxTRtlbiZEz8cO477Xy6IK5qm
VZ1zyI6ctL0On4DKdzNHB5YZsfAixEREt5+377iF0S0maPXPWiUXiPufc5gE
C37jOiSx8a1/fHP167TR6B7MYjBuVsreZ0P4oA4zHxHJJnPlcv09+xwwbAui
ZuGaGVETdg+u1M+K7U2xb2p/VVFeyGV4AIj1UaaXHSHiR4H03OexlaDPnrT9
szQ9cp5jRHDoMVySh8cDQbvumxSL4rmqRjOXLLleUIA5EpjbbT5y9tJNM9NV
SP1J+7xM/yJtFj4LD1+XeFzkld7YXlFgqfJcp7ptzKDcxGS+pMUm0QC8+7NQ
EkzZlcCXj2MIM02Mo/ex/bNWMWo/XjMSkK/OGB21fbCbUWM/iTF64mpUgNaE
jiaAB/0cpt88ZNMPlGJBio026oRJvu1I2QP/GEe3tq7YXxoAWeFrf0drnsD6
JS1MzwP6Sibk0dNYesJL0rlqdjP8QQNh79IfcYR5TyvU0hOIUxJ+f7S0rRDD
iERj/bD8n2HPDuNoJXovUC3nInhFiIKYXY92IQ7FoVuQj42x0/pTVXnpH2E8
pt044gaiLghOpQan6WeajdxvNIP0kENXOGcXnXR9tNPd75B4T7WDTZNdgNtu
Ol7/Bs6RYu69dS6DQqDXJ8W6585l3o5OgPbj2cjN9JYj9bsnal2ruZapLBCO
JJw2TxiaZvuDUYvINDvHAzERQk4lUpKevz335JmxZ2X6pXFlzFvbcD52nPCB
bcYrgevMDVILJXBzK2X+kHlQ8cCbxkifLuuqtnpiygtoteaarXDKjqjRt8dr
kdZDK/Tnrf5q7vJ+M9BFCnhoVaG45aHkmhgEsmu7Bl3OMMGcVHYaFWkjp9Pf
wPr0t6hII1uqUf8gKozm3CnWh7WQOlAJdSOAi/iGluE3WRuORN3ovFV2OzEp
ywqIRCh0uBp+RneBgGS5otnl7bkS8lKxqAy1/k2mpx5kA5vvbRWbanSzde71
67pRe31xMsBa9LTKzW+BlkDZOddan7O6VhOLUFRBn4V2PdCcSM2mx3w3Fjw2
17rnibdAx+7tuusGXMb8FWalFo5c24GfjHcclqkdWu8DtlQIVqZ4ahp9SgNM
kiCGOECP1iWqpMXlutGX3Dd6znetIJ9VJkqRhJ5GX2EjpPUkRHMTLk0X2px3
JlF4WAcDOhCIPh9JCKMDbqWN5ktX0DfR1Bdnw11QL9H+m+yw4hVOKxsvsEHL
HX96g8zelVG1Lonwui6jrhtwNwc2wUmYBUxncwoZVLmtO7hFVJG/Mmmik15s
9VaayMo67MAXoI9RTB9UMgKXoCY9mXj9/Abot1XL2aXH3P/zveRFdPeIdDvw
MPFtqqKDpP8OzjwE6iMyXNLWhywi8l9Y2P26UqXCTnJGTwnVD7zuxR2/aQ9d
3VxLQetSBd0MTKlMFOGBycdqj2PcRjbmPHz7wNCD/wPkLB8JxnnP6o4ndrLP
hLiLnjOQNReR1ASojSm1QHZpavDa+CbjHin/QYaoTKIHnwwSJ/hpG+Tn73F5
KOvs+hxOEwF0b2Xwlx0p0KmHmNuMOCdU4XD0MVu08MfWZPrW1y3RxwQs5gTI
8w6e/+bvSrCXEZYqJvLUmextt7WF1fZT6tBitlP4iLpf0GCc274zMHmwTh7A
vTdUaXf3GmeuUSxuH9sV/f2fJUIkMe98r+Fdf4OHIU2eceJrSNpeYbnoMcnI
v9n8Z98gSpzNTsyxcxKwlEBa9jhZySnos3Tmpr70WcovFrgoloedm1/Qg3fz
c3sHaeCPoiMQcGKKCriU1VCILTJfB2lRe9Xj7BAxq+fhQimgRaS1wilu0z3j
wijeNkBSvmYCLX/POfWF0bIOVTps5XRD7Eh6zvcTp+mB420K9Gpieu+KusmL
ZBhKYXLFCgVRnhath13eual0j/bCJIMFRHEaPRbSJA79nMmu/4jLGbU+5stL
Jd7XxS21rF/Njq8jqqI+ggFXLMchz8UrahVfqNW0xJC03oUkLWqJk6cJh/ke
tPOnPTxTRPeYc0Zia14BgGHGfHpTOvgT0n5wWEfxj7sH3pE5tiM7fo5GIaz9
+8T4d9wVWLfm9TEPw1ggjk/hqappCg/UtCuDv/Ydx2gsVBPKHMntLiqJE9co
wRsfv0IwhN2uAzre2StAqA3XQjatD+FBOX8BWf6VaI0ybbLQ4JM9SpP1CKki
Nt5+PhTr83dokE1f7Fb827KKPebX0spE3QY534iz6BQtIvpOb+SiqbLIlUeZ
A++NcNbJRvA4lFA0+UZDmxVhxpuYCWVruNhELS42w+t3CW1rF5sUlb/8dd3s
CUSTeGdnH8P/gnK+aMbjSTQA4yv4H3hAxzBoY59eVMWRtVCwkf9N6FAvwaYu
9MQhhEU9/md0edO7Uv4K60VDiZoxawqncsNFqpcZXNIUUk6ohUDbzBnhwuhF
E6pEgBrHHav8/ReYwvsgWtudUm0kRwM3sKpjTrhdme3ilHk9NTMreza/yj6u
bOgeCZ6N9/fs/vv+MoJ3Uqk7SMNo3jE0c44mHa5ncL7nE5FekMRulMehzrHf
zZkLGnQGPe0CKAUsR2hUdoaG5oFEWGHSSkM9InO9K6TqLoyYSi1HUurKob5g
InWyQwX2tMVdLxWbZ2IhY+JX1XDhZSZFK5kG5/jvLg7cv45ZNtE68Bs4Nq+E
VtKn/+6UPC46zFcNR+0x4TZQPGJRlFpdcMQSA3qk+YnwwgWX1FfYtE//y8W7
Z0rYbROH3TXkONcG0YE1abH8W8anPvlPX1dgRcmgMVc1w2GS56XHWwISltc8
f64ZkhsKp5dKceYwB7UPz5DpZV1LxmHUeAiDTPObs2ac4umCedQ+8hB9vLQG
q/xkrCF7oTHze96fSsAQhvZbMEoeP5kXS9tiEbZhoMjxcWab7NX19GX+7Cee
/iUFqwdLE+ic+RIiKm25//W56Xg1I/tXbVp8dEMlsy3pqfzlrtJEi9vA08N3
EahMfZjYy7l9nf43mftOtCrUA77uTLoYXab9cAv6JRtt+Qo0HkPvyZubBemu
dMuvLdud4UVBRehOyLZmE6K0XMPVrAZEtwTZ91dmmMXdqEBJ6vKpqMzk3PHV
jBBFes2+Itf0mC3CETQnX9buAHdl4QOQSpY/pBdqupHZ5JzCrrOaIOsuUben
fPl2ItkYY2TIISne0AfvQplEQuO7ML890Hokh4YxPvgU3TLqHWMHTMmSmj8w
hJptwmDkzvmXlh1XYYKkFHEJ0lGETkV0mYdDeXZRlREPIfnTApboC3sErGNp
z5M0MW2+Dy60Nszo+ShvLSNr13b73KLDRcFcY1hLFa2wtx4wliX+h+32EjFS
rn4KEiHoqJNNxxnJ9gwJAyXHAktcRQ/CnAH2lKkEglfPr3JRNB/Sh+Op5jGP
tnyWoptkQaW1VpKgiPQM5tqBwn1izSJSSs67it3uaajWTU6q9tvl1FNVPYJA
IrWC40HssqCDRvREzLETo5Ov6gD2ZNH2Oi7faoI0BDBdH8U6NWa2iXEs1AZ2
UkuTGFh7NNTamlDO2YCUB85bTXZXnK5DcnQ/0kmXOte3XfQrPjNkxQNN3pHv
xIJ32c09LTqGIoHeX4vjs/LZW3n42oLnJ3WubYzHpTPUxMD9wen2KVrPIvnM
/+DwNQ0UT7DRbP2nYqfuTC5krq8F5L1AbottHcF7Y5B1atR5er2/5qAa71dY
uUMAofQtV6dpTAB7h4MqOhXrsZLv3of3Amsd/W6xCO+ri+U7lBLyzEt+Yv2t
PweD47X4RrbBLLFif9sh8xybJU/cBwDBhcUP7JJWQZ+xdc2w95fxjYGUUEcj
STRihp5yFzK4rSUxfJv0ZGScTYkBzoYWdtPbpd01ESu1OaeHpBUS+CAj4IsB
dazVoDZglrUIAtcBsQcMWzvL15jezh3Dw2tX4LNKG6fXTTSz2+T2r71+6+CV
DHEBdJg3Ex6hsxTkda2kseLqEhbiJVM1YqdsYOzkTO5SDCbLahpZOJ3yNY9r
exaXUXpj6bQ3s4bbHcSJmyiDtYd7N+q8gcDYrikQQdj3arY1pmTi7s7L3b4J
To03L+aqd5/g3rsYaizT0RNcafWIMhEM87aXpIfOwS/N05G2AHLwDv96lqa8
xbnvECrUBc7OD+vluDEFikvXaYP3288J8pw5TXPA3VJy6vCmgk0QImOi+SMZ
dj4MxfeueupElJbbZatdo7C9MChdyYkgeYiE0GbDytG0iWSBsP/XBSnHiVA/
PxgAwM0+dRqTm3lQkh/TyM7UzGZ7+JcHRph9aVa+vexfMVCF5GdPW8+9v5Br
4MQXH4N+QHCyJW0zrvH+E8us4sIe7SVIe/EVkvn4J+2c5KvL65mKDGNHOMWB
d5tmhAuKSBn4y9FAfQ/psRdEizbnv42JI71sCdibDL+LW98EVnEBqCLqd/Vh
Jy5+MDWlI6GmwfWtu14lgkTN/ocdHz+SjOgADuiMhRyYUHyezWylj8Rdj7qm
v2R2vNLrguHv7v6kx+BeG2QZpqKKjwAA6N/dAwWTntSKm509BVkJlJa6lHlR
ejACdNdTouT//kAUiF0pGPMDdVv9JiHVBFLRzOx0DivkvNFuj9Pd4AFlmdQA
NV6kc+3qzjrRe8B+KOs+YvmH/BD/jUZWI/1hUfy9m9IBzBptsRyrHWnqUF+S
iwLV+y766xQ6htVbLsBhmVhtemA5rSlww0Y0vNmzM4q/GIkk5h7z78DoxmsD
zZxYhhsHsZAzWibBrvOXmTJzqdgv+lgWd0QGNN/V7/Jt5BZTaiBRbVSQkHDJ
aj1+kCqMLmHVpNNAhzkKwM4ZuruydVZ/i+tOsDSQgCwUUG8M92lf1YwT9s0A
g+PxcAvrfcxJM/frwXs1kwDzBQE0vnRgmZR1OYuR8hYvH/iXfaC2EViQbQRL
fw6I4BsLZJr8DPrczMegkzRljoNQJtvhMFNtThpk+WCaV8qPvqXnlng6xWXO
45n3F+nYWVBX0zcH3TQwrln+doEvQ8rCDpqWMjpO/m/dBsR2jB5I+wgLXsOx
ugqJWWWpDyz/Qq9IpaNNw24HTCPMOX1Te5IT60ZV2DS4uQsf+/HDmjJaX7ax
PMRromnHPV6NKCXD1zVHn0H8x0Z2iFOJ0rfOl9Lh0pd4ktoA5Ic4y776Kyox
wjT3ZCYhLPamS0668qw87eTWgdHCMc4psq1Gxqy+W1l/n/tsSNh6acOhdByo
tiCUCn8jsxt+GNq1DrCa2aYWLmQjgb3lbmJBbDY2wMzEqwV5Cp2Hza8w7mqN
bB8vbbUgxfe5VA69etP03a6GQlIIvu6MtwgsHjz7FAQWTAIWYGp1t0t8R+mN
W5YrJ2nqVT8aqSVJN2pryclXb4fGgxdTNDbKJdJJ6pV52JTR4xzdI2n5ku08
MaoNX3xUTr+4FB50ur08aXbuuoEuevGlb8jgghuJHwXIZmtyuLfnZ07GD9pM
5jOrtv/EsKJftfuG9MI5vXy8oJ5pdj+7YICrC9LUzc5+4+ROjpr3g+USbITh
8J3eccOgdBVO4o7ZzCouEio3LA+w5WToIERd6qimSzMJ1AqEeFxT5vYWOmRT
iDQHxhKGrf2DbQ+G+qxfMxTH+e2fLjkcwyDxSsxqsVRg+5cJyuWPNQS5NGQd
b6jvXdEaSzJvkEoQjHJ/DQWJMQMb+u+jL2bjBHhvB7jOtuZ0RdAuKmXnTm2u
IjIgQd9WYS/krkyv8u1x2KgCPmAKfM8cKuRitpWwbte7ozy43GW3bSd8viFj
sxeHu5wNkR8ZW8qKWfEuhuzmhg3C7jCS4KM549hfTIlhaAla7i2rShUrklYw
+8voO9trHVeOiJ8LEPVDv+lJUhvLnOSAlep24IY5cYDQqeAdOZZr1md/RItQ
BAzpAN3cotkcXxptQU89M6Cs85iVKchvd3oNag/mczpZ3Wr8+SshTLF9GHHH
4dP/KNdQc2n2QfEISK4NP7F0ozlIVsM2f+XZWH55pjCBPIT2Ac6fIN5SvDH0
u2m/+zIej2s+v9Y9Lp1lzuo+FomNOwJ/FIbEybLLxFDRkqqfyZkr/FeQF250
kvqZzepaaslYMEXBS7jpJwFm12OdxVbFW0x/rBSoeLAbTnBt0d99KFbxi0yh
eqAFcwAa9qkYSvApfnJPwOpFZTWBkCLWmFDFmi/nmfHA8ZIVvYANIyIlCHr+
krMCFTVShRT4vVByOxWrX5kOmNxc4zjKVZxLdvhNqmLEpn00owcWejh5fk4J
IBQDF9LJk9tNIcpxbiAz9k4zoVm7SA2j7fSbt9oay/1as9+rSPxHzC2LfxN0
3/TnqTey2bckY60bslas/2ygLvPbRy3bevBLwrmA57yWMe6bK2qUKxAMWfiS
1vN3cQuLFBRoMchn7WuwhW50SNi443LBorpBXdVGu3VRFICREfKjz6KvGU+Q
YjZobjaV+YFB219R7I55PfByKWT5BzziCoXBMr4xfxIGeVJJsePJ7Qhb6FAC
zb+tXKC2tl7P+ktr+rZR/h2+SDzQIpupxPAsuFFARzcDXUANkm+YYh/iNsUn
gP17YkwlLKZa4iX4KyfYW1AA9aeuLNtTrlllGUeYsGdEGn9xDf2Gh1C2LV8j
Vxu3e+L1VFDe+Dt5Ix+Jy1N95DzFfSSQH7Y+hAb/UpJURsVYfsZOhRWkxqbq
ky6qWrE0t18+S8zIYy6pM8WZas0LFkoCRKt4JnGEQAn9LncoJCgFAz/B6kpS
rKN380sw3kxpwxGosmnUPST28UtEyAuUwNJKUQIx1CtjCBNKgOsJuOicl0Vl
jnKs9tO6DHExaEs4lnjMJrnz6UlifJ7EwRq0srCc8gSfbNWeZV0NlTCOxV7i
1n+NfuSqC1OKoiHYb2Tl2uG6TxANRPpGSuyi5MZad/IuGW+vKVrvGwh8Ubwr
BR0f7HSjA+bVlY8jh7yICO/GPTFeA3IGV/RDZoOMAZ6+aALpnRIufNtLQA7K
zGUZiFROTi6VySDz2gGphw16bbFsaGOjMN43i/n6W+2pXBWSem/rlYgxEpGI
Yz3ye1FuSrcVjyzpPvKxhZ23y0i9L7yrXRAx95zajvlA18DpKlkOO4RbY7cX
unV0UVBvxs6mIDXdYSgdUX47TMfwRNeVzVLbVBeKuwsH6zzLA6upbmzFs0bl
0OJCS19gtVbmmB91/WMRXc0IvkEKNbaoSB0WRj6Qu86m6EIpAiZu9hbu9DPb
alzM+tgaflOxrtZbJ/yqI9bSoHc8Z/O6gE6ywt6ThUfEkiIWVxsWL8WGWhHN
LfEXaqJctF4pUoV9CMy0bhN6+EAWVqXcVi6o0wAjvUVI2l45wnFFd6zbcfPD
t3cJCFSA+RgPoXaq8c1iZtJYzh71JGRxTRU4Kx6TCghV8lTSdllqVbDZxyK7
kgtXFdBITnZhBSWJIfiRdMxgiatAVEAnFJ1yZahNM49aY2HdWZ0yLUHIm2rD
9LG22JULo76pQSI3HbXJ5dNmh1FCeyzmc9L9/bkiIHe/7Ew9vYLvjCObEM9/
GI3KyF/eiO/qiMgYTpODref6StmEgo9IjyjJ8UoKgj0Z0THCGCRpgy/IAxHd
Pmva7DtjwvhAWg6Nii0bgNR07gYDwNKJJuv5AlYoa06xb9gjiuILHXvDl5NV
1WBeA5DYj2h4kkR8zXcoYv4jQF3aiopP3q60eH9KwVWwY14+W+Hy9F8WLYBV
ol0BtPwD9lcSErP4SR2LxmKmgfqFFX8YWy2sUtK5sk6mRv3zuV+bcqjk2YJS
8GO+hT/Ghla/Tb+LibALbysZKFiuXcvjYtBJftHZoXaKB6ynHUemXJ4jFAUD
7lw4UpJABCACh603rMeqFvX/2YXoRQcDb57bPf1a8BVnKJDkLwWRph8y5pPy
0gK4d7gYMy32M5iaccxJU4+wyftqXyEBCeaHJqEE3jEG+h1dBdIX+katMLWS
meTcK+hfMzjecj3rnKyJfUnJTLsBOFY3TqILVpn9ib1uXousv7MnW/ua2wuq
RSnGsSG1eGl4to7+1RxTRQSCdC0wGESZ+8NvrSXdaWcV8M4gkonhRPjhmhGY
IUcwS2zRaALyqQ0Q0VEGC3lqHBltHNeEx8HLgHIwKbLhp24I8RcNRuLfK+xK
twpjdcpPf2L+ECynKRoZCu3pEIQcDLKMtM64EilyERovmCj3Hn5Z817bnh9K
V/d+XgODXZqZEKGBAaDFHCXw+jOU33wqWdgpUnXCtoXtP9+nw3ibdZpBrnfl
kZmraKZOtwklqb1JYbupWzPknRbaUgCt5ddCkPjITrTdIs9IdVzbX+KlZ9Sd
GyXyKJCLN5F4IychdnH28zrvy8QbaU/A6LLx6EaL3DdRcRcSI+KiJXMj/P0r
n1iF2+eyeAeF/fwDqW0iIRM3AC5t+S1UT7C19VAoQvQeK23/2LyvX3n9AEc+
c177wLycRuefHAC62XF24oQ8diHbXdsNalhCUplpl4pqvrXT92alH77Xis01
Jn+QiiB+yednFlvWInJ6XGNM45K1Amsj/CEAEYKoljevjozi77UdAFrOHS6u
pG/efN/IRI9cTmvXLARvuKYdcNwES9ZDB6kv5UDiV7tluaLmDKTqNqcvFWaH
TbUD0zfPRuZBsSNNhkA79FIl9sxf/KfAJvw1sQK5nYxoeLwDN/8iTRMkcc5w
Z94yT56UaY4768XmwGDDpCgDxfcbJ6m79VqWdoRtlfmsP9WfoMOC1S3l+ydU
5++mD7rtODMCiQ8sYphC9F2BO6FdOh3qLt7zlyEX9/NFAoQkLgJrg1z3q/vg
EGw4SxlOlawnyddiVxhUh45kwrQcVE/L61ZxacfQiN9FpkcPgBq+GuOBrn5S
gY7yh2+QYoY5M5mphv68zlqWcfAxKboVvQryAIO6kDXnT3UgfbDoVxfbGC+K
o/hZkEgy5QH8F1AweQOA2jskkN0iJofRevJuC0ZvEn5W/YBdqTU4zxh2B0qn
/CuA3TUaMIIFYw/x4Spx1jzFRv41fWwkO5RjzVaPYlSfhbvTjrOCzH2wpqC0
1wwzW74tDFDkB+Fulj56J5BCGRq/eS4MqfaH1H83ClGK/31v1Cs48Wg1S2Qp
rd8WRk5FXoucqfY2ALU+oGQ5/7Uct9NpOLPZ4hlWCSZHcDw4PJNVyHnLdlQY
Z6oR8Fu9VM5a70ooketQQSo4Zxpl1cu0HTQ8lb3r8nz1ySWyf+cI5B7md+V4
PBI1emr93FaiVasGLrSpsVJswz5neySsUSiMUZ1WnXpf1X4k0roAQxS+U+BE
kAOw1yzOc17FXueGRhC9CmiDgGWK9lWY/bGWFTKTbUbnF+ubQcJusbQjMis5
W2+IOZ20cC24kb9zVLQ2pB9JU6HLaExisMMjN0PmJ0L8Eog1sBr7A/VBRzCm
FMcU7APDms2uS9uVBPXB2d/zVDoAq3qrUVEt2HSlpVvLlOa0jxwuPAqW7IjM
8kTaYdMYVyWS6lV2tOpE/hE4mfodJpv0c6QfQJlHsRBUPw/9rfkhh8v/uLRw
0xnY8yKXcpbpqK7PchtaQ//YHGuSt85PW7g63RQpZLw3TELwNyzjBJ9U34rm
pazCFw8QfG0n+xUIDY+py/0VyYyrCG1RLF1MyFecIquHYsQWrp6wH/d5iZoh
jdFm3wzZE4cRpKoSN405zHZoRIfvbDbNGtQAuVtugDc5X+d2CwYmoH2UitxO
6pubn8DxFW/GMBpJ4yj07WPP+1L2/iLafihgukR3nPl6xEctdT+Q6YAkLRxJ
+sz/s/sPCy4au5B1JPNoTClcfU0qMR/ElmtRdHFrhQ7E+8sOyvGmKvnjcm08
DhOpqulwHcYQDTAPG2d/1tK3W7rnR8oA5QJd26HlTThk1b6iflPZsMgeZDpe
E2Un5LDOzlOpKE4ObrzNikhHd4hrPvG8HqzaQzaZ+IsUaei5qrCGk2JrNMIn
a44ooIjVam4yoKAtTGBuTfnuB67HzGEUZj71j43w8zrF5dD2prc6g872a+3s
Gn5B4RXpm0ujGYuZOwsUEri98Wxzj6LeAcp+lhudHy+z0i/JObB0bc64b3q1
zPr7YlJ5qB8vQci+dnlZlhqZb/D+cBDI8/xH5f+ggsgoC5NcdK/oS85YvpB/
BAneUtixPvOA7qmwtkpRLUL39HwKfAkDmj47PGSeklr3UMlm5WxXEBBT5srN
WimvZmmQgjbxLYOW5c4dR/zEaL+lwq0tWoKJvO6AUYso+TPjzcGcrCK+P6aI
fksilv0BJ5b2rPNAXdbwP5U9aTMFCPwxXoWsLnlsZFU1DRMRmX9bsanNAIiJ
uQ6dH2hskxSOAFbqAZF9JfCJ1zbKSunypkZaRNz8UEA+tp2u/f+Kwb6Yf2+S
w35T2pz0H8Lzfil65BBAKHgM/fg86aArnWKIwAGJzfluZ9a5LhYtzRHSdLxR
WOBj8/ObnDwbJRP0UnfssUliwpIdgPfRhd0WNMxuZWbQgGzdHxGjjbBM6OCf
bYtyeDuqABcnxZHq0YDh5HBKzy87UrRCtXkISIsLfXUlmFrXhtXbfEiuSaeq
3qxHCjYrAciPcdJSvFawC7ddgPV2H7EZenNCEKR3Cb7/AehZvZyG/iRQhFvq
Ylb/PT5824VERs8QiaK2k4q33LKOhpTUqum9jwkD+aoZv9h4Y3G1ZBcAxvdG
XUiSNAE9Fq53aPAcjdpC0ePb+yQcWk16lGzSh0pmxEGmvEsWpR27KPfPTxMH
74VxUkEM3ZhDgzqlWynvCCRBTXLWNTN2FCU9dkhUQLodGtYpCmllvKYYtcR0
CDnzgtE4wxgnEIkMk2S1yKVDIuIf5dnndqnplSJo7EW55BDvTCD5GA9B4ank
wCERXbOKqSRWqqSNbsjW2TKsxrD1kwz8cWTYXK9xsqZSOCaqkySi/X29HbTv
PF835y3AK/u2ab6LnqshwFfImm1Xi9UGSoMWNnAy1wcdLE9YR6VqFmpULiXW
mcr2lQOZXvLJ37wWJ58HgT8eb4TRcLb6hKJ9r4qQi/Q18M4qL/a/MeE7gG5a
qoaiZoLtUDIsozJ1nkOeSlUy2giYGpECjHgHYed9xXNd/1z9aCBQuHa11fZH
Tvoe5r/jFUI3qHg2yOaqbyLjBryVFcEnf21dQpu2iWLIfWZIsQGledDmeQUT
Y/gPq0qA4WV8w3atFw4UiyVzs5Ks12vkN+64OIoHSclsf3/P+vrCXA0Fnrp6
Z3LH4LjeiKEqrBg3NltmDcVcZ2rKFYgzcrj+M5ZPeGZ4SdNHKOg3pKU+Emi6
MJQuINQI/8rnws1K8SKMXOAUUEISWctLDnRdN2l06XetNTSHk75FbwJKhe+j
NcOg5RjXW+Su4xOJVoBsbHKenUFzn4OpPYJyHQMP8/dvdPViZ37r3UAbbI/+
7IWTLcrrBZlS+jVE910RwrqjomAU569Yayh1xGgDhY1rNwdliZ0vhuIFCiob
zi8a6tYMLVh3hjt5zEGer1Hes2nEAYhfxzTlF5zg7erQwfDvdYePUV11TIsg
p8Bmg2MBY5SrgImcvEo5HRep9f/SFierlxhqbW7OE0d0De9QIZcHeGMA/1Fx
CMFGV3gGpXFo0NAuRKhCOwuebb6lZBmJj6rLeSSgxY8lHpM3P5XqhJUGs3DR
h/nYPShc3UNMAHh5bliTWsBUtyu3AScqAuDO0e2NSHnyWzDOqk/KX4tChMax
jDKM0pFrf+r0IXRK4RiHTqvZ0AIlAxRGAe3oLIR/tDGTQAAvuPW5PaopS0Bg
NRzCX/6Ogy1PDbnbwysj5HBEzXTf1vppaEO5Hlv2Vdshb0QNDNzhi1dT2ECd
2St/zzR1GQJCsZTX9bFFiSE7b0b+g4VraOY5K7idz0EI8GSMMtkFAAF6UjF1
2NY9cqdoJmR+eMpLMN9nevfsn1+rh8G1zyzUbKYdWTpF8YC1l9ahMpuUeY80
E1bxsM0WfraIcrjfJCZ+a8IXUnPADRHNsGwz7dRAdKVcr9JjS3MB358IPoUI
A2zSV+uuy2z2Ite4wMnKiy/BnrRdOaP2qxjPCB3axQ8GsVQjyGpmwXVrIqdq
/o8HChU47K/kWfg7E2HoV/HBm915wEV3LPnPFp1DcBThpmqcnPQUdKzr/HMZ
Vc6DL4fXKeVpth1UuJQHiq07NCAHRWNiDMY8YbPIAtj/WMwf2dPoA8LnSIbl
o/jWaWKiG3A1nTC0b33zfX7P6ETVtNQzUcsQ/Ljsrjxq3cbvYU2qHOuclAf7
CKdm8fcpUkdjHQPUmMIvQal5nLxJ+14x9ro/Xw2Qpj7UrJhSYPDJIojV24Ya
zVwfZ9nho93kC+riE9lW8dxJ/LQwFIXnB+Ytx5E3J4MSTZgyrXxhPLzAyuyD
7+gLFjr3B00VMjX/nENpEPcR4MPdVeIv1IVFI4IF2DsmaT2RGxeLwTHnDEjq
uonjU2sF6oNUpulhGlvWsYBH4D06addb4TFbjsMRgY/s20NGD8ZJWvDCBAad
KVr0z3gM6qt4An7BmgjnzkcU/7KbZDl1ctnsDHO/ekPB9xcN8d5/z+7fLUn2
bWBtr4k7OGEZ7sh+8ENUvPAJ0jCljuHkDV5qaZ309DH/hmZ8ixm5NP4GkJBF
/XWk69uqsKnt0LfzURlvet7bLYlSx8ZmcFzv2zGPHgSJwOe0X9/9JmzQwR3N
gDITyhqw5Km06usGLiJ93Li5dcQOBKoK/bHLp20/ilWaCMU3gzH8jo1CipEP
F/MBPGczpyB8jAOt1eUjdAW5eUk0J7gLxgdUauIWfoi2cgxQ41BXIPnIsCcx
9weI5tY7ZPg2kD6FmkloGLr6RK5kA96FPjifi+8OWwtYYc0vkqg2/04sB608
2V3BhX49HR2ului51qxYb+TE9WTks44ErQfwi+ImSXVO8YGm63MJbjJh1ipG
9PB+YUT3s+FrP4qfMW1o0k84JO990OGK8WMIICV/qOM1WbTQGut7JoAphfrA
+miAld56Gc5dgwzmHbDcQkf7s0t1SMPomTgMjwE17Fdl8qy7tKlbDMIkQ8hE
1FSLyD6mpDHyeD3JpMNJQkQlzY+pNRpzHCaHoJlrgiAqJB6Zb7lifQvZO9RO
GfKhEEtDJyr0cJ+aR1HVJoImnXrSrMTOWT0H6NBbjCcFSJ96jNaz958aJyk4
SzZAUaOUrMemOvFRkiERLmVI8C8c3jqeN32KdFJvJfV6sUA++vxWSFaUOnxO
rEMwUqZJN2YoGdlGydJkyBKtTVVVxHUeYKn/tSCpgRGJFBxyBSiW0KIluubO
Sbec+sA+K7Qilgfn1REEvIFfkEcb73opNr3AUPZ2lYeULpKWRlLfw4OZkSNl
8lez/Am8WWqCkwT5nUBecVNQi9Fkap5W5bg8vh7WOgKD5i5ba7/618Uru5wQ
yEuGgJNPwR/P+DA3rEJ/Kf94X0iqLu3DUC3AmGVJ4aMuz2PtclyueQVKLrpU
v1GhkDvCdhR6SOFDdK1AWRZHap0aoGXB/buWFxbVD01CZVUgDMfSsxvqG7k4
hkuZ1kTyhgzXIR9jOYKRz6HNqQbIZEXf1Ykcl77J1Pv9Rl0QpyLdBgTxZqe8
+h5NA6DFzqMHqvq9HQbpcDO692sEiAoml6oUxB3/Oys1E7ywJmf26K5Ifejv
lCT6wsJhN+5+ywj9633nSCMXEPBvKh06f1cNnmCXX+A0tryefXQN4d4D2EX7
ZYEHxHbVVHRUOh5yJk3Da5q/x87KUzRKMD11QHUWOOqnqAfN9gff0jNGF12R
q9+8sMSBfWKpdT+FG8NxQAuxag+4h7k3QHX4Yez4yGnSfrnNMLeQaaMQdkst
7Tm2CXtxk7Z7QegwBOLEZz/OKdzL5+/+NP0orvJeyV7NTdxLVYwi+vJB3qdG
L9NufVBCiL+E8ZSW15JCfqOHytjpYZPYJFqSwDxQTFMzbhFpi2U7MREo6WBj
hpm7ag5TF1Dur0DNviij0UTsq0zIG/uoJD4FDPEXwUFMmMCZklbZ4u0Z3Vjl
7QaLJiFJnCz7yGpd5wCiP87og/4Ik7RVqHpp7EagPOzFwGzNz/wZi4mow9Ce
MrtvNX22BbESa/GHDGTA2o64cWGyJ/4eaIKBBOciLSLDb8HmsWypoMiIqYws
G1E4HIPQzXajsYshc9nfBGUO9zLyCBiKzA1GorLVFFIpnP7C6GADZ2HeA/XR
FNVMGvWEyrhtiMlLiFKGuqHWz+uy+4Y/z7iueLu70i5x/+yDe+vdbCdodciT
g3H37B4u8WgRPrnmWj8Td5GTF+VsajDorcBVQ5pZbyqPB/tS4XD7RQFnAsAg
/QvoNJW2n/GjlTFFDkFO/vtyvdbkTtM40y/d9hEd3hTbDiYK0hjLntRO36IE
K8OoDf3Rz5Tzgty9PA4Od4rk0i7pXQ8TOG2JRP8C3zYBCgCuh0iCdEB01MnE
nCvtStpIPanZ4T3od6iu+enSEkYp6AjK4U+MZ+HZOhcTwsVS87+Pp2s2mQeu
gzpLQnERiIck7YKZcWHXIsxRcmHlDsySH0kgW3+SdZFb+KoztNdxcqh0SIRo
269dpw+BuaBRJcGTrRtQ39FzmdZiRYiKXk3Uo8mtowrc3JQObsHIRhWMbwhe
t3ruMlkRunAkAULZj/ayefp8ckQNczhLVqkPHMcgRY6ZuJXp2MBU5T+jxIjf
wJjXM5bIiCvo9pl2P/K5M19XqxiffJ7Xs2hn/JOFAcBRKf7AF9428khnHnQT
nHnlnIYEpm51g8nfXKyWnC4wvwNfy7E7Faw9rEnL1Z9dCPvdEIUiJW1MDIWl
rNxNqzs9I2gdY2qqYPIANvMp0Cl5htY11n5NSjusxiXNoK1KBOjHMKTcm7hd
Z2P4OEvgdK4x6QBAeoftIAzRV05/S8mh6Ijo9By4w/aaMvV4yzPON1YTgHQV
qF4qAeVdUVolVNwb0+miTtU1XdJVnXsGCCl8XvPegge/LIslhKK53cQUy5C6
B5/ZlUyZKDtncFI3SWrbpjjPsBtJQ094SypJC5LWmKQWPwQRc3NPBxxth5ol
tX6UNpW+iyYdnbkrPnjzo1Lt76COU7zeoAfeNfp40a/nXRT2nJ13+S6YeOfv
mHbcC+nun26AgOSbOI+4y1kEvr0OmOonbdRZK0tzgUs7WJ8mS6YWN2k2Jfcc
juLtJ85dtOiRfjDm/WhcZLWcpZmJ/YYNBWBEkq58M9NdIw/WODOMcp7SrxsS
zEX/3L7q9PWuLpQMvKSFHyJ9nC3aVDsXApP+Kut6SgccKF/diVQ+z8EMtr5M
JhpkR06CxHLw29Yckbblff1mVvVBaAPPEjlyffQfAgTQBkZqUZ4Jn5y+tC4t
BYGK0TXi1cf0y4agbOE+GkUy3QbM1ie6Su4OiWMlX2wWd+zT/RCKUZ/QmkCV
G23Ne/2Gh7tIW5kPaUAiGfufQa+ssSV/RWDUHogrW7qhAY+HdILILeMB8/6h
1l/vMtrw5FTsoYaRIS/4KL/78FNOzjekNv54zeL8s+Y3Eoxlo9mfxDOQ4VXC
1OenU7fZ9o/OWaUkOlwCcYIBoqZYdMHqo7Gxiq9eW9706cvcKzIFjVaM4jQ6
Y6UOM8ppVlCKhnNcluWTWN3zY6geEshzjNegHXs/5Ll+xlN8hYahRQKy0ohz
ygtLfzV6HI2ke1rIjHUdD2HBZBESwR5cCnNE8cfowgxGuGKMvlmFNVypHkqb
F56HrQchagDQeN1f0vXXs0OSeY9nS6pgWiC98GmIOWwdgvJ1ccc3AcCZiw6J
0/9DNDWU44FFHw/EWcYTLUtzvlt2A1b//wisQZ1/hV7yOAdrt6fSTQ8ATZ6I
2PT9BdpKQTC2ncXlm9rpDsivwgc+50JfCVKfn5jrxWp+ektcbvEPhI3DfCsg
W2cxLIhG3tb+2I4f65vdKnJydPAGKESy77CuYEUbVe5G9ti1kc96Lwzn2ZVe
P0D8LpregWA2NTGZPSFdCR5tzD4AUpEokK5x6Uff//OIzH0HRmnI5WJi3/UY
UQtcprX1v15acgbtYaaBPS++TqL5KNyaouqhTYpLiAK80DqrVOma5ciQGj2f
h22wYuObOeTlduVZjB3yjcxYrkeLdYIcooJfvTUKajJHNzs1/nqgaKytLwaR
Px6iDpimk/zDeJl4KuZGaWoA+N6b7fskeyxKTHtY/lQ2XnjadwRB9TIyKKq1
V2GjIXp/hG0FbrK6muYIjR56RjDspDtdgtDheuEVLwSKLctEFIZBAB2MEP+i
Pb3sL2079SoutaWCBpJtJUz5FUjj9H7w3aHu9GLLGHfuNtm/2QDM7vP9n/cj
v3oH9Uj+34uVw+uJNBksx5n41LgE89+uQdM97FocIvMEqD7G1/TKPjFAFjKE
4bNLqLWhfVoUAzIto60GZbiWUOho5Q0YUR0g8OSZAX0gGzT1SAdeNfARw49g
Eg8FN/3587O0svUNXLj9AHfg2U9AiUjJN9bpABWH+QYSROiy7giHQ3Xyjwbl
yD0VntvSN8aRHq7bEQEPwewHyhJ349g+Vcjn97nCXMWypfd5MgadzpKqFcXf
hB8gddChgQ/lYkXXYvSzkXwO+SIRIXgJGuAsuWEr95ycwWbvfMKD81qlh3hV
Ukt0IZxujLtdL1XPt3KiQOYjLGlvgoDJpB4QIEZwXN2AvrocfiULDuSmaFst
8f2fngbviXLhfEMX0G2H8HSrLqoBVcqCf0R9R2Xz0zIDX9juc/OvVC3OoS/B
Ul7qyPwYwiO69Yoli2vjSyfw8Kt3j9nXpy0ghCQORUKyFF31wbUxzl7g6+iH
1lhNM4ehHMwM02u8PN9+yFDYyDfvbiNeTZr3/n9lcV6o5kFJSDV7XZNCCejv
araTTaFaXZqAjsJ9GKy0PnPmbd+jGF4xj9+ISuJg9AxqcpueXmdaRgnON9tA
k4y3rhp+Mw8aWCg3xromiiVoAC9YbnicmnM2UmqKqt594FvYrYmHz4E33B1j
aTt0ai4WHooKFvaWiGkiXXmXW822r5DPbcT1BnGqaQu7l4BfIpHXmnX4MSPJ
P0nGOyB4HddwEzEdtxwHe7DKep0PQpUhObO6roA1hrNHmE8Mv12NZvtvuYc6
gLuPafdL5xGBFOKJmorBoENoOFF/xvMuJES516buGMyR4hxT8JDlfmMT3iCc
0NwGaabESFGvcFVeyuuECFj2Tg9mMYUq+QPaE6sQ6Yz6RqkeUUGvFCeMHghY
DXpzwbFu33F7vfGxiV6GdfjA/DpVL0AkigS+DFHsStR1vHVEf7BwKn013TKI
xXb1cRftFEYuFRR9WfV3idioSN1ls9umLBQD/cFiEasYAGPaVhlUhE+NU8Gy
ZTGoOaoiuRrETo64lP7A7B07xdyqE80p4jo3rOiY558WEiHQDvTgeigzuVHL
J303bxSEfl8YoCuuhmCDG8QKkNGZh0kO/pwyWJjHCkT+xf7Gvuj4hE5Y6EKc
j1HpcnQv6Q8KzMzW86t+bleeWDCpfJmWzJVAlQiwVaEkRhYeSUrW6W1H12bC
Oe7HTsbExI61V7T8Mk6swPX96z6X2iiSovDOh8xuGOF9Ek9NPrVCnbj7QLjh
oVPegO54pkPBWBuV1YgaqyR7Fc+tpOGPhwc93jMyPsm10ZxjHN1ZXE4sB2Ub
tTql8G9qxaiEVJbGonlYXf1aDEjeQsBkqpOSFAz9+AgnPi2fnSJ8HbQIRAhf
9mIRWHrgHFRw+K900wDKa9sdQc4awN8UaQO7VT8jyzRdKWrY8rdlZ/wMOn9h
qBfupAE+xnuEsl/QABD9+9yUJ/z8+EfszTvJ91AB7Iz/Vbfufr84+xIylYjm
u9fBmuV8cAfZ8VFVVZk0+WICKEpSWQovm1Gj+OQBGjn3mwJ+yxxfJJT5bxkE
/TwxAgPP47uRFHSV7Tr9EGv3yWam4GfaUqef+/emGTzIhbjjwmHFaF6pF/cw
mbDESawLKpea2XBhw4FkuJVPwIjfTGYcmhjNgTIFLxeyavb1/U3d4AmWiRVu
duwx3sz9KJUudzPh/ALufL0ZeQwxrbA2q0ALKIyOK4S2UwnhfQOtv1sYVcEK
vsYQEaoB8ldFq7tfdQkCg5y7LgjRF9S5Yj1Owkn7HRZuwhIfMQkwHu93BsuS
rASCZqJ/SZLQEySevfpt+o92HfF5yOJAe3CYsJC3JaY0IUoQ0lTfMR7FDHpR
C5MfSuJiW0+fBKd88Sflq5pqQ6Ki2ptTqNdJMz463QCRZMRQpOayw5IuF0oc
kWdeBEMp3hoQ33DXpDYMnlLI6jMRiwWEkPaoswpUcfjpyubOlQIiqYLkwz7R
hOaHKPpVTSCrQ6DGc1zQ2hw25lx6vRfyBLAXahcjSkfX4D+pFRg9Vele7IUG
3HC8X1qnOHyUx+KILTmoKPnvm1dcBE4a5cMga0VVhuSVZEdC8h0qSdCFF6SX
e1/QnPGndiJlpRbk7dEVdPYlJw8hXHnQujN5IroPqDZrQ82ZOLqfTr3s3yUq
rkJlpz85PDcvVt0tBjUS2jbB0ovibkMu/Y7XWby1hBquJpSSH26IEOo0vkNo
w2YUPD2bU7KtZ0nEQavUxdZdh1BDV8ySPgJzho720T9/ptClahCJVfqLeQ+8
Myzn6M5Oeyo8GQB6fl5qgBcZdtiJU7d/5YOe5nxfePeygqlWoDhUfKn4igPA
BhrZcmti/+lCr/w6RONpdS+r949Nqtug54tDcAoqthgXg1U06d2HYuf0lk3m
3PXovdVI/piLqzuzEPJpYadGwEUWPPtHhAraf3MjSkI5XZyfoMDZJnhjneuN
sfB031JnncFvU+0m6LSV9Rg7pn+eXodtOt0qMH25FUea/i3i9il1+X2WTpeN
2G8NdlsmQv68ar43HRLLcmTN5hvucxSvzMmpEu9nfM4fai9ZQUJ2Q9pwjatw
Js/j1PCGckl1kLYabUlWa5BV+FhhmGOS5c7TkT+I7d3V4j/PNIfAt4r6WqlH
k4SrwWut6TMztyREfc98Fg8GsXcJ6Gwk303nG/EyOkttV3tByX0pi79sG5OV
jb1PpdlsAS/UhtUST8o7af6CFK1Jsy1O5qZZr//VPsAr7+ym+5t+5yPdzeG3
2eFSf3CVnSk776N2ve9ycsCjMLCVhpFm8o/F0JiNU87KmgaqRXjRgrfB1z0q
e6odBMVuKOMbT3Blkg+4wYv8Lqvpoabwb4iygig95cEG4DZCnG+0N7C7DymP
zi/ywTGjzZgAjcMMPCHQTgmVl3NhZUaSsXx8/OCDiIdYRmdAPi8UabVwEmZ/
3wGnR5PvdmtrNL768DLpemrS9O4yx4sLj0Ew1BXFaOZvY9UhJAzdGbxDCz0j
62nrYe53nFaWbE7HxDntaBPxRG7C46YvBWfOfX04JNzdOi5OnROXjnnwMK6Y
vxWLzIygZBf7kW2Xb9wkrzD631O4sKHYAV+sU4tJnkNg1gxwpTm6okjcOUPP
6UEpecLCJSgjD0ZolGK4jeKc9i+S1SoB94PbMXA/+2/2t6W6HRSOA97eWqbG
+1NuB8hecUNis63+T5NhBj9u0G8ZkFZYFXYhBDmTZcTaMW9Y7io5LOILJ0FY
bDLQ6VssY1pPHT0NxA8qVJJgznnxsOwR7K6To9RDCxgJFpgIX/lP4zv+G21J
AkIc1JDwcv96Lsoak4XUZbFhpu8rSPWXm0LKvVtEQFZwimZsAEnGxvTYbqD2
I81vk430mm7YhN+kZUPksOXyfw/tRRNmvmc7m9l+dLM5ZL5CplfM2qoYcJSH
jUJ3mYIX4yVYpTgsO45uCS/hMty8dqJ9xhlCsZ1pnaeM9h5OC1BD0EuVib+u
jIo2sRctjrhg9MvVSArVjHvB+ghgiD1mDytLzdMdtBuHL2r8lOgccW/QlNdE
d6J/18W90qS+4URHug3Bv0zekoe4/m5NNaw7hSHM7ZekTQfcbgFwPuLkz5VD
NHAKOyv8iPuBjyDuMYzxjTfAwLZ97396TQ1zBR3YMmH6GjwbJUC5ByS6Ic/v
QM3TS4qndNyuP2VOftcZmQrM2SUeS+kqz1RR0XNVuZI9QQbzF6eGxGKNZoH+
7LUwt3jeo/D9oH3tf1GDrJdIwsSNNcPv8d1LWqJQYeE0se1u/u13FIAom6E4
wEK1kEqwe6J3lM31pHggAahVD27RZAbAqEsdnPY0Ng6qf3Xoa7SC5T5+e3+u
2jRQ2cI9VymogGCm4UsIPMz22XkPMSR9sUWVdPL8SBZ8SM2HrCaDfpHmR76n
dlfA7gULHbVtvR8u/cNOr0Db8x1OEMBwOf4U16p8zPdNRBtp9K2H7Wjy2xqX
aG0qNc9CUs3YKySXDJgPRKElgIyoIyK1Mb5WT71Q4qxl6UZMGqPE4nFICNKp
qetVzzx+GDNztdMaUssHMCyMhNUZH4Xq7qrL3Bb8eSWmwUSq8m2+BVrzaNTt
DhV+nRC9/sf3lfMbaojZXtQRV3f4XaKd9zyGN2W0npuXb+qbAz80dAVGRWxu
OY5bYQiDPrWPpMgfW9nrDqkE2QabcU+rAtzXPXk3MN//sX/N5eyUOYXe6L2E
xWu8qLmhacQo2Vf3Us1DXpknxHMslOYFwVHYc1RAOK0JBlV+hoYzHyT3K0rm
cyT3Flvnv2rWcJmXuL8kqWxL1+LdFsLGpi1DTkvxrIbjaLBizEn7zBChP2si
J4E+PhRz07Bp/mp68WrFaGcB1VTJexTl/b8XKx0UgC+F6wSw+rHoLi3D+YCn
KrULZedpvC1FJm7WXmH42rkexKDqQSkdixDaMblW7cF56pwCKTUyqnENL32g
GA9NkzHqc1x4oimzt0fBMF23XdysZxl0pSVpD/mGmzU1MkGR1cciMOoY3U1S
lSfqRNRCYxJdShYjX3mLKFEgZVhH9gl10KoUUgVz4QdCgktXq1I0W/Kj/FGG
28g/iZC2XnZf48A3Fxg7ZFHmDvWdHYMJsltn7WS1fjyiF6j5+o1iGnTwasoj
BKxzKpawUo/jFeNyGxDYjw6339pHzPJ8aC636mY2OafLeQO8O8B8UVxKuTk+
G0Y6D530mdUpSZdziyU5JW1g9UUt1oUgPbazyMunKTBhE1IZWM/biYBH3y0k
6p8740ScOtGhgsb8RPHgMVnGkYS7k3y08Ukbv5jilieY/s28qxHgzn5wgFUg
qDzkne3PmJ9o2GaE1MN3PYmXUWZsc875vxZ8jh3gIB+lMgsd9J89bADlLbr1
cqwXo5iytm/38oKs+/O2gTLPh4TSGhGSTdTmJIVRZ1HHBLR3EhgG/bBlWJAF
D9nwmsyfFaCLhZveIwmBedfKFRiPmwPHZ1Jou9EpoSiwAF09W7QVvhyEQTL5
yFgV+wrG9utEIWia1ZwqgRMGHh1H619E1s9JxQjrbi45L1pQX2RwN4BQtvrz
VrpbHOh2aJJX+oH+SAtIdHaA/LAwM3qSaDCoZ5aUZ4CA0a/ETINg85H61iYA
IjuTaQHT2Bm6Ea3VYYObWOz0cf1ZL0k9jMXHFfhdnT4CVJXDAxKsC4Uro1pG
mCd5FrBN2k041lfxOUeAWW0WG2v3vEvyDn2s8A7EkkD+Obg962uXeSvmS0uU
2z85VJnuq5/zCDej/rY3x0K9EPdmxvRoAqCCVuPvCeREswzimMRun6LijNRs
9r46V4Cp5GWQxM1noJonqPZdsboah1h7krb7TVyJsuY8ZQvl7kedhuYW8KB4
5LryuSEkbpgVnIWdmx2GjllUERjqDMIwKpPMiY3UvFGFFiftPcPdUMvqeOq5
nxI1ZqX6rKN1rOEPiIsHySdKFCvNloLh3mjIZRKbLuYuk9eHijE2hkPrZKxo
bcVDdwd/vGKBFhULcKwMA77z5Za7LN6xdWlMPZY9P1Y20PM1Bpg5oe65mod4
zHATV9nZBzoRVOQfwhIq7Ni5FJuCMwBba7dIakZP446y4W0zwUjnfM9hBDAN
tzfSVctcz0kLXQhTSxVPfvIqozLGD2USVQJKTy3mpkPrfkvv8BP59M8CbjIi
JAYQpmX53s11Q6YjKHpF1tGj7JJQj8BNMw7OvfJi2YEfT5wx6skBhT/GJ12b
bpWcO3SG3/jjkbLhpigOWLhHFuw+XqDu50VfF5zpyjSgaCkyyHsuVwx76j/u
67bqTjSbtFjs7uQfGEoMBe8xA1twTAoIQ0sP7cpp6G4JeoZ1RetNtJ//jYwO
Q3R+1nAIeDv7Lx3oHdmxBbzZAi/K78Ej0EngZCF4cYXcPaGfwRo1ckW8Mdb4
Mn/AI4OK7i+9lXWFx2OfDnx7TJ3gCRW8bgUJ+2+H21d7Tl6v6dx9oSZWz5pc
UUluntcSsD2dUgjR6pC5zQEo7QugKXznj1Y9pe+uQw4QGLxEmC4nt3JIzAgn
v1pwSLj9N8C6yHphE4J6lrF4jgwcvh+5Wh9kSEPl9wkD5FVPzlqNUb8PyIw1
RNoqso02K88E/DJGOTnD7OFOsQQKDNdrTQSGRmy2EzicJ0fYpGdjxcENeKhQ
3JeqtE1RA1UbYcyA5QOjZOtAWcz5HcnWW+aa81PXH6hW0jhkjgoe1JXpLLFk
4I+BlygEdhla4xzr5x/wkG23ddIuCZyHDn8VWEjrf2G0uALDrqf75ty3/mPf
g9JD3lV8Fi4UNSKiPagw72TfR0RbhL633AhEHLe8wc/ORFj3CbLaRdjykxye
NlA5BGL6RbtOFssYeIkZH+Rb4TIiRTX+q4qbrL+PN2H1YyFnAye9xMW/fNpx
Qqz1leJk1B/mP7sdQkaR8NgFqT2flPIzhGJx+dHxdGQ5mMnJD31MpCF6IpvC
8G4B2EouIn09771CuaCbWf+TQj4aV53ymMj5bIqD9dCULFe7VqyhE6joN4gb
bXBCq9Q1Xv0PZsLIw33R8nhUUjBK9EilX6u8qBKJb2AL/+fQa7zlahPkd+d+
4aACYtoEPFzrkJt/mOAkYyh7bA4hnD8vKfM3Ux14IejTOuBdXMY1odcgH8zf
l9P4ho3opqdcVQ9T1h0DCOelLHDMuLGujN8MB5ksZTF7W7zGEteWtnKzV7Pp
aLAMhji1I9vpC2nO2+Mf7vNv2oNRIvRoCMX53wTGXfLJIqoR5aAXqbcLonLY
A36bPwPmk0zAi61Kqd3BjTOiMuKyB5A70fK7aE35fY7kvInzaJImXkcLsUlu
VhQDmSry7JkjnJJ5NHwdU3pKetOAJgVuyCZu4zbLzlpbveKnhZw/nGHrPW5c
M1Xz8UEQCcau31CJaYt93iyvy5fnziE6VQjLxRsj+AYwka+/Up/gFChd5jgm
PsRrYOf7qSvIKgFzHsS84+453yshIonVL3WPzNjDXajTUS7tQSrFfdpfu7Na
2kOxwXixgVJ8Uhe9a5dNnc/WJ+n/VUwccAbpP5ijvKaZPH3R3yPdZe4d4wHl
LDNkoY79nNN9hCeE3uA7JTjWiiAb0V4of7J9h9aMatHfW3st0JIEkLbuzqJB
fXalVKmsaF8oRWW6/VHNezshU8cSIIGuuTij2+o1gkgnK1CZbcr7FWBDeG9M
TLJZ7CmB4U/2MhxPp+MKdDr6fc00bfUNCd9hDxTUc/kaGyuKopXLYlyXNScO
DxvnGYnKaB5F8Iihw4UUL3TZPSKrtD8tG/MhRHeCD/D8tZDHC/fwSlF2j4bB
rlMrb/p2tOgEyUaVqNKb2RPuUloYl14r0TzX86F6NnX3mVN41+4VSgnm2PQT
GO+jLsY5F9UTupli+u09P/7347bToGpbIS388bFcxc0Yvmfg7u8H/fnR40AM
bALFyMwJK0lJDWi5yq7mMJ/pgcJ1BS9dghVbL2G99XwSM4u/woqDGLzoKraD
0jTpZ/7Mwvrm6BhnMDQrgrAjfvfwMGibbpnQ0d6KaJ1ArAg1i+0F0imDpgMn
shm4Dz9b1vhEJg6cshlgUDDyvi5TEzbz31tmIsbBqI6ZH14lYSQqnDjdS8sC
kf0nAGhVUawC3Ppd5OZnjyWzQe2hpGglAETdm4dz73BQ+12l6Z5izPU6zCos
/RnjFKJlvN/h2WPQKdJVw+SCFCxTNVMJzm1amaIi/sozKg5OzL8QLMvtIZp2
/QSLWW3p6/7ay7dXOyLLoAtT8q5vWWxGCfl7ELlYktNgCA9oda6MAg20uz4n
jrjzb4urNfla0NA0DAyRefPuZe0Dn2tW0nohOCzcrfv95LmTGoMsO5aZQvok
stWa4Ur8wyFIvjIrJh1FwZU5+fcKYtwRMInmOmj0GxSbunscfzbYxpJaqio+
AwL/U/rMtguXpiE43gsYPfCYqeNXq6S8ATHy43o3UtnQLyeS3r6NNVQQmZqB
D7LQUdOxd93wEDQk3dGaV2RyVVvwATSWLiofrLH6bunX84C8zexPB8zRrXqk
3lnNGNhXnqmB6pY8xAUR6rQN6/v+sq8l2E086cMCwZjMN5W1VPLvwCUEr9Yb
GHs4iNVOT0lKhO0DvdJdADHXAFsaBMS+TxJoJyfpySNzgo+HEdk/mbEHBAxI
L53uwfkvdTOurS+B+/c8yCT0AQ3fdgZGk/m8mP9ubUQp8iGcHs+pTEtOQz9C
rX2UF4pv2ri+ruWkzUnXLffla/zc0K5CKc2/qyZdIVE3+wRX5iR7D4VD233l
YvpyNDUJ6+ufeLBV6Uh2k4DR9XOlOsv5Gf2xiR3Jvv2/eKCVL52L07srLI3t
P5nOGLP/BewiRPYz+gHioenQ3+BJlFYo1u/NwnmVtYkGY2woYxs0bp0rhp0N
Hkz7AIKCecRLq1YnI+bVUBY/Ef0ku1Wofxe5WwpoXB6RZoj5XDZsPF/SGIum
BJbU+Sv2Gi/hmMQrO7tSpheWzPB/xjbk4PRC207LOQ+cix6RfS/M4W+02daR
Fnomx9brDd12Yrwj02sxY/CoVwSD8oc3f5p8/SbmRB+kOO1WzxUm1AZh7GoO
MF3BorYWupmrFCNIPdAhwzmuAztw0iGKZndE/ZEchLIAHWVNZ6ARD11IBaYE
sMfAJWK2ntwoUZyOuiflCK19aMjMz1S2KaqANbsdJi1vuxwdXodd98C5rz2R
rCWQqC6o1C5RBy3aH1QLG9xqzEOywk/kp5m7xs6NOSgckX0FP+JMStkCuNs6
btTiVLkQJB5V0qDEE/OWnPzsQScW9UyB8nSynBCs3La2sJd7mVP+jnCjRZ5z
iH9PpYtUprnXNY98M4IIO1iZtxeW2buQly+f6a/hNvAFT8RUrSCU6r5hxBiU
1FAzMM1a70fLC0OzSHkqglAhElTHV+2lAjuL89JScv7//LPxDwd8F6ie7A8d
OT1frE6+3izR0pmVh7qqXU9pfJYdZLDzQ7SGSvx2uQKVdB+PnjZKXmztQNxT
IY4PlCftNqhqPW3RSglfMQGtVHSDUhFUH8ZUAy0jXqPapWIIAW2hvEeLr/1T
SOZ+dtf13iQrDFqRye3MFxNMpCFpgdHggxr1Cyz9xDs+rBD8vEvA//oKBAEa
oIKunJRoMxipvmfgxmt4os22Wm765k7onj2eTKY0WZE1IhXGmKNZdyULS5Zh
WsASA7nhJVxtRYYsM7TgYY/EeL8Y1t4V7xxdZvtOlH6Z0VnTf61nEVKldlbu
DxI+4ofDycw7I5iMGKbw2f1K8fDJyMjayULqMwMY5FpwsWm22AYEn3lGZmxD
Te7HIGFps+5hN3IROalEfF8O6unYcIpU/IAScZXh/OGvJx6FRiGbPvrR4Wt7
eK1NQ6bHbdMxZUZmO7nLKWP+YiNiGbR+trTujubJBEtSJNE+JL0Z7VMk5LXv
2exMGoy8Dv4giIY6KE1lpkxoDqgsG3Tc+tNIrPUOy/t3c5E96MiYArBO9FkZ
5cTcznkBgp94lT1Fq3B7ph7RG7+zCjXLA6vbnM5LZJUDkGICTuKSt+Gqknu9
lMrwuNm/ANX95EfquUqgikRZ4a6rmCg/jWcmM8MImgrfCsweGXA+ldikmLl6
TX/YJl2N7bSkrJ8YaWIGD5dIASn4PJGCZ8WmCyxadJ8Iiz+ijOJCQYYSgRhg
BvxzvGwfVgLDoeJn3xSpbq4PARDeiZttO/1tMxoGeT8qVOzDFrg8sZXPiN5T
budqtuYWfh5cJ+0BYRpctA7tWdRpPe4fSA9ig5Wr5VZdZw31DoHQTOu+siVa
52T3qMoGObk6F5F6f2GYLmmxtcg/ueHsJrujYXAT5WnfWeKBuLX07yFR3FgF
9Cn+sBYZqbPYoWjvAeJ40ai/vqx15w5rJRGErTFHxFlH1uC7d7huqffoBOxw
ny9FEGXxPIgCqETGns3wyhd2EBHFpuNSR65f0lSnGILAQH7EsLxeODZ2wVuL
YeAW5ff91J0aZvVYo1gfohW0dzB3v3yB+7vnn5UqRAWtAgSIaXWU5INJ6PMN
NH3NlZhv9JCeTZCF9XJXMoDonSomtAkOFwEborHkYtX+5EGchqaeOkH+CTWD
qlavdbFYVm7R6l3vdnKMxen6JJ5GaiSD2VOMvmpZuWp0YQVrKcwbSEKqrle7
0LFiLLwcvOUN3rcFIlNgRlDDH1l97/waiSvKmTdF8UtkL+uB3E09+s+1RJ4Y
aKedbDIcr5CcaTwEinwdokCbARniHEZ8LXluZBkIv5DXe2UvZplW0FFokuY4
BISqeFR2+8vazcdJ3oFVGPpC2kJCLqYKAC8rBC8XHbtz+eORuulfW8DqDvBO
izdAZRkL0jcxghNQRd2xVtLR+qRlD22qyqJbdLJ1vEDZU9HKfylxVn8AcUjt
hHcR7oRLW+Xdm7EMkL7AyNuQgUyPBvVNOWHIw0EM7yVj+bQLhadB/8+VfLI/
48eUUTNfT5yK7S3OsBpApC5ZbeJPxTuxVQ6RTs40NkmBKn6IxbDzvQKsyvue
wA2A1guHMSTAho7Vvx8AsV9dl2pTRObGqOPs73uo5DQW+2Ys0T2qEdHHJuDA
Ndhc7TieCgxZ7SpkHxtmEXYXU2eToNBcqnm/sw2fMNLn64J2BavUFkJm1Jx4
RC8Tunz1CEZ1RMeoXg0Ld3QELv2LAKk24L8C96wqRfbHGRjTy7VazUIah37G
GxBn9Y75vhrgU9wdP6lPpm8foRfPhXItqQRp2pCUd8h723EK6fv67H6WB9vx
Fl2FbtrnLEsYRSW7UTvFRQYgXNENzjuz3ApyJvRQjxVil2ikiLs557ya++eW
0GOq1Ss66fgYe0woMqD2nzazohtM4eWkOERNnvz+PNIPV4RxHNFK+ArNHkLz
YgZCzCvjra120gBISwuDciOxG0ceqBq6q6FnKtbj2he/DP62GZE4Y9vbf3Zp
E3nN4cZWbct8WHAOnAwG3UkntY/DgDDIE9Y5NPQaeRWQyvKEy3lmueZ7PMz5
M4NtzhrnhD3AdguEZYe6/IdDa7CujnUEfQAT2DGTxZCVCI6H6z3Zr1m8iM8z
MH/SxSwatJLwBrQ/6iosu9ustEmmaoUSR3pI9sMtwL0uaOn1IhLzo+28JPOq
oclqQgdzJRwJi2mefIMwR1Jwx0sTZmwHy0GgTML1lSKdWC6aiFdbKhp92pME
cPegQBefgHZdUdBEjEkvm5Y3QFRptv5IfQtaxLSl6theNTxw1hDl6YRUya4a
raQvYx9xgU2fJ48iY6RIai7DbvCu3FEJTjCTcPlVaQlAj74e1yzz12nMSXu3
mS7etNHwS9NuGeh7N67QuYh67w4WpNYpfuF9DP7KZGizq9NZePAZC7pK5Npa
2TD5nWsx+Sz7O8+cPxhGJRQyM/68Vrr9FHredE7gSimh+2E8MTEhv2KUoxzH
pRXSCUtlDZp7tbZyDsjG7OeHv85L3XmXcrztGK0YVeAgFacWtKD5ndgdw0Ot
JtezcfdZh+4FMkD3heGZ3mXiGeJqn89zrrMKrEJuTQSa2DUKcYtu8KjGsioT
g3zal/KTgPFc1xU4T5shZiUl14Dk1ua1cd86Fc2GKXRA5v7LG2nb3Je63XWa
IjBuJaiFMsYZxAgJASPCJFPxnLrvhee/0xfGQtQqmDMV6ZMM6+Ledv9iw5Xe
RJZTHDPvG6/sv6fMeHsPaiBmKDKhYPSroGgcUMUo7GkJ/Kl4sOpY6dqxNjBX
pqrqxuiLdXwdCqtizt4i6jAbEVwOA7wUMYnE5iLMNOe2E8PzAKPzGDFqk+Il
jwiKSs/SWp+Z2275jHAPI589RlzGxV8H9LYz//QXNApf740di0B3qavdZ1Ul
gFHK37j8OODxo2AKl4lzQ6TwuMFrnLtyLUwOMweClZy3AXg0gEPRkv1+OSHc
tRdcj/riKl3LpHs1thRRtv/Lzc/vLgBsZz3Zn667yMO556VJkV69vB6/OOhT
4yNzpa0yq+R4tk/mhKY5LAQvhcNkTyeQukQVerqs1+unJ09rGwdL9NBrv614
m2BMv4O4EXc6jXGNdramFnml4nlapPE5Bt1uBDBEVqvRlZv29LIQ9PKRvXjp
alp52pQaWwyUQ8m+Iho5Swt9Lh22wmFy8+I2t++20xpQwXr9UQJZTEWP7/tC
8oyNOjA55NN8n5jt9ePHRa/eb5kPxmZtILKn6+EL8/Ih8MN2t1nA55OPGiz9
yNk8QNd6+SGwbXM9Hmd4z7y/QfdCQf6rQBpWyMYRRH/Sa+o1Z8242bA/0LuB
GQicWrMrrqSeA8mY1haTSixQE46b4ovEtxZG+zm8jBuMSuS1VEnGs42ABrXO
5PKOrrNGOEJsAiZpGJECSvu7e/J2cTXRnXzc2SgF8ELPRg7ke87oDI1aFO0O
Y3m6KJ0KHD/4oW/7vTHOV29duFaAU+M4wqs6F7aBbk6E04ts4JW3LCUK4BiO
df1NmQBNT/UA+c4y4fy+8vRkNZa4cqvi1qsF/eMPt2VgO+NF140yPWkfTNxa
Pv25OVTfY09jOxnv+2QWof2gBTLF7DTEMjX5zjPhvs7HWbCiKORaThcYRL/+
sFtsmqySLY8D9sT6vo0T7X3lpwIkXMPkUNYAifc39EMeHJcBUf1QrovtZYNj
hL8U3OrZHNLVXf59x8rjFNTjZoYYuc0+t4xnVCOHIrvvQBvGhc7X6dSGqBWW
hj082FcjqFXnoCfkCgpPg5dWLL79vHjoWibQAgy5Sic0XbSpI+kG3As7DOpZ
5E8HKw3vnqD1CY+/mkkjg5HsSAKkRkLqwTR14VYrq5RTjBITPHanw9r0mB15
xySRh/CM8/E7qJfPzJ3nj6dwlDG5KB9hPRbd2y/FvPCmJAPrcc5UfzFixgiV
exoEbasbUaLiQP88YWh2jCfx5Cz1iJijIk9lQ8hk5KekKAKmy2jTSZ2Fh8GM
UC9GYxR6j61ooICaTRn/O2a3bgesyGFxk77wsXTkw+Y5mnJwNeaeP3DAas+/
ID/y268uMLLd+C3rCRbAjnPRv/B3OSDJUktCdxndo0sVd7pioFgzHVZYJAVy
Aau+CUHSclqJsYBt9pdiulWWK+TfFEcc+GudHbMpqIUUgrUVhPCEn/5yMHNb
49ma/Eoe6UTsftJlgWvYL5uusedumEthPM96fGoixjYim+K2UZlvwa9pdigZ
4tzmeTv3oPWHidndsRd46XMguIW99cX9AHYb5+avofZ+GTkb6QjTwJqp2PYR
y1MN+6EkNYC048OA59r8PrseryBf9xAXyyaSdv8WFPzU8YlNIRhrjRbPPsN5
tXTT0x6GLkDnHo2rfGG4u3ACXfyXgiXVezqR5Zvxty5ihNI6rq6DrC1OclUK
e4RfIvMEOnpiO9G9PHhbYOlpRrcnwvj8ufiUitd4SfrmkouiebOn/uvT4K+h
Wm93zFt++tlBewZLi4gHM/pbdbKGk4C10xlyJJ/+GRiMKbk8L+Qe/Xgc1FGw
BznGn8OLBZiJBukL8HmhaFz760it2QI/1jp4fEitTS5Cri40/pcXlKLwkbya
0Jq9XQqqzesKjRnwcU+vQEPxq/Wuwm0J1PYHJw0WbGDbBq3KDV+9TQYl/imt
KSSazEDzQ6pxNLADsysZRYBBQeQsP2dvf5QIx7SF888GWARlpOcTSxi+v4zS
rMjIQTFHRqXKOBvfBF0Huai6zzaQGbTvacaX80JrXWrUif4XOW6ZHZsAFI5t
JcigXds7Di3/pbkUV6+MnTWPTRNpxAKmV5yJ7f7g4X5siiBsNxT/yFUaMrfT
57MhZOr7i/ICrfR+FOMUcolC93As73wlxWCtTaJHgIM8x8ELvRo0ZgMDkPji
5gijoW2qYQPJYuTLDASYRwooOIikpXkfFOx02ottgfoRVlPfOIGVvxK6dG6U
x/KrKnDqSPbYIN6pxv6Om/R9TbtcojpU46BScvQs9qTmHMZOde4Bmb4Khf9C
Bqca6quXiF9TaxAzt5S+U6PNAvLeqaX2JZ2kbCO19dZqmNBPeh+9r2HdGs/Y
XWqFIWeMnGhUFdGWFiOXjoZo4SIfTmIKo+WJehhISyCM+J24MkXU/Ckl3DHc
ft2HDxoB/LV77KiP71wsc8iOoOAxAXtisuHyuN4fBBRZKn4ogk0q6gWS1jP7
jN9loVNVD9LTZJRa62P/vgPqeetg6Nq6LQ1Pb3Ho3LsYfV4kkjsvf6GPO8Dn
UekibxTSDAbT2k/O4HmI58pC8kcGLqQWSaBAn35mV9OpUmc+KSLp+N/E//WV
O63wkWk5eubyRUt1iYWJdZfZAQ6V8surf0I+Nj4A0ZyZplpqHsgBWhenPL2/
yD3BqKxA59yY13w3c1NZotWgmPYZrzeeeeDy9PFqYEhYq8J5WL/rJLwZkIX1
7I5P4WMOOtSSMDc0svSHWtWToCwUcCWuG/zoybdhbXCuoC8z9+UwZphUROnM
9HjGMjEkQFPvtyfeG2WJM65JJN75fZboIVW55Q7OufwIEtgTTftwApc0o0Hw
kJiWHcU1u+YWqV/cJDONnzBzsACANMy7R4txVf4I02MU98uKcqE1ek7CWc79
6wOjpqzMVORb+t5QNSLZxhl4291htzE8zSF2Uo2UetrfPSbYCZIoKjHv4Owf
37Nd+a5gL/1MJ4YE7c9xXyUjDY3R/RWTtd5x9H1o6caLECDZb3YOJ5eY6vS1
qu0QbU4abXJ5yPECcHlO1Vy4Cxf5EVFawPT3Ki9aft7xqCQFRVnpfnUHEnQn
sMOaLagceSlNL4tZrzMpPBxDxFd4IN8xUUHrp+5UagxiWb6mJF78/6ii7ZWJ
ZVrY+N2D60eAN9aDCqwwmvBwPIn7wPI89teJWJGqguXeaiyf6bSPNhYkICD6
jg3vWn7lw/aylpP8whY963FKSZrf9YaYwtaxYuaM42dSiyB9Uc0sRZGYi+Z0
ajdGZ0XSvKdQMD3/0lLBsozl2nZr2uh5FyHCyRWe5c6ll9jA1rVM+455ImkK
HnegGNjMdKTBn8dQmfluNj0crY1iH4k5sAZkHxVk+2n7EWfy718LOeN969fj
UXmuqJTqTButaqAPumzJ5TVB9vJJXiaFAqIMg0hlkuX31rWPwFfao1H1aEBV
sZCZQZSi8A6GvKJwooXOZWnY/ty59ceYGHmyvXdGaJO+Yh0YRiITAulU0VCn
upBUMoYK2z216lJdbOyKQ5DkqonuyPLhgDwKK7GMWhlWAIQImYONEnAx2piE
tv9tEs00V5lFmSWYi9e4nBRphZYlgSeSjq4YHyGA8L02bYTA188SBSGWbCpA
Z8ZXVQAxN5sqb7wLoAEbDCgS7kN3lUuIQiZI+DDkv35jgl5+d5zGE/g9OtaO
peO4dfBjQ8xKyc1xarlFUxKAaJ4LZqi8b+3ji5JZQ2uHG1aw3056Xu5J6Cno
sv2u0FcT/o40o3kuQmOGvJ+m0wlhxD8xBW0GSdqCRRyf3hP2IANxh/cU0G6i
FmnUcXV95GOhZvMdDgSEUWBQtafNkR+dwI+WTans89Jsqj2RbzWjdN8LJyPd
dXour+xamAtZorRA9yhL2RNZRtU6COditZSAjL76RZgO7yTYqtUhDIhwgJns
X5DJ2EHiBqj69t4t2DWaJUTIEHqir0eJXb6tNfj6iYYNBw13vpYqkZI4iq3o
zSLwpgBtPY1NgL2bBb/0LelECnU0uczmdARtS0uFxA7LtBLOHY4GSAZK6Crj
BN7d5s0gWh42JhnNXF+c8ZCYi2w/IIaMNU9d+Q7t2qedwgSNxmLQ1mNPfKCT
Ej/PTu8irGWLICIiTPn7MXv/bJQfNlT5/U5Tr1ErcOhEONNXire4xvfxhPST
cwL7U3AYAr3qJTKgRd6L2cUw1prhlOxYq8muBLq4Ar65mMJzL+BdgbfqGC7b
21hJ7O1QFROI7d3d9GAtHASfzbXKEVkjsddkLJlOm6+vCYB0SdYklhYjEHqM
v5DSsWwVj0uVrTU+os/0Bao07Cr3IZY5a7MUPdghPuDh5o1N06IYtjKWhLP7
KS9swasWA0xRNvUtJZaQfrTPUPkJXZW2HWYoQeY+ILAFZIBm5MmnnIbQmrEM
x3Mx3Yv5F/oPkYxRm+On1bjzurLhHcM/riwNuyRHw73i07tcvjeqO9hHDuWd
wHFhR/+chFv1/ZkX+AfjiIWeSsWX+rFDrCrWQU5rBk23iw1HGK/37sR1UigO
I6NXfTO6BfnO1woAZUyDQFY8yA/3q02XAdmsEJYxViZXasR5tC1qsXHbsgr7
WTUm51ChC1GOoOYT982ne51XslqEFDr2zpenDStdHEyLZq18dkp0Py0IpWwP
uEeNvo053V5RqR7dSvg/c/FIS5BiPZ3gKySgNs8bAUzVxUukxLlYr+/j696Z
cTEj0Eiv1Wq4AmJRFteT8uosIosfTfScrYHPa88kUadAEiV5t4xJWVK8lfM6
4ir+eJFeJzotOBwY9ndAx2+YvD/8+7hjZbp6AixDCW3ZTePBycvMuL9uZuyU
JJsE1CtDE/ls7kO81dmfrPk5zWaMBxn4dfdruApKW70A3tfnPlU7ybsDa7HV
4zEvVZgM6epJp52GokQQdsJz7ymdu1D747bwsefrt/4rpzmNQqCxTDjMq2y5
hL6S9SZPzUJPxYDLpUHvvP6ZgdI3SNjegza/lJMUTKhDItW6/yMrCQ+siGjn
Ydi5uN91qQccGMH7DFXSJszRGGeLeWvT0nEWWrGeo2HA+p3trKtGU85WCM4H
g3t+JdTw9W9wow+htBB9u6xVgW/IZXCCaisGahMr2UMlFhhROiGDuceUy91i
4RR9gOR33JqXirxCIV12ctHIzm3DHpYRmiUh4SqJ/8kOLWAys0+wZHB1kWLM
I5oT3iSn0Sc64lG8beKSCTSD2vjNJPY1HU3gkaG1mhXT7kIqe5Nafz2wDk3x
Eutz68NjFvc7/KViAL6qbkl9rD3MP8vKPcKoOaPck7qlpFrpSwNcOw3TqZaX
z9Bel0VwRWSQk03QBLOpsuw8nJIXGH5F4gsc7YhQpGAa+8X0sOyFcFgxYjPG
SsH12fbsVIy/JjKyK5kqDTk6h3EaNqb3HM39KR8ATOEeiQVR6+dAENOjXJbh
4DjT0x9waAOyAS02hnSF042CpcDbuSTG6gwLP/hn66Ws0g44wd2whbG5FhD4
l+2wvnugp050un8aUhLAtxDyKRZtL1QJqXC7gLeQugCuVk6TLUAI/ZLfBiua
Qg+WPYdJ5Fq+IATVb/XwzCpIL+OxMiPQNqRvfGkeSoVmIw5LSvlEnDw2XPKf
2Vk4siXjWMgAzsoNES+QArrwj6DPG1hCYiMVXysvgknq+YZWbiSj9LBeRUl6
IvXIeW+6Lo0hmbOiVdvzFJLXJm2gExCDmb1zTsScGmRFnK39AKNZQvIYT9F1
NZiZB4+JsBx6uBXbRBRxoUM4ObajRv3eUV20oqo9nWq9Agkk1CRtasX/H7cR
OjxXaJSwpKV1J2zB7mMHQOGwEglDIbiLttNek//5+5udFcA8II/4p7Zn9hf2
xJl1TXPtnHIRyXRAnTPV2W057P7cu4RUP0oN3w8RAImJlYXH7ylptrF3kG/7
Cwqv8LvIG9aM/PWuX6KZ4u55QmXvH3VY68kdtrT11+8rHJ8YUy7mkx8JD+Hu
83RH7wtxzoJBXqERuUw0SWsljAiNnM/YQQJ+xPYw4wJ95Q7424KXPtZRJFz+
Val4dEzYHAo7WqdoKHeacSL8aQKpHKEKUacSf9QyFEt73z3DqeJY3NELbk0d
nluLAVAvnh2LkhZw1t8IM4TBiOT+MuQZbbrscOn0g+ZVhwfABQwhuvmsikTA
DUdZflnId2OGyHKNzJKa1gXhjZA1JRlkkyo0WxFJFeIHtNhIaNB7aEvsDaiM
2lbXaYP26vkHHg/Oj38n/81TTG0GJoIfI0BUhERRGmNyDumndSKczKJaeNMH
YExV5ovjI42brgNX+kX4PuUl7pFF7ea2iRVTBsEVC0gMliXy2U+3qju2kwiu
VqYi4GZ+WZsFBhYNjI4FFwFbAilD9TbqwCxeWS8NCtZ++zcyLiNNw7T2tdtM
dHiFMUvDSrhwIYpFo1ooHfIKnAJSF8vaGqiFOSP/V+WT62xmmmMEQBLxULKG
Fz/FbwV/T20iRBykS2Vy2HEa9thkv2T3sm83zmsgVOGh3YVDWM0m5g71Sp/P
w7DgGkDzvPBM0fJZWeGBzZPON/Kb/wpN20iOxjY/9hNZpPYfoj6uz+W5vSum
xkjTU1vi61LdVG6GEPvNqlSxiKNkVOMBM4/a5auXNYF+pqr2lFVR9CQZqA21
/HiqtoMJOX0rFxgwLlrLuUx1jCPbPatulf6w3TBVMp5mMy8lIuRDOt72pjga
FSJY+B9NHy3q/pOSQbvLJdp3amrCpJGxTQci/hiZifXfHaz4FNU7+exymd1F
HgX34DHhew5qO9Amu2SnMkKQgN6B11WVYxwPpHFshhqAp52k8GrduKWYGktZ
QzICN+qMBy72pIJ9qv9kB805vZq63WCt1eQ00m6DEogXgNah7iiQTKxnwrQ+
23wABVUVgn2pA4lmFCZuqkkdreAqimIlrI11a9YOoeaKplk38AX7KmP/HWE3
btUtXqr/jDUn5D6kxJEPz2YM3teHqy1gv/VZ6/XjhfV40IZdTMlr4YYUBTVX
FPAw9QexttrR/te7j1zcRTc2CHvwcZxhh6hlBXRp3AGg8zus/JewA/zJcQss
gde3GFj8hvBpExUBGHjh+S+lg3vUF4EF2lTGmsOz/6MfY2knhgeRCla1ji4j
HOa0eFpNSqFru1BmoO/3E1H6Fw9VJNT6U0MFzFB2Gt2K+dtrsnGmUl621qJx
NMtoItKccbW+rt25EzhTt+DmcetRZPboTBRLxcdZnmMXrl1ewIDEBRJ8sYvp
pJu8/QH+JHttgNk+0IXpACKhd/wOmIkkINLBzW2ErssXvV3cjSZ2ikJF8oYZ
W0EEHcfJYx9dyYhISZ26aWnGuh7kzMmT41tcGgxucuft9FCt754gL6wIYsQ+
1lMU2zLgCFwlLkjJnqFtx1c2jnQBAx2L0d4z2hJfKMRqYAGE+FkkvmiRgxqf
ozzmVe+KLOut/4Sn6EdUTQtqRh/OW7HD4nqrOtR6x6k7iqlybkYQnzuCEpCv
E6DEyG20p1C6bsiM06UnW8en7G82ahvcUuw3e16I/Jn/A+CX6rgix6HHiFm2
yUoosfZy5dNXAO16mg4+ngwsCTjZfiRbnfrQpS1FsFxGhq3lv8iAy2wUQ/vV
18J1nVb5kcj7MTKQ7xr9yCzoTd7JDzYOmnj+pblcBMfEitJLm/rRh6YHrbIo
xoDoXtqCTbCREuW4WQG99iJUY9goEhZ5yridOuZ6oIdbBW20KeeP/PGUIMVX
gtbxRw0v88427mhYBLyDbo7gYGF7wwtHGsVNPqRY+/gSQ8hmykrOvB5J0onw
ULGyFUoJgcdt+96kQ6+9io02hNiO2+HUivJm9ooFahjCcpa2J5mELUovjUEO
hDigg70Owc10Bv0/BeZB0i+2oN3MNrCtdWkx0Wfk8bSz0fY4GCS4B2X20VBd
JxD/z+G+ujwHg5UY9nPYnhjtkXjwH50iRG1MRHuB+JuTs9wbf9Vx0fVpLH9+
9GK4VbatPJlX6NZln2qhmn/0OOjK70zkyLvKDgz4KpfVsJ6LPQ8Ywbf1h0XG
wyZ8VgXPPpvzAcxrwTuQsRy+rHHCYVzWT7I2UjEyOx8Nj/8a/W0Q+UwEJn4L
z14xtPQRKE4D/Gk67WuIvV4+gewA7RLobI8farvAoyxBMM+4GacTt07CCE/T
7zC7OEVgWW0ForAMc9IUbHKOYgl07496fWDUMgLe2MDmuG76ip+RyHpb70YY
1cJwjlkOGVPEJoYqzwLgVix+0uBsGUuTiUQwMlwtVFRIyygZMFHsvZDw0hvq
MRBU1lCBF0s7ey565yZXIivIp8vwrlqLNtGNG1R8a077w37th/UY15LWEIC2
ENLvOSnbpBxBVHmU07RmJwBMFeAPhbgBRyjMcBDzlC8PZgBnvfjtA177ykYd
F8ric/zKqJ6jo9B4X4PB2yK/c9FvwPJrtYKaibYuIE5OCFw4xpXWZfr1jrGJ
AUCY7B8DXNwtFmGhvorBzKbIGBBVQ3PELMf3S7yurwDsrmYRj/tye+FzE6bh
6pqn2ExSidVCRtLThSCOJkqxoKAF7wyARXZRlu0wN3fkgQurL1gt6L7lzYDu
PoQxrRLVlUqIZ4/+Q9856/t5q8QQAK20pfdsVORaK5oCAsVkWtHg9hpX50ii
dY95Ktf/q0pAww5WBJCwt0Jhk1wuGrbZ+dqdHlG01gdZOgX/6/AgkQBb7t8e
jYVXRWTimhLcvTdMZxsEVZj4woQWT57ZxQjhs1RPb5e7zYVMr95Yii8XqNpZ
YnDfMDsNimpjYZJq4HWyreg92W5lco3MNTkh3o7TmxJ4h+T+RkPxpycLn9RF
XQUBYN8KVK+7C8jf0ycIQu41sWphZlGQaRFgyyJFCfrA3DxGDu2GpQbHYLJs
8cjUgoDQc8tzBltz60L2eqnAy1dfb9F5sJQVkWlfYxJLnwL4UYVeaBGVFceF
DDUi9vQK8axYHPpOCNtxhJfDgBlPAvge3pmVDeHOMtcdVFjx70FxCS3fQu1V
am+KQw9CaqwwD3vUXsT5XIuC4wLDq67k2OCj4ODoDq+jlYU/mVEcW5glXXQS
Mcl81IKOIFsQqSIhP5s5f3zS7Jm5W4RyMqHM0lvNuxtg7h6IH94V+S8S9RCa
hvx/jZu1o0ZxNfNKzsiHkOxmTH2CVLb+KbRHxYCjjCudNZXjH5+fwGciIGNc
3GTPVSqdRlmLo0HxW/HaM3LsN9B0Y7pJpwWgkn0ACZjx/RHLJAB2b6p9Rn2b
kOqAhErK8NUKKw4kzN9FosCTzBYSh91ZpgjCyWsByBckOsS650uW8vm0mu93
EQRHq/ZQVGBka3MUY+RPwOmMJr+9cI656bKnJJMpx9Y5xnkJBvTsyF6FihMK
9wG+EE/p/2bz2E+WvN4QoHBFKLKfHVAK9TrCnl9NeWzPAGmIUHXJFXjBEimt
+P4r600EM9hLashlfCxeb7/PKpPv+mf0crWLGdTmMRqYvFI9+NyomGSqKly2
ntt0QjvnvcZDxfpgbgwLrLyghiII60PAdvj4E62ZWgtYn1O/+GlG1f0SephB
c81mI5GI4wEXP1EDeWfYynbBlHE7DmosJ8b4VYWBEexc5iJ1YPaKTV0bGybV
TZhsSdy3jbmYoXSBSVda+pRiLtaJL+/fm/Na1UD9eyXsRoWYS9vhS3Ya3y3s
SfRprjvsm6lPJ1S5J98k76LfQnLt+qZX8Kts+eGvJJMjfu5BoHGdMKd41Rre
xZ0fvSqDNNYkci+iYuwumBbmiF+my4MRisD1AmnqWJWKTXLgWas6emRyEfi5
cmVcsNOywStDqXwF1Upte2pbQnAZzGQKy/Pl4zwaY1JmniZtNcb/M+6DKtRq
NC4H6etGo08/rfekTLmkPaYoHkIODFx2zzsJMIPJl7FqoGudv3JC83c0HAAh
IVgT8mGPR7/7BduaP/wYc9aPQoHQpyojIjrOZavPbjt66yTBFdlVoR/0GtuA
DVffqelyVlDhA12Mr6LYV52l8g1czMKyKx/k+YpDtXB7YbaeZm7U+vhCWgSM
djIfh3sEmGEXNZ2TEpEczceL8XdxVR8X2GnWjnD/yGqsTAOURu1C9Ow10MEd
kw8HCOHQkXFdhqbzagXCnnDFnGvrMVmBRnDtB62NQeiJ2137JxYJiiSn4jES
+SssUfbAeAUivgA4oWUo7vAN3DyFfC3LRsgdH82TjtncGQO/G95yFEjWa3Kq
C5rndcrvatQBZqwa0MJeV1z0SS2IIrPzeaVNiJzN7t1DN7Ez7csPQ87G+P0Y
46kLpg+jOVhqmC2xBzp0wizw/KBkoDDCPqZd+AmZKhuErQCnllz611b/4mBA
pYJ5JSKzGRPGDSNpLiWSJDlrG+Yj2juM99bX+kRACGocv4NgcTiPUAaXmKm8
Vi+kBBMndEGCVBUSv9CvGEVOIe2yXH2iTdKLvvDu6Pmx0a2VKet7C5+2KBji
/gapcbEBR5DK9RxfRXVkKAt4b5yFBBDmBBAtzXW6gMc9JiIdThnRjPHx8W4I
TsLcEYZ9jowK8CtRgbt+3roh/1BQ5wKMvMb7/Yq7h9TzDhQdn6HupW07LJXS
LYUdByIOvk9PfJzKrjHOn8qByDHp9wMJay3L9owPYHh3ffTpnyayyqj7f1+R
PWM2gZWPW4VGmyqh4keVo/AxA6SrJdKTEBedfoBUHbcx6yZppLBTcKZG0FVX
yUjNbHd9pIA2ZO3osvDZUl1mSBz/PY5chNsEjM7vHTQlkb/eY6Qg25WsjvfO
yRFt5Of9GQHOA5LwGcwufFcWN9BK1q3rSDeHjLKkdTocIU6Qk3x4UvAyG2F/
+O/Vlqjz552AIzPov0IsyRFUmuOysLUmr/vnlMxkOOAKZ59sNensms8G+5Ko
Tts3/vKqwZPFfE4fS6s66Gtcoo/6Itl7pLuf5Vppco0RfP23h1lMOtNqQHRM
oSRPlGlY+PpJvA2sPscn2uZpsIGalmfln9VNV7sZgL6I+ZKbK204XFSjwkVJ
yJvFcfZm9Dwoj3FwVzQxpKp7z8XbnP09ZU25OWgQ0UfpSsbCAejGChmqu8pw
3H195BmRvuFPIKAzzusbgGzC62rvKIPTUIfBSUJEpTPnXb7vYM0ZcHFDbsDV
6pjFWwlhVFZSVj4MyZZnRZ7UA21v+RJC+qnJ75VmlmCi3SIrHB2je0UdM3SH
V5sEi7SISez6/KXkuLkUCsLT3EIPtT+50vr5AOFEg7f5J+GfYekqtoGpqzi6
2OjVMNWyZ8TIpPfj9PSTt+p0cSuxZE/5KZsi+KrCAtCR35My2CWzpor0ykGE
ZT5pe488MEnt+8bv+tqAZpU9QTRmSS2BOSPIZu/oef+rALlM45nDe73WViD2
3mZRFsSv1/Gut8eANnB7OUrE6g/aLa93O7y8Br30Z9uut4UfZcinOI22BZLS
SxhKYy2Uhruv3CVR4mS/2z/FlJt6J7Q+cFPnIBYKxQcak4tAbPqjSnO6UJfU
/hok4U2RSfffSLOwJQj+P0MIdMdsMPfL3Cxzva4HyNCxYxZgD/bZ332m7k2t
SESL0tyOwuvC0AycZjZYHUIvTPlUKuEXF8y1LbiClk50mMcRjk9gQD6N6VbX
JuPwh+V4NNHp7pDlwjm/OTVEQiYfDtei2frt7yGfWTHYXHKm0AYeGkfH5XTx
OyNpTRCfmQP0HUEr/8OGLSfQFfVVAJay7foap4P26QrZb80v+0LBGd8hd8Br
ovlinAStIA3xd6hupOsCw+TuA8Be2lb96wPLBRMjipyojEkEUdSRaTmu0reC
N1hutrKkCUTMwvRkbjc5ywFSSHPGoW/E6xJyPEJWIxdTpaZm9Z7H/wsNDR7G
qZfVve6ylpEy3Mt5RwvVGQC70CyLrxpc2ckf1ZOukvpGHsIlxg+2PwvCGlai
44bNhcC9wLpPP6WjqtDSkkqvlf+dZ1O+zbeUmnPA55zQBnr7IOuFGD+4CUap
hHhKaIhLwREXb4PI2lCah9QlsiyICgDLgkW1spKq0aLmDYpYeZ6pcNTTPvct
XsI7LXjWJLEFkWKoz4fY5s9T+BrFjcd0v2p++dQPL+6ZgNQq2L3BfjP5TwKo
KDhW7wrYcj+3OdmRCOFZ519/xH/ektmc1B8VKPuHuT36mKEdwaEu3HELIBg/
ocsvSs9BOxPOZqAu8Zi4ETuIZ7x9cJDQ86QS6flOdOdI521mL68mnBQCQS0j
wQB4keJ9I6w1RqCt3I6+oHZfaFcp+iF4Rh1NjO5hR0bLDLEufLCEpqNvS3Wn
uOz2CIdsL+zgP4nwbquxkfqtJFugvn9xHIWe/8PFcgpMX/UroN4u7BoZCPdj
UkJSAusthrfEaoHt9cWu9GPxNRGA0aHQrqAVuEpeleyQmJRl/0c8RckAH7yG
yipv2liV+jyaZCJsB1Cy8jguMYciqW6zsNNj5cBizskekb8O8u/QiQPMMy7T
ZbFvRAQ37XlpNC+HgOgcjMkR58D+PZKfbvwtfV8bfhqmVxoDb6Vmllgqo4gj
JprX2CqToV6aTD0VNOBRcY9cEqpx7HWb1i5BoR6IABPAK/hlQXMf/1AzD9wI
lK5lLlMRrhHwb3TwSU5hxrdav5PqJR3Xltp5CrTqSbGR14fT6a8h+iyt24J4
b52XeIMzgy0B+dE3lSBfFh/noFRodgX/QQb7Pf1DHmW824Jc3ymG8DINxT0f
yveFLd3xV7G9Nuvke+xuwwaTGm6st7A1DBmsGX8F5BetYjvI1BsqWWm4p9Mt
dZR0fEBbiiX3jiUjGjKMqWTpLHH/k5/cDy0kSDTb7h3U00s7R9jdF8AjbhkP
ZxlBwMa3tHRSMS5h//neHE8NhRXbFsNOQK6KNUeFo2NCDTWFJk5Rpjfprmrt
ERC/xrcL+w5D6VicsJubJgIuPcwCSDJ5nNojLERm/Pl5y4gRfl+ZOxZPNSQi
Z92VCL+577lsFGBrKTNQA/tjRgCoRkAm99LUZw/a5lOEvcNSxhu5vqvhkpPc
h4im5uxjf6bf/1I7bIGaEZfmzgmY76CIlZNCUspfvZ2HULKlnHJzGg+BfwMB
CbgpoSbfB67j4XbB55ncrLHB8Hp0P+f94pmrZRMh/mU1OuN7tUE7rKTz8QNw
xOOYMoenjvAvV34QbxKjy5QVoOLBWSgeVUC70TPhNzJTkOZSCj6Oj127/j+H
QJcaeypMZyU4TTKzj3M6F56U8VVkOPKRZUADwzw7aJmheMB0+8nNmebfgpNx
IQwsj9SE2VnBurhmY4AeL5oG0CoaUIZBEfTgJP+sQYZJ2v8SjET6Mvheqm8O
VGoJEEl0RD8QRkAfdAChEPbdmPhwUgeyavnZHGnDU0qD+LtqI951d+kgGQbi
152WaPhb/Qa2PQO6gO+HvH10AaZ1vLlBASk+ybrTcBfl+Q6AcUGaMyP4dS2c
6UD7HgjBrtrL2WXpUYnc+EKds1+SuZgcoXyom7VUm0EYAVQ3dYGMC8CIMt8S
BLzPGswzvorhqpPif3jw8s/EJZAe3O9dd/AOQ5jZa1tG/57DZ8jqRgpiEzrS
gqfrTSgvhI1Z15sNGr1mWTTULf8gcN3KPy8kO4KR7mjG6euMfgh2HD/hRlqm
2nEsr7sT1TRSMgMwg/+OksiFTp/YEHqbSVkiqjuolWzvFPPrbWw2RJExk3Mt
moJ16SOytJK3sQ723QWssH+bjjQOPKYRnbDryu3JxId/DrQx+WNLnuohM2MA
vN5/ztOEAzIKTYVmtJdwCzJlH9vh5DlEWv/ooo2UjK9fqw/R2bL7lkNOF/oj
P+vMKmE5PiavCJuF97Gsu6sMkwWh1i6Ng/HHaabVypWUTcSjGMNENhOR1Br3
yA/952FDQGKIiROJjlm5nxaxvCrXK4VoTia8DujB1pyK9FeYA9dTJyUkzljW
lgSgihPNkKKf+kBDJzu2rGO2T/523YLneC6dhEw4A8WczPwDM62SFjUhWzd2
oML6qp13BDStxQWL8I/2pRXlb3zs/01IBei58tdv1eVmximVALtJQ4FIgbVP
TAfnatwDUHBi417bqDBH0uAHWU1K1AWu4mTgsOl+qtmhSsYlZmzrmUi/KSHa
JSKRfdVKP8ucbXeSVo8AwSvutsMIEi299mTjbnZH6I/Nht0t8W4MPLrDin9U
njcQje1A52BFQDyCAeGumdg6kTBegN0SI/tY97GwrPSlAU1A7PdwBCRyuel+
QmJbD7uncS7+r1qQbKqZYF47Q9Alx5CPGqleWKAfh4IczHg8cN7/CP5AdMIM
ODQCgCFJdSrjYcd8vvxWCUOkE3sKGuyXi1WSCAvhe6gFz7GVuKENPcalKuy0
OROwtQ1UB76fZLJKDlTwuQ4FgtLID3fztUbOvFctSXC+CJK+jw79EqcHqlCY
boByKKnbRQQAwG4WRsnZUXs+PTRbQHQOst3VzvBcmeeEVMKPeCNYtjmJ2+uO
9DF5BBjKEe+tN+p5Q5xVS0AXeUQvon0o/JSPx9brZFSivn88NzXEyZQ5y/W8
mxOZXye5vnc5FnF+RSNn90TWVVFffCEpPfJBtnGIU6maXvX+1GA2/+oeW9LL
E4t8Y5X2JPo3cgrtNQeHPlhn0uKEk6a8r9QEruanlSkCqBUockFBKAPQh3dW
JKEBNKqWIRFisKmcB6fIpNYmJ0XqATyb7Gbc2FYAiP2E107OLbGhsz/XZnID
zmPcOtTWio0GWIQiXl1ahCjzT66VWOccF041uCxTDad0FMnsy98oe2G9dieK
A4ViCkZgXjqLls4djYjYl9xDpq7xwmkvpyZiakAphM7kALoFPwzVmg1/RE9c
jMZOQgAz2qVEdEXDjSy56Nq0ewN3hWzQPZeO0Mcy0gE3/R5Vx0aalA5uD++7
xG9katcpFnvo5COIz7VQfI0K6VTzfu7Nr3aYtOnOigW68DqXR8mFNTCu2+vC
qipKhYF/Pnc10zqCHJbQUKEgTraCr4CYfPTICYJ4oOZLpeC95H0Dh/dfMTuh
dPpxN0Z5LWaOI9QV20M2eR2bfyMmzQMUm+UTcnb/J8P9I2QqxTcXkDFcI/Y+
vzrNq9juB2W74fP1tPGOKIbDHP6aX5eijpV4He3oGXI8MqsNotkXfYMr+3Pj
OO/1v2r/+8YvawnpCAFN/rfZoXHgRSMxGv4T5hMOkBD+KqwhjbhlyR8G+Yyp
PT7jxMp9UCvg5NfJv8GdgZOmIN4LcUJ4Q6YFyuYFDAjnQUwQiqATwD6a9JUV
YWQgQXckdi1AZ4vJ1w0t2rFz0OVD9rzFEfHrkx7VrdvjKY2Da8HzOp1vBmfX
MtGVRJ/a66z1kNEMc9MSFe4xy74Qq62527e2/mAJNEfs5uYNiD8KshbBdxrT
8GAOQxEzLoG8Voq3qUFhm77iAaztPW97gA74BmEhWfeQOmv28IKPUeHJ0BBx
6MjluLQsgk60PyKk+zCjv4l99g8HHxOZEDSPgQZYQDcXL7/i8SU7EKhQloYT
V8jfqqTDDbvFEvxsPZ5nmByP/kJ4PC5uQvtOpblXbfv+9HMRKP9kHb9IwBJh
PWNsdGTOv3HLWeQj7nDYCkCBLYqAr9vtoc2QrBNSHhxPNLOkrGCoWQcSzOtM
xKG+r02yWVfIZlf8r0lBz2QU1QerYQbtbDRquxUH5nc/jerl7y5lqymjMEQu
5YCLqCsxTIyX1HV2s9ZzRtjit6+Kvs5EDCYzGeqs7eSyrM13OzX/evmjkRL+
r6G5i8xVMv6Jp5guqBBv4v1Rn1o4PHIyiB/G1WpGXdLXowLqaUKmzpjLhr04
98c31n2XsffdSqon+2jLL1JQv1ruQGpO/X9BP8+uUq8RxkmZe5WzNUa3C6wg
+XTkFNl0rV4nT0M3bVC7/hHJvSwMiPGsEi6XzGSZe0VXPzvDWIM2l7BYtllT
z40rRb7DIr5yXSQL4598Eamfk+87OwwqX54L1oKfkjKYtFjdz8E6f6PhIgxv
4KtGuBn/InKI9NB2pInI+rIqoCyiF7FCFFXpatxmfLB5hNZBB8um+POF6ugL
KCjSlEiQ0A7jLTvpkAFImRAPqmwb38rvrKq4idFlkCWFftGJBucv0MfPBLD/
fdtVt1tPeIkKrrVyzah96ujUr3dejwj6BfYs9QfwlpdUqXpKEJTR4f45hP3h
B806YcswbPnKDOo8pXW3/YnyUX9vFeqceFYEJSoUexG9NWHA4Mco9jZSoUFu
f5oUqtDhZPfQlubNylqNKuzbrZjAyFAdPbhXBvl/TA4bdFtMueQ2YPFDw6DP
pEIwTJV6KPhchDDMNwTCZfLhwjtHLVCzlY0p+u1P5PF4wSbc8YAN3C1FRAIQ
4uWgDg6GHoDLoBg8/i+27w6EkFeGxP8cEI37hv5o4bsnGj6ku/0Wv0JfkpDb
ThgvydJbUHdVBfI27Y9QYiycrZos5oOkds2zkBIvLwnSkQzKQXmfyWWcLYaK
4eOISmDE1H2IH9oXUq1OYytjJbo9z+wOfPXF+wwspiS4N4GLlDwPo96cCeRU
cnpHWEdNFvx6FqqT/IrfQO2RqpzHxk8LvmZgEUREGufekXOsOrccoVhpL2Dq
bxWsof/U7UgnBEkTWeUzNK8JbKFqhdOkHcOaE3fb8dtZhZEJb/RaG7HkMwPf
dQ1pgDGkWrGepEcX1KXBMUpyXGaeY0xvr38Kv47WcMzFbR9im5GcajbItvvm
o15X36Xe0GIYc8WyIesfpjpHxuMypHucjlgX5OkZ4/WSJfthiAzc7FtyCpEr
TO67OmI9bKQ8NW7Z8OTd5mqGOwFhdM2/TiLoRp3N6MOvCosBhR0iF16Np/sM
hmfe2RVA+AhqmnBzTs5ktGuBIdqBHD5dffUJfnsEW74VKmSOp/pCeZU1UJOj
GL3pYpKuc9F56Mc5AcslU1bucMxPkyWUBeeTZKWm1Uj5gAHjlYzz/OlFFfVW
PCyWBhuS6/CqoWfe3+YnlffSVIu133SuarP+TwynWVnII8IneTlBOBB88VFk
9vdJyhOCXVlvvdPavM0bkHVU7f6WK42KlssyDH5KlHsZhbgMordfvNadI/Fb
xPzuRwnLd7zCSEzMO/yrp+i8dapuVp3w6lZo49OGHYlyzAGbUYDduqjwHYVv
NK7Aog4vZA4OGYItFkcI6fIRPQvR6NqZ+OQvoF+2WEIxNDtA255C1KL0bgze
jL6pHj4HlHNviOxA8BBswxy0Loyol0S+1/WWdVh0OiYhnNIJVILck0tQ2TeE
qAulNDnx2GypAMvIiXvajhGns4KDwQWesMONi12rF2DEogUSFaFGFkyJarfs
sIxP93rTp3TvSVn36QV14Ftaod1lbnAUnTb9A1N1iJP0pwiKHSOZzGzKoYmT
YfjRlVosPJtiFVr9pMEUv0afjDG6jL2ZCJczyQo/raROqRgKLOioKryjRMQN
skDYOR+h+ZIhWUOtFcEIAKswYZXPcuou/fH4z8Fp0GhS1aDABZlpz/sxa5KX
LW2j08sUxtL6QjPlpO8MJjEaFOel2xWc1NYdlJW4j7A3tHHpqf57XKRlOLw1
bdcGtjKNDB+OOK1dyYDKwbbQf18lGxX7hQH4PUt/ccPUcl/sO9ZmG9Zfnlf2
ZlGbjnv3OTCpbEsT0Aziiznr6ucylMtaBmbOyxiwLdWt9aWgU5mYGFSMYaIn
jdskM3pxk1hZVz5Epv8vNFgut27q6VDa1Ur2Al1pAquFw3SjbvbnAB8UD/3A
7OsckRmygqpkXNWZcjNFseXwPdk6x7YHRvnVZfkJ/yTSEWdCt1Ys4nqhFG/D
MbYKpAOy0xDOnoBGIusuAyr1yOdrzo/9tW5694jmfuhQ1YRcTUfIzlteNES/
kZY/wtR79KDfMA9yseTo2WOMq/eDcZQGDjdBJivZ3FE1M1svc1mkjxGNlC8I
JpTdPSNB6VRHHvB4+GUSGYaVyzJaxkzaVk9wlzrRkBlQ/O/puACU9vFE9HzE
8GIyAW1snd5fOrcJVJlvqKx6TNaJuzo1GQDlUyWcL8Yj6xsW1NPs9paw1a4w
B/ssYaNNKoox2K01c045zxFQnsdDYoDYaAhEvHcjjPaJqmk33UWdGac39Aa0
dIzIwWqEz9UYNTkScnbABURDi9wPieGkL9KxhD1lBtFFBVsv4QGZE4+BQmnU
n3YbJsjmG5BWN6TV4Oj9bFUYBirN/lzYMIx7oBVLhyypx1GZ+MqKAWBbGcis
a47tsUc8JYMUTuK+rr822vwXY9RTYg5gcprAQxFxgo5TUXFOtTGiRzlBIXP2
P/V2FX4aPFxK8xYq8Lg6OJyGS7Jac/5QMpUvefpqFSWulPnNMS5eRbSOI4QI
DZ+UioDHKz7ks0c8/xPHU6rS8kV32Pz0G9xd64NBrW5ATzQzvbKVNQooSU8S
BI7bOFmVeqIJlD8FufFVU/o31M5nWcqUo+eks/ekYzcMOBdT4gzq6Z2SSoZU
k3Lum1+gGFb7FXYJPCqVZQVIZEXuKXzu2rWSnVfzpQYV+3h5TTkS1KUvyWHt
yA++BLZrVwt/BHioA0oRWHI/tUDgoZEtJk4WtlYqnAllG/WsCILFtBpt9m0o
YQHNISmt3wzy3fwA2SagRuAiT5tgvXHUzVS31rqccwOJLYPTqFJA4iNF14YK
O//ZMfBbK+wxdKLMW+nFgky/tNKgF0ow7foMvL35ikFqJ9gwjfBg4sP40kPA
mjvMayFB5ZXYPvJQHNhNjycVFBIUdJR0mvqa3VCzPyKhDQaa9ultjrJLceXN
tCNlGeWQbT00YihuMm5pirAZ8Eq8bcsE2ahVwYD+vMZyhiwyErBvEi6rg198
OAYBS+uq+urpQ46F1mWCKeo3rDOGffD5bhes/HNPcfhBIiLSiUcwSXQrCbMk
8hRSzWWgPKEfcgaRmhIwa1qiBZ2QoQLN2giWH2qIzVzZkdLO0iBV5eI/ohSi
EYhml6N46ej9BH955erL3TVvVTN18kqJMvMOLwK8A1yZZITkB/fRT9rCuVAX
qYMfeJQGAfYpKPDrdZL8Wb6xMXYByS3yd0fJoGuqreXp5Sr0ZI3FTfukyaYl
2dwqqaxysiKdHnaumVofnM5kfewXrrJNlJ55P7KPxa3x21xcZbMqmNwkMpze
KcGETX1cSD8PwzvydoFC31n8EJfbaD7Jfr6Fnivv1fCJ23wCguCoo4LExkyv
uvX5CBGKpUCtO8ZVD6KjF73GKHMmNhjBnKqRaKokMc27D5j8wKr9/bO0WRqb
8xWUpdKZcGy0BfKPcNcKxB2lIKUfybTkc4OfQ4g2CPL+cqHwlb+/1ATOUAI+
agfhzY9qczmryi7kIc2FkmvaP56udPgQODYqpp/PYTJbUpYBwcL5VerqrN7H
DQ02yLI8iGg5GQv6u6Zn3gGZWUDIYUNJVfhBqUOGx1sD8B/fnWB8JwAh5kks
Hj8nOWflHdoHI0gTjRLGmENZyZTQOxJ3uAmCy1MOxdP06YtKCclA3pUHN2nA
2NiVBOOb4bRRp+Z6KB/QV1r9LdYmhSVLmMTd/HjhRage83mKSqvmY1o2RR/T
DHTWW5gpG6jULIJmm1WEQ754YTBWRthApC4feDRSzqxRieEHKF0RSo9+mLfY
yMGtR2pPb+EaKmevqdK5jSsUk6biCNEZqeUhJ/Qome53XCaPwQJ0qQzo/qzJ
jQ6CMjniRA7ssL+kYs6PahFgStF73vq3wyz2amlqe3SFjP0hK2vIn6kdcVmh
TPiielCmX+7oGH/3wljCz8LFbnh/jh5NshLnBIS1ghkqTOQe/eY5Z+xEJuQj
YSVSlBUAsa61/UzQhvsYLPZXI27TdlZwjphAFQpoK4EM3h9PdoHnblvSFN7m
6TH5TmwqB5fv26TH9OFI/JIJTRXF1fuhfNjiBmGZwGiugfzUV4pR8YN1g9tv
0OG7+xVkA/rVGptMxdji252A3O4GDidNHpMr9C21mwg1Idruofqfj1XLRVmR
EH16SwDXd2NG+s51CpMowQexSw8TuREdnz65faIxFRrHsbO2RX4kE7rRWUDK
m+N1ySNIXw1m5ehg5e3pruyBksaFcpfOBUG85TxzxNl7aNP46VTQSM3zuJ3P
+ouGNnMiqKQCdgPI/fthu8trSyvgmdEUDGLgik5Rb7LjJX0wD8S13iYkhqUn
VMx0JEqYCrwe2uGUr4I6vCyMIDe55PUy7pbL++I+XFlyEdgB4x9Z/lqDL+Ru
O3UuO2rSYjUBPvSnlyPn8DblMwmS1kAogvUyvNjaKfdwlK60wgC0filYRShm
QPl6YGzFsUFWrsBKJG6n9VNfDjJqc5f4NryoDQ9zqICSCQvO+DoTVg5hibTs
sOAY5GZKOobxpN558rZwzR36iFrBWJDpqZWp+U4oxMLPZ13iBrIq+oGS/R9V
cG3CjRc+UpjbK8sksu6HWm0uFfhfrntwhdUzYzGLGHIDzva5i1ILHJyph0au
arLYlNYcA/xDVe+BbGj4kjLeQ3sO0xEoov0j7/lo82M0fdoRipVSF6EzfDPl
LYClC3oTbdqNuxgkPL6o1/Nr2TSPlc+WWQyL0agoRiXI7sXZyYG9F7Pz/nrn
1Agiy9Q+hNlP72Mk0Lj/1p2nBGx0OpI4KpWjALjNovmk+pIwag1nFl8E/3nr
onRyIP/FFOapoVhMIduu+8ZlcEJuCXNVDHGiqN7/yBkBBsMkR5BoYzVkZ9ew
H/liCyWpouCis60BlFDE5MCVAuQz82pmBUaC1Ea7IXRSvKhlWxTwAigj+tU3
EK9nhXqfV16pZri0mZ144K+wcWGVBAO9BTUH4/wFoA/RvTYxDmQBgLbJM+7S
CCu16QuX9cIsb7sQQZ/3kZUWwaWCIe9d/Te9UOLKnQ9+2WwUsV67M6BW+SHy
2in09K2uOZk4Ao6/s1+BsEZ7c22ZZmfbCa7qD0ph6vdoZOWhftx2b2aik6Ek
BZk8ZoSJAy9oDztfFhfOuJv8aSrO6RjkBLduVEkKuWTSRYv0S0vWSFpoPqpD
UFqhpMXOfErDiYPLv+P6jEM7JRrjti91rrvImuGstRNeo3bRPBXpFPnQFUHW
pCgza5NUbvmytUn4QAlC8XsNauXkTSTAfyjaRkvBE8Z7vwhzFljjYEVxCb2u
uXqAyugYAxu4PqAamgj0p5OR3QyDdih/uvQnC4CQbdtEZfTX67Y8sVpvfxqw
q5SqUz59qQv3QNLe3SJVddq43Hliw6l5DxTTNAF3+CAzy2xzBQnxqqklV+wD
i+0kGhY8bdwTGSMk7ziIx7a/i08UmSL7fTfveHfHPamkCY5gMCSsNfOj98Ny
FC9x98d4dlFMg+JDW4taA8ACXDEVqKUy6VI71bcpmpjueRXHxfWdFCJvvQpi
DqulHQ3c3UH8MU5dfIUVN217GjDCW4TziUW5OonNgC3Gc+gMYjXX+O3x3YOF
8XKhXNF0aJK6/DZbL0QYokjlyTCMkrRreGbv0rtC+D9ltT5eO2SjWHEzE4sz
U9yIWG5/agqGPQTe8x2gJr/ma+cWHiwAX36y6XLzKY/nH6r5wYPHtHtvy1WU
6QcNfaXIaDeVqhIQZoGho0Myx8Ub8BBXO0Yuh4/SFAAGjkJMFjJINaAZDT6w
3MoGkdb7qe4MPtkSpKobc9BPjckrnUuBnSbi2E32iYOn88U9+kwcuWVio0oR
o+kc2JUEmyunwgFV4LHI/BNXKdaQCF74aM+Z51wBObXIjyI0LH+ZF02Zva3c
Wb8hKiNrjJ/MdYu4mztUbh2LFJRz7PCf4NfLO2kcbxF7KZrlS9mWvHfwaR7q
gVw3qbwmdlVdGvgW1uwLKKkUXGWIENa4OaNYrjJ3Md8WkweJQdD+TxUUkQYV
f8RDKVwfD5fbMdNQ8qPFnj2Z1FxMfYpxhUjAL/Vn/aaV6gLobswhP30aOOIs
fZfsJFl2V1L5WEe4qPI6m4vrofFOQMPaBsS6dMFiM3OY0Yfm7KvLEmR+sPpC
wULWhC1QyAKjoOCHqyYrssSOKswM1tQsj8cP4kIIoPrV4buf308ZQUO7uatJ
3cRQC0qfrrGDjMbaM6JRHGPLClYyII2FBn3LaW5SKVML9+sygndvW8epufWg
hb1JzbduqOHPtikFS8oT5W/qxIfq12v5lgqXUwpc+fWUszWz9uPSx7hoPGS+
xZlGpYKen38P8tzUwXHDdSAnmfoLtmpdIxuPeOX3KEoq80fEPOasCKpzS69f
OPPD8TVaWzv13KKCX/3Zu3oI04TexcsZ0EcxOMu5sUhqeC3NckPdYqW0NzbG
7WKyHcaNbFtzZ5UV2QhJfM/UwH8U6NAVVhGGXidH7nUaUbtbypKf0MraVj+F
9vLBzJCAAQFFmMyiYihZ4MH3qahdwBDGXDg9v6R8mO9YztZHPXB8aP8wykAE
PWAuarUrNhBd1ojdvwuIQEKJR1PW5mgj+/JIo00cSkqbYwInG8lF0MqLcizn
wHDZvpgeCyvqTq+J3B3ILdFtXHNEI80o5YF/CSB9gXu/Fez4EF0fAuKzQvNn
up7BpjnVpevYNt2enUGGoEvWXfmuSb1JFuAutu0sh5EuIi3k4pJHi3vGyG+P
4G/UwVmpisSwJY7pOg5uRkAc1oHQhrzFsrip4T2mREcoaIlx9nhcEm1j9/g9
StkLj5sTYXApBeYRuiOz5G7mXcbXD+x+EFc9jL4e6bYMySChKWyym0QFi4pu
bWi2mw/TRabtA/alV8Gz210icuAdu4MhyU5ylKRa5jhWr2+IAuODeBcrWN2/
I7c8die5pY/6qiOi++FzG8vL7XLrhbm4fYU/QnWHRjicUuTBCxBSZkGgNBA2
I/dP5t35wdK+uXWfoMO/iqhbkQSXaUpwq7xjHmf54zzU0gSZ5moLn5lc76kM
79maVd7DOKB/s6g5uVR7hcYcwXmERGwGcnangDs/6j5Y+sfP3iFE74VXXgMv
m1zlHK9EwJad49k4GpcVIAfUQQjQjopajAUPGlWpkG2SYU+IeTQRc4TFZ/zQ
FWKnmB2+wvFVI95HsFWFOKVgC8SKZh9vJUWAm6wMvsiRqWpI1T3v9XE1eDTL
VnYaLOIioioU18rVN7F6RHlbzOm9djXeQA9XZbq9MSY2pulR0T2u7YzQTBrP
cbErQHVVNIpVF3HL/+O77zlPBb4Z7vxaaqveqprGoHiiBF/X8yoUzhGT5Qu6
A0+/CmniqTYjZQa8g9ZygxSpYHclsW5ZR1yjdOrL1+np+ECQ4/trEnmpvFkA
OdcztsYN4MObJ0l95BVq4LS2g7q+RgeX6m9TEMVHqbxLTm1ZN2zGuJnLPUY/
Hn+6TJy8BEqDLtoNOXtnPc/tBY7Qg3Bqe2myYU4iFoUMTnDqB/2YHfglUVek
PPwPWdrjQWAV347TnqPhtQJyBaJVjXlLmGaCnbV20pOh/dxtwZ9cXZwOoCEn
xaKs4sbWkoQwz1z3K8i2n1fv5amyRiGS/hf+QlHTFI4mxfYRKZ5edpQzYWRS
Z3hPjf6zYpVcbJX/k5bSHlh/N9dLPQ9hw4hdGRSnftJpImOHQXLuX7IbgGXY
99DCidAY+FK/ecROj/b7c28za6Qkyxw+PVPUxFEACJw4RsEH8Kb2xL5+L2Wn
4bjngMpUk1LwY2ppa5am/5v/dZ3dZG/ZAFdYDKHdGbyiz/VKQuGBmsDztGUB
9PHM+7/bnxFh457R/m07I3ohUT+/ekh1i/0zw0kbeDizH2KavRQhZwRabV2Z
P4u8BeT2/hXFFHTVDbA11eZ4BYsWNw9xKjnyr6jT9XvcChB1/7tvO8zG+3rU
n4Lp7DVEWZNxwTMK78glfB4iRMtSNgj7IXwe8EwRR2lBK4KGs4Erq7Ztji8a
gmkDc+0OfArlTvvd17cfpw7eN9LUVbDFNSymuWi03A3RgOKaFIhAttpI8Fs2
/XSC76uE2sN69UUSDWvDNXOQkPif2i5ANd07AqulgH5mb9ETEMPu0Hqj9p2o
acbw1ZM0jV7XPLbiiVnocprjUG4HFlge7aWbT2uDg3xMjjqa/jon1ZIlV8tQ
nd3w+Vs2gILWL91NnKyPaGTM6avRzKl28Wmn7NGXnlhZgy/6g0quM9UyvqPl
pNHg8BYQxK+FyJpNuEyjDCzfo9JcUmVIuewIKivzsQvB8yhcXVy7wVRXfUD1
fExUOdVXCvgTZRD4DuhQJ9IzCYIZTJCkeFVBnfFR8nnO7v12AzJzo+z9UAV/
hTJ0HPyfxqCO9kMBkBGXQmVfkxXvEOiN6IqtkZuEio0yb2W9cqJ4mmaSEAjZ
BwXN0uH+3MMwKU7KnFeqzMnA8tQRy4tDz3wXm5rTyj7sLeNXn2SZLcaXsNd+
jFm3U8rEXXBjVO+yyAddGKt5AOmC/tOUColRKrYZawT405sPoWNu6RwxzaMq
jLGzM69vIM8fUpVqeFKnnyxObXkRqZIuds5yg8HSXFkFL+E55EWwNd5xe4X1
vchGlZMKEJ6FBIp8lcvDabriBJlEhTPCUk/viuClqn/v12pGxnCeYlCx7tHM
00QvmLbzhug7p2SGTnFqzpsPu5FWN8QjzE2aWzTe9Q5G8NRRR1XPlff3fDJQ
shAfJLhWZhPTcIp1Sfa38zVrqpQ3xNOE9cDTRp32duvbebuy4+8TyLoXyPJx
dVBZzAqKpwNagdc0szT/o4nErD4UWKoqnG5J2CL8rZgo5T7tODAqWWbIvRLN
iyJx1jx8bXmxZR7aNiywb3oPqRK9e4zSwvIWgzLqjXzzapQVp+2AO+2vm72c
FkOXuxJq1tXteyb0rH1AvVhNndBdu8U1T9plm7ppnh2oGf+XA4JLpUs8W1Eq
olkp9WKGi7yd4c09zT+nbcPuPLTvIBKbz1fI7NdbjFMlRFxZagHiJf1weyCx
5nf2Wgz1tTGonu7O/lYYYPVUHygVN3BKYVUW7WBP3rMmxlBnFhLQVIEvdSYe
Q2m45hT0zNCB6RJ9fm7cOqbANWogC+rP3+xnILpampbLngyY7LbsYKHzVx0n
3H4QLFbSkrAjxRE90FX5ZnjKkdIH5PVx8nQAeoBCBUeUbuDadKnQNLff9XU+
5pTn6VFVqaedVBfuML02YtJSCEFobFOJHsy23cBQBe9Ny6aTb0PEpjqDNGVz
12jLPVB6aUSyr5PURKpMTUL2klj3Rrtz4LnU/Pbs7Nu7EqhKmIgJGYb/Vlxl
zyFvhb/TsbqUBdKxBdc6ur2r59EQMzMO1+F4KR+b0KY8qlmXt982PT4+Rpce
mJ6sQKDgzynA774UzZ8YXQoB4yQcfQ1Xxnd85qHCcesTGOxSL4JiZLDX0QyL
PuAm/NSwAjbzcN6Mi+Y5PstlGvGLLqS7BUkdPuYLtdGXX9VTb3o1MpCRaTQj
SWbOi3eis3X+vkYtlF6S3x1fqUaC9ODmgyOz3hIeNbCTD6P7AIlrodjx19ML
sLYF7/9ocaLokLwbEolioaaVd5qxSXlFzMXul1BhyhOsHrGf3lhy/Zh9WfIJ
+eQQWl5UBGHK+iOiDy656/pZGS363GZyOFTi56SwPh+AFYX8fAM2OqvJJe7h
thn+65f3D0O5xI+Ctsl5oCW6lj3dFxjQK9vIynBgA73PJTR2c7h00/wxr06K
tAtbMn62ESb4CdC2PTxNMymauhlyJykfJj4lS1j/+A6ZiLKnPQD+KUqtXiXX
KeryDi3eC2j6JLnwKeK93fuJH6Z/3YPqGcLnXcnKQffL0sEAV9fV+Iy9dQ0k
yK4oeTUjLgZj51FoolALRtrD1qrS/Lcg/syWWwYopV7eDdY4yiSRY3OrmT/U
Of1rrAYl67pCkbmfJ4Q4sRksIyx8mmD094LSzO5MQbOLetjnWqH+VaEHej4Z
cJ9hWLQNGXCF71BkwwMh/0/mDCFVOGiGXB7YEKLCALa+0jwP2zfuZPAbf1Fx
SH/It6d6CEJSa1lrUWY7Cwqd3pDtw2HApUBo8JON/lbipRfOZsorz5Ty7vNr
Gm5gaROd0kxAsIaSVhuKbMOZUpJJ/zcZk/Kj6bckwQDZzzCVZXni76e5Vuw5
nYf7dwf90WmIl8n+MqL+VlEYct/5bTHFhLdIzVFdVnUS51Pxcg3BzWDMKHAq
5w64qKONTiFdED9pJOLvTNQX5nLWXRsHO//FI94GbHnwVTbnZpAl1+vDTcN8
1wrJwN3j0BHtKhuZxjCrwL1JY/2KW51VqN65i9PaYcisshmC79HKQZadRJij
mMgkE1DPghi4K+Zh4gtlkZjWu5d+FPeYRkwACrTaGPXsD3shkOLl2BdPzOdk
28kfpWls/UETGcnlKaj5N9J8huC9T48BDtl8Y2ZqpiQsxVlT0gsogYK4mFLq
soF0ATSEHnwSamCGS1lggIJXAcwUy43/TQ5n0X2yCFRs74A0/J9JuEkldFzM
1mmXaF6Zw+EHK4si3y+8DnC/ODQJ3SmYcT/ubCPOj6YWsT0i+NMtEVWUhj5E
432gb2hwo8n+KbFyyM3mxKiCIEyfjLC6Nlw931CaMFv/pOF4ETU+Es3LrLcF
Mw5U07vJR7X5ULxtDPWTtejyQR43GDYhNXCH47GUDaUyCgfKRErLeVn+HWG+
tjInjCvPUwaHgKjl7ThitCnUTMrol4Eg46HjTuOr3KZ0ktonZphRTY73NMdX
MOAn4oeqZdxIdGVZ3uxCTAqSV3fOq46pMMivWMVwBr7zt1J1o2G5lhH+ipIh
TsqOlOfc6k3Vsr1CrSVJNJM+qHLfWX5/4cRpr4xNmlGx3zd4NH1mzimDoINO
BdATRUFUJiIkuypSHDODdHwFDK+TguwvmAfjxmxCQldp1Ij0bSj3KJ28rDNW
MNAM3Tm9OELk7bWBRYc59/pNdc5DvzpgMDmxjCoYT80EuCPeLJcH3sVSX7QW
3sob2sVvhy6AWDFInjNRh21a+nXA7C+xkaHw79xcqv45VFsF3ZYmSstjEsen
fE5aUP3eIItVgYBJkr3uw8UAeE2Ovtt2Nhv2+uF8jY5yZv7fZR0m9bf3ZKFt
oxknbVokwH/1j2U3kJ/IAkF1Abg97ukC7DHk3Skp4Pzee918zbMXa6bzNVAO
1f3D3Vq1q4eXE1+gMLAuKK1sO2jS3bO0SXkgTDVzLSWrosuQa19IpGRDeHr5
ssf1nf6QG+JeIX3GMalazkz+8Pqtlyniqn2CCgSfZDLf12M5OxMB0rSGGajj
pvoEJdFmUNaeQnjo8EkFhu+OTu0rLcRBhhneLVKjK8J46OyPGCN8pyUFE/hY
9Wz50knPzetbjthZAY9eetvlNfe9lDW9UY9iGjp56JzfjEwpCWX71DnneBj6
OTDD9J2Vg0PGT0GI0lEXOsNcDn371Ef3Igb0wWEP750KFIq3e6GSq8cbkcA1
AJQK39f2/sJEhaLGcAYxCoC4z3FQxaIp4Va1Fbx2vf6/2zOumkN6EpfaHGwT
kPFS9Aph98+qdtbZkdvXHl/x9HL/cCDMwis4i0PO6qyDfZ8amqEMpLgwqGp5
qnX/kt9H77v0DYO6MB8X/fxLHDXvVkRvgn9KdCSI6WSUvhS/081U6y5YHkQ7
V3WcgEi/Q361ZGa1qkxtQdelXdl2TtI8gzAE//Yn2jpS78CJigD6qBXKRaKi
nZdZlHj+JdepoqdKcj0RJXJvXUMnoSwLoifHki63ZKS58FEIIJBxbk1D+DW6
kzUzzfnU6YSa5mY4bV2zE9gvCRAFm1zGK/56z0UOAas802DJ4bQcSj65qmkz
4E5i5cJingUcZsb2ikljl1Zp82RuvMeXMaayuyGCHrVmK4hXg1ZbUNUPkvA5
SFlTnCskVRXmWvjmz/wlkpMzKgGou2Ck2pvklddgr4Fm7/hzGyX/pMiVhu2y
l/+MLYVeol+wzA3BBSu7bYIxjNkSk8h6nOQvP9k6CMyToqn2hYtzAh1LwY4l
DAEtVxuXuco3Qdq0Vx2HjGdhJqmKbQYrDFvx9hJwO0ybRoLYjFoOTCHC6Mhe
UWFtKZOeE2s5ireiSmu9o9JmozKqNz9po4Pn5RzsqNAn94G1qdROouW7jc1a
IGRkRqYZknrcivkYz5fh9Sbal2Tq7YTFmk00dfwt5hlwDH/uwy5WelCh793g
rpIjv/OqaTDevbpqcy1kP2ZNZkJ795BD1pFdH8pMGLUxrTRnh/rt7TaBxQlo
cfb0dS5A3msfDtnR4DLGeDpRWH4RlJPT/NErSgx7uNmzAjGHA7PMrdBcTNhp
MIsD6ErEjvhJs5LuNFBBxxiectjPWdUm6aSVwFwwiaOX3AG0IlS68wZP4yh6
Q69gf5YeuQ+3RwPcR2pZL6ObpwG/VqHlUdJlUV8vtZ1C1uMt50kEi041EVwS
t5XwEuN/8Ky1zaIAn0bH8SXf7y0p7etcBMOTlNkn//QnV1zyCqJEX8j+1yWp
38jZaWp6ov/2sgw/Ebz0N7MbygdHCEFYtxt02S1D4grE9tB1aPp1lDBCIYI5
pUiNdXkvSPnLiDGBPXxkB5dzbM7wztrNq87alJW2G1FPbNlJeH2UZwZmbSGl
E92TrvwMpkDEXRAY2XSoISn5cfAGM0Y+zvZS53xOb3BrfdnTveHGRUEtREws
Wq4Sb20GksBfzbrje7/IZXHEWHAUwwgy/WWUvApm81LORoN2EvA5rPLCAixk
nKuMyHcY6BrgKF6Ur8MJvRPWthydIoo1HrxEwTCnUJsLCxFeLe8CesxmKBF9
Cfiv/intpmsaqnYaYVX6YB10JkOwwFZP7C0nmhiJN017CsXjVC2Vv78nnY77
CHITr/VJKYGhVX49efZglzlkACftiSYhIHUmjDmB8/W47w2m3mZs5r0MdQzN
9v1Y2zfE0Mlrpm6mfvFVuSw0B7Qvq4exU9Om/Oewb21XZ3JBuasePiZPSgH/
WImtc5Bye/J2cr5LPfqxaoB2YEwQqPUE937r70R2HftTd9x2tnSFn65HvjfL
aaehGI6Ibw/L9z4yXvPxdiUGyh+9GTlzEjvefFU0T2p7/eND7sDEYe2UaqVZ
kB1VwNxjzjjY7sjAh0eZTywh44fsmg9pwbPNaoSPVkN3KGMF5bT4TkyXsdyt
+FpngKxyuzhVtYXzKBTRm29hiqX6sl3JJnuwsfB2BumJoFePitvrJj3pp6L4
BfSMHVTWWE5ndF7KnnAbCav5CnkgPFkEf/Ee/z7m1AnR2FNw510Lt19OFTYm
a4MISE1RLh5ZKcORD4/w9B7Dhu08kWRV5rKbrv24vQpe4yeZvaRpTbKAagHw
cNqaP43GXhbpy4NjLPnL9HTaQ67Hi9pMsJIF0zuVZhj8JMBr8WZgqg8iJ7Ly
kGWrcvxvKklNLaiKp26C732BYJDFXh7tL52ls5Et+Sy+JCf+MlFeMZkirCIT
x5PBkCaFqJtSqj6xXNX1lbdYwSMjK+fW28oUl8T4d70sl6dSfcvGyg5I5q13
+wQSemT6jiH+9hr7LW70fsXEB+LirhVnFwxWQnE/qoUDK0yaYWhvFZ4BgLPp
r9XtEfIClJxC9/7KjeuMBx6zt7HyI/T7Yfhe3yVLrACsc0/TFRAxvWQN3Std
gs1jhgXEfNvrDet96RHu3HeNjcTtJ+40zuOwxdFy11GcQ0dKXocd8+FVMOdU
be1zUwTppxwFFX5DSLSdrmYm5FU3W/TVDEYunu1KOljXD/7UuadquHYTAvfl
HY5mETO/KH8+B8OmWYKF0F1Zc4Rf+OrbZ0rUNWKiiVJseohwDf+XyJmpjKiC
UIO79JDiSzUl+vB9IS4NcIdO0lk9DEafM/hu60DZL4p4bY0fegwTrHzDcjXk
g7K9bUmaODpu/yikFDCfwEimJfpr9drL5uT2k0JPY5Y7WkP5hTcmkr2O9yaY
X/EIiXOPKx8x8KYdFSn9oHOANRlY9Q9uOlwyabvpxfd4rTPOgjEL9jXOh7er
Eae6rleuxwwcXplToEwHYIu2U+d9P8964DkeY5xrrb5rUWl7g982/xcWWj9y
mbGkmaBY7HIhwfLxJ3OBCt/EFrtjDaSQVRfuIiwj0Mx78UnM9+Q4OuI5zZkR
VCWpjDD7N/Vb/HztM646t+Xn1E7tdFDsuGuO7LTeriwukuZCcRRDyASnQ2kG
mD1ee+8F7Pvg0m2pvP9Ff0cgJIgjX/gdrlCrHLgOAPKFJGFuqu4GfIEf84ls
/dUyZv7pQ9GY1Jytnsk5ioMxO7Kb9B1G/LRVzHFfAIrnVSB23N45YhsfHTlx
j7U/0QCoLfoxU47Cp0/FsRdImfUV+gwgrP3TKf6Nvp6AzQcR0dQc61r73WqI
DJv4UI66kaH0cnSu0YiYdizLD45firbs8nPesvys/BEtxLG7KJ8Ejw6D9MX3
eVIpWG8pSJxnkQm+DfANeACx8Qc5u0hjFDtKRlELqToAbz+YSKYPoxAisNl0
CKmga9tsKDpcTLzsny6htnywXK5AXP9oXAZUAUmS+djG2dSAlBQ0flcCl0Gs
koOT8vbm0fFJCw+4vgnteIMZeXYEcbqaGiQcSelWjbCsgVDKVbg/ve7tldsi
u45Ve7uW1JGL2WG0/SzmKaolNqfiEJm9xl314/f2zov/3W2KKtf5LbrfzJRF
TP0mKvdIBnSn8ohFRxnAhln1jEjd1xw3tt2V62RNs4GgrQFvhpObskTsm5Hd
CYrQP5+VJUb3zUSRWCi+B2gfPio88+qCZ3R137QeyWDMx6DplrLPMkN6GJ90
dThKJX8m8rVYTqMxtimnObPyO3/ulHurbnqAv9MRdDh/6t8KpkWreo+exNGH
mdb/85gzbbl565IMOjgnQRypFHBgvCX26gTARHyRWwfnidAAav2CbOOeaPhp
/FdnpHWbR6rHVslQxnp3uaZGPxmjF6wOHRJZej2t+tRl5H1/UpIbwZ5DMF3u
F8MMgU2J+xIUFQp0FVl8mcGffeZ/+gFSH2VXvBre2R4IPVj9hGAamcytHxJD
zYBxyoykiBo65OGBBUTmrs1Do47nmjoO90ZWid0eRBLNfkOqs5vvdzg7C8co
JQ6ypHotjLD4TFzssnjXqJl4je8/OBA50N8Y/5EbVVkhyNiCQ56RmvlRj+Tx
zD+H/XOt9n9OkLNgX1eQAfV/ZDu+jJHEnJE/CEuArAId7Cqtox/pFkY8Tv1S
wob8RH/vF7QTlfhoseYcjWpyNzohTI4B2g1komimFUBU/P7AZIAj/mbPOKue
JBYn7hFoUm9AJwnwBSJWGRtOrYrgCLfzjk2TUs7kKVdzgkU13nBtGP2XgpeT
95kBU63Lj66LXMOgF5zOFicFsFs12Wdwb/ETDAWgWQcQXmKqRHBihx/bg+zU
d1OATa8mXi54dSDgU/cp+1HW1phQ6Ew8Ho/dSF70wsJK216XDvl+FPgMiZXa
N800wKPUMu2c3pyjlvEUFI0lAQg8Ega2DM9YUzuqHVbOOTPzq76vuNeNehrm
mMy3oz+NINpMqe66W+VBfCgUbHdM/mSSuQUWYMdUlvY7GOR/IUYjywPk3bCK
cfTBxgSjxLs4mHi0q3ubPY6PH2f3LCB0XgAOD328RmARmKwh8wdEeZ5aJC1I
5dluBgXQyDEP72qXrf1cvjYqd6YYMP1E5y6viDF2fLNjOeEsi9y7+pWsKfsu
PF/Mip2LKKc3OhISItEOyqvVazCAwKD/JzoklOW8l99SCvNQix9mo8y4mViR
eZJRTN/ALWEoysnjDNmF0b50gNWtYfg2cyN2Dp+PFyvFJE/CaFTsOQ9qsPOz
n4dYrmu6w/bxdtXwvqFKPup2LFzq1sF+ofuspnf7kksRcYmyCMNs80y3JyPk
oR5aoJUtLuR2zPMvi4sINmu+bOdwJznlD2NfZiEWQK/8+PH5LZi1kd/HYtfw
8YhTC3KLvprGgSQCkYNeZpjJn9jDtD5PFlBSr4Oe38ze0KigEEwHIMiziXuI
xcrYcN1vVmxanZMX4TXFjMG81tolVWyzINEwGxiWSA185bGLdKosRH7rYdPx
MexaOWFNWaXSZl4rsWAodC5frkPU31U/ZmZUIW7KkccioRzK7JyL7CtZGMpp
kT9u6iMqa0CYhuoT469kANNxuhKFHp6NR4IjdUynThpT3OGqd106uvpDAkqW
JuA7uge2GRsXL9zyZx6TEUEODN67Vn/k3tlV1P/XeLSgzZ9WnswdiyiP7hK+
S3pfbxOPUaGseZkfKR82Gfei8ryvfNStLWfuoo+5Aooov0clWhChv8UdZn+2
Fl0pIzwyG+46Nz03z/2cfxxPMsnBpvpDYdLegAjNpKHiHomhXADYF6kOOzqQ
ppq1E9HHSwV8pS5czc7hstyzM4YijinWU3SAL/kOtm4DdzsO4GEJ8I3xSpjz
D7c7fvdUq1LbeWW8uKtk7hVmEm6gwWOpMLBZikuKAjta28GZ+fjd4semV3H5
hMzoz3hAlOEOzwW2ZlNG6EigkWcIoPdmI62q/Sdtmzg+QE5sWtiXbvzGlJhD
lgcpOzQqxxiXTh6mkjtf26uR4fdVdls/7Tv+71FrcQocy1hSOUeb/UWwJuw5
MPg9Q8kfYSYdhMzKwIvYITEovB1n0mqav7A0I7UFyMZrLrauSLGofhYMwok6
SO8EdyYgUpSgxTwvQyxyz5QI178VGV+D1RnH14v9Y2c++E7lnY2dz27n7/uH
b/BahbEA4JEC1V+Kp6OnUrl1wQ/8kIdG9J3NMWhQ8RVlFu1mG8vTK0wHU1hL
uvG4AE8n4sjAcIZQT1djetXGniYtxSgGVUQWEBKDQOqfA30rsaD4rrVrI1HO
vMtuNr7XHO3iAMQCP5vGoyPzXyBqyj2mrRb2oQV63XvVZma/mR0n5mydZYNi
x8MSXmcVZxyQsVoOx/373SMsWmVbbbejwwHEqPTPZLd/zzu4VL4d3y0eXOlg
Ecs5nDaPr1Og1a4MtlUjrN+ZsoliPGDkIwiEuWv70AjTlmkMYAZdlNnOkxky
gj1ZgiqNvNSSGXfw4LOGXTOK4Cuor5Sc9meKOXEG3jGr1A0i28VbKFdgn/X/
RvymWcmO+q83gdxSvBimfsHiM2EN/MoxHeWdBtwcuteKCBKfXUq5QuPS8fGp
beOhswUcnpsunWGRWxJGsnftHAcHc34MYx4+UhsacyiOt3a+v1Ko5EjgmP3B
59wNez17UvDVbVdszv9X46vilNKlzXcXf8QkrNb3NxCy4XAHYeyM6zRowIqx
VchqAutvaDWOSxkgHvRwhdDS5ZIgK+AP1B5XLeBqtus6+2hQABOCOpb4sq5L
Zd4oCMbOvpzO3VNf/I6przuhcdN9QcAnzwc5Cl3wjyhbE92a1Gqb82lDmfd0
uD42vCTDUvq4GeObtbiW6xZmlH4OAmSSlfX/+MN5LJxvNiZSoaACBwXXml/+
zM7EoLkBi2qnvd3+33JIiORAYqUHGCDdNIl+ScCjtHVJr6UJOPPJLP6YQKN2
iehNuFsj/9ACzYayfw9aVHnBgZj7B/7a/mjL11w/VqkeINMs/EYiR8iU6dIs
3aKViewNfpxH3H1G7rZQRtuYC2UU+IMH52suhhBbEsbJJowyZnt4JmEf6LAV
qG4nV5+S6ydqqhqVa6aocYSDFgo2vR7fMBmWyfj/z0O4ppMR7XfbRy3N4+Lx
99IgEo/Z+RvKXZDuAlj146cuv/ATD7wyNRkW80q7JXZObl8SpUtQJJ8WrsNU
FGSzCZ+hdokZiPtUSqPvyz6NDeljJo2OLNtUdIz3cBci5S8IxXCELUJo8OI+
jRAjGaedMWoupq/q2fR/rA48VILOkIf1UeJft5MmRjLOXkTNCnHMpD7wzYsq
jewiN5m9owK00Dc29E8m6OStAOm3jRDxBCqVxxYwO1wfQtGkK0yxkSuYCtsd
xQqlhnZT99nS4WMw4kR4QeFQjND4rkRIsiVLBshLrINI87cKzt/fhfJ+k81A
fZtmT4oMHEaMFtiTeJRPSMZBuLWfKWtTi6Y3hJ1ZZCo8WET4/ktBndfdnxUd
epuA8aM4jPtew84XZCVgUE0zzO2H5HrvB3CBt0534t7rsw2GOHX1tB+3g3yl
WdiUbSlHzzDnYmhBfWGmXragfB+WkwR/idxDDx0lGFgWRxkaBdMHCjZmRGC/
pEsaWMao1luzfy0WYpWt93N3g9xq23LM6s+d7Nm/ZCoYHyWmbmZITGxhXXkp
PxqWED1YFu2Db4fjDS8DGWrbwZ5yyS7QhMdNhrfVaJO5O6QocnqeS9PoD1rS
+pwu4eXvNerKXcPvtfcn4oE8qdfgrJ/VR1DykT/QutBeXn96gD3WeK3B/zJz
8n/odTvZcuUEzwh8zXJRQNdXNUdWD5s4goSYRZNfl9cQ5KbwM4LiKChlM8c/
LUYLQeMocl8FER9/1wtuXZzcwlJ55I9srTE3OcCv8u3BxMyzmsAbmVT3Zg4S
TRZCjJF6DhwQbbZnAz5FFFJmsAk+zcmIWFK3CCKIxNEvytwEv+GHJQCLQsKF
Qwt6qpYnO8f69MEyEjrym9s4ISz0l5aY19FyKtQEAvUsZvjoe8QPmGhkerwL
dOC0+J9x8Pr7rypl9mLsztDrXgUMmTfrXx66InyMXwBZN13nb7M2/WYxL7v2
CmErMd7TAqjx/2D6DMFCLFgXkI2vSFY7bYYpJIZsbwFwVtvLbaSC8fQHc+H5
XZRcDPDaPfrB6AAu5QBIdBY62qxQoomtzC+VzK3wplh5wkD3CK9fZqjv7Wwz
+xn+UvK1aKy04XEWKFePeOCECU8GbRaVIBDoMg4pLjBEMcVNBFC8NO0cSe5u
1RwAELzjGA5yz5uoYQhkf+Oxoqr9H17JgQmrxFG0UsNHOfORIWyKRHnLHLTT
2CxDeCH4BcXJX1WGKQTKacSWOl4leNfcCmGSPun1boGMxk2Aa1Vwo4TV7tnj
FBzlI3S2zxYQkmq2K3lrKLIKYRf50yHdzPzO/1Z1LWQUFy92yYvQm7tBkDsA
HfAargV592OuHcaSJhFcsuXcudwWv+hVmHSnxf9VCSR/dUgIK6wmk9GmrMes
fFWa6FkHLLlOZePJyqnBIKDuv60enSTfmYKKYqyR+4ytvRz7LMv6FiC1YX2a
qSA3XNLFHozXLn1OnFnE2u7mO2GnKSp6fsL2IYRORBCGWvTDy2FX973y9UYP
+qLYRX3IZg9mfJUGs94QJF+PoCYA6NXaRzYXdfPz7CuA/UJH2ga8Ja1k3uTs
ju4AFdRgEc1L8+SMjXq0sDf4TCSKZBEXwceeYL66ZmljCw0qRJRRX/VXkgCx
R4T8I4NxOzuiZHVXIVQw7Of2FChFWl1fjgvACf94+mVHdayWpXBGHBfdkz8B
UEg7sZO39543yyd7r7H+lXSZk/BUXOC+b8ZLS8SI8zUc7R3DVxr3Z4ZEcSEm
JU8Ham7bU1CCcThEIfSHHE1wGt917lZVLNYt5J/7NcluHNhQY0soWK9xHhXl
zYRqb4zMdZS6iaw7Lc7v8mnFmdDufUy5RCUthXXU2BhQDKqz3XDxmCbR9CX4
O6C6+Vj7bO8rSoMds4UmdFElpVpKDCAmsPikuYiKdaEKaA5bmLrl64TUR+lm
DRVmfy5H1h6oYMxSOkBfg8/R1IrJdTk/dHZ46Rq4Vr6R+7MYfLeiQ0VN+Pox
/sapHYww+XBn6JmnkSaZYQ5/qbyfzr7y9OcrENcpp9uHXD5lhP2mugEYjoJZ
BztmT9DS7k934PayMJhIY0PJXq0T5x63SYm1Gn0qdyLJybJ+h1GTVfNijb2P
tsurREuW7s3UDtlYp2hovn8MhjlthetCSztT4SnlhEiVOszZMOYvnMC8QsUC
mD+RH+XPOMg6uqY/9RWMAus/yXf9CjdF2IoAnEMpSdEl+LT1yOMxhCGVpMQS
ctQeqFfquhmXmUzPyrDiwT7oBRdIBw52JBXW1xbUAKFd+5Ah7w26MCn4HgGP
ICoyCvWTbJE9AtfxNZDE8+1ihOMGsqTqh/7OPIhta+du1SgBPd2REq3IFtLu
mBN0A7vXSjS0G6Z71pB3jX5HbVKGIRXBFB/qq1tkJVExPDM/TiPEDTshNtjb
CvpZRBO8WsXycR2r3ezrOSTsCbdHPu8S27ArDOfZIy58W+Hhlqa4m+OoGXRp
WibE538d25L8ZDECcQCJ0Kf3k0EGcFVMX+QILDBeXbUwosXT/hEovMH2Ys6b
xNp2tSaelPPSccFDHvC2MDd6ZGPzw828O+C/9cqRfod8LLABWNRlNOtkEzQv
Ca8mltrMQRlrRVaI4dYte/CQPhxx9s+5OyJ8RPPBJWUQqDAmcrN6R89G27WB
MIXP70Ai5BGXK3j29QcBd8loqXVqg2iYuSI161gS2WEnEeFWrhpDi2G1l2wn
vwLDZ3TVAkRIYRhimmZJ8u3cr4FTDPKN3EX6WJQ8efCsiPJ+Qenajrmqw5lG
YMP0v2Fr3hGtxJZU2Urc0NSEMQc9sBRe7DYvI6XfFtFO+JBN5RAA9RzeXQpC
J1xeXC0y3YHfimd+LiZ5exS9ojsxffFFW9TNMKrcXik7Yh+3DArcK/fRxzfD
Ho5++bWy1Ktbcd991S1Af6LKsO1qd8B/Ks2jLJBpy9C/VoupBcFCUTjGVEcI
wPgfEOrE86RbmvJ36zUvcA1SCQEyRw1T9kVIssTpw4a0SLqJd+1IGlrmhLln
LgGeYp4jg0Qk8fAQehI+qXrR1ru9NiF0qdqcRqNDmpF48a5PUvY72qkRuo9s
9OEwoKboNBXzw/Xh7/lKMJeykEbLdH2QhlA7uNM99qmneZ9j0dZJIiA4ZJbb
d5yvjB8flGJx1GuXtqfiGfYXeiVMSltlwZYCEKJTP59kYkEsfuZFRgSvJxjc
1BvvGRuCXbzlcI7dBJmxT5/P0E9m2EeBWjeQdrAmnJ6D+BKL2cScytWEEl7C
iaOTNxSALnUizY1S0W56pbdbKQwCxZZxzX/omH5tJ0QYuUe7uRGJMScODvYV
AdNkCe7M0mggaJdCQugnh8wwadBaH0aamzwH+YDFPMvYlKRHlXvdbatbN2dZ
jSk2QO3xCVwHAzBAql/GNwx4YrN44WJKh8XkNps2JsHH+YE8cuhAgK6jAoLD
h+fWdlp3+RIw702vXPex647h5rtxHDC+CHP06x0m1cWxtQl/YFSx/Kmi9di3
hmL8WRbF2uoM3szwMfdfww/TXlpXPUotoGO27ySYpreEDmrsc7rtxa8UXDD8
lFyrDXbQFpcvUjG82DDn51Ct5ZFHA2Pro8DSt3r2fysbWgv4HHMzQO+zBw9y
RNajL1cvYq8t0pczH5NS1JPhFXDUdA3/RWO9mhyARTkNlO+Jz7TCDr+Ng31M
bmYvAKpXWvTHQ1z8dd/R57d5VKavIfkdcCPviZr+ZSAM3POSb0lIVHH8N4Ur
l/4Mks6qOYL/z+hdtGuLr8v4AzZvMUCzA237dXuANP1bYiF6RjltOCTbwkLC
/C3WbwP8PXlgr9rZUzoQ60oVjz7ZHIUTeiQxC3WVO6zO6X9z7YCo01oOyuOx
XcLfUFkqcvpEjTZmoVeVh7mbrF64oe4RsLLaBi8+zGXkQamBj31j51Lwao/0
ADcMIX7Qos4mIcLXbsHfmjE3//viuUIEx09YMsEXf4xtwCxDyvPv0klUMcyS
kUccny8mi3qeE1p+jH6TkiDGIn3hCkFXQKNUbchiQfjcoP2NyXDbClHgLvwC
WdTH5p7N5JT93IkmhdXQeaYTx1HL3amDxIFEDhxCPImu7rIrS+PTr8RAzurm
p9lWoHcfiYWYE3zzLxcU8eBmYNzZPzffpbwQ6M4cTPex7pVz+GhZyMyPKF7p
LPz2fRSKpU3Yt3+8z8o1B/FLs979yavCMfIWacqY3gVVsPswkvAoxJ9OE/Mf
zIYg6u4azj4/V7OUcGko2WbXQnjwO67F0YzNrNoRmvGrVAp3HkLA1KoVjfwM
FoUFTnbuJ5OzKl7PbUUtUByPV+D1kU8480MLnHlhJh/Ow+ZDvgfVgeJFalm+
jvpKVRZHkZ0yvsW5FxJaRa5uuBAEsvSAFj30N7LDWy8ldHeaq99/h9tZhzCx
bHtaLzhkrtJbxWdKc/JoZ1XF3d0XJdDRekqCJCalLp+uxV6T5Hrqy27MkzOp
3B5MBmJiG+TRUTAm3HfBhJ4UdAgVfvjC/81NDmF0eQjZt91mdPUfnR99GlZv
WJg2ipNtHPRiSIdDXSPCMN8guMrRKcMJ1ayT3hs09y9ABGv+ptgX2iCr4703
fSnXrtaORcIehd8ZIpTDueG/lgdrVy/e7BKHSdE1dZEyaeSjF8KrgkpSM2g7
SyksKkjK1aMQAE48yQMwowweZED8s68BP+MTWrtd1/rDA+h+nruFvlQnOS74
E8BSxiWgHzZmiNJKwM3gvp+cvYMr6FomC9rTICXJGBQdv/AV95zrYmeEerRR
/69XNiFUar3jmrNw4+p2HbjEk2MGhh6eYhGUAC8HefGDuIpfVqQP26hYrTQr
eJTNo1y9Yj2XUNFdvf1aQTQsjK68O8i1asD/mvH6KYbDdSrYyCBonGStblql
ewtpafCk7e9qhKqgy2EHEQdY0qgGidG1SwwPdOJUSZXwXxTwKBp3Sa/0O83h
AUxqaeTVBtoT62AD/wXFrhUnfAP9AadCO/W1QWoLhwzJYw9p2tFi98MXSy0r
02vdaDNHYb/+5gLE5L9sB/NrTERUOuXlyTAf725rwTe2JnKH9ET5va2336+C
cMie/EzDLXjJAMxHyAJwc45t1gnkS21ty2Kub8xwUh0aE9gUpUeny+3pFkfj
yYnGL8ZVHKLiBeUlJjP4OUGA0YkHCYjQ7x8NXosX7KSiLIKoSu3AjSJEGyS4
QkyvnybbxHjsDd567NY7abDaNwMSwHdHiBCEiyj55vWERts5xGYeIFO8xm4w
h8z0rzee8nxzS1A3zAVLtd88rF82uU6qhnEPC/QLxYLr6zdFIMABY1IZELC8
VjTPaM1u5USJpbprcQnYHTjWEub36eqaxb7baVUW2oUqyi9xPMFUz5vO9nYU
OKvVpx/KCZNjezY6Yq2WWqINCc2NuK4ysZrJ5OJgLPeG7q14Bb8b4/7+OaIQ
tR11J60HxkFYbs7CLOvS7M1/5oa/L0C4WmgaIdgYz26bRDcOmG/55fQejvft
D6oBdzmyhCrjUb2sjCixXNmbJzYmgibSt5HzlywYdzZMm/Iro4g309GWJ9JH
PpuiY0ibzpJFMImgAES8VnA3oQNZTfoolMfH9Vy+esmndboIMXpwOVxOwbRX
oRK7CsLn8mvXrCjGK2ocvBUpDBx6IGas8/lyHkD4hkP9AViOohmZMdxD++bg
QXEkV1ly+BjLcgKXwlQVUqY/95/YCFlLu04PqNOMDHHAfoE9sGpR0BFoWOih
i8NeO49IAKOaQNyu2iFZYphVzXhBje9l9yQKE/W8vnHGxcw1RAVkbR8n2Dxw
oFXmNZ5jxPCZ8vHvotgudvqZgzu4zcVsWNpetkWSanZCqNdLzKbrm2oTX/RK
EAMngJioZO0hqz9JKeZoGd77JqG7zRkVc3mBbKdObxaO3WvmHhdSmwTirZ6s
QmZoWVg7Cvjv/R7trGXUuoJ2MdBb24PFlu/BxjeRhi8YXFBklGhEtC2YyLkI
gpEbjHOegp7A4ITcMSp+56aetn+gFOHNTcqG9viBSVhJNJwvOwiycPkXqL8u
6oAjviC61kryWs03XUKoJUzFWUJWUTfl/ps54SxDLXzvCjWez5lbK2jBRpie
2fYJO69Xc250ujjqSqbIBGvXcW/RPmRKvGNehFZaLlixIRS0tjSs3szbhOPF
NbhlFGKuLTwnzkRoOdN3FTjOIEkSppesOTUor99sXX806j7ughRPy8bTMC+n
SGvnKUggAvQXg7DCSdNE0iCS2HzXXIzkIGerq4orRpES5+tk/vMvHhoqJAvo
ClRVnorN7BtZnZGb0D8mMow7SwH6H1nkIfyeDILRrk/cwyeH/g9erVZFQSb8
UuWYSwktts7YGc5rfGFxtE9k9WjYi0A90ovj9onrP1S6uatgiWvvS5VqhxEF
xKatziPEwQTUIOkBPlJ1D7w5yUpsz4DezLviTcKQpsu+0k1s8NBLRFx/zLah
SoDuC9qPE+bdI9h75JJQOKvRYCMsfPF5MyHWYU94iLr95bM5C15ONipKQUIz
6/dTkukDtPD0BO+0rX/Vyo/yXHoRtFI/CXFym7mlM29g6J2tMK9+FHsCYnyR
CXIx9xzgyzG7sdgpAT8D2yeXrD0HAt2wbG3X5L/j0Id4n9BIV12hxvUUEdX0
kRxUbiS75uWGuZ2Httq8wTsaiBNNBJMJbtsRwIDtME7MMWS2kKQyhsxsVWv5
dh9Sd3/EsVaNLrlHeLM2dgBRfTMZJhJM+MauCM86RlYISoDWqj3LBg3TNErt
zKfoz4AMxIGnwcovmYj32jLRtnrFET7yVGr2Bb105IkJYBDJdgfDt0wdacBR
63tBhhCJ/DUCWGx1m+qNSqWQf13spxX5JYZS53em2KdgGjBoWVp0E8iSFEqx
6/qJLhqLb4XaZPqAoPmZeiuqYMVl+uutaEHUdyp7LsrgGV7ybUQjeP8nVuDX
WReJ+v4NLwYtK0GHAOEzizP1f2uKEfmgAjBz97V5x2FbL1aUeKSfHBs2KNeU
glNOPqkLlEyGEBXNq3ZUWKoqpiv2VZCnyFKnmNRUDw5J9G5SIJFUA73cF2cL
JZBm8cC7hoeI54SO23YLCXFPICzFj/aez9Q0co9zyUF9v4Z8ag1SuqLNW3Qp
IZMA9URgpR2IKJg8/wklY7TmFBfEI2lmRxWAKO1qGQX7qy5nSSI5/FaG13Ab
wFK7ZklNJdCMg6futF2oLQ1rutkuy1yulSsj/uppUM/gmY8RxAddyIBHvVMJ
e8ZyzHdswLcrdVykwRNqtrFhPfbDvOjxoIYKyzpxh9D1HEaeIh1UkYL8D4HG
5dy7Br3rV13WVANc4wRuyxbFEK13Rp5suZusoDvd5/JbpPfv5bTS7aHP90w1
BjO9Src8G+CdQp1LpSTrwdoo7J0O/jOAk9jYkvdJpKwJa+Kz/Ie/8GcJFjhJ
7eEssTX/fJOQi/LLzGwBYf0CH35N5bJdJuJO0Omu9Gt3TWyQDk1tIVL22cq0
6yHl+M1HpCetF7aI9HxEN3fxp+0PQuDbA1c2ZBBQ+JYR9JG6YpWoXPYVT9w8
kkisHDnt+M8w0U9dcdu8OsMbw63RdcupuZzWPaDSTfRsszJvTD+csvjW7c23
AugosW/9E2IgeNfpwlC6vuoRndBGWAViIZWhsjnRc/kN7+TXrG9qzzKvKPNH
YO7RUdCBs3WzzANMG6ReMKW0lcrSymqpvXnZhGV5cIloUFY9lmwH0/m+TMuD
3gmM8xpdscBxXJXCNyGcrTDOtCUQ4dzqYhO0AArCiszCxmmSeZ2T1QRUuboq
lE2nRJHHO14BIjKLdLixLFyLLLrAQdKkndeV0lCJHJ2N0UvVNN1kj75xoqKM
PF9YtYC8e7YIeaovJJ2AZgPcCwTHUVYa0EC0bvGnZrU6e5fi+pvafnCoZSOR
z4n+dCHNz5yB3sOuDVYCFSWicCqHqVibFmJr3Jc4MQGwlonuxEDaaChD8d24
vZ6xrk7ktNIrokpFUs/nqxHGoXQr5jP7XNlxS7xiCFONQorslAdNPLi84RlF
rrIyFqIO7YkzFaLVLOthP2/MKHnHw8mrv7T6DgKeuVb9Pcno1eFFW66PHoFO
gJFDEJlrgYqLyOYQYwkJj76pyDA2phVOB4WIuXy/hYdrm01cm3O1+CE2K0Fj
uDa4OclL2hp/v/TT1ffZoQCuGSuoKHP8fxQrMz6KfpszLfflWCEDR1Ev/Lf2
Bc+SNKlQh2WBNuFHP+MajLHUjygdjHN0OZBcUcoNvpKBu8wOBOC3dZo3IwRo
KKujWYgILyyEO10ipx3lGG1BJT4AQsPUSqMEvF2yrjSfFOAMefeOwnfFcrIC
ZR+cu9Hh05SuMwEJM2aP8OGvYsyVKRdqks6RfBPto+g54eVKp3tyzEBjbWjh
nFAJZO08EeGcoGMTnDg+fhBAlErCLgRX1gtkH6tHsjxGYmQ14J03ogQQ+g4W
btfmnNqOBPiR6ZmaTpdXSKpSPeAExfiPgZuDLm6n0gZKOJjSdI/hm5iT9I7D
cXoFE62I9RNiN4LyEPNW2IYOohbfqikzOTBIEpGUc3TOtK27XO2smWqXO1kS
GYsGBCvtGM0ZoN4cghUg4m0HGTAcb1VrCfqt/pagblpEX2IlR30ePKRUBYzO
rByaC9M5S7XNZuuZxRe7sNZHO1Z3Tfd2V210cPJ86Zling5kwM5ppJZNb8Dr
A14M7ULuj4ObDTVaK2q9ri44DHcrFQLkDvoKn17+cjQpMIDU4iRVBJgT9M68
OaX0h0oUv4rjA0SXgOUdBWX0SZN7aayFn59Ubm0UEigULrM/sLCGVcLIkOg4
MMOOYiMDh/giTS5OQ50Yu1I5cal6ZT7n8zaHqfrNb03WXPO6YOxoaYsv8sp/
+PzaBpr+LvyrwkH3u6clUFOmP5L4ZXxrWMwjrEImFISE29qFTdjh180HRKDT
AskIq0R1i4gNQ1RV25JrzjriNAoZ1vm1rZHkvAvPbINRFAUUJgZIaVX5mEjD
N7lzBtuZimkZbSZcN4IsnJXzATlIdH8poYbgkLwbs7mn3Kvy7WyDZnhergDm
L89jFiyt9VEfITDTvXERg4Xr8FljQ1X6NyyOYI6lmECPVuOrsS9YwmVtA01i
ehKQw1ZvtvAm99OFBY1feQrjVDqYiJ+gt7QZ3mVk9MS1HzO5aLQF4WxPNBuD
RowDwCsCylXZlK69DjIbUQpOk4UigqjrScx9HNQxtPsdhvzI82JPUsnXJrL/
jioXT5iqaSD8FproFPWgUHnujzcn62rl6gswZQWdD8SqwGL15S+rmIMwti4q
oIcdVZ285fImbEo6Kafl8KJYeO3hBSzO3p7wP5FOcPfqlCO4oKOCPtaL5vwA
2K7wgQ0QSB4L0ka1hO5WG1h4WbmzWLgkfrG9L86EsAKgkSvLcTB3B8I3mbEl
K+6DN9QsZqnB238SJVwth4iMyVXgEMnH9LgzpqfMymIyQW8WCLlxTIk5Vcf0
b4vbZDDJ6gZnKid5aEbJHgQ6EskCzeVvE0cXE9B/ilJVHpSBdwBkqt3dtNvy
OE4lt3cM23oMI1HCGWSuCHQmav4R7qz7hLZbTrYVONnJLAESfU8JKn2zGpa2
ma1NRrrHI4sY/oVmWwIRMwX7PBzP+nq+x4NQrI/M3m+Bh44bchzesSJMQs6I
xgaEzu4syv674Opr1rwVeW7qXwnQ11hh4Q8zhBr8nJrfG6rNfMIBrbShDNKY
qE4ds8v+PFunQzP11kcq/EZaTw2KiNj3r8ldkHgWut/EkSkSd+tyCxEgW04Z
Y/DYIrokUXNruHUiumUiubRgNeQUilicE+59qfeq1CZ5HxeoT8uOevixGiXn
/UJbTR1iYMSTjUeKHDgjUzeblzrpiD5OcbibcpdwJxbAOwLTvviQzAJiXyrO
cnxj3AVd+0BzU+HcTIRBbNuqfn7uxXPmjJ3iR8FiYisbCiOmkinptJPZb6AQ
t1aLwaBWfhwVyfUeywGTmv94VdokqI+3j5vWNzgMJqgq14kOTuzMkQVFBXvW
Eoc+L8FNz69bVnha5nUpiDzV+QMKDBafaBOBRo+8tRFmmW9EF1o3wTIcYvaX
XLRPkKmceZELAflpwq4JsDyem5Z06535sTl51VtL6MJYdKiY4XnvZ48AvDPW
UTlHbh+bdxbbD1cNqTUBzGQitYsoudJ9Aek1SH8GmFLo6q/Q4QnJbXn8moSc
3dbJKLm5cRw+fTxbkWFsQd75FumgCj0CppMHBijkfcXnZ0b1hHFaDdLS7W3K
wSCCrTeDajt4wVNESDX6oUZ2OVeY+mYr7L2WLnK+4kjkoxi9o686J+jYZtIp
+s54ww/5AhrJavek7sfnqe20sxjAcHiVISUTJYO+VFMKLcrJ7AJh3n1/KQnS
jyKV3Ai6umbbT9KTlXLJqYAiRlzf75d9iH7vBvTpixUkQ3n3UwbbjhjbLo2l
vVBVhyvOgYQQaZ3+rhY5J4aBgZRO6x0h1OJnZVbpKXgwZAqW5xgssaLdmIb6
pFyioXyqV8yb2eP/Vj7yfDpKgeBANiEQsqzY5so2k8DvK7JuWGSL6bKQHTWu
Fi5aGUtSgDxxj8KeAkNIXwa4xc4EtvqfumwED76MaP9AWMA+4YuxZx8jfwhW
rUYlvYZy+S10yn1EPnPT1yy9ps2168HWS4ClJK20Xpm/NQPW0Lt5vadvM8zQ
chZnxA7vge9aYR8gsqaCkTiyg5L3Ohrf6Fozamnfbiz1IgVieq7WOOyyodGK
+qZRcap0DmdvSdYjhxSFCwuHVQKRfOQqrr6/FjziOM23U5eOSiyeVXAorAtB
2Rp0bQv9eloPHnyUSZYTfz8LOx3+NF3N0ZgZFfedABJhgQ8NG+irlAsHc3oq
b75I+8MMX5nn8xQvij3XSeX6gFZNYZALvtrm9gHiR1XfPESY4sRNjpymRFgc
0+RkFQpHz5GI7d7u+9F+D7S9qvJdpjuWt6zPJ/yI1WzJ3wAB3a6kQJULOqZX
IN3J3Lh7xZ9dUxI8SeV94C8WyfJfAxixaKNh3KFG271rNbt5aWU7FYtxw7uJ
Vc4s64YZQIsIZNhOLjQjm3sBHFoTfCET1OmtQGqtx/PHerJznmi4Rwb4aTJG
Is6csClUuW2fRGC5zAWMW6gyIT4h7PIyU5QZp9XJTrgDdJRaXwmGh3qQQEbp
zWvakovgtr8lbbx4gc0kYhrQnQpnMX87i+ame4nRLnmWJZyNEMpWL+zErwP+
MC6+TsQXQlxwpS0/RRPkZGUnmSkHenrC1gsAuz8I4ffguztVJ+GP/YC4G+/6
A/Vg5655L4FTtvffYyhbSUI4dVkCj5SW4epKSvgKGp3v1OMSoyps2B2Iimft
txCzt6dxv2OVeg0oJ4FRGAdyCtI/SdHKW/aG+sWKA1SOTCJt1dXpG+ErcagL
60WCDe1+r7XmF2QwzTR/7Q/ASST/YkxhmLHxLQQz2E8hCzvEpiyPaV9+pHdq
6nu6zMi40gvSA7VesZjCuQcbTcVUuslCY+ao1HgTEF0JVoQWpUdDOiYMBeTQ
UV6bkGI4mIl8ZN0F1az2G9qR21wCEt/QlmTBdwHB7ih4yc4+KzBsI6cSMa6w
9C9eAzw/5HS6477tgjSQQhyBdNzQ9Z1zOj6WPXKwrzolqq2iyTI1V6aeQvx2
99qiFC+zC3DRKqUjKgBcUk9U/yUY7XEjs2Eh1Bs5G5vQJx0TyuIeM53BCAqK
KjJYP5ZGy9mL7b/097/fmY/Nk3TLL0k8m5eIge+XqnyOeyevzZgmUi523Y2a
q2DInnIpvxQHN29Pw7weBywDfJUUDdOw6TKpVjAEPTWUbmyj7DZSLq5JUImf
tWsPTDYVB7w4FxQuT8c0M4Kx4OftTos+rC77hTaZEIiuquW/Cd619RwkrudZ
NN+mWSbpfUu85B07X4kQX0VCtHg7yTKoKZ0zDb8U5sGPn9YUpNqkCofX2LFI
7LBQYXWo7mOR+OkgMsmXmBfFgoiq2G1m77EefU9EWuolvRUhsWHa/OZkp43H
lZhfIKMjXf+Y9bIu6K0bBnShhIsiFjG+o9yfOkV8dYL7TDOooilQ+EPYiS/J
HreE3g8X9UreO4G2PoxjO9b/DDhHf7enSOFsi1hDRMW48JKSgxbY3tsn85EN
UdvmS2MigMRkS9YdutBA4W5F8OW37HWwc/3rVI9ISntfvEPPIeqedTrd6XiJ
HERk88rOTpS2YLw8S9BeBc+ZRoPmuYF6R3exHRZMJeRN+wtBitxumP6G8LQH
Z104LvZdDPv5Aa7eVKyeLPbgCtyn0oY5L3ADoVMC0wNFFQ6rIruZ5la375KV
2dH/Js14vkp84ypjmETvXBkvH7aIpqItWpQWNNpFtQQDKPpmMIsw07Rae3ES
wlEbJLQDz9NeZgFDd7MbePc0JCet9fv34T20l1Jp568TQ045nkCcAyQXgsTt
/lyCvreggKAITTHIjknA8QWbynuEt5pdW7Z30B4Unds9doPcKsAqd3JfoWyd
+0VD3XSVQh/dA1BQ3rFa+7nRzjfJdt7fiz0YCdO4xlUGCiU01Wy3erpfTy0n
wuFbcI657+q60t/eMUEqVtpg1Bs3sW00mzh/K/f/O6VXzYV4gaqu3bLxw8xd
gnFxJD9PgeENjwJDR3inMO3/0OgNG2mEKQ4gyxswCbiJiBWsqmats8moW4EU
leYOck6omqaYGPC6dDG95adJ4U2Q/9wCVf+VCSMlWBFQLqA55iPksKJl/kFi
A0XXsUPDpf+7TqvvqQkYRTkAui6CQWhx8lxFo75GY08jhcyP5FVpGMi/DVIo
KeQg9jE1eGPT/qNS97wbZ4obIMQakkZQhLIqayfg59YFsy1ll0t6s+SChvGG
gcZ/jYzk4sNFe2q8zgP7DeAKg5+3a8yAtEdv535KelIxs01UXpxlFFqGkE9+
P74OfoMYmX4slMhs2Mh4te/AImVMCCO+2UE9p8Fn4Wds6KoJx5Vzug78Efoa
UQW4V2thxJifFkOpXJ24wX9NvFm4A8xO5d4pOO+ommLN0MYw2L2AzOX4L4gn
3SWYko63UmlV6+g3Rcsr6waCqZrlnD3DARS+k4lDuWbacMV0fJHqBgjS/gP2
RczHTa16A3f6bVMvPHeN8nY4SoA0I57D2vc/vbEKHQR6fHXnhrKv1TiIPOsy
mBQp8ax8TYaIzuuLns0/yseDrnWJmIAGlhW4jDQ0I2lCmL0k0mEV0qQxuTvB
RCzQHu+4zVjdSXRhwtLXa0LKskReFd6TQgSo7AHY/QD+jUJo9ncz/8uCdAoN
op4Sa0fmkFF9/bCdDRsCQa7Ez9bbHxb6eoXpJNRAAsuEq2+Ybg9fCzWhQOsj
EgDp4BWqCE5/aBwO797VZxLqw1XULF97k7FGvk0PQ74xpZWvO1/QLW+PNFCm
Eg9A4NcsJnNslEH0mEo4beDdQuWB2CSu3b6Ogat3O+r8+OQLZqIOh2sD4z+c
L9smU/S6quH9qyABfRvE0YoqRKdiBs6bZhtA40nWW9VCdRNQQE9aB+Ublj3p
+OA7aHhVKe4Jn3avNl6x9VmNC1N7AN2JliV1vKr0HtAkye9fD8lY/ibt4vKp
E6XP3J/cSc1+Bot9phRSRFmlUq1MT/vTUO1kTTCwLDRhBy2qZHFQIbSBl4l9
FwFC2r47tB6LhGlXULy8LApSpVqT/2WliKNOG8cI/6rFfpWEgQ3MINnUadL8
RoUZk4renh9cSB5/8VVFRBmhNyYnrA6l7hOCBcQB9WROp3o7NrrtvU+M5oN2
6VqQDkDtVwVHXmPmukCt6iWzsBjlfTVA2u8auBlEURZ2PNxkVHbokX0IzLff
AWwZXy/4BDuNeMhxc2b6SFcBPbVRJVph3U9JztG7kq/CrB9lNkk61kWgm4p1
wsY8eAxh9UVUKTXIxC7e78lSTulKaKumXaQlMci2cTWLW2v6Ya5BGZDZxNwz
BCpkDRCUcCBUqurGx48hY7cEaJetDPMmkTjbP+szBseldIpKDdgqS2HMa7fq
0LNTI1cB1wfs3PUak6R/pGjAWWItyo+kIWhOqraqe0oHQ2Vt4oIsIPBlCbf9
8fpEqLf2l1mqb1fmOg2OiauIaEGjHIPAZTl+b8AaxaeokUGpdveayhdn4TqS
A1bSeeTgmI2VO9vpyTQ4+nvCewTfY0fEG/DonXAc2Gzzgvc/9LDKNv8EixvR
Opxx5gIcdBeSRCECXDLBoCYIVh8NpPq3jEv+ZimE3PfjoW8wd8PKm8AgdeuK
i137ySJay9XNB7fcTd1FMmNtIrAbakhWjF2o1svITeZ59w9ZSdqKNPullJ5S
hnsqtmhEJlHv0XKJILbGNtcFbHhUx1VskqQhmYi6r+zO8NnpXXYnuFsmF0DE
uBzroPsh4ou0sekJrlPRaJvLpo1YDf82ck4rHomI5FeSn9AU34aMJKqZXp0H
w6njAwgEGnF+T2vQaPvhIApKRD+6M1JFFDpM4bwY+20YTMHDMj27LmqF1FCj
ImP/rAte4IA7b2w9fzfg0AJR8Dywu8zdkyq64e3eJDUEKNw6/KJfz4jCSwb9
NHVHsVs8R7CseCeAtIeISGCBOQ1gbDEC1QavDl2Mk/wxmqxECpW0a42XyVML
mqNaHD3i7AzEepZacKSoiN33uVo9P3buZR3XAPfFQ0VlmF9CFGPJfLyRSW85
sTpQ/42kxjleXRTAxMgR+xMJXXLQCEbmzh4WmXEDZRqtz0E1jFUKHIPIwjTQ
7+Y8fJaNZKRH7hHO

`pragma protect end_protected
