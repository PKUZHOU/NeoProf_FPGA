// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
oMkCfA1weN8J3q7hzHwgF0CtC5Mj/A4GexWDzKJzcIswrnHPkNT/MafmHe/rKTF0
hCS+0GT04HWsN761IXwPtJKvj5GfkXhhtgMsrsfkZtkMp+jPfxSvNjCsw62pPdV1
/5b3nlKKoTM8O8zZMv3THNoYgX+eYPXNHo1SDrUuqau+JbLIyV83vw==
//pragma protect end_key_block
//pragma protect digest_block
SfRcbTLr/hrYd0QVoAIH7GjrGg0=
//pragma protect end_digest_block
//pragma protect data_block
G7G/74ZVnz8SzrjV/RoDrxu+UWeK5U8+jmezjkgmTwfRd/6HQesXr3f29GhrM/Kg
KoX5/p4LbmJdGYHb+vMSuGNPa8MdwpAwo6wGRnj8DGYHjuh+b/YCjqegHb/JXZh0
qeVDmrZEophQUZTTvp5h8H8aa3m9Uhty5OlFEUXpDsrun62gS1G+1Tk+wX5IHmbv
ue+NqdOct+/UJ5E//+yLt3+uxY7DScA7eg4Aepk1syqaFe9PmWgDq/7fisrWYDwW
j4AsZtrpEhh8s5XF50QeDD5gAFxMBS79sXAGLakifdd0Jhle3LIXTm0aKdqrVLLO
dLLmH6jm/S0nM1ct7DIKRHocMsfDffJ2rmp85p1nym4Csm9IvwJszVET8eYS+3YY
MA11RZybRck6pEIPa6kFReSsuxkH+TDva3EOaA4fpVuDnviRlFlXLqpZ8A3eWkBk
Pz2UPu1/pZYdqM4ABijim3RAJeFT7UHEzT6BUjmL07I2FY/gAD7ybR9uU9xmyBlD
0R5voNDa5AOYtHqpntSyU3gZP2lGEfgm9fUYFETYBCK31OLvnjk9NnhnWqTXbk5l
ELW0aDGpQduMJ3M9EXFdSTcfLWj/cY9Z9tuzVdAxXR8HX4lA4NA2WHEXffG8s1bx
WENj9P0Nx4iawBT+2M1h6Iglg8DjhEvCL1QwgFBxEViY5QfnlzZNhekWXjqUT6lM
tj8fU3fxM0qdCBzzpMYpdWaqgAVhOCv23O+Yv680GS2O0Jt1NsQ00cvTIGaOpHny
Gp7EqvpKJ75/ojSGF5epWbx/RdKUmvxTz1x/HcUJtAhoKGQ05+CXodj//VKTY479
mZ56JYmehjFabS4Y1WvxoNtFmywND3UHs+jLpnzLkTU2PYpoQuTr/iDgXWiCzlfi
vKla2Z+ldPaEGp6Rzf5WvcpjOnMHXwQie4DUTwu1ol72pvEqtaHhb3WoCfYFGBby
amdsRnLpfTRab3TVM4wXP+0Wlpbu6SDoJ0nB/BkBTgmyqLy1XQzeHWzcRvPxPRPR
bwPN4z128c+a4Y6I7dL18voJme51p+P7sO3vqG4CyyViOUJm0lFPu6p8dw1aEqcC
fmJEI+Uehi3Bf4vxW9qp1N7dzgDG+wMY/oYbuhMzv0SaE+CC2aozmVAOUpgevdKE
eFdJ5R6HIhJ6Y5Nt7X0LH2Y0SkQzWRsUIYuo4ifFg1mq2xroCaSbYwfSSYZ9wzn+
duR7JwyYG5dQxtvhno7jMm0gMUI2TmUb6QNWsnbpOXPEsi3q2rwPi69Ic7VWfwny
kyDDZbXnAx/aWxyJhEbVOXCi+NG62qliu29UpiP0fTZL9QmBwmMs41F0SD1Bvd0r
eLgdCBy/Ar00XbfqNWsho+BLx6VO5m0ANejCc0kbS1SmFvAETqcxs7bwf7h9Qfmr
PrhGhD24qkn8D9tblzrhD0/D87nqkau6oXlBVfQ8cY63yrktkIutT/BG7DR6DBaQ
kX/NeuP0HpdtOJA2P2VXMuEexajoDoLgNVaSopbH+NqXmMM3o0FLKWfZ02KnFQ3E
5S/9DmlxTd5BtF0aaITReTD9aweboFhCygCZE2vQUboxFlrijwnBPDho7eAwZ1+T
rJs8jPQ8+/vyfJTlNIh4Z45F60uAvOtfgl0Mt1U9CWTDT4c/Kb7xeGB3JJXUBesg
Kkmk4W7KhEgJGUME46vtTkQrc5uRyYeH2CxgcNlo5/thTw4dxFKx2Vuswq79WLRy
yKti4+veAhiOOBX/crP8/s0srHi27XWIwBQNF+5UZiGoTvXxKvkekDC7qrmYOXqS
e9kuaYz8yWALPPNNlFsDRFT8JPMoOdg60hAigqDUyGFmtp0uUwwM+6vVsKxV8K9l
WQ7IarwnIuEIci2eNNgWA3xdcYEtDRXsZX7mSNx8x5rmRahdKqXK0Om5Gz5R4JbI
sR06kx+mIgqQ9vB5V9g0Ph7zW8jrKpyjqI91K7aGiV5SZh0OeuZcicFuzp9/3aRF
hYHaO4eA4CDXilZGnRQU8zfUjkdWwr39Hfq9D+TMSn0wvYI8kLyC6e2ZYPwjkF7D
nAAALSpRAK6fHOMvobH4erYkY29k/rlEOUPBC4s8c5OcE7jT1rmK5rerLwKGHEe6
MK8GE4H6j+M7SVfg5yWWu0CaIIfuWxtQA9TEBGUmsxdbIpLGE8AnI4m4UCwVz/Sm
nKR5Oqw8LD+h1FFbFVcX3szzWUuMa66r/PUnbh/jyRmE0ZIPxNoYzH/J/rU5gCFg
t/dU6e5zYHwS3MtT2CWPryuwLNzpYQSkJFHLsG6BuZVs79E/dwwK4j0D51YpuYKd
/qiPZVNsxzZ390GSs4TwrbdLnI75N+tjnEkrQIeApoh/XNo0ijGWtUwQUHIct1TB
lLlNroLctf28ld2GLf04FQBy3hWOV2UeQz3cR2cYoI7acOSRZCN0BEvKHlcIS9ke
rZMDrLwKCMS2+myCVZ2pO4hxfGvZ1FjVQqBO3UPRYn/W///zF5yVSIXEB8lYYQDz
3gtHl9oZNS+bcIEpszZ743lwINaRe4p4NYPc1yVA5id4VNtX8wewZzwa11empLj4
EUF1k12rYmlP8fec/oQvW9EZjNuDcEnOYcNy0MZVSV4UsUs6E2+gv40UuKimw1WY
sUzdJyrQO9xus+M2KKuxKJ+H9LyICaQ10dkubYiKWER6oQLsVTb5i9KwxseGZfwn
sVT4iU3a36krO55fMv7iZkJEUiXjcsoeDxC/JwRDS8uEUrnEj0boYgXCi92zogTK
aWRsGWwr2uj+4Br+DT3FXJUoUOzMqqjJJg5AkkyW1PWNg+qVFJYIacdfrIjmupHQ
jfdWyDJsUknRc+EWoFFS+BaRo/QKnFntuXBf8IrF0RxXExTkzmMZpVheO8t6Cwjc
ykggSRfjArQ6xbqYbb2wZNzfE5Y3AGZoDreGV4Y0/IPpxCThVOjaCwTk03C5ce7A
TT8d8WIHuy2PZkC4EP6btbwH3Qxer9BmOZGtxP89YN6DDgqfl9RPqmdGZYwwvs8f
5SvxsspP2jeC+IbvVAsMIvIZpOvenLqsC5oFBLNpvClKLxqBAdRtyZHgUEJar7wX
klfWz72EwatSabb/lV9D2S061RXyVwWJa+LgLJXoXFefIs45mJDfwuVKlmDcKpsj
5DsXDVoOdKd+URKW2rLsyXFL6/79m7wQgJgPuVr/iVeZwQg73yFuWJRM5AR/bTcM
GsONdcCIjN5TsqEUlfMQuUQUm0nIP84En9N4ZtbuJo4JEhKZJ6nDrmlqdvC+yHiL
BdT0qvLmSqDbRa2Zu0EhTSuRJCnk0HcASeVGW/HCavrzggct3GC6JTXi8yN0VsSa
C/bn9ODZPAClCDShEMRVJl764nsHlFkZBwWNUDWPQxh3ak98zCbCCN0WapU2azTp
Pe49849rDlueLF/y930uPpnMUmv99Plm4OS0LlNgRdl3A6vqONX4h1znfmWqZAjX
Nwau80w9pFzOMMOQSyn7K0XGIY2UHFn8Y0xrRXD8zU6OZZmcV5Hyc7GGmzJUMvby
naKsAuwPf1gKhI6SWYF/6RVrib1WPZBWeGOnFT4ebicqRBHY1pSLIR1IOY+y6eik
T1Kwd+yMiZmvx1C5frjdTchIwYAxzy/K9GdHOhnGhViyqv5VY2l/to/lB/88S2LN
5iPUFEcg2Mt2Yd1iA68PDWRurLVd1ka18bf+RuYP7p3U5uyEUsI9ztEL+PVcDYlO
wt9RSmTKlDsJ9y4jIA5FpIW4ASizvWY3KVogC28nNUIthryvbsC5KoKhhdLkecdw
mkr8Q1QuUSc6BC+MtDTgJdQ6J7Px31FYNXo+3EIFOpiJqg7MrF1m09F0kdxTMxcB
BJCyjRnLrJ5ZLAy2uhRIuWwCBwcTJAggBoC8bbEACvMDXlTPTWv2xksOhmNTe46a
SVju5C1CvY8OIMSZoxRITYYZcl2psXn9hxFM0ReZRxKcCDeOV1XIE+wmxTNV8vaz
6YMgObw6N3f2POCvK2eA5epcHEd/UDbipaTN9s+BjZwpKT1UVRh8E+hPtf+zKnKe
8upeW2S9+hJKDwHsCghhQV98hlGkRltZFNKADuF/hIQeU9fI5gra5v1PF3Noul5L
9kXMjnK1zaEFCqDvMMSx9UcTzNSUPvbxx+ghbZU1dafcdryrV8i+nllBV263E2sn
KtCXSMCKnR/JYsZB3GRkYLN80SGm0I71mFDLYnKwCcRDYW/nHEIOYnY3Xs7UD0tw
xo0n+QlhlYp++AICabkAVQIz6LShBvC7vQT3B8m642r4PFhKdqMY0JPGyBkqQUGe
IkmaQ0ZM1QuQGTKcHoyU4E37YlppNzW8jmey3UE/pjQEvk0FsJIBeQ9gB24QMyJg
UNrIircQS75/OKc5wZgTBcKPKJEfkEbEdraeDlKRFq2VFT7H278OtTuWU4O2Zq0r
DqVNF64gzT96YSuhVDX05WTwl2T3d5Etxq9w/F9YqhaH1ZMIRPk+a4yCUkS+CLZM
Mem7R8mVxuVIR+qbk3kD+UCR+kbU/Ipzhph31b6+dAcJ0SKMgzc7QgXkNVgd7Mip
6MRtXxA5YRrqeik8wPjSKm66Myw5gAY2jRJfmhc1B69j+HZZLT4TwJlIArTgpuAE
I6s050gcgEFLG/tYLQ97s8br5Asq2PAkyiDmMLg00O+VOofcgzIJyBILyTTBboK2
Z8b253EhXLj3Ap9LylZP6CouRga8/BnPc2WtbID6/vhiXFQWj+JrNy311w8Rc2jt
9X+bx2rjDKMeLKDiQz/mSrJXb7ms2xr8SAQk5/lHr8D55n2IwnLWyD2b4Hb6/Phb
mftTvhlM7jHs0woopndDJLyF6PbwTiu7zBcUzLsY8yQrbxRF7Gulq2ZF3Koi0rdH
A4xtVqIdgTgYQmX3t97t5HYDMwWRxuMafH3Tdx3uiSui9PwDn8ADXLncIHWu1FMU
J3tBZpTCayG4cS4p/ZAWdCiYQ52tQxyCft/lYqdfcuSB9Enqw0VgtAXoKVExvcA4
yiaCVdQFJRSmpGUhv6/HQbKy+TVi7enjwwxOply6koEyg7YhT9RN1bP6zPTQzPPh
A/T56H1YwsoUpXcDGSYw4PG/OiH/eCin7DzWI1/pWWc2z2ysTa1GU84GY2FwI/9I
BL2rifJwrcZQtF3dVYefwTkW2ENW7oRxBC9sPWFRsmcFOATmCg+4HVARQdJOhGeZ
fNOXTwyizXpetMQQhHmaRTHsVFJ5ac+FWL4pFGmXnKQRYC5x2TCf1Y7gG5bAlv5g
tkQ51qEOotjNfC283UwHhppiOZ08mPjhSpUn0amlCOGLlzMaHn5E25npWrnW00bY
Wa9B1mExiCnF1zowALnH7T/iGsMuB/Yg7mYWv1icpsvyYLUJ6JMHtYXFxv6hEqvc
mGin03cqyBbTjSzSTg0YRlkusUKgpoo1WCYHqsGLrA3JOyrhFmZpzFuKTRe8pc6o
sYvhfY7tjrmIK7nnwvP7V585ItD7GkZ2iuvFGl64FWYCTqp6R35jUSdILb3b+G7S
fPyeTkUsZ5v8gtfpbV4ylsOztwJD+XWJ1v1eAM/O721+avXhPIBNdiqxwLCcOxJf
lrawxYXKsPNylCpCU7r/o5dOhh+nYfPQE4OX+3gPpjwNSHufp07d6tkSWtPYrYrZ
DO85eiVcjFvkVao4bYFPB4Jh0/lrRg3Iimzm8Mg7d6mfZTQSKNpm/akofmHmP5yO
88IMaOfDkm1kuroIKVT14M72QigkfVGXgpm0k1heQMOtUVnOnyM6UsLCpxwU/BmD
g4FY31rUoatsnpc488bPmkbz4rCZA0Q3hnQIUQBN51pRayAhECloHjb+MIhautQN
xYbJRdCc+1wdzv7Zws4stgxHF60t36YRmLBsDyzVou/hMDayFGCFbk+S1nXgdj5j
NZXRFGHlg65pmzmTFYXBJuNAyVhgFtJDvW9MulbwlnLHpwCzHFZpK3W+b2psIcg3
hdRko9tUBG8B1PT2gGQ2z/HwJHLXOcOtnmMvzvRWpZNBHmiDphEefFypAS8L9mmD
Spt3PhmmaI5t46G+VyMZo9cAeSzxKfekqhza6k96mGULpWQVj83Ug5MJqnCuBwsq
e5Wdl7Ky8dAP+UD/cIEkY6bT024daccKFjVxAHjZLeBDo+LzTepghbKfGPBJp3jw
6qPf/KUnVVPSqONup+JFZnrPeVJLjLvo6y0hllmEr4OYKvlIZ2Rd4AVBkVlCKt0b
H9HUATdQ+HHlzqoNjjaJ8JJ95LWzsjnvkud5PIc+HnSaf7z178fqWadnfGeSaT1R
6LYyXPoEAASiPfENd1MHrz7J4QK0gTV+aPKCa4vn9IBKnPZ+a1TwAyFf/BaJZ816
/vNlHT3C8oM9bgpunQbnCp8tZUsj/m7pXmQF78lhfpr0u1qYcXmxsjRsww+1rfyP
0Po7CESJsiYVeG9JTzixo1rcUmJvfDHgQHVYdMFoaXgzE7YNL8g3sJLbw8RWt0QM
1ZVGQmUDGtRNJLOCeJQ0GJY+VmC0TeEJxZ7bHN9APVGPcdL7Bvy6ip3MN+K+1l3c
QFc830/L96Gf1AGNc+li5Aizg5duu+bllRgigHOX+Kvsd4FfsUw+fvffNjrFREVm
0x9uKBlHOJRKTi8Tb10wzA==
//pragma protect end_data_block
//pragma protect digest_block
hzSnoUeiarmXPIWDYCo8x1knGG4=
//pragma protect end_digest_block
//pragma protect end_protected
