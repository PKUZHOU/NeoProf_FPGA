// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qV4+/SNEDvgU4cHDJ2g63dLjSMMxaG9QEjr7pdgaB+26SVJeQfjIp1uhgdJ/xX/S1+y+OkRZYZQn
XAfMAZ+YTM8GBOuTxoDVXSBfMqOA4sxd+3/q0/IFd+chGVeE/SvlyUsVoMHyHQXmaBsowGfJdmXA
IdX7rDyRUn1F/+IvYYjqJEQe9ObxbkWMzr86eT0FdBSzAwyLBUKSNJHkYTBUck3y2t1Twr0KfWwh
hl/PG1rpM1qVfygXFX8Nwyj2itpqy3Id89F5/Mr0l1XJAoqGTJcNjyCkgSzIMK8xsZ23dnjA0+yA
ZrIjTj9HoV3/qL9nj7B3BV5GXrvJ8641GJYlGQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10848)
amPNV08n5rK0oFVLdcVDkVOpQ4JiG2WKEiK5eMfeEBZJhBHX0vuNfQnRuKc2JQTtzkxbKdNcVObE
xpzTwxmz4YToi2cjd9/nWVEDfSQQSGS07TV0GqFllIwGTHAB2JuCjdex4lttQ88QKpyhjzrcgNis
FP1WK5eKg4xyhIUXZFShIv3+wfDJlBkRyW+DwmH+PB2wIftaD7/3vmR1RJMGDVwpewTHrcuYqf6l
G6zSx769K4l6bwZvek2/XmwAOCj6Mkq7iCbmQvt/0xnFS2k0qbbzZk/tkFtMp6cGqS0UFyWQnwgM
7W1w0D7Z/jqnkqaqLtQ4wKa/32AouAyVlwPBuU3n3NEkgIE3UVO9u4C/feXjICBAmE6ajDyaxVVn
PxiYUyVrza8zZHvHAOqCxLemltgJS28UysdoPNc32Jn89wQymlOK9gc3EIyN32oOz2G71a51csQh
PcB848YvuFkCP+MbjQoe16kEJs24iVCTt2rod2I5YoolINmVFCjVlN5fgpgIkAe/NwDH/Vg0nVGh
euouU44qJzvng6DT17+cR7vbGfWr7jSp2+eLMG8kbqjJWR/X91J4qsaaDj8y2s0rSPpfV7XDGbfY
wlb2CiM4mLWi7hJdNdNzMoNTao7iQ/P9G0/YjzoS04pHmgyYpQ/V6kbZFxCrvrkvfTEkXEHXvi65
z5gID+Dr+LTJ6ZWN4wBSnIVLeFSuD9F2kZdvwY61MENbW3lhh1rmt0jmO1gW2ENUnrrZ9neScHSy
CBIJIjIwL1UPYemvKJT/kkONAU6h7rPMOhQc0fs+qUMibPTWaeqygBO+I/YQsXHkGZFWLMPGN84g
IzQqb+3PSdwYwCXJSebVoIimKVuUWA50CyT+2fIozUiSx4mDs7goaD1eJay7/LzDW/HHJ1g94W35
t5dR94aFETm5VZxspBocdMh6Bn17byuBwZO/hcpz05T+gjnt1OZH1qXaYRHHqwq+9c1MYRRQRwXj
8F2arpZUvmMFA0WsmuKifvBxXMae3lrN8YDmD8DqkVEVwalpV86ZpaqbnIYixKRaU9D3SAa8ubmu
OMDPAyPxAo8Zkw/vqE+YQbBDdgQu3OP3YqUYkO2XdhO8u37qZYvQmNUocTaR9d9AtC/3YzgbHrFd
kZZ9H3Gy8iLDuGFXKBPBgCiDKAjjd5EOAlLhtm3VfUV8amwpgvI8SK+kmBPYw4nzkE35yKichGEP
dKZ5h/GJpx6tBBszOY989+i94JLxs1adRV+rTHuYFjsseUwzgp6k9uB3AbSQiAEl+xYPk3N5o+9T
ALcbJR9/ZSm8eoys76XVWulEFaiCajd/6TzKoAKWLfs1pd8WekAiOnhcgpZuQcVZ35F4s8FZ8Rw8
bgYQKH4/MTgXvazVnMuImRKNavcapiZtgjC6ood4XlLFnAIh5ClTRho/ed5UdbeDsP5RKQ0niLle
PihPwuZSnOCPBhEYz2DtSEbDd/N4PCHfi8VDeWpOfagOUC+pmL3Z40sZlUkj/zKJnbTER6qJ/gKN
/aCLAu3anSpUKn3cN2Pg4ZrVAH/whxKGAhLo6owb3spz6StyHIxZrwmZ6tVtQzoo+X3Jh1ZJ02gT
Ygm7+NNmkq8U7e6MmQY/kN8OZ1u/x16FL4t1UkFq7zyuM6HGUFJhPHPrm0jF0tTF1ZXyY7CoqthT
3x2+8iigsIGlqydH1pFwdwaSvf35MBowx6k4QdNHSTXUywa4yb1kfPWUyOXrydA0By/TGezMNhKl
8LlNZKGwQvJPqpaz4LWF5Q9/8QUEZVasITQ5JxC5YWTjn9cS0E/5/PLtmsBZp33NgDFEc4A7LeIh
4o144Bj3smfINAw2JlJLz93ScuUOufeto6IPWChpD405IFP4glpKTFjoB5e5DO2xmYRlz200FANs
Z/jwAP/Lm7CHxC2N/DjeVoI33c3tu4kOLv+y4m2LU2zMnFcoypxR7craUfhH7ey7EliNz8lYgq3k
IQD1zcAzYu9QvkcpzOz3st41g+s4lCQ7xmZcZnlxh3yKsyMUhF/VZu+6X5chi+9sjEXQYXhcDU/2
MS3Z8oAA5uo8YypSFRsCE0M+mBPztVzuQUALsOIzzwgX6wMQBkxPTHY/mGTPlAlXQWYHFfwD1Fjh
Vl3qo8kcuufZwIlu0OQ+tymf17/xIdYWul1iR0PKGz/RHbmuOgbAhCNqvyqyhruQ3ZFd6+DppgF8
VQhzLQkoyUO0bdt8s2WZJ2iVh7+4QpEshcZJcUMf3zY3EHZ1nVvrJVYH9TLdtGomhStwDNGqIAM9
KWun0d/WpwWfB4ya2gInxiHE/ZVTt9cflKxLaaCe23U7Uj0soM+EJswIGUX8G9IdRrTw7IphX8qV
CXl0Lk0Vou7P+J0vRkw3t+V5XeZxOCeDhLy4UTQFcxTa/sXjZK6wXGj32gtKEhbIKaL/FP77ojlB
kVntHjsG2SgrZIR6QH7/2kVEB8d5M4hJXLIfb2K3SnCvw/3GFAsnkn2QkpJMyNPviAccF2JBW6B2
z0dsC4LXHEHTjOXYw9G0xuczqoNPGmN/uebCfW+iYH0WLq8GbgMTe6frsvRtPTpcbsyPJzYQ6hud
ZWimusSRSjibUdtjDL+o2e84eii5aIXm1nPwaaqCvaOzA3epfbK4YxJE5bkKMU7KInsLItLfbb7R
qr1L5OM1HFkr8YtGiBg3FOUD7hE8/3Qegw4vjlbqJ5BD4vHX1F6YNZ4Lwkck3BZs96W0GDV/g0wy
LZn145fz0Nl+ea3zHuaD5lEsxVWx0asJuC7I1/KteHiWtArwxHVNH+mOXTKeH7kN3nnU5aVAVK0p
ulEg5blvGY8vJXqnoZR4U8gOldVfSRPRga1bwvaUFXzJwFSV6zdUjOFMiqRtHmBSBFlbFp6spLzU
g/iWk82Zlh7irUIvxw/eYHjQUcXyJTEcEheR3kam279BxDSQaj4dKzGpVfi91jRPa07MdtlpQJhB
BC6ZSIBcJSMcHOpG6AmBTapT2PxJTG4pjIIZTN0Y8P/+x+bFE/x11RHItq0/D7jkQzHRVOouBr3u
WA1QXk2Hpgk9A4rFcBQT7P1outW7mtsYqnRumHrhn5Xt+1ZCmLGX/bSQZhoLEngLcEeY/gmjSubD
8/8vMUGvScqpzHh0oahPbCwtExGNCbR9FjIf3+oK00SgW6kPsKm+Ai75awuK4NFyGOOA6OJPaIft
AoKxoReLfvzRADhPgj4jpJdqlch28val5AbhTHvACCfeRrBvEoWbDsgahgPKtQZddua5h3vrOb3u
QxzeOzZ65QcHmP6wJEWTdJJGs5DaIQwsAF/PIc9IknkgEYljjvzsYI3W0OevE4HJLtNMsqdjE3Yv
ry9lF5XaQqYzB1qZ9vqK7R+6NFDrS5bR7iziPkuGPo/D0WFgTLe1QYHcL/nv5RNBHJiDO8oeI0PZ
rmK1OQu96xJU1KM7vj/y3EkW9YF7KzfR0vcc3uGeZJ29h5z7JW/Gi4X16wAffMQewvvxwgjBcuNQ
NcAomWXCfOjoXtIcI36UyXUKq41xsRrmq0ByQ+K4xfZRansTxtsFntXw6Xti0rq1EvjxCLt2ppgl
mI11fMBIVFwAZ6ZZ10OluOhav/GK5tSVNxEiS8e6rSG1bC2nCPHBtChhqtFZB8l9o6skGUKzXcZh
OiUe31iClKk/TzjMigu8pmsNqXW1MWiDNfyYnYYD50Z0F3gLwu8BeHn3rFXM8kXX1JStHhy+835z
zQkrRdD8ZNQctbOHsbpPOjHf8l2bvsFNRZUvQ7gr4U4Uaw+tX9WX8DoJU+dlWha68RS6kR37Pmqj
HBQOKsuTDHXM2px1UsnfaKL0Ptr/yrbMpszlisMObxYF/HbPUrSugLpXgjQ/lsa6P8AeX3DY3XQA
VIOKoG2WFM1TxEpUCkvUBWQ5qbRGW7EOZ1zaN8KIxtwckMfh7c02iBB/yVb3ko42NMpv0Tcsyc6a
3TuDUyib6+u/AFJpY+CbxagKEM9IbmtKHUyDnNXhaihJNYOpAvnUgmDMbzhfel8k2yA8vRX1AJrH
tIW31YvITDyyrfAJHIAhUyg62AEwpSo1U83U8uqdh/MnoYNOBveStvIhDg8Ai+Wk4oK2VJlfJx9n
ljjTg8RHvferyCqU/tZEq/m8SrkUfgQAQSaAH6CEWZLtn5seJHjQtkVERcD++SIp7OaodpQsMKFT
Q7eFcpBNMFxfq/8loGWkFUYNg0Cospy21UiDxgJSdFi7Ni+QRVcqeD8yE9X1yyJj2RnlNsxABycc
6ffm/x1y5jZd9pM3ALr0aUA1690/ZjE1nOFDyKxBKChgi1uSCaDqPu5tsz1GUxkbkq0T8sflgNUe
MMQ7Y1O2S3Clv1lz5FCpPEPJmP8J11dBrcspj1oJ6u2jFVIZEs/jXY5fnHY5o4z2r0Rym6v5rpnl
Ljm75qa+VVb+0dAj0956BYVdflJa7iTANlF1DwoTLJsxQ30g2a/6tvEHvVt23ifZa27J4KxD2hmQ
lraXR3Pu86P9UH0YuYZkHMqBJAGN8M+zMllT4AoxE+N7Whx59qpvP0blhqUMFYr9ThQmPj3DLXVR
PPBjFgxdTXrVaMjglZDJP5UTklIRefPUkuhg+Ot/I7a93BimiscFoWvM3/sqy0Ogk3KhJkBuKmW6
znJVqj7qPx+1hu4fngQll7DZzz9qGzWwvcqb11uzT24CNMAx5O1ohbwCRV65WBbxZRAkKxhiFPxb
1hxyzUm4z+c+gi0MgU4gjroP+HJFKRuNmYG08lbPbNobSC/OY57X5QRlBs/wp7rPmUSC/LsnWzJz
1tE4A6IVItnhkBHzvR7Hf5IWBFRTRYl6Srup7/T0LzzMsKNFU/9u+UD3vftNL6zfv02r/nrHEhWp
Gl5kJmCF6jwihVn44Km9ToXp3eR0Iqi+yciH/RvUY7voz6RVy3WWAvn6IV6WESoOZ6hVmTDOU72l
UTZw5d60x5PtUMgPR6PIQRwbWY9nq1If7cB1XZ70l2V9Lry22XgoZvIp4zUYLXXvu4RoT0jEQldZ
2fJGuO8h3xG5UKHXVZtevNRDL2u+N2XEybOVPJ9dYZcL34DzW9Ecz8UEt/vZ+5/D8qpr03XYpsA/
x+uy9GvJh3cg9PlV8SMfYOf3XK4r366tNlc3qVAWPmqAFHLdFdP/6bpKISAEybgcrNxGhzYA0BTP
Lj8oAgAyvT3g8VGjkxAfxl+PaBEnDiCXLRvU2vYGO4uQK0SYKOuu7Qreni3FpZrgATDfVrtZFJ9U
NRcNZSHl1Gy1m4d1HXz1xJ32LPhT+Kk9cIM1uFGjExLFsFQYCKnHHcXCU19aMtG6VMCDlVIv4h9r
T2n45L9T84Iji3e26xV/E8mFaUd2dAlur9FQLsCsc0Edc3xkL0LSsJ2lpR+BqmMFVECh8SCB1Tt2
zvUgsvHygs/XjpszOnwXFIFZbAManAz0lOAee0ThdIm8QcIDsp4VwLccMpvQqEiwKLiT2AVYykiK
3mu4AHZqcM3ZHldkzJxw9PbzdbVnIiTdrq+IkEr/le/0SI6eys77KmPUhqYWN7ArAqpsgsH0gTeR
Dkp+mWF2DV/oaDmmwKHHw9g7HrExE6vFRIweVm4m6kxT5AsZT2X2cAJd2L/7sMw2GvF/f+ZxWyVe
8dc+Qyd0XSrg1A12rFMU09xveMYD1ymDxBy5Jdv9BVtBdMGP0hMv4L2Rm9Ry9z1FhG5SENsbhUyk
9M//pjekwkm2QYDSFokKdqIeKs+lR2pTnR0Qd6T+p8zALttPqTmjsXYSBrV2klOdPI6c/+vyYCkf
ghyERvQgRHo3hi35DEVhgYImK/5OLoj72BNe56IDJ9LQJUHKfF34AvoTaY3heOs41O606w7X/Hv9
rldWdeDxpCWpid80gjzC1r7GMp6kOIAUZhkcsrQs50L5zWTNR0bD7YnwO/GVrcX+V61wYWjTYxtp
JxNSVKDy5eiZLaUtyYfxXInhJqd5S990YMG45iK4Jd+c1fjATD/HHlonwTqb2GBRF8saGp0GI1Ri
KF5vFG98E+mS/FFve1fGZNnH8pXPAPJkLER3a0zpraa8rgLvQhzhvUokk+TSfSjGrCWgek3xQGxL
dUn4LiuwJBOb3g40EdFnrCWtnpZHUhsy+H2IaWpATGLdkASxiuU5TE/6PSpPTmAubXRmWDYd6Ten
0AuxJ2+cftY1Udl62HIkiRUegOln3c6Q7K0Yeczd+5BQwiG/EwpMG/rGba7UjP+zxsdGjee6LG1M
/h8bwlxgxdk4WOUwmm1o7yJ9idbCPhUb5q7BJUpKeTjE8lEdGjDD/aIsZsrTldzuwfQqxHyKosb/
mTqcOO6Yg4l4ammeRpKT+hsIe0WaikrCwlU4Mqh5hGyvoAVpgpjpYNgfUMAkBq0/ekBLfccxoEBR
4vHqFd59oAaT4jrTzufGfYULWBuIYrX50Mf/p+0GZnlfuQcA3AXepRl/qFKWtf5yxxBEro2LPZMx
9kk4btjVTobVyl0x6s18xcDPIUQ7u+pvz6KfHhpomqrB4H/UqImx1tEm1bjJURjN9DGMRAz1ALOp
nWDIbwtvuKE0SMqhWmPj0q2zpoL/J/X1I9QiRbKwy3zTJCzusdx1IuBicRKbGVZZFULo386lhw9r
/k7QwQ8DMj5M1GXbHTvy0RRtUa4QhNhtXHxps6uEoSSOZdqHXIrakRHrrQVkhBeOYRLe9Got/VFn
vWJ85GTGkShVh0fosZYdLfA712gjtsTKeyx8QubPNrCOOlfB0SM12AWva550YHKcMK0vUR0vjVUk
NFT71YZTCiiQkOWK+mPp18Gso5B2Nc5B+ZeUhq2+ZY2wP3MjWOmRdyWqFO5rMN3fQLbmgk8dZRJH
Z5R5sV5dvqfNiC8sYRAvmW5Xhh7FHXzCWjtS8BmIrVdxINpUNRiyjz3EsPrnvYaIC4jyA7m+JQ9n
k4ZWsX5PsiNT08QovHzhRXtF/msLD/md7g6N2NHqY1K1NCoVaTslcIvA5tKSGOQ17afishmzA2WZ
ob0ei/EIYRPEuZd0n0DUP5pMnz6dX+aow/536XVIX2un7s9mG3+HcA9LOcIH0Uyzs5vm1naEv7A1
Gxkux55SPw7KXb2GIkaEIgvuUvzpKDVNz3on9X6qJjrXootfykehMX8bKAFN4BrhZjlblMJZtGr8
SxoI62YzQIMvbt4X2Y0BdV9khGFl3M9qe4g1zKW6APxVry7bzfd/p+FhSVEZmT+k5f2lVBiVTwLR
fJVUx05Yy0qvS1Cpv6Ckf9e1Nwe1VX3sLGnLE3AH6NPsRd7TTFX9ii0gRTCeGaPyyeQvMfHltAYR
KSidjP7z3k+1dISpE3Lml6b6HPZs33bYTfLsDw8OIUvp5DeHXijfpCOJCP2p3NvUB0yLiVbx0YTw
4pIrep5Ivt+FaND6amDTZDxA+rHipdHhFXj8iaGqV+0c60QgQu214njuzt3JHaGNRomz4TLfWj3s
oMfTD2mpWVeSznvAu8D16WYxNX/byh7BDbl6kCh4fH/2wnEqGdhBx0EajN2ulYb2IrCd49fPyMl+
ILno3FdSPiI9ln3aszDa4zTpH7Z0u+s7ic4EWzgM5Z93yBQPqSi2gmsI7EukcLU/vDCJVkf0d7PF
uYPnv/tuO3gaNiHYPUrotJ5mhncm/+YddQP8KJ3dYUrnh9YMfJeWKgBybOvSAS8vXaR7KvfcaTpS
6kKc4DzwGKGTGI4+1FqoQF1O53+/cFuOuox06ndYWJWlKDLvhYpOGn4KgzAwFinr/VdlGjnLbjqb
ir57+dG4Q25ZshbXvXq98lYX4/O+dvUqSuqZuLJ9ZUHWf6/HO12CXdHsCmnzyf3g4pni4uo/Oix/
S2PToMjx9W5vpRxQgy9i+j97mhB8tgJ5+prj7mc9gjV/KqENtbnubFOPLgI1uf/Zutkmw8Ufn/1x
pGiLUiLewb6kajpRZvQ6uupc33mJs9haOgqbrPmzbv3fxrAz+yVwxglM+oTm47SuKvl6htBq2UqR
tU31nU4MnwR1Ne2AW7fIuHxa4Nqn7eq9gHaM2LdOJLNzvl53IURBmzZ9h4QwK918DEuI5694WQGJ
kWTq1aKKBSIuCFsDZIfb9iDjXKLlwxhzwkcGgPMVVuopIZwMd2tapWufxzpFPzq+h50kU0RJAL4O
XT5lVLqgXRho22MQjzo9FyV1XargTVrsx1ljLpt5JQt3t8Qege/hatm9z3nwJZQX8rCO8uP3bUlM
8T/NvKQ5AgpLEpWYvTWExGWlkSLOJYbeAz91T+YSkbroZSWR4T3rS/nzTRlTJ6YrUclgz7kStijF
sWtZPGQmMBbPOsBaH+9ed/+PhorWLxdwk06hSdPvESXmx/MVhkmmYEZhHJYv26p8q5z54qrSV5Gs
4lp74uEe28RXemh9Q4Gw0EiWYV6uwp8Yhb3lpV99AQ09xQZdQO5YJBQ0XoUPRRHl4GhclGfuQVCE
cDbgQUYzZJTBYKgSFu7KMPID7fHMa8fPVf87VaicAlusOBSWC8L6Nyu6jkNFJ07UJF4ab4Zeo+Nu
qUbYSCuSbZUZDjrz3nvPzE8/WHJunKPAbjuOC6HptGjhulOVhLD+NM2la8CvrfpdbyV67sDzu81r
ySm0HJUOyfBzYIYINM7Ykj6HfI9B3VhWzjYguBnvxGCvr+sQhAXer+yIUrYhfE/7X6tER5kn4o+z
n7j3wiA+ATLGwYFuJ2k1FdcGwlZNUWuK3VQ0Ft3tF8ztOiwrHJqBMgcjJP3+TDmGthGtfUtJ76FY
NqS8hxXV8ImZsvlH+ds/G1XmuswyqWhXG4f15PFQVMGc2MmjNQhiKtCKac9eOXjDMAFRItdlJVQd
M7SrSWdLdjJYaLVCRUQtV61kihRjgMVVNRCmgdF2S/HE3DRd1fG/4s0qFxXLHi5zgyo1rzyTLcj7
+ushUmoHUqafn0eq5fJQ3cSc9leV9mdbv8zZXUToOdjDYnIz39aq3fLxqIESKcFcSG2tjb3LZ5ZJ
fyx/uI97J+hlzrHaGJghSqavGkGHOpDFzsjOemvp2Nf4JrWj7i7V44dDYtjz9vVpL9y++7fd3nJa
7IZKu4/Cmp+JLyrf6X0NDYy2nX/ZTWTyHQikAY7IYEuj612EnrxK63TmdADIyppndiZhXOeejULX
4dal8hZePQBikZvrV31q+7hzgYdgAsVLsWn/Ih3updgaKtHT3yQGZrNH1WUyfe1ecHVg2twrMJkC
TAaep6Fc/clssjENbanqGoOghFCu+Tj2qVJGGyzzD4ZG3jznen28Ug7ezseShfmXKbT+T2dwUDB4
mgUG9wilPjeQgu330Mtp/uO5PCERCYDRk+yoOk/rvehRjUifE/t3L/UPw0xHGHMCImuWk4uacSFs
ZIGML+zAzH7xQHo0hQuVag5qBX+vIN9zSEA9QqDk7fuyVtvfninyLEZYV2846APA1wq30UM65XUQ
3YgeiDk3KZYhGPmX7ZTWdiovaMh8Z8+cWtBdvvsVNwInQvIvucMfKP7qwTHBnz+7PQS0tzzip0Ft
PHzGm/lGN+CkKWbEpE2NYCjN4oEvhfH7CsZR6aXBltEFrvrUfiqxYE+JiCZRsOE7wU1Klx7wad9q
bzUCs8vdDrciN8Zb2WWfjfbesZyaJBLXv4w8D+OhYQvQsKu6cahlWpezh/uxhhVG7dzLgKNSU811
H6wMVqHxlNAZOPx2oel3+LuzI9q6ZryoMfKdBOwdEuQq3uDgvkkunwvGGumt6QkfiBq71FJ84VGN
gdDRcVQ+1GZxmeGGowuzqanrzyQZBd03gJMIcl0ge3bPNvwR4v1NTtJ731EQCdCDH2BADFvt6xvO
xFiwkEvQ3PAOzPtJBP2kdTn91+oV3j6bOAn5xL934drqUQeHkbJu/UCfJwu6Gm9PA6ekK9epX3KY
34Fmixwv+kv/Fwq87qMQ5qDN9p/tojkyMioRbbUPgjdfwSG4U1Mjj+sE3lKXLaI8CGipliWDdu5F
TcVl77wWVOffUcS5t9PQQK9sAvbF4UPTJYE1gfTnZAnCE94S30gZAkamaRdvrfQZc0f94F+ItA5l
TdQTpNeGZW+yNnAssCVE/hXWgBIkoKL2MSPUCYBdt+N/T/CKmOiVF6+ayYcYxuSbPXnyxOLzkW8n
eW/LE0tN9VmevU4dSDz2mSYzBEMUb8zL+90x4NWoupXr13RloveNJkPq+m3AZxSd/GzagE/fIIkm
f9cy+PYhEZTK7KZI00enFFCgWw1xMopmxtuvzUJ5z+OnzEGWXkfHTdfJ/iU7dVpzBItarZMttn/R
Fx8fccL5A0p4t2WQmR2kttm9uC/qHKqsOWmNsBSEaJBqhjcOAcVLmopYWWDnRQUJu72Pqgh5W7CY
DVZjJpt9ZTfYSfzt+mRBFT2K0WFA8yKu4uKV61l6k5DEKkghGchfGqnYChb9blXQE910rW6ExnxV
osCImQXT5StSwQjecWjSF14XUFzPrQGYlcGmm21F8JLMNepmBgRBxmhUfwb3HmjyIK9btrX3mvb4
PjH0HVzO0uCbf6gvaixxBq2yMM0V+h1P9b8BGrYdMGAGSZfVIiW0/oImX6SMVrm/iGnSodksYqM3
btMs7ylEsDPSydqPPMBmOlBBAI/zWRudcdJiwYhuIml5OMP9Pg6dLqERYu842N0OBxExaKsguIQW
nlFjOi3eQ/NYPYdpRvNQT5goakcg5CCrDBbrS3Tia8xcQAovOuHMvE7mRa5TsqmNFCPSjTi2cuz1
8x7RVB8XwDtcxdmxFjLc5Jyelv7lK5REZe3nkfihseFfL9JTzwTAdI1C+0oEKkL1787GGwLyQJgw
TfxFmO2ZhMeAyqzBj+c0Uh0Wyhc/nPGyMuCCVUWayulDUKgzJu2UqruZKSCePThAXvaiUP3e2gcQ
Pw3bZg22b+Er2ahaPs1H3dv5foUQQ1OMXcswqkQ4CcEf9aBwSU2pyY9V5RpDm0MlRA3CTc8SyGGL
ssybykGF/heOlmTRUm9M0gGazgVENcy4+9mRluDWI4zcmI56DZcyTJR0aAogp35J8b/OrnxlysN8
gUUrinWAE7k7oEHPbvtNDNGcSFAmzZYDoyX4zC/0b8EaRPdvmqQQnRhmrHym1d/jogTY4RH5SzX8
ll57awnIGC+WtMxqf5IkBowhVwndP9/IgxghF8a+UPumi4H94nkQVxXFMIOBm2ab+MVatA5fQXSq
PqjU6f1Bu4LU+L/WuWIu9wiTmqfwrRfJaLdlP4PkjkEIawh0R/iDMHsmA7KAD9vmDIVgN54Dkmht
I2wai6cARmeNCCBMiwc0qvqe1K2chP9a5lrUiQ93JLb7heVv8Uw2tgkGI+Z0JNPMqvXES1772WUh
taucGVPXCO2fOucg2I5hZyJ4TlENWqf3YQoXssbuwvj1tVMaYeGBwiOajoqYwjK+LAzlaEZMj9Zi
O/syjBi3bT4XWeaB5eeLGUJ1/KnE9N+znRNjwrgf8Ogk3RzQwu7VIaSa8KZyTGUeCj/mL6wgxvk+
1zvujh27woeOxr3kczt8+83Dp+TdTP0B9xMvrMChMppj8Fd3Y2ak6XUfDxpCQGZeEWeE6LTBABvk
hQdoA3KvjYY781K1UuQSPMaHgkfbJ84tr+iiL/p0jyRiiXals/kOYSJ9d7ShaZ3iuH0h/qvKfole
LWZQ/ayJZOYVuPjO1tlnlvvWz9x+rSHy61WAdPXUMEUAn5OrljdPjeHY3UuS1kf9PTwH/Gu6ZgaA
KeVcXGDhi27lcl752Lg/1oBENzydV8s41jqOC+OAfuDwcvPcG65TisuaFlL1hq3m5//phTi8T6OB
3yqFB2SECuoohvVI55VCB0zYXf0H11fpOFAvdvXe0poGnSadsQjf1uXHwdD7QCw2fbp/oGHWTPvt
FNjCFj3GcFOJ1N6lZcyKf9wOVcUNAoMb167s5MNG0nmkP03V+xoLl/eShFiAIJBFi5hpGIsHQ5S0
GKTtT2BNPWPhwHM8PF+bpFcaFYAZWW3uH5dbirsBF1dpnOYXHrtJgPSHM3achxhBKr5vh31iN5hU
Zlf6HDNiaRWwoZf1niO1X3mzPdwHkqOJlh/v2XEvyV2gZ4dXR+tRtFWEZS8nRVktT32pOFgAM9ju
OKtOeHUiJFZM+l8Zy34uYYrXNABtdhtoCvzeN7w1Pt3vHasEaX7WS4fOlzVtAwB1X1CykNl+RJPL
bIF78fST3/wWpSPFtNV04gZEjaesJKZq0RiOzV5/i9canHzBBfYd8fxoRzD3pZJhn0nPwllcNTj5
445QJM4squgf7RXvem9qNbNzLVxm/WaIfHymuQe4GVRm3U7+qeoACf/MQr9KaqPaw8SdHEdmyQwK
oaZse1P/I+sItf9OOIYHC5/UL7w6Yv7p95He/E0Ccpo7N+c5RDoA4gGXvbqecIxvXgAxZ5FM3FrZ
9DSQLsuXk8yISmifgIigM/Ce/7encMh36ifcS49mdzNk9vZFWcY5mssawSoQ6Ok/qCmgZL+iLi3L
o5oJYFuduhNfUx9v8ZNQIwJQ3lwHl8y08mq6Pnud3mXPzwgUgEW2r320h1dpQ8zWPokUt54iambN
8dmgfpmh6KW9kLmxmZrj/DiW8Y6EUntm9zJBfKm9iQAKJrl7hPdQSBkbVnFvOP/t+JVGOCY9onsA
ItgzZjGnHat1KSwD59ZwGYlOcQnYm0jtos2H3KOGG0QOBxC+1DLff8H7e1fFdk0h8qEr3bK6y1Tl
VZ2CseQAKozM7E+YzELqf6irwAJVOglJxVhTVPN3BHJWIYOrPk13mhHFjEZOnAq24wYIjTqlQhQU
rGOGztHde9ngbUyteUww/91Hia73L2FjvzFBmnGaeunXrBc7uw3SqMLGjA44N7aKjdWdEI9Yf8Iz
u71KK0SYNELfuT7NF4MBku9IfIpX+avgkmfbosOyFDlyP/pi/3oSz00dRv6Y+ct22u7LDmJriwKB
NFeB7ejY4KfMjxJfSjaFT5za4oAeUilsHGXeSUJTAm+ET04sPTQ3qFxX6HlalE9hLnSSoJ9s9N+G
TFRdG5wj4VDI36eIK0efW6TP7GSTVXx+ufwWJG5g1CvxockHgdBmWzJtDzPlJ9HIUmHf3KUie4HB
V23SblodzokUnzONDCP1YfPrCvNKgvzd1+czY6eEwZpjfgmNL6ghyLiSzMbXxL8xhUwyEjZM1Cmi
cpjTXbntkfAeqfR3jPR3/NOiEf9sjyaowHilm1m4jbjQEfIAZMAtL5Fn2G3O1fNLfxh/ZPnEp3Qo
fsXrSk0aOcSYawojw597AoYQgklNQDrqdGoGyQaeHMnktT+sEVfsrs/NkqXnAeAWLOWQs6uV/Kj6
jNuvZszNcHZqS7R/rEjp52MrxpkcT+NM7Dc2Fy6kw5wi45rhuJnKOSh/e+SnyZLR6Wze9qDnq/It
uVNYM2MQucD1D/HcCchz+4HqCkBky9hzrWmunjpl0KcvY7tKhxw/hVvWS8BvETfCFJqGxxZ01xw5
4Gk6uLleCb4xej+RTNXo3z1+WHA/6jL1nIFbvS4THEpCHy4rNtCB8Su48mgsd/633Y6Chx9JcgiX
FGNEngChJHAWnLrXV3j5NU3+XZKf30roHOCWgdDPmrsikNoCDFQ2s2by5r/LR7jVUgmS6OK3MQW6
BnD38YY4KWWc9OsuWlD1jCWBraKLBesfN9/omT+4LzzIK8CPY/pKhDBIAQNFWE96Ag/RwiO6z0Rs
cPBgDYhdJztUXIPW0OElH6zkncQZvO1FtKRWFPyRgcqdIKav2K9TCcP7ccirlSbryJRJ7/iU6DYa
4VX9Ll8BLwWJSgHIKBoLM5pC2O1tVBSHljEtlNrXwJfgqcsyYXrynsNnUdnoWOR7pPon7FUo1+6T
A5G0XhE3vbjSnmqjXbdi8Ol/hT797XwzrpIIDWRVgHAyzHXCDmOX+2fjf9sH0rO01270DZtmg8jq
XUZs2rNKtSOiG9DiPb33jlj+9A7Nfh7A13F4Bx8BYF3cWU5T1eeSi9YnZMYoYoYBRE0PjiRGnIu1
xqr16iPVBMEBpc3QW2Wye2FjzXWzfzN28ZcmQUg/vfgiI1eWf1zc3ifsetr7joSwZP+QcJYwbBK4
5W28I5uu1h8bfu8YfolcnjH9C6moLZwQwJGzDJhdysTUspL3xE/84f7ZRsIIV7WrM1hELhAtFzf/
JYl0bbGTewmNJWmr9JKydEMZiGM058xIBIQEs54aL+D3lLjDDKiKBZhe6RNjPs6+7yWDBPccoq+y
S47tOcaXOctLQKcKic7QOgSPb6AyJ6G30fwRK+EahRYudzKte238gjYdH6Drbek5sPLr7F+m7VKl
MUqX9csRwBq1IEXkCrY6PqTgVXqx9TxNh0IkIJ6SE/PR99qj4bSvJDlnyuf5MIqybYHyFUTBlQD+
u0FIjeHsD5rq06e3fy3Yjs9BrNVCicQLdwp78wcCghAg244qeP9X4J4uQxkLJNcJGPR4O29i+3Tw
EEgeFedUmN/R3yxvhyvclZ+V
`pragma protect end_protected
