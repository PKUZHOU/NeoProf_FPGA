// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
1Svep6rNlF9YQHD5UmCTgdT00qeXmiAseWWyALYLfnClzeiXson7wv5j0blV
U72/C2rvIC2T17FcV3YCC6bEUsj1GEdI5mFtDn1Xdt+HLeL+EZ8NX1+ZWTJw
7k9OI1PA7ClwSdTVB2YgrPoVYje64bHg169lu8klndcSBNOrk7dvycOVjvZL
FpqPMmJSI41/3278QOnJdh4bGa1E/FyF6o+TEoY13OUf2Ok/DM7z7rjLWsDq
csd1OyPoTfiB8BFMgOITBugSfBKrnODj0fs5w77jGQ+CnwdatO0Y1TUChPyI
w1g/eJd2Ks2vSra5db6ooR8ziiKmBrI0IqfSjGuLeQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hDmFgLAIsqJuJBLAnHDmWBbICMod4gGoRusU9DHJ4JvRackRYHrSykKwauQ+
gYARO8TyLiploNAFa9NHyiH57FilSAnqn/3hTnxG4ormVk+XPlC8JzUi2AMA
bg7c+TB3b400LUWxBSg1t2X0fQ/P9Tm9Pgvz2EO/PKJkKKR/SVranjedxzus
2IaGTxI0yT1rKXbDmFN8oa+KPQ4MTLhnwvpNYk/KqjdSIahrp+P3+NKQPbrk
Faxa+UYlpNsbRNos5wjAimQG6V5fABKxsLgqa5xkIAO1TSiLI+jzR4B40uUb
/oYGHRAC2fF9k1YHhhhmJd/m8hFxSC2d50fnP8IPHw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O8eqAJxQA5fu/xg1yDV2Gd0yyAv2uRxPhDT1aryGN24wnOuwSM9zsc2V6Wvi
B3xh0orBJkwaxUN53lHzE4EfJR4nMGzoMGCG5ydK6vVpt5KhazFMcm+AkDz9
rOAQMSFvFFO/6RJT4G3+icXd1WKOseO/9TEaU0Zi6cC8QKcO6OWiQCjIwHkN
o/uWje4XSB8R3IeDihMBFibpKMPR/ZLih+gAQJF/7Nv0vQaQAzoGpJOocyId
KI2s22ZtdoS+tUQPWW6BgBXBmS213/71j4AeOc7hXJg+nFErswooWxTYVp1x
Dtak83HMJaHxIQxyNMnao1iUKQCeAt2+LIe+Y7wPMg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BmGklPpFBi2aMjkmHuImFx24Fv91rXdzQaovk5TARZ6NMIRNwxkfGz72h9Ta
jzzR4lJskHKRKnmsO7H10PFy8rnIVHxyA3YSBMMsXfKqHUyBr9yUmZiflara
PaPA8esRjKSoZxzWoi3Q8jb20YmBbnb0ugMoTYd9QKZg+yaqoMg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Sx8jUgZ231HnjPPx1irH7j/UVMPj+/jZGKiWYHthuD0nQ87C0r0q/Kyfqso6
hCImOUabMZGOzkvtDwOcaaCtNGNggX6iDTdTTNw6GQA63Vb26sJZoFrcK10Q
HSfYJ8tPM0uGUBl2XQrDwwy7Q2raZE2iu7fF57W0xV6aoAr+b+HqGYU1HI1j
sgrIg9G7r0JXtk75g2fJXwvMt+M7X+jwwMkc0jD+6H1sNQ+EU6fZjyZ/CLHm
1xNMZsbiRlaeRIWO6fKEwZ3qCFSny/u7MG/DMPE6aHbbCbYgnDwMybRVc8p/
9oppmW6Db+V3n45A+6alxg+J3WZW8hZtuXb9AuI5YoU40CrabE1nZunoMeFt
jSin7+OUT2usXvAD0HhCFti56XZBBCA7zVki4ERhd6rs5eWaQWDSCxOZhXwj
Sx4sLsUaHCCDZu2BRpuJwLuaIoqMPvtrC+C0lg44Gl0z6I9ty+JLlP4tBrXl
JPIGFuNUYtVyCGSVPuSY3FpLKWeytB5W


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J3bE4M+zMiKCa20d9qR6QG/dvswJ/XIDq0Th/4+AtSmw6IAu3ddKHMhn2dtS
YVjJEld0Nb7wrBerLPlO1AcYHV+UZ12qSaaSnRCEWcIZfvywBedPNN2+mx+g
+ci1GLmemXaLBa49J9YmHYa4Tbb4dqDj6/wz+m5Y41vBjGvdND8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ka2XjwAO4LYvRSShk26Qkt6AwzanIXJ1hYwVRaQHrUlOLFV0VbL8Umxbu42K
T8QY+wANnHk/WcwzV3IY+XZndBH8Zg0Fn57dKjbdl5V9ZZN3sGvtyUgaa+qp
Hqf98Dg891kHLxWiR4OBz0Wl78U6hMQkFvZELWFO2Qh4q1LfvLk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16704)
`pragma protect data_block
qbmzqrpWoT5qJboqCf38UmBQm+SWmiJKHYM7f2c+2RCBUEy1WbJviYt6bK8x
j+FDjKCQUuziM8ii+lVVzf0Tsk+rp4XW5YG8eq7vQY+yukFF21JF4Q2y062z
jTX5Oo7HSvP1k/UWiEL9vKjdCvhPr3i44kxHGIxp+D8Xr+s4GTry0vH/LRjI
edXwZj5HKK8K5F4rdUO07ekqgoXay0sW+fbGNIdvQlF7trV2shqhatWP91pv
1R8PKgD+nE0mpnGXa1MaN0EfwIBrWRLUBjSKl5UNufWqvrh+LtQaD43dtLAl
r4aKVz6HcQvY5joapMycOpW6aINZJP/jP7R3ZBBFLZWUhgDrJfipRBa2p0gl
qOkKc9T05BYPVh41lF/azI4hyIQ3z8MEiPH+zBgJJ9eRff1JsQSjnK7TYYAT
aRiOmKJm92djKcMr1xRdWhJBDs0HX/Ntd9rKfbNv1UYt/nWoIEpaCV6tpauJ
HuItBDs+c+Q5ZVg/UiLrhDPUdqMFEoE9w0YeeEQv8RBONpE/R1vpJyz4z3Wc
Mg+ew1I25AQbvo5BQOQ2Fq+f/6oF4vF1TRdybYKtg7yJw23h/P57KQSdlv2u
XunCIQgvFG+ap3jDwXHZRn8TpYNN3R4LTkiW6cA9GkERkcSUsfnp4U86nSVK
0pX1gN90MgY45VdxUO0Gj7rnI9uCZcqsj8kQZiTIQNYVMmER0I2RyfA1dB45
v9k6Vp1724Ok3odKovY/15AWwVEB/xueTJKkJ46CgEIKtTrsGAMMijDAFJdC
PtNVu96bdAocQo0g8kGXcHQ/Q7Ado6m0v44SxjNJtYJGJARopt67YZuDOCGn
8R9urd1Oo/9tUIzEMkMDlgvFR6E64ArCV5jHghYjt2x3/r9wKiZSAQ1sFxMm
U7csdlEkZoFjMJZIZbAo9Yucg83H0ZurHnjkohGUtrSBapWU2ovIY/JFt0P1
ZHigQyhsOduABAo152uvzb9xQYPoAhAvHocRwwz0yf+9q9yfbgZpNsfokcUi
WptHiD9XCQaX476Lx6hhbsccCk2FUNYjf4T4MWOLYxqrc2WYFx0s5gkKr8cQ
kCV4cl/mTpGV3wOnssZThoyzRVgR+FFzdOnLGWO6g5jO/W0gJFk+iXYCocKB
0Dzrs7BxSShVKsrzWkvWt5+PGv7hdbp90KG8I+BlEL6UzAjp2ElEvgpbXiml
cFoVzo4mDv/R4JEE4lqs8jAzk8zdsy7IQYqZ6zOmkWkXn4pM9ySBqiN+an1S
uSUMJDJBPb+i/T2V2VaPm8cteGa7zyWkZxrsNy2FbmMVtc9AplJ9odO/1lJZ
ZTmlnQo06XVEs5R57gO4qkpVkcy+P0SXdOMksZ1wLsUlXfsc5a2A0wKunjp5
qUjkweay+ePwEhXykxtgig+acUzj8CAVwMSQleL6B9BDb7RLDz915kR+sFbu
o4ydvspSRFL/lrTV8yG8NiHFwzloCD4Aj9gkkNbI/FxEynq2TydBhF996d6B
NB/1LFfW5AHC2+CLn6EodQYW5PNRgureD5fWrUcqWX2vZT/cc7pnUmNk58LM
xWg9BBPpTYuzjhsnKe0hC7PrpteCohCA9BCq/Vlg2WMkqrtazBcaleo1MDQR
liKjzOtZygD4UDeVpN0kNO7xlzeWPCU4fpHTtyNaUl4l3lH4ue5WMHw2nctw
ucUVUnmQASPkBXaHVu2RsdSqtdhX6GZECZsIiv/d70sFzV8yeARft48Ez6rY
njK9HqN/ei90gRb05XJE4TcHvG+cmH2czkjcDs1tezpXU1EwgeLIIN2vQc3e
+qUJyM3zGEYgzgXqqXJshnyQ8wthN03y3KKtILOZh5BMKU89qmHKvB5DR7+5
oaKYnULT//ZqXhXE7ZGhNrrNQG66u1OZ6+tjXPExFiWRxOpxzQgnVpgvcqBK
h7dvscRgmWRc1U2fkfoxV2bgcPTjzHhjo/lEKNLmSnB4RfzouCCd9BW7KqeK
8B3I87s7lLgKNp0hsmr69HAbbwctLccqvts4DArfyhnWN0eEwRadmMqKcsQM
Ik1qIIJ/MiudWIFz/2d5TmVtHAHAlOjMCuZcqRaJ2wk2rPSpRydmEyneurnm
a+1yXR2Y1nXl07mgJlOQjot+08M06TpCGkxR2czPfHmd+uZFtQTJLSxvPVDI
u7uAtphQBz00aFqy9mVPZkmSC1RRmcRkVsPlfaHiUHQuse3uDrQlszGqdXm4
itaUjlrQGqe0gW3chYnz2ILNH88D9nJy35lOXr7WSeCgQWksLGBV0zra0H2Q
5m6QsEPy9n+lU8dDzTDhhsaKls86PW3Uxdn0cyQY9mgGpeqktRkXNF4pUcuX
2PHnr9zvYTmNzpIOXzgEc7W3R9h2bawXvQsUVyAnMCy1BMZ1OOzwxF0AZziE
9R3nKCV24NysD4HqG+aixedlqJeyWU3wNUg1Zky98XlN/kJ0ChMQjbQJsAk/
vYBE4JRni0ZirfizHARtI48YyCo5rwOfzllx+niusLPU0XTQhN2n/VSQJHzT
pGfiZ6MrN562jzAm+DiO7bMkC3n7nMZfGZXtKlgJp9W21FfYqN+viLyKd355
a5r04CScTdjZ8rRTr7nY4HKCxWiM3MlSmqS2UClv77MkXBULC1fvLHkXoRjL
m+oremR7yYzo4Pvpmw1nNoh1bR+QqPmjQlp+NLdUU3PgId1R73SBSBBdVhjk
X8qkviTgcIRpTmJbuEQzl88XTHtWcTe7876LULw36aE5+GbUoUVXTSNvkoTb
Rk3pVfg//sj6FFGPsoi1Ll8VKP0LccvF1GSVqR+f9eryAq4FcUdAfd1kBV4c
uMjAELDa+UQdVinZztBmeuYxC5admtTxZeCUc18+I/Xc3I/y//VgPn/HY9Ct
QIjnrKr5sFn+CoLHrtKuktWgMlms4/Gi9uxczUZ885gU9xDXhbhWC2jMIDhF
Ot2PWQcwtiqVt4/v9Uf1CNRS74L5i/lT7cluaig7BB41fanzKQhN6ZbjoKme
G+qUxHKZx9dqnZA7FPjTu3RvKbf8DUrrxxKQD91GbqVI772ZpYCsVUjWuIoc
8McZxDXBcCc/P5lYLUZXv6ciDc1EaAMXFie8mJaJWPkXOAHcvRniJo3VGhcM
8TksVTn2WlV5ZG2uUlXHCBS94id6Fehkn89LamT8nuZqLbm0IPhVUcSsG3f4
zDSdERBisCLVIWoXnjNutpu+0VVGC7RUem3/cF8yfycpfOHL0q3SBdXx/JGo
JaSkxIhqY74unFAn21PVqBuUMcIcS8xolh3gEbGfGO6TFwtYNN0Ixd4LYWJM
tNgm2AftzP4dYM2CwuD53514xTZlETtBwvnsiDseRyrgXK8vMG5sbm9tlbpY
ZUZcLzsA98zVjZwrv2bnVng5YwRRp/rMWTppFKOZmsB5Umuf1IDewx5uc1L1
tLouGOfogjOFjFsg6iKUdDWvG9cB2uBDchBkTqg+PrEq/1k9FAGmVpMWKwBu
v9pGdl70s7NUykJMC1hLZkZoeXGe/ztmdnMkl5wf+/vSjVJajc3MdiVVGucv
3XrSe79yNJE25hXHkKIn0TmLY+m5Cl0F66tp9TqOHBLIRKpuL+CvCaAEmx8x
OqVoFkkmAAR8biWQGYROwDwbnFpnxUOZr5j+Smfn5alG8GxUcJSRzYfQsvDQ
pNUdFSV2PquFFtLd36XkMKgBUCPpWAKh95FqtlzFzKTNzvdKMrU94gfxfHm3
wxBe8RbsAJcFWeJe5JUweJENltHnhq58x4XynNjUotGo+ap0hL9HxHOn6mtx
GDB0XY6hbQA6ARYwQ73kMJNswzrbXs8jE5JLytmOxMDag4Jcj0p3WDRt886P
HRP90MxkV6cCZ4303i5KFIxHGV9GNIvN9dNhx1RpFtXTH5WNvohYKKY3OU9R
Mm3l30ZxNUFoukFg5Il8e6GnCuMhDyYVqR150bzOfMsnm7qH+3GiX/f6X0Z/
m/2/xbrccOB8aiCA7/YqphBEZH93y+DMle+Q7ocj8qEHh8HLN6FLlts2XjEo
nQp3G7DDdbtSzLO1yMtBAYQADwoSbhJiEK0ZO3pRsTZ/ZdDIT2ubBUvNJ7dQ
1BdzIJtKREIxBfTi4sqx6V7dm7MhYU04Xons92HVTybn3zKulWpgOI/cjBQH
3xf4rAZcuVtttdEmPl330C/VUqv99q7HdYxEMyuRr/xdnaOlsPXegyw8jM/K
up9g0EyqUjMVp0EM7s14Gt6qJsqv8GX07icC/4HKaYHOuOQF+5cO2kxZbCJ/
3/hh8TLgmV+8EBPX8AvvsY/iVPp6lawh0r+nvY2VYtxmjscV0FYPW9Bf7A7o
/1H1pRTydg1OqPcagNd+1p1HY/2i9USRMRbOYwSrfp6i9k6iGE+8sjaK67fX
eH9hZt696XjSdX04935sPFDzhs3k2nLf+jgAqGAhyOOnwJrMfj+ctV7vPx4q
+c7r/+QRg3UbZ78/Gojh1jHTigTzwIE1luwTDC3g3Nb8DpipkufWj+/kAQcK
xDzCZPGzRO7lWbHoiMPhkLzoli+hBFiZ3v8w7YMLZ5FjzDI1c83ruzDjxhFZ
OJki/bLiENpy3NP4Q1F2lL/l1bxuc7yZfSPAL0h8wUsps5wonu4t10b6Ysmx
FLDS23dorosJi+hGsXvMdtwW6t9DxBbixxwF5VuTwiMlHIRcFuHl0JETdfWR
gbqQP8tLBqfEl9TrMFTP6Z7sgjDHyB5l2eORy+vad+1RGCC2IPp9jVckvOSz
mhhGjeucFD+p7uS+9b2/fl0m3VfhEjYtjw+IluINedFNE5glmmSluA/ko6AQ
PcJA3cwW/iZO2opK4R+Bc9JmE5Q13pN0J27/ul8aqOjyUtvBiHoKtO+dV9mg
OlhUge/cXyvofSl8FO0RHa4rXqoy3KM53xeAGNGdeSc2/sOMt1/0BKpJY+Dd
CLK4hTyACR590KiUqHaiPimLTA7m4RDtd6aaZ9cm8F1L/wUyQTPMjeIpDjUb
0rxhZUbGGzPFiAsPLbGHSW1nX3NyqqtRWTw6aCHdwg4wWdGePr71lZhNIJUE
kWHuuYq+xER2BbGl63MtvJK14yYd6E93ppHb96EbQbwRBU5qEcv/vizwAIRM
JsYAnQq10yA+QCMu9PZ2X8RUCcBDqo9ERyriaKC7lIfcqAD2LfLE44yGTzKg
KCCXENskZHu5HkIVaFCxJGKgGtJpiIJiY3dj5ICYCVL3BveshGBCZ/NEkiNL
k5QgN7teJyJxupAxonrR7s6WOoW20b1GQP3ROcw0psyqsQ8jTocLWM5lSRoQ
W13OTgeVnkQMSbrxIHVn+zo9dDvUKQd658ZnpmDgC8Evsck6nIN2IOdKkkIo
l5C+IdkdBsSKmuRjfrOiJXED1NET/5tTG/qvzpK0e6XmCIxx2fqRdvzd0IbU
wZjoYsvrjTOjhu00RO/BTqTjm0uV9FT7DvbesVfsGP72fIJDq1RBS+WTBMaS
PUmaB9SpL6X1XICDzDrlL18aaSS8rijyR7GPmx+ZGffMftbfZsHrI9Y8C3GP
h/fx7rQJchOUBXjnNrhMP2Q0GuDxsXDrKHhnrUK8CCZB4EEDWES4knm8Xs/j
lLdPoC807XFHYvvRo6ahxlORozXA5LskoCoxvnkJi7Z6V8/lf6uSNIfXXquD
p3clcoi/qwD0kKIcYtqO1YKThOciOoZJ82q50dAAeJzIk6NxyeKFrTnnj3Kh
YQBeIzE0Q2LLvUn5wsjazN6M5V92k5uYTAq7mDw2ilClgpzORMVBgcIdp6nk
Jt3yJAufXIL6QHSSaeitbRq1tzp+DYHeje48lFh5EtYU796PPBLSLb6ussfH
wT2QaVZvQ+RxLCQgPQdqz83llbuA2IgvloceK4ThuPpfm+6i77zeMUz63Z0i
iOybb/LHqKCdk7me6W8PT/cgUKSeCxV6nvqYszWDQWcTOYgLKcd6Ykz5qHCi
q8eVFYQUU2mM/amwzomuQ3C5iD9OJbLWgsG7i6PiLQyhmwM/QkapDmonocrp
m+jWEzRQlC4ebE1yHmFKvV9A9wm7+GIgMlKOMtWalmD83u7uXyDR/OzBS7/h
ssmZbHT5gCed4ukJDZxG7z9DR3Mm3pHIhYRqnKb2rFcuh2CRozU1ffpM+2Ny
iOMgLIucG6p9tzvRsQzn3yl76RM+rNLzBdaC6YrSnhcU0H6pZYLKOvzFc5wF
rPiDNIEMiIEo4BGfrMvGXa0X4pcFcOGpnaoqHtaJ0akEJtmUvWUV3eDa5aqy
H9yhhJByamzx3t3IEe/naTdYZZAuVdeiOVaoPoSgwKaS+vFQpYj1iKk9Tfoe
swWtuaojEpqfNhD5ckNunb7y0IFCRHW/VOlKrVaQCUWs71639X0faaoiOYGG
OoIk+aCLzbLA1RF89G3/3phcL6SDWDe8/HubrME+rkbLzT3BHwk/M+2AyPhq
HCnK/YTzTlSSmpwMCLTOrk1VCxFn06mSGTsheL7oxZid9zEhmH1txuXtWozq
OyIkiDgtBBQNnWkSBSh3ui/jrsPdYYNiOC7+YdvX0vd8/2DdLolj5fPhXpv6
tei7Nd1HgTm4Vz18bQ97jrbJho7XBj6qTB1/smdfSCOilDQxHKt6pIBBTEfH
oL94QK4qMDXq1qfard2h+vPQZTYw/pn0+2mDKefiDuVsx+k4PSAv6VnVqiBk
9YyGLHvcCS8i8UVH7VL/0NAtn1vaOH9CmZTE5F64Q6Lz66FoxHPb5SvQYFoR
CuuTM4KT54nqS590ipC/jzipZLkfMlfNurRIDQZNJe5LP7cvo40bnOTvRADe
785IOlm7wPO7t4LK2t4MubyDW3+qDFkJ3Hy+fjT6Q7PIRksK+nEdb8D0q0pY
0rFKy21JsERzQu64L6kAQMj9vW1TE67HVoiY62jKVrOnGt7E+shPlR1OnbHp
XBg6h5LIp3+qJ7BnW8X6pZYnCgastUh/sU4RLo+JPPhFtLaeyuY7HOUTNPvg
dAFQdf++cGOW/p12s5Y+ab7/vNn39Mh2yV94Z4rufDiErjRA4/sAzN/tKrfW
PZoueJYt/1vLI3KOXe9F8CVjmtN1wbGrQG8GIQJGMnvzwCt79rjbNys+A3nf
xPE6xLiGlLq2c+fO7LGL0gE+0P7XOqNpMPe9mdsbaWrQIBNW4nGNu3Wpu3C3
j3Sln5d9saqszTKz6jA+PLp0ahUabkYssZT50WlJTkdpqgurQyGn7cc1N0Y3
w9vmm5qnVDfzuQl3PmY+FEOWNNbnHw0bYEok7s7WVI5HYX0cXJhv2i9Jd/xc
03nQWtcNpXZJT6E2obonJczJ/K68wTtpe0yoZb1Ve1yNUQ0XDl4odiH2HqES
ctn+OU4HZNFsYRL+F9KdsuYCTPOPrsJkkKOA5GjHNqBhKhWFq/GQ/y3Zh9CE
g/XyzQUfKpAW5T5ED5vHu0YT8DT5gtru7iAtDExvGsfgcylOowTWC7Jw3Qgh
5nyVkuq6fipN94iLsDCqV5flxipCAayZ4j3qV/BULrCa6fDFD8oo2n1nyz94
UdZXjHVV33qPykKM4NrD9z95/r0vtXP6hjrseX3/g1fjI0fJrYJw7Gcb4qYQ
Z20cVtgTKtE4gFf/hLosRAdbC36KkCQspOqWE9thAm22l+PiWThy1E5OHXcW
roOohh82bKHRxlE5jKwpjdhVNLjl9j0BMme8Iha+10ixd3SKjzVi1T19G362
c671e7aWM7mX5qRulYr2yiki0pk/WtqCGFQrfnqRQSEvwvn6r3qtSpeAjCqC
jwgy+qU9OA7ZJHurro9R46Akv8ei1mx/AVmqIMXpFdH2StG/9esdMLFlULKF
Xsh3M7T49cdRK/na4hC9xy1DPRFZnUNhvCDt5xOJvIw1qw8rpfVvc+0MxvtL
luLendRWzQiV1nksCfuIYqUAb2PdL4FdtClBQXM2LSBxL9GZGILY0B3yR9eP
iLJce5lMWyGsJuozHK4dZvq2hGjcKPp/+xNLNaChh6yDUVUJL0ORRtlkuXpl
Jv+zFAojAMMLMycGaU7jWgSC4LTXR2wJDc+y18ROVGmqPp6zI5T22DoF9lzX
QwBFNw5FuB3Sn++JfK12M5rIX2dfbiX6vm4p+mVSoEjd5pce9dv7RqZuZdP6
WseJv0eGhg5WsV+58b2h9WotByQN5yuD5fC8/jwn7912PxwpIGSeNlgOeWug
X1sMecRF5TwYrSq2aPZ6aGKXj7WeiIWTUmCIJ7mYUIvJmeH5mSHpFT5qruiX
1t88h4ynHlN1D7o/Yx0hj9Jwpa9+Aav3GMPqis0hUvVZvupvvaIzguUeud8Y
h/r5wZEiDRSuoqnia5oTTs2krPM05+50AyFgtLlpjK/GVTivypKI0Je/YFQ4
1oaXaOClCrQPQZEhZ9LZI+lbENobZ1pNjrHE7s4Q+5i93bMrRRYjDVd7sgp3
pnButExDNqiAVb7mOvjiL7gNtLK+tvulJjHtLwmo2z9Lb02VcZf05z/D0AFk
L0mpQYe5+WcpJ4Uf0Z28W7RHLBACfa+XQOgnnp/OW20/sKzd+xLg/5YST/h/
3gIz5FqgIX3XoAFkXZTgSXBcDJ/9dxRUjdvJebJTwaxOaoT9AUtHvkg01oMk
/2dMay31RdIKXdnVs8B1txOXV2OdKvjsR5/0Qm75Wi8zAOVfZD8SiplgMcx8
w7l8lsV0WDFWZr48WA66TnX8yvsh7hcM1UEBnHP/1HkAsB8kJwKj+gYb9hwx
/wZ28Vw9cnzWvCspBMSvC7yzvH03FuqLttfqb0y9PyQfYYFjLHVKAb9EQFB2
tOiRyeJiMpe7TW10UO+Uldw/g7RNsX5GmDT0gOj+bScWwA2IziBAbJajG7Tq
1HhBv/QpkThlMyVkt41v1VF41eAy7ppRrLrbzOyER1sWA6CIXsu/5jmaQpiW
S7gwz86BwzyfWQl058CK/VnR2KEw7oxGFrhJSbgTH0xNeoBn8Ei/0LZlQh7I
ftwNqqNYwweHgs3YUFrWPQ/U2wKZFJgU1ZAOSwhTQfLDLmd+HjOzgZ1GYH/7
wTlGsESkcOSOrchQ58Oq6CHI8NONA5HG8xuivAbi1ul3PdKGgfewEfWrLmB0
7ep4Up9nJmXkqVnEZ0RF1CFPClOGQSbGiT0Vu9RNRee8Pn7xKQ/RHz8+DKtY
soV39C9c8Q0mNdU2M4t9tyqXgTU5bnqk9tv5PzANT8fsY5kZYzud+0eYPzhW
pUIu2a12/r9xG0VhKI9vEcypaVaMxuDp3vEEKABh3FDqaFQs9MKP/7nM2seb
pv2arjnktX+vd23ZhYcYHaWrhKHS4ZVyQGBWptKgT3nLVBF9wLHdLqMsQkP7
wJxxh+PEMl7hnQxNKsrFNbcG3tSA0Be+5suWZ8wndBE4D41rtGtVt3Xzwsmw
M+TOkt5I2doGIy6fuhH2zIJO3o/2/o0cU9D6uVkfar/qclmlfBHaz3TkKEUK
oUtVSRCQYx18HxFtLx5kxrsilBq+IOqETxaQz0yU9OXO35E1CX25lflGGd9w
yz1jl8w+WvB/i7a+O0Rb7i73plSmVRqN2K4IXn15Z0FeMRVHV6IdtJmuJAAU
AzCimgUA7BG9vLJvWkbIVkLb47U/irmfyJ2QN/tpCJANZmGNfwt/OfnmfGm8
2GKmoaTNX+msCUv1Rl+J8oY60jOjuGspy/SHTsu1CSDRU4slFEdWU2d/wE0M
9qYDIrIgYFCzh+EQbWK0nXzIbKGX1Hl2NiReUvrkp0zLL59Pj0wQGxuSjKys
9irDscrLwe+Bp1WecoKdFzBUU18ATnXBsyRU7QkIZf5uTB1psUAXD4+L34YI
v2Vb6U2/tWXMP28tDGgEQiuoXYRPImGhgWhfFXpE4ANKIlLbqDzMi38S11PJ
8c0936dam7Us5Z/b5AvHfr87PlOpaErNofBRnbTSFwYGl+oJApiJdZ1Dtj4o
+xhLUDo8ScBDOmfZSEsstoFTwhcGUoxdUM0QzsgoXgeGxZJ2228NteduWDHd
TdZKeg5NOCFOpf0BKdJUQtdRUY9kQJnijcxVWqwyuqeNuDA/NwRB7CsE5ZFE
+Tj6lfkpXiwwyQ5s3PLdZITaymPAxO9+3OrcBmET0iRLDPq42vVBO0DUaJrr
hZUz9SuTbp0KSxaEBFITq/ZwiMohgwTX5GG2Nz39EGfl4yzhWXKqDfGkAuy4
p47gd7rKHbnttmQj+dlWNZJwy2sIzPDxoYGDZBE4tioRMtGNKwDXvRTwKTsK
GySTPXWhK0m1W3dU5FJgS0xMVatyNu6z7YKxlrDyagKCO0R1rbY8sJhlxRKL
u7SlzuIBq+1W7LscWgWBOmnbjOwx7ARb8Iy3/Mny1XOj3fR/crSceiwrVRY7
n6KU35kCCzA6D8p619CtR94is7a6YdeTLVz9hRmml0IbAtq04bo0PYM5AivL
GnO6bazKdXG9auumMQQuOKhXyifcPP0M032V4X9D2TCM+fu8A1L6UfPu3u1R
gMbbRuhlO8fe2wioTMTAOvGbcJnlp0MRv6CdyPgOiJBbVXDHj40sAfg95+kJ
S2QsYN3BIYjuOy4Q0IC+IbrEfBPIAp5rD2pOHSUBeurLuav8tVCpxmwkRL/D
b9ago6yMq3jnbMtcsdhJG4JfLTpDCP4h7roGoo7Xs275P2DT14bjRlQD8yZU
Y7GBGhsfv+I4zhUeCAWSoRiSzikex+/Ha/EJ7KJh/yPMAIkdn//gjdDDYRcn
Kj/vQMAMe96r9AaFdpA+X+XAUHCjP05EQZ7+B90FOJ2dg5v+zor3inqh8/10
b8CGFbesLwIazWhIJfcCfEZ8MqJ+VAdDNMFJKtLG4rdEdvy4KW5ep0Zveb8o
Roh8pFSBv5vbHy9PA2KMxi3AHLxyAfAZvJ5YHwxethvxOUzkVR5z5yTAYfY5
yNpKhPFkxAHct5B0Cabzx1lxtFy0gImlAJmet7VE3qh7qfSc4jj5jiDdw84i
BfGOG0CtLSR/cRSmRThErnBCCKAUxVnJfES3+KlS3uu17ifUHJF1RcDKB7zx
IXfS4Sb2NCVTJaNDrnNxVNcia2gPNoeDFbS55Gcn0TUz/iAYmppbN74vHIqr
9oeDYGLvvV7229gDziPhgDu56mXe7bhFa+iordvTBeGvDUMOCgxmc3IIh3Y8
h0/uhQVae4zZQhnlB4+fEB5Oin5rqBED7xaPJ1CrDftcqagPCp7D02Xk8o1l
ytMXFra8wWQT2DgHbCv3ycVfFdDDZcUWbnCL1Ip2/XLh7ZGOCyeDbzIJpTqk
HShsRTda4mTKb7SUcSfUxi81is6DqjrG8ilFgcE0qFNhRrFtw+67UybD4Ycc
rZ1l7fiHxklXmxGV6Yiya+uTAjqFnMK9dqJ0bgvQiMFiicPe88WsR8nl5w18
nD5/4bV/MtDfReUUD3B1KtQy9vbcqVgI67aqxeTBTD+K9pCB6x0rIHVc0zc2
Cna5NpWY833Jphs1syg1wuz9oYJHn41cXUA1JIl14GyjuBxa1HyQjEUTDlzS
rFfY5d3AKINkFZJwn1okMW/9/AN9Z6+CpRwMXUgk38i8Gz3jF1KwpnbxE7Kd
Nif2JSqpTYO84gsV0ZlzgRYvSIsjDuSORa0Q6xSoFZ8bnnG52lfqI3N6d4be
espnbW/h6AS44tmbOEfkgVkaRVjS57MGR7o48TsWikxpiAxQPSTT692U/4+q
e2zuS4UH/ZSUeOg+A1Y2s/4sH4vxrV1bwxCNXY8SYGqIf1Irsxwh8Hn9R0Db
Nd7i91DOZI3/J/pxC1ZJha0OfTL5MdUc85gRvC3NiBzil5JfMRQpXaqQzEKX
nwnLZZsXHh/tbxoTYm1lddL6ezHRkmVV4uDcmexPZA2CHaNjDcuBqFlfH3qZ
mF0D14RFAZAo1Y1TUCjhcajXcDyN4IFoD5o5a3gpX73hA/7RpHTJUTk5fs6U
wjdszFvEtq291uip5zg6zftpqgPutAwQedhNSXJiSicGDDN8ii2PeIfFRUvc
agXgzrGTe1evGu0e2hn88cq2KVxlqq7kpSLzXqb9DYM58ICHJt1GyBuFspnJ
jd0mqPgbr3qjNXehmxbLPn0HJhx4i4sYTZ2b94xQa9Ohc605u2h77kVLj8YF
iwFVofWIXvHQd+oeERABo5P5zGLz+cVeak7GF70+2ODdJQANhtrknXeC6wEK
TR27Yp0AH/CaqteMl/Vn6A2C7z+tu0y0TQIU531mY1knlY5xRWcLv80UFKWG
WN9ZaAHPmjQaRDu5IHO2rAsSrb2X9Xdb7HnDV1w44s7VtWRL7D1sjWDCYQz/
tLJvRXfiZWWQWi0IkKLVVzwmx6JSgz0Uxr1JHQ/HTPZWJfY7hoomz2ZVgjL9
HoWL2SB4jeSm/tVVmdjZCrscC+6+9Z4y2dhN6FdsjalVAyy2Lcg5coeiBBhi
gFQi7PmL+v5CUDyf02utvuFDkAUGzvvDBXO8nGHkO3l598svY+/92McCeP7U
WNN6g2sEwyTq7fFi5SVZ+xs1ccxwitGZdGM1gyz+Lwc4wroZdL2bpZ7RFkF3
ULhKF8G/tMUR8XM587nWDJTig9a8HFdQSKQ+1VXOXRX9gHZCxgWHfYvNhru3
+29U5p/owAiDgN9dR4Gj/cst6QjuHJL8E0Vt1nZErBnkW/exG+lOdzdEaIad
NLsd0rBDl3SQEXwNL+bLk8DJCyjDiiW4tzqNLLoLV3ARm/DJ4K70u4C60Fce
740O4ZxRb88GYA/NiBy3q0uoLDIfLcpJOhbESfpuL7FMAXHfUnIsBfAOzvio
UaaUtGIX6d9g8MOWw2AZUtEV048K410yk1Qpx+zRWhC59EXNC1Ik22jidCiB
uFLwVSMx93f0UgikTIT5nynmx/NflGjdT6DOrZoBX/Ekq7r1gh73Md1k2czU
NOpgc8lpBGHHF84nbncgalwe5u0oBGIHtcOy22u2oEgleQurwmRGBu8RD4ha
HtA2YnpNQ5i8MlKSFppeldGYJ7hkwHHiJlrpGh3CMUHrEZRpXfKl1yobUMFI
CygUIjkyBJ2A/ZM3VpcsYpMbPo3179wt/o1FHTuPYq4hvSATCO+HtzgC8bpa
EBlV6FVoVWFNivYu1/omETf21mjH8pbLuHGNbh0CzJsbidhqqEbh8qldmLlI
W06Xnb25YbL45cI3BsoyrvmoBx52usfr05nfNvJFNZICKwAJxE0huM/X2527
p5YkOxR74cEZ6dbgHXloulGVK0X+4oXSgteQHfuSr9fJn4zsjbIaGp1yZ0V2
siY4q4o+/oVBTBFj2jl42hkkQo9F+xBTAWDJRGE8MpaoEuRZyqVSYZsZc1Xk
WfmQBsDfLEYL8UeC9VfmUp+gcvRnFV1LefghSZzUE2V5Pf0eARlnGqk/7OAy
A2sjIP/govZmY/bzN81pGi8MGnQmPKA8X8CLKj4WgZ02WDyRys8dk0HbASAi
jN2anjk3tDkshx4NIBYspy4BaOsW/+bb4kZsUZI05pBv6xdCBmOvKl8Uar75
oZwC7+pqM8h+19dSU80ZAYDAGXLRZAxKxIaJFmuJb5KoGK+jKOwv24a8FTMV
QMHti+Q/PFmAaTYJFaDfjz1Iea7Vzyt1t1SKSS0nZcfmNzUAbrA2BGCBPxhl
p4JRdnQmczApszNYam2wNnN0ClAFs8NOb6LAeDh/i1MScpyXg0rp3yMQAeZv
/gH4bP0NLaqW4SiQj8DwhxbCpsyVeOxPc7izl52SRBEgpuD+L71kqgxVkzmN
ObpQ8P+xsvhBZSiBavXr6dTgVf20H1YFXhO0nOyi+fg3ouR5Nw7TDuBM0KIV
pQXQrMQUi/fTWGEc3dhk3aYgFgJX8nvOXu+39eQtzlDUkQvs78tzgtWXIoCe
Zb6y4XbPhlhGcs4iA7nwz8tOiKaEW2F+PxUUl7b92RQp35wHKioOdgYIAtbB
RyHmpaDcojNHpkeXOwu9YlnOjOgNOTPv5iuUMEgvrGzHpuc8fBL8J0EyyLCs
nXQAfhNjd5CjEzf0pHw+77xueJrEkZ1kE/lOz3SbXgnXHDmF6W3IOePysPXt
5qvMRK2HPHyBMmUjF+OdutFvk/HSyESd65qfJbrYxL+RAHjfHTHwtZa5sWBN
CgRjD2ARq1zPLhPxszag1kwr0j4WuvwVbuXVUfPBZdMXZcvKvvgNaitP7H9G
6Gi4X+cvxjzXLf9CD0TrZI7lb1OBj+qnIDY2CVsPWqBIPFiytmbYtthEwmiD
U8ygXq8Cv2ym5eE8iltnCZ9+xsW8SL4QUesCsxt4kOwOUWhco7zxMXbqK+Qw
tDj+GAiQqy5oT/uE/InMvwNQhl3ehl+Ihk8U9Moy1mr0+xepPr3hMLvq3e3v
anPLucMOiatSgOpA5h8eTqWZaDQ+FtUYf4g8gakmR86zC9p3po6khPc2gRxd
NN5ryyCOgsr/QpiVa4p7A0jrTFaTF4BZWg5G10M2IrsAoHnDESaBx+CCHsil
n7/xtt2JxmXUcmEU4JYJWd24Ehhku7oFv9bx20tP7FxoKc/dfN5SJiqLTauI
GznsH5zkYJn0sVJmvkTWq0jsLttgTaT2N8eeqFGUD2gketY/ZutxwyYwzKAm
G6bgeZEmou6Sa7SBTjBzSoOwehfFOM/eS7Aef6VVfT+BImKCTGNLTJ1jQFIQ
kzpQcgARpds/fmcYyB49aybUF2l7ZVRpjHbbq8YtJjsJQb6FErUe0DnxxQ/2
Ixx8z5hTs+ggMRrFFaRVbp24MY8psPiQu1rjLtWdefBk6A/9dpa2cGaxJa/4
MWwviqAT78DmIdk1mQOkSF7bO/hVX5/W5XLZt3QUPHAAXxwlSfNTkiDq5RY3
arSP+RUOU5ZRJRcrpB9DvBc2vejTOUZgsyzsbyiUb05QEeMAvSpfagRFlw4K
CJnlTebogo0t+oO7baHqzoDf9BtQYgy4CbpHvuXd0zL5Xrx81fuB/UZJe1Vg
aOMUKYoOIgEr2eOhLlaTBRMh2HGmjawe1ejrSGsqNN+0YuaLzWAapu+/RsZU
y6CDRCae8dKTSljWXaqZqwCCaWV0eO858qZTeiKHY2Z+o0w7cHrLHvQhXCzB
anHBCzxp30NHc9l/NtKM6Jd3PFp+Ohx5zP/2gDrWqgpqAluEp1RIqdSBVWQU
q+B+ezxCTQZKV7d/rAjclKGroayrPXnUDFdS3v27UNk+spRsf4gC+OiDU3mt
UfQgDnT48VKOS99x1ohXhyY6IHm5E6MriSg5VpoldmYFbKGAkUI0LGTfh/q2
mb8zq9ObNKJv7PRL/ASHKRbvedPnrAbi6mF7FYu7d9I6rdajx0dcVyDwM+1E
4NHcmKZWQcbQyCZBb0kYEt+UvuECw/T7w0e2v8+jOOrQdpymluDCWDIG4qB5
lj2U4I/xZQ4EUXnwIZTBCS13btkUKaTcoyfm3zKw93CD/A46ZVwgsOifosQ/
SPy5oU5gR2ZctCBuCrsfdD9vb454GlP/vnCeYvTVNU5lB7pYrjN/SYNFAFkU
AYyHQWzsgcg7B0DPC7iyYqmMcXneQLECc07TXbqr38oklMKR407iP0Ce9zFn
wu5UEBLmGVTo63rBUYptKuRFmMGcYUZwHQ/vVHkpaWuyO3nVQ23CGxqRQ2/h
BQREGwCv87GwLGvNLs3RJv47TOCY4bGvbsznl5YNR0S9zF8ry7R0OMVEFXjS
4qEfieFx2GmuieRHgvwFqhf7i4TAXve8b32EbCerQf9lXrgNPDywhE+g5sca
du0aFoTUrHPo01S0OVuqR6ScNpItwRdwxuoQxx6FjgmDfES8uc7naPVfl5d0
de5pxEPPES9ZuCvrRzhuBOybQMz/3phEotjTzL/E6vQNUy/dq6foJ9g+WbQV
DsQO7eGgfmdZszR40k/SNAxTme+QWF8zZFtBLn+Yk9C2fUggTA7gXbgirdlz
czXQHXGpaGgNR3KInnwZjq+JN4z6ZM3HiGUwoXsrWIMXuadJYXJWeOMKsTjQ
sv0ZXnHYqDXFH6w/VomaJJQM9px9t1ZD5kAX0ph0SX5r1fmpoYfe2pg4Cou4
X5mfST7Xf1ZAI5fhsHehZKTZfHlkn43nrqabRPXNHlU/vlCRKc3IppuMIKCq
Bky8TO31TbuvwWPQqWLCzuti9O7s7ny1cKcNntUtZegKn4AoqnCm81fTeQY4
z6SEu7qRM919ZPyY9lopnz4CCV2wJ8VSQ5qywusPDZI3LGdivCun3ln7vukP
JVFq8exuNR0vORqElDG9TYumLTpuHRVORQkMBUg1JfwvsZHOj4xa7/+/WyKx
djo+iP2k9sTKA3abvyy8ezyCOd+fxs8D3eHOumZE72xmjj6jCyQ8iK/YHbjI
napevG2KkgfwHDd3xbkLwT/Rg6vRvHKTs2vpVZlRs5obzHDYOVma095Ri+0f
tcA/+Dzqa7pTj4+OKdXCfqWppWIP39aLI1XuH/4/SCEWFKgXRfrz5gn9d8M0
5u1Qal1dLVYR97S0CFMp0P/NApfGjOFyi9PI4+n4LkKTKqrnIXWcYOBbiJ5S
YQUaXjG96VXXtsCpYidh9PvOR0AvUcq19aPXw6OSfojqVSbTNzbnKcYjYhnN
56KItKdtq+jRBWz/R0rSmc/KOLuGBUR8X3GisJf/E7UYFux5AARPG7kGyEdb
6YM7AkYydDhtKfxom1W60LlcNprN8jHaIXrczHIXzA249/UeUJaejrlIHNlm
wRqbgLz7y3FIXLd8F1zpkRBlQmQ/jxx35Yh9/G9MMTRpbmbPJVHKVihx+7UU
tRkQurtTQvJxxlPYumw+CpblSm8VhIthX//emtE7OdlVM+S6G/SqXptSTW6l
G65CtEoZ2Q17Ea3O30J50HIvN7cDoCccMHVNj1BWhyzZX/O8mlY1kusovpeK
HQxOtmLYle15q69Hp6iCAJ8fAZUP5B7/g2c9hkKyg3ffmsIYpqHxYS0bBiC7
DfS7/yt+W5GnpH9lLHQJuqq0W89PwwqzG4lXgG0z/xaYI7SyMfmudEo/XE6/
icJN0xHeSvWGJx5HYT3smOh1SuWLiopTmyUpEMaOykonWzfrAefZegt3MXgL
oBGrw7MpX7dsVJlkfo6OFhw/OAKNiWesr1rDOPDgHe6UjMQr1VkhwtxzhQ9k
gOxmg+CBOLA48VLjVTxwlSMmm8rHw5y4vJq1Ysu39hw74kFD//LrxmXRNne1
GW5CAIsA733V4lQgYduJbEM73PbL6DytO5IdDAvh8ObwwJJb5WxtL/8s+ndg
+0WPRyZgLj/is/fU8ySnVdiaogwwygIDKvk4UG1KNVN/tRk9AbCoFW7pNIrZ
71yJ0WfqWxvVsoEDNFCP3lQ+wWFxdbmDqYOPCiWcriXPrWyA7pdVxak2UwgE
S3WXVfdWiaGVwvPrASWDyLjHxML+GBVp7pQ2zgBJLA3f6H66Qy4Xj2Lt3Axi
1adzFC/PbTQb2VmmBNUBCEcb0n/1Y2AxcJaFgSrrEv7TLSv8FoEGH5f0Wb67
acClAedon6vmKkWNUkUbaS8YyRdW8gh+53HKcEcevpfF0y8RCJ2cmxVgV9ST
nUloT5SCmhtw97B5yGuf5W1Skct3uBpNrtKkZcY/rUtUHXpDXTPkkBEkoPK4
3A5W3E9z9eIKAFCa/0Ul2PSYN6TB8gNUlhQI8NjV88f3iLWSqs3HqzmuHBck
L+o8AvEiEgJuGgmC1gDZee7SF52qQNsGOZnjtf5IJAuCMeF3xECTSePhS5TC
XlFcoL1bbZvxWDhHGS+o/Mxo/AVGxvpwIlLA8RtVZ/qLERkw87DTdPoD/PON
sXbCRnq9aLkDvN6iH9rW7pnePFpmIApjM8mzvPuJBDhAWsaatj5R44f1aOGM
cNagrjjUUduruMZdubOAuAnmEVvjuiQvNiV0IjwCw3vfjerR9WMqNeyosKnT
ftDT9uA9qmM7Rb4A91MlEnsZBO1BT9P/O8G8D4vHGpMgXJ8DGgj1ZpGewea/
TuVbinqnCIvFUPfUhVo8Kv6+2zShtZDDZXw5UxlpxXl+u7iT8Kgsl6w7Ru2t
U+yQ3AN2HFykZn8yB3sLCpqc/G19g696xuDsYEazi40NyOOMeN+rtDV0QcEQ
dkxda2IfTcdHbq9rRbksk1QXrpiAHGJOFz5LbaiUzbqAD3NlKfg/LHSzU6aU
9grf7PJzYVzPj9l1yAuWG24cQam6laa+iasszGqs8TvpoAsxzJw42SXCpC/L
phL/tTe/CBlclI0cTCSnE0inOdWKASVLgBKltmIVyM3NPjS3+jwSck5oT75g
wn56QVrvE6CNWnJJ+1XUSZM6j86JUT9QylJOhT2Uos/sP4O5OG3Ga3NvJYKm
N8xW01vifKund3NCA7yIMg1Y4/s1N/16vXCP//u+JV16bifb0RHQIPrLl4FW
xmajy2ubQSeRjzTTBLlcpo1uc/8WhA0KcyuBwYKm+zNj5P4UpYSQ88q0yq0m
IcKrVyTSQQmnlmc8TJi0kuUddDQZFngg5ajijPeIHT1pBZFvmTibpNKchf94
83Ooo9/tfUCZlPBiz1UihM/mUOvykx9FuGgVz5sfQQlXroL8fBb/Q4/+rfeW
Quud9QTo93/TfwQxU83Oyc36jN4fLqZh50SrtzGqy8MfTeIbHg5oTuyMO4PN
6A3xoVgrnQUVndWmQPMded+twJj/qlAwr9rY4E7xb3J+n0AFmocnp5yBWh1q
1hXeqGq56hg2zNXWEGmxn6O25LEX62KkfyQhNymc823Zqod9on3Gu+xA+aw+
+3vZcvMSfuxSIlUyzbWbNKKMt+Ez/GmttJiWyzsPLVZkFRx/EUgvKLtBpYI4
wc9EvCB6CkuaquJmUSmL/uwcHJfbz/sEuv/+NTJgfzgjiLxYdxYosAohc+Qt
t7emDqMjK1Km7Ry5F9neu8P9N2Z5CO8lstS82O0cOBnceKG+T+c9X0Clfb7o
Vd65lz3+AnkoYx+CijFJTKBVemykIP/DngJEZvVS2kriX2AfTv3D4O3wlBIp
rZiq8ZSQcNE1ZH7swjJg2z9wr9hBYlBYgNwMJY3ygv+Kg7FCbY8cZAsKmo1+
lfbhLytlzemuXcnT/jYqu8L+wFAqTrZhyrZGNJE1E2krU6t48xgn/4gb7Wy0
kPgGdHPRpIRGj6KrfgWC+N+Ezwu8TE72xege5zGT0XREGweCJUn/yLzZhiOD
zWpkSD//kJts+aaEIeQrkdsk8K9C3yPgLsNWVF1Xqt/5YlSgUBw3IonYQe+e
/XBa5slILGNTi3l9LQ0NAgjJpPU5S8JHKISwPVpIzPc1aauE4y/yjcAJuNiN
TqY95vG0AyaRDHEKgGArA6E36LpewzL52uMtvkeBDZMHKXCoQIBnXfyl7tBs
WIL/GbVBsdNz3T8XGq1JydWqYl2zD5a538rPNAczHmB8bj2AotpAypj0/rkZ
qBm0a+PGTJoyYfZ7DFPeQGPSH8PvJbubZvT9JtzcmFxzy/p17/+tG9dkwjaT
ZoxVQKaLgeMrdh4h/QwU/K0Otd9FqBIoq7cw/z/XebV7tQeSkmsxlyHsWJYX
culIkchmQXOf2V3zPdE3sLDOHiB27NmNsJf8E6fo9hIm9UxKoiyoC3eI9g3H
lsME/fRUtUWAKEMfCQErfSWsidvTa+5GLfL+eVd8Gh/oUFrk+x8VG2iu1Z7E
GpG6tCXdt7UdGGoB3mrazXYmncT325xuL3u0uK6kG2XZ/Aj866nZNzrnqyLw
LIM2JwmwG6E3qqQSPaCN2v/P2K9qcX7tNyzBpyADlArXLfjLo/iUPihDUO6p
LMfdZgOLIKzils3kdaJjhS+mFj1tuh/GI8GVewkP8Lv52M63LAIt5FvlPZk8
5BJDtR92iS6bHzpyCgaxLataWMTpHd9ucYsLHnAZYLlUp80QvNJPh+j+FRx0
I6B6T/Xcr2un/E+OMjWXvUOGXozVkwgQkD/A4p69QeaIxAtB4IR2ytskdFQe
f9GlUWo4j0lOI+VfiJhQbpXqX0hu0ZokcP5JGXYH9r2u+5t76uUGNIgCHDhT
b1Sr0X/AwwKEZy6J0bHNJCBUMY93ojL8e9xOWKm3ct+0IM+vqbsG5LYJYu8b
sF/0HJOEgzD/r475/3NWe4p9EGUkxn8vUK5u9vZsndr1vPWoHIrx/Khs9s6h
c+kuboqGmY/c+7+h+kgKypN2QsQQY+uAFAqemzw/CGq+s9AfbGXITdpWkygW
n5VweTiVc2NtuVrKiGVvRrbJjjuReQQIXCFkY20/0iL1FXaF2yBL3YpaCECh
I6kG+UQ5AUp2NiBfFlHfDn2rSP7jo2TDaeg8cPZgJ8cZ1px159FuOffeV66n
JY/8xeNiZKVOSyq5qWucYJBkZNipq4pjaqXbxwD273XpMxeJBVn0YIFdfX4d
3ls0Npxbrh10gXSMpLPc13cu2nEOwMziALye2Zw8NROrhaOVRniFLO9hnQYa
yPxbe69+A7i0D+iQ9VLQttFowdvPsTKSZ31c7DrpJX5CQkaMs1qvNP9XiJwu
Y/CKvU5s0zKi99q/Y8A2sJIPcSQ9AZvC0pVHUZ5BkB3xhmKl9umRlcO01/ho
GsTcOjO4hE9TAfl6Ey/+GDb0KJueLU25H6asQXweW8TH3ovQpkMiBQoeuMo/
owCCuPWCF6Un9x7w2oGx6cQHow0yPwAXqo5OmAU5jiaTADep8JViBRqAZSkn
2s3CNwK92KFRbOCgVPOmjBRKYqMGKYBkS3PVsb32ytUlakVDGpzOhP478cv+
C6ux0BAA279W5Lj3DTiCQ4NoorzNJ353g0qp49pHFMFBw1qXFnd3C4F3AtZr
vO1GhIsepmnZqlaeppiXkLKSA3iAtJI4NSSXFYK+91H5o+QNNMoT6mveyun8
gINw2y9i+MkRm93ONw1uytBGYh77ZMgBuxtiJVVKI/EDogMwF0nonjKOwpXz
J9WHAGNbCgzcwdaEt73xQQUfHKjLDQKzUc622cmDYqdBHJURhpmt5aDjWQe9
s0rBSeyYKOwVOI+mMVSYLZYfL5NBMmsUwJ27ktmvj4gHGy57R0GNlwBrdspS
wGNnSqk2X/3iUeueBf85ba2xOLBgObAp3fHJoFv7dZgZlTuCr67VReO95Kcl
ChAilwNEDYWaAJFjSoHenvth4OuxPHdef+D1iMP5nVkmpR44XCLpB5Zwsg1P
l1B0P4VhDqq+oouemYZNUJiSEM4VFsuSgLWwPuh52u2RDb4/aCO9AUeG1LQn
UAxOPNNTa/UviDI/wxtDGevPG0J6PlOtA0JPxD862VwtnwdMyBuqMNO9axLL
AykczvMVtNzBwECyGYPKh9MN0B8rx83E8djmdiqT3mX1wx6ihjxs/6tVkFJh
02PgxKRqOSUMAC5R/dlub0ITyBCyaa0G3YxTuiQUZ5rcbzii3LIYyGDnmkaD
bjmcAYsTawas8WrshDz+JuymQo9JYHXjGFq60pVBdU7A0vp49XOnVNajPT6I
huJblACLp8tOn6/fMWO0v7Inj3jAI0hieMRNWNyEOZ3o5yfb+fysQCEoOe8w
VGpq3OXxXvLYTYKG4Q/10DfxxE1JxuXwt65bv90dh7jWd0r05Dmrth8JOxbr
BKTZvbD8L0ae7zLTx+71yoRD3Bwyo2v0Jmavo7Yfh3Not7QuJ95nxnfQbti9
YyooEEJlFFYcJ3Ds5+uVrrcjOJ0viK/apWx04ybHVl+rQ8jq+iJNXvKrNgkS
PE6OphSdlEIvXoB6Ov4erdY0RBHZHw6IzgXb94i8pp2QenrmJ3FFeDEI84wy
pJJa1DdwBqxj4BN4m+jmemAXi62ehP1jIlQJu2yyWCMcIFM6FSi4pmUbq7ZM
F3+A2svIE/KcU6rRUgBUs+WAx5uYMTkzbtNqeLA4iXwaUw13+KfDS87VKuir
wI/9kz6y8sRAF5Zf2m8Pl9KiO7hkzJoIjBRN5ucJtH4Mq3jThMmuiBWh7pWu
E60w4ytOlZtEyPgNckD6Jnb7Iwa9ZloaKoBJ32vGVZXz3QRze7Hg+l/xiS1S
4Bb4knitysbi4rfbsf7jQ+5cJAzJY8xgalRucd5SGcpFR72TfXi+NNvBJ+c2
rFYPlPCemIRrM2nOCH9V5TWs6oAqfRnU0ZNpK03bQWdq/l2f02PY+HTD6KGJ
DWw01fIkJmSmPQ7xoySE5ZoDbdL4113lidw2aDEeyMB25GpWaP/5B3PeW7Oo
TZeIDt68PxYbOOFe/V0oK3/aiSznmhPzA/TF/V+kU84WC0kTbMgTlIQ5eXvp
/0HBEkk7FktlKln5aPG2VnFzJy3lUCvL8VHZJEYbCOUFz2Kh03gGfdXv59cp
wcIIYWlqW/Dv5GpVmAkk6xVUwrLFSIBn55EHp29jiv1A9QNLxbxcG/UwbQf7
tuK9mHepASWd

`pragma protect end_protected
