// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vVJfHJvJUWLUgY502d30sCvM+eGLSy/CrV01Cq1PDZb8aw7zA+I0ddRaKGHvuURozegvmW1fTECb
xi4XnGNGpDmfeyo9BGjgVNKjVM1oYv7OIw0nxwRIbc34QjbHWh2zwnqHN13hz4BUEpzN04NYYHyc
UIlxFQAjx+6eNc05wkOTJQtMCi580wTA+9bkLOPGywbxH0MqRtD19L87OO2RLReRXZAVr6lfzyAM
/FVmU41Kk34kEHq37IKsjkx2NgikL0ugT29gIuiiG/h2jKoC17xiH22H0lOkKh79FQmBGQ80axHB
5DnwSgAFiDlJRrjafi6BWEREyH5cOmt8TTY9RQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8768)
tmInEaBNcoECx/QuYOt9ZrxNbLHLYRGZ4ulff6hzkVTnwmuHyl7Tm0O9RVOJFxlvzAxjwrxkQPpD
+HyM56YkcZCsuR0oa1JQ6KpSlRCXE9eVVYMiytS5ZwKd9DqreIxWcQb/hxoUnkaNKCkwyM4H001x
2YFEOGFdh43cXmaon4yoTVG7A4C1W2wCCMHeKxSdrGZQgWsQdtarXqcv2hgNBTGhas80us97Hpeo
vEn3EdzywMDOMEqQMhlm8quQIGf3LDCdCHC6Hqn4kKKjtaA7ahuyTRfly+XG0+4U2Nin0NIypmYD
p2xshY08kZUhAkUghhMtFU9xudUGw6Jzg/rLWhc2m3fzki0sxaDyq7t5RKXTCpqFHzmDGcE027DA
ZNMad9uIfe5FgkGQnQdtwbx4xmFOz36JKqKGVvHQrw31nJ1DRFpaKSf+58/yPPoTnKbcxNebI5Mj
pL4MHpU8Z6oYsr6EUgSHaH+Vu83YdOVNchhaXOdWt76wQDUEifxoWx6dt1//sAtx5eOp/lRD89Sm
ToNphcPEiTt5OVz1vwwiBZFNxRVkHX5f5PD2PO0fWeMTAXl0W2HkgLcKJ1t247xP7E42IhfUlAjk
0kQVX62m4u8MrcfGvZXt4H+69PrD6slGdhzWvmnPg4dgfwHqTgWjIng6oUbhOFwt4K8O3fcifQ6j
vn0+1bl4SST9LbJvv5d8Yi7kJe/WIyItoMdBNA9QmmpVE+NWcTDgncllKZHKiD7FYVQ6ly+2lZFa
+kArvr24SePLZ0O/GqP0wv3A1IKoZ3hCTy/S9Y4rmmQcUGP94vE2juujr75k1tIntWR4NlCtpV1r
qkeJH0zQUABMdq5tD6tzkAK1LDFoy9lfB4IDy3BnSWGXOLx/kk64a4Q3O5UWhO0AcIwcCOWH0Q2J
PIOw5DtzpvESfTCDC0me0T6QzVKBE0L5EE0QqgrU1M5MzszdJzbIelAKUO+D57CDEsj+pgS//Bbj
4V0kKN27TeJSVFzuUMqzf/bETRBhUT3IXhlquj21V7eEoDh1qptUXjpX72e3D9ZPKFbBGh/ZkDSO
q1a7FCoit7tn9rBUYwwFRWGe6So0SVyWV/FQTY3hQLwhYMCxvm45YJU+bM+VtxtGaVgnW4lmhNXN
4Nn6Mt4Z4/iQP1PMz2OAYc28ApJmNhgufE5kLA1yZ8bCr/vgkRYaXO4EEV7UiP4zxoddQeBLpS0X
zrSFNGHwSjJjeBnP5Bocu9NlB0V1PKwWLTSzSMMM2gfD2ObFggDdT+T5nGrNnBXev8voRIhUPSn2
c3MBzFfrnOMTY4wvtT9Pq1Ud15pwPH57lYsp58pJRYM6SNJfvQOY4TAT/8BqPcBdmZKjPEFGamnU
FK2LMoev++Et0ZUX8wDeG8MZagPUki8O8fALsRDyoqdxCxaRBafzeNUcRRSB76g0RSLtWSc1SpHy
JSx87Pp+rQAA5KqFbnUpjm7Xhz3N/z/1sG8eMMZkEByFDjMm8nykd93IZUGPyO/UCoKpFJmNnLBk
F9ppF1sycKXntj6MuFWRC13lj/U0AVPKeJakFrbGO/m1/h2IbX8qYa5EvafZ3E8O0821wq9wdUw/
azmE12vTlmNj47TeZxRpoFnL4saz7+F2Bkzd+O2I6QOWJ9c7uohQy7ughemQy3ArWVYYRP7/eqr/
wwo5ZCF2uRNVSQ2Au/MdXPoWl19ByOIWluF7s/sLD+AuU9HHGCNehZ0NiRpvXcgnCfv/CEPa7i4k
94Of5YTjnz4utDoEqqeToufbcNEam3/lzYGY7N0JN42b7Lamu/ifQvoZ7WZLN5fWYpNe95QxHhMt
fqW8i9GTYA89ii0ffc87UuhZJmGy/OM8OfhuF0r+qWt+Q0opIPbKi1CeKFLaBMVtUWctiDxfM1yr
HTOoooR7Q1tHIga1PAFT0jL8uZ3ZP7ukGzXOu/oNQI58x2GmexPqHnGAQaaBJIMcL13dmdelUg8z
A5cPdjwXgF1fUjXSyC7MQIKX4J6x+PW7I056M66/B1vlwfUiuDNSA6VfGBNoJQeu0nYLXtaj7/P3
F01I4x9LGGnr4FLu3SfKc6GHhSea9JGPqxYG/2/fowmi+l9uoNg7PIW6NayTMMYrU8jp2zZmEEqe
n4EpczdI0NcrKgfS88uBbswfHZ983t66KQ9y0MIGt5kxrbmrYEZVSygPDv8Gk9yHvszGcFfwSTBF
PNChcZXpk63/gJHwAkU4qpu6TIgcpAahIptjwKb/2YdI0IlWlEb+tXAMT19BzCUzFlC2nIkXGcXM
H6jgE6oRErrE//IXhFqsnvLRxDK2S95bU4o8lRrlp+JmvZOjfZS9wmRfgFWirmmOZrCd22XxDPX8
WvzOzj4FAMDcqIIaPto0NAtJOhoFIFM488wZca4CUcocATk2RflS3yYSH9aoGc0meGxaJrqPm3to
LY9tHLl3d1hR0Luodj+qi2s4k6tjNb6P9dVI3ophLhHmzRysc42NuAgMI/u4+cAPUpDeVL8Msmy0
RHYc7sLixDPCLqt+Hn5NdhFaM4kaMPqRj8QPNcONicFtXk/Qmtr0Dzn/Xrr93d+AoSl5uJoD9ZLO
qtIT4jYcUh6D0SPuNjaNh/RMSTiNEtpWSwAe70zytiPPpdswmgwlanAqyL4M7Eh7lFLmmgkGGCGW
CKD17jn+qZuqof8REMtJyIefiCNA5KpdvsMwzdxNf/Dm3hnLqxE/P5nllYGQV0yNUAbSdZOj4K48
8FQW9FP89ZAcYwc8OHYSC2PnnB7oi9tAVFLub1alC7FLTHxknrHZs1y9XASVv9zZGclsVwg+VUzE
NTQsQ2yuF7MlW+NPb5GV89c37QKJNwYkzTL0jrSmHp+x2hk7HgKallBR78dBl7nMiV6LvisAB4LH
PGnCBLS/NEViFOyD8WlPBKsoLPX0ADQl0Aw6L8gtVe1axkZJZuit++P0qJsZ43mNyfdaBYTBlVde
Yke+jF2iiAaAubwDDA/4114P3nkxYBLylmVkgk1MVU3ChxNddYj3AoPlYkOE0BRjGINlB1MfyUKX
1C+p2/BQXN6cm56GCvs40JspCGCdeYTfUNlXuzGCoNYpNL401uieRrHxvvpB10NEjQ+7D1jZTaH0
tbXmd/XKV3lChjcYsZTq/eHNqdKPzd2y6fYY1XRR+VkFOCn6C9r07CvAWuhGPH3ZHqrcKiHXsGQ9
XYambeCbeg2UB18fkyE8XBk5WsRDyYfJisQuVl0V3Ai0NUEecYP1HVjW5/KWWSD2MRaLHTYdNVVk
YffQhvuVaeqf6snqHTjd9EoutCzJq5QrKKG54E419JCClSSr9g/8A15K8ZdkM9Gie87hSy4y3G39
WhjjYgJNNT9Bae/RUWMZJi87DRhZoZxfutWlQVDcIiA+RtJWdd8ojWkKwB+C/fRyO2KMgPtVXRRR
4U25Q7OJ3k0ogh0YBDUS/p+KKb5oRo7duu5DokCASPo66e0EBaOAE01ry+QaTppXIj2danTJ062Q
j3KRAaG/Qp5WzaGlp20e5iqXXp18V5hikbsuewG//VlfH5xYJBTE23XbSFDtG21XO8hpx30LuvKl
5ktuFw/eXuUP1b4i2pB1HRB900/T2uyH3+GJN10Z9/iYiKN7Us+b7XSK2rTlUB6BH0s9vdDIYuo3
8vPpQWcDzC0Bva2zKCB5b2noTYyCUD/e4PJKri96hZY2YJoaO8A2gxzKxBg18pImS22qgXYPH0FE
o/LhNHlgg+NetvueseWCRhN+8gUOEptBdq08wlkE8bk9de0Iv4J5StvJ44lqFPlxaJk2GS7/bBi0
x7hrR/HAJSj1vlYxp1vHV4iaEn4DPOfxxZFtrOj/7zEs/1fkvf/GSxhy1W3JBNNgU/a/m2ALHK2Y
sULQbhyeyouFNjD8c1llSiXiAOBihEg7+6xDXqeNFa0SIgCj1ByUdtESEQiRa2TrONmiAzeMU2IF
Ks+WTzDgn3cNO6fi27Acvu+jPE0bV3WHi9Cytt91DwfPhXs0Vn87ZiaFhLE9rJ47oK/NkQ7+xWcq
hvD5vaijeer9A+kuTqEy42S1c+bHK3LFSN5yP9xLf7pG6fIMVzhErOdyONK2sanC8S94uy06ee92
Ls7x38sATuoMKW/4Kk+oG6CiL1m830Geyvj0YetxD8IF/tHGiryMzTX16aYNV+plXrYV1jIuPH+r
2qJOTq/yRKp6e9MdYWcytJeAUOSx7hA161kb8P3XqFddrWCFYT/bhCLcQO6mX5XWjgCcIBT7vfrW
KluYb6UGwI6pmL9VLrrRULejxt7fyS82TDs6cbLq2+CdvvRPAsEz1p/ZX+lEK2LPTMWWDNiMyNCI
APINqYWYbD2ykD7nbyJPoVOebw2o1W0eEO+qHg3chzmXQpFnYOZKfdVs6JPlDRG5pccrk7Kgpg7D
2okEoYABcJRavwdpB9tH+7EsuUwjuL3i3aG+21R+ngdavktxmG6qdD9q2qxTgWkSUqB40tCZnIN6
HeCu5Bg+4WO0bHOTVPaX6UZDP+z7js5dYZh+Rf0bby/E872Y4XvkKLAAEB+h+PkP1mHDRU/OmDEA
vt9WTPVyTiaxyfPLch+q669iM2/+k8gzlOs1arENftLUqSF5Y6BpbsOj+SQ2b2oUopPofHnveBwn
wVyAJK8RcRLBR1+jFgdEEkBQbKoWcBoYYH7F0y7msL344PmP2r8mWRyWGaQKyHSSnCu2Wm226np3
K2YY1C/R/U+LI1Y+VpYcCnAdGn+hm8xwEaQUHlp6CvlsvU7ymWixEjOkMXBz29IUcVKHYg/ta5CG
ZGuqj0oo0r6w0iFEIAbJR9McwH1YPyQ6FvvV8COM6B4NbteLQL+VxLLDlFqXx93bgN65MSTchNF6
b72Mdv+Zr7Bll8JBpIbCwwUT/nyl9p0LAFnFwhgasAm8HzxJVFmMlYDJaolRXm7Lrl3Zw+1tvl69
jxaQivprRIvQkD5G6mgTn/QHbqE2/4Y3RHYbtCkvlovWihgqw8Nz6/5F0DVgT2GC77ScFFgHvsKL
MmhL1m3vrnY7PRqK1yvcoUCC2MICZraIK16pa3PxGSkPfeWd7wKmA77t/slTEFb8prHbjCAKWC/b
e1ILNSGREke8Ajx+brlRJRCskaRYMup16gC8xlLNyzZvaj7BJP2BfEx1t+ZXhY0N7/koiuwra3AR
atsrOxHpf86v/rLUboeiXZUf7SMb0rBV15TJvFn7fdgubEEZbb5a6kZZ4t3qwBsn7/Kx6UEdDuDg
tl7QKAJS236oukTIXTO0MuqzvUhCf8Y0eVUh+tCA9HIfnN6EGkWRRSd6MOKZKh5CIvUYlobHCYc4
OIckgv9RWUB7rKnSn7AWv+9CriYwTK3Ev+3qY4L2PGkC0B3ALFf5OO+EYcRfPGtL/V0Cq6zybSXn
gojbEJdmMu0+l7JEcJ51wvsMq3cUy/QKsYYeOzZonn/NhEiByepCn1Ow8IQAKh1nEbyRisZU1GT7
vpqQ1cGMNVGSFOH+T0np5aEfQiy+ysEL7Ux86Qabqy5XUg6Uvkvkoa5Gsi0FUzHCUSF3jkEslsx0
cVMR4x7ecTV0mrGUKE1sJUsAtLWWmU4KRrKoKpvZQdbYzW7LhrNXVnqVeGuwHUXUcvhUoRoW2frQ
Rk0k0ON2j8317QaIJ10k3KVM3ughFf61Urhi9Zd+kJK0Zit+mIoGu9UbBQXFLRaMXkAIepRrXwOf
MjGfZlURdjfePxEqkLkGvG2BYFH64rW5bOZkkYHSIwmE9fYhdZjWQDQySYMYJRpcjbYw3J8NF16m
45c/y36zDfaeAXrqdUC48tdw0KC55MqPHObhphaEF0PP+AyS5u/IDVld180inPncWdlREUSbeqFj
ijoZKyYWt6lsgvl8VDVT51hYNOq+Jg43Cxzz4J/8SxaAF7rImol0KyStd3RTrP9r/6tV04O+CR6O
P0tS6L+vjC3kzIOz/qkGskDtKqBZObRY8mxlOn3Q8SzgqTIwosdcfBy8r2hQTq7noyPjCTSzxjwW
tZfC+3+rKG9y1KJXyBgYhTljy76b9scySdhhYIA5HdLYJhEWlvD7zHrCNLmvfDnE6WOqvlCWBmj2
isK1dFPtLI65E+oukFbMbdctzntxFdKJ3kaKnyTOYhpUunF+di9nZiPuWdw14jGme3bXVpvNvhcL
LUbgldczBcnBbIsDhEBYZSmIYitOxr3LxlIy6ydwN20hwtz9WSD1vur90QOFBppBocWCJCww7R1U
HxqjOQN1g3Rs/Su41RRQshT9h6vWbvI7jc8OrQnII9DqRsUlaGkaTXqwbIeM/ASnSt78ohwle9jt
xjlkdBMGdjsoIUZOdinUQxeVqZnUhqLyZhUoSADGhI0KrRnBifJxPnKz3SRldmSYlLYHszZ99Bc9
In/wEpcJ9KLEKGjwARKi2CVlf/5Al0PDaX0DNLAScwr+ApfWxMbPl9xtO5xScQDImojol9NuIeiP
NU1nevAruOF4asHv72p8qm7Fj70K7IuvhgYHNhgG0LLzcD40XDorZTqGyi+nSepQdYBVLtGdtSa7
KeoYNqoQQmBPedBRx08vOKj2aHBHG71/pbu/9MdAZE3bjFEfDalHQ2jpXLjZM4HCW7qHp7j/b+js
RtoD+Zuu2fhjEMemC3scZZ65OIUt0Oyo6lsuTektJjmnd+p61cgpi/MwQ/oXBUdJB29r3wVRm9if
DCRgob60fa+b9sbZCLS1Js6BK3691lthrtYj9YsIf6pj2tMfhL7NHy/C2SrAHD91u5wwEPE5rZ3q
O/1S+vcAB9gNeahPstKvbdwP3aqiQUDnilp9wUxp6FTsjId8Hh9jO41TDBx2RSyAadLp+22jpm/q
vq4xrp2vZk5Lcs72Rk2wbCIGQB+IqPSD0YQDUFITuCIMMBx9GRgxDDuBxA6CgAOuc3wRdjgFCboT
NnpA0YE21zLoN1yS88n1zvm3aHFHSysolNXoLPcspIyP5IiSMQd9dWF9qQP/YyeNbULxfJlmrVVn
aaRYKzz2b42s/zSTzKHxZIL/NZcSp0iyXou70rqA/eu6lUF7B7vdjOpbJQwiY4/ROUbwLKbFh0l6
MOJZxKJ0DFfVyLztKeqUb5gdwUqPqoAXBhIC0zdLk+COdFvZHx9S1O0vc0rYqBlXqgedJo90sGg0
1QjvQLqEczthKIIYPrIkj0McMqRkFVkSFkuVUsFC5M9KA6LfgMGHFRf8EfAwk03ZMDqSZHYyZT83
LRmHZJxEMRYrv3ZHxqcEiNTiw+BHTp8lX5CofW/oLfV1qtgzZcf08wpQveeqbrRpGnUBL+IE2K2w
o96BvY9JKeDlWG8V61Eq1uX7djNnQhrHupLoC06xAneDzPDukzz4Vq4UXeavlINIhgicy+gUUfys
IidYiiBVm/5zlGRmA6M1JNAeKOZU/DFanvzIFa4Fi3NldMcqh6PEhxI5bRtFBnGPRp4t2JBX3EPS
tunfFNV8u8CM9P+8dkL7+3/7BU3VmdOQj3+K5oy3aTldm3NuWHuIJ3fyfvSBEkwkbp4SuTUfTgIL
pF5MNsEEQGmeQ4hRb+NbzrTU5mtzm6WW+tuTuObmzg8CbmjByt8EBpN59z2mlaCgNqwcEhBUXfUU
sYeE5A2iOOV3FeoAxIVhYqiWM4ALvKgsfJNyUJEDfzYvmA3E++HzDmkrQfd6gLc0i0W8HeUyM1az
FhBtCcETE1/O2bAJ9Wc5cTLljiVnLxRGN6sI6W2bOe2Jxj1MFDjOCMqNAp6pdzSXhVuoxy2UMhyi
AZcFwZAboqT2hrTA90Uj2vkOpfkhMszvMyWPs6fpZtNHBTIgp9I03MaNiX6Bmikg0laOudaH4qSE
CTJfsAFG3F+fo1oL1YNQQgxSpo/Y8Gi3cllwXfEq2gHZLsNdEdQgLy1ejDyI4TgmysgswFKdXH8T
nBXoPn4VsQwo7u3Q2f/EbW9jGK0TTbm6Lgo3FjC1ahuFyNMvscbgGdR3fmQ3o7TxK+7vG4mSD0o5
aZkQ9a+Fy64ac6D60GtxxQJGwVudjVbwwT41QpJSw+49JZrCfDEY2EcCNC43bphBSVDwNkRldmT3
0NsuvUdUODpnER3D/9MgyKRyn7iOaWgh+/JkizYv4AmEQciy3ie47l4dYSNrCEkmy/AUZ1WcZ26e
rMZlqxEw0jZpxLPHc/QwGimayNMWlbawDKVFJ6jOhHVRakUYuEIKF5N/euLAluuEcTN9BhNucSeW
fIzwDBUT8j/o8TSEiLq9z1Oj8qDB9zFXUPPNMQ4CNaFbjwcyoTTPJOv/OcSLYl4liMGY7pAC7Wyt
Ejm7Sm12GLrYraDJHBCLHgbrpvXlOh5tOO+jkbgr01BsOBTwFLG4wGtTslN5GtaJWMGoPKCZeU07
Ke/iasMgCwhp18swibTgkLWS02WLJtp9XfHR2yHIC6IzZehzr+cdzzmus+eWU7mAKvemDALbaBWp
JkqMS89QfGTALkBur2zSZsxlyiS8dpcnRs8TSIybCsega81TewGImpaz6TrETzOT0W9x1tRnNTtG
WoZHdh6D2Z3if05O7T31/78BGXMwHSxXEy5B35X/kQyIUs7eqHDpncoGmCXSje2KHyjNNhKr+KJn
ZwAiy/vxDH1/AOAHGkYpMokwJkdIcoe1ZTXDnRwkbXLVqmL33v28NTnW6+jqo0MEFZc9W9OQXS/9
Pn7psYCcetBp6u7jyA+oe+iOU3PYRvQYgU5GI1iou/Qkm5ZPLvO4h8Hl05ADKoJZyGldiYQgnkaM
boxDKPn1taaRknkt9TmMzB3yz8eiOovLAFVWEbgon5u6AOhvMRXHHGZhwBZ45DP0aCURvmDPoeCH
bXjm7Ta+NPJ9F2B9/o302ZDOfGJijhGJ4taUc0NFfvJsk00GHeY0V0Eq6s66lFNzKpxDoFU3w6Ty
ZRFoHgYniBYAquxFyQCZc3oQ4BgzrdpwiDMi9oqxRNpQzKUUbiXhjKD/119sK/kCT6+MkiauW87H
3QKtb4vCQpgBPkE0cvTpbRJKwbzlA7CsHv9Ng31gz/ONPuLOBD38RoB8RkzOdpTfDncgVxjJhLiy
SkGSlfv9wZokM6+ciV/cgbiqwmuXxDg52cJNmPMjiUwitpOWidm8EFpX/jiaGTm/S+xfARzNLpLV
St4m6fPd6ijkQK8K9uuwDLNisbGQRLNTkttheZ8OZ1X4tEHH5G10aVNB7fAv2r+dUUUYUOiaAqjk
/Cu250qawnF/o7NnQGliru+qvYGGpsUXaz1L58tNFUP/Feny4zmZvQQQp90cGQtlNtGSmo0T7LZq
fqlSi8Sh1bTjYFZj2Zz9n4rNZ4lthspUTwjBfnUoz57WoeJuamnQK2nW9B/DSfm1d/rDfgNDAMW3
tOL5bIDNmihlTH4YFO4y42htGeXGHpQNof0G5s3rCIcz0IXOaGFdZiKFnAaOq56fbmEilb5ARfDk
zOOBjJ7f3cSdvcIm9I/vS27tI2tCn2+PJKb0NtmssPtxTWYJef7IdsAd68cQkqdAXmDSIwoDb0tE
Pytk54G9lZ0WxiRlvLn1BK0hV1BrHYEsuxoBsbQezwkI5U606bp41cbjic/9WKdAT3C5t4wraMbP
O9TKs2HMBm6xy4J1tsy5PntT0YqE0wuD1wU3PwHLzL0laLDYKgJqUWPDIoCO4EFF+re0jIpV813C
WwGqUd5PM0yA9CNJMpsfD48HA6hNb7fRZtCJ3qZrXtVrooNu4RMHkgL65aZKt4Y/4dJ92MK0u8f+
MEyVkPS3uQWxDzRlxk+Qoten4+5l/+yUggzYKUfn9tRSqfhlXzUEyjpc0kUkpeop5m6CDsnMnOxM
vAtIId70QwU0ayn1Xcj7tg9w2XF9aBTg7FmNpll/vpj+cyP6vXRONVCaBhS48gsjGCALOi2l7EfE
mz5YAJCzxr5SvKpBiB1ICqpHWDAYOXJrm0O9eqvaJWVzNC8WkP/MUq5PiZX4KmxiUU89xuWushrI
W+BJiHemm4oImJVCbgMixjgkaVmLwuIXNZ7t3oqcoSNuXiWEjqVCGMooV9r/PRpEet5/A8ZCZNZe
O1e8n5nZasKTe4YXR9hYRWOHZGa2uvxRI0UQC6Iz+aMg81S8187ncjmW7BszkPUUg4x52+OkafZE
Q7xrLRVMIOwrQyIn8nF+SmCBe6Jr0Psn2mwWqcs4WgotM/gS7jINs/a6BPssoTu6QNrtZiEPcDCY
Rpsns7elHieM0oJO60eNYfwIAwCO58QLD9NQdZkSFkQMxcNKVKR525b4OD15wwqQIEZhidITuKep
KenlpCfczKf9aez8wDn2PgfSfeXXBeWTWCtPyBosQrkXgvY0LSzd5bYtfqgTYA34R6dZVzmlYjD/
lGN5bTcq83Tt6jQGTCZPlXowdJ+NOPKrbp+QbjaqJSDAhGXGsktnIm+XLSKMg6bil50/Ob8OM979
E1CtUG/OJJiIMB4Cu1FqGGY956zC8uhjcOiJURpkCIUMIWe/6FzSbkeMI8MbzWZtILaB6D367V75
uJJSiIFZIJqaHNFToon0XMnxrdf2UzK0SM1GMby4PMbYDynVJP+BIS8xA7PI0jKgROl/dYgE2lof
PbY27zrEU0BaEhfvqlLTZ2rL73mS+JupFFxppqX/CsYDnMFjD9DNrLasDk+fElF505xzxtL75u3g
CrYIFZP8Bpf7n/QKh9njtVUBXQXGrJdvQ3HJm+Q3LtOzjdup1P8V4t8wPVSzyP8skzNJ7lkS2bqF
esyIyg1SoagRKDlURlpX0mb2J50yZMXKHNAFDUIaz1ChO/KVt5DLDjTdu3iRWszgkyoTDbxAdvTs
jLRI5mabc25EjoCUceXFkKZNJmI5d8w12NCV5puut3+tzOEbcL9oBjOXIj5xzaYqB3GFTndhU7DF
EPL7HOUkL82AWztoJqZOzpaXTEGbqLrVhRWB4iTQYjkoS2Y+DdjUwLUiCwQ5hwtf2sXwLTf+IdcB
eju3E5xtcg2OfBRuAnNUtGUc8jE2NAtLxyNT2j5Ymxg2dsduQ7b4bTdfOogNx+2NGomzvv7acsgl
cG9Ngyywqo5uYuf4TuAA9ZecaVJ2fWHGCh1Rw6TTet6vT7x1S6HWwSwjqEaNStGy5JcXnlAvTQOV
e0EXfjTd37VQB6fvFOGCruqx85S1FjsDOCSgOTMoOdcLagP+QIErcYNWPGzeCegTe2Ba2yOasY7P
YEy/tkK1jev8W4p5lvXeyVnaHrCZvv5m9xckhFwY71m45ZCIwXwG02Y9+axnWp59f/IyEByRgITt
+2UnVl/VSR7EOy72FO/DOY1HZzEI+uT84LXvkW3lBjYfUlRGkr+OBM7Yh6tmVCBKgZsnYUVi4tGv
Y1MV5Ze5EG5OhsoZVKuzRCOD6DTPyR8SFV+7B27xJ93RPI40YkNMmlXKSDjLPHOWEKTRzA8z2dnZ
rX7tvBA7DElHdcKAnMqcXO1PWLMgmOhwW2I9VTSKInU4iLio/n23sIC+WMdYGeeHfahVP3zO346o
FzLo5ghyVJG8SwF2XAfaJ28NgdAOyzBAsEEV5AT2QXNtKBdfd0YNTaZc3Bd6+yV1hw8x2umwwxNg
KGb6VTPYti0MfvDof4Iy+JV/lJzcLYKdKSe7BMJVjLc/2QE56XlcY+qbz1Ijb9bJHT5ABWhepdcL
Dx0xhMt/xuwTp04yHkKpXNlASTFeyCRFA+FXtj2Ew+AgEyJIprgKCazXH1oydG4=
`pragma protect end_protected
