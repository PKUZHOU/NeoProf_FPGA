// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Rc9IaFJJ79Scv27EgP4Jsoe6BKoYMP4N3nkVtgS55ExZCxoRCjwFnLZRKdnYwBCS
D7wI0rl41b63H2cEx78qObIf2HmeggkwD/rQEjn8wGBiCxqPjkhWmhV0U7q1Ol/6
Hi3sVPD2mGsoJoFfM0TnORJOhZRhDArzf3+ItWjmz+s=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2432 )
`pragma protect data_block
B2ZxaTK/DeqaalIWHrXXd3zEbxI72C23fdf2ffHzU19v/Le8KNSuzRJUuS10a6yx
QLi6LO2AhPfY56WRCMLAzFQTKb9dopOAJttuXZtXFuNptyukeq6lEdMU9wYNCJee
qjYwjMQM9piL1CDExj2gj7p8T7TeW/0o5l3ak1iG8LsEhPLVclvC373xE9mHxZhP
wFeKam9WUCTxvHtLfHJCN+3K6Ff9pYfc2TzhfFOAHxgbdf2GBz7YnWMYe8Pf1xPG
xAzfk74mUoDvPVEO2LoS6G4aaSlhzSK+Ntj24fCCtSJArSyZnkvnS4ezm53RKIYB
6qTwT5IgImF1HTQ0MLQre1AieL71Rx+zTM7tASyF56NA9pDsrTBdDQkZnejvky9T
wE36Lf99tz2Lkg8ivRImKBb95k0KF1qqJzJ3jIP1YksvL1E4kQf7gQSMvybai/30
/d8+7hbwSG3z5Gwndgc/R1UaUdcp9h5NSQ0DOnPvYk2P5MeiI1j4+rvW9YXymwfY
ndRiostrf4m31IalK5qTT+L5wzT2ed7iWbPeZzciC7FA6Vdfx8pIfoz4nN3ruDF5
aMWPtcsXkRc3B59pEKPY72Kre3whny3YcL9GH6XQOafDbAjhryuUOr9IFDPt0iBk
0AeT+jQ49PKFQo5wgQ3io51ATuVlYnF1Retm4WralZ7iaB7/+j7gtQXeeoLfZZS9
I/gnmjinM7jcPGB7yxroKcQ6R4A7Ws4Y/ZFHzbj7ziEWQCuk9Dn1crdHtCzTAnOD
681GQCUSh9uWJ+EJfh+4ZopNXDcxpzK+NBoG4pi3RGWHMjT6O3hwN1NMIKMQm8TE
2XOHWmE0erADXisRCmUEho1nJe0nuC9RP4CXmfUImWk12jLZjmgiL0e4uNzKLlZt
BpfH2ulU/iE32MZlvaYK9mIcS3gQSF08RFTCWpbm+eV64K9BnbGfTgg3JJiUbeJg
USf4UMw2ItL6HAdofpEk4673wIlAx7X9WKJo6zT5t3M9a4cOdWzgnruLIeOFz/ok
q3SaMn+qDsTOVwrUGhMMU5aGYlGNdy02rixh/dT5Po+sg2tCsxFk6452iSQsxCOG
lc3FMx7rypx30B1KXjqgsr1spnBNXGCiIhnAIjIWgVAmilY9ffO5OAQfmB/suISr
K8lLNBuX/dqaJX5di18JPePV2EgC0ps+cvh/qoOlibgL6YyaiWoeM1uquO8D1EPo
vpTiC8pw20oAPIc7nSK8NIXRhJdLfdYOeGkDj8vIYzwL2gE77Cr7xMLju7ig86ph
JAGo//zvQWi5gM2MhvOgmBbLaAlLtLLU+mgKRrXplp62SUfertJkiQMHV8Z3rYOA
cVyJiHcTWJnyVvFUUInmm/ApR79ZowsMiaDJm84lAKlUUjftpGMpZRz4pm8Ya4NG
RpGeB2V2n0vnSnR+LADi5+cwD54LdlZubUQ8hsVCt1HNdto9K6PEtgcUdDCDDP41
wNgZhQJ2EH9FTduBVoN58Xe2PMh99YKuWolGR9SRlu7m/YXul8fPlrpP8QY3VEJ2
MiEYqxaA6wfnXuhQRu/DnsvCAVrHw4yw0DthnnWgR6nSsNKFRWUN40Ph3JlvElAU
91EHKzVJyyxwaVMwBIdJ0cQ73TNjgkGrK99darjVqt2ADmsjlaTZdYXkeqm5aQRe
h/JOXQqGIbVBXpD6eFmeIq3yY540NlQCcvkNK2keA94npYUY0bFwnonL+jB5FMiS
0yua1nit13cckVdBFu7tR7HVZLhlQVt25+g+YecOa7M/AwecVp1J57egAc1fKyYg
KM+42KWhC9xgXPcKg56phcruTlh9yPudX245BLrB2vPk70q96pv5Uu+j7mdYn5SM
CozW6XATJExa1tYiK2ZL3cYZnlwMfw2+N6FExa69R6d3OD3CM3b0xaBK0GHGTX4/
up53rKYCE+qBPVXnLJz7C7KWVBaK/fU0BoQ8jzPgp2noMhhUbT8SROpbzW0woQwc
OpSq2S98kpX0/eLPxrwM0OZoWNU/rzu0Twdl8UmoePleGQL4WW+eErjFIRfWaSqZ
U6H1HANOgYIC3Vtr9KZSZJ2iRdaKprJcBZzadf2BLXeeddIAOCyLMjDixuQBhEhc
1OFa2Kq8r6IeOaNAmudV78ZMbBeqHMTf4j1Dj/NchqQQzC8eYW6WnU9CB9sNEd/1
YuqBp90LlJHOUkMFMyQDcS/xLHcqz7RMNGgpQuG5P1ErnPigFoJtqErtLopXHh50
gmSJoS7SEk+6l7KVJYfVW0hxCPlgNWHhoRgeLYsseMtOC1qZfRG6HGe+wQPTsxta
m5IRQjW2XW64Av47Cwcen3vzAjhuy0cu2YTB4/uY3x0tis7Dcrb8S5CpP3b3hvMH
WP8c2UNM7qERYzzLe3iEZoonju4GcOMLhpuLVaZDPfVWbeb9MfYZQPZ+dEv3GEDD
LwlzifJbU4vfVghjBjeVBUM6MNvOceEE9Rw8g4Jy6K7GgA2hkXec+ZKluDlOB8wP
OG2mAR4fCzSpJC3CbhEQX3iS32S01xZ0WFp7u+moD4O7yUQaNwKzvyhkbSEtCCqM
HbP4OfWlhPHMitOOalGI3A+0pKj8I3Hg9DHeyAgTdQ0fdeAk0kXnpK2uC5047wt+
ORC8S4cDTl3aLvoISD0ZMZoJbs3DPBvX7yVlnU/X147IR84e8+zSSgiBOpfuJJm2
Q+ZH+kPXyY8MJmMbT1UeDtc4VWE/CI1E2WYnzQ28tB1vjJbwacO7q9bWrUsOT4aH
1amJsC7GO93wA+/CvhHG0wuvDbP6eMPUS4EDc9wNT9cI/2yMIgcac1iTRpv9p7aE
pjgtJv2f/9aaT0hUe2eybHhYhTUP18O0fN7NUZJHrZkRA5Q/Xps5AcI40D8ck2gI
m1wj8lAJLuwAkfQojOFya4XqinByR0VVI1aMSB5n684O7FefPu9QUz6idGzLUSum
tb8g2QSbs8kHMDt7zXNMA9xVJPRUAVgU6Pydx1aycsMIgAoDhiHaG/l5/QgJi/ak
qfsnDvC8Ljw+QBp5x0kqyl2ftupEAURr4xqjXfn7MJ3rIHHu0UabX1KC9tce1qy7
KeKovm6M3/v5ablkEqrPNdS/l6A9MtjUcW2lExGaYTjtUkgwQtlgHMUS3+klXs8k
cEBBa7+ovtROiwKvx9uUeJxZ4We7vs8jj5A14/eeP3wXa2iONTJlHOCPIrFVE3QG
FQwadavoLb/oY7jiSkcLf6CeZSDKDHzv7e57G2HMSz0=

`pragma protect end_protected
