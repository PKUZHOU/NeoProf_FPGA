// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
U1ezs4y88k6s0oC1TcdXgzU/gy7ximOrnR/BvHqtCCZwEvXAidZX1g24Zpa1yhZB
Ym7GRRc5G6i6q44tI41Zpz3eeymSf9/+XoSXlyhguDVHQFqLXDpNwKydyqwHy7FE
5sSnqkS6Ntoeufn9LBONBr364EwQZJosxZQ3P+qjxzg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10336 )
`pragma protect data_block
Sas0at7qzdTg/euIqE/Lzbx0eZJ41e+JVWnyuOprScTO2NN3C49oK7XEjdzmslRq
IynPYwfMVFdd1hrTCnTwMecHrOT8VYQwIVQ+0lt1kmz86q5YiSGL/IpjbUxsRkQo
TBV7nOF2CNz+ub/Z9i7qfeDcb7HXDmE/1f53TzB1JmSeIGdDeSSA+Nk0Bwyo991E
dsUJ19OJWDWxj2nYubGFsAtH92OZeDLT3cf/bHzhSTRGrGfv0XlLjNK3AaGTz+Vf
czoZ5i4/DzbxmByJumtCjbkgUkxzbDPj8RCQ5jtEweGTtTk0M9pryeXUn9rDLlh9
jbbdksLafxLuk0dMQCWR3wwzgBd885TtCTcWjjXh9JPybpBKlUEIMkQO7O9//J6X
gw/hh1o5QfWHxDEgzRAtYBqwBdjna+yhdxUK2a6ytBPk17Na4lsHf2YYn8gp9UQ5
Io1yunsNEvgH07N6IzZVRM1nCDynCik0gknmMtoX4a06/GnhrwwqKXojedgqhzfK
gKxmxY70zYNhbR6+9Sg9ju1bGT/ip79U0yIyb/KX40aZ6Y47CM+WnNT2ASqJGYxC
1eGkTZYzqrYeqTIyTBuSfINHitk+ivLcXIUdRnbOJBs0zfxomP+vJu/t5zGziel3
thA/84cFvwF2gBpE1kP2w+9TZox5sS63kOfwEe/HZnbUJ8YXpBFLgr3WU8Ykai5/
bJJqDb6YljGX9MgiaXbuLX+Gj76J2zBEHMkf3zTMAb3Clh40RKxf67ke2yWXWZ8u
gbY4mNlY7vP59udHoMuNY9TVH6qwvv3dpw6UekVq8DgUWQTsEddJYHzSt2JZAFrJ
7QxydLf6OuURard15Z6sygXkqn7SSlr/GnFSRZ78pd01Fb2IGp5WS0hMmFMz2KdR
oA7XTx1Y/1BhnaYQu1NzqLP7Y4Mf2j0Z78O97dmQU837/+26fv/QFUzwUlcRVqHS
4boj1Xj1YrZ6DEEdnSYjQjTWnhmLgc8guABhKhuejms8PeWc0+k7mCngG4+5yVut
cY8dO2Z5/LRpLaU3aw80AfzR2TtoSJ/lZv4cSKPQC1i8Y37qQrHZwW4uSiK1hyLW
yScqhHVk3D6VIjyR7SHlH4ylmb8Yahcch6StKm+bHdgWxEmNS4DrXGa/2TpMOIac
uhO7LGexhzF8k+YnhRHv5/LdUyvWWBBvsjpEMdOUwyLtJ2mS2H2crSH+E2dtr1k/
qWxY2SeQpyoC7hKdTzrZ3uuUO99Q6iGYBepkX7bxxvTa+WKlm9NlzfVLWeIp6vWl
/h2GCVC38Z9xsHN5lB5zB2OL4gneq+q8xq/7D+qezbZRVODqxCLwYiRKdPiy5Q2g
gb9wjD3Dx8bxlecZyuK4a7R0dd0NfslNyoa886nTWNj6W978RJXVKRfNwPZwQA3Y
iYb3rMzztvucYWSH0v7p/yl9O6yZe0xGeb5G6ZPIxUZc8fBoTJ/EdMVfZ1qwMF4/
XZKooX4HFv76v9YjBYe3ZxlLThup/AtvOjxHbhdAjWKcRd24gQLgyJ04MmjVNvQk
T5VZJat3RfcjjAzBFkMVNvcBszG62i865FpTSVvVivp8R1tcNnUR/qXbw3DMuBbM
j15VUWqjjIpPm/lziFlbShXmp8/DPMV/9RxQQYAXdWS2bhC/2U7XIKxAmOtQmqCT
OqgfEY0Y7a65OnqbMyzV8H3FqOA8G7TqXVpxjd2gnrWyzzrYTBcACIUKA+lfJoYb
Kp0bW340rFzTIidJJ9YeMkYr2BJjn1d4X2+Je2kNuExfVN10TRAW1mvHs/S4NmLK
9ryLFpYTqnXLhY4/85dMhOyd2Cl/+8WE+N2eXUf73Sdy2TQvVJoW1//bw8qLHXdz
n72L8C3Ey+U+kt2ZjCspak57yjdOl16Pb3rIscBqFqgyCP5riC8TyAl8PMFVKt0C
i/uRxUiMUQZfY39qjaz4yAcgPLOzlxC+lhYuBQSb7p5vhcsX3O936JjC+HQ/486M
rPSu6ERbrr8XrD45k/SaXjlLFzUD6xV35yjAau3UqPFzhLrTQ01yVQIPzUdkY8d5
eFXS79pXHnhNc3Pd5sPgsqwzoiHnckIzWWWTWOkhZLaKq+5sSzWzS1h05lEq2gL+
Zo1BBfHCZhKZfDjLnxkG7xMyU9UOvGw5c1gfhcB9GiWdhxsvL3gQm8HedyYutxQT
A5fQbOh8JHRUkMnNvRoSOO8ice9HjDVcjqEqPCwGlYKFDOprrpmIYMi6Zbz22nu7
UAigfd7ksrk3YgPIlc+smfntvjQB8HmReysXXuvlImuwP1WaAb0Mxlld+FIpaNZp
gQxHwiCG1ccSgyk7/+J2zu5m79F3cOmWclJXbhxRF4hk1JBxcgTbrEVraQG0oTYN
XJkM6L2cepubgPjp+nE95Z1eUX2ewUcwcDAv3LkpVImkgHM38pOS9vBxzGNsy1k8
2hTBKDsQXYjH1/V3fJfA/dafymCnXJlqTcI3m0PJ6eZ7bMnYPJaBrKhh7Lu6+wD/
5nrESkKLdCvNmEumAl2yGTmD6Y/JMEHGYInVueMmnrWXZuVXRy3TT3HJJm3b/DIN
qLgRGmw3+t2xcgl3KdUY+zuzyUn3DxUapdqfWvp76fO3uWtT3vqtl9EaIvAAtp53
9illt1xmL7+kGsQ0/bDXC6hgjfHaxV1sMyzfA3zvWkKpBUTyaO4g+nrdQWCMLAi8
vR1Hj5+d/cKMuJxN9040jytiEcpSpIFJbcSvs8zjsvFDoSQmL8QxpueV3YEE+z+L
P1qD/JYhhgc1Mq13M3rodjUjVZkOn7UyInLW86shbqgFNOhDvps02KgLhaLGgrX1
GDrmKxlfwTWnPm/4vJYS7/rcmdOmy9zBI927ZE7UoY/+M61Q5lyLh6fBriMW01yN
ozKoqn/+Wq3hJSqkfMbmF6O4URY8TJF4WXFMcm0l+zB7qV63BZBooLTaKmURNV7B
LqOPym2lwlutx55bExDCdi8wLdhlCLb/EnPYxmcr4LCVb7zQIpAvx7b4sjUEGNmQ
+b3JnHlkylRaNjIBKRUP9RuBWqXskKKWxEkuGmVgGRgsHN6fIzw6OTxsh4FkgkJw
by5kCQ0ZjEMmZF0SveiJEra4e7Kb0zlqOB3nSsbNHkPpgElb+rLUabYI4SpPQe9A
cvAsCw/4ZdqEgkXE3eLtLJD3D/iMsLBUZ8tcJw4gZHFKZEVyxuCHlGCv/CzxL2dF
0s6+AzulIxWdedsej/VQ1vFwdsM+4Y4IWgkXLPE8DBcd6qqxGGoSZNU110jMBq26
TTIX3Gf+qdhH5OF64PbI9sFTVbCC++IFTpCjv3k6Gbnc3SJVNeQrVm50kmeIuBMI
MZuLaye6uNkDpXRt7Zj7SpsYy744B+SihVMawzqg2wRQsQ7TwFg845tLUSoXrsvV
aZiUMuIbUF0RimalwtmlicSX2FcmlJRIPXOd0xPb+/wAbK1cBaeiuWLZnslONUM2
pzkeRfiufDTHavGCcNYfSxAILRKBhGZJnlAzTSorqTBRMEiIgfHuarUkMX2c/2JI
hZNhYj0XkVqG1nS4DI8WkpbfYloRevc2wHp8xXUHkpUYvxD3+LmLP2crYddIufLz
bkAZ3Hi/s+Z2sWsCYrQTbR4yFBi/C5rEKE9mtyguAE+rVpv5QMeUS5J+NmI1wyzH
rCJDZ2bcH0CPSaSYsilWPv8rVXNZslvwb3gTJE4SbaGwYd3ugGhlW5ZqtDEkENVj
20NF3Zb7J9JUdTouL17E4uvfH0eM/zAIAOwmDjzmF8W2R05tjsrIIYhjQ5125/R5
/h5nzFxD60wzk9HRzFYUJ8M6GEc7EVdaENpAc1qVzqFZjKmHeUABbI7RMKzF3ZsY
ftIReJyrC36Jr2pnw3MPBTiGYAhwPyPJD+MIKZtG/VfcNF7yWc+TEYPgXFb8DMFp
zfzGE7ytw423/Gju73e5Rjq+KTpGiSjUKYRffHUAFBSWUqL1Qd2G+9gMGmoqsiqg
Fbu9MTgxwDh0n2jkEEeu2CTGqlE6t7Du9fEXMWMUQssGmVrVOIkLv3gUVmrFdgFe
yiEiceVjeXowPJ68lKi5vGNHvJoWdjHqs3Bp+RsNWgBW0cc6Fzs5di3twjYa5D+3
3BVqLtRck0wxVqI7SXJxzqu+4uxqo5pZWKxJqmVHMMy3EOkXdoHC4ptmnyA7Qhix
lbyjNnflOEB/dRRMFG0OruQMmnIvW2WJpk2z7Ff/5dHUC/7zGXHFQa/76moa8bz/
LwzhoJJw8u3ZqniJvXgY5rjGQeZQIQ6Ga6+m7sr4hfP13xhx1jFF9fNJUr6+jCqQ
hSCMh3YVX+TCz97pO00fJhrB/xoE9KqCTN2J+jOBjDPW8ThyKlRiaIb7qmgNKEbw
0gWD1F4EDF2Zj9B7QZ0jv8we5q8ZOMmwUZzTMiNKfsLPx6mXMKzI8vblZQ0eyNTF
NLSAZdlMZA1Zh6eVeU712Qqe/VNSnUZ4bSureYzfgT9fZDJkIrEc8fEyfwOATYiQ
pjb5w3YND1lT4roMCBCnrhcSNMe942KdKdL+MDi0XqSLbJDlCCbqE5qTZBd+UfOE
fbC+tqwqwHgC2Rmh2ez+Sk7UmVc4BRjEO0iBDzGi1nIuM6mmcQzfEMTOfJ31HLFn
LpG9jeKWJfeLRyDG0wI+uugGcQb+FDf6nJ0jBVYFBmds9UYQ2vLdJB/q9DC//Qvp
5tDaVBX5Zn+3JKGs7arsxzzi1w5hA9CyFbrEgs3osXNzcEm6bqkDoYej1Mq/H/Dc
eSrRUcWUqf/LQP069/U6mQjiwsI4sItG5r2oxDOF4KD++jtlLsuzEQ/cGNmJNdKT
HjRHmRqNCluiariCNyGeXKNhtVJcUgBJJJhLYiKLnAWOD/tm0X6ZI4Il0EpzOBKO
HzQvALIzXoWV5ZdZKqzPzMiJgvZuEZEVM5HuPWYMXpEMTXCsXDe3Dr4XOTajAdfL
leMKwERvoPrb4irZG/ac2uFGCOADTtouuy1d9pSgCuKwXqJs8enUseKaSMXoNMhQ
bX7rI+f06QNNUN2nCavgHj5KQKB14cLeLNk1Jva+70Mo2GUWO0Z6yxQKWFExAFN6
7I1c/n0gi6tfJt80QoO58POazvKLjbIRXmMoOQubnvgsWdoXqMBwcNKcv6LfiQEi
huOn0ardhTBJnXEd/yPHbN7R23SMKfcohwl+fYemd69odcurPNeJSZus5VyQFMAq
dT3tj3Lk02xOOK4NyIJf04TgGAHMTiYIqxgvFdHPFa2DnTUrO+qNwzLRZFEiJr04
oQMZFcloZwYKmqw/MIDUv3h74cMTtShvszgTSe7sVkEL0MznHvbJbk1JplZC2bdw
mzkchPvnr3K6s9KK6lfpCZDB37XeR9xWsdQQ1UjUZ1zSacVwdPgGikvE4D6Sdlvf
iAPO1v/Vgiekwl8qxdmfdTcOKSr7nSOYIvbOdxWBIPLuPrA6UwBphapcfy3LK2fi
bB1WrWbF329XQsx/f6V3E8AIlgB472o++NY8UgStPqrfQWvqtEGR6c3mhYaFOEro
X39cWKBNHNWuAFxmnpCauLjNgDoESY/DVT02gl1QEdfPs6xob+F/bRTTcIYdZPUg
HVXUEZYksNsy98zTG0ujEfb2xrXWctxAUH263MYSmF/w+Em4AR8xyVdgSPxuy64T
sMf+tC2uKHXY2Odu8rsiPJQueoGCItG4i1WyYGPwqKphFSmODDT2cyzQAmSy0jBG
8A96j3m0PH1GhYl+/2sJs/E9Ph6bU8mL04aVSrQaIH4Zhd436r/s0APk43KLM8E6
aJtnXJz7pn8nYuqF41/Xtor6WkJJbmN9M8tZVcSVEfiaXjJOjPFrBWnbJiVc2HxO
64zk6BjikqQq1eEfdsoUkJEUe12C5ZeMNKx9Rg4IDtqCVx3/pWnmmeMKttNZLrRv
FcvpELeVz/xuUiVcJ7/s0kJvpwlbAbwpJ1OYTcbLU11cV6OlGUGNv6S+/IZSiZ7Q
+c0FL7+9J+1bj0eLDYZwevoX4GQifFBz3rnoF5tKiru5r03B+8Y/weMTD4zyLvUj
1YpIIRKQnBMwRUZKuT7d1TMb7QWbFMHrnvylgGGUhNGv4CJ5bcpQpTmza95UNYfU
Yk7nx3/dGedKHnsl2SOgq7147xpAXBjaFEivP9qsDKCk0vuuMh7Y4aCtUu8uzhvP
m9YxNoZEfhUnhtihYDeGmFo+F+sQFk6GBx2BykBtLORPNInxdZvHmtaCSeo1EnhA
18+/z5iu1/F0zXsIRH0eIPCEggbF9MczYcm5vsGH6XaHte6ShIv435lMFL76UEZH
WWhe4YxPZUmYIiyQuECyGzE+Nzuxsa6HWCQg3bVUTQowHwPryqVGxITu08HablAI
qxCAAIRmg/z83pS4DwzmA3roUt2NQZi41493dAWFbL9Pazdn+qFatJIKDnsKWZVn
TC56lb3Ir6eevGjE0sXob0OzYdHS5sAlbUib/BxCK8BQ1tGTDemO7Mv1GN0UMmrd
3nA5c1XLkiTcGu6h1ufSiQvYUbSQqiWK4XuupKa/cN3ZXoMLhvujcJYSvYHcJ/EA
97cxEzNfWxPEDyBfQytY80nq48hz45DCpcC0hb05ecdB2Cdl1DHdYaoCs6a1Jw4M
zk54XnuBnEBta9hsaR5o7UQFss5aKH1iCd3+mo7bOVM0IA0YTCiSxTrLCJgR4vPT
tlrYw+G644/yVF5ssiTRZGMNN+L44cwg1rpe0KAQylS3UAa47cA/XIPtLviPOwAi
JyQKYbn0XVAhI2AYHtORloyUWYBNPp4GZbTK/iL6JGvq89ehC6V0zrcaiQAg6GgM
e40WcSDHyed6eSobg4DADczH2AlGVfmvuyEnGADnbZBm90Vlyn+qRSPbhrnqi2oR
sH2wdSaUJk9m0XhwL5b504kjceTHR35hsAye1JJZ6Ns6kYzkIdkGaHrwBPO9SC/7
kxtAivefEIkBra1gN0TwlVDoWynK4fqAUP7h+xsERPaZ/errzzCKtlnTOxIqNVMd
n7Zm6VJBdulTx8VOBQZ2+6GjJhmpZ6fqjBde/Mq8+54X491bTfXZNyeYN6/cxPzT
59Ug66g8lB/Rh3aumfRmvwdNUIRSnB0STsl4ZDjzOtbbp1Adz38PLJNJ42LXVa6e
eFqRJjNHAE0W6yy3E4+Ym/6UZyQqhxivtbinyfpt1YQ88sed9U76BEqtMkchvvVV
IX63b9mH2SWK2HntEieQRdGF1AMMNM3U/dOYwMU/KhzKgeA6Yyd6xxJoDjn8QkGP
WXEFacqtv8hW44r18SyrZdhN5Vh2UeSdxcX1gQazrvW+niYdOTHufm3qvikeuQU5
4xeVGYtx4GDxJwOd39I0De1XsBCj9ZtEIKPKQwFvgOBXk+c0TiRBC8YQ9uq3ZDu5
nDN7/ekIYVHCQyNcvVFue0UwP6KBEsOiV0YNVqt2hgIeaIxGIa0bAG7Nu/CSoh/X
R4ZN5JK9IDPKBUOJe1WvNMVVz1q+VexaHbbQeM0KPT1idMk35iQVDdXqCGhC8SjK
N2YWY6TLfzHqzr966j6PeJgzuyyWdfvF9Ll2gj7hWkzD72LJyrQ3q09EXESpKiGh
Sc6YbwtMoqfJqd1sKQ1UhydjpUcqrWnHCuYaQo9oFMrZsdeJ4DQtXccO231EvUOj
8qQnk3OdtQOozR0FmPdEbwdbr1hmK+5TDYuxWX8halLuyqMTOTxOa/GJrlbB+n9c
6btLyCQ7V+3Zl6+0l+lDXYoLckDmWEJcm8fBOIMA4pd3EVWfXztv1BzCG0Qnzb86
A3DozKIDeE2XgpasPBKCEGO4dZD27R0du3Y0hp5wlbjTfLRnuolEYv1plj38EN6T
E5Ii/afj0xh6UCmkv9tlPUATaU+nfrI6TGfmNsCfBCrVs7PlNMwoaWMhYoc2hohe
ppUO5gHv0yc0kSbge1UAT0S53oMDAXf7FEOCwjbRr285lZ610fm0mDPO+NmBiNEI
ZZ1zYLT1xbJBNLIXb7bbWz6WMfE6SUBIwvopwP2ZE4WVy2/EPpS7K0mPSwIYouIW
cptExxLEarYgUIosxnhwMIKVK5iGxL2EyReiFUJ+Tva422PG4H5NCnH2x8RvOTXR
AdDNyKvIsgqdyj/OU6w6a3vqLiPiG+5Q8xxEfEOz51A4XofZhptq43nnrkB/q0Fz
8o4q0IuS/o9By1aftWWBvZ6ylGRVYzUBwt0piTqnsTZ/hWrzzawxTD3cLnAjxKRO
tHN5+K3NsFHPIUOW/qcz9tvYWXAfTjVBvmoFQ0NJfiOGb3zSWMDZBCvY2GBBHf/a
WbRnCSguKjwI/TbeZIg6FZ5rh1jm0khsKVjM2vmNOanzGqOa/CtYCdhsIip7xV5D
p906XKziridjSiDmMIKsEy+YwPoYP4F85e3OeJ/nI/hri3sLYCZ7SzNpzuiq8shH
xbbx/p+vFm9EVtyQI4QGjmRzS4zmRL5ZAGiiwYCxoXhTjk2WkPU/zvv8S+os5w9S
wXhOhMU83jPGBfGWxGEuEALXW7WNKNV0fsIIzcQ/sq9va/Vox3wOL1iXUsjIJ6PQ
1qRrlb1DTf7a92KNSOYCCs5n4DBE09pOiAkvzHWO+onoh4yhVsbS364B5kGvTMx+
Inj4K9zDn8mMSz0COzn+xVyMIxGk1KirmRF4EQ5GwAX8SEBCC+xz+6a+5uXj5hEZ
khLHXP9s0isk4aaCXF4xKu5wlbq16uOJc6Wepj0ZeKrOQKjyGW4km12+9Fa202eN
M2bE7EWRVPL6j5Jl9hytEoFAQHmb0+5lrVflN2Oh/p1UXIrFlMcyc/xL1xkaPQfA
Hu4JLk6PP5aLWpfj8oT+eHw+APOF+nxlKX4QHYiUqyoMptGmg1S0cz2Zy2UjFOJf
peA45RVz9xzOH1zsP8zv6Qox7NOk/KHe6cHIgv8NxK56Lob8GaWypYGHIZdu+IdO
7FidxBu2VqXdCTorseXQxLDhhpyfkHXHT1rXvew4Ha1Uv9JvjkCqkig4hSJ3PJb+
A6Fjts0hAEU3cgxtFxDIIuD3n4HhN+TPpcsNFWe835FJJ6aEUBU8BaZY/puiwJdE
XTnYd34Bfjxe4HaBzWM96es4rDa8vMvoVxe3QFXKd0cnd5GqcinN7Iq7WSjlhn1F
jOMh2iC6pJk/nXUi0Rslnj2CDkoa8KwrN8JLIZBXF+4HyVwxW99AaJYo73fxf1DV
K2zTUHI1GYFZ3J7sMBYv9UPD3QNhPdPjBWmEIbcGolp14LOJijZkUoZi4r9QW33T
N9pbGklnPlgpkrDTeFY/fEci5Y9MKYL0DGpfqMFPE0xS+vnx/zd9efWo58VbiwgN
/Tass3qpr9YJhixqIQ+QuRf4FZ7RZbugO4G8q0scSIm5kFQQ1xH6YIOYeiRcI4PQ
9Er0mP0/ZWYrCJ0FPSvEJr7eLKH+wux/+EeLf7bbBN2ZiztN/h4zL3Tbk6f/hak6
bmFpfS8aQrd7lnuitSEKv50AqiV3o3QH7xV8+xoN5Uzs995gkjiISEBoVCctwbzZ
f/hIcavsSX8SNHeQI00R4Ugm4okog10hDC1tB8Ujj6f3der222ybo1PsmpD56pkN
Qg53Yu2cEnxZU+vuybxirlGfiwfaqmquvOi3t6Pvi+0O0j8saZhxLValiPxOyu9p
DyvxYhm0VFFm4aqYM3xT7WzQ7dQ5rms67bWgWXwwBSQ/wNsnA2u1xWsLiOfK0XzD
UHpzx5WFvaCKLFWyDum/WQru+LCh0XijogKPGwZQ3AQ4DwX90qZ93cEnADZF2IyZ
as687OqLn3W5NOLwoly1pP510TCJWvNhedMYWxGA83aRXg2m3bIrJiAubfK0CFeg
Ih+xBPRw2OLTgn1+9qjkYBjI8W/CyKCD+ZBp2I/CiS7opbl4bgM8LcMjL5sJtQLp
w1nf23lVcOiDlu+szYjkCpJI/kZ/F1ihB05HWTSeVZ4cj2iNX3bs+hFunqFmrd+i
sZksGiYhzGnK9SelDmiZPknJFKL9WYznWAnbi6McMwaXbEa2cGJQZWBZOxAnvp6L
FIAXHA44TFzw4uFdMrsxPUNd6Wlk2xqy2oqiYqsa4Z8YiDyWtTImcfekXpqu8DzF
ruv4MsQ7YkzMPkOyoKDKzv+TB448xE1V/1/T+W7AeTvyjQyT5kOC/QXLb5eRVSHJ
4zxM/Or0P05iC3YAIKH77cdsiWHZeLkFiAcjfRBqz/LtH2Jl8YKEDuKW0W8pG6cx
WL54oX/3gD4hdpfLzGvXstS4zjBvvn8CUkjoWuRDLwIrFM3o7B7kzykr6dVIhQk8
iAI6l6gv6c+X1IfDaj8PKCK/udDdk518Ex+4g1jdMtNw0LEPf9xiwWAUhwbplEvq
AUemykawM52cbLoTlGrODRKNLKJjVUdDQmvjFLwr2U+U82HMVIEBjZ2s1fttyxnM
PyrMR2sSK+r2PmaXZBYgPM+Ccrk2dIsy7L71kf8LrukN3i+AywX6XayjSFsv5Nua
I8RcRbUOXzSvrEYXlq75aTAX22Wfxc0YC8IQUVlUArkMPWEUz83L/6h++k6ZZxQN
gGJen7q8DSHmwGLDJWBA7i/Bqw1jvBpnVsM5zq77G7TzbyYwzSylhXa3UJwxJAz8
x0GKaiKe7cnm7sd6iym4b8zkePW3ie6x3JeQ9r/9eaIFVykJf/Ze3a0cgt91PqPU
vcwh42tojBVvrCf6cdY+cVLbJ9UFW6MFYWPvrxW1sZKglbp3r45sOXR2/vrXu4+/
HbK48R6tt/s90i+K/10KeeB8kgbrWDtk5dtTAvyLJpwqjZtXPU12xwSWe0lfy7Q4
vhL4L3UaXwScA6v6mecaeoxUx0CU8kmAjhQlARAjLTesY25h2DvSqg6yzM9rFfaV
SBPiO++BOcSKfIbz0e5ZMqDduTTNooE96SonyAwXXN/I2SP5anTlnfmOUj6JZfEo
SWHllchdPbGc46CF5UVoIUA4pWP6tt0C9N5D9buW+L1VRbKxQHbMH8har6KbJ6GF
LRlg3dnOZTWxzSJQXlkayE+zS2ULnGrPS1onpWI1iQAjJAPiOy1qar3MGMF5fx0V
d+rsiTYzYvNfh3FkH/t/I37z4Cqntm4fDhxhif0dM1u30+injqjT5bxwsmJFFg7x
2BPJ/p99THSYMbMS05J1KzwJZJl0wBX2JO3ZWkHoDhg+TnB58Edx3bBeL/7IYUzY
e6M9bwpQkvbNMCLEzzgIkyYIEww06lZ4S3zFxT31DlpnXnJpRSvkU9pmA70QmDmH
z0qe0235keJF+UALbqetF3QDhy+DsLMZfWuZTaSyHGWR12igIlsD6359m8Ockzq1
Wrbf2lUw1HDHWJmIPpKoFxMXF3mS9rrqc23dGgFT0kShrSHkLZZNGn69F2v8yAnY
gypOFxxMsdgd+6V0ryVjk/E3EREDueRoq6vjDr+9G369kIEnXMxaV1683JHYvSax
Qe8fmOeplaNjdU4IBvXCknWoYEWGEqVflKgm+dxPafDN08l6tbp/CMEEVlUkzDX0
J7kXdgt09q0FlZtw2vnScnr4VQzE3jkrBhvlZhKjSSaVYZm9+/KmayZ4aTYKQf4S
AtkSnzcI3BhfTT1IakKW+cDpAx+zhyQ6KgMZFB3iPw31ipt51+tZnLAaGfR4kh1n
QAbsRQVE06mCmE4AOsQnhKTfuM931+w28+8Q0Dv9uczZYp+MFJ4ViYRjvHmX/CEL
reJnFAS5uZn7vCvgDtIjvzZtsYrxBXkc7j3f6cgU9raN1f4IOXgJtjAPB+GkgqfN
FHnU2X9K6JGxqSNIdjp7cYt4mTbv+wjlLdk9gl6Pa2W3GK15BbnKgNiPJHfRKmuZ
5WCzPusKd9BQZWlE4ua+YYWJimalZhVp1jTrGB+244YInS/RR2cAArmNmfvS/uQv
QeVaTBE1SsXeDfYn8zROzBl/Miy5v1R0BJrji0J9IjgHFQBEmoOPBoN12e9Nf/wu
YNyRddgCp5mhz2MgIsqh3F6a4KLAdAKa4EP3JDiEEbh9MK/5bLsGPkX8/LB1z4jc
V1YjpkwnkPipJ5QlVx0XGWJsPHcZ+Vz3N70AAcddmp41RH+e52k2hGVfOhvTq4ek
dqqxPAje88TS6PG09CNYRFkjSD53rPVOaE5IQCIH0DkHXykoS9tuBoWUGjd3I4tu
1hQcgZNNYYhIeQ/3id+e0ujTA8DjuER2KId94nQfD45SfZvYALQFGx86Yz3SC640
4mvHSn2O3bblA75F9RuHmuK15Po5i8NpyTwl3jGLSb2iLbO3alKjHbSXBQi6W8bV
jyGD0l1YgP2DMu8JfJ+ki+dWVgeHKcjH2clC9o1jdvO03siCv3jTdpfeJV+Q1s3K
RJ6ixJqL8gucjQ3Y2rhRSI2EV9yu9bu6sZLTpsDseo8b/6CylM+fAsbcmApAyQx1
Nr66Xyqqf1OOeYwOboqasAVvcJyC7RIV/D9HIVyq5YgEyewNGLBAtpS3kEysrb1o
rq7Th28QjGAwm/F3aGBzOQLBkoRsMHnBaOXKEUCn94k2fDN+XzgQZk/rG/9I6D8/
4ChZ4ozMIJeT2n5iaM6ZIjEIuuZThCwueKD6QyPtqZsjMVGvN/71arxiWcx/tm+r
wAAo2sr/CqIcLRFoQPeMVncGH4xzHngOUSSGcvgAIcrNNaq/4h4CaiZUwPPQOrac
x7oicXRPsFloutLEXwmA0BIjiRheHyjdXvyESxrGGuZOJi3XTIVYMuJKpOnrXlDR
0RXQ5dvfFuYJgmQI/KVWRtHw2zDJIaTIrQLsPkoV1B1kq7Ew9zSui4q6lkhZu2yW
M+iGo5exbKN65rOKFu4wioS/VqOKGG8NhuDO4bEPer8Yxphc4wlZTbvRKF/9mkKR
jIbpodyvbjSLL2AiH1i/Aj7Fs3I6TvyWOzBtEHGCWrKheiqLiii90y2tt8Zrmx/J
TbMMgO/ksRyKcskRkyXHVmqWPNl944/o6zY1QbQF5lajcOj/fWk2+v7L3ORXsPp8
7GgUNmw0gNe2McY5ygC9EiVvPhnh6oUceE8XbqtGJeuJKngrP+tftggxMg/7fvbe
3Ex1n95HBEkrzxOYXmWQSfWJiiwY9qeLGLh2klaY2hjR35BvoJqxoOp+TP1rYvSd
Xg7s/tQNxvqD0drbop/9AcP7AbUDiIaAzgQAi6ym+ZBBsV30A0AFQ6R7aBN3BTdK
072NNQ9H1UN5fy8DvzOd4983QHxwzFkz/ATIe7t0OZCBim7MDEjlmQcQ1Z0LweuS
HPattNkFKoe1Et1jBIPiG9zrIBqn5aR+FNnGm3icQbVsEPgUqA0Lv9t9iUTyLoGu
WsvOFyALz3jnLPoFsQWSsRxLNa/A3nccS4St78dROf2kq4i2HuBC1GKd0C0n/WHr
gGXu7pdw0aVDNOFeEUNSVSJkKBaVs8a+rI+UR5hsUIjfbgRc8NmzMPprrErIxNLT
iQnUGpGjUvoPE/4gll3lR+syATyctjiz2CprWCy+UGaYq1nY5nRn3a+zIKTbKkx0
gwcNjY+uFlCu0dEtVl7b8Nv0HOc5hyYOkeH47jnI9NLBQP196G7aIt8VT4xpTbFz
Eg3EZ4CTozWyByBmTcsJeUXI8cTcyn33zCSEKtISuWAhESswO0Ltr2GJBqkyG+du
sspwhQNdVNlohWcaFX9aMrvyWc3QH0gjyNgdRun7Wja7/0J5tqEcPmlXJFtesVNM
282IRLNp6dRwBlBLvL6griHNsjSL9/CNqo/sQtz0UIue0DJNOJFZ5aLkCz68MSdJ
k8O7xPRNm7Hj/qEp5qJXzdUTHLkRevI8ALBnuIWHwEONqHaiKL+jhdk2Z3ctjEGw
7NTpSlEorS0XoZwzjLsqxA==

`pragma protect end_protected
