// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
XBKSJfgbtupwfpO2DQmHzDqVZCjwgwYTKLKJUCNhlP1CjvrPA1XAVj/b2sIzgetg
ePt+gXNS6duQeFNY7788MZaNniij2CHh/ZAyZnD13IjvhgZCCDycYv/uQcdWksxq
eZVKvGaa3FvJ1HCwapeTaPTreu4ZyUwZHy9h1R+2nzA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 3792 )
`pragma protect data_block
/2v3ZJRriFdpf2sf1gNS+rgGrN1vh5A7waSzIzOZNU7GJpJH74bUIIh8nIm3qr7h
2RjiraSu37gQJjKj2P4vWL7rAk2LlnrM95SE+FYN+UKArZ0hYt/K9wXzCca+YcY6
BF7ipYa/lqfY70sepI1UB6sqmgk6fXgBiZ7Tt3FUk0Iybe96g/6RWM7uycXU6A6L
jKabAPdjg4I/y7awZys13JbHaHvEANz/d8v6kL3BVWYU5MjSAlIrEtaFb7GC29bl
yOnoFTTJi1FYzeR7El5bPrqt4jAcWhAOM7dWdxTd+6Hksw6mrEcU+IDOMtbu62fT
usMMgv70LJqJVN7LlhplLv7UIDXJ66P8lU/4CbGV+UvfDQmGrwBHyS3kgPfMD43a
pvTGNS1CdKZyiTwKRElOtht4wcKP/mAtk8HHcUz/4lg1pdGKEIk5SSIWXpH7BC6W
C5NC1H/5FJ33kV5f+S+PrNVWEiv93f/e8+7QBivIqjU2qPESZx4U9tVCCKM+CiEb
mkEU8WafCOgbpfEpGvb7ule98qgZcCmsUtp2AFsf4jSsbY2Tb3WoBNqbLjALzy+A
J/uEG+pzjE1/2xlRsVCnXHvLxs809KI9eEvhb/RaBYViAtcZRvQN20In1l6/LzHG
NePwY5uT1y66dMKbyAwYhW2+0FLMQ8ymhDpgeqNn2NA7PehJTwRWtxNapDjnXum9
D3hg8JfLbw4vKO6MylnCeEKUdIuGV8yrXcKjUE5503zLXn99VV77jGpVi8c2uWaa
GuD1d2Vkx+3c6gVpV2LiTE+KFxXcG9gEO+XHd0uBN/u752QPynRg3mtAKEXhdNXy
/LawvAV0/lqDGn0n2kNIKFecSZD8IFCK30bW0zf4dfYqFGy/fge2pR9oZXU17NIz
znr3Y9CvqYmhcfxa55F0aJFLDsVQP6xd+6dG8p/AdX0HhKPsdvGKcOwlX81KMhO0
8qIVtsQXuAgaMZha7JZbSYduQJLDKYa6Q9v0xKbSY5o0wQfxKmY2vP82kzTzLjOE
kl3ab7pSSD3oZsnVK5l5bPcIih6a40JdxzZ9VaEyiXZCv61ids1/iJ27kI37KWst
S079Zw8vDvPjNUOtU3ppiFCPunvHUSjwHO4qos/rVfUZ+c+Cff8WOVi+4thk/YsU
xhAQcMecUs5l30ivDaH+n5K3ERVOGK9mhRhna0qS/pFapd7xV/GNIz5fJFfGP9CJ
0CFXKEozt4EOwUNZV7NQiL17PIjP+izy/h+w4jFCE+Ac+HztroAflYOBPDWrg99h
g5mbL7svyJu5gymv2DCYOHDzogN77b7sGNxG4aV3Sc4z9zLEIEEkoTlv8g00fqw+
Lw7lF+mPHyzCQAZCYVDcj9z6wpkeTElP+eXP+c/WE+S8SA68w0bvH+hCilGnzLYi
GZMQG1i+xQGLkT6VPYGLywTxFBXuUz/TTQS2qRZnEgEvcRGkgcUU/5tZ6KmKHtXp
3DNr7sqqktdXmmV84TDUJ8NOKuZWdTKXP03n5lYVGIljhZsoAxUFqrCgHvAHN9nQ
TlRdgi0er5LV6bfHUh7BKE7doIbm8xBzyJJwGpx/Ydj1k7lzBnRv8/l4G72rY1mU
PoKs59rNtIM1nXN42z78Y9HPLcDUA2Vkekj/lJKRUo27sAP18WtzpMUv3pO1tOJA
K3GTUfLQY/Cu9vZbrRS+PTtzqVGulk+297xYeuWe0hBofmaB7al5DPqzYqXUzhJr
ZbfmxsExf2ZikIrvvqCR7yE5DegwcvCOTxqYnbCuECA3nt0bXs7cDbTS2yAKzbie
9KdsYPUBmxrB2g56zi1nh0d1FpkrQPfCf/IkI+opvsd8aiepTiXIeM6zMeKIMdOv
yj9YC8e3bsX0qINo8ixpXFjeU84qrkDQwxbYicqVuhOo7NCnFEx5agKt2Jcaunaa
IHrwicaEejWoNLuwV6GV8AqIP5BLAi8EiQwJmdhc8me2KP9pB3opK7S4IWT1Pbjv
/6RO1R9yaxDWgoMRpQVxvhWJ4F9jIm/ta9llvBwdW9HnhPXHva75DpDCzvpz1WPe
bwRmTAJ3MH2MfpIU39zUvpL/0gSZz4zU8GgkFYOGIKjRkPlQfQwz/d7Ry16twy3b
e7RzeZsIg7uxScezE0E8i0i1FYlt+c7Iv6dT4aULikbIbOwgp/FgmmVXY1cPHXQY
QBasgfvb0CWQnCHPvOQUqvLM2rc1zkMJ0ky/2lxBz/3C4lxuiNySo6v5zISqtPjP
cfFwWboizSNfwbf+OeuCTUr57IeS/gD1xlRjinx2HYSLVQoM3yQ+qQK+ow4NzeCI
uwWA9VtPUzi9hpNVZwhA3nEnICA1yhX/PWh+G6nTvagEpQxUAUuB/OCrvf/KICP2
KHzO+nenWJwZPVvU5vgg6wW2G2fBRZ4ih8RLfrdaqtamwah1HwtgNh/xQ1fzbCNL
CVJgoVtE2o2m5QkCB0amOfH4dCFlZ7Ioo4t3XGIelpzSV3aquZ9MCzenZluvxwqo
W59QfjJLDuBmC+zL6mOdW1Uvmcw/7BzxWq1dzn5Q0vrTSzAGboJiTa29jTsSCyOP
0+pKYyI8hWt13ove/VTz9Q6GaNZQMIXi/rv+EsUDpkhw4wXoG6Nq6/yiJ5giE63y
BNN1tRrrA0XiM7x0h0g1j2WYZQSaTT8BiEwXsrhoiurd7ADWCGNJ/+DgDgMqEhs4
z2em2fma9DudzogzClQh61swOIiOpFQ+Ke91JjuAMSP2E8ae9llNs+PKLCj4hbAs
l7QpMRvvhRNEV4O4dDxtigW0VYyigLUV/Y7285J+cqxMnJwE41h8FAxO+B2E36AI
4dUwbzNecMZsa+R3GnUabz7Mqz5dbTCekKtGvdxOk9VVSBg0+mo+4xnVIeh+kKNR
q9UHFhrMycxUcmqXNdlcN0bhGlPfwTMXkN0bobgQCMpUBnW0KNRoohCYr6FUljja
oj4H8tU7TwGc3/TIql1t2MvbEmKQrPdl9abCx3lsny8rrcfPBJ8F2GWDRHCBWwHd
M3Kcu9FjsihUiHE/0BZXrBCmdCm+xGos9vT5vLXRA0EW6NAUm6/4you/ACbmUa8+
/zllfR/NDb/mbA54cg38K2s4IRSviICM9ceYEbI1dxEsvaIi9r2IzPvQA21D7noZ
Q3FBPpSoIN2UhX9Jy82D3QT/M5gHT1b9WH6TGBft7YGihIedTWifpZ55OdLNxNj6
xix7cp2Y7xmCSG8Z71OrsvrUzjTkBqvz3novXPECm+5XKaEU+O4qmHMgcvJs0PdW
SPaLvI1sHz4wrUWg9ZOGstondtS/p3Z43rfbDGlHIYMYLE4TwHr+nbO59DaoYJpw
4BuMwm8F/mcuXB6HNWW8tjiHdG8qZXA5A5dYSSHcbg7a4vg9K0NWRatuxartQD+F
jXL8c2WcKPhBFO+9RU5GT1L+Jgs56CIXnyeNBUlNcYG1jpXKS9sX3qizvUVgI40J
e/3qmREkbfNTnq5UAIJtYAvGFF+JDCkHTAbt1A+UZ+kGAOnWBnZT3R49uNq8DprF
+dJTIbEhc4td+CGVeA+2KxVYhvuh0wcrUrA+il00U7TcaspU1o2JAp9Ynuqb5Soy
okfEeUcDCQ3gX5nQan95nrR8L9aQhabj90/yG/t6ASPpm0FtTfU1FM9jL8ZUYVkl
Uy3PnH+MQaC3gLtodUmMW1MW4AQHzaK1eKja+EvEfDtKfwvtK04DeMsDoN6yNFHp
ulQDs9+jvrtTLjqqyja5gktr4WEeWgR6Ye8CSizcuxQA04K2swxr2gWsbyfWlCcA
x7+vqbYzG8LCe9EIkZts7Y3DOW/Y6jPCWV0w5c31gftHXGn80KmDNZtNXMHhxK/X
IgQZmeEGTc2nc87OYiPEa+Mfr7dEBbMXNCGbiV0RNj3uoXvnM79GPYagatThXkFx
XZiliwJ4wtzp6nu304KWid3xtNB3woGfTZ5ElK9dvIhQ7aopiQilIehIVt+2IyPl
z8ebAvaGUMcbjUbnGILkjXdzMCgNsRR9Ntyjw9E+7dE+HmeP5IcGFpAwgNCpIWXu
iiDI/kXYMzx8h0tBKVflwhARps8xjZCxOXopv5GFdAgarPsTv0ZHv+jiy7jlwylS
XEcAGZupkcis9jTdticIlkRTgd65qN+soMhcctZ3J6NBkyRUXtDrdMU1tcuX/jHr
GORDkna5tRmYzsF/uEvrJILXadWahwIbsozXmV/5KULWCBiGvuykRIEQJlJSFp72
MP9kGCSEWauTnrn8jdzPmDGsY2hf8XM2vf78Vi+czF2JQAenabFdOjKHgW4qFeZT
gWMjTfcTdnLIiT1oieHUUKKjHaY5ZeDQH8BcXvRDzvQUkvSQWHuIQjBxK4UjECUw
7UMI2awQ2knm0t4p8BQUa8fyNFQP/6IjFBQecKeJiqmgOgkXvYz/+8l7WgUywhMx
yc6VzG7IGPyC9+P0/JDi4C4W+aiX4nMM2bYWX8qAQ4pUfTldZUIBy7lO93PnraSr
Tln/es3UmvDjgnjWgTVZ0oDZkdumaUeanlYQPDYL2zt91XYCXXsZMMiXBWOCEA0f
44jeSIYStLS1WAg7TZjPOTFEm8bDrmWJKUDMqogFaMZt738V5IgLH+VLSEXwxPu4
gNc3Zs8fJjJS2oqx6ryhGeOTNCGL9VpyAJweOKbYsS+6qPyjUrUl1aOXO12JYsbl
5/ZG4aWmlz7laUHWwJbZba2WWUYlyPxsnpN3gcH3roWUp84LJJP3PD6FE9t6ZcH2
hw3AsxwJ2G1JPjTLOyYfS9x8cqI+7X0DUUo2REpkEhJTfdWqT9FBbOLunpGe70c5
E1iC6RCMY7T0qeCEPH/aF77WuaUURBj0STehON1P5nHtepnLPg/T932SgGhlaszh
y/ZIcjKI5iXhtll7zAdxBhrk76TCpmXhE06OVZpLBA1oZfcxBEfzaGTA2rXTfhrC
YbPglwfMP069E6LR6DYVc/3+wIEJJ+7TUMIkNzofR3pG/pSrsbSXm0pP15iznZhY
AgxkvmfxAfyhCm3Y/zHUjKRywaZzI73tMNnlaoJoXkSY7rWRlIWl5/8UtVo2Dl3k

`pragma protect end_protected
