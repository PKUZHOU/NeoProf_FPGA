// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
edVIkmeTJt23i6FfuGsj5/tEB+38IUmlCyV+f/CYOd+1pufW0sUSE9xxCtb+
8vc7fdeCDraTvn4fWA8j7h4S9d0SQvofn5giO+IpoAeH2nPOuq6ylTi+wtEn
H+qbe2b6XkaMzhG4CgNCB0mIP4xIkCW7T6MAmy0l0x5baZTdz4VEEK2r1CvN
4WK/Y7mMcp7+EWsUggPWwsNVeFVHhLwQK2hIcKgdpM1Jih8+Z4nP9CtXRen4
Wlg2O4mi7lL32xvL4J0MMml7M6VX1bUsOZthklINiH81CPs4jpIGeFPm43I1
KJslad+ACIYlG1VgJ4pVlKrncKYyAdzhYTT2Pqfdxw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
M66PzYAY8UY/a30tlNltpeHOUptScKDi4uL79ViOQvxVow3+GhEUyVbc6Zoi
rtv2exo6vgx/XJwBAB7p82CqJG4nrxLKMEo5MqF4imyx5HK35ILnpay/QYtr
/iVnCWrXpSg2POtuoEgBuLDljRqLISJewjOakPwecYkft2jNHYf7rhG6zapZ
jQjUh7qXp7Tr5G3C58oA0xO44wpBkYyKV3DHzww0VnyMexbkUAldicBAjE0o
RPWoKYnDUvBIproxzkPHLwxX9/DYEzNyLDxnJaX7NfD7dwDNBgxLZ72qAYnr
YdkFc+ACjEC11jqLX0/exhOdFuSqmGf3r4xkNdDt1w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mTVCDW34LaifqaiprpEc4/mu0ujYY7lbmDREKIl0a+BYNAuJOpIPsvulfyd3
FcVbADBSHhZvsvYOOoEato8xIHyYcTs4sy26F+BuKi8SRp4KPIMiaqhsYnog
z3EvDSEiOfm0AHgyH3kNVktHGEQ9OlXpyG/+1Rk1XZI3Mup8FVi1LBTeBPek
95yd9Q79nLqslzzoZw3KWiNt1nG9EUqrc1+ECgpkVzl/H7UNzQsbBHG71NTl
ThoYhpl15EBDm3LX6l2Rg1rf1pgq8tm2tJhD+XLOV7JgMZcajdYTJ09/+h0l
JL/5z60eINRe6RTE9ZWYzE1kd8rLInRRZ7dAsE+++g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kVo9xQsoUqEAzWRMnAJ9DCvvwJ36uCnsZ5HpCt3RR2gba7DNmr5JQtHRJxYv
09yI9o2wkMof64i9XILg85PxVcg6/hGreQXOINTcjVWSlNuoFWAU2836lYe6
ChPqoFHecTj5+NdxWviCNh5xABJ6tN+1VkewGwBOUP5ush4WrC0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
p6INhRE0Kdh7u6gGevzSJ0EZVt1vX3r2KliCTxbGJPRXbyh0QhcQTJCpprSq
clL6YrHFsq26Mjbe1/4vduEezC8HeQVjN0OUSzdxH2kSU7gpaV7/fuaC2KlY
xM/ozu1WxOZFH3qQIfHPKDRDgY0J68hR+dxKUbZ3B3892yGJHcuGItmAwgHm
yWxX7PXaF6cV2AHZk6IHG0MH6PArG5Sy6+Qm0xMZxW7KZZZmNPcx8Wqx32ZT
2FsZnyvE64gOXgDSxwEdVnldZpVxAt4MMPGIZd5IcuiflWwpDprqWv2Nw8ov
K/QZyOWQFcYgDvPEZjeHibsKlbElOfKHkOmY6t56C1gwUG7NwNNnMAGhyCxG
IWUWCUXOFy4nZ+HkV6E+6ZkryUJGzT7u3s8rOnIZMsw8XFFR38d4YLhFiSGL
wXzOzwdG4/xYYEcjWYPqqrmDqDFulVPNcIbH6RrcieteOocX1+ZB0Tod5M5z
0K9JXoBdBEkTfqE8z+YvImRuWZIzTYFu


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dovyALPbvgtG91TEMfRap9SGzM+uG/hJb6TL89NdNTvF7rit4U/bkGskwy0u
nOjnX0q0HhUabfPAJtFVIHTmxVH0CaqH4yOFViZLBQz5IU++6Y2FTTPLadPe
/QXX+uuPq5Y+dSlRePLy9wz4D9JQdrNwUUAUz9py+1grjP8Mieg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jvYWQHTavGsT9rNW9hZHuqK13sG2ocna2LMzubR48MfRQPxfvAqiDlwbQLzu
CKium5dFI4/l5y67Rp5s4upZXRh3X0lOGL3J9BNdLuBaPf8y+stNhMuGBGy1
AK0PtMMdFpXBXTb65IgQr5lOfUkQP0gSGAcE/1FG7mg1pnL5x/M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16064)
`pragma protect data_block
jWY6BjdrqlytkjxpOfkGK8T7P0lQ56jtABAB7TEABVgSpSEbxANBF3g7frPJ
7Kcgtm0vbOdcW9+c+vjyutIHhese0PIPxtvbaYB/u+v5Pu/SMl/hPf2MKiDX
tMpkfl6zRL588O8oVISfyl4YmsExQnIDChGFWsAokNTLi3+5Xib2LiudavpU
US9Q4x75b36HzFkAg2zZQRcXJTX3dJP5Z4toIG6IhZKIiwa0LjrlbWX7sC06
NXfeL33h6tYPOt2lhNGbdZrEboczNINofDwdJFbRtoA6DWIxFVdifoVPzt1w
XiqI6yR1VW2Gm5ofv6kFHKXwQt0UOrRE2ln1sW2RMvE5XMZcduvNiKNwbWWq
PFSF++JGRQUC0AjpPMTFIpBID+6ZY3920T7r2yZMDr4560j8ZsmgjL7eF0m4
w6p6dWUgVA/rxOduUQOp+jIqR9oHcxoIy1PjU2Xl/MZwiWayhTzl5mdHMAV4
aftKmFusIAhtrMXaxDoh1CGC7v3jGEHtTY/XK17Ik8SjnJfQuDa/eQn7U6qN
ecLaL6OMe8mXZZmy+2cgBVbSBr4Prwzfd6SFlQskMLbjVFhRcre6NtoTkbfk
bcYfkj/22AMtiAV+h6RAYgB61ZhsmrfZeVjiihfjHyT7tLmDGzfJ8GfuecnF
HcATDvghMsZcohB8tvOT/wdlyOu2Qte+P3tEUOowtdTfjHaiyNWPXol0UVeE
hs4P1hT+oX6A5VdMQksFkSRUfU2QGRXvt/nzxwfNmaWBfk+7l/rpOQz6Rmeo
RgQZtsM1lQ/rJVs6ySZJ/aN4vKwcV+SNVqpf87xbLc6gNNxL5BPSw5uKuWKX
0hzAPXY0ey9B6/0dsroDo4+o6hDMEUr8Us7fpcHeq/PH7Pm9B+ryJ2KgV//V
gKWFb5yXsmejCKfNa4QWga5tudKVfcE95x3dsGdNEw4WornZk4TNMM3bH5d3
3IQaum0bMyjDF7nbsxaEJx+fvIGL+MEx6s4GCYFBsLiawvu29DMuiL7he2Xq
vbrns7SXmByPsTsdBZy2j0Of2jNQZS1FhCRM0u52kXdbcmnsM+wcbzZJJv0j
EsLHJyxjBGukK0oorKrb6TrP+jLyE2zGaKpWRlkb1ucP7o95RcYrHY4xKPIj
OahpeEnXIa/wWoypyMCpsneBYMFSlv0R38gsP9dibzxuaYzCokXwA+Uu6Wjm
Fyz9har3EwFjsMVW7nxSqbHpwP244ruLJW0tYwNR+eu6rWhDnDW0htMgdCyG
qih0jZFjW0AWaygRG6XFFwkfGDeuzk+m8oEjVE5q2qOzMnEKWSrSSooNvpi3
hjveHFj+QFXCf6QS7hsfIpAEJL7wxWKHVF3sG87lCPASedFVKMvod+lY10cD
EFq65i3xmvYK6ZNbYAPDLeAUCb54fyqmqpKgzkTghUqQd+vwLnGqc7/oVZb9
FwluCl4zQMpokbFZOTRldZbwdMQo+2bxVHVTwRQUb1rJqRnvNao7HntilkSj
meD17bt9AybjR9XRPR50valpLIf9ekT2YSUL6W4FTbuo84TM1hsG2/4ehGHv
Fbz0ulCFW0dLtJPN2lwIlHkAioK9VTnRtwXasFqc5hfEXZm+bFc/jALulY+R
TYJOm0ic7Ft/ceRjdfcqGODXZVHzrfEneR5MwcKRWCBAfkfpFLfKFJKbe1kI
dQ6TswePegDCpMFHai1tJ0Hz+NvO+VmVfh2OuHkCIIqU4RewbX63v5oyEkg+
Vz7JA88qojXCBfutpitXqaNR6+wlILiNRzmoJgRgd8G6vcELqp9mD2xl0uO4
qSZlLtMpnSyQNlwmjxEyAxP7f1gU3WQQ+3Ab3Rs+u28tsmGMNKV5R1YGxbCR
sPBovBgZ3ZJPbBHrZpfgSlzFGqIRU6bHwcrmxHUubePlgLQyoBG0MYDyglaI
AE+Cl8xIIXkjaPlzBRgXq2NSrOVsPUvi2qbw9QOZWWorJ+y94xYegP0Zrnah
GpfAs2OBgVnb6KDTMaHhld7w61TzKonJEE7wVw+d+0wPdk0JWT//6cewb+Cb
Xeavozsay8Og7/sPVQAWKq2kEVWXkzqKQiLmeUZcMbChbxOfUcRXue0mK1xp
o9XiiUGa0Ufdzj9/qku5anE8z8RQ9X1CrrOmGvC09hY9DGUYtg8CrVQlPZ2V
gG6UVJz6FIDUVnrIduP1+VtasREXngRs/TElDCNTBV/kN2xFs3Kq45wZzzJ1
/yU8KTjV8Wx9+8CAKmnxtwrLNcgFeyUpvd/uGwWHizJizKtNycsQZOc7RsCD
oWDnjqQPvviDp1bMg2ucnRw8+Cw0BfP5gYnuX9vgsUqyOQIlEy1f5yEC07eJ
j5i6GwUl5yZaBd0GYiwEwGOUNG9ozzI6MdYLC2S9P7Xzp/gd6sU6V6nxP3QG
8jxxCnE0jxhTZCTaVrw9/ivzzYAiS+YVB0VZyJZpJqMVAOvjo4QReXi6zZew
+WaXFaNnbi5aTRx+1XrExSA4Y1mOJr+C2qLmixwt7B3qy2Ly3KPn26EgOso1
Nj5ACaMx6ibNvQW0141ARTTTC1Ws4fFJK0wpcdnGz6zz7FascNSrNNiCJqBt
mZuIDxj2taAIecbQtj4URN7+QA6MRh55NpDY8GBGCXF1YYky8KLaOw7qJr20
+lZ+sUZy1lllvQVyTSx6LF6b4rab7B/tRmNEF7nJd0bIuuujexfcaZgyTpf8
GsOZeW76+abzYQzvRfiVotriD3/N3MU9fb4LC/kQI7OXoTVHIb09t06kJaez
Cz/wSC83RAwjkO9QPXVh8+BhPdsvfykKyPSo565YotAXhdV9xV5/PFTyfHDY
rAQvEKRQ69HfvsSRwKKTRKylZ3IO9gtwJ/cpKSjwzdZRufN8rgK8zoaGcnsq
AkzCdw65nJDNDUzLj07ZR7PLNx1yFaiCD3OBuv/VNqDJb0Wf9hCKlB4Zx7Dt
Q75f9/c4nod5mfXlCYXsZxucLdFJt0VFP1c1kI8WMi/Tv6U8vNvBpzzyKloT
ZdRLc0kZsCh+fWGwWtOZdtYyeszKled8RtZJWvTc+2OphV9YlwqsB1Im1dwn
znPfZ8wwNfok8oW59n+nu9FYBstJ6f8Sy9Qztzlaxp17EHhXNhuyfJlWpHHk
3mBeuOa+m3KpgHHqJ7PZ+osZr743DXSct21UK530zer36K/qR5+Gd0NKOzRX
DmeJ1zpmG6MRhghacrdrIJQRrX2bkzZpr2jPon1KREJgPDbauhzp1wLatS29
1zinQp7VZ5oFKMIqxhfVAU8R6W6Vx55n2ZGJKsFmkB1b+/pCPHPC3EUb3M+q
e8aHilfUQAkHhmX6BFHqL+LHiF1H7GL+Tk3ql2Wv7Wf71kblN1m0SzotY13f
YH4Mepj59SS4TKLJL3IkC0nbjLancSO7f09KwGuw4IV0HiMyP1f3e9hoCm3k
/+51iXKZTMux5dqEsd0HBb+QoemzDym1KJCuJij3tcwRiauJy82/Q+U4N7Xo
lMoX67kN7VqXytMG2pCoWFYZlJfZpJf+fWFIDbCyNdLNvbDJdGMbNvco+tqI
10gjkq14zozUrg9Y566D4j7Wg4/PmwZ6p4jp+jwhovYQR7QpqIVcPrCYqt8q
d+OGazn6Uxiz9LKzFuzT8oJjk0YwyQbqty9VrjeKQM61BH2mC5Q8JCmmU8f2
1J0NYIxqrv03g8TptjpbWSnGqpw9g+kq4KO1Q71uOiuWSk+slOepS5KHsRj6
09E6BlD1Pgiy9sUyy76T/jmRw1plPLsfWRlNznCNo839a0zfGJGf50SVdJBm
va2RKNy3Bo8j+7Exv4E0EEV/qa06+5yu5BVZo/k7n7XjpQzwZksjZaLDaQSp
AdAoEWJsPZoqAI6Ianko58NwEFNEsfPEexM1r9m75FS4fmrobj3tvZ+b200P
ItGl2DoUVLDVaZnqsTJgUWRV9TTm6DrEUV5wr4twslY9SoOm73ZEqfAaVjDf
KG2ut/0QoAcLM85ceFSYhlGx9Q2btl3TdaBgjX7tQ6G+lzx0iivNwnnrxHeY
v52G9ACoGNGJ+LUoV5lLzOkhOlF6UqGrJ1beV17uKuwd9Li6Bk35T/C6aJ17
IQZ2VS4eoHjM4ESu1hjcrinhst8/Iqo+VAtItbQRlnJgfrOQYtdoLR6cZ2gI
QgtTyRjBJeLW+smjq28HtcnZxQ129p7GwflItWpJkW4AiVB8sDCA9LWV9Tq+
VvkCubyAmNpHC7d5u+A3MO7V52iBcKp1WLuqdyXuUkvePKYrfyVQRdU/oEvK
IGO+uQY9xm06oO+else5+FP0vorlzLqAHAcf3sqRfgl0MiQAjo/gmHRL/1+A
uNp3+TpG07sywnbz1l6n61ZMQhY1JQUKF/lWn3vmW6SRZRjt7ducQr4rsFcW
JHNzyESrXT02K4XaTBt2YOvHNCt/hudhbjCj2dP7i+HzM1pXvChIsQRDGp+5
+iCPNzNr+Y7p1PD/0KHClduRnCrQ8OLJYddv87QZ+ga76k+hh8UddUrhtATl
m54jjMf7DlhZiideFhe60BOGEx3r78cJahJYxy1E3EX1N7yiuMOhzjuxFdgy
UYYA6h4Ak3Yzimfx447K8QS2SliWJiAUviIFrS9CwyUgAAm9WuE8TTmrDgkz
tk5N1SzyW09vJ2DNGNy7zw8UhJEBA5PDs4fsIfRHIrP1wvovbwf3+r61QMdV
zMaCigH9InAMG8BnhnYq+imdmVMazWElKShxpgpIWErrZEFR/bjdx2epUzjr
80W0yLYQn/pP/k0atE/1UlJID/T5CufCCAxUcXk53sNuj/GvvB3tAV7Yl0Xz
dcxHR27ZfKJEIpY7UWDGIT/puJWINe9NpFzjXl5MTDxDXJziKfPHZdWOh8ti
TfpRBQQOWKH2Hnmolg6HWm1pflzq9aPvRO37Bu4rcHHc1QxfOASYGGR91xxi
WZywt9OQDuhGyfY60S9WCsyOULeYQ6QaUEUhhfBdbdnh9qGkWEHy76K71ylT
j71ZZp5/h34KiqekGgVV9wPud6sEeifOiSQTxhK0jBY0TtstBfb1nmHxMWGd
+tHXeT/8ZjPwkZDWxXNyNP4rABSTJlcO2tO510NaMPWP/E7b3GZShJYW4hCc
lfDxoYZaM6moBZ3Qy2Y1PIEJbgz0dnqjh5FCxYdgo3Eu/xjxZ45/XRmUdSOb
tp9IV3UBwtuEWwb2jRQCt+VPEX0cmIMPBgrJFaZRjnBYs0xIp0seHyeV1Z8p
n9k+hMrLijK2ruXNSiEkyEEMEXwH8Qj9IG5zIPzxzP1Pr+e765Y6AgGt9N7C
wUF1uF2oqPjK/bJvjYBe1PX1O/D95PWz1ArUJFplo3yAmnVJCfQHgQgPpEsQ
JuK5TrW5+v3T8Hf69NhMRbNm22jBCHN9a/cakH4A85cFbux0VceV7G2vmdBF
gVYF0UnjfDHxhlb/vRFGWvzMWnn4sfjgJMT9nDTAwmHt9umIvSrIkJmN0+1y
K+FIMrdadsHzVsLMNTVRH2uplnYGzmiWlTux5rnk8HNqhaCfO6ifbGX90yCF
TauqRHdzETQtD7unGlhntlO43IJ/8kuxLMmQ8F1JQiOnhi+ELP0YnXpaZkmC
DHeI7IDcLGwdkuHy1vSIEmIsKLvsrlP1tr4FIsBIcblVqdy53e/PnshdqbSy
ozsLUssX+XWRkCMpFXXCSOqEMZM0stBLmx/ECbVjyAmXfLEVNaXhVbNkgLp3
CWMqxp/MfRLXgjMHTRcmqVj6SeSdoP7ZJSYzOYfHvaCbZcPXAy4Ku7ZkVD7c
QwX65iF6euXXV+772OQViJ1qwhSR9TcJDRT44qbVQyfLSEWku33cN2Bjof8v
EI2UHcTFHzqImXRkuWrgLEBS4sK0reoVGISxE6b99XWmRZNmgGkuujAUWJZo
7P2rXGOol8oNxPng9kYRTWuUPnE9RDZ8ITruhQnsqRUDYte0EmoGzAKKnHzg
OuqmB7axBPg4cuXxMVHCRs2RKgvrpxlnmDTLQHv2EZHerFXY6Lc+oU5/8rH1
jQWVECl7i78yJlBqywB19vGZRSt5hyLILMcWyN5lsuQ4KtrGGnwZJsxiWFm0
Z8jRU2HMpIXBbF/L97Re8FX/jmfvU9bIEXQvSIy7q8j90f8KTdTzrn6ORXkt
u4xXtt74pNqqdRniSwT7HtJnAJvNUobEQq/1tRLa1SoxjikULWSUFGZBbDeD
hdqOyTfYqijPRexd/VGryqm29QsEhDgiDj6MOrDlkS8YBYJD4aYYgDeMKeVg
2xHHYwJdRnRvg+PGeDr/ZoIe+KMtWUGBpCvj66+AmITlpIZpewTPTPCbW1EU
/KBYinp6pzqzS5/GyPbxYeOSdcxqEa3aHcxG8XZgbsDrcpG3uqm0XTBMPyMx
Xy/q1JtClXqeqXzUkiveBU/SrgsPScr0cbRBTz97eefNgC9WjHrgI8cxXYy8
AvEtDIzmyIWRQcWbSixnNoFjqMUlXIzGI0oWWcSIr8GgG2xWlyPTEextJsQo
nj6gmDuB4zM0L2EOMldA1PszJTjp82JA/AuOuz8wyJk8i3bAiYbCCwodaKFt
YVa5AotkicF0hO6WG+wLsGZyJVF9AgMIbc6tSH0MDeysMje78F8e1fTwui2L
oMSpd8yXWAjubusasw4Vg/Sx8xf+KEi2UIiqM2VjLlFByANXDFHZLBayQ7dq
sBeKoEkKtf4dT5SVHj31csBEsMvamc5wg/nyZ7IN1Yg8RSJtQ/2BHX9sjV68
MNK8sSJHOwOgpPF5vj73o4spClXgQb8R+6R36B/1AC3ooMpogs/RwkPAy48A
jfjQbmEt4/BAdpBZZGE/CIHx0ht6kfoMq9sPU42aeWT59ldXUhvjdxu0bzau
0GOIrs9MfnWndLN+Kn6rSkpykWbyRWl7RoGrNNEcHNqaG3eCHH5KBhwKrGVI
BpDEIiTos5G4QWaj4vbNNUS5QLUfDv9mONg1S88ezk5fBzSQQQ/qUMSwWNqW
inFWOigiYpWvPXOjno2ZVLtQ2RKYk78jvm1eaRKR/B8G3dQ7pV6GwucnriIX
4keUsLCYbWb5jtlsdEFdu/2rRGRxM2SpwbLfUgQRvVWVz0a4GRG9a9Ny3Dz1
i6P0xVk8ddYEI0WlLyC/9U1ZVFs1+NV897Se4wofBQrFqin3Atj1V2NU/rjg
rfR5bUHAAfbeVi7f2PV6bCSzOn0a4j2ppEcfyr/FyXQcKJbd9mK7TQE3B2Je
zGVgiWXzGLdTIMzAR4+qxNBd1Eq7UU54mwToVP98YvcS/s4lz2QHJm6l/yJ3
vODWZzza/sGvJsdSYzX3Fb8oQnjLR5LUw5fifE9XnOtXuCkCMjlglBPpm3e3
i6A3rtdtXxwoM5yNsD5ab1GKBzzZ4f99YYlv4Ij0xWmeJCCCCXy+M+aDPjQe
V8ineN41Ha+ghyhYn/8OURm745ZMsu2zhF5cSOJgUd7K6bB32smmyBjBycIe
NojnSX7/CpAxB1mRIlft2CK2WB4TlHcCPuPswReCl6LMqvWuXWHr805LWQWt
D0PSviyGbmTkNhWBog3LLzw7BKynq8SadNhSxAJWk+rPLJqbMOcpBumIpjOL
wgQkkQXJTptvPLOzgOkNdJFcGc3BgOESgfFkkmJcjY4WDXwu9sjb1k6fgbL7
bwWN744882nDNO7OOtAxk6g1qLRaXFXW6C3WwZYpQ4Lvu+0XsqYh0BARZoc8
6taf7ExG/BkcRL2moQTm+6BjHkSVtYQVdrU8GAfE0XtZ4MqNIQDd2nirI9PO
6OwhwX14KeBp8+NbLRES7zsZnJamDq3btc/BHgDkB319T6gDvsMhFj4zoKP0
czEVXqUTp1WdWgw5kAYe9xNTaHWRDgeqvwg7YrJ5gsTwNTOTdsmATMQMN+l2
au/Rs9MAehOt0rEAcNbsYVfyFuqMxLzYKe9vmUNaqmqluE5EVTgut2ZClz6Z
ZldjbFVq1EZfRDP5qFuMLGsMETU6E6eEIwac381AsiA7CQBD3W3rCO0C2LxQ
EClzmQJ+RN79254lEVPr74Q2rvmi3r0Yo+brLemxn3jkjPXlcH/cZFC4M/MG
LyN/+s0WooY2SnpKmf1pkqSUKHlTmbRcncu6H07nckMXNtF5k1juNad9nVCX
UnibWPiKuqnNz8D/6G5QDW8PLOYkak7kr/793WtiU+ClrkgEj3cKcgvD4aJK
NTfifYhQPVMiSIMswFrZgkAHDJK78VXcIEKY+4bmbqXbpJRHNfdmaaRY8eTi
1eF6PeISttgorpLjaD3zzQeoJ30XCld31GSLSx13MnHax8Wl5dh+rdp3srse
i1y3eXaX4oxcSflmLUOvqbuZBQWI+IryOKwczZnpXIfCV7r7g3/XLqmWCANz
afjuYrXA+AEvwJbXmB4ll3KIcB0JqFlE/AgZhQVg4lg034sk2rWo4YoDNMBp
Ymn5vvkXIEfDp+aLFDkU4Fuv3wgsX9ujwb9IHiJ+YdhQ3AmksTyEVIcGRu8a
UzR1dE+gWRJKw6YYL8vaWg07pXKxu9bBdmmn8c76aD86oVyuOebiuR3r/nTI
lsqWB6MX09PVEYDKWWtftaNNhZwW79OUeZxBvCit6A+zWk4c4EjzldL2G0QD
oErcC9GS4lSKY+Ek6MUcOTF3y1QV8DKjz+MvJ34Kab40ljvh2UJouTr3wXBH
W27FcKedR+R4sWUbbo+6DsK8pKzsioOA/09BbJYbTElnyOwZh19kbVIpJdNm
deTH9uWvjeY7/SoqcrY0KFEhGZbjdBPz9snuJdkma8So9w/UDezp2VfD3cvp
tamR7fYzOtTdAMXVtMBywy7XtOXQQOtk1iaiC+WWRjS1vSF2Rnmb/efPnnju
X4S1+H71YBg0Tuh2skaJRCV80yFnFg8kiAGy9Td3O1qEV+0czk/W+7sIJr1o
cieiVh4+WWKqr3We5wn0+kTdQ+u/4pVWb8+IHIoeEnM7A/8p5h1A4aA60hLB
A/gnH6OIRmZc6E+iLbPRFCoZmhyqs3g6HQANO7N41rrAfnRR+k8Xh7h7X4XQ
SGVvv8FECd6i8GPb2TFxvq1eLuB3wuR3atIzWWCj+F8ZF4jJv1kZKk2ruM2D
eHA9dDZ1TrfOwXqBYUuHBW/9eQpCaiF6zJpIDgE3x1gREYy7RKlls1PhYNYi
aT9UIrpgSif3P3umje8FUjtU0RyCx09FK5phcSk4QT/LcWhsHwLSLVJ8MTJd
+fKmGTtP2E6UisfMPLjYXFOzKQIUEsCzfHJBHxPmxdgXlMnT3uM/0BIN3KsI
XXWLx9TOgsZuxPWTo/KpVZBBFZ4UqZ8k5r/aSKIhuQutl5/NOuoKhL2yUnr8
Jwg2kCqTGTx60cSVeMlP0sw2KUbfN9l1P4BBPDk2LEqX9rIdsbXpIi2ESQI3
uy5WzY1qrMBod+avnrLNdqAMwQaMxOPxbgsCN806504IktYzBmSENuATjclj
3V1ZImZGgYyzbRzQI5f6W/0xN5qWegiH9Y4aw9ovGiZaCWOqF1HQCTArluPg
tlxWI+zPmtRVG61vK+qk+UH/oXqui87Ign8i38LE4U2nESPhU57LCuuSDWSb
h0qsOi0/yePk1IAb7JcIWRXDYFTAqO+SzSV+zZrswrByOvveppqJWPoc7By/
gNSF1s2MUPHNsbxbXXOJ+wS8Pzdtwtp5wGIjX7zM6/cKRsCwNpTE9dXLgucj
p2c91wGCsNAJ0wgB7t9LLOMY9ccALgNqNyCbTAd2M5RPm+TFQUJHSZdHdjyV
hwuN0SlK3GNsHgObRWprFQ8OjyFIz/5X7flrjZv0+NQFhvJ0vbrCNHWaJCU1
nLU0qHvxS+5XqSTMlJm6zYHG7BZxMnRwCtW14VPOjoJLuLj6YNT+36h+xBP9
upPERsG//ijQFIVpB5ufTg456H916p2OjBs78C8bjfv34ACcwONZPA7sstac
JQwl4rTv3TDY5k130S1DPaHfBs+eA1/O3XPrOE/In7xeHRCkr2d/QvGhS9h1
dlJoAqxUYqXFkc7fcBg7LFQvqfSMjmtIDIHJFNbVlkqlVqz5QVyuTLryAB+2
jsWFptbXaKLkzq2yILVYuPuV3um6R6up4+RY8mmk1eNRoeSdVeDovJXrMWKX
4LiDI3MnJ8QUDiXe+XVBXdVTW0bHSZ2ypilD+zYrYTnB8Fc1XSHy8aDHhb1Z
IXBLnNEk8a2EUT7usK6iFcbkRl3faSCRbFIJjNBs9E7CgQ6qm+VlisGAcX2N
GoeZqqdOUnNmWHGn+TI+JJh83+qLQwYk1TOlYlrkk1/SjEKBuwKZVchTnke9
IORHEzoQgoE9RP5UqdV+mNGrGTBDTD7kPf8qwv2ksw0XcwMkUgEISApskq23
RGgmjD08LHiDVmbsvmn0FM2UmwL/SwI5cDpWQplO5/RdeOTVV8PyGHKe9XKY
2lDXx/jPx6eF1qS0ZxCdMuUeEofFcq1hGErwvh8M+2UvuGrpMB0sAPDykLWf
a1lg+OwF2mTIEJ3flKRdewuu6QVMe+Zbyckh5NmiJVrOfIK3W80eGFkGiRhe
vIdjMJ1cl673uQDjpa3deFZbPXAXwHIXZ3BIQWTHpKHXUHCRt5EG761mWJum
ITePtXQ8bK2owycWx4DkhQDNOf2wCG4j8A4rqCClPtlg7U8+iBDYTD5tRip2
U9hkDws2iRpXnZ06BO6szqEKBVrrdPM0vucpIf2s54KDN8fBMRbtrXxuXeDO
gQbJVBmEqBT9Ngkn2ZXzlejJ/76MIqQaIi4vVuX3IHV/dZBfXXHkEP2ZGs8+
97qwwQRXxMe/L1hSH9NwVWNejC7D3GFq2Ho69gsAJ9ejKFvII+WfNzSmGlm4
aLRI4yhw5ksIJHa+IPYIanVGi2d0tZD0qDiBwIwMZF8NJhaqgqNR2qqmSoQ1
w+0N9vhOZcsuBrIjw9eE1VetAuJ10sXK9tScIMlJq3FEHZC3hTbrCjgkukkZ
GUKmN+dajtQ851HafL359l6eFgtFVxbFqZJuj+W1bJDkEAlj8Nqtz3I7TUKq
sEDtS2vwvbVxMfwgws3tC3OxiXZU2bFKe9fEOcMiG4zpHHYjsDCPj0SHFu2g
YE4wfNIw/Uqfth1rCW9AAz/9C8chm2Oun/nRaRt17EnXAjuf5/q+Yj8vLVZv
iyNAETVipsQyim/+N+yRlJmGB9tC6QxBW9OZ/3csTCfb/0EI3G3MBer9H3un
bGiKbeN+JYHoBhGe/w/4mZ0rRUp/wVsbdoVUpKWJVrB+0FSmeu4UR72JQn2D
0HjSZq7kzyMZQVkeDOtoERC+M5hBSIK4oR8mwvrotKLoUFipC7H7gON/DHQi
33sb/ASoWL9zU2Qt8Mk+V/IhPgo4LlkA1fYTi1b0ZDk6pjjY2g/2QFCwD8VL
KDNj3jU6iBEhLbZfg/fvhxgOOjkbvTXBXiPUAo9umOiRl5q6pDRqgrh1ks+q
hGyh1MofllCGi9Zl8BUxCvCWFCSVBPSYKadFNEMBRTNBjCnMDCxKcU84Gibn
ktKevFGxPHjweC95196OQvT/sIUf3eC0uCM0mTnkfhrPfK9hFdhxgEohTXaC
PoCJC+UScyjyUZtlnlforauAkkn5T9B4ZngMRQTu+YrLgz609q/127dL3Ps1
FdYvqs4QAlnQGsLmB0Cd9cvHqXfpMjsEaXFjwSnMsl2NKh4/GPRCq7fl7T8J
Hitd29ArtcHWp4sqfOY22tJuVZ2cBQXiWiB8lRv5/5PNKEJvS6GFYn88NDkF
6nXZKlJXYqpQbwymkdb+W0rXdsVgr1mQSK9DBoyJ76q4mqm5JYwZEyifI+ai
o+25WVrTqEYmPGHsn8X/Oh9ihVtJlPrEpuK38VGO6Qbzaq0MnNG4XBa4p+3a
gXZ5ijbyoeN2XB+mipj8C13pUxbTBusa82m3JFbrdKhnTwndyBRPrr0Jd0RR
iZMJxF8Hq9PGynVuj8kF9TbWMJCrdSToVFV+cd1PJHNqsOmNMCaNqa6TL9ks
9n5BRO55SMP7w2m7z6ynie+cbyrc5cP1d7HR/0HmZy5KrXGjrOJb2CfBYN0Y
49nR4VU+/ucJTzvIp1l/YwAZPr9nbRK9hMK8iuuyn0/YOIAh07EV43AKsmHs
SOHsEzEItOnOXCwsCYJrNM1aojzM4XadnuzjSeDATdD0ZPeaNfyEkgMqo+z5
wxfTR4y+92JuU4IC4u0Kyc3KL0txvSw+EP1egplgeo8wZjTg+f2Q0kBuuMK+
QBuQlEeKzwYmhMfT0EZgOdQiLxcDZtzhnRUIENt/8UJmgMQMuN/IFZemfvno
1hWcLWr7aV6Xb4DWxOSQvw7bCkrOPyZa1UH/qKmsFT1AvJ1QL0V/yBvzc8jM
QosgNvLbOrB4G1lW18NT0iMoVGj+jOTKYZVX91Mlv10RkgQztJZOrWdl5NnX
HgyGQdfobNDDCADQKoCvSwRcllAfYnsemLFFyy3AGHHNr5TMgJDI1A6qjvTt
5OAxrFU5V7/SNFewN86ECK/+OTvn0+HwuT229uKljy+w0xUSvHkG+3Tl/wP0
oo0re+5hP0aevyAk9JCaH9n20ceDXeasd6qrPOLBft8mAm3BaY1TReloFY4i
37VnbuvI7P0KZdurf+lwtSpmVNgl1NJb7obYZn5L2HwbocQLTESuJFRbayJR
iRn6uFBY84nuNtCsrYBm48BqqJYfE8P4Sc2NIhlw6YzDAtTWZWZp5nAkHIKd
bbiGLdrh8ow3P/cddlbkCGTKbmvuv/L1z+Z3Uqb8ERR6iGCULiWz6GsYlwZo
IEAlRGlbkNpDUY6iGLCFhoFL8H8twdvjdbuyvq+TEi0YDytF9RQl82JMdMM2
AL5QpqYUv2MuGZIbuh238sz18S9dcGFeYkbBW/lvuyZ6u4tC3gnJ+oQr85AZ
8oIDpgNS0K6Bb9hymzEY4HhNzE+T1jp+PHQ/GYpC85ae4xR2T5U0qDL5yY4o
a0O976x8gCuuHjzW8xribWNr1QMvyM6WjZBSLk8Z9uPWL8KLs5ABsiDxOT/c
9MjlXfGswxoD6Ph/Ki9iIlszJ95D1MFx360RSIsGucMJaaPoBjx5nCY9Wojc
r+2ormNGYGANte4sQGrw8x+Hv5GMmjpalTUhe88VTyMv+9QAnwY2aMRkITDJ
hDNjhGacOscVLSkXGZSZ8Wl2h+qkNun3pgor0I8Pe9vK8ob9ZHDewQii5MdS
lgOPbUeiJ/QvcY+5xt3XKGUbgWQ9qkhv0WFabeoTz3m7SpYWvQhK+DroBLfO
XAQVhTvNYHQfAMCQzHRbEilCFm9F5dDLEc8pJ2HlSr0KRj51ZJBgYoyxjf2s
9ToRKlprOQUNi1Yyvlite5/AMfHKD3KB+ywrY9aSfhq1XE7Y2+nf6kwOO4pK
ba0Hq4xFbUJvVoVmHZqCYU5aAk9gQbUWK0dhXMIFgj3J+b9a8AzYWytqwH0p
Ip90Q/HhPxbmkJKoZHhGI8Kr7xFGDpv297t4QQ+xm1eP9xD8f9vdbUecLuYE
VosRC8LivxYxFu3pgCyrt/cL0g6ZQeSwPLoPkp9tYk1yBkn5LovY6bAMQePV
99AuN6PaAnCzoJuSFEdNq4BeVdG8smO3Dm8BBZrZQbOedK70EfA0KBNkF+Ag
9PbDnP5Z8xpSwPQ6/7AYriGZetYY650y13ogDJjFzy+nFh5TuixrXXuLDhRV
rmFlWvLCx42h+v6hNS6KrwAj6GyES1L0rCMxG7LTl6jTdh46x1OYKpU1GkPQ
hORlZL9y9Lo6+rqyyDOHEJAr395wlB6kvW4IjLuU1H/RvjUI2U7cG17tTI6Y
MIkPxjqsrn2AgACZy7Jm/+4s7yt+FpjR3hwEDcogqwvAyImLna0P+oZ1KiFp
KjmbijOwl2fMvbhLP+xVd57/BI/lD26OqPVOL4TJG00mM6vSfJj+OKop5yXK
RaNVLNJOk/clL5srERv/R46tP4rDUaJ9v7VjvY2Fd+R9Jrcwp/3slhztAQ+I
pkFD/Qe+kN5n4ba8ADYIRNqBNcUFNtr69vKGIhufykM3J14jO1/cqcg5bjFh
nI1W6McUfDLqzTHSLVMySBuF/JwEO1JVErSUXSkcrMVGnSVUOcPvhTFvM7Kv
6RZ7+cSAYKmjWblvFkFCuK7L88S80ps12Qz/eshAHL5bPCShAqlQaO2v7+cj
NgNysu97xKhszPIdHfCGYLR1YRNg4Iu8NPLXp2WCX7Clc7Vc304+RrFmTe40
YpmfiXPoXvnG48GSTDQYwJneWi10LFRLkv4hmhsuTLi2OeLK8B2/bbBOhWFf
amNq9SxRdCNZsDeoYa10b5K++Umkn9wZG7ldwZL4AisKoOBz2YNabg5lecxJ
O2g1iPPnW4xuU5vd0/j7NvkmmJZoCuHt7sVVL6N/G4UFGHV7UNvH2O5ER5dr
2qnB4Q1a+mPqqUAR3r7mObnh42GfHtFdRoR4WKvp4nTomQwudqTsHpsT4kSf
NqlJiuakttXV98olJEZGzXmInCYwlNji8Fr+CbrwJMyosU3UiTVMqwx6pcGB
udJSasjqb8xkYHY9qTSmhb+mqtaA6U9M5O5TAA9+Zx2nK+WZQ7NBtr4Xdmut
CPemOk/23vtaPxt8u8XT0myhOvxHX8JChzUQ5FVQrRfgdnr30+GEKHt1cMEO
tTLr/qSh1jnNNGoDHQU2Q9yVx5IGsbsspKEC+YNoKyIR3g0RWF4oA6D2j9Va
/a4uDiZpRvAhKD0CF9dK7d0rL+vWm2vKUJ+BSJn4daGoSX1znc11ed/pmQ4c
x+aY10A4nVYEn8FNYqf9D2Ju01wiLeDAypPn+uPG3xjdlxhoOqzKeBq6Y8lG
AGCywyizOdJYJ/Nn92YZB++LS9UdUuz88psG5UPzJmk6ehXD/ThhSq5pC2UZ
9IJZpz7zGOFhD9KjDLFXKtzlx909h1jW/qam7QVoJZUwPmiufmHqVmPK7+Ka
hKjc8ci+KJAC9cRJ64h3dET7XHAhA5T/X3Cx++HU+3zRPcquVq9LOnImGwCj
zu6sXXNCvUZXQigr84wMsMr1OeZ+XP4e7aHJ8ecJTI7VLWURFssym+qwf8ic
kFc/JNAsO6eb4IjtK+igDDbNrAv8Y2oyByBa59CBFPm5wbRS9v33sOW3CkQN
nH5/NUy7WHbriBQnJyHPEvvn4iV5DCVPxd2wGHrEiQIElM5qh2V7pC4DlUER
rJ8BhosH7eFK4XRNRt1ADV8fKxwJhPJveyPW3O/4R4Hn3On3KPSDWaE7k5PQ
wirb9G3WnD8bwzz/K+du4DnZoDYQCQGEufIkw5tYYyyyIBEuu2v02G/HB0Tx
Ju1nI572DYNHprVjbSRD+NDabdKAHZF42gKhGgm9/ytI3dXY9z0W9iYlIfrc
4YNdwLT0rvQvd5tI1jb1byWSKz5lMfTCFxMDoKa4mB8kLEknJhOsouDfrVLP
Jhm0tlv7kDOJJe65PAuMHQtH+RLhlnv5/EEuVeKnpcwC6t50FbK93Ag3hXwy
mOtB4GesN6ruH5hFMJDph+MvHLubQTCAEK2f46XsTy3dS8treud5OTtjA0Ck
751x1e2cIVtINHQCb67XewuYCzZYDswFpphs6luVJQdl0S84AbPgdOQkmpzZ
2PFH1M7aqWzntA63pE6h1mmG1WwjYKUf1sld1oUiulvz18DGGQXV8EfckR28
NAiJckBmPL3X3TkbNEg4YxnarioUcHlaSNJ8urR5m31qSr3zzhtqeDVd8XAO
/s6mCZ5MyS5/Q2aTxGgEOvC0AYkk8I0Q2aIfiOwxsR68a8w+gNHY7Op1tdYf
giCDRstAFNsQD7Z05D7ngavNfvuqHiXrACQ8YTGWlcBrcBeLAaCb6ri+erPy
7I3GbCXy3rfbpErhguuzPvpwuiT+Z795OLA534uYBLc/93CdXK2PH6iF3bky
ROSZAmOtNFOiongos/QKMAJxl6X+g+dSHzi6/xhmoI4C6TOXoWBB8hJFHuEe
vLvBbF5iz/E5ERL56K91wivwibnC+440ZM1wRBqMBFXP+63doPK9PrrD5L9d
uZfKTdTtSBZ4aSsukqDpRz+UYEKXagZlV3FE1DxBLF/smFGQQ2XablVNJ44M
v1EEhYT5oZi3QfZWwMC8Cf65s5r/E1p2Cd3UAXYVZhy2rXo/bvrTT+VX85Ib
umaHskNvvp+QAACEmnqCSvdPrkYwnGaFjNDBTbux0pv607prKur/5B7x0Ujl
8u+/XJ+v6r4WYCml17exMFXBTMn3/EGkO6S/O6Cv7ul8e6X95MfzsliUHKyU
r/0PIy/TvnkxCiqH4JKny+DEi9P9t3xX1CK5eE78r1AKTfyce90oC1BlA08W
YZakgGK/btVQircNC4PNFuGCtoOw2Jdafui2ppDgh5l4K81yUmOq2t9QOLIZ
KtnPtbKxTe9HHBlbFVfT+eLc9QxeMV3r0c2Optw6YxfuIHMkqeqrnMui3XBR
N+IfJYHhtKi0bYAh/z312jwGN4/0iiHDe5DTPpIueO9fSVYqfwDlMqPwYzf0
/PY8AjvGcmmXwNjtibGEFINqO2haMnSYGew/IgIBPszQT+ppjzTgxcABFSnZ
ouguwDsJlwrV7+MnyC4imDfHtBPw4871a0tpEAdaJOva2FIgvgkHfgkhcj2Y
vrSG4+dWz3EC/lIhTB29ilId3UFDj88BHg+5JSjgqoA/35nO2LSFLy/mzPBq
hGrvDrJlERHaJKq/JuI1VyvQySuHT2JvlR6ylUY0Gwpf9d8uaxsz044c2F2L
WfI9Zzhl+ZQ/E7mK6pS39sSE8DYem7kopJ57vf7pft11C1++aViePd6kTlnt
ipJvb1EdQqyimpbM+ZtMnaT7ZWR3Z7eSE65J+WP4DUZR2W3QfUidxQK4GaP3
jKKZEuWgm8DtVsn8cgeaDqwG7b5z6XmLSdo/NPhROJqhh3Y2rG7uTs0wENiK
z2PaSGd3adFO+rcSoEWu6W4Yhp8zFxCnIEzCtp4S3LOfoQ3sejl69iEt3JQk
GrUVjVgwIYAqIilcnPpXzbDIh3cr9cf1Sntki+6HSe0flun8sVbdOPkLpVFF
ydeS630VFSjW8VLzZHRJ4iNpkuxxzF8b/bmjMD5NHjdYvf8joaPG2aOBKofQ
n+zN0d4swQBpD/8vOjpCCtq5KWLxKvKhGgSAe+I+3QszjrqKjK1kolIr25Uh
5K2Kx4Z20GSp7azuqYXJau6GagQPY7hcZUdqHvC1oOZmBerB1+5IrNQJwBt0
G6iFTDh4P9lRN91yCf+7tsQ4Xz+6hLFuOGvSU4iOl79R/6JC91sSj2nnmsJj
Ju49QNW8jMZsHNFWqqn2P/NTr1gf7X962RvISGPo6oMi4Q94pWntB0qQoZUc
4P+67+EoG2omAIJaMc5PrJEGoAANq8kK1EUveXLcAT6YBkFVY4Dm24voPO0z
pMkkFmxmpzpd6ipF6MB7c2VXDGyRV0FRkWqZ5fSoTAMjcoKmQA8mj+DvAXsE
ApzYvVdQzoboWdAT1q52a0Slvyp8RHElwhLGYw/RRR3/U7O2a7H+sXWNPJR1
jkVNrJl2JaDIHGOqkbvJsxR8ufvl6rI/4H011Djzrh/XBk6tqlWhUFdh159l
HtGCfS6h0puVK0n7bzPOV1f0fLcgvdF2qQIzC9jYUB2VOAcNQ6km/lS9WnnF
deKgrWc7y1e9wpLRfcVQbo5mkSHKEhCwx3m8l9+8bJv7GFfOObsQl4ITxn9e
zdBUVt2l1NZB+tXaWXTaIxr3eUYiPz/XQnaIOGa0N/SAD3AuV/whQGgrDwcp
jYLtfMPKalCFx4CDGW76Gc9mrgWwi0+5TOC9yGDZ6FMVxru5CfviYE5boD5R
LmtVzj1YmEyTLoCT37YyFHcLa8cJ5iBGO5NcPNu27BJc0Nx9xXibZ/r83e5D
uD4QKvBwkSbTfdAyRjlPuBeaT6ttdN2RMEZq0/9BMeUwCqcGvs9wa90nU/2X
TmadJHiKL5vbgnM8prN2CL2732VFh96viDM1jo5oWc0eaVM7bQy4vFwu+4mj
j7XJLmgMeLLea0b6WivMwBVUNi62pFs5+7FSQaF3cDtjcAR4Ne2PrqQpAzVW
Rf5F26M5cfCNN5wUXVfTz54iJZlg886bcMaXTSrSeuWbiWuxQGuUoSFUTRaC
AxjVHia1/mjCSXXK10U9jQUvslITCigLQRFbaO3SM8tiEArdxiSBFhMVQ3UG
Egs1rp6ZZfjp3+u6aex4GNeNzT+EsnRt+6BCyvjKovvZOhY7Gubz9c0C1MUD
ZELbf+7ynV96CpBflsRs0tk9Kofc7G6z5Q5P1RkabuEmvxYLNSdUO6puqmgL
N2UK4+SD1PH1T5SaQk+WBi4OPwDrXR+1crVP7Gng7ezBCxN472g4U9eWjxjJ
SDjhEssEMdlZOclyZc4jn95f+1b+3IqCmawujKNOVBnCkpRmxepHk9aWq5LL
N8lEIm1IE8VVfLWUDb8qZ0A9KQ1gBm05gv8roSodXGwADwz0xifZsYt1HZkI
BBvWkmtUxs2LtWx6fehokGGoZDqDIe8D903oC+7fHNBGQe3gGQrkMn1H3JJR
ds3sWRvv5ab8hU+d2O64v3gaZHkXHlYl3838g/C9RMLuC9ZdQO341F/8iDBC
fGQ/a+U5ONMunhQYARynizKm83QsRRLb9cZ6bMXUHFm3EkC9hYG6ss/T1x2e
my+Dc4hDmKTwqTJf5wvhkaqrOzww0dmHW2I+2z9TV5hQ5Z/DKrD/PwyA6/uZ
VszdcodkSNuYiTbSNCqAc19gtThZRboYbsvjSqaiCfQWMpbRwektGvpr8Rxj
w0YNmqgOyA1fhtGPP4MCwtgZChlr4Hk51pN5o0aOXNMVcvF4HaobqXLGKKQL
DXvBvTE/wQ1kHNRpuZ9weiwA22P1cJ61Yj91iXDy9dVnJx1y3OS6VMDNdihG
KLR8PwP1jI5gxHHDHP9sJfiV/7hefAYfjy6ylLy6ogqUllLGsjrqTPhVqT3V
CTZtyXQYgmygMSwrAqwAvOQJMDHMcsuQtwB+wOtxTA7B83TkSkbxsbkvnSey
Z7UvAGDTQ5+rwZP1oo9Ecsm4MFNSuujeFpu2kPnaKU640d6SqgcMmM5QQMeE
K/1IV22zlwmws1L88ij5Rh8hEkbMXsP0KpmhpkxeYhsXY6+s1AzPXBeleAAN
Aleos4JvfFMWUUIm7njVoa01Q5/AfVJzBHqxRYoxL6T8/ctDMQ0547rgmP32
zw2n9dxhm/LPrFEFtsdEc3xdZ62fbGs5vwAXSP1/hxv5KjVSbLniAsRjkSJN
9+zzLVtEqPRu68UrljPZ4fpNrUkt2xGhYggb9J4lTMjuKd3EGvlJBtx8Hrs1
D9swtLXZuDQH0/JPTCc+s6admqO2PcPgdCi1VWyIl83O9JuEvTm0KsyD8bIr
P9h1UA2J4yW5u02+dU9LCUZqYYnYmTcB5uwhBdDk0PIv5I1zQqwu+yz7sTb6
cNu3QuvbmEAwXR4heHcy6JD3x4DjomnHyBNK2bL4OmC1Rqb5t0jRh8j1sU4N
vLirnq30dp6pQEPq9DsY/OMl/GLLea9NSR1smWSN3xF9h0YPKlQ3zji6U0vu
OmfiI3s/pHVj9oJjwNbLDtQRAJ1sLugnrhkWg6eCquLdzbSivjiy2cUGGpii
ZoHE7eSyZc1GC1c5PI0MBPraayTiyLVU8FzJU8UTeM3OyTOs64SvAJF3R+ja
WLnjxxdezHAHNPzqEQMC1V8hLR86kooxD6tWdwXSTQ3Iq0hieLU6nWzsTIX3
PgN1fSvBjncd5AwTDKdK284wrst/y5GKhsFqcnDVF8NYHQtSg1TC8JgAWyM3
X7nBDUJ5P3u/uLRxuMi0TB4JwMsYqrjS7sOLuth3BP+6aAs4IFOXqZWl7Tjz
OJ/z/DtJsu/OjjU4NPjvu8ayFuMEViEtJ4fK3KdsPLZUmbMYM9ehxsVtISYy
+OjW6Ee7lzPNAi2jZKQEhqCEEhbPw9VqDhpGs1RINHCLeJrZypLhnwflwSn6
NGuHIiRuJkOiHbAsaE3/pfP1VUudkko+9yeW74sS2Bobdg4kN7G07QjgYFSb
wAVdeSbFxkfc4/TaWEV6wX85x4a0/XEVYtZyPVT1a/fm7K7pwV4cfj8FE+Yp
3i3D8Zm1A/Q2Fvs7PBB8IKbv8ou0WAFYvvf2RHdlngK6Hto9yJGIXLA8kvnE
Ac2PEBdayuUaWyNHbHeZ2MmjDBOp8eITTE1PjA76KqUyusMdxAVF1Out0Ozv
3sUySd2//tD/BV+CQx7wrHWBxO+f5K8S9wuQ2B3QEuuIUNvqLPvt9J5yjb/t
lxfg12J4qX95Fxelr6azmOwjDXt1RoKabOQggU502aT9M/iUU32G5zS/5Qb/
pqK/0neNbR57VM4rVo39PDLFFHUYfRSXLPrC9clJykwcpxbf+GMH7ZZ69aUB
YNlxFiEyW41YTHhNPBu1kRTbhDaPZU2gqtreUrNgqPdzbgO+YeGhbXGyyjHO
jKnstTJ8Jky8FVCAQ8KmP27mk7u+gU8H0hqVMmOoky0ZnGBFWh6QWrr0vaO2
353ALS1agTb3Kmb7DvrtSyUse+YPQNwpfVlU8aLduuC/BJBk7kep2eR18Hky
1xbwXWVmmPYa45xpY3fLIZUQ40YVyOhX9qGE1joIvx5C/CTxY2FvxrkIGFLu
UwOxcB7AbOpvXv2tZ6LgOoCcEP0BgPZ72Oqv1G/yQY8TUXPgccq/CWhuuStq
6fo0Sq7BnzUkZ9daKnL6l6Zm9cn/csUUZ1hZzJgLDAhumSbS9DUbhfFq5UNS
huBgLOhiaE/B71S6ljKcXUowYCh6NAhILbE01ZJHzGa9B4s0ktjqE2ifFv+N
HxKrmbm4UxQTQSu0H3+T5h3350YIHnDMNZVHJ+Xaf4nK7tUGWvck6bfwcV3U
JAzK27o/hSpfTDYwo4GMRbE5u0yjJcSAfqx/OWNThkA7OQtqz9i6kpj8ELxi
622vvaN0zh3njLHUBtkbbCCyeDozx1cP2sEHN5CuUlVGvRCarWo5OvyX6mne
gzUi5KHoIzLpi4WGhriRMQJbFJ5cJ0Z9CyzWPUCViyOV7VCgi+2d/poGn/P/
uhrLjtP/SlQ4kgNjnf7NVkmh+1E5KgFZzFSXEJtWBOB5kULF80WDldB8F8a7
WqCiOtCJ4FUnzPs2HgmyVkvw+s0DdD0Pd3BzP3Tjx3+fs4z4Lwh2K5CZgg4X
GJnLMvHsMJ2u4UMhmAB0UMSw4B+wcnAaLxn8uWR1p7ur4ZH1yebFZ5CoYrrw
eAWL9WIAQC3XjJXA2P2fPzUZdHLMV9XaB1zsLjTNNA3tWwijHOWZ9cLpBpLT
1slNK1PDlzRO7RHluUwaQT8K6qxC3xwVlXgKC63cYywN1DAXDpKT5rCFuWr4
SLAx2xji/jtHEW/iGge32YTyFeyj/8BOOX5NysILmYas0tn9bPD+J3+ohKEc
/eoEHYMTPXSdaKkXDbOTv0SidEdF0t60bHj1DOBm3IHKY3ykMRe5Gz56DoM=

`pragma protect end_protected
