// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
1rKRIqiv8T0MPbCLmPRxQDjklZ5isqa17E0fUlBkxkL0d3yhy6GdGaxfc7ccuLTr2G2qRnzywtmt
Wy71zQx/9vQuqB4YvNqqEXWyfHKOzDZUl+G07PWLOIpMVYEjm17xxxM6RouNY32T4spAHODD3USm
OmqJVeaIvXZdY4rcju9wBuvf5YpREXxk5WatUwlZcjSVYY2RYS+lyPE7i26jkRhivQp7DrC9WoGB
P7u0PWc9Xu8ePjQdtOdfg22L7p6xkYJdxJyDJAr2+hnrq3mqlacVE882WCGDisqeIQbqjdVft/XM
/Zn/tBgWuOorIoZENFIYsT4ZBxDHCZnTt1Qghg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 32288)
zRkipmpLcG6cLoCOD6G5LDBf+Jxg+SlII2ySh0iJcW31eY8oHUCRCAQA0811tR0YZzNYbZIYSHCD
NAeS5xTlPB3kiepVFJaUGHabhe+bQ6D662cAFfqfm8ywJX1uSheKV/eFNWGE16qAPWMDsROfOlk3
EAkJnuRU7gosfDLiNpoyzpU1rn5TwClx3oa7FBmQ0NPNDCNgy5YGQ4MrMkvmrYWE6y3yqD8JSWeE
11shri0olgwClKFTBHXeAbtinA7QSogfF065AaXMbNJfT7IBLMA89qZQN47eLJF+DIsjE/Jm8SKK
RxC3yg9oHkss89JR2B3AAzT4kC3WhLz0GWQDPGuQtlOnaXlCf3M/4hXwVTnc3CrKBDibtbHbqnpM
wByT9jo/+ZbS/GlFJ+0JbmqZosUO8Mp5HAHV1DLXLObYBT+8NDZJn8A3BLWKEmtWKAN7BNhHwQLT
3nbdLWiBiHuLPIsEOJmJlTr2JG2IRKPkVrwFF+U64usYef+1LBqbk1J39vKkLKPY/CU89a5YtIN9
3eQFiqRsiMrQ8eRCLeWn+XjQpMTfLHKJRKQ7q0xENiW+Cd/YbctLBEgQviqmpSd8orFZMjiEjZms
G7T+caZX5b71LOfOeEY8L/l+k5kanGQUEpH7sRPxokqNdq6KsNns6KhLjuf69zjiKObkl5dKyXSg
24BpuA0OFMjC26TO5RFX9J9wrq9Aw3Qap+tVSQmAV8HLjgvZ9AqPx6bGgsmfFLaODnY4d/RRGxrj
+TEIrtPjDH9P9PA64E9MUvn5F6syZfIchlFZzP7MPKvGL/Q4UEs92sJqQxMyr5EnBkuzYtY1kRTL
ZOGcDhxPsKO7Zt5h7xJCFQWoVaus5etl/kWGBKITsqDbFK0gfMBKPO36Ad+fNmFdiTJx17yvNr+D
WgVLPwO5MOsjnxKuOmXPJ4v6d75c+Ln+tNgO8DDBi6AY9PM11ck4morWDr3QYZWi+Rj0hm45WpXn
Wp+JVq59OVKMYu5D6kaJXs9XMI+sL7SEbGiFkImnRPF5ey/qziT4vzItkU4FOKF5MlmYyhOfI+V6
55yFA5wK/+wTW+QGZij5lfHI6GxI3/Ga98iIIGwj9zpnI62qaohtSNB76HJf7m7bKFoUz9pTljS1
JngC5hAXRMFf8BM82+qgJWdxZfdHZWAYLGDtneNFNCxrlGA5uSB//FNDT85UFQZFT6grE53J5nHU
9x/xrr6f53auDrfTR3+FaHzobFrP4s2cwCa6AMshM1FlP9JCF7Km4tiPcvcm7GVUCaNVj8/drPxy
mlTLmnpcktwOjqMLQXP6XPdvd8+KFzHUs2Pxd8U1OCI+BjDVWeMv5CQGuTWgW6Xm60PCcYc/OiZO
hVvME3QbVG5jERf3crFU0zSZUO5HILLUJOziHEeiCNHX6csqKt4nHkBwmfeW5njIczyV/mAMLPUy
xB1dLAv4VadHOKzxihf7Ot/wsLmidMSsGzMKyPIUqM4EuBmBW6gbUefcx/2SFpGd3n1DbrmHORDJ
DavP/UW5PhAnjRVZFTOQDIwsjg9Ay/DcMyOkUYptnv//47mx+keCVFjHaaKGhXV+MQdriMflOygO
8QVf9MoY9n4WK4E8lqcbIKj6ON3+d+LXJ86m3hIE+4THV+caytCwLLOqDYqIiBwcvCDQfX5ySmh7
09S7yEwP7gqRDYGfhAcPlCL3KY7vDsBlWh97oBZgFKWEOHRqmduavq0/8fOr5pic2TsW/0eGZnjr
+L/nQscOPuBi0/SZ3caybsKTNMt0IFuGCACgvisViEb7urPT5dvLluUCb2YNkW29B3nHu8iptZwN
xp49wlsHzI0Cl3m6QcuqzbKL493gfsiFfPPwNoreELw//ennmbBJVKMS8zXLpMjz2AE257YNo08T
M5EZ/NYUErQOar26cGL/d8yhBoaBA59uwsbVmwXKSOic+U3gVgrnofr0PWepvwe346V+4lqcfrC/
/Vp1HAsq/AapL+koNJ7I6b1anvoCh6hUn3A1DqkZlTAF2oF4halvbZjd8tUC0YPAK8yQhYxYKMAk
SH3nESM00Tp64yuT6G9XG2S0ROPv95X45nk4jHlFRsCFDVy2NXikT7yAkA5PjnieF4llgllWYuCG
H6Q9nrIPB/Fk8eHpxC0geIkXGu5/xi/yaC+KBy41Tr4MQ53IuMZUCFUNToMoWFTSOu5hcBv5SERJ
W4gn2sbjTihLpWRludR+sjvOtRYO+FjmQbIUHE1ES0PGV9njXNQ1/LBHTa2nIjAtMdugAPJvQMCz
hcoH1eUXYw6A0FdFjBEhMZhbmFC9M/jUsoKtYjBVnAA+8Jhv6L7uAakzA110avqwzHkRrukcFnz5
s65DclD8jINDK922CHGvuTC4PAzImps+GibCn5r2IbTk9MAme3i6TidDGL/SqI72nJgk20/2aaI6
89eWPjdA62kQgR3km1JsWcq+HpajBSyD4YGx3CVfqnkokIpJC0wSLaJky+TGjIA3HlyHBRpXpIun
e7A6kCWOfN4urHJTnEXEu0q5E8kxYI/rxZPVg1Ezwcy99lAWRJ8KPDd2+BQtejBQb+es7kDwcCzu
UL7WrGR5+iaffW4htzAcrebie6mB2KCTd/Luoh27/m5ih8DVtmOTwVB9Fl0JMN5mD7akIZ+VJ2BD
2DJgy1htEJ4ckt6zok580xLzc9d1Oiagmx43r1lGECdVquAnTN6xyWj4bHY1CZfYSnViqOrJvycL
DdTrO7ht1SeoOt4DpptKHd40mL/+DapLPUac4mg21cuEnZJY8/Td19Ap7iNhInrCJkbQKU8JMz1p
lHKvWAcHynauEBlWEnBzVTjBHxjDLJSZygq3X2hRNw/TZvmR5kQrTNBc0JA1kH1FsOVli1WAGgG2
HSZYPm2nZ4Lyj53REQyRFzoBgh84LEUk3R2pqnCGsK6HjBIrE2yG6Bgawsqla+2LoxqE2kH7VPvJ
qmS8vYvd5EZs3RjzOa0j+zRAefeflLXqOloVTNxAlnPa4roCXnZnLsFDmu7sUZMu+8DPxeCJ4Kkv
3kAtoi1ZgynBzqs3oDxvaXAl5rt0EV27Z4TP9IYZzmu5446XJZLrkV9gU7eBTHEg8OuVnVa/YhGC
+Vr4fnJbKDe6G6oBfv8sjc4tTljwCTKydcYE5YgzuZ5TOxo0bJ33cz+ACISx9Lp3fnp5JTqCPn2i
wWNJ54DQsGMtFts1KIUbiG51OY37DGxHrcBY3h5oa/sWICF55oPdXjzsHpDeV8GZy1LZ1pPk6DIK
TQj4Nq710G7T4WA9iqEc+dOuPDmFDau/LgPnSlKQk1X7LQN+OyYaGMibq2yAg/lFp9dWtBdATw8P
NStQIYbvqR8q1eCKuwgfG2SNNjcwxQxp04wuC1rIFESz0/IPbfhiCEJni5qvJufALoBu908aeDbC
cNcDUeWCdOxC3Xe1R8oInYTIDh1OKl0kMRNiWZfKvijER6zrLfdnsDWy7vxWSbumIsZBFC/Nc01y
+wIM14eh+TCTJsfPT2C6y1Z3lIjDZyHlCBlZ4qQfubz6hog0x+VNWttyZjsB3r/DvxTXn3z0rX9T
yDvs8mwNPLk9ckQH/pyucgBwLbuFB/mm0LgUKweJiNQMPO8uI6tghXlXBBPXsyVPjki861nXNVmo
EKGJajlJINJ2tr6HdIrfh0yb4KKCnhcETTE30CqAvYF3Xu1U9duK+d1w0hPxRab0EQvUFiATEAra
yBwffeJTSJ7iuvHFnekAoadRBQfwenahb0MkXviscF4F2zttkVz1YlF8hqRZRjNToF9aZg11KKTb
jOoOT9CVWS/ZRBx8WMzOrQCNFqEyJpYix1YXS04EghUeBwgfzxk87W6XTC1d4K2VFpcm4MUqT4B8
wC8NvHAbAQUlxyce8L6xYrPYrwobwFfz0Fdl1i4ylXZKc8zTuLRaZyuUIGkyBodPF1MW4OUIfJ+x
32rZD5+4YjunbgqatR1mcw1HvPBqcudy5avmnDn/9HnAYdiVDeYIMEPZZdDFNIA44EkPT74ATXkc
uIPoL5NtU4nhHT+M9igsiNfEwXqrSyvuetosEXMEqTEno4f6b88LGiDWqkw2INR75F1SBAF5gH+W
ziEMUviQ2fPiGOl6OF69Lhr7a+xrh5ohR8N4X9dPvWWWnka/xjVp1UM7QpUTGpYJgcibEu/wx1bF
YcFJsWA3mgOIkpP5r5SHskEIsvzQaRBUleT8iT8XmcIAKH5h4tclQ0hMEPynBVOp6vC03F5wuq7E
CYB0Pv3rnEWlsrK/JYWkHE5itMGf/c++7M3VBnpMXk0KK3iA+sbbpH33rkcX8lyYsp9tWW0xUCEH
JvxuSNiOmt5Jx8aSyho5miEJa6EnSosWr23pK8nv436bt6/s2RhOuW7TBkuh0OVgzXqgllhu8EuK
tgFTP0QQ8p0+ryKojZWFLHnfHceEjaHk5Nza1p6G+pLVmX7RxtX44l5bbsVOBviGLIq/drPvE9cu
NDtJ43CRAU4i8W7SRoNhNl2mrpJ7Np2/bS78MpLa0UnUDB7XiuE2Q2sS1XaGJ5yoaPj+sKcSSJev
Vx6ToKTBUx6gJmBXk96sNupofiI2nfOmXowcB8jxgMib9QNqNcKsl2GGIeM6ZDBUNdjmK5iaPCi2
S65l6Cm/LTDjAvieSU69KFCO4xWjJEk2ZMkD55ozZ1r6B1F6XBjOZZG2y4LQwipk1HN1dIkIaVQx
mLt1O4wEMCHL8TmvYoho9VVZSpmagaclKRKSIAuMsJ29alkdBxncu+aDVE5JrtcTJV6g4Kkp0nuG
nQUBmHfz78DZ3qCF+YcmBf/GYN4JndhFR+U+UOBiBI5rb6R9v00gbLuT3unTqvJhyW+xFCpf6p2K
19X+2Oa+/9kceXO/MvcnIvW9dmvXY5oXYw4a/2Qf/daJkQsCLX7Jvvn8aMp8iRwc+BMR/LN9COI8
CLz3qw80webqs51iVzf4FRJOn3uQUmGSpIWvZ+ByHNDWO1+yL8uUcm4HSE2VJQn42uWen+BsIHpi
GoBPO0VepaWLCBRe4jWToOwA0f0xlpjqPWudMXphtQ+STgBmcdY1PQ1PBG0ztugxfZKLvC+f1UYP
WIxPpgvT8CC0c0/lypcRqSWgmx2SpQJtGCDXGrWLM/C2WOLKODE1VApKdbzgWMG2RUCmWdxV9aja
XugZ/a3Nq4pLGLVFhZHkpx1SwMgwiKstaTin5PmWpZpe8EW8DJe0KSk9iPfYb1DOTJXzBjUcCg2H
YXuE/GN7KUaFUGVyQPqEXVC/vzKdnlivpEfW0+rY3BhNx7U1+NglPaa7aRYOtkR47V7PzVjuKR9i
YjFzjdn5C3fAubZNE+1zM0sufsuWRIthBZsAermmuLNJvNm720DMsfmCDiLsWjQeE7cggpx/C7nH
D1yYKGSjkd6gdu1rrXctpqNpQYoHDak+LgyTFXy0R93Hc9XAp3+a+Ue3f6o7YnO3/KVP1tbGAhKc
iVR48ne+7Oif9DfYivfdvW8Z56aGa8neVtJxC9R7PYLhBrQm8AH3dbOvEyGoifZMujcXCmo8T+zI
O1n+UHEhCAjfJ48GPfu9pz2T+AkHmORRtzzlkTvelGHMXgBaUWZFXvIwvn4kWgzy7fw5iUxFemvi
7Or+vps3sS46MMnQ0EzRQS6HYdWzcXg3//9hibpM7MNNksJSwACAOtkGetKwI9XDE1zPVLjFeFfr
u2xCvod4ZJ+iJM/RBIKexSjfQAjqsG9UADGa8RENE+pPXRShk/0z0FcaLtm9KDuFADrcYzwGXTz2
Jl2TEr7cQL/5tc6lAEdt1efY9tWAwtEgz1lWIVCZP3NF2eW6tqkMM/Pr1oULJB8l9YloCYrInbW9
3hChhj7c0cFUqq/3yBg/TQITpsuoPFke4qlavljk7qNf/CCOPjhqT3uVGgmP+k3Ugi28sYQJV6uN
/tWMeU+kgn549NbTBeZ0oV+3BtGgDY0fnZ3Z9k//uRXrFG0oR6YUZBY890QrR5l7SUypF5kvS40W
5Ukw9uFZAAjq9ocq2UiHenkVnIKv28DENa2bBcsId2KPulNIHcBOeExYb8xdzmlHbhfHmiB13rdo
4KuDfEOq+OSP6moJMeS7unI0j5gwMPpEtbMEi0IGfYlnMpdBhlpMqdXFcsctu99BxD6lsV5Hb5du
aUZpArw1g9SqBm41/G13KOSuyzJ+8J7a2jxOeo+91/Mpvm4/KpgdlYsmRFIFw2+kwJ/CzToFM/Ty
kYKMH3DfDBExFo7JYvvQrwlXDIfQQLiDv4q2+dtrLpCRDiLM+M9AzEbD2pkyc3BEPKAKDGs0Z9Xl
xm1uVJ8blymf07YACLRzgtD1HIaRLgTVni7MvF8ewPePRzFRifO67kY4UN/IwSeQCvNyHy+zU1pM
TlOwuh4PpNYtqPWNh4eldgBP2+3IA2dpUttmNQZvD+vMKUnn6Y0+ADQ7SLOCw+HpZ7dqyZvJiYjK
HaDmHG7CJA9GZ302Fippdp1JZcM3xCwhKT+5B4p3d1kuxJfYEWlB9stoSpGY/zVTcTxkqHFld1SR
VbWDjIlsVkxYjnohajZtu/OjOmtDg/3mSalVh+5wqZC9/DnVMvwhngjpuEEsog5WfoT6BDcc4meI
sKz37nu015AS94ENo7v5nPVEy7kKjmX179BJ2sxHRqmKwbQpAN54bFFX/VSkswwu7+Cbgfzl4hRz
oO9ALwDcFzhasvEshvemUr0q7CFMAJ08PhLWa7ZrvDpOd6dGdlH6Vgh4hMIp/hM7RgkxlsEvnV/e
gkGEf/a5IBtyyruF8H57yWWH4saKgwEB+RSurfRp5mOY7vgAteTtZ4TeWHusbmXbogduw1cZPn1R
bM9Q844gERWIiJuBypanIX9/HELuIkQi/+XH3HouFoB4281Hobt8fTBDBhml8hDbs1CgevVTMsEY
74E0d35wuKsBOnWKdIEMQB/X0KdmgkwKdnJqY3Bn95mkPDSkxlJOSTC2o+3MyRTcqGl1MzEoco1x
VOT9aznkqqq+hM9xjG0dF0HJekgIAOwIKo/Mcmx1/DvauQk0v4tNABSOdixXKKkH4zUhkMeTvVzL
U4L3YCSWvB7eQoY+Vu9bt/w/657X3GsxbelMZZKXmxnljYxjhNhjzouxJOeRCwQpbJpTOkJATidj
rDrkngFkxVnzfq7J5rh/aSBNY7z0lbIg0aXk2Hvnqoi/jccNcyOzy89Y5BkDkjFqy1p9KgasUgEF
dj2b6vvYd/3HEUJ0pe9+ssGdsAcDj8PB+F/VHIi5oO/52OmvU+zDCEq/k579txhbydmB3yc8FSjE
jda1MWPMG56juGEIqdKnIjckV5GpiEc86pFSAXuVbPri4MqUjhSV5zKoYrmNMs9bB5XaSrIGFc0w
sTAhuHk7Pee0HQrlICD2x20QnrvKY9qnAVtM9pw0iyf/coZc3jSWYPPGjkI4FMa9/ML0koolnkt0
bf7aB2hXQSsVmEV2l1tQehKXCGDAdohjj4eJ9D8mqswPL9fbXrZLRJsODcbuw7qfd/RuINRk7QFC
hdxPOITMpUvkDzls45yRNa8ExZTVChxpjfIP11QLGakDK2bGMEMAR5y75X3eo12y8JGI84PmBCnc
DeqOVFXhK+MIJmHyWn/zYtKEUz8MZR4HvGpU5zUiJXL7wPM1TuJ2mzsdL+YEWkqNUYNkmS13WY6H
I2T2pdgT3zJ1Jwr7edvts6PNsQblOb1BP6Lcw16Aeeq9g/HrRCK+5E0FE4DlKjNZv2qqWNulPTSd
EJFVaogtRay0qEMnd+7pubWv70Ub/bEr9NHTkuik/9EpGOwyBdSSmb/H+4DVlbqNt10d3WYnDKOK
9+hUI3z+X0yq8eq2AWysfr42g0coU45l7t1L1c+FUKSaxMv8pEdfzlidLn+2KQ+M7elNu0THiCxm
R594/ia3NOEstQOXLwf2dIFHUkql85UsajOnMsnw4VqLb6hs8+4LRKy08AbV952msBSYXSsuNjE1
F2wNUO9b2SOngHBJ0SoiV0So+yEIEAMNXvJItt4ZQwCdWNEdifNAEvk3WC2uPP5INthZwv8aChNY
VT1DIeKR1sf2aqpvTqguVSNhzT27+N9qF6XSFTnMVIrEk/RYhozYXJPy8+fLj+dkmPEF3Hm2CSty
YCyQTxMYP5+qk/QfMfDpi4eGhkq0gzSGnHYXtI3E8/2mLY0TA9ztzaLbzIkVU/T93q6RVXxhEKEC
iSs6jMHSkvmqqtFSlIjm+hJ6iN/nLwdGzuOaJsJ4xkohGnGlAesBtOv/zQCPw797fc4XLSm927d3
46PfLH9w13t9oHBVT377qkfKwxNSAE8pTYO+cBcFm0vy3V1l37XZSetcXN+jqI2kCGZrjkAYrPU1
7fCVAkKwv+TqUwtN8SevbVu7++AYFyDnmTUHlXfXlKpuXo7Tq1zoR8ng8payiyGE/cAIOjKarj0z
xVo5sFLaqi8bWsEsFyb3u3GTFWx51j/1sBYnyhULhLBZun9lbVHqr/vP1z+NNk+gPjTV5/usFs+/
+GA2K+ksd7QNY7m7PV98S6uFdSXxpA/bLeOiPIbfHNe2emwgb0m5XtdyDCoUrZaR7N+peYUDPy6B
XgFT0vBXZP1Oz32hu6x4pFNV33ytEPImLPlHh0gjflPyYMIk89xPy5w5hIYA5+kSC88ielWvB9K5
T5iPhIqkrkAaylAKLDQJlq+XqTaYzFz0Hw+y4x61xcwYyZo/JMjFpF7LGdmIvlAy6wnkXeiB3bst
nFiDCx9EeMMDpBiWXDrmi4dE8g7OvXIZNZDGUaGuLS2Ese1geW0hN5h4ddQlShbtsQpKjW+93NhS
tqU15yugYQmFJic0i+3rvh0WfFQGnArIKcCVDqcnpOngRhGbCassy/xuI1xwaclKeErV4HbMY2Bn
oCxN06M4hdf40EqFJY/bSjitec/I8EDVKtwb0+PcRk32E8tSf2SFoxyNF1+zpUsRPZb8fXRgYLWI
IaUwQ8MZ8fZcBNjSToP3vzEa+30T71S5S4RkZbkoXYwzN4sh150upHCVQjAsEi0B2qGppCaKWyqt
FH1seqNH2pfXgnQj1vX/fdJWE1zuuCgpWs1yzNDeDVq7fMP0hODnbvluRx2trXJ8ubDsXM+RpBEM
DT4JJ3BNj67QKc+v08Xy32tspZFQba/GC/3CPmjakIFdgdGcXRHxPXnjDH++S152PecsPEsicnua
dL85su88DTLgJlqDxgdZNTe5nyGKf2I/a3Z2qSyQ5CMcq4Kzi2TFfLret9CkOvRcCmJqN7rlD8dT
p5oHqh4r8AH4YfHSaeuNPzVVEI9tCDdRp5m1yCbWYSoDDpJJVjtNdXAN/ui4RqOcFXciMMWZ4tW1
79bvL5N/xEY1KCU4iakulXlKLN4ILsGmsG8bcqEZCsBhq1s2le6vJAdnIuFPDPLxofcCRvzrjKLp
w+SPGo8SlcMi62llIgCKsxwGvh6yg0ePeT8nyZtQK5ogBLYpl410bWwzwg/wa8pDeJYl4K8N+hH/
sCJY9AqWnOxgY+O7Nc2zozdftUMUEoL4ODjSxIOoLcg8KrAvryQLWmrU+dxP7H1QrYcBHduuU/Fk
OzmM066Zd5+Kajs7rZI3RzPFCGJ7gsaNRVLlWt4myKErU3A9uatrUn1MIUl6QQhBI/eT/yYiEHa8
USIdTIdY+12pbiog60Izz7xpI58FPh4GrgqF5/IVxrp9hm3Pky22ix3OJ+QDpFoS7Efg8RZMfnpP
IURzdVgi8lpt8ZKlqxskYEjnxFd8QUxE/NBkpDmlGtm0Hq3AZ0saT+jRvN8d7bZ+XA9rsuOOFEAT
scpUqu2yAlu0CIwcrJ0dZ9B222oFWP8hXK3uVsmAahncYwSx1PEwoKoml7VxO5/xHEUniQKV7144
heuW8WGaPmhKU21nQBSmoplL3ztzEocjaV94zu720zc3cguXxUorKo1q6z9q2CbZ9KsipEjK+Zqb
US+UwZH434FgI1H3lFTa3rZqUFcsQp+Yi/N4gTnX3D3J9e28MAVq4NazoDj/wtLnqdPX4oFN16w2
nAru+RTny9O9yPwXZwd0Ft4QrmSHAwI4Bi26zax/FbQs9ceEg+O7SmkoOlOdOAzLEIMiv0OPQxeJ
5U1DpHL+5c3Ni6Xtwvq87XnXmjzrJjVIQdtmIzL/jPv4/OiUQAhPSZYZjrF1jkfz8TPSyW28PSOB
6sgnDGTqFDG+BkMJGXzFWAz2E1fQi6xME5aIkaXAcF7QfY312xDmJuf0DqBkza5HPnWVDsZ79Dzh
TjPxIbZGmfZCdpnWvXISwAN7r9HV8EqazA8xmyuS3ZP27zx+m9p2VorhtpMvxkOJJVVppCTWHus8
6Ine36WtOJ//8m1Im5bfVBSUHlsxNWQljLX0WpCIZtuiJxLcOcRlPAaI5jZQCu/XKN0wGE9X5OTX
FdpcG0Dk737yvRGsSxfjV28TosG8x+VGLYAMX3uE86Aw7E2yEI1ODp8uZI9kpmVpn5v+t3Hb1H3o
DNszELYgAXhfCKN4sxiE+oUFn9jLSpdD9hgDHFSZHFVk47ajgQHL8Zmy24b2GTSo4HXzjSCO85S9
5/mSiV475wSwUfaANSbIkndrK0Dbq185BxMuTPdiZUVFIayiTjijBW6w3QvvhBo4PsrMhyILe9Kz
5/FpHLAWKGIkHfJ5RU8SM9hCSJ6lIeMfIDe+O8F0EWFO/jwd/g40BbySyquIJjg4dGRAM/QOcpDQ
KFLDZe6p2si/9TH7yOwvvkAl70QUmxkltfk2v0xFnhTzCSV9vKLDpM1E11MJ0jvoNUFQIiO83pOB
AbuRFJRBpViw8QDJP1miBKt9D2e8QP4tiaSua+kEP2EKn0+FjhHtZiV30Ka8OAkY/p7i3aljBe9R
mUEPMr0QFLc9mbjfSvZRfNi/BFcGC0+xIRjWYB1q5fOE6NCOam3eKkAmm1wHvUbppiflh2+3mYjt
ZTA+zhytolOoZ3NC3jrCDC0VooSfe9z08oNuYhG1CuOTXq+c9AEw8mXAzGVdKTYRITilvH5o8kUX
gSNcg6C/IcNPK9HZ5SFnyJvqwWAwK2qcSnmH25BcFm/t+XG1Nw4c63xVwfggioRCUS6y200OK2Tz
D3k2eRFpAu/6YCjtrUNdDU5/+Ui1BrLftRntp7MfTZ4nBbkgOAqwRIr70qOK7+InJH9YOwFUnAWq
gXuUWJfT/q16IMDkOYctYiLGxO3Hh3guazU7BTOGPB+yBPM+EmIB49UoSZDwGh2cdOph/0uQ4aBK
d1eDgSy8gn4/tFGlao5r1U9xPIET+pZAx73Z8cE2CoPdcbdVrXvmHMMt6mLJVgCuJcpY4P5KiCqr
6ZEQu2lXDMVvj1lDe2ZN/HZCQleUOOO+OrQu8E7qtWxIBcE+7IaDl17j5z+uqaoMs517T0bO8O3G
33c+yYIhWI76KSMTnxKwxMqVvVyh3VVRFoPbNrnnzfhErHDKmWwdJXGLtFdxS1txSvB3n9d2pSkH
Vq/eEOOo6ut/l8BhBjfYv3mxy/lzLebCx0za1KtTj5y7sHFNGjRNuj6oTQo44smSW2Eu7tgBwJt2
LXE6qzOvd4MXpJrbCbJ+v0QUTZfzBdUiMRwRjt7jUv4quq21njuNooLz8ATNG5c5AkzHWQASWQ69
R/LckOOvo6xT8cuScMrEeRBMMg7iOrz8E+tuGESpGuo1TUzjsTU0Rdj2hXKG1gxInO0J/fjQUseP
n5XZ5DDJWvdw8tydzBJCbLFETe1HI+3+LMIlMMcbVzsdol68ihRR1WCx4iiwx+aKxYDhqEK8XNYR
u8wA6wrzS0g0Pf/2SkZHOT51QeO3dAJJSfTUzNHQ+Z2AOntHn1ffosonbr0VT5YiC8WI/v5JURdT
2G93QDwFJ5gcyqKHbEB4qDRnzEB58RrKFs/KMIzVVuA9f3zeRV4lq62cuL6vq+K4y/WaZslgJ3PM
FavIi4fcV2bNsWx+WCk7xschEmrCHT27ekuPz+rbpwcppO6pAcqSYpAdwT5rwiC6vq5fTTKXR4LR
SO9OrJCEtLdDeQ7vO22ZLZTJ9ydH614MLWx1Rwgk3iJMylqZ1NvtlwZUV7BuGecQa9+z5scjBMOZ
zT6K1CrCKNHGD3Uzzu+lL6Em+Vik1if0P6A4n/8BKQKBr/6Eat6VmTn8vtZf2Q3HEIYxPXsdPYj7
d/87W2yp7sSo16WCQvacohXkIfhkvHkDcwq8cQZYCi7cxR70NqjQQyt6WVQVTYfljpwAAiL22KSQ
P/CTUobFhLJbArCWUHHETFSzQ6LNgK5LY/ixqbMVhRebC8tCCglXDckYcGcD37mkkygrD1iy3fV4
BZQy6MEgtLcnHiYrL1ggzN8BUdJ97liqx8tUdCA64lQHDCF41mExHigUuxsNJOySKDw9CjctXSDi
c0cwH9o4y9viKxHl3ayTKocO7dnQKNNeifC9aF7g/a0d61CbBdoACa3/y2OndGuc12+nuiLSzPrI
sbBczTZ7u6mF5nI21pc2V5Lltq/J7j3vH39J1nlJcyMaAC8qEev48wsudJnaRKvZaqxcQVzVIEUB
5L8+RnGiz2aV4EMwAP5bAFCewfiNdaMNdHF0vJJpX7Vq9OWjDILTkdH5MhWZX33D0EqdLznPp9dW
Xn12kZHqEE33c6sc6nDK7asWq/s8RlrprSzgIJq9rQHwYCkMTQty81/J3Amh5YSq+lUFcjHFtwHh
GFB9zd6JVenQvmE787fBUF7JvDe0ymE9qytebJo8XMsUjV1SJIRMbpY8hPNNQ+2ziFhChDZQRIoC
7BifnhReT6VROHuO4umEXcgUxVpGw3qipxsrjiTDYZ0FdMI46PMpZaQCE2VnPD9TpkMP/EbhbYnY
NQZ/VyvePXzE2hZXPktaFIBbHHl2SiNAmG++OmZN71HsGFE/AWZ7Nr3MlPKfGXn+34vg7LFkYD7r
TqL8lE8Kid51znY/fNW13PUiNmyjXgPo6OzZihyQMQls7+ni/DXcvOgpZTZtmneyyuKccf5dLMtl
IqGfjxLwcLRCg+/HLpBcaPnQjWsAsWsgFCCgCjaceWObPr6BW+tmuGTpLI5PPnGCW0lKr5ZToc+/
mt+JJd0DFXFzFMpK1lfdasYPnwkkquOQR7EH5B4J4mqKmxK3zPgLtVQLt6a6KQEQNPoJuMxl9Qzf
+sa/G84TWF7wIisNdYa5Pnc1+lnmYMpj6jlQdIqQxxRRfvKIYC5v16WFmIe43yAG+YpJ3NjMterv
31VvJHYadLm2AVVTgp2/TDdOmFcBJrJ6oDWjcPQJMmVQIRdMfARr/wtnyt4Cfni2KaqZ+tS9gC9+
yqI0Bw/hJquKnwapSnu4qbeapu+X4ylPopYHTpLHtmHwL09IWN1GYTnn325nOk9NaVaWOr33m9hR
qdZAC7EEKAlL2IoXBEs61kkZaUDo6uGqqNazHsSD+4yf2GLv+pKYr7S6RdlJnru5+h+pna8/zgGi
abXoabtkiBq3W00DIokJldUngqfGj0LiZbsMG+8ULa2gCDLIMJjKTBrvnKYOr3wiFLSnGGQaadcX
pUGk32T893jHfyvZTEuTfo9YNlKxMVh6vwT6GczFu/kycZAn2047OfTau0RbXbrIZK0lEpWowkPQ
faNN/2ExgdaOTiQlP1JwFAe90oxA5qlTkag82ox9UClANOxVgfwFHDZterHwq7eA7feaiSYQvseP
TZfwtlOhdAvgIS5XK18xg8aQZmeqpqrTljsG3xzaIUWEAOGlc0EzRO0qOy1f+9Hhutz8KCfayjpy
d6oQrQyy48z2dUJc8YL8hXQ0l1z7tpHjEQYcxNW649TH5b0RjIGiIKcM72F4YVOepzKoPrkqc1s7
Mrm29DQHkLJmkNASIGBFjxGCraa+biQcxUUQZdXrFfjkR5Fn7Rnw4igE6864ofvIiaBh9N7yIBmK
Zogw/VfQlRCn2+OF3rs5PO1/m7W3KK95Ly8GifTlyA3wBHyxQ8SnEhM9yI74oXewAesC5pn5lwUw
9uje7vfEVpzzagCtt4kSKaksJx4QQF+7L7fraumFv3cyPSfm2V8MgWeaf/fl3Edf7A/Yq3rHNRbl
WFj7nHNj7fwH8e4HVY8Swh7nD0lKP6jI6F27blfXE73zNoUfz+FPyqNPY4ygouLtPi8+eCy+eQGB
NoM+SLLspz/e7wyL6NOFr9Nb/0SKq7kgecEM9WGpY0FJ/ozjw6zlBK5sm14T8VnSaX3idUyQxDYu
2qg7YiS+pchSV1WXWyQypPxVXmDkkPihn7XYhCvfGVlPGMGR/39xvrk1cW4f6q9jK+ejy1QFCwNd
o7U9qesTbZOsTFGHlXT/oCYzlRdw0jd7lPAOa96Om+wgVQVeKq6/iwr9DzdoWnGmq0oGE8xlMCVk
2+U9bXQYVslslPSdJkV4NdUlGt3txii16cY05xHWktsXLsGxw0SSkb+PF2hdVnaE0T/RQWua1Ki/
fvjOIlYk5VvKi2ZceSvmU4+CM7ql58mP/3yaVYfj3QseoudnmgQYX02+eBxETMw87AdYgdkEHbKu
+RKrsfOzP0ToD6dL4W6QNPnXBBZgqsWVsFBdf+7ZckyV4dyLHtoFnQFUQSBjyyMAfKg9F8PkXOmy
ZNEIvXslpHqw88FIrUE5nzT/H2lvDPKR2jQSEZ4UE9BqwGX50bBvDSBgyvIqTVsc27eax1hZfBMI
WNR+rUhAWniJAf6RDgu3xfn6Trjvt4QUr0mIRdfDtApxndvDki8wEchddjT4jJZwsdjJ3ZuljX0u
T5E+J0PttKcMh1crtDGJUyy/RhKVqUfqyNWBJDeNZDf0pXJYKV2sZWr3t+FE1KH/FRTAJ6Ry+P6o
QuNlIbi6qQo0u06QlpKHqaq2c21CjxSOAQ72A/HKqyegG8EWb9F7XhlNW48mHwYXpeoAJFjqNiua
OgHKxiHL/HzsB3OIbnwRD9LuA4nbrAy3ohxhk+0JecCWrI0oGmnfZ+Yqb0MxqdbqhqqKYx6NJIW9
3ileMLuiCfHqBA7Ve4TtpJW3ApphcqlEKi8raveSS9tgoyhZAjRHiypLNxj0jHPbi1GQW6jhJCp4
L1dSt4203TGBZAI+TfwAaWFX1a/vUhAHXbZf3Q3gmtwoS8wFDjG/8GJTIem8i8/fFWk2TySW21qI
FAPYB21xmGqL+FGQ6sb0l4AtQOF2jbJoOQuOHdtBJKTQpX4Nk+x11KCT7qfK/DCOWuAe1KLLeE1i
dg3ct8jE8Powr4fCgk+GEqzDSA4NnsCQj8e7ILBu3nrgOiJ9TIcwaNKNU+WVFJCLIOe+RwbuLgN/
7uFC92TL68zXAbXT2bOQjPWjogVF6vXPnW1MofIyPEyswiWWq2WejVrRmeaSAywnWdzywMIlCn4o
GJaTJDUYy+vFtIiRc9foeWPametDqtek9jlOjIp3wK8V1qHyteS2pnz17yqlqP+82ZsL/+pPeTZW
PbSIRluUYSTRb+Q5ECod92ZpTI6uNN0Z6sM0FOWwL5SiUofJYR2ADMkxHrLzhVqt90Jw7PoEFWXC
9+UbJo2YUO/r6xo7vYHgdBY4uZGagRe2tYCnqFjLaXsv/7KF3/YyTZS7cb1L1Swc9PqMPDu0YieR
JnPmGhZVwNS/vVmkIcwiixvGYK1O81rWE2J9HOqeTKmhtvbdNjyOC+6FHH5Dk8r7iQY5yNoZ40MQ
3NbEo9fA3aI53S0W1XQSRPCShiLiyKISz5s5QkOV/xlhEE9Zmg8sRYa2HgB+Zm4SLf/aX6DUymbb
4ZyL04aWWSmaLqaa384nqeKNcT/7gbe7Ac4St8F+A/yWMtffUnDyV560xyESrNGYOufpghT1rxCd
S9Y/teYbpZmkrm0/efX/tPly+psgPGJSi0PYqQ2WO7OxOHpoCDEdxzgkJxKwhtQ56E6CVRLIJXT2
OK/7vNDVbqqKZCa7VGKAwZ8dQNEQZaHKursITF/Ewya4BAqfnTDlHcOhMkzcKvwhMLZGh6imb14Y
fRl9bB1AMUreCPttsvh/aKVN7KCTze56kBP2RAZGoG7oFYfCJ+fvfOS2HMrPHey14dlCIJIBDb/d
u8vKyuV6TmzN021RXpkTs8QzzO0rlNhynbYXXs1g9zBTgcV22dhDRR17gXInccaUPALxF8mSD0ay
TSiuth4YfycTBum1BJ7tOgU665FkajmzPG2LwZfRTdC6P53qewC9Vdy9S8YNCe8zfL7udDstsFgH
X1zFpTU/wF1LuuJ1vf71FNDMJ6Fp9TuuiWXKsNZqmlw/2a1DBFUvJlWiZq+PhvKFlIkjOVky1DgY
P5GOGQxDixm8oINpMe/X1lqF+aYfdL9h4YryfTgKMFgUJ01UzjSIyEK+5Z1Jn49UNC+Ti1mp0gdS
aRW0LDauogBYwbevrDQgMWSk5aHAXvFcSYE8dRiOxLHhVr2XG8h4zPFlMIIevPllgn8Qla8FXwQA
JfAYw1/RX3eO6C72hBCmUS8uF82giSlDU+/1/Z5eqH9mV0UlsQoq3bi0vLMwuQ1B5Ruz33V6UpQi
PEgaEqhTaRR25OuSWm4xYFG7KqvYEUWGXR2JKHTYCr1I4h5BBFCoXdKHynR+iLLgNioU9ZGoZi81
x5bcjZlz4gyarIN4m/1gcRRMS8IaNf9mFCFIpHbQbzdDRvEr9R6HVg87EUJcuvv9xAanL5n+aPGV
yw+XPSCmfE1Rbw5DFO2WlaVmP2WLko/YsvsViHyEoMrh73QUksjvmbyXfQ3Gv4pHyhwPZ+LabnQ3
74jtbQcq2o/0W3TYPP5yjynY0ZuaLYuiTyWIy9GoQd5SsFqvM5LbSJUIjM5CCi5aHFSp6SKpkEYZ
oxE78lixBKgHOa51dbY3HQhjUSEZIgY2BnNLdxjpgDmq4SxmJPcT5rUJ1JauH3tU6SZPsWj0vL+e
YYqX+DQQiogwY2RtPHe2+0+rpCrc530gsTOqIS0IvPoFkiVVBEA3ZW5p3dZoUUeviG3+ZgeQYjuC
OYCnqbtL8riko8GvQFmYcCrdDKW7wJ/ypwY8dgc+SQkenqRf6FFkAQ5fsp52AFlzzj3JRVjrirPJ
teSzWtoIjWAdqjLyC4HMXu/fdZYgoVtpRw3i8Dvwj+cGRC4wA9PXge9j4JxSayiLcRiicb2wK8fk
WEUUjMeS5Hfjjn+bZm2W6Sf+Zkeg6DA4bURDQ1E8zPUDhOOd9wh7cpY0QVIUkEnq11Dq9zcPgtfN
EtuYf0coIbaQaEs3CHeRxzK6te8JoD7SojrbS76PgfV1fatlOMkEAuhzE035EBXQLwZx5SAnaHT/
x2vLkqgb+pRhRjcRMQWhY7yJRXC7iZpXKm9faBv+2z4g7FDtv9HdkXoWxfYL0Fe1xAR7+iDspl7R
F4+fSSu4dSH6bY7s+Bgb+VuguSjhHPCrrA9fSR4TCtj/7G/0G37ZGUolQYAXJ4QlqjXD5pK/05/X
s8jUJ9ZIr9co72jN57UlGIEkIz8QM7+AP0GJPrUV03OP+ZOeY+9K1s98aZz+cs6fNRuADPxlRsgO
XBFfP3H9f2rPNpPlQjhLIlx+mzXyd3TJDQ7wyduaxdUKO/3VN0mVYOZ9QSeFTwQvv+ZAaU+pALK4
or8PTMvITTMnjHGoERmPEWkGUrfqztuSWE90sTEVP9me5GF9zqnMqD4qIHNkrnjfJR37YPjX5Dc0
obmjB5Q804Z38HOVInJyPZ6rke6EDHlj5xREnv+/8zbeT6wOqj8ekZCE1D0nMU6gDY4GPcXb9h3P
0pLbcPw/FXS/a28bPWb6i91yTRZEJLoGMdrC0AxHKshXLQmQGCfJQker9xANKlMwBeDC0Eq9pFxJ
eNRxPGEZmaJcFP5G5cwwbIWqKiI7LsAhPXgiDq9/MMhIAOQMgTwYA9s8WWD8uMH8pHjapsO1a0ln
ZUR7SMKSmg4LUNb0AvRDtlpNgufJA3yKaSpqdvbDO3QA9ABbC6B2s7VEZLWEBwjDYYA5sXtkmnmL
hCyupMD9Rz5+dnp5xFthq7EIhx+mbVULHaijsTT15RHS5xMaxITexP3tx4OafQoK8Q5fzW2McEtJ
A6Zr2o7fjQW9BveSEpPzkpFiJin4YQfD0aE4HFty8cotdcmt94Q5j6493crx/IQnO72tSuTmwb+z
rAzX4ZmjAgI1bHVf3TysXry1ZJJMxENHXs6mZYl6wCy77UP6IP123d3SyTabRfsCw/K1e7IcYDkK
BBDJMHycWlruC16dnuWi9Gq8FxFNomxYxJtc1u+IDRFJxNzsAUAZhnklLFlNJh7hx6vIm993UaI/
MREU3meD5Q77iSAVbSHgXriGHZDKWHQ7Ny5ljeyLElHNMBbOU4NDljhjxBPC85HUJbOcRFpNeGhZ
qzc1Y/r9XUegRIp+7QWsFGPNEiZhHzPYWz87uJA0DsA51gJ9+MC9lpyoTcHxHiUxFsJMTYrySu+f
zbjMSve72R0fQrawBF+wq1B4O7rFoiI4D6ZeZPJeq0Lu9IqTsCS4UmvxaAY/uQ6asZb9xqt04fRY
db+vv1Zpt32iNMw9B+MCwiwcugxz4C0sezCgaOifUZnSbzEo7JvTB9cfqRqx4NInivU2jqEa3b0F
xLYUskzclMcjb1DheYdvm2cR11lRwQDHnSxNxMWaXpw6wSZoL7nZxOXlcbrHK0RgVTAPdZX8ih0S
3QSNdWnPbeWfik40UoOk0wRJPI2TgIHheSIabrN/hDwnMMOXW0L1pRC9cmPFRlWZalUjtVTuz87A
ST+AdB7leYT8usw7krs+5hBdFyaRoY+vEPzDt2XGnMsWvnhLpTqkrnqwwiCFD6Atwz8sNqmK0RJV
ELcxiZwEJ8pkUnodUdNRgzzLxEFZ+ToUkuqKz0lzvk4tJAYvp5FBcSb2k/YPDu1rlMjTbH7QBYSQ
wayhoa1bZB2lro+lGP4qTZzTeyz+4VCY7k3HS6hmTHzpokC4sIlFaCio3gBH2jQkYg9jz7yW6hp2
A03MAY8WCBg+ohQzxeWEdYNXsel3gE8GmaNG3fv/olg1MGFoYeYLdCOCSSpXl6YEIeO0py4K5EG5
rqrKiz48uFPiBHiCKHBQ9R06hC45/oYX6drRdsmfgSE/DwNOlzz+67+GaYjpcSZoee2MUlgLs+hx
yvi1R/oV8gUU4TizW2Ijz75qq7zBhZttsW93AJPPrlU7gBhFjmfmswoYB569R1YaNxj6XbTZXHaD
yOpoa7h63K9Uw7XuXmofpN2hlNTCp1F3pwOt5R+b6xSVLWdV11pzaHRc/M/bRKiNnwN4jLxrX98U
i/2E3YXYqNw1dyezuv1oYPfu01Tf4X9NeLFl9q4M2DZw08N2x5X3ieVwQ+gAorGRkhfhOz7lbLGx
6eNRy+NaJFKxKIr1BB6Ji2Z7kSKot8Md36Uuy+RHifLE8bVgqGnrEXnm1hBRSV1/63iX9V+t0Pkn
M3CSiHgdgLvEcyk9sC8z+Z0IVO9rKuExs4Lz4PyX/2/VBaEB4/P3SdUf/ouSTsDBDFTui/3mcOWT
qMuWkKMI7LD4QU7QhX2aW0hjXlZJ6qbipkLvLjwVm4X2dutObuNpksIFXRfsDDJ+yDjZWgCgeuMR
vrAoVaqbD6NWsKPs+y20GucglFSdB9AR4+Bg4Sf6oqNOJgrZl9oxDR9pEPKjVuWorWkyy8LvBKGX
b72Df8lC23SogAFOa4i3Iu5Ora3WrKXh+kTpQzFagjlzcsA9XphT8uzKuSErxsMPOr+EYNMn6nT5
L5dhgPwA6EqWuhD9Vob5zmf6aeyov1YcbO5QptDXI0UNH7Blo2fYTi3Q7/PnEPRJayV0hmImj99D
cudYjV6Mzu16wXU89XNrmsp5jfR9+t2t3y+WT5SW6OmYGWPYW9QTs/31mOz5AdKu1htsdl2idTrr
2SmqjuEDDCa+Zk5a20zwu5vT6vtOtjuv9KHKYnWHFWIb1uZZchLsJ+TNNGimfgZpl2dC3tQclPZm
8nxwdL+5MSnSeNgQo7zJq9hXE+cyyQKU2p+14LpDHhviwQLfB8dIrgAKPn8GUBKYpNDgNPzot2kx
2pvi8rWawif4jC4CTSG74MIdirfh0LwcxyU6otAmNvv6/7QfPlWfQ5nvqkzWDgILwx/H1yMr8vSL
Z43DnNpon2P5jrUra9Lno8sqk0k5LIdfXMgl6gromErgHqoyimGtyDg/DOxipK1sFeHYt7k92F28
uPOyd8kEl8Z9jSMe3mcykY0eyQMeCFnyWaLvWnkpnePRqSVg504IZIIDUOa5zCzJRzZDZWmHNYkE
29oLL72S25SyljGAyFWAvVJjxKRIIS0PycLJeBT9TRfEKrAvYznxlrl+UuBgVLYpQrkxdh5HT8gA
cJFhtF4MTmzQYZieR/2FiT8R0e4xb2F51MPYfib/f6rQA238tY5xtPSNQOYfEGKmNc5maDEs9LK1
IrOZKVC1KcwS+QnyueRpoogl/jSBFLn9JqHIRWPLQ1N7BbrIXKEnWqCvJg3Y1ydDVEatyO7UqIbc
w3t/poVhS4pbxDXSNt2qVzqmUu0L+4SjbIC3vHZhaKj3H9UzmdB8JVXTmxvaVbLwPNVBL1T1/tJo
pTN7oEJYIB5QXIOePwrR76EO7rZoONolbgWeFNRLpB9qyKsXov1TAhZ0wBWPA96tyS3YhzP7zWW3
dOUJLfGTdT+mQx4p7O0ejc6cPVWyr9a6ylXAS415OVRR6U28KrRgUyeFbpb5KPNH0iAsfx2BX17c
Ilgk9qUsSYjp6fe8FStFMAsK0gdfEvslIS36zU42XEF0zdD1kXd/BXTJTKbNehvG/gWw4834f2xf
N/rGDEAgBBqe/nYt6x8Y9YwIDK2TjdHjb6bvOTBFvh++QIYNABHHtm2ZBMZysWF0Mu8G6RdL1s4F
uY/Xjksst6M3BFPVKtqAUm0NJy0y3LlAKpyAiIAYQbtDpU4qUrykCiAxWzBU756J5edCEpAG/bG0
cKXsMFQP2xb0bboC9l/0yIECgvAD7pEoQ1LjT6BnMh1SL2U5P75WIa0wo47IlbJeMzh4cZAM9HA1
yIwLxf0/BdBybX887keX6q91BI2kmCKLLy/qi/TLnUn0brzwKtQPnr7qZBYt9jeQzZ77q5ktBHA9
n49zrSrKzCzc27KU847rrWHgWuLrehjVc1QKlcVGJpNL9vZryu4cvRsZT+0/eGENHGONGw9aaMab
CT9s2PxQ/xKd6Ufwt2VsYls1xiZ4cfZsVl2Ly62Cnd+b7dVeP2FoZwhwdu/1zt3JiP1OEmniOMTo
xWl0EX0AP9fp15pAfSEH/MXTRmlUQ84Yv0OrfRJidPdNVYiMvrmfZTL2Lyo+UWTHqQxGT0NT5ZcW
bgLLeM6VAYw4PQmW9s0KNMR+TB8pPXR0RrPmbxT06XSUPDMsmnYvLzgxUWtotPlnFp1TlmUA5UHi
JojgTATJN2sRd+Gutsp0+www/ODduX3g/KdyUX9t8L3cCw18nS4pKHOTXGA/QdgIy2V12jaBXIYr
E8el+XDH3WSQopOYM2vc2FiQ6+SHI9AXBa6OHrvxpf7S7VuSMSFUxorhwJeyR27InO6xJoAfQXWT
TSDRUnoH5UmlReme3wpwmZFqHrQVcqDVb84mKy3lI1+olce/ld/hmvBbbvWJHPugp26oTRDi9zWs
DRPx0MgZRRYNuOTEhQMeYMHIAGvhtmvsG2zOcW1XfS4y/mymrdpvOpCD8QROJ+l5naGrFZuv9bBL
bv0XL2LqJHW/71geK84uSIBX3cIRS4fJruEdXcP/ClFDI0DbsZoNV+buk8HlJBQkour2THdkoT9H
xnLeLafH9wOlhPGnW1t723VJkyYdUrQ83aj80+8QCa8KlzI2KVZeYtJPDspb26RD40w/WR3is0aI
E8X8rqExUy0w4D7MX8nZBD+pLeJSv/Y081AjJl04KEdg2gec+dbd6eWoPmrmt5JPN8jh5foXI6f6
NGiyFAdI1FGgfCDIFu0YznGyXq1xBtcb+v2CfB6qhMj77rkp8uLyJ7RhFKUxlQEVDqbACAMX6O+7
BV+HFWbo5CYRG4mztAVvn1fLL4pb617zgXWVa1F7uVDEgUBYOcB/WL6Pc959pxvxfuB0tC4VxZ41
wBJ1SpDc3+evuYaGrfQjTnA6dFNn8OiBdtgXQtkNZ+zVFlE2xvT9rn74q0UNIMFPINcXUPTm3DOb
TzcAZYVuTeEGYesb7kL8WborbCxszkM0KY81NzzjfTNqqjVSUfFDjq8hUhX0u8ir3urDSyjigsyS
5XhwJMtOWa1+X5WmJPGuLXbB9KvoBBX8H/yWfaFZbKSQnjVUKIBORkZm0k6vGo4tjPWojD4/xPG1
bzXuwj32LVZX24zbhSn/EsLpZ7bu/F851zHRIN6Yq1tPTPO+xFea+flQnd0V9DslFB/MFsvKApfb
zV99oWTvIbNM67b9aw2VseKl37mNqAzGa1u/8EmgODlxjl6ygFYkwjCMlMZhBoXsX6XawtTfpopn
Re4dUF88d+ueyGvaElpuIqWzlVf3L6A+TcG2s2mCRfXzGJ7oroXd/1ove1nBAJ0zq5rYlYoPdhQW
dM4Kn61ifVLKcgG+qISq9MuMFY2bgTbuKVrI/QrUM9MmOp27oiqZqEMqpB8vU+Hk8OHxg0vwPhu6
PctV0gWsKWFVk4DvuH1ybyR8P65Nnk7pbXtiPyV58yWZvr8JFJxSZ1qLSAFcL5/I0+mTOsKXwAhT
FAjNvHqFfcU55xmPoVGbLpyIGXkkkoaP8v6LiFgGnWZWY+OR/RiO17fxONAkMYtdGATTWl7yW6BQ
g5GcliHkYWbg85h6kekH8oNOCYxQDPgl+YD+pt6Y0moQFT+YIinRiMGZ+gzdCecfDJTkQBuEhmH1
kf3Wjbl11OzptqAwVg4IPCcTndvvuryhmrlFtz/kfCd4IKqk/R/2jCtDCGp4+yclCGllF4oSa1mB
wr3cPFm/Gb79+FO9JinEAjgld05UVYOa01LZEQmRXgAbbKyOCsfaZN0u4qf0mSpXTGNcX2h+4cxo
ETvo7myZDYX/7BtCl1LLryc/plLGn7W0LNr5d5/pA34A8kB8PDjyIQGB736ABOK1baTWQrm7MSaq
hsuAN2kt+Zc+9+PHvDkiXNwd+3/Pi+aCI6ktA/ix+NLdvTDrOieuJGe/gke51RAbQuI4L2XaDhag
/pQ0my2XUFE4OfdQYssf9SKw1YEICcOXU5FpgTgZ4NGTPOxngW6+Y6mfdJSaJZbAvH1d4hFgLmAO
eGV7gTZzXP7d4Qp6RJbbZiGPDIQ1oOyQ+4GGNU3rvBmZZfb3B53iVkxQzBddcbSWC1wa6ajrUkde
v17Alce1u91JMYPP/mfXMEv00pj4GyjLB3GyHp0Na1CW95/aBoR5u8iGXq1gdjd5PiMkzo9QUqUv
snFBWk63KTj467uqKwfyIUSLho3P6yZOeUCDVhOp/hulLaegwhO9fPniVhWEAcHdz3+XkDBBTUSy
h+fIdTArNSUWLY0iWUfzumfKdYXjLW9c2Y+j805vhFNc7r1Makkic90eYCZi4np/7FDnFfJpJ+xc
VDhyKzzEmqlLF6svg4T06w13yY5lToo/jOMUOEiJu9C1mfyZt5rAkbC0/Ucan62v7Eh0NRJZ8e6b
Y4o0KP/PXj/R4H7S8vNdpYnsf9YCpedBqZ/nclYhDoWNRvnfzVxKgg7bCiCH2xEyI1aKnXTNmBRl
ZTF3fZccarK3d2TH6ziyt6dVthi+n8OnjhPLbW7ke7IcBQRau085KgzUfUn5dxeZ2YOo+TEutkMp
Uqw1qnsNJlk1G2CqgjtnC+S2wbyEBaeKeBmPkxPErHY/D5A6FURphvacvKsV+g+BegmuRnE/LAZq
L+IQxTMBcceOybrQcLwyAfkc6u6Cx2n4wUWxeCZ3AwSMbGtW7a3rs2K3OwcBZ8rRbgzN69he6I5G
mS34VE2AvrZnRdilH35N6ZjJe7/KK80d0v3MYOUHTKzFmeNX5h1cSBrglsZyGUguIPkrMvlG3W1F
w/dLX1BOp+LlrcAd3CUEMKWbQMFT0+vEOnml5/bmfup/j6ZwNXt4mKoIiDD0okHOhYDU2C0VNsjL
E5Qq5PVrrYxxB3JAFFlCKqFfOPOrNoDmc7N+3VHCiA4hYGUgQpg+FG74q/n7vcIl8MDcHk4C5ZXQ
MD8vBekZEteWyLf2deTjUK8Uk+qmcptsbxW/zhnQCgRXgkMFLSa9+HnY0S6t0f+x/mpAHsd48Mjh
upc+fSSPkNhOl7z0Jl1nuUICqIlxCRTfxvULD6SYO5B8UC4vcfxtxsVHq/mkAgSmHWqg9UMOKXlJ
cDCHtqTYAktfJtyyBgjxQ8DWXof7RGq1x/jilgI1KcW7nBWpwQShA+Svvt6w4hxqHHPTT+2H7l6W
Is3Q048qXV7cqggM91R1ZaRmwkYIiAG9Ukn61y3UVxONSabZg5flhj6VBSmceq8cCs6MYkxdN0V6
J5dQNttYbPDTgXMb/EmKgpSHS3Vsj7D0reKFGCUcvX7KUsCwFX+k+IaHb1dd2iUkjNt+pzcktqHC
opzlxD/UDUgtMfy0cugP3VlO2xH3BIXm37W7D3gZWG18x8N7WMmPkHduzUzy/LwCVa/1uu0yOOYt
L16g8uHWzLKd7+hDUcIwGaDLrxBKJaBZ2NODFMXoYp5UVuUkw8t4LeYlaifChN5ErtPhQIH2HSLw
OrlRfXSChtzaBdHo5JHZpHWt1Es/DgJw1p+sMx0/pjBS4RLmB4ogLVRz2RfdgzzjJG8zV9XmYN0M
w2bG3nwRvWF8Xi3XWYujqpuSqP+vDhN4pmc64Dvo9rnlhNEk9yVy368h/kBszrfL0JC2wvB+/h6Z
tytLb+oKMVwNm6xy7ClHA0VkMlA7JXdkpDT3ddUZAV1GZLK8FwklQkZ2mF3+mA2KryHcuE+Xae+t
EkUqVnx7YrJgMIKusdkMDIU1C3+zQgVgiAA7avW4az58eWn/IXjDockOmEQLUqLUHuXul1uo1DE2
XiJb1ZMJYdTqzuUv6RxAkQVNesP+O0l9mDfrbNedUZueOA4QxosPKRqwiV3SJFEZ4XmPATTGPnte
ohokCTOkNpCM0K97nyTL56W4MSS8PtJF9E3e9+f6BGY5wWBlWeu66dbgxC2W7Dw/tYgNSINupao2
R4qoSi3rtIJ0YOS1+e93fJWp6F/rKjIZaIbKZnDo2SnAS3WIj206hbFkXGfSnSbEZFSsgTKuBbWl
6CChHGSu3Qpi+HRQnRVdl5Qp6g60IDbMQE7ndydkHXJZ38XeNQmB1RjrGGaCMzRmHQtoDG/ewsaS
GkqIH2L8lP3XhGFm9mPlEuu16ryOLishk/qx2eS3P838PfABmryD/o5CnIKidC/t/FBI067xcBzV
e/OB2O100QbVEK8gJvGxJs4AVfXwsI02M9mauukachlv9RaqzlQqRJiyRfervUBtDKYa5amZoGr1
7gmHsM/MNqzsWQ1S8hpcxpgAWvHHfg1gYXx1aQAS5olok2/Qoh5V8xpVMYL5TJOS5wG8FsDEF8CQ
0zTqfpUXP25beMQjPsDitF/tAHWWe+y3d1yjJNtiFMAJOOedaGH0r0TUEmjCYPYUEQpv0y2ZJ8Mg
iTt1gS7lu8p6Vaw2cY3uHoFwIBXwVfKN2grBW4PvByw3+l3WvINdos4z8zAQCUj4ejJJzlyqJlwh
ouYHiY3pfvROpDnwrKKU7hxqCdrF69OHyDftVRHhCsgM75BpCIWf3hOL+pavzbuZIYbHTRbmfuNZ
id92hYG93fGUF4sXZO0fF/9yyzbspGTdKREKbbLuaZkLj8Nhg8YmkJlSiynj3wsljGldYojTTqML
suVTmUVAj/JeWhWcVR+su8ghnoAUAvHLssF1/hKC26HuOn36+RIZBPf8fDOpRTrlBSN+Fb0gO4SX
0dXmUqS0wIPBztOaQ+neTToun7FzYFnTGF51Z40xQkuxW+23MWHnNbwra47Gs88Jgna3lBZBT+Vm
WwIKHP+R8ADb8ohSbHS8+dbUWL3D+qRN+syNWnhGCnYd2Xs01Q/ubfaK77pPghE8+N451ogEp/P3
pwGlS5+gjqVYsTHuymnZmt6Qv3CbjUFt9paOAFjdJuh1lfRdkpFWfSI284OMnAIGIY+fkD9lYEuE
31bw6yywzAhfuAfJI2UOhrA1W+vIrzHJgY38JZvHcEXKVU4crDpG0V+fVMZHEaPgGaG6+0LsKs2K
+FiAXDnAV9XUyost3LDH1wTKtHfz54piu8P598/AEd5Db4EthOeUMUvxKMSAYtTOXd+PTRdEMdu6
7w5VLdFbzcEWytr5hoP0+aAqsUGDp40rMJMJ0aeimRuOtXJr5ZMdstm1c1cqtOW+LW1NXnIXO09A
sg5P0Z1n6PqI1DhbhhyBbNwGpFQvUTxkBKz/k8GNgm6OGxJ5rY/s/PO4bnR7Ay7YfRIJ0iwAqm2e
H4DR7vBdlnLhJNHDtroWN5MdNCJD/3l+nJjYAu4P1OpSjfxfqrItX0pOfd0YPbRlwRuz2qxKVhSp
D3uuV/4LlXueAbJYgwH7PWEz46HBIeSVSIzcHmcZuIsaAzrwhP45UIZ/r7XVhlrwt5PATrx6PFSO
uw6plUodTCbyHk58b7852UIVXBqFSWL3T6hAFgkCzDHCxRGAG+PxOpSi9Y5nEZDY+zkwsYawl3pu
ynmkOImlBxZSFFT0Wq5kCSM5IEla+sTEINve8oFZrG9rkVtHfhF/dXGTnGwn9y58v2EJmFy8nNkn
TS0dBO1R7rR4yj2Nifr53NTI4p1Mcs8RxGdmQ6gDovhBsFx/yJiVaOWT0Oic7bF36otDQJb688Fr
dUT1aUTEElnV4qLnc/EZR6OrzAPqsI9lAyS3G6UZzzr0LetGJ8qTIafnZ6/KHYWKbHii1W9IrkYG
FzRCxt3xfVAn3va8GtHGY+rbJC7z1tXbVTBi6cMJmjxangecC3RRanQzIm/YzeC3pxlTRD+m+XcS
Yd8OM9CwuX4OrvskbzhqWHbG4rewyvbCQvAdtkZ8G+f5AinPudMCLHxdyTXexDeNJVE8VBM6o9S/
SWIe8oRnOCKou9GRpr9tfOeQ5g0VGWwevifEaKffM3qozMxd/OZd/btDyOs/s3GcMByWM3poWdFn
gLMY3zezzCGsf14DAj1c0blvtP6bNFsByolA4COEDD/2dVx7FJWp6cQvp8rRTAqZey+eWSSQO35c
ZhJNuI3aqQbTUFNBM/ZFri8EVfkkos0eGL/pnqJL5YD5zc7CURQ4cUKmsmSxrmnQ9u3F0InlHw/y
F3RYbF12ZOMve2/b/e2PBWupdS4XiZNKIKC0Z867lJR14g4V46nxsksS8IMXfTFL+8pW+ixYFS5S
RvavinuhuWzcv+Snz4zEfPJ9ZBCNUC2BYxzM9dSEMOcYfeHsjHOLLfkRwLrzjOXqB+tcU2wPl4fT
GEe5yk1LGTRMbMX8xZKLIDoXSWIOS8SnfVDLyiTg2BfF4OX0e3HIOszFdP8ztSKuZKcqoPZb8bua
mIFKBW4SX6p++J3KLlM4CuDd7d5wud0VuIMMWU4hhLC/lAiqabLx6/NHM0H7nPAjxILL5ReKlGhe
fz08J3nNww1KxfhXZqiGmf/kysWToAiQKqgDGaHLbbO4bXdzDWIAq3peQHUzNsJ2jVD8qfwmo5Gm
bRNjX7/7l8rKiG7sHK1b0EiDdpW60+NbLNR/AZqRdixe+wIx+dBx9KLNgHuCgIGkfJCVADrKMNx5
05ml+mBwNL+xFX98KjRFrgUEXdPBim8+q5PFQgg2GIodIhX+Q109mPPIYlftwcKGamyLQd4kqQL9
di3258ek8rsXcObU9UYfktYE7NhqR4LZUShcS/nnzgJHtFu4V1IChfSsSwpHEhJXHCUwfDl/a3WV
k7AeW2lzsMtbBCu4VrR1dE6IwD3b+q4VVwBKL7nfZjYGQ3iMemMJpLRPoM71Lgz8MUiP9il+95jL
Mv/U9ohXZmG9/m8RCHqjaDpU9ezk7VBNrv6eSTxwhXplMN1kDdJCqXA0iDzNiEi9RcsZHtJs/t/p
WX5uOb9IwpvizNDj+E1wDdqP88kCRZMpdWULxgZS+0SNMZZml8F9vvKwAVoBCtPJmIR++zILkzXa
NZlrC6aKCLZuaVLqNHy0NIyXp1zc7vz0lTFnmpmSl3OYFYV2avkQM7FPPAclmpYFRdNqTo/SijjL
ixMNZL9higMVK46Wb0Yd3x0adihM4lGp3octZ0ptFI2HsUHb8fizh3/5H4IGVcpVL9ZYUJktQRaT
PV/RaFL1Via/vwHSqNTuOjTrEQoo8BnrmhasvGVOurNOVeZgguCmEkTz/ipqLE9tvAvgbD8CaLvB
xcTd/g3b4tt9Z/L3RaJT81O0jQdseqmTztPmehbrMsuhWxtN1FiCb9aZjDrXYTbihoUagwaM+ZJy
R5J3ZynCI7laVW1+42NKFOpDkhQCMKK/ugd2o/p5RUDYAuaQZ9RlufBPaY0x77SjA9BlyLJcmrJd
Trj/l3h7vyTnbd0RhDUJVXlsSjI64o08YiM8AUXr5gr2UM/a9KVdXfuAZhOSRUYvLUqr2cUcG9pE
0PwgypBS9K12Qjt879G5sCTkB0jsKMM0nZz+TfteOuv22+0Hdmq3E+POqBQeRRRdfa0cUpJzC0Xu
r+ru/EzhZ/Fd2VdwQV6dK7od2qaMMsN9bIbsL5dk7SYWvKwd1UTbU5pMOjjIpdsDK/i1ovqMaTxP
ORkErSdfBlyW/4sqPy+Zy3Es3C4E4rd5wfY6EoDIX1VocpqOAg8l6Oubs0IDcRVYi1X37l6Nftyh
Uk8SArHfXpv0sSweg9ur1J7bPWrwH16tXc0LKLN0QqFdEfQfLTdDRZ7vJQeCL8lX/Cdh5Vz5Uwfr
e3nvQlndKarO0pLx5MNMJRDtkY07D0HQ6uzthRu61PBpDQT5aybtiAiDRggQXoHDfCKAkseRpltL
JK2d9qvCn6oDpnaeVmxgKLY3ult6WZZATnqmKnnpc9reBAXW5u7d6g7yPEDTXiAhSUudRYF+XqaT
88N656KjamToDyZBm0MWfaUutOZAbW7Ekz0mEpiEOR4WI++Dus7BT604ykhHlx2A2NKzDt6cKE45
owMmWb1+hqvfXgwsbvY6j94rUNwr73wCRyTdf/UcYJxgtfoDXAb7wF1b6iUiDhyEw2sbGUd8Facl
k/TsnuFKQKc/ZcJ9BWxxDJsHYqMXMp+ubopQCE28drD/QD6GYjUI0I6aDB04+w8V1FrDQjiOgcub
eVUgha478yP1IUC0iKsyUJ063sFDvVSTyGgmq1MtgiEMjSD0gmFh0bFGMQMdtljhnifhNrrkv2wg
GBY6PMcjstsSTZZtovD3HSTGSwbgUzckPAt2+l15aDBoETs9ytTjxeQowDM1yyQWAJCp9dGwR1C1
s83Z3YlQVBZcZZEK1gj2rYQ4jFufSiRgtHvCfvWTflDD4UOyAgTupXOTs8UGpEvUbU6fCr82JJLJ
KSwL3iK6xR+9G46ue51++RvqZ1xUGSG5bzHYziRPdDGD5Z84m4BpRylejJmu0V5a+eG4B6xH8IMr
G/aT9zoMkJEvrQgluqha9LdZpFUQJ/PnaAGJvdKTs1a5/iJvppUJk5DuezIFoCRTXdQrgFW1marZ
JgZMcQE+IXBCNYNZa8RwuZ1EvJdlJEoE/P2NmVOW9i72cumpRpXrMlvZfNlstilWhz7TGgOdOQri
HjrR7eysesPDAQ+6ShAxKK6WJmSTIvgvDg06Qi7jpVaEni8h1eINuzEwF7J9DsSzv+ljVTZ27d5o
06Z3S1aumun1fm4CiTfCMhK+ElJ37Ltooxf65uzO1iquF8Q5pHFIySJ+i24PTjqNVc1KM7I2Mv7M
MUW0+8z8BmtEf4iabxe67uYYkF++hi4a/1TA1y+gdV55iiCqpEK+v6rRkqoJk/J4Oc9Wf2CHo4Bz
NDcpwCLEhEGBJa5rLup0ZEJPNGTZQBE+XRUqTH6r2+Ik1luevA+T6yq5dPwIF6biYwxtv1WR4HuZ
BJvROchshqzqC5Sx+0OpRNnHcIv5mvIvhtNk88JkyZJZqPfM97QFdwNs+XgbtF6RDNnGKCdeQHUd
oE0ySdzylBLW4EYVUpCKfD/68M6S/OuwyRLnoMPHZGXsUjyBsKj4bKMxiePYdrducCHkifXtods5
+Dov4sXZTf8vcgnrxXw5FxaZdS8LJdsNrCmIrWsXw/tFPeLgG2gIkdJg8yb746zWy1m5/ixlvgFb
6kv2xRFcrb/KvwT2Ubgegqgx34yGMHaU8OKGWNTopU6NZ5sbfGlqkktK90mUSHLTsGPm09lhJ2cl
r/i1nLd++eXALRbTp/Bt3adeJLb4iaketdTigiyCF3yD/U5g0cU1RdXuo/JpGB1ZXymDlh6NjkKt
hrTSIy0PdvdAErS3Mn8f8nTxP4KFQQtZGk8Zf6Ad0EE4dxOUyti654dsskzdH2FZyPlswvk/SbJy
4qgMur1N5tNi6YG4hT7mkcZRLhxUkrZBAqWJmTWE/p/VLT06672pJqct8kB76ZWbHoeJLkAwByLQ
+WpMd2IW82Edi5KyvCBpIDJUviNYBL2GDTHeyFGJ3w0uT2WaOR86XwNBqM5uDnd6IaTXdmUjtXzy
UWjwxPXwW6PvengWEXH1xKIgZduGQHaGAyx0/bZ468YUud4sjbX2l+dutZput7H6Oz7hikJM6Rdn
DGVGTE9dPCjPCjpAHtpfhANrtn8c+45HXZdBrayIKwOkvZEnY7jZDrgZzZWG0O57Txp+ofgJKmef
BZbTLWnKm+RJUBfk0o8lXn8cQLkw6JPC8gHohAQm1MfH3ctTfhmk0GY70hi5T5Ge2gWTevQQMQbl
yiLfDAphHXzhKZ184j80Sz82rw20SVHLL03nraWN1u8RNGhr3rKp4jwV0+IeSmtSLwODz+7S6kIG
hXciPYPbJji7CXiSOzhq6yN8wWMwWrKjSvrdOZcIN3iB9YkY3s/Vy8CTQl4l6XNgEviuiH7lDlrq
J5sL8eNtflwDPBES7kw9+TgwhUWb71VjrDyDYYbpnlsj2+WDTMQVOMOj9+oNc4Nz2WhxSNmvYJ5T
EsXpRKF1oRjN93i1WduDhrZVtUTPSYp7kmiLrvfBvg/aQAlhi9fZIzrc0nevZPvQsEIHn07Jis94
ov6JSef83U24TMkbAg6q4hwlD5LhXxJGy4tKKyT3Cotxq3qdf/kmmo6wSOE+RVR/jNywfmNhl2rM
gnF8ye9gYghfm8Cz4vhpz5Mt42YJ0DYy0C23gGF2bC3J4ofv2/Woj0tIhJLk/B13xfB5x5p4/mmn
3rqTagTw2tahLx6/KNd82J5yOzTR20A028nxpog+CkpLg2jQSnL6O++YIcvu6mK15Jd+WtaTmU7m
3VZfQO9syt4EECjb+3hpZy0H3fV4LGQiBzpS821p1nOBGv/PGeUS7aVXfor/nJZTjVIn8gM8RhO2
YKI45pHpJNxSI2vp9CXo+iZtnH6G+NEFuzmYihaFmkVlYkAuVIpGdgVH0qODuBSotLjoZJ8kTsc8
5nobFsWX+N6RfQwJd9YMw5h+gItyo/msWPSarvpRn6hBy2wnlixD7EySZMM0jew4dA4FxreDPD5V
7dv1XpviXhrwrOjrYGrpdJyNUVow79FRaXSnOJvbTkzger09N+xDjio/0Klt5t9fRwdlUUk8BQeT
QOen8lvyY3sxCGmn66AYTOXmgZNlqJ0ZNW2gTfcH2CrcK7kNPuVBzLkWAmU3MUK6RgJf7lqPE+VK
SeZQifmj1dqg6PqHBoz+iIKS26FikojK6XI9Ht+n9ERXyTCp5Wp4dA9TCZt0Ckn5ImWdeZHqIkde
87cinTLad8bcnDXJ7VMS5rgBblXI4FZ9h86mv8aobbGFGu6MZVYiUdqZe7S169rVWBJUP4Jqog7p
2U44FEFXzopDwJLAwUYonfrk0QATMZXAT038wAJsWu5Kb+DXfeEcuuTyFhKwfRUKKWPc9E1VC1wK
aQRPeVdRpFeX6mpjRCsfPZgv2FM6gCMiINSWxMvj6JbUgLJw/y1MT+uQa6PKDb8E+DnBEZbgyebP
TT4uoxiNbIPfwGj6/oQ7oEBfoBkgE9joed6lHe6QxaZwQbOkvrp3VKpERIstkWnwLYQ6TMj4qWVr
zntl3bzmmm7hU0xUgugpW6fBY33mr20KmZJNiFc++XJIPFA6Xb4YRqwynAYCoJpmQTYgK0AZIKNl
otmCZ62FmH2jM6DxyBrghe2E1QmnT0z658O/gDXSiiljQngKQWD3mymupNGCH6nvGR60nIX5EFQ+
2XHpOfOqlOHzXoo+qi9Lyx5mfTH8NPCeLOT9Xt7lHHkpz+g2qqZQnVsmHT5cLrPNoxgA7VVfYY7D
roxoFbmRimIj3xEON3lM2XjTqZHphP0jhdVYsAn8FRB4bCzWpWqqp8gBTUeDcUx0U/5s8VPLNegY
91hTo2rmyCg1E2byJqmJB1bKZvIZWWFZ7ZpKQrwZmnkaIRDM2pmgUnLY1/B8uDIsFxG6ikGJ5bv6
rNJYO5cz0Y4UVeQY4TyGO9Dm9OVdyQR0FIjxxHXWmoZ4LaYe4fo+twVexAq3qLYHOVGlC6fXNH+b
TWIKFzn5ZRsHyUKvm9+7pgWPvrcWQE+AFrqkOEOoZt3IhheIhXZUjB3RkoEqN47tyQAE876gZkeF
7vMGO47yDvwW0Jm7SeY37fMocjD4fA9eT6fkarTwxZanKxO6XQW2/Kofi8FxD+UQF6cWuaQBBXRa
KMSx7ys5AjOofUtyu60lQMmtTgFXilfBscEjFNXARh4kgznkm4oyKBaeP/G0+gCQEpR8ckEW5Opn
siLsSyCQ+IpOzaIZVE8dY/3UqcZ2qHJpA8reyzg38Mza4VE4xg2kl/qtLYfM/xQNWIou834zxFSh
nO58l1vUvKrHG+D04/UThcQ5mwL8wPzZmcIKc1VAhR7bd9gNS99/fztHH/79kkn3W7FGB0GqDSdV
7uEpihAq/7MvvNHR3fmJOAtzdV/4hqcMkVKpwgAgmpcTHW9SisaPDbrYsQdEU+xZ0z6qeAzdyqOg
cuy8Ybfq1pe++5gPb1YpgEc1FihgehJwgVSJU+h1dJBh6FJE2jjen0lb4sr2X3Z3SWzEBI1uPaHv
VJaAp609HA02R2nZAiXEFThToHojzzDl/UBgjOm8rSOmjJA6FzhGAPzAX3wee/4J/wOiQPRnPKFb
rtwTfrCnu9B+x+U9kORr02q0eZAzCE5sManzoDE8borv26uEULTWsRcaKNkbaRZxX5a8d4grAM+L
jlHxDze4vbL8YBAItlF6FMIFWQcRQtVSUNwEwlV3+HfaLGn9Yf6RqtMjozrJlneaT/H5mDl0lwc6
rkn2dZMAG1+B2JaBeuEnHSM2iVbwZPD2iYjW4+U3qYuCyLv/jyc3LUOnGI+zvslyhaWXijX7TeEg
udZXtV9X2wNBjNZJt8s8yaxCVmGIr+QtQBzJ5RFPtH5NC0oM6orWGmXaRd2T0J6sI5aIZMvrnXrc
OqXcsiN3bCiPyoIqMNi+hZXKGDvxggO0BpXrtecDrEfgHEzLaSHCaogNF8ikR4vjI/bLZmSYb9GI
oNY5gjMFL5sq0CcISv1X/W5l68xnooTdX4lZas0uI1SGeMd5yMkQdIsMsfcXIvae3Aa6GbUA9+kH
3iQntjBAUkP/g6FJS1k6wk9MWr6ddFFRMhlgAxE/xCsLHMJ7fjFNz5px7RlojLA6/4w6lXNRdDUK
gA2tSgYs1XWs5sGMTHm6EPkg6p8f8u2l9DwNRj94mhxVplKp7ro7Ib/tQP5q2gWcsFpZFb40+NDN
0o5GVE1gdMkXTOkDQ8rhYnmQzOe4FKQVb6szu4jyu56LluIytgmFrjMde/GFC5PfcdfyIDgykNMf
kJkRRepVjL0WWIZ5kzZOUMMNbei+QOWtdXT9+RuWYVM8rOEvhUEKicjacZzHzgXnls6WsOLnnct9
lp2JX/mcpMUOVHsoO63RjwqJ+NQMF/BFsXoqK6XrJfxLke2BM9JDlwcCG0LAE+hHN1MivvA8MDES
Awi/xquD1gnUUIxDnMLwiqQu2GhjQoXJjygsjH6T5VlZriC/Rrq1YBn8XIVX87FSlCDKdvCtqT7F
lTKo3n2dAbzKEKemn/lF+uh3T9tRymbxRGo1QHAEcl3RmzBvryIxP3B2mlb4j/+dT2GePgh8H5jm
2ZMkyQTb5xYd73S/WTsn1nuoklH0SOddufpN1YHxD/sdoQUR2KZwUu39sRro78FKh/G298MWWyjT
JZCu+qHwRPXz7ExZI8jNgkyPaLR5QD22M0jBKvXmTxiFp0onb5oQmAf9QpBK10eS+S89HTS2/oKG
EesZnlDS0ogG7sgotP9cZoj/axmnkRMDS8vg3Sl/ip8gHE7ZC1wAfQZKbDPepa86el1MXL2rUSXK
DASqQCSz4RWhOBg1usIFTkQhDL7Jzw8v9ydOnJJFnwHLTCJLbHDWZhiMxaNRcO0YCPuRz6CPsQSR
GY2t4zz1yRifaAz+m2zfVnyR3KYDuhUbq/+6GJijKyR+PpJnqe0fgseI0ufAxsLUGOJcs7FFAxcR
33e47oWZ8A3U0tsVkeOQ6j7kkgeMBHN3j/ccU5mo97Q4vPNEisoJ/Gqg+FQl4XZV0lsznQbG/Xbs
ZQUt7LZjQV4xAui/LHnJMToDsgqcUIKLHTtsEt+pQIB30R59de6ASc5pvwHmI2Gtmf+2mr0IGFSu
24KJzCGqKntVc6s86iewh7zRJ8+RufdRJSJqvrA6rpPOTG0t5q6nONyRn+yPCLDCpwwk00sQLGJG
x6nfA6Gn9+pPgVrZ5Kbx/3lDB1AY+JuMuUz5MIpMymn3ObVJbsPfCv5M4/RTW5BlueRbjuC6rt7E
ByAfBQdeIm+nBZnhcFkCsMa1sL9cyA8g9zvCEBGMTxmrYApQwxwxqlpCmL5DErWZK1dLPGCj3jYZ
D9t4ZgbJYxNHKy0+SpQ47fAk6oMPI19BSzo7nYJZTK3dzVcNzrowkh0i1HAIEGU+emSAEebzrdUc
5L0Ry4zSBriskUHSQHi6cIBGkB7hgZglVX6rOoOFlqQXcNiepeqVRaGfQcUoCH8zMbNv5GHMLRx6
uC0pkM6Jjc7mbe5Uxl6BlF/cxYqzrthBZD0qOcfAoUAggMSSqoQXizZMHTh2YFymlWWNCf7vkxSe
F8lDP+X2s1ypAKEkgbFQvdmaiQNNtGW9XWFXvF3oDKXJqP8eC3Ryaz1JTTZi4/AujRmN/xn3QdJz
j9Ey6q4RXLXlpf7QETV0vZHrjH6JE4KF2XJ0CKRdq/1xK1qKKELhZOlzqZO7lqzv9gu9ZBoEctsN
vhRYF82gB0ASpn81/WHPz7157P2EPGIgqJVLSn6WADccEBe6OCAa5wJWxnUsjw42ZY4CmTXiyMoC
EmObcQnJvXIg680Pi2vDYpZDmB4GWcwkao4DP0EWKCiMC9uxlI0cYVTYWO6QR4ctG/1B2RdQD1j4
Ky8YUFZk3npxru2hjYIySY2pIrfJRYo8AcGNMWXV/U9eDWmMl4uKdbR+6h/v3rh4vsy31ZUtEHXX
zUD0C1EWbOy+f8nmv564C12mVrvGGI4aKOGN8oOW7hmBdDb92CLh5ievJjxO7HuQSpAb1f3DrO5s
SYJCqxzorkK3C1ZDRUNy3uEZ6S9UA8lYsMCGQHKGSog64JuwwbfpIvwdcpWxUEMSsDfFXP+aX8nn
Kx3Pk5dzyeC6HMSOShaREnkN764sqqhJFKHao04V9qccpjhLygpeZMZKzEaK8zhlmkRdQbvyETNI
nkxgQO7ME7XyZi11VAjIaanWBSw7QfMDbz9z2Z0qw5Q2RLn5nqjJ9BmyZlCg42eMi+gzRRNgtf0F
gZpGMlZTUEzs11BU3PuTwniKy8vUOg+ZtYamYJpli6QHrhKB5gp8YU5V4EBfwTwIicPn7/jS6bWH
YDxv0fK5fP/ZVLxPtrtQGBPPM+Nw/WJ0y6uV+KKeEclC6dL23PAXyb76DxTVqlfAaRoS/Oz2MUVb
OZ54FYF/+evZscdiUCh3DY7nQkuK2u0M/o3SO7Ow6ND09xg+P3L6DBQ84ZDDSJ1ikRWPAWkf/9aw
M/YiV/nOr5KfoSmGYgeFs9M2R33yuB6ICUYgP33hvmc6851DgqIJAJXmhqPojCE9joTUb/cYCEzQ
pjkheVnpCCZkL+EqaQLYhSaXj4MLpEGRFmXf7+yakQ4YeQ6haBxjofVz5T16DEdKcA2G5ADS5NLz
HWHBxsr6uVjQv3P4QcnvTKSy9z8NPr7P1/eL1wIvpcKlR76ipd7KnnKUqE1jlbG1srJ5qJ7ulLFh
hXV1VPD3veojBYDmlpP7RC9nz6Ueo8/fDaGdMdO87epvXUgMPbnD9EyGUoid4BLoGY5dqAxS6Uow
FQocF7WAA2eNZVKAE9in04k+hIp71kmOL73xZgmZKlxp4WWklioxCNe2ENDOGmJ35QhweC5U22Tp
GTbmAjpJ3uRxIMDadk5N7i1lmv8HhtFqpFnqc0mRUgoqhVUD/N0PkLoveGmKHBy8JdjO0/9HwKGy
n2QmO8TyL7dLQ72K1OqFrWgy85t1SsxHd41+jYa4gepkeiVbCw2REkUWPcS6Uo+N7q+7F2JSa1Sj
HWYrY5eUMN4MMeJxMxeO1oToMWhzqcGOhz6ynX54A0yFxRzfUgZYBYlZt/gHzSFkR7+1eOg9Z5hL
G+Ioawi/se/mR2E1RD8OgrS/RUWdosrtFXO4CF2c70k+kX6Bn+koPavKwKGaBsOx4KDF9gYMK3RJ
SPjGXB4NJhzi+Nof5RW2838yg13yRHLkru5jcB04vT5lKG6LKc7DOhXr+t+NQZAmx/Wz5PVfm8uy
79m+Ua0nXsJ1QVjnmKZHO47nMNdHZ1pkmW9lonnFE4sv04dwArijWcpYSdBE+FOG4a7TPKRQMsCr
Tb2Omx2gK/6i47NOEhOVP3/G2wfwXRzDWS5C9AVUV2llZ0m2QPBahqoliMI89tFJ1Nyw0oBobpC5
Gtk/Omta6QS2gO6EYguuvy1xZ5tkDYyK7oYEx/XqyChCFwW2XOduv5wfVKACZj5lguYmw7hV3TZ4
QJ4hvIQKSeoj/Y+d30iSRBqmnfKvpFNT/uF+QcE+Y+hemaJlWseqAuzxzn4GHigdY0PU/fzJjadM
vV+VwLbkvY8Lsc/a1W+t8NjOVKAApCvL2+q1yFTUjfuipcSy7217B3jecxK9ZdoJHkCYzgTw/70v
noODvh7dYlCkNRMKSz1yUFO3CRcjUOK56Bu8pFgQHIhQl791Q9YoAEiol5bE+l7TFgv4HJ8Xg01k
hMd8XrYZ40AQ/682zdERhdPwXrZeWQdzSyW1jp06P3ffcBlrFaBFJDnCd/aS3F55W3QzkbyMoYJU
Y4bZNedqOhyCozkUkkNbermczQ0PAXMt3WPgga6cqj8/xwWUikB/yGgXTzoGPswZCDNAl7F/Ij2H
BpXdlg1wZVoHcehWmXTaUHhswArqn0d+Qxo/Qy8kYvS4XYUfHOYTwdn9y3gc2M84DQzR7dFWOkJl
019zQ3oocko9M/KK0eMw33le5D+hNILMaByUZ8PJccHcubb2ZQ2BwensQZpNkCuyMFqkrR7M9FFD
V3w6mySWX5JTLF9t0BbpgLjnCq4uW1krCuxs/qRb3+xvpsNQHCj8a/dwTMbr4FxpwCiHlfcVDQ4N
cgEyzJpHj9YaLGYUSq4w65Lp9UIOQQMYSjVuEk6/ZgTn1wTDfVBExQCbmlb6FyD2+1GLbwDz167B
bZ6WMdfPRcHB63XMbG1iUCsAF+7vjoyztY/CgdSQ46zVKZaJYKOvLhACjfHzrW5y+nKRWQXLG02k
MEb4a/sqJzi7HLgoqrWwzKRQRAVzQs4LlIzPsVZoK/qlf+IJupsDbteY3nMOoHrGB+bLt11ekOV8
IYRpdevCGPizwxg4mRGavlxVfuHSX1qxldhB7znQliDx9Xu9ntLgO2MEI5wUlILhaqU6YtjIZSwu
daJuBlg+4mZYQBir8hIJ9LetnWTJ12L4FWIR1S5n7LKMTsfpr3aJY9Z2kNFsqiNRt7md46ecDQu/
uRd2ZZCr366yG+/F6hk2zj8SiJan6e3W7NgjodvHYsqoBiFecTX9OpmEadD2qN6PhWaraVC7txNO
0wyi0iA5GzYeVc82uxp6LPPkNvFEVXhO5vfwHOsKjEG+Vt+d4JyLjdk2+WenmA0MAwr1XMjDUZIS
vFGo2cK046LIgFD2fyuXlTa9UCXsnbvhuNMC2EuKg7Yfnhd++EQDh613NEkPTisSoM4Ni58l+xOP
62HCmYA24Z0NIR0w5h9MpWEa51bU9lATEJ7DYXs6saUVg4dxyzKQ8RMVaioGd5T8ImgMrEgzuGRd
FY6Vui/lt1ZBq9vrxcUoHE1ACy+B2Vswn51Tkl3aKB+eZPg8biC/9yAd+4fqiU1iqwEo4bEme1hC
yrpu0k9PwHGis8VF2w++bmu3Icb4jTW9uvCRi1orVpdgX2PKOIDB/HrplRoNFZQ+V4nNQ5jMwllj
XNh2wq0IzBkaCmwuUEwVp7rPTDsNSzq+w2jdEP2QW2Uz+wyTaox50lrjIn21LPmAZXaFFW+GALgp
icOnIyKQDWdlBu3fVBGhLNUCf18xcZH+BElHK3TOenNqVIeUEY903HOxbAY63TM0xaeJURebWXiQ
nJjAoFUNdrXO04XRgj0dwR9aoNIporfRcvHtGu7K2cFc+JlqJVnajEpbQb+73JEmW+LvPpjtJEZ5
daBWyRrc6Cwx6IH5XQv3stuyjT917grhsrmcZQfnUOxkQot1vzCW5eZ5SEs1/tH5AHnhYMD/RPkr
0YuakqXiIZCRA7WahThi0zksHn4/qSBghUUOuCUNTKuCpqD4So5rU8IlPG4lkb1VLCjlDftfYPzD
OuuZziXc9jwuhCpUs7gtKndfR39p56ZKUxi/JSI9xwtOax2wgyAj2Xpy8iCR8kFsgUHvZjWQ527W
rg6yBkXrBhKFGQ0Of5ZPDyRUBCyD8ha+xhzBQwzRJLPM6EqmXgBxvrRT11oKBeqBz9HcBBOvpBwl
iwf2+AQ8EI8u+mAUkipCAdxN8tnMM/J4MHXscg4Qv93N8wkCFmZY/7T98OZ/tpDZHzyC7uwGhBf6
AM4lWTvObuioRj8V1j12OGPG44yMT5vhBLrBU3siJt0a2oUfs4ODSGUdbTHJIzof7o/vsKjlyVaE
Xdd/PDMkpER5UFnX8pdRQqfVFRBQA7NueqJuaBsHCuoZYl7AL0TP8PBOavI8CN584jqbl8lsm8m9
v+lLzHjkrDbtKkw1AfPOsmGY/jpNlSfc948gBKPNfo5pfXrOyvTJmp1NJqZYA927xVQYFBfnDkYB
sOQO9/4tDgdrK3EUC2BYsrRNmGESkQCxvkpBFr1Wof6EIqoFmgYjHc2x6pGY/CzBNTaAbRryOFy5
tGMRu/ggVbUUj/TgGcLAhIU3MVhuN2gAKuHQ2J8WcBtWvGL7Pp8WQjZNTln+NU84E+SUbHp9zUsc
FzxmKnLboii3So0NMzxiqLV9jeRhKwiskPUEHvB/1q6CyhpijJCWKy2t53/1lMxGZDak7kQsPCR1
IxjD1oX1dNkWa1Kf5FH/X61jBBh9v4JBwK4GW8fO695oFX5zz6L7G1Z5XmjudtjxUdk7nrQPVyX+
ea+cHtzzPQ76ySG3mtp39t9OFrHidvfPqeyd3CUThhBmk5qzsSAZuyL7dBPHsRXyFFerDhZVwj/i
azKwTTDDV1n33OIeeAlkTFnG6fcnBZ+edds1IzhdX8CcJ+lt1ENXSkaOGP3ZXuuZojaLvEQNQVRA
5W/8xWbzinPFJMPMdn53PDA7F4hOPUQxSLLjQzqnYqP2JhXt1zr6+6lZgP9a2TOP/9tBOCQu8dTY
q6/8L2YJAHuOjD/A1CL9mQ0cK5SIZ5CVMa0iKnRc7PiA4L1ACeM43VmROo2burIs96S9SvACzNVc
AqIgHsK89kKix1E0cJEyDGMVRizqymKnS1Xfu5jPcxAaZLGxE5zPhnS3/IS5uuZZ0voXdiQQ7XC/
k7xW/5qaDAUrJr96qtbFn834FyymsK20Pd0pPb3Rnu0BGM7ufAtMfBe6e3Lv2l5z+1VI4Fih4p2C
WLLDeTafxHuTlciLkvkgLR0f8cEM9KbYlIyFuHwZyPGmXK2BS+FA9Xp4lacePlr2iDtNJ0w48v+0
7y1TtqsIPt8J+Q+CAMDAoktfnnzpsHUau1fuMB6+4tfBIVZ0YBNZCM7xPu4kXs7CqU5IMLkRyion
azFtQ3sM3umPXBMsbKUqUxSy7WK0IMIqZYV6xO5fAmHJH3mSnxFN3WxmXRd0ofTB97lqEig4KbMr
ZN7g7JE1YoOkjItjcEzQKbaqmlFSVa5p4hPoR1mwC6e+9s6OM8G+MZo2SWGO86LZlY4eJwneSoKO
R3aIj3I8k8VzQyM3si0wbKOG/F5ZMwJsyrOHZqvRH3VtEnUGfDK79m++yXo1dhEp3kjncoGzFAzQ
opF8bV5ddn/1Eq66VdIwv4jfvQWFilPXWsLQoM99HH5TQu5WbU1Sxb24cScLIYzMf36XD1hZyldE
ErzaNKniSxTvmTTwQLxLaKGBAJ9iZeWjQYOg8L18RyB7YLcn1TTXTEE9dGHOJ803Jbkure1V74bb
M70Fg+t9JRCdAxqy24FV9NFGbb493JnJgR14q86tyihG4tGwUIxPsaAEStt91ADyy1SiNe9YlKPN
kJ1rJHjEgxKFuRnZ7f3GytHGUmQuNsqrm/sQiX3Lec2PTKrpzrJ6LVPqiIyY3SswV4aRxOTPPL6b
5Cn8qmOaIBlsIVdJfUOLqd3ovVVVlJyoc3Cpe6wW3RXJZ1FrZnlL/hh7UmDaKm0KTlSa0eACWoZP
nyhXTSExuPeSmp6sO1hQL/4WkWz8LBAdtqdBtXaYihZAe3ejehjnFmnsQTRU4fXYoNFvc2572cfk
bPjHvu9N0tmmIFTDaWCkoyRxwFHoWNcSUZTKtcAkQBcOhXsLDTBb4cRbRvNdwqqOpMF2064dioTa
vpmsDVu9lWkwSEarRkA0Q8avLCd++XYnylrYMfJ87faynjsYgJ9YHE/nZOkTLRA8y5zxPw0MjtQD
KSayJau9kk61nVj67Zp0gvTpVraSkOFnaDgduq7rnMRE4syvFwT3GRE/1aw++IOo+SJmoVoUQl9C
rhQVZ5LKQMs8DMG2EIcN1FTLiVouL73hN5yrs/1jKyKUW7aQlaTbu3f/aNXZIRT/N0cDbJWAczzv
PW2bXFj8TmV3fRL18nSTL9I3QGC4RO6NEnRmZkr176WFNYBTy7BWRuOCIU88BB0sTbImCvl+vZ7R
26e28N9sMkccZjDsMZnlRxb2kuYZUYEjagKivfP5yywk5ATAHFvRWsPAWmcyAdTA+1HjhKcg6KM3
5XsvCvZf1722eaDSkFItYDKzCo+uCAAeFjseCQZAn5nzOB74VjjDsL/unkc1L8Dax+Nw6B/hsAnu
YEHTcZW5rQahyvRbm58BcBKQXTh66Lz69lPZR0hdob4vU2sIZzH4J/ln959VPISJO1YHwN0xjQgz
EWscEeEyoLClOWQZEveIcJPr4XrGQAMECJGaJPaecGhALGb4HueHN09yRiEDcSbfvmWd0Qj8Epsb
uuGhRIJ9/LYMwPTJvKrQB1cyiWZRoDSU+N30/8s1KIYwSfISWW1Hcv+10jykI31DHH4mEL9BZges
mLHS0dQih3SDgX5jF8+zXGHzLakQLkz01F7BWgJplKlLPDJaDtePq5txTYTY6aGrwIVPO2Ds4SOW
ZuBlon8QmS+G4YH5gtGt53m2yangQCyyTy/C7s/RiErYbBwKlFgWL9pblnNxhbP7o5J+2yrlMaqw
jGs10WY7pSBIJLaDd0e2R74/hEJlnEibnkvYMBmJtBqN98VW1FZD6zYQBqUR40N4tzgwXyUK2iH8
6HhpG/uEc3JSaH1lxQZjUp2rohVS56Gj+1s6DDv7OWZJk92Vy+JNc6LBagTMlLXGtxgWpGTI+JvZ
VKc22IUSxdHAwit3RpF+cc75M0KmiXyVhsbL93XmKGRBcIVYVNueyGlG7vFlHAOjnzzF9vmktrea
8OJMXU3h+TpyCAHY1jCTUcWLRWvTwokSvlTQtIxp35nR9NVHb331u0Tesoh4b6/G8qGKRbT2kIuG
cIUvgQItDWmalrBrPkemC14zVNlkh2OJ+BAd/GvGhHtejwS9x07M30UacJG6hM7ogKv5dd8uENPT
CbrkN1JAufgagnfboOrJSPqWzuqMYeGzxfnxEPEt/FZU9Kmo8e5QT6jcs1mOY5S08DAkYGELg3LI
xzoRzC8zs9h4kCNayjHiG1db2GJ5wuhoZ/EKFqi5ug2Am6QsjhsDO4p7+qPaMgFtKWkA2/rBLIOR
eUMk5VWmYGkvMtKSV77qnA9DJbtqn7MeWwimPeGwfwezB8sPgl8UwLeyeiriH4MfARMDChra34tX
avllRFqCMEdlrTkbpBYCbG2s1L9wKmU2+TDsRbGv+TZCjjt+vV7YuYO0P0s/UUmmL8ND0cG1cdUw
EPA15SWLObJbLWDkEEOkZ3r5xWCI92nQeCRm5LsnzsftS0y9+EH/3FpQbyORbPAeY7Bd5J45wscQ
WUw4kLYsx7kQ2ASWVBND6gd27IYVJqjHvBcqbj3dcXMBqKkXcMX0U8eI73A1iReL8oS3S+5yZW3L
Ltmt1OxiuT5HAD/B/CVCP47lVcnDtvNw/a31KoZw5rT+IOIppaC7uCpAccNt4OAG510UHCav0C7x
fV4xRGyIeiRc/l6SWCuPjwgu/CMOqs0LTw0259IxL8ClXU1up3tGDrTRsgzSfQxEnBgt7XRcsxaN
JvkB/mlpUavG3BvuEw+c34m2S/XQf8APBNAdyAyE5/H3gMZYxgaPu6y8V2R/4FCqrH8cMYcxVz4o
XpkXKurdx/Jh3Eufa9fEOZhBoZWKyk2T+ewrg+4lSLa/hsn8LMfehd7FrD4u6kiFZpYerruw+2u8
Kpn8jKJNetCHX4eexvIT0DraHjhIAw2fNdkNi3HHEKtUE1oMKP1RwFNX/Kw9PyC2rYJo8JgBq0f5
1Q4iwj3khTs4kXWef46hZEkava/gJ4XRngY=
`pragma protect end_protected
