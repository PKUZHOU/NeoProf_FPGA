`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
nYNXORRPP+c7jMSNT00LtU0qWwu1oYpWUqut1YyrgNWXPtyHtZueAeTFHfIxbdZ1
3G8ns9AvjrIfCDpQYIUekGrkVhyJ8V3IVfzRzIpwX4mGsIN9Nbobm9CgeGfOwT8R
aSO6zDa5XV0plkG/vp0hMnLUa3Ft3sYBN3DwmVs8oMk=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6976), data_block
Wb8FtYPh5N0llKqlvOrchXzF3kk3lCHJFz/TPgSDxV7/s55BzwFw8A6NxhRNEjH2
SRR5UBqM9KZxfMRfHOAnXOaiyDiItiAi7BJWu2JBb9Z6i9IfsJRLVg0DeSQ2RVVJ
BYWJk1y7r2BbImMtwy75dH4wQZccTG/Orr1dtSF53E6iy1Ill33wSVdKvaUlyOjt
m4ZCYJVN/krW6TpyVps4o+ac7m2wnedRcwMeSOV6G0RgqmpxFfWiTFGmUS7hungx
FyQQTf5+EBRLlt77GrdahXzZ/KFvy+3oTz0ja1OKkRlxs+bEriTkrGnnCgFWE9i4
lr7MrKgas708TcJnbA5bEtzk/xxe3B5d884K44A3oDmr7qiAYXbqUW6QfgcueZyM
SQCcJxPMJJex2OUSg9upocHmCH4XyatWIGFe+paAyteWgEB6EuD7gnYUYY+qb8V1
5HsMf7ivem3r8FOiyEC2T221KPm4dIs9F2m5mbk9TF4nVJvqJCMADxU3ABjGHBaw
0our3awLvZMp47eGATRU+f0x898JOYfDCm/S+cI/dlKIlrflOZacb8FFyaLI//cl
IPhl+2Xq+DlKKA0yX4EfeLT3tvqYAyjfb1ByZ/rF/SgS7JXVw1DAHUBvV0JWPNhs
ph0afQPTYlpv8L3ZR0PRVU/fvE/31Djd4F3g0P4DRZFNkMYE0MoAPdSpXFMKdblb
xFAhc9HYthCyekyVgDSQhJlAlUnsl48G3BMBkSMyOkmPKymKb1n9/MaiP5Pq1xmu
Dp5OnStnKT8gIfd2H9PxuEaOiYej7uaSOJQwTaU63mxQh8E0xSjK9nwMQPOKplTp
w4KnQAyzMnqJNfUJKiPpnUv1wLmt5HbEMPKFqnhcDV/DmqTF4AD5Y4MXfFSyv+f7
MJqm5q0Y40uGIoBLz7CpYWhsIV8IhIX7C/nUshvp1FT1QJ1t8WKd+W+pEsmoryBw
pM4/nYlHErdZOVb4yWLu2rT7m4OekgrXTnaF5Dam3f+8FgcyNL86BMKYcpeGvQi6
75lK1MNPOm/ZvYwmw/vNte9LtR0wjw8D4ZroGPrPg8afZwZfBdlL74BRhPA5ZKIs
KF//7NuHturT6VMs4YutuRYrk65o4tzACyoBtuGjZ3w6NknTgdrViYJ2erSebJJX
IhR+q0ZZIGR9F+aDocdBHxAE9NrsXWEC/XYDIIHQaO/ZuD11dJdYJpMj3gRqHSX/
1/460z1jijNPqDnUTF2Odagzhuj8z43TvFTaH+6nrrTNYJuMI9UiILyEzFCWhkar
k7v4Q2BQdI4kUoB6bSbh/Ga3mkO4pWa6MXqxra1ToKGRP72fXbVhz+F0k08+9scM
CS1IaIQDal11FMW0naB+KnqvV4ZDxJ8vhKz8nlwaUSllkcchgC4E84m7CEBHFYQM
am9Dq+Igc2QDxF1NRUlu+F44OuzgiSiR3If11/RW2d2IXhgcEiAFIB119ux1MxML
g4AshMe8MRyYzLvbqyy8yBTztZO7IdvwpS9lpSXVwz48g5rnpHBDWfDNSYSe1Y7p
PPETR2AHVXcj4nO8OHonYG81rr9hqcFI3zOHdofUanYt+MI6qMJ9AMwecRXhSeQx
GdbSYATExcvRzpVEY2BNcUh/e+HPOhW1ldYAyeNL2YpfhhsXEczKA7Cm5w/vlDWs
4B6F/PYnuPD9bxj0qm6Ro8fnWn2Np8hSXQdr3FRqnWftX6K+2iAPShu/Nsb+sExD
A3eDhdGN8/+h/7DOxS5n5Vo+Pk52vsL5XCLSzN/gjl3zTlf+gCod/kNoG19SyLZD
w2WvFxj0tS2Q3SMkWufPKvvWfEtJp/7fK3AxlO2jF6kOhExJjAB4MGcadZi81blw
ARMWCksc5CvxGBQnaaBEHVJGm6MrFP8S5XMFrwFe959CyFk4GfGsjEduq+22FUyo
Vz3SelYCkqBF2TI5ZWUmMOwym6x+SENfIghAStdhabQRgSBKvlVDBk4O48tfLSRJ
DVeaVli5JeU8aMHp0FKOETx/dXg8XiNLHBzmiYNV6ywF6M+BNzfTf6NUsjuxCXvR
xt0er5RBfzzm92IhwwLUElgWNI44Wku7648xDc0KAa9NuZPwzljoYelIEmYpCdWT
aVAasgrklMJnrgAZ8iCuNI/clxo/tIDFlsADYD3GH2qP29xI0o+yRgqXDhwXqWZF
5pJVUkBiZAOJWT5UCFc/W5korV4KWHG1YF96PNDSLTw1WOm7D4JqEmmYydxaFFT0
/JWpBgjkJ1Rnjx7mIb6zO8Krg4cMgk0GMw/g07Rz6zZMoX3awN0q3swpdtAztt3+
0/Oucmyx+/HLJH72Bspm6T099A/+70HR8dGUVuerWCyEVubnWu7Wh7GpJTuESuvv
PVkMaekc5eg7M1ViXYaNBVrc6FQK9QQifIttXJE/iICrrW9NFf8w8gdgdLVd4R3L
OobN3QQXs4LzLXqFewC3l3C/o8zxRHMdyEndMggOi+ukSDhOr6vdRTKN6pLL726i
IPwnifEKam6i8JFnA7Z0pvrf1o6p0nB/UBXX3D/doCaWzzmYGbjpW0czNaFvHMyg
3gi3h9Zz+FjII3/XwkH+8UhglAIOJmyFwBm/VS0NvrYRg0rhk78zM318UitxWCZb
6L86NRmhuZ7+U9mmVwTcVeRkUCsDM177j/C9EbSVObSPXLhsBFTQT1y21fBLtIYG
N5HRW9lw0V29xKIbBG9+9EYlgRY/GCP8F01sOj+Xtbr6foshoTkyV4bUQTw7VHtU
FvS9jpF+dUjsPpad2RzRpl23ARMoKLzaQCdHrJgF9R8yf4SdzNaYDNx8bNZHJas6
kh9UfvO229dLdeeZHVQwB29hgdcD0Yag3qcSy/V62OqXMvFiUjH4Au7aRongoeOJ
SRdZVFuh5ViUZpZz+PsFl9zZ26SLfajdA/oOQVFO5zdEMpjWDVc8JGCWh/P1+2Fy
CDlWeCoTDSrkASOdQRxi1CVCrkS28sre/w81UqIrNI+q7IpEZWtCXDWH7vJcH9FS
9ldSW1LVIE/ZCos7RSWjzkM6BwVx1A0tC3Vwii+V1v/Ve6GfsRoMblgCpz62eAVc
jQI8jyLhWmldMFiR2lSn/ddOx8srIzOWMqpeha5We62MIbNhe9ADZpSqPanXAqVa
1fR+rUmRCO3MhK0hTRp6HO/xFjqRuzs5O4xx4I2U0o7qEHmmwzS6RvpdxP4lqb8q
VEpaXx7QFnv+zvTQp6H7tgCazs4qayEVOH4kz3G7nitkwMBpvjygtfU6W1S5t4xk
0UopfH5uVeHd3oNlP2t0CJMggICwh1VWAniabWGlKtQQF+EcE597pDFDD7kSaghJ
W4vQ2K5LwSySyyldF2BvG8gUdEmIydFVt1TCTgUbCMDho/bvAojwKg2qTEraZxLu
qsJAU6zL/Bcnneyk9jA8mxPh31kuB3gnOurMjF+Ky+Vo1NZz0tr6YJWgAddKAmQ4
VFKMi0rl69ST0pBeykfjG8/3bmEGPOZ0ZC77JKDuiCs7sguECv/Bo2gqg6jdbXds
jiJdnvmxjBQtI+oO/WQAhDcLdKPofmN/YYuuaOIQUX41wvaaanLyLxSWX6HY4HMx
djrGsEZq2bAlFtqnq7YhYW+ct9nNxwR7ODVAMg/lP9FFj0+5rcEqp6j6aur4solg
uzKItEw060yXwEiBBXs/tUCoens2cGE6K8fHY09oJEg/ZXpbIY5xsfVKq/98zoNp
XoHL8R2CbMfn7Oq4ocygAIn6Qj33kUtqH0BSOSPTed3+/ZSQy5LHtroSLGpSxnUo
8Z2nDKDZneLIHGSwmYeJErklWNry4yVA8WNfpM3g9+pLggwejkI4mFnPlLWXol90
5/BH5eT3cDnelp41l1LHzq/F1MzRzBl+QPBRq+3fMUHOnFTwtSNvpG6pLVvnEgrG
T7jN5ovDAAkDIPle7efL03XaI7PdIUtlSc18EhkPjtV8h5p3g3SMhqjq5/b7/FNM
vdPvyf/v3mUi8Hq0IK1MEzOhHXGKt+TkvtGBDAPtaRxNk/cYXhJIVCnvza+q3WKY
SiYD5ext0nzZsqG8zNFkoeW9iyT3M3NxkilpeBVmkyiX5Z8vOx0Wz60FJ6Eazi+V
nhOEmSm7kX/BlrWTqiYcUWxSBZ7AGF7kVbELgzQrRaNwkrNE0BfY2gXUryJmFNVY
JLOQ2WM+v2SEdOwEMCa5Ih+N5oSQCTMsVTNww6UOnAqMeVmaJaO4JrjBze4ORl1n
GMga0pepB4IMMQ2MuOV0zn1MQdifF75Z1hF3mVIxU/CSCNX0xTtZd5VrAJ2ADnKq
e5z0RHhytPkkwzGeBTgr7F/iZn69ac4Pg+lkH6ha37L3HDcy93/VeF/8aXNYYbvu
vVI1TVJcQ9P4W8Kh0XWe4FvhXzDlk0ogHtBj87/UfOe9oJBQ6Bzqv6d+58pyB16A
/li82DXhmpk+n22cN/pM453f2gu8SM8M16GWoZLmBGolzye2usVpi2B1LrFr4qJt
0rE93AyVHtaJiJwCkMtx4NQuASkAY5xUJqjAkNp57QoALfI63396chSwxE5cxHL4
c5kR8fBX8W1NjRwqTgV2gQt1S/VbtrkWT4Z+Gx7TUCP6w81WTt7pSjZ6M763i9Sf
x8LxvzdTTPkPwrdF2sy3Xfzs3+vtNWZTIkkokAZ6UIU0BbxXV0UQrwE84VTmh6Nc
Xray9vi3MHAiFmBanC6VLQqFYiLk8+xduYRHaluqrv/J0Ioqg35vD8vLesVFEzjN
ZHHPsnSNhUr9adaU9+Jc/mP+n9Y5j5pMaza0LMq0G2QHDCDLzguTWsx1p2jN0AuG
Yn9hiUrFygxUjvg2+YKqWfxLksp4uvfT8HBBONOgo2lrf9V12BRp/rFFOQ8qmwoH
1GqdcqqfkgGrL0YBVZoHTS4z4jWwgfeUz2x/XFTdELwAOu6eQTuuYcdK5+Qqd7sv
eCGTxCOF8PTTzyyYYOUXi9RQm8bLWsjpC1AqRFk8vdUitc5ZFJGt69GPxCzRh6X9
c5HMt3T2gavU1R1Fiuj4W6S9Faw05chZ4/qPsb7TpTgejEpmy+2HIjqu1xORd+WH
tB7YsILjFyrbbvykLywlLIDSWfttOMkHT40pYUlyDdy1nRPsTvWMKE/UgCCjHG0u
hy68D9rWByJuyogdMcnRt3sXRKQriLSgg7UZOzzPKLLdR2wIk1Dc0Ld78VTUyWeI
8l83wGSOOHELiMoZ5I/9QFBnpy0aUWKbBdH1/DI4jeGkZrIvJMfRcQ89SZRaIx5z
5luuCsyTwwLOQPkqc6J5qUQvqlgX39Tpp1/TM+832mMDqKZHxp0I6/Fdh/WWCjVm
000Dz2WzttTsOUzRh8+WlE1FJgIo4CCRxUmErSE4NEKPlSl6LFY3u/z80qS4L9/2
nQEsWEmYlsAGonRNpXRVkzgtA227y4Uqtcjeh5xnQJOnHG0xIEmlooOZ7A1UK249
bjDmoF+8gfjm9S3LkB1Yx55ePQOzMReR9qnpVoMYWvslrcklP2/bk1xlk00v0bZD
EazmOS/XVcg/Xz5EF1Z4G2cs6kN7JCsZmBeXiwfcaA8jVl/MNmOz12T1BYvxy2ku
03nf+4aOh71+5Hm52/iWmw+nKAjLd+szGQIgUvPJLpTjgMTsvrhnqTN7jjOIVdJ6
sau4XiwC64yfXvNQub4t4wwfoTb4MhDakRShJaB/pCnH3OlK5D+N+16Z6puWzEUW
MnciA8WvOl5YCh19xUucBgSNXOr5N91qvIrOuLe9vgrX3AUg3fOoZj6M8T2CSBc6
Hgar/kfRINx5opZU2Y41TGGxXRayo0zMaOb6kj2yus3oBrlQVNYpyLsgF7CWLioc
ChFn3CxlVG9X6prE2+fhzpctEGHwUDBLHe9GRSluEnvpeldYBU+4TW4wscyKEgFz
qLFYCYDPyLI9DIPM9i+x3ewgwTSSAV/7XueoBYIRu9HSNwU3tI+iUTryy5v2vcuW
eIannyHiFChY8x5kN+F2YlF82B/HCSIQjSMLQAB+h7Y8hodlIuCNWjUiira2f7pE
LnE5SnzfIWG7aboqN/dMTxYGAKAdL8pG/Pf72LLRAHaBGBlC9CwF52pjJ3/cwk2r
YSMVIClw13pTqvLUFt0dStqnh9dm6nGv+do26stg5JYY7Dv/bugyX5RvoK2zxmLW
7WPDqeG320fYQm3kxfcMQLR+QUCaNFEFG1oC3+y53Z61KLL8BKUIRKRifXjm3EfZ
v4ArsWvttxhflZVCWthBDdNhwQnzEmzv3Lfun/7+5EOSr0FGbQMerYCLwpPmX4Ng
pgBHXf1sHM88uTDtvN4AzvUdL8F0MDx3E1qmom37zRmZTdqHPG3E0r1IlQown18g
Yrd26X9x+3aoxfeu/WeIoaVYYBjiGnzNGToayo5aJvpDhUuckQ2nfGwfhggW8eo6
JHZJ9AoZB36/E275LpPao6Vp6kK52ujS3d0NScFnhwL154gQYDo7r1nVw7aYo0j5
lxwAUePeiqPM5LwLjbklzU1Rr2ARwmw8HzpqHRM/CS9ry+U5M0jlfztj9kSiL2wb
/Qz8gQQhtaiNhKMZtgzuORqs5TGh2dPda1076JjN9jaZOQfNyc9BnfghcZ59HGcD
iG1nN3FUTncaC227dxgOSckaHPZjdPSJkfRZyDOUcQatlFvzcovUIB9lL4KHTbXV
tVKnMxbZeQyL9RKN0g5Zthvz/gelQhqztw2TgLRSV7VlP2jlbPZYCitp4WkRDJp7
AwOD2VbaahjFrdVQmlJlkRLdU++o/RSmuoxOQa6UENGeKm5TBq+d28OEY3HdU623
0N2HTn53yLtgAMGzHm+tT/Y8OGEcf3Sv4EzuUTBN/x84JFYTPBnz21EYrecHElPj
cUZTX8BMZ2ImtCKY1AWPhok3Mkc7dsSZKJmta+hB34bmdkC9jmDtVKKB2IBdSsvj
6PwRsbYl16GUs1/d3z/frMLNy3k+4ASEDXnzEruRhbb6x9LSV1p+2K6WeO/y5vVi
kj2rSba1Xytjy9KUwadQ0JDsqs1KR8noa2E/j3pG0GIuknwPFnqRqnyJk+bH1vN3
io3FcRkoMDMgFAFVy+XZ5o6+ukRJ3btduh4vfB9eod1vK/zT1JrNw7estnknJU82
0sUgykp4k0p8/hX7fVt9dPo6hUYCBUIlz4ue5jdxON/7N9VSkSD3Iw2iGN+BGyQP
FgyimxMVxi/pg1m9nxKj9/AiW99wCyj+vOsrMuVAmpLDsduu1bGnKmJnF/GMoE6C
ZuoQEYDNpnk6UDjcpRfscxtXiPAiUhmHM7T2vQp6rGwQYnD3dS++WHglu1LVJbMM
J4JQ6kLmVvaiHZob9zeoa3nndZSjGguubB97vSfogW/fieG5VrSibIXpMhR8fwv9
SpIwv3gKZTIdkMTXZnLLNyjd2Oxj9Ws3w3lK77iZcD1l12gpmIiHJHF8vve4Oq/X
H3ptALhUgKuFlUiW0MfPdFJp5ri8F4qPB1SUZHJjgkJ6+erhwJwpHjM1FSHtqQZb
QeUZknUgNRpselUZ9OetQpV4kqhhhyDFXUh7mcw+edCXt1lob0Gcjh+3CI6OXBNa
2GJoGhrY8Bwwna0/vXRa5CE2s8pD4Ur6SrUpHnv+BF2c1VqcCSyrIex0Nbpxlnqo
Y7r8Bm5G8HzhrqiVEuW4+4eR7XIB9x3o4mRuIBQFao35WgOc1ptlHtnfAPQdDhIO
iah9Yz9Hvrulis2Kntnit5dbxRFRNqCgfw/pLjxanQifXbYTd+iPag6pouXT6xVX
mKixpdFlb6X4ILugNE4P4Jb0IB3E5MfzvB6BYQ9NOviSAPAPqOSfAMFsgzK5Jc+K
xI1agnr4cjjEM7BvtsGhvUZVMsNbpv5gnKBl849HCo90NYwUTCMN4Ebrcy9nRQfL
MIlK4Fr2Wt1qklIy8RYAJx7zGnjunfr3UR3X5wSn1xB4so/TZ+lsuS3iqz1VfT47
2zM/ZBTuhBq3KUliFhwfn8A+iJocPSRG4w0rOnnTdyzzrYYZmkdpXyX4jgB/B63C
Lr/KujE4i+/Gcrk7Qv+pSzYtjhcKbucV8FpZuPXc0F4DyNkjpo3Oyo318gYmIhNW
357E/y3h0OEnc/x3GAL/5W/mylTCT4v1biDBXJrCrx2qtUR4gVV9hrklBU8zjU4w
lG3/+9kSdXmhQUURxAyUsk9rpz8sTGXrhxSdyGOev8ZT8QlBBGQkPYbQSpW9VaVQ
S7S0VQx05jGV/f5unk5Mvg+y8PWPc4/dbkoMIy44R2kYV0QxJV3zaVBY7MYf0bZy
cBYnVJ/6peG3oN8izq2JfqjL3z5srfqS/SOIbJAEC4uaC22ju7zhKLsaVnrq4mmS
Dbh5c71WobFQGvh7q61RSJ071Y9DvXf0+CVa346jQBD+m1SX+E5c2v5XS7YKCyhK
W2vVNz/NYNZMuzrk34lve3F1YdEK+Z+DQW2MKrHSzlkp7t/GdM0/jPDJlLWyvsqI
1ZD0BgwL8btoEie2ZesQrjBWQmp186z34rRsaCKQuUAWZDv7Dm+txEhKPBoWbHZt
wWkQzclFfub2gg9tgpkdG/emkMpIOPIws7SVURljRiskZp2Yxzq0S7d9YMDlUk2R
wwVlpwn6KE95xkuuapWXb3IfcauitLdIVscpQyRWQzuvS3n4rQxBjv74NYASQppR
fgyLP+abCuqT41ZAMzjxOTGAEzTly/Fkm0CFlqIB09rfCFEtE5rgAZIWTTiOlYpJ
WIitqeXpNoHWs1A4KXXBksc6cvn6F4j5YvUq2+1nUEXrAD98DlQX7jzuivpQVqgp
/Cx8aE5cj0IusysMH6+UMSzadvqaLspSTy4FCZsY1AKZyFIQCRloGVaKzf/u1JVD
l33QM63mEENP402cZJaSUZ+DaM+tMzgyZt57Fx9O6WqCttYYhM+8/6PR4VTosRAi
rDWT5G3fkXnmhGLusuRIyzEvPQkEjjzeMHkCbCBVUljKXJSOH/edUJOP0E5HmBzc
NVeIslAR0B99E5Vz/J9eiyr6mNjALxeaw1ggOBHEuFUcEoyHShWNR5N1GQNHz9k/
kxq6XFOz04WUmsCtRu2zZHcNAo3xPFyl9Z8NzKkiG+8yrYJMNhUFS8YOv+3e/bHv
K5mikmmOw3faxTvUYxoyL1cfK28Wh6Nq1ms18/YnAM5HKlgYJr8CCWSUSy6P8WV5
4bcUc8F/dLVEx5/HBi5oxuxc01bK3gvmzW1grIz98e1nbBJQC7MAGGPrIV7xilFW
NDR7+xqN+lkgsL3ol46DCr3glPx5U/7BceM0WUQrP89BGuXNVbRiqVAa7mb+hg4u
W2I6GbsoFNmZ6v4T//ntTQ==
`pragma protect end_protected
