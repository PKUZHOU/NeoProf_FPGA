`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
jTAojb5b7p2kuUzafutqrJLkkOxB10LLdiA3WSQ4uwnC2Um9crN6BAC7rvaA+Zkm
LOb5q8FWNK+iSJcLgx3wSmMhVi1G4dbbLh3kDv8i+b4++ZCd/B/pOhbtb5ZjSSV/
AMAoSB8Q33YFHaui5bFBZnn19RxmjXpR6te8+9WccUE=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 28736), data_block
tMi6pmZbSqK5YHqGh1W3m2LNRZ+SQwk4gy9ZW3CgVwPKJzahLU+0UhpINfzC0S6H
WHl62piKWoHau2gqlQwLSygcabgxVTKgr1OQXMsOKkHxQKZVz4V9JJ7B+E8OQb0g
K12Co8suLvEyToCFrDEHHEUbDikjxv0tpXFPxBr0XogspZ0e2iYIyD3mhcVqgj7s
lCPU4ZSjXTATevv7kMg5irj6NXAaYo4hAIFKQUX9S1ETWB52KhbiWeASwgG4Jlul
fCTzv/23cqNZcd0Bg4zbvciqW1JHRedt8X4O9mB+seClbOHcQX4twqTwCt1iAZHQ
5T2OHrGUgAJKbDc/SgaTHlhStyw9CUac7N+eL9dYyks0cyK8dYcEbp6t0WXwZH3+
coMVsdvKfQKfeGPtpYh8OBdYw9jiSwmMy94AWfQ3Opdfm08tcDPuYuRvb+aksssP
j22yGkft1jlwsFKyJAASml09MjDWTIExRj8zXWJRVkWEhiYYmtmcnk9U24vMTq3O
FmFq/BTHWjHY3qgIVN22WEV82BRyRJF5c2Xr52/JIrqAi4JUP+/0Xiz2JM500fpC
p0/8oubGMzrAjd1DeyEDHG+bGw/+gpIad4hIS85zBduRMR8m7gP/52vObKwYSL47
WHWNX4/MDi2nKdXqwWNhijxLajynTI27inxzhv/tEqEJQ6WCPH3G5R3fUBysv4rn
7GPVnHMChmtN7KYJ42WjGShq57MXxbjRhuLsDoIHyMpo/YYervMRO5VmRXHF/guN
ER1wTUHNR4UoLIEtE91yuxG7BGJcBkTRXO2IjUxKo/SOsmm99gEAHL0n1pVB+uGa
t+eRXl4tHNohmQ7QkjM/qGb6Sa3ShJa6daHqVQ0bJKtEavQp+0tqswseoaPIvyRE
TzZwfOx3DNgBFyjtwM0bcvBoYq8En/cD5JJ9PU4kv6YSXm67v+gCbXzbOXGGjMxq
UaHfzAn56F+H0g6wNxqyJy7JzyFL5VjAfjyjk6HZfzN7G1RlOSGETFNVCTQB04bx
DhHljpMsf3Z1Sn2IoJC+QDvQFWJ33O0kFP+tS2jhMiP5Utb2m/4jQOP9SokkFdFu
opDMyH2q0YSXSaGFx6zzk9UeoFozeNFD7IeUS5PzKV2SX72SIMUjkQFtJP289F9I
Z1/Y+fHW0cMAW1Ok9YLgA0E0IqhLMfWf/hYSGHHi18U7SbzWEF2+nQ5Pu9fikZs6
hWPpbSxducHOrtEeCMVs0lBldFDfupqEn9J5CTNvLgpryJaYFAdyLjViXnJsIQIL
retVXvTOz4Y8ol57uX/dRYQ38T/0dxvRkNCaSzTpKMRaq28Ddp++9/MO8Zrj0i0/
jVG1yfdsVRJQ3t/1Zazxumjd0hvscZY7PZWhwTpDqu2h3VNxMgmR5S+XdhLXD0p5
BoNCbfBEpWodlcWd2yJV3bcCKNcyOpHeX/VFwSYZyYfXSkn91h0FE1CfpZ7rAAyP
yk+R1N3PdZmDeUCHVl6pQi0/i94DcAYdOUYkULG/Y82ZoyhqUIt9Mua6VVma819s
dYv9GaHCuTiWRoQpptmbcPyhErMpo+8POEMV7bJmg9MiEKsrfaj5Izsvha5BuXKD
8kkQLDTkEDYuAYLaDzTdHNvAppU9bMzhvJ68eD3w8N1BjNkLXIGIy1UBU/6w++xc
r1+TXFUQ+gB2wdyVg0BvM/03GhGHqVw+hhDEic8dxxPrgh8qW8k8OyvsB9ZSTH/C
k85fNaWmeif+MCQSZOcFx5iCG6gv2oHVXNUsGaahWlyPbb29TW76y3C+ELp3qtzR
QPX3dNCrUAEOLRgfYT4XmLqvQ10tX3F+yewG9EZ8yvC6QddzpKr6mGHs2exmBtIA
Glv8pkV5ZhxTkTIQUTRZu5ObhmpVDNnw+nT37W2A3WdUw21TATs4c0Rv+DZNQWy6
9D2yNbtSCGD/RaMl2y9NoSZm78ZGXvh3xhcabWgf70haLOkisX6UtXGtsX4KIqmM
yjltcdNY4igdPElV5k526GzBqXAP002RZzorF1/l5soQxQIE1l7lLSb77pucRc8r
6hj7Jo51WXTp0vhUeSqPgtNd3xiX6oFqEpMhKG1NRdKk7hZa9m1gZkRBYJINbtNv
BmhrQH8DKqHrMUEGOnqHh7kopkHYmpVbhQpmMRmJAHzcD8r+OOUZHRQyXtS9Mobr
sXf119I04QR82XYUrqU7gSQcJ/Md6Hq8vl9Pk9H8E7fdGOuQcIfO4mdZSkxpwk9i
e9fK/1ZxRnZhO4HqiB4WYfXlqgtNH4AYJti1RB2RDMEKI64nY5iNlS1x18DQdBDR
OXouSP0sffWbBvk/UafhB6HIvg1xW/Sk9NFakqi5cFD0J2h/aVHDZ1dkeyBsy9OV
55tvpf5uUAojtvIRf9EPX8jjjeix9pOKnVjrncIXYbeOAbi3m2YXT3eGCvilb1aQ
BL3kux9OaThGi1bEQNCGVYtiq2wuXoSctnOUgOe+mSOuGolZ6kSblvtjEnuy3kon
moicxx1gArqfhOEiHuaHT5/Ei+gYECo2f1qKQsMomrj/ueWBtySD63Vvqg6+CCgG
mXRsrk2Ir7CbTBHIwnmzDv7zoCw5rcQlgglkq7yyOWij3lpsNykTQreaNbp5/vP/
oXBsXw5u9cHK5nT3w+RL3Uu4q3fcT7UsDX0bHjO8FwYmJVWwtyzOJ2ma9N8egcHu
NehHyM10GI8BWTH43FeJ/UAuzOPQyWlWbl2XnhFK/Ini2Su7I192cAd4vS72N22P
+qrpADSURy+UnXKeALBFwLDk6Llh3oKty12fwhRFzf7NMiJsFnuR/O4Xwfwny42q
oLnnTkObxKQmikHVdMfFM1kxSNrNiXYhvOntNG0seTKsNm15W66wirAYmBEi6Vuf
QC0o/Yl2vZHCBz4pHHK9OQli6XgnjsPeIzXROcdVmJ/G9rZsYBqCst7WZYk/EP6Z
HAsdh1VQWZLbhI5pfLJYxjmXtBbEch9AIDY53lBLlawhWGWXy8j7LyU3uW/7H52u
If/v7eqFtFl+KLKH233Ubii7b5SiVq11yjk/dYp2fEo1Cg7T1PsD+V3ZqbKwOhjR
7D3w541McvKWvIoEdCFSzvFW2ihzFVrqpA0LC2NRfem0vCl7ZkcHj7Elr2rx0Jkl
Hpb27vIWcH6w0FhScgU32kdO6atzvu62Q8eHeWsRtCenyttuFnnk31QcVwBQCwtg
BC5Hicu7GqBUBxF8IVvWgQzErf+Ymt/nsqIxe4cQnDmyrmvnSagNuUMw5TaXT/g5
Amu+jIeeynYlX3OfdlSyKqtRuDTAvhR6Sn6xCnFzXDP0qGb+eoI+xXUOylp0gL9K
fJPYKR9t/0f0qBYpQEBGJr8gslR3E2E52Me0xzpEeLKw5CweqUFWB+FB4uvENkaH
GM0ub/HRk+/vdmqSNJY1Q41Q40kKhPz0lqNvDdMgVntxR7QyijXKnVTE0otW9F7m
DVAQasUzy/IWBkobXgpXPT/DLNCPAVJC4yz702J3YjZ1AGVoP05bHOESALORkJkR
07Ml2amZIsOz3OPQlGECVgSz2WzeljQrtRlBnopuCs3XLs4dEALLg2Jd1cMPp06T
PmwlToPjaW+5gEKyGDJAbXu1XCkZBmjXZP0ELxJsPpZlCss4MUjJskjLGU2jHMZX
6Qdbc05Zc1fYGaTXMEDOBj38ikHtBHD/DZR81SPPu5UOgaN7EI9nB8h+Nb+jXF9Q
6Ma5c+wviJREd15/UuuQN5WPUQ5rZFpk7XRf/OX6oFf35q9RwYATGfUI0hInmrGl
ijDjB2ECIYmCFJ7ginsAtSnJctL1Tb2pq2rGf32VGGPT7iS8bDNNNoecoKsLixXR
t0w3M6/e5Z58cl0iHGj6FUB8yQPtjcWzZsRLio+XZulBvNnvWMkECsZYwR4ppLDX
E80Mr7aOCxoLlFC1iRBjKoZ84RFi3XwlDPROCTonKeoUrcJTvVwE9nbNi24HJIO/
l/YK8X++gdVsBWOvzE8T7fOvx1M4W6xxDciUQM263Q8L7IiWTrQfNKfsTUZo4c+D
lib5x9PrTgkFDTwpgLvGfFYyA7xVOetqkg8wad69o4y/5wPBp4l5iSTqatPauBkH
RvDZL4twmGTrFYdKvOtP4KBQKoW8R+rS24ambcAssWugilp86XqAisi0gQEd5fql
p2KO+hFRcyGeTsy2BndfV0U7/IkC0g7pgoojHfvRnAFJYKeDRYXSYI5hGFc9R4D4
wKOeSc+us02BQCdYZuaSBkAj++nGLDuV3iqCwKC55RNlao+pyw4mB7Vb3QpnCT/K
lNcf9lDIrfrpIFM2FxaxRdm4YXqOYCg1/6IPxkPBgVkeL9WyxPdD9kgGxMM88gxe
JuQXPostsApsXVUYbOSSY/lz5PJcP0AcLNZAnUrjLZ9kCudm3xaYWreOU0qob6M7
N2zVHkoN3oe/qodG9SUiIyl+hwenQXwGh4YXw21pcK5WCumZpnisYEfziTbd+56+
3CVQH9i+Y0QF+nTcwi17LyrcmuL1LngpodHlnXAZwVTh2icfmUZ3ZxlOKNZle/Wj
4FiDUiw+57/LTSsHEuWWrFTw3wxzb3BuSR3AlnBhHSnaEAMi6//znEVUHwP1lHll
Rz+JqGrvTMHiymd70XuzEYa9eSJQTF7kkbOFTLBG+5wnTghg0ImYh6P4FtKficW5
cOiGvJuW9TY/M6KRW9K8Ypisl5OMk/ObqVW29wBUVMKfZjFy/JvMDuhKnvW2Tyv8
gR6NtEi3f/JRVivr2RhTublchljrxMTCTuchEIVvmdJpgQk5GtXSxHq+xDehtOPE
07VbeJiP1d+VKJcyJ5gjiJNw9Hbnx2kJUckK8CioWlQL5VCTPiVAvSTcvnAdOiot
SSI5ri9kHTMEyRDD383A7KMvpV0FVVD/nGVo4/vdlSXkaTzJm5zAM258uvarEFxS
tWk9r13ZSlXwMJ01vbHMiNVwgNj9Wfu7CWmo8v35LExYBwkgYqrwoJ5W0M/RWIQh
++ToqzDMFqOS9HZjZjE8LeuwECWA+qBgB5ug8ssBrqzbSQvieVb74f3W7P/lU36Q
qJ3fMPAK2jRVCqqS9wAAcnKVBfG2ePZ/ziOnD/ZoXTay83+RHZZcZabt3pW6tROr
zY09wIsV6udQMmQUle/MmHkcQZgeEWJRhOuCAO2gm5E0G+yy0jY/WGC7EFhyFNZH
oNNGA/2fLXqT0NDfw68l8jk405p8LaUwA1R1mNZVLhQOeOPLhfnwgwoVz/NOMUYe
Md0KEidaGiTBK2UfFmwI4UcYUvd/iqJIOpuurS+3AKoT7/jB5P0OWOjE+KgBvZ3O
my7YWonR0B8e8a8MIc2xivAMat6j3SoTaz17tDr6kuqmzwu7J0/8+cEfEzpoYFR1
ReBxB/RYwZxs/99a6Dz7Vf64v5LrVKZkQKPRlsuzK+R8SoZp4bYti/HPVs0e6eQj
nxJuFueehj2UlGO4ZDmH9N2dN70VWnsTAbb7dhJEXdLMM3paSnCJQWTDRcsrX2iz
2i3IXkO2MLvHcG/O1fU9IYoueK0S8LpanR4ZeMShOYqPi0WgFen2vBKDT5u5cLKW
UlD8xncCz4WNRoYLmfMQnC7k/Z4h2iS0lAy4yRZkueYqotPaMsgW0Lpp3d3xP/EK
RL04mPnKMGn8HIzy5BD9d0MiKqPcpXaBG5A4m/pPRWOU2gFI/e0ik/WExt1SBuo+
leBzvy2VtRW2j3XfSesRst2wIkHNt+zL8d88qip86KPOJkFFm+qjPryd+0paQv6v
NXcbDUzKWbXMb4HhdQ/chxhBvt6rhdGztT/POC3FeWIRUuSeMXPBxPfL5giyKt6u
MnDVzcpfQF4FU+V2cxIvwLPhNTRt/FQpA3k9WTENsxllMFolxS0YGByInXL0q5R/
Fy9imeMZYHKX0GC2+3EIhWet8hCxo1FXo7gV5OFTbfK4a76NYiqepSt1qdRfuvk1
/r0DpCOEmTTP1YuwDOBrLjMX0AC/vFoHWq1GH23wdO6uYttFIZVA95kNKsnVI+oV
kFlxhucmDPoxbiZS0FcR54PvUvcWPAHIDZpx3JeIYYRWjw4zDexsf0shZgPT6Jj3
K+7Oxpl/SXFPTt5ykEFHBUl0HodlzTTeGwyGfUzzwiIXJVe3A72QZnB+0U22ANai
pRyuwMqjFBCzis+uA4lxJxJ/JAwMiZtSN3K2tu20y49f1CVXfXdr+1fWsUjSCMZN
rhark246lcKX6Ue+r3eOAtkqAMGHhoX9Imjm+0Z54JEEilei3duxnSYiYwQ48t3+
NP27qPTuVLUBXWgs2XslwH+Tt/a/n5nMn8DPmz7utNTmczLu+zHVL5wkIFGF7BfW
uuWqcxOW3Ngh4wmC2XYr7Pl9qeEIu/I1pMWUeURmn4gu2Id8gxxm+jt72ml/UbAq
3tzBD6JmOR66v3iyq2IZodXh/yrflMAYbfSoGas3FrmhEmb/krjabI66jE94jIxA
hVyF7nAdBJvkIvv5UTYvsthvUMLyuYgn7ly+5QY2YBVthEbpXLuDoPTx7BN4RbSJ
db/5b4+3CCSr1Kl2WA527a01JfnrkH23KfMMLwIHhlsIrDjJCq14EPJGlZQOd6GQ
nPx61DyOY0GsAs4CSd6Ley9Gs2tBIqifZtp2XnvQ2f5eg0WQYiOVe6GhmiKroRTI
kQv/00/4v07l+ybuWftEVcz1UwMgcS87SE4ZcQegJPqbePogVg11p0w1S348kx6m
c5pibdkWxMeKMXYxS8UtbuFAfWdDxFOXNHcb1dc7Ceq5g46Xu8OvMa1Uimb9bube
gtH6e+9209ob5iutVak70mRHPV7iXxGPgUKUyMFzV3z+1m9MPaIUlZyPO1nNrJ6N
TaJ/OpdHhMfODU5iDa29IcNaDGXNP2Xr3zK1uu9vcJ5KUda9grNWDJdxvtjC5e+3
qh7iRe9EA/j7IFWryS1ClRYiY05I7xd5FeuAkfmd1nclyqbXweFPXNstIiA2kERj
xrM/o+HU7IJSkqxpCUpy8y/VW314VOZAW5C3PBkL8oC4pWx/qGvJnwosIuuJO50E
bATInes5h+dTtt3pXTK3BS/GAfW3XD5AtTd9/t2/6vbM8PR2/A82VgTJNCsh7thT
RwGusSJcVyZ7SMV9wIrDqH0Pq1At0aofCUyK/RjcS5dzaiwZOnBs75a6P5yiYQDL
VO+5hzJI9+YwpP+2cXJCIoPTDT3KJFB3uVNj5hfCvOT/rQ0pqowGI2hIKnSzMQWW
yvAGiaiguSnbREM2EmCs7/zYlFTOpe/2CDPZ/sidE+E1EGUag7Ec+OPI3ki12ofm
i1TyCu5Ae9on4qN2Rhba2LMfHneS+iz1qeMLwzxHfqh6x/SE2QRZIRemL2yHdn1q
5M6HElSwSE3HsSeAo0PC1aBFbwaMh8Q/H2ct2yUHyqM/tE4ZY3C9mvTO0xbkZSwI
egxlL+KvhEvKJqJOA5S0Jb/jip/24fgfa5F/CDAgCL87wZT0j9G86wlE3Bv15qwT
KxeZErLT5yWfx1X1arxq0lW1CXpPJaery+t7XXwA2TGzhqF9i2y6ltzE2Yhn7U1+
xwtIc/PUHOT+ES/MtlSFjEjGFCVMiVHQGRjsiLcsQ/f8fnTZw2c22K4SBnydeQ7D
3WRnMBPrie52FH+yS/JJT+AkLScIm3ZtTlVS47axbnna8NPYKGPsv81CEMn6Nmme
2HYf7EZsY7/OL6DyleoBzGVetrgv+1H8dXLKqQy62Z+fpHwKH7dTwgiS1XlgHa3c
RhnfzBMIymKpEgzdzUOWNZT+x+51oseUdLGpnrFmx2ekKFU39n+XZhpCn2qbkO6W
gL9XY9xYJqskirgjtfWDbxFiRaQYwCU9NpAqxo73Rn7xYkLYrOwuMc2EH2sZaX+K
LqzC5iAd7TTeGGFYKXWf7QO30nOCtEyiPtYL3xjAAUQRRZYlq+AJcy11RzKiWvl/
221N/3Gz4zAkLvlYrL76OsX1zmqTgwTn6YHXrDyD8nNK8nJ8zTTI4zJzdDqcv5kW
6xw0PZ6uR5Nswi5Su84HbPboVxf3hVDSkLKcef4TRQdwA0C8TOTRAyIM/ZGQpKnW
eO59TAK1R91sOoA5F4sldTwA/6XB6ZVJQsT7no2RkKZZnGTSDZnI5pvH/wYFClVA
fHkhLBmnjXEgpO+3beN5aZRV7Jg/99imv0/agDDOJgRWVaeYK1q9H5DNufmp6tW4
7mfIE8lYCxcNce30Vsk9qP9g+hAPGdKKl9sqfvrSliIwgyjhT9wS182WBpDed3yv
0ldL1r+d/9F31fad3lAgVjvETdPWCyYGY3bbdSJz5Vhj5JEzzt+F4gJ8PKg0nv7P
oyAMSSVeM6hPL82+dii64IHFxTrS91Ko8TTwYCYnFdqq7j52MZ17WeccOGAnYReH
au99Q3pHlutCWBvraCwzaGAsk/WOOUdnFXYwOt3ccl5HgtqorZV3LyzFyepYVau4
eEZ2Y9rp5iLr2xhlvEzJb3DzkfmLIWqwFLT1zPvzxUfqzi/Swq3GfMhAa0KU1FPq
c/4vV7oYwVeAIpfOO89atlvUwUJEPKUuqNmHxhNxfZsaSA/xN7J3iovWPGuWA9xs
CwXVf1YL3FQJZ1WMCrA/Nq8oVPgWROoLgh9xi062sJ3hV4784PVrhxz5L9VWb5PQ
8YU7bGbeQFxYb5pIySfr19cCeQIB9WxcLOUGx7g24hXWNveyO+3fQ/0KCCSI6mo/
p7Bb+Qy219WDq2VGgAhPt0XXeKQKtR6chTSmLjMCxIPzT2JT16Ct3tqXTNVWFGLD
y8SqDmzYOb8RQI5xOOCD25aeQdKKGDyp+GJCMvwuk+gXkYWBr5LbZWuV6nRWfQ3b
2vhG8Yk7vCkmPVDXIlZCIxiIHBW4McA0lYzuXSb4fAufRitKMaBirgVexXIsB8Tc
kjI+d42i8nZhRL6+hV4J4LiHBBXjoXQc86pGfMsK4jf23cYtoW+0PaWT6OlLZt9Q
c9s3ptnx6lYOM/6XFyfEVIQLSprZFONxTH29xOXpqNQsP+zuRr2gqA6hMgB6ZxLb
QWYYR8t5Ux+Xnzq6wy3qNdLlcTlFOQoBZ1Kk3TAgQXj0Crgswns/DCdr4k44SMsD
Tyj9gw/MkSA6lcdPK91lCsLiAIGMmw857MrBPHorwzgoXsJYIs6FDKbPYQ8hEHlZ
IWrkH7weRm7Dro3EgkMynu1n7hISfK6RfJYNu1U7jEd7AmgufowoMbxxRLncH11T
hf2m+Gnc+6IiTqai70IsjDpw4Huuv+pEHBlpyHhYBanUaqug0Gpx1E9PcfF9bwEr
a8FOaaWsmjyQsgogWim4x7RbSmKbYSXtg4rrA9OmYtuyHY/7nnaZpvIAZRLKjD8i
kMvNr8rl8V0zk6epBkMXCUH8QF9NaecPjVyGoHeII82vzUc94Dz6m+4B8g6IIh6k
amawzyGYaTjYiYGqhh07OnJavg0xSmxsw1QKjMXQCY6eCxU5HxASfGjh/1xALeVy
zaUBva/DiMCuUw96OW0oYOB2xczU6tzXXNC8nGniEIpy4P9/7SRSwtfbItsDkept
ftZ+BqbvKq0YnVgnHlk5ns925AyhGiwFfau7W8LiUtZZxqDK5U5wnx7GqUrmkonM
u6pni7pBF8tDkIDHoHfPBcuExUJVcFJkyox6GlPN9yZl9ph1p1x9zGQT2NU57oUP
xh9xjMephw2hRG7OuOJkubVvmOGI84r69Js7lZM0mTpZiBqOzdwrlJ+HTIqHf5om
gPAadq4lu0NRkeGqpkB/XxyRRGlJjUGZQMtAz5ryYGHpY6jAqlxoTLvJWzUt6I3n
4r2IOoef7eHSEJN4oW+lLVYnC7ybVa9vPkp26fBNRNHW61fVEXeef9xkwC6H6BJv
8xBXvp7W0JL7LseM1FNqP0Ju/fRfJTWTq86cBkNiCyavqGWReXK0IWiXDIbeU1uI
4j5F9VX/LjLcXYcfyvXUoxK9dFgD8bjsl+azba/5UDRe2umH7CmcTKXElpMwLNoS
ILOHOPbxfaJ4j7HK30AzoZpz0s2y3dk5uuTlsm4d1g7jz9fty1mB/t1byri5EGGM
UKWGwbkvOe6JQvLwImBoz8ny/3tG6IhZMyJMMRBrL3a3UyFSUQWrcAftUqqEswDv
FwoNGx8JSZznvhaR56ySZl/4VC4KuwRE4g3/u10xk78+aNm2z3sPW+/LXO4lHtAo
4AFRccKhD2GZ5VkECdLNgMxoxK56KaA09i/iK2pOuZYJffJ8r47O+R72n9MwnhnK
MeseAadVWAKqYxr/mMY6XBjOLEsmbFXaOa+UpyxnOOEH9+3cVVYuJ6HMb+y3ykqb
jcL2vql3mb8sfYLnj+gsyi5iMz/B+vvY5MYXbFt63Obo0NNOUBGTd4V32x4Ur+R9
WdHx7L4qhUc6WRqUrL2nP9WayKvT74HZ0TdztoJP1TtcjD1IMAFJQO+UAN0DFkjx
K0Yl5nL/qYkh31ihKC4shRuyYxNblzlcL7TBuVU0Aw+DIsbFv6FTV8nQCCOoQqVQ
Dydj76qF6pD+wOvSl9vZMsGfy+IAxbSxiqXVyJfG2RbC4IRyFgpjvzy83ghwa39o
7xCCmVt6tMje1d7MM7juqLkCWkvWi/yel07wli5lVynXDUjn0aKCH2mdpmsOZWEo
QHXlCz69DaEQd7p0Bf7nEgyDVJvPTkNSrGjX6489Q/wvTTcg/0v41aUcI8fgXO5q
aKgzpDHhr/foaGo6TxK8OSZ9oQQF8qarrhyA62ylO7bVdkj2Id+KQJAmuK2fHaWf
zX6wr4ZsSCma3SQfzf02KgFHyiUZwxP3yy568//oBx0/3s5c8csRrSzQzozMpQxp
2X0pOHccyDoKnbGJKjneqsvujEQyvqNaLfbz06xhN1wVMQsane8XnHw0IVbb/EqX
3vB3q1K2GiB46jVuBxaEAnk3r1qKV7CaKlkCmueKmIMF+7cbLlsFJrhXk+ZsNrA7
5r9ML0pLBKRmjCmtVDMEAMDJyAhArij7L4dJt6huxXcm4005wEH8olUbaL7kcKEE
oBwd2Co14dRwKXPnVCofzl0eZzEssgjm1gdTCk3C0eySRfRIDPi0R2HDoiPNe0ao
SelwGjLjqZjsQdp26Gvga5cslGdWtoVxbGd6Gj5fdaWlmcOS0Bhv28+Z3jCgFjIT
OT72cc83+TyQ/iB0o2eT1Qo3O14NovNynh3ZjJc6XPILEpAapnwx0n6Kp7nqvKaP
U9oeCxzJrme2i2GeVv3Lo6fOZr/zZA8O8POqFNoPd/eIlz2xmxfrf/1b/u2AE+JI
l2fMvYxMIym5b0YkcZqT9sIkzSBy0hvVHTqCw+Bk8anRo9nSygIFFwfkSoRVhRxI
wjH4QoAT4P6FCb/FPT6skgu51UOEG3cnOX1BJryuxOIb82u9uw03Lcr8ow4TB3TV
XmiCjvubL9fplj7jeuUUFfmBYs6B1hTptco/nPfT/62OEZRcg3FqyJ34sWKXmc09
TtHE9GzZ9VyXbKOnvdWn5eoTz9+2AvSfpCGPsDqmoTBI6j+2EhuyD4VKhIKUOWZV
MEd74jBMD8R8X+UZYGi7yD65/Y0j26UvVsjrqjd/18mx4lBvPbk8sO5r+h5Uc+Jw
f8wA7ix5lPrwcukHFRUrPhioB/lbCBqstJjwfrmQmDrJ2yzNvNOutKrMuoeMJNQW
XiOhnQOUhD3cxXPgyWxCK5Dj5fw43BGpHZcGoK5dXglXxTXSlAF8heYW2V8G9j+7
xkB0PL3jIbTcxHX7ru7XF3z2qnMwo61brR48Y6uqLDBlijTcW/hlP81dh+ai53mL
MjaFk0MWWBa7qG1ZNdobWZi2crQyjtZSPqo91GcuF0DtY+1qTVAS6wpzkjUxGW8z
lahHFl0PX8vgLzG7T8zFqdRiMLdFZmI8acHfsNmcfgdgP8IJfxro5mIfS0gtArxl
wIWx7aTS1xKsNuRafTEqXkMs7GRGknCdkktiP0JbcUqKLS8sq5XzWpYsZ8Pg6sTX
dSNYPHTdH56QZuTOxH5wmb6o6NmZu8AW3vmDM9BrZhQT4V46vThfrhG6HzaiH4oi
oFuM5W5DlW8vOXVCnUFZ2YK7SV6GnY+E0CX9GWgWiwS/nPQ6CP4LXlW4yA9yDhUW
Nyk+zwP2vvTEX/VC9e+U/D01Dv27WPO7HDoPDL0qz/HbEsFnjJRl61TEAX0lscqC
oXbxpmnO3c3l9lKbHRorRTKbAEIscrQyuTrQRzwQgmdtGWaPEwDGU7YnGIbvfT3G
9ZuyMKfhPS6wVpFBgD5oDtxgQZHvydH80cm3wKWkJ9buslLl5d38/PDggE0w4CP+
SkvgtZyIdi7Cq5+O1nUV1AjKslHm3qE1jiLU60ZQwOJU/SkLEy5CfdDOqn2BI8uK
tPRQ7eN1bXxAvP0yuPJMblAc/RzFLayBQI+2sB1ijO4YSUteVRA2+8U3WVNS/v9j
w+yvKF0vFy1vuNVg69FnhbXKdniccvcFTMKzCtbjtztJjShEWIN0iaYrJnuDlcem
RGSAwELVBFrHGT8PVzxsM6INIOLMo7vrKPQgIzAqEyOsP4Vlh+FKu7VOz1F/KcEi
ZHUVEKUQ3MuAkrfOwZi4ziNhHFg5q5dkD/mQ3njyoU3ACAejk4xmMF1RI6q8ZArA
dMT/y4LrPLngLGGCtTPwQ1jP7cl4M6S3ptAumeUBdf+kLkYlBG/EuwQS4lIn96Oj
3jHlvauivzSH1YS7VnTlX/dS5bbQF/R31l470XSGjGi+niF/ZQm28zS2WFS1MpRt
f+ZRDV7vbFRXgB9eLL1dEFY/n+VfuXxVn/3flmVTrT9BpPmHjIV9M8xCt9/1wpLw
L4TjE8djsmI/5XjoKsiMWLASc+LKfTEd1OJ5SDWmYR0/ZKimaWNvH/G9SvJUdQDr
tj0DxF+tFpqaD8hdzVr/aj9i33xq3aiAZkqsuXdiCWGPHesvT1U12Z4X6rACMv64
xMXss6c2PprrCeEeQi0bSrRjgdNqIYdEmgkVFWG1sMyYyHhee8msmtz0FTNFyswP
fEfkTRfx7n9MiR9x7xo17bel6IEEG4ww8rhjBF97KMmfGI6LjItbJgjBgQp6L9so
+b1Vh4QOgDlLjWnpgNgJ3fIIM72qyGz/D3OoXvnBAfS8YwLJSmG3OBk6mYwFjWNW
kqDYhb0516FmO+ICFfSuBQrS3ibPQSinLCv0jKExZRJDjKrreO2HTvkS9Gs7kj5Y
GTVivqbbR17gr6/+Ebrz2h5G4R9F2O1Mie7eh7bjq6P7gecdX42WMEI+8fIWHUX9
i5YoeId3kuEjx54Jkr5UULdq1OPJ5CYHuz49VZJK+UHZucdyXsivgNTmiGA6NZRh
8cQN68AO3w75/15AVCHJIMUH14DMD9hOqZQWej8rHd7azhPGEEp+eoABJg+XES1G
ckXQp09/rZE0xZKLZl0cjLUBruLF3E0vI7UjnBGu735lAKmPIyn2NrNN9QEuigvb
0mk9LzG3UUZrsq2UMEkqDPqnijxTsCX3H0fOHzrZUJgz8HNKiZVgV4+JJMY6buAr
AtTEL+8d2ZoDkOSU2KXPV0yg19c3pHsI3t1toIJoNxjdIkDdfcYosUb/9VaL2SkO
dHlQdA0VnAmrWivE1DLAJQ3pSLxJdAr1TPJtajTpTGezxbUluqVN/g8si/p1bePb
gQzAtDzKBLwxIFmhmRQnTozTSAzjYwCLIItRggm7bY9OfIQEQ5D1wnldPhV/zloj
HNZ3cJyf451p/Tq/yrqRUPyofW1VZ4LvogjS2rcvpA6sgGHkrrEGZv88AXNrmn5T
6JIpcVNezFartP8q2P8gIp3v//XhxWPV3o+cQSgJ1VO6Zae7l12cbmbZK2NtWEo6
H1/qhd/bvOPFn1SYLDomx/EK2wi8agkltCS6hz1a9GJXAHaLCMWvU5qvDufq52vU
n3030hLAux0dgOxCcR9pyvJ68dmTB2ZGdvcI2cAgqFDZ4EOJ+FDaIYo5GORW2dBD
/+e4tSLZz5dkwgtKfkYmujAfOB5NDOpq4RhJuQDh9/kSLA+9BpNGPaHzqzGEM3hO
J88/Nqyaop4M8Q2uAyNAka5lWwlj1ZCZaAcIBVvPYa9HMCiPPRdy/Gp0uBOmfItS
0/4FpJMZVw64Px+ozDYLZgKRBb+Li28AID++4TFo/BI7Nhsiyep67n/FGrhaf/dE
Wk8PKG2TH4a0tMA8VyU0NFw6cyHADU5G6/lNAQsGkX/FtciAEhQVkTNd1nIEEWGK
VGmpG7fGPiCCdjsoJIPdR4wPHOi7SrEQj+hb/Mo3bAk74g1mNSGQbYZc6ncuIIMw
40ktDRN6qq7rE8Qv0LBg12njB2ayc2fb5jVclB8cjxIAihoKYoVuv9R48tt67u/a
2MjrQGWn4bNMCu6qQoU8U226oJIr1ywo1SN5ifakcnnYEiOMHqlV7f3aQfcb2bd3
3lP6zxJ1lAQAxO6WjbCZnnVJss6DLcbHJeFSHFaDdikNbFqXuC1uXXtxU3yTe8ZN
D3kge79B3NMpHSzg8Mcyfd7oRSDAj0d1baZ7kAoYeF/b3cqTdWxkWz+n6ysddOl6
ZVaCkYZTmcMehJOEyhrSJcXHIqQF0AD6ol7Ks86V3MexsGHTsR0SurYQE3/cM7pd
2KnrWgHBwrTLkr6Y2SEb8bmWuNaS9xffddoB5JqbzHpU0DMvk84VCwcGscovHOGg
iR9Fhsf5VV6xkSinnsm9LI+udeb6MSnAXP68IOgtALnoPAuh4KuR4vVokXIyBxwJ
1Xg5C2Rxy613KlxTw4UBy3OgBNgK8so9TVNG6Zqk6zY0e1OJ9WK4ozXBxiz8LkWR
dpbsBXFo/enurR2YPgbZKdLO5oo5jHTL/Fixi6G41hrUgRAlX2XL8hHg6LtWtoBM
oedvryrSPEQ+8CTYuPKtRCCUhisxm5azfCCNFBvOly+x55u4hZori9CTSX7dArtH
gilXEmAqEjVgiSu5Qmac5h3BpExlmY9KqcjFqCykfETkO1hem+2PyynSz5BQpQPG
o4ioWI5cvgnVxThjj429RcD4ndiLXMD0ko/xHlip0sSwzMZS82UMY75VVwTMnqKo
xtSPsMzCx18WbFk7yQCd4dKiapHMBRSbdB4bJO1k+hKHQSy0G+mjky2l0gfaPcVh
k21SCHFuEBPy5Zkdb9cCvhHT7diHkKtef3XJnbGlc1YQvyQ4Z9fjCz5h+Yx+UB4e
TkfcWn45KS64V/CikPVqdt9I6HqyyHuMjAAc5ZO5K2ZhsqJ4j3fkfbHfZBBmpOcP
+AoGISUd8oEpPspxVrdJhiBKOCYYA/NxuhhkV0F80lXMFIn0FtWDRq41UqLt8z/Y
1eRcEzyxqLiJEuzIyzklZht0itJklu6nL6NkP2oxGAJ5o8S2MBJo9PNJ6g86Y3Ok
NC18PTjrtEtqFjrvNkyVnDFAmCBbxwlQMA3vxazZYsQOTc10lh3cUTeNq/CIc7qs
F0c3iwQE+l/YMHTgO590b0HKStAL2POEVYBwSJ6mfktob5MdXT54yqGJzOZINRpa
eXCUuRxWcWkg0sbpFzQc3/C0cGVPAKceRLEJPRobEJ9kGZ916Ftv9iDhZ4I5SmIm
ITfPWKIxTLOKjs8D16qeQWKizX28xds00RyfMYvnBwRexltzU2XpRfNtfMJ2YSEb
IT9doPAvx19kRfD7DuWalViTRjC+lPpgYxva8IjHh3gL+QsJ9vkMMVYFw5wd70Dr
RS4WR71YNhM57NsGyOYlNNRikNBCabAKA4zn2IiiMaPDOtuRiimk6s62ZGSHx+8n
hUnEK3/Y8RyYSyVF9Jb3GYfJqL6Q7sPdWxKKcDQLqsTnEzPZ2X8XNcjJmio8SVpO
o4y6fEbcu9z3mttLtZEWv0aeMlwjtrj08gkehBcjkGj8NilVgfzfvs/Z62BId4WR
xzCyJde/Opza/ZwqVLJeIKqngxo93j4lCJglxkmrI/OUJxJyGYdhUUOQx7uX/JK1
8+jZg1J1NTujmIewiUA78GTgd5pnZpgmVA8x6tUcQGOe+eKj80xzsDLfAo/gIKbt
ZUc4x4+BgV9EBX3g7i1QG7yETOT/Pd+FvfghIHpzMOiZHsWYyXWZKDd34uHiYUPW
8vSDHyPbK4crh4iHiVjYtYQtKXUNoqcCeNqTD3BZSFu0kGX6/vVwx2BE7wYA267s
vwyvgEuOY1PMrJ79W4xcCdR9dlSTTBq/IoSrd8a4mtLbHq9hy5ATdrZoY5ruLLc7
8Q37j94ceSyAwjFJk8VaFlPHD/w9GEAPGsikMJDpLRyNARgh78pwx5GLNC3vT+bd
dGJJ6BAEcHDlr6ntiOtM/v1AS8GX96JSn99Knvitd68mOxUZrmueh6NS6APU2TI3
WgcQ4j3Hx7klvMJRT/yV9a850KRjpCU92GHZrQ9m6PyirdMYQXtMhOzdVC76Hmj+
VNWtyyO+0kmu6hYwlWSO/oviLX/r/j52pYjTh7xEltRewILxAQdvMlyabR7wtfMb
Iyf+Dach9pDdrIN1THDDsXBGx6JK2TRzDSby/41xTD/VqNML9zfP4SiqbvbrK0AI
yAD4xiZBD5zY8LIRqaIWnhShD1z8GvvJlX1ze3G0tv/EZoVk1Z0eHqYIGgODTLn+
utudzu071oP9cwbAfoLEcbIyx5UNTyieZU4OoDmG6Xro+ieq1UfEwiG2strrVUTX
UP7rArypUWgtusIEhgHfo8SE6JudYHux7x6YRz3oPpoFoH4OZ/AnCWN8lb57ccp8
irOkZjDeD/fvAZxuD1tlYmE7BstD4aMdrnqUbwBKNGuyU4FvwLnEBGBguEzyHlge
BlbuL//GRmh+4YxYVZkeYfJ7KV++Mvp1CV3tnR8dB1sU5uJTXV426/tFkxB6N9pm
nMCwPkfEm3CaY+SbfyomAqXlvP+GJtIlWKaoyifWVMChHqIZRKclmjXUFj8dRILm
MWwfsZzBUj5M9VGdo/yshribiiqAm3onweT/M+xgl398m7nOrYiY1pj1E4TKOe2W
dLmMymwKYVkvYQi0V8rxuZ90DhZKWfJaYS3Ay6vREJFjqIsHxT3fEhK8Vu7FOPPD
uYt9pNMljNY2R6TtyotGWOlT2Mw3ANauRbTir8HP3ckWTuQaOU2I5nNVpRB+oOIo
QgIQ/VW9gKKTps8bUF0U1P+0JSWTMfxBhAX3gl+a9GHtTFxeAH6o6QnNCwzVHICt
qRvdGgpmeigvruLNuMcSdtiUYX8Pf9ntG+lMOHDctza0CZCPCVYU4ZX4gvSC+IbN
f55unoyRGsdr0cIoRgkIM95Da8wvFVe+mgSHwSm1A7HtfG0Cv/RVClS0rBne/qPX
KIeCVI/NMlK8O3cMQ9+vHWucwaZvRBXXi683RMrXLeLJmZfJj51lyZGGq2OKhy1+
LaBCnVjqVE6SJbYXZ/pZQtW7ofvxL6gkzUlfCYlXReojTmEmXHca2N/U7NVwKCBf
7zC31qT4omiduc94YIwvEp7l31iFMKHLD7iQpaOte89IModC3nXH0iwYArRF1EJy
3eVFGZz3ffKq024BK1eiiw/N4UvNUGQirnmnBerD9lvFBokF8Ovu9sX5NNZdZeRo
iml7KUiwOfReNNqTgV9I43xBMurgnYZoH8tndqf+R/cbx8PPFk8Z2u8uzuKBs+aF
5jmujB0zuRGNPjElN6jiRlrlWvfT+3lhqcPT1+vaxhvQ3DHUHmRzmlpFGAN4PaHs
8zm9HSWEQNsZjjYhRIDWOXEfULi8rUP4UIjIPhtfwicdm52OYRfTCGjBoCzm5V/X
hCPvHIA10rOHkuZEnxmDgggOvl1FyavXkJAJUl2t1rc6JlGNnWcjrSW//0H60nza
T2k2/v/NdgoqvwVmRlAem3xU9YmQvJZFtXYZergheZokH9Ektvx+cpwctp8uD9Ej
1tVmTNoLmVFnwJ/43+krNz6q4UVLs5fGRcMGgdbceHAKTCR6YBOFOYDxqB98flCm
1yEuD6IVoCLcAItiXbWASurgTdkaHZA/jZFaWkQHTjU+m3smw5Mr3rfVKp2cxg29
vhM4LaKL/Wa2eN358MhHzl07NIQMecOwKPHpvg49K7k8L3eue3Rv+aiouwZKlOrj
zZeyLlaEZrKiVZ06X6I5VvcDGTxLomApl9jaXpaI0YiW9CpNThj8nS5TT9Rqsbm5
jv0ZdqodLAk3Yv6GWiirjVPc43jCzPn9U30ihfC6UdBU2SyfIa5rS2odFZA4T+Rv
5ePE4SgNMlY3oUGosAhOz28394ivJFG6iGRPE60XHp7Jgk9P3412ZI2BqHYh9z4r
Kwvqnwy4nvZL4/ek8PRc7Ro2804LdJgKcJA6zhYXphkMsU/1hS12vXLALl1NDRex
MB/QLpLqzvJ3ccUlsWvfSjWFyq+ESuWpdtd2K/TmCh9YHRu0IMYRgM0haWR74/4o
sA2XggAuXypImlPr2AY8OlIxQujyrtK96ME+Jcb+RJ/X3hMUF3NaiKjztQ/qW1AJ
V9bYRMh9rm03eIstNaUsYb8Cu/BiTaE0fAK7eMIMvdVSc+71Op1QypDZU0NW1XSe
GcYyLN8nt5v+QKmnO2l7V1uhMDQy2g8A+Vj6Y+Zp13He+MrKVLPIv9YBkR1keob0
9ZST2LCxFty9u5b8lCPWqkf10j4zkiqvoQ/ZcB1tQTVftgbDUUsFYAcI40TxEk3I
m5euB8LL56opf1NRAIqUuJVvThOUU+pndW7aEMd2gSL5Z3TrRpnX9Xha7Awssn2s
XWxqE0ME4fjuXc02frfYVdkaaiF3EGcrzWDWow4h1o1v7uVirGMjIxwRZdrYDrXD
egEPklEI7TVawHI+zbJNqDryRxLLrnCiM3hzVL0rHZw5TzAwF5CdZymJil9NLatG
yTxGTc0m0OptSHvheZN1R6s+DrehBIih3pwu6CN9w8i0CqrTDnCPkGGRKXd9AYMo
SDuHAq93PmG9c/yB38o7yX6VTQTmwwHGYxGoa6WbEaWTKjOR38JiPJMNc3zeIcgS
GJeIAgL4sEwjvG5q6Ms9t201YvRJ9vf5ZsJlI23ncru+2CTVq939hvSUqOxZsVn/
7T745iBzHCs+9AOpkjvfluBOBIy+csA9FgfOylQtLSR7Sy+0MfCgAOe1rmGoMuCm
btYBmD4gMk3hPYD/oHwdhnbsDVMtWIxOOi45M4VmObmILWg96izyZG60xNQxYdhW
xB8zs5IEaoIU3ISmat3GF7X11wTndwA5KTj0No6DZ+u4VVb4aq2s8mZETbceDeD4
uD59mRAYXhroAORZCzZwr+mdXurb3HZYdd2IU4rSAHWgG04v6PMF4MZCGxCa7XZs
oQm3E3mq+8iE1WaUDFWo3fnVu9AHK4An1izgZoPSyGOyPA4ixwiEtk0rEhm2Da7F
NpYauQrtXEHSCEqfd3uG0PiPAUV40c2Kyh/O4XuwroDu0bgqTlc9dXq2ALIteFlR
4tkWIhQdwH4IXSWhXz6Ei7QI1KZpPHfX2zdSSEVQlpz/rsbdgxjcj8qfVAH9jN9z
eaRbbrebgYjyzm5ckSscWCLpmZxe5R3q6RGnbdyrp69SHpieaLXP1Fkkb5j/NEFI
rBb0HXSLLzfbVgamnYP6fDoX2wD1j4yGqvYC7AzZ+PpTaUR7sMsjI2/b+nkQvCf/
o9/0nYMGsOOHTMSOcwYt5MhsRQbi9THgK8uXAy5r3Ap0i4YxFU6uUzyD0k1zl6as
DJiDZw8ZYz9sgxBjOOLxBwDQNtzAJxsk47hlHeLaBTZSowrJ4M5qWAl6RR5SUoox
Z7maJdNzqem4l6k5Nm68WANKsks92IDDQBKxS34PfJVVxdF1/4BoDvTerGimDde2
siDrLpPdoVoMteYwjLiTpxl/tTP6WTzskBZQMGbB6FPscntlUvbqzvG2lpv0WZes
Q7ytkw/fbY3PqyeryVozZQLJwTaaKZQFr5C/ikS+6mRdAdUDNWIGtk3dsi3O0j66
MSKQMjVa5kebW5wY2yYWAi9hpnmGuOSuqxTDKfImqxauodaQVUdi+h9mf4/0Chtk
TQxzEn/DjYZJzXdv7/sv2iit1MOAwTDs/EqD4WgB2sE171rUI2ob6d6UAYxusYl3
cdkX/HCFWpxzktIoWD2MYL0WJJQDuk5pm4H1yn1IcLFmuAr9Pj0efzBc8SHFypxP
ARUws2FQVN5RDJo+f4KnBuM0VaGZ2mFNyQWplwuAyaAL2TqFebPgddnr9s6dmj4Z
9xMwonKvlOV9WSVq9tdSJXtQPuM1v6JgfKOMnJpOTfvBSAE83C4RDAp6he1D5bdY
eZOgwz1Vizx8wEQYn8GwToGiHdZ2TupQ2G7TDepMfQz/V7XOnbR/9HFUqiv4O2Rl
wPe98i6Vg61PqeP7W1/t0aqUWbVq0raJ3xROWcb9mqGOQukxZsPvDG3NXaSFnAOO
wmZjJTTbnI+yLo8FUBm/2hnyOY7qS42f2aQc4S2g6NiY8Ly1gMeK5em11zTozC5q
0qxMvGEp8YutLPQ5XcDTIrNF+MCw6cnyONAsa3QIwoDmoa9YUTMQ5VlopJSLc2GH
ezidltrYJkvdSLdl9HR5EiXoytwQ0E18nFkjsFXZBTMo7NJ21ByrsV4ebeLPuMta
bTf8PshnHhumUBQR0REHw1WbeKZAQzOMIIB6mXfrstIvlXbYrSJz27G1phdnTbM5
jR5qlVcSQQl1SUbxZukGXCnP6EtZBwmF0DxshDswqlLJFfbCbm5h6pSoYvE09idg
EtRGPwj+HYujBuzw2zPRIp6XskbLVE61ZMtC9uUb8CW+fJbDv2tsC4/tKTjTu79G
KVL4hsMIiys1kRb15Mgfu8ZTkiFxZIiqN9/C1BoFuBHFhO1/KE7+7Urk/jkXNOdf
bu+UCKdeHYdyvBCNMHCQQHm69SZXEA73zvAPyRTEtWlbx4xoG7LM5p7BWWNcj8Jo
+wpSpTf0tBP1YN5stiMEaYaS+kFEL4Wh7UZvuaK8W/bU4Haagg+azAMwwe/fNZa+
xhPmvPj73SIxc/lD1QNqpBuz6oWe69a7GO3dbIKq/CC+MfA41BmxsT8WmuKYLSq3
A3lsbuNF+h1lxFVRXfRLJgtkkuxe/rQoe/u5q+XNAVcctcVVHzpwJruD0uN1v4Q/
tPLUsb8+wGZyjM4JoJLQqrZt1LarLTsjXfHFUA7M5h1ILJR26DjHLK+NxjNDs0g5
pdUuqHqaEuwm5qVMY4+qmzOkrID7pH9HQzDbb8lKbKaJ0nKji15H/D8ay2ywq6nN
g9g1qZpWiuQGEqK0uK/N/DelfeRYzJoCi7sQFut5qYVagaKyJ7szc/xSN5TGl+UL
ARbrcEfRgs8b8fPgah7DIPFuIs8SYSuzzEuz5JjkMTPhnLCO3s2rQQKVMBEF30/B
MuJkmitZKZEu6s2AfkQlqU442hMo/PeEGw99xprj3FAMSEHIcMPNxStpeSPRuEP2
Vdnq8AfjolVRTdeEn6raDpvbv7OzOONUq9kf3EVb8L3UHktpfeYXzk7U6kjjjaYy
113rcD02xbd95MrHKf3CvxEfvWnNIs6ZnA689KT4NV1fvG/OI4vmEH3nZmEqkTNb
cetd68xz2o/n9tl1SHpoYdc6aJZDvQaCvgxdhtLG//sVTaKy7vEPG+QPbSJ2xgLl
IIpFkZdjIzKIcLVWZitNluqDm1YiF0QiaI15Ch7BVotuTY1fLwIuwSbwUsOTtnC2
jOLNObw8RXwgN7J5qgnLrLn6VaxLoFo36adA6pLvTaVQUABbIvO+MBlOL5jL2mW7
3VHcz5X9zuO8Il7XOTAOheYnJcbsGi7tJPj7cnGNy6nCEq2Ru/ttrmO7v3qL2GFf
dgzFEd1k4O1BDtvs5fldoCvorgUYRw7jpq0m5SniedtG2AvGm9sGEpd1qR14hxA8
N/mfbpMq1AQMBXXqTs8kjTh+AvkBSa0/FC36PQ35Uiqm64xtBk+6noj5iCpPO2q1
22uevK7sczhUC7RGwqxKrH19YSZ4wVfnz4ymcsEzPiuUgcuWizSPnPtUX6xTtQUK
Pkg/NELTNCctJv+QAv5YoSQ/eiiOt6IwsBQECfzi0eOBO0teHK0e21Uiihf6myfD
QEoEvqD/9Q088yZ5Lzt6hCdCyoDVZU3wpr1UxfG6vBbJ8u5MZyOYKPbMjyNdadOX
+hwj2DAOeuGFJI9Tk+0TH3F/5Jot+ha5qSzntWQq1Pu3DnVFObkar7wTD38k1LO0
kKdfvWz37u+b8lZS1Lq0jakxJDd5iJr/9yZJmr/0JosmMfR7KQyNN1d99/G2uB5P
HmlVFXwGrLW3wCigNHaGvPpf+s6Pby821VqF4zS4GgJDakPPG+pO7qOtT9WIhpvX
5Nj0Q4Kw6ypz8cHghzXfeoyWz7ujMgC2nVixMnLwfuQB+dMba7Er61LCXgtJygvf
QmeCBCzIdJ0AUKXGSRHv4zdg5lBhnst9Yvn8IOlivn1KXP2C1XLrhps8UXBWOLvT
Qx23BPW+QTEvqIvIqiHPtT3A2oWPtNNlDCWe8FTGiMpkWGvZxnN1IEmKncwmVYCv
sO/XXrUqZ8UyQ8BfUaX9mUVrUXE4ouuqGHDSGe1TuXRNj3qoYtFfus87Wqhg5vde
fggGY15wH3CUSdvZONKo2oUUE7swjSwy0I/ikG+T24OjS/fAX7O9+e+ckkct95IB
pTBmswLMsDhLBw0cCFBFsvuEF9UIYQF5ERPw6jcngivaxSfpKCshMriN1zOMoD+O
7NkdX5NykTVMthRbrn1tntH8vQHGfbqSAwlYlLiXhroc60cL3aXFAvWitQMHHVXH
/gXFKSed7CkCPi+MjYmylU/2AIMfObF4etSU5mM8iiW3r94eHbWDtZIFiFe9yB/j
e24wTeZjEW2d2Zp1zPhjbHAzohfDfaGD8UFQbyOQAjL7iKlHbLtyj5sPPL8bbToD
yY/TYeYZ2CSLFjNVtq5+MaR0noxtkXVGBpvCAH/NMoEx8pG8lRDSPcr3lcol/oqk
5zUVD140PN0h0aWMxz+T6YS80tJ+O+UDbylmDXfVRkzLqq0I0KdG5XX99TJM4JN6
hCHOs2yKaZz46qlhBa+zRhANguxciNYbo2ScpzonC1gy5XDlONBg0ZwriuNSXTeU
HWL9UYmaoLtgSXFivbKVveRG/PbUKWUaIyHQS1u5JatHhLV+FGF8XOEMZbAOVKKx
eFP4aNg4lNL/5PMJH7TCrbLnYhgO7F6bkhH8PQmrCwgl0/gEodtaVGKu4FVwxp3k
4OJJSv2p6Y5ZlogPwlOu07RGPTWaM9kwONDFh48264IXhdxFionWstAeKYsjZpkA
dKvRps5o0d5k8lZQjmfX6a5ex8xaAtqLXvrLIy/nZ9IGCieyy13GYC8g6ehXngEA
uQXCRRlJu6vXGL/xL7vQRZAPopncjqSbHoA1suM4ukO8cnY4C6X/qaz+D4dw105+
iegXREPbrzkQX7jHrNOMlqEgA8cRJpYPaDnxK/twcXmfKVrYm+DwRO5zGixpvE1k
ko1L09IKuWFw+6UcErto/Xp9JY8tqXY4Pk90NWrLbPv55U+8+zMbkudCgOg0wDTY
3ntzoIJPjBGhHVRPSMn4Fa1dpu7a+Omcl5bSOKF/4wEXxXM0Gc+wY4WaCQYrNDFD
ymU0ZgsKBL22u+1smbxRLoMtBW4RCUMJGDLRzfYb7V6eU+beTJtqt1vHF00repkl
v8Uot0l7CQBc1Qcw1J9m7tgmYqXQwI9fdxqeLpxEVycXeWPETSpfF9NroPGp/syQ
koRVGIShiEzYUE9IL6EPGOjKlKNI0lROUO87GdRnaCH4KhPPXOlk0hDsJlv889do
E/0PKsdb4FN2eYMTgthDKPCC3WvQgbVZrQ2NYvWlzYt798fvhvdNoGXaGba4RUBD
AN9Xth9QDqKLh6hi+ODtnLgj/2yJrXpGkTq1MndlmOTxngq2pUDl1UeGrlExI8F5
ewJd+UzoIDSUweWzmHi/u/6/il5EQ/P60j0ZEX9sOS75zKvz3SWl8ax2t2oPSFdG
3OYZBCg1+Zt3bPOwktP2oZMfEEX4v2U9nxyrw+hHdCP5rNDoxS6C5z/gf0yuNT2d
zVceFTaZsUaAd5r71ApcspZzoJaSxYIYkKfWYVO1E5Dm15f3rftqCUPTAZQ74dmm
EgTWyHw/1szpRzJu4Kr+WjWYoYpj6Te/TAUBdFSCDbndO/LdU9CKi0DTut0brnFs
eKF4XAg86plzfl21vqjNJlsmn/sb648A2YiNngyMLV8tksDy18wP/AyIWokMVUHN
j/kcGqHMZNlVU3CLKLSe09yt+FusOGmjUahG3i/vPezs+X4Iiptsv6n4wjTwfIMV
xGEgqFIiW1fea+gI/1HKwNsypv63RTJ1Zsm6nj7QYIS+J8TgWkb/SDUBe8s5ecPR
CgXg1FJ2nMe5Siv9yN6akEtLfxdm7BlHSevlT+X4lP7IQKVcdzAslW3CCslkz6JT
ca4Bsm4iRR+1r6tDUHrHv8UmFeU6M1oCc1n/L7RsusyC8a//eElY8C7/7ruw2pEQ
oyUJhurJRdU9EBAXE480lhMCUv8Qdj/YjQ16J7KhWxjwvp7Hkpbe66LwrPWO7tmB
aiNtXSEulu6Z58NBOQb2DwKYV6NUjdbLmA/hAdszCEtfw0voP3KIr77In9XKlXda
dvuglYtFVDSj0sH/1AjwpjYpBWgvh5T2H1TS+IqtsEpWnfV05GdMcBmF4MOwSAHJ
Lp6XzIWvhI2ZR4lAImAXDQOEBfvIblRwcdx1Mh/shftfj6KMIa5o7vPC3sG4wH0T
tnqidHt8ql0zolVhbvyHfZKQyA01Johf/v/kzIn7zNdONiv7tvKR3T+gDbxDUEXB
Py9bpDPqIMXHy36Mu77ZbEr8FpmwHjGh/4IKAa+ObysB0vAFod9I3vogm4ry9C53
Bls07GTvuz1smN1F5rgoAlBvqbwmwDaZ7NFCV9iwb7iBMJ1U0+sXF04OmmJz0EIs
6eEH9/oilCsf7Rbb9Kpjil/+g4MnjxMMzb9bML2Ek4eP1STaNU8P9zbzWFxpJC8S
lrD0GmfcFzJumYuoh8ltvB4Tni702XyxYc46sXXNo+MM0lrUQ0WsNKquytYOCdz+
fjAt8eKvyaO2E+E/XC/MZoyZYCvnKHNvhCwRaZg4bC4QNc68KoyUZ5fXhkxq27gW
cq3LITudALWCgXVjiwOAlfJ5kj4FWnbcURnp8t14dLc76i1Hebdj7rAlFQYiUm6P
8jikt+sCaASrz2nL7IrEcycGbcTXNYqxtGYJI2fNli8RsAPirHQ9QN9PQ5AriC1O
YWjVyMLtgo8kJsBAH/BGA0DUTkh0xNWTZ8GTF1smNrgtKNcrU1B1hrWd5US/wYp1
TKQUVS0J4YAPu/umU0MFY/NzqmEhPOkLks7zonea81iS+6m3ucofqv/Hq4ByHoPC
SDNxoSM9xxVM7uMNgySbk2cPgvSJ0xAKV6oxQ/ctiGcLqIXdeoSBeKOkER/l4Zqb
zwjXdiqRBSU0JbHc2am91rPsEuDRsVLa78rZquMNNRCGx7loC8WijAbfojhrdDtK
K1xgAvwlpK10+6629nYTGl/ufxG2HjN260wk1rdrQ/ObgEOdWZjt5qxbkBzQwrr5
tbBRVNVKPqhfyxG18tYejb24Pk4/jVOzihrcteluEPUpVWbQ4KWOm3w08U140eTy
889p5pdpaebbIRTcyz4WbwwXJD9FPlVoBtUxVSGDLDXmQuBUfdn6rSK30+TWW7Pz
3v8rHKzAmHJUxfL0ma8Kz3R/j3zw8xZTfajddCWG5R89o/8EKdj9xTXEgfK1o67q
4OZDQrXWI0L0gMhokWWNrwWCjdAD5/DYRPc2+U2zFqAjbzfJ02RrMiYBcflo5weE
m8D8guYD5QwMeNW0UVBfFIetjecz7ZMTEPcVSTQt6tFrDkrIBUNDne4B1wcepnSE
T0UMikln0EUAaAeHBIsfKiEwyfYKA063IuEUTFTV0yDEktAMs6qWwjQvbDK+w9vt
b9+G2KjW4cCxuqF/Qf63nrbBcYOBJqlvbm+E4g2VPkJ8gl7djQkpzpDS3yC8wlQR
MBhBv2uBtc7rBxt9TRYoLVDmIhniwQGnA2B/zLMNDAM65ych3R3POT4FOfoHn5mk
dXUcwmhjFPMZxVfTlO1OdLA8QwXvj8FNit1bQzowGX75bTdEZzpQl5BwKGUZWQB7
bxiWeoWCmsNS2Lu86epYtyfapxq1SsJrwVuTQvBZ64GsfYYO4VgNNgkqat/eKRR/
L5z9BvydMZO/k1iHIVCEr/Nd7Hkmj22rpeKwpuUy9b+UrI+nfewBaDN4ezrxYBWv
nkEZ5LZzLrvCIdWRdv5a4X63SAl2g1aY2dEC0vF2LvEWx6JnBjagcbLS/wtlZJwK
YgZ3yBH48Mu+T+IDNTbQC4l/+/c4MxT8QLYYqSLowduROMdk5aLTY7UQXFpBzwKC
s9XMEm2xqszEWUWTYhAyLmJtSoepI1sjCTkf+14p8upLtAmqSaS0JciZ9dO9PEKx
S+0CgSaEG8VYYrg6YsWfCaWRou9/EypZcAVUoXF617ukqea+9olELgIQbY31/v6p
LhuCBxkE2ZbHYRlkrMJYhaRkjoKQlHswSK/jcSlPovR//F+zbJ7QJxa/4zhgyHAs
3rtB3JazgU76faeFmLfWDjcwdB+Vw8MT92dD+EJ6ZqnvusNVbaMp0R0czLPHnaYe
0yq6eVKEWpSodKbp94PDOXukfvjPw+Xgqf0uC++YDZhYLLsmvPd20Sy2B9BbDnVy
sbb1LkUjcCgGbSfeF9Xf8CSx+CprR3juAeLnvWjBmbKOAXDZW2vzXPkG17zl7GH7
S9zcuAOu2aquagfA7u7Zyy0NirOh8DvdqlT8nj6GnY/0yxQ4XENTbpkxCfjcnR2l
ZeaL8V6Z1842na6yEJ3TMaU8ACIBMn7Fbkyk1EzT5TPJEYZLoUn1qn9hg5RyZj8x
a6p96/a3a2t85QwoGg/nYcl1pkJyKTrR6rkp/ac8+FgLyJ/JO/utTe+23fW9nO2F
aDVXxJSTvjpvzCJ/m0vQ1CWTegk2jHG+v6gj1Nw5tIEegV5lyzqbBqeiwzit1tWc
l+NntgC862j4waKGH2Wp8F3rB0kXOLQscOtP+TpAYmMcwOa0xMEmbsqjtET2EMt/
NFo1ilQDVmirRjgP0gjUhExzAAgDFfAJ3ApLJ2WgXLl+r0arDId5Fo7oEdPi9HE0
AoB2g6CI037qJ64LXEOvymwjuFL7O9tFn+4o4hh1Xt+m+AQwGCuZNM7iDS4k7iF+
j27dDn7ZkY2x9WQvhtYqh+aS0f95MOoGSYf8tgl4plyOiq1nX8M7ZldVSruCJ+eA
5IMXr3W56A6YSXZ6u5mqEVlYdA7mVrp+a+EgoI4/Qw+aZUvA5uN5LZPzW5hfTh0C
asmxeSv5wi1W4PUnTWATQa6lqYjS6KgMkNMIsyL8GuhEMrDyubmrI5tjsk2NqTIB
nZtlVqTHUGBYIsWGlGeyuZRdy5YoIPqyjI4Q7f6vzmUquu8q8D3Yp3tDB5fz2j6l
6zs7ePH/3es1fDwgQKO3F7UvSlzf7zDFo2coypLQWXVRlTgCIsEBdwdgTbLbpDx3
RFp4T7p+iJJ3f6Vte5rimKiKuGeSmlRNP2l6WbD/4v+9znYOwXdf6k4f6zBRWGtE
oY2luspJdwv+5b3aBiMUVj8ExzurMr8/4VuaAt2Gc9z/52SZu+PaJpNfvmNKMlTP
PXg8FUL/JMdPCJD3xsLZiim48Kx2kJHvJ7WgLas1YbdqiQOwp0RWNv3CZwaTm0wg
UFGhNme7MvcH1XNFY9G+B4QwnAIHaN0Y4Bc5FZcwc5j5WRzjCKGmFLvE2lA9l3SQ
AsvFqpV/AODDQiPRV7dFIp1HdDBJJUnqHo/IKcP3nzIPyhZpIW4Cxt2edjqHMXaY
ldZFCJPrvTMbcdxTi+0yA3Ieg617Zp6ZmLGnjRc9RbKEQS/Qat0z/xbAm/QXw9p0
gO5C77l8b2PZ4ewwPcKxA2ihSNb/Ex6naZmyYF3X606nxHCnCqjbjHj2caTsmU3b
OvSX82HLWfyt3HCEflnKKyGkiFBDBwEJt1xaacBgn46hfcnUAtYCJugsUPTDX+3Y
rtdobPDUVdeCssvHTzTfZBEGEET48kt34BuYMsmANqI55dJbDxEIl5UN9bn8NtPU
+zScvu4eSScwR3Yd0lZj5AKnh8j6R8K1DWgDxZoIemYw/F/rOYocjHqkGZOXt/Hv
LhX4KTjh5v60CW6PdnTxWQL/jRJ+ekHh2wu2A/su78tqzsuiZpeZG4+SrcFMKD5X
jOueHtmtk4/zFlMnT23+ZX36fhZ77RctnV6l1ZindSAPO2CM1w2CWnNIdi0EtTRM
zjURipj2UvqcvLJ4RplvcJYeX248mAi5S1mtclo6awY3kJra5Y7wQvuHZsNBrNeY
mrmdxRjbbgNZOsBBtg+UrqXQgnQE1Hio5yU6rbmgjp+R+wH93pqXWCB23A3gkx+6
C1WYFLXLadPvPBEfLTem4lkieCEJvtwVp3xod6vRfbbRYs6mCdx8p1tNx7uWhtUn
PX4EloNYyAzy1IxdwVII5TfXZv08sN6Q2QO+9kItw0/xX1zHn1GP9JKadVW7Fo1X
ePRvMxLOlvwtnb8zIGO8ADNjte077kNLH3c9qxR+G27siBsblACIghp0bCZ1aoPm
hWAKmXi/I0llAfpFYWQd0zwx3BAsF4V4T5mLHa7BaoMp5bHN1CcP46wJ4OJQHfEN
i5Q6Tqo6Jolk2tokx0HkDn3aVIx5jDKEdmyIBT2yLataHV/hfSVQksowF7mqNHCT
xU+BntQh7zFC86B7w+Py8JhUIXEqPF8G9NIY1IzYSxGmkepfAA7HtjPnoRMj//Ib
E9G5Q4EDtwBIPCBo5oIs7xtnUwXQXaNzWSfyZhZu6JYfdnu0QhlRHxIcx8SAuDq6
IrkVW0P8EIbCuO8CDxa0hHSpjyS/Fa4ri9RR8FP7WHXI2WL+TAUrvAPQ32fl23pW
Q+RN+Wtd0GY/qRyi3ZEi8Voqw2umbRgldnHZi109094qmoqLgGS5l5QZxs+NL4Ai
FJZVZlVsBdyzn9CRM8rpIILUIT3VJyRdVwYLLi68YBTYOzgOFUPgHZ6kJNNI9LMB
VVS21ojMgHmkmggGtE+H34C+7j+UuLVdbWNDvTZ/yVIsMzEGZXVofsKXjdlVSZK8
IOdEb1dLjEp9g5m6CMN8u1RgPVQR2HhJReJvB20U7aFJYXXiZhFNMXXt2dFx5yo4
VyXpCEM/eKrGActJRfULERjl0KVjOiWQv0t3XczaeFHlqPCegB6az/SU6SiC8pRZ
W6WJ4lDoeTk/8NOKQxQGkpvxWKLiVxqHZwoRmkYMfvKJ8leXqORtDoxjlSu1K13N
3Pax1/WT/IfnjMJ4iJ1DENm5L9aPDBh48v0cWaeBvIBNeutAciDoEoIE6q91xUPR
fNTKGNVtE/U4UhE7FpUCPDKOTp44uUDI/V4koKqpOU3NN7OvMC3QxmzQ6HLdMWHA
2GlJRnWVJrd9V2rN3hASPqatabVOEugTnyjursBZlpNA1KvlUUK+PflY/4CzHcqZ
fu4Ps2XEVMfs9wHw9yhnBxu/cOzTz/7skZ1fadmco5Z0tSjnKd3W5LXme3yiXUoq
7Rz60ZaFkC0ah8LhHXeSh69p8gcTAT9lJoVw3/iKVQxJV5IkO6gmmRG5K7a+tUxK
9zQQO9TWmFNCs9htF3nJZ39fiGoKVQ7svXdg3Vc7NuzMQA6FcIM023qgvhsQ92x8
rM/6XPHIyHr0JodiDhYScyi4hY+cUVea5W5wiyJvujtIG+GktklAMS/CzwfwkPHN
aoebFTq9aUOZz+VO3Y/qKQBLEFMatnYIl4s6k/nha5j4y5JEJSoBOxGNrcLSYBTd
Vg5Z8Qn2SJ8ca/3Y2pgjZnqfcO1xC2Htw9FwN+sCsG/LCKh8BRpn5QGJkkSLHTgJ
hp/LoVsXsdhrxyVmIOat1zGJOdzLagWVyHGkVVY4+fFFLC6bn17GEzo46/BqILte
W0zqzpIkj0A8dXtS/ulxPZvsI9B3rotXeXcm2/y5K02BqJqGzAxokji+ZUMt39/W
W/g31SPJ50QFO1r+sF04mz39tyZFspf97bP0BhRE4uHzUcc8YYXwmXyyV1w3MAuy
uqQaPNFFTuEMBQPd7QmnQa8oCA0zoz6DMen0EPELOXH4RFL1W8GsxbfMz79z73l9
JZoElUCfdFbghH4KDvantnKq36qAmLzwPbNmnbvVG2hSwuMoK3CuVPIG/MCUv9/X
MHLzLSjE7FlLB7JTs+5TONYV7WQidBaDxVVzV//5vpwGBsyNeyhdhmL1h24IlYEs
kWwb6N/e419yBSgUac5uiVEj0I8PpKtIX8DS1TjLY00Q3VAUyduVginvQMtFn8Hc
QvoBXdPPjUY0808Tphj357iodGlidnHp772TjA93awZBjCHln3f3z/TUp5QwGSCK
gyTahD5BEW2OaurD7815diAMKdyTkzZIZM/o6NXgSNzBCO/NrdprfA4BzczV5jxH
IU/kxn/hVZctRI1pxr3a8jl3xOJdfbL1G0cqsoOg+DM+m65b3qtsBvCsGOncl/PV
gyQJxbNncTTpmqLp1sMUhOrAjGUpvNhToAoT1jxn/NxdOVF4+WtjgZkMDJJLBM+1
bQR5GtnKh/QXy2QRI2rBpmqJw5iVv+2QwvnRL7pJaiI2AnVUVDs9DNQztwknuZM9
lCTFrNmyAmhMEQHATndihhhxG7y6oUtRwyREIN26DfNeTKnye3fDTzlu4dQsGvj5
KHkFeWqT96UNT4l5kl0kJC7kgzZqkSfOSkUwWlqG97cF6fBXUGOKkhGQXvEYx4A5
VQNwWjvd6Cnn+yRuI3zUdqbpSJLp5dudUowP5TsozUp0j2l82fW+dxn7G2n7UsUa
QNNLrweKvcQPCLvPmd1820WbGiFTM1U/lN+84BNvrIotHxnEUUSh6gKFGDTUHWG6
1rWqEWd40aXf7AQB9YQXIokAlLGYCM2zFp/tIBDj+3nzdAYpStgLdE74PPsCQNkm
18No6ZB+jAh8UZGuZ3aPZ47X5NmYRiCkEp9mWZWMoAPltvWphGWwknHB5ei5sfwZ
opLOw8XUiFlVasMejC0uKs0t3lhbtPzQPEmbKB9z5VPCMQzvvmJAwKsjrT7YGBDC
3kqqcUJHRVwxTi3+kct7maPKq58hZolgzmA4U2uFhNevavZ7eO07CSZQb9k58kBh
x+4gfq5Dy0tq1pL4v5ov/BgkAX0b8v27PQm3Cdk+k7iviziI9vrX8fhSsRakLsAR
sBPcykjxulUSTvNldUnoZlRPQVuE2XG9ts9Pu5rJNy/qwxj+4hxPmwJbB7O92MlY
2EVw17PUlz4NXTuMZ5cWl8rwff9cs+WUlGut+4HePQKLQVyUdwlH1LkfevP7Qjj1
PIe/b4+/1aFE1txldooMC5sh0XRH707k5/OH5BKjqWfbnZttta1htpwofYRMQ0g2
D4f82q5avb/IHejMk/3XTvCtbifSdeuuN76LF1Z20GJ2Qp8M9zHe8HdvQATx9cbm
xZ9t/NvlH/T4gMwM1HR5VcuLOWCM5HqFOevPMUFJ1+yWHxnC/+H/fWjKsXOedR3o
jj385M+2kWDgUWnGmf+h9hCLsk+cTs3/hUnEMTT43qAdKNEXAmWCLFuKrwHr9LiX
tuDm0KUUrrSZPq+p0o0W0jGe+FPNUmhCaYAOWkPwM+do/ALqCQYnS6xfnUamcFKX
yCCNuhjRybR/+GxfVUkX2fwU7ZlIu/9N9y9acwFlhDpR8FoLSuf5AmfPAWKCXiht
X3GARz0Nu2v0OwKwSX+mez4EM2AySH4PTEZ/R5uzlZusHkP1DvLdg7g6/4slOtye
nrwF6ryfMUzW0hCLs41ZzkZP76tPXzSkNiRk7TkDoOUD/HfIBZ3u+WgQU+hUbZSQ
qfJsYrvv0y+T0iqIjLOx+cfRjF5bkG6ioxuWUvmsg2GsZR/FNSvMmVDjd/KqYAyM
yn/gCgUEptjVgfZwjC7+D97lDxvB2ij62KWD7jyBgUC4ENIHxjKkCuQ7CSGnbHYA
J/wyGVdcE14/QogbYdGipuqXtSdDOtIvk0ixFPzaL/83wUsS1chJkaoIbJLmxEGn
Jt1r00QYoNnKMnMfrtSC/TFEttwmVp2/1pREsk12RxwV3eDzrTMSC+U57lgfAPo5
0l3b8t8R9JLP45lu/uHajq4nAbtXQ2G9Ku5GBWor4q/BTDl5H60Z4rUezTwlCf/9
EK50Tx6bisWc398CXvRN2kgPOXATkchnnoITi6IxweyM/VXjwB7u8XYSP9YVDUAQ
0aUaRB9ao4KrKzq1vMsLBGGpREtk5aKjCXc0rnN31erAGZ7sqF8rVSJM90QVz2MU
QNjyj8XvBqW+V+H8ktVr+w+rgGSNTevAaFnpweutRU8ZjsPc6mn1dC+UXSNcFrcb
pznp26mN8aRDqrQMtTdRA2GyrXjBQ+2qAiVqDVFGEp+wOq1vTDBpZemuuRmXjly5
GxcMjm5e9QqOiQMPVSA373YOdOwoFw0awauMJdzLSZDYen0b+fhu2oJ2s12JHVUV
TJVWbP308MC550RYGuMONTtsLtScWq+oW5J0Fpydn/HTkBZO1Zam7yu25K+7O4SO
mz/PD/Hm01rsFqB9oBTbNymFgeAMl/elMxGRjACArRuWmeQZmU0cYMVsGUijuvLt
tUphGqFmPyi2z230nU4+g/Wu4SAHYJI5nzCwt6vOuYiZg8AAJR+mYczQi6Xoymr6
xQGb9Z8UoPCJc9p/iB1WcWDjIZ6tVStnUnUkyB4YJZW/5nj7XNMK+L2H5ff5+pYs
F+sGXPAmQra1LZugl9R+mxnQGfSPrAT0kCEkQoZq9y+I5S0/3iPDjpNVcsmpI/fT
up7Gs+z6Dj4IsqrDkbqrVpBzW2fB7NFUNgpu/paic8EXqdUm7aVwjF1PtlduE2e/
zfQRofZxyE3Z/KUvRVpXzsekWEwZf7edOy+K5blFVS/rilYTS0/HqFOM9dukvJ7k
MtaYTQt3NS6XOiZGV6aV/vUUPfhrGhZJO1SSiPEXSYQIrI7KuPmYF464Uje/gDf9
0lc4QBHR3alzE/ybOGE/1tCEiDy6/W+GO5nF7y1nQHKQJWrrMkc33vRl1AVQ20Cw
0ZgGHwESZHGSBuCCM0qF1duUctTleiRmoUOTpr1r2tob9Pqe/0dGO9qqO5GKU4hf
ujQLmFkGH0oDFwWKKphD8YdolpDMy3XfFGDUJ32Y3iCdKm+1qfIOjtCYeDrwNtrA
Onp0T7qgXhXj0JPeIQ8Ib/NCmoat/2Z38PVY/eVAjjYRf1c9WWREUnxlMYBFJMNU
bggXyYDN27JHgWlAxHcp7sV+PqBBnG0rtkkG7CAtQY6R+o96QP6qYBD2y0VJx/Yh
q2ZamIORRTGeBu1aNBekKevrE4B2UzdTA5QpyNIy3s+SDWycWKj6/euyKtg6qdvV
8+6TMp6T7U5gO20AH2It2efZYNJDK3eDxIyKXbfogt+KILmmlOV2okcq2+yXx6+a
cpmNLSImzDUr4hbTxH9YyMh3VlEdTvSFK+/H/f6KwIMxuKNei44V0LRdCWbpxOIJ
YzWsHIIbKFfzH0LJHZ5xY31DOeuORTS+v1Of0M3kHkX0ILoeXwQGrI2TFUKz1bOd
KPgryE0GYKo+aHsfQd5IGaxzilzKTtpwTNKHM31i6gx+PM9+GcIvxUhOZoOKz+rU
s3AJCGwJHOO6Z/LbSxF/Dlz1kHURTFdPXbVUU4150dTNbDWVeiqza9Zv1lDU5VP/
H+tdL5y4TQAMnUQ9q2pGtAzDgof7QQtARkAQPH3RzIHzGuQNlrAMCIgLCZvejV0k
DmwKp1uWj1MHafDYTX9HqU8QIUf2m7ssLngfQ18Os+mjghTkS0yC3G5C8jf5/wu/
QDJ4xzd/0k9mYpaNyfPBAbaDOKdODPhnl9J5603b5hq/SoXN/evz3w2YSagsM6ZW
CWKJ45zRoUrLAZ4OkSCwoKU0j0RqHJIZMQFN/gg836gSMvB65q5ILG0QtA2tSvxU
it1+FQ9hwFfmzYR6DLk4AwvVQZvRo6RnhpitRQb6QN9uNlo9fFDG8bbpDSDHGd6T
dnb3Hm334klrqo8iTA5piA5ih0aI0psDRq8mq9i960tGL78ikO955yg7B1S8rNeq
fwyNbMjdtaxa/3ExRnI/5f7+mLsa0rbNSIa8uHdRFBdoKV9jILlONd4ROeQPJ4Je
WsERp3HZ51T6AJTRFNt5mjkTOcYCKGqk6k/EIO/zQWm6RvFRFB4tbu9iPDDC7oQ5
+1bGAjhsOAXOsphmurapzolBWCJ/IL5+ZQKvAlay70g4HciSldLBpHf5pmUAuI07
MPeRF0V4fiwHOr9z99P+ZCiUcMO5ra8xQrI9W3dR4wpaP3zgFomPRmqyiCNIw1OW
AkzjOVgFcVi86o4zLTVhZ0WbaZ2wDKExSdmo0M6rTy5CzYEK8yFXa8I7yKr/81w+
A6lXKhG5D9UTIwjvirtjPdq3PwWyj5nh3u0GvmWGi375xTS9BFjtlDT00v4b6lUG
UnllCs80TGiwzRmUXi3w2yLowSwja++IBmK71mfKuKrlv4jBatxwXo8+p5f3BcW6
rQ06D3te7xQ+3GzCFlxZ7VGH7IrVOnBPBPE9vWUEJRolsxmtfuJp0mNn+eZ5vuiD
nce8nB5x9dos+RTfnNNGASzBQSXEDXfty+WIlUet8xS8IBz2RD14jO5YmoVuiN4o
TkydWbTTqQE76wP1aDNoSr67bwNKfiwcK/PM/ampOAMMZdfHnjPIHx89Mp+h76Wp
RE60aIXe+0fsIQFLATcrATjU+BX+V3fUjIcuZ+6vJRi6S35Q990JYqjNSslmo91m
wAxNrk0nOgo/occ7tpOaoXnNuHcTmdzATiIwu83daAwGW9aq5QHDLSpkqLL1+zkC
FHsyURlFF1NOauS8VSR1bVAGX+Qc56UyB93tHF/7xbv2bx3WeAE1s6vtkkxWAuSX
R7rn8mkvUzioJmDHO0Dyo0Exz6+UOcYPjHDozD464RAbem7B9O0iYzDBGuTQTaM4
zK6q2FPVaAHWJFeCZyys4am4CmkiwaMAtUqfT3AR/NjknvIDGOEhwl+VUb8FW7CF
J2uq+EO36X9VwpeUdpYtDpOnwVbbIs9bqbCo5xoHLCOEMiXS2WA9a7iMf5d86Xog
6t+7OoEh0FuvuJ5b3zD/dx6CyvCFl0jGcHsYBXLTahXNdn30qnNUr3U9LTU+nim1
pVF0R0mqwS0AZB2ZlU1zajSoF8iyyf9JCrcs8dEiqrNEZk1s9tqe92Df6M/3F10a
G5vmLOBxqIx2UheyI5J7CZB2EfjISceXTI89dcShty2GUJpefzHTSMObCW4QZw2O
w/qzlvpW+SLNpJeY44GIgFMCbKoOyy+p8IgHzDBguTsLdBjheQRltfsWbtl4lOaz
0NwdYQguPWA7SNaIpyqyOkWpCJA4+lTLMe2nUkL7zW2ZblN1cf7nn51lOo7jltN7
us9lHtTI2XRav1z6FmGPnOSHg0+PtzExJ56KnUml7s3JbL4fhBjyPD54H0aQBut8
0kjJuQvm87KfyVPZCbQvOc4eotPKsEI3aqkDHYolP51NXqsG2NpVrtMzvDMkADAn
4bxWz/94WrcDhYu7VQy8RMURebwXXP7P7LqnjGAZ7aAOqRZTmaQO5xaWXwKTACDj
iQ4bEqO1NZK+5G2hPSm59m2xPCkLlCeT19tGES5yJn0DujBhMPPideZL2DCvA7e+
aBIzkPZmnLWoyhtdJAeUzLFNIf5s3o5zd1RbkCRAY94iNfUiwl2hbwDBhywZhdO2
7o5BQZfTgEYXNkpyLvrbIjR/9L1AlD+vP2/liqFBx3xLQ9rTsiK++ABDjBqgw4gO
hZyUlpQPm5JAwHryVjemo9No+YVNZgEeQckG47awIOWZrhVwlxXi9pK1hfIfJPK1
HEyLcSfjXSg/ewmvzRqhymmGMmgGHQ0/0RcXnAI8nKOPMv8P6b5kshlHmSUyWS5X
1pAj5FuOEXGcYvjzRhKWM8Hxc7NQdnNMUMGYR9rEPbtMIbINJxJ9/SoXsB04edJd
wbKXZFt+I4+K4s9sm6gup6RHGyxYXLQI6Chi6ewSEX6+AvxRzNMjJutU18UNg70N
DjBvCNRrs8ePEYIX+XKVG1PQfaZOMo1LFYFqDK4VUuhfQ8ovYrSonR2h6YhcSaxT
ceZx9ed8gjp9D5mfJb4P8QgL1wOTD5lq0vKGG6h/JbgqjoTT1ROVu9O76gmemXGW
bDtPqI7gXLL3Oxy0hDxWEUY6bATD4LZ1g89BWIbFbRkmNQyOuPuhmhWivEvV3dw9
w0lJFL8oK0sksOUiiI2Ek8IDV4ly4bkUmJcN35Siehw2NEqhMA1GlWHcZe0QYGch
ye2jB8L9hQHf6bLvB+SufNl+/c2sLvNvLozNcQY9aNMRP5STmg/daPOHc6vHHPE5
TIAipHF4294mT/B7oi6nu6Q7RcigK+MmCj0LHn/pbw77lHRv7y1J1B/GviTQ+iig
jKfmFI4IbOsvkBsOxuFkh2CvevopQ+gOOVzZaYGjsBf21Opffz7xGgZfvh2XH6zW
P1ihCM5SgAmyxjSkWhMy7i1i53dWD9Me+QsJUEBDFcCxL7/PEJ/dXyS9/oU9AY/B
QydVATDv5y7tAmVhK2/3IJPYeW3qXqNEz4pFLjGamFsTXkTIIjsZAiLlqOOaibRv
w8lRzRBTk1IifydqnZ9Xp1zE43v0QZ6Ezie+NLDzJT0VNzHGEH8z7zTI6SAMa6uO
tsjEbk1XtsHOBSqbgbKbRwfqM71MHwMG6UFsXE/Nj3W6xPUeG9wxnN08d/XAkjws
eMLjNJ/VpBDv5JPcBLzgC2bVnKxZlOkxhoYGxAkHC5YR7/4pNptqrUO4evMlTzHD
OVEKwvV0UiOfwCyTNoHPKjSX8ZxtHOyaY6i7U+GiIJk9GyiaGnCW5TbJ1Q2PcMV9
J83b7bK4aji/1j+UtrtDvcW0hsJT6pezkcJyQRqvZh93OxjLLcv/xoKx7DdZoZzs
JrDCwlQ3Ik7idW72POtnrf15EUruw1LqS/clziMqXkpuNJ8qI793S47uIJtgSGjs
Pv06ovUwpH7g3PHwGImS6z3pJcx6rRjsB8DvXVoDErDmHuPxOqlRKqHYhiLUvdzp
zDn1DM8tiZH3+0NJiSF5yh0iGZ0tQqcTLMAUOcHURPqMPgp0tyhz2ktzWJvRZOBN
4gCa4DP6k4jmf+65Da39ZaFBiD5kJRsk8dAjlRi5uShDZFesRfHVq7aIPNZhWkUc
tdrOjwnrLR9Y4bXShoQVHfeCjvh1j+fHmbI11fjea1bFKfcPmgVjFxLpvB3z6HfW
tPCdQfSl7zvRf6d6RvybU6FqX51AMAopoQYWl93EeAbuQ/VQDYmkd1dIdZ6bq9ob
lqarcarKgEvafbcq79pvuTIL/Eo2/teGeL3xAC49u8g1wFnNiYDiIzLQqyKLKy5J
2XMgkpfjhcmIEmO+0F/3lFdK8QHjmO0uzW46Kd67RfIzIRZgw2084GAfBUIx4hU3
l0WG9ys5fCeuoQCWJPzPcdlDvI9R08k3nr9UqggkFiSBVdlbPl8C8nB9nZsPSMGm
ouoziSbLHprrf4GUjb++cHGlLBsNhFKVR1hfW1EJMyJGOYZg18DsME/cyh13FFur
mSFvUQXq+ovtXfpEeHrK/6lpZGNyhmCgBu+A4HWuMaxGpF1bLhlrbTZtNuNIYpKT
akMQpcKW4tDIArSamPcpLnYIlniu308LHugC79g04w4sPSRhBIh6xq8TNUXAuMHq
ELrLqdg6s6tIC+QBNwiub2gmy2x+Xr6Q6nWUVUGB69DqkIVH/H6HBGisp00GGov2
+89ocsMfe2QZT/rijbIboYt/81kbgIM02owNLzkUW6YpQmHyaROlHCRYq/BXE1M6
UW64RLCT7OZQr/em3EFHCPBc5OC4J2qp1Sk1av00dct2XGqtzjilPmNbGQUArm7U
sLZfn+Q9BXQVka30gC13s6abFGoqwdfYqiRaqbKL2ojAhZ2Xj3IlW/FbOtjzBxsl
Oc8tcNGu4JZhpwlAQVSFa8t6khmu3rpJh9MYUasygwVu8EzZNMIeAdnmEco3Nxq1
DuYsvO9Lv1ACNFwk1ovq6yxvpGzkWjiMgd1nMl9kIpo2bf32qqgujy4GmZA77Xc3
7ToiLxxkpKD81DKCIcyc7s2BoY/CtlgtRJvzlaw6LKTAev/muKuyGqO+9A0DC+Nz
5APKipuodAtaKp03zspLLprfeOboSllQRr71JR+TnuDwd6RpzeLgMo7bONKAKTVQ
21gY/+T5y6mH+jWqoVyOx8BmTwnyRADist7QN8Mo5/k=
`pragma protect end_protected
