// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aoFsEum3bG9B+jyN7Fa9V8y6087l4wFMx4i/IRuH2rnJQ8wagOPHBRGFfoEl
9gfDgsX8kkkwieGCK0Ew7Gp+2E5bxJDRqHui+/Y7h61KJaAGVE/rcDqOx+iq
96d2ZzaxoWNQrTV6QCzSIk+ew3NQNGZtCzgCylr0wgnOAwTB+JhaM88+jpFX
4Dtfhr0lgc8bUdBTJa7Xmr8+ED4Jzxq+HQBkcFYaP2DSmWdVKszuyiZw2K8t
XsvgyEmwrp+FhgndDhxp43Z62rg+YSa2H6gGXy3K0pxxs7u0dxrXNWopXzBE
6ZGt54kuEacAfECijRVLTqHbsht7y+1+6Ze7H9dgEA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hOhiIdeCS8jKuwqwOTzxW7UjBQK3SWMof5bnNLoRD65h211yVkRyxOFkwCH2
pIPGMsjCgzdQU3KZxSdjN4gY+h3TpPw7Mp1VqcyPmmENlX98Dsl4frsyavOZ
7Wh2R/UEs5nt7y4lnn85ZyhfazDPvdzRi6eEDKyINcJRayWnf11cV/Vjmqx7
RGuOuBJc1rWZlhjJHBCvaKuG9XhhZuDgqbi0AKj9ufKZgs6r31b9ksij8NGc
VhXOBbqFx/utH0hruKqZOFfTA/TjzvGmPwwjXWd12xbiwa2IA7RbY37hilzL
e3ohjzKdqFisiQDTiCNqabryMFbmzs78d/0gxXNxlQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J0m0yDm8HMNL4AenROg/KkPMfLuWmtybxf7cox1RkWNll1DaDGvA9Ukog8oB
4QflZQmZF4Uluq1ne08h9TCj+m0U8ZK/jOC5szhYPVfE8Lm/Mh9r1T0HKDaL
D0TLm8twa5o2oaeiBSDQuWetr0/Ij5w4WOEmNKiuZzMs0DjiM0oEbbylxyN0
O1H9MH+VduKNptVtS06DAmPRHxvAOuF65n1ovgf8R06ZyEllQ9zD+YOlJWfT
cAWCMuJjup6ZpuZXc7lF8wlMuj757ehGjISmv+o9hxkzFHTfEnYhfOTKf0gy
ZF9f8UmrYjQtxfeGopkcdfAdnEC2PLwEGUfGDXIalA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Uam7Wm5BnVErYVkzfgSjW06oIUgznmkUyGByEDeB5+v3Nn1G0aiPkxaEUJJV
WM/yl41TRPKq1NNg+B0j0i+vc/aP3HwGvxsd0VQAUw6UMghb3cSrGj3o1TWF
u3eB9Lqakc7woZDKKczRosiKbWfJqtSatonRl0J9FCqVH2lWJZo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PaavSwxhxxur8ec7Tnjc5tCgId1dCNlNI21cV+c/zfWHKjJvdSc3eLQcGPBC
vf2D8eIgbfptEF6JiCrebt14s4Hfpl02qnOKe4qJ0rDMgpFm5OfDDrn+fZc8
/WoAUMGI7u3YXzlwgc4OC9d3Mrp/d8SVpSFU6kehWMLUSnVveTsUKVjn1NfA
KoFLzRat8uaGyHelWCtv5m/EuwpihwK5zdZKZUgrQFi9qS5P0kQT5yTpA3aA
nUM7Cw9bZflG9qPPYPVMLkK9hJYbW3GUVuJEj5Szlho5jElbcB/o6Y0m9iUC
pUjjwDtXBmvlmTCpLPhZX9/9d4tLcU0BJ//XExuFhzSfRhkI7+95qZLYXY3N
PxL4wzdRtOtY3yvfypjjSUj8zVdx8OOFeklNe/HQMm1o8fef7Z83N2O9RLm2
poiz7f2k0RR/2HN9V8k1kKiJ0hJlCuR9YA13egJBG9R/HC2mI1O5oPaOKs9u
lLGFbQ+V6LtAuHBWoQGAZvYYtrYds9KE


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r6woMFiGti5UwTzST0VQEa6waN9X6rVnuDo68hm2v/aC8yJOaqxAHHUEz/am
lvFk/sJ2isZICoZSUOLEwfSEFsjGp/7RopVjAaa/IsCimJOO+M4U3CcV0O4e
9GRVsJs3e3LBAAoTGRAc2i7HAnu8jAiaYZSaKFdVxdzXPZVeG3Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PVzCQ+pePGt7KMsqbV9pr6s7pvxfcdQTxce8yxgyOGMJTCLv+mTlLcjW+4Yn
0uKgxv//CcdNPOCwkzNp0KdIz680WVl1YpXBOON4kXZ3tAFCPn+qC2hU7z6P
N8pwG0zvTum0V0Mig/3XzGSEpGnLKYZNaSHKX5pWvuJjfx1ZTmY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 66800)
`pragma protect data_block
V6q93lgzXYjJS314gl7pTFNjbPKiny6+px/AIXssbn/IlzkSuhAnxLVN2ymd
mz+a4r9ss//wpdhClOjiMZ60TVgrh40+V9AOFRtkZWyb6fpqwq6EM5MvwUlA
5PgRS4N7/OeHy44HvSxH8dZ0YEKgXKYS7YMWSAcrH1onx2J2rmsa7BmJg9sM
RDcdfzUjcd2L4rkDr8bh26+xaPHf5/5l31W++Mno8elz0+UeROSBQ4P1TmEM
yeh539E7qRq6VLSVJRbh0tMJ8d/GRVyitKhzvoaU4RSA9C5VyZwkGwRp/xp+
hmmTOCNSAQdw8nOMG444wJ0tZIWPOb7GQiUkeRyc7Ic7QkKQW0cgaehwhaTc
lpElEAvHvmTOJIwRO3NHpqigICEuDwwc5e4EwnxsFPOE33IEMzotzsaqFj5c
X/DbgqlnJf7DsbH1M6sre6MQRjx/+8wg5yjinEpnCgJCHVHTvmwSmGMv9vXZ
TwjJ72sSmgHAiklRcNwtS/Q0HlmEmvk0XfHmtYx5wHXEtZdDtSx2K8BHXwcU
IEJ8ynBj24mirKRtw8qcvE5lb4d6AJrXQkAntI0ABmnxplB8+jrIJ44xBouN
OCfYRMyF187BZmyz7pn/HUs8i9agCmPFB/RU3J9QeXSocxe0x1Rajht+nKFV
swM557E0esAWlBEr0n/eMLn7k70Gjsobg/yh45ZLbVSrsdXvvPRUKgjUzpuM
YnMB6iXB5o5FxAzRqCw1x8WqQx87ttV6VE27M0XZDtiSU927CKiPtDFE7Y4P
/r067RYwY9rnjSxKIKneKizzluh3kIHejWLSEZCf5ZpcBxvjq5vqVG0rtByf
2pSo+byz+ubHXzEvijEPtVfTVc9EE5hC1/1HCNqQ0EezGKZ1wCXhfYnTONwH
gjME/yKr+zgqjhkQ2JYe5MJuFda3oVOkBet0ZBVJvkmL6w3ATKHm364iY6w4
SyeyA2jftn2xobn6PX8WhHczQa+SVwmUC57uDid4nSiO9GpRW7G0rdyeTcW/
mZhsKCGkmnWTE/NplTvHCFSj3eXvnw33sQBdExbVMBxvQ9b66jWycUN6ZALW
lRqCjtgKQdEb+9ci32WQn0gPS9Tqr8wtNGBsZZRyfWY5Vfl+c+KQxBfPzQJI
8Bvb47CyCrbNr7Uvg25qJo3AESyQj1envMclJfFfhMFfkhf9w1ccSkXAj8Tf
vJGyRJkDUmQ6a7bRb4vRAEdasBmK2jjyXirnF+zjqHqiHAKd71tO/jC459Yv
Aiv6DMvu7Jxsn4huITOk5Jxnr6QpagP+m6/W/luoZfg9Ycx3MMDGWIE37MlE
uhEoExMcnbwQoA4L+KDZaR3pOUWtSWBI33VvsOhJ5WkhUbepKg0VLLY67Qo/
5Y+GZLgsbJsSk/ssGKm6UAIzrQLc2YqShfwdJq7eT+ptq/o4CRQ5zlDuIsy1
dEJzCU+QmMq6h6MjGvwybsEnq8Hn99Cic6KToGGwbmWFmDgWOvcOM/I21isJ
1GKMY+jKFT6MiuXJuUrwRmNtpk6xIHlnL9Nlyar26g+QZZ1F1F6nQU/oUE/H
6U+WC2C3OrPGHovgRUg4b4a2DC3iUzx6XPOyUyOgpcTc00EEuXq7D3h/XjIw
QExiM92YCAcssO2O3P6ifnyUq4Wt1Bb7NH4s1L0NoDlO12UpzdnAt81a5X6n
d3/kjjP14a+8wy3yk3CCwci9aOImD2gcs+sthI8oW/acxjz2BYPZVlzSsgqD
NDBVGw2gEGT5W0tLU5w3VNU2NxdmCHFTwRnvUkr2kVUCGysTJqHcIfht4x8t
Xwz3TOypQv5hccs40XLqzJsyACaZE4LiFc9sjAyr6sH0+6GKkBI9/5qH0t26
314dP94qV0H/NjM5b5v64l5YzgclzSW0ha/2BDhZ2ftDDTIk3YPEibUSL6XA
n8FyB4J0eaNwWbgrmAnIgh/zIxug9jJ3C89/Fc8bd9pSNKZvfPc+VJ0sMDZe
ej3LMmJsR/RClEq7L/gY8Rnw4DPYRzcSrxL8BDfx6CfOgmTJoj92R4NlwlK9
b1zIOtAPCPWFhFcAiVA6ne3SNRydy2jIhgIe/Pbg7zhTDfkIaINtL8aJya5/
fkmsJKSHs7ZSYS4enwQBhSz6OLZLvYVcUnWBSe/W1CI4C90YVcMXeH+N0qRG
VUjNh6bjB5kQWpHJLQ5PvMKhUoUPcE9hHbnJjywPx6UBGYH5LNt6XEZj5q+Y
drblIIitlSsINbC20+R6L+unJUBVClZI2SUCVcsjLLSs/5cN2unDBO91RUiI
FMcWH0wiWJKOmGIdR7k066jf0GeHIS3SHpbJqiH8gZw6P4X+SlmrX1ejMwyP
A+DoXLt5Zr2Ex9eGegIvKqm5Rk9yXqQo0/uvGLGptHmrRa1fREQI/1HbjVKj
JORMQA5LgR6+9VJA9jRv/psYVJh7HVTHrduT7U5HVwZVMMzCF/1U9ikAh1n6
+l6yqAKQByHCiMK/SjU/UyLeN7kmSfZAFe3RDCKQ/vtZ6ACP6tNu1L6fUqK5
+wpBy7gVAhqzs00cNfWfA8Z36dJWTiG9KJICiO26LvzTf623gre7P+TRaRdZ
u9XXTn1PkqCnwQrFa1vx+CPZYfG2U3ajaCz0lbBXHrmwAFh6hRtjbkYqr6Q4
DYzt5xKBYXKIbb1MT0857Y8DKmm3IPB0agBZCjiXVeH/KJGNrDIG1vMhOCWa
+gsVifjOocQWr/LMsulQVDoP0NcTuxotc/L01oIdr5JaPguakUWiYdAHR4NV
kNowce8XTgwB/YCDWKqlRicja9EMtbdeYpYg5WHzAcj6qBVaNbb5K6mGENyu
FOfS+FodiqG0XYrcHYtgQtYXD8XEAqLoYQgL9KPR/U1ogio7qAhGfMYOfykO
XV7EFvTL0J0Mk+DSdRnjq+mT2/89hMz1ow3/ytwhyYGNYc27TViElGpQL5YM
m0n7TGvVNIU5YOZRuCU034+FTmGgpwJZ2HJeo3/bh9nztopz69cprMS9cINI
CIbiTfp5agJx61KmR8y4qM+F+mad3t3yPLMq78JduvG9AqwOWrc7AtK4JvMj
nspw7dNNRbEBj/1jXokYaAQHE25SK3SdlUTeqMr1KTbxA773PM/CHZOoRBh2
7eiJddl9dkjlvLHaBzwoNm/6rC2t0FitXW+mGWDn2aW0l2xiP59bvExEew9p
vXnqL9GM0Ao5iXpDF5+pQYopKLbaoIb8erfOfTdZGajO3hrPOOkDdQ/eA3Ny
9XSDoEmFWWR69q2i7++VOP0KusSJ1oPtoos93bOEpJfOmA4Gx/mvNMzvUD9c
KU64U5p3tyqwsk410ILaKv7N35QK2vkGYqNxzKeoxDoRv7Jm+iguW+Jkb5oQ
L1IFVLUcsaF2ifOlhDivAUrT5gLBz4CFwAdjCyrITeyuZLyL9iYJi26eNYWW
2oRy+1zw2ID5iPfUVByvvYLpAzDEUXDiI5ncwNkJMThqMzZKwYctnfZVFyJm
hsTplFzvyUonqINodx6jcgBkKoS80XkrkmPnxyq9AlhhH7dhHglWfzNyWxAQ
d4s5puGyjJyvSNNfR5Ooi/e749o2EajwoeD0uAxgWDo7aB/VXWwp6hoOk8M4
cEbGVP70teicQyGNlHIp3IVEcFgZaqHvLXq6ZNObDLQLq2fOezgneNX5KhLB
JnZqTv0qoxV6qbmLtHHlKjYoB6T/W4MfP6Lg7T6PLaXBp2fMNP9NTj/zmzR0
iFSdAGqj9AkQvdu9lqtRFdmYoh2En/6JKYzQfmrpBvaFnSnpSlxVEG46L7td
YONlXSsWMgPL4eC+pPyuoRx13CbaN3D2vfiW3zE73m20eTtjnlYjANjcPibi
uQ6qvVMj20UnZ9tmONXwD4+F1Z+qm7rKWo9OmqMAfuJ0G3DQZ8KlzF1Ln9n4
NKyFCAsevZ52NYYTxlFYAx+dlbsvPi37e9vzm7M7L9tnGeFEE9jo4YYaaPYQ
HHw7lI68ukzIovUlEE8bkcnhGLJyqZX7DTMEm1XymT9ThAKpsce6o1K1yI9w
tSDGD1JfCPfzm7j6kGbEeZy9eXNNn+iGWSDwBotBT+WDRJkUEH6JgIGE9ebS
w5SBZ+r3yQ3fG0kAive1VaiCdF/deTKoqVNlgI9SdWMSbPcN1iOvDFLi+v8c
ZzMJh7xO3xRojQ1zLvThgPdYj/85Qzy7Hx5YdVKXG672aA2N7r7KEzCvkMMp
1UTx1FkWTU0e76qt8s/LBeau2ap6aTK3Lriqd4hyJ7hpaEdA+lAW918iKzve
jIE3ravTbUhKhoIzkoG+OLv5Cd3QnmdrfGodh/W3IDrMM3679siP2e87BwIA
GG0jl/cKwByAkjdrQerRuS7LYB7ekadVs0SHxoSc2hTj0YSULGkwHatdj1XU
mQRWrtSWGfArpNCwGLOgtwMxuZmE9/FHLu90ydX3vnX6mARLRv513ZNQ2it6
AqVy2enH2aOQyhTdp1qCeHDV4wS2d4Fqeew7fNSHpk5/GgbeYul1vT0a8dC/
ECh9SnWwY40tqT1KcXW6sfCgdjZ6QUqx7A4K4j5DSc0wDja5IdBImAL1zZZW
QQYmGEucLbCTF9PwIvQxaHv0Q0uwHqf2Dnd4w0ZXZeobKoEh0kcPTEGVNzH6
vryC1Qnc68fi52AmN8RDzbUC1U0cKtIorajZRy93tC/gIZ3E1/k6adY2XpkH
eKAgd1vtuS17G1jvNvdbHJvJR8ODOfpwQ+WRsQrWrfRQT/zfk/l6n21A53eK
2PTPMFyFN/xE62HqoVoMqYFeXsFQ1hxOWHTqPCW0KT6t1X/NyLr/N2aQSaym
+cCGu9dqSIW48vGgoleCJH1lAyqLX8YjEFx++UhDpQ/7xGJa9Op3/8MmJlMW
8EOpZAOgHSF9YDxciGmF/AfTRQWGgZmyTH/AJEPRUESS0KkhYdGR78fg0rZC
WiVx2q94ue2UTRFb7HypJbgvAF99uqEnMzP7Nz8ykXvfjrIZzwY4LE4VGgGM
JeFr/3t1COvSXRgJ0kMf+X/0UXzqxP3N3cT3m1Yp2TKQGPSiHr01/uemmKHu
tbi61IfDWvVPlW5TSWR6+1GZx7Q+8d3RFOc4qcV3pkq7RfHEDMBhqvjSdNKb
xZjI7aopR0udc8FIGDESDgmuFfflnSlWYZQm/xd85DK33SI8Hog9jjgr38+a
Zx2sg8UJUsu60Ma3z6ZYxJGpdwzHSQDZiGs4jgqmN1Ync+CbFCGxk21B71br
1hZHEL8+WqIoya8rhfVH3X89EV+gQdc8XRE0A4xz/CyfEug86tV5y4xDFN/3
nXNbTEvEQ7fWfQY4qsM1RRJuxD2NO2PmOL7u4P7jIyUwv3PALso5i3kaN4TA
C2t38YBwqw5rxHAwzGOVV0j3F58o5GkdWvmlk9awqJaKz1i6ywN5xYQj5qY/
mz6+Jnc7LEh2dAtVXZOHxQGG0MNEYud7WTq1vOcAO5YI2Sxba7YsGNrfInNZ
RyTUJzwbxmzejjfZa3qbWojAbETjhmqnZyCL1zBSv/b6XCgJGLds3Q2Ac8ls
J4rQ7q+2FBXysxDeQ9effpJq7TI8sVubwydjtWAemNpF5HLm9NiikkGJVEQM
mrE5zQkWLcA4jsR5jEEiRvmUG81tLhpf/5l2RxNES9n+sG9VB8FG5ynBzlZY
eUZHbRJwgkRW4U1+SKEkzeSHeTkinGaZpciUyZny+8ErnwjVPvAqlkOwajOR
P3JdWP4nAXXtnpdW+CaBBgWWV+7J6mKym3LFCO17lkwW1NX+tqKJYw4sr2OB
w6yW6747VYfL6GjimOyXBo7BVqMUrrSlj8Noq4wuQZHfQhpFAri0QT2mUWPE
msc+ow+6TtqiefeKHk/25K4DP9pE+gTyxlLTTAWVQb82wO3n0zwNh6HgcDuc
lBYpLO2lXSODFN8DzH921HSCJhIhxLTsawNi93MhIS+4mmfiEHhe76CSnHWk
Y927RwpRjv8mSwdkCDL2WhGhVD6zsWx23AdOd4R7aHZQ4byPwUjbuvyABIdi
8egpKFk9JM5jeuSBE+atg975Bb0RMuoFwmvYRfledKN3HynBs7dfjHGNMQpJ
DLCvpQWMG4fjj69W8mEJ8uY+hiIuDKSF2AfyX1MA1aql3aaH/oRhkBKl7Vm3
x/lDNP0VTjrjNl6msklKm1dt2tzxz6oz7r6eiDdnPlohrb7EpHsQcbw9hkk3
FoI4sKki+fFZ2zQVA1YWmOmPTs8BWyNdaNKqjNfNzQdWknHuu55H0tqgi3L+
uLNMZtt4UugGnu1xk+3ogcTMagXNvpoU2kE6qvh8gSBtJrzp5k1ftoLuPC0j
fxNGuwzg39TtEWHOWvZ83iCCoYjk4YrN35js0vNdNN/m59H9PAO5HHbcdq7J
B48tP41SPSKl9lJHBNA81xRB1EdDa/FZ9kV63wELfmV9yC6QDCFME5Fn3chz
fzVNzJrhxbgWv9XB7CokUzJf5Ik/sJtswPE4OdeRaiwEQ4pHmuEc727RP+MR
zIndk6L5KfDijVuMe3ns/gWmRftxqIir9tvxkfYD4naytkwghAr6hEVQ0crv
zF2pfXe2S65sCIQzC7vLXasBIf6Qenvk2pggnigQtCPdLfSd87QCRECiG/OM
k5F65MvIn9vD8O01tnR0V1POwjLCskLfr/Gs9SOdL9DzJdYuVlYewnMw+9Rb
oxk3J/zmJB5Z7mHjIkVHGvdTCdyb6jpZ23qQQMFIHFzLULKWi/KfZhYbNfpb
II33VEOijvpsyj13ObW9YL6RDkv01Q1uAN9oUUNM93HCPn8I+oHZXRqsreGP
lO/hua7T/4G9PlgfCFmQfHHmVX3vTQWKzCYLWkUM1/Mr1hqo4njJ3DX5sZVM
cXNfucUQkJiTFaKiknXufEDaqe3L/c7WNNNL/HpeDltBE4Rnk7//iRVP+iyC
lGOk8vXI4k2qVFJ1iiLIgIyih4/5N+MX7h2grzrLYsuGuJ1jvSU3W6TrA/mj
12klfseAA6Q1c79KPvCnVNQ/N0KYAXLs30ZktZNMHo+hdOprmJUDNZvvWGA8
yBRR30Ah6LpCWHNdXuNzmRr7TEnLULLlQhiz1Qy5A8jwwxpo5Cc7Kzt0fkb/
QQjxTnmaRRo318P+ZZe8AHnlxf4Rl3piXvW7JNl4bauhly3UoPqpSBpvNSjM
91/JOs51LfkkdR8QRVnW7ozpaADMjbrKhU8DO/PCNHTqVDu5IR4yDDdro60n
ERpekUCs2hD6iyz8XpnO29dENRhBovmdhd1YibZ+WO3mQujBfnGnVfI5ohGT
VG/CckEnXrUNTaODHt07Ok6g4srt4VUuhu3pnMBAXhtv0XkFOGoa0uh0uqVB
7VK2WgoVNGNSor5g91AaKF5Tfh5ETz2PpLINYpUqmF89hvPs5auENjiOnU2S
98CL8o/ZqMH/oA9PZOVppc2Tfo1xqvp+bC/VePkfRMTBWUrpMUha9GOYOWc5
UhPhSWmUv49bXx0BposMHsPK8zCdDSk8LjV7urHuP53UkLFfhanqqhhVfJUG
5FO1QPqfayYJsRs7FDmHiH3carnTpVeaYCTyjCp0j/wIClPZ8GSi1Ex+tD9H
+7FrWcsvlJPQ4eYCz/ZEbCH3UOgabmEtEjYOGA/Ir/ioJXSvV++P0PT/BbRu
XZJERuXdnTeWSlzHV5R22rCfItaiM9ecPm0iJgZhSotgX2DrQ9s2PdlvQ3D5
YRvLRqYQ+20tFw9dyCPkXwZFlbi0pq+Jq2bV8Nl7R1riSZUYYq4oZZsYVNwR
PlVpRkHKrhkvnaKarwPRXie3TFUwzEQbr9hMRkbkrRhXup0xet2+yICtyoDB
fAT1VvD3AJAsADIk6o4oAb09W02Y/q6YZgLLQu4via+O+gejmZ7SkBfuyf5G
DZQnPmjb3eZRDbV/4lRcvPcEaN12dckKmLp7OhnpyHXWdMVulTsP7T2onEhO
TGSeD56WCkIoS9gRzH9PYv6OQYm6qHVLJTGEPVn+HyKVc9CKuNNYGl11lZCR
xOAnQPV0yAUL/ex4fJCw+4LUeyLRaqmhhG7z9x6VaH6Xc/we+aRZlKd1g7i4
Sw17EUmP5V7ks/By+fnKNV+/37Q4o7ybJo84bVwca6cRDGMuHKPAiITxk+EN
bC8iNasOJ8pDuQrs8udYJSGx+Cngvs7vK1oDXOjrD4pi8hWVUjsCGgFFk1Nf
8DIorjtrziVT1CAQGgaH2PvEz9xLywjc8BRKMSPxtbBDf3Vbu/oSjiOPcJlC
ivYdr937KeS1cbgC46JwXgTb0XEqDusPRE5FB1Knx7BXK/ZCnPibVxMR6cj5
l3NTBT2rWFm/4MEjl9jDv3l3u/oiUdbWGWsCoMhpr5te8SPwt3brGfuZVxil
cumJQ9hWyLwTcS60g5cLD+s/yfD53nDmbxNLBaAxwqCdaaFtUV6moANQZRhU
/ViYAD7dtKO+UirSgKlQ7RYPIXhEimOxFDZW97TIsKvN12Ph6eagxdJRG2jy
1VdiU74wi/pc0sBm5W4J8NH9qLlDnmWDAia5rhkT54WQXX1Inf8pUhfvca2u
HJ7LbCfly/BlwaeEkpZutIZI8J35i6Ad0xcuaDhm3CEsvjnI4z2ZNVQf49zN
dHxCn+CWwK7Cxsmf2MLpKKmv7dswM+BMF6kXXebfoojenZP9j42z2tzujfc+
gmtXA/Q49NumddyfrN9fLQrie7lglZ0HEUwuv2741prF8U+2lvNi60Be0ZJr
djIhoMvnkUjU8aGiePOyXKTNT/7QpSZ13Ofdd+fVVlWjtgGKQ/jm19SZU8RM
+7y7gwa05pBKpTAfB92v7mfw2C/YxSqpW7IWpVpQCyyRbX3lYHph3w/c8BC6
VG1ByOPc0CePV9rTeVbF7R6INUNmZ9DhJLG5XH9qvQJnwUn784YPNAV8w5Ky
Gb/jZ0IyK1RV/LwkB4GU+u3Pn78T9TUoTrweeWjWNoNE/WilCo6cdpue0JLa
MtBOnHt94/t8VawdYVYc2E5gaoU0mVFmdKqiNQoPRLpSANp+7EAu8w1iZaJL
VoEQXxEiRn/ldh+1IUuNkkqW9QgdDRI7k4yL/TP2CyPmmLP42qw8hhGP3ehu
fSdlEEiUHZXsQHhH9K4wAfrb385/BguulayM4+ap8JkJogXyGjkYSglmDALK
6dSWfaC4PevPtK0Rbhq/lVGCNdbJcE/3lHShcqlvyW6mROFcXJOow3jk1V5j
4qlTJ46LjrRX6Mk0/336c3aVxoVY3VJu/+knGKV4Goqw5fE3PGn/PDOeXBrv
/5lH2mmNTAd+NAaPL1dG335mj3lp4Je3vY/JeOMOl0YrhewNSTJEoQCGVcmw
534XZAbr51gEEs3jJrwaN+nH12B+WPP3XcneOf6Dk+ev7ncolZuAAQTplkEd
MtqCkQPoCQVLDF7i+F8DwsSi+tt3ymyTa6mw6A/MPoDMM+lCZ6t1eN2zATw8
0dty2r7/3bsGl/pzIDjsyx8VtsrLHieocmsuNkCbdrrTX9/yI2Z3qo9ezSyZ
XQzvD17ewfF87hsMy+D2PFb3u9svntLtgUCKYAZLXueSzoS20rSsJy5gIL0F
696uW+Tj+ydVAXuJZLucVoxjZTvvxQv23hiZnxF9YyLvx8EZrwS2uDF6RXfL
q1XBkoUvRIw4JiBWnnhi3GJv38+V3gzNI1cV6/3lmBVlDW/9urL2CLoytnjv
mldIR2ccDKLrM3S6uPXajC5UDexUUWQj4wOgzLl/7MmbhqEiHgMqonJOcrHT
4CnoudZcT14RhvR2UEOWl3JXpupmbBZEIKvcWlorY0BBWgInyUY9Sug0pSOs
q7TDhU/lR/rjW23hzHLSYnLvokjtv2WMg6sjgoLVdy/6MAGfinjxytNhg+Ze
Rl3wk0Yar1UGx/yjozEQBCOffFsU13yVBNbehunhgM7hOrBcOmBxXVBz8VUl
rUniy0pLtNERESqjQC25+8SyATUdAD0L0AOj+52yaRnLRiolCPQrLx6Ab3T6
ANjw2hwdH3TwGv9FnwYhdzdsNYmXgW4VnlNlyYUbDQqqrLpBzMzpA0zUpcCm
Dq2mRqBsXvbBuVnx26/QdLIu9P8EF6E46SlGw3mhozefD6XdP2W/P0FQneH3
sx6DF6ejXlf5Wh8dIiFIG3RmYmLLxaF2NisOP5c2fJe9CWcgduUHq/dXbzjB
VsGX1DHFfRu9JLAEW45ftZiTCkncuaGWtVFQvoIFVHJHgfTVxRFI1jekVP7Y
yzgdol257kTeK1id5efX7sTzrXnX0JcVZZkJORyxPxD7IuSi6MrOJ9HseDDL
JhmEDJq0xwhpARWNz0o2KQVO1kDufp53PWC+/uvymns6WC7NETxPex2zo/dl
+Ds7fd9NxTiuKqVRLTAOPR8/TtOdiBizKwg90Q25cnPZMQ/50RYxKRfJBScW
J8kUwZNGBIj6bSjXnbp4QxefVaPDLSs7ql7r+7ByKkq0POBOfrdp6h/pv6MR
Bzd7SVYcs5FU13rYNC+ObVWl2s6ixg8f7CZZ+tF9DMcXDVaGEbeZ+TWY61fh
J76Ow9OUYttNQ9HkkflLZidP7rJjj9hPhqqA4TPnAqA6iJJhKbwc4CQULm8S
+rPPmajDlBpawvmo401BaPQT5Out6kxIKKeGDpjy/daryo04ebBAiQN9JINq
wCrcOqawvqA1WHscmvnPClSbcticEKvMriFiD6Mw88xKykQZPWsYjayIQXB8
cHOywi+hFEw08LSb+xozJ9hhZYfFesV1EQVO8epku1bsUNCDE/tvXzhKS51w
gN7pTmWUGAbjRDF6FF3DMdOcOqLeMDloEEERDIb6tsVVAcOxa1aGzwXOWQCy
F4ahBPtRwikuCvjliE5gffCJUu4qH8l8fOLobB7/aPaKMrrEzFvvtTD7OhsJ
Prp2633KukkBpwBwIKzQEoXf3sO9tVLOn98WxJOwPAI5iyAhLoWAzJTOk2jg
RoEj9dQe1RCSTXSBE9aJdj+kHUfcoJRWXw+CrJKZSBA1jysvHRKvdrfWE1I1
8wR8es40Nr0qtLfIUmvYfISqhgM1YYwe8OrGqNMlV5n/Egkwtlr9E6MzyS8Z
sW9KlKj/wfaYNeIRm4LRJggz/dbeFFzY4VpTQPoFLiiSPJs6u8e1s5yTFv/I
eZdkAwri/B2kjwkK81/Z6rQr1SCHG6DTi8hyLsOOfkZZtTZ/ckHe4wy/hMwG
7KbQ2VrrVwRbv08WyZRFbg1hr/5pzFv4qX3cYUw+R8NRAk8/HAmEm4/y+/Sk
bU2ZNLp9Q5/UQFXIAETpHwojvhyyRfgNrMgv6EYNVvJb+Zt5+wDmsH9S2lXr
okoSlrozKnf9n/6o+wLfS5g3GuZWi2iN7EC6wd6UhYyWLCK+iTZrIn2PxFHB
EQhmhlP+pjAF2A7//N4UjFoSh0d5MDBoOgyXOG7TdRvP/uOZTWBwugQBTE9J
CSa4PsZfeXsceogcWuKf2Dta+GNyGal/Lm7D6KLWNpZRMeKpXRzDlJ7+lLk0
/iPrBmmb5hYRX//zvD+RLZrNbGfHNxe/b0kZ4tCJoTnw+BHKg5kPL0gmRC49
8Zh4pCF2dQkJbmGKW8OL349z+VujIymCVDTW2ZrJugJOViYg9Au5Cfmy++eE
lx+JIZF0xQMG+RosuU/jmGKxw5NkvlnY0xnUEVKgPikrAAEz5qI1wU2JUxMx
dAg1KFYxu7ocv8XEfqlBMzqkplFWmz051kg31EW3+uyAbVY5F5PMadEobd3d
F/zng0SrCrFj6tqXPClmDfk77Rc44PZF74Z1s/Dj1LOsSlxw/zJi9jUJZ0Ko
WmL58GInIF9pYOJgICuMCcSpPag3LVrugW1VAluqEbMOXr7WuFsbvgxHQzzA
slt2F4m7Z2eY+MXcse7SKRzAtI0P/d3ECs1hbaXfs1hYN8w/MmNH2plEm2Ji
AE16igM2zb+7bGbvUetrBBTzOpk/8Tu0cZYyOyuMqXJjblaZw/zw0hbFhWDz
XIMJ8rdtM04YBsYU961FY/QgLzpq0+TMr/uF0KJl1EPqyDbpq0yhzvr1Y3az
kYXcwz4LIZcW46Firv8c6eqV5cfY6I7Rp2VeBWLmmUydKOn3JU5RDp4opeCT
rL/NP5vnI3JImjy2AJgER15pBI9iDlM4ue40+VenzsAZFvLk5Yi5tzwuKmfn
PGD1xizvXlgov1wFM0lV1MiFQ3W1vOvRQQSU5K6zS0YTqgfMiJeOh9klFnaz
dGjeghitZtUpOBS7dfXfMga5hDOuOEmj00EVR5H0HQxqoF4lAd52nkK2t2vJ
I8W/pkooUeOI2BFWYLYOF+kWvr66hgRFEqDwVBBYEUBL2kqXrLVja/TO1j1/
V69UlaMzmGdz3wM+gHhJKk6LdwRAgbY/rPuKyWv2eXBDhyzTq5VWtPIyiRkO
3Tu5HsqpNEQgc+WCCm0bNLAYXdS9YXAfEN9Ns5KnvgoHXDheHUr+t3wjibRv
yxPo/RCc1mkYjS1v97v6vcFjJCmi72970DDG+L+Tto+v9BFEXjjaci2QnURJ
Fs9oZfqSsFdXde94MpRz/gpa/xz/QhpFkFY3R0lILlf0cRRYWMxZM8x+ycbD
rNSTbX+yitnORawaOp6rcxS9PfnbjDHwICYHdgPr1CAOzEljHoZqNywTNEsB
Q85du/CTaMR/PbtwhuoWgeL1ZZCwLsG9kVd9/W5PiU3TKwqI5NlePpxyHK9o
brqqbYACcSHM988X2nQsPvvuYsrZkfFg0L3+jN19RNM+eVOnRp5KaTGS3wqb
ZLuhUnW11RhqEIZuDgwz4m8PnQdiSEsCdvzSqGhv4VplkJA9mzi9VsIQcE/G
hpo7YQ+eEYzsN7S3/G1YHZTTFUMyiCRGKkxvEDzcH1KNZg7V6u6lreNkcWZt
1RFvGk4kdYWoUMvJFWsbKQ13TIr1n5gZgtaHNVajmGgAoMlMdSC4mvjKdU+E
HJw7d8Di/ZHdNq9v18x3Q0xC8qWEt+dCgrXZvl/8LsNzyRU3SenYO/jYNUo+
CKyTNr7E4dAz6tQZ6tEmBS1lJV3gCoC/uur/iQp2pOcFYixeSP+qr59qowBW
P/OCTaIDjRsBbE/6QYR/7s3AKG7QJ/RxK53p8OAsYKMPhNjv/mrdA2f3w1nK
EVEX0RLWnG/MVTjFSBAyvS9VPv3FJiDcneo0YH4YTzv/hiMbSNKdPh/LloXu
RDIMxqrpOZomRRg7ZGcPVqKoDLsLCCJu/m+yG+83LD4vXmGZ5mMiPyUgYrUi
R/n6XqViJ23/T0vnVgEW6wWB8EAzCCM4qBIPV98RnJ69RuQ05xkkfRF1+R+R
ElUuf9OzeHdRJC/Vlmz5beFF4u9kaGk3XREzRfHiK4JyDF+B1nyGhpdV/nUb
mOsZ8kjCfUrCj4a7aaPkTcRJUAF8D4LO5u2HbW6toLHeZJcOou8ozQsxuybp
tDr1Uu8VQ1npoGiNuukVpJUCWZNeUf8XwgbPZuvyod7oRD2P57GybB3gA8D4
IyVnKVrz4eXInnMvzZM5tXy9JOc0TB+MZa29mHclGHm3h0xC36sOOENi7D4u
s0wJpbb9D2RYcTGwpeyAVyvdxvgkGrt4COHJvX60Cu8z9WAo8dSpSb7umMcc
c6sKP9fzTvQ5Da2GgSc0VFU3cz7JHgu4p1cOSGBWNhymqCRXuHKWcake7fIw
duhKTic3uHMYv/ta5cCm6B92xCGqVa40AYyh6FusFFkhCUCTYPIrFHf8LaSj
CbPDy6ZVpC6CEAbYJiiK1x4NNukYJhCx9ZJVnv3ZJq1EW4f75ZFC/9TXL3JK
fb6mhNoFO4E1BpCdiGATb6VJU/ZSPvgST4Z1OAqsSOh1fKedgqNvLt3ay5cK
vfbx1y7kWjlWg4IH6iGZi13zB6jNfH+PONX+xIwnryCckm08FruYL772HJ0/
36IFI5c2b2WpgMx0TrWJpvhUMRETvEEmXaqRPYD/wHGFnt3cN+eFyVG36soD
D+3IN91YVFrornOFucwwrJ0F9C1lyR6n90nesS1x/ldPaR2ikViOVAhjCIpm
3bmvLPNpJMEkfe2EBST/wWEvypMgQRW4EJshvwjb8P527xzitrdDTvMGpBef
6HOr2B7dhRefsGxrOzXfaqNg35ikuTscHqxXtXRZ8b36W5kJW3pn74NeumLP
kaWqQAj5Cl3cOzFZZ9NVImp7pbRQXoPBRKqVIN0MH81F2RWHQyai3k+8/zTy
aue37XvR2GXB2uX71r6zjts8t2A2Za/oruh292nrG4U78yp8GEFvWr6Pt+1D
k0OESxK1i67THenw+lxwYjwShmnhx7xKcfhSGFOcRi8lNT2LnK83BHhqlL58
+6boMB5vtcxsqks7B2ZmKO4mhv0y0laa6t6nRLY7IjYi2uRDGMVO46Ati182
JWCMFOc5vTlqNBSAt/t6G4KMiwOhnNrmS5Qx1oUT27Y+S4rxkMvbtdngzOwf
SxujG8oT7joI9k+RlyvjYYQh4OzyBM+kHXHGJLSyrwjcHbAZ5Jfq0Uyo5vbw
65FlO6e547t2FghBTMsZAeNm1Oc6hbDXf20MPlzwUyx9eSIU+uqy1/ioM7Px
6D243EEH0rpPH9uWX0ZFbRuXanG5Rkeq0HPKmAnVNHiKhZj0AZpa6+w14fwd
jdyFPA4k3ipV4ggbzjQZJiOhhP9nIqQF9brCC+TJWPrA9ifAF8+FFew8D0LF
IaFKQuRDbSSRHd7ZouCgALQG6P4QuUoGCl+/JS5D+hWUr6tQsppRGS7IDsDh
IP9axHAJ0KAx0rXRsazz0+HOLdP6D59KLgS+lAIenxadfZG2e3EgHnlkxm28
RbIuX8/Nguv9Z93UR20nCPJuQoaHPge2LWDM5Heu28RkmAeATQnIKzThSHYY
9TgnzzukAk/IdmlhYwcG+YYWlBZnojkp7zFOs6hXFTH4loOkPW1O5FWq95iw
N+n3Vh+EDpW/0phTSw2Pf7a7Oe3e1/1XVFjrrcaPfVh4BYjI1ibxEb4eflqW
7abFOd5pXGUkZERxb3hlOUIXTJgM7IxBPFnoDwdOINT/m3xsZxMISsAOMCRF
/R8Xjuzk6Hdkukj+CHeYAdfBMyoJv8fjx88LgrOvGFVWXPQHe3/33//KuQJP
hsmbOeqoss3d4cc7J03iTbUnYi7JijxM5zK1QfuVLWxAFvVj8Q4jpC8zCrFq
V6jAW2okp2rh6gW+j+TAI9QjNp+lHdfVY5e2Vu5rhfy9OCqkrHh+0Q4cE7Zn
HG88svOGx7sYK2TJ7W7xEdIYPnHVwNnS4QrWpDjFuEHnmkHC1GgP4NvE/xcZ
E85BJfvAxskPZBj2B41IYAujMXzXaZcJUISjJ//QNg38p0UMJP00IuMpQvrg
Hc/1UT2v1mwUPcKa9bDmYnyBu2U4I3P+mC8KouvltgSR2mzo7t7389D4Ur3r
72CJz5q/79lrIEYTJxJYChwsmb+zTbkqVq4CzBAaZZZRBqAOw2dHHNky+EpG
vAOdiW3KXQ+jdsERFSaJqq55/u2bcOCZR89lTzuETUnDuYgOJdw0UrAbieUB
C5V8PkkKlwL04z+BZ+8LT3YVlyNAQydal21gtf6bTT/KaAnTIN1YqF3ofqlU
DNfbuDi90iDvYbM8PZZuLfysQjAFiXF/1Yi2DtUZPNzJm2wv5mKQoeBoOWzo
1y94C2gSUfNagSo4pDGCIKXOyBWHla0W4tvzcT310H8kqxXTPrfXAoE+HEjw
d8s198MtqIkKVPk+FXYi7vZqQcfuz9aVWNrKwSJl/OinBh6XlDENB6+GYazZ
4+JmpLhBgGvueB+OSr/qWaXcUJXB5vX2rcPpVGyl+a5kt0Ho0jZuW07G+CEr
bfnikqaJSur0F9C29qtM1gBZg2sY4vWlnuNu+e3jZwh++RwbxPReiFcoyBHD
H7ooW2SefSNCDZTscYGjv44d2lmv2vtPriaiVIYHsRpRYCcoDuGg3exfFWrn
UdLAjVqr8LprJzisqTt3l8Etaq1lUQix3m08JMC/0c7wtkIOH7i/llLruc/f
qgAuGHO3Cp6fN5P1qXiOk/3KVJW9RF2Ha0o3AoenLJO5jyyr/IxRgZBef6uJ
TuuufmLLs5aNIPhNXOfQLwSqHKW3+SEsA4n5r87WxZvOE3IrUCansxeYs8Lw
doHdLeLGhvyZT0Lir1JZNE7Nz38mvJCAmTPXdywwsCsj1jU+Ke3WdfKRJH5G
l+2q3mNojCTupEnqbwgrHamhXAZHB7RwuLpJirJlmDO2obCq+mpON+sLJpiD
7MSIeqPxaqOK3fXxi2nD3DjdDosT/n5JgEWdBw9MYIoouKUlZZ+aqAWI+x3T
+unArfOCPVSareDTQFkMuN/GbPQuuUthmi1GBuOtVfor9YpiwlkytPmK1sqx
vslTOU7RizT1RHZCJkfaVoHdCRfeQWnx2Dz1tSFpeKcC1jwNHwMP07K6cnIX
Usnq+h59dJnYC3s8LYt++u4opkYWw6lU+gUhhpbqFogGO7xON/24u14EvMWE
aZV823DLk1HF1HiEULsBXDOWX/tHVUrKCAsMgnsA9SJ6w2eszoG1JAb5BZNg
DtizhnbLMZQUpXC3PqZniARiO5eGRDJiymPv374aO7G389KK35nvD9cOKb5n
TYLF539nWOiWazqTm0ZIKCTwre8BMavVXdDwJ8sAg8vANw1ex/SXpPAuvHqk
32bytr9FqO9IALGpRbRSPpbEw+NOsa89jBP9bR75sa3UqF2ifnXMOBLN7RH6
mOihOHCT1lZ+gpSDPwM6qxngfh5IjdGyMi3OkQsAK5845irwFkBsPkkBIC3d
sSvCHfFYMDrp5jBk7vXWkqSsN/PW4U3n49KCNHo+i4rF2cSOZ5XnYwLOtNGI
mb1fvgN/PRvb0Sz/za8Q0XxbNtKNcn1MI5HmalU+Rc7oP0DENTpH+RDCl52i
N4gmGhC015u5vx7YRS+DmYbx1mOH+runInwH3As9PEEoduOppscM4/YVsC01
IgVzMX4Mj3r4zXKo2KWVVyaoS2EXXQXrlrM9pfLwPB/3H5b5LJtF7tzVkRRO
+dAIvNKgJ+2Rl39oZhTQrY/8lOxQlwtP9cBCzZ1qXJQkhtbJ85Fah+pN+aP4
R9nbytce7nf+dttjawQssq6ryntdEVl4/EdzElkggyduOVlD+BzpUxVr14bC
tae7+XTE6oA66zHs2ikgGkV7LDCHGX9OzrSeCHEQ9inIqJttIViC1UUke6Yy
i1Lgtv10UyfRgkBswOdfvKj0oCKa++MxUbfDw3uHh7gNpTqbabAaJsZMJV1i
t9ZKNenigE4QKMJTH14c1LVmzs1rLZCpwcYw0lOKtIJ4DQpcCi5cFHTtPm7q
TU1PAW9L6r8IVgZ7wZAFtJhwfpKxlw995QMX+KXPS1m9bDwPK7yMcn4iqOl+
CreC1nkCnH788CH7Q45icYADzfcR5iSNJXNMlp0nzQaOniT8/PJ7kvTnqaRE
lUlQ+GS5wojnGfk2SCc5YwtICE9pm2sFbWQbeRwv+vK6t9g68sacKOHm5H0j
iNa4/kOvD157v6c68wg/jVzeh8QiEQl3mK0hxZ0XMyWrl4J+6Xf0lH09U1LM
IKM5ZUnb+f0JrL1nh8XU/BZOPz5Sing1M/Zw/Jg745O7AQqU/1BPHGiyUwKx
WkMMuhgltN9GFFgb2g7gLYcb423rEXhH5gLJdl30supzYgIktD0xHn5gmK0M
ufbMVvo9oUJ+ONN/USB3aaTUom5+F2Tm7W0TrVdqvSOSSi2jkDdxYqVOkv3I
7+eV2fEQUOGpX9d4ceVy8W6tdT/frGZdQmEjUnKlfUvHE2BZMTEPTMKkn7dP
jlrbZhdJNvrkAq1148qc3EqCN8TYKjuQi5nJjGxHrIM27CTFWsRMdhaRbI+E
bMN7LC6UnVsj97uCqdHzqsyYmsXwRVdtrAddv1y19nBM7a/jv3LJFFdjxrvz
6SSFy8/PNMU215cbNC/BdUvR+bE/YWF4W7AmX0FeR3wdM6E/tjqyKTSRP7Py
EKsqjd2tmqMNFUR71lCcQTTirWJ+FpPqKQKNMyC16H1xXLUZTUAbneeiGkBV
6i/mlr5inVEn/hj0pK3cPiFlPZXPJ+frfbuo8qRSVjPXS6UuAwy7zkM3qkhz
He+Ufw6F8FMlTHLLTlwCakQvkxsDNJzEXWmqbnZgM5rjrA+IsTjTjgw8dxca
abDfNr8FNjK6t4LzBMfsPSAtHyiypHmRjzP18w6WoRi2cqS9rSptmBvtiScO
NfGX4+84cuK0HnwlMxcoSz8MdGWX2EMjbKT/rjJUyJMS0c4qAhDWWf8iH+db
2LTXP/0aS3bu+1YY/FX8q7a43a3ztGmXKTJ803Uwxce0EUkyisUCP3W5350e
7WCGOiwvYR80fvzdokmxu4vXZZ87GDMpCKG0KZRblk/cAIKE2MI581BMF/Bc
EOSUB44jUZQzI1oHQrsGxcHK8or4Yu/bzRMXrldb0AO30XZpXLUsY7K42pQM
dGbQXZ195zxZosAU+sbgMSEOgVSvpQ+Ji02LWcKR25GjgdTt99mSuR2PdQT+
zMa6S77IMwbw+EfCCp/wBW1FC94S/SRsFRjELzQHUQNs55QIj0aCVzys0rfm
C/mriMWTX3KIKY4vZi+ejNvU3UrUcxVG1FRCzhJybULuo3poyrPTt9gM6IUX
MBwcDQ7xNbExVsVVjFnLI+YQWKI0l293YXwkv02B5TzOSpNOEmWSg23mEKSl
6OAoIzhNI+fZkYQSHWEH71qenhmeS1h3iceMbxpkRb84yjRbGY2km5M3BW20
Hd9N1zny/ZyAjVEqhkATtoexQ2e53z8yKfFuZgUt0TxKj17iWSvo9BE2U5bv
lg/z9l8wHx886T5JtOn4HYb7wJ3VIWo0IdOy6oODDyCTSC9wWzTNP3sWD6Mt
CKn6JzHu21b9ZN3xwD4vINEN6vFdiACOnSD0kmAiWfIRTVaPkI6XqnwVkZIM
46T0gqgNy1sVaG/dMiKKlOun04YeUJJHdhURt/8efzP21hsV3wHx91+qO/sy
BeM9ocf95hx1M/zfDn5VyFxeGAJva3ilZ4bDxdOlSdBweLIUQYlK8zgU3Izs
z/pXsRGSygI8okkvQZCqPAjVGgD+aXI0FHG8UAbJBmjyzj4UiWmToq+p6adO
8kKjV+kYbhRJmEnu35Gh7NXdSsLL7Llr5Kzff67xgDo1repFFMh9Itt3XhRJ
Qorjw/gkKqb424H7XKV0Z5t3QMZsdKB+CJxJGtwRhOxq2IjjzwmqbxfBskcH
ZX0HnzzvlJRr9eVBiX89UAPv3OJqmky49b3JW6zW6TbLTb3+yfZGyajGiLUU
Qn9ZszLlVoJZCco0ctdUK9xBSff609d1KxnUgVX/djVmv6F+d0FH+GGMGtjl
KZYqRqjMZEFAlwQGtMG1xv+jOKApnM0dz5rLLp5SGuhjOEekVrOXvcGnkMlh
fJOOetLu2QJDJr0BHjIzttF+IxapboNkpGpuz/YfJKdpiYc3i6ODlWxM7SoA
zW6nRlDq9cLD7spzIEEgdH+fik0VyWzgET1XiAGHGFYa5HxUw0ETfpA3ia1u
YXH68uEOskpHce/KY4gFa8YMaqDz2lJZEOpc9sX5APuLIoEt2UdJY2Ku90oa
o+TUktLUnYJ5EoTHb5y+So39jAx7m1QcOZqWi6JzD32X+iV7ZV4rD7ZrUBB9
VK3Qg5Uvf+GxvYiHcEHxbjmqKG+SBuIoR7SKx7TJvmVhfH4AyxyeyJTobv4I
3r5Dxb2PnblbStoBlfXzA+/dnBay2QhMTid1YjpsmURuAj24LEFzR7Z6cNHi
/54tfn9wyaQCf/BrQ6vC/FnbzlFq8UKuQN+paurA11qzNrOC9JOt6O9PLIoY
eXgHLkX6N5m3Ag+wGDXgG8in8WW40PRfUlpKcgAx+x5cKQb/sHWUtjX/RYUo
HTXHWJSZ7CrWsxOaj0bP5WmpD5eyjyQZpukL7DtX1kS7iwbjSrlWsQJNjVj0
AIeyZ39SEWDe/j3857XEui/OUIgJ+Ky6msjXUBS44sydZEzlPx1+PW+P+EBY
Acu8QNXyKzz49UTbt1PEUL85HhBx7WodeqkqhdW1qlo4kJd7BVZhXbdnTccB
DMgTJONr+E6k+G660zrn0iHkC5SoVrAVpvx6GxG+xAOGc43ef1wJejKjOQAf
RAmGSNTShyC8jAXHELzlNj/VGYDUeGVJ1mlQ4cSzj3bIxQTewWO+ZM9h4aK6
M2X6gBC/fGlnLpiTFmlDrTZHYVJjvBY1wht6LqiRpzOpBZsEm1GfhWU58wuv
t9AHNWiXoPmD7vr6UdiIaCi8Sdp7/Kbd+0V28pDyZJIJMrSCwJVVP8WyKzHn
2BxWbzQYBLH/NaxmWOj38gDANQq8EiDTjYVliOw5Cf610aVhWlJbT2eVGa/H
7T4dqTlJE+RzRfyRV8Jkh77BXViISnmUTROexdoo/DcxcAa9IwC+MxgFaen/
Xz2O2Jqw6Zt69qrS6vC/WTcO5akBSDwqLkfxCwfUB5KulKtQWZPfBi30Gmpi
7jV4VRwqIpreopQO+KQdzXMH6ckYjnxaY2MMHLA6AxpMTX+as6VGbphNfZKe
yRQchG+XwFYeuWEbZ9QLlonsIusokLZgJE/l5cG1vHWUyNXa/a8JheSQF8RG
Uug0AqzQdaelHhmtbeP/0KxsqTVqpCiCjjC0rbDf2xK/MAwM9ltD6k0lYelX
Z21AyKG2JGGkKOVzG0kHa7fH0U2hHk0N9rXa0zxJkvCRJyaTCnLOIpDQNLf1
hPF8E/Z9EQf1tgl4hUaA3xZABFh8HWJXYUgOiUO7VJlP3FGTknbUsUK1xmNL
vDqQCVrHKiZ0readAqkBkXB218zFA9tiQdcZjAXKD3GL5Q5HMCMBkoL6/WO1
eXl3kGF1nRGAC1SdumVB2IEeN6KpRpg+5tVrzyL2W8kbuNBFH+WUjpsVkD7a
ylfUfm5KbgjA3znD1xBQ6c2vOX+Gm+q6+CwQPL0OfwmFtg/Iv//IAEdwS3M9
7t4TQnP54AUVVXn+HNEHtw10HX+Is+eaxiTuxLBOia5cSltJ3ahlOCOheDet
GOjMn+xLa4d5EFEgQssg40erGpZTWc8U0JseTjlIV06ADsXU19ZgrAs3TOpA
yCO5CXKLKRpWgw23VmjYSL6DNtdwc4ydhwkcUZ0Q//pld/5IriWHUI7c3er6
pfpJKLhy1aUdPdfKT5TZ9bu1UqZvgAdZbcZICPtyCsb2osYc7+omWaBG4s9u
J4gmtRpbHDSf70ZMBm4somMxarbKuTIfD0relQu+CLRHUkqnJQuwrHDWM3qw
jExC48AZIse3B4O7zWb4ST45Wq0InofT2L56IQGdHhMQnUPPj2TjHTnrGIiB
vLe3Q8jwDNci8VqzUUhv4pk7O17cH+lW4eL/D0ATN3rh6iGaHlZ+bJUgRHLV
aIGziY6rGlvtMH6qCXUS3OAktkEtA8sMiX6CfReRGH0mpWRxep+cxehxLEnd
Ct1pnB+L+kPsUaqmBwMNhWZSZw3n+DgMoqD421iFqcj8C4Vru0HmgLvvyN4g
RTAUAzTe7GQf1ZjtypJ4n5cMcQqSpI1jGsBYh/MYSMgkIqGHTf99/6JiCenh
pG01VYIyohAXHIxpC13RTBgaPrAMJBGCdCPfHmfZOBBIMaTxlgQIVhEjQ6/0
GjJhF5QGjVNs7z8TQsYRtomvXyTEPrIbmvsmempwO+khs9XpIX7T8uwrEvJN
EEDIF0j3zxtvE359nMK/bH28IOL4x0epJ/UIPBWvT6XhaeT2enGPffTW00nu
kkwtjBtyvbQeRTTv3coOteXeNGD8BIAdkXVM+jPq98BNwTTEbGr/AajXXsU6
Sg2di3r5GlXgrVc8fhLqb6oRUV3R5usOx3deUdrjs7MMxMjN7apfqUAVPgSo
haUFynw6IUtObOsfSDg8YJLaih99+PdTy2WVlO5jZDLkyIEhFBvZcGu1E4NE
G/RVFqMNc8gaj7tX4aH4N+P3eAUga6uvnZ2NKYo3Y9HroqN2cBu+Ee+l9TMb
pCV0QC114oE2PhXRW0uoCACY/qyMnG5U3ltDarVE64b38JEwBcYG+C7inqcZ
eFA1KeQkv1LTWepaKReyx0BZ2+wYLOSnv+TPZwfctwlL404UUsAaMb9eu7iB
FlTgzERRWAUd7aA26qmg7udw5W/ADnkELxhiQXRPpr6+HHg+UIxAehfpxmWh
nP06WFt2N2+8XAFQ8M/6srNZcHLb7LyJK9xxEG65LLBYvhoY50E88ynidT/w
AxsSlOyJUCflpuKs4JdVnnCrwFkAqrRw+R5qcXXozI2+FdI7HYjL+LqZ9z5L
/u82CxsfEmDNBcrq0pn1H8P0xo0gWWGeKIdcfd04okl1WQnfrJBvKsOm8vQZ
c6sSjY/kiHSkPLOlgMK2M2R7fX39Zbh5E3YS1t0tM14sOPnT0ZyRy7t+9zSp
myvwaaThD28wyqOLalfatf6B2sD78X0olA0DHawT2AC3tbS0JsWsRL+jvgyO
NrrlJDz8qYDGRt0p0Z0hfiM/99IAo34MklpaoFlC7Bv/kCNZUOgTp9QwuMIW
iCYEN+QFczSABnLs0WF/0MeHJBV4qRYN0EzSD44/gakzdy4ITNp7EnxQRZLF
DZOeVa18HokK+3Xm46652GizmhC8PtkGEGFcep1fZcBKcuZxpDnKGHKtr2l8
cAmIMGsSw2haFGP6uUq4j9ZiMusMFe3JYU95gIVUvAck/fc5wp46CClDFGuR
m9n8eT/AkIC4m93JzamUsOOCKe5+PPysYVH+cyWf68Mw3fT6L2cBEjmFB32d
pLGCMG+xR6YEWv3DWDxPypBp16omZJvY3lAwPEqe9ikuCIL6qz7/Qs4BfT6i
tWT7mudunDqiRU0sCt1fURco/vKnjOL+LdYeNZAEo+lUZO89w87wulyJtxbn
zTRhMUlPGxcHzifxpjP+YL/86Np/ihhNbCQ9xR9rSK4tqlCmTejB9d02w56j
FLyxX32lxxDzscfFA8mYSjJIEHG4ovAZnxsH3NoSKLC3g1q2N7oFqFrkXUb5
H27ytnE89Dc7OGJoXXJ/EtVrS5AMUNDaY5hdxDrBoiFB/SJMVwOs3TFwOkgv
Ws0LscqY4TMJVVn+QIXgs9lUntTZhxCgzWMg+jmO3AVDyrQwOsRAFrf0KYf3
VVPVByqup/bbnOYDXTcumGqcuY+kHRIjrElZpZFs2kubenKZnarcR0pui+Sj
Wb4kG1gFaJ7dt0d/k1tBNLqfRLKLS25nJTQEuvdB/9M1v8P/pqWoR063u0aY
1psA8TeOdswrF1+Q7f24eY98KmkeHO5fD7QBQAuK2hNFBSU8pTUoF+0xhth2
as0xBXLjjYHlOZdV0Z7iO6GIa6MwrgRObEPuPSot+uMf/VS2w/2YFHZmvv9H
+iyLHVZFEF8ZrmvVHb/njTtX/4Ggtj2wfvQsb2TAxbKDvt1g4UolW8JScQ7L
jvhpI3yHUP0AOYru9D3RZNBvuqT0H3fSgSf1hwFH9aCI7CgdWjnOzJzVoWY+
YqUbYQIVKj31m65b3kGt9hOKcaS3voCN0b/ZGdpWiT53gsTT3ZarAjXr/OaF
6/BqYheZxu3fig/Nf1Eo8puCFp9t1cNBhTuGJoFrwolODPcSDRVKQtM7RRGP
oVYB3OkIqh5e7SYY2atQrBFLYaKizX4b28iRs/KxamZgdfLtZ3JG1xi4/c4V
fbloyEta/pZ9NiT1qAOuOu2bY6NNkAMGWa9fYTmyuzZ3KjKtbzSwGp55JKg3
69RI6kMcX1VHozvhFOjGGnQt1wQeq71/ChR/6viZFXfcZf4/6yMJxSCTjs2J
f5AfAZsjH9wvTHsg6r8nsXA9qoordddm4rtfueSKpi2o+3kugOB3ZMtwIHcb
PFFuq8S0xkoAa8t4+wunupVzeBPV9MtNa+6UjnPgjiPsnJZhuKVzc7qcUHJ5
rmqRyTUrblMoMp7OZXW7SyvEW6mfiynJBypQC2bxbSwwr6u/TNf/D7dAYEaR
EnLon7mR//Yd/DnZVbh5VsQWNykPrS5+Sy0PNzcBBaJMW60QTVUH5YCNQCFG
KfBkOCmm+25zcBekX/y2B6+l1ZeFRY2QpsK+rTq1T4CzPciDSSxwonFUMSWN
L4uEf+nq4xA0Nyl6fpbN5cyDhTQxagfKZLLAexB7y3145zl8WVDEftcoBNjk
Pc5FZfdntB5FWsUD3M22i5ZN11kzb2hEOApNQKWMZ9WqolvmuQuuGyV+fAG3
+3VojuUSdEqT3eFAtUtFyB/kaMfPNL0q66q8/kgYKKEkTyzaaAku07RK60AN
e8JDwM6B3WIyMVl19wN/xaACuNccpDVSZocbUTCwp5hLSxYlN99dEouadQSF
cWgrEcnh4Jz9VwfaAmxAoiO5cxwL9eVWjHM+ukI0UKE5BRe/V4ZWffjbzyF/
ohPhvQJVuc3xPYuA9UkojnojdglzZSvv+Hm1poO26KJfMKzRKhCAJet0bgyq
KuXz5vzIdUrFT92kM7ey6izipMSyDivtUBB1uz7SD5TfmkL3ICFxlHoi/8Ku
tEkj/O0Wb2TZchHFdfb+DJqSUYBNxmGhHW3E3j8lkLiD5kl3r8v0Wj0axEzX
KpRJIp+GCzMKy85EEgTeNKXOailwE0E0d9H1bvEargmV5f/eA+X28mTjFNAJ
+Se2+ompDEuOpbNG6F7F4zxCC84MXkyqRcvxoUfEiUne9QMiiyOfC1yb/koK
P1yPFUqTlBKvS8SbY1kpyX7hWQWcpe5qHymCXkXfVE4+QD5JrfcWHR5npuNM
Of22Dcg2Uvt/rC3Ea9we3GYInsy7ycvGEr5HXq/VhO1dfgBSHHZoIJBdRsiV
iBR83v7mBIxqxALhQApZEgMAnAPp2bcINXMqvVx6M2vSzoGU1JHbOjgOwRkk
fTObwcrWt0ErBlQkXtz9D31Zmfjn7Dv8fwT0BR6aBolRrKZOl4t+fkkrEACX
2Qzsbh+mh8/6Wm/R0rAMm9aHtxg1Ks3e4Ahay/WiYlKIQ+WTQHQzO2FF6ynC
HvbdN0AaZD16tS2X5QSLlK7od9huMq6VWkdfEJVjS7hKfN5KKkX3Tm5ZJTNk
jK8tnjJesvhhswevKhSS9Ir4SxnhS8Fq2ppntZ+N1p81TXphwE6NClJmybcy
E7Lnj0F7F5FF2ni0DAazqKY63hshVMudKr3WAr5ScjaNz9HGwVMCCuV9ihQg
9ShoM3aaPEhEUeRWvluQFx0cH+4Cb4qC9DaeVVXAXeINqoajymLEiZM/z3Za
Bh2app41y+AK2/8ii/5n2wIMVY7zfejsk9aycN5cV4q5lk7xMilBUI+wMGQP
RvsjstOFrIUDiZ3A4ypY4cmT1vqlluMCHEC4TcwNmcfnHRyi54SL92fj1CTT
MwR+5BG077D9JSXIIFW/ExC+mLv3/6xcsijVWe7zJoRolrTXvQHB1Dh68nJe
Ith/Kjyusdz5pIwtcwMjYgTnq9ja6G37v9dP3KqBzSkNh6wCCDhkZcA/kvfV
lBIWTAWifdeGqosRtevnWQ3RzQ7HuEzYcLj4gwVqRBy7bOtCyrWMoIvAmAvv
whjSHzl6b1v/BEmfZbINFaQ6xugfSe9zy8NlPdxvBncXlGNlv3vbxQvcOcQG
JJ3bVJyM/sO1FiKAo0E66Ic/8Qo9vs6owwkzd7hWja0pu1z4HvQFIoErbFKZ
MEPSG8CUgS0jYSZPStVvygbdVFLczIFngtngJtU+rUXb7JmNosz0agTL3MQE
9Ul6R4ZOklqRGVMfy9yjosupFFd6ZG/877ivZgl/mNMpe22WPOuGCThQ2SLT
6dr4bGqO2cohuGScH4zXABjV4PhgMqBfbW2F8K9pjXF5EomsfaiHZUXr2pWe
yBbdd88YRHY8r63gGMv8Mmp3uRwp3QP5VfyWrkIcOOha7cUT6sEo4E/ymbht
QPdxBw830qh7aaI7fjOLjTf+pXnY5afBq3r6bPc0kfvETUhiyhGtHlOYNQJg
S9KyMd54pFLFV1RIb0+dGDQFcr83Mph3t+Uzlk4BkkXwpwrcOx8pAR8UtAUS
pJy1gMFFqrbbgljI9+sOYmfaHjBLLb+kHA8llHBqndaKjtPWKrIxRiDt1lWz
kIMtYcN2mRDqBm5zfnGcwqmxs5C7nclg3K3mjMVUT6plz5LqUBUz4Y0+QLjv
GxJP2ZeyFZZcA7cnFtbnnE7A2r5DKexES8hZU9bdD5daj0KsgvKqdG3sVSXE
oZRp+/c+Nd5ogCjC8w1QYa8K3VJQ+pOzDDCL5ObpngTpL8sAv8CoXhd4mVAx
AvYs76v7iubeGag4R6y9kjBHo+NjJom0Y1c+iuhotXmfgVd0GNerEYEQCftr
Ptve8mHZD3gRunAIXlEbtndhsCjdVoxUpVlysnLkD5tbOUta/QAWsdj/7VXF
CbwM3lgRrDqlwtmX70iMjHQlFak5m3yrxiY1D3ZRBA1gR6Uv6dS+zAHIi1Gv
u90SpGOBkZaTHWkf3ugOsNmraDK5Q+jcwYrZMDdXuX5L3Bgue5uv8hFuKzxB
x+nTrNH02Mkv2DdzJz1zYSw7xdyVD62xlbz+STaafgKW+Ys1+Aye+ukBAFUg
zekCZsXw5lWMBQjrhmim2DXOQHIXMjvhqc346vHkHPVWOiO3YfmUYVj3uG4x
LCuQrDJxPs7HEtffy6D8hlnK/mlThz7pwXPmplHyx6dDW5XNE/Ohtm0L4KB6
Wv/w2wcdz8NOyKScTLOwXxInqFcYzvkRRHGF2ODa20NypcSAnKeq4mZmQOrU
JnC4kpCJCs4tpclzCzVGCxCDYRa4+jigFBfWVbhJ3S+ybEK39qX3xsiuy+gh
CD2fhUXSzLu3BVlkOHDdSgzxQhBKem3AWRKUYwBe0MNV8tYEcRDwtHMCVpQ2
pthcOBEFOeuS1FOo+BwgCTQ65yQGklerfDb6sJBXVhCZbVrVqBWYEc24DRyr
c8YMJBLrjhHtJclyv1K/u+qhIrP6tDiT1gYvKTbUVvP5D6KBz5FQxOMVq8Ou
t+HNbRr2iX503p4W+zbEm3RXdOBJaYk0M+J9EYNC8dQrcvnyJKdSSG63Mpey
DkmFP5V9PM2SKftiljjtMnZIR2fD7YUO7gYt7Ogsd4bAR9IitbEPFGy7c6cx
JdtGiu1WQCozkT0bj1/wHyWwpsj+EaS0CP7GdMWGz3tkAUJZiNQZXYbkWfBk
4WSnPgkwayl8rtLg/AfiC8tFoeGAj0JqFuVl4wSho+DPz8qk5weTWnurr11N
ieLn7BrdvRXiPBDjwXu51lnbTAUGgi+n8tBVhElrih8jPCRk/43wDcXaUwxG
GSdLVl/E7+VNM+Ri+Gg3Dg9yFjlBVhQAxWCo3nGSqxPCpmfTmJCnswnOgFWQ
AIQacNb1H0myih62U4f7Md6QVhKjjftyIfVs9vB2U91lR1qhNk9zMhdqNUZw
01wXGrfVZuyQYzG47+ajID4H4FQwCDk+j7U8oKJ+zvJc1NGnSjgbCWTp4Z1M
sqQrCVQBEISljK/NIsj4q56HHA4o1nvm4mxainsouuXz55+VpwQfrhcdTUOF
GARoPXyboOLQNy8rReCb3CP7yaUBl0XaABkoqBWq3zBHmqpBmPICBE7cdVua
vrAQe1uBc30/jyWMfkZohKK/DMAvSeIOng6BeiOOSdg2d2AqAPjpQ/Awcpi4
BkxhkcQHQav45hAHJzjJ5R79p7avX8g28MN5M4CPAgBPZN4M7yVTW9X5TLqC
Tw5xjP8ms2sPORJ7jgahUgBWe+d5L4UZn0bsWDtnDzMN9WcjV5GnuMN7z1g7
nFNfs4eN9Q0TXRTbw8z/LA8tSytXLg7ASVp/9FP8kRcDdeyi92E9qzYAh8np
r02ljUWzcSCswdVtcmbn/UPveIF0HyFazA28sLyCabffpqJpDSuXNmKitAWS
yzLBWbS9Kq0JYGlnGB1/qAvO/j7BguHTc7X/d8bbFNju2xSk/8+MEs3A7z5Z
dEQCgLxhKdC5U4N74qXkApIsPhToe3BIIG6tJot/RVXX/2Vzh00wofts+2sJ
R5/zi+A4n+xGcI18LKA4a/cbrD/AfvvP3E/whullUdGWn2t2+nXMgvQYQ+1k
A+/YhasiBQc+sFKqmcVBEWRCvFYdfu4SJ5dkMIUnWdBLf6qfVqB2/Crhpxrr
Kli/dpGpUS1hderS56BdcGu1A3hgJaxvzEVL5ebWE71jZfrxnrvnB1W18T+W
BLP0ULWjhgvFWi9SkOGC956UnbyDKUCD4uDEyKXdbPlfvudBkQWuDtqDvaHe
YcWwByeMKpIVYNgShP1tuw5XxpNJvWmrImflm29mD+V0TTz2JLqb+T+9CYpO
SzzJWHu+j9zZCaDEX9iE+zeelJE0WBtlhgxXKmS7Jt3Iq30VxSDAbvWVPkkx
6AnnioK2v9RaiKyxyQ8jZ/myfnptyXXfHBCT2fku7EgBBdqWi3cc8/pYf9ho
n1w4B5Mby+WGi5CwLgGF4XiLpGOmR7GpFKLlvhdlGvMLpgC966Ff7Us0yerv
fIxMYOLszaAIO61R0uZz7xyzkwS45AbfKVtOfTFMJwXZRqF9kW50Ur+cycxK
lL4ua/ywIv7edT6De/cF7IGBr3LQ5LpSYMSqr9G3ySmcMKgFDkm3rrbKZy4i
p2ndYgZZAIZkXOCkGaf/d/3D4YEn4Iud6YxQfYs13ChiY7e0FSCly7GZOvxO
f7akQ+e1H7/pt01fPOB11OtSwHOA0S2wroo/ODYJXAI5xcvp13zdVHCwUV2s
OJx729ZZHTVzpq8889d5uVeUezgmwVsxrNdKv2qCKmgPu5mhYfaJTe+Nn33z
iVrhonPFRSByeDVlTfVkLexu8qJ7faF9njmTrMgdmF4Fsmt4kkajieaU7SLq
BNBRJxV59b8IiwWY0ksOsnU8mcsrnYaJJANkWFxhr6dzLXkSQaPZKQrnVR/u
ebT6oNuU/XacO2oDTnktsSyWa4DDqn47UkerbshPT8mmdPo7V0PorchQOy2g
3eUvVqV5BQlHI+Nuz+jLDeR6FRwGDT0mHrxKLjrzT1Lu720LO17/AH1jBV+q
kw7zyXYhYT/KR/rnEBT0WC2dul+jevwU2DmkCQBd0NDgpxdGva75shSHqzx3
DYNxD4jlVkpISqvxjN+mUBkf94q7X79KBrLD991JEnzerGX6KDnex/QRR9DC
WOmheYqqFjhWDRmv+9Bxql6eOPa7mgZrUGaLZnWucHeKyQSFDwkx8CTvIkIB
Ed9NUkQJBflrJ7+BGPI6tFFOUhzg7TaosvepW6soqoWKaY7NuGs85skP0QVW
s7D6IVOqdPC98+28vX7JOOmFvvKikiXboQcYHnqm97n3IX2eeHHk+8GUcwDo
5z6i5TerJyqd9dT5JUfJwtvOk4mISoLRSlEe7gi5aRxIbwV2mWHFPXgmizyi
0F0yXqy55PML5aOkqXzpgN6GTAif1jVn05R78/XB12G3LCy5L94ClmYeG/9s
pYHGGt+9dMWbrMpJhDxDLFpDoWI8nFoq8z5pNY1u0uNG16t+H1p3WVMTsRM2
hHb+/pdaWoK7CyNlSXI9SF3h6RwFC0S8Kzu7JvQsKsb7thMueQDX34NdzLOG
hI6Kz/H2MLuzyi3oSuMuwNaOnEfr6Q5p3PIli8DM7Dz2jbvkOEE+v9Rdbp6S
zk8tb3BCh04JNkuVGvKSiqNjAhCX324/vEb3SyWXjI0hafmMrxG8rZEA5bgL
qdH18xaQ9E1FpZTSupPVDGgq4Abnqj2XLxQ80ykS56Kv/Xez2YD1mgiOMONt
RZlS6dCUYKH3jqV4PcAxwQaPx1+lq9B0n85aJWUNX+jDzXtsSGM8zr2VaPKH
qJ0lu6UfnrjKs14QpSn3Wi4E6/IEHmCU9u54Y+eO6/y65JM7C5rzIHdfJ0Wq
FPOLAmT5gWhnVX7ObRoVIRunMG87KqDZrATuwaFDmnHinleQ1VjrPYXstZsS
sjArGZzAHVnY+5EozcdSXVWXv6+GpQpTxCglAl1Y6gsYXueDVNW/mHcJ+1f/
iafjjJtQ7z9+OCEBoVqxNcTP/PNA8p4M4ne44bdriqdUmt10pW5Ape3kDWn5
Ehi2SxfUYqBQ9ih+Rd52GHzrenSCFs/d3dBk/cXxYwDBAtvmW9r3vPiU8p5M
LPY/IATdwEgRerqACCQ9spLfB1mTPyrPXvb5iYAQijKwS/KSQaLCMyyUlomf
mgm51mOZAotui//dKPEO5LV+uwj9ZeBT+gcgUu5XtIT+cMTsKEXK3rngaz2n
VfwjCt4YxP4HW9E2fyHBu8OHhsZLT2wbj9PnUS9r8R973SfUrhEkW1z0aYTd
CupspQSBjXBPvYbLNEX78VDjiMFG9XDhVsquxsrfXxzjWei9Md3yJuaBvnAL
2pKYkCMK2iNoquU9vA8piV5oel12rSIPeNsbP2ORxsjDNoqNZHHNY7KXJTl9
6fxsiUSJ+JoSKPoPxsujT+IN03KWzSK6Ru5qcT1ttf+S59wnvdgd1IDXcnIH
8JzPETboOQfnJAZzIb0+cKWWZBFh0LnxPnOdPvxzseV2gQuSpymF3O1C56ob
a9qlfpIzeXPU6foNyLCJTZDaedPsCxhx1L1O5xTnY0Q/t3/HxW9jT35X4IwE
20HW5qSUkVwEZSsuNXVgjY5DyHezG75OYKmXSmULEH8qyY8Pg0w9qgTi9m0h
2lUMGZwm36rngDzD+LLs1xWGpkNDbviN5kxOL16yVOpE59h6QclsOlscwnFS
SwpKkDw8H3zst9Kpx1ej+9MJo0vGf/n8Z0MZMzultDpe77f307aWT2n0ZgCp
afrL3lyz1SLF4X5o95eyL+FM0ZBZxr4C1YPY0XJxR65nfVjdNDjNiB/Zz/KL
Psv9HJ4GKEuJQox+LIgseRVamPUDn3h9nu5Eug7iXJ37hiVd/SUlwrBddFP/
CZ7xSChZUgVlAI0gwaSvWmkiP32F4pRkTCQ35WHsJ/ZpND0UUlI31wf7gIGX
pTshswdyQqn7ZPWR3EnULJlvFMUdZsXXP1koe0Hw9F6pCpKTPgufipXX0jYN
Tp2GkuKFwQQ96tGjGJyjkZvTYXG/Q9XKdrUrI8LVk+plLG9xmlwMSnoDAC8f
BbwBOmOpgUrxJpf0Pm8d0uhqPBRVsWZG+w0P0qUZTKoCpM8QgHTddD4b2ZA5
HBICRZJS1oYPp5jN7KlSJ/rtq5vqaQGWdSSZERj836wZmG4GgqSSI84ZWcfd
Ph93o7cQI/vGEiadgOEm9EfQo0kQrLHwzaM3Pfr2iP1yNOgB9Z6K6+CnTT9W
dkT90ydOHX3whDow5JCrYcdGeJuX3+PNeOvdTcIqX2aFYgnhMGA0+Q3rPvvE
y44kGXltRatxeku5TA+sLzMRarovz5jmTunX5Yac6ZWomWlWBiNctmfYW6yt
FXOZJRMK/RoLPTRBMUdx/cHml7Jq+8XknmXSEtAr1uxWJBYBWKEn6meBcbNq
Sr4u78swWL6aXedln5s2qU0hLxNgenMzFp8xdhwRMLxpXIVljvz5Z/RhxaiL
PNxRIaAi24/N3F2YELu6S7EvimP6kgMURNKc9owv4KEIQpbfjsnA7+ec4Gdh
W9cYoT14wuOGJiQjEQLFTagegGua9FS61cZQSLYB410CgovUy7nmq5UR6cI7
eXHLfNwCjdN3uXcoeEwvOfgAieWb8oR41M9pPCh51W9TDGMFK26Aso8M4o3c
CfxSIIgwEAxtpphH7txwsnSQk53kpJXOcQKLfRIN6XvThJi3LThRKDa5e2Em
yDKLhWxASsPk1ihfTvnAafiAxEFQIe1TGm1NUkqz96hAonpyCQWbBNjD/nIe
8MzMZZXpR/ZPYN5Z6fG/M2L/iI+Z8VkMx1rOwTmJbSmK5VUPD/iTzetO2xO5
/+OvDajMO70SMZl0XZ2VwVut/dElaMV9kOJqSA32E29dI+qVvEOUo12wZbDl
gTO2cB+tuV4quMozvCZIEDz9/fMFdbsGDoJcYVs8glyN9M3cBpVCTrBKEPPP
FK/dsHlYHmwveGKRD77fOOe/XfHM6fvBTEx0jESnM4XJ42r7mh0Y0zEN+CZi
YAESBNZiC+7MwXG/maReYknWuQo9ZMhtwpunj07uvrt0ccyzQu1TJU9X2Ofv
Rh1geqqR7KfsUN/l1NIR6FekCwSIqKIe9cAsMfHFS0dXUlhY1uHAGR5H1Uss
Wl/TklPGtLZf8xH2Dtjm76OH4wxhkhUIYzaVHryfHXHx8ikAE8fc9YyzwmL+
Pw289WKcxKsOH6HDRxr7IGLwb+ElxfN4crrWzmbYi+0lSJJl24TrlaHbCRcw
aL3Ld64320GQZDjayfGOeJImC5E7JVZyAZFfZx6v9bjOjeBWdS07+vsd4mgs
rUprrA/BKZwxlZ0N32gtPhWQWeV1z9gzL0TcZ2rUXcYYd0zwg1VQCivnP5SG
ud2E6igMf00rXte+GVtVOitetCiK7V7f2ZYx/AuMWnxJFCm6drzVKu4qmMz8
dcR9IPBMO+KmfV6Xvr6Tnyj++e8ZmW2U9nYTmQqp2fQWOZu4H/LIubPgFJPa
MJmVrcM5ywkpm0R8q0PkKkXAf5/e4xJh/TchbXHSjLjmul29EOpCOgdZxax5
j/0qvdJ8pRJKxfSY13PrpPUpzERaRX5KwPHefUUeK4FJgU3yOcYWbIt3PdCP
OJ3DHa2ZP/ZPC8bw2hF1uNSmHmbaBhTVtgTW0m9JDnJZx6skUWSlC850Qxg+
y89zePhXfUZp3e1DeQvqAh9PJGLsgwWgXrbWbi3VXMm9mM1lGNKssJ9mgXRw
0ATlGqt9iYmTmfNMKCZhduvUDPa0kSHZvRXl+ndraCoALezLkTbRVdDD6L20
lTGBDZQ0+kl60CCti3cGxrVTNfnA4ia4yqOWptSNRfdtQVabt9NTuSFamKMU
2sprLropJW00erKPmcYyKeLLkRXTlBsErACL1pAfeXhTWFnhz+yMsC5hRw76
omW36hNV5VDrPCXeA+tLdmPDWgqCFzLmU9uQrt15cp53UbUiy9Ox9k+/kVb+
BfLX4otdh/1ffEtxJlfft1erN4VrjRgjKm/HFQRYTfmfbuquC6OHW7QvSIuD
2eMjtBAvyaM7ABJzgL/9dspIhmGPzVjmgPR6t872U+okLEBiGG1SlEYMLMC2
KdrFFrsGmqShnl8XbBfw7eO8DkPrdjh7qekqoGninfHTTsuD0JBroDKpjRl2
CbCpjIjeDLRIIIRbC4oxKxNBxBze4zVGP5+4sBXI1rJJqSToSsOGsEiGfvyQ
bVTl7hgFVz/18akke+t9aRsKtBL9koVCXrq+jrE9VWNTwtdH5ygtHmDZqYFf
2ykTCadmq4tMUk1nudHj92WAvS8+/iAduM/PkpiHoeTGB8f1jZuIqMcc5qjm
f7uLh030rDuAjvB53L/MeJuKSnY47jYSr7TK/ldyJF8BStGsBHKBKK8PewCW
2NMASBKSTh6gVzbuwSR5Z0MKmdE5Ry3/8eQ85XEMzXkMJgMiKmndW4Of8CDG
aaFMQt9CciGsfzJBVcZ9OlpO1jDw2bwsJjGNA2JoiBBsY5yOmNOdHK+4LliV
/+HbQLlhIShLu81aYCNBBjx8MJ1v8XZKEqjjiyqJ6X4SFyq32Yl5XxscYzUP
a1YdFgxVbn9JewxGOI1BDwKF51W/YyKYldMRX1EVbbGwxcBF2omXhesgkESD
wQlbj8WrVcFP5BGjWlDaVM0G5Qf7is+UNTpgPzEstu0cJ5p71vWGceT1nGaM
iABkcVMbeP4l4XRq7dBkmGXnRBxgqjGfTUApZ3oUAgPFrBjvTxI05zFbqxdq
Qmk8SoOF/hm+U2MzajLOEcNbQXYuHLZr4Kz9iWJRRegaVnTM5HP5Y3dCvGcm
uEkcy1h2/6O8HF9/bmnO6VYz8ViSWJW6SdZ6zncH+adW6jXx7RzPllxoQzEM
aHndWePc3ohlWYfiG7WTFalqrIyjXT7ZwWfBbo/iSQYM6ogHGhlyZLtdiGGm
DTlHfR0HCNL3UCbdZToIM/HykbuXrCKKhOZn7zpGCKKPqo7HsO9twUSVnGSG
ceNWdEeX4IF9r5aZXU3mxn4wkneBnyAiqJ4T54Y5WlPDhzg75KG/HwdY5lzd
8sSLG96aAeMQ5RP0tk1wTtk9wzV+CQT4ShXOeDsMsMPL5UhWbPG15KhIXt0H
sqt6rDeyGQnMHCTgmON72axaQipm9FarhkXAHLWHTnn9Y1k69aWKYUhDKo2n
aBCh1CLNKiBeIe+sgfQRz1Jhq2osPbWBo/9KKc9R0DkSRRHU7XPahDyDHPes
Ee0bdXuAxBEqbMmC1wbDvEJq///rF9BXSu4aOg0Azu+vopWQ1bGzU0XpK34b
QCEVGpGL4gGlKq5MlTGK3z9FkUxyeOkj7Gp+nc+qOl6m/EkynWKmVPyzccvv
3RqkevRwvPTHmtwDtb65jojav/SyxxMuqMyg1SBgt6O+bmVkX3ih0T8424hH
9LjZ8ewvcYigdFusH8xg4Q+hvMPcjtUAMst1K8t9TC1zB2yb5iD6hm3klVA9
98BaBino5cnTJlzglIXwojyBV2KanDhxGPDqebmr/jrBSAUOJ8qiY7Jq+Ait
3TZUu51HmFW0VsnAC8DumP6xQR+NQJM30NzF9CHrmcJBxFHn+5DppYsBboo7
PJJf2hWhjgIdkBo4q3ybAM2JcJx5jiOhWClyX69oy3wweRdKYMHWJXSU8Pad
pO8m/4A6tWLEzj72MQpy1o+7u8uh0YGJtlF3ZhGHvagRaVCp9BN21GcLjACy
UxBFH3L1u2nK8kpUOL+NT9i/OIRNY8WknJCFmiXAzBunK4xiwkL48tZa8mH1
/C/lsMMqxp8VLC0bvJnm8cNnkGG7U3Qf6TTcWHViilpEsBox33BGhlfqDn7a
Kx9JnB7UZIZygD7kgXTX77BgMZKdSNbY5r3mykUCaiejEh8OlMj5vtsQb4KT
/jrRmuuFjvU5EpWHIFrcF99sYxRiByi4yN0SCKtM2UMgSsv4mlNNdF94w0zG
VZ5UlXIEXqpTrgyWntPxtF/UaXZR0arSrOG7Ml96tZ/c/vOl5krjmnYA0Icd
eXjHaIWrKbrzzwQt4ECy8V3xaPRKUQwtmoh8fNm0pcBTxRhxM0vFcX+KgmPV
omtmN6fKhtvv+019Zeog4lNmosb+pCx6T3VQqrFVOu1lUt+ZFWvDB4aUxrU4
HMMlteG1zoXdeS/JX+AN+Ixy1q3QAbjXFhWIKHX7khhC0dW021wr/t2ZYeTT
NmETnhucJWL763QaOuKZ2IJGhL68gTNiKCeAZfi7ELnvKXZvTPll3WkLAQ4h
1zQs383vdIS0VD6gVNY6ECBKmVwweQnjqPbYj0EcDGSyF3MwWgzE8E9pJH26
GPUjd+5Z6kzhDCByLgHMqhTTPP36oIyoKx3UTE7dlVxo/bmfnF/Q4DdzmvHd
rr9I61K5fUpME+uvZZtNtX1OH6DiZ89TA3x8xYp/XUsYqICVPkdAFpr0CEpz
FS4JQyhzlX0sqS/IJek9q+LWL4yNI2nPMXzWVwmluvwO6mj91E/Duc9+56BC
JweLry7KEuz6Mb2piwuAIk4vpJl0YVafQTKx9Hj+xSEjZrunYboSIrSBxaCJ
utEMlJI60g9lGhZAKpG6qdgJ/gqD1RpAJiaG+lwVV7zZj+GRgcvrvo7w04nk
4CNZPeUgtmNKoF1h8s8TXmrEyc3OELPXgJMfbxkrwtozWIHDIdPUrVjB2ntT
r2BLvg5KAofysR/hFaaahlAABOUYGkqv46rsGNT89//GPHS0RlYH2VCUbYZ/
R2t6wuPnEEm7MCorf0K9124ARTkgSsXAQ0praFacz/pELkViBisCpkmtWpFe
/y7cmSWji8yd+R1sIcoRTFh2WnawI8aLYY01cKEyptiUwjtd5PHTUNUT7OfP
EsHGYKaTlIRCXnOwKjLpJinHK4ovWovm/+YiGCsLkZwWIIeijeh6eW3uPvXK
rUFh9oQRkIlzsZKPbk2DxnpjUskq5f+o8TUxBYnqMZl+50C0+hBQgc2OmRJW
i4h8o3qIGUJvMv+uwAhdekg+v75+llIyIhdC62MLe3ZsSgKoS6m87C0SqaIs
XA1hoJsPVEw5+8bNyQzeKnHQ3G1+qZzaujgBmW4bJoQQA4rvyv5rtzJXRjzN
kxZDI0o2Ivnppt1bZK4u4MOdqQJwRqSDmInEfo9yJ4hO8uxHSJrxcMDX4szh
YL/B7ApBuT8hqxUhvvnE/XDMICrqlLP/LxNeaXvO7TULXIGt8+6IfO6v7rPY
1Jict566f0D0/m880KN3srOVHXv5vKFPDV9opQAr9bu4H0++gI0VK+rOQZut
pAueoJXd8+PCFqJwcGXEVHJa/8okKYpD59xgnX1oM6WIhSPpS1tAAaGcxGUM
+0rEI/hKDH/FC8nRAzBVk1pPeWnKN72BJLA8jczfI3PLoB884T1AgyDb7Y/a
b+gmRZLGJMuuJAiPp14KSczfAMx3Om5/iEPpxqG29lSNLxgIIzfrlG96aqCh
KW/mOrixTQBVFiMHm71IeNnaGhKNAcUauB8eDsxRkvl68PGZPrDfKqxZ0Ou+
suToE7XWq1zniYr9jF0s06pI1W6q4Rmz8YAAa+jbJN4O+8bynB214mbTETHu
W441nM3pXYTgN2GQznweTe5HIWOYYIqVrHG2e2XR7wb3AelItAo0fmSj5SX1
Yf0NZQiHB7uKTN5TrkF/RfQxYJKios/lgH49w7dlNEFVOI75TGaUxMrigHla
PTLxIgwkE/optbSC4CJgY4GKz84sCtbrpefl+xeOmTmGdfhgQlBJkN42MPld
fYho7gkgfHSfTR5wGhLLjVWuhGNzLAWgY9buw1EYO0Mrb/QN+btePCKTvKGX
CKiizZ6fzW5bf98AqKsnxDOAXyV0Bt1yPxoVpY0OMSo6ZwvRR6Fo9q8xhAt2
HgiSPwa0kFxG5U5DSyYTP8Rupu0vzTog7lq5qoM3WfJmNkgO876vk7jtypZW
r47Sthc/jQC5egNnMxhUI7FiykW8AZGiryBVK1S1pAYo05j0OXjrsieNiNIl
Z5zFbuwwzBbcOYJLaS7naBZkHgmpu2EdW5BhWEOWhdCSgp6lGN+jx5Z3aeIe
5tNpk3sg9njGptqCHFpg3x6HTfhqlbCAWyBpMqWfEsoiz/D80RUDn9w6MSVK
rBF2xck3R553NHhHYmMiKdLS0+W3k4N1Su8uH/GIwQhgew0K446NkjGft7RJ
yMSjmhLCxbfg+WRgvt0j42SrO10SQGam4sZBFpqQ7xETrsDDWnTfY6KIXZUz
0+G6dGmF+1Ly0ij/WAQQI6uh5DWD6FeleLPCy4SlALankYs8b2mY0gzbWv1u
OJ3wXUxU8UYfyaqWM2QQu9EN90kCEAcPl9wVtmWMGdBB1xcL2fgplRYI8ggr
PzxTJE4hKSDuM7fUZEX0Ad7m18KQEHVeGubfXFcsJY5WyXAiPtFbLijILUQU
vUGOBYD17giDRKw5Q+mIhLGh/QRd/v2EPIt+u4LIgRtTNa0E5wENVS9xRAqg
fWkus39GpPF6JVtk5LAbXrR944zyjDj4AZ6Ddl9ZkFpeQC+ZbYKB1KcvAK6C
k4Yv1UBQaJdGw+SNMVenGaOR6PwmEsN4XrGkhFmlFXZiUlIVrc535V5Azped
AEkpMVQNTyd2OYwU3Eijjmo8n/eSjaX4Ux8kEGh5NdXONKyDiIpiBqWmiaJK
CCrnbMd5zJNqttdlfNRZ2PnChdB4nnbA+GlqCtvNmjm8RDnHlHRyMx4y9TyO
bpokfD96MFugpUbGQ/xzHCBQtVFPnAIHHfle6lvcZnpWU56TH0AKVsoAPuUZ
FrBIG7ciahxkPh30inh/D11RCCjauDBaoZG7cOm2O5TI+X/y+SWs3jAm7GN5
aAQeavX4lNW+GS4wR8Edtn47iJq244ctMxKm9lcmXhhSFL4aKS7LwTxD/3Sq
gPCGyiTCuKIV7CtUcruPDHcsFIV9VJDarY43mYr5Xu2VZpcxRMq2DPIMyKgL
Dl1eL1XY8bpnMtGlVti2Ryb5ed/ULgaBqvYAwgZ1kN9gS7SMjUaS+YZjdrcB
o9eOU5NsMX4INZsXxf/ZHDJ13EE2CIUGxMf/z9gU7GXWK1xzIu2MM63mul/e
NRlJRm/qhX8WCitsrl8XrcmS26/z6onb57HZ/mXN0E5F4dhfqJKRt35441p0
pRHYkvjsXse+l8bZ6FwoYbxp+FpctEBdJ/rvY8PWaQotLbjOxQts8Hk+yMSr
FS3JRtkYbLhi73z2SRrMh7nfcx6PJxN8hFCGrmJBK5gKRJ8drqVqQJx2j31O
njAIceYs9pUY9Wk7gxpzciDwao01Z41RR97O8NJa4WUP1g30F3jNgGEDZtYy
ECPauqowkKlXY7R9TG0YaJOxiiaNtdFoEpsIUEzplOcE3wfHo8KpgfEU/Wzl
f7pBsNwi9OdmhoMW4/5AGhXiFhr7D4na1ygrjNgIjy8A2WFdM4Qi+ntvKLFR
ERvjXeXYXKZ46HYGtuDzjoTfkziZRXX3kxnYQUljMgUBDEO0YlQX1/knGxzt
7a58WLDmIx1wPjyT4PMsPY/Zv9qU4Np/7lMnzOBKkdYaD7VwN6ITsNGr+ocb
CfHLGmeZBfDMu4NxN5CZciYP5HlYYHdVYgueegCapwbtTSQVI8+vggNqqVi/
wp745AKIL9OWYYmcbX1zw9uium+Eq+499coRzJsfEjFLz9EoUR+uleVFx4gj
TUG8bt4M85zpmWKnrmJC5lAGkM/kF4U+yaUlXUfTyGrLibr4/Z9SBLQU03eK
P12Dv0xxhAh2nYz3lm7u4zGiySOwi9Zih5Ld6+N3HNRPw3NrAQtBg6/6YyJ5
RJy7Q7732+TJ/35GJ0Ku/3CXXETwxKQ8WtjXcL5QPEJl4k2z82vG28gOXGw6
s06O5sbJEaLIHGbbqUpX/+ZR8nl9s6uAW2ihIWrhjTRL68P6wQMtw1uhwjam
RBLlexTa2COIIGvjhM5Nea9v4NqGyxIH6qjG98GsRrgsBQiLRirXLogR1t36
SGREnxtUnmrfV2AyEcsqg79ZnfMattxrQnAnN4qBaLUQo7Pi8DCkY9FLeWhZ
eCffGITfDTEzu/hsNEdt2CdfxjkcDddf71OI5YaIpgyjF0kRd57nRg9AIb+m
9BH5HyIwV3gFRxYZa4x9tC1LbJ2RVxZYwDmroASL9/+VhQ2LbxIohGld64oH
qeCFr68OKamoj7ynBuwVRBHo6Df4NVghFJ5vsM+/tiVg9Dy+QKFQIIbzCqKO
cSwz3+0RETYlolmDrooYRLMiUICiTwdx7rbwDxfiM5pBJcWW1Z+2sklvz2Up
GCnsurmLIKiJljH0DfhcdDcIhrUp2OFPURyvruUXydjdtq+ATwdYoXntMvSM
cqMRlLU75inmPY5IEKpD+lsF+NrwyGlhGDAYSBrJQmcFEzK3cSZSBTJHLj5H
Hw3HvsSNSAlqB5MEn4Z/1ouXw9zZdnTxyUPG4PHCYa/jorFiAj/6OEAaZPGx
fZkpgPOlwJwAqboKdKRwjCw2/bWp4AN282MNPfrf2K4K5WhJiRpuo7EKqE1J
mHgmrUWlsBSz3k3RkQTy7hBxeI50nkijr3iy4e4h1TlcBCNR1UC1PrtlBPwn
mcMC+o0VirjCNPJhpPugh+1iQtLP4OosXJg0+S7LKU99LqIJWdT9dikjR7CH
0RlOC7FjRz+JrS2Jxeg0vmfdAKF0qNtAJ2j6kpFUVEkDcOGceHjMqUwODH0f
zOikcSQl0qopTuf8CSSaJfPm/ntg7UsIACOr7v4aaBdxvvPU8ka5vI6iQUkd
+ql9iKDLktIoxggcN3O5vnq41UUME8YcupDvQXOXggUtfBH/Zb1E6+49m9W5
So6FHFhaHzOoOaScDMLkMD811+3jqqSndQC3PgNKWsPeec0nWgmrIg7Pf6SA
kb+go2d/m+H6TAA4/aZtJjC7xJWPV8Y8V+lz62vcmmAGe5Ro59vWIqW5Ndnl
p8J+YICSDoQ6dfd+fnrkVzUDRQfE7YaHICjPyjFfdc9HA+BKOTC1IKF7YIER
YdFWSTo+KFYgeutgWUd33y6qD4mkvAFzTQhpuR7mv7Z9wo88M345ZqIgirvX
jxfaejqWlYKsM1IHDfrb++iSSp8tduo+kp2qjHyUT8blEe0sGqEIPm+tcVeZ
onxALHTHUv3ZCnFesDW8Bb+b1gY49+X6yaSp5i7C98iGwtdGhkwfHrpjctxP
Q2L377nh33HSPdZLuUDJzcbUv7/1l2X8mt7USbvVbfYpP4x/w230bjpG1cPc
wDCHAuac5vt/7w1r8DVs84sg++iIcdUK9spHFd8bkufCBVHgyyDgBV1XIVT4
Y//dojRpjas1JTN/rTO6PwbnNWGvbSWwI1SnhbY894BkZzRn2bEz6MY6uKPe
Lf3rdqbqN1dgT+VHpBFYmKT26YAifprzkYVcxPCBYT9so0XzYetxT3Srdo/P
eKguJO09RVS6qTh0elBy1cMYHcnb+/HJIt12/WwGsQpWIYuTu6wlzZFwPapu
e6l/wTjh210Fj81A8pDJgblxvWlas2plysoEoFMaINAjPs9Sr6SdS6Ul1/hQ
dOrPkCzqbDd3jVxQsDAApEM5eV4JpMnq447BHP4RqFGbLFy3jyP2oObv61lm
96dOzgKuCPWhgZmxyTTzlPs8FhLu/UWiDXFO0p+THjUROCrPpAFmpqwCX6F+
qaIlipQNx23V4urqkxpvsxIJo3ph3Eq+fYG0wkoAJmRJM6xXuPEXiy0/F3jd
PcUeWvZfRIPJJ0p/is/YRKi7+CTJtujXXCxF11tuTh5Fmowz14yHD/u/mrA6
T3vKfOLgD5+7vxZVaxCIjya5WSCxfLOX7uOvMNnPEv98zZI4QgQUci04aCDE
P8JtFSN8KG5Q0XjXAzqV3IGeRz0sp/AjXk5Zl74BpC2ZOk00uDjJp6q2N6DM
/JkLwJkpeBJimahPUj53ZwH3jkbgYBwlVXnGq7V5xyV9J0t+PbuP0DlhHKhe
Y2q/QvKk4ieTZ/Qws67I7EbdnY7QTTgHLNUGytwnTVpcrEPx01hkSKT4Gyp6
t23L4P9pk6izk6LTN3pmflDBbs0bFAiuhHq9Df8g4BkqLYa54iThIVjh8x4v
bF9p1+JdIn9obh8FTXInwXC2giGaztprlvXPxZ8N/UcL1ev1PKGuNgvDOeSu
LboiU+Ws7233Mx+T2nXRbdYwZmaKgG3hs9vsqiRQPew66KHkZnvI6nE17g93
Z84Jf1vuMNG03Kea+/v1tFSnF5JVj0BIJuBxOuf3CyYklq0X5K+oILi0qvE9
7hTBRv48nzZWpBWALATGZ3elg8+6ZO0H2PElwuj4iSH5Cm/RM/Q89csuC6tP
wdT8B1tvcE5hxkzvfRtOBtxJxKym4kGhsCYPXHo4nzrUcye5O+d8ANilB4Sy
2IlRUmpncug+d17zGM9ugUCKT/37zaPmuhuxVbAG7ehygq/STuDTOZg+ngn9
ci3ndG9BG6qgvnm8iBtkEzuWOn3Jx8B7ubpovi/EuI1nNjXiM3/YHVNk4m2T
poZ4PFx1bhrQc/tmIendWBpz77wqVEh8x66hzXl+qX6797KDVdgzZd7Wv/Rd
Qv3DYlvUQREctSBbGqCSs+AJFT/UmtmosV9uUyAjLBNMeIzd63OlTjUcPeWu
ngfddFKt9aD81Rdyj1pvPJfAYkSkBdf8Tah+YBtPB9vQdvC1vu6N95oGVVE4
XTRHIN1rqVyGH33QHJcaVY/Y+Es/mtWtrYyqtGzBtmXbYKEagdxV0/T991y+
vURHjU++yQXjnDqSe+unCBvBhYfQOgNiuRLG6PrIN0tuxNk+easaBBL4MRiy
noP70jw53qot4oXcRiAnBquHQc5sghXq75vdbqVazmK1hfPQvEfCsixzRfnq
eg+6bsfm5xnO7EMwCbazR8d0LQNKCXuNDI1pQbpYeuMnuzwFOqxY651dGr0a
dMsscssdXHoK19QZRddfM0XNLC8akRrbOVOKjz9jn41T38/VDWsVQq8HoyTI
SBGufJHgWhojo1lJlRuh24vanDb8sejtHC7y0HRVkZvT5pCUrgDIfn1Oaomi
jrnZVwv0C3D01lhMICUM3K74I3cVTsih+7UegUZ5wnhMJln2F3OqASndCI6b
c0brXxoS0uFeQ1Ut85JnR3J5RymGhtZRyH5snmtC/qiFwG26MwKRlgqFJ19H
5HLixK8lzx3TppAkY9QaRT0yWA5+w+D8h/NU5lLJUFdaCaX7ONBCJWIBZc+S
1qvr+ZVWVGFpFNxutQ2vyTsfFJDcu9HBnyC2ql+fiUjsxPnpOZhzaSQDNeFN
oQ0R6Aj3ybqm4+XgqF7J+YpWTBwy4FrHTZaFErju7XSAg+o2TiBbZllVavet
KZiUvhIe+LS9sOyNY5PJ/rzzffG/ScW256nsUk4DksfyQHlw6zSQZUMJ0rqQ
sysDzc/CtV1UCO0vHebgjGGTg1fyBElgbOds6IBCYF9weR0sG+Qrb7IxkLke
ZSKHLssb/I5ECZB8Jr/9QDsjPflryHNuVagKm7CZAWH+rpazHZP9+djvG3dR
f1bOH0wMgsnFfWK+Q+CStC1bRpmBpO2jXCbZsXHbQYQirgK5RiCbLVixhK74
KLDszUyFduJElKKBXW1clpwA/rJZqCo6eG9UnS1ZXD3bnqvfqLj6qZVX7wvL
dxdc/UsYyhZFkrxKpeWOS51e5hjwBpQZQ8IMn2uiB/pxTIQr5OLFYn6/BGXX
KlDJ9K13osmlIJX497HMByHMResdK+Vzcpz5YcYrokvkoz0MLB4W/NFL6g9G
bDSovYTG7sJrPD5uFs9XHClefUs+ZliwkF6KiRMgxiS1nrUV2G89l30PpFKr
d9BYxGa3v5z5bZS4ThuIOidCeipeGkxSFpdPJypjY5gRfKu1QtCXYJZeY+RU
f7n32UQfheNLtudCmQWXqhbtEgmmJ+TbLA63ez1KUu+GrghHrNFtq9QewAYT
eYyJRLNIq3fvexUGcLKwG7cInaf+jKoEO5gCD+M7dm0jNsqIXUlAolFXPso7
DJGYp7fbFrSC6aOEPoboviUMnTMiAgleIlBvydc+tCjR/7ANeld6eg2OkIPI
xKyaLr7esCn1AYSkchXiqlofyrZCo5C3KscFqW8peu14896tOxm1p+YuZ2ew
/982rgtwGTrvv8/bFRmzT+pMKopBkgW9nANZPgHvaVVjR5h82lGJvb6T1BTy
aWAbn9Fn630RfznQDxmPb6BIAmy7BJu4GeMduEGoQv+/VJoaUQQpXZkweD1j
ulxoumL8fBmAosNR4vqiVlqLAxJNrVMjuXtxHu4wVXtTxcUq4XTy0V59bTxH
SXnF34MjSSqMczET8seWX4n4Ez5OVvmRhfRTSmMi6mRMd131EjdvigHDaFTs
tzG+OsTa6R0z7B/VQTZ1w8tqnRmesSUIRePKD1Fm8tH5PFhnAJu3sVg/huCY
a/rjpKWpSiI5Vbi21atPBWd3PltpFV2RH90owywOROS9PEU+n5HrJhi98fvk
xvxSxpoJpVXYws795oUdXo6aQUxGNIzTO2qFlO7gmMRurDeDeke/zQHeItkB
2foTbQ6pUeGEEO6ee586DZT7CmEfW87Pz2dyqJHbuPKiLEfeKHnDH+w2f96g
5+a06pB0iV+eSE073iU/Ilfoc32aX0ty2p2BBoRr59eoSdGIEXlGhVVoyV/h
aoshhmyCKIioJIVxRqvanrxoaiIum64u2aaqLkPeodlhYPiNmuzdh1NWFWTD
hN2mj1/5uDJDGX3sFAN4+MmHznaAs3VasSekRJADS/UWQ96ZzPRoU8Wjqp3v
PTXpwRXpallzk8MMjr8S7X5KrcLKYfcemaiTY086yKanuW/SVQHgKMHsg49S
sRmPb1LwXntYl7/biAbnnHGBzEIiV6zr7VZKYFor0eell6/SDgv8YBT+sNGj
eTVtV2lkAMgkOJfYQHTZXsYHJA+UQZHetL4pA2/Se350E0qfPOE7B/57tJOR
U4P4xzk1cgBOl6+l7AZlOi0f6a/CtQjUEGYhl4CYR9WstGjlCkki5Skn0DXU
TXC/vBWnsa2FAcMZsX+bqQ9VhbfYlgrOgPQL6ElbyrnISWgLMPovTvyBSyK6
tC0qSuzpYpDwWwPTtatPyuGE4Eo+UdX5CO4a2/5wY5YR2bc0HKRKnT1BXh2o
A5uEBJ9TwYfc8OlUKlx3Rm24AQhtvC0mogAyWuJ9x/JlnLHGHnC14wwI384A
ZcEtcvsg17APk/1vMinQbrl+XhYBw1MZV0dzEawNt6lUMcjKhBz/l1h4BySx
irOMdIKj/p1Nj4VaVjLs2jUBGmjbaTDCphfpvFwwSn7qOCXh1KWTigBOTsYz
cBXoShLuqj7YrDeRSi4L2lFeaiL5+NT8nl1/LKTJoureXDssCUXztXKK4zjY
90uNb+X2jaBS9lLHqVvTOPZbP3jr9DdNZOgvC5BETgw8jZlIr8FYdlmxLAZz
bsoLiG0yT18FwuIklDQRITT6IwxPzEXVbEZdsl8WtJC6phC/g9JT5XyCpKPp
t59ZrW45V+BFlcXGl0k63TF4DYjoHeAgDSMI9F2QRmSYFd6IqGk5mJA7DXGN
1spQeYMsY0CKi3iAQfdTj/xstqYfI/BRZCNh326GbIEbMDdF/0NfJPGeLXY9
a+WwVX1BxjlgKvqsYZWdt5GCTbWihWDsc9xeoncc9fmGATC3X0NZt1nHQV1q
91vQ/hEVTyMqTdmuqimEJfZ5pGnCzN1pcJp23ol+XE1QlWzfSzAgYfsrNU9/
L8T9XkcIp6zmrCkMQ/hbuGiqX5yjriy8l0+ClKjpzqtqHx0+JVC1SpXPqDND
+MkVMq+P1AFc4OEVlju8+uww3Ey4qe6pPwdl+7GrNwpMII5bUVG9COKglh4d
PpB6dX5OrqQF1RrdCn6jnrks916CpQv0l7WOfNpuPWRwt3xiSWlD5xUE2YYV
LEdMJ4m0n96ugM6jBB4Uy787muhRx7/8HYjsY+xqG/pyt7y6bFSqwbGBwtaz
trRh9RsLaKhhoP1xK78f0V0fkrxHKoWse+QRd0ux2nQY4OxTxupkapNqYpzi
ybjZVSuIxblm3qPKVe/+PLVYYHq0buVUHhAnodwVpYbaL06mzeUAS9Yf72L8
5MYwGGx3abw9uVOoSEqaBgfXIibJKqnmUqojFHdSVP97H00KdAvvZ1Wy7G+M
g15NPv+50QuGxXAGZjVJnw5y+x0opPnX8rQ01bKi5alkqnK3dnGGa5H2fajp
G2lhOpztB8dTjfNO/whb/1jVcQvl1A4mzqpJgn0jicKeWCM6zNqzXscBNFHX
8h4V0SW1NQFmDwqpIMg70wL/SQgLUelxEB80aDD8NBprKQzageNySZyMSGyx
wl6BXJxunvLCgewlCKi7x2sFWAjPjm+qPP8U+1YC3bQya4at9dszeKc5QFuB
3l64TY3yfd/n8kZGXLvJv1u+BjO06c+gY/m7LUrN4bEkImuzg933lqtgbsMD
TjRmuHVMGaaJWcw0MnqzRdFHlwFRsgsM2VI6KvGxJij5GpftleCGAUt2Pydj
/Swj4dsTEp1uncGO28DRyB/7wgyh4dUrZiEM5GrXBC7B7CFTbrn5TogfxxTP
VMeml05SFupRaGikFLAHasGpdoSzJMm1SjjiCf8KAV/p/lEje8Xn1pVfjLp9
+l3gRJk7wCZDW7R2eS8VOjekpFe9SYEcEDO61AMLLd214urv86qVk1L8Kg2T
vOemhUfdqFfEcc1UAvgWVNO4DYZ677J3P4ALBGDxBTsTpJm8m1DSVBTZ7Rcx
sFMURCD56gBeuQxnUnCuWkaDjr6Fiol7Y1YAmgfzWCqQob21N5hCWlAtlaTg
2985EtZKnaGzKAxwgMSKn0FaA+q9esdk88aR4V8HsXLg3L3qzmsQzWj6FmQV
ooFQU3SUCd33FYGiXoExbeYYQ6TLhbLQXcP+Q+aMMGrCdzVPhqrEJ74443PE
xbwFQahK76mwvWoQZjjc8fUfZKMatJx5+GWjJUXPHuv/owfYFN3NViH1RY7Y
Yny48sl4A96/hnI7igtldR02wcQZMSe8JDoTw3dDCnZCP24g5EYOG+gDKF4N
FocvRidXut+fdnvjRfjC4UpKYXQVBl4Tt7A3RloODb2H5f3FH7d0jPGtLkgE
yKNFWC/QIYzdl/UtzjyfjjTPqcTcJ3Yo1sXO8DtHVA/JjpEUYbagowQ/BQou
kHWYlxErrLsYnOMr5Z7BR/r/9JaNnsN7xvpStFcqp3Aatt/lQ0XeuCeC4ylH
GV5ZhclrI7imykelvAp28xnQ1sCf6xdz1qcKQM4sMwQg504wC0xF0/cWSiUG
QGMwgkzfNVNwKRPlpjeqDq4Y6e/lQiuuHieOM+OvyswUsyUc3Swlgf95rYbQ
kbpgmngBpNc1jUyqBwClAeaGjCdH0nrrieYQr3rXfYo537DTEVfDJr3Xzakd
QYpCmQni+MQjtEBeJ7rhxgqwdAf5nief97H5ZVn++yr9iH1aGsqcwMnWELnt
uou0c7iG25FCiQoLO4tiDkTUJF60Zaep05YBx63TAbovVbnH5CCEsF8pxrtU
FxcDg+iRNieYUMSJwIZAYPozxGLae4kkhrnKZybzww+pXQQPnG2FUE5ptmfc
xfga5CwW3vEB5GEAr1vtzRoqWtJf2oKjjz7WvQy/Z0s8J1/eQ3/g3BlzAxSU
WQhHvAWw3SfOwAP846jz4Df6IA1tZ8TXIVugCt2G5uR19kwYiMlnZZfIYmA5
h7pUhDpJOeMQzpCFI+cf+xUKKUIH/jmRCurhYWalo8SONYGZ7wnKNOs2CLWO
Heex8ggcflwPow9STA2cSVWKfH+An6Ua3Z2giS3gTqaIe3Cz+K1lv1BPwWzn
9pcKQHjiys7lRF5H1iBL07hLR8DfYEIwslPPXFfJxJ7KEzL01XKpJGL1tLwl
MZQi6lQ+9M2kuJxTzU3cmALe2D1XULDrzzP3JnTWEV91tJ/RTs7HZpJR1Wag
X9cXmd8rBQjcR14mME4phny9XuOXLOhuKEQAxsZ0z7KsXj9iK8KxESwcgMgx
szW/NoGjPfpas7hB3sT75ee6YePI2Q1efiKrzM3SxHa0YvZYX+SzypyzZEV7
sNdybxnioArB5l7aj+GSf5G6mHESe8aCItMpe0IU6EgRmIqUUtyOxn+1EaP2
PTM0f7EXuupUE2bF+aT4TSo7Nnm9Dm7c1C6IFsEzn+PPhWGsRW8KcfybshFH
p3tEFygplj8HG8AtF4sViqB/TGHvx+XrVQL08zyOmSbUT4xD5a2nbunWu/s0
pYHf1DCCfX8zSMBRlwyPUR4WUDJ2heYqUNswaqFW54xOqWx3y0a8wWoWBsCU
QCqrImsQgCzyFfnaFIuB8FQVO1tJhr9aP9R33zZ0WWJ9kRHrcORPhE+2WFyh
QD42YoEw3nJorhv3H2tMiNDEtnOxHcnRDFTqPzahEvZpjv/Gk8ilLy7XKqkE
XshOn9YBirsGL76J+bbTaA4ZznzCe3DOFs8+UroogvSFW3QZ+yFiVDQl9wm4
OrhO6BimAM1oFWY2p4OLQypbI5oHY/8Qyt9LAW7/Q2/J3fsz/XrH3xqsckvx
6nocV3m2nosq2XDHx9H/5VQAjpc/csOGWcTN1gyjplCrMte8azPlRe9nL6cL
8kEsrFO/tk+8jvQHuVrjldRJpWHH4Etfykh7fa31+0dHsotxAbZwYB6+8oOW
kyc3N8mGZI/tVvO/cT+zfzC5K7DqdAnqvyoJusY4Hu2BdXDCtEGRRF46uFiu
1VhRBPuglk9xoBKLnDEbeR77ZSxHnNsVwdeOvdA9fHSbBs/DnE4VTtZ+qau/
OtL9F0PAcZufs73J7C5w8Mld38/o6mEnusMd5m+TfwwDwFq16KzMI+ap2jkG
Tv1VPUqlPjLSfoRkuFlHX6e4gzBCXp+1jPwHFNqYmlYUS+pV83g4uNV0FF7O
49yc8v5Wv5QzIVV9u/O8tcosjO/yOuo8Ny+OaEMhAPnsNHfmIpAB1vWPvf5l
bxuFKmOH70BLEsXb12ngGhVzwhs0zPvXUhOG3FXiiEWGvuOIQB1SkdEtqWCu
YOiX6b0Nu+Xzddrxe9Lr8fx93/jdp4YSh/nfUX8V1XTmV8UqfMimi1+h5x1C
ydznvA9HtlsC7+WgqGaP2Zf869JMMg8c/NyPvRxSbPMntGvDtlhkmb4DE13t
SeP8IT1MgZqTYW0JAL7gJPzx2jqauAJrBRJhLnPuPsJHaG2DDhUGdNyBQLJy
65n3ZWlryPJi1nKn1W0HAjqbifzy4VvC0Cb8Y25UWTC3Ts3xpd8vOyv/YxPE
TrFaI736VN5//Apgq3TKmCbXUjUDVRwLAEGJ31l4hM6AG9NsrMLZR29lyF3P
OGpJOKmvtZc5zFonhdEP7oEnyZ2SJcVZTP8nS1Se922sbn4NMSp+g8DP90fl
OfZ+utwBeSqPGF7oPmceAfKDNhkF2WwT+DxBAHcWJGQRVf7iZCifqp5Odn2w
vLcpvdpWzuJwC9cQBMAJQ+txC7lsj9u6Sc+Aes+DM7d1YnmG616cKtPr9zOO
yTw2Kk9zHimOLRyxW8LhHq3mLcVpUyBKKPmAKbZ22DLAxyi+4wJk9JGlmM9x
Mx5GzRLsb9FoDiqpFv+l7GdWOj/gWe6jk59aVVDxVLHgFD6wJacYxy4DhcZv
kad0hSWGJbLj9vVl/YZgNWvz6Wm8wOSlOlIdrG8hRCQwMO5EqPjToQ0WyWmV
YZWeIwbjdKWDco4O3/GMeAjmFvCtVMmVuDbG0Gh6r+f4jQFjt/wV3iA35tVI
tsSSJd70YbBe2Cn7Gd8kbo9Cu5hxEotxLDXMS32188tUsAOmXJkViyeDPZlC
ImOuoZtdaDyZNcgtadaCqeVR02qJ5QIufOquEU5CdG7BZVEZOX9pb2w3jlFG
dj80mPzUW3mNUHqeYaNrjcxHhyGIbBtQw1PyQaoUFgO6O2TAg/rN69kv05ie
V0h3+gKjEYJVbyoXBJsAYy5kkw5yqHbfPWADOm7+EJisu/d1B6sanrnT4+qu
ul5my9I1XjtKC3Z50MkxKybmdZExu+31SR0IKUFLJ3UScLbujWpkAGOuUtXM
jHhPzicyXXRY0vkfB8rvykfNQ8P+Rkj8zjRJV9i0BGmh97LaxaHZETsrdRli
7AurZquzc1bpvZeu9IYzjlYPkNyyWKxgzrOdYN14nmn6ayzUEG0JMXpzkO1X
Fc697lU6Egv07O/u28lCSD5GbIq5G45Xd6ENqbHkJsf7wkM3alFPOP8pFie9
KJk4UlA4k/9xjuZjQ1YeAdUv+YWLAV81maMJaeoYIw1nHTidaNz+82hgSSJD
AEWlSywnnuM+ER7elKCWHKtFp2bMsZaB7rpnUGi7ZfvTRK37IZcrTM89Oblb
oxTAndIAqowTBI3ppcI+Lo1M7k4dQ9vy6xhnDFQ8wvuIQfKxSZtRLpyUUFxm
uJUAeZCQrQ7g7fQZ3CiHwrBGYsN7Wg2RuSuY5W++Qp9v+yjyDwqXQ9w8mxDi
6uZbBuFrU+lNgLDtCRSDRdXZI2MyvE4AR52qdy5DnUAmOX2D+K6CZeA8g37h
XlzIBmm68JhLEn1CPyMM4vS+h2LIR5naDj9m+dXhS3CA++Y9Tfg8i+JCc1Ec
4TLyvhpYX6zClbx5STwVO8nPgEp3gL0mD3GAfTfz8kRBJNpGFk6mpt1OcQx7
CNejfCCrFRj0DdKhRLpR6daY+GgojArNIft8c5SLeJ4FDbuTFUf6bvRMglq9
GVFZyOcuvmat3/RP5KoyFA3rR0lzcKoHscoT6wlNJqP5Ok9afPYMTK392Sgm
0bF8KMzaH8wcJFwPeCpK62ureQMgQICZXF9NyCKbqxsqtCOoYg54O3iVEDl9
oa9Ehd5tTwDsoHnEpWHtp6WE9PgDKQK9wy23YtiTK8+cwLrGYWTQm5HIpjzS
ga6+HJ7jzWUD7+OLSD5oLUCdjbbV3QtvhdVksASXHxupKeRf0Rkdzxdw9pYD
rNrXbUQj5HAGHfDOvzXABDXHR4PPIYSLSwzK/FrNTYP9/X16dSEcMqKuD6Ty
GUUaJ4uu7nhM94Z/cP0+IWgSjD/zfqlyorX4TSH3Uo21HFr35YOEQDrSsaJ0
JLWJf2cdQtb36zqyAE9zeqLWbd3IE9t3BNBgxbSmCfwHzodOh9KSZXnj/geV
xVBLhqkkTlkfz/XtCGoSOFXU/dKd/fbnLTxutPYeKldGJF8TrhAWFvUlwxaT
OVIA/942UzMmMqw+sMj7Bm9khH/cnxRh84gHR8/ncakGor0Bz66WWMI84dy0
wEmBVFJk4OWL3fCs9LWPZi1iVgox+G9Q2wx0F9JLpg+2oYDPm/E3ECjHg8K9
hsf5nkFtZbOdkVxXVnNisPDKV9m57OnUpFrQ0uY9jwBGr61+nEBYjlvSX4W7
cTM7mldaKWw47b8nCZO60mRYVBHIkwnlepgKX2cqfASYZOodr/pjkA25hZfX
jN0Ll3XjDmmeehBs6TW8kz2zCHIFK5oJIbBVOtPD99Cn3d4pzqd+YnlIKHTh
cJ1VNtk/L9SnqfwXSCkxSXFIm7+MMOE+aGycfjXsjHP/rAIut3xZtQ35kf2w
ja+GxBAP4cn5vUNQHSyCbvBDpE50jnSNvwMhIBbkPbYdg/VTESSin+Mpy/Gg
yAf/Rn2T/oPvu1OyyC9bemDUGF+3PVZ117G15QS4mccQMRPNQAtQual221tq
/j9onBnzVYGRyhXWqwUJP/YEbA+IkicCfovo5I3YZEOPyCKXPgf2r6XQnr7H
47SXcjRv0p7F8H9TitKKTiRiWE2xyHMV+8gqTX0fW3ODW9LFGkQ/swsOSyLL
iCgEKf3QjF+gaA3l1yc0LF/fg+nPWzH58vF/IuLJdr/wZnRYiG0AQQwgS/vq
ZRQ4cEK0ylXn8OWsxsN62jueTbZAdILydnGkviU/oa4yJQ3W6IhLU4agTOB2
4okGvPh4SKhUceoNXcqyCMbwArgk5VqQ+ejmon2eSqagjbswGvEhfCFrF3ye
Y6kkv+BYEdaaFK8mTv6Jblrf35XF9B6hVyZSbtDz8oG5WQ+OrFZzYAc+X1ly
ud0haaM+Jb5zLViftZLqhjxpsDfvsgjGjg1NlMRCgqtMVfg/AFXVfxpj/Io3
fMvwmpeUxrEqW18vG7t0wIfWM9PEuBR6KROneXeGabaVrU0q+EEav+aLukNR
VZ1OWAGVSOxs4yIdjjjeoiNinutwAMsr/peSeQkO7eE0QHZe4uM+AJ8ZATJc
mEtZFujoPpg90+/Te+3bbR4KyEhYnUlL5mrqsZmEkdiyelKS7gStHfBHWkGM
NladzqkNhOxE2W3TjmpD+Aev9XPEVa83Sa8/4isKABUCdBddxDhi8mNCJr1N
58vmhWpMg5fYZUvl5zHiDOu6d9wQyFzYob7iUtqPEfIZOSvjHvF6c6UWxRWA
MPUsQKnNBcrFKwtlRj3+9RpTcmru99PT4T5jilDKXTwF6OdcLrXWn7kIg/a0
LfY41WXF6vq6EOz7oiOuWRnKw3B99qH5CYuHnOvlGRlg/nVlgy6dbopD++Ew
kPn2hNenYtMty2HbGAAdrismXIqj/cyCSEY6JVSiEwhxdMXo+yyWZ5AEZcY1
qUMO8VVa5meiyWkfB3OqTmLWHKdQZey4TKNTuDx/a0jcivIdUn5fgqnflegg
tM/+nTPiKe7mpTp2OE1wobwZfiZF93+y3eU09gYya4Fvpgom7dg7GBLqqADE
aj2fB7JCx+UFuVBQLACy3J6rVTomzyiRid5cZqSvMJBzfi6Wsf35TqkJH/5L
XzMhhAgWxzkpVHvi2v+LnjKnNOK1q340Ah1oYQr/ZOZNYlJbQQqaP+/DXqpq
wY0hfjt8BwgarzryiBbx8I3JjqcPqKmOK+nfGjDDeJ++H7BHs8YH55JeIRnf
Fsvr2OPyy2iICXKloxxJYrdNY3/IBaKF5t0a0fsSwL3HjgkQ3DJCMK/T3I6J
DtUgkf3OwEYQZsJSi7uZ265qtBHCEFJ6gGCcyq2L6eWA6pyddADSoUnK4lOp
A1lw2bXC+mN5bSQKW6fv6v5CESXfhgdqex8cPWOaX5QxDZYO4/4Pw7w0VjF2
JH5W9IBl5tX8clVCEC2/AkmdzUQG056OS4ADdi82FobGAC/MXMLUK7QMKV9a
PvwDr7MlGzmm/GSETkkcSpCybRuB/PzSvY9NbShh5ksoO6mF8nkXZ+OeNKIE
oWeqrL7OEawYXm/Pj10qPXE8E4gU5uK+hi/DMeOxO7LavjBUa+w+NgiRrrGD
mNbOW9ImyyhAR09Vpf0OvDG652r/7FYtAeebRHKraRyKWMvo+eMI0SNlYjJ4
GgABSMhABEPyv9bTEK+Hxl09SfThGtjd7lsMzR2EMEN0HRQ5nTcrGKn5QzOG
0MT9fevvy0eubPDXU1mAcOT2gUsKfsftejzbllsnvRn5e4E3NGzmEjmjsX1t
NLlC9OrMKCmuEvgHEUYZsPaExO/CiF52dw8K+Qg1rYFbMi3oZa7uBDHTFpnh
GEYimyihLGmPAHqb/px+AGKaoRJfQin5Zdgtd3pQ0C4cQj7hpAnvI7Le8Yny
yeLc1m+D9lAfvwwWpb2NbCbSu9OfuInr20mDpBHG3exRvmboPLMN29C0ITCj
wq2PM9jC4ljj3cIa6zWYYQdiaJi24QzPgKcHzsiHIKTgKGLLLNQAgoee8OKk
BvuO6RVl5f7L9XwOl7EbSHeuuGq1fSJyNSQgGTkwjxsH3/OLal+ACKSXH+X9
ukHDyJd4BVdcKctnkK7br/Eh26pnmrrwouAeU+nidrJY5X2a9b91IKhgKkg4
Npkvd0DTVXkHZxgGN4DPkZXuvESwz3Enn28wphsIwNuSkCARfyIwy6bn7wcC
ASvnuTXJ1NhaHG3D423zynO4OL2a2ehc2ww/s8RRW8Je0C/0ZVZcmWao8Ljb
w2XYzfVssRfVxdfrJDw3WXRQgBtPCudQJVnxcP4u5HYaf8hVE+ntRRBC3z5n
BDPr5SuAAs3pAuz4l4xVtXP3NQx87NUB8RM7feE1kD12i2qLXJp0ms5zRdWO
ydJREGf0hkFdN0OG8DWXrUQNDQAb6PeJg2DIMUVvksManc7iEDf2y4BHquKZ
bq+y+UJS7REBCtQCM7ZWwRDgEz+6wD2N/SEVB2jTEB7HINVMU6GWVYUvEtHH
Ac+EMkpQS+1mUjzpDOgzPdCr2B1jVgrk0T3CkktgHBH0eTiI/a2zZIPvVG1D
ASyrxaPYrYdqUgVEmoClpPqP0H0FgbMMliFD+EL8GBuTnIxOm2cZF7Klt4Yc
TWwXKUtNObcLe4WWYJClr9ubqwknHQF4O7jRLGCZ6XiZqKnGb2kSkrkHPBs4
OzTNrnrh2/zUIJVIhVRtT2CLgcnugL5sKNdS0t0171tKLvxCWslgNLEr/6HK
rjYyiC7oSzAKBP90r6PJyDrRAwEQsUKwT84yYeQzMDtnWmNR2czyJ+HoLBOY
CsflVjw5B/3G+47NrPcvsFo8JxGm+02l+5lt8Bxv+bQu29UbjxHNnod9boqi
QUQ2j93GqSLfw/8iePbUURWZxgnugjBJBkmZ0qMasLlSIZth7jJMcXosfarB
12UO76dhuniQbmFkmFnTA/9B/zwBzY/stfWJ6gtp+OJu3039NdWQDFN/ISsB
txJA6nzjEqBo7yNwgQRdN4uJBo10ZfuIzURVgnuRK1luvUYvK9aUdgVriw0Y
Iz/R/I8H2W0k/pYTClH8tUGeQHAGxilWsTbxQ5vPMwNw5A75afRGenHv2AOp
qe7JMf5Iupd53Wnp6YDGQUN+Jt/zewUPh31UupxfH26NgraOO8R38z3QrIg6
95JAIkHlTyYY2W/wufDDCaIZ05mHBEzxo8Ag1QbSTlOegr4+zWfztaMkkiYW
2A1SwaaKRS+49psCflZFEuo7pcPhSXdHKsGswHzxHzWirNlFmkcQBWJZqOK1
/k918GAOeC0l3b+0xKngBjd85i+WVXWShpPXE07YPVF/u13ghUD8sZjk28j+
8jw1Ml8SsRRMXiSJ93YvhGW4n0QBxHALru0Ep8PCqByLg2URqJNvOYxsk+cF
RdJs36OLu4hiUTUWNjea8UMVVMeXHElF0r/DdelsCU1SFQPzDj+T3/FZ/+d6
6t5a9BWI6bTOvsqqYl7cAU4rboAm6BQlGpvJCjgxgbecAygzs4ge+g7mcPLW
hH8TZMMjXv0lxc42SqcJzZtQ6cRdmJQqO1DbFVU7Yo/jL2kz0m/fpJlnLAeD
/CTPXkJd7SlEetLDwGzlC3BblqtTBljMpnW8Y54eHi2UtU//V6TJDQu/NLI/
+XXMr2KkrIddjGpcSky0kkr+WzWZb+PmdjFmkxdVOCStfW/OhumS9q/UDFZj
3jpuz0CAlFRpkXTavd9kPusRi0tcejKlDM73AmEAKbKU2s+L3FSVHlDY+Wtc
qYGA2NWfPcp/hyomtyW7B2wyyR0A+LAkS31vtGCdhCleOuIVTx2XRgdIPd5C
+bieM60m7Reanfo+js0s9eIvNA+SYhvtoUndi6aT+krDNzcCY8UYS4T0DFX9
X+YgI6hxATX+e+EXbmUFZ/c5gY/KOhdGucwJX48SmNAvmnM1Uewosi1fRNbt
3Re511A5xjaDzl2lk9L69gCYhYW76fISvTJi3fDDOLrzhy9NM850TMKw0v4/
WoJVMBujQ35RVmtM2hIJf2ZEJ4yr6CTtfER2TF/buTq/x4rsj0NQunT+MVUk
MOsZ/OK8eomiIHcrwBj08XByClQ1hvInk3L22T1+RKpuc8jeprCEF1L6sRr4
whhSbtd51LzcqMztAVkUqy2hZ0Moob3yhd7K02drapUS6q8EQAuS8egghk4z
KGj7qZQDhPcho8weF1G1ynD790tdZmuhKZyJJWqci4RBD0nS41ItQnBhHeex
0y2mrgdoZy5cJz18DfM9/K0VMQIN36oSoWhNq1Ozqz0k/QZJ7UXPharQIapg
ARVUFWhATC/6rHSi49Ksa71pt9LTmFGPD/KaEEeeO1y7nHB5rrApPywjSUZ6
tN9C/sCFo9HupShQJ6mOjdkN2f9uXi5wQNONXFSePib2i586Jl3t/Mo+xWN/
HeL35UnSGPnJQ3iALACqw6Yaang0JjXb+9ccDfgrGzvJe3EB14nPZY5+EPOh
cda2qa78aK5d4xyUiAqzOvxkeG+nhEVObxgVx3zpxp4aJz2FcUK4ZsXuamLS
VGmwQY/o76I2XeOc619oO4cXuYt94wJrfpWvrkNuA/YK5VgBaPil5GcOtooh
PeyKk82bbaTsI7jtQBp0NqkOr7iEP7aD3RloGSS6uCas63zn0gggr/89UdyA
YZj78B3ZPEpjXMDpa4F0cE37iQKMgtHkY4tYHck/E/pBLMYO1QTSRhb5vBYi
j21F1fVx1/mHeZ1XOwLNj65pu/TJ0YLO6wU2BrIuhP9NwRx9fRrWRjzACkmQ
yh18kPw5bwf55Ld3uOA2ht7QM6y8a1T6a8bLFEim2jNOz33oReFGMVCA3czI
6gungCh20V1y8ZqEddkXqLMnphHi4lyg8shehEk1KImq5g+jg5rl8orVRoqO
im6QEJAbmK4pizXKGg99hAzbm7ofCM+N4obwxJs2xRLfDVEu6iybw+mzfRmN
N2sVTDemEjAudS/bYcU2GzBca9fY/N4zJa5P67yAu3plDHI6HTH0M5EJUpFs
s/45p+RDrZJzyum8niluOx8a106385LuBEqXTL8f3KrrVBbyv1L6i8IiJZxU
Cofn/RhfuLH5tCKGZ9ZdrK20QQ6F1YH+o74uPxn0loC8xDfG/H7C39KfYl9g
48hz/IuLAXQ/9+7GPN9uZZ0s3S6H+E5HDcPajjfkg16c1q2aH1R3s7RDyvn+
XcrIcG/Cbe44qil4Y7jt/hgJsx7WsobZjJRtjrUiHv0Pc+Z3KKisszwUOSyg
uvUjJbohQlzY8WEplykpTDDtRDQJW+QeBDwJzjAntaZ5xIwVF9W4AKJnMPQo
SNODi9DZiXsPYzHY4mGLh/U3e7xDAQgMbjz/v6wEof5liR+P29dyBy8IQpf+
HcVhd+lL4sWFaQFDhg2BOJlTlq44rl5bIAYW+SkBCPGwGuxPi8J0pLHDNvcP
CDpLtxHTp4M93epsdmLPJyYn+JsSyRIRFyVnpdOTSdd2BqzF6dR1vlGBBIhw
kCwMtE5guNZmBhVExC0cmhR+98BG+e1Veh/VSkZhpTIVFgtEs+0VAcrBH3Lw
/cdp+usZMq+UbHmcfdCyW8tXcPH0RAmvQleWnJGy4q+oN77MjPvEU/D4qBsJ
+y8hAWbvENXgoUGL0ztBulQMjQVRspw6VOAICjvHD593/ShOYPjEUnncQUKL
d5z/qFZ2jcNGhRQZYY9exQccx586CpLCG3h+zfSEcJmsoerSYpW857Moivuy
Lt5IERhqi0iZaqfwnzdgq/fHcMhZBT5JVXWXGJSFSc8YJ+Z79kgl8X5YAwKZ
K3va91wN8y/J6E7G17LDSv9r1SwI1zqj5ayliNi55N4DGGCcyNmfdbrP9I7O
YEoQn3qq0HEsYnHUQ8Yy3CWn17vzZfiOH1ZA52eICgMEfNwwbULbHnDQS2qW
zWLv2vXbUQcrhEFzBBQ2uzhKC9XTPicfzpOoPpJSsViI1aIBkouokFb1y6+r
U1O1vOSTJrfLXjxwMA7gqmZTdHUpcsZcer4mdxhUptdDwZCuFdau1dYpiZZu
JBZEbjascNuJk4TmKxQ5WUjTcWZZgzV6kwdtN+CyHmgLfRpzqAkO5STTgpi8
1FN1ezsZWgeB4kATqzcfV0K05gZMEJRlyemFBiZtFFbtbTLJNzMvnUzUnn1t
oMghIMznsIycOgjxfziErl0JdjKjsusPfE/rfkMTB1NwBeScKAkcfa33f7OQ
OLtqrY0HuqXyQeDxU6hKeyWIFiOVA+HsKtv+u/zfw8n1wxA0Iz6plzvCTR+w
VaZlRWr79BkIMEY6pYkW8uIqmhVWqpdD0Nl/rqTSy0g/0QZQUg8xNPhVPP4X
88IEFgllMh9auDI/1q+vVDujuISJZxCg0wSjov04yKIMnKLzOVy9PbJbB12R
zdlH8gukzIR324jlQHvmAiJJBivhWz6rZ1IOZBEaBIzbDuCm6eyWmwwgK3HG
WGHpaPK6Nx+W854/NtwijTXLUHnmiZTuwVtCL/9yE+3fgkn1wBY+zZif/sdt
//HuiSVDcl6TSgyhszGJJ/kLEhTm2Oy+5+XOF8GGnp0jAaDEUo0W3w4s9FBi
9Suv4Xar9U+FTmuhyEKWOOkMBMCha/ZvYp5pAbutl3G3ZxDzSQTpYKlKe4Us
7qbcprKw5bBy/LwLMomO/v8B2JLWmAiXLCt5yaKm0QN3PGo5E6OzDLBoWXE7
gCiz3KIpoK1tcjJUJ3ChEwMOFWLRNSz/E7jB7zV0V4FudUkbMxDIg9VQPs0g
DUzSxFbhcv2mhhO+AC7x5igsxq3xLCNoyYKuCs2sbs4bn75s2bzX5tWv1iUc
NHQZ7W68lQgfJzFExBrRDGYzFKapDoXpSNT+Ycu7tGGOTrm4GgBHHfSqy5u1
n9D26Iz7p9KzrBgoZ0u0y5ZFX7R10oqB2jIo3H4LoYKkz3Hv6FUQs7jKmVWh
XI/xU2cSx9q9LlZbm/IttRZPbR4L0f+CJS7O8TbLCo6S6LnluyPiEvMOwzdZ
EV+sDHpFDCB+xeOZwMtR27qBe5x1iDjhq8LdRw/E16h4g/IE/FGhtVq3eiRW
51ycKMW+UJBe3A6nCjvczNnAxa4QMLVGr+uLbFCW59nXZ6YZMm0rtM9xzUBC
zP/niKj5MZc8UblWkXPFOF9SWpy2coSWtCgLcnDTMCsME/Tuz1bIbLkEh2Aq
mdC+QI3FFZduOABF4pxDenvae2unfLCVKCw90v755TzpQVMc1fHHm7fegXUp
5fjIHqKLiz4Tt9+SbfyvWE2Gus3aaIvtH5z1pMlETeIXehBHz9J9RYfs2MRz
DndEed4LdkV3vGwsJSf2MDfTMI34Fy6NbTig3hIDG+wqlFK7jj14nueVA3CQ
EbPJEJwoTXhFJZ56syAxNEgNYcOXwuadHocQzdT0edmmUVUH2ZfiwESfTzzu
crs5t/PtuENHJGMeLOY8IgUhRCQ2HUdBIX2V370DM3NU91NCxTH5q8U2vNXv
GnfWrb89RIdx1m1qaSEDB7In9hdME273hcRNmAy5z0ylVN4glJkOsHtSQHtB
VI+tz54zSHzmnGv3g7YmTWK3lI884EZfo2MIuXAJQbWnPSKIAL2M/By/1geM
l7TVgmr/B7H7zO5BphGP50I75toDfRuGLOLZkbHcc4zr1YEqjlBHsmcbEpTS
JG61zJpPiuxSLTtxBshT4YHzC+rIPj48yoGTY+2YogloP068YPifCe1Nir81
IsfetzrSFKHZ71iLZCQbbKqEdvJk1KhVIvhCPMIPDzO+iswocoh2ppbfnErJ
q2L886zlQUnwKkduSfXX3VlW2i8CENBCzNdufwNhkXTL0elgc/hv+X9l5apH
t5iurzSI91eqLxb+jZJWg51oTfL/uHxYsV+2axXv6k6TixeCiy5oz1PFCVfg
wZ2jG/Mkz1+TRDtAeuio5188kyCLY0LA+EMR6zt2pomO2rboWvB9mxsiyetA
Nj0ynj28weZmZy0ckBvlNFappkwdQ9PLh5oV6ulX46ql2fV9krrgrv6/XbYv
kBxXep20W8EvojLh8CUYFqezf/Nqp0W7Pv7pa9Ywe6FLhWDJiTX61K4HyUgx
/CFf0XAK1n0FllRd7QbYzqz2NPqFwv6k+BzY7eh0wxwF9nCWlgRvQekShzfn
Rv1lFyOV1uj+iZ/Wnkp7EhCOtNU6EUAgw/CI7v+b8dMrsMoUpV+ygBMVDfiF
VOo4HEqQnaKN3Cdh423m0ZYHAMwO1OGYdGYIBRVtIQtj03ufrl8jwS2xDe3c
v4t2TswduCJ2MrX0pP1zRte1lIs8uFsH/RbLrepNXa3BhXRTnEQ82HGMROD+
bcA37uEjDvYkz3rG4/k8rPCWMJ68vHwIaA4YgYDxcCIPYfTE5sdTtAyj78Pa
tks5ofELqcOaT2MutsEHUrHJD2CaqjVQJ1eTqHbjihmu5UHrQiUgphI8BLnL
ultE1F8/H8ietKFKYXTzph//RW4ovFmh9kAm4w972SmTBJc0MGiHKve8xlcG
g2YNBzJnoLo+bSjG5OAWph+KezycdTJg1+Lp8Rj0Uo/kBlCQKrP3XnGpmLLd
ucAxJJUJRPnIVzsmIZ4RGpAe13e8PAGJxttbh670jlG4SKFpxdkY6B9LDrNO
I7QvwisET+SkbhLnoMGvf1ijGQHBSo9GuLsYrZ3ChiCp3rJsRAiM10PpxP2K
DY82F6Hsa1gBbMsiuEiN41+JlfApdNYH0407vn4jBipbf6iLG0Fhvg6xps+T
JvLe9IdV4wvdKQUtgMGSu9Zna6y4AfGLAC7M8GKS1k3zSxoBLdDahoA7foGA
uBMVGZY8qVgUciqugfgxbqKcCe0xY/YW1KbJeWNnnWbnX2wax5dXyVu0cdmx
fVmtCq0PnAkoKpCD51PWUf7j2WEG/MKz7q0cf6rrHtSqXI0JIXs+2VNmW1rM
V7synfe7lBdHYSi14fqDUXPbyQL2V08HOYAczlDfHRVSu/Rzd3lWYSwHNGco
lalZQLwUTxAq89O76h1+sM5mXQC4AEQcc83c6TAXDJaKxiXRWbZtflwrrIZI
mHGtycHy/ADMOoU4MJuigDZnZZ/jGIeRJupJZjlb70qynxEPjcbkOV5RRItV
0pK4Y4jTLzZ0Ja6dZ7Q++sT/vbfROrhJdhP5NrSIrjWPCYdgAC95JamW/gaF
9HjNC3taWl5iGzk+CybaicCa0QwpKGFn3XYUkczwcx1Pur/oMfyOq+6Grytv
O+UmtbRsG61yFzuloXVC6O6Mwk7Wy8QCXHILK98tZ1UeQRekVxmN4dNMNFRg
CYYDctiJvQ4SfXk9YAnSBpyWIhBFaF40KNzkZcVyV758Ltv/eVnD1zmbLMMy
DNXmZakmklZhJI5Ztk5vCOUE24UgFK6H2GVb53yy4TmN9M9JxHRMLdBVKNsb
EssN/PA0dcbVt6GWbBSPBToLD4SRkNWyZ+cTace4YTTCKSCGvlegojW5q+hz
Cn0BVndZRuRmQp8qZffEjA31cNy8+muydzr0uMMNV9LOcA46aMX3QAUby2jv
MQtmth7PwxghQ5oxQKzZDv1J+TG5Z3l3i3nH7g51a6TPG8sNYdyCilGJRWiu
juEzflFJlS+QQKFHiRl3BFluONxKAPg9JhzFqQtlnL7LLbJIhBAzALyS5qUk
ds9LM6wCvePBDbfitPtGb3sysVPIPPM88Xv5gdKqmZFRnD/Tnpq9NN8ApHqU
Zm4wl4WUvmArIot6MXu8oCG3/y5H9c/avCPolnqSWJYxmFaOiopkDfkzqLTh
RvKJubSIiRAsdy3+3rvno78JuuLiE+NHeET35QWuPr9tg4iMWMh2N2aGTPvw
8m2e5grwLT4rB5bYmVzdImODMBG2NO77quoKOQUN4krM1SRQWcihmo+h6VEf
eZRRrzLaQHkeXeGg5B9jDLeIuN06kpyz4e/FNwuAX9YGDGe9g+TaIncGhdFx
DqGaB6YyFAO2qHjnoplpOHf5B0ebliMtAgImNwmHnSasRpyCaauEGQDyftFL
QR3qRX926xa8T0o+CKcp5+zGpubDF/4n5jq1DTw12vZBClCW6AV79xjoGMk+
HOGZQyBL/gIyHRVkFBB4+Ak7xZiFFFLb135rTGs8yt5q4/3RLz3Y3tE6ENAl
rIpxarLMrFTJr158FpmdcyRJmh2JL0aWV2jt6LnjCHC2a3GzpXWoEvXPz6+2
TUMLEUfPc/YA7k2Q/xEiPR83D/Vn1WtApPM9bcwST02w0bJHW45Kc3JAlmx6
Sp8/npHnV2IZhVjVELVtAbCdYQIM/+YT37VEz6WHniAcRlKFyKNMINRgzK2l
5J7wgmIsBPU6pwjl4bBW5hIuk8hYx/GIMIkygHQ/fJsFtFUfEqh4SGu6KAD4
6BpS0MH1YJZRrUN3Yn2LE/gMlUxwG9cn9IdLauPqYEAvW74SdNmlsIx7vKE9
GnXbQJv45PDbVDMj7RpyYm2m4caQPihQlNoaJQY4fVk2QDLfHyBAEfIXm97R
Ihmz+NE1gUivKUFL8OjKuSn1tDQQla9qINU/C3lxzrzxLAqnb3W8cXtCmbyC
HI2MNlAOc41ArVPjpJhQVruLCqdT2Y3NYtz1k9/G3Q5PYqSXwBZl2fulrpsV
Yy0TPzJRF7TIZFKbzD2Q8wBdySlHxMky23m38rPKQZWUPyLK/6hB1RyhPJG7
osHJRQK5M2vdyqKH50g1UdaHLBdh1twvYw/lhIXqzqlc8DwDmKwo183/YuEV
W5YuZCNtxxv/3cnJk9YKcB91e0RvccjtnCs+X/pef3fvlY5AKMp0GzC5vWrX
iGNx1o6p4Qt3mRmnMkNlqemL35fjg7OfW+IXZrXL5pC6LjgeG/i4aT28iqYv
wHMc0PyfQjC46vJx2wKNH2AdvDISZA8HHkJjpItEB63dCu5Q0RJ37rlabakK
YtyK0V59eR+U9gAaT9ndtC7iBpNPRzMrwCRg+WdNfYML5vSkArIJ4Sk0FSIb
XlK/j0P63sBYoDkO3DFXDffm1+H++x5NtO99+opf1eiQx74B+EDJEgofH5z8
S9rJ+9kMO1y+MMZZl6Ppj+WhSfdz+1dzCGVM8GfxW0lC2qwQiuKm2w+Pv0C7
LIxMiIfNqvBnaM59Z2M+21slvzJnqF7cdXYNZSzUlsx8pBEOGD7rvk9BbXfW
o3VxZIDLpOEB5hX2+5ikseisYlrnlk/GhpkoUwsHLN+pL+GOoNKxh60i4pmW
GsCEiR7Sn4lkL1pSPjS+fpPITjnf54U9J4VzHtc4nMa17dnxlJvdf3jW0OHs
Y9oiNzyo4/G/U3FuYV+q+ErrZHI7rlqf+Sr0MKyJW55jZSmSQL5k3XuOzXes
0id3asTltXpuzlR2nh2mXq7bWKTDOFjI8STZfXqAMluT1fDY8Ck/NyxugZ5h
MaJ0R1aXpNto3Yrdr0Fc1xHYgitEMmXpHSUO51EyY8Gv5VPFYBl+kvCNJ13l
8U1KgfLoOTBw/PP/L3QJn+Dx5nT3CPBJagVhREPKvKvvGAZNgpQwmGqyO/xZ
Fr2l916qboZRfok/guHGzd7KfETYoxaoZHdfsU7pDjhZ/IwLPdL3X8Eebxgk
Yi4EwPJOOTmo0AHld5d9fORaTMiGg8NKrXLc3D/tzmuUjOGWMlu20fTgfF00
sF9uTrsPX5ywWiKCyQOMo9oxu3Shqv5CEveIpplvCdNr+V3K/xqkaEFhlYUz
HsAye2R4HzQCNRvGK0a4ztTieHypQ6/wJe1D0f2TC/wSUYbIp3hmGuIij7Yl
ePlBMkxtIgZ+hBjk8C3gRHlKwWhXNKPtYEAywroeCmi5ZtnzCi00ywyQYla3
wyvcv7FwK65mewcswFJpy1cJ/IpbWpC41cg+ndD3Fr0QmbRzAUjHLfCOjtUb
tSiiBSeqCtmtoe7W+0jwahYbZipRp1xAjMoY9LNnB4QyzzLMvh0Lojq6tnsh
pPyh0qj9faRgLkwQjHgrX53BGlcEuL945PvPpNiq0lZiDCTarN1u3NjjM4vo
gzfkNosbO8jnHGxTQCaEuqlM3VXCs9Ay6F92qxqcVyna0tzhdw98OPinsIgV
TS2P23uaNl6qappLNVbxw5kwedIc/66FvWdiQ7C/CyyaHVvOoAyfJN9/8h/z
VgfS/1ipfP7SkpbwoPear5MLrveieJME0QGw6E2bHVU5i/BxJ+3JT5WXIAny
HZJuP+XipGiAl3btM4qV+xIwuo8vYKUzrXxwPBvsXFOMMGqt3zKAtuy50faz
U7UAy1g64OeEn5NNlzbJ8soNKxKYubC0ONmEn8DMgGHNQBfl5Potomt+/4Qc
b/TcAOlVEXBKm1Z7xZsIOFAd/4DjfFwrc+KqCRAPfZm589fdiXdVpkt2TDmT
Xre1j+k0S6UHjxe+ymAS68aZ4QCOxcWGXBYJoZeF5bjwzfSRt97b8rVcLhVR
uVTw+XiJYbGkJn7zT5OMRM/hdxHbbCw8Scai4/mjyrM+f7/L4123phgWCSmf
qnGHuPKlvFQCP6u+pjr/vOJbtClCvzoWg9/Kw5/L5dimx79S8GYyjcAqwk5J
UccheBT4hn/L9dYpDz3+6R4AGnlnbFnSmYpxqwL6Hd38rhfoYM64DOC1iMei
BhHfcZFtiSsoW9WYcggFR+1C0AAijpzhQC3TzwXP04AyCC+P7YD3w1EJjuiJ
jbLy8Llr9KkUng+Pk0I1yGk1UbwfBvJFl8nXep0aMZORmCyY9omxmfG2ipqF
xgg8lyx0Be+GhZ1D+BSW705a6m1UO7fXVo1ADhKvWyvvqtv1mAQGgqVnVoL4
kv0u4qzghHIf1MreNdGncKxzL1SyCRh8E21ld0KFsAe+7LxworGGeQ4xsmiu
i/te8wAslSPGukoV+CN6Gm/Tc9Fruw3kQ7rFtxqMyDhhV7gZtyCnL18rGuBM
1Fup4rcrfI2mRCehCFsBVs1/RY4dOqN6fj9t6AVIkl3iyRVXMMy7KHesayVT
xAlWjzhF5HambRghg0jGB6mkQ5yt7r3SqXLNDeXZq7i4TFPhziN3QssATalf
aMJ3A0HdYUzy+NvXA357veJ+Ch7QW9c0Jd3XnpIiAS5UncTc4nzI+EBHSZSt
NKpC6YXc/tpMMyGJuS4BkH4BKOj2WbcvxQUY8nhnDysrpaHB5f+G2mksk/V4
NFdaMviGYRhMCC6O6dlrpT2ejqKRLA6PLkR4jHypPMn/BTBe2Cr/eZBVDy6n
xk1AW6vtRAjo9P7r+NbNIsQ6Bwq4ktBO0Ncati2xLs5bgRWU6hMtYuYv3892
eTbGC3vE2VCvzMMZKd9J6lOFPJkS0ioaTm4cDwrdF2ZKhcTQZRXCLrFASL6s
ih8gEo/vSIiP/sk5vJmicjP8yhse6Ibx4MuySqVHx6qmoRMROLB7UahPml4J
oCTTA4tdbJ8yFsPzLsUPpaSEQg559fvTAxtIstZKpsb0SU1uhXSakUldX5kY
3+ctrRCMLRfEqNgm97QQuSBkKGSUO/OXcdy0QuyLRen0H9Xv5A5D5uP06DP4
irdckGN5xi7vCT47px88vuQOo3GHnjES2hu+OwyQBZtDywEkUkY3A+nuztuQ
IkkawBzbpZvY7Vsfih6bvohfjLUhwFfSqAFodtQ79iIF/WlqN4rL2PkTdx8Q
bZCGC3RilwdunCQbXfdrf7MQlTDWFBx6HCLWEOppSTCbU3T33FkDBrE/bi1Q
C83KK8F8huAvWcf2njLKT9FoiBacgRK6deL8qb3LVdSnQ8tv2zXRlsIMQnZu
N/OQVVdtDwC/AmKBl2F2ipLwKzpWM7Odrj7KrR2hxgoyJePVuokgfmLsY/E/
MmvRKDp9+EUj0VsoVC85Sxfz5FsdyusZNn2EOKi6q7b3USBe26WFuDnElVVY
PSJ9qar2PyXpp3mdMc7iP+2hgpegyu3a7K+IgD3oKy3fKH609LwXNHAydB9y
RK/Mz8txEF6UW6tTx87BtG0RwAtV9/ENoiyXt13pChEpZTRqC1nmnmnZJOCy
LqjNaw7TqwzwPa6q/bJ5pgEbQCm92KVR37urY0VsFSXfLqeYlaFSuhHTZpnq
PfrG7c2I50oAw0pX0XVfd5YHfMMa8JTx1G1uKFrRlnGUNWEq5juRd4uee8uy
Zy5ye2zRRJpEjNALV+lUBVlhQraQIhIexzM79jzF6WdfrTxhicq3vhhpl96G
z9jgh3suSWvIEu632vd5nOciSHyMX7RdQ/8F1WL+zpajayogVLG7PnGg8oNx
klJZHDooOYNIJFtccom+8SsN13891YfmvU1goQNb7Q08EETSHBaUxfP+sv2K
rX/pcsW1uPuyJjscUIZIxrjY3HNiDd6tuRO3uWv+VddYUA1zjR67Oh886MsF
Ixed1VO/hRaEi/Ja1SBysyfHTwq8J+03eQ/Gwsk+7iRpM74CAiM4UeOBICKP
NJangjZIuXuzsYm0mJPp/vsckrxJzj/NZR6dI4cpdX/0ZH5/jtbH6/+H7fBq
a+pZhMdF6v8BFB/SybQstmIPujN5ChVwkxlVqE4D2eUWvXrZY50W7Ptelrep
FtYjg6sMr3KDYqann2NJMh+kqyY6jM/AZq21Zf2czUrPo5bZHJEbYt8R/ni1
nWg1E4JJiNSZWiORkidUv+id1VvT0l6mKQtr6uL8Zhu4VY7KJUJz96XGc5YF
SZGPluGEdQPwG7ur4gpX1bvC3nDUFqHUxvGS6XyGFC1LQHqJvHcvGcjYdSij
gmAjkADxLIivQdu0RI3C1os3t7ulFGauERK4FzV/ADxv7p/c7MtD7We6EYp2
lhrEMb6B7cCFdJ891/N0hKgLJNfijbMcnStua1DtK3TGs6EHQiPZEk+ycM9l
0Fo9Q8xVxvS+gnTW9GLttH14iQ4hPWjuPQ8V6L+lWRDMf4Q1DMOw9CJt0Zly
kvy0vYWI64i5shWGn0JAhfIVzX4HiUkN9PQpl2ubYTFes4liblGgjeO2kZPw
Itz3duUAx4vo8vzRa0//qQobXpMFRB4hE4G5K2B6AWr2l6s90bEaZu3ockmL
Y0wO7l5qtbPm9ZhbGS/uSJM8KYO0LIZH6uKZMjZm2iwAmuyB+Te6KgFPfWHQ
tmuuIQz7c5J7zenvKCg/R7nKKu7zR94QZgu0sJDmze0nUeZ8dozvKx5mrVkF
20Zx+a8iyh102hLBVpE48LHpguWhN+bVn4dQgiHcC+M97+HfNiUOVWLwOdSB
01pyjTIHGg8Sw/8UW8rIckT5gCVUhR5PYiLeyz4Emw6dd6Jlquy0op9r+4en
OYTQiNfJP5rC0pFN0z92/9tARztsOGDTx89Qs6bRlFz0sxmCY7w1zYe6XIVB
JBeQPaogd5TCDlKtIYufKYBEJKm6demJEYg6NZ+Xn2stdU0WVBoi6/oCkpWT
+5AvKfpoIM8+XXtjJmocZFtegtou0M1YUUk2JyVxf3jUhe5cV8BRC3oynxsK
sZCLMyFxkMOLJFgzqg1CAUocp2Rw8Q68zhIaxAjJBqA6jYkeEYFKPE/+dcrP
YnX6vVcXfjo0LuakmuobTnRTwfGE8ahj/uIQnetPLQQ3IjIX+n2Rda09Hk32
49CiiKUpAS8NOg1RyS1hDQ+Ciao7BatV1QFA1rOBWiTHfDRm0EE3yvVRCXbg
i/EoiSGrU+DbQUsSxwmkw10JW86z6We08iRYuuV7+SxOHWr3C8RReK30htnW
AZ0UsxCvQlJycEz61aWvsilEV97RKllp9UF7MkylyBY+sGm4BBaAIddYUpME
9/RXEF44WEM6EaWfEkRlKGMrWt2mlk6fIhsXSH21W74o05YW9Aqxqmcx9iR8
9xfUDmlf0BjDucdWKAk4cF//K7LXZfbRHg3/99K2V9rsAHev5Feu8KJ7xacV
olYDF4DO9z1epklqE9tiUyhPr2jw8NQ7ONhqYmvYlwMxb12yPiOjFzK1IqlF
53YlzKs2sFwt/Xrj8tDQygSMz9+CgFkzRvC34VM7r1FjkiQNqjQm2b0ku1F8
ibG7/eAEXZ3D6kPweN+mMW6s14RytlUi/J0OiQGinYwvvhT2+SQPjtMghpG2
GvRCI2q8JbTp7TFvppqx3she31ynFInWoTkqx3/ZaJ3IW4sTbKBgXNmngg8a
0QMpZ6WniPEX9I8wHVnfv5PqrB9uiQn8ABf+F6xt7IixFXDXH+k1ioV7mOXc
gckeyQlbkLKrJJqzKcP3NUQOJxxtdRkF1XTBxdnd+4Dg1IP4zKwUdpTVUnxS
D2mCTlkyLnfI8f4KW/ZSk8uFsFLyv/QuAryFanbkDM3+bXqEFLun5c7l+2Rg
0X+T2m+sE04pMPFTzaeO6gLpaD3Lt4GcdcEL7fnUiA35iqalU6PxUD2Fiw6e
gik6TY+6vG4L9ef13YuFsM2/E7/izXnxdMd6JHwFImf6QxxMC7akbB+ZKJ3k
yJZD+SWYyz01RwNmT8VE8fdDDPzB7Uo0uzoIS7ddyMgfAPvYMOX8uZIkVoOo
xD0cX33p/bGhphZ95HkXGUVDnpCbxBUotAo8Z+V0Ln9c/yfcNLwl/LCkxJ7p
mRsK8Ly51cg/F22FnwZ2CyJhf98FhnDRc69yXkRiSYLjlKQUdK7XJoi6ORCU
fVFXusda/xUUX8edep33k6nB9leJUBTnTUzhAsXLlFUPJmoV8kOX0L2nQo4i
Im+j9+oqClrgdk7QucRnNJ44Lry0gdflvss4PriBwyDAMlzol/cMRnbKnn+v
tWpAq4SiEcN0/ubTgxe/lLtw1+/YIdfmqcXnfOPlo3qdl3inTGSBj7BjRsvL
uBte6oM/wbfAmUS8D1AlV6bYRcJoNBKOejT29P5qeKeZol7ui1XTm7mPDzuP
muXafRqiQWis/Yj4kANTKTxGrMENmZahrtnloWzySfpfGokYCLQemhKvweJo
oVEtgAg80diU6bHOSr/lQDUsDUiHjfir+HBZHCqmVgl8F1eWdqFxPFDWx/Qh
kne7RgX5Ho/9BcM+L+hTq0a/JCRJQTcHxcQVRZlPGkmGC0hG2bhHBfKsHEf2
mptGN9McX0Z7hQJBz/GUSYQTAZpXhIdlNEB3uF9Mag1ItYDyGZ3CtcysOPCF
UEpq6wt1wMHipK/MWWzkFQmQcW+E/Xx0ST+1UsUx89utuUbAv8TFKHOk2m1L
LbgWX6CQxAME1nQevhWlvD0QK9xmsDzmVjzpUwvd98i/VcJPZoBii6VznIZW
q89HCmq4hbo+82YO4jtOyvO1UcUdiVA12w29UUHukDQOajicceiALSrQBMFp
Xu2Fw8gqz2Lpw0SR8IUctvgM2FNvPPFmW8UR48GjDvw79Mg0KYtEcJwvVnpF
wvFIVGFxgmC0NaCT72YchLScs4NO107CzTqbaZFAp20bRTES0hwZdzYCagDL
32np0rk/boOyH7e7c07C9haC/RL3GTS4208KklEr2hgIEuTUQz6HGnH1Fh+A
r1aBk4dlFgR/0vTu3fMqfHPn7SW6N1jfCOVTaq+nRv8u+i9aolIPBZs1p1zH
CCgjyLue3WhwzOjBcU6KTuJ401MPurnqTQ4Ct4fqZiXXa9jrJxIgL4MEopak
eeh+bZt8B6hKbaXCyFOMXfOxzGDYm+sXkKMGDf2mz3B7JVhjgpOHf/RQi07x
Oy4eiWDoGiw0wXmnZY2YbiFaxpa0grsDppeLu/Cr4dnnVkOfaxW3/T8vUX+b
M9igwhVXjNzW3KO+Z8J6BVSt+SBpmiDV+r2okvOiY38nqvHK+sIRwc3KwMKv
du2m3zunOtsjVyY55mGDStbM+s1rO+7Gb1+CwhvGfxnhbjKtrMtscKN1dC6f
yrJIzH2NNWL1Cs/yu1+VN77JqTGwZhW9rbC1gEjjqU+AJaGxqoX+hkM5klCF
eG8t+zrEIw/eYO0juQ3h+hk+m67l8WmRTb2rUbgu4OQAHLaigfO4WkBTC+PM
QyUc254nqTix6bcCA/YI+O89OF4bAaHQVEyOzZFVmW4n7YjSMwBcAJhA927b
QSPf2ZBI7Zksl7+0POy+lzLT4JMS86RDQyPOF/bjUHbIK+44roFhFL+Irrlm
LGkSRNaujleqIpIxWcI4EQWzVCzeOzLmqZD04nUygrntcAD+Fq0SAOGeKMXG
vcnTtgMCqYBqaX8Db+BhZCpsRDwedjCxGJSHsH3FgDA4DuD36XgqeXheOL0X
8iwB3Jc0Y51dGfY9xPG0n3AqWr/z7imtP8Murclfju1LVV1cqPbNrz6cQCcv
+6OFDBAYeswoEqyI3mRTiAP86hzAMLxhVxnfHTeZxeGAxF5sXX7YRBwg1fI9
cQRKYEGtqMa4SLRoYbTxF/rP5QjUM4cSuFikW/VsJztfk/npI7gmmlk+1naO
+7D3I7OW/4X4qxiWxdDS/a+8TjajurPpCamkOO+E2dUmEVrvD4PNZtIRtWkM
kcIPPHEqFcCMrVVSgGnEkuJv4AK1PjATmlXVGfRHn7ttqdh9nSNIM1TbnppC
TNHdDP0AX/iBKx+MoibhZRa8ST+DnxuY9CfklirLzmJP4AsKJE4ntCnBqjU6
VT0nY/vcD2YNxH4Uby4YADJ6s2v7mIjU5P8/hvsTITfeIh4FsoaRNCQ/dU4D
gkVJMBJGcZWBshRmi3whOBiScggFNSMyEgPEbqpoRs0qrhvn4Ievhcte5Q7j
ey5xkeLMX7aNH48XnO1KbcVEWQasAJ0eJ8MbS5Cyz8QZRO+vIJhfYwPYYtsd
A7wGeQgS79rfXcEszmgQFTXk44FcuPtTY4TlzF4P0iL/qh8/zdGu8PjRV+mI
JDO0i+wr4pGsqScxf5z/a6AubN7aer8xgtkH5FuXEw2IzrBNTRmAmFZtvAJA
LzwScQm/Rlf6j8y/ezu7M3oWj0BkuCCaJ4eG47j7AEzZphhc/L6kWLo9FiPq
TOmgrRIX1ZWtJOHykOXI2qpPO+BFK/eTcmq2sBBcXKR0iJQzJOqOo5NqD0Jw
Pvulhdhxv7CwfNs6OCsfS5AznifezdYje+WcHBfA39pzkL4PUv00sy5jkuLL
sHr09TTX6BX/Rq/Zm9yQHWtl9KFXkB5htbjsSYL/ABINxIiT3ZuCSyDcpDfN
+1fprHYr0rpvigUfZ/wmRxKwA2svN46GpKopgDmUqtCJLkYwXPmgup1CUnB5
WOLf/dmvvqdaH7190V2sRn+pCC3BijKi42wk0fCsbumWM0HjhgyDN/IwcjDH
8McqSK4CpYpmxGQ4e3hQ+MuTJX/K+4/Cz1WobPxPaFjwB61QwaneG/uWypSO
mwurIsTwEwW1AxFinnRjsmaZjaIXzuaeb0Fo/kihUGn2QQCiWMsvZoOlFzgD
Pu0GLfF+tDXLdinx6IckPL2kZ/venZ0z82Ntgjhfs3aSD9ZgK2fHkv0cfhJ/
z4Dv2JxHmsUD+avGfxzpxlvVP+7Sm7ekHaDgRQI8oP8uIgZPUJR8wWvnk6f4
U2jooq2I+DETN72EzzlMtMV1uxBC2K9Vz33Rg6j3Zn3v3gCQR2rjf2w7vf5O
ojAd9oNHOOGJ3HCiRwnqNfRO1A51vKS+XgrOgQuDcgrJxBuWp/4E55jHCH29
8JUAtT8Or88T+JHO2w6QJABJXKLxYCV/BqO2DJ5xemUNzPYsqYcLzWqySOVj
lq/CMZV7lf50/ME4So/X2NbjEg8exIokKQqb9B+qE5Fvzn6X8pFdTHptHWQW
j9f/l88alYZ8z8Gws+m9anTm00DukVRUz4od2VmjBseJ7OHJyPv6fZdVvXgk
zldZ0m/VU++1DrXNTPNXDR9pNSZgAfjE0ODUqAPX5L+2Ub0E232sVMJCCrqU
opceIOqPCYDyFZR4s3aoSBe/pcGVmeYsX05yIL2pJtd18MvqF4ASYWDRf0Eb
ydnup25UAsNPBBtaAU/xt28xCB28Tq8qlBV1fuRWb7T38Ex1OWMobgeIruY0
Q5NferoRoO+obM3CGV7XkE9582e99J8rBPOjnkAePWuZtMkW/JUQXEXucyIr
FaMa79z2xM/t0tbfbbSFmcq1Hc9yywwEzVT0oC/HqzO535cS6lwVFkicAf7j
FVzS352ag5zbmxPwtoXo95MjYGr29okb6BQnNkjSSYwAFfX1qRAcKP44qTWl
9kVK8SMAVO3kUAoCSO6qHof90pFyZXgCmdNT1fZGexdRzfTM8Zs2gv6b+PGF
f0akh+XCwqfiEctjkIsa7+Opan/fPqvhZe51XLI17PV6UyUGiyIY+Fefr0qL
Iy1AC4/GxHneQb9XMUx4dtV41Vtiz1ytdgBg0l7Q5m10F3ShbDBiPXusdC1Q
b1hC7Ka604M0K9EILNU/TiDu6AuNm9WZKE1vD6ynZ4dnLNn5HtN66Tzj4iA0
qZkn5Xz5+15+3VIIVR21ND4or0QFlOqHw3cnqPzX1mvF0z88Vud5XDNF/ify
S1M37dnINezWMLwZwQDoPuj8VZmhzXYVmgTlUJ3KUpOcHtXGfK4AMaCUtBds
OHjAc2anJicykNFdsAcZbCpFCvy5E000bXns43A8GneNxf8B1K97SuwkoVU5
IpLdNF6aOm0OnRvF+WEMJ40MOfX4gsQcLIUEk/3gfddTF9KLF+5DxL2Pj4/V
bQycvEfuQ6VnbXJvPm/gLZTBeD6dGkxgO7AQwmT0k8C0Z37vwMtWoUGl0xRZ
M+03+vpnyffKFJ6ju3WZgNnuXe1LvWivGWN90vtBZd56I5j2ZlPf4zHXaTZY
zA8ZZdDwo9yLlxJM4McvSLoPrGbtGzplAZ/+usN3URA8I0xm8FyNyAbxk2Xi
WJWtprUiJO1iRENWyO7iABjEW9JXLTiHE+heYe0ZLz+IAU+Ko+2Eo6+a0hRL
taussKNCfEz6bG+dRQBZH5hdjc8xbCln0wF0J+dJnHVUDnD2SVkXgxo/887Y
+Qw0GXIBjSkNgpI+Ejbhe9/3UQc4wfLEXG4plcRGgjS8imgDEi9IYYMl7A3G
et7dXxOEV5krmnIABWgqqJA5pTxNa4GcHZ79amFg4wfltteFpjH4SSIhQDcJ
t9CH3Wohl93QGLUzd9jgV6WKmyHqq2ATeK4fn227py9bJ54y6/MFVkUV8mDt
UVrjPCghQ8QMcZuNAyR4CrKYdU2+BQHO/2NemYedFwC1cZ0mdeOW/0mTX1ZZ
sxhT+Q2w99nV16JlPnKTB8pf/zKJy2T7InhptFuhzY8f6JJgFrgxs7kNgShT
XW+cFR9jpJB2c2+1Lp1WxfMicjfgSr0QjcjyXwioYAcAlia/wmAGSZTWDHbZ
BoTOFROlFngBzVpLAWke0giOhAtXPWpPFgaRJ6JH9sUtaGdejB7MCAONDqRF
PDbeRG9B11iXxBxRqIRIx4uy7soLcA3l1q4ajOrLGpn34HJLuIaszoV5N6Jy
ZbGhw6kkNmzOwa8nT/1xof04AgCkeRWHCFzfUtaS1v2nBgZ44pK13Pk3fNs4
v008nRtG9UQ98gVCB5oPH8lhaNxC4slY5hh2H3geA4g/rcWcOcMqdeLqA0Pa
8HCr0OhbZxfruYnNUbUyhbchhph1YDBK7vNsxo3IzCqo3gmgCovdUjvGTENg
RkvyJhkWF8aHT/8M4sX8nArpxvDQAohx0i7cNKH6WI4belQg3AWXQs7yhmn0
rJLOHWY4pgasjS10pRHE73npyDnb2U0lOD0Gy7bHg2tmunH5gpZILNie4HJu
4GVkWE5x/ZY/Xt4R4eTmgm3D4pGR479tiI0TUPLvmxH2XPPbbcJ0iFLWIHbV
IpejqRAnNuDVTtSVtZI2JgDF2k+hDiD9Du9DB5COi/E3KrBGLhb2WSbsVajU
tzkPcGEMKPa89cthV6z8hOxzYvMaRFKak3xNBpy3pfqd3XE/Re0ZJ3Y4qp/b
KkRN6FdbJX4TMefiJXY/l+DlW4TgAyDg4nv7M25pvo36kHLs/LbTBcjhMODw
cB30dwUDjgbAhifPOXLBH8FNf8bnfY1KMOraKX7byjBlAION0RRW0qn4An2N
Y9mcsbhPo8XkRoO/JlwSkhhdPazcrPxs0AOFm6sS7AbP/uIb3OtwNQSymsfG
AYg0nKD+xiarM+1cHSjul9pI67YYJqxG3SFNkftXScMFwyye7BhnPIVtChc4
a3QTbMCwVgzyspb4Dm3QoKMzSI3x6O4DLjfm7rZXY2sFNGTxtPhGVw0k1iEJ
cm4MOg9ZOxumaMorkKOBDIX5+1dgj9uATbhAseV7+EuZudDtmUPz+tfj7Fhk
ovQ0Q1XK01j4A3YtdNjjBOKouODtqg8lG3gakBtoCyG95EUzWCsIDiifENS4
rsmwTqJgWAdNJXK/8hf2B8bovJT8UymIPzyqtJRKJQAm0OlS43F1Pq5rLdAT
biVbSZcIgagVUPz94ScaTUA9juBvKDyE1UVxe4OAEzK2cGVj+dHNsUWiQp6c
nF3Ht0nZkSShHDVktCJYI4gfE1kyPLUbXRBrFt4A+ZOED3WV1sX6o3+odLKX
jUYTe6//xaBCi8eWhWH0KGnxiH3Y+lawGiLy9E/aUwHGoipS1XTns95ltas3
c1bkpC7mh9YrdjMcenXyH2rS+GkMGe1UQBgBFvEkM1q71fVA57K0DCk+YyKp
7gqNtY4cNbS6OpRXwxYBh5b0rQkzIx+/PxvQTSqqIqGOKd4boJZkB6VyjrS5
AIPgywLr0A101KJdp2m3sOXCd0AOF2A5l09txykjlrUNQBW5xuQnDYb+Wfg1
EMBhZ9MzH8SZGyy7AbXnzhaVEnpezskLNWuszGRUyYduyLkwyvE5dzWsMtr/
l99pxJMiC84qXndoJ7qSX+3PozZIpPOTaoY9yl34p1JEQwyoMsF+nhS/jTEl
7ZJkCFm/4wZS6kM1mjA5J8dJtcIklVfSVrP443rPd+5NdD67CENqOON95L0k
LcuRbgKw9M9rcRUcnN81LnkFmndfxa8ye+tmT5Byc7LckuKPVJ4xaKoeCwF5
SKP/s0vh0SGG6S0C1zue2qhs1pJojlbC3Tv3lBRMUNs4gOa/zcIt3urMh30N
QEdeSuiyMKOoZt5LhulMscad4AhgZ52+6uBKTXifdZ0SebUdPS1WMQap37lA
TP/DKHe1NlyTS0E9vQKs3fK9dzCrraML4N1zEi+wP+thniSIp9VO9Xidr0Ad
96O9Z6jmwuq7bcXf+9gZIeGxGH4iAcuKUUtg7Tbo6UJEyV3uaYs1nFLm1mSK
VoUBeAYdln4WF/g+RHyh1M38Rlgv4qJViDP7r81tFh8GR0wMKPrLZX1QOI9Z
dBCt8CRS6ys+IN+nDyDeJNUfb/z6AgLwTZUI9pyheagtN1yMXBT2PFWsinM2
+Re6Cgb6ke5+myllZC9Vj1fiYdmzhHxeM/KD4WZVGYGIJckFk6jPR1byayZu
TlI4JFSN3GOze2O9VkGfSszPmIOn0lDQNwIxCaKY8e4cXN/Gpb+aouJiKmG+
HHPIUSytjX01QRvckVAmEW3+4W70GZ6HfLW4xVCmaqgjAhZvnMri2HzDoc7C
Dpt6GNCHC5XAF6lcyk5XtX/ghhOGgHMOjuUv7yzQ3dbBpdIuyrfn1mn3K0/O
w86AjlWesueGud1onFyelEORaPKDRXS+MgUzZ/cvDAKwYZcpBIoXFVyjwh+H
47hYZJd/sw1xa4yRBgf+uXwqFjAOrI9ScQ5dmHkt9xLk+jMtcgRnIfykpV9d
RHUgjhlDEKPmQdhf4u9ss2IFoNLXh7VXinISVPf0pDuuV3IK5pLXta2JBia6
t7sp7gjmQBUANw7J0P5rvJwjHPcv7gZn8TtmZ5TRFP14bcAhN7OXiE+dZrDY
aq6kxsDj8FNBg3PKHGDa7sh8e76cZe8gsfWJAMWB+vBcdOOwosUINx+tRhhC
qQIL8DxBuxdJIlH7au5caKukDKygTrFKpeOO1dMHGnmgS2aWb2Q/TqTJFnoJ
28UlMcPNlEgHhraXTnqytcqZL/DrVWgT2N39njHaBzaA1k2YQBpBKJGKkl/f
slMhlNfxfQ1+5hNfQOjEmFtD3JjOVQ+1NllznE0O/uwdhUo0UJeln5w50W7b
G+eJWWwGIZTgW5IeGmYN68t56eYSAq9or8mQ4AVqKTx5b6gMfHm1tbpepCL2
gDGufxg2mQ6S2efMXVHwUYPn8HNa6tYp4rg0oZ+bHa39dPZDeOD9UxkSZEw/
pYX44yOwlxcq1t7loR2lZ/woRM5B7lVTXTWhKwkoSKkQSmncdJOUB0IwvMAR
kKv0L5On/U46e4ouITnieYdqjYfa8tEF2YnHg2jH3Ge8Lq6ThTdVAKSdCXjr
JpX4JPobDX9iqkXSEpPY98s/PEUdrvq1LEXwX219W8emzf81YC4CMKcGt3aR
SWxn1LddYoxa0WQBVOmkyfTcYmWJLgUoGPz5h404U8kvSW2AtSXWc8TwdWvN
HSxpgW0v/a0sRv1ZLzfge8hi9JTdZR8Ig8i7p9VwvLVst0HYKc1uiKuc9lUF
XycVkwJEAW7F80FT1zm109FllMu+5kKW5CS+NI0441lYwKlbVvYleOpP76vM
RiDMvwA9EAQqnhs3e63pzoQW2D0H7hzadJst+vliP4/ZQCJVZr+EAeL5nmCJ
APz+z0DqI4Uam+cR99uQIrnvRocprCXlBvcg2DUKoeMpRwOYhCeDWHsyhxhI
2A6FxtfX09hjhFkf1NbweaN9v6fiWbeWBh1Mwd0AXFMQbu6Eoy9KO1LGDRJr
DJZOqelmIp44ZeUfZKyMXe9yd3321zK8mgjpYQtqAcuV3yENmXAiQtKKDOPh
rLRdq6k+Pg1b1gVCx6PIzfvDEE9o391lUkz/Y2qRQ9ZeI+PEQHnuos+S1UGn
bfVEbZ4X3LSsL0fr0hNcsCA8s1gjiY9WKwycE4dmjI8BUALt0utrRMziG6rz
Mfhwifldws8TD9PS6aOUgGD52R7+qoGHBtZnKOqkajvgbzpXkR/lq8/ovwh6
X9Tg/XrRAykjVqi+uHQS320WJbSAB/ONA2FEJgML6fpPEk1IFuXnLS7Kfnik
kzYwFLrOUH6eClefevsURED3lUiWU9MPn8G/XIKMYeJTW2F6KJbeK2j433OT
wsOxSAlaEt59aXzCBSWOK8QGQVuIJmZIzoqtjAhIYleoUVJelb1t+gjU8Cdj
V0a0/C7jwJlsVhSIpm3dQ9MRKTIW2xrKtK6fIwzNP7zfyXQ0yakgMRW8psiT
gflmjtIqL2RDAat1AX5JJdTrNFUm+XKCJI21RWWPs0ciLTnqT+kwhKrgYHHr
ASY7WmpjiqkhL/XSRhETj3mwfHsSs4Ig3CMoM5dyaSrQfEEIdup07kVj5xMy
1b8NentekoxEU1/hNYaR5iDU36j+5/xWMvKdAG4m88zW7p+iuuiS6KLOgKff
eRv/MZ/waraySSVIlXREJFIzJq0Lap0Z/+C3/pA0i1umhan+Nu0CBYhX5PAi
cTmOBcUw1eAHodsBHkYxX0QI/gO+2CZSWgNRWaWt920DgKet7ZvFTcNpbndK
USjePfAFN02l93NMD+mP9e7FHizc6+Vli1D1LfAlcj7kRvJfjjBLhjynuDs6
/JiOJGAY+RpT66q7E0q/MZM//a1agsyGIqU3wXokRBRqnOnKTAvlEiWn2dU1
MDqjroIXuj8vf5VE8UTSAc04xQeARw/PuX+0hHGAdr4GaerstTQXvd0NdZBA
7NYXM9+QxjQ0YEy1xhObbW1TCk34o8z89+8dLUwbDaYK8+zpibcB69KOWHZO
9N46kCAIvB0J49Z/oglncEGfZyTccn103ICo4ouFXkYlQ5PLULk/r+BkOdyI
HtQnfPMInDlxK62mppw9wEtAiGBr77hKbrv9P4cUGcBLctRW38BqhWjWCLPx
PZMaTvW1684jVmtmyBQt+pt6ylY+kYEvWf1++SPUEF96ZaNljIytQStHGeen
0S9IgE7ZeFZYXEoBvd6Fc9jZiczaQqfjPNpRvUbwLU39TUnnZXWdxUmM0GXa
K7KrCke9GdHCL1Z1hnK3FyOoFVXK7HFUMcrSbBHZ01FzwY+gSjke2esgsTSA
XE1L6vVTOhtwsCftAzhRnLdr05fRQNrDQT3YaXMp7vV7Ae5l+6AMPRjJ6/sp
cdfOl/TeazwofwJIk5AiyAKrlkXRgkD1V97eIrPaGcezVC0vgZHipAOK4gX8
DjtngOIgbuH5XU8w7cgXtm3/CKchcaMXLlGBq7FiRt8SpTDcIKHWXL4J6Zid
3ByrHml5Wnqfl1i6VNpIAA0YxE0QgIlG6opRL7i0L1E1cn8jT3X/LizyyrhV
5KracMQPG6hQtkQfEfR9tdgvJ+r58X7WmUkMQ5nMZAfqNWvgveLS5GSZIK/U
E1WyoVJ553+9ccXcVJdiDI/vR4WFMUpu5/0QexYAAd2zkU8SXUFvVNbJwC3M
0Kezp1erRzumiH1p269+V9c3R4j8mli62oOCkS9KjUzYm3B7V7yByM1pDdd4
9AiAe01vfILHL2OCAkNFLPOPzTFARb+WY5voLbVmTC+f3enhpZr0dyVhCj/U
+dGXeuEUl3bQkKKo6MYFxeSZOgzPm6pf6PddaSgkbd1mcqqARNQDTKF1gL9F
WAfZlCHcu+sFRqu0jHTZK1cflOSjxyTj9OoFVH5W/3+kD/sEPSAK7srBoT1C
1vL5iegmMZgbJuLc/liqANW7k5SlE5pnMiV3AzmlxPWJOJLLJCq0oDNvsDMa
nh8+Z7cPhM74lGnJJZwya4bY4DpJvmO45loARvGnE7EhocJNUGatf59uo4PY
tY4NRLX/BFGa2bhRTYiyUgWsZZ5uPgaLtpWqOROFpc0nfsAdjm3R6r6aaOGU
AUjyJ3RlkPvunKJskFyOQKzQO40GlhySVHx7UhnZiG/BZkD+tiRUWzYLFjtM
8KwlYZ2RjKCMy3sfuWaIw7CBmZgqfR8zH6Q+RYYnFYLJA4Sy5V4ozBc65JAR
y4WOtjaqXXti8EoY3h7g4xP+grnpc2+nHSRAKbxIuGXlNOVYHdO2x6PhbHiU
Fk2np4UGTNkh9Pr9IOgBZKuwNmDUBx9pnYonniH4UFnrSSq8pewJaPtGAadT
aKE2YAvNjAMwjTP0vOseEIB+3XA8w77dWw0AmehTQCmUsTAKU/g5+Bwv6Ls/
WIROb80XjjYVdZNJwUGFkxVnTmR3scLGjkdOvptj5XcioqEFxp9t/qmtrGuf
G1icKpi5r8TxFGTgvn8tZWdjc1/xT0cs4Ko2gqYs+wwMVfk2lERL7sE2jOyW
/nVjFjxxORezq6MTDO8FaC8U7VG/1g79Vl2F0imjk2m8XBLV7p7afIFow78/
bk/gFLAjuNx1xwDiBfPGiPtYocHj69mnKYYF4NDEWY9o95WKwJleN4+E1hr7
tcC8My2I4r/oFlqzNiCWIOJb2wsfeJ6Se/MkKoa7bc0dy4JzaaWb+YTaLrj3
KWuWTwjKad7jfYF6gt62z6i8xRQWbWo0Y2l3bO7mPP6VdpSX12h92g9O0DBo
amrYFPJbpAHKSGXplVlQO5v+P+2XEBgVoC/4kW5Cp04IQOnjMUnkBW+Y1+ar
bfEHGGZPrs4MdgfY3AymkvXuqDqdCW6JDO7YRw6i7LHmO4gBpusbV7v7E7F7
Fe79w8g6C9iCCnlpbY1zmtAYS6Os6+7dL432vC20XSU9qvYZKadLqQSWMZ14
TASCybzylEJX3QCfeF0TYz8PGc7KHpqNVTCw2P0RsxTmexpUnLhiCoOZJOur
eXXynjkGYYN65n2+3wrDueYbqmfpAegzGn0XJ109WUhQz1Ztg79LKDR4/4S3
dUTO8yLzOSvy4taEFRvMKvHDYQt3No7xFcrwXtPeTwtp9tLhAEYBa45vjgCz
FgKGK5b51ITPcXhHXa2ZwqJ43q/2chqf8lpJ42cY43fNzKkdeoXFVYjk9RH5
S4mheD/NKsasCIfpQn9kVO5OWGL2VYNsMIWOcwuEPJHNGV5RDlfPPCDmKtJ7
qqPEnrv0w7PrTakY4dbc3i8jP8x0GRf/Ecp/8PkWP4gG7RYlJIFIF6nm2a33
Yc59QvHcRcVh7xuo5sj6LZ3X6ct0u5onJyZrBiqt8wwOYxjy5YE+wsdHEgwV
EzLv9nmkLck8p87z325RiUQZSVqEEP32l2pdmeh2v0wfvCPw9mNfCstnYoel
UMyb2eja+zUNvV0oRycVPsLY8Suj3yMPTZauPK3/45TmrTE073hqAdEUoDDL
NyKw4bQYVGMZ4ny4gDTgc98u6g1JaC3Zjqri1f9/Qk/WYBqpsZmaahMb6dgh
hNhxbpfFBx4i5drlzLU7GqWpSzOi5QjoWrCHvuihA3HyOo8oaNm/A6vs1iFd
Tr5fNl2LwZ94CpbTfDIjJX48D43w3wqdyPtYUtqkqKhPOqV/nBoWVDhDipTm
Hysl31J22rCfrMRcREiw933cexVhR9DrAwTLCFsyO4MEjbfVLe1IfHp9avz7
8Vzj7IyTDhO8KSIowOPBv0E1XIcUEIWE3sg/VrgTPH3cwcIKnMmgrzfnKVYw
bKHfFctOP3W4NmjVWgSIifZp+tEV3T9EmHFb1IUPZpbkrFJ8H1XPLSp2mIjC
IUeTQHpFTnLPL8vWQ+FYmyOHe7brwxxzCcoRSueX/mKdKM3wXxdfTsHGJK9W
OBrw4E+F/5sZ0LqTdm+XzH7ZfvlHhHgAuvzPzH55XfFfw5MQBr+Y6lA7apGa
kuG135/3mSNQO7RxIZpBj1nu4QPz3i1sCQvqj/0eg1e+3QmMDSq3RRQhqhgX
wKRBE9kNBnQw5mD4v9lKf/E1GVLJqoUQC44/cKhetk9PZw8SeDJHsyEB5hwe
OgcFnJTSvDKS3Y/6pc+G52F/C+NxZeqTC4AqEy5kYFE4ouRn4NZUAO+S2Q5E
A6sMQ+2ttbW9tA88BBTKy19Ek2ovE9a0ASXsHux6bqZDHs3aoq67EipqKMCg
dSyPAI1RsicNtH34MKjUm2EFFqbLGRB2eW0a714SSjiZwl4SjRhGGFE79krz
XyJr8dfBTFLaeePXuzUoo9cZ1I4oFU+58SM0T8AtL/pF1qi8ZcWv6/lzv7bU
RsOVJej2v80k7hEupW0gOkz4rWW2QCNVPFJ6yfNYz2FMjdH/7GWKYUfkoBPA
hvR+AdsXEbDFFPiTDOQ7dmpmMdqKOgdBg83PFfWlVFAsojPqYyZs2AUaTGC4
XzARMrGREfgfyvAopsRq6/G7FFsoIxl7AYQKibkW7S1uQB/2IXnvW1dNqARo
3dts6zIvjdgnqJdKRx7cAGx9CRvia0nHi+58JYbtDa0fRI71+qKVrFZQ4YIB
x6vmW8NoX/oZM0uINlsLSCWlnvaMT+217QjUiST+uFGX8cLYooStMBwYqY1o
jJhth3dyrYmGitjRq3oE5qgq31GXgvBQax5f6CpEh7DpGzzkMWrZ9C959XMI
nAg+bBYXbkQ9mIVnHLatr4NnpT6JsKuwMm7c1t5SICRV+KN0j9lUdEn8KlDE
v1QD4GWlY9GeZ4cx8Mp0vmSjG6/NFsGKOmmZsde+sMO3sGRHRuT7pjy9hYjh
qBWCH85bhJkJscvPMFe3eKmC4aQi3RL0hK47G5REu7IdIrRG9rbsf2zSAob0
SukdHRHPYVXuXlF/nMLtUP7TXPuhSwSYukpn6rJ7JJHOAP/oV5o+oSVW/A5h
Z1acHP8S2uohqDE5Esd+e4A6bnKHPuDwh4vlb+t40FxlzvBGq6pp3zSEBhUX
w1inkGMT7ApwRhVG59sx29VSm1H7P4XpcZ2b/EU7OPYF7Ph5K7THS/YFWA1L
nTdZJXgOjDaculvaip/vC9bqOoFPh9DH+dzTvj4qdxVstASPoK0VVGZrIPcq
UhUfm1k8FNNkzDX89AZJ+E85PdrNm8h92wkV5i+r22DuUzhN8gWyDKPWUvva
28OYhMc0dh8hdcYVJb10V9TwNOqN3lBveVhEOA6n+OHXMtIOfg4SAa7mLEWe
+BcY7iq0RwmicoLLFw1GzmQeQ0Unfd3Fxrb77keBQmzyuno7iM2PkyjDNeIH
mdzv3YCw4tOn0rorryFeJ8KAgN+ZiSEFJekb0RRBRs40vgJTdkTOhWnyzhZm
ys2IRI+VA9iXLto8vdoENYkWrtCQXkqcBFkh0GRFHzKyKTwCujotxEkyg6hl
xTq7c8s2jVpobw1RzIa0uhoB2YCVCFivb6dNsvNdEqsBmIh48L7B/8BKD5vx
NjnbBlSwGtAGk6RSb5tHQtPe/RY+ZLDyyHRXP8L7/h8gVDeGf/pGe1YTzd+H
ZfTg4P3P7+nQs2RDxUbI+U5SUUNBZiCafSOg9FXQ+hos6RgX2HdL68t5LxFL
M+Dy2jvw+S1GHWZ+qs/TsdrCPiaf1+hYe4f8JeST5Q//v7jWxPEeV1gaTA8c
aRDOHQ2fuLu5q97QOCqvktOHr0DkZfiMpO4zf6R1IpQ/ZMIDFrgPETdLj8gW
tOn7oEDxf2p55Tcud0VvLP8i1c1ve0cpJWcSlrj+wNPyJAi6Ezj/u09vZDPX
Y4tAire6cRW0Pk7KkEj4NympV72ivlbskk97btv5aOPe9Xo3DZCxtiAR6lCZ
71aD1xvpkjfIa5fsderDYDn+5nUCfHqis9GImAUvYaeHwNsNm6kj9Ljov5px
IibC/rPg0MR2SyERQPcMvUPy8VqBoAAZXUTz+snjGFgYFqXagEOnwO89TX6v
10IckjVvxEuU40YywuxUWJLN6cIzpOr64QygFL78UDAoD6rYGqMhdGWaQSst
vOR0SP4N/Y1VX27cwmt8ppx5TDYNooDAxxKoL9vqD134G06Ee7E5+dUwJlJu
iOi1ci3SaJSWiLwk+Jvb3wMbFnpOoNxOXyPykuwpmx9kQEERDJHUr20tSOoj
3nGOW3nwkKWXrl79hWjip9xrJJ0Ms9lulIXSrY4jJyw5WuYSlgmvX1n1ohqo
MVDWvy1Q02bTz5YKwcwIe5bUUsfseCZZSl4KPByl4wel8qhRGnZE0JcuYQgH
j2Aphw82XocaFlLfVnkRiyXK38zwP+DxmQHoYi4BxxixfNbICPnH1Et7vhwP
0xXnDKevkT2BGs3BY79dtWje96a7oe7/gtBCi3ZWgiyfInu8PcXj4hrYixp2
Yn1HSTzk2G2E4ASosdvBtsnxxVS88OW4D/GPyr9qtMZf0hOAeLZOSlqKZd9y
R6EHYvsqVFChL2AmiTILNdOBN3X4mXlmMuVnWi/4jsrauUR4kqfoHtSHAAMd
2oz5UuAyqkyh0cgXfpZ5BoE9uy+I7toJKdVF5jZs3fdh5DRjXMFal/3HMUhc
iBBJEuEJB9hy9uodhzvbudtV0moWPaFvannlxut53R1X6p8SH9u8QnmfFGCv
j3sXspfpLaz0vZkwLyYkZniVd4MGP2eL9Jqs3UIHs6EDFUMWokrz9IdhyBGf
D/b+tQ6LUkuYCj7yKHD+1pny2Z00pwbfuhtvi2xsswjryLqBF2ExYDnIP97t
YN78T4rOOKVMvaxp5HRQZXD2l8exk2wVA7eXORREh1oe6Xht66Czcq+JHma1
9c/cjaXPyFmdRAQR9hhON06Mt9gKnTuys+kDWMCkERJxyEDWbTVQoMvZEnzI
zFRy3J2KACqYt8Xn/BBisjOWVvh/op0kvzLI+0yORMH2WT/4mcpasthFFdUN
LIChdQGAmOEDtr6xfqvjEail5gBD2EZvAeHczQ6T+i91TtoARsb25sjpZVjR
tX/xzGVtvhXRHt59cgfXVI4DSpw6JzjZQA+Cfw5bXOuR6y3Z5g5MpArQWouN
/OCfIw49QRzzFx6w5DgZhm/nXjKGEcF7mhQGNSQxYCmAL+ttQGzUpQSG/xve
xrWmm0JYWPmuFPP/dbarodDMMMvhjqbOrTET22oVLAg+dNM7ZE6C0jcyqS5d
5PneRop7MnxLm3nNTyDiEFfStyg2vhwHBKVw4EP8sXolNn4XM28HhkOILE4I
ocp7wQ6asXXmtgmh+5RK3KPgSKiMA85RtZaL+ovTO4MGppJ7uONEREL17TV+
wajdMkN1fw1lsb75nZLXL6Gz4l1puoq6IpXcgFVntgKgJJ5PHAMso4S/maF/
DlGP6t+BRKr7BfEyUqH2lEKB51/Pl4fiJfXKmoVpFW3NB+weSmJwi7hyF6Uc
RMmNrg7iz03SWNH5khLXYo+CMAtzOU6Adgb/GAnixtgUGY91yj47ohUR5YvR
SjhhCIafsVzbk/LCCS20ZIavdceZpSEIWcqrXZEKnEeDLg0JVGrPOs07wDy3
jKUME9pHJtOnbYzSJv6yrMO8TjynlF19392hvLFLNxy+NEQxk3wzwatwA7RE
Gy7RGuHpEcRmlxi2Q5D+ZiHKEjN9CKbfV0HzwbQ6RztdGdBgd4eV1nHXAx25
lNed80HNIOQ7eeOmLHT0GsKLB8ewM9ld8w69XcwuM55PVfB38g3P93ktMk5Y
Aa3hq8ZfOPvj3iZbVrMnxvuWLZmQ0fVICCrCB9R9xNxiwGJMrHuUrh3emA92
xQkUha3DAXmn17a+qU0Hne+f1bib9BsyPC55KeYco2DS6ZoZVCGZ18Zxyc4j
9yY7LjmhicAlfKiT7kdfxLOPQbZprwcOp5sbQ3omHyLGjiWtx+u2X7DjbODr
s7CuKaHHdbNn5KS7uGXg+4eOti3t/me05plXrTPZVmAgxh8gcRd9KdhTgI18
uXz2PQJ8UXcnRl9x2h12Z8s11t/CJdiqu4viBum8NQBHjAyQktKaKWNN3SJX
r+oQ+4Rspj+NQ+/3qWvFF2c6Ln0MX2Hn4fZdITcUOLR+cbdzfVcK6cvDaeFP
3XOFrsuasQQn3efyXx+iUx7eHUq0yQB+BRLC0ls462X/NAmXVVBj/k4g07wd
MEL2c4wCJCfCznO8pv17c7+p/DW5MYwaHlfp+3SF6awYgbPAlX3DetmFd6Rf
VPnGKLy2XPjbf7zBEHBfCeuMA6SSo7kHVk00lHFhhSrX8BDxgSfarwHZ16G7
sOKs97Q3b8h0P/8LphA+leGem5yd9EfHrVgmgspoiX8japXG62CLOTFUK5gX
ZrEAfLhKnwiyxUdXk8gV5W7l8UZ24cDh3K4guPPatY92UGoU9eL6pR5nhj1z
GASLgBKeG1RMByIAoHCcddQaak0oYg+pIFkortabCoAgLHhjwWQ8JIE/xGzn
jnUNvpwDU9Uzk5m9vXEgxEXKQtxFdeRJsu0Yc0zqoO22uuBWllMpzEVW6IOA
sO9RQWpmJBlL6j/M7mgVFXMMCRvqzxLqLaQW6RRLzyfMezDepaCrlpNppxWj
9rjY0R4PuBybWb4GM7bhH3zmgVy1hJMHyl5bioMCBIBu7OZnGTavFT5SS0ix
fJSaL8tEjtQh5mCZWqNRhL2LD7lccBKtpjx38CYT+RRmK1G1oDFyX3OhUrM0
39GKsd5UpC3TqhJcwtol6uh0zrBllExOvZOnsTm3pDEM2P+gK8WiNiehtCDv
05/pzaZtIvuo75/OZFaOPUNY5/V5OTy2uPrz+A1Sdid3eawSHvVvAAt9hcvK
pCz5XYS1jfuWumsgTv8UgP8g7B1JDj93DyjPBaxOq84EjkYSyJTew1XSf/1U
uTY1Z7/GXzkDj4DMCpPuGbWT9V05UntkviraveOGL42sxvIDcBOHn2COf7Gg
KLKf8HTn+2KCUIpi5gMZbGFrDCCza2GB2YMsfzKKX7fapUaNqfU9Rxb5pPHL
zbxF+T4GgMBAv+LMGf5OVrAdUO18C5W+vJSMbDOrQAx5OGFSfVk8qpJ7NX0h
MEpDA6RaHHK3N8R7TPN4a8KAwUlhp9t7NhLHUrxgyzosVBdaXV2gv/GDWGJ6
1uMwJrCedKflRtXzfDI9jCxaQn0NCo3zs4yxovgZVgQ6XWy//MxCzz3hUCXN
llRN7Oua30segOywTQSSlZj6pQ4/0svdhPt6fDv0dpSjo5rrAzNVw1DkQJV6
atVKbc51RjGWTLjgBGTvHAVFmJm+f/YXsp3qs/tnPTyNQ4e7vbN14PFxM6m2
neuK+JlSgbimQgcZZeHCEgoxiznEwPmQ/aL66bT1IhyT2QksfcndBfnZ3tni
I1OlYKCnGg0PgGcG5NUy2zCSvKOSSBT7Dp5hXJeWV15Zh9BdrWHOrg3oYGZW
emIS/Jo+D0ndo+O3Ah3mx/okE8SVWqgpkXTBxVhrfO4d/KOWsY9cGZ/6OYm2
3Zp1RR8eKDz3/QR+L+/SVB6AsCq/iXaoDabH1mvofrMNKR+dSoKCmhTyQIGU
9WZSS2ZYq2wvupy0to+1ip3/nsHChzcTyLI++UNUqReAeeqsEbyRH+/AHbHD
zlwckbgWE8nqQ+NrM76sPioTu/4fQJcw8PEPJQxQ5o1RhYYvOkCOTEsh6RGM
I39ldcZmz+tpPixXXAeb1u/e2N6RNVnhPDvPTEZRVmj7k8RwKTvT7r5zW/q7
bZIYMiUwX3SYWurRPpyZb9k3Mj58HWhyyGCtoCGZntjQTrO61h62m4NZ8gql
hmGIKou4V/WeqaKp+o5h1OdzvH59mErAYEV8PKzaw9fnI+nA2JuxcNYHDlOj
xVxWlSd3aGs6L/rCBqp0/JU4hFinzCDAn/sw/DQJUB8rE+NtANNGTKB0dKWQ
sdbiqwbMcpTSMDq6ceJ9eUirTytOHKiqAebNRzOOrHmDGhF1cR7Bb+1zEXZW
uqBz0Qb1QUu7lfFtaUYVqvWCLqFpO27BX6r2nbMLdR6cswcT59kmqxGPhmW5
AlfToURkvwFLKv07hRnIMFeUZzibG8xMWBXkgLOzq9lRZvjEuzU8pTTPps6n
EU23BcKCR6Qiw3BloAKCNmvNNso/w+KU8RHd/PB7yfG818Vn5eJnJwddUJ2E
w1d4Hvk48S0y6GbwZ7A8IazG8WrJXdzeuB941Fhy1G1c8DoL8tCoxkEdVL3C
cPEJZU7OX/6Uiebeeki/nqepCqns/GnHRn6uGLMk20O5D7fxpwHHWnu15e8Q
7Gf9RNpMmzpvGVdTWbKBy2w0gRy92afInppNqG19bdQRs6QT/yOWih/vjhug
dOvmU8GbvZ8ZxklBrOh3C6GUVpknoA7qN/at3oQxi8pgNu29VI04k9J7/C0Y
iHYnPzx2zBXG3MSfG5y0n1ARZtcnbk+R9P4Ke6K8BM5s8IxITNEPqEe14eXM
1jKFV8nFiNnkqZllzXyjarOTIt3KuLiM5Ts0C8j87DU8jr0gPJoWrV3jQCb4
FyC9Nq718aOr+T9Gjex/0EHRLnWcMrKAzmH8Y2Dlv/Ekp5QuGyFdqBMnNV5g
2vIonYj7JUlO4wGMOnl+ksgvy/G9s4TkL8+UapNlScLAN94qWa5rg1sFSYLz
lJ37R/4QadOXUJ/cCniI8XeRWm6XA0WTQPTypaEvrjyf+nfY6AsUh2gCr/qc
bB/fg7BLpt4RgrP4jfRuPTQoAcEnd2fvuUWteiA10Wlf1RG3xmLH2rH9mhrT
XkIkM9vHY/zOiQ8R6KkbHkzzSeUhLOVLLkF/+mdpn9uDK7A+zd7WLUWGQoYa
U/4tLne2wDcXCuEXN9VLUZ6vkPM0XVQ3m0mCifhXQyFRe+7CwKyeA5o9iNXM
WYjJAmoBdfsDIqsamrx01aj51pe2B5CIby6SokHHKaqjhiTmSiQcFTexWK+o
rH4VWXHatjxy74WJQ4Fs2n6+BeJDPiZ9hi7MmgMt8nLB25KHEn1LbgTUbjH8
U3eCV9xsCEdTYZlHXGmsyzbd/aVeQtHbxzi5XxIKofH/7OBNI+DrOQEZd2iu
5oD4nQ7kOC+YsKJlpzJTP5P/w4M3DBppm+qKkP9dz6aBrYxtS0nZMruoNS3U
lj3givTI29qjCyEvT99fuv1H+6nKdFZIT9snMa7hw7ZpKR86XSNyIoZPvvmn
2FjEthrAbMkTrKiMqEJu74VvFMUfIQeQH3BDtmVzKDM0AQTCyoQ6wBviUYSk
rDpfUovjvb4nnKESKx+A7G1BBO71BFVNsWY2T6wHePb59oHfyFyGD6x5yYp+
aIT2FnDd9JHod/Nzgmq0lzWEws5rw/upXbrowtjijgzx5eJhMMnaPf2Xnzpv
e8E0ufS08G63S0tlJ2HmwVsk3PB6xLxv21YzM2INeGyQCFXypYIaPJ2B7K6Q
RiMjuWr5iQSjYe9pXJAF3XMy9/hWXOCb3rh+SO8OS0yJrGXLOMXI9BjC8PcN
AziOMCDauoczyEWJhQZqb4KPRswhEszXudkN+yK63ixHd9KznMxUhni0Qbeb
a4dPa138EwRUptgsqaSNoyJ+hsxMGFenB+dryVZT+BFN0h5+ihrZMCl4FUld
uU+mO1EtA81yijL0Q1wi0lyH+xTOC3vBnI4WSiIdmOLQcb9/27gir7RHQU9A
xUMJxZpzBtREGXUW51DPStzGPWW4NXsJ57TuaSTqnb2tav+BAJfeOnpWCqZQ
zrjs8M3h7OfmmPV4/ByiJuKgDQTKRlzj69e6Rmdx40tqz9JT7ZcOi/2n+9lN
AbI+wQgfIarovXPlZX3y6yINpTDsWcsfjdIpsGRN5HvPnpeGGiyRb42h+hXL
hE+RGIkYiYjsGyea9GAA6kBy3D6wijy1uKPtFjtbnncprs75IrwX01nyhn5q
yi1DLCFDVqhoJrXB8a9SjLgP9xFW/T8U6X53ajD4nN3IYthWv4bdP4trVNdI
9Ef+UxHugIlb406PiTJPKhunePKE9Pg4HxVCuPn3AxiCiZ1qjQrC5m8IPA3l
n5WjyDH/e+rTfYZ/43SqK2gn+H1C7YTlLaT/s77jnjl3YC2ok/XY8FN8Fhfj
oKDyStyYA2PQJcTDp1WqfkrxhZgin365PEpj+ZN+gHi14aLRz1dCC+2cs/zt
K8x/qHg2MG6pMbNcU1pSZz86T6ClsdpHCFmYmFT41V2jA5TswLumlV/9DL0c
w3YzDbHjhwyMdEkZPXFkmwZSspSVBgDUMjGoicWowEb4hQNZZLQII6jQ8YW4
WAmtrL6tAAJmGCNpSHo6EsXvt1VVBKdna8jVG+WbhB/83/huCvJrH0gSw/DF
oGRFQXMjgatLm48YK8K4VQTotCX1fuDL55DOvI4Qsiic0kVfEsCHT4tqRK5Z
TW+KWrwlr/zCdCFmMtKkQIzSA9x8Ha5ZriaTpIg1bMGHZvxcKGaEZHUmF82S
LQn/zxHShdmzwENbf+x1Z8BOMDKxzh0yrFpcntVCpkOpcwwYaE7gUjfq4YLN
o69UfdLA59bBvPKopruV861qJFX7QCJJ9bj6u9IaY0dRYaZ2v51JygTAU+WA
4yfcxSIs/s15V/z3wL9Bmcr2TTKlEiZR8EcbWHZyhmArdgxIj9jf9maoLO+2
od57H6a+Hngrhw3QXERTb0vnY6n+vMUmfzgZvoOKELrvNzBEX/tXxni6Ihuf
bkIdp0cu7TVbg7zEEXxvZvVHtdscu2UI/5A0aO4maHX5nj+EjbYH3TnRTp9/
xa3uuSw4VpDi2gl+8XQvvyj/zXFiBOft5UzwXm1hlFqbsBc3jDSDpyoQGWOe
jLkDV91wL9U7odMAOw9ogdTbJzgy3yz/cInn6sSzssus4N1Wi0oF6nfAL5ZK
QRayCQFxwqn++pfDlYfrQRFvj+JdR7ZKblVnv5EL7EOsBzhvKMImy0Vs39BP
XOFlegr/9EqUpENKhq2wOpcNsi2tWshesT/V/eXsvsx4NLH6YS77DINbyyYK
LB0CTK/5ba1D8tccibd4K8bXV+spA6mjWtoqSULvNxII59q29R3POEB3WufJ
spYHpiKvnESGRwY3O47N5zhvOHOWRoZ8qLFZcbzaYkVNmt7D/i0+AdCz0EfH
cgB+a2S3GMEjM+ac2BWQG7zD+VoL7fPjbKxIu0NdvleaAFR10UPXFHQggcpT
k7x3ZKdD4x7awxnzIG5i1qKOMYHezxXZCfBk6J5trOB8USmyIgePgOUixI5F
i9lV0SOMTgkpqdZtllhp5knOJc+gI9imxo1HCrJbL56vBj74XvLHShoNSlpr
LzP57eZQBggy4MSIWw+fWJZW12j/sYL3DRU1jSk4hyl/YKPztu3nXYbWweb0
rFeZJa/eUvyEXX9H7mP7vUkDjsHgIclzVVlqJBXqyOTnViprNYpU3JaLc0js
5sFk1OQXhi7Dw0P43CXBPEpq4p/7IFVusMFsf9QHlG8rIqJIupB/42xdzLy5
5NRxGuPMsCaLyWOPaCk21NVxxxfBM9FTjfGBOs+/hCXxJv8LVZpW2q4NGLAA
+2qiaukhII3+EsMOjZXpFrCMX7XgMZglGZ88ec5Gd7XkEBKdE4e6Vej8aLLQ
newzjxhuEl6KJMHdnlNCD/onYgJbDTu9lfYxs+DxcfzBH9vjmOwWwyGRpw0V
sjWkUAV+2LP9PXMb99v3QW6wd4qn5ljDXOY3hOeZB3VX0Xo3wMBwKfmWOfra
44Moo/934ETKOx3QB726B7GPUgKY9TdrL9QaEbMsPGWgPC9dEa90oEZK0cKT
D/pnROSZ4BSV7N07Wjtl5BKBYQcNGw1tI7plGu+uM+Puhs4UYdv/aCGMOpu/
Zi7BHHZ7cq85XutM2sKYxcnXwqByLmvO4tRptTXSy1ZvukrJNtSmtQ3QK8kA
0t3/wBiOghxirdeNfLfB8LH+Z7DlWTzCUyeptoHWVBnZFjaSDvJBbjZTOyCI
ZOUOMamClWSrVUZHOyySIeK7Nz8=

`pragma protect end_protected
