// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
WmIW0GnaqJfPDeej89HcTdBA6uE3W+GKSxt1G9aqqA1I/O21X0vJYTr3el5xMCQG
cfYcX1aGOZ/QxzfrfZPNd9UeZVuFd9M1OYksySIKyxBpUzKmQuv4mZ2eWP63e2AM
RVjy4I3QvSHbEQg97FXgGKlXme9WIbIbKQVdZ88yBx8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 29360 )
`pragma protect data_block
Ymu/uJboeZSd0ScM8452e9PrNyzcyU6F3oj+PM58dWsM8WSFClnwjsjL6Qff4Zlj
tXxmRp3x1YEQoS/dRMtDGrezoS0QeQN7MqfmFD9Wj8WKF7N0eVUD2G3n7hk/RWcS
p5jLIrIoV3Y/6GQyIcGKBDGcLeNHLi+1Irz/j9ge7QwoiIEB5Rg4TZ6qkPvJCsjr
E2Fs84ax8eLOattfpE5CQ2GKxrWeugutD9qVsQ3BxI/qRO0f8GlaCn69AXxPzq/E
uEsCL+XZsQpUSTBqN+/6WHzPjKFO4YlX5WDaXewxJWoueDxjkNZj8Rou6CM5fxCB
IVWZh+u2kGdUdZCuBWa/+htu4p5kYnXETXM5QEO62ajklb7eUaALO4eRnzxDfbiU
6tYodkk4ZFZCnuEamvRqhbnIH4J9RasAHx6QrcUe8HeW+MdUolMaCXMbKQaDas82
ImmYj05MApjJEm3gjaNmnfPMFUHqFrytOPZ/J5/5RsAmFw36OHWtdjQ3b0xEw7Yk
RKhMSXmzBtwHVP5kGip0d+Va8+XbZwOxLMqUyTU+OZvwn5rJPICBncWr/FFW5xFr
UzOefsdR5svNfNKGMxc3WSkV1tVMSXxewlUKnYbLeEJuQ/mFDp7hIAL592V+yOKn
DxTs0WcldrnVWgJ/iSbehgktGGtDutuNVm0Lzue+17bc52DpPLidhTU8ovT/MGGg
7G5qKVGqBI/8ADRgvD+iG8cb4lEyBM36ox1eAoNt66t3ZhISpRARU1IoRlNgPP5r
AVSJyG3edxR2BDqr92N/eU75C0GHb6zFenlLtueXi1IGGG6aoBfANwZ7C5ygeRb+
w/4vVySNp9bw7DS19JG4PqN49tyFbd8WEnN5fSD3W9tArbPwQkXHtKOksjpQGpZS
d94c/bLpZFzYMYN+mrEB5dUJ0ffPY3fl30yLAxaHFqZt93Upi3lEihLTg4My8hQ+
NXPSC/GFyTSv8kZURqhDI0mgHgy2F3Y8LOSXXLWKBwn3LGdDlW2svMwh+IiuchpU
4zq6ELAvzR8Sxpm8V3/EKw286sRs6SIEOMFYZO+YEMdUGTATAg95iDw+dK4WVk7J
7TOBNm5JwiEQtQILqsbA4H+QL6NiE5XxWx78UcjliwnbBaxmHSgpgGqIushywJmH
Wrtknx4FeqRp+jiUZqVykSN/mi678AIyPqJyQ4fJAAx21DlrCFm6Fl9HOWaEdo4v
RBt85j/2j8cUbcAdTsW9t53HpOQvXRGjmenr+esDXK/8CFnA7SO2wMDzOqc/u1CM
PJAGC8qEQHPDVuRIqsIYbWYWWdtYG1WA9dIUX4imZaovWR9A0zX/GzD5iyB1OYbo
BJGMfKXJvJrbHeKcSztcoPJTaaQ44VyPRlJi+Ciu/o3H4jcrogbImffGMuj2Zh58
yo8HqBhkxb9T0oE19Rc/CVL1Y+0HJxMX7ErypoLLClNjc7ZqjauRIOOLsiUrpuXf
mdKPK3deZpxpR9+Xp4mUj5tz81+zdsdH6APM3pYbGWU972igR8u2vxiahKce37ys
2gVxvi4lF+55kiRa62Y2Zxrfjv8ET/OUZP7aM4ghqxvzoN3iX0YDcweGAxWY8bc8
I+0ewJ6Xrep8f4w2UuYOBIyvoJE3VEFkLQ9npFtJ0chgQJvwhEsrkfuqd6nMwcFa
Oa/6sHtbVFGts7Xs6acpQ9ZPUkUIQguuvGm2uebRWPxfnI/3v/EVCQu7HjW/d6xu
CzbRdFRlz5P/sEReoTBo6jyHc2h8btvuwlsoOcUdZdRChP2oKzXVXwh3yckwG9wq
cY4KxJHioOY5NvyB236x24zd1XlMoelpmr4urcV+IHFJG/Bdr3w+v7oRrCxJApdN
QwjVhQzuj+b5nT9+YEnLwMt0UZnuJjzpqJ+3IU4LUVMvasJEhQqmZq/ers43Ug35
2yiuYyqxner6DxNbLxy2FU/CyHedcT9vNptshKm5zER7GuF8Xqgb3YNVyCGGgtrz
htkX9tLzyaNmATQ8/+Ul33m86q1cOXPIXkpPbL52c02W6sUlXElAVYEyjPmQEWr3
iR2GFl2wsdVCXokDfJSnttNabjZEsdBHskbY4ONZBMQug3i1KojVgDKyt6aXKjPV
SLPLfC7jX0s4/zr50imRFjlvM7/xgDYpIIVHRa1IVqEOW356apFUtJpqtFavma9O
0l95CPwQm5uK7Qo7qWcMrYz7teqB9ETS6dAyJ4VCVI8uA1G5gGsAJ3YxSwSMdk0/
smm2waKJM3BXqx8ovZwJe4sAPfvPf7z5r1H8lg392xvopoyfl21fUa1Vd/hMT37t
ByWtvVAH/6ZxuoN2yAIvVUeu7Bsaw6OglSQeCSj9CLPuct5RgrzxJ/u4rgobIHwr
awUwjPBmHWCmvHa7v8oWtViRLoyulg9In35VDQG4wk+YlcbVPUfBnLavQ674WQRT
nv2mMQN4wNiFgKN+zKKz65LxAGk0JX/6nEYmGmmyjOJm6g3xG531S8iybci+Up8E
KDjSLGoofm7UVMXxg8uDzPqddkIOwH8AIyduFb9FJ5BQ6NVSp5LTjev1Kc3Uz5oK
oyJI07ypAh07/IqNgjuIyksqO8Jxo7M8IOPCyKOUEJT4ErPVB1OVWSJVThDG/++n
lV0yL7a5AlYjUDg7NdsTXUb4iAZ08UQAggq9BqqjKPSzqQdfH5a0pEjnuTMBeSAL
vwC0Lvkzfp1XKVr0b/KQMhyDsiEtv4jan3RBIaWtOhoJx1d6GbN48t3kr/Dltauz
IYHCiGDpgiX1bKXeGA2N4iQPcq449FEHqiJbMjVeODGa+Rfo36hgybiz2pQkW+y5
DLhk71jyakAkxpx7ebjis5cz5OQJ/UDaYRGp8kbFpZq6L0CgbsS0gCcvc1itsL+e
Jl/DqEBkh5xMaitr/pcaEdH6v/ZLIN0mtpIl1fKB+tKNq5tWMYBEOjfYt/QaNKVu
n0GE4qORB+FCZRutvX6Y574/E9jdWgYyvO3YfUbl5PLCgvbBT6+bjZadThSD5+Pe
Xv4KJlxHrjQIos+RKOJKTUFPuvZOcJwzgo+uyFNtMPRONo+GDNyoYP5ekP2OrIkd
uBCaub/sALPxfxvZct72PrlI7qwUfPwxHHoyVe2JBiZfK91HVrvvvdhJmbeysYAp
OyYO7z/T+0kvPMu8kLY+fRTtJdTkbzKHDEIi8Z18xZkSid686H8w7P9byfoDXtCr
AVgVpU0DnHkL+8kNCj/wj9f7ICaYJ2+fhrGlhfBmZkrXWJGf322x6apKeBkLR621
dSHjHGSF0ESkcTunRN0yveHpdwoICBnnMXBPzz3NGzUDIwIzP4c2n5czYAeU6wJI
2QjZPBC+oZf6pUaog3wNrUQzkXDom9Jr3Vzz5RvxbNTSSegVc90mC6XrVu1mhYiX
D99GmnNXGfIKs2ClTNUZZ+XOTPq2wJ9h9V2BRPxnTsRV/cklLWRIhnkNe3ySo37I
8/6JUvspPVzgzhmDnSYkGKoXGQvCKLMIPlWp26dNvnueTQjpxxY71A464ods1C9p
oY5FFHPb1YvrDZ1VzEXheDyv+owmbHdVZS6LeX+TnucQoIY3rc5KIoke1MWr+Gyh
oVc9ruLBKrfbdsM/AoF3WMCEcH4Lu9rlLG9SXM2AU7F8Gc5jMLAuTeP6KRiQ3sd7
BA90eYrerk5qkrN1hlVQYqldEETVUW+PODUpXBRRqLMOjZA+iQrDOs7+bsvjgu3Q
cQzxiKIZLFrXgwzcFjcAoNDS5z4FCnEDtbrKLu0D9W+9zWG3A6cqtFG6YI6E7GWl
YmrZH7qtSzI5YxXCG3dNpAQ0pCgsXWtxfLqbEwrYqezRmBY54FNfwvHrIXVIhy1k
FqYF6Gyx+P8vZEheGGleGNQAy/MAThSqMFfNAhIXzKph0ubG6Md6WqQWlOi52im5
2IIFMpWL9MZfB5m0Z3e9WEexyuRJTcjMBzps8G146n/I6cE+wpz5i7IedeuyLoG4
14Fp8EaUcf+exYDa4hr0hxQyqx0vUj6yroDXmDbBcX0Vj7APAMn175yrD0OYXpNR
pZLyUC0TwHsw4hF7OkM1teiyn12t/qd7vBrA7NYtVvNGO3BTqQpjxClQKRyQavjh
rTJ+6v2gQLeyrnyPV6iSst4utsjsA7HU+LNVLWypkxYDvS7HPzf1NFo4YLL+Y07f
z73cYTX5ibfBJPJJhF74AZG2yVyMc1xX3KgQ5LP+H+qxLEKUafuUZEgn922sEh2x
vCzG5r2GHpzPImdrJhLzWYoYVyvLidXFJBaXyPu0eHqkceA4wNKDnL8YUjqIvXdm
mgPuB7WcdBtwhH5QJCk9XJhgD6eobReMq+w0MfrJZfPUAJ1AJ1XwGisFz+8fX1az
PTqRo+D50M8jmOMeiXFyve2ESdQfZqTNdeZ1GWly5dPYf6XY1QD96lugbfziZw2G
1o8lWFtpHf94VIaQsH5pP04nvpX1Ab9epe1SIAq0gszmtHrRHvbuYEEJbOYV2qFt
NplrFNes7QQVk0KqxzZF3FfAGyTGzGwzS25z9NimAlwu8m73dHEgxLIsZMU8KKsD
1SMv9aAy4JTDJfPsgWpsIFt+bSPLPqynGC3CdG+VCULvHyUnSgjosmuxei5A796Z
tzZYZt7+UUkH4x6+m9CkYG/5CFIdw3mF+bsUf0cU4dQmkTvpCKOnoGn33Yy/H7uG
67IcE4Svj/Oy2lM4sjMsnUVR1J2mnQHAqM5hcryyqRzTes7hTk2ig9aHYYp+DfzU
niJT/Xz2wv0x0IcmidPcII0/5p1USsKM+WVMmFM+A2GB3U8ucAeJu9gxVHR8siUx
hIc38OtgRPo8H0caoFQsid8eqyM/A613au9DcziFKUJ+o6Pgx2L+TN6n2Fx2DwNm
k2S/t/9q5/e4ccaI+Tda9Flh4rUXqW4zguV8aD/wU50XOrvrbJaUlX7wjj+Agnt/
y0FVy1oDNgmjnHu3Oo+GUDHv868NXDBsSIxmAEaALko632hhNDNYQK/K+VnHjyWW
zOXti8T2YvoKM4j05/mjaBJaNoF2c3bDAw2dR9kAHWFJbvEOpocr3qmIaVZJTwre
op4zAyToLBHeG5fJNYwJRi+t8kPPz9NDGJoXlayhZD3yi3GSJHpnJpB3frfv/XYG
a/dkkH+F09qFwutK034EnBtL2U8bybADhO7ito4z4bBvEN+d3hrensuNlbs4eod7
17KKP4AgZGcgEl4Fv3RZJbSm17I/uaQu7A4AioL8Hqa0UpZVhSJBR5jrzeNvj6uU
01TYoN9l91fXKZVR+4/3BdCGV79FVsuHUplwQc6Rklx2eKqG6Cg7/gGSDVGwZk5q
jSdCgv2h7HTy2VfR/pHsGWR28ZrKKLHXfToYGNElnMhVwzOA7+OedIzAcbrgcV5k
Vy8KgAvmJ8AW9x2pXvd7FWlrVFcsSRQoyhzPBYad1UVQ1Cs4GjVRquL/jXLJNQ0P
gCW+xVBjCcsLlzn1MDtEwxVsAZ9C/K2k8NIAGF2d1PAMEVCm1AWYrXyNbpMiZ5DN
hHKhnB2uE40bk5raS3uw8OLn0IRLIb2iKNzsb6+BDZU5Omw/NPwQgntMSgPtDb6j
7vApAz0Vpr+hloEz9YoZbJ94ob68BNzPAhvlSlafcVFOqrk0IZtpmwdCkyVK9oQS
TX3Iw8zSqkiusMqh6T8Hua9auHB7nOHSEm6Hw0LsSOnGKkMFZ5XARtFU3nGi2GpZ
a/vTeVPXop5HYnG72lcGmX1kXHLbaVHqvArLofT5+xxx6kXEpA9o1SdKXNMUPJrG
spWAVVyRkyVhfXC42VMBjZseqC9qSJAlDR39xAz7HQvHVy+aSSUDCnozCpobBmtQ
qolTcAnT+MWKgeUJawGcpg1WlHTUKVM4AEmUVs3ulMOOkJFJlVDr2dkIR1Jv4WsO
HSYny30yZZsAQoi0pOZ3P2ZsvPHOreG0JirNhMYIemDbwKE5WSeXuSOmGlGoHtCD
XdEc5GqMqeBpwEQa/rVEuduQrd7npngVlD/hUlybp1z5J2YTtRKZBZmXp2vg0mHM
iJg5IixE/bMb+iWpfRCkJsK0TEJWzRNJlZmn/mkiVVeNxxvO/wT4AkYmj2A1gNdQ
yKOoUjV0KSYbZq2sygEW7c5mQO7MUavoaoST4WcTkIU8BnJQvO5PZENZub8I0291
1S8L80wjyQoVjXOdfm7W1k6ZrafUIF6C+VgvMKkZvbCubV950MinxH/zh9UbfQ1y
6DMIpKhc3tO84pHH/rBUlNQPEdiPQj1N0d6Ti83GqfKM0bkZpwjk5LL+mws3Urdp
ePyTY/92OqFEXdNZ9PQtpNLyQh4dnb39hTq4NG7kcXNPBRsk/il1owNuk3twcYrx
1ccp4xKinzQlT0Y6hS/xIAkfFLKywIjpRqwHQix1egcWpauGEdr7OU6Vlp4HxCmh
8DINu1gaMpkLtIsWtpvrWpV2KAHL9RnyO9o9QLGEeUJRUYgL8k4dGZdPiERWUxLq
eWtkJ19coBQCJkuNgLY0IDTLy8XROHY8BPLs8161QPA9pyd/TS3O7o4LWoeTm2pA
rbZ6PerX4Fs6Eh57ClMWgy46mogaSDAy4BQrXLPFl5Tds36HdRqeFSA+i03mbEXH
/0sVyoVxw+aS525cn969664lj0Vx1EqUXlytlcpyJpCTq47xwNuhqWyJNHe8K7y+
0XjUUStOA9kL7CUfTDlEEUJroF9LNuJAZEbxIU3BW97ZM8kgBsCdLHGZrfg9i49k
d2NIRASMlr8JTRkhAYDAREAyZpOuoJFXR9rBxPU7O9bMzu7aWrBZVmYqFy3gEDON
UmBNTM9Iu79hOxepYMqdOFKTVuPTePayWQHde6Mi1KkLW7lFJeYxRQNQmaOt+mxN
JR1rZ/MmkW2prgYhq2TjDjGMt2jSNlUjBJsGc+eGmFutx4hgFRiuD71Rf5fJqg40
8cghWWWKBJ8NtUEufya2rfiXRZL6vKMaY1MdVJaF26qXp8YI8LHGM4BiP4C1+oAF
w2Drr8KUdleUPgoyUeLWJP8Vwx8ocPkNIr/EGzZgE+OVjDflamfARcquFLBqVhzX
yWkRFiM1QTynDem0eJ5E/+RnM4WPCrG8cEmZBqwCQT2Hwg3QfGCtSLwNE4+tJGl0
J1U5wGZcN/GfA778bs7mTvMoShoovkBxaanCkYZ3q5tFm2OzfAAF0zqZjLqfLNDH
8aEhdK88UnS1QCqpiBF24rF954e+S80/C+e3RepugLnj5vX3p0KrBCbfWYcqN979
/s0bDvdtrmwNdzZsmWyzWiXIuNZPrsy1d9axo7DqQzwp1WTyfk4EP/b7foIy29O1
wiKdQiLMPipThhfCRUZvhW1Wyvjvpcbvm23pTbt3zJHp1zf/Mhps35fkRrf3tq4c
H1ZQs6E+Byo7ghtToFUCAX+6LyUa3v6sbJryF7PL44WmYY33WADR6HiRWPsyxRSb
t6fIUcMkXhFs8qY6+t02RlsSfSPiEiJAM8zF2SyNKKn3JOWaQ4H4px+lLa5Y7v5V
XtlR1bUX3WM0XuXR7ClTEnmzV75G/pmUG0lIBr+m3CNnwh/FOXNRYNdMMgd7vyoe
N3x/hwEsGsmSirQe6xr4AC6YsYo7LX/1U00z7lK7abywQD+YawuuABxHUMJJkY0X
l5zdSyFFCaBUOgr+RK5IqSTHM8gJHJ93YikBQvPHt/e03D7yIm2Hszy7m8AKONCM
oe/4+qzz8+GwynI7ov364VjG2uCi9C0A5PHwRG5r3E9l/UHoHMMchSD1bjZBNJs7
l/Nvs4BsmL6V30XBQfkHFSKho3mMT8qG1Foc5P55neD0EByKVSCLDz9plNodSAlE
anMtQFxuTlWz73oWo1vLE1oHzYaj6jXFbJZairBjcgcLBr8sgaU8pzb7bxFcvoZB
4jR92a5xhPhegv7XIJyErBB10rUT2d6QSTQVF6udDYbIEie40lp2TRVGaWLTwJlD
iTErbqz62UyerNUcaCYHID98o3eGIOGYRz00oYye+Wo8ARgKO6gFwGjwNcdO7YXT
/+kp3iLc/6HlMm1fVQIvn1CNYy64rwF4FOvQIBodDdHYQg5wi21js3AgWhSrY6BP
vdAAQy3r6hfsUglP11eQeyMhhEwNidBIApbftYivGEN4RzapovnwxsqAptizbtoa
d1RLmHDMCHVBQmB3XqwfOPMSGhIKgYMh7Kk8kIG0Sp1JHfdqeZoNwHZiW25y8vnG
ty+faVEHrCFtAsUt7yjwUZ15oxu0dos+bUGnhKVwDqKhUNp66TGkWp2v9FhDbXEZ
9m9YuKapnJJK6XX0J/2kzTX8BdimtFDtdCuxc6BjRUtBtBk65pxFcXp6IHOiW7UM
Eb09ZUefHzCpXB0JUMKSMg58saBatoHd8mZVBq/o8dFvUEbR/a8X1Ar+NFpHUrQD
JLWP28Akur090DfyRr71joLtM5bfI/A+6/nvpYYJfaZGtwk0FwLltF91qaI003he
X/ugJSkV/2ru0XvTd9B4S/8SajeNp7xTzhhdWKuvrfENXITLBSw3mQeYIKsz55mA
oU1ZIQexDPkK/Kiu8di4IYuliVEEDqCMeS6o1gzpRSGF9R9jgiJHIcuDA/m6JOfQ
ndLpzVJnTlsov+FUT7dDvql+/DH6j17l5IPDttLQkK4wBfAOdTGgDCsKJHcmH/lE
alKZnCg93NhkPpxxVFJpriMMbhikm/FXYSEv/XWs8AZmlSPHBUMzMYvkaOXnxhG/
/APYJCtzbeLaaBd9mij2VxA+TygDVt4oYTbpgR7qIJy19RFMVIUyB4cgp+ZRzNPG
U9xX8uw1p5Vv2keYjVNNx4VZqrtPdknGCv5m2bQqsbr2HvADWnN2z8uoqlJc3cWD
Y+wDw3SHRnfKlNieqmQ2+CXERHn1MZfczfq1DGeTyMBoqiTJK1gzZAX6MlKKRx1H
a85DyVEO8OwE6mPqc6izVPbOodOyVfg+WdGkKVG1kUO+13uKrlJ4bC/OsQm1ojks
FZT4xl+/pMBmxGmN3mRakpaXGUvfTnXcqZ43fsAb2EivsJRaej7N7R34Yw3BI8Gq
NfrVCQEceR2VoDezba4MuyuqSnp4htoDMo184SgsI2cpjAnPYqHIqd+0Ownf+U3y
pCe2RdjfLUk91LkG/RHkOi6CkeTs/fXg6c5VnAsWAb0mYDOHAuYObY4c1py9VxR5
rX2wLXosNX0CkwfRNoFSrwRbI8sgUP9Xzqj2Ev2avFENzvItERdG8iUbn3MEalBp
BL6oT4PT3FJbVdH2/fDQscHfEsiPUfKujX4YFMSDCo/M95TAqO3rRKxwYiDoLZ8E
PV0JV9nqsN3D7IV+PhsoLSQtmHjAsJGYtBRmCqDoWfTy3WDZabNDzeWOQPuFm+bt
YjMKr1FxwevFHXUAKa8NKCaAR9sk1UOeMfH9AN+l1aG8yFM+x9zn+xV00vu5KeQY
nRYDKCvhZmfiB1RFBx55vXr7mBYQniUqRiANb7AgswmfZqqdu9n42C6UsvkYC8e4
T5BDfv7VX0NJGhkHZNAndfFKvsspxpQZoGapeGuJGcE426ZQ6BUgXqKygdu5G+eY
eaAx1JBzm7O7VVN0jye3rMmsL4di2Pmr87gBT0MfFfyjt28dYGvB9SN9HPxIqrc8
Bw2cUST8gQ6CF/a9W2sBcAwQINb+ctbk/kt56a3nH6wlQcM6ejmkkaVvEy9CUSaE
uCWL9RIzO3xV/ij0R1FNGJaHecPj0g9oCG0nagEkqY15Q2C8jEKXbCzidMMkmgL6
Gc0ibOB4rAawEzqkbAveldpBgMzJfb3ewM07hWKriUrj6Uij/kq7x1oTfzUfAP5z
xuBMunChnM39zKU4v19REb0vEg18x2MzrOi0gtG7PvAlEiyZs3S9TGPotpFP68HF
krFiEl3M1h7kzxjEF6VlWiZ8VEwmD75w4BBIZEAsmQ5vWkQpkyhWUGfy0lC09ene
ozondd0OwRugfHtZSYgDdqZV1xw6Smg1fp+zMVJtRFPG14YeJe13t1wPlOT2NH35
6fox8JP4dA83HLwNxRM29K3c1RKhbDKXhMvbOd3irGo/HCglnnyYjEv5naFblahL
Odi7W1LthrA964ZLzCgt0vqdQL/Lr/cvpdresRD4hjW0YgrG3XE/IP6y1wN4cwsR
LWHfEKVf0/5ACgYiK7EgmJnh4jTORd1II2zYKbEvRAoSwgFPJ4Ieg5QdNgUrPySx
9z8MZyXn24L/e4xE9yol1zZNrioaDdxOZmw2Qnh0qRnKv7kigZ1G+BFr1vVohXOl
+HLk9uGWMhNc59qjjSkDQxYhbG6Tozn7hCj/ZRcFnuejp8mWI+6nOVv2kAyI4xNh
wMecWvS7V8T+c/sX8L1l27ZgvMoHyFtVCdqQ4h8fGHQ5j/cCl2QzxX2p+RtwH7cP
ybLL1y2VIEftIWck1eKMMkbc/MywtDLY/FO2HeiM7rh5+XVPk4sURiGJbuBAW4Bv
p88Vm9qFJmrMqD3zhEUMR+rYlbtsjZ3lJ9ru0QsgBnYGu4VQYXZWy6JJUuPqa8oq
8rR9ujNCyiGL8iXQLhOKJsyYYimNSmL+JhDSV/Dxdm+SPMyCFkYXp12IWQ0EB30K
eqQBG6l8cLGPbyBDtUVmtcFbSlYcF2xg1p0VW6BzW3ujjjqJMSaZPvsYZp7rsPXV
Ocm0ASwqY2+CNEvBrgbCMbxoOTvzbmHDVjKI2fRCplCDlkA5PbcblziwBKVOo0bw
+gw/DkBmRLgeIC39tuCQ0EnC8KzwpLxjBl9LzaCSLa0ZVoW/OJD8MFp6/y+r7Rmt
1wZ/qIOXIR0z6uzWLfH4MLGVKEGTVlZjpOAv8w6lAIJ9e/9XELodfpswE00YfheH
m/4JVJVdKOq7dByjOl0MjStnHFrsaSDouuhwwWC739iITqW8Vhs5wdq+yj2ffpoG
BWe86iKidtNsaeb+ZDWiaT8aoa2LHd0WvJA9o5h2DbYDwI5ev9pwNxilOlX9bg/e
11rxwnjveHoj2rt0FCFCqi7ZLxNalla54IXZA2vATobkEmxNvU3hGCvrHtg98W2B
UdV2b1N1IYlThagzyYvurRE/J7Nqfsmi3fXDmCOC+1sgZF/DDe2idfRlK9RpJIXS
LaZCFdSAONbTuKgpzXKx8IA3vJkfnKm6cUqScdPieoQKg3s+2cALWt0dyMObudFJ
wWKhK0Y0Ic2BmxfnwB9YRKRnZtoQpai0/W/iV8CFDDq7CY7WJi2fRrJUr6FhJ/DM
0cBWKgoFTTkwntqGZbUZXkWd8nJM98/t0dNvnboJTG3eeAfO0EHeF2SrHXGAq+U3
+uD9Lp5VIT+yJeAJjLZ3pSjfo8TWcts+TObU+Eq30in+1tykMMm5ujtdf6bApD8X
9goM9ev5VRU70DxuStF+R9NqI1U4MRvBdUuhV1UYUWMiuDELnSvWz7AOJ/CFBwRx
mLAgHx3Bgr78nN+o/okwpdcPGm+5TNWAhqfEVPRhjldjNbhG21WMSBbGh1ZWb0iO
+lOgCh83nMHj+eFad0jE25ZOae4XVsHt4p0SaLWfRmf0ud0OA2hsd80YgUHS6oAy
cjpMysNffwsZDTHGVTZMdqErQXth3IDjdkuI3N1TnTBb2tyHQBdKYrkuvkxbS1DF
+sCmZ2AbSMD/WTxUbhwc4NnUQf1ubfyL4oU7oLu/fpMqLyNyeyMhnlwM+37c38eh
l+UPZxkNjs/6QTwSp5JaXmpYVEQicucE6WFQA3KJ4TITH6FqNt8GLLNaKPle1PRn
REH3aYSMDSdVypTT9Oe5oJ8ZElKK4ObkxVnEhvwyyeUxhKjtTm3xgFWizpoT2mG0
tP8a3cWk8XatQj92cBIDRcZn8V8rcE43WvM+fGto7+wl2Iw2bY78budJvJNsJa/F
ewaZpLvLJvVG61GC1agz6IqxxjruN+WrOCwAN7D+iWP/J6n63v5NIWGWqgEpuCmd
JdpkH+IQKPRC2FggSdFCO0k+3466GWwX8COWWWrGrSNKbtxzuYp4DtqdIT803ELA
quGS/tOE75LhAs/SMuK8gZ0K5R23brbbhwCp+v1oAGp54/2U9U6LsrbLA+4+Xouc
jM2Q0Zhlnwc2wQ/5b+dBZBkSfJGyS+3pVsaGd5s3R3NWVLt2IukAoX7Uq/QEKj7G
Xi//geSBSmm7h2e0ITMA3uu1/IrWJ0+vMuep0lhfjUlbmGkJrCCCWDZsrFGyxjy1
F8WfPyRx4mq0qL512LO/ecImLpAMmDUcwEyovE3ilGgGAvb+f8WSilwORjtpAy+K
+vrOlVmZOyfEsPlC9Udr1NAEyRdYcg6/oncSiNfheQDEpyZtkGpFgH3CysWs7d+A
lSssFo/t2I/bFkuKCbG5iNDmAljMf2UTdjAxxO2reF7nr+5pNwN8jdc0FkMn9/qY
Aw8zstHSBAZHfh4RpUMnASa5B1NiiP/5k2+nIAV6J1K5zvyeEfG1VR5jddMDQ4bn
jr3Oxi7VeWeE6nGjMePPYLB6XqQtuEo/08WdsB3QZ0KDGpaldVUdmL7RdyRecqyC
v6c5FfWiFdtbIFM+q+VT8EJV7Ioip0xGU3I9CEvdJS02hI8QN8olbDGYNjO4BXp3
NqVUzKcm7ICnvdP+Moj9zHMapOPZoLDIbdRav31sgsS3sCGBniMjap3/jeIv2A5t
riRfQ3bV2vA6Z1UjAxDaR+92Bo07rbj4sCg+hslKB+Kgl1rW43QzAIkW064N3C01
tRDW5XH9Yfx8RUA/7XUMVXSKY2OB1DQj6jQ6bgCz5Q+KOUNprnfdCQC7B2pvx0Wu
UB4Hjg3A70CaBSxNXHpmqiK597wAe2TuSWoE974C/en1eoIo2rBBLGA+mCgAO7Ho
0n5k/oloS0vOvHvkUh01hKFJ3dJnbdGODQm4yiaQ38YmhBT5zHpmQeuogkjh0ZI8
dA9TZ+lSUOzkd63IdbonYrovkwRYhOOSifGQHFJBg1vXL6M1XMPOh1lLBmAVVVHq
OFhyQ2rPPtAaok8b+jRAutvshpP9k8nubqYvdJycd74dFVpY79d1nFCNzcPMIN2u
PQ6XXefmUK9RcMgMlWI/QMgwUvarjZx2oKEIcCTNGUQpU/l1b6Lt71Funst5LUg2
/BUS0RV7HOt82oQt65V7Do3d8SRlwFqSgtTfUnR4mn+kHeaDEqjFVVhUlBnKN+oW
i1WXYPlS50aUjPuFLmQvLHr23vuXOBLaHg8kRVK+BMxB/5TnWzqTrCl+KYahnvmY
8EIRrec9GoFYexC11iumcBunJA2Qfw2HWlDqcyRhOC4W31iOiXjLBTZSDC32QUIM
j0gzMsC8yD74d0Fc4UNbQJqbYSDKneSErNMeYnwEXT+bRuitqdy84X8EUTFc+fJz
mxVoJjLETcNKka8l1EXF7dOEM3u58wxx1rNv6qWX3ie80CMAFiDbYowl2Hqdgfc4
iJXHqMFT2PTXUvbiAhtAnVxnRGAxi4CjEo4pvf5gsO+6idTYrPJCMUpbECjCcJId
uaIm+ovpHcGAkNgdJC5S/lWY2zN3tv+WwfZZBIt2ynRZoOtzm1ydPag28mIhoM91
9YvRUQ/IlMMLFDq2HK3vFqtP4VeVW9b/SCO+etKFBzK1HFvE/VYNn4nN0YvprQtv
qGsGf8kW6xcrqBVsrtfrTw1fEDDmZuUQ6IxqtRomA2oCRoNL1zWAeaVPYi6dM2+O
OqfrSewG50u3Jf0+qCNxcpXjL18PSZGFK7Wu6zyBWOB+PW2pwtGUX2mzpdeXeWNL
g/7cBYAP8CpkL3Oa5XkFP8tzPH881zSxrYk0sw8DEmZ7C1NLQlQEJTGxKuKkAesd
FeV2/7NkwJGJVsVF9shsxRJfVSVZdGW1CfefB2Q9HATvaRnHiZLtb2u7weU1JGgL
GeYueeTaO3U96gW9dM8eGfavaTQh9ImWxCrIwq8r7sk8sLemBs3DNDYsWNwMvkZk
MTH5t0IcLEhCJmX/VDIEbonK34V6JwYl93qipTgB3isHzI64R/ziPDSUymOiT2H7
vR+ml44m/xQk86ykpXUBt8KnO9SB7teOdzaEy39k5y8gL6UiiLAn/QRBxmuQrCY3
WMsH+yWbvpv8HdSeBnOn7STobS5DFeJX4lRPpZqBdmXFXbJMSV2/P1UtZmIutrJM
orWc9fJJAUCEZzcUaOGpwvStdvi4dWOdQlAuphPByiKZjcJCIf6drFhrIamX9uun
l6uYX/YRWLIumYzQS4YxB83ij7+4HAgSpaHLSOqYy4FltlDq5l9D6PBW4S0AlnPl
D9B4QSLn+kxiqwTD7ogrDmrIr5QeMKAmDSaFLL28O80jWIFndm8ZzbsifoPhQV1Z
F3LjIsxEXQr1a4CTdX/oEfl8rRSNyF2S3Z4NHH/uZFOpgpxwkj/EVM424NuoNkqR
e+8HgGFbTUsktk8LB9WKXmlklTpon9yKXVYolYI6GopCbHtWo8yzBDMVgyKtHQjp
JRizVCNyy2V9hxibXcYklm7Q/obUJpJ9IIVHja8D7Y0+VK2MquGRLfrU3ldnUFrd
beXLev9HZrxP5UpZ+5XGCaDHnLronGjjtWVUehFN9GhR6mVG/jHKjH5iiaxzH7Ma
imhF89P1n/b9t4Ebw7KoLxCy3r5NsR/E9ncT5THXyp3GYP9Mfayq60P5m+j1q+qc
QvNexSJmeDrh70GQvYxm2Go82mg6eiISTqDC6/ltH+Wajm086UdXPlrbVfagty00
SeyJvJXlrLqpM7bRdE0t/J3byp+tHUs+aR69hM8WZiEt11m7WdSuw2K5kcrk8YpN
SqH9twcX9yGfQpYx2AqDMQC9GpgSQKpUgNsvo+92LUdiiiRiTDH9Hu2uFbjFDbli
81Bb0dXE+LC+NF7PioReAAKwnucjxS281+tL8G3dktUWFUU1jz9gecB0/AAY9HN3
QZ+RhU06tXBXKspig67Yai7hffQLI0EC0rY3Domen4rMZv++eX4ISrfYg9ryx93/
M5JS/gJX/G/1bNr63beUAgU7WzclhqupzVqqfz4QQN+SW3Ir2lMN9wqwgWc234hn
KNYhbq+I8VKQlnfnZK7IkfuBHcmwsd+sKnKo0VJ2/Gj0LxHSokgnYtSQZGkwURPC
SbMKveamzfTt1/kOfL2ANPZcBd2QSGHwDxwZfcWHglk7rK/NTtyRqZoI61JwT7nJ
Lg5ybGkWEGkJQCwSyro+OZgQXlBfozvED/kyftS5Lkcs33KQYvW4A/SjZTeoEzR9
jpAIgUe/X2uWlZh9PBFKQdfoFOwXhyNv3M8YFgD5ldHSUCUIi7i4uNMYEjFHjoSD
cPItAqSeCCXSLSBY1KVXS7DX7Ge3R1TATB+QhcbCK/VRf5BV43zXRn9TCXwOuPjd
tvzns2CSU8rMQdI+VoFx+DNpAw6gnumWhLdkyBVnhdv+Z0NIYert64aDxqzE+M+x
08e1m/a7C3qodj/n+hT1zKGm+iaUMuJdgB1oXf2SBp7A5atYVjakCDy4R1lAzZuN
tm3HIMjuMJ8yJiabAZQrBIqx3JmeYQ9i4P2EdShFXGzvAyF4VD25PiGvc+uh2z29
iTxDFCBLogAForHksGF6tidiTaXI5c76ZrRa8ZbVyRKEOUZBkszDpjPCOHBWyQiI
wTY6yJVuXGarGhGW3xT0zQRFmTFwIfu0gGmUS0WXAKp8sGVKLsHK5jwZqX2j3S1b
OyZBZJ/+dDkIUFKCiCHo1apMXUinGf2KUrt0wWNxccSE13AhAAR11EjoU1U6IL0S
P1FvFJo4lFRtvBl1TMUfUB6h0e1Z4xDkQjTeSncadNw0qC/4xS4moH6GMOdKQYGq
Je4MD34MCIHgGx5vzbeEVfz5uEtcaPLR6+dCoL3UolF4QVzxmfv6N2RT0/jtwMGv
/d48dJ9jwUeukPvmj7yRSv91jjLjdY0cbxErnKV7ZxQh7NIS/baIYIrnydi1/e+G
1hJR8R/q8A1bf2on5A91+NZra066Per6B3noNgwvjKhs6B76jaqTlrGoKm+rlFUU
y2NdOpUvfeICk2tCJt4537856SgEH0sxk4pJvLzSUWw7hyqgjQx4AeC4ncPxjPn1
GnchLFqGjOkO3poOxqj/rol0yVbJA7ZZnM5fW6qr7ag/ALv/WlCKgejk8+eif93V
MY7aLRKYVi5+2xbHEEFwpmbDx1qHpEt+mxAIrN//mJfZTAeMsoaDYbMSjOIvrvJz
bVsra42ymU+rCkDI3bZnxM5GDxVGDP2iEgrq9TE0/U8tYO+4Gut4sZWmx3QvVnny
o8K1RLiNI5QoUrCgsHEKpCkW3rT6z3QEzU1yZWxahHP0ql7q5lEwV53bXV1hEChC
AnVBqJ/3d9UIKLQC8T3CM1i5DKSwnz/06q4FetNcG6a+JtCXJQGcJeerGRmiVKEl
+yq9w8jUbc4bmDhp+6TezLWV3d49y8xb1mCjel7PfQVP5BPbg1skIAZN5+Ua9qGc
vCPDHWSRKrJWF2b6AAQBM825V/XYZLWR6gZVgU6HMsqONdQCqr3YcA3IgK/GHYHI
IodGWsvatdd0Hi9RSrM+mrJRL+kxB7AfT4G9QZPlzrXbMbbc5hZ8AFWmhTK9FJYY
5kRwfPufAPDWc59APUNJ3vZKv9EgFmmuDnBn+d8gDRmob58EZJNNgWqIBuLUyk3L
97ErH0ND1FcTpaXgiNQZBrf+44eGYbG2jCgiMr4PtGVFzYNRXoDpNLS9DIJa+Gzm
BzH/iV7XMrJJJ3MmUKV7TkKNKkAkKf9uj64NKYJngafF9fCB6ipV0FdB7y8Z3c1o
TfHkEEpqB2qTRznsNPmhUy+TM6NhChYRGDxx5mFOszBYwcn1ktnes9DpxkE1+yYu
x3QpKI+cKTV8lYr76GGVoHKmH/AWrP+0ngBtmN+BDHYIFE2K6jxtehB0Bk160mSA
hFzPUbCaOJ2hVjwkVdgPkXtLvMBLX5HsJdFO+Gc4qFcYoPXmh+v7v5aGS/cW7NGp
p0E1jnFSjr+CH/O7RciZnfLgvL2659JOKX3mODOv0zL/4vRPFIuF2dTR1V8zZKaN
u4dpr5vUKWVzGuMTRB+Fyl1oYzXkxphGT6naZMUlCdooS88IAHgojIutqLvOysBr
yH/I8MCdb4qcw3EMFnxMFAdiUcf90+7A/S5piSdy73bmWa0pmNlL35yege3LAI3c
8FCx45Iaai/LJgSKpUs6LBkv7NneWTj03KX/52XPLwoYOEOpnhTE8Oz1gTIu8Qgl
Rv7JCTH2s9BxD47yxMt82d5YdCfCnL/HXjxzwMXsdllT5cphQLCDfBG/p2LwjhcM
m6RCRTggTz9cfgPVrqWDsZ5NQX6+xsKd7CUfmehvX+hxXa533ucGTge5F3/p2KDY
qheIsmJiXYmo29bZQj2DAYWf1Poi0savKTy2LHVYscvcffRPv9n5pOmzjInQCMxt
3LVt3YDQSL4o8DVxKfcpEvundthGljvsvy7Cs9F9HHZMcxRNWjecm5eGZa4gRQl7
x+0TgmotMxlxIehxcX1ARj4DjPkE/lfhP2uN7aGQ/qnri2MJZ6jrQ3qnhdsCoi29
YfuqPy6iHb1qYmRzPAeCVj4MbKNkDgP9lcaYIcL9E40mJc5SCsygCFgWK0O//P3Y
CwOv6IHF7L5HsgYlaHq7vWhUHI/KDhyMS5LxzCrSJpYq0k8O58Pu2WHgLMLardHC
KMAtwnbv1KVJzwX277JXvSlY8t15mnpP1WjeZ09Lawyjb4+td4JO3NxBEfSLpUnv
3IfqiGhauKku/aveLQm3IlH4YOjaXai0GIZHieY2kWBKGuJO2s0S0e8MF1jWj738
EYvGmr4vFYsWr2XBTzZY01ocJQ7+x2v0Iwjd/RULfCoLOyBbQTuNmiOZPiwSfUlX
4CMrHi2ubRyw7GTqTB8atXYr8GdrQO4hOKcvI7iCpTQI2dABbVhm21LDx4aclzAE
rfdC0cOQlEe/oeLVxcuRt97glUxmjV0K5XCuBdGC2tp7Wc2dmv8eQBXLRL7xwoz9
CNP9bLwXsOIVzXUukq+ZIv31ApYplQ2UmLS+4C8FkRm0eHqdHpuBot2lFYhkt3lP
x4LqbCMtiSCem7x2pD5uDld1SWv30v3/pw8n0w2L5ZDE/bx4zM+k3e6euxC8HyLx
uIwrNgq78/7NXsvsGPDOWElXm/jfNdYSNX0C6YT7UTyk5i3T3zvAIOG2QIugCnYZ
O1gUb6KRuW7puq6hpGgqzACqCUe8b/AzMVXRm15IL0/OuMMTi0IMepCqZwyCPckb
2MmRV6wYp/F2z+l7Hv4DxIQJqa28ZqIz4F4jqrjU5S5sAPz9Xy7RGuczfy+7eTx1
9cVtqkuLCgnD3JfkO8kZSSp2XTMPi45iksDrgGL253wzl/Fst7ddGKfs2UWgCSZY
koQjMXEBon/1j8F011fuJl8IX1MjjviD5y+7QaRKokMxHu+cI52hLaOvr3f8ynzF
8WfnsbhpA6ihRCHJgX9km7hXw69KfPe6ZVtIyi42bMsMuae9vGKMouzJH96TPB2B
4Ml7JstjOEDNRVk01l2vGxN6WhVmoHeiDc+EVEz97HBOEHlf7rrtQGevfU6DkMdd
QzVBTK4xD5xyUi6G/Bdd9rW149CTJsLufWxxvg38P730s96iyX5rNqWuNEHyuXoN
/Pm03sfG6s57j3LBwl+T89jJfrI7G7eyUdbprhFCuLx/qrRBsRnTBzIJegYLoT+S
M9x4JR8EW3qiyH/Foa90eZ54Mk9pmPPigg90tcaeg9GBq0dXbfQc8j5gn0cfsxo6
gbAudhyMm7WuOo2/55HoIAvvP44/UI1H6ITFy6tTfYCd9ZknsXREG7WMTCO/JpGD
amL4kSCzONDd4BJP9o09yA+Odjm7FHA5vIHGpOV1a5mkYwQMDKYKkjzsMHKfhKIG
AbDDVERlXlYY0sXHrVY7pfvEYrZF4MOGBCzLjDGbRIzWL6/5rW1hWmG6+S5g6gcG
RB8/7WLfn6Sz9nEz/o+7S4LzeZ+OBBnlOQQVqznlyXAQGpHKj/goXBt1gWYrL2d0
87pfV+FLeyz6CbLKnaaBZC8YtAVFs3QpJfzo0rU2+DpywqB/4hOHUycr+X5IzalA
YZTGLuUAABC8tBAdsIL2jpI7Q6mDv4OdVXhY2NyvLLBf5rvnZ1qWZOPeZkBf3+c4
YIPiTQ9Pzl3KmRP1h3q6zPBharRvew+T3LcgyNe+IJ5yIDNSn3FaZWu/MKI4cjdd
WzlOVW3HMvxKxAROrWKPeu3BA3KVC9ZKfvZPpt0zmEAKodw/PfPClYXg4H1CsPEY
Rws3t3WDOBf5H9Icx824rZtfQFWrY+/xsxyJbVbfr0w6K2zwwzvMrqWPv+/TuDgD
EeDhSXmOg74BRv3N7fRaCeUhysIUp7oT4JPYRmMMGTFUY9jjW2fBna+bx8Sqi4do
1wdWW3LejiVwiv3E5dsYQplGbvZXQ/pcmf1lOsqW4JyUfRAWTM/Kc8sv4G+6pLqX
1EB6vWavocGjdr3CugLuBJL97OQQxgtIgc93Fb3ZzjdkxEQC/OMsSbQ5n913ivR9
NdVL+W5UAAVb5tSc5AW7JNeXiAkdz5Dga5e+fnMva3GUSuBcgtEsL2tvieh4UH20
MexFWPltUUZsDwK9kL/dQzSS93Eh4aR9vaSiYdz5ek6STRTNvdB5SV8Bd5m+16UF
iVL5azhXvvXVEHnDM19nFAkxNOGuUQMk4/xlas3sIc7iow9pKxlz5eAdNRdxPLah
ILHoBaopIW5ngQoPDl/ztl/PSQxJd2RmEumlWSx1tGGToWHKGfSCkUCNuU68uBqa
s8SDIDqLENQMX6Rx1aL/bByDh9BvEDP3ye99kp7Vh4SqqL5QGdbjoXjbW391t+NF
KZmOuyaP5HIIO+9ttzs4dpksG86G9zT75nQTbazYFobHNK5CL0730LkD7nIgcj4X
VoN7gV4YEUbf9WchJyazH3cCsiRIpJaaGu8tm8eg804azS9VwK3AMw68ZuGKa7VN
a8uwTcMkuB3daLtjtPNwimqa2mFWDyTevwB8K3rHr5pItJc9Rcspa4d74Ne2vLR/
gR8opCZ+FuVXo3N8MAZVRwHC49sDD15t2F0lR6lSYk+Euhj6CCY3OV3E70UWHXrK
c//BMXU1vzPCNjT3N4OmWDQa6dJl9yaDOSiWLxZUZtJBYSyi9I7rmoZycIgBfFFa
lgMSEX7SVBXDMS/sD21D783tEhutobMGhxEnqklIVUgkh+uALIUgS5hfOwtGijH9
amhw7em9PLHXTL5J2O87CHr2LGAv+jjLu3CvVlAKYIgJHXYKYULwAnlSOSV4iBtI
Mh262CAkjvZlfzD23vZ389F2+BojqHC4nE6JHi8KHXAU7z2pD8dsgIfD58ZvMVWJ
8VWBeHGGiTg+RlTK7KyerGGNhhkUdH/c0r+EbLyQgcf08Iqv4mDQCNSvvnoYRi39
f4n19WniC98c5+kGRZeIplEamY+wAGvKk0XmwmFMTlBrdH0LT17wnyBoymOJwN+X
1D1RpmpOox8VWFo9WTDhgfkew3qPfUmPX64h/hOTDgYFS1jjdLPw0pL3m2o3fb2r
bGX2qjSzKtDyUKkJbdkbEZiwKSQzRMcbZVwouYuptT42saTsAnbpOyQy0K+I6x16
Tqtp6aNAOJCfgtldDIKGP2d+txOKmkJuQgFpYTP2F6UjD7PeYXLcTPiGriSojNBD
ANKFWYMthL9OETdFR/1hxfAOWe836vwX5HO6ar2/WIbtazkHsjDSvQN2FY6oPKH5
a65pcw8cPtALj2h++sfqr3fyR/kuwi0RJVMfeUe4qWaGJKOSAD1EaIeft21BzIcF
+ERPEX4GPEtvtzzAL+yIGGUwCGZPkiN9Swwdi24+JqrotC4qOLUp/5sHXaywhRj8
zD2oKOxO2qscXSWpsoX7/5S+rg5JAsBgMT9HHuGsX1dFo6/i50qlCk5vqCeHBmjF
OdeDt6acNjEa4bq76DpuJ5AR8BJGrrzeFFZjHB0aIe9MHMqMk1oC6kZIVDURfU7h
u6tmO8G7szzjtlrjajftsj/U7YS/IlTroE+2QOpKdFLjdOqKk4IWE5HDeHP8cnug
ERSN+SBKU2RGZ/bk9IaekdLZJD3hlvy1fZWn2rpg6GulTkk05R78IroKXdhBB5cb
1As7GSxCQbaSYlXudnvp69wDkLf5ZsmDRrw9t6CEPBw6PvRAPXAKoJ5ak9aZAbw3
r+vvZ5Bs0f12HiBKuW2RTBvXXnU7M59EiosraagsMPpVahsldoqvgdlbkNEqGY5h
6hpOAubvYSHpufUtO+lq++8PHDhjkOLp/ar/hIMNMeysUx8QxGOMb+IKrQDHiAHh
WykotkhSAbw6d8a31CYRe1g6eveKuFCQ9EoU/I0w9tMFomLCbLfhhpGy+rO4E0zG
+mZRtHsm4GzvIT5+2Lf1VBrBM11+6WfvnhoRMp6acG9YvSi8uRlJuz73qQYqrvnv
CLAdaTX/Vabcz+rP2eXuwVoG0WCUEfjZwRTYULOtbB0ONPwVhf1W/d59SPO2FdJL
2fVL8+gRd+2kJDpRPSfLrCVCaseGJwafyL0IRC2fMIfHm89A79Oo0Adp2lThiWbr
yB2dY350Dt7oSs9nQZ0cADjXmhxg+f6bOHmsQmpROegneqyI11Nsagk5IkpiGvdi
1rsH7oT5XW/xmcL6+TN/2HGAmLqJtfQfguWxl5FG+p0fcq+e4yWYolCt0JR/lfnr
SSBf6T1q565NIhULpYvLaFncGFuIsUm1PtLV1phfaDkECKDZfQtHdUkCcHplvJyh
Px6YG5qzHPTJT8XzE81q+r4l5GvTmK61u4LtLxnmCTaXvmxsONelbJYYEOXNWKYN
lJtG6UiqKjMCgz1JmpZcW4gScuAR6utQGLLpqKDUTlfBQq7tf/fvx9o+F9WuRI0v
+RBiSIhtN5QqATHIqRPJbMoHlpCNxEDdTa6xSHSUMGW35KPGyNWQpjppI6v4UrpM
eeDQwyKWILh9VtjHc3lgknRoXpemy2e/9tmAThnR2cE213RkvWGGINj7mIqdes0R
cQO7ud5+2g/nbgosQQe4HQOmrNhUHQ5c2v+PZpWjDXEuHlyvLE7M1qzeaVadY7GS
/9l57cFZ2ydVXXDq/unE0IFiL6EvnI4RmmwFW5DBIUKzCy2JZVIRwWcr0nJ7s1aK
ScDOskicGNadxIA2WNXyEWIjV3qzzLIqLw9W8GC/GhBm84WSKvZDSBu+rFvygDVx
kvUlr791tBnrUczN7njv84PlmcEjNJ/bU7MuzvTQZ0KjC3puu1+3LjyCRxzhcN0B
xlAudl7Rj4FdjQN4waUN3d5dlNgjc0tBHQejb5VOQVnxl1OEcIpeNWDN2KRO/x6m
Gm6zQMb5U7XwAitwgUbZhBY1PkluOV869C9damylSU+b4HWeBIgW72MIbLBn8l6Y
nCIJcNuM0zSXFq2nl5nLtDMTKgO+zbF9T7FJIF83a4b2q8QUS1Szw+mupz78hGvR
8ThrN7DNC8Grimj+lucIk/To+ONULdA+C1hvf3e9acd2K7SExTWnIpdNav0dkrXm
dArOfT0et0/tl2HvMEyP8+d22MdkjjEln5PPLXknBBmkmoD/boT3nuwzRoRQHNbu
hOdzH6Meoay4Qr0kXHbwIMj0Z4B+st9ieOeGZmgaS6S38EOdfqUV2yE2DG0aZLBW
08hRu+3uLbqrI7oaIJzpw+Qj5RIZR5iTyZeKGKw1shF60wex8kCzmKxLxRnyYEmJ
VISy77a+5Py1gTJY2ZONba2Dcgo9dJecu9ZNLRXMDIL0WnLa2bfoMmSVhlvX2+EI
JrpYYd2j9WiIxSQ4dEOd/YOlx5e57rvNWHPwz2Upq/oMi4yve0opuP5x59Y8nqZk
ZmOPUaYVXa2OM5q18f+XEO4ARznIuIaANJdJJE0TqcmbHGcdUmbAgtCLCMgXRdx+
KcfMlq3RC3yebn/yIvo7hjwNi1ihUEele/uk+UklWrvpbMbVck2hon+8DKa0D+8i
GbY02xw546ZqmLDhBcCoOAdhnFSsVlFgjANmoQnxkNWFve+wflQLC4gaA1Db4s61
DYDQ3CQyz3GgUo++gDfrzA8hU+ndxzTocyDTL7ddWEVSfetMoM0NFYmol/inShre
ASoV3L1ZK9HbT7Zlu4ol8htx2OCcLZFAjlAnw2tYKXbHlopuYgH0HMuJ+HPuYeX7
KbCZG6HVs39AICZlch9DZ11lJbaKEMLXZ88UnrKghEGGLxLTyGwuOYVHlDcagYtG
EqT6NLTBFW3yF6WlbL+carxv5xPYlKKcc7+zxrDdjmLrYL/3JBIFFlPmMTKtRnRl
KU/A/cc3aTRIXXT44OsfMP+cieJSgdyatXRGKRpv2nmojxrTNIQqzopHgC/MB/Ef
QZ4U4s+NCbVn7BnCg1vAhgXPemhS4ji2nYQxfQvjyStEYhne3esSzMy9erHJEzfv
xdlxtwuW3dAZYh40X7chPR+zU+Pg5G7GYXIr9Ndg3OLDTKaXsjEgN4LhTQfVW9Ja
d2n6iIDaCbImnJ7i+l5dh6v3SoD0mJWKMdPuPdGS7xCP/fSMIwBbZ5YLk0UFPExK
4LrDVUKKmtYIvj8TR/6qC7yA/WYh7sSvUwbQJ+K3IIcnwCfqJDKoow2e7S1lM8ud
h0Q+BHV7xqeKlU9E6ZYG7d9qjFEtBknvgTNvnv4iF6Wd4H5jdLK+AcxL4I46NQtc
h4gg8rZuzHl+wSMQYfLK2Hp3Nv2tXesaEJz6DwHBlFF/ABCauXTb5ZXV22V7dNvx
gIBFr7ltqLYxjmpT8XNdhHYugHdmlGa5YC0djo0cvPhtdOY6mtlPTmL+fuV4Hh6M
lvfPeA3iKA563bJYp3ZIz06oGjkHeduodXngoUcDf3txsD4CR96NjhHKk4PsZvtl
2UVLDdzrgZa3TrrPbVBd/SiQA4xkTItf8jgKKd9ziaRF4X72VETdIj3IRFu45X5/
2ZA24ZfF5im/tLynvAUw7cPMiJIsTnDWhmHreaup/ftoPTkPYdgG5EXZHU0mTmD4
ry7L5ULsulZZuwCbn9R9w9Y/2yhxDRqcwNhGZP/TJRhJ62tJ0XgBGaaXA63Al84n
GKosatccdwa41/jwF3sf3J+u1mu75n5xb8cn74EjnI67egJDx2N+WcGUoVaHUUYD
dPLurC3AlwrCd+TBJSoHmXejnTzSgIolRtek+SVChMVlgIUk7uhUTrUHblhClAkT
Gn3ONHKfo4u1e//l4mf3US+oXB7Ev6+7YPqYP79W9gjTIxXbLNFwc9FjDPODqc8C
eIXaXlTWB505lxgtM5QJ56G00J/oHFPKV/ZUcK4D8+9mqwZ2pd+LOgEeaL1z0mPl
Xac8kcWrt/iTwpxeP7jZOp9HNMGdtzTdGwOG3NQmBnB7CNXcQHcS7PlrapMfXxeZ
DEVJeaMgaFo4HsQVym643vv2pWfygsRmd0kPlIDdHTTv7bg6qgDjDz2ZEzhbZWR0
JMXSplkLevtD2OvyYjD5bndj5iMmMU33pQR3vQjhrw2tZgNm2PsAsVT8GzFld5rf
R4/J5VM0tK/kvlua03ReDnFmZqgIHbY3dOpVd0qRQflirUlOc43KW0bteB9MOrqy
wrM5KWQx2TZf37pt+kyv29BvThfyw2xYSGgSFRPf4ZVzQOpmF0uU8fH39hsDLQJH
8XpxWV+DAduxor7v/GCDRoqLkfXJhLBMvGE5lp6cn37MxkHQ5ZUj0plo68X8axXz
lRXzBKEXBtHYVH01Gj0TgQGGEejqeL+IUDT5xa4F2K40FOBQF5dhnx6DsZitKX6d
lf+x3/7W5Row1/ApQmShljliLr9xGMaPu/PiNw8Cxz5xvDNYe/++orgoPh4StDw5
b1E+qdRxvyRWVQb7LZEDBf+t+WTpUxugxI37VZH5Wfw053rgjV5pTrdNuI1aTNwM
z1LcBcgxbdbVM7/JhdX1NfyxncmqZZpFsilqvHPsjUHuMxMfPwPE1yIaSf4TuM9L
8ohL23eX9oF/3lWY6wfsypBAajXk571gY00m4fQKRdGNXCMVrU/TijC+korHBPCB
hL3Z5gXa87Uh3jjFsKbtuSm0oVbPYtB1R+b45qsLa41RUcr8YFiHGaut7bI8e3a4
wv3JGc9iMOPQNE2AoxTXR8nHfs4XqOLHN6H6VL/58Pu2Dxva2kaSyZRQaNKuDPA+
oS0M2McmgZDWxZSNxlXjd9FICppQLjCO3G/Z7hCWEu8w71Mv2Qs/sqjZaaYd1m+m
wdoA6Ug4WTuTx97Ce02nsXqm+x1f5QQ5W39PSe/XrviG6xZHbSbBNO/6D4RmTMZF
7RvT4BgS7Jd81JzQW2+xeoNviei+kbIgxeRqzCOjjCq4LewfT7zsFRDp81cWYzxB
pd/HHt5kzmcidUJOhisbb06brXPTugTHvAJOW6DZpPsI/fgwsG+JlOGTcHY6i6Ev
t3fcELh+loItYgA/Naxu3GqLlYlm7doTAg3lJ9zfDMUdu9BwC3MEDBV4sfi6/y84
Z7sV+gkCcYmoyO/SDLVOqb5/0/Q6xAZmMaOxwM7233zUglVq00aZwzOcLAeRQ4Qu
WkV4fof642YfKpcp12YXiEMlhQcqDQukPacegAe95gvYp88aIbpk5f3RRsOMCPzt
8vH/tiqhu2F+zZFYvrcN6ojksuFuGbFCfN4OOLJfewgLxHlN818dTLcgHqwa2agL
dbz6jW6VyRXTCtXaV/gAqp1VyGvafcEeYUCj2MzGNh6LngsIzvtxwjQ3EArRpHs7
9y8sMAG8/qnxKZGxaF5wjb10uXBFHvjkp/EdbxJIJiq0EbLRXMy1XoB1P2IMsQ89
anFN09j8ctDtmw7pJGxTe2cHnro5z4JsL7v7CmrPGUH5hEyaixZF53tHxVrWdtgR
G/OvH1yp/dGhurRGKFglAe5SsIlSednoL8ClBfyibc2Hbg3lJAK4y96WZw+Bx3L9
bE6uARTGHcmIIUvGoDRr+l5ltias0flHM6VFw/hT1KYklp0+T2/JX+5o1VhwwZxc
LG11jnhsf5D4KCQivjarkKvlSFQ9wOykGobxm1EabXBfD3lvxjt4lB3p+n789Srj
wfvJQhJ3KJIvBE+IDgWOn45ZRM3wlECv++sVmTzaCBhtEQ+Jt0UmXByAyfDz+3BT
pq9eQ4MrJRIqm9B/P6GqaKmA9ldgUFG/vqBvEUhvk0ZN5CUQovlyVzI1TEUOgoaG
DM76JkE3x9QmaoUAWwzkzPFR9LHOCJdAhjvYfeqySHK4VlPmjzHGihyrnE0WEPvp
qT0sk1QeMB/hEzrfKzj8N9jhjLvnV7hbqa4OkSJOiryc75vD4A89HJp02XKIwFDw
CizCdv7MQet8SeP2DhnoyxUvBFu7f+Qm6TAdhT0kuwqYyPcagviqROkBOpAlopnY
JxpxNsokIAsLpuM94wsJFlS1E/4mGI1OtzqG4h+NVAe67L1d/sQWKlaPyN3Ql39Z
/X1vdLF3jYWQFvUUiLd4SJoeDlTC+Jtv210t7y7F6rmcLEX9s0cuDJriai9aF8Wi
4AnjPQ19r57EV7A1nIKkRrFtTlWWAWJGcN2df+NmSPWSlAX/LrrQ4thWMBZ24WiX
nOIKt5jUU8K3fvFPGe5lu8W1sNx4h02S3WdfZGttvyohys7nUAF9cLzvPlHM1317
mgiwi5nzCaSJ1wsrDkPdpHsIJg4QBQUiScycdYCcBzbi7WZzqhFRydf7HWR0e9Ot
0dsPMUK8a6iZvtAgHXWmTJBihMrLnSrTwZfln5F1KQesri74A5MiDZK4o66wdm6G
hlQovmZU074uKsr7ugYR1PCbVZXGXGQUavm3Gkyk/JYDQYhwYUsDEc+Iu7lLPy7D
CctS+21H6LKBStuz9X3JbprCQwlxcDOTuuT/+pQM0ZcR3ELpjRTuyhKQOGT33Ote
q/mpLszCzMX+QOKTkRDh03sInjoS3IGQVu3rTPBK2ok/ElzKNRj7gGtjRE/fLIiE
CpnhDM9cZKvkktuiAylbeDLC//d2m+iLw53k7HMG7+nISdiqLPF/LVBdTFW32Hvm
jZOImDwNyxQ2VsdoKtKOcAXZYF/LC5ceh+TrA5/EFRV6Ruy3+1sreeeogp+1BiYA
576gtjJDd9B+etmZR+8jjC9kx/+CbJ6nokkfd5CtFfiAJTN2/dA2WM44C5wBPGwS
3U+2+2PbgyZuRuFPCpFaR6Gr1AHvGCzkfH3d8akGYLLryAVGolNdqp62Te4M2BUx
zx9d1fR4ym4rQ+TeXMfxfXnlMFDlCGQ4WJ3Z43JIOd1hsNoZ9sbAbhmzaLZyDmjU
oM5G1NYLN6HJFQVCP/4cKRX5bD1oMtZkwHdQFiJIii1T+2BIO5VKRJJIfVpWpDjz
j9GsQ4CYP0bkDFC+2/yJQNs0cdTzAAQqRYJ9GJPw7nh6lxLxT2/0fDY4UfHKMDtg
zcgi6Cwcqk1uLiHwvsJthJbNH2Xj3tcSmzCdxawGvNrcxlQgHOxrjzi9lN2j2uv5
DAzbxnpTOqm1tDlb4cn/vKsg8cdnDZBnFISqYSueLvUmyJfUO7XUktmvAFSDgGnU
cuTK3215yXW4UlY+tAoIZwcaGH5O9X6ffobC2aWyoOKw81f6oaV3iKm/hqAb6b3K
LnrxTHoBFyAvfmHgnm9/mPC6xMvpJKZ93/ZoyVUOPcbG4P5OH924/nmQgyM5kcj0
cbFAEDx0N+L/aoMLetSo19Tsq5efO39Ap82k/LtEz1ttWIpDcbheb65lFDN6JnIz
YhMo2KEXiMWASvLXY81wJBsacfbjYBINXYOhidw5ihIvK5MdUXIbolOUqRMIQpUj
fYsi1ChX6GNH+rG/MUhVnt0jWrqhdWYLyw3JlDg6qDTYIlrJzzm7CL+IafXzfuwR
Uj6UdXJIqSQjlBJ6rzBgpc+3kOZk4fraQrhGs8FqqZZ+vQclg1RIUSi3zGzzFGur
VnJax+y+cnUnrB8AfIdyP3siwRf9/RzFPMn+p8quDd8qtyVrlD/mz0iSpeDLuJJw
Uo94+M+zon9L8VdOsWUOuplCayeXE9FMR/uH+OhfEVs0gRBYaczWeknWcbmPH6Ds
ifh0T744sAAT/poerqnv3k1QwO9Q1uXyx+jr9Kzk1EMsbWh4PDpNfwGpraPBweV1
OZ81ZBsTzxkLdCsdE760QE666Dpc9+PCEG3elB60lIdEgiW7p6WtQ3PV6W7HZVAu
BPMgRFbAi/CtoOuq+jrFXHV6nmSWJA/+aexznkokymtOxtQjnTGl0rpbeQKBFGrh
gyQ9fTxKOgElFEe5b1ZO2wTuif2m6mLlWoknEzeabAh1gzdYFA6mOdA7L6i8rsRL
WIjGEl75xswg1HCX3x9LCV3EJJRjYVnRocFhnMZYA2YipViR+j/Un1gNcDFib8q7
dWPGS+ADGMsiVp241XSkrUz/pFhq9Yt4s/GMX+wQjMhDEv56bugvKV/uMM44L5PY
p7ah9QAMpfQwGC/MRBZsExTflM3OPofWQ5k29sEbwe22ahcMk7/vhnfECWdNxg+X
6lqmI8uD1NOQL1e/9TXcw9nG1F2bzx/hPrudlAI6rd21b65OVVfDtbgsU8BI8C78
49+05TLY4ZU8M+c5PLZSmN4dmj4FqWIsJFFcbfbegMJlIMJV7zGPZW/u6u68aoT4
3LP+AQZ2+kjUq4q9FdnViA5cPPdKuv5o7A/+gFMbQ6LG8l6dsXj2Xlr2owZi3MMw
MQuCdiTGzOBL5poNwyyFVT1mGs/a1Hr2iWXkximL38PBAp4Z58Xr+I8Q5t5FHUn1
NHKgiRX7ZB+iPweSxdQ4HD/pAROtGwLul/8jCOzmJNiBlrTB5JE0RpX0UoOO/JqS
DBFGEQ1qbs4nt3XjIFCsiWPdI0Mklv1XcNrME5R6393WhUyIfmBXpqt63/3S85ll
Uxut9r4tl1WAXpxW1O5FHwh7DbBl7r/VVzJUwnRn73sg8ctkjVWtc/Bf/dLMSPBE
hnoUH7h+CCRxgQdl4USf6dnzCaL50T2u28BWLSV6hkTW4LoynlIjI1BHp3IbHk1y
rMNbiqlO2u89cjZn9SWldHdhQUTruenPuyUHMnnkW3LPxbsWqmN+sjn5m3SHXH30
MDJq/QRBBM2akrF/QHAMcU08odm0GxwOlo9gnVSAqCyl2uJUBCoGKadPu9mvuk0B
DeZkt4HpfdD4RkAGOY51oeIkn7nNBys5wi/1+Q+XiNxGsa5ebDYmo1nHXN76ngr2
86J0OyqHreRK4juhQaQcX1XkpzFRVd2OhNP9bfZgtykd5O1lru4z+g4nTF6QaPBO
vkrLJW6elX71J9IJXTIRsM0PmWuRk4sh8BDI36eFjRFKgURtZEjv5e43RiN2CYr0
NGjsYRfSd5v0OeT4M5VLelpsF+wL0JHAatIOJFS9viZJMvYGyMTvuvA//r61uQPD
+0t8ZNnLAehPIBTv6hw1Axw69qRRxz1PYLF2gt2GM6/+b3K3YB2iKEF+VwxxzxA2
NJE/jv3DFfGsHoSQ5RZKt3NLerkLDufcv5+sF/xUyYXB7uuuvzwuBR/jUgZfTFtA
ERbN1Q/k4yJ2FQA0vMUwfIHh1tKnrUsUJRzxfpcw4WkX0PBnEJuX3TluQkSgj9E/
d6tCd48qs00sMInizd6O3b8RurOqNtwv4j7i7uQyLDfIthm8pcx1ub41Jq5SAhP7
MDF7ajCVl++0Y8VTkVwFHvexsPExBgcj4Vk39b8RCJ38q0U9pqxj9AbsF+IZ1s9v
8ayEurdnHvYZPgtqjF9R+IfGkIW+denXBflLCyEJxfuSgRfKVuxBR+1CvSJYrFzo
SgjqYJ5bodDzaHsc1Z61UwxIhxSgKjtu0h0D23+fVqp3aCjF0gsPsCxO/w3hsfnu
sdkx4TIhX/Vzw2AnY9DLlTg33x1oLWoZAZSRe/WwFI/8JL3PeLiZnqXXzexgtODy
UTplKXzg19QfED0PZtAUmBgWABcOr1164uOOv0o+IwewH3nUv9JKc9zR3UQV7fqg
f0PZQXtXlCw7fAhsNLjjv0tXI19kyvRFer7qifq11BV2qVVitDD7GifeoXZGqWhs
iOXBqvjbyXE9EkDEqIy385kt7J0Z/HE9Xf71McRszdAnsSSj/3la6M97FLj/wB71
sz9dEfkWw73TdnMU1MNjiPhCKRtG8/OwEwf+TO5vSMB6tdM50DcWEMkkREkZ6krW
MkgpMOk7Oe7qZS8HGHMVtAybc9t8jmzHLQNf5aHzM61luQ3YFYijUCvbJIC/sZjP
v4tVJuSls4glTk+sQWT/a/gMw2y+q9IxNU8Ggh9KWcUxg9gdViwQ7ta0deDQpuCc
CGNA9yovXrTIX72AcUhEncJQzYvufzE4ApT2iEs1F165pZJ9+O5L/HVS++uIB7wU
RD7v5wHgnYUMKcyiO/PX4Vfa2fb6VcVBeQTQcmaDSZsRM+m2ZawmPoi83QhlmJTb
QWLY/cE+9bfTULsAYpKvL1cNJoPT4YU5HNIHvEixNWzXsZdbV7I5rkVwNvjb7ZNK
ysHX5wcSSycdut8ytp+XZs8fmq9vB8GuS3aKlmFyeApR05JEkmw5/TwaOZ/mJUNQ
woy+9zKtkFB8BSwvB61cmG/9wIIfY7TzIRViuHCzTE+YUNd+QwEFe/XYOlSIdOWp
GKK7XS+3OZzVXkK+bK7YlbSafrspD0CcWqAFoyllCCthj6ryo/biuAMtEngyGEGd
lLyee3XrmNcsTH6TQysd6jkl6zwvxQiXWg6RRx5ll+0vAzWmvaidp6pRMecVbkxv
ZVlcvnMVrBTJybeDYo2N81KCSJcPfSfq7VRChcCTQOTeYGQ4c8HsaIeciUzv33dZ
e+zikWZgs9HjgYrK+7w2MT0n/7grzOHZZnuzhQbRUuN8GhdlWOcfwuhJO3NveIBu
ctBNupI37yvys7pADgIPeu5RT006qqOGhD6QXe/r0G4Sjat26QPtFq4q+FUfKmYn
rWyllPNcJh7Ux38Nkj4dHRT2dSuFarj1MPJ7D8Jct97Eh6bSrESMvZv7jQ8nM+GE
glBLSME00NDiT4r8fDNaN6WRdNsWC5R5mmRN37KlmAS4mSlxSsn8pYSqRVQf/ecT
zTkM8XkkcY+CP+REfxTCaUG77sARWnh9RpMyztEbPPeXjzY93nZyonaxv2BGEJDw
dT7qBMQlimEEUNPq1b65skRnJzBF4Ktb7DhqEWz0Q24VKkm1+StEs77kfheoUJx6
ppBQo4nBCoPo7aiQed2MqrAZ83Nmc9RFQXYdh8uJRvCNspxrlc/u8QvSy61MdKo7
f65dPpiWH1ixL3qjdP2rJnVFNhRtIhINjj0mYXAdLmpyX9+HtIwmT1g/GqK5lK6/
NyezABMDGKiQGZVykk/fb9vk0C+k/KCGSxQZZpLSgtZjidvrIc6Jwuww+3Vtuuc7
h+0GLDa8T3NEh+jLMlkTZjqzliz67jSddB1gPwt5vHRMZ5uIRKri1NM/3ggrTnOu
FSbbcXLZl2QGqm/ealoPCxUZbgRjvDxVR6FKt07TGIgPkBhnpa4RSey16FRrfTTW
5OanQI7+GrVItJy/f1YRAGfrnT2MsShotA+OvvJ0MISB4UgpXbRG5xtCHBVkedbX
nzhM5YabDjhUoRxHwP6/b08vXMJRIOpnQ4m17f1m7+kyBhesGQIy7CN8fSGChIsj
4e4wHJVgWUshNXYmK98axfNp03zB3XyS4qrax+hWT68phMwQUWN6UCrJtgAu0RVP
Hcin6aYHAeRhcxeN6GR6ui4JpqqEVhEp4baaNg9FDHag/Oh4mgfpdv7hHgkCQ2Y4
pnKmCglb6B2ZfmtULMe/uujnLXdbFw/Rcumou3zLtALtGNrgCaCbLBS/sWyjg6kB
IBYfVn6zX2O7QYX42oGWn+Rvg2vUqvmcyN99g0+WzwUUIH4NasMFgOi1OSLslyJz
io29f8bmIEemGF8PAg7qCUUAwFcLlNqFstDCAe/lm4CW1zFOwsMbhVkA2Rj0hZgf
TT0BESR1qbjtq/IyTABSaYVBA2+Nu+WmJlI0rhMrIzK/Rc8YmfUS630z9pthgjX/
OIP1esqtRd2zGfEOfC/4xniv66nqYjCjsxgZWd+1Wbkj5Hj0baOYNsJuusm/z5VS
z0woFxlynEuE1JSFw+ty6JebFaUf9qdeBhQ0Yn/eQrLGJr/g3oe67b+WHBsYxriS
xLGTDQonMGHRGXbk/HdVsmk13Yc7udKKXA0tKCZUMda/sZTrFXxUoXgEjzdDudCK
gNUWUwkmvyq7a8stRjJdnkxZqNl4i8CScF0Uinw8eWiiuG4ocCDo0jvHZrQcrx/s
qxsB+LhwT9IxF/duhIxtgV2S6dDfhXQJnp1vjbpew9QEUdJo+W8NmsPwphSvtGdd
nAHesnzICntgyoM39WL1Uy7nleptyx7XuSXh/ag5VhqyevefNFv56scyFqsf3DdB
jouSVLOccHZFb+juQWbsTny0Zt0s0keYpztIYc64VEYg1w6xX+NbYmF5OUfYPM3G
AhjIOq25Lfi6iz4nYkdZAHl0WrJ6hAjOYDhHE0bx6viqJcJTn0cbsK5lO0KKAeV/
zuW7+p0ClFmQY40yRSGu086Xt8VgYL1/++6GAW/QQedfEobgxRd3KKiTgzue3cYP
ylqiGYoIVAVKWlj0LzVlXsW5BY8KZ3G9lPMIjUD6RsFt2ODIHQ31I0ChGdP7fmV1
j4ZS++EJ/RDcs7V7Y36EtrH82DiQHpDIRiXzMy+RI0uYdUZbPUDKVBTdQDvoQGZZ
z1agq/+0hePwrTm0FwO5EGNekVKlZsL7e7TsE68KqnYeayLKi7vYBta9NOqs4NN5
N7YjQsrz5aY6h14sFbUMdxmEyucE+KP/Nz+E4mBBU1pZ2aTlGNDytic7ot5h7LgJ
X1FrdmKngmrEdtmVXFmruUrNTMTr60I6u4XVuTfvA8w0hwCa9KhC+lVEf3h3qh/j
ibG2Us2pbN6yZBokXtEn4SJFQDHcvAcLmTZYr9h5LV+CdHzNpulWgH6H3ksqsBr9
adjg+of1oUUa9cVSUSDaOfivw8mOSJghQmuQGjyMzA1YIC4sax8cQPF1BQyY0Ry4
v8misADrbnf1hohOYHeyxcvZYjFKa8CrCSlQmeperT5T3X6Q7AosgtAXFIocTk7b
EnvzyxvIJvMaqaUL/u1DSEcXsLTl65H5mfF9jC8NaluirJafa3nWCDeY5WExJOQA
UtmWcyV4jPqEvxUlmxr88u+CI9XBpbVlQxXiuvjubJtFl8A4e2nxwlJTLfOtASez
bcANV8PmqGxJ0TTscEh2d2fKasDsdpcZjtQcv4BQ+tXN3KKDY+naPQx2BtxBg0Ev
BsoRcTZyXhJUHlbDnA3aTg/a0ZeUc739zStYwtdxPmAzPdfa56xZOHAx1rC8H2p7
60+ebmqbPs143FDQxy1UvSHU5MdiWViJLngIj8SXGg/VDJWpDT6lo9NVYf/7NXSh
M2fA/AJHeRutO6HdrunlTml/RIRtd+Rjh52CcLpPnuhQiHdtOfY+9u4oofIGNJ6K
ZylYeiGDHpIjuUe+p4RVCugcs08YapPfhH5x/GRlcIb2Pj0rdr7o40x/XFNRGk+y
rzoGP0MJwbutSpMz0Hk3Ys2CjOTov4ydkxGhaAqNn67lkdVcPWdc2shJRJzIiPRI
FcGZHZFM463WwBc/Phvbc3tMWWtX1tra7pskJLrd/aSUpZEA66mt1sZR+DBHbZCG
tgGhFsG9tRzi3ooWbAFu4LjmRt0D8OdFEUvhy8Ercytee2J8KSGlZJZbg1LQq2/E
wWpyX7toj62u8OH01ocoZ6AEXvz5G0X1DEdu34rnEsjK8ff1yvP6GWiW3Pf10QcH
dUlq/gaI/lQFJPkBT5EGtuSy0+f0m7YWK/PGDi9V3382Gv/VZMjw24sNrrA8PHFg
vycwwwtINkKMLpttMlxPi26EIwbZUhJIloBZTPr2Vi05pl4ezE/QLtLesFjpIluh
sbjLCc/V3AWpTibsUM59I54AVc3NzBMEu3CIFHSSJrotoQ/JS+LsmMO6AJ+omgqM
XVJFLgsgPZAHAJrA02GRMQL8uNehTuuglz5fGEOdACcjHvl9Q90bCAJu/a2FrVyW
U8Arlmuz3kmBJDxMD+JeUBa5rCt8IoRrXKFFYcaZR7E+lDS20tZBr+zSMfZi+y6U
jbzDgfI51+8bPupOhY43gkKwQs72U4tUglC67sIGcPKmw251FW3KeRWAmw6JxT1z
w9DviNY60GinQSGluc045Nz/xGsb4ln8P9R1u7ePoE3hUYHa8g+5RjYHebp1lFB1
rRuMwkJcbznHQtqrZRk2y2Drg7Ptt9elFwSK7A9DjxrnjwsLJ0LiBlSeInofXw/D
s9w9c/mOyJD3mZUMszfWDCy72g7ZPBDi2g4CcOLVjuNyeNzBls4cna9DTUCM5rLg
WXk57pqxgA9hmYRSj7yohemGRhE43fX6DZN/YJi4QzaDHvABQlXa0LKkxUMyGV6I
60TykSu5bwFwlzw066fAtRjpAhtXOyBW0r1mvrr6wlqvqLFXlu6YcKtaBk1bfU1X
fi0DXRFpIGICwQDOii3gI3oF1pQUO6VAagAMi0X+CqpkYeXZ4CuX0rGC46niJxMo
LfEVQ2wE+M5LauVCObX2/jhchpjXBL5nR2CBHeXt6z4Qwe9J3XKsOfalJG8+t/vW
JOXwI+2rBrJq9Vl/3eUSU4UOGkVqYcyCXo9dqz8Whdt1rqK5EJFdF2ebOZBdqOfq
rCj6nD0v6bn6F3f3jLsTgIexqQHlHMi8j43oxgV1O2nOuclHuuiRfckSKy4ocnO7
IOa9ccQYGIIoONcnQ0BYmJXM2KgFu5Xy/MxvceL6MjlbD2UFG4O9mfEdbvBpMNap
n5nyP8t/39wIYUuIY9/WdIifPVPDrV/znyUhy1ShrhWUzZ5tmkn8aEpd2cQivnU9
y30E018XsUCfxmUJxmPycRa9mbu9aVCR1VHsLpAlFyQnsY94VK+66SAj54KPKgYU
hZ9c3lJb6bXoopRsr1F4ayHfofzaiGT/U5lK4AVeaH/ZaIy3Apf47jPbkLKcgh7c
XscI74pPaljr6U6lCHpU4FrxdD+84we+PLXmvHJ21qVy2gKnWrNLHBnAyaLZocdy
wuKsTs32JGz1ZPixXXyP6oa2VQibEtuCk8wfiB27UU+YT9rxekOjk1FJiKBTkY/Z
E3mIT2IlyVrRU6EIpPl1aGmTOR+8oC52yhfDA333sqDX/PgbLewy+iv3S1lujmSL
IoYysc3jA0cL2j23GILB0SPJZmBJHnSaZWeKYRbXzIo5NnQBvZ6is5MLw6C+ET0/
NYQj6MpSYqMWOLqWv4STzs5mC0O4k933GOjfBC3DUoTjCzx3njGW3fyrwJWUtHpY
M11IH/j2Tj0Rr7kVE6+fZvPWBbOPtw1TJbhLgbmxwEkH/wl3rY5dKaRXYNjfAlNO
Efih1wnXETsRB1b/yNITdi/0Dk3alh0Fybbpoxb+CDuYq34ikLPq7MHxVnC2LSgX
WsJFexY9cmZRI7DOQhBd6sIGqUXL+NLbKRySEbGOElY53ytKD2evH4X0/M/Db0K1
1U5v1knBzczirXv0xVl6bMS2gCPGfden9O9b6ut5nMgiKfHIAOhyUGWXQcSxPvTr
oRGVUDbSCPG/YB+WL0pEN3WQEL/oE7lKb7j0/Qaeboj559hxuS/03hkxN3KfNJRQ
8EtrMOr2fT1LxLojpMRaFTQ+uj4muQpTJ2WXNyjkOOkIG+FADIo4lbCEkwy8c7AV
0rgPpsjBlQuX2dzH+Qt2mI5GHYXyoZZW61AxuV+Jj+Vlwq+9rYdKraGDbkrb2R4T
Cy+H3Tuwwp8oI8gta6f59AgJFGlp7/vR9NYFj9z9304g8Difb5/CYaC+Tn+FQEEc
eWcAreXVB/eNRWhE4bkSeMk3HyuCZuzrNyUFg70LeklFgMif9yhydAexTJNeCSut
rg3dKppgLG/ffH8IhRJ10K1ZBj4XgmqTQhX1tLLYhtNoOpfCN0I06kjiDRxQ3g8T
Vp114A+J2IdrKp/Nu7CUt8bo/cusqBT1RLV3711jUwaftNm+2aq0MOl8oM9DGHGY
I03WQf39RJSyh91I/sCxGULCWtFIz+PrizYFfrqwVTuLTW0wHybHQVD2MCC8cwv7
ApwN2tlMPpIZk6WpYmwj/+XAIRzkXRMajNs7k0FuNSZ9lydctH3Ijbk7DNcxLh1t
JATPDFJ9x2zXozZ09vCFkeToH2ZeQV0y49wFltyNOqZTLyh8ohCJm7bxpcvTw7PL
JMz1eSiCIws7sqfUQt6fZqz9T3fPEDWI2ljmRRM7kwDEid4c6nSuIRLaqCGU7+D/
Osqou5MjAshRYADIKDdruluJKzklLW06iJ5UXIQh5S16+qHCAvvDFAMaf4HaQOYE
b7NUUeH36/4RQ3+VEU7z+fCr8MnD7mzdrsXYWeTPkayXCVsY/jbFAD6+u4uc0WUK
6dVcn1Rw8DMs66x5Z9PUYRlVoxdO/jfQa2WjH5031WyIpirZTf43QDq1u+i71OA1
uJ+HxcG8e5LtMDZs+WDa+1ywg/qHAxwwDnN86cysj/lAC4BlJtE4pklhpmPUhivz
Vdtr2fn3r3jqNx8kVO/GKY8wwrVWcYnMpQ4BMEgd91xcwG4QM5fyGUWRPdeSyrpK
P21+TK83PgwOFJ07VQHNaDLTaz/1NDQMS0m9P+qm8ru1Ig+wqv4xdbnHxhGEWSWe
kx6HNhX2xZfValCERoMC4KusnoEgJLBW4ka8CyUyEV8QOy2aWPvTBc/jzgiWI2KX
oM9j3b/1uj3Bx48x49ijpRyVHyY5YK4FSdCvk03K3V+bTQHF8cnX3uUHI5XKo0kr
qZPZvXZnpFKLd/3SMLwDH5qiZtZD54tcg1kJdmqL7xrEqtRNudZvKlNIMml8yurB
PcAo9/OkxDiRrPmAESaHWQjWe6SjfQB4H0XyCd1gT4/AT2hNz61on6GQeOsTpBJE
u6dyohUN5lZdvPiHUpWL7le7WjYCUEdtM/8JbaD9qgbyeZ7B4vIQopVAIzFFt6q7
bnOcKCcn3gZ45KlBy0gkL3p26xrLT4hvq3LswW4d4029R8tN79nN2VS5tyQZWn0A
vMGnZIfb/AKc4OGPFdOLxtoYpNQf7Ppnq3gtCL2V5E+QRrRgKy/46A9QYveDTWNz
guJS2n+IVs4r0yDge1wLDesy/tq50wK7puxhxdn7yHEqGRD2TMScbEQgdhljo5g5
U59Uqt77yop2TzX/6v1nV4UeQ/P+U9HAW8GxB//9JmC/4L9tXxLb23l3Uap8dsCd
Qejefz7Qv9jg7AE6omyqg/Lx7jGVaPG7Pg6yFB9uhnxx0Pq9O/3ERVdNdCgQtFVh
EEgkNe+9sReJgCiPOv+YbD25f0dw7niHEzWJlXQhOufvNKMnMttLt20uOGMVMCze
SvtnA4DVQvSFPDSZ2Z0ltgEFDssHJnH1eQPq5fo1hG75GpNnvbNgCPMtDclQosW0
e9H7aw2cxW/X/2sswKUd2RO0d53SCQLSHshgvcedLEqOseA89OZNF0BVy1g8x6QV
2DPsDrdZQVNZwlLr8k/OxsIBF9t4gjd6/lDvNpJZd/UpB5+Z7LW9pdfne8XlBwFZ
4IY92quE/+wV9+VwhmZ2kQQPk9Awtwgo0XusWgaZO9GhMnY7g4eHW/ZhRGD+sf/L
HXwM0tANM6CoEYSBGkUPYurWq7aO3KVy4ifraDXycJdKGJKvBUoParVUsaLpYzUV
HA15dr4GshLKoNqeqoHDwWhCFREw3EwxDAqK0Z/+Qfe2sFNlzTZAX7SbdmL+vBi3
VeoKlxF9DkPdNzzvEHygJSs030dTGHASR5OSbQL3reLhHFt3lCyC32BIFin2mhtT
9461fUX8iuh9jLTRMvq83su43h6QBZJycAw1khjFxQYDTj+FGiOBe8CO9fbZ7E3Q
J/0UBaGMfv68e9IdpB3TsOfJ5LSb7I4qNp2wnrv3nUDJPKiTeAjz4dnCF+MtqJ9M
8LHkMoLLofwqXa36x1cnwglkxGC9tli98jVrR6kWM3RodKylzVLv+Di4FX9OrdT5
vdBJedfuk7H/TLkjoGSQoBR75FC5KVkpvw9TAdIIy3rmyJwcIrV3P+QJqg9viEw2
rou1Op7BO6ZBWkonwy2h84mWlT1gKLHDwjUUqYEX6L9D+jgJmvDzBnNf69M9KfUj
wVX0qEDLh+AkJzyVOTFWO2xa1IlS45D6Fqry0813ClLGta57tBnlMkmHpUCcH+3f
c9yvIJBVjjS4FJMetsXHSSSeUj7FAdYe+oqYCF/mahv7IvvM/YaEbrhAtVrFiW57
NM3Y7ASR5uaXcajJk850zPy7SKloew8dX7F6hcO9PfFMdM34m1W1bd9U63/jyHCp
Y16wgUrg40z+0iOUjRetFPv5D8Suii8zSA2ABOpcy/W7h6YGH0JG6Ebu8FmlrczU
IsFeByuHsRNtaTPAXoxd2TupC7WOsnesr5fI+/IFqpdUADeNYserowNbVTxa3QsB
H7v85rVuYkUyl6AuLyGKJRiLFN/sfLXb4KAsqjRVdUCwg24nduLajEa8OYMyYdvm
fR0zf9/WL1mOdyRuUBNGWaXr26/0FdpJ3LnftJkY4lfxl6nwShh3QN/8vFu/nIpl
H/ufCXTVRQv+EtFEHvZ+hN5itCtcKnunq5/eJJAXU8DXzwz/1+UE6DOdXN0vyhkj
TLN7uLHvdn59DUMCJfMFNJQyTrIYMBTqpSunmPKg/U/CIarKs/aaemX5toyNmguM
s/zc27iGVMkk8ZaSkdYoLxH0CfVCb41sOGgwT5eDOJQptMxf0BD95xxTx4Zla6LW
V1LM3gqjB1F3kYbCadi0YB2zVsNKy89RVoySWFY6EAPgSevBw9AJ/1x648Z8orzJ
junHXsWbFbbHLTR8fZo+BPDg0SzMb+Tv2x1tYs6HgoDHRK+zKRvh1Vjcmra3IhIN
9qFcWHjDr1JdHXZ8oDQRsp1/XpNztYWrQ8xp6LQI8bqoBfVGNbwqLQFsx13KOO5a
W0JtqtchrtN9OnearmcICW3MCTPv7vrDHRwIZEmd40N3pVpp8/Oal6jNxgZNxUL6
QtNkyhwrhBxtThqWlR0Ge5pDlMJVXGRt206gH6VZYVnGCKEmScuFbYRVNdmNzYDi
EKucEjDNN4sJxqZghrlmTtfHFGxIwCaosl5Pmr62bxZNpbxYTL1tH1yCj+Z9p0QC
xfykP5gcx3GEDjb9cL8ZAJ4FdVaCNGi3rrIl7Mi/OQU=

`pragma protect end_protected
