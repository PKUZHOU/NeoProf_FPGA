// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0jqQwBQPYpKXZBR5SHEDOMjG4+0JSLFbJ+OHmWYUsQW6ixMPR5RJzlaibWv8
2n003fFtq6FP70VEnQZRkp3ERZe+/SH84nGIy/0t3P2gQU8ommFkOnKURddk
7EayOzlEaCLQPFRlp0Zyh27aslSP/PFN2plTYGelgGwwKPw8/3wdaIqfVSeF
g7cLmP8QIIAa/5iNz36tGs0eU0aw2bkL3BhyOjDkoTNFCXDkHyRGRmh7rmQl
lrQ08epH9c0Y7gEnkUA+hlvO4XNjRjlTjfNbzE7/RZ1i1/xqVkvHSa8U1lzD
zko3GM3M7AhwwQ1QG0uLZ5CmZFkfFpdFmzHp0aGoGQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gQ1tDTSQtqfRJXl/lXRV9cVHI89nCt9BYjNsErJIEp5eHhmjqJoEbZfAjb2C
UtLpCFt2+CSU8k1ReYC8YThE1yKoE1oE9hv/Oh2nNiJ7xHUBvrSzELjNFx8i
27IsvborJ/j65Rt6VviWDNOIQAfO80h1xotr3jMT9URN0KJw49rr9RBvcVN6
gWihpQm7IImYUdGpI0A+VgqOa7z4ervrnT29LsR/StGZgzIaehllxCGof2VP
x/yG5sp5cjGQmwT5nmCZrgHFQ3yk6xhp3tSi0ilG7JOIgg1FwGrKkZxxIF6U
CmldnkV9RuhlYeDk7dYkSHYkDMkaqO7vHsBjV5k45g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iXZ1P8QNmOFG/Nar+gHEreRMh1eDZnq4vVAdGm5beU+1ffvZU+9PsVb4yf2Y
x9LqyHhKZyYoCdJtmCs8d8ZexCYoGVCzGZN96CNReXfCBJ8XAWIJYyZDBMBw
HsqxxdU76gGE0sHViQqaBSPTNVAl510kWDWg07SKt2HFma7yoGWwD+ejV9DC
jcHp8VsYGMXdByNabj4WIrO0yyeo4yWwYR2/ySYn5dsSrYFxz/a6v1X1/so6
u62mXPW/2y2XaO54HyRcYeylo6zzHQiI3ZKnCDAXXk0WMqJw5Qa1fUTVXzQE
SVJJPKIhjGnmKKWB90JiA7bOV8lP26kgr1y0Q2oG4w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tG3v9fn+zU1uYOmZP51nkOYmRxPiKZSc0xw00eamalJlPOP/nsqMrUVBve1j
2ZOONJlTBiK5AodtgQJv/gHfW5V5EUUEsLB7+o+RvtIlIjv95U4BB/K42bpb
lxH4iiqnwECNoasMXtTRvrZydBIKfz1BR+X17FDPNfAkXtSYbUA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
El2IuHnIczhmFflVw1iFQPC7L7RzjmdW5fdbixvcgTCOWRfvgwB82icXXmFd
Q3FULJeThc+aQIOUkdgZZsRxJLTPmgDLkBKCpl9nk/927Y1W4fpKNBVG7JTp
BiJIgEdWRtoY4/bB76qbruMUZUwGuN9ZMca8arh2udqJAJPT38xMsq0vMm3E
p2ItO6cFYAyMjQANBfmtvPyxVEPgWKV/MGoD4QF+DkMBYCAC/RNpJJvcPP8E
2HV+9KAd53onwJqhad1OS7Yp8w/+4SLJnyfrls9ovW72iHO503fcXy5HzG62
eE2nr655QLTv/a6oufHkUfJRvyWewQHloId09yTzct0pK9I9Hig/e/3GZEeN
jH651vTWhkYZwWC+0KdK/91AzM6wSOtyS//LdVN2ZlH7W1o6a86Xk4okzEX6
O7QFmtx2i5IfYGNMbjmjv06ZSbe/DgZHdPig6gCVDY9bCScQfv+j/UpsP0H/
4hgq+aLzdjQYzYZ1QTHyC4H3EsBeD/Bt


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ckk3qLXR9GBpnSDh9tvUMMWU8OueF15Kfy3KTPBg4dQZfbfC/G3IcTggyIqv
XOQN6zd5ZoF+ohVK9C6DJberQpQ9z4mlTfkQJKfW+sOW9J89Xu8TYTLShhWX
b04F/Lc6vWFOp09GElQy9Abil37E77DQcqp1KOOI44b24SQowZg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sD9W13E0qQGnI8IBoysfTMQLu2XlZGrw/wwP9OC7KYTyJEnhTBTBbBMg43U5
EbZk7aa/9VFxi0kAmKCKUagxWiny/rkjKHhWuPusgUoIFFIIJlnCfIMf6KHV
hzjTTIXwJ6kt3VAg0BI3Znr/+3NGXkd7QSJGVRR2Day3T3p8q0M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21472)
`pragma protect data_block
zTGtmODr5kTua7i1wb6Nq8Lu/nABtEg3O5skkuC6+VEPyqwZkv7rwKsHVR4Y
oFaHiSrVTKqbhzIzKLtcECJI46ECH2qqHfHtX3tC7IpOfXOY7dhMldBZjs77
XmYNUHOagb+wcqLDn0zS2w14h/42eMc8ll+0QN1JLFXz7ONkNoiZoPLa7G+5
6TchE3wS7UgxMTB/8KAJL2r6n5ZwXgEL8MAhPxWxVg3nvyh09E4L/YE9IOzW
g4QCcM0/vCYV10nJ6qdCMVM4N2Pzaxu29EYcofKCBkxLVqNb2vbOqDarCINk
31/gJ4lpfJLiFXsOG2XQkyUPCzlaLYe+62wQz5rDDoI18jtnKhvyqASK7HSF
mqyHCymxPzvpO5lz55Sn/pbYMHNqijfiIMXAE87a+8Z7zReFccRPQJF2NGOp
hT3nAj5cDYyZtcicTozorTg2/0KHFkYa8vv9xrcHEsErWTTgW6zAwwl3jHWl
5W9J8Atq36N524ZV5kZ3EbteRdeo5X+MAAb7J0+EjWuH2i6ht1ZEdlX9l1/m
d2uAXQZGCaGe90K6aci2dsuTK8a+x3/TA7GsuarqSfC2BLAZsaKwv87PyTaT
sH+fIWT6lBR1HEv14lfgw7mxu/V2WuuDoQ9whgZWXYaAryoBadsNJed3h0jF
ZxUUaRzQ5YVgkBb1dS16cB3YV5JhBNxOWO7eSAdJrR/bMaEB6Ks9XbYZ9p2R
IfUBBbOWPNifPK/Bg4IPdCRJA4ivjEHZbnWfEBjc9I9v+i4CqISXD3T2tBC0
ZJi4t/hRKunJ6bIr1+3oXHfD4B17V5alvmYI9li2mHhU7pXouVzBP6mNqBtw
xdwjdviAki+8L7LRpwx1UQujNm0ChmdZsDcMZSVh6B/XPayCWYugBc2UWt70
bizfWngPsBbVxEZQjIWndm4Kh/ultlXRsXohNH74R3SPtKBPPRliAQE532Oh
kLfdwzugnVdB8Y5+W7bMxlgCpZQeoyTpgHp8nPHvoS9WoyOwhQCR35XX1pkt
x2zQtWLWr6QOyo8Bg7zak6oBwmTbYnBExVTrbGkiRUEOunr2u8K0rbcdQyJq
PwH2DpTAJVkjjKbQ/eDjM03+IeU8OZwgv/FVzr1Xmmnk4V3YNF/Yha5NNo77
LqSnp6LdgKD0UzYTzYGKh0Q4+KqAARXgTsm+oU6sETNAIojQfaKGnGLpXQ1o
bL8/4fhuFnb+uETgic6894Jzl8u8DpYEa4zQFDzqXn07wSnG7lb8xDYUrqjp
sSmj61C9+x79aF/iMkXE0tX4+Y+ZBRpeDYGV3LwlUeojp40HgnIbEY3idFDx
AhH50hFcEGeDvPRjxNyKaWbuEYe1sfQbDPcy4Mf1FvhGSDvyxlTNoVS9K44U
fSNecmcYhvgNxC+acYYtrlL4Lryvh0KDOTDGH4r7Yj3TsUOKFskSHnFIOriy
FIE7kD6VtkIQIQFrImK7rrl5zR2mqEHAM3xgwW7aoL4yE6fFssMg72DJGXKA
rLwTD//oDjxFO7HvS5YDt5YAcyBKdZt4sMh9z+o04wOmyrq8mj5ET2w3t2J9
Rlp8B1TBNJYWvcjzrfZc+LzyvycRTn9ug0ILKrsiPWyndppoBmL0dOmfMZSV
Wdwl6+mwKDiz0p33x/VFmbNd59g22Hv7N0r2c3wXzY4UzjKatMdASXW/pGEw
45ZX0GyoYkow2BEbYZOhvJZG9+PWlW0a9thGi1FZX+Zi8v0Jx9rp8z4sycFy
apIuFZDVqb0C9ozVhE0nLyfPdbL3T6zMOd2uTiMmxpVp6sICgvINTvtLtc89
KwrhPW0TALVkDuxiNFqddJR2JLZpz5U2WbImhh+x5icocm1p//ybfztYrbn5
6mHqs9J+pDXikX1mI1CtVI+g+DPbPvtgYjOliZw03+4/4+m8vKW7tk1h0mqf
nHinFjv62Qq6ngXRcAnNkqIi3uXBsOjtWSkYcONVe4DbuKsS/mE+BeB7TN68
dK6zXyOhznG8jmnocICFiPAWrA8HKOgrsRdxoaV5hbSbtRqUuddwjQegOwmr
Zv6lRSQixHYxD3WJp4AbEthjrIDagpgl4+AezX263ZaR66NUKF+EaK1PfoR6
ZiQGRTLO1fl+xwbvGsc/5RhkE+9rKGhr2cUdqnAj9ZU/vbH8dAcYsAwiFywH
9CyROUnn0mwn+mZzKkHN13SNUNqOxU7+gh4TwHPwerxjgvfGVpigZO12PCiE
8Gk8+ofNDF5ot4Q6aYsIcCE++1d6JQf/tLYDoInS+v5O7ejNp3vjSGnoeIcX
BF1p707+HisjGpDtMp2egDJiFDLzaROt7LxFzZpnN/HXBOY7+Tbv10ZtDgdH
akGPQiRq0jGpDHZjYzxX0SFeoe+fq2B9YIqDEMLmplaT5Xf7lYopFhdSVX8Y
zDe+vdhUb3hNadpt51thUC5SF1RE0ZDeri/OFSZa9grLX8g3EDOJogKFNMd4
88mwAci13KSzrbto1yycYX2PacX2os97cr04IFcofrlh0QsVlGDKGrJAOr0k
KuKIu6GWbk3l/1D1OVAPEEhLxw1K5jvxm/jRzuOMtWUlLEUAcH+/718h8J4K
PrBukpaqTKpVyafN6IrNiu2q5A1+cSHeL1SOsM++EpxJERYx2c7iKZUK/3lt
70dx96Vr+xeOPj7pG9YzEqOuey1mz+tLqB49DQQAwrWxfswyfvkYHYCgCOcj
rmYPrYtuDTDOmluEiggfUDz7WNMCkE9ccHm2XYG+kvkYOl90UNPYbW6A/cP8
7tpZjQ3KtGRKgLHIkgqcsVDPZw0Zui+qR4iIQUL4fv90fTfeDx6KoIf0H4zu
vPzGFfLFGylA/1wdwOi1O9M4bTG2j71YUrHXbe3Gn3QQZYR5iD1UgyjOXcf6
mDTJNeuuC1utVvU9+RtmDpmzWbh2Wtoi4sqSyWlkav+4I+PbuKZ/m3RRJrIC
YeJW/TmHolxgG5sIYV6167Tu96QIKHzVQt2oeMYQQ+wsVAC83JEvEBuhbdS6
GhaOqTK5AHV9LGx4j+QONS7zqv/0Biz5bqpne2EVJXHg+WbQ9aZE5QLoTlzd
xJ/Ow9HN6Xo4cHfEdfuFTTbJXrNaxUKoX4Ho0MNvtMIMesw7EfOouMCzlqlx
lMFaz1te6sQWxmgZ230ocweaaQL3m8r1NPKW3PChYpkWqOakbt4OMo/S6o2t
yjOMdzhH/EQ6U5yAzXNcIOzVoKQ6P8lFBGvr8RmjuyKt9j2mPMTYDz57M0r/
6pp7P0UGF0MEIO5NH1aTbxnjV2KLbYl3PLbP/D4dnWDXsu5gi2DlIez7n/fL
DP2kIK1hLloYz4xzZtirJIRi+S5vS3c+PpgZ+4ivmCqTOougHTlCgRZQh355
GfVOjudYswvoiyauHoSIFlP/9VDL2E4Qj/yXBDxTis6Y4yQSJVvCR2ubspKq
5CclnB6YsINSkhpKlX/p/4nmh1r29qBdQm5jkMmwuCfnZzbfuZh0XBs8RNTQ
KmK2IA7x54exzC8Mcc4flGhhG4c1tihMORDoqmNyhoBQLzUGnhcnNjhlKVPT
HhLKmaye6g3wqUip73KySQZbJBjeDiiHeMeTv/+0+Joqa1RM4jbThWeGGclD
/rkxZHsYkJG3VqblA7FsUNPIPozdVeuiKbMn58Xll74PbjwT+k0PNkHBrZW5
37SBRIAUP3sSpJsJSwF/8VZeDJhhMDuJxJk777DwIC9nB2mrXrmlZ/8bR27U
H7RH2O4smlLL8mmKSVpaDtiaA1eM73U4FtJ6jNJljPqJbbXGygX+qHAayYuY
2fgaFltbBDdbpi+tpaHI4Hrl0GD3/3EE3eMWoZ6w5EIiC1be43ebkWYkwMqg
AYlFi9k3+jaq85vY8cLrnC5xmwHh9M5tJfWECUTU/gwvKrAzHwCPYwkKvIYP
cb5W28L3NC9WYKOHdVJlygbeG+EFg/8cnSeLIvUYnpUPEko5RxWnh7DzZnMS
5JDCl1yGVKQGhTD0Zzxj6lULXQHtFg+kKnQOo/QhBc36HQQFZJbiHnLGUt8R
a+yjScRk+1RfCrlY1ef8FyQ7+qQSziUIKaiR+wrn+Pheni9qDlXBSJtE9xog
QTKJsLLPl7RkFHED4EAstE6o0jr7U0EsYFu5jDpHvI4E92WrOfQR5LWAb1fE
/49tATE3xWp2ldQndCrwKDL9xpSzDM6boFTmiLVBJkyPL/hN5NeT8H1B7jPS
2aW0LRWRVmdRFlfAH+H2MF4LYEV1y2MaSJuskZuxtRtk1HRmynODkzEcbMvN
hqOB2M9kEQzz3cqNSIIgqwnr0cjpy0EswR7X4ZLLY99woYTn9D/F3Nwn8WWT
cRwmZ1LHN2Cn7lYeBvIRu8Uyu/m+G4+JcQ4ufIMCZ6CA4K9Koygz1eKqKSgP
kS/CBkiSoNn2MHBuhMno2a8zL5/Hq+4tb2KF+OryMuw74h6y+7zTVjjiYLn7
FwRDGb8Kto8lOQGvjK5DAIVqv+/+jsIQjKO5p5EfejGF5MyE0W9wCcNsAnay
PBcGK/3bbA/B20krwlWPYOZpQGmFECN7bjQKYK+UdWWGZyYU1D3dxA76xX++
ZdFCcZyqsNoOOZ4m+cSzkex1UfyQUKXYruKjFQlOYWPcj3SnJj2yrb2vIjAw
cqejYPKp6t8jcA5aUw7BDqIRkAtm+UTaROz3i2cFYpBB50vu+wkeuHGeXkrF
2xQV/44MpwakB2dya5p/OY4QEqf9UyJLGiMALn5vWE3jAiovEgedB1+R1NXP
3zUjwUcGTTN7osJ8yNFQeBf7lLEgm7PNCjxAlELNtLMiVKjniaXfz7MjrZjR
RqQk2lgBfVaj/DkPvrMshQGXGMZRoFrDcycuiJTtYzcLSrZEMnIKPdp/1YSi
NrBV9oXsoJ64nAiIp2H3m42rOBmOGn+jQotZkEJQMspfulPsCHKnw4Mv6Bq+
2Utj8FfpstRTTBUsVgpeqgRA5iwQ+LgWR1PZLyRwHPIuLj6QnLwFY5wn28DB
nnuKz41H2qmv+UG7WoILmTK02wNchVJcxG1VKqRcqiDDKTgRwYO1Cvx3ILVz
TR83COW9uBuWgNSudZ2ZADZf2b92ueH3WDV6zIHXOK5MtUW7RnoGkzSmDqkn
seezKJiX+hAhzsoQufWCviAGXLhGsAIz2Ggxt/Oy3AO5DaDU9G1L7BuLJla5
pfgqsIEuzU5frDdjjmHSf4z1RlWoTSQ4PgGzUrnRazexIl4VWnC9h4r/3BlK
Sp8GgcjshHRVAccN6yBtphR9w7muV4X0f5/6Td2UhI8Gb7ZjEiQTMtzwbOeu
xevgNI3ujoDWJFHiPFNzPUIy+5vBzgBuYIY5N5tBm0GclvfOEHVaCLl5NmMV
wZ2rLjeCkgM3Negm7OUI1U8PpAG3ZuAg53kguCx7AQG3PoIVDSKOCH6WcUvw
lc2r2pE8O08uC4eyEjtzMv7Q1BKyqPEOtdWxBsG4KdEY/4oOLqYYIE7rtmc0
LbfsHTE8ksBANZ8JJVk4CXuqg+5oCbTCeoAfEuSSOlFLSQM9xe5hFkhEy9Wz
0+3WEaTcyxvkK0BL4eRRDptOX/DKVPl+tIchTni8fSIt1HYAH5xrEux1UGiA
LlJHe0wu25cXuUms2c5JcdZqayPSsDdldR7EN0bz3VxrpbUMmFsdDJy6l3Kq
lsHDYtGD6IJxLz/TRI0LpE14DXwhLHiRvuVe2/1IkHeGcIu93movu3kvw7LO
DyxK6kzUJLD/kzCC3y/jGmU/NHY2tHDVeVZim4Ch7ZqjXAR1nL/a8k23TRkC
sr4AiuhKOxJEVArlgL9Pw/pKHqivdnasRCqjZd0JOjnxyDHf17+oSMCQc0fp
A+wIfAmbD8Ff5gMu1/7NWD+dw01qoN/OpSdxLXi6yXE3OV6sXTNk1EMbM0Wf
O1/0DEl3FlftQful5BsyuJKUX754//pRyQ3rdjT/WudcHYhAQx7NppGVMvrE
EkLrWuPOX+XMJCKzdenrtGqycctFTCgfbMxikvEiBHqN7VLet+gitgcFq9NG
qvGLuzuoLJh5xdJti+O5h+lonP/NdYXKfTSRPwNbizo4FQv8UmWIdZzo1Q3k
AQ06VFrwqYRy6xzqlbYDY9ljeRUAp055mF+W/PmvtnjGTDlAGAZAEoipi/1/
Klbr2iCm3Mtj86xG6oqKBvvas/dU1hK/6E7k7HSsZ2s2KOx0fPZ2rMYs5gyG
lrtMczxMkcgzGxeTkWyya0DC/RGQeOlmDekDgersx13GErT9GJkT17uBh4Ay
eE9h/dJFR0xcPxtXO0Y9BWOpL+Hg5GlS4ZX2midyy+KcbDFaEGcHoRfR9cfA
wwUjPejGYm3hVx9vd9GnZuY/OvZCfseHtI3lB4Z67R26DrnLd2Z4CN0IMbe8
U3IIZMyL/7hOvsBHzO4iTjgn70JZ+4MWoOvZMtY7Iu6XZ+b8M8L1dP2SklQH
+jIxseDMT8ZeMMRtvkB5oMceGgBjiABhXGZ89sbG0ZY5qwDAXIN0Rs9x7pn/
N1wxlosNJICXkVhQ/wZdS6KAvj8ay0CranPRrYgKvACJNDJg7HYP4ZD7vZDV
faby9WaEKuR6+p3EcCAXf7f48wD6zqO/rWgzrqi73adfQwJDjCokS0RmMzgs
zEOn5Nc4M72Lyb9uzI898CVzf/OiWLgxHK0nquAZWrI0+vDUVb9MvKfU4fv8
4otR4DGpvLPrtX9DcvWKjPYla6SOkRjuv1JFln3S8nhtMBMSPZg2kkD7R4Gp
A8uQGFuKjEj6Gftkf14jeMYR55OWPs1cjqu13k/vywPkkVxF/tBElgsMBgrr
GOHOV6/uqvclWzpYeSuQpEzF1V6G2g1PWawdIVHT/Vy0uMsN9B1iYm2CElKf
wrevNLTZBRBHtmdTAN/PCReYXH2FhciMEIxmAkTMHCBnLLuAtkIZ8I5jlhct
HcheG045mdQIdRsgv+qtgVQTxPuYSHpzDSJhDuUxbwmrELEA4OmZ4aUyUFPA
+ZKU7GXD2xfRFKBjz54scnkifaZQfcxBuVZcUWD3chzxBN4iuvV8gXy4jGlm
4ZCCfcBsu/XUYqwdMYsbzTCCU7XzldbTooKK9lUFM7pwLWev2BaH3Qmm+M28
OElIdVxaOtm8s0GvrD9ANXmrt2UMUim6c483L96ex5GzIRZ7oKkDN6bjvp+c
vy6gRzHkyB8ETMGFYhHDYM3aux3MQe4rnWBML5O4ZshcQ2wVHkyo3T4XNy3n
PrnA6spvHoIACz2bK7rxBEaLhFbR+g/fM4lfgi2ZyK7CPqwpv3wE3Lp4XubO
GucMBnBHbISUY5A3c2dsutb6RTb8PrQ8eYD+ulyuvtRMIEgKEPHQTeFgLOeT
uU4MrqrCF5elAhvAFThLM7crKA9l2EcLYTUQUDWwHnYUwfA+htQbAUZ3nA1t
bBBBosiBhWO7WMNpulVk1DzXy8QPy347j/l6f6o22BEqO48LyGxI4UiXHe5s
RsojTkezQR72fTQUN0je8Zs6qRprbqdT6kMaC/ru1KYRAHZ39LiBe5Zfy0OM
i7+9SCCh72R8sclPQI1pooTphj2MLddz9VGUpd+hFmbRSWlnGtTzcLCHW0Uc
fGWBg5XTv0FyGjpbUNVWoCwG1p6y4Ebs8N0+I2SSAbletNwnIuBcvH4KmfE+
4BRoeX6tEGPf8QhLVK40uzT11+bjvh2uaOWYL6rD1c5AYMgOmQjZMgSRuqZo
x6NJ09j2nGVGIx6+gxtbud2vu6nJvaccNAVcfBNCxxOmJCAlCmm1Tcq7UBAT
OqhhWg6/hOxoyKvO31c90ov20wNqaCY/kDGq/3QMGfcO7jb6N1ZksZp5VwSB
qT3vLlerz59YXrhy5oflpKwJlNP/zsGivE3E1kTRZ0chHFdvJ3qxSH1svxuW
7ZWyE3Yn8CuLIEtr2RDFs6wvs6qmghXRKcQQvBH54Z4Yfm3elZB4gVTB8NmE
/Mwcp2N949a9a1BM/d6dfpb5hcZrityqOe4amWsusIbSsKfX0HK1n30rpeil
yjfF8u1lP8KL/lsGA0Ou2arUYCxiti2eOueDANoNFzsyOExa72t3RMmAHY1n
jgj4BPRG+LFbdQhxuGPI+IYwVhEDyI4SDgmSOtEETYOtRgaoXw7GW4ycSO8p
Qz+nk4AFs2TEyTiCGHGd9xHxbK3+aoHjL8QmKDGBuwLhrp5SEpFJisciSq3T
8o9i9Chk0/YihHjOUcmnx7yYFAydj1Ti5Z5ceT2JtaR3wHIs/ipgTVHm9Yfk
0Skeac931pwj9sE7AoQuHKJ8Q9kaLEq5yE4OuWxLpDxgEs3SKudpVF6XhnZc
V9rYA72xg2xIjVyFBfVP1wmhmz/IztAEImMY1quPQuETVKlxqB3zIwUcvx+d
9RB0ho4sMp4fbFY2EPMINENc6FmoTkzM/5+uv9TBRs1JFuq/6YbFl4/k+HB1
uJLmPIgbgqTvtobP2MxX6euZJvtEfxqgxfzCQ+P5ilrrmzXxhcTXjxDb/lN0
uEu6eUHEasGLlBzPKLnDM2ug/k1hlQC8mVlCIBbfkKDirHDnTj/Vf9VWApji
r4zxWspn8GQylxCFZnH+2ZYiHEQe5xMpueWkQaGXVKMFlsP/QKExeAe0fb21
5pdIFF6KJsUH2g3viGT/005f2lDUWybqH6knxdoUw7JFYLx4hm9Zdv5WKN7E
rtXLOM6sgUJtBH6cr91IQHSpHIHRR17XoSNBT9Lj7hdlFG5t6sJEGreSZ9O6
wtCcuP+y64t5Ic63RGN5YRXz9oMi8Hcu2pYsA+TL0+8vUXcgdy1ADTe0yJwH
3mPS9yJntryet7bUgwDbTEfMqX9FRfnFeylY3Rzc5jfewWrr9L35sCtFDkIs
tfJOCkGJkJVD5zJWBgCIaIYt5Spk4pzNNQxj38oIoyvMnLb1SoQ9y3lPMTZr
CArOc+HkxrWyTqdDJaTbOmEsdfPA3cwTtP/xgHqlvRV0XI3m47Yqhc8RZnJC
Ri/3vll2B7uwmWhIbJuUuYzKC3kigxfVpcfR2bHBT+2zNcD8J3AA19Rrs36O
IysI3iDx5+0hLI+Fz1pvJskxrMcAA8Yl3sCYWlgOayl2QtYmrRByYH41LoHb
CGZjANDqzoZlDufi3rIhqlmkZ5CKABPq//lO8n8EOpDrpWNx+I16F1HqrYsO
z2PguHDYGymwLhk5defl2aonJKaOE8rgA9ByXCJ1d4RZ+N9Sef+Z+42DAEMP
uelzzLbIAUaA0Y+1uy3DDT4H6eqhT0NEu36ez+WeS/PVvzACvFocSfR1P1mX
vujmAWjvlKB/mXsgkVPQ3uOez5YEvc1kc0+/0Tnd37TF0UCg1oUZr8DBelyw
pK7H7hiUb1TqddeIPsLOlJAkMLDpLXn0nXcIrCHlaVRyplXbst9zOBkE4jCS
8Tkp+c2gea2W/dO0tlLXqnraTS0GI1GiJ9ral7gy23I/9LS0mE6tVWynk88j
hFgsJVmC0J90sKLzO1camGhGE6ki7voOPf3fWvXuLQylWTZP/aL4ktsQlfRy
GDEtJhnBucXp3QJDBQY2yWzXdjDBurfQ0RJivSPGOx4rBuPEIne/LrqqjHc9
CNTVVuRZKNo+xNUUVS7lzgnePXnwOMTKPIlLF9PCeEYfALY/eeFNpWgBY4ow
i2fOmWVgdFlikVEMyb74Xg/veEqMd8KRRkDu+DnByh8qumKhJHdkLPh8pPNZ
BWsTFWX8vZjROCMIToZSpEHvrniTndGTqDUqclpKZVLkVC4KN8058Vu3vgFU
F8wUf0X2gUcFXHpgtNc9ynw/QKy2LJ01ntCdq8F89TByg/cwS33jpPLXm5CH
49XnoVX7tlJu7YEH72kvY1Dowk6MF1k7SpIJ8KBumPq6BHlHolYD7DLUtPhL
D9jzoDdBB0efz4IesNMStTb2ACuooBxIvy68zRs5bj5gcmarM1jP0WZbKXdd
z4FEZZ9mlX5kLVQCDdxg5UgRqW+1xzE42OIVx6DjoiDdmsQovcy6RrmGRVop
VkNU7I+dLcQmIRQBlkU+2k/fGfAN3v1HaeYNiZyDNQlsvIMun6kYf9Xk3ut8
OLhfF9e2efG0fKWJWGGX1sQNsC7CYbSQXM4cY1b+ZGP28tpPmQP+JXgZtXOV
oyy6ho+jtgQwVFoWjHfv363vetnrdX7ysaoGZPhc9BdHrSPUg+Y96P7MxEME
AwJhyfzjXnGwxL6ID2TeVy61rDO0yVUvkxGN00MFMOM8kHUtoWVeXnqGxA8H
pTCfaCVbEnxDwZsqS6ObX7KhL/iiUHwZz3JIT4bAX+sBskygm/ACqtmB7osz
ROXfoiNAzORzS2qYxWTbZVtUshx1jCs4ag9O5WWpJFSfdXuqFag12tTWS0F9
pLWV9EE3731Z63alDM8TbBx++Kc+kZ75ST3NkdvAA5gGETZNGiiORe/OK2Cv
h7eYdgNN2rG+hMUExubEunX1WO+8IdBmlxnNIGybj7pn5xPXfBW2aYnYLrwb
O9euZ+FHz2t6J5QQq1aN+Hi5/oFqYrVqZSTWnS1KjxpELhQ4OK0pDp6lQxSy
2DvZjanW+aki2z68bkrXhzZOTOU3B7yu2ivJ+R2X2HgnUTVT0Al7J+ukWg7O
HqFLCq70eZDP/Xqutt9kFJTxGlIySA40lQGImyMSnr4mQ99FzTgJb+KYnPUo
0R4VG8vGVp4KCatgKalGXeJ3Nr4wkEWDLxqY+bi83farfbnP8RcVcPErX3Hz
fmJBUZJCFPkhHDZD8vu4+nKu3TVN1o8/4/QIUGRwA8OiLFsIzgaSKWvJuPhg
QpN+LLWEzrlcc7y+wIBYyplSOr4lMw5K0JUzY1ZCsNcfWutm6knMEBYrA8j4
8TyzWQMafjz64+VS3mZVXWIesj59sBF0lI1JqkjVZhlYrB7hCH6uNlZ/i2hI
dk9Q75BhgPVxxOpDheBZ9GmTZVpPUwbia9ocAeNpTA8QMZpRjG5htEg1LXZE
kGs0ysOqucgLgO4X7EuPRzUEw3Y+YT5zcxAOt31sJB6pvSbfMQMPNuRMa5zu
AQrDUOP8NCtDYWMG9Y2lKiRi+PDmy627N+6Hj7n3UwZEaGmH6F+DUY8/dl5O
ZLw1Sx4vkMwpJJS3Pl2wGWIdBM3egDT1D5fAc2f7o3hJcAPnPvFkl8DxI8UH
g7K1XPcOS36FFkPkVprE/dx/JmVDH9AhM9N+GC1wmwaPUYkgsNT7XIOj5Yp8
/FnvU5Y0avWhMwY6v6PqbEwrNEWcyGvtbF4gY/KkaPjUOIOxPtUft/lv2ERY
5cbzHA3PseQ8EAT9vnKmWBjevXbUyMCoTAw0njLZZM9jmDuY8cMN2lkt1ilg
UztZt333avWNHYbdXVRQUOMTpHd6zSrFS2KyUMIyHyATBbMUykSusHaQe+66
vkyu2Z2VbTst6a+/4bGaLtz8zM3uuqi/b/lFhcKh4X3dj9CEIt2Mxy2k32sH
KxkgvdHN/CTkprRxnNnCCMf+Z9upTgNrD3mqbDe41StovC9ZmBZZLGHSrwJg
tbji8xWkfXCzFrgCtsfojcjCxScpOoR4aKrke2VPKV+/z0CHSsrxpLf+Zklg
9dz5gqv92Sv5FCcJzVel6bqQ36o0ZvhqWtIDarU67YW7tKx6YOXM4YJaZBHy
ggMjfh5cgtlcUgs05GZLuYS//qvqUh22VF2LJJvVaeSf0RNs1kRyN3YCmCie
i5AvDF+dxkTk04J9xKEGtGr0DEpGOstjD4goZ4MRHEf6vZqreeoYIbdoikCY
kVa5JowwQtp7Y2XxfRF8cXsG2rg30zchTK35whU7ucCkbW5i9Yo/EifWYD3N
9J2CuJA6fifmKOT+iwKCr+TxpaQTW59A3n3OHgHQ5RfQLZ/H6MQfOLfnejNb
a6oIl9smcBzvUKpfxjImj9CgwhaKpcGOKtGDHyEGNZhg5OI0hMaQy/9tELCi
oI/wqQBx/a1god6ZJS9c0IN4nY7Q5/SZf0BlH5BhC3RQCiwgDENFBEHOO5UA
jRkiL6j2H+ZzGzbPc3KD75Kh/uuqQO/bB67AG7LYnfgpw9B6EOU9KhK3DQsL
8ZwSvYUCkRBcqTr5d0LblLZ/TBZ6c1/EjV13yIWQW475NuckoGUDgXURKIhw
2SoJUiyCdzrSSlU+UwmFi30Q7cVfJzZWoTZsvan5Ff2/TvZ300xbuOFCosep
MIuqxCIMFOqgUpmXFk6jprKChgsqPnD9i9+nJwz8qr87CoppkWvc0zGZzynC
0TZ/XGVO2AB7fHs6xpDpJcl9yZ8EAAJ6JXF/2OGrxbHwyYILCkhIfeQ1ZgLQ
FawPt4xkAuevdprA6eGDbDR8EfOgJhKlD6kJnsUImonf6z13UfKtvMrmx1Gk
IA/gl+7pkNlR533vAZgW3hcPKWsNp3Ar7jOQej69fYe+ALmsyEacNIsAwskp
46gGNm+Mf7fR0NTk2f4+nCAtZ3VfVizsD80sDATAzqkmubDPha1LtOGZcvC6
jurtzkOIenxtDUhWsvKa/TeFLHq1oeIYVVvvgk+T3pJeegYhELGDrKrNjZiq
gDOT1IJ63Ncr3mLVgNTQ+5vVck0ouEsWfUFZhXxgME4fTguVFV95Dx19Sf0P
S1WfuSPwaHhrV/nEn+6OvXL9G6M+/ubCMZbi+FfTcsigoTiSpxIW8ejpJOqZ
ZMs36ioIonPoZlKP3NkSENsoeQUeacZu+1gs96cd1OU/rM+ZCG3hGOXfUyn3
mbaoT6sH0TpuILm/UF2oZ6MNmItf56KgmIowUrZb2qREIoEmXPkqkzRBXBgt
BqsbyCf6DlGaO3c0fbYtoOVdlG+TEX/DSF5dCxvLeERpViQeQ+MCoRFe0HoN
sU6mPC0Tq1ZJ+B8dqe6DJV5VhN0+81bWvwr7OeuFTDs12/FU5Kok3T+BBYP4
sL+wPpRDEhsNICxRqJnaIsQahXO+eCFXhIG7H/inwGm2+uIF/8ExZT8lWzE0
ZzNxA6xwg8z7J732PJJNYbPWS7gCGg9D5p+1OFPmfnxlE7dpynb3XemDGHPP
UJEOQ9bbC/c2Rewe8v0JQ5D/MxnD6sIMeJa9WHgvjA8048/Gajh+y5vCgB8D
QubZDvnahOmqzit6th4ajfiscKZkSYSxDwQIYL7Z2ZvL2MEB/I+5XItR+2yb
K0C0Fh/Cic02Pb0P4F1sBtXWWvpO5FWcSVE16pksDUvo/EZUaxXK/VgbELxK
thgqYiSgZAt8s7yw9ualTCPNItZjYn3eGFWF05k4Un8sK9hFJHvofpyWp6b6
2B/op3ayIvzeyRbUrX/f5CgiO5RfKnRyoUVZxGJbeX2eiIYKSKdhQ4k5Yaqt
ThzB8ULwVkYz24G0/rsGAuXkLDiOp/DjRemv+61vTXLCcNP6Aytt22kH2J+I
GPvOdSs0eCPQTFQCsmY5eTitk8NP89CpcAP41YTJxrxPvn1USQPnBOdyRCxB
t54R5k2SIWe11Mpr6+KMVLEwoHURQzAar2SHqAiB1VQ4vGq6IO8cN9YhESwT
bHgsGmJq+EXm3PQ2aFgskUSP6Vwxey1oki9LcvogwewG8Fw4f4BMdissmazI
cmY7IPqArsEKc4Eb8B80ASBvbmg8TK3uBzPSc9GBzPwcTlIJDmVIrxpKco6+
UDmMGxsVz4A5ckSfD0X4io6mFfP0LLG8zkvI4X/Ro+lGbQclJlxOWmstDGcj
L30pSCKb19B1Xsc1mLoic1GhVyo0mipbh7A0x6oy6ei+q17ufxiwqQk35MXL
+m8YR0yR+4v8hmVDG1INDqVol20xCTcPoYdWCOOdCry//7QU8Kx6++ALDG8O
RSx8JucmQvD0Pu7tO1OGOW0XNcM4g8nEq88jornvGyCMwmBWEx2pnEYxyAcQ
e2v9AE28OIaKl4hHbqABXPz/a9++pXwS9T9kDpOx4e+MkuuTPwIY5CaGTGpF
0yXZN0kCU+s1shEMpkA8vB0qVSBMVFXrlisbhc8inP8P1hpvCxipMvUaRqBc
VMRkf753lpVf6YvVu0kof4u/XImgF17GueDpqWZgsJv7+G2A7ro+AIhih78F
+c83KSKPYv4GvjbeWi7G7lyZgHtUtu15+8EUA+2DswPMEUdtramx8qkmtKLt
WgQn29sxxVBplUzxPILOYdPkrsw16LJYLxRKi7ms/MUOAfYGx3fiq5umqBmf
vsKERnes/FDaORU8TxCJPfD7wC12ab8rgbt26NlPp7jhQQxasJyKhsH5DqSj
CIu0NIVbyHeM1NXhIiZh7lpbApy1j+RNmXq5rbwOZpeIk0RUKOGU2D6RpPq7
pFsKzBQVtAimInUh0NOQZRUS2OoQSJyWihtezkjg7PAOKuo5ErZLCJJtn7kH
itZAVsqjgZcfdAJZgJChtINSROgFTwg9jVwMCM6MyG8onCvBp+N2XUw2X/wl
vQMZZ0QogG78UV3BUdmocVXMJG1rqmxBCUwpElvBRZe36g3Sj4FYsnt64M6t
IoXAVQCslBwhf6g+YT4Bt4VJvh3M1shBJ7yE8TGmGf+gmc6BLRaJdyo4ZnQw
nxS4SV4TOEzVG8VjHE9D9ixHLIDlFysU8rvvcqOyDTQVmySodhTY9UEz3S/4
HLqldYocWmvgVdBsXpDequaIHsuQDB7SkGHUBi2XdTQHKA8d4GKuSYGk21r1
hWtGawYO06ynkU6zTMMqcmOUB15bWQGYSRtLnMV3rAv6Qwt8LSVTGzY5paKi
BfKPSkYjPbfYpAhhdLihzER0pEHompB6gD0UE1Zl+TRUgREwcYwEXqqs92EP
7RiwT4e1l71bZR9D2CKS2kn6U5UbBTtOmXmy4c6z2pcu5of74CeZZl7XruDt
KuX1JmsC3UE5zsx0U2JZHucHddZR4+4ad8/MwBPMOQpi6UsRrzRbP8205HEH
qqv4bDQ4/AKq7KvWhCuVpUMGFPTB0QvDh2zRWM2RAZCwRHwcAHED9QXpGSSE
c8tkqMyk6uEMsRRgM6kqy4JLjtcBQH5+/6XEKqxMWWNEgKZ1m+hpKV5qfgvK
9Cpf+am3eet+0sMwKOH6PHJziqxJEJRgGuo5Mhj6g+PmKBGOoJqaJ+7hHNYY
KpA3cOf/F8eOxlzVkW4BhTj769BCFw47cb6K35dla8oZCVNIEQIp+3kmOT2y
qUmcm0JswJQTAbM/uAcfGJI3wfI7MFLfn4mGBXQQy9bgXOl5SscGDQx4PEPZ
7b2rBjY79ZY1i9Vh529oX3CKDfE65AO/i2nRUGrBaOJr4j8DiJtvIEkexivg
0PTe3q0fETYLaLCz8ogywEhE9VBFxEzJOuOpgCdhbECIIXo6U0wRWpMDZOBx
dTA/NXK8pfVZvc74kKooQ3EE82V2cZJakHRkJIuo408MKrRxLex9AlMuOseF
gCYTsw6uTRJ3FX0wkMf7gUfmUyPRcu32VgE+e37u6xxNsEFw8RKybrIamwmr
ZgiyRQNrGFOUnrhCHjMvdchS0g5ypBegN4r79VO4s8uLxXWk6Jb/lDOvnRTl
W7IWnJagpH/uKG1HmdysIOSF3wUCHcoRJhUjdwLwMHv12uyFNa7/rRMJe2Dv
Gne41elkvovSdcudetEBzpXZWGNtLWlpAhKiyYMKQ1eun4IcocIdDb+7g3n3
5j4Yv8LlaSqUWiwPGhpfovcjUi0aHVeU3UuQtStRaRAkG25bjy8zsj8s2l4U
IfVtdFYzfxMPsFB96PAhTi4bXj9CmHjFj6qcESW/yaRDdh5HRtaLEgaaKH6m
+PzBq8mlDSLtk8drzkWqzcqAUN1WTplymGfoFN+ZKkOpYJFp9bhxxnF54K/R
wx2NbA5s5cZncZu0QupRlPf9NEWIK1Q06oSDtNvAz7JwrIsVWg9w5r+KTaeB
mTdWxQzB07N359eNOPwnywNQtRfqGzVCvRWSDphqPcWd4QSMt4z8RzLaZTOH
BQ64J55zaJDCTfwMs3hCrtB9KPPqJ14TqIOnwMQCs/xeV+pdzOjtJU2TIqBa
a1BfB9KIFq65NSlhqYM4CRzSW/n5wPHbYFLaOXkpOWjoidw/+5jKGjFfkwQE
v5pRGCUADG2O2w4BlwqMq3OyWFCQtoNl8tXtKSu1L9nf2U33WO0Z5kQP2bcf
dNZr4XMNpQW5sUY0zxJokEJxZYaIle8gWNz/fvTzqhoP0FrR+uyhOecFxwnx
TV8zKe3mVXMPrVDB1eK3gly95u0p0c0oa4HJcHk7m2DOyOh67J5zeKL0+CyE
+bQlOapxY8+L6nhEqVrRaWz99Rqaa2HvmEsKrfOUO2QCODd+N+NQeMaZNI/h
vh6A1WkGcPx/N7Z4lvX38AX/VjU57ZpDjV85DYHhVgavxeSEQS25/lU0pnAf
cegy+wmlVbDL5ztoMbd4eVOanp6zLxDlkRvxhwwkJC34yx3GkSlmOV5bo+DP
1NeHlcVVqVE9rVij5ZGSXoL/P/k+by9uiodw9cag53Qk9mRE5/Dp0pJWz9wD
ztlVVT9Gfxl8aeLriqnlwdV/LvSzCwMQ7vpo2MSPYXMbFZZGtwEJyZPSz1os
+ML97jkxA2SQBZhuWflMQ4Sj6TDwt/nU0bkyEXiC8IOmp5Fv7OC8EC6Vg806
ZYIwHSAH1YOtS6FJ/rfmEkGXp+eRTdZZ9Js+hmXuiAq7eS5nucbzrZRXuzvL
fHS5C6ZauJVngVi2pXQqzp1vdEnfNpA7NTVxpGPMtdFuIc+U1hwiMscwGizn
1Mk8Qs0H02CCfldtiMCh6cL4oqJV0CRIfOnonr7SCsMjr9bzs2hS5j+krlXN
fs7C+K4xziV2rySzUq9YosraSKv3BaEOulqO3PAj83z2bVNcq/Y6n//sk4TQ
n3Z5rDrq4sWTjGeMh9RUkNZ6IcTbPXAPzyt2iZL5l220U+9gR5Bu9U0JiYIh
S26cv6oj/BSR47nm/jBaLfPeSR/iSZOgBdeeTnh8z7KW46Eczyfpq27U7Nsw
VJ9vWJhZlWFBuXGnkAOdrHqpYksjiNIsFXG7iKcTIzp5QougOXGqWYc53uqN
JkdFCMdfOtx/OCmtl8Bcuh2DZTBSayqQJgUCqH1cYdx6hyyD/f0eMWllJnX/
r6DYUy754CrWC5LYA8x61Ee+Rlpvm6Kz7go/+Xxz11mxK8jk368RWG5juuso
WqGkiCQIqogZfxuZU7SqOR9sOXVQMgnZPzzjVvCz3mspnBQkCFIVURxGvhS1
EsUX0XtiIlQ9eJauSIpAynN7Cd/0EvJDuoDDXC850vpIQt6Waxhq8M/bcMRi
AWod1YH2QVrFkDrtFlYfmpcKzlzlXs5NGj2V6l4Vw3G1uzBBZ9H8/zfjMoyl
7pyoqoA6oESlTNhPMwYef0VdEppEUm4bJL+j4Z/hDn9AWGMqM3GRuMch8Zh1
x6AuhzWboiTGBroY21BPl5WQQ5YFHS6VqGeyrDev3V0tFRy27X7DLek8mNsd
z9V9O6R5cyyAOtvDLsMIgXHuv5fQzrq7+z6c12V2rBVRiB6XNvD9d7OE37oP
r1Wlt9cMpEV5OgaxXQ+DyeAb7H07GUhacIxfSlW3wlDnX6VOqxqlRgzDw+XA
bPnznHvS+ptNRJAeKG4uW8JzC3ij2pTrtl3D0HLDoaVALhnvou2i9Kh1jviG
KaHGKdfneu4ERffK62iWV33LuPrLAjUO7LJ1Qw7ehQWoSR6PDEEfv7YJqj2T
bz+OpTsZhASLnUIinAd3+OsOMYFLt6dKYYoSP8AdwkgW6Y/j8xPE6QFj3WXm
XlrhyuaYNYpsOF+7L8VW6Di2F5BXL9WNBCE40sRSWg1vZ393y9sFfATD1gPJ
0rg34eMjl1EeXma4GLZL0iyqgemUICi1fm2nCLYSswqvppS0WyOAUq18a4Cx
djKRVBQyxkSEOxOHwN2Jd/UqFm5jxj1imHKywctffmZE9QqZ+ZXZFfDUdzeM
8NudI0t+rrI0kiN9SD9NRKDNDb60RSpXlieLAUHALijMbsyzjMTALkCp3CbT
1DU+69Jfn1PtJxbJ8yGuBvF6JOVOEvA8RTFuuw19Psu71aOYuVnOei/14DVU
7DsmdlCZVVmt3C6FgTnRp1Kkh/IIW+2zZOfBmHZkosFgeKYAO/KM78kit4NQ
L6n8yllmAH5BV5NYMdxA2UfTfmH4PW1CP/HdqwFpqoXsK176AlBXkcQEDgFf
JO2xPuE4bS7c2FamroWe9qQK3dwdoHR9dB4dB2cX1kWnC0wliT2cn+93cjjD
Z81nNLcEPQrWGU6k9lzq6a/CS0PeF1NdcSsCztm2/w+L1JLKG4wtKb7PD/f4
9/F8v/LTevMVZW9SRlV97ayPKS/lj3NW28k7AM2EiTGj+1mhxzgf2CQuYGLJ
Zpg++wMyLc+SI0Qlk7TOAACV6++Pcz+3ewSBHjFRk5tPNxS531Y1IONMVSlg
H6u9LWcT6+Dm7qxl4uSbEgjjN4oW7rLk0kRE+7fLaVN8JK0JnkENrUZjE7VU
jG6WfbR/zeev3YAJXc7LCxM+GPrkNJsVgpz/q9wIeZrc8aHTOd+C8SCFpYR0
c687HAS+GCrz1yEqbb1jzoYYpxw8bctZPY/UFHl3OzClgwqY1n0aDds5+jEh
qhHpUOFcyb5VhisRxjeXE4IW/pUdiIPTLr5ugGUAk6+yNC+YBan0we8MCiX8
HepO0OB+xpQwxSnJE1aE2zGJ+fm+K6AOeiCyttzlrAqzrNFIbbA3tdwT+GmO
ewurJad1QRd8YChkDkQBPTu2exG2qsUEIjWCjl6P6N5yCnOZNFJ97q8MkTfy
XN1klheQRSz8n3WabYmsAhYMxfUJZ3EWDO7oqjn4QGGzEt9kdo6nLSBrxASQ
kWhUZNkQkSBW3j10aU2gYx2rJyKDWFZ/RywLz6bhwz7bSWWYs6TRmDnEwZy7
mbnTZ3AHYDvp5ymgnOhsW/9J+9zknRyl9qX3Nw5eKwvdRlfVVM9mdqbooVNI
MjRFjAuOu+x69EJUkwaqXlzfqcn3h0nEulzdTsgsz5Osmhkbztvcgeib2tgf
dGUmQaDOxFf+lZugkF5nC5fuYlhciCaHGLEqtKKdn+g3oYCTG85VtAiZcU8h
KWQjT/cpQDDdl0gKep5Z3/UhnCOt0Bob/ve9VBTojb2xO7Oe7L+jTW1IdsZf
evt7Q4kFwfouzVp0U8WYEp7TJLKUzzOBLMpZShDH1Bc3VazfzysMkmkQQj5t
ATfcuy0zE7JifhwSpqAfWSacYPOlHm9qJ6dM4WjVbUVjF2gPArEDLG0GtngC
w5/vdE7hzrgP4Cwm1NHgaqf7jnQZdLfeavIyqhcYc4kJftQPNXXuvfc3D44H
KmGpyZSrTtLemh1ZirW7JYickPAZ3zk4c66kiN+tHotIupDwCoY4Vree+4iy
OVCDFK/CzkIBrLuHhB3dYioL0m6niuaC9sYegfnMpXWcqEd5cUqe2dzO5iBs
6eho+iI8Mqd5H9ZEBhgB26sGhv08uZCvPovV4q0aLDTbAvwif4K8q63pso9z
KWVbZ3g6mn+CZHVmqxuRkLO7xiaA74p2PlczWnvRDCD3zbwg8pVYYmubXiKG
FFqSeboCMG7D9hbufO9SQXDQjk+FUnnItdT6WcOsm81LcvDfMMT/Goz5uIaH
QdGP31vpTIk2VdmMf+qkwHQ2/ftZBtfa6rcQrID10jzI+cxiIamHMkYEMcOl
RsxhPnwjlhITagLH45H0ZeDziI1P8oK/9t5qcZdJ7rvya0ns1Rz4P+S1iHBF
xEIX5SaYPhZEop1g5CPHsvnNUVN/mxp1CtigZjaqqRGQZfOOXTnjjw7sRJwG
28c1fTlzUvUtqCFe7vzXq1ndMnRCKfhxxhBM94rdpqIogeVZO40wDiUitbho
H7A6Y0h/1+EIN/w7OaR0qgLcBHyc3NpVWgdlH3sWlOeGC6Lb2EwVJvUxjzLP
9TLRB0QZvTmyLkMEVeJSm9haMVDlBu+VUA2uUo7LzCeiBBHiGYI+u97yyspI
/E63H7AMipf6Nwi+3tQFamduyF2dFR+axrDRzx4T/M+2UT5jMIKF764oPdoS
gJDD2W7JPsU/bs2rl/lRv+DU1MANAlowNFI+odvpoEnrupSfptmtL6n3E26H
yy/tsZ5ZJekngI47kRGiJ71OkZZZXO9VwaZ2aaXC6MfrUh6byxYEB23v92BG
QdX/D575XXEGQugTMIegZGDm1jwAhzwTppemH6+FPhbqYPVh+BSWvo8j57+y
Xv+9R35TYkmRKQtqcWbopJe5863quPdkSaouWXyOeFIWnpp6n4Y3jjx6tBFI
qv4wE0/RUcHqWuKaXKtHgMEd5ttfNgIJjfrHTtpfkz7f/aBnpfv3G/RtePP9
STRfYBrgzhiJiWlpbivTTM5RJMdTbKUYPOkdqgoH+gWtJ365ZsxYbsaZ0K1u
wyrFFHXunIL9AjbcX8Fe7CD8faQkv3rE2ZX9/qfb+6kwHcLnXsZywcm1wN0o
7zDTi88+C55HC31xkEfIPhVNFFHANSwaHYaDayttZjYjMBy4JcOQrq+aFY4T
BXaKb81EUfGulBL1pc8oDk91S8T2/Wj91TLUVpfc3fxitTv8PrwzCo19cd9g
H+orn2zQN2OOwN4583a6CRAB87QGeYDlOCa5lo+CFHpKsyEKJjP6taXrooT3
el/zjYig8MsMvIodnOZebV/VixwLL6ycZ5LGadVu8LiqhOZ2hcjMtmFLzZI/
lBOZTJ4LYZwDuQ3sY/M4LNCWvhHrVGjuTwarf/XHhhdOiWNIFSt27zk8ZDI1
yg99HtRgKl90OJSC3Hv3S99wnaIVPqxiQKnI3TBp2PV8o3O590bsdveBUC4k
4CFEpzR93jc2QOHrf9mQs8BZAFo+scfUtDeNcXoRDRb9O43P6tcTYlAf+CBg
Kd2iMGMSQ+p7/71jhw6XLg5rO1u9GLnjlgTo+GC8ShpCMXqcNA0Ybwy3kSaf
7MIWZmbvGEvG4fwEl7SsNTVedziav0wHCZ12wwY2kJcZfjeGH1bqIrJLFPls
h79PrDvVF3aLbsRVHZExRktlHCaEM158cg2axcdvZXPKyfHccs05YxJPOZo/
qHR5lEFqlT8BW7I7KcMweRctTLRZxU3zQCI1E5vt99W8o2Ye1qVbq2sMTD69
AAA/zPxZtJrBkLtQFKV1Ah5GFA/WJ/wQFgdY6FKYjmq9wW1+G4tLToNGWr4b
YfDJZDZhtcVVUOe4vGMvTj24o8yaYC1D8zGKNSfMv3I6haTXYyuIFge2mUrs
2qo7w6G815zKGeE9pNIbCm4GJA8WqjaBHcqgTeGNSCC4X4FtzUG1/Zzno8jz
fUXDQ69+LvZ6Lil01MvKvlDUhTEDEv+8qntox4SmVYK72rfgP82/HcqYjADm
k5RMgkvl48sz+M/3wrGD7coq7AdpbyGSyUxqCuFmDnYfvQzyTlIpC4XCsIfx
1HCMG+tGXVvg1qwodjU3u+kKeov04ayXV2H1D8FCjdn/eE66Z8mHzgP4PUSc
1ikYasCsy2AOmvm+1Rq5Z0JF2rX+0/KrzlHMonXVyFl1P4CpbiGUzrFgp1MS
cLj0uF2SXMMW3vICu/ZWZnTreHv8976UTD7zb2ZMJOBIFaqp/APBoMTIopSL
kyuQsO7UB/lW06t9ebuLsKvV2JU8joHidhvMFWAtiSeHCIVMLYcbKNHv4O2F
40zt8AbcoDDNzWUW5q6tXJq/SnGp4MCcvldxBNR/Uyz8ziTzdHdAHvMOecx5
YbvOTNTVOoVQ4iDfMmMs5kL4bH4eAjM8CoHWiP7OJJ6dHuB3DV8cUI8EfZqX
mWoAjO8WuA0ChV5Q2OWNY4ux5mpyC7xpcbSWGTiAN+3EYjqtSxFswZ743fAd
R2pDct8Nw81cbAp0F3NFt9BVPtxC81UD6nk7wqljbCq1aQICheogZvQqYiCX
Ge2tjVvkPiQM7CUh3T350YLF/QD7Jopf9cYm3FsSuL7HYLmJXJ/woY+Kxwks
Z4Tu+vJTXOikARHX2279QopXrHzHKmFL1gDUedReGwe39R4X2n14XW9KX320
3UgfqzUzY4LtMm2kbZ0BDPVslZB0rZ4PZ9waDPVZH0Pya8eM25mAzWz7izJG
sESL0+1jgae7IRhenUJh5GLzGA8G8/Oeqx4ahu6u+IOVb0eQbC9+l3URnBBD
8hiKqMZ6bYav0sBYfWdoHRdn/K3aellLOtHgbNqp0rcNfvk07QfHLjHbRZ46
M3rVydBP4mH61Jpe/w5FbQ8K8vkx7t3aXgSgIXZ9pab8cvi+lw1TWZrGKY2S
LiIDnuclkJktLdApwVG/mmadLWLnAja/PJwriUQWVs6U2m1nw/XOhgaxc6ca
9VPUws8L7kI4BNTq4asK/g2TUP6JdxO5ykwSH+epp5P0HyMNs1dheD5+wJIP
Er1liLM3pi80jCG9roELt8+m9KdaugaHW4ecfrYbq3YTHkjoQl6cJVQT9xtw
/oc9wGeONL8+nKMEVEXPSGJoqRsWLeA79yXvaF1KgitryRp8gm7Hf9HEBo7A
vsdPzEMoa+PxwYd60Iqo9zxD7h2OV9ApjFc8XkDgBvrYN3ksW7gYp0XuDIb7
SHl2hRsWMYaXqMAQozp5Hq1hc25sjvlY6QcRPK/3x7kFqBvut0OZBDFEQs1m
KksWuM7fy5skn+ouMXUEHP6t5fkMhNh30nIcgPtdfU6VsU0dYcRM8HmhqsFb
X/KMBJv6qkxur50VvpvDKYjyJ0nT5af7TkJVk/DQlgvtVK6SOlUJztGeXHXp
z03RzLmyvQcEb60BIASYIxHUitFmQwmfylCCQgMVJaL1po234nty9ViLabNC
wC1LyZsYmRIfD4VgNZ52HH5+qYtWrsxrtiWn2U4C3mergMJ9E1QbdIWQsP18
b1PuTyA6j512VIv9eW65RJL6jkTBMc2tIjiG2JR2/UjoKUlDHoBYi+G1fEuU
5H4HhjcXHsXaxpTjFjjX6+lSMQrJIe542XePkQvb5HrQ4YGfh4h4+rGnppkN
yOnlXEFZESFJtULNELxHksvBC2X8n35HdlvhPr9XJYbYGUVphheOBCP5VC1b
VSnUY6IB1dZ7aXtAhmDV0W/cxQTArs618YDrmArTrXc1sRJLh+RtebYiY0Vx
9H8QhVqmsepXIiDCiogs8+RFHIJGEdtbK6BU1NqZy///1g4nRLTxYJw50Aqc
lQpqUX3VwE6Dg4XyX5SqV4VkJEcyiXWgxQ6eo+UX5WyPUVyUYAlkRy3WmzDm
CbLSekDcqnVMT1HTJzFaBMQbvfJVESBshu/cojA4qwhixzbk/Q5zN7jZIN/3
LxPcCGu3O8cPax9ZqabCV1qAoLh52FrEXs8ixWBAYQofbs1kUzKsMPlYZVtQ
vsPcq4iA36j71h43V144NxsCmMMM3jBGvR6McHVR3R8BQITbbmVvPP6EUEaY
S7+Ty+XICx0SfkcNypRKaVLssauMIcZgTsDwvAp2qY+3bUHSml8M3ihUEemf
WTKvAWiIj9A7OpDqpvdIMeHJnVvcn93wAxK58Dqs1IT5uZE2LoDzq+63i4oK
IcwXo5jyMTXtsM/LcPzurgEGI9kjwL5Bd7D9MBOgC0e8XK8btthtEvd5fNY5
WdposQhZB27Kbkp++P1Pm3KtwagzCTNOcEkgyoyRrKGYhy35NhfagCj+aMsE
rlPw+8f2znuq1K6jigoIGBS1F1zzU+fvZKt+6BXKWTL096gekCxTThl/3gT5
CDebj0dBAdwtvCat1njabk+voQ7lhJMJw2+AJVroSNBc+g42mA0te4RwCQ37
JXkfTgx0Qz2klHInF6TzIAG24ZOliD2ziG9Q67qEdBLpqDlR4p1zBJC41UI2
LcxZ+6UNIkcmaRh+H/snAlRjLPM7O0GA3Z80t/Frn/HRIf515nc3FDbeeFIo
fIGvbaFFFECD6jMx0vCnS0E+WW1DMjSWlilvc4+MDNOCIfsh2w0BC8vLvpV2
cSLQpUuo5TssZBH6lsnRrQ5vJH72P+UE5+9/556PcNYMSaIk3OubYOkCZvYY
HiwkC/Z1sHUvtlR/Vqbzr5aLi44pCKjoz5wRx6womnTHUvetrjBC+LzQfKPf
2JRWWR8V4EaH/tpTgwttkUXKPwfqVCYf33mVTX7PxXKk5ouy1JcsTuvlzVqD
N3YbUCFZPHHsc/Z1465FhZla+RG5g/0bdSNVZNpAGaOQYjfgYdUO6rRZvn3w
aNoDFX5eU2n/tEG9EspOJxIcuAeiQv5BbwmCl1CNTj4IVwMlmoYUyJC8psU4
wAGIMWDZmYAs8+/XfWdNnKReiALubMfylO9ZLcPnVVt2IS4fOnLXLrYwhhQ+
ADBMM4UmKGUvVEo5hin0i1a/X9sK/hhKhbPWN785dRb1llsQNqIYa2j8CIW6
6V7Om1KQOg0Iafe/csScykGPklwHzjvQapaRGxh6efvP23rsMwHui9Yi0b7a
du+aDPLwn0yMst3bcx267SzkpeKTXcL+fkQOBuJHAUlfR98evmGt3ABGS8sy
6uBSwJt1wbYt2CUMgcXq28dyxx0GzbPGqJijwAhwfjrTC6fG1ij4553gaT2w
SS0TysR1WmKNCEhFGicbzvs5QF4Al/21PGhr/IFppuGRTpDwI+th1gKJmkdO
wvjgHodV+bSIVBfQoikxrKNT7XFhXwDhUjXbPdX1/XI+eUYuhKXM/Up5QCdD
okuJaPTM2jxkz2E6G83oEyqeUWtXcB8F5r03ePyC84r+NKKJ+7o7AgwjDSAg
Bm4uGbli47GPF48JJaSQounSKWArxlYHuslPj6lg+uCYFOAMKhiEvxvci1yC
qiZX1GA4IgI0bkdBw3jKD1ERMK2pci+YT9oJn/f93ec4oMqHVOcUEBCS2etI
WI28JcZ07PejukCY7y0vrtAm3kroBwlf8UgANlqRSF4F0/unkSm0Yn11D2/D
dnEsAlmVT7vyaFsocWtMeCRroqOrrocqxQqd+OuiopkvTyqgKXuUcPFfSmIn
hzDYBVeuisVXEcDSBjWEluntsMGJq/wCR6Nc1ACb2rCjQchiNflcm8WiG0xz
Wg0IzL7vG9Y/ra/0Tdh0DRWD+N1wSKnqhfrCJz3w6P8AzyJztpV/N3ZQzbpx
NPvTUZW9tH8E0lKPoq3F5nnc6WOHUayf4tLyxakX2rCqE/NBg89n+Ih6JdH4
8LAuX0u9YBB1q5XgtZNbZdnn9cPFpC9QLHYGsi2eeHWU/uS1YQP9+SGmtxix
GgFu7ezTgvihlAwU044rot5EFB7n8QrA+hzHOq+Tys05iGH+HTuSvxC1Ct5+
yqYG3YVuKJ6Z2v+3ZaS6R93Es1gh3wLYn6IXX/cQP/CDcwdLenGwoUT1GJOE
PLCavNMTEYrvEw5G3D9PH1ua3D+cNv97ujyXv6roYUb9mpJDOWvLMMKQwiu5
d1pGxu9QWJSH5NE3VTDTI+NXfIMtfm5kEtdzyStIKsqy+5yIg7dI7fAJ6kK9
qUdZ1JA2H9jmMsloqQ5s5DlLJGI+gxXSAmxdIFnC5NClbcUSgvWmEPkRxtGz
m3hdLtGcbux2sPbWdrpo6UpNTR9flsbsX9sKSnm/hfnZqoPnTkXwXPHpWsWf
bkmaAHeL51wZ27Nm6CZ2TlkKdklhmWRSlcVb0tFsMdnWOtss+uUeHlJnSM81
f/5/0tKpPEGAIZGT8JTkqglcykYX7SwZRkC394EypmbVBk7dFc9mzoDc4MSE
yLRbcD8IEeO+wJ3qbgBzX46QsW6q/tIvWVBuzZh3om/Z80Xdm6T/k2pT2PyI
XBpWou2ZADiA2pvsRUpFNj9+uytLOo2DjVwLBpC8AFsBr8oQ5wQZThFJp+cI
Bx6d+onGR3AAeva9axKSiJnAifXyIpcdXe7a/XZgNhPCVCZ8pXuomUL/WqpL
/Xcz78mexRKB2g5L1pY4CoTMJCLAH2NFh128qRRLmTKO1LoDzFYF/5hUg3be
KUbr+zlD8M94g3OqMADH1hUzShYqYtWTtHD+KawQTaGENZIOPn6NdRqkg02p
hzJPrALW6bhYnrhMDK3eqUAfwoiu+5n29pzV1MhtzYx/XYNtt2HXbtJfpvWJ
cewftOvrzclDrouB1FSse7JO7jdWAwqp7YamA44fbFcrtum03voQaGhGKFQo
JhhTiIr0nqfh5hTxQ7DZHe6cWVYbwBnyYbDbb9U4ELfWl5xa5hX/BP+KX6Gg
HvqeS6FiE01l829AwqE/Zrprqtrifs0t99ZQvLcYqwls85azsCfrSJloeD8t
nHZmL+7oBR9/jNcKXYeIg8/myTPDOcmNMQeyg0+58QqQlMuWX6v3U2tiLCt1
y00jdGPLVbfs6yB0LP0asd9Rr5W8rMQuBqIwtc6mRA7oS/cSqVc6CQ2CcW6E
Wp9G5JEp/x9hPmbXQS318BImiSO9MRX02wZOQTUUH/JHAOE8KYRjOlhC2xR0
kvtjFkOR4NPMv1VimWvSbFDYSC2R8tO1q/GV4qMYsLN0sM5x0YlYpbg1hCyF
b6CcwuVVFUfJiVvumDyieNMmW45ALVcDxKneonyaXSJTEA22/p9No14cgt+7
tS8Uck0l5QXn2tILqBaOTxOmPpI/qDodLY6uQwZjyPjSEq35EIcc81C4Hfed
qwSsKLZPjcS2lUb3ywiGVMEZmtK5utTYqNBTycF19tJckzUpmGMajN2qK0oa
onjyh/cex067IDJRSV7jt4YsRPqV564XfdMMkl5/uDwLFYdd45wKmTuZjX2C
M85tPYKkSuPeCjRTNfehcb0uFxiOgju36vXHngBeL0MOQvg7/d7x4YxvJHW9
hmBZQjq4CQyDdEjogmnLQZFOUTl6oUswlbIueYU+lZ63gNv1Ydc6I9O1R4sq
l+zMUK3fjkhZUULXI7T0b+wQhgkkYUZ26vpfX93miqOLHJ5yVI2HbKgjTnuV
2FrGlgEE0jnxuAuPil/RWq11loXCCUiPbD82l7vHJhW0i0sh8wbEPG1U+HSd
cR5W+C3dOL1b61NdoBmjU9v8YgzYCI9wqr5dHnn02uyg9QGrZ8Kaflh4Of9j
8W6a7yFzmPRBRtfIYxyCktiBk2xRx7vzh0KFbX/IoxkFQO7zvxsdeNsqS0HW
swJZiXxtlo9iPPFG6re0rSG1gEFnoVkwi77XXiq8Cpqiz547SJsCTEv+CrAw
7wJJvoESIfz1fU2cYIfNVb2hU0Q0pynhx4HhepDDU01lGxQ5zJ/31qspUyLV
JA332w95d1rD4gl4JqapEy/c/Eo5Vn6kTcBNsSTEHdA0GI2rM2mMnhBCNpPS
lXLsCMp5BQ44SL/kmh20aYw5GHKm9u/52oS2gRsuKVl5YbeOOH2N0gDfmhQ2
iigyqsjD4+q3tE9yIIrm5OKmcqbv2m0uJkjgkfEXsgrvTNc7bEmwOWMhFmiV
Wku/zX39MCfP+H61nYqLKlqfV/ICVQm+0+VZg8v0jWDQABdZ4fdxIYLvSVhg
2AHh7Cx8Hd8OAY6/8Yrbx/JHPXsD0OGRSgMbfMZf2o5jKQ6j4W0mz/z155dd
kRxi3VGC2/DoiLISNa6m9kV8KWfOOTJmfk6TZjcoebaa9mywx1Eb8oSrY80i
4d2mS+KaEYtT5yphZ1qbxTIyctjIOLN8iElSrqwJb66TBkNJZBehvzov0zQN
yOXvK46DETddj1iaHQ1/+5NVvNV4RbYJJYgl8+nig/ZwdQTYSvWE6ueipNCh
eWkQ7BEcwkTIA3CqQqcJOMLlWycg4r3zIJyQirEKWon34uI7/iduN0ZURf5r
uAifUloO3OLTCVe5ZJ6cndbh/k/uOVMvl0TExRhP5Oy1ZCX6ZQl4XoF5Furt
43COkobNgwY3d8uDvNIusY5zfqPdDJydK+4gHyCCEQh8TNOc8w9Z3lrpzCl+
D5L+eHt22o6ltqnDjP6+JqY2AY0v6XzyHEh/5QIamYgcD+IDoAmCYMhA1Muv
bAHi489SNSangx91CSCUpTvcjBLOlaSjtz+31Zy7iczEq0/LxgD27EtzJJb2
4rq7b7RTnvMG+S/XVJUJ3XZLf/xuGTMUyjAPqFQTAAajkyzzD668HfO19i23
yPG8/+JJCCldNIWf5OcC9Xku1ssEagxOWhDnC6dg+T8Qxvsm9xXERsKEi6XB
KiZOOyY54BD8bpfsru/QPaUpICkH3sIQuy0nDckPgAyZn4zD/w9HKBcpyJXM
ICbK7ABTQkV/atAj/xBPvkYZhF8TQJrcrWRTlj0Y+vgK8484D1DxH0FTZfS2
GHj4UpirJORHP0/JJoxsr63m8YMdeKE94mnzLfeetekOlZMFAxZuHB0D6X30
bEzctvDCQ3KN/EfAdAWlvGEd8qP4uUurDmmmsN87AUzD+CfPTssVsaYxR9lt
axb0NccnpeuDtOEJJFZyHtpPbhkvrqtkZPd5AjoDs2lJFtbeW11pbJDcazEN
L799pjhVv3h1PmYKWQC4mfP6PoyrnlxU3wXORMWdA+RznWA+rwn68YZuU+/Q
KDGRbuWgtAB6g2UdO0YCzHVYCaL1TtwSlm+hUSiEkFzDgr2k69pY/8Lg8KfH
nE/gaLMramKGVnfsFZEi1kyYAB2IP9Th9y0uBGszH4WCVHGM0GqvqPDikPWQ
YBO+F9CJUvlFfEnZ5yrllrfBwQwHt0Hy1hFjGb1OHu+dcHXx+u6dV0JcusJy
8Asd8I+u6AW80TPiRer3+pAAHP9W9sNv/1a7ZlBSzc1SGNpVVhh1hsY9xW4l
pPw9BkUWxusGLu6E7swVD5ZpyYB+OEmtSmhd+MCmGvRrtPf+w36Ssfl1vwkD
m65BO+dV4w==

`pragma protect end_protected
