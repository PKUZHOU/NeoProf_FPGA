// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
kQJFIO6thg6CqXoKt6fejq6z/LuaRbj4gtcyADs9IEgfGQcMVf3MaHLSnv5DulYg
YZepaoPYkVNFwpMq1c76RBG5GdBWSJ/kDRlDZAKMHusYKBMMf6odfjs97ge8X9s0
Sc2diUPcDns8fPBgsGAhXfaD520ujQz6KQHtXl8K5cs=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10576 )
`pragma protect data_block
VNsM1alYiKkHnZCREBRItMSchdyh4YwwghkWii5RdjIu/3R7K7Sin1qRuNaYDHbl
CTgyg87LXecTZabp5o9JVm1bKl0zwdKVHCpFS/Qp6kz04+RlkU8lPEDbqXOmBEgT
0RKU3C/bwbDd2LWqfcPExY3xtjOcxlZh3wxJ3I9Oy0PY+QXIPmDIjNauSoNR0WHx
O7SLJ5QWe/2nbtavtodDMfDfjOM6EIPCkkrofRAgH5+szPfCzggMoVDqd4vhxYcJ
jkj+6wmAkkfNC9cmzHigV/89G8ohW7fG4QpCn4SkwgR00CIDTWBRLZYpUayitpa6
h/YCY/5VUy0W+NO4XIhmb6NphGjqy3+ARslq7bZi61ygTCuir9fbh63D6ra9m1L/
oxAiyeaonTghpHd69WnJEIgjOJv3pmdv8trcGfdoCYv4ZPfRCo1Rl6RioH/Tw51G
CJn74+JYSffS06oMSCFyGOA92n7OFKdSBKfCIRWndXEJwWq/EwU5hDflCc0KLoxz
ZiT8jGbfzepqgQgOrcCE0k9fC6EBQ68UtyXJKVCQBZrD8yClKuMsZwyMwrgP6AeW
fEDuxlCC8vwX3JacmhVXOYKtc8oljEUBGipp0LvGNppjAFnwwmo8on6tWmDYK8ML
p1koKwRxT/OazlPFYm5gsQ4Mbc2Aqkv0HSY5x42X4a+RMGmVy8TjKHlizUmRUkEQ
w4+SrD4XQIbtfOv9XaNBs053EXqb8SxBYtxnnOTFlnq0SRthzBsoA5TKUTUVNh3D
YNq9tkFxmmnn5+NmonvBtDDTJhij2ioYZRvLVtsCy+NZ+AdDDkLg2xTR8FW5ahrW
Q0Ve6Xe4WToStTqs5CpmB5XsA9e3BKygljfIaS+3zmPKhDV3vvlN11id8bxAoPct
KDLQ+RbMVcBGNl/SYECRZpxSTcbBTGXQROGZKtn/+w7o4NGXRGCuiK8bJY0BNTWO
kukb7XLkWZ+ocJbVjDNQAqWMjJ25burPv9ILhh5tJbSsnH178DlPFyEvVqZe3+od
26lXIZWICsqLXIgzp6P+y3gfZU6POe4uYhUbZs3lKrjkYFjnxR5UQV6u17qhJbmj
bUNH6+QXEsT1aGhVzkoehkEgn1WmCsibheMxxuhugXT2q2JMKWZazCp8xr/bz0dJ
mdls1zganRld0BFEgC5SX7yQW2HcYA1j5Qcom4cPICvh9mDu9eiafxrb5AHAg/wd
OpB0/dDJUEdOnvh7MhavXKHWrHFyZ38zhlBXHSm7vwjUYOKD05Fy3YWfTj7TyLVU
06uIsu47k4Umm0wn3Dn/EXgrZPWW59v9/LV3sEr+KB7ZXaBrQiSTkwIYCOfBWwgO
hal2FQwRVpHukSTHSm/krxH53l2hYdzkFZZF3/mWEAgTigS1zqcakAPWTYd9No7N
ICYFCWP0i+x7O7pd1PP0ezrP6cQ30xITguGuP8RwsxnTUdANVDN2+6DYtuZJoy4Y
XzZHP1wNMICgEHKDTi6+vshGJ3Krn+D8kNpHb/uFxQxoUVtIUzh+6LlGzgO3XW7S
uoPA3FrM284tLpS8n5vcwXEVHod3BtG2VS6VvGsYQI7v7g4vd3x64kZ+HfTjDT4W
avEyhw7NNq4rWgbQKndOPZ4N/ZxfwboZbWVw6lW1XzP7R8QKzYFaCt4Inob2V2ul
57brsmpno5ZF59EDp7lzyNdyQLPc/qLA3ZbE/SZsmAx3OmCg2ElR7mMlVgzr60B3
gF4nqW7Q//13tfqZHWq5ZA3lfb9C6VWzCl/IMf8p4iCLmXx73u+l/E1jFhlM5D7t
6nMKDggOueAcYTE0jUb4G2Yc3flbwhkpxBmu7R1JRE7LtEqvgZ6YV3qMePyHy8Le
+Y7ec0RSeCJJBRq0BasbnrEqt1raLB98kwB+G3Nuxm23ikupFaNJPNWk3SBvOnqg
CW3wv99YFgT9Qdw1xUX48iuvANiel7PhsYSkIKM2q+oDuIfKxWDcepGqK/Cj5LlT
Sr/sikpm7Dqu33M1JDVtiINcCNw/z/J/pWwuqfYCociRvolXuNCAvZPUb/PbVzZo
k2N91FBTQ9AUAOsIHJS3jX8hUQVSKEmhJPNSteWKx6NYQfQy/y0bnggwkDylvEpe
uJwSbDwLi/ZEzT+OjpdA7WZNdgnt4Nrzh1bAKUivG+eogAhR94hjzD56XV+yVQo2
CCRtdm4Qebp6ML+USXP58YsQtV7YgIo0d3qgFG3AvqbncsApEp1Zpr6svt/zAH/Z
Lg+5POxKBOkYKn48SncBnUGBeMKuPq9pcbMPbCoB39zpDN7PHxBtyPu1rTVjbUX0
62H+D3raliG+Y93CsBVYchLhwc6v1hvV5fomDi44fn4/nhxP+xo5egTh/FjlDKW7
STd918C9mrEQNu+qJmsC/rkL4q0VJN8vK45MA0jeXoleTDZTTEE9UoAsLh3s+oIi
iBJGsGftGAxxHzOE/p+JhJOKXTKSC3IOHG2PTEUoiYC4geUaPRvllonsovGCNnIn
oy6MdbFPCr135Igw58FB8p34gotpRTUMuX2nouWrkr6e+pcELyODvqPYFmGQ66V7
OsZnbTAaD1jzVqOIOg/F01Gorf+sDJw4m+UcWDlNPj/cD9M4LKFr2yOsHwn7tvL8
e6SzW00ZteGWuNuZX4qzCuvqEL5vH7H4/sNLpcuvZurmIOzus3jLTMJ69XTnm1C6
C760MGt/80TSC27TD74zTgDp6T2hJrT3GKIQy/NcWoVZB2upYRgcXoUvPFweP1/f
iW6NeJQ885hptHOumMuoy7mEhSUIxxlr2JLN1m4NjqqVuaoi9MNQBPgaLc/yjSCN
ad+xtvtZrpF/5hjdI9mx0ulCKC1dOPJg+Rl0IGWXqr8LQtnl7Ek720lKM2wQOfLg
N6ctwdfQPmInsa1Nc3CZY6XY2hVFM6F7l+rsWSEFe9b3U+ADdcSEPpHOUaDCYNVh
rOEFMwvPbnFWTOR636AIY5zGuj6uWzp8s5hPVAg3uKs1nn4n5B8NOwbRDvqM/Mv/
cJW4NNv348r/53f10673g1DvvPZVnQsZhBxUIwa6CfOwMnfMAm0IYSHF2plDzTeS
9h1Hy5VTbnVLEZbZI32E0Pq5t+UEAyIdwa+XQAculddh9r9khQUNLgcLDlSjGPxF
LN2iebzoNoz3aFCVocF+ilIaJUzdfRSyqFtm8IWUtmvBJ7G2x4oPpBAaM6YEYnsE
njV6Vm4dzoViwI9FauJtjmae4WcSAHsyMxw/1GsOXJRExVSM3fBRBqb53GfORi3k
p81/S+iVoVSIdlyKq1rs6nwGo3aPc9zh6KHs8UvWcLgcsM1TMFFdOkw6FsAD3xLX
Jpw4QNdySyLm+XZ5CAK6CckbZF+96KF0d+QmTzK2XRA2Nug7WV52W5/apmPMg6an
9pnjTqKYg678YEQZrVvs1RhsHmHzhKq+EC9CjbMAf7hkW5xP+HhUqH8R9bwpIadw
RFP2Bed4/FPAtQ0cdknmTdsdfnILt5i1M7/GAOO5jPBula0eMlcofL/vvnq0mUYR
Ap2CvHDRugO9L23YiByddkodICNIu74lpXg7tNSlHPH4RUTVtlwVTL8191jeSDDS
wSPQTJn95YxpS1lu4+sK4fotL30P7Pj61XOBRgh1uVnlYRh0Ar1JbWrmGbQUQMr8
BDXdVBwGkgAYlL1jMLFu5szlU5FA8Exs311ulI60tEI+L98MKQ8R4/3c4Q/UxkOT
A4iSRLZx6EwUsJi44elqJOxazvQfEjnRquA1NRHksbG236hHFIsmNq3s/vIfHVof
Telrfzxvwu3odKXFCyGdd/zRjSz69Yp1SLz+iAkcK8Bi5mRgo4AhjwBBWLg3DPkX
1YrTdIN2wAkKtWHMr697/0wx8RDQJl0nkfKXxL9MipXoR+A9y6ItNTZdf8KCtk2T
wwaFS8ERCxLip7EFgmdNVml92ccJ8dAfpc3Xui5drBds5KK6JklpT+MFo4MpMhAp
RLSAZq+dp4RzOtnwlZzoKCdS54B3WrYTU752U+e2oHppn4n84ilYa1WFh7DzU2SW
m4yTrADpUVxMMXH5ue5cp8I+sqd+4Wh0Zg+DuMLdAxeCDsir3WSUgxO5HLrhhBF7
b41ck2kYKxxmq2oyLyL0EOZt2mpSnLv1Di7HR863LNqNbZs0R1frrysssKAptvDC
oXRDPBNtyJ2eX2iPjfCvTgn4eM6tdphx5AG4GLQtTLyeymF5Tap6mv0BCeM3BID1
MP+ehlYYMrYZf3xqZDpa6iL1QUS5lYYFNPJYo/m8duznFtmzyJzXicY0RISFbj9w
IzDpzY1bNgBv8Lz/+Fx1TTrRRcEgVbY8Zr4s+KFC/UuP3bGDbTnLhh+Hg/oTdqUQ
JrmilKeUzA2Dr70SOTNgs58pywRSsr3/s4TNol61xcIuinMUSALMrotMwyN6j7cr
nVbOh/OeLtiao3YaDEsMkwudOmzLjUUyGvvQGSa5J/o4/2OnPwT8UsTXcuPePiLf
8yIOiKLrtVcP6QHZC0Hj8be1lzhGludmhxq3RdrJqeYTn7Se85BSVjAE3mLyHRt6
7t1EqnDGBQTyNAenYhsO/mT+ovp2nOqSQpw6e5tdlZs+2y8tDQcg7/iJf9t/k1nm
WmbuS6pTmNCe62OL8oEHrz6tRc2JgRJyMVUagGGXYnL/GQdfTUItMOn/eAFMtqeY
aGDdEADoy6lOLmKZqw7a7BSk8fpImVlWq5Y0R4w4b7b7cwLVD50oqjmQKTBDO3QB
+b1lkXk2oGnS8OcZnT68qiC0pJR9gwJybMfrxtcWVaAWnrCHawlRBAhAdN6S5toI
vTc1FS/xPLGMlddn6Ln4PUNJZCoQob44UCD0e01ObokLXkfOFeDQ2dgLRuEb7jKu
V+FLK1wr3/0ISstwlnnohah1+tGMgL+LEegZ+aP+MjHhqRQJLCPOF6Osg765f/wS
IrFqSTkcfUoC7mhC8A4Ps8s2Bg6UWr8LSMJ3INt3mGDas5pVQvw81je8MunoCX3C
UIEIOSWOrSCpuTwNPqg5AWxGiE8ge7JdJaZ+29A91WwTgEH1mNDbH4WUTGWljgmz
YQloAkb/nmJWTQIrtfgzmoeMs9jPut//70YaQeFuN8ckxQ1MgxWmXM+A+FftOw4e
hHtVrUftuCFrejeh5+P6O6EVV8wNJYhIGrLqGg/voRaQEpeJ2lZs3pmQualRrfLw
0PsUfLVvOC/G36rGAnmU7YWzx/VX1lFXGJyz6VCeLF/Ua9SULB1nOXhZ/J9Ul85O
CPT32/Er3FER7xgcqjTr+tzcxfIPPd0fIF1YX6bNDqINW4+2l8IQtV57RwSUHcsu
yfAorrzgOEYLWjCJiG4YbtawNytNt7LHCNrzXDVw69KDmWhFRjnDXRzdzZfhIImQ
7mEU6UPI4To1yiOaA3X6gxr7dCqLwL5YTSOxyv+cOU10+Ru09UKtZsNjTDulyGm0
4+o69QuU+r4hlCJTeHT9HByTqq8ZIcTOQLWW49pGdNXpz2Hh3R2GqvLmLv0Oy05Z
xf8O4xBpYRnRc0QKVH1rYWUS7cy4RtBirsvDS4lRgIS/30mN2AspaHy3FJG6YJFP
GwehoUx0uBg6yDBk7JnbrqKaVD8jZYgXzxNVPWbRmYA8h7w6+OUCZmhO6n7b4QsS
m8FNWfVTPhZV760ryKqzLU2Fn3wNBfG3pNShbWG9Jh6dEeISt2nwiR5fjD6HDO2d
YZz2g/SGgTlq5zAvQe5AVvMFAOJ+Jm0lsc1J1P2FCjgTZbvVQlpKEeV/1cXXyP+b
T0RK40M1QyubUM3AWX6w2Pls0USmIlKSTtrvV4vcL85DV+CjE0xxINakkvAxHJPc
eMZGL/AoUb4daL5xKzDqQg7+4i6XioSVWt3kHcGkApWIOnXQB0yJt9kLQgVg5MR1
xjvqPHTNH7ZVJrE4XJYH2RZxVRb3tPmqBR0ONwVAfsJraTJxD6SpZX9QbPs61+fT
BC2l8pwwwjjJFmb29+TKAwv7goMKgkioYq4AjsYAf9IThIntRCgDmUVVeoqZLmUB
pLcmA2yFVjt9cdLGAN+JY3bzfor1960+dm9TZKClGx/gjQzbc4K2cetz7OZEYzI+
SWEdm5YEOpurhZHFDqMg6OFIy+ZVPNwsfw0maeRbbo076osPqXaJuQl/ny70dftT
3neJz8SqHzAWoi+6gMkx3lPmMjNDoaC71EiRC9CoZjeF0wxX1b+03j+kblq/zOiV
d6VsP4Iau4ulYjnZ6tJHbZpDYxBbVQCP5m65KrLpw5/93Lf1w5gjxvg1QJSQBEiN
BAQxpTjOxYqWUE2///CYCm2ffIL+aD3TTBnjbgEUroTob2VasxWYdWXgBuK0DKIm
bF3pLBID93V0sgOPL56sUQ4vpb85sB7ZcQiw2jCU2hOIV80ebAw/lPVUpMOYYIrj
vNFFAWLoyc1n1B8FZtRQHHSTO5kyFtCiMtyxRlvqe39uoGmN1I7nYvfaKuZV+QP0
9oqru2ydf0hx2r7wJYD+aiDvBSMmJkklioclqs4s2kcHEBtbVoSTtHjJz8ATBX3S
sM6D1FB4C7IUtypi8v4SUgHZ6uTnTB4uL415VGSzV3UWPFaUEmq7Qyn5oFveXSRo
AVSiZtDE8WxjS11tY8GS6pQvEfDhNZNgiifi27e28mSyqai/2Pffes682zYPsWA7
zypcTg89axRboo6pMGAuewXLTdPO/z+9EWOti2KSUlIxu8RSXZp8teVYalBZAR1F
j0qdevpkJHBMvaNM14Pr0SubKxYop6ZNdyAOq0hy5xtF/6N5BVBtFn91BQHtHkRK
MBBCdxx2nI4QHUsMHjcMVHLjw+Ac77VEbU2/x0yElNAot6mvlb7MTcOMEvMv26Yj
WSsejrUpeGpWcShCYSw9K1wKoKYvoIyn4oKCjo5od7tgPSbLsiL5E7ZftWUy+7R+
aFjlR4ybBAt95kdg+HGmsUbPUi0GmBsajzApFSkhG4xGqWJUtnl4e/yDU0I44BNH
THKnAMZt2aLArH5GnbinSK8rTuZxX6+SeE1m997/bwIqk5kLr7AjPL+c0MXcvcrW
Qe/N6Wq1h4/K5FtYoGfYy5wxFbxkibOmcLVPkLy5B7+5Zfg3weAO4R6BIYZ6VdCe
04epF2jCkZHQT6akQT80jHHu2YgeY2j1pQGvDYAyAkJ5vaFCRUhzGXD42XV8A81F
8Vl6r1jZGMfvgaRRxhYcbcoKTJHEv3idqToAf0HHKpcRODQs9ACYqgXlYIryXyQE
zN3GoagjEedPUF/I13JHocgo/+l6fn95YqlqYbHpxbXC5Hr14u4crv05yAyg2C+i
LmM4ToK7yzorNZMdR/2dCA05fpSa5S193jul5m8A7Vv5iGjywnpWyQ/MoYEgfW6D
VScK985QiiKUI/MKECwUhHwRT++SU0XS5GNKQVJVL/xmyQJYrBAeOklDqUalAyO0
97MqVP38rMvEfOMtZ1tkd+5ZS3KSyFmGL0UK0hhnNz4Xyr/KFz9A5MNYknytdNUE
EMEepMJS3WRG9MeVUM7yZrfxxbaGly56NhCMlrMWDKYeyWnsI2VqGDuRM2gLkM4J
gH84gp/34pegbataYxR1+FMbczJZaLiVW0KZkRbU5zCWxRNPOiYalvgmvTIWxXaj
EP6OSy8cJeXQfbeTPfiJ0MfFKG1YBWEWaMLr8B0XXrjwck7elLRtqVwzneZaNZYn
7pxDDHq0bfJEGBV5IZetmWpwFVdf9Og+rAjXYErG1eJXB/Ym5D2dqy1INuovNdDO
POmHPbegHsc0GM8oZQ3fTQVlVvAcqNd0f9Hq6gxiZ4m0VFmnHcCmxLQHg+qDHGt/
45IfQny5LFoQybyBE0wkZ3iv7T6kz5on++eitEDtBttfrJVYu2Aav1t1XYUfZg6r
1TGCuIzv+TlvU+Md/yT4u1TgfHdMCVfLj31ExQRxEL3RWYEgyFlzoie/cA0TpS0K
7e1phBFq1kWhYYlBVC5ysA5W/NW0VtUM40GGN8fMj74MQfFRWdWNJMwXgAMYEUA8
dsGtsp/t2/N2KtmwD1Evmpt6UcFUsVcqPkY6b242t8TCV0QMBJwpjmSc/sExnaws
oht+AdZp8qpbpuimZcz7sIa8o8N1gmVC83hZPaslHBNPznnZgc/+Avr//9Ws67mE
yb7JLvQlzzIgi1V2+RK7YCIjfUw1efvuAN4Jh+RC3HkTxZPFlqmUuTzmZiyUgxZ0
85l8VPe1KxfO3Hrobg8ph5Xw02JpP1C1TyMoMxjlmTIIAkNLeJhMQOEttqrbmwrv
GwhmCxDqdh8gb62CQKkUwQHldyaSoeYCZ7qwNFNuIw/La+PfyJZuYYuLh9YpXEpD
+oTO20P30YNf2Ee/8gX2o3A4OaO93L9OfZaDjG5uJc4nAeeWaa+LI1vts/NJu0/p
7sEF9kQH2jQWBO2pw5ZIUJNUAH7XxSmtOxy7UWBfzC6qi0pC8fyHOaCAMjRNuAJd
W4fj1n0exVToJCay430x2JZLOQPsjZ4OTa+VePVB6LTCjaD7glgaUJpKDr89GbEq
HRai2U+Ah5Z6IWnFotIlWZkewmMtN8MKSFUrtqFDlESVZYfmTFJWSyNS1e3uVI+P
CjyMoAVULPMqAjAdF2jjcYfMDk2RM66B3s2dJcmNsBO4UrcYMCFmx+UhVrQz5DPl
a7J5KuQ0uCxTnB3WIZcKVS06mDl0Zv+20siZWD2nzhL7JwnaFy8xscXWTRImH7JQ
CEowTjPFQjJbJDbQS2mradDUsLBC+DFf4uVRdycls9nT1dffZGlh1v2Ln1vApFeY
qmN6RgAzXH1TQshdowZMS2jcBx7WkdVimfz1QC4WrcBLHRAddyD5ATssVHiKoV12
Lo5kcmGTllrH3EdVMCiRq/en/rO5GgfXNj8OLjDc6QHMl/K2kg1XWJa7QeXuDP/3
gjIEaRt8gaEtRwQWa0Z6Xe5qNUCPse1/mpnhgeD3DoY22k+7DgAn+3B3IRY7dveB
vZg2l29Yqp+zMzV0rmpajm+On2n3ZbB9/oG52nFUgxRlPDi+8q0EYdPnfpu4XOja
5nFqRZp+hOJodHhktB8YvIDyxOngmqUrtKN9rvmj7h8zgdqExmMmSKQ+ZAi4BOtO
FGEUj+QF/adPhX74yuOClBMA5WDVwItSXT1fUDdvHHQbRoR68GfDjPblG1toff7w
/P52tHzO8Ei1i4RtA1rrdJ3dYOZuUrp5CN4Ff5SGD234PpZW6/nu/thGG6XiOpK/
O1hxJnJCvbaDbXXOj5TNVUWb4iC+hFgHDSaqthub8wo7fsr0nHsBZn27ZhBAzO2a
m8KRCaERrRLozouKpNPjF+NBlQ89arXQZyRGWhTo+QHGLS0arsoLauepMFNF8gtt
vnlGAqSkZNRayW91wSYJQGAIz7mO1F8JFFlhYPUrRQKZi+Ro9iV/tmcD2wYDPIs6
c40qBHlDErQBLXu9NWJzfynE+Y41XAy604tdPWi9ssYiuGeVJj5yG4CwzN3AUI3x
sFZtZZ04kqPepbbb1+nc0ycKET3pV9tb3WxKH8H+ojMU/Rw8PdUS+6jqYWE+VjU0
maFPgDqs2fz33w4yPzM56oE8Ejj1ceFbJndv4gUlnvPCz60kEGaltrNrORlf/tH4
129CECbfPqJJqUZTrBVo3vdC5m1oVmCGBt7XCORBlVMSXHfGNIK8JNpS3fxoq8jF
AbueU1KEIoPiGnzldrGrHoYr5CkBqyoVCbOE6VOF0onzDZHeKkVgutBnCeIQmRKb
vPYej/OuHJ/g4+54UlYVPJLEmpcwpaUe2Wm0XrvTh59aPUOwh/S2Hmbd9iqN+MpU
6q5uQEX56A/mh01krfbsn+ladVBEiDJAuk8ynvHexd4lSAjT4AtCIWlWznKuXlrw
b4xlxXmZdbLF2sJVkfrj1xO4cSSekpiAXOi5w5/FHW/Wi6j4AypsdfvHHjDv/zpx
LVPfXS60pgsLFhPu0KBnr1Df8Ve1u9mZXjIQnIWJwCuq7qWTyN0KCRIiueovStfX
OKXFdh8EASNSPGbW3HoqP9E5ux9lnWEBu2Yuy4oRtODiiAql8e5ovPqdqIqZZa8w
EOybAsYr/sgBlDGSIlCbeR+npxISwW5JkJ02H2ComIzF/XxI1wLY1WTilM+yqvBG
Hgv1occ5hnwefojyay6zuzbMCUxnagsrgeGn/AbLvVTEnF++1AbG3pngiGqZ/Op7
fKrQ8yARE19cALVHrHxsA1RoeQgrMy7WxR5ZbgMWeeFCTLoG3bOxDT7FRfxv3FHc
JtSev7c1B/8fscSwkiMJjmRAVBHbVSAEY14tZvS3ep8I7oPDPuYwu4SadUiYO80Z
N94nLl7c4gWweo3BhBN6sSsFAtNqeyHyujMPJ3tjgdIuX7TmNNtoMfbZzKv7uMLg
AXNzmV3qNC5JWqNllKBPVspFVovtAhLe8O5XjhARPaZiNY5cRd3LgiuYOU6HRdB2
pB9RWb7aAqQfPs0KSAerhotsjuXHC70sota/0Nq86jDOzROIHOoVLkIjCXN9zb6h
Rv1J46Bzeo/3sOOYiqAisUONBtJmCq1SwllDuQ+mQqLvcmmCg0ftKYNjB3Gkol+/
wVqOoePfbEOmMa12bd/oikZyaC0z3VglKe42uT6reeyrZfWBBPGh7/iX36bgpEAB
s2dpWuXPzIwFm1wPlGCIHfkM+A9YQusp/ScNlqseRX8ZMZ4cu0ABS0OksVW8mu49
6OZ36pRI8SC/PslesRYNr9Q63N7v4/DD7aXPdS/Nbyq0AtyZQx0MuHb1OJyNipoB
HibfjvSQsxN//wN/n6mBAaZZRJUWTPxlFpw/KvvDrCzTchZtMyEIZX+Klv5ait11
FInIBL2c+9nfVtbtoFoAmK80cVzzZtOZyNorilwvQ+wsPZaGxT5B6gtMyH9IAsiX
bepB6jzXn0sHRVC+K3wdPWLOPszgP59Jf1H3INET84UHzG9H9/kFD/llXIQnLpk2
RbOLTeAequZBYbsk9ZMgHEULidnP983VZqhIiJRlEtviqLhDl4oo6408VF2/LiPB
z3JkO1s29dDCnjXvsSoQrd67KTn82idm4g8YsutbI4r8uxRWqPgT2jmgpoy/B+Ei
Z6RNuFsKvwGe3SW4KzHSuNKzi2ZsBT547UHZHV73iE8PcRxFzUGLxDAmAdwgdJKK
kAXn45xpkMkWdG3QVuA5uOSYZBLfPQV+ymJ3C/3IwPGlpVflCa4hmwoK3NGxYOcd
sq1PA5Eej2vOo+oNhVEQs0nB+PKvpg3nmNXYpDqksHjkfgOfogM+P6yq7CQwfD2l
Ko7Riwz5j2gHyRecMrpDdUZwb4Z3bU8A1rp5dwW85GW6qLuAd99xQIHUFxqJ6ANW
wysc4mfkWVuTOWzqWcbA7r/EvTz3iCXV+4Nh7jgzpD8Pt4SgRKMAvzPJmCleH8aw
z9Z4rcfHtOR8IS/e/Etz1Nv6kD8gPh8vLlSBRprMBpaaxC0fLiWQZ65UiagHc4nc
KrBFjLxnSat9BmD74BREE9Bfl99sbkwf+hBh1QoPkKW2Gr2V3nBrbSfm8WCOUqB1
gOZKwYrCsbi2I8MKNT4WpGlnh4YhoW3a8eWVymIosDhrFmupOYR14KhOqe2UnMau
zO9zoy+1taYLY5TifJjk1Xjs5sybgHM3lVa1U746XChrg+y7KgIhKpKq84ZOiWHz
INyQh01BxPul6Y6UNrezYJAv06Yh9izj+/G6FKhSYZyiR/QddMXpXQCAXJpAzXUV
OPO4CpCSjp97XFXg364ZTtufqep5AW/lu6Z477xv2boYyJduZDdcl3V0LpvEZb8f
BqVdbPyJwdda/VUQbEl7oCU9e3tqhwDhjtflWSfawQdEhBpc+Py+l6CzLw49JWDR
0tFSHWhBZyPNad0XRhpX38XgwmRYFOyxf8YIB+bxlmLCd0AuPu30O2lGo7a49/ai
WfJoygXlwDGmAJhRnZoGCJx7EhjwK5H2HQS2BEvBQB6/NgL1aHIQB7cCeUBAf19a
blj08FxzH4t375lMYfEXqMo1QAWYDGVkkhkBQBLrRliTSA0lejM25ZpkU0TWflz2
3Ukt/bTVYQqguqk4oqzprNNCiS6BGsCHEb4Zy0Lta7KLgA88ygb1J5TbL1ivkyP5
WHJx4VdkK3ALBvDftFCnXiBhpDXDncaBWXPhLzJvP8B7pZNuhcZc8iUlN1kJkwtE
H9Dy3T8kDq45OBzKYaa8zl39kKbZ7jrv8nYbVQjDVN8bVycVvenEDFsAwHFWW7p4
dZTMqfvL/eDmC0otrKebPdXA2aPaHi90ANs2HaGYThp0zc97Fcog/2ukqOYmDaX9
r5J91Fg633NRWMqRxfiha50+LsQ3C+jz0iKfreeQDn9VITVyFl328ITsbOV64KA5
x32XtTQr8/GzdmibFnL9mdwcu8F7+zkD8s3AY+8ghvdWMxQgvdHMi5bWpoUKO0lB
R1gN8AXDClZZz2xog0YYUPqIaXGi2/MhPutvtXY9Ew3sH9aIm5sx9pAdTYC3xu0G
ww2sfgEFhhEF90GG2YjFOI/liht5ET5sHR8oJCQgESdnXEPLlPSwtVaVEBc1XNEA
bEJRe5yXiNgdoT8tNyqATT9EBp14xNqXntg+D4fft8LtJF+lcaF3zfjTue+pOhT8
NuKnU7nUxeuMUUbns0AGSPuli4EwlH4QYHvoLSG0vw3I8V7aobEExQHTtnVpZ9n3
m4SFAQw5xtEa4GsoxM6eg0iJtfcGX137v6YWiLVRWV1ciuGDq77iLZuidPOk9e0W
7jtCXnYy7zrWAlyVGFT8fg4llONAb6DDwETr/Gmk8i3DJv7FftTv7Cthu+FmhB0P
UcpddWbjqnNVT63ozzRQcJU3KmONdXekSe+CBAxSS63p9EliasCLl7yC1mkCEMbk
3p+Sn2rcROqV5K1OTYHEKZ1HyGzcMUshREdvgFeYc6BbdCz0XiyXV4EJl8NfENKm
8L5Nr0xNSdoViOVUiDiVfDteRz4Ug5UPrqvSearsivLR4RFPV4G1vflRML5ua709
xueVa3/g0F1fmgmZLdO7vx6FSSeCOUroqPfpGgAilnoW3arh5GZbCPacYR0WZPtE
z3FJneWR//T1/XWKrNEGamBardXiYYoN8sYft6ob6JY+2+QAwM/bF1MgGI7Hml50
a2M9UJcVX0nuhQBHtwIdRwuETJYP7Ad78o8yBOvqpKwXLFWmhCmV0fPiVUfKjzkz
fBFHilyAJs5R/tsWG934tn05xKI4SQh7Pf2rSYFSnMuZpY6LIRi6KgAW1gb7GbO7
PO0GmHUT9a9zyeVEbAXqA5UK+LHpPItLg5W9CYYHBldPv9ubsA8QkuPq6OHnwjHC
psCPLOhF92Svl5aRvIbLIqNvNKAninazd22TXBaaKvILa0KYGHtWg3ruCQeqwoAu
okJ6AKBzpeV0D3ieN4rbS1mmVbs8/Fox0QxWs5F71YF8BLL206gzIjFLpxHT4lrf
UWQF9NP9+pb0Ynvcma2RWG6+0JwU+cLVc54Pr4Bti0chQ6B7GrOeWJ9IrW79zh0c
KH/lo15jVRtgd0fSVAHBadOJusbUum79G5XZXP25+80AtTUiazyxfEW/6OUgSl3R
zjbgqOAlkAbXF3srN8tqPurqgVw7gDmrFr5zTgxtVaufrB2uuDwoN4avhuKEMqlL
3izUHgrRQvxmcHkpWnSEZTkj7/jz/FRlrkNRVQ1s9pNUVEC+UQ6tjKfUP/32XWiR
1Ks3ICjb70F1ZhzyxWStVYVesC3ilq9oknzEtIIvsNbhM0iZeG2l+cyAageE5/o1
RFYhfx/2COOAgAjqJy3yH1x3MScZBPjhLh+8TCwxbqRgUburez+45g+vx81BAhfY
xxpwMjLhzCk6WF6R6j3zHDl4zRWndJLR9yAMJGxbVfm6sR0YoEM7ahz6Tv6z20RO
N5Tp3jAAhff5DgtsfzWJPqpisY79aGizvwtTfJKV2TTETVixmGTKqjiEdywQIx08
Ub3Df6SCcE9KqFbkv3tqoV4XTHJ2jTzO30mFebEG7OMCXlAX/dxOsJi90ON8EtWz
REgAuD4KhmxW+0XiDkiyzEczZAeSnH7kG+j0IThoyn3mgmb7hBFfwxXcAQvRXtBf
CQaUtaW7wE2DYYvFy22fWw==

`pragma protect end_protected
