// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J+A6yPIvePE3nNgbpYe6EshqiDNsH7YLDVWb1xW3VYvaRLfaSJzvjdrZDWlv
nuH+aucbrLurXid0O9pVxE2bKXTK+STkn+ZCFxKIiLX/I6QAKN1/CGY6Vjbb
Wagz2E6hYEMhPAFK1GzWp7e9fZy+kwEnFmxX42pA2AejbZVPAXDw0yxH1q2X
X5d87S+59cC768/Q79fOG5pROU56fFFywjllUj2lnQs0tTXefrumYjtuT70S
gZRvP4bXY0B+DeE3NfO8iYZI9Y6nHO2loIxjGxG2zqyFMqzIw9COqW4d12K7
YnP8p7L3+NmPrC/jTnsIunl8Yx0BY5oCXb+o2McHDw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WvHUf/O4nBJKJrwy9i1wh60X6IWQ/rWoiDRlOmIhugcvzmNocqbmRBQ7V4dB
jSSfH4mobwOO5AN8orXEN58MVfhAaqv0QMp+cg4EI4gohXRHeum3wFEeG8HE
5CZ5bBrZH/Y2kE7tk2baZiScXBt4YVa4rBY5PNhrRqZVmd3VovPJ6mLFtNEe
RbTjt9hYbSFkjir08OxG929rtaj3UeD7do/aSgVts0GA8k3ZW36BDhGUXBvt
Rk7qrNM3jC5qXtVa4OAbcxIIZu6qhF52yikQ+fVK/IpdlAvtJkgBbpEk2PTu
eyLq5m+NfQnkklZ8MF9JFVizsTimzPCRvS3vLz8F3A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fiTUzWGohwVYxN7gkMJrKL2ZEQgBFAfuO7oAqL3fk8gwgR9tjNqYnk6gZx2e
jX5wOotrQfYquyBBPmU44ftkCFlVX6sBGHDB7sLjscp4RshiS3YKkNOEewOJ
Q6lrpJRByOhfbC4gdDdMxRwPgdbFUD9bEy5acE9WU5osuCR6B//QrmyzebZa
4yi22I+/F9WXQa5+/PXsTzYtL3hfbKFI/JiZwaCoeOf9Ufd/ko7jjZFvDXLj
YxLyDXEf1DBKJRU9FObg1e+sMCrdHUnCaafrCZS3cJwUSBXTNDlLJDjqr15S
EVTTTnGJH9+B9ys366Qr1tJHzyGs1QZKehrxErZ3Mw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jAtCGyYplkTOQ2d+LApQcr8WmgG88xGCOcHuUPu9RPbBAbAvtkAhX8t7vlaC
dnDSF25qstfwX/Gjskn2dS7FVFYwQypmtyJMbSsAykHyssiW7+Uyga6pNll4
6GEmYcmXQq535lzldBLfz2b9CHbza6a1KOONU38YLvyqo2FHFwM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
NPXa7nvkDF0RzNIczAm6w4tyKEpBJetQxGmg9Y1TNGszuQj2EQo6YWfDtA6H
E7a3yvEgCGNji5ZueJQ3cvxlgFoVNTvRKd/E4/7IFOBeYPYFBhwoL0P78QJW
w7oEUsOZbPs+0gZWRO1x1zenmAZn77dVu9FjDBHcspNhpS6VKaK+CC3xCWi3
cxDK5KdOPiwDWm7wUn/bJfrMd0V6QaNX8DumgVA+wd5bc6duHf9pu5yQRw21
pvqKtZwJMpFUsJSJ4UmkFtWW9ASSt+UDXQl0APyLzgNvIBGULNkfIsNhxO8p
BcoswLfAy+I911FKT5xicDnfpsNbvco6aueMDInYknSwOVIxyjkb5ggWgMLZ
Ok4AME0xC2oMKV0Q5Z/9z3XMo692yoSGGtxXGxKFcEgfWs7QQDMp8esWZT5X
YqN4pzPGSL+O+jv5i6+hsfXol3MU9mAfq5Jca8z1FN3mqdaEZj3LZBZ/j+DH
osPsWD07u9vR3o6h/oTBoNMOS5vrzbaK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
I4gkLQR42nwGVcBEK1O0RRVILiOsTHqySG6Y6bq3JHQsl+6X/yW69wRGBgbg
0qWoEg2KCGG1ZrGuKKLFQZvAutzYOxJSW0nAwciWK+xKqciv1O+qLYgaQHzP
lubCpweSqa9HsvxcpUhQqCO1g08yG/NtmZhtSReXc0N12/+y+3M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TsZV4N+VaDxHUzJtlyt7NRo+eFv+mXV3WTSSKxOJZR6Ce1ktnFAg2OUPhWUo
+9vkt2xBZnMPZ0Hfu11/0k6aXRw3AMAZsB3roQNBy+YW6zZUYEHLxhcUNdEq
iToGLXp9CSHnecK0eboiX8bJ38OE9qq8xP3jjs5nwCvZlAgSEgk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 5536)
`pragma protect data_block
OAQqq1uW9YxvTLv57WWd3aAyWf9t2VyKhTEq7NroptcePBbiZA0OE6TXqiR3
Q1AtuPwc7xYScrLARF00xBoCQ+ULy4qmE111a+nFZ4W0nwfqcYmeKUfio9BU
KlhYHrRqyuO/iLLOwiZFeiAVTYOoL3/Ft0Q2jBjPl4hQQwJZThkJXgY45XL5
NPYP6pTYIFeBXQW5wK9rtK4jmxlBicrnmxz8sZgclTwtiilSohxPDEIYpDK8
uGo0ksRTt3XvqJKJuid2/JzucdJtF7qJ9yFRJcbIRKzQRPgZgPT0v6G/1bqn
bbibZV452C0Cbb0eqNLWrIrvcTu7jdwmDxclk3wqk7atNBzLidSdzZNZyXUC
JYQ8byXqYZLrG4rtI1dFX1P6NkKqehp9lIm+ux9/T21oZOSMR6t8dTstW5oL
itPlgQv6LIckCSIIp44A0giZ3ooBbXRirtjJEipllovVf5UDS8kEnf4kNl0/
nhQkFTJECXVM4swRr/sCQEel7gWpUsq7mIiVA+B/B/Ua/Mtza9VC2x+wtjRP
K9kB3Mf+MRhEBhUgnEF9L/G9aDlEx9Nc4VYErPfdyT0KiAayz+OnupVlVH68
Oxb5XcIF0QrjZqSbmagJVMXn1VGt32N6g/efE5FoAsoKyiWPvK6/N46V9Jx4
0PTQmYf0DvVQKC4QfnXNdx5j0w+Dpk/ZgdOD7ceX+d2eN93d9uke0Angnp6e
Rxw/5Sb6bsgiNzxeMYH1UTJk55xa9EjrEjZHndTHt4dcuIjGUht8hYS2nkhU
TBoM1u0/ejreji8gdXCxcqP/AxO3/NeUSmrafKkyHNdDT4/xnW2SwUTrr6ZU
NgqSDv3mDObXNjwwEa4PiHaULi95nrqjQ67r2274EmV4mDcLpUKzsk0QJehk
1HN0yb4WlJ5UhXjS/Phj2A9pf9K8O5el3CanVNu2KHJFALRLDlGtUPETdhFO
odLo0+xoYR1+LGla6uXzW6P+e3rGVCIuIAe51K1KWKUjwx7pgEyY30KFRy+k
SKwhGXNm0edk4nNBYy4lqP02WtIcBU9fYwHNOXMFZMsnur3OLY819ayDirfM
w+hbzMSMyv9/gIEOVzofn4NxnDQi5ZSS65uYy1ThqUFfnKypX27NmTXBDtgw
bWEvqiZ2jGEOqctbcuCVcUfC0r6f0yoN9kaVksS535cDhtDNCJEtBp1LGV/H
FYbz+CkZFVyXhENKfoObgmUB95dTBR6/dBv++akrWYAcmvytuHOBRw9hMHLI
VEen3y6FgCBDXI/MPbxMs30JfX6MSe+QSVLoirArpi0cc4MR6EIuozG/ctua
5dy7KnxrJatwbuhQlvAvySxGOqYFKlWpgIfZbFJnmbaZx31zt9SdPB3oVz1U
J5eegkqW8VsEaoNbaDvwFLQf2zEuHpsbKyglzx6d/XL7INP1Mu0Khkyb7QT3
2P14kEfAqFSrOdjFZ6FHenCSWXzpD+y6cCS1h6KCi0vEfGKF/dxLpyr7CIkB
DZjAKgvzWKPW/3A6wLYbW5BjBuYzH+aNs7kQh3jyNFEIrvBOABs83bmhSlZC
x1jdse5g3Si5wAd8KfxioaBCMII4/Mjoc8/Y+M6Etu7Q8IK7C/BbgPlGUWol
cjQ1Ar4y1Lc7Xa1YNt499kW8TAZGGOKgxs4FZJKJ4vNSAsz/1visFkmai8mX
JKH/bJ4vBmByHCvgOLDE4HlEPHd6KLTrw/BUykoQOHqyFcyfgCAGiv/a71Dv
EE6YNumtoiq9P4GfKScDWBIepHv4YPReW8SWTQRq21AMZMMwwWqzSA1JuP+C
08/wFrGMnEyIVkHIVhhzn6V6FsWipNiO+8erZiVpj03zCP/zaNXpATUgtYcS
XuwJwzJYG/jS68C0xckABqgp11pzthJp7RFEDu6dvOteSqDRVOvfI22j9bM1
BafdVd1FxkuriZjPdm9vYUtsCTNOTda4wlHoRBwZ649TjfABiShyVFAxByLG
vNoUjtZ+pS3a/0komPb5beH2MncJS3/QqzabuplHddBBiBLfMMg4ETBgRB7H
uxFmv+9+U0lNn0tdCrjXdeiGIDS6BuokQOUPBNxj8c9BAfSxbm+AhW5nvayo
XQ4DvavzVn6Wut0qriKOFfw0gs0SxeLiRdYyTwitRhN7VQnkvpEhOuRsvNUS
fio0hCToxk1B0oSrXqnj/XJOO3EYRNZX4d8Z4se6+WOA1RTD/hFmSdnISWrn
hORW4sFpA8Om8ra4VswjLwH9/dPgGJPKW/2+xQ3VfkhvUAJnX6qoVKMWq5FA
dWQC2fzcwgG1wK95z4/OQbqWQbkdv+2M/aohKTkAM6wNgjoOflwvpRhI7WQh
S3CGuERucXWEPAhgE5Yc4x4RRIrVZcXEOxomz2HwB0uQ1o6OFJBdauVX7O2N
WKP2YRys3WoXNKGRrptTmwvr3VvCCXXQW1/rRoF7/eNMo4X1Ya+JzN/pntgD
T5eG9thpTcw7cKRIhrE4qYTQ5US+QPOcQefnikWp5ygTnePR/xx4hbjZ2VvY
0L1ONU6JRGNKZlNwMoOErX8NnZ2aQdr0G29vXUiduzC2D0YPIrJGSRHnjq0P
bTPMIHOG3wl1XimEv6dZMUZX2oBnT5egBspGYV3Y57iQuSD1dltSStTrbwAD
pS4nSGxh26w3EwdgpqoLkOnDVuB543AMtGch3E7ck5dI2EoGt+s2lg1ksETB
wk4aMGHVFo87FGBsfu+2cpov7Jp9G2828oKNrPYrApfu8LmGHiE5isWpmhdF
eYjTSHU6fLbjThcZ5jLvi4DKwCYzC2678T+pLgIbMK1faXTj+QVMuSGfdeSW
6d0a/kwn4IhM+deXdBevdDbNVsgEhtiWiMbSpcLzD0xB+bAYqdJiKJWU6/1v
bh42+FJbVp+EzuFF/vHRhy432Ld+jQdScTxbHnkaCme2x/ebJSWvzjkZtwgx
2g9ZLE/VnKRcbYMr4YbPV/wFfdvypVR6h5AG0YL8RUAUUboERnK6akvaGKhh
wu3gEUKWY/LUZ4G9HdDfV0c2Vn9VgaGbOjgIAEoebRN+D7y42Dun+GyzulKo
x7HIN6LIf8svK3/dL4ErGRZkog3+ewcDXozG00CTjo9MXT4LVarIHv8P4jDa
1Sf0SOweEuDKQz1FmWoQw1A9s8qmkuLz4HVKQI68sgA3Qw5nMqQWOFyINIO8
v61p1LaNz8KGRgvgCWKwyhFljvipRag0B5CnUDnAn59UrH1UyRoeqSmjCGAK
aMxI4WOrkiNyGH1yonPr9bmJxuQbjjXtZHwrstFa5xKNhZm2VG/Zl16QA1MK
TrQCOkAXoUuw2PGYcR5Yvr/DmXenn6N1Z2qVzPJQSuRhcmZ2uCZLkTQXXqtC
E4flwqXGgx5FnkTrF8mrWqKBm7dR7YVGvS3LkIcQchQXIJ445CWp19q54mLe
nvR7MUEGRDzFPgEUtS3r3FtSceNHrZbByHjlFNpD+y+zpIDhazo6h6R23L/x
G9I1yqmSxFvZ5Evl0OxNMBJU4vaR9jRA6/1LorCutgis7W0YktNasWZq44v4
iBDLbIxB9c9OM4cJ7/Qbij07GEdttWVrx2pgNI2a10KaryjLZtpDIyf2ErrR
S+XzFbjg8BlsMvVg08Fc9u/cSaCkTPIG4fvpeIEY8EcuSqr5Z3/5uvJEVLHP
3jfZz5SdWNIYcI1KatuGNiCrsoRaCFRE6siEkiHrNvzPSGuUeRVQLy1VnAug
mv9HxrIa+clhDY5X4PU2wIzQ7O3AGBIFx2bFRr9xUjUy29Lt52DBjy5g7rNE
lJEnP4l7Gl1GXjpT+MGnLVotCh6OBeb0QwWPsUTEDlnngeUA6TYB2HnFEdIl
MS80pPVd9yGf9z64N4b5nrZ2RVvKXp9CwTRtSqjp/fMW4h/Hn1i2MNNLFS8U
uB1VbgbiWR87fE4oDXiJYWhrAV7fcdoHTYILh+dDov2P9sZPeEt1rgWaLLvw
8XzRDyMhsysKQmgC/KjOsmUf+nBNLY4+HI1G32W8HoRrcsahpWi/jNW1QGWq
Eib4PiikwF1aGbrvOu9yhWOdf/FriLs1uMnufKZHZDrTmwY81NuAkAW86NMu
361dlc49VJxoP5kCG5GuaYG/fue9qrRs1I4AAqP+J7MOVcPwIX81i0xmwLQ2
f5l3ck27asef/migD0OnDLQjIk/PedK5TlsZCmI1OePTX4ybMZmrLuUpiiVa
f6fUG7qu/ouLsoeGgLTlpcXI4zVoXZm5wgOFm4VF2syfeHB7FC0TpXRK9sbp
i+07pd2j/AhheytYHYx9KqEiZRLanqepq5/ILB71Wx8vPs63iQlWr/SuSaxV
qkolM005VkJ///uRjOo+Z5eo/RdMFSdJrYcZCUTIYQ9Mta5bGjrf9fCQNL05
kwaCH0bnsC5YxDFsSrhDigpvhNhOcW35ssvrN31NqEGZDU5DW+cxpB9Y5eg4
mtoV/b+K7ufeFyJH7shYeNLGWy17eND1rSXVG3H0D7rElMt3/+dUcFvbJrhs
FJYM096guE1YEvzdPlfemG+f/QrvWVceY/g/M4/jBlEhhi1zBvE4hZPNeS0Z
5gk99f2CNo7Ds0389tHh42UfvE11qkfWTFcnGIDN0467aXHnL48UKAob9DEL
lPhJnGm/Ub5c1pNuTlqbGvu1w4LbF8qz4+dSFjZdBqyqtvIO/78Mc4iK3mU2
m0vFR9kcIjkwPynpSrRqKYEcYf+li86ziRb78bVRVu7ChETNFIhcEn8ZvkHT
UtRhC0diQmXuzy1OAl11BvBMctoefNlTVMIzeiyswpMgSarZP507i+1kO4/A
xqjQyJM3R1OYwLDUvTkkQgnsLPu6NxLv56DjadklSlGmOV7rYNSeAFsrx3O8
x14SFtP6oOVS02ZjFPOqNVl893sQyzdoPLE/nruzSXjPMcSzSTILeuCm6O0q
QtanCRIT15BCDRVQkhaYWVIjhsJ6CeUpkXdpkvPSzf2VruEJELAtiIVcaOnM
evAq5MwUp3IfmWsCMLpmq3wWGx6ZEQgqrwOjNGbejNaBDOIgkTVvuSWhndXr
sI8XI0xnWmJMm5MzRoNQ83H3I+RPLaSOgi1OQWssmCqzPUwFdBVOC/TE0LLz
v1UVI9Bcv9xqfzFcXJ5qzxFpX0UkjpQNmfjQlAjunW8Ec4iRO6r5fChp950j
FHtHbMXYPT1hf2n+rII5GPzEzzqAI4KFz8hpNj91ND6SEitW8DMTQD7FXH3f
wG4J43HnHQmEvTbtswDoAtjzQq5PGZiByKSrkfpWZ8PGu8q8+GnqN7LP4eLo
CML3dDro2PYHZ6+848OW0+BEzqqchiWp60Ic8pkJTESp5bbwrmjXdW6fzw7P
l/BYIzcPx08tFSbK5VISUVJQPiWKXk3R1orzyvQn+aJSqD4pOUKLVCLu7/Vi
kC8DKzk2hi0gMbemt3LQ9q1H/UKiJi1gCDv/3D6/tMYN3TVbzxcdWx4r6VUq
fsdt+1OXLat7rXPH86VxeAd5ZrB6W9z2GAJ7A987xw/i2OOVNvB/l5eqmi8N
hNPHHH3/OmwlIO0WhLRcP2zWyU6xTCWWtCuFjWB4UrPW7W87vbfwjQZhSH15
dIaWWAiM37g/6xIC0l5iggnRSiZ+KzeOorvALZ5Eztij4SC9WU83rOyjW7F+
MIEztGEbpAr037BWSShNIO+68ISUYkx0dloiU5U5tDnGlPSxgb31z6r7pYJs
KuqDEIzn+LbCUtkY7r0gWygYbk2JeNrx22FgTZbOrv1vIB1y2nMrdA3f5z3/
Lot8mo9foUykG2eb4/rfkBkxcVr6Vpfm4bcuPQZFGizqBuiqPdVfRUuKY6mA
NeNKc996L6H1zR1bBfYzVI5GAFFLnRNMlBZUqQXDALvNkrBlGWL02KQfzUy7
eK3GecagzwDFaVGCRwHlyMgVykFz5emPGfAHhZ1oleYoYEHsXuqU6FCrJId6
fhrRmeQQhHiiNApc61eXuT1d0s0HRJkzspv+ZezX2TNK1xuv3ueKmfr8H/9P
3Anyr92cGrYmx3fZDWK1DZAQLBqDbuA0MGijKrCg3SN9xW+g7kcP2Gi/65g8
3e9Flf8xWeHbFKWO6MKUy/Olhq4tuSJGYrm1g3Hkp2V6Lxv0txBHgCKv7v0l
gC2E5vb56SCXMvDECM968MqR67hkoGg183Ly43nP6fYaOG4EbnZFuh4UvJpI
6HbJUlzXcMCS/z+QwqtlGM5MS6CAAA6rh9jHvP0EN0HxLf5c2tzwfeX9IETE
hxmK+9fEA/0rGZRxzvp3v7XYKJhGdqeVUAthTnGvM7IUUch5H2BF19hXcmAt
vGWys2tAu/UxKAELA8YlIaKh/qRpVZBb/6h9Qu/Jk1vgjMMw35v5ExkIy7nY
fYe+dIZSaW+H1jzkDewC/SUS2jiL5qYauV2+LAmJswDeVPESTf9wSdIw6mqs
5B92cJylbHRzQXIOVXhEk0cGdPRltxCNJseQHjcpzA9GXXo8mPAmrNxsbsj6
+Ej3ggAlsueIy730Kpoi9+uAHnamIhMIE7OWgOF3Wn2Kqfz6buN32/kIkM+W
1oyqRg+TGI2IvSXHKr8voqcw8gpNjCpAaNrL95UI9kOzUb8aKaDIOiqwX6pl
rP3b/Qf3WEivQj8pkEjsMGPSeB9ms9nnrFuOjScsC4Y6/ujtNmXUTpl5wgrf
elrTWErC0m8KNi2VWlE+wBpvdBKc1ilSg7QKKA6hFneWMJel0QpHBBs69E00
0EnUuyCGXi8UmNyNaPo6yzyvLOCQom2KaMv5Vz7z62Jnu6FQoDXiSatCNRlT
ledtnUAX9t9/82XW7OTu+uLWJLXC9vowCO0UxmDo9T0MMbouxFSAtxk7PTT+
6kCqFc/oRk5lb7pXVE1oTObmQk9Y1G10bFNHPCMYvNL3TCdV6yqVV204ytv9
ARUop/BQNgkB/Ky1O/qCD06EdkWOQOq+2ZtXJFzD/P5lvhXJb2KTXDsTl759
2xWvdaS5Li15ZA47kKIL8fxCFnPue6DvAl+u73fGROqBnLkDjqziOJLsoKtW
k0JqB8DSOpYxzXVOwB5kgG/Rn5RfhYoAINaomoh3LhYbMJ4yG7mCObaeuZen
FSD/xkHoRdYA8D1+mxX4BFa61+rHRQqhju5ASbztJdZtcvpSCMJ0qGI1ZelA
7x6fOtHN7FHUcXPm8Zgj+SVQnW9OYF11IuW3q8R2MkFunmtxaQapjFJP5jKl
wahceE9BNu5lt7EOz86EG+LBTUl4baantjfzrZu26TytteYF24G+paXMpDzj
cAx6zN08HJXtjARW4O/ZpaYJXYCeo+DbmSUBtY76hNsXDqp6uplDxPo66bHC
VzN81ZeaEVvkhZGBJgsv0Zjt4JanbEcDEwzAYHDQWZv6LKbpSEldobyj8n3g
wA==

`pragma protect end_protected
