// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
yObAZFvaa5lvVzrAfp32tJZs0/4VtqTnQvApBZu+yY4zBo4nHzmjjczp72RD61JU
HDHL79yz2AyPsgNG9Wio4/XVFWKWe4ax+DwTfhQndut19HdX75fwglXWgGLecAza
cmWYHoffyIQWQFSqC8cYP+doEYZFG2H0/KxH/P2dVQQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2160 )
`pragma protect data_block
rf06P8l3kMZfZw3nNVMwz6X0YrFhk0VXSDgDoQmhw72o+SrKtaVHXuUITnWp8Afn
Zj6wHJJ5wUZMEKIVyLMOsVUkXUbUW5/SNE3AOQBRp9mtKuTvYmcniHSLolXKZdrj
652VfUYB1EGkGOCVGOZ/3V/SeJQ3wvcErvrbmpquEJeicGPxPuNOiOEB6uNBl1Qe
f6yWwSOWkwsjvzbObNHhR/XF48CLfen1hPJ2Fz5IBYaWJirmlE4tlYrKMGe7Ydrk
7oV363is7HwMJLY88fXwLoD8yLNNk7FuXHqngMXpB2UrtPIgiLlm/fjm9RXnpEoQ
MF1SpPO/xV43Y+6At20SM/PpsSNSikIGBK/JEIFJXswIiyrqc3rCEaGIqiau8cZi
WgBgkkV0CmFJU7V7E7lqlC9hf5htvFA6p0taYgW6dQVRIpAG3LcNVVX8as0h5wd1
TEitQ0aVWfRkD4Fs3fsjqIxk7eQ4UrS2ZnpLZag8rzIuFusB3Gs1KjFSV7pWukJz
NkzGcmG+czf5a7vhVEmDnXDxEqfjekcBHwUDHrz2/REvVXES136hyZGbH7p7cChA
x40lB3flhoynoSqPQAqUqJB4HodHLoW2HAbuCjxHxRNi75F511snb7gFVi/99gdY
qMsve6E9zAcKuTk6EWsmUD0aE9Pdl7SF5RWFX6xe4/6PPjLsxyMo/m0c5cKXOWXL
fOqp4hB9H0Nb63Mgp32tVKJ6cgL5x3NT/V5XzO6WIfcJ9x4XdefQwNFIvy1u1q3r
xJqitI9bjRcTuTphRHffHL50cMG6l3bqG0cD856vZ03U4k9zlOTAfXHmk8SWIaKW
9fglzyylCUGyIpauU8ZFX+uifNGethKQEffq9E5YOhu6uxF6anI+nO3Ugj5rEpv0
jtAoj0eJpRGSvhJBvCNtTNjPb/b1gRW0AG7qovuo1DfoB4Cqaupo+tpsQF2UVyi/
tYGb8mPFq5C8gjq6VUvR19Ody5oyDFO0owf2yQmIf3JSm8CVOvLNAsuX9i500GL6
VrMF8oEpmwEfgxCUD5f1ddbzkklAO5ygXwLu41s2wKRvljz4KUKW8rpI+4IUYI6L
EJzGlrhbUy+DLVFaYn8iYorWaNrEXSSLyDr3Bu5syVp5Z3WqbgaZ6DmHkgOtmpBo
60M0y0Al230iHanTkNXv+WBv21+ZZjZnQvq/HL/0b6JU59uCZlEodADJpPNV6427
MeTjXXdr1a4nxmNs7Vr2rTmSsM9eOnw45/OLLjG2QTRJg4m7Fc+QH5Rq59wyOKQK
I1IHLCvBjrTitI7MKfyARxcZFAMMaBCt3rz0fJ293LH52JKaHmqi5VUXqllr81OF
qL4dW4DXerhdSekeCQpiOYmduxWbrwYGDHarTIs0My6/iRQZJdB7xmBp73tDALxu
jIDLemM7EjNIRh8a/IETTyuOZJTku0i5A22pomMl9bZZO0qT5S6/Ama8WJaIT3uE
MjjvJodrx1J5Jo0yaX2OokFjdyif+BHmLLho/fS9G2+HOIpsybKS0+NVaTVGiLjT
NkfR+s8vJDHqJeH7TGegYV7np4fuV087Idbjz80I5FuI7QAwlDS4a8+NKZzhE4Dy
OPbv7oN1kTaW8sxkaFIf9hD0htwTUN1l7dCiJtJ4rwbuCSUSaR6p2a6FsxO6iWTa
5KTMGBDBQ/G4z1skjbyFslFrYf3mXCP+IVB6VxKJJwyXrC2Ryf6CB1vsclObBKsZ
RllL6PkBZNYinC9Ergcn8qdYWcLmF9CzQqNctx0XM+gbuvHC7aCSLLDI/fz+jwZ6
mhtYAdFZRvMSMX5ZKfuz8lsh64JO+JcEG+BvoPMVNvlIVhBn6WsObe3r2ypvclA3
fDTg79eExeuOABEUou6BYGi1yFEPvnwbQU1xR1BWlWeKI2c4DpYwL7pj7xUX//oY
oZxs0S8l43PXazFlThY7aMh+34yihP60F4JiX3GArdxUh0FCe+8pRyT1y3JHL9ym
C/oq/uLF5z1Fjqrcao/z39YOpPTbCxApkZGBCogjAJn9S0C0pkbGiPkJlrSEdZNs
pG4sIUYKay4SByrfu+oSG++RJL/BCfXrd7LFtEl+7ZOnw0iRutlrTuofpUDyqTVA
LZaDWCeSjgsoOAnjhGiI9L48jUDrAgwU1ukkN8ESL3z4d77KfrhklQicnJrwv37a
S3Cb9iDgEfVjJoxaqdhWRwGIANprScCFwkpOlIzFC41W/bgnEOIDGL3hrMPU/3Od
ThK5XzfLkTGIgDa1K+crn43TQuENL+XOuTfZfQKRjiDCjOJlLqCYp2jFMed4St9q
UAJ6i9k+xD9owSWtuyVMVSJeg37LLV+r3rq2xiPaFErJud69oiN/G4TJQpsuHFUP
ZMJhrsGyNMr4QeU1ne7EbWKSWBQC1VfuCW2Uw/8xiu/h86/NXvNZgiw8b93u+9X3
o56zeoBiIvLAGfoc8PeNvgJKFiLz1f7Or8tJByiGZhh4j1aeFiwGvjc1L0lKLzP9
Mught/VzibvpT9jaJBL7JB5wDnl5lDIRpr4My7mdpkI3dxBCoGJR1gjBZH1eOSrQ
Ql+P0CmRSrE1Bg3jVy7xYlQTG5FXHM3YvSmb1sp1VdYPTTL4tw1iaLswnwCKNRB1
uPg4MXDJmYpkmTra5yZ1w3Gv3+IzEV6X4/+kicqNvRpOaj4gDERj6QFqj+cos3Wf
kbGWDxjqz03RBOdk0sqNsF+Tuz4S9IDOZT0d1vpCQQ9bg7dCUiPPeLE8LtHO5O/y
IjMkBLn1jSVmSIYJRFZz0RorEeR2MobKtJXE0dsJC+1jaAI6sjzOqwJei4D+PFCn
Lbe3ZyFC8xJl/OZjMuNINwI8JJsPwsO6MMxRZAX4as+vN0bYWleakkRzwYw9M2+M

`pragma protect end_protected
