// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KDXLIf4ZiV9h6GChyq5aNvDtZfq61FopD8H7QQFTSY4sVQ2zNo0m1s9uf4Vp
jwBirV/Byhe5VaF4FXzSLoKJttZcYNXS4WGn2GBV7SWynAIm/zBxVwjTbBU+
8vD5rzSsK4z5D7oy+aGZNVKWSvbdwZ4KEqamtLtQpHMigos9QCD5A84fE9ks
+JILAKemlkPQLMJxpUH2nL45DABg74PRSBvD8uTTbDl9RBLCZLtiyHHUqOJ+
bqzEAZIagXlm+aDHz533vFu5R36Yu4LxKa7MEi0kvQIz1ESOyuZtUX9yx4mD
pLVe4BgfMkdeTn8PPHp5y0ogN7/ItSnFlUb/JUWoIQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jr1Our8n6MCrkkM6OdbS+84TfOKSmfRNm54z5BBcVCK6vJeyoLMNisvbpQsN
MurZArnf1V51hUzw1xbAsevK/AriPxmhmCn1jSQnNWBFc95gOl5vZbCmDytl
z1eDSERXLFuKvBzx4LFOJJjbMKYgF5DIa9gfEtB/dWh0SDS9Gu6QjrOshKNQ
Q6J0VIvs7jrij2Ejhk7UNkDco4Tj0PaS5qEHFtqyHWkhfqTfRrZJCZ/6Zt9R
6+m6YRvSulMelqvHsgImEEat173fIAfYcg405EY6CG7aKCMEBp4s1vmiVSfE
VSoJejTDVgqvhY6thMDwNwWSQ5ALGmjJxoXr68lzDQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
C3ACdvhraA/Dx9zVJ1dYYpr4MulC57eBRwxcaSVJbZUvE8ifPcG5968SMMGi
2TAVc9476wLcia98HAZBaHxHRUdkM/rhB63RUWiMGXNP47GG8jTkM+wV/jfA
Br+pxsjhbgqKtEhobNwjuV/12KJczlBgdNHY4rNP/naIVIDPJqdbcwnvbMkI
DXdTbwLLSh5+4aju4HaWlIKSXTEDDQaIW1W8BViYZKA96JY+ou08SkiW1ntv
MdFX2RLPLwX/ORoml7644BrRnRQR9ZT2imMRWRMwEBzWnglpf36gu+RWMmsQ
zhYksXYh8vu6yIuXJqi248/Mzm1BYktYOnWS5KrJIg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Kw32H230DsszcKkcfQmeMXtFxnf2E0+5wub5vId7Bl/1d4kGgFUqRKbpRLRe
2RC5sYbPpCwEK/G3iwWJlGKtsyPVTD9W0snZkGQqSsXMlWiR1fzWVZGxcqy8
NUHhbxAm72L2LQASsNzS8gIqtuWSjezs2+FNo92kcnsV25jADmE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
jewsD3Ca+x69WgrMajZDygdSEzeeGQuTM60aGgwGx0NAkyhgHrOmoCbZ486a
ICl9QdzsqrnJFoRsgXxQunFynIIKP3wgkrnnlwPcV9Z/YgEOg++Osq3WJwjR
p39S3kmB1dFa6o/K/j0U05m1Oh1/t8nL2KJk998s8RSonSHXiwDvfSk5ztEK
4cjdPMA4QVhNrm538xFrSx4zn21ifGaftWdUsVuPs3tleGohKLpMJh8bjodM
58T83G785bLflUL7llrcIaCTIhIJxnkCmuRJnLSzF3aHFVCTo4INfQTcOGQ/
/+PcBvNIc6bGz5laEWtTITWaE+qJPHnsDM6IL7MRAiiuj9XpSUrj6P6+DubN
xq+EMQEqvvyATwVJabgYHG7ys7zNIbw2Au047po4oqqzSOOVzLi6uaTEDuQE
K1XOI3n2lc27aWu9pOHAJj3z4Hh0m7GP0nGKAzo81HHkV2Ns3OLuZWI3EP94
3kdVr3u8U7nwmKO3oWaR2vyPbRsBh6U2


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
avVqmhuhDooo7ADQuSONgtx74HkwgKhBGh/75hDU6X3vBBzKz86p3gzgQbwd
OGikuCHmrRHbtIgWMbEVhnywCFhJDzi5z8vxMLr6N0hdDGoQNOJth/kaEcm8
6qh1HyhVP5o/GsrLGdn4fOrVUXJJfcYRuW31vGJxw1SvIsFzFNk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nPI4IjzwD//k/gGWYbGyhlCSLAVwejo74HjvUGlJfM7cIHtcad6sqS8RdjQG
NVYbPy3YujW0Bs8gicvLvPWed5EOgcrLvZaHy9Km7YjVQFY4E+4+f2FBrKtT
xLGN9yNqIPAzeXQnROe+lPq2Qcj07m5jBoffVpAyOmwTeBhvq6E=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15904)
`pragma protect data_block
tHC0LE6QkW1jwe3wmwaYygMHJNp+ONKddLl2su96x3vpoKCCqxIlM0nsNwcp
sE6BHwc2WQqDFYIdpnrVJdY2kVaj/jy+nRGOdUlYlOUIoOTP+rKpmpnjPYJa
FjkbjYRojgem1A6k3BKTmccV/S16ZW7feniUZ4M4TC8w3cYYMpr4nzM2yPBD
rJcjRcZAR3LG9oHgiuANXsmec5VN3ZnITTDueolhoZyuZ28iyb6ITC30DBqP
6HBr9syPY4B0u5EGLuneoQlPiAh3vv+kuzniOJCs2fKbbH2/LlAgcLB2PqNT
pZVm/gpWRGzZWK9cXf2U3QYo0tb0qJWuw+HDB4cjXLiaMIDR3y3Pp09ZOzfU
mJW0WjZQrl2aJuXTioyt+Q8L3Mn8FzJU/g0ndc7Zeu0o64t3LPpa5EJDOw/5
gXPxKz8N2XxdePii0ilYfi/f7TNPvTMt0fzBKJPNPOe0wC+TFrVGbiSuEze2
uLb1vz2B2vW/yA59j+GS3Yz3V45QkVJ+PcAWOqXhw4mcv9y0GEGrArohywR+
a4owG/6MtBvlWPU97KHA1wbpo6iqf9D5454VYhfinSK2IefjFB/sVBgKf+/P
nnswECu/fQ9hcXEiilZUq6uCe4EpYKzZVxoU/C+CziUWpxzzI/Eat1r2bsFO
IpxIBmLdJ9d/vplNPhNsjs+vNQ945Oqe/+EnAp51WNgVOqDZdxoQTs36fn67
TgjNTQgSFaJSt5QVOuPbMZUN3/5o5gsMrV3ksZQOwsqvy2ik147HPIFFYnlp
TfontryyF5k2657XK47zJ/qsGPAvoEryOuVmpro3RXmjJQPO5hz6gdIUQ7Kg
XgXB3w/fJvN5yw0X4qPHUONt1Ref41uIRvxzRlQSJaotk30Iy4z1PQvLKmCT
AArKeZ+iniA1IynypIlyYu13dztHnPF5azy164246FbfpsFZzCtKUzt/dPKB
kbu0IRQL9wvolprLj7YGPRkd1tvYQg0YUUo3b9IIUfTl+gjWnHE2y8v7CKCK
hSHzlzNjmWMcXVOnstMUjyEJ03KqqlXUPKGqKOLKfrcwQ33LpBnD3YhTxaIP
2WcVaRwvxL48avW4EKJuykJr7mBVXQZVuqHuLWxube5yI8jAWm3p6Jd0bkIT
PsGd+CdMP83l1Ak0QYPbi2MXb8eXA/LRkLDsJk1L4zYf18doL3z0OP2n0ryj
5xoi2tKlvObk7zp2j9S25ojfqVp6SJdcdjTPsTsZn9zMGNWfd1E7IMWpY9ns
mHZTMBpDuuIdBs8e0FMDnCZ4uJncD7vVX2MS7nxNVSMa19Hu+sz9+tIuGwnm
mn6gzxYVmJoZk/HPAe/O5Q4XD05f5HNzYmaEj8Y8y9y9n+gJ6T5qn3/ypaVY
W9aD2ne+/YMQ4GQZ67kibGDwvodVzw2L0rkkZr/E7KAtySyzxb77NFupU6eM
4gp1m6C8q1t8ckJrL4HICOI73oMMMNXMm71xfTcaX4XK4g7WZWfHa1BBYpDO
j8Pc/earDNQA4EZ6L0mYxfp8ZhSIkdZTN4cyj5f+tsQrh0GLZosXY6kQLT19
OcS09xjgnRAcWsc2ZUnmZfHd1/L1LY4HJ0BRFDYsHfUr2EqYtUQiR5pN87nI
+es+RsCo/1IQMmXOmE4AYocglKQJZPuXOhKsqLPk0gpnZGBFoUuuEdQPxqrQ
HIknT3deTvVuyykt6LvShwr5yQiECEPImKLfjhchAAoG6W845+Ms3t/nXBI5
PqB29r/tgvOMPmUvqRgNjZauILQY5U52XY7O2LrqpaUwdILqcwYc3yYVTJnn
MgKDiJ0qXjLOvFL/8HDLXFx2qPA3CkHF5IGy8rdVyfeKI/olFieyDo6MR0wg
Xd5OI6P0Oi1fm0UHqDfEEERdRNg44suhmeW+8wB0/EyVBqx8tkOz5Xi2zZW6
tqQgQD0hTHcAMxRa1ZPmE6iTeo04IC/6M9zciK/QZkCO59p4VrM1V/58vnO3
/dgLW4gUSmTSrwi6VHVAigeLJylp6Y0ILE664a0Zt5+DLN+SLXiOcSPs3B2S
9mWHL70iJzhy8bSC+4P5uItn+j17HXj2DZ89CTO9kGVN11DZdLbnCdAoJlbt
UuTn7f4jUn/vONn2JEElIWVhM3doEBPyAa/f5F8JietBVH7Zn7lyn1gvdfX3
G45Y/h73YDnaLkSIhY6O7clJENcbq2ASiqbweVl4TKDR9zJ+EbXVNoWmeEzs
jTLh6ljMlEn7zWjsAis1PNrTuq3CTGRhVT2ZJb+jXnZSbRsFbKLTO5M5Yixs
zxvwlhCLdpfG9mKNf11rwdJVGtJLAoKuOUt7GPoo/X/VVMUw4RVFWWqMNdD6
Mx8Q2++ODVCj+4csu4/5txs3GxM/KWx0pv0QhmjCTeXKS/JDmQRepTEYS69m
VbGmtGLOM+dq+fDsX1zn2P3QbT9gHvG+OyNz4jI3n0SqUb04kpZiiTP9Sl3F
6UYpdY0GiS/lRImgU3TqEnYsOP2Z+err5SmssLY6q+2Y7hmCLZHH5N2ULxqK
H1utQjS/fQn5xv2v/DKheNBTj9Qi0trtouChaGP6jpkkWAKGq8dM0NXwloWL
O0xcpU8ROC22Hk/izMYiNA2xkJRj/pN5d/zuZtwHF1tH+PW5DOPVUQu72sGF
slVvlHyiJ6o414cThAHZeEog0x59q4hj8+Y3z2KgPZBkbmB9ybWIt2sv9wmC
XWFpQSZSsPWRLY2kgfruCltVzRSA421b+7Xc/dNrhCK6nL3JEWu6ppwuzQoB
mWr8yGOeZ/tAoXsgYXMd36ozDzIhCTKWxGARpXvCh30BMVdd03mjmzFGbuV9
jFop5cIGrgsj9gf9WZtjTXTNnXnO5V/RIpg/csF8gDllLJXQARoO8WKJz7Q1
N0vP4/kdgvrPX1NqQe9/oWAdEzlIhqk4QY1/h9gd3PYVQNeEmv+WMf6ogrP8
AkqTg2eTYt4g8rC6qHIx7jpYEjl9GezYezFqX9auiNxvXTyOTJYiB7G+HD0A
FbRsIawPyBPlSHZEYaAVe1o354Gi82TkT996xcCgaRHkZWN1XH9ASUK4eTHj
FmIWmIJDuV+oRC6ocS0FqG6aXSKd+CTzGdf+KnemNeayxO4xfrcXgyFXJuuT
HgFJmtiTT0IMQnPROWFmeWz10ryRfXZF7PDrS023EmMLcj4afGBXCc6uHklP
coW7tbCCrnnStoSi42Rl/Y1YkX8iQDuyiSjZYOwkFlzdMIXJri4inuzVZIY2
3XKz3qtUiO6bfvJTsN07//embN6NNPnGrPZ+oS3jfBtkqw/xoJzs5bwC9GXi
NPsauYMxECUKBu5m1e+KhJnH28eOkfpa5c/AIFEsbr6IFAEqDyk0GJjNLpo4
htLLsPuifg1V36haFXRA2h+aY9A5qFj5W12GitmZ3y0o+tyiCLPjrwPFWmyb
0bzEgCncDxNMoviC3ocSv8AHw3u/1RHawphyC3Cl9ulHcQ8SPqyWKrpQyfmY
RjnZFBnzb8FUzZ/J2GsIrjxzg5uee9qWnkR2TubrrOI6F8rJgl1ewHhTw3vX
hVVMC4lHNSNV1ZBtgsS7Q4dws6pVbaMKL4QDDcwV7r/E0nQjKXsyASfEZgCl
RwHjROoEJafY4cGD4w7zWupbA49ojAEp+35xJcAryBSJgdSz8hQFGDue+Jg9
rZWFGaIFe/V7o2StILgP8dzwbIMe96UWy64yM+qtxtdBRIFRZ5+JdEwoFeSn
oxkz0LynoAdHyRlxQ6tQStB2bMC/iUKDuRZ//7TtwJj07LUAiL1ZFvYCvsqa
24EED/eieFXiNlh1PZK4edrPuop2cyOB08irkQFATlSZfrzdgR3p7wMGJ/sx
10W0scJHxnFXZ9CNLtbafJz7WJI24m12QVWd3/DeQIB2tmPAgTq7DtDZDHnb
LEtcEQZiyvQd6YcLFwu/k8HX1Rn4oSQfvRYVqmxwoS4POsMDHpaYRKwgJ8Vk
8LoMQPktLjnbnw7NNOS8IBR8iSfltRLoLvn4xr/dz1JvjXcAkbI0GB9BEVsI
SfDQVbLw5C8ly1CVPy7QX5akjJzv755ZSH8eFsXCl5Bnxjpdn8BNk2jKR19s
//ShLvm1rBhtqTpSn3Ry6JXVhSBx0txLor8DrUNn5vlq6PklTuy71v1IUttU
2qoQbeb6q1knv+u2m/TQPY6NzYFiDKv5eRBvCgEl0fqf6yUUBR/ZQlX8R+Im
vQskTguxjBZxn5J4Iymw+QGFNpxEzbc2hVij5ZWvUUj/9johUSaqqZT+oa1o
u1ymA08ynuk513oWl6Y9M9qUGhgdims24wlz+PEyB47pUBTHUNYg6hlb0EB6
nfhr3uUu44Ektc+6OFa6kDjBgCkbrMc4Cv6k2iRkTt1REOU1gMMpG9M7otwp
XQm0H5Mff+XpVRhlOKnU3TzZE6V2WG2ERWLUc9G8Gt8Lr9h+Q7i34V2RoINA
zuBspjRsBBMrEM5PhfYS/w4mdfInd7HJg5/gOjL+jCxS6wdwyLgPz+XsaB4d
kkQpIUA5jc+ymDyA21IM43IBWFuJtgtX8eXj4FdldgzUiOagwWQyq89UMEYI
2HoezRrqs66nd3EdUB+xIpmCQ74fddNoMJERy6bdZx7IGuGjuC6CL+5M6re3
C/wqWmVrmoMf4epD4HilwRtpccwBJH4ovTzdYi2DtNbAsefIXdv4OKhvw75j
yrX71Ufpz+2SjNPIQjOrXwoFtTqJ0GYQsbDUqQFLibxz+gTFkd1f7DhdN7FG
iA32gDSwloitWRWld/8m69NpkqD59GFnpgqamQtIhcMkZ5f3leuTR2cx83BQ
CekVjAW3cTK3unv9qhcgmy1k6xMOREYzJfe7VEyddrq0viGjOptsJWPGB/mx
ycknLbNjnaUB1mFFdLxVI1CERlvFsMCrYwV1oN4ZriOv7bsUNS8eMnYAos/V
3a1jkfQwztXmvY3GKxHKyYftOBW+17E/S+johbSBJ/2KdOlXHJu0bdqcvzW5
Qrxo/aD6qYK8ODhLLcdg8sBrY/kVebz65wkBw7D6hJmEElvlGefKnBiejzSn
5FqHT0bVU2GdarqQaguZ9UegzmhTB9yN4Vj+6aVzsnz94G2YxmHB4ETrB/tK
V406vKMg+xf9OHiay8ldoCYAsWig+RzVhlh1MXfvSC08P6iZVDzguBzOdsqf
BkejEbZr4MZwH0sN9ZWPDQHsNQ/WGJv5HlYaBBE6V1pQgBA5yTQg12PRpTz5
yjAmt1Lo/s0Gc8WcokYJnaKNE94ocSegk06Xj0ejhB63RGUPodVhkdt2U6dd
MHyo5Rx8vhkZicTb2Wkh+aR4nYgKgh1osoYPEdaimqrO/yI47Bo2CBCGHPDI
AJFGTLWfNnOO3YOC7Uc6dacExTIw8aAApRjjlPzfa/lpkE3O4CLkHoZibBFb
BKkiEzcwy9XKBWW8D95UkbkmlGCK95eNsZbYERfg2mbsrhCLC4nDs/01J9e/
HjxUXG6QVv9QOiDrbAlwEQPYy0izypgsM+4mITZjot8TXTeSMClklbRoVSo7
vwHjx5JrTI16WJ0yU1mLSAMYWN5PLMy4cFxT6R8mFeL4kJFhv7nZvk8z8h72
aRCq7KA/gAGs3F8jEpsoAsMrYSgItrsPkqz9aJJvFLos0TXIutMOKoNZL9aA
Ol/1AgyvVlFEiVOLFpaZ0Grv3GuPPTNNKJlgsiAxO80TpQgZIsvyvZCyhYWm
VQy9qt4DS7E4+b2a7SsiCCaQGBYZThMC1n4q3lPJVAbCBP8NkhWnTw7jQIrS
MsYl+t9O8EhrlQSN0eRW7n8VGpswvn2c//6IoUbGB9A/RnJAd1Ge6ldZgcBY
foXa6QPMCq5cEGMl/u93d0Db5UoU28Zw1aTj1z1L9z/LgTKvhbAh9GIhQCFi
5FglisTFQ672MwuTUYVl/NdVNEmVF5iz8JNZICEB5dPiOyFpkHOhHoqbktbV
aFsues5+nQnWpHwQw+epSdF8NB9VevErenP0xHafhzCSJoCBvtL38TUypek9
81jzKKEugQG6Oike/s4zHse/aHfleJ2h1MxyifKJNYPHoGXF+51eSLu257N8
Kfq7dICv/q8dYz2YsHK562PN8spHZ1ym60F5blDssGR+BJR/FN+K7/yvLswa
zP9OSGoul4z4OpX8hPFrlofGgIUj9fLgN/rzi4h9YN6i1RLMsqWumnQgcpFK
mKQx4HgdNC3UEVXcWVY61bPsKJGMOxQYMcgHSLhZdOZOZ4Fbuan9ml/DV37N
RgKVGE4qYOCetbTiVF2hRqKdE6uSP+NLbPC4giw08Ca0BUcBYRfWmhY4pfej
jAnsBR8+RxeUu3tlyqSjIjAPp+FITAU/PGmDZfmeHEYCRCmEnEIyCwEZw66l
H9sLMedCoksrlYN/RDA/GGhKarOHoTQIW9JlK6VG36hMoE1c5dPIkO2UXOjR
jmDPUvNITQOyDMKAW0E9vNrLgXb7nc7RIZsiEaBe6HFMbXuef56VSl8JReN+
ApJ8ta0UcaUnSEf0Vyp+Foor/NSqJHS+68jhH17F6EF6YyRzDWZUE+9j3J7P
XkQ8zVhGwoKOPJxPKsrctgC0qSmZ7X1Gf98nkU2S1cwaN6jThAgtk1s2jtEk
eNa8Yuom7hwTlQqV6fG0jwvAP+Wd3ihQErDl6XwlCABXDqXwUBsj/bAzb4Ck
MdqWC59GBH2leNAtamErivQ1lbaHVsWSC7RliVR8G90DHDKa4H/vtXQMJr8L
CSXagz5djW5eqDXJj0et5YcqLEvXTsWzo6MNKODtxWLdzeosYWfFh05dFU0h
gNv12wmLnI6ZvCCyLzk8S4cxJEEvNbawtwjQo2zXBuWnC0qgQTFsMPzyAvOp
o78qksw4BjROnnqkAfedqIU4zctBbw37qVdHsLgaN2/tlViL1Y4/LQSDGvpd
wPJQvFXuLLHMn8s7xv0eJYPZGLJrPm4da5mZhuNwTD15cySdiEhR/cJLTKBe
9prfMP8GAJZyzElQWyoaJV5TzsQ6loNTX5eOgVIPbHfvYQ9RB0Ua8thZAKLj
fNguzDYFPl8t2HScpinz84e1ChiUyYoCCSzJ1s/tsgPGVCuNXaNBh9a+mhte
wgIizDs0a+GTf3w5nmOb6vLGMopL9T+IWj7/N7oPMhHUy2mhk87At3fMaLZz
mpsvRwz6OC7Bgs07mz/2JrgXNViCO9odIRCzfzQsPygCBlm5+yg4xQDKwdrk
eYsV4sMTyALcK06+ULzSCGq89JBI3dauz0Ce4OCKb+6KNP3DCcAUU2jiNqmV
LQRtu23qwhcBRoWAqOEC/dWow1kWQ8JwdnbQike/JI6KewdT2yZl3o5AfuC8
2aU9LEN/HV0QelztY8kjExqnh+D9CGM4XoTjAhumxJg4fYENB3bSE6sfjOH0
/ylX0pmaZB6FjLXsT9QXPOgZqdCLux7AwOtyhtTXz9GAWZgJcQbXyj9u0Pgo
n9lcRegU9m124TsCQrbT4H4QAcs4uDtzRcElj0Kpp1idrCjtpI8QLmjHp4Y5
Ja8xPlhZwM0ac842tZru1N0tBbVMaucjp6V06Ajqc5wo+HUjzoSh0bdBfcLS
wM15hwh/AXT9oHGN3KKMpvMDjxyVsNYBVIFwE0LjvuyrVblqxbUAgpufW4sC
BRio/pzfBOF0ms0+opWlZ8BToNuYWzBRu2zj2lZgPqttgyhnIihNVHV8aE/W
kaWv4Js28eVrXvA4HxolHIXgJq8CscZq9fw8UhWkkk5pN5XCIBhx2eIShOF2
FAxWcyy4XC36LzqDyryDjnpJY85189ZPdtM9ilWAgDGmSzI4H3+UlzJrUpAt
PWRbxHkapTFnPDPjOMcjKLaCynHyaGOjx3C/fQLx7uxGR+pvWOd9Fodem+gT
QOxaNuTLY5e5rFTGO1Dom3KuBLsHqckTS67Ecukh3jqkYCCPIhZ+LKNESOLY
OGlUPUfZ+dDzkBuveLac3OJSRPr2X9O9L5OR6iMECURvE4cj99+F1fUNeXwj
j4MUMcS5o1HXgul3zMKMgfct5rgN+tLo/R1TZe0nXsfeag4tC4QdDYckDXJf
yVjLQiUpgS3gwTcFeLYceK3DFafsifn/d/wRGZLJPgcNCAGlR8f5YAU1iViL
u/4wtjxJXgkbeyxyBhskBoBy4op3NKiUbHXdrVsmd9U9Cz3DPerAo71pjzvd
YlK0jjUuWTgcbFmwbqHAVvWTIo7xYyl0D5q1WGYIuWNzU9L6K7URVuES+GQG
BD2h8gNBr8Z7CSHAIBLKsS62zjpR107zYjvi0OiSHqGMe8xESvSQzh6r3/0m
kqqdU7Ds1I48v0Rc/6pgjrPI3orAyvIjXfHatZQYtg021irt/0TLX0H7xn4C
MNmeuLPObs5lWPKf/9JHLw5i0dFcqljl/MMM1jY+10oh8LgyXOA7t65z2SlP
034OD7fNo5cgJ5ZoLG3NiWke7aYT3j8cCdpPeqhBlJ8NDM7lyen3Fa2FUUpe
crY+RI/HqvMCwExcZ34mii9dKjleK0hwXE9iykWWezQVDzkem0mSuRjmjomG
vk/1QR0xkary/4F7NvL1Wsj09t8urRsiaE+pv0wdAbQZsqhDzjL8mKFOxDio
sGi+OQAnyrZPotcaF0d5LuWA2PyJDUOpf4NH/0Zt1dAhjguWA8SJmUsnbD5m
NjAUZdbe7JqlvDAmFgY+yJnWOMYGVPvkpdR4aBeB9Vjfvv86F0+QXK5atnYH
6cASkCKkVeevtFbTNXWhfLy/3V14WpivLFBSdcIxdpG4lqulRxlz2pvR6g3k
6CqUU3n2N9CmWA5hEmrybK+km9nvg4skij5PHcUm8Dy9QTOdtUiEgcwEeuZ6
J2/XD0/XUQ8ryQzAi3hK74AHGkLVmpHNr+7YXlRzM4HW31NKTRRjklUcb7y1
5tM9MtA9OwAgdDRj1QDXSti75w33j9jAghnjv5wFF2giDfc+G4subdEirm0I
1w7qzsmX/uOi3PkvYIpvun/EuJAX4EIoLhcUUHxHGFXrfqUpViJKF8fk/vW0
rrMZFqM3NDoA+lGdOymJasEmTnPzIjQaNQdOW/Rr0ybVkat3/VsT1qqXmvQR
/sTuHTlaK1MXLA5IJO+cLt431abrleI1LRz1l7DAKGCFwftIZeIuTYGUucrR
/tHZ0ThdEeInuXYUn81d9jUZt6QjAo3ziC/pxx0Ies3LafhYLfPHZUPO/au1
uuWDgIBSwUE8e2Tz3Z6YVNr+843I7eUY/ZBdIhpgVRHeMQM5fM4F/onGj6Z+
AZbN0+ugMDRqbKjb/I5y3fAVq+ZADkZaNLupv2uz+K9hV+bY0u+Y6rdxxpwU
dkqgtZ04WFCURd7OOIHN9fA4sPa7vz184/xXMfiO9mbBH1X/hP1an41urKkW
J7/9EqQKAaSmdYwq/cOI+lbP4PZ35d77PsWjC+4b6Jo5r4ZX3mW1/7PyQHOK
JQpx4IdBJZhHgHtNoA9pBG0fAvbObgKyZayuuoz3YUwfkXGJ4Uue90UqNeuq
ZS8abtkqR99Zh/d4G9HF7Z0aBvrW5RTlE/0h+2p8HqJMcQYp2soVC97j3/UE
KDVBM+WZ+r0SQM9rk1RgGkeolX7BjByzQkn6xyUWFdX8oUIlPk+iRc5DRkIn
g0Pj7tYX9jlTk68/FueUeAD3Ae0y85Sm+dMuRS7zCr+3Fe9nUe2Bxyg4eY6Q
DD9tLOQgLmkbq3a1TvmObmTyPElYQmvCCH9SDexVClaooulYu4l67rL+fx9g
QLtEyW+bxkEzLmPr1HXcay7CTLAg52wWp98V43RdsoHbf52fI3HVpKj7L/rY
21DYiud3vziAhbqI7aD7j7feucVNCXFcWKb2n2xCGlI5qVLvnYg42GjRlyuC
xH6G6LS4kMqPcCsgODLqo7lvDhWdQ7GR4DMuv6dgP4zKLseKn9zkR2tSwWNE
PtQO9CrkyS1yApJG389KcL1uqP44Tgz1Rqa6Qb/+5dXZuCs9uBUVh8t75Ede
Zp7M2zdQz/jTI7nXB2pMQ9Evwe+sOla5lxbAs5Iq08HN6e79/LNK/sYqHvOr
Ljv4ejQL5G/FYPxqI58nE2MkXkBST4K/fxMZjuwrJUEqNIT+/gsZ519y6hLK
PixUB4RAU3VptH3SOa12M/zFEf1d116mCXUAxo113VG1g4Rj2thmopLGJtMA
MYtphY02D0PqxkJvX/l7dfEAQjypufOdEK/DdVqKEJTyj6v5j2BWoSjOhgqu
8ZC4eAtKJzp+zzzPS1PbUtOjsUseYd+ZJfAUOB9xVH17lUVsi/8wjWtwomLW
84leau65kz0f5O9h8JQ5bfGQkh/O++pkNbYWAIVU1kyLtwWX62doIEwhUEFJ
tyxM0PI0dGvQkdBV7dI3vlb0Ux6zNHpCHNEQDPkvHQe+0AcbNxCgvJrAToit
bWSPD2NHid8TXpX+jvakM/1hvegmTEX10yxKGWo0ks20+GDwo1CkNxSlXL6G
9QsxaMGX3ij3GFwlBrSbSbEtv9K85y3LOnE2/BNY8OShTcNkFUuij+Oz8HG1
yCsPrS6LT0ERV6C9LJuFFu4w2nS31E46qAeGlT2oQ+pdEd1hWKFQyv+XB1k7
IzzZrIJriInBmXq0+8j5S+wnXPgv7Qn6wS85mNKqLvz3crR6xYTfLayZ8cid
8U2xWRBYEXlBBc4rShwVbAAe2FP9/h0a4LpJf+c5qY3EjB8wXkHQ1BeL9OYi
QDKUlIYzyTgujo3drQvhbtpy1T5PEyMHHGuYGTEHw3Yj3Ru7L2IfupFHeUQn
+4WX3SinwtsVojJl94Bsv7/V/a0B4bx4vy29vOTkrgUVVluYsBN5ouEIznEZ
pyzngaxGORF/KKtZY+BsPgt1yiRqtdxvtDcyZr701jm84VQ46TwXkzfQDIqV
igxn2FoRKFGrUR+nPjpFsLfpc1GP/3JKrstn52TcIVlJZoQVNLCs+OYkt+rM
BO6ajZfctWogDSLgGVpQkN7gQPwBne0DBUOC2vlKoWx9poMlbWjUljL1VQqR
LZQUyCHSK3boN0chOjAxACmDYTBF+orqzq1p3Dys0E7nnqnhtnB9tBDQKkfP
QKNNqLZy743JgkX4adOy3dwGBuw+pHaCWyZNuRfYTFW+Hx608zVKSe0sqCGJ
kfSlBsEBFi1EZdhYyOr/DK71cagOXArH5uaD4Zpo/3z3xGTh5tQ7sOupry7y
19muFoeWSCs9wbYq1zEMZxY6g4oH7KG42QBgEkqtcPm8g5JFjmJI0uDIPaSp
TxEQL5QRL1nzlDtEFW3nSkKous7Q7GMwXEcSn+c5rbf4Gj0i2wK3AEoM9b7/
qKz7W666+h8weeU6B1UeN4mY565FezOfl4EdoTcLuybNVIzCyUA2wY+WmQQ3
54ESY2b1Yl1Qkp0mCNfdbMJeqB+2AoMbkf7/9GGajFZKnzDwBJKpkzTQpHhR
PVWqIfAEofZR9HixxBcm+lNn9F9dOj8OC3g3R964HrpXAtgOamwgnMZtacHX
bKcSka7Svhz9en2T4C1/QxdqPhINMf/RJHc89TcIfJ/D3GMDRJkeNJueklCa
GVD6B3dcjTqjFdokdaJeJek7L2AWTVId7lvVBpUMyWdq940jdcxi6NcRCy/f
gjj3BXvcWZQep0rl+DWnHKwls2p9d2ytNRRJPA3i1k3e4ZOju0bkl1kSHYkW
WKcawl6kF5DQAAnwFLs11hkM0SXEMLptYqAyJsyZbTFBBAhyC65CXg1XJZ+F
y8LR5QFEuJk32nMNAeEihNMhsPT0mZ0Sfwjj/65B+wxt2Cg5sVIK6jJIlLIK
UwsnJGYnzfxdIT9qMRhqdxxLYUN3BnNuw7olHzKTbpWfBHN5b61EjdEUUnSd
edynOjPIJIy7jtMWk4aBxrrmjVxIXFFnSmEs+I+bO1SzWFe9Ff96xJ40WZju
2hyNHQAHC1kNsdEijttJg2JZGB1Y1II+9Ohljt2DGrOCvebgrnBEzujVLijV
vjEmAcyBdi9Fn7bd2Jx2CXsfgEDvsKjJzfpXbv0BY3hqlvix5DNO1XZPAg4e
PmwUZPdKTn/ncHNEnxJsdMjM9bCl6NkEI3UEG1PMVn4PKu8Y0eQ1USs8Y6Ys
cnSX40frmed85As2Ik3OMqFkiZK03OJ9etKqGZ9vx2foFqqJmnxZ3niSFmmu
1E3dObUuJCPGaJ1CE5UwKsNZ4DId1gA78edHAE30C/5aOVaRbDMobwDvRp6J
oZcCmIyfkHMTK/ypdXbBVltDDhpUp1l0+Jhr4CVI24LstHDvjnrb7PWX7uVq
BCg/mQsYcpJDfqv+BG9E+CS7TYN8GbusNiR3hjdXGQVze2c9kmGOIkjRaNtz
rr2tVQwtDMONMl6HL5EtPh1oN9VdnEquJXHU879baFFeWH088FpyUBTlEnSi
TEFcYi3H8j9b/Ulmo3n+OeSok/iFb3fOuMNzrymKQBIXu3oFcktj3ng982Kw
MkplhiLXjHFDFci5Ulzr+jZRmxOG/RCeYCL0oSePoeeW4saxXoKKRt9iX9TA
T6YZciyt1SPwwzuLyzsT9aUdHk7rnjIK6nmG+PUTIClr1770+l1FfsBLBSVX
tPyiOARlWgKvTE68Y4jSQhhqBgjg/3FnNRprfne+OjsL6+z6/E0BvYVt0n0E
Z/izpgFgr5HlHH06ERMFm7krMehwfAZ5z5qyn31YXBK3akid9aiHiymoOP62
abaDvvxuVyWMJ0hOtsG3NzCXWFcvn8/eNo3uBM7bVPTQPpUMW3RphkR+kPJ/
gnkpMPT9wlkxbsFBjxpSe5cWCySoGDh/nAGCw43aUFzDm4+gzcOdKEWVwn4o
kbRIFeR6lbvQPDQ5ZpAgzp08/p5gliG6KKUy8eF5QUEKTvB1msotHRaKjYxG
57DyCGQqSsKHQkfYasEw9Ym+s2qTyYiTTbclpfpKthLXRWzDkcXxakD+Mx2e
GmDJMICqHOI+fWdEO319y1FTWHcr6pKhcZsJ5cqBXI3GV/oXPoNbe3TMZzQ+
ovy/as6eic0T8KapB4hRXpBiu2CjZAaB4oTQt+KDmw8M77+YJFm0Wyz2Z8mW
1nLtYOopKMgn3BR7ZtL4g1gv1mV/uq5AeCYHczMv08KFhibkTBUcY38M1f6q
KOH5twEqEDJs+yknSwzDPvkG6A7vz2s8f2iDlGzHI3FBXFOfq90kmzTVBL/t
BScyrx5fQA5suLzyZIpYvIF8dbDxav6BbuD7Rh/cdFV98hAqfseGtqEbcxls
FgdlBwiN9ORLKDBLEmwvej0KQ7FcrPvhKhlVEJrW/jRotF/F06HOaUkIqEk1
YGhYG2sa/CmzN9219eCKBFw6Mwz8Ni/sdk87x7BPs0BnPxM9lL6xHipWPA4I
Cew8UGXgSi1QCme5HzDe/I95MFqlvGt8XSv+Td5XrYeCAIr2H4Y2GrE/ZdFp
zBsO/AyhU2Ip3y9WriUkpU49Qa2atfOoPBk0DcXCCHN5L/f76oa3Pex/eHsQ
Y5+zTxAr6l/ko8LUhcxjx0VNHBarQxfDIqtlGROg5lPuyaACBvj75QTZEwcz
flRPFfFF9SkfU3j05Lgk6RcEY7XnPhbzVsxMYD6+7f87Ta1SoG1Ck1MP8BuA
LHOuLJbY4RHUj8Ibk3a5IOa7BGx4GaH74LPFE6RTk97aqqZ9s1ZDIeHlc+Xp
R2BOgJ+S9vOnBLyKjqrju5tjisvqkFerof+zsxuSfGwf+VJkVtyXUW46lgL6
GIt+klnOjUewbkYkES25e2ZWYvFxDJmR6mIyUwbBA/D5YgJn3nasxBmXIkKB
GZYI6R4FQ/4OKZ31dRoLFAHmJyOg5MkyqEtDvTUDAc2b8Lqk72FYQi4CHmOS
rME1+dxmaMR1ALHjEiFClAdSsfOLfwEl9X50Zz6x3ZzgICgaHvEVAFnrvSTa
8MYTABA/cpVIi7m7fRbELc3TNRUB3TXcEIMjmpN3GZy/AIIA58faUah6e8jD
fCu/jOmqGCqklkRhuiJgqewZNl55R98U78Bw4LUjiwn3maWI1LxE1J9cj0U1
LNKukrR2QBRMX76ylGNIfKkj95kDloxkk/QqxYkaU7hrqlUOM67yvCq6Ufp3
jX+fKMDLJAG7nBnHyfUxaRDt+E3w494tl7rm+Y06KC0tydE66Dm99rhHtp9p
A91pI+NpWP6kpmeQoQtRvjg3trantLFxWvQOQaHkUpRkvMQEOAYDyBfF/xc3
9MyKdbogJ4XB4Mlxuy1x8ZzSKsAcOszvs83Igj7v5o20Xd2/GObfEGXy8aNb
E5Oga1oH38e2KNsgtMKIWND6aWazvIKfEGcRJLeY+93JZsibjrm1hdt0EgBt
qTaZkIe8U6rL1Yd241qQu8LuTKYtg0WWoIjZU1ocit+ZdehoDkiekQi3eBSK
ojZIG0EupVezBBUeKLDJzSunOame16xFBY0XFi8Y3E9hfviaEgcf5iHl9bLY
HfgWtrMkNZU6oX6JBvf6LlqrAsAmemJdRL4iBc84lOrBvCKkPO1w9Tr6z0Tq
Q/8iWsKWhelS+yf3risCjnAp9hmklsqrMGOEg9yVBGXi7jq0HHYfJ2nZtEGP
zKSB/gUmemFgKSHlYO7exuX/Xs+HLgeiZPAZhKYseCq5hkqgW+Hr8x0sQTS2
xzEHy0VFBqNyFOQhtMTL07umOEAesiVXMUBDxP1Xv1FSpY8fswlrAcGoM6jI
s/fmeJxD+Ay0s14kcsCaeUNF8VjNVE1CfG4H+c+YZYYl/Ejd5O6QzWV1trCc
PZL0WriMI/82jYyFopDQuOZ4xpkFD07R/jlrkP1Fx283OZcaVvasABLVvDgF
eI7V7twFstUvg84ejEa/mgedF2IqSrkTtixsYJOHzmtaNtDlRnwRgmBUreOI
/AnvLWvt7l+XbEgi6QgfIwo5cZ079hEcIRXmN3zBdSq5i4KH80b7FRpl/p0j
x1GHCfMAZb0gkQ/Bn+B17X4R3dnRQA/Yfo/f/eYQu//y5u3bzqzTYX87UHgg
fFMmGj9tYUCug/cWDGAYI4OSoE3k5gDRAs3aDGV2uohUCVFmtDCc5U17uHlL
syA4s5BjpEFluAoMubt+sqg2VLtJY6tZk8V2IKHF8AA9PoaApFKKPDxEmJVr
y2/HDEFxit+0iiwE/UCc5xLeo5Ic6IUS83N7YmBx0r7vgvf6pfaftGH9Y2I4
UVwCvIU1wBaSfrmya6e4f6qnF3O7/0iwk0ODYmK+rCsP1gxU3RXgy8NN49f6
UN2I/LNME5MJyFLZjsNFOyh4iY4krRl7BqK0TYiWOBN6J+jsW4KROjznLPGe
Rk0HYPpXrH9+laNRI+7j2nSm1NHOWvNsoK32Od9ofxMIrwgUI9k+GJv+l3XC
mfBBue+jmKTlarohF42rAz952YocFWiGe9KY31oTDO31zXGHmorn4p4EfPUt
6Wabzjytb3wDeX7dOwXVs8oLeImnd3Jb/Q4vHrtbQ1FK9SlpcXwtZiUHJegl
D/vlwVil/7RVGpQMZ4lkuZ/CodpJUTXyujRugRm44ihKR7YJbaSiTQDLqyOZ
dGIAVaLSxutCQyAP7ijsUFworBfYxHFU8cDJNMATTlJoOX1ch4hkGgoR0mEG
oIt3y49X3KnVkFpb03gjXhQTCM7qo7sfQTFpPikewEeJIJq56lnP7qY1cz9/
PJXf8Vwl73eUtMPWtSWOcVKyrkIZ5B558gkpI9q6iSvlG/Mqglao9mGGqc2I
Mn+HNy5XW6+xc1eRatpXWzh2GzwcND5EUdtm7ZkUJ1FDT2Jm3zWaoPl+lZ2F
uugEpZNEQtAblnw1tBO3lNtqKyGHG4DcbgIUysItuFsOrJAtlzkjj+KgaI6z
git8FDnUxXOQxBxqZ+FbmnqZViRkf7Dpx7ZrFdN1qIHre+xbLEwews4EtNOE
FJ7Nu3o0dsMcalEM1HezAkjGLmUU51h2Y92Jj8x8KepI8ADpoye6U0jkfSXr
woPqlDysDzsEt3FtDxxd2S5zGkqPWvVczxZdPbEvuUmxFDsoGJjz/BNIcAXB
X6WyxHbwYTsThQwzhodlXn4AvVt+z6S+Gg72ZSoiQCLywNh3s2xn4Q6G2Kl2
lxFgR2g+mnJDppM6tnlyXL6JcfgRF/t6mnh9BwisX8UCWblkv7Vb6D7I8M9S
7AcDdRJuivjhFh6ixUsmpLqI0SV5rzHceSO40o83D5bUc1/j5SBPgQi3+ace
RdslXX9wMyiNeEnEYi3eEege3nFZmEkRM76VSBQK7AF7JLlCYhV7X6adQhbE
aktKPOlWUdCcGskvTGzNAEHbwPbrb6I4+j8Og0xlOMjGG0deSJNSb+DY7mHe
of965NHEpcupa+b5BlP433FSKHEpdh9hNI2t9bQn867PPeomlgCFQWKuoTZW
XL8WdPyRf7klX8Z81CcLAKZL8Z3SXqcBuCXQRi9W77AcddUuAgyvVhZcd1Cm
RlKDOUEcdNyxvAHOM+r7ZEuKk8Nt6PDGAWZ54C6mNk9ym4Ailyxe7XJB01gH
y8OFrWyJFgcEJvvLfrbB5XLAmdnpgFn1P3mysJGyLpiSys1wC70EtF4YYD87
QALM8FMry7BDsoPIgNCJnvUhRLApoxjJYhbVsgehaxhWHgQy8dnsQHoU97bE
+r8+CdJyeOG2Ef/LmQPmUJLPlSHGkqYU7gh8m7wxPaC66wPGoUqqxPI2NIb0
31+Al7YZVkcKjUmzd5CPNnutBf2c3iR7j7KUDNByueF9nbHYZh4E4g1HHPwZ
hdC8Muvm/lDSnmkLJ+Rd5mV9U71kDgtwM1DEiwnUAcvWKY6I1ckZfSQwYHm2
QP/uMnofIvJas+Xhb+p09jqkMQkvQktqRlR4zYILQ/6pUMWTWmQqwB3h8zib
DYlEAoUAXhRiTyumUHXjkRpv51lgq8GI5EysQl1RiR/tu08FVaPEf3Cu1pkt
ccD17wRddq9KNsmVKPdSeoCiqM1sUE3gMhItObhgqlGnmrYS19h0eu3Oi2f5
o/4GtdnM7Motewzmd06yBCnHuHnQOh5h2oYeIS65gKGc2mMWEFGlrusdg5HJ
AJxWA9mMjbG6f4QMOF6OjfRJTm19jGw+cpVKOnTicVoBzM/s9HUsfZR6GrDX
UahfbaEJJEY7FRPBq7B+93AKSyZb932AVkZHLXgozWhqLy2A3EWllXByQiSN
QjzjknT4D00OJfmozwqxZceDH9Qv23iZHkEoj0lKm77FKHYnbWO8Yn5H8sPa
iQPu0iH/RbOC1PI7Bewjf9wJ2k2v6wPT87J1/AKiTrQka65mh2xMifz6zBr0
PoPgIHgml563CHztjmBY5XHxDaZziRc1dxmY8JUHCAX9ykYac17LWLJvm89j
KOv4bXOLQYB14g6M6p8hZfOx10duuZcvlWEtOHctd/vKplkM0ZuF8eXSWx75
zlofWCOzKqgujNRbOReioK5HBGrPuzvbotx5YCsxdGkHpjH//aP0fCu62dhj
uler+P6aawn/PWW29hABuLsAZ9iM8xLwA0CF0cicLC/GxT5F6QLaLPh235wn
jLWjXcZFFBCSZ+qVO7Rnz0Np4YjKmERLgevcPFeKTxJfWa219cl+ZT1OnL6g
IzL/QZZybnzN25lpW57Ritf0TSbU/J0rPRnY2xZXp0EcWhCp16ZAf6JMjws+
FlYCZ8hYplTEC/rXX0QU5viNMzL/4uUlIG3eLil/1P/UFmSe5GnKK2SAyHI3
RcQkgsASDkrak3hbvKw4ETWKVe1NLS2MDeKW55wgeR4kbFdx6Mfq1tXTNdGv
nt5tE1ubiywUrcdJ+jl26Fh56z3eO5UtMeucvmEh6O09bFce+8G31NQGmsVW
o5OQEZBUuvhVI5kLds89zHM+p2rUMjA19vBXYX0MqG2xLZBOuobZOWL1vHRU
pg8vLhAyzw8VpCwFTcqmLcxJzOvjYGZWsbsOs9OaF31BvVPQ73fejP5YnDaV
Y0O/lYyhnGuiX00lZdC4/28uVcURwj2t/otzjvkTOdyHiltkE0yovNQqOgjm
QCNxmyVGHxPbWOwHz36BCapsNRRfO8jG0ClB2imJXifsrNkVgg+GOfKfwsNu
3vgUeQfogYAddx1OatqObMXN5FjYeV/YJUnDyi+Q9lN/kCTRN6RcUDuGh5JS
gqZaoUT5qxN4Q0H8j5TQntlpbsOBD/po3gmI4i5wS+z75Lc/HtEfkMLdudkX
WiuyAgB088F7erRERmUp66JnhaRGeZ8awwedxyWE8wcVABYPuNH3bj6WMN8W
sKqbl7xBmQ8ayOcTGDex0QlvSKukwPr1v4AB02JaZEP8fiup9gHMkDZfxrya
UcMzkb9iGlJA9iZ87jnLndaTtZT9o8UrbWrAWbOEAbsjxxSznUaOmPRnQpBY
P+OO4OgG6jHJmar79QQ5TPbmPqyMraPiqj982qKzyV4zJMF/nX12ROqbBa6x
xMTNnkbH1VIpJT9d7/QNy8Nr3oLZEQu7rZ62tfmSbRHRqHCS+vuW8hOQkb+4
kMJqwYKY5A/5CzvNpETpkDfoaSTTuW2wz2TkZhc1B0qjaNaMLaP9HIku/pqG
ZqLO0YVt8AKW6c7yx/l6fCoGcEnRU73bZeLR0EY0Pl/4Pt+pTvTsaIwlPXwv
agOeuXs5UlMix4tiIFMc6VRoBuaBGMcrZ8MypjlM25u88tSQn36BpiQ6ZByb
dU9fxD9WZkEX7rr7R5Se4gCGqSSrfhfnwxUtFWglADTAi6DVrkOKBUVEZaNW
NE+ZYTAL2i2NuRFhe0GysMSuTazxO7AiyzIXXqw1pyx3egsaoP5wOPjtLu2d
Yik7ouRPhPRcRM5PI75oTlA3pct/iE694OLUNbbA3fwoLzYpnIQBWkD4evRn
osgffd2YfHu3E/sGEtRVRZIvMIYpkb1RSXpSpbkKpjrldgZYI4YVKgQetRAh
PcPexqteABmAF0HM9FW/Me9+3gUaWrz60MSMpx2Za3yRnlYXWbj4QItdID4Y
O7+bSpBquOmha/ZU7+x+EBMCyDnqK5pNKfAqD4xC9p+oKPPR9tuJOmgXQl5i
b0k3TleFDBQmko42AD5sRa3pxhDkJTmWbzOB1FyUqpB+5rAurFXKpjonatvW
pmvKWAvPrkggXm6toWIbKn4KXGyUmJ+nn4n3olR/Lf11EjvdB7IhqkLHxmki
wFIRZmoiE9NqQMWD+5pnoop1fsQ6w4RgAcMOib+B+Ns1xDqERimOj/BRD93Q
iGwnni0I1IaN61bIPZ79gj4zjcgr5E0LIn/l3wGYdu5oOQpkuOehaGj9pRNa
9RsuhfwAT6ZY47dnVqyJHsZOLbYIok3C1MTpGvsnwW8e6uwp44DGV4MPGF7+
/GzGn9zNUXA94bAvvT7hTTD5Lcw0Pl+rCPv6wZglQmFot+LWt7ulJCLL4856
h1htfq+1yQap3Mdd0eKFK9U1Rns/jKEk7Sc9wQNYoS/m7fJRMVDnTzBrTEFR
u6AsEHPz/JrxjGatXMgaEM9LnAmN/fm0vcOPblC4wQ3IU1EkSKeW5m+qE1Fp
mdxLcPVTpzNhXYjVUWuNhNkEPJ7roGUf8sMAnktfngTA0mFu1NLDqKCvwr3V
viP6eKRF8LsDxMV0roLUfisqMK+4YkwD5NqStqGd9iv3Eg4CTUyz1ul13zui
ZNWppotwjWtBF5Uo6OXbOD+5FcP7I/C9XBC6zSKEt6l0BNoJpitG+PxKMcJv
BK/1r7YVbClEOwRnT1ff87JrRZY2XlfqLT3jmoBLt1mFmEJC9zlG93xaBrqO
370hyC8xp1H5FYzOAay+eb8WCKrvkuIV4f0WPm5EI2fzHmlmbSvKiv1KQJyH
JrEfWkvX9HjtzJKCfTKIGEIWe6Fz4APisnM4oYG8UO3OAZyOsK1YBWN50EhK
/cj1POcIzdTwllHeMRWSb+lNpcwDXP/Hw4dw5GAfUFvRqCdMAd9gj8nYao3/
rT73+TkcL1Qz/jFvWTnxEBDQ7BX7ToXdCY6TjTw74i8HyE0zCCPcPBpkwXGu
2CLanUUVGrr6xBzWK9vI5r848SbN0pYXcy3mTfkmzdkumP1dlwC1+mBiogWL
tPYBMmAax2sG0gKtOI13W26aM373ANbj62vO4SFB9VdCC0ZxpZEp8WMWxnRU
S26tl5n6iiVmRRJ4JHj/oWAaqniNXsPjQLHjPiwZlkI1b+Y/Q6kCXw4g7OC/
WGSXVf1tdOTwqKAweHyDxb6LA2mj0kgYmhKGmaK6++cpmdAJ2k4K6lybA1dW
bzs+RoS4P/h9z54KFsB1twYn4sVLFJwgEhESd+ojulV8ht8BJzA3+73qRh5I
DJhrRSZYifN+cTHnJ21weO32cy2QsnI+XDdvWhUWuPIB8QBxU8okvNBvM525
JyHcuhb12CCO2yWrSpR6CluThELzP072B1Ve0f02rJcrHRMR+afAjkSXCFeR
cTsPI+PO+QAIsyVHE8Ch6Ebr6YyvilB2myS7KsL9Y4aaR/Q8A3W0OEI0Fn/Q
qv2I+d00R5eYqDt7giDjqxuYW0HDTBwSQC72X+Dk0Mq1xsWQqS4VwIz19PEa
H/aM28eidR+wWB9OBHX9/dTeEkwNbT5A5vdQVPgP/h3kmB1UYutrNMcklSmf
Krk2nGB21RtMrgP4gjTP8BveYvaJLJMQquXDUlyuXMBArIz1iiifXwhBoK4c
+UWsQ4KeQA+kf+U9fNRYsGTzl/ZVxDQitWbfYV6ETMkQ9gaYe8U8mXr5VkIi
/El494m+DzX3CnWAYtepu5XBaEmcFA09TVeaoZ8Lixs+LLOwWnp/x4wEJeBt
UYM8Do8WzkZSXg2U6LMfZoSdAZtePGHmHOiWoaslQVSvrokvNBEd/Fk3e4qA
GA7Sw+gDrVZE8lXy9S34sRtAF1eWw/psyNlMJ8FvlA5VzkjeepG2MU8uePIz
fZz6JQXPilFydDyK6xSXFYflt9bitnELIwUcGv7tAczxMxDE9n5YI4eoe9za
9giPJXT5QYt9GAdlxEtXHPFBVHzF22UutZuUrY+winUuYGwA0x9lykheU/Js
IeUreMD73MDYPOFScD2yjISNrgqTtajX0wwmU1eUGhZEb9haG4QttaqojVfO
m5iG+cyqLUlrpxGM0Aq7hLPp3ykBDvdHchEthHOOJqaTnEcSzCmRpiKYagqy
PWxbrzU4ZJjB8T0uBdwuY7m8rIys4DQdEsMH8wVEMQR+IToo0lWKqRH754yR
TPOuFW2RSKrHoRl5Q5e5GrCMjgLu7VsliX3P4wKBT8WYj4pTxbmGcPJHPN+Z
KxRpnDMfZaZlonQbx2P2A3YBKA==

`pragma protect end_protected
