// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vnSl4DyjT0UORv3pV1sySNepveU9XacXj82Vfm//uOrEuie/YPvsTMeWWUBz
Ao3ZGibRe7M286tC2smEI6z9IDBQqVV9qt8/+yO3JHckF+dTUrT1Gdk/nLBL
ZUzzjkQClBTnXZSmzJijCX9vcbAarndiIU78Fmv/Dzb8KrUvHjvcclaj5HzK
UiAekf+UCwgKgpDlKdk4PJ4yaHbceXA0SemRFc3gXpMp0jcc1yiUW2PdSjJ8
Lfo5jrSa8hwz/+uYtXKPtteklzDzllkRnNtLPa75tV0rpYqHfwFF/CpmOmAM
jn7SL1NAZ4qJZtCrzy+I027VbNzK8J3gpuToCwGwfA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jn/g06YYHDKI1pJGkVkW3esyDByi2FQRpYF7pDIzmbHjItAdgA0bQ/ofXW2Z
ksgCrxttyeX35FqxexYXFPO+Im/xJpEkZVKKDU76JKomm3tqaihmIjQPToGV
RTOw1e3AtXpvEPkt+7LOtP9JiHvCQj/aH6ZJnw3TZzd3t7Q5XK40nUvTxyEN
NX2fjNPfGeVJKIn4b27O8Lt90xnIDs1Ca972ZMkVD7uh3/FI9FNDtLENNTkj
oj/f6W7IrGJBV7Fzbm3kMhYQzY1L2ieRYxOF5cRxOd95Hzxv8QW7Z6Quqs+E
2qVoNoeFDAJ1f+2MjgqzEScgifqD5Yo8gZIZJwyyLg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gK6PO8bVHJ4HT+HoH3cEUzE/R5LVrc7LV/LMGHR2fUM++Yu/PQcFm5vVr5WP
wINAZMwFGDt2vpp4XppobyherHo43bpRoQyF8ygoug4lQUiZGUlI65lrkhU7
ALUEHas0lFEwI8sthHcHE249cJmIcC8MlJVcKiBJoWVmHPEeQ9e8bfiqOaFN
bFmwboJbIWUHSHA3gn5gJLVDbhGKyRhXv7jc87h6QZXybbOamAF6GokJHIrH
8AtoWBRlNZC7Bq5yL+YcuQKV/tpzHs2nfwzix1N8VhauKggr3qlTg411PK6F
krlySrD54bKcYcgBscBgwTfXpTDQgas8TfQKOIH3sA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IZPX+sdJtkzTF695J0Dd5aN0lf3KSmow/+IIkQ6pp5uWf/iWqe4iYPVT2Sx+
R6KtApBaIbtzj5j4m83ompO/31cqjQy/r3qX8pRrpNjbj2sfYkjtjIBeQGAi
RnqEJqyHiiYEG2bo/2mIBiLPe/0moPncpIExAJ4WsVXbgU7tlC0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Y+x/U17qY1f5/N7fVU1gGs9+DnVPEKEUpM1LvTW4kwPyUDlJtX47mDmoFVU+
v7w/6kjRNH/6Buk/wpdYrOI57NIEoNyu1yaMKQAHRKt1oWl00qMFS31dZ3m2
Fco/Oz184rmj33d+cxVDts5L+Jfq5ln8FyMewu3Vu5jhimgBTM2RQCMhQgtP
RPqjJlheXcqkHj3HJJaftNZTefgcCgIlxWlYizIg/m/xOvITNJsOkE3PQLj/
5AP8rmSu70IuvYi1ZQWeWM+StsCIkJ+mIxkBxBj81v7dM2orDC6Jkv8PsE+g
tOE1Oe8wT9Uyro81/MttzqDKRh4Oz9Kp/3pNFK9lCSpj0F68+vLji/Xp1HxH
/ZXeaa7ZHd+b4jb71+lt3VQBXel86DAgM4Te3OOX1xfnaCqsAG4m4h81n7Dz
N/KBJ/MORy4jaA4Uoxnd5G/nszjV7aIodhGTjL8PsKlTK77UTZPpz2Fb+rge
GWvMcdRStnEhzHEyk9io9HuNrR8xDrU1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tS0642kCHaodMRPgpjQYanGd7YiV71LHAgFKSAtCsua0iBYDzZABnevXv7Ur
WTNNo5wwbPWiFQWP/uEHQjCon7wzDkzdh2wNZsMEO9oxrVKo7EiMmaIL5dgE
rWSDUxT2MpPQAIO1W2wV1CgSNoTALiRiA0kJbcQGFxmBjkpz7/o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VRliduI9ZxDJUOsotYX3jKc9qHcObtg5vsQK2k5DmWWYX6/Rb11fRfU+kLQX
X/OS+zGKke8PO9WDd6bV9A76YYYnZCrodAjxRWqqSC4OgMWnR5PN1qBOizAw
ElwUTghNEZukbpMAqQ0duzUZXeMbU8ManWM84DzKDVvdXbM4fpc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6864)
`pragma protect data_block
27ITELGK7Qw6qnohkd6lvjhDlKGPN4Ovokth9Cd8lY95eHPyUzZTYvfnPIkd
eErvtcbrfB8m3g40pUKBEvhn/c1Wm7eBXuUcwWw+GD5fioOLF8ewA5BISLlP
u7JCIad2VSYQr4IND6+tbj1CWqvRA2oYX7JQRmaz7oKHkIv613MsBmdBnKTj
8OVoJaJGT5h3+XV9oJViZRULzShK/DLqNXFCD4TvUqYZ2RBie9eXbC/b9Fgl
3Ta8eeH23Fq4x1Q0iylIRKH+auzadgD9DvJiPzamWA7/0HvQnfFwh8cOCUqN
5cXMqsnv97LCXKsKHYbZ1elAum8us+tBsNJ+nBe1aPP+0GasaGIfKTzTVb0U
VfR+35V8AHi4rQDbqIiJGcK5qGpHhKz3WsXfqj9gLAfc5I602+yclilUSEPy
162QfFJb0Y1CoUXf8q1d//ANQQJtB10DqD0hADtZKWV98g6G0ZVnd776laCt
hqVjNmHKeag7ciAtRm9ii+DHS3F/0GhRYbzrUKKNYMjdwaLcQdfj7pLV4A5f
+WKjC3eQVE4i8cIKOUPbR3j2ZOcr0XHkmHQxa86d0XBzYGaSAsftD8IJmCcD
BV6PJrQVulaJ2kwGWnIKuTv8sNcy2k9tCwfSX0Ii3cyYmDNRLTCIMhhcI1Rg
HYGAwX/FiIs5Bs4pFJHmCtJL9g7uXFtA+03pmLB5ukRI7Ra63nwysQb6KmYH
I6sgVYKpfDLtmRxGhSgeFCXZovwyIBV7/+fPVqPI8jcCeA/fMDBcaoiCqtvK
NuhYXh/zdyuTwHR+Y5l/0yC9z+kihcvTGvD2hpeRvFr53cartfdWwShtZsoQ
Lo4pWu4D1vT1UwCLOx0g3OMPqiHP6U+Gfskew0XmWZ0Dr63abt7STBhJgAm9
PMw9lakr4GSE0uKbC7jzsfjf+q+SobDaozK7ztlM3KNW8IXCDFC25IQmPd/x
RDyhf0SbI77WK1HzpJ3mbXck4TvzFnhsU/ZQgxDtx4LrewCUtGd06Px6MxRW
OdiIO/1sPz0qlgQBv8JB2Kc+J9rc2uB8NuAKNJVxwXoq1ozFd4/xRTii5j+O
og3pdSYP+AAv4Ih2nIiN2T/L6w/R5uPQKD6zk1llGXvs5fXlqoDGxPhlEnS0
03VbiHTr9VHfdjSwsQz2I5WLjaYtk13pcmEOEb6AlEvJ31zk8QMFMVA/sKQC
Chjw/rjRtLAyP7x99PV31AU0NMmZ7SdkpEoCQ7jdgcv1nSQLf1/M5rByIoIG
pJ/330K8Cz2pUcsml8CSWQ4mqWVBPVPekRTJ1VtcbBpPPuSTyk/Mpgn9eD/6
jm4Ek27xc0of+BgTE+peG9Q4wEBIb1MlSHFJH/tRpUheX5NAbkXeTSTPvMjA
Cl9kpdAVlGttBlWGoZemtv66boAZNHkwSG8BfZVCACtBzT/b1FbBcqPKWgr4
5YANy6j+w2LL/ft9oJ7CIuRwTgOR6vGmwpBPZhhV40pVodFc7Fnemo5gy5Po
816p9mfpYZWkFts40NWB/F80oE/ZMkWObiE5abweg52ibe3O6g6xTwRdngwF
IkKW+KUFOkaecHwduSSb8osKuDrFU+GQX+txFHHBnecFOKJlfd+O9e+3GvxK
ZXkh5wpYseTLFbVZdEY+vXA58I78u0d7my5LSu3Ls/RbndAY4pI5CKmsuMzH
cQZ7WaKob7PHKuHlSlt/EQaJoyrev8MU2jNzD/pk2Xp0Q723VtiN8FlHMm6M
HfDcIS/KFUr8boGTYHofd5rM3M+/I0pryckJYcMy1WTLflcVrsZkhZzDX35m
9uPDZ/tdRgX0RGd/isjS2BkkC+CyrPjfMiHKMbxKojmbnQOtMdaACNJEKOi5
7bVUzxfB19P17EbuxXqWIDcSxPEDZUQGm15Wkz5ebgDdw+I9n0f7r58PYIDw
DXvNZZgzBHQ4Tlpt9hl0YujfDj4bg8hhj3eouot1QjEqI4aaHETT4IqzrSNc
LnRm8lTdseei+bIyE9EKPIljdiLHugHKqTjWoyZdRwnogC6l8aaVUSIf9LoN
dlGlUnSmr0p24WGoT328hAss3NCf6o6bx9vdT/tK6UhoEiwvf/h0Fo0izj2o
w3lz9nxx9N94dZo3pHll1wj+/coaM65wp9uV5er2rfY47N4cRopyG83I0zu3
sI3tnBFAZnahisBQdChy8lOwob0qufCAKWyG6UWj6Sdd+6IEN948FawLBGoj
LBVWbk+YyCtbbt4+aY1BaCTB1Zi9e9E7wwnNwN8q1hDSnwE7NnW13Ys2TZbt
NhR3tZII3lKGaxsdG5+w55gvPiKKyeTmDbAvC5yy1W4/GM0zjC2cNq8L2zJn
Kxw4PoOautZxDlSngs2g8E+Vi/Ss9J1LQKwjBOcTXbjbfPjMX98OaYNlYgiX
BvcTLqdAfKAuQybIFNUzI6vQ9AIA05Y7SGCLDQ8YCf3LCBnUUPpJBpUaAuP/
o/FtHg9mzZpYdkTZHE0AEam1UUjHm2NmLGOILoz70+y52OeKM3boTWolP92y
BpzjdWQj6lZERmEOiQNRQOFwwqbxdx+vvduRfgZYCvc8YmfFz09qzK/lhbPd
VCTLsX9wuV82TOgqXM5BwqxdEzXMK+XGafXRDVdILbQFuTBy00CZtheLy8xA
KhfyfrIiGoViFEppoCyIq4hGcyZUxj6E2+YLZaaHfOJ6VJBOKSBPCH6fZV+d
3eUW0bVZgPKp13Yc0Bu+NKQaEOOVjwDkiLkyxCPguMB6TS/dPHCIdcwjIXBa
0Bnx37Ct0RLWMkYtuXIzSLSdKI1WgIlXA4yKQmy6EHJ0w6JlSDGkbNBjgP8U
DfeJP5demyfAyh4JEql6tv1glInh7Go7xAivgob/tmGFmO8FnTUWXJqG4Y1c
PJvhtQPTxipOdHxRGDhZ5WDgoQyRe1cK3RWJBPUViL/yWmmvqxgrJFv+Emfj
BL69HGz+yA6XzQBKzDKwJJK4m8Wk3S/b3+pg/cA9xlNxpQvD2KYtzur2a91h
byu9pXEEVlDvlGej9R4Ein7R47D1k0Hkz4BJoXagXNJ1X5k0d+Rx7GsTMSqe
x0nrh+pmp+mGxXCoNUQRGQYbXA85S3wddWA2tiRvoxaDNlD2MueAcTngXCIv
0fPBCaJWNesElS6I7pSVHGfwEnHsP20Fh69Pd2jDuln58HSAHwXQiZSJCaJ7
umUrgJE+o6mDV6htwpX3piBh8AJeZoHJnUvLxjB8EblOmUjd6RfRqfKKhiD8
++f1qWRKidLipKCo2RCHd60Q3i/kCHLijtln5C+EzslI7q2g4criD4GDSrXl
vedwvGcYB0E2gPMmIjxyibaMohqaNAE5IGwW2i7OWhqL8kzU4pn6VWfYAzaX
K6Xe2hMqNdEOxVUKw2NUfW9Txcec3Sg+DRqFMs3q8vU9QgqQC3A+qA6H4qeq
oqYf21n3LupjuJlxwRnylbF6JoxH/D8qFji3iBRfWvTAeykrsH87ZkuSIsi6
RsAzNTLDiLYP7a3PEYwHDJGO4X8uzp/6JGHypiCT55UBi/ZEEbhfxEfqhA8B
DsqjUS4tN8StBoBqspNNY/auCVICcxna2x8jgs+bGL2v/eXDefUFw+btEF4y
akqbbHzprAslWOL3O4px8aAbmZZAlSzxHCwcZyDjuHcejPRznEtZbwUktAxo
32/x2nPUGFBxS6HjMde/zeq/nrPcIL1im9Q6rxNzw8SFchX7WUkzwpLkQXVF
EREdZYqJbZ9U2w3WqFjNXf95gKb07GdOrJo8pLxUiHOOcqlGjmQN7iho1ijq
wZ2eGkckDSJJqhh+qvmiqvMWFuxFM8qOSj9QfONe6RINcvOb8CAxsmIlCVgS
criPj8B57iTdBwL7U7lwydeG7jC3yJfMVlTwnlpNRRNdM/L9/zZyAybLviq5
9IPOm7ScnsK5ftVt6QMFUubO7aozcxivjFETsup60lDkXrtBuQLNbtOyMgsW
fQOX7uUm23DxmwO+FkdNyT3Sk0VkhXIUCI2wWiV2kH6fNLkIigOg/IcA4RW6
7zVKxz3FQQkmxfRZn3vYRfVz1vVFPukbSpYCzYr0/1qL7C4TJ1XEtLb7f5s5
fbSZU7owjWLxJM8AVf/LyxchBEaLlhGXHj1hLFFomTebiAgIqO0qxzRhTSA1
FP2cnHW57Ks7i/h24dPpUbm9T18104l/UBTTqMht126PrCiPMeDlBT+AiBZB
8JO+A3pNLyIeG97wT4vDkB7WPHwT2zhY+L1zNuU8X64X08cAnxL016E9UCRc
r3pxs7LSrq0g3S0DwYk3YGFcoz+Tc4rnOmfxSk1Ey8bk/90tuMwko2A0McQi
kx8whYtK+HH/XQfRCtyo3/z26XZW9VHmScBhiRXuHp8BfvmE/wc0Exng4h/F
hQSKSxvI/N+Yn3oBeNEZ2x6cgnwiAqEeUoZtw4UBiXv/xUC69iNfkUNyQUDN
Q9vKTum2EXkiCOrKzG1qKPOK1eQcXSGFBJ/1LV6KKXbEITfyX85D35949Oos
JhNOa5DaZuKpYnZcUIAo4z+Vs6e6+FP4LnzNqm8crRATvT3P0vOPuW+czI4A
09wFERIFPirJeY/330bkkZCNbWgUFtUMOMo+10+DMH6t0nZYp56o3H9WroSM
j5FOL0Zy6EBeRSUAfusW5DnoZd1DkPmuU0hz5jTuFhqM7M83/vt8QCUcKMXw
mbNFjI0KdfFAI9sf10LokDmoFAnKuT7syvoCNvKS+O7YRTYYAn48UpxevKu+
clFfHp6/Ak+c1WbHpJJ0fYGqk5KyBqVWNWk6jW1WG9Rh6gJTf9HaMxsMWgRN
mqFFxomYnyv+VAgCGx/eSCm1/WwZ6WQ1uAfBXyzWUBgidoqZ4wzpDeAHqKDl
4XwGw3l0qk+w/0aMeuLBaldrSnbjG+8GaTF4d8fv+DiBCiRb5uFhkOFmqJX3
RAVQyfA2uzwLK/XqmQHsVtOJvHyViw2ct85vwtxBqGuQyNqzQF+87pM1ArhG
TtwjnkjGh2P679Tao4Qdl9oEFumnGpFut+s14zt6hx0TM11dc96dZ5bNSIVt
GrSkakSTO71lgQ2x8Zb8zlFy/qdzlR000CXkSBtx9iLzck/eoxH1V4ovs4vd
qSiTXmXFNCDmmbyKk5D6NKxX8blelp6QK+4DNkbDzamLXtycJUBarcCwe4C5
2Uk48VhzuQeiZkpj+VUR6tZBR+oNxAFSMg1ljzqLp8HXUyILxd4gj9wYoU3L
IH/QNS0LCj0eIVfVCTsq/XlIpSu2fZ+VVWCKMuWv++EeqV0u2ev7TqCj3Lvu
14FCCLJy/l1UwOhgOhRMgp8PNBhZ+usH2axqWg54MQaZ+CEdZxPXaeBCRdOQ
FcAvAiReTSS67uSEjuT15/IcgCWXqSnwd8u5NvRIPZKoLbiwuYxU4pTp2vCo
/vQmcLgMmkaCIKmE9WnzWVS66xNQNZrB5NYxFtB0z7Mrj5g3BCHrryfYp9Ym
2Iyr1g/3+cj4axnuG2As6tjjj+0lb8Aj5t6ueYTmFH2aU8kOvI/g9GwUezwV
f6bJv2pSKDAxXEblNL6oKMH7Qz/taMHllidAnPBEXqTUMQdJDRQEERJ0pMem
2674owfO0c2ZpPw7xU9Hptk10pNnF0+rG/Hac3Z6+uYjjLPQcF0LjN0w0oON
dqqYNvLhkdH06VSsRlgFrIu4Gq6dvYJBVK2OqDvX1NriGrPqE5mxcV6R6an5
Ey3+ZrQ7vFNYLc/BUlZhxS+p2HJfnMbmWNjesw6dQJyDMBh6xW8niFGl5nDf
ZtMGVJd4s1l+cx27AGmnA20D/4w09XdCAJzOG0jLBw4psAHmxXblFf3J7QGw
rD6y5gUtcg54m62Px8q+e3T/0vLWR+Icrr0fghnE3Wc/mK5xEKMcrqFT1TwB
BhbyU+vhnFSYrFNQ0Pl7pgilJwBbeSvjAdSEMRmru6QIJuISy18TpVa/kcHO
bsnCH7KFef5exQlhp7WKCvqrtHXqjaXz71BbMF6XonHVpC9hIIrX3fcHoHsm
0PUessbtDt6ako3xuXTwlbofKg9A7movrRhCb/ReUp7U0NtjHSdgCqAB0Lea
PKxEF5J1hUV6IBbqJu/A3op3GZTnoY0Jqay2q9Mp/FhL+BbIipd702lLq0R2
XVo9C3P3T7eBLSmyf87/A+pFWd/5UezHHI6VUgDnQfIDEdj4J96fv2f2Fiqs
rwHsCtvTGVdd9YLPcmvu8s7n0jDUPRjDO3QdzyYRhtfl/8uykdEY2r/vxode
OPcPLAKrDpG7P39HfTSYI8ydLQ6tIdUNhvARHy/ArK0M4D0XSdqe5QjxjZwc
CaLghXIs8bxVSC4HoUxFq8KbnxOCYOIcJR+fYyuDcfcKTSzUGBM1k3026ydY
AFL/PR9kQxpSy8J+i2hgk+0JpeDfto3a34u32/RjDzanITCx++XGI6IKYEdi
UrQ+2dbBN737goSlLev3ejoCse+bRGqU5LU+w+7K7Kl4DEJGlxZTYqyQmXQs
jgDBD0Dju69BUErL7llpObyDtlXkOZHtk5P8Ah8uWy3vGn9p82w/YvFoNdYT
auqH7QDu5inQseogEbZS/ymj0G4wQctKc9uuQmtUeEpJklPNEnIcy17P5BoE
IJOTMeWLRwkJJPGWoe4FnM/FgpJBU+ilx8/EN6tXF5rkXp9kIDZYpFCoeZrz
rOJAMZdnDIKTaWssT+zirBQ43koD9ZubFR79+n6ndi1mPcyK/JxKA6wzkr5C
omaO9xsyLBNzTbhFtZ8ImpRDodtNMnFEVSXt7J/TAHPpfEwGF99MxINjmctf
QPx4RYlcKFjR1rB9/LV6nSdYuIGZURep+Y6vJpPSGY62P9v7+MIm0PhChgk0
45hkt9i1VB9t2TsjPlU3XREiai9g+Nv6vwphpejJCCMzgkUgJbKBoyy1srYG
CK2dDUkgF50blkeAA4qwM2XqXB5q8DhT5weePBdybHPuyT9inAWAiZazE9ks
LNicztOgRrF0UheS0cqMDlHqy4UwCvvqxPtPEpA/29msQO5OAWTyDI9jXRxo
I9cFJmuCLhuKu4zbXf5NCLEYE8NIcYwYYsWPc7RrqRJxxogPmciD7rtoQIZN
flyrF3yG60huAafPwmSTmLyS5rH39sJx325V0CsHgNlH4tjFTQgHp2NLvN+v
ze9maj63QTWgUXopcwtoYmMmEmRbNs6MCVW0ffI6CfZw6Ls+l1LtosBgUIuK
FM28TW80KM+zVFT3bgrCRipAbgESKpSw5iKkFGAgLppgUVfYBEhe0WlMaEhy
ey3MArk4yjlgu15eWIn+nqt5bLaDkMqPbJH10VwLSHqglUI45L+v/bvW4i3Q
yJbUU9lVWGa+AKNXrSbBYJNtnAAECMvJ7ZQmQkg8Q5qwBtnn0IIeQq1creHa
yRGdM7yB5Rd2T89umVhyav0/DJQ+NVyx5YCaEkbxgMplttbQ9ASEHjo2lGJh
9KygwK5DM7zbyiH15v03Pl4fAMJFyW6yIsKf5Hk+/nT9IpPuXg6OAbCc0cZl
aKIGkx2NTJPo1GJbcpzzvn+4gxaQE2X4qgV+alCIO7nL9jKNQHnuPlMbeFke
TAoT5E17+F93N7xPOH/Ym0BoMIQkL0euvnDz+h5YZXrfzY+ivhzKd+/gFsSa
UN7if9N/QJU7MrZk9KHa+psDWQZEtBTcNeh1lKBd7uzJ35vdWfk7hstEZO/8
HLq9Bc60CjBD2mRRSZ9XUbgNkPbOHfi2clVeu+qjZkPyR3qaOQ01ADyckfkh
obxhCU+hOVQTv1yRC7XyInGnkQK60N7mBsAZ7L/x0i0lYLEX1t98R1LgUXJ1
L1DrtYwoBpqvAAkLC2hZxo7xkKdP/yHbxKyVy2TYVhGk7vBSa+F6P0tmH39p
x0oJ+Y+OP4K7nPjMZUt+KwadWU6uqX6i3U4rqlaOafiVBq7gdr8i24KOdaTG
jO6ayPBNUkDLnuQHrzgQ4UeqAW4XxlVs8W5xnWiEYLSic+HTOaKE4b6MrlUT
HLEfhLbxdQTJC0stc1HpG3VzbTBIGoQbf9pXiBYNFIl2ZDQ+E3c7jTVnY+YO
zNyqr5tXMq1/+unrmv3q7Iada5hV0g7L675Anr06gZmwXNcv5zm89bpirf+F
Xz5pLaSEEtdeVWV53DfwUSpQC8mUE+f3o3GGWmejLixvy84dy7iF8squoaL7
vMaXAa1o84XTUr7CTQIcGNedqcVCs6inPVV4kRAypKzZqBagzoHrvgotGES7
Fj5WiHa+cKr9m4x8xqqhSr7+d5qLbY01+6eZyO5EX1H6hT0nSeLc8K/t2FzF
XaJH599Yma9dFeaanRctlZwdhd4ddAmZXHOKwYu2J/eo8veTHHJXF1jV2fc8
gPz688aZ2yMqFHbM/5p+S4FQgJnbRxKnr838sEpsc3ONxmeykUUW36UeuLjZ
257l8OoivPRUtl6WM5/nwfAgUnRfoeFs1M1eylurgtVy0Ek80TEM+M5F51+c
/9CTAJXlswbr5EahdvawHqJL4OhyAC+zSL89C4H/wDUKEV7HJqMQ8AdS6HgZ
0ti7fKpFGapuMuVECxpJtx3wK9cPWlIuAgEdbkmAnzN6X2pkhVTb3juzqZqi
FCRzsiBZzXg1nSkmxGHlwL8KlOvmu+xNVZf00C3gQ5mlHklEf2MGu/Zijipb
pfLCVjnleTlPDurGOzBhWxUglj57M2pG4WCE2zSz7yOpCZo7C5RE2NuSTkvh
sft2NqaucQcvzYqlsNKv/C6xm6opH26Jjoix4+6SrONzM8sEsWYbxPQ3P5Cs
GTPbhG9E88u0/kxiVjrPQryy84hlwq9+NFTv+NlgSh/9HJj1jVazrVeSi5JM
UwpIjl34GI/pCRyJ6S8CByD8mxAibZcLN3zoOKqKXFQoDruUc/E61LEMqy0k
yE+j6DjJmL95AEaLSXjJo3xTtdQk98e6NUYFr3j+EQfLfXH1tGLxAbRwUC39
G4ptIl9GkW3j+ufbZV9iS/AgzWfvWkFkU2Y3BGai10ATr2z3onpR5Bmo0UTf
9bARobV0qCgAH4iz9jmmS9SHyGTZep9PjNXVMafouwzT4XZI0dYSGdHGnQTL
ANmFNF9BFwLVCFEPYlHwZuxWSziJOf9g1sWIbSOVyn2Ivylm1oGgjgCPMhjp
CPUjqKVes/rf4OAU0xlz0fxaCs7CS56e

`pragma protect end_protected
