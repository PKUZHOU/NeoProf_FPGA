// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
24C+aon8ij7noAKK9q2owQkZNtAaS0R8iDLC52ymuf5y+lFK5Ae+Ya+cFBLdCQk9
2FsrrC0W4A7m26h19qjd30CAjYbymv42kZSFXqjsAjNsaHKnsDmYbXljnRSC3Fhv
8wM1mFeLkmJn55pmWUa+qdiLl3No0SnKRtsvtE8mOG4RNZXKO3EdWQ==
//pragma protect end_key_block
//pragma protect digest_block
QArz3L/m+NIdd4ue9lJwfBB4NMU=
//pragma protect end_digest_block
//pragma protect data_block
LMraHZ73hBmhGt/Txmg5ilIBXo1pUyqHmm3W9kv6TfW90PIPH53+koSs/4VDD8ve
dysTiYwPkXAoP9A2SIRxGySTxcvdXWcwPA1G8QKgNg5NOgVv+gfw9pgQosbbA77z
YsHdVq59+PXLbiMBfEtSptoPtb1gla966FNT9C8/0cacRSc8Dn5WwtKP6KtwB19a
/oBqV1MnfbzNjJdapZcpbnxZdkI3Tw8r9xpcgodFiroKY4aa6LxgbNTXUHBJOw+5
+0wIZrR5IIc0IZwLzl812tAqR4b9PyXHFTSnsqHrq39O+PnwcYIA/xutIp1mSEZd
3w/TyYnOGhaPYGwjJVmKtbBiJJHdsgsEggqRvzbKnJ7UIPfT3YxAXULnaeAht9Nf
0yUmIxACbCDAuhPxuqtqVD5Hrodpu9yK3kvIDk0Fd11M6FruVbs4HVX9RGEGCXuP
FrkkPaVg+qtC8PvhF5raVb+X+aae7yaQPH464auqpzHUfvA0yOBDr4Ka3P2if98q
j+XZO4u29tz7yK1ANqDF59PS8GKXezP7Q6SynsoCDM8g0trefGTA5D1BeJ16OW3d
4hc337xwU3/1J7VswjNh59hOb7iT+qS70sePyfpLW9oUkFCAHOEkJFxn3NCovULn
jFuFdLHsnJrXoZBJAYf4rrKOnhJfxq9kOHLxb5t/UZAXvdcTRkeQmG+zLdBOfIVO
PZV4z2hzkOuFU44DspENcbwUaAC2GFvVvHAcvCo7Kdw0Kc2UhD8/JmsBA2xZT1rq
9LKHvicK/NazZbTe8nBRgedYDP9ciugWqQ7NNsODSAbqd3c/hZEl/112Sxpai3Ef
+xMGdSow4jO1ewCc8+sIvxMV3XC4n8KGAEU2XT/bMd+MlepmNzgl4yjavVwxCHK9
Sz1MSdkgQCH/IVVyWXG7ytkzWB9s8S67Q3y1n9fiuU4P5xpc78I2P+KNCl43FO9R
Rm3ak/UsmWyTo6fTYn/C3VL/smtMg40QFI+6CUnAhsZeePSPnOPpQxUi8bL9aJIG
1oDcEe6UttTlioi5gShcKrYz3WmqyLEZtqcx3CTTp76I3gjDw9qhzinipqncnR9j
b1c/4NMxL0AyOu9c4pKRdYPAbRv9SYWaW2Q7b7wuzBF+UhK5f+SnS5kt5/B2uLal
fhRecy4KJAznM96Ed2TAbdmzVACkr2Aq+b+3OFNyglwf6GaDEfQD5Ik4Uz4J3xiC
vTkzH7GnGDGl1WyVf5KlJHtgVumhgyYKxY62yQ0GEBM4jQVnbl15MJA3bsI9/qf/
YMCg/c5JBcSBuBNzo4os7NIyzin0I3WV2KVuhm7SMFj4lSQeXh4//O0KtsN7K1oT
+GpmLjRYpu4dedgGEeP9Ao6wOD4Zddkv65RZWIr1yHsoUl2vDIYZVaQ4Q8/wkp3Y
9P3qg/A/dX+LRV2Sou0mGe4iwPOQi9+HkUxEvpqwd3XC7MG4jTQpx66EpjH41jUH
6KWwbtKlxY51piccb8vrgs80rklie9JGqRBvrB6AjXYqvydKLZbHQJ5kSFYn35/I
g+ueEVKVhgIzFOsghKFlj+9XdlAJWWsSM5dJ+4l7Eq0n5EX9otnEPe5RYLPaNePh
q70zSryuegbyI8Aw+WOOECthjtPICVZxzgQPMuff6fC+fSTzL3zrcfgaUcDQwBIo
4r1gcFPyNxOVPd8kO8j0g6f9oIMM+7BzyjvV4eKrKJVnYQXJXE9zd3o//i1Off9M
LDjZGGRTzW8gmn21AhZDx2rnshfZOx9f8m9zCkVtaEn2PhnFX0g6H2KNTB6wm8QE
dsPG/yM/faUtZO2PACQV2JP6DV2rtjt2Fn7U7ISb1QojUchkA8lWbMTygWNFZSgV
vHIWCg0S/mJkJ7+n4zywR/nuWvzH9FnZmbFapaCyQWRdbvHX/LOv7mgaHrBZnd2s
6roS3dqxBinyWJyY+Q97dIDqm/RgAexrCZJwcub4Uj+HaXr8mOq0GY+PGQTkSCCs
TDxKNNTtkNAZyQxsDteQiNAsHsImhdKYUENFoD6hqBt+KgkwoH8eJ7KZICApTdXn
Js1F7q6EB/2Z5xvQXkufQQslSHSOMOoTsRT1vsu0XbGQMVNmjh+VhhMqFm5oAnoC
MYQwFFvpVzF8hSCo0eWPnrwQRIUmAMmnC3J/YyaS/+k1by/Lw+dfj7cCf7o1lnwC
2zO1ZaeJUuH0ybQAfflRDXCpjq7fyXPhHEqrfW3YVMV3uRlSchqY43E7s+CzgO7+
c7PBJVCBRCJYHqjEg/62JD9Jia0dEo+TKslqacmTYMxlg3ABYog+Eo/XnqeP8vUF
Mbcdff46VylSLF31nS6a2nkhclVQGfTodlm+nO0wZIC0bEpfOCX/DhoG5ZmQ7uR8
sKrg5bW3PfxE4i0QadVPMyZeYIrRV5Nun2JBlC787bDlA/qFnCRTH3ugdyetm1kN
rnyO2zCY++IM0SbgkzZ9/UdkpBllIcKB59HUMPSc2lqoQLWCLgokaB0dgW7r96Ni
OFU2TP7kXPSwTZn0lt24gTQkYaKEJLviSaNzPB8Ifwtrtfvpr4pHieRXAopERpyS
sD7lctzA6K0zxczucDgFJaGTfI3o6ke6zajSBiY9A/KMpGdZT9Ds8nv/3P6azsOo
YWWQTkZlYGXts9/XWVkAbSvbn4AucXFZxIaEaZOmJPdC5w7LGNVuxKU3tJ2Y2cBC
p4YZzCZK6ZFFNNJ6BikRtgM4XdUj+w5yPMAI0rUuw9QBS4sqiIX+lYdJY228jSW9
rbgu++XJDjAZd5S5CWo2mQtNb57hLRh4lTfWPFxaY8mubc5YZLQY9dFSOX4Mnab9
y7V80cPousK9vi8iBRqJuI4dsp0byWSucaVD2SNcUKikvUwvQiHA0FZ1EE42No6w
JXKUdwBtMfC6HCcr3L+JVJ/zjZm6RI86J4KtpIlA+/c4Vc2oWKnAYdL1iQmBW/Z1
n7b0L2924URMpNCxqOsrT2BEtmXOwy75zNp1+dtbRv6R/sNMpBgYjP+OpLOq0wdP
J7oAhqap9F4rq8zvHxIdqKgtdWcmZdCoBzs41GV0nCAMKb6TF7BjUUcng6owFo7P
XJOYTCYldbh7Un3X4ddexCb0EQrv/LrIXot76EHKfBb2GqVswkLkLrV1RYN2JIkF
Am1Te7/phHb3F4lbovn/+vHh0oA4IJjZ5kl+QBZlqEquLo342oInLkxKmvQppsuh
IafTC3oqCIFH7Vx1R0AYO4tZ9/lXWU10gpwiJa/6pHP04MKACjMysOaHi1ci4sWi
HZWQT8R7zifBnNMkC3jXnX86BiZL7rwaeKS7OZER2R6l3ggmOogjfjBUisRvC8cg
GVEyI1qHXVyuvFPc7VjLEnZQTYThXBiCErqI6P6f1LgYBrcBTebUGEFM2Q0rfvpx
vrru9OBt7r6raR67Isgda+S6+6KWSCBOscWYYYhKyKY9y7iy7ejSalybq5INNdod
KLUoNdOiMYhFFRA5J5/FripieoJsE4wEHDSU6RMs/kAghl0Y9ryJ+aFC+DGBx4/E
s/zZ6o0ZqHT3FQhRzKO+uKbjunTLJHwmcG/vL9sH8/6pJWANrko2Bx1DQOZTaxAm
oAiIq3lauPCRhJYyzTg9yHhEz003meYgZ9suTxeUL5kcssriqG78dPnZ/mFpVc77
86hqxRLIc8TX1mLoEpsrM+ycZ7QhXvofMlpEqXdlpotcZJROYrrO6oOcHT44TgMn
rreKuW4seXdICk9eBpKADWT+0j3d/WX0/NAxI+fpeoKOPQXYPL9CTE3mtmr3G1a6
oINoltVQHvi6Csgm0dKRvmUD29AYf4XOZkgCPa1c/P83xbxNRUxV6rHR49s/G2JT
14jnMksmYCVngqaGgvzRdLwobf2w8CZFigog8n6noy7z1kVasGO7aP3TUc+C/Zem
vwytehpOUXXkZOkp59s7lZn9j5rDi/N3V8EV/hVThrL/tLJXn67zJRx1iClXwM0q
lPbbFgzyl1kfWFhZ0JWAOZgRt7/bG2ewY5G9LMfH/ojW9uEUR3U5QMbTbnysthRt
sz6dH66LdtLyTpnKb1t2+UnXbx7XXCMgA6Hm3ugU9PjkqeD5knOJqF4QFhbnAdUg
lnRGRkTs3IRaa84yqlJlaOQMNprRoYR7aNj15kuxENxALxsSqA49dAhXSNr76I7b
j3Vv1yNDMFo7oAFJkYWZ+Dh3pICfgZ8VLoIjCtfa7YNWJPdmUgwI2bzROrJtQj7p
UnDAFIMtiHFWY6z6V1XNSmcS5IdUmfw1Il0IxZ6Gf60B7ezDtbZsMPifcKzeyP80
bmudJAb5xFUyqq0xKQvFf7jaT0BHx7WmOHqHBaZdiOLQHrZulEgOWlAHYQ1qBJA0
YyCxVNg7KdVxp9HmJi9hbDQPZciW50rgw0cLRi2UZ1bRHiVndUNvC70DZsaPzt2t
0Qcr5k3+gwlkTe+sZJAaeTzjqOfh+zbzPpbG9elWa20Suw3kPD6VtaDTP4LGLnJ3
5eRCDG6JhxOq5pfmjDifCv6E+QvpI81sMpjqCzxwBrMsgikEcty8uDAGxJbuaRyn
QnWhEyFCML9J4c8Xc4ka/EAJUIfPEZtrEacJk1muCgUKeGBHKS9G8oUtRDKfn43k
8fKmJuwSSU4v+3PRm5cRZ3jC4BVWV/RVXC/7xy0aWHF6hNUpQC8n8YAbfoujiNDt
dSWXbbcr02F8Gfn2ZwEcJDGI87nvf/49ShyZJRPkxhhmUaDUMbfWI/oc7vLcsR1H
UIZvXauacdbEocTDCqrdDo44+kPfd150YeprIzgFQbxDOPKAzSfCzjDrLMDaU+Gu
7YPMAi8/vk5UI1BI2tTlpTq8izMLteDSgn1OTgO2Za9lHB4MZY7t9imwT0f+5DIO
wLvhlikJ1/z4B/xTzjeVwiL4f3gNO8HIzDalGjO9QfeFzk3aWPrERn+M7FkOaXx3
dI6GLEVKp3HNOCxEirJqXOG/c9EbEifUFT60HQGLsrDQyanX6MF24EGsMs0ojmdF
T4nV2tz8bqhsdxwkK3URFgVDHzBuXzCmRev+dt6UOJGLJOcppldj7AVVAhA4qRy8
P8nv7xEmaZ2vf9qq5XZvez27Of6n7xuJtNsOy0V8CC9gxT55aEGNoD+ONUbfG6w/
ailMXS0BX58o8NAZZubdl3EmGJfHR8Ce4ZaI6foKW03EEa8lqUL6BO6zl9JZf+/t
n3PpCkDvdOmxj6HVH8P9w9pMXURm5iaLu7N9Zv6dF1X0O9oLY4hCUVZjRY/zMubS
A0Ut98F2McBIOuQwSA1QhOqy3VyMFt4au9e1pzAzYyufmTn9CeRD9TbHGOKm4pNt
hZBdQNa2r2r6cuCLg1O9fl1zBnVoPaB7oIdG7zs+PPwLMQHvhRQVMehxr7kxFWIM
0GseyRF1BVhljnFtT7Cu3EJPj+hfx+SGIdm8Mz+xHqDZgI+wJbFpusOGM2RaWMwC
4JWah58n5j+hzNVgmqRYHu8QDYc/LHzbkEp7yYHir0dcMKO7PqVfXyR5ruEk6Cxv
Apy45lH4zK7JSYsVmRjL2rS7kMfz0l5VYntvywa9QSi7XizlGYFWegSn1qVNy6Sq
2ArrMb/Uk6cvO+hWZX3W142XvU8RptEls1IgW+Ehv0ThEVjVfXwLIq4iwjI2zv7c
61TblsyofQg0pbenUD/ewxXQpZns7ZJGdmbbjRrDBMLBKEtFgILcCXXbmfwMVH1p
bmFdvwBh+vGmC27+jXT7pBKzIkqtbpEpX8Yv3Crf3/lyeY4Hd53+FqZLXkZC+lFp
t1AGuN6vnSQN3e5/EjWEXMl+aKePXTTaKgl/Pzlwr64Ts/cT3O6mjZ6oX+K6eUTn
vB06Z6RxoH2mEq5QHvHzT+iha++bFFByRu9V7Prj0yzTfpCnjB6fM2WWv8dnV+Df
xdpGz5EGJZnWAWqqAtdf9e2iWxM9x7MN8KCCGcQhQVqj4bPz4ODhClbo9RFZA3zy
umsubl7qLFOALsCtYO1nfTK34raEZqsO2cl3KCpmRac3aF91aGH+1s3uWV9dTw7x
VH3M+451owuHQX9rkeOXeDzSuaUEepz+CJ+QELwajPgG8sF+b3rQxqp0Ur5ny6Yq
VzchXhuZPbxqzB2Ob1gf0TEL/gUr1HG6lzNlDl1BF1ae43j6LHDh18FGwd2OAyq4
3+tkSis2+aYJ5nEzI4layHKL+Nbt/7fboywP7+Vhu9WqJiAUypBXYRUlfkdXzp06
U6PDFlvm4EWYFyvnz/cr03XwoFL4segUVJy3cYdM/dVN7+qUj96IsJ+Xcl0Instl
c6u4Ji7osYh39+ck55prScDvtQU8a3bnfg9iIg9THieZw/lB2YB1RpuzUVtddpQ5
qwM2IcwYAQavBqzUFKiOcqwcSrHHIxSFmZt/Y/UxMmImyHTERgNxBF17hPqTiSVX
Mu6KG8jYdE5VsDgF7oEZbzWqF3zw7Wsn5XmAKU16/dxjZjmi2IOxGgVkkmx96NFk
Er7wlf48or/snpX9zerECoj29bfqwww6jhdQhY6WhQzvK+nxmhp/gNGsML7gkgcf
XQISYOk9yMp6JFWdu4XBVcTNgod+N53mBgNZ/7uXnfy0F95R09gVmR956HoEoPxY
MwQ5VjtjKADz0s2sO8cuA1eMlCDFUEgaI4KIYgZeg5hw62VMRrgmW0xVLEE0WXN4
ptXAEuR4p4GY8A4jfKRmjSZlXqvWWv0wAS4iDcVMYjTFjWxLE+yq/MIokIIoNWsd
LVCGWqlp3RWd22wHR2CODh/DWAkHz0dpS71Oj8QvEOl1vvsVU2JrAnZBgPdOgOKo
LWTj0JuWjuwkelrEZjmfCuRFSxeMZx/EmEOLRT5QNxqCEp4dHYJ95P+aS6bxC+TS
/+uFG/VN+bN7TMez4GDLuh4jndfRqgWd7re5P1kqTec5KgjNgbgG16S1UjBfXadk
PYt1nSmS9doT2goQKouHSCFTlFpD7k417zEO1u/z4fdZH199ciX0GbhRvSAmx860
D96zjx0fwGGC10t2ggNkPWSjlBp080uK7GxbS455Zt+Mut5b260S2vwiNSbzFKnI
K74GV7DOGPa+mQXyGihe6YNfV2byb3TgBXPV/Gjk9P8B2xs4Wrrb/0wJTMyrNM8l
uhqAgijSMLwbt+Q5ThY9hEZBNBgKIHMh2zYAa6syLXwGPw0R9F1oTS4olyl30DpB
+ucs1LXg7ICCM9Okdjvd50GX6vgU0m/HavWZmm/NBS6miLiirAAtnGu+KRs7v7Q5
TcXeOB9C8myeI9rEuOqRUierajrDC7eX/3UNOcW7jWkyRGefkSH+W9iAwxn70MGa
su0hcTIV2mLOlD3Q22L4EjQmR+0v7/b5RXSKCtnm/hR+lge5ZSAcw+CENfnBfMXc
Rn9DdlwNbWqwEhAW4cuYjBsFAdUBv6xqlhPNLbMLowXSaXboT7NCUEkxVSy6Om+t
eSUi8Foo/rn7f+OHTzJ9hpUnLsSf5U3XyLSIVJUZ0zdyeXh9ym9/QSnhQSyGVQZk
LKSuUdePe/Po005WePJHnfj4bmyf1+MBv5APp5ksFzeWO+WS/ugMGs8bmGppSJLJ
ODPyYaCOvUWElktCeveoR4XlUgiwIFeEz2H2sAhsw9PbLKgh2OzNJPp+azxjsS3P
csQQJTkMGJ34Z6p3aCDVl4fpGu2Y1z4PqcBKQCen2SjKHHX+GPeBg1pJoq8yR8hi
QoQf0y5Ds3tpgOF+0OBiG8NfwPXCPDGqA7y2//Ywp6L6y4qXq6NLZl8Md45tSxgF
xJayaf5HTFaKH6KeX4sSlnswJorVgK1WOI2KRYZo3lvlIySuuLOpp/TteQjxbZEA
vNrBGyZV8QxxVZqQnIETJghJd1gEvMmG0TxQKR2tPpVntNnc7mdCCva0TNPYZybO
z6ldlcG40FL7IxUuEMu1j+dmaHoLTpXty211rOe9HYCmf0CadNxGS7HErLW2fgL1
59r331H76lSRZpDGHePD2fVVWC5w/Zpp3cbkdjG3UQel3oibgHwyD8A7SRl1FdWW
WJ7F1WSONxkRVI5tjrCUn/KXa7dAOaSp94qfdvmDc+xOe0pU7BSWQqInrQgorq//
+pjYPKB30tJuhB2nsRs/S7PRy2ycQ+qRZRg+memR3Upu2zjcsVX/l47G+fbg22fP
4oLMaltpNNa6ouTX//S4rCZnbWI91r9Z+Qk98mBUsutr5P+f3+AB/J9Q50SVT4p5
XAo9sH7pvtNx8Nm4r3WYwSMYt1ZC5btM4SC9qzoJriwcV6WtCUCIKePAx5FybwU3
35wwMkPAIqB0VIuRfREVxC87Nf2244VeOBvtiEMGF0PLEv/D1oms6j7zqVrmJJ3J
fzQ86NeQcaqls4w6N35e/m7XWu0vc3AioI/QOTwlom26VRDpui/zFv6x8DP7/BK1
bAyyd15xruWVd3Tm40wtRbpn3jfYjwv3fhF8BQb4ztRPuMCbvIXdk+QDnkr6mngS
sb2Z2uHlA/u8NlMO75ZDu/exrdhK73C3u0+2P1WrgoOXsxjU5850pJ4lD308FZg5
0cSELs5nrVaQ1Xuovxf2YQwXlbeDIb7uEaeQx4vMFpPBy3/3/4u3cm99d9Y9RNk0
8kwAJP67PPb0VDthrkmhZaCDSPFzp2C4GeZDqxz6aFQBnzCavO/Ff7TtP92jOvwc
W/aTX9fZq2WMSQHJtpQvb/X6qsxH+IH2ChPtSYWexkhAmpABW3FfXdTqgMf3+9qV
GFXnLOg00umxRHQATDGscveTVaniWrtAzabeMroBWlzoexTpisNYVd1M0YxP8/MM
jhZtyzLbkl4uJKrSIdWGimnDaYNQUgIqog3pZXt78QtwmPVsWR7oa7Q6NjTO1yMO
bqUSZXKa8gWdPhGFqA+MkKERaP3TwaZI2kCGcPSu+2fmDMro7Q8bmTNN0yls2hD7
uPMKarsv2g5DNJrpvaWksEJDZm3qtKH+PDibrgbOC4AMZyBgtA98/w35bEPTwXRS
ErYvBrDPeNM4M5hWOtAdCKQhPmr9KRbBdbPuRX+rpYi9/itxdkyRcS88dWY17pA3
TN7+jJ/c+zOnGdQQz+LuRXQQdLqJ4tpQpV/PIV3F3UIj0m8Ji08rg0iR+jyKUJtU
iBSS9RtmafUMNwSdgsyrHd4BqVOPQILcLY7KMlwO4Yr7zv40x1NM8dUesSt4uX7/
fhwrdGil6JjT+szKwsj+zAYaX0YTlLLWuG7AQTqBdE7sQeUe3KntTDmQJO+BSNXS
AZ7gNHFrqcNi6DHgM50Bzudakqg8Y+o9zA8sDF5QLLXnydJG4YJyrizhKTlfMvfw
z+vJNqdUxItpWIdbI6xwQrGbwYoHsUoxOKx2ud9sOHk1rFrgcllg4zOLEglBuU0/
UuYE+NOkbVOj6kBT/PiEFivEk2VdwGkni32J/jrha6GtnlYvowIVTpdjt1/Hz8tg
0MmtjR8JQTAAz8KANKUmPbl95F+YyqtxDGE7OVZadOwD+0Ss8bQ9arHw7fEbdpMz
Ei0X4Fwa5ZBxAmv2CaEcIGxPgPlMMTu/gdI0V+oL/fobR8TPuzO1f/1wngxjNC8V
VN3miNrwO7suMs+NGbwwpiPvoX/e91G7wY7kvKEzTip8rtjSXxNx9XlxmwxX2qee
hgoKP8KVTmqsbzHbgl6s5BXnXq5TrCshPt1Pd0j+34k15vQQq5gp2gvgCeOwUQxV
C0ZFAKvx0y2e/D80z7GeH2uv4axePdN/lY33jgeWdbIc0ToZWIy/71b6QsnSZtnC
26SgzvBcR/OrfWpVnyXarF3s3fIspSrmhL/fbEAy12xTyv2lD6ncPlP+uul/H1j1
qeZK/+nAmkfnRqlzcfy485VVV0Qbyfxfk/p9P+CNLFSwnMXV3fuZ+0mIyGtrYQZx
wZADztmXH5negLSKDSihuRZVW3GaE9ZN/naAOof6P9zKrIYNq7PehlWr88Sef7jN
xYOQBvFB4uaj3Qzefqf2kXdDfC6j0ukSe2M/nxQgyXcPUS8onKfJ/x+ijjf7ic/y
eNMi9DrW/FBoC//Tp+Qfs/GOuV+/hKBDVDfmxYfbpiWrag5D3rOQZUxa8yEewuOu
SYpsQBwznWIX7KN4G2zLYGIpkNVaTYY4NFr/Gh9yAQBHqrMUDIDTjQyiujmsl+i+
GZtnRCVGZNNsNC0z+PNIUYCGdfwDmpXYfep+jLtKM9yGjm52Nvup4DFJZZzf5QIb
TmqpegXoohx1buu/Kmw7soeP+sJQrb27PI7Z6xuwnkFnJqqT+EDyX3uCucaV4fO5
scZ6c5C1jjqI9RJgc8YFoseGP3fcbZITl2axqr8Ixxfi63jNwUMWpEQg8wOfcFyD
cl4h6AbVN1O30qb0fsKfCyUz7+xHzqTzmhij0gW5cIaR1Uw/vjxwT1FNk55W0WV0
kSREJPZDp5uc5C9C2EeDpy2nGtFtNGE7iUatnqZ/SpTNGFBpQaWYJwq1p2TeglF8
IekKQ34Vj1ejq/D3DIZh4MDDF/9jjv57syWLB61Tj+PKQTHsfh9sOHUF45O54U1q
lqM0rdyc0ogMjbKwgtRZr9G3yjb2IXa4XAcc8ZAzwtf2us56ISd0P51VFmYU2ql5
R8Tq/JqmSs1PJPuTU+Zc+CxbXDKDs0OWHJMNC93hXd8PsEXYApj72/1xL0dB61N9
aLKsAvamr2i433mFi+QrYFq8PX1zYRrv+8h2KZwUrXBMjWSPLLC6II0aDrC9ODRa
YojeJJVOlaqVr5W2yMS4xi+z0AqfxuaHGNute/9xV7JjQa2DQ75OisLqaMta62FM
jsGtNiUuV6vuedh66VMD2KPlcC8ntB1COFpw50WLRJlOHqTCbgxqL77Ps+SXMleV
0u2ER4L3JPW0lRNLCDm+pedGN8tME3PFBbRwG0uFG1ke1BM5Q0ylp6TRxqgT0Mj+
LZuTQn2waEXJUA2UPZoHRLluSO+Ut8Re/SanXXj5bBETHgxOO1JM3NOrTwzGbGqr
qUdoG4E0taGLhSmiC0UeC6SiP+1AXLpf6fMBVoNFCNHLmRXyAzj5zirJNogRf/wj
WPgKTq+Tw4YXu8UyhigRyTZUTyLVSot9I4kjbjKbHQrqv9pvcySsLPnmu8Fs+udU
+RzAjVknW6ivto6agxGeWuMllGaSCpKUxrReMMOqwzDLH2kaLIdLE2E5oPo10pZ5
oVW6jO93Q94xEIYzpTt/PVi13YXiuwv9hCZw1Fy6kN2I6n6aOqr9GokPFs3QeJ8p
PFJ+jGfGF5/AYwZXpu3zkwV2w1JLhOZSTKT1gqVJi6esOmVGNWo7c8fcFgzyJ2sM
HnTTNQwntHRGthGZSqB6P0wyNM21QE80/j6H1RD/TKF2tmEzO5Skc5GsQaqm0skG
uNE0n0hP7jDUeo3+IIXfZZhEhqqkTEV0dAQnaLwCLe1qfTuT3D0j9uwdptIovbGF
fUX2D4oglm5fZbxPMG57CAgnq5KCMeUEKpL5G8OuNFdn1fL5R2LT1tNloPXahWPl
oqTsj9LDUNJHNho2DUNvFsNnMKgiQzig8SWY+XAPelpxEcd/9wJLlVpdUVNeJsHA
ARH8tdAeXf0m8pBD2nknOIETxtJo1dlnhr4thNXSiBx/9YTu31Hkv0SWFEo2rroL
l4Nvxf9pC5YPPPA4y7FpNnQErQ1YM1IGfHZIViTStYPfG0axkXyGmAzzIrqfQh0F
zyom26QKYrn1/0rA1RTTc1jkzb4tV91Kje4yrAOuG1b4qmKhwaIWpsz7IeeYGRXr
VE+EcY36HB2AlVyZTVxh0uNAgoxByeAJp0tXK/a+j9WYyxLrFE6L+UrfCeVDIlV3
jzjea/qzLkHeOsyrMT4aaqjhdUiUjKppWj1i5jK+yHp4J+9ly6r4bn369vegg7yQ
cgl6KoC4gUCdmSzpEt48an+1nUNlG4H6NQnw0TLMz0IEyyorAw6x6db7HM+yGddi
POw1vyref/Gi+J4KhFALLhIRqdTBipC9hPV1D4Vx/3DdYHWrzALL0sH7OOorQ4zl
WsCaoEpDL7t/n08bUM8t5tK5HLAZ/54GVZxC70kmxIKEAwX88UTwxxekVoQNe4Xz
M7+r8xrYp3uYmdOy8gQT3XX4rmVIuHix5SybOZiueturiqB1mPi74lt05sEGkD0P
x6z9YBo2iUszin2SRW3BFaFrRlJKhWREyR0+vluTQ0Bhlh2DqsufqEK2lmgUSFmj
y62SrHxaMOA7bdGUNGIu1CK74SZyhfckhrF4K0olnjjutBS9KfKzqssnc1YUfZLA
eSspNPjhAQgsiMarWTAanp1S+NC9wIRDAaiwodrLDv/VCP/U+jQXmUwX2ooGpjpd
wLK8BEtLLXHAUhQ5em0/KApYdvF8wdp7ToIeXp/1BbQdwlznJWLjIkdE+THWysYP
T72S7HwoDtczmGUr1XSxZoLrUHNFkzRX/6FfrQq0WH0tn4/Bsq6yI8iYW66yqxJU
euj69iRA33oBiC6rHgobLCs/S2V6kO7B4RGK7QvdDbxUyxojD/QJ2rmQlFcsqqVR
T8vX2nEYxdpc4rFcGbD6e4q5AOgENn1PE6Y18iKOORNU1MipY9l6dv6fyVWEs02t
7G3PnV0W4o2VNdilXHXac6Cdz/Grdr735uH8YdxMndsG/W8DjngQTrdVJrMbt9qA
b5PLO0npb9JTQQEesaIwDKL9nQQE0YNzAcpIvG8JZbwMYdBU/rjlU3n2N3g+4rgY
4hYgTSO7Oxjfn+DKll9O2VgQ+EgCK0zYRVlLqphPdQpJ0yu2e3MsHhnCErZNPYD9
5Gn7SQKI064ikhEPVlHF87WKwLwTOfxH0427HmNTMLqn0D26NEFam/ZO+jDN6EM+
CvRDqWojhMfwLBAv5Lb1j7t4R7hhV+oTr9zmEt6aLtT70Qr3RpPOeo+Hp9yy5bY6
+mVAF3sw7zNO775RxrM1Y65Jt/K9wuLFGzNYnnPC7xdOD9uZiiqXVT5GsZBMJoVs
oYx0qB4PB7q0JTBxLyqjHowWhSjTmk4FA+2lehSBhgtewSdaweCyd6XsRd0s1uPS
LHZnSOaLvDh/MME9mqStSDa2rPfJHe9sOSe5ZB2IMLRAM1DnGkvQOew6aRpidz+c
pbCWyUQqJMjWJNK1DozXFk1KRcOeL939CZqDx1zs9Q6uplpRq86jmSMtfzmSqnXb
StHfuzdEyIccHKeMwZHBv+6pVoVXXhT7cAxTbgJi4KHn7zqrHVVITHfZGBn8i76q
spmMj5es92Py83bcSLj7gyuKcPKIfy06kcWfPA+cmWSwu9ALb1s3PAEE+iWDLUU8
plCwW8TwfHsXoo+kJRs7usXN5EMh8R881jPKNml2BJ2epWY3Q5FKYGrcYQBVfhk1
2o5Ce3NHvQMGeUYrppc63LMstBHhyrnpoukuwqi9EUWlqBwjswzgccq9KBKualpB
2VPOyzQdlmBjYqxjMgOKJaS8olDnRoK/QddCUZm3Es0BwxA42M6NMP4KVUkQOLOa
FTGYYPliHYyPUfBYeGgw4/Rimk1Ei838OSKM2Kprc6umZy2Lvk6mpFu9Oa8AH+7I
AC2iMLoLSYoc4VCeykuriPH3GxTN1jOqUZKchWLya/KO1I+CEyq0fLIE81N1bZr8
k2QxgpUkHCqpXuBy5Ne9c55Sgc/5p/4+Ye1XxF0oGqyggFboI4joH3pEjYa8UAxv
B6vqfACdyIgsdglQMt1oPAx5eGXSOLg777k+/oZEYW3mlcA6M1uDApCz33R3KRwr
a3+42frlYpwcEARp0SYKj45++EQUYAdz/curdvdOqRis1q3Dfr2WL96WMaVZKJWj
u/YplkHZA249UtbE6CX5pYT/AiEf5qubl2o1IFHpuFTy0/MJT2SLH4valIk8eIZa
4GFNFrhNreLV7c0N3+3vdpn96L7KPQpCMzQon+lQ/wsZiJar2KoCvVEERqgyAXUt
yB9PxB4GrOTqTOVs1FqNaRkcMO/SNjlLc9uBuWbDM8IsUR8e9qX+Hf38TttjqP9t
PtATTOK0K0oIP7DebLvcaPPtR2nSDsMZhFLG95/nVYcc82/9zaYhR44BXUZYIisa
VWduFExhXIH6un57dx8dAdRRkMBHEOgPDrt0g8EHmaa9b1DHqP0o+EjIFUG46lZ/
x3BhAgiWlFXsDxuSVV6UwOlRyE9nRja0BuXQz2DNzGC0UakChPfIIYyTZpT0hre+
VQ1dhSPE3khus0bnuM/cKFrb9Jpe1DHAx9tkf6Gbhz6AnDlJdBuM3mC6qzNUmvcQ
1saJh5UV9ffCtnFrVegr1COEqFbT1KhgEskwAmlshYgV91LLz1JnsluG7I2r0EzH
9umZ7VzP1nU/MQR8zIK7e30KevziR4GRT8AiVGeE5dzTbrW3jJYv2m8EC3Gv0sW4
jrR8uSjQI/1T93hudPQdkeSQU8zzBqMa9Zvw4Gls8/Ii5JCCXgZCjeHpLhAQ4vaI
hdK0UaI6zNXdoTQjQ7QoP+TeyLRhC26lRtCzcR8s1oPB4VOMKx+vxnnwd3f6kS9q
MdFJj6LVNOhi7CMv/h8DyRzLr4KEbVIOd1qB9MeK6b5FjYfDNNLbwD/S7wX7dNzg
jdT5wsfx/xcp4qrzZnxQzRlpfbZL7Cfg8k7+PbwdVjgYlzEn8bqbAAysHNm62NWN
K4s/jNkcNc9xab4N0RftEgoVngbdVPBP3pHkSOhI5jz660UzdSd+UZXu2sypsvu8
29VRdvob9NHvhaDDIt3wyp5sEb15UtxArvpfRxABAjohcP3JGSo+uo2xXrEROffl
ZaxLkzMxiHJ5fWi2qxmOXg9sVzsTyZ6jhDbnaNkaLVVUQ2Dyn67rIAy2betUaIL1
lD5wz4JdjJb67PSX+N7Ci8gZ3E+Wfm79t+4Nq5aaGSsZ0zFrh3iGVkZ3GAFBUauz
kTSn1qmBL9y0AKFtPM4fK4LmB0NFtx2g5ckpMMyNN4LHeCOKF7TXk1OjJ47gLIlV
/GLzAjWPRF1NYYwMn1mS9SPYnNBPThgbgNLRIfZ7dNl7e8HXx0ZDRFwzquqp/ZrX
PS4BTEconjVfaKjhes80UeFVU/9bxSkRHZSTyC/v1l2F3ftiT7BXM6SpuMmb1cOz
f/gzqZbX5JP3C0HOaHWMXmxzk+ZFuyJgdA1Y6InxnTpq3wR4vuKzfLu4s4bf3LHX
oyRsQXdLo9F8DkYqVUAUiR1CgxZ7ZOKLCkDgHPidOECgFPAsK7lhbgjolNIASJiy
d8QrKvYe4mjxYcNX92rdxrW7wJLYincY6AUEZLOQr2/mhsuNLazIWpCL04X5pivR
iyfMEQcaMdDsdJsjOlfnBIR0nJ3QwwPjA8RK4ngez4VLVw2DtetI83kYllfJA8rW
jUMxXegcr2ZdgHtoacTYQh9Hzt6pF8XRHwRO6ib9APHsorzdrZj+sgF9M0npVwWR
D5vy8mUUgDEUJE3XZ287TqIiqV6tMl3zP17YiKfJrX+UHBg+e1wOq5igEEfhXGjC
tvQRaA4Qewepo6fUn/rInWYEQnSBfmtbcgtUXfGnsmrQcYR4jd9HxhoSY7UqVXZJ
9Zo+nU6n/5CVZKOKpuRzejrYUMCY3wVFaGhuiP1BixhbJYIqWRufGgCIUONeOgE9
NH/OiWKFXuClHEFvsKZsKjnGKngLI9Q7603xspy4/vyX21Q9UO9NdToeW6fi+1po
RXKJ2ikFyHMIJa1Db4fYZdY0MU4Pe9JhLtkH+8w780bC0giuw+TLpTXAcT4W7c3+
e7o3GEwp35duwElpn6FzJ5kGMn4JNglr7g94BjvHzX3FWz+TN+2GtysE3h/wN6cl
Fcxw5JCLV4VofKwe4wJG+AnwCJYE7DhVJXXvsVbod3ONyXCqQfebpFXXtAjfYEV4
SEbqeP/b8uhBArJk78QoJ0o99RCVoBpoReX9I0OMKyhhCM0jmR62ynP2Jq3Pul+T
1WF8quB42wuMM4Yx/rSRYOUke4F2NOuR+HAxxJlXN2UL2njha3JKDkQJa0VLaWqP
FuoF3Jc03FqaHH4NJ9DshUrmsPAJK+ois74TahJNVEqE18g3Op1r8WxtpHXO81fW
Q4EFntp20rjMMgrO884wu1KacNQ1AzjwYE8WRz4T5aV6I7z5Wn9zt+YzS2WeNQMa
tmBesz6wsNg0LljxOq++oJvqeXCKywmhrECbpituKEvbD0vM8YjsduEu+eicma3P
/tUjHWuWg37kDO/cSLQJ1s2yhdTOtWTm9UvR9HMoRoP6XKIrsRcPDXdiV+0sbylj
etsYcSVLuloB30wAV4kJQTu96b0aNpG6qthYlyg1fEXyucQKHyBrvka5oQDhEBnt
9prCjKvDsdjSPEDkKmshaSj9UNfXLNeVw8GQTPl6QdnxDU0s19POCS/aoT9X4T0Q
E36qcX8uIpNXR64HUDTXEI6brV2zrYEyEctBapI2lxZry+R5AgUrPFFTTv17XLD2
WjVsPoC9UWzaaG5qqBfTSuuVR5RKbudASrl46EOegPntSLydOfQnr6T60pGrj/l8
6fDfZvjV+bLrIG9wJfjKeQjryb23CDhybQGs3BE1BqUqpHHfSN2oYeR4b2C3BUy3
iE8PYWmY27RZ1wz/0zcmi/Jv9nA7mB4NvcjdpW5xGS/J2frfF5hua2VV3VByORh/
xCHorka3UAWciXF0CUr2GyXSon3clenZUairkfg8xF75VkDTVLmqUNAvKxkWQJ5K
HpxUqJxIOtEW7ytpHJCNftt8r5j10326dt/rb4h+SlT04wK9EE3y2j1lgtVRsVfr
uUIlugGgjQm/Kqd4A77nmnDrPB5/qqdUVhWM7rCFNLGUW9qHRqYjvz1ZrljVS9vw
r4QfXw5WUdctQMM1//1O/pZmlv217zDpmGwusOE41bwIFLhNSr1MTd4rNoVSm7Ns
fQXSwo9cXaF68bk0xDqy6YjTTIxZumW0T4zWfQrIoAoSJJ0bej2Rha95z4jqtohW
qKrdbYlUERSkGE9cmEi/DXMK3t21Vk6WlKEc6vQqUt/FcTh7VVLb9E96rWgnMnP0
uM1du1KiSxy8vQ44TpHkJlPFvYEoQkzI6rmRKMxPS8v5Wv3vvnVrYng4jAGUL631
WQN21Ecoh82IkeeiYvR14pa1Tn2m7zMXB/ANzOxXpZypl+RuOEtLM6X5t4bDoec1
vGe7ZccJ7cyc0pkrJVBMIJ7dv2cFQ/2g67ntdnqxPkxqabbeuIhZlPio4qDotRdu
bdpaLYr8oF3qd9WGsdYehCOhkUaHTNmKcNm3/EuSLdt4gE547Vnp63Q4+rIlVoCl
YLlSxojQ6ZX/RcfiAlW4GrHza30cMoqq03NRiCxU5EGFXtwEDxIDaMPVq9szW7XP
+tD1NhDI3qNo2qce4XJMUw+hpjc21sZhjxNYHX4jERRVYFdEOnSbt37Cf92nknsU
9dVTgrBIWFr66zvShv/sqsdEu5o8yimZAkJzlTZgoGK5Y4qCektxCeY8yAyvZKAh
5PC2sBLPuKbUURh9YR3G+f+G/MrKdEQ7zR81J7UWmBLunhXYzyruaEw5fjaQsLxY
n/VUObTCGn9aKaYeDy8eD5fEnrITjBTsE7nn2MzDXFs9yB1xQbNT0TeK7+zEdp1G
OfDU5WKqSqMd89Siw+vLMaI8Kpp6oO7ndvR6RhKSC0XcAmi697OqswzbrYMFxhOa
KI4R+b6W3BJgcjbs6jKthjLgPGod9jEmDCmsaz7oM/A=
//pragma protect end_data_block
//pragma protect digest_block
3GW8LZv2nhLWWayzNvs69ydjrBQ=
//pragma protect end_digest_block
//pragma protect end_protected
