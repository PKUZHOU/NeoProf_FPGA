// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
anos6BiWJcfw+3p/O8DLAZm/SO+UFZEzi4Y+JBrbCjges+Zpz5xUqfh5y7QBvStE9buUFTGJZsOR
f3Rbtna5pKJkr8fR0TuC/AFp9q7a0/1FZc+EWuo3uu9lfHQ2D62TrYz9Hg7HS6X+TCfoSZ7t/cCj
hxOz0YthJP4lMPNGFVSNaDvQzNkmO+YN3yUr5RHSL7Ujfev+BcgyB8h8f8rkHSyxqhF/v5Nrr5nX
Dn71vCmuoT66IneemG0KZlMxsmC3DMFyFoU6q+ZrtP8+HFHiwpgGbOiU8EPLX2QmJ2ufBHDYoIzD
PCll7IBPBf2QSVUk8/XtWVXYqEGWlB6JyGSlWg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14832)
7n1nOXRfMD2rY9+8X/UhuGCTaFxfGvQ7toPdgTsyUrcj+aNN6fWHRVvYNJEz9ZyCNFl4iH466rxS
E4+gCpPCetFyz7bInjAVzQxfU4THMAfUCOIJ6HxMkp3MyEfmbaNT3p8zuCMwd7ADUCAAMgIL9Fmy
k+KDurQCXmtCC9N+CFzNnLlP9movQzVsW4oDI9xE8uyt0862IVZAq5CS1ilZjSNQ7o3gfD1baTkA
NzP8JwSL7Q3YWuUV4bHMrgA5ajNbQvfj5HescMT+ugZdprmCYv83gWoCOG0OVDIwZQGT0WNC6nEm
PniHScCK6ymJmgqR3J4lQhnO03/LC8pdEIKLF1ZrZ/NzB65hCBABr1gOz4zy5FCid21avuSQje3x
nDE/khweyYeeQhjL0JD87lk4e1WyHgzDtwfMO768ioI/TtYFRd89z/9dv+oxMX0Ph55JOBGyHFS7
oQLsxMrhodeJZ0Sng5m0rFea3ycdC4o2rSGzfPO56RauNceoDn45GhcFxJYEShgI/1J1yDjMw/Lp
K+0lDtlqfuPKVWCyC3kMxl7y6iWN71YrlqMSxCfTOMpxuN0YrmAYcZo4t2bk/z7NKVJp6ZWe7UKr
YmMDxQHL4OojupgEESjqhlzTDLIjcHNYwMhdid/W/KF96SHCdP8G6LRDnluAzJnqBOhUVf2agfbQ
GCEfuOwZA8zjECNwCPU8Otbhswa6s6rwUfv1COBWmLC3u8c/xnKbCmYyANykgVvPo4bGlqvs+ELo
K7qq/S5fLu8Fj8BME9AMZGD5WV/048M7aimFMykFmmJVbqIC8JnM6Tprqm6/5L0QpU2NnEhkb/Tl
0Y1d1FTb8WklSUZCJK8gfFVUaM6oB2+6vunVoA7jQ8nhAhGG82xy+Xuwo9VwddOvkTYQY13RSwb7
SudENcb5CiHPZcw6Xj7U+7f3LkJdTAs5DuY9RkNggfVFx10DMdVfBY/gkv71Sxn93tu08vuYYdfS
Ci4J9p0SVK9CoiVB+KEMvf79GqOv7zsKyYQyKxvikuo9N6AlUAJl3ryg3OwLCM4OnFebcWHduNsv
tHgC0Yxj8yDtdGeCjGTq/J+Iu2WF9a6QPR+Gy/6c2hteIG7QDLiRlMPfAYLvgGNTuu4aGdccVRFJ
800TlfCATni7OLGzGhvqUN/pK3XTb+GJzhiSMFAjjxvseRj24NoKgolDPd0XcAEzQPLDMdtiHHSl
EIoaILBLCdCe6foKvs0s+60PFKdMZkKlA49TgzFrHs+QrN/8qysrWQSvG+9HZx1vb9iwpQlnc0vs
gB4y0inQ9J4sqYD/Z4d+C45+A3DnwHjni5t91q6Hrg2Loj7Oud9cF9nPhjvEo29i07458s46etE5
FMELuCucfMcCQvyqEHbe4giV9UlPHiYgFlsia5v9p3u4uK0f5JcuG1Jl+rSiIF+quMab7UTu2JWk
ju5UU13a92e5te8iHy6a0xENVqIugNVzPVtY6euwC/vaJXB4u1tMiSfYwVlc2uLUOepk9gcAFrtY
2ZLT9iQZZrpzt9AMesCNyn3a37Q48eWEd7mnlZKVmVILGp/R6jnT80rMZ5XG1BxT6d1A1eJRcQFQ
0lJQ+cIePJUUL291zfthYAB/7djZpNaH/xNXmOM1ik6SuuRn6aT/WPurUagYY8SjikV63pbeM4Pt
nFF17kkX0GuYPG3GQtwjoipGyaSzvi7uifYdog3GVfDaJ+EAbT4ci+BZYyCjdu4V7l9yfKBQahPn
9pOEhv0Z1wp87hJmjBevGM+cz9QbBCivdNTNFmWD1x3pEN/vPtY84kX7L8YIiSVKn/nXDUwCF2q2
9vZvzwEmiOkW7BA3gXllPXl6KPhk7/PXAtN1081CtrxEXCd/MisewKfWlcTxpMBPhC4c1ZuWKiLn
wrzMzuiJpDO6uMzC4dsBMavcbUkCYFxyRebZqnPgkXGuYb7657wYDRDeIukrG1dLiM2Q89UrjG6M
VIlWUU4O2QVKbABfpF0Q9u7AIF/Ka3jdN/NfKBbSSGpFC0WTVbKyq9kA3XhtrefkN0oTFdhBilew
tP5T+lgv723A+OZMTybdWB9IWVRdhWIjPDjXJvzhDXO1rcjPWL/GNj1rp79tAG9XA2s11g5gjt7u
Ty7DdHiFwegYpIhq67KZcclg+yRgUy+OiO4ubE2yD8CMpH3Nsq0pKScF0oyTzL+ksxf7BLoe2dTs
KbeRD8dP1Lo/NobsEccEquV5YStevh6Tij7eX6sRV6Tno2gEb3B1ljq7zN4Kn8XyBCTNAZvbFQHf
eLVJVGVXULW+QBLh3PWrokb/f3YcwEc0f+jheZI/31HOKuFQ0vQkfMn+EfPfn/+bQHpcZ29YdBLV
HUWopw9kP35k3sEGR5t/PvYs+xRyAFUWOQl4V8PIDV4OOZcMiHCTJQeNw4Id/4H5ffA+fdiev6/d
ok7/uckd9dNNQ/JMDSv9e4POChmMViaQMCkAxB9/TOE2sC1koA3hISEBfaudwOH4rx2nrZj9AwGk
DyUQq0xG3pXnk9EBHu8N6XSdDLnDEfY1sJU+aiy1QceH40dEEYpGza8oonozSOTBQaWXMeGqSpV6
cao7Rlzpmo4SQ0vfHtKwtkhM2cEa6BcgLJejFxb/lcN5i7Zsf3sUS+bwwj7XYv6VuG8I2TxhyExy
7YReUy4mPLEho1b7/rSOOmU17vvUHaQiKtaFiPZZvFsVTOe2KZz3wf/sI+RtvZ7jYgFPrcP3YZBd
i4P0O3de8ephk1AqqR9oMZBhPjFTpXN+EasPMUwW5ZpR6eVFicsb/GmeVuAUzCTTDpWV7NpmIQfm
q2QVLkUp0TOa6NWPdmHn5QWOdEqvk5qqSDK2DqSdm+tjpnhNTfpd0lc7Ye/t1jB9Ll1dIpY3OMei
wJqUH9SHQumTY8rY6XuoAFtawdIx4XHMf2zJzvPhriHgDHfC9UH2ZVngMApfFdR43WsBkgjsPkq4
6bNxRcS2ldmHEqf+fmiI351vsEkV2JWaKdntyN/uoDjDu5X4iMfSOWKrumU9SECjIu9Q+baYixDb
T3qXb65m3/2hLPqIuJhHsBk40MhquEAwGXQfQuxN8mD/PounGjsqgV6M1iOkdnV2KPFTLOyXOKHb
zsaQBFL68I1vDFwC72Ma9YYHzDw1zSmno3vpWT/RVA1AfT5CDsM2oAP2MlzLkFtPbFecMIlkSXd4
C2KNFTKaF3u+FuUz/Jt0Qrf2/OoSJ0pwgZdwByrKmer7Sl5xCZvv6dhyrNOrE7UwvlrVw7H4W0Jk
uAlcH8i3gAx/bQrRy1FDaVv9V9kqYuL/jcYKQEoY9IvoLOUSYrBnWN25jXhV4EnbTZwncdy5jjHC
z0LByTxsbAITbZprKLA+qkVdCm4pcOHlB0k2volWDg0Mqa/9W3eZahyF3OSI1kdCaD4ayVzoXb73
Z44IF5N2Bwk7XDmjK+lafRbTwgwFIgNBBV4dyQ3bVjpBoHcZv/A5B+FEpzuT+RyDqRxMBeWFM9Pb
kmP/gZQZUBcO2cJwe9RHs/E15alGGEYG6nNVbsRyoh+N1IoMbCRGKR4MXEYtisBAdtp9rasJcJLm
Kzma8VY+M7tW9ZaYIb8GZMh/vcMZOzckHz76+rpHJKZL7zJED0BkiSqAOve8koz6VGxDbuZ0lM6N
IpM5h0iYdpX0Q5utRBx5TxHWRyJy5VjZZ9Ack1jTZNq22S1k+MPyqLsUXDk2ZPYJ+Hrb/e99Vbxk
4zyoP6IXovYrwDPkhbAOc5cY7TmMwImuZ7co/RAOnJAHjNdNEsM+gaZpUH+Bm89wYbnZD6G0ZPhU
pXzbjAy9vQsWYmMX4vwr7htka9DmF/JDTB79iQQdBg1xI1Zy+gLnLoC918TvQR9h9izwyF4vkvm2
E26iCWR9qyVtMeZrA+JPvPit4QeyCVHODiK4aEfLrAWyZ8P8ViNN6+N2/DNIMj//eR+VmbTYF3jE
tq3UjuSeSb7eFssCDoQ2v0z8B2HrdBiCp4YF5TgqQBPofXHdrvsAWBlxSXyVgXTEX3Yrgah7oxi0
BxE/EhQCMZlojfNJXSxGbL8EjVC+wp6BVUww85m+16ddaTDaX3VIC71WBgKjfx5uUuFnOX0xNtzA
paVC3QzaHuNGU1DL5H4cMfoc5LruAFQYFoI1bje/ZMNgoQIS/NA55FqeWqa7+b7567A8uAGOatj8
gy9TrjGmj2K7MJ/0YqYBeuZHOyWqh4togMtaZe1l6OdqAbioguS2JJ0k8QO96a06GaH26Q6vcW/J
0quiJslWPHh4DRJrx0gjCYw8WLatga9PGe7k7kN02zFxY67Xv8JzBUyqRf0gU8bbqs2anUcTv9oK
lc3UFE7i8vVyUhNGvHervbGWlsPOYhjOUVHq7gd0Qjkz6ozoMpbzVuobmMhLzrRjf4H8AMZ9rwsQ
3/j2cyKoJqB/G+tMKEaR9ylXXR3vG4EcSuyGCljp7/EAYI+Uf2HXeAbLxCJZl+7nm3gwjtA+m9Z3
U2eYkncwWLEwRIdHBTMvrS1wOuXDaezPIjdORHAHeBkv+2eWrj+Xvvps/SDd18f6lZItz/YY2Ri6
Lc0LzDVZtOMp2vfqIG6EZjuMnGW+o7RInN+nN47rQXZ/RtsXASCBZfAjlWRW5sNahWpk+OKymBA3
Fs1HvkdoIPzSFlpp/K7XvSy9UJ5xfh/tU64J36YJL4XcVYxN0t/o5UxlZ4udnq97mUHDckGC33Sd
TIY5Y+XHseLHlotP9YuQOsbHOEBph2XQsShQTBvd6/KiGsFsexKt1IcbHiWzpxk05VETGD2Mo30w
CswwOMTEdhHl/yRfJoPC0oJS+NmDl9rmBUJjIUnaKiN6NMl9Xn8vDHCnCbWiDPh0bM3yYk3mhBmF
/WZTcihDMFjZ8UTK+m5wSkq3iPG3xCqd/qZJxjQ7zADa57abRIIA+gNTtlXBR+YUirlnpyDu5yPA
MZVeoN0bF4wwJZE6/iBSvSGqWQi4H6TmnFxgTJcSeo2IgBC0wPUqiSYYbGMviNVMiCsIHe5LdivX
AhlJ1JuUN18mPcUiWpqIaPkgzLDWTBcbyxn2lbA+byGZaH58TVfAtXP5mfWIQwfr0ceajQyUTOS9
JRb0KUkrEKJqcXjts+oKPmDGF/5jTlhnd/1lczL2pZcIs0Gb4A5adRAgKfz5nIKuvNSo1Ivr8t9N
eGL/t1fU8OcxtcS10P1qJS/xv0quZe+YdimookdhT2GF0EiGgqQSHJz/qKvnfunzfWBIeD6y5n7j
RyNrqOqbBXoTlSzdXQarMVUSbiJbzL4wBcb3pp3kDm23cr0CdSrKW8EgNwdMe3oisEIWQGyT1YAp
/4MVYawxEOApeEmZEOJYO4y3I3tX6DfKLMFROk29BqbNHBczxLreDe5XmgTGDeiddicyOTBWdWeg
B9RwVA4wNLjeaK/7xYXCLqe2vux6LpDFt44OBHiDiIc72qxtD9EpUAsfwbq+kKz/ZKb4YOtXEPHA
hmFwgvbY5hE87GlZjuzDLXSp5Swi0xARQPmX/l1DVPlQ996zcg6FqRwfKjEc0rxxZSKWS/HIy6Ss
oz6bj4p6KpMYoQG5yHqQ4vfiRdBWLI8tokPpTUplBubfonN3k+r4D209cjfk42PxGFrtZ6VM22/8
oxNDgeeO0axZ2EuNNJ5X4BS6UQ0odVLNS7s/vEJNH6FrexoJtEdGsFyWnwlPzkPQYSZigsA2uABm
fLSm1nV4TQ2c6VVWC1+nV0Ly1XQNyuyHCd0BR8Zr5mry2kQv5KzODZ6LwFF8JOdMtU08T32HG/ID
ZyAPzv+CQ+smM5Znofuu5GAF+bYznZpem7Ni+jS/kne/ZWh1S3p2dNL1EM1ZS3T3JVKuYyimPyZ2
5n/fB64VQ+wFP+6hyLmC1hYq8vp757KCgQ5ICbVqYf7sAte/EWJuYhpxvvG/zeoZjp/A9MHJeLIv
jPujQx4/movM6e0nBXq7CKV3grr2CWisHAxjAtCLhGclUKPSFfgSq7I8UoBNpO043HS69aCuUOWO
/9kfZfyCm28e3CccHjuzdBxgbP6b++Ln6BheyiO7oITWHNJbWg27xwtf5yTR5TduYb7RPGSg1q7d
sbUuN+sHStrwLpuvNkqWll9pfF4Qrcv3AxQ8dXTHAoUrIuzUZNeGgzhR5Ko5EbZaFqM05mbLO5Z/
njx7pnWPWmyXb7DNQFcFaWGtLlue+Ak765kxVC7DxhAbwmLFQAyS31EPR2pOq1YrILsuQF2WylpR
OhbwfqmL04yTvn5Dnwtj1ZhuI/GY6XNkqzxWIZtNDskSibX+fYYDSrQUf8Qn2olu6d5z+NNV3qxE
4wvniifOt0MIMbvIqRVbBLDYTntT6UP69zo0eZ067RYgO/hNli4EkAn9zxDwK8I8UC7MmdKzI4LO
K71p56XsJz4LnNMBvE3J/wds10DWKP5ER1j7M9E8L0aoIzp7XY8Ee34Ow++IJxBAegGLvu3BrNeZ
yutqzQ2lwF3eMxK8YFppM+r+58/ohcVJCw6ve8VG4DhWnsYdOwmXLGvxo+Nle+r2Q0ISRNieKn5o
H0dqNw6oVm2tY2fJvwX1LxI7hzmMqnHD1OhYl7LEaTgXCp98F7wiJnjYWu2ASIn5As6Q4LPiG4ed
lynT/ch/SXQfO2ZpaSbMEj4vr7toarQGr+bNGwef99sg5hzYChtVGtkBIYSO1vQKLcmG0LBXvk0n
u1sZq8+vKuFcqndm4NMUc2Kjc1e1sSbvUko2q4wciJgFqnm1f6XWqa+WQqLtVfZkTYXN4V8pZ+p9
W8BHAeDjQzAz7DSoziTtIe1SUeCFKQye885sHAP+8aUjiLVnt27x/f3gSGfHQ9xMdS6CKc6rzev1
KFa1Hj5mmzB+eO3ZbkmgidQy9jM2zgSA3c/dH6eJq88CgVHj5peTl9WChHwjmNgLkVHCkJKrRBrs
pnEBpilDpQs76YDgJP0+riHrUi4xh+DfnTj6/zXX9726sHfrtR2837ngNakOkdIerhb1d8NAklJ9
gS47Se5dH3oL20R7b1njIW+60u8NdO6aTZQpFdaLc4UEDPEE/vWtXfiA/lJftfP8XIP/dVl3Y8T8
/fgVC3s3KdgofE7Njc/2NsYIsWHv5QKeYiihIddxcL5Z0V3z+L4XQHog7ElhqzsxbIrPo+uzcr5r
2fPTD4otloiI/N7xdcVself0oNiUNk2js/UCf3gbWEpNwgM2dCEQ3eJpi3NJVNvlTSdLq2ZrAqA5
460t+/+T4YvB8Lu/yDiwG+XWPhjwLy8e7VeP7RjUHNCNekR3iC3ufqAglthq+ZxdZOvbBNFvt/vA
CS2374fptE4sJlrlkKTPiWzNLBunQhW/vaoKT3bC5JQjgpfTGdp3mA9LMgDbEja8/eFpD2h8pTM3
1LgrlxqLJJQR/bq6WDFVsZp5/QqA/vs5ftLxBTePZG05y1a7CldCgsvhObN7FLAHSI1uq6Vml1lf
mqJNLt0lP/nK91i1DnefaOBEH7XpOqfVxjTU3TvzI5olteDpkcs1HclxoOWF9jlgUsiP2sdLRqYE
uWLP2dqLE3YOKZ8YZOK4W+SsdvElpBz7jp2wy+2yZKnLbRNX+V3x6ymOd/sm/yFmiBwGW1mqSkaI
MKHEOMywMeFgx4rL/xvgE1M7MAzpImCIuSsKHkFpyFvJfioSlnMuaUEnMzqWFG78OLWAqNSyx7Jw
FuVgn1pLbw3wPFUXxbC/DNFKfNZKHDalEs3jvZma6H63McpvEIyLgOtP9Xd2eNxJYdGlxRsw4SMJ
hoCBlW+r9BRYznC2tjhQP3yiwsH9ImflnsMHGUGq+IRX3t0wHbbO+RUT8lDk2cbOtk42SUIAjOc1
DliAzvtmId623c6vuudoIGrbC5RzSwi3R3Gi0Cl2NralVnfWO/DuUza4FSG4XsCFR5PlSXL9qsDN
MRPdiDip8AtNsJwCn2rYhDAY2xeo1P2X0pUtxfuekGTO7a4HAWrY7ZN8owpRPBn+KUMpAU+AJ9wM
myTax2CXzPoFzCq+dXDO21eGJHRnPpBUdoMaZnRBT8jUVoSc6jzHQQl38eqxLKBSsgFHLBfbvNsU
LFku38FCraghm0iux5rhlJeUWcoOuNyWQsa6JZayTResSZ0metGbqL2mD1TTMWZ6TQ4o1Kt5r1Wq
elO9TB6n0djMrkxuzUx/lmOSHFxcK7HjB7+/m+fhImEHZcGEHehvMd9t6BOaRqhUwHbpc/h1Bqil
OTk3CxOGWIkDQjcgJdFUsuLpgu7Ra8BCfPVxUe1+biEIo2DH5gi8NC+ieL3AQ2dKbG5Xmih4FOgE
npXKDul5A2WKquwxDqGEUCWCa5aIUg0NKQwkfiHtKKEuybj/Q+torlGpk2dsYdxiTwiid1+QzfsK
j4cGGGQnM5uGXDnhLItPetkhS5aGq6A8xvukSuGukRownJbktv3xd5p1rQVxIdiLSsc6Y7UICOw1
6+l/IxMv/l1y019QGGbZyMD3Oh+e1riui6Wrv/Ehb1eHyIHwi1Yd3bc4FABq8Nue77vkyv0BsJCe
OsLIVkaBCG4QR78cogoNkJQDap3+IpYZAfCg+ZL9nyxn7OdjNJDQ3hoIxLuBabdDmeuGM85rVjgo
rk02nD7kaPDCul6ugrNznMlRk7sIYFM3WV5m070QAzEOndSja4KnhDZcZsCS+edfWR1CYR5oq5UK
qFpi7K1KQEiCxfK+5DMgybKFnsIz8clJaKrM/ztIv7zwq7PnnunsXxbFlFhJakyZr2x1hxAPZPZb
aY3URgiBAD3lDqFtqvfjWTECewT2uv47ORJTdX+mThyjEMjy7pX0xiw1UM1GDWpEhMhlhHesGdyn
fsv7wcNeYQslVb9SD6v4qGg4NUVSI2Q1e4323Aam+6r4o1zrlag2i61P3dgzHs8jKhgP9B5p6Rwq
IKTNIctpE3NSc2G9dv8zg6qDw/mTywsEYlOs6Tsw8V1no9k1zIO16do139bfeEJPVrwwrLw3+41P
oY8ctY7yRlgRbQ/mukjIyLFIFeoe1AH/n0GleENqrr/kIrpGyq6Qh38qcEwrW7zQ+tqpk7rT6y09
P9m+4gUdT+/yG6bPxE37D5MaH9mbH5kBkw718vvpZBhCLmWaBzrA4c87MjzTJBCn4vDBlswdD0h3
Whv8ArEoOsmP8TrAy7UbY8Bt8l5MsV9T40ian8MHu9pS2dkFhZwXwm3qqaY3qvOD2WGuX5RZgyUI
9nsgksnK7UKeFrQIhRYjBJp+z/wxbBA+wgExvR0lsu/FnNzk8yM0lCzc3OhQ3H+8tiLezIQbTcYI
jmfT52CaaN+P55GOAd2fJ7EvWmUDsvAoIBDWy6fGmlg1dl9eDRF1FsxZgRrwkglhTz//xtfMxNun
UEmDpveeVbPyg6GS4RICWcp+4JT0Yxh8M44lley0o/ju1sEIcVsosw6fHaP4Tu8nnTPzjYWsQDFt
ZxUJhRBdwHyInAZiz0a73r6P3sGuF1vEHcCk8INlMNCWeTJnOdhMtlH2HFWqkSIuYvmMVZDxkq+T
20t1+iSK0j+dMuk/RVvigh7kjjQaAvlS65x/10RHK1tSKOnZmVbInPzhox34d8LLn3Cx/h5l3yQZ
5oL9IGJdt80KK0CwOJ3/dNBz2mz4/duQ95gWo95jzvjVvJKxPvJPCFzX5PMqGCPsRS9Dh3D8hnsj
QFevODfzHG7E85akvtJloSLW++Ci1p6dC+lhBcADa8Qv3DVkUN15Mi+AS37ZZSpbzuAbugi/ovqd
cwZ0Niuo5l08ERIMcyrjvmAaYcJEXI1prVyGraMTKLmihAqSiRuTPKXIhhJbM61fApzCRa5QTTo4
XIlzx008EEkg67tg/uVBgRXBn5WV0scN4f76i84/jqqDKthpbbVA8xTrxZpRjsAdPDeaKRqL+0c/
YL7wD4yLCaNlpUvsu2Ld8i3dYY9PG7NFik/49TLOa1K6A9+EVqdoZ2k6gk+8nFd8GYgXTdwiW3s+
ajTOccpZnMGQvhNGVeXMJ6+Hb3XQwnFGUjG9NU8kURsnHrVechqLB1/Yodh/Rh4r5Ej5HQJu1Yxp
qypGBMVT9MdDrfTDNeCEF1c1V6XtkxdgZBBhVofqbv3sHAp7w5KOqL4AAzfICOG+P0fYiVQT3AiX
NMDdn/LLO2xZrgI2KSZAG9sEdkWAabNEdFnB8nExcVgAEsTPeY8qj7/hloKTIvZmI3n1/BeQheRE
lu1uIQZC/E3r/zvoVBZgAMitDOJZvFtkvI7qFqZ3zluCydXzMWEBUabyHIVmtgC4x5nLN+VQTsgt
Y+G/zywVRAOPevl2sVsCjCd/EDYROwTuxM2/dUV9p2QVEsTszutdlM53GEjRLz8+cJh0O4Sui5JV
5TCshAzBvio/EfNFC0jxtq3wpD5jMQIAteFojvLjrheBXKgUQ8MErTxVB2MLIBq1boLQsITvAFRg
PDNspRI+f66we1RvDRyWpjP4eSwH10+LgYCAWYI3s02JCos4PnTAsFYGVXccF2C5HfRaazfPhlhZ
P1E8Twh/qcfkEjswGC696zxqq6O7ao3sWsT0NBsbvP8uD3SS1dayr/xdwsixU8D/wHIb7FCgT5xl
iyn7RZTSpewAc+YjUj3P5XYFbuFYzBu7TYIqfzV0Dj1Ys8F9XOsnNnr8Lo/pQNz4W45mVR8JwISn
TlY9YoBzPBmyabtU98sEyxfWrIsE7mxJLdfzWjRBTm1nlj7XAb0MbDBeMLZYaeO75oWXHjnDgJcL
r80sGbMhQMb/B2u5mjRtNE+MLGn1hFMaDx6Kh99PgK8WSstG+RPxITB/M1raxUAEMG4W48OEIaLp
Py9mmYH6mEDMPFbBjU+3YlHFqZvZxAJtgEp3vg2Y6V9pD7m2K4gpRcZSOZbBjs5kFxheZhjyc/kM
1qvwOs70Wqjxux4JZ1vZgD1HfCDgZPOYxCd916k4Dud9nN8XMcBy+FHLmnHPjhAUfKdYCAYIefcj
7dxINDudLor9jp81QAgPpQoIv5es7kPglzgNVa0xIipGSVVMFk13Th2OrZxutFKw9sqdD0Gt/sBK
KfKRct80q/GCGhfiHe3TqJuaBS2GG37iN7nX53Ww6wzVO0r2x6+g5Spfme/J95JMOtQF8jTPtYTI
nyMWxhqSSrzbb7hSSQ5hKBc7FDil6PWlPDSE4k3ZGMeykavBHzfrFV6xlw0JIkQAP8bPh6nuPcNx
ErkSucZzHT3H22oLQCAWsQfcPT7kCEEgBqTsU5HPb6tGvHYtJV+gdhELuhYqZVasiUxJ69OILfg8
pHzVHhWWFtAbCadwEecCiUHfGwdcMzaD1lKF/DfihweEE/jDk+0G30u1+007WLmRjLbE/I9XKohr
RApfgv25OMpkaObfy9de4L3a1XavJlzFLBwUO0WNrwFxhthVJs2QmEIwcWqBI4mbhCtY07eODdVC
ru0akQGs8bBbWGFbqL5fQXsPBgbP6+FY6ykAnWjosWtVh+cWh9Y0TwBgBiU7X42v/mSj1KhdVzYP
sGMW623Tty5meTc8sfxg3Roph/zbPSHdgNis5d53TukBnDWlaYppj8MWjf5z2NXIjyCTNTN48RUt
0Ezy2E5pXTyq5cfP3bRAY6C1w2Ax0QJNliVGbpecNhhl8xQvrZmt1Ib3FN9ZIULOiAinEoRWbeNu
eV7WIVDsTn5JCtwo//Mgoz31k+1avBNM0y4LvlR4/72geMjV04gVyV5VArOX14Xjg6TLLdOZOeoJ
PKz9Cg1O32PNdIbOv5f5G1js5EWgrO/fy370herMb4xsAp2OfDFh9TeaCr3hnXxqawUKaxC3EK8W
hlDgE26ahoDyk5SSFNqgIkG/IbAJLag+W0LL4xdzX6aO76JZnrwywTN79qM0fE0kum4Jx5smIKwH
kjPMIeZX8TF8OhMuia+hUJ8xi/iNc47mpD+IgR5UbGPBTnQEnPR3qFtk5dBBSIz1U0cTOSV+qhcs
dsC/FdHLNg8EeTTqpzs+GZ7fBnQFzSBmRg7Vw8pbtXe1ZzSB13wPQf0RKOZjHQFkH318zIddK1T8
WE9NkXjadyUGtfRRXS8DB3zMFKufmdxlPo0Z801Q/vowgzk62VODP/wQN99NNLixSYLd1bnXb1e8
SLmEJSWFIcAuP38ZYrso12ic7qLrOa0ZawUV6iCNDWu4EugX7p35yZXBEdDtrn6wYFb8fYdhKf8k
mQzJW0pg/NmSJeo2fuXQotskOHJPNRpUkdElOnbj2HzEBBLP/MAXW/3thYoq4YPm39kbHA/cRzu+
jczDB2KngCNHf2RmMndiVf4xdaly3UFfvxu1ieTQ5F2Aj2zI9E9W+l5YLSQ5CmLF9UDwWxAxT3cr
pePqNgS0X6h1HUnnniAPI1c8H96/pDqwmCBqYacc3zCweOVp5TtjvtQikVVZt0nKqQiTJjtMw8kC
1hyGBZVeVGsqGvkiF1v7QYuYGI0mp76xfPivVW9856VNe9iXgwceqCyfHCrvi+eCdH3AY0ZOExO1
a+P967HUk6v78dtMy4TLU0QmsKLRUKrkCAqTkKGs/qRl48euUG3aEoQ4Ofgig+Szl6gaVBLHBGH2
Em40zXM+lOSX34IS/T1WNCYkvOGKg9gWfsLNb6f63T2cO1OfXxZ1NTVxtASRVNeROLJbqIlZXRBB
t7m/1VvgE587aBqJ3Yh7j7+1YQ8OYx7BKpMjziRPu9xAgbUEuq16xmQnBRJ3iAjinAv82LX78xgx
fnkLFCXHbAd7B6lRy5/QgY64erQGrdY8kLTy5gsShP97YwqErH5hfLS1UMB9XLqKcEj4MIKH9U56
sjvWibGmzY+73TEapbm8PtVukkgdcLt1MJb8LGOpe56K8dFka05+/Vz7ewRXGW3moYpzNZu25kEY
IWou81iI6pec8s5ojLVril5BmVn6BTAKhPM6pal7T1k2PPBAP8TJVrr1+mY78aU+8uafGeFl6j8F
fn2BEbTLzaLfPFVXLOGOW+YUAaM2n0MgCYrg9EeEr82tBUcs98kgIZubq8e0WRW0ByanGVgqZ70z
q/UB/cPLTxF5pLRlPuy7kQUuBfNv4f92+vRG+TBPnV+b+/Rijg0QHAvafObVlMP585SSBZ8am2TG
1hjemMLTfuZAT6jGIyBKZjdrAHT5xXpVozIgP4y1lbcYJ+io/tl8cNO1RvjMwXRQ8IiNF/Wur+sJ
kt3LkC5DGMM5Mt7TxGD9F7JZJRL7rKDnwOjIFNTJAbyYXwPkrnD1cCw7gZJ4mNuWIQrEQoQsvbxt
Ut2mKh2/4RuEzjEvPhvltQH1r+68fJUc6T9cRRXrV+gWeSCbyWThVczzV0cWcA9xPOhy3H/tgSLo
AZZ1i6+/1onWi3KUW0MlcwnNW0Qiw5oGwEDqUAQMPicPjF3cUQB7TaewmJO2hpxF/Ll92Wz9wCbY
Qof+wTizQsub8ZhVeOX9kQZG+f/Abb1jVVgaBr/53Q7e4Bb8+S/kjsSRdDfFzVJV3FD9XWrA+MKb
/G1gbQ0C57t93B4eDt5eTclJCLwKBe4lGIO5sj2/qD4QuCoqzQRSKuSar6CgMwq69Hy8SV96YtNT
ByWqNwlKUkks4BgPbxpF6ht/pwKp8g3u8B+46AZz7DCXFTV6cuXYFDOcnVunsnLzm13ohEAOsmYR
rh5tdiSaIcGDmR7gIIsILX5HFYqP0Tu193neIf8x3T+YnTMq8kOIKviof3lYhSxhaHFaQQJ4bONE
EA15eXTqJpdoIhk3lNziGtVztmwn4yJao/SSxkAxs4NSFcA8WMI20J1FidrLexBrHNsfFSV2louL
dxDpyJYoQNcRsk49xjDPIw52IVtrqBLMkV4lBvL3Y3YBOBKhvnvt6Gfc/mwENSbvpPygfmFW0+ON
oGffMSLN/Bfl2wQcyYdwHe8sg+eIIOc9VCW/Y6fHRsXqRCn+8iHY1bZPy3M20SQspd43EcktekYl
IMmLeG7BhOpdAhNPOPKtNglPod1QyXtoy7Rj+l+6FmG88riiT8/5VCG+9Y6umWQxfNgltoJYljba
q9jipKdmDmTkGhz2G75EFkoXIs9nK46F4qD/1Xou5+SaVmHyqD+fHYyBXs1hL+wBfa7Kh9eKmwob
rVQedZ3s09pbWGT+qIL7PdqFnZ0xS7JkFvb2ygE21Fxmsy8hNkg40a4XaZXqNuO52xRPIfHSXMKu
VbDCU6qGSh9ywnrRfzpcSZ+xGn4SA2exb6wBUTwQ0kCaiUiHzCpZMq2rDagTGpEIgTTmYFWLuJDM
31rV3hKwdVEDw5qQkC32xFZG4TnfVPDQ/9riAs0T6rZZvY7FlFKpcpWYdVaFZ7wfpqKBqJv170Ad
zkxtIJgqkJCGrq78NGTHPj6146XH6YUyuHT8if9VK0KiBPrKZIy+h79mK6Sxl1/lqNe7rA+8+/kV
6l5aTUSUtdpKRaX8tZv8WcFsxOE3dsNOUVvHtBptZAVG+nuKU5JnWBl/qC7iGdl0ThdzV225V0s7
adWQsYaJ7C8RTfDQJanLPsJf8NHitfBJnpU7H2d3e4K/4NYmNAlSBtMSUDffzYrFySNkYixfXjGK
A/je9uRu5Cr6oS1Lji9ykVl5O6N2WllyMgpkCvtxyrfpcxgjkourc6Mg8ojdlImCVB6tpWy981lQ
wGzgJdKFswJVKYO/WPP24cTYqb5tYc6CzbggbYSXl9hfS+LLhofCljXAE98m37QeIPV4nP8TUSMi
BkbKjl2jcdBF0GP22RitawXM4T/j+jRiVzIt6v5koaw2Se5bskWWdEUMzzcpU9A5H9t8yxcTPjXE
LLFmD1YU8xaAUVynlIIsGoIlCzr9bKB2DvGgjoYMe3xOIwDUkRVEBsCR0oicY+mn2xeYCOJ0DUVQ
rB2t3aGk96x2YmcDCpoWi9CpYagU1/9vq1CEB8lxOSv1lRV+GWzc66pciThwJbe1opGZCM3DXhX6
HHwdIDHcfczz1H7WMGIgyTPG2oqPDqKl08Fw4UouDFc5YeYJzVwZFiD31h8+GPd64SudmQ8l1JKz
p9lSnt4MoxEXpVSheEwGVbh8eQxkR3UndFu70CyTezTLDrVHwfjFBbfB7EhxA1WJ6bWIX+2Y/kkL
VfTYGTZnQaNkoX9Z7ZrgfULmWdLAaWrFSXzpDQc5Mwv7Br/NJgej5m7p9DxHqnzrmHN5hi0SC4+8
SLv+pBDkQFCqlwQfZXtV90QS6hG10prH2lH+lvPdbXHTUY7gCfuaOa4m+2/PucaJypya/Y0xWXbu
b95nXjP4Y4q9/P/M+1JlKn0Kb/pO2D1sK8P50V8FiRYv4ld4yQr2VMqtSALo6S4f1TimIdhDS1Oe
pUuudKlxJy9ll8iYXdVlRnkK4KY84VfHG/cwwHm9khUSs2i+vDzW/Y4PREd09+zVTlJB0YcnGtBG
++atW7GbDAnWHJuQ/xgvvBHRbpbnTkUUJQd1S/QqPDbf9uGCtk43u4PaOoyr9zSYaQ99CEOmEKWt
8gqFgTt2ub31j+fDP61sHur2I9/SJw1IBMXIHYx2DAICm9A7nY3hcpPpWlCFXv/9GNJMmGY+RLVK
DHUk//bjQivvnmCO0SXguRv6f0xP5fgO8qaH7xB1H3v7pGdhnI8crrjfmZGO1kgiGohWOjQJtEgi
Spu4+K6g5S/Ct4Hu6d+EjHx/lAF7fC7lIQWYhN0JnCiuM7Z1oy00xQumk8F+kZD8atYzzw3trYst
hqH43ozRq4bB98YHkuXtbFa5LaZgry/Sz4Fux6S7M06jCT+zyVaf1RiHJdWRdcZpBfv6Njn7xI9B
yt7WvH9xrB8dltNnUuSVVFCfN8SZ4JcOWLra63MEJ+duBwFvpJ5UH2FV+2WfMh86ihAFRCLb0WYQ
yFU2Twb5TJHPGvPR/yYhynH58Tqg/FBPmTcE/JLv2MHEZVPONqKSvrO9j0c3KBU6FvdU53jeCpXr
EZjJvpckAw88qgjOfTwHqKrdMMpTOo81MW77jDaUcJaUhI6F3z1yLtVz3SzfbcyEz7IXVvSWGhIB
pewk7JMZ4WWExyOU3Kywg1Flj+H73rwe0dZMzjg25sMBEhf5c5f94nMmqoxVwQPMRIYtDmLsd0Wy
BJedDVIiwir9FDI/X0tzi1V18LY3S11A71+8AC4uBN18ozlHowLytUA9VP7NJjMIvSptZ03RFSIR
2xeyF7+9QvKD3x3CbBH25I+E7RGuIt5xs0Kh/zqPiIpzKGfbIdRxq+s7BMP+G86TjmiPzW6kC5Bv
5oY5isQoIMq6yC3oLRo3vBPIHxuW1gj9302m2xdjchFdR7DhElnhQ5FN/G7KO7DHpkbwYcngjcIm
WbTluQD1Fje9sGQl5V51A2sz82feo5emFEeFxIJ6Kyk4ONv3HTRt72x/LAUipN0K/Voy1XHDpB0y
m+I7End+M5I8QxSiQLz7n6DU8kWVsXPKBCovcHBaBvjG8u3mf0k1+Eb756m5yOlS1GJr2JhzqX7y
r0eTBCDnzP+jOipPDrbekCoM4Kq9AkzDKeSCy/Fc0Zmf3iPNFSKFfpKjeYo9HhFh0iQVjpk+S/Fp
FXzt8q6wEku1uI5GkwcgpmTMVVz2TKfCK6mf/ND9s70gU6YDVRs2ZzvVQa3cCwKbAVTWofjMYkEA
KyKtGaMzNL6cxmIlX6QYpmv7IRBnzPpSYut8g20sYWSwZoc5R9HAmAkjBWve1ucAlEGnxYOFL807
D2yf/Pc+/bVLplSfbP4A2pbYiWi5q++74oBZsPpXmi1y0Myw9EOe6dVZS7fshjt7KqHCkCzL2BJ/
Mvgh5WamRLvdc++b5EgMVltZrWatRryzYMeEcd9B1ipVCvzjNLEGV4cI1DYKxabenhFDk8xnB3xV
KPWXXbP7NvcLcawZuglLSZHiwMwhBulSgzmwvCmfclGxXCl2ewc8zxHXgojkOM53quciFsWjzI+I
/m1eSe2G2OL2nwrMbxU97f7gXv3dGVll9CmIgkQtnWyrv7zfc7oOQ/Kf7Vc3xG3HJYf7UmF6t7Mm
2Cn1nMxRwO/pNO1komH4noa84s5XCJ29bb0ChHZkEpmpMuo040tSPtDBir3KttV0y378LogAEqnX
o0+O6L5sFFCI5sL+ZywXFhaf2StO+FTAoZsEpSGmdWn3p+oyw8tuaAmI5C87TzJQX0MsdotNkXCZ
tIDm4n/VwRSG9xYMadlIwpXlgcBwksGR+XO4is3ywBPiVkqg19DsAamCtxZRKqk6yFgEQsOXhgHT
w8NvN90hkofVNra1BxAkZ3jkkm/eo5CclGNfN+xqb4/TZAdaDFZZQkYqx6eNfCE3cy/6zIfz8n7K
hbUo+MKPbY74XJUzoylbfRlvA05YQYQCRFEQEPetEEOQVYlXXw0EHObdURw8nveKwmm3SNkm8v8n
QefBWgpsJWE/ppcIvW8AtKnqy+jkRNZsMF/mWJQ2FaQ8IsvKlOyph2mRapH3tGMcXXOJlGJjhOwq
7Rb+KYQJrXo/1HNCKEH0YLW3/G4FV2EJC4Zamru4PpwI0lPVqk/pM5GYvGHdmvEXwrPcIKGOL3YZ
vTsVCSWiHk8FFeIvYrt546dPUwKCgLC/fFDSqCL/rP/ZItozLfzjdxqdLMQJ6fLnoJW695O2XYEX
7lVofHVruRCi/ZFOq72KhVbDT/Gn/dazi44ym3jGOBuQ4da1msSdAjzTcxsWoXVgzju/AP+BFflb
vteb0Ck480GzcrBzgCnJSTv9/RqSfzld8smfN3EN1QBaXdj3qugDOo6H+Lpy82Zh5PnOw8mfEfPP
GQD6Sc2Fm7UrHHNgCKr4RojZcpoiy9nvyrmzMEB/cWpIuerzAO/IpDoSXu1Pq7TngYoUugcMnIjY
NDUieV1FBv40fPIGq9ryRANyBVUcPejc7OIaKjMh9cqHkZOVk3nQFjP7KennpkoqOd9g0rNu1D+s
sLWRfcsO9pDoKeficCG2W3yBrzDwMUqY5oYARanQtHpwV8kLQfUhhJmNA2H6muc/WzmYIMnPMKs2
VpJNCXkFL5F4uHFU4oJdJHYQYCj+uKGipCEmjyI5fh0ajfQ+AkRz/y4C3cHGbJTz7OGZgEu45/Jt
csjhdAmQ0SJ7KZx8BgJdfRAFPpH1F9nkAzpmN0iUomlCoxLL7+4lA+xnZh2akAy/sQumR5QByWv2
5NK+bfJBkjjZNcnoKmVxPGW+I2hhLA5DEZ9+D1knEybzs5Cl8gWdOwDOe7UCCEhYi5by0usCK4y6
bbXl8hc3vvPaYdhmedyKGUpzHGUN+/InKe1Cqc8oCPSow4B5FtHvh73dza2kpbggHqsLygf/Gw7h
iF3ZhIdPcWEqZva4rQy5loJLyqJiU5NYDQJ3LPjbwVMTQmJpboQkqdoUWfyarltltQeYwdwHH+zW
dzeJ4BNsvgjkgYV8OaJvyrDtsY1zOCwGmVh3Ul4TXCttHhxz/IXymIqdo1jrpGDnQpVCRdfPc0h9
EhYw/GQT08GyuH8kenCfBCcA6jtJA/0HESh+em6H/SBWqO3Oga65tKDUqiIidOz+z63FzwmbPfxX
/FccR7lcJjOhQ5BCk9XG7lQtgP5jjhg2C2iEep3ktrsVMgzLVy4aH8f9Vd2UcO3bBPnulSityqZq
VqW/4rydj90vuLr02tR3btS1FI5Vh9VYutSL2C5HECjkJOTCwm4u3L8L2QTmm5MxSay5i95P+3Vs
EJj9i0afAhRk+hsK6uSdyPH1Q/EwbjH11sf57C/TcRNYHNlNq58rVBsZzQqtgM5g6f82eOCNMg62
PVLbiNATia1NY4NpzeGIseJphntY30SNMoEb9grny4b97DPv7FYvfbpy/UvGt0BUTK5PCa6O4BGA
gZoCEVt2K82mU6jIzmijBGV62Mid3Ou8PQLllGT8pzLwHW4B/X+mcaAvH7d1+BLTyHNTCC347pVL
uII1qgm2wtvazaV2nCsHgeFM/zKUGNLM31PaBDp8GwJq1ZUZlNxlqQ3MQL2Kdfqb/BLJuAqYPPCL
7w29wk+N7aUc0Q6soe64Vf9B9wyprECYnOpfRK1OKzzGWgHkhBFW1iVlsaXqx+ePZv2borG7tnmD
ZvkQWmKA6FXHwnwIeV13Fa4rigZ8uZi6IQNBMk9mLDgYf1RAwfI9kOtWTpoW+sxwzCO33FDJdcOz
rAve928ct6vCOn+zwdfF5vFL/n9VAzSTe/jVHi9yj+Wl5MB0KZW0F+6GdCL97jeP2h6Y2IqQ9buh
9FoZvcCQMiDSPJzzqJU+6n7krc9ewBe4HtHVH3gNhlfKKGoeeHNOhOpyVpiJFI/GTuIxp45/gcHp
dXglUHB4DOi3dnNNdEtMDjJtBbWbymo9GfU+EbzssxO26QxxdJ6/CSKi53WA4DVUVlmo7ExRpm2R
x+FysNf5LBnMNYhjaUiznQcTXsimHHGPWZ/DUv4SJBSf1OgWBY68AMXe7Yk6m/nBadKmXPQLuqQR
FqzEdWg9nGuQcVMwFCddwBzz42ZhU9PC8lJHmKb1x6oQBSbJwMcX0si4Kvh2FVOZpp/UnfK/2+gJ
LS7w3dfflRyh2BL7Ka86gB0eIHdAtcHNjIHQcJoTRm+7dmNlQSDTcnnYSFUDxiTNeV/zS3+jInYr
uTr5vqJyi4Pv967fXI+Cr0iXFwwZXrM3WYv25dsLOs8WjLubLE3n+HW0wB/7WokotFXy6mxnAYCR
Fd+cpT0pxEgqybLfkLNt9/hxkFb+hNB1+Cf2Bxya628E148HF99/yyFHDJ3FcFI7PrPyA/T8dCUu
HmvssHHd/zyfFCxJIKfqSBJysrjjD+DesS+bYDvgEGr1nreKnQZQGFMwqN60sYYxgx+54YFmSxvA
gUIKOv8O6fWl6idr
`pragma protect end_protected
