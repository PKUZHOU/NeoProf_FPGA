// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Mq0HG6dmt80f8SUAow+vF6BGCX+Ikklu4xhtgxi6XcDiuT99bMxfkDlxyZKS61UR
36KJjPQytmiUfiRUQQX+G3M8DnSEWPilMdy5CnE0206mttYOM/P0Jv8ybT2renC0
/AGtuLOKaFNYXy3rGOu3P36RkYMDQv0dyetMliPxyb0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 91088 )
`pragma protect data_block
5d92VhGUq4V7ip86F449BQt2lD28FT8TMGD4RI+W41n84KHzO9GzUxWqHFSnrE9e
33PZp9uYKSodEsSCCdfVHQtM1Xs0LTJ1anV4dgvJ7erfPKiWG/T5YqgrEaUZLEf7
ido64V+3rNcF8FLbF+OptzDKQWr3VSWFOvS602G9KdnE2SiCdmBkxNd6CdnjaysT
SmKTxcTLKr+vJOUrz7b+8B60vM5Q1W+sL4IG8Ltv8BmUy0vnOcQre9TFYMUy2qGB
xwNNinNMfzUV/dVwIYU0kr8EPIORtCzJZ8zC1kRzCzgMx7d5vfKx4YyaF1z30q1w
gnM3f7bmYDfIyOt+17C3SX/+WtTgxTxiISrewOqO1Tnybae9siZ8zCsBBbGF02y+
5YFgmvs2jAUQ9CnuQe+pCvoS6b6n/nqce1u7Vmtvb+HUjXwRiWNCpmt/VCBI6MtQ
Oy7yNhSS4QTOKhiy8d1yaT9ZiSBt4ehGbgLa6/xdskGlRbs2jPX8CHWv7gjHNv9I
KkW4hhd9DvVjhz4JO27YRtav6oxXe5l/4w2q5RQtBJbGGJnsWDFwPNB61xqUv/Uq
oWZSC2v1IzJfkDIbQ9h69lT9p+d57vLuFj5bU0pFRBFDydQ8FETTeDPYMzJJEobD
ZbfWlbs6DIsC6tfVwgXW6BTXfQlcg2kU2VSUgUiOjtwTStnmCL58Yci4M5mdDj+w
OacoaBG57idvv9xpjDVxdOlWPqPFJkkGXvVqVMYFMBqKLIsVVk2v+5iBwuMMrKKD
WmWZBP7qHO77rUj/YzlC26M9acpc4jopGn6xGC8iWMSET7+1rlxnBZr69/F8JBZM
8lWuYlwrMWN0C/5riF3zhAx6rVoKeVYEQt9wGkhWqaX8ea7J/ocl/isTAW/z7YH1
yLTwmihvGp7WDz/I0Cfe40Yva7c9f0/obcruDk6txG8kkIMiLmFwLFWfJlZfScHY
q3mVurUZAu6tAJgrl1LF32/q+CX+tIgZfVlwds49+TRNY9YeWwEiewSTn6whAm+3
TU3JHuD2RymhXICnsD2MVtuLIXGg804sS/sKRE3VS9Lv2HTgJumkYTIjUqAqWaQ0
T8My7WFmNm+CXdufQ7fgIcSBa4N+4ynOPtVIQbs0xxrZbKYUC0HWyBOnMvYFrEN3
u9DnTfeY+D5JB9jh+MS+bmBdUkm9GDKwOUcrOxeE7HBxUMbHSJssR2vYmsDaMXbc
pqUM1Mg79xZoSTvBymGPTZCpj6O992L9ikXrzo3/pWuNAC8te8681DSPhw6c90bY
N7fIdDq7/RjL9rJl4PbnfUod+KQnnLRpJ2rcCyc3YRp7pLGPI30yZOwLBvozUPLW
Lx0SJxJpK7w34H1DjzsGDxyAupdX3FtSU5oQEVRU5hjlGwJGmWam9iCEuDtEgaGd
VQ3Dsb+JyUVRCd1iR/tECQDT/Xz/F1Mh/4QFmAjTGkHoRf95vri0FLvfKuudZjUx
qark3Adc1S8JMx+lZz6E+CUD3l0bNnWjtEhJQ+qE+Qyrn2hFZeDeA4oqvaPlS3Xn
6MQajZPgOcYQVZchtjNTllTVulcdoVDp2ajhnDzP2FDV5D5iVs5FHX5tY2v7iELr
TTv9hdU2CBgeF+2d7PNRyRSfoBgQatl7TUcRVCHKEsgIeiTmr+cdQIQXfbIqOzF/
D7pMVjIX22bS06QSjXFPu30whJ0yaZKdeUXCD91TlH1Wy9N/lU/AtC8DMm2CNyQz
Xg/Rz0pzOwTOc12QT7GYquhUX5QkI8m2m4XVgpz0ciOTGrRKhu4yV+mh/F0tE4sO
Skmv+zTW3J3WJDrncfLrEuQK7vP1VWWxEtUKP1bdxzrE2rDY/0ZGfqStdOPWwQ50
h82WslWtlmUzZl03LYDdY9oC1/qhrBIrqgO1SflE9KZJq8vUOOCzQO4LKMhNEdpf
6RUFShpS2cgf+trtm8HCo6KPoNcgzQGCzRsQQcZ6mIIvNdANSObqv0be0+L0yFso
saYB8Y6fMC7m9A07ONluYqnYV7WTQvvPbTHugjz3fh3vqQBcXLHFly41dXQcK7z3
chnt0RziIZhdQx1CRbeh9FGzRO3qC/Xt6apCNqBhFpU0m2g6B9D5zHvonvE7esDQ
Us+66KrqYcIyblnC03oyWRhnwOfXWVl1vemsH014X9EhMefGJs35/Y0JcyMXPXhf
flRxqd6X+WjIrmg7k3aH8I74NuJp2syLOUeUIS+ohZtZ5u+hSqCS1Jxo8XC/xziU
rodeBoavl5iJQEX+RxccGguSAenGUtEZHDfXC2jj0tG41ThwSYnskNT4oEsJMzQA
BMGbM1X/P4QkGabEm4rj9wExwOiIir1gqZf2nOJs8cf4HyRlMRo3pjPICT6ynMds
lwFGveNco9ULKwfKmMdtHaHlN5Q78i7aYS0aoQSfBRG8HLLNQgioH0iOjgTWsgK1
LDYM6/GgLuAUKnZjYmXdAzSq/WsKNIdzTzrkhPgfJwpY2KfpWsImEKSTeGZT+m1c
Ela8tz76Rh/GINZ2SS70YayHzjrzdI4PyAZxGpNoF1edmxiEIFYoMfTSZYEisZHn
lOZqBW9sRlf9LR3YJLVO37akLc1rGjabhQVurAfxCuu59OK108O+Ohdxf+YoMqYM
oNaoniUuh059cktDy2mlbxDpjQGo/VWJROzhBbab2k/wOZhMZfMKVDt8mzD64Qz1
5UTkL4d7bVV5gszOZbriCPW4NnW3kMr4Jx1gQ/bP3ourCxpHsWp1ZQ2H83Nz6Kas
PYrKOsDAZtdNi1KwvaTAwHD3DsEZ4MfA4NbdAyAVmNpsLgZeTK4CrtDNHZhM/pHA
ONIRTxRL8kUoufer8IrNgfIbeIDUh7z+JMAvkFXb+h7ohQ0/QxW2ASmFnHg8qJQC
Cl0CWuxP4m6fpJh0FWLKrundXUTlRU8RMc15uBskxC6fu02SxzROKAwbghOxI0S/
G8TTIDsf07BjHiE9SzzvkHyKHJxFzT5sdQ82cue8N2siZjnkGqL7Eut1ncd44pkT
FnZBQj/BV8AJXkvNDqW2EwmMIRRqK/gBaAZ8WvsGIOXey9N4Wu1ynjoC2PxepdRL
/himHD5FWulmYPKhalk9eGQ+/SpCDfqBaFMVJBB18LemEyCmxwb0DqZdrDAt2Dlj
HaK+U1flAOkdHKSLpjP8D/dZ7EDTaRBAroOPeseIFVoH6JD+HLgzaNpXf4ZheRtd
ZXw+th8x0jSNxVqT9FywC/s8rWp9a25xV3gTikNbVI9neQhdmRrWgjqOBbftV2nz
pfuCUxRLCgo9Bb9POG8RP+LMmp2mvsFu/7kx8AYzFalniL0aw3dLAjwHy1CCWmkQ
YajiB11S0cB5YNvbgQ5d6NoDAg/22bPIDvZRCVWDfckEGV86Yik8gPxN/6DKGSK0
bOkFqfMZeV1LCSVKHIYF0qEJEzr7hJfju5ajrRt3KaqsHmWA2MikZFSgoqx5WAvC
lrYhNcQ1sFsaGwVfZDpwlJ24JuB8MQL6Wtn+1/uxGsRt8vepRJhDRtF6YzI1UwzI
czgLFTpJfz6MjP7CBG/Vxku0lkuLXQuqgTwBcGA1FfN80JkQNSntSZqOsqp+tsC4
f4g1jlPV0z06D/OPg50Ulzx41abbSgPf1tiahImdOmLFiX3ZPMi7UOlLm49qsNo7
8AzC0irO9E6j2lnR9gNJZLlPZb4ELTaJpHCZSK8X0PzcBpCjEMR8B9L+eG/ic+eh
amGwi52q2lOTmdFu9L93Di3dI/ELKZYdT1cwWzCW+D/htWVWcrnkQguYg/q2ZdCQ
CjY5yjNkZ0bDOEVo8nwvSRyyKvAVUrcm4PT8agDXsGJVoqOmRol7oHoFBJlMYvfu
E2wUAWE+N+z+Z5stqwVZhrlhxexL7XTDJe8272DqFLYQdiR+BFjLJsY+8uXJgCnb
CuesLUcXBj5zPqhYpjJOThyTLx702amx8Eke+bslHXyXLT+4keEhkI61Doh0nFgq
P2ag6/0/h+EnANrIGw8zPRqF0od7993zfY+MsNBlY+9kkYefuJpGPSFuIyxeqtVT
30lzcNb4YXG2p4tN2c+Q12HgHOeAzc1g8qw2bY56dhZ6u0FUnhVOFTYOA3ZomKx/
55pok/XreLI8YiMXig3+0Xfo+HyV6fq0Id2dcepRCtT2AstEJNTiPjB/1qQpbnVG
2MlE1O8AHhiqYOK3q3YPO0u3dORgJm3TWI/uYmDKCovdK6+olm/GaPRR++YUKCDR
T4w4oHScH0IdyDGIwVYPfxM8LAEcbuc6aKRUqhVo3Sm7vLkiJ216dtgd3lXRBNMO
68JonHN2aVSz2M3WaseoC/fm28oYqwkqtOKH69nYD+tNefcWcooFFbMcineOb0hL
+P72gFUukmT9S0haaUb+d+obV3uhSrq2Y8R/iERbbrQ8dLB4Uc9HeEW5E2Bx1xga
tmqN54oFWl+2fcVeW4Q9eVhLBUWunVN0Y7t3q/dF2lP+P66xOto0IO3pHgjmg6My
ts13sVfGoRhp/8Sd0l2MKztGL2bMtIGkkkJDZYlbS1PuBbEuiuhI+488Pn1McqcL
lbeD+D/CjmE2EJmT4nSO95WR5m+Qt4zB2ngbQQXe6VNWmrYHo7Np2dKrs8M1j3jQ
B1jGl6Ps74y/KVQJqoJPJFWxQuAvXd0qXe9nDk8/yGIqUeHkBGuaIva68IP1skyQ
dS52AGEqHSSEjHT8JD/cJpTQk4UouJjgDsm3cMpAs7scJ8iO0yyZ8cPh+vRye1ZN
J50KY1O7pGx3yU8WP53bYrMHIlfvOE86oyCRjlOhg5gIykSGWDi+2swqedkQkzJD
ICkxBCCJ2hZBIHtVkdY9hT7HoPuG85kaY+zVSzMfRD6zYyPpfVI75polcuxnHTqS
QQC96xMwRxNYiNHXfXcaTpsVRzTiSzMBCahbjtLTFP+ZHJ4bjprcRSv26t3U2D3l
hEkl4cJXLScbSnSgG+Asw1YPIHyzqV2QJZEdcvhCKV8lV/G5DT+Ozefpo4BnQl2j
4JrVfAe5tn01oP0HXp8McPnGB/QgJWyGHlWVwxLoWHvZ7wXtQJxyTjH0W9db15sS
RwKUYP2//OaIDDSaY5RrgqYS2uvsV/C70X0SvKdow2XPvWZH8jKiU2OwxDiW0uy6
Hi5bwkFR0ifiVq2cWnwbLtmp1BpQ1Iv20Kx/sS7dmsaEVCTpRsx15Y/aquovla+5
6jGj1v0o4SCsL9rDhHcrBPbpaGAsRycgCg7vO0o0A7jnidiOsKWL+FDNc7odARhw
44oobm2EvZbP3bffoAQPzJzk3bm/vz1IfZXYxs5/SCTobs/Qzegq13eFo1rR8WKg
78Dy6YutKoazR95R371QRcci20rCPvTFi4eSU4Y93IUk4EjRRp8r1nXiWB0kdyc4
pTeh45Jbo6NGIjiJlADEgL2EUvRBBhgCMMjfoPZQVn9DDbP3AF5Gs8/o2pvfQpD2
V+KW2FR5BeRrwGR3Szsxm27+uMwQs3VZLjHBMx0KEWVJGfFFqrIMbl8GbHU2+Xns
oAeXxZAp1cng8c+V9jD3yVqlEczpTZ2dlqJAbUO9iPkVPWycTAvk0+QG9hrnKyh+
ysFgs2ZmGC+eAXUV3BmVf8kHqwQ5UyJG9Ghq0tR24ZnlFkVg6wFq7vix3njJIJJc
4ScG17S+4ymPfGvhS34vYVS+rjiJ5W6eMUFdE1Gp1rZYFW1Hvz6MCcVu1GJ0e2Uo
ZAqcumidHjjNxM9MjWUnYgtkn23ivQXFj3hdv+nWfPwPPyWkyM28vZ+RG8DjIpxy
O0QnCSISdsxtXwB87HsfuQ7VAvPMWLa7zU+QD37kWrhtQorfC6BO3CevlZ+AdNd+
it3C4b087wAyLNA5AQ8i2ZkYNgIDWdfApwQfROXpC6EM3DbmcxmxvprZv2PxBgGB
C0dj4YCb/FyhL6YCGHRJu5T/JxymQkA/zRWpmJKTjGiTSZ3HeXFNFxywerjOsVkH
ziLyXBrwEmCj9xUQIBvn7JeDfFkXWl12IHSZBKUl1CcEHIfTfZLdah6/AkkNwAi6
9Hdl5YKvR+MrQcS3aYVXd6tooxG/TnLzW6SxSa0cteR2wTQXsJgQdXZ+OA+Yvlt5
VWgQbkrQPegBj3+FssFzrHsGuGzhSEuJxeiDchkv1z53cWi5n8wVU3V9KO6weAvO
buyTMSaj7PP9/o/7ZcekWyF8uKCOYKEoQWTwGnA0vUmfItgj+W2eVi1Vs3x0QysA
Wv8TvGFY1B9lbBmYShyk8bAw1yacYzcCtVXhaBNLBgARP0uwcwhHhp90JvRUPvyt
aLKYGaHmtMX3lUGnVI5AQmeKwveBkD93fkidW1I0FYc2Ez5rTE/dK9Uyyf6KVl6Q
iRGu1NtDoOcJk2yI6cj3tGNv//A1PUYhT4Rn7dXfYmZwUSR7dTJXJcwWk0uFtXqe
AYuTIQvP3yGtYrAUBXwHHr32LSpBGRyuK03rtILMit3+Dq5cRO8oy1vrB6p6TNLD
7/PEQ5ja4yJXkmWrkMl31ddl7i8Nv9+Zd9ol9g58iLcHBTdnxAgijN85IfdveH2A
8dh5YTYPNkw4ZW1DJfah+PmXwdRV8ckuQTLsOTDW6dEzIc21YZSSGvRNyFDT4G+6
66rpLdsAJVaAVvG0VzrdutciOF+WTp1aTcjDUT2ntA5FxFu+oCwNhuTDwSX/AtDx
n9FLMufTysrlemGdLsIG+ZmlXXX4ALTcacECGAMJn0BHvR8fA0tsUaq1/Df6v9ED
Kmyyg9ZOHzhSH+te7IeGdgQSM6avM5VEkDfHqOG7iPRKtJjGoF6ivwuQy9kOJNfE
tn5k3EqYZIo++CsZ6f6/DcEd3OYn+bwYOyJhCSO/ooIebxqZCd3onTR6AGkN4SYz
oSARAX5qld8sOPG0+DzEI1oJ/4P7HvBBpbKzi0ngN3kYiKGiKZbwBdCGO0qNepD0
pvoAKvq3HFBrL4kYvrpfQ5h8f+SmY8pqWsFBidDx+I6WAdkNkWrp7CWz+SnlZ03Y
Z10mW+wrUw4KX3IlNg0VRrsklQNIMU5PykAeYSlF5x/KH3K/MnKgLAcP0wa2Rb5q
/t/To4no8H9ZUE6eZmxjaMh6ZnjOn2PD916lpfM16x40/Iatguuz6n5ZEUJ1kJQs
Rc6Nk/wtp0XdPM2HHKyT1P7Szscq7SP3nQSdm1aGy7ySmPovR00Qd+9GaRyWc1PS
dKoWI201dpZaq8RYVgGmhbBUTHjRJThTFTengTi3g1qt6mEY99SfqkLmeyGSFdoX
KDUJbHPHuDtCuOwnwn7Gs19I/IKG8EUVZbkEsICtWMLaB4m6xgcTaMOCs+K+V3ak
0ZsCqwVtdCHXvJR1feFqJfPp5u8khom7qMTTCr7gGKGiBloqI8VSq0Cr4I/RDrX8
jhx/pgKLuf40Jnse77Y5Jbx/dXwNX36Go8c9TtkSJpuZnDoP9GH2eqq635wyrOpl
Qbeb/uB5hDVFIAwDw3tTqUKE6eFjVh0RTUQfrA/UJc2jNGUuAiXq6t4GA+pUvlNd
pbgYvIa71cQs8libo9Dek7sYbZkrdEzenjhHjHgANNB/EStalPXzJrtAy5AOmcmn
BnthpZ+8EVx9o6retaOybkiCDiR0sH241uf37C4gzvPEBJEGbjfDEEEBOsw9HuyI
NbDAtfb495OS1lj/z9Nm3K54wqCtGecY708SyfFBvic1s3U2T+fvGCBzNOKJ62YC
B51DNW7VCsWNJ8jWnaKJypEEftKatfiMbLUQ9hKQEwK152dw7E/yKTVh7TzRDQVm
kWELFEjmLiGLKnPIHL7k3HKX6b1ut51tbc4EHNQ9lVptTAZMkvyM+7DQbi4BAzbW
UjXAlvnqifm9UhehAC/I5S1S1EwTJgpFLkK+c0kow+QEN3JpR8PJ9oC/W2wqSCPp
sdY6RXcwPdGYvKKp3flv3mjSt8DfjC7A1QwZMz0dejBSoyim15w5WOVJwYjNVKfC
8QzudPFUHi3F40FV/mtaLPK2g+1NVnCenCypp1ow9KpRYers4ElgP/W+LJiMCfJm
C7oeME0cstcEDD8gD4dpRVsb0zkfzD00o6k2C/QfGoGwRB0BBAU2/c/SsUS1FKB2
Pdvw/QHC1sN58N2lPkRE4q2hH5wrInEiwsZMzcATScsk97CqXz4PCnCrrgmTgNfs
uqrYmixiS1Y/D8cf0UC1DRqhlmIC+rWy7aJID5cBnjasQl/WxigoiPj9duPiyv2S
aEEiUCG3RnkhO+pkEOcwR6cwbJrLkQ7jvvAgHl9XxvA1AfYqjkQUFU/kYSwRruZA
9BRVC24/84B5s6eixd7qGnG8AmJ18hL5QT644WWh3AU0z2SkERyV2BSd4FNGeNIS
IvNSWZL29QIeJfA59g+QaMpvSDLr+wwaVVFyjX3wRolPwXKv94gfHeQHxwPT04se
1bnKVWG/qioLG4ogcjv/YSDGP/MJbNw4J7uVDtjhEADmR/EZOTSXuwNkIsT1BIwn
QfycZ9HH9MG0osA5k3yPAlJkrxz3MV7Md2XbRFplXRDqpw2zmZNcFZTPNORsPVQQ
aXbaZ+HvSF1uNbfXoEJbJRB+Tt85vYrN5r4bD/EFd2gVYxvcxt2fOoxEtr7oMAxb
IbIzI1nB3eDJaRohCGCZvQU7cJbNr24Vgd7KRSP9i02upLHXla8/39jHZUwDPOxr
ZKFTrYH4c/qzxruUNIIeO87TVrXe7SqLKkJ2Xqkxpyj3sQMOYCeiOLPJM/FxCKez
gxzstfWWY23cXe1uOeGz+RbJlSuE+kiDxs0RJd09ZDNmY4AxxDvyTi4MJDxfBQZT
/YN0uYwbsv9k+359C+aos2EBjqg44b7LTEIQRI2AXoQIIsft68umyVOdVeOr/991
nvkHkDui1xp+L6mgXWAnXI8icHHHjYp7lmUNCvKHKrLFfCvsZBHVruIs2cIMI0YO
g+ZOqswP9BjDff/8F4FRCx7h/L0EWySrOGt8SUzpWWNkHrW9UBR4RKQR/zUeXSwB
OI4tRAOw+1JlROkh5bZq+J0SVfonHTWN+oR6DPl75lgkJifDHDz8pXDp6GmjQmRr
EHqxeRcD1wDQtZsXcot19x3RNBiuRBiZYF8m4rRrBOQcUfKwvax+u5ZRHT+664Qi
6RRRi/4VQrPyXQ6DohnWgLO5krP970XRob6AnKv6rJLUgcTj/62gYSaM6eOBE06p
m1fCdxGaZrxJMIF4A8Kro3Kd2WP0hmxAHoiKx2PORVfKp4cHgkfOwOTf8tktq1Pl
QPyhh24dgc9qaIVbvo7W3wjJMjlU+tFnHvsTLgrW6Qc1r7qdrHTFxuLPseDYGcCZ
tsHeAV9cQ8M+S8Sy5cbGPKn5/qcAAHxtwDWUaA+xQY60eZxpWsgwSokIsmFqVMpb
N1OC4qdypZLOizOqFcN14KM2h4frGuIX73pfbPhkLpP0vwNntmbnmmUyMW7DuCuj
aMQDnEa5EZiLWobUklBlDG7yMYeKtLkQi1Up4b6A9QqpEpjW1l0+qIgAc+5EQyC5
Zb5CragDuB8cO07P2JmEQoDb+q+WHlMXYz3TYpbF1iX6WzVw93vuPJDpvkEFVwSN
BtSRTy7qcK7YNDRNAMG1m5KSErAwATTvdV6JVO7Me275HKwck9N35Poe98dZ7/xZ
gv+9w0SLMGMnn/P8RmrUiYtz2liOZoh18rhJ7dTLBaQxA3ziyQ8O9PuzqU4VNEqU
4WS+zVJFnC76flzQB4Q+sxEDIAd4rkwt1gxxxj4VV1L9Lb3kxzj2+RfYv3+jG54n
qm8Ce2q/EOqpxZXvMWp1t00HLXpSPLvOe9neRc9F4Xa50mLRNUhk43p1CXFX3dcT
dsX7Skyz2mjue9WAfqDaFyzdmLqbKrYHp8MNwtfeusWWUM7oNMp0e7e1mMVKYC2t
lrxkh1q/GBssbUAV88jn7tXz3A5FtFwnzt5PXVmn8gaRfmJg7l51oIgh0FpiDMiq
Z0gQHaoVqaccgciC4xRs/BrMCcJwkXN/sz56z+sX/OAhiynRzHZWaA6/QnVXMf76
6klveCCN+OBeJaTXY9vaj6FGkAJvb3g+B+9o/XQlrBZ+xo1FzxKDytw0u6498eZy
2qWpV8jFPFebxUSJ8WQJbPCBPd70lUknovSbEpiymyKAW7QsPM3hTaDUBeL+5Ru5
g1ahclfbLBhgkqr+A49ht9RtWE8dHQKzJ7BYkSD6FESoCq8hjF+axFwd9+WeWPm/
R7p/ZvEfgO3s+BMRvc/UmiGKtuCXwrDJfmSiQ64LReBEwRffofboSSH6k+RryNv1
y9J7HGtdfP0+3s6QFLCvzMnXW2UfY+QHsVLYVQ0c2OAUW1esdFvlX0X8GFjX8m4b
v5Yszgbn8J5MA1IHJFbNCY1QvxR/Q4S5RnCUvcJbqrPrCdN7V7SiIhTtDZCjzBb/
PrjNohF2e+kGP5su3TAZ4p2qZPR0zeVi3apdF97qtYNiKlVJtT/3ujY47ofoj7ro
oNQ6yV7iuKEkoeVv+U8jAE40D2L6t8SLjDs48+QJlzd1y7CHtbJmkolbaNhB8Tgm
bb42nac3EwPpqn1KG6wrW3P/znzFYpo5f67/xTQ/PZkzjBXsqmpG9xai25QBSldE
M6Htjvtj/MNu4qk6Zkn3H02GubbytLCej8EZhbJVEGeCDq/kolaXJnFc2PPGwSmT
l0AEud22UUAB0JXdgFzAYc1Ow6ykwUUJSXp7D9l24gQin7iw60le+L1oVwC3su0e
1oG9UNOJvqp1YVvs80xG0VusUIrhRBqA1rmpaBWQWjpukE5ifYKGXYHpbtS5idXc
adJ4SP4ihf7JpraMHpfj4OmPTLYF6HJROFy/1DWDgeULsTtUzgz+3RqszSx/EtjV
8ojcwvLR32nU18Xavx7gTiK/1L3xb63kXAhLn5PoWSDpGbYQprr+PrkRWcxVY9f3
41HRGllXbuWRmywnkp+nxLYlJ4KxE7kw0PAv0kJqJ7Lygdvok9970YV5EkDFHego
XoBJrHl6n/1qjSPFob3YE2diw1uobRfXMmOuFfMv4z5rJMh+nClU/gl9pLOt6BGM
L1wqchJ34uAgCiJnMWeOWFeuMxsh32gJWLkEh0hqvNuf03oZNBWKEejc5xZJkxrc
jqWAMeIElSoHEqvuCgxXPKcgvSAxCVLDkPuuO1Xenl+6hnqXG+vP9RZ4HGli1xZu
efx0qRl/MsHaLfgrKb5gBaYTQRjq2hzfoHWf5uuAaCyXJ2/Cxz0EwP6D3XJ8qO3D
mmy3uW3CYXYyBPvqpaGPGwZ8b/9eslNu9cJwsbdKIIY3KgM6OcRDMPs7Xc3lmW7H
52BF/ooXWqriknZgFYfXN4geIbqSKVD/QkUly8m6UVs1a1U5w1s7QG/ZsWSbAE8q
wvtcpFNWo71tGHV4Dwokwwl8wBe0MsJZjng7zyXI8BE61j0ovlU8FyrmJl1ZIO3O
LMfqoIfedTa9grhbblMbz+aKxk2ci6Cgi3u66WRR8NQELVUM5g8OtAQCTn+WOLKa
G1nL9/zV+TXxvlIDHzMpvDuQ6i8MDm+1MSd18fHN4q/XKtnFHfc6TtEFefPTxJAP
1OukKLvtq8yBddyD/jyezGI2+liR9+CrXTCDWuSZNDlBDpeqKmnubiZDyCafHB1y
Ya+U66XKRuFJ8xwaxTZEaKmOzrB5iA37bOGOstufSUXClhW72G2oPTlkOYKHuCT3
kziuTk11I37wnWh+q80u0kZux5H0qZYYnvnzpYQ0JFs4OC1AbP6rwxe8k4NBA9FY
VAWOpH1FUNugUC64q+CKDRRZXAeY86uem9szxsPRIBrW5K/YtslBWFu0n2QM5NjH
6+VL+25Ri7yFlGM5o25Qrcv8cw0yuas19E1TnTa7liz534V3oiLqAUghMRSgFphZ
qYyTHSl+kLfMLtvE9DAkZfdOtKD270ZO61hRXMsjrgOIBAXa8zIMHMG6m2JkDy6D
yJ2+QcRHYA79WYQf6LLspInF/j8wxVsU/wyQYviUymWGR8Puu7IsZbbECS2c5FPt
7KjKcDvIy/lF6iQuZOgcFcciG/CbsW2XBWF9XLXk3KEj+PAYBPxitcmHPeuqgJau
JCSqjDbJlNJINVzvGQ8SmPjhQPiBwxggL4PDWubdUvXjRpI1ZFWJQL9Zg7YzT57H
pLwfecamOH1MQdJ2sWaNzPTBCxJlaj8OHg4Z01wNs5fLDpLbU7HSeKCVYORNoaWk
O3yQpLb2CmOCmPuT9hOPbmrBXpXK62astWTkUW6w4Cw0hyU5wgFyyFv0T62+oeE4
DR9RPZLMVo88wdTKgznaeAjtGSsRE7eJC6Sn0OjlqCNqMyaepbrJIpvZ90cCq39+
X/qWQqRNMN5c1JY9PsyGrbpOY3pa01/DZfKpy94DMmh0NYmCIgQbD0McXPlgnGsc
ZFr21tLjaGuAD/r2eK07lFshG7ZojcFKqmBrDn4RQin3xz3a64q9UQctrpxd1m8m
iGW4qFwj0nnGo3lze5qzrVcobvrVDg7FjzCSwoXjyQ69u8GFb+jApXHiWYQZr7e3
o1BpOQGxfwMHEHYQveZ5GU2lSM3BZCzsf3fAFgIKLMCjplQqr7JGcta/1GAmkRlP
nJ3NFAL/3ts5QWNXai519cHGrBmoYm7DIezuwXc0nDEO/ZZcCNL3l6z12KK4ft/d
/BjAkM25kF/+PNp+KPiWHRw7nM36uhK26yHMj/VXuqF7gYWQLVykvuTzvPNNzXI/
z5JCBJ0kbvuh01+x2cUrQz41ibxNPLViAYjBfWx+0GuM1QRXwkX046BySJ5q3d5e
w4+2oZ4mYFkaDVfNQBkcvvYnOPUrdPuFY7Aju5rJnPqUjqv9A0ZA1jaI66K5uC4c
pIWo0pVPbdGmRbuqmmsCj6S/fGwZCQChvUKKGdiU5PCs9/U9z4UHKDpV0MI5+Gjw
RgO/edtfy7lG1e4VwybG0P3gqdzM4nL+ls/QRX9g31zV+Nc9JR05U6FopVD4sIft
FQM6zM3aJnI1zvRSapta+NNdYZifAwWeFmPjp+Gg1gkisSMiDB07O03zkluX/glC
nhW6a5OyM3wN1rArpIBBsQs0suPN/lLXxCKt9l2jzZozyym4Yp2eBRSA07OFK7b2
P9YH9auIf0DyxvJmB68JA/dsQxXKJg2ws924mZ2E65/Z/qN6iyW/tuNElxTzxAkE
dGZcsjDNCS2ycP3C8IWM3D+QRv7MjIj4HKs/pWRIdGTb+mrkGDId9FezO1+8tpi6
8MzDCDpNMKPY3Wk39F4+A60qR6mxkHzdECzwcpHUSTkfzaQ+4l0Y107IWgguMwvc
9qI+tHmAwvjtzBuhX9cVddKpWn0ZeM788cFc7STWr+QfjEeQEMP1utDMheYYgMqQ
t4J6SUAxSHA5FjYGTTwgJ1RWs38pypZE67GpprFU+3AVopwzsDlPCQbzEHTS7l9B
DG10up0xzoRmbKSSmCYVkAVr72Hr7stTkOab4bWjIERbSC2RownwmaRYE6L9ez1j
rAxxUwlDMYe4g1zA14tLgxm1codlSzpil0eMnInLonZuYDNjRb03ASenACNPtYNH
dyjWR7QO9U8hmbf8c7LsS8k+I61T8DQ1koxvKrO95r6To3Nvp+3nbgX5skPrq08D
UyiQ1RHHI46QUtzC0v7je5v/i+BnQ1lOBxMLhg8n7dQK3H7krHMvE4b7MKSO7JCu
kBdtezrIPyJ4k1CiVYwSvJTknpdZmjhW3uV5QjiWnA+DCIXHt6C5FHJo+JapxkgV
TKopWcSEmXA+y19YNMFoPKEgBASFdbfYippoGUOsd2daD8NI6/tKNFizeb9WuXb3
Mzn/wr1xjdsFYkV3uMa9E6vIuGVl53cAA4vkBfe1PhJv73YBV1tkpM97QBEBg+Ii
Rm7yaM6r9CbytMaClMO33vekmANxISi3XFl3bhruQ4Z6x71EpA9Wp8fpSht2WHbP
qLkcXfQYSFDJXqkV3OpNinAC7lze40mzBObddLzqd6XNqZVsjX2NTgdsHIEo/Sc8
nydqX5BOZiLsjyLbrVXpXiA+LbJq/Rks7snlYiLeDKRdmzf3Top7KZvoMQ5nE13R
wBn76oYX3E6NhSUhkjG1iT8bNx8USkGgJkopmlaBiC5VFDf7JuydHeaju/bpZKJO
+0MiVKeGyqllZBFtCnaUiAy2X2eV+4e2fLT2EbOZCurhpT6hKlimBl9d3/P5/RJY
wiM0BNnGNrLBoJPH48eGhmTxKRrWGl6xIoc/xXMmj+Tu5Lv6fVJToNIR0iB0Jlsr
Pw2JryB39IXhSgiJqk1aO1DY7Fc5hGPRtnYNVugF3C0T4eM9Vr0NYopEKo/vKgV6
cuSWZo8pYxS9ZjkWY0zxNVbZd5l9o4wsvye6x0GKbVfeq2dqerYiZ5FiGmnBiME8
3ya1V4vmyPf6Sle1397nxgDf5LMxxmuq6lOof7xKirKrFLVWUMPnepgAkUkWIZa2
KjvmjUOj4HGnwFG1C7wro+17jfWs9VjwOHujP1ondiNizG6Pfu+ZmOATxCyB4abW
CAZjvOn/prkUEHV3N2sHO+wAMKYFhovhYGuuex9TM206HnIhKUD+yAQ+l2Kup/Mj
v2vPKX8kIKjQ6fCaT4F6fl2zEXavF5TECO6rFkUDuAj/tiSevbawDdA71rUIIvL7
ubYtAfxDpkYCR1NQcUYuRvWY6bi0Ry1YR5++qDQwLjf17pHLx3GSAUgu51wiJUKN
J8++zJkGtRHCn6rOL1pRtpXCJAwfDAyeuYkhtdi7b8+LsQVjXkvK0tlgDbhggfY0
IHcWrFhany8EB5bPgNhf3RuurhIxEctfLSwTz/aj4Q1eA2tCNYuhmJIPis4vVLXd
XykIW2ne3v2Y81CERpIytdlDq51QAlXiqyhNFlDW6QOxVQh6lgWwhEZx7GumRm4o
vy3b29OFaoAwdx7iiz5d2YfoUBK+scgpAsxrXR5LzL0HeLj8kuQXveXNEzbMkbkY
RzGty7CiPXB7xNSPg91agxjuLvfNzwydokuRnK83lRN0Kfc/CaY6NDMbSOx3yaOY
e/8JiEXA+7+OITAiRZjd0QRIi71wVk+BbngNYn+gOmYPFahepuuVMP6ilSTDbVUD
xQBm+aLygnDxFAo4l+LXyZgIp2Npmm1jy/XgoGTUcUptt+tWYNlMJ9Zdf2mwjsPF
e/oX/J4knVgd5GdTV+89pUd+hz5KgtUxSCAPgb5zEjARXaxvWWMJUSNIKt3x0jxp
STwFxGJOuriyOARcuKO2gx0+7ZvFVu53Ier2eVb4o7PxWw41ZRSs2Kty2aEtIl0o
6B/D6UNfi8Bcik/MyjlX6eBAxJuC3r/+G6o4F5OWE05+5TtRLy/QRZ5GhahS1bSg
Qw5k/v4CYImzpAd7CrRmhDuDK+PXKbNTKLiI5MMrIlIIUGKklIXeQTaVzPi1A7i6
lWWPd+d2EXe8ylnEDC1NBP36H6u27FOpcZYiY9aqJAr+fhQO2a8ieY7bh6OBaWd8
OvGQ+ODeyRr9OpKMTAshoGRrRhPmZ2pFztLp3ffJ/cQ9BJgcmdjrHDnsfzVgyfCv
oMPxXy/sqwHvk7WKsf3PX+KLG3Sds6BB1N8ZiAKpBGG6AhRcvDDYVAnHIe2xCTPt
3g1G7q0qJaXH3pTWHfMiiDjsiFGE4s1NjXhz1L2zNeBWOJoh995e1yj2VtzqXSFy
0SMjm07BUa1YZ+o8UuUBO6bWQfXngJDRb67p5GzNuJmX7vFOCvNQYqJ6EJ92rm4I
PSN3Gh4fIrlOoJ++S6Kef8USw/eGonobHFyGWkzo7FEhIDx5nnuzKWranMqz2MYE
rKKTdEhsbvNApv8iEo3e8M9xlsxXBfTrr7jQFsmKjrDVJbZpWm1iAMj03Sk6gF0z
clOd3H19NuYbBG3zKZRWaVGo+1g7urypBKhIoLJ9iLxRERd5X6xLIQbeV32QQwMt
IG5ms6qhVzi0R9LFT+e/aEhwKYh08lvBo1+bEpMx5q9R32+1t9HFZTrzDrBBlEWK
l0mEIo0zhuhAScfCfZIwcLu5oKkqcSDG1MhzLyba8URvfISkXWsgjArNnf0UGE3p
T55vIrSjCKnGIFpi/bYw39uTjdYo/bGSTiRxhcy97ucU06YmcmV3xWy6DytCptoS
yrhN7QAqST/NdhQXxRZuNF0LfsWOXPupK9ed8b2G+YC/Y2bVWFmL9hX1RvaIl9wG
ERwSqR8Kd/EtUH9mJmZSXBdI6PCBTfB+mOtm8Qj8AJurjEMKiVPavRFn3zv/jkPs
yYsXfN2O9Ve/iIpc7/TCIr1L+uixoA9ZZMSSqaL+DGcTu4enSB+NWQ8LotF+m5sJ
TfO8VOoWUAANnaB8WMbjiKvyKbIgxyXEc1KY2Sam14Q3Kjr4iV2dgYVusmeCkN02
V7DXwKekYjfzBvlFqawhUFt5odrhQCmSmc2q6SYC4JjbAMDONNXf9QRZnrOe6OPC
Q6JDcyWrAL/UiEJJoSLXoGUgj1uAPF0GQOz7yx9FLb/ZwiTCMD656Cyl4eRQ9EK/
FCvl4NRKBOQ3pg+hkwJuhqCA4kxoWzMuFcnhzQ3RMenGmR0G9XEZLH6GvA/EllLR
BZW8goHa359FzBsOCFY0KpSfxCOIquDxlws4hkwQ+PdX0EHs3wvPfsEXKGpoDBmq
M8tbbfDcwzhn6zXAPVrT7eByvCNkBzYsCuhJroA9Rlw7HZ939vv03t2Dk3zG6IIp
odVUhhrzgZRcT9uf9uUMiPtY5kYAEC47YPtT5krc1u7OOMwgPxII8TkhtBpPb6Lq
pxm80RmEgM/RqByaeD4hO7G1hETc78cUSCNq5PcwUugThOYTYgS1LYHqYLsB+EZF
vyMmMWmOmQYAPMUJFQBCg0fFa/dCA+RymI7FgdJj4mwniJlrIsTjstysDyJCkkyr
sL0squghTkRaErEIzDcAD9txt0zjkdlcQwDE1LuXhHdJAdgdLem70TBZ11cj9i6S
sXhWO9EkVN9IQF4g5tZwG/gnqD7DQNTO2XeetEfwN7qdVy+XxC86aU+EFclqXdYV
iEAMlzudPvbp/H3OSHM0ZhAws/skpeypApTzg4msxlCGD6xjoqG3V5BVq05niT28
U8nb9f50vJL91cyP2dAlEIQg89ejXrSTKjb+qkSaVx+eZnBtS8+bgOWi01COCjqR
5QXPKDVTLxOsiMDYm+wWmGAZmCIAvbkNGF+D11WyR6PPE5wjhRiXQu+lXCDfPkNG
7tjWYqM1bSEJ72jZOkLY667DlLbmv6ecT6PIhXK9Wa6XnnCnM1e7K6RifdyaAZq3
SI7u9P2qaKmnPkr8GW1Wn6WwX7Ykdr72BvGGZpzm9czjnvmJ0zA5UE0OEb5TTqbP
lZFVagBMU/S6DTqbOc7UD8/Mc2X3VPJzVcDusoL80IocHFOMeymzT15Bv+8dHVJm
qkO9DhwtgENUX2muo5zYQKwK8TUPOnkkvOqHQWU6gH9bHqrZZbxXheOGOvBFkdbl
KwKyqawEd5/79im9HWw5E6D5N3iLoXMNFr8N0cihUDzR6OaXWyLxkVtyBkWuHDpr
3vnHovraEG2C3VEevmBN8oow01v3cLgzlwMUBpE6ev0MKN5Ip0dTJ5I2P36VoTPK
2vqX50HT36dnAZupzVmqfvt3WvrVyQaYDacVvAf1vKzfvzgRUws59RITVpAL7WF0
e6zbO1BMyOmc7fqe9B9AAg4rz2bm9s45aEabM0l+8M/hlla/IVWYAHmAfPK9DLkl
VyEF4iAIfZFhRkfAX0iWbGp5WTY1o2l41QjAsFA1c/1R3MQ6EkgPIZySUYtV/aZj
c3v0yCRZwR0AIJgJcSHrPIHyQ6EXffpNTwzd0ptrE4jQq+qb/DWwbmhqaiuuX0TJ
dL5rgH8+FXBOt5bYcBN2amVOWer4UPjjNnFwJt6dOhRz84yUaPt0jblEwx6DK07a
cGSQmH4S1rwFgTN4UYDhFEe12KMPj45l22L50qxYChwF74UUI3EVSWKAUhkPE4zd
SUHBd51LaIFv5+1qeXd6GI/P+AN54M0mdRVNf0yA/QHAudTI75CfamwK23enmpa3
nUdFKAELPiy03twUptf1A6MpHbWE1DRi9NaKLXdlZanqU0T8ArXO1d9UO+sB9HCt
I7u82276vHYws7eiduJ3XEYyrY33zt5xzBUKrftaaEWxjK3rKetEloxNKQuOgpRy
whmul9UpE37FV9MNvoh1MwIZeRW1f717FRF61ILqOVhwGOng1wNUyQwy3k6rdy55
aTOry5q93FaFYMtofM7oZYNGPBzDemNzLsUq0ljYK+IL872e0M2NfCJ4Rmz9Tf9G
YNXD57m5QTL7i6Io6lLZ6UK28Kn/KqPnWWvDZsQwq9Ub0TmjLVpo70SM1oz+A4Zo
IUJtZz08L1zJkCuRhMwoZSawOsa8QvJoTMeluONj8LSeiGH7WGawgJ/fd+9F3uUw
lXxyJP5bP20lyf2NLTea1ZQQ+2M8qB/d11PPmHMo1M2/mreMQXQvghU7xgLAw6ob
TrRW3lz3erfZf0sx+wXgmaobdN6MPAn3JLCW2c3gtI31GD9lLSVW6gTQuIf1A45B
O+1mkjjns1YsSXTyI+lQ8X4b8/gbQbTBVBbrYufV0GH6Pq7OnpK5geIbbEphxWPP
+rZbp7mHCxNxiRUkeG1j/0Eq0w2LBt5H3btu7oOvAjE0Y+mrvHrWMF9Y9nPShnRu
Ekh+5f5vLAyOk11bXIrCUfNX1wQaTWLwM0vGMN/tJjsnAkcP95MNDwRdmwRI/v7L
qjmU6VyIe+nwYlow+iX8xlAvypBHIKnjv54vHJ+2zD/c+/qg4SJ1E7fcW2OUb8+O
KHhxlSfI9ggsp6SUa/Z9dfOsMO4/v4Fet3QptIDI2ig6sCJu4z8/Me1TQNqkFsBj
36VUQo8ZGe86BX526YxiZaXE5zw/7+fYnJYO2h5mIYvR4JcAujflsjmbz4+xYv2H
SkTXTZF8KVKszaKyDk6G/vy8kBctPhC64nEZBO+kiKiYu+WUD8bFaEVfdxPKI/Ji
HEIBjwQEkMk8HVQzZp/hMvOL/eEl+2AlE4C2ym7DMd8YdFpGJMI/kZAiBSAhX4cr
g9Jadhtpq6HkXQR49mDcw+VZTTZZ2LN5qULqu11LUEmvjOWSdIZAw6FYauvzNNp/
umgLxDUMR9oJI9OfgpLDA6r3y/2rjyLo0U9ndy04ZvqQYD29opmIjMi0x3p09TLo
8U4Lvi355jkb0w4IoXm6nUyf4RUClpxg2WngwspH7eKxol8T4/NTaxcWxLbhv/GA
X/RXZLgqZ0lgXXqtk5IgpFNxEFANcynOPMwV/ycXZ5H4XhyFYDcmpbLdaLnfOUy8
symcdWdXFlUseIIS7WRWZVofVSs7oKeeV3Jtr0if3jB5l3tS37JhoFVxTxM8Owoc
N4ZyrowrqNp3vx8CerHDkpuSppVbRzXC2ka/kPqWrX2GB1xktPlvZbhgE/FlLSsu
KNHCT/rtXnt5l4si7jqrQC38rxNM1e6MGBy2+U0Br9QikXmgygQHjc1okuzPXDkq
hp7NGKJxiWn/kWnbuPe2tSaqM9GninY5aYbaMPxGSxp2TytWbn4jQZrBWBT/vpXw
HFu2vsTT1mBLvlcL6yeLsYvNI1XBbfF3omnU4cFSk2m6Cukpw90OU5d++ycDlVqE
k3X8pOodxcnmH3XyrtN6L/hLSNl3n3th5yOhBcy4zw/1k4Nq3pfXcc7QxJW0eazm
ytFjMl1yUaKE8O8+PWLU7FgHhaoa5OvLn6jOiD6a7q8v+mZL7cTPq7w5aRAROZoT
5S8zxt/ruz8pHK8NluZf3bHYhI3inSIOt69LNXu/LZ353FVnT2mVzUBahzdbsPmG
CIqTl8okWDsQWK+yHcDnss/o3pvS36+aGqhZqwNqIsRtZvy8ofulM6J2f2aZdpaX
mzc1SUFbj3NV/GXaJ77KHh1HPOkR+K/vwRaoalsl+G4zplNYoJTUNnwkWp45od6V
PNpEDcO/WL87rAw7CnjcaOZ6FG6dKHMAvxAk379Ff3sBrs6xUMasmh55nhFQoA1b
leL0zTq1/OLIg9TQL8nNSfJv6XSqfRddQLmXZRAV9f4ib9twSHEE8B8J4jLPrWmx
Mwt1RokCoS1vHt3RPiGQbqtd4GB5yWVS49vlrGRncgmf9wnSbJd7GzED82Du1fGx
sl6sl8w1Rdw+/9UHzm4m2qtSTdrgrYRjmiRhxMKXqgpcTDkDvH1XoML5nHfOruaO
Ekcf6Zhzur1kARqjul53ZT4ebeLzgnmonFToJIIRw7UC8USJ90oLvGWLyhiYabE8
gQU8u6HeraYT2V+NXKrfGjjyN8BuZUeJpDdqxh0mR3hgS6YCQT1fTjsA3TI2uxP2
Cer2SqrmCUm9LXUDmPGITUpaOSLPGl5q44FF7XMnLG0eBrrT0FJYYf3UksnXXAkq
uaQDp15wLtMtaG476tHGRMnjN2mHza1JyxkIv4lZF6XPgMOupRAJ1ByCJzPfNf+Y
Vet1hay/ahj3QcaYtgjAsH3EuUGfM/JFXxY7g7OEY79YuRpcvcQnEWc1B3S06tzK
tvSJJMOp1FO0FqQE/mE94ypEv78jMf4wTnjSIQ2uybWbaDNzYycMaV/QTjrSJzvH
OmVwPr4klM311VS7Z9gytz212gyiKywrQOmM4R+nxweshOh9fAdDlk61z3MY/TjV
5PbtyMi/zxMtyhbRvFdjiEOG/h/4tOWZv7y9PohXM2gdB6RcD4BVsdDgYOSQAYs/
TyYzxTKG+WkfMmrP2GEtUhfXdtVM52xDy8Q02C1mt2BAj3vi2mrpuMnd0rlmbQ7p
ZYC5TnX0XMhE+DeasRlbqaQzNsQ4UntrdgtU+QpMuMWkKP1fc71uQ2veoIoJ4B6o
63t278mZOHlDB7Cco1FzDEM6sIJZL+XgC29hod01fY3AFY0Wjvl7f2gIcbNgwLtx
jNT+ATTtcwrlo/HlhhtbEagNPi6EodcDwISbCL8jkqQeWSXXRVUoKEpl/Z9Ck+x5
aceViMF7JXi5UT3b8CrPGmdBKXFDZEkcle03AGLifTjIXoxWScMUtxB7v8TqWKaG
CLtRIRcAVg1UYhNAcE+THDIye1yeE0zsl+26MIZQ/P86CfC0mMXqJ/SXohv4igUA
B+W4463UQxV3FfOMOU3AWKudpPUIbDtR7R7crUUVpezNWJ7CivZDjEG+aw7Ovr5a
JOdPN63/kc1KtihHcN2XTSFEC9rPyghX4o0DYK9BBM6R+/9fmXWnnR12ZOhWms43
iNbzq6lC3JIE26LnKfqMeIygXzKof/BiBssx8NhNmAVbqCmEpuRHv0ZTVs+DNfdr
EHAjxKNfECkXYKdxvPicIZD34XRBIBhQjJIxNZPYhNPC6UsUTbpZ/HJ6c9qiwZHV
w3+hB/MNU63u+nwgnyOZ3rtqc+1KU2z0GPTn7my71yKi7hq8/DAu4QFln2Ns2F2u
rrOw6qeZKagV3MGVULKJd5paMOHQi7IXpYVuVLMDGJNSxEmeQYyUfVqKqcGN2QFg
8W1Pf0XWIM6OicMdoK30nbuBvABc6uXnxjiBSzAiesD+0nGjOfRq1oLgd4mh3iHY
4QwCS2pSaT5+0IoWqn51xp5+PxcGGH4I+wEvjfnCHOmE/C2s4m1o8AFucnVv+pSm
FrmHIheCYuBfXE1/nTvtMKNkVCcQmO02yCLHOA0wjoLx+UV88k2G++6vjH4eEurX
mSV25C9m2ze1ez8eqR89Q/zaDzPR9ilIn/95FsQNgUSr3qi9f3IwPfBytM82Tknx
Frzgp3/lw0p1C1aECLbWNKt+sUEViC7Yr0c01v6EZIFhhD6Amwz4HRxWenucvkw2
lvLDImcEky0PbWzhuX5VOHExBvEYesSlpryWK6vwILWTGb9xeQd/Kb4YUSskQPLX
h2a1i3e6I4dToxiaEfmrF1gZqAqo3XhCowdJicCP8QpI5o0bNtT6+jWhxUmZPLvL
GwKex7YvIn06H92EeaCSIw/Vgq+8lLMilRu3Se/fo+4LUThggGJo6JmXKd8HLpXE
hqJ9O92qlyrDtcW3em1HYnehIHeq2ov5l8mtNy86WJAFfaEfRYtiaxl7nJbQmwsD
BfTBUrK9vCDzrpOme5YyV1WLL+nbU18OL08TDpLCrOstHp/QcNAAAJ7r2CMlfyYV
DAXQuHVJvJ3R3u6VFfTSfkCIIvj3j+M/CMTADoLnlQFDolgGswFps3X4ziqnM7Q9
WdVwyTkohjhoCWm5I9lNT9ktCiEHekDSa+RD0otbjdLAvJqhK00APeMOj3/xnoTU
Hg+R4kU+DOlZiK6Xo0uLehGYisPWcGwoeJuuNR82PhPpWC3ES9Pmsx2jjUE5Qyi8
L36DbOyfWeDXQaNqsgHhsQDDFYjyviMe5czxa6B8jGvPbphc+hQcyeEDvsu9RbEg
qFIDWrEZg4kaLaW28nol95DHl/YV7n88fERayhmnYUmTQzAvlXodw5k1WW2LYa6q
ueIm6LxI5/ugE9V95reBx+ebl/TNpK5wRXSAtbuoChYkZbuXtS1tk9JuCOZtVrvL
7mcEhZWGU9pHpRAQQWAPsE4I8r8RninjKJuvN4KlDYkOJzOVnh81vnDl6MXZdA7/
E6rsmxi3uE8amMMnJ0BVme2kX9I3qJHtaorkY9wj5q9Yd+CW7OnecQrF99I7CKqW
hZq6F4RIDdlc458xVtujs12S8LR//MSZeYQcPeDPuzy4YlUw0ie7qr//Gz62MJ6E
/t6Y+7O0pzloIpQ5+R304I+C08myovOj3yK9y/JvY9oyLpDQJaCtlLlx/du6lLrg
AHfi1QaLrBiQs7aPmgOvb8+VsWOsMKxa2umJA0rkjZYr6lQUkXTk0OoGbT85+kGt
FDozCj6Maw9Ti0gUEXg30NQBR7wOdePjHY0fO5EdJztemUcs+aEzODbDP1asbHCs
R+FCzfA2lDH+/pfknCeI0TWNfH1qdzZQiRyI3tgMX9p05xQwjkBwvZbb6W8gaFv/
45uoEK1BdWZ4pK0saKHdPdSoGa3P6OMV4iv//3oyQ2arXhk3K3BUlO5MFO84BEwi
BlFjxYxP7DMDR2tPecKFny/ivnPC2xtKGHyMuXNIJD/oqkR/RHlkF5foVs7+m05D
01jX4qkeVioeWBsXS9dDaT0RTmiDFFtqePhfP2AEBDhR2rPSUls7ZGokL4C0SVnx
N1sti1Ly46iTdeNtzCughxN4YSIVLFUvkPhZBjr/bzNkgGNZsndG1IM9idoef2tE
1UN3DoU2qLAzdYep0aOfUT/qLSolysnoDpT6gjJXsllN3XwtnvkufoOG97Eblki1
Sgq8eqVbnTshBYTsWdBZ3qqP1AGq0WEgj1z8pwA8RD3D1B8Obmld9u4S+kEg04yt
vO4Tkis+jArD/a7ZeqoutWPHpIuP8+19Ppns5dX0JHhPuccfHZHf+0c+uOl4jZyC
qDtbcVBBNzpJVEHNFM25+Js8NXZKK1VEJpMmC6fk/1//dYeH3kagKLVzPEpbd2jn
JT3bcB+DOKO8o4eTSJTN48o6h/RpFnbNnO0aGLoa4YmKBXddGaR5pRLrQi3ZPZQR
awiVlBmw0ATlmTFw0Qtue2v/TfWrsJyu4x0d1l0rUc2ag8pwhakP3Fnb0IcOg3Jg
Ype6cAEa7JdC8zW8dhn+R0+pkXvK8eZAZgQ/C3MINIjSd54CqgVUYKKXJ4BuYJHu
8JBeUPkF3dHePIo01LapysT9Lvx8XOPg7jvWpsu93ACqBbiz834dR8ZkVKksd40K
XVPXUtdhmRYzwftp9FXVq3ZyeoGylnpCNWm02zd63bUHLV7fvoRD9D3345/D2fwN
iOp6XzPwu/Pahr8Wh/OiL2v10Ellw+sS06OvFkPMFCMujUNVBz+29phHOilP7gPY
BC0977fz9ye6oP5N5uaYazLW89k6NiyYp0yyiKKRR6SYbk+3YXodlfqnFXTA9lXa
UQX40pDo3av7cj2eHLJeb7SlEBou8U6cJYiVpwLtTM+qQ8IjST/vclYj2jtyIW2X
4M1Q6I9Ed3i2CB8ON/C2A0w9Gl4Gor0K/RQTSkViuwC/JnPDZeWHv4kiBr6+Hym9
nGGnI+tt9PjccdFXhmmcEcks8zeoN9PDwte0mdcvQuuWxTYG7etkZn0TvnHDO0Rv
GIyvaI+Tf/j+3iZHYq6KgTDAmUOQSzRvepC3nRug3r5vEMDI7RLp9RVWrL/8OODZ
EWBVlz2cTUC6mr4D9cZYvtB5d77Gr8U8oECoi+cUlmnwdoFEt+/KA4ZzNAf7JF0N
xnnu4meLj88v6HUaj1jGUWfMJfDxbCHMkyjn0pB710Sa+X2kj4xkcvoN0v47671o
kiTMrut0+E+mkgCIuFPm78sYe5+J0ZmkGnl+aX52wJNxKbpN4XsPOLuBlzvjd0p4
qoX+xHllgXKzaUZpbKUfiOOAupAYNjO2esd7qY27GGK8o5Y8jEpLlHI1T3R8/9dF
71LYtHD0zCM/2wdc5oNinmheytmjlMXQpyEtbjA3RhBwech6EBe5u+gg8O7AZbNx
eNrKsUdQTcGU0gsBj8tCfcUVdUKmUTsMWcRJcup6KC8pNT4Q9mnFLtRxXaBR99I1
t1Zhj75QloSqnXJOMakH5SINCJ7prFI/WTkYgKrhisjaRLHCJ2/4DlEqRsK4LaPK
GkNhaqdeR7xy+/sjY/M4bblRA8MhKWgMnJZOTGhzG9aJaoV86bWvSJhARlB6t22D
kMxetnqTatOfLpSbvDbtIwBzTN/VNAXbmTk6c1Ie4xYABSdHop+qU7nX42+TK7DN
ud5MWJdELfDY6o/SavzMPguEu9jp0MM2vZ5c7Ur4VAJa512/BGI1rA9euGZIZw5F
KZ4tBnK7PANmFGunt2QaCPQY9Qnba7EgWj0IwWrLoNBXrxo9dnLjV+Rw+aO0nefN
eG9Bl3B63q/nEtZMhVhf8nxZ8iDlyhYkIrcs3H+jUGstFJSDWc3LHcTpUjut2Kgb
K66snkifr6Ykwv8Q2NyQ8rtanZ2vFgFYNyxWcYZXWX8JbHHNRQkvIoTm8ppDHXBD
sZsFPGrT6wQ2x/0qrRa4YwR4jesUOYuo31Lz1FzA51erWNEvYy1loLE9Svd28Srf
ISxfeIcq8StsrfzXW+Nn+tm4xrKZCphR6nyANHIs2CRy4qVLpU9SHJNDhkhqQ1l+
2oN031Hmy+LKlkDj9EcqC8kHBnVHajzg+2ePSIWtobYQMKcR9+bsFP0G1VVzmskq
bwgTYNdasq5Q4vNEw+ECW2ez+Ro9QILYGzT8s93R76WS9fHTNGZduFmuMoc9e7pY
ETK7SroL9FEFsdqQd3iAnt53BzeXm16QDx1Ll6akmtMOmHklBRI6Ghe3rOYBeHdQ
HARL+yV+HgWkRA80rwWq1XdbxM7E2REWaBymB/IINKboH2Ina71zUEP4VYd+2IXc
eeyn69AQJrNqLl0FgYy3JexMbK8+iSWqnVZ2CAc0XcFw1K9tmiivWi4nSMGXjt0I
ExRBU+utJhyaMDRCP5024FTjx8jovRHHhpii8HJN66sYKnutm4Rss/s6Llvc7yet
uqlVi61ilveZN9M03Kfyht0X+z6CU0Q2vLVBYp8O/dcvOlm4Egedg0ayhOWvfDCl
/kTtUhkpGmc15YmhKwDpEmblFWg/aePW6MywL0tjcVcS8zxp+aNm5ZGMXcxOHf/X
VeDq6pGJqDODtJ6nQ672BjqdRSKagDCMzAsEVKF2Nuc7D5aJzVfVb6FfMdzBBFxU
zTapdNAkjb1dM+4OXwJjZgpg07TSBljyPTstaYNA19bxRd54bEto8qENxBr8qKvN
pGJsfP0opCEAbpK37YCodj3KKX9feoMq64utGepUF0GXiee8HnbqLJTO1PaNEemi
Z2Xc+V320m2HwXhf00/o71DskL7MZ05+B26uZ/qBxXo/JDCOyShyekStLCtEaWiN
ma3TrHoh3+Ff+fbXneilVb3Dxd3St1iih7/D4B55BA6Tyxtb39Z01+2iZWsL0m4F
dNdDYkozGNj5nl/+B2c9aQtva1wKYIlTsvMdjjh5hPqzwubGWBMxThV18RIbZuu6
NBffZOEK9cC6ym8au3yYS1vuYVPwJNSLSuD3yq8euVuYS7HMshD/go9KBoCWpRFp
JYQMSeS52DdRaKibNWRuXvK8CXjemmRjCaX2IKiMXLRU86iszcIHF5UC5xMf/17u
T02MsUJuj45ISuwBIgSQ5425xxANGuOOeP0s571nWmRmrHhnjSSKB9lcUejpVJcN
FxEeDU/8nUIEWhCV4MpSeoh7GXrCPUqo0XHRGouRUclOpiPeVL1+mHRlnfV3NGkA
HRdwWi9OnZeoR6M3iTPa7XgWfWinh5n2O7ZrImslCtpMvj6CR7EMkCFfShZiLUeQ
OVa/YrhYZuow/iEUUOOdHsTKeM1O8YYw3DfiggW5cDEhalwL0KwDBvebDHcQGxFz
fbGP/MeJXIbNzaWlBLcuXv0YOyGDMgoig3ewWID7m4OwxwCy8gC1I31z8SOnXdGq
HwzSxaG+JwYffDQENCrSJngvTbCox1u1D8usyRseVzV/p1/7QnJ6jMLvPtQWE0M1
Sb0eMRZeTBQjhPO1AJdJtCmQxPCn0Dm3aTJwm325ku29veEwDlTqqlZB1s39RX7y
I9piA6hBhI7zJBwTFej2fWs0TQuMEcTlhiHiGN0wI/mVU/843LLkzeoTmfudX6Su
jm0ilxY9TundW9mh+YpYIcc4w02Tk05CsKGB0UEnQZnT5ItF7F9ibpc4Gv+rIzuL
BnQ6yKR0fWWL0c/frCJOd+1XmSjYD+DFZM+wkXes9hnkLBTF8Uz6CsU3WLqNCATW
95KivW8qJYlSf9VUf7G/psse3sZ7QDOobF+NDMXuujND+VpuKtkITvsgvdQ8Q/dF
1eblR2c3kneNMJdxQaaWh9x5RdYetA4w19nmEJ+g49ZzhFjFD1Q0FzDezxhCpZK7
eRcWo56m5Ind2rWCViA6PHdrYpbJl3qIdbPmdyPGYgeeKzyoxGDrjuyKWvEEIDI7
iFvMe0JwsMV4Gar97SqzfKkMKJbk9upEjh1LTWlUUTjnXQrZm9AB6MKS1jMSmQJb
v5q4sz53DqupzDCdqQ4ajo9QPLZPAnLWAphqTL428TPUo3Fwhtxf6XD6btexAp0S
btzZffbHtGHZwGEIrmFJGPeQToIeEXoiX+YEM8xhUeInbKgUJXYAe/rfAkIb444t
Ocsl/cSB+FxA9nA/+2cJ3DIViHc3rOyARKqDomNkBc7Qjkj13xYkARZI7pKEGmA/
UJS+P1epslHWcq0U/AAFegIAHoIuSmU6VaM2d73GMgW1BPmyftrJxs139DXXHRgw
8m0mVs2e2RbmocBHjOY/RyurBzM5b66tnFKM4KipKOUBTKNelZzGdPsO/5VB/X5u
zUjsU+U/08ZiAUilwr9VUPq249XQynKJfeKa8qYAyAvz6OyCx2HOP5cBZp5tRgTK
3oet0LRW/qgEGIe1D2pLlxdkN/0hxUhoFhimebuZ+RDaTTdwTNTrZJtO3nHQ6vkW
dAUrNYPRyN5iveXrnc4jfKgdB6juTkX1b8Xo09sO0aHFiHUP2WBXO9qSLIr2Q73k
aXiLfOEY2ccUNiYSy7P0Js3e9uzuHXKFQqnuU0klOGeaF89B0CptpvNRbPytdcj4
6ikXDsrjGyWtTTY44xSwlbCF+TnZHlEDjkp6cumIjcX7gJnseLZ/0v4MPC+gi/Ds
/jLmr4tnX6LaFCIChtj2vweEBaEbY6z1iiEjY/ECKN9rhejXjtFrZe57Dcdfs0DH
zciPNR672P8yaALu2Us2oFJajWFA3u/esCbZ5p52YhpMxnFThvlWShLEd6epX0Zm
LczD/HHKAFfSKk49kZgqAheqzapfvkBgkBZgitkGFw43hUJVihrC8qKkaR8UMYFQ
jNjzc1DUqFebwwYXp6kMNBYoJE3MVdCeIYWnXpozg3XEnwyY1N/A8SV73cMwhshu
5mGY23Z09aohmOQwQ2NGslZxhbatTVBXbWgflRFmN86N1dyUEkrHc3CqC3Tc2xjN
UklVT4CkbO8QhNojZA1L8vICX9Si2+t2IEtTayLEKdiuB+y187AeG0Rji/+wE2gH
FIk+mDYHEAamYPYuxj4usc27IKkwNnQlx6m2PqleENsNMJ83pnFro9tNsqF3jSdd
ZXZhgrAW/hLtkrEQyDhiEpEDO5AjpQo7R+8sS0GcQDAs9PPi9+ws9rchKK/HShDZ
FxMQvzmIwzgrgV0MR+11311wSgSlADMJKZ3OiX+epqrMtxaMt6aKKDG5wIqnN5Id
glFZNbfVUrzJbUgUsCflptEKxzyadW6XXv4lSAiq8093n4ulIbMKlS76+siwasyi
1Zq9RekH3NdWAzq27I0iB6UYpNKTo3et0LwjHymfB6AgnPlVcDbehrXIlKy90rhn
cggspur33y4maqEahUsiZlmfP5fHrceG8RbFVNoJO9qauFPqm4jn4CoqGvYLOlV8
74wdaNtRghC31cDt3r/GNNqDZR99G/oqKhN7fiV6x/v4mrYc8KcRgnRY2wu3fEhq
nkl8Ufd0mQt+Cn8O57vj5DrocO/55laEZNWAwIRwIRNssC5EsbVlzjFKFLtA7mPI
eKBW+yP+hS0G0JHDsL0rU4rV9u9E2TxzjETdNI/Rs4iqxtRiBcq7pPBACBeZDVRf
rMtl8MILMgQqm0wFPIkMWNLZbwJRVhtGH8VD19snBWKT+4yL6FYnA9/y79ljGcOQ
i2H5Blm19QfHaFh6tButjJ6mcKrX5uAxiR2sHeEFCEojomhBKjNZKDjWxPyZCM5n
+2qpEQdEyUoHiPCXmrtRtSUNCNTNxHpjkdKysUeLNGNGJ3OxtlBlotC+7kfVmTd9
itwGhBwK6NOhmkHsjD6zltt08Xhf0ToYCSAbUS1D4WM04Qy80AwcL9vfiNg0BaVc
THLPKuUK711+Ay7qOj8AKSVKHUvxlMq9apBu0gOj54gKZoHOjSfsCBwU7PfLm4rM
OWHharqNLJw8aLBlcxrNKxeClX2s7JCFuzCJxaiC//Zc0LU57NFEgBLw9qOUXBWX
4YryBNShcRxq9AUwA0PKxZEy+p4rTTE1O6rWuxFAqoT9p70WgTySvosULyUcx7QR
DRShYhe69xxuFn7LzsDKPTjIe4bKqoNed0TS2gVDaKUkgG6Q/sUT3QrQjV695qvx
xPUlrY/EGej5L3kxAv2xBv1E6Mgjig30Xh/4M4vP1kiIiDjTJoRhEGkXxQR7gFy8
aHNs77JxBk5Qo/3OBrSgMlL5QMhT08RlwJuIYm+pzRb3kYd1AXeahAFJ46jTxCc4
bvMf4fEnRZRcOo/5SltW+xq5jJgax+NXqVSPm03y0it8Po3X4c3VjR1Izo3MMfgB
MvnmmWDJthxH/Mj/mO7CtwfPbG19eEouDDZHt5oyC8CS6GNOLmcN8Z5LcimArCNw
jtnH9kn7pZPtpzCXku+L5g51WetpJ+YrlU3LW3SxHJdUr7+r+HADYB57RduXoVfc
182UAkKKEybrbgZrrFxG33NL6aD2/5HZ1HBCaq07FsaTROVenW7+Milpnm4aSeMI
I5YAQl4f8PDetpOyUcdE4fFu+oiKYw8Z1/Y8g+dSJmWP9pT1zDOth0TJRHsBr8z7
OE24ZBWILYglWrZ9vMzrmL3WJBeN0lpjzQnVjx2+awQK1rLLqyW5c1Sw2MnQIvbj
eLRRZx/25L3bh+m5HKp1/HA+JGCmdVMNzYg8HJjrd5fApuvVAH8YZraL2Ou2H8lP
ZQDpEMPDSrg7K+APjtjHly4HR8hUWeCvvWb4sC74rA/fvW4ckiMh6lgcBvw8ergs
46dXuAfr/Vq/abRUNvm2qFDL3TNW7nZrYHOkQN/EwZKTY5h//ROpNGe1itXNI/1a
sM4hL5cUlZtELsp4wfxxQwR2fxCWjmt23kdgs/e4lLdbePMztsH1IjDU7oFtnRYx
gu+cIZm8ZapWmspmItXb8SUpUB+QMyspovyabwhyy5xbUYNQxvWObfJ6BsWJn44F
dF3T6gcqIDrf+Qn5NYcEq1Pc3/T3x7h0gpd4M0PVrybJzClWXmlZFPGpOA35dAKP
WJfS50hFRf/SvkjM4jEK2PJyp4vo+9QlapSymPhId7+Toh8NmeWJ34EIah1Tg6p9
FXDpezhPq2jfe/AqJ6WKZ1YObGbWKrJ2/075yqpqdyGuaQsdOngsG8k8nVkzrJOV
6zO6btmwFpMCcY/tmj6cS1NABMWfdeLtcGB/MVSLfIbPViufbTRcef/gCHXwJbIF
gcsbBMivqOsDPGa9gfdm8IP8CbbZgOuuJUuPjpvHhqLG7sXNSBWK5Fyf9zonZfk6
cWhdh6cL9dC2Cp0vwp+JH8YGYFc+q1vQvo1xLPJAGPWrFOyAnVeMatSWOG9vnbgA
EnKwhFjIpHkc98yJOrqtRlQSuHX/qt/92voF7RHWMY57ZXNu3wWYO/ZOUV/9Bnw9
B3kV9Csq2g09ugivtogginNB+yPvkb4Cf+Ix8JQZVj6oTlpFLTvV1KWQpdG/+32K
KnTsYwTI3t5YMBr11YVSoieRbzVtneQz5fdUlbZHAMgnWA2rZZzrwQAZAecCJ0Q2
At83BlMf6l5UgGYg0l1FhkalNciNIdJcNurb0Z0nrWy41QgaH2Lq3x/b5mkEbP7k
YHYw1F7pmnai8EJPp7khVH8yFYtpi1yEsBRKFWZzIYELzjy8zUegXu8+PwNgcD58
OiIPUTqk9bAKEjCMr8p1kciM0lbSYrSLmXifb3u0215XHVn9hqjAJe108YyxJy+u
cF2TC6NBFqyGXYpvWYjJ+mpd/HHGSJm/ta/ca+M+gcqRDPaA8hE2aAAWONSOVLyY
LPJYvJ41UH6xzZ4b6byFMQxezUk559lzuMMaFnM1rXbUOsil/4u6jhCvXR7qx0s8
J2BW1w9wCRd+/WKlqiF0DZZB1zw395cmkcwS5AC8DLLes3t20Y2PpL8Elf7JDBWJ
ILQ1YIpjMkm4kwfKii9t9Aq8YTLUmS4RjRz73ReYijQZEeM/2ZPCKAmjWrJTrhOI
ymniKBn2jFwhOUfhR3Mg2vwFXceuBkxBwv7shR8C3jlS/zunXJhPZw8P/VIihy6F
+IfSHPBUGeacKuAbSJZ3b04GnjOpppEmBMEd/aec0XU/ZAjsPF7FX2mLM6uo0ZKB
kKU6poP+EbyFdc7DhUme27XZefyP0k+ykhfMn5og2dMZk6HE8zKT4g337RlcSFkf
MH5fMCVZL6N2g9bq+MM0w3uzuOhMBUF820fEK+saw2OhnWp9qUmjxG9EwBVvmsC0
68V8dTB9kftCOOQe9FAMdXyeW/0IUiI80VpqwF7MFiNyFuruJFh7z4qye7RCzWyA
JhGYCqigOUYk4FG9ntsmBkt2Ifwt809qBXSDiG3SheVYWNJCn75IDF2ZGiIppb0a
NfXZ56m8tlG1pTmL+6IE4M0Ckj/Vp6dKQuYY/xQql/MkUx1w2Ve6zEHEg7mjXa9D
mR6ZT26may59557ppC0R7MsrMZGlexfChEC40MRyAMUuvClL8z/M6JnjZXZhHFS8
Ph6UBnk82Xg3SJEf6yFcjF27AdhcZ27lxHcXSMS2Avt62rjjeGbBdAXaMbhchtAQ
x3dVSeFTl6FVvy0PREvOYu9z9g+0x2d9gf7af2FBAw2ar7BXTmaNy7QaE9WIaeJR
SZ6o6nTOj75Fkp90vtCT/zH4szce0GhhQlY73ucfn6Ju9rh4M188uK1IG0h2SmnD
2RXCGChLF09i4Dq8OzuFjzhce3gjFe2024h+99bsUXk4SBAqv49aOnKzVagZjJoq
ly/aLVMfJ2BNkFAlatlvkjSWBijuSjh3BCGhFUuAmf4lHIPpHcaqYbEvyqmw65Te
OQIPJSG1B7AmiDSij4z0rIxcs1E4uyOWmCmVRsDslbTByd2TD8AdFCZwtxRxUaDI
f/iKcKCPzH8JhQCAEkrqblJU6nFsh0pil6/HEhaOsrfNRbgkDdOINPEmVHbSTs+Y
kvirkpUqznXGa0OOOoC+Jo8/xYNt5EXUbPZ8/vwFFeFFAcTCem7DxM4NM25LZpX9
kbYxUlq3Q7aNGUz7xGtNgeo8OSZicCu52nyANmKhonYROsLAyzo4444/z/cYZrNv
UN0Z0i9a01QHbfmNQUEK/3nndq3sRDdInDeIq+yNzQXd5DjwYH47AszQ3lQLCgNc
oS1cPkL5MT+3aGLzqZeeuzLh4lB/nQnHGwBPBNQuhexv8wJ51Js6YxzXKfOK7tCN
qhohmj+nVJrkB1WXBvhZzMq3pw/gA9WxUhdAkhiBSMo3LWjdPnf2YKf/hIgTQ/JD
Kx7P9KePDzSiKHn8ZoGQNKkY6/CR1lTs/5G6TXDy7hvXlq6BLDGTII9oDqrKaCm4
2hzDbCgtr4Dzod+mVxUEXlj7XnfZv/BlThiJA3Ov5suaL+1qRoFw8RTopnEVtQ3+
g+QDJhhZTLr80OThJlIORAzaO6E+5jhFghUx8COMm/gThBRmje1qDu6E/Hd7zIKR
QK4+hJnHjAiik5g9uRZoAd4zZRekFAHBCFiTE6MAzqqDTRpao6QQlTuVmUXsCj83
Ra92IaU4FSm/CzFMoe7ijyCsKVWi+hwk0+Kio4MUA4mu2Gyq7C1uwuV1banA4QrR
KPWwQG3G0YnT3PnFlgHAHjViv0AY+xXNIawwHvll89+aeXoAEHBPAgKAWzOpUtX6
+UCtEIgSuDny+hC9o8biX1uEDxzSb4uA4UKx993+V/j1jNhNXkaPD3RjomI3Kqpe
bTlgEnU7jH3L6GO+tZopbZ8ypRNJL5hFlAUxXr2E1vXGkiU+/ExXrOXFMD1ayq9t
TbONTGXBCRBryRb/nPDsvMVxRgWxMNrLNe3sIPP/i87KXqn9uthnhldLRSRdf8i0
Eh8pMrKspApIfKuGEoDPOkarbtcyP9KH4hzkhyZfPBZwu7eVfW630xJ1+4Y0lomc
s/TKAD/wXBelNFNbzTWbS58ApKlpIZzps5nX9nkleXSggiExDLIuEmRzE+ONz+F3
MkRYpX77J+kWrUSrVIvTHXm1txfbVC0gJD9p/uBQbihY1Q+nVTi8ikO897hja6dC
LYbdBEb2kThPIbpuwc9hf2efCz4th7BSbZXsLcLxib9CxjJ4CqALWCpni0kGyPRd
oQuaaTxF2Zxr+2FbGl2QjQyjyhATsmZujr2dC3mQAK6XNsXJlsSM9C1IzO+PVXk8
aPj2aRSurTlpS/64rwQxOVW32jUM+J9gdu234fD5qrB9nhucZ8z0tIT46xnrNdRM
Wd8zg3G2nc1L+h2ZoQHaz+CAvgN+qFnPh/98o2uYvq5W8xrbpj2l1anyoPuMpuP2
bgBpNNlfzUL9gZiFYbVwwfsluhiqW4OFACPDF2TCaDzT4nQofFMDyzNRCTmULbFu
6nwMQwDHwFR6J0hK+hL6C4zizDu2bEta/CelynRvecvRX6KnShn7WLBQWqCRi/nG
NE6yVY0+0JT/wuLmJnB19rASYaCzKu/7PI/VtjAULpG+OtI0lPsnyOcaEvA8sMY5
k3sBz1N39OrPR7lkHon2A01wifBh7Y/qsYAu0sOwTXZI4yzzpsZduty0+B1yS4LI
zo427d5xsZpVZ2NNpHmhgrua8ZJqngwkBRu87i6Fa+jCLIAx3kto90wVn+psAx2A
tEMtKibwhNi1mToA2Usta/G0vocq3V5OBbNob50YOrQzVgKUHTVGSqdll+e74NXG
Y8GNqOAqS3FuwimI7+6RBkCCKz4/Wzqn+toSd7IKXe5YjOwOy+UpNFMEp54YWrZo
fj16mtEny6bIa1wSd260xK7fqo+zQN0ZjnAG9zarA3Tn9nb50rLXV4S9gYYMrxdR
tGEDTj3/ZcBuRk/lOb3mz+bFpOUcgmAPuNlBXLZ2NHOe5OSrJlXtjSFqDPu67D1/
dCvHZSCMamnoiQtjHOAxFvmwEmFebEmyMW5H4QWb+GuXt4xtjM6SaLwe6yf9Chnd
ApHQmlOfBOH3htbifuZPZP8AzRiDZqJKJg2VY9yAvUicwX9B0g25yS+fITwPHvaS
7V4YIy9Oxa9L3gG0D6rkoqSkg3ES/ltnpq4vBbpUenrBJwr4uR+ky5Oyro8tQWvm
8QoFKBA31s76XzysWzG8ENHM/wUz8+nMbyCAyfFjDJQ9nHaayVbXQNUhP0los2nc
lHMmDmgXu8t/8NVBgnzAxz1HtZVrfqrbU1Xuf44qtG0o2Srh3nsPoEgF5Muzc8eH
qRGlC/4S99A8Ae6i07mNsJ2fNtL4MhnxuQ97LQirt1XA5aR5Uy5doF7sxp8f9p8U
2txi/gl1CU9qeqqR1uNmL6+hp+vVea9EoSaWBgCD51ijH+vytnyfUaqu5cj1vNPj
tpSN4e+EVI9TSNx+TDxwf/iJFkf3BtRuozR5+W1/bVT19yrfh6qkHkbvOwdSwihp
Cxghg/tN68ppl+Dnw5AMJjzSB4a3yKhfBgLiiPT7j9jWlIG0Nb6JivqraHLJfBpQ
IFSDCZr1z2BFS3xWnQvVB5slxSkowcDxM5Mvz3tgklPnOG+3bGZzwgpcU/rjoUga
IVvZCLzuX8/RMcfp4Os+JiUkIQiQZjfK7MPbVYvR18C2VU6A5Q1GeO18AMYPQZvq
m32S0W9SsjPU3uZMlg7wD3IcIxWHLOwKjb+9j7fN8etiwYl508RwJa2ayhSeul5i
/1nGn8kCoZSAHedFBQfpKBFqm7XdhAwQ4Mfdt5sAzzspaDHRNk5Yc3KyESuffG9i
vOQ/bkTfqNaGnbIfq16r4h3KDCVsnuqVotKSuHxikh2Y64JHLKsFDW2DTRUOPrTO
E89PPH9oR3ZgR5kz+cHJ2lCQow6TEgdfQI8Petnhi9fkpjJyI7tVyR/bpvPK/W6Z
n3v22CUYEnlAFzMo2D5l9Sxs3aYhIu+wBAxfZMLISGMNwFhEV1ssRf7kv8tJ/ugG
muqdHulO8BerngZORqTPTmGo2a4E5OSVpNddHV5PIPUD2ZvMc50Io9ExEiOhlkSa
JDtz+QBEXyN1R6RKHje5NjX8o+FQyLKbQauXiaajzo5cHTdi2GOBx+mFX8UZIdXZ
FknimotYH0+GrKNpIH4TqfqO0qLghVco4UPCjY1/OzwwSA6cxzWVJLQ2WChW401g
OhBQMC3jTOTkFyobFiOhDBwYN9NF79F4NcJRfXQJObmOQ/OxOupc0VOlpcyQlX4O
05RufldgFnAUno48Lz+DPcL7ER1E09Ww+jB4a1KGYDpm1tstI6T+ZEDFHgcmAp1f
N6vtXYNNG/+Ukk5dlLdSMlh8Grsdutqk67ZARjCrv5erlHUEp0k2r/vQu6wQXLyP
Bc2h5rb0+NG+AS8/iq6mIwEY4X4mTxICtIvw7blcRggIQ4IzFdSV+fhMWtPVVug4
z2vDY5cOSx6VYmzMuBBGCNb7eAz4mUlwd4GinZEmxYZ/Z75XpqWIlOM5U+yG0NX7
/LdpoNVJlcxZfWVj2lkXdsDMPcH9taxi9P3aYDT3O72v8WZuk6cyIXG3fsEWd8Eo
YvyTHp4G+3eAZD+y381gjv6IR2fYPRffxms00OTyzPKh0kkt+kmjtrC+gOBfzFVU
dQ0Rv/CB1vXSAFCa1DPep+1zfxPLsqVa1LjmKMNhV9vVDC4f2jUBFYbjYWEulPO9
8VI5XXwYi08muznxxv/pS8L2UdBdozuFFAzcDWk9T4ed02jezYUhMULXEwpjd9Qd
fGpeSaMn5RjlJ07KcrQIDfUzEoYN+ZZO+Fz42yitR8JB32BoSvDwqrzM9kSOg4pc
FLYIWenGZIHZ2nLQDudad4J8Is0lxKbOgc1yh5d1+iPXx5bTKgiBOIlcaO9n6kV/
SMaEg8BgtjSO6548QSckTWd1J5TosyWExj3KnqRvCGpZ1+ZUgkx+MngNKGiTXiYm
tjyE4U4hYV0Pr5im6+lEjAmW6DHYvCVfA8d7au87m8WjE/OjRoDJ7W28X0VEEapS
btzI9niucW2BO4GmibLrGunkgaGYNRE7myBQSFDm+IvQAym3Kg7qe9G+AhJ5YVbm
BZveIW4oZGRBzSVuuBo++1UrhL/+ZEkSZj3oOitc7yII1PA/DwVKNoXffhpXq7eu
g0At/m1CocBMqcswr6QUP9TWY9wdgjDwQINzG2vlGUqQZFAQy8WEvoIsED98wLgL
P2FlI32LWemabGwQ0x5MStEUixN+lRuIa6oVKRFVrYiA4wx53w5tDmLlp72Ty3jy
GEmlP6ast38ywwWYNcrklsFH6HEUv7nBu6s6+oIfG/gc3C7lmtSPowqVKL/CLiti
baVzWSHwlfMm3iYQ2qR3oa8B3v4dWDxSCel7cwM9Soz68txqMjmgR9cbKtyl7YlN
u3oBixAhi40tk0FuDJJhb1e75oU0Ml/nIkYJnBsIcLy5S7ENraMh0ifgi4zJOrFz
1xgWe0OXHPYd8iWdQQRK0NT924OmGgJWVgqAa8FvRhC5+omZc6L1Xbm/2xdPijtl
YsCzINKz2qfhlw0bNq7F0jCxv+0eweNh8tdsGSluaf5ZEhJpnZ4iqh2DnsAWvfBw
pnLZf3xowNgg7oZn9X99FZJAGqXvN5ShbO+CWko++MxcziUOnqS1kasrWuYG/c+e
ZXZcuYj7pWqUTcC76oCbTNnwPNl45iBZLPGtvw9OmrgnaHC2CKuNw5a/30Wb9o/a
gWCsFFqmFjXPFtMfsBh0g2iPgx6kYkbUqSpMA6oHj87633bUPSLLjz+zeHE6XjLX
otQmibKx5CpiB0q6T7eOKl8nHwRH/HiNyenGptbdqqRpTpuJXpPAOcdGmW0ngbUE
3kJupJM5fJrEdRLdN58ocU/TYfwstzLRv0bIamFBAXtp3OMV3xQYPPTJvzotG4Z6
bPmX5WhRT4ef2KwLcuV8dpFwIs+DR3tYbwkir0Ycwt2RVSkFPLN4+Dgg0KqlHIW6
0quWl+QUVJnXxGDC2BvABE/vb3dqQUGZRLkbuxVPcUd9jBJZ+vpjlR/999fcEbny
4Nbhq1wexkODFNXMP0QMLWkkEqeY3eN/Oxz1a2FYhK12FNqRo/j3mOai7kMZZvs4
CqBAnj5OOV0EM+03Aj1NTLDg0z4R68LCXCdE+pkpbpeymvcxqPqZC/MLD/CXS3Fe
QrsM0UjMI5FuWaZIZgHcnxov7uKLqWfKFrTEoWJNursdU77/T2PVq6dEybfkp3wQ
x8JE6t/uJTibsy+vUXept27Tj8fhrq2Md6l8Um/a+t/thkDJQZHbqBY2MdOiqE46
Nqc78ozrZo8OeeA66KoQTkrZVFyne1exa1dizegtSEF+R0jZ6V7xUVA4ldZMQnQM
vF16PeX6kYptGQnR0lSbL2dOjbJEO4BHKV3EWorYGNAvYTESpOkT8phLyE3oNnsB
pZd7QjpxPcQKMbK3MwA5gSHnQdsn9kO4dvA+Rv8/3t+V4NdE6fZapFkQvjJjwaKf
J8W1kfnGq2B0xHLZekzHcAj4aR8H1VBtDzuAVMIzjWFfTqfpA79MCGQOOMZZ3Gw1
qn3t8ir6TIGNHj26BWVdxWKOiVyxGAjNx5pN+aB9B6qDFtnpAYWLHaojcXwqLdyl
ajRU3xRUeIp5Kv52f751HAsmRqmGob4Fy+rL7MBnQQugASV+rpH8HtG781ZzU9sy
8PshpqRiqZgDXiyISN+EkoakljBHfnUPFjKSCt5iL2DoYRXybFAYh4k1Adn95wVM
1xSnSrVSLjkpLNZah+CvtLIJnyJ+YX/CEEqocERrofEXcpQ9108diPeVOPpTlLfg
3UF2/FtgRFGcVLOaVeTUSKc1EOjEaizSnGI7kZUugbayjtbt26Gasigm+Gm1ZPSa
MMjksY8TP2eMYXnZQtevjYT40mJekFXrZZKjhkKQ1dFXKqzGSQ7FAiprIoHmXvYt
PVY+Ht1te1sj2Q/pAV6dAHOr/xczk4PPbFyfIM8de4GdGbTlrvJcmpSnn7GBo1AJ
gsaIO0SzBwPbWNOHtGCvUhTgGUMy9MqZCxURFjmMW98Zuq4ko+ZRniHYX8izHS9Q
uLOUOzdGT+D+FFakx1fjqelEb2R8EQ2pJgHq5HKWX2vNoalt4zwClEde6OzzYy86
xBneAWxQUju3l8RE3cWjQpnAdQqiuLEjxLjvu53drfYTisB9Us7BscXS5b2Enpfg
snMJiEEBcLCdpAQFV174TCs6YwbLfuiG9CxtkM1pg9eLmhaQxqadiHDPkMTy5Cis
VeS0b0aLwIz9VMs2UYvxEECBAvoGRjWnqs7b3MrL90wyBe9cLRfyD7RyASvfqQwq
ph0w0OZMgoiABICFHttTsOOSvVoXoj42g2wC9zXJ/tS8kVw4n014hA290eQZKvpO
sY1Akw9C0Jwuko8iLGeRjKIxu0eE/Vw2Cm1niGlSWdgDJ5KX3Cc35OqcgsS4FwS9
Nmoix8C9KvGCHoXbuszl+v9lCg2IHuR5EtMOArUoX/eeZJhcC3+54KisbnnhutZ1
OxWV9TimTkJnlMPpSDi2HT9W0UZmqWFJjyDGUYkIkXOLeAwPUQftdkDECP9H9X+u
naUP3pwY2PFklUTdMCacBX67WimX9t2lVpDpX0uzyMyFfP8IBg31gTm7E/UfF/fK
3YnC7/uzhfvsJdTqKo/934xcOeAJvA15O2FxIyYbU6GsgPSd5+6G4I5iNzvquH0W
bMkdDdWTaQCXB34I3h41S/TiECc76n6sae084S5oA//nrvfAwEEmn/Kqm+3dr9Xb
utPb3YVFpxAxCOPD1LDRC9vMkqlYbpmr3NeNMvsP4R8dHkf3plkRcSkxkKlw6RZ1
FtI2ueC5DK6RLcLVSBmNd6XBWyCxMcNq40JwHcTRA4BlQFBRg/HpAZnLia49Y5A1
pGiCmGJSMu4Hf56mvc4dNW5cCgDc7WUR2GN6qR1w4GsY+aJokbwbvnf5i3K7eLGE
AmuUt0wrfJUzBvMf/PtNgienaOG14t8NdaAiq5B6wNE8ICgljRAfjQScSzMto7xA
gy8oztb0GTd8TP6sn/+RrceybjLuntk9MwS83tyxF66ltaWj5YiAr/Zv/xM0bt8F
/aeOiW2vuVG9LIefWXCv6VQK2FTXDc7wR9Syk1L0wJd5mw09MDp06N554hFFR2eI
wTSN5JiCD13VmHkFfNAkxJOwJUXtSwVqdiqze1I+kHpo/roN76usPC/pHuUPwVTZ
XwecjgNvHlxmQO3YlE4FfFkuWzZnhn8QHQtuwBmy881lbG+nez1aeZ8VEpSm2xYn
7RagKYtQnjZlQP9HC2Mw+wWRlWNLI6YPcQ1vdEe4qXgZlMyBL8Ja5Ks/S0LONllj
5XHnWFwVE1UwexU1F2fookiUTX/SYK7jyxCtrVLhkkegGBQ9JTmN7z3p5cey47pz
yKPbyqIbZRrrG/GRa4GfVh+4EtFOegVl7QG+6TFN8vFMRX7Q3MDOYCVrZ1IU3jQo
B7sINsAIrq1xKhz80hfIHDQhh8q54zmtlwZSGWimlMWLYZYPc/pJUppOjWk2D6Jf
MuPdb7OWqh9qwlA5jxkG1UiLpyESJMTxKvaBtwhQ/n0UdSRODrZM3kNArOevMHoz
yxHW6dqliWhCgAi0FttDBQDhk40SN3a7aoK7W+TVNEKRH7FDfLjJTXnXSrWS4Qvc
kvonNEk5iUrpUH01UnSBXPXzdumhNsbxrZWEefPked6fEp4CTKPBezeIrwsMmXKl
0D4jvtNfvt6mmsKUEaxjsktE5li2QB7ZNRF2Pg9bpiyzqBhle4p7Q+4J/37vdKXE
wc/9NO9PCwOyYFR8iBSupROPQGFFzbnAyLWTYdxlQ03Y8ANDqLVnBLErCnShdXgo
5Ki+i4y3OHdod4Evl5ThgxlUb021lhntWKk6bEgq1wSig0YaltuwGiElC9ATJJ4U
C4IsVp+2IX+CRPEP/HvxcklTc5Ve8Ya1quwg5Ke18xRPayOMMRCJFEngEu5PjK0j
qyDz2MM1j8A5EnXjActMOSK5kyn2+lGawYOV25N9w4JNgzdBvVs347UxQU+Y00A9
vOjb1ReMGbY2yc7rtBSU/K/lKLJxCkc3TbDewTWPL/41TsUj/tPgrk4N0KeOLr0/
Bza6WUnRNIJ7Rkws8y/Nl3jAE0g1VTfz0c95ZH8gGZ+wb4ILBCNMPXw6ekJBoyY6
g1E7AwxFcs/1MdDkv/6fAFeHYRZYvV3QGFx/RKwLCfteAkV/pyULyEpIlLH5I5Y9
EODlVciy2Ogcy2ym43RuVqki2QVcrRiQbUcWEkRm3/LOW3WI+LWhDzGN0af6ivx2
USLON8zbYwKr/zLKVJMVr3awTSrnlp31DGz5g4YBlLvfVnQF5s7a/ZOTFZZpSXeL
/6Okl1mfwIDHYMZY2NBGCtpBhJcZlD+oYEkWp0W2gjsrTIJ+J7GutdrVI3dZKhvn
lj5reFaA58mYSoeAwhXFJz7cxkfBQ6D2E5AlH8fKKJ2fwzlGJ85jb2uULAHZi12f
cHBvuqyJGqwj0lp6EbETTRaaruJtY1XoBz5vU3ph12p8EmxyCo2uYL4y5oll4oFZ
QeUe+2D1g2ZIxVCEMbB3B+v2ZsfY3E5DCGlnD90/IOvDjLrJ7/0gIfB7C3HUtORL
vmBRlU08GIFlHU1+JnKALYAd83LVoVOYestu32yaHE87BSbP0otfNMWnByu8UYlT
hobHou9GQePZ/PuU1WAE7kYTxWhvt5jQFb0g5FeVGMIG7Doo5EnbI1qxypIqqXey
r2cjeYgqK7byfWIwCa/tm/Vt4ZxAlOUs190NdaUrK9miPpyqlaiPDmeG7YX4YnOv
F7s6ecJhScXRTjZ2LP1qKA7t919JiIH6VUMSRNTPFyHKDE7k1B2Crz1CqPYPGh+m
+73uyvgyAwQzQmgstmJhPyr+9ahOQncoNpe9JroEGINJp+g5Qxe7I5x3GRTLqwKR
GjWakHMJ5QJbFi8PqOlSvnWZ1T88SzYe92sW2ITan/MEXTLY0FkCaqiFQrMGRp+7
cHBiAziaxQsZOA8RgqelWWBMgt7Jy4C/jVKGs7TclXdq46TQ8j6EDKIdUWF9vNo0
cXbxKLtfsM5uvwfuhlYrOOsSL6pG1tSTfiFMCcNo0ywwC/SnusL7O/zbmxfc35hN
9w2PysCU06JxI4wtGrJmqUZEWlRFftdCdqF/8OZJK1A4d+avQk5IuX/mz9kBnLXl
g0xxKR+4ufHyjw3TMhxjKiQ1Zazo9VIoUESoJFxMRFVQAEv8NEZq380JLWN5uSek
oB9oBBbPDM6p3HWbtN1b4s2QP3Cy2a/TCTY81Z6bZDHFVJTaTmyV/rRDbYdYzfmI
uEFGb41EfJglL1VR0N4iycGX6r26mVU2cmXQFvHdmte8aKnZ2KFBR7wrZtUr4ale
+ZrDCyDuG/18Ug7D1H7aKD1QnfJunu7WALdW6VwvVhaeJbOwbgiQEN2rA+rcUKDo
LIBEvET5lDJTr6olBuyP+UT7kOayz6JaROgWZ3NTPh2OzZGcAsjrKAlV6w08QsrM
21PPwuvcKDhPdfBnGj/kXm5HeX+vbiY9QhDGwfFadESnh0uDbFU0EyPcCekUrM9V
pBoqURMShPkf8E7mKQd4zc+ZsZ5qchlzCrfOKSc0ByLdy6zDi7yKRTY/GFgXy/Lq
JPu/WdhUzINQl2p43UPidGvxqKtDCj1eFbHMQD0ooGTuQObq6MH/DjbCGEqltall
MUZDtbmPrZgADGTxv7qOG3umN1fVW/SylmGmhCJq7AtbQ6jZReHIyfSE3JIQEMe0
v+l+8NrQ0NA7UjpNswD6REvrTUYJ93Cz4KnFmZ36Kl5ceASMUgVylWjahkJS10yf
2FTf8NRq2h4ip9IX6MapesnPRYF16IckgtHNh8QysR3dBMLsvcLuYzwYxlLD0NOk
94BwprL3jfbfICjAixzxlsdVnxHqIOM6V24XYYCtrOO7zdqaXM2o7O9FK8lpSpLp
GVJec4nXbC4oWW+nC1WNOeX5PH7C/gEZt1rJf+Lp/+vy8nsadUC9Wzb7DN7I/wqC
XqyeGZELbCTzf2vuPT1V4E1AcHcwU/9Y3g/IEXAlksaq/5vHL981IsWm6NIoMIpn
iPBNS3Zaglymiq9pllgDnSvbPIgTwHVWBOuK9AEUheRGLzMlmbFYL1FnaMejF+1C
Bn0gyOvEfywqgbM15cShbmisgC2ET62AmyagWpFfj3DuzFBJmNRCODTmQUQaCtXl
LxO2/FInnW1lEEZTxredOpltffxHQ3idzsJGIdhhIB9uNuJRqKrzyIEKGoM6XlxB
kM8Tx7JOSpOIiluV0VLH03ynwfgXk/aEwPq3f/808moHv/9nKsYTYX9igTsJtV1a
gMLkZ0wcDbbLobe6YyeoTOWluHxA0lpxhfad56bPZLKEPfSI8KSkyMqPwfCSDaJQ
ac4wmKXCzR3crxX/op+wGiFyxszR7mx7ZkEeGaQyvL7BcfgG8wUtwatR0ibnYxNq
gkxIG/oQKnfLZm3Bj4tdREWMX8t66vPal+bi7xXZBofr8DlqWNrpMa3e8kzMUHPc
lS0LenKRHOmf43rsqr3FoGxAqgs0sgf9SqYDsrSbj3FilkpUgUM4FpHb13hHT+Hq
LqOcZ428RfCUCJBTBXZJPx/nwA0TKjnb3o1uR2/KdAEY63yGd7k5S/elmo777uwK
3v9v7C482Vxv5to8Z43OqrBbGpg8aM/XrSm6BwWbZ4r4cAAv9jSoMfV2/mts2XGN
/Gds2JawmXbKrQjQmOokPf8R8L2nilGjlr/epeO2OP2gXIVJZdCHBYYR7w/KAIAu
/gpnZ2Cuu0qHUX4woUT9AFmIOxwWRvfeDNzakkW1GIbTJJY1qsQyOa2BZtuxUPYG
INoShJrWcFLlxM+mFOqxEF+pVKl5fgP0uVK+8GXtXNCQdCPUITZG2uFrQWRa84q4
dwjwB467DAoZRuiMq10DTf0GGxnnKp3jSgBXoFzaxcUO4wmdeq1Yy9I6HbCS1QQj
z9tuK8rINRjsaASFTQ5UMI6Dt+G/mAwyD7fov74lQlD1Xi+TNy5R8KiSrphzSL/c
/ovNcEZ7N/qTFbRuJXkqlQ9X2StPkBtGWhtiy5w3KpSkIKIwmhWoeierrHdhlCvQ
YLeDeVxJ+uipjxS67fWV6m+8fXF55HVExU2dHefRmqVWRVSap/1cvAHke4bbVtd8
oJBN45aap48T41FuFQxd2pcRSHw7Z4XbCIBECnW8f90oygaudJ/oFuvFr+lUArUa
kjnVodyY/YLTuEaRbAhWYpRlyFbpYYsVTiXdgQES8CKNCXSHRYO1sidOlh3hMyt8
/xC7/ZC96VqjnuRvDrEh6juJNZ1yjszmlJsIP+HHAjwHAT8RBegddB1sZ2E+DbSq
TLcCC2tNtqT0MyL+q09dVVcFvLzmCXjVkCpVMbLHimEaVKlNBdMKX5CrojbyCqYm
YU5wa7w/hy4FL4Ue9CZh4z4bF5SbSEWJfYVC/ACl7u0stKG0KJMc1bRsOPlWgc1a
+QY2QHIb1jkve1wjqlp6WQm2q4dJsE4kb0YZjB7FSrlzNa/+CWoTS3vLAzBGpYSp
7cFHk5W3UTeLe1wVXAQnZrToD9h8Y+b6aVkG+vqIqLom7+cus7x0vJMdkPxAAZWB
cFkK9ZxEOdbhlElCrHHRRW1cpXcvAZNtsQWekn3QOLcwfMb7TDDGyR3pKhfx/E8t
y+fXozGxSGI2U9jGH5uRZbpSrIvAAooqCn0Emihq1TFyaL2MKkUigDupzPcMmJde
Iy07t8WdYvrK5+HLbK8/O1sw9B6wJucB5hXFzh3/heKB171JVhj6D1W4UMYd+l6q
p7AziMs82/3l2ym+tT1buSFC/ctu8M3OyWpqxd1xS1fxdbfBLZ4k5EVRPkbVjpqc
U9tmmnHjgZ9Y4L2xQVxY955AQg+Epp+TkQf6PJBorqwvRklBX/0Yd9r7Qx3PN3Y5
aD7ZffiF0xYjl4nazD6WYq1o/alWgMyUIuGRmoJGy5uC7jDBXQWvHMNulRfaYBEr
TesydCKdGs9D9y+ODjS/QHoTXyrCJcSTtCrYLelHIz2FpW2KWDBw/mDsvvTbEnTI
2Tn1KOuLb5IJ1VNZeJgPqL/UE9eGQy/a3d0BZhWDqZcYF3GXn3aRW9KZJHA49xcG
iFm5WbRVsjVOKiERKNmMU7/AR1k3ez9MbIMEGncN6JUz2uSz1QOpL6s8kJljo2Gf
2hypK/laFitnXV44UFi1hmm8HFQR6rQuzmBaQiKg5R0lZT0ahv+aNq9KLd+9PsBX
+j0I+NvUq4inn0Tg21+t409V9AMXPudvCl5LD9rhI0SwLIEXPFs3GUdzrZoyDyfn
KymP/rtQn/dXb6n1rx7rN/UdklI8/fBmBWnUT30bvzHh9jebnA1wtzcAMyBxLgCE
8xakNYcM3i5lO+1kB355frQgqf0E4p6VmsqNqvB0wI4Bcy/zoBHQ4ytkLGEIX8it
1YgU95PYGMN/5268WdY0eRBu2c3NqI0lE6SjLOEY6jwGs86ZwjrU6h16OWzxtKIJ
1qSvHxHbSAUdXInKX5d8Y0Fj8MnGFBJgBcPi9IibUbUCj/ulGE98NGrhQJdUuZs2
eNGY42GIQJ5a3opDWx11BRl+jBiYEyiR48UqdnrZ2lbekA49M2out4THszPK/9bh
q1Br+D4I2/5iSzDPael9i4Fl5flHevb06d8s2gKEauQZriaQysYhPKxf2QqkEY1v
FcoC5FfkQKTvfwwygIshhGSOp/kaRkhEPzqXf5uPBDYsQgHoEGIK16+ns9IXnqWZ
/qkwQEge+pzHH3Is1REZwxT3r05DzRZ+LdS19buP2noTzAjykQ62HZknYNAXnBT4
f29Hxjtjkc3XedhAytyEp0SwN6uDsu4aG24S1enkKsT+EnJGWOq8QNtGfx5Ua3np
QA4a4EeoN/+UrsFKum6mhvBSqh9W8auJE8vl9Pl2sivDYXrpqOabN69Xdm9Iw7ie
QFqLDlC14jVgqxafcgOlH7cKGYLyxZg268XKnKszWtgbbvjnUTWkf5mDqcVjDipR
v/2LDh07NQW03+TfRaoNLViQUb2xe+mZdXcNZloiCzwFDuf8Qj9K8QiiWUFYKsHy
Qc6evfs0cydsDWJj87VQ5XgwWuFSqTy/mXeSS2BUcNKcuZnVLkSRFjt0JnRoYiUx
OP3xbGNOBU3U27MzjT8fDSoqBwOJg222G9VVhpjydKfrKgzZNUiB9MQP0pyVKShX
0Xp4/kqY6pn2+KHq4Tqe/NcU3Y/NaoIajr1PkAeivEyhjQnvsxGuo2mK+YAz4J7N
zhZGbONvsVVwXA4K+grFE4B//E1WvnRNxvb5dkHOHoFLCq8jOmEFO/TjY8qexRWq
uYvjtH2Xu7f3MYJDqXQbXGzF1WRtVDvYAowG5nWVRYbMYnbp0CvB+HFHW8cZwK1z
tGZWFGlTf3Z5qKwbNQqgANU1uFmjyLPK5DcVSzp7L9KbgSC4N9f69ukTawWkpNit
A0U+7FgWfCWfmn3A2r2p4IA1hr/iMlRtnUnY2GsAeRSj8TvrCjfv55COT6eL/7WM
iFme9MMVicyr2w4dJwr34ILfsISR8qVynLDPysuY1j8Nv05TZ4Xm0gH55NBQ/6QS
lX5fV3dPVuB9VrKWK0Bz4btcdLrQKn4uo1yAGMItDm7Q+BCXDvnnuDQhbZSN9F2d
gCD5zC6lokdsj4Q6++ETAJVUpAzJvnLdAuIp8pNHVAv3wYAZUD1f7ishe8jKSJPd
s6X0+YXzuxe1EYld8ayIsx5bLU/F31Ia6/n4wCTj/kW+v/jLpB4MX6o5P4ZxL8dX
fMjVIRuKFMze1T+9LO8vh2dU6pmuRU7NC5h1MoQXW/VSZB5/dptTZ4P8rbdMWO79
fjf7hnKXN9PqxidpGKdhaEleiPjiGDG7AFHrpPQTF99uVPJk1QErpjSwms3JbGrc
pNNMcxifqEQhmgzGnCQyHUnHM2a8LP0WamjwJVcLOZJXaAy5vmHO/GKvc4uKAnIG
SS2m5Fx533DHxoSpKkiJ/kIFSrxm6oNHMBUL0N3iA8TRy8oh0THZ3gAfzvJVdxxa
D6/nPGjUhdGqQjwnaSnez/WNENtdR8GCX6n5Z/dLsEeCawB7MXvjyKi4TlR7qflE
rfLL0fG2j7RcIYGja4CHY0fSRpheSDsi/16l6QRqBniayJPWFl3uBLb22lnbnCR7
y82D0sPl1ma42ytHtycjpWfhxOewjQ6ejq9gfd6jFbKLs4Nmu2/0XPi1C3khv2UN
IWyNYp0h6cXjdFuJBsQ+wxvM0HsxgiDqe/96Trdr7nfhAUxTA0aLg8hhehusBOYB
4N6FlJsVtspWTlFxfIakz2TVSn03VBw7AAuovUEMOpnsnv2lBFn7ihlhB1JxJtMw
+XiJRey/6wPSArMKa/t6Rvgq0mIsputCG5ZQ0xJuR12B1rpi8EhOWKz9iQHiJw6S
yij6AGRL7lEQqgrJV9JyDdvUHBGcTtwl9he2/P6DVh2G1rB9t+Gq1eTAQxKpFn/s
qFaB1I5kClVO4K71dU58ecz/RmgA4pbxfSG4RDSLfHj5Clj2n7/HCev+YLY5tdU7
qRs67/ra/yByDlqPl/UDocTOQikc+mKE8W1NXKmvk2b1scg0KbTvPFv62Y9xWJwz
ZW4yO5AN+XXGJR54yAaSfQjHWg4eoNjydcsL+zl5YIRjIUXC7C2JjrxUhArGM+Qh
rjHXvsO/1sHGCXKRLqLBK3GIFLovysYQoZRW6bJ4sHqjJChKvBPv+P6MSRa0jPNH
GwXnKHxO1guHi7ScQZRKLBxJpXi/xtcCPojwNc8L+NBNcx2vF5T7sVc0HDpSfB4A
Vf30uoxB+Noa7pK9YSkGdyADEwBzeM2XxGf5Eg/501Ik5u7a/Vka8sd9Ra5xAWum
X/eA8f7DmOmEMq2dwWcb0NYC5tndVwmDXizXBzTgPq/gQDIiyInn4m2bKSahJWRN
b0KPfkCch29Q1OR86lVuWonVqwPxOP9bMKrZ4iRpeH5OKDoR/sSXUcVT+TIySV34
deQJuOoqNj+ot2H1ZOaAPF1T7+4hoWuBslkOIRJqL182Uv88NNaSkrPMyH6kMhzb
9JGRpyCYcNg7M8BS9QmupbWHNx95Xahc1kSTn60WERcS6hLB95/tYVOBN/ePrpr/
8ksUii89K/yFU79DmiSs8Fh+dIPP1yVzy9wl41gvfcN3XfmoI1Py2Eoa/cv1AQVv
MOv+QTUzDkYOqQtG+TsStRS18hmO9nTmRbM8ovOdtt46n7LUdTShNmZAR8FFO0kh
6AaORBFeDrQioA3WkF6JdZfVggGcYkIYwPSmGro1O05+P4kcs5+tp0/bT85NA4HT
EAhjAZ/TUf3fIxe0+78tccPiK4ns7GmCvBU688tYPRhlzUgP/qFh523vyx8N6xYC
CMeSR5V72V0rv0LD/czjIlqA/ztT2UY6FAEp6LLjxwlbw1aZk1QlDQ7vOMriDiEw
d/q/vyWm51EFVUM2fHtZ7GOLFYFO4ZxMgPdS5XO+ChmOyT3TJG3WH+RR1sEMwyQT
dnH+1Vpxo4TPUWaVh8CuZOv8BjZeRXlM1WUbmYxF0HY+GD0KvnKi9gU4NvlDlFIL
SFpI6iCRXaaNRZDUdC5XZfZGOVsFhsDBv9tRDDxcFg46YPFI8BF1vMO7XuWDLZ/8
jROCZOvLoQSa3EfKdsq7//CiTZJJ0rEXZfpPzbVqdVcNpsTjNlFxU54a8NYW9fYy
vU8D1Sm4X5Zo6w9PxNCJbyDzruPQ6mF5HXsTzom/+aWu7gkfpl0jTbcC/0n1lb4m
8deMm1Q8I5re9dRQsVwEDC9Z214OukxqsenzX6Y+InMkFpD4+mKESwmBYnBgJM5a
PFm1AElfo9Wjw/yCc2pTrstPR9WA8wbtpEXUoLeBqTUUdMSt4XsUJhSPp37CDQQ1
f+1gVr6e2i/Smhsoytd1L337KiBeQL9BSQt7TJ73NqASQdKmAASYRbjZoHLTbkX+
ladssBnMwI3WG6Tk7/l+1Pop6SqEcy88YjZDaAOzVnDMhG7HSJlU7YUEUU1JLTvs
b8q2xSx2MxUVAx9s5a7hxzMgyeeO1aqpYe/N8hNE6LvyTYtDYLekzKTEtF6Lla98
rdP0HQqE0Wt3qlKXkDG2I18isRLSmjTx4Zk8JrrQjYRkL/Xw6N/ILfvWLA1+qVDZ
Acd+x8lXITfLq8W0fRna1axTOwIMWuwAOY8PafJdoMEyMkawg6n2HXcB/Fa3kHNf
XIP1Ey7Zth0HiEQXrLJEfEV7UnVu/0h12lTdHVDFWIbTXNCFkn24gkpgJw4BLwVf
vCpvB5V1qSH8y4N9YT9W6NYxs93hffCoXWkqYFOQSyxl8wrWAclZkIYx77WOzyC3
QRKMcjjgPRei/mxpZ0zSQ45By6dgMEScd54RZEQH6bXoZ+Q4/qGiBib0Z6JRjzRM
lGhA9mTB+AMjGgGinhByW3nx3U9+6J2pOmMWOf2q4E4Zu/hs6ZgfbvodmJtMYyXd
XuO/QbdUhF+mhh19QznkCEWlJ6FJm8E1SHQAKdeK4MekdLghl9Kp+fDWW9vYD+3A
+9SahWwnPkZZEw9Dvrgwt7jfLHialVilINlT0uWQWKBpI7o51wmO5re9WbZiJTOG
G7xRZyFt2+QLAJoWdNTpNuntD1Ur36ozj9Q2sg/UV6gEjosIpPuw2dutuQgzqIRs
pryQ5U3vFpNovVNAQ8wonVNFGyV2ArL4xWpX7gyo8PSuoZtHN1EgYawhpznj43IJ
xry4034lST+EpG1LQj9ktVoZG/7+iq5Jo3RaYgq3qoxinqP1GtpzWLUYf0UC57Hz
EpTvUbkqbyVVcgtQyqNQasFryoP6lDZZvWOFOigoifgTtz13kNoCQ0PgRG18vUOo
YhWYH3EuVTexEUdRoFTNMidZohLFRMJHT9HLoeZ7QlQT3COh5TCn3HjQsNsK5mPP
ic49ep8HhcfYAtb6uaIG59sj5OGw+44SYhRsIORAzQdfM+UPS/r8bETT1C4DydbN
jw7bSwpRZkvq+aCsCGCeBqfE65DIr3Bp7PotCfXt8oyHiMTGYsyPH9R2Oj5dvx/Y
ykEO3339+DdlRVpKYOKWKLyP1x/WVcc4MffPkIPkLv4ihOasCarcF/L6rcJsLotP
6RzZaX2M/z9RojMxMtJFgQ7ykFT184/DuP1CW/RmISdoIP6wKYD09CRTybR9RMZO
l5HFOa3cg1D8sx+v42X/l9o7dBdnEnApfx9g0TPkCaobdETU5iW0Phtw6z0CeMHW
1hPPoSYsOnvxMQQ5ZM/cZArpHSFa9rXYyPaIW0WGbnXE8s5rUEyzXuFgxl1RTeVc
+2fkfSP+9UP6rx6MFr2bFsT1z2kWAiUfkWfLDMNa0ITXwXGzqQ5PPg4PSB99WNUJ
VVLdh6ym5x7p2EP6vfaq7mG7jbzHUxGziqQhnHUsLcKKypulSm54KlkkXgtLnioe
M2x+Oe0yqOIxAIVMwXL3Y4ogeWCOYzeCPqyLl33poNOObddIrNuZZWvtDfLu8nvF
1gPMQFO6Iu/7Vzvho/pXy7nSZazpyD9qzp5nCksFjtih47WlRmx+NkhaurKEAfDx
Twvh8da7i97kWV+pope3B3JUYfJEqqCqN3j++WtMVSmPSfiX75+vdwg7LsazEvlt
ClxmspO2lClUnr7WZRRJwhNqAGimZ720Qium7bYLeODx2HtK1iGgUcqPgBu7wHUB
Dk4ptBzfNKRPMcvrZSlGL76t7DPf5CNlRKXq9jz7MlBo3swyEeVVIMZ+mH5T2STj
qWF5QTQp4VOtzgibAAjPWBUssnhpW3AFPu4sIdmbVN6HWL+kxoo8ju90VxxeeMh6
nzy+q3ZUCtsfaDFBkbhN5BhtTMazF7Ly897yikGNRdC8ksozhkhWnUWA4g7eIIBm
J/PCoOK618Lp3K5/nBS3ZKbtE1+7WgsiRbBnGdmKSPRFcDJg13Uf+L4xkn31jNaf
u3BZXsZyxY7/9Eo886PRRnHGB+zSdtGl7WHzwYd6pEw2OIKu4F9D4c5REra8VUD3
g4eQKzgpY7MEuCz9+vi3HD9LPtU9iqUWlTFnHMYTuCCsuNOQ8Cs7ruEvh/aiBGL5
OR6fXa6uKEeJeqQ1Jeuvp2zdys3UjuD1JgdLt6F0t4TFnfUSxILO0iBNbP2eHwyU
GBd1SBHqmuq3XWbHhsKn+f/W8wlZAvgzNl2y+/epLLKJrgqJ2e4ls+RYgsj+wG+S
QZcoSwjPgTFMJbE+2Wjrxw3/ZId2PGLA4Am74LqHTLX2SmdVlfgX0yP0q3G5ZsWu
Ga/05gYaZF131DMvV3yeO7IZ3DSGM/dTyvqNIB0VBirZUf6ItGdqPp2macYcqJrE
iBoFkfnpvVhJVRO4+1jpW0hA1OyhSYQAiWCkztiabvO7wFAFa/F32kItYwHBgGpl
ck61xIfX+Ty5o8JSuQ6xh4jV05XzR/CANQFgtj2nVl/uIsBGLqxaqOBuNYKU+Ylt
3By1wMfB/YuAcMja3M3prmqrdxPNIruOhFQNVR1vdWy9Deaf2jCcSeM1ESf4A4IJ
0QwCsMN+GbygALXc6a7f6HYz3zPnf9zCKRirJvZWTFt3Abpehl/CG6bkPxiaTtM5
qiURhDyhTETmwSHursKDiAU5k/IYpSvxPk12fp+aa0W98QDETev6EravSsVneebn
kWC1uI4Zh4FfZXjIEAXeDO5SK/vc8fVct548289m/KuJXt2gfFjJIDJyoHJ+Mk1+
ZesUI2whTqHUkLSeUqk78J0mj5eRJXGiSqto/2zAB+JCsRZqAQh0j/g2rRDTqqda
afYsiYkd85MuMNQflSHIWG0FKyW36Qb0yq/H0ndSV15kFTMqs0SYQRJGifHWNZu9
gSBpsa6pxrkxaLyD9i2PmkKOt842GEnGmiFMcqHWX24kMTh3Rzyxvgi/yQZ0sK10
gQk6LDkBgFnkHhCdhQDo5DqSTTCRhKHNuMgCbQTc0J+101QXHOFSjcxEJBtI8nje
+JoLcZq/DRcx3uDliJUvdBRtQMMACP7lEdZiQiI9KSdrmzS3MVBut5UDZYA2Ght9
+2hH+XNfYNkmevIfUg82xuZs6v7L7czJw1FuKNwjrud6b6D3qyu6fqzhXOqGP3Lr
e3wKnhym+z/pHbk1A1GSCS1swUTX+WGImxUteZhlXZjQyJsO0ikx07iwOGHxdTtF
+sep+mbfWqQmzD7XXFnstqDGszBQ6AhViXYw0tCxLJIevJCZJkqwhccHYaLj1IvX
JESFGD/+twqygiOxvAn/g/n85YhEKgQojrvOqpwsn0K3rjN/nySPoi/8iYfHxikf
jYd7R705RlwDKIVZ/gls32jnB6ZxmMVj3XCTO8j+APMs1D0nubnAwOlEMZx5fltG
eiLOlY68YjaaQ7XEvsiyCmnN/iCh89I4SWrVkpS/LFTVg3GP3EP5jzrOcwTQIkz4
PByV0iKkt4rTsPVf+biUmLpIERSE1biLfQ8M+8gngmu0HWXff/NGLXStpzQlxfsa
Vh5F+MEJ2nu6HZFaxa6XIEaYH0hjpPDbu8bGdc2zL4Cd+Lvba8w+1n5d95LSAxSf
zBqBVCjg8eS2VUI6cY3jFu3CgFKzqFbKeE/TGhUHmgIst9MPtRGC/qElL5HOnivR
InIOxiziuzWKauvlIvOz+f8bABAAZ5eThLE3ugV37uxpsbotWZ8A0V/b0Pa+ePza
yuHdkmnqb84CPaTySLzfnCO1UTrbNySOGBlJSgqxN2YtHkMUhVrKcwOBKuS6aY0Q
Hfb6nV0E4lFMMVuyA7+pskcaJz6a/tE8KICOYYQYDMy9u8xLYFscGJ65jbhWfq+r
KviG3gn9/IVpqowfgCn0TXcRdlIjohvtAQBS2e0ctSF4U6PB2m6IRGDNT9Qtvgev
cwvFj5Th2XL7LL2yKIN27Kjwzi+UkdSy95EKuLGZZ9tls/FvHbJIIyC4wvS2W1mc
QzUHB7gKs68hIB4F44Us4l6N18mbikdI7ral9WQiaMtgr/FNd24ez9Qrf2n6TUiK
m1UJM7VN0fvG4Jrh6R4xMnNVha6eaNvyB/GaSW/IYPGHhoC4VBiuoQ5+tnS1Vf+r
yLkNrugOMJzhk6FF4DAuFqDmR0EUOF97qt7t/YRxCphUGrvNVb6DuZXZL+7ucKVV
wKg5holOoGhs8SICZgZGyWl+wD6plgnWElKXB7muLncabna8gdNM9H+gbndEjT1K
s6DGEKqwQ14z+3A7+OkVHPZ6WDgqEdh1w6RWyTz0DaRGkxdtCOKcKCrpT8L62E2A
DxN1ie6UxBIr/t6ooNrWg1AQA4UenBDaN3u1Hs0ucTAAZhy/QcBGEk4lyVhk+634
/EaYiGy/S1yvlcxmSMa6PlRa9FyUY7UPzoFEFDtYyfC2oxGqOwg4chIiVy8LL7N0
34M86+WbEemxoqfi0n8O8PDBvp+ofDM5i7AfuqOF9/4m19vywejQOmA3qj3c5P/+
J9yd5aGwwR/WOyL03gjfQvKtAuP1UCl8i/wx66NHS/bPEmImq6kWuZWZ3cINYzJN
CPUFWrZ4B5HApusRcxVeeLLrscQQB++fFHVy/CX21qPfLRcsjFhahVj0aD4DCfr3
PqAuLgqd/FopAUkysL980UzNqDmQ/efz5iBt1Y6MDwzuzARcub4H6gbxPnNsCV61
3IDZ03Gd9TkyMWy6xE30QU63akCaW/uEZ3IXvvrRUiXIHtlyGFYvZ+2lVt4yYs2Z
GuCPyYMTiG08CiMT9lXLCaH/XW4FfrUznC4Rlbexu1hNk+SjieSFITKRNadw3D3Z
gXB+deiycuq39HGOfILSc+Jkv3pCkgpX27nfyGCD8/WYDJlAQw8jbojNY/IdGUmB
GACsy0TjTDU57xAcN5JyFn1jGflyH0xMXl6mmKQJ7a9HTfndsrREn2miFv5N6aIo
W2fZvpVqWEOAb/tKJhOao01wMZZF4nwfWNsjYkHUnwUQhIn9gfWPB95xgZpR7RAU
t7Jpy51NZaUVTDNAMJcH8QwIcfFjObqMsZLBZozCGAPwD/SWwJdmRPOsIM6aUQvu
H+aNbBKQD+5bgs//9tCNj9QtUCSllwbv74+M0y51H/0XVNWA2dUZZzMmx1XFubMj
9kRJvl9CsmC701Q2OkcvsgxhDbFHDkPfG88GNm3CCcdjwVWvEe9l1mHbQedMVIFF
I0f2Y/Y8mfg9tCd83rrOx14cJ1PrZbd8UpjtiEWx/ml0zwd8SlmKmlPKCEKE5/JO
Sw1nTH+I8StAZSCnKBGKJ3kFW7Nr0wdvaNvrN/B7pyg2PK+raGA5Np+LyrEn1NyM
z/O4D74xPXgSiLrN6Em5uPJxq9ppaDzD6zBsYKwmDczv5zyYraXlXDiELNDXYrSZ
PlEXZKTRvk8bGoEZrvxmWymNadUDMmhsbdWpofOJHwbRxtFHeo0eShmZ/bU0suqm
qmWUEXDN3e/M1J+JN4Uy8PN6HLVBkftCHi5rCno5zSruKCUlHpAjoOPznQaZHhbq
RqXhHJBHWJjP7J/4fomRYmMu/J5RDUDt/xkiE7ZMDuNDdFwwtLK66M7gz6PKk16a
qimqX8BH8EeOyL21zl1SLDGFoA+676zjZ5um3tdcTu2r54XM9z8sluKGZ0WDdPu4
5kZDUUOijTHmIC/jShGrAbA0b7baFRKq8XnoK7O4K/wKBTBwPhRmj9uZElen6SaZ
PwN8vq1Q4TKZu6UBYCmBg2TA1PLB8LiD2if5vUQDwDDxdmsrvQysDiAWy6z4wHSa
kcb6qK5PXg3QdSzZIxiTfoIvozZk8d/fAbjS9MlZ8EK+UCbw4GLIbd7G3O7KoNka
pDHwg//29baAbx0pIhTYtw5WLmPtsNt+UiUsjD2ofrPxwhpbij0XADzeWMsF1K8r
0SDBoLqQbpXHW1B2KRYtt1P2J+iQSjf5VAugDwhgCf11p+sNdqxU6/X/luo7ja27
j5eI4I+peDnkn8uQLsVaaGk3BOIn25Zm3nD4WQuChE3522+9Fze/L0y62/EnxAyM
Lv5Dbi/LO5Fz+DcLyNoVNcjEuZ7CmafrNxcTgtnleBLiHfETdYVy+PurwWRLgvvP
w8t3Wz7xxuBWy8P+QOgAAdUJ9krpylgKZBb5ltdn3aFnTexmsu6N9T/K0GD/3Pmf
M3XfvxODMv5UprWjP92H1zmVuLjxcoo88SKpo804rhpD+2SzKFdy/cFHdU8+x8ny
73F11clcqmtszrGfXm2yF01qTAfjmxBriEhZhjYPUgHak0z5DmFH0VPTTvmUP4p1
SNaNewWHtknGkhcSLx3pvyPl80lHJXSwhGP/fPnS9UqYRY9oeSkz/yeJGu/aZ2T4
YurZQOxN/t+61hcBwkg+IdBM7IzLCBxKjHvew2q08KnKdn5DTOnvWMjUFNZtftg/
quIzsfGpgKKBk2VjWxBvf7pjUoWa180g3/uhDXgW36vL/PwX35q0f6F0n9FzL58K
j7fsJx8uGTy1eJk216zt+zdcn/uLzXmfrwt5wOvcv01vDBNuFLwAVAM8KcPdtYi+
6tU8yRKvLVAEWXMR4C2H9C9VbRXOVWInBLeOjCAs9wdLa0TmFoeD8uqeDb5tzodO
c3A2W783N1w2mAWsXkL+4FmI9kUtrTegu9YV5WGGWF+bo0J61Ck5CQYfM+mQHrT/
64gjDIQ2J6QZ0dauix3e74DsS2QZzBnpPtqh26DET4cqSz+HM1/9XqGPuyEwJ6U8
RMID2yP9M0SKuvkeYskV1Z2Z+dEi4T26JfR4sfBLbFn4RrWMPbHNkizWj2FvFVFK
ZfGkVC3auy47KaK+YClHs39LH2Jz9hRvqpf8S/1/Dqqrk+Nd9ZM8BCTqEkrMPj4H
sSpMQamqp5fkHN+fEAWDqo68yb+oOfxArcAZhGNGtHSk4iIeNSBdtLAou85rG3/K
/wR7IZz2BJg1XXALLTGoW1bJ2QaPxcrLuztjyb+ZPFlhEWZcuTN72cuJ0Q1MwNtu
9X1W9w30Joie8rKP5ydUcLJ05Xep9kdXMeed4BGxeaaR8e/ifq6Iu4Y8IdsVwPE1
037f9YiPzoVPCy1afgqmzQUCoL4gwdS67C1/TWEIIsNvJIJ/9bLWyjYt85GX23VP
7froCgm3RixZML/dUk4hnmokcKCNtXJjO4iZw+WJD8at0FoSf4WPLnMpDDQ8HFr9
AsEYRLw71kpaVxP00cyodILH/NAPao6cOll4ubzHZiQHW2//syuJDS0qB5cSodWy
L0q+IJbLb4oftL9K3NoeQ8Zuje86/u/sgQ43/hCwlihn5f3pxPVCLRdK//pTmCHu
E46mxYiBmh/d0tSCAr+S5YnDm3ssq/AbDUWfIFR7WmKOI7KwprLCM062h3GMrrFR
kzYlQkIF4+1wlVMq2E2tTrrWx5hsuiYC5Au6nFJqvdGm9NinNZ/+/QD+Aqo41UOW
bKsMR+4DhAWmqV5O5FjN7oENlfevCa0iZi7nX1EOyBuaHE4iKZF/ElRkc3YPr7SJ
nL6INH2BINiLaLwcudMVbodHCB1Dv6tHNVsbjh3bjCx0m7+1CjbpAIiIRg22p3jI
X7E2l0ctVQlY3wqYJth+/lj3RfUJFNbxZ5Aq62C0LCwWcX4OdRe5tft7WJOVZmtd
cDKUFZJ5RyJ+qr0IuYQDrswUQ7KCakELomAGa0zBT52lbV3iIQb+zPUSle1fUG3k
B9MOniUCoQxuBIZrjuAQngx7OfxBv4ksjaq82l7tBg4933Ie+PJYlsAoYhed6uDB
cO6BPQDsqJyCxWvqf1L6462Bn/oWRd4TM4pOEJXgcbk5KJwZXWWfLpcwD9Nhndtk
FqELTVrDxlp4b97xS688N03dQBA6C0g9C8nesNtTd68Q3AfAbwDWfBycOrBPW0C+
KlECYsu7NvyY2DkOi+1aSTbgCfM9ifpv24fbznL+7Tf+bGmeyLzjwtINMmp1bmkP
YddNX55zKTCc89RYXD6mxyNM//D2q9DpepiSOuc2D8DgaduQnYTpvKtktDdl1PtB
wtgMWn6B8/GKjngMtyUNDkYlAI2FQB/6Kz0QOE31wQ3IbhStHTWzXZtt5y5B1X3Q
xR7Pli3jdCTKEFBsJ9FRdKKWbgOtKx0HCdEClMuC138DJtHGw10Oh63IFY5yZaSj
MV32t5Fw/nq3XgvCWSrAO2nBQBcH27LGePjSNAIJr9c5gZNaaCEryqDuZJD0ga8z
Hq8HamG0nQyz6Fdrn1Gf8PQJYAruWDLRez6vg7b1QMDP6Flsp3zrI2EJkx9Gw4Jz
G4eZdgn26bf0hWgHh+NCqLvZU+Px/EMibaSIb2kme693SOMqGxqAWtyxKHs/XWTO
IcdisOzGqVC5dbKeY8pT5DamBaZwXGGtGBn/ZD+R+42txABhK6zL2Gq+VHG71uhb
Rn3pt8Zza3VD8EUm4d7lkwMLh9L7zqlffNQ9GredRMuo56a0C3C0BD4JRoHO7UBJ
/eHeHTkSaB4ydT22nZZjwa4gz1DdrQ3IAcDSyvCSElb44fF45/s5OrpP3Zknwz9v
QTS8UjpJnaoxx5S1OqU9KRxhORfcZJrlYjn11+4Vstwg65kRQ3eOPOFvJQsOvgq9
YGmOsUbjBehwfWWx6/jm2SZRYTAiqkvxs0AxTePF4kSjpU7v6zrI7i+b5TGONQkV
m/lBLgA/cxyKhDMSnG+XlFUf9xEqKavzwUuTA/W0oaAl1CwdsEAQnG7LVec4eIIO
5TQ4ecmTkrQ6up4QE5ielqZ5TydrzDxyfNxkKw9mFQ4EmNGGUkchy45gRAMVpsPb
Qddbn40GV8ONOMyY2bTdg3muYZZyfOluYpgVg/t0aGeVSsdI8Rvr+039ZN/E05LJ
6Iev+Sn3B0knHk98aKdq+TiVu/NRX/c/u/UQpRzxhSv/GawNB9YE2XiSQZ5ktLlr
ETyASO8bZHSJ+9E/SeTxSc+BV/xEKEYwlZ4YoYn11CnepMeVFmJ1myv0YlmbAjLS
unmVZ0+AnHv1UL0DDXcta/3HE+uMvVUDgvOzTMeicJj+UAWASRNauDm6Xyw1r0rv
T0bjpTFlyvj/t3FtdCewS2WrONFXNtMQolvzAA6TUtRsdR+FwwwTkF8rrp0tFMG5
LrC62kZDSr86lzUKFSPT6lKR52OfZHFfMzvZQD1r8T1WNifGQ1zUbw+ecptw3eWZ
y0Inln/IPl1P4anWvhI7fFM+/vpR6nsFNkDpO1L4BRJuyn8Brz4u2q5qm12UjiT4
IP35Gx0pD0eNGnlYzVOazPWBxalQz4Pj/7w8gCEHr0kpzl+hEd/5Qcx8kGaPKRM4
gfdHHUaTq6mIS3KfcKgQaf9ac02vbmDdM9m/3kpgqOQDAjReM1nwW9+cl3D3phoH
FLH5MLRkRLqVr4eUkl7MbZY4T5ZUHyRE7GkrxR5dQSc4jZtS+2fPD8VvD5A67UL3
F+jYEcq5npcD2nEXNCTRp3kOa4uwxokSRlzd6aOfR4xbFg4ST/O7Np6lVEPwhdrO
+q7cgn8ricmHib2DZE8HEbb8AS5iAHqsJzIgK1JPobVIcZh4d1Xh992wb+XzLQ/w
xrKPAGwx4z0lgA6pH8BfApaixbIJh27nNJm6MMgCq6ivamzHcJfDEDlOPZPldSaO
viRG1eI8N8nA094gU34n8sBLUsVgR2AiFJ4mAzYMgi1BSUT/c+FYqeWGJJ26L/cP
GXb1CYcJ+fY73t4tPRV0sjSa+Sggw8M0q/lP1VETyrBEVrtNy/ZW219mgEeV8Hpr
+WtBi0MBFJGdHSomyXnPrnF+kksGhDHJerTorW6vUsNDnVi8a7ISq2psuX1db3RL
18EsLmvAcT7frKAssHNDfFxax8TQoDPl8OBwp5FouPDstBm3Vmbvf297H5SNTtRz
cV37iwAj9slr+a699tII0z6run39WCn49pwvMYAWnE/DDEPzvQVM1xwQAASvEsEY
SuM4pc0tZ5R74HnkKMBhkKD7WXL6b3U4PuMGTS0Yt05HCYrDED4k1/mcumhrC2fG
Zon9J7yfues6WKPXfhzwPq2riJKO6XoN+PDib8lNTFDVZJREnjCCYEbySs2ihsE7
tdhyRgsMrOHA+jGEr5w3TeqKEVRk+fPuho/opCP6PHLs8Rocs5/tkzMxajq6uTIN
CmgOBbUo7pXkhbsjbpuHnXrdHtg+oZoSCl9J+83pmsDVwWonShYzq+FwqEFzseJk
EBqvOVAPQLE1J7D1lqiHL2ViNueHaGAtIMWmYEk9rJ7z+p8NN1Xp9xc4kbQp22Pv
XYmxfJF5V5R9Qe69MnAnaaTxqfyEXPRKbzJ0z957i9Jsvzrae4KNaTm9M9LJfanZ
e3VE1HfykJd8yRuA59IJvfbUO7qaVsds6SF+s8w3O2wamywzm/oRbZx8cJReREdI
vB/AoBmd+3oPxypcdGgza3Cr+BRzpBt9SlqLiVRR19VxNbOITOBMb1glOdyJR5iR
9bBA2cGstfXSXJ1TiNv3kjXvvfCQzOYSWEtwEQuzziFLfLhfVzlpzfSFcBIw5NPB
Si2RtAgoq/jBh0UVeKDRlz/zhMSFpDso7OG53gdqKUFOruSGBM2+QhQ+uW4sXqcj
5SXItiEZDxiMDDZuFr1bqSd+SdGWLi2OMLlJiutuzgPb8qbFTVWT4fDazGCs5M61
meXHi7jfOoX4mDzF9hvbVZ9UuuzlSlYRAjWCdCLI9rB1hqzY+Yfk8NtB596RoWkW
5/+aIQlccchAWAoIoiC1pTVVk373leuqKLBWxxPQLkCdSgga1I1K5fIV37OguUXQ
ZKFwq1yHMQxHqCMGgzFulBJY4cCI6XxIc+Ba2FjKzUg2XFtwm3RoFpUgXI/ykKtP
4sOcPqT4C16Srrv+VJRPxzDzfrRFgJTUZ+7CHODrY2xhPmgsWiDxU40N6PSV0EDb
6qNa90Ugp5J1W4KJRWU99+VsYqKANl6l59uWZ1TBycZY0+kGZ+q56WEBXKXJz7D0
M/7GIyMtP+YoFYhaVi3AUQcjmgE7b3sBMtuM0Du3+qAE3uQjOgmauGoGl3hrxRCY
LsuI1eQ5di+xdC9HC2amSluRXxhDXIV0sLHraL07Y9g9jDb3wreeQwDMCAYh/4GT
8i/pdQvJHalB89+HvNNdTyWnvdFpTgqNouue/Tsvwd/LsfAQfK/NEk/myhkyrDn5
KY+GOftriT7AxurTDrXNie9NbC0a9UAj55UptwJR2OqjCSn1Lq8nkboLREAk2PT/
sgCVSoTYh0kqET2FjmfZCAx0nmHMtQ/Ap9N6UbSGoxWvvc6LFK9aNViT9O6N3+xo
BS6n/LWLvaaM8/5qOBqDmfURf85N/zcV2PFpFDOzLQGz05bRD6Xg6Vi+D1nEChfP
456t0oFDioHt9VMCkmXBy+Bm/iLs50leglCdCU9aTGpQQP/I5SSG+XqKB+nTQ6KM
c2bXTFZvs4UT1typKnEfhL1Swad0dDnDiv/XsPRCuSp+r2A2Szj+NgcpIQon1Dtd
7bA7gtZfty+hIQcPAo+J+AOOtbNhsKKVEOQcHu5QH4lDXE7Xaja2Or68386RSJ+F
JVwvcOy4wO7SAgIu+VhyKYI/XGUkfwRBP5zXChJbQT/JucSldM9tb6Mxew4Z/4Gn
8Oh6Itcl5zr64hiqhmnm6Fd4V6Gwq9lcNP8Ly0IEfhUXdQo52YgHrBGU85II6bJ6
IpcA4MNW5VjAWIGvhACjh2UZCfD6lAX7BxKInfKNLB03U27hxmZ/2sdMAnHa9KAx
cTuo+bKfHaeeAvL1J/BhPfgVQDk31XUy6UcEhgUpD3baBHeKaIq6Rnj+LlKOd5Z1
/77oFdoLDz8N1NRU2rYvP7ybzun6e5OTANXpthlHQr0fIeD0fYVwlYtuJPMJ5SQy
WoLRjQdzQWGbcnGMhQu5pxPUGj7iATjXXDcwmk2/BZW1F/Zv5B0XGzqcvYcqh/9H
Y8108hapBj+/RbeWVw6UWKrCZNndZk0IKWfgsSvKDZKBK0JxkhZpm2S6fRBaYVgb
YCp8n/hHXvb6npumObAaYUi2Y/LyoqgwvABLceS0lY4vPR+dYwX/UROErLIGc2BR
8QlO7n0SyJyoUZDaWjvmNjaJ1C4RSCABXQe7LSruM2884cjEqanFwPiaPX6y3B0q
4bBgJR0O3P8vCZuoMRrWx7j9pgz533i91XMvV6qUn4z4bzSg33uonL5ouoq0mN/I
/QHQ0HlGScuvAw1VQffKSx5XVlPd8CD9LwcXPDTUFezU21CT7/TFQuTP71nNXG+Y
7T+d4QzLG8FHlhN2QGjXOPvVTtrLxp9zsi5Z29UqJGlDbIG0I88ynuEkxufE/+SA
Sjd5rsaS/zSVI7qU1A1ATmB/oKWPpYfpicj38WKz+21t3tCArWn1MRsaOURL2ptK
BTVKIoUnjDANMwjb4IPGt/AH1ju5zH6kRLGOc/rOgeZESTEwKJfiSXkey2rTZaRp
7K6yCP9+WSG/YY82s+CHlpR2heVPP+mQdlorJUlT9qjtuGsniy+to8snDajR7ghz
WHam9KZgt6meCk6ntgva4/m9IaEFTOg/ycttXARChy4h5zcqPXRNbBEuQP0NlSPt
52lOvkDWEMPxtG9B36CbJdwqPYG9LsgMz1EgiI5QxU9TaJl0dCJu4F304HQxAFM8
cnXFfTgY3EfoqLs1CuCJMOQllC8xTHbMciCbS6fRkwHLaYQ0ygeDthaKXB5QdJ15
oSCw5HawDaOVIP273p+3ljR/Xx/0f3A1o5/AVj5UULWfrFt9wNYoIQEtsAdenwCM
0dHePXSi9LTlKV1rHfQPfEYkYEOv929qa3VxPHxIjcgsbPQuCAXpShYjw6G4otxU
IbhJPY0L/QUmQdFObAXRyu/i6hLreV01lf4mFVyNBt+xjFl2in0luLa8EbrWPDKt
wMVxhw2JfwrGWZwfgNZuE310GobAIC/mKs85r6BmIqh2loqxaSUp64sXgEpEfANK
WugZZIZPsTCZFPwW/6FVn80HN/T8E8hOsift6Fr25+gZfGKuP9FeSJ6itZ58v5Zv
+VLaUnFGXco5JUAfX6eeJ/dTa6XUzQa58Pz+YBNAt5NUEzdOVdiZUKZVioNCc8FV
OfErz8HTeXRix0D2QoUAB0zxUwUV7L2sNXpE4R9YGJF82+KDrBWB7eA3gM5dFObh
2MIyZQf0AeWwI1XTHpRIPfs5+yWzE/io7Ojsm6I0AaVZXVW4o8Bnnr7sOtwE04nv
NluKZfXZU1g/LxHp2DnMb7MWYKjPCum095W+gwFVJdcBmY6dsey6hBtaNm68QCgY
Ldl28S51UI3092U4QMK/x8EDzffazbhlV4uFL7NBrNTf3i7KKnSnH04IL8LhCL5v
vVBRbnd1o8rFNkK84h9jRMbCdN2LelL8p+HH20wq6wTDeuRAw98cJH4uqNLkx/8h
S8NKacV+PkqpYLO6lubzIHrH1IT2YYFRELUQswsNNJa1YwjOGpdou9K8W+MZn3R6
633sX/KqKwG0gCe57e7mjcz8sO7BWDrbb5kSw2Yl8EWSQUJ6JmGnZAFPwfiyYUCD
w/kZ21QdPjZxpNGcE5jACHCdrCkJRrCZ+dl5IPr5yJ2F5AIL3UoCF6Vy9G+ZdXlc
8Emh2iuMDdxwEHH4ckTrY/jSWbjkBjhAn/nJfzvybMdj8BHradCOVsNLwZ7HzH5E
a5WOjpSbq6+lstIKF+yW7BCG8CdYlq0HMVizv7z3lxkcLFkCWtDEdjCatlvrZ+rp
yB/aKtjxRqMf6kcZ28vVq2duNn7coMNfViwd78Yl/YT7RIWzRIHdjzKmMx9CfH9b
8bKcszQLn6fPT7gPBMITdyVzbbsO9+jMjqzvv7bWCHH8nnLmgosCfixE4BQJZ6Y/
AzU5iIKEZYggrCKPlQI2ncDvCvK9OJ/HFeK2b/bzykshE4meXv3JWAzwYFVrPAfk
iQvXEcndjEFVF5a6Fqaa7K5kr3EXtnBzeBFwbVtenK3G1oR1wU4V+xWFYZNX1ZHt
EHi0jCzycMkkiLdnvuN+9wHoBm5GMqutUmqQhcoD/SlirNRESe2OhMVrqOBv7jte
KoIXTeM3+UStu4MHPepxMtL1n4HqHU9yn2XbggUHY7GOAqgNZefAJcl5Vq4qLHlA
faB3HnIvKHuuXFvHyzZSJTdKV2N9oB+Lhwu05qG4h2XpbhjCLUB4lGG0EXMge3Ng
N+uWO1kGyfD8sl6imGQRgy5fDGvLnU+4j+SekcJOvEpkKnZTYPh73awrlSXWKG5s
ik4u6+KuPmUO3ucHWIyyfjJ94nKibYNmZB02VNCKFyDYOsxmT/yihC/2JO/oSRr7
9iZuyKDNUS+WQQzCp2+SzlPyMOMF30AewcpiAsRqSEgaByS/Xl+S9Jrj/14E+W/1
S9+WxCR86OJD8xg3UEyrZaMuI/eaN4DFGTBvoWY0ms2iyPi5kk0QwGllBjQt6g3i
IrH98eXRKd/vsZ+lgNMowACT7JH0gedfO77vf+tbhtbo5Xmg57k+idQ3DnrjqFNx
wNmLE2YvM5vKb6Gbp0qJnBK/piwCgCyZ7YY7l1/rKUS1i5/5Za0czZisiIma2LXO
hnVViOevS60pBXNuWlmSS8KKCyBM4j7TWqOsf95T3LqVsFKM8vT24lA0RmCQK2ml
NFbabyDlevpwH42R/OrbfPtJo6qoRPd28KL+t3uKIPJo8bBqjoDq5NYDcldT7S7/
OL+48BU0SFhsff6+i8SDbOb2ktrtZZXsiGNyFFD/xfVLggQyswSPytViZzi1sSeT
kGSBEU/YaKvCCrH2v5dr7T7HJ+NyIH1gwMuvSWzpRzCbWU73qKQJ4//GmefJv1ZZ
O2QrqtUEx8AyZhdxxb04rO+kU/ijFSjGofCl948gA+ocpsH/ipSVqKxi9BZeFlHt
CtPE9tVhWMwzDPpfHy5ZrqmWwE2zu090NQPhruNU9hw2476FiEkl28yy4x8PaSN0
sADtAy5adx7bBMJ1Dlu6Q+WPXvZl9ZeTtqTOfVNKL7l0fihz4F3oPQ7HmddVE3uv
2VkzrXsItN8/eANvUgKXuwDVQRHXvUVKE2c4h3eZda/dUTsBXvk8EgMakhuRsO9w
03iq/f1mLk7fsjHYHIqQrwCDs+nvSItNj9fVLaeIHP5BMDk8wT9tDzQ5tGyNsuu5
1VePQOdlzX7NfcrypAiNEqlk5KHxk+AvWjUE6ByynsgGq0UTEVvXiV4lX0vRqD7Z
O75HbaaUUDvxZXzsB2SHwdiuBMcK/CiJARouBDEbwIALNl7uvfAfKsjdPIQu1qu6
q1BJ/OXruoMrCKcRMh2cuWdwKRQ1za2JR3ZBZs7OCX35FHcqCd0LHUGGbeKybA09
icaG3c+luq+T5/I8wQ7ZQz+wodPMpZKFvVMRCZD+oVe/noQzuz8/eK+Uu38zd5Uj
jGTp0UAGlkAZ3pptgOyeM59+73+uZFQ7djymubWPxyYYEWxlAMvSuyUBr4QcJ/SV
24G8FlJfpCWZCvpxuvQdzUMxHZTbNqxPX8gqxjbgViChTv8BDsROelbxniM5D+7C
8bUmCiRnYO8xYpokz49zoUIX8gbUBGraida5Y3pzh3FkSCLL0T78x2bZXemlDzgq
C2bqnJVqN6+dD8Jar/KwmSZQanVZFvV7dVen1wKzjI1xWLuS6BDOzv/6vAF992is
9bGe3L+tozJYI0Er+Vwb4JEQV+Y+u9ISA0LiMhwZT0K7/Qfu6+ehhwY8ym/yMISW
Y/vhu6cATRCEzHWcVOhybI24OYjssWfF16BN/JBh8jyIHBtcLujAKbqPadAjJStQ
Rg4JbYV5DouHFjC0wL71dh0iTTiUireySJ6yiCenMeW7gPce8CdoQDIiRpRq9ITE
KHL2SIYvTAHccOEP0as+ZTiEAmH2WAuX/X+iOoF0tvGhNmNzUb3wrh81VYTa8m2n
nN/wm8+v/dG4VnNcMDEKWrkUnTQO+wnSWaFVsUw32k8DIUMJikxyAbz9tHC5LvrD
u23FLUnwJ9qOLGMh16TKyuZiDe44CTMkXodmg/3dqN713mHDiQzrm+nyWE6CBMdc
PgKxLKhgvq21drqDK6wNBkVbjM56iEbk3UUNjNqcqw3wVxm/KUejU//1/SELfn7Y
b44SDQFUWNHD0Uyo0Wi7CsPYzEiF0YMYwsn3CME2XQOQzPYBDXtNw0TiP7qMPerM
kqMpHe/PcEZyHB2MUOvZGXgJdvRwZaQLZlnOWfzM9u9ZHyPdURvGHkmw0SiIQgVx
eoA2w9H8APfIGHEsqmD32nf41X//FF3WaZycr5Q7bA7a4//Ytf08VDgUFM+puFVx
0EKp/ONR/sHI9SCJyJcVU84gLXggCEsJqwOqGoejv3l5uMrac8HaJ3iHhf1IpLFo
DM4UnEN253nSJmwoEF+2CzPHLwEiS05h2cgw2botZuVcg4cPYo8wdSOJRtc8ecCr
HitdhDl2Qkb/+rhWijnQmHPrxUFGqlvMwxjf10YDsrYI0o+i4N2v+xkh3oVi10dR
6lsjQ06dlR0Y3GsOBtZbYp1n5U8r0bD+rp7rqRRc0zZ7Um8WwGCjxX31AHn+7sqM
um5BIen9TL3k/EvHwMcNDIQ7UduAut9k5psvbKNuhyFhsqxCwkH1HR505xl9JX3b
6pOzHk+WbhQfW+Gck8iHQODjwZ/qqvtFRXgEsYQJEpT6Xub98Sk1jZ6t6eQ4BwwK
a5LXwmVOYDerHYDYjICn/TT2sgFWwCE5rVvM8w0dSwJwIpHQsgTc156mNxmj6Jwk
izhWtKhqgYwtaRMmazl/7VxWRVelfG2P6+UK2klch/lZa1XD+49Y8Xplqcs3EyUZ
SntcBYo1TxNlmMpYsU4S23L7KQZSwBgy/gyAnDQEOiKTpRIUPdpmhfYqBNC2Y5BN
4IvlXUkxjH7Vu0ZDkG2XOowsXb1cGCbwmx+HRWv26AaRj9qCy46VhaaZQx9/puBN
XLcMs2zklrAFcoKKeWSapAM1ez0QNVdJL5NkV7/r3LmdcC9ZelqeTAPL5ju8fs3C
vS7diu2i0a2iv2yBVyPmf7t7Oub8M3Db10baw+VgUZUliWgEYfOs67eEgmL0w1qL
5QFwTcAZsA2uMOIAGlkyDb9po09mQXuqyGcmg+hY36FTqgZVyNQhjsR7wP9rmRP3
VQaR4edambPjUUqiAzK4SvUKkMRnqDqJVJb3k1OLAkmmp3v/58wrLTJZJONN13lL
/toUsRGFeXXdQiY4eQs9PgBSXxIZ1mg2iLoamKmaSJq0wNK+Zeg5/cCpyRc/dIhr
csbt/6s4anxlMIuMn9gqIWxaWAFUKrMbqEa0LM9zsDo3zsZaSLJqBP4jZZMh+AbU
JXsHgI42SZvD04bMp5j8mVrT44/X5L3MZnNiT/0xifHTDyYenPCM8h2cFZKl4Olg
a5dv0EB+bjO0SkHiT90GvBj9ZwIXhOXKrFSig9ygx10TiwPtj1aN4sk7HYl+BcBi
uq2G/k37hiFjWghkYkEdcWRcd3R+fvGGTCecEhhUGl+fik66M7UzVKqtOvYakbob
yKd6Iz4P7O0OqS5+wKk6zqYHrNSNEQcHewB+VZai0i2PARTPqchdZOWJbWp8p3QC
j5kjWLi0RSXNO01C4VTGCRy1ajXHxlzkFlLLmpU+1d+YPdHKpl7MRfNwkJSQkx2o
R/YdPZj+nrG1iiemjsYvFHnArdLL+3jsutXPiIlpvvcsvueIvRzShwmI2ui3QTyy
aZUPPnf0GqnVnz50bhq0x9VWJEg9LGBdRO2bezVWb1lEKW793QEAucPj0TH2vQSD
rYHsbdYa3M0sV9BcOOIhvaQ3AbtdhFdw6qdpRhE65Zfci+CUBu3HoZC/T8x4/9sN
x6AJUHMnDStcwBR0+B68kwwASVjdaxqLThV2PgYmqyEe7QuEhYtnGJxe5Cl7W+it
DgkcDeMgoosBLCs2z5z7vaojPUdfTM4r+6w/r5VGkIqfVtoiuar72cPacavJssim
79mclco1SbugkgokB+6AzV4tBCvGfjfAj6PSXPL+SX4pBPO9te4I3ndb32Uz9x+5
gHU/J1tCns8Ajwdpru8VqUQi+u5WRX4vY3sQ54hurEslloNgCpC7gNDCNnmQr0qO
/ga5Nlv5O2OSmlMCIlVnw47XdffmIMyg9ruLWH2ZEV6bUxyrqhFfln21suf8Fvxz
DJmcaGiAsek+9AwcUT+aKU+eOUWzY9lAVvK4sOMhCM1oXrDa4oG1XgqmcZDNnehV
vfHz8I6Yg0GWE1FUIt3gKFGdFtkdVQmHjUBMe/r/hFX1Kd5kPXQ04pyZvj/6zgd7
pSu7L8qRS3URmeux8tCfDvXZNflvy3hiVkqXkSlVgLAfm4YlMRbJwQbtukYvBrn4
MwfirH550sTXYIgfmicpw+a1BNkFfsj81XjVPbzSIHWWNW9KCj5n4z634vgyAz9y
LTFidXqsP/eqGfUSCGBQB2RGs1vch9alZoReBqw1V2fATAwFNXRk9x7SLLqFNYI9
lq/w6pFL4o0Uav+KOBZWxyT//OBBHxi3vojRtG56RDEEGrsusd70LiqOw2Tf79XX
nIoCG9Dg6pA7Wwtiv03n4+BoImzGf6+0R33EqjlBZu15IZYfDKirCPnSjZm4ikWc
1jSwahBLtJPlMY3Kx5PCkI7hzs/lAnkMkpWOFPI2ACtsRYb6LEg1lsMPmsUlywvr
+a06ORO2ZOsZl5k5OLcoB1Fo7HuXoIXahOv3ItVppyk6vGzlbmiFmplcDhg81q/v
C8d6g9quevjkz/duXh3C6a2C67aouqRoaDwLczMHMD52z+aHeYbrkzdSThl5DzP0
mbFCXv2NYv6gzoIiYeP54t8JXcu/5Hl5tFo3sXqYduCs7Sgg6U5z9Wvq88k2kIqO
Qe4CgpsRkTTm5gry/i5s8kmR/ky3b4Tq+hDTnflI5sPRRsAsk6wpEqdT7xhx2tD+
NGYC3KXK3va4iph7vqmaDwr++nTR2Sus5NhYKfyznWWcy24jaxoaRLK8OLCZuZ/j
/V7/Co+iSJf6L5Cn+ARCus4WUrlzs3jNpByZafbGAc+rGLEWr96Kk89CvzHw4y39
z3ceXvqtzCUPsgKUFh/GJ299Br5oiEGMSCvfoWxMu3XQiwNMZOaCh7TZgX6kB9n2
g/dwRu9lw2jR9IPckprMNaNj81SQw9h6lER+CUUvHB9TUBGai/Uwz+F01SZpKEV0
cPB4lubYly+18aVbLSRlSiPN73DzFkoMGLl01zLhlDkSS0uD5f6z0jcvJslyRLwQ
FEhO2VaDFYBXa45PI+zkLvzVjrMKwieSJ1tjutxGV+gUYjX3LHFeZtKw1AOchspd
79YtuT8Nw61pHxNNzp//FDUorXwE5JHE+n5Tp/SdkgYu5wcYMIiOf+ij+I/fMkPt
mYBlj3G8LFXG0ZHo7dftiBgeebJcO+X81HpPu41YRjLTZG2n07GNHZnDQZzt/h0T
y31rKix79NMDgdQjw1dQaJevnSbWlnWsakaCS22ygWAhi/BoNcb57iOEK0sd/OZA
dvhLCHLyGEDxVWeZY+fUOgooIwg0isP4PUO+J9Xtr6takrm53ILh6fsIiQsCszvc
9BgEDURrBonzXe3IM87LglUw6j6EcW7l/C4ikxcfXrikVeYQsC8BHCS74v7iTKKQ
/3nGvckn6l0cCcOwPW4qM4DdxLix7+PK4qNeEjC9WQTuhmyTClWp7MVxIKiHa+Hi
rAm66nLRS/jF1kck0yi7GGtCxR7+jTFPdQH3bxNMQPP2nz1A2I7T9gHe3mlpy/Bp
oo/G2+mTPRNYwH5YbJuCDeEAs0iPaZ7/+x6w5K050VsgBbHISeKEnp4bP+u1Sdnd
BZJ/GvBbqIEpwy14ekeoeu4Frlgy2POfBe7JtYx0GUcdZNWL0ZsB8OFYfEMGgFjx
Je/1TaIMzzxi3lV4K1NoenrwO9qrD8DjFpg4HLgR03nogw7kCsGScG89v2tEh9Sh
5XF8V+GDYo0lCNhEznRbYhg9wW+IKgBUGzBFv6P6RwN+Bs+LE7MB0iocwpPWj9v4
lfckBnoBmRsM5O30F7AoayL5eRwaN3QKEsMmRXRrOwFH5EwdbOREae1dL5u5g1j9
wmRXjVJP/YmFS6yM8mUeqTnBtv06L2WJEs63o2lfbL8YKFACy5oj+Hjyx9/QcsID
scA0R73KCMSdjtSoigFd+niqrDWbptEVOBYA6i/cRWB6/IlQzTKhsqZZp/xqgB6r
n8/Hs0QiG2KizRVEtbsMaI2/SCeg9VQPBf2g3BAiqmtFf5KhGWhoPXV4GT+/g1SG
7OrbEEOijBY0JohIPcdyB9sl0vJNvIraRe0+4deyWADtJ71skhDQHXUd04ZktX5a
3mFiFXPoRGL4puWyK90NHuYBUI+AHlG5N88qVLt2391uzqoI2DVOC+jw6fMdY4hY
hgcbCxVOv9ub/UaNt023Kz9dq+SqLKXJgXt2ZjdJeFaIJL3Km7LHDQnx6T1l/88S
aKXgLTmmfSa0VjMX2kO4xO67yP+GXIxpRn5pNYGTYqqhku0Qdvq6ovrHmcZ1ppV9
Q1IKCkeEyI2FxSNOa/8TgSmZJOYzSe/wZHUDiN0Wn8//WNDlaYOZU6Cx5In/+QJ1
T01bYvrs/cz0sxjGSRnGjTJv2dqQ/tPtgt3DG8x+cUMoLd7bDQyNHCDWB6ipOhAj
4hR0P2RqxrnjIFrtfIKUc/pTRO30JQfF3i9NmmFHsoDi24N0kfQ62kXCUY7nXPtO
48aHTbomPoA2FokD+3xt5CdUK0x37kaOBWOMzb1K6iHDvBQV0cDWsGsMTomLjCpe
ZeMEhVrB2pmZ4XbHtlpAR1aZLr258bEPL2RE4UYUz4U++h0Q7Y+sfpMlP4lB/aD0
uIDzFAf2BiCCxi8lpgmjzfaQkMirU8/UKw3LU/39LmaseA1l4BkD/0dqQjhCVXda
5Mp9SsgoChQln/mqGaYy2QInL72vJZKOa7r/2G1kjbwZr66lXs06bJUD3z68LZX5
CRHY78neXvJ3Sf7kLWWvVo4IpMHKZaeqPi8nroodKHF96A/VH9EzKR7SXk9K6+YL
sIkntNpXJgiNd6L/yZenTtQ/25QZA1nwD2GbQGVDtKAsQRe0lwByc7h3OudRMrUA
TcGUcG4w8Ci0kGlPpsaorlU4px4orJySPxxuG9puBgP9VgkANpHvak8gLQvSABmI
+U6HoIF2BM+4WcgSU2xsLPXcsMLkcMaeQPmE8iX6J5i5nBYK4U9HBnqW92/IxZ/Y
BPpaTItMCL9L7F7z+PNOvMVq189Gri4Pv/a1yGgItlQK34CcSC1qcwXD3fntJS5o
bMhy/oLZgybipt3tXCrItEpos2j+Vq8z+9nH9Ld9raJPicK2D0X35TniV19uUOWE
ucstiL/YyiNLy8ptybTolmcnL5YjOcAq+jmaJpgQ72t2WFUqpBvzb7tT+FolHIf4
zuCVW6m9Tq2Dm9X3kmz2Bk5H8yLp/rWxNXBX8l3vSHBzsw5KrXt0Ysx3B+v0EPJi
FlVD8AOOA+kdVIHAMq9dcLrJoGaDsOy3cpCH77PRRhbcjy9HxJthZsX9RW669d23
+EYDykGp0WtBIBCbuEYGogtTZmKivWN3uDbzQ+D7LWVEgwBqTws+GWAREb1GSx/1
VQzZPIdN/fx2UYf1lHoQR46ccEe3ecSiyaYQ1BgWdvyXsjYHyQzmNOcQYf9WCj03
ElUbjLCvw5W13uKZzUKypu2T2pkc734HWW9y7lb9bqtPLJoL2le/2+YHvxGjbHft
+kB/JWL9QpCvkwCPgsSlQjfRO2FolhVwnGoixrTyJGoXKTAHQifPJVFe9U5L8mmT
Y1xmxGYzOfAAoo8rFhXdgiyaipHamdkb+KhXL7ZaJfRMySH8M0VVaVgyLDZDOBEw
taPemzikaoxTfLA1rC04C6yQapCT85CKj7XCwvvu9MT3uiXA2JEWptPBXRhQPTGJ
7XVdDy3kuJ5ByymMLb+WloaCoK+D6Nz/jqMqLogadiWqI8GwMHuHnlNXa/PJ8c9S
B9gitHRiHix4F+J0Sj93TUH2Qb+JW7/J/s9KS1eqD+apyyx9FsG2afEiaQiUcKHt
ua99glBmT5CXZ4/msbuYs75SebD67k0g4LAPP0dlRjx3ulYf+FWlFdHvN77jHAR3
M2VZH3iCuID4QRV+zRDJrGAW5ITgG3nnXHrtR++kZXdWSZmlELSwP59WgiUeLwhq
HfXW8RpkrIH4Et5CQcKstFRIthaF7u5w2+cI0KNp+5AXmk7rdBTZNkUFCkE2m8Mz
qG5HP/7xyPXWUZFyzypJoyL1qD/bKcpktpbOprSAl4F9E/KZRILMJ+ydOqfB5hfq
WWYAdgaUsKCtZRTZFn54rd8Hl2VYuv60O/WE58tnEiTorvXjHyajoVY93rgYjf/n
VZmMJUfCjkUo3EaIE6MqJ1Bx6tQxa5FyK9g2b8nDUkxfJAN5uBPee3yPNEzO58pq
zK66OMTsF+RpS4UOUqymFw+7QD2vLunvHo4MvnLghLsCw8OXuYykVel+u/72OPQI
Jh+TtKIJDy6u5Ms9euOBMWBus6w2UkIcAcdPm0JmHUe/GRsyjXKb+ZD413FfOKA8
hObC3MnFPF3QeJ0N7o+YI/A2mx6+6kUEZ/pv5nW7g4MOoLLzLs9DwX9ZiitTcop+
Z+jCeP/x/3gvgbI0O6xDQpoub8p8GrhKjgXlA9dTUlb9CkpdcAVq1p16ZkckIVk7
IOpZPnOl7pvq11OSUhKT5BtBsGAI/Muo/znk0cLaqyS0wbHA5BK5Dg7K839hun9d
0xWwMJH73l8jx9auYnmuax5s9+XvHVH4/GWT9oyRObvhFqKlQNsAtaczFXPK5raS
LTFbogi/E0AyYkF0veVfKaWMxmIc0RR4uoEdDykmCoZ3b03V9sKfw5GJ8sUwRGGt
G6ljhCLzXFLTKnZaQMamovKERW9Hn6wsLruAyfMekxXrOnLDxrdgkH1+vRDqW88d
TM6DT3WHxOUTAxQ152Bd6NDFf8wdKZSOt16plxUnLFO4NIYjxMOPMwW1t+XeCOn7
m//ioaJ0EObVDKz/Rbk8MFVsIFbmLvLb07gAnS5W+8V7iTQzeP34kma4F7Z/pqVF
fInDXwVX4KF9T8xMlko14JKSfN5gr3qgQyDypXunoKmTRwRMUP+8wB03SlHosNVj
64dv/hxBUVvDBpvx5xlqofrvr9qAkT2NynOfPASMcEYNCFvN0naM9uGBfHvFZJV3
cTBffhAMVWgbeWKrvl7R22legWOyKe3FDpu1Eyjdt6OTQIoFHriQIWn52avLZn3Y
FYkA67ebyVeRv7U7ZNYblI6mSK1rDiZ/BWbgoNRO/GOsewvZ/G1viTpLUBr1WFF9
IRUwFFVTUUT1gDcFJ2NgxMKYaFcNByPM5bIAe6yrxnquoCEFaGpYah8ixH2SdySa
mRSqoqrP7jJd0T5iibvLbgAdUJlKEz5PruhbfcEbm0Sy3qyFHGB8LLVuf4nNrMdB
7LlID5rNeFYeZ0J6hNLEJDI66/214kk4yXXPUIVSdh8cxkpoxKi+CmSxXijLYak5
aMHFidven60KH+vtbWrX6w43OQ64ggy9Qi1jQyqflt7npS1Mf4nooTRMtRyrw5YD
2/0T2VvNiVhE05rB7RS3zyz4zBHjO3tJJm6Jl7klvXoOmT75FrazZZLsl6/0YHXK
tsYwxM6CFTUY6CgV8JV/AEEu4MULkx8UotiBjTQeB1iO45iPNPpEy8Uu5ekK3Dan
xNL4Awcj6Y1Wwh9GKK3wH7WXZmNQnwcZp7Uu/xZ7AXGCfozPSgx2izI0EaTLnnul
JKriaxuv1c23z/8HmK+vqis4kFWWzaPO6qG1BFXlwns4ZnK/dbl6Go7Tb16AXop5
X1iFz5MOcdC6UvL2GfPn3SpwpWHOedvSsKLg4QPdG8aamCxdHugsfVZxa/hy+UtW
suSuBYQ57h6lGNzYFyzBjFNGpzUf7C00zKvvT3wF9CW29SKQ+JAt/K+G2AAZWTad
oQGt9/LqODawr0A24XNlrQDvjuAR5lqiE0z1ClttCdFWe2PR0kyp/zlXUB9oMIjS
AAv0dGeDbb+mK9GrXhg9KuRGLvHERGHgHg2Pqk9NwzJEHI06ImqS4FHdZf5iPFzq
PCcerr4ghNHdvPt7oE035gRxfqfSNhWYEKTyQly6fwaTdSMg20r9ORhoFR3aIjc3
ukg8KrhAeVVJxvtrRv1clouX1EtFRIH9YWiCeHMSFeGBFHRBzIqbWbT6cT37fhYU
jEShRcAiLnTUhWHKXaOMVOUGY4K41eIPqxIowTVP4pKXKxfQedIFYu/lJriRP85A
JlYjq/PQ76l5vWHwVOeXL7IKVu3xEerZ3Bpr8HYCu6X+2HyxAZd4Kcah9wbDv3zT
LGqMAIf1raMED5Itnw7VBgN+yV3f9m0lhp9ja3DDHh2cK/1bWtVNBD80Kk9bYI33
fNSK3Ik7wABny3+GnrJiBGOy8MgP+eNIzpXFS7Y6rIZV+92OATgSb8vdjwOa7fi0
vZqIm9dqZIej5mRKFs5IjXNYcerPegLV8KkewGLVf3qrWKn1ZFf/b3sl4mDaXD6p
NZSVNtlfYn5DxLBwmLdty/AuKxMqV4iTV+zNULS+A9e5NbpkiRVsIg7XwkTfKdnX
cRbGAcXN2eCyvuXnE3Rg9E/j1SOYUQwfJ5yMJEYdDpK1h8gylzvAJXTco0SHEF6z
zY664VgfEFehZ+DYjOqCYHD2tDfUYb7mLbgBrXD960F25As7MKI27PK33LYzWZgs
iFWr7TbEkK9zQ4t2FO4QayBf8CZhmKw4YlqoDm9rBQIhqdTqJHGAtnCLYBZCtUF2
0wsAMrPEsLXgAWr3NGxjR3UFk58ai5hRZFIZkkMlmR6NwfQZJhuolrZLgCnitl8U
LEb9jvdLzuhMGA9DMA4h2ldmF799QNvI1Z9qXbF/MCc8aVC660zmtuPc40ZjRc6J
nHDXfDXzRrCVT0zuutp4k1KlMk1/0dge4y3SekxG2G1hCX0C7ubm3Y0Wn5sr11Ct
MBRQnhfnc3z6sLjvkKStWwPeqCxP3JBCi689OSdC2owup7ceg+2ZNOTShEW5Jzjf
uY/0WsNNdsmEX2GIMSEFWDwwmU5WQdBGeJ89wZ1JTV6pM5Xr9MGr//+j/TJSj6GJ
RmBIk6+nLLnrmaXuQQpDIshnYKGazxXIPegJcNxEJhpZHcUyQJo1+z8XVfFH18q9
tuYegc27UVcwYKLGRldvHDz91iLk1HZ3pivCRsle1SjwmozePh+Qs3Cztx4jfjoi
Vd4Rm/EKTPO2Eeb6pvAg2/dWN83XceLYz2XoMdhOeRh6/LKUW4pmoyKpLtD51X5P
RBSwE0QP/ve/13EHn6jg3B2Y1LBhpcOC8pdepMngDUwA9y1KWMuOKaA/yxCp7BpT
6YEea8AeXE2f4tb6lF4gpYR4pw9gPvrecdsrdCBuApkq8yRZrRw4CzCxaQc6QycO
RsM95Devcq1aLho4BcBQ9PwZAF6SRAifT53y4CGxkn/gveYoMNQWdlilF/TstZP2
Uk3f+IkUPxXDHDHW8jFoxV7s0CtLDeDOHvoCxfOekDL5zIpntzZcXab0fv62DNT/
xscmd39UVk/oHi7iyRG2Uwdy48CQTt600ovRweIAsmXATPbkyED5AyhlEd3X79zU
lm16D5w8krniac+Mrb8hourvD/UydUwE/9OzD7HuOhKZXXNcm5gm1MQh3Cwxpq0/
f3ZiG1lDERQmasBEa2cSW6ds7VZIebZ5YCDWXWubGTgjpSy/oMeww9aCD0tmdrgU
QjFhZfkinsF/Y7MJnJfnM6Yix2osKtVQEX5U8//vlqa8+9BhMwPjn1DCAheuzwbP
tkAFuKVmJ1ZXwUmFkb0eLFiu6Sfe6KazYgmtv29YV558GT/kLBP4Bd6HjtVI956F
gLqqQnSF4cWkXkjteYe94fvwC9UDoKbYN4I7PF3ParuMhwng/ebbp1MAEErkuiwp
H1VcvbAEClq4f0PU5PS+Ilcke2SfYZchhJJ5dawQ1SFKj3l9qvVJV6VBNW42vg75
7h+WeQCxilgxcQbcLmExlXNRUQnu69MRMkmj3rj/DBoTehHGmfIM/yP+Cs5UxvaL
TpYlkkFtB4qWGqcVLZRrAtjUehnHH/Cnq7nf8zqLt45ej3FgU5CWe+ZHX9jDxGGr
5OxIdsKuhhP8nZt8kpZ5VLhffvXBbAYzJ2/5J/WOoBVCoTnOCPEeuZw48ZSEEOwJ
U+E1LW/TDbF1Sz42aSLPqhNiXHGNrlPF4z21M8QNHU2SW2w83C/4pt2hDQNi/fWC
r6Uf3+am1rlkeURdN6aKVmNQLcyVe5B+eJ73g+rEAAQx9Sxj3onPc4sUprcC0cty
C2DUz6a3wwsoaCXD3XiKLAs1wO0Ovv0DmuSINO/lzVyiXhOK8NhzKpFwEN0FG2J9
BMOzzYV+ZcKcaXf4B8/D9MyWSwADxI0TiJRRl5NITY84FySKRudkfXRsAGCLGLTZ
75gnRInYNf3H4WL9/2Do2bJonnTYd6ytzqK5NuhXyR6QaHTD427jD6+wjgftpolf
3fj7iI+GmVLQu7uxGOGucUZ0OdnjKAn6x18Y0lR8Wr07hYSIx5e6Ai5r58GlWqz1
Xc9LTJA9qQMWY9CN5KrS09fdV77IIRZU6V44QvBSoOggdaaHaOkBQaGXozHaAz2l
gA7mNkxFKQ50FK3O42CKHkMDkgaV9LtoybhkW3F9ISHUxAE0u1fUPkD3xD/XVk5z
Xf81OIQeo6FEVDiRqikUPOLFEftMc56+zTF9x/vJIIBoGLLE7zqJhXOWa+zWrDfj
tgLcerrkEul0AppzEk+akE5omHPx+sYytBWJ0UeCew7rbOcfzH8a8qnaS+cakL0D
HRVFUaE48/CiokPmZtAWyKemEPdPQBhm1TT5yYIu9vMS8a1RvsQ/eJLZJbDItoM5
yq6U0cWMCumCjkrobyK50qgKiEmlm85M4ai0czEQbV5KBvfhJ530K3PUQqLrSWwn
ezu/4U4tuF8V2Nhqpg5n4hpjUaXMg8kmPZY9zWP2CcyJ0s72+RFJ7CPXiLIWRc8T
O9sZZLlgw88fwRAtx/rdGOP0jfHdG7pllpy2cF4Zk1xGQYUpeW0xGAVqpf5izNmu
9TFwUva/vS+HLNfLWS0zg7YAyoFzoCYC9I5NoSy43s+mPq66oJGM/WbfjLSCWLXb
satCHLh5icO2xj8XuEN/jj0ozsitWsN4Bq7zTe/ftPmDA5Lu1YJ5PtIuZZGc3T5z
y93VgzAVM3sbPCrdjK8kU8aQ3TRLvatW6A6s6LQE0PEIPUQtQX4B7PXJzUjkrD0s
Ja7sUVBrw2A3WHKDAo8ux12+PJfAyglgI88utBMjO+lFzX4857mZ4BZ65gtEu1wZ
CsiiVkbPIqYpShBqmn28UsguYIeBMAdNHnjce66Lao8pc7C8NTn/Jxds3ZAXGxr0
uBHo1JF0EmU0Orhprp3iqbo32dK8Ja+BGz8jaGeWoTYQF5v2Z8POR+enGCRt+joQ
r7bt9AsQq8Cia6AWqhapzAKpSdu7SjNBcQXoAuyBZp/7qvBqVAvG3JOorzXT9lE4
Frc6uzwX4058r9bREWyF//jOnr2IaGreni+rlaBhQgE6kGAPE28kI0UqIgS7BKuO
soLjDbtrSfINEHxf6jdX2MEtbEd6BPXAsvo+uHX7oS88eNBAbRtLIn4OonRRahU7
eAXVOiclR0f47XzujUNBL5A8p3INlwAqg4Y7xTPzAv/EUXmH3uWq7Wu2GyWc1vHD
fC5PniVydzZKQ9X0HsrQyqFKk7gebMsRjh9mEJ187jJouiXLanT2Mbx1J3b2I2kX
GVF9ef1liYQm1lJGqHHwQPLKgPrcZ2rQS046q3AJDAIdgFcJ4J+TYfge70CrFJI3
BQQKz+5xGEwZxUOCcVcFXNncq+Z9ojmP4n23K21+C+bhH6s0AIu3ZL3o2lwGosvd
Rkhjt9jiyQGk41OIGhknoY2jTZtSJSjH9q3pTohtcHbQL5/AGAoSnsJiVLyAMO9M
hp9m++50pUUvkt+MGwOyj9P0lKZEAOdDX6W4G4R6GVGn+kZtMNh6bZw6QsBSeo5O
Q80TUKIog2tNEPLP/NYFG9fa6l5+3TipImv/F4OoJ1kruTGs41SxqZ5/p8eboVDM
tsaCHGxDXfld3+ufem487rDljNsc7hPZ0beAUUHEI5llOURsMvWZZF65gseGJm9p
tS+q/svDE/nlh9zKIf6sxiouBHBHk7G1rP/Hm0wMkjaFYqCTNGZIYOtgvOqnMF+d
04tQBuBoSZBqLQ4m/p0qNN40czVmXD2hWdKkQ45qSxw5FW3+LFOw7twTPmeJCNyK
+DJMMeNBPxOpZGgplxUR1AugRbemda5Yb39j6Q7XKpZI44NYqIiBbPzWjRHrPQn5
2RK+ki7utL+s0xSXjSC0uZIgX/cCl1bIN0SZfPIHKkcMDavmmC0pjzqBUIG4Yapx
0641Z59KuA0MgtIvCEXl2HmMi+Gjf+GRMTNdh4kh18ywmGPUlUpQBmejLLHPBTU/
0i8z9+f1Jl9I873WNXo3O2HGZWhsGp6MAh5rDa3Dz5Ubj6tMo7Xs/Iydp3DlIxPd
0sLR5ZF34JBPSPiAr1JdFgGZFF+FubxrLsOAxvmjoYMhBNvYcrJHYq0wnC8gr0Wk
4NvAtLo65m3gv9NjTdw6JekCWRGnHCWjEw5kBoXkuUH3l6FK/2eu4vGfPQZydnaW
jkIemzbdGojTyMBE8GC0WMYxKrHarEz6mN7xQhTxGkC1Hinxww9eNlcHYgM45MVt
kOcIPBR2qDDToL4UKQ+M6ar4tQBh59jaL7LbgKF20fiMNkTs174mAkH15gFoJPsL
dRqU1AViR4HL2PNbFEL/FQlRiRH4fF/IaFcnTXNLyEqb5cc6LpBSTWgVaU/bMZQO
xHtVR8QvqTuqRWS4ySrBjEpmAMKp3O4/55hDMUjoONOhxK7OiCy++7chxuQNNnUR
xyslqNBQSO3CVAAgo4PIAplZz8nluWNbZAV2Ke7ju/ggwmLV/aUn/7w53Zg5Xy7W
+Gl5mx5b6kb7nSi6fW1Zbf/G/iE7JRAWhzQ10SRepqiEv8bARsM+pb8gpRnwV+2C
l2+FQhsLylYPcZ7HYpbpkzdzjwR1Njlo+ey1+nwp4paHDBCv1YVes28gsTKiwlBp
xZ3yLJn1KaYL8iN8xjrbkpJGUu7cfwk9DHA5ejShz28gb78hNMOqacFCKrOUR8IB
qS3dmsBx7fV6Oq2Oe0lqq1NQFlQ2osRYgqltxCypy4U43N8Ts5Yh/SSunZqRINsB
FADQIDYLG9EGTGf++M1u5i7kuULYoZEo2S0vAt0K1vGMMC4yB5qZWCgtr7eaCt/9
5BXCQtCiMY/zTgIEhqz3AFgSurjwziUWpwhJIpD8MbCooi+9bwyee5Epw5Ku5lbj
p4G0K0yvEhgKSkNLwzOh8SBatNHUpTwwBAKx5r/e6t0wS4GVzhElTLOw/N23OZ+E
69CzNfytMUHDqO0KSDpBOXdP4d4pgM+hJVo7lpw7U1flcwylT6haUoEgBmVHhnO3
MYxaMjUH2qthFvxdc5+CBsI6JelU7wM6E62fN5Hhs9vIFqKva15JzSKaWz2pmK7/
Kuyg8nzre8fs31r5Dz71DugLrCrKjyh5IGijNxrcfKFzN/X6q8KO9ODSLc9KJrvy
ANEnCn23zl3S2+jAbHTRL2a4Q+EGujwXRKhBYson7P2q1Y8ThNQwH+2e0AkfxPN2
QRjCvl7ZFhH+ZXOWf7oUsXafkADSfCVfLK17xaOoXTwlVZOTsS/qYUm2ih2Kv34F
xv5Uec6H0V6kUg4Bdd5xBHqjQ329FKWHbVE8a6+2HEFzEpr0HUfILTjFTeUFGDxG
NurciplmYYO5/Y0vxIMJhU6npacl+XNmbY1w0tustsr5lp238aXK5QvE1Z1dZjmI
rbVCSQduAtX/g4WQQcTM9Ggt4PZNcIkLGit3p+Ou+W6vHsKPc8A2Fu7KIRKijqDa
R/SpYFr1tqmhnWN+da9e4mwvuNQtwaugqXiLP4bNaDGACIeVvOdpdHG3Z0y/FiI0
owuRFSC8lJPUCOubOv1hgsvshRWV9RcivINq9aK1DGq+w3E9nv69eFKBAdpd90HM
/Kwd5JrHO3/FgOp+Ws2zZjX+/4q02Jq01BHjGLqa/xI7YsY/kqUmEbAT3d9cTWBy
Wr87OWaj2JnURcQSRbwolmXFQq2AHEHmRCNyBvWb+i7APC5Arrj6N2zi/u8nLyKJ
F5YfriLvSLk8ND/ZSTww+qbTwJPHRm2yXD7D1N4XmXXOXmujOL5Q0g1gRFHSQ97S
VKGfdY5Ht/YpK01iTyhI4/TvGs/m9Jac4J5kcypBfKzITzPmrAqdJwxzDxt5HUPz
vuKc3Td2fjys9WIvTixppAeIm7qwfHGJ3XZtoynpm1VBVuukSpt0/9EeeDKBbo7A
tmYSHhzJeErEZ8u2rpSY3z4Ws6SjLK4XIQVbazmWf09ke9T5HuI5TliwFvvZCYiL
F3u0E/okprbHl7XApFYivC2r4X8uDXwsOjHEbgKBJu54D13KHJ+ZH7MG5Trt4gxV
uuTdqqXPRqVa/eoBLT64OAs3Whqoy+eB+20+z4UifXeKtQoOBFtC3O9acAIrCjG8
qh3bQH9CT6C2DOzzHzuIwv1eICLy1/2W2T0P7Fkhd3LrHE5+xq5inNRdSm9hVT25
DPVDLve6Jnb4zTFLFqj8zOSS97xTmMH7PgcLt3OeijEr//6FPVO+eJ6rJSDHOwmG
EbgMObhpstjcNBY+kL4z+nLl0701kYDLaSLFh+iiyA1jwB7h6t+4/PcDrPrqNo4f
O5auL6g6jECmZ8rJewPzaPekfKKZDdrI8H9NjYDhFSL//PUXUDgQc0IlIm+KGAse
+J3k1ngfcCu3/KbKrU+WH0SJs/DHh/LEETWqbhfolMAe8xTYNOhXvm8w+IPlxKSg
AqEjWUYoL/+iQ3F017x6paes4QTbhtBrbRZFxekFoCpBlYpvuK807lSQ3y6ryJ/I
o0LElbp4ZfmrVrgOyII0D7cJMp6TpZhFCLBQj3HgVeUvqEQHmEW5Q7O/4zv5lyfq
rsECtkpGMwHu1xYzE7iYYjvUr8ZFA0mSL61GYaAbyz39GskOzb87qSO5zhgUT80h
amG6FJ9wtWjRj0DonyxSba8gNjuu24Iz9eBuNfkW0gcOi7q7kJVgXFtlydo1hQZZ
kW5zROCJlbME2Hgmerdes8yeP326pQdj1o1mcFxA2N5QgXCgnDtGS86sPDCGzJM6
bmaSJmQWG/kYysg2fzEhy1oEerCijx0Gx5ChnCjJQddlGpIYhLr9ZknVL7WUUDp3
w1wHdrGhm6y6xlCikA0Y5QwZEVKLUf0AEVIIX7gRL0Zbe9Wa107Bm/XA0mTl3NNM
nYhiNdQTXhAiSRKpxYL4FYp9Vht9KpTNaHWYadgF/ef6U5kILkiep9FnsoJvZcYc
w/ER9WHneO6UWXpFv4TkLtcgwQZu/ctKA0o700CEBkXMOIT5F/YD1eBRpXx5tI0V
VIvcUboqdus824DfZrDtjdoJ/Lr3LQow0XtIVR/JdSFhJ5njjIT+7Yqf0/hY5rVy
80Ohs48FWJX8GU7Q+PBA9STT+Rm6exJf06I3BlnxueXFEJCiit8HKsxtYn2PlINM
RgCL35nB+PxSjistEQJBbZaFumlY7rFxczmoHTv72u9+WNHWcQKec3VFbK7ldxZ9
RZsciqtRT5jNfvZ/9UkpNqaWksb6D41LRv65sHAFPOMsv7g2Qwl7Wfi1E8E38Pk0
emxdTFo6qdmmPfFdU5ak8TMdXTSOt2Oe/6loXzffyBVbBEUKEcX241EOi5EPFl8/
OzKKXVrN/ymt4YAEugVzCp39S6TFuceJGz4Kj5276e6HZEMU/DpVScjRHsxQOQa+
iR55YtI2wGxWQ0RpuYSGWguXwopT1/9M2CmSKiD9ghkxyA0dLXFsZYtw6SXiviEj
fqcmmPNdbq/GzplgSJLkL7itkTrkMpmi+jAbkKTQhThDO27seosiL2O65jx5c5N1
kh4w8VVNxHXZwaeuCth0iLeLR7V5AXWKnaL5PeTpF+9eTBVYj5wQ+zkYyLjAmCDG
dNn8A5kRdryUY6so5kovGsfrRxH1z8MSZgqo/n4A1jJr7J+/uDSUxFxR4v71cfua
+HitDxKDm4OhxFBhhbByjM3+DIgsVxF72Hb1LtcPmNsRApEIi8O82AVhwVqoGcgN
125g4w3gc6QGvORaVu0BxORRYtqyWUDsnpnMnVpvClzPwUteCTM0uOgOQEz9IbdJ
ZW5I2UQ0LyWnHFVuvQDiQvYTRSMdzx+oisKOi4lVXjG8QnXEIeIfKTtEnvujkf9V
7monvf9/9dwNOW9Wyx3+8+LdDJPuJMHDQ0S+uZOga09hzY1d55ZtACfO0PjVy4og
yZAOfvvgxzQ1zF2BuzqOK2g13/Xsj2vIV0jx/L+u9C66hE6KHYdKwUle1+c9Lffd
PUfTZCmiiauMj9mGkwLsqF2h8+F3xe2LswZ+6sUwGCBajUQJ+RZLtZ0OUhOV4H1s
xV0Bjihl57Ymd8xbKEUPia4PZOQqbiYaaIQqw//TJhiV+nH1NGvZiDvj4IhVNs9Y
E7rXPoL1a+80UFrlgT5wWA/pEiKtgWjHVAGLob4CMIlhqI8Taa3kniKvbwYz8/SC
lsZY4QE3ETXg9DFv/HiXvOAczstyjmb4YIN2f0JKDCG811odQ6iKjWgSJQrUe41S
6t7LlreP6eyQTrZVFaRlSgH5cEN4rsuB+ZyKHO98B4rSJJlQYV1/RaOsrcYwiLxE
SMTxKU/YS8xtI20hmRqQk9jek3uf+rL+8Ff4Nww10G0Xh0/TPhOlARAHCVE7+qnf
Gzx0CBuMAi5Pr9I45nRepqDInvVYpv4/ZdAiTyBYXdGoyUIv6O2VK6JACe/nzIjd
ZAjwzencKtceDlkXVE2HNhI9h+mklOpdGHDSB1oLh4EyNB4BGKiFYbSNmkxPA36d
boyV7x/IrFWfiiWTEP3o+JT1WWEDw2fUhKfxvrrnRhC5umqdr3oCx33QMyxq69nw
akXTmPcObI0WFqndxxooGpzNvvKlXwjq+5TkqC5IVU+PA4LrWofonEkYqH4bbvaY
IiQlxhwHu89xHUzDWKfuMH258IZdAIHIRuJDyW6TQ1ec3NXpCXH6yjfM5nWgZfqL
4Whd+wcaQ+ytdiNfQUOWptvdzD0Md5YHrzaQTCOoZ1/c9H9wz9jtHBccyMTdtBWi
Z8XetiUFUpWsStJAuBMTM0LK+SYTafpLMMTzYmqYtbQ0RFnRLG6OciMMKzhoXH18
+FPvwNHUV+FiqbJnJG3Ebebiwfp/C0QlEgSfaiVYCS2kZ2tVEzMM2y+8B3AlObBm
JtxSk0bMcIYa8RCqqvG1X+9mWwTXwmuCvE82m51sE13WzT+B89HT2nBnNooDMWXM
WqnMz3I2j3UxtxdeVs6jWp6wzK45Esvnr6sThqcTI4aNmudtJFHi0y7whJzUHsSG
pRB8Mdt0LfadJVipkjSTuCwZSYM2uAseZRzkaY/LpBYZ6qkbU+jbQ+Qsq1YHK2tb
7+nU5gVRI8jVu+p5xhlvlaLPGlaoZRGaWeaMBv8Dzs4FAUP7CrOMZpEJ465A+Cd0
EFO7v38pznkeES8yURe3LXh2Y7zpfKadffJPcViRtMOqPlLFQA4aubGvUS7VHzyz
JO6KVpRS065ZQSMKY4ozd3Dd8H4d7o2OOGbPt1Mi1WfM9deRrb3MWitxYmvqEwVT
gAunuoMuFvbmSx3cb10sPmHInlW+wTp2SXzrc9rqgD1KfHgDzQZJIla3dU04iJzo
1e889THNDmf12B6cSXeqE+2NbJjxpAHBv/kqoewPLwOJ2LFXZgoJ9DB8n3D3vtxz
sMRXWEQmgeEKkIG590VnNWpEvMgg0pGNEG8PbAE8j9Hbi5nUA8k9iXdolx172sVG
tSxJz2fNIpdsBQ1p7nnhk/bMbWMv415e+PdFa0O4YH0VoTkwvnp5nWQ6ptwdwEHW
m/sTkAG6JZ9Scnt97CuxVW+8R9MVvenOGFhZRKnf9z80BZcFrA1TsE/MXPFyXhi6
MMymvJ+p8cAr3JrMp9prKfAjBsnfCjHDZP2SVDnCgDU9UOyeN5x9TgLTjfJpPWUi
GPTG8ShEEN3dySYjtmJzHN7/DYiP/DkQ/u//ayDssY8QkZ9lFLbvID6UQDvoZmnZ
FCZ1weQKjSyz8bhjjE9usw0fVO8Ow/0EJaEOHpivmk+AAokvElJ+pgz7YHjqYCek
TuxrSR49SIXGpXnGjcxoh8S85Wdqc+WZ27ub/SdxV7+N6ZtpBlr40wFNawtjxLun
0VB3ujhN5D4wtXlVW/Ym6yfLBJgjfuI+sdhdPkCTwUlAPgQ3p9ZEWgJvkrqV3oKD
np9rHIl5sdCNZ4AxhJCg3gmVWb/63el6Yw9TQBrje0PSjtDOA8OrRxrl1M8vEUtt
FX0v3xT/fsu20DH+cixwfZJD07wo39zMOlgOJmVGITWuyt5OlIKknAP6i2aOt30w
97Ej6xEA0IYOqxLw+6lz4iT8AGVKygvpHjRi43Q2VZqRhRyo/rc8J/407FVSDjVg
P/5GMEZX2+bfxSdoxrLXOj74vf8a/uGxSoDd549FLvaz+Hih8ewgUAS53PN4OzV/
Wu9Ogw3cUisyaXijTxrUnYPdILXK+UYojupM1aJOjcdnafAOIqbq6M9oSOquFhZ5
qvXRsSznBlVdiVMbr2Gmnm9IvJnQFNeVyQRGN3ASUENQETTqBQnMC8rO7FF+374S
WMa8S7NI2o4DE2sWiYY0MBJtqlnEMlk9ckiBFtj4KsXotACVH7ONBzgMVmo07Qy1
cn3IF2aWhLzUg82Nj4eGsG+TfqmChJFg+e4uU33vyQwDq+hgVYu1GHwEbDSG7OuO
L6bSX1WZ28qq2i01mQhN4OFMaZPpJM3wqDiGRzo2TI7M5dFtkQApCZJa7KU75WUF
TaDJ4QeJ16DTQP0YkwBNRZvnH2hRt380tBSPiqyvjFewzPfEuEjRs7GPS1mZuIWj
7g4RJa2WCihiAcmioIDQmR9f6ynuiDOX9dQ45C7Fxox01RIruET7PJwJ4d4QS0mj
XfbYik61mU0wzhXBWnGrs/6/zZt0C2oHdmUSHMROKLsMrPVpSOJaEEUADBb7eI38
5l5mp5igRvsjjTOEdxm/V1xzaGN523mTCyVNQ/dIOTdytKSfMs2IEHiByI4Ewy67
Djg6II3+B0+r1YmIK8Kl0mU2+w2U1ekEwmsDPuaWpU3mPCnURs1PWKF7dC+I5i9I
EyIAFxBdqcdhq5Z40uf37TY/HveZh0Qrv+m26ewjrJ2WodMZqdXCV7XtN2dzgRaQ
/aw19RZfsaqHmtNDrwEDCS00j33F2sJrm/LOjUprPvJ/P9ImMixsptYsU8MCIAeo
mRzIrLAsFuL2GjPrgl04/IzJWf0jgLA6MJXKqv1rr2ATAum9NQjpHmpaP1Iqvrda
Uf5i5w8ZNGS6PlJH7mAVpJZrM7zCISbcYtoh2CNRmLHDUg84AreEMb2a2svrSh3x
X2vhv6gumyvYAhMTMHuNpYw2wXphFyOvgim3PYxM9xzOG8WeTin1VFB4XweykGu5
/uJ14Y8enTKV7sVu4Sr7MsNk43l6ma66lzgCvBmctWs7uZxGZmPGSKBq1lVYW/rS
fUJeT0rtkaXgs2HESEJpLb6706T6YwQKgjjC6f+F+Fum/k5lHsRr0mYwdLjqE7Xy
VuBSFSN+Y6/olnC7aty4YMCqhYyiGgRC7TyKk7NBTx0bph7S7FzTV3iuFq7cNW7E
Ux9LDrjt8E3yTmyfnb6yG+TTZvvtMmlihHfda9ivDx9Bsuj50XsgQjFFgTZgZVBs
LVBXZoBB4sk/hRUVd3uwvV5nANQBostz4NBSuWOry1yCJyeNEKSKPVZ5ol0TPOUp
AMNXbtiLaPJa/RXh+Zzbfqm46jk674eC0XZU1+xMZ7h69Y4yWevWmwJ61Fvs96Dr
MVDipLFfgtK9fWY7T6sm4Bl8C00K8c8yGAQGx18uYpSCxMOYYYvE1isb/Z9as1Jl
yJvU/cntD/9pMgDl6WvBzawSs9fTk4VoSTqNjaLUumL/aqwzeUuVAhHYMHKe7oj7
3ZFI8JcfN666mq+k80MZZ4RcwILN88TUxyyLf0wAdeG2fB4PybEfS2ZYfOX10W9T
mRejCH9WRMKXTBNWYRxv5yiZWKKX/9KgcVN0AbOZPxY//gXzzxZIIztGIhFCI6Rs
acpQr4ZAXErpreQZV9vstV1riDg/6g55v9RBW65VU4oeN/ccK+yRCRJ03EpgFSPm
A8xIQtWXSKCjlj4qM/jFaQLu+dU9HcVRrMrVNDd2LAv4rDtJwymH9mSN9PwIrzkj
zJnVj63BdslGolVMhJQYueRIxzq4Ih+SAQ4eq0DRjWYTOWGX9Y5RLdzWMyRGMEpg
fhl+h9vhdCHtgSqWa6Iaq+c9tiTCJxizGcOfGZNYYUnTONH3fQm81gIwcmbI9Aj0
n+UIxhQG7oEcVz0Sq5dZeClalwjMD2cFx0OFEl+Pv0k8RPNDX+sUSaaI+e6xiGSc
0JJfOHN8EWfjXCC7/ss9g3v3FB/v+SD3JPhQhZ2gv/mWI908hCFXl4Ub0WyNAFk1
YoM7bvzJtv9A+w2/C86OuHQVB9AWwmA9BysvlQKLnbklFCeLReEWKuweTWIyzeKS
SmkKxHgkCwaiGeQWOhppLQ64eLNvacnT+4TpfOJiRIHgya9DFGCr/1O5fm3ZVJcg
XKkgxYuRUy7RWlK4voYwBTNoQCUI0Wt2ESZV6889R7uIbFkvSxk3PuGRlmKVg43S
X4nfsMC7gDAtG3s6RmfMZwlsm8FeUOXsQGyk1jM4eUrRQj1dWLIStldIUvx/UiLZ
iD6BlB+HSAF72mM3XB5qSnPoqH6H+86b3u+q9gjs7zUaiQIKhXbL7T8aaqg15ujo
UNM7Xe9Vc1bTrl4mrpVxCc7yskPXh7qmyCzZQPB0f25BwIOUMIq00O8O4k1/Qjco
pDBor4zwXy87BGmJkkQrOla9wAliwhcQeBE9KZC80vPwV7qrD+sVF07UxbbLPOV0
ULOQ/SYj9wTHjgoIp7nh+5Coyziq2KveCuhQyTptZLc5N/RPrHMpR87mGTBDw09I
yol/Y1YGgHxhkauE+egmst7GJe+mKHkPRPf0c/Bv1x4Go5nM3jVOBm6QFV83BZWC
GZBG+QJFqbGgc1XFDPGZ3Ah4rhrwQTywVgwWauZuqwsRLYjoNEmzJRTkNywa9txD
StxdT7x8R0Oi2EETnLbXxYYunU+GC0sjOAziMxtWrDLUoz5QYZ30JEa3LGFanL7D
5KY7oIVETJnENi4jqiDXhH1EhyyHmjtn6fh+/ZyIZDlFVtMZ2B7+fLompBMN7AxR
ZQRFmnDuqDe/zLCOuMLTLLDfXcf8t/uq41kyS4F79wdSBF4VZYel047rV70uISzY
z/Hj69SzIYUn1B94jVtsrL7iYTRXaBMO8cuoRDXzzyG3o//S6E83yLYo9RkEj58u
wv8dSc2mOyUC95Oqadsr1GXIgXDLz8jk4wPM8b4EApr9i0SoBmTtSjj+sxN1ZUGg
gjmkW6u+ZUZMqzV2knv+6xsn2QAo+Pmw/eQg0jQQA0PQdIsCeHhk3+cMCEs5MS8E
WlyD2Fd3B63wuGSSkDN5Gw6ugYzZUQFCbjqwHXw2Hg3ClMUkaJUpxR7FhJ+b3s7N
zBXTqzU0olcfFIwEkDoL6iIir+PPiGmHhFJSd95RCQuz9jpzc3ViYDK3cJeuAVvs
ABKpO/GFSl0+Jl/aMwa4lU6jXuJiEuzNBXV7WGQFF4bdo06IHd+2A/7Fy+b3cIo0
xe5dJOwhXaxC/QsE2g/AOLQmgn2sv88XxqOi06I5RfkwYDBF32mBda0ldjpEX+4q
2dE5wlv9MM9tiz643gaO1cOyJBzgzqiIKzmwxCQB6i+umQMBIZF4nLrKwvNl62wC
SYVVSnw7Jjlj0c87Wla5oZO1LRxZjI0mIuE5ZmczIw6lurdincMYabHE5gp/ufvC
rZIaduc5UbOwccT34ZUJPMOj8PRUGO+tukLLD9bpwS30GTzXbbUCbPiMW6HDuOO7
FwKpJ86I7RTOKNTeFdKX3pebJcKq6yPnopQ3sE3uBnbws8bemwhr006x9DONZIss
b+vu33ZVAJrGHOf8QjABBy4/Rta3cP3m5JX8zuEHGFzeUCFJNEDQwQMzUV9ev1u9
CYUM+GMBjBYeoCzfe4Z78mgnstH3rjWRB6Ee2Ij0955dfXUzyC2gkzdX6m91hP1a
4/DlEKGHqGmQIolOM2z0ueNcsTINGqj7PD9OyyO38Ul/XzWFSxcCU3nb8UmmrFQI
B/wsRhxinPywhRO2X1vTJsVayfyd1/hSbaYApN1IDwRYjqLJNGJOYqsvAgU5NEBB
D/J18GCpDEnIo/BlbkQWuUAvY1P9lSMkz9hFVdtMrweeNpPf0dEOH/xmmCxpTpGw
kkJ/dtbBpXhUI8lfKb6NMGNSLYvFtXkTnhX9V92JavdUKd9RuV2NhrsfFsZt6e1g
wTmq/G87Qqm6FBWDk9Tb3WAaaJPKPV8gc6HtKNOZ7Qm5CvTSTIAk3Y1ZFckhWnBo
Bio2de2oi+Um7A8kxSD1OEyOL+KVb3aiJUHWronCpi7KOqDwr/ZkhFBepVN/6lv8
wjn0T0E1P4Qlm6DC8f+Ytzb0lgbvJG0XHA9XLbZqKoC0TYxcrqptbREQNzwywXd/
X8W7/CFQ10VjKOMCk5HrbrSf3O994AnpljY1HDTJAnjLV0DZDP1uyr0WafEGcQGO
/O+eHWf8sR+2123VTJV5jWtgwSs/oGddXWTuclbwkAc6YUDf5k0NNtPz8ZTVDkrW
CzaNwWvJFBzdidXDwUumHPlHXqMTwunyNdFm51KGKm12t2e5z8GugIgDgWdNf6zg
H9EViEN808GaqUphO7k8JoLziOR9rO/6dX3d5uuSsuTAZcnZeJGnMwP/2lo06sR5
t9uK+kEpvapSBo/Fh7M5cKuNJNF7MMrnQ6qQoBijL50I6tWJII/W/Q6PfzQ3mxkE
oxF8EHxdxzCiTnVqcZQwP0jeNIKCqeGLnU9Q2CNG8PK5TDPPZljK1wDg0uHbOWTI
RhL35pfJgb7B06w9qm3tsBf0DrijAleOOyZkBAA3ibq/oUjgD9ix1XWBiQjpSGFk
yoLSNP/s2A0vXLIEQ9o8nGW23xn8spS5UwECb5G+Tc1sh2tFAM9cNaTxDKVKdlsG
JIVQFLIwa0c7PsvsTpivJ1qlnBdtuD0UrrJVbQ9bPF2ebzI/OO2kB43zJMUxCH0m
047oH8HlySLOFg2B3QP17/UCO1Qz/++MUd10KNtS2TOoBMQSlRORmzcL3TwPaBER
1ole6sJoheshcnZpeQdUGb/L6uoOVslAVWCOQ8EHZXbo9K3Kb3k42I+u9RfDOhIg
lJVtWMmJEJmnTQM8ns3PxUy9+Rjkmge0mzNloxeKyYpJf6HTHDBjKmpOQjYNott5
yvqJE1AjPeeZhWSWK6GUZ0U4rIRDQOkqYC5LMoqK8EzB5gah2L2WJfb09l3srzVk
vZlIcwz1qGd53SITXrKuZY2M2nmKHK/ekGJlpJywEl4VaXLtj0qIoE8J63+fzFxH
ZYTT8aF7VVNxxTNfqJSKUz8VeC5krZ5cbnuqLFu6Ha3z5T28yY1EFIMW3CI8T/vd
P5vcxuXckgVYgbF6ZXMCQmiHAFM1EPwTMFyfJQ/YAB34lNoo/1wb3d5bTCU+QYZ6
HlB6NLv3D4CGgfbJVGCZnkmnIIsXxzsPRhzN1tTM/Llt5Uj+6xti9ItmwZ52evYP
2fkLq7HKXM9+gPa88R1pQIQ4WfB2vBmodj0ebt6QJyPVyz0sTRauD5QNVgUu4mrr
B1XIK9aPY2RMHv4ohAuJqoRmgWK8meuLhgx5L33eF6BHvWJFOafM+X57kPdE6T+G
8LwU+6AeF71fuyo8ppwQyodZzjPHQJJAhkNlo2HOWkxE8H3ElKf+hHQ2ZYe8btFX
BN9z0ADcYF4dFGMeeqtbmu9Pt53Ug1sQ9nd4NEqK0bQOKLyU6UZdA8Mh5KIUtAwa
dRtzJfDOOBAA3BSpJthY9YENnooPcbQCrNpVX3oVaxugQ5FvEn7wM6QBtLUFmzdP
vuT7CDqIqn0XJMIDMYmbIaVCgeXA4qZoFl7P9zELTjwGZ4Is4+aspBpVARmmPrL7
j/dTHAp72RuAsxEEcJ0CdG1TPlGuVVNASv4uxRCEWeLmB6D9SubWB8VBIhYT2sC0
dbXpcf+oUPyucri4REZydqBSh9JYOWYmKPD4hF55OuUgTcmO0Z5eIM5qOsEfnhq9
S4tfDaWrKM5ltJqAFfQvH0HfjnRcxE/D4ImrpowY5+I9LCXrcIgxL81hhNATuA31
QUQtcBTmNJJN0RE280ej1ss37ziAeLUpk8Y1QcAYu93WMD/j8lVPp5J5G4C5AG/e
3b6WDQdj4lMYYYM5pdA1+5yKAF5UtwnyRvuc2PhJLwTn19OGYAp/NFWrWc3iJ6e/
WNUeJ6TprvfR6aDdtmPbM6rSrM/X43hLh5OwJsDMTu0ctz1mEJaRx2tkBKAINl1O
PBqDH4t55ZGEElseIFf546ixAqqXRIGCHGXX9ByBN0ze6eoX9GXtv8INPJ9rS/oK
9iKHQG6fVs6bjQUAn2/UGjvwt/GlsG9+GfRBoo7vU8sXmGfU/1E+jLbFWkvkRHsi
F6K91KADXFfMB0eAeFAuQ1zpxlGhd5IMsAgRWR5IG+OqUg1Qm18KD5QRmArKw3CD
BSc4XKEyShIGW5FMDSqkDWgTyQdT0fl5Z1P7Jwmc8gpsCFcqPTeKb/izOW6BG2+1
Dcb9JuYh9vjGK2okhXCb3nV+6hAALuEmtEBQiIpq6Z7qsQQVJaYEXGET1bg9xJHo
a8Rp+C3v6bwXOM9GQeZ+9OxGy65HbEqL2PGZsVjCVjF20H50e/qgXEWrVPSjSxij
vQfgfVfOL1W0YDgVdwtYkJAE5mujonkLx4PKSM6wFim5flcYiupvs4odfTU5Hpp1
l7ibbd3KJ1BpskWpNO/oW80IH4+jPy3ef9/xvwXgbLi9byWl+R8JDksXqcVQWVUY
lKmU7il0MlWMVJNePgcEYf2AKReS3LlWvznQREi+SVPr4zGaBdxqtrxoEDCt/l2P
ThLBra1Uh85NL1w5SDc1+sXZqj9cIrdnaIB8Il8K5qlM69RRCHAcW1aRM99PI05t
bgtfzyaGrZIh5mZDy0Hi6zVzOq7nfyNtuINZAkB7stFoPmZt5sHV81q2lSpbMeKv
3viriER7R7/IrZQDqdNCIhwsMSsDjdKJC9R6zXQtf9STiGtf4IoPy/OUA5qL8SXy
YnayFzEiZa04bpjU3KMVLYg/Wxh7RUXTcQQECea9vJsIevtulNxbyV+qTKVVnqq3
xFQBceihxbovsgSFaQE3iQlNA9gFvh/8PtuWFPh02t9FMSPCSDyvUsL2Xt39ZV+c
hbVOnlfJxLYeBXyJYdh8NtEn845foxn1Gr+sPqo8EuWN2fBi6FHDFTmc8l/oEaPd
sOLna1SiI6ShwX74fu7KvUHZL4ThP1s9o4E9pVOVO2ci0/KFMMzdh0q0WGqkabMr
qF9cs3vy/Wq+kq6qasGrtsZTibXR9lYatgkr+FLVqDvDp1SBp9pRHuuFYd3Q0la8
r3/x8BdfqzrmQhVozPaRAH3bv/PKx10rhiLVXlJluxJIAK81AO05PgIFnSETWSu4
vQA+cfBIWgV6KGbpVP2VK4alMm2J1P5CQO4JOJeF8uI/x63+kIWj4guHpk+kIRFV
IJPnjVmqe/2PSGdy2zKupH+ntzbijAOU6DagKtMOF+hRkV9X42lcunLmGv1hEexR
bB85URyUXEvstI/SU/eWLrA8am+QkI18HG4pIO81vwBSs1Szzr7dIXzoP/MpItIQ
WvH8HK6UKMN8FQm/ztIeF3c6EZRxYRL82dBu11FdzV/mzQYj7o0CS+4+2ueH9gZU
2MTtLAFY8KZu+aAGsChcNFSZTlJuwAG2+O7syxDwmWpjzKlsI5DoxZqJMelJuLxS
WUb/is+zYtHsKKPlYF4TFpUNLow37XKUaxtqp1NoUnISmCP0zM9OlhvSwSlfl4w4
Nzj5tK1kWy7PzDf84jH9tCpFtXtwZ/hnBWj5K2xhc0ubd4IVcNH5xcnf36Z/ltHu
pN5HhohQxDzDzQQTiQYrHJ5D/3U/FyKC7PNdKlsNZQhAwTd2b/Qos36lQpxanA0+
3/aw9kcH62Xbq4hdYIQ5TQ4qKefvup8PaBN+5jNpVwaloXZR7OvziW3Pmb8DaG6f
oJHt10Yx6OJJfLFXxYvtdBtPs5tDUis1gWfn7wMGCyg04c+rNAJbxVPSyJpvyuo6
gDzNu+2DeYUJ8jhr+zwAIws5MP5YVCGxzU6AAdfAfzAZpB6afYrh6MiA4BKwWYtm
AF9MtLYdnrZvK79SFPrqZg4CltyoG3vIc8D1ZXCFhh1xASlY5iYn9Do1ZxTM8SDO
kkYtCo1OaM9yr5OiEuUWqCoJjzR2ZkBlkKC5z2bpDjLHDIvEuCCq0LSKrM9TEgr7
2del6BNVXCEoLUsDPUWn0WE6jclsjQeAyPTBN8x0HVjeHaCyU306EjBLmgG6rgQI
2wNj6bpn3hnbWBkdz93Op9isKZ93lwR/kwtu4263KlgHV6UHGOSHmunytCldern/
j1dY1QwLQVUyf4dAdpNZFzcJgOwNB10XPbs4I14T/Z5t63OJFIbQMAiBtotHhSl6
9bZQKFOCoJGksvHfhS0qC9SVILEcIbGpUUnSnOeDc8fLDwkFq2BSAHn4TOa4eJvS
3p/rDXzsglbQfXAZ8aHYmuy51x3LlJtn2wG/+DVXciMJ6I94XrHrnPfaHG4TAl7s
3ew0fXALDkqnQKLDEHtwWrFt1wSb05v0biBAC5KKD0WiNSpkyf1e5A/gQtRSNlfT
5ubnveEnWelmxaIWlWVK3SrMM+InsRIzvfYSvbrJ8qMzfZC1Oxu6Hr4/gOWnRWHX
2DykLv7SVogsIHlMvIR1Q9xE/8BfmAPV9xI1PGjtoa7Xa+AnoYb3G9/+nMmHwIOW
xqr0aoDYpJuT/3WqL6H/8n4BR28LRADZG8z8yBKtzp5yDQisTwXnpjL0GidI63i1
0EZ56dP42Hiu8h/g9+ohOrVXBjd70TFMp0GE/epq9kG6P6KJGq0SZudzKFbfEM+4
2z5Sb9uSksIvaWivYBPXnFHBkyBXVdY/SK+a6XlbLdfP9VTQSMohVz133RM+PVA4
p19RPJ5skpmH4K30eTtctzxXhm9E+BbgWWpWqt9/dN+FgqcNmhiokKT+zYChNe03
KdWXAjX+SItMTmebKch6WVO89DGaQLqOsYCrnbA0PZP7W5sL99GxcRqw2ur1i7qh
luVlW/y3TWjEm9kYuG49MP/tiKR4uNPwjNTUKuugeQT/5OhJ1zlkDhks5hthrUBx
0cp/URWGaYQL8j/PDWv94961bkn2CN6vucSkyC7gzbjs18SUPsK4tVZpYDHsjv10
gHXAkBP8oMi6zHqJgWLsL0tAF9yEA3WVNKcmQ+EqHlasSRbY91ePmSluu6phWqfF
+9m+gMY5atk0SH2RZmleBg7hPVFquqh/rUmgj4kPCCGVPIoRRF7rtI+34k3OVgnq
fGvMIZHIn1nXpRCTdEHZqoL7GnTiAe9TX1GCr8KeB6XhgY5C/RUQ9wl49OdSM8Sj
mgYgdtJLO71qEB+fNNO4r07nDCDD6c79IVPSWs0DiTAu6OK07+vqEJlQcs7+wa3p
UvClQng8M3ugDF81vKNVXk+hGKpreNrOZpdz4mAcr3kDQYa5GpAK1Y6dPImrJ35W
aHHIFtWOvDnlcMxdfn23OFMB6c1gl8wjWFmUtSHbIBped2jMSPcz9icAB8pxSG6K
AMmihSc6FG2UV4rhb8orEA1/DK1GChWzzAO45EZaOPPHPOSgKyzRZ19DwEz1xIt9
e8fBvnQDrhDjEuqfZKIGnkLCugB2/ORJ5DPG/roAosmDAXUyOssY2sJ9VJNG8m1y
MQB92uxvOsxG4qxmpk6jTmMjpKwQVaBHmZr/oh5HR4yzn83IABlN6EjJRvTXSiJm
tXe36W5m+7NOFEJB7Me6QzpIWFJmFg9JZx9+c42lWloAavFT4xx0QjMs9zSmsRf0
BM7jtBnpgtirOdEHDZiMuRjphIoOicpSJyXr1GQgUKVxe2VmJasWL/UzC5r+UYAm
UP5Aixs/td3cwnWYMFb5xxLjnw8y+s7J6F0pbWFXeenOCFlaQ177bgbWFoPAG9Ea
vsXlT5DEQEgRdClaZNT/z2eMydHcR4tFZr4Y4Bi9mkvZz6wyV0MEa+9zD3VJmEhL
outWYkr2dMrqYRllVZmYvtOR8oE8DiHN4n2tpaJjhkg93uhKe1mZjp1Buaaf9MDW
WQiDA5NRP8oivQznLRTteyXRzCGNjrmGODf0Ht6hLjuWIh5rB48jNRjdcqZBVu5V
1c5dtADkPC7NVfuIRM0e/FbG/2DtNCdH56xdCOgivD5DYAxonYdwBAWRi8nZICOJ
zdLKWRwhjYdEuDg8fEyk8FTS16VREjLMsQCy5ooSHwxTG8dsnMnU5Koq0BM6jteT
pUJJqIdXSYWz1u0+/j5WqVfAOT9vzJruax/YhB+6kF8xpPAOPmky+9XopRq6wFLh
+K70l7OixFtJXfIW+ihSHFZj2lNYvYJbtkdJoS5BB9AP3m31IndkfgWDuH4WLWef
BwXR7C3TzYmyvoYnUsWTONKxnoQvWNUofQzC/E+BFBOiVYJhwauqF0QyCfusCGEM
w8zB0owq0+BxYHWjeflP+zctJG+juCAWL5kdhH2lUx5MWPTJ1WwinjLgOt7shH/V
aapW0NqVXcf6oRGP9/gTxBa3qmLfEaAEqUghszrP4NVBomcLFy39UZhUq6uJLKj+
EhedfOWby9c4fSuvTETcsY0JdEB3OiGj7/1M4WiW59cGtmHojxj+9WzaZ5Lxriqy
2aEFkbH8DCgyfJ1ICjFt5htwKlKxic6PI+QiQn8jXOJeto5TR+9sMu+sS5/r9Xy+
Jjn6m/P7ymP8pv0ZhtFbMkInu/ghrH4PUIwgPNBSPhHQXSjCnPai8BMGixb7fiZH
Y71MbOv6H9ofCJgi+Fz6tno4OrAfL5MkXuuqvSqummb55wT+nqefRR/oFt2zM2Ei
p+ON8DSe5nhlHKad6MFxu9aC0MYB8I5czsmqNT9oJbs92soS292/IS3Pf7FCjhpr
1baLOYH4QafBW5pNkXxjrkWDUHQqwMn+fW7QTX84SKiipfqzSPUOqehnxZj17aJz
1WJNjCmzzC3poQxVWVbCb5WpvxXoVmmMy7yvFwIWJgjk8Xf4pNp6qKe0i/t5ejel
Z9dlPvnfZYVpJ0pGlvfAb51aAjaQ1+K484cR8GkHnm6Ev08NQqeFlOzqOGsfbmn/
O11lrRvKXQc3afQpNMX23HMWRXVzHm8H5IM6MytvqRg4SzAYIDKeOfMvK7DsuBpR
0FgTF20JUglvAwy6XhNyM0izjhN0druysZwhi1/7etfVeeCPtsqk4elckjqr2GEu
S+gPHPKZvdSiwCa4ssXUEE1994oeBTqQcVfZ8D1DqrjQZPIlztRDseCgXOMCerUl
sQOkEF9tVDoTqfSByYOOZXcn8pABWAYQxC/qsJPAR8vU6AHH67nOPppchu8hY7mX
bkfSpmw5649Z6arClCRXawoWqom11Md0mzyamAxOhCSbbsfwU6Duzt36EW34ig4v
d535g/ypV23pLmNZ9qR6hn/FkwKB2PBrYzeAXb5h5tNRHCKNumKU9EEKrYI6OGZ4
sPD5XwLyXO6JTRS5Um827O8Jqmge4rFz79pwxV1kgKG+vI137+8dj6iXl+jOZuVf
oaavNT+b8vyond7tIIxL6e06khsSFEl9/X62O7CC54y+iZbKnY11joZg88CjhpU7
Yw4c5HCiqR/8Y9LqPDb0sXWEaOoFsgmqYKWf/oxOnXwozaOnCWgPamm3nJfWjzch
lDSBLc1DTslPOX40fPFCYy+0rW6RcoyX19LBJ5Ma832qfziKT+F3yzq/VPmF/EEO
3Pbi96a1kMdFlISHrBW9rtGFV+L4CMpsqrKRq3plFivEphZ/H23OGllNO7Clv74a
sZIfdtqz5ZNXEWm+nZemcgD1KcyIkYCE2Qa1nwQcItYG/S8Vhl4+nL4KV0Jkw7Ec
AUnHfqXZ/7z4dTugklcD6RKzu+NvXsxZyjxsHOazYqhpBuvQRv+OihXr7MdRuBdA
KXx8IgujXek+4iKoTjKS8yvbkVUQMXF58EGQi1RG5ooNv9vtL5FNzrMZjD8p0TwY
9cySb5rs/JDjQ//+6Vhrtpr9mMkOPkWcZSP4g0+rA3QVbNjY5p5SVFv69bB6Vvv1
T7qmwSX5l/B0xMR+r09ZK0M1DAr72rbDRCvAby7/s0NYlfZtlDKNXk55KX9GUgVg
hO7WbAe2DiWgaWq1pMSFy9vdBPFYL+eEWwEc+BCjffDDrSVRMiOmuQIFWOHeiaxf
SnPN/Qj+j7k4V5Z3hnkszwRVo1a97HxK4kgrWHKKQU+f9nK7T/e3SCpJo8MTQuDo
vO//jnIh940vanQ5FmU8LP24KXGuhABnp6Gg3Nd+wKLBxMBCgyXM67zSNgTLzqHZ
iOinM9R+ii+T0FpfLzvPcxZhxXLcQYuS8a5LDMlxwEfX0E4Z3moh/sXiYzxeWAZf
C9Z8VM2FKlhh0jk3zRglH/4KO3cr2PIJ6XtAZ9R1SC9PrCYOo21P//fAuPEYpa3I
7vXj6kadt7qHSAOaaGd+vJLon2al6Bdbo3AlAg78cAfKpil/SI4pFKrcfSUbf1wN
u7cILDO9RomDEK5Sg3VSAU2fgYbLA69JTS4cJoo4GVn4Z5G1bFQz+sxYTgEbiqWH
LfoWcfCxtL5S7NfvvqnDEdChip5/DhH6rL2+7hZJgiqVIMicwPa1vcjno+DTi//F
n3aD3+we5d5SYkemPA0vODL2KDN/e4T9V9Cql9rMw3Oj5rjJvpSw7z5SVVs76aMh
mHeBTXPldwzHxrvT0IAVmoHVqjqybQ52OA363w+piWyyhbwhgsKisIDfUaWSVneb
/m77MwlZSMx1ePAdseXeSBmZz/Sfv0Ku7RN7LLeRO1G9CUVqwa2kfy2qGdTiUV/0
QFTtOR145uQ2t9rN4ivXWoluDZAtNNOqj+5GaXKmtRyqp0GTYwXBhr12kpN0uzlw
ZvVVwGbjG7WUfLcMkYDm7hDCcKlxGexZDnTpKoRFuWM0PdLsQCbOzsYau7nvUMte
3lRJXItqN4Um0wJJD+kka6SxMpwDOMsMZc7kUXjNhZtMnH4uH5sUdsdg1Mw4sZBk
fik0Jrzhm3KYOe9B3hjL5XB7PDSWtaS2hjaky7liK3lpS5ILy5/ciyU2yJWfWhnV
4UaTY40CVNomUTrP2N/yx3EVUdOtb2pWxnOH5JJOPo9S74qsGn68UhAOaxcjQWJv
E9kPSAUe3LYxqoensGbmYDxCOlfZ/Fo2r8pJ2wYEhUM5y/MWFRVcgxV+Yxj/SZMb
DSSLgEJJNRPqZ6XyTnUbZpCFABuKnx1SHbN6/BINiaCPEy5Aye4GM0pkanBa/S5C
LYMptwg7aPyR/ouunrVOX8DUCfjCvzBsk9g2UQp1EtPwnWTCJz60Qu4vVPulmt5X
9aGHhjpkxUat9qrh1GFTBLXYN+5QFFDVpDYSFFDyDuZFkkTo/FLHA7iI6FQXB5I+
7bPlhT3f21yQwWF2lw6xLsOp3UpdLVN6cKokVVV4p9lODNzY1I1MBRslLvyt+mZ2
c1E+l4AmOYKcFSUN0Z8nfdtjy5OUR0uGhg58JZIX+KuMWYJEe+3jUSoUloqumdBA
fKAThO3HJDh/B8m5CxppovKRrT+bOOYVW1VQiI3CMIpILWYc3pkDhpvfdFX633bz
L/do150H/lgIAoBDhR8Z+eU0+N/Xa/5DOX7QetgqP2itYgdFYqd0KMTYRukYhrsN
SHXNrHTE6zqqhBjTHZLAb8E1mfvFagrx56ahIh28nF2V5kRWIjkKeNBG3OchC64c
G7VnOuQndoqtkAmBC0ZawSLPLxVHUxvsX5WTlwtodAKTCK+HvvvNHSMvAqbMjFcG
8pt7j2U/lUlA3hbP/gHORBZrg+lbZo0p66IDE/vMuThrPL67Mghv3BWwMNMjnPPm
IY8BsKqc2tYugktLhAN5pLGeBa/JWdYcedOU4Vg+4a8mu7ITe7MP8GTV6JQXWjXp
NOkCXEvFMkZc3l/xAVPr3wOGUGNXPm1YambZJyo30zJPTC39FT8u5ZoYSzo78/aX
ZNFkIj66v55TzrZvYZ0OFS9enxPQliaM/f5MGT9SDNERZ3GQMojGX4woBYGNVKjf
iSR0hQnPYB/Gdw4n32q5y8IwZzP8vuuCmUmJs1DznrPcQM2Y6ucjQF+O83AhS2mS
QJ3g/yFkjRymMh28zszRSf+GCAWYWR1gUvLMyXtQYHRU//cqxrJRT9ZL1mmo/76R
DML4J/qqELCstIpSVfBd7Wj+FeeWNssicYVPOA2/9M6a/z4MDZMQ23LPSI4KDX6N
2FNLOTwbDwYaAwNgN/m9KtROJTAHilbHjnpVRt+DnWdY7XJY5088giwocq4mbfxO
YSbhxwNxoa8uFvS2H8J+xTDTiiA4+CJXx2BEZfoMJrFz2tkGwU2QTxIBLzgm6sPB
E05IW+wlblz+pRCgi1weYKEE7r8sr0NokBHxcSUPut4dy2vG/X7/iDkrfefDmHJp
3yZJHYN2h4qco0Fvi/gynwVyHBzkKFvsfnG7/sArfZz+mA7njy67DjtP7CbQ7Ib5
jH7Rp5acsGaV6lBMKkYQHcrdLI6FfzUUogjzSAOaUWgRYwTQB28eWTtlBDqB73v/
etfaMfpErJJ8dOBzxRg0U7ctDQ2wXAcvtLllrlKWfB2gXxgfsbDbiyfqfDT1UujE
sRJQivyQAWY1YgddjQeaSyKYOUfDw75rR5AEyks01muMzzzbGI7IEHNaN5jO79eR
izsYPDjfIqV94iiL4lkYB4z/+cqRXiwYI0pyg58S14+t7/Bs2LwqIR31SYQjF/JU
vVnIZkItdLlYp9ORiY1OcXsPKmzwvCwN5VnasSfd6PQfol/vjWNPVl3nAk0EG8Cm
K87n1xJTqN7zpzbXhdRohE5aOAVqroCfi/LBNiT1CToOzoGY1uQFFNxaodR3zOPw
uqU43IbvZilTodYIi1gtDI9J2zxDE6f/X9IG1EhPFuV5M3xMi5X9k9GlCRCSpkSu
yWWPSsryS3wXLxSegAsCBpyORWRk2J+1dBuGnhBLVEKGb/qJYqnVS8iY9357FHUW
feWEqFnUBKvpvN0dqI68EkUoWacexojUnqZF7Ttms43EDcAqr473f0ZykJSNV/G6
PU/w+3Jt/c5R/MF3zjEb9w1qJVmMj1mSE+2BWQ4LdsBVcmfCMOHnZ8m2BR3NMF8f
qb5p5+rUcJZ9zcOPYyNh+Ko27V44lc21sceZ+Dv3WmUSBVYmqvceSuwMSnh9Nprb
OdW5vpyxQQNlIkwqS9gNOCanmo6+NbpI+LyqXYZWDEoNEWsUOp4hqymXdQ+CL5CJ
rgmQ/VNGrK82n0BF45y7spN3Z3f2ROi2vnbJfhWeru7xI8ZU80QAIKeOJsu4lBLQ
ucl/SPt0B3IcETlbP3J5xkujiyDWDmPojg3SjJnmna+bGgrLSB6H4e8ElXaLckZE
C1LdZvYVIFWbrD1xD5vpIxGecYkCUxKLqz33fwD9H0vSpw0ZGXuqjg47Ec9Ru4NA
uHFNlhxsrTu90VFz6u6zC7Ty9AgBCDkn/hDdTjIOmXJo+o9foqgoHNRYb5qUWH/1
32Ekx8mmtqXL5wRFPNXpz+Rzr9LtjIJv8nwWBQ9iq7DhBZGxOm+qJvYPWwCDc1NE
99aV922MI+ahWzLL4TuAAHq3+FU6dLlRh4HVn734NCswvVlSGWtn1y0xtEK8gWjS
Cy3AQl4L0GEtzk2pB9e+GLPtVD2ATL0QXKRdtA/1GhLofH2POBIE0zOMzGNcBk1s
4MJcETL1Ju3uWsfd7p5tQGyN4biG7T+kQR/pTCuDxJVBOx7hBlBK+mN+B5bKDkOI
3F/3ZU66VRMid9ryTA1QNHIy2kxjHW8nyY3fg1H7IwcX9Q5Sm3G8ON7nIVVtxTvC
zx/UtrdH5EntNyo8JPWY2s3nLplI3B7b5S3RRZsatiJ5wT9tUwt8soYENjHCXUFF
w9WViclx4Bo9QXl+RbbcDkEX2ZhM+qOSl3iFapUpoRsY0KRPTd1Dh/0v03MtAn0T
yMq4NAE5Fk7EP2/lR2WU9El1QXyRz7kvztYqgIna8iiGdAm4AgclOprwLv0n9q1G
c5BPXa+JmCVqRajAJD8jcQJOckrtelqbmk87Var/PH0xVvyAOdIzLqIjlAIBiPJy
GGjo5UU5SZqJ3NsQTqxJHoWU6VW6qeoNwsMQsntlEmcswQq8Mub1YgO1iDg7cuMf
nwXM3+kuZS6E9Zo9pa4S6MCvfalRwJ+5QzcBb4DuoPH3XYQOVeiNmqdzwboDVPvu
Hf0cYtcQU228jUEvtTh8JFeRbK+hKBuXPbmiws/iOskkRceIGYZYkGvCIKwrBlD2
8JZk2vBbFnQN+cMJNQ299ttEDOxJx5A99O7hKeAtS9tEZZLsYwTul70BrJre9beM
1vtg1P2UxqcWRRqWgWqAzh+NPtRXIvFD0g4mcadYDPeh85ZPHCKl1Q52JmjXo7Ok
fBaXZ/gJTKxcwocl2BQV4qpE4a/3dPfZR1IITgKwASNlnXaNLhXrosuH5zdRIckc
UxsqUEN0y11T+QpX55aC+RHyZVqFX2lDdkenJSxEjTuX21phcKyE00gFmftlFI6a
omwaP2Cs6vMAtmIL2WllKz95Jy8PXh2W7lbsM4dnqhjD7/1ydmFuqGflA//Pe4SC
/c2ulLB1WnJUAeRh9aTAniPqCtc1hmm2fEkZRTENa765qYGiqV+BKSYkiyIzfkjO
Yj96jMD0fYDB0C/dyxuPJlqSKRukEJUZ7CK5TwHSGe3A1qDP7rh4pXviUNg4N9bP
AVEhZSSeKykHD489Dii7NZHv8CIp1dKLatE+pp2d1s4bYKxJFBWqcD09aYtVfDtK
vrRzVQ8XqMsVjy/PTA6SJYoomX7eqG6vWAaCkwhV0CW4Saj5pDY29oJftdMMp8rJ
9//Q4kwRCnLgBbGlRVWMbmPVjKQZJpHaofxg9Na4WsM3wOUcsOQcloU/rgEh6zgl
MJmaqoHLD3VZtUA6hKfmEW9KRDl4xB1hUvg7zHZYavuZp0qzCLM1o5FVNo7E97U6
PKyiKOk2u/RB5YfSt4SA9P+B9slag2oGpbdj7PVEgo/IRYW7YgeBQppksVkJXm5H
ZSRR8LUTcgPlEpyArK9ntnkJjNdcGA5IHmqAhwjiM9+tvGn8RNmyDA0dJ0AKGePr
NmVAKrS5ZVspmq0ms9JQQMICm04VCX8ctkPs3s++byWiXlevlyL1Wu1293K4qRgc
SFAmOKgIwllg6VQYepPK6fPhZ2hthqh0L7GkBBUVHJWYMA3Z6lGpTRmGijJkmXOS
MI8br+KSlk5RwRzaT/YMnFAIN2ngqpVX5Vu/QB/MjBK8c9cgA7iAmG8mjmWwtsUb
UEqcurcPg6vum34d9JG3b1hp03wKnjXnRC2rV9gNNehd3ckV27ItSAcOjJNgDMn8
bJ3bUkfMmjmejIbLjbZ2gdnzCH5YfVY8SapF3AexGja912OrtRFeFFX+P+v5x245
yX5Iy4XnYClpc35Mw4kagFkyRedlhatFsaYLHK/lqyU8mzYcuVmXnoJ7PHLflzj3
YXJ+rGb5CQORrx6tDDzxwnRl6waRb6fwUr5r1TqZCrCkhzlry6cVzQkxMDroc8vC
oAWIQ6cGKvWrvvJAMoURtPtUTqcyFxY+n99DmOmvJXQ/wiMXNsDQCdMCg0z2Q7zE
qJYDfmiitiTnbmxqv0Pn1PaGt7NvJhldol9A7FZPFn+R/MjWqJH/oripDoEpSeHf
EipwqxqXbqBUWRiD4mlNIIDbuVyqX279S9UOSIwbXrYk11OgPOneUDI0qexL/LQW
xYB5LZQiT6anCDLJk3RdyyEOZrRz2gu6Q7RxGJyszFzHCGMr03GiR8UpWomC8phc
1iirIIbUg9anCF4euuqP8YUSKpuTberG3IIh8wjs7VYd9IcgKml8u9Ei001PfhjT
6xY7pm5r3ern9k8O229iy2p8hh/+vzB22ZAU5pzpBQ9vaqBhzSQTrflJMJE7hdb9
gJn6t90fssU3A9ZtgOMXmBYzSjIT/lav66ZaVKd82fy08bHHeu+ef0K9Ichnx/+0
wPXegiga1/Gz9qUmM4ng7UzXL6qK0/9LVwMpPyTIxh4HOGTRLK9B3uFsrSDQAlHO
fqkQSKck6RTlGEgo3w4d37nlzh/mbRXlURUrv5y/9NnAkS+Uu2vB2R2+fT5t2cD4
DJDVvtV5FbfBxBX7xM30+CNT+7BPWYWj0hxfD5109D+51E7FbGQMM3xebBwY2lYf
d+wQ+qp5amPlM3Yo1KkEblmji6/m34N1arUlwdEsEQpWAZfO/KGLVxk8GwDMv5k2
c06F1HXIBLEbSnesvjs6QPzFQfeLGO5QoeWf9Xk2Pb6BUg4oiGMep42uzfOnEBLT
8+FicZJJQ5OGh/MaOcImzLkboR3QFbWoJx0Nj95Ex4uzXfooul2Pz0lYs0C/Q87Z
QjTTHULEoEoVh6FG5iPezPVqgf/Yy1NCki2baUi2NPk7LYEe5P+OE/Njiayaoz7M
J5/3ISdNqLwUECwL255xP2ZICAL4gK3+Nok06vAkuv7aCksDIS/V8ugaJp5YiGmf
nKa3raUzL4qrWD4Sj6VBfooEKYY6iB3TGVI6SR2xaKNoLikrcBe/3yWXNjpiLFEn
u/I8HPYiF3tNnqV6nsmSTUIGsSokvg98Fyje9cgF4zJb0Kt3yW4QdwDToYNEy2vw
ta/rFiQRLGDN3Hhmsc+9rrDakCtf6MuSC1mWw7lAfk8AB5QEr6gQkEaGWbvz62Fs
xIVYNbmWXBUD7wqtxUwxYpow7MyBuPCwf4ZHMhbYX2s7crj3ajdRJf3TWRdwd1hD
Z4fHV7xrxjwu0Gh3BkCluF/w+X4AyjhS2LCYrDV4//zp1eWVuEtVmjnuC6cXdKgU
X+tZ7L8L0mdbLPA5aqpc8r9F6HhKzVBENtplfhHScKe0b6dWkR/MZ1BUVtI3m0E/
RJHS6QIlnntxj9ioF7RskfVT4We7e1ymvO8186QbGIN96w7YgbOdS62UtXVRG4Dn
BRXdWt2d0TBO12zDqndJ390yIiuePe9V8CsKIh6XETFfXAr8NJMazqrB1FjX9AY+
ZhzZDi5CIgdMftvY+TuSOpzQEtrf62YoIUN8Txsp/WObjDgpg/1l/BfDCtWI5Rgq
sk/BYcUG/QjM+KuZkllmxDYnJxb81dD5rWDdsgPUlc/MIyhl3qpYewoGoPcEzf2w
lJTJx/e3eo8woV8RqrTA8wWzGPUcYORN9Z3VBnwYdmGXXAJn0cTCfqeEAfwlibwm
YceC83xYoV5u5lhUKwMiRQC9QZ/TpWkMw8sZZWX8FyRs5YAgvhkCszjdPg/JDiWI
k9bvwCTXi4q7mW45YIdzAm9JYp61VS5PV6rjeAnaV4+tC/swmE+CrP9SD9wVYxP/
nxclP9gjz10nHa/9C1Z4lRuiMik+Jv5SB+tVMJchtbwuBn6LFa9ol8NskBGGzNJ8
+btu/OKptusCYwDrA3M7cwLnQpsj0fJLlGvI3yWKPiESPbASqN9fOm2C9wuhXGR7
Jl5Mw2HmJkocaL2OnONwrZ78z/mU+TW8q2P9Da/RAD8Q5cGAThgmsjcZ+uQiScfg
x5Dj8/qd/4XSdn6ZUGl2R87SVBsrezWpuw9ajDE6eHZcL5JJiLHEjEFQ54Awk1a6
OgwQOEObDYBeKWDMPK+MdfT+kLLztQwcymbSPMvoQcwdkqa/9cp3JKR7dMqAqXdN
I3VEggSbER/V9N0nCtGcSarafVJD4rnctjrpyQz/aQuYfnjvV8HrYWKwPwB96Q61
GMRjQVwFqPmJWx/rpIF9sA1JX/RO3j5emA6AkHXnYV6FnZ49i6RJ1mQ6H8cfS4NZ
IAw7RjTVt/CIRGEe4ZJwauyoLAOpx7qZvcdbgjTAbgGMTtB99oqmjzLVfiP0vHjo
uKn0jjKVaNtEDlro178MQY18BHzJ0EJ4v8n/nTBxf5DFx8ccyzsoMvpiUdwE+5ov
rLUoA+7slOfFuA4AkuMrVL1NnoB7BOS8YZ4wFkPQb12aVbeqNk82UCSCQ6jKIx8j
+BomvfFRME6l5OgpWidzgFvOqbBUTsB5zSwGW3bwiyZTvn1Vq5AouEkdKza+hni5
q+xjuKKwi4vmEdsmkY0h0YNEfh1uwMwfF3aX10Ho6sIKa18gNaxDGfdm1X19dage
7cFIMHDhcr/JL+bSrJX8y672o4f8QitmQ5vEnTdmVA7u57vwiwyBXz0DxdfdV828
C8MOwN5li1ngT/pGV4vuYLyhYyyztA21hn+uduw1fnoyjejv/2YrqBzhpewwHK/M
WOoZ6v8vRvPvSbxVUO/ZoZSTQlGjimKQOuePY/piz7gEdRvqH6Q/NndUwW6Xi2WS
xKs4FHMFzSHQts48Mz44nHn02C8BxdJl361U/jPkCPK2YR39ED7QEq5yJ+3bAVFT
nYt/ZotbgYRmJnVjCHdrHz52kHumN7vsnyqOHUiznE8qMKJmXziaTGdH068U55NI
TwNWPdnPlP1ZPDzVFSxAumj3ddTm/AS/qVWTpWh1BE3xX+rgnogXdbhozTbIZtir
Wyp2dslj7nkKkLaOfinM2Ccw6v5w19ZxsOu6BPBUmxI2+VyIBnJAl6HEl5jqXnN8
tGddhPK8jJHRazWJiuvQ1N2w/nyDYFVrjP9nI19PDlB30KlLMpgXwgaAg0J/nw6L
ewYQTDpTzQHTjfA45qaGkpk/bfd1XMtYhIs1tbqGhg/Z4P91AGig65Mw1Xe3rBIf
UxQKssCNdD33sMapZqcYULqMUJ9TNdzamJNiZ6elG5xDcetTz2C3kKvR9pderDSV
CJ5eKy3OQeDPoWDfdOP7iduuT4hI67W/lo2ZinnD90TjQl3t/7FAMO/4YKXpjtzq
IFn4Sda2+uLeb8B1/XhZLkAzCC+Z7Ciwi1vPB4p+R3tnDU7EhQx70mLPC3er/R2Y
5Cfhb3eYhhPQFvlr/GG7V6AAWUuhUPjiqZYgtRv60PjZ31l2lsonjG6hYj7dMZFc
FeIag6WAkibyy8hVDMQRu0nIvGW7wlESqvfK8H56dDkyxlOyMGqB0GXIUs4Yq9W5
hXvtG00VqSWNl5eTyHk1x1iLfuDM7d7ivtJ6WEpOTnDUU8lKeqnQMRq/bK8Axoh5
Qgkr7wDwAB0RnsZ/MgZsIbjhnTn3tecEIIT+TcNIrsGx54ejmeZ2/Xb9VkWCXrqr
tufZmVfZRwrJt0L4ITWJ7s0pql3VfPxw7IA6Hl1LFKkK0RwuYiox6GL+BNQnyH4E
qgrsoUj8+3WOgDJG0R4JoDym4uxLad9Sk7ysrrJP7sJn4TTFq4scd76BnLsWFpt+
BE6CTZAk17L+R4/uo0/VyywPxFyAL8UlSpRKwGRbtcqD6p5dgZRumzHR2Cj+eybm
JdArJ+PLDoSNtfiFCvxgnRSqZPgaPgjUaGoCa5ucHEydqWAEOCJMgxruJ9zoj9/3
DONFi4XVrWcXYqSDLWE0nebIjq/5Yi48sG5syO2JJdSMj66vhPo1uit3o063XPGo
nEcArs+fce20bMZV6VXilFRFi0lSBo6xJXyKzExnLc6yxE35o3ACO1lf6BA0zi8E
YH6IO1ky+56ypJyhDM2SKldDb+QUw3zzYSYwBr3qqE0eETnRDd+GL44/CV52Y+1u
O6qqmrGCVnd7mqbF++3ybhWz2X71EPZbdVZaiWgqIh1AyfMO+JhnPJEdHKk6p79X
7MLHnqjGgNG8wE95GnD7jseyBUaMHDCvgtw5Ou56AAQtS50OnGrQXuVHBg59v939
bbAbc40RZpW3nHy+5bnEcfFNVvmncxB/A5edpw7EPpfCPZ4Q25MSAN6KElhjib9m
RY5tUbgATrsV7emzrJm7HQQZX00m0oVJ6i+fQu3xd+hS7mD0Wz5+hyquvvsuoSoO
NpogTxSQv+o5ji4o185YL+eT9eViuUgYdRYb1TZ4kuhSpKbFRB/7ZiVqVbtOeSHQ
vlC27cUWFzYlawLE/QAQ4QjkfZ9oZkKB9mBceg/peSuKv2s6YHHATLMcIVUBcGoI
n7JU7nN5T1WRK4XYTAdkg4wrmEkU712riB2pDIGb0yqrpPsjC3lx3W/J7JnBqiwN
tomKsdx2BosSmWjU9XTiejeKCBP1AvRmplpZZfxJKnpNm5ahlQQpaKyNq0bSYpsQ
mcqjbzlAdQF8pgoGYMxKVZkBoMNF5Stx4qcW7VhmaHKiMWnLyAm70nYT2uPbg93H
Sq55tDR8kOB2/Q8mZnsPWsWnXjlzJZYdot7yL7W6NNx4t/uIFSHND8iALbdCOTfM
0Tn+k78QCbENcFz5OZC3lYoeL4rZ0+xrjSbMJM1RZgXZYD5XdFhR+m9AUnwnk4UW
KbGjVdMn65Dge6ypgd0ZVdq2jBuR3n6fCRRqU7ppH7b6UTiK1K/bByj36S2ccHax
BNhGIN8ByYYy3yNg6/7QM8XZ7spw7wf+sGI35a5xHDPqQwFB7j8TbXGGACmwWjuz
M7FLa4D2PE9n/4h00qOqih2GVfpAJkOMWnc+Bo2UTMevn2TPliGxGQf8IEPn/zk3
RdZMXnUb+qw2BMUgPG3zxfCoJ5ivrixn7Rw0gmvOOsvP8+7qCK4m3yJKdmJZYso4
AJFQa9CoCxkedJpvOR0qFbOC2jwOIoyHO/HME/90+mqDiJO+knabWstTXGcP5CQo
zuyK+14Gzf8GbX4XEMtg3gFfSxTXP5/Ri34KBuc2Q+5/xRjM5wYdbjhJES9bI4HW
U5NdaWzTi3sgTYi7/vkNihaleWYAIy41NYGcf8HhLzdImqE2YOpSGwDPAPjHbhY4
BEeDM/GXfd2zD0bIneTP2TslMYfUdtYrik06Ugq0x+ga5Pz57jVndgcVb7mMtXP7
eNcwOF6Ou9lYHXe+atRNBf5/q7F//JqfLjHkzareJl97XyvVo/7nw8A0szgisXMe
eFlrVYigJNI2QBxFpqPyAkiTbqt1v/TNRtL1BKg8rGEu2Aec7NDCknEewpaV/K5g
e7bbaC9CChofAj5VCvCNI3gyfU59/9tAYq+D70WBrsFfsdR+wDksZcFqPRmnF8VV
B4hJIrapV3YgU5jDJe9Q+F0yo48rNbedldxXXY2WmYYlDXFEiGzsWgmkN7iRLqva
Re9lI2+5dUD0Tru07oz5oRGtS5T+mFCG5IUZKjx7X325SQ/Mouxz3UGSSkHWZ4+e
nKO0BWlzdM/UPjmTL0Fi3xL1DGkXNk5OuFvn81cW6AdkNfLlg+88M8a4LquUkKu/
OsOSPXoriY1vC9RFBgFp7+mn4O53+7QJwLIfwEj02/xHUWCI7DAuuPu+vi2Jak2q
hSkb+4g1IselCHN/X0ucmF1lNnhVflAyK3q7XzVcqr0lwhKnoIqFkOoI1N3M8JK4
RK1ayQpo8Bon57lxTinjpN2c9mNgWyS0TnZ0SJaYDPE7cZlUsyrdenVIIICeabr6
LjhWjQ+E9dBcKqn1ERUpu9wNCJIJIstVAXPs1KGx/y49an41WbDFw9yaCyBasXSr
iFvwWX0Rz2ZYXuFBkp1dK4Bkje2qyxvTgIlSFTNrArb6EwDZhZyYk/lBmxuqQ20h
gEy7S6liDp8GrhIDjaT6jV6JDVJEh3h5kBAC1FInQfkwj5DFXdGEhQZCjaLV5DGL
Z/9HKFdwLv6f5q1tlDibRyo/T+1L00eapzPnKfWcyxU+8hUdbHWRJqFB97fwTWSm
tFbcoTV1Kmid3tDY9vsSoCE7svvWhh85Y+LUHo+MvkZoCcU4PHmvmKeHxMrr4RBc
t+Igod5poJ4j+Hh+DDxjx8yk7CZ24jgaKeua/ubQQ6ohN5qgfuoT5HpyVz4+JWiY
RRMp2gAWtJaAlKh9nIqkPZmuT0n6EczAevRT7TUV8Ypz82Nk0pO2K0gPd4GGYZdF
f7inxHzc9Z5QxKaZdbFqULGp86bzuoepoZ8ExktWJ3DHf9WkA9l6c/4tS9P0azxB
bx4qM39/AqbrZMwyq6fCRWLjkQmB/GxSFGElF1UVFqzu28AbPpwsycezjl1myOiV
TBIg8WLLyP8k8v4pZIkWYS0BFjiboKJFdE1AB6npG1To85I8kT2Jb8SVxmQ5vhv9
T6Ajat7D19ZAW+JfRtW1U2meY2OQrbmBxMDJIV0XlAG8FRBpH2rMZyc1MMu0wdpG
JtcbmYkYmZrpNtPYtDIDF1JdG6N7/6gy7Pi51n70LCaZtxF0vjT/1evcSs/8dXr5
y6vbvQwfMdqxxddV8+XRzG1DR5vLXE+xAylljEDStWO7aAsMMVhhCDNqy5CrIa/t
hlZijOn0tO9IFETT/hOEDwr3jPNISuK58aZcTlDOmsBU/2yLWV/uMLRDxXz/Jlrj
IRs7XHwn0lTJD9HdBBInLNQys1qvBF+ihgqZ3DDzEmk2UrOojTwNkJQ3ksplvC2X
sOiy60QSotYjFLH6RgbiuFaWmb8e3UgqZHikiPUZDsjmHsIFkNIndoSjCTCsDzzW
8OZfXX+anORFDFhHpNDWGap5ZHe0hG/143qmzPFJ0RlpG7YUv6UBza9VPVJlC4X7
IGPo5yFxUX5hz3LZ4DDZnzpnleL6pX7k1eYcOjiUQeTSlibl2GiNQMJxL+lBoU90
929M6BG2JOW0NlhKI0jWfXDmDVWvCCRFRIwbEpwhM+/Q8vrdUO6FoxSKEtrnUBn5
dV4T0+yIaTZn7py1OJresTKuqnjACK/Lo4isRaIQxodqTmabyrPOyCGgwc/l9X3B
76FzOzpXGfshsodEe3eC1HNRvzMB6lBeQTZiRB1sZmjoebTGQ6f4BZ5Cqm7ZwOC1
flshk9+BQPs2/jyXj1qFyeGI8NIPSc+4sPL1MWPYSgKDcG0fSK3C8dr/Z2KT5HUv
ag+toNKM7C9pIES8O6SCfAAfXUnro8Jd4aCT6JWSmUW0k+FHrgAgZEjLywh9pwV7
iokiP1h+r4gJUTilx3QZMwxW34uOQRPivGV9Vu+3x4XPdmCwcrjFLD7vadORHkUc
uQjszXeKSGX9grQinPXlG4QApeKg+cmzxCzVEC6kOtZyiZnOLBZsz1HBT7QzdLgD
UCGZSjZWiJskXExo8QPu/GoecvMKM39oSZFydIdsOS+ye4zpCi4idBc38FYOc4te
igIcllJ8m4f7fljS3CMOtryWcAuRs7VR1sDzYcL7UIyA9ZpbphFOBr4+xtadLqgM
M8GiehYYBwzPrsQtsfr8nMlfcitMQRF9V9vxobVvZi9UVkEBp7gHZsRJyXL+pXGJ
WYDffMTTwMLZ5+4Uk+sO+IY5ngdb/P7q74hk5tc9JjbyASq8fuhaJDW9AmAh8yn6
mYo5MW4NmNj3gABWXM8a1y2KoGhGmhaOPd5QK7DCUT2W7askJJYOjzpgj1kKVrti
W1wqh7lUx5y4V0Asuk1w8EFiEstq65NnXIYkLfWfAHGv5PtzS3BkZ+eh8OOUGS/r
S1P/hF4jQcO5RFBZiigjXkBSj9VQ24c/na56dIlXtBbojK4R8Zda4ps8kv2FnEsR
P/HHltOlpcq2j6gXJZ0RPmMnFit52pahMX4s3IucvTX88pW4wC9OeJh5BBlz9gte
u/fYOU2SOkcd1wsq8ambutjdYcvERdDSGRYqjPfIiGoMHgn2g5ixxC3kUDsEMxdg
sWJTOXKo616k5d7ImYmvSq3/1IceZKgrUjBEeBctooijkYJ1BHNmGlqgoZP9ZPMV
a1z2HRiC+KsPyQMswHhLbYktXumQUtG/ak+EJ9Q8RhGrJNht9IpCCUn9YiZBJBhZ
y2NBMJiI5zkc6rqozmX4PvZTVrJ0IRnDBkUR2qTM88fizSm6CHdafHx7TIdqd8CL
c3U//few/ZPdEPDhyuJqAXX3Uj+xx+D9yEpkDxKiB41/1bJVdchKJ3W4w2e+5MTB
wjW8gWFL6DxNNQegRs8rMpesDq4QhCmhxStrsgv2e3g2NSGSLDfhpRjlpmS0oOHy
XJopkaTvsKhEtd0OV8EPbvNaww+fNgN9LGQR15DV+tjTqJb8ndg9+GFEsATbTPip
ETLmaH9UVog1gNMaf1IuLiGfnxmZT03pxh9H8lQDg8L8WlBm17n1diWpXuPc5EKR
N2IU11Yf5msu87y1cRozT/yZSuR9aaXmkvs9uzFMHybQNpwFye54AR34q5K60cpR
wZ++7EsP9nygYoC9F4fRTN7Mao2YOCrTG0AzNnCTLfzwCFM7tuAa/NUeguHL3XWc
wCePXi3+/MkUx3rW4DDdb35nF6wMjjqjwn6B/smXEZDQFeDjqHqOPzZflCXVqZM+
3W1OnDieL4LklRJNg/FwZDTvVsiHJU6I2Kl3/hFaOCNb+f3cjQ+Iy/HtG5w3RaYt
XMdpMgvpRppRc5JqR000Wyr24yp1hbonhEfPJPNB2joQmmKr5gIUSsVE3EEnymZ/
N3WNdNaIGH7u2SZ/oKtX5+xkPyCpc3+jwk4zVJQKl873E785+mnj6SYMuMmhB5FB
AA5axwizy4s46lZYulWV0UeXikgiJa0nTB2xs9NsMdVWHfai+iHKA8zXQ8aYBYNU
vCKDrRh1uqKhSnTPoxxozqVu0UGvmQ5SOiTum+0ZP2rr5cjbSG/whgfWhdSLi1ip
Vv4Fd/6ae5MPe2OAetzBTz/OqDrSJE81+qakmYmIEYIYJV0BbdQugxCNnUf9nMws
nQtL68e5QFUFh+JerSASQlES8mcTT4hj3MNXWcqX6ITPZY+1YNl0NRO75axJkQTR
pH8si0TPCjUEOiASl9MjqP0vSpRviKZ2rzP0+8zQvdR67SzZK6+rRdxCZ5XRv0zr
60ARl/TcCMFSK1kUI1ydoECwmCCGgGlqKDMw9oykveGc/my+il/9exa1ryUeQALd
5eHPPSJF7ieRriFox6DKSwdVu12T/xMQRkWzsaKl4MrVGYy3O28yuvHSwGHV7J0Y
Qo7Ab439v8qt+9cPvb83B9eWK9DoA+4Oq2cqLxy0jiENbvrNQeiF8DgHSX+PZ2fS
1hy56DOU251PbAtIfy8zQfSnFya6Udn0BPegua3WR9NAXancag2CyfOw5P0Sfu+b
VAowk6HK/1ZNRkWqQyDTh9UOKoYFOKeK54832cMe1BNkZbUAw1vtop+PzkoDH96K
lu+YItHxvCheDa5qM4aySq8zAtARUkldw9r/JExsQ+VyXvS/w18jMfg6JnqRi6yr
Q/7xrQzJmi2KjZoDh1LlRj0+CSuUt2nZNMM2n6OHwHr1tJOWAanZdQp5TXZea6Qb
TXHVniTSLMMxxpX1+UQIxMnYFo4Hw7f6ww61//U7RVe+VZYZt+2JnE6ATUOX6US1
pHz3WQ6wyCMbfV8EYpZ5SZjfOG54r719Usie4Gej9XryisRxDo3pQSYt6oARItDs
40EwGIp2Lu8SjimOed7YtP9wDhaJr1YPQ2PUgptDFmRG/VYKHxLP33qIpqIjCUw3
9v+xsbDP9sJ33+NjQiV+48BHWShPsfA/cK5zzmXEtND4xr5KAJTGQUM56gCYEV27
i3NLOHxC214Wkw7WO3M1Nm25sOY6VSWfh7Y55OqPcPr1Mj7S4/Ij2FRzb9WdCIvD
FzKFiiXIE6ZNDkJssvKVFdghRIqFVqsZz5sp7UA1e8I1GNcvwogVD8PIM90Cv8XK
3xkDFkEPXydfyWjKxy8ADepsuIw4ENfIXKK8AErf/Xh/Mzto3fIBwH0EauBiUHbD
6HFk7KxVKFk490Hm/mDNsosoIjvANRx7Ge2YppN6buTzhbiiS/S060Edw4xARePC
VzqLw6yEQlEg0kPdxujOzjUjtqBylxJTuTa4LOw/pslWdFqj97uo5s/wAU7W8rAg
/vL2msdrKOgM5LfVIMjO2jyJGZeZjB1b4GNucGs1dV5/oh/ATWJ3vKMJWNBjdTf+
vsie0/T3CN6pUK2JhLH6bONNEAHsfq48ANANTvDdFJiEe/6O/YRYqXTgECB23+KC
J2Aahr6xWOPhM/ei0rrGg+KBFdDg/ZOj2oVb9pn+4zohHTjmhkcqJqFt3pyy94xZ
E0jNhVLkOe+WpJOMiqVa7dqlEXQfzj5m0iXtEqsra28ye1Tz4Hs9IOvPIkUwyj5V
r1Nl5DvadHl99dgRtV/jL0KOlZPS+C3Gx7UoNFiMfl4l8/hXdjjXQVz3i4Yvh7Ad
NSTn3L2cg9hqJ/ZfppfsLtHjv4nb/HhQmLIyMvQpKxHAjCREAfmrb7GiszC34vN8
lPvA7NKAzKhjKA0PBA4gMr1HEjQT18X89QsWpYLpVP5KcgRmNhm7EXGyf6B3mRAy
C/wOqn/s1o0zphdxD5yYCIpbuk6kfnpmqiPRwxsi6EDjFBVWTooBPi+DTYYEnEOO
yENrCtlaXQ1Qc/AgbeXvJjnAiJ9oP3HX85L6pd0xJwfpe4hwPevhomx+k3qBbpip
OTJEobPyFQbEZMxaxga/op0QnNUZ2PDSksEDTxpG7Lp97VyTe0kdCRxRRvZXIMjs
oWR0S+afIwX//wqAQz6r/3sb2hvEHwvcQEn0cfPhWyUaMQol1DufZeR1Y0M+9qs9
S8FH3vQRWWI0sRlH0uqcm2qdKwONi+doMSSKU3Wvn8xRxvXDpw3QblZxl7NhV64s
OMVagZk4KuZIQms8HgTdRt4Gw+c7iJBuG6O5qD6klYGqDdLX3ubVAwbn1ObQarZj
JatqqFBkDQK+ta66463nRDiui+f6w+WEPcQmJX1zzLVCD+EtJleFxUJZ6dBhzeBI
2UuyQ3q5Xh4XQyFuN6OuWpOOJVaha9Bjyf0JsaHo4i3tij93Sn10adiz0bti/b0N
bQT16zDFNU4adKUglnlaRtZ3CH1ZOH+i5lILeM0asjw0X6cbhbRoFKIIXoA6vC/2
5amH62gXkiatQtXpVjPRZsnqUd8Y+22uuHnymisP+rl6zzQdH/VDn9UCgLUQtmJF
9/ctPah1NKGEnwdMCxzcIuX20t8ocedwMYPOajZgNVnenTIOeQFZC5pcBgcDfzUX
5qN+j15fxpxoitrUGYqBqyLj3zFFDQPHM/FLz1TxATlf6jgh8xmHuNjUyfDoS3xO
YybVAa+MB81Brqt8/VToXxP/H4UXmdmpwXL6ACeJN9ZUrrfw7fXZaHA8oyqpU86j
GQy5SSHIU5k99b0OuHOhKUbiGGUr5vGNwc2jgxidS5a9ta8BUF3HpGmmHoXjh5Jw
SaU9qk4yKVaWFBK114Qh70zvjVN8amJydlg9cBB+1MwkAqmB06esRMDx1w4PLerq
DWR9WyXrlHv3USUz8KL4VU0nxYzv/CDVIQRJl1U6KyinsKPv1UFzEyJLcjqJUdrZ
tn/Pj3divZ8Aqp8kB/PmXkd3I2IZ6J+P2eky7jfRquUxZyv2EwdEbUt2FVvyQhGP
Ak1w0UHXhPJtfzJGknRNehIldqpaz3ylgIdDYsUL+Bm+Jfg5TZKqzzQ1cAqQEyLo
CzzvLxfNAviHG8t24OCIFNXPkta3MCnEt7a6eLgVbDpZr5yRu1UeKSobthjzASho
XEHhRvvkC/8fvfmu7nX54K00G04qlqBBQAy3gbNEYbcGgeWh+j5UoIn+BNjicWZ5
ysVqLJLc0ept1weIzoVauwperepdttFfccoUoJ+MymD0H59iuyO3OE+mC1OwkR5J
hlQPLBU/c0xc5he8P/kchoni0hAvSCS3+GkmUjKBfZFMTHFFs4fh9slQ51Co0Kvr
TJ6Jh/8zQ+419uge51jD0B2hXHXzwil2EJEcWWJFlnWxaRRRdZK67NnETCnMN+hJ
ikY5aG+5pb4q+2YNjaPnAH8NjubGs9nE5yPIDw6d6iQ1WZJZ2zzVTyMLn0rUz1zB
Ijh5t07HykvzZRV6uWv3c6zeOBK0BCLF+sFO2x3Mx22Is0sdD7BGIMofTMZXWRJb
/3DAqHWPMXhbTr1o0REVxG6XLD+A+OBCl37HbDYkitnnpLx5SH/8s9ze6l4JYKpy
6bdTArldyQlROysI8viFIUoaFuQlLBO8iJKn9cPaAGGP9GtetjfcMBHqy/HeKvqw
6GGGmm8Ys0LqoD8zRfm5lKHZ9hog7Q/064T3SeoSucMVurr01ckoqsiQHQkPFF27
+wN72XnYRmnJQCAB6fRP+uW57lP6Tohn5vHoJwejxDveGEUApt3k0rMdbESQeEus
JqpkWvzuo/gTJuLGSvDxDHidh/bMcV9wVDBQsc3Tjka/mmhDIgkcUymW4UAiJBOw
SzYTR8rhKv/ZDJNLtbO0CjYHjdCPtvm11fZxcpHzfWv/JT/1Iq967Hg0MFWZAizx
5lnAFC2HNCH3qy5fTPY2E59O5UcsVvJn6lm9Sv6RE0eGKEzRzc02nAZ4QDN5fY95
hZHne/yhVgppCiNVBvQEoXO582pvFg4tb2CGolqVD+6N+Q/MuiI79pLgDwcVc4E6
5eDFcL58UNXaO11llbY4nLYVsBit8hkHqjHJhSagQ//JmKzFu4nyFkneac+9a1Zg
h0+jN91I2Tye5qX79X7wav0TdX9aoytsvzb9AB1P+xPbBb1ifYDoDymrpSEa+fja
IFIEgqHh3uiwkVXPyIwzdY6qJ3aDo99+B24cRA/28dbwZInSGe8bb4QVfiePFHPu
UfuHKl6DEcDNH9UdrNWw0Dg2QVfZmklL0fe/6k5GlBel+1IF1rcI7+o6vNSxpZUu
i1iuBb3KFg3rAZMeNy81setF1nB4PAd0vuM2ZmYVra3UqjwmZMQZU8UfQ2Tab87L
CjQAeJw5WFOH0FIuldqR/1h/4nYh77s4UogOSJ0SdFOjl+TBBzvV9aHRJDqiIVWu
/hBiAA4lG9M7d1DwnmX8E4jUvsaww35Se9Az26ioXZHs19UX+mz0FXA7ZNlBm6D2
p2u2vHht/mcHUkoiWwyLp2o103fq9gAg6HuMPU9HhqvYWMMRIbjB5XXQbDMzDWXp
W0RF5VyKQsfx+f04HSH1j3SnIM7g0USB6/M3A0nkTE0dvgE3u6NV4RZht2BDfJL2
gImtB0ztbJ3/YWDZ564l1YY71BjbfRroDmOeJkmUnhqFRRnTapwvhhk9Axu+4b+W
RoOiNOGq3P4ENINYSTl2d7y8e2iRcS3kQbQRQkf0KUAQBIQhZtZp0zAvclNdjyTt
6kHsRuGBGw4hqYyf/gKdYuJEZ+0CkQs9rqFqM3f2XqyPVf4FljNs4E8gkahzoaGH
swzXIp3od+wDeA1sC2oeZmM08QMUDg33fQfcLc0jAR6WvaogybOhsFLDDZc+8Aqd
/CmZwvZ3G7fz5GMJuG6ook41iMh3E7R1FBVo9SAMbYAhFMD3hCS/2NL0daG+mxj5
7rM4hgMS0ZuxsybRlvbpfLIN6d27c8PWFRiQgzVMNjjtbM6kHjr1Le2m0aM+b7E7
NMj+Mx4258W3gmTTAi948tTqpuN9CkYLr5Ju9ay8o1iafSEGaIlytZHV4Q/D2vLB
TNoOGyTdy59vRyLUQpfIOjHcS5+m0ahFPQj6dcSa7I2JFZglPRqpnWTKn1JrOc1j
9BMaWVh4GtCP+Qjew905lXd417MEtGopRgM422pDk4VZU/12HFxA8mWm+E+z5mfh
0mW84TTLHvxxEa7DZeLTXY2mrXObDi4SQy7QKoYjReiMMiUhV/e4Tj4VwkUaSTxz
tGaXrVP/mKUDzsnK0tl1Sw9yepA8DSIcDFlXsoPILg+Dt9iwgbkol7Ea3zu5pY4v
exeNdcPOUjEPe6fsCtV95qqrNzeHGYzKsJHTqVhoC6ybzHtEBl05WPpcAx9O/1UY
NbNDRW81PGQ7lbhOmT4mk+VmmXtEmFmvctaXoIGN3nf8p+xSkjp3dH3jsDWm+GJn
iLvzBaOxveP2Tps7AqB18DX3Gmm+M6WSY+PM56iI3e/V+CC/7RgTLjEYH6W6haoU
D+cQ12HQWeWrHYa9VtaLmAP9S0MPPIfXG0RgptBjLYNA5O11xsIcM/DsfAaUIziG
6j9tXSZ1Drwz7NqdrMqUW9B5SY0SEZJtSJJXfxs778Ud2sgGb8kVRiL8RkkvTVwA
aFwcfwx63Te8yR33lXS6Y5adiejxVXxA4tePADNzlVJ1LTWTknhEObsbrdLebIPR
YMXGO33yB6/6i1x2NHrxonQJV6XKtUk86bNb3muz3hpWv//js5pSNnLu57Qy+nQs
aUXDxb3tJPRRDrvMAqpGiHYgLvPA/v6SEMr5eDCJ/ggsoEM281rWxGVcyIZjuom5
aMnvN4jpZ0NrvbITbNnDvnATAWyajLi5PZirEHqJff6y9WkwBH7lsJM6vJGVcOiJ
rG47+jSFwhYG2ReEVhIIE+KlERlamtqpOMkU6JCheNbxKNZ9l7Nafl93f4OJQUW8
9NcIwWDLwYlRW3TntksmRRzyfo1HGRNXJOOgjo7Sf7jFTehTylqgjhQQ0xthmeUS
lQ7sRfvrasRNS+nb+04H6KxUMbPsYZh1YeOunc1nhu8phkgqRfMRbQxAHHCbWpTX
/fIx9F1rcz+sQP6XWsweE1gfTRqBmEOWdFTR611oGhD0skXBIXtxYSkn9TsOdCQy
68tzDCaHKMTNimK6xKYQ7mSv6b4P09WxlHwia01X98BxJYZGhqiqfjCGc1kRllK0
gJDqiWKYBwaYP0vc+FtejGamOWO58tXa/shLW5yYSqvLUCjZWmBlkGHTavu/qwXU
QEEfjmbr8HZ/LRuq5wtf/ddEjKftEV/7aYi4cOHIvXCDEQnDDbU7r08M4ezvrr0I
TEN85M+O2D7Fcb4iH/ipYzDpVwxj2/3QO8BsYasXOd4bb+0BeeAqB7Yp9dkgQnNZ
z/++wJfy1Fhup+oX+st9Ad1scyOkRPpfDQ6shOPMSUy+ZlHAjc8zR0PRBqNpGJT7
R699OowV8IWnWYShmubOqnQdUqNxCMaOhnqcj7sPflwsDqdwdJMtVkqeoO+UI5h0
fQlnr5aG1t2dIFg9/cHWZ/+7QzDj98txzt4vpflnREY6ZiOnv5SixvoHqxaHPA98
D3+72GnnuDnQqku7xCbIh9kL+WMDDdIaeHrVWqNVcCBSHWvDi1r1CDLiKmN4mg/0
2FCZD5ICknfoyHD2BcEGSI2RMRlvs2dE675fn8gF0neAPR2MB6NpCz9v15/qDYXT
WDQ910HLt+f1B1miUth7BeQGy8rQJTGa7aVWFzH8BbJlh6Bbg9PhAyWvtnzIHXt0
H18BigeUiQSsAZTxbUjnRDBZ6eYmcasmYcV2Nof2zUF1FZfEN6XZS95v3wHrOM/W
1jxWTBUaY+QlMzBds+H9O8nPofj0NCKMcGskBA8MrPncj5s91a3OirNPLwtqFMEn
g/b4V7azxk5zQruSpPhQPErxUGwII1N0zPraf1C8HjsxUt4KkoDQ76SPkdmwwg+J
YZKQStot62Ewwohfzd5kOzLY5atj5nSgkCmH0DZ3KYeoDijwxEsmhnYIooHleQl4
fdn4XROKVv9kHbc+RsUo3eShNn45EEqlAwison6fTQ1494iKENwSL8e1n4sbAngy
51v4Bod76y/2iZqVWDcQLnkhvhEC0jwud1SNUIdU5a/2f1daCmVwXHt5P1byO2QS
h+iLwl2SmopFkfcWawjzdHGkXU5wVO419SpLjHdlcoQtg9E4dafah/NcIjbB4sR+
qqdRmWBgK5gNiFAzK5gir8nRf6zjPG95ys6l7rBypzPppRKMz5auckAydvOeCQvo
gNipjtv5CLdqWKANFtxv+bZKb1nacfH4tDW4ztfs5vfhhCMK3H0WdSp6GOtpP291
SipZWiJiPYn9bkf4yd2RrAIsnBxVmjI1GtmS1jUeuvd5fSc+fsG93OonIp9Axyj6
KHXUw4MOF2x6LTCloXEKC18F4nB+WHHvr9R8x4qWXxNwDRFdQcSJbkJZuDu3bx1w
rb3QCLaSpc0XxtFURW3f2S1Q1RSVLBPccspsBM3nVXkonmz89fOFGBtmQgnNNq6f
NIf2lGrcmFARNh2Stqr8zTdeNEuxtjN+c1h4AKMW1WExZcK/d8Plz7dZyaE3T7JG
K+0ZzlyNG9L0tcKnX5Purh+voc0RCBK1TMmofeGB0bY3I88cFp41BAyG6EieUPg8
qEe1AK4g4TMD8Lmo85Yfc5YD2+M4qvcNGol7cwcUKcoTiIjm+b7d43lXPlQSrvgF
2clb4ix09EZlw2hKIOyvF4AFqrccNljwsgrWeru4XGxbPnjope7n7vY1ytKNQPRR
P2qXGGxkfCSTYa31Y6X1BB1Hk6Ks7zPT5JKjSR33sbXgiFCs+/kueNQi8IfeavhD
JL+xl9TRHpKsxxnEsmnoAJlXXWOCeV+k2LFvzgpXGB+qJ/uIomyB6TzkT4nqhyXL
6S1GL1nv9wDDrh6AmIVZmKasiJeLCx0K4kbA2WZAqZ0wLV7foNzgOWukEqXip8ZD
DpZ6seOir7pCv27edYk3pKVyKN7i+DwR5XF6sIQaTWFenUSlFx0e8yrbFhCwYdAC
AX2OvIyJ8Q5FPUDc76zwg86Bo/oQkUVWOzTnegU9jVZoQkaWlAUISAu7aDdm+51G
TDGy7kYAu/BDcp410lgxiiHaX7IqUJbKNcEbacR27jphXl4toKB49fyNHy6GKGmP
Q6uJBbCHMzJYaLNfy/MU8wOUJuFh5ZWKcM5Chy+SiqFArJ8E5S+c5zMMZ0O5e1Ry
7sqKi1zsilHe4fYnwPeeI+bayGM7Fm9nuaMNnplLQ15aPmgNMHPKOyk9ddLKXEtJ
y1uLN45qMHSITuozh3x48vLXqkXxGkb2+MNVTz3Hy5/7tbU2x/ADRqtVTtxJs4K7
ZpUV82KrMAs1mncBH8rlVnKndApsNrxZr80ipM6Mb4IFr65rNpsy7elA9EvUDgPO
DTXTSwGD8f4f/cECoy37cHyjhcPc7ewFWkW0AMn6lHp7oEIUPBOwa4XJ9UVan7jW
ZM5r1aHoSk2TQnzI9PqklDJGdqADZa3OCxbWFkhhMsm6PVTlzp/KxWUyQSFbtq8w
csvZAoHb4aVdSBDFVzZAKAaiJ3JcRkze8hCmlGvvAiHH8c7Nwx3rC5ZJcIyIrBhR
gqFuPJsc38uttFnDLVff9+MiaQqchl89qerJ/MxD8VwcgQVz50AmoJzADKXruQkB
/3MeOouSa1DoqktelMAPO/d8wsA6aYyaw1YC9f8UMBX+4QPjA55ju99Y89KlcOC5
RcKmxb4/YEXhBDAq4FkRiTBCUMjz+ZF6KrYFaxtoQpDXfdZ57cmsmxNhNnWfW0Ja
NIaG9SmLB71qDbN6KcmHSj9nlNsN05dqPknSjUJpDr/X6qFU0PzZC0eIFycpudzh
CdGI01XNrur569KsScdeJa5MHM8wUIovCevhWi8ggXimDGLcOvSjqBBr0E+X1bIP
1MouDFqj8H6CCvJb1iah45nRob0LghyT4H71f/plLcDMqsyUL+L1680LwL5XpjsP
GiZvUgpR1VxDTw8iY2F4fzF7xYgdgUKWjlLgta5xfqoEvkKtWvsEtSkGSij6+UWq
tmm5nSZhRAMXDG/clUt7SesruiBzk996fsi60rVbwfMoMMI22C6owtL7JWCDqIKW
iYEOxDDZl3LISBhsELuog3U8RG5VeRIxAeH+MlZSoHAzAghvCsFzjByoWMqHRiIV
EjJFnrAyUo/Ca60PAA6LgzLszeLRL+tSK91g9ohf2OhD9UF+Bf9Yg+iaPPvQd45Q
SjluoRnL8gZO7646X4/k87KuAm2vPjwrtrVVyb8GGQHWye1BFQVeBZMrC/CbsZJ7
IST3Ez3roSMpbe62Cw/KZ7NcxrJlkQ0hO5mS4YHuC5/MpzFEFGi+P3512PYSwJGr
12NGRlK3MCFEdmBX+YGk2b4oGMMtpc5+QEfTPIlyZJceXSXG4TxI847i/VWWla/1
51bCQWBytre+aW2PJy1qdkR03IyR9fvMaqqrYn1nEMYZYjxubgK61FqsK4uYOpzq
WxUuA7mxHJxEncrKhilSzv+gOEVtmBAQZ+SB0wHAAnub0ALwYBWZvj7UXfe7R9Gg
t0dUmH6At5MEPlbDjXteZ66oMOFrYyyOWAKuvp3SWlhn9M737dqo5rG9OBlcAmcg
N/Pjy1YDlypViEztJlywVvF7P+eKieqwjgisarhoDkamjZ+CmRHRcC/qNq92X0Qn
jaHp2FpcMZFX/g9iyUb7oiueviZWabR1MkInGx3huYA0oOSsu8XEKiyVkXAleQdF
ajwKZfGKrq8xjK/gfpRJN4XPTufaOJh8YLyW+g0eNP7M99N39Ubz8JlD1TdBfC7P
t6D7uGdZkRpRGhubIRLEtB9tFtDHW6EeyyCHE5K198VZ+lnIxwR6AquE2fpPKaXh
dBLhmAHHxBNma2bfnmUDCDE8Z7b0ot/5BylHMLLHzbzFqaXCOQQBIGja9F+NRviH
9t8M/1pGk6jO0xLb515Zu4qoBWKUaGIMgDQYZ/Ql8fFc/u9CVvfKCINlJNjQSBey
DtsWDnE35vQNpM2xuV7iScERdNMg/BLNm5gzoL+K3FNOr80VrXbFa1hqti3Y0ysQ
9S0cPpR+WgB7dQD78zpwqWc88tEji2XT/yr4cpYCKs2SSPEnHsyVQlNYy/nr4cv9
oc5aUlXLzwKKTXR01jX4BGRMhqOqTPMt7c5r+0Yj1rgD4fG3MpdCOhbVSfa/bEyU
E0uMIhNYkP/40rqGcSwnErV5gOKAx0UPBfCnzlH47qAJBNMK25dL7qptAC2seHjh
hSnYLv9lojHWXzsAZ6qkduQmn/JoERGvFjezbu1CTHF/81E4OYlktaRu/at0ioFr
XT0u+zVm8DEDAx9+14KzUm/KKcgq60BivOCqgMakqDtpRvbpbSywEnxZzlIPb35P
1M4r8mLNhpDgfo239lWjS5grJBRgiLjhCbAJOLz+moSGnq60xRGkGg4j3V4tJrO/
paGaTl8HG93yaLl81od7I9QQG6+EqTEMCsU/coTALtuVStlaLnTdEhHzb59SWtP0
DPp0csXcIGSQc+rWt24JWSlMjOR23Ux4K8tDLlWpqmHe0CnkY52p4AFUDWKDFR+M
vSBUo9+1vsHFYe+1GwKXsGtr8zZLrriHO71UyVbtkq4YzbCBc48RTBTnrEl5J8r0
UlCRozV7avDHhSI8ZnljjQtmKXQypp9l/1djClJ9dIZVTmgDgTE6XjquHfGGq93X
fA236vOI+gk0DKddY1bX6RJIffvxtNRTZtLzIjTEqbyyKrOiPZhjJlTi/m0tOlOo
1OT85di//WESCbin0AwviXRR/tMEm0aidzoTZA1C/kFYH7iMxG587w8qsuZt7yvw
uqgdAlE1XozwGhYjLqV84wrFtKMam90EHqFwQ6faKeG5Sju5BDizw7kyl1QCL9iF
ohCCIuUUd4+33ZPfi4PoPLQDMscIaNkpITijfCFRmUuLUdRxo83bI1BEF8i+IUwb
Ra6mbuW5O54rEDZCd8n6mlo38vMY5NpGx1bO3mhtHzOpWCzbuWV0C7Zu07azM91/
e+0o21MCrjppMUH3nbijaU0IC5O8zRCjyltWAv+Y3CpzZCjjxPjQH4vacxdGD55V
W/+ezKLfYgKuQ4LwqVa91CODoLftuNNE3jMOWJLFK9id9MgOzQJJbEbbVzdpa8Nr
RZqy/sOOH43djp762V1L+W9qAlnTlbHG8BdW5wGP11I5JudiKxnjo5hEJCzXstXm
7kkjWe56GxL8rUHFO0YpFYxVpIp0jKXrO/ucEU7ymZrFJWVnPaCmhTnsitxwB6ed
mkR5uLIN09q09mN76hUOlI5pxluSqIrktTMOwU/mx1CYnMnQzwVvRO401r1TBx8Y
abEUYKChCxQNjNSGsZdCTJwy8oV9CWkLo+7HK1v5tPzUjPfbAtRHWOYVTr0MQFZp
ipHQ4LHs4391252MxdLxYnqDrlJupbDnuQgQHgLYAWuHsS+mlxv1PEOiST+3vEXO
XpMMlrI1EAXjuKoTv+nrBVoTdd+cEaS4PomGg/hN/7eVSFywGQ3sjzWuFkKgU+NT
UtElZVk8BcNHFzh39E1y1lL0yRvxJQ9mtQcSi86U10d49tC3M+ghlGqBtee8Fgy/
H6XNpK2Y3ssR8snk/eCjMFSik50Z3Do2IsjnPSbACHRq13ALzNOj2qWjvueVnOsU
rIBC3eY83Covsir7QQ8ehFB7Dp0h8k/IEIz+83wrIhIjlFzW2YkZ6l6bR3ioZtGU
PL4t+h3SbBJpVz58Z/LNWCKFIyFk27iwS3TwAQ90g79gSd3KcPavxAGAI2/oc+nk
6NFkwGtC/SUeH5DGkwhNj9QqnVVIn3WjvrPV5UhKDtro5ggEjk2VzJ4/d2Lavsny
cNf6kn2dtG5XAzmFYzoRVP1qE5H6k4sCKKuzGd1HNB622IZfx8qpdleDlnbvnXAa
wSUme/sAWoi6k0OSQIGuc8v7A3F3WVXUOd8gIAROVLVDJbdG+lSaxSPpBJH2uqTp
MjJvvHg1YbCYcJvjI/Nvv5VHpPof84IwbSIYaRSMWFU2TV3ey56klhzcD3peL5/P
wFleTrh8vTZG/bq5OKBp7j7NSYxDiCsEIdU/4h8CKEHiu470euE9as+HYBMp1o6/
n+aJW5uSPqjRGS1/jT7EV+WDYAzBXl4g9hBb8Sp1+nO5cixQmposLHI3nIB267SZ
PMdqTEFw7sYoJSEWTbSkm0sGqKkFAQEwRBhR27/dHoeoXbqWIwVnxgY8+8NEUSAl
nLLU5uVdmFw2s0sC6Cb2MjSeBi/U4PvueQRhbJr4+anNt72POHCfUa013n1J/LT7
rZXi+oKnzMhnAYpk/EmSsajnaq+kMjouu/3c9s9n+K323qL7eZFe/MhAHkQBZPOF
5y51BNeLOpBgH6yNhVnxkrWzphvuO6VPq6fgG5rBRmStSZrMD/4U/VHPFRNPCQ5e
mpn1HX0BMdn0Llj6ix7q6roV9u5jv0bU5awGagVSIAaotFGw85aeeY9SqRhqfDt3
nZ/rTprjPwiBR2ijC1DCmyvFJ8TSKpFGFBe6ZJAV5sfVEyLl9Bh2EvsYQaDFEK3B
76F28kWDFOyUG23P8M7z8AkAiIjT/3ICXy9jr7aZncFrU8NKrvL9NZjPvRQ5N31T
ISuYOiDqcwyIjfJB7isedoXkXhgGe9l1ZWPTpJv+axrLzvI/9zlPjAuVHq8JmuXJ
HMjebTDorlFwJTZAkfqTuIGP8KF+/ZbNSwUp1vwPGoUJawOlZt4YgTm52aRXGjsN
qr+FdFYOM8rVg44Pg3OtsARvo0id/hBHDk99mGMa534glEo09uhfa19h5kJHeLad
TOYDvhy2Iiv1ZwpO6tirX+SAuZr91mAvh0U91fczDeSVMNpBXCJoJx6c/ZscVezj
O/HLLJOns8IgkbmwdPS56P6UYxcXHPmH8b6dQPxG79g=

`pragma protect end_protected
