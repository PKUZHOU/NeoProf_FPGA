// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HnFGP8n91opRHaiU2pbpBtrkhfxRLCHMLnpTB7lZB7HP29Tco/NIWBHnm9Zm
JF/W2VzVKw14Xdk7MlQX5ACIM36HLyOXTsf+2IIrvORTmA28vGmtIFXfjYxL
8gxdrK5q3WaXZDMu+efz3LqHcF8+idec3wJ/JVBQE/1Clm1Iqcr+kdJcGpSs
5acbyEBpzzwYgRqK9C2EbBRQGBpmHlk9E+06NORRkqo/hCCHLKEmqVfwBezF
qhQtG2BuOJgGnZ9GAlNOFCgjIDNGV//wbQrKIjDQUsqLHliiNhpBSNKiTrnQ
2v9OlKTB0Kxch7gC2+mH1Ynq7zE9GVJJFmyHv+k7XQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l0eAJTplZX+OIjJSyskVziKCdxt8rRRvSJZTyTW1T30DSLQqkcdy2QNFP6NH
jaxBczGKoS5yJlF4mNMniKJo6pxZfDHgTnTIYgo+lKT2m0lpd/eWLKR+NLte
upwNMOL+x6FxhukDtC8HCo+MASel09RHlp5oMc9XlYsUvnqugZ+bUDcP92b2
IwAewmilnO1zRJdRC7N9DPkK+1PFMXSDqmplREK74edSah/uNxByX3m57bye
irjLCgDc6vzkvgokHoOmEUMySMkjZ1LBoCeZZYUxIqj5rYtfASGJcalosXgj
pTAIBgGZf7D14gajW6XU9laiCvPyVPw0d50MWC/aFQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qIAGUQQtiPzzeUIo+6rOOLN72oQgZ8sfNrMpobo8FvRPMTscHD9ZOWlY8zMS
rfNzZVzmoGpa/r1Psy90ty46bpK2/8l89w19xOacML3oTS5JbGRICKAJAEKq
lsD6Qt87kUPaXHmZ6QX1x1Tl7C4mF90CT/BABmiaMT5C1NtQBrWErcOPNZV+
0LugooVJx/nAPY36YeOdhNe5ots5fmdiF84ujGTqwRwuKESdwkOyFw07X+oS
6DUa/kiuX42GASkwed+uGm0bfCekOkI59b2OCchv0tuRuoWxub0AVEMB87Lc
/kZCsr0j9vrp530RlqzuSnQYRMKR4ONkFdpe6ONtYQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FYTRvuxE8dqSA/KKGrZWat6ydEv39HSy1iU8jyL8fhSzceNWpjglPtmYluJ8
c0UQNUU/U/E/jgIQLhhNa2xloH5PsutFeAL5E3cA1iLM8NPBVx0pW/Z1z9jf
QQX4+/xiq4RVEoPGD3IfRXvJot4GhKfutF5UTJzEqDHvDI00AaY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
WgZ9vTJNFS1iR8KU6Rw2E2r+l6AMhMbJq4dLkbNBQYn0vzyzyg/mieMSaExZ
DfJOf0yYymD2TyT1spGDIo4BX8x93jfd78If2oNweWfl1GIwsHnxvJH/LjGE
sctL8kOG3hiiAOvKPCeXzhIhUZL8e1MXQMMMHu7bQLtvh9qGEgS4P9viL2yW
eliwa5AQkDKvTqV0xVcHiSJEZx4eK1hOEufRPsnkNyH8O7NDGyV/UQXdW6dQ
5Ykvk1hZri1D38z85MJGcqQg3LnyFluwh230LpY1SNWjmhAFPd++kOpoF54k
13DUDnn2lCOCkxhY5T1cB6I3nCCIY4ZPgl5QjrNzzfuTOH0jOxUEJEu6REE+
yG9AmDLCszS+3jdiOLC7Fktp6B4d9bpXKR7Zzhb2Yt/QErb0UXCJ2YTUUKPG
0wMWF6EqgXHFLHM8x9JmvidsnWOf46dOpyqCgi4ZOXv75TVJqxPTqnW/vZAs
MJ03N7ea0KaeMU1acr1EHOY24kpMytpZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ocz/MPTA49wDMjB7OBTt+QEm5ige8M5UmDDWspwcppG/hyqZ1X2iOelb9kdA
1Cn4xH3HjlNDXwyE2DgO0VIoz2MeABQbSmJKMB9ogw52Ixu4ghpS2J6CkLZu
zEDMc+VpRe9EdhJaWiwhiYsXk8V+QnJSZ7rp86U/3fVqAxuVSE4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gw0hm3THA05eDLOE0kQyIVc44n+idBm8xXCsDFRCrm95/+b5hDTqZNV5fxgX
9ShJIaAE7KiRsx3nrqb8jd7qb6F/5VO7hUYXOdvm9njRSHXwxMa1rBNtWoMb
3iOCusaE3Lee+NMq9ooKrs98w+2vQ3vwygjrYPAI32tClXmFaBI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 37152)
`pragma protect data_block
3+FBxVXU1iUbJfjbogq++bZigkqdevkGRWXi0NAuI3vj1HD3y6829VT2PKFo
1jI20XnE9zwkhWT8C3NB7HYqSPljpiF6fT6FQ1KT77FSn7gp+HXJGoVelXjl
xC3LXZ9nc6SJKD0uI2FNySbLREncxD8WurF9EPQbdd6FuK2uopcJl1FyX9fj
T9K3/8Sm0tF680kwSPK9MhqhqpvJ2ovKWulV0vCPlVKyFSoeEaUgUF73QCwi
QnjYq/L3Ub+XcahboMgcDpslHEI2hyxtdaX6pdiY1u+g9QXTTRySEo5Z2l3T
H3dB5AbCilb7Rs1jmjFFreAqPX2mN3NndrCChLhMTVvlFUl0C0oHrIOMATMj
EVI9T/9WU4RCFZmuQ9pmJw42u8lSPZt6zM/JyfxKHEIqf/b7i2W1SuCMhEZn
j6WP01M/HEqIjsux+CTFZ7rUlC6QmXVoy9TArtXeZJ9pwKKBxABHAXA+8ViM
TgXPgTYS+P8YdBG9ZBOJpSzkM+pyw5HR8SU0zvG6UkaYlbyDEXpQBfcpTUzW
oFABZJI1ZAkW1xCwkbkb7zpie1nfQzDqnbNcm8C8SfkMrPzkG12+IhBQCpSn
QNaSE2zRP30s4mtSTlnQDLfyhiBYVzbEhldjBTxKQKAEppyjk2kguCmbAS6F
6FQJL6+FsQghXe3ltdG1ZMxptb4QFvGBV/OwpcT6JI17OV6A8sefqGMS+5kT
zBMiF8Wpy9zLZ21RVN9XAit88AGRYo924KKNakWRDhnESpDCNozf48c/rNRH
r4MtfoMNcT0pRvPqjWCrONWGb4sS69IwacFc82ZvSywXrnUFEqEzeJrtpSag
nMXrIrM0lRfV6acjMfHMMwor8STQex1D837pcizaEXfB+Utru5/04HOUAi6w
UOnWNgU6j/cABSwL81bSTSSJ7LbghWdV9HLddwIFHv/ZI0OtlS3tHiubZUjv
t+5dkKC67vmo80s518JOVM6tjC5kYNGwRy9WE6DU9TdcJVPTLqSn9L0mfu8C
NQiIvPx7Zuu4Cmp3UxuaovUb5c5AMkS/jxySKQ37Z9J29N2S78qK9BuKrGdC
OrG5WEGJO+wNQwtXeyUXr/eyCktoi68vWTMyyZUs0JnwC8MYLFvu+VyPOKte
xh35Q4BjGaz65E2koQQSpUqJfVZmtRwazXK5kQdLi9LkKgGbYo6S5nvp8IKn
aoE3m2V766LEhHbKXanaWCrIasRtZxdTQ5iwmN40JcRc0BxjeBh5uvmeKXQR
VlfuMQ2/31NaBmpEops5FCG9M1LSgMAvyeRqc+fuWsz8VpxYU26e8j4GDUIY
N9leqPShd0cp/Z3HV1CJ4xQWUxzXqk9hRwsp2YzwJ8oKNe898XwOQGPbSuFV
gXYMZ7+nvsZ8EAozNSK4XvKdRWWl/Eo/51YdJCk7NbtNG9zQ/X1Tc5Ha2zvV
Ol9NJJBQ6D9EIwZGiGnq/M/ZUMJEcNDGuQh3A8IpnNWHzUsJfzq3aCkvIFnc
V5v0Jc1/MktB3PfKo0XI8Qd2kgntwj4wRwqx6dR5sn7ArsLGSu4afKiyLwxi
9NUbTVBF5Dum66aaP9w+c+J/eQsKkT2lR4OLzKUgGsfO5g8o/+Mhad/zMsYs
T6CfgH2OPyYbtHwZt7yicrSkBIRmqqN6vAYVs+vzNhThJhjz0UAPzQq7b0Ua
mH4X/Fc52gdY5FpTu+xdtIo2hVJN3eFczbLQuPBfesGPqNj2fnU08p6OLXSD
0kRwpcabxljHRHZCNJyiRzcJHAW0mJKEte2d6H8ZTij0DwPE/kQqxrM+pF7P
tf2NGcQwOeQovA1Fhdg3iyDE1bKsBjNuRCLgM8nIAnmVs5Kfj+SGty+YnCs2
cXQCi8x2+b6fHJa4hRHfRglAYTLZoBcrpv+/JJYGD+ovY7KROOeaK+IcgdrD
bjuOD4uG0+LEu+uCcpwKCkYE/JEEmm2ge5xSKCB/j/8L0p7w+c5fnW0BeKnS
w7wKLv0G+ytTDRbD7p5zrfgaXWgtX+YNv6fF0CvExd2GldTYPUbj+zJmsE3Q
+3En+O312XEFYstCeI8h3ZsEoZjgsOG7CBtAm3J37bGvDAISVdgECA/0MJ0e
qWJ6Rk7y8hqy/fVEjywv6dMfQxKTTwKoDWDLyNUqhfJvpBGLAOKBily/JqSa
14JtWH+IDtjdbQ9A7l57gBK8oFJR2IvTOYKZSLQENhxxg8FNOOBLzJfvRXyr
Sz+lQTnFlJ3a9FNL2LVr8bPa6aKY4a9ee6tUDU03my0zIDViWMiWLQ216kgT
5qdbzLvPCmwZv2Nb3AEBa1CJxxBuVZgduR+3kNyPDeM7Sb8gueswd+P3xehU
1nZkaA+CqjlOXVw69pjVZ5AElWmxo9TDT39HRWRyRjdXUupkiocnKkmucTGY
9ayUcRodC01f5dHFjp24cKWwU2YPulVmVfYFBo95/fn0ABBrt/KB1U8spI0A
BrzCPFlSiykJ/RP2nFsNCo4abgQap+z+YPWT6LBQ1dMjAeEN19mL4x4lgKPY
cBpUJgtYzPgbFnVPimOT44OwIoyWHZALOUi98WSvx55LZONR8r9vXcKzSl8f
cYGsnPpa1WC+6Agrh++pAb0txGLf6dZkmqCeoIRag+8YqhKj0yMt7eXLsR77
NzGZVfrNUnD7StJ3d6yVzLWYTPNagAlEVEMibqYxRSpaCTboqoUeHyc+p59S
/kYSkHGL1L99H/KlrrSc9Zj0IWYkC98N5NdwMq0wPW7q3nz16Iw64LKks6Cd
zbGiJ61yYilX18asDuP8nti/AZxw3x7JmOqsjJf1oF4H/YW+yk2PoCSf4Dd1
/Q1N0wWaw/SCwKo6qp7N1VLybBeH3D+KmfgdvcYe3I5imXnycEpgyldEPNH4
dJx5Gs5m0/dJL905NB+53q5NPuCTHf95LyY522tzU+Bo/FGdzwIqOmWHcBNf
FUICb32R8s0nmwzpdFxzCswuaO4YrgfHYv7+ArrGwEHCKDpedQGZ0yHKKwlo
jS4fzDPnS1QfcWmtqymq+cFablgKEAhppoCBseQdzdAGY2mKqGW6k9749yLZ
eTz5bZoR2eub2nm44gwi4G9Vpz4QhS3EPGawN4Bsk8e/T+XksiNDQmeFVziP
bcQeKng76jmrEFa1pAEib6O0I4niCP9b6gDw75NG1RXGhwf/I8QWilp+eGZv
NskJvporYX+p0g7fQjaZDKouaDjh0VRDXZx6uuOc75WcfxL1W3F7VUu1HtZc
V4rosdDpL4ePLZgs5d2Zh9X4R3051Yh7Jn1GNeczvpijMu3yqDPm+DAd5K/K
xKH9zeAsPuYOS7D2wXxaFYGoj1mCdT9iZZLaRgX7BsJHbYSr5qNijQlehilQ
n6OFWqxVh6pMXLcOUa4UItJaai8zbTJyudpNVswKDpFdBFOsMExz7jP+Cycz
Dq0xDzqtkLvxliFSzyBxBD+d0SyvodscJ924q37bflh7+7YlDT2R6aZFvfpT
xPpvweYuEiGxN7EAPdlUDSzxs9213uMpd9INBvIEaiejEyK8j5BvNTNcRT34
cEcq8Eh3JB+cu7FwEiAef1n9jCuL8gla5kHNItrNlwspEZGm3o/g/dp9g21F
RkxF2tl2+TRknPidh4Zk75BrorZNXq9slyKUBwYOD1voTCe0DUzt/SjQKiC1
P4YAjOnzmn09Dx03rakkpjVXNnpAHeg81t1vmY6j/5bMaZri9q2ppKxE4afZ
tw1IY8wyiQda2ayz74Nbex+WLwCeohSNXdnBfmQVjyNdnSLVnZfFxF3fXXiC
CEUv9klbQy9yJeNaQHy4p08+t7l51XHLZxTjLCfXNDcQZ1H+UfMKVULgyt5j
FLHjKIgiD9r41GXxIc2mh4+SX3XEFmn2Qzw3lOScNnABjC7VqObNTgSSqAEe
5sdTylPWHKz24Wxt0uEAKN5My4rXoPCQeJ7jfUv8qCqwAErYizotdgvfEKCk
V65qkS9KdbE1DYhVMx7sahdFxRGu95mVyxMt8TGuPfiM7PzraGFdhGC7uDef
qABr3C1UfJSHd2vtbTJ8uTmmlt+P1PFrm3h0jtL0j6kbMp7dql+EU6HJBqV8
sT5Mq3mcDlTuOYo26uGj34mXLWX6mj0ic/rVRYZFHbqrd7zKxUslGeWm2asL
KcsrhEYmMNXcutVcx8umN3uMR/qIo52LeDHD3yJVbbJ0RHL4/k5Au5Zrlppm
5VQoCndZP2U2UJAf+4fAziPG5W5sKP8+NxW+4I40hKfHMQAzDzV2SSnnjMUp
Af8bk9XQbIR5wdHmDsE+nkSiVQDt8r0EDcVy6QKokLEDEMO+I0VAE0uI/Xqf
3u9wC+ly7fvEG6fZbs63elJ8SaLryuftWVumgc4rRr5cuiqvmSLSWSkgCB8H
Q5qYtd4UZC9SUyqQgyiDjBc5Xq2yt5k570F4e3BN2dn8l8ejq5NcveHLS8+I
T9BC4XJKJtdnkhFq3/z0umHWkkIsH8bUyoKPOVsZXQGypwJeoLQa+9k4QIOM
SSIamVTEiSlQlTdTm7y4Wo7Btc9EhoTXLFhpBgGpxarcQFI7L5YS6I2WmSrt
GCsoQiyY0XVsMeClF26Jmkdfr53fFk3pU/99KpXmGk2YwwZqK69L7lGAB4Sl
2X13pt8DifvYXjSBl7BZT8LeyZ7aA/7DXOVHcfIQ5xoNoAUk7P1etxBY5iHh
Xr/hE+zGRaR2ePB1Q2NMkf92ZS/TsB7Be6r7KS7UfzD/ncQNT3eedkNTHqcH
8TVI6IC60UNNHgtCT3DlEq7VkD2/ZwfnPAv5k1qwj0TubNObkexFwMH0OGgM
GCZIcLLw6sGyihMDzCUTEvZcWQQutSdBxexMh3xuPOs06spSeTD6YNH9E7Rv
Dd8qQGUMhefDYJKoWM1Mbk7kd3uHz8eueoBnm6Ffk1WEyxqv2ZHA17xUSv5l
9KT/LdiEWN/bd8GP26a5QV56uo2GnmrRyMhl6H1XAo30BjjS2Fo0OYNskDio
YWheYAT3CAYzlhAhyTZEJ10F+wFrJ/NDcdD5IDHeOcfiG4HqG+8MZyL5gf0V
PeEf/bJnu7ZxkpJhTOHdljAGHEGrxJdDzlv1PuVO3z7I6sfz5be1MTSS7pGm
0Kug9tO8P74ek9qm2GZoNrI4mwSbed008b7UsvsZnCLe3hdyxMlDJK45sqW4
/H/XBIn8AZGNILna8/zDsYO5KiSGNqDjTsP3qQV2hv2Jhvqk3skJi9+PIzAY
6nlvFsYz6hrOnPI/zQmJgv9PcLp1zNQ/g6n4X18ZwKs+wMgq9SYE597HRpYc
5EH6PXldO3MYYGoQ51EUsYa9IYbKSEMo0lqJd54/bcbaD3s+VS+W26sRoTKv
uLhpHCFaE1zRaRK6TJZSu9bvQLITXfob+bc04liq6h0y1PV+FgqmjJjsKLGe
yw4WPeyZQgIpBraWf6jP2AxrjGa2oVI0M1/QzNDeub87iOfQ9HxQdzlGtxEx
tcLGmTTL2/6tqh+1lWVZylfqzprYcDrKPIqshmfP6ng2g8fEGdOK+QToz8CW
Lj5matoVDEL63OGx/UIT6vrA5CzhkVfBxOuxnifDF5+B82NM1in1J+mJkadg
zxkyCIxCWS77OiCoW8F2aSiKVzuZ2fFJ4HyWPP6qXpi3N/arfLHmTsVCOPfD
dGnDxtbDcCltmmWvwpsKsMzbAU7o6ekvFrl9z6KVpy4zpyd5KKSJL3RqFO7e
TK4EoUOQEGYLq8mxCB5mMQeIkvyJjgrM1LwVvS2X7LG2lHcmEw/GS2XmoxCm
Lkgr3ipal562r0oFYKfr+IjKSztz7LpuLkQ03eO5aeWC2sq4phcipWI38z3e
vwfbpb3ee216nAzvB/nGmdKfdo35KXXdRc66zheNtL05xBtqMbTLowi5rqnG
Cx/p/xwawM1zjwGjXatGLdD0Gm+5s6gUTiqFoiNjlZtR9L68wPC8bdM8oizG
+K/HnOOkg+foARK6q8K5FHc4DfmGZ8Vcegydb9yEEsWG8mR85N9Cesh5kU1P
tA3o1NxtP5UrxoLqS/OzvFyr5u4fJ/wHtlSbEXWlgP6qP8V1QoQ4++JAjcfY
bkCazGZ4kULoR3pIdRrxXBywjX21n8eRZdbU3h3C9tlWzJlQNiFZwYGqV25n
3b6yrE6gHf2kLbkj4Vcdf9H63liWI/H/5XJJx2RyNpuqywX2doyabc2S+YF/
afbDamzRNxJ/ygSRcs2ih2Mhp0DOKQSGAtxrNw2bP6/a46jhiPOlI/M+3Y4e
yHRiBUyw+Jdx78mLTyzJFkuguw4dUkjTSu03fvIX/dDCu2/F5YHngtY1Dswq
OP4s8uGk1QTE/JEgOuZB6mNPBxiOCruSxeTgfPqoOHu2LDTmXHUuXAZFkTvQ
ajMdt4ZMRzD9vtoI2085cV4uSD/E6ISGZGC2jB7jKzCD024RHkBgoRZ4hXmj
P1djsHkkrK9kBsYZd0id4CkyBRxipQUZM4G6sc8Huckh3L6sjaTx+3IXCgta
xw0jPMDdLO5oCC0X168Ehmv+l0SvkNqSjoyY9vMFX9tejWGK34/IiTMSPCGt
+chLf92VTbI964TSBUdglJqdoE+srPx99JJO+VV++BXzAM62ZWjH/sf2u0rO
l6rDa0e2yROhjPH8I4d6mz/ucl3zFDqq9lUDVS4TDjIPv3DZdbzDTYlY0/w9
O0vGcUjen9+t/7Bq4LvMb/L11JH/ntQpngqFkN1MXGVxPc0DHZZpr1IYv6Ol
y9sliqFx34kl+3YYxaoy+W5xOO5Oex6vlJqNEkIqk1IZwEIiK7HVYMlyzyjE
tQa1BXxtZjGZ6AVc6qzwcJJ6DwIsoNinsUoQ1wX20Jg/PAxfB+RR+MtJRKWQ
aJSOBbQorkWyc/WtZ7u8ZGANdrNDF8AdCw1BKZzDnV+rUZtXIYSH7H8X11md
p/WJj1EIETsVcOAzfPJNY2+S3W+RWPC2ZprXc+mhVMFhBDDve3Kk5HJaGRkm
i5hnTGsUYd9C9vckud3VTbUisVzMqn1W0nywkDslzKhqqU1oXZDh8RzL8/Sb
cQcb5fEJCIVPbTmxMHkbPZMxkP7f2In7RR/OCavne6N6PqXbO8ZO4aqtxrTa
lVSs7eWxpEst9VpcMqRfNiGeN9QpOXAulWx5P5YruxeqDo5aq5le4gyvkBwd
i2wtMZAE7IkTaAbjf+5EP0+4yg+Bcc5DRZgGcQ4PJSGn4EFqRmBMv1+Y6b/4
DDfemz07alc2tYgm7gDfp19nMrGySIIDLPMTKctRPvuFu23GkcWbhzWQFB9l
lkP4FGkdujaDl+il9c/8mkKwk0OPyeQZQRK61U6hp8RCETh33qH1epVbaZcV
L1QYhjPiddnNYQALhptA5a2qRLjvi0/MQvFDxziB7qt6oBPzPi4DHK/fR2gi
0naq7hRpRcK7Jyk1L3RRU3BEFfgz8umaWCM+k5x9w44e3qJnaQhsNtOhhYXR
8CpQgOn0TEhtqW6Yq/SrJ6h5ivf+so8PxuVhj6Ed4N3ZwJlrkHTH38srx65C
W8eJd1E2/gXwjxB37uWLHrwWGQ+zAsr/qRlLdyow+IiIipiMEFZNEQZ8e7BV
jUkMGsF0UsyMh5En9uGKZAw3E44h3Zy79Ba51x3MoAmvezuarhXLn0GHWsnQ
x3Pyk4BbrsFwQTXl6bVjmWg6RKg2ME22Y5v/YBQwCD5vNEHH8ezwxgzhVGI2
W76EQTWYswYrd8lWghMhNULrCCLdEU9ZuEgkWWBjlEYJl8zWBFnpJxYGSG6J
9jlqXTvLfuSeozTY7WGcWjwHk04A1MspX3fIaVI3cSH//3Mbk3bHmz30WKR6
wxYvTVjRz5rXy1q1rjBr5N7H5RApGKcunvRx72rBAwJCHL1cneImmCEHsBGG
MVia0xr7YHh7/OvAsFidOL1XavhTMRFzaUOMbMueVzPna0r/1LPiJsgXqFKC
OuWMz4dh05oPkoQuLrWUrOQLD7gOvUsFCz6Ao5E206uzXNpsHLZW0ITNII/s
7qcGIhgskyxGGH8sqLAF+p72ijbtsAi0qRVr/AtWFjCQVldJ6y3BHPzPLtPR
8/uRfHsYG8Z/obcfsHQju8fqsOdlfoKSxratgwIT9GMB95D7Gt8/ldmOV+4j
T2dM5aeYTyDPs61Cgklw68pM4gBB4jHdFZ36sGu1vUQ78BNlEvnWj2FRCuN2
c6uX1LbLuA2wl2ZQEJ4PbGFsfbJDs+KSESZAb75iO7UkdYlXmrsweJSVE12f
wiDLHIT/z8t10vn1HpYNPRNY0eSjUXNCFxiw6EkZ6HyrJyjEt64cT4KL/doO
t1o8WvYuUMwMR0svp6ocGAoBWNGPOOwbwelGOu51+Kk+pTcpFUS9aSLbFhvQ
Cv4jjW84+Ay73WZj6lnG4MJd7/FbX7J2IFBm0ihjp76TnZKT610A/ARfhDXj
QHv9f5AkIJPQr+9FuRdrSESMCQNwiqtBUlS/yOBLCeLRkEV3NsMAzgrVq0YV
wMpU4EKdB+HqDngs8o1BjQ6Os1HzOzf2ls918ugMZLLaa6V3uh+CUiQc64TU
kV9K4+1Qxvml6zpcTGDrfXPYALip30YiqkMVIfHESM/awW0OCCxRoAfjZVIB
VFpf8LogLzjDQNX+AAxvGJ/S8i/jrbY93iWJbsMg5S+4rpEKlEqviL1sQUhs
QIlaxUrf3+bNRg2IWWljo2T0md4RfHG53TWCzcExyyg5JkAnqONw0icjqcXh
hd9x2lw9rNzjaIaDyYaA5iALVpPpDHv1IcjpEO1HYgEFZGzShJncgW1NKlrY
P+rj0Kw5D1uF8Zepx4iVaSI6OKPyorKn6pQUT74HVEy/MjXi2MnGw01Jz9og
3MU2xeuBU+9aKBEDIEKSvwYTw2j5yhp8iDCM23gMaXeZ8QeDBPr8vJBBavpP
+QqK+pwbp6b+c1i6H17VkmlgGn5qc/WcgO1C0lntY7nJ5yIC1+K/RrBFjQkt
5yyC+CXfSpaucGYZZQJGwC6tTzC0/rbEN/xSKQt++idpjMsFxu9CIEfJYxJH
jZfvQWpt2AueKYxq8xNOuThzs+f7JyGF676hTfqVlbN9boDsTRkP7Jq5cEW3
BKYVZRkmi52SJldnTJ3qvkbXrTdbPqB/3H84fOEkB7DkvmwrXClVAsu9XNrK
qP/sZ8q9FJ9wBH6qrKpOSl8RsZPbkFSE4MK+CYFWiBzQhQ/aTkYqqFWrLgKZ
bkIuPKGjoc7L/cqdje/duLA4JmSEfZzPATN6P3NyM1MkIM13Z+cYkoWZ2M22
0V8gWYCU/SSMH2ZRKQCNo4PnQK52NMESvmX9t420+NsE/+DW9xIc9KMACqU3
KOXN0fNgaQq/cd1CVWxGL4aGGBxelySaqgqO9dLV/Iz3FTqM+xFw95pqngsJ
A03eAUIK+qsvn9LvsvgOw6ZZ2RU3Qh54jhWHZIV3ndLDJs2gfTn8L9rDzYe2
vzf0zH8MDizi9CaHpW8itGJZssILxh8CVWCq4Rl5a0lKK1xh4fOYcpbQ0OeO
Za9ZOxtBJLGd9eAE1DGKeBy5oPvXY5D70q5YQD0SOuTUcOzjCC0WX5D8f5tV
1ZZhBVWw/32OoHskyucFq2U21lkKTRH8pM1CVPkubbZOScNk1pVDTQHmstl2
PXqHN6AFdune9wVUnzpgr4eaH5m2She+XsySjKbkhUMAr3VXG9fMJnH4qKa/
WmnhFJVBSrTzCdUIBIUJstnuyngQhAXMAB/+d9Hrg7SGOqv5bnDTomuNMIjl
houQKTUTECup9IVqel3+/UeiCl9tdlKYLQXXE42KIvskNsuZ2U1b3DyAaoA6
py+LXaqvWfADAIF5wUSdw+eSgFGlm8dqRJDijKxa2l8ZpwYn5NuP9Ou1d1xN
S16nJWfrwW8sgfnnnZE9ILYsryNi42FWXgOKbt7w8THXgT71kpMQpSSl5S5L
x1JUaC9QqciKffeFh6Ch3qSiK/pinZQlfPAzP8HoaNMkQYvUdQzl4FKmKuCL
eK5qLfW2sHJ4rqfz06Y7iaFBxGgLr7t4ckedVOLmFJ/vUJvjZlPuscmTUq7I
3L+QKj3V8296C3DYQ48fGoXMCKDeHKN5pCJFulcNxIrlPKQ5Ttb2sOfq3xkn
A06yEIxmluUdMEp8VWLgSclA57d6kHOdK+S0Xv9bEg0jiwLdyte455oMjFVU
Gn5pbcHA7eSlh9uB/esD1J+nnJ62EhwnohOV4PLhPuqHu7+XPrRK4/O3T2yF
u5LFW9BG7H8GW5+RNsjja5swaGM05X8WihUlnLE6G89vX4brzsk01XtTOYki
7eYAakj6iQMk3sPkFi4fkFKQ1crwByLeeZeVOkm4kuJcmwakOX/Mw4alXP4X
FFR73O9jhUQ5UI2DN3Z0eIANPpxPyHvngpXVWhifIpKPbhoA0zN83BX2xZIh
mkZ+byS5P4zDf7fZKiba/EK8sqXYrF0BSx+60eTLZvRuJI+6Ul5rSfMFvQB8
gRSteQREGC4ZAKDVzIeaw6Fa0BK/KenOYBccnwaDO7ynwee5ZcXC9uxKX7M9
rkat4idWadjq6MrhQ4tzNMof8ugcJkXgwgOAd5O4YFL3Re4hjR37DvjtfBMB
7N346+UUiPAAjY03t8Y+ESKTZmwH4/D1pFCYNwL78QDYApShKu4DUIRkCJHg
PwRBx7fhDtWcAEFUsgAGb9K4j0x4aRZXGE7tDiErL5ykShBQqR1EjU4ze8In
9RufUBn8C44uM30/MbGqyXsYSvKkPP238ySF+CmA0zWTQ600EPySc/kyMYJk
lGLmLvrJw58ZTAkGxpb2KqZd9Vw0+abMvVthN/bnbAeJB5yeYGewNBiDoxS/
xgQf9mDfc3uaMCU9+/osSj64UNJpe7f1DFCuSjvkdhmci0wUdhdurGfuaMWW
J2YTn6jiicCe2d1iAuOesgUtNuLoP30DyyLebnG2FUGgE4rIHuQyGtRwCGFH
MVpXzmXykS8Lp1gYAj7uNeuukDPWENjWnufiqB6+LH5XwqLpj8p4jcZQHchw
JBnpR5Sdjr09TaZSsOAcz0jfGqQ8n//RtXr4DmIJ5VGvJLbgPda7JXbKlftt
tzDGUft4dVKStmjOOHE4kYOUwDBBujf3qKEqLNy2B4ZQL7SxqhY2rymrJZz0
aQoYmwy6ybyhsNSojgbGcxhVOn4mBpkTOfI13vjtOOHqRh/bdmKc2liOKgmj
RJ+1bentzing0ZqiEEJ1QV27jVZH9tXOU/q31sPiAQrhNHhwx8RjiIFt6tpG
TEK1FSG8lNx08KeOzvUG0qmlgQti3kKOCIkgVwDAvUEJGv/jA/m5wK3pIpQB
Cz4RUa7W3YS/GM39cYICUWyvv4m+aQqyMG0iEZ+Ck9xyeBxHQSsswY80fvTn
fl+Z4XHRGzjrXD/hynyZJUbF6MbUni1cJ4JUGNNELaS+IOhMqyDRryuHYp36
Z3dnGN5QTfI1JX12UpaFGRZt68/tr0mLeaI1YFxobgkOVhspYCoxqIW3UgI/
ZXA214HR8q44++1LlqNSjzHLt4ympTeGlOpM01EAl1X0KEaB7O6YT6ODA1kr
lrVQHPDthbBW8MoxdVihqLxr1jRc+FOggnUNAaZmLSNCKH8W3w4pm++wRpag
LG3mwWtgbP1542+BO+xQXDLa6SyaY3CTHNu4HwAP5awt4DqDje+cq4XRLMUp
dpMM6YgXtM0AR+wZe4f6x4//fB4igELRd90LBw7th8N3NYxODpbiOPAIwdJh
D5Nhw7NVbVXbZVAkwlKmrvEXUQVzZSW5VgeUYsfVQuBJnJmHMWKm5q3Lw/Jh
EMuOrlfYa2JogIy2yd2aFaEEZqRUYzLNprWk1pRFaGi11cKQOqfMH+fUNT5X
LneYPkhfhUaisyVwMe02ad4fmmmAmZtSeFyvOwGbs3jQD6CV6Uz6EZhNtFqx
XZCA9YXThaW91uRyN3LJHHqijC8ihxASqSQIn5VUTWPniNDWySt9k0fXzeax
087neYGX/Kl0J6r9v0NnYatYPQdG/DU2f29RdRvRHzsSqIK1kuXGggk9odJT
3GkrEvSqaMcfnvQYZJk9tNkGSQAMSF9/5r8U2r6GMoM+bxtnhpCoi3VsX1kg
Ie+X0lW77p7MEIwqP10N1rUXtVfJycO5JHnNwB1DVBE2v1lxJbom8VR1Ls8P
ihCA96a+iIHB9z2jcDDMZgOHFdu0n7y3hNr8+kRKAd7212t2GJKUiO0n81Td
qJDc2N1862Dz+0DMPldcwd1ZDR7JmjgOYaDfEb/ttZjHaBxb9Dx5bJOWgcyW
Fd5QZlP2Nu/lnPI+zbPlYe/pyvrh8IH3VLovJKml7hCAOtg0ESguwGErQ3HI
mgmN/uK3e3qNtqWmCRxb8ZLCov2psswfuqIrMSOglD6HEIS1KuK02tM15yO0
eigjhya/kvztinIls+hRCaNmEZazl0SWNvMAe2YiQiPYk4l35h0QsPSXAdMh
R2nDB72PCya3OL2I84jMUCewdZFSC4CAhIJqIqKznaAJu1AksySwlA8jYveZ
8ti6uBe8ZeGTNfr6Druxg+nWQhsiOBK9SCgA4yvANGRom3PgDZGjUcVDxwpg
E4MJ699tKKGTcBsPk0MUtvIokVWo2zQeeOrtRQwyWmxPeJwQebKxW3NbzBBu
EmKLPGjef7D3xtp5W/q4DL1yuRFtFREXZMKFKD7wuf1l0O7+V2z8d0mDMMSH
U7xFVA+bnbFGQM7vbnXXAIFqHwZdjsMJxzdvo8mN3BCj9PktTvw8uyIrFsi1
mYrfXIKvSSIprWPZz1YRrT00iYp8kD3kUN/Py9fSCQOJo6noW1twabcYFAnJ
QUb86oEpiiDc/jnLxLQIawkh/XrUGcDnLltGV4YUvWpxlIa79dVXpyY5GhGg
QyvEHLBUd1GcEKEO3baKhNr9kH5Lsh3NidHj3ll+XuFpljwKQaLlbGYCyu3W
q8B5CztFiWI1dTd9u5zO2NwioyGDWOpbInc6+MX0n5AGcqORWBEeJ8GLqiSH
y37v5l3j+5WT/bqzSK2crQQoTJTph92kTcgboLhvehN4gR1MBIqKECV54/sq
k8hBXO/2MmHN8e4gvr0VH6h7abfTmefwZ3WU1Tcpk3/OW+r7t4sO81C7YpNS
kPC6OKRBh2Inq7pSNRT9aNWIe15OmVSUhfaGly/hdJajI2zDaPpjIl0kfslf
9eHNu7cB4vU0fAXxZwxTpSq0GcvZ6D3cYsP0iGShZRinMs7CAMaxapfwwltO
kHbuGDM2gOCIzULkqHVLX8FPE4YNF4e/UfMNgdcGpxK0nYmfEhZduV0GEAJw
cJkb9b2mLUo2cukFLliYr3jse8t/WviYfIjZk9XmKVT7dMJCiF53oTLFECR2
9LwNSmVkq6u6xB4DiOMTO9oXWGIvCPTofoy/f27V9RUK7E26ubjDSBTqp9jC
EH/sdsDg+cSJ/7hG8yR6xAlco7UByopCQpcpypowT9VZwd5DMnXoPFE09n1L
htHdjbGIyzIacSS9xKc7ouvL06Gui/aTMnFiT4e3uWJoTXhrYJOX7NNnUunx
odVGJVvRUZgcErRIOvEDRHhZ9GVPKaJzcXETBUjSCK3JBjlmhU0Q+cOEFUQb
dJnH8BmahEQ7t22hEGzfgdP2olYci4MmoOtzUXWflYZWoPXorGwiJ4/i7oHs
QfyCiJasTK7kmIVl0gN0/12WTT7QrPFOdGaSzT9o0VbPwqrQ3OarGF2Im9aC
4rlf+chgjI082PzlM0nysSZBYpeJJnRCmjRTDmjQjrM4C3hDV3dZEu4yL1L4
2TtBtR83GPYblDp+6giFWdgPlKiFQl+FoP6YuYK/L4YVmcSdQUT5DavYaDl0
xcr1mGCVv/HARpW0hPZBmLttahF08wQ69AEDLiVnCjrirwysD74GMCCmzwnp
3Hxh90pzS/t77mABRIVtiGGv/FmE49in3vmyXt0vGLnEuptC1emaXW1ycCMf
z3/JqGXZddZg8vprYGizQF2dDQNOSlT3yA9GJa7jjnQbPJ1H6Q/6HCrsyTN7
h8eZkRH6WYiO9AlQR9yqVtqEfQCJd5cATxeTkThS6dHG0IiB6ERWckB6kKTM
fiBX7kkOznDYWiCMC98FbIupvR2FSr7AlVmLTr8g2RkZ3e2U1gjpHkriPYxp
pKDOVuXVUkuDDx+AXpOQuCaE75cNnLP1o1uq1UhLoVd+9HRZghAi4CMYz/fy
EBf04QN2sVHabrtihAJG8MyKlmH2MteELNEHPNJOPvkxhpw9tQHJj+ObTf8j
DrNlNe9gFc2DK6LoBtKIGHiab1fBVYisqo6ZaOldiTxu5cqhj2Jjp9oearwA
NhIy8dfmPfuSPHgxRtElxm6EKjyHw/1cUpMTYa6EyEi6M1TFloCQxGG9r0LO
wVO3mAhzSLtPnWbu6jn/Vo5Q9F65V2kxT9RSFrA+Tf3i2BgBP0M9KqlgOcNR
vo1Hg1XwubAUrRsLHhmauSYzQawziO+bhiiVoQ2a/ZvGVL8ll10p/Oz6EBeU
5IbmQACkzzR0Szaw5Alm3sp4J8pQCkOLwrVZ77deQxUWlrLJSn6cLzyu7Iye
RYmXaGhibDUoWUdndEnTraUV7rJXCc0iOv2WLUMej1Y0jU29KYmW1AaPuAkd
PK/q31XJKBwDpywzo2KxWOVGii72KZZjpV8d/CqvZioqApo+qS0btqsFixRE
Hvf0qq33hdXii1wQDuhX5Ax54sBGQjqx6DLRpmVOSVC96XXojOBKSaUBsEA+
GKqqAzb4RG9Q7lwH4K7nr5DL7GFnzxz3SIybLvhJCpONWlc4ghfl6Q+3t3ma
LEzYJOTCpF4PxtWMLlc68cbedF636jcHMQ4MiX0lakVAhG8RZM2QK5EXJsPg
MskO5Bb9rc3KNzJwHyTgglC1qfhYZnPcSm7DN2FQIhZN29ObuWI1CRbMEuVW
JWFTfS+td12YsceT9kCFpOee2aR45/+zV5nvzR5T3EfhPvaiBrf5+2jZq+mo
9ikZwGMrkbyYmnBRnyoYDGs4lsnfBwse2OeoO1qcF3ZyneymKaoK//BND2EV
MNsIOuWorD4O0KClGbU7wEW/DAERrEhi1KkQuvu8mOG6gcE801gQUhLSkGF7
qG+5m2I7brMxCQRO4yGXlaAmWuadIuDWqRKthi2RQwrprdK24Mwsp8npStqF
OAxYEpbPFTBu9Hjo1J6daMvKPp2hjZ+EyL9ceMySCO4ZqT2TLTY+X8MdfoA0
gODiZtJ2Fob2mNstEy0swSmFLlixo1rEfQAkLbM+8CeUewmjfs4fHfD5Ur2p
97PsNE0Y1Up/RHnFwfYAI6K9JQKeMCNk8sC1ZX4unok88SP+EbzAw+JrxFGt
XqyldByGoDzBJh95b9aZfOa7xaU3BunlNidoVbS2S5p478EWLdWFobpVff0J
7xsrEoTeCyCdfl4f8bRRUWRGQTtxMH5GBIlFmuW/w+lCWFiI6cbQCEGvkxqG
RMk1VzbpOlmzRV1Wm2U3tKDJXJP0xsfxj1f7QlsHEq0oE5s6Fm9NthAqjWVH
2wKDg4K4A/v2YniC59heVwccHZ5Bi1kSzWLobE9b+ZT3Wcs9NZZ0Nw6oIIr6
NtT5Azh4skcfe1kYgh6hXh7+LO1Tr9uOVGJZzmXSHYJYjAggKn/SBiiZWCMy
OHtnRRPPHsrTWrtYQL8PZGkVtQ6gnKa3c27B2moVoObCjaEAfij89o9ASRBK
SlW+wjKyl5X7ej7UnRMCT01t2c//pFYjRDxUzbYz3kbt/0RLvmcxcqAPU/zG
GJ1oIy1OdW+D7OpnJ/bDed5F0jxOmoym8hNbeETQqX8cdHzRNcTkbchPwkW7
+9bfVbl4JGwxJjFLT/SfK3qwFWkBIYjDzkd5zPmMpdzd0967QkDJYZ51pCZ8
+UWhosa1TZsz46gaKrCnUqS5bdmFlscR8S4Uf6pe0GT7qC/mJ84UTmdMqo1g
13QI9+PWKcET21MYXqovIbXKebBuviKs8N6NibAlpU0F/GYaxPMh5mpKvcZy
ZBVCDYTt+1jS9xHmuAfknZvBcxMwlf2uGssvEA12ZOMgjShfvxpOUMuqYhMO
tVgPpnSgNWczgcFN73Wq/Q1ME6s5K6sVJvr/4lBmZnQKZj/R/F2s0V6KVpWJ
oXMKwmfU3wzqxVDtSdACWfD6hVk+Kq15VBhYo/eLfd7CgBXQ8g+6swYwKm9P
mSLu4emlY7jt3LuhPWHtDhoVPJ/tPxlaP3xaK1Rxrqqz+PI84eGD2tPAryS9
PQsEf3RwotmNL73VgcSrx8eYjN3g9BzVdUSL4wTvmXVVF9Cjg+sF5/NYogfh
KZcHSDZXRqC6A0nliv9xciPVq2yTkfZxBRUiC84U3JLDKbqgxnooyRTm0L0o
x8CjbKqfUYlKSVJQzNGs490NePAbeaPzsl1qDUBjFtTzCBjhEC77nRtM4z3r
t7jTbMmsque0INI5+h8puZ4dOdbc4nGWdT9bD1BWTDRjyF3jXneu2yrxO530
oDme/qApudzklnLPYLC55HrThRtogoRNJ1mZpER6klbWjowzB5FU6YUMrsxe
Q55GtpLXkebtSUeWV+1nBZhhoys2HJ7jScFwz2dlQbwTBHNCzabAkHtS63h4
dQjLZxWSCgCqJvaKe0WUUclMPVkqDn5qlBQfO6SzYeOE+ttzwbI11OhKcZYi
FWPTzEoLQAt4tUfiyfCHtIr80o+KtH/5qv2NVpdvXafo/bjdS+xfbAnW06x2
xKZJgxcUSVN3LfxbUYLNGJMZh2cTrxg6PpckPTygjobS9INtBLbqDdgtSOPR
2gnNjCnkSu5xA+3Dp5B5KY7KxokRXlCtAA27qwOAm4zEL2t4fbekfc0UFX32
VrnYbRjejhKMbDdYJ8zfiq9etJrqxnITlTlAZr8FoFupAJHNjPkP7tD0oSIy
n8NcOp9KkU/nWGAkKg6nZWQiiFMlP+XFnRsf18Qb+zptMXh8HyaZ0pQY2rBO
2V1S50myOgsU4/WaZye1cUAZJs47s+LpRbQ7qATeGsDhgw6SIDucm/Q4ZAFy
TY+RF6InBGWMx7XaaQgwoBdQyO7K1t148v3Kmq4UvvFM1zFGcq9eGHfg9vY8
WM5rjnFa2TT/JX87fwpjEyxy/Q1K4+L6vBIq5Gk89jZsdJXIsHFawYbAcQYq
tATQKwsVWCXt7rzlYlDAj8Hir9OEUyMaICVP/uYi8zaFZyfYSuXTRP37qY+Z
v4Q/PAdoosvdXTLeiPiPiM12l/AiMp46CaGPqGKh4Y8thSXk8J8rLfYdf9V9
73QdsYstqUhhcitBPoWHzJFY65jqi7k7qSHsGdV26rB2X0TtcNKfyPePTae1
Xrc/10NX9xVf6NRNIY/8OrO6yXh0GTs4+Btyyy6//IEmSfls7+1OdfuWo4cH
tssR5JGaOudiUWZa/o+v+qTYHYhy9YAPFIqbyjrCe0CQFqPbUKe9SuYHsU4I
j2wT8cBPfpNy6496+2In9fykuTb0iwsPiw5vWz2LVdN3j3jIprLyXj3PNpdy
6c6Q7FAMgrm89GSK3fGnduKGrQ+vyZcgZnsNssFbwmblVI3+4xzzC7n9MaSt
CHTkRkHcvX/atJDlQ7o2yTWhAYMRYgSRLHoZXEm3zEBqep1o3w4tExtCwgNr
IGqDJFfkiZ8eVbjUinBb0HJzvpOhVHIrGXG3nI3nfDXyg/xRvjv5aT2VW7Xj
EQkVrjIdT5f3poX92snQkwLLhGd1VUbMhQ4gzSg5JgcKBc4QdRxdUmN4KbUv
Q/NOrog7XdtnGbUMsPz3gmqx+RWEa868n0Zb5bg9ecQy88ew/H3Z5mqY6M3F
EqGM9SHAb+kX53pdwnhgHzj83MsrsJLBfy4FcJxYnj48nbxgD9POkwR9847m
Wr+85MHyeeegqakwajuua4IFS1/M1ianL8g9hjOK8amyExJhhLnXOuzJtObC
fRqiZZ3/N6WnT2Xm6z3JdTHpi8IvED02qLJjRP8UDAz/Wr6VlZRJEh4Slh99
vMBnHB+HvwW6ao9FuHJfx0WLSEktad8rrlmB597WoK4MYT4MxWfZfc/Nf8MO
32/tn8h90PeW9UzavQ1E5zkUXRt9r2+uRMS3m7wbgXxEnb3MW98RmPil+6ba
W8MrUzUBTqOoS/UBff9SrNJgcb75d+kbxs8e6nwVnfy1HwYuoXNkxGHwE6Qr
qndisNTctFFPf4filllO4TQJWl6mv6nnsXO3zK5/Ot6oyhYplXi4yrHehdBt
FjO0WnVuxbmubVCJ7ZRzTJgzrfWjRiSfAlzrYj1NbEQJijSP0wPH6nzoZBEP
7qTdSClTv91WNxPZoUdTSyRSFl9SrAHoffz3jayb16moKETyiurtIbFTwde6
QuaYRC1eMVd11uTkhYlSEXYZhwAe52u6OHupxUYrT7QU44aGZ2RG45rqAxXO
bPYMAaVErH+HC+LSKi3cHVFNUvIMFXgvttbDc6Whj7yvIkTiZDJ5ttrA4fpA
9rvqnXx+nGO8qO0nCGshtwiZWCxjwJgI9Lg5coVxw2aCxfqhVTSemty1eKHB
PY6OqdKMDflgOWCWEC3EcMnhRm/7XVKdWU2kAjVWg9b/T6SaIjcZW+nxj3Re
Yo7gt5SCMrvnF7rJwj7Yo/beMhowQ9e/lYw0pzvZ/R1Fmpc3eYcYrga3ZtSe
keFj16jSnvzd4yTtQZCyFEXvzVirLp0vwr7R7fQTATKnxAKod9J1TtukmLTn
Z6h7ReGyKkSgle/Ntt4lSFSqBAEWhkjjsHXxMykA4jc50FfUuis8QzMtAIXG
m/v48ixxiAnCnZt5hLOs9G0fBZdBKOXmhqcfZ7kmTDBXYhgVto3+KvkW6Yju
kqOAkmNGU44kGpkb07kIoT879jZJ5fKFeX3tKfMsWNvrL7XGuq7C5YS0Txb+
RLLW7Jp7PTwxWLp5TtBMoukriPUZE4SU0kkT40UEBiU/Q9xbX796vEoTNpu3
erdqRG+bDXg66Y0xzROS3KPdeFdUz/qDwCe2c4DSF6ppFd+Su0TZbkpc4R7L
iaPROZJ3bRx6SlgAV9/q5wbSDOJqTPoEQjul5E/sejjWIhb+YbuArIWdzpqX
WrAnQ9GC8wVssWNdrKFBhwn2o82WVysod3Qdyg2YYIDUEcX8Oiqpr5724aOO
5JarnEDWw7KqSzXuVYtECXsaFS4oQbNDLYlOroP0lQJ4DkkPAEl8S92hJWyv
RVdTK37aPICrVV7SL3dejKOCQvICPDDqqM/Kknv/6oXKyg9rTZD5uyG1J0rD
4O10tk7237czCsfgi4PDoEQOaoBDpouuOEFFe/fBKP3c4qRNye+Omjt0T4o0
D+CKE+GRWudZJj5AitqcsiBKXip+WMfWZ+EDL5y/WNCm0DAgcV41p3dJ3YdQ
WbshP9qK2pMzHIRpBKnAjYS+9CJxR75uUD4MsTUQhnS8PU7Vs/Pkh7OkXxfq
QREmnWE3/Cqtdqmo0Bk0PUHVWjODmF9FD43LTDRnlRVAv9uqG4b1rzi3172v
kLvgCmMPf0wZ0AdaXsD2QArSmgXaDMxWl7XBXav3jf7cIhNxSWcZF8u4yZBp
Kx2hqipNrHCzbo6ALhOohsdWjBfSU0snaGLpet0Mr1As10+3cp53jNSFeZeC
CH5/yuSQwEry+lKxbyEHpa/R3G2+UOcL7H0ALZNgpwgqEZjduKaoah3TIx7W
7c6RZhpt9z11qPwedbxTBsQybm7VjjEhIUzWBAMtiec4CDVj+PcbO+rrpHxy
zRPN4/xLP3Db6e3Q5qpzShX3nSL+M502wjC0kTfTGvwBaD5cFFP+VAjT7qua
YkbexKZMGgvwyH5S0CohLf2noQsNFTGvNcZHH0SjDdK/9LQOa1de8bxZUtVD
3zZx+EDwn12CBcMfznhsueqPNX+n6vN25vScbiOB0VrqMhreS6T49kCkynpU
KD/Zqjj0OoCXhYorGtV4H7gd1XWxGgVSDgkjCdDIcUDp3SIhlMPKZN1kicql
ooWUCN1vR3/UxVjuhW0hMOFRf9xRHPnUylfqiRyA4BWKewo87IT3QRZw/OnZ
CzsCmmnf4WkzE+TnhCGA6dVrlg4l99LrIxJ0PfI5HZaWBmvMopZ7Imp11w6t
uEuSh+GeLuX7P9rXjszUH7Zpgg2ZYK7A335+Lcwqy1ZSZqiwI8pvIoFyiCbT
TIxW65SXb4HDoGHSmYaBt7GTybrdXfaDsoSlVfiADKceJ13kq3I1OTGd26mw
+qA/BkpHTj9U1m++6kN3gWyrFw+irc8FFYRHMYgCUe+hAGySVQZODa2ZOuMS
zevNnTNDx4/97oc3EvnQzBn3otscqxPQ+CLtDtbahpVRMxB9GoyHR8GF5Rug
JSI0PtS4IEgS3L4XYp48sIeltCYmUaDOpLjLwi35uKWKFIQIDCO44zdTFqeY
zTbl6o50mUnJOcL/V1hDD2NymzYzOSaO8jd1WgRKRlx3B8IWw30sB34YkWVK
bgv3Tn6NxqaNS5uYfpCHczIchPiJJx9qFCldj3XXW3/4jsGo0t2+06kEFxjy
ucSv5xyXhtpbHzFXOLLH5/UnL2jrmgWzAnNyhktoSkCWLLQTr2KmxN3BSxVq
fBnfB82wipTnEhS3vsqROCFVzTzhbeicEIHZ7Uc82tN8HY3IgfLy3nraOeRg
22pvzUUUgQSE9zfeCv+TwcNbYjjT5Cp3OEw29MeYkWIUDbV3Kg6HqjLOXQmO
aHnHYYzuCH84qzwOwvIildO0YsZTWy1xAN29DlDIU84Jdnp+M5WmwAAM4GJL
nBvU4oZt/HR1ySFf2EF+q8Hlabd+AfifWGqh4YL65+/Vrre2LGls1fRcqdyc
mmMcYGu7l4pWvhUwNAcKwJmQhuuv7HlUv2NgnTKGDFPml/znnO195aHb/e0j
ER8BeSYsEE/ltAMPbs8XiuZKZZGJV5HNBEjVZAhM+mRFz+/ZkLG84vTgrIpW
I0Ao1UHA+BE26fnPkedfWUx17gqwlKfNmWwdjYwNq3625rdW8Y20LRDUuGqP
O6uQ5BI1aqgkOIxHMhFmC8N3+p9AztjhDwOZdUwVYgq895sB/dzpQwnQkg/R
XwCLsa/RdwjmLf+9WEjZyjt8SnkQe5aO0PrTLQz/0djUKCO1IWMX/Sz2EEbq
D7ACPYFDxwErih3jOVzfpXJzLgB14VepeSzc5EaY/LszsDRIbkyegTgSHxfs
v5ZiBk3/tefryAyMbENRuj2DP54CaI8ufJ/4EJGqpeRAmUFzPIR92tJkZoSw
9vH0T/iPFlPqJoodlfYfbaXP4Prn5iYagfgvYTX1Os0Q0smLaufkBQz8ItGD
rpHVclBV2LdrxQsS1Xx4o4hMpP3lQJso0RPt1o8221DRLONObMMiecebAHqS
oySRC6I1OPSl8lYqtaF162bhA94lhPEmaL9R5hF5ZfIyTmwV24d7Xs+IQl9q
TeEcPewIgsZjUMDmPZH3Eetx+n5V1/RjcAYk+e8gpe3ERkkmWSIp7gfmrnC6
VRRgLMonqpUgTkLCjLbLPv9NQoGCp9IJ+6aE+rJHB/eYlEBwCf9yiwiDAA11
Q4+x1f7zroxbjqeFsyDt43BBLzcC4TGjtXD/OpRc9ayZeDB764Tg1wIUb0X9
WHZAzgnWNxhX0+tNa2i0wsTgJ4TB6LjEr55PFltucUs96SioRdkHnBsCv/pU
p0p2IrXfe9PUAvDvPXI8dqx6wPkAovgNXaWyL7hZeuW3aAy+O1NU4xTSFR56
fb0STbT4AF+KejIvZO7RlR3cU0R/4P/EWpJYpQ7gJ9z6YwRTXWyMQdbsy540
692Gc8G/hiQhpBmDc9uoJVEUXBgGNoIsXrWKEdIgXK/euBpagyYdV4fSz2gG
p5L3DZ34UdfmMBX3v/o6UHWpjG34uADsf5TeXreTtElNcE5b5Ofa2eVwv5OW
D+MSHkvBevK4Y/SdUkrJBSoL7YFDyMkF1FPJU0s4XeJKRLmuo/xeq+8W8je/
yWtKjmTX7LazGjot7T0qhk9JCke0wTpYWpWu8PwdoOdpuqrnun/HOA1aJpRu
kLUFClpd3DUAuEWmCDMzlVDMeOdCCUWjd6Bh1RdBxpgex+OAvZFwLk6ksEcR
3nlDMb6ftUMf/xawFi4XsFPVSyG+i6kBWgSXQOzFbFFxjbUhkPdBXUwkjhz0
ExJPxGcRBY9DOklhTlGiuDrduzj0kEo/AR+/jIrokP8h3qpD1jBELVsz/JEl
Aq4myYXl60potkuwsFBlMcgYjV1rPFGgfz8IpOBxx4xWFzxQ67Pzupw1ndxQ
B/fy+dVbngjaNMfwiPCcgQvOsDQN8KxpCtUYWoOAlufAXaENIfZdiTpbKL3k
RrbliApf/0Pg/IGibZTWRCijQoSQSRHTwFF8OMznwrvPKRQSpIKpASJ65AjS
duGBInaIvu0pFAUhs42Rdh5SP82tikBY+/A7+Qph8YuPwpm1gINGpVYMAZxS
ohBl6dPrbPGMugqEJGbyJN41Ws+j7iFMhyFmY8tSp+YqSE7JJWeW7MCN6U2j
Jr85hFO/YpE74dcB1IKqKnr9Wb5Zb1oPqGxumaIBY5nH3Z8UKLOUwOKyblyI
snOqYbnb9yF3zVZ1nky46o7v5+tGkf1R5eaMywyOotvPhL3X9tj8kcfkisqS
6fOtjwlnkgxN+cLIaoByF4xfhMIi8eLvWPqnVZRndn0WgUgtahLpHiVxd9qx
Zwen9NkVq8BCFA4sDX/OBxckgHZI/m9yOpXYQNl3/rsS7niMpavmp+PfqsyG
oYRPd5ytHukjiH1PLtamnQLXX4zEGz0wl0JGsk/1QY6TV1KR5cphNWYSIUU9
fnC1UsTu1tKp3+N/z5gYQ0T54Bhxx/XTEWNOJkyJkKJg2XuHmnwpS2robhaQ
pNVouTwgiQ2EmTH5nJ293VmM+wkrcx/LMuPry6BpOuQ/2vyL/gqzVfrSBFia
aTT+LqbI9Ff7uAoPVpWnXZLbUwwhgHwc7yMbjP673HAACjI37al7qIfXXpHZ
uXKQCwF9VhalL16Opr5tTXwx9bVTC6AgoHgf5tzXlGai3pMG6pLmBiBnUQhX
q+zZjuZ12TBmYJuvs2T0+eTosY6gYi+GBDf7Uuiho1nShINb9tTqXRofdB0L
E+VxVdcaKLyEeRReLSWE9j2NvZT+fzBhW6FKskDhUOBSA8i6SnWcA1nUta8S
8bse0I8TEpwpQGhLp2rVZ8MPEpyvTIX5AVwy1JJvU0/DVCk3cmwT4wlrSQfF
Psulpj1xsREITfsNqX8NlacAm1FqzYcadarrMlonS6vo4EeN289kOq/0DiuB
m4DJNgXVWPMpOpxPbURrEyW2KbPaLzbIf3iTEKj3m82IC7+m8nkqfQnY7zBA
jMICcc/ud7P+EaIE21Cxf7N+0ROYVYPy5ywVRI/K/PsRG1y3+sv86CDCYPh6
I0pnNsmT8OTg5eMpyKMac1ACMp2NnCNBrXVMz09LesMHf7k0YyLHYRmLRYJb
cEOo0bHORNydKTK0jbhWlWkXSUeHGiE/GnRbFworl4gXVL/Yw3sHDMvrhNAb
Ho/RoLUzVA/8Rhml0lVezu5JBe3myJYrraXjrKhUuF+1Uj8v2y2Bhnfp1u4q
V/PgOdWFF/e5rs53clm2rBrzYFkF+eBg5V7qc+4WpMHQrLx4MkmV8SidnBSp
uGg10bKJcLy/cTkGfybMCmXQHiH51EfHxgYp7FZQF5D3RwT2bNqNoFJhxa7N
484udtEvGkoiIoeAaYzBg3N5mdLYM0a8P0BjqpYx193RwN5HxI2zkImm/d7q
elmnB//jvq4GafPY9XDIapWxv8+SPHAPAZOI4Ar4orqIFA2SkiaxrlwyNkRc
Ot3qAr4TUEZa8SKpXvCBd+t0R+KjIMxZtBShgawlKJMtxFvu179def6CNl38
H22g8GaAhj0pm9fnnpy97XbvDHFK2C4UzzP+S/AA7gVwXLhqIcDWhmdj0MuE
5SJITX1wcOHJX8F2EHbtq15EUxQ9vSRkYQZ5irZuDY9gom/y3oOIX8DZkNV+
FyVnlSGsQ4GMjCrby/qJDQ5qjJYe3J3GQB6H1CnnmvpeGMcFNh0LWoK1zqzw
/h7+aGDrxOmyvDpks86UIdxfllVRonDJiIwoONfVhRQhqIb5iNgJirYzelJ5
F7yyV9oqggiBx34WXrBtIB3ffDEzGoWLWBZuu7Q5sItdaN1rVpaKXXIFi+2u
rttJekfT4PwRJ2DmKMlqq3NbYRzFm/aS2YyeK/up3w0kgd/8Ilaf4IYY/84z
INZDAgdHUz9biHguUuyZZAOh8Q4URc7JuSpezegeMuyix5qG9AN6jAy7M3TX
Rv9PYlFcYQmUnVA4pgjrtRf+GHUZsYm246S+dYY5Acx8ipXszsUueVJ3WXfF
SVPnsWs/82XeIvusU6oqo//i3OMtlGkb7bgY6/yt6/enT3K/JJ1rx72fmnu8
0IcCOL1Gk1PYY/FknFhUnR+bVNWLu9Jgnx9BOQV0x4FKe5m0Qmxp7tSiJ/MV
T+D/EjhOZDjqspH23Ew3W6nXVv3Bux1234KgIhjsdc8FjGn4K6pUC1EjsBm6
EE8ybFijbm04Ysz40QhZyQV1yknFA40HZRy5QI3glIzffSzNwZRl7p+KSqM+
jopxdf6lAotiiISIWlF0uvnIAWqfTLsuLplydGRsB6nWOV9rETpS4gqbfk42
/mWhXleERa2mFkpuYHrvtTxzLHw4+k6YmlwwIc4y+tC6SxlOWh1W0OKIlyWm
9/STCqdm5rVsMYiWDmjVXAy07hedGzxKppvS25PIeTDQIxVeKBXBVMrJtNjm
NwJRYBY4IRxGiTSRZQhquYHOrQLKBJ1asmGyZ9oKQqYtSwGVd0qsn5AkqmBu
1XgYhsnEEnJqm9qxeCVvb8w+QimzoOmg2ubRIrxp43vz3XvaMb30/VGcgsEQ
Wg9zz2pqsNi/y9CYhPTZc7hy+D/ofKBhMq41mdUImvxa5cZ7xetkzTXvpwbe
oHlFEtBemKesPFex6M3ygh8TGcvEEk+Y/5cKzJ70J/mpy0mZ4226yOIQFC3n
+Oj0ZnFKFURUBh3FxbjJqJY7HGcjYNmEKqxro+aVxKTYYOsNSjBW0V1o4xVa
0DrJNjpzaI7vTCkm3S3HJGpgd80o+NPnuPWfj9OrHoIY33iJR2T86BAUe2QC
z2+ud4QYPgPd3rp1dwGtUzbtEFqhgmGss3Fb2EPdIavZ887gFNQWYv9LVMW6
8Rd1v2vV7LwwTPXARJH+V2N37yLIc0+dqq8S90GD1SJPuI9VEsBD/3EhOz5J
5a5Vf3VJHwnE8kmwEsRjw8NG8I+CmuE9l1Tk41LwxsEdTatz5e9JAgZ0DIL6
cG7JPdnGvAGnIdAtVW3P6d9eedPpglYcE2uA7qwC5H3R97t/0tDfTPmin0ft
zoFjICh/wiHf5EN12g1lYHQdOuaG2XUbfvtTX7FLLjukYzp4q1sqG59NrZ56
BO9xvx2foYYiMtGz6c+gxC5RPfu+0dXwRbCEglVWDvrZYLBqXBXVNVGdO7KQ
1NO1MgvQQnR0K5kv9dj879O+L9a5kuNwqR4bWbN62UsFaTatXb5t780fj9Ir
K++Gvezdcu06jAt8nPp/iPZpSerc6yQgcNCKx3zsg/CxRE4tMOxCaW6852A1
0UsRCDEHVGwEWp7NLXKRLLOlx7YzfJ/3ZClpSrJPiNYijtPI7ivdAHcIiBRU
GIlr6GWLRJHaFdRqHfkURvcvd4zAYt52XTi//79aEG7/O7UmdFEyOPzhrIj4
LUpm1AWyw28UWxHhJOK+/OSp+gzQXCeOqPZ2qHATRVXik6xLLEqSLF6kifjd
2HFxuXAc/o52h4UuQbVXylcoflhy94I6mqQbsZWV2lokW7ErZNH3G6kOj1Gv
UHxe/Da7AJvq6rV8tO6+17LyL/UPii1Z7ehBmjgb6lAEG1U3K6DCUp61qqfk
DDDEEnM3Y/MKOyb9wNYKnLQisygXv6wBiMXn8sCL99JfuofUqA6ZgWsiZuRx
S4/GQHCHfm0DsR7N1awiAKyVJJO6JVamecFZYoHcgMBuaz0j9+C/01H/pG0z
hisMWczevhPOnJmdig+YJ/yUNqmTK0e2E5k6lajxKsg33O2nbSKRMTZucQaq
vE4vxEyEStvfmnetFa58EgupgtZl/4SmCrOSEKkr9ogBGe2hvtQUULLcGQpA
rD/wENwRj5C65fxas7CPIYW6QOxycoERzEU0N0uZwjw6r4fuJyL+6Oz9e4cc
0JfEBRYk7qPMnI2NnQA/4hAwJskt5W+Le7mro1CB5Gx5tnxEf0j9DtQSoHNd
TTUP7fQlTd8RsK8kF3IWwF7X/AxWNwgE+9PVQS4mB871/RTYTi4anTl1JIN8
juUnyyeWjjAJeKedm5ail3hZxq2PYLMIlrR435DAzqVb9D6ZE0vNFnk4+tbt
m6LXAB9ODXbu7mNZSNRDCXcnz0/B6iXrEM9K9XTOxw61kGYkP0jySDbMwfbm
bmeIAKL4CXNnpMkpNPIvc90lnXtoWJvftCd+MJwYDnFvPwJ0BuA7BglN8zEm
MK5u3H9xcqQzNwcqvHD74eYDmBvUqFrwe+gN/oAoPLOt1PDcsuD4oJ80hKB1
yqJJbUxrDyQoqvm4rGOLBlOuGnpa1Huoj9qrRJWvtgZBTw1JAcOVpp1UHsy7
EoPbTEZX1VFTOQEqq9RlqzqLgJdGFgtsOVsuS47zfSs/38pYQTmlT3ew+3M5
UEXdupQRAagbRiPSMtDmuS/PJAgefT6S/v3EINMvFLxG0sHwye4Pxy56sxeD
ZOwi3bWQFaypwnsni2UEcELdgM3f23GTTMYHabM811qq9Qu6tE5fMLdNjZZN
BStaLz1MsV9jeQL1SeeMvwmyiyWdUsAN+7t9GidKAEz2hjYJ+N5nts0wkipo
MqJuv3/lhVaADAqnN5AEtc2UY7H8f1ktZdcdXJHFCfYEu5IGk/o4F3LlHAi+
3n2JGZoIzhad+v0raPWO6Ut3B7YJ2gtFg8hAvpNa8MZv7gGixxJHnjQCSuP9
HOQloHeebsmAL8/LlpiRHucWSHtM0G9zWBpJiTKZ/4OXztUCJe0tqQPXu8S1
kBNcTJjTryxnhx7Mmup1NTpmeXMCJGvzFF6usRfMrR9Tz20pIXH9EfWclYIh
t/SAB54TKkw8fRbqQklC4K0qZlWBbrIQX/+BAezy8u83MOGjg6Tt8SF7g+zZ
rZBsK0w0thbrza+2EOI42lOcfsFhdqKcnpE8l2s2rtTeF9ziqkqgL0+FK967
XtWcsbVHwlr4DEW6OZ7zQFVRP0zSbsd5ahIvt6bVmuX/oPrvbo7d69BKWX7r
b9/x6QxqeYxMvd9ENyuIAcdvP2nwusH6wRcqQzHDuGx1ynPmADbyMWt8cLNC
agX7zSs95D8zb+xLc3ifZbAoNKi8SjcjB9diJf0slrh7SjQIj44cxu2HCmoc
k0oS7ZSNSaR16a0z50QoHahSyEkKBDIaB4dOAd12ArsbnsD3CFK14UzEeAY5
udVlXdnwQJyGGXUTiv4BgE2Zn9pntPzCIcJELx2bOrIxg9fpGTCBhnQNB/R/
oIV0PT7PVhJHh5QLwKJd8amvdtmJ4S/IUHIBUw6FtFNZou4GQ7ra1kvsNWYD
gKCCnpTABH0Juobz3/dfbjCkikOKw/Y36XUtIguD92RLhowwkRNKNMm8mC3j
RnMBykvEe0MHFApVpDNuDjWmiUz5fATFYbj9qk1TCxKDgrT1ppd2G8x9Y0JG
Ot+tldoSWOxeqatwBExUmTUEzwncNTbI0e0phZ6zh/+cAgFBy+3Tx+/dgOPp
ndru6t3lvXVR7BsqPuUWV5APPT9+aSWoGgAmu/aWmyydHgSmONEZERFfxs5p
embC5kkps03YwLU2JN9IovmAvRYF7WZP3yrs+hMUBs7uN22yyuxPtOADKs+K
X82unf33QCOYckOFXBWDbtWkyqiKdVtM/GGyAM67P/LH28wpdRNyFdv9W0ZT
PkpR6E0i7r1/tZ11yWRzl7gaalMMDOevRdYVRtSSFM7rkUiAWE0h8DvGYVJk
W21WGjCIh3/7rQ5SmIg9cr0ew74+kGR4f8MijQUlwJoaXxWW3zwiMs1R/C4+
w9rRn2fraiWpT/vioV4cS6fC+dsEAGHBSd7Xkep4W1nWDMf2RVXyO1gA7utf
jZO/lU6p+thOI4rdnjo+EETFzFha5dpfIZqK5GDfUYSQuLkNeov/Wx2a5Bim
x+sNFtHVMFIjESLmprhAgwS6JMY3kCa2keq5jBM8UbpQ+e157ooyMQ0H6aVe
KWU7AEtCPX8WTiL3JHjnqNEseIJLbzZYRy8Ft139z3ruF87Aj+OS14F+vim4
PVGhXJ1oVzTbanSQ7581Qxx4FCwtng/tjNInkYMS5kaYhdRJbkLYGx/fhUqN
e0Aff72YNw9Vq03yByOsGskZjYITNpevs/g2HvTNfw0eFLgk9uckPbvAC2dr
MeWJZvw+2+PriFclqiB3Evwx7yXcS36Y1YyiRVzlND7mv1jsZ7pqkaLe+YRd
4G1H7CyaGnXKvuwX9cshtqecnmrwWXDxSmolnFQuEAD/rTePylUxAKcAspsO
G3w/JwzGQdXaY/S3pTFeSQJJzs1tuvmNpkUGcUNi7hT3+25DExVEuiBofa0e
jwaLfUudsRt5/HzdPmQu8uWaEATGTqBubTZN+5iHYNlFaT6grlAO8u6+wR+k
JV7Cu2SoYvC1JQaHHLnFUCfoXlBuEiv5fiywqyRCTiMUTzfOqS35tqQvJTtB
H7WVa9UUMwjhRlcaTNoKcCE5GtzX28I3BTVK3tJHyTpPSkJ4hvjtFQTWc3Zg
i1zp+ZSV9ARXIfAd+/uv5deWNrqmsfn1VaV0VPBHs3eZ/Mtio+3y9BHNyAwL
ffikS2HLKVqF9IzbImyZVRHfhkeGjSxBCKqEt1nthXnSL5me7/IYYTcJ5mOT
2vqnQPNF0XPXUMf1L14yxSvvUHTLVlyivDtj0ItZt0dZCkUGooJoc3oFCTHh
04UJ1bN6NdNFhiG5yOIq9l9HDpTlQlpzucnxP6Vik2Dn+ZZatDprI4IBi/k5
43aIz0wmIACZfo+4s56BPxiHt1IlcTjVNuQgfcRMaBLp8TVdSsvZtJgmd9az
jMyLLTA2TDU0tbJP4FOX51idB2Eh0R2iwiD83dmFHmtQrmkfXLqKmVO19qy9
GZoPp/hhzYBX/Y12b9IrYffhVxGX4zBKqcDUAtJ8LKUzW8KonynAS902dt9C
tINvDuVJ/wCmGho08hNhCPr0jL5cwtmqoX9IIcXM2AMd/f1c0Wu/s8J2oQdc
hg7GG145hBdgXQ2Ydh13ehhAFf6bADonRof0X1/7lIS34x0rY0MvzkHX61LP
h5tJJxeIqfWfwPDADzwFzQrlKhIrfXct0QRNZ5uUNU2xTQm5zYakMtyLf4/F
Rm8OKGFNjGBl6QjITwI1h2a7+O7aYI7p2vOQx4rVF5SRbvvciVEAgl75Wb0P
Cp4wsC1tIa/yACun2bsgzahXO3So93d8561fFi3UpTn5dT8Ud23dCKdHxinZ
HLqjTFDd95aQlxZzztKjrW1eQLjMnA/0dW9ooCNIfib8e71dCudy6G/EQd4Q
ShpkFIfDdAMdes9IwOyJEL3jcmc593UyRUN5y9tgsZ6IVNlzf3aKlNW5In5Z
uJG2RCYPXTnh0tMN0ohNUb5YuUS3fyHsJpz1HeGGnPbbmu14HTrZd/mvi1ZM
ygS2ydJr4+iiRGjAIBdWSKu6nwdpxlHX4Qx9Fj4Wlc6T0L6PbjDX6NnVlQq+
mvi/QoP3/mTpQhsJDnDbRRoSpJ9cgCsO5VlkYf58SWUKahv+nxN01Wzdz4Lq
zkcVMhjSQxLDOzXtIzQ9vD+symsy8/NNVZ5yu//sodMsvgwPmrDH3F6z46aW
vmK9TnTnMI8YLzAeKWocBxxiF1JhVKIDXSxeibIfEZj3XEjYFW3+A9ACfXTa
bBF0+U/sbc91YEMkj1GCPKgem+YZ4xxI8MjqDCYhXmwul692O1ohg29jDJH0
ns0DJjjnkPd1JFH6CA0Q1JF8UStgdQpoU2YFgStzonzxoksuvP37QQkSpzFu
Fwk6padLg5v6+XNg96N7buxgJtFb2Yf7T6cDyARyjxdMPnPhn5TXeLBpK4uJ
wS26CCW9FWFZrkr6SuPzB3Qr65zbPcuYZKsjnLClEEu6u1zpP6aVT8Q9LC0M
rC+54YjMpOK3pdv+TOGoqWuxBoZFKw63lUN5wVcNHeb3UO+gDV1iy/qysMDp
/E3zdFTOPaZdo8L4eBGI7zyy+bVpWqcyDYhMaj8ShW86cGFiBXBD2tN3LmZn
YrlVkrjWCHQA78Qmmjt/tpzmkFGEtsWjJMXEKAaaXVKtyL940Ojf2WYVdioF
1zH9eciRjoL+UIELDO1C7PMeoEkg/F/odQuKzjJoTFH/62Ff42E9C6eLOQ03
4YrHfRDJ3bvyY7Kn7mXUFfv54yNbkzm+geD5mpQc3HiUbr+Jkj5otCtNjEi8
HWChJxwf/HdvSqOyCMdT7IUEOTE85Z+72GgBHrM3vKVAOmsoII2RxB0z8HHA
vH05I1YTsqyD78+L2cHLHT+FthnXW9MekiWhvpMMe1kc5f2RHyES+CFIkB5R
7cxGykRRrf9k+bHEMrcVduKE+KuyB8gs02vAIRK41JNp1kobYs7qz+N1rPR3
fxH55DWYz3Yui+TbNgr7TnbSqk+2kZ6xXFQQPsED1ZbzpdodGuQPGW/55cHv
VxjCr9A9H2/yIn3/sOVe71BmnkwS19khX8dFcHx2J1FmgPfr0+RhE8fCJGWe
sXKpBk2+FiONDoALDj1evWVsGLwrP63vpKXJo+EJTxRPCnYld4lzMY8i+zRh
ku6dwbDPxMcGzKTPB/wlfxLuOvuPk72C6nTrEN2oirZXszOQVfFIRHkYzQDm
kxpz9iNots4K+HqKkyqBVXS+IJAGBwbqsqXsrAYHpvwClEolrJMBt3xUbe90
pXhJJNKkEVsqoBc6sQznYBcBmf7b57BN3st5QKImOjpSpb67pu822jmtdI6F
5O9/7b6E4BNK2yWi1WAMJzUKQqac78v59aKb9UkFT0vSxhVTM0idXky1DCEb
IpjnyFpAQlDZZ1YXi6cOYZ2/V3e2Vc/glFSW1X95bmKXkl6L+aEuSYArgnbr
7J/vZRFTkDewfAf4lAtX6/kLRb2yL8XXetzEP+ABmtBatqXHFph+gUs2aB1T
IJjdTgkhEzHWAi5vqkpRQ/o0uQ2ZsWjtiDizNRNLNNH1DMQMf+6s0cMc6XmF
Xr4uRkhI/Q2TCRo6lhaeZ+64pSi0/lhqtkJgP4o5PO6tNyY2fTOgzqbQz6uR
W98Mw7L2cVtOTkmoZvU3gjYHgApMDutMoXMu5XGs/Kq5JxOwpxj5he6ZTkfC
2Pqiwl2ew8moUhqsxD04xvwT2Txrjmx3ULwNHn8D+c2mH8qXLpEMVNU2yyXY
0rRt9o1Pdic9oHeKGDWgb1ClPD7O/s8iu9yq/ChHNpekyz5s+TfJ+h/kF9R+
gnlFaLCdSjhoqXl1I6jrn1SEFaoXoph40R//9dGQIBNtOk6v4w0XGrNBG0AH
L4cpF1OhiGevC7ayXb9RXYCzZ0rjIGl5CJiio7LogXoK6LlXaMrLjaHyS0/D
4Jzb6m6U9gYk437wa6jLqwTCI6t3YtaH9uREDPy++6IrR1TvC0ES9jeUeGzy
Oo4URCIwdqa+MV5yKeSsnK1QbywhrIsp9ShByi5P2aBQdsosDQOgpcT/r2NV
+2lOehKle+v7wHdb+Ekmc+1lVj6EFJB8AJR9CW4OK0hT97ifziRR/Mw3xlQj
ThsuRpjcC2Zz+BIDrpSS4NS+lwHyCTN17Si/fM+ebqNHQxU6OSMNS7gz6E+T
KYXRvxE5KGqTpI6qBu4bbd7tke5VzpYo1Jv7838/bY7XDMU/YylfRuLuZ0bw
vmS2Hwwe3GWP2NgalwoIhcHB4pO+aF2U7d2aEoPYbFoJpZclBz0S3K/Cr8KK
aoWM1UExedpuKJKiC8f1JGxdUlgEPq0H0QtGOdIGml1ZBthUXWfqSKncs5/K
D4oJtTWonSvrFq4y/BMx7V5oBbS+QPihSWGZgGeEYliW4xDSgCuqlWqCZffO
OWwUT8oIUuAdt8Nk0WyZd10z/Luo5a1yWd11OQMuxx1SDnnqDr96yYDeXXCr
5BRP8YMIPazhUdDLOn8tmmxdnlefEqBT/I5coTS9KzAvT5nTIkHWUn8T3qsW
+n6UfT0G+cDcuyataw2Ugo9IJy9oC9PrdbvzirLeGw4mp9quWtXvhLYnozFu
B92guYJp2rWj384sNVSatCbliEdgzF/Rm3ubbXO0bW8t8MoszJLyf6baeNPp
WuCJ6dMHPxVaDNUD98Qr1WmUvXJb/KAtHnN68ZkKNOOFB0fP0aKZbcJpZlM5
guI/kxRfST2AP62UfFXiUlTdsktKiOOiFZtIQZuCShaDYyQT3UMH5V8nAff9
7H/1cq0l9qaN5Dc4617nWxT1Pv8bsM226fi/i38Je4gTJt5Dkt8cVusWuCBH
iAIG9xymr1jO2MPPXM95CyMSbXJm6l5AHx/SKJykrbjqq63MoxTCpqJsRRqR
ET/sRPZDHWj5+cIXRICQj/Hn/NYssjekjDTy1ABxz8zwvpnMvX8nzqhqOQ/6
tjAcHTd5WCB07qs88sQokDrM7IdYoIQuZ6twIjWuWe+wOJABrBfegB6l0Aw+
LIe+rWkbVqXA2db15dBS64Ytu72bs0SBbCZRORUAhxjwsuxUKxNZLG6hltVS
MF4dn/Bva4z3UYG273ZbarjvefLOVqsKYn+OgMz2FDbZlqiZ4g3V5l3aXeup
+S/E7tUT2BV+f47Z0ktsa6txIyp27He763qsjkC0Iag4fK8UHzlUjni17G+y
9F2MCdUQyiilRqFlslKDi/H7dTldmHfI0MqqOAHA8DTzaAPn/lGGTU0jpA1h
nilcBXYWkie6gCOCJEvZRVLohxbopDV8WBSgNwt2+Z8AsE9D7ZhjTbFUG86x
pDb75ey7ME16NN/UzP92OdIgZWS0w5MFIgRhz9xB/cL7LEQbLGgwT9tme/QV
ElbXvE563IvOs/mKOkgP8J483B0iUeYDd18UhE/7laDNPdERVYqJXzrPLWxn
8p7jJaCRRoGH8wM1cZFBMPy6HO+H4GAnz9ElnenYK+d45CGGP7aA22R0GqlE
GigOov5SFAC2vvHzOrOmy832cDZOX4NVQqdE7da6T+CK7D/qYnIi2ddFkSWe
fpP6V8OIWv6osFrVmR6rY7rZ80iDcZgRkjNAXwLC7ZqKtCrAlCcr7KZxAYIx
b5S+vOMD7S/j+shSUdMdGMOGWtQmkbSXDSIXbeF6+IYzka53PeLI5mKRqZVY
Xs9QEkqOnwmRPyWUPWgGAYtpS0QnGX35vjgGmr2e6jotKkkLupPS1KUre64e
lEgroHghbqresVG2ki//75bZXhq3P0LjVNWwYsnkFZQGc2iBbfuIRzhW44SL
wlMFgI463pqeMfDpgC75tu0dAe9roX10GcrUPHwZ2Aqs7F6tx5NpX3t38jkI
NFQz9rSy080GIQIY60LzP/dR3VjBvFMQd1h38Fo/kvPMm0qgwkFq0btwtxbN
Bs9+kA1yVWi13Sxii43yo/LRHGTmhryeshmMrqSAslnbPSGv2lj3Spz7Sg17
eVB4/9VjaeaFskAq4w+iODsI2VQlsk72IAAEA3g+0H57c9i7kvr7musaJMX1
LNqOS7xfQbVAkG7QSO6x/eZeZKVSbnqF/nO9H4f2Vuf6XGEfddszUb6StZr7
W77lJD7jtGx7buhbQGQAWqttOOsnPCVaFzSnyEQfnQvWfZL+d3Q8sC54ljfJ
KhFAU7j82ES5bZ5XemeqZR/lZ7NJlD5wJANRcqiNPx28EeFlhPpnyFAe28xv
VdZKQ40aJ0a57j8X1Wm4mozvNTHrxE5w9+lsGE5JckMBpD8gFWFKMdCl4I4E
0nAkVEdnyh3yR5xgNGqRBuzClsPTBjRj6s7qiDEJfl1Vz93HXPeqriwwB3Ar
HkjQfFztdaAqtwMXvcRYJvtvTP97xl/wYNkiIz7mApuCKvWHIVtFvjL4wLm0
JK5uMQ2GHJTDlMKxhH+HSpI3R82I803OffX0EVpmOuUS6dZvEOYKT1k//bb+
+LROMIel/cGpzHRKi5k18EK1JkfL8zFbc15x9tlzGE2gJsOYhFuKp1xaX+1C
CfAtE5R3ZiucVOnyFUrGW3bBBjMirh3jxAp3oGgIYRzMWokRvFLIiQ1Me6Gg
in+wJa4hKttjK/Kzoa8rfVRpHrqJhvcujmU5G6zboAreDO+KR/ZsMTXreH5r
W8a0K0XSzDzvXlj8cGN5JPbPf1HTdOUgjGyH0qDN65hLLWFvMl3smaUBG2+N
2fPFmIPlbgdIU0N+iGLLhYLbDMui6H0oMkHaUeJyRTqHjKxj0MQY/JU38HJ4
S5iJ4Qu+igRLd/VcWU7Kws/DkBVoW6YjfqMNe2sgKrdUhCgII6zHA3Kqh/LE
mKbPjtH3LTC9VTT+HowjZM+LhvbLI16zWwlc/5ZZS18JrEQ654brjk/jvg/s
30I+ilyjruNHuPWbFfrFGPtxeE3Wh+sEjliUz2AJ6Pgw10+kln3PGSeDH77d
ZTIKOQv+NRsqwmnNdSSxBEjsK4reQxIpVpG4InF1IFLpP93r+0bxPQmoO76y
+mDC3nP6xpbKqU+3KsYChhTANRxgsdXkHtMRFnkiWNih3yA6R+qtmea1/Co3
W87esMRiswOuE6NJYxYcI9uTw/KwxpdNAff9tBdIMwrOTYNFkZ0kQNWDThEj
PO+dgn6A0LvSnmmDLLVwbJjb9vH9z8aV6AYBloylN01lAuPIM/Vlm2PTqgE1
HrwrA8aq6DBma0bu6T670nq05t/ZBg+rIkgXQlDfAPkVUnxtbnbE91SVvJar
wktbeYeb8EXLosUohx5BOq01dq1ARGW0JhORtzCnNp6BCCqrsjZb3Yt1aele
0ZgmgQ9RKhLcWTkv+59dtnTDRNnDbjPM4ttbw/6XmLaraIe+XR6anKCddqte
NTh3bHiHo1KA4eALcuvzfHFvHlLBH77UbTOkuciFDeqWRNz9JV3+Jh8Nrj6O
F9fZz300+DldRNr+2IRavztPR2Sd4IbKbpAGgSmF93oE3R2u6O9LjjyJ0YRY
R5Cl9xatnInJa/NTSAVND+P8aFfakIcS1Q0+eDFBzDT1FLvV/H9tnVe4qae3
VttY1cLqHVPxjaYX2Ip5odklabROiu2IHEUelkDWjcbNv5RFEwrY7RXUuQ7g
FPf1AjmaNjAPtMQm4f5noCBRbU0gtMEWtQ+Auq+O8wmf1OHFiLfas6ja7u6q
YJxRcdQgQUEZBAVaclhyFhWRPg/nkXHejMpcyC9owIgFMBGnetL0EL3/0pKZ
JlBtVXcqi9pgHEGZjGrjJv4vL6SkLNgNTaIkoDIUjUJ2qYlQyljMk57IGKLT
IEtZxJTynKExhu9cPstH0XXI306O37Eh99+QKBz0FDt+Gaf2lBzAHIevZiZ7
82zDEdNhIf331sfFTsxMtAZ/JnN6OD9FIgn6Vz60zDyOXet26xqT6cyGYb9J
HABfyMdtSXiw/PJJ28DdEScwcQOmC2d9QwljPbHc3jZg2SO4QhfO/JSzWneb
Kc6WS5EzzHlCS7xyHextrZ7/YgEk0Z60+S+8q4yeG2Wra73iS7MwWkpB/D90
lsIUKAPWJl+ckcd/8mHR60H6sQubstNif9Oa3wBU6OF7H720RUVVRRggxXUM
/gHbh38IdA/gYjanlf+ELTwxebFl27YtTzwKok+bPPFUdlC4gpYYLVUudZCV
eYbsKL398dD0gNiIN8F6oCbfP2eRJZwJAJdJPgentFZ250fFP6IyjmUwWULR
ac/18pca35rQhjdHsuhy54r4YrWJ2+xyGyERFBU80NoseBMGKhzVqtAjsBJi
VOKf3Jq2I8ndHEY3YU81V5NKi5jmYQX6Nt1yq8oG6KvoRT06ZZMTxxgy2YRz
aX8mAodpslrnR8Rt5dftGcd67bVklYdrH6C8oYHX+zYo5eG40f6P89GZEpjt
3puGKw/QVsliVfhf4QzOiDI18x6WsMzeDe0aB/2RVdOHQZGo04Ir9jDlVroe
bTVMujhWLZk6Z+ukj5pvP1muUbOWipIIADa/HiTew85oahwL46R4UrUOja2u
CKYQTInVXnlLzTuhHPaddGCOmzrqJTlVFwlyJA1sh/sTl6gIdLLA9Z18q4XP
JfbK7An+2mOyLOvaDLbKTOMP9jw/mIUn7+RgrLfnMdCqdlA0MuFGQP2/YSFo
0EsdCN+34p7tj0PEp5zGq1MPgyvkXU8S7SfF0dxtn41c+Ek2/VQuMOB2Acyy
MgvfsZ2oxcvfndGscXKb88VsYIKhSbCRHzbNkBi6nXq4b36HS9lkQhLFloqW
Mnbths36oTo9mLEB9DxO6c+tiFKkSaCqqD9tOr6GcKpt0sVQgGIn6qPlzX/K
zgKHiC+vGHJMgfpY0GglknKDH4ih8LHfFZm0Yxg5/NZCYUQJTOaTLANbQTTn
L9NLGOTEhn4hkU3rGRVrXaP6P6LfStVLdyltL8XQq7TTS0Tg5KxQv1Xiq9kL
OJu/tHMjkWwE8OVdctOxsGMYNdwEFXp3lFYutZAOB5haqp7z73rKyJnARNSA
uYM8f6i7U9We3MghiQ9nfC+h78BF+qBQDhXyy3eHwZ4NC2+mK9kQHHkXyvI/
IBzCuC1uUjPdijhSf2s+9E6Kpiu4/btLoZSeJVzQILPadxdLR9epwAsplDAk
3I+BCIj15qvJQD+cm7jbPQuH6bTvz8km5tpZtza1j3bXFI8Vqm2T8A5jdzeH
FKOAyn3H+/5SXI31AA+/Ar/x784afksqw3MXulIFdi3bXFnZZ0/kV0SeEIQ7
WhMROoPFqei6Yj23o6tZog95lDcEq2JRplYGB3jJ/4WsQrcPojHkO928BAQZ
b/GZtsi1QTWggmgusa7O3mH/4nncz1DXnz1Ki45T+C3iUtw9XPzzhTAlubwS
7MZwqu3LOj8PESIQZMnZyjHQO9WktNw7ESgJ1paAh48k4580fp3hogTpll1S
BXVwlb7r6VzP2Z7I4fodYPVw+7poXug7w5WuO8iUqGaerUXyM16Vx656ClQ1
ayaxbNeGA1MeQBLeC+ACzWWXo1fbjbt6hsEShlAGFMxfdFwyzG8Jzx9QOCA8
nSVJKwighvAB7d4jldTFkHUsVBjefbwLPo7ianx6Ha5hC37/wfLx6L0NcBSq
wtWXr59xapW+Y/k0bSCjmseqU9OrWtD6EP2QB7Lg5h96eWwwOGWH9FrT53kD
UwWFY8+l6FTlFO6SNgHx4VmXxGxr03FfxTS/wZy1KhmS9M/7NdFpCyQ8Vy1R
28z6MlOEMUpOUXbdtWZelKUFOrNiPcKLbjyqxPsZV+DdVZWTGc4A5nwdhsyP
9HZ1YtrvCrSjPN/oqZ0+kPyoBm2Md4Yj0zCusEqz+pP/aHk8WRZA5Bb4dXIB
/6HlYzYuw3omJkNpdmniJVVvA7D/FYVFRz+cvTb+CdtgAm5vwqEAsYRSj86Y
AXj4l+JI4Ba+gPA2NmkBnpkKZFN4apVjTfOqLXoASCxz98r4pnNeflinZTCU
dVJ97uGxEggsWxzIkM1EyNG1ioaw9X+Ue5ITgfT+ujD0XPZ8fqyii6tyDfaS
O98Zb3I0YKPuLg3fp/GuQPelowDFnCp5ZSrUTjBVc00SnzIE5Et/EekFOBLN
JP4KfnlXZKXjI6WtZbu8MTjEVrNeRkJJGzyftqWC8ykpu8DXZOTvagRMiG2V
4OJ1FY5prvVMw41cpe3ffhzphAyzibbBZDFw9Q6+yytey7fKLcM9JVAKTl5n
2EdgSavhNK9a0m2JTNS2NulF5DgtzHqYQDQ2CIDvtuJi+v/+6r1HsHYUo0JW
XMKwJR0ZK7YqP9j6KGzaNB4Vqw9XvqWnnrhWBONjstPtWzAwabgKWOuiNAva
rMA5MBBSXvz2lOgWmuNr2UvT8sVFS2xNlUIJXAk1/sjPKe9cs/qp3xVeHcqw
Wh14Fd7fi1nrDFZhG/5SVZ9rJaik96W9VAiRW1a0hAIWdlNnXPH4BN4CIPOk
esyg3D0IzQqaK9fcTunZpQjuaLMX9YhISimEqldOFUsbt+BNrlbfvtBQKDRJ
j9gygLE/3viBRzns5DNvml9AnKfnWReWLnJHbUbZ16YNN3l2v2I444D70Kq7
j7fawVE0l4sUMdZ64wTTJOH/kbQse4A1lJihXc47URirv8k3MeJ15jkdlzEU
riBNKmUWsnd7LYMYI09dWioCR3dS9NRWmndmhLjb+6jYph3wDO+dL3TZ9LV2
NBHs88IE69mPZVbUgn+v5UY73fE1uGdN9JxfbXsXMLT08QTiZ47flK4ZZlkz
brRpzfcYuOEF1sZ5hPoOFjTvsznW0uswQvAWe9dEFiGR7Sc6fCEkNggZuLGf
VzZHWxTz3KMsB1Rnrxq4MVQ/B4thUpk5osN+XdczClyAZyGnb8kv4ymxlbBf
q4GVvIB0FWrW6iDlZxt0/HEmed2DXks+TQ6wOcB4az0iDq0pGTXogDp3Xs5t
jDTaKoYg63sDWKXx44MT85pw019YuwvkIRZaekc/YDtcQAKtOjEgWz77af6e
SnhhtlwweXPnrVUknQ5qstHD/fFpkCbVQUDCb9Dmsc4a4Zjy8x6Dd7ZicDPy
NGR4plIKr6DGm+Bmh+x6d2tywF4d/wLnm8qknf0lokKeHfGYQozIRGDE6Ooe
bkPl4Hy7j5X37QXA6Aw+JDYSzmuMd5YxT4oOCVUtFka/xLvdRoQGi2zXAHDs
lkvE8LbSvgTo7XxxO5mYRKJWXbmvKS4im26K7tj9L4paSNMhuoAwrbg2lHgH
qwW/fotR44CftJY0lIiKFgDMeUoqXZSO6kmqWJMo7WPfJTr1twf9lhHbiVJL
KHUb1wkLTGNcUHKQIHITFcma3FALMn3UcRYr2LI8yKJhoAqtq5qIl5sy4Dv1
7SvKx/8kII/XHAbJ9N9EtB3UXN9QVnKyJRHZmrN2EliOyiRUh1R3CPmb393I
nQCw1CBuWWriibilqakJnvx0rslgrpW0HmyYpXz4RpvQ79KoNis7WhiQiAf1
Pa0/EHLfHPdptA9mDHcL8yMcGPMG1dBGnMDyIZdQU46HRiQQkYpqKSNxbJkq
yZdHHZl9N9Yxkc3neUA77CpexMiMZTCfyaV/otYzpa5/o2V5FJGSWj+sZglx
O0LFxheC/QKoxh6qSz40yZXNcjXb/kHBzKDGUmoEpvpimIrBKBUIA1CkARHI
uIt/t4vhjI3IYo/TjMUtA88KL/cTic2arRNASmC2WoqCaD7dtNDrXhBUIX56
whS60K4y3F/cjR93XWIO3jolG1iBkzQ1YsEnMcoDMzsaH3s4f8CIgkH0e7+H
NZN9CN65QY6oQzcP98gEozBLdtektoq2ExZvlJz8ffklLFucOGGhMpJEnanC
JmcZrbDKS2YZ64VmlW8NoAHqw3jFl36SbyZ/aLnfv3rlQb5hQc0LD/fmH2OA
e2E7XbUzhcb/V0EWUDIjyf0/EfDC/pPcgotaGxuf4iBtpVJ7nULxrGTKZpLs
ddRf9U2D6dxQvg75bdAGgzIiM5VEnbDfzCcMesa4isOt0zYHFpJCyEb9Hkyu
8iM7xlmU/cEF3ZBovICb+5ejxeWzaWT7Bvqigu5G72YgwIr8vED6Z3YtlCFg
GWUjcCqV/Gs/Myw3/yUG+PPWxWXkU0z/W6cu6QgiizzpijX2HNz8RwXwI78x
HpvvFV7J4z6hy7h5ahttEBXX9PUcyWXdqBYOFdx/QGZeejYb1O/BH3+boQxC
a0JoE+rUWyvNJ+sDNpTlfTTLP8cKmCtydwZjSyoJP2hUYUWCj7hwJAshEsx5
3T+NgRbhM+84Nf9AypyWU5uY9nc25My6qNIygbu1YnUfRCbYj9wyLxwL8c1N
zAdBQdwJAZLRuhjxi+HonbTD8MzsOVU3yH8Lczb3STCSdro/Hk+FlDwquf08
CPmLIPGMqSa6IwHPlOLDXrTThdi6tUIHQp6g0U72Z1MhJZoYa06eXykNHn56
IJRw5xk4wuPVYyFuIb/x+av19MDz79s39k4uzIfHHpxID4o5jEvufo5CwgVP
qQUsFZgvGQ9nM8lpzTmkZ/uSu5i9MEDpDvn0FVI+kOoHCNOu/xRnEudDdadc
rQOzDqa1JS5wl/Qj+jQgrPnVOb+9CX4evw0JOxpsmNc0xN4NXWOniz4TN4BO
8H4XNFzEzNN8bYGWCkhMBRFwJw7sXa2QeUHuJiEG4EGDkklS6Er93LK/ssUx
gU+8tfogz5cDeGZFPVGu3pmRyrXn2zkN9jeseFVfHtR0z487T9N+UK2RCex3
LBhheryMyp7NXO3Sawb0NZ5MZhGwiSGjA/4QDEiVb5cglrAkaLnbUr+8FykY
DGtxyA+R6ZJ4pjp4PYVDaPzU/+rKgpCxpfC3Z95JmzVBF9tHj8A0UXJPTyVQ
wO5MYi+kzDmIIDKuL8dGAh4ufruggVslLDQjEhEKTecgpSpb72ge1zPqkamK
MBZVa8obO+hbrtdMNjxRibr145YmKoaKEkVdMelno7z3e53BKHxqt7krJ/Jq
HVsVtzuiLhdpbPlcAlQ/Y8zc/JI1RbdMURjTJz9i51iLW5aIcHgNu98LRiSD
6QU76YyxGksgPd+ALDgjuyYucYwwn2tMsJ1lj9kjvp3ZJGp4VH9iuKcFMwNZ
IC2fwkvOvPFAm+72zQcDLwSvRYsE2cmrOwdYoIyR+82xuCBSAkE1eEFHO16s
KVmgbE5/PXEEGaqSoC9zg826Mt9xQsus0v8apOM9pbWVDY2jtAqqEG8o3YqN
p3hELX2yuWbMj1DVUAiBDerYm//HI4Ecg88x9OaWqHSFBEqsOhqAbRXLtGD7
K72amKM+K4IsRQeXUDDfJoEFvaPGQeFskFLCyLb+wMOAxwG1nrJpb168Auul
hdTu8drgTUz1PU0XYAGral6lLqBgFV3bjaJGw7HDbbMMRsCS/EteU+2egd+o
6J0RK1sky2GPtUsBeFC58HOCeGDc812oS8yOf35LJlTODmtWDQtWaYjHMB6q
AfjVweRPBRrj9oy80//dFB60/rOYbKIk6766tyks+wZbp4aRB8l9CN5KOkPd
iC+PFtG0DBz02IUS0LCoU2Q1hakIoG0NUWNWdFnJemVsKv6Li3tNia+AiiwX
yL1/Jk/wB8Ay3qKpzI2z4EPHH93sFIG1aorKzpb1vQvqyTJQ6qblbWSRK7ak
5X+BHCSQ/rNdZ89JhqYeNVa/skc+3dr5Dk1zKhq89fkirVNLL+pjRtYkO4EN
AeHZDh6+HxBYIzw6kyx85wKY8UG9nH+kI/oaxjEJKw+d387J3VV9TOpOnp+T
J8pQx/nIMkiHIKHA8Of63bePLhdJLVoARDTPm+qqArT1ZDIjITVAUHk5hYYm
k9KB4XwzG58Zj1gUpd1OfKiaQ1S0XLDobSnUPDPEArtx6N4yKJcmp++0GEHL
o2+9Jhq3f40og3hHhxI6/DCiv65NiHsy5s+1Uv/UyG+c1hpD3VEsai7A9EgQ
SZdU7mxrlfykrMWnIcu4Jg4E3AkVX3BxWiC6PXT65FU4+Yhvg8ckVQnVbxhw
LQRbYqpqEh+8q+5DsrMliRULbNS1n76NyKGZKAYzmpV8DiTsvH2TOZMNcog5
EzFrxnL0ar/6xrJCHuz/qE0e97jlc22SIKEAjipDjdYaCHAImYhe1NpbOmGl
3edKwvcq6YCi3LVYQnrTtR2zJKOamfdaP7IFXkJNh9iosvqKNbvhFLOKjYfK
L3M7/z89auIpXdqUiih6ROQg1boKVD5tkYR31+SqseOCJIkG2/AdzKZ/k5n2
33uxK7SEXq0pZK0L74+t4i8jybLgebpBx3sajiOnvKxlp4+cesB6usiXECzD
xWNDJw5DVjDVosWPp+9pmloExaLC9kknvZ9LRCcenZw3epK69Oh4UHZuuSJ3
ZFbazqYE6GMVTSPj+l46S5WNa0hahjEX6k3gEOnBY3FD8NsDVdMtVZx2ETe9
8TXxmWCCbcGv5AE8B5jQsWKpulF4hDo4LJIvhNnMlfRllU7CdFeQJCKSJoGf
ajFPgFR0390MFI3zp4Yxh6yYUXox+VsqWQ0TZSKRyyV//mlE6fBFBKsrlhrR
h84sZlt2rIjSmqfJprLLKGosUR/7FzQbTCibNKvMl0sWxZNOmsrlR6d8Pe7r
2XkWyRpwCxaynZOouDLkwNvmueIO7fXF4aWGYwZjdcG03OYYfejLYXh5HGOS
+xgVZKPGrCvX9Tr490ck6mIgxcKpbSaGcHZtS/Lt+wAekmwZKbxaCpdUwYFd
1VfOK8kx85G6Kr2+85y5M4j2MrJ26denV7NbT3VzpmR8diBUFH4eeDPeUVvZ
ApzCry4kWsQCRHFD8EHoS9RePYev/sKYDn3iQW+G1O1ZaKU6eaTJ5rqaRdAb
bmHm9bdibDOMcEZy2DLzo9Jl6UnByVON8Ck+5G6yJGsoaF8dt8nO5d1Wal2L
LBUMqeZVWLhKtom1srZFCHTXB0hPX/1RqVkH57ActtOTn4O+/9fZw/XPjNPt
JSrGmHQVVrWf1zu2wixuO/WNILxZBWbSxMESAf8pa63O5JkviXIFA+yHUuWT
OC511M/qen/cqWYrvRrmADEjVRczLlQlARrrgZrJ+y9qIaQmMQ7MN8gHnJad
gLi+IdnIFBeNM3rrH3Qj4cEM5O3VcTfuZxbONpJzTE7n06nyN+RQsfKwpWwO
Ieq5QEnq/tMS9Zxbo0hTjhv/eYaW6gbT8pA2mns6coNv+j2tPHgu16mGDW9A
Lz5E+g0uAd+tJcJgJLZLm0ohTkd3o0fj1L/h2fdda/Ztg3e0PYmMip8T2njG
Qt0xMrnNjrd9UI5fUBvldL01WIa0IY+UiSN3T6wtwxawXMa11fOQER6spZMo
N2B3BdJkks2Od2sFOFh4FwcdxzeK0z49ubfjkuVj6KOkVTbkqPJ0xr2IDX38
adeCywhKh2Xsd36NSBnOp37q7hudcqQz/lsDExeh3SucdlLLoEf4aXNNptOH
S6y8Furez3lymKUoSxr7HSEaHNfGzAEzP1drZdS4OltZ/DRxxOXtslnt2o2z
E9LoJSGBrDFETzHbbyMQ8VAbc1dZfmWL5ktelyN66WPYhTZEZV9shzScEapu
Koi7YBEmgYE8fOuVaK0XpX2hlrH/g5Lc31BRuehJS6+37bo2DG3IYscxc0EG
vb4KuMEFncYYQnPd0ekqA8YkKBBbJfEzYQp+CfXI4e/GHNzgOhRw3WtMNyot
5pdE5X9JYyRm0iLg8PGDTXDkM8AGVPWqcDpjg+TbS31KHiZNAHf12zbH1wUE
kZ3GA4Y6X/Or3IfrNk99lkCzqbbwNMnKYagCzhC8HyegFupAQCYowNRgQDq+
Ydg3Q0D1++6wMFIdESZqen4vyHaw2UNdKXpLZCHQDFvVVMt5sl/dr05aldLR
1Cb7QAlkgiXqhifOxd8NgYTX/nHBkCPan6H0HCb+U1UK79I1R0PYYMkZr11L
fjbdc+XIlgtdRk8fRe4o+YWUpxnM3W7Uj1FXJ2SUQ6ZwJyir0i3O8LLUWzel
c/BKshxHtYsPR6dtmSP74k6+hrDc2DoZshlWwrjzNVrzdHaNo3iDQN7eDl2J
GGWx/l4MjFr85b/7jgIvCgdj/iPRmg0m6D2VeoAe2mVwyQcAItHSzCa4TpbM
i3Xt/4oNxDnfKUA2XDYNewlmmmsh7iVInffvyTnMW2DIR4W/WMMayv9PPDye
fIty8BgRpSuI5XZLKcrtHPBmyKgeZbb6JULX/TmY7dm2UZEQkZ8cSf+tT5os
E+sX7Eers+Y45G2kN3a3tvu3H9i20i0+fL3hLD1BkiinnJW9xGU10+sCpXfa
U6yV4Sed+vGXd32bRINSu+fXmVlD9LhpMC+qw29NVi+uV5g06TrU1g7nTSur
3Qd7GpKrXDX3L26/Zihc8t4D+Tg4MutVoicUTyGvxu06XP5sdPJvnfRJ6XlO
fHMde9iU3REtMFkYhTCA9b7ilN604slPX9/6MxYEpFtJteJGD2YOP1rugoi0
o71IbFvzYxFc9haypelB6GMY3tx3rQBbfc5ka0xyjk39lu1GhhdGhHpgmUah
ixi/L6ual9vr6BbpUpYV9w/E7JSOoxyMVO0bxNcP4Odq59UV+tb7IsXFHpQp
Bvx8vIzSCdFtQEHvtzDYTDtcikVy/3BYCnrEoGAgoXbr00B23YxSNKXTSDnq
hSOS68xBlagoSBXsw3h9vdo9gR91E6tEvIKG+Ih9Lmpg2xP5zVJe8J3rVttv
rBaiEfO7tpy00fB48Zfte21QJBFr+TvAaLXeGlq7GflPG67cuUd589KpLbxU
SCeF22N4QfXr/KyHMfQB4GbVK3JKhT0dEokiScnmddoHlyElYfmPwYy/uLSF
n6Z0IBiIBXOtPQRx5OcQH0rSDW7Xd0yhDaDUe+7Wopv7i52cqNJ/1/ahQGrR
88G8enxrGeL42j+a4XTLQX5Y5FexjLqRZBiTwhMxHj4+1bsci0iLx1F/ccab
SZZhPeNA8PurjQKodqN7cUh89C/iMGMKyNImdpemMIGk0bvojcI+Ny2Dim6K
8bN0Lo/Svu83/NodhwPrtDf8ceX2R+wq3ilpPdqWiQ7HvWaTeWDnfYFiZLAy
GmqA35RHHH9gUDdHaeTmJuF2AeCpzgzjNAJ2/30F1ixrH9rcD/S4Pm+v6DMb
eeZB2luuwSiQh7Y5VT7uzoin4FczQzkN8Wf0teWntuwwVBK7jWysjBLFI1j1
wC+4Cm1tHs1dHQFJ858HA6dBTQpSV7MYuDToTAv9KIIkemVQX2qcmxWqakLf
W0qibTDNpudE00ZSpt9KjfGfUoUMAijyug/TVwtzv1AL3TKd/5rgQ2QyooTf
Z2oQdkRDOdSpWZaHhUOzmPahOt+Fz1mdvs/+NzIW+XQRhyzS0/LDBTb6Pg30
V3EE1zIRwMCpEMXxv7YrU+/fahNshKbj1eEVWdYYT2HTA3X/Wzj1TPzgohn8
GyjkmuOR8aHwIGmIDRLMEEBPrHybueWCGKgoq9wQCfdxaHTXp28sH9gmvilH
cDyjWEyiNVj05Ij/5h/kHgcDSVjGcTCxj6daTUj0CLnQ2NsLGPre1DhWFYB4
Ik+fMhxIwYGWFGqq6vOVbsqkfSTLXYfsRf6XERKFNGlvDhdf7VURHZvG/OXO
1hsUNpvq9hYtMzf3bCpK5pMveoMQ1O5Yy7jYUKBM+oaCtE2Swk9ROQkbTmo6
mViXDmEy82ZlScWvocph4zjAeSVss0Yxz8vs617nuTzfYItlXbCgweBi49ym
4XavaDzBaoVgXHNcvEQ7dZE3a55qUOZfeOCD3NvWTbyx3I09puwrDuf7Olgs
bSNTTtG8yJCaxY64OnylKhOgsEvtkH307zlw9ErZrhowQmh5kkro36PtE21c
wW7HMHCcKlnz9Eo657ZIDoj6jTVH1IJJbQrzrLp//sB7VIiQ89wJxWEtd3Tw
88XTgGxfuJI2fTZI12fROj2UxED789BghEtHqYCAyPkInJsdskdUwVNw+0zX
Wp62gtreuchvwefBEdVuWb6sVeFlgTKmyunbk7gduWRWzxCuo35lBhEY1LES
ZS/Lq7nPx+ZiDfa2Mk9rU+ebohsWe63zyz+N1XwYb3uKh0ycVoIoumdIWX8q
ZjGrMN7BP0F5Qw4y8qfuajNzedhhM9W3pEFvWR5vFSSozYPAi5obBOFK4+en
ajHLWMo5O49lm1U2MlHHwU/mBADWKk2DsRTDSw1VgHl2F2/R+Qaexa8qdt7V
5L2gLwMkIwewje9/kacUx/lMUNVCcEa+ueuIpsPfcTjtQyHfy8La5HtZqlkM
mYMpedvkRAs2pucdDAIyvIzl6QHNioNmXg/j18LQD4HJRhBCbW0AeZyBrC7S
Tz3Fc93bbkBMmKdz0G9hdWkgfQmB1bbYc/nIdUoB+sNPy00dg+ZGF/aO1L1r
hh/fnU6lVfSalWPWjZRTFdB1+adHCI40WMGKV7vVv2k1aD0fokrSX2TmCubl
brodFTDZsRKhA/+i7xD/AV01Qhu3VNByOIpu1DzTTftMWkO2Z3WSIoRNXPg6
SzyGnfivDcrZPnVhgkZPK5vLFBWxIOb2Qv2zOrsBL2WEhwxJS1narbhbIQ+q
Zszweo/3Ztr9R7G2COWi+oVS8/sq4KK1Ipe2UBrVbQqACKeaIHwki/9Aeiu0
sTykWlduI1tZ8PkZyGX+vG7Xzg9kMYZ5qcMEDrLaEXuh1502yy1CmcxdsJNI
/dJriBxnrb8z/87feRjQUvcA4a2IOonHBf4SQbvE0PvWnUeKN9HJEjwTKLPH
WEvhwpadsghDCPmZZ12xhzA/z2dUiHBdLuirBu83JuHaZzMppcQUVcEmXwsm
awRAZ75D0FCHrF9/Tpcc284a4Z4U5dpWOiCeKCIIAnbIhuK89tthGJDkyhug
2CT5Liqhc+nURvs+VaRxGlFqK9qsvc8RXDbtFR+Xy/ozmjXnn1T3crs5FPpu
O0QkUwXRS+Ap6knTYKUh6h+dWGP2Dw6Ymd4YwfbHFxXq+KJkxdT7m2uFqFeY
InfBPlXr1t8JfUT2RUNyBHfaIwAVb3AhXO1AQ46DtsleazcCID4lPSkKQ/jt
VdZBjEyQRxND7jy+vudEWuSpzDbieecSgEL/z5XXetjd1en7bxEiyUPZtA5l
OULCnt6tF8cQmj8hemR2dHbt8bI5A6YkVj3le1nFeSwYAYydM77mW5VhsW0J
mVKWH2TncZ+S/RWSFS7tCCc32AlmetUZ8D3iFyVkvwiT3ZcTC3IEzT8Hg0qd
A663u5ACOGhWP6sysM3J95BpGyGlaqefTtdcsU83pMrXG+hKkmCOk+ENEZOj
vc/N1Kwvhk7VOxu3eqairS1w3V+RrH3jKP+gIwrmzTfv+ycoJnUFKwkPNMYX
89YwYyFsCH/PyAikzAmg2RmAdJUBf1sG5RNuYpq4gErdKd7ACAjDrufWuYzB
qJ0D7oenIv6thKP4FhxopO9QWtXbbhGTlD6ywnUJs6uC2zHc/a1aQV5iAoWA
dHpRZQEbPziwqRkz6QqAAhTxPwrflMQVZ22ETqig4914vex1EKxMDG7aeV1c
kFm9GX1KOPlvvKXjHd2mGCVdWviZ1GfraYYLEXoWcFXMCJO8Llmcd+V8lBuh
7aZXikUQMeYjDi3bXsehchrPR1EOrmKUeifzq5zk0IfApzXAo78MeSZQRq3I
de0Lcta1U99JXMEad427T3bCX8CCKtRSboqMskoqlz5knJ3IQZIEBtBnl95G
MhYb4P01dhzNDX5WKkaDqsE4WosNcrVk1Oviz0llq4wIOKgK7RcOUcscAQZR
/bjHaMNUmS4F5rZ+MrkyFDRJTfhb3XPnRGCqc0DORZ/7KcgTR4fAIHnLElJU
6KZZV4JcIkW+9G4R91YNwTvQakSVLt4Y+549AO2xQoKayakrJRJDiP7cEwdZ
UsfrE3PaPiXGWxpqzs6VIxFVyNwGwRrcAKwhaQS4A4KX1qfBrmPqKCgeut4j
e6AdhCd0KjRaRmCa7br3e3weCLj3fAiZifGhZ6yNzaX7quh3mJv9JFNUNgYz
YIcb3BpaHMEZpCiBVsE7AdbYaEpeZ0aF1x6IJX3jGa7sFueCfp4bOFoGRB6C
dhNhQSSimsNUFJHReBc9oQ0r/kY0I4Lp4ZvOIuJrQnGxX92yili8PeYBJ0mR
bzRbxNIxIxLgP+/t81iVtOgyXcJ8/GEU4UcFoKI4Nnzh2m7rQChzSR1WyXmL
Z4DFQzCF8t41EcJxl0u1PiJmoYR8MjOQtCDZA7lToQxlHiLL63+gfPTwWO1O
QH4XgLEhThCm6qyegTvplYdhvzMfdIszX3nxJyTfJU1URdE9TiJ4MV/J07+w
ENUetZeEysHs8vPq8eFa7VpMi3nrrXPX9V+6SLBbZr0RqHy/txSHrOkFsQ67
/lnGFsqMEmdsiOdxtAU9tEoqzy7/gnzK2vtia8TB0uz/ys5lqezDm8NGO7vf
Ufg+ZRrIR4S4iciLUlRDN0Gqp4rLjQT2i46QUiF5Zy9cKe3xntbbVafJcbD6
NajZYBbW3BpV9OGHTda2OTYlI6a3TJCEukH9jI2dqDLx281MDz+ozEPrRnCm
4da1wc0Jyexlj8n7IWgTYOT0zKqQJDhydM8R0DEP5KeCkCBjM8fSIkDD3DSk
wc4VY/H8lBToHaI/ip55cS8JKsdpLyDpvLcyLHYtxP54ayzU+Ms19AHtxrZu
0CQWnjZjaSHGn5tM8x639zSPmEwmfL8CltmL+im3lFAoKpxunVl+ovOaTvLD
4kygcsodXe6j9ID3XSesPtftmFZetXMUcoXEuSU71NpzEa1Oo/cZ3Yk9KSXe
bCSI1QkRil2YlaiInRsKyL23GtbXLVsGgkl6HP9CsRH3qmj/T6+2n4e+jBir
+eSBBy87FiWqzRDj9Hg72M/V/9XoTrVueiitilUhkwXexonqWsC17DC79goO
+Mk50FAnVsn8rt+YkXbJy6lWZQOJXBlVYOmOONRWKH4Po9ILa8rdJt7ML36Z
Qhcti1mTSnTDwsUMUEh4QuVy67/yIPT82aQrJXVjwkbzVw/9LLgUsw/XFCX6
u/gGp+7KEe9P1Y3w0uCAT5wztUCb93PnrmCdCLUx2iNjFVEAqJayizM9/b76
cFCm6ZIx6EBTAsrlDyo+muGaOKRT0ALmHCBRAfPpW/YDUnGA7I9G3D67OIoY
omswQ35cggNwal0uBMNoYIKKPZvEzqP0Pjf7YwrXZgsWn6Y7t8OE3KmVCT05
pkvRV+VoaHgEzAXQa5eP70AGHit224cMPs9BDYpBNOGQPbGs5apnndWS8Ml1
CNgAF3zH6YlmBMZhA9TZmY4qWSZJHIQ7RnuC7/BavQh4MB3NxaZFFNzKTWig
m2Ng/Gc2FQ5TLrWSeBlGzIaVROM7kj+W1v/pmv7r7wwKDY0eqsKzLMOCBuuu
oKKRIyUzT6knigUBWOmTliRJWU3Bh53TOdCdW6XC/uY5Q4O1mYChwywAB1p7
p7ylne57XDAmd0fIdHSxZjy03GGC99aWrhfliHulcPvkklVr3p24M3gn+xqM
ulAlz5uFwAeJrfGj5RhsUZRq4kNqbiWbjVB8W7V8Sx7KEqX0WnO90Hb2gbED
LWouWIEcNU86TCfCwFIw6GiCBmIZJ1zzwaOYVorFTzrKSexKrjzS4TeA6wMY
wCWCRt4zTXTciR8M4xgfPf4tORe9RPCTbd4NY9xrhe4unofDJC30gEtv2bAK
j7cKCHHeb9Nx38Q1pE114MUrgrPVYFsVK7jPU5N3EC26ekXJaNn7nHomqeOQ
Po+swzfMm0mXTRg0v7fQ0Qn1iLDZw/DOHaPDzjclLeD83neY3hA0kksJd75E
BqEFmoFlXIof2OAxek/QjVneAzFWLcLoJYNWKLA8kt4YJmQbpQV1ju1WMRbZ
VD6pGBLTDPSbQwvWQfl0irbp6aD1vliXWugN2dkgQlHO3JLuvYVJicy4FiK4
ULag3ksxyHbT5jf/X7BwI5B8EiVsFTL9uVPE

`pragma protect end_protected
