// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
tlZc+XKe07mEBWlmEtZS3f0/952KIllLrV9hJvbADw5Ai5IbH/2qPMX4RH5G
nuRwwTu6AvtV2qc0u15DTaMb8sILCPf0lrSR8xYYTZ7VvQWp+7nFrBATo+KN
X+w3i9lJ+o0JB0LZaOn8cuio3wZrQHHYVwmEkrf0qfBpHp3UFe6Cbf3OxAK5
r+IheuCPH2N7zcZtmGm6EVKhT4LqnP4tr89d/aH4tFxaPPCg7MfSAWhs06p9
v7qOVkgrAyIRMkFK81NOypun8HjXWYOLttjMxyuoQmyMdkmculUD+p9HktsN
mL826r3UtBShCVzflsjNPrSOUvGByDc45q/dgvHDmQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
po2GbpWDOvzrD2rvfXKdKQrGf7W5W8jMc6068HyLs+aPPCDW1mHoUQzB62YB
ZW9YkwK4FRLUpAzdm+ceZdDvRrj7yEQu9zpq1iuJ3vQ1aNKCRatWSiQ92+se
uTfI8t5FPcpXSscQyG9/dj5gYfsu6N+T972/DDjIKQrFtCfa6NjzQ81w31zG
wxKR8VIq3GeqUK4ZoJE5XDXWAsABs+Y6aEv1G+tkmApvQYSC/dkIh6mC95sx
wq5nfFxS0kOmDWtor0SHJDm/qZqmSIlWQiyB6K06Ue4OGcC7Ka2HXXbq3BtT
276dVrMqo8hQLJa6CW+BUpcPiOB6p5rWLxBXrEmooA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Frbd+s/JpJfkKyh3CMHJ0/0SyAPUxY/muNWzX8PoZH4Cer1rOq6Vyi27CacY
nC9ukcugRTxWKBUhk6TEg448NRz/Hk13I8/bkHUDMi3ZucyOKjxrRQPG2N77
etnLQgF/9l//PGMQBT4AjXFX3hxKWQ9KYvD82TIp3rPPzmF1+M10E8REMRUm
+901qhnyYAPFPVDmb/ec26W9n3TvvoYxUjSrUkg6igDqxGiAAo6ulVboyCGm
i4qHwtjKXWaCcsXl9rGxiNVc0qVmwih3rlm3iMxwV8GN3HMf9COPQ/SfUqtH
e5y8+l9+Y9Nu7VQ7ifVtvMI++xzjxVuDUeloDadAYg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RNcX3ODJkbWuWbmFY2/lxdAKZ1tkgF/LSQUJxX97mttuASh4CItk7XLrPrMb
jyGXzoMsW/4k6sAOloAAEmETlCdAcfj0Gc2Y68ENwWKwbecZHr3Peark9SY6
fGCGzxyRwyYg2oNLd8SN4AnmJQI1qu7fPdcbxr2VSO2PNUyezNc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
sq9athGaI67ERgLddh/krgSagr+kFn40WRyAJIZP0l4mZ9uq429aHbgp8Lb9
LbC9J8qVM68j+Y06aYUJURJcklR1w0BaZFor478PZxDINu2O3hhtA2bB1hfb
LAgVvoY5C5PRvkzVMsFM4T4ehs7zQ6MnIlHrlfHNzLkrNeBMSeFLTa0PpMP7
625SbAXA1CeJPrrIru+NQVhbxgDdrLXSksmJ7vULQBfNP/D/jVy9hVFZ8g6l
EkI1uTH4icCYbRJR3sBHsTHaByKyewfODONxSyuRwbIzniiXgKPmF6AoZ6vU
q6IO3cJlYwYdpPxqrnPne8r3jRxkKpQu8vfqDjsU3ftZNaS52I4arTrPRTg5
uD2Y5D8Bglrd2P5ewg8ixZRWnsWWuE+qbWwlE+uX3xpgvLHMIYXj4NE8zDrM
s6wriXm5PTzk+814tNcGHD+zp3sya07NFr0Gum/yXaWLfN27AvfQS3SQS4Pp
fpJRTaFlye4EatuvH6oWqkmoHLHRCKyP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JmhAF0Z3A7pLF0gyS3DwCmKXXG0JHdqKVBOg3s/ua1QKkQ78XlpsKViGRO4+
aDEAEficM7JJomZQIR5tLbKNvhiewuWXKsCLDgd97+MA7LleB3P4AH3m4k6e
2NpD6WX14OWUvKbm/DSZJDky4r+7jpe/4OwlgG2D0IppTRxIgas=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YZzEQfLV6a/6MCDqmeDxq3nnbeQq/4nNOX9FDrfK/nDmdyUOTPqE/ob0+EiA
AK0mhpgtmbFnKuNwC+8ogmAvJiMm5jcC9TvV2GFIIHSTDGGebBx3lb0qFWof
oGZtv1lDsArvyU8ivjMEFe6sdmNCHjcebCqjl95YGOZ1qYy/3as=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13840)
`pragma protect data_block
ysJhenFFWy8Ju9XVDDZrXEyiXh1eKMLu2rwdU2CRgpM7NVDO7D6F0fdPwVcp
cLl5YijFJFkjeYiO/cpsmwjy2K0Voe/YSBWnNrJ03qLrDaLRmS1YWJ1ESqzT
mrbl552nq70sJo/03oOfPbui8O51uxgPGMfZVWLiaaZsAhyKj+O0FR8zdvMJ
PMcL6zGyV7SmsM1nc/+HNjzRrlArLk9z9bd37IXTAjE6tr+uG6O4LAwaWfUn
oVgdEWsJ1wYNuuv1pfxRNlyRmLNnodUuwy8A0HBok/yusynYMEGE97GaSmCQ
TZKInpAY/GwlLAO4gU7lHql+LQIX1VsKM9bf7QB2ihihBIpDq74WOcP/Fzg0
v0Qt+ioWtczuk+AHp4MbKDbP0yTLaRQcBbPVEi/4pWEeWyHyqOahBCp4Kck0
SiJbrM7+VxFP5o+we8atYZ/yEWqDdpPX3z86mmQcFlnLYIG7ljfTfum2rbHt
jN//QJMJHZP6gH53Ky5AKwBGuWz+Wo/pbcppUWoW22gLpNQzXw1HxDx+Q/VF
MfiJE59QNOabKdKWNJ3ImMu9I2/DtmZaK84+SkFmlbajusxUKsnfK5s8MXgL
5Vdmf75KfHvHb71SfRsJWbVIh+poOi3lg8bJFvWNcnFrZxKi1ExTKQ4YUScZ
6bOE/Ijutkz8XCs2S+7GiTnhihUOBvCjtlUNlhsCYE2JVWEWRmB/MdClD0lA
VYHQ0K2z4qPM25/yj4KO/g4dmoGej3AyTtmgnFkjxjDZX8Vo29yLdwhEPU3v
q3M6s68+jtFz1pWFcd2/WLSP3FgN8DAYAmpj7qzbHpS9DtmudUgDL89x5hjM
RIVesnidljzvsZiVmwWfuwy7jLsln4txWT8++Qz9viNVJ+c0dnpYOmscYSz/
TaedhkXIe7RxPAj2Kf/rrLhiyhD7ScPOj48NSN24eKJufAjcV9xE5mpedQ6Q
vQbVtvYHVIogfPqFw1z1cz6V0AlyGsZFctYa06nds6zvf2HPA8HErH1cYRtL
g1mlwrwCoskfaizvqN6J6bDu9pOlwO5fT+sk+SEzspJZBvFsrPqP8KMR8jBt
Krm8XXVBlJgcxvTJI3XG4n8LXgv+2ooVPTt3e0rmuJca4tSVYQoOeZTWfHah
vB05+oGPqoqCKeFXL7JOXwhVCEnAV/Oz7iuPXuirrV9tahJ8vfsYWZ6qrEDW
KsP7qPu7dizOYWjQ3Ljm6Dj+O2yQeYPkHlkE4GSHQIAAw5FzgoW040UkuFo9
LdT+UewwrCysWcYcWr4XrRQazgZPXWZcv93mDrF1I2wTdLR4Tu3k5jI+qOLn
RNtMvFOcdkXDC0n4i63BlkxYOxRlEcD065+DWzDIE4/PXvB6kbbkAg+SiWQe
HvV7wsPSr368bkkouwVrP9UdyrsJRfCZEWNrNggsxegNWnmz9DKOPK/6Eq1E
8z8ghhBqDcLg6FOH9a22Os6RCA+Xgk7a5tOlyTCBwbpBP5Hu4eERxIrrdbfT
PYOuN/0n42yvO9wY/+T5fvO5pRm1qSpdnH1ECXgkGiuuROQ4stFUvaLByCeU
00gyGog76e68XxsO5oOthwY8ZGjsY7pFwVe9cyyOC+RglEFAOQfdMVWhuX2i
ByABbP1ewNTNw1XL5QABCu7PHSgCiz80xkZOh8HOmwgAX3nLNzPndUWS13kd
fp7HumUVmrQI2yuXuxn74af8T8akzo7qwVKevzmcZ2wczwRWW64X+YEZT7uM
LFE0Ib67a8cdkPC2ZE3nkoCbHfa3UAnFNdMJ+dMKb3AEPnZD+j0Vp1lMYoOf
Zg9MyFdvHXIkefrTjTESgQPZNPntwEWvB+Vt/KKKzhnurokDnjhtUDEtZCV/
iKwyUuQw9+xzqyqsMIO4rDKJ4uMmu2E6WFowXyGPUFY/SJcK1Jfj3MyUkQaj
2XKuhubC45XlCL6iL6eh5TSyeuaC/qMYjr6KuC49q1RPuA5IYjsqJiXC3TbH
EhxKdht6LUGg4MSUT3WWILHT+16f0Gg+LkUBp7j7gVftxEvklupnWaEoHQz+
Sx86e4sSmirbZCuNvQhk0TTIrJlkQefd2RSBfhfE9P9moD3K4Ij4yqKEv4Xs
Q+Yc9E1+F7xPBp//K4iVox990DoGy01s4quQvgp4mAK02hpT79Dba2XhXwIv
f43JYVk/5auNibyY2QMNIYrEBv4HQB5cNrJQ3pVoKO+f517AHbLN2Xq3I7gD
lo4XkQqI9QgOawfOBtK/fLgPAy0HJspoJZQI2fgt/V0wAQ+HYVnw7RsQ5PQL
Vk6KJvYy6u5deY/LZ6/Gth8TLpuv1uz4T98E27PhOUFoJjXjthqUeTjD4v+U
D1dRwehxQUn48F07EAx1bUPDaA2WoG77xw1fwvwgQfOvcm39t1HCaldbTIjh
bhEXIbs/wY0iWQVlzvTrkJ5wwNMjtfUosJTPIBQ2gfERDHtga6KWFBgI48zE
a+WJH0+Z67JOMDZhxrb+8BSJfJgLtzWVwvY7Lyf9koDgGwo21JdgXbTwXBba
31rEaxWmQp1ZxVYcanwR1ororuS/YBCAict9Fsliy935C8KEqUoyKIEaXzhs
k2BlRgtsX31BJRb/o5RmdD7gtUYc66l5VO53ihqVA6UR9SxHS3xG7Qt2DEvG
cHNOnA5ZFCs77I2hB4duKe4NkgsGwZtnjy3/YJuXkVJNwE6ALrHbwExVvnCO
DfrvVb4IluaBLutgIqUs/N4E5xLL4R0b4TvFXB1NNpUk5Dx4IlTzCyOsy1Le
c7xPIug8GGI8+XrMZTsWZL3b0bFcN0JFXYDXWyVEatcJTDt4wTKg5tn5iFvG
ojFYEqq11mkF36/obhm+0ZXLtU+fRmoG36TuX3Mb46zCa6LEfItnkb94oCyR
NmMHCaIttSPISg4CFqLbsntA/TB33mqS3NM6C4Bgdm2sQAtFxoufvyDO8f5w
uhTiEJ35Mp3rIhI5fdJHQW8wzM+t+M6bvextCUjXbnPsKrQkSCVtkqyD0F/1
4FxFp7RFQBe1DjHxezI9mTmfh4ngttD9DIhvAQMHPM/OhiAHmbjULsn+Qvjj
FE0J0dnVY2U+piEQaPLXExRwpDZ6Xbd6huMJR9JUshmrgNdlgjtP625276pr
q07vD9+DrGkZCukyofKz5y5QeAWeTrFfnFp4KAIdljspyWsN/Wjwn53XB+Av
U9z6YY6Ie1IJDmgRDY89h9lminNILuyclaFQTWWm4sY6Ni5gOHiPGz++AxqG
x401Dh78jfxgH4CaFpfNgLd55NO46T+TXcEooIxsFTm2VRA05/5RH6Mm0ylL
NvM/7w7z7magSB/AbkDORcq15poPwpoDde0cBbyDdgmKq51JmX8AKZOXVi/Z
ieL8te24QtqJ3HB/ybV4hTerN8RqqRVF//SzoVrg+aAQUiSUkaYiJhITDcs7
NrH43N3iGbH9dcM4OtoE+wMIkPrHIpissxmEdFrS04WexWkSj1VdMmnbEm7v
HuEysFR7LitLQIsJdVb1LFnjktuVrSaX2nbS01GMEMDhcC6BfoBt7XE83hdw
Anzi6OjlczP9MNcKxD+/xCw6NRvCGnd2i4HR+fMiiCxygKghRFzYg026Wxo1
NPsHv2z/ikHaT+uAHX8MLbC/gMr6uTdwNVeie74qBjSQn/2N9yZMI1aV1/Kq
UFmTtC5D7OpwaJ8gJbqnkMiv1dR8mUmplN230nYnpYBAE3F+3TkjEq0yAwfS
JwMv/hbc72ltX8KHq64CALnaqKcxAebVZM3lcc7KI5SJ6PQtYAVObAfwuQOn
v3sfbDYlZujQJ5UdTaRKLZXBuPCBJ8DhSfbkN3dpyAO9ce75HxL4bDumqCTL
EwSlrKRw8GSXh7LhJng6Ofk4dfd50/Yd3BHtBHY1IhByTn3qe3MGl6HKQALo
TPJazkDQv0iYq9RQcv1Ovp9eqt/AisKcxMiuW5AebiyW0UeF4s0FpDo6Vw7l
ZOBLmN8ZeVYzpXBh8e0G8Jlg76rmkcpfi8hsnb90FyRdH31VKH+yw2mz31z3
uDooKfRKNWTLtNVwR+150m2xp1IGblC+2lAPwbUk4csqsH3bgaB6qICCIm2j
PvEMEyE6lR2Zj0HuewNJW6eKmtLWYnqePH0IvNMaWrHewEHMojuifXgjgkjQ
Uvf6/ZZzPOBXQ+U/HaelBzKQXw/ddFC2OJ4A0m1C2JBLGEjW29Exq+eAQwOZ
GRgZrgNikdOLx98iTKFrcknz94PJ4Pit47i0407CvplAUtzAGDdg87VzcDFE
ay36CGl2AVQj7c6gSOCw9IIKmBb0qWDqU9G5r3s6BIZVLoxS7RDIed/oYB3l
Gqz/n/okzQPSKM4sH55hc3URNUBCer1A8GF6F0HPzd19DMwEO1b4nndx7wwn
UtK+CjcK5NVckdC8ppOtOP9lfd9rINJKjzj5VpAzpHCLYweS/rW+cJP84vSc
sQLYqdzApuSkSTnS4lDRQVsago2QVlLm2l/5DGvz3/1F4ZYTgKPEinSrrzEy
k7HTQs0Ik4yVL6bVYMjh+kEYcFVXUG10RhKlHhAZWEq8hl3JSw6O65mk59WU
tOGswqy7+XiO0r/YoeyBGhMUl8TT8zSYWNoDix5yo5jR5P7cIiZk2EBJnU+N
B+7tUXTekuB+uONc6jkRRu0rPCy1IE3il65xzOGMiDa8xyXGtf72JLPEIo0y
FQZhv7sQ4y9MLchV/t11PMeLmdP+ShUkXABTe3+1baFn9tXPEJ7wDd8xNPnr
ZswoorNlbJD07ogfpdSaRVuXEtjtaxIyO1mELzohLq+7g0/mTeoX8SW86Jfi
nXjBHXdIMAyoEGloIHiGAVTgu/4IU3yfUtiK/57VEYKGUfBGh4fKVznwMpb+
ZexC7MRw+4e9esL1YarnGaNMWyOmjICfn9nc9n4g7a1K5BcPA2qSq46kqvia
nlwHZ9xfvr8HkJOVJrH5y4ItlIUbzqNKwfpN36a68P8nMHedsopzKsIGdsm0
5+vU4tLT0anBRE0q/QpLlJcCuw3GrrYGreW6zzEEmMo+uOiYdQ/MvsIqO45r
rFSeRaUi1FX/17jB+zCtMPqwaGCuxHwxWf7+Yqeu6+qmNEVPvWmUpd2iVine
0CLogwBfmLoSgL6hKrqJOchtf20vdgiUm+5x1pPrqo4eRJW/47rpRTDcDKoY
uf0s63EwC8KXTchhyO+H0hVxyrakv9eh2Crky1bJxDj9oaEz91xnuEVt9JFY
9shc02oZ2+8XRl+g8gsJZaGUYJk3ZdeAlq9ZKbuIAtxpgeMhAbP612o/auwa
rWer8EF+9kfEHERPSrdYLcpNfBFQkwP6BN+eP+e3mrVpow3RI9U0MiANMsnP
QPHbqoTsaYi/NutTDzku/+8KtBCNhqTf+m0i80QTrfzwSjPL5nPyaG+8bRgf
pfR1QD775V53wdXFPonmPHnZSebP17ZGNvMFtUaZymRIgsm2QRCqjJl9t3Re
v7lIRU7Sg+DNELss38PIGrYZVhB+bqMn7FUhgWfmER4SylVl5UozATMPQyr3
UHjpI7eTO15qk7OkbAK33Y/8chE2AdQHatk72TZkx5SDBCv3QCH5zopk/63x
b4qh5DhV/70N3MYjw+ZBImqpgiwt2jV9ebA97Su1Xio+9P8lxyMQkjKdYWv7
ibSykSUs/9nRUlEZpx70AQV0IPS2XNABT8LoAjQbOyWCG407KVUj3tRTdlJt
nQHW6TEgdHjxn+G8BF5fuRlRbEQyNyuPzfNPswIXuDBQX71Tc9dyC+VKAFQz
ZgDS1jnC9TuY+2Bx1neCx/Ag6hRjk+2AW0HU0tvFOKRfGYlgG0y7qpiK3OL1
nFoI9lMLlNJurJftgrcn+0Z6lEnDoMNTegVQ5VFciSIykyChPywZR/eTFodt
0mIDQMXj6kR555Mm/ri7/sSyH/KhbZe2H9LM4KCysIJsOZap+DK14PpkLVdQ
ntUI2uRi7OkAZ9WMfxzvsEMxc+CwAwnW9wUlljf19Xf873CdZnitTl5pgsSt
nuN/kCa/2pI+oQU7XYaVrarxtXPWUML6MOb2fPqi3Q0XkxWyGP17KZoXWdqF
pz4Dg+N2KupY90b2jveKqsYdcID3RCohtZ/9otrSkApXcm3drhEcjkTWaLtU
6pmEU0bG+rDV+Wka2ryGrPMotVDFVh4LxMv7cuk00yjZMJgmBOM9ot7c0Apa
qZWiS290TpgP6bh/y/T7cp7gyhIf//W1KHP6vWHjj/Bqm9Yfrom5FXS8W6EE
Oe6K+KDLeXFqdE/nb5MPmijHtD3lplIJQg1sSFIhPKdpAX69sAbCj4nGwgf4
59akGYiH9UOMSffaw9mMIOnRogY+3ZuTkeyDhmU+fx5aPXJKu/6d3gDvG5e2
PAsDqTigYPQC5IS6fD7IdVYgjaub28Q5aEdCuELCBdXbP/KKKC246vkcnqoI
4tT0GewioFaDhOvV+quENq4r14a66rqRVT/jO4ZI8P49/+TZ2MRU0PnpQsxt
mF6BCLoJT4RzFZmDWwgfzRUdsHY0Budk7NHlCDWH3ckIERLY3oV1+O34yEL/
9qdfO5swFdXwpF9TfIOMdoUmZ15rk9SBr82KMcYHovBJvWn6KIGQfLVk531M
1EFeXAIS+IuRkV/A2sbFhJR5snBnzeLpxdi24J7y8u4NG7cAyGlZYLimrT1d
HIAQrTbr4BU/PXGaK8nG0FEq/X1k8h7+MYEZH8opt1eFu/XPkYcaj8VO7cmr
9zk6Nl0c15DS80LeHliL1ct2KdhEcKPuXujsBzVvJDfsYkdazSW8WHUbmTsc
EqTnXnWxNCBDGHe7ulh8qFTTAyRr7fIGGmVETeKvG/e7rrPq7mwYb/ByRjGs
2YfEE7ccLNlUYyVgHH/tCV5JUEBSJ+/68CcR+gIPL91BKmF26zIdUnycvV7C
UJs8wO22zrXd2vgB5iqEKpAOBszkx3rCJGJkFl/w7cq0/0NNEf54qSGdki+n
pMhvvMjboRF1ecFFyBa2+ucxSPwVY40vwDTQhr4QQZRt8gPOsVMD+ZrM5gGQ
ajXuaKrz4LxWt1xUOwrpGY21Ez5OcZWPxxmS2Zn+3lWWpOwip8jclUFWOmd4
xYeoUOQzxTMbgHJ23aZKyRoZuPFIxwPdo+CB5c8fg5yGpX4u+kNtxvJjTsdG
XbxypI6gaTDq0bDNsbYFB28Ea3ROwI/IkK7UvWOSdbv1ZWuB9rDKjLPUSb2B
30OMr55Qzpg7XtvW4qqgSAPOdoUgiKxmUre7e+Ed/VZq7hkFgv9827Nu6h4v
BdHmpvfW/nLnIFpWEbBg2oQ+yzSVcATmLLY2LwecZQ5xWKC57JqjY2R9zxLD
/vk6QA+s3Pl9X+2q0Re4omcuaSn66TZVd7wKv8vpRh3oIO3qmweGoFUf3aDt
r+9Ukzm2BofBCkBJH+rC66bLDFBjF5lE+UkEeaG/2BlentGklVBWzqw9oNZj
DAnV1Q9zawBWuRHb9W01lai/5L4lBfK7TMVdsVDCWFt27pqAkvTpWHNnViJ7
278SKYqo0+eGj/ciLMJXRvpdglMXnszI+dRbjOS/sBXj8kK8rPVFztdTd4rY
baB1CFK3O1UcPrLngLT2aiZWhkgmVSMEEl7wU7QjklttaO2nxhfJhJeUN4C/
nGkLclhI2PeOciVp7KOO2ENy8iDwcNB07Kj6/PoUeRa1ocTgdb781nLmswFK
lrUsOR3xgdyHUn2RgeLJqCT8iVCoE5QFSIPYOOzb/r4f4MfoEx/6ahr/oCv+
aiGAPnXpCK7VYm8HfzH/SuVycJK40x7ATs3XKxLlm0gREiGg0sss3xGqmrzV
PeKbBMJ8I5baQq11leL9Y3lgXSgQz8k4WoJKCtCGOqOzLzEbujtRqJdVOHrh
nIfLySBU3jbwESujilQ45IxEWby4Sz3MnU4JYV39XJAYc1XL9YQSlSl2vsuU
bKMevg4ODAJDEVdd5dxrxf5+yajFbEwllP750ouctDV/K3jg0vQWTVzTEMbX
AAte8ooUvp7ed+iXD64pEkrA+cziaOBdhB1HpqG2YKb/nuNsuLJ56HYUPGQh
/tw7E/N6FKA44mVZM8BMcXufTzwvh8heMxb6dOo++4YNOzf49w46KtUqZx8+
/uNk8D2KDm0zrgczMDjnwwma24AaYCSXePERvw7MfhZ6TYvQ4D38cF4x+Gjg
k4+Kky8iHTzVvHM0nK76sw6Ih6vHqqRIrwoSF6jDIFIgpMBiKS/I/vNwn6xv
Encefo/+Oosp3Nk0WFXg3WOBVZvNEp3TR3dX7zZkx/bJm8BVIRyXs1Wom9yj
zShfWylkD8GVN+yz8X1aPIqyW7VbMJgHn9mOc69653pj6bwiKVZRMq56s63/
amP/wRHHvon75XHqJ9/cKvuBDP5ontjjm2079yAwsk7mK0ArOjdvfFF11iLm
LmaXExHMqqJLlPP+OdEa77k+UBlSclKungXSSEIDibykjwtL6qEke2GPutiF
KpfdgveaKkw3iRTrVItIoTExjNNJQtIpCo+3h2UgPVOS0CeD5m3qS/p/pSrF
5nPXtiVS45E/toIXF8D2basKbqwR49KqxsJ361cNtJ7mugrxbXRfetLpg82m
cU6IDzXJc0E0LYEed8nJyx8hURCsn1SLDIwd7i3HczQ+zCQ2XRnbJ/F72fuV
yRkFpqkNN9CmGObPrMscThyUlXp3GBY5Pf1FWi8F83dWfa4XG9CCHXbk37cj
LmBdpKEuMNeSZy7in0zsAFfU+gmcH/x3GQw0yPRaq0HszECjlX7ZXvTBRy8l
pke2HPjsjRXHZttpWg/S4VdmBcq/q/FVItWS3k/1UTrP6wg1uBKWHP3ltYh7
+IOQU+5xX4j+ric5ijmP3obo1mGDE2p4w2VI5P1qEBOHp7MEsf1fTK5E28bj
v7jsPG0KyhzkR+hOEimHqISctuExIqcPfPclak/YXRvQyfFNtHS1PInn0um0
2U/q6mRb7FJbJSigTIWQxi2Yk44EU6YN7TbHQSjrKXPE44k8SJfXrdnMfsAo
R8dIlBuJjRX+hBEePXqNYP6jab2WgGaHhlz+I3QF9tXUIDZ6YzCuylmqJVOG
n/zLLJ02xQxNyObZgtmrb5zNWgFMLKjM1htsxlo4OadoNFBSe9wHV2coMam5
tsYdAbIO/ShGB24KvbrStPXTqEwh68ykOvyafmsVf/jk//NhLNWVUs5kX1Za
ZgwcjUw0/dU2QUpm+XuLrU2K1bhTl1Csd+UKa9j6E2W5k9Xf3exLpFf2cYGq
AiIvmmQ9KMdRzC168g+qwvHnwF/wRpfBeMeqUT8fGRI0e1iHk42isEjIsFgh
nzUW03Dy0UBnSk1FX2s1aN3X4T9TGZoStPtLfzl2wcrfxF7lCAKcZvfjutz/
9ImBkBPQw58fRCD3F/ozHw/eQbe9fkr5w7IRqYdUaBTDBkMG4LaRW3CaJ6xt
Q4bZvhCmeEIggPK9Rmbe23OmJUbcujhKjj2ll7PAUm0kVtg0AFVF3gkz0A0A
3XDYJwKxmNRXIzsKmej3wudlBydbV2a3Dm8cpLBnDFKr53G9wb+/nUO0qkyu
aIOTeT3+t1akcwKQYR0N3R5MRFlFD/4/kDJVE4thG9o6W5Pzw5YoJZ3LOpHd
oTknzQzT7TFbLKb3rE7Pf7od6Ib0Yho3RWknChBT2F24B82Zp7rEfIlP98GS
ACC/DBf5gUlWyv/DuanVBB2GRg4ng3RE9YuAVBTAy0ep9npCdGITf37MTMVu
Q0XauDgRvaWRN0MQNgxaqrxKM+D5qvzQkuKAN0vGWUAfAkxwAgQl84EwLisO
M1ggfPKfQgMFtKGqt9uQHVGokRdWBK14vy4TRG2McrGzbTJudPU0PWqZ1ksW
/OLY9dE3GyF6KN0TSFE7T7fC/Th7rOSKQmq94CZ0hhcCJD+Bp0bDN3+5xzGN
NFUFdUSZ+jaTFv1/P9DPFMBG+BKoZ0mwicQR1qBYnQr1dfC0oSfuWh344jcu
teXH9/qTQUDgo9UuK7DRxM63kJv9iDf0X+qjCKtB0DVwD2tJNeka51BUiERo
AnZ4fXOwGEQd+Pxxy2Ahw7aKeyoc3mNc4i+vRJfDkFOG95iD0V3lVdBfHwQg
5Nw8AGTtP3VZR8637YDtuVd4fU7NHL6dFau7UAFDx15aTKx391/K7/nNwgOm
y+k4li2A8uN3HHFqldt8FF92nK8V08Bk+aLCDzevomZ9O3KDXGEz2WTEvzPS
U774icL33jOn1wy01BHI9Hbz4jo75ePThGSKm37GOyZPPqIK0GADmiAf9Jq3
bXqvQinGOSfGOkWdsFVYKFH/xVsPPSv/6jqr2IQUK0i1Nhk2fpzLGKysrdyF
KRo7kZaseprUcj+W0zGQpNy/YpqW/2ft5dCZ+GX+m57xsBhchv1R8aQ/LSwk
ZuPmlbe1TbQKeaSOQlt5dB/AT5yLfKOAnIhVCam1zcMp/cTrs9Rf4M2siVoX
beoTUSLmA87HI0HZEBP0f93CoDw1MeOAe6vGyp9qxrqapzgaqmPcGatrcKMF
Dxau+b6AhKfEv5c/HN6g8Y3yHFYKjELmmPbFFrdh5jeyn0Nw10Xx2sM3TTIs
aq4FQ0ulh6sh8SGM6yU/ViaNeE6S8aAKOPKmroIuJakkfG7s3EvzbqoTqa4q
KeMvlsnPaEJzO27Fw60bPNAnEgbw1N5wdQKEQIH1ONtlGQ6Z6F2zG1yGtqIa
8PW0bg+G7VNa6rlsWmvqMt8T9H+lxkkL6GnyERZNavo7IT6ZB4ps1pjB3mYt
CSjFJ+tQw5W84LmVA/cIpJARIrV7yLDpjaJd9RmMUybSe/E7Q1VjnLVdrNVl
J3xiSq72ewKz2ZWS6CfvD4k0SVSMW7kLTUR64PdKGpuiIUPLr1MEcGHNcIZN
mtZw1Ep6kGwTFYJ5PRilCjfgZa6WwRwjXikKq4qM/lz7eHQzeOlxxNmfzm7k
9pKsI4lGwrOg+9QTq58nEtexnXs5iL10EPZ18d2y4gRRfeVVtcCyAtwfa3ot
DLeXcV4/i3FDaBBwhoeD+wksUEj3WnWo6WJcDWtUYphCIHEQbDWR8ERVGgRo
We4yyWu7hXmHoMeVIHdJM6Xr6eNDC915TD9sPM2PJgZcJqovZgvzy739AV8z
MRVcR9HGWKppxuJLzXa/YAgDKQY0zPU3/CCTQB+pVV2gEi7bYVxMnTIbEVgr
sdkq61cs8ypuXJqVfIRdOVUbGKH6zHhNybo7nkqa1G8dR+mFuwta2lS8UE2Z
4ld5PaIDac4DQ21YOH0Zq0e2MoAXt0hGFAYZC/9YVA6AJUrE/doxk7jlNw8V
NDgeTDIYMeq53hZU6BRgckwPkR+N4ijBrBmN2QGa2+CSOcSc+z2LKBJH7R47
xxmvrzMMR8+7QXL4mtcHiibRE84+AU4Io822BXsTIYoq0M6ybWd2tG4lVAYa
o0LSTyUlhyOA20c1/MQhg4jz8R6MbZjNyF+cI/t5AjPC/RLZvL3ma7g3k35H
9110ySuv0zSpaxd/ZYR6w2RG4sk/iJbywTLBVJyQpi1rb5OcUZ3ZUvfHdTVc
rzUJjs7MIpHDsX1N1eO5mYdlbligq9olNa0SIQOjZcKo0vWAOiNJ9+fJE9P1
FEhlnD+1SciWLzbipFeS6jsdUPQ01bv3+88ZPi/ILT5rLUtmSBsMJR4dI7s9
bMipH9V5rzldFVh4btDDaZIjfNejJNOzMErSY4JSf0XGwsMJOjLICiwKGJ+H
XENXx2pM660JcyJL+v4/gR5+SQIHfgWtSdiBipvxyVA0yjwMcwMK/YcSSZmC
BunVRdgIDOT5DDnisq1Gj8cE7BThZkX0FHyp3uofFSYe+1RQFd6pBzcmFFEg
c1yPqjUwtuKhjLOrsucRf2KNO94UUt5wIZGxARaBa/QjBSSVXEfrUybwEvqe
631d4+A+d3qHkWArDR2dxdwY2ttly/7fP9jBdZnqTV3yv8H4IwL5wvx+qRr8
wydIbrvpJYIqAFmb1Lj0tqRMOQglsTDSfVN0lF1Gojs5gq9T7OhrQat0MPpi
m7heUQxJjFe+V3z3bBKGmYBRQA9UblErYONYbYfTMiI6CwPH8tNn04Aiy+wy
mxr9hrmFNZF4m5DUOyeiTaNQYz55nzEgDitMqWEoeefaQNG1hRvXwNrBW3ZW
mKyJ9DEHinsMGaPo63noBQhdj5mc8evwMw+8lG/MPBO+wILPZD70UaZxLdFj
ms4x0tPDLkdxPgQub2UaA75zsN18PDOUPSFXBZGcM0kObyh8zRbgtZysdD4m
IyW4RlcR2KrCygRqsWM0AaZbm+4JqME9ZwsPy7onQtzZBdQJklcOWRUgfuk8
1Q7Nz/NxzqdaUnIO4NQOHoF3uGqeo2j47nNAOUjDorVo6eFDbWSBccSD/teW
ntg4vanz4tAnaDKq3UJSdd/PP1owAPfr4HgBHLp6jn+PYYIJP5ldBmeRGude
VG7/xAlZWqhvI4LQ4DUQG3n3Vc36nzpM9gQL+Zjoab2w347PgNyobwT9MLaH
XL9dEeJVRLLu65qJhtRuQLda7IHAgrQAkR+gMuG9hnYcGkUTfH8F1SVvOR3v
d32aP5cVRKj63VLTHggBmQLgA2vd4OgFctSgPyLBhV/n7fn1QuiUKvKZb8d3
wmZrNobe/tXCjQATeRoi7PGatPsqMCxAKiEgTq8DFvBtE1ufENXuagS7Otpz
Xux0vWSulqRHnzNhJqR6b/M4uWsTKgADFw1J8VEgRIyNcsyh9vRUXhrRmlPO
uxCQBElUWFCTcILeX5pM/TTChcFRxsODiYUvMVxDYGfMhAWqZcqemnVevmaf
GYPhC9bFm7gslt2NkxJkUzrrE10S1stIBviDRpJjtI6PGaapkOB4LOBfk7uK
AF+RNU/8TFU+4Ge6nCN4oWmWvrfOdZR0bgoklJhllwv6VNmzwDqfsZPyTQAu
jww/RrF+u7MlvWeHQFIaTE94HPz1cAnlNdTGRKZeaQmFhPWyyG9qoM+41jqz
YL2vJjrusP85ey093/eMn1vCALWUrMUgoZS8dfz+Xn+sRee6kKqUJjAUCULj
BmdzOCAyd6p5HGrN7SLrPQnljtQbVlgf98FBzes3Uq+xil5b1O3UgMoeA5/k
cCPM3F5mU1OyH5qmDnHrrktRJ0SvqEt+TirskeDqxkTvzrI3G0/w8rXTerku
K7l65ZyeDX/GszPfqxi61w3llCx5Q5WNVRWOPe25oBF4wOrB3jmiXeSo/yrh
8zJYNaSC/HoqspYvqAcuWBzF2jg55edhrw8B2e6mKi9XGlpGqt0tNB/dAv0O
MWUTbqhSgm72rMbJboqD3UPLzb6t1Vd8RjCsveJOBXOCfo6JGn+NlU7zxcIu
ERPdL7IIRTDS85rr/mwHtR5eKW2SesaLaCDT4lg3xOpZ7gEp5SUn7TdKVlMd
0pnzwntjxsFMBN1ZCuH2MlTe0pY70yCTRYMGk1G05SBsrPMRgOPLj4lgDmem
C20QWJZEuQczkyaUHfx9Y9PT+CmN193x7RAPgNlu4XOBZ1RCTIoIA/QGaHTt
pqgvaFSTc7bn4kHVI/QKOur1CHWJw5x9Mtw/d2L1yromLtQI/4atExUA9ll/
W4ppg4+5G+HRgN0Vo+y3nRhW2fyOTaciX3eaIxwVS++wRRJusrypIcExkrWx
KLofUGpPvnp2dKjC3N1RWGbCNglxwIjSBhrHTxCNGju6gB7GLJeov7HQ55Kt
gFSn2LETwUleOIKBGVulbleSIZ5pFNUWG9+l+HZW6isnDTVwNRpGB4uiY0xa
swOs4u/bOVQch9dilLZh+hRAsMjTkr+0opJTjjCWukfDW8Pal8T2VMa3pBHD
evTXbG1H9kKNlstYxHaw4k2nadWI9gqUuimi+1uAvg5BF93+EVeoe0ko29ec
XWQwE2I/4/7ELefb3bi8Okb3Um05CTIhXE1cmA2CsrFtELQs9N9/dcg1962m
jwRB5f6ObdxiHXFmPeyg+OO2ZEePN+lwAxyl2pnO/7TmeyCb6HMOmYKSZjZW
fTr//4RKImg0j2xnwLRZN+DP7XDE6zj6y7zOYnlb5481Lag2j+ladjjq1aHI
/FRjLuqfYI5R/cKF/dXQYHHm6fETLzTWHt20W0XGjzOmobK8EwPaH3WUhFho
wpkJS7KUbyYDJ/6DgahmF4U94TapMbnBZBswq85c9DwyZRXDjqygKz+jAFN7
MuAKaUOvyt9WyssVAODj6gftLEpYBSllL8m5lu1YM+Fbp8y4tD1qy/0BkRKp
ixUzckjTF8njqZrTV9E77GANAbE5CM0XUWYTdtJp3FQBVhY7Pp8TNMHpvm2M
NSRw82ImnJob0Eq/krIvWlZzJbgbOmULGJD4FvL779EwUJepEUpk7OXZ4wsI
XxvbGKh+QdWYEORTV0/1nwPtJeDl5hvoAccWG6dXKTsygQiU06Sst8lHeh10
DldN7PpUSHu3NDdffQ0laBTdC3ToNmmU5WXk47ECqoDZCmUAGT6QKDgCaISj
LVfqd/scaKuFLrHu2zA+hi4Kblqt0OrrgTeVRLG4Onta7BN86EeY6xTnn7RR
leFYUamgM+E6Wrcoa/U4qzGr0FZyvNE7UOXlLuzNSdW0WPj5FzF92xOnie/d
Sj2wDs1+JG2/0U/SDVNV9NPPbaSyC0QWFauS1eUCIZ9i+kcOlzWOWSEg2xjZ
hpFXEzvzd8pwbT4DKJqzU0ech8x710Pk8S8S1LczjKAlOvgy1dXhpO4Th+zb
3cROy2mbKOZVknS49gjk+Il61/WdPPDMOHLOpaB6c3hDDvgzhzPwT8tXot8j
L7tvYgGXKOve5wE4+9eYHTdSTNs02mJBWijFV1/QztWwk0mEgoYHtHX53OwS
QvQ/Vqa3JGxWFLYelGXQPg9tx2HGn/SUVlDMBaDtZk0wB7PGUNRfJKFDOg0g
28z7krPA4Xl5Lucvc+OeFBK3gDL5ejA6eRaCb3FVuYOrBIV/L8E2ZGYY2gM+
X92wZg/R8H6yBkQlCOEZeEGWFW+NMH5XA42PgsBiLmOvzhKrpDR8H9wwIVkS
ZnQOwuejAqUoIS0x0kSlYd25YkoMTpZUixbQdkCzmaF9BjDVvVyTcKYPhdM0
pCZIGHS3zKPJ1GYtF5lEk2vZ2PcUJHbKvSjvBGloRB55ARCzvPGZd8h7FVIW
8PGPwd7XbduaLlUQEbBf7ujy6CRKlT0u8OmDUiupdIXfAiN8gcTVdj5jOc2H
WJZjDt4p6uRbJI7FxPYvq5aboLV4rxSTuDLPdx+o6PN4GYnM8L6MY0rMBeLG
xZSe8537dNMgRnoEpQvniYagWMIo5FOxAl9KANCzn22I9qnYPekExK/l8Ch9
+ush5/NT0LdDbp2sVqE50TOBv2sRsiJcAe+mNNe0nOo6MLWMpoxzq75K9zvF
OB2vhRB0QNyJxljN8wIVFNhHWEV+w3asWM5Y/WE2JKQ2BQt+hBPiHvjk6nZ6
PtUL4d0JtIYGz4yCtgs0URv5kjrsfeOxuFwiHfRrAWYwUIEFwmV1ZCuCK+DH
TduLAw73K7jeJvAf5UFvzwMmJ/NOBB0DeGf2rTwR35NWaL4Bs+l1cBNOpk7g
bbHkY/dF9zekLAIskKuCO4J6DQu+l0CoQrU5dPx1aF7nsKrkZHMY6C99N4ST
orJEAhXcCbqS9mXUGbMEeUeh+/LkEgCX8W8mUYkupF4Q3i0djvORZ6Vi2RZF
T5VbIrqriI9GUUD8Ev0HP70MTKIDOnDOZfQh9IExxDQqVnSbgfNaAqZGEId8
ujXutVMLkXVVJpq/BfjJyXKrEV/EXI/LbiPh3qYkbvn8Uh7766CP5lWVEOd5
wGsW2DUOU60aCfmZ1qDCdjDhzOve8UWIhpl8qD6mBDD3DVPMeB3b5IMDWos0
EP8ob0W1ft8poEX5DaiiaP7G3sCqLjXGMaqW7UW0De4zKQ5/0/AUZ6QpXiN9
QKp1Dl62w2FMgwHKK+x5dz2w/GQ4uUY3nFWLzLTzPFTl7bhXr7w6jsEBYp0m
hgdk3cgZFDRmGyNtme3enJ7eRwoR56o4daPDb2yirVVog3nzLbNB4X2bkcdW
rogbuOT/OkEY+J7IujEx6hm1qRDqKGATSYxS0AGFA73o/AxoNzSqp65YWrRw
QL4Ui2R6owY6IJ2EVP3LQcBwtMcFdqWFdOa6Wtfyk0wNWdFA48QkYaQjUypf
SnYs5pCWw0gUFV0862PhenCt5KBXe1BAPabPGja5QQl+7/SdY9NE26ok9Yjw
EsLcNhMuZgIK4Qs4LCAQTQYcx8j6qEwFJLwq0QFm3/JlRAZOVaWmvel6AAMi
OYe5PRr5HSLiaX47gioaVV2Ml2VHmp6ppJ8gPFx/dulUBQz6kiGOboIogFwH
9CMAjAc5wlpAL7S6jb8Bu9WGj4RnLFoZ53x3wcQH8iO/LU44vuDGAe0D06XD
0li0RbeOdCBXmqS1/r9xtRfsidrIpLySDC9b7MMH7QNsZ7eaqFUPVp58V18f
7LmxSNgs1sOr7WgnZ6G/KRIAPrWMN6kcMgjeohmcIckTezWn1FP9V3w1IC4f
dcYF34KhrTodJ0kFUEB4qN1/ZRwdZknpuRXHC23+6zHf82AHo9W3y13Tg2vc
dHOG635bQwU2fMP/lSZG0KnEnW70p6Ww8xjLiFC4CO1uH9AzGxHO3TlWqF+p
+zKbCqOspFaOx0jtMG7bPGHM4G7wJHLq6FSwRZ0BpASckYXr6pQYlkNy8bH5
kKArBUtzIWU6YSpYMk8c/p/phcLqiXmd5aeJFKLdzJDquCKxIX5oe2ouGvk5
oEK2lIttSsqr4IcsXANMhCWz9HYxh1OGCDB9mFi3GqfwzXP5gbPckLkF4ymJ
48k1xMCU/Jbx4eEZ5VPhwMM5OjSUQqLv8OnuAtAqa7HYPJzPG/EjF8iCd2mD
c2CVA6gbzjq4kkEFQ3ckSgvj3NCejr89ujrJFjJ/W/LXWQEsvL1gLQcN7/Ru
EsskqN6zX1+k/T9XME0sBsHMOstVbwmjiTUrqGxTIiBKKXyeCGFgaHX1L3nL
LYdeTxcBLyphamnnRROWrGD4GWRte1IAL97w8nPv0czUlGU3/kYmJsKjeStT
4rVbHBbj7fYoN04tVaGT5rDU7AWbq+O5CrEvSA0uldq16U222LfWHCd86Qbx
4LGUUJq0vN8WiCA5MB0l4QxQAfIzU5Fc1qCrrDyFxkQwqgeJXZjWs51p8UFX
ilNc8znte2gg+FztEqZbkY14edey1VvDlixL03Rx7NyWGkSMOFfHYd9DEif2
RGsIutl23J8y5D8WiTGlhgO2W01qmKHFxOpD6knLW1ua0kFW+lUP3Pflp0uw
Zpz7+PnZR51OcXUuMoD5DvGlsoxA6+3z4qZl6S4E/hBThwIB5juBFhnV1TLj
O1ByHxDtq3mfKKlJFY+7igSXal3wA5MVtcHn33tF2Ea9L2uBiQtTk0ktvQQn
Vwe2SUs1mh+ed/RyMgeUek99ZvTxfea3m7NmBMOgyDWLaVgUvn9T7EAZ5oxS
3gIGzqKZoKoZONflHhhYehBSGziXXepddPEFrYp9MONEG+a/xNrhc9tPdgM/
owRKVc4zl9Sdm+K7oRzETum0LVLkwrDQS2lvxCUvsQJslMJnT351D6TEpAZK
2fQfq7DUJDj6KvtkbJdcAIi+rfUx5fTHf4eE//ZJjvgourWR9eLp264iK3/4
xfysOSYSXYTeFd9Njm5T0eBJZGUXkj+7fHg9yr4FGPH991TnarRNS3jZIaR5
EfGIkERRTMQsgdT4seTNkFl1OPuLN6tQnNHjZDS2yi6PYpiABlaOhx2occzR
DF9y4yEbPFM2FBDqMzA+S03oQ65N0QJm88b3a+FlRJgn5JRuAj+Sdd8Z8guX
0DBSdKg7rcdDfmqRrikAJ6kOjNyt0gkzxB10NbFiCT4iM/iWmn05NwvBErPM
0wNjhb9jlwa6fDf6IU9qb49FhMrpUu+uil5eB9eu/Wp9mRL8MzMtmlZJq436
MfPRSxcbXdz4NRpEXJSp03ls2hqzQlMAtFyCBdvEQCoUmTMdjRUmezEZbUZm
XsM9eM7V7FogEKdO6rdBjOMTqb1Y+UYXRS9MrtpWjXlZl4nLwFPtY7reJbj0
yUNsPk+E2UoVLVoniHt4robWWcOSPGcrlBbxWZGE3zNXQLrSm3HgYdaaMYxC
sSsAI8a6gyiouAOz5bkK2YgUqR4Ma+fuVLdoGUbsNXyiHMbAjJ0f0GzKBYRj
7++8w20ScZM+Jv63uqGLo2Wzon92JDasbgK3BJT7JjZEuCw0XcXkg2jzMegz
RsRY8xwbZOu+CQj7dtn7PvhDE6bBdKHqs/456gqVa0tI6Hic23gCvzp2vXt2
vAVs7mFymw0facuDLd4KTBV9KBq3cMkIMxgGfdFk9620c1v+u3HBgRzjmjwW
zPUO4/HaRcY12MufdyFy7gNDmN7BDe6BjiZCG0VJgGneXlEg08NDyIWK/34G
YsGXLfGg7nbCsYR5PzWKIKUZ6/RwVkwFmA==

`pragma protect end_protected
