// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bYtT/zkZVwqyV82woHUdNAOIB6jauEMQrjSvNlra8sJ2+7WvlUHBln7loJQV
U0hcG2yh933axMpZz4AXcBq2n2RaaXU8tlAesuFiFOehwr/BLEPmXuRYdTtB
e9uI5xS9ga/ZA1DE8Il5xbDy2zmUyM4Grc8elSTPBMUvEXwWAXRbWccmA9VL
44oSkeRDWepGuoC1rAilZg+Z4FC2llgdA+a+pRzNrCNnuaORUe3xwf8cl3Dz
eCShWHPKaA7YR+igq5vz+20tx/pGXXp1M2HiM63z4Ie559G8jSGQalIwP+Ez
sCGDZfcBQ3ls442fs6TiltgaMQSH00RkcNe6v+766A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XxG4MhL8A03SGkuh7YtSkDu2BzL6GRblv7cq6sN1NuHff1khtV3nHS3hgt18
vhQAVrrpWQvQXGeeqBwvtnHHXi5OzpZJkJz79+cBd0KUxOw8bxe229go9Zkn
/vPpDt1DQT7C7tNGW3L8UuroqORAuArQ78tyWHF4Al6MoiETKNiVaCL9D7/+
HaT4hODWHjYhKmK2kX4+A4ManJBp6ThHHod3Ck72hDx5Wt9HCRmXZ5rAQ+Lu
9uNDRQeoRv58k/7QQZ+btgLSMOBCM+1zWDW2lEj2lXf5ukIJzbqodj6UfBVC
pGM3MmrGtk5mEoSxpAnc6l7uFyLBaMmQYBF1nw6Niw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k1QHBaRlkNv4P8vr1t68VYS/U2Y75QTFxz6eGLZPhBxKRYptF2ybUoXxAEuN
7cyU7drQhFMn0S3rJTvyHxt+HdgUfgw5bibg6rhoybfkOqoYMvhW/brjTdhn
19FyNp/NH5QxjsofnDyh6NfawO9we0wEnvR6I9go1mkToM/4RnJTdpkAVLc7
rzBocYMGWJw+VL35coSef/SX9G2+QhwjT2FbL/OAglN66sngSD5KJutXrlHx
vp6GpH5osjV994KfHPAO0jQlfocTiimV2owTTZKtEljfEDO1PDbyz8nq/luK
Sopa78jk8bl2vhdiR+ezMAIfwdVbKs3CDjwaF5e+Iw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EtpVZan04dgGF2VhGaBUkA7Q+jDruZBtA8WgLkBmVFScVjeX8hsz2D3A1Quz
Ra7xsGcckJL40JX0pGf6p/+JUpyyqKIaogZ/DJdFl6JlgpYpMbC380XBOXMn
EyiGwxGfKPJsp8iKvM91UwqHqN7g3Bc5ZEpD6TffDksmYQwxqgc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oESvRVXqATmgtlWLMAv5hL9TH7R8FdM02T0TrOWNFv5f13tqBsmAAdpbvQQU
Dfnk8/s5kpSUs8ZTKDllv3IMZ6WunDbEKDp66JfDRArPjsJ1n8KoA2qd17gP
aJuwHy42wNMvBNG9nBRkbXTMp2Fa62COq2pVB5YtqMZb/VJqftaj3Fh2Rfsb
DwXbdy95I9q/BAQ1u+y8qR/ATbbbGcHOURkKjfbfcGX6LQ5DmoMyPVrxH3sN
peH6FWG+lL4xUyi6VOSJiP5Ck5yXPNwtSGgh2aIoCZQ2GV3KXK6JmqjbI+dB
fqkBPxb/gM6i+dArHkKBCONkV3OYqIA05aJMSo7BPOf6u1QVj0KmOwl8L1rP
CZ/5xB7esNMj4PflATZN+2bwIiX4DuH0VZTa/Qg4vx8dgvvZtqMwFHrhMa1Y
IpTXBTlNjNgWDscP1Cu1itawWyGuEVl9+eLdPLKPhtVS8DiZY3zGuGkL8w2S
yrarFloLcqgxsgBfB9k7ZWHLedQydshT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rOpRMYakZ2Q92PQb+vWVqpMz9IVHIRphlqPIaoYQFnHborLRT6U6l/VewQqu
IXxzJL8P1RrKqIK5/TW1h5S4juBLUDLP/GcGhA9qtbz89zTOJeMUI5uC1D6g
9LhVJ4v6rvwaiSND3Yy7lXQiwEyNrkHJ4MZshIIenzH771UDtY8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rXJvsaGnyZDSLZLl/PIvDodmCMLDVkwH1EoY0abNv0+xLNLFTIUjJrc9oE80
sXkMNGgIlP/n+2P+rIyu1WUXJs9YsFupXxyEqfrklbrVrFEiiSQ9lZLij6Zn
3geRRVltAlUC5CVGwe+dKrfNBjQfuHYh9QRFVKVCEAKIHfWMAQQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16864)
`pragma protect data_block
lcNDRnOoRQID1R47xkeV2f3nU3MJO7UpPQKrGCj66e+JA+v9IUetHCK2Vylj
TDP8yfHb1PJLKB+WvtZ/QOi+MmQIu2rrNOmCDJtAXfgLpZtb1TgGkLsYeNDn
yC1SY5/5KqiiLA7P3TQGHE08G2jm/cDTASiLI0tqvhqP+Nl9ZHEeKvn6F8lN
rEI66sMC02CTktbfJg4g3P/4aYYaNTYb986+TXhO6h/2DLaPW6glswhCj+8Z
iOxMMge2otWafIZV5PDzY3vAZGMZQRUTqjDVcKuLhz+s0YXXw3qLhZM8+2IA
HHpacbPMDaYkoM91FTbouUkgstV6g/nOZ36k7PMEgilE7OOqTwGCsNzUV7bI
xfndWPgU3GKfQNbLevOifMQZ67vWUqk8/b3jrbbLnv2BaVBIsdwyeFx22ZqY
4Np22gf4UXCBoDx1tycIi8QTJa8FKV0yf5KdAiWNHA83Y45rDNeQ29cAJqUr
FREPuyRZ8sDZ96dL2WmfCYZMGtqMPTzQrzlTiPOzXEz03KZzLqRO8dddKEXh
m7N12JtTtCZvgwMzQ8yuPBD4OSY6eFB+f3G69TV+B7R6wJRkxfnTXd1P6PFM
yfmBTB5aMSS3C3hfC3MHureEPC48iQYv9NLlsHx3iaOMe8R+sT9JnHBZ7vRY
UtOXX2oupWo0u1w3dTWAZwX/dgiFFgncW9yGzW6dNVIhDM7zG7mY7Y5QtUA0
Tje1mt8edmCZzPwOuwC8DzBBHbe4a2Mvji7/krL1qE1XqFqqFN36wc9AY17Y
U7AUfu5U6pSJFP9CWvD2HwlFRluGV5ZHVoJc5wt0DCQz+6r5HHzPv1EPqFL0
Gvu2nV3NqGNlUfziBS672SjePlAL3fZIc1IE0QRf2Tv99SLCywZpiKZ3bIJW
shCA71vcuiDHWQLzr7pNbrCAtFY2+eb5162EBzhznfUqpIjqSuoiERd43RFv
E/rCheNK2vTbgC8IUYd/VJA9WaaOnC7Ohu+UEBSfTekJ/WJ/J/6OxqchGA3P
HYOuFvVcRvo9hpLbdDWxMDsSxtyYQQ+al6Hks+Z1/2tyeoXTR7CfIsW1E9YF
z6txkGO1iir3awvNkS79O9fpPaddFE/wQcUDISZDIEgHwDPdY/vt8zJUGZw8
Is3F5+UmN9ie0CdyPX+GmMRwPTe9T8xN6eTXpCn/ywUQQt3mdXn4f1w+YKE5
+XeNdLIIAFgbCKtD3tRafU6oU8zJ4kZaLiFx1n/X4VbTkct+gkRGGvhbn49m
0iSEBcBrnAOkV9sQ30y6tFhL6X1kc96Q1flRjwHxo5APzPKKjCy+a5TPIK44
5jfPKzWD5BjKVJzR9iOkEMm03nogrJ876vNVo32KS7HJEs8/TDBs80An+9I5
5cSP1yjBkR4nYumbSkhGGHwU/Lfx+VputWggOYvnWZJMYQG8+xTGxV74L+9Y
wNSaBA8AIzvlJu7PIY3+BQNB1yoicxRLRLPf2EWwgn283PpRNIH0h6bwdZ3k
A6MgIWjt7s1OUUPL+dIOBebTprfDnWKZrPi5jbQVhFoI9gbKZmup/5AdGaE4
J7KMZQVE0VJ/a9+rK1FsCspIDTjy17ZmYJpvWoqbvZOOq9OvI+rifIFRo/Ba
hQ219TD/Vma6n7MSE25uywagSg8RqlVAn6K3uej+Ps65+lmOgzHJSQpRXEJB
aRy9gXC5faoFJZUnZcsodpUPLxmbmkXhu8pSoW0e2ntCbxwen6OO6eK+FQmG
fesWrS8a3FH79CYAzK9YgW2gE+b6CZNNGdUC0f3+A2I527beJw0EhhXoYcpe
dBv/QfjPZGCwsfiAHfYnrGJ8o5SjZrFXRlz3mf3Lwf3seh+uYdCKzpj5YnZ/
WHS9fOOoIfUNgIMpvX0v93E6dO18IO2d1qQG/61KV7fwhEq6BiCck6hQapR1
o88LPZNdFaH78mM/mLf6mwwu812epu5HmCc+WlKRTk4qPG8kEh+NwoRY0WtP
EP3PVSM3laua+Lm0zmtBCbTm566FkfOT1x62zAfwBbtoPln9PaetXH4pjCjc
X2DzmXMeZSxkuPGkvM7XcPuz1CTCWjO2j5qv2FEGWe6BagOHvGAdyrLTyJjx
JWKSFv8bYhqSd8TCB28Zrj7zNSwv+16qRwjBZPs/ePCqeAos9Pip7VJieUK4
qV5JecVnwEUsX+k17/s8JiYaLI860iGcXgk+2CSzvQ5dQxKXZtQf6MnduJ7J
qo/RcMkxVtaLTIdrH/Fg8CmoeIUOM/4iUZmSSLZC95cDPyiDKFvCtvwf0r3B
WQgO09btVqoVIz82kc59C19M7dnf91jd02/jXfUXwAY4rWZdKfDIw3+bYP0s
XlBjiPEFeBUe4eMc9mA+577V3c8I2t4QQdZNAKC5eG7X+okT/gWg4aogYQNZ
uvCNqgYt1JFyQRHvpfJWtMVPngku2jVUCSdcGyp3Q+W5+b4xZBrIK9eMoHKk
kf7pSQsPH4TpTZz4lkPsG0SMbaqAQHa2BDNd5ndK1S/gv+IPxfjz2uC+qR7T
Z7Lkv6tkPhYXL5ii5I5VB62TAnlEMKeV+DdKTEJnNS2csSFcUGf2/qa+nVuq
ENyZqnHQUllskoS3oSADBMoCHu94Cvw78yss58JG95woFcIa0kCHGWl3J5DD
0AqpmCFFZTU2DFpPvuDpJLPeXcWbx8+O6jNOQFcEknC3OZTa864MoPXDa5o3
NbHgq5qYF7dwVbvK64u3t0uR/NiKz17+VyJnNxMK8SnJZ23oeBGxR1hgCVJV
xe6nKpfka5Te6nNthJq+txmbRi9MRNl1iKs11J/veeLhX625uUyw7tG07RS+
5bwuziSbIo7j/7aKq2UeeetfDXwX73+4GhvhoPIi3/JLOnYIbpf6pHWfd5oE
5YWfdYpdG1agF4Ai3pt8SIQmTtHuQSZJbSZl1DwODij4vy7e3xzT7nW8ySvm
taASWe2e0f74VeLA4WXLIFMDtW2o/c4CH0z7PKJB+r7MqSIMw557jKk9yfmJ
1440q/qOKtW4rDI13JFiRCYvgaVmUUzaXC+odClGQc39K89c3r89jh/yeKB+
0Aadn/a3DehF/RK1gnqrK1TfaP9sbZ5NWMWLJCeKpzv5mi8yCvqPO5MI1Yf3
6MHCndbwHcWbwReFihEHcT0jIBHpdKDZ74FwaE+ISVQKPUQUVSyI5d152CNI
maphlJygahl+J4FodZGoW/5FYaKkJ4uhfJo6kMX52M/tVHlZ+95asf7jtrjr
g+KyOmsfPUaFw6FzC9xsV5KGXN2Tuz6BHmj/IygcgBagtR017QYJrHZ6b5lM
mwU+vEHPHfRfP8TfhOnHKyKC3Vi3fWfR1gsQ3Tm/pYWWx7hyS9Jv4eznEEj/
P4fhz3QkBowRKHKy5PTHkvpnI/cWstS2r7vtE5FYw8TaaSIud/DSo2tQNuoT
zY87AGi7x+6NsWMjX8GZZDhRhrz996/dwDDKxJGodYPpusXbMQ6VjWvuoV99
9PnZ1VMXI9jKTFyCP8y+bbs3Zn0Rxcm/2EEqOW0cOnwvh4ervpE3ysHe0/KV
zvxDPkq6ppLtqV9iV1ZCCm/0ZKWC+lCE2OPHEsPtRUb7w/MW90arznT7Q2VE
IToY4DCbXmJAPFOFGvXK30AbEuNQOM8YFTxJtnXlscIPT0e9/8TM67vbPxvW
1HfW0LHRfVO4gGoViJhzS+oRo3OaRKltIfM17dtAP2WHTjLAyLF9AtmWzWFu
w573ZaOxJl39MyMKra7MidO5LXZoTg0Z3Hm5S3TBAOWw3ZXqs1nd+lRMb5pG
yybU0rVDD4hsl0LgTueOSsvlMX6mDlG7AgagV54hoxw6MO9G6I4YZ+Sn/jnb
HnJfrzNUM6RXGvp0n8L5bAuD7q87ATAtYKcAHDeZLBDQ78W5Yo4rEkZJldbe
w33V16C5bMJzdIJJkKPPlU9p6ZhptI85hIhPd+UfQiwhSHQNoJOHxzQl3u1u
/jojvwfuwCtt1nHuPCvidXevDxq5/gh48Ckfmmnl5wcrGu1SYNaXaE+4ZrHI
szmE7rdRhJOmyw10+XMqv1MzTOj0w+8KtPTbOcnN60Aw05iyoz5xKvR/jnzo
msC0W8uBAmhOD5XQF2Nn116xSvBtuNr6PnpmuLc6rOa4huDVp1vNw7SpHgAY
Hm+WpoY+HLmtyyn4QYr180KFLIfA0LGAccQuYozvFPVkAWUba+oqm3VbDUst
qMtBMmf4KUnfIrDw6ezZNuD/4chhgWRmDeoDiN/1N4Y5E8yl9TRvF0oYGuMC
QY1N6hit3NsSoFITnKC7bIubUD6NUiytPa2ffmPVzv+mN4BwMc6/Bl5REUyo
loLZaKwVwvcAFyogHxVgf/UeW6c+67Gq6/tZWXwV/C6uFqFv/zsYqMxgv7Fx
OuGMtlmioSd02Fgiz8Y2fuEWwLN5/C7CikezbHu7Yy9nB7ooxj0GxmpP83Ep
rUkFNsBNYvSYmSPYPBNUnNnvigdGBcb+wbrsuJ5rYlFNk3CTjHmAoBUmVQ8H
gi0lSR3wCv6AVarSo1shk9FXevBYuT3vcB1Zo8TeTi10b69T4NhRri8HTB3r
EuWsxCXyGu94kK4FXrYmomvYgxm9IpYJgMHSpmYCh+CxkaVJBO9zR/L3vOfp
Wh4Btdmou0cUsOuQTGwZRYAY0F6Nm7UF7qCN3Br1THCfs73GorkdFeTyXQ8+
Dk1gHvyRJRPkXkE0/4qaMo4NDLfCYuppUKgq60vsTQEzJhenN5sh9XnsxGka
RQwz2pTKH3++OTbBw0E+QUF7B7LutYwIg3iJ4j2NwHjGvOqzmmZkBm+YLT/z
dtgw7diaL6+LIsYlUKw5ai+ezH7j4yOFt+Rn+sqjqACkATUcYKx7R5o507+T
nhZPryIpMygOAxVBANKLM2Hf+wh+RLxBflKtz6vqpTqvPt3YfibBth0AqcIi
pdKjzZkii9HrIxx27UasXsCXQpWJ+FxtTH5+u3dAUPPxdsoA1J4eGYNc5y2o
vv7ZgPEKqiktlQLmdzmxNlCjeRnSYvnUp9H3Rp6khgYt/WfaW15y4G3EFL+0
lNnFL2+VIWtg2xUo8N013potaASRb/9y31BTUHUi3DG1gqXdUcGo31cjuEVA
7xRbIR4rC5illmjVY8KcKXETBd0fPLeo+OazMQh4qON+KZYpSpc3YnMDADIF
xS3NHiWli5pAXPhkO7uDrxcLBzbE3V0hXULvBrQgvb1E2l3cwctWkIYGGA8L
fG9r2PsBdEZLpdzwSllg8M8Tikb2bdNdtLJOOsII/UP07o3vu20G/x1c8ovy
bRCniHtklqZAGNdexpsDeM0BmU/aZm5ZJyolppTxvw5RSpg/RZF0N0pzZDI0
oDAWEZfeTmEZ2sQphy+PVm405CrfqHWwwQhRaCOq2sJTBrhwQV6p8HdLaFRH
KT6orfRT3487GLgj1GxOfEjs5VEC12qY2vE0hTMCsyyqEDuurlzD+Er6kGwQ
0h1oJ4KFz0fL9Xf+hdiSfPuzdqA7qzLErNEzQNAoCaMX3zlqzIhJJMRQkak3
/6jJejNKeqcV6D/XrZiRr82S03UHeD/dVl/PcWO6LuSO1rzOi2eSUhJ+6ey8
XSiJT6Zjp58e22qEDrJyCZ3h5WVDAl2uL4RBxwd+8g6GRtuRrd2cVw+F+a1V
XCQ+zp52DswF8+nOUjBf9nLftq7RdLSgdRBnsgVD860he8C8pn7VS2LDiWGb
i+ROFhTQ1bd2e9AE0F1L+jVdlk66Jkn8K0Q2dQY6owc9wqpkAbg2Gh2BLOwV
sXEGNmF7yFwWEPa5djPzoNCpuW+ZNcbxtbQoJGRZF9acoavycKxmYWqkCgd2
e3otuLB0f8apiBKD8fo6vOvX0VWhP3Z7A5Jv6XAlekwmiRiZES5NZ+1idIIE
gMBODsMDvs5Hin1OuOmITdWslJSlYi86dFYFboB+DCeLsoWTCu/rTjx8eoV0
5UDENP5fmGlVGz0vu0cz8M59mKqC/eFUU3UHu2C8a4nrZaulcW+RPp1oT3Uu
nsvresORlscHf9Sfb6f/dpZwdJajhbSDxoWNRwB8g2Oph40+XXaYDhQZtYrA
IN9cUING73Itl7AFGRztlt26tybPFh+mlxicVyzEjj7W0r0oc/fLcElMFAn8
dPXc7O8trtTy1/Y5rxx78uVGY3eiMpDitHWsnU+ZZfb1hyUykf6584OwjMBl
ATFd59m3GGUOqHNE27RLSbYe1wZ92EoP3KX1x0nSYxNaQ/SNhflovfbemMkR
Ux9xbpI46pgNJCWQWg9jxhFSwzAopGnYV6gXAdzFWSylE0PLc6aOiSGzV2WL
LTucz7Agfk1Mva6/61eOZeqoqjJ1ZKJXmO/pVhc7ncBVqKtkZjHq7S+a78aK
UzxZ0Wg2I6QNVbAcQaGofc+fSBg7gmfi22J7plUyC0/ZQsBTGplJF3FKPQOU
DlKk4kzQPCCoiUY3+q9B39zq8kd4aHhzJbgv206h1L9/DIWfTpKpe/8E4OIk
NDponFo6Zruq5ua+2/pVnPXelYgeA3gnnhqq6qirzpmxb5P/ELXHB0hkHhBL
QUK3W65aLch5l4gA+vxbhHDnowt/gxBvcRVR4N32bOLOA+0WMPfxdJYn/crE
/ZXE848stAtAy47cQKZrBT/OZz1CdGrezyOuK9iVLhDE0IdBAfAcDJxnb3u+
4MIJqSudFvpmy3rHcruXEpb7S7wsLVI91ew9l4IX951drHdmjbwDO4L3pk4J
pMWFn76OXNGuJDDpaddqAC8QP4APg0BN+GmmOFmG5FprxEKfiid0sq37J9r0
aXguC4QsZGkHprpuikxKLhKQ/+Q1p4rzsLJFYZgCocRj7KP7PWc9mLWDvecF
SUAvZ2HEj18GP77ZFhbzrKjnMYbQ/ydjK9H1sUyEQjGT7qZaUgBDIP0p7aSA
EiPggo82e96t29Mb9lH45p+cEQ+YmrAKtlOU2wa/UcWfdq0lNGnKAdGmCDHp
DTVszARC7LMj1A4yUu/1/vMz0QnfO7KmY9icWgtFglZuji3MfuV7jEGAeeDi
xup7OgkwXR+hbu67x88b9f5gLRHzs02qfGzVDWNwy8mNqMbTflIuzfCQ8ZgA
X0b+CfIhpRxMGEvEfwTSHLe1r1ScQhBoELh7skgnPmc67EbjgTiQPiN15dpw
6+Hcogs0aDcYQ5IFKdKAhhOpLTb/mBh8ak+hhRxAwj0t7L5rrOz1TmpTdzLJ
6dCVAomPO4HoMy0dNYzAabp2Sl7mksINldjScEZSVVYbW11hsKiM/HqPpQIq
N9yUyphombGeaD68Xrcd3nhxJXdUrpMXzljL4XYp9ICHbEXFkn1x4kxZEOnH
V10wN6oZaoLRfAbSi/47shjGddDoqe0+tfdQRinyoIC+SvvYTNDxlFnvrNdp
HOf+oX/hdjWVzVzZjQO5Nw8XHt6u5TcWeUCEYuW86fHLsxu7eoxaWwL0nmPs
w6mdoZAe6nYC2m/lDdi+IIVdlee6iGCTgON03UjPZb7/mhObx1uMtFhq0cBi
czTS8OBiJIg7SIKg0RzTQDcjGubISGcyIYuNacMr76GAG5bw7drLjDU9MgKG
qjfnzalHjKaUZdeIPzl2xyepechKE8kmeAsKTVFmv66X73O0msKKq8R0iLpI
xsxMcRw1lXK7ahEDYdrl4glyBXTD0z3rJNdL0daYFdlo7INGHbvRPVKxitlR
gnQllA4tPHHm1Olma+lgFdkpYAsNFg381IEgjni/S1eA7MseQZSMKlErMaN2
QYJOqIceUzekvXz2whY3+KIES4Kj+5J9YuLGFjc9hpBa7hAZwyL6TpuR16br
yxbbUk1pfaJzadhfF2pGyVMUcOYJihKaR16yQDNlRWvJwoBchCACnsu230wa
hWeOd2reyYa1ybm9e3MzNfYvN4fuwZsUzR7P1m4roAmjCcDTkIs51TETa2DB
hcpMADmXdIBOEaREH9BGUNKPojt78vqyhO/XXJndrMrwiaTl3xjPAO1Zfvbc
labWTYZtgxFoO54B/MIkluSH4/o6NbUh0oIXI8NMOvwdP8stkaNKkvIAFzPH
keqz2zHLIgDK8naGQlnja/Hu4nxyKLmXKCpFKnQhbyUm4IRuNIyeeUVPIXZ8
4iUqLfyt0YcMvZJV8zZ3JHlLZDw9eO/vZUBPW2uhSemflPdXkjhH5MTvsY+o
KujtoeOq3ZhOKoxK8N4XRx5iosp9ydfyNBXZ2y2rQwNos+KIscw8B5VwnsN4
ZrGrIhtpFzuhahEZhVF2gKCyo+fqbxuZR6L/4BFTAkUfw0uLjeQ4CRtGSTIe
GS/JusE7P1AV0bum5Oti0EUHvigtfJbtS8rJlhXVMmlboJ9Tg0/WwIcw+LjM
IGDxLXUnoqGgTZ/zIU0d9g1LFdCFKZtXUI4n/AvM+3EdL5v+MoV3fEaCF8sM
qopaRmjSLvgk4iJsUiO+3PgrCfXWsT1hPBhs2r6SS/Lwq9YQxstZ87zQcdc7
6bmXtrgp7xSlROCf/6Jem9OqnpGSifpw+Pn8H3g/89oXk7MVIWn6jr2n2NSM
WAfAj+Nqv3BQ3J5DW69UTHXJ9iVUovXK2CWTCR71IAWS+8yO6aFSoa4ySYis
2eiILKzsimeMvSHjIhTvKLjQ+lummqHpjnmYqvOYgcCaSUMKC7g4ceio9/Xl
v7MRMSpV3O1lIVvWDns6HDBYm0gN1jew7FnwvYXCrv8sfwFDIs+qi8FSC5hG
+cShiWNjRLY5CNvMzNwGviby9Zk4D32i/Ftnd+01sooFyEJUP2ZMs76Atz0B
e4tZSXKLR5yCzgOASUW7L9OQt8DxhzT0+gzhTWyGeNCMIwBtXeuGz6lu69HY
+fMobDPCp4PQmtQWvCqd90Ukgw1/5bXhwxgwbdON7pTUPJdcq9wEVq8FtvmP
+Nb8WnPpxug/Fi1Z6hHG6nnnkn/avEUrNJTb6GX7HE52Cf8jtk/yEHn87FLI
453ML2aXjx+XRe80VknPHnyWZtlD3VisCJdS1tPbo3VXQ8hmxvZS0bjgHTfi
tNKm5PgWGLPEPdgjoYcyLgeP/sN/8+unCR1zv+vInBYJNo1bW3yJaDVsdgHs
+G+7ihuNvxN98TD1ZU/VInb8uvy2RAePWm1tXLTBiQRx1oHVhSoZStSGCWXK
hmOHKMkmS6ECBqpbo8a9S8/4NC3Tia+LJMwK3QkCkGSh5/oQUUbJ6/lbBnlK
lT+QVleuh+pjWBKeHKRTWeq3HCFCVEhS/GQGqNiRtGyAlDyUFq4MV5w5OcyZ
NLI11i6f1tx/+QCLQP5h2iBPxoc2fnGL8nFfgwpMuZ5bLIE36EEWzMiZ1h7r
FoL+Hnx05wTcmlXh6ct/wzkAF0cuOy3R2GpGsKAW6lb9iuPZ6mOawtewMObB
gSTvhVHn/2s8FNXqbehwG9xLdsG2xtinVSIDW370glpsFhVGL4NV5LZkTwxV
HtWsKVP3DafvyWcaJf780pzQE5Wr5l69ge4iyY31u1iBklteApr/zP961q5C
UTyFaRoFZhzshpuGB4JOykt0I9Bm3FFuuHQcvrKbreEZPQlR7/L1HsgdNHkN
SAukv1LPX/CqCqtTU20r8DOd+e7byZFkRn5bg/AbBjS/WHlgqMFj9LjUg3wr
IuhItFVkJi1tgRN2+gVTYuxkeiPlvc+5PjrAXq/RFJpp2R0OoppYiLBieDrz
zvd/L00XWsF9aI2fjyIZfL9F/Mf+CB1IHQql17kT5pjoqxbhUgU2Y3y4+Wvi
6l4uHCU7BXF31BZDGcLWdSsbKheVhJagISPBxy3q1AytDWHgpxbgT+aSIXmA
c+2RpMo352YfEUPpgJbaCegfC9HvEGCyrQ3D6xgH+8cNh+2WSLpqq/MQN6g6
bQd/AschcQaMJg2MwnCsOqkoShpMYQkLHgbOz9ZuOrmXi26Jtfp96rT78VJX
upEH+HBXS1BUrJxr5rxu41s/zyWlJELqLTBFK5QcOWqU5Yr+YakdtJGiSDg5
T6idcUkt6/z9zvCgr4V8iSTXvXPp3lVMnR4ioHgKKXl+grtQ5bBeNIV0OrkP
xrRG7tvcKtnJ54nEgqXKzdQwwrYYkqHLwW2l+kodjvWaHxU0580chiKbcITm
D6/j532omk3Ubsjiw5UnqgvMoCkM/2L0QD37FNA6Av+FFhMWy+nKHWgCi+Rh
SUA4cgWO4gWN+QCqMjsoOexRaKhu/7OiQJehvqNtp7r4lTIzsSKpJbJ2/ODj
WemQRwpV0PwMEulI0QYHTkkWvchg+QzCqQM9Q1aNv0VdmSeB9lvHuJiQZ2qv
XcKD8P+ZmH74ZgYA8YPSS5RTyc/2YJKIPTsgqrSEC3F+gTKF5L/5W3fPTVS9
WDeeux9ZF+DePvt8lC/tGqOQiiJLIVN9pne0KETLb1HCZVp4iWnNo3o7/mJ1
RVtfUO2ewiNcVjv6Q9zZgFOIeqY6NXOReJod4B9UguZfGygG4ntVIOsvPFfj
9bAsARNC/AEcmQUs2wfSmnaaxYkSGx104sdmYcyTsqcZdbqo+IQDPHvzGnfp
DE+87Zo1s5pfvpB49EzEgWGSqYo+XWO7Xd5tTJY2yA0jHx4bGVAb99y1guBi
p9GNgUu2sQNgyBHROapQI/7wOHTUmH2VRxAL4jZmmrmccKavCsMyggpX3ei/
jahRts/mH4vap+JCHRAPYYIK7AwvY9xrnrRo2i+t1vyPUVaR4bDgaQK7cP4F
h03Yd76hiqiZ6sRHbnsmVb6lgQCPb3uaSjWr9x+UM05NzKDlJzqfEjrnwpdY
tWxXJxNvAbZZ7DvlvCxXHcx4iXIJiL4Zq+qFEkKZbhk98vthcTdyVSPLz5fu
jP64+bc6zUdLAegu4EwORJ6tuoYVxziQDku+Axif03gBYtgfp+gFDolZdQj3
FjexKf04keYosm9dbx3he2bD/ifIBmTaU5JV6ZFvs5hwvwFGaPeUvQrXe/2q
88nHvpC005fY6djQGwA4t+dDtiZbz4OB6mDGPY59C8NQbN+28BGY8BcIClLV
Lu6LZDP/Z1h2gdt8sQGiIqyv8fUv4TOIVLayzM7lVv8JGMhUvk2ozKu2DBIb
silgecjiAe/sURPKIFZAEys0v6aQhIApbkj9z8eLoT8CrezXbERCHHVxzApD
S2AYVzCrEwaozAHl9+1khcDwc742a85mhNJbtmiGmvKgxNP8fzrAPMzJ64Aa
1q/6Wp5rfUKx0y8aGvcOGmBrGpVEE5ir8s5XFrIreQokSkDnqaqFKZkM65Bl
eFMW8V7niDPTdclJdGpdftXjaqto3FLTCCnZWi4PXRWjOOnZe6buBsea0k7Y
03464YMDiNq8SJ7l/hLLM4vg4DdWY2WPkBcCKRpG7nyyFl1qHHMedfRkTfdM
BVa4Wyr5ed6dXh2saS46gBxyJoKCEAL12uIAB4hTeYjRXdYWa9zXeCILVDT2
JDmzc2EHI9tu4Fk4h2EXp3Xgl5XJvh1ZG4a2rrsEQTZcCADsI0V2pwRP1bZc
Ha0nfseCBqmE8LDKlsBkwDkSP9yRl0PDign5fmv8MxAH644j+otNyLBRIEQz
wMRo6RWBol5/Ee/5VEg3EOJJAUTL5OY02NN9P4gA6oPjXu8ljD4OGIbGrpZk
62FXorvFd7sUc34FZpNvcL6nQp3IcdUlpFbqMarZ6BdCOqyLAhqY1QIb00Je
peN63JohGASCbi6uqVS6FHEON7rFuL2qgxQoS2TKRRxccf+J+f1NJhG482/7
poGbCdlWrH3EJWEZzzWKTOb0spPgmZuYXaqTLmBb88202VMJ0FsB+sfrEPCG
IKtESKYT0UKqa5Z7c1yuyr/EeNIy2guJLzmttaiOKTsKlI5IQMPzlkeI3Hkz
jVURB8WRaijod3Kuc0tAlipfa3munO0Oe2L0KDi093/Swl+Fc0lwNXUk/J+v
JLCaKHgEN+cUPBIdm4T7sVxqJF0NMbcPtYG44wmkQ0xj0149dUOThpppr4Kz
faG5UZwyaI1GHTTrOzS3UDRcAqjZp7Pnjoco7m+eGZZMB1kiQj1PuHW4LhlA
3yVEbIIO0Hn0HNd0DHYkMVPsS7UolR8zZclT9pa3zo4tEbw23cGNsjq3jlY/
Y6Ix0tV8np6o5mUi2k45KuHgAcOK0uh5VJZ/Dr1wKT3ZK+mYR+EYRmb0VJ+Y
rgRTA0X+XrGz3+rOOZQlVHbaHjZMf4Cjp2JP1zVgE+BqQRLPmh2aQRxscJfd
jNVwbeX6MDoL8jAJQPhJAiNc5ME0lzjnR5R4KMruN03nx9K8XHb3CCeA6F81
gTs0BKV6/mlSs/IIrdKe1Tyf0pyotOl9BhLp9WlFNPqm4I7o2IpyXwotNMWQ
wbl34zBHE0Rfp5bKBHBB/x4CRjAkKio09iRsn5Z0Z7iP9J+aZ9sP5Q1w3nVM
WvU7tDhitGrs6jbBabQK14GqwGXM5PNP8/wnz5yszr9UZHXWpbOwg8YGXndl
BdV+xwbGjSmF9CTeqnwXiuEY3T3uIcW35fjq9VzvDYgmQTJ1+GdYFUZ36RwW
9yJp9fVPd9tpSg9mS9KHVdCLJ5q7WVFJimXehdtgtBJkYCgEUpspvfNSz0FU
1fAybFgG5KaLAy9ZAYz3BH8MKzoOpnZJCLpr0ktR7K7Nu7LQYbNoprRgD4UB
pUXBwwnHZ/Vc4I/bDLd8FvED0ncXiv4PgJRPeMft5rUZwVimVOcUlbCsMPa7
vTEfnu82FpcyV8CljfWHDeNDfniaI+rWz/GEwEw7IIgQQQcNwGgnlX/pptgB
iVeEZPHDiJmNrpBcZui/mqbIHQl3Xa4VBN1BPlqttQZuifJMgv/7VKjwjZgi
6DoRHyu//8ZJXSEP4FIqFcE5NNEg3a8mWalf6hZ8yhDwFuV35OpstRtViX3F
u4tqPWN22LwqcELo0tsKrB4FAWfm0ZvYExyMG4gkNuv3vDffx4Krc9CrTsIn
5SurWf9AV/U+We8PE37YSwSsNMFrJOJbhPYvnOkoNk4+2EhS5kJbydReaYQI
BDRBS1ipeiFMQiLM0DupDa+R2KQJgmkacErrm/4k8ggUke0/6dNKjQrKuce8
uZcmD/s/tgAqINadlA57QC4/z9Wf+Ei9NCQ0YRU3hh/gEoBTFBHe65ERHXt+
5JMlUFlNQl1XIf1C754HVFTCldoceY+r7cyfsox52rsps6FUGvdzf4M5ryzh
xdHML/rqT+A27dpfj8FlUazwBeO/KplCLseajmFJJWHKcvdWE+70biCVFQs4
jHLgie7EE9Rli89ZEiNXUILnspgQ+1g8fZ89qRf441FSotKLjglAJzaCYSRS
/Z/u0vHNumLdIGtXQFGvL4ktqhhViMxbEy4uC5swYEOE5YhGgU9Gx+HJmLrw
9JUiFCSLCcHINvunl+PcsrHet/mJGjxijwrKH72NSlcrleSOeerrD8XPadcT
9qC9vMh6jA/Yx/ujYz/THieU3bIUYYz0c74TjS0hfPMTPlCXkrx8XOJ9ga8/
RJ90ez4BsPi3Ivog5V4U2mRnW2ZzjYu0AckAhIiVxbdd6V2fjWscmOjm8Umm
3pyZr+Fzmdr5g2UysJkDSYlJ4BdY3INGE/p7bm1xfkzXll7XMK/gJe8rs+Ge
WYmT/OemzVsWbURmEx/5n9OUcNISzV2WuVp44therFNvQZrpx238udvE6GNJ
RhDNgbVQtwMnRpjYcLvdFBjySCX5bFrDqLm1ecl+uA/izAgaf0lnTyIed8y4
eA/8K8Pumt2AV4Xvv5Q0tCs8FNiG6Lv+HufCq13LA37PaRTbdfeZDesIlgT4
vL1dX9/65oy2ZewiY0Pr6uOinbcHyvccSqEPsYHJL5Ytx/h/qLp3acOc/VTD
yeqYguqBmlBC5YnvSgILe2UoOtce5g/jjaYcqj/nNU1cZcxC6SqRaN2qwpzw
E97eKYJc26dK6tX26bWNkeT3nwxhE+/7rZ1u24NZm98iDovvunZAxXGIhMIo
4hi+mKo1vPcJYjDZ1bNwieZ1bHCpnCCHFyDPlqiH6jaOScwMDAKBclbjxsHh
nwN12n78BjK80RIMidX7xMhySr38Edbn0cg58NH7oknBLQJs8Mp1xw6hgQ5h
WqolkdDSQtlQnwgve0UCqjBYrs62Yoq6Iuv76JmVhWKjnw2bfuqppRl8fCo4
k18XLZY3P+wVlDtMhpj84ECe7YphbAZvrQVsp4vglk+ifnsfjfs9FyyWB+F5
rLCzCbcLZaoyCR+IvES09BocEMoF50S9N8Dhc1WclQNX5OicDq8MfE9h/yCv
W4C6DwBhWTN8W1zLpcSldJWDb5+GPNsMdxM2qbz8Qf4p62j6U9fDOmD4k/9j
fRzhaaZ5jc+yIPYtA59ZtY9QUhkIux+QFohHSoJ63WGnKPMkkj5f0dkfBDwg
5Qv/C/mz1qQJKE0peiJ1DusTYxM7Xn+kzHpaB2X+akxmoJ+C8mvcArpGCB1g
guIHLjjKq5eCOzK7m9pKPFHab3Q+peGJ35aGbEN5SytELW1/iA6ea7HZSdLv
9neliyr0Yqj7ll7A+MJJwds9GsuzTlOBUyFnRNJhUhJ3UAYAJCoA+CZCdE9I
iyiYw5O5NXfVCUNXD4ylhPApKP51hodcaAMUHqmIETKiHe58WVz/iC9gAlN9
3Eok+jJZSG+rLvFyL4/ZcqgMW5ytSpCFqaIiQhHtAAqlIRLrhGhPBcmxAv7Y
QN8cW/10cdQc+7rBNfwwTV9cgFRxIM2oegyPc6BqV5b5T+tHNIyhZ9CiR1jP
ox3gfW5rC1LEqH2TYAT8Qb4XbbN7yyZEuLYtNlPuwWXDjnCzgL43NQeP6yZ8
WnVDgu878Hk9TqRPGgTAIEkMLmeb90aOBLRWeu1ODqRWBWG1KJYI3fiRClst
m/iFdiQDtbFFGao8313aq6oITWEZ4gZ1fvfXc9t9AOgymUytUp4a9NA6d1mn
w6nsLVOYbrrDljSYfOTZiEjtdezhVVqvRldmNIeMzYR824KZeSS67VMJOLEe
z7Pc/WSAd43/4+By2HTaKdbSqCA48yXw//MxQ8qxFf/Ku76GVLYa6kWTcCBK
r1QLxoAmiJXiSVL1AJaFBgIVfFo7KJ7Z7mEKQ63OcYOivx2lz+cCoDxQx/uV
6B4CHxbi+R97ea4oK5Se49EiywlUtkhAsgPRIM0ZgjeKuP5u59dizX6QNYrX
W8vDIPxC9uP65fiGO5JuWYchTBYttPMC6WE41QeLmPRJmFD34+uNetay7GDc
Y4aCL7pWx+74phFWZZDi0//w8iTwY+tD9Eb+a2PtxoUSoSFhGpGm6MV5RQg5
LziTviaSALZXOa9Am7y1YImm4fmf1XGYDZ9u+fDXfF/1tNTUDUYLDjU+8vV4
1G2uEZKGiSuTYjC9tBynO9zm2SEA0a+7YVQl0kov3uqDs3ffG5I2NcHRsEsW
RW7RyxvC31OvOfutPhjSOrh/BEOxKMR4MpyP1g/80pg+4tCNZSDtJm6S8wo7
BRY1eRsAI0GtnXflk2YFMz88JvBH7tCyPaf7wg/uRfeIt2Um8ZXQY5+XJyvM
nRMj2SedLj31oxIZdKgIhNQ3zt2IJElgQhC5ifN4fgovi1fvZaq87DcNmeBr
6gFcQIGjR+Y3HAz56fcUU7BoaAeb9WURl71/WdxabRziLuRHDrONuYB10ARO
EzdPKR0iTGJNccH+2+m7nl33oRKEpMqr7wYtPIMZhRvQRdgMLOHCmnfX9PBW
9QV1ow4nSx0e/Pqx7DG+EkEgafPVbTN2VYl0ACXHGeAL9+LzA23W14INmIYi
QKD6cxZTa/VlOG8/hlCmx8Uhlnyhl6mXkuLUotWbB/rjbdOgB9nrMjGZAZ8U
z9xRaFSKC0RsQNCKL78GebejvS3/QPPsp3QOGbYn1LB9ksdNlz5bx0jyUHiH
UM8ykzoOHVBrhG87mAW6dy8nb9bbXisCiPOViUQJuIIrBnuwa5orsbQzQkfW
cWpcRuPxJ/0nc/lMfaByPlYw9OG54Mn9FNSsTdFMDJMuPg72E1YR2V560emh
0RH46Tq/POqStOc+rAG4L23M+35gR23803La1CSP37DCDvYYldbNG+Ag2v/q
6aiPyl4NBUS2t2fei1Z8xNGc4P+PjVz3QS5/zvtHHqkMd10D3ueECnK1p3mG
PIeiZBC/DjiXzarZosHk4+3eMRNd5DtaBjNqKAQcJifCrOPk0a6Nl/+8kYk4
xR/AMCbjTu/Odwv80Vr+0iOtiq/rXGfdGEPf8v7LL7dpgalR6VAFS4YmUxCZ
AtgdG6gHtNtQSInZ2GiVFBOVo8Im1mT5+i4aE8ycpHVKDZXlgRQ0cbH56Vxi
16o0GupGz1KvAAccwlrB/pP9aAdkaKEKzO5PCU1IJeLBFssHQ4vUojL/oAqa
jIeGWpDp1UFBdS3UMWb52m3TmoKw873wPib3qb1cl89A3wqAajZ5hVMDKuNN
W62J50nEp98FjTiLoz4BeN+TcDasNtVRAEfmWjl0tuDq8u2o3fokF7PMEI1m
wyaSVJpS8f/f6DuAT5Hr8pD7T/E7xVT0p9EQj3g/Yx54VAms2Lucojus4xS3
csug0e5aiYwKO/qvIiAM3X8YVjddH/9df1kQuqoAPWuXA+Bma1/KtJx5mNhO
FvEIr4T/Kd8sdu3dmNjsiL0zf25K0TuD8FZOoAj4pjvp0a2T5lLfQGOe/wMr
K0I6UTgIJoAvXOAQ6rJ1bpoOIEdFZtXofgUXrgxfTFCOZX9ctLUQzNgwv38f
mJMK1bxbTrR0RZ/oOjelATSuhF1X0PsXGJLHrZPbm/bm5zXgaNj6E3AQanLn
caVgGczV4P4i4he56K+UU3j2+Ti//BVaXrtjfky6AcB2VnZlz5Y5hPiWXUT3
KC2TDd907XjDE+WdgrFaV593OQgfWC8j7OYbQoPQEtfEfCHuTQi74Hoigqqj
W2RoWZ6SJmTN3PrAK/5p6ujL4L3hRAlExaWACTwJQHIDyQhlRHK2RIJfPBkf
uHBYdv+ftQHd0XBSRS8pr/2/BwI15nQrlxSRad9J/erBMRUV7gMfuA4xXB8C
SQHkQMLfLNwX3YydgTjGXJSAHTEvw9GrVPrsGe8qq+VxT7kcnWLUAnB9jeMV
MGBChIgBi0VjvWHIVuaidB+SB5rlnfRaMjlTGzVNyX/vNyhDFx5BNloEcoFc
PBeAAPTp5+m6NAeClHvD2jQ7aI+3on43n67IlNd9zcnN7cndIfe2+pM3ovU8
ZXWG1zjBWUwQQ2kPjKWrZWi7nNMOvpBH9Dw10F9PZot/nYzs5p4Bh2WE/nkZ
Hc2wbs5ILdDgUsC/kDf5GMmmvU/8L8OEzUC+iYEzt9WtHShnkwP6tj9q+hDI
yZW44cEsbijMHOM9YDREbcKMRCCo4OjO5HJ+NM8pD0GWyAznU0Rnw6FH4Xaa
ZW+MgTKNhFF83jgvkt6rBjgpR/VciXczurRL36OMRyBnzwlggcCjp4PbnnM/
sUnNz38y1TYtEUraIQjOIaDj+/h6mw06qJYQ9hBxvywenaDLEZlNvzSZJqC5
/etQe4u3+XZJ3qcCMXLhlnamLYpMl2uFp0U+ZiA7dhW1jnLT/tyPpG0bV6em
MT3WJgyRKZV/KG2GnWtWO3dxKYtgyoei7v08jvtdDCcLkYATa+/LcXFSg12z
gR119nUjUdnlHJvEwWyg6at3X0qzfqfKXVibH72bCeWQk0tnm1AxvEkPlJ6j
CGiPa5JG1TrKNACZEzN89yPCmHPQ88qIo9Qf9vVsRu0MacIaQPJAjesQN05P
w8nWAgWfR/kScpCKsw/MFVY/dEB/raHgdI8ScL4qgr7/XfBDFybiHUzkNqT7
YY2rAemiwoy8r1N1cF3yJ8mGRzl7w/25XwpvthTrhfvqm1yOKXsSIE9bupIn
sICiTJfTt5sVGcOnacwVeA6PuUdnzpjReQXmLoRrcB33SbCKZcfom/8dvyfV
jPONfQ953mOweXwtkjKJDSwG2ecLVNtsOd++qWW1GzZ+AEfjqKWyaKgugUR+
ebYvRuZaoNOiMFzuyosPSQjhX6CHDLBsxTHBzq0Uds9xmoIgOhn4k14/1xwz
hgeAUTwO++nO9qsZZYj+fMLRFXOpBnVWjNWuIa5Ey75jppoDsA3FrtL1iWe+
46yuuX34wcV0axJ2naQmW8ywTl1951CHceqA3Ll/ey0u4xtxJfDRRuJcGK74
1OFzetRRQRK8UMX5CyqFNrmqTHcoJSau0Pz4rKXlZKt4Pj5mN30hrFDqCYYY
DxzpmoQGVAITg9fTotVEyy8EJV6s/afx+/Z/49Q3gvPeP2kG2ES+3iwE1RAy
zbhiMvWZ2eNzDSdBHwNR9G6+j9+X7cU5//EOcMNybSRc2suXywQ8CURc7DDB
74GbdtRi0jgT0XLaNwoQ5hB1HGhXsrSINHC/Z87rbeNMkxyS8Lwg0PnIQQpd
l1S3WRB3x8MH9nBkSczAimezKYaP6xu0h/n7I4XEaZoVORYKEEQbmPvvJFT7
zLlyl8aoluXKfia9USqs7orRjl9rtDLqWO06ZNPcRvsmtEzMXRLyNWLVcCkI
5SHtjPQPzHz6LHX3dhM5JfCC76cVOWZ4tac8pTYmOYbR0VSPUxuoa8ySHNPZ
FS9UR9MrW2sBD0IVAL/Hq+/2L9B4kp3fL8V+ds/6ZXMmrsPxIHd6jkVTNMxt
XMf3wV5Y7XwGXqVDe1DVlYzNAgS+fGtwgTzKK+U8ZmYXJC7P8PeWmHC6Ag0c
Swl8kiCzlwqPOuHhImtzETLNfbJOw22fJLLQk2RYhRcp9zT/37gjVX4viULP
FMVwa5X93x1k7U3pqMmWFVa+VMw8OJeXyDlQYGmckhyd4xeZ+FXi31Kr68N4
Cyt4KDAnx29PFUEz+0BXIpmvqcZ2+NDsSt6olXDAvLGRqRmWuU9NAuNM7Bv5
beP2bpL7Y4RmAPOVKXSYq+hbUOj5BrTZqgqHwKHQzQUjwV5d+Nv0m/Vp4H9H
BoVal1lLBQIfacGtCh15tAgl4j6rOAN4ZognZ5n33hPDHtydTSx+ZDlQ5/De
x1Q6C0lEv4HQ+HDGM/WtlWrsWy5SkIkzXOcRlKxJ008RMTL2WjZGM1Ya6ztJ
BjuhiEk0pPlLTBX/m/wR35yY/jprnOiG32TlFhiYQA5cfOwFKyYEAMkUIzIt
CusL2iIo7Emw9R1mo078DvN2Y8gIZyfwpVNQGAMZ/nNCSw46D8pqjLqMcGnF
NDDtAI8heSyTFW4rkMFB4U06iU4i81QXeOHLxVWy95mJeSaLCj3JZchKU26r
hKauzJZalutG/8b0gIJXv6ZOsBnrEjxxmwEsWpRQ9cBy/1shx3PQYQbKbXJg
ccAT/HUv8jq5ubVOmwequT52bmiziVoTPOd8ID/CQxzKgdJIcyTOioyCRyrd
YkkNLlc6G4FGTceELV90zHFgbE55EX3LlCBZ4jUIZLVtmCvF1N6WAOpvSFMj
dyl+wR54yEQ9Z8GxLb1+TArhWa3fHKJO+NC7dax5LRw0k4EAxI+rSHZN0Yuk
UVCxLgyxOdi1w/WV8HrjgFWtQX2KiRareaEkzR9FrpdLj0fnfPHAlsCS+REU
oLJUISRxRGjLuF1oR7cTOhPMf3GxoJS/01sZASSYd7+9xlHJOgUs7ZjSFyOr
FiMhpVSNgrcMiVWVqc8m0FZ/mBRRZzoH1nUN3wPTAOO7eczc2QrcVvscCJIK
f9FMZQVKRXp33UjzVF0/qdjb0KPVuxCLx6cC5Mko3PdL/h6Qr3NWCkMmaYkX
sOPH83STPYsuOoDa1P3Ls/PQHBvX/qk1LkfEZMkDoWGVMrTWnBevlwnkigC/
z4AqR+UzPta7vfcj8zUHbXak+D91jPCiHtnOUUN5ngLJ/L93wDyGzmPATMF6
YhXxMm74J6whgnD2PJXFcCh8nt4qUQmHCEIGnkplRiUyqX95Ze5siEnnzBhn
teGIri1Ta9LpRcotCP88Q1jQXkdewMzZJY1nm4uWavC3ZocClP7Wh4exdN3q
E/217Nlyw+UhxLoswxdShDBcITX3lQPOQvp7J7Fpe/91bEwY7vHPAdcDgDMY
Wn1h4rPGOFmwLW4DAB0HSuh2fFqh5+sm+YJ4XMNbe3FZs0vmYWY7kFGAazQr
qqEZ8xOvNgwBrEdR6k1YCuom10gnjrhZuL3VaxZHOVbMRjYqMGX0zjV0ofER
MXHPZmeyC23WoxTzf1dgelMuIWqX5Fv5hIoev8mLaGnS75CvLhK3Ga6Qi251
7SC0qmrzV5+QL1QSor4zCO+bM20wo38QyMdpkpeqEVDTkmjlTz8nhr0WNdlB
wUG9LPUjEz7/SSnbBE5Lnwso8GoEcsPZM5ZXmlELb4PUDMQPcq+ahclFF4e5
zQXHAqOmTh8xG5AnJtJZQoHx0SCCJ0aMPIqxggfNuvk4JwNZ4MLnhqzHS70s
QgNt58IM5ziL9GU5OFRTegJpU5E565Ec/xmzGm6WIlTITAz/fu9Y2/AvSM/z
V2iku8zilkkCXfQfUB7w1Xpolt6wYe25Pov5PSgCzVDYkmAhOjUetdWHBi5X
bFwzcXcmJPbv4acYYqhOlWDNn7s5ZsAwEqrufK0lIVVORbp5qnmUtMdxGrK+
dQXeE26pzoAMQieyvQbRRcXXG7yeox4QmnPejsfnDVxW/1Z6BV60P8Eje/Qu
8MW1cKr5o26ux7JVT0UUEqX2G3s1OOH8XV+dZGhlow1RfeaIOzitV/QCljt/
2/2Z7y5ykUN8mv9TQFgMjzRsHuYucemYEmO8WQ2tWoXIqTOG5pf4zRHAfn3c
bfQrzrte967HRTDtXyXTKM+l9poOLNvh1ulYNqa8i+pqGBWaRzOvWIpVdJ52
VViKqXhYn11l0UM7fCzoFO4xgDipz+HosPZi1g0zbXxjerdNC70cG8Hc7zjp
gcogs9h6X0T5DtoliN8qviaZHmIc/Dam2+DCzBLyONTjDErjjJaTw3KmU3Oy
9i+jxnXsu8TWPVVMS5hkkAl5r+5sbkBwLXViBj6Iug2hbXZpvUQe/2g/DBRE
hgUQKMOuNfI2CuORcgpjJmbgOf1MN/+qVsQdKjmWsfdiwO6wNgaw8nEXSgMA
JJ9iAOWVrggmHHQz4Q8LpjBsT3nYXC6aj3iOxqDwCcI4gMCNYlYvbDBZGOcW
w7KHYqqad1bHyuc3/EdaeT9wBHBZldjrCHh0iVLtllIJoZP/pxs+DIlVU8CK
VRv89Co4DWJapUTl66pFNjCnuQnRSkjSjY/uWYQF53piWmQf7fJKW1mLnuOC
0+5T0zrcoUpTByoca5E3HD2YaM9O4W/+nkkD/OZp3j2lvIip8xApaSQ5OIGj
dw/PiKF3lgo4y1hvZst4wd7XRF2g1JCRVjrXcrWhsoHKWZI85NxCFHGLQuZW
zkDHHtBl8Uqe8vPm80q+RmdZxTxn1ZCQp2LzKhbVONkd5l8GUhB4ouFwFmSK
/VA0YCvPrgyylnvS1OANyCQnIxt3ZjZ06IO8pHzZ0q3nWvq654ipcNwULh1j
uvn3okLDzeBxUGLOyzLhFMh8FyL6TzpI2MUwOaM3HEy+dhUb+4VfzUtuYJmy
7DNVKdcv0dx7y1vmZn07QLuR9bmvx/7NZyZdVVT+FzW+rWmnjq3ImBsGUyUl
fuE0lOnnhanu4ofJT1ccYAImPWjkGkw/e0f5fMBcz9k0zO4ASvQlIB7aQfBB
1dd5dRfdxMXTsWgeMLyoHc4PmDlO8hu1fPwgNizlqLdEGgz7+MbaZhsKu/fi
I3au/eMZb8Ogbc1jUltbLAkAIqkq39jGvk2apEcrfoVusIigR14mdhvlvRyI
cSaPPteIS6CC1vT3z6pL6pnwPsVui0mJA5FSM7dHZmezxIivy4p92vqmIsIP
3zXkt91eYVliqQCUmW0n3xB1nbe6XyvbLmRxgQdBaop79vpfzn7kOmYHgDPU
ZPBESn7ZA80IHUKnUBtBjJTZaqRV7nWdG3Ic28aKLyj8nJfWM9kaXBwBoIeG
/EhKKEHna09DFWALEXAS3FJJ1oBVMlBNCTDtuWUJPsVocWRYDYYGJnuNzXn9
es5T9v7SfT4pIWO0pKzmI4U/lfU3aPg6Od0n4OydczDpiJH2vpkykxqrvMmK
1vKQlCdCdmw4hZyUJOwlmnHIloZED29UYoNMp9qcSmj13LNADS58unM2Pfa3
0OkS9VcorGavxvhaLIXEUTfxcxNwT2jvAe+AMptTaSrqfYWCN9mVXAbY5Fy8
cRNB4ZXQ7yIQM3ZzYNFL9byl34hbtQ9gsiczFTT2avB/cAHZ7c9+q2SuYSof
5XNN2tfHCnMUdws/EnAMO7usd3DyLUAsxGpNqwS4/XAkS+nYQmf9kfY1ncHG
2mRc/zCKA65qo9xCMDXhj0FWHY4ku1tj08QHjX4SPQBP65ydTlZH48gRLjzB
uCSCeskwxje5/5d/sQEQLtmISuUGCvzpNg0PWy1Qko///iLFnFAn0kgxOduB
bwqJQeZgr/jM4FJ16vlJsgVaRfON+QbqzXicQqCX6r5apii4+89MsusvYxVm
jXgOINJ/U9FFEMCF+ObAemt7tm6oWoQzHTCieE7rOflPEA==

`pragma protect end_protected
