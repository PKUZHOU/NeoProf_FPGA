// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
DWBxDm/uXfLoglj1N5j2yCXz2FiHctBXD4b6jeKCMZaNggUHbQkkTl1QRTW0yhaa6wk+TILlr9Fs
eC7v6KIx12QX2TpCUuo/6E9pIytKIyKeHkHc3zffi4ZqSPqzPmAS/JZJ6dN1kIUVhGy2iIJAonXq
q/KRf3E2WklKpEFf4gQ4W951eDcOHFBo0n/V7wEuSdG8hx80w2opaMlRPQDhiRbjRgqaBjlCcN9Y
RzQIAa7yNgOwJZEc4eCb/f7KNRFEajUGy5vpHkLTl0ZMMU14t8Oy6Df4CG6P7ZbrT3tfXyEGF8RV
fpBve9yHe8NLXBEa+lR2xbdPUdk5at4Z4+qcTQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5920)
0VNwSRAHamRBpUxr9egO4lnxR7zPypEVbdpqJgZMS22LnbQE0NLvW89tJQhVGrxAb89hpGMibxj1
THBtVp4vlsAyEBRnQRpcL92V1+f0eT4UymIKZCrX4ACUx3PGT0+XRw5dSFcKSEm7zHwlPTBBVtZB
H/uMuwhOzvcuHU6suAzWx3Yzpe061/UxL+b9GXV3EHBeGtYBbOCgOCSqUyoXn80yX5vlk90uUJN3
Uo6o+wTA4nQPrvAk3PJ0K8UzASf+vqyIUmE+3saVEFzVmv8XiX8/OTQkktBbyS1gcGChy3l0R/F7
aZKYsnUd6fRERHkhbdhOT3NOVN7GcCWshAnP3Rzk5upJrTit+/+aIVufAlJEK/uxZ2w/Y5dUhxEz
YbQQn8FCTPUk7NlYQ/sykvVAc+tIcKPtME00Jcg8qlqPMQakBDHzmDOih/L8E4D9xBxgMLfJJHaj
mZp73m4Sk9YczHMfAztoTDXdtMX8yU5uJkEILkJJQlB/cWIqDBmrKXpPkLJSexjTaPOG6RKyiPy1
uQp9iL12QA/VSwjNqwG7BzoJVbJVmt8W7j1f8ccp5bYJ3BQvzTixU6+2opstX5jxzw2XOjXOEFPW
KYlUKpWCrwHc742M7fS0R4EzvF4w3G4Wqwjc885TsTeiF63yms2ZLhrVa0q7sUeS3yi0O/oZUol0
9xMrENWnxmXsvCzP/Jisv5FL0OmMzVZHEJZfFFSfdi1tagD5UEx769OSkBaW7n9BYLk9VDpGjknr
N+24ySIquxN8O3vrdGpvKQ9iMCuk8RQbX95T1QXQsDdNaeX+BJApY4CTBbAReTc6xYLCkjcIPE3R
mq9krKSYMxGguzuSS2rqEHwip2SMnaaB+Y7C3DKF488AY/mBeZ2pd3a6aJIAWWKbdUVkB6CyXzBT
wsBLXR+FtLrTCXD/f/ebUEkrFKdh42nNjJ1+ReiQcGtPdVXhfdq8hrQegMK7YoFeGZdLMZ97+wiF
JfVb0tSJ2oN30L8L8gsl2D+DygAXBghi1jpV+0lblAdoue3C3kya3NgO+GyzSmLlfUCiqWDdr+c7
4Kl3yqJpil9Im303dYU5v9IEt5zYd0UOvfdqQ8vQNQlvdwVvkWoZg4twr9WpowOJFzk3SH8d/KRz
luATvwwFc7lubOAs4L7ez/7zt+rexsSAOd8zpNsIicCjqi18WfNL5m29Gd9CMZ23oDBuPmx7WFhT
bTU3O3DI7WUpi6VQJ/6qlkSfXgs/maeNN2i0dYQex2NcZnoYsfX1VkQh4StGHyWFZKKsJ+fjrkmC
k21pOM+ts/ShAZA5ggnvlf2T+SmanaPQIU6jYl6AjeAnbLIYOAqgzyLEo9wRUQ+cE/wU78fazCra
gkxXkughruQ1fo4IpC+e54+pxozQ/Zdn47T3gDJS0R7Ms75mu1qBkRntYj6Xd0JQr31/a3QKeJh+
YnYUB/7eYbS2q2rC7t/gsouMDXK04OV2R5xSfl0fuypMPt/MF/1jxFdx7ZQBtdWzf+NHLqJMroeH
kOZmmxvDrJD76ucdkzn4TxhUZpBqe2YijGbM/NWTktxeZMeBkjk7RO5G8TaRlTzsgXSRvsy797+v
2o1YUOf6Sye+LUdWnbbQbwcXUG4CMc3ssA+bYfS5SemXNkdwxCsKBkaMfrVbVNnJj+hvyWrzdd8/
xgllBTn7+2aw0KMIQLGvr92Z+wAAalPX7+Y78hpM6uKlLzU6HWkR6zADLnpf2VAameVk99jmeaaR
D8ne+ihend/7m4bueGz7RCbrQMwrldX2BrENoLIVB1M0SgCiAC0KhTmUcL3ud0/6FYffdXgJZdUd
eoLtKxqOSBSRA1hJrUgiROkby3o2KAcKJLIXdvD47JKVc5zv1EQzuG8TjLBYyLkg+wOusBB9dEpD
C4WhsTX2eazbP31i5fVdvH9tfwkJkHOv7N7UU5JpA2DqevECULYEGYADM3dPRLNEt5aZBPm2COOz
t7NhkthVvLnseU7Ia6L/dawdlnEiUiYHOJ8bwzPHHyYrF0xx15ZwaP0Ht4S0+oGZ/LJ4W/r3gYaI
3iYcG70tovQyVqlg1RuYeteZCyy4dxvwjEAKWzfh1mPf5JB93/oF+5G2XS4CsNBoapMOcwC/CDd0
NuEXX7FCsOerGoPCMXato8h6RHh7XwgX0e6LRGQQUSAVz4mBt2MgHAaF3ZzBsRCSE3itDz0TuygC
J3Y/1A6I4DCG+s6kXtjrS3U4ub4dI99c2ffGYKMAJwQNCdEAH9n1xzaiRi9PQ5ft70YbCcsCH7Wr
BDH700OHHYCI5RPOyCIXRyUOoVMdd8VEQpBwKU8Id8hn502Wu34zhNB4Jus3+ulc/K5h1GCZ+bq1
7h5yoE0JxTQgvxuVlB7Po5hHxWStPYVU072GN6d4J88ImpwHqjYn0LHTk/ObCHPvI20/oAztYELl
9p+FfSmXOJiquLE9DT0C2E4g2Q4DHPq1QqQlzO1T9SKZhwK9Zr4+m+h35hfiZnBFFhGRO+MF/Z44
iFG9i6S/CRqSgCE1JsxCU3brjJehQJP0cA2EQJns7faHy/mKV3pREHl9x8NCqMVQjdcquXuMUHYx
Z6c8Gh0mAnItXBxR6SFa9JQNH9eZ5vxuII7jR5PSy/gk3yNc0QdrSbixsjpjXd5SgsPicbMXoKrD
qNEKqvWHA31DdeN2exEO+jIHIvRsFPI/De/i1RqSYjM8KqmkobjbMueT1U7Kv1wdKZ9JJJkfMh9i
2yGAELwMfuOvHnt/gKEetB9GVGefbH/Kxg4aFgOV5jhY0ns80gkR4Tqghzn/TSZWOn/Jtbum3MWc
WCFpeJ7SAu+bv0g9IiK2onqbF+1Gb+PbjRi6mIvDG9BHuUhLDUATLga9lH2kfVZmS43HA5KZT03W
uL4N6toj4WVUJnu2m1W6OfnIJJdngPNmDgmw2C4tpqIWtLesGcO2JJcqKg3X1oS88vjRlTb+//xN
n4++8IiE7FJbgDKLeA+b95UsD8O6LABLEn537v0eSwThbd1mszq+u0zfOqYBUTLXdSeYUmr5N685
lrQY2vtc+ZAiXs9K2oHJd0mOygZGruGijrNj95MDvfmlF4KPYt0eYhHYFwkXA0QCdlo92tt/62rg
d6HOu624xXiB8vpID10zOjuiYz1V3WGjkjhoDSoObW+zRDriKojO9mRjCbbTKgVO0pI7fOmvHfhp
cXNrVAi+pznm38pseqyUgaVoO87qZEN7IkKfvGpH7n1kXXG5l5r3mO/AZq/flhczpKOYAq6jOoDb
jM+BlrCUVXV20ziQN/JX90cxQksbR2czLRSKxqHwTRti2qn2dwF0dYCL99iQDN1RFadZ3ttGoei5
n33FQRPBU6nv4Q3pxEMDJmPOtKkxH4fsau4fBZA/Ho8IKACcoOkAHic2qsC10o+e7LlranrgP/kX
/G6Y4v8cH1xmnlZLTIL5VoEcMEfoMaRyeBpDoHs9/fUjOMSyL5/N1nPQmAD7pmf+49zzkMZ/7wg0
huVLeXXDrdlJ0brz9kpZIOpooupP1MqVHCQM/7NlQwLrw1qmfvO2ZbV/pTerIabqOFpiVFP/EUq3
HfqjT0A2sxcw9P7of8t/1yFgEEec4RN7mGfKTS6mxWv+gkh3VJelojdBxQPjQezLp2GZco/fTeHr
hPMi69wlfuSy9mpBoe5DxadkpZJYpBm6fh5A8HmBV9flZcWzzi8rCSVpvL7rVJ7hgoClz7mlaWce
7CmJWCb4ndfkRJDUeU8E3nvjfRMwNaDdiczc73JS6vMTX6tDtla+hvdT/DdkzYcQPbZRp+fCTWJu
FLmnlb5OCIVBO120gqCrbV+oC4bl8xUqciplu6XbgSC6GGS7CfYtUSKz6btDJmbZ1G+0+NeyCylI
XrU2rdwmDaSRxFcDpcTAUt3stqzpLVyAI/diGczrtZjDfpBDOywDLGKoW9q/zfAHLSplfiGu7Z2z
xc6bot8+qA8TrkNFmXaaWsqhCwIcdRFJtywxJx04XbMS1H9TR9gpH8SKfvHVBayBtMbuA4z0KFJA
/gaxxPixMa5jVLxU9JCs6HTQIctbNDKK1jSw52kGuv6tOetDuu2wOfXTlseW88dveLqlEixrMjAa
aduulR3jCQ+toXnrCWpou3bTpX2xJpIzq8HcnSZv9p0FsYnu7imGv2J2QTNkl2yzM32BEA++K8cH
5iWv06f0WwPqKhgNWB2+9k58bD7dhFaW5bI0Ku2Vu2U7eXYZdeIIokgBpMncjZ9PW0d7dA4bNCZq
UfspZ237y6LYLlYok7vvfEZ9T7XiCxjXOSO44iS9806wT5ySwugOTmtRTBMYGxTcjUX5AoQMkdCP
Iemhp//oSz7/VnXJwAxTk5TWH1dXYG5VRw/SgXa3s3of7C92dFEvzr74ZFpsEnrmhwEcYN8r4L+H
iTN5iBaapAjmI+oi4IMVbH9fXLI6UbdSNfodxsWbtnf6XKLVZU3KdGaQlXKWmjXl+9jqgiGsvjDQ
ki4AMZQBnCNT4Oo8rfo95VSjnkJUAS/kpNmJim5zLzCR0UygGi95+gUMAYNSo+GVoN+1yEkITxkn
uFPsvTVrwR2hCnpnmRI1rVLYn5LrI7E3pDJ4e55My4NTtMRy8hPGPVfoKcyeVgyJfNDajnwEcgKZ
eMCXQ7cWrTJK7GpeC3g2EJR9SblamSPNRojENxa+Zd3UJ6Yp/QcaFKQAB3Gy8i2YARtE2Sv5wOAF
2ijldPGGVd386fSfVg/RwCOztcDWCbYL+jKb9b3qTWukiWEQ8OAqTIjvQ9PiaBkYbxyBlk90c35w
HKWu+UvOd7mFPUPxlLXpXUZXyIU5geJkrDsVf8+KpB+EVScvIDfwrW2ifROUDIPCNQmsnIwfwkyI
878nU/F5FcusZL5ZuDMQKZops39mCvh/1TlAS7lXyBpqeQ5yymJSJyYd3O/CaVeXWZk0b1ymKIyz
mX2DTygy6sJjrmq1SdMLPxzphopnhDFcWGCYQSzPgHscVtlvO3nTPYP4TYNcPdQGvHSEPt4tJBiQ
a74gz8pINX6PbhwJhlAJdXRiX/CrXgGKqTEZ2w4YI0NzZSP5BVJPoFvJX6pw/ShhgCBgN6YyVLg+
D7ANUVzkxyIzgzAqNWVTvKd/wNMjqaFF+Vtpy/M6y3glvdlFfOEOsuD3d2V31OGaMXh39TOe5hwv
4IR3K6GzZy1NrJK91UN4SDKUh2t5NGFf3n2Uk+ao9Kc53jmP1wIz5f1BCr5zHZQXcBDlvSOvPSxN
hsmceK93xV7CpL2oPzh+wDCzY7sRNgtjn7av6uIUReeZEeAwp62HCaspUx4U3abQwFWZjYD7dpXc
JLW+p4tA1Zq2ie/yoz1O6OliHW44BcGOgxhvljF6Ust7yNnHFyPJDohAq5Koj/fNZQtqJRD8ZG9r
ls66fAwLhZ5RXc/3DIY+jha+eVWUtM2Xxc24gy8E2+Sx70NW1u/B0D/N1YvkgWd7IWDXgtrtnPLj
bzcrGoIS/NerXuvkwYwoE2+eJKgVYq4zaOWIAJNkyT5WlTT3bNZMbiC5CECWStFTHUXkBW0poJyi
XwwzZnmHt5EkBQlrGiXMZgdDg8Gj7NKrBLfpAfescSbqbeV+QuPrcjJxOkCuvd9qmQZYzq8piICF
kAlrO9xo43cIGOp5UjtKiz1ySSPpvad9hNf6b54tsEDzUWIfzfcqNZPYEzqAktLsnaY7H4fTR/WP
cF4ZKpeZmTFt2ncnbbAelEH0A+P61QS5uiLb3b3uJHnI8E5Itm/rHEPMGqTEmBhqXA2wypKBg8PN
3j/FO/JAGKT2zFYdjWt43f0bLYz82oGM2l//5q651zH5IM3fPaeOfvCH48Lyyg1PU9Wicd0i1cDZ
JS0UULeWQKRlLYn1auE+dcC9CPKxSjV2sqDp6dHFIZo+OXw9OpKO8OE+iMMfUQgfZxHVZlgaqSQm
eimnqWZXqecBZ4YlpGYGt/suS3SAuU1hV334wMZVwSlxgGh3Var5MFX6g/lhNDr+cS6jhkzVcGV6
AVJZfhhEw/TldVZOTPWS3RG0644Tvqy5AoCBPT7zGrP/kpZTDdr6/PtpGc6HoNPUnZZkQEYVXeQr
/Aq0LTnJ2ccOMLwfwlWDbyAw3lbEI82CvYkFeGqAEaamtIjXBYA9rHxLeJYR7mPulQ3sCBgna3xn
X/R24B9fPBUb0fmCby3+6zcdiUT+HKwzbWjhwvVPQDO5zGThCYBd7dk90iaGFh0InMWZMCmgWbbt
6LYrM5qQu/dJvjI8KhhYG13GGfcxne1/wwDe1eE78Wxqbe4JjUEXYqnlHot/+J92s6JBt4wQb0tu
y+hJPXudL+lLMsTqM8TSmdCLQTerhrXxqVvMRgFIYL40WNIAqGsW0ss2S0uIohNPgaXDrn74Rq8H
zW1nNHggSerUdgRbyU3mLM4ZZONoY7ehedJMhSLGxoFzhah0c32tJ35artQVfG3on9rnS3Uz95sX
uA0Ti1vnWs+1Dc2E44dCq4jF8q2Sv61XLxraY3HHfN9EnVpDdp6ED6LG3Km6Hph7vAnI2F+p1/Nq
tkDPLQyRWJdCsWj9ZOzXVlcub/mVlCY3y8RnjWlsnbZRb1OpfXzXQNPIAJFWKGZ+3pofBjo38I7p
TU/Lp3X/2GVjYCTbbAmTipSh7V3FtgySJbo16gg5TOCVe0VWcOxenR5lvRblhStiIglxkhzkoy29
38g7ED7Xgt5Cbv95uYsYX2YLmxrs48FV8u0y7GYPBOwuu1jNdFrllBv5ADTidxAfxPvaypiqU5vd
kGiM2B8vCHnworEHnmYNaw9sXI7rftyvWl+Rhq2l4qSPiPf8TL96iwERumV/frPLrNV1RR/q4Fdf
efX5JDQMyni3RSMJwxuuIdd4MuH4TuwFI+JHjn87Lt4uRHKlPM9VB5hxsmXwHGh19rrLo2pPNcFX
6wfsvJFmDEM7wjIcFPnxmwh2PbQL6jk7rMq8KitWrraotTjI+VFG0ZrnN2ir8/wkE0Urz2qqCmcj
kO1pNABDn4A+pjuB+JeMHlO+70bZBfv02nWOXIKY19IkoXDhTpwm5JIeN5q2qZ4Aheh6J1v5BR0L
WEim2z77qhPpcZucgVzM2/Zu3PubMCJTpQWTk+Lyc21voPPANd8aOKBz+YsDomGyQUpiv8T0xS0g
zoUHHcP59hU3EkOzZXx2vn3WAo6rUJ/v66ghce2bmI/CM8YL1c1EnnfzEcXFEbztptkeYVmwANZZ
nbN1f2LfQtrll+65UJUHrZCxT0MVtFsYG4A27E08waOii7ht2t4hkdAtnVP4tAfpMve3YmavRlUG
CDHrdAuqDVwHsj4oYY9tzcUjwq1mEOkX4u8Zl2HYKVJF8Q321Euz+XnxEc0efGwDw7Ep4926GN/+
5LvWarXOHkV6wm6mWg1zqFIaerkLqXf5n+nz91KSIKgo1rW3dhIAGsEyjiOxVVgQa7680shha2iA
juCS8AmdjL4hj46Sa94oaf3PGRppakPfioNozs2oZGxE3ZuVcqEvF2YyWAvpIxxU2KT49R0hAmgs
z7c42EUKDY+k/p0kxN3rQqVZk5uOA713uLfpZqH2HUfOPyYpGir1zsuiyVv5pkXdNuwTyfcuMR88
M1hArVUtheloGC4YoBLJ4JjNtpWp2bQmQqhYzAZM9SZNexNiQhMMqV7jeW7+B4VqGND4OL762ZdX
iguDefWwIE0QJ/Ah2pE8nlCRw1b1Xrs+t2o7rAuIaANEgYbgAxmJ7w73hCHjLzwL+1AO3BTLMzfr
uC85fmZT9YJ2by81R27HQn3oe8tDd3usgMAXEyxHC+UropFZXJ5J/22KBkUgns1oDBdofvDlvIV0
6/6lBsx/RDWdevBKWu12pbLsZS2NXxQ6syIdwxIp/YJoraXS3W0V6s/fe9JQcKl5pA==
`pragma protect end_protected
