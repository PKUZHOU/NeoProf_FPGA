// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uIcoRnv8nCC68zLocnfZ4sFGQFfBmX3DCPp+c3uvlVxyiqK/+XpWSJ+sWcBS
ZL2fk4GJlqq478ZDgmY3HZg+0GOJsNdcrbRMkG9MDd5tO4NTwzYCLHCGxGZD
F7QXOig8veePBcnP5njO+kmNQq3utW6sRgG5hhyBp54Kz3IpD1/gV4pR4Z0A
B+GEooGGnDErYofCCkq95wgeHNf7ykZNY89Itspbdq5PWcOuQeh5L8e6er+8
jQYeHMpcJ6egQh4tdLopcQ8Tf9fm92M/ApU19o/WW4dRt1KN3Ej89IDZtN8w
9wgzcgdTY9Q129cDy+p5RL5oJWVR0r99qxzxks4N1Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aiMa191yADaUhDxn/atKYP7EvX7yITJq0QiKRLZvfX9D/sVgNjhBignrEyVJ
7XKb/pjXW7BEbrNlwmHHLhzuMf7rcg2D5A+wPcoEfbTtwh8f9Vp8VHN0PhmD
1zDQAXfqBtd9Bx3H5ZVdJrhhMa4w2LZPdCCxte6Vat87vXMzA+faAW1O8TfH
XJ0jbuIDT8uHvdTXgaIZR+dh6DBR3L7gb5Tj8jqRzucoxdEu8tzsVQRoJXzA
or/B8vA7QNuR0Jj6ocCB9blAYeZHfPA2Gd3h2A8EP3crecb1erWLFaMMovUK
tJdZ2B4YusjcUq8BnKvuqHDW72scXCOu5AnxKUTmNw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fuZwLNo7qjtaRHdQja5sAx8M2lA8axkvLq2xNb1FFJMl1Aoe6a5/QNpTAqmB
6GL4TyXp/boEl8T3oPE1eJwL8X4x3tdmiCjN5z2iyGnV+8MJeST3Zu0XFqF8
W2s10QgtxCwpz7ujzv4tBXu2UW2yyYBkkswYwU027lZX/lVQMCtv2R9Ucyn9
OkQ9zAQ61bdNPjeOBOQLl2a2xmF16raBRlNAF5eKm8koHvSN77MOdlECc3BX
Yh75DAXUgsM0tG6K2iv2aOTqsFk4JWJakWHxwvSzeDeIuNSkk9U3jZlVIJ+y
r3uv+AP3Y1y4Ka4+kfhFfxQgm1Z6qcYJqOEHkMWUug==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NUHfXxuF9olPnUW5tg5jpWBveTqTlR/7mCtSY7Eo589YCviln7u22zsUQ4D4
wCrpdH+8XJsDxjiKtTSACRMAmbDSO28+erBcdHRdqRj64MT8eDsuUypf+gD/
8IHmh+MLr7Bt1vvzBdJW/OCSuPD1QPDI520A6j/2urGZtKCALjs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
kqUSFZ280aG3dh3pye6qFPBXHwKfFu99uQIdzWw+kYX5SN/pcJDTgdaqCk4z
RWJBJy677hJx2nFlskr6OPDu4jfZDEJFuGL+BIqyQXplNLCr/8vOs7WIKZ9D
h9n8sz6f5OcNnTLinO+WXOpHGLsL1QXbuSBIwva9M73J+nb+Rq3SUxDNqLnk
zTBPTc/8e9LJAu7ebeWQVkqGpEhsXQsEBac5XIviYGaGS5ZEqDvoVfHsOE9m
8erUlP+R7lXgKQ860QHa1Lyv5Qeu9oLf8wcj5nYajZAOCl8Al7JTKukztRv/
qqASGLrShBM9VXG8494di4X+6mxSG7qjHWz2/ixaE0/vARD711+RwZ3/v0uq
ASwWAbaZhyBwA1uCg030VPOAJ2tMFODFKdvpglLyk/em50HtkdDmFHwP+73Q
RFD4F7eWDsnQXhmIhkq4XXQe9DeEmQA3szOBZzVP2mxQl173o5Rg3dZvJfL7
JwDQivKUQuwdZm3DcRXqCkccVDmcsAYH


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tJsYHpqiIMdy0fZadzMZtVjtQTH9xUTeSHGxKv927H+WBgx1AjotwYAmvwHo
LAka56sOFgfBTGF/oKEU1A+4PvLzSAgyLj8IN80JyvqlvGsFjehTKMpqlBO7
9OLeE2y1+wzLqWFh+dteMuOooy/7hQ4JNzkLLdssYJETvjrF+/M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EzgxIARRdRW78yw6dERr6VedQel6y9ez5eDugSGaT/przKT0z5Sn2ArmppjL
dptxW9rZPLy1KSeUVx/YV974uuEdE5qIEyOp0Q6NYcFgHQG8VG8eJEWNubOH
BwGxHbgMs/d0mq0mWCIIpTIzza0wpIiK3RVRfKrzAckGOHGxcTw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9024)
`pragma protect data_block
S95RVDZIddvKG1UCFedCHIEjPT1vt2MzodcDnZsqlxyymH0Ff0/umTJR77r+
Ur9vfDUZ0z6V4shHJSwR7cvAoN6G3vgp8+oUzqM9KW7adkd2A//mkUBU4njx
XP+aCY25fn1R9FDPVjg/ce4LWBASFOaKLZxIDw1mJwfE08ENLmM0WYtEgcPU
rmQvWkxkeiCjpyAeUI8OjDxgJSO/LfKPcK2aVxCuqd1fY3s/YqbKEErcd9xG
fHixrbc0Dr90lzmJQBQIOTB9asltzF4Z9DWLbHrdi6DF+/1DPR2xNUh19UzO
IFE6BzsPmWmx9to7DhnwKDfapiIUFs71st12s4KjVej6CDCA4JIrMPriJuuc
QiVrPK6vhNNLWiVY49uvDa569cPIOauk2oNr1baeA1qaQpHibWyxJ1vWIwwb
Iws7UEQWS4LnqlhY3yik/xayB1ZuYlRXHV8ev3943e9Uh6sX+dA5SzvcRGXc
IWE3LBOOiXQyh9rsUZ/H44cMvTQ7+Du+NQBPpp7ayfMK6Yh3LQSx5or2VpUG
x3LetuPHVbrCsttOpaDyv4ZCVQU0NU4zysRSFOKAbEdXE0puParaUM7xVv+x
h6H05x/XyUe1r7KISc1/uFsTwWfUJt0dFctSIVXBfYcG+oEYA7No0v9ecwrF
ibKPoatHK2a25mV06RYif6aTxOQLOZdf46iAXXhnDT4Kuz0U7xDlH1mi2fYc
MH1FTnDYXJOq2mqfwVX1S+xyuaEGzSgCgDNaQrmiy6Pi+/O4KoZo1nzs076P
RY71hTnCdJQS6W7HTxny9ZK/S38Qw54ri4m/AVm/1Jva3/WS66rSaEgTYsfK
TJqOWqcDL6V1cvghpuVDKlQrepsuqw1F3/gT3qHNRNZCt4V7XxScmMpr14al
GXYGXkgFn5hgnFDym/v2sndCJqwSspu7W2UrmtWd0sCUWdWPMqG/Sd5d4L/R
D1n00VdJGHXmheKEJkNJKEg9hHWBZdxYZDPQnX28JaX/RLm4tRRIDiGqA/4R
YgdZ4mch/jNtg50YSWeitlsuId4d3CmMjwylAbYXLAYPWaWlwjXHfHmeaZP6
KPDe55N+kX5t1imzHtyA7Rn7IpJiLc5ZteLL4VskitpUI4rK9WpjaZIQgFUd
mR8dMtf4RSJ0b1m0pq4wal7xHYLfa8vmNsWRFFEptS7rHp0x4IQWf3SzZOMW
UU5BNTh2QTJoqlhPbKnoor3b0MOKetRGMFCF8GVo5Z0W6gdNJG6QZJAyeP7o
+wFTFm+6wBK3ZebHFReL2rdo1By1Uuefx2tzA4hdsjcXb42BAVl3but45HA2
XzKw8+aiJ+/j9n+5ZLWWp3B/zSEoLk8MvU7v7tPMnjwPI/PUwTyhDVTXzDZB
aGHm4P4T5bY+WbaDhvPiDJnK3rNOGITVB9ZyferbHOjT2VbaQpOjQb1Klsz9
WiVKIP9TvjXkmBnrWxsgNv6/bTLHaqmpV0dEjDFwPKGJQnlLYVCgQzUBia8G
68NVOulCSevEdVE+jeqKGYQP+8Lx7lGXXcGAJ+TsdYLxtma/hK/T3rmeN8EC
tinqJkATKEacNnuk84SI2qkLEH5Lv3PmAfE3g4ZYwy/+OH3DerUYgZYAuB/b
DXf1XYNgbXCPuSiFFhrKV8FlpCWUtqFyVHhZc9B5M63BFN5olKO1coDwT80V
dbw6tFbVBH9F50e8cn/JkQDtmTQNOXxvHsYrhCbevGE+e98uILJmm+k7MZQB
zEZcrKWENkoRW2jlXj6LhLBgAwBKo67lHfoInXYWVjRun8Jj1CbmpHmWrf8T
cuutixzDh7Ka1alDcT01tjzIDMVD868kwa/V8s15CwLZ36DB9chwl46J3vhl
K7DKoiRogYkKn74tqbvORMy5Fed1HtNDqWijDEsL+QZq3Q0fdWGci5lDvfEw
KEBjccdaKXyee3vj5tOzly3qz6b0ROWHtR2Y7a3ULLJ5NT+nVUP9RqDhzsZN
rkSiudOqj/TPO3i/fgoCiUd/oQbclGKxZGG5nt+LwlqsKyL/6mTGLoabGV72
+g27+BTmvnm68WIqLhG+yAoAHXVBzMtjoX2hiI53zByFtsYYXPFBycQV22p4
I7VLMlZG0RXR90dv684oT611HipFpgnRG6KNGicqGuLRaUI+Muc4mwwcxA5B
P0TsHbTq0f7M0YWtvztNJaCX3kbPkk4YqkekiRRxTilskN7lEaa5M54401p/
Nz18eL3Jlq0O8uD2Lq0DirC6r4JYy1EtKEOWXJh7YTro9XLIcp4YoBtfTX/I
cX2XvGUJd8VaCzRqgpk8yw4g5cq7sILVxXoplX1IO/v8N5sv2EhFw/8b9+DI
Q80VefOxz5yJJeO+w3LBKXjGd1JRt+ODYZ48WmW9gLbjgVy483RGBn+SP1eO
8wrSVTaF0Ld1MW9QkVCWRJeiC5xFwbiKPkYf4petuZnQ4hKW0W3ahJ2SKugu
dOl45x58rENg+miuIq4GH0BMn5rGnxhGIuNsD6juadHpfieEzzVYjcfbUAPF
9Mxi2VGaySV3/L8LZBCPvdJbBgxt5rkHBr7QJ92gRksN1yV+U4r6N/81yzZG
j8vD2D/ICtYQAudZvmA3VPXvKdcycnOYmqTe6g9MeF7OxnTsI3/PDdPooUkd
euLcLrl5if16kFx3qqMwZPptjTBx3xLKb+sEb7l70hYlD9uZcFADiGPBWncw
PNqvRGZFEcLdbTYacnsUgELiDwhfh/OlMQvA75/USuFBvon0O4Cs4jOo8TwH
59fWClxdAfKFaS4NPpTEJLyLdRS7pRJs7zBnzsbsbglQNEFfMUH3233IDj1U
sowPzvR5UesWFW8aO70KWgM62ZtJFC2XNuhF6Xqe+9Z7ORY9gL0fDZPHQYMu
+PqqsRUA4uIelV7ISIIpvmZcAPQaumLUZxIpeBB/tLmhyKE6L1OfFWihxnWc
lhO4f8NaFh7xn0ueGgujUK4Alxfxbrm3hN0+BQgPIcJq7lte0hO1m2E+CIpX
NV2LnWXhqfEbqimpWeui0hzNn9Sdwb4uo1+EUUFbDbRdLk1uUNP+SeH3JT9S
uF8NGDXvsY2bJuXzEc4haL+XIVffRlfvq0NSF/mIev1iyNUK25a2Y77gA7Kp
O4EO8mkfWOY7hHF6OEdkDI6FHsggRGG1sjzRnyrEVo0aTYr2Cff5VGNMwuJz
C/I3G5jvD+hm6aLZObmXG+2Nbwq4bWDzPwHBmpuUDCAFDjRlx1ly3jwvYVBp
uHEZiucAmi9FHGQNQ0XfzX5XHcNuXRl9ANe00+9/jRc8YfsDqohkQzfC6/Sq
6uFUTzMGDeZNlSy9i8y7mYnHDKX2LbaovUQ16c9Rcq3a7jRDgxtJVcWtyAEi
Q0pztbv9syMJEZE5wNYi3L3Q4NQhni7PJ0nLAFufdCsIMivozH+TG2qbKLMh
q+zbk3CXrFFmFSbyeedwlkzrwXZhfHjX1gmQ90VY+mPMj7axlFYi6xdwuPB2
6ps6V6p9x6ovbixdN41kYABNPQog+P+k6yQTLlr65DNaXgo6om2rLI6tuvwS
s16gasz4AVYNFlbRqTceVZkbv6WDkLWapNp4vDt3BqjwV/Qsnzc8J7HDWAia
e9layFWvkJbqZ7gNjq3MxZATz7pJymPitKSkNaspZDQb4wFwavE/evpXflno
3OjsqzctR6ztsDFyVxDQpLGmWiLrebkZkqqZHI1+7xFLrY2p4+vEGIl6VEHK
HF3KQrm+ESubWb2Xkk0RtHiVuMN7kmR/PFKDcNVcDTZIWFZHP/xkmRfCK1Kc
dNwdMr2JiUOQCx4/F9iZY8SPVqQaEvT9gJu9YVKKAymBIbvROmML5bCrBEcd
fzckXSQwWzQH+KAHoqKPSSnaG2CbnI2YrOVR8iGOJcbVxu8DSQZVJn7aN00C
MRlk1WPR3mW6VBykba0JHzf9i2bYS7AQIg7mMy4BDVT/xayDG/LE6CHX4zKO
ds3WnXbHSeZuwnPcHgJP1qrm3MWia/uxcIXbFoUt3RJeZSd7fbAWywdMz4+m
yEwfhpRVozs8bJrCEcyty3XPYGZ0piRGWiB2KuRKj5itAJjlhTDArfRAttVn
7PeYs/ofHqZtVt1cQHRaLtKTi9JKiQgDOpvEH2h7Cx9uy3sdFe1SLRoZAFHf
tJO+vrS9JqNIzUd4itVBNGAcx/IVYvtRj4jtNRDEZgdxcdTcuInkAzI9Myw0
+2DL02JRf79P/Iqdh/sb+sg3QUyFsRQRFQbiSm+l8udqCM8GxZep+T22IB/6
K0BsIoUR1n9qJB6NZSwQu4Z0eD+qdY6S9OwOpZX7SkYX0kMIMgF4iF1QMPZu
Jam/nNZMSVNb/VeYUwEhIz6vn0jdxi36C6peckjqRpe6kwl2YxpefBZQr7D+
JNazSGqY6VvTZwxqi5aK0fR58nsOEDb9HLzvIYJ/z/z542jiYJfsD3m7Lwwz
WMCAesG1qomb2i5DRAJCzHWovRf0TYGB8R3vDcqf+LJU8BumLl5cRu4LdQYp
whCRXPjQNRFcK/sImrqDZeYlLPp2tB9/pH0d+RMFgOYvXal6vI44WjqT1Ngs
pe2cTf7XoRCqecsTDRZ/xNH2uKp8OVL2Bh0bwXiaI3IJczEm4TE16bU3wCT2
6UuPKTS73YecWtF6PSula8PZiCilPoxHMYmeW3ePOh3JLGBG9DfAKokaKI1C
UDm9Nx3QMkECxP6/OmNLKSksL7qZdx8OGITYbFyeJ6vy6d0HCQEZ67kvunAj
rc07Lr9NqOO0gfesMlAF45CACsX9d9sOi+cT78ocwbP0MADW6VViV3DE/sGX
PYP8FWxe9crcj44lcH67xUQEiiykyCaFYLxXIVrfbLbak94KExUfhMokbkTG
WDDtpIlNW7oaA613Dxsq1d9SAkOZRhjdAcK0ePDXG91b2FGTLwlk6O0Z9cfM
DrJ6MIDbLyNwG0s6PVM7KV2Y8W0Dp4xOYDF636pQn1eVncKzrE3V7t2FG2II
HsqfQQsXBRc7bLIlGUfB1aejB0HQ0yMLQYvOp1G6bcZzD2EBpPrIigKYFx3C
w16RoTulFCp2yVfVWWe4GaIwFJ/GoCRvUrMr9YBePZ9T8bCZT8A9KhFnvOqL
QHPhxU6RsyWHRYwk9m+Yos0HGgQKCQKXGso/vASbwP337f+nCg/KXa/E6bBD
2SovwlRpcGLGUuljk53tuJYzHCXivwnyLjnfvdGr+2wJRVHZzjcmtHcf/UdN
i20gfY17WdnU7TkLY8WSJFqAjfKhLJhY7e30vE6HcZ9oiisc5MYJMPZTzXMx
mCLUvGWNsJnmBcaGnXZldzHaKKebEsbM5BmXs66HUJUtaobtyvwseKjUT+o6
DVUHasvVHWn3IZkB/6MjNjyyzOmUcGIXBaWhVzfXjwo3c7mdC7Tfk8XHR7kc
/KtlZusguXvXulZexdfmHGxhxdruwnngBL+Z5iBhHabrcNCwcyffOsnk12Ul
f4wah2qhp3MXePfGTaDqYe4jDmy1KP6aggQnP0F44EXimtWspFRieyynG+Jo
TDmcu1roB6E8ZHcP+pANTvNGASCvVPCZGaWVp2aFeTM85ANStflNJO9enaOy
H/9Ozn3Euuhfrc+v2+fr9b7N5yYQj8dH86U43DeKbjZsotUYXhocKTlvo20E
pCPpz4KeScceB2Uc7k5SFkRLIgxosJVe6kbHebKp5arID6A6za+BL7/7XV5W
nYCHGmSmj64FUKDCQAJC5j8S/g6+OHHkPncRv1YpkH2sntV618VgHQ88S2WL
/7pujLZ4gJrOxx7Q6521PnVHUOLJVSLNnaXkzQpiEAfYlBR+RcMQfrLQqO9A
QCpPxQhxYSfyPlfyvupMjZu+UcXGYVo2JpyXQLpdhsa07gM8YhwwIXLw6nDv
QIdR4qKlGXpqselxxZyGkPXhKOmD4zFg+NH8lBVmilg8Sgfmv3d162NSmO29
/fFJxHeeaKbg2Q/bCkmHODCsgFKuGiMgAp2xKPICz/wknG6kAJ5fxIrf1qWZ
R3a9msDhog4icBWGgyineFKkZaojD7bDtePrf21szliYnWJ76lST3Ht9W3uG
bqs/1yPBI9cffYGcbNCk0WfxioXsXdLjFBhusEnNCcCN/dnR1g0Yo2PqGOb2
2Zh+tqaFQHZci8ta4cc0UP3+EtCYL1dBL71SsBImJw4+7IJ0uS9f74k+7ZZt
8wAGm9vi6E4tE/YMmM+a+IrNpHUg9ZOUpR85VXBxmuDGYwY0XOBIdBfNzpV/
5zCj+2aU+ZTyWpRVtmF6fNgc+qIw8LE58Z/YlMBfXCJuAJ06H/23p2t42VPt
s6MmthIBc1BjS1XlpDuDLL8qi6hdwEaK+LXNDiUyBdAT3f1RKfOSOOZ40tKg
p5oE+/Y6OJp7wvqCHIPJr7HOcUn2TRRZ3YEjnIArBb7xtPDbd5LiNnCe58Co
h5LCUcMiYepWBKiSoB5mYqVsf+bETNH1KUqDPu6IowTPNwkG+PGIKnGxCgm3
Lp1CptAAN07zLwvItaPU6NrAe09CCi73HMlnMSBrf3Iaf4kCVN1Yv+/XPviA
8GkoGUOjZ5LyurNbp8MBIDIQf2apd6F7h3qumCD3SlYfoeyZ0ScIlmzEbXUy
ywbvuh4EnQehoiyUX6DAsBYdScxyGzoPkmi5Jt7s75OayPkUGOhyEg1GCHkB
cHJDVzwFFo0Kombw7XmsGRtI9j7fKL3CJnmTwpjQJnZ9yfxywMUs/rGlDKq0
cVCo65m5uNM0yituJuwq4VaWoDK0IXgG5SNEZIe4SFhVfvac9+SjgTvle1vc
vq8FZKfjOBtKt2V4otlr0Eugaqu0YcYsFekPPSCQDgIo+ihDo3/Ak8TaLvjX
nTW7o0r0XzznkTJfMgjACFzJxtYIB2K6izcmzlxrINwU6q/TJbZ3V4rsVayZ
TYtmp4wTIRgb2/z8ZKQhRpEDaRn73MSG5huHH0zpju5/ZLW5kGYHRmP7GFkH
emQiDcyUPmAZE0CjrFYL3KJu/sxJC+GxcuJ2IXF0j6kbzENsbwnVAJxIMrJD
7/IxP7fUJtrezK/rsF4ue12Mlp3/ZNU9n74yOAORr6KYnWonlvn1w9QdTwd7
2TyY8xXrvESNKyVQSNmkb3VPgOt4GMmKSIPj8IaXlae8X56+eJy6fraIBQwo
OINaEgPTv8Ak8zelpuGMujCyQWo42kbeZPaPzb320wUzd+NtY8zo2YJYDSCz
IxfkolDiiDZ9iJd2ydrmw4ajVkwa1gxjoOUD+B4o5lAVxHFjm8HxZJUajUVQ
Bd/YD2izCCi4BAQviKFkl3zPPzP+yTgAsTg1qB1onlOrkFwHj5xC6N8gX45D
RMRdo94lGnhAKbpiE5T6iRoVas1KJoatNtf0II194xVJZmGZQDLO1WJ+uEwj
SUVACzgeweX9sNy83ZMn3AMebKPk6TFwP1kRZsRMV4Ykg3XH7fYpkn7wwD/J
lSFOYYAJKbQuWIWxFZ3rMUF5wmn7LET2prBUAkAUZr7WQ9mx7sEpXApTmMDD
EB0K3Sg00Sen/Mc43XVuNVkU/nB1upx/V3FRvHSscBP7M+p3KhOtYQyW3syB
uosW6h8N3mNAYsEhwO2/qzHqYGEC2wo4d8/3ZGr1zwwrqGQ9D0n+W5W6Jv8L
S/3qRWgJsA+JPbJ8L0+UGSzppRgn6Sss0rCoa32KN6h3lHmMO7UP53Y6P8jj
3fTpUGkXiKGjfewyVa6O0XslCkrb+4gcDsfbqTuereLuhlF/YqhBNpx8G8SK
pOOjkQx+xYXPXs8R7hWddm7pz0tixRtTXeUIhDsZPv814Y6aC/sl9V1csk2y
DqnC8U7WKz0fDr6SC2BsbAZYBN2jIe5MeMWfy8IQVuord0IkgcVD5C4hJzhl
3p6dN4c/+ZoPIyVUF5DsvazJRQ1ZGY0nrTBUkDjD5q5k66kI3zWEbegzvzfY
NZzIaYBE4lC6FnXPLS46BhVuAc57yYhnsaOdLVbdkvQCk0b5uDuJLbNmVk/p
+LI285iQt6ciCWWxX9PUt8wXtoo5jbWAxK0jdy/ZuGydNqZBsfUn7VeFCHp5
LtcIs5Mhuq/MNoqcZz0hmITwPwi2YqGQH4A1vJN8PHx6c4249BrFN9pVFrQx
Lzo6A7SUNPqA1WeyDHN0TtMFCGSQ4ojE9JDQYSnIk7E9sdalwTm8iLJka3un
HcthooNnLXpES3v09mGB7maGNy44O73TLNtehtmD8cAAP7FLlocUmVxSXb4J
pIEEOVKxyqdGgUHOGDhj9mLVHbewk4KJi6WgwGcaAQUirbbA9jx5R2qHDwhA
120+hDB6Vbt4HIp4FdBbYTm9npXK8oEFxWo6dZv1MgDmh/xpaKUwJAHkRc/f
MurkgNu+cwjIp5P2Z3bCfRUZACccbt2NSy5HH2CI54IkjQiC5P8o6qm4iRQv
1ochNSlELvdKQai004xet/MM24yfeCDRo4KFB06D5znofwXo3vtkqbAajFIV
REOeKEZXNXJJtHs6zKYZ6oqA2AoEsCNT/mqSX5Wo7fiTKiY/+kB83JQKRlJh
8HFJy5qflIqOIR1F0QNLuv/PYGz88xycpx1Amhh+/TyLT1j5G+8INXlHLJI0
fcfGZhIG2G/7HYrx8zcRgO9NkgluMiA2XOrUGl4b+4hFKnQlLFoeeDl08Ngs
phPzUwktZfqNRU1W/TnF5d5zFfqCd0TJFaKRsq31T47zq5RrkevgxPTynqSo
BcvkI1Lk8As//xH9Oq5kDrskP11RZEqe42br607L4bczItTfUhv+HhQh/J+T
u2ZlUE/YlUiSH9jbZMMdZ7hd0ia/luTzeuSUddtX0rpnUSV7iu+w8f/bDTm5
33N0bQpaapN8Ia/OLblQOdCG3yCfzMfEJyBijRJrGOJ5DKcOzbi9g/b7XX46
MM9pmgA8jmVSl4CD2YvBBoM/r3WSdgvvlqWJmR54NLCOgrWK6Jb+ru8NS8w3
ij8obhf3r/LKbUZcswJjNxakgHRTnhxaarcFBFnvDKR6QeSej7k7F16usYIR
fedscF9KeJY0BVzvFqvLdSkO2wAcX8vNf6BCMk9dgiEjJ4gn/oR/VY5j0uOd
YntBmFdRFJRTyLM8OwF1RH6yryrw/k5GXoLxz1yPw+ibtQg8XU3mDuYzqBgm
P4fHXf8LBZnvhu+WePOn6qkT/B+ZKcrqoucTYVeQ7RNyIxkOYJXz5FvHHjcd
DnBGEaa3PvZJ3O0jk5NCi10SwH/P12WJOtiZMVZCciDZDx0gF28V5Zgd12Zv
q4MYCyxoXfLd0hRYMHQtHqNlOIF0Lb0zhC6c6atOLmwkoiqxF60bb0U1Janb
HveUYimz8fFvsxyb6dlSwXQGgd25Q6sC0k/cj59hBGLYhmDU4upnCc2njsPc
yiWH2EwZA6WLrxbtNDI3Ef0p1ahC1oRDdLTMvOnmgfh0ukaEsxwiW8XDo0Tb
/iODs3MMXF/DV51boTq64BGcwavQZjwLdy1y43dlcnAh9hzPybi1Rz4H7Zr8
83I5fKMN2Y8INfoETE9va0dUE6Uj7JwmCwtu4mgYtRldSfNnYo4qZP3IU3j0
jQGYqtnHGYlu0Cft9Hc+Oe9QYWY29/NeZXwKpmsvCzOiHJiUOo8U41Yc7uTR
wQJ/mRlkmf9nl6SGDSptQ3rtyKII5xaDK1pYa1wM6YP+QopsiN4BwAescWpz
MAqpZXycNyrLQ5Yt9eBKSU7CAENrr+JiICKrbYMO6tWC9UKAA1MFAy7/WHWM
Camx1XXkMYEOEhSXREpPZpIFaDOqkdBl+30GyWcnMn8B8hemoZRWACnAz21l
wTcOosTykfh6qH2f8OQBxfv1mroPnMYPaODPIaPJy51xRVVtrSjU6NjPH07t
GgaAcYLnMpFBg4fMQHi9B3P3E5c8cw5VSyx0S/DnJhEazMeNkbMxEyJkgyrH
H0APxwrxYMLi49tXps02JXbBJzJMAjCNaavc56fnZq7UhbpRZE9tf6DocSwq
mnLNrkkq87GFz8j43gTGZaNIu5a/4Ws1IBb3Bjo5CSd+FxTR52P9s/7mngeC
fN+4j1N/n6sGBDdKjZAoMnkenw+k5+suT67TAEuS9hiCG+BzDZoqiAadbQlE
PnaK7cdk0ElXk7Y2cx+Uit6bDfnrMJ8eVj8ACF91oVYu/PUu4+N+Tcy+Xm4R
QkFhkKPtzxs3nfQi+XWRisiNpRDSDPo7+3bRaM8nx8SwzYc89dZiZx+H4gpu
LoO6biiaVnmyf3qCWK3P11+yaOD2yMjplGbtTC0xEQTzeziCW8S4QD3IIgs/
Lm+mIP2oGqUE324+dbRzvVHpl0hX2VkkkGN8Ba8hbTlByQemjoGn/xSQ8Y7s
e+iYWBjrCUKBNyPXWYC+trdYe3exFVwJxjsYRqFe4udPPz3MFlAJ5x4MO2Ih
BB2dtm9IIFyMGlQCV17LzT6SxIeRARHnnchlty9Sw7wBHTkWcl6C4s/9jfHg
JPw3u6YxriyqszoGHQ1+6DMVgZj+dI++/pjT//F/4hLir9zGAP+n8scq7eKS
pGWhao0Fx9uJalNwu4GVSd7+3/KPHXRNGVr2ysvg8/hQCdhvBPggrZG/fWWf
gqRPrAe8ytO1SxvRs1JShKcLlqwAFfj8btjBqKpPDfuZ1KAFLT9AXVtoqE7K
tJQejCGO0jDbVf5QquL+oar7fQzuH6TkScbWUCMBvyN1uRDBY10dRoP5NZWj
FBtX0vePqWOlSVnKkdp7y0wC5uZr9Q9hrhYnfEu/v5pU6hi5D+tPvgdVschA
QsI7i6vRziEA0zp4zw6RKUkn/u/4NV5PG4FE6DRBVuMJ/X1ueOBYi5rswmn3
TPBSNKVSWNql7c1FeVR4ufUSGN/CUgJIIYYgWl9HvfEaStGjXvIfDJAuTYQd
hantqYljaB6fnpz/KzMm4QkSeexwfZgCajw9wxuEIqhEVHJ9Zy+S4cm9K1Bf
CHbO7ciYMghyI5rDPmSdD8pbdK/PZ0m2uCkyWeDGirzHuYgP4vVIuOLxj51J
qBCYmWV+PruJiku4/JXJrIcg+TsZxrjY2v+AjZyorginsBDhgMuRUWFdTO/u
J3aVFMnK22g7GhZHHyVJOYapVQzUdXL39CrA7m3vd6r9Pz5CbQsConZstKsl
BQb3NxiHzORXOU9l4xsTovrvXkBLz/VxjOPB2EvMhWXAwjpcEEkwHFIHPtXs
nGpcNCQZU6M6Tay0fH9twosV2ogijuG2eWaQMFxQgbjMEsPR7TLHIZBIr0jC
AygPMYOYmWzRthXyXFPkPXULl1fhpTQhRyfKZ+y3Kr8yFBVkypivs0p6oby3
szuhZzbBK3AfZj2lCBSGn3M+5HD82xLatnjuKYI21tGqg8OAuB2QTET+Qfw6
dNxatuhFfKjbb/9cqwdOT7+mLM1Iwk5lwf1ZtfDWavvAqvfwBR9OyHv/cmFO
Bp/LPFBaGCzRy9Gn8C7YKKPiPLOD+DDWfNQRmoBljYj7y8aEXMdT5vog1uRK
3v6Y8dXmkTthT6FzzL5qq3AnZEDScFjpU9URDS+KYoWBc7JNkBUinTg3PEjz
57JzIfskWeKMqJK54mKEJBlarMLKSnFjzo4QZ12FEdarFnMSWR40PCaHmrrl
KpLoAsnyCE2dFPo2V0GNdJS5ktaj+LgtQA/CxS4J85s+kWLFAaW6PI4baHWu
b1YZFte2xoT5Ie0U28s2GtglLoQAHfnFdHEwBLv5EDHp0l1tInLuRyFkvHj0
50DxMnA14EPFNvOzKAtOxE7nghQ26xyga067qGZiT7i3U44QIxCXj8AB8pmi
apPQunIb7/zeoGeCIr0gtLOuyKRI862JNeP6+mX+tPHb2M4UrwbVDLEYVLR3
SvxqBfEhxwCwp20qA15FPSwOK2WLhLTtSZz9AkVZ5yyxCKKZTSmUN29w/SVo
5OWHaYmoNHPOjELS5KPMZ+J1jg2zJTV8p9qiNYpnvbpmFBqHP0YdpF1/JSOI
9mldxA0YW1m71T+qn9t5F8W7MzKaJ3n1U5Ps6jAVEy8zdp9sPJMkluRIJfER
QBwWhiKPyLOkOFbouBzQW3DCrMaOmCvI

`pragma protect end_protected
