`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
i3/OCLYJO7ZFua3QbjmZQEze+bvgLsURbTg82VX5SGPTI4Xmf7O6Tq2MAu/NG3sB
KtLK/dBjWD0upgRw2yDSoo3Ffghw7HEEnaWgpuYHblCxEAqZQax47zgwtqLWxPAy
iuljn/H++qgasB0urqTxB8bGqGCSCt+rnpj0IA/UBvo=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10416), data_block
h0LNJiL7uD/X0FIM6TCH7EIrxuqSJrEiIUhMZ+W/ZTRrw0BJrh7feBnLGF9eXL7W
u75GWZASawTv1IlBAYwm/hxFwLMSaW5WUeeVxVlXMQr9viQxjr//YGDP84MKaY8Y
uCjRW/UG9Gg36M1Baza3m+rESTj4KRRzTICQSOiWe4yHdxeNtkiC72mt61BdEMWp
XbEyuvirfMLuZFvQk8dc84yL0w/73RqMZG8sznHQP+53LkHXK43Y7iJDSyi/s9lr
GSXCOSaPDujiluRxe1ONFmC1JyBUPi/b1eTvHsotJipHfuhmB5g9Si085Z14wnKE
ILUwFadPcqlObbtQ7+7NglBcsB010PibI5SYTk2zyTUDaOlIvMRLDbXQRdAPEQnZ
Y+hUU5t7cIZAeRlaplvB8bjQ9uY4OB3MPXEx//2dhKf8oErOC5Fd0Jb7R8hr349E
nrZkGTT7VCxq8kg7bn4xMm6Brp2ab/LTRQZOAP8V0He3eTfhycn6wa1M/q2VlEVI
jhvGet+Kp8oNN/aaK8lmI9euj6gMbsW0u//pY08N90QHyfmxGkyushg7lJUU+be8
KQFkeqjSTaRqs4AYmhpkUEL6+zkL4m8l3gnVKYAidf/vNPJyxYiwbmuhOYRkZhUS
7OuTNVjgOlAC2yqUx6oOWUK3WhxmjErWSq9dCxTO1bKvLQnAFcn98YWagW06TQe4
+nNMUO/ZNjFQd8RqNEq5AmNkJmH53R82VIhhUm3MkBgsC/PGHknPOnpl6SDOE0UO
xWrww6/t6fzTxUwLHa91LYrY73YBTpqhtebjHrU2h1IBt7Vbi5fNrFDCTVefZAQF
y8VgEyS8sihQAXiEsKgBa3QsQEHLPhonZW345DnzimjGNY3cjnzzRZUv/F8V2KPk
5Pv8JY8+7C4DCi0tXG5uNB53jVtBM9Iz0oCVRnIeCbIK1QDxK8sSVdUwp6cFF+gc
G3B2hYvsyQVhJCt+6Vu5z33ZgIMJeYqijdoW9YJ/ZwL+xSC8UZl16CVooQkq06q2
LYsDKJJEUBdBmc6DtMekuX0YmVx3v0EWymX6fwtfLOfvuf4xsI7YAP2IAdpPkQqF
jyn92jmpMli3h5xkNsfYNamOCAJaZ9Gnbwx0mawgqPHCaGji+Clxrb+yYnnMKSaE
Hg6Ql/lH3FmgDpqPx3dEjv40Rab7o7lpac30aZ8FOWMKEffjCXUxHrmoqPF0axai
iZY1riJOcz+7nIy5Vkc+dd+7CyHbmeXuUA3pZqAn1USPDFCCGEpiGMQ4z5/61JdM
waWN6K1Am4/fahXMtoThOr+Zdm6IpLxTaZvEP8hQC9uJvihlph6fNxE7yt4WMxqS
9d/+k8o8ExvVDvtHE8yNBwH1ZQ0HjqmnzqaJGqsue3HwZiW1iJ7gZO7O+1w57OIo
ee67W42czJI3TquD9NzHgL/dquPiXJORVJzN3CjdKRZn73KdsPNePV5nOJpET9QR
DMTpziga+L+bulwD1Gk0971fHlastW7zaxOSB7447C04z8ct0vO3w90z8jSkJfgj
BEBfuqoI+/H02soFdY0OmY+KBvMxeyDfmUzqIIIGBIgJSyjsiCgytApJcS1GOh07
lJRpEe8pdViJWYWcdUH1YVosMxDvdiAVplUchCFqtltcb25L2aZOuWEqWtvVx+0Z
jupennBFXC3uN4knls06ggCZDi748qU7BinfoKwJcGO9cLbuXziYuuZqeT8C2hw2
nRy50Ag2uVyokD8aggF8duxna/x5J6zrS7lv15F6xXGmjn/F8AEK2V34a4u1aJMP
nIzbeGpgscfxtQ6lqSCjogs4Z+vmd9bdIR053WDNKRHYBG285T+M1C02XyEVA2PW
BOg7WikjswyH3roKx/Bj+XP8aG4NUy4GDhsqmk3NmOHi7FyEpyj4H7xa47hLu8W1
MyeYGerwCSMbFK2DFDJOg4X6VEL5ia+B4kQgNO7eCs6B2BO+POXvjTYW0wG9tHng
BPfxKRWhf+EIHUcMfbQ43n3+kNxHZUj1jE4GLT7UXfAKso5qaWQl6Xff6jFte17Q
F19IA4k2rkXIhaxh8FfdnF1YVmAtRxSOXCR1RMZd3dfQY8wYpIIfsLVO8EornET3
s5Zcf47r7VBNxNFkQKf2iiPEsjMxe06B2Az0sl9BOfK3qOY2a3lyWp/qZ0wQw/E8
8ETr2Eo0gasvBNvRmuG952LaqOGUr9Lk1KH7/Y4r/zzEAyu6Ee8S0lI8KYtI9zsH
2gjuGwbPTKVpAnTDYUMJxBAirfO1eaz7duvUuypRCZ/ZsdTiH4nqsM5ioynEC4V2
bmfCy8rdGXz/5AHCFq5qpjwmDw4eNpc4dLhEidq8A1Tu7DQDDnijbHEP31dJ+YxI
L18sKcDaqfFZcaxO71BJ004pWSE2ljJiABrTgje1CUO8ga7eMsD/OsoGcfKV7NIv
go981ffh+2Fe5MZqhFDC+OfMytUm72ib/Kick9J3BHc4ffI4difDjD88GvWKrOeC
/IjZI/1d05H7wzjBLrI5am/KqD/9S5vloqDf0T4nmRCQtZ1lY2HbN8o722o32Zp0
5CpquT/Zw80Wo4bOwT3+UT3zQRi6m3WLk92RWNIcSl4Q/KWxDz/R9s4OZ/PbWcxx
kkdkt2rFr3rUc70Bh3WAv3aU7MmG1kg3f5qDN2kFD6U5VEQbX6gvTn8uSTExahtr
2cGAqv47XjYqlYMzQ7T08j+4C26b5c9NQXx3WF2PM0u3hAs4mUBBxHkg2drf11hw
WFgSSnQ7D2gc979wMVjG+hKn6tfnXMgrMM0gb+8KCPYkIcfgSXuyhx49iKwj7g5M
J034lbZTHeCjCkWzKqWH4NU9VdIwpEW5YThcca6OFmRmKfSeQCqjVBH0BTh2cXLE
cUGHb5pcbZfoDVuSjk6vQB/JffrO195ioLdGuIsGt82tTJh9zHvlSc6eo7yiE0Pe
OXhMPusYP6NZADx+69Zq18OwYxhAOOnnIbWbivUTTd4wah8rBQbzKTlKRH+N115K
b1MdRWJ3Hb8ezCmReFbCOZVLyuLHf6y49e45jM3IIuPvRNm8y1UwSvtm2llDdcfm
pvDZSlXGF3hB4dVYbb2YSzi9236lvY9935RTXEYR/rNjm+s8yUESIDyLfx9oqUB1
b3I3un/AJmDNFHV7uiRGYqqBCZHohROme1W1LxJcCflZIwTYsZ3N0QXrMk9+hRrL
D0TTOFUgY8SLBI+JaDuv199Ps52rq7BuCk+wQSpNVxQBFXKATIiKtwRm8xlLJcv3
0426uPQbUWxCm3Giq60pNRjCCXPWGGpy4JmSMfg20GjwFn6Z+VxCo3Z3MxPhPbf9
YpfJ8eDxZnewDOUFKavEMR0J2hiexoovfoeEh1TNsWBpG1H3FY2OWQCbrHO+343a
2fy8VWgqeJCutMT+0eCUa4WzaTizSMaa49onWrNabXdP+5KFlD4mvwtsjaWHq/mI
r4dA/J3FpF9LLPbD7mGpv/6h5/4M3fWgBcSlOrhEuIMrXOQ1yFfLvkHivfmqVXM8
wUEOE6Oh0WrHbIU95CygCA82+VAMzdJwYXR1PxRi9ELDtXrylNKkoCYZ4C46TJBV
UzleLVYCcBue53QeFGui4H1A0Al0zr4u5825DCNtVPm4WHcgub8RKYVh9L8kDC6q
XrzWGqn4ff0KqM0r9xzuGFb3Nu8N5IEMl51b3emzegIP0AEndk4coL9YMDfvQYTw
N7XXq2KZPBLJ0Qwz1uFs8l59k7hXYXigGHt9QxP9H9Xx19hWJHJD/jaDGNZpuqUS
OZpcgD5J371/ICBkrAkuIKTxmy//ucWRWBTiCHtC0D47TCMM0EzdyRpHUxZ9rMf4
RCLme9O/78bgOAU4l9BLiO6sXMZD1d8pYMBRB0WzmInXV3LnKhOso++OclNfL3/m
T7xqhE+m2XopyRHUFOBRHUF3qanVG9vmsJ+8d1iUX5knhPWJ6Zo+apf6Sd9PLLyA
g/tLHUbT9+neVmsYWlq8d4MGkuX84DPk9vF4B5gF9wXDR9AtRCPAdHemdC3hz0Gq
00VDbsnygNR4PLHtHyrpxJOBaLCmHe/md74ptcecH9YTSSJxrrHXRw6OicQsN2cs
gvJqyjZQKukDCJg8v+rQ7nnpi9OmFCQI1C6uHIopOC8koJMd057Yn+hQxgc1/J0k
dZql2BmICnZrEMWg2qFwlbmDjJuwl0xe1ApgE4RvobXgunqj9hkyuzIqkkBCAyYq
1UWRpeGUbgVeQ+ZlKAwnNiI99XLLQq2ZM30B74glV2YdlZEvW8YdJCSm/8dLbjhJ
SOk7fWWdQWC0qNcj1UoixhGIHSQ6gg+yrNxaFQtqUGDXMrd2qmBATTWJAzOdMIRG
2BSjz9fNbgnOe5oFc26ipAs4/UncfPETOddBLzB81HqCeZ+hMLB2Oc3cN0qutavt
i/A/4Vn/Vocaota9Z697bNQe0XakP226/spVEgoZ8pQMtAW0qscj+aHtDZ0q7Fot
mSNJ4b5CZ2cvabAjix9DOeU53FjENecQd5gR2OOOi7Jw+JwzifdtKfV57VA2ixJ8
kHMPIw8YUlkEFvuohlmFbjcqlxqL8YfDxG+PXgJWmUEdYrCBacdY6nwHy3gaHSbP
PO7cwIhg3+04o0/s4SX4yZlMPPw5DgDUE4bf8oZIilAJpw6jF9Fb+HQIZesWsetV
e3rH6o4BP8IkUhlDkXTauKo2USZ+mpqRJHNeoh/Rrkiyy3cO6++cVUgt4JrAVsYd
dvWE5ubYZWtXaHH9jri/fnDKwAIKp6/uLl7rVrS90IxK+LOr0FBEfy8lEkHOGJ4M
4ldCht9xd7zyiP9eEgvILbiex6mofBTSowgsPa5ujtYkLYr9rfBKc0OY7hmO5spr
7kfmmRdYWFWNnpqQnnp3bwDjBZxlOY4sICVpAVrn4Wopt377QuMQszP7ivkQD2A0
wUzvOnfvywSzEgvm4XSbROYn0vOWSP2/DwiVZOxKnN85piOnZk3RspBUFGE7Lenv
jeh4v99fc842jIUTebhve8Ptqgk/z8LULIpxCaQ+9hKxH/j1Sl0D8OhxTiGzXkGZ
b4kJgsuDt/shPPLhJamMVVklQNWAxBTKbzXpdJTcBvI9ugGmplNPJAI5wB/wsswl
dtRMi6+De7SaCyV1NGjNLKkRyCe8jyITmCTiUJM2sfA3BRFaXwRjNBzWUKkp697s
TkILh+k2robS6x7BHaki5fTCBLqOawIqaU34WM8XJJBCP5xnBZJ7gP0/KdgvXpwI
Smdc9YE3koAK9WKUbTPmMwizAviVccML/ES1t+bQiITq03YH5ZcfGykI3NneXuG1
xMqajr0e7+NEM4MN5SaqTlHTKmKtgSR543TPLfdkm2wGj6/OFoRAEDBY4CCdRe4S
tGhentLQUW9m7EqrMP7cM8kLKij7XYfulBgLU1DVorQhxRYAen66NzLIuzpeKQRR
PL/YTQyHP4zWGPeHgnEm9eqxfccMnq4Ni+9rSDe3opD56SLNb+MmBvTuerq4ZHJ6
m2bNS3FlSJrGapbizC+J35rVmU4eB0qy54Zwy2bk6FhMsQtX8HQtXaw7pnGQmn+7
tef1MqVoWcbYRl9h+8CUkYXdZ7lx29F2mWVEFQH45dI+JK74dtQfxrCEeJ01cudd
7DWwNhcopBLFkwdygOi+zCfVvvqVXYyYhMfTxvLPXBNgi7G9TyhyJb/3XjyFlHWE
xXZDakz76SYy7+kS7QKf5MyyvxdEMaHut/VteszKSNvSKfly30uRHsiicWgeYW9D
ukvMd9uXfhqE5+h6t7giDVyYBPYziH0PYnkjWC/1WdF4yZoaGQnCowLb9QvtCFZm
4jYd2pI26K4BRoMvT9/bnsWr6rFlb0tIS35hcDILKZ57JjBFahsap9MBOSjGECI/
geAjxbK5d440eydOHnMNDuqnX0SF9hGgnVHMJjtM3dIi7KGYCTDk4+ohdUay4ML7
nzpZHrxNAgYiOylc+s4Wzvq4Q529i/ECr5T9qyouZ/YtnAs21Jt9mNuXb4rxzNJH
/X6Kbns74BcUWaeEsYbT9bFzKLSf6+OBdGD7yrWYBxzzP/76ru7q83VuzDwNxcCh
SVMKbgfv9Bx6PVB9RqtrDzS5xfiCmHJAddxpkZ8N2+OSVaZuaSCxQW0jXu7eVYk7
i8r06GiQLfPtLgA75IHmjlb1aQ56pNRsg0kXYUodwW4aolk696+n0XIXofsPJPZ5
XtpP1HD35cfN3PAan3q/9SQTxhc7ZGxmOJ7KZXcNCqX9Z4zEYkSvT/+94zxpNYrf
b7AdfuLw0uB620dL8N9du7aoxv0qaYLiNEyvCBgarLFbdLR4ohZAddJGWcWUTgOQ
WSP0obj/v+b8zaYyZc8ky5vQ3MpXaKqOMMQg2Np/B1NTEt6o9XTFRB9in6N8TBkX
UyLcZoLnSsoN3PtxRzoQbyMemTRoaAXeN8zZWyELEvnZuQ5W1zI3O2Vm/UR6PpOJ
u8l0vxExHcLlUR/EAA6UsfltsoNSZtWWxRIvoR03jw4mHeWEwUN2HQpv3j1LcmVe
WHkhNb6x5NO8HNgMR6AphZuPHs4C5LNKNqjcZlI1Ej+zTIYXaibHG8XJOP/DlhxE
cyfRFiayoRM64tX7VbdS3llqHHfA/7gZyYisEvqmc7cU8c1IDeqBUEnImAzV/+AE
cux367Oy55KDlrgwC/AZ/3LKsp+z24B4r6I6FRAGwGEO3KXkZs6L4+/RIF7ybm8u
BUqZhw1IQibsCBaGIEf5u757DfZg4y8yotgKiErjlG3soFKzIC6E2HGt/m5HC9hE
fCoy9OO4eyAYChPMux3Jmu5o3n0OG+KE+ej6ss742HQa7ZOthwTrDaTKd+c+YNGA
sEBp+e1SpTP8XmA9/4Cv7xjoiOQj2G4xcvRZswkmlwVUNxRDmQyW47TFAthAU+x2
RrHMvsXlxkH2KCdiKZR9DyctxiuGJVVIaQ2K70Q6jDkPe4u9ydV0+MBRHDUmjZeT
tt4bNMLsK6SpY1xuqIXG4og0+041IAeSa3ulQ5VWXyLA1BcTXGlLm4IpZRaegd7o
D0yFWDsMHGta759reCQ9ckW3jyhQWsiXeV/edurPXtLFFVtlL7sCdYEmxzhrXObn
z63y6qof8u0EQZOT+ZHKzz1zMcbShzhGavxIra5ODdOBW/2t/EdmA3HMGp/Gx5Kl
nV09rBByRLonhpDyUWSRKlRbNVFT7HGVL2icQK2yc9Eg50EZtK+NE56aOkRtZSWd
pkVtwEXFemRovE1EpGSY6fHR7hmgwFjdE4ctgTZWOLnqwocBqfrU12IzFTz+8AEh
rYl+oXZDRuq3HdxV/u8ezopjUdnnvmEKRlFrN5IiUHk5K3PY6sENGwUiutHdWhDu
JIo5NIjG4nKI3yY9BI68gHp1AUx634/0C/NpNMoCcRBwQq6P5XGSV2fXLA2Le7eI
tOu2Ivi3JWpXR4QNkwHycrm6LA4DRLxzZ06INVpoF6YTZouDhgVKwHFHXW8KUOTW
SpBvnqBwgMOqhKCPyvLwkVp8CDi4wgcsTRgZkKgq7DlcJWRfSadysZ22G1SpVCss
keBNPfmDbGXdplOMJjsLNdQkTHS8ivrZ6wcUQZbehE9ch7bXP275a3vurjQF3jv2
IWcHq7CPo6cxahuVOErafFDdOMSqZnPUjGi/VhOZZtAcotiCUkXizALZ6+2Qdb6m
gBfUKoPcgaFn9i90uix3CcGIsHGL9ysXSJAk4fIYVnv2HSPg9Ut+Sa/omXGYIUzJ
zDePv/AL3kJOdRFKQTwDEB/obxn26dUhojy46bD7OyM8m61E+HW635kdpeEW0kE4
Qy61cyBowhAFQ1EWMRJvPZRxwLoiFb5dauKwfb47xwLpQ/nEAMVxx9349Vhd/ZHL
BOSm5LnKPUtTCmFm6fxyWI79EZUR/br256g2Cjoo0qpqn2kRAe4SI+M2GdscHcug
eiqPcHSBnXjjAKM1AoyeEMOCzcKHKp8WNHpZaXEgBzcIa/WcEQM6a+kdODKI2NYH
fsUE+4SOmVNmPOH4HOjSVIBMOcD6fqf5dy5J8ZOBRfUWV27CKDyypvgtmuoaNi1v
uQubX9/CgY7aF0zNoqGqK6iVxSJTOCuB+FZIrGSECYnBulxIoLx0eyXs/X+/QkoQ
rCY3zZPJGX6HgPvLd+J1TOWeXH+EFXcFtkanzyIGI04AtFSePBlf/eflNSLZIdTX
/u3XIxOUIqWjO/Oo6OnTpvd3Ivwmf0KLtjJ6K53OwYtsVBOM5SuGVCgpzrn4leiz
ycmQ6n1Bd8GJDXseiSxzLsIfw7TjsyAWidPjwy7EHn/KRvfhJZV80zY+ZRF+P2HY
RgZ2u76zmONe2NxDB5vU1iuOVQJL6jRklzjOmUvNB24RxF+zjbdSKp7G34uL9DF1
d4zN9yPolVV1/WXqF8qKQJxRfjJrQp3MMGOqJlSBpidHv5PDf4WnCJSfPVrbVeVy
YOuRu4EjXoNRX1AVgGx5ZyPOrIwb8j3WTI33xPgjBmZCg1ooN9JLMF918E8iUkf1
FhYSnuFBnjFnPRYKGrzwx4CP3PFVNRfqKtQTvMoSQwsy4gfl99SRc+z5fQJNlUD3
db/t1MJgKC0xdNabfQD7nhLIaeE4iiSKDlVqumDnosteu4nysv/yYUiBDhmyIKn5
r06iBENjwx2SdWrAD8EOjCWPDAgggTsy/ZiOPnhBtvsvH+kv+xEQs4uc5q7S8MAO
3K24/2VbMJ4CxlW3f9nM3iybrAwV4IrEU3LVlOi00UCzl0H6BWG5J4pCFsUBFGOT
vQfDi6adWZ8I9oIBaEvDfccL3Qh6gF9EdBfa0agabJkZ2AD4cXbWFkMG8sWlorX5
qQZBeUIYeHm3UsX0dhfEyD50E+BaF8f59xaV7FkgIjEY7NmRCkYBLb/kI+2+UZ4h
Mfrh/q/j50ge+z2twJM0NyErBWvSrro/DifFK0VhQ1r8/ldo30190xdTbmy9Xx2/
MVA2U2Kw9nQHFtRBGf4KJBU9xSeNVZAvVyw5qHLVI6asnxSudXGeuWUUblG+yg22
P+njNFqKi/xG/Io0yz2TnvXoNiVauaqCj46ad7ZBNGj7AdWxCJTfm5dEzRSuDQZ/
fevhLTw1nQhXOtISLfxX+loiUgws0XwuSV58jYHb7F3MMgEPZ3kp+aPGVB4XYJvA
U2HxnXaLr2GVroNFbe+wKKMxWTw0OMwqY/IYQaQ3l4MxC2+1QcRo3y/58+JkY5H4
QyqHBnSnYm3g/vKTGwoQn2bY9y4naRmrtcMzztEg3bB9xcop7EYLgB21D/FHtt7b
BjfW76/XfQ6VGpEbOMvvH8qcmP/MrHrKIBi2gh/yhyArVd6KQkpPqrH60aS28PtB
bqhtyqAc+9IBCXda9yL12i+zcr+dDMBrHlemVj7fsfhWacmDhOCuzxK2K1nELn6s
0OSOGJDA0p4y3wB1G5Zq7JQzGwGbpzleSRJBuw29av1oOVzPl8gaYFWi1wCkVPxd
J+izL6pLmuVnxFtG6RcarBgWRq/UkWM5yq3N28snutuy1/8bIwnncD/UiEpXZ9kI
VoxPv9xL2ufv3xUN+6HZp6U2QwkQtgREYiuzt6mYHz4fF/ZegdBrzR0dGk881Buz
+42taxGAOfw/V1AhJsqrECrXiAbzvLYOVKuydoaZjEmkVpDDf+MRRuRCrnw5MhhJ
SIer0eQTGK1TModdqdabgzcCdIScJEGj998BvQqHze5UuG4a2bU7ipUHp6rwEUV2
c+gi+peXeq9wtrb6A3O0T2k5RX3dKR8MVJWOEUeuBw+16x3OxOFcayc8MItvpA4N
KH09MhB2ko9S+yOZqoIkz9sBiykLFMy3qQGDXzwihorUN8/461TxQMVUfYx/2j/6
z9Zl5u2EZ0smDtHyvmCiVsB0DqSsoUcu0g3zBcv3oejYwsqEnpIwbpeXFklNdJ2N
HIkJXUpGtjx+oBhT/yDS4RlIxX1pMcPsY1g+81iQAfd/U/OcsCqa6g2hJqxniGsq
xLTDe4OBZjSlIcp15GWz6ZDOzDzmlg6rsZsz4u6G3Drn9yr8N09qQKkm4882G7Xx
lruHInoL3FPTog8Rmp9L0w0ymZSwJ0kho+7HBQJMqjUR9ly4jH0lYsuVjGJ2HZCT
74iFziDJ/1GcYtd6ED9jDgx8kIWo3Ltn6OEr/MkJQdN35Yl/44mQ4KthhpNLhEWX
em9JilKjiIl4d6ePARrmzfsWyE6cGKvcL2xWmTbywtKXEUsGSI44Q9vyuRqKwiIt
ZtcG4CZFoL9w0w8mbjP45Nsk08RneXJclYQgxdfN8+A09k4P8LwZfysziOl64Mja
xBI+NcJxfoeeRRFjHJUZ82MQRfkatpZPJSXu9Snb08FR1zd2741YgYzee4eLaquC
RitdJptWK3hrROgZbmL4EbueNrN99ZHGbZzvrerW4briUMS7Cvo3+tvIo/+pvlQH
MytrFkyc7i1iwCRJTAlzPy7TH2lSoG2HuU6Og09UCbFSukjMSFrVvZJqJHa/AcHV
V3dmd9zezqrRVxCpHkoBJE2oEj3PHlm+dIOxmBoO1gvbdejccy9xRAeqEalDedhT
cwMYZdQlRxp8495QF2BTSeGrKpZlD/YF8aO8lrcOmC6SiDCmFF1E0KtphUkj5oT0
XrIlKEIfpQBFWY8DJBrMbKHNwQbK7cIHL937b6ziE1ggPf1SvFEibvhT31qLXp/5
sGQ+kiy8Rvhz52Hf7YmTVVy8apPzS+YYlATZF0fg40Xf8r4x5yUqz4/RBVzJGqff
ypWNQTRGH2Q9rP1+qnVJZ0aVe0JVRSewd4RICjV8mhIY9HjwahjLiAWryPjL5bvM
7dtr885Ym0gFtpzMv0dEZSX3Aq1sK9FHI2y/5j/jcSywjWdiQhvkI3nSk7uZ89Sa
jUdTpTD2VI4zOaUAOXZSoAwT2A2g+RIdRCmVOwg9J5rZGH7yAnelkA/4fLFTiWyt
JvdG6BYthv1PjXLmvhVB5haPzZ/YeAcYWSkBgeXpNI+zHzdF3POlWEJGP72B7R+s
APgH3IWtwAwz2FBrV14XE6LdmDMEUH5j8pnsSDPBZOD3KhXMXXZ0pEGXWSQmckOR
JQT9yDgOArh1QCT7594qK5beAdRLp15hHfLzJFo0JYuuZZBZ9mookavOR2TIknJJ
eAZoujUZyIq9c4SQwmUPfQj4cCqLolI+E1irQUKufAmxO2ZIx393BKCF41K2d4Da
Wk81TpUKjpiFUu6omuCn1G28T6tZwqDKDkH4RCUODkjngpwg8eeICjW82HeJoKsx
t5o7hSaZaLMb6HlkOA/nfuOFdSnjBWKi6gT9rhYK7DdFS2xvNjtnsF8gemd2LeOz
EM4VsZDUZIMEj0vKeoH+DFFsKhw8ksrCOJgLWScV6SeqorQ9wFcYRFQ0x6natPn/
IRLDxEIvG/8Xs2kWkSuSPLCLLxxWlRNYWFvYHX8F3mDGk0fujiOZbAmajtDNqZ6v
LfJGb/ZotYVIu7cJnedZt3c/vZMMDiZdmOjSAYuPWFymwPEBUnx0zi0rt8WPfl5j
4TUS243hMx9kWU3LxB00w6NzvDgBwsx8cRapNPma2q76cGh+xqGkxx/6aqbZNDQ5
f9wv2ABrIkeOC3KIlN3fNY8+RHGrQavXR3Pz9n0SGNSQ8ztapRRN4H6AFrbucu8Z
HUHXcb/Nca51vmwGC9k5sIbhTZxgWgd2xD9Rw3XoWRtnpsSBNqlpBMKkS+ZzCO3Q
IrfQ4QTQu/0MkEQ+bVP6rm4Lbsk0mQ72SBZQ3V79BFR0s7YXyxWWSqlk/2bD3X4e
B2SNHDOAAKKlnuQvLX8RjatKNHlWNcOUvtuvSyTakCZo4ti4CI6mH4nMob82kxCP
dJbbsffY7/+rra1A5TxnNm6O4A+k3eFHN4y2DXBmywL8rjAxAE44L9xy0eVVBIC1
ugKfz6nIkH9rrUwAKeBuvlCAyiZjyRSp6dJUPH+p0ZyuD9nvYz2oWDaS7UGLMf6y
32No3sHUiKOCPIM0ZbxPedakNq+kkKyhMCVSFFheYDlQqSjm3wK9JE99iHqsZZOR
sEhzoSeKNzJCCA7WYAB8D+kn7MxpOjuTQ4o+Qdq1b72LEF8FiAupf618i+YFtxeo
YyGf13BmKhWzoXPmPFMmfseqTTIXJtiIGjpthapRrHd1PoLSuHqAu2ZFBoemutGG
WYvUpIrXU5xTbxWs6I2maYNgNA0UJF1FR4oBjbG7sRSEjix0f2cFDRXJT4ufNWeH
FwDiSkGPJKRyxZM6gVWugA5y5Avhqt/EugjrQxf7rU93wdRcCP6waR/jIucTxfUa
Nf3aHvVJnT0w5n1xpEUtzp+CG6hNyuzz3KrZgqMVof7zHg/v1cPTuXmPLfzhwVY+
Z405p8OjBLf6s1NdEMkvfrQGgDBggfM1COlXOwsz1PQsLk8LKNzjpecNLNCMX30B
xVdN5koWGVynKOoyNZIHkeysrewMlLKhOC1VmSXT9rIIR79226bmOgJmL4Wy+klc
xfnW6mEV0NzXlfxtQWczLjZwXLmXg+415uIsSJxRgCHw8Y3Y3QOU7L03mPvAdQiG
Kzo5KJxvqhkK6HIQngnZhTwdvC/E8O5KZnnW7JccGGSBqJuY/8MJlzgpH7eMKFso
0Xa5kD55iZ7BfdjRDU6+DIh8BJKWFZ7RIDY8UpmlpUrwPiQ7Wths0vfMMEN2IT7Q
b7bbcDZ134rAy5uKETIMnFJEwBYEpvaK1PntBF+gRIi7Rg3+YGVptDpQSB+TMKhP
/IW+PCtnPQ/FfWpJy58JqJ0PhXnHjW6nHukWk0tJX1tAPTICaDNk5turNeAPhvTT
A1srntPS/4Cb86M2gCEfKAhorOdx7DhTQS2BCQjxCDEjPn65+kNzYaLE//w2/vDG
hFB8RFZ03MMZjL2DaRmajs6Uv4LFLclWjCoEZE5KI7bHqIJPaeC+IeTEEWqX7RB2
+Q4TThDdOVJRFUpixi8K/YBXjpL9GmV9kDJJsXsEgNKKiZopKg0+3VwFsVdZzsnh
1Sqz9jnutdz1uAQEe78gd4gcBXdJ0iaTIj24Z11p4y38Awm7qe/i6pKiRPBs+pih
8ykyR0TBoG2DMJ7HriJJ2Fv7+rSQYu2MQwTkMGnuWBwgP6dWv79bU2vMo0ey5Ll6
vl8F4dHDv5KpNoGutD5BUu53zZJxOSupR3eGupEZeeVSFJKqB651Jal6Kp/hw+ww
cN56yhX950VpevBC7LjBGla34gHlEat91jw530U/zP2drSAFfzes5BwiEU76OUCw
l00B6mAa8R+w1zy36sk6BJwpa06DJwqRRD60y0iEYEhspXfOLLMW2/k06xMRxJRq
UTHjZO9ozbse1BvgbOVG6Z1RVTsa4K9D5A4Yp9lszMEIaJ+0YDLoVjAdnQ9pQz47
lAmEgfRVLRoi5zshoXIWs2FA7tz5SlYgNWZ0oDc2Z4KqAlOOICYuCWlUjFO5UkfR
OzLeWYGEft7ldkCjSKeWw4sPCsvXRBLOCSGIoLHvetOJEuTBQq08FY6urfigz9Lb
m8VPWeWp1EoBjCxEiIOtPhn4CEo+FaUlRElB9yX3LMraBh38JHtlXNup61AgoOwl
reE1fMhXvjct6IEOwd1XzDBeiPZNzY1flvjp3Zo0yfFbOhs5zANIGabb1irtlDIC
qUD4HVFRaQlFLjNPwDXekEg5OvuoO6K/C9EZpQzW+Eoza3Zs2+SkkYnlZAoBJlRh
JU3LrAdQ12FtJLFhluMbpfrwjch4rLmcY3USRn9oMX0SUJIcpmmsxFHrpEBmsYjz
8HsLfrr4lOY6RCYgSEenk2VlRf2v6OdahKLIwI1vK5vuoEvkh9zt5SexAvv1DLYl
5imUn5ipZwfg4YRJ1Jp1/KRDmFj3HTafWn2H/uxXZvlBG4ptrmCzaFRBTAfd1bTq
`pragma protect end_protected
