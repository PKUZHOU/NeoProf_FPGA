// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
0rJMsL1GL/8mLUQfgHSdbDuAahJFOo5CNQSgM6hAGqD4sPFSHGORUNAaJTblk8M8oLrzssFFfmve
RPnv/4ROjCB+I84Bx+HJxoXu1aOi2ZhkItqYS+3A7wZHatNiOi2ARM7ncvAdUdjaolQOv9XzYjbT
fewV+fAvXBfNgolK7Rnoam3l1ydGFWR+D0N1JclQmkTFhm3COQjw9GFeOArXQ+NahRiB70cAhbBV
cua1Zrw1bB+oVLEWZwwAj7MbAq3AZL4eIZWbjhSC1k1Qf0yMCnZQHg5OP+SPdr0BPPtWFYIEabGi
AjLjGcu5z5Fd6R7vKGK+/Pgs3iE1N9+BS9Y0LA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8544)
wmua67TdGsIGpiZmNWK0iTSNvc57cwEQEO3LcThsMDkJj7Xeo/laLyV/SIDSWBQiiWlC/MeNIYXr
4GTTQlGxElbFvuiMymrMAZFgr1R0nYqbaR6AjIpL2OF5ffAc/qXZlfRdRZFZlPoNWWANsYD9n11C
o845Q1BChiXeBtdLKz9RihDn4i5yZiIKLS0A2oUTzW1wcY3ebibGt99MRce6X6EXJk1awV4g98L4
w0EYZJv1LQ1uBCB602zOuws0uZHBgf1uKwjKwfRfynUlhLY62tUFWyRtmFfAd3T8THwj1icUPxEI
EUoC7W/seSDRPemUoUZ0mv2f5woMMeZqLFWwRignSHkbghVLXiV1qpwUN5cjy0/Ag/r1gxlUDoXQ
HQPSnfT4SFr721+xpc++nXnN6YmYuXNf8gmNu2yrhdYOG6uCLFUxwJxfn8NXw7+LQr2mC6XXLv/9
dc17izADejnAmyft/fOTSRCm0uwxzviUn4XAk6ybArnhxoIq2a10mGn8A2lQ6TKq1uOF0kLRM4A6
R6SfggvotV75bo3KF4Mevm/WgYOL/oN+1JNtj8dXpQOc/vJ4VD+EO96fpoC/pgjxHk6IAP13zhwj
9035hKeC+SzvPVIOw7M5cGwaxw3B/K39CrWwMBYuB0AFwG/5iAxAclxNXceXiGWcCzp2Qi9WgGgt
FggUtPtSlTVZBwYH/Y/VPkFK4OdJ1veEsNodhIwynGJ2CIbwN0Xu7Kb8bMNr4UR/r+CElUexCiov
X2X3zr8nOyowusWJ2wbwWMMAyY/woo2nfroNiCXTGM+ge7vFTlhX8CVqiDlWv/FBJHasjOWcg11Y
Lhniwp5ezkNN0oYmEooTmfMZWWHMg1zpbxNsVxH9IiNhJbrlFOv2/OlwgJ59pjhh1oPTa8h72hgH
Ix5ExxCgOS2mF4TtaOb6IFd80RhXLC+7uwBVlRCcexwezMB3ukMwUv8FisFIfGAgQvpGCOjz0Zl6
u0NT7PcnHcuZlmSvVXk2+c3Rzq6hyiuhzTfYwxZ94obgG7kBtR/Yk2fhaYDuyYJASJTOOw1VkhnI
zk+T9ntH0fLTOT1HO//HaHnvpQxDMSpLIUmRPyDlpgZrL/O7UBaOMSic32TVxR18xh85Njh3oyKD
krGIqWv1lGdiBLT+phh37hPXsggEXNrP1vv1mROIbLrMggcs3Lqqwe32ykpWJo7naYKaZGQbRj/a
B+WfxSm7jw9aIpko/ASLjaSo6c8JFkGwWCE8Z6C2U8eilL7ACwarUBhgMWoK6AzQQ03vPEhArnik
53isivggoDjkn1WaJVMiJuucOueq6J/RbYrkgAIR3ydFeUnvGjj7Pw3tQaV0gpaNAS+IiSKF9Bpw
dsYfYI5rLCl8BOh47fm4BhoHLD1UWawW7wIoJm3OkwWQOZMgZF5Tf/y0wGZaMLT052K9RXIGTO8f
LgBxs4WQfzKypOSAdyKvZ074NjmvvjgXb72CkifmptCOEdu7Ev1musFHf+9VMoTd7saWXVWQhhx5
SQdKZI5rcIv26SGgppQWp0jE61STexgjnGQ6WK7FVSzZ5tPo6IUXlOzoMxtCKiIXDE7OIVM8Eazy
sRFl7U6fw7SH6YmZB7qbYwIsC2T86bGecySN/5xZBok2HPFxUZg8WTeC4N+p9UBswYMLpP3jK9iM
XfMoqY4N0c3629nBX2rmMSBq2TfJKkhb9sD4vUXa+YySCTwaFpeQ8Q06lxv7o03A5hWaUvscjNtt
Ou7+Bxnm7HGlRAaxCovAHS7N/xDw2/GQpUkENQRDzg1P/YMB2YKVam5xWX0ZvaKuHcOf9fRx9L2h
nLXl/yBjHBli6NajNnW5dayuMlvcree4xtIypvhb7VbZlC5GbW/Wgwp1qavjvzVihmycNCiAFHwH
i+UbfVYofkKNRQsAqW37tqVJatH84Ry9HO4i9accmaBQhturMfgXPjLmvxYKJ0Z7hZMDjKXZOnuc
Wz1gl2gTbqzjqPO2Ryf5FqVfuMDJwWdE0Vi+hEALVup1R22YVCL+DBUkHreRCtBtBIJezeZfHpgq
9+tkKodvdGB+GdbLLQikBT01tQaYuwfGq+H6DX5yB3g3LICk3HioBex19DBapS/DrsgV18Q1GxU3
GyOzkqFGfv9KGU3t09ccaQO+CfymBQQZo5PS8DWm3jV15HtqYTkaQhLEDZ7OIEaPOn4diQUumCHE
TTWjIwPU/ts1nGUjyTb+ZOIn1d+4cs6cvguvzNFI0nWTOvSrWHkouMR2VvnuA+brvXfgefWH0wIR
pGjwQwdn9GgAe1VT2sxg9jAw6J+PUWPjbiBHCaCeYZXhT19xJel/pxsULJqzagr1e/76FAiPHAx6
lfQZrmiMXmorVd98OgSb9PzcWlhVC/qr9FCdajH02Ei4VIHpv6kQOvg2B+F7BlTmkcD3P5XF+t+D
4J1lMZks2LioWMotACs9J720VII5DzitS7Lt4RES740Wyb8/Cq3c0D68oHzX+iPGk0JFjciJ2j9G
KuNzvKjEVOL/pfyVhiRCdGyCdZDdLaZq7/i1ikHnpjd7/oWmIOCr6BwxSCTIcPBl2YGuinjzITZo
bAVgVMkNCLqx1VYEnzKGq/Ddcmcn/ZkCiSsLUVmf6O5JMAnZ1rM9IzEYfPFXIIxRDX9WuTF//4qa
8/FBosUdyQXPTklxjDbU/lNHHA8+qcPMBH8e5L1SPjZ4YnLqcqmG1ePQphdTICLmGhrpJC/JwjWr
bk8jdIw5e18ME68Fs0jlAmcCBQ6DUmVzxrdq74wu5hyyfv29yt2CYMinJ93tjw6oxf4iEXB4mwri
DxPbcj6lqH3yCSGC2tj77aSesTwKh+n+f+82Ll2B5B98bE4Wa6TBwlS/94pAe0PY7GMtJgDMd+dZ
iQRSVvb+lu2qBwa/pamxUc7r8f6T3ABXfSMBiIj6Kr/1fhy67bVD2GMhS4eYF7WaGdXy5HZMZ+jO
lr1/JPGWCYMk+cdOOmnkc4kAIs9AtcuuX/VaZs9yQ2AKbgRuu1VKd9cf4425gsQCrqg/4n1Dur07
07uj/eUCZu6/xkUsyCdJwZEpPEE9qEeaHFQNUGpcRJRE9k/xOLlrd1/2z6i6x5Ou9wOmdUWjvOOu
C1tZ4vwqQ2m1/obN53OZV4vidQy7f3EwFHJUWzphT61kxff/SMyAaSpb1wWHZA5qUYqmqfZd6dIf
9Bm7PUxTLT45cZI7xHIMkz7/xfPwyhyP4EOay+vsXsTA9tr97KDg/ojzvXw5drjklAqhYsb59v6J
89EQzSNi2Kk8OpNEmzqcQoKlTXJOQ71F9myj5AcuyXFB8q+A8dFaxcWA50X5fT9GjUT9w4Ej0YVv
IXh24wBB4n4sJlGI3+HJOmQoIR4jWontxxSVQHoUfgRqS3PLnTRYPke1Mg4ER/s2g/k4XDwoFOw9
uUKIa2BJPbY8rY9WVrnu5J9LMcZXva8MsomdorQiu25fxzxKLyouyonVEuiB/wXLFNEEIR1yBSqb
XIJcQC4dVTXcWoyoJVB1napZkfS1SijsobYXFQ0yREVeL+3Aj+ClcvlyIxRcmHZH+7WwV1FaiMj8
ybC3tHJhNQQ7StFxdza+Sp/LURBxLoFqvzm9ghi7Y4BLeG9JE3k6019fXVHecWc9YKappq9a5/EC
SqNBj8W2CTEQWVQODYcL+Ps337r24nydHzViZVex8nBn7sVX+b8lQ24N63+uyfUBnDQvTrqL1pHi
z5KpKUICd/cRYXrtQtuO77gLqdH/FDKeeVAB+VUVp6lYySyriEHxLwxbaAJ+5P66XHzzNf6iI/ZK
nVxRcFFjuMQjDT2bOIhWza9hYdqKk/DyUwUas9zrS4C1D6G7+qFpbchJZNoSfbM9inCvi3eGWruJ
k2VnmtZuSqKC25NiDFc9h7VBYenRSJNTOi1NutLSC7/4EfckVjDpp+rtLK4gTR68cEXx6GoPnWum
pNL7Jf4XkbYFa+lhM5qzN3PTiB+6M/p8X4xl8QrHQp9o/FgKE5mywNcydRatRE7W2O/AwGeinLC7
xoDCfLfP0PVki+aTcdjzJzcBzpX7JB/Tn2rFSpN0VaXZglJikwPRqVP14KB9z5cLiOmxln3XC6xX
KGA41Mihy4SgBuP8DHJ8Lwx/P7QmP5LUrSqTBOzr2dw7shy5vpek5PAMQio/VLf9DIyqbMCQlH8b
nzXg7aROlNFS1Sg/q3y8Lu+OiJ46XYaML1/8yeG6VLdvMwQkmKik/8q1MBwEGoKjNR7fROGW/ZDu
/eamNtV5vPc8WdK6s1U8FxMaBBYcTJKPjpnKajrXjWrBKaJT1ZF4UGNCFauQqwCGCyRokubOa5Ss
jURTowdb5EFFPp9K4sglpM/GFqjYE9p8AXsFy7Oi6JnVymO1e7pd2qUrUURh71J4yQky8Y8Yyvig
a/cS9eBL9Or7+iyq7i1vzsSFOJbhwdPao0f7zGfXWSCQ6KthHYilfRFqw4cEDucV8ueBBAjHedS6
QNj0n0DiOJ2bO75THLIMPDw1t9P28RJy6nSFHJjpNI+5CYTmomltW9UH+7H4SGW80CAppmxW+vyV
Tgbb2ifV0KLHGIL92sgZha4HtQ8q8+YU176c+SO0hxQx0dlspmZVsVsbRUOuYKf23k5JRmi8xwzw
MluA3oCyRDtWShWjsS3fU5t5sZ5ZG6iBlf91QhU9SCZiDKvsjjlr+o/MyG1QZnfzablnxOlwGJ0s
5JAVn2psPpQpdgyvGjqRi8iA0wdgqvfdaS329z4nNUY4JKjaok3rqRJNjBmkUjPYIWTR/zuQrpi9
kyDcMqM+EtyElILUu8DPiz7OYjIHnyp+MQCs8nX4pIOFf+T/5ag5aK3wLk851YOiSC6c7xuPJS8n
WuCn/LiETTgRr0JGC3ZnCtPv0oEqnJjnHStpdG0xgdjq95OJ9fZYamk3bsnXpf798Qo3jN0JtoCT
j2KAAJYh9Tgqkx1Os7o2R++vK/IxeE7De0+eJ/jKlY8VsKWqHPp9SflcXkp4trXOC3pAYsx5aSfs
LPGkO0COhNpo5HAdfhqX+02ja9mBHyZNS20+5KbZMMVmKUlEzdiDTK3GlxN2lENktnwc5lTandMc
p3z7rHQ9tvcSSkUDN5VEFChCTrouAosnOwfV51K7T682N2IbNajQVMSRWXMrVC2+lbLJdaNXl0h7
NtmyYucwdUDcK17SOKBM7ZDpouZPvVeg3gtyokWy0Vrm6AVzfflqfirq8FOQSsZHL7nhW47LdC7o
c8060RDNPogLiu4exUzcaLmxZS5G1jELYyDEV5KQ35mBWKyyDcQTqi5hj1h+69xIxPdYIQeDXKMQ
EV0RM5tYAISGWeo3mQ2b3oODRumIEYx5O6t0w31ANypP4gIlJCSCDw7o/KGtfrSVF7JMpSAL8BHh
KQ83QzbTTBbmQFgXku2+s1sW1secNzNbgaWBBC7ZQ69e/ZUfKz+eo1v3gS3nWqZMeF7F6yScwtyn
TwahgFAqla8tzfBu+BYuGyEk3d2vsIhnAwyo6MFrtZhbcqryE3B74bIBW4nFJrqyEudWqmfgStck
oXSTO9auTj2ZfOem+HgT+YtZkCL42PdhnJXeALnSEKf6gH2/KTGMMtmRpg8qgt4BcqqRgv4ISvML
MJr2518SntSYgDXcTXEQ0lawn+olIUpseK6/DHT2adNStCbgg8abH0VLGCnVZRr2a5ukFSTK9zWL
BgiegHHQyf0EZScHv8YoHG6IqCdgMJZKx1G8h/EfgK6Nww0CFN7ZqKVYBAUzNGo4VoUE5rOpFtU6
5k0ARugUtZLkgyKHJcvVz7s5TM1jLdyetFgW3xfXJeM34zy6+ze5PEzKvqIv+JnBP7c1kL72LqHk
ElqP5vHC+kc50SNzGhw95pZN8FTYS3kbaN+TlEG6UCZoA0ao6VnPntr8zfkuPCgOViWQpJKyenMp
/6nQU99rE+XyJ4KMBOKKsCxsVfR5dZUDEUtvvdC8lLREn2gtLmr2t2yD1npGwSGpm64vQD3EyV63
AFBcKAZy/hJpc4Kn3mOII/vyeYrYH72XB/Vookf0tt2zuR16vVqPb7bvjsWRbML0H3iYtIF2A+jI
flkBCYpTx+VZ0bSNef6OjCr6D61ae9py9smlG4LIpcfuxENXoZrihlsst5MqbCmIBm55sHllnygs
xuqSCHW4uXby2k8U1a4NiznwTFg51AAQnIdExhjyVP/ufZToSsWWKVON2wvvVDwtGiafjPicXM3M
4EHgjbaJ8FhskX4diphjevC/mf1DtJdLeySGnGsrlEWbG3RjjaNU2Uqpj8bUG69LJtT7LhW+2Ab3
aeGObfUc8T7rXjMoHAPH6QlSNlabQf9huFlNyPpkqsKUkOj2uUQxLrksmn0p1fCq/fHt1EqJ5os2
uJfW2bq7mvG2D84E/Q4Al4AUyjU8RU+MC+kzy5xyL1CWLvU1sFCM4A5zxpSOEYIhVY61kDQqXF9f
Uxv3AnUF8AMmFw7OFPTWTjMpDuNJ+t3G8UAtPgf4Ku9onIGvawzTaCQc1ayu07LlNtQMbQJi/na9
pcxn9IEYaLGv9w7CYUlU+6P0CY/sx9UpjRnyC2pySKe3xIIylZWkKxYKteo4xMoIJjY4RLjBkQ7i
sLGH8cS77WQMv32EJBgP+khXf+Sa5rUg4PyuSpcDObBUSwSsmWMm2/ggsFLb2dCno7+KOFZX0VrI
vSXWGs/2PZJ1Eaf+RzBBV4PJf4QdLxL8WrrUVmune6LS5eWH/NCbQig9ggmsU1S/QEpzA2CVTaM3
P0qSCQghf0nOJTJYsbVRpojYCcLlrbcM1l7QjTIoh1tJu/nPLItnFyeCcC9f/xec6HBSEP4t42v+
jR1xULeuBxN0QbhGEwAfxypBTsuIJ0DqfSAzmOFrsQYrTp/WJG5y3snYXXZ0lHZuVXtxYkEclrpO
EE1gfgdDBjamErmer3PlCkMgDedM8muP3d7UCN2SRjEXsrRSXxJyXV9uf5NSLJLSFHQWJV1hB1wk
M/oiZqfx9s8KvJD+IQt0uqBRVqEfQFPKX3Xmfyx2t10zfCz1QcB91s6dpXPlzh9iCFHW5wK0SywD
H/bDt2cSRD55N6a2mXk+obCqnerer3t3aWESGKkWuWxosWadWcvk17Nt3gaUOLyGU843YcdPllTN
+ZaSMezr8J39H9t8Tf7/IpyubPFnG6U0gqn5slTmPpOoiOoMF2xc5++qJDkac4dwOe/gya4yyon4
Ofrlwki8RiGY2S+fX67sOzorNSkQ20vJSkgoS8Fy74Hh/rqt7SH7lEW7l7R9lrA71BIBARbBJymU
lylEdWKDHmIz+HHYtu9K5hNFjeIfVJqvgzUJxU4jEMLarNMSVpqqkVpCShUH6RZrI8sFUOfwEFbn
n4RjFzUIvXheRIik9bcifgSwzIEnWMDez4WUEPBp2jwnSkj9WQyEIVeodPcbu3PR4aVXEl/PqOzf
hC5ZhlWiqRURtE0arJHWTobNC8IcSRupho3FrxI1ElATiB1aM6stxw9my1OWTpRPNXZeuLmcNDBz
K66ohNZ2oPRRH160dxw+cgab+JNocJtNZaGmxXBlUj/13UfJDaj4vdxKTAryXr48c7ZDFBx7NqdY
suz9rRvwcjkvG7vs9inIwzrQz2qR2VkEJEaK4ONREDRu7a5+a2ImUBzr2xTO3rBZrszqKWyfL0nH
HlKiRmCYKSkFW90tcF59RXZDszkbeOiLGmPcx6ridhEKePbh4RAH2Zpm5OQyYtNqTQLCy82UFr18
fg+Vzu8tK6tTp6ZjxNhd9Utx1leeoNYJvHtJlCi9PcHvHcMz6Sv85U6autp3gi22a5NTWOulVZAS
5ZpSvtxvk50q/tczqipoj21XPy34bhtj3xBlswZyrIGv7wuNoNWNhAYO9z7RIPjDDzRuI8jdsuZX
rVNs9NF0kp+nBgI+sqHQEIxSgk2riAozHELavY0d5vwQIjlnJmv6BERehirpXa3dTQ1l36/3Hs2h
e3fQlJFkil2KKecag95HZeX4ACNktUGyhOxmgnW7MBhuaLW0Grr2Z8df8G8UZZDoFb4hCTLhk7YB
7rTvTCwSRsy9Dij2kYzNA4owLqxTEF3KfniwK9maGxOsGMcnt7xPfrQ/O0ENULsjzFX7jZX1TB7t
KsArGOCyX0LdUDKXWcJ4RbQI1eVCsvqhQyckyeGoB9RndOaPAq3luthMqoE7UVN0XZflwDi7ZGDv
/dmLbvytHoFNu9VAc3gCa5ueCngI/Zw5M+x7B4ir8FKK0Rhd5MPX1DeTDwgKi6Qh10zwda51zc+6
LqpLS3Fj0boJjGKavfxZP9OuS/cV8calkPlnTxAJOUEkCx++YfFOijMxIf3RwsoEYBb45hZV6kh8
yvwrAmwTEkGzRjEmaukcbpf6nCzT/aMxxsGJWwbjHDXijPO6icwJWMPcG482hdKmTR35QjjTS8WY
icwRD7B0iRIpTm6QSIZ/s/zz6aJn8pIeJpWSCWa6SFILPQpbM8Z441DqrCTbhwHOxrwq25/d1dtU
n4zmddHt1FMhAoRzw/NUQ3tII9FghbVA2mm1FiTT2QaZUIbU9Yg8QpL0Z3xl5TfUkt46jr1uJXEk
Bt6LZHyZvYo6zCCJqewH+Qh45ACxTEQNIQrgDuob70Z45zlE2nrgWoKw6Yx6GVftfzchowZDtgXE
5JGVsHttA28PW99lGKgFfpyM/BdLwsWhNci9WP6FBpNrX+bilOETFw343kV6atU5QmRohZT7wC5o
V763vLzEjI+6tgGWIhGw0CJM53Fk55owl8OQx6vFmS8LdPqsU4w/mFa1tokOa4fLn21XfjKfbriY
Og3Zlvnu4Q1xR07cqtwLkN2GCD69Di8IsaQkpyXeGh0BrSGIfCFotYdYgX0oov/JLcVfqhY4nIWv
l3KGF4wOWYdxpDogNEWg+7uqcHZ0AD5e2jmsH9sZl4J4UO3BGlCGBV/x3ShNaWsUPPGH8/j1QAJr
7COUYU0Xa6xz8+4nBMqP9H4CNd16QILNC29ayVRfy4VkgHQS0DQQFKnZ4fOnb+nDeSzYNrjIDVoS
Ca9t8LnROPlWOICmrl8c+a85pMyGE69GJM1sHcy3oCCGObs8RcUft6aRGeMqiPoovFjs1u6nqEWt
gXAeqAaqqBEzgLsqSPyfxz+1wSY0Yn9FqHdn8nXh4fDi7NKR+itgXYmgW3fSNBTtEMj9R8YFtRIP
1571wpvp7WYAwWAug4b9XcQgbBE2b0dnFL6LXMctqWcKXQiR5lIlVEH8mTKnxrDoPc/S5HPLl2cE
GMwXe3fkBlIpIet0krycoxTN7oP3R7aZjJOipcwAoYE3T339XGRYRBOcAC333S4PEsT1Sg/As6bL
TLtWFcHErPIgP25Xf4xxLqYV4vi8hiupa+xOVl+INcLqKKVXp+6p3tldGG9LnyvakjxZtZ37yzX4
lHMHBZf9uIhV2jyGSqCOS0FrfkYj9Qtxfm7WZnHIsYXihIdsa9y3YUEGiouoDDb4aqjJ95iqViqf
CO9+FV4Rr7qTtlJRlAN36acVddHQGTQWpcll5UbDglE5le45Ud+04fC42U8JzTqfm71GGI2KEFCH
7n0hGkn8RMrOHBIXnSFwZ6FbWqhHh4lm4SNGv+8yQPKBHjhfR2INWb15djCafYjkmMEi4/8cV3AI
ukRbn8nc2nbg1zZdyU4oUVxDk6Q1GAE1J4IoWiSWoLq5Qrq5M0jy9SwQN4Z/VhQm1N1srek2BTC4
leFRYbQOTJeRddTEnr5RhM286QwdtcU5oXdK+TGRbV4QsQbwHTBS6/+Vte+UGa8OVqeQcijLS3f6
wCQKe7jA1gB3vf3opphnZKW5BY1ixJ6zFrdKI/ad2teUAOcgMlAhL43NKUuT7S4cQv9a+o4+MpHl
IMUFYUFUSaGGPihpa7GfZo78NuC7XdF1Xz01Ex1eI0f1Kn18X1V157H4yJuw3yk1lI3Ycsg9Oean
b6CTayz7yiQagIo9YznreDb/F13w4dmveIJyJnEjBwCogSxSsyTVP3nTOhNjjEv0gtwAS8FTgqwR
YMyMLMrTaLKF+9xCiWdNtmXTWLPIGeChfnBGArrl/hCsvQIp/G0M2Ru40VZEgH452sOd3uyKgAvo
zK4PN7UNEQ+qJUK/sEGIdGG322uot2/3y20wRHxNUT2Wslt5WWeLvPBAE4ycxiiR3iTbQBbqdL/R
F0MxSg3kKRHcgN5kbLkXUFugshYFozJAHxNW3CoYp85ZNLONuglYwYYV3ESGcbETXsXDhNQZUVMh
zJ1uYA5++5OKs9xGfKMZlH529yTlY1ns1BdmzPpo4Y5QHYn0Zzv6x6q2w/d2DeFIFHDhdqhJyq8M
Yo4F4LRLcNucPEgod4RkL7eAwveB/o4x8PwJIURCISWizgNOEep3LxkN/wimqET3xz+WysRbjGaT
w3FdHZYfQNklkDT++Zx2rRzg+Y29KJiCMpGRgsruePPWkAkPTimz2Gg7YngTjSynA3nzevGKU9cg
bvkFzdFuisZEN8Xj75CyHhnYPMI1VnoQW2M6twefMv2lTPV7VQfplQTREbaQVzYCrMof+jwN1+HP
POrC0joDV+WIlaSFZPOslfOrPpfq5Ho3O8ZP18qzyWhhTJUTAk12T0nD23KRDMp0ukH3vDMcZNBQ
eGTrx/0lzwMfOfWnuZdv/EVdhLOQ0jsuuKHCIfpycX4n0UB9xWl9XL/ZXbAKAR5yRiO7X9So1EhM
cFAzwk1GYvxToTOn+GARBRjsy8xAi6BFkaxUvOBXeX9lE+AdpeJ9l/4qgO+W5zzFJW8gnCcopfYI
+duXjqNvdFGb8gszZSVm1Dm/M7xiHcXPTNt0QOmOX7oreUEFHW/JCu4bm3SA1de6+ATceb7m4usJ
GSOymxrSQJX7PHbNokQZJVgUxLQk8L+tOOLVmg48Dwi8xrUWUGQV1bHJyiJSKS74Mlz+xqBWeTlO
19e7XPElsF/ApFoMCCqlXAM0p9DabErALAPTNQPDvwGqrxXbMz7/MM8ifflZO7Y7hgWRYdeErM00
/Y1WtArrVa5ciGpHWJc4qqJIGjfeGNnPD6shcTzpbMUiU556oxHcrWvjLQT93oGCO84106LEcyPL
IUQeKeW4/1cdYMHOS7GqaH5vImbR9plqH54La2NDKJoC8+uUejFfpR24Q7SiJqVj/WirEjG/IIKw
ZMqB9zIFS5TkzOvYU6Bc/H5cp7M+w5L40VBvYM1Gi/wa7CV77dE6RI1pbcyY2KLWsqKntJW5x+SM
9Fr8tSN+G9pfDAE8kYj/0gYPZTr/duqAhMqafvLxhaG65ZTB9V1R2WQqhrpBXdCG38Zwy7ZzFRBq
tpCMQneU7N+P6jiCmG5CUqsgPTWcCckAiEsflW7Jaiz1y6M57tMCA30qQ5k2zgg4PfoR
`pragma protect end_protected
