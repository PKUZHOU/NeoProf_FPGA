// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
yDrTYa3HHBH7w/Wq1krrkqvFC3nUFw0GujJ329bY45EfUwsyFZvUKZ2reODnvwozEbhYJ/NS5gyA
LoJrthMAJBeBI8plK5g3tpMWZFgo7+MG8u/tOI+4CDNqxa6hdLyfKlLDpHEoNUEwy6XL8CLu8wAD
8CCg+qS5/NCo/NkptT50Hvw/pczQ3LkemAnxzZcA7bAeoCLgaU863qwjJJAerzfiptjk+PZ5wU/C
xIqZPvNTR/OpfUxTeTrMukwSV4iG52hldJqoEWw5M/TxlwlTzUuPiWcRWxamrcB6Kzd83jJ85ytz
m//CWLTQYd+zkU2iv/QdtWZfgppKYSGT/wm77g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 99808)
8MhmgZ+4q2tGL4Cnks8rxyTf8ZuokfUdTen6InbRY0c85pPAoF34BqXwWE8QabmoH1XzfGs3HS+U
8mvWYab2zXP0oj8i1NXrH6Y43brAAHPzitDV9dFTlPPgpVq9R+jJ6YexBqkofIq+CoVbfMTHfQ7w
5ZVhLI4k3fhRXJBuvBg6yZpYHno4X89SJbOnKBhwwMYtM08ukOZHuf6YuL2tPtfeSiLlKsoSbBgC
6FR1jQAuX64bDoKipSWz8it+n1R796T4ud7e7YoWiz4W5GMoYXQTIFXlF1KmWTCOUY0CRq0B3/ol
Kc1+wgTfcxx/6lYFzGAKDqL9VKKp01msnWYyzwTYDN2U4eanWBV0LrnvG5LkDE19nn9tdgzB1u5s
uctMvlodU48cCdbQdO0HXuuscO9K9DdRRiq+KAq4nXx/dDuRdaxIyMWWXR0rhSr3JZQiILGINtVj
sEl5tlCfRKrnn4Iit8fUcyKgZL1rcnJ+D+nFOPtX7MkqmQdfTm/TF0WthZDrcrbdpP/XCJklNsSG
thmhD+WDEl2upMzGhWC0ZUdJ1E7ZaYihxPpMumrVcChaXizCZAVYLzEvzEY4omT7/GZrhKndA/hK
xLu8w6AyETMFOjT3Pj79AUz8vcyYU4a7lYT7+Q5tSFqarDJNhvKfwMxw8Iq9cfedwgM/Q/yavgix
SCmiwUasBH/2svuz8Tj2FOSw2Qj4OcS5ptIvg+gX8CR4JAZOdLdzo+3TpvQMRbPuXX+wQQvDqX65
/c+fEhQJGVGCwEpTL1QXaujsjAwEGZHfQ+nM6BFrxor77mQwlEzm4Duvs4wnjak5M8t625hVumV7
++/uyS/8MJnhOTZiE7EeUdx6VI0d9Ng32R1dBWUbrEfkwzrjASY4az8SHX8/ojc5WrnskSU2I8Jt
52JUWL/KnIlgrnQXCDOm49bebVYpxJ4x4CrgiV7wYAKQxUxsaaqoe04/qJaBZ5ZfVRFoRheBQ7YJ
zjSphW+cRNQnSGboNzaIIMnvmoEZGAKHkM+FqrbQZUKNpZNJqm1fwIrS4Rkb9roUWoFUIU8jClHH
flNwkI4yY+QjGhEu8n9bptcP95N4GIGwmO9WT1rMY5hRdqGqTzwKrtLcG26Vng2NoPpgcDy+VYSJ
qSauVXqT3kdIYEprhNAXduByCjS2EphDHAegim9eZzLNZjNLvHz59ybOGcMcmnsqRmrYGrVc8gzs
3J07wnnWu922z8q6Lf5pifbxR07yqyXnAO0KQ99ROKUI2y3TP7wlqeil3PN7MG46FQr+lyKr4LPG
4G6N+R9NLX3Nb0lUPdZxWMry6/FwI1MkYqzFFm1H6R91XaorENzT/GRy5Dj3I3XiNbpW1Q2jQF83
sGUV0iGyYYoApP5rwXWVGHbX9V1B3pHQ9JA2+DfVCce26Qbycn+7D9HwEWmf+Cu32aDAYXDqgt61
42HDCvWUlzUpi8ACt4fXyGk3IE9uCu6C+Y45UVkRxOGzswikXRCydG7+R7Bfw1V1jrwSKbPdgZkS
moLxYsLSLY3kXKPwaLVwbwNMhD3xDaYfDvoAbwmLe/8fbUG0CsezAW6Y3RtR4M8wAB0YTtFrylYf
f6Udvv50KgyeQ+AkgV10/RuTrX6BttLoaFKRyfrlp7tYP1cKTq5Zbhj3AxpiIlsXtRD+3DObFNux
qS5teWd05noYvuRJI6wL42/EXUYzbP7jS19ccnssBAFIDvhrRq4laxZNmRQc9rKsQhPa0gTYCcEH
XJUr0c7dnzf8lskoDONUjYJkMs2dOSKFRxmkUCm0RBTcdI2vEC56vuvmjIkZsIcuqdklF1FaLTir
QeUQSGgVCS4Ar1TkFAdUXZwQHFKGu0OjK/iD2X4bG2G969WWRfA5h3s8gK8DIre/jFLh6Lo9KNMH
kjdFEJvsSWBSVzXzN18tDQY269SLfSopOewuVF9ItQebi7wma95mDk64tQdoKrgYvJuP2kErgsMA
tH5DGU8Yxm606WNl1Qb3DNRQmNMqTe4leWdYQt2cXgi5x+v+QJBE/YkO27ZC1Lqw8Mkz3Zvi94d9
5UeMdDbCbcOy/+gu1lqoSn+VaCYG0A18UqlJcGraJT9fCo3ot4K43pmD9EDtNNU2IVc/qix7902q
ZUgSEj0lp4XfZuwHw18yJYi0GCCFJseOqrJzBnJB/nmn6Fq4/wG+auirntzxmnSL9Tl0InTbz673
F8u9xoi6hjvSdjBTSRZd5OqkavkJx4vASA59jnd1tsHIuPUrBvA5zmHWXzfXnK0GbLQoVLMdHAmJ
kHLIs3gBp539CGRF/Zj4yBTTj3Qm8lVNJ6PItpq3uZUlBBjjXutOQVGW5e2XHsYq173QXETYLAKX
thBoW+zm8Ns7+Iu5wllkI+GttoIJg2QsrFsKhUL4vPDGPQJRWHw8Ws38uUCPp+sRqQBSsCmjhGKP
UmZe1wmgZPU1OfzJ7dMvh6A1/ES8JXT5NnlLUmrpS2N+yv94uUCDJrIIRmWPy4CsLsYUmqlJxvO1
g2DwrLiop+a6J+LRnfqSEbYAwJdHRYeVgQGl6tsWvG1faH+XSWF14yrVbJyFvT3mJWP7MM69IalY
wCfrq0ckEuH6HS5iACYPYmWyCgKzyS+msYMFg8MpE2FzmXX20pgEohb8t+aHw6gWBwxmvOdJ7jOh
Le4v6K0IQ5TNiZZ9a8mp84E2byRu6TIr/xPUOtCiOGfZVP0UaJhk1oGhABpcHOupKORJb8v+UjrX
/e/fEEhkKWMYLKVGSc+uHSYR0PzlQe2QHKz++fuQlfrA1wAUWqC0NptNHIjhloWYiYF+XbMnBOlc
zaf0Q9ro/NfIkpWNdGSVgDwrPw//bPQlMTrtX9l7Q2XcCtvampig7aiGmYKvSQtRDJIfiNAw1xRC
oIdItBYmGQkHKhAD4THQ8c8cqWOe2Op2lZag/NWqq4vVZet9wGStT7BHDo72GTJjSYs6XPyEdNiS
6DxB3FTLfhSltFYFIcictdWMJAi5K1BBe3kONZYi/LqNLuYEUgZ6lc9EOQn60nhJOv0XXOqYaO8r
Q5WapiPosnYRLQIzu7PxdBFKmqoyGFzWK91QIG0YG27F27fLvYcJjmmOARSQpm3CFYsHo7W+zw7I
f3q+p5Rcab3vXk8F7XRiDHFMW/FZgUhaBYJoJHy0iQW2NzXi49S2WpWwRDUGQr4kZR/bwUrZRTJM
JwYB5/qE33ZoAVJdTIkj3NC4xoNyRMYWeIlEaiiVgURrarte/stoK2mr/yuJlJYkOYgqmMA8BDm8
qti6hu6FvAfN6e76zeDN3ycbGl4f9bp5ej8OyxbRtjU9RcwZIdNrJu2HhmqOodGoeaHu9loI7Ezd
bpx9nEeUwVoTucDk/jtJgShCasyuopJ3FHOJi04JK7zTMlYdBBngLhGYYOPimf4C1EyPtA2E0mNp
gRUL6chhQwfHvHHXMTom7CKnTMCHcAJ0/VrmQ0EeHpKDs95lI7bg+EhWIXxtDC/n5l2EO7CwZ5pN
ToVwlgs0r9/gb7uVOy3fOSLx5OD2mhr5L2nFbrK0rYh7TNVTfomdYHrsi0NJJoG5QA8gWATVsF48
lOEymaczWRe9E2AnsBMXhepPNwm0MVL2EKqKqh9FSUJJHxSWjT7BAT5lf5KFH+nW9ow5Qbl5Dmeh
iIZFH0m09MC+546ntvVIbO74jDgAwAXZqdsukiYIcEovJQEOk/6pfsmRPZ7mQOLL5ZpNZ1uTLhWJ
5OiEUzH2luE7WonkFu+2dcKDUkpo0txTRcyiCJcQHyEMohvQ95IkLpebkUdXpT+AjdPL+cFaOyvY
SU59R5vF/W5x4fwp+ZCXuHAjjPPj8pq0uz/onA91GYyYfSmNd4yGOV6uwNAjNcFFNkZZG603ENKq
4t8eZUI+ewr1jc82zGxLjmSc0Yf6M1VXGw3qEO21TcXlpl2B5r2Pe7QA2wpIXPt6mAo7q3Grc5MK
PF7ckO6zvtUlYIwsEeqKzMQhVnPBtUOK4RMs45TFuEzp83BKwR9RfcX9BR/LBsq7ZzQpLyXMKVdU
ur4R+Dlx3yqsct5tBlkhUfIrqqCFejKAv1p30jyXI4VfPRsIlNrfS9gttxrBcvJ6AzU53mMC3F59
t32p5poPWTPFrruPeRMhePqD9kv8qcNGtQzUSiySqmVGmtsLWAIT7tT+8HVBJpm4G5v9JbBygs9J
yUWvrFbJZrZ88ZkqyDB+ifNmahblE6J2ByFRvuIqXHK5WHQp6j6kGuKUxUjzjx4hLdOd/Af8X2x2
5418KC2MNjkLcqbu3ucd/ecX+7YrZ11Kg2QO641nnigDgVoAYFzWH7V8qeUFTwVMvz5qQH7JDOOI
K2usnBqsZBkPuagOl/FCY17v7ZCG699HWkwDSoyC13A/PKBT6YL+vWOWDlYH5cSsbVyTX/z2Xv0l
yqtqt7mf89CcXz8KMRgD8lPkR5fLAA8NdnCBJ7i3tura9gsD1KyoTM5gZcPQdjYIB7X01/c/SLVW
eXJf8YjsVgIQRjuqfkiSzdtVWMiAGbuKfraaSnJXu3g6anFchaalC1kSrb7sAqrfFLh2aHpVfKHO
0EOIloAi1ZyrXeqidy8kYYWnXANyZPGSEDIM1kFnY8BNTkTxBQR92p4ueeuFWqrFsEMcxAn9BzxG
0PNAaP/mVlTmnvcDjJD3sKCiUVkxNa/hwmtoSoKhIYt/JHExsJH6G49tOcnfr8CkOGaxQwDa5exn
gCDJSfcGI7w3UuSNFqiIC8Yv0/AP9aLaFpsbewfVdQOSAPiu/6zwJZDUn3jRa6Wjo5v1Teno0go1
SDzbJ1TkXSNZ479m8Kh93uOs53BuK3F+nH3obVaMTV5Bfzpl+zQhRsT2vGVl7iQo43QTBKzCPFhW
GBIylG6dAt1mGw2YWYbR0kkkCslqec45CRmDRTE1wHacavb2pFdpZKZQGYi7lZzO2/4rw9xt3JOM
eIh72hQVguGgwYTAG8GuxRKUWrkJWG3s0ZpfUXZGEJICIkqSFgmaOGCdhQbUQCATCMU9USpGSVq3
4hVRVDOjEDyEpR8RdnsiFeo9IRVy/auwi82DrOiq0EqwEdp4uPYSKgGxg/hj2J9MdAkkAHjGX4Rs
rHwMcY4LO+KUXNjNwSX+iIc3tlBCUfnYQ/izVdh1EpSjNq3EuVmXEiO7Wr8iBEyprr4Fu1i9RwPq
Mx3uvTtiYoAB+rKzaoNeIexA0BPHCmL0eE49hYdrcJvWFR99C0udEGfUDtgLbX2Ypghsag6diQfl
yP3160l4udoAtFYKfp4aHIghGGoiQ1OLVG2PvJgS99r5AH08ukXS0A4MuWOK6UhqnuuYaSvr/AYZ
yxLkxIqcrQnOPBapD4mz09Y3kgIYAxHhnsg7Oa5MGupGlAEZFeIOFi9EVfA3biZ88M0ij9mxSvQZ
hq50auDOqyGKdYslFnzIZ5K5ZgHhYqSVpMN3mwVOITAfezAXa1afLE+eFRRakwxX6RDEVveE4o7v
n4TAUxTPdeePrSExDMeQZGKrJN5I9eolUIKNvtCd7nWvcipGWohb+oKx/mHg4r/wB42vj6fYPijh
KyC2sGtxvLyGYCO2I1OOFP02nHmiWeQ82R8EjWmgnFPVw1XvggQWqnGlJRuo4OulmJhlzUFQnpAR
mKONTZKYR+4yQ7KPsHL6rdl8eyzOcEDHJAnO1mTTFx2lZQRheGgJHEFd4jvxvIORuwUay839j2xV
n1B8uFteLh3kDjNeQ3jsMgL3kYXa+EOTVEEDJZp8BMSz/dtpbJvnHs4BlfRw4P5F44Thr0dG3Y8x
WqGCch/Sm2Zbv7Xlj9WmFDd6AQQgJk1davLF0QwDHe+JEwSeMJ+xj4bTjobDI39yYkm2AUjpqJNL
qUjBbLE15U/4YMb6Se7PX73d6dWFcbooA/VhMInlbp4eNh6BL3GmlxKtOlOW7mO44nGjk+fB+VXA
mthietVy969ltfYRYBZ3KjNpTycfxhY4z603bY+HiFBGS66DVgXZSvkqRCoZUrYcjjiwiwnVoWOe
sMX5R8m2A4zClBS4RHo18emd6lHEnLAM7yIcr9NacvAJvZF1DMNdyQhotRfRYIvnToeYJy59Ere2
sAH1x7LV6V4phMjnGt2ASmf7ntwrn3En+5Ae6Y4biFZryIxLuRzOLdm8YGdWd4g8DA9g7rHuvf+0
ITShV/UablRHVWSrVYYxN0VZ8oqkcB/Wel6D9tA+ZUHcKld7R73Fr5qp7bR4p5BkJ0CH4/RZlx0D
ePbwRwC+Vpy2U+NFukmi+FLI6ZDC8i+4KGiNughfmU5bu49eRhkNetaqKyO/vCQseDjVEFFb2KXa
X/ryqStUzxn/Ufu5zDH0ccw4dIiy7nd8D70h/Nz/0YP5/xiAngRsGgk1+++8Ew/A101+1A0GSjU/
XjaxP5XGTZjt/BpaRkttBWqt3j43jJIZkJMdMCtCC68XFDYtS3K4ZcyODOTb4YOuRx2ywfS2GqIh
GdDW1A8L7T+DyeEEV2zdGWtWMeg9OIuBJD+9CCRWTKuHt25FxIQMER8RFcqmj2NWTJ2UGrxMkRbm
eyeT3GX0ZKct2W2SkjwJ9TaGBKgCN8OWwX2j1/keQgfn7hx2EC1JatlGb+hVahcjvXJ7Qko14BN+
6A4J5sLy1Vdd401bVOQ03gc3fWTy/iGmh+9uzlJmNHuPSR3gkxyKUp+pBAPX7XRjCxwvN1mvuZbw
3PXy53GYc0OVW6oNQOwJuLK87i+Gzg4ZGdDG9+xFnqz8cE+BiLhkkm4LOuL97se1p6zQa5UHcVvS
iFgkyDNFEOkekZPr+1Sl4MmOkO92LwfQ8m+O9cTU+F+4migHrPqNGgLYCBuaw8D9lvBpvMRlAbds
V2+4Z6gkAzFqAUJFxxOmu13RMt5JaHvfun0/Mi/lJ647CNEQ8TJwyQWbUBfmPH20oz5dk3jE9v9F
2Mdr3TOl50HyHRm4gPSRvACYHzG9fWYrjD74vyr+v/FFqusqapRDSG0czXxKG1KWO6Qxi+JMNwrW
KPy9mEvz8NEU6pX0g+RJZaalYfRg7DeDtRESENz82HiOx8rKv6UkQmG51ziH3GreIqqU81mWDjt7
mL94F1MpUehCrz2MDprFP/s5UztbBclafRwFWhkfz9UrudvUqWkjx6NIk0TWsR2VD+/JbIqkBPDt
bqYCglRFA483y581nJzF1feZ94oKapZHehLVqZn+yys13ZcSUpIO0TUkoa44OHKkuCwY9U7KRGyV
hah06vfmuUSycGJe9dMhf797qQvdJwofSxNA/a4YhHbANYfhtGKarGjP6g6V4HbKO8mdU0d1jGGb
tWNKygxq69rWTOnANZ62tPOU6JSZf45xF9OMOoLKQP9Y2XmkaUky6nDH5eTQgfrIgLGo/nt32KfP
QRzsFnt61vKXGM/O3N7AZ9VA2ON0IZR58wWWT9kouu+vkT7Bqh+nieNXfE0/pIJe0KOjHAkbuWvO
wbxJYA+si+zRXy/9u+SBNMgKS45L+l/7WABk8h3ZSApCDI25LHiunRySlhK2D7iy4TdLZDC6Fyaz
RIkShe0ONCMO+35FRprwb1qV1r8u+2XceC/ZFHoX4McCnKyRimJm9VQI/2G3ima+qTFJflh0Xwzu
VMeyHsx7tjX9ceyitKJHRUexxou3nJFNU9jbL5S3vikZIYhnXT9GI5tfi4azv2d1wbaMI9PDysxE
0V6MdGHcl+kJi94OiUkslENIEgj4G5OdbnfyAyhYRjfFQh7UFSKsmY3y+snl6QDz/X5mtATpC1d4
QC1wWmhzm5S5Oycaq8kkXACjplKibgzdp7+Q5vv0gMrbbz6tmi9zkU5EbC2sNtYgNwyqcbJNf80/
819HFoYl2aJ+BnWDRpE4cq0Hj2fvofT7FjWS893o64wgnRQdsZR9PlLNavvYtDnnQGA2Feh8ajT1
f1sBr6aE+TFo/+305ffrRmTw1Etyx9TubmSw46Miavra1JltvLmKaRB3J0lAZOyzyfkLwtVORSTw
3SEPNsKUKFaen9mrzyuSqCZuX+F3BP2T8gvGP4rXzXopCb1CMDt+GfS68TCrtsc1QpWAZxquAuYa
vbBi4m7jo4BLYDgMMyEM4JtkCVrQoKPNLrWRoaiPXRktLcCsuAhO8JcNz5NETBlX8/4Xp/OA+LPv
SlPFbgXLQUigAr98k4fc/w7GBQxc6aRiR693osulYUb+p9OCm2jVjV7weBFwr5lPCIqyy4Q7NnuO
seyMXDmT+ONxyNbaHnkHRubeYJIIb/YaO7bSSzWPFx4vZ2+kVcVZ6dDcdlfYYexnkYFLGGepmzfd
/1VTQy9KwaQnR0zF8SVFpxHwJuJZZkMQkvXVq1B7CJiaIixblOkIkxeuhQxlrCDn4gh5FEb3UBl0
/zhEcY+yAS3QmoNaxYlMLXZAmKUjKE/6GQtZ65GDvATY9bkoiTxovkRNLX0vdsKWgfzDQOsQZ2SR
cPsuDmL8/fUzMGm22OSfj2ywPcqtfESkH/V5GNVdR0F4f5BkLHLNRIlQOipW6oS8TCtlK/FbRfjH
zcXuH8qb73+JuTSkFSIc5/lVRLvFPYdCkQQTg2c+HJqr3/5NvU7IPwjDja44Z1ByIg0XiK+3Ckz1
fYIS1KCTrSuP27mtdoepe3xEd8SoqK8vCIlZmY4qH8toDibl0sPjg5OZ49LZdbhnVI0lXQC6e7At
jnIL0M0ak+rb8cvgGKZacPM0dMEC1Mn3/VRPPQjZR142N8bWcmLUp37tDKbF4/Y4DRNZaLrAxhzR
+Xwr/0pPI2uZfm7dpbo4q7pqWoIvBDc+SFPUlNn7MFObrtKvZpgwnBkzUNI0t35aULt6GoUWbwCX
mG4A51EoWzsUx47wjwG/z/tOOrf6ypoEQZItciKY4wyvI1qQYUjd1ITwHFi/ocKcf8SrfGbB6K8t
MdoFNo47XROgOHmgkMlIaz/lnG4l6ji5VXUIENz2aFXqcZ+q6X+MhpfIluJGrzoimNEG3NwCMjEs
3ST3l84lts8YZyqW+r2mbYKJVcVEg+SaAkpWJnip8HgA505y+af6L+BmOaIjvqgZNrXLR8Kmti7z
SQ6HJoIU44j5Zi8JBLq5PYVJZ42Yn2xy1dOWE/Q7yUwzPhyk+Qjqi897drJqP9e1NogbVVvE7kkC
30K22QWUPVWS/TSt9xaNwBKFWYlZPg7/8+hkIL2/RRlM0S950r3kSUrXsIDoShxcX5rVfNq39uO/
d9zoUHQiYgrWZiiyHoyqzjGivj+3gdbrnStq2akp3wSJ26+Mtxgb9oyL8VZEQ0ZMo3dK1vt3s4CO
8N+G+O5WJdHGwxCrQOGsDda2Y+WrsyPthTfzP4r6F1Ma6PrVLeFcNmhVAUMJSO2yJDFr2qlA6mgW
TNwAc0LNF3E8Ws0yzQhBVG2Plw/nHHmpNsfz2m3c0FeMeNVkOrL/qF9Q6g+MJC3nts7Ae64m6u77
3s4Q/Y0zvo5AdMxRna7ukad/ynAcuQhkb97rNpXSEEyWptGifPlqJg6f1qFbiJgkpDGGYd8SGkDe
FdlgABY0bEIOXfsnTFfL6VMR4cCBJsUGKJk5/8E+hr2alGIIkwilRbC9G3+ml6GTZSXCeEIYCp3Z
t+7b52HKP+9sZwGH2/6zteLEufxXLFkvmmqc33nm/9+m6iEclZ2PSg1TaHfdKSqwZhaeqUtYnr0F
Nyd62+gEDHyRT3ejX2+8gDFSdWOiiSllXoBw18qPmuvB4xxLOV6xSECWTQKT9ECsNjCVPL6H41+y
PeNDN58hvOuP/zb313TXvN+6C3o057Jcfz+ICaP5UgYzgAGeUWt5Ol0LI8ncnVeNauBlN8H17XdZ
yA15iDdHP7Wg6Oa+3Q19z+63hXnkms/rf29UPuOHIXsMT7e4Iv4C+RI8DIMa4+qRWppgkqfLkEj4
qBjN2F8dG/H9TaEWrRaDsgnl7Bs7a6ITYGOJUV9yvHf9Koh46BPbD8ljn6BjeEM3F5INCRhlEAw3
JskGRvRN9YoZ8VIXw4xtFTz3eihJO9PQN+ia/r0k/Tn4LLwxs25uzJNsjyYW/D1PGVzGHraSkYyZ
hpB7zNgGIstWBxRq8qEAFbgCaEmO4L9urozcMjqlo2qaartILvd+rz4AB7f8sbY9ZH05ak2CfvRW
YHIyEJ/UNPSYdHTzvUySpv81xxS2VP9grWUOGkBEdthgwh/aggG+ASCgyVrsGlbqOb7DXouhtuwc
vWo+riMFNYHJ7Xuu+XUP0uILXKKNHCyrZ8oH7ZYTqmD60heslgYVdSKEse1I7dVJR7wYg3Yjzrnh
MfQhb37oQPEshbvnl27E9vKYsKLHLEoB1/+fSYoZO0wPVjdOcHlSDfB+1s6g/5NORtQU+B9CKEZm
KQoXizQCLT1/LG3HqO8IeWM4JJwUm/k0j51jTEckhUaLFCFqgvpqtkuYUvUiYgA4QkYiJEvgGS5J
neOPMGcioh2eU86BW7UW8P0oNlVWe9zxozI/qZlCWJTu7mS83sUy3CPLWPt9uJ+6aYBgU0vV9F87
4Mf8jjNv1pM65nZnzBReqfYmJAs6CWidljJa2waCscI023DgytfJP/gxPfBmkkgu1NuIy2W9v/zt
VwhzgAQ/tqA9sO03OwCu60AQ4oCNVNUfTFy5vYiFznsVuiiwS9U/2nFZplxdCe42+GvfNCckOfea
L81/EQGuYBK+u7vycvfhOd/RWEm9+AWTdW7c1SXRfsF4d0HkfsBQfDn0xw1j3lu1g6bVcGepW4sG
EQU0/ZrWPMugVrg1tbe8axU2ScjL0RB3XS2oKhZMt2uOY8NzdHjih27DRBhegWJxEVy09SJCRR/X
rrU6w2mnYQWu6P5T+ddWTyk1wSYHLzCaZodhCKDDZxiFyzLRJNbyFARethXa3l7DDRtHinsLH2+u
EK2AjKbsZddVUUwJlA3YcfG/zJyEdnjyavgXh5oMeDnI9KXPRMNidEVVvNvihr3ltC7+/WGJIIlj
UStBbI9sDyIWNxZdjVCMbZDsZoodJRnitoChgDUT1qQ/SbhruS48pPRNxYEmJQ1E0+BhMF5Qncrc
LM2EjvEmyFcxZnddX5/M0rUDtUfp0w9kY3yh+Y5zwkWK0iC+xkzdm94VhtzbzOHilinEl7POM+Vv
alOpbBG5YSBiYOtjeCrMEfNjk6BmcPtBT6LD0CjWFaeWE/Kk/5TgCGLIx1V4UauGpq4FFuHHOJZ6
aZu2xSMMZj49zZs8ujBCcMRDhjr4Hxatd60LumNA88zVUCpiy0JNpLuuyp2eQY3molqLdnQ4J5Lw
/P2gnhkOCdRsjANQMb6sCDltlCjqFBNZmXRTzR2l8RoDrb+UA3Eqx4FXyATV+UBSWUCgOy3CGd9v
7lBkgGXTDB4PMWiLqBHcpnWAWf7GDPfUKWbc1sCJTUFk9O/+xXhItdG7ihiQ0eSBoHazaoss/Mjl
IEFL4SZChlIosaZQzVCACYtnZwS7kWmPCw5odOVnruDLJFE6Xe1sA+GDNxKb+0yaBRttN9ZqE95g
euOoyfwzYtOAbAgBInCXJ18TVd9y5tSs9PykKBUXS2EJbV4vRuEk/xQ8li/7R5jmgKIpKm5pg3fQ
kb5ipqF9UagXKpbSr9CUvNG8mCg1s541Og7Q7WKGNmXXHupxO7eBvLkLzKm53eaUJV+GzRppxH0f
0r6Do1FUA3LJKP87JKi7+4fy/I9FDo0Ulzxb15h1/kGUDOIPe0F9e9ceW6YA7LFyTmNQH2FohfQM
F3uRPLCSYOamC1dYyqrqRZto5TqbUtvr6ewmziFAhtwE1MeqrihCfQVg+yboAhKt7ZuV6HshMhbw
M0zohDdgrGjtp0Q9Gb5EK7qurBA8HtcT5AP5nlQPBzezDnQfhBoRz7xcfk/jwwLzhgbJ5f70naZR
WhmyKUePrR+w2IOIfm5b9M/a6MZS/Jx4sdDgLMAesvwrflUhwm/5J5hWkneOeQJPqXaiRGE9FcYp
NYshBQs/g1IQGUyW9Xz5BuLgn2yeaLlBbaXAZLcCh9VI68/POWBxPgWA6dplwPffMDpmDAxjbE6z
z0G5ni9pAgMf9I6gRmhkyHgiotQdnUlIYsMlF2gk6c0i4bAGFvKP1Pf0d+2ERbUtfQbMMYvNo7Ne
opp99ho3FWsZPUjQZqVE8Jx+n+idvNCu135lufhHgf6gdMF2Kg6TTtem3HDqtp/r8WodI0Et2mUA
Ay4r7ymXRJYmNn7RFnAemU7ALW9VCWwNGLRuuD/c1ghS4I/CQojhNMIAtOYvza5rOk3Mp1vUDAWr
TRQIrgjbHB7vR3lLnPE2TkWPKYV7BsrDyjrbk2+V2likxcZn5lkNvrRHh571WvwPdXcTd7I1VrYz
irxZT3OsduUsiny1nrYYV/Bq66Y5csh5KgsYkrQmvQfCXJO8s/gxnIqMGrRaoJNiCdvSZrgR3oCz
CW+Vmc+Va0vwwB7C+I3ybtSYjB5+AE6oicKqFwyZti4GAiP2NtE38pVyZgOucvcMn7LZbDYbtEYS
H0DxlYDHdHEyRv2pmAzJHxoO4U855kzCdLIDjuBBOrT0lzwXx0+eU1qC6d0NeBY9QKvH0teHwvvK
xA73cgGe8rzrumrc+TvHqomPhRE+mPzZl5U3/rI4cD9+a7sOoGV/e2cDb2K10PfdC43FA+HjKeQP
+oknQr1Odcivb+8whaRBipEjERr+12Mmf1rViknitqjuvjHsexqO/TGSR3c3b0cAEWnQeqtI3jgB
BozFlfk4cFyTy2qcfDZfnu7uegXK9amCJ2eA72pQYqSSfOLXPAP3fdOPN7/DDGrRNNENOQwQ7Izt
fiVsgHBFt78D9sTLvznIacFwGOYu1FH0KmjaMVltpDfyQotquaA5sZJFrm7HcgSaZXE51yatRO2C
LdUwGqoro5cowBvzl6FrwXsbHsDVf0EDDpVacdyOhqbnD+elF2ayBWZydoVaC45TtHiLaACep/mY
QJcW8nP8GCPVI4ZsLlvz2lIoh7DR+pDRf7osmHLg0JqeISnvGi9K6U8bvFCx6GIFuDJoRYYVYjUt
QDeefVyYRVRwd3HzQOqZjZPy/KifclU95suzsOeWEfHxosiVe1cbKSUWg4fMPJ0tCgABUdmHEftI
1mU775jUVQHV2wjqicbmAg6htQL1/RQqc8b/BMpfGoVgNUF1oRduATLgsa95d7hKAUEiYznbPUua
DZ5hQCL1URW/GHPDlh+QFpLJzZF8NutwMe4hCOIEiDjTB+EYlMe/Wk09W8yz5XDe1eucgpADZ3uj
U2vreLkc8hgGOeej+ANNjYteQnpXhc2FPCI1qDGq9Ui9oM/BTLpicq/mXZ/OHgdL2EPsy3nk+yJE
Ijzrrbbl58Mqbi/6wEWuthuE01VGx8N6VI6GEDXjLz4KbAUAzuVBbvz1rZPlBHp+fP9abIJJlA00
COD/PIC7+oQQgsrk+dEeocSMPEi3AFu8Rm0Y99SgOo2iurOlbLeG4Msag60F1cSnMBbNjehsdVNn
UPMN3+Y060/UPCKDOtFh6iXfICZvNxdtOCbl40Kmfj2IL0+CDsyyaQjYFHmivlCRM7QXW5C/Tjds
wo5shV/ZZ+AweDoMu2wd/RJ8zgta5NotUQsNpHGwkPxpCIrIIOf9tDlyL0Ox8H151lFgYggZnmyv
e0Wsgx4X5SquCUAGFv/2DpCKNDDgTkO2BpM9wemRjHrWT1eWP6JDTt1oy13AFq0mA0Kz6yLY+FGo
+n1tjCQ0b09i36Pgp/4/kTimYVs6tnywlZtvFANLr/coCK1UhSqBtHL1V92AuA0XOQs0VNh65lJE
1dwWAHjmIWAISUyXxjCvEble5NSN3++B0yo2hyiKjaCxh1xwLKfmp872oXcSOamszq8KBKp4RU2w
h2mnwtaE4IZCyPrhp0+GT2KD8qzc9FQbstJepA/qjaihJhN/BNZ8AtDTwMiftMPuN3bq8Cdl6Sb0
DKDoLS9X2kDxHqz1JSaPlNM2cDyKQ7zPlFyImsjNxHsQcoqwnvjLF00ByS5gOZbPgeIJbA0KIprz
at+FNQMnoSCgJ6KttSoVNOwsDUjo02ubnUzLSVnIiEvzM+gsYf2x9u0SSA9j0bUHHfiZmQBXt0uZ
0gHB1XebqY7D0FhvcFkXgQq4Gn+xSFAFto0VVghK5nP2mxdIemoc8TWKW235Eh88Ear012gnxXnf
qMq3eZv71NZ43D1nTDMP+uniEWn2MFQBtKv73fNP2uX2zagKGB382l0qQQgCB8bYRBeXufIr69cA
Wq5f1xViZCLv0whWf5Nn7pyyQmzQY6i8T6YNHDVjy0V1+HJQb2TXK71o9dzA9uGztkv3DiADWenl
+8633hLyDBQ3NdC4lUX6g5O0ywccqgpRNsALRjU9GKRLmSVgY7sTmlIfD5lx6t0v3k6A2tsuuAhS
N3CzX/S56jIexkpXp8jX+pzR3DzdS3jQEjmAMd7Fa1+MdC6q+IChO1X7WhHfgQonuz9X/51Se2FE
uDv+zVROEMczxs4turb7A+HGxKtuagv9rS10/ESbPfQhmbzXijIKAjjc13dShtJXFsUBsIdBcB8S
Wzu16ei99IaVdCrl4zTJyRis5yZPmoa5avvz26Nbk/8mZtmerVqZsE7c4FFGSTKjS3FwPR2ZZvRA
Q4BXiI0ACVP7p/MMpWEDW4Baj0mXz2cYb121xytJbq6d2YV5IcEWutO788+3dcWu+9+S0Uakasdh
IsxHgnNsdFxtoGCsVRNZ/tCtin5g7KVtwewIdk+YjSxuXWL1dkiXO6+71uwaP6PK6guaeR9HfKIm
3eHn5il6OgpXFNtBzECBQPKZpih4WEGw3Dyp1NasVxpbQeKQSlGqkyYppbmJCuPYmsKopSSc2LXK
qIv3PzNKBtcFVjO4SAmUhrKu3as3InqBqSoqx2HuYJh9CGtsfBfrn5WXlPw5K6oHF04/VoFl/2E5
yShaPaQGPe5h1K08UXKbTPHFl+a/JKosD7L9tZaA/XW3E7B3fY+6DDTYakucjiWgfOH8J37ZCHFc
xXmblgI+UXaj0sjmsEwKMVfEd1VV5u6vwZvHtpHL60021/tB7XFf3fqoe/kgpHrkRARii2UX9Tje
ifxmTJ5dzTyIdyfWumR3XQ4YfdOU+DQJRJ+TCgxe+Ns+kye1UQDFWDF5p6z8KqDt06dQDPI7+3Y4
8DBWA4c333NyImOPpNmWDB0N2RJ1wSrqxSYdNI9JWZtmdp+KST+yyh1PSqVDLqnLU4QkaYElDiQD
LxgnsA5h1jPRQ0t9r/FTW11VflD7CwD3to9aVqQm6+nDm/tuwEqwftdeXJUy/qpJh+QycY+pGH67
BXFlID5gKVkHbpTSkZr6Cd7mZoI+FtkDzy/1f5aSli1+ONw7zTjI8hpZjpBk9B/umWPERLGbs0Ao
QM1oJ2jIuTEkU3KyTccs2WSZclNN0oNhADhfPx691psOKwtYmah3DWF4iIgxZRTiccJ6x36FbytG
PcsM6NAgeptC4gjeJve2zhrpTBFh+eZzw/ncRHxL7IkO/y5WnqnJeJq5nazSDHL5XI6sSV8hJrqx
0S7mOQbc1z4nEXaCVNsRTHAll6NGCT6LakF4Qb69WzLBjQMZWzNmGFV3H3827bNrH7lMtGL9pze5
V4KcV9Oj+fYOyg6+msnMldImq/h029GW88uSlRAaLHyzBT0jtrhBmZLRP+pMiKQUcwjlq4zoNHsv
acOZLOlcmt/OkOfKuHfxpZj0poD7tIYbp9VyVZ2A+mdLgXo8Ycwrk/9Sia8qa91fLx/mMjI26h1b
UUq3pQQcGcfYmhqHiM/BsShxu3zO6mWxT96iBePORpRQiV6H0rgIE6tgoXeur3gsqtzzGNgX914m
RmGPcONY+OCYn9N6SHTB9/i+O2vltXl3XWylwBBACeozygmWSohq0htMxWExAbsJ4kOCUU1tmGPj
gEFXOEq8wZvwF49W1Nm10qzCIm0CUwztQXhW/Q/4bopY3alqBt33KBV2Dpz0QsUzP4//YFt5FaTg
Vo6NxBreHM08OAhKhTPdPCfi0cTujp5lA6UgJ/ipxbCayPK/DwgCKST1Jw3T4MJ2lcgQSk13sE0d
gm0dpBFzftJI0GkjreGN0si/bmXBF+1KZpg92GExKpYC6Iuf67bueMnoW27XLUfpsIV+EEBN47Vj
3j959w4NxHCAoKSnNIbqv/yo8UnUORexh1gU+xK7Ci5CwS6uamIL88w+ruSHA2Bb6vhRWMqyrw7e
S8jNrtzWXlG7Ujyzop2QmUxmqPpF3OwP6sI6xgT9+wtJycLeBvMmDwLonOdjXB+2bn1PJFnb1dW6
prh4ym7ut7u8u1u7tPC3M9LRDybZ4njl9QqalJ7PbDyj8no7O5ozI2zQNBpYu4oATDRIb5yPQv3l
JDzAm9tVHWH7YN+/gYEhNHQG2ZfcJE1eWE64v3nDvELdIKAbN4TtChqyz031nnoiuvQRNNBQ5OP2
uj5EaR8Agh3Uxl0FNyMtNj3c5/+3OiaKU6PpmI/hjLCw8J4YCSNz5uGN5GuH9KK42tsqiTecESN2
JJCz/fou2TyovDHMu5LMIXmCGfSPLaL6YkP1m3w+XmZLGBbDHjCB9f32RwxtNUa0riMuDJ4QuHT9
kajBWhPdnv3Kjxf9ZwUE+OtCTms+4FGWcetGSiK/aIyz3UYhrjkIbvjFEmEcSTIC7GtNjxjIaXcr
B5yyhI8nSr2SiVQ1gSygKYc4XB340E3mzg7J979iT3HjAkF2+eBRHt5+PPHCp+xsygPgUwmbzDd4
6DzIwoGBJI0eI3DKedupKef9fzZ0mlRtC45P5/+xHGdpJ/4Vsvs76RBvU3u6iOYjHackule1T8ji
+mlyLl24YUvCmVv7TNd5ot5y0lR5RHo24GE0POBxCbi8GMP8kgZ+X/gEO7ionA6kySIw0euhzwNt
XVH/Pl+wsWyKh8+vVvK0+TpYcT05cyuVTCDEMBRG4aDKm+lf62USSk8FTmUZ7zQrsNbP81ZMhd06
Zxo66D8j6Q87u9gkdheqYrgmgXUNk3zFsHYbCI9+fUbrQlQI0yAyk5d164xpeoqGlSN8XwroFMXQ
EdZCB1VrE0eupXGl7/+DlaixsWuX0qH1OKmcat3Rui8/PVVduW9D+WTQOmq6fdx9vB3V8TBoEzRA
JjUV/Wci5yI+rit4KQCrpAauZm/7SiVy0W+53kxAfcZMzAlwk+PP2sl78V4ai1hIO8lp8VE+cD0+
mH9VjgUKzGZCim412YRkVoqYgFJpOlS7+XB/gQZEJ2py17l/VftDzkHWywm7S5wEITmr9TLXhfTB
kFiTfFOIF6+DhcSPuEDbpRo3px68O9JzZrqmeopvBjiiT/dEDs+tPV80DywaW/Y1IQpxYiLyEzU6
OOxkJezB3QhXPOQ4RXgXbzqcIAmnVOeAjL8lMImtHpvuyEWnL1snvJHQrFavlV7NEEhiNfnRo3xT
t30IwThtXgvEMChNvjRsfx/bEso3KPumLfx9Z0rZf8svbVqC3zUIamcpQBaGsx8znpDAsHCjIexX
Om+ZLBJ/Jb4GTrfa4zV02jGRFvV3tvPH5hkN+PwSyYyNdKGI22+Uj9AL4I9nhwFJFl8X1iObKCkr
61mGTRyAymeHIKndbf+1UnHaDMWfWD9sMno/afDglDwObvliLezu/rKy29ym8adkQDv3W+Zs4Pj6
swonIDCkAI3axKGelGBGUQCTbKhs8/08xhgzHT7oh926Al/3o/OnWx4IlQB3bRqLCzWYldLYOzUx
PMWAOCS0VE/qhBhxJRUQbk010ih/SC41w6oyK0KMI0iNVEIf1g/CvClLuQ8o0pizgGUhWLxxx6ol
7yGOlbUjVS7yNRrADAXPqoskqOtHcc3ZhonLxbGi/sYnFJr7pj+S7xCLkuIPdtSBtudKTNgrSe1p
FNnEv+Hc1F427SRFe74pyU5Xg/FPZa2QYkpmWF1DG/S7Vxv+T7C6VwVcXf0JmQyJdU47YWVKaiBF
NmXZHQw9uAEM6+6is+7mjbCgD4sNZ73hDMhcP9Qwefok+tEPBhV5/MSEtBEiBZb/IgxjcXPOzEVs
V/nR8TEjgnsdd01rbniq6mxrYJjkBcyJ8zd+b6qcftr6tuk8zvjKQ1PB4H7fjR1N+0VtZ2n4KCfn
r86B0t5dyv8jNUrXx8MYk4TmqHqVAtr5qDhpf2WFOcrJ/QJZddXFFVNttNTGaFRusVVjXp5y2Csk
TNoyrUVXD3GxwGkDioArSdGO2EKx7RqX4SPQofCweNkFgcn66SJ8GUk/88JG6H9ksEjI8arXa+18
tHQ4rnDHtALWpbJ9ibHs6DFPtsIzdfbv2W1IPLYmPfhT/eQL+Lg5PwCB+0AHGwXeE/mlrHnRmXKV
Hcukazqlhk7zlpR9KwRzXuxqc2lDvFA2uEhzz1JgXBDBL2ye1eGtA9ic2jUnkh4LN56RsyEtkTcc
GNqoasjCRujBNR8c9Nlslfd5HLmJLaFF2RRQ3ddxEA0vcapQqMXtQmGzFeGLerMs5c1CcGC1Mskc
KwrvqQFQE1SNu5A108z9ogANh/yVfFJtx9CiORlNnPq6631wGpGbl1mDTAETGAgp+dycC/qVOsjx
q2C+D2by3EcIolcYx1HbfjMO84NlVZWOcUFM+YNggkLDmgu6mlSqKu4d6YTSAqwwypCY9El8p8LE
tD6OFZ8sjeuphSEe3RtEa/yb2IDdievXEbPyDrBn6164zMH6z23ZopZeknmI5c3PJ0JjHAvOthh+
sFarZPqMFny6lgnfmh2Bw6V37anggVVlVMBPqrYTfh8SiqIIcg9yHlz1DMiletQ1WXM7vODV8NtA
wYNLn1qteuN7Oc8c5GJAZfrEaiYpaNVdpKdjld611q4qBeRTeTApstYKkAv1iIvLh2EPoJVPkJXR
EPqlHsBLQRiU/XfbcaN2sgn8NQP+xQTWzDq5Yo7fdkjZCaLWfmsrn/rSUH8DF1b37Mud4MQhCD7N
8dJpWYpPrY39swWNAYL081Xg5boSNHVJm4TZ9nNXhceyMYN8Dru+Gq9Vmed1y9/k8nVp5+Tf52vm
S9BBJTKEYzi2aq07whKC2V+UmXPmaY3SYaFjwa4Wr4H8uS1YKyCesuHuBnVrSSPnLMKJwgQ7oHfs
8dLxngqHWvZcB+SdNa8zq3HTaxuJt6am6YLnKbf35vZp8EvyCSDkUbSUSkRCqdYqgX3RLiq2nHmF
SnPTrlwZjBgpVotSefHGbLvK5TeLAu1oJlGrfaXsQdQfLJeAKSVevuLjS12U0aFJMRoyMGfN0VnC
kZ5iHqaGNcsGf5tByFWnfHxD0kLi2auk/6jHfWTw7SwnjhmSQgDuWeu4TqMGON6rDedQnLP++Ivt
WsTeMms7qssq7BaeBCVfUJhKLjE0UbbXhF7JbD9fhAsf4fPWUsUU93k7J/WUalRUj5daX91C57Wp
gjX7rJKlBfWC6KM9f3Tvgv+v/WGws+tKPE88QY0OUqNR/KEAZIOJMv8Ylwi2Wy2e0sz+U0B+bWOc
xhl/ghi/Dyv5JMWuJPrwBd33WkQqrzDxfc5URgKldcgq/5bDXtbv0dulVnVqg6hVCJ+PkytBV3yv
r7qhYtxwk+aGOgusRaTt4KPX4UJeKQr50rYpHeCUSjzYxw2qrk9bp9xtspkDxk8MW7y+pZlJPmxF
1Kmnkp/bfU6MXo+tiL/o8O7hSi7uIJEMilXCGR1M4mdqoKbUZY6FEwcDqyaiReM23NDtlUshDFju
afoiurZOpMclfpO3CLK4rpU33JtUBgbpGsXsH42G+dTEY9iZjVjCehHyND0L659fPBPDm1LBhXSV
OqKcgQaePzSmpw2euJYicy2vKGOixUTA4XM8EzjAry2q1hTlbcmqAc+cnFh3EBeXY8ri7hxtYFXD
k1fdpFpdx+kg7wWbZSSql0TjiAb8T4LF2urvudJE9CmZMBxdg2UrxQiz6IU5chrr6mwigjoTOdqL
ZS0Ty6DwJnpGP9ZG3N24viAUtIISQQMswuVfgcPtNKYGYAuLjXAWHWW9ikFlUuH1Lw0gWM8ZIbcZ
O/wV5+DvmA+iF9ACtJY18bJmpzXpjn0ZVezXNZWXZzO11M1Bi5sZH6CMudFwFyvU5HGYn4r/4dPr
vYcA//syblmGFYkOvwI4vcUsJ0QdJ72yu723uMuI+APi4S44gDDOLR+kMIebuvy8FOics7Dtgkwc
yN/aggvYkOCzNzYq9Wj+QH1VJa9Y6ATqRg8p6mwGUNLvwe9yg/C4z9JR4Zm8ccPyujKLpCdttkUD
YM9vJFflqfgxetbDyZGNCyu4szzDLlljrYGAlfa0DgauhnK8rOmSQHYPkK7fp0C9wfZIvhDl2dpd
fAXxYbIQsCgZxsjhR0Q59WA+t9VGd/vCfUwy/Ec6NKeKO+JaWF+nqgmF3xHf2Xbdq3ghsNlpKhjN
UA9JrzTrSkeoQCbH12zdJlv3nT7FT8kEhLT+PYnagtheUipo5k1120/i3wImKaFgiBwLA9gnmK9T
kOMuUUnmVGAMBiKq0Npsbztg5FA3B1ZKTIUkZdWdp8BJs9uyfU6IrpyAToN5PPbfv9P7lXi8AZ7Q
hG/ol4aL+qQCInAK5OwQ/mlzxRRL8/kVgWGhQpJu7ki6DMB/ot69tsBwKLjKn8/v0IJQXODzGQho
7qh6/PAquIgQE0KOIphco9cFV6ntQ5FUsDikLPP838Af8olwOEAGKmDU8TAhoXj/0jpYDDbt51gn
a3nvuuOZPxOUGcAXPtiynhFQ2qENTSv8O2Voatt/LSvWuoHJ9bCwCs0CCTy8PH1bu/dG/QXKsKL7
AmiguMeoObdaVZCUpZ0Xm9SWlwQIScHecinlBNFGEUUrYvdhKtA4nBuwS4oxX/6gVcw1SylKeuDT
9mmHxClqCTFWFvWgX2mI2MQUM7ghjG1AuHvJajCgsekkHV6gdVwtaSU2oYkVE559LTO6zjwa1qd9
wk8eCyr/SbbetmPMauMDi0swkZhEb9cXqsD5w8RGeuBRd4URXNcl8Uo50PbqXKHIeY8XsGJR062U
uJg6E/omnJQWAWuQrHetWMUQfQzgjvBzoerTslqMLH2aAdc4rCMcC651DUiOXGsjEpSuJ/owZDBk
BR1G9NB6jfllJoUkrPI32scam5KWNUn0sfYW98aHtGPBZWJrApix+lezwhf66IGJhPNGLENt6YNr
BqtndVWSvzbqIc5QIe/7j3Lt/WO8KDeTW7MEKAkvHNpU2ABuZJel0CdN9miVOYBBC2tJxNMJBwpL
XiLqE6o20bZe7hq5lwC5yy7xGKsC9ZiwfmR0fyD5nUrEakANcFZgjIdW+B8DhfroTumPXSiEPTQd
/K+53uPolytWdwM5MafwoQgOgj6dP5jLGIPb0LLR2jvnfe7tN1wx9zBEVmUKoUNyYnxoKDceQcyi
ezUqPkXW1w1UjoQSoxlu9ZyhM9D4ZghZT51kSx4fq3LOqS01Mg618I8nw3sIRvNF2bwylpM83lFA
WfuGZ5s9s3Umn0ako28vCvw4HZonT+HOLfDUE6RDdHZ31mkTPswW0cfjU7YxzncTONfsj3/mhEU3
+vSJClIZ+mPM22vR9KRN6D2ioF5VvhNpHdt2HFQ8FQfWXXtP8exRDBgGKE3ZX/+uZaqfCMcf53M0
HW7xmmUtVFa4uIqBbwAemnv602wAzagIlpwnMdBfHLnnGiBlHkk0fdSNp5hoTa51peQmW0gs/tJ/
d6+tLKyInGK9p88lX8ExE0jyIj09Xp8+uc+R9D0NLAEGbFlBPyEkXzdNepUh6Ip1VadACZdsKdzX
xw6RYgi6IXilfaE8xVvO7fveaBQNiwFkzbGEToCXmsAvbvnuxe5+dJuUKTYlSidovvgACMR7tv56
ODJ+5/0nSqZ88EgybfiOsmPDNoCoZCS4OgJU+9ZIXDxMj4ngloMBCIpXH9bs1l5HpRfEzk7abBaa
l8TD7QHXQg+6P43Lg3nRStJfmi/t7CxkoWn1LuDoLGC4Df7lCEMDpJ3rZZbVbFg0RmXxVdT1dC78
tfL4H9Fp/6AlTGW60HsVQDC5P092/P740yJ29tCC5VZgsKN2qBGuakio+Ec+WH3R316RFQorNsuv
fnAyW3wsCO9tmK1Gdt0m8w4aBKlWRMNTsXLwbpIuH+VL7/pl+Cz4dzoObRX+uIChPEE0KtfiT61W
6A9m7SqKtMkCpTGSEEeZhgmAAWX3fRUV/XDVMPUioQDSgoN1T7Jm5g2i+39lq2ltA/GCao4Wg0UZ
LsX8ceYX5Rv+55N5sqwVCc0hl8GeH8Tni/6Foo/LvcVJhC/BIKoFu0Td2VCIhgWhQ3lf5rPVmDcj
XKkGtA59XsxjPPfByD9HrJJVEheJ9eT3JVKVmo1d4igT9mTl/83PA1hRGGuE/RZzA4YMpckXzjTW
Z+PjAho+keRIaL++qloZwz3YIM8xArxN+M1GJKZ4xTGBvBdAiOwVr+Fcx1wTcyENXP5NPWC8Oyph
fPMKQsEHm8PTPlFWmS6wR4Z+WYBK109aCWAtbRK6a2QYj6KdMqdjrzt21JoIDcGuudSOoKOvDnPz
5GJMy+3dwwjOH3I4Vtet47jGuRrg5nNNfGptjj4OWN+akZS9yfC8DfH7wtFOtpcV36qjLLgOJrpx
K+enSvDU6lcszucZqywdT76ZBQvKYbraU1kH1RVDSQ90Q10zM97mbIGpjb+aKqGM9UC+0HYZO5dY
Tq+TFqCPRD7SkVW/P1bfWe72UqkA6Pi2TpoCRoeU7+kJKjtg25tZGdl9veEXKDBeBPYecjaqhHNd
VrRuLTyuXqZEcW3Fg7J2CiO+ivuBSFMpDuZy9RMMgc8mxwaAiXDQyoRfl8vmO3VpxVSV84ex2LJu
Y/unv4SVD1yu0WjG+Jj1xxNC3B4NZ5r4vfFWbAAyPRASVsf63asf+29GEh6BxE3JHfHoxFpQOiPt
AmdcmSbRsiuo4K6Q7EpTSWpxm9Ihsi8z5kUNv1d41y1Im7dPv9fZQhYUgW7hXVOSzso1sDq0nZaG
mE7kiob586NfWX310o7rYLpRMuvizwSsbP4E+m9PJK9Jsa3QXwZrX+F05SiZEEYo4q5coWao+UIa
+dADMtPU2CNhhteqCGzKj6uc8IEaapqG907DcLuSqHeZKxl1eCHzXjTOBl+YdBQisL744PqBY6WB
dL1h/dFE6kQHlBsWtHSj0sEChcMMfhjBC9+CcYePm/KNTX8DamX8kj/duEOQVpMSWKru3NOr1Lto
WPY6arZDTEbu+FVNMzKtZp/8JrXw266yxHOVL52IRV1FU5JOy+rENa6F+dYuYqt1hl7T18uY/uD2
OslHpb5Ff046LHJ6IAipFmvaqGvwpCiT/6sOk39Jfj9mJxFGFx1yJiX11R2G0Bzd1n3TSAerZ7Pp
zAwAfVkCvqRQAxMRNnNFv3LgTTcUdd9s43liaPiwwPYbdj2jU/7UPWu0+s/c4YNH+SatCowC7FZs
SgF3CZYRvrf2naarsxXcTIFZ7VWQmtFhuvIOkkBAH3wUTCk/GzT7YVovjBb7/b9/+onxoq9yVrCb
YJDAt6sCkGTKj2+4DiiL0JjdDGMr4CUZG/lXchUm46cBNGHcziuddWx7yAEabm1UixIEztko+wbW
2dyvQ5exQapFMHOAQ1B1n4QIxfJOlmFSxbcLIjon4VVzZz9CQ7NRiEGXHZihPmDnOU9EGrtyoHWa
UMWvbKvtN5MBJ+FSJ2gOCnFTPH61rN+jU2BkWLvY7PcGDTAFtQTeVUTI+NQiIiGYY4y/9wTUSY8X
LwpY53K8j2dWuqvH8ZTcI29ebjaXdFvTwCWbCNgVGNPEaQ0A3JKo4K9ie/CsLWF/CahDTiFdWkKH
HXvHmLOrTT4UfF5NCPA4LXSQ2dKCuxbVUoh5u+k53DT+WZyMy66N6dWCZb39R9q5iEyC9ejzmiw/
G0Hw2vhlz8ddw2gH3TADRpeHC4e5s/qWTFybfQjmfMKIjftQIqr9YZS+PE3nEJBE1kvecv/jFr7Y
JzjLkvl7Bzc7qB1FCstfjHZXzhxofu4HFwqbx7R5pbA1c4wFqOqvsJ2LRYlX7WfXs4d1gOXaCcyx
0IlkAQF+aDDg1iArXpqVMQQJueVxKy9GWlNfC2KuIQH3I7JsfhGR6O33Usq21iGfV4+tAQ/0khkz
7kjp5FvmEhUDY9d/bBSEF2RCsMJ6kefuNvxtHbYAyan6eaFMeU6ILZM0nrn+kb/Lx3IpG23Uc4Uj
njLWgH1BbUnU1/v66MOjIAc/SA9LBgusR8yFA103jXSYWocjGBkRY03ZxTLQXV0kyvHSDpjxV0VH
Fnw/L6s2P4BXL0jvYUQA+MnCAnffGwbAMm0xi/Q1DEWYT39kfWHM1bdmGI6jcsPKqgb41sT6swkn
NjqsjsDI3rGftn1hJhozhzJTzygxOS4JWw6yYX/tGcJNvo4Lhu3LqD61yiBCaJZOI3Zcdbara0jw
ygGi0Wk7FZBtaMD5e/+3gnbaO0mrvkEmzzbiebIv8gJ/t0GdvRvC6z+vlfd3n/TqgnhTmFXEnTVh
v+YmClu/QkX2i1KGDs6rQZHBVzjsef+UIzW7IiOwF0BzboUoqNMzKPyOWh7Fuab5scbxV1kt4c/5
KgnKpLUsblr/BoR41j65vhi5EeE9WqR6yALtUyICdCw1q5yp5CPESr2AVXeyo496H3BfmvBqfRd0
DddRz+/AIpO52fP++drlOJ3Tw5BIf4lB372bg6l3PhsY7R3eWjri3Jk3hYnVvuQvUK5/iYXG6MeX
fIDiEXwDZDilnqEfm2LZYnsfPclXwyMgINAtDMDXkJXsnS+zyjPjEuyK2bAdcn4PXk+Jq1H3AvTV
sDjb6A97b+Crl2uDjN5lh57ay56f5v7BveSo3kU+ocoglqg4yBIX+FcLUdvK4DICuxaznKldBTyv
y7PMKYLAYOA+hEORdfC1NsQAAlfeHncyS+x6jASvXF3QjeiDOjS72HSeQQv4s1+Nk9hw3n9MliIS
+Z0ImHBsqPKq+2hriY2O3gloSVPhHPxhvPDhcbFLe622/rJhIfpPc/byIGPtMyixPKKWvs8/JLK2
QbuckpkvOzLWRtAEe2rbIK9/gvOUIrDJ/n/640Bfl4wYrGrZt7jGSG1BK9SIAIG/2N3owaylHljy
c5nhkhU81JXVrhyNNaqitOioKMGifYsFZuN8hfiavK9txlmxS+RcCNsCmEwLZoMPzmPewH3X2U4F
Pzx6FwNdRxaNNu4byj3pbsBIWrW7eTBXkdYVb4DcN086YbJipJcmSvP2uoiYCu/23mmnSP8hR/Vb
f0Oz6IaNHiXQPHmDdyUr+26Ox6CyKGXWngPkWufLun+FZ4YG6goEHTj4GltZ5itif2+EFf3ylWgh
4JtG7q483H6PUePfE15tKTLtVGOd3g+x/mE1hHb0d1ZZyw8ovajp/jdNWE9vDJyQTs4esKj0ls54
HsxSLLMuxBmopFkSJL9BSeN/CsIquPrDf56jZCb5YL/hnVTIfVQzHMiOo6wsxBXl+FgBWwsBf0y7
cxvAOC8+pjT9k8I9MlW+/n3PFiF6oSTszd42xIOj63OPJ1NcB93t80BiqC1il/0OfUAjwMa11ej5
XEJTdH2ImlL9wQo2W8wJ3pCB+ebRPg4TRwNK0A6SJDmTTBeSsViUNV0+m+87HoU5OvIwM2g8vyHz
LteyJPhN8k0zL5P4LOUCdz6nNHDd9QL0ZSg3oF0LLZhK1F2ZrwbHp4tWq5ob+3EjYl6xVj36hRme
4bAcordRnPIJxMXigAk4zMOUs3JadNyXsU4lMFxfJ71FeTylj3z0ntaoeG+a5aHLn8qtJ4BAIBBF
wuXHqKQm1b4MyxjhBo1zvKJ3jJ4NCfK++lHf4/IoAFmAdZECjNKd1+A+mUkxTX86dllLJPXW6LpI
wLmXseMj7ey0vwSAHV3VMT/llJcb3VDSmehgfJmGyjQe1yi4Z6wCeJ8qcHPxajxrrTnFWlL+p8uQ
agHNwHsl4SmZHZEtDUvpp1AKemoGJ16ab3mzLi+adEPEko72JFdKBsBf+pIpnnd/t6p4QlTB4yTo
pxWYrgZuVMn/bGCzTyV/GmfagFytjQH110NuIwY3eeBfopKz7w1ZfJDm7V9/5zZ8WrN9zLYZCNPj
YmzIXK8TQhSZ7bmnWdbMA48+U/P1F4SmsV1x8TzI/4w+5I9rPQ2inI/87k3dAtsKNZ/vBBFdvQi4
50KW0hEcMUCPCLbP6e/W/b2/5iP2y2oJ+L8D+/igy/TX8Qu2ItNJXxHkNnGc7Cyjw8W5HQzYXV0J
uKyCcVbMZ3fXljpPxCkgT02O8o5RlorajMTCArFXrYmLEzq488QclMDFeQl7xy6op/TDWeI18JgJ
legRdPMT3KvJJ6z99zlhKWNWCsHghpV0LBUuZst0BYrWsImtdDIj/yTNOeayvge9VSV3vzmBrlg+
0+GJXgsEIhdS7Qrvtd8NOIIzg847deZkdtFXZ+okpoTavm0mlQSEsXlrmGnnfv7OCDbB89qxamLj
9GPa3+JwZBJvGOoSTwhRBmFXqtD4NiW7cF606/oyQMCiJTN631yhPi3tfAQBiYN2SE0ZdN8BX+E7
U22bTVqoIUT8cpGeQn6Lk5hnOP4AfHCbNrqiga2D605vAkyhlVPcPc96HDa9GeWgo3ytFihNvZcy
pvn26hVsspZoewfn/DbFWCd3UdhYhf9xw5D2GUzMgKly886KzOncgi2IR8FQqtibr3ehhxLQweZ/
kYK9zZsv5q/mdqsnGjNCpSywkILiCB1v1htZ0bjDBG6Q2KYADX/TjWMXamxdjGnx5KmZlBbaJ6/v
BsPIC6YbGUeDP+tkoWeYmeOYlDGrv8CcI5B5XCGQdiUEraCuFtPSwVnrgTLxonauKea8gBPtweVL
UPa893Ke9NqeYHQYcdwMYUJd04TSeS1pi1zkkuC7PifSFayN5hIJckCzoHo1B02kpqZwf87Z69AJ
eKqRoqvMiCf9x0+iAmTaVtJL2z3gl3O4lr68SZJ+9vdXOHT90cBPXhTR3PdQZnp36mLAY3LcIpwD
GbAel23jVy978ah3l3xd5jEEH2I1AujffQltpCI2j/Lfmdu97x+TURZL0H5Udyoty9Oyi+9MaOl+
FpIuRF0TQam5Ae0s51BLRwKMWlWW1H0h1PzgZe5BUqH0r1vylrS5l/Mb4ebe78b+me/AzaXy/DYR
XSEmwe/MDmh2AKiHEscoAP/mD5/QlH3pensWXpTvJWISHV7oRiSBM7Vbn3hjZQJhNuLCYE1PC1Io
CNTXCc9BfPobPLKf0FjzS9lVNb5BtS7zDqXxtUbqjIE3iUhE32efs8ur9WCReoZIUTICbGA/2g9Y
yo5tW1NcjNBiq0lKjVgFVkbHNy5PLwCLwK3WviDcL6xSv/IYGJdHEanx8lU8z+cQELbxg2fi7mKF
Is8F2//gHMotfONAtqBpBGj61kR9CgpCikboTWW9tWFehfwS4o2GKba81AP+dao8eLbZiqcUdjCM
2MirvNp1PYnERX80r63xC6B/cwxv7zUfx//zS/K3QmvgWVGZhtdH6jIKownzhKNR9zr9wU/5NURg
NogA32dcuEoCgzWhWoTrsi7+HsjngTBgJ566rjwlsi4zGLV2GmabCHV9MhxeMuzZWEA2Gpxh/lg3
MeOfxnN3aXaIiaoWhkVbtyTCV/Swo36SNxf6NI3fFuqeiATpiGHyts+Dnc8GE+muwR35jvQWtsT5
c7ggUXPE3o4uGhrA6RgOr+wojVvkOhZof8gevxunkGj77yX78UNx1xdDuhW88Zu6IeWJmajQOIwX
JiET4p6q4XRwtsS+SB2c0eC3OGqvW6eNVlXKBeI/V0iYTRkdiNZaPEStcC3MkfFGQv8dfDkLzVIo
+peYVJqvTfo/WMU/z+EmLooxFrPA54Wk9qSKeuVonuMFFxtofsI3ydBKrzgLPrDtIqgmzeDaseW0
FPgRwr29eAVL42eBwkAhJUSXpYikTtiErxwO0+Lw8ix0DxxxeZbmwVhOkIlWwy2nR4DJcf5syj/f
LL9GAz4e56RWgb36YdHLmvYhDvMOPuXB/OyJKibcK4hYp9nhkoAhCRppOxODiv0josTUgUk7hnEy
kG2yMU0ZxtdgWKQUJKQyT2NhW/Lvn9Mf+WJu/C1kH3mRSlVDRCcDrbwUiq+Zgjsemwf7rOrDt0Vq
itep92H8PtrHQDu+0ZBgQiaYvrmYfmCqM1lAQMbR9UjxC4k369jfwCTMACuUTanQ11xPMKC5jUri
VTqTuDZGr/zUXSLU39tSmkRPfnfEUTW9Ra9QRWUlBMjPadRZEI94g1JTRNVs8uUf/5w7YG5+1x1X
VunvMj4eMq4Y4TiOJ/knqvKE+xtdPWMkRUqEXrHCCn9xuSnyfe9hK9i0FBkUf+sDmSvp3pYCHbx8
NHkXYSSiZgLrSnJU0Knl/pYMhfvRbitr54YQA6OPRhlkGk+MuZIxWsMc2hn0C3iS1nQAU2YHHJVC
oqCT42+rw7a2OejWXVgXHhnzjMXWDQI1T1rgnlRseq4aIrOOH7bsJHT8O48e6XNz/f1sz2wVD9HC
j9+6weH03LtDv1tbyayRa7CxrGQ3H4tQSlT1PJZbWKkFkCA9TLqEglSbmVCJeYVjtMnhWWzeP48E
EM7u9b0flqPG8yRNtYl/FO7XBtnyRDQe5PktaWebAS/AF89bY/wyDpDgLhIwIi1geU0APdgAXZO9
qkhKT0GhuttBl5nBycVtm1gN62F8NdKoCvA8FPIpEg/B0mzqtHTSeK7jk69yLAA2bHOaBQXcMcGp
DSQIGJ4anX3vuQQP9Rzi+pMR0EYgifJD6O+LUCj2BtG9gZOkPq1QDNY4WWwNpnM5qcgH/1WHKbHW
B8TZLm4iWS+vxrTOYh3bIlu5EyUX2dqClEhsAHksHqXjfohAAcQ3b+6cWvWKebdBl/9kKnd8UHWW
RCTA+8aQEFU8whvCeowsonla+jQ0OhiEyh7UBsDiO4GFVTLKbcnBKFI/iX8UzfWgJRr88NOsaeEC
Q8xYKoP/68o9jhClopFOueleRkRoAt789DyUDRIqsWVvRnwPQd4WuIbbKZwxU9Y6UaV+hYpH9S9h
ItOoR7FWIyd6W35cT5ZWVsN6DwSngBvqy/iFxYYGGAPl8IN2GL8MnPVwCgF4/aU2ILrgSHKoONT1
/rwlbXLDjhAQ2hf7YizfscW6c1v4IDJogcGqMgkuYEWmxoNKu1Iyk2v118u7OUqQJLDDf41IaAW2
OvRSS9aEegAf6sJt1ha45tOQGTu7DNKQdmna3uW/5Oy3vYit+dnjtmQqzxoLA9v6Xzi33xS3OvH6
GvV+jrT3QrTwkZwT5Nu16orBc3ku8I4Z/AIPzlYzd3ZXHJ9MybSRqkEnq75p04cdBzQQ5hkvEWxO
azmtznSXpJr+H5CIFutJgdqKEMyJmwOzgQ6BGQ4Hy9LOc96yHdrHhiNNJXTVkpjkWu9udzgWoJIZ
MTrhxtI6mPPspSlTV9ygINFAlOn64tCmGtE9+Oh+lcEbdwespKI4r+7iyjZVvhlhNvDA1LMoxejM
WwNnYf7bL++ei3rG8F9IhE/gRBBU5CB0J4ovzQLAYZeQnp01T9ysUdZb0R8x4UN+JlJpajYMknXc
IR6/0C9ajYh49ukarv9FyNRiiOgzvBn+N9rYSxTB4z9+w0RGpCEp3HaVKrMUVCI6928J/mat8Dzu
RE/0+fa9aHsoBRNC/3S/WkASTr5/Zw+1nnGsk3DgyLkZw7ERJQ+aWSeYTEDmDe+sOoPRzyyLsY/K
m4EPaj7cCmc6OMNdoCQ46jqO7QwdnIfQss9zEAFjr+yMXpW4wQCWXSpUWUhHq+mISJqUwWcaknmr
9pTi1MPEeAxGdoVILZTR2AqqcPjgs061QxPa5ZHNKxvfLpO6NCUWaLDjqN23RXW9sebZ8f9E1d6e
nBfmZliNjsMmfdZRtXbtn7bkCxi+pVfg1WZXqvSiMqIv4RIoCzK70zQ+9diUshCua2550RLNY0oZ
DRi1LwkbXUeTwPpXn5gOgu+ob5J6iCJxs19qXwtSox/lilm19uK6pg/mCbn1G9dBLZwg6BBjwky/
mGeZLzbCXKAgT9mMCXqyQyB3ACf6NmbwyU+5AHnlTysYadA1Eehh+IKv7paBM9mFut8gVHEK3z86
0QgIksX+hjiY1oOGctdvPdXmyli0L9o0+tdU6rTIqMge/7j5ouYu3FO9CI93o/BbNHF3FedvkIx7
ir+a02b8X1FqUysu0yBs81arnc5PVhn/fXnjAspSU0Q/yx80OS72OE7RhEu6jjJj6AYW+agPSoea
xVmqcITGDD8KHsc6nB7knAkF09qJy81dmndf+tDz6epp5+uerJAJgXfW/TRfSIUNjdpaQM1OmS8v
/GQ6BWEd5mquLwWbLEyhxlVr5q/bS/rB5R9LTUmPFECFs0eCz87NMLfr09kQAlFOCiDQQUZ7M8F2
vgepiaFq6dY72dGD/kvGoYJ/7AMmQ34yEp7qTHVn+NsFcGqJHMlvmtaSqs0gkN4ZoBSgiqIpbj2h
SB+mk8awGMjOHeZuc8a5ekWLV8kQdhQZP5WIuRZjUZeiBbyhJLsaYC1HSlsJHKdqX6iLQVTF1TDG
evXvZjtdhsWeeCTgC2g9sXK8PClJ/LgdqR39/V5LTU88NCEvuWPGPov59juyfaHspJSsLZEL1Xrt
1q0Pgf+pEjrtRy0G65qvCj0TXZyRP254o3ox14xxlFmwiudAjA1jH0YKauhzHyDBv+7DkQebndOR
AIgQJnQ5YNXGq5tABTQ4Alty1ysVZIBxkWxTXR3l8PBjPvxfXPiC0WWAfJXcc5s7StDOQqQa5uKf
vm0EbWg613MG4KWV4pjzAd/jsuMeH4tLrjgXnAGpyPBxQtS2uH8w50M2zC52l0pPhjSe6uodS+Zo
OVyVMW3V4cO8dz3NG5/7K9VnPkDYKuM/m/Fj7Ll7wEqHjbzSCYHOrUYJ5fX5rkZ1p2d1elwwXngQ
ynUxrsFxCnolMF6bODrWBhbAU9t8ndKAwBs/vGTSlFOvP6IswB/89sQrrqGKUnR5ND+oPrNIklce
a26ixQjO2JEWD9vIcWiqvyD8ggssG71jCd6nQRx4wLoc3V/ox+xyrDVL3WDqwdQdd06lhquIH+MF
6R6aWAMVtgMvifN8lZ9IRCYhf7W3cqnink8gxHb6Y3O7xSkfHUDRwK1pWa5f59EX48D5TZrn6lyR
IcZ/xQfo58Eqpb2kAop4aqkgsEs6/Jd3aqAbDEvUvRn8CSkUL7VwAbBmEgjTdnXuZ2CpvDki1ce5
WZt3GCHHM2sogLANM5M5RjReAyYKWcbcEF82/y9UNSAXdQStMm1OZoPYiPF32a6ol8LFKqhew1Hc
190VnBcfgRAuUcX2hHNTzH9ONdCu/OUmnOx4IiBQ3lh6CJKemmWW/lqFKokJR3nv0ocielMhYXA+
6PGbCyBLpBRq75vbclgYjFVSLMgBSgWISYTsfbxv8LGpHwFuQR6pBN4tTkCHTVgQ37pHa2rkYu50
nXqBHh77sYJ4BcxQwe0nKD0PG3KTnaNah+poIFb9AcHFXgBa7z0tX9O+ky4jU8T3jA4dcIZhpia5
uARB0E+bkahjCKPP7ODkrLUOaGFPPJQm4cdcweI+0xGWxVgL9aMNh435YCZxk/BlFhji+6ath8k6
jxR7QNT9QoEHEYxDcbooqCVmUJ3ESqzFAvjhMWcMHBVJ2K6R9+7sGeIYfP5KCz6tDtKqfhfJwArq
CeiGxGt+tE71eaCIZ4Vq06+lnqLtHAh76100WZL18lVJEQpG8GIUpT77xKQek0N0B/geyzF9uQkt
4OMx3Q2iQgcBK0LwIxkMQhxgIRMR6GsnwA59UczBYlxUQhnr0b38Fe+G0fIagaoyYYbxoyePgll8
h6XLoPfPrNN7t7EV7fjHUCw6MTTIrwt9bXDI/8J7yTSrZPjvMCUAyIRSBpuZhzOj+kchtjgqPlvd
E80yIUThtfubzj/JCYqXWMasbWK9Sh5xyWKuaxm/CJgZP2FifHSnLHpwIOFJksOc6Fe/pNFhgv+3
IkFq23ABReP9Z7RqnJn7Za5Jt2kaXkBu1iTuNepH49CbTyEWLMNUxPAHUmA+83IC9yTkN1qh7PaI
Epuj2+Jk01fvT/+Eu1Bjoi9GXMsMVm6sQNBzStGnTquqOKCQ7j5ie+W/HrVBn8HqeLCElGZ2MXCi
eOKl4Wix4ZtXNyW9IVdXG3umYfg9ES8VeJPgvWHRp5Cqlm8lgyMVjuuTBVvHKKoZLb+4n13hDsZo
BDSlJC3HtWwwYvi2l3ud1E/W/1/F0Hom5iLd2AKXZaQotSHJ8XjFIvnv+oFksREWH2sF7+Yzt4nt
gWlwObvL5Rhi1OypsqSfWL9hhbdgFEXOroP/BsYT90iFlds71zcH5bg+6LsORAlc2doxb2k8qMGe
nPP6E2mnIYeecURWwAo12QroMHTgc2TFNA1AE+Q+PSgsoJLCWY7vrFcTYbWFEnFWR5yQOepMD81n
WjJvu+CBNRfVcFj02zadYr2rhug0s9aGyqvvSea1IbbRpbc9lZMqAfxqI6v13LDCDTJ0nVfUWHb/
limIpSq1CrY3H8Dmfa9cYRu0/s0Tu3dlC2Z387gkt86j9GKjJJYdYIvJd/L9Yr5DOfcOQG8bBbJG
GRoQ+i6V3tCGEaWq523INv68sy4N0apoU+ftCTLItac4tlb9WrVxTtn0/zZ0tnaPWqaBDQVVPiRC
On66K/gaCqhM0umcl3rb70y1tKkJBfqBaNDmKM+S+9otgv1nhpv3c7XK831fwzpPh5lmlcUp0RIn
yfB47h14RaCpEmkgGvV1Wr8x/V26xHpVclb03V+QzOCahTtIgKzyZ76KqPPanJ3tIKnQ+LN6Ni+v
/lzFAuDZ2d+99sEbui+7C0Fkw5txVUCawlDv9obH6TkWT+Bl/tRGhdWqgPme9DQFS8klB+HQA82r
qRrWXa0U/NMWnzVGvqaXq2jcpTsf+rr4XK7s63bY5w7oAomSpfQXs8MtSXLUXIYKtXyl4hcpPyMi
GD5Z7QQW5Ltb2wt2htfDJLJX1WuDyd6MLioDa7ptzrIz1+WcezYOLpdfw8oVzVmUb/AcO3MLkknz
OAIQk85JBG+scpoYE2Xf91w6BwPSG+F4R+40pdIKplyZA+FrkWudSTnXOv7c+VnnYfGrT9cbem9L
v2j7ZrRoytgHX66q3RCX470jiDoyGxCFpVGcXhGKQGK+OzndvBi7HntggL+hi1x5TMn0xpUJfHyG
cZ3dOjdbUci8BFPVbx9TKIOKgTgJwzbZPOV1nE+NTaXkW0eJ+fAQoHAR9MkbyoqJVdii/+bPeThh
4OBC5s6JYIQ+/cH3f5GOZEDe15/Nq/ozAZX8f/l4UtqySKsfjyxwjDv/ub/WsZx2d8LONCkxghJF
FzQtmvkN5tHBhvLzIfXJG+MqhBu2pwCqaCA40RFDowu0ycuu73lU83TzO+m5YLmNhzQU8uUhslwk
qlacqYsqKuFEWfoSyOkRYFB/H4r+3vPLjnMOYwPy7MXpu6VhhjnbT8f+OqOCBbdLtZhOwlKadt+M
ig5KdDrHvvHcPMmUzyB6D5JtwyMUUAMk6cQGE24rFBbrOXnylHN0Gid6QJUwaG2B06ASK8rdm9BW
fDh7jGZsUJabtewkpGtGJihOtpCpBI8o5XEbVYyk+m9An9ZH7HNQ81f0copDmOE8VZim9BaV3DuM
tY/DpiA9ZsuK8gzUhSRVZ3i+K6hFM2o1ZIcqw1/5lYNP4n5gm1HJ7JVhSJ6YD2mthl+44adzMIQr
S0hqMmrmzNnj98SmDxGzYAhBorbVxQYumvegWVRrEvKEllEDKTyiviintSiAD7FjDOxnTPlradTt
jmPk2csdyxDKPEKjt7eQ5Otvsm4skPPZXTeBs6TNuqwZxkNvwctT068oRX/kUXbJ5fxd5Xxc3s3Z
aFbA9QFZrbcMy1W87hIx5pgXqq9OEvYxvhq2M6X4pmmR0p27RxErOvthJc7VH16l9rHqNrb4gG3G
gBfJHL8YxrdANhYnU4wpjyg5DAZJf7+5SAPv+ydYpSg7X2aMIpOeUWB33Rydw0J7nZLh2ItIDx5a
Y3124sp7ctusHaDQAumzKjv+MsT0HKJemOoWuC59iQzwtuSDWL6BvFwahgH0IiCcIGoaJCgJHZgV
Nfaxt1XQrn3Bzl2c+uiRUDeABoSxHDdDPWyRWipQiHiRnbGI2Ssia3B5TYOvuxZKpQPI8/9FYSrs
MO0I9q6Xyhxe1J9QheY5o1XuavPqTtE/npSi7+/Opqxnx9nTMfxyQwPTdkyyVBUtRaCX57UmcpfC
+/dJUHeIXpDlYRdkSykgN3NUg/KnYA92dqHjHM4FxZz9+ShUJSlNOWaXmbShINLsB/JZgEzaxM5g
Q2S5drhPHqGVrEBf3s3nyD7NUrgLxJrpT+S3/nhVOaFJXNKpItWgiDy7C6KriuNkvUzwzN4az4aj
p5IZF1/Ggk5/mSNGOho8BI7H5iBoNSyXcSvIci/MtDSbJwMNZaDdGyorljUJauTA/4eUMv8WIkSY
NjZE0YHI9gF0cT+KQjrZ0UjipgaufiX1vJrmPrkAndd68FKIU4XH0ANK8+z4D8z7TTh2fzla+6/u
ZXlwgxYJ8tzCKE+qSwPyJArdDRNwrMuxvEzCnzUKw2UklFEalY3Ai1d4yhHyhRU5GSYvrZ4SAtlc
nMXhAalFz5cfE3J8qw1nGb++0O+hSyOCDrU+/m11UCKwk4bN8bxaYzJFmmPmxsoRkDyI1UCyVAea
LMXnq3m8OxGz+Pf9HlSoq7EPX48YtcSXLALuIEjBU4HHM9jeBqGaW0HGJeYTb6HAWkrjdKjIKElc
y7FzLtrpwlwf75+R7/+Vp0bAuVoVZUJqpE0l0KWvsn21s3civjXnI5+Y+hdiCJRZF6zjSTEI4Bpp
hLGKyD16C0W0Zps2MavkRxWmGGLWJXaTdT8ow2RfAKHBZ6B8Z3ygIRgT75We41nkJNdZe22WCa5W
yJIKGt+uGTkqy9jDSwWbWGnDvJFALnnC8Vy9UEYg+Citg2h+f1kZOGMBB0XdSql2BNnguoodu2/X
0XyZJXzo+aXpoUSnoEmFTGxNEg7xhKQn2mef2UxjoVQzy+7T42QrJDluGEQ8phVaWdIH6fdPaq66
bbiEDZEdPoJAKpz7rfLdh3e6eN4parTlfY6kfpMLbJqZTNEW4JOpeIIqdq2ceTCE69xiVydRSnQF
SvgkCh13x52mKs0dRBzqt/dRct+g1COqrPuO96JDlAh3lubby+0pYMYEtPcQT9Gq1vAr/xbpglAp
xIAg41VbsDlmALnm5a7EGK2R5Dt7kcVVDX7wMnkxMYpS8gv+qlMw5+ZmHXVXsRNqfgzTAFd5Aes3
+3AIegKiRSJ5uHhk/xfWaSFYHaBEUCvc/CLjDJbPwWrhiTtbyrit0+0Am5GztjgXw9BchR8mm3/g
qNqvo4PX1YC3bAAvE8k1G0p+9TBdwqJWWNxOKbY0ixflmHh7eBRRsnv8+8AzrBfGoeYD0UQWeeg3
PcYP3H5tWPEiBwNZaFCONGtbLCeMJB1q7LGCeF5O7QFzUQfzRQrUd/AzZjNwgwjF5mEpGFkJST1b
KIv15cG4UufNioMhC7rrxGH5zwd9wQzC73HwGd2CyILdVgtaCcMbF/E/0bG2B3Vll0IymWxBr4no
YV3ZtbfkIUyJkauX7+8OyzGAwvz4r8PcGlGN9QE4tKWyp/kFeM0s2uGdetrAL2vgT/2Jp/5KWPsj
jMAjuN04XuKgqfaQ5zbL2FYAI5TS6pDwQLxj0cf6Q7qWEGrGVBQyGYNmkjyXYru3lK1kaZ6m3IrD
AZOhR2AD1De0eSlTVyL8r8aXGur897Qn9rha72tML8iJud4wIxm3u9p+eqs0sdBb9LjaaaZhCiL+
ZUgCSPdKrrBkHoz4GcJVazqb9mCPES27FFDBXuDmTPwZfT76jo3zlxPHjD0NMvbJS7Ot1F9EyRKd
9cDMX8Azuvl/fdrLFmcKFtqtlEf65N55smhwB9Op2qbNYrGFr2EsQVA6dtf9ozgEgJOLIPcp2pb3
yjDyXPB2dE+sOVr3RStn4An0HQHWMJCPQxVc9XXV4QCvTBZnniohF2fK3b4Gkd8eQ3QwIiw/Crsy
q5BqlxMOKvMIkjoPJOU7lJC6PYctrBWAVyO50sN6RggPyPQjtug5dn+tOyZ4DOzwW/QDwawaMVqF
WT7rGyLo/50TNdadte9SLC45v4fXFNDCd3rOZaXGKvNSrgAaHMU6jgLE5v1Nx6mrDjqSv6iXeqT5
oIKNVMgsiFOKs4upyrxDhGIqYKTrj+QwpCUSB+HnuIkseLAFHDCYXt9XAW5/LN1YvJX4t17ZAsY3
XUHN8SRmLujFAbSIwcw/w9Zozk1A789GkFClQQxoAKesxTU3ju4l0/VvBc7HaoQDGSHuTTxSR4ex
YuEXOoYVvuPwTEbTpmvwdy995hpqNS83PyCatm1d9r1gxhHgB00k0unP+VF2erRgsB9q/OTGrk9n
PV2SfqqvAXrKWGEAHCC+TzkbulqxB8rYDotTNC1+YncXdjIijAcDO3nQ8Tmali8B4E85o8WOV6Yb
1Qx+mSlHODGqZC3scOXiYxG08nMPsWHKrigsvPxiQnxUWuk9rSJ/VIeAqel2W9hhdxQHmy0KF7YB
XEt73S51Dhy/mYp6GK36pN96PPjkQkvbW3IAieOnKkAYrGZlT5z0wJQtozZ0TA1vyW7fXQ5R7kJE
z74gj3fiybGsyGcKEMxmh56Pwo91alD4dAikt1PJwIE4EJ9FryWKmHyOXb1KOdQa9cELlUsSGt49
iMfdVk4rR2MAwUVwfcTq+bJUbdl1FyK28qokmQEV5x3m7n5tbySr27EHHKpnnmmHVv4pEncE1NAU
3mOqaY0gKTKfnRjV48Z8DDpDIlR6pBp9FWWlbek5BpYITor74moNJAlf5RxTXxdQIUeNdtWbztXg
wetHwG9+7ei72IQT/FFlvDhQoGYS+ir/pG6AwxJf3rf0aW+jzjeqQ9vt21nyLLjTm6yTB/yX39dY
1pwAowdSn5MUjYsE8Sf/aabvPMNXpq20jI1DHHsQzTmO7swCp9BWWkx2H+BLBUICXUMBu3K0u+r6
JNo7HRzxAM8gxZy3QH3ko06KO/uDWNEkN7H5AXq3USsAWh6RJ0jE9h/EB+l57awnPkoDqgBQzmU8
kmI7lzHKtSn2em99qL65zC0R7tFxHbUdn7O2jA9ZCSB05/6M7uJ39fUQT/dNa8N9zQ0+Ur+XL4X3
dcRBB3tDGrfT+i8+C7OBws5nREK7pVuTqUY+GWFZ1cJbxakfXA4iYfw3MajVF0P5jTDUsR1R0SD1
E2KZbKxgQlJv5dm6X3qxgK1hIaz0l/4SBV1jFAuO7v3eF1DpOyUlE0v3ra2MjiccukZHUrxZ5E4x
T2thnD2i+1EnfViKzPX4gLd7tvDv49oYDjhcYifqHid9BtlI/ptrY7RitwkSWzwwTnzIpfRnBWpN
yJ3tNlG5zTcZvonW/S30/i5NkoZCVj1DjkFSo0Cpa9JvfFaGmQPxPM2/LqkENARJT3TvBbacILrN
/ta81XJeXf2UiCVbSe4feDBQbLVgN/DZU15IxBboD6xaQ2UQ8M+nOW8I2RvPPMeXxCkB9DXRvGjm
Tuc10m7kdqzjZ0PTApZ+nRt4jvwTrmy50ExYE4AC+9rmNbtOHeXGp6n0X84JKWU4mkq0ieBlNvrh
B3DzdeHlIUtv6+Fw8/4CwoHsXU0YUkceMiXYL9n/g1nx3zBMEL447CGKEiZL8HHQAkiWt/d+qOQi
qwZbxCF4uu5sJg378CnK8nd1+xmg2jl0kymCXFayXAxKtazzpbuazsftdaDYaR4xmN2UndqTFPVj
ZyqcL5Tw+ire9A+dvUbH/6Kcmiwdfixd8FTkYAwbUI/vYDp/fRQyJBprfatr5SqBHPt4Opt5VEM4
rK72wF2iO1w31mUMtBia2Rn+8FFh3LKkQk1zd3d+HTJHEEKmlI0JsR4rumixGUeIzCg028nVpSQy
AOXQBlDBmkFCJe4LzS0/RyI7ApGWnUS1NUDPKRO7BY5aXG9PzvI8c+4MdE+LP76twGiyN8dxtj3m
jJezeeJKVcNjdVgHtL75AxxKMH00bXWptTBT+GTfQ2Jf1xAP1AOtr3hvt9bwBybxDIzraEDPgKtl
zJ22wjWKlKNdLZ0KjLH4tWJ231Vq0sL4z6BjDmx1GrrNtL5T7l4V0yuaQmXJv4teZ1J/2Qz6SX8M
Ur5mkwjzqYpWWSdJgU6MEovXlqyNO887UrfwasmlTPg/RF1gKnefBD1mL0qAPQEKQHNDUlsxHazB
0ZFLCpb3YeKtaeCqYRhojuRR4LX7kZl//3AIAyAP2zheDfuJOiNYPzopwFCIxO8Yn9dOmLcnqUSd
JA8UlJFPZVu2KSNDQ3T64x2wGWaBCae+kO/31nldvrrU032MAU9kMdXDY5IH+F+jBhjSQzXePBkF
EZThOdnTaSrbCeEa5yBC/Zj7Yx1sUvbWIilDWjXYq9C82jJ9Amo0JywSkUeRwb+SIpeTb5Rnzdw0
dyDqp9TcvBJa/rxB4dmcEFX152ZQJI2NHVMFv5uD+oKTFvmwwjj0eNIZ1lF46TGQX+mHo1UuG8F3
b5ug955OPCN6gx9u9vNDDz96QH2BrA5ZcjBv3qo0R653wuYUIVExyv1WQaLHvHwl6FbMmP2eLA/k
LCrM4j6wNQ2LTpcijFv6bAo1H5JmV3oTU6A1Val5rdC4rMu0aT6lVLdNjpDhBPgJx7NMh4XbfDGb
5OMi129EPgvcSVHN/8tJmzvY384PCreL3VfV+NHKr4HXFpuNKHpopFlVZBIdpjqqmEYWdQGqeLkg
vA5o7ZssT2h+uFyCc0Nnthdd/fyP7aAzfPiO8ApfZBaNa6NN5Y06DdNHUkpXZg4RdPS7bibi6/I0
T+elzsU9fs/6y8mN0i2YRfJDzA8qWYA+AaHHNbsxlv9wGot83q0JRLumpKRsUGejwLnl/yr5s3vQ
6Ab/ocyBrVTagyQehgOjoKchV1qAamP44F5/xdWFA2cORtktFlxZlqyiD1qO0S0rzOAn1oS8LKSK
8g6zTChKJIko4/jxPsvXfGFq09Vnw+LohQ/MS0Qzv1KRKj/4Hn9anXEcH8USynjCOJpWSlbmi4Ll
FRgMDWQCghMCXmJi+T6QB06m7UEaTyOiOE8vAfM9MoHfQlR8wtC14slKIsoEyEtsDpP8jnDtCLMz
43u5doBIiAcCIlFntdGeGAQD4i5Ulz/OAIajkZeRIMdNM7f8c5oVay7Ab1pUy+5VE9y37fh1tXb/
iagy/Q5V0CRqfVbx8brfTWWeSbcBPpprQiBLXuGSWe5q4RkrBnQsgcrw7lpS8nyp+s5vvA148ocy
wPSqVkjpC6UxaGfH7hwInsuG6Y429vfhfgcNLQjbZ9eiBzsQN25nC1HJh8d/j3oPZckZEEXKCxXj
+tZlDee7iiMuQdu0oofGFdm7FQ4SvQveyig0DyBqWFY0Ylw2ZUL431+cD2IR1MNusYxaHhvpqh5F
7TARM/xw5V8lt3P+srw4cK/+EqDZ2H3OGLxmzpBOtVSnNTjNQtIXx9WUs9T3M3wUtov+WZvW9tPr
yEcUpe1oEaPoJyaRoJjDelJZGseEYJq+D8r/ff3IHgkYyOKhgvotjOXiAZLrum3pyVk1IyvHfofL
elzcbu0j52O35ATEtQ6mOTymnNia1Zjr5+WDrJ24Kx+2OrVVicq5Vm+Qdu86awrleqMpSp6LFDzf
Q8ussO4wuX2MF3qo/6oW+ZrUmExFkjvHQXNp0uIwvWSYQHeu6BeRb+n6iWXyyg1VlbGcTACCwNzC
eHkjPdsK2pqC3cECLA4F8gS7xrzr3IfYKVSJBkHAGHFcQlAtvJw19fCYeFLGiPKygXg22930xyAj
/v9bLcUg/Di3xc3GfyKVOGLTyI/mhivra0KCLfZ8X+5tGwBPEHC1vSjc7yOEbSXsAwLWg9ovC8Kw
YczN5VOZaPFMT9HjOh2UWa+fcld8YJ2ij1dC0Yh2xmBiIKbgcsKXwShMvtHGiNA+/fWjTM/K7RBR
feDJ9ETb52ZAszw5E0r67Oqx9WhXXxv6OieVwOh1EKdOVxxjmLNSyg5Vvt7g6fq43L1bG21CovPQ
cMZtjUEX6NRcbLBhlganG8RQE4+gh93rBt2L9rSiJYpVMeEXJLLlSAEmXoIq5Z/yWTRqRp+BdJI1
ClxnXcVkBSBd6ZQpOy0Q3Fjttg+n9XVEk3KhYSqFP59RC33NcZtfW4CMQ7XmcomJSGgBs0Qa4A2W
CQ+4dwY2C9udEyUPo/Gv8aegoRemFVqinl5rKOjKu37dJUb8/yIYwqG4CmVAXRpEl3a5hh2jLCu9
SoLJLbq9FKAr9kWqd1zcqRAwUkoU7xe4fZLmAV+VrGHAw1tTCL2gtgOlVMoVjIxvFN5BjgiS3HWt
R/10gKdYdpOFBiA0blKD+ULzeEacx+GnqNognyKkFG8+IlH+AWNjvzJoO1xbQDCoQ5VbU8Pz8L/Q
IXW8aYTpWqWfq2+CwY4PFuRVgocq6Et5tgZjtqpPKAOCI0LFOKjW4YORH7nZJ19CRS/C3rRTAjJ5
gx+c31f3c5+dOl0SRSqz+4MWGCqzhArVs5lJO3SuIIM0GZBPiNULAX2qDMbR9cLWer0gCjX02fD3
u+G9CVG/uCmKBKWtoLRALm5p/neHY7SZTr//MidTpfAbl+bE2/KMzFF2reW/J/GngiSaXnZuZcgw
haHDK0c5u0H/EDZuqRDZShkUgG2LRVPgVcZphp4L2y2ddj5lg5blNPIrNZGHtVVyKRLZs4v6HQFx
gway5m8DLrADXgd7Ut+vOIbMvUJqAsJ55fUXjhPxWwAh2ctWJ9s/RdamcoUSPz/RjlnArG2s1+5o
ZkiVy1cH7LQk8pO1lWCemekBluej+F9XmJ6zxkzw4VodNLtDL+wMjuHh72spIY9AwJWl/3Idqbwv
+TQwKYDfZGWSmCjpy7RloYgTDFnKzk/vP0CgovdNC10mB8F/vDMp+vvNst2g/zsw7sQBKFnJ6zI/
v4JkE0OWO+RlKQvlEW6sdLU8RIUzFaDgp7g+NSXjxvksf1PgoKeubBjcEBy5JZ/FNUxaVeYRc88V
lJxAgC9oOwznxD5+mKRbP9Golyp5zgktsVniYIzYWPGyhXOfttDGcuqCXKlhGYShoI46An5h/Z8e
ZtAE9lj5kptkgNrgvjOXsZ/pCGHCNz63kn6tnWa54NyZmZDNdGsDJsigp6YVeO/dC5O8yzyJFqMg
sSK1dbFct6LJjvznIWroiaQPlDxh/Hoj02f1U0MjWtREuZbYYnSAPE4DtQ/TCF2SWeSkI+wTgkv4
KLDtnpKIPn+WbOfAfYGOwIYZE6HVRCQUt6xXd9lA8yHf4F4/QJxRg6EbVkFJTLZShorFXbwm2M4x
7jxIlj0OFhxawZh0KoKChXArzRU14qUQg2ZaUmKWPqZPA9uSuJih4HdkDqiCgu7KlJDTlKAn0O5l
FEiC68tS8L7ZrN/TpGUwsXGVoa0k0eVWfot1GbIPgVT56OaJae2omKiyZKQlLhbz06fODvqRDa32
tEAezcFrKosT9zg01/TrRo2Ah9n4duL5EXLi7PIWAhivVFFB5zNDJlQZlFDqkA795jVfkMCQ7hBM
vvdkzs8H5knaaY+XfchH6NjanIBXP4+OMF/0AYlFwy+Xs6hkubf18Q/TvidKGM/rlpUNP4BJ19ce
N96auyzQOtjWXAqK9CN2n2mo9DdOlX0+Bwea4bTVQXcWAtyLM2PCjx8K9otZqKT5Ut98T0geGozQ
uZs6m5k2fnJzokOhHE3QIMsxKEqeuPVJh4SchfB5C0PWJBCBxfjRbhgjXNzwT/C79aW/QBkcdbHE
fXEeSVE/HFwa6pefxUeSh40uvioAZrLw8VkSsY32TMv0GBNaMbBcTBZ2VBnUGSaCUQI367BSKv+s
8GwgeSDvNtDBfGivQ02DW7/mI20kOUgkLZn89gedlLJDDphH19ncyQB7wgP9XaXTI+ngE1C4GFe7
eK9MjXJUP7SyhOsmB3ZtJjylxp3bGx7vgxjM/CEUcXCTyjQsPC3Oni24sFxkaXcnj6I5ySNc14Lc
oszIM44f+xdqpqCxP/JxzuDbOESlQRXOw4fBD+jgCaxgFYVZPIp9UOtf/hcHS4nPJfkZPSEhI3RB
qmm9ndFuVPxrwzKheVwISCj9df0ztek8yVp/mOw7vFQ+tJq/Ar1xyYUKrxImSWB1vQ+NVHqEaBcM
+STHi3LZmnw7S09SZ5WLjKuGOLoXPjx5wn9+QdO0ymkwSYj173nzeMjcwqSCXMx/ZdqS/4JK5VUb
f1XP9L76NlL8mHnEvlfZPhvbPsouP8hQLphGUn8zkGP6JSk50HeUzkeEAjm9NvuzPBMPrxzq1tBB
SyPj0U+7xDXtNrGOhBWZKGrIIhRBsSqk70RxVgKM8LCwgl4dfqXAj0HTycXQdHvaFoQTYTtuA3vG
lfFBe7ddp3/kJpDttV3KwF6Dlm4KcrqO26lMaoO5AyUQIyixKzQy7DcU65TrEE9r6PKAelJzP1lD
uSxY3xw/ZwczxymJmG9oFgG4b8cHUmDalQ43VPHoHWflb1X0s1g6myD+8iO6dc3k6EVcUiERU7f6
bRfPLj1o0jJKz+Ndso4Rei8lQIukbVs66qn/QKt5gCYKgknZZmKUAFCniMDIRLi9nOAJSo+8eEkO
Yfct4vx6UHBLfcrhH4z353yPx0m5uKJnU3zoCGdOJhhC2WILxmZ7JB3Phi7U6fSJb+UkK9g/hugg
ezyC9luhrnXxoqV6RdqV8/ALFPGUHcUmtICkBQ3gFXI7CUrMxVOK8DpGjv7XcNW85edOUea0IrMI
a5R4yCVqEPaae7a5aID9SZ19M5u1wYfDtdQxfHmbQT3kOvqkdQLPYEdRbJAKuLWth80lxL8cW0VA
Sqe+OAb6K8GCWLRokCmwmAdHtmEEYLOpwrBgfQDFj2QxjPT8UFHIAa6U45nQKZcahkHJr2EmTwYb
WcGy7hSEPsljyEx2RRiHqMNV67qF8CpAhnfLZCYYHBRxrvkjlHBk8MYJ8h8lhlthQ3Iagk7ZEjIN
kirpMBhH/acTymZAklofyCLsenBmiuXwTD8XClE0Pn7hidWgkXSuhoh9JD8udU3a27J17z3BdX1Y
ZfDX4De/gZdK5LishhJKTq4XOU99wHTwwnD8RRH5OI5rP0RzqL70e0F764rRFwUDe49BjLlIBMp7
NCSp68luPVJynBRNs7yUKgqedHEX01mQAyXUKTbr7GCX9v3VG91Ay/tx+nknoz+rQvh2FzlMTiM8
IoN/QnR57jmNX6frdqPNdDEp6q8v2Tz4WHN49cg0YnpFuCOivaXQU139Na8O6I/y8IKYK9z9FbRe
DDbRUJf19WHUq6a0wCllgPDuf4AeGrbUj2ct9LaU5+TOphsmwKSntcl+gSVex/xjXo4Ku648Xkv/
Kp4GaY4xkmXve6hZ9sbpJyQQzQ2pS/+S54y035Mjif0t3wD9c/PIbfOTErwb2kG9rT9rxrk4d3IH
czIXLWhLtx8xJrqEG+qw6UaUypUP8oz6SKPpN2Hm2CIda83kvXkbk6UVjS33zCGV4dfGhseF7Kin
9yM7LjNRugXPjLbcGomeEbdBbOxnj+m5yM/mKp7WKqL1vE8T2T3GOF5dzY4PhUymIbY0C9qn6Plv
sSA6CaXTKZCXeq3AT91ltX/9XWR6dFW3BNglHpqEGl0vVLAKyfBUZerPqO0ysb7Il3d0uVifG2yW
13obYp24KFLZ7zXiV2cx+pn9YZ3TMvVsr6dD3iCQJWqlldSfvCyQLa6XndclL67IsAV962nm9UPk
eE0/XQaU0eygalpS0AFPjW1u0kNSlQyfbGhfO9o+qWzMsawrVuhe8xPj0PiV421MyX9+DqvwSSCm
3nkc1VUh69Ew8n1sRhTHJuWgDx/quClnh24NKnMkMgo91d7vLeY50ZLLo2ND4R2vqWtjqF0KQEa5
8lasRIEwTUGmAGcZ3LIW+pi/NTxFPcDFrSzNiayBgomCA/YfdPx3In4ANtJbMPMR7yYRF1GskoNC
zyYhcEvkiDtMAGlskr+J6L0gEiENSjP0OSHKL9IDvrOCPC3FGGIt58V3tKupDnwEQZMrVc0f1yiP
44GXtp7HmpQwOg+wf6MAll/wFygBCUBf05vq3mzZH+ahrHOIUXK4flZk52QVfS/aAHzAlOtT3e15
LwScVxG8r0mVFOx34H5nEJwFtn4p1RyMpK6waWAOobSSOKKjByn7rsO7CrIuSR3m6XOaN5LzhCyX
wGs9e4ye5yMTT93y8p4dPqGgOluP61HlSBf/m+nChLqd4/DwXp8PE+DJacvYQR6kw7iHZcpAYSxd
f1YixuCHUaNxTuhTF+ynxCwNUShn6u+B0q5F5a918IHoyP+uy+EMv5mhu9HF8iBYqC0vWLh3njyu
trzeUoqAKz016K0mrCgO739h8SmgHNiANdvgUsU83qMi48Luq+K+mrmLTBoEHXB5HbzkOM6HxQtj
ceeABU6G9c4GpGQPW1mBQ5Ye8BOP9ueYSAOcFqA3NmsefYKJ3B6JF03lqQ7wY/5DX/UWcL/Jgwio
+MVz9i6m2AcZl+GnKHxSHhukhFQTlYSm6NqgIGB53dWhl72n7CHqS8rEhHs7SvNgmZpvuE2DhnTJ
/wg8mpDnN80YtRDY34ikkGLLZ1siTNPSCAX/uqHLFuNuVHDAk4rGNHjRfPjU4g3bqCcLjkquCfJW
IIe9IMjycasDL+O79dOQ6BXMpshAhr4Ajg2quDb0hmI+8sw0EVcbFbGILrv7sIVCQTnJuiiNwqhU
dNLj/9HGINNUOr9rMjv+68X7/2bkbVJGMRfc0P9UITYoib3QXPnjDV8pG7VVsmPqDQU7eT4U8QWZ
XDqMaN5Ten5xqeBbDenHSJZzZAgkWAk2ckbXvq5RUWDXyDultS7N6FwpO/F1sdLbpcEeh4V/b15K
qMo8oBUvyRnG5xD+RI2SSSTShdzTZIWj28PWaJBZfvBr/GuRF67kuaaJ4DXqAvuMdSwjc2ClhGLQ
pyO2CYrRE8KmmpoWdB48RshF4NIr8RGSfanGXvjU9M30NVBLD6NztRhCjovrsQ9IW5hCcMGZPj80
Qo5qt6ZlacnW7ZI2L5FnxA+NqC7BdzkmnrX9TvIqBkM2DRbBCSuIfnT+ljKxsGTePijuNhidT7wT
RxKCWJ25CCLllFQGGAFPrLNM9Srz6rBzlzYXkiMz0+k3B9NS69/RnzhW/xLLRti3BzKTar7ZQKTR
I5qU4+ElqTzyn57u6Euc3wdLexIiWqsBHDKqFgUWLxrd9n3H0y35FVhS0AEQQj1DkVj4sT84SfwE
dIPowb+KfYiSzhsRTItNAWnUmDE5YqvCtKaR/UZhFYwdHcCdjwkRperPbOxVV1dJc0ucxNptjua3
BBd4mJ6mvReoMdhi81eP6IMW7mitCC8siRt0JUAl9ddE1zMRaHPcmJiB/jZ6VEQz7/pJ7ZLn0jN4
DVlKPbn9hbiTFLOHtP805ASwWgF8y+VVCiTK8JIG/5nyoA/INtvKVEDr6aKzAly4HbtRpSmL+w6M
wFjDQ9C1r/acmiGFg+3QaaIppnxGT5wxYMhoBQWPv9Kq4C+esKiCny/8zLekTSDXJBWMdGXyfnr2
hR65pPScLAeLU9PyWIuBIte+/yTa/dzDBGhU1CYJsjmJFCv0oiSt+Rx9tKjSptEUpkZpHMV0MioJ
LMeF9wacnBEUxFv5G85Vd8SLWa6wBoiea+st32T5tWYsugqLqFgly8yxCLRZLHcKN4V6sFTUdDJZ
anVxExsROiBx89VaCJq20QYbxciwnOqXhdID05hlTO/Bv8SpphwHyZEKP+fuaRV0+KBays3UZvUG
pObiCUHuukvbHpo+269YMridbyGs7tec9Xbl2YkgI5SQTgE5nt0nbA0m4sOhE8dqnmVs/AHz6K0K
iAE8UP4hprJs1RxiMrig/lcMgZbAB9DZrOFxNk+jZOARNsF7qd6Fe7DZx9wWScm1hOmJwrn08LwN
x90U9Xgn7kkOl1dbE5RBa6Kg+OYpDWGcWfdMSxg3FdI3yj8Wk1ZHrCyY8o+0BWVgREdNqZDYbBqy
VyNVgbczD1M0EzV5kbYs0un622mfbSmi/mQfmQC8bLYpWaEINTIG9c6uCbrSZNHXqykeH1X5p9f1
SujXfqdFsRFtFojpDBHq9U8JeY/IFrdIfaObwOJbruUL32TSBU4P/qAPgFaMDHF/oSGITBVnDSpg
hvjpqr+WTphV794i0Q3CVIDvQniij0IjLX+cfm3FL/MEwZqLdDlhU+Ehmp05v5H5zh0RVM9vMpam
2hLsNWPk82aBA5BU7/Hz2CDKdy2SnGMXzMS/lh0LFFFf1WQfg6ltEE9w59473xqhXCJXTOevgqq1
bXCEV+Q7IF6SYD5T2/4bsaGY2FEHysOsjwYLex7HrArBGuUMMnF2VYpJLE1klWkrwIkdJQwvQD4u
xrD4fwLLBS2w0gUjYen0HY3R5aLoNSpkSa6zpKW92xDTdcArPnTiTvx+UecxeXhgT8FPduPcZPzO
lyK4KTc5C9huLmglZ30B0yI2DROTAdR0OS9U7zCsqXB+seKWQMck62pqcdkPRXWGESZLlEzN6rvH
IIdgkruZNzO+VXtZ6y/cgsRQqnKjpK9K8B8l11T+rmGY3un+ZZVWeR/OF4FD7Xno0raQyjhYq8H6
BzHvhEXMXh/40PDoWjhx1z0JjVKRQOs2OmqURU4P+ewq5nN5gzUBXi7qprdvfQVPIxUYwBQ14d33
2XPWITsK4ypPCgP2huAK7DZ6ZnBc6uptlQM9WE7X0D9//tlDn+oByrH4+I6X+OcFZziakSv9GJcn
gEEzVnDd92GzVT4dF5xeBGsB0g0R8cE108SjCzKXt118pOdIQ5tjKQwH0OZrBu207NIGthMLy8JE
zZFjGH68dUcErXgwTFdXadBotmgTn4sv4gCL9ZN41TgpYMZPShdq+CLPEnyLBQ23TnHUEQr21Ouz
YY2ffZmtw9EPC53iunw7FzxANZ475VS1Rs55/pd/Lb0ggCAYd0vaxfpBwvGIe7D5Ny+Dp7ovvIzP
LCzgfzOCNEY4d+UK/tox+km0HCdCtcR+ptw7tLBX2Y8lfMXbKOXjuxgYzWRyx7HstZZSgLI2w5k+
InnwNXDipfS8KbICuOpkpf4z7/WksE6dXeGS/5D93Fnlb4djd1q7rZBko1+xMChkWvhyc6HwEXyC
RWivNiXkaU4yyz97nxic9S4T1BcMhRzwGKar9G1MHWsumUkBvFvmCdfei998SWOKiBfEPPi21Ivw
4Fct3pH0+hDrpmZwfrPVZBkGFDs5nihZYJwjC8BT5XS9W125OhLHGvhCZnYa0bUtmJNEFBF+Vyeb
3ciw1nztQ+nLq3KZKsVnYlV8Wmj6SAoIKSRG9GG6gt83AaRzZM7ESdS5/618dTAKbYRPYqt6JDWX
88yqWcQni4L4QfAGD06nW5F9kRL8UBHYYHbnl4vELqdgNsyhdiuLQs6Tpxg1yGPy2vyfMsDUqxhv
ocaoFKXNw0KC16C7gbQchVsgqdX6O8wV2uaUWK2oHuCT/uogdY45UZknZT+RKAXhT/WoEWwLGqus
8sCKV7dX1Wa1mjGVh79M9vVaKsn2qjsPvU3INd9Vg/BpxJ1bBiYG3y64ItHu+q3VR9gpTVD5+zv4
bbjnmEKy1WVw/BGZZlROZ7WcCNX2h5CbVnJBE5Io6iY7i1xQlY5INGymqR89w06r9235VJAKy24j
wnjb0tpinFc1mVRTLT57ks8eQyJhIbXTM3HCamXzZ6IqDaHJhanFdcoTLz714dM3M9h1E+1RlwXj
aL94+2oBmA+JtfY4EALo++z/kKlwmfISIIQlWmH/t3DIlpzIDgsvyS6GLPQ7Vzn3kW3NBUP0g5Fe
Xd+E+X91SkHXkt9oiCu+DY72Av6f+zP2+E0ADNMKnTWOG/Q6jCvAsnVevNbhLuh3PPc71D0v4s30
h739aF42bKTnb0Owpr0YfdutW9YKhqw0vbFI7kiXTET5r7an5jjqEbPYTcjUrw4gbbGleb4jg85J
8LltGpPw2wjzE/9tst/9x4Oj5n3TEbT6R3IxYV+7No3309ZzkycCIlKcscSQxsWE6lfcOEDMFPhe
qCtje4U8WnbrDiGSlTJRIdb1hgfKIdxXrBL9Ng11Wdod7+5w/LnbmWtwzAKAf8YVqtwGyM7W6YF/
iQWqnRRZt77hYtq7CMTciMAoz8UcnBof/1VlK3I7uXDd8GUzaBNNFnnuelCZG+YRrm64i1T8VR/z
qfFnmMyl716p3zdTZGZFbKY4MgSwufSHBiWi458+sxo4s1wnVU1B1GjMILO1aUf4+m6CBKVBG1Cv
x4bo7OChGgPogMmDNlajUE8bzmwh6OgTpsPwj5NV0niAgD4LTe8jS1Vkkg0GnEhxfchsi03BVrpH
i7MTdhNuq1MDY9210o9OJaEIQyN7nZ+XYD0ex+SDlYrdRQZsCct0vplm87jx6wwJESJ8aihSDvDr
dWE0P2GBnnsToY32RK1D001rtaG7jNnX6pXdkWNSnc430JSsO4xCAVcVZXJ3JzbGRRKYtoM2JMOC
MX0pVvkg13alKkgnxB7nPcKrbWT4qQNJrJlRZu4A/9rU3PpaQgL167E3MlCE8n/aJ5aOTaAQ3Ui2
SOhH7IQNYdDG5bak8qdoikwuS6+F+Hz6qSXHAMjb/fFKzm5gB9A0wDfMoQfcxJ/G4kpT+OqQfuct
FTGp9SInnd6TDu5GY/HK4d9DhMHSfYyziUOyrUO/r1r3cluFJjWYYjaqRxrmvFoau3JuUVSt5x8J
I6Tpy5oZPrKe/7CIuLg9oB9bkrV/W+rMh0yUpFCy9HGvr1sTJtWLTQzXEK5/A0tAjppCh4MzQvSe
oVYXPQzV/b8vi8pSEuILYMK9PNr0pHKMSVNc4Xn8SpALLlACcmPUlqsf6hhFCL1T9HrzG35oc1d+
tIzoYWtS6Z6EkiMZwt21RjS1d5qXL+3e5ZPuayd1ktIP9Go02nfCmz/iiXP1pDz1sxdqqAmzEOli
ueMCb7du5ce8QtF2s5U7G2cuhYfZcI3EzDHCW+QgbsUOpsb85bwCV0fcVyZspJraniAVqwb/Iz49
UAS7OyymCkOOhveAE4Pp2W+96azCE+meVSZFujEt7Dd5WeMrKAas7Ye9fS/W0AmzS6ghhLKNd3uf
Tlw7CUfP9hrkU5fFBGWEEcu273TaaLBFbosXs61fgEPBxzOrVA7fDTNXnaLiFSIiC6ZjXDqvxg1S
eo25EA1BRxyYIIIesoLvjGy0L7tX9EPAlnaaQaWH0bVTWhPDR55wVFdOU5lf3+5yW8+Y/MJKSxYw
wRyuq+gDiEGOXEYzWAX8NkejWCixJtLRlTpqcNOBacA++6H7lvhb1dF8QN47GSpbMHQmzH1XLnsV
25H2GAZCpHNrfaqoUVYudWWBwd7aIvsiuzqkUjWLqr0CtLXnd1Is8eTbrcL6EW0ymwFnWWVb0sz1
nN5waMyErDaeyEfz+cRPWDoOCuwTvmEuAqLinCEeUBvvu5f+1l3ghLPGe6lwUkC6Ab9Hj97AtZ0e
bAoJBx2lWm7Y+iyCguYGDUQM4B93AXoltQn6JOXJK9Uc2S/gcthMxGrIJrms7ngPh4aeLlhSFtRS
iU/Pjgj4RJdhzKnuAecuY6aNob/SBQDPNKjWxHMbD45OLn0AgqZv1HhTS1S9crJeX/3Csmqh1Vss
gZ0HY3rmlPoxRYkgW8DgADHJ0hUdZc1IcZc+LLFVXrgJBvyDWjU80sUAX1HZKA68rvofsXpV3sn9
w4iYK0aLESKCEcZtCWAJ2E3NSpLIwY7/NRhE1zHXv1Su5Otq7rIriMJ/zWEhWUl3Lx2poBENcfkR
7qXzBK1DgYv7/Sgge8TR+BqxqAVwMzoaUFwCDjk1BLomKNKET6oX1vqiPCdZdwKgb33dFAU6RAyM
J69HkJhXuY8addg4qriVXJlrphqIE7a/Pz2V4n2B8RpuxDSbagDNId/wYTSsh70kTYr/AoWL4E2c
m8s+BhahTQ+VkLHTBJ8a9G+1cNW44dCtk2IEllY51a2pnNRSLdrE9FwUCocJKeTTYmi3IQ+fYkqF
XQL0gGckguvYNKZrXYWRzbIAQhh2nW25aw+qwk11GlxKdAiwP/2RkpHOcqDNq+OGbETn4for7C/l
RFyqz5viGUjwluip8qxSf4iSA93RDDQTpfYx0F1DEk8T2m1gDxftXEnNc0Ss3wqtjvdx00q/I+m6
mDhE7DVp5PC3NTTgQd+1OSQ3tERQyyhxj9wsQfWz/o3ODhFuam90HdXw6GO0sQRCHYW5lndAGpnv
tfPX3+Rm5mQ6xCFmCScoxjFCN/0A4C7+ParCevVz0SlzisGARwKpVzIQn+iVxysedI4F8VVpLRe4
tjlWXE41vHfEU4OvLsP0JVJFQT7/gyrVSfz17+xt+Rlr3DbTRgN0INeNHsjAZ/XuENZamsx7veg5
AcKjRlqfiT6pHeME5ufBFIu6ljuz8dgvlKnreGsCTQLqhJ4NAwT6BFzJDECKQ/Yuw2jMoIDiEbby
73KkOnK2x2lQVZR6KMYWiNE72vtSZiLFqyz95DCtw/+CfhiMv+5Y5sti2x6rxw9SII4HVxX2JHbc
J5vNsgMz443EK0cC2k5N7Fd8j6DsZlQfDSXQ/Srf2+fy9DSzxoz5ShLVrFKDhA8Y6DRxKMCNDcrR
c8APQAu5WlSHfdf3bnarMHdWCIuz8hytIVGxeQuUZ65sMLnpPfbAFpLaf/Mx8d+ROpCnyRAB05Ru
31x/AIFvic/bi61SB3V4Ubqb1ka4sRbgw8yD68+1go9WErf4THugksNJx25mZREvMe5QlTBG8Ute
dnFPcFqgfjOKBpC3Ii7X1lKZq1vT/h2r/WQhkdQFhCV5b0rdwxsjfon2gO5ne95dnLJmAcZikVfw
XdriyobavFwLztM/pMQDKzboGe/aQZzFTX+yAiiK+UMI8Er+X9CcRTcSK2XSpGanMezoSsiLIpZV
nfWla5IhlBXiDTJqcOaRV7amOklyujjNs1GTp1m+ZiBRFDSV4aO7fOkL7/9HDymYQ/kdjmKzkiFN
3aS/1r9J9GNwfWyG9d9fDs9qp5rXgI5xH0X50hUV16HXaL4ZlfyyIHgSA8StMGvN3Bf+jIBaQ9TS
xlbeOhv+1k3+by6HGaAGtDXj+1XnjXr/8fTt2NRUU2wj5Nj4VqIpSRTY+UAnN3tSZ3f+KCQI9KbC
2WF8bov6OXszcVnRBSUmfWQxyZIr12pVUKwN70jvjWPuSh0Si/7yI/hTRtOsNvN9vJDAhWd8eDNj
w/sU43Q5wbwj9u3uIVK/Pai/KSNXCDLzTtgKaLL3fZ44a5L7hF22Q7o1uBmFs2YBt074v+jcJPEy
y09U57De69hlqJd6RZRDWpJUVsTMouGx89JXJsXLf2s8KLnNUfA8N+yHh+VR8oKxsHVfSFWme6ez
3FdejJxlg+z4wjBB+DRaQnYlyEafe8GVqEdw6hEm7GGMxy+qdvAKoLPiWbFzBilR+kXTB1CHyp0A
vCvBRzo0ZME6tAT2xFztGUIqSE8vWSfIe9quVb0OIjultxp8r9pT77HYOjB3QpvDH14iE467PWQa
QyQtjETX2WRvXpgNDkpRbmlVFxY7ZU33lQFwDX/mCVf8Jc7i2jsPCn+jbUNqFSoX7ccjqONsJ77r
8TlAas1nNJ0jS5qUrYYo++Ip2ZH3ybQk773hcN7gNY5AYNc7zzTVZdC0I7x9jyWNsUX/cRyvOahq
VI8B7DyrpFVAa31hWegiiHO9oIt+us+CMGIwKP1YvsRmQW2ALEJWPFftUio/OqHquGTAPs/5CJj8
ZJSHWf6c9GrCwdMg9w0m/ZZsT/1c6cIbxAqMGs9219mv1Frzt0pU/a9Qu5wMSPX41iHOkszD0Hd5
+o/ia/dc+NQWloj53T2i1rFpSVYxkGKW0sRvsnIOQPLTd2/CXz/fqoW9BBeDhXcOqHx9VjQZHW6f
AqBq1jNVa8wfnJ7PDdg2ZTDlNqYYAbT04vvyNSM7ACbrtgbNCwjVjT1Ba+0jwCI/0NpHcTg8c1nc
pT9kAnlFKrCAL9AIkm58jaF/Qp/60Jc8XaUfL5Fo6PQzXykLwHytnxT+jkfBYs2qzgr04O/1wOuz
658gr7+7MOs6rHLwEzJCrYqeIGOZD0dxobPxgaHYH1Ci+NSIf01nM2AXZp0ULI9eAqbQP6Ry8dTC
k1rXzrUssqsQrbBBZB1o+xds28c+RrbskDRftZ8QX0bBcYPnOm0WUm9Q7dYZ4H2rmMZy0co2v4+o
x0uqcKFiv6JeBzRpOuBEvYXOu04vriJ1duWi56C7mhNsy99IUn7+o1oH4drdnPBnC0UZ4NkTUKpy
8GvdCdJSlAKbOe7jxAeOOwWAEBsXf4jcK42nO3CavmG95UxVbvWHGMcCtrc4m/xLtwF25ZNqWrYx
W9NAOqQ6CR+Oo6O6k/dxrFSSP/6AZUeouHeXOX9nJqQAMArISJCvUphzCXc7yC2tGM3IYs/CufIj
XAofDlXqMgJ7rngh+bBAWAziqzhsNruWS9VepB8vGY7KsPltkwpb210FxJSR0Nxv0/gNB48WlW8w
4VIarynH5zzW2LuBgYIh2H3H2lChRaRWi5UaMNzp1FBhBlnV2bZgwjBUfcwt0xyOEX8KyEZ22m45
Yrhg/hL1fz3b0BXmmuyXmSLR219PSlxX8NwryHJyk4CLOaR3jfkypWjMrsgSA+CJOyrw+1lScbEb
0atvLPpPXZMqVqrN2uUZTaOks456JjodE+yPr9VKdN6xKpSjGOjIbjgOLqBpO8lzTXK7QLjpYxvc
wnzHuPAJre6SWD91BoROeZV+t5fPyqZUkuvLqsMVJFl2sKGrwLNiMB8ETNesF8keXe+aYQeL88/H
9aAHvHIfjgSK6eqkbEq77Y7wiZaCXayQa1PEjLao8/BdyXDfeV/qxm8/BFTVp6E9fx7TZvsd+dR/
NYzzwuICtwXjaO1LaMc/SpI8LHmqXlH68sHmj2hJzL5qHIx8mnvWGTyuAAc0QUl3CgCxrnlHoVHn
JzTGRW1kmM6lOEK1C8ngE/WagE2EFzipMSgwuRjeROau4gAyt+qmGuXpA1jG9wDlIsgze+HZSNmM
wtPqLgoxY8gSZxhEyLmLpcxwTdTL1XGQC4NJzX89NJV/OPgBKUk06cMWb2YBP6zCSpkKiSWsgRJY
oriGMfgsL16Z0980rIq1ACWXcED3bdKZvlZg+OsnKohYCxO6A7N9u4jkjgAZ1iDnLIlrBu9ySNMx
NaReko/cXIdcD6EA8uG0i3kf3C5wImqPsrqaodlhNd818ZyA/DYP4uv5IB6N8pA4IkX1MXZc9fpK
hoeSSINMh5T9JzC0GX49ZWsqje+jnaOFldfGctszz94eH/Dp5S7jQ6R2y1nwMfGTEM9d9q77A0rA
pWLjF7b8r8TXjGVBnGsqbRd+C9PJxyZCtN1fqXNEGrVgUcQiYm6nLtQNM1RQpWY5u7OM4OJ7QRJu
LwX7KwUcCuUKj8zFX/uQZzcgtJNt+zTirotgB1ELmrksYIJo4jcg2bm47vMcK5Ril2bfPCPQBj5f
EWyq4FVx4FCrQGzEmu8jQRFa3ViZ7NBg7zjUjFV/8aZ2yis5pM0dFUfu/dFwaAm/62EjD+PsNeLe
4cke/AFrh7VMw1XBDISZbMcqCfl4zUcOL8UlriHg0VJi/i3ZCNbTXGQXekA0uaLOFMxcsw4NPzO2
qvC3Ymu8pcMjwV9ViLWnrs9Dj3pFmmoLVKklDeIwlEWAOwxv7w+rzpZAg/3m1sDhESX0D9gOYzai
2ruQZQXydDGDPv33nLCDsDmKKq/xA6vdQqeIqW2sUrOvnv6QtGIR0Sm+UHq91SLqlgLmPXW/5rJ9
gvUZj5Rg+6AAEn33BYI/zEYTq5s4400YPBeG7QcPZXrwb4KELNvdOvy7su/WnbHYkYpIOjrBpL9O
fM34OcB9Og2SJspLdqbIRdft5+pMQsTH/BT++itEDcs8MbE48VzM+aPJbP+2yLhGu2Z+Vm5Ktt9/
66y4xBmcQbgth9gZSxn9y/XbQTsCCF+c5cVvwDUpgQo1po2lQumIEsqz9XnwypUBUFLPMYZ/SJ1V
s/jlBP+6kqUYTVa973DZEcKUZeW6Qpn4QEbHdi4x4E72LfTzS0HnSCc4sm41pEjeE/42GFtvaLjy
z6MQa9DZWPYBCLXhLei1O7jLVkixIFmydo/ZVrxGQCGI76vKl0zlWteo0TCVXmFGYo2iSRqhYf8Q
hF4c+N8kVIsKolih3aMmh923m8TBtTjA2uqJwbPKoKaTA+gcuVvxZIzmz5KsxhovcLIMAm0+i0iJ
sILNyCa/D1xZHULoDFuDWb3mRF5yOZFpq9Xr2DujohozgngpDevkoJuXSAFFcdoT1mORUlGBfC3n
70x6GtCkacJQgS5hOLptzp4KYeD9UsxiE8/rvM+q9VIUnnn8jw1pODTv22E0HCX+lOijFoIItBcw
D5Q5TXcTctK0QRdnUHWEvwDilzsxcbpOvauD7UZMe74C5sMQSUjq5UNhu+ZFe9stimWwxMh11hAb
VJBfnerwMqcx1+1jZ5zsOTj5C430ozMbO6TrprHtr5vgsyEfHlShD8a94wTIRKf10uRTO9FFSQee
H0raf7X8BOIDT8rq5tBG60Kzx3sGwbX+eLOmj6E3c5Bc2Nv5G82gr8m21LfBNuzUJt6tZMOPzuBv
vHpmVKjBSnlJZJM7ZSiquo1fwemut2hK+lZ7y9EVDZxVnB6kJtEWKvEdezM+xFD80m0/aQfDPzrC
e+cESNTCudnEuS2zwqWDFSSDEh0n4nNHsePFIkie4jey+qT8c1T6bz1k1RXPXOT8SXV5beUHIGJ7
yFeH8ojiz0ihfSFhy6OHrTZlpVkVO5E7n6eiCmK5JVaRjvUmuPfNPY6tpTmyhJG7RNsgS/8RYsED
vaTYjEdhev/k8/tyk5+whGVM0ihWoA8zfQFgDYQnCa7mHOVpUzkpObyBX3GHnER1nyQJR8e+hTa2
dzxS01ecJNNX9r6ADMQMYCPF7AtoMckPfo9ZGdcAF9C/6/5R7rv7fWvxaKnQ29r0fupkNoH66MLT
WbNh4QvvwyHDY7vyIVZanoXhC9XaFI0/AU3I8KkPphTj+HtX2H/bGjb7OYdFwAK6ShFf5bSZwube
TknGxK2G9RSTx3w3lUIkDsY6MnVvYep4VfBxXgcO5mUq+i7/TOHETV6Crqkc1+yzOshYWRARj+zG
6wKjCzIb/q54+3+6+p8bk3D48YFWN3N05IRJckNSV+KHpRJb/Bpyum0oNkFDMGRoYwLGMnOemKfz
dkYiToO0LMMpIFvKhwNEJNUMqXcIDgJwrvtohLUNbkjpoR7sVLavhfjv4GdCIQ+yBH8UPHkgjRvC
fyoHfCQuwIYQ1yvfpw9s0unnSk5msBzJmJah18mQ4zZpu1PatlHA4dmreaW0J5TfPU+TpNs8fPxn
75Fi1vSAsyVMvZ7VGj4BvhThjWqqtWOJDxV3nVZeh+44iTBA75cGzA3GLk43Cl3LkvZIRm72aK/s
+SmzBrdpJ+DCOZt5GmuSinkHKJFJBthyABIlSDdjSceQGnDFTnD25hoJcEHaV7APkxxvvJwiXcSj
yxgPUgbgQHFyIGOcsMOvAdjoXM2bdCF4ZLZuA1S+WElJXBj2BBdZyJZLveDjSW6rDd3zTiDtEEil
JZwJbjihxcGUjkSZLR/eo7NzMCuklZtje7wMXnQ+S/WHxum1dtO1wB6sZHKgVliDtoatEZToITr5
W9FHqYKzrfdmnO0uWH3hycjkhhza8bgQZraHAtNMkcjxWvnuheIAmmFdpS4PpE8cbOGBZpXurjhl
cQbyCTQvwa3NVpFwxhz+tW+m6Ozfxx2vncd/pu5cjI1ZuH2uRcI2guAIsBqVk5bJ2ALRPNhQn332
lIMncQno1Us1eJERXcGnhV2Z+S/8O2edtT2kS8uczmPn+nmyo+j6Hu+OyLJPE+K3XaTAJGmP/+1f
1moP5rOgBDnq6A7U8l3gS9sGVVv+Rxwk+5T8eCTveyi9P37QrsLQy+M46/mC/auTA28ieaI9IcZK
PVjLOY3bEBfRrLdJvbKlPQlvPStd/7kHQ8w70G4oiUmFYDs7MWjeNYr15KPjTQE0gEU2KNQQTsSx
9RvKQMQo9MttlOLMR+JDlp4I6ghlx+3iYB+04n2MHdBxNnf4suOg8CXJ6UpE1wVIg4chgFpRBhaH
M6TPeNZ4/cH9NSCX8A8A8m62WvgNFl4To+LBEPjVM26aDpKtvt0o7pjQ1JmqZ5UH5CiyiXzfZ/+M
S3jQtVzeBKmlaPjW1dZRGsmkRsYEXXphJpLQdAurG6UuYJxVRDOG0lR/dYFnQV2nLfZeYzOVkMov
pglFlzYDwNQDamjmAuNxK77ozrxpvtygzOZAEgxurJd8zTJTJx8T1hOe7Eh0Z9l0fbunpgD6mofj
9cgTd4kuhei9BOMZhPTNyHhntTXZ2Ey8Wl9nozXJRnM3dNBo7yLgaHdJ/MENd1vaA1U833d6/LS3
jlDsDtKJ0XLK5BjpllRnZnws4hcyh4KSY8sXwQK9ENmAXG4xM0GXej4BTz4ZBuHMDDREMidsibr4
K4Wo2WKv08i2q/s1zmpJu4u+Hor3kxCR9jJ2e113rOxoCjokGKs3tdVrsOGwPrRj4X3Fae9C60/D
GpOgYBg7B2MT++YDe27N2yMj+Kvk9pMZgqy/x5Ub2sgrFssMEUuIQd9Z5edKsiGyMmcUPhlODbKE
vnrxBGacF/iex6THnq0c4kc8XUnaznkmC/QeOqoU6f99WlON3cGFxvuX9EcQeXvH++FauuezYUOs
pRCvAd/y6YY93fZnUGTcxOhrTInGEDZMLOk3Lus4foBrOaCiKl9JoZb1ccHuWKzBqhyfCSvJi0Tx
XxfeqLu+zWIjMcJdXVf0pkdKrvS9JSUUiF8l2FZMkECwu3RmQR4LAK+bB6LWJfUzGs7doWfJxjwG
H9peFBtuYJibrSuEE3RqtawKuVV/qnXN0qR6YVXa6jYGBFr5TKY3yT2y5sa2VrOBhPPYKhQNUYEo
uVXZ5DAm1OiihAqWD+2sy9qFq7pHBQNVTL0V1KwO2Tn7k7gZgsnzeoGR6aJawRM6yfJ5gYWNfDxi
yud9bi/wEcOe6pmPsmW51L5ht5wI8D6aMN3nxS4WpEQ2N7uKyE8NetIjOlojxC+fD+tcPl+LSzAj
o2/SuNZFtDBBVbnu3xhgCG9zm58nh40ByT5l6l4rZ4rkw6CxoJzCMCYTD5mvHr5/8PyUPLt9Lkiz
FufI465gxeB/XuV5eS52JE65QMIKcqPNfide3ka35oUHrJIAYssB0Z5uRnCdkv9Q3Ap9t9e1tjiN
xecHjN+V2Dg2zkesVSIF1SKb2jlrEU442nEP0ZYO3HCUzfHQ0c3cnOLWUudwk03x2FC5Kv+iEmVE
TETxhJREqYTR3pCX4gQJ9x4d1zXqMFI/ovLjCIHkMk0VQi28BFbegxVi5F0tgs3K5K2TtRL2sv5j
szmYpNLOmwRXVgzHq9ThXL3tItkWiyy/aRKiT1UWMcnkVH5GRxM/2SO2w7p+BDZGwHpvPP3+M59v
zWpUk95W0C8+8q6F5B+cbovNe7ZIt9ne77M6sDTRUK7Fj5f2LNcWo4ZOubYtJZoZgNmDTIH74ALB
LKlnY++g+kOJgXeiExiwGMEjQXETC8VZWlaYnMQVlZvgF8WIYcvK4PrDRMPplGCtPWAuRwGOKdyk
Kay/z8MNKQ+xkIiiD/SeYlZ/WhkOctoF/LFr8ur1JauIRdkVgxRZacNH0A7Ck5H/3XqCVQgg1dAY
dMl8dd0Z+ROzAJxDWtPBrSMVfMiG9KcCi2VMCWYY2vcrdwPMu1qnl7Fgy0fYwKp30CSCYZts3mWW
hbJq/JM1AVJed1kIp6606l+GYFzi2uo0rxOwmRy1jgHSmhmOkPRhNk+ovAc3uvFwG7MBKqv/cZlj
R23c+yjsP1c7Z3s9ptOZZG4UNhXkoawoF5bnUiboorqta8ITpI0YnoOhm0ncR+lmu6XtISfKcb3L
impPTIxK8vak6y1xLnbOaiBfUJTpWUEyuNs36UQXj+Rqgf+xsp9uABTKrzzfX8MPArhLIqTLTN0L
98DPX4kk8+IhO7WRmtDNMw+8W2IeYdeY64paAoVdzBytrZ5fzRg/gm5FJZbg9WeZ4n8jR19Tb84P
/eC4RNqtyzaEO+CJnL8gw2VFUFPNMEGhn8DS4093lbPUDWD/W5P5Oq2gyFSI4Kv/iBdTjt0mMwIW
XVqQaJagHep9BMc/PmJAoWN89E02mUqPYaxv/MAUrqSkV7WYKChb5NVMNCDnLwxojQsj0VAO1DXg
PIII/Pfj5aFO39Ta9floaZ5IwyvnAD9gBgmI7EPpfPaXRzn15wic2Slb5YMQMap4zSZYzCdr8wGd
DOi4TMKBYUrW6W7eY934TQFKs4PJLDVejkSF+hyb/KD+TVgnhL/h3jXC6S8GwF+RyL78+t3EZLKn
eaC7jwEcvem3aKaBWGim/MbkR9LMJEcjwI1qX4CUYRQuOpQXJVnFsGJTp5G1Fg3TeSynGt2WJ1dj
FxCuvdoK/F9LgXLprR1UVjcSQkBFBFc/LQLn3oC/l6rOsXSXqI7PXTnYXnb2Wm1JWxQ193vszmPX
wAEhzmOGsnGaubgAglFtlTZdCdZA+AHFLehtDYY5+ax711VWeZZHKBQtU8B/ehVVK132FHgTz9an
0Max7Yn+y3bJTGKVMvd8s9bhrBJX6e10pV54Ywrrm5D2hMufg5mf8zXIaatuEGc4kfmX2Mrfr+J2
IYIT1KLcZuLcraRTIbSPfbyX379Et06h4GI6246mXRkJZOSAPOreu0aRfY2QQT24jo5aJKiNapf+
RhQptAsCozRhR7jDCm1n2OeBhu/RHx5DYNTg5J7bgeyvShfrQeZ6MGACVkCgnmCeTfhmfX515kLl
kJ5x7V0xaRhK9MyVciwh015mXy+EA0sOSHFOC783TAwrM3Y/tE0zqZgIPdccqhW9WZjbZlnSs6DA
OFXR/QdlH5khpacpyNx+lj2b4q1cAfjwNWOYuUBfxchQRMyleeMQ2+Ek9RoroHOqmmwn8Vgo0vBZ
o0N17CCDDiVPQn3hBjMOzqY9cpMl30zFWfGE9O0KgRPpG96ryfYzdFYtTeatBS1LA6CcFVb/QG7W
q89Z/EyVqQgsaMmHHpD/Mev2xw3yU4KJLm0EkieuRj3NeDDJifgf0SwSWqE7ZfL5CS2yHSSVr/Hs
ri7VMXqXxKip8flYzuuW/Wq7EX3AFBjbfBrC1zCCSwBiGhEywY9MekudORlzDeLw+tgcNGNcN31y
1clGM1ALH3UNB04CrLJote+kFVJGHk7qwGzSg1UBJzEV2eGchonhHAmMD1JjcPyPJaAKXjzM6IsL
ywk/KmwtqWICq7jXSXNcbNTXTf1Hiyi3sjCA0Fdp7hOF6yRs+16pOr/X6nCS05Ihc7e02XQi2QNg
lI+EZsb4Vti3piByjYFFGOP0tIuezN/5cLf5As5owpakKHsSWDHmEF+egvQ4PKyF2N6gyIlAfNmC
pui/Q6AHXC4wtNI73b2Jnug9LuC2d+6zfPAhQXAkJ/rRfuG4d2mzsb9y1FJYWzfIG+2+9AYpyJnP
WQoVI6JBIIKMM9jWpzp7PN6KT1laEUKpYK6ETbfYLfApvedMd42nXC8Hc4En8uqQACbltCPkeQX+
MU06425iiDFm7EAmDjqemJ1dOkiMJbTLDvobTeQ26SCx8AAGs3dAhLRUuBQbn72DCzoPWShn3KZo
MC0GQPbsof28RGTfOhzTceF+cF41zVW99QqmMVtDikDE9j4hau36PDc7l/hlUAIE3O5T0qTI4G46
G2mNnppGyaYYcmYf6kywq2k9FUUNhmS9xwZm+rl3WfKn4r4fd1/bEnJauXQY/AIZQ1zS4ClLIME8
yxHxhleX5DuwTyT8RAlbjjlvGrrGlDwIfhhxbf2Ag+4bgVStUBHz8FJ0Wo4rsrNXBlAvtfcseuAn
/o6NgoC6mI3JgX+gpmr3HhA6YMNxqujf5sd5sAl3g23Zs2BLb4Uf8r66z5Hpkw+IYuGNHVg7XQq0
EW6ZK+iSGY8vvuBNSBXkHuNkNY5hEuhUvMCGOERBhcLkj+1VkO+DDo6J8/0yE/BkdiPAs6Ia/E1z
PWlMx56uG41BfGZ6GgkMTovxgSxbnY6YEx4QMfBcHLHzTpftXBQxZlOJzA8aiDAxeRO0UlhGTAfv
phtfaRHqB7qz9Bkjhgvv3/RItUsrVzrjU+nxQ5zDRiClcdNX6L/llKfwbxDrjkXihAvxifQxTw3E
Z6X3WUz6RgZ2EMJ13T3/LqWEawGkWh+zUI1oybiJwgF9vWmDiLUd60Yk9EQ3b7SHD30VNLNV1Lnn
WVn3/u1EY+aFYKeHRDNziGUgL+Md4HiAs6Q0HEoRk9xGwX5xCI+yItve7mjCzjUWhzEc0oXIqgtU
TfsacZgRpKM1V+mbbDKMBkUIVxBKy/oUm9Ne2vdayAZZnqwoAdu1iPzKdZv1WyiQGvP5edGWcdFg
Xy8L0wxznAq+kg4XgFOBtItu2g+OW8ybRI9j7569nRgj0LbFd0b4EGUywvQIV/d6HEWDjY3na+13
tviTPB53ZgIqh7louq1sEN1IonmGsRk7o4wLAiAakSLqLrz9XsvLmSr+yzbQDtntV+BElPsSt96N
8U7hkdpoXDLpKr2a+a6WeWtAvR51tllIWeEIusTt2u1vswsioHF5mdVZhG9LfqSNL3ukASl1DEKD
jX/J2xB8gtTyjLhuMuSJ6OzI15+rTDsDFXTXf7Rq2/0gm6CfpNdXJISHw4ioz6YnG3FRhq6QrsMC
D1SlIr3n8Md34XTFDv5KEwcUk9ob8v4NnhUvJJwqLJcZh/Y+4Gl1M98FoCi0dISfTsvPmHVv7reJ
wWTv1dQj1A3FTrTMIRiL9BmNegrvsjT7Z0lKoiT1iTEDcEhMEBqqhvLDqmJGDKlA9ptiHfwUC8q6
2bxZRyJqHUNvxpHvOpWGYT2d8S9raGPFEeKBtiwxwzykS2lCpraZ1uFGFv8W8Iwdh2Q94ICQ2tbY
IZhqgeKVW9MUG4pHCOZuRz3nJGxQpk+yk3HiZLIKDvJru7ILeq/KlbHZIXqTERajGmkzXwCY35eP
TvLpV66ul+9+nUj3S4vCGM0ZoTvCXB7onDAZQZ5kHJXlHDfig2ILlFuFMUgYGijCRmMymTgiEqPU
EviS30NFsvg6B8tECEI4sq2nHxJIZT3dqwQX/B+NH5n2phEi0EwjEmOTNcrXxk2yM6MyMOAEH1qz
vNNk8l+UvV7Sn+oijTbekCtQYb6EU9Qv/rll9pNYRu3sVW4lKJEMXiS3eY8tQFyxMqG7FeubKKgy
g9vXT7HFaFwJjRxkbf8WiGdMcFoUzGPS9lkzmBTK8x8YrnGpZA3R6RCqy5jKqkhvYwGQqTRN08Bx
JbeN+Xq3siJfMicauT1fm1BgsdNW2hDpWVJzpE4rXXTbUfPt0ypgLlRQsefY/K/lVfYRCUvCNB2T
x6KFDj7Gs4GRMgkJVBDwrkMArN1whFaE+Lgof5mXD/gEsxkACzNnDZw6Yu5DVXELL01FK6+QUuzN
SJQr/SfOK/7rBi2xTF5VqnVlk/D7UuIqR5coJLtOSLEGWuNIi1nnalJTH+k9VseBD4UhwgOeuA/N
tWsGYtwrHr8QfLdBgRDNW1WLTJQl01YYV7saZA6OqlxT/+PawppLIwLzoyAMf16okTZPUCBS7BuN
W/FsXczdfmvhdiJavLW7FxAv/0LD+bKPcDm97S3swla5Eeiuy6+zOzwlkXhjSUFA4+vsD8c74Qks
BJpfSA4c+35Ml/6knWhBjlaxA3NN0ZOJ7BD4sBzboslefcOQlI3IRJsFvO5YSc7iv6HeyAnL7ieU
35T9JWEUcn6aTjNbUKKUy2D/Bvv6RI49wSHT1kxBkgN0BQ4LbLe7TwdcFAnMvIfouLyls9SVC6Lr
DvZDOjmPDnnTfrbeeT7UrY0MnrjV3AwVUcgeFDiMJH3SS8hHa9lmiLCabrv+5OUb0AePLmJ1ssLo
elM0lid+am1y4SsfmpaINmVqaAlkGChh7l5EtpirIX6jQNxvSm7UR+Clt2BNF4xT0RFxLGBGQi51
V40i+nmLCdbV8230xI7Bw6ZOwWNgohXSKaylUzyrJGn2XbyB4FsqZbDsviedfBIp3d6kCSFvjnzG
/y3yVhM5QeGV3Wn0XzDk2bAagtPMolokk4IxrqwcomX/espDVSeD3P0jrpY1Xvzf2uWwWq6YNlNO
t7/w0GXAof7hC1P881fjJ724K/iN3QCdmOmtf/o36hbSgxqRYUgRaYf/kdTicsHh8jMIYin6x3xv
+4OneoRWUOefCsaCokj1t6Gu7iFKccGhwRhnPD3CaDFUPOpyzNemwEfrXD8oC5w7eI5+bVtIPMMo
3UXG8370+oqSwxrMZRRmljJ6XVytlmw8Ga0tkHbsIvXx3kNEpRmKGgufV7Y7P/igE5x4VMsPjfhN
1Ti664lLGugKEmQpYiOgc/DLe/r/tYLBlXFr9/qgCC00rnHt5U41vFYyxgPZS3jgMemQa0C6LKBI
uPxTitl4DNSEGHf7oW/nP8WFuwn8UOQUZXFbQ22fSXe0LevGcWjITHGlQBYLtzgGNMDkPivhntDF
e7QeALOVsFRGymTIgzhMx8mqW6y3gHIhMv3kHkhePgJuQ3oJMhk00QOFWMC8VSIm66JmCDTU7TF/
HpszWAeInhJvUa1+8pYH+UPonp5ctSoO3h2WlHuHVwWAy3d/sSbJruzCOnNGQpWec3zHvVBWfBTv
JESo8c4fm19yhmWF0ZYCaUMj71qUnqd3PwuTXC0kG9Bhd0A/1ypWC988rohgQ/Af2ShlRFcltrXk
XUQrH813bNRy5uASLf7Vwa6QuQc3y5AyxKQWDE0aA1hPLk8y+lzzpOKJkGLcFmTMT3Li6hlunyJj
HnL9ZpJEsAjL5JRvoIVDhvGX1o1gke24kz89E3OrMVAMS7cUtc6VN/f7VXC/DMeEjSVfG2xtwheL
WeCs01S+efz7gdU318VJw7b9NbnmChGLUe3lbAqKa5BgVKe9ETEDnG4sYCevQgAWZaKTLZex4O/M
lVPIWWRQA5EgsIV6K4du1HJEc37nD4izDpRUg1Pl8VKkkjL/vTpcMBiLBTTyAcHaH406cL3KDiRf
HIYsSjjBbKZ08j0tAijwDE04fq/DCuMzWsEl1Xb2ZgUl78jIVtXLjg3mXZ9MYcIhWxMfOw13He9B
2AN/CocDTXFk2XV2EHvYTvw16AzR/or7zjQU4Pbaa0N7f4GM/gP9yWvvP8IBFL06T1iHUGtTweHW
2QyNj4I/ymRdAjCH0IveOX3GH7D5tTNy+JEauxBPt2zq2uU2IobgQlFxOI8w+/5iImGM4knPUa4O
K/q0stKRJuERAx8Kp2TPKTBHDj5qEQv6tmMaoifZvpnbbh6B5K9+CVk9/6LkHolqjql4GXemn/s+
zDexAxvdo3CtHkwiAUd3DULLm9zdAA3hEDn3fnh6ZFJ/OqBWttzAKVFvmXd8DA5EZ1lSxJaTGQL8
1bEJmlLCM/n7xtV7uvyaR/kpv3m0cOv/df7PNag9HAU4XRJy8MYHSt1oI5OnO1R20oHjSU0v7wEx
BfPQx6wUYkdeCoNPDQkBTU7OXblWSiJfcUCtxz8Oi+h/gAvgN4pGUBAEMUhDym0jbvewyJI8xp90
ggTI1P+X8mwDodrK1P3S3FE5gMTUNhW7Bq43ayzP5rZS9K/9hpURr3TIElNzg3CKeuEBhJfY7jSt
RUCgRPpE8I2Sw+8urOqe806AMAOTibDJMkNVLsGlT3U4LxzWzLNLHMyfxc1st7CZ+EreHH6if9Gt
Z9+Gzhcur+LsilGTYgHmnsAibjkol5TXpdu+NRrzlEBnUF605vqNyBKH8fNQ7s4zvfQqQw5vOPxz
edznztNN9pONZW0Xc0/Xo1NcFhryPSzI/9aclflyO0CElQB+bO+4fqAH+MfKmBmoR4WfnfA+/pT+
yApP/URxu+5oPfi+Vo4n0/1wRrFmvwD7qswxGYkhn7SzoGZZhT8tUmqavv4KAA9KrmoBN+QVJxdV
UOxTbcYHWYvjWNNBH4yswqzer5EzXj1Q9bYV7jYkaFjLJGohmzwyDoUhBEbdcSArVX8fc0MB37QK
QMHE9PRLM9Qjo30NPtyx3Vpkl1V8SlTqQrG9wTcly50DEMeo3rLO+KIfSSCjUvLHT/RywholDH6V
knb3RZ37XHvVlblcGZ9AFZ8id6zFbQq7U9qf+bJIYX1bTk4W6ZayxDplLY0uRBQmqnReJn1258Fz
EDTOh9GFtCO6JWr01ygNjOh/aR/d306vuBb237GurG42WRIKHxoFVFZDqCG3FQToMSG4liDlvxvT
RS4gncMQlGbBKcO1Iaap/xkNFKO4t7aUmAdMd9SBwHZYYvYwwfMnISSOoYzNihievKXaWm5Ermbl
DW+GLDQqjXT+lZTb8XevaP3WTMC8r+MfvqN1rOIAKJ/xMk/97rMk4/9i1D/fSZAj1GoMHKcVvkJK
r/0lZAtAFNsQPuQEFQZqd+g98+cJ5bGo5oCjmhFSvZedMcI+PTj/a4tTcXuCujd8TjEs9YidL+zr
Y5jwNjUHId+8W1jGQGVSw2NPnCBy9RRGu+QFfG1JFGkikFy4bC+0devvDMLuZ7oiajq1iNS1fHxl
prJY0PZsBlhqCqO+YJmXEwtH0NECw1zOuLUNYYOnfxccHEdTUQ4zyQf6iS/0+Ir28ho2bplxidNO
NWoRwgpdP3eDyFy9NdCJGZ1QsS3xSpkoXD0xxyKBTfQsUhmylxf4SDA5LmICHKG/G2NP5VtT2Nby
XwBDXytTTFviwJSxC/IEu+qZZt8EJzQoLGDNTmCQupvPo4exS2PKEhkxjnRSKTuwMAFUQv60S1HL
hQaZ/4PeYFwrgvpb+Xtuk/JzsMZcg7XCuFS9VWvdbws/tSa3UMx3T5NZmLI52lcGaQcilk5CQZNA
hnA4+KE9E0VZVOZ47EdAnPgFv5wdFQmlPucsVuv5/Sq5plejdxAugw0STTDse1ln5v6OkNMOcpeD
vhFdT8ZkDyzi1fJtl15iKko7SbTclS8jaMrt9D9Fn1jAo92Rb+jbeYHLuEUxXqZrSiHdw/o9A3sI
I07riGzr6aM6e9qEdv8V+OXNisYcrJx2JEeQHqT9w8/IOb+zAVpDwAmZkKtiiSUw08KBcDkKADq7
liMEO2XgZKT/oEZCWTt2OAn6dEywN6j3vM+f8o7J+iaqFc7mf2nlbXuCwV78KgExdG3HzRdA7AUx
50brwCO+/QGnriO0XPg8g3o3Cj07cCXB3ZtMJZMFa0aBc8AlaPV1aUHHw10TdSjrXqGnMpiUJT+F
amtbXwyFOttrMicylpBqRdIBV+sces9P6NScIIEyf4RTOfu53QHvWi2FHDtIh+We3RRxbKSRnpUD
eeS9iV1LlAQ/DIDCBNWHEMiQidmyzKqZ1dTUq/To5Rmf5yQRbY8aCsFflMZEAGpuoqdQ2ixPo9oW
ou7LgPdKs/jGUZHEx4NTQR/b0HOibxm27wZUkQjLHTsy6kA5+SseTXYS8KSdTXdYyUFK/qteDi7V
Q5PokUf6M6eX5iJ5eUIzBR+pYkAYkJ8U47hjMeK2ZSuo0fpuaW4i03mkiCs4QpN9znbqTc3f+1XG
r5TMU8Y4Yed/Nbvj0osOUBdix+55lkxQHHaq02KxPQUROucNUTtXihE5XAhAoXtPnNBA+x0DUm8G
AW6HbcAqoSlg5KhJMgz9LxQNwonW/7KVegP5+m+TrGoKcQl+HdOWrQAnpD2GE9cJsLpKky9SMPET
kMUTU5dIA6AGhpcoYnOZqOGu8SrasFlwgC4MInoDvnqcwbrmgoEfKDYpWoItnOq3VOGzgfg+TxA5
Ma9xvYD60A0r584w7PM1YjbH6U2Q4aK9s15K9inhhd1HcEyjP5g2ak6YDXznSmfZW0bwjZsSEkhF
0Q8YERQYuzcK/v71ml1uSq3WPKn0LSBHqHKiifB9XAG7bjiySP5+zev4evKK6kDkeR+o3KfToKuf
EuvFeci9UrNLAsAhkRwKSLW94bpYmPRwu+FyfuE7niPrWekThC7YpTOsBg4qq60O4azZfPTa+u25
yYL8iOIK8YWdShMQDtcx06ng/PxiZUG6g1iXubLsohQGGJcjEmoOfKMqTkbhrxYJ5cahvz6YMGJ2
Eh05ZQipedpgO44RbHneZa0twBdaVF8JEmESh2mqmpeIC/JfEMu3PH4vV46DtQlkBAHAaFfsVq9m
nKeftsm8Ss5dTNja1qjY2BP4hJFExAAGzyWUbCdz64BNHIPTUvTx4zwba45H5QgyzF5XacuY3Cvw
n228sigNu9yhJUjBGOTm9NFeg+wrMPiBcbFLVyeGlYzXB1QD9yzWVbVaJIV/zUQmQjcYS12wR2O7
Su8el87KqIM7gNhXQPVv94y8aRs3YUp0feyPEtJplwX6nWm30sfkbOWyFk71DPIifY3nzL17z7GC
u2BsM2zR6+0yMTFp1Bacb58UjvzHPbCY8NCwtk8WQQzBbbjse6SdRrh6CWncRIVExAoWDDX0Oscf
skYI4WSzvu46/ssKjB87XwTpt2j1qY1VjAoiapC40n8bmoRR8ZrvyFtAzF81hqSmClRYZCP1jsBP
C4F87DJlxQAzlhCnvNWCvau+tWUbMNmxFdGcLE9hNzAMIrRiZaaHNHRuoJWU4rYk239K/YkNIgsb
8mIjQ0nmrfSl6vQneYAjNtEh1xySZiR4hJPPlDHTFYzVTnCjDDjtVyXYS+lVuucUGoQOx/tx/YKU
9bsfArbnhVr+elT28Vrh184O/qCA8mj1mKyCe1pBBGZ8Y5gO9UL6qu9ribibVeG5/3ll7zDb5t4N
HEEO7dKsQ97JLLrDx9ca9tTY5zg5pFFhwgpoDfdxVP2GxdKTDK7A9WcpAYEVL04SGr7L39JZxcuF
0JS7aVJKqj/Y6vD8kYD6drr+7jB3SG3vIJ6g+jvJaDE09JB7KNBy1s4tmC+LAQy8LFBzAX1zymAT
ee9xVDwWH76GBEZO6F6mxhDo5zG2RuQxANodL9wDIkaLEtWDlUWx3874BC4GSVL43UmaRNSq3BuU
0Y00Cs2W/Gwj09iuXsOvWy88O5D1PrB8uJLaakddl1p01DzpYYOO2lriJHNEgnRkL6otnveCqERS
op8FCOdUcScEXlVrQl4Lf0hNcE8fPLwhVrQgERNF631ZvYHOkBeTKgV8dFSgsj/lOyGg118JReKz
V/QlqN+b7Ri3i2cwqu7o3Zt5zv3fREsPQwRrK9ynj+xlwUzwiXFeGtRhP+KcCx4Vtj9rVwLJbqUi
dhitCw3e0k4iaHYr82LTSm7vZlvL/1eaBoGvzHk5GXB/4lr+dFKS8g3boGnvZmQZZXxyQkKF6BaS
sXuLldS0BjHKsKMYj96r2opdLyoe+pvWVN10GfcT6XXXwZPVVDDmQNW/1/jE/Dcsz/1kBgFFL8Sz
Ae0gKG8J/edjjs5gUrYoGrg4CfY4FsUOXSet6FHLrluS3ti6PBfQ6L0neDIcebX77HI6B8aDT4WA
R/Nw3vyk2HWzM7WnbY3gopHkFpib3P41TBMhSRxdnRzeafv3s11wFp9s/lN+z0uGiPsiD6zehGRE
f/jB1Ch/KBclICUv+XwIXpOQA1xo1Svmc14aDdJdWILjpHl+e2Arr2KBhb3RN6rzXFw36hOQWWDA
OTClA6lsVGXN4mEnCq3XUwrYN6BcAA381HTkmFEWRqEybN9TDBbthypvzUXiGGYfvi2GB9QUc7jb
0gd2nhIKL/guqaTSL6YUtQzhqyUf5hATPfLQ00dBMb8VU2N36ZZPsvV1jx6RfLs9tzZ4+suKjby0
+usi3op3by4Hs8cHX0wfQAJnMxJK9fhtNlaKsp7+mH36NC5v4ZZD4M9lVBO58OvlxDOrsrmyJRjh
xrmvedWo2FepX1IUTaUn+x3zhTtMOlacyokG+wut4Q6AJKlS0nGk4xQxWsukn1fIGV5Qm9D8FcMx
/1ks4KnwBEfwEaEFXgDf95bZS+Xz2zPKik9RG38YiIlPhOdtH5jHOwtTgoZQUwCr8I4xvHGmoaKS
0uGNc5XuAdQot9c/oZ15gVFwuJJkkENu1kYiodO6I2SbZ9qzzOK700t+cI6IQsI+sTl3Tl2EQYql
SnDgxDopScaGNKjXZIwl+dcfYL1pQ/LU+K1M8cAM+ZcObhUPfK20fCgYIvtscZlaEoAIJB7PFW/C
H7HYRpSRfCfJ3TrxpolrwtF55OEQRV8gKUJo4WAsHX5VLbnOTUbk5YbWFLGxXvNAGdPX9uYyFy5Z
W8W/ychV4kO69EEoyKnEn1k5K+1+XkRY5IiXa/DWFIjHrWQZKIR/vyYASuY4rzNe7htDh3SEZSZH
DootIWFdbyrxC92ZwCrc65S1RhxP51Sl0Nip9dejTXoh2XUHAzhgHDBoe+xbqQdOG5m5DCpph59B
NSSp6OhwXa+/8aAjbNOE7G1TwucQEeuIetUXMmq9/ZFT2Y4POU1W14VkieFKe+5YAyvuLq5BR9iB
qSqimbsjcqUOLLe13NIpJ82BFPr7tPkLoecILoTjr07mpGzeQ4e/iKntwU3hTKvSdH1MlX0dK49x
lRD8fX5GB0OyFFKX5FrOmPP4MNDg+CEbaAnFykfcP7gndq/aaWqFeMcpw7SK7dHPPox+Sz0gslaf
2wijmGC/c13bYPayPGxbs26Un/aTn0Sh0EuQgWVM7/flqlC+sFrkX5NMG/w3xG6MEZ/OEm1WNOj0
onSHgaaabmtuDcaJLNxh0eJ3OA9vNiyaxQKpkVbw2EkbfV66Hmv2nteD2foMZ+Iz5Ri0EHiJyZl6
VY7PNT5jelMKQQNxyCmPLZIYNMQbJD3cG9+Fwo9qZtHJq7Vp+8Xg8Yxvx5A12Gj1FB+YAVOBsgVo
//DV2nZLv2/5NEgqx/eJOxI9rnmUOve6fl3X9f14Ke/NsViXqMgvJ7EjLVy/cwfe1C6iL3ZmFXEN
afXBYMYMcQmim0sC53DQTGnoCTewTFLb+CTcki89ZZKkUkxjqNzPefjdQb8biAIWrYY5Dghj5rVG
t1V96iqy6drxaKc2Wa7zxZGGMCnHQ9EZhIio14FV08Qz/DZ4UR495fRBpszGlB4ARa/t9ddTsfSD
5oEawo8s7Ih71OYAPtee/mGlM1EehSg9YfJjJ14vHfw86oN02UYBRa3/pjUNmPEFylc2Kj/LDc5n
sUWRtBUDnCHbMXkIDyJXG+605wTNezNqhgV/mZP+xXUxqgv97u40TaKYFHKSSzlRzG0usJGsVWoB
6tuClGRKw1L+2Hppb17H07u9fhe2OB2So/mZu58ngkS2UvFUlnc1LeQR/mj0oYTAwn2iox0sdsmx
2NKlhVOMEbFsbHKs/QUCCsOHceY5oKiqXyL31qejpIOI+FB1CTSJ3q8BiG5dACl/qK5sJzxVoGOv
k9kIHGsT69v/5pb+Dr7MpsWOZVEC6G2QcRqdy17FlrFnmZ67nXqVPsL1YPojLitYWAuPFXOp/glh
H0gtn8NZT8zqHv/NFRp8/rjYdw/RX9S3PkIq+j5W9cCidbbUtgEt0PmfPAs4UUinAulNQIQkoxQ6
MhehQ+1CPU5tbSvzNtTmx9onhc3LwwEjPoL6n7h4ykiBy4/CafFen9Z2PEdEUVKlBiX2+i8SZpb/
gb0oJdba7Uk92r1nG3kstQk9abmBGrilT6uaRk53riKw7jn/RdCOSdJJ/2ANturQfm8GKa6Vnq0x
7zAnINctKz+jRJ0PZK+cHPljiqVrKLLXgMV4mMCUVQ660b+YGsWVAFurT93elhyJfi8Je5Jz65Hh
Tx787SM2ALnal/ekqFFbx/ATxzp9CPQPIhnsc2lhildGzTNbvUE6MIV1GIoYBp3ErwJGag4i3FJm
+VukzPLnmIsfJ20OYEF7Nlh0dZpiEUs6fZ84LB4MajU/oxXxFJuhMdLYMf495cPKSnZQJSC7nvwn
HF0yqM86Pg2adfl2q45g+3DQ1TtNDXCBM6zFgPtGb9QQMjsS2/dnlQLbNmLkXpqEvaXu3SBh2vlz
HOwvnFKEEk2sCIMcinjCsI8rJz8WROBxXvau1ohEaMsVXKvwm5bdHgqAhRu2e4c93GjRLXGDPRJd
ozeA9uodsR6NrG2I8fhAAhtKMBJay7w1EZVvyxuj7cIKgT48kZdF5ADeYQZQhyhXRE+ZIAKM0o1+
NRnRrxnSDT1YmsspugqYxmtqHICKCpgGiMQnICYlBp3D7O6hJ8QoGyppSmo2P6xA7HYhedoL/vV7
sve6fBCUvtp0jmP+0M7qy2HoUqJM6Oer6xXUfz/UuaHHV5FO8YVipX1mAUW8+gB2SkRfvIH3K7sU
qViyLx+Mw+rKcMAIcQyqg6jYEeVSGVPzHhWajCWaIplUjmkJlhv2EujHg9bgV4Zd0s7VeElNPdXM
+Zch7GQxrKKI6U8/oqUjjIuDjBrNSWjKzpzwPlpNf505T/3cMZj9QsqcXHrWvbbL5sfervsLMNo0
KxroLOMf9h899UaGB/h7vRT7Gq5qGlS9tAwvlSlTHG08n775Rkb39P8mz17Tu3ubS5Zj+peA1Oxc
MbQHhRo2DOYog3mHvqUAf6g42CHhXrjhOJgAlOyyFSPzTa9yEnADHECxA56sbZCYzxAc5QP0F7hH
k6l3Y59I1dr9SktYujutu+TvSGt1/WbJWF3mbb4BPJALxb6teHTaCGW3iluMQDXR3e+vMAhse5ij
IzNiOIA2wmZMdeq9/XV+3nxmkMTwiSkPY0JJGfYdD8iT56K7WKHMbZ64Lls65OZr4RPISc56JHqe
n5dQJIHPFo1sy+BoFSYJC03/d8JaBFw7TGB+3SWnRLEc0REXn6FF2Ad4hFPY9UJCc1J5Qm6RB6Og
lDK0eLwxpFsMjkxUOfSMVVQIx3GnxCDTnM9n2gBvDM6njpwvrYCovzAbKAOHO2vfrFGkrG+1T0P5
L6S8FAeBwkzI6YCkLjrfjJocslqpNWNc7AciGD2AOQyIVRCNJnHZPlHPdvh8zupaSxIcbWRvbkDG
BGU3cQt29AXeKRBSTr6IEXH/h7FPyPk8dzSs43v5I46ELl73PRdHzC7CorrFY47HJ5LWBVV7tktI
+I40k9Rk1MFY9RJoBMOhcANb69Ys9PgfaK/BvkjZaZUM1I+L4IVXV/iWEanTWXV8QDZwSEJZEmuF
38vMWgC8ouJW5fyh87tblHmXw0Xsl1k+lHQrJM2+BKhotp9hdHdaypkzTISGRkW+Mn9VZ8euCSk3
voWXxIohtZfwm/+9cMtn+Gmx3NX6oJbCggVpknu9NSyGNIIkNvjthpZ0XX4pc6gtpeZlVS8VIy2w
eKenbP+v23ZeSsGmuCAsQBSyZoW0peUy0MG5g7aS5K4IaL8BmybEQPBoFiiOtovW7c7OVxjnSxxQ
Zs94lWdxXJRcyqZJ8bWiUQcn6ZemODoPJQ7a3MvrQq/cujB0lY4r+YNaY145fceEVRl8LDjPVYSV
MnYfP99ynvZeXG0wLtmvBy1TVdTZaqRSUV+NDHP2fKDdAl7OmLBGIT82S0sEpjefENWoSEx+hBJ0
gwHpfUz/jdwRYQJ5NteGR+MqzkEv0v1LfKBzQ/dmPl2q/iuoEMeARKDw2L5ucUKby8hoSsMh1HHO
44HJixoIjpoMjzrnpWD8EQnbqgpp+3tR4hlKzqVbSPql56wG10zr+g7j0RX468KxPGLtInr+tnMd
qX4gQ68lStoUVIMMC2pONlZ9+uM4tHpwZli17nz6iLbBCSA2iurjYwF1O9b54kVCFfj/q39kpJJU
XS5S1LbflyJquruuj7pnVooPBgPt4Wxu0LaeKw+cbrshTRQJNZNleGXgzGQwO7D+JNAJ7yCQyey3
+AobZ7A9nmmSTlIgeR1Ne4LsBZZLkWW1IU8HXrH+TxQ5hHD4NxafTGFmcqy043MxzVWCGH51LKRQ
JvLSfFZqiUFWapKmZQhGtTRFZwn/b8gB4ecSC9Kta8QFrAvO0qvFcglWqX7X4SaaiGT1TvTPPq1s
dwCKIW6Zux8up/gUzXMWAoCWThwD5wtbGoRM45O4sulnhl3Kgwvjk5aeAlrvvDeBQF5Hgug2kc7+
7C+KHpVnXmozTMQJLDcQO7UqLL2y7W+zv8o9aK2CEU9+XkRYPccg8wH0A66FyxRRMXkSscI15U/J
bjjFQm4n3wY+kvFn6nJz96rNfTCtTaBi8DAwqo6VILE6j4RWGR0MvD6szHYrAi9dTkbrFC5jjON6
Xb9scyizS2Yxusw1vxzKsHgzhi2S4Ank3UEYq2I3n8TxJHQUHafiFe0T5lhr1BKCl7jKFw/4Po9f
CQnr57KfFQBio1+DMXlty2Xm01xM4qiGP3ygzalOfwduKILxm8s3+X++JHSv4kssgMr0zVtZNcJW
KVMSJ/j/chK03QHA803BXGh8TKvc6zgOfZXDaTMIZvYMV4l3uMAi1URmFSaBUUsOn5fqmIsuvZcS
JCkCLarOJE0n7O5egVL68Vq4Tlf/Mj6T/mDOoFMoCZwfudUeNTshHda43fv/bb319F05LqBKfflD
F7nQ4/MeVy40j5PMgBZDlC1/Dske/W9u6OZR0H1zgzU/Ev07QPpuX0rVgMRmILHKCNcsgj+Hkm2O
yQTsojGUc14RdhpL533fv+cfSv5os5G+Q1ZccQ6y12oe+2F4v3wSnpTZ6r4x1a7ZDevEnZ9zQAtf
jJgS9ivNr5YdXVRBdFjpRhhPEqbORvsiEu52kZgUDA3K33MQx2nZypuP7B0aO3Yf/2Px0Ix9Pp+u
Wj9n5TWL29RxXPZMvluSzDO87EtMgplBVZAkSrc/bSFZSFVm0zS/B+noXaTJAbiqAzjUUKaVfZVI
Q8Xj5cq9P1rLi9zrHygq2qDdYiW2HXy7AzHeXovY/5Cg6+L8hEOuH7CyJVcvfMmzRJjDgEO/sbbH
SLyYfkpQ18tB4qhcoMiY+rCb0USIOseHX4yVmnZV/t5RMbHxr9MSr1ZrMfSwzmFq9Q1DA7+zDkUQ
o1OqSBSEVBZVKqtwdMAP/TqcaWtgY7OHD14QsYvLiH7MKj90XyhkPCSoCfC7DfN6BYKegbQEmq3Y
V6JAj9IvD87HocobTYyMt5dkCqpT3h43perbmnD5b4THO+Ma4hF/0OOvyWhMPzIvVHEv+J4FI5se
PfaSzHt6EyZuqQajDX+uwEvl5mx3JjAUmwLmIglWZX8KOOrpG9NODDQY0WDcDAUPujqH+OvHDPsC
Nj5oRUc7moGebSvKMduaf0+LscYDUO1xGl6PcmDL5GsBrn+CmgF4HBpVa4bwcz+J0xFwEiJgA/15
A1VUttRNuPYLJDxMRzdmjiEa8udADu/Lq0xHKnxzhsSGkom3P/b5StLA+BtJY5gJN0F5FALYGeHB
TXoxpQbt/kbd6tbTiQiNYLKJ9Awzv6pil2sLDAriAvpVOw3oxdThDFf77VKZ6ugo1GxaD4dFRZzm
nWy36n3PwAzj5UDiplFSizlnFo1LERYmArSqdjnygwu47gQvG65QfAPvUco8jlw5EjFwo+Y7FgdX
NMJFgci7Ifo8kDRRhVDkBiMy+MyhGMPqoRVnJptlDmGuyuMjGDgN54wW2VJ9kLRwC/YWYufjY1tO
5ef8z4ahypsXjjxuYKTthV+Liau4i422mmgfUfWydc2sOeflnUgFaAE/pLdrg5jBvvNaC6/pCYeY
YXDSaiLxlPuHT5iyl97mtP3uZZVxfUMPfBXmcbBt5Mf+Hr6UIUWSRSGs7SRXcS+CiJs3lefHWNwv
qYQOWhnmqLyJmT5/rvsRQC7UUyjWcBEXdfafNjibqs/QVK674dwiosK/5ujuLbxdROBT/Lf46eD3
SshSRBjBW0La+kU5bvgqrXO0Tab95gB/x/hfW45hL9w1KVlTrnRFgom/oMMoERiEeakkGUgDCm9k
nRm3FjeUH7BUDpGBt2DUpynXMKZvAwIjA5e0czIBOLaGARSozS4ktvgWvTW1Xz9pp+1c8hRWBMih
VD3rhNJbe5ut/XX3j5gwZ9TvRRcIYaAI5d6I4t2HqRrI7qxWbbPMg+M6JOszq36bMWtTKvHs77Y5
GOzofqEuB48LHEbzvajPzk6uPGVtNvK2BxTF+GAiTC7S13lNeKEJ3js/k78vB1DrVYgpPgzOoD72
tyDpJ9uH67FA5SJ8aRYxRR/JQ7pt0rrEKmY0aevOU7zSOGwj54J+cYIMEDEhFKdlzlNQj+wbpqC9
WaEMyMBbPO7c0f4rzCY/a/SojIIWpuPVjwwxIn52SVLgBrdmX1F7PUHFtkXUngIQONnFdaXU7hNC
SP6RrCZVTZa5LYTknBmvZ6z19EyzHvLA476i+5yW04RBZRm6vlC5qb3vdgzluVsLrfAJkWTn6/Ml
GkhAol4BtdjPCrzXm1ywS9JSDMeujK5QtpuxWJiKy3ka9ZY6zSlsDCRhpy37cnwKcxp+tj2hxQNi
5za8HoG5JVZPvAI16BJY7vOrjlTQyT7kw+Cq8WrKcCgUi+Bf0plTeF0Hm0s6AkSD4A/p/8gpnztD
A2PC8o65aGhug03b0IRay/sueBdO0D+MMj3BeDRubPWhEgN0YpAtzZjQ0RCha2DwLPFwYgYZMnU9
QVaiiQGKM/WkDDXYhtdgzxKEqEYI55vOODKT11Erszow/lhWJAzLR988gs3wOrmny5nHuozqHm+3
Y+97d0wSZB2RHr8Ek8sxfcOVOyWU5V3wcYi9/YWA7GOQAUwwqL73LKTQyg6rXf+FhUx9gNlz+LkX
vIkXEHEZn99LHZfgoSNri6Y90Vu3LAD7qHUGmQBUaKfd9Oc7+zw+nOgiAwtzsIGaj5S90cgpvuGQ
nl3YhIOGkD6ZFk1QCuv94Z4cBLGrXi0/hEpq//B7XNNpUXnNYML8wfL7+rDgs3oxf6jeLCTaFaig
P1czXgNakFxJlnRETfKoQGQHli9j5QmbmSsY2Ql/oK5Wfe11X0NHLA5ct/sd1mMR6paY+axNGpS+
C3bnS4pbZbTgvecOyCo9SvmFZ7wSRKCFV4/5KVeinBKiKSiFqc+tbGV9Gd9sadbyxiG5D4SQmzO/
DWrJKOEdH/q37hUm+suHwbRJjXnyScRcc/xOWwCpWdaW48vUIpYMnntx/urL4o7rC/2Q/HrM6B6A
MOkh+EHErsbRengH507HmJdITC0kxMbKHwRTl4Sybk1Co5tjFGuaKDx9NeyUbaPVkezMX4CG7GxQ
LCiqgd1+r//m40JWnS1NTnRfgE4Lw0TiMZJrlke3/dn11TclEbDO2BPPaMB6qfTTDJzMV+yHKqZy
iapmzr9a+VvC1MFY1GUHG0ZIRLnklzyoeLqJ0eFsMVetwf2wvnp85d4RPGYvgxQbYNHdRJA6eb/F
EFpBB0jaCOrmrcAZnc2XGBmumJS5V5dumqT5UuqdxNh6hvmAoFc39LbiuJAu50Ulhr7Gl2MkMlr/
Ta42Uy1NmU8amhTUmVjYYSU7TbnD7TOZ2i4uRbVhqqKBVIuwVYdVz0LHKTMRIwncrvs3Er8SdZTQ
O/UHYdE33djboYa9z4xQQucQUNLCEhMXanEnryYDNfubB8ouBcqEnlNM7ltPJfgTT5mflBysHe5l
WtzuzdBn8QuIxUkQg4uspIcbVqi6ZnCdfq+iYVAXquvkJCW6P1iMhoFJV3ShKz8+MK1qP8kf6z/S
AMDvmK+gqelyXfxUBeqhLqzzuQwAHNPPwtkiAqZNWnFsoodPSZgzmtXUNakJyr0Pxgdl1WjToRQ3
3Pv6rCXz1L7ExQB1jXJfdTJfEXTddVlESrOFxk2Sf8VUvsGOIXC+MVmpAMyF4PL3fT3u2FZ2LAuQ
dCgs/UdbkNIoS7uyWd5/fcXTWZrigMnX3gufnRTI+G8LJaOABHpbkhYr0qbfEPpqjRes7T2BffhR
LHk4b3rUVZ/Gij0B4zdeHdhsaH59NBEhAhvcBqlXKKQvqUiHFvpKofmpKvDQemKbkfos27p9kWgo
JuyunuAzX9KPsUXkb/k+MOOIzIGLW4unCJmA0E5qnknI1y6QVR8OR8Sms9h4mipI+H9hnuVR+aFu
WaW620k3q6zoEtcqVJTlhEVfZ3GBs5DyKlkr38g/qoXEl4Z4G7lKY7xLkGD5EPA/veOOhlsAEQuh
fmAA1n2kJLQ1Sq7OzTdFgJY9e1UGbUb6z+vIsACoOyATxgrPz0GEC63kPxvCVhVLriOQe/ubLlgN
A8MBICFfRi476Pecr57Z9bLmv6A9jd7+TMiQozKvzqp0h/OR0zrtA05hoqkYJCuqRUiQtSmK4fjh
3s4Nh4YTQ+Dc1BeVuZaEbD6qRUv+rTQ2LiujOGRE78fyhByubEdjzVx/rCaJysjl8foJrNVlakgh
iSXSgIeI9/AwXxuGyPShJqUaLpYLoR1NOVlKc0nCVNvgMPYZF/ex/oZELhZnaJVyUqlKAxsGT2z3
ja4M+7TEDqlVi0aq7rMOKf07+giW9zVHT5DjptOjU2TyxNCIZ5/Ws7BSwfM+Oj7le8tw/Xs1ohwf
eyTGze/GVnaCP+ODGi/QLLgEluM3u/BGREenkSNv9ATDP9kMB9HPT1zM63QK21GBdxRThp2TBHJ4
J00eBfTlGbwSv8WiNP8HmRzIGgRzEFijDwoX62IY5kmaueNUBCpa9gvlV8MSzywUh4Ra9DYQhTcd
M55vyJY9EpJonrgiT5cJB0M8792rijrlP57ik/+v56wPCtGFJB5UHkml22YE+IpSex+yxOCq0Uoz
NjjeBIATuSJuRbJ0PQsaEIAdhePGhHEUswNwsbpiEnM9baHjalxGw2rMcLe0B316j5baHFrUtus3
I1SVV7U9fzbqy/12C11gD+s8JzDaGdRXnG9Qhp4ootEJJgZLnS//zmiEX69DWFIBj7fGfQaxuJeM
e+UcSzPIOnvuv6faxHB6tJ6mKWOVPXS/rwV+ztlgrQfXpNTltDc/mPelM9e9GdSfkE8s5pf0Deoo
A3VnY1yEwIRmGepv2yO/pNGO4ownJZre04FjwLnNH0+Jk+KhgZVqftFBcuSBp+QrAqR6mvZKydF2
VVCScPsNsRhgyff+xw9SGjggVUkgN7YXtdt6RGXSbeC7zVHEajhRP4ASsCP9kcIUyC16vieSOqYc
n33Iv6MLI8uesfy79jxxbA08cKJsVtcrq+Hulh2i/Gkm7eBv/7xZnxRlN7Ufr2ATOnxfWG/IUFWb
MgF0K450rnef+b+5/vt5XvHVCD2uQWTafpfApEQkFLpaDK90iAr2EP3vcobT0Dk4qCyX9lGiDnmg
64LukdbkoRlGkbTh7UWIOa54D0GsVfQOCCi8/X5JCBv3uQVEXJgSPflj/V1/+A+YhW9eR3/ZMRBo
DUjPg4AiHKd1L45B9qq7bdNFtVAo41NFHF5AwC2k494ikch9FyfeUTZuHTOaHhr1a9/rQBVWX2HD
n3MQrZSMBpN9rFTeHAe0aM8oN5hReZ7JMwLfOcWGVqpHOAYYQDUwjiGVcTuoT5Y8ynxl3irk0L0l
CWOXOzWtwBH7G0HN1RK33oQWlXd6KVn0gx4WQEXbjnDNr5AJGoRXHRS5YNOdipqVmVF2UMIDxlDW
sf+mpVeMY81qJHH8BuZ5y50so2sL32e5x85M3jtS/VnEC/bETCCtt38OTbvgBCdDOhv+GtquT5is
FVGhxg15xIq7fjM8xbUVO0D630LueGUv8cVH5HDEbWZq2qXzt7qNb+4nmywirYOkEPuJUAGAiSWS
hxrzcnlkJFsOyxiXQhZck5fxtssoMgE/OrDaC14WQDGijUv7uyJlT+IAUFGPCCNJqX+NaG/x7Bci
VLuuKFxWntzgFVvDLT88cifBcHJUM5JM2p6UYpjztKdSlnlzO7lq2f7xuWrgngnkYAgW+gx/Mpwd
IkNS6QTh37lshWTr3i8ANZhW1lzrIyqJGlhcaT9gM0urq5VdT1DCbhZTqGwUwdQM3aX7yGa9p/6N
b9quUuK4Kd498KWJP+YHci9uFTc6ghgxMFX1TKEGNlvw/RCRoZ5E0SOSNTVSBhb9ljOUtTBHW7JD
9/8FxqWR5A5Yy78cgLbMFArkV/yWpzEeKK355YpZDTNMJPmXD+GNHwAV3qGQMcB2spt5d4oNTAAu
MmqHlIp0k9Yt2g+gEPavmw1IrtjPGzYOKX8sv9z6m4Ex8tpiHaNqDIY4nBWShGk26cfVaFcCEyqN
1XYz1+IJIZSg+dAwf8fXMe1dR+D22mM8UC1jAw+ubCMDk8HlBcVZsb+LO+cawZgSU8u7TCS/1zgc
2B1GoEhVL1qJhr4ROwGzf7pkyITvhAirnW7nEtxuG9Y8w84CXGHrrkzMvuOIt+2sjyr0qCG7J+JP
sYQIOS6ST3MV2ILZMecMmBfoQsOQhrQmMx8fhTf0kOL90RxSEdLF6iRW70zO+aNmcnFig2tXM7C1
zznGfHXQIW179SWEu+YpB6M1iBJQlizs9sItV3h7EPlRiIFmR/XEDzelWzEUA8CI4ECeWhb+NjGK
W9v7NKzz7q2ygApkJASr6VKKVKfz0VHBHCiQHKPewRO0nq1i9ibBhPbfSeeFew/MlDsgw6EGS4O1
v8SmNGQx+EW57/rIEuQGztfClgW/8zNyJYx7THPe2dIXtVwiuOC5A2tA0t/3McH5TlYoXvI4D8IQ
qZfaXSqpXTY8jIMEzIvZgfRs0CdDPdS2nJBczePNZnAW1gkb+xqyKG136fHcNDDmaTuFCOk7iGjP
l1k9mMdMj9PCjsCHSzU7Qg8FekU+ekSrm3fQ1CN6eK1N3ztoRsBkQ9XjM+0H9oU7Nt4g9zVTmorh
HcBrJfa1yJ2weAF3Kz9NfOvFbWLHon7J79jYJYkgdEtUd6KZ6CUi5M8H02nz6jXBFiKPH0ki7yRV
Tq53Oi6j1X6lliSgNAbUWYXLDAsJBkMkXZdcKu78gRnIJXbf52xsizYORPOJV9DyHprazyp89wzG
WARJBbDyX/f5W6KalnpSH4cn+URoMzASICtEA62ElD719tMQ5Oz/L1SjL1EtW2yzq+fYgudyGlnN
374tnQb3EPVfE4CN8RWZdfbUlPiGNmyUqI6n/ioq5ydHrPhmaDxjxU819qlAjkzW095aMmunAbmj
DIE8gIIz4d2b6pRdC63lyWhdNAtLXc1cAndg2zIWpbY9DROiVEcIhOmRlQMdgf84RwabJguZ8XR2
HGcVxamzgxD7KlQjNxE6iaeNjZo5yXUR2dQaBkEXKCr1WmZOcp/T0cAJPx4zIraZV8kNZ3RN49gW
r42S2WLTpESsjlSy/85I0/ho1XM1VJOG9I6ubx5Y8oVzZjL8AyyMUARpW5Lowmfzwvhabd/YhegR
nsOoF1MvHF10u7xQDdEM8gwknS0EqjJz5yf0el8W2W8FzCzNt0OgruFfRYM9R4W1qWgFsZ1mUOkI
DzlhRe/wiqfxaVCe+DzFk/6gbWByjvIsGb+poPDGEwOj2DbT+B+7q8okjDyVs2Zf3PTTnWES6oQC
fUvEs1NVydF5tWqD/610J7e/lUNwJI/Dgl7GVAsTatdi7ZsEw++VFd1WZI3eKodqeLVx2zMvGLDi
ZAlwdXiLLM5aRbyK/sbcJFSJEruL+JcAz8/6Ug2HbliabV31Oq5Xvyu9zG/+wZrJMrdRT2LeQ/+r
Oc+WgCwl0E1JFPP317vknMtqw8t1gnJQOIACHccGvgHHy8AoIianXkHTw3BWOt7yMrJbKDmvayL0
zB9BxgI4fjITUtDRZ7WFoni6VAB9xkb7XJ0D2vp0f9ByvEnS4EOiQ894Q6Lj4HNjr65C4BgkdGw0
JHi6KNgrRkU2nQLUEkwHzLCsZ7tFVJMece1ZQ4Qkp0uOj9fju5ITgXCtSMYk0L8Vv40V5GSlBKlY
d1BTsmz2DiMiQavHQD0dBS5dJEKK5M/WikcVjY58sjdiPKFcU82uRpzMtmbncV+NCbaQvO/yw+DB
y5RJcbuU8bHX4WSfi/OOzbsxBknNKLUbscIlzNH7PJtMtTIGxYaIw0VINpdu5lVVGx3xuvIbMw1Q
DG0fUjMIMvo5SaJSfoo+v2sPaU6jxAA0YMTVpM8D8E4u1EySt13UnFe1EJQ0r9fDX3LxdvVwJ9AE
vaj6/1naq8OOeeTbp/ZCcJfPPPGuFWLH2BYLc9Q/z7zOD78RLgid3YlXb4BevC3KTPg5ayIcINRY
vjAlUDubNB5wCfHDCPWtsIVpzDUJ+Fh4ojMpjWc9puQT7IPGua13iAoQtUnx1H5Bm9nf7QTNM0jK
0MtfMFXO8sSrV+1xcmFml7leVyWJPo51xGv0o1vKt5Ua8BNSd9gpStbP9sOG+UDrqCrTeB+tUtus
Au+w1KEevaJILAau6qArRmvDm3aj95/QZ/t6Kg01iwlQRmiV/nrxg5qQ1vBqaBfsxQJmY+5SKuYF
usbWwH59IESnEhV672s6n6RexND8Q7JskS6PPtNhDxkAGM5i6NjEyQnjCTQpx47j4pxBViTCAZ2T
jVr7/Vx+anX99QKbPDgxCKPYGHpVM0y029HWlLw9pCfIr25qA2MyxV6xzZZmsn4P8IAGbuNe1/xY
lQ8DKEpb9LU6tsn8FOnvek1DlkWJSKLsZw1jc5tQ2ulo+IxOr5VPn25Y5oa/JE5F6HLfMaYKTQB2
8GhPQ0KnBdybNKMUi5/1rGr6Ll/NRYQv7+txeWjWIOfAka9BahzmewMM515SVbopjmpJLpQGCB1L
XIlITQrf+kXlNjzn+clbnHi3wvGimrxBDTVEKZbc5X4NHlEtVGm70Kd/NdpwE2BD+oUmROcNmINs
ktdCSC0XSliWMPiYGwjQGi4C0JLwU7Ff8vWvkc0UCtR4rIQDr+3rgtQ/TYSdfh1MailREaGq0Vjd
V7taVEZvnLlKrvvPg+mO+/gcsaJJ+NON9BZnH6IAQogPwgOA7KfxxfmnOHq8aj30T0Ti0siyX4NO
+R4jU0DRTFc5E+9bRDD8BeSnsPM7IEUrSdoHEsmQM6hP2USDnBsjYVc6qbjnOiJzFhzhjKXd/F1/
bG9XdcGm9Qp2FiS/Gg2gFQ5rO9/bqU38aDv/mfJaFMDREk8SUlfize2dnPScmfznSDSpD7KhLLIE
qI/xb7FuEHyv3MrYAVi26TMOmO3Ej41Kqf3nr+BljcxMo6cgFnPv5KVBzgniS1hMp8mea0hh/WtV
9u78Qn1KeTKywcMLSGChU3RAW/vZipbfD8zMOlAyuNDko445ki3UTiJ3kiVoo9ja9fk15oFuhGvo
3ppCaFltQMfOvlTfI8ZR/KY5TpzNqJgyoOcjYb3sDuIESCDKfR0eJHhHpoOgxLWddgV12EDMpEck
oFS/FLKidapjwTa1Orj8VCtH8rVe8Yxajyf2eiY8rs4+tkzDbPidsHBDgD7mtYKSHjhkBpgeYa/4
Ropin7KE+JjwYMC41oSsngytoG1mI+DcoeisZxi9a8rwoRqhedHcQDPnxLaX5JhArMRaDYDCGuTc
Mfk8bigRV0xe/cQvRphtlB2+38T2IGUj7E/NNS1gFrlELqLkg/SuVMFZ1EdjqWzP6pbhtMvh29GM
kq21WPv8DS1KVZ9eI8RCj/hK+M6PwQcj6KbTsZ7kYpYKiF5+ae67K1oAf1azQtDGp62Sl+JYwAcf
fqay+ouvVi6IBvjeT5QFF9yXM8WCg6uvLCvNw0xaTbI42gK4HgjyB70uUIN2mDQBRI/TGDNYuE+7
edxMLmgUW1yn8qV35lvEZmK7sOOgKxFs8sWDLkzI+8goNh9yqRjK9x7bPEE2epJGRkJF3bLw34fk
SQZxKpvNosPXpa27EVGUvE3OXLUO2S45N6Ko7gvU/WqDoSqUctlzcJhfGE/PhcHxbLifYkj0cOZY
3x5+fqerZIT4ezt/CZOo2uMHkmDQhcevoQIEkKTIL4MBNYqmHrtUSPzg2lNblSKYv2OWjYEC/LRo
1IFFscAQg/HrUPVhJ+oMhDFKqqYcJlj0jqqvjKEYTG3Bp8KrgIB2tTjE9F+BHaczLWSIfMrxMkwW
Nu9xvLa1NQAPWZmBHqxFI5HOlsMru1ahiQJl4zsobC9RVoDQ0kb+TnLxBZWMkhArVztS5U6Ddx4r
j6xMG9ToTuyyBs/WBxQkchbVWE4Y7aTc0veoEny3FWdYkpuH/VeZlsopjdXtl3/5j/ue0dx9qVjh
5geMHNZN801puU4B7N+G1ai2koDoc6WVJQCGh2E2Ifffg8KsxNJ7pby+3EIJ3tRDnqkFE1pDt8/R
tPh0LdNIM4bFodkrkSTiSpD2qfcEFGfl6j79hO4huWXALSYE9R+P0pz3gnSG48gBI+Q8jhPnQwp4
W165086zg6vz9KYzKXcknJLEV4KxBGvI0jUsJdZW4q98GwIMkHSKYImWRwmzfPDYut2mLuSFgehw
KWZU8hAUcmO96V07Z9BHLCTsMW/8zY0OFaU92VRROBrJ7xz5glebttnHolGoyuHmq8qgTynFf46N
kJ7jb3cVULdjHAA7LDUA3WYVziZAf/wmYu1nIRROpIbUN3HYiNmuYnUqdUtvAE9HwinB6s3DHlYe
7/79SdOCOTfVXMOr8HF+qcBz7+JNbcjV4jy71b5Tl42d1KNXQY0zSxm8AFZIk12uRDQbHHQkbiPO
cT2YEb9OIriusdFhE/+peBCVJ/hAaTv5iW/em/axZzC8BEqHVgFL+zK19X8uFOPpXkME0EPxkaUN
7VGgVW+WXUOW7zKnlUzkmKW4Hiva5Nb3KwdMNLntWnwLQMUiGrvkwj0pQkSnhOvRh4nySmSLco/6
n46AiW6UZFDPvB911LGLacPw3LMCiXM9JbhXcpnXrCgXM/u1ayWK5vTWXlNgWkcqAV33cEAp32Ul
3jm5x+Vn8a8YrQAJpE3lBJ1+3pbGnXdL/CHj53kWeSdu2Al34F6WIAQ/MdaH3YTHAaQh+dPTxAhm
EJgblI8jSV9DMQ5V2rh7Ma9h1dnsBLCrGJE6L+5clK2h9CCy/Qc/UVt/WYBljaBNVQ/zMmvsrSR/
9Xbq1xECM/d/Gk+INQn/0n+ogWS4zqD4tUkaRaMrPxn2Yzv7+2WlTC0ZYcWLjoLrPOPuDzhdHA7L
KQKxZkh+hWQJOjJKXYeruhn+xuxNJNA9YnzyWuQipSWZ/RdFu5PdhRxn70g+Bhd5ZGVCwm/V3sMg
Ne4nqYxylGwouh2wg2u018KAVi1u+yqzlc3irbXetOzfWil01CHkeTsuA8/pCEcWfF6VKWPEKDJg
TVxE4CawoyP3RcCMUDNEAePpp4lAFmBgEdNKIUqaV1nQiJC1n7HXxWhKhDy40Uq2fzpdCdXUk4PB
YqZqoMmtHhvREivGidsq5mJDcXYXQKU8pqUR2GsfDEAH76Ghq7t9KaeZ7fl333RpkQejeg8wxLew
VDJM5J9hSM3hlQpxhZkALwho95/nGd+KL79Wajb5eIXQNDNsqDV+szZvDFiS7bKj6d3xOUZc4LbW
pKmo0hQ/I/A32renipZRWBfsH8ELDW2OZT1zWcGeSsWKzV1/DHb86sKLGYztbR6iLUkP7u1nktZ1
xTNidO5Gg72ECKTAIJ7n3IVZ+PSbtHI3AmbryKf/4Nt/YiTLqcXLHX3ZsuGHfYaogqY2pelANGnO
4SfFq8Id8SAQI+yj1gOKuZGF0jF89F05JaYnM0b0G6jHVss1cPAP8L5fPKM2+qnm+ZxueJ4gWIzC
u131OhBih4yy8IRaYfqe22q8qQRxRSBpCWTYHxc7IDoWisJQJSpAXH2SlIUfakIMS3Psl4HAMY5E
ex7ZfdqCDRsZCSx5m5EhqX/4pG+Rkjn3rcE+Y/PCFy+jtuCs7+zquYQvS/5lA46JoXbCwA263eu2
uYdTy1505Ok8sCnHpcmxFv77uU1HJwvwf7vZPL+LAOWlX9pCwqWkvOqNTqQODbVP4u/B/cQKvwCx
RGZJtjF83O2NjYNqGxShBrzR57CpDKnHH+K9QDQKVoQ6yqWHMlcYCrvoFOzTbIqm014z2+bL14wg
6W59BanejaXljnjn2AqzxqRcJSlJXLg/z5B3aQHBJCb7X77e7R9XlD+t5o5M0Zt4qVaz4HMvUaRq
HmEHW7P10qyHnaoeb3Pb46ufI3jSZOdT7HXKKtPKtgDg8P4wfi7dkRqDtEfyxVoi39xu2sg/XoAb
k1wc6a31S88YkZ+RuTe7zRz/7Eft065vjJb6OnP4zfjobc4nNm8KsxCp79L6FY/fBT368fSDMENg
iEej4OZuaZFFqqAFMltx60OLebO1AAui92w0IrfW3vXM66EqaHRbbhSvv3txW6qbDoWjtGX8Z3Yd
AwnYjR4g/GrstsL1GuJohLUHKfYwrWaEPqOhMYcf1G775Zw+hX44Edzfrm5SMyRRi6fbRQTl9Ltz
sV+UoceFatO+V2gudN07klMgpIAvVaCx9ztDseCvbHNvOTyZMLSXnXEbl8ab6b6JOLxke/yQwLtU
np6jA1QYkhnrpJa6Zytzvee3FU1u0kkllXI09Ra2lOPhDjTfWyoDi+Y2gPwGpYY/XieTZWAo53TO
ayRRqHRCrwm2iyy14IjdYU4tyWnK2ukDcMaaGOAWRVSpNQErIanP0MErcT29Fa+BNWZqeort6RlJ
we2ik6d1GrhY6EDQkdmBgMy08WQHHW1YcB8btpxFZLwRuUHJIIozHPkMIZ3w7TFmy2/ltOfSuO4u
KQR6Qa9xMcO1DDJJUhdPzyQyyvjtC09cxHPltme09Slh7i6RFLEaufuJuoxRsaUyxw6INUlIvFXZ
9+SWsEQ2Bnmn78EH/daeXxFGSlWg2lxMPF16jaP2EmSVKTWoPO+BLKgzbLoowdZmBHB2VKnSXh9l
Ix9KLTqnVPdxs+IT2AtvZH+5BHUHpMdVSIP5JZ7b2EUpqHJP4imAvNaU6U8xNrBS05jk/WZHPzKN
lO0/nYoF6w/GLMebrvUZuHVrtCQfwVXZRIFWj81VF1brnTqYmG0q56itMgU+2/EASqRP2Mu3LOLK
fhT0BBwuVIlv/ZQrpptuXjDi3i3FUgUj3frZuHy31peTbmBD5hWbnzuzFcdSeoJYIMRwtLKhUl26
iWox9a3fp1zzJ16uF1QKq1UlKnm+0BGlsoVyWRVPQ3VL+FTueS6i9G5J+LK0yU8yOT2Bljq8NxMu
WYEz1kr6I4uw2IYxc7aAUIOtCtv1jxSFKX6FRM6HjzWAVgQPmSO5Bbcg/wg6L6mUSYFS0yOwRiDA
zP0a+wmfzZlo38c/empgBN6zEcV9HYkdyzhMDLUCf1It+88H4mSJA6XWZoi4QuGrEEqMLyLVf3AU
ixmBfv+EzY07jnQewhJ3Det/X7UNLCbPMTlmkg+pViE0Vhh6fF1HObC5xYrwSi4bkuV7WS690GHB
frjco5GXlpTiE3xRkC4X+iUapCY1h4sd52B7dRn+YwkZtNa/oHk1U8otO/BKnMg3F7GTm4olilTy
KJ2tgRxawJPwV4MuEpnBaT61jNbVNHskjVeGtHkkxas8wVYK6OX5NUtlJCFg0DSAisWQFBb92OAs
P/1TZJoxtRx4aArHSV+D4P9ffrvKdD3q0N5z0Lb8f9ueku8P53ItYwmt/443W6sXqHsLFczFsfYS
Ojawq7wURTcNJFAREcY5sPwn78qlJ7+iiJzod/heF5fyVNh2XZE4HRJGx7t6KQHaxmEFo17Uqrpu
0NG/F310T8qSV3fpD7n609rf+tyc2yp9qXzaYqKOSDzC4seRKLzSslroWJ0L/GH3VHQUJxeUaQcb
NIIiBgXWuD1zApEAdGmYLpFEq9CXnsoE2G10Ofd0LFTvFE6NJ/6rsjn537rHNBTPIP515mqPHfdO
nu4em/8hTZ5whzzZ80y/nofXtfhbgCLu2ZH74B8WhQg41zZDx1kz2l1qgZ820Ly5s3IORjCbB+nI
PMDv0SSYMO2o7xyhxZ+LuADoQqWAKe0FO7TcDf1wm2Vr0nhph+iOoMjxhTiUc6C/eAC2i7KdARhN
V3CzRxUypz1/BkEM/LJzMcb3QLIrMzO7xfbrUKagjhcy4xypRw/pj6mMPfoWSPfpWmnSr8yY5nQf
Lv2/IUjLUnZgaUzlj467io+4efig0R1ErUwZNprjQDaOHWnfbObbjz3NNDxBHLmlAHx79VQ9gQVk
P5o7I1C0gMxQKVflWEQSqyB8uLCPyjfIUqoSK30MhselxE3VDoHqZ2R7wdBzbojMIHRST/SD4Ucy
ar6cx6Hp983jvi2DY7mL3FXOaaAg5x3iqu/7imUaMVSf2godq8FgxuRaqUaX7pPUHNq9TlMJv8wF
7O0r6u+BnYabXsgnCmzx/AZYeA2HvBo31K9tz20rL713GaDX5hPzx25T+BIe8VKD3B0LMpnN2PbR
SNqAFj/99ePO/jfxCnkZS8Cb8onXsTgQ9aGeQDvCZ3AlHf/+x9bbBg5Pd+xdZpPiGEFqONBwmvB+
bf/u2QBcuD0nPKqaRcuTKzKgOqPb6Cr1OqGsqAMLLjusUsYibxo6ehY0OSnBHoBFS/ZYh7jYZAIq
xS9y9OVC/G6zOWlINU+gw1A8mxOOftrl+ohvOvUDiW3aJybIi2CHqMLrNjOYPMP2E79Jg34Xs5vb
utADFb3s2UWZUdnOymm0jbCq2j9zkN6FctWjw4zsHG3173mKCjERb60mtqM0AWJgqqAhALHaWuQi
6o/FgCnske0Aa8OZ02GkOX/0jojoCp8dF9/NCnBTSpLkR6fQJVP/KBJb9M6UMDRZSxJGzRX3/kJ9
8Etcsg0H/RmPye3xO0Z5qLDOktmUiia+Cv60ivKVePqCUnH54GVcxJw6cEt/mbSWePnYj+Umxr9X
MKcPfAMbtQgk+12TVqngTT3g6wuETNJ0dR0LKZ+2pZT+BTBVUb19bsgImPhi4xh9JFlHbqTDJRgh
UkISMcdBpq3OH1y3EusvMYkiG5geKfSgsiqtxfEugjQCcSAQg+3C6hyQzgtSuyXS2NWwur9NOX5W
yqeZV3bfik9hbJKs2XPTjznr8JiGCiQLBPmELMkkkZksLUP+qsoQyKZR3QrW/shcLNTLUQOLD6HU
An1LAtVGMg40sZUW+dNoDu9sudxcRiuW3nO1DI9T6Bc/y9BmIQ6K/CF0Ym2O7BHKfBEfTtJeh9s7
1tJXpRbmCfM1JIMuHAE0PKB9+5REuvTgJZWLbKdUufgc0Vw5hw5PoQm5faW2eMJ39Phfc12b5pQ8
4gghaXSQmeYUXPfuZsxdN3iVpDw7FepTmaEntpqZgFr2Gzhw0tsJlMnWJ9olVu0BE1Bakz0IfeLw
bRff4JWndX8K/fgnxajpYZiB9Le73UWAUjiXqnWUfBAdoXq0iFWA1tt0cXohEp45TMpY48GpyIap
0+e/hbvksbcZ/hHtzlVjBkwI9xUTMEvbdcr3MBpk2DSdcJJmul0Z9+MDqH/gYlFJaUXWk5+aQGCt
qbsLv4kjZIV/fe3SX9ReItNz0vpoMcSgJwN3nxQc3enNPq1bKSfzCCXqwqKFOin9ErbHn6zfk1qe
7l0SRkiqecAOYVNzHMP3+zmPooYFCogpdD1mGIWSAoWBpjhXqvA9s36oUDFo8KpMQnm91XpKklSX
z0CWsU0lD79PfsoNA2e1AmFnUh1hmKiSHq+mUo06R3oSXHXrcRn9zQq3EfiLFJh0fwBcF9YOuf5U
bh+RlJIyOBgLt2O02Wht1eFDItlG0dLHkXWDSbxLTtk/vNbFGwGDvrZuPmq4iaBv2j25Rm30mcac
xQWMztSFJmTLkwIj5rDflF54mka44LnBEIV/7Sodg3bQOSMuTYWhXUQ4ZH1k/yfLvoUgl5g9PgLN
lNm1oOsfU5fh3769i29TTO1qxwjru5zfGFXPaTm82iCvd00dtXrK7F+8id2PN+NEo2kw4C5inIKB
MV0tQ9RX1cw3vm0jtGY52ZZ81N1sYHIPD0iYsNNOBT+840z4zmNuMTTVOn6e+wPaBnSOKb+3dcC0
rcmOm/t7bSxaZR85iEd/SeDMQ3lxSkW1I7Hss0VC6yeeZHeAe9TwmHqbRSmgny/OyaO4F0yvNXy4
Chdhi51CGKUuSW7Ye3sYSV+tVra712uzDqXhCFJVcP/2J/jJmbS8X5fizc8VQAHOMO1OPYy+2dSk
qNN7oOAxy2n82Wm3tKWu5/udkQGeOv0HeGXDuT/v6JC3ff2eab0S+urtsIQG10tX6+1azrIARMBh
ZfNbS1acJXUcBxHAgWHJ3CZyQzgBlyyYku/Q/QMolUwbQJ2IqsU1iO/cY72T3JWHHrm9FvyhKK/B
yo4Wm4sNeDOFojt4RrIQps1pLc/G7jkLCrdIIisrEnF6tkhozJU+v4uholRFYV2xYFkB3nFR40rl
taqhUmic3wbcFsyh3N4jEFdsFH8ELypVJtZDNAO1395S1+OBa0hgvgEUxwDgfX3OeWqrE4POmpoD
WlrT+03/40n7w8MbcsKqunQt50bCiCTMBTk8plOYIMncr3o1rudK+18eGU+j9PM37W0q7AE9yy3e
A3MtcxR2DkxODVyllotSN2yIVjxJkUS+rmFT0YHETyK5p55nFrbRmb8yNh/+Kc7IzaaqPnHek71B
Ma5/eyRVejlFjZTCa78ee1A8IRLwlMgFPAwKC446WQbxug7Ve8K9gRVHCeCqxiDV5H6H+V+/nHKT
cVl8q9YX6at/iDEld+zQSdUNaQEevJc14jGx8udMXDFAp0If1CdG44BDemr8K9No8+nyW2So+Q7I
Vnl23SIiN32U1bqrHnw7zKw1Qa1BsbM9DalSVEa412T2/AK+qDk0v6rgz7/8/2DfPbWLkoP15WkR
N8hYRVuTE7vxR1Fm1Z4x+Q2/8OrJXGzb9rP8nnxwd3Y3XiMSVMRz1YcgPcuR/1NcK2jxZsvotpGF
cb7V1grR2gxIlTZWuWAEqeXcTYqWJ0bQAfxfE2rwb0i4eDt/UnnFhg0fnujVmHvZPJ38Eh+nT6Pa
nDIpRNVuGOSS7WXjOQHf/ob2KEcZSuDd6nz18Z8NBqnX7jZ0iGIEMFrT1sXmYHWzHFWDCbca58nr
e3NBMOB1znwguPpH6QNIg2JkzsfWZRIR90gaxq5fqBQGmBdZf1ELebanSsXR9qdI+iQ5lmnQREoS
VQ7DLgGQOZKcDEE3K/Q2h8Z9kPEYrh6y3Vp/4PX8P7WmxCULLKIjNSu/Ue9SWcEdnOPIVwLpwefp
EtTP/jF0e7YusZFtR6k2zoVAgJL2SvCcjLHOP3zQ8BAKlt7nQkY0LXW/FKFQvqSk0O7a+IU7B3Tr
95qm3YvJhiSCxd7V3WWkYGRuC4Q728jvpGwBU2RY3sni8xFMERcR9et1P0GuaztOZUr9oG6l8SoH
CRaUS0lcKfdHa+xaF+UKzhRCjs7Hi4j4ZroulvRkIGJAHVbM8tRSL3mChdX2FCRW+AOoNjPe9aby
UytISG4jeCVQ0MNyIfI7pV9uwN6qkywGFYfdXmlFYmWgqGfyrn6vR8wiI3fG3nXGkZAhLZGwoHkX
Ob7K/m+55t9HYSNkCm5Y13bS7J1v9hVZrzaPWMnnebLog3PUAeXw2CHOmEHm2jxtsjiatHRLYSng
gs0dKMwV5XGLYQCScbQPdvaXojaS9Bd63P1BMo6KI8oUXRGWu5A1MDztYJl9z+dUVeHaFhu1cdJw
zQ1yRUWkz0fDNRMqaBStJtzpcXl+gl2KB6KV2LL32TgepFrCjDN+8N53pbPqPFw3lSxJw34E7iW0
uZS03kmaNQswqwkxe8jd8Uh+E+B25MnQFEYXbg2gqvjZsolhjNxMVKKcUHfg1NxZX9v6hFGJjt+L
fgVNSHAY7cfHa2mW1YDYH3YLwmV/TwJQEO+OjuR/4P1e5m4IHMJDHyIZYycTJpaSVNLdmkIU7gKE
3ca2zryMnXaWOAPFyNsNSBB6p2zv2WQBvGTNy3ZlXBdtU9dmYZNxuts2L4eMNyboQj5DMC03hlpI
nRzWeCzOtxJx8T1AW9mOeia+qYx6eyvYFKkgYMKJ746t0U986zyDozpdLLBkhnBO8lEywIwsdlyE
x1TG6i4RtPL51xqnMh4/soEF9FYxpXkNJHrun5xHTZ/pBHFkvvytRHCNrALBC4AGJMDbUd1IJzt2
l3l/uCX5EQb5YffvE7Nt1cDBAXY2/3BqRfQXEnPWzzuvRatFIWwuWu533WWYm7tKub98NmGihHXx
m/xSxTK0OrlfxRFy35Mk0rfQDCsXEzlQy23zx95uQnmzcheXv/YWk+3AKbtqWGTTGpzWGzPugwP8
foyYYKjYahzI4Jh0FTqfijim4uHzC4IpTuoFvomVNnutdw304KZsL22FQdha8xviPwUg629aB2on
WlAtL8HEUurXWDE1xqm3qC0GYAnbr5VQY3G+bcL3upnofAAwF2oc4JZhf1JLe4lYPjj0OTJMoQUo
oNVWcRpndLXNBotBkryYRRGUbrY2aiHNCk7CZTkUhWpdXj9i4kZFF5GXC0ezv082xMdr0weZneVe
9DFMd92T5ARqjJGUjOBOaZsnuQ/HYWugvD7xFliNr1A+BK+JmVxQnID89Gv11QZh0e4tJsuM97Fa
SIK0ndvBfGtz9TXmD1jpfhKqPhr60cVSPvCV1stg9wd9gi2qqimAGLlSitzX84dZ2+r7CDzfuTpK
vtf0O8j+CzbXcOqEjSB8dgFm4GN5FuyRgGWI8y/lTSnHvJQq3tO8rcFLxz2+QURc8EbQTqSjx6Dx
gWS3GLrgNLBy163mtAoYdd2EtXIYBdc8LzPrRmk2FHjTTYrB6VSEpMBL5VvYqt7lU8gLNODYrIP/
YhfEDp7ZWpalmnUyoYMqxlxWi86L80NxxLvZFiOwX2G641Tpy3P39fw0aBj7GpdCDpRYV1noTRYo
iXeEqdOXCZGz7XlLLGjnmc0E3hWc1G+oa/ERrVwu/VWY7bFqBpoXtFNcO/4SA1lPHTsKLsk7neBQ
3HQHKGCBa37ca/Ru6JHwo87fnEN1v3/ikr5JZjJhkNgZHnxgViswebM+0umEzucZSlAnH2oibgDU
UpGPXgtybNH4fz/xlD3R2fwLO9kpEvWOFnETS+deehCzNYqctoU65EAvIujX8gIe6AZxuQlWnUFP
3o790Mptxw94afaMQmN6fbjJue7mNYE6K/IRWPei5wPtSl1eYttH4U8FujSeCrTSvVV2ZTo/uBee
nOcufqenw3tz8lubyHvpC/3ArqlVB/is8Pp6/ao46p8m6inuJ/vc0zo73kCvRhk3CqOFLO10QO8t
NH6m14wO6JpQqNL7+49YbDnLiXsIYpGflWwL3NQHX4faq3KoVe1xBXmtLbEopGVtcdrNoIg53O9q
NU8s767ifuaOZ/AliNwhrIjfsjYovRkIEsUDUE2NYAuqJt64pkUUI3TVoCUqmMoxLCgktZ0AWDIZ
wgBILpyfcPXiVrYo2uH7mmTx9eE/DEbaYmnVhfmM3zj8vKLZ9/Xhc2deD+jEVeWx7px3VAiLsyDc
rT3ipHM2OOJOvQ2R91ZN5k6P2v2cGLTBHa7Aft+UZGD+8AQJhW8m6OTYN9qceNLyXTLi3+LQJrLM
BvoODWlLQTCTqC+I1/bhZqUIOulq7rIktAwFcWnFoNRJxEX7o3513DKqx1ZMUcgghdKA5AAMxIYw
RKbfHBVFpgZiCucX9bYHWnDKeW83QxqcHh31/X+5y26xiexG5RV6IDYZN9xwdpu7f44WVApQvQ0O
a3e0zRc2qyewTYfzFYUOC25v77JSt4sk0DjjZKFu+3hrgroKL3ohzofS8wb2x3Yn57UC9GM42j1Q
uKpijl3LuYnbx/wlqloBHTTuIlGJMplk7NlzFHFb963rTNeXt5Vwgp8VL/6iNQ/sOhupXT5kI7g0
PIO4BNry43fGyyhLSC+sLufpXE1Ol+z27Ff7Yf/B0zYML3/2mCazz5rULdQAjaIKZZQZ82y+GcUw
HMr5UZB/onSd9f2wm1AoNse92Gb5g9Gn39p4Rh4MNUg0lQiTssQD4cFNJk1x+q1jU+rsxjrVLx56
tFdMv6akDkUoFURW4k4WZKIPTlO1ALe927u5xB2OL2jNaRT7p8kf9YOzQk6vNNxQ+9mGf74GH/o8
wr8Lm7WaUVpk02RjOjpvKl916Ga8RP0DG7F+lCZZbEQCErH/PYsfroeDAQx2/W6Lr21c/8Mgbxzs
w93zNqKzjFY4wE2Fk8AFlhevPH7bXFXpCf3T0h8AyrOWkxgF/AOexmnoloJyYO4m3OQEj1Pqy++L
bd9kpLGLfyKvZJOE06toZC5dejgOoO6KwS+tQfE1KWeSLqrpaRbst4ZqZM+5vwrvQWxPGe6eQ8UH
pFH5cWNIErkw65LGKZZYAUS7C4PVPaWIbGyPlmvZNqYNPPRxi9Zscob1mBKYHToYPcCZ6luc2euD
f628WVNpnQL5fQ8vbe8wYnn3M1VaY32eAHAWMeutZqkrbEsMEq7zP0y1KtihREYWU1duNvQalCvR
eqxhu5PiXnN8h4boXDXrl+NmWmCu+XWZw8703jfnvBL6EJxm/A+bphJdrcWow2jlXO2ZaZv7Dizu
GtsgSwuOHflh0WXVkHbt+E50xxpI2WX+WQHPZiNb/Y6KknD2Sj6ZtAAl8iwlns2S6S9YEc+O7vKT
pLeL+Bc9hueY4qr9nTlUJ3codsTpChkdTVeWuwcqQShO5AHWyE8XnleGUs9curHWbutq9G+uBHd0
LfqFvQNvyhHEH/ZKYdwaTiRNeXaOVTCCQGbpB9gGzUMwryNhc637b/C8g6gni4to5kpfmj9zo0Zf
x9Xu5ibgZju2zwKpy/woeKOg0gQVfOvsGY2rAYfMXFiobHCQhUI4m/7PsG2S37TN4oTOLl2KYsTc
9mtN9oupPGOup5VtcKPdWGMQtfQRcO3H8ezYTjCv3swX5C69d5ocJsjVlwi+5KIWO1Fv8lU3mMTS
tahKs9yswPxeJUzRZPbFkpyaiKgAQlyRMNOy0hXooXd0lp4h/lwrdpf2OYT4PnzfYIOWqiRuM/Fc
sVPcvJe5FjiMElW9eEgzufwkTRVmZ+1hOelVWYx9eeMhUolKgePWb86uWitJ5l83Gnryc3XYAKAR
kcXC85VZNeaUz5pbT0JpZduN7M3Q1+2RDR6hiwwlD9KB89yJscAD7oNdz7Ehn/rEl5g4jGONZdtP
mlK5jFZTBx4o6FFQhZS4df2EPmTtuj/aCWpQ25ZVsI2nfmCAR64EGNmSb7Oxx4IE7n+01GSU9+oc
6fopEzxcTV7hAmWLgbZCNe8beMw+6mkzL04+/bW28b8wPhBPWTXZ3dYgeVroDr06RJthyzRWhBNN
P330KwiTOodsqwRnRhhrHnZWI45iNO3sOiX1Ryh/2Sc3I9qZGWjbFsWuX6EDWedt5X3AyUrfZSDM
F8AzyLlL4GlXM8VkSIvUU3xOG1EQxLvzyQDO7b4Q7xPKqKAEaJCoABcTaNgVqlpZnTIeFBdJk5m8
mOoVobIoUu6aU50W73xMZh/DYIvrKd2pymNwI+VYR6x986mlc9ImGKgemo3Zfdb3xYHzG/4OQ5Ta
woe6jSqrsig7PmW6/xyWAB/YDmN5xXs+xMIDS5nlh03gAWg/Wz6GNQVxgY35wPV8VZfkHXTEejIn
rV5orll+HIr6rvVx+t0xojB9HzfabCao7DfpipNHJhCcvMCvHsdwsAnEnqoTL0PVeLBUhxEvMcgO
tp3ektKlRP+eWgjAp8v53un3iXX2uRfDBwkwLPAymYKVXspceeH1ErQfUB9HQk8bozP+p4AjHHaI
RLCPWLiBL+CQgiB1I5I/zjBlpKZRxlGJX3lF2CPDufs927OiwiJ30+iVINI5rcK5yIvGHAL0D/f1
MgxqlYQe4wYCsTkmtenxxKzYSIWUpOYVpFzQaybduNyLNBz9KJiiTIU8j6n6HLEPGLDVaY7fvCTN
z2M0XE9Eex6Ynb7pKvjbTRBsrqir5Yv1Dyr/Sn70EZ1PuIsLdm8wpxXgR3R6CneMaqA35FLuDQ2/
hkdTyRkUFqXk7cB9/lDjY+quKuahIF89kDIaa7yGyzXlMmWHQdlaVtg+SNA+1qwRIeC6K8FhpMbO
3EC1OYd/Fln0WNvyJHBncxfIyuiQkEPMTxlPvYfQEYmZGip3IlZiwYlnI2aEy5/FtSMmw6fzFlLe
tZyRkbM8WFUF0SZ2k8eAPH3RV1PSt0KkOo4oWVIW8nv0+d4grDgYLwbC74cmrgNl0UWjZzaoK+hF
53eSB5gk+YJxFV6oPeGPQ9joEpxyFfa8f80bKU22XJLK+RzOWjVJASLG2rjVXVCJAcFtDuZhU4m+
u+XeD2OjIzTBb2X0EHinfAd/VQeX1mKx9woaA17/7p816sFEQx80xriySaIVpMpQsuadAukqqcXX
hSqh3ZkPTcWT3YJT9lDe50PNTfnlzwvgMRDNsRFyCGeFWRRbGFYqavDzQwwPZCLRI+WOmH+K+ot3
ZgPbOq5NtuIaco4bzn5whIrXBueSh04KTJVMnFHXH11DAKUqhMRD91LSyu/basZHiECT0wX/ASOF
+U6stCb67UvmIeKwttjaAGu+dnEMNk105Pb/MwlhFSmBWvh+/oDCRfyCXABS4NAs3P2Ud8eRY2F/
Ppqirrcz4M6ErC8ZDOglJnrd5CIhjiD36D/uPeSw8axRoEjCrLbUHJ9NmwhGjn3vbP0ysWLHONIJ
leKapSomCP3MrTg8K0nm7oFAJSnBcG2x55IKl8JdS5iVO46UazFWsiyc7YQFHRYHPDpJuC2G3bM3
SaHOrMKfGdFaDQR6tqexAMoJVLQbWk3MbKtVCLLgjB+A+qIVDM4vWM41PD7D/rd4pe0hFBJW1NLJ
fO87+aR9qMWtw2e/d8RiBLy0JM1q0rgjLwtSLwSiFVoifWuxwSUOS9h6LhD2L/zzwYCm85WjMhqP
Y0RdgksIidH5i6+S2d5tT/G82SRxN8NeQUc/64VYRwK0pifIqQi817er5NZWbHBfuEziB1WwXsoT
MwVmlooj9P2+rc6KUlIGzknKir6khmS7EgpTJWLH6SDJMCOfZmgiNfhE1cNULHDg8zZvYus4ijUh
ZIThqGBKLp1J3t5BhpWJiqZr+VAvyAwtpPx9iT4AmIslrWdfZQTcZemcnnUDqaFKiUkCXvzHUMJF
z5ahBq28XNUQxZNJ+0uRw4LtNA0+K9RrwezY+Gh9O26hzmTiNx1XhOowhMx0EObZZBZC7d6mMcyb
T2fk7ABe9GURPGluCGanBUlg3DqXhJ2UHgn60S5Bt6wFxDIfGuI7hQh5ydbntEAC3CCIJv2JZ0Po
SS3p8drK04/UuoP7XR0VroHsy2yoJ51Upt3Nc8Mfy2b9tyMi03ob7klXNkRmpk3z52bEaBwuD/Fh
L6d+etBetKpRheESdInWp+R8WVSnsbTcFGymuzelqKagX6QnibB+ZbHAkkYDH5AbwETTH32X3VuR
JbqQLXBip9LVESblODoESwdgP1pNOtGdnQkNWY6ZHYRVisp2IFnCRfzf+w0WCz7QnJPc0/70mLWo
htB6prHB0Nzt7akKN1OZ0Fk/R1r5UIvEVXix2H2EsbW4NTkEct21vDNMSC1cXYwAYDYXvLT7w0ML
S8w/KqM4ZlGSn0Hwo/DPPmEv8YvBZTLHHEI4Av0pfux6/UDiw/pU+qnin6VdfFxk631h5B91kliM
KvUm/LkcZibX5SzhN4SOicbRBxeAIgXsAVNQj8lSBXZ7aFwK4AAVOolRGmcqJxOHjwe0MaiF7jhs
m2eCk/brXuyMyIGRlIfLJdGUH4BgUiNrLx75Wbe2x++NDtnQTU6zYlY6aMy1EBbLV4rMOfb2eSki
5jliYfAByaxnXfgFGjuYVYWt3nhlVE66bHVE0c6/zayHTPeyTqBRX8doMNymjuwTB2B/f/sGv719
AplcPQSVhkzKqKp1CXKWxKeVQlvsyRViexiDVJ0g5IXiFakFxIg5OV28kwtOBHU6fH9yu+P5a8LP
IgjOkirFU/kJEK8V/QwG1t4byYyNGeeBNVGMA2odazJiHfZRoefRE4I2Roo3AlG5r9HnE4CN7GpO
vq8/McdJcMvAwH1EqK43eQ42dlG7HVz29zoB9ZNAan9Dtnm6Ch/Tglt+IvrgxpIWok3+c+0jPVEC
UsiMbY/ySlxYNVPwZqLpqHivU2Dtj+RqDCar84YQpYs1LYXCBS2PyrRRwLueVvblFP0v2Z/R2Quh
vkGVbbd8tR4aSRg8a/Y+yql2qMGm7MmJoSiLv0SWeZlE9U0hsD4kIdzl1v5/6wXR3Tnb1rDA8Hou
mA/tiw71YWMKaNH+OcskGqP7NzIcOtZmcDrMocfUT37KU6uqKprJkQZ4ikFdACWQuzMej4G9ZM1P
yxMDEiZzVUqZ2dto04euF4r5Vhl0PbQpjR3/FVGbmPN2FXu6/Ta8xi9NtRYG10+gH7LPFx7DyvNh
wZkKB9A91BmXwLyF4kcS4uOE5wSGYakrFwWm6mJS7hVS/8acHiFpsdEYfGfvJI3moVjCY//rZ5HK
qtn4yRSbIgJlDAKJ/nJ/xhnK4WZyYZ2TvgF2fZDMZCrBgRqNATT66EJSdG+bzsmlqOpxtND7i8VP
8jfL+Lv1+CorFWxpvRjiM4sfW8zxpCYP+rarfD5p4F9AXI7FfOY1JnQ5rgBp9B0TotyNhk9Hc6Gm
E9SPGkKmMU30WLKqsUViVh+hstPrKurCQxdr0BG9VZabLj9JiSqRjCYMDHyyrlyBBYqBPQ0bTdbY
884LdBQ11Uj6Y6OR/uuj3CzeGHBq4F4Zl9qZ7fH0vaYG4/Yl1etp3T1cZghBWVYKrFmS2xkBSDPC
rK6+xSwsTu3f9DEKb3lzhIv8oIX9tvPkJXVcOH7g5V5oxDZ8G66y9hJ5XvlCxZQcNCpx7SPVBXV3
tyDE9mvaDDrRbJTy2CCs8l1/LCOUNRw0dM3+VFdhgY4JQADRGCa6OBwBUewCvnfIOI6BeBAl47su
N7z91PeUqXyLVcn3qxR7xolbso15XfLKe4n+mni/00J5+ENF5uJfspACABzOXsjofBONBSTHtMrk
PzNAne3OJ42zDpU6XmldJiPWh4CDibAKwzuUbiP2aWCvQnceeGkQD+YcM5/K7F6t3/NJphT1GQf6
n9LDx1YH/9I2SfaSXpUGgPlT7k7/1xx8rqLBMVeeh5ppLfglRM9DowPMY2CQi2Y3NA34g2j7F6mp
jMvCjXZ6PmIdfP4FHKn+RjeY8M+g8zJBXsR+gGWkeekSKEEBQ6yofsrpAHoH1Hh7bvDBEMBUfIob
BmPnRjOY1o1RGUj/lr/ce1xO985RyuTZspLdnYNYS7jq+JipHjxQGMokitXfth7BBjLxL7q0XrrG
hBW/mfXSYgJUhdX68sNyjnqA406mVV4pM3PcF2VFGC28SQO7rRTceOgU0eg0W6sbWohADOs2glOY
jOPSDHsGUMRt+b4j4COI91ZuRrBrxj3XK0s8BswpImFVOflmxPwhPdeO6F3eb8/aTrVDvBGPMIzi
9I31kxtPmfEdUkzVDu+4AFU3LSmboUZQVYam2+7SjTIOAMIvFKYEw5e6SetETR+5+hEPoWFlRCZ7
Vg3Cu/t4OEups5heBmz9wk8qSB4dRhAROxjmjMHap7u64Ngl1R2z3CxCMyeGcoMTrRbNeRhwzLdz
UJTpQd9MUajZ/AptTTF0cIJm8K5s4oMB9kEo0nHHPFVNDumcVAniRU/x5Gp6OPimbohCEDzUnsDI
lvSmKbYUU0wjNQbkvYZZT6SZh9mJivS3P/8HJsKNe/sk8xMEVnneTwGY67jivJc6bjgYXkDUIp7G
tZPX7WsV38cjJ/i5AXc9NB3h9W9yQ91L2+kJ4rPqWhLSc+H0ut79Y3+ImBQ0SOxz1xVdhynQvu+W
l2P6kdek/NyphKr4Lj9sX4feHwZmIEzd3z2oNe6PjFo8xnR29TrTEJbc7bZf4ScQK/arwOsckPAp
mYJKa0OJYTrpGOO+iZww2pbzU6VTryOuAEwNkLc9HKM26D4R8CnbX9a5fuP48R41nsXwWyNGVpcz
KLRnfALyP4iEVFHcsRVEnRwCj91zVKLtHrgewtkoQ/9XFDyQhIUBoBSYKlHqjtT8ICnMT+khjpKz
COp4qu1B8/0nQxcy95kJ1FgfKF9d5ZzAW11QFst6qmZpCQ+ov78b6UO+KPB8tqxNDV3GkpHJgedr
vfiYZ9LUbEEXqG8jTTxMisDXKv/f1bjO/7ekPT9ig8EIzFiAiMQqx6DZX+zYQJRqO8dWNf0rg5YM
JG8ngPxGCy7XK9s8M1qcam2uRI8gBzuO3d/XUsm3rSpefz40+fe7AFtn1RrCdlHh8s3/5cTzbFLV
UMPpfY5mV94OgXw9i3cKPWbMq65OEf9KL0dBhIfHdwsDaKhIjhz09nZS3SFxJnIlAvDEYFPxSZmd
eOPDbmOibhFMiatSCQW4WkuHaDi5dM3fh+Fo8YQGko+SYMJbYnaZBW0p5Wa+5d2wifYvB2xKPMUa
7ZqWwoXg2mHG5f1bGsYwW/yHrVLY8lbMCgh9IngENhDfxMoiJqJcJXGkD7D74FRe1on1TkZBYTx+
2VBRAwMnbXcl4qkUTINIrQKBmkHDpIQ9XslYwIlF5jJZGQ6OeBuw02og8HYWfVaGbyu4y+DWckN5
ONUWLruOcTrqu5sAS8nowOm363flYadB6ngq4Lk/oGBbWiCcFEbYeMMwn0cx+GDdlY8MF7DXepgO
ARNG6gEAoSAr9ZQM4XC8uoVBrRNJ5o0fqHjqzr6zrOyZTSmBMZbQngUNaKsAOPw+5859oKU3iyzu
4y1dgEQ33IPEw+Bm3lPbRnv4NxYpMggguGhhdodTlvJVty/IPLF3T3yJv5OUQh4DH80A6ubASWBF
WlWrLSkLLwUdp2jbN1Vs5+ieB/m9uDsAfdzbjVW9umKb1QV89+8i2/rN11vqlypA/PHKwlbq5IA6
7ZBewoszKJo+kCKmRPG+5Vv2cqL3CZrOYGVMLsr9XcuNAtk0ePTz9AYfQLxVj6fGgFzmBg913Nm/
ln2KXmdYCpmtAtnyZdXew3UAnlb0MqGIlkvpmeeRGbwNQ7SQn61Jp9rSbk2SN6IgnAvmV6kJtDuM
B0AlrhwQe+2G5lNcGPxSlF/AbX276NiQB7gfoi/hJHwVaBCFZTV5mBIvpaVPtvNzkJcMOJnE5ZvL
GtwaXmoztTdNSs4KyAMn1X8iWlwMufMSPazOPfsj+jTBH7B4TXK+EKhk2m6OmJRWJvtFv3Pn9Xd6
HScMlg1HWe9P8dpk48zTvsWyrCnDdbSEPFvAbnPpnYmTBfPhSdmNpHyD/6QL5OOzn0DzbNpJSwQU
EVqRP7prkH2ryvT3acI7qkypqVXFTyC3zmFGYZ6eaZQJ43OKXvPjb3ReYRTNuGqB2e8wpbdcE5V8
68LvKQ1ptYaojetzID1FuTR73Sz+K/9aj7dly98Pa7sBUkZGWJIKtkLrkK4qJ4xXp8EPX5qj69OK
g4ZqfVnIPnHHcn1pjtvceuMq3O4GBw0hSV/RFTmj57B05a6Q+3bRILnSiDOnOiOeJq6TDcnnbXHm
qAhnYZGnqsgC+gyUS8BJI3b4dfBvy8pfFArDy7GLmDUaQWspmUJSH1Y885Dt/QLhuZ5ioYT7WATW
g52WnNvFste2y8ocnMlmvvYvB5+7Pr73TS+dfl7irNz04yhEZn8vAMUqYmBNLM2oM4Et0r/8UNqh
UVaVMfh8AJBeUtAIxZnrGIzUy7gJO/LLeLL/s5bJeLKaOOkq/dPUuPDAoOUcZDojESRL3yWLkxBN
QiDgCwY84nfJIwnwX9tcJH5Y7Vd+lHXf1iATrxWA7W/z1hJF1TioxXtls+6Le9p6ByzxzUCZHDN3
+uuvN+CO6uPlfPZcSousgJ31unSHpYaXx9dOMJoKA5WnL3NSgKFtf0ORx6cZJXIzUtqw0BmRsNDu
mk5slPfLwWt43Bh+k8CR9YE7NNNOMnDlb7O8DxLFQpE67Q+0sBmhuK12mpxchGGhfX8+NrPx7s2w
935Ob4Db8tX5mXSOtec9EG8RnFiGTySqYYmLK53/kG8OdDOoepTRtcTMthdhRO4FVQz0EA+eCOZL
924TXo+qxptN9rSgGZ0NhlhxxFSIqj3tL/n10Esam3c2070tlDcM1CAD9cNHlJWkhujFsmVL96dv
z5NnRpZCILlhhZOjVe3c3LwU7Rhxv11+Cy52NlRhEWc/sDKXLI43mdGKroBwgeI7+kiL95gckV0r
g5HE0zVXi1xta5Ux/CDej8teXYS6pLgYIWzxOX75RSYtYZSvBZ92NKirMCqyIeA3uncRWKKQnEJc
EZ14/NyHnwR5RCooISzLTKDUa2mVrHln5oK40A2SKdL6eVEAaFvSLEVE6sLfM1hBrNt7EWqQ0kBz
/b/+CPAGBDIjlCvC3uwk/BTFoZNKbWHQrRoflHDCPETwvSt8Y3ZcYOD+tf+CRpt9vdR+H1CPUmUE
BgV5OJ9HwLYAqKQ3MBSkm8vjkhGn6g7h4gKJPga010ivoTTM6wlSjKuIz8IMoYIR+h0px9zH1UPo
jrthK8h4WFujJdsEWCwEKEctgnp1B1wPH9Kvz+VTUijK8r373k9Mga4lEcrP9bYgBhGSfEcHqME/
VMJI7ncZrMDqSnKejc8+tbr5wZtw3bQxQgELwSkS/lInQBNUdIH3w1AJ5Klh73w5DE45HoLqDnpj
tvmaKA5F0QyNGyG+mF+kT79I2hMEToLyXLXl9mIxSDxNU010eIjdwvyymbuGYZKzVRO7z182tH05
SGSNhqF4NYkvlea/F5TxK8PLaGtC9uMzm4aIc8JRFxSq8MsdGPjbMIPnYBhcKN5lc9UPGXiFuxjJ
kqvcML6UYlMjFC7gACaYLaJBYlrbSFeXakEOAXVwtTfWhmhrpMGm3yOUeLAeKstGIDoyiHQVa2W+
rNt9yGh4mBcO/EljyPpqMsH/JpeYcQKHxXQbx2NEV9oL3zlyAwOrufjkgoQO2bLNLd1WZKcjEEBC
7YTjMRNZHK6SjsA6/ho1LBOeCvindMMRh7Z3kzT1vXJVpf4zQezEy6LwjKH/5buXuvgqEd3sdMyV
aHzS5wlkhOdemd6Jnsus9qlEPgqG9rQzfbzTh+vRZig8cPoJ5QTPYYiPGMtTF6sjLPE9rkszBSZ1
9GqJGXNHifRYAo4tCV8B4IS/rJOVgDrrdMP/DE6IMqAAx21pzTNKhXj6mvde4leIomPL3FM1VU8y
jWTtCBnj9xdnqZmE6PByoMZDwPDWBK7UXDyUZz89iYhztteXRkQaqOp+jE6A314yNAyOSjaVZxHe
3LIlUsHPdpyyU+zFmnHkdFu4z+tWbqhmsLnWUoZTRfris4mynUIGjMELNKDNcksMz222CEoydybS
xMXmjc3/RH7mXgpuyLeoZQo3ZTfXGyUumffz3VWKi1KlyqJOXdW5sWhIanqp38J88P0ySBKHeXzw
2j3E/v9u3XIWuxMqT9y+38wHsWiYdFubQz8m9WtEQtd+S7QV+Aoq/cfKa0/yP7KEPNXGP6oeQOFy
7UXAGzYJG1UmJ/fBV/Dh6bwsbZO/7QDD973cwzDL8Ygjww76/ISUru9Ln34nciz8Zv+mJx+mYfcs
tc5vWevsyhiTXZS30xHv42VknIX0csI5XLcVvKYCH3HoFNLfwMFOl6BTfFKgb5bhbOmdGxG8o+CM
ERrYaJgfXSaV/Qa7j/FVhpWtMK4S7LSzI19IepqJLbmO/I1RsI4c9BSCfL+kxf/oxgWxFd3E+Oux
lXsXPOSbTblZRWK7iRG8UThXsFrsgc+8b6gX5wWeeYoonlmcbcLzvoJ1XauU/DJ1FdNT0giYCzao
95EZ50cLPr8i5sUsgn0qSL7K77Ee1XoYtTc1iD9SabUg4An268e8QSYglOEoTmIydpInTtD3Z7Zi
qYjhwQE2drLCiX0sXKBHeSWONZIZqldd2gWGWnXM68Dh4nweifi4JUzddNOY4tNxxZtQLxmw7vEG
ptWIDY0/tbKNfhMCWAxql4SZ08xnlHfuajRRJtRanEJD4T0vEF5wMhUJ9mxbRw0Qlw8vHtg1W2WK
rHUOPJGLUAgsxQyxR6TnekzvTEB8R6Y8XGTZRPLZIlHIOFdda1OssUoh0acNw8dHgSWmbBO2uZGi
OBJNXI0ri+T7pttaijw6iEH5JayU7EhCUdh1SPP5DiE+hp0CsNCy8rAM3bFstFCnmNloTw/yWaJc
nZFbZ6Ej785TLWIoFYq08eSqN9EF/dBUqXL2jhXyrqK4704yI58HC6wE6U/WDMjjOqT/t2Li/EaZ
xGeEEVsRz2FP6zWVPEpfqQdKhY7bf9MwuLjaAZYZchLD+nAUHvGIa55TtMtOQRnKw0juaET2TewR
LCgaUIO8U1SJMHCPVEOwXy0R9Wja+g+IJhCaSIpY06gi8Iz96rCKWGi3qJgKrL0AAPgj4F7lgKdd
XKVbI6WUq7aXX/jcZkx4c2eIEA1pqXEowugs11xoFxL3nMytT2lgiFBVK7PNPBuGYcyDLKsjgxNG
+3fpHVKQtLR9J7Jrmnom81RG7Jgpq5lFzzC41WLc6mPsMPTUXZfYwHZ/rW6nyqpKEeOPLnOtP1fK
UrKuE+3tAjsZH/IkMNIC53jSn2Lj0XEkM7MOIS40s98S/5c0hCHoTkHws0KofnSl7lSlpdViaXIT
Z94FbrBNY81NAKGzedYGOQM2rnZmJHXZaqYqubovDXcojk1W3o8HldlJQgcuLtzFn8jvMOtDJfxf
KJLIzUobihL4p88Alg/EtTI0Ezs6T03BgbjZK2WRHgNy8x0y38NE5nL7Rao68PPBDz+sZD3b7zen
gy9suML899b4002st5w16AVSYw7+gZtstz83ySo3HMTc4fvpx3ljNw28zktSwqdh77jhqh4oWy51
qRbi5vkW6GY8f3YDRtUKAmvd7JMRZ5NmhzH49fpk3r9pWP29qg92B14TMpilq8rVltpc0YQsP5vg
1w1xYPYe6X2o2OyNy9Wsl1mrg8W1naqDhjeiyj7xFHGd5Ipasw/QA8RZsZ+sLiKz8s3jPLLPuh0G
osFzn4rdKxQ39uvSZwemVEf07gL79nOW3GdKDP3isEGKez8NGLCglKKLB8gufxH5yH6XH+Sh8OYh
m6GPo2uVL8b1nxzBuEUN5vZbnpOTFIlWq0cMpmOYH8rUlgecBFJmuXDCPgfyIp141gZalS5XPcnz
/iAcLuBNxiFUcNsDXXTxtKQdrCyTjxLiXhoCNVV8d0FCGR8qin/gwF3KMbNUmoCt3LDQrOwctgNn
cjZ4M0pLRFGmBTDLIGS5vIT5SRHsDBWmVlJCeqBc+cYC1PN4TkHbs+yyiVNQkyo9YmsubAK/z3d/
LkhBrtuAp8RcroW7oi1D4aTjZU94/d0mXjT4PdC/FhOb5NGxIb9LdBQz58fU/NStVXczXLtLIuA0
uB52aB8XWmhj9YbmDPG8Cv3h4uhdh/M4xSFv5L5nIiSXTJoU0ZI5UZkRmpRKbHK2OxSLuLVmf6im
ZjLoyjPZPnc4pKAoXVublXdHPTycdpu6c5+nBMP6swWrZdMMY/C7P3ZWf2BxYJC5DDYsQwTMqEjF
p7yHwrrGKMtZhhSNv5vBFGZruBM4Gmx7EntYHxgi0OY93csghOfsnidXtX+wPk8y1YpRh4TBvDtD
qS5Q5rSPDzbsdkbFiVljuRKbbELW3OJ1yOM1BBp/v2Ku8wMYP7wVWr5V9As0fxbIpwjP3QqAsbDa
o/fqXkWSEnuXR5hw4kS0s8NmqVOcWielwIX4d/75N4fGaKWYchD9QIzLJnzG32afyezLF2rKFPoT
vT8x15SyIBWd6HXhsVsq5/VkJj/w3GqcMtHFZF8yIEJe+V5eprJeSdKi1dykG7le6xuLi93z6sl/
ODkTDs1cUuS3gV21lwmUZnqWN1UcI9CEK+My64wXgKRMGcCo49yKsOBgNOw6MSPyeMn0qvWyjEz5
cOxQ87XkpWJksI8HdqBZa28WIdf7gu1qldDw7xo7GOBFv9mxQIvDuPjJLBhRSzoNs0ZjBr+sudUp
tDc7UbKjyIoe5QS6vSIZhMQAVxZb6yBsVtxboz+bF/AX9ChbZgiPLdxQJgHoyYrltNL660y8mDRb
YpwfhCjmtml8S+0sS6NUpBvciYlxZrb7mxCTvgMjvyA7NnKI97y4YTE0wAh1jLyf2ADHbGJYBviV
BLNwrQrUI1t7GCYzlxdXpK5+J4+eCvvuuxyhzFsUhJ9cD/Bz8nvNiKlTWhgWryM491UgbSaV62H4
OQQkQgEFdXe/U3qH9kfE4MET40OZsaDZaVhmr8nUVDnvbPjRwK7/WQR0s7XdpkQl+jJQjdpws3MG
mJItgcz4+hbk7ICS/vyzGBjoYpKY6vbnvLf+vOZPj7dVtVytk4Bl3IHfWoJI8b+zSLtdmWgJsxpz
hwozwb8OGXIg928VL8LhT6qbtrsdyMkFMjWoXl2IDFp3BQHmpe0TMyymlNC1yDe7Wu09zQw4L5/Q
/V2nz2+HUWuGNx2rtIFRPFQcy5vyIrjYpZXFBQueV2jlecoTQhLiGr83zzBk1M04cEsJ5G37lLiw
FjhPVoxl3K8z7cd2K0gvC+QUPkVd9HtedljVsLIWyBXHUYbltze5by2RiGvgip/Um815SwBYLrAj
YR4koqq+49utlIcPKNWpXVZ7PINetAONfYOqW/vjUJ46zDsLi3M0r4N2W+5h8xm2C3lzuCFxrXxX
HLH/Y9vhrkha4PzM0HIvErKifsLJ1LzfICKL6p0bsMQqL8hhYMsohC72dbwnW+rkkbB2xXWLdmA+
nTwpFaBTm5xlgJLZWiH6dEADnJU5065fAd4YkssN/meDK8ugqyvGEm2eAwRMDVAV/EPD6/a2vQyd
rrjh9slhwu4jxj0vbvi+s5zvTJ63lTxKOubsWVRxfqTuiGY8jr2zWWxZNQQuha4leQqf/X9fw/NZ
A5VLq5oQgziuSi6J5GswwN98R8/4aSsiUhuBqEudGA2aCa62anQd6DjSdqbg3QiC3mOcu/Tr5bZU
2Ya7V5Qc4PRX9tpnV+PR+uBxpJXGn/1D5IUrW/rRwibCETJS5WJJgrQESU78kzktIbi/Izcqe1KA
4yjLGA0Yn/8nYkA85wfMAd4Ok6xJ4Tsf9zD9Sal9kAXLrivTmu0W6aJs/nvIDnI7hiP9sqpVPwvM
TPnogRW+yWX1caFMHnBNl1nf2XYo/ZQlZ3B2fVpwgFunhdoWz8yAhFD02HZ8EFB42xqHzOZEaI9D
pWb6VSiVR22mwuy7XBdsrikleCRcF4KACQTnxGzzCj/z78w7H89GN95uI8FJYyQk/osIBszAcrvw
C+DuID9u2OX1oCr3bi8mJTD7Se/UflZxwoFa6h/ejEQBAAE7vR6wkda3hT/An0HrOpEMqTjq2Fmg
wn6J6QIegd7yGxwf85iNr7uGZgeJZqW6V9icb5VuegaDetF+9qyYfpEDMMfTt8YKwvFQZZZuYeiK
Iu5F4muWJRdF7ZSP8TFWCA+omxyDFYHSD0lMA0JKPw/AjJPv1iV+LqXMBw9x2i7+0++tjl9zamzd
Mq5WvgWfSJsuTWQ9tbllkYUK4j33M9O+CtnmAepN0NNHiGs9pTyapLm5TAHFW8bq7F3gSoSeDCNe
Y6Xdqgt/6MvvH0Ot0Z8jKqzJlogwfGJbr4t9MOfFzDxYQ95+BXeh37PaYkIjPEXh5viKK3SEK13O
NkQ36B4I10atpaI+jMxq2rzww4nMxiUGu3neD059DEVB9+dDLMhWWlD+IXdszzWIyb3jwV4BZjX+
+xKiPxmU2YhH2r+61Y6zPj/VUu684Pqz1EIKyq6iu6yRYHDXkkh13yDXWtk9djRHj6JDl1YtSOed
4xJEaiRyzqywV2aqB2yocQSYF/psvKz2lmk2Q2qA9zcBg3+SYLDTiAgQJ9rlHJnNs1o5e4dM6ktA
1PHqllQeCc1EhXeixueSOKFkUnP868mQGbrRFkFX3zZlIMB7fWFwnc4IWOeLrqn/rq909iuyyRn/
axIH3GMDMe5Ftdc6dZh+XwqpR/VCHcKDt6R3nuNfmvQa80iVF5sKDxgnr6xN/hjmHIRfgp+FIurD
jZt+YrXSUTNg73q/ixdXwT1QbeuJONI/+tmBjxHmHr3dLzxTwypf/ml1X9c4M7rfygrlG08j2y+h
FzHvdBYXmTVkO/J1kEFpvlQAo9pHqQFBxWFXif9gvGkcoHrcFsDMinSLvpoo92FAWesV+cF78n6Z
86Uyc+ghDuJzHSBpSayusDD/gQCgLfvPThpLwzCTfo56OanvQd9LPeO5IHqxyRAv4yDHXQd7FLMW
2hqsqL9EZFx/H/j5T5QtrLrKCVQIgvyXOclGuVsvjtnwb+LNCgsDjCLVynFsbCDMtJgdKPJwndyn
OM1RqK7wnrbsX1Ni7NKcuc7+KAyY3qOFVhxBYZV9ZNAiuHZ6zNN9AQbT0p57m/rPMkwV/OkHeZyU
HOo0QshfXIYWGF62TqGKHQTkpfy7KBxeTRos2pRumH8e56kh8gzJ1IoQG4vQuB0ERlQHgQdhLMSL
a6VtKRZXFyz0dSo2AuskR71uoLLspzU88lHnaARGCfQIdTGAIv62Zkl1pDdGb5n6fVRqFc+b78/r
L2THUZAzA9T2HZ+r1kTN2eEjN9TmFBlgUHXWuiZRvLOlgmezi+nEt8d4/OmuG7AoTjst36yIL63e
bST0csvfIIzu1Vvu0au9DBXo9JdSEA1BUzbuELGxOLx1AfHmC1oGPYYHQeyP7VIK6gimfst/W4rN
sUqyqqPKwWT+QPocHuWynz6eMI4AXbhfoieAYc//ZkG9lVFjJRUrFyAX5JKUg9+lrRQJ5l047Zrg
cbqFR0w9HYFVvG5VeVrTkSw8vdChD0UQbVOAuOqwtr7LYDL+eoR8gWng4395klfFmmeePZ/99P+L
evsnhM6KlnSCgPr1Jl9yrFdYQG8ItsW4Pgl5YD7huVTc7b/Yep5PXHKKSNwVYu4l29HlavhdnXAg
QVK7EJHtaxaIwC84Sfm8b+q+NsT2zwCKdyV2aw69uTWbehDojV4o2/4kGETkC2xWmBjiAEuGCywK
wQLyzm4tJtTznVJaD9x4SZRFSXPZLXD7UhFdnJjGxaP6BpibcK1vrpKSaRe3yx6AU5rX9bkSYHxT
FdKPJpi1ILB8SF+MxB4Xx2I1AZDdkSNVMn/sSjc8X1I4d6aka7RHO/GhIDZG8F6h2uhdOjsY2dVg
i4+nubxz4RB38kd3q1Rrq0lybcmiBTJ+1tp1u6Wk4EHfdGxzhNkvtBnAxB0HlJ2hVOrlZYbKGHkr
fYgxtQ7knJdz6ZieNqhvosp7MikSJNmkTWiuItWVruWS3qt31gNQfzzvwOaCzaHJFudWdvEECmXG
ijwefMkbr/ZqHTLF5QYDRC8c9SdjC5CPysSV1HzrDCpFf1hkluCKYHvhOFxG4M/DrSJrdzshYpZX
JZFXr00Bg5eDgssXMzIe4+XbIed2BQQ7aTgOYTo5LRYUUZsLpyRLyKY6TLLgqAF8OLTgK4wHLUXd
nV9qcGfykkpdL3hyz3JanBK5CJsm7XeZJETarfRfT+Q/x9SeY7dRChmO4EeMEvnbVjydXQ8al6JF
jdOJpM/miYTDVGX3jm7Z+TNfzNZNpb+zUys0mLrf5+YgDRG+sqWbCA9JP5kIH/PpYdv0D2ohocG5
/LS36EfSlUDw+QmVBoC6XsuE0RmV4BGBzDGWQ7QepHg8hmKLodD2PQS7OYQrJqvOBhzJUttRVDzx
+D7/UPl+6mFbSFNxeoDbOfR4pG4CaD8v3h6HFYdvEkAw+SfyW9EGYnHMGF4jXZXeFtKAenSRZl5W
9vZ2LJxVlsgQZC6YowzHsty+jmSxN0jxy4jD4d3IwklSWlKzbykpGTmZKKd9+LkGOZdPjIF4Q9Wv
K2gCXt1W7oyOEjkHFuhxgWiRZg0RRT3HNYQQDmCDRj7EFhzqVwDhSkduL7ltwE0SJh3p5LRR/Y7I
gezUk6aSKDcz87BFekkBwzyxVj/wtvlzsbjgdCvd5dFp41qzs7kiIS6fIJPloaiZDsFG+96lp0FY
murUajdBTv1gu68mIMgzEKToK6zbka8qE9v6T4g5fvAIc8xGeR73mZmLexjTrbyOE5aS42Sh39ca
h4ImoLg4MGQi8kr9jbBgoeRuDyOKszOWmdzne/oSQYCbi8Gx4otE/hDLnoh1keCZ1RndCY36drFi
QTttX8569ypADGIA7QUL6HWbhYi7psER7QJOvDb0zr2rwlYU3/Fn//sY1Mj1XMzgaHzUrYiRrsjK
x1lthZHhAvbmD2J66ER3s9zXWYWE96ij4GLY2ARtmIhzsrm/0eRMCg3yrCLDzo/Cs6BKdcHYMCZk
dxG3J5U0Cw82awLxNggOTkm2tQMX3R28u7chvVFkxqDTY6VScXUFbCtwu7l5s/oiehoP7ZE39sax
i7jCIBPM5pxrfiXgSjzM7gvu57jfF7WuMOu3R1pSJU0dy42p3NB+CsmHZpMIoX6tzztdDnBaodaC
jqS8BnuVGRpfPytPW7ERkUlkSytv+iaz9tjETitTpZ9X7jbakwZ8YrA7H9NayoymMpH+ocdCtcUa
U3pz8H4h+yrnTilEvtjt+6zHFapmHxJ+cGFaKC29bCthQuExVR+ENdMxaYiEsn8tLcDB24/7Co6+
6niDoJbF4Nj6l50cr3XUliULaDJczvYmiCbb0EKfCdj1yzB5Z+8d1+GvYA6zSdoWjpHkNVXUF05D
5TTgTWZ6qfCvWfFjuhpovM26rnp/BR/w5yYK2k57HsK3QU+38ammphDNJ2SYr8S2LwuLjU3nw003
/FZE6VwDZv9N4OKFJIPH4ct0MTsGnqqwPwgY9ACCLZtrbDKrsaQaUK2jb/27Pg7izBD6J868z9Ws
VP3FpVdokrpBF+iwHgueevzH4bEtsTag7Nfva426+LtI4BDkOSxtflEYcaVDNB79tRJO1aoKxPX3
zaw/T0J6lOnQUFFeqPh/L6PJVntTscJ+89vy6AJyNuOncEvULU5A5Qq0YYrB5os4x/pA/fxn++Ox
7N91nTnyFIb0SD/0DU45MrQNxA0CTr1F77DIilQ6q6+a2aLEEKxxoSANo7l4i8vgx7c9NKadMiic
KSQQrjKN07kC9UzWRgYldEdHHVa93zEVPLkzIdWXEgxQRPmEX/uz6j9L5rgRD076z1sfnnQQD/Ad
99Q8KLfo1+BHbeWpiYpxnwevWfSUXBhNyVzsBffJ63VwkF2Xv4I3z5OJ0InyRiHCrjD8FYPQOeoB
5tl4PQNUQ8dAs8HOGBAs8zImjdXL/AR7o+PdOoUp0vI3PDlm0dpSl4uHzxoAPDw74RJa79DIsGc7
PlXsXyvzDSkWjsxUvjQsy6TYITG9Ld88vplrdY3nC6uA8G83x8XuHJk0vrfVUuJeEfDAyvHmF1FC
bGjOTxecFtLvI1drhsTmbm7jOqHrmXu6gK9YQKYb9D6/1eP7A4UXWmg4MPTih2uOY31OwwHrXOqD
xv4JGZ+yixHLexoAJnmXQXp6tOp5yoeieNH43L55v+DJSTaF4pC93lNE3mymOpErYnZat1/Q+5hh
jPhOBhIwlbYRb7+oDrhTTKGQyl6o5Scj4phklpudN5N+2VTdCgxp5f9K51D/Z6Q+WiAvO7Hj4cdk
dJMaU4rbRy0vdFYR4knlN28ABg3yzEE1GnIS0UTgCkZ/r0Aj2h1mpB9JUJHwoGIwq4/RsxaxPKDt
cXrMGjmgn6ioo+b0Fyp781wHl73XMp6CzlPv/hj8MxgPrUhyfjO5k9BQ80KmIVZMxaTyTLW63f1S
T455T1olP5BAwPuARnvrmcO1lDze9cuVyvtcF1z8I8EACpj13HvS7znq5itip+UXFCPbOXKW703O
JCpYIL3n5/5a+tq+9qQPNiamfMgkhl/KDKBonLFfTd0IYHNTwLVnM+Y4+XNH7iE62oXHHpcLRarx
HguGJ2X4omPcukGW4X/D+Rh9d1vxMqVG0e8w6Y1fJVv6UXW5t9ADGrTo66LNAABCNhopJmIU19zn
baUV+qpptiIFY4fisgT1QbT645p3nicKdmv+GIN6xG82wW+MYqMh0MUCS3dNvshHyXb9FqjtpRy+
wR6q46YI7UTdNvYpCYHUE+hKTxbysvkUByndUaL/fwYm0cRSd5wjHMhhDim0ac/9QzfTWpYN+r7X
zLIO9/Yxhl/GDIaNj4pJA0g8I2CnJpmhjmKEKpuCilQ2M5lLi6Bs5mZYEeXxPXeVePUA0czqt5BM
WxsHHaHF8EziJz+HxpLqYV7wfZV2WrPTAPdLdrqUTYlTVf2DIcYe7hzjdz5L4bCzFPq/JSY/L/Pa
ogDeTcEzkK1M8t4cfLXtcks/vVbALCxHJkfzizzzUoHVavysLThPrzdf6eVtfKlPoq3ixDTzmhjN
YWGcatO7xxgiAaNwk9Hi71Xr4F5C0deceQV8phsNQQ+M3SIsx7l7KH1FcdtQB9PT9IwZVBnb660h
hq4eQ0hyb4kR+Ls3CBiPXJsW4LQIHLkk3dyVJvHBKGStz+PW0WKCZCZyJYwPT9IKyO9Z2ft6A3rT
wSu9XxRLlRUzy5LDEwMDJOtr2xMh7s1XbqXnU5bRFI7NqfyP9K+8BnkUT4QViPDOnZDXX4DFMjC/
BhCVaWSMfBdesEpff6tBH/jtyfqt3Xl13jcQEXaIuDruHk/0kR8//twVrA7uda93ZPooaJ1orP2e
MwJ5IlxRUWQ35DoUlsjFXS1XxIjxKFzaQcwUuPTLDTFmfAbk1mrRae4ye0qsSzup0/3k/fCVf8nP
tb05EfonZ8/lpNQvQVBCcNeG8lS2jl9OdEaAKEtnExFHQ3N18lRdAASpRgzOPyGWVI1mqd4PbyYh
BPO1G7o+OUZOvZy6Bv4hnRrNjnEFgdfdiqmifzU5NhKHQ43YyABKRy7YkPoJwUGmT47pycELQkrB
JUdWYn8tGgVRDxFbI9GiEuKxjn8u09Cd9cLLRznZvhJpe9QRT9rTgZB8C6AGry880K4CRpJ2eH54
qyLjVE99o8BEA6AmyLRalGkzmh+qbmHfTEXRuSqvPLTzs8WcznBKFQpdMPCRmltLqR606aNNhrb3
8LWfKLChxGrTP4/jM6gX6doIaNzUH7FO5WWtstasN4efJqUsNPNWb/VN++ruuSOwDzmHbzqE5zul
UwVgyeOSbfhsA+JssdUywZ+w6pAqpTE8P5TaZL6JjC5fCPaG9GaOj9g+rX5+w7XvI1xk6VoKh81+
NWDeDOWYwVZkd7UX4dm8OVSy8D9RHLzAuzhhYFOBZdCUIPhjR37j9Y8L9jm7tfhLwvtG6mjK+GMY
F8w3Ok5vMFmf+7PGnom4uE7++zsojba5okhgsayseXEnJU9z4Bc1xyXweIhHMr4ytEgkdioKXkBF
a1qxZ8rA2RmndDow4zeRUk0go5eySxpKV54GE40XLVue6gEm9qhS/YN7u06sciV8gGdDp5Dq1pG4
4W3zF/dY6FwqBbc5Zdnf5oohls4rBUulzo3EahxmcQEf7SEEi08P6besO+UjGmp1eWlXdHBvz01Y
ayj9iig2IKBgU+7B11QlZPIdKikJM8XgxVwln4V8Q50tQXdeimh2iSY0BbmGCtCRU9UImkVowpUc
iVTLwlhnm1dlSgqqyKOyJGlYTPj7q/Xjqt/U53Td/8Fr0ttbChX1r8Dp+SeToeDQXYW6UKTZgWhO
sxVVCaFCDkKZ1N72ZBh1+4QiKMPcjqsm8E5N3Y4MUkqimKOwHMneg87hjRS8kF3CiJ5a+Vf1LPrd
EHa+V5Q8MPrpsyUCtYJyBsTpv1RkBNP6EtMRiWSSJMlASDcQ2VN1Yq1jwXShhv4jRdwZrxB4VJMh
RLrYf0rNbgSMBZTkCYuumLFVU9pyRb202gR3mvrTYMQQjlBO9wIPLw73gpLeCY8ZLysnn/3lPcHH
iaIkTFFR43eXp0Dd6uHS+BpVDB7TCrBqWta1oFSfZDLSS3jh7R1d6u8KByoFi6sZfS+qL1kjjxL6
PArDtX9bFdP4DezyPrWpu+AQdYSJ06YfdAJ/CjCSj0FUyMoQnlZEV8akgwkfip3jV9WGJi9SyqqC
0OOrMfl1V/FxHX6hvlnB6ag1CNDJsl/vYQQ2k8m1XR5VMv1feqviHzMxvvCzTrsapysQ0kaf9pxb
+dvBz1S2fIb36vv6jDVGXYnyn9upVsHL9mQVVB++DvUSZWJHdydER+xSURAy7lrucC2BRJABhrLC
LOngF53ykYciVvi1LapjKJjZGNIM83cyoyoa5BoInKgPcVu1idD9pp+J8wmpR4Vh0VgW11QsvGG6
+gOka+c1wk1RcbvwgMchZsun9AHXKd8k+puuOuBdxIfsA1YWA7WU+iKuWWD2zILIn1tx+hwUPI3U
bYpRE1K7kJ+p6gjA0QKDRqKyv97RkmT6tGLuCI9/P7Mbf0ZsaB966m/bD9AgTTI/Lxf+dTqvb73N
DJHxbwvZm4tZFh8rQoUdjySKbWA1UNZOhb7y/Nv4FBnbCpdm4FIuKtqPLN/ZFoHypeD112j3cp10
ps1YN81ZN0XI7fIwk9EYUJaAlz3s4muU1JiQEcU0w4mZ2krR/CyWCG+TSvkVBgUr2XOoihDei7K2
wqnKV09qAzFKUPMX+SOf0jsv/0DqhwicpasOl+vkTFtAZdeaS3+xOiUGt7U8droyZWXRGwd+jfw5
geacflNeUw7GoUOAB/HV/zbJxGVgo/P2+H2TJR0YFYSNxiwyPtkBN4W346QLeOcMOevTqSZB8Pv/
6oFMMkEQssrtkWGqkC1UP5VVhUOGhfGivbNIomN//Bh2zpEY6QbptwRdlgpAAs2oZFhOz2SOxwVq
QExAf57Xwfmv2WOLtiG5ZMgY5hAWs43j6CPp7OpjRwYxgZlIxEETBALPzQ8+4g9Rtq67LqHP1Vji
wQprSmL2qCOpR0U1mhmf3iYAKudn3wq/JYdSQCtUGgGlylwtcldSIokJ/+Oy4G59qEs8lTYWCH6q
9asBToK3aeW2y6DNTqf2Qz4InpvvOYfnGv5TDB4VrAVy96OWGVB4F27u+1VxnugJ1P0deVdfVMel
ukR4Od3BmV6lAhvvhwqjS6F0GoRUBy7voz2zVNaGT8wpg5GLDMWXo9h5+Nap2RMG3gSsYKfTIf7l
WhFAjPN20PwOIy6r05wopcbGnJW1MYLjeGCsF6QKdv06kGgji19qwI9ebsWhg32HJbpIoKZXz6co
CIakeMxXIRzSwvaD6l1GSXKtJd2+zvNRE36OU+YQA42BwKFYegT3UGqEfHKNPOoer/IhdPstNWeK
YD8XQExZcs3S/YVOEtMPeShWsoUZuoGAz6+8OkJqtwbmhKLjs0S2uNx5AVmLPfbq1ODMXEuSWkyr
qo//TnebCZ5TGOfL6PH7tfhmHnO+Z5Ca9CADXNNfLKnsvrq7lP8LJa6uICi4V8JiLRXkihPKcrUM
mL/GNGE8hwwgtxfvxODcyP2wzyk0IMZ2hTvN2Rk9kWhBEmOQlBbPMcL5T6+/TDW/8TA9asi8s3Y8
A1L1bLzQvHgoPMPoIkJ5FugaF1PnV5hox1VlYE2Rn/zpH+hov01Drli52gYYDARv6saZMAyj7qz8
CQvN5mkqlSMVsYZVNCE067g2tA0z9uAD8RcohLBzKILgYojXEUFL8RqdEkGMXSGhac4h8pDF7Z4N
pRhvqMKzH0ps/6RZ4nar0PiFjP57dR+hnRAkO5Q/sMojLDa57TEZtrrBfXWTWil+Gd8vILuv29GJ
1duU5gjBPF1Vq1lTWkGKdQFDWhSA0YBMKJ0RYrQ1EDO2IIYwS9u25oG85dPrmTkhFQ7d2n9XaIum
KKICk7wpg8L+XBWs8dQpVfHDWbrdyjJwGQQ9lNTAYxdq2GVNJBWA9r7pXFn5j/rPwfGmP27YamD1
0v2bdVeFU4GLRvtoYmZSORLJKpZ4GNjU8IWR6uA9H1zOJ2zHuuNJJT78NsetE4LJwHBnzDIODWyi
wqoiFpzjRv0EcGQkPai7J6BHMOspN+6KqfBYBCrsHLalItN83I+GWLxkVzFPecibJv4eFuLMtBqE
bV8rjDZ6mfnf0kRAZnCIhI7KjW5vPjz7Hym/mCFnzk4x7pAt7lpuehqVaL6PAyLmAObp9JQ3eOWb
e8CUTPbKIgNPR6HPZBnmF2KpGKUdb3VD7wkFSDCHyKXReEe1fFb9fsShjbaiQpmrkzpWCEbm53ak
dhGllUtrbvfnbps07w+BtcuNc9uwq4Ldr6qEpFA+9qXJHFHUU5rb3KeWyc3/m8JKiUyW9zgnz8Hw
/w5O2Qch5P9oIgeUQLwkzTXdZHG0xfIL+Il/zVXVPDOn4v7uyAz+dWanz92KtBOYed5lGDSNNHoF
infhFlPBvLImt+JqCqaf5Qn9/CTXjYwnMRtIQL5wwv45EVncWIw+vnYl2VPkd7J7HqnUnEgeWpN6
bOydqHzMnf3Q7gsvkQ1DjRLmyacTstaeWxlBPJN1jJukp1Nca1RuEhqSB79dm5VbK3/UQQnVLJFQ
k3mn3k/n5Kebo6jWkDHxrXq4Tm+hBunCAXL3j2Q9sdEOoxooAL4P0LRXTcKjRPgZZS6Lix8pWXMx
vk0/agVNGL3SM/IiHolMeo+BAJLQWojfUsGiLuHfZIn9bz3QbMEWb8VBpyuDmaKh28YyD0fRqGxH
A0oFH5Q9Ka2cuwXxS6FDmp0kX1xwTYsWp7NxCWjeGfAFju395PHbBX+i1ise6OyCeTpaKC5NPuz6
W65T6R2bIbBX7gkPQs+Mc0jLxGTLrWp2bg1XwFuP2O7RfM2MNEjSs4Mx7BmcJTgxCzuycG90LCXW
aVAcEIhvUmWHs9htEuEIXDE8qQthM5CIXdX6t7sS5iOBbuiNVIIHWd6rV5xicoy2KzgfI9n1M/si
0tvyo8QkVc/+jfY2xwD7oAR7GJsCUtFPlmunyNw4dmFDWugevrbzNDVi8r0CVKWPVLA6dBaDoeSc
YMewsgGzRp9MfRcGwqXcsu4ikob29HQLCPStVt+EWZCYOg5dk5GBL5MqvYRYtbW653BXxxaXT4Hk
Po1YMseCx2pBRYwjk8nHgf/jnXTE2rCz0ucCI+O+KkgHBfnrqasvCUgP6LoPAk/OYMRKE3byFtOa
Pl82OOTzqASiMaJDDlM/x5wW7MKqJC7cXz3F33dlo3zktQnR2YzrOy62q+9ycY6SY6wwrMO7DU7A
we2g4HDU1YDqckVqOs8V0dmp/dJTqMp94WSFQfCIV69Q9PSdwTr8ftNB+uWxQkmQ+7BJZB6cb997
TcoPQ2MjS5JMjKJHbvhl6GfSwtwFGgUwkFbxKfVHMObTg0iZ97wi3s+qB+x2NSV0xz83uyWPzaBz
cOkrnld1O1X8WuUFjmN7jVPNsZ1i85ep1TzwsFCKKEIQVOTsv2jEK4dkMqJevj0Pff7dQ4vlI1dl
8MA7ojdRGiX08hvw482WcECYX9GUFOw1xmc2neDw87SSfDR2yTD6TMfkJCXdMRHlcejhuDud11wX
QEOh/RRpoQ9idpxvCx9SSw57CpVbp8g2fWQ/ONPphREnZ1p1zgQqWiDFswB+hi0++tbcj9xS24cE
0ldE2/QgMHb8+1BzCIVTJWASxcs7zB2AMOD1DLa3duQ76shivIk3Pz0ZmVocUmdeRRGsxdCW2wkD
mpMvYkuY7iVgUBIRkoGZfmohElHBqccGipb2UmgfcuGuPRT83cHf5jDnxOZqNUURQR3yw6pG2BKX
K1Ij2A8zzULTasKZfoeOyI0bMO8O7NTIkIuPl1qrIxc1R5D7VX3CLbeoRYp8P0TG9MTWNSYEsBq+
BH2UtLt1ZboCbr4A8UCZMFMb3zsmdr9jS2zXfbJZNuT/GhvxbfBq40Adj0GNk/MwZmJEHoNDZa0y
BfGtZZxV/ynf+C+P7ajRrbmGzSpEM3LwYHxmEGziBuTVnYwbDTE0EUCwD8LmkgiUSdFttCCol+f3
1DuF1wh+7U4IOL+Ly/lyVsFkxoy4JyY5NPp97wB0ilSXikv1lrkTBahRqm/aW9YLgpxsG0KWrcZ6
ZSwirpJYWhff+qUIpqWixTI6MsyBeQL0dP2wZd+2YY9P9+0dXgpTF0VAY+h3VOIynwc1FXdqyYtz
jjL61uEYrJbTeFo28TALNoRUpbdT98reorvZ8Ilyw5ILENuwmRKHXfydJAq3okMaDzRshmGHSJ4F
qM8z7Q/+M5jEzMWaAGvIS4q9nAqrkXx9VeYLGAVvzy2d4Yofwz4o56DREkkCP9O4SzrX6aAU5upR
OAxjXUZtoX092wyf61crSggBt2KZDr3bJ9jeE6IUlPG8g/FMUV8khxPvGtprG/Xs61fqwmpgwmvf
cjpKrYf0RyZIjkBhs6CzsieOg3ukqVDzQKECAUn3Pkx8Shc3ws1bSGLWBjIL6PqYkF0dkQ3i3zCL
HjHLgHkKqEplcSoBNL1DZ+uhGSOKJCwzyszgdHWn4UjB7KKx6LCxmJFVHi1tsgOS6hcA+xKQ90c7
VpDMs8kX9KVhMsSsyk6L64Y8GOneoiv1DTUhgeUmyrDwvgJoev+ueLPylizUssd5i8Ci0T7yrwxn
mhNwkx1KDrGyUpa+04rxxz1PddEorfMqW9PzMsQZ6sGhDCvlEdPisb+LgYKu7RVkHVy6DP22Dj5P
RUYgQ/eMbLBiTjNWuXRpTEim9O1q/24eiwMj3b4cd0daZio6Wh82DAOJUv0AB7MNU0aJsvAppJPA
dJdKwkldva9iKVvFBk4LDo4xi6eSbmtszcNDZZTfIym0EuM2AFimUCjkpO/u5ehz4AQ/TLRGIIyv
wWkBpOLydbAKZZuzOv7i0iMXOn+iNPzF+kk6ZRlCkvAAR7WV6fAyRMu/qNNxcsfYi/phAoac3gLH
3/3up1YMZSXMXcJBsL9gEwetyyjXxfkak+whRRy6vN1B8gb+98ba64BKPYF7qOp+MysTNTyXHOlm
aHszkJhxp18vQp1cPrq3p0iNShX0dCcaRxwZUbvYH3jwfWagwM51+cq0NgqUwB/X0zhubB4b+q51
Y0cI0LlojlvGXD2i3JXbVlTFUuhMhb4cRY5gKRmHfjou3c4lIN2sld3CxrMefO3N1JpwaWzaTXqB
jcsdvAyWsHQ391w7F7yPaTr5Zt15UAnsRzEJgqj7HrDttqo4ut51wPK6YQARZVwdBk6HApOFojot
tgxa+fkLl4Gh18DMin2RHQ7sJ2Fe58yNGRZGGhcmJisJbBGF65NjM2qRVX++UMgcuHCx5V+ZDbm8
paHWb288vXU2/WlgLEpb5EbrgDCER7X8Rdwf4/bYr+wTf+xdPWX392Zy1jurki72eT60JQtx1g1f
rHO6BEagbl8oH9PlSe/UYmE1v7c0SuHe5v9qrkBoc/w1Kx8nr1SBSiraq37HfD0MAmRmzOfG2S+J
h2JhQ7bm66JTqc3yc1RJip5EAX6We6r1KLVzesSI91iisN2rqZsjFCg1p/n1GwCWKu2W3glkBEuZ
zJwYYYUJRT4EKjFwbmvtFJhC004IhGbLz49opKYj3rWr1vYKWHmkq4eC3jGniF4pWHAjoNAsJcbO
eGNmUPi77SEaGkA/0zzjPa483Rl28yZL16w+fXlur3RIycC1Vj+olOf/xpWtnf/aQbAOwounX2rP
0V8+T+zvlulNdXf/DJlsX0acNL+eBNujzQZLopEPFp9eu09qfSyGsuzUGiUjocA3ibd5nUren6u0
NnFD3HtVv/5MV7tZw9iqCBxqJycc2fHohibhppkaFiLoSfTjRASgBL2k9UMS/xqdIjJVOjTCdfSS
+E58wTviLmckpyFmlhphtIeiYxdGtqMg3ldqUeulhpTgAiQ479N3LEpRQIriX73PE9Fe5b6aCjf5
LxkkjeRThWo/3c7kTiI49x6U2zQjGXvQYaZgn83cQZriSMSzjnuZTWZQWd+/W8/mbNJvVlYWFKxB
8waW3VacAzlUiIVa2dCewRuAJus0IWGNCIGRu+35rAQu3jATcd8NDkE4nOGwPHfzj+7WErcXM3D7
YwBky1P50Q0v7Zgq+gzWXtkFnDtmeqTwPnwD28m/68vNYTs5OaeNDrikeOgL5rVpVU/9saP8YlrW
su9dtkYSHHllZIQGAGIve+WWg6ol3o+abiUlXKt+8CeeqLPUxP6s4nk0MbbQXs2aKOU/mkRmmwZU
3u1iVejNXCLqF0Z5qP/Sl+vsyIXiC6TMDQ19CPpcVpV+MclQB/zOirqf3w5GCct/NxNQAcM3pj0F
YfZpjd6x7QnR7JGmMik5AxNrhY1VsK8g5hu/fkg7QggNLsxYI+ly83EoUFYjDAZRPU7aYX7nnloO
Re2Wsd17sThCpit9pld9lQi5m82KlMNUAFCmKOXsaT0ZDg0ezUFt99lSvXzi9+Pqnzs5ORFq7gvH
FrJJKuBZMWzMK/3XrUAQm4EsW9t/kVdk7XuIl+VVfcXA0R8Ro35mdEbjInZNkbCqB5SWgHyrRxGn
ZB71fRkTAxisdYtdPSnE0PsVPZ5TQpsx4nCNV9ymtJF31x1CRlNhyqq8y5ezDm4fx6S9YG1iN+yB
x/GZiXQQzeH2E7rXiEecqQJNx6DT4iJ3SsJtFutuaK+Au8ZH5M9DW0aWi0wCFvRusFsyEUiMIii/
Dxne3Tnp/hEuAUqHqLHH3Xkki2mAmwczTVU9O9PAmtzH7CaGeBErpLGCZ+Gmb7NWWdlDGSO8gBiA
vRb1yGZuK6zsXWX9my2w64qOS00Uez0uMi6F4JpxlC9taiVqJREKD3Mryz+N9NSEVqdqVwNxJyig
Dr3TbfOC46ZQFWUTrT6zlgLswLZ6MDCyorp/hxqyJOurNNb8NkTnRML2LAiakEEQlgIHGXHwduMY
CmtZw1sOFv9STa5EFZ4Yc6aGb9GEBrvh/ZRP2VBQxuEOkITI4SLALl168JXbLBzWa3zZELvqLqvx
lH2eFAY5bnUhr7RRfQBEOVbcFdXK8XXRW8/uB4E4ijuOq6qwXZE4OXwGr4OioLB2Nn+u3dB2Uns+
BHKyQslEOpf/xpiQR94P+oKoJsJuElfZa1pug7ENPjjsFQVJsrHrF5RdTT3rKB5MrEh5Rad3Ax+g
jOhIEZr7LEjKV9zlveFFDoquRZrZlBrGQGz0fsG1vxo1GRdePuqaLkaGM7XDCrZc8Fc8yNv7Ik8v
mkBbkNT7kSdhYcTYGd55j9o2D5VWc5qela6smPsEjwApyrmPolGXVTDK4x17qylyLcLmqslnIrb5
JObccVc/Xvm6birv5MltFvOa+nQwDkDFudrcObW1qVAUHXQ2VAgNPQoPFEOIYYqxYBqDW0e1egeP
sHIZ5arnAU/4A3B0b6krMuQmWG6qTsU+urD0J3MP/af53PM/HwBjt0JnNygGHlThhl7b/Q0V1Wt/
TAzNlPJYbmeTPgkepyNdxT4lPv3hR/aIkk0jLH+imccFuWt5Q0XvH0oIYEav7H6dEI3EMA8YjqCK
GwnFDtaKUPucUGB7ZqDeVWdV2UaVhG7kB4pBwQNMHumICeBPovKUCCSfD2H6Z04aM1shR2WfxmB/
sUxa/1tf4OsmFQNTcBpPuA1J7/pbWHH2PnY828K2vUnZq73COgRvW7H+MHJN14aVYtuv/OIJJTz1
djbn04v5+ulLmfyDK4N5ot48meADnCWeB7cc6oLS3S6FzcIlwUNT78gU56ZOGoIBBnYNX6BugwAK
O61R/TPz1jyhhd1/0wbCeFT+e0Pj7hmbEkfA6f5Cm+iXCJlTUonrTj0lZTKPsDb/jIVVJIMvaiH8
82+/KTIZJLH7z9TVeiRTIH0+0yNsfngSc68s3vvzdrlAsCe+FOm421PupHQB1TxuxH9kf3+JiI1L
XlJk7ZUj3d1I7kmCX+1CczOIp9FWza9yOwrdacCmvBrFoQwZrZ56wNIaP9+Gf5MpqfRG2kFhIyic
1PLNtMDwfWWdCdE1+p1fK52ORiJZIlOvzW151t3JksxpB9mwKR02ItinG+i5EJz5a1vqJW3kwczR
PLOsCQMCeUmJM81UBYwX+DuS5FQXyjoIwSAxAhDjoF5YY7mUAzEmCNZZjIYn0dKh5lagf2jkWdhh
OorHD4iBKWwLSKmd1APLVVynEP73hYS2nnWYdjeo0Uz3DmeAVowIOepjHFatJNDvk3x1kUbEgmXv
JwTlKMv0Vsk30vdpk2y74YB2292Y7vG3v8I/6O+JINgHic6zfYK3WsGl8ZUmPVsltuGJV+W1JtGI
6WQoOtzvTfFRhXs94R+r3I2wpn5HOR64SJuMvlBb9vRcVLfcrzp2q+rEiy9w3dq8ccWs93SuwE3U
XCgIfxawXXl1563LH3F05PX5bkJc/mAszwi/O7a/GAMzBFW7CmGrI6NgAqXNYeSkPWNEK5Rp/SQo
Gt7ptt2gGYiSG7NFxUNcGwJQCSBnvHeYCgY9kQ3KkfAKQuUiYhQHJaE1Kjw94dc8BTyeMOai12A6
JkFyPpam068fsPTW1c9XiYRKP9uNbf5BiRMZZHl5KchTmh1ytrL7wB88popVywKlTGZd1vjDKQx1
Sa9EMIY2U+EWb77Mu4DaBjibxY9xqZX9SwGdvUk2kFoX1BTkYN69PhLzRjVvFGB9xyiXydycL0rK
OrXAEsEWuF172RSTHW2hM/wFTF6XJb3WWLggSmRwTlYnIomM5J36KF/LZtYzjvEfFzP534hgOVQT
QJ1xGeRuLXFQ9H0+Xjg0NYdudkVsUtHvQg7HOF1GzhHP4Ho1FiMhMN6zRbAJ24DZtyHT5GWmz7Lc
SJwT1lpZ6NlXJBt2w2HqtaRnkTZO7lV9jKnRTki2lJPFRgRMnnZEpwhpWcd/mj1gmLqbckk5Ej7y
A7ayi94ez8Um/s0zgHZG2ZfJ3wTqBoxN/u7bzwhT+37sN7Hm4tuEPD97whVs+vXoyYaZ/jNBrMgq
WB7aTwg3cIYTnxhzmouf8/NO++F2b5UMi7N3z27BJcUeiNvCCfbOMIviCGgOUB4WJXytNkwU0gQ6
JGzumxSbQrdaDvUskuH4jrxEB7ClzydsQ+PrP+XOHONT/a9xuHV5EWOyriaJs8qsePGLZ92F8q8V
cRFC7abJEchng8cILnDOw5/oRDLr0Xk5L/juPlnwMwb5w9p1NYgnshW9ijv4r9rFsez/05o2L9En
4ogdWPx19hc89PzUvPyXA4riBjRcPbpTWOLQOeAX+3XAVN6snLp+SONIYdzjQa1Q2hSj+3Ex0/0Y
1TnPuF89cVSsxwwalbNS+vw5rRU4tGMqLaKtXhNDtHNRsB9dK0CnhxL3cWLHaIFQRKbTDe/rbSu4
27ckt778sJ+i6SFGJd8SWxQafYCqbsQSEPqyuhi0kqPq126nsg1BnobDGPtSgIsOY6JpNlFHS+9G
OkESn0AK/ZxbY3eHaVDY9L22r+9WiBecIZ7+vGpCCKEWVHifS0ck7myvyPeBd3+gHvpVQNSptXfA
RnpMJdTWk1AY77HB2v4ESvv5ffjeMXqOl7J1E0aqVjJb8yC0xPNN1lDLGnR3d5y2yLXYyJPXgNUn
6EaGwjGqqeHj4Vzs9orfLe7Zua9KV2xx89iP9wCzjM1MYLNeVlhNs8nyV2CugC/oFgW8PXHlUj7j
fDFQ+dDKavZwn+dz2+WUeKIavk4PfPsvS0pg4Pt/7aUGsGih9N+Z7LmIpYHrteyxTYuQlCKXHU5a
0lfx0v0igXEdiCd1XPqdmIlMsUENlltr/fneOmC3VN9fcSjG8OmW2aZu2GRyUHMvqXYMKS4k+LO/
9hTWtx182beMAxNOVnR95DXr0NDCCG2U7+76Zp28fl4vHCbQVI70Zct+Jo/uCcqYelB6QgiKG+lv
FXeYwSSdi9XXqjo4xnh39Dt0wuHnUEgw3Yc/N5MJcIDuNi0E3fqSpQ/2D0GOH7sYeWI1BooWbpTs
9jl98UXgQFJENbyliDAqxvfq1fBKfSkYZu0ORYJlKZLHqKOb1SOLbStEvMC5EDtCI7D+1MOM8HQF
9M0HG9983ojOw33j0jxyloYYk9+Ls6QrePLyfAE3JJGBBH3r1jQviukWzlny+guNNE2o/nTx5tqR
m08Xg5Bzx9L91Jsg3pVo95deZQPVe52Co3tjUFQeHsN7sNHQljOa6bKYtsVKTXbtae/SrziMLK9S
sFKLSnITxu6zE04dPcQf9GGjhtCQWeof3o26mXailXRAGfaR6bEmRtbwyQE8rXftv3P/et9Edeuz
QJBANiYg1QtCKFiLAXwnSsNrqEXOwYSdGOP0EsnPZZ7rrYK1DxJ9AnEVEKqN4BTyfKJnFBmc3gC+
IbuQu4snOhbJGFJVNxQawJUOgu0BJEQarY9p02TjhA5H6AHqhq6hovrzVFL7p69WwW3x0pWjESN0
xGwboNDrVy4C4VQl+AuhyyfyJhfWo6rOXX17fVpkNfwqTj8/SiWB62YFErIrREEs/ClGno1tdSrj
7AFJts86DgzmMPtP3PZMOTKBelU77sjpyJggX9MGmNzA+SsTLEo5xAIHoQ4abFL/vAF1DN5sup46
3rdSS29DMNRAlhT4SsTMaMV4POl4TDFOqJYm0CPR+mxgsiyXdvy361Dy8ITGlUzvLbyO5zXfwT8/
RJei2POsyoM2I8HAtuYU3ZbqULcp7Fx00Gl4A2ZzVM0HoGK5miteFi1SIPLv2EuZh6aAUqGeR+Li
mbw0YBP2ZIVhSTng+c0p9O4P0PG+ybxXDW67eB0+PMzNgUc+WfrOEvsXFgXA9pcSrC8w8HtIQesY
tfDYPjGUGTFfzLm/9ESRa8XakH+lxd4+gAGFRjxYuPSkKaW9RHa5bIjQTSmTxUr2C0eFlqSZxHK5
r9tsHBcHxwwx97GravaqqIzLmkJ/HIW5Kwfaeau8zg0nd4cUq1YJD/XVVHfMmQrFSss/KhvexuSB
84aGIftihaZ6kSc6rJFeUoO9ECiumP1tSqOvUrD6YVsYTCxl7eb8yZmiwENpAVUNIN4fYyxOTn97
wcBhDsKQ5sP3BiM/f/tQ74iu9KleHEyi/z/40sG5UrTo/Bl9Nk/Hz+Ysl2uzR9V/D2/OfMr2cMWb
8ktyQmm13RLtq/xoRRkY+lAxfyOZwWlgBLc60DtmLEQe3etMTpGBMiZOKuEPAxCGL28yibcCtacF
XRRGXHbDTMr/QHzp7e5oiQe+z+l7GoOJubhzb3iolM5I6jByY/jEbMCOhZ6yEpsRr0DhCHMJqriD
UGDskSoDFVrfVrCBHcOtaBUDMma2F+wUDnmwZW/x7qFg1z+whmA+oJ4MQW0k+3tJrrILf0mxCKG2
rBr3Gjz8eoM4U+El3sb4BPyoAa+IKNve7pX8iTvP03wBtf9gJWIBEDF+cNFUVUBddJ9f2AJS45/9
kRFIyJEtqO2B0sFXphr8B2LqwsDCxzkdi1Oht225KKrArCrlP52RD4TCI6l+Bkp9YEwrE+NPvwR4
U3TkL18JEogNpwDc1xWgGh64vBA2AQlKUTIOyecVnGrhZtfKlLR40KlhkC09FVrJfTqoRf1AVNBD
qJA3fLKe3T/EUPON2aEmyf6Jw7dscTQEDxfNKTiyDhS5sf9PQ8YVLLQ2gDyjRsTseXf3rzL4EoMl
gUhEMNESPB+MuESU1kxpalawxSExVLUyUx6sxYGGMP2tuOtC/bM0e/z325lxTlHAfsUKnRuuvGBR
zWy+/Klokbmg9/sJYWJ9YLAtC1r7dlNYQ0JxbdW6UuW9YGQeO821H3O8TRGpfqXcdv4f7yJtpswO
6+NyTg2iWLnxM5ugML9XQAzJdxPADZDQw1FmUePpCHf46YBZYHgRGH9CM1VNExNVHC1vtQ5nlgiY
wXpbber4OJUugvU2xl1uU3qfTQzhyNkfnrCKCBAVb9OOpDfEhBy8b5i7nukfYwk4u1Ez9WjlhRma
5xElo8h3RkbieAK7eii41nqULHlNRxlV5/CoVCGtJ0Q/XV77DXg57a8hZW+jbViGfaKQlbLWPhig
MXaGmwW2NHvZxa/Rd0S33HQJsUyqQw1XUg5ejaTzv3F/niaVkzFcvBZ7XPfVtrepfAORx3UirtNB
mX8X4th9XCDus9bG9U+VK0NVPvOJDwm6IqjiEmkGtNIgXF8SyXCB4EK4cUZfR4474t+L443rQdyB
+ino4vqIfsJ/H4ISfLApCF0u7PAyhP0h3/sGYEf3AOvwDAXTegrff187C8/HLMTtDmRtVDCCzv9i
2P2TyF766s+h3ahojQ+6saUuoZ41LSoS9I3f39k9Vsqj3V51hDnBNVLfnYECU/84rdVjRV7hs0qs
itfxr1w3UKg2lHOb49u5a2T1pKmQMYTut1WQpM1N2f1rqnoaCcPL3VeW71lYkVzffOsM+GypSo+V
Y7YkP9z6g/KD8CmisnsnBPusp9Fv7ZjPu15FUDnA++Gz+DO+9KGxDFFq19N6wN1STi2TLbc+AI67
3n8xw+NCcvMuEOVo1FqwxPD80k20HTcFSYe5gj5qV5SUmlQZaVE2vKWPhVkTM9t0qNEL/odEAKxS
1INxPCjn3NCC8iVnFfhwJKQGNFOqw78vha1SEavGykHdsGdmktZPw85f8Av85gpB13dXkkrwzWyW
ZrMhUx+pkY6VzxGiebP3INZKFZ3WIE0RQPON1Y0zCNKsoM+N37lJFG2C2p1cQ5YWF7oeBh57XM47
4NmEbRtusqO8Dh27lllVxntGF5872yWF73kv3g9dp9M0Gi7DB7pSwekZuxZaUFysYm/xvMsWE+Ts
fFet0PnF0TDx17NxFFD14UbaN0s3LXtgpoAng+7zM2SxZvaDbDzd/ghZZSuExdPprQ/R49ZDv7y6
Kv69rbn31mmR70eji+GClgHbAEpVwUuX5STtD+69htYZ7OYwt+00DHNJfzJ1Lf12O5YKIfb+Fchu
v8/IXYIxF+FxZ3XNBUvcZ/IarTUwEUJxRj46LTdSU86gCrtp5jLBkx0xEticSW878j/mN8e4nmUU
LEHK0CPU3bxl/wkW34okQo3wgAEtX31W/UwJTY5aSFSwq6deTxp3BmKcO4J/ol63EUqsgPVqihkh
GN8uENPRonoggnYOHjfz/bJPzooR5fXdyK7sxbHKBwWOwHuKeWg/II+hwEw92xMJyXBvxtMaM4bc
xiNWeaezM31WFwAgK96IkT9t4XSXgSueCkhHTPA/17VBAEm3m65cztZcVwyEcp74RycOc9QUc8/L
B6F1kjtZNDM7iZESFR1DfZZtf/EtTMpY+8BwDx9cgLHz5LsqK0wJEE5V/8RFgqYVhWFxcQrziRDy
htsIwTFqRZJZs+ZAYA37HHMkWASVUIVUf94f8sMP1YyFQBZIKyCTVrhzRxEN0viPNFO6Wc1Mhfdm
2euTPw4XtKSoGwLwFKcFRLf6cDo3wet7IOJ7IasJLRurDUBdM4SsiIWMf6CvJ/WxjQVnUFIq7OHS
4qYYz4Hwcb/UPCOUTKDsQ5dbd5vRQzzdIZMRhJmH9+IAivqVNWYV/nIo3EwrHsHNUYOh2x1hT82I
p1c8Nc+Lm3ACSLXrJBoY0qKct3WAMTuaZINm06az9EhAKyJ3mHbH1IuO9v99ojT0ej+VTK805cUA
gcx1vvDN+HasfxNgSa6RG6XGEo2zJk0AEhNkybi6kMpENcDjH/OTP46LOfs0Xi4hqZ5BGxH+ly6O
QEvSvoVfVwy2+FD0CGs8Rit3iPJUh5T1hP5VgeJh/0nMt9Mndfmt7ta6vJgU1x1SgcwTV+BNlFqw
69eubARvuOl2HAv7jI3prN3d0Y3M6LvjgZl5nsULLOPQTnSe5ao+gXOZHTSu/khuQe6LGsICnZgB
sY/A0dj6O4VQZlCexZvEstnl5Fl5vZW1nHoWWxmqZntYaHoCmdUajPB7+47r0gZ35giTiStNCYoE
2qRCLVjKiG55JNeXR2BCyJRa1XqDIEJey9tSnpV86BaKzT3DkzBM2Wzp1Dd+AtnWGNuQv/3ekGQI
hCKZXI87kgRAgQ2Ifp2F/BoJchdvHilaXVqxIukRWxLby4adU6tf9p3AXRCcd+ell4OpGdrnBU0w
fyhRMYedTqNGfVNliUFV0aIvcko+V5EgPsWTKtRI2aiTMBd8Odf6myMnzu4wf/TkaK0J+qiZk9Wf
n5W/D7X8lot3BvqWEkpQgipV5iUtUYCxi/HinIQIWZQD41tjRTjrY5aQk2u9BbbDEHgUQ/8pgLmf
yn1bzEvjVFqn0z4KNECOW62QlE3ZKKDT/2eD97Punb17inr4Ihfe2qTUUBO1JuQoVzAfq2l61S7l
oDMzM2NoK2gY/zdWuR6c9HitBbVxGPMVdMeS3BBbFk14OpH0ARAnv2HdGCthzwHjXX4J2EvtjIEL
Yv11RU45GskAPPQfpzzLAEf0Q1f9gC2F+J4xeNku6HnMKwtImsk51bcJvxpDxpeYlHsFFRfhFBLg
N22SvTWjYb4OjwF8ku0tmlikt/wxUam+glMeVcKqJeHzDIcfbB7SGbX4X3uylQPJ3SrFpk0ZFthe
a8jhYRR2CxCmjJtG9hevxwKx4GUZ5xmg/4DF7kBjhwrz3b/oDZPaNjLpZKBMWTmn/0NVRUEdQuGT
VNgElpmGE0DR/QpZeH0gDPoMsYkT3FBsx9+R6tvPbFRehSot0Ji0/CxI+64EzmKZPmoUz9YgL3Dl
eaQE1b9RizOmPXFZhVPZCLJoUL69UNPpdLt1QdRI1Z6e8nuZc8vkoYdC0njBdA7/uspaCWLuJ9xx
qxrQUpgBaoC8wH2aPqE36gR4cLJnKEzB+sryJu9cbFNndoFfraHCdx9A9jP6w9HUkBodV+LPJAxi
gx15dE73Rlvo8qadlaw3g8Tkgb8xqkSC3HroHMAHt+vhsP+IYortwbAu67TcyKcjLpMfuJBiqkup
otE7eR+EJxdpa+YFrtMMkkjhRq7I2JzzPPi+QzNlDoEDiHuq33wHAwxlyw2IGbaZc5h1sVOOCc+R
4Rmn3kLrdrR4mK+q6t7IfSr85vAOyt1DVl+FFDKUALfw2ylIRFNH/lOqVbA5if0uDPqCmuWjN1kE
w6bGGWr+yM8I6wHugZakEGst09X2+usxU+Q4al24Z7iL2HUZRWiSZdI0TcTwXrAHIjhxzx710q3Y
GlY9jkLp1itiVaxl0X5UFGJCvuMCF9aHQce8ED42y/PrhZqnTzzO+DSj3+7BlmwECLvqvYSZfBA1
RfKGgISMfHSdz4XKIyFpT2ytle1islgl9UCIPNKGFiPiTIFvhoixkQ6KMRxZH2NNewQZAYB+bClq
HIITUekT/RFlyIQpb+0tirQTVPbK8HwMRRFXrNfSELOTs3k/d8Mj+htM/jwO/xfCulw+/yez4HSA
FvHiTL98leIK/CAafgrly9tFzJfT4EOJDquJ8F8S8iqwwPrgJf0WcWs9WLcyFDCt1E3iebOLzX7i
8gYqGjJYzotBkE1/3JgsBQuPS5xkJSdAxU3pRr4hedZrdCSxuq/ugsigwi6Dwo8lv4oNOZKXpUne
oXVMAQpGVIwqZxnlgDe0B5nQpiSwSvRH0WuAB7Wigi+f1vIDBG4Ou5fnM9eD1STJGLsnar7bT9JP
Wgk6af6pQ8XQZUkkgQxFqnSUEZ2XYJVSmsMKAJ6j503pr/yjZ8YaRHuhkBnINY5MB5D10rHp1/gY
6WA6Skg3nju3Ouw2MYTERZvmFoOElPtpaOtU2JUB0VMXSlxm+V2XtSGsEc2nMLC2tGU2y3POi6qQ
tJ5AYdmZvP+y6h451INDWw/Z3I+id4jb/rOn0ZK/63nYBw/EXHHN4tQXOVV7+lySD9tv3qum7haD
ZL9k162glBwCLRdFcJG0sftZAPGDL4sXWEeIAAxkiJnocPxuuIr5yif2+vVF1gxYzfQwlkedno/l
drsDd+So2LHMtNjMg5ApQ4RTq5adOl8j3g0GLVsFu/m26G73bceCiivqlKAtvj/D0fHY4zGHfPHy
hH7fl1qHB+6IAKkOCZkzdy5h14ejDPYzJCXRXxXcWOmh+WDFGhTevi9QhKvgrfiTfnXalSA5vaVd
YA6JdAXgNjGbO7S7n7ppGvMLBpy8aMtSmr+AZ+Z3U/6AFXL4tpuNQ2X5SRWxRBPiwxhfDR9fajH6
r56Q7ZLcANXGAbWHbxkBktfRow1zYR4FVIOtyD6RYArZc5I+ijTxtuF6HEqEAekpgJZYKXhbwNNJ
brLUOvQE9OT9o+L3ethl4gbHPNZDYFl+7R7xCpT6jG466T1+gXKcDRlRep2mkBrcHAD9AFpnXXrn
5kgwWCcF7GsBfb5jpcizpIWYDcQ8eKPCX2azzKYPjrBoen3PcaxVKDT4OKUaXzXU9A07r7kiW/Jh
W3ppXp5nG5TAFqiGAkDSFhmNj3qm9PLUKrbKW8c1ivBrANzNl8Y1qVstmOt5a49iVf7CRo6FdNzv
KG15rE0vV9Lvp8XUdkImePp0DkUJVhaLn58e5HTKL0QyhYga7ORqqrdRvLVTbHGX9zVvSm0PebkV
9C4SNpELfeyqC2Jn8Z3k5518Da20UEKnW/eCUL8bsKOxM4vbSeKIvxqr+PUsHehOchBTIbddeAk9
xGVJv0Nvyq6rT1/egwFOtrZ18FfC3ulKuEFIdQ7QRl4Yo5S70MOlgnrSOht04pWv96qLYyWaGInM
KbbXOlgRdtuZxk8PIVbMFgb6LzkzWomEWcqKfDdrigM83b6j4W/lDwHp4ZiB6pTPW7DIEYOH85Xi
YooYTvCy8adGGtmo+pkViuFx6JWOQJO7QpYBfpURdJwSPxlHR3zL35Xo4PP2lHlRf6mg3C0O2cJq
aFtwmYlNRl1nOnLFW7djGy2DNmurJCGmuRTNmCk2bvTg7VjE8gGtQ0wiuEtEhCzcsovvsQKXdt6m
7L37agV1LdgO0zqwkkILnFSLI65MDGdUPH7Oi4JerehTtB4qU+jbSwxro9snnSthJzDvBirjgkj1
0ZJB0ZHAqPDl7giSKNUla9CEOrf+doKBz1P6XV/NG1EDVnT8zqC247lsl8F6A2s23kPzh28lYHoE
Ah/J8laWL4Z5LHNpkc3+3o7C/t0ywWc0ULK0P4DxcnLUNcsXM0PyAGzOncpBJVfm4XWs36Pr245t
KRKPH7kS/dBeQyF6YnabKesxWOKcmlQ/t/1TshfTEmK6X771tHoZXFuZw+TW9CVT778ULp6029oU
v/Ji045hTTE0sKBXpC/EbW3+8Ec4cbePSYv6F43UFxknmNRyck5HfG+7K58Si7dG87Gu14zuJz81
nHh/5J+6kIz7dEjSUlVOiyKt/lX7ikwkPGTlKmidNDLDShk8ij/P15efMcZDdSzlcW/S6JqE4lrW
S3dpM5E8os7uCJz3gvAnNKnvapMJaFpUIdvwOE/QymRY/ttJlEeD7ichkBpyf7WX6LlnaHPNkKa5
fe9bg2LYqxRKh7aGrHpHqcUaCXAV75f8JoSa+/i/eYA9l7z4RdtmSRWmLwWANmbMLunIgUBV+umX
MBZ4GDzAeNcDax9qJLwYbxFmaN1DdcRmPwE7w7ehTueJOdkgwdO/ijPMO8GLWzfkxnmSv6ivabVv
pjzOxIxFCsWSqzus66B4FGj3lItz4rtENu9BpQ19AgoGhKtQkPNyzQIW8qa4ptszU/L8JINsBLq/
/Q1yPzDG1EBht3v8wlkyh30lS1oTU8PRNexjtCsyoGBQ2GeuHI7FfuDrrjF1APur1O0Ke3royUNt
mscyC+TfsGwltpZBiuN1b7aSuogGj6mOcf2YxJrOGEGv7P8IJa3gAXFqezFcXSBfc28LHBwHbHGx
goMqeAp1EavXIFrIs+fBuDjCRs38V67fzWscxzE18nscPjBCowXnd5wglbgNxg4b7c1TeUZnTSyV
Xjkg9vkffIO4MYH0geal6sxtK6SKr6VZpZgPNqIz7ilJx2arWMpnnq5VQuL5TsD6FmhYEuBt0K6V
ocaZKcx20p4Pi/3u12jDC93MBV2kSGIfO1Ys46kS4Dr8doA5OQI6RmUcHteffOUP4gvDJgrZcFft
Ke9Tem6gQj/vXCJej35wAfIUijrq4oEuDb/zwYaRgt5bwWpRWM+3Nl3qeH7fp4bxC8+uZfk6EwM5
BwKWmP0QMjs6GOtBczkk+HWkpOwGqwCmntYsQohbG9tBm53jSe3gvzgc2krGexS9kssCusVjrOBY
Mg+BSH3snP6YlP0k3Wio2/OBXv3cu91IItG2JssDMX9YbjqFSUBjECSoku76GBsXoYz6fFLck0Xd
keWMerkXNeQp78RkzZbRBjNkbACCx72cFl9RX41cVGMTCucqaBKz5DNrgTQiajvI4bczueLq1U+8
GA1VjcJ/XemN7iYnjSvDD0kHdCBQNgpwHVbJzPqXt3AlikQiZbrhBfdA3SNA7aBSnZapO2nxnLkN
12brsICP9vtKpktD40DKCtvUXp2qvZxPfA0bx75qMMNI7mAlCdyvNN1GXF75chZ6df4CwBUdaICI
UQXMmVEdlVnLpUYYwDiGZ/+4C/VIQhPNWX0Tth4AVvoYiF3KgJenfS4qA1qwdfrYDNaPPz/5+HCY
PLuet4CW1rrVK5GISmO0A04qX4mAHunaUT5KHukQSVI20nDWtPjLR8J1Dh7Mk+QR3BCm7tY7kiwM
uKmyObfY3vGEFNz/H22JOrMeRPGVABMXDGTHa8NTPBNw+0PGX6d2rKj8bzlJjWG5sKemylXEw01g
Pu06zUNjaRtjDZHgSTyF1gKd6C1bP0+/kY8gt5fh3ax3UgD7XPS4wlWpxWJOVn8Tzo5T28sBZMUg
jatxa7tlCmWAtNv9UqOIA8UdRQivgSEGvLVs7Jng16YdO54xF+BGuHuroO2M3O/EjuhW8xygDnCb
0tAs96cAw1LGtkYcuyPGZ4lL14wvrf+TrYyr1ns+dwVKXNopa8m6FWvI/ZCR7J/YHlk/Bh4H04h7
eZQmY8+3eU9Ix0ZWHNej8briu9v3HXS3N36UMG1AlxnK+yWZh40boT3goR+UbpEfk8ZVfixBUL4+
ES2n/q/jAVmzaQHANTFoQdb4HpkzjHvbo+v8ptVo05BGr+sR9YiV2stOJzkrDRlBwcMHJRbg0X4G
dbxxzOrDssyqNr2+Vxn2J3rwT3avo+RvB6K5+wCkozP6giGf1jFuo9EOFjrb7nisgG2Jacb9deh0
CU5cEpoa58YTzbl+LtnlHkiC8DqCCAP2sy/XLfMb+hcmhhh8Yx1+U6Lw3in+NZyox7Aw1cYkQNyB
IrUPwMnYXW3buBRiEel7PSp5PzNWpnE37FDqtJt/l0dQWmY7LvUPB00L08gKeAEp8cLRSYCa3XlV
HPX5zvYlK85hQbQHmLoACRJITM8EB6Czi/lGSrSXDXPN1C+LOIPUmn9bb6CsbmDo57CN+IPM32E+
pT65SZNOsxE1hiRB8doL0RTJi1XNiXUtUnpYddOf3kLVexMiPrADvf47hlLeibD9bybUlX1b7mmT
ZpZetZ5o2tdAOo/ypO9oUWmhDsYNfMz2YT6r6k0CZaNPOJfVj5bDACU+aBtAO0xgJ4Sb8hBHtNkw
nCGRErm6ZNMhIWJp69LjWVml7fmUbPzFbdbesrQgnyF6J5Ht11H1O8XP5i2+KacNP1BS73G1C/45
JpRqmkW08dLNDC4+Zgg9aCBkz/SJTMslGuPgb3ppJWknMzNmR7qg0AVkrqv06FLAjFdnbJ5oLyBw
W86ZH6xIYaRjCNqiDPGfH+pH2QHrmyOT9MAzvGigcfQvaxObtdvgn0Ej/fGp5+r+vuq6nfNyJAFz
c0xeCQcjs3ufGAAqpo0uMfFhVxJUEXqAvLj48Z7TICoHWu8odANRWWS61I/b9E7kSsCS2D2nKGE7
QIDcCLHeB3kol7QtmvzJ5q1Eb9r1luqQZSlRHtxnb8O2YDTePDovIsfFFbZUlX/hPCplfZsyMPmS
gGqG6FqYR9OfyY3FYn36UDC3gZdHXFZIiBQcmSl/OQH2QEzEF142Aa+dHcVpGvbtgr0Nge9WfCBs
K0N+L9yTfpt9pLBWFyXatQUrlCbspK9R+Gjewe7uwIPrB0U4nDRMK5EQUQyx/n9v+hIx+htAvvNr
DJ345XcvSjA/WcCPdI7evT6rnnsXRk4e2p/tRr+I0WJRtkQs4a7t4b/7BnQqJZ4vvMD6xRFJ2R7E
Jc3vBOj8qO5fpoRpnyAqaU9hXk9H0VMXqafC+L/PnDPpwVj9pUiW/ig/KYVj0qYJgLo8Bzp7GdOX
Awfd6SGhqfm/vNCbbU7PVTkf4MCn/kBl/lMEsrsEom7NSlJApni2umgEcxVr6VZIaZi5oeybCbIU
7KdGMTGBVtqrIdoWxrx8uJdipXHD3qmiHBOZj/3YMZjd1WMZhsJlPPUWRLKhtTtaxbqqqCirTs0S
5VCvupMeRjw//diiC5S+dpNetptEKFWewB/6+Z0zL1mKiCx9J+AK+RsKrUhM2rbHPQPJVc9nfqLV
fgpO4Sr8kXwxa52DE/V9kQMBUqF3C3OXFGs85zqP86ZjgbJZ0a4Es1GQT293tifjsCfGvPgYzy62
uMGvUSE3MAEdkk9somCXx/e9k0DjmMhvi+CeMroELmZYwOJdg6GXPK+OQU2Nomy3FdPJAiAfvz+u
d5jEXprEB78izduiu2njcELMR9QSs/L1LduP6bWs1Y6LTms/wVa10z0hG4xFJO7AJrWGCKY5MFrd
W8Sf8FqfDaVV9PKucBkV9xX2jlDqAZeIbL9nYH3meJYPOjuvsYfbqPpz5KFbZ7kxdORA/x9koQMH
Chbr8bwLMJCtcjfHgR47BQQzrKXoCK4rcjg4z/BOO8EBQD8wtwbvkeRqmmnRsPkKWdHm54b2pujF
dH0p2oIEmqXmh4rKFw3GD4BmIx8oM2zBESzD9jaww8d26S34BVaUaeGRBIpgRSA+/Oy2RqScvW6l
uPYyycdLsoqF21Nh+3L6tUVwUxu8ioePjbWllrnzUjMkOdcwaqSlVaD22pUqU0irQNVb/GQVX9IX
Lr/TSxgcsfsLLGa6PlvkhBQURUy0SJHgAO/VCfCPQwtIMYm9s7B2tFBjQaoPzv/daIRxluY8Ji8q
jA==
`pragma protect end_protected
