// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
jdCp/Nhb5qBwD+2RTR0DVA/1gPM/NoquRE9VgnhOeUFuqVCjvJE1bRDIWGTJN2l5agPlkfpltut2
hNQnR+byZnC/tQNg9zVmKV7dR3HlcuulDTQ6rhkkF/C4FBlNzykndMPbwaTQ7uvkGYE5hT/POLVQ
iEfMrS/RQ4PztJq+y9bf3Vv//IBNwqeBSvUPJneg0M/8Cc7DRcqrmtprRqNnlirakcP0alELF35a
lIfdr/z6MgdIQ0rYyrqYICpD7Cj16xk8nAgIKAsp5kzck90ck1Aq0VzkmdsGjLAy0MZWiEW1rnYi
pCIK7J2R88RKPFVGU93rkTNvXUQDVwOBSAM9AQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7408)
/HxRv5dfxu/mJS9xUTvsMzkB6hfM+47DxRGYwdwwCDv0eaNnXIVHeBb7N8LuV4CCWqpAYyW81uBR
Q6TwaeHyIwYOG9lMRHdU8YEwiO7pdvJfW41g3zkwQHQZwHGZhU/Q0m7MAGlKUdE2BlN9OEokWTIu
n4J954lDu1YA1jGSEEYzanvEo8H14EN1JBn8TU4SlaQ9e9BagFMS4Yt+QgMso2d7BEWopJlYBg+g
sHaIM4HNZg48FWtTyYdkgqETjjqQCeR3+kmliwDaJoQBnRmjD+uDb1tMLg5y1RdTXHpFq4A9Qokz
IkVWqHiEJdrqUsIL2BdVXV66fKD1dXAWJ+92m+RgPyIK3CzXIXtCgTmpgF8WOAt82mQYAbjgnbCO
vT2z7NW8lNCCiK7AC/9ojSP5eNAij5lyockelat8onV4RaiP5MlWJb1I7TEab/cMRBmTxKu5dzQ7
wQZgJHLN0peDpkqCd0DCbtXZFpFNohoQrX5tp9XNPWr1lQl0qbCpcBuFPPELw5YxelsXPOq880w/
W2QMde+BNfTX4ujVylPo6Wc4nibpE67lEN5N1bAlsWOYKVMVcSTg1MI9tRML/X6jbQg27cs0Vvt/
RAAR8ZmluRdJzROe54bYrzTdHYx4ZTVYxD/fHxcacELko+4MD0XG4M/3wxZ6HpknkD1ZhFBpnOFn
t5cV6W4Cyuh5U8GVUVeJZTNjs15+DOlwJPa8btOrsGE7gWMAKjKaQjO+yQ2zLr77+EX+L3zYEHpd
Siq/cf+tMA1yqC9crPGO06AY/TI+q2nBMbmBAZYooBBpV5sp84mNJ0RFuyFzZXXidcLHhC1pSOlq
iyRDUI9vAd20fHCojwFqDONv9Xq0ox6oAr0+LEiseCeO/v6yOy0hCsAxbHSyjpzCclHaehASOwRl
EOSnciFnaT9UNVEf9aTcnFi4c6105pwMzDUdjPRRPmLKN0NKV0RApNs2JwYSfJjILCzwz8k9Q/bn
q3ia5t80a1P5c1vHs631kbUZoXuo/F/Zl2SXYSTK3md2F8Hwjpt5BUmRXDIR1LWONRl9vx3cCvvB
9WHSI87OTZ6kV4QVNv5eUbiy3L39fhTFXxyGYqK1nRQYte+S6yrzjjAhz69VNctG9r32ZTplvWYU
Uyx4do9tt5XKNVu0TxfIWs5Xh50moP0fBeGT9iHfpzlLOTWfE/OvMgbzwD3CW9hzRyEooT2+6aQn
wuYJtiBdmYzKLF/b/m8yJVyHvA8jXt0nR/yI0TD8B/3XdpbQJCxipUV0RaLbgjPxqGYCDPANmVCi
1d1HBldBgdzl9+yKRDJXJNQfsnXFyTnpm4HPDgp7AAhN6he2jx2BFmJPAPFo71C21lc3pDOhkD8g
p/Mvp2/7+jJ8d47cn/wrH38zUnVz83B+rzfSJ9QjntZkPXvysyT2kOabde83C65cWFUm7v7wZ3LC
ch8YPRhmtQS+v2fnMpW+sYS+fk3Uu4nHhtCw0yiy2SBxij0JKm94kIXJuc7TXSeskPz/ad8nPewZ
aE/dlLaIWAXwQjNKzcceOUjemXsKoJpV9T5D25NAoHmX0Ocyof5oNdwVfTEcb++gIxCbfy9EUfAr
HfQ/MSugjcaKq9gV0C0Q5kQBAtEw/k+sN8bg3WjyPPuAU5EfFvL2KOK46ynzBlyPvtpgOeTVRPK0
8yubAWiPqbmipctX4GY78/es4HkUgAlyPKDa+w366acnyUuR7Ph4PxBE+dJBe3HhPim0+YZdPW8d
PDiQYjwu0LaQS8q+S+JKBOV0+g8o1yxnrsrt8arq4JI5iMbd9sBolfMdlzBwhaw8auuRLZmT5yj7
t1y39qMLhR/yJELszzi6v98Jvld0Hf4duhJrtbUuIat+NnlxLCYfk9qzTkc4OtU0UTZGgwBAJvUg
EZcGyspv6nlls8Tx7xyz8MGDnZ7E0F5+4nZRroNMurSdYqkWkr32JWZFGs1Ozbg45dZg3p5bI3Hk
pID3KfL+fna21sX+1cTx3hvdsbnddDKXPk0qXCViyI4xm3u829Jd9Yf9R6dRGIWrWc1fsKiKoXkr
+qjiMYkqr/jdCE5QWXxF6aNISjVaxFTFNQk6jPTii7/Q8RVP9IEb+u4BTaSDTs3671KzWxLNh4ij
v+n4C4xCDVB/R8ILJE8IEQ4tA5JE8/TFLe8eidocDdVhQsZ43kj1iCCBTYkRGcIjrqELVQuu79+m
/2kGu19N4VyywKH0bjwot8diysohr4/Vg1qvpC95PyU58vppQjiDGmJ5bYP7UzuWaQGWj6SLLKxH
Fl0PDzTX86j3QziblAhAuyHPnVZyczMRccZ/uCynObr7liIwqWrKxwt3UXxkLXQilxv1t8Y51ex2
Tc593bwPdadeiD7pmXDZFJ6AiDElMq6ZM+0+wjmIquN9MILjjrU/UV+5CRroctIlSou56ZrzeEoK
3ZjyN4ZA806d5t+gKugz/PJmkugb5bxZb/2qmkd35X+Ww/l4zdvoqhL/znFW0aqJ4ymQhHiUmvXW
7ipFQMYXTU71W80Tkx30dWDH+tG3ez2RJGf7xty0VfQy1jsyd/tUdXR4Wsbp1N2muQpXkiXuNTHq
ZtDYo9cuC2lhMTn6vKO366kAwvvr0OyYvHtxTzz37BxUTkbwrpyOruaUbcutfpXZHkwqnm+dH1qV
Ddxcm5RjlZZq+NI92OPVUZVZBHuBL94JkwKE56A7YjPKJ1fpZaSK4IT0smaNMFoXvJJgKIun4gJs
8s+O+9hbxpHmSyBNc2IPCygecoW4nX1eEt1Jj5fCr/NgkiZu2+YG7bXhE53ab7uJzepNym/HUvTg
XuD9Zl1vK6USckLaESUQtrXgecPqRfhoRqzRGwmRi/TBNAfZLkYT5oLkQYw0Ur9QwP0mX/AWVvZH
qnrS8U1l3q1dT7HVQHWcaPJ0sXBvu3v+Lm4LAaxhpnaEPBSA4Z00sAMBEkXNAoKLi30OrIwmwEm9
rm5BljhEXCwYJaQV/4J4NWem4wuWoj27GuPEiwZ8MDZYM9sZy+mHBdYMAHesKJSwaYHs6xbPZxoz
UNNKP7RGySVMbrl1mMX2AoiuWQO3JV0PtFaYxZThZxcN69KmW/mFjXpjZjBwG6uCLA8uA6H+nan4
WQW8hvEVVD9Aepd/qzKuRb+dDQtOF8Cq2Ru2nBqb/9gvZMeM/By+TLnOX1AVGBm3V1ngVom8FVte
tCBW1eTgmL3WWli0jjKBzxPA35IsbqKtuKPeCDvRnH+v3GVbXMKpi6/EgnjKMoV74UHKGtKkeLPY
aEO1v16nYopOX2vQeN9OnL/xvInSBLhniei/AzCIc/ic+CSvPRDzzk0TLUuD9f9KPmLOxQCWaOMW
pnf1kXMOC2PZS0Uktcnh+7XcvRAAfpeno3fiu12GhqdF/hSw01BuEwtXhxgqqDAsBmOi9R2RUoc/
VEjf8tLeObPcojYZXq+qx4OfBUHIazEV29oUxuzbkE7jLW3w57WC1O/r8baMNEq8ZiMQOzY5THPq
Haxc4alGIQHr+A7iuCDRHSArKGacmneresQgGJVzNFE1l5rht/70n7HE1wTq4KpVCRK7KGtPU5vp
/fvbsXBMKuJecDJoAAPWnSXTEERglvos3Altnz5wkWzB9L5bREWLgKNrEM9g9tJtFHdreFiLR7QN
Z/lXRyFgTnZLkfC7xPYWcxNYhzr1ag2cm6k5DD1iaHI0SkLLfuhj2imOrooS6txxDo3aYpQl9H2z
ut4QGaAPj/dlSrOZ2yQ8iQ2VQOZklVd8k05kS299F81PHDsygDosJDCYWKyOK8BHIRYQ6Zso0z6I
ZwtusyHiw/LPomwwZfFBACGiwVWqFxp7W83y7nxNdW7CY+MevtTp+M6RBUC8PwCu59I+s6VZrl7q
tlEEoQm3JkG8P5VMd4yMPejmOrTL/0+hQ69x6YX3wavI1afJvNTM/1/f/gDKDwsDgXcZuxF2ykM+
0f3Q6kquowhlItA7WXcfn61Q10s5I11SE+8oi9yU0UOgsevRp668UbYxm7u5Mo//nv+N0ssWQtZK
0jIvXzd/XhEjcAF3OrrZiuPpyPAZHJ7Kcf8Y9mNoHDvCaG34w/K4V1jIEYZ16k96VhQMiT45Aj/z
i58xRAWkCozyPBAsaeVWJQpgip87XzBP0JKd5whx66o7OLqKSef+6IgY8ZFnrbqL/yvubUuUpRNa
Xw/ioLqxwqWBlxWKZ1NCMEKvyVCZGnmU5CBjLpBGucHIRiUmgAxaXnKKkldg2cW+lBWmwfz3/A2+
bAw5eGB/19MvhYwy0IDOd41UGeb1Wxc/gAuI6yj/a0YhH09peCUoLnx1sjtQes/jmme/Yy3h1CBT
PGAbZEmwhwNg5526H2N4b5F1WEfTNx2TB34KdM5VNQgx08PQqjRf6P7M+TUAP0KoAVGIURsnFdkN
yASPTKxvih51c6SxCZVuBG5wsP2U9V6pR0gHK6kcaWzH0CeqyAMiwLvPDPJ6viArDIcd1F6zN5Tq
ACHmiWNf86UJtUKieY90+rxNdxF/GfGaMlvU0SmcQ2pdsxNaWAS7Pj7m36g0/4f1uOrAJt7QHKge
U/WGj1iG6h/O88HUpo9ifgGcUn+ccKro43bAhXtyE9owTUw6Y968kHiweOe0t/ee6FVitGA3brW3
UJHpA/daTqtPgK3lZRaNMUgq+FCWDlN9oxxEo+tWIRV+JRopbSoGkSxt3PPOwzkqx1kfXp2W4Sdl
7LeYfmqV5bQTKM4BxZuUnt73KDvaXP1T9GOFOW4tzW1mKuKZ5XA9mnfnfSFOP6lNYujzPCfkenp0
X17OssA9+zap4jF66l+SGpoyz+EikAHbHoQtp43FvQvZ+D3MET4d60akd4bD98Cl5yp6ITmd7zRa
VNloczHX2eQ1cRgVG7LcGLPiLE90lo7ZQBU+ukwqSDZ7tSgsq+u9hxWFQr5jn5WPdVROin6lJuuD
nfJNXS/QGS9oeELqSB9W9jCz0C/e4vSRid/Bms5J3AozKz630+zHa787IkcIh8JfvbZHPY+iSE34
xFr7T9At6E5LFm0REwjyUWfEArRAv6qXCpkwzqvs9B7J6DPinss9WW33PVjH5JwJ//QZDP9SPZvN
zNcQB9t5ox/x6aTlBXGT1E2BJFre6nwEzcwFZJ3fUBlxPDZ7popG8594siXRM433+sRfyq1ItDjC
XOwC7nW+xovIccqA3CgwMuwrthmn6zb+rF4yW59PmNv7SrYq0vtMouwDbxE4HU5G7PsKjQlg9hY1
Sei8iUA2m+VTsJdqNH9D4M5M/W24YgdAZVzegMU5h6lJlgBHJXPPAonaVoDLmXvoED1W1fYxzlqM
oNbLQLXlxy12/ARwhMFvnvsGcEG89Qxv3vEEw991rCb4zLxVxVa2cvoFjwdox9We/g26yDJe7olF
pcxyyRMGKrN9RPbRgHKcdLcDiv60jvMPRVRrf+sVcImQrgE+Qys8+Nt1yLaZUpQP5W9yGRCFUeWD
DSJR15jqCQrBWC85zE3hvxZZKb3E71YE03ynA1L+kTn7SvTz3/iEhR9m8pbUkErhkGlAUcE3yjhq
K+DDwHH3qXCq0/FVvIobM1la8IYuzlBrNG+vgOeCyEXVlIvTNU7fiLEAWAhc967qe4mqpNGe7q/E
PSgAS5ykE6n2ges68qMKtaoun2D+JnjTv3zEKhnkMDRfmaHXzwyQ7SfxxrewNX2aDcMu/HCUc6xu
Wke8IUhjw8jWWtsFzYnK4bz8scGRwIkgqUI2qLqpRmbs50i4x517vEw50/XW6rCDf97LIzsjPjiF
h4zLsUkvJQ4ClUXAa9i2Lpq7n5Jv+DGJrXJF05ibwowia+2QouYiQEnvlALDGHLSldQEM95TG0xU
aNwZ5chFwOdluuqTLc1ocUu3SP0qxz5OfkhHm/Kj7BVnfWZagkValhy2NXpMZUhfL7afbTHpd3Qi
lEfa04X40VveLZVFUkU8vQJ8ASbONjMh4TkHTvpMdYVj0yagVhKa1FqBbzp0jCb60XL2vMDyXhzH
fCXDNlJmTjH1O1mgUtAdJTzlSwXLjAmLzGk+JcNsZXbJ43xZKrcvnyITqi/hLQXOtFp+IMsw589y
dqpcMpOEEyOST6lfj1Q7hELtVbCxNSKRz2s6jUwxwBQRY9QDzHMm9N/b8RJcc9BGnhJepne9xiRo
xf+yN3a4yQNxZWq1oegOfoIPLHbC2bo1xlIo0EuqReW8zOIBGzqVBBD3zofvceSKqSeMHHglhJzC
+3IVGqu9joZ0bnZmhN9T4NWiaE4YGHrlokzCF9F4+1JfxZIHBtqtGS6kLyfK91wTY6jx/GPhF2Am
ANpAoMrUXkE6LdS0Iof3HAaAgMQOHWhUGrSWTTKTOd60rS5TkqHDx/dJdZh3q/7DxbbX6IPPb5uk
2faiz29e4gZQQEOcpkC2bXciuULvPQEcfjrWKTeCX8x6iq4zHOsY9dRi6OGVDHkdoEopEC7jzbSc
zw7NPGyR7GOue3/ToJfJ0IgMt2ptoiYtBpbsTm8ehdascosl/HCerRnoHTW/ugg3KAL8HliX/KP7
9nxHGhaCb9NPWSGiWq01fbpYB1SzEp9D94u3EtMW4sRSfpXmNz1B8FKztf9KKKQBD7wYGRXlnI9z
EEz3e1YjG3gfKd3M19Kk6vhKywf0v9jDW3Yi2z8jFn44CPyzb2pIRortaNff9SqFWfAXxm3A0koh
60R62WmAPKB6IQCPEzcs+SHDnhqOEdv0W0g9w5i/94IkMN8tV1ROGZ2XSux3lEh7x+rzyfNqh4Jt
vRt/dhefqM1TawymlMIy1AAAIuEDtQ7heesJdXBoWuzFZAXHk0wfaTn5Q/HhC/CQJTK/VMBVDL9Q
DsKARdc1ivqD3v/GQF0wMqIYFtmvUEv1393IsUGXTdEwMT2+ZPlHbxkGAGgGlfKkvSJjWABctlEO
VzWv4McnGmA+0bGEvgXPpUJlDLVFr9b4VgQHp+XckE//c9zmxnp7/rpJOHjjKH5d+uS5Q2zYo8Hz
Gacb7jk/BEIC/MRvm3m12OM+Mq5E0b4SiGXvBQbbIiZ9N2lgzP4m7xTY1GmyDC4bVvj3vhKBKBto
9gF6L2BYm+xJrsv+F1D+mIRs6JOAMvEwqOtFySLdjXPzOqpgD8YbDh/D/VKyBzeYzlAcKEEs5Qs9
Qr8U9GNj7tE3Kx4SxwK51KpvLXX7661f8qwWUS+B5wdI3ouftszAb/558rr6039Tpu8J4xrdsMS0
Jh4QFfk7mc1a0R1Ye15cZRm13Ku/zJLZ4icly4uxVaCpM7pMJ7ndDah5rk7O5EFbAh+b+tcHEHN1
9fHPtfnA4w0RUSix0Fl+4wDpKWxINcyKUyRYsqCrjDJyMNW02AsTj6ylNr38LoyR2EhCgOtReR0h
fEnGVtIvKqJHt+XQPkPzq+UPmC45di9UNTIqZe61aVtY2ZnJ1sokzGjTpizh0B4yYYSaMEfYD/md
xc9OAl99dK0MK2w3O4tdgrEeu2Xac4Zr84LE7yCYRCZ6r0uYDPktr1hj+MKVAwVQXAj89bP/5aIz
ptsGexvNiKtUKqXSb0vbnUO/0iOOs+P3Vwagb/Ylp5zbyZQU96rIfNYbjeD9rGbUF8q42Ean5Iwh
SCM5wPGyVso76muw3a4UpVz72cj3kolX3dODAehwGuZLgrn2D+dUCDDz2I1vYA6o/rk1rjEnOtwM
lTHnc9hFR8/BUyrSYroeYK28LsMXGhaBMq58Lr94xZXJKdr9/vkmmozPQs1sO7vht6k3dbNTwvud
H3dbJBAz4xNSuRAa0Oq6hTSueouVyhiwQM75F/900jODrkhTU70mracuTbePTszYEXion4USOaPa
8u/wsEzYsimVODN8cwGVvr56pTxx56BmPAZK6aB93F6xFAPKTKE6fkG0gLlAHRV1XZM7Xuz72vLr
sxGNnCMAND0Pgjbnh0jii4ZNkrV55+JehLcbx8QnlxhYKcnIU3PXgtIqZg1wJ2npIHt393BmcvrF
gnHp3FWieNRngaBozor22fJ8JRGZcvfFscvVqTX5S0qO1stNf8gxJ4KbWKBj/uu/1jcg1PECOoP3
od/YP39UqCC6gRqnYjCGH73MJJD57n7pOfj41NbY0LPYf9vQK2MJJtfSxC0Zg0Ec4RhdMMKEYI4o
itj6HsElxWsKveXGlhsOM00uh3U0vsXAhmhaIkbAuls3NR6VMUn3HVodrLNkXaBHyjCcCwyRTxSs
6T7PkPytd7qGqjzNLAPj7qaR+TfKelVPu6Q1n3NQsACxVEYHhdgYs/6pXNCGNfZ5gmv4c1VQqSNB
2dLpn7kv375EMf4mD2XzN2Lb/DBM+NJoIU30rFqve+4z2tgmSHA/tMgWkqUlPmtUPClLkFyUXRFq
itZAwivkNq24y+01+7+XHoD+dNAcjsNhcWcTLeJ5oVYOKGzbYhj/jLuDaOLfPQvWK9aHmLQ6D5ra
O011EZTS42LI6beCpFEvx39Sl6QpsZlCO6dl2lgJjjDlYvbwQ3Zq/RUdibuKPR7t7htpSdJvfAg3
0TFokQLp0j6S57uppYbNmP8vjfI5lWoXDRzEEGmCEvUq4SMUpM89DEEB6t8UfCvODeYkjcx+I7m1
LbfKn3NRRZMX+AeP40h0u2RkCLfOAjaNn6U1bP+vlS1Txyov7uqWpQTrvyncG0q1TCFqrD4ZKpc/
D3MPBh3H4Do9pn5papsKJlyyhzGX7E7CIO0WzaVVGo3KPCMSP5v5TB3I4xw9vRuBDFS5EybLCU8l
G/ZZNtX7vwBa4sa3pDRav7dHLJnbQK8w4EIARaQh7cYXbgZbPiSgTfTsu9tcuuTSle7VRwfF+GdO
+p39J+3b8O8n5tGcMSKZQ7gm9drtYL2Zt/w1ps4xEl0IaNrsNzdWZ0G/AWFwAjIcXM12102CHOTm
mJ+6oMr6ICWOmduVnpNwLZGGyIbP1H2OZKXG9I9k5eLyUHSw/gAonBQlGkyT/M7cOwuqS8e2JNYN
4MkMRUFy9fP3HuoBkM+FKGthKYOMynF/AzUeqxar/dh2YwjWoVzv+4XDO148DxhLVbgLYkEjxAK8
9K1/srKiGG04a+gAjLcm5e9scvMF0ox7q9uZ9ZRgSnpP3uzKVGgabLd1e9B6K/xW/tSre4sjANFW
mHOAxKlH58IL5c/wR3z/czrDSyEXFP65OJSpqAhsHYMvdKhaHIv0rIzzqNEz4oIWoFzeAyFbLY+t
UeDmug2bnMYSQW+Gp1lncvHcpJkuvZDLHPxq1KS55TGSyiX8yaX5QK69yQmvzPIMTTbOj1A7yq/G
J0pUbGP3OgMO+fibeh8XPEbMGXE5yHsXX6Tap3T2LtUETP9FpnUSjVGLI5hYNTg3n+mQ9G7Nt8Yi
Rp4Hubq1amCBqdNxhurJHItGZmOtfrfGSN0JItDXOdrxg/cLZ7NxLmuAitsIxrFPZYaczPnZgFW9
pvseQx/TZGuLgLKsd8uyF3n2OnoB0rUVGEsgH6fThDGUibOC6TdPjcbE3+syaDNVGHRWywypRyOx
/6jMk5ntYBPcmfQhV8EDAucl6UR89Bf2SP7du9KabwEg3iGqMMsD4ewDQttbFo7AsABl7tMyF5hi
Ln6adClNuLvQ0bdtyHbTyoMYpfQH5Xd3hxxxXoM5wWaS9t9ZHBcuHBqXPkBGOckPAGBZjE7SBWAN
4kl/ewm1MqB3X9b9cwncg/749PQ+RLKjZxv41XcPGOBeW1Nfkw8WYb119DMpv3lPJhDM13Gmvz6I
RWG3ogqhoTVxXz9V+kyEg6pvD/WLz+Dncp9n+/XTQnLsmF40RIbg6KJ+gK4y2lqeqpgwrPCw3ljv
hnE2/XLSvGi/ZY96sL95DU//DVMasqJ4AvB9++GhFdC7R79WPcLXAK1hG5NMkIypErDvbb+tQA==
`pragma protect end_protected
