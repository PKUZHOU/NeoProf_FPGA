// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nFzaEPKo5ThQGAhoWTNS/QrbtTvvWUXQmsj6TOJRwWd2i2li/8vo3XRg/L4h
9j3iaLco2S1JLje1SgunguE8XXBTHbOfYHgBdCj6ElARo3DqkwG1thOYrnhG
+H79XbBKB32R+hNoBy/HAccUs+yXIjiCRTm0/ALzQ4YO0ejgVCzABvSwFzU4
o+hz5A8X+nOuFamoHx6dTlaZIP+m9JZ7HFyIuz/RRKXsi20U4kuKYJkMlIWA
SnFpo4OvMZzyawlAVyiZQF+SLibtDcuwR9/qlXQbmtGVNJf/VaAJH6EnQjSR
ZF/j70kCS5RKYT8cQ80X8v2Kp2NGCMsFCeQbReUnUA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lhBssD/Xngdg1jfVXkllBRHbMyrqpTUGv1VXpByfoToxyKq5UeHegFWPG/xx
J8X+/QqWjYB7WUG2pG5aZxAxZOmTHVsTDUxpG9fUkulNJtR1HDP6ElzgBLHh
38PRxU2ipDArKH9E2QnhX8cJkE0e0/Sd7++Sn9CxhNP1I2tA7cWUTL/yk3se
WdGhGOp23qjzP790UXI3BBQ+fLXuBvOG+7FhQOhqsVQ7Md7KLY5FS778DgNX
0w/8/1muuz3yBeuMbqy17iOlf3KYIWsbjByxpSa4+cyJ7eBm3S0P65hnQ5ug
WxUeGcCDoPOIrc2E+w4K/I6HEskbOyllcdy9z1JIIw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YxQcjt2cMU2mpUjzEUcXu0ncKDFjH2V10NHGc1ccmlWIgWu7xtmqdsDQKsZx
odoDcYE14ZHVgL/PUMKT+3p2PAIekttQjMDsU6YR5egdti0Bfkw58Owih+TO
GAS3SRO04bnXp6jirtMYhGr+PSz/Iv7B3ZuvPl8awR7gCavLCAtR23nSxpB/
3OEVJSIjUMgIXwJdwbvE0cwtZ8dcdYlxNGArmYcrKMnAipsSoB2dvoNR381N
XdK+Xi+kUHc2pyRkkk3BZio/TrzoBlzdbfyN6uVj+e5hEU+r/nD9tzIxwVUb
wA8GSvzEH7vKct72PqitDUFMIzryU/TSQmSwuv7+iQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kt9HstJt78AElTi8feA5vriot0BUFVBjFMVjwVAvrAUbtyPIFGXcct+sVI4z
36B8q+G4UnxN1yqxD6hftQIKEGYQ68IZIuf8mT+XjW2z1XedqZMvfZ4JIu5P
cUYjAX4SaNBvMODT95KhEOwH83pU+r7m6Wy8l6/qviC/vAWsAJM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
hUrX/R5iog9bQJHhyWxF9SQ7bPhC7yW0hdZTAjfSDgDNTI8AM1lg+VaorrIC
kWk9ejXMiZrLTkfH7BPRbziuQ72ODc1RMd0/09WwCNBBItTGYBQF4KSRfLfm
7D5d213xYsddn3YiGAoNh3DKRfNVs6QebYsVLE89w7SqCDxXGAR8RgKnUaM9
NkqWKAf6nz+0d/zGLqRJMt3i72M1IDJ0nOMIfmqrTqPU/Q60dYB/eXADYs40
xlAIefHVCrNWdnI+z7qsSfQb0LfD06n8hl8Qu/rEU+4DI/jszoIius8rWbmJ
pAhfkH10yVwi5+TcJ8oGINQgm0ElAz256Ad/MKrrsw8FyU/jSz85UGGwt1MY
dIo6GOpsFLVL78rdDfWgZUZPBbQnNnt2/BVLqsDolXRTPjSBTTLXQfMv8pKL
UbAW0dTtNR0cMxbo5remoCjzvL9UwY4M6SYizSqzHi5es/Prt5uU+bjByGhF
WyWTCd3SLqoZC0Zdgw14+Y6VxdVK9BjT


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rgTjqvuZc/KMHPA/3JZB58uMUvz2t+/yUME+GPdXAzrCOX9mlCIsgGDPMRDK
Xht7P+YHWsM0vtKe23e6BX/5xQmTwhanlCESKxbLZ8TnP8lVzNDWDeUl3TY8
roJ6jpejAxX7AMw91HxwGVtpYl85mLB3wGQJIxwGDjSUkzLw7T4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Qwxzi+wQQYQJrUwf+nvO8kst0+nNUNuaU7mcSe0BHHpNiBX5xQg19FpsihYe
MjAZNY0YsodXn6jWGmkIYSS2SxBIQqbXyXX6kWAFEhqpvDQW+RW7TXTnlRKm
4x+onvcaacdfBVqZOFXqQYdry8GU4p7BLbChoDORXlLLGWA+eko=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 72288)
`pragma protect data_block
sIwzUMBUU2QQQRxKqxxsZisyjEPUFCLSsAc2b+dyjTjdH3BEttnXQYtXJPXc
Uv3/8BOVus4JxNT+ty9Czs47sZxGLdum81xph0bFLV9HHN1kGdacqYJ5aqHv
gipBw7y6jYRvdfqq3G/dQxYiFyk0lIGhnGLooVqhVReDaU7mlaMYiIkr3Cb+
hAwNjXkS1NYGhNDZojYS2cNP3WxQ3NgwHO+v2M7v2wKnZ1ViX+FmKajFXcQY
slsm+Lu0nHYMDvJM2web55yZRNTI2KGPdgPWbvm/3MtM74DHdG1fkeyY/e1x
OpQCIEGox1+oP93LjLPDL771JhQturBH/E19+0XlSxFYkhpXMPuly3yGLkyN
YObrp+1zACDOZKJfgIeizh3/RB3mHZphuCzQef48g6P71Sbpvn2QjJVr35RQ
jND4S2IJ3l8YCFQ3wUcA/aa8vn7tiI00azPplTDbKFSrlywhOIgXEYka7FLb
TGbk/xVNSd6wYw82drIzsC3alG9Zmdbx7blzM73RY0nbTBLgUZv9Rq1LJf31
ODCYDF3IwDRozf9ztPr+Pb/cNznSmcZ0f+ldP5gBA+YDza1zDB+pHdWJEUSO
87QbZk5K7KDcCjTX2Gwv3K07ZMvwpgCAj7NYa9kmPT1oPOeSWxN+lcg/IQLB
qd9V5fJC8+7uZmkkmOIThe7WnqfUofwJHs70cxAtITTvyWHwc7qLV/36t1lb
9Yx/fllVPnFNydTipeOX1xUMV31f/5SFuDYWVSqttMQgaoRrUcmf4d4szOAk
yJ8gxQwvvMD3PIPnDextOu3YbHOcsyPjwyLKUXYTetIR8WfnF6qZpNRxozJk
0elOhMH/3vU8W3cYKYDK62tvMYECJK5+ariTHqe1pQCnKVUvevU9i6L4SL9Y
PMPQw3farDliFNb4BWYgVagdndmiOFB4dsZlVtBPQKNWEEl01iWopqCvPpQf
S219GdsA6zwcR1nwobdnVQ0mXNWjKDCZHMYx63ZmbgcMYbra27ZsmyAx9CWh
4MEtZlj5pCdfBYM+avq8Zca+3wzEoUrU3SUXNCFI9KBgcCyfYzZmiSolfNiF
VII8XU9zzY8d+qZ8knwtSMTy8ykdU2ZOHRnCKCs9IngNCI4V9Kf8Wqt9F5z9
pTarYMaRdP+jFcNGlCMKbsK+RHa1PXMucF4ZsJYqd5bel08gAIkLcX1fqm5a
aw7za8RaKdFIrPlWvGYOnTvWmBJTwe7MUHYArkm+q8st7u361ged10L8dSG8
5CXC+K8w+zai6r9XmN/h6J/LfyZc5bnBEEdTiOnt/dJSkoRqMLDRbsc0REJ9
QSNLjV/85pSKQT0lGc0XCGsg/LhEiGQjcxkpkZgOeq8FPcgL3oCIuxJlRigd
lVygiH4ZgZ0x1ZefkH6R5hOC2hx0ttnbK0F3gh+XnPBooEmu+uHf4bF6c97B
Ykrxuh2y3a7d/HWSj5jZiH6SkFejbg2krBodArvlOktbIa7/rT0hSt+0ULXo
LzD1dWiksNpavdP0iPU954qQ/UA/EhvXfUso9vzWAh5wkjwjDIQSDKMm/3D4
MNGTr7VWqMffSwekEF4isyQFM/CLvPa2r+kBTVMZdd5p3ZgGTTqq1ifnrgXA
v9EPLL9QecMb5mfyz7eFwYD/rGO8B7gO8cSStpQ9BqaEJSwk0M/N9PtnZgxw
dd8OqIsC4raLQkqGaIXdS8v5ERzf7wIVG0d+plchUaJTSDacT+7lfym4ji7G
CzdLyyQaYf/EII8torQPw4ItwsfVJ9KTAVcnoV8sm6k77rWeMfi95ix90cuf
gdSk3GzvbMdANirW/jO1TAw4+ADgZtcPm1DWu7yeJrfaibKJ1l6n8Ukv4mBU
qUuzSrihHF4xcBfx/5lQhCHa2DMW4Ip1GSBaZVzq4eIFam8IUeIZQZuuN+6x
j2/MqYoEUu7FRwdWP/rYYXt1idUTZtSB5Dy4bbYh+F9V4Z6qNpLf/Ohf3eS0
9I/GQWhELjyIqIY0TkJoHHTrhk3bCVqD1eZtP5kFwv61Yfgh8uTT1yo555e7
9vC006Moa+ZH4/z3j6EkCuSLkm8BFMJvKMsNOzyKbrxe5eKogvDlGcx04FeW
B60AkzU50K7YpB8a95eHJo/arcvpWAvwh9ArvUTRG80FBG3tiFrJGIBFVtY5
KtgHwTfqjRMYm8xb4sSpkxEbLNe6TZeqRq0wacD7ScgqSjdouR9xz797Ja7B
6fsXJOiROdYBpoaTJTdO39rWaqsDnT4md0hbrA1UAJ00Nbr3MSq2ExUWtz79
xp95pW53k+80T2Jw4220VWqPlbhKW5H1miW1jixxQmQ3plC5q5Fqfi/eXpPF
K6qEsR/VYhSCmbom0QlPvkKLW4+gAmQ0gkM2I5+upYnDKoQJE6AMRDIh4yvs
auT8ApshR6qWUpVvMYnWvDYjpZuaoqTDDnhBXHaYl/Ew9e8IzxBU0tKIB8t4
H8pHAqasZuSzMab4EddXItosWp0Zqzsu9KR7ybUQ+x81Jk3HRdy33vkj4tf3
C4DsnKH20wfkExuEWHz83mleW2TXaGZnpsN/BD20JdCdMn+DXlpIPWuwnbkG
lXI+S4C75+4tac4AmSpZ4Wr1yWqMnaMT55mzzJtHCjtGCQNZsLuvxEaD+oTf
Hx4TskgqvhzkgY6In0sRdT75NE7GeImKIiYSIL8mhwO3JvbY9pcsChQF2Isi
EJFLVP39ote0rDwicQKtWIAoxfwklVdSVlHsQupr24mQLP0s2Albt+gRpvXA
8Boh1poyvdrCbC/oqtIH450Yn4Pn4JNadpFPiIpx5P5+ZWqgpVbTBTfSGJtr
+jx4evym7Jh3BdZdNoWhPHzzGFdsx5TY8SJmpk9NgsIkrEEOlRWT3qa7HWEq
Tlzx9kbE6/R1a+X7u4vm0Ix5Lu6c8p7yrgwfQbRbM/+IaRiQ/2s6QQ1ZeGYx
BF9L9b/eI7quIyOpd3eCGl1V+GZ+lCkcNsrpIU7WZ2icMlRPdZElEmLfWVHE
LinQ4vJAzFi/DHJt9fx5ePdJ3rMdPT2a71OnSX7pSJqGKh7oVp+MB5BHkUEn
qSPLX6Q4ubTdqie6j4Aj0CraZ0B41zCtxGerARrRcUyF6S68WxZ426ZKSPDG
3U588bZctd4uVbNT7V8+cYxyORDdh3T8tYSZm8yc0AnpMawvvrvnTL4x19ai
Hjgv0KAnrPemPxaEp9cXJF74IXQX8SL4tSDCgsriRWJGP07NsDh3RIaKGLBb
keweQ0OZavAW+m4f++TvGPHt1E2N1P6Si8TjN74f2HN36Z81CNU8kQUCypQL
WA8o9LxeHICay424s/zl2jk/+XrSJo8axOsVVkcS/8SYgfgi7P7R++p9hA4X
z6LhUUlpHi7cVCic+gxmHnzWL7ZriVq7nFibqS/5AJUM6zrSGoR0juIhaqip
PcDraM+wmEc8+jTIFrt9d/unWfrvucEFDl8heT/GibnKKsz2SSIUDv7qczWG
Ee46//AJO1DV1eeLm+4op8MIS7AMMSdi/Yk8oH1dFcrwPINF6iZ/96kr2N3r
HwOYpoNApfZhdefT8Y6Nt/mq9k3m8FWYuVxYJE2vgjCaKhS/QuyMIKGZ7hyI
8K1P/waObxzH5HOjgV750Wjs+o4IV7bmV0QIrUDMNlzHA3MfrBrS248rGHHZ
xztMrjE/mPM3RPzRAG+Yit2JKoJ0n8LKHdHOdyi8JIKAe++hotfqjKjyJezW
EXoU+YCScui8nYXvhM9O3nBgS+pIGM4QI1doEi79CCpio0lmJTRHmXz07v7J
qSOZwjMZZbHHw+azqqbba3oT5lMed+/Zzg/rnp/j+AxsYMkcNrpOB5ZtwuFr
+vA2+R5ri7n3pXlKQBGTlu7+dL2rU23eXR8gQUO7ihHobzBckIR08IoyDLJz
TJYtvLfm+t+8IHztcdRC6NoEdLSd6IH1F3S+245+trX+4KazOwVuIHvCdYGh
cJ4Ku43SaIsYer4DWZPpeIIk4rxCj8klgVRSl+bk1QivDcHSJjXKAw267zqF
2w97p8GxdtAZcuSGJ662K/oamCxKO+sfavYPxQk/W4WHXCH6dsRRWlaBVn5u
xkuKPZPnjEJblwlqrFtm2WUirOi6TKJoR/83pBpKX/7cYU7PF9Etp0BiHyEk
BT9nKsi1RMxMEtQ4TopHgWo8uemo+JeGT83MQbPA/SJwziWFC5WMowGlujRj
yvlwHsmNUxst9wjb+o7edRoKtnVg/xj0/BrsgjWJLwJxcbFIsxk6W+LyT6uf
uq8crRiQb1n1P60cMnY0ZAurmCMJVfRCtwhDVzFNGEusYxtJnc5UudHDRVkT
+Nh8srXYVd5AXYE2cfp5HvNwfkXYA0Q/ppW5JWwDA33SuFHqE9OD+V1U5BJV
CsikkDFG2k4kexSxFgMkdITlkq1tFdedJIlVHs+ZPZ7+hdJoQCLqk3H33atd
TFUVpKKoaGkGNbU22Ow+wUScbDH0NFgQPyRFBgIvQ2JFUlFOkrbGUBf2RJ4B
W3z8cSJEXoic/K9/pdtNSZZET6AZjSZuhaKJbqY0HvSG6jxRVwbQCMc4aHj1
+I+zEkUR6fddNc7rqUiuxqcXnsUzw65s4Wcl3aZo9eooMWG9Rdl8Yxpgm4ew
CahGQbQDEYHlF/zBzJ5y5UDxBr1z2+8cy5mtWI640ZOH6cdQOaP2gLHtOTXJ
dx4iLFHEtzrumr/QIwWuPrD6wk+Q3KGCLqQjLB7CPStvbCUUiY+65kI/ucFv
RLFRnbPJpGC8dzsdJ74skFpLu/cTlgoTO1aYWdqK8x5kcNQ8UP2Kw2OYFxVt
bvEYp+NQsd8Y0jAzoB78vsP+0+qrxDv1JUCKuOxgZYfcNx3FZKSEnf/5wbQv
rT42GmZ02kCP77WbzHObcBx4OS1sbiieJZB2XrwRb+x/LQgZ5UqBGOZc0gaO
c6+UnT5fiq2fNkMsoZOlO2RaCblO3K3CKQknLCxtnJps1blMprE3hqp+rWMY
D8fIMvtOUFCC6RJ+DEyyWIEJK5Bn5mVztPXkzFKcQV/Ck4yDDbk1Vg0ZjKny
0bhoXVNpaUqRCn8cWQT+XQIhU5Tvo1Ap46nGC5VkRHyWSoBCABRU3oQZPVsP
BWjMhwb+43EOKwu4LUd+XLKuhsnCPBtO8HS01sOBcHbMI+D1YE+7pL5c9ar7
6eowtS0fkP78gXMkNoFwFyTkMJoQQSPSAwipun2avMyoGlPf2D7XJ0lYCJhh
2tA/d72wekSesdnjZgA9m3ZJB+EDblJ5LeOTuRoaGp5WTIUbWafo4Ga59c54
LJRlHL5rztZQ6e6zdxA3AsnauPEeZaHwYCdA/JwXTU+8KQqAkf/YnyX0Z1DP
T1UDIAK+j7eaL5se5d98NPLNTNgnA0u9s4PJpZUN+PG8xQ0Zn7XaEgl0SuWF
dAd3bSqjM5dVCvL9tcmnTbIcRxlYPWbzVfTaPmdHH1oQjm6z4FyqE0ZXFlF3
GIgZUYD81KbstGoOaBG8zvGUqaAGGWKRVI0kZu09d6HLXIQU3PRPkuwN++HD
Of0mplciYRZXQ4Y7ie9dEtWMMS28RZCcbnCGKwmnykeUiZ/iCYndta9nx/eH
zYgO89dpUsrRi3Ppdd9s0xpwIOfObzGwKaFHOAj14DfzdmADDwnwlXVuwN/N
Cjz82TFqiRNbFUDJ6YILpE+29GD+gZ+Puzw6Ek47hrq+aqvcBLsjkrNYxYqC
y5zUHkljn2XgI42wjejxEwBDwmb5rIQqkzhCJAs6lkLYMv0jtiQP4fjBZuXW
hFHIuYmbh3tvV72w/oMxJZDpb+s4LyzX5BQDNCn0UfCw8gtmIK6WrcoBa1Lm
P+Z4ErkqQFlEJIMn6Vv/IJ1JAladDYtottI3g7g3/0kGqKhDu7o9hm5d86RB
gjsutjogm1txHa0B0hhTljQx/tpkbaWQWjAA4u55N9EtTjoKjpr+FKUu7DNt
SK/615x6v0HXo6nz0dps03ZS0ItS0HwjZ3DrJUOYchW8r3Y/60qOIyG+5Hhc
ja4YOUOCjjagJbwIASGGpRQC4cH8O93Qtb6ENM1DHag6OZPhepmc7exSa3yM
BV1YwuXL8Qx/6rBcfbQ9YSeMD8cbJ3a3MufIAbWpY1lxACja+DqwiV1bc/IY
7ZXpsgimwPcz+vy+yyOWLloh6GVpMbcQP9mV0NlkdYSed5PsZERUtT1mhLRn
Ho9L29Ie/Wi+XsU+csSEWdP4mgL6k19erLyXEng2F0mGF6j2uSTeo3euw2Rn
kBxx5rpmszhnhfs5ioZAaCM0gft+vI42RhlaVsWHlQe+yLrHO1783WEtgXsl
Vq44JcqaXxeBd5LPmbAAMX9g3sWBMjNySi4Uuu3jfA1VBdlaotRaRLdQw7hX
iWPnL4rqoqv8EUVegJmkgE1lodBoMApxGRyddouXQK0jsmbsUoLOmL23bm+9
NrFbOw6P/tpbvRFnYTe/RCp+4f6ntwRDwugh0Pqff1EryTUU5x5oH2zJLs13
G/ExJD1YsanYzIgB9vxHsKDUKX5o1hvv7w5Xwk4jXd0ajroaBI7j6LeeN7iw
v3XI3Uq4Y0oESZCeIBi5g8bsGn6mj7QP8Y+oP5P+NpSM+8NLxt6mK4VKr5Jp
MuEW52RdIDahDvVjk5gDg9fSDRsMy1P1MfsaFeNUwvy4EQp9HH9SX+LMasZX
WX2niLXzL2h+Tn8nwnF+XkoB//N9mwI7nnOhTWScA0fAGINHjEcoREu+cyeV
78xaLrg2nWJSAuEvipiFYPZUxSU6Wr/WJJVl12B+efTWFZPwnKlMnq7xm7nM
wY24ZTKVD8Kf2Vfn5rkSI++ODNfeed8/ASaXJUB/Ba4hSqpcCWebprhAn36P
J2yJCpqJQ5uRZPEYtqbvotkplUVcrgfk4O3NEHi1fUreWteBN3mqOTcpc+ZU
ldZmkIWfYqLaGxztc3eyiyPzHeehiiCRjEE7UCy0kZGgeGpDpMsb1ohtiS4o
I5PvWRglqjj0sgFTogqVGww8a9DFxqh4X1/87tFQ6QtFSJv7Q1B15xySS6hA
wtXDvWZIe0CmDCKpzpvEyXrkchSIURfKn7APL4wL3fP9FHTjwozbtszooh9g
8Lyc6CzbOw7+QeszbPuwI7qTB7axMHe1mLH9XcSx3lXyChn8v1LvCB6Dm8MA
A/IZ6klwfcCdHJ8iQ3SpH9ASfJQGkju9v4Ih19HX0htVETa8x6Dyn/EYepUq
feYRjePijUJG0Gw58xFgx0E9XQ/6YAPcSIMq5LZJdSd1J3doFQED5G9Ow1vl
uhxmLb44ymrHa1ErBO9gXGBFi6Em6EhuI1Y6XVC5pO2kQhRITRN7BewaYlu+
pdn+aNsZSwZCPtug1ja/rF0nkwHIv+UhVLvzypvFP4L/DmCE42ckQc7WBKZ8
hfDXt2nLC7LNocN9pP4j6qcLBB8xWPWKtwlfzHpkrDXbE70L9ZkpG53FmsSH
NENvTcsATWRxB81FZhKVMxfcPr8ZUIucy9fG7arhWJjZ5K4pjYvDfLFYkyZ1
fOo16wOsMNE92tPr0UfmYztRlCWaRj7UKh5mbCfDDsq64nHgiRqMUMmZMXSa
UpZkE3ORCJkwrYu4kxErvtmggTYYZMr/huhA91OlHcuMIMu92uS8CJWQI4XI
xVbxoB1pZ1zzqGObX6+ape9nSHPsWiVzmrhBKlbQ89NtnStgGczi/6V3My72
F1sh8tVAqvakKPHPFrYGFn7XHZFFohTcs77VqnmOJGRW9WDQBb0Amek4oWt7
utVI9WmfQoWsnt3PD7eCw6NSfcI1zIbAQqZmK8IR15J8Gl+dfxMdvy6/iStf
BsCxY6DvR8+duuYPFqGwWgiBHQzeKrRqVO9tWutbh9oNb7p7k3IZm094RzXL
Zd7R2ME6k1ddUNAfWDDImhsWqvoosShtYYVE4mmDqEFdCnHXOlck4AJfCMg4
1bzI88u2ho1M00faSpidg14UkE/SdEwYiV+vwJh2zQLbTIcwbDxpyuKvOL1O
SEk6JMMYxHAL7cG5Wa1W8AJ+aUu3Zv+ZM5t+oQNwcbxjgeIGlmwM0TGYAcPv
80pl7SmyFF2+EhHnoeXVaA9cQTr5X7fLD34gJ03MfKfgdW/7yNU3Nkfr30cC
i22S3D0YM38a38VsDUeioYuRQ629gQmTk/zF/nX95gYPe7SSBOCZzHNJ+L0f
ydjTJrsrFjfQTdlCzi4c2L+hERKMqLQpOR2mgPNAZgVmM0wHrRnUAASvNUxB
uP8z/2wRSboNN4esE/NnNHsW0+AgcttHjVQWPBE1x2oLEZrrxBhO2FnMwuR9
TGh3ssX0loMjLNmv4CLiCVPDULJC1TTZ15f4EsGs9ct78xkMFcTRFk5YhIuC
lb70pMJP4iUuEbqh9egXSP4OdlJhqodCj6DQvGGTbEmcejS+x7xuljIoEWd6
tAFsbyo4JZdBwVGYrkblq0I9CcYWUro4PH9rWZUd2/8fZgRq3snILmjUIC4O
40LvIntrnVioQ3YcyKzmiOIIMuCBSAkatVmv5sCi0NM85sNoG9UVABEqrWyf
xeYOmT4qwDPNDGn8N0S1PvIUjC3KyejHYkboJ1uu1btn1XBGiK2LCGCr2E0g
I1HK73AMfHmJJQMcn6Cs7j6cnwNUXFpjYnBeNGumEbK6q+XYxIPgOFbSrrEH
BvztAP78G/s6ti8OH9MznpJMdo9lxvw9BEHxzMSk7Z5oUiaG7jPha0eTZK2o
RhPmv+WNMYaQDg91xWOhf3MsKPtE6nO/xZtlqGOBdWxLyRLBBFqyicyHtHGa
j+vVx8hLfCRLzSlTEkn4KanXcfdNsfCy7RCF4+eo/9qU6fPnxAwiU1vJmlOL
exRy71uISueF8URwyesQaaf04S+j13HP9YnBw9HdrbPbEUdOjriw/0KHLWPj
hhRkx1ef+E3Gjl6DeiTGSptQbW3LkVpXyUQD1G6Mk36CmE0ZqrR4MS0BhCb9
B/O6ZuxYvSxniEJofGtIjpktxW9rshEz4rX8Ju3C8rnruEFxWkiqLzmZyD+S
jxPky1LhaXJ4rCdFqWyo9KNEkML8P0RPoX9+2QSsduRIuXRmH4+yEs2X+ZOC
J1z1mI3B5JRiqm551ZPfueSAl4MrvW5r1gy413+n+/UhprumXpUF2y6Bq25F
2lO08P49XHjtjM4QrpbP2HvIQrdVc6H6ME3/zm61loBQkGswUvkJE/SovNHh
AdZYlONQT5OwLfGXj5lu4pDRvbOGO0Z1fSSHRkJMSwmcATKjJ9JulAp4ZOz5
dJjb1HuCJfLbAE/g3b805DWKCEg9Krbbk2NyeDE4WSWrvBs4iPOHLP7YT6Cp
xf1PK1/9W2E5yGiAWFoXcmfRaIFib1rkyRX+5M9G7gP+VJoLTaQYn+jW6Cfp
WHr0+ypsUY2IFs/rFn/wzyRuw/MF1xkbKOeEFNqU794CFM5p02nI/SdxMmuN
1QfQ+KNWlLKfwQEVTU9KTtYGqb7oPzUp06xUARAz5+iGlppeysiqnsAUpSIy
0/g9P+MAem/tCni8II7BrgXqP8pizdSBF9vPUFK37BIusHGof+ajd32ZekSN
NGytJVBKiEkHdsa47TQ5HJPRh8NTm22lE8UtpmUYWUMOOqv3DhITBocn0Bly
Sxm+WU5r71OhojoKFFz5iKGMfk2LbEohFTPn24MPaGSuJx5kHjc0/sWzHOr9
OKeAYXjWWRyYI2vkXmbHn2BDCUcuI+F0gexcE6CpORiVQPxnw/MJQ8HvvINi
fc/41U+Qsi/11Oc2G2ITJUT8K3PGO67cUF/ILr0HCFzlIll1LDF7a/leHGUo
iHxYLQMJZDpqKpQ5fnxugPhD0Q3qQAxpDt9lB4sbwX1X+8p9PZvZ5O9glkin
vMEIWkvrRmggtfH+mJpxwxqYfLeaf+N/HK6PUZeCj+tSSMWn3znyhccQYKhg
6r+ceGUJurlvRgCwusM7VgdDkFNHmq1JP1p5KTEmCAqtnrgPXOKT02cnoYji
HpT5AmkW5Nim+eATQzXNtYP2UMOTHKmoQG/IoVDDvWoq2kx58KnOejHM8xoN
EIPyQGftF9e14oU/jOuJruFKXxzcB5sDb/Y0O8LzJKGFKVpeZUf0N1h+qlSJ
ikIvLWIaZxCREeyxJh+G5Zda9t54KJwaBuycmPoiZ9yGTytXlVwxsCO6HFl1
M/Pp9FwebsK3NRCxwuyXijhqS7YmnL10iIQa5SuXXLbI1y+xjDwEnkxGu472
g2we7HOxNxPJXlzzSWSr4edH74ex/uQ7hf2LR9G/bH6Ifdqd1/pYLmROPOBO
jZy7b1H6tV8WeGDVP6iIAzpkYIFHan2WvGWHUUmpFEEpbbo4YurvAI/esNcN
7P4wZbc57bXkvTK/T5f0rJmmpgsFiHki4d35KBnZIH970Y4+dJU1ez7HG5sJ
PvoUzRNArP92gItrTBlWUB0OMz3CB2pe4wgW3rjc4kLujvCVw8O2/6P1A38g
9lCWpGAUAmU+vT7ZPGilEwlmJD7IsvwpOo5XQKkV212TWQ/W0VZ6NhryRhbr
MAI4DDEcz+t24JW/m8ifX8bJLXlpRaAWvhsODE6X95kvt8aptbMDi9NaE399
2KZzV6W4OX3DFpmUkWBRXDZmX9pdZy8monsBjHPcyC9Ii+ia2lEqqVh2hcbT
U6aD42MLjTi4A8fRQ8vLvEp8juPe05Hb+O02TftlOM4OE0PbRu3FHJJSWuTp
lNhrAMSInjvofEyu5S+i22vVZopT2U2gffl4JF4pi9Par2acLJcpxYBrp+fQ
WzHpVcGzpbyw1FM5uar8O9IVQxcIlzlKsBWB6BQqJxKKnWFna8sRYFiJu3Nn
Je5pHQH2Kuslq3L6wIz6IGZ0TJFrdB9pUwIeyTx5aj88986DKW1rta+uOHlD
GQG5fQmRi9kbv/NlbuVb9d+BGGKrbtHdEQvUY4vMnA7gZHXiMJXGPkvLeli2
9Cgg1euIg15EqCLftiazFnPxeC+sDaz3a4bTlGvYp6Qh7ccc1aDEsViovkcS
ssjACdbr7OsLzfed6V9rznRd6RV0HfKyW2dkzITA6baVFBFrCogVHqkMVV8v
ccC7mYNQRfHXzawSSPianptRvfYScSh0Gc1ahg/T0QoDYjXFCqB51P1BCTC1
x70lWbBCce2OIs+H89zjyFucmiDtxmO8boE3NA5yLFKIxEcuEClH4bBeDK7f
yJ/vwZR+WeavjNvikI9WmOkqT/OB0SH6SHXHvj0aoKVYkc+EoGXdmHRuH13X
ek7LteHAanxNH73fnrIfrw3VV2xA+L1460L7KUwu5A16dmEfpmN1gEEA2mzp
/tXpsApGNOVxgoYIEhPAvtjN14p4eWima7IIykdhm6sbVRVuun88LFMWAnZb
J+dXk0nptPZMkfilBiLC/l1b+IyW5rUZqd83kMwTzqWeOU/bwOWKx/QxpOS0
j9QbK4o3fEJPtd6JUg4wCcNYqIhZcnquA98PHH+L+EoJOC2touZKO4Ij/5qP
1idfrhrZ81Aw9GjUvjFfkL8apKkEbBP5GcG+bgA5VXbrjSAM+vP1Ztwc3fb8
CrgH1gXR4NJMNEK+aDcpnaa73izogW4LwKLyOpQ2vd6HYvuVMRAX4OD8nyiW
MUJC4FAX/+KPvuDQR6Vn1tOkKBIxGsMG00kOFXcsMYMy+c2VDq8XID13A+e/
pRHebOEBA3a3CzxQORJMTr6xA5I6203iAVFT2eCbwrO+1xdOR4zg30w6un9n
vJA4RTvsfzkH3iAFGxikinzLUS3Rlv141CSHOOUpXSyIV9c+FL31cpWfpX3R
ECSVScb6N+zv1Dc6T+6NrOn+FROUZR2CAiR/f+vbr/k5Q9Dq85ypNYBfBgAk
G5vpE+mz4caNPXVJwAw2TCE47W6Iby8EEIA879I5970jnEHto5EJN8mG7BFJ
cHkXYDd9HWZ9fdyitUyPykUz1aM3nc1ZYpqgpHIhMk1ZUgdENOiCnumm3gso
I/js2Xinaw6DOR5tD4dRoHxDUHQLPZY3r0meh9cyg3GvPvrE4G+5TmomR0K3
ASDX3ogNAZGfihyV64xy65uwq69KfimsRvmUx4go1zgs8rXniNuDrtFFbJuA
1Qj4zXwy7n9gHWI4Cqf185v3Fj0/xT5f/Dq/kOM8Iaaqkeste9i9/SL9YwoI
GJG5Ml1OtsHcr6Qh4P1kb2vsQkwWRY8KN2d34aFy/SXRfKDiljRuxmusDK4C
CeRc1NmMtCxyX7Baxt5RzvGfoGisqJHUAtdaJ57AZqukitLk7IjOyjokGc52
CIM13ZOBrTjn1elIWX1ffC6XjnwbBHIUcNEO3dDObE0NVo0sk3JemD828/bH
7WCe5ympyH73QC3lnZWXTeC/lROTeY61mwxFvwui5/ttXVEeEeA/alw6TMOg
Lto82jy1JwxNaV69c38Oc2hOKpM9oVSxf9/790PAWwEEvmu6lJ2+RdA4gKZe
KGRPQhVtovkoN9qwCjgYW6O49lIwks/dyY74a7hFiQP5zVcwLKBPiuseU46j
AC04IWIJatgt5qBKiGxZVnBB/Cb1P86Ky1auQyLliwWDZzA3OBAtkn1/h7PM
QVjrWPlpOn3Hhw94DQyRdzLlUrY3Q1UWb2C2uDgFMl704fudqfEOYNShtZTi
RYkuy1JJzloFmx3bNrb3X7H6VFzWCh3qM7l08Pg1bIyRzV9NeIZ8xxQRm8LS
msP1Wn5xsK1uAEJLQGI79EdpjQn+CyzKqkfZnm/YL08eOrVDoFgnt3Pw2gGW
gyJ2yWXupDDaaBAy5LerIkcmO7nj5LbLTg07sEILTRItvzev56eGqPOkEEOo
w7R2CnsveJfjKzpzjvnIT6qF6YMQrXQ9jLfuSB42S+uqrzdNvqdv2jAchbJ6
Lr4f/CMr3SXwB33wa6pgyEzxUkmh/SzsTSAliHXGtOnv9ijY+xEo+QyaY3xu
ZczVq5N9GcVZVetvRL0CBoVdpigAsJFyPJKEbqHZoC+APcF+yH3XG0EcGc3b
mfnT7q2k/21f9bFh39dm2A4FRyo9yLG3L8WDcz08cZCiEFQKL5OCNbf6eRWs
FAAOTw5lsUZbcVjbI5cCPSfpEc6v4BaVXavaKzz9QC0z5JMDeQPYZ5NMr4VD
SinHXxbRuyivRg70kZJxyQZQqIuQlu0juF/uz4hGm5u1aS3ShcgAuLL1B4Sn
Z5d0PdyxMcCMsQgqQX+kZU2S+VHUjPHxZYRPypIe3d0cZ6rFRMrNBpfLft6d
0AiEEd6cAU3jhV2vO6ApIB+1GNFERSUKhlzFaL40YqtFQDmOOK8K3jzM/SIi
kwou74y6pt3ZhPaE0/KO8lk3VUHyCCIqdWrgY3SL5FXMJWgqF16SAnzuLvPs
Cebh36H09MprtwCTc5P0nuYzYJ0AmK6JMQk/VkSL6Su/hmnVa7JDgdRWM7bd
j80wv4+9zzgrv9w4As5ksulV+5aad+Gcr1tPwvoaDjLSKhebViEHrz1m1Jhi
GyFlp/82ck5tEkbborYaqxeX/xIx6rq+j6lG8QwoM4YxXhQpAl1ABsotXeBG
IDaEnP6rofdPd2nZIM/8Z7tk1Ah4aPZefmrOT8fZRyUVvsqFLAUzfh4EzTvB
tQGS11nH32zyUm4WTBfcxMgW3RV0+Sc9+zoyZ0TsWupUj+31kl7fnUG/Yx69
qZJf9Hzt8Wz6tGlRaOQn2PZ3nTAj5iOC9gB3qdzGmMT85miBFXBe7aFlrdne
OIffcw9WVmJEMJFt2+gxFd85I98Wc8K7noMVEPMs2KomUc57L2XuzA2cKmiw
0Ae8DTfM/kLDs/HSG69kjWbo6puZrihosWto7FhUQcwOySOpPVRcDOPKzKHU
Db4pZR7Ee8Hnds5URvoandk3LkJkMboe17FskbgqGqlRC1D9C+TL2VM6LeJi
WE68deh4AOp6kBI2GCJroxe6qM6phSLVCnPPdTYBlyauxAd+6ur+AKVWyWC0
0SUb4uLYF096wjbWm6yWsB3BtBLd9s/uQyBkM3/JAyTAkkQtA4rVyaLJKZe7
X1tlr/ZuXPiRMlClQ74zo+FqJ8sl0WcY2xOBNraLAQclQMGb8fHX6TfaQVuY
X/FNcGEHEq3+TxIXLSwOLUQkjflJgvaR6DGu1gM0IqYxvJzWntH0PqQProRn
p6IsZ4+LjYwIRGkTZ60Qq0yvR0UP+ALOUxBd545MEPEOhFN6hMGgdvaFFfQ2
o3M/wS2lNDohlz1vlTpG73mda0bUyBjymcKlvPeXvBQiABaQjIkyN1odn6v1
m1GlpapzjneHK/vIgNXZYQ7lLLnBbM5z4A5rg+RphCXKglfhFqd5m0pMm0iQ
hVdrepcVAOXp7nAI5xdJSdTAdj9+dKyYO/Ochz6TERC68+k2ECJ2NdBU/6oT
fTIWcVo9egSviX3Xk5SiCrGjFbWTfTgssedoP/ingsoh2F0UYRtMpeyHNtTx
7oVOgF94tKBD/mVkQHp/KKy1dXLh5RJfzPGyYR3pwxTuuiq7RHLo14+yFJ4f
GRW+UZw9VgXIEiF3Ip/NL6zALzdnqZAUg80NhdnWkND1P8oepmAVH1y9JEI6
EaqARoT/cGUlASSxyzJQqOhQ/HjGpYCbgU3K3wY6qGrQE++d0debKbeDuRl7
1khjanwcC9C+6vjCJr8gMresviRvUwqhPS88Tz+mhKZz+tZni/oYEI/Vq82L
sUPIMkgDeiD7d9mXNSfwdL+otxX1NslXYTdU07MVEhXMBexj4QMIBwBeADdb
kpl1nikxIjDeJv1ymBINyV/5Gqn253UEVBg12SnkpR3JM6qVKIh7dbZw+1T3
1KkxBVx+HhIgBTVwkWtX02Q7RGlaOYx7tr9EWMnGYLzvwSXP4HTjQNplsEst
QcgN1YM/7gmEO/0HIt5i0kdxUH7OrgLW9Afs0xm2SaX68QBiYPIUvn2SOaYb
0hSBhyY64OfYgYkeqbYm6JUQihK9cdN5EpwreJpmgsJNVTfFIQ9mqvUHzAUj
jGLwyigItSyGC8SlQJzwrejO6xn64sA81pMwmMQnxHaHuJ1qVaQgkdQdGxWx
C+hioGlqobjZSZfFCh/4V5JVgiDtkJX72WOsWLVN1SxRFTgsM0N5yv1PYleQ
mwGuptqiA5is8EYua4CHGxKrHfPQczXxPD9GB837zmYM1WlQ9XefrQtvj4mC
dNWZuz/wWXqza0pUjgOnqDttN8VkglzQ7ohqgnR/mCSULDixsCy6y0HTaoRq
US7jJ/GA0cFcpFHwICBttm2sYsdb2pk5SV+gb/+H90+d51LPmih8hyJ5CU8m
UPGdOFfBubC5CAmQR/JLs+RQSDrQdUXfGXL8ZRNR1BCNkneE7ikUT4vBRIV0
VObJflSdXWaw5+SmDKa8hphb4/3Mg7L6pRXbUd+Ht6ovPaWtSQNz+8df45GW
Ixc7Cv8B93iUfrCkbNklsGcrpNGNV80+NdeiByIUxXOkdB50vlYdVyFOb8Ds
Ub0LWa0/5Z+hjgf9uSBnK3yywGPejwiiPDCBVbBTyTR3e3lp0dU3t3ZJzSsQ
R/+DRu5l2VoEztuKGeNXORov6o2gx/cWY1TiHb3vibmSkrd1aA0QZ59LyPi0
ht537cc9YHHUTz1tDicamzx9gdsPSOiy/dfOXgia/Q5ow/ZJ1hIJlFKQphqB
Ge6EOh5ogZ0JIdhf9deGQZU7tZn5zCxpYORc3EpCymiZURl9GxQQmAVGijk1
IWdtByk2tQFiv+sqiozemUaQuyLEgEpSiTFzRocvDNvujt0HE+Lkr+gopDAU
YyIfEP1do1dfi7TbgBOCwd+kHX+rlDyillAb49p7k7q2V2dC9XzlU4UuntR/
KWD9Yv5j/0QFL8P6CRL5L4bLH2irraJejBupX2loIUurVHQY5jhSTXbO7kaa
CIQz2z/K1syONoczWcEN1t17sr+LzANXRqvZGhI6o9L6mTJQKSMfuAC1E0KD
j1P3AXp6xaT9m7V+eVE0vh8Wwr80bhuYJHtqctErclg3/9VYnmIm64v3X30U
taX8R2zR3bLR6apiaPiMZy8rBAUcFgGmoAmEecmq+Gpe6wRBtf7yPkRASDie
SWdQnTsi4yqOLaiKG+x3q5V9eMIewP5tV9fAlHUrx76yz8x0IN4t7fa63wDv
77ogHvLGwju303U7y7k+BofxTxUtWZNjMngefFJphA3oa3X5FdoA+bJdFVOS
dhmSILrarwFu/tQm9Qb+dXjaew3c6z8eZSI15OPowgAq/+ZKzRFF7k9PbfoP
t/X8dVAhRJPNh709gg5NB+jk8JWivyUvnnlUK8e5/ezHiwyro6gUTVIJHPYq
6RJjTXUkIUuOtIIHKBlUzZkrZAd5D6Cg+Rzvci1a1Nyh2OrQK8kckxNxI4Wa
nfsa5ETGytvpDB41umladUnWjtpUzrZ+duFN0cYPNdfeCjhxan2lpINDbEZz
IUyDLts6BsK3jRC+opIS9zBS8rsfmOi4EnsFx+Mr2URhDR7U+aZa2TNfmF+g
rzp7X1CfObYLwCp6oYyF8m104MfFxqHuYP13qL6w6E2/7BHiSNEXMNFfKDtC
heAFJmvljqvoRbvwxy0WLtVekJ+16ZEHaWjel7yDVVOEHKC/RPx2VHR4HFG6
k3ibh/M9GnKLtpPIc8q6ImdV7BNP74rG5086KjsBec17GCp0szKgtwr01x5C
wk50oKgX2fm2pTLIz1kJKcQzsGZ00RdpWgZhtLo+J/+w83JxU9E83VydyR37
ett2caoFNbZ/sBGAwePR7JV0Uuj6SUrU6xaEnQJiJoPqoMkOC3cXHQpUl2C1
0eC8HuoXqx5ZTA4nbapIcmZQpAkJsm47H7rcicsdRervriEdwLnx9TM/g05y
Y0Ay/C59IogvsjbEL128UBVTCFRkPD1STRpntRqGKk0ZonI1OgQ4+ThXSF5P
0hnEW63vAyAdL/ULL3VjMPunu3U7jkcuVgNcWd0EoE3N11za1bt9pV4uCA3E
HAPfRz65oXKP9hdH7aZthu4VFGeMk7Tsg3hp5rpxDW2shD7m6w84GsQtmVt5
f9YkieE1vDwWogpx8gjavCi2b6xqQVRpwxijWM5rfUqluRdQh/fP1NrwtMUy
1mFtnE3rd9eP85He1INk7tcWzdZ96FBBQEuX+llqN3v3ydsy7rMHLxZ6enWK
LhP2LE5sb/6pJH84M42cQE2/dnUW1z9dFXcQDv2qxdF+HCw8KoctbosUlgvE
h8BqrWSYMgelt5X+nGwKVIcpFX+2cLWxPn0A6PUDhMF266M8/y0O0EjC4Kzn
KJTD918SOBQA2b1lqH3bsaQdZ/eUm5NkzThGK801EvMsMmkODWa1iy8ds5H9
+HuRIaKJb8KLTD5ZQWdci+8wuU8k5E3ZcEbavWxKa2Ox8BeP9ES4DA/kmoIP
xrqqToVbrglmUdATg+CUA8TCCj3zKAznF/Ie6/F0n/01bXOlyGUnyKTThvxv
SFmc/ooTBrrttD5AUWbacBnzxuKtlUCT88hTHHuOMFutmR5yP9MUSY9dFXkU
VcCOFetj05Cx3yyGPYPzFUKfomSpjhul9amVKbak72DZkzR8cqzuA5uATRAP
ztAZCQ/bZkVFOCjO9HmUz+x1qMMsVQo4N6vqq/w4VRwAkOIlC8/FcK5ZINV2
6XbHY5LSxBfLIjs3Rpa/uyQ1/VTZTioR3/RzNPb+slx9eZV+zDD2W5k6tN+S
nEaqw8QpiAsZHebxzfZGQ3eseG3R982R8OZ98elTqSVH62IEgeSDYwySx2Zj
TMfQ4mKPT7LnxpuBSP+shirAjBjgOLWrOQJorSYWkvyP5hzKU0vsHn4xakFY
ZUFDzwRxeQgwsmkspw5lNosFdPIxs0u0Z3zll5gHm04SOvCL8cPduQ8Cm0p8
lSshkEbxIa2exJieijSmcuI2rpCoZcTqIT0PmJFjuScJb5nxB9tAgP2yYfeZ
gfiM+lTFn6gsz3BciTxkA2dKKZHdgFN5N/1trAT/jaGsiGiwNNMOQZklG2Or
YqleC9s8pNR7UJRPeCYWAE7dkPghyG53t0hei0KuwBRNc7b1hn61BNozNgvt
6QAly4Bjau/j/qO3p4W085AP2WcAGaL8zxyEBU1Qouk+ku2amHTF9neFSiIA
KCkgjfOjTK+6h8GctlLkr7VZznALX8LVIHU3jVVXm2vROlarwMfPouP4D+3Q
brYz8tXHxKeqS8tFKLaRFeg8fmgGWoWS1HUEjac555fctShA1/hx8uOPOTdh
o5ufRPSnGR9EYpzveAEfyJa8CdsUwUaqhF00irvhUrYi7RXWx/ziMqxV8bYn
27QyKfgN5/BLlntRlGgMIC/Lc6cc8ubwkevCTWmD9l/N0tBYBfwFtD5uvPwK
RRxfmZ5iH0BX2ZOHtmzbCULpNcHb+59w1HH99VAtm/f7Y5NBPmi8fj8Eyp4M
snqaEojVfQnoNipgzEsEAMfrk+nz5CU996JuV5v/UejsouwqpvAUIpi5Fpir
Pw37MZG2L8SCoPQcFHvtosaq/XX5yhdeVVC8ixXYkSMOZTsAlYSyKjBFj4Bj
JhuN491Znwi9vLy0BBvDmWDw8Ff6cbC4wkVavpzWiw18S6uiuy+lw0IzEBjn
azrlGAmEUvPTCChYPDivNu5mZds3ibuuh0caOyEQYqOUnYCj03BpCN5jFium
8GvpuleXrS8uMue5Tm4f+5ldwJZMCgUvsRuo/fS3GIqwC7zamjOFpmE4c+RL
q7zrcdng4yRzlSakCBSjOUzYUEaZl9nAzy0Qc2fpgHHjuVvPiVgiei9aDFyw
e0Jz2YQASs0J2U/eQilp7bujFdDfrkQFHrD7J3UXj3z8xQA8tnekpRrT7YE9
7wPn5PEYgeoCI4NhW310j98UmbXZjha1VST/sNL31Ke0HR3/t83xzIu5J/9J
Xvt9txP+/1+pxjhmky5LL/tJo0a6t6/2etFp1x9tMIQkdtqYl0vlaJP/phwt
H/AH5fk76RWdlEpDxX8mZEfslK5s+V0afDYZHBAgrxmdgbNn+JB7XpGZAwli
pzlQJ+zJs/rfXrh2nKy/HWUiYyt00b/AE6MNFihrJltty/AWyfVTlhY2PM+x
X9ooLfigpUSmccNKYb+EHEhsdON0m2GaQAoe8386ctqrs/Q09ZoEDWbNXsPd
BpT4jE0GMe/n3C7MSLCPmUGDI7qnTdFZUjsdSbuEhG03VamGyOHFaysPnRWs
D0UJ53MvUhWoiLiKse6m+NTkgpTWtP2PLsA0HFMH3l58RTtqXQBjIbBTkIin
SCBbfSVZYipwKPHQggxj8caQ6ss3K7Chz5lPsMDW2SGPmj04+iieM8tZv3sE
yZDh1UgNFzyLipvYnZtskjQHUmPLzI8iQL18Jaeyn+95L3sBKycWpipkIwmU
/zN9XakuwjfTX/yKENKll26fG196vf+cIW8KjjWBOOMQP44E/4Q3mjTVX+vM
vlh2LzTDnXEu7A6qv5iWcNlC6eC9rtoELcfXath4rFj9hoHWuaRFGQ4j/IvF
U3vwQOJayLpeADkVOO17Ddiz0pYZhujTpJZ4scWWeeeu6a34ST3ZSWCOo3lr
fiROnjOq++QRDt+ctlwMUjQlscR/nzLmrm6nu23VW9KGXuwvkZOZ3o7DcB3b
5UKtl0TS2iOErW05uojR0QVz2bw+enLhM79L+prpwbV90EeY1hNlMIUlVfhh
m5SuHLa4x4MwXdY8l7h2QvpZtVmAnVtYlW9cKAL0angcpmXFS6WpTug7X8LB
66LMFPwS/zxtpUf6J/vrtDtIUPCFaXVphbXsRkAgOsWdqmbdaWSB2vEXZd6n
OR3rKdnz/RvQoNQa3z2DgC8vESMjXyoOxtBoX3VFlgK7V95917lelzEAJTJk
MCtso0l++DhDZ/t841wasxaANfRfWV4IuqJqvc2zUNSJLL/9qEuoOwUKjQfj
9+D03AsqgBQTDDz71ENuW5Xn1ZW588ETGvUR3n+R3E+EkbjO9r4VIHOIBDgz
dmoGO/hMq+83DVYZg9YRdElxsMf18WSDeZ94moIxaQ9yrdjEAIvWtTE/Xr4O
odqO4aOLg+nKqlpK37Nmdwie6r2RsSX8mMUCrb1mIGdcxfC0OcRyw+GmZ74a
wEgX+pIJ2krBETV+/39dwBCKG+f2EFoi1KObemeNF+bNC+sMUwI4acYcla2i
WCPX3SDM7cDfQDNgTfysKpEuWqahlWGe3ByWPfcBfnJuhQx8LpZDjmEAOxfv
zmZeGcG0S1Ulv+OC4GOcVZDfdwaFgmwXMu4SX0xJMMEYaAQRP3SOSvmPDfu5
lmwNP0wUuAVD42i9J5edeVuKmP3b0WWnDt+3i3azjj+sg92ON5EFqWAgccLP
0P/V1V6+RKGgfJOZt5x7j70aNBTER2unr8Dt4I2utlf43xiL/NXLpu2NzNmV
7ZswnlZk9xf3LiY17q75blUgq9MrUCp5Xum4aLBosST6qR7GwININETulsee
Pt+SJhJbF9Wb/L5km0We1UiWDhE/h7vkvEteounL6ZJWWh26zPXiHnF325we
oCY0W2JRgb+ZGuPY8SGxI7VcthZnh+c2OgraN3lngwiHGgzJsltO1PcE4WLV
yWz/dRsZu3khnO7pewlNp8yG88DaOY8IebYhITNKtzzw2GDCF0e0CZcRd6+q
obgRVjYdqUrAE12ztRkU5DK8IOYow0+Nzl0qjpBsCpGzn+6Mpic7MiMnhkjK
74R83AnnCI4Z2Hl3sI7s2zEFH9IVShqzFAZqKqglnqaa6O6bvu1DMMWBG1Li
ITPlTPhVXo1ds0ZpPARNxY9MjKEWq5jBwqo8aXKInq07ZBu5iSKlTzx945zn
97mcxII4HXYhftGv3o6yhjFtAlLDge7wnhwVaeAAPwioCJO69zsWpmKHEhDd
T+wgxa1jKk+2+VJkxDWQGGgvQLIcidVC9WgzoFuqp4TMe9Ww3X+NjhqfK+qG
c9NYs0jM5pRG9BasmZoKncwtTNQwI0FwS62DdTL1079FP7sK3KAKc6NUwquD
AtxB0qye/OaJ6FgesRm+BDkhFzspPLGvVnzexW3ITNWNcyhhshML/oRG0uqU
hmve9m0WsxrxGWkXWyHCoK9gByF7ow1Oi5QsYeiVTuU+4XwHHyLNhvK8iKNi
pDY+4T08pKQogiob59EkSeKRKubLKkbQ0fJx8fxFQb5ZHmkMCySVz9BrPmpg
QXB3sHVqgzaPgKN7Quwiho+ZnzXnWv78BBaJ1/osy+Gy6MBqpncHJhD6x9ZN
WwonMv5YtB0o/WNh/lkBKXK2v0H9+iPSEeKk5pV8KkSxH/Vp8EyjZX177AQ5
fyrorFOfFcmXF4EFqmmXsXjS5bzEBkzdGhlMoJYAg/FTzZgnnYtEPhZJSjo7
RtxBVaCgfDnyyw5z18bWHxR/0Ts+sztPVUnYfbQjpLjbWu3i71I6k4ZFZqYN
b9iJ/Kc3FixxoahQb/J4fQRIz5sWNxiXMvRfbT75+pAfzoRuEG1SGWWAT+Bs
tiNiJlnuSVVco6kr96ShSpd+nOFsF9D5weNzqH3Tr563nNmnHjiirNoS90O0
FQulOqnZrdZyxGiuTD2w1oRT5CQTcUUdZjhY5ZDZOhDPeLlenIV3jRwypmGG
JSeB/K5hdSLiIDu5DAXuIbBmIdxoS4APo6oXB1FpRNfS6O85LiVGvNlotO80
syCaPVLYQ5ZvUfECn69i/tUa5VelyLdLl179gyhdEhcD+yd6aYRgsQ6jqcb1
ndiXozANtQdTS2S0pmcyxdGXEWzU3VerPu2DecfdhHWbf/EOCvIZPJqedc3J
gSEpEQoedxYwSWXHwPPl/SaSMLqulz9znECqhytUjKqdM9FAuKzJjpbPHD1C
bayd6xaQLWyIBSxCyXADnKyrc8VDGq8vSFFSb1eFP6VuH+UhqXDOMODpg2mt
Vt+DQALPFywdO5zIWjczfI2IMIqqetOaEB7oZIR+btzt1uwCdpG08TB2Ilnf
f/oDwaBmwpORurhQV474QmRsZDx641e2w+3Ao2vJLZ+u8KegogPLpA7a/Hid
If71NCW3EGYvTLox5ZlOYTCXNNTsvK4g++fzE/afOvxOt7qeaBSNVL+0OMJ1
E2XGGELiKB6qarX6fejKlnjAYaUZIWkHEIPg7xtQ0acKTFlwT5OV0zIMGEZD
fsm8tsULH22JLf2x595hy6UZF+Ri2JypKyzqYfMRWyACM0i/ndWhYtxiOKla
jcx7KNt8rVN3cWBFJi+v4RAOmxLC4NSFbEyJQOeSqqxVr9R1Y+S9aymQZ1GW
v8qO5YitzMLKV+l9/R1yQmi011HM3wuZ1Z51+2Odq/fsANmd2OeRLzaZQOHm
On3OnjAQumZtIa3ICdKwWFNJHtTPyadH1zPHKmMYuJ4sYA/bsXzu8AgbDD1O
yilq4CFrhrdhQgUJipuUGMNS8YyXfZoRoILmh5zamfuXxvwQC+JSGQTW9h1m
gotXvakgM6p4YznmDOke3859EMX1Tv76ec46RbqSoK1p+h4JVW1C1VicTp6u
jDz99ddy9mDrLsCkASczECWrTUvIF4zkE5o9anpQg9rGqyrRmsEA606Kwxmm
63aSZVi5O3jv8pyPfAqY9IvlEqcn0h9Mu9748cVHP+x1xBwAyTVNU13ZVTZ6
fE/AxsVGVaqNHxu6QQZJEQ6Dz6cjDbqivEXBRkfb086J7htxJH9EgIP++VUa
iMgrThJX7i+9aRcjUEcaMNPFZI9TM2P+gLvyoDfiot16b0avoNDua63NQSMq
pO3VfgRTWYexGaXwE9PWbPoVM84v1eBJ+/yo2KvkEO0yy49AzBqRzuOjvY/3
IQv3WRY4PYgc0y8DmrxtWghCJIBs+tZY42Er5Q2iWQ5aFAfmCBa5YoDBRaew
CvtTo5xfM6NztkatZUfKIqyVEEYnb2SSsq/V4ttByJ3jlBaWkWSJTCkd2pTi
xtXD7RUrBA06mrbVFhWHu0w3fiEIYdkLlR1JCRxqd+3ONTC1WBTA6uJOJKzy
j7Vi/XE8q3tLVKFWMUcTp2mQRCKa8iYxw1GlXZrl5/ASQZGW8aEpxiZejrW1
u2QnSSoiYB/4w0AskMEgbRc9PKP/xJbQwDXFR8+RWjLedOyGZthn13XZ8usQ
xtgQPkdbs7df+v5ZDT1USbMJN45EEB62KD8JqPplqNe/2nk4r82+cCxJyPdt
pYyvlv9ymORT2HzpePZLiQuOWg22TdJIvzc+YtRsV11YVwk7PGbEOqISvSYt
SxZ9MGt5szcTC+Fk8TXpnUzv8b6dRnnPBRAoc8R1J372BvCNBrQ0/rLMn4lW
bYBlxBAvandts2RmC1TgZOVUhSgJuPPeAwcB0TunROy13b54dD46MTQHzu1s
9QaQrNoELoGjEatRw45KY0vpHoSOe7GSfeJgyf5CFk101i6B5qo8L3YU7YEx
xd6mZ1D5i51hoK2xtSsVNuYx7lA6D6UV7qjRzKoFW56RtMxIcZ3U4eS4W1Po
3nOB2vxGr4zRpNU8/R2oZBNcB2ia6sZVgpQb9uz8aKKIrnJeQNzvWLh4vwCe
gAVvsndEzqq+fYI9WlWR8lBsD5OYG5Fh1+kfZHQmAwWcFTpR9g7ICCDPXMTj
+XNcvz6fn1mv+rJSULYI/KgHrwLCkBtiJfBshfk7gOr38bkSqky6HEt5EAcT
dAXkRnfOM5U/T0p4Z66EXe75EJ1289a1ufHSMlJA4zTKWXKh4NhbIWAZ6ppQ
1JwWSz2P7p83dMFzUsRaqzTqn2LtYxw8iARPau/7XwOHFqONjFhXWS6i/8I/
PrVTiXjsL2QgoGnSxa0U+IF5Ft6wV3TTCekKstx0sInBpnw7R0pO4uTsQJzS
AC4Ytc27cgnbXF7X0LDCvRyEC1oVse0kLLJXUnTaq2bCUAmwkJL5IWmBVne2
z6XGKFiLnT8aI2+E2iJ/Z1p3HtKOOV9E7Lw/wdnXFZyoRe2pAcH4lqyFR+Mc
/DIzs/zvFBkp+b8Yw/1dgST5+auUvItWhzb5td2sgyr7YL7iyR+XqUsBERgk
3+E0AteNkXFiwbRMde3J1sgT5CSyx/J5KVG03YH6paSD2lGC5An4jMV8rxMc
m0wjiAHfwZ3guGFpkC2ujluiR5YGalrnnjEwDtuzPBI54sLWr3kg7/fOW2cZ
DTyl/j67OzIYsCXX97ASmo9QfkIFgRZaAoRHNuvKtMSBAoMFr69zDiZX3rqI
QTT1tOke30OB/FncBsAveu69R6w2zeSzeQbIly610t1scBpU/L8wyOgZN6Q3
JK2zC1k6TfVoPtiXHXb+gUvbwp+k7yDTPowi6zGxFGhPw4lYuJXRBb7aEQfb
ypvjyWjQJGhvUK+D56wVUu16MJE8LrkUTUcdFtekJXaejp0+g09XrwdM2K6K
2P0u8pym2ye+aCPBkSI2giGMjPPUrGm6LxDT17dVnjrw+yciE/dgpcvsUcWn
6qs2gtmI9mimMnoOPQmDtFNK1fGrGYZDGDCDNMCbU7/yMSiY1drZI8Tua2fb
ManFAZqQWU7gU1cym43xaDrNAzPh7J7bsTR+8jDLcG0T2eTe5iM7Hni+tiS8
rFyfDXO0TqK8qbjKYywChDe9Zs9fE3T4d10xu2yEGvps48qb39OpnJjEtUMM
oivQIhX0rjkQWQ8MC687w1cnaZ1mG7RJ9CfY50Fxy8lWikAftA2cicFH7itj
8+KLpnOhE7lN/2mA94oWfXPyHz8R3PFQHWGSwFaRPxEMIvf4ntYiIySHg4ue
Q5oWuu6UPveFbiHNBIDw+tZrfBd8CQEiGLS7oT7daeMWrhng0ubJNgPpMHoB
Jojvr8Qp545ma1gOvHFGtQa5cV0EVbfumoJkhOfqadRKITJaMwXt5YSyGwWE
EFADDgo0Hm0FQWBkbP40cCDUnrQDalZSyy4Jh5lvticgZKrjDpfZdwKJwVZ3
QVjEKPsKOWWH78lDaDYshLEJOCCvHf1ayKw/OSzZrUU8VEL6Gq8rcvac4kMp
nfvlnp/eHIOJS0QsqxXNG1n+vPxIoMRanGfb6UeTp8yRPRdON9WxnJusVqnr
+jfyET8ISyM2fh62sZaoOo8h95uMLsLn02NTdI5BOMxrtdUgO6ilSpgKRY37
DNi13t/tfdJ2sF0J8P+6EX27nxea1NGgbpA3nb0K4J1A/bnB10a6OT760wPF
nvmOFrxoH6kFU9HTqhJEVXUcD7pByQQVikHWIHc8Z9LZK70bzluxQZE07g32
omI3FC/6balqxj2dpYS1odz59+kzOa5W5YCoYDzZIw0Rk1XIzIHI8QLdG9C5
ZpARbeo0m9I2mrYruXJqs1OsEV34CtiBYmVJTUSRaNrggZnnrV3JYzuwHSmK
/cYgb7Nudqk/4BVWYGmA9BYP1Rf3TpUt1bKmXWh9dYzaOSCBJv4kYwOCcNW0
U5qDf4k0OeYPYBS3dYY1cuNwYpVYAOrHU1Q0DX5MTDOg+SsI8TTQmdh66SLY
TdMIKYd1G7qOlUtEjpaICqh6Cmh/H3gBls8Xhfykct5Sf/wkS/m7GmNPcVET
KKGaQ5wupF2t1mjjec+XHc9p5TW4FlhZFB6huAWd+xyUkRI/+6AHezHHQ9N/
07TgIe5b31ECHxe2NEUOaVJ1eTaXVG2K9L/wgVV6zjf2NDQbWlFsZ7pnwZ6k
wYnoFxaOPf5OEnMPKt/eGNScScY9Ps1BIRSoJuWZpDQ9PhkGy9coq0JxSUDu
jubA4jkthw3pjcK/wFpnhmkghYSyklLfdD8PCspidckugt0pi+zKhA9SHwAN
8x4mWU8iTNdoIM85BOfhDREbQ5p/1oGWLPpW5n9acdK7IGr8TRNR/sa60rE0
BK63wLuPbDpWWRap4kjPSmEXfUb0WW8//gHekhjEiNtDDGajvmlW9M1Gkivz
EFkRR6qB4r3C/yjBx/tRLKOfeLFXJlAXOsxtQQMGdo4hdqb83zEl2x7xXfSa
f07TCcedh1QPP4rxMUoHF+5Y4mCKZsbTBnWHn7QN7dkOh20AZarOmIbjsCS/
yxqkC0qJUbiUY65QThu+4ZSHGkza1tBiQo0/S5vWzFouRtkzrG+6fgzZ6JSD
lBt031bzEhShQvrngFOI6xOfRh6q1afKOoR5j8Mel9rA0+M+3/Ka3Lb3Zvuy
wx3DkLhu1VEpTpyLH/UHCdKx9L1xiQXbIEMu4ZsdIQBcsUb1tZKukxvpu9H8
DUVxx73/aEU9M4LWXFB9aL1u5WEH7fwOE2nxhiOBnBJUc5iv11eWdhUwD/dm
9UwPCzR0pgWcn+s8FKVbkXs4OUBkS22iddMb59gbsI01A3qjdwN66WbMWqqV
/oIdimS9sPngWXmfTdJ+LCyewU/Gi7aaZtDRYwFHZ6P1VlL9rstahq8PRPlZ
ckWBzFIMM3qoXxTGjHjkrPpbhheqpRjGWfw+6Kt0TVzUXaEAARrLhJxwpVq1
c7Xl8nLst2gTnWL8sAyVh3kycfbAPFmwJEBDrOI3oEoqzVDkUCQw/J+a4KoS
X9ICG363nbuXKLP9wSTV0jGAdKScHLBUh5WMbxkDzvPy+8uAxuxXgQz9fn4J
I3kEKhQD1eme9wAsms8ZMONHX32PdR97ST2LE19JkPFJH/lA4RUnSv8s37Pr
Ie0+4LhoXF/ZkOXfwIVPjG9ZpB91FS0nzzARCQu6RAesM3dWbCvJNn0fPlSA
8WISp0L9n9sTkfvfS0mgt0j/LyOmPqJ2bHN82cL80PER7/aIBG7qnebVbcGp
1In1xMG1EsW0+TLFUS5XrtG3Y3AtUlYsrMsMU/L2IpliEYBZkAsQz7Zfrf+Q
uWZTlWFVaNVlu/23BCm6Cqq4fuCJH7BP8UVdH2vMt93Ldc0pSg/fNHR8Rei0
9taRI/dDR/qqcjVGLufrCuluvGrTk4hHrak9FPn+nbYM8kkg6n8IgeYAoZHH
yurKN2BcPqa5FHBuYRp8nPBB/YL8XXmz3S9Rj09AcFfrDeSXwEOXFUDanqlj
a2tKwckfGFdHUYwm5PdD74WE+BLGfu7PqvP8S5f0blvbhV+D3Yhv2lKPQnRA
Kavsf1pfzKsCCEj7TF7WnJbDibhaPZZuwgkOwXcMW8OSyUwbKBJBBGSSH+nh
+F8sEpDHUl0Katp2nTawMG8U4UJ/fXgOEMN6n88k2jkhvkE6ilJ6d6tgs1zi
IIGj8UgRkjoHYz5X3nav1LwjMF+XTlB/pEBSoHI+dQDqhGY3V43JVio8rKrR
2yuc8xVVpI7Z0Gp36LFeexpfGO+vT25dIyGNFAFpzngK9dMcJpYMLg8ezJdy
14Rt6SmODYaY+ud+HLpR/x+DIUvCm1W6knC8j4FP8F+/aLmHkxsjD0+9rgVb
/9sgkYQchZiAdb1rTfkVbX5hiH5CfDLgBlZR4GbqE5Fz5e6BgaRDw+jnN9Qf
GJgVZ912X3T9Um4qI+m3W6IvIXZASKJ5LJr9DkOChJ3SmRMAvF7cYUIUXIs1
G4EMAT41Xnj8zpVYQhPAAxWasVLyYYphZQo6hkdR10NSJYIkuVsdD573MZv2
tSQs614WVl+VNsH67O65Lc7AjaFch30Bd77xwhKOtP/ha/NoKqn2TcoQ52gn
ysR94RcazwKI1il9So8wrPoOLEaFlreAotK3cti6inJ5Wke6K7exeduzjok+
ymuK9T5uRu1irTdvheDEEeq0tZkRo2bGC/yzuTzCQj3zKrsljLw1SrURuwBr
zf96/664uAQsbqursGrXsrsZ1LzCKmMz7SgQC9stCCMJmHfMHWoFhI3mYrjq
Oa4e7Jh/nrxREfWpA8Qk86oJLRh6pkvqcyMjnXR4RbdGSH5yaCX1f6XJTy4C
qMneCH3G1gQU4S4dWVrA5R4ypfKOs35fHRmq0L9LK+pGTGZJfKoEWuTs48qj
g1SlGN3pAjDCMyq7sh+XmwsFNFTdhg+jH5BlAQboMJUIiHiuKTHy9ZD9PBVB
w1c1/odpg8qz/x+0ZeuQOJ9f/AjLu+X6JX8vvzuXCRrAOatmZTT7wy5FFlFk
h2XAnJYOQqTPrIEovMohbZBsLUoEq8fVyHSg2fo5ccoYaM/V3YPRQ5PmaN4k
sBF4GGFGk7xMg0TatMCvRzRFsnpr3ZDKDMseXIaFSEiUuCd4xAlMK39WE02t
IVjBQI8KUmgNI3IQkaElSzmn4a+btKFUMgqbJFAh9gjVi/Qj5W9CovfTK6jG
kwYdjWWMPTqr8oCH7Iz6iarWH61WJhgNfEdQwJg9oyyNdDlD3AS/LMbCWGiY
rY7G3i4OXJsgqoWmb0dxRoKYyJemUt1rp4M4j4T5qottLwNFhf39/1MuuECe
Br8nL++fIU0R4O7PSDp6VQ2j8DQJvREcHUO2CO5ZUwQzE4GfCg0L7mqnMft/
exJnab6w/ShkGlNRpVjpP8rZB+slvS80mxkk6sQcUCKoielDBp09EqnMUk/p
w2sNHtB5BKM9ot1p14wny7+/mQI5Xs3txAKvolBbEbSjaozlDglkixicjSDG
XaZm0rzelTI4Cl4HcBf3WplbKlLNq8+DMK3mzFGtqzy6JNNBVTBsqsEjOvQH
Z+AhImQ8iXyB63zmyXF2WIpWsZbxW5GcQ1t3DhWI9wngBmdUijSTUfnGgkgR
YObGrt0jslCs9p0ZZwPwudElaevahnTaRkSHvUOB0QYSs5r3AS6G7wrYVTWN
PrPzfHynrFBuu7zhCa+TpSMWbFYCd+fNoEeVt3GjjTLA7K+41mI4ECDYreCo
DxKrbZtW7BDXvpNOORK/jlhlKsRZUIgt9EWRLkMF1JXvgttg/tUU3EVBz3f6
DcV4cV28I2NwZaFkgm0358ZRxSIKx2agxIWKlur+hf/sQK9+6d2jrRP7aMAY
vy9TOCUrsMLkuxTtQjqFz6nyO3lyZPp1i4ooELcWX8UzswcNpHp6ZMh+gEh+
lI37cqzm8PClS1bnTF+BE/WdxvK+ic2lKAq8Md+bruHrj3W8kG3P9mjW1xdO
5DzxSgiuRYtpSgiH5iR//HlHmtCDO/WO6IjU5WFdXMua1mTFUblkDQxQ6oYk
GIMP/UoEvRl9BrTkFdVysHECtTVOYTlShVKMnkKzUFP+lgG5sYUetiLOOcj7
gc5D+4ya8sjTwWQiB3+TOmlf+iPp7zIOqGr3khz7ii6zI+tGPw1AwcnwQzyF
zpEZAK/QkJxGCs6KOFl7oldWDodl95i6dq5+3fmjvV/vi2t2e23M/QFulVxh
fq39Wr1NK+/X1tjoYG6YpcS8O1a1+Q1Q/vg4jYYduzfd/u+nOT59vBGwfVLZ
wUZHEIMu83IkE9BoSua9aQwCRsMYSbe6v1nEWBe3CHSsH/Khsfl87P/I9XZx
o+Klj3cuWlL8fht++O1snkwP2dU1c/0SsjBKkkkGlNnYTAjnjrAjLqzNEKnT
1QVybWY/YeWvi++nzZGiLoKPrjnJ8yrFMO+6uj3018o8gWmZqxzH/YZH0gYI
tU1oGnV9oM8CMuTIJMbq0QMWiC5YSdAbLIaqQR2055Imq5uH3hIpgqGa7xXd
/L3BPqmMbamr4KiO6hi6Br7wH/+l6G2wQzkK2O1GDle2TQXwp21EM4BJmShf
CIjImAz7rDdOnCdk7cx/9BhR4igPqMZvS+MKUqtM6YdYMWggFKqIaHf4+b4V
5IK9x1liZFyrc/Pkgx5nIHimYZXXpwaC1kgtGivkxF9kVhvReCjt3fqS0SD1
U5ErKRbdpLrsd4s4qTLzLceZo9Pn3UXFBhqo5yENYXMmF/cD5YdUQBHrQjUK
lS+u0LPpfRSIWaYtwgWrGWM1z8axcIdQu5A+tCuwqK1RYGqX1PGykFnR53N7
wv8sAVX/G4D3DSxVuK01TaY45soLuGrC5aI6zpdIjGcwlJVyvG5syQ1H14Nr
LIx/x6MiPSFhynt8aux27erYdSVkNGZpVEyNjoouP+x2jO7Gackeql1/TSPt
6stJgddCNYT2Igli4Xn0RVo1LFD0WFNlLBXoF4h5wR1LbytUGvjnDqu3QBiz
lPxSYpI3/0i5Wi/+b4vDB60wKxmfnHlmihsTYyAsj+QLmj66K2dvE2dtL0yd
QJXrmy9k44O5v/EqJE9Lo6uNOv8ezot3idNUJEOA1HTNWfkTgy+1aiisGB0P
AYPiwmeiYuu+zRIP+X2xwl0jpAJhZ9c4Z1zOuKCXmBexFsrkUjj8Mt+dmQMq
azJZfNsutxi4j5GS8xsPuNw49Kz+9tRW56wJZOEcpMNKGdHayKciZjOPPCDC
Vzb9IuWTf9V8tizr/vjYdFKK8/Pya+mUkJ2spGN9yRk39lYyMqR8i0s2QXax
ScOBvJlRf9aVJAb0tJilG+x2BUBPP+J/20qilK62Oluu61Kvv92QC+UuERkB
lqM38pZgV9+gpXpzUClidYGPazQVqJBjR3xWWlUJS9Bl/+ylwb2sGGlnYZg7
e1vLILGbfIVlyDZz0xt7zs4vD+yqi/ojiGORBa5yO0uYDyKZtFN4aBxbIuV8
1z4NB92dfAXUc0S3XhoXGn3p1lzGzrRzHNbRbclRfCGt7Dg+hqsbrs3aoHUi
ZZBvcpOVwYNmHDV07biM/5FgO1DTC5Ua7LeUK5gRolS0WsSGIBYlQw9Nh3jH
nS8m3qFnRXE1vwRQ5su/cpd8Hjmavn0ShZo+5fo3QaECCUQgdymKxDRqRUoW
Epx5hLG0u9lCVZd7SJzDXkFMPCRk1nfeZzQhhNG5V5bUBfFdmS5wnTIf7GuU
ya+gXRfjsjI06YwleUYPTezxiap7PCHjDg34C2+BtuYRFUwsCJD5UUKsSsOr
NaZc8xq8/N2Jw9qqrWCple4l8obiyCZQmlIwmOvw9XcQPCC9bxcf3fDhBYgJ
q81lcTUWw7wk3+NJE9FxJO56xue7kEszjwwdvGUj7qZasQtIhnVENe3fffaW
qmgMmAoskzK2ZxlHD0ZZVEeV7JaPPE5UFD2l+QAziiMR5y9PAHe4DYHITZtR
5DpLnwJxopKSO+pdmgNRM+lnGCq0wzjdq+b+XP4BAOPMZnj2VKExEpmFeTZ2
gHNX/d3W9TLhPym1alLLmNEerkrZWjs0E569w7KR3VGp3AFS3WwUSrz4ix0F
uhWw4y1mjz+zhU1+vxTptwaMsCLCk05H14nDgaGvn4R6k9jQhi05mm0+2J/B
rsC/Do20phBAW5lKObZykRtNMpiDj9JuUEyQJTExoRrLmSxx4UzQqxwTbWgI
57fcT5LrH7UZxyzGsxj+CI/ah9PSFNvhtc882La7DikxnsRbQfpZilSXZWH4
rGQ55DP/Nm1C9Srk+ebuaLvloAA2OBCpNWICBSU3ZvU+iPKwuT34HU2NGcBX
ZsC9rqr+fEyWfD3nb5MXz/7+cthr1YQJvocQGa/KzGHJDUdYHfc0eq62X6u0
VVoOagwDYnxNfTCQhzszCNvAYw5UUXWTT+RH3Li0rgD/FaCB4P3dfKSU5Es0
zrL7yIpqiuAu1aBFt+/47364M3WXBx92C1aHVoNGVYWqTVT837Lsc7hmGouE
Q7Kxn0CllZwSvfhfGfDr01Dq7JGAKF2KIb6BQMonepLvJZUE52zrRN9uzDKt
qv5EYNzImlYMAnmMEYc++LQPWNcMUbcV3WxBm0B8h9N7sXPbkSlss+nkd7FE
7W3uBb2iSN5XEerXs2kqkwcpDf+uuUr3uU6h8Jjk4qjnX3F6xt1T3pUXMSXW
g/HP1QpQOHOjpkt28CO9JSFeiiN4+YWRXKztyqXn0G+f1ACwkjRqH/15q+0B
LdF79achqgoj5tA2NUaBg7QhZDL3LGlzxZsZu0HKDW0PCi03i0jlxxgGToRy
nXCaYPx+SbV/28m4lgr8eyyBsE4f8YzhqoScSlCEmOTz1tj/pSly7Ku5ckn2
AYSaqdRFEcJsYgIUPWz/Bgpgo9sSFGjA8X+iozcJJT9DRmTGaa6PnAmppJZp
Dg2+LPKap6Q4mD+W4eDs6OqP2bs02gDtTE8EoJxRpcvdFC7c6hjUQz+mLjX3
1oJeCb+OCr61YlmG44Gilcwwl7FtXd8NDSDcXEq3DELjSajXCFJqSzjzblGJ
l4uH37c81PEsqcVmUPSq/xPZkd1fRaMMZv2oXHg6XaxjthD1rk23YGJFem69
2dTiRqBjYRRPj0X8nunOqqgiC6RAIx6PUtryNFYk5BWBFymRTjKjlrtsjCQ7
ypbE96tvWoa0LQqoGwpQd7n+ZdjpuSP/FO1cBagi8Bnpayb73tFpkk5KqSvg
MT+auHtfwn69mvbFg6XhbaGD/SeXaHX0ohAHGtcd2h0cOB/NKUrXCVxESNRB
6X3xFCFaaK17drPF9up42GitPQarL6doIZFMJC+VYEjflMyijGR5EfZ24Cmo
6BveTs+3dxgoqhOYzCgoLRS32ml+sIeaj5S36i2miytFfW4fkAU1fvl0wgBA
YCNnwBOEgvAztCGt1c60bN3LDhHb5BZcrD7st8P6BY4WYuma0sWk/HsoqcgV
6CmO8k94cAuZ4tnEPlyi9EiraZbqdDr6oNTiCwtwCt2tqtALkXXYmAIUh5B8
TnitiL8feQIvAStXKBmmu524knwioju/TOD1GCDbAVfps/VBwM1WuJ8DUj6/
mrfLqZpNz76s6mIl8zk71j0ohyXiYT1PLWmSLx3W3Z3qdLpYq7RftLF785ac
G104vlGqzLqPVCfJ1ymuAQJDQxNuITdhEK/GcNj6OAOgtMeL2FuYCmlD/3ha
rycMmpYaYkV6QP6qhdtUkSY1c6YVvQ6kWBrSCNPuO62xIOVj6htU51LYYiQu
knFcOjbXsKFJs1k/2r520TLm0Jkls14T9JLSeDNQYLUKYdGrBn+1Z528HAiz
tkDmJJ6SdiPrUIhvjL4ktvFxMOuYvF6rVmhT1j6s3w41xptQ/eLiH+5TROFF
SSgnphqPbXVOTbiN0DJ/gGeSh7NLnPb0IZACq8T7cTLGBGohxATU9DhmOpbo
xBVJvM2FT8fx4KVj4bT3H//V0hcfJSsy31Mrot0e84ION4NhaHHYQPI22ZZ+
T6IhZSVbkmefzjccRiMOI9X9CPcZMSRiiwvIhGxDFRNSq2zwU82LCj5Hgl4N
YdLMH/x6A45Nr3KtHOcBHVynmk45v0XD4SCTE4bh8OwHCVoRcDFypmEKD30W
fGZeR4OsQdKrKSZPs4Oo9VZ21eebeTtB/pMdo2PWOYzreSG7T+QZptJdkIhL
c/M+StQEtjZfTSATJGKbgEBIjDjkPK+f2Te3EzGZ8sZe52dhm0w16yl4klhL
2qAITAlYbV9OgOz3SEcpfzUpU9xlFnaVenmF3dLKhfEVYJOXyJm4XqMGu/47
bpAB5o472m8UU7266583CjNgda83YhAEwu/xjGRPnL60/N/0eLc3Jv28Qc/l
7tiw3ys+MW7+vlCK9JCdQeR1WHxrlMAc3kjGLDy6fYF6I2JJ6l+hSHDnk9ea
Cvr0zPKcqxjkDSpOkGEp5m2BKXo224LYjyzWL4hTSVzR0nF+XM1LLN200KH9
1WDw8rsVJDKa3tlN2IDnv0QbHZH0bnc0sjnQefkE/OQnA83UfhTVDgqrI1xk
7lPUU8yLBgFVHR1WqwHEdVADwv3IjWw1zMLVKbmFIohguvmIok+VNSv4xY+J
A9boXIhO40fn0YGNOWaIu98X1iZ2x9YX4qMrIvDjYF0r91NhXgEcXZuRw823
jYpu3bmBmgkZsNrgzRJbhlaM7+NiWft1jtD90encPFXZsV6kkrFkoNVzWp1v
5s2TqJ6ZyNI4c64gZAZsp3+hZHcCI3tVELQwgnbzf3XjDwxOxlRoAgm5tQwS
WWXkVdYk2s7Q6/YcxYKVw8ac3K/Fc+7V7NputR7aRWwC5t2AWTBWk35Mw8dm
E9o7UqwLQeJ4cONLVFfVYUK1ly9c3PUvVWoDYIT6O5UNpwaS7K4wEKzEBAD1
puTUbjR1xJizrBMoQI0axUYhzy1yIiOl+5aQ1II7SwEuJfNKdV+pIGL5FIlo
0qTQsB83rnmDh5SuPefCm+3x4bXZHJLmIQbdlLPGoHEHO6KRD9eCJpq96IPd
RqCS8ZvDoO1Dn/QLMmcJHXEANzONoAFYIaSvcQI1OkM+7F136ZSqGvcwwmiW
EniNfO/DzUS1f7abfRpMbaUZMyGBbD7wk/UaSxnSMtB4krTnE6wOhg77DisA
Kl9h7XhW2IaBt1Lv3amauBIsGu3PgX/Y30VHbbl5KBntoTG26fYExPPtIBG2
dgXfUYQO953Ekhqkezmsid0b61F5/XqMXmjV08QV36RH6YqTQ4tROulqCm+U
d19gFfixqJQ9MS2IjGjRRLymbAtitnP7e/Mte/eAVx4vmHCQUbainYOvrNhp
FPbRahICs2VhsO3pBVXzRKoPlzRRmFe1n5oOqcQ+ofDj54QhcgLPbtTTZgr4
t2MoKMFd75C25MfocSXtcOpMRJ24pMVyOA7AVUrN1NTaqvJdUELNb6zlwLBB
dymphDiXyIruaH9V5TxRsCu9ECWUv9cflzN2MtyfgnB+eNDQzE/iXCQdGCO/
5B6A+bfGdn2OT36GCIC3IRslTRW459hwLKTlkv2+pMcrohzHk/ViK29whlCm
LixiPfQXFSlA6DqF77CChXYPtfDHUTINV1dWfnqvROLyNBaQPs1zVxB/wmyB
FYBDdUxWuzMiW0Cr6Mc3//WJy+lsYg1u+ioM84Ii2ktoSoqmv9JTBZxbyhJR
gJgIKcrU6njXyjhCJMT9J/5sak+G/EusKyFMml63vLeQtfTMgrfpWzfagLM7
sq5Vx0na2unpQnQlMfJKHjxnJuENeQkEovULo099D4hEEOLHD0BO5ZqfVTE1
OxIPnHTby3uHSzjZ9lhLe1oIl80h1VP8623AOl7EFE+tmLxN8zzGo5+RfFgX
KmPgqZpw4wNynFs/YREuvsWukDvHKufDqkQnLK1hKwLTKdfpzmhbMlA1AxPi
+sohPgzRmO/gftfFNdbRor/55WddKS0Wd8UTgGlOVAs9qU0sTDqyHMlWjjjx
7Dp1j3DhJy959xavS/dxDWLvhqRqSiqRR9mVqYkl5Pj9m3OJfqZA6yuaRaSh
+8OK2P7GHME+1KZsQPgbM/DhoyYh00NRHP1yN4bzzTzGbayL7S4fSkOeY0aW
W6GZ4CeyDITeN6/dKs1ZaK9CvGXR1Awiznm97pVcKkcMRCPH586XsH4OWnvS
rhjpAWfNcKmkBcVoU8UT0nYe6D0ytF2IMlshRz4N0yQl/dB4VvqjmyxFUziR
HIxNqI4UO6PunrC+g+HheJyZ6IT8KYJ+of+OCWDMcWnNFl4TDbfJaZUAjTdO
2QS+k6/vQoZBAILdUbOgcqs8preiatjvWiXdCLu1W307Kd3S+PQx7cubBH4+
E6yw71+xWwDazIUrzwH64kZE3xAGlOx42rn8DP5Kfy4rVPjFkCtg3Ty41N7b
eTFgJTct04fs6tngsm46Hr4AJsSwVI0eTHqBD7i9GYC1AsutTsZ7uJaRrXXI
3DHXFxTA4SSajOShESDsyYgsz87FkPaJc+US/NFqfTXgYY8Ly1dmltd9oUmC
igx8Q28KaaVoPpYUcW7HZbnjGbtYTm2monwwQbXH0pyomcIVi4ajTngYl0zB
t2HgEGYahcfZ2hM/nqVqEh4mSEs+QFxP613+C/Hr0zC8RbOFY58LfDFPAi8/
RGSqYFCcYOggXiMUgswOk8csRm53BJkOizoYM7USAZregVFqI9MdzIbVPxCL
40qQ0P6xFZfJxUTOCtI40C1IpAnpEMOHD6r0y5EvXbYm63HKFfQLvYQki5pO
A1kOU3meNKi96e4+ntYfrcJG+OzViOdEICUoV9x4tAffBI/gleBkE1su1Gur
zUQEfLcSv4Q66ZdW80XXYddps2wn0v/bsv+43PtOOJcuQRWA4/GaGWCNuoxl
0zPf2BHM2HWutmj9tTY5AjUZKdGzAmwnJQFLE7UVGJQsPE6BuweqtEVacu8x
ub9dlslkZSsRGJn8AosTbKqmZG3iun41WAZZeX8LYI8HCXZ81FMABDh0djOk
FAIHGyjGzlenLaGSTRqbHVLpKUXXDc7fvbNHk1+JcNOl6w4NtVnLZnKv0w6k
Q8sGCqjrI+sFV7V2CXU4JTar3ZVGZOOcdtCY6FhnsCjAXzBM02vGQiBRZVEm
7rUVsv7f6qR7lH12JiODJHpa2P3dK2OX8l0lIivcY1PLZMEtLESi696tKci0
tXtta5OZ+qOjlx97wc5ALI7+hXllXUvxVqX0H/2dgPmPDsZGOADpLkFKgWLT
3rYv2zfR9IGBXesHczoaFflcqjG1wTb6BdOck8fEymDFu/h9WhyRf+HSwFZ/
PSJrpHYMx+cPJnR4Ch7k90fIyo9dghEMmf3sT/buGnbRy6xaNW1/U3JZsIcI
cpLuwJU/BMhdX8g3JYNO94avVpX76Bn7/r4h8SI++N8fTxf4uKVe0XE8lf4d
ID7DubTEKczV7BFStywbGes2Sq6ugWfRXZ8rGRUv3tJbNEd6VUYr49EG7USh
tI1CXM2338EIrcsOxuMX4ERPrLodrZDqhO4UGBSzRgsm91T4+dLAmO1UccuJ
e2w5UVOaxo6EjC4fgT46gj9/i1oZC5WxxNEgG9YUElWBUiz4ucXL5YRUMelg
/k+X6my/q3QTKvAVGRA5hef68sZe/Lkrkvq3ntehKEWQi+GtpYbta4MSO6rm
1BbiHLzDs+k5E08eWkDd13YITbECDLnfXsWBmVWxUFAjFm696k8e3qeX/WXT
MytREBe1VZEXkyTXBWGdBCeUgSEdAdcOpzmUPnYLiqWJSTKng+hzCOmkAK1x
Gy12pinMt8hvomgG007kVslcMNZx52z7XtchkL52MV+yJc7CDgPPWS389Dl7
vVpiuTVrTYkNMwaTn0vbqN9PRr3Ey/y6a1zLL7azMGqzVEaWQ6kOni+tmcPY
nXkFiqY25XMi9/C8XEDAurGv8EKA0VNz2JUgrsQeVDOQ2AY3x37XQ7O4kD22
BDe3fEieYSwjDSy/TkQmjOIoHqmtImSB01t+6KdT/ZPKXOG67eCTVypFTSYn
NZN2XMakbTqnOIIfolNu9b/lQpYAdWxPTbzTzZ6Cnabzeh96kfHwzpS20DXx
DMTHoEB1su0uuA2TcO77nEISRd/Lns+dR5UR0HNbNhYCU3hoHLgzzNH1Hl6J
mgIIMxLYo1L9WEKWmFD54LkLhOoTZk4+STdpEQzStiAHdWp+Qou6Pklo+U2J
infHBI46TVNwy0Sz6qeUPOQALq5gTCn3u7tC3tHHwFLG2qYprYH0ZJbbqGZA
D6mdC0BdfAkFq6aOoGdUGJmUniGxcc8PgxkX3yTPHxXwY0Hqr+RQJfGTv+id
2L9AmgOQNUuUr6SmjX35aZqjIDHpk8L606iqI6oL+HGJ1hW/ZE+BnLk9Iozz
BpJxKE700w6VvJ2lVekFTlF3WdKme6QgUOp5Lkq5+QlOKC0+SyZcgxfvZ8rU
+X+/ZSzveoSKlse6HTqYGmyto+vDHBCgUDAFUWuyghFJXjO0PSRZIJmCx+K5
bqUmObS2kUKzybDyDUELE1Pd3a6gFgsvH1sIqxUQj8gqKvWy9d6F7CxgJGyA
dAfrLu0UlF1QQPp39KqSn8vs4Z9WNzrXrUXgwocJwFETdiph5+sKamdi2siB
HIEEWNvaQzxM9KtFkrnf/VmNTnHEQq7e7FoOI9a+NdRQ2J03pehHpte6hRZF
qHhX0IFqtNMRbD3yEi+oWEs7OhHYtBDM2/2v8GwNnbv9ebq67M7rth3P3toX
reIZAANz6DoBChPMdrcc1YHOv01eDXYkZeyvvswRGHrSQ24LG43yiOb29oaF
3Nat5aoP1EQ3Cbj208AVsJ6Zt+1c+OCxXn42VM7+l+6OMhz7q3wSrbbmPCPc
imE+ChMj1nkfJSTC3dTNGF7knTLaheg5h4IE0aaahj4czIP5Ki9LC1/iJvU0
x0hcozNGe9ceDPzKYabe0PTrwGcF5K62QJrFxAkVHX7dQuNz0mlJ1t1VmQII
OUUDH84CvAq0Z5xUTXG7V6tz+WHv17GjfLHWpqKLoBmZUAVE80jKKZCCxaLL
XPDoCB6cpv00YqsMU8hLGxCM+5/I+ayLDyab7ET1U9F/8b0MG/6eAIHcgwgl
MG5uAVad/rtKtsN+atYLgfAKcJ4UAtuI6DuPJRXQbDzUntPq+AcIXACWfVaH
ZT17SzVwZnrz19hlKFd8jP3dmLv/PYZt5B7PHOAm/OuIq+yXM44sF0HZKf3s
macQqvE5VZRfdZ4bEuXO+ukSHaX2UHz+l2Z+mNRwt9Me1Fv7wn+Hxmb9cuyN
lESPNBIvGVEp3AWqxL0VKm270PP3Q3LNlvuXE6oeasRVQxxWrtD6VhELxj1Y
Z3O4e6AtNlKJU7TZSxJKxRugEl8QA65Vl+D1c++urTEXFFivHeUD2BqgJTlC
FlQRgyB6Qx+UZd71cm9BmTW4715fajEbHZjtJ0GmUbORuHctGu17qw2rgytN
8auEsu5pdqfxA7KWl3jkn3KUDzHZtACNmbz1xjn207dfiR3xZ25f7/m3m3Cy
mbSfSZ9X/TrlWToL7UulkpyVnzebS3loKdSj7B32FB0ROH6Pq+mNf6dWt6F0
sbRDJXwhMsxEmxoMFLVUgFqMUNTemjNWdkJDYyS/D0C5nC3wP/Ggtm1RJe+W
NTj8zQonjtSu2aDtZ82ZmW79LzZrHRcMSyq74cwMXwwQwylVOrQpSaqsaY0O
nqJ0kl4eWKhqYiumXpPBma6gwjdz7Om0xrP+bhIPDa++cyvDbgeZSA7c35Tx
Q43wxHo2y2tNkyfxIsxdBRSqVkEscr7jweUZe9aJYLp7KUtqKrDTNZTm4sbt
psXL1/kw28XTHXd+gsAw+ZMk9AJevQe/nnhyRFMtzlCrBEgbInhh3BjMolVe
4SD/aSADN3MCXxCC3qnn51wi9eTZRMy6PAl3C7TnrGC/5HCwch/cMD78waut
2BA0YHT2WgtiIslwyOCIQANkDqC0NLWlZHDPnxUX6zTGH0v0Nm00l0SXQvVO
UO+LA/U3gI8u2Sw7GfbLFQBoG2fLUCES2ha55kqrs7T5Kpyy8j1cpaydSevT
lbAo1NTXXE6J1MdIdFejnqQXuvD1Cgactv04JArgGUvnlsiXUWd5l03DPGvc
BimJUZ5uBOJd9lV7WEv/k3H5pjv4dU4j/dvPTZ1wKMtEOl1wOCDLRMH1JqA5
FUgjGfbUHNGwV+ptL2k99BpQkm21tQin7JmGrHE4oiAgKQDWZclra2DWUcK7
egqs6yiVT9TnBjrETNTacrCgRkh/qxuCGqGSWLZtwdB1ZQwljGimsUUpUl/p
lzDl9U9Gw5E5ogeztl4fOwXaD+YwFN93nwzfTA/GzD81vOBtbxkQxM2QlX0O
jZWw+P8F4/W1dU2M40VL3hqUdvGoYiTn08blfo0mJJKIcuzs1GKo1HLq4ddb
iO0VeX1toTjIjCYvsT1TtUvvar8RLls3G42Ajk9pEdADqYd3XSXSgugSkpJ7
FD+42SeR1EYXStEbQNXUC22xDa2oWELfoA2RfiIEdPP1l8urYkmMlhQstEBd
os/YJkHRMALOhhfvKbC6aL1ItzRQeFP4Hh376MFKQAr5iVDDJ+kPRvCfuyt/
mobyao1N67DemVJ5y0oJ4i0A6215xUKj4G0TeZhZN0rIo9ZGcEo52WIRvh1m
fO++XJTN8/dX1Q8BxgPL/ToNeKpkYMZUCBr2Jmuwgxp+a16MfCy5YO1nfnKr
Q6Cx/CUv+MjmdWRZ8JYkVB6vsUpfYt2Xd7xp3VLQmliCnzIdtoj/oNHgCZx1
9S7Y63gQSRSkzD/UaJReWBeXJYxUBKVPqnV0woudUQffc9ff1HJW6sq0ImsC
3/cGfkiMML1agL30pjfyJ7uihLDgcFKeWyc5rYO1R6eG9F/MPJwxuu+0/cWJ
RvZKSjwWZEc36YCIyZHrG6vn2W25WNrlzkyogi8vYeBiDB6NkqCVtBSXBn+B
lAk3yM9oLA7O23HPed1xb3rFh/xaG30ijW5fwwy3OmSK2vkYZtqH6skVxHHO
v1yRcbRVBMhivcSSjEaL8wSKuKBTyE8aps8sKdPIuaXpqsuzXXIvIEkGWeB6
uuUdvUCJfcesdMe6g+x4sbZDfeb8DdOVF1oBPXi+SLm6wQEX1HLztE9k/WLS
Y6UBxcekmWdBQ3wPnLm6aRc2yNPUVQjoxSRucZyqgGf/PTJOsXxEB2kJS5Pz
B6HjgRGqmSHENYosO6wKsgfl9QNsdBkEdoJPYcyyZgU5lEImha3PsOr3jN/Z
jezm68JZUQmssYp9pAENQC/bFZxZwRxu6jpQXKCjqQBN7yTlGiSYXokOhyCq
w/YssB+OQ5IxH2R8wzTu2rU6906ZiyaeMclSKmI8IIbBHtO/HH99AQ4ut0za
c7u2t+ExtHaf4viYBp53bPUpsbzBWAlhWUaEfIRdRXR6ofRMD7944l+fcLhQ
FF4zia7k6XwHoMl+U6Nbe9y4RMnVn4+occdmXUKWTRvba07cM6Z0AQcAs06G
5cST8HBQNE6ZIeu3KOLGiEaNuT0E2NeU3GCS8eEYV3N9CNhqlbCsNaZHO2sZ
iSNxQZ52IGjK6rEmhu68tIwKSHW/7DLfD9pbWV7SHCQEg0B8WgcJZHW+Cvg8
ezb+iE09XERVp/LXX0Ho42opQr/F7CYN51saDDjudS7NtkkYf05nazgjxXfO
N1iljENplss0wYgcOPVlrVSQbT838fNCcAcOGKGE0AtrcHpc90YQsP9TjAG3
VUVTWwC6XGtsPCQPskJxb1T4iNnDWOfIFAfKA+Y93CBlKGLHdldSG5EdmIQD
Z9s+slkdjWPcqLQBecrQtsS3x+GfD0QFKQbdcUIgZAGykngch7CwmDmR8iMs
vhbw7aBesXnQOcV3VFnGZg7g7+r93AyhKmJ5g9toPnq634/QNFdwQrexJT4U
e/Hy3K74iU7bFJFxxl7/NbzdNmcVZl1G/fw7+pEV5UU2XHgrho3A1tv1kZen
6wFdEBtG5dalNlc3B9zIrPLxVTuGdt0yik/Fdg2eUIcxWUHnh9qDRVKNUY6h
11ovJm6Y9NVHk1+BSfya4wyMgws1HeqbgHqHhYHL7g0bypwVnrVHVDM0v+iG
lxK6WvTXVjGDLN9cr1RR0Gsvt1mqcmRzI+gjV0KAQMXwqCBMLm1fsrcmXWKB
9NWAK9dOY3KiEyJ8Io5FVs6j0CHocjpGsSoc05JH4wJMMLxRhxbVKyOQpQw/
/iebTZcHZY1E7ZJx+XZufnsRRrddDaBywillCbdNDynVba9KBEjNc3Wt6wM7
MbCu5YKyidcdo0rHocFOmYap23CvaTaNxGFcEH8YGRahIw/63RpfeQGMODmF
4lixT5mvKzBOIgMIxwtP7L8gqP36GN0tVcPkQKnJ3vsWqDHJ3bcrDK1CWhxL
j7y+qsv5Z56fbnCNWuqA3rpOeMh5cyRZwHqaTHxMIPqtXsRoiOGqinJ3hfOZ
jk4Qkkpm494DmNJhsdERvmn1fzEXED59VQB2K+CLD/ACjt8EQN/coJq2pZ6J
f1IE7X2Ey2HGsRzA6WQALpS7HkY0T0ysmsflmjzcSe2zbzpi9sWAitj+UFoN
VwDQ8cDdAa3uOayb/wlF0+Dz9z6JPOnvTzcfsZmuDZUmpqV6KE/iaGFiT2iK
BVICBZbHPrSZGMY+/bgGDyFn3KeM4qC5/ZfMl+zvOa5SWbsHaN9+fZe7eU27
unLnb/BPUmqP/nNsnTHFKjjQLFR4hiDw3QziWSLTeg4+rRXg56P90zpTwsuB
hg2ekjZXIX4UPeKCBwkQ3BLuv3KPUCRgExj1whbGiRCm552lHQqRwVVzuX1l
UVZk3WqsxsMxlrD6+wDYTUM5cinSfNBvAlCwKObYLr8NrBmbmnuPWbXMXiqz
OIDNUNQgiviHly3u9Fo0SbneEN8PcXzDhtGBHkBWsEx2SGIkpAfsukCqChSW
Vr0KtYdPB7G8dZr18/AWF+H+t9QcmkbQ8QzT7OABQ+J9atSskKfBx3DRGbXa
J6+tDugDD7BQTxYzb9NxCZPaPbGjJGfa/TwB7VnEz6E4ifcK+x0grzcDrQmC
zWhxOApk1WgDf3oAiTEm9LUUkNETClLVlTHKp3qHBA8JcTbG6HlBcPzYwrS8
HoPgodPJjiCxuUJfPGWCeW3yc3aE6UqfMF2tvR2vdX661rec9E30SeK+5t4w
sER+1mvIbbFqmnPIEYJgNEM0zdwmMRA+nvvg79RfmzjzCEQ90FNbud4SE+M9
mcD0lwSchRRQA9ajCX6JamQYPP972nAryVPcYgEGlAqSIJZWruVLz6yDMHxP
ZTJm9PM0SnkI1pSrKrqH3lNSP3/+qCtTZj5OfutdxfQFbnRhjjc08zGTasyi
W8Wp195LYgdDiHoo6lWPWFJOKlFCsGCVCJa5al0JKpBXUpxrmaNsXJOukuBc
d+2Owpr//XO4pqHBQBbBmkvxowWQ02Rjom8QDgHItiqVcfx2TwVTNRO6MV5m
xZutrL3UZ11QIfM3G53LS2lGu+ZU9Ev+9efMSUJPBjVPb2WMOYlPi2dvqRis
+9NQU7hJmNU7wb5ZmaGfXczhiSGR5LpP8iUz0VDHssK8rH6Vl5PF4ciTCxy6
wTmcSCmy9jdy0yew3OrWUVQNLSalWeDhmNvsk9bXf/P8pxKf9XyjqsBSK7Mw
u7KUVvJB9NNU8RksJOtzZKKQPM91MT9PL/623PNipuYiZw8hqBjsMyM9Kq77
GVKVJ7wDSpeBs4L4XK7b655NGyyka2Am5MrP+/4PiY6sWUsDbZBo/zNeE3me
IwghYgO9+RTHg7RFKnSKAp1hlLxRz+zPPBUV3LFb43fWm8Nr5aG9Exf8XAmm
i1u2BKewSHQevre3h3bdX5cA/u7rsBYCsUTcT7N2dJzQPsbnOeFT85+aboIA
ZMwrQ6cdWoQv5sKOBs0koD1uT7exPJQPqaQcCGu2u5y9Lr79Gc4NXgaEB5ry
IzQhPF7dQ4Ry2+eM+tvZplb2IUB/GQWgV0OQQW5vPG9H3X5iLUU5hPfiLebW
7ieOL74arpGR+8wtaeKMN4gybf7i/0XHOdUcCRh0wKPYSsLMX1exEm659qU/
V8x52uAEWTdqOiUF0j+5lQ7mdoFkGGtBhYBu3ESlIwolxUOw3FWcCI1r1tcT
OxHiTLczXRf2jZZOAzNg+HWmKFJBZk/09zVwpfmH3pODiu4uD8dzWiEMx39K
4obPBVkHCJgxiiUxxlhevNGSFrtDxCgmPjAVkGw9MWWBhAIkC1IpfRnPm/dQ
Hd1mFVJDfYUOy7hnRrNmShEXd0Eg8Mfz+xklB9GKvWvI7ahQqX61nWnf9QqR
jXaEdw4lh2jb+KPUfgpq9X7jaT2APqohhbeyZwRjpF8MAZyJNR4LXJkCm276
BtFJHLp9lAh5d1cuCLRSS3fCQdgD2M0a+c4cnsfZXd7jvPfiilCut/QYVrZA
AGYIBqZzCSWSoLsg+iGZDGnKkOLLf7BdIi8YZkAj8V4UY4Ghg+NoBhvDsUeA
50vLbNPII26cUTuWsMaBqblK2y8ohTHnfF3x3oKKLA3HCSGlUipZAk2hYshb
pd2vGpyJks+RMx2x88JOY39KLaeHNREq8vHznHsSabyfRW+VBUnFsd4HKMDh
agWCoBbKg7pXXoV24PdhxiAZQw1bvOi/8aFEzFi5BtvcpyY3/p4dRg+uv9D9
RbBfb4RgISkmiHnm+Fjhu/Ps7cGn2boHsUTR3D3wZlxG44CupsgreeWyFRPU
uJa3vYzen/gqApAz+I5+pV/zBIHcPYHIcg8jnfWBpPjYkV35MwIP+92YWjER
HaHJXNa9+YO+CViWo1kO+5tlwPLTL7NynVOYkNjVVTuxNAh/VnDot2Y7IYQc
GMDj4zXfL5Iku4+1EymoNHDlw36W9dUKu5sWVG0CgMADZxRTWsTdr7vNNI5/
CcK6bTaNUyo86ycBv3ktpFJ02If7qT659GmNi0AUQhlwoqiB2meuUjX6CYUD
p7b9szxsrj34cleukdu6MRcQRkKjLzF/fOneiLb8A/x37wZwwmXicv2lZdl5
7XN/SGIC2x32G8MlxbrohfNyMT7QWd42gIn8Lc3DLWLXPrjMz6lJ2ahthL9D
rb+EkPN8cPK6Vw1itAqp7WfE9LU8GhZw3Tn6GH9tdHxIzZtV5MFRBuE37VfO
M2IQy3BMvvDbCYyNzfeYXMCNTDzyhoZMeXMYN9fI8Z+796Dnkg7hDHHEF+/m
KZvzcwyB9HF7x1mibFmGu34Y/Rr8Mu1+sN8DXsUdbMpxmvQg7R/oPa3CNcPb
iEwEGFaSxyLoaYsd2oLFd3KV5jq1a2+bYArZ76c+RzU0jISuHZjBBiPyrWqz
cMnqSr3ZpUITuzelSb3hbqaBnyhphsd041FatKnJe1QOG+hcyxJAsgjf7uWz
VUVgB+Cuo1tn/IP3ikRyqJTOcxqHQM66kGy9u7UGNGKOOBuGQaNWHZ+P4hC+
tbenNmM/Ayb2jvQZtZK4enf/4NIx4icFlRILtBNKLpxZy+e1Abv+fGoChqDB
qQrNgPD18Z3mJhYD1vwpeTgUFn0retQvYjuNcNrkQaI95dRs30pUHVXn2nHu
Kl9gVUhFQ3LxCKqwwtYfOlk8ELX8pJ6zW2n+PSXt3KnAi6fBe/yeygIyxKVc
yJ0wVJeVs+NcR9bW1WhvtxMMkA188T5r4GtoaDgA+gfgoK0JBZD1F2uE30aI
CSvpGkluQ4xGfmraRbvPANA4PZwj2Ey1Ucv6O1lqKypzuTpYhcys9KJ3orVK
yhE8UuABZF0Hb8r2NFJNe8n19XryiWKZheJp+fEN2otzLwx6Rn/u6MfuusZ9
451J8a0agIy4h2TZCqolIWRvPsp3GisQbTvV/oxW6YA37Er5S8YzmX2GlY5Z
DMt1TqGW6Ijd1/PRnVRjDGfn3XtaPx43WNN54CX6sNkV61Sh3d1nQV43jc6q
5MaBhUqu0W+/aIKDmwL7MLOaZz2b3ZWji4jWJK0e7qD/AxsMDyle7L4DnlyC
J1L04qw+4hDgbU0XLU6/a8aBvNq2hj9TgNOk6Nd/y4DwrHsIAmA6HHmsPDY1
ztq/pCqhLLZSaM45lhOrWwq1TDhF7DQBhuhuaks6x1Q7JVre61TJTLr5mzY1
fPgJIA8wXTvxPHnAN69aNskp6e5WWsOufiZNaAKJYYAxCnTAw2vXJa9r5QgY
N5iUM4+4ayS5RNAFY02nwAJxeuHv43G060xIU5l07HSm6IVVggE3Z2d4MzF0
KO9581IGiAYKcRvkwDZgHmhYcax+jThq7rdaNtV1cmKqtYBBusK7ALSA82Rt
LuJgkuQOOOTWYiGcJHoiYeFJ+ElxiZAdmRLEyQuQyKhmZt5THGMkz1TqpXGg
V8WG8PVcttvnMDwsxAYAp8PPlS8ckrbWmbE9TZsXAEt4OCCpSJeLGVLZ9Oe4
sIHzSdLEW67ZrWX4GI4z9F+IJABwmeR1mjtw2n8E8dpmURNE98TTDcgstyRR
Au33rY08lQCILn6poCf7NFppjqIWyUGQ9/5SLYe+47ZNtzchUi4iwx6DfrHk
IzTEfhlnMI5JKnZw8TKsygFYqYG5FHuF5r1SdcE7Vh79zr9VyNRXJVqlxG8z
kXH83jmMIB17SJ/kpsFfQ819hyds+mUKK8Ye2kLnafoXiDUXPQrJyzu5Stnd
Yxvxed6tXqHemGGFaUDzbWdMTBX+SPRChre8vBv5GIKygNY5gNJfvE9sUKfd
9Pr9DG5PC0C8ixJ6CuPqGBgJRi5rMvPDCvNsZkROeP5UWthKmldVOZnUZ+3s
Jz90Pai0gwyr2ZNn8PTA9/08+Xj5QvE1BGaSQp5UBrC01l4ryJbdLdjcHhwD
A/epxr+B0LrO08HSuj3qzgyKTPzLs75cxaa+0eDYOES0Jm4JTMGkQNnYC0h2
xBBsc6SGXT15ids5lCSuy/LtwavBVeh3muN9po0O3X62Y93G6PlqL6STQjmv
h2NYHwGLfKy509ybv2u7B36xZENS4GWdjLrnCPGKna22mc6JXsSDc5jz6/k2
106geT/ruLvJyOr+048Q7Bm5m3onp3+dUrLIt2mIZ9FyTkBmWPcEzDGqNC1m
+6DVd3/2eZAP+YmZZ3LQC+5dYgKQ3QRo7e/eBLRen/8/DB9VUSpcGkVhEYyb
REALihzxxIsBZWAGOtjrjAFtU0MGYdZoo8RBpd971Wmw+a2PinvK6BEDMkdz
fOdqkdRvTM5MKRde8E3+LA7VOlLA9AL/cle3xmV2At7a8d9vOPJAS3dYKWX+
9uSWpC4jM39JwZw+8LKB5NQfAiPoQKzF3Q6kCR89FrNswYneF85y4Fa7nLKm
rZ9ihaeudWw96GRZoU2SP9b4AkEGxkwkoso9t69M6mj3HguXDHgMmgcxz/j4
Tz3Cgfh9CkD38lffJna78MR6L6Qn8lWkLUsPyDblVGsUyBIN0jRgbvpEmwLl
ogbhNVEsVAG5UZqFgqUtZLwAYA9Qy5NfwvpR/rPkBBXcJtDSmTxO9PYfOjOH
QjfWaQ1kfcs87xXcoKZl2mq0XOuvox8cJMHgcVLmqm1scVdETK0iWxIewn3C
wKByC+SW+REbpMobuQrV5gnOM8U4ocW1FHyAYAVIlRm2bd9JfAW/bhcUHBks
unzyMRWLuh68WpgaMd78rb9Y3i3HJYzzHjrV1ykfNoQOW/humdJXLocVRmRQ
MJSkbIQ4EEHsfyLf5Xd7pVOTtKmAZVWQ9o/BZwl0EpNlmO8eGNy/gY5vSNra
NsJBIvmLIc94vooN/MvFjkufrwUe9Un5LzWrVrQMq/5CsAMWQa63mLmwPwu6
J14XwfJhGO1SCuGrmt/bKlp+EExVkGgNZISvom0sHLSoJLs5TrCYSTBKl5+m
SFq3bDm4qy5XvKMqcRvywob8h+75qNvMAm6a2mYD0FEhtOM1Vj3V7wPj0iPy
Vdancl3k4AWfOHHUSMHYLRCBZtX1eA7L84i7ybCADLNIjYHIZCJEAHsjFuUX
ZAA7/Ga5dlUni0igDw674XuydkmxKTTbWWQ36+3G76z0TcJZbGSvX8O4dP0L
MsdIvXcA08FNnsSbxvOgr5sSdSL6j1gKlGRXFQvFqBr+R1esogUeBuxY/0QA
NENW2Qwm5lQuLwsLUfMzX7s5vC4nppIs7NuFrQbdzkYVTZggD5pG29znYDq9
RN0CW6xzRJE6ApWkQ8zVSbcZk3Ujpd8IZLnnajzpqIiCsSDSdR9q9H8oTgge
GbDJphfxLKEXYy3FVucMAsUwgdC4SfTSfKobMJDC5iXkP+YabBVsvilUt8PE
z+eyS7CwziMZtD5QvY0acRa5CkBz6WS0d8vGb33q3K27QUfn6wyL3qcqQSWs
rtb/zWdMiuFrIa+HbLh1OalRjsTm945wbTISn0VDn9mp77pdInWKSE6X4TjE
tbPad0CVj0NzJ5xa06qGa/z2EexwqKYSSyJko2wh/vegGkf1tMIsB7YD2nco
SC0Old6Kjd7szrU5jOXnvymIsiwru0Yk5LW2Iy565JDl3lVxCPnZSdVLL6hI
thJWjpRbuxUdJHnrc3ezavI7BVD82rbFSSsZ5Ij7jKdd86258Dt6fxOQE70c
wsZOx2LvF10KStFjiiILu0wvJ/Kl2nKs8VNY3GeUOZOdm5cLuPDv7lpxiTIX
RblFSbj6NsWrYllrRpAJUBxTDI5BdicnjsWyNYCj5SgKdv25X2ZEQtlqHFQ1
LkDUQO+d4IjqPXl01uq5snuVIX/1anGAxag/2Tg/rSm2GHvEvHlYv29BIord
eEf1DnHBmHsjP/W81nZcyr/LKIxLA9c8cFwARC/h7tNQ8zUkCusVpQ5wLg7N
SYBwfGwlIPCORpZKc79p3+achPsuXkvP5FK8bRRlkEFUgZnFTkleAzQcfL3H
nKGhi2PYqD2Tz5k4UPPFq/2Z3etcgLU5lhCBT63beTnT495wsKvJOuPUBi5B
vsMMseSrh80Xzh1AxLi5Yk5qMiA1av0yuNjHgq+/6zPcgF4bkzj+4NZpjW0A
Zj5O8Uf60+BjXG0OstQUaGn7wZF7dByfkOVyEQ70fm6zft8QdC2dHsvi+eJ5
auh5VtYXmVCNzsVSPo8kYpBzsqkgilGnRA4oaeNYgDgYztZj4XWT6MueLSOx
BRdiEx4vMeeBVwoJ6iQZgYaw0bk9lufDLfWUGDUf7l7kLB16J14jG8X93vjG
WQx6N1Bk5KInLms0kNOLjdP0mMgCjGt4pJ6SkAsYNOwoV9u2p3Y1UjOFRZk5
ZZfpsmIRwS33H1YWxyEEzUHywgi4HjXExJvTDKwbqpBNO/rCXBBXjS9N9FVJ
HkCoRo/H++YSfWoBc0Z0I9T7Z5p8VMo+Of8TFaInGcpKGbBkYdVYEBBrHwus
AeoZeJTui6/K4ZBAhffL5TwMtramdv6UDe+3HHBT0gPl7QtIE5Cu6JyCHSHa
oZLzniKjj3lACo7w7v6eNJBQddew15TIv9D1QIOlYdKwse2cNe5bfpXtv8y6
kyvVvnaFlQ3Gc1R66IT2VkIZe1F9z0ZlfbrshqKkUXfLnSmWKeyzfOlNfibk
rMqOH59yb/CJbwIfy9uUpdgmutJ7DqOyjUwoRHemarKeS6eKAhrCCteH/GOA
KdTrB3y6RB2cjPejJVsn0jg+iL/GmU0eUOcbZO3J96/oaorZfh54D4gFAEWs
UT9ySbWBuBKhUHCmzmTuixYuNt5hX6yoqksY3aPrfM0LaW77uVnLR5VE9RD+
AkcJ2vFR0eRAM7+05q0n8tUfezh4rUvnBwqykyT4/y13m3vm+9+uqKuGKDnF
QjYey6qRapiQxnoDhIG7xUm8D59DLgDb5ihg01efU42/DmskJHjX3ZFNHww3
6mSQ5XEn/eFHaawNTvXc7lLlx7iPpwydhxnkI25o2+DHX8kD3l+1Ea+GaRv5
ErvmUgRB8g+rwFArmpXm0M361VuDEh1XAB8spwI/RhHWhePBp4uB7vhkdJvQ
RvG6Khi5a2eSaVscNk4GK4S/nnorJ518nUlUhsa9T66rmIA2twz/GY5e35a8
RUv3BaUoe7Hu9qKAp4rWE1PhMfSo5rMb63uWts3lU2pYq1kVqI97QUpcl8E0
VXxjhsulHfWn+63uqRqzRwrL4DwMgZxkp485klMWLDxGWAGsbzIbkX1TOxmp
W9f9VLYP/89QxG3hl3dA6anFOv6WZphRb7XYOLb2p4QDLZjPKtvtTPNQVPE+
gf17VlK9q001yfYT3OupABAPFlT9U8hBbeyG+yZp39KsWwbz23z5vn/7eKuA
NaM2xLJ+rHdctAcVZmJNBl8FMURM5vloyFUJM/RBBIhALMEpF18/tvuCM0fM
ZFYNKf+NvKRgZX/N6uqlyf/PFgu+c0m81vlUUDB56eGjjRhZgf6ZTh/kPhBk
PVclKJ13tfG04ANOXxjKwxYeqzOwhz474VYUW/Fte2Dg9SXMoim5mqHAIi/t
1jI98GC04eduG8QSbCGvAvU/kZm606TrrMNmfAIFIwLEgoycJQmR2JAAVV2H
vuZCFU3UNCUXgfIcU/MDMF1JdzT+LwWNHDBWYnCj8WMbEcq9/DZ9tQAZSbYS
1hA+1cQ0Gn5lgGaiyNzVK2sXQ0LiI3QGNSFEEwR/uVped3TQ3pIQvxxORgix
ZE58KyAXQTfVB1e/HQduBWoMxKsrSktWRtRrNqJHr19qJXsmTS9WMV3DyZpi
7CezsmJpIn3skKBfxh8UG7Ee1Y0RawbuV+IM1lXaSy/cHrlWYo7Sn5bbiHVZ
pu5sC4c+vZZNmuBVLT2BVib/xtjwz36JnsKdWGcMKHWZYCdDsZOGGBi3SY/J
XitPAQpGC0lXk09J7f8FIcz/SXKDz7Tx9TKCPN9e6zC+heV3MWlGXM+Pbn3g
nWlzZQXDKn/nJlAlhXuXDQlRvRZZ2NV68LHaMML4ZxDiJPWojWQSKH22aLzr
8zofhxshbZttQ/lFHVWoxyYXgCklCgUVGYw1FAsALaDUcuRiM7THSdIn3uVG
kud8InAxo9Hbz8aIaIPnCgkzPHxRKVg/ZsquZ1TTxiw20mketgqCqeYPyZCW
3FMvt7BVEoH+D92ixUjsaq+dYNB71hBPXnG7ntEEWTfgLxIGUagA7kHPVZX6
oFi1uECcesmtfHFf6FDFkth2Kz1MZiODoDhhnimcm8FG54nJAO7zHLCYhaFP
MdyCVj6YBXhhlgcoN6OXmQgg8RU531r2f2kY2HiY4lURG1Wgfoyptwis+FNU
9Wlfce69n2MEM/z+bCegW+CKrbowlTMwyC2DBg2dpmBKQa4AZcnLeIvSaBBp
siuotSOcTGr26dpnEER8kv9ZLdJyTNbQqunBXegtWdcKba+iXzYY9u7KcSpY
7IvdIdBoW7Yb1ou8EH99pfAbLwHa51cGG84I38DdpLShforfZzsGOMZUwmx1
DNrGRsYFEnaDAQOS+Cwzh1ISfNMB8co6LdMTpzpBeR71Vf1BEq0xb0Wdms6P
F4DuZSa24JdOBEQBw8bmwDGU3s7rYZC8oEKT+MBvmXbjsugWgnajITdfVQ+u
gVthMEfaTfGao8JHFCNUoy6CzWnL0PyJn6INTpfKf+eikQMWcQz4pxtBC7aU
iYEeDQUs7VZ9Lzuo7mXY5sTCLAjCMo9/9iUHl68huoD9cq/Jm3HDL2qvGKve
8mEdgXkZCkuM3rvBUpZxdrlhz20Em3PT3jGa6htLld/6QQr873Wy/RCv8v+3
quTwtXMaS5SFuHHCD5xDLADIlPUnkZemPpSdYTeCxEt0UHvgKpuqCvHXrg4r
VxpW7nMpW1rD7+/3g7W6vwH1pp8gcPIu5iTMnOqGCoq1zJgBFLTKP0L8eSEL
zykWO4vhfMnp1p6GzQPywdEoWAaJhr4XWvJWq44MWkpfDwBaaxHmcW4mu9q4
m8wu2ZVqFQpaHhWT14ZPKY9mBiCuhmD2JmkC/f8Lj7dwN1eMo9eJDpMVRMUr
Wwz1+8/bzdbyqXirEgVECR0bLv45EeEkfHB2znH2kOjSW0BFO2qEcArLmOov
2FtBsjotKy7PEB/beWACH2/1CtcsvOUw5UeA3u/ZWM8OdBrJZko4C+AL/xGj
iURkpxRkMP03sjzaLdzLsDV2/0VqgdQIrbTjKM0JqPm/J0C+j+ONqpWW+yU3
tAUEk77zCd+kBOvCVm2+LxjbvxSu05eyyaNy5ey2s2yefyZZaxKv1MTupGvr
nh5RE3SNh7SREB/GZv9llTY2Es9GMXltAE5N6N71j+xfYAt9RAhLigkOXsiY
rm7uJxVAtVl1ynEvCp+E6RKT6jyDkVFxLEY/JsTrvn1+/myV1CUal4Nr77pm
OsoNJpdVX70F5tfM0napqu5r7lL6wsWMyfb0pk7y83pIyQcZx+rByXgkuud2
yZJMUl5q6FKOa/Z2k+mWU90P1Xqz/HmpAfWF6cNCJuyuGupMLfwxgRlnJUQt
lv3gf3S6RhYgEsdQVj083sVOzqi+IfS22f9lNGxDU4UaQJvxXOLvmfz/TG5s
UExYlhrKLunm0jX5SCPMubSqdsId4lkFx2n/61Sv1l7SpdZtDfKahnshOfDf
gQNoLVlZoSF23lvjgYUEgvRf/68ERLt3i88dMoy4tN9XU5fOoL+/eHdfSxVC
yv8lXV/G27IMj6SSjCM2gPPcyBUisNIPaIeNTYb6PDgupw4XXBXkzxCWaBQh
vRQdy/WK/SUzOoc95o6+iwpSpwNajucQ6pt7P8OtZ/B5KGD+s5DbYT9kIj4o
e2jeyjQcj05lUII/7LLzounhLnfkB2lgdFNbXyB1yUOvYhMucksKZYEaOViO
2dNjHCoBg+reT2aRPhx9YFfqC11JjgZD32H/uWlRPvBAduKLFaclY2jYObzD
r2r9acoyJE05hufejJa1WjXXYCuKtk+04FC6eG5k0ej5gHQDW4YKkwfe1HyX
qYB65yLl1WEryl/jgjZ6xg3JEAA8fTZgMq1XjLBxapw+m2EvQ3jelMZoc0R8
+sDfYSLxUdm9t37DRbi341B0eKid3yiFEIt3JL2M36CggM165tsMl5Efkiue
FlWXhV/wmx3pf5UvxibDSHU1D0OtIfj4KZOHsyPsGgaeJxPrO8zwHsV6LxyF
aOS0iW5DtIeoM4quB70FBUAfYGlH1VbXjTWOCF1KimVAV3V9C3UB3MXSQTx0
UNJCOJF+ywv8eavuAn1N0AuTlHIJ94CG9e9NV6BQrERLsBTNhUJgxZNZDKrz
Ds7hjaoKF2JdBlNbj3iZe7+WVq9HD9/t7IrXUo74Tu+4K6EeUQaQhSe82gtI
2KtzjzFPm9ezmsdz/W6vRyMblvf556N6ufRB5LMvdHjARgQztV/c/Usqhl2v
hrD+gPwnXY8BzU/+6YiRKxW2TZ0aGmM9UngNaPt30/DpeemrInR9ttyRcgxD
XcU+pE3N2JNH9FSsS5p1fWlkmxFSQhH4vAFF+AySACh5vJijkpxptT9X/3Cq
dA9ZkGFk7VvKxYWt3I855xlRd8AMKRxf2MU/nwQRXVH9eHCVjEJsLGPuwcUa
q4dv3IShFaCBmcbwYJR2kkXoauxaNCO+jVaY8ebKmiCPK2M8SXeF/pQ3GKkk
YS0iLIEJlOqcg+3YREa6ITcW6X1iQd81QUvyfs/gXy/zwz8rhxGY+e5ObsS1
IX+goKbVA4UikB18qHeC/DsQprrX+v8W1hWKvOLt77rG+Hoj9qyFz0qcDxLz
ZOjDWFsLCvxbexJqYyc0VMkIR6qvloGH56JNN/tDtO0aP9ShFQPhSTYHxWCK
RNxlOcJ8tCnFHT5IycWWx0natHG4YBviuivJu0AnJruItotFSBhWZC91kJmo
sjyH7L/Xm1HH3BGRiaU4i99Of+uAWkS7LmFK+OGi9jSB1GpvoWB/tSXePwmJ
opp/Vzk9ilxMBAZzRrO5/rrR8hGoRmKERB7BJIT4zxVdSHkKGs2d1W/duWMo
gCpYdEOcfGPyKQf5+QJpZBoEepdTgkEoUmP8F199KW78Gq08rPPVX1GRb341
wJXEFhGxh5V9v7Zo9kkn5w9Fcfz5mz4pXE0OgKXswZT5237+SzAr9RkAK/28
8EedMgTnl3iCWTO8IFnCINkzYP/mA5uSfOlW2pPgpfNrRpF6ERwvNUkH7OPz
/tbJXRIDsxAIrbOSD1Jqf5DczsuNn7SUifdgh7Ld7vGMJzXxf5OvOroLFZ4z
40E5bQvsJjAuWAx0SwAR4GMY5G7DzCoDzODDdh4r4gaacfwTrYl6Jdh3wO5Y
0QpK66L/51PpaNlXV0wJJ2UO1i12z1I4zF0nDYNdzAek2LlK/m6wH+LwYQNK
9mfFBL8dfl2tuFi+dTnAUuWcsoMLH3nCZuT3+KeUdIkl9YweMakZo+H6bi3A
VXW919WrvoeCqobu6JlY58+Rm53gJFpIh/boqpHIK8vSvTM3WV4gLaIoLq78
85rDvxciCxX+QkqsqnQFC2cK92IC25M84kOxT+qYPpzV3TjcO/FSAhd8gydN
FFBd5c2zpBJV7zUEz5eexTDnQlgfpgt56EtmrKHrGWZQRUuDgRk2lVfASVEB
mSlZDUsg+XYl+g/d4N/x1BeLtg895f10XvJo3YLLUabL0EslOz41nVWgn6vJ
4dUNSSbh7haoXjjqrZqFoYGXFmfzUjyVi8pGvZDg2cSLiYmcGG/4la0Byfq9
bqPwG6rtGzFYH1LB6XsbFBI952Up4fCxiy6bV/Gc1QZZT/MHM2KrypsbzOXg
X55fZxGCZRJAiONWwz6s3htPSaenku64jQ0mM8yzNebRHBytQ9+poYuLf0xe
NnVaJWT8PrYDkasEj7+jeXMsJpNEUJL18xvTiOMSAItWZr58ahyWjFXdbi2K
0XSwv5Nm6D13hWyb9mcYvWgeBrmVhGGSlKfvpI5MBE8gMpDC2sFSUPcsomfj
sn4zhi389yZ+BLK6EBZLPclSoUcSDh+5GwhIeyPeQCGNBehJXANf+UFzV0I1
DRbWOXUstIrti6gR5JPqZqFvLXkAhpKnN9rNtC+o7P1RItzmlBGX1zw63ou0
Lx9UJ7LW4pAMFKV1TEW5Gi4bQWyWnTXYZX1pYkgX7gZaqJbJUnBbkvr+od/R
AY39y9SbEEJMWcxK+FHaZagFY7u64DJ+gZZQPcYWSktND8JH8MRBex8gFO63
ggBmQh5CZv06RRyDWP6A4gqDsxOCLzJ9/M8uABKrcPT4b8lltl1tkAIlhwFz
KdrNLDUDojXy0TvF+qkfFboMb+SmJjKLqVQAJVyBGyYYNchxeblQ4JhHVx1E
A0b7qubhuTmdbQZFg2C7Ah37ST7JUTqOse1uyy26autRSjsd/k0Z7I1bNvkF
NlZ8DTX1nDXuOlypfG2NROBdGeo8Y+WBpRMLgmn60qHNTwllGMj1RwQgux1V
JSYqssgTWIi+Uf4xNyoRKkegcdpNNv6Bbe/gLlNJ3ghPU2ARN2Pa2kKYQl0n
jd8r+k4XakstmnZtP+UxJQ2K83TGCCiioIuJGr8qr6y2QbCFZhMazP0SCPoc
clA7aMpj0Y05ms793gevpzVvMx141fW4zy/eENHgfJOCK+a/2O7lYUlk4RE7
GY/8Ny3RjGiy+A6djWN2KQnJtKP5dih/PcKqjqzGqwz3z71Xv66Pk1CIfj4D
yfKvOcG1l1aFkgGi7y8Ye+UhMWVyYzQVr1uHZp52Nk0RJAyzePwppE9Syh41
Gi6B2va4T3dY0+yJl9dpFgKmtMe5X3YQRqnzdwJBqB77RU8vHdz8YrfjuRU3
4DrWoJyNOD1RZsjehlL8b9hdnSZUqeJCySYwZEWM/iwgKssXdhGHBVOKXfhY
m2wVkd/pBreJdxaUh/ColtFxRjzTUmBsEkbd4kzu5UR0m+x8ZXnwQo6hbbfX
TbJ52sFe5EPfTCKpM0KHcZpm8GnQgqu2MwBdr7gejlV5ML71ptthmwFlU685
vbxtrnVGcvtN63zvfCU26b+zOd14KZVwjYXZQv7FEQ5Ie1oQjbKDA4vS5ckI
bNO+nHJ9t+iKm8rP/btl026NWbXOUCX4cTsJDfSICR6X1gKkzzcyjNxXOIM5
H5M+t++eSkuyZazQQBmjF4TtN92sm+ZNJDabbALl3rQPy7NC7bQFacAFOywh
VBlvZAPiDI1/MVV7ksZpn0xyRB9jKywTjOpAynvKTMue5SGv+ZBfZqcqNkmZ
HTtLvomkN2wQ6kxITatxn0buQ7kYFa4/bBC/JvbLie8dHcAt6dBlQFWSJUOC
0pdQm+iC/NtzVd3CZTAnDWjTh8Enir1BBPkgNl4TN6flf4bmubDC7S1m5M7d
xTlk7U2tcniz4kkgEJeWkFfUIiagUii9P6hYqYWjMRRiO13LsL1+TdG3jvDP
CdX9jZGIr1HiGOFMVQvOWUEt0dBIwKKFMgNpYyAFhoSWXqKDuupQQnkC5HGV
O2JgvovThfSqfskJKf/wiJFkzlAwvoB6cOoeBMhdJLHAuCcUKOc0HzUr1lHI
AUwq6vijzzEhfOY4HEWCPCYiyW0VIsIPpyz44oINh9s3JXglEreL/lVKY5P1
Usw/QguZPXJi6H8xiBOdmMTEK7gVqPHVUdTJbvGbRni2CExy4giX2VqOI1ZY
wsnUz8Igaclz5m6D4eJQ0YwT7bBkmUOqNOrEnh7ybQ9E+hpj86twF1eVcR1i
evaSwzDlfBhMQFG5uogWjy4cxYxLccyw1VmtkKs+ihuzHQXW7ZxfwgnYSfQb
YjfAM4jSbjlsVOSkeMiLkb6Yco4a5c9P4tr8WXGoGMNhjQ57qDV85XeTywI8
GO+0pgd3nDE/5YrsgQ86TwIDdSvgO+KUb/NPRMb3jrFx1z7BXwBLmTTj7g5B
bXhhlQDHn5hn0pq9ZjbNgWrX9FEJ8BXeNoPMWZ//F288bvn/GP/GRP+EPVB5
fsGPChdWiQKu9TCmD7YvrkspEG4NfFpHbqDbxFj9nSVH2GcUiSmYptZyb2f0
so1EJW1dZXas3Yuu5T9JD9jxyLSS7UocuPgpZBX5pCD7MJIbCIxq+sbtnrI+
bKEXs2dXARzNyw8LkWYc5mcchT7SBeYTj8qgY2RZiVpvOEliDi1ii5jvnoBs
5ZZSDLmJXLB3OkOy0QhkhkMTo0NgwM6jHUIZEB7/m0IffWF75ejBAMnlv8Lb
RhwQGDotaX6qKMUHkM6ZqPkQm+wSPJDyeS/dw0Fy6SMhgmi76D9ltOB4fwnO
rWGmevOt+vUMgY4YlD27htyobKPqohL8wmd4eb8+nr8szBOlMzdd1XH0zmsz
+9ImpeK1hYDvga7ep7Wd+INdDD2E3zvQzJk6m6UmCDnRH9gs6KQD9NbKb2LD
MFvlPq5oSce9yIBf7c+SBfVnFXYaYuqrdSBckT1QUzV/J3avF1TV/TZKfefp
WjTflY8jiUiIs3+/zDiiykwWGAWNiXaGnwVC74VnVx3Fx2Sr+me4qmuPZeWO
5p6gnLsI1Sjx6Z8tgSFDDhD3sCsewwsd6yl0S3sjS2j53/BSYi8AfV7cFQwR
RxPzVBTr/aOsk8QeGwbsF3j+iRIy/dU0AFDAtdUmDIpqKKmCC9pAeyVe9hQU
yPw8TTr/upQrkBxfS+m+zLFhlZYTFGCYo9JKb+5DOQgmhgNtikZGMQnM8AM7
kaX8VEDGvsZg3sOswX4w9W/zZrIgG+gXjq0QsA8ohldxNB3wNBa9UEWviDxt
ROSWFszj1pDhXpBB9K1bOrYQNAsFOFixYjYh6+vzVHRfqNaUuqZhZLTNj71G
l9AB3YB7XJRPGcNicX09suLHkiMEvINdcuCz8O8CecYvD4lW9do/0N42Oozz
r0VIOJw8VzSBIJpLuzzWpsm9F7/Nzbc2mbpHX7oV1HPu25lybJIA59ktAjLa
Z/mW7oPX+Hx4yWJUMdikya4ocQApty6i1o3W1N1MkBOpH/jzaMIzybwOyhtm
CBmCYAG2JuFaIILod9xZcoYbq86DnMnZjwZvsqdlC4ckeqfn5Z+2xsTsrRlv
EL9Ed7BxxYndcP/5/lsCjm4f4SEfydNJFXjkCGbw1walawK+D4OSo8JS502o
tPTkr6Df+XoBKK5bjws0A/ThCLsAutS7bM0KtwoH6LErevwYTo4tjpv6Pbaz
aUgynUNyHZYxy1BCkXb5adbbZzr7kfzKP8JCibyuImlQKakN1Yygt+36fQx5
JNccNCv/u33dMSd+ViV1RiY+x2OSnrdsQPxiGBC3EWXDTl/92ktT0IXbZtkV
9F5fEbPStt9blQ2po+J+in7A3WzD28O+iU8N1HjJmeAW5sbIuH+STkwQX8J2
MOb0GkN98SzdeRJdKb7l4VRm+sq8NJIaFAcAvnSrLSW49mDeSqFHljxuvcb9
F98718lFZYZdSqfaccg5HXIf43qjxRpLdZf9yJEl0uAaQnh80+MFsP6oUAub
Tsopjnm8PNUaTaS3El56JlsNwFJPWy9Gto2HGz0TDzcsbblLXtLZGNYJMNp1
JuPlBl7ftF4BV8zjB3DQCZc5NMcvAdmWII9tsEfpJ9ninHm/t3avfsXpX2Sv
LxX54/iUJZ2w1FVeJzZvi+1KPAy0+ge48Sim4iYIWnmSm1vrTkU8H3MmH9pX
mr7IwoC5hEtd0Xgfz4gCxGOygODjrd8lxkW+W38aAOaMUEKDqOR5bHWVtGD0
6PJ/BkEZU/0jcHkLdPlF1+YwkWCDGiXueq+ujvawOTPcPJBwdkBXAEY6XKMv
BkKEvy45erwyvbcj4D8nH0d8sNZbz+MWAq3DhTfZGrVl891o0azUZb8V0AtT
R/8VXlqa4YRtJgOaJZ02IUkds75AsujsG+s2zoWZvv5KQvMMRnfRhEJ3FjXr
MVzuyQ8uM0BHfkqSH5Ch9oy2KuqBMhaKSl1SFKBU2qAkxhlMxHl/3Iq5AG3v
rxNFO4fQaSP/po1HosNNt2JJ9RkzFyiPwyhSpWFe0yoJnqHutOIAOuFnN5pJ
39Tn45KiV5lmFVtYl4KrsdjLTNoHwF5iTyjGtNkEXORvrL3nSmyedvinIYOQ
RgADhrUQr5PGgmTfnsTQWr/EQ9EM9ogoemEZUxn3w/MCeUdwO0QL2AYY+4mM
UX8/z7Uptyx+69Isxbo04oX4ROo9X0qEb9Qkny9dBu3M2CWr7Q7dwSFcJRaU
zcdWV7Kdz2y+sC/2maIeQVuEWABsQBp7rCq95D4vPnlkOLYeROLVC0yyw9Se
SaCt+hj7nuZuOHrcLtHr97D3eqGLbUUYOKLQ9M10LNoly4NI9kGBWt6VDgSf
niokUJ+QuRqzxM+ceW9E8acMV0Y8aAw+MvNuyB7PqeVWww5NEleREkwh+g/h
xbGbkfwShUelOhvHVU4mOojewEQdIgsMnHsd8e6NWK3+ASKByVlD8asIFz1l
j2GLLVNRwpK/2WQ1//fppJqZnVDZTjylRyq5lSr1ojw/ZOcfMOXh4nIXSmTm
jwOrJU7zKlNj4mg8JCHI0/+E6CXEyb965NlomSylDeO5YptfGQql7KDyTcJb
iP/tNTiPdftftvyL5KaXXm4RcVJYUmICmSGhgaMWfAqbwQjdnabapsL90T3N
Hywl1MtjK96TQgUJyoltY8psygVY6vjm52MUJJ6RAcWuaihnn6FuIjmQ4clJ
2DNvJ8z4MyWfzVXXwgtkI6AVE2o1Ow9DOyfbI7IR1Sl1N3bjXbalOBjwZMtv
5g+COPMo68Pv2bSb8t4IE/L9RrmWg7dSFLVLpGcrrY7uJnehHo6/qkzh+DCZ
HydV6mFKb3Zsex6NVXW2rBKsXoLwPptjoVEJ+Wq1db1Ukji64eRD1F8i0C2Z
8WcPEc3vtg9hiE9Wfi2nxNPXplSEUfpqk7Sis/Vdq78UFk3y32fZ7hbt2Po2
QtPMW0Q0P/XDGOoDHjztoU0FgMqzr6H9JIY2d/FReXesAyPy1cHS0822EjaS
hwhUvIIFkiuURY3nzSXkXQsXSfWv018DaCiqSMxjd6q07GZ9Uj3UJcFUqRgp
ajzoi1hV0OxAEs2/EJ8v36lnC3DuxQcxW9M+1VLdX6Czz8uU79JlrLSUEjEa
2111BJJNpuPmDS3h9b5ciag1u2ocKXxC+hOsjVn0WgY53GOdSrjQUwzB7O/W
kyUlqbmWGymVRqC337u0QwdopKh/G4XXyyqt0ahQNWY3Nhe5mpTpH7NQQ6G1
qdCffXE6ULQgPeorTwr5pNwtd95bTOISh9R6/b+Z/wUsbSa7F0i80Sl6L2DK
SBCik/TJLKQjBMe1AEVeufRehtCh3F05kF0brtJv3fi/5Tyrh+pIyenvm22q
7bMpnXBFy+jGSJHYGXTbG9ZR1uGskU/FK0cuEmYVnwu0H8OrFTa9nAbxLV1z
GrP2pi4ZHky4p6vQHEFZ8HrQAPcm0N1LNoHtdY1pvmHGJOwGkd+eLHGCQG+w
xYTJfdn2zPWlXtMt+NRpRjyToMx+TqaBbTa9rfKA8XxN5bXIKy9U8U0vQ5jW
Et7aAtyWpfzvfSb4keF3UfBSGVekuczuTIR3DQuh/ocwyRqdW110rwd1vqbF
qilB59Xk7AvqlC2H7qLut0ghxqTBA9lrkVAC/CZg0aNQ1H/9hETmCQZ9fXMw
YfrgZivWXKYxHe80LVlKG0UZqENi2gg/vyDVji71X+HdLAXspLGArDBcQ00/
UOK0NlchWlI/JGP629bWFGUVtXo5khKmRbztLGIcrh5itRgRMRWH5m+WV63j
BYnxkLS1ocrch1ezvAaQLB1/mRklGIGGJR5xZRJNgO5pyxHpy3HcCwTiyPnW
2IyTMtJsJZOnsmDRXfl81koeZ9WDqZDm5pqP4zLrU/bfZfj1Jn/QY2PROi4T
xTzhOd1ITT3cXPu77a4Q3AhJf4LfvbqPqW4BP20NXv0rwcSUdI8D8y3wwJRJ
5tI7Pq0w2miFqTlfluNYJKqvdXga/kUZsqKo9H1aXvEcTeLJLXCeQQgXfrNj
Cf/WppTpM119YqpxoxGWNo4cNFtumKM7oDGEx3vKvJ7HjSGXToUs9WHfp0yQ
LvRi20yJ5tlrRHIjTLMRAJ4+kKOERF9D23VINe7i+aFzFukE3vcQmY1pJlPW
TalhDAv8QKliHm+I/7qar6fMEfNFhQ8xRmPUxTeNpPKKPWx/7x9NyZN1R+O+
obmWsD1lTdVeR7V6l/WbUaORPnxWPgqvsiqB6l1Z+ENlNFdgBzh+kYLbSBDR
BO53ivHnjngON3ZNDNEZ528M/5rsyW6u4ryGQUhJqdX2r+kp/efC3hqTEGtZ
6w3VOLphLhBeH9HF8M4UYa21t4nNYbzed9rcqc4TtrRIFtmty0naL8y/FWZB
jCa0Rn98WDYnsYvtoNAMjAdMI369ZwvSPx5GAXwr5ktDANEFdcaeDBJCBK/v
UYdXq5Cmw84lXd1+yPluw3ls4uQLfH8vlpXYv3Lr5V9wF8lFHPeyanfk0OTv
NYNpKH0+DiLSALqJyKg2U0f6k1PeY5qKnVvybalF282my7rSJRXrJ2gMjhOR
EfcFeb5nGeCsaiVz+aprbLXg3Ms08YGmpZr7lJ9g4FBLSkVwGF7U0bU9oal4
6kMVODFglyfi6WsRxf7GvvKeJafEzELlWsZlBgeSwLmR25qau5aILXyUyUJg
fmXpCbpc2upt+tlmOIH+/rCvRHsSN/KiW5RbSdMdspBtGr7ChoKmdNIQYjrx
aRlziCDSJiiTq22FXBJr8pY5VqFN+0t55hHxxl0WViDT7WtsWufWf37+CaPt
YoACqjUgx35Ivcwa/SLVPV5XefswqMRt7LX7Nr3jGw9soXjEIembmyFboN39
4pwcBjDQlXhrYBzivesrnvZMYuVMCxkE0kxzfwiV/sIpk5Dea3eeUWBj8t6j
XlGi0lYgSdCDk2MRIT9mZxwFZKMT0h4KJOPVTOiGzyUJQZXCPEs7I1Bv3+1j
TwVDwR3LBiPmQwfXyWix8Zi8TL6MqRNUIJq2dqdW68VKmHF5zfZcOCYWqreG
08PivDa1Ws069xoD+6wGYqnM9t/S4VgomaJIKkdN/zeRoIzBKYgJ0d321ek3
8CscXoME4sUXKilyNAikwhBYMVbSVf30IDqAc9eZcP4mNHiWjFqYeeuM0/QP
1TZmmAF0Xoo8kqlWQ94wVCtPuXxuJM11gafON37+ktPOdI5Eu3AjHtHjb9Xw
BvYpZIl97GfxzhLXgrHEgWHuPkI8sqdlgU8+XVjKaJpUlIps/9i5COlloyzO
pS0Q5ihNhK8VgKcpC5QnE4FPTS2HPCM6cM1d8QmTK1fSZCttv+i+a9971KPO
tj+AAAWTTnE6mdfzl1PQbKXfxlu8/WRVQNsT3+uI2djSHOtK28mNtio+g1Kv
FfMpKUuOVLLh/NvEC18HRnUGjlOggyKj4lhv3e4tECZl2LBtXW7+82ajYVfj
mjkM+tJQgc7jUQ+0lYZXxg34SLTptWn0OqNLq1oMkJLIruh7nlxey4B5h6+f
NA8N7uzZpwtYGWUCrx8UGB55YQJqKpVrmR35GEzbig+sn88J9v5HT9tuaaac
0QY6coMpqHeXSboNy3zTdtyqNNzD3rqHWgq/oHkiyXll7XYvehUfyaJ+QJWz
ZqQc9a+rXkJDN6nPOW4RrhyN+Vs3mXzLDTgxnp7000cgIAbC4kujtZQe2MGf
H8ZSTQsEfxc2ua+bNrdsGIw6Z1AM/LuHjKE9Kw0z4R3iTCketNNLoA1q6ycm
05tOnJxybOJ7c2Zvsml9OUfMGw272Q6Rhk6U0EKGqiUrn2vsvwH7wwbHaZRi
qM3Xkm5SuI1dRY34Kbdltsay49wWIol1tmyim0xLmAbK3M+tbW6TvGT2BfSM
o6iSJqm9LIjsXhJj73WPb0QzPpleumgDTY7GfpJTRE3cSpGXD2xmNEwcnDWY
b0pBRD81em8Z48D99nIc3PufaHSPciEd5ZFEQY8CnFSjVorzMjXu/RQNEYOi
Nb58yfyMFayLTInJPB2xP3hCL9WtZMNZw8SghN1dcGsPm+cmcvoZRoSt8RYk
ZJ7e0GQswtwkDNmeW42aJlWTb2Zc/B6EoraILjc+2anY1kwxZimwqGnqrjPW
qk4ALmq5iJA3Ku5CDRo2lGvJU97AbWxvSVNdVeuNnxJaE66dbrWDaDhOUMIe
Kh+skWKm+TuqTKX+P8cKXVFnqFCHEJ0HoOkbtvHGmHqq2dkVDMRrdRtrfoxX
TKO39x/4BXo/si66zriKQSHz2Tv3QuSFF/64G/Gqpkk8t16pMuRiIi2scxpM
pAj/J2bCg8SN3asJzrsaiKAoTPybx4ym8pkBwldH5e9hBKK58djYB41Rq/s3
1rkRdy/poYVyGdqJSE7I22zM/IkgludsKlAieOnFlASLP4MVntA5UHcHYQpm
wvhdBS8GckwM425jZuV8u8g1HAgnR5zZctiR3vzniMXUUylew5WJa2appc3I
KjkmiyJrmKvG9os5GIWUS0geDVePXqf3wu6UywRqJWKlmHlU+/axpwsYQ5cY
u/HUMuLS6cB2m6RR7arrB7RhuSl0DouiLoPB604wSsxJOpll3yEDPG8OhqO0
1kYTaJbq9tqp/8UCG3cR9t9Me+9f6Ze0Fr2EtiCTG6CeU7sqVkUnMViM+qlH
qoxk9kDqNt2WJhh3eQ8BtDGhfAPWm16Ecy6B2fyFEcS/7/2yzEU0Pkbr5O4V
g95pCEW/W0dHgxhImmi21a6+JE9CNo3OS9S/EG7eRcDn+B2/thgZPrjBP3cQ
lPQJKSR9fpf7DKBhdT3O0qOCfW5n9JJL9SMKlHKK+jkWf85rrLB6ACOOjx8t
W5E6hUKR/p6igPxURHBMxNYC5l318ciVwYNoHZLBSfbA0lfNGXrXGLo20k0m
N1ude2ay8R8EB4DhCEFwm6xOIBzzAf5EU3bebi/xuctNcJce4JhCC9ayJGBw
DQ7YWQeMnUzcKnT7MR7+DuXhz23Jxs3a8aWlP/yBf7LmKKoPsmeTYC+rAxrV
fvE+NarK8XEG4RcdShdVFHnN3y/A35uzsJStcJHRy+idKYOX+Ypf9npPUfZ0
8iKpgqxHNThlbjxA21qefb1Ck0bxH1Exckmtb3nc/kRvBBdJU2hbawJRoTY0
pCYYiJb6Pxx/iVxDvr+nsR2z/NfhPy0JlyuT+lOnltJBxHMCW5x1FZ/KXpUQ
zJeyVHJbjYhGrNdU/FrpqoGxFHC7BWP8LBcUB5Cr44AvTV8Bc43iL9kGO8go
UZbAp0hvVlidguk+WhtSLCbwqIO1v3T2wpTQ/cGKKQQlPIBz5H10pFbKtti8
Ovp/2P+LUASHDnM0tKb4j0tKJB+gi3yIbwzPbDa16fWpeclQQ4qPFJxr9+8V
BpjlOa2KJ+O3N6ozslk4M7o1wwThHRIfoEuYyLXYG6+RReNW3eapORq+izmc
VKUbWsrWJdOCkBkg7DABp4XUu+d88aEve1AxKoAQo1rT9pf+KnanZ+NnNKr4
C7033bzIxMjMTjTn1KCPI8WVAyi3YNfcPjhjRsn/9XZaggX26HSOpZe5XC+C
IkmJkJTsoVnmDcmLxqpqO8N+TjQS9mi2ygbC1k/dKcbyaQaQjVdHuOa9XZHn
liM7vHZeCMnrrr7rwesRPGxfy3Ndtft4ZfyS/bZw6iuAOrc/BCjtp5dFUPTp
gu4FGGUUA/DORFY46nCM5EqxWG7IFfg1jDorxpjd2rQ8hakLVjVHTd4uDGAp
tIIncy7Zti3NVb4LuUwmRbPlNRfaklNx7EEQrC1kXSnbPRI5gOJDul2y8WJN
L+utr79nOARFVK1hvwbYi8ijdZvn57abyIGP+4miT/EWnQD+Cxovghxdz1xh
jm5ip9VAGKtR5jc2ahCvymwvgHvwU4bAjUdwkfAWO7iLtTk15oQODtXfhMuI
nUY05xp8sif6Wl/WEfDb1wSx+muw4WLKWXMIjQn1Zjw29oqJQaz6kNA+co5n
41F5nIN9VU0P555lHgLmY55p8ZN1N9+NZkrzgnhaF2pcpRAjfZ13/usC96CK
yK0MYoHk3Z0vlX1qSQv1EmVEqlCoXUrNXlXd4kJJvX9vjTjJ4fW40kGyLIzA
3+EYYk7LbNojAmE4qNQfiR3LvLTR0JTui7ft3e/69llm0KirddWvDD8qLnXl
aQNLe69CyG/LsvFJWDLYwoyeZHjDUPd44aZ2Ovt7nNAmEZ8Qvp9d6a/exrny
HmivW5gQF0zvehhNlj3a0w83S7Co/YIpZ0uvgkwBZWlpoeL1Plvub/LbKx4b
ap6eymWBTqHA9o6y7T5g+OwdyJQ6sahTGEnCmWO01LWTfRtxMz5wV0ZhmAWh
xQFFOjYmehpmVDsX8cujhBbCeBFfiVKQuP4ujtOvQsmFMd7KTNKJCSp8Az1H
jNEjgrAyQe2GOGqVpa/8jmGdFAjLlNuEWqx1AhtY3lvXZOlEsJqMhHW2E6jK
ocxYkuEbM3yKMkt1vqqZlYKV8nQ2t7kKYh86DSG8cattQrAAounHPOIx751u
gHFl4sHrZErx8gBQ7mG5ERmbtxbvWY7H9PVfr2rGosEaAa/8WyN0NIV3B2KM
8cTbRAVkCKESj0y6p94+XbnG/DENKXcEmG7BoVb96LUEySLbfmR4ZI3eCCB1
J8V8qIC/rANh7Uuqcnxgv7JmRg5ImmuQRZwUaUdWgod1RuvAD4blTboE1kFW
Updsw1TJSNgwqtu+c4OxwIFv7Cuqj4+UHx5L/4K1XeB5f0KKRfqr+dWGD8tu
mfNE8P5CLQcQ5VkOQ25voYOWt6IvuoQA9nK0g8QvabqFNNBJmMck8SFC0kys
hXk3xiLfbMOoBbqkgWOyGpxkjz9m2sqvyvspxn5i9mQ0RpEiipQfaoKDfRXG
jAWFMcFnhhExcena5EZM2jgplUX4yY3WsUqwpLj5Zb3N6MtEs12XZyJaw7EF
nXVfdJfwRT6ERRLa+Y1qsMnWsBRtr7EGwrUHW0z2oc09dEhByRisl4T+X/H1
26nm7uijxImIq1oxyrurRF9d8EseNIhC69qQqK6Tx1K9npPTITfzzS8qUMGf
xgZM93KrXZcgF/zrt4+kQ4ZVdKRhUva83dmy9M4EAU1OzDwdZ6XOV2cEgCrd
TFCpQPWVExNN1N7tAcxVNlYXWt9Ax/lcqAyK8UW6CTmgbUQRqxarWev+lJmO
Svif25luLosLDUOBng2j8NF7Zf+KBWpQPthAR4B7T6/M29qB/0yoqeVhIrwF
g4FQ+mWVG51ZHVnJTvWemge8IfJFRi+dF4iQgewiQmUkAwp3QSu87nz13Ar6
r2IKO+9tqIQyeD+G9Zc7onYjmwLFho7aVXcG1TMEPbEDSLZU9M4zRPnv9AiB
Rm/rbiK+f4eoIUDcW3yob57M5aO+MIuIEu+Ai7FtYVKSx2DyLuzGj3N39WGM
oOwgRaOTgC2q5ZDdja28WciaCDn8dPXGDndfpvKQPkLNEDeJhAhLNgR8ONOa
SnK1Je1KiZBUz0oU2yOEtoyWYpxZZDLYVA70DLotrC1NnI3S361BGOWMFNEt
uFTc31vI+sc30tnSfgzB/hx8n8IepSCSIjuqOUy5mg/oSF1MtOWrdpqgjb3m
Qp2AWyIknex1he3bNBXevhrxHElXQaFgRTWpVbBvPvMCUcqGPrlGpvHq1O+z
BOvVA4rc84mnGVcqYy88+Ni6e2mgzFkIWy0fpk134SgQccOh5/uE678uQeL9
s4rDoRdifuobfTCWWTXmgmDWtfLM6tajAMuHUT+KCEozUIuQh3BxpLcdV3Jy
QG5/A3mIwKtrV7GwmA3jaroipWWvzTA66Ls7mnF5+uJRRfZoHpV80WIjEean
fMEYQGEuxBykQu2l/Bssz7CiwIOdLji/pyVWPYcKJDxRoOKVGt7bI58sa91U
lyefzRCfYADpfbh4/bIyy2adw80VHD11FViYDZvBFIP+mu/7yzclc6eNrIK8
PsWcg77dcJ+WMtTE7ENxWu4p01TB7GYdFCG0F3PGm6dKf0kdXKVOwJKsbaba
v1ujsvrcASEUIpoagfLNPP1kJzVSOs0Ibpm/+5f6RZxl8DbI1pYS/hfGRDX+
mJJReS6BLqYPwzkFyUZeB+AcDzcZjdEbdrdtfu0OyDiStZ1IBjDYOAcZigNH
+ksD/0RK87I7ERWJ/fBseARu/ataQD+jSveKYnJF87eXotvQ1s89jQrVWTio
/FhAFSTPGOzWoZ5Pkj6SukEU9H+KjBhVWdWsiBTWJ2jDutZYawhRKBMhFi4o
DtdXHyD50WevKBBjP5DNaLYkb/ACEYEVwnpmziWQNze/TUsVAg8/odrUVcLR
uUcPfw/SrmAajejdDkKCaCjTVwaj6/Y436wqu/DCAL4rxbIlzfWzBMigWKpM
2qI366X7bVcSHjQRgJCsY27jaj7BfAuC3U8JetjaYrHzV+oJUw52Fr5/0ek0
m25rpp57WJRTkF9parymfFSEYEVMFJMgaatVJ5QacAI1jIGZtcrzKX63iocc
WyCRzMI4pZFnx7mmyGU3DGcgEKSiD6S0cid/kNI3t7WKKIoyhvQ7kuQsqrPb
m2i18rGSTH6k4q9IJzfN82hPaAbonyPAgRUGkSvWoI1/+aUfRFO7G1ECGEhi
7G2L7g1QL83IVoBfcIszUdv+fi7dU5or6HlTtO3YIm28bT+OepNhKfyHlb6E
e6CI0mCdRB38pxQKWPOHMGhvtY21CD1gxWj+BOPZmVHcOfwDawhfIi6oqwIf
6QS7321MB1+JvcYGQAqf8I2OKCvj7jAeNi+am+KmxuvLK7Gyb7575n1VryFn
IDfZihC0FJ+Z29J30TTPmOOLVNZct347Rp1k44/afUSV3+3QVPiJ81yoDefl
P6P8BB1qAEp3fvF179NQ9wcmA2hiTc/4zNMFP7TxOqN56YgTXUzbL/MSxbbV
NS159fvlnCJQgy0xU3VMcYDi2+eFJxmB7u3EmgLECyFfzSAPGiluYqAVyKEw
yPL3WdbGAbd5kPpCC7SLHbmXz1ePJiIgPC0nR5le48Ya3Xah6lCn5/u4xDcu
hlMBc82ug/CZJ1KKhDRF/XJ+ccvyG755rIMLxXs/NRFUJssDN+tf8mQ+CcIE
3alsu33C6uTeuyrc+Sv1KTUEZMf34p/mczErD99VeiU5CJ9/iDIBeYSKhHtr
ftRtcKFF5JdTUsv9101lUDgxHAyFDqn+Rj4TVVE1FUC12o0f0wenWwvXetsk
qZb2p5rJCCZkQK1KEMwQRyv1En2tTPRPeFDt1l1HdBGGyueRP9qRDigl4fjv
uGE+MYchszhWNkL/AnGVp5Oi+QJmKP3Cgafwq/6zZ57p59ISPQ5vN8EsgHYc
CK5ce7sJdMGCjFw2pkzXYVXC6Q7RjaWbh9CLNEbY+A54Bu/MUgmExPi6QxOX
NkRcWKMgndLnqzP7NyMKJn3Vmrbk2bx+lNjbNJP2SNyMQoGSS94KnRI8n1Vz
ua9RGdWr1KL1uWa/Uomlt5bcDriJ9pYEv3uFL791aHcuTuGJg5acm26fzpXW
5vDYjEMlmFC0P+v/Z/e3TwENJZVnafS8ggIsnCHHocdiUQivzlf1gtxguEO1
gOS0ARm4qSctOHJ3sO77n8EProy9u/2bN53/aswEXrHYodyDE6VdsNEitJk6
ink6opnp19WTfbyt+VvgUJXswiEgjr4008zwMFIOJq66QtbEoKpl36Q21PGW
zD0GEuWNMqvVAbIksUXTYhu0Rtn8LcHt2Sl8SqjOOpvRnCaMZil7MD4gkaC0
Sh0cQafhDgirnHxspzqEvplq0klkFhdhE9cVMOOOsiFBbT3oFrucwT6QACSU
NnzBp7qEFbjS3VXSd51ULIiUoFuXuvGh09qjX847SSmm0aj6NvPNCf/T/pKC
tZSbGYe0FXBbx0RS/DKS4GInTFAt/RHQdtlqPyRIonSy+2TfXwi4W+3WbVqA
yUA4JKyuVtRFufhTqYcT/jLetjj1uumMBwU7T6W/r46nk7TbE74AtRQGPppt
cwJZBuQYwcPyHBVVInF3zULzChMFpht5KpNekf4PoCMJaWA0ZLgMmUunbkXa
AAb0fMguRiuVcz+gFyV99e32BfNp02DbkdC9dRDWbJwQTIJ3Gj2ycHOhYHHZ
LNrM9D4hN1rnPm9LEqh/bS4Qbl5lFZbGuRdLGZ0Qnc+xyHtAYOZ77zG05Mfo
Tl7V4V0T9v4+kenRq6Jak4kn2JCh/Aztz9us79UNVcb9YtftUWL8UtRXD96n
0GBtesIE/cWn7Ym0zdEyqyeDiYtw0twUK4LKTlIGb1QJJlFI1VKzQUkqBJbg
HjnFntCsbYh7d/4hRDjwCuK5gH1ldSGvd195y34hvmb+oRJiOUYt4K8FJfeQ
MVwJwSpVK396QisBkuiAfKeT8JcbtUbMK/LrZB7Mli/Pw/Dk8snxQEhPw97b
nz2ShV2x4N/PIdJYnd1omvaTM88p/w72VmwgAct3ZSbvOHc1gt0mx3QjpImp
b66tDvhfWK27eBzLJ8eLTJ96UPhaRRtwrPixhdYoR8o/EpgwUbc1k0G+0Th2
9iw5G3F54cBpxZ6f8OBEwTM1I1YdKpv86AU28iNkMn6GAHi+3XTXEHSzmlug
AR1cSzUlJxxlnRfzNk9/+X+4QQDlPbvIFnzjJ+p1m0V5716wCRdmCbir2Sba
2+agQ3JLffJHQ/qyCZ1x7SbT4VVE5KzSNsAQ2gJ/Anu4v6G6/X+2hvGIMkjG
rmsGRMbvkxPjJmPrYwGsJjBOZhrt+oLOf3/+Yz/Fa1O1yU8RGCBOv4PHaN9f
p2mpwkjnOBFPMc3xWs1jPzchQdVpmN++2DRoRVxwcwPzI7fl75wxvUArgSfj
HgBvANHoIJI1Pbhmgr7KzP/bwgoO8btWVUWr5bdIrAocrglD1WWHpFnWQAlQ
cKXPWe+RI8b8CXkW4XEnbDwP0qTLgMZRPKrWL89Lg4n6fXYR+Sxyl/xilC4T
bcQAYW1tiJmzyj4mq4fulEEyQAmHncP3oEVrd/fn5bl+l5CxvefPrUushFoZ
Fyf5xEF69RvNuNC/EF6aWvGc0KRwAWHEJfs6DKnvFpUrAVObKd8iGykAtbbm
3IoXmrPVIKzTF3TjFS4yRK5IGav5m+qh4pZgod9XDqx4nwX8gRa/dkb+zrAa
JIcVlbE6dA+kQde2hdiaAVfJ/phtXCouaj5dectH2UvzEhWaClP9unv+SIYS
KGC0nbHuTMq3fgOasKivjON6aIbeSTCRz1bDXgKmAHsBgpbLDRnhA0G+zK0Z
mr5O41qcntXwVfrD0duEAV+yiky81tJxukUloCyz5jj7n2YYD5Tu8hDXEa0S
lfe/WykyIobDO2RP7JO51G4nnrcfG7FHytpnyZQbL44mHvMES8kWQpgRyjV+
OVaWjY9x9W/w5ofZmx0cYV9qke4JTl5HZOdEctz/btwiESPRp5Qgcy+KM03L
ott8kbkZI2YPXUnw5Ag2pGbxEV1Uvhq8w+IY3jjrI+GaWsbYDrryrUvTeXeK
GizkgqDIvMNMJ1yXzPZ09QjKq3K1lDRVyxEJJOaY/AtNinpVcGV+jsF3VZLe
S13Zzv4VJg4nkj3UdUNL28S0pKLDeKC7hkxVLiUEAwMW/QkqRmr9aAopCtg+
YX6sRitWjaDPOOvrvrtUdyXcheeQ53z7lijH4rG+l/fEKUTPGZzbwN0s+GZq
Hn2G5r/ZP5S0pLAZIsDUrjlrRc9wjBxtsKxIH8IOR307pldVBrY55HntZsaG
4TGk1LwhLgc/RfOFTvyO7AV5Lu42kgDz1DRXhIW21fTI04AuM96mz8uOTHXi
Fr80csyZClUP4aDoRtk1eoLfD4BIk28IRRA/9F3jeHz8On5VICvJaPQ6CpaW
yfdvFn7LLM13iMwQBVEw4lYSuGUlC5YUx+iLWpDVM6wiSbzs9xq+FVueSOXg
x7tNBg92Rs5AlFIDUbhpsQrBy/GWjsVg/VmqPVpD0yo+/SlSAnCd+HwN1kI1
KeGy6yck0Dnzlb9nzK6bksg2GaCEZ0/EXMrPfQOuh8oG6xdLxwmKS1yRAY2/
B8FS9/4y1mI5QtXrTphkl6UvdTOFcmVKs3CMzm7wXZzQ9b+GfPBWX8WhMlTK
WwZro59xtQCxlsdJQ0JgOlwDcQlVFISYp6j8LgncgbpeLM8p53uGPz3ryZM9
e+HWBWAnY4ilfZNCeB3FS7k6KF6Kh5D3b3FhS44lMkZgH4YY8vyx8gJYOmTj
g+l2H/TrqMLd3e3hRlL+mVx+7R7gWQRJMiqi7JpbWcBrZYSGwWM0uUbSgcqI
5VZhb9jlZSkG1yKLOW/g25MC3T47+dgosKA1ns20Gcp+jdVm4+bda0/bwcm1
WOTshYitLiSWGyNjjlBbq6g5NZ0YYcwelFdiv9T9qTAWviO6YX7wmih3UNuJ
rsDVar3hzfAexhei7g/2oN4/2/H86+B169skixSK7uA6rXLxxMMRE3eR8ds4
uPdnbyNU6gL+j/wndDXBPyBaECcQyLAkzkqVAeMdcovv1C1n5e0uQyT641ub
g4MoCdGYpedrF70muwtpfBKJMLHl/evTp49WMqoQuDIkZXXu9Jn2RcfgTtww
Y0+ShZvINegFHQhF4XEjYPe3RPiZ3sOgco5GCQfiIxESYQ0IpAEBPDeAWM2r
mo589ZrVCKsptUjBPav3iDnyh7VnASRXTa/LZi0LAKKJ1B/iZh9BCBgg8AXY
EOtN+dOP0h5BLkpKs2Y2wuX7iW64muu6ma1v/irThy4uQaZ/RX5zQz4lUxdN
MVB5vLoFZwB0I7Sd0Wwx2Rx/MfH7r5VfFQvWHtodI2bDdU7TgQHwyYAkoxFY
CJ+4Ca6qaehjg8ekLvYslL5OvArd6IwNc/d1y68hRgvUV8EG7cOKp9EHYp0h
N9R2T6zPGeZL/LFS7Se1BlICujpEB1TLzc5x8XfQ525yTgfDJPqWuUaSTPgU
Ra87OqMEUaZLZkeFT854RmI2PBJqt5bx04Es+pjobAd7cOIOaDa+fa9YDAzY
VokGjn2/Ef7EAHtrrKtb6VEHQ6XCFADlSmFHKtpIaGR+vceOaA/B2LQVdwmC
TYkNrbeX7NTdGMLTB/gPQA+enZs3+zL16i91e7Wyu2eoseLG84WVOBUv6EEv
Z1Wl5zzOdiXkd9OlL0TfD7kK2iOf3vWBSppBjs4po6Bl48ghq6cBT2AGp68u
hJVYkJRJTnjZ+aSpdi861qbFwTSDYDpQs1aW/le6/eJBXRu50EaXAG0XoIUM
O6zRmaXgucvGh2U8boXyhkZZ+HqB3LYvWoF7SVOWizXBOwdMyvajSOdnFduT
0GLWs7lFof4+1lzzIdjMxqCDliTlXSGY5/wBySM/oRLx0V2rz4gx90szQbfl
ljwRFU80RxuuzQHhYwt2A0gNXa0dwj1trrc5k96ty9XDM4iZf94Z+W8VBSnI
eeybDuMT/NDN4AhwR/pU+WJnMtZ/qutqvKJqnP007uewIZpun/zb29MImJvw
Fay01rt4fdWB9+FgnqC6F+Bb0qHfzaFOLa9A1Lqly2r00kvOB8nuDjneaxRn
k717A3mQcnkTW7dXZHSbVC3ngwBzmXivTzdAr+5a0HZE4eeymbD9kRLxKE6f
i1S0ClluLwCOIFx4rnZKViMC4Nn1SZDgXaEfqX69iV6eOQE5wfzdD/rN5AkC
UPSdrnNVD8D2GtYsjW0rAVuqySsIGn1EzNRiwiTsRp9/LMTqP5ooJ4P0WWnR
J31D6m9i3vLPHz77H51wG57FYRdmMoLP36bKl3u6xoYWFFThdxWMN4Fmld6Y
YJOhjQFWibRVXKEAeZQat6Q9i5oaZ4fDvuet1DSaZXPsnw4I6uKi9fKWSSLl
D1AVelZ0RoaeA3nQZUzvkSpOdMdsTVZK0b9yx7I3geo+DdmV6qnECSoOCNwN
Qcu9isGrLUNEgVcSOnqbYn51pC5Y6ToZyHzZWaGyxn1YPDob83MgVjrmfPYd
xhppI2aU6IJIi1042svEuGRGJz4xr7tXTuSNcOkU/A1aYe6nnq69e0UsaNEu
I1BlnfIeDORZvD/7WGvw0IDzgBVD/1L5UeiwFTbq+YzY/FI3xRP3og+sBrVu
fBwAPLGsYfO1eLVhuXGEQsJnGherEa0welvtnGMoQ1HShbjIDBbmq61KfA63
MwMaAQj3v2udg0Abc11tlALyDMek7SVmA2JMXSixwnHWIn08s0g+Ylz+DoFg
LVBWNgYzNcd1mqIluhJVyIDKWdBtHK+Aw22/h4hlbQBalJ5m8ZJYMA6OC9wa
tFpCvSuEBDuZTuU14S+/RpSjaW0QgQtVSwy4+AZziJBj3rBZVSopABRfJbVb
+tAoo+2g0nl1w6OLOQbHs4Mzdo6bReGp2FlavNAfcNuJKSVLNTD8JygDADf9
ESFZdOYOLmhdUPkYG3uqedzXXkebMMeRNAgEtu2o0nCrQje6h3H+jMUn/bz9
LjIsPiyXqwNIW2/sk0wVMPPXFzKfSWGMsmuhcVaXXRgyM31zcUpi5C/6MlfY
108HjTVJp4UNMfNvP2pNEFSNGE6c+JtIRyfJfbIcOA8b7fev/XxVgaXw1oJG
DbwScjeZ99wKE+zZCA8W1eMT3baLSglEFbWukxv33bnmj2H5a3qcjKmpwp4Q
MMoWIyjWXk9cYmK9BJNx75NYJdOtbZ9WOIimleoGM243yQnF4bMMCz5UwHfN
5R6c/OICCrDBkk34NHXokfvo475lBSh0WSZRTak6EelW1qKK3j5lilJSPXaC
04fmFihK8nb9q5hjR4h0P0Ex8GQb+NPe9wNnQPazCzjS/k0oXxJ3OZME03Ov
brF4tJSQ2qgMS6epiKfHICIMhQqIBlXwbTiMUx6tg32SjfcT5KBjbciHHLBv
9pKZBhPskd4d3wrl8rSCueCEMywXBFfGwwz1wSlQAna8B8xS6N7+RyTtG8Ww
4ohjI9xv+j94bB0xsWkgGcJeBakVtFME6q4OkIVEfGH8XZ+I7LF2nxjl4/t2
uvK3sKzJchNEM5XKNkpDaIhSjhf9MtJR/tFeaN4q9Tr6XbHB2YX9QjzvxBpg
XiDnlyXcGJ09ew43d3RnZHXYtgVfLciaHUFAoU1Kl2/bucm3+dZsIAntNnzl
Lc7ec5vxKsTVovP3//k6pm15ztZUItNyYRHdaWbBj8bDl0PP+lze8MpKTo6i
lORz81wgsip45Fxhwh9kjFVmVHkTipXwhvLnyDCm3D0xRPL6zxl9iUWyHKdA
nhoTkbjnSwjNbBkrRaA69Jjho43N2mLOlEdHpke/f49aEe8Ca5nHlDGncumT
VoxJkrbjNuvV9d4L01HIVVziiWV6h11VFKLR1aaTDkuhgivMBKYBl2oR1YqU
RKqTTViQNdXYjkNGncDQsp18cAp5SUY0WIIfg1GwP4gDNxTuaR5r1okNuqYl
/608UfL6lzWoP9E3QC9dMB5ifNaTo8w5CPQ6SPKFfnHmkEiw1RxYikrG/fn0
9iQiYEgen0vT1hCTAm9Z6zCjDLS6JjOdQh+e0OGMJFHP8eAJ/2uO2xP28ji6
afCS6hE0CYmYOhXI7sJT6krc4eGx7AXNWyhAjbMno6JqFzn//op+XWEcbLCw
L2AGFPGQCkQD9xxlBL9uQj2JBVl4hHmnnvgVZpRuQ1rMTmBN6iOq+TYBgabi
gfvlnSkiyv5SpXwMl71THCbnvLtDYeLmi0e7C7mclJRyvOBC+C134Mp9Qd0r
GLEvY8sSLR3RvDtIciq8EtFWMRBe/ALirBpLM4dIc1rdqeJfK+A9DSIOPGX0
2PriSFgI9SFv4I0NIhS4WkWesNteTStQ4ywEbkfwKFTruQwIPjbAAgy+64lf
XfqqfnMmmdQV8vDcg+M6Cp1eUOzbQZguVwZHVJDEh8wPioWKJJdBjJijm/nk
MEKI4syriWesRrTpLTaKzG2VkF71K6a1PSDfQPobM6n9V+5Sv871ffFbd4Nc
yv2hAD4FHLdJ7cXETTyg3gZQ4/9nsFKMpNor5gY/LI3XHJVhu+l4znAmSVA8
KFOZFTc6/cwBrncCWq8NARjLovn9j0bUjw8uUltgHrU/N7yH3D1C2fx68zSc
Fy3w45nI4Te/O6vEUBGtmoaGL/a/18OGvygcn4yu845tfoxG48af9CsQ/cZq
KYphGJo2SEXjgPbH4mLZ6IS/1PHfPzzNyO7uviZ3qewd9OBxm++rr5ghrZVZ
OgdrM4SU4XApL2+69dgjc2h6w1thol2UDnTcWp8+6uTlU7M34jHhgDz851ZE
/qhktabE2MDOWeWbUewU7qkqoNmPOKwLoxJ3A1PcVF2IoT9HjbGAdpwG08uy
Xv4M3SurZAsReYafPKf4tj322LeWTB/brZBe6/kEv0LmxbWYb762kGmYc05H
b95fMn6KycQyps4rZ5gRNk7rIGzXS0bK+7G8o+ctynwQZF43nvCIf4aYRdBl
3biQfQ/VLl/lXqt1v+BqVuwgI2CFwrM2QMXIgQ9Xdn5TOBpFLANX/2073G5S
LuYZqdq5TreqH+jPg34UselI2vjrILIa3Zw3ikG2puSqubfIxJYuOcOkP2F8
82ArMk3JBKD5AAsXjjWzI/xF2yJN+Wx4nJ+TqbY7vjH7mc8mNxoI1R8Neo5g
K7pF0ClkRsdqRlSbfJpLmL+o6M2CkNI6kYbmFtOUhp3lrv6vWp/crkuIuB8E
ZyBrI1eyq5arnoK+/aZvwXgIMt1cdL3v0ef/Fh6qDpIIeD49uL4x+7ugJRQy
l0SmR95SOfwmvK8db9w45vJGTLcecgihmTlOuyH3hTjXap4Bkgxqs/kuOglx
JFYD88rgg80j7sBFi5aXdhrD/gW4rgc6m4ubzl0/A78EHfslIKsRwB+Alu7d
rBlHBRniUR0PdLemnoHj6NnVMISBmdnFN6S45SEY4xpsmb0si+FQykQ57Rdu
raX3oWsV+bDRm9PxtFfYK6e9F4ehXNKaeNv+tmBFYP93kX+Kg4Xw9WbV6EEO
1wMMKKjWrfTfHdX8/COvh+HmyXSMDctQaaOxcnbOKGg8HWcHTl6Pim1Xi5Fs
xeNujxhVFL86byQcOsIjKnfvkl6DALUWwH/z1X3EIFXeTnlc/SEwbgM70Lik
sScheZWC5Z3oYIOhkL5rvOQ514tL7YPxluvaG408eloRQ5EiuKlgMCtw97ez
bjaH8TF5LaImuJNq3PzFNuPAWzxpp7WhkUT+u10zRsK5G8nF99Atj/acZ9gK
AAHKJJwBWVybX5W0d2wH5J33b6UEScuubjH33x2Y4eXBsUOTXnd8kq2dfAbd
7sXVjNGYZH5hTSHHebBMlj/gfI1bkpnnp61EPNZOWB0DmsB+N5DpSFhuTbOf
Vpe1LgQIp/7KgqiWU64qAcb4z2rb3dB2WaWnyfXbJr/vz6RnIC4VQSLAg2Lv
aoBx5WP2hxRFc056mOLXIBtxD6QohfiqKW6Jma085WxSNpy9XwnWjNSw752f
OxI53BCRUlxwVBelmw4Iig24Yac7KXiN56G8pW0aDl0NXv1ypQvA0c0wrg0m
7Wh65lqd8nY+YOal2To8eiH2ORG7RTd5vO1rzZXfUAyoMEGurMQHtlVsjTAU
zDpYhMXWWE+PEBtZeJb73BsbOy4mg420G8lDkkE3axNyA78EuASrhkyRLLoP
RIiwXhnAWGZrtuB93CkFo91EMNP4bjSWUjhLkTM7+pvYLJmNs6mNHuzh3/eQ
EnYRSklUpoPhGGAPcY9x95M7n2HAHkVIsGMdPVvGlYUWqFCFQNHEi22yMO95
KFvPSjvw0RvqdNxXE/op4rGXtooHM2FrA/AaFIlNKa7oiSyQEGEt1olVRHZO
1i10akJmoOtg19GeEIrcm7fVMo+atmyeEvOsDCNQmDvtobp82WsL+B6gwx3A
KOa74xP7Z5Hy4JINtLsndVrN9fLLHi2uINfTr8MBSVRbVum7iDEKz6yQLcn2
z3+8LU5XM397UvvEGfmKCe3ZWS80rYwOhnpTQwbLCpqTJdQn70HUCtdwr3Qr
RnSeltcpX4EvV8PuBkgGaKPfUDb4KodELCGX36Dd2CNBmvpIHwzRH9osLI3Q
CUPXz/xD5OU0GtgNvdaxlgeg9C6A/k7xLc36c4u94UL2kE+OFwydMUxOAGYC
JnBl+lQVxJK7iLINWbQRBD4oF88HB0sdQOu/vBuSTmwTF35SQ+uuHMgjnon3
Ycux3MaI4RjKHidftxAN1MmozfNqhnIjikNEn1dbAke3nGfcFck2VUSe+CS3
d2QomaFyfrwYmCoKeQQ4otaXIoYqsI0qXZU+hOZv0/d0ChRiKG/Zi2UVbTxc
YFWbihQHE4H9/VGImNt0YQa/OziyqQzX29Olgw8IZh25j7poJZxhBHAjO+xh
7IqcRjewYVGj1y1lgdGMaXMBF7L/vnG+1ax1sW2MmO8tRqCshH1kMvakQiFb
8wbJ0hAE+qybuQJQ77vBiQaDDG9c8LG+Vi7anOkiL8OnfI3fKQfIv4a5gdSU
v60SWzTRqFEbgo9TF6ncGu7qrPZ0gQkzHInKfhTeRijPqgWN0TJTKi8cL3Jm
6FpAv+pkJtxicCWB30ybEy3F96gxyLNXhzEXlnlpGiSjU3z8a+NI2mzoZXjY
lqpkVS5gmmrxLKPL3tW60jsElVoU7gKxDFVdGJ41hCLU2RXs3X0u2WzoMo9R
TsBVqmzQxo5fHePOrta1HAavjT7KVwmEVUX6lqEZcPB0I9dMg4ledBe8bH6X
keGk797lll5vskR+O1oTjFBTG6enO8OBmHPuipndy/qb/+DBfLdWov61ryOj
hMcYD8zFAj3viEy1K4iHNKzUv+kZ7XPYZVrJVwecntM+M+5Cr6L8XpKd7NS/
V8WinCTdiiE2bR4u1bvUos/N1UCUnGglc7DEVY3vC30NOOReCLrhZVNumFbr
9o4l9Wc4N3mC7IXEs2aZDkZV9xhvqwaGDmT6iTrUUfYiXWdyU4OT3nLpGU1V
bL3zracmNqcBjxtIj9g9mgQkkUrmYpYQAT/H6ZoIZ+3P8nhsanCcx/LsXAaa
Fs1f8obiVQw/s+J+Ip7eAGWFs1v6c40r/aEbk/czTyRBA4jhsQndccC95lZB
jxuVECq8hW2K5KlYylk9TNZTOCu6gjQemPW5fw+XXZ7IxB1yyQr5eITP31di
4giPKoayQStQ43K3f9pjkVOn9BWZjEa9s8J/hAu3resqO57InsmQGTlGMJYS
MsxGp8MOnHZ7BH/ZOq5fCPROxLjI0LqqpqA37boq9gq4SQdP9jNQdOJe8HAF
6zRQKyHWXsfgI1I6xEh8NDWpzf4WixkFem98CG/b38mLVu7V2qCIrB1GPEBo
hWF6qPJl4kpDryyDiVQlcNUDbrH2DjVUgKO0LKOgsksOvFboxBLxB7w3D5OG
HsWVDXZ0ARqK5Dau5uR+z2wzbdRMGlnX1HB1fbT4yDRnUZzUmiLhnGWb+WUY
PB+Iw3JyDazPe1eMTroFXQeCGuzPbHZs/z00OHLrEhEhxa7u2BaJek5tdjfq
Er5QNzddxS6HWu6qV/2kgXc8hGjOw618M+cnzNiDe9opJUG5LcmmeJk0bUN4
50hfM2k4wjZpCVrhXQjxycEV4RJHPevdzdMgKLWx7JPxojDFMnLFfa76n4cx
FhVXWoVr8TPBNXUvMB0nxGoMEoKdgLxEuMw8ONfqSxaKye9YA/LyODvbwHV4
/nQtC1mKEmZclwxvzb/nCIzUvLQ6vKCj3CznVoImXBn3CE8n35a7qZAR2xFt
c5bzgEbkmtKPkHUUtRANaQTERRQ6QsqI/gV8+9Qsi0gAW+YaQVlCgVdgXkbp
roMNm4aE6AmmavMtFbTI9oMgJXRWV6Jn/22UOEOcRMGPOyFbs5aW3tOsOvjp
uYl4XhXiKlYnwA0pBpEuLAQt0PTMgzF7i2UsKJ+njxEE7Npn96M8SI5MT5qT
Rs3AHElolfjrIWfVUJOkLB7/yLI4JNqE3FemYouCuIewC6v2/CC4MCFrswwX
58aFZmfKK84RtDpr+EOLMmQtZAoBwRjR0DbfJiIiPH1GOIpkj3v6WGgG8zlh
W4fCY/kgILF4sV9O2DjSRhKSfo28jqjmk1R1xIdjwXs+SCGjqiFbdTu8fk6T
RwCNXV4296s5nYAYYUk0UtySOK/D7N4hgCVa4THrw1Ms9b7sgbUZNbUesZQr
/zKsH0rzYnjzsRb1eYFjNPL4SCmXBtYGp3slg+/cs5Aw7EqbGhtu++amgmDD
DTs1LTuX3Ry/f9XdrRlpQgY2AQzmwJ0xbzAAv6cHkGOTKYcDUHsWTqJvkSbs
HW3cNo52JiIKaIP2f34VmBiKX2Rh6F+e5wVKDX83qUiBR1vo8moHAsDkYnuJ
37kpbuMKX3PNStX4jnClRO96tluK/b+mDPpYyTcjqnCxuzAuUSU5b/ByYBhm
2om+LPE8+memDno/ozNCWwPFIkN3UaoNPSEkENbioOXFy4UwuPSw7lFgaHkD
87KHXjNMqe2Yg8sYm73S6D/pu3svBdPlK9DOWBKL4mO09Da4Im3J0Nzi/F3M
dTLtvYnx+g3jGSVr9CbNqSiwpMPm+RY05lbPhO1ZxYuDBrbKAL4jip8dD9EN
frXzMFU5tylbfDQQrAek7NWM3XxlVUhxiy1gZva8eAEVAztblYUiFsRdT+vV
7qUyuRGJWuUAf8+6GBWgpckawyugaA23jfhrIsU4cFkbmvDmL7kisKAfSN5d
2Yfcxch+/HM9H/NeghGKyRn1kkNPA3fALssTp9zNSEgllY/4ml+eS8xjcFqz
jc4QNx20Ii3WEChRUWeLMm9wMZu1J1I5KWCUDMvaohT2SutFYN8mNsKuAqE0
Q1XoaTEQ0jlIC6NP1Kpm1vsPOIdNcHu9IsgFEsyH03MVlhXLTPvMfOPBZ8l1
FVRN5Bn38xXC5+iLaE9WYjdDJFdiQUCT+OM9HNqnyoyxPDFm/NfCiSusUw4q
FvemJSBRTEGr77STnri5IJThqaubhXdI5LURn+c8e0XFfegzkyWQ0jMqeceF
fX5XArz+KZL3Lv+BTh2EplsIzBfk4JAzdQQXPS8Ix0DgjWl+ihZ4aG8dbmXK
7YMgq/9MmtR/NV07uhb3vfAIQwiEOteeOM17sA5i8lUcrZ3pzsSNnrxRcN+9
AylKpB7XglgdoHXSbHz4rSaTGjimfwxsU8KtuL6QWKThNcHHrN0obkHowWw8
rFf+/rvqhG5iWXGyO+XBP5S1IyTpUS0g+3dTcnnhOF8x2mN4iaUHKHvweo3V
5Nujps+SRs2uX9Zf0UxYIxTPom2j455zwdpgZ/YoaHmPcWzkqc1d3Czzx9PF
5Ks9ePnAIk0+znyw2cECvvfAir1hLNV3UDww2UyPjFEeupSIAifrGgyUWQ/8
8ybFfsyl6tCbL1WKHGfQEO/qIOdSdPvR76NtqXEBXYsnN0lr+735BZ0PKaaB
S6QLXb8VItb7hJdRRqNBLFAI4oSLfF2jyCCkcF1MNebH7Lqdgp0WbWjivfJC
Hw+u42ezzqaM4f89lbhvYIFRmSioCpmcPl1pn/gNdDSPPASAJtoIxv2+qfgd
1v6n7mrUO7CDjwpDINiDugbpBtMRdMDhjctW3UkwuNVZoKLO3hfXAIcXm08d
7mmqFadXbPIb6F4s/n3a+vtL0VFv1P5UchqbqK94vGIzeilIy1gqsH/C7fRL
bdqUc8arE5KBNS4JMQQj2QJkD1MuM0dGJPfqQMI7ojwRKrxxl66xFg0OVoVL
dvK1vUyOYy4OrnUuVuZbEqr6LSZsAW5yNg2ri7EeuMIDpdgSbLjZa7eiYc5w
ytuzIztgJk9kylWnHXVGGmYVm8CXBf3kpqH6+Q9bKAAh2us5ZmtucBnXm7CB
69ifug2sfhGW66Xw3O7dqpG/mItVdaU07XeIq7EWYGbFkrykDqSX7D3OGHgh
HFXo6+rCv7gd9ChvpRDxgxZWjqVwm2tmjWBOntDJqkxnW2iVXnEksL3Wfarf
HG/9+6ZVVlHFkVEEQfpSmFNuJTSmq6IXxUboODWNVn11+KWIoqIrbfKU9JAO
cCvL/a9SdqMj303WA36EiJl9RCQ1MYYF/APvMRjnsczgb81Jpwn0O8reLlfz
4q+Vim1M/uQz8vi5wbGPxoMjUQnXk61bwlTirdwMgSZcetKw8h9udWpA6rOm
95bRYWn+zvVISc2sZ2p0luPH0qsN3HIphanbZO0vy0WKKV0PqPGOB9w6RWG6
JyKCOj9HYhF1wGgC1eR9gd+7y2iYbbmNTsV9bNNh8Q1b05/DzW/0Fdba5GPz
oJCWuxT+uV9qRjMnFUGA/LfbMyGiPiq4DSfI8kZiYyGt6ghBWNvcDG1HNAxQ
N6UjujK09wnUuPLVKswFRU0NQz3pVZvCRSrkAPB4DUE/eP4L+Yxr7zOv/N0z
CVhcV0a+kB1Izv2l+gQvuygIIBO498UcpzZWDmPvaAddHU7zc5jHe285s6E8
4dkB6eZAe3m9OLtAZw6qcnk2UVB2oG2UVfURGsrZteTNB7gHiNxKY2sBcEI1
5SRMimG354RvPr6vIuOwd9zuSdeZKNk5EmN5G3SER13wag7hAb5chwihXs2r
X2fmp/MqKY+66wTKn7giKFC+FXtiJW6qO/Zt5kobXy9z75U7zRIvXwiFMUez
2Mwk5OsNYrhIFE72OLvcHOCwrlGjdbgZe8LbyRLo7KaUtbiFOpXXymBubz4w
w16qjOnWPYWPRw+CovF999xidbM34X34AU9L93FBk2DKXFkY4Y9E+Ljfllor
mW3Dz7iK/AN8PjrWRxZQo5KR4wtlYiTVZq0YzWpvbXxQq2OeCMrs9olavjD/
nw9MkJZvuRjD80MjzDi4Lx4eJypakIhEQVfUNV/3j6JgnBkxIgaTGI2HZm8Q
NEaAR3w/eURBpfMEWiQG7ZlEfr2MCnDiQS3mWOgQgNcoReNnpLfg8e22TqVy
SCvjHYLyo/9lbljjjqvbaPKNqarB7kd7erH2VIu3q082f/h/mlgc84cykUJ3
9xIdMRmmDzCxT5hvrEeoHOwoDYifCgn/8Kpxl7pApBL+mUC0zVgafsjexak0
7OOGOW3SDSrs8nnEGpjlc7g24rBXiDIowviDduCyu0CY8TKCMCzTjhGZyJsI
Ypa8aMwtVyZVDaoyTYx2aE2g2JeoQSl8It9tGFkxXBQpQH9EzlYmPbj9EDtx
CKcvwi4bB5I8pvlQwBtgoQzDfb+Y482QfP6BBIBTlAK00wrvNa5gqMdky+cY
o6hasLLK6R19DsyC7WJpB2ZBeTOPFC8lCV5ukKlLI6ga6/ovrz6iIDJCwdYk
scOne7dJbqfMsiN7wk5s3vMZIhGut8PnN9BcCONgsFMa+SlAL4sY5ePs7xn2
Xy9EVIQyYP5peynVWJQsdNE/T6n5K7VLepVl30EKms/PszHnZn28kuITB0If
/SeYInYVLngZkuF0rgBsvy97AV1mmQschpTa2iwAXCU1GIpvom2G4Dip/gfn
tGYIXoCyS3ITMkSrySOUki+YKbvvz2kYDT+S9n1A4fexHbzs0HEozoHcS0La
xj+zkizJTd45RNZoXjs3Qv+STHVnQMX/Y1bZQgHxmiZlCZm1hjtK88TQ/j8K
LJsXK5DA0WUBD7xALYwJUPskzQaI/skqNP6UFzLRPVn38xmceazanaAVRhLy
+3EvVqjWXu8sjyw3rWtzuKsjE5nITLiuOT727iD7CneqplUBAIwyGISuWoJO
E9PSFPuJCY558txG/Q3jScipue6+miOmFJbsN4bKiGYKPJwFufSTR9U1GgMz
GG+T87Po6PMnuGseYD5OsPlekNAUBAQi02YCOeN6QR3zCXWqEkWHU2wB5ip+
0B3x+lblDFMouGp6VQA2Mh5Ed0HnkTisVKIuR6AZLGQN8/H+4TtAmCpBc1S+
ocq90AKM6he9jiuwyjJovlGFZz0ohae/NCrESzN6RUSIqD/BquP10f4tWWGl
Ha6H2ToAcQsbBLC6n9lmOXKN/X/T33ZWQ7mu4G+0JGSLAYzakgUR5niOWNw7
l9DENT9SDz1KSW/JKGMsAY3hy8o8HcJiHIP7KADl0fXJ0OmQ2oTDA+6irN73
NHJaV3tQaA0JKpuJXii8RaYGntioF/f9C1r0yjeikZY+ITEWaHkCWwo5FAJE
bRL+9gaf2yKsk6XFgEZ3i2W6iVhJS4csLzQvfmD8cGknGPBXuMQWHgFkxDhq
X+aQxI2fTzmnzdfqLFZCR0siU+0fICLmJh0X0B6cK92lRS+sFTTDFBVu1/SP
hfjnRL2n/kQoxFRn//nwkDmFd4wzosGX7ED1EzJqQGW+SajR9d+vSRrInW21
RSEO6f9BnEl7a9vVksLtJfKHQoAFQE/hEuX73L8PXkm8AW3pdbOajPLIBsCd
vdyfMy2HVjfP5fWFcGjUyhf0YBuVNnhrMFVgvOP2+Y8JaKLKO3E3mw/V+f/s
6Rq8Jq5NGeUeI1UCW+McE60+9cD9hWq0qa46v7wsMa3KB4PMFAz+Nou0jnQI
fFhc0pjHOOTAYQL363NO8wZVi44ddIj/wHGIZX5g0oguosmgyle1BbCHR+Vi
e1c4lGW1KTiwCOHklh9g5/ctgc67zljy7hZGQI/LUNT3MSzkoSaKPUpChmpO
r2mvXoRc3SoDsQL93nMxVt/I12PE6mQ/dHvK0rXj0LxVNVqzoQTTeuEmj+Vl
KiYOpHRS6xNOxgOqxar7jLQjngBu/Q8k58n141xheU6/7V2qq2JO0oJ7JZH2
TAWx205JPqZjWC4mxMcZ1Bm9OmdOh+Uezr7qYd1m01/7CGo1iGSSuzuVym1N
jmiMeAVjhiuhES9NNrto5lOWpFe42pGGczv1thknpup/PZaS52ehfehbienW
Y0u7O7zI5EDdIDrcr995X8wuRPCrBGoUvWWLKWtEiffzvQET2ntFRDgnTpzl
Ia4B4McCY0yA+Nj+Ux5vCekgkDohHVU7W5AMYrNGJGvjEaBl3oiG6C+sm8+f
VW2PfPkQGE4rmexvNxdFQZVIMDWwX9RK+Ue1OEgInxhj8PBqfm6oqNy7/cpM
2T9/pIXCtlq+mx7C65RhmSaSOMmxvLLcD6dXjTSDgQ/kSlIz4JSE45bZRv8E
6vcctLs/x/u/EqZ2Jf/loEpkYuTvZRS3tIxGNwORxy8GbNpYgKcGSU4DIqpT
ZtY0+gXyR7bTAv6k8Z0BGgCN66aGGmTq2sHNUBdlSii1xVCy32DRePQTXGCD
u5SfVzk8zH9WG1x+zHbjzx9N/Iq/Sk96GiwkKJn0HOTSMIS4Y1leSfsO22gw
HqK1RkIZg5H3L9Fi+CrXHO2eca1VzWlQ9wEJXL6bz9Juo5jhKZJcrhK0TV44
y60DqupZeQ4kFTSSbfah0yi0c8qsXS6WxfPyp4cD0RM1X1iU9QeOzSvrkHM0
GZSq2svOFsMkg38/7IR0/bUXSFHfeg1SLVRw9em86vvThNPTvwvHseit4bT9
mz03oU+kTPvNEyiFiqhqe1EVNUzDeSn1hMCU00Tci9pFfK1SzmoMMiSPnJ3p
tFiAT7da+DwyEsmF3KAY49Hon4OqeuWGpOJbFla9mF26XKgehLw/efM9u0Af
Ru38Iyc10PIKBoUwzg6PXvVdYTLD+PUYxmGCk3PxG552YvNsUKZkgceFacf8
BCBZYXFkqxy+bjvVb8P85ZX5E9aiVYQj+toMnmbHbGlwXTemW1EzoWCdkZxX
rDBmP5GfCEeUCMoXMI+P6SV4h8l77tTmla/6SPO+OGP3gIPXj7bChT45BkNp
exQE3ORbohXmVUDbWhsPyTBFsa8AhbWfrBVE6Ab5dLxsRyFdoNHYhfqwfLl7
QnvRgluljDi8OdoiWPzAj6tq6QpFx9Cf6AIYRtsChzQkX7LhLUuoevS7Cn+v
Gqyxi8NZ9C1JD3hYveq3oWtTaXsILgBqmQToDeO/5V78wQtkqU+YHLO1lau8
Z1gfCPw7L6V5GRLp0KmkarUNspr0teDfpjJ3OKiuXRTcOee+659WnCFvRQk4
d3Jv/bdLEK68VlCNJEuVf2PnlaR7MH0/wD+qANp6VIA8AfM+HX0MX5PbjlN1
jOc0OAeq2t+PYtuKzZBcniJ2EqSuifhvyHD1GYA0sPFx/Z3rOe6w8E/JSclJ
f530r265HKrMfUTdzdGARWwEsJREUhE9QeuKWyA+UbJ5iYK7r6H8h3qr+9L3
IOBU3vdkgZD/LmXnFee86cmRRBDYYP/T3Puj0lD7unPc1/8+nS4vlIBRNZCz
zW0k6S+hiGaIGReFVvAPUktNifJRxfW/BP3nc6toEMyPpob9gh/CvWiEX2Zg
2F6+kmAcJGWLjowUQfykco1NR8+puMLMaBdwBTiNaDzOFDAdSFOqkAXnSmZP
6ODuHMbxAfhF1mZyl5KoC5dyvvDyGX3LzyWyZInR/5bTw0aMKjdKQYUw7kuj
3HFdOWJpXr+sT++s0rt7QIPFWlJU1YfBaPKVjyFxlB8GsZJpNKwl1tBGqMOE
bacz0R6ZuTo/OcS+pKhAVbzd0SzObvbEzDeneJuvyMDkiVdjicnCzfhO5sR8
lKZztRGtWT5LCePSQ0DAc90OeJ5aulWLIRaMiDEP31Xr8i8sD5wnxgl0LhcI
UCxekX1DvomsbBYQbBlGZH2lb7p8574+0A+PSmV+vQzZtVIFG2q8D71RHsmF
Wohh6prjgm9I7iVeLkrjNEqvGmQnxjZBUFSqBUOmOIN7mP5SuvnXusQDlUOY
JHaW/Ple0zvBOot05d6rxvYtmViNUtF6hHeMoihh3HrK1LLVHUNmPUwbzRH7
mJ5TgJnESVc2SpJUaKrjzzzhu4CdFLOMV9ujTmQSNOYHUMa29zBvhZ6ycGkJ
0UC0b+taSlPjsMHEMkrh43d04Q1PSG8WS7z8Zc0g397ARp7ur0BSNuNONbgk
4lHByJBTkzSjfP1cOn/q8iNzkOVqHpsWy/HV+323t5Z2B+TK8rSdC/7Sc0WS
tryKOHJR9VNsX2RzmNVtzEbMgjKh19QRVlrR74/x5VqjduVGuLqFgb96s28X
CLUeqmouLyYy/pltA9Zx0gfWYpyd5XwzMI89Qmh3n3e3I31xfY5bwCSQv83L
ilB1EKJfa0Ekqx69sV0RkRULouXWBfOkpcu0frGEhZCvzmjnGl3tji01/B7e
Pu7snvZv1NvUbjKu9y6FIQ3DRqQXPe98VSrmea2c+A+me+Pnm6ki3humB5zS
fgkvYRKwxy1NX+nVXNacw2EzX68JQmNtKgCQxZ6tNX+0h1OfshG+dgXQOCAo
/eq0FFYJiBqrgw/GZpVFAJ2gfPpzDKZcg0a/Phz0VUmnGSFW0X9Hqpr5sFaq
2sfTfU+q4ixJSiIT/OiKN5sohrs4GRQC38wIP2EAlDdi19wSGZVNkDGd/YL6
uHAEu+nQcF9T3ymyP7Ln1KM59h9+Vz4q7Dm2XTbD8hEyRufqwR4KCuzk/Ori
VI1wpBuOvIjXqzO9zyJ6E8zx5gpGiKFYeoATHEzqbnhX/439DfLVETk5P0Vm
+qTqna0tpCy5MIkqh+D7QbJPs+523MDkF500fjH4qQZlFhl1y7FqR0w5hLl0
kMLCFZtlFdnIpXMEwt1j2Qrht7O/ZhB834LGXKuYeY4n8sdiXUUgUHZBTcW9
dJVJeUXIQhESavplccie256iKSbBPPkLxM0r5NFLv5zfBq36dseCeHKl5kz5
btr7FUvoFroo5oD+p0Wqv4qFkdTihgpJszcr6sMLTLn8qnh7VkfF1mgy0vRa
dwxpXULIOOC12nCjp1Exizt/Ig+OSrZ2Fw41o/IfGrtvRsKwioSrXsCLXAvA
LB9c0cH05EEL8E4igbK0omceddsptoQxHvrOJZytttzwOuyfsRZcoNuLZHQY
HzL4cq52rQXV/Umm6hPkd/X822nz99UKzl8td2MBBmwoEfcSo7svnLpY4tLh
Drk9+TZ+J1WD0a0XvGVjt7HK9UStxnTrve3zbkgKmPLbHupaHTrGZLLibx1Q
bmDM3fCp7Ji7AFO7J+bXhXyRS+vwm44PZtzgdlSanPPd0yHwHaZdnXABo5P6
T+NJiXioC36rL5InlYBWt//ulUGwuezCDkOjfotw0k2dt3axxK0HRyAR8FdT
eb30FI4r1nQrCCJEADASywAWiDIbbwmsdgWaAwr2cNoNDN851Js5RLjt0P6v
oNpMcagX+tQC7LE62H02OQNRALRhonmTPvWHfInnlphnMGDHCv2u0i6VoTkk
q3idfsOFLyrIXGteI+gBsBHk7FuHYIT8GzSvnJry3wTOxowkzKi8/Thh3iEM
ULO2gEQSQtfltC6edHitfMytD2rwy4PnnhGND/SmTe5Iidh6wYgr02mPNL6N
v/Rcna/14HW7AqsOTjQ4iaBMFL9FePKrN3n+wZbhBI6aQ2aUbNpH1tw+YM9x
YLeh4KmyTyfJb39JX+5j+tKHGlPkQI4Al/I8c+F/GItS6KoKMkcu8bna4IKN
v6QpBzVMuqDccQGtzu3Io8sJ1f0ZFCLs3FEgYkMwEWZfs4jB1XYFtOuzqVsZ
H697krkbRelfQt1g9128MLM9DMjGXKsZ6K+WPOO6MZUQZMwBWCurAq4ootWd
dfmAzoqtnVEJ4iiB/OGp5+HgoHH+EHhCDzIRBErVJJinTAl/oZccDbUS+CA3
a7rj6NteDdcES3F5Yg9bODOwCfMpH9xz2SHHC+lZ+9PSvf/bQ2hlZkr900ch
073QGtnbAqJ0F8uWgNh+ArSrfIhtI/2pSTFtPcniK52rIEogqX4Ij0qtMuQu
yLnygIWAztvSmh3bYbd69mCgCx3DVv/QsVy77MM1MGqBksQUKoQoM3y3J00R
bgnOhAsuXLyaJDfC6M3uR1d5wt+WjJkKbyPDvIMdA+nbzmZeX4RjBJBTAhR5
RvdRFNfsRCf2Ak6HXc/lBvaOe8c9yY9XPwSef0AVUYrZb3DaH0Zu3YX4cvj9
aGyJOpyU0CbGeryQf2dgb5/ajHLwNPWBffoAUJOoT3b2GByAB5XM3c/rERe1
/XqnveNkpVU5iHx8rpVHuO+1SgwA/EiY171tY1lRMRjQb+RybRvCdvdikRtn
8TYt8lnC/rJkBCP1Jnd5dLsXgc4dl6rEXRLMON12xgAvlWWIgcrn5eYlf3Tn
QnIPmp6mcyb2mKAPvHl5s8yh3PTA59FyDo+n5MvNUoj3aok+pa3uIVjd4lZq
ISgmPy8bWjeYkT/OVvTi+55ZXN3IS1zNoDaGeOGBu+rRmyK/hd2dG6ge/MeW
oW+MrnAjpPyEtOwhR5h5xvlcLqrQiyg8n6zCtaAbCelUAIqhGAiO+nID5RNQ
VK/NNQPqDLGdJdHPq5kvdOT995ggXUAkWAONbrFS+7oN0o+v8dDsO728YOv9
+2JflUXNEeOdp67/fW7tza1e9RMl/RYjy4O16b7MMqBSssRulXHdtxjZxUgV
f4JnLamQb+IHvdJy2Hpz0iUZ8gOUr9565YnCNJk4PIVIjhbIXb77ebzM0u/O
31yxZXGzoHlStTTqb1x6Q4kjRPZYlM6UlajMo42F8wDLsH+721HMsobvr3k/
yAVq7aXuRXIIa7wm9DTzZLOSSdnN8cIPDGBa8R2oSCsL7bX3C4/bvJCFMSxE
gXdfwpDdj+7uzKMW0T3LbiG0l+DawtJAsgJRaozlRkCAO6+bQY+S62pF31oB
VwIf3anlWitUNs3wTEQEBBNwkX1Ms9y4jk0IL8CtWEjSgzgYyIIN5EgYIkNl
g64YSMT7r3+BwwYxbJVDiQKN5/iBKTz5ZQp0r9tMgjUzqvZBjRtL3nA0COfw
YlOa53eGTp8b6RQoACy6tVZPgFD1C6+iP8igIiwJX/VBS6hD0gfqy5x4nk7R
n0Nxn16kIm8UdKQaKxGjsW+TUySsVbUrOenSkvuDShZ7oCyKLrxVyf8sLXMC
/zB9RDC0BrdFnhYkIBgRYAm17ImzIejm4TlVVV9gTP0SXOTyJc0+jtQcIY+p
+QwPXL5sCTG3MCaWm7T70mv195vN7QOVpitZdX/UOvBwhaAVRD0nJAg7p0Si
raRnUF5pJGQhC3SvdHatowfSKcS+qISDHieawrnd2xw9uLLiepXdd7cfAQf4
AmAy85FGnOkWscMdvZZeoSW6TNEfjx5bnnOU5uPUBb3nhw7GWumAifiGAQ9F
PawUxAY4LDtMNQ+Jeu3lakGI1GXv9gynRpBRKVhK7h+NQgEjnqmmjmuEpFz+
2/xfUz9e0PAqfwfvRVcjcB48kBCV6ABFOK+yu9RoPkJ69dHMVngHflNqUwsj
FG8BiA6+6VxzTR7F/1nMbschE/FeUOL0YwBXasqjEcRohFPUMtL40780dhT3
vcho9eBKwDKaeyU+WUSE0HnRIpQaHxiKubiRgvynHvocx2OoWzsyw2Yd4hXS
iTH67KFK7Ss/lRp7RXZu10HmkuhFdvO/kOKiE0Id3fLZJy7eyHR3CliSPEJv
rGXVZaBALd4TDX8ScuXtvyradcxCuNmUZlsIdbGSOnwsrmDuy5B2yzyhHUIi
1cIomzraQij0oXjEald1Ub9GUZBzhWRB08R+1nm+Vq6QDQMPs0HrzqDvOryL
ITZ2irN5GKPqu5emMZ/e3nGa+iEcGCqUQGxbOE3rnlhT2+6EFGmxr2ae0AMf
z2qJh4dS+LmoqMyhJsgu/27fL5gHh+MU19iZNp7Rwfd53P0zpHPXsYH5//C3
3lRVJ0t+MMOAc47zaBJxmWyhGTOBnc1YXEXKVaak2bUHnQ0pFFR1wawDsq3k
6IPmQbS2d/ZBRHq6eleAZ08Bw24m4LZiZ9VLaPq3YD3KLf2P9pvpP6mzyJPx
z9YGky+7288jMTB7kK1zwZsmHijHlF/bvk42nnsi+nJwDUojPhYtQpzdmKwM
fWEvx16CcjBvGPEhc6wsK/jrOA9F5qbits2UQr7MNp2YIJooaGAiyllykX81
EvTyNnn7X7MSpSxGV76lWzf31kw+KOlIfMovmRYEs1k/0OV6DholQWuSTiFb
3Z+lNET5kSh/KZXgtzg0IAeBgMHVPZ1eRKdWNbhDYRgTAbu/MeRWIqjhkV/v
2645MvshtDuP6eLFjA3jYMPy9bo9IDXsjaeFnuP5zVHGaE+X6RWAVLGzOKgr
ZaXnW5i8+cWKquVxW61O25Mmw+db9XLg/qAqqoTHqOY9nPDHqrxx61qu/ZIY
B4IPugMoyy4uVCf33Ri8fnQYdZSKd7HgwtsZijyoih0ptShAL8OXxZKv48S4
+qM2IE4Pgc22SZ9WeDA02l61DCbfEiPJrJU2MyDCF+rACiNHsskUrOYiGRS4
/BCfI2aQ2BtODOLrgOfsBnEOCEVYYsrVvhHCVSq1mZsJNkln/y8HRIoUcxrJ
a2Ik8EqYXR72+9znZXNIFQXkJ+YeCIM4d2rINmqNMoGrBKW3CME2l3JAx+PB
NBwfc4wybDrotr29zcfY2mn3Rh0zyzoHwxoUWS98y4HrOqm4TQ9htC4hxxM3
bTsq97XKpgwFyimZAqLoC47hVb1NFx23hipogs5FTnrz/BKugA8fXrLBANuy
kPDyPUvY3YUHJnVAPOoVl5UzdfNca3sM+NsY4Y/43itWVWs9wSi6tFxB+KCd
SxcBWznkitBfZIZaatl2JATuEVJGFEhrkWC9js+/caRoZqtHT4JfohetgCOP
L1umdRyzJ8PtB1zs8bNPOUsa3Y7Q2uWEajixxBwm0/WavT7C3XcYLtV4Gbra
8WC3yfsTOAa8C4RbAExvDuJ+oT9qQGtY6ZcgfxDC+8ezFEJfaGdfbQKXCThG
csSEB82hZcGfm/DnBGsOGyMLsWe3MGDYBIecBQPg1h+/L+Q93YNu0KsztNDW
fjFnLhnH4C6MOac3+y6wj/3oKM1X3hchL0qV7mXXgqZ4zy/B6yJyy89nY49b
kKSXjdLTmCE6IlPgSvHuLAKVUyXvPIbQZiuWk3WaZTgjut43c2yGPNfzIYTh
luFCSNzZYYj1rrRwypNqQ82PT+eb5Bi+xN+D0OCdpr3bXq6HdS/iM2t8emBF
j2GC9n3Or7yD5++7iT8hUGzlpZ843p9CHQg4o4AJEaFtigYMrlfVwjJMHqf8
logHrdQDW3BNi+uc0k5heLQoJdGobJ0DSTg6FJxn82v0fccY9IXyo6rzwVgn
akkHXhv6QQghjOLcJSbhqB1ev8tuIY/pjTiFaW9GYm5Z8QzhFy1HPLxh1Z1v
cMLTaxIAKedHmjHqg5C0e0a7sC926qzDM35YH8MjNhIkZKrkalAKEa/1UUYO
IU2KrDShAbvggF5qfTTiileBH55llgay84fNahmNo/d6dxmw/u0ZtSNiZXD5
zmzCHFZ2JXW/Nz7nz2KGE+VyPoywVaF0xF3XPRDCMANSSSJ9sdvJKIg2/5kP
0uR+J94p41K/PHm1UimLNEw43XbNV4TDNwn8HYUM8QgOtFxpdBhIAZiHZPBj
VX9VZrB+XJRS3k1WXI8OTENLuu3KAGq0RzV+0lAurpWBqgZ/E17eCpqPjOoU
hjBu1NnQvZ+MDIANEwXFEdNQj2d75VPLg9Q5r6O1kJg73iqdmXFDAH8sEp1V
YH4P2YSYzM4V8fKjqYvZxM+NrJEZfSkd3INeVMvEGfa1Vi3Umdftx0fRaa8s
eImknVY0/hsy0lD0fpw0q21Vp/6CjuYl+9QlZEzinUAD1Sy9sxYg+BICg0pY
mDrldwsSB25e4HIaEYa2GcAKzOECeGCHw9oVN2gG4+JVhgWcnblutop3o3G3
eGNlepyDBLl7az8yVxczy8ocWpCtJtrEyKERHBdoNhOSfR8c26Dzfhw4AzCA
3YKcCUvIsjDrvM7ls/KSHgwMx/Kg332wyxaaIR0hUc9j0ETjAYymzbJLz462
AvSb1RdSJlOZCw3cYjcUfKsjtTlXV66HiZlQg7CW+Y0zK3kC/tw2spbDKuuG
++IrJbqBbjYvgX/kTEcREyCNbGXLxyXQWgnDCdZslQJO2dTrq5PhsTsVGjs2
0b+Hs1MSBKRdhTByZsPazhtWjiSCbMisnuHR7MJcTca927n8Nb+KLHMEWH3u
LQ93h4daKT3JHhxtgRab6g1povJmLaCiBqE4aj4yu+RocVT9RTjLjX8e22Wn
v8Vxcf3U1N/AzbPNNdXAH55LRPJCai0dcWkQPVSnOZg0ZZVo+3/VZE5y1F0g
TpiAgPDZjfQVjdJCe/vJdWGXV8nz1f0isOU24uCunQN0juTn8QYHriUCkR//
12BkcrhwLZtWvZnJJXT6e9zB5unfIMNEK1SmTpfDSn4pu3lYuxa+hll5Y7CC
DSwsQ/MYpZPaNRBz3NDmGLt9/kMus55ToZdkSUcok2Ua8cjEbjMuZn7J+wC5
x7Gh1MXNEyugTQ2vo3E5gvJH6/UHy3D8Uh2JSeL8tm7VZj5agzD3RWPLDqIJ
+QsT0+oUXogV5JBIRSrNprMxEDLbESb2YTGh8HTEdBSmgqvrk6AG+FrHzEnu
9VCmNnBj44GbtB3/XAm5/KPOL5g3l3oYp5q4YiUVCrEJPCsqJB2hSNNnEajV
73cvZebRisEWn9akaEXTOptZxmnRF0tJoUWntx6egi0qqx4ZDnhZypsTI5d7
srSdbTUggEeMoYvoo3owAgK/IP6iY8GAKzCREyTBgOwhAclOkzJtm0TOZnnq
QewOIcpwHYp2Lu5aGSbDkXlZi7/E/OXym03Jf3HOTA5IApJyRqzwhPKMEd3V
P4GjBZrAvtcO6UBCwyD12OxNu672f4IHlngLK39DDEvgTQwFvLYMOSZZj1jf
z2e3lFxvyQlES3C+CBhE0MKacB44MZPF5pkPlR2m1N8opeNitJtg7h4EJytW
JlOCmAGWw6IozN0S0fdZt8ftVQ/jie89EreEahA90XQW5JF9007bQVF3yIwC
AJEQPxI/7G+MkS0dLP3e7L02HOwZ4LVQHrW2ARV1erm6rosmWWpshQWaMC9y
+JrGZFcXvogIaQoVbP+PcxY9N8fz5WLWpBziJQuYnqBXC3skpwvpwamZSVlu
YdSixn75Cl1Zr9Yn37kz+3oQGhicHr4GTFjP2Ihg66fygMUkOAYX4VYDRZgf
KUAkHsEOYtptnnMkkw1dhZ/EvU17ItAMBfAeyWpgPsof7nfwL2DrO13oL5Ur
8e6UDFV+JtYKpYUiyAzHBjoo7ldfXOQqZRWkiSKJfbPMSKPLWNWiAhYJ1edi
oIQIYDfXG1Mri6+nZxjw0MUIuazHDRRd/bVhoppEYgu1OjieGnZUMWWlXNo7
dW0mamd3ftktSNi6P52pYCKGXcYUyKC5+wdGT14mE1OqfJ/8rkAmEm0rybGP
i92A0K7WCZXaP45QgiqQ6Oo6jVWEuBir1sMipVj8YhbU8+NS0EvETDChQFMC
4joMx84AsL05dwxutVo5ezV6SpDQ7N6IcAC2LTP7Gb56bQ1JJ89grP1DEd7n
ZUkwhKgyPmJNyJ33xD73txgZuZ/zx/STNR8vJzN+FjMUAK8ce2I/rVBYec30
qsYZgeE23XItOGuwFsXOYGi6q2y5QycMPDHVd/HtDPxoCw81Czmv8umZdPKZ
dxZG9D9QXcPTG/nmd4m2Tpz56iRhSZaRj928jQdK9D6MsDpGMe7SZXrcttks
s+x7l/csB4sMNa1EU8tr/evuycK9FDSuzCGpik8fmNHfk/nPLlmofYBu72JF
AI/EftaXgCvPDdxu7gEbH1plDdTTT1OmMsNZM0nA00xQS2TkZ5TYoIpQC7+u
tDcivvy+od3y0bUcjAQgw0XtveumMRm1wDHj62BzTQMldtbHzJENK10QDz1/
O1IrIe5REZzItXbFVRjveoyExjgFHpgkcmVFNMXmlgnf1keEyRav0r4yU8jq
wfMwfjdED+FepX/D4t2CcT+Tm2IovLcyQa3EFQeccDm8ttV7wqXlBU57DNYE
7VD7dK8aUHPI5T9z1AV5ZDWuZlgg+abaogV2qNXuufIQ2Fal3CLFxDl/Kzws
voHQFw7d7CS8HU5mQceEOXlS9HBU0M64pfToKOgySMGg/wndflDwLQMCXgL8
WPMsGXLGcJJ9kCM5V8zma+AmJm0rlDWoUkK+Sfqrg6o+YWvRvE6IB0JhpNdT
gp4HlVSWBEzhG+9PvLO5qKrlhyvBUyHQX0NF3026DyWJSCheUuslpHPE/131
MqfLyaslQWe+qHC29NCIDoJYfvdEvdV3ZZEdH5nmU+fGqoaqgmc1BJsPCP5Q
EZwITkqcS5iNBom4YjCoU8AJrYfzT/2iJvQ57AFYfAtKEEBDj7Z3GYRkor9M
vHlPvitvCwfwd+RjPU2PDwla3BP7G6SZqjFLRusogFaJpmJQA57l4IdojRLb
4yxjsqDwotldvVngPnf/rhzVx0dAb46oG/CAmEGf9nm8oNJl1HkX6ugUaOSo
vMPOdt4ViXrljiRsiV9ye/NcfNbBuvyhNIPinVhc0O4cbtSzBnBQhEiDX5Pi
z9G0yoV+rFql5uVV5EYUbbRyiZhfXWWAu+/Y+9ljcuqu+diLtTpmrl+fm+T3
OTKeM1btU5s6sCMl+B7k/FgR5SpR5RPsBBliD3eZ5iYBJNY/pMCFbE3tD4sn
T3Fj2yiA/pT8VaHf6xTn7nkc0bbqjfv8G798zHHY2HjGzH9uu2b7dEuQydf5
NZ7tUwtUPidbt65C+1yV0Y+YXgrRBfR5dg5ABoR7+Lu4O5dKZdK4si1RLo4p
hUuJsAB5Ub0u1V9naWzs9kT9gneVhP6J7+KcBLw1SduHcZ9NpjIvS31B9OvC
qTTcWBwbJAxROjynFNpObeTAaIf99Fb87QibF4IobVhUqEcP9E6UYAV8MOch
LxXnlEWHv+CG12RiI64kKaHDQ1O1iHDmi8xBH0myyYvbY0wbVwNJJepnxabP
dnG/dFpbk4Q6DEbN8auHxQ9wj1T47hRsBQSDpqi6kO5OdLGYtgAA5zWqSu+R
23JJEhyj4mj633P0i0hOTPk8Z7PyBfZsKEbOmptp2OktaTbhrdKy0QbaFba4
K9IavqIg3NyS1+h3slxEgUt87eOcq3D82qmCzrN0MBeSohhdB8LVPIgWSTNd
hphCCyQ7FAcYJdm0BZo5T9USgSeMPm3mbcl8ifM7djWvR0S74yIG1tDEhiOW
n3KIPvVM8JDeFSwKWdHYWjVHn5iGoX3q2GoIjC/aVrAEU8eTNAtCaf3OyPrG
oG5BhM7rFPOMwpoGZZumBJFP0AfIBmWE3pKyHnidJ/hlnjvGxzOMCndZ4vJs
gfv3WSD7BJu+CUTcWvNXuXxZigox2OFHuJ5Y4ym5+W5Mi6mi8cmK5suNaDNv
ryXKtXXIDQgS/s9tp3KjVALLWmfBxlEmggcB4GGEZK86/g+pHRvYyBXgsCUU
0z7J/1fZV+L/Yl335KqodvXwYbY8rg7XfBsTfnJKN4TDfdA4sJxMhdNjwVcF
RMMrtLFNkobScvhM7E6hV8EbHvAEG2zQhTJBT4OAxIbRaybZaztoFsV2roiD
ktaWAoOhtju96DFUvWnllZEVVkidjyD4s2KuBJZtPvAi0u4EcX+KDyUNFbj0
wpTi4+LgFUvGDZnRZJYFL0iF6szkKvz9iMfO1lbJAiYrO3e1Ke1F+PEOXWlN
EHNCDU7Uis47tgWTK34/CEvPx52oaJw7MmspmbKDurxHM9EGcPo+KUNkJXOr
3V5IGHIs7UUdFfJlOuma7E1goXTYhkOYIwO8chG5X1hmlnR2H1+HnbjYF7w2
mMrhArZHX7615eUusYbmTjFw9M7vPr7Me0yAQ/XCbxH9Q/lxE8rXssQU/6N+
Q50DeqGS3hhKxTtJLMaScDh/FB25h9zmDKVX6GXESiThmhpbQ/suQNauhfKk
J4Y/+GamVHmamdubp+jMoimsaDKc9P8Jlwn7Or2B9XweN977oZUQYJUHpCot
1UuFDUi3Zquy8Fbf/o5sILUI+pJsxxgZ1DP5ta35KZBPnGQ0wVh9HBHe1wYg
z2nPI0pIos0m1BQlqaXjXnWexkVLv6o28vff+NXDs8882tiudZIXcbR0Osu6
lZCACOdvtIGU1DGFrmDUWNxq/PGqyfeaTck92PuKp51ssDqFBwjgtoxIujap
XWlHpR0fnvRugKL/zMtZ62UT5VBeCKitZguz60nFB+bDiN3u0Tsz1IvGZpeQ
H/QqjS9MeCc6rX4ae6eEJWxmfUgKlKj//zyRm1dEl/ua4KDg46pfmxk4/klS
itdGJaIM1gzfVh4uPMvPjHmY5eiUDTSBSIm3kOeWaAjxpKAuAOzX0LBLB5mq
BGbnCHRw8HZzcP4hRY5fbUMiQtNm4v+NrltHXw6+zByUy8HnvxjYVF++ZSxT
i06NfPFhQuBtLJX3ftVGZTy54OXNxmNWzMcYozGrY2KwAGe1a8hrap6kSpSR
rQseQ25kUzLw8dzPIQJiwVXihgU5RDCEUPzzWpnOPd4B4NAuQjMBUoHCIoCj
g1r0eTa7Yreom1VGXOWgBAvk7nt446l3G/WuNtc1wU9DBIW+N3j0RJ92VqOZ
S46zMT0NcOqcPIbCn1LFTWcQX4mh5RKnzYfQzW9r6YJ1Wq8IV8CZT1C5wrGT
szeRjMBigdffbqWRZALTqHeLryN8gDisvnR4rQtrt94WQrZKTWtWVDjcjWAF
e8XhIR11nW57CKN+uTLOKRIThHz+wA4v1EOguDDQwCFHKWldXxYgg8x4UJXF
rVr6tOUJ1Mv/PSIJOEyKM5gReRx1yvm31oTq8J+A/St77gJvr33z0UnaNnX0
qrjqjtMkvsPD4d77LAVyU/89VHmOSrKi1To8gOUNOkmrzk1t+kKuq/oszZj+
pwnoqlHJSMWTJ0LhiHwy9j8x02XYQy2kW/uN+b0DwJK7WfjdFXZmRTB+MILN
gLs+ZE+lvUvQWXVIi7Vrcm9Uzv/SlfHnzu3uLpnY1z5k1hgzfzaqdGEZvXuz
JJxQHjCa3EP6SVhuKKQJT8U8l4BNRsj6fHi49ZZ2BhU3eLY156gVo0jRLl1w
BsbA6SCpzUqQBv2YK5Pjgtp4NsdO2jnJ5tcVrS74ujOm9DUqx9aSuRVym2h0
969mDJFPMmQcp4KkY0UvsuA14Zc+MIoqyIfhPz57n0wvIRAqvd0PpSt+OGNF
y32XxhxMGoonDALOlOBSnEW99Hs+ZnFR+YIvsZcSxPlnPjsZ746SBlVg1t3Y
JVgTkoOBHuAcw/j8mEFrxCYTizUK8O+Zcvu3Q7AWORLEE22wtxIKD9eXepyR
v0g/kMEZHEuBItUnZ9Uq9B5ACdvZgGBjAXW94PV9gO9jj3gBX/JhmZYVOEwH
uLn0+ZSeggltf7cbHho/6g5WcXPMdcxBSPFlpXULlIZdu4+X74bToEUJy5jZ
cxldYigp2O0fBtMtPT7eyIva9fz3GdvDWj2JJdsb5sPxGGly6XERZ/AkwdC4
71G+vNoPK3ACiNlfH9NNUnbqG5mmOCyaEyFoqfc3UN/oIv4ZdlxLxMvL9QPV
u1TlZNk4SAd1xy8VOOvlylximw8qr/uPYkhlDNsJ569u5/aSm2Ra/FgJ/9jd
LjicNC895WoRzH6RDspG3LA0l4KytF8zMS5TuPwr12R52cHAPmhs7Xw9dVY1
uRYdMd0Mk77aWHLGX9kFpicrlS6eU2I/gvF0A5EBn7/CaHikVg01kwSir+uN
rVC7rGHUGsfwFwx0NvHzvddrc1apUi+Kjh8g03ZidQmXd58+uRMVN+sqQpFQ
ksfwQHhpCBURlLNoHKolNmfi

`pragma protect end_protected
