// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KmpKhQL4UjU4FVlp0rQblTXQ096q6d+kNxX4WfJiz6dbg29q9IpLAWnu/xT1
PcUowTN6cNUgbjZE+HyQhFdatQpORie3ZTARO0vnTc8G2JLmKwmc1cNdfaEF
K26bwC+1VtmV73ZG5WtbkdmW2J099GyD5BBZ2jOQt9iDaauBwPjAZGofEOAU
fRJElmpwT9vOIJ/C9J5R2KhhMBc6hPFzDVgbCrR0FYojSL/eUlMqOiLI0mZf
dE+U7IZ7OA5NVongAjJlg1EMLQVlAfuswf8mMtmMrAqUSiuuIPY1S4RSXgX8
MCFHgoA/QlIyo02fw/P2ALlBAmOH984E1a4saX/bFQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cEL82CvFKJ73R7LqXIk9Vn7N5UtiWs8Et9UXVXGPkDtgm+zUfm/Kawht5KCr
0y72ElnEUduFhZYosA3mWPkV+33cGc30uvWqu7vpK2OYaQ79FAh2wn+ft2JK
+QZRU72T3Z5XiR4hkAglsjOyt+Wn9QA0jA73RKr6pM7SNLl97aQb3URhX9Q7
+BtitWDR4P5j3F+yClyg/9zS89W+0mJPEW+yvpTEIjLf9mPwFj9oEClHrozJ
JRM1J1xpuK7g4L/wZ/Kj8LqeqCo31ygdskDSmS1yRGp5YXzRmgYcTnFHU2YF
Uk5qaqTwWM5nEEyPY079b986gBKO9wnXMeOvb2n6IA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
V+yvoqN2ae+1bSpQw8TVYeRZc9uw0uJd9kugsHh5U5bGmqO7H4N2ib465KfI
QF7k5oAtvkHZYwiaW7osZw1aLbHz9i0L5Iu6ubjnF3Bpk6JkLI/WzTUdSnjC
TuRTRZBs/UgdiGYb+r8sxKK7KvS+rIWpZTceT/l7dNM5QbFZlehj4790xjKB
iFAV6lfKq5xRsyw774zxDWWcJMwmCP15a01naP2B523S2nKdweqSqV/sQ828
vw5QKKF2aNOIr+eZnuMKgm2wp1PfbUiAq22Pzm75cMTy2kVzFkKpkLFxPH9L
8cgqkEE+sm/RwAq15qdhx+btU38jwiVNCGViCzSk9w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
S01ErTCtXZ9/xNmKJTD2plAHubdAdl13IhxQgN0jjeNZT1RQtN0Vdoij9UUh
TlwfZqGG2maX7Ye/ddGMi7zS5hzVvrglPO1nNSDzedBwduM/fICkX7AzGY4M
RoTHaq3zBN0xuGQHQl629wrpXckrlKDrqb+jnotmlVUMkqenNog=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uNMpVPIqE1e185kGADDknJMBTumPl6tg9dZaTaQVVYaeB03QRYupD9AB4nFI
k6YlRoO9GXNyXPgt8K6hq1RJj3emVYuy/ZaFWP2g0g3jjZkdaDGJLa0l4q+6
V6ZHDIt1LC1bRitfQn33Oyeuif6iwHBX+QuySvhm1ngGyFMwcruecNMvyxJ2
6N6DUj7GEkyR2Kye13n4+ENv0go86Q1VcXw599PEMj6IPsVeIQUWoEXW9wIn
L+9vfRky3asKmm1UJgXZGr3ayYNCfVc7+Sl8NxfxnAmR8Ewq4BMKVgkYo5pb
3RIJQKP3zyOKm2XSSvSexqI1SFc8ylEiEJs430W66KJm7ZFSMopvtZtdAgkn
c5bF7j9w5PhTsoF5+arJ95VIU/T0dptPdWsQgnzp10OIiB83PJgQJBIEHm7m
ifmgrVbdg00y2SrYiBHR1DRJNq38oM17qZ1ZJWfv8WoBnsDzFbJjjgvik44I
oyJSSFUIausnrzh1wfuOnaWmmXYxRizx


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DqaFMMfEzAhBo/GoGpeNCZj9Xxs49fM4Rg4WiIljaGcno+pxXTvuuSq/DYDu
LLHRX+SH5mW2+NyTGLIizd1z6bX9T3koXl9TLVB2kkGMmmNRCTSEECRCW8Lg
hMHMS6UL+NxrcmtMZvEzyhXAsGCoaBQcbOQVTNSdNDG7HuPaTUE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
myyjL8QpJo8FW55CblII7uAsN8gjJhF4K7ePkBiyd+4s3OgCwEZZky5To2EI
i+RuiEXWXAY+cov+UgdHyV4enhkIc1eGD30zBqiqZfDbibbLRVU2aamitWHE
+LclPn0vesqOPv4LusTWamtucO4ZOPRucYFNaJOUmdtIgxDkrEc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11136)
`pragma protect data_block
KoAGMM0T8yZGk1yPut6XFuFu4vH2uAzBGS8pbm/qt8O//rfQmzrC2jyZkitq
RLB8azeP1Hr0mPx1cWA14bM+8NfVfBQQ/w4CyKcIJOfbD1lYUQJi9s8zuCNv
HFCrlt6G6rUFsFIMJgYazAsF2QUHIS6fv566BYGiseL688C+BJw9Z607gjPH
bZvCd80CeXejXEOxDDGEJTk+vm3jhHS0/UiBg5nVfuA2/tE20C1EUmLH1cPf
DeoGFIG0J3mqJcBoIz8MhUeSaMZYSGpbd4/wjaYXnVKq+UmK4GH52g0sni5R
00dzHUtuQNQyiKzvQZAq8isNYJpWqU3AL8L+dJRoB8vGHN9a4Kj7fO9kKIqC
BIMrQBo9xvxgqh7Z5C7h18WokAI7PLj9m04mqQrKHSvKxrnFs0aP7p1Jr6A4
WhVji3FAimuCpdb76oH/wPM7ic/iuQsLmOmwJksdP/Dc0M77G0h618zIUsdo
fjrm3ISF9lDU3NhdRUyfbzCt0kIp76DqODwKTFIx4Y7ba5xv551dGBXlEccR
5iDzktmb3TNTewP6vRrdw0rzsd31m+dMnF9Kqm5Ht10GqJzm7WMgLKJ8w+od
CrExr2YFf2d2ovo9XqhG0X+KgLdYDfhhz/QIdv2W+dNKOjLMJqM+poXEw0ii
LnzSPe9ec7Je+FlmMLbiG95YiG9jk1f6HWB3z1WI9P+wxqowFmzgTCsNbAKO
J9IpluQ3H0cVLUNUj4/ZjaatXiTNdxCVzI2yY7ec7xotLSmP6LbJ/vJ5LcfU
G2tGzuqMuB1daFRszA2DtWe9wFOCH1KPMw4rmSVuceLiq+zJgldtpwcP2Q+N
WSt60YQpgF3KHVvxem5N5ill/fZrlZuh3EyKn9k/h3CLWnJuSSndknZSCHqg
CKKlZ5Ed6THgMuLhd0eFVO+jqkGPIDuhVy9d1veyT05WPnXRdoMgtJFrFhdK
3eVOls6yfplxoq317Tn9MX5kdesJcW1GsRAlGN3qZU+sjnK4j8SbS4pCoPYO
72d41NgGkaIOkDpLELkgK5J1F38I6oI/6fzbqgnOcv2KJ33AygnKxpyABcj7
f405VxUhgkPUP4p/20AUgah7PRvqBy8a++CKRyLbquYgW0UEVeIYMxG9vQa2
cD7uevltKGPEmj7ERxGD9L44KVXIrmJNX84apf+rWabdODUxLxKbBJW9d5Wd
XIFRQT5FBZDRsfi7jRpFAhxs5fKaoqgdiOH2AQjJlxa81fRya2paQ+Ip8bks
nsbu6BozcwXrcJAX+hir5gNcZeUN7DAM6ACmthjuTW0Qa85TPRQnsXGcwhDu
1VdFeVp81xDt02s2zRjYJV/Qzfn+HUTviIqG6hujToozliUpYJY6JV43fudZ
BdcghnNT+BMNIMtjYJMPVg6uLG7nibXFfjWxGaPBQGHolxjEVJikoYH2+IVz
eSRKYEbSmMwQKCE5/8DcEuazeZsJ6L0JEIl8C49+8bcicqg29R/ABcyzBvlD
aws/38tFXzhNtXr2xxAKnf7nXevpnYsUCvT7X4c2IYur5+bjtI+WClc7wHnB
bJrM55IuJmAqzVcDpnl6Jvyyun4+7Igs5SuBCayIXYjwt0YQGZEoFaWJh9dZ
qoXBCzUSYCgS39xn6L+eopW7AFMnNdpyMcRm9vz1OpqjkA4amhWPzdac3tBX
ipuXSqmFkUI6VNrGpWH9xl7SyuSngeupR+pFVqkHKOI4LcODTHZv56i5P7Jj
CyN6T5g0SotjyN4clIZmfR1gbPGSpOAQjvAxBf+QWjxO5kBM9GedLYi+S6Oy
3i9J2hY9KwD1CeRipRWbEKY948KMN11tlhIR7f08whKZ4T2tzhwA8qsFOfuy
KTDcW93c8SLQuCE08qmqG+iRnJAzVgNNH8PSnvIu3GFdqcLmaQO51w9+PsFP
CdQRnKyZagioOiqYlhKS6cTKGxKyBrE4I3zE3KUWy/9Ip7L22l096I1+KLmA
Mi6WZ0RayWDLPHlR1s1mp//DmjFagXANSvBpy8sWaF9uR+MePsOlnvYdt1cN
tjpfBd1VTHiRxqPvWs2SVrrmLnd6/HK6/MBIxl/15y5N0o0Q0IM0cdpct5xh
F2t9RsVrrEDTIcpapycyP0Mw1afz46wsVo/WpY9/WR2UekwiHPiVN8sATXbN
AyReR1+lyOti8iY53QEnfb5oIPz1nBXLDeLebm7qs30PWgkw6A8bns5RA3pY
JNIxf7hJQCzOUQviCPTVtPvGa5r5DTOjFdCe/xWGl9AuwznLnAN1DFliKdZJ
iQEYQuw/1j8maqkMq+EYy5x+s4hOF/fTAVveS2WJ8H5KP+AVHLqWowe2N64A
9fD2Zz/L70YBPf5wAC0ErczQKN77mYoXUnXkgzGetMw1dW2Un00NF8bZD1Ok
Gkxhizc+Ty6SqkHNtOl0Gc8ewhb096xVY6hiVgUZOEavQhiTft1kHMMFzJka
D//ubj8Pwo6LIWwLZgHzk+pbKgjlJVdjBa93LC5SS/r45yvu2vAEIyb6reYH
GtLBWAhLtR4JHexWVtDeCaDtuSheO9Ice+Zf1qtZcoHxVEG1I1NMzWhIrFb3
jaIJbdannX0nLSmdBaT3BS+5LFMB+fSfK4Dn3OIdpIVKtjxHHSnzLi+YGGrl
izKl2xEpZVaQoWOgHLxLgVk3sOER8XxGfhtu0Dw/CNN5kXNHzJZQg7lsD8kC
c7hhS711GYOhyvLQFU90CiByoQZxtsDzqpDQaefsXpb8DM8MJXkwTMSEfEyq
xAnCtcFjoYib3ws3ACc0YI9R23wf4IviQOJLdB8FkVYehKTdlJ9nXAnDrzl9
2IAT7TSfAgMYgHYlCZDgAILJQYzBIxZwe9wn2ZvY3DDjr0U7FC/VMGZZyKT5
OWZzCV/q3SUVyiI21I6+UC0f73w0Hrhd44MkOqd5Yt06NmINoJe2lrNOkspI
hDOPH068gjSC07u1CnNFLTzLIr6ZbWbsLp+jEE3IiMBIPWl9me3YLmV5EEdD
cyQ7gF6STWhwX8LZUmL3Me/NttH/s24awGC8KB9QkAhSq/j4WNIKdc7Ij/nK
fDlA2Rj/FJQQ7DRN0xpHQPD4d24kEyfi+iVwv/kMxgrZZXwZXW1omAglsBHB
ksn0jcIHy40qcOCIAcD2ivwr4lvbz0M0aavcvORhvHz/dzZo1ujtIoMtMwSS
7a5mAwRHCD0KKuHeUYIPAQbZDBlR3rl2QgO6IUb53kCQuR/8nyJrckCJTWFJ
8I1vdQqe3VEO3Rn0YNKCaBU0cBkTU4hqotWiutZKAXme+855geeSymhMT8DD
IRHCaW+lO4mENo1wqdgxXL7TLT0b0gzwXEcarPI91FMPxGO15qyioP18f7YI
uIY3CYjdD5eSPprW5U3vJ4LXgc3IFe1LOTbxS3bzNceNkPIdi1azF1WZlT9E
TSWlW1x8zWbOrTJzSjtIxUPRzrdzRotYrGd/4XJDb3evJdjDD7Wi352lZ8/E
uG5UfXWXsBQcW77I50RFjJJ1NQ9er3itFw4DFTaVaDQGBoeygY30T5s2Ywa1
Jmqxd+PxP/PKvn2Vzn3wvbJBL4DqyYbT82jORCnl8zguOZpcyUnicCgclEiq
nxhui1c1bWGWQAnGM7PxI7xCfIo5d0WGHxSZL7v5JscuHURGzebdIY5xdNQX
KECCDtVVIFjSbaMsM0bZC5XzRlf9uK7c7bsqomCmryoGh0lLrhHveIVEJKJI
EJu2txbv8TZh1XAerJ/COgNDoU1D5S8453qBbG8sBR96dKdbIOlhO9WudIBs
gtJ/ORBvrwCPmUZnxdZU6y3YYL3Fk0NhstGy5U+sr/H1w9wNPYgk2VetQmSc
VyuqX0mqVmrM5FqaNH6LYzn2vmNBrdRKcy7UgOmfuH3pmjREPiL8+P2WaGkv
fFxwL9ZEm7FYFcCphLrgBWFisRQZA9okBZzkyQQoBtv+C9IJI73bAAg4TEWL
UhCV8eEetg5SOgciaoEd7GdXGsS59RMnSBt6ZsV8q9bhxUIBJCWuuJyjQz0l
gzwRVFsTrpqgkE97nHiAB9lrq0w7G+RPMbsBSvPmnsjCd7Hb0C07kbl61Cgv
akhtdizxkfGdVOFskjX3ejApFF1uRFhrm0qIRAIsylekaRYnqwTR66qR22AW
g9J/TqZCsQbMyo0yUGgZRxyUUlk6uHIuyCqKBkwz3/jd4TdbgrNUggS9GRmE
jrpcFgAkvRriNWiTVTGjAQtecLaYOgTCXwoDuyyUMpB5T1965DsyzdA6/piL
tmjhAf4C9Q4W7kMi0B+IwKVlgf7Hj3kkPMvIq8iIEwOdxjpXgDJMPRJyvMDP
vl79dG7nZ5ILmb1p5VMFw1OiywOOo5iQ4z4QrLjX39dX2BdWrDQiLyzaWI92
9itvPs+tKwpljeI8hBZXDAI8Z6KbVyYMS+je53CTsSOUuzXBLMXtmWEYjBKZ
VuP5JAqXb9s0gZDI/hsKRy+3yUZatF8P4IDEHlWCU1aQs6rTIVNVTEXeaNUx
8WMG/xcoQzEHkg1THfibylJ3ptHvZbPDQ/KRjj+BFvernayDnXqcOcjAHuH1
uu4BpCHdMtAcFBo7maW6EWhJlnrCZtKUeUG2JNvNYiMYc/pdy5g1trvqpvzc
V2mLMnAtJYFaAJ7UC69iKV8UNKc6VW0/m6YRXbh0M8ffs0c0yTa/lShbWJj2
HEzmYlv0TYuuzulm94CPYvDksQYgU2nncixAQ5X9fvvI8H17vPaz7Zz/cKBZ
iGJqKSn6iqkXWBcNWM/XyWm1n7/q4jVQ4Hn0X80oF8KcxmjIbpiLKKR6weNu
5oItrtL7Xlp0YSxeAmQj9/8LE1sgLhORGIFCXy1V1q2aPlYvSGs4p9XqgTD2
jd+DrXZsbqv51crpaISVFRcEz0tQs5fGiTza2zbrIshkKngPBJcJgeUFAEs7
U2xdMam7oQfeujwSYQ6nxQ8Vvlt5yFk0BQibEoL6MR9go5jZS6WvOcsK5w/x
HyNFSqyLGiDTIHc4sD9v6AfV1RWb4K9gH9snJ4koLSecDq6FnIdNpBj+Oeim
i1ZEAOl4HoWypeRsY2R5PvFXt+EuXwXov0WDratD0orlP+OnVHIeKYech7J5
DpWFIFOOxLhl4T5m7ebXHJDMMwTtJJQe+Dx6TxtkLyHyWXg2jErwkqjzuA01
wJGL5IQh53pEhYWshtHL3QLepQKYiG4+0OXWT7DSarHY2yk27iY1M8BWzRXZ
n8RQddkHVGy4AZPOCocwwW9rZz2SqJSOHaUGnfDxCQ73kf64u2XO59miTeq9
aWm0vJCpbe8RnASjMq0pIpXWvgdXPRdcNtf16fz9chhvFBIAyNUHAfMSJwoB
JFKOPXC06i7onFUXH4gAu0KW/Q5eWN3YptsmwEMMyHLrJAqqmbVxchBd7c0E
tAS4aAOv3NvpWSVQDDZ+TjtDy7i4NS+j6Wj/pD0urLzMpAkBJoQhW7drBkPr
znNaS8kaBsvmTtgeLt2Kxq7KX0eeuqZU4mds2tWNhtGp0zxQtHVuYn1P3Es8
NNU4IRCJ/tQvOhvgGHAR/e/P66HbPygRm2YPnyijXyuU13b/QrB+1BOFxOY0
3CdwhY59WeV0LFTHW65hbRoKC986JZ90JFuszp4B2ocKhT4mgUqF3zsiNZ6P
jBpvZr1vwvUiQPptOQarPkluB0+0gRUPuppT0x97PYTr05zdXtTOoYJB3Jhr
iYj2S3p8vHsGPeVVG6UCEiFNsa7wKAEoYpVNZpETw0BSWE5d4R8bwhmu7UOG
NweCvDN3XcIrTBxQP4v9cN0zics4PaaG4OxgXl7Ji4iOaQqb+NomYfA94WUV
F0XIN8vr9YPFOzZS0joWWrrqlZeba116jW2BBvY3CiuQ74X7YuVuqrA8DQ/B
CqJ//S3vV0CMnpgQ6HJ7CmduXlQtfjgeBvihFHZ8C5cNleajw/NSFl7Pb2Qb
YOTN8w7fg76TNq+OsicMEaMYX19+wIfAfPN4KgZaLoDQr+oEbcHFKesUOiVM
aA7afzcjVEVPAQEGyLM7a6Ebs8nshzszlpOy//7D4fdWnGae9ZZxa7dkPaxw
BP8fX0SeqVkm4BP+3+zFzagbZWiv+HkS8HUQ6eCDSQHj/TQMOitRi7/UhyFz
rYDz1gnxyCs/0bbGszWkIVGYFUr7PdqtYzbTZM+G5rzVMnP04uutcsDC8J50
mSUklChEftOtzaL4c1/srGHrLRijmZVFyiOr/r8T/Jp1vkTKLeHFG2s0tECE
WpPsekKsiifazpzHuF+j3fUg/CsQFT0H2BVa37xhhDVJx0hbTdTZ4StvdNln
YmxK9i3ckRCTj/xE5GIIXychPdyIw9Jl/LlUN57zBOGLnG4iHDeDT93J43Bb
yARXHKmpUB3YUFOIZHPv32OlKzMoTt3DD/v6AmmVGdYmgzuiXP/n8VTB+7vt
5ExYVM3wJSa/Y4ZNXfv4bbbFVEKhgigI3aLs+g+J64ogJWC3VFfqf0U/KyHN
cTYCBNcUKxCUSlwOas4C6Nu0Ay54Gw8gPs42qaTfYiEEflvFl3yq3/myStTr
eD0/MPm0F9owN9Y54p3yLxw4L0gWlvJ2YESd+H3HKE1JTnmwyvnOq1uNeE2j
peh1ud5bDcxH6XzaL1J0MjTVYo/ShWHsychnfrloshB0L/kD9waLk/iGYdzR
29RepFXwnfkf3DpoL+ApDO0u/66JXfgzht0m2sHiCGH2ODxp/+qW01tPE6kH
YTDqMWy2nk88bxw63G236R/kitqDr3GAqlMgRfigpYx82xkHhe/OnY6uDqeQ
q1iJ3cl7wMnGm3YumACo3U6pNTqoEHO7hYERGYrfX9tixQ8rzXUy6K9WJo+P
1E2qmNnN3/7u7+H5FD94cACnqYZXWVRsRDEW07fQVhpsZEyWs9s7LwaLbkCV
LyCzz9RgUhBwUe4eZylpyEs4OykaGxn3nf+Qfb2RfNDrEwt8JntFD/icjtX5
qrUnJn7I47ZwplxAvPeXQkXWoHW8ws3x8PWjLxFo3SUXJNv++RMkZxl51h4/
Ldckp8MJpjEpI9THKFkqoTM7Rb/UexkVnLCWgDXfNCdQ9fB4Ye8aXo3PvKaa
YnGiOa6kfRx/n98EOFag/J9GZFSDaFYc74JrJmAK+nPjNczz/Q+WXiK4Hd4E
bsNGDLtAAcaANVyc+HnFqdDC97483Emx8P5jDrmjtPC9xLapz8lL9Ij2cLhs
MsQMX9iuR2G6G3UG9sBPJ6BbHuJMi5h8Y9LzcccMjLjxZ12+OcVgKcISNCIl
VxfNroJVFb2yaoECZQqKa9wREgucybCfvFMVAjwADVZZPl+cjIZmXrSxiQAk
HY9t1oCTG2YVC65JVUJ5hQSRNHPRZgM/v9cTH0Em/sarnSCwApGzxNFi/a5A
suzyv8LWhZ/m/pb7RW3U+RgisaFUKsjnuNwSySFqD1kJ85FuDdaW0qN4hqzz
hZHyljQ8UG4AJDiUzP75bJA18Zw6yZye+nchjuPU4pLl0vxm7kNgbqQYEvPA
NCu/KGwqrIWZxcXRQ6741rnMs96ewnUBLgondM3Zxd67oQ2AvZPb3nlp7+qI
ZzWJ2NrWPTde2x3Jctp4sUGIU/+Zsq6fAoAgOSaaUS1E377e/2n8J/84YTpo
ZphZzB5t85QorUZ0cVA3+DC6qqUVmNYAbw+/nvklZqX9FJw7hm1ra8/+ITPg
kPhsE6HessmL4UA4tskt3zX8/bHoLjGdhN+cyY+VhJL+ITO7lQfEXQQ9tlfX
rOEOInWulQtyAbJNgtWUYkdkY4DRAhoPkqGIetjFVM1FtySfkJwT1mW/6xH+
+IpMnj6HttsEJ9KN1e5SfSJonlfPK4UKXml3XPeXeh+ZOegF+3JeSeeJFaQj
SIhcCZtpxRfZdm5W8vT1Fiaa+9tSs8L0mmnVKmUUzkZ0h5I3pskOhVksTtbk
6uYWrLoOhCcCIAuK4vnqGOCnLOpHgS3DLkdG944Ftf0Sl7mLFxYR3c8wweQr
uw2JTHerE7BZfA45lMa/m0XkV2ko3QfTyye+FR4BHQuib5R4KP0H/8J4lCDW
gzKLc3mMhEdvKl1+bSfGw5Oyz8nUXdFrg8FvLjqgy5BsTUk7v1laan5sXRAi
h0Lgu/yJr1Bat6s96Y2I2OEKfKLXzokfNepsdNdWCAq7BjQl+v3iCAn9bTfZ
6ijTfaQ/Xk9HbdI98cy+QPkwF8QavHHzogazw9s3zDTdjki16OOPv4EpsVSG
fBD/7zICaHyeVt6NBVdIjGExXeNMOrcXF5pZBq0JLYGWcCRnK2aUQgDI59N1
5L1h6H+y0FNDdVJE0Ba1/Zb6fqD0dsm01+6tN4y2WYZGeFgK7OITvHKfMvh9
H0l88Idh4MPRox6c6WEeem8A9O6HdXTjbgW/JJP7PbG2r0ETr/+jOMen6kit
hMwL4hZ2Efnfu9udP+nwYNuF2boIAv2eUoNZL6jOlJu60KWMF+X7LenvzJ8i
pR7PIq1y8UQzIIK/hgdSuGnSEvvsBqGfpTQE5U8cBJpbumKNfhgj5AgGuupb
Z/WsXo3IotcLvnPSQx1Glvw/14RxGTq+9CRyzJpqu4DQfGZl40Vw0uKTXrqp
c6fEky3QeWyJdLPC9qm/seaWS6X6PDC1cTClbSKt5ggul4kfhIopoCs+PCZ4
jxZ2gVv8AWocy5muGBGeXYxXG/cKmcnuOHubOLIOJhPabQwNh1Lt+1UxTAwj
kUd7FyzsVw7DGrTj9MdQMXDCRrrz+jii5ihPaoDu7xp2KGy1I/v0l3+qMhEt
SQd9WlUZxM+Hrx1c9lntRzmesef8pWJGf5dIRw12soh/ZyBQgDDUrQLHQKyv
Gu0vlD9EPsebEeN+cH2QwXc4aM5ch0LUwpbZMw4X/EA1hhsQrYCXIXgNnWxI
RWlJeh8L09LtbgdBAWsYBWA8AeDopDhFxN7RhoJ/C32hoU8Y8C4KIaJc2VvO
YYSlvQkDmFnxp6Mn4RS4aCofajEQZRVfiYZwdmdJvfvDXXkJqIPMkgMHkP0G
67AOKPWzk7pufV0ShhCTrKbI+x46df3bsc3j9MAkIxRo4zlpMa73/5AT1+/T
MVhdsPI8I0Od2Loh14p/2i178E7XhYxblSVRVhFD1L8BiaSzU0zoNk73R4u5
5c2GebUzOI++aVOfJ82PPd00POTzYxUgznYe08BkoweGIphL7mrhm4FVAr+p
vGSm5Zf3xkbzRkyJ0LTmlLq51WlSwkiLVxxhxAVb0Fa4+0XM0fBbJfFw62wR
T/CJthfdg3YllcsbMo+CowYd6ydW4Eb14SikSwdNP9r6KZv0TmcyIITLcBgC
LU6zV+WJX/ODjgl6MhgfyB2hGWHd+p++0vx1Mx2sbtbeTlGRpGgQwCNoczN/
Rzzrg3ipijMKyxEIjV/V2z027u9hThKgT3OqG/v4wzgE/mbQzQy/5k5k0Sgw
vTSnNvw095d533S9lNq7l+1DgBwM6aQB9MVKi2Ot7bkD7MBXim+kVeF4c+fC
ZNdvRl8WncLfjGFyWk9oIs1Dq2acbXMZSU4UelcTEylKTwlgII6V4tUL/5wg
eDsg6yBeY47QFCJY61/r6nhOgwxovy3alzyA5rBRevt3858R1/aNFN0SOgdf
WXF1qCTpg74L/rS2EGjT/lIacNLvAQhU/x+JMUG2r6x3ynvV/8u7gfiAd9Xx
ydW/kL8pV1Rr4xRP1ENjqQxbXbBC55FaECZgbOLFK405Y9oV0NE3+uMSJqbV
aHodkuaOfAsTQaoWkC2g1gmYLi1IJnvD/tPmN856D96Bu+nvgQTG8c243IUk
CZDKruila9vVRk9uDLXagytp4Tep7C/0c9wVr0tV7N8c3Jy6ZZ6/Nheup6CG
hgK9u5/Bxbd2vzbCpXCRr9YcHPk2HIn2ttGn2k5b53FQ0PdyQJTILexRBivV
QAh94c5wjjm7iJazxRAehiFIxyTlR0bc2vGGG52CmM189jck4ckMvf9hjveV
crWgXWqpF3C7cSw0Y9uzDqZctMH4cwmzM3OlFZiuYyxSK0hDENxDwX6elO9j
rpuw5SBvWZafd862TGnGW20rAUOv9zj5iFcIHmJ7n5pnWszDY2cPFcAKnJVq
gYWCPuDTlq0UBmgR8phVDesSwRJsEYHdpztP67C1gKwhQl6D/W7+z2nhhsvF
I6BWWB1+wf2VGJ7+czW9FGsUaGf3vqTDjJG726Vstd6xOu8yXdvNYl2BGOwZ
drNtbn7u1JjHIf8tzy7ajYfT9+CidPWCa9hBufntccofX3BzdODtihNihQdP
ZPGoGSvvnZUJfJA2Fn2eOywsDitW3huta4jZ7rsUHz70OGt3yos4rd0HAVPR
IKLw0EsjRsKQdbLWDCemjEay8imGE/MXjiwbfJVQEi2TGoVKWmX/s1UnjPfz
ELDclU5r968F2+6Wx3wjsmVYkzsXPUBDjex4SIbtnY4VZYYbtK0Gg+Ylun/1
xbzztjO09t136Zuxu2mBkzcDT23oNFXXZyvqsCxxDGiVBjulJsoinFsTtlK1
9kJOPCbYh6ghjQtJYxDvcxKiGg2Hox7l3TjAE4PYfrvMe9Lwxq5oO+eeuQmJ
Csfwt8bNce1ADsootGu2z0PHD24K187pdvRUKxCmXn0txq8QugXMzJ/tF4JC
/2whNgDm269PIS5DCDI47bYue9RNjS1XHZztbELbWYFncfsVt2kcaCuyVdyE
FfJ+OdnpmLdquwlHMYB4X3CRAAdCXFL4KDqOARYB2dnlrCiFyB76IL5KGCQf
sInVM1Y/rU+ZwWjga3yAvFFofwVcBlZl6rBjJijDRUfNOe9z/hnjtb3WlyZl
be02KbiPlbvPEjodxnOXnp4DB0z1cindGQgd5AynXcZ+2Cs1YadkgAwq43df
qRhCu/RZ0H7YkFfv8dNiwuFgQUrWzsOv8ByxrcDjOSeul26HbZ77PPIvyDR1
CyxlyInQ0Y2gqTSOq5UMWDqPd5ppMD+w2q8ccN05+OAPcf8nYo+VswnaV3Ri
nNMFnHFl8uWBwmVmKQyOX+qxpMTMCKPDJoWiS3b4F0R6xvtkxbOVJa+b+Y20
uEvam9ZPGPRWs85lsoZowoW/YLgssfZpztPI/UPsxLCFJutm2fyiJQ25ycb9
EIUWxJJRcbKVCRUIdb/tt8UBaTCBHeTtkhDs6bxgd1JPiZvltIO6D9LpQVYK
TwYSe9GCvapDB0gRD8MGB9lVXUXxaKBSBivdQ8ZAmXKHK30Jif5N5OpU88XW
5rX/45TuDl1ckn6GNT391PzLvTwVTIwYzpHStgvtix5hxdwmI/rJOkxbtzwd
+DKPz7lQfMbXlY3aj7wu3TK6vUZVq/pC4+bB9LvGrj7NkBCtc4+CwSBycmA4
S4HoqfH29RC9OBcRSQr//yYDdUsdLlVI4MkixTgwVKc/pN5Z4jsEujg/1BHe
NFm3RB8y3jbP15d1+I1RmUKJEM+fHodVhBcOE96hNO/JuLoZVYu+lqD/uoZi
aEWDPZz07h82jszyfi7h8E+MUDs3hDqwBWyW51oRXBLjlx7uuNpgfJSZCEi5
XN655wPyIpUnCBhwoAVNqXo8m4LAY/o3LHYtTvV/DIEmETzgCVNqJKmB4ZCh
dHOwD2KfzThm6wWqT2wr0qBAcGMlQqFgKNfdTfeFw8HvXfhocaLdifjDQGIc
9V2HBiAkBTtNixsze6sZOF7Z5NcfWAJzTPdypJvRUzHPfkwlJYE2zyK0Zh2v
0OzcYnExCI/RcrBnO6671MPzp1duvdWn075oyRln5OFN0u9GRo4/2iA6iBew
v+K8WHv9rPOjBTnPAF/YTEms5YrV6MBYdFZxffwkmFs27nL0BL98HP/gsNh9
LQzxxmt5YRLoWMGlZOH6aeq+YC37P/aeaZWIwciUZFwrFdwMNzRMdITuECzv
qicEXj4ZFG9rYuVXrnERCVVyEWXv9HQbM9h0tklFXJRV4QnT8uPHtkBXRVM1
4u7cz9Yb2nTi0IE5Kh7dfkIFxcd7/PJtc2U+M0DIx8RlUQqPtI7q/W+LWo8z
rVQsbuTWKhaU3t5Yu0qKEXMDOqvTL0km8ODMjDZj7V6MC8s8bvOursu7zB1p
gEt/Ld968ENkh5RFCWR0G8nvMWx9w8UsxYK2CRra5Ger2NbLqXdILY3mcnSP
D9TIu/1qwhNKAIpE21B3G9tEtd22YukrUnZn2g/a0tIN2oYUFXrs4Z+HjVt1
0uRwBcSegIstY14K7a6MAK4rHI1bk1NYRI6Lnkbi4LEfQWlwlF72JEBIu0KI
HjmqKv3ZWEk8rWDNlkOhHkXn4Q6UFITrbCB7v3xDV9eqy8/+QVgqaRWQvjsP
AjOulq2H5ZK6GFyWxUkqUAL0of2aRjT/hq33qCVSiDsesrXeW2qvsUlKxdD6
WJrAM2AxZpV2UT97ab7LMu1ws48lqr3hwJ7ZZUZ3C2wqgIRLW/JnIB7wTZQw
VQLKGhzh4ZeD+gv/YaXOi4uS3+OxO3ke0+XrNicUNgPogxq7r1NiYGso8B7i
mWPbH2rSexmFSQBKpu7FdZsLgxiMhzyg9zsMjrnDUZPkNoGGjEztu458p8XA
QDD+cdb1UFyoKMNvEAWRCg7QQXOtQDO/MQRdw4yaulIqoSTqZYFMS5vbU0ps
UpKb7ayNxPCRUQTH3srjulHV4xsvFlSpbhOwgW2gHL2eJRp7lsVxI8ivGo5+
bpI2AAneW+9Gxj1PbjoRvD6vmhREewav6wfdROBO1GKt8k2RLqGRUphUKyIY
ZekhfrzHp69hduJ4HoSWaZtqVFZpiAPph5y2l8Buo+tJWEvO16xG2GKEhFJL
MZW64KbZlq7w0cAAwlW1nkdiCFV71vvCnlFkeuYTRqUvKuzZHpiXmTOKOuC2
IaneZfS1hbATuMoJs1Bc9Wtdt2CiqfjUO3/VfZjYCWrCQZ/Nw6NkTU6lswPq
zeoSNzwgh5+DRPndvfjQmbfSW/Q5bxP3F+O8gEzCayytIpj/rVrj9PhftGDu
6ZXvFtoW7/CGUGBfxB7DE/nD+6sLjSzHJF7YXXjV/c5NC2Hm33BQWG7rus/y
GggpFs/tcuvJ5zrQ0iW/yRupsaNjnC3MHWYbTl8cP9q6zY1eG+lo/NBnk7nE
sw06gGMS4RQr8BtLEEmRP7o3vjDwdjd9Y2Ic6CFuqXoR6EwxYAKz3lQy3ws1
0QZmF17JbP/amnISaPYK64IbLe3kHD6qFp4nQ94peZ5M3jzudqLWDGKG5qbR
KTJLvUg66WMBRdjBzeKyj07XJpLhQm9sZmhZ3W44tNJSIZgiBGqRyskumt4G
4ElSinRNctmUtRyl32ZFUfWSTc0PFdOfuVAtxzCQ+GmQKqvZxtU08zQPfI6i
AHK4+aiaNeHc+DtkQJbQusJ+dXqu8VmRht/wqGx4kt6aMgC9LI7CNgKfmOdl
yazQ1qBSdWUwZzVcJ+XXSrkt/I4Ex5t4mcq/vEFoS8kcMTYoSz3eXl1a9ujO
GetzW8Rb/2u/3DaxJwJ4RCDhBL3FB1d0dFqySlxyunSWUslxnAQ88EWwqcjV
TjjMbG320HAW9yX2S2L8q9tOwpA/vwhn6bBY3bIDAgztUfKPMcvo5Jecq5XR
WdFH+PTxpKlqpavBo5VHylDxcXmbHwfzR7J4bGHXoUh38e6BrO/5la2wNd1b
li7o2Sb9c6nalKjxp9hpINHtoTcS7HAnKCa5vRSji5j9W7Cm80pFu9I9ir6v
0STzMGMI/HZp97BU1+kPn4rtMFNayksCS2dyLUDFoLW6Oy+uJmL31cvHw0W5
26+GnprzgTZFWjwhZQiRPkTMUCbh+H8b6dqymiqG0gNqf8IQVWguYll2Wq3y
UBOP6iW1ZtRViEegBCxgOa8zA92vu8+3l3b4Cj4O6l64rvvF/ppODWYQlxJH
Ls8Fj7KzeKOn322uV5icl3zmHwSVtpCGuQDL0aSoxn7v1X2A5qu8tlLN5mgE
Oo6DPDhNoCWV5HtzahuTKcZgW+pCxxz7lujYCLP6+7ku9PVOVveRu3Ve9H18
if16znispAXY63x4d2POq55JzWcsBo1r/WrXrZCciIW26jhcU6oRihE5gLul
nkY9tT6E5YZ6AyzwOgtbANHU4EuzENx+u63+x2znpjVhSnaidoAn7XRYJ/Xc
27ef/sWhO3VMe2kVl0piXc9teSLJsi7GiDDOC7AFwbfXML52fGeNrnerVqA0
ux8y2u/Yhx+71Pz5h6oqV8Ag44SBqcmkgBUP/sFpjm0tqMYcL6GwQ7lWl9jc
QsXduKU/hHxSCFxr/ARAEaIy65pijjvkrzRESMsKfDn8+dJ9yPzRKntI62Ha
ouuB7M2i+esNZiC4DnM+Kyo9w6hkZRR+OG9iWuVM4y8/hiVlNl/4TplFTZej
TK7U/mbswjfF69cs2Zg05Hebp23ETDsKHuawMwwR9gHpl0K2mNVpNdjopyXn
unnl3ezzieC1hv832vGjP2G7UDuuizu5jxEGCH5g228PB4SYfKmfSuTcKRFq
m+GGR2NElSW9hdREpPcEsZqPqecyp3+mCNoKBXPjgCetVlZJYN1s27wNr0TY
/7K5Dm652R/bK/E3dy6OH7HkWkGUm5MbwbSqpAnAlmX7Vd8T6zhlXwkuzHzh
jnrUfSOdR18u+86+5CcWSB20M5hbTNlDCRDSDWu1iPSBCSzblIR1OnUOOkOH
jk1T5wzzAksQ5WIA2YP95R1ce1BR5648FnKXsNMUG1ouP+gObpMKWnMuxqDu
i2z25Rtxndyoh6NakBBXWUNkJtOSPekYeH6PdPYpowZAoJVrzPm/sArfQHPH
VH2UuM6yYW87lupqr8tCyjcYs/HwD3Q9xgVY2oiVOEiAF7Pn2MB1nrwhu4QO
p8k+UCcDsTMF6g9pTV5kG8wb0m8v

`pragma protect end_protected
