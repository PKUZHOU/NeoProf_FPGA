// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
FhL4KKeUjQkYZBDsF88TzHeApxd0uZQA+W2pN9841EcM6gXhOWJJR9Xt4LM5Lwuh
fqmbE/AvzxB6BinbyAu1JA0zLZcSuEOsKfdhHddBTQjik0uxWuIAGaTFpNzfbqWV
C0Zw/3zu5qw5Z+U2Sckua/+MQSX+GMutXhJCjOw1XIFcU6UV5LObhw==
//pragma protect end_key_block
//pragma protect digest_block
CJkiVetuqjAFIWbM4WYdM9Nw3mk=
//pragma protect end_digest_block
//pragma protect data_block
y+fZG9c/pIoMwumyHIUqhkiTmwZlE82hdvElcAf0k7L/flCHNYc3bVEZJpMJnfRx
Jatgrbp8OEoVUY6L1yALj+hXCbPUKJ42ihyMoclEPQmryzS8tzB0VYmV2Hn2FI05
dBvR2hzdCmAs+W2tOh/WXBtRJTLQdqE2Ur+BsNYOw66aPH4Clb3iEyB09f8IQDtq
Y7SfIqU1NA9nSCAvnNq+9ODfUOZclL17bV0/DsNTsITxLPmHhO3lmFN1JmBtvOVy
rCYaOKZ/MUdjrfTrxF1bO7Xj+obwrNUpqr1svMp5yecz7hUw4unFNf+3nWRUXodn
HC/vPzGrRLeSRmxtOzUR9+p0GG69mm6IOJvoHuFjd69Yzc+G8vqsI2wKAVvbhXqb
sxdbY6hkmByePNu6pctspv8LbTZUnDztw9TTgZaonbU3/OTlynzzf/8tVlsNfkQv
cuubwlnTXUhACRu/iytGxr5/GbT8TkQe8DSIsODgMGfHx6jRFOwdO17AczVkSXDT
BH88ad77lFNGv4bbN2hbRwcsvUxjiXGQB2kKZhQRLgRr8feIgNw0FTqPqjMjBvTp
OFWuBfcrhC2EXM3IuHXfiN/Rn9tcNjJIMQY6SDFg5/WRGyDclJj4e7V1EUyLrlYV
IUI8FbPSLkpubhTs0LKOOF5LIkhm3QFrZyYozdMNyEU6TEu5/9sQgwUj4ZGQ2HJg
VVYcGu4KUU/ctTFviqMPBj/80jyy2ZrPAABPfio0ob9CcfE+qA5JTm51Mgyd/BYP
8guBsWKoHnyy7tYxUFLXFBgwpucSYSaHSca8U8yVGb+kDpYPHcrw4DsniCNgcq6o
BGqRlX/vCBfuegwHJZOxy7BucoE/XkImqjAT4pQhfiiIqQdWhfstRTwlEBAelKyv
JKnJT0dw7gzMbT4q5nq/Zd/aKLgYKhnLYd9wf0xYRgILUOrt0iJpsEHkgPEyxhmL
NvTkG4G7e4a095o2ojbKFwjxCqvgKV0KnjuS4c0/di9ckTX8O0MNQ6t/J6W0FPez
mU6c6Vz9X2/4+fxTybQIf0z+hkR1nNMRMSrvXvs6EnaaPrs4g82G4WHnjn03Zy8y
EVZsO/Cl3cW7T3P5tS4iegLYoRVIT4iaOtiACeXMm+8ZrvEoogEktNIzTLoJhE/2
Ho2nprjp740+NtczqXsovLckxEo2hQu4e/BG14gESC6Sn+bmqeObrjAgAcUkEV5c
vpZczrePBeACOuZiu36rqD5oPcFFADqMdfvANL9yZby4AB89nR/Cipkq6wZQxJrX
rYBTMcsFVVbvAwE7kJ9TLiJaXKN1N66tE3hLujLwrOKr4nNhFTLJ+9kbKjXYpgtR
beM55jd3POrKTM9Sd3lMNzRQi6u+j3a8xxupprvkeIFIc9lrpZb6jMbw5SdtdFH+
AD912gNOVjgDm4RFYFY2MAyxfruPj/ZHIOc2cnTZ2ZJpyNG+WS/cuc3X1c2HXXvn
3+xvNWrc719zwCytSOVurlbUjQ58NqtqnRnxi1XjH3ZEcB1LlC0l061sur9LZZqi
kCfk9nzzUqNIHqzh1i9vU4nadonXs0T5HAKQ8LCi8s+yqVNQeXfVOqpyzSZlY8Xf
kyfherbltp9otdmIu98LHg8OSaMoxyOn515w2MM9zjt4j4KYNjuJnPHRM02Incpp
2cielxoZRAZshdOzegUxXZG75AjFzSaf4auxX3s0wI//LY6S2UzAWsrgJpCx/d27
V2UBrxAS/wFN7jomnPztqpwwCTPsBs4VjQVQcrdbopq/mQa3MLvVGwjX/o+CAVjV
pNb8WiHKyeeI4y1UpquF9J3Pat7JWsbDH0RKV0Ihj4B6ffgLGn0T+GllBQM8zq8p
VFJWKIevp0wBgT3DZroPqRYyYAIdfX+vNIidWTnUWhRrghHIEMG8VxyWiNw4a2Ex
0GRVIVMd6HLjSEHUmpc3tR7HVFGhfF8S5NbiL8LbHb9U8RimVUIClbudH86X65eQ
LxVUiMp+QDRMl3VrOp1qMem7PWZrQBSOflLy+9MhHGV6xJ0RPlkVKwZnAFZXDOzr
fBr2izMtJJDm6wcgz5YbVsPD9xfMzVPe1BzJc49EcZBoUIlpWseBk41xaAlcRUnP
I0Jk+m4alx9nEWTZ1+y99/uoElSR1h+HdgIlQntZbDC7gWhue8aeqDaPMsA8M+Td
p6N4byCL71xbmVep9uAAXTmDAC3iv3kuXndjF6kKA4NsJ4G2CAEWrFgUZ+SMWr6j
DGq0BO+Lyznkg7GK9wXCSQNkkl6CPak2DiYB+QxomOjGWPki1pD+ViaUjwNMAYB4
2KD+cIU3nqvi2Ww/LDLr9/O+4jIUeOsoWajwRKZyMitthZfxsmHcBYoJ+4JL4DQN
dF1G7PkGQxKjrFsLQ8oBYWqdWKa2ZmGz0TWF/JzE45vVSOIvZ0lqJE0gQyHiyw+b
Dk06kEF1d7dKd67Y29WMJLzIpwY8/5NBVDGsunyfOKemOvMcKMsWZsq0OENwhh+I
WUxjf6SXpx4YavqrRMCekS4rJxjb6nxzh3UxvZxoyRXa4kLa+ncANu3dTnYJH/jY
8fQ5Em3ZJxNj51vVppk6+JVNGnJDfFwrLpH5ld1YhKlOhabVPdhvYpqgDu7jG8Ba
CoDLU3mH/Y7H+Rcom0tn5IhyeVRh/U760qAd6QTmGtJnqh2XGPqy8PbunOF0/ldn
Hh5wSvBCfF167xBXG8kwVNDBkBqcUg7m5KxXp4ufvZFmM3K/AsJ9lEhI2bFyh1R7
UGhkwRcrco5Ee6YhtkNUGR/+JuP1D/D1SBoxPnvwVmfmJ7JasxhzDgg/j6ifoaS8
foXcGatipF/+Ie0i3xWRw4mJDYOB7PVnaL2G8naJeTGJVYRUFlmEHsYV5i9n4xgu
D2MZ37/B9qjx3mFnS60zbDf1Aaik2yju/9392neeZsLr08a20JmhUi8y3pRuBPwI
F0cTtSGsihiRQme34JWVXnfnEbuHFSXGhheNtzyLGREpBuOuyUcKVqDi6ayvTfPh
1GAp+u0K7qSQ9jMDEVmlsayDjOOYhzdq8a8i2vGizxggGOXvtEkLO/DSxdKR6dO1
kcGnsJvPuS8U0mmvqiaScZaSBbmVnZnMpp0+C8ymLv1ApOmN0wXoLClfbVvw5BIi
q8bVuQivm4JzoY92uGAN66tKk5U8g32ZxiVVtaSr2CObenjSpReu/r1GKdiQtd4M
dtlgI12gbmLBatFX/ug6rPLI8HHH+M4PSnwVBI24qnLYtgN2FE9VS2/g1k/9AKz9
p5+IQyujdNJi6MBTE615WPGCVBidxJSu5P1k0z9ngMwTgTr8oxvX3llqk3wT8TDl
qdF0nNiXML0n7eVYrgS404Jryg4OLc45D4S4dwLH5yIcCNnbbLgisPxr8YwT4n7h
mWBYGc5/aYmZs3H3OVgYpKb6qLaRIZYoKSJuSCZidg4ivhbY7VwXgVXHkasEzzEY
34vvTiV8Y0iB86qeDfrezKMIbImk5pHRHt/xFVeUHFiZYj652aG6PS6tWqML+uj6
KW21QaIwkCyM/JyhLCsj1t7W4EB0jp2tsYScpVgdeEJVN82I+JViPmRQ8W2CZTmL
XNQCPVJXZ1NysA/NoAVu2Fy0B91FQncChu+TwOws0+8wJUwPYMjHdh5NSDCDmLW1
KOx2gD9fnIFrZalbA9uDw/Nl3Wp5XP1GjnVSQZ/BPBfNqlA0N/eextk1AXuQu55p
NJxRVmCAYSFFPyRdgee9gG3qZoMRUzugxA67//I7zE7Jbkuq/6w8uBbPZ4gb7Qlv
Tfzik4jvl7GpzGMcfWHyb8HGOqcctdC3h+I+8wXcumY8gU2ApRscJBbJszJjFCiO
OFuPkuycLuMerAbG0yeyYfoCQpO0YZvZpn0s646G9eZUUOhrZixUqT2dVNTzRIlf
03SoNKVl5d8U1d6N/bmQnCawGv8isL57Khf15uHABV0227IaEblaiJ/ZKOJnO4k9
mje2YN2kwMhe32sYW4QTDKhfRBZ+Z0Vf3qDaNutUOlDtnYeSlMwjvDBd8og0BVlo
o+uUyoCM1U/j28EFjXc0IiS4rdzpSFYplh056cisu7NEnA6L9j7rEZN1n7La41Ga
ieo80To9mbloNP0CfH0Wx6lg2klTNQfrc7MxinhLsdhU8lyhSd4iKHMysnpel/n+
QyVCJi2YEN7EJbmDG7xgjp0bjd5Iqu3TgEB2510ezUIb/Y0q5SdEgyCviqrCpfEu
dvxeJNKPUEdFo6FK6Y/uhRkjf5b7MfapFYG9SorSXfVqWEoB+xwXVCZI+5+O4jeH
yEznDlPbKtyaDlUe5ioVyXDdOlegTFzLeNDceLiJa/fUQUkXJL+eL2SSoVjhHvN3
B9kgLapaNrsTogzZjGI0Mo93pSchHbztJq/i2O1FbEyLgR5hZRWcaa7C0IrbK34l
fLGH9FrNztPXDunIS/+LPyO2eYn+g9sy/hCzw7BToAn52IugfZ3H43Tb8GcSzp+a
E7P9zWrfULwj+8uYWT7MAsHXn9ijAHzyFwhSxSdp9mGX7c7n4KVR08PnoLc1dptg
jQeVJHbS0smhKR6Pm6ak98uDV7NBiK3gk8v6+jzJlFhvJb/XQ+QMDWhi3TTqHptD
7lPYcMwMiZ7oBJgB5bZaTB+nywO/PeVbSpwegjlTlNxxJhBUClYJoqgbW7MCFqIs
V8tJi7UYtUkrYM0NdnpoD2N6weVGVGVPCIE/DRjzG4SXSfxRx44wdJLBahv/kIKj
a377Ba5A8yeMfUmI4GSe4srjy2xNvYVlortHJ13VOBLl1GN/8nAy9hcLhqPJjAQK
Bzb5etzg57SC/m4yRuoSrit8NI4P57IBJmqtTG/l7xSPcYqBg9SeDtnqU9+Sl1rV
/7JYXJdxurohKn1SKkx17gA13cYpOcN3ZqFnV7Leu7ifE9LelQsNHFXmKk7p4RV4
5FRBiijqY+j6XtCHjzf/kY0j0LugzRrXPRIa6uFxb6cUFjcHhVGWbGkbZKUGO11Y
BmpO9dS8A2LaXrY/PTOU8kvpa0M8/rfP+YiiAYPxj4HoIIMyYKWSocn/G68yPQpi
eUWDAF8btNC4e/ni1cAZ1OZqzw332KhYAClAGarrYvs5VdxE/TZtS17CA38ZV8by
2I6zW9VkMK+RYWBYB8btsI+YrHgY+hnNEJ8miWA0mRQWbwIxoV8VFb4Fci6VMs5U
qxuo0/5+wmTrsXBpewkIjR7ViCbFCbZ2o3bBiBeDr0pXTUn6lXH3cN/bXasQcvLV
PC8w44YOWYaKpNLWitu/G4CEnoQUB29ZfRQzEENZMM2LnR9dy3u2rsYcoPxhodAn
p5jPk3c7w8mMRFwPxIOjnf/bO3MELCJdUzRJKh4AGgcbhiJZN2l+Ghw5A/c5ohQJ
9CrJ0rmZ8Chx4u3CnGX3vmvpPqD5eAXAl3DvKhdpocFcAyeZ30g4a0PXHRWvva5f
Yc3sro3RbG+FWNk2YICGpzlVgNRR45LULydQ4xDeQI0BQYjTRs1qW6qZC4S9D0eO
HxJN34eG2/OXloPqpQxpoJIbonNNsju+MXpemQRZYiVLgEocSXgwnc68ASZOA56W
OqR6GLZ7mStjPSVDyAqlUvIfP8rz3jtOOA/Hge4SYkIl1gjT3NXDzUmQpeRj4TTB
nsSSGrFAoOnio/5WmEbZqmZbzq8uddexJ/1hPXDBAb0mnwVOcs/IZs0sVCjg6m8t
d2RVOPNhwGDGHOnFjr0p+tO1rXkv8AR2bUB5DFya4kw6BZWFvnUKWY+SdfASHMYw
H3HEM/v0BmhWIXoN0LeUvl5+fJVbk/7Zb7zFSsiWrGh9nh7nm30X6zrAmrPUDIo7
e+OCDBo73ysRU/NRbdzQY2YZjntdITI9t0FUxovpNT8T7ICyVFQfbncG6wiUTS9L
7Iqt+KI95YvBf2/m/4MGhcxo45ZYTXWqSlnGMP7sQTQFeVfSuWrfWUbLrHWHa3kM
6GDhmoPf1ynCKwayGrva2HilxQPzjDI/NUmzPVnnMvWBHOao51+ngOfYO+AFxevw
QteGzkJN0pBmOH4RKQ6Geh3DHmoRw4rG5uV0T7YLIBJUJxlGH2Nrv+g6CjFzTLuJ
T5uo5VM1/Zk6nTqtL7TxdcWHI+Y+7k9JMRzStW9UKspse05dgTGer2uc+Qo8kdrh
E6vFnN30vP2FuklQI5c4k3IdbzRUKqIFDIS72BlqGg1jwEH8yuc46QZw8FUlf90k
U9lpP1+obwnE9LwNCbTVhtDvunyKBp6829nLQzHl+pUm8kPiccAQTNsZ9Scg02O7
B4S4s1U5BL2P6ht1bhhmyamg18199uThSNX30QoCNCayJNTVe98aP98/ZuYz3P44
i82O9WHr9xUZZIUk0X3sIDbY8NHIvRgOnA44WpI2MAJI3HaylUeC3T5dcLop71CL
HW7Lt4IOXGJhzoJs2TjkGS6waI5ZYIUTmKsrwnzufy/BgW0/zmNDe+8UyVzzIflS
HnQVrDoLY0+NNwkEl7vuXNIqSmO9Gt0T9pDOdOxGzi2aIFPqB0XTP5Txuo207/m4
+7DEKF6ImLWcK2iXseCh9q+PCy4hiZyMDI9QdToM0DAgPvYjaLr/6erI+leou9cP
0+l/vPpeazyAAMuGLAVongSXvym5qlcLvrlkVO6rMRGh0GIf23DR08mOFa4L0dyv
pJKhjTUGr+hJU/P6xrLsGAT53aewyYyY/mui87DY3RS9Mxruegazf0maO8dY+vg8
08QzlTnEH2vFgpQBgNRCw34AFgkKuXBQQE2V3AEfuA3eRYLxLskI4t5XVeLm4fuO
rLORji9Cl9wcxR5f7Sw4vq4OPEY5ZLfs8bcZZFhNBT4TCOAZrKR6RqUGkcBt6Wuo
AQa8hkjNRoMaSvtq4KGRWTb4eL4GqAQMiBDdgjwWjmxIfKjiP4ip9dKNsrkSbvNF
GIIeSfbrgK4iwUdwOEyFozmsrA+StqDZawViFg5g9vawpLNXt/p+lHRyn0kYZlwv
XtXmyqOcAz6BAAX6BQiJVHq20ZJlNmSsjGLEbBQZ7Pvnj6sYAbxalnJwJ4tbaLP3
jM7LsX7tx0JwyCjKhH4NS4VoA6+Ifi3lvNCFqWqbJ+YPb2BVtESFo/RQTHqzim+F
8exTzVKW5XFUsAG3WLpOUaro1HmLZEmkHOS5+8VPwTR/7vQUAbFN9GDnEeWdTkkh
/DXGsdbc7pfFUEn+Tj45/Cv/4l6cEp9rv0nRh1k+zGn2sXioq9rUp3I0uCEcaoPl
UrROGOVKOPGl+SBKTrNWkJceI8fjEQ0lRIGPcvBtiUYWjljJMi4Dkk692H6EF8Qn
Ne3cAWCwBpJln80PR+EAh22ba6ERFv/8Qi2OuYtTSmTxWIjsIfCmD6+R6gvr1/wQ
9yVYVG1bD2/lILOYdtjOcCV6QLUq0nJ//vlRoYoKF9Jikx5GRdm+J/EUqIcL7tMj
hnd0RQr2WNSmOxMsC2x03mgbdpphuGGtoMpWWW1AMwrGxSaTufq23Lf3lyYHcazB
h3JLU38yQVlN+flzmEDNgZgs9qwnjTjsGg2wrqu5W3aQqj2VppSiKBNQihbeE2h1
7NlxFDT2jk1U0wOIXQrMhkotKulzZ3NACTrFbtChrIycG3iI6nVeF694wf0fEszm
MM4wVH0hKORjVcJsfzGRZYPSNShcctUktJJF3jj3gy7I8bQdVMQLR0qQRo+r31Sy
4zRHDoUcMY4acBdq58JpTRzDWUo3jsF4Q7TmQTS29L/cOana/X8quTjQNjIZ1G0Y
KpNnsDLonu9zcBNiybmmNbZZBSVDUp8yOX+2o31WuWOE1GO/KCiL/HfKow/cpXxw
B+ewL5kcJ40h/KMpvpNXFOXdYLrvJijkDUB5rL0nGJC2dtEt9DJIQi7kBFdVb3R9
CAKD72X+9aQQ6F2ZY9ES2LcFN6RT/uKxopzSuIGRwNvTmiw44Cn4p9TCXke+7iyA
HieKrK6Gf48HB3tNpnAQky5uDGkc/wUGP0hqA+EvXr/wPSZ7HDiDK9IeG9o6KAOj
9Z+Alazw96fpxTP05nhrE0Piz33H7iAACyy4AMGgDWD//X5XTtJQkAqikRsgs7aH
y8Dsy4PwQUOhKRdiL+/MFBluK9LSSCy8Wn1THYiMbc5OD+KU6hX75+ODY84DU6NI
Tk/HD9uT3dokeukfle+TN/Nk6i2YhN2CVXD2W0AvpJPIwSH4g4Xu6dl3aAK5aI7F
MJRwD4IHob37iB8B18jyTkevOEIVvwGyM7S5b5ODukHTUJAnQC4aPuder1vGn8Mo
16xkMj+eAm9PtfIMRzqAe/6utj3w30vGmeub3X10u1BZO7FzAt54aufk73QxS6/J
QCKHbqd1CdjenKyN5s80aCOlVUSLEvjyTWM5RGe+GdVwcfh0x+lPv4x0KGHddK47
jXYBWQKJn8iODoOIrGdWB3y5ozfQv3j6u/02kdTOkOijvHyJmKPCdAO5ilhym3Ao
hRD7JcF6GYF+9WrhNtvwtcSFWhnnuBDaWbUQjUKaK5zdffV0N02f4vV3o0IFzGcH
1UQoTgvCSLuYdk6aPUK9hNOI7onWTWlqVsd7vHppVVM0xvh1l6fs51BhJfn9YMgj
IQBAVgJ4j00KtrKBZraVPhFkFO5R69qE0b7orlmisNkwC+KFlxih77dnacPH+1y6
91wFfIlodN6+EuK9kWTm0+VjbRap8Mcg5P+UP9El21E6H50O/I3x4dxMC67/6+/t
YkwN9XiGaF0cCI1Zx0THLU2wFE9MpT4cu4QmsdD+y+5ozAj7/GpE4KJlBJkP3shp
2A5j3gnixrQrM7t29sGv5aG5H5rDc/NtDpaOA8DdPqCz05gAn3kyjJw5VdYWYHe5
u0V2VVM+eNtYDTvsOF83Sqxnd3grfWZ9DZbiItzpIcU78QSSxfGcn8M97hSCguf8
jTFHMqJrY0GHgF9Sfkruo9nFFklo786YoEtiBGSXnmgCgiK1Kg6VYkaTkYothQaj
e7nA3UrOpqEpZ79v8LiKjLPb/PB5KHeb8+pAjtnxobP7lDatwJpbYad4vSLRAybP
4/rSDlbx8gkLlYbtWBBMghADL9htY+V8wF7Dtha5P1jaN7lVAa7GIXeUdXkjlCiv
cF/qD23IQP8S6XXVdWbPIazHSDfbVJPQDcs8MAo8rs9kgSEETDKco9GcY3V7gODG
q6WriK9x58/8QpcbJXoc95h6veIm+HXoRzRBMUvWBPDsC6eqWhOFNHSxfOUpermG

//pragma protect end_data_block
//pragma protect digest_block
A45dFmxQdAsHJ1X/kNGETQtMb0Y=
//pragma protect end_digest_block
//pragma protect end_protected
