// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Gf+BncnLXX/ygM+ZPuMEjGUL2GE8I/3m/sT3oBna52ejwDFsCK5vnkGIX/Y2zJyE
NyEdvuIVy9q7OpOucoAk5aStWi68ylanQOu1mPuvHxwPrlBnpJ0TMBVbzH6mEw07
8VIrkyi8q8sdNenJMZ8gZd2nUWNBzWpHC4gXJ01+KPA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7376 )
`pragma protect data_block
e5/dSKt8d2hifPbC8T7lBmoyyCcOmbD/xh3vjNL8u3dIphZRl1C5cItaj4YYqpmO
dWA2FgZgJ6Qi/vHBpf6IVbVaYujrL/h2RN9SlUXP1aDOLQ+Ydz2D49oC2uugJLfU
9Zs4Kqs1QgSQKFq0F/nY3iClaovEINPONOe8Y2pwlp91Xm3wxgVxe1H1r4IJhJZJ
dwjd+d2ce++Mz3ZK5Yf/ov7tvVislDleg7gY0OHpaXfpA48hzhtFPek2lrE+WQxX
FWuobiZNYJm2z2ZbS0VjzjgY1pw/RvYs7+jZc7Q0PN7M12n6yhKqfGeWZU5DWVyM
QFUHOpeQNRba4E7YH6M5Z4mda2UeHHMz8LBDMnAzsA7Cuc22wKQusbR/3s4hp8x5
L4NDVfYpjKPy+thUgUTN81Yv6cBEpXr4EXZNpoFhqlxOh+aXhiyPgT9ReLykYqLh
1cUWkbCJ5PUWEXP2l9gpFWSWVybDmQHKCERhVIw+6ftpZD4FI6Pw0X04+2UIpNB2
Yv+iN9rRsP+0KzgxIK7n7+2wfDHBkFGJ6gXg1ExmXvcs+p4cVTAptAnkUzfWl/3p
+LlwVat0Y3DVPSuMdCG+KszdfZR3GIhvTtPuqPa1rSzBDV0LiWlaKAAkhIHSev7V
kZZQvEiXLX58gaetJXmy8tG8u6WjG3pa16IvVVm80dpuYxb/Mq2/L/1+wIlV2jA/
CmeUh6sL1fU+5cBK0NMUkRetCRIi8BcrH7ufvFNvlHkGXGSB/bxO69aTRPkyn3fD
H97z8Abm/pkeLnoFmFzREpYw7L3szS43FsKhqqfTJfu7CatEOPIULFAFUEYD3k8r
0vUVvKldv+I6c856WNsTG/xk9OLr4mZN5f0C8x6+YDwGhS7NJmhxC200cUxhsP5e
+DtV8fQHutjFUMPPj8CFAFpCkCVUJ+hPIy5uRpOc+5nLAM8RKa4KapwYsrrReF59
V/rV2efMpzjyqQYokNpZxQBr5aTI+jWdUHbKFbbYeEJ0g/v+Eic/kzE78+INQqwe
ptqkzWwIUCb4upF5f1d7+Euce3gnrHHWGHX6JVUg0w5I2qyTJtIUXSys5sPSyvCV
2n5W4mzGFFg0Z3Dctf7zDkWuoD9wdupGSFYKcuP41k4dvHcRmwAGOhDynLhciTJH
j54OAKuwlGutiwplx/EmuKCcJTzogJQhuYY1U+Ss8e+EJlIS4lamo+t1FdTxxmG9
jKycF0YH2t16OYakG5h0nXwJQCP43RVNavMLLhHhc1gP8huXdnhljmh1I81rabHM
QyJb+F3YhxIqow1pDxZVJ+AR80AfM3UC2QJS6HKlBBJqG2QWlkC59oRr9ycsdGcT
xLTyX8Fln1TMyVwUGMcxi+tI2owxcLVvf6LgVZo5DS3bbdV3x59qnETmc21iCKIO
5JMvURUORB0sBD2qy8MtX3SLUhplAvWrehbfrI+yCizJkpFnN2Gr/IGvYZsyvFM4
LhFtuWx2ZyWLuVYafZfLjwkMj1Bq8FRLap+oYYF+7082l4Dg0NPsJddVbtpcQJbO
6bpW/H1Zfu4K8vQT//CSu3xo6zKqjQgfIroC5y2EdBXkyeDXlnEUu/120pZ1hI2P
jnltHCTpn5gZRNBdquofl/Ye/RQBr8KWbEzaZbOrhIfeqlwgaD7kWmb9aFTV4IGb
5HlM5ZBvQmXmMeWcbKuXnN9knMvWdcEMDcmH63mjL1/0PcuJhX/WqSr+MXSewFVk
w6NegKGCD0Z41uJONNsIC/R/Qdq+fzlSZt9XSn6wkCFfv+COqfr13Xdi45uRAEE5
+A8x6SOuWYI1XBMclN20NzbFviOsCpBr13GosS2ahSXNW8+Pw4xT0wrwQwLIsWra
WOwB8Yp/RPp5HQkSt8qCijezLXwwMygILvL5cmx6XguESE4vEhh2J0dO6qLYF1/F
dWZACa9LXQnw2KNxqD206CMEDDQZyLeZ0581yJ3z+UxgFpVOg1iawyYC2Og9BG1/
gZuH7rbwKteDu0f0nqxFDCRekxFB5zT4mHKszEtSh3pdPt1gD3ouM+6t1v1NVw9i
uw4MVsbPJabNhfV0KtzljnvO5fgfG6gfLvs3qf6W4kO/0QzFEzxOnN2N6rU9pq1G
WYZAC0qu1xQKesgV9H+N1cbMQFUvlVU9SCcXYpTPWyGjX1ZQvARUrSd+ar8TjcOj
lTbDpz7ADyzPlybyuWOIZni+64f78M3AjcBjGezKm175dvscV/QHzm0+srnBOT6x
6YgjLMDjvfO5n+xIdIGpN3T4ZLlSe9KXGAGyd0WIr0Mf34l8XyIbqO3L7/s0L5Qj
fJccRAIWDCVoh17BMymG75K+sLykjIgJ6YclDbe46CGl0gRX+DAj6ArU04MdWIad
mmp/0YP+yjrb8J2SWVxQPHhfWjAKf8q0tLuq1WTeZ7hexNHoL7O6x9dHOjxAIOW4
AgaDxPutH5WQwM0muIjqnSxlVm6/5GRRrcK4+BLvZpAX3mUhNrAtC0yqtKLlghE4
bCf1jI0Z4obOrjEpuE/W9Gl6wq9tHMwymY9+NvbmU1RM5cKOIlG1tJhY8R8sdfdL
45GZl/ViH8O/r/H+jQMKDuGu+b8SONHCZTptmamTVJq2MiOwmCyLRkVaZc0n2b1Y
ykaaPIsva2S7riy5cc2ZcTBRgUMXJDHvkLttux/wU9GAv5tRRjnfqR0lwM+1+nz4
eOEGMQeGH5+XjHFSGugNYhazIhMSqdMSMjR5kXXBjd599VJbPA2f5B4w5/p1sWEY
3pDlcM9N4oP4QCNUyfOHENChjRivpxyjUMeJbQUtHUPpHFwuC+8GXYK0mtyhd3uK
GjorZ0xN8RKWiQo2/T+WxCZD3J+yjIRJ7ZMzwidx0G58kdqhMJhu/asp3f9jPPkj
hvCf4aQeBASO7875QFWqYXDeskxSAb+OAI7CgtUD/GWgWO2hGxJEzLvkFWSCId4D
EiQb0zWMesFTJJFBU+5Jp27HLqXtAo4t1upSOo+VEXIneVYpqbIXVkThY0OOm21u
bLlJAjd9TOWBPG2htgScjPzScD6Z+4IJobVzRW7UxnZOeSS6IGwoWC9No2XOklWK
7DWEl4T/WGNnV+AYsBnZV5+kT+FwmtFkmzmZaroxC64Bq90DQmjxNl6IyzgYTSDJ
RCK+5yrZ7hGCTdOvwvIT5OP2S+XQ9ZY3fE2BQCRmuAxGHLFLKCLzNqdh0cmm9VG3
Nif/bMNl5CNQtY1Hr911JDe9yZDhIMNIG0vEWbTMpDusy51WTu5n+DNLeOEh6rq5
XaNXMLjeo+FMaEVAsbVhaia7cz3P5vxgAyFxAWoaJ7F+jHXFgmxd/BW9jGevj0/P
QHjz2kKXZJlAM92V1ZSDgTxR9MeT9+Sc23PFdvvfNHjOv7huEwmPX6BcqFDsCIJ2
ITzuW0odfobmtIGF+FF4CwuWAADV0DSaeRGi90bdV5Xjcqm6vnk/Odc+z8bnP+W9
WBgaxnApKSyQDOehiPGnN7zHqe9pBDT1x8O4lGTfAIDJyH11BA/lgXcshRQO1XSY
JdXOvzFcWVo41y7pmjIl28TbFRbl0erM+ppR6e9Nn5OK066waR+5YFvk8oSp0ZaX
+NclnrRqS8MpE5dyWQ7pdhpNm4jP/B4obnkpWBU3dYmhfjJTSaMfGBZGswo2u+M9
ENHs9xWdULmH42QM5peidfyiQdFtTAF5n9TQ8xRgsDM3fl9yyyT+V0Y+M8kM3e4q
EIW0eJHZPYW9pi7HvgFna2dHqEIpIP6uIRHTpbFsTu3mTkh08PKq+wLo9bwPyr7c
6W/OuivzhZm/E3MPV4wBI3CiEfqpS21/up/Xyyx53lb5G1GUr3j354oE7Cwg/6Q0
ay9D9EFYQgXXMOzQ+dsVfWMZhbdevjx8soOWgG3ZBZ/2mEsZ9pGFGbgCk0gt2SvE
Pod9VXrkhy6WzMumaeLY/pl1jco/ZpAchRGeSXbzgUeygW6TQkBbHZpWl2+ECOyO
WibtGa5K6bHuOcBUJ7EMXBYTXvhTljX/7WQDvotnkItKOGgHTXD8EdehTjwCTseO
1YTNpkNRYQZI+fC7B6+8aYiVSdXUxX7Ya3fWFGjeDh3zxGNVWoKbchYI84sp3k0o
TDtue+p/O8JU0tKMh786pz17G16wZK2xVtGJs6k0jJdLwyCHgHSKZHR8+QNJmXqB
ggnEJcrQj5WZgHp57WSJ4ydV7BCVzKqdQI9VJK2AT041XGZ2gqVEaDgT9TNtTwQo
C1L6m0Q4SXCXVT20HUKDFVbvJfpFXGkY0OD3gn7IbN4RvfIggIoaNn9LxEwtf4Uu
WDTETcKOd61kmoJM8UuvWRAQuEftU+f8rQWjSSAHzBgrLKWT3L3ai1mmgr3gBh50
yAPXVnTgD1DHYZsYnsArLCaJV9p865XYqx97QeJ86y3FZ7AKDh0tH2SjYaiDBDEs
yyjG1BAulzL0hAwcRFXT7nqlh/L/IDF0nKKSc3LOb4KNBKTlr7Tbeaqn6R6P9nFD
OnkmsGg/mZBgRg+NrgPbntK34/yfijU5t/+OG75HBE/FB8LR5OC/mjEGp9mdil26
B/zdZz9vfNV77YqFvVttezGGOFk3VIRfyTvihGs/M7TkzjSpBB4Kp9RNuBCZl+2R
MabPdDxAWhVi1wAZsL0q8EdRVLyYm57YpqadNHpEXG4J2N/VMmbOdStbjJ8mEYck
FP8xY7OSR510fxA/qqIvkN5sTwlOt2KmaN59RIbb8KsZFpk73mRBCiEB6rH6T8Co
Bzu986z41aNO3Juq9RHw1CeNrlcZllSw+n6TTpR90VjeOj+4ovuDuNpeMYz5Xsth
rJPGuwfHXDuUv3iYuq0SEatjduHFVJNdxJ+kW7EnQM4zyt/PPRTeFPBfQa59TNzh
nkJJjB673fG7TjCbVidQ9t79+oEKZtZgiBBd5HE4tXJ3dkNPls64XbMZeoSO4VJ9
ZZtE5TPsb/MyU6PtBT697IYFJubL0GKc/QNtDdHf/4b/npShrPwmpIr/exi19COa
msOiUBlO1dnPFsRb5mUKOBcUTYHy36hB7qafFM5H6e4T1TTo2d0dkSpTdxNY0oQR
E5ksE3wDHtI5FzXGoIFfqxwT7AutXc85WlU9hjEI3sMzX1TOFzITc43UV794BelG
wdm+daYViVUUGqsj/Fl6drwI/GC5+OlqBKlGNgmWEqewqQTKOzk6ZIsN5w0bOEm/
yIAMie+Y5M6pjXIocVY7dWY33lqDWO8+nzY6nGE37JmRoLMqy0DwZmDh+d1WsLyq
5s5sDCmQTAz2q95dmIolUDGIwZ0yDda0pADKC1101RzqC5dehWTYLYzE8pvH30lL
0p7hp+L2PYcqxOQa4bcve9ccl3CDVmqKReiwAqxIPmS2FWekelwmkSQuNRWCccfW
WleqWeuKZN6xXC0YomKtAeGn9fERGMx+lDcHgCqSYZy8IKcRgkUYGMCnoDe56GXq
OhKc3czWT/b614jITeei1sZCl0CkfmB5y7qwNHlFYTk5ha+d2kjMjm58/njWnHKH
B/6zU8rjRmct+WJ9P+Rw8SwGMQeSalznq/S30LWg3cFbNtJcg3XcQAU2O9VpezjY
CRfI2DXJEfTR3m7+opogAliwNrxv/yrRYpHvunFtMUWPaxi/NtI02UfMsHsybkJ0
6/F/mGLbBM/NWq2wEmCLs6s9ip0it2bh8k4rpFg3j6I81J3cvRi3KtKvrTtFXvmO
DWmlIC4ytsJEchWu3WcQ4mnBjpRXHa3gISEZpCvx4kjggAde5RSFgiSNupWMAUfM
sTJ6awv17PLu8O1HYiPqbgX93qHErxUWfrykhbbyS4vVzJlNrkGA2ckrMQtul/0E
eQjJVW7fjeZNL7M7wNhenWK91h/rP9jVryBPniYYW5P1uDKzC70d1TIbiNKQE7xF
G4xZYCf2i5U3BIHza/cHRN9MbIuly5Vk9at1epsKvoomYjalIbGcqB5ory8B6anC
Rf5U0k14ZQTNx5ApQJOVXK9g44ASaLXX0QMOHe6+Wg/3bypkjRYMkXMuRgRyGZaO
StX7jxNR9QkEH0a0E1BbjfOHdJiev3VXXoaQWfqzHydJ5Rv1dasXWs1bZG/WRZAT
EWRP6SBSK49FIG0CdyzIMTiD4upKE5fWlxQlzJIe7PUcEPnEb09UKR+p5QlIaR4i
ASRhL09Nz/ZRiI7tSZJb7x7UsRgKdM6FLVK5Chl1VdiKN/GTFsY7hzas5xNjIvnk
i3lNiMzZydiwhJR2VVphehUyolwVGNJxrqQQKyeypoiQoezftYF5opI8bs+WQkR6
+pT/g74pHkRO2Eg+lgsfTZQYSteUT8PyrtLQf3baexEQwBPD1xL8aH3rME/jsAmV
XZnc9dtHFVIqkOo2fAOfnB3qMDDDOY/Htz4Eqz1T/esev0MHOvf6oVLiFQbFp1fY
glM5/QUl7N/PyWsZmSZM8FUneIMHbQo009lOq81nCnpRDPJQyrJbgDgkJU+XvV5x
AVu+jHkW+lVqfsb4RT4WA/7pRHwE+mhxW0KIO8PlKOygPezg1V6MNAmEvcFA6UCV
CIGAAeoKGJ4FpJAp5CA+aJijaWIinMOi0fXWxtFMPDkANgGJakHcKPBSW/ymGsc7
z50kC12ldzEhyy3XT+BuQid/vMVfSr4jK+0jFeX/zQ7O5+jC2r/ajfaAEkoBRH+c
XtfjoCXlwaJRBRRJzV8qqwsL08+t2RxUaNOqCSfydX7sSPTxEy8xIFCDrVDkImH0
dSE70u7cIX6svh02caPOa4zPloea4XXN0ButdNtvV8DDyTqtXyeL5Cf9ZBU1YucC
slL8De1+IDQdofmR8WpofwfPioRY1ytkxf84XutjWTovVCbLFM8UrSzWRviqgttx
meox+TSEsU69109oNXvc6TzHLB6iWJd7iU3bfWxUH4iIbBbkPQM3OxtUnn7bjSVM
NtucMR3jDe6igqjnwvB+dY0K3bv0IfEh6RaospwPRuzS1K3rjNRC/kGA7j1syy/d
+fH9QbrABwiOGMRsA7XPlcwHkoDCtQGddfDNpCHC7Md6StGQaac7Yu7kHuHEMrkO
JzzCpxT/emVnwq7RcJ26TUX9OvrJKMVGtRGmDkN3s9Wk0Xlg57YeUoQO6SSEhgNt
4iHXg32J1BiRTnJbpHZafrTBlHZ1cBEFkGehrtqh0A0VzM/732yzB8ik1KjHbohw
KO/mtgSSuOZfLQYMZ0jj8aDdFy5AQgrO1LLXoRshcX/NkMYVaxElB9OLkzz/GrQL
IZM+e36OEpHhfNMSokd9sZ7lCdfb5TcqA5C0tSJoexqGCbWopcwXWT0PZsseIKMs
8Zs0jyYtoVBD9f6UiARooaPYdV3fWWmJQp5WT7KsUj664xwdUcPXW6LtbrciPEQj
OBa0yx8zYxvyWtz5xWXobs/E8q/x6WluAdeXIpBqTw/ESm7NjfjS+51IGkB4BNwB
FL2z29bGcY4YdIxwrFZBBP+VPd4bDSVI281AfrxAEZRU4A6Te6z0OI6c8lpHeIj/
gRion7z8H7bM2JI5d0Mxyn/yTqNnL2kgf8AHyzoAMfasPZvsK2hrdfrkRd68cQF9
9OEV2KN9d0HcmvhTwcNQ4gZkPGMv8vCnKnTBs0xt5pkq77o/G3czONA0R7KfXm2Q
GgvLth9pRl8OO0hjU+4SnySQPSKCIROAKZkMbLhhm34kxXingWTlxo5nQG2uKfKn
j35mlCo0+kediwzJb7UR/l5Nr/b7QkYahB2xmZNT5Ivxp4Or4hDnt7zdKC6ppsWc
N3ifMP/LyAI3/vU4v4aWHxDbW1SjK+9QKHwAOAwDJZ+FiVUi7Iuef+M2sVWWYsab
YpOLhtc9BjoHokmGLjD/jc0NvBXtjOeXiZbIyieON6zVfyjS+8ManeGlsEvcjLoM
yoQKFJk6+591A8Wih7oy4ZCKJ1C4nwQZAecP6Ol7xZqUh9IfqJ9+HH5//q5hk3PG
A3e0+jX5o1edfxbJPzCP4Nt/Urxm7lkVNGHKa0nQXcPKVw2V+ZrLT01MfbNdbdgO
52WUunbXTJytlHlR5RtsZQlk5uh5J7x0XTtO16UAdR2Nd3+fUAn1Hip7tn6lcXUY
H/TCEhKsSGAlzk3x54EVAaSHhQHDEIxfN+ofQD6TMYiHU/3CzybaiWFgv29lwyZP
eodYyYwbeeeDPWKfQXJoKWirwrjiDdOKZh2GJjAdLMzHlB5nK/mzddarulmDOojn
5pHG82Je/DV4xAxSHCqtEiHcsHmjdLs2s1oCqTklsWdn098f5N3PwWbvBQqV8aWy
NbCd2luFhx7n5317zWsfdE0z24lvUI21sy2ma7ype1Rs6OG29PBM3RudKN9a5oaA
f8BjPLEJ6S6b3uzvWmx8M7YheaKGaC19JO6w2zmAupW446h597q1doCZjt2TJSlJ
wM7zc8SojZFP4+Ie4JthnqmapVHkwcSjdgvoqrkePPo7TkfM9/3bk3gcucmUdrrO
HZMySi5BG6ia7TCvPfQkZbWRxz/ZHmTqyuIxdotyl5rmF0vt1+6RbjB4/FZ0hVTM
PiATSlLYN4iEWy6UskPCI9QkblK/GxlWuUPM6wTaMlV4kXTSB5UCspzSBSj2Si6j
eVB76aH5+tk2xKGGmP3tTjrfledsjgMEvzXeMxxpCKtz35nGHr4tVTPPZytumN9Y
xys+JV+R/bYTdE0WvTAXIToHLanRmGMoxD6Q2Qj136lErFuqO9BY6FaKVUcQGEVa
JnGKv8ukF6lEEIvTHYWyPFnja2rbjx3VZ7PUshxgnukz/VV046PVf5CtOXR1Vxrr
pdcvKoy8o2guvZ+9aMJDtnnSysLdo9a69nrCpvvnpNemyNhXD1IJ1+jR8iOXpnXB
xb+T2u5oPcigFHnVyODKIwKlKKiL+CRm+MOvxXnX3Wu0NftroAPD29O+fP3lKj4q
/2h7jzRkoQyRTfq53sCbOK8IflfQu89q2z/eCaLEbd4QAfICnES7e8bkbLLITYlV
4bRewM2o0jXGZn0LgJ+0jEdk3FfTyiLQGvEDbSWbDDW/8EkE1UE9JDfOMJCWRdB5
bydV12xm9YhdGmzZr/mOCDcXHMJuKfstWsfLZ/mzX0wLxpHgdYrgJs8bqCGOQTrm
3JevwrUJiDA8ccqUwErIquT36c7/P8KMa/wUb7KzkUzcJH1utc9AIWAF7w5nIWrv
xNg0JEryyOZfuUssB/lSOwDKaTg9wCgHDYMPgMHXQZlAxF6MFBbbFngUxAkfzXR4
a01U7t7a+GGD9otAVHwHR13nfMZrEN6zhfCF6vuteN11BqHpra38jehZWJx1wxDZ
p8NPhAP5Lg7c7nyj4Qk+5zKwtTzhn7ZOSIzpg240SPxLT3rdukdCLSbssmw0NI99
APOewNs5VMO6I92hYOLjhZNIrzeiMqkkf6Yy1O97uWp8w6x/P/h6FKYskViDAoKr
5YSkep9w0DBCDPZPA0zl8Rb1wLaAMzI/4VIIt6GX6RXMI2P2hlKlSf4lyIOpHvkZ
dPWfMtVD6EsB1/GG+rhKs1OVI0T9kBPE4g4Zxb01RAGursKXv4h3ECn2RD6UDZTt
waGRFli5aQeTjqL6tjax8BbuR4Ku1H2VtXKM2u0OzC14M418xr0ruxM98MgG9Meh
F2NbAQRYsJaV1JM0C5R/NlKi7s/TUvShZyg06gvtM/6UUjTM2Nme1TvKhh0g0ffr
zoLLfoKQE+Zi7G891/Uz6dzn7i9dpIQu1MjK0Zw54PjCPZ9lZxgxeGkn0D727kBp
H57vA7nalgctHcONjOD91S3vJMz97u3LIxuyw/SYxg5BskWxKOGDs5uQY1He+X05
ywMlev3nu6Py8r0MbsxCpUJ/w5Op+IQxWna7XMv3Qnw=

`pragma protect end_protected
