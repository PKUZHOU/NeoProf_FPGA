// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
rkfAzaC7ZVFTUam8Rs2Oz04BK1WnjYV8PqUHV1/dBnkjnduDLYBY6l1DWAkakgL9
tIRJc5+J3HQnHiEDsiXjs6ZDs9uVKmP2twHkoUbECK+kQ5XVlKcwLBoXUc5vLMuF
cRcdunIcTACsdytgIRs1NqAJfhi8eupir2E5ct50230=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 26032 )
`pragma protect data_block
cRLeXR/BKbWN/fBiovJugc79PQVd9dwJkgz0aRku/owPWm4b6S3tJ1CS8V5E7WS2
u2+WTSzx/wW5ShRa6Xwiu8xu8owtwixs0ACdFg4PYXE11nTJyfRsSbHVvaKpkiUr
pisb1/oFkaMrQfJ9I+dXYhZowZ7iU34rzFS6AA4Ca/t2ypbhSNkQNilz4uOLgVC5
Z+EGL6cpTJjJM3gIc1QYEIyBeLtuQZYhDYRnnajdUIuyJbwPpAccKZtTauno/VPG
r0+Gf/DAmTaOd6JHtu3ePE4uJRdszbZgx+1RxvI2dB5+euoW8go2L7Eu1+d+RQeI
smlkG11sgbS43V0H73dH/s4hKzSBUMyXZ+p8AaYJJb0dS8nmhxG3AECt+YjwlwfX
ASNlQAY2FhblZv9EfnX5qz5eXlO2KoqFzYpbl+1sc6sDsMqQSoJ/jvAx6Zh3RyiC
Tk//WlmJHnmoZoNixMeLPI2UK3awl078r70SudwHBq/MAvrx9mkqh3a/o7ozGrRi
jPOihQio6x5qgBH+Bu+2KvaX7TencmqGvAobyTIukTuNxtVq9b4dZE0DQI90/ssY
Y1aPzLOMOoGRlx42vhOEmiU2uos4nurgS3rDj5KVHXcW/OwPcpRp90jwHYyA2sg7
gsZxX1za6Joc4EnZWpgf9g3LWSnKvHiwfjBNWK3Fnzfu5YXKwwNchrbtsEQcrcvY
CEd/WLupmCfLrxLKDKvshk7IkgRUJQn3Cnx9Lr2cOywAEDC739IXVVX0cs7Uyn11
Ci2Iws2PWG9zHe7094hNnDBQb448yTzrYztqsPW1olgpUJA9u9PgFPkXa7FK+D2k
Y6hA5hWSplMOpzS421Tu31z38akEpNv7vZkFMwe2yZkprpkfRsjIhnLrE7LhA4bM
i/nOZIRSbB9bCZU6KPKq5sdrLL8jX16sOiZfX/xINjjgsQmCINprZ3RWeX9VmCDN
E9ny6SiNPrRlep+sDFo4EmntJni6JCla8QWZQ/qeOcR7kPR+paXr3nQbGnZFF81J
sOc0LohvgTNo8FH7j2B4IpSc9x/hBWQirvlwFRBPkNj7ONe/eas1yJMBKUSUZved
XKvd5/ZgXYcHnhb3ROcoAf7NHDcFnS/wOSeqyHYZ5M87JHhDsx5heyoWazb+S4ya
R98bO+3TcRFRKYhNaS2S5NOHyEr/MXtrX9MWZ6ziF5VkN9e7UP2caNvLNf9GBHLE
0u5JSgQGZZIGgOYnIqsV3YNYY2rXVNQEgs8Y/gPYdAlVSkQNzkHoDctXp71yGJYr
OkYnoZ4lqC/KhuAe0wEa1dZRwa7eHIufCJPk4k5cqEvLX3cVEtrmdsEqd7WjMzvF
DF16eFq9js1qSKrYI1NhvvDDWLTmDWT7/q/7wf+3873S1dRvs+pYLtogjsWdcdLJ
tuOSrmRB8b4jXydKNQGMoe+jTaT92tOtNzFqxdTSOrzLrLU0BO7EzMPlLgW0XyZ5
LVIEjF60jaVKaGfz3qpOY3FPXNGTAR2OKhPP5Q6cZBZ64kadhaTxCCFbvgzoOX8r
yM3YCcibhBc62uuZ5XVgkSNSCXmlW/HBI5ZXijLEIgwqCorFby9mFlPRSzHASkim
0fmufWshqLKram/C3aL5TIn0/He1WhE4bvBSYaYrr0Uxwkrdb4djwN8ZkI+vbqHp
1hGI2siZ+uY5LjZmfcE1HNGld6Kcx5llZVhJkWZhNokCXLSxZLi+1l2302KWCLtp
i7Zz7QY9QhzhT6zRHBanmUQsDF2XRJQfqYVy0oIofhucRWExC6888egTOvh5AiK3
WSqm+RDoFkhZlMqM/ZFC4DKw1hJdQqcQ8c8dSJaU49UHnztNO7WAJ7/kVzu9ocjR
QdHxc89f69lT9HAcQsDtJXPowBZEqK/RkcUIzS0nD3fo9sLawRv7uWE2GvSoyh+i
MSrxVZ+IW/M2IuJDF2pcXf4rSzS+zaVxmCChlzEVYjFh8IXEEAIQAcPiEZ+kR2/9
L+XGKbdw2tZrZfelOIeHVnSImUSJYI6erfK8UshSi5ji0y8QiRzDZG2WUHnok5ZP
zMapNlb40huWjMd8X3G+gAEgLB4ry3m661bK8KpYuC8RdFd12wF4ccV5w2dNZf2B
MQKCR9YjcG3eV8cwDKCfWxny0W6sXuYSndYRKti/vbiZ2ZlqFfqEsElHNf9jazxt
iV6mlijAHF/ZcOml3bqIH2BsFCObc63BBxxY4VQYMgAIxMBupXDJ/6E5KRe47deb
XLgHX7p9ngPggC9wxzQCbcLoH2awwdBb0+S5wOa4nHsmm/ZJLlBz3ars5Q2XAP2x
7DAZBac8BWknQ3v3XszBD9O9mpG0/+379xWDXkMdREBnnJYF9DhjKDzDpPRwprGa
szdLHE8HOULOpJQ+14sex15e0gE/Vk6MmKt2k+MSU7EOYw3db1shWBqTVnokwCTW
CQhNG7AoT0KX8AM/i4FNKotfS22IRI4wyJBgrtzXOzi44TcCfVvHZD0aIXEP9qtC
GxMjlKtqmb3LqTUPuXz3q0smOIltmYSZUkSCWw/TVlir0YfDtM6H/sTZv88JUSSM
IdB63kiWu/qShy1OHEJYXBy5ppJ7jNPIHlYUbdHLJR/ywNTQuHs/Z1a2DlYBGuXS
EEDVOggfVsHAzFFM25yW3B6EfPV56ddKlyykYQSpeyc1zzqlxlg5+7p4Ynvh6t9j
mtWN8Yx+WdZ+v1DtupcJf7Bo84Q588nLIwEVzhboPVRKkgLjcw4IIM/+fB06SsrF
1Xkv+tTC2RHAnSDZvDab60Wf/bhK/8Ha9kdB7VFfnXOaFe3mbQw7a0+FgxfkEcMF
+KSjJAaepQnTOR/02Yg+FWnc+CUyoBAwXjJ5F0PrHygFybS8IKYvxPpD6W69eoBc
VORi4S3+vuljMpLZXX7kp4RYfuvsrpMyP6RrwOK1CNghteNV6PV4RVTbrsqAu9o6
VI9fYJwkm3LsDGRITzV6SJ68/DVLQfrWge8wdfQbgUcPRmoqVGuZMvhhczL400gv
1kXwPPDe/gAQKCD7ZaOegXeS9NX92KIeEktleaoccxpRx1B+V5bUwkaThI5fOJ6Q
uqV26dm6cF565dyfaGgXtQxzVaIGwJWdnfoiSoMP4bzQF/zsnKOKFqyJBnYtZ4eG
/Lz5hDLS9G6NQMQzxZp9WTCK8EiH9yRzWH11DH8WlzQe60lySeqMvZM14tbHMhj6
x3IWoxHLXWRECiACJdY3J2bqZAFEsW42lAeT05/XXNBSQSLd18NAfk/UM/EJPX8O
7lhLHSPK3l8T+SHC4VlonsGNEchil0TejzZWMwHzrbxrbxXkeua8GG8XYTZ0rZYK
Vo8RxcP9K3V8vpT6elBtkIzNUm+YhsWOwLcLrOgo6l7T7HzooWhhHyyoUMUUwmml
Ellp0dUJ4IMsTA1saMWso4bTUYlzXrbPaVdbQHYQjHPNumyEBc177Oq6u5lfdm+n
njQ0X6Qu4xogcsTD5+AqtBx4YHY+qPFaO2MK5eFgAx17sgpzHAIu/m0/37w4C+Wr
asaHIyJqSQUKUI5obe5Zu4Hzinao8aY9p3JVhS5reJ5IATTzyyyWCdjPJwriUqrN
D42EI7BWkIjVT4nKIcb+D6h4u6iGPCGHY2UpXkvx2dkzWRD4Prl4Ohx5CZenGzQ1
AUhSfOzwP3SzDDdjc98pWeADvPIvJ2HtuvnT6Og3fM7HzRM009troU5uvobK9Ldu
nxpQcNgb4i1nEFXdjL5D7WJArKIUvM8yZDjMar2GtMbRqW8w2dU4vwHULC9Qbrjj
jWW8G7igX6e/dAI9sEy0YLs20rIqjQPlum8yPP5tsO4NC0zeFCRBxL5qaLlXCXil
jD2RO2PL1VpRMpEFeR4YSv1DEsHvpyKmO/piGyjhD19MqmyKJobfWlZC2fkUwsdG
S4ypTYKj+nR0llKiZ7aCET5FeAfSzcibQNEIO3LdVPumCOA6/JXeybNf9WIADwhv
02wx2rtTJniHgJKoFbk+RpAUZUvj2Gm0ZeBlqYkKTFFp/c2IDO4i27ZCEE5xBCUo
g1xQ/0Yr3UtM6aEf7QU5zywiBbX1hJebUZRNtg/Fm/BgdhdIG1z2EHrj8Sji9ZlT
+weGkwkF7CMejqgbqkH5ed7seIiU8FfjFyejxntNWrNXFX31pN7IZ+coU/AS4qfY
ObQxg1Wr+FYpdkYYFKXPWgNbAYVzaX9IVLhciANmw0v3YYHE8qst7Td7ZmG96Xo5
yA6MrQBZQ8f995chl5WWJUq7CH+boChmsxTfo9Rz5cdTopbJVKtDXRU7m+wN2QyL
2/dopx1ruYvDOa3D66Fisc4w2yceWGE1xnIpe1XCsE+JB+ULH7vbmNMthCgIfQmS
IwpjHPJ3wimNd9dfhc+QPwlvRR7dxmnE27Dz6Anra77n940W5tGf6cP99ulQ2KoP
dJPaZ6+Md8V9V+mSupEAv16+A3q37tAFwYa9SPusCtyOEU0NPpecqUDErRAqR6kh
31LsdVm8s5YFZZ35LpQ6ez+QQrUKwCtgL5Mz7HGyeCW1XmTfxprHh56gsZMuFxlp
n1CbybCqm8EZ8rTccrEgK1MxM2yFHHR27nxwopgcPZXuoO/MBNHoqsHEFGhANk/3
LqSUbVxZKoXsDOHQdpiT5goUgmzo/9poS9PkuyQKqJxE0tmLwu8o/Ql9QyHGN1J4
ozmEAODAj2ZzqCgIwWxwNB0E+CBxSEC+LjCCC7fDQfVP+tNW26eMfpXbNNMUfA/H
xSzuqy0sBuXXQtD5XQxKLdOycyOZjPerFr+LuenM+MhNJ4glz8meJwd5Kb3q8pTu
C1lPNv3kaXZ3YHN1VwzLMZEgpJRSRZ3/ZvuIKZ5gGDVCrK+7r/cJv9LYxOFtSguF
P8qQNcf7Hw4tJHOKPyTAc5W60YQwCsmRuvY3eTNEpWFOVLzcHPbDnJNpchHsZWXw
wczBJPptAJlTfaGfv1L3v2kT31yb/X/9hdrSCqm3GCAkYFK2zoUzfv/RK2efeTVY
P5wbwIUWgUy7BYXHPj0QHxbIdv5rnsieCyXk8W5RDapU3cM429v5/5+VhNOxDZYG
MnlG7zAWwhU3hG17RBt6nVZA4XGXROdJKzDD+0tiigXValbqEDBM17t2RO2bXtB1
iXaqTbuj6bNuOtkpfzfNbWZoHMXEEHLU93e0luNayORxniacCv63GmtYP0n5euWr
rN2cjn0P2iiChVtpw/ywLf57KoNtlWyTA6Oeyhf2GuI1pDawUFnftDNospr8z8kX
U/6D/8QSZUBP0stdkHVDzPMQFXNf4qPpNnVSoV5hUl/JI7XCN92yCxpYTN8wEcta
ASeAXS+5DuaV/rPMTCvZeVdpjebQmp/pgWcXcCAXUL7rNplx1zH8e9I7xopl4+pi
CKpJ4X9k2KrIwk+vrnOjoRuRGTFm8qB+5OEwxyPdenrzRv8RHIhyY2aY2GW+HIB5
eMfrIjQRi7AB1Vp6GRexZAkQt9f0per6UOvFHOF2yelqnu6yJAyTgn1JikWVNycY
TAL8bPrrmFkhYsZdlz4ZDl1H+6epMC7ICdLIOlY0AJQtRhmH19/0qSAIpIMgE23p
YTI1V2uWsHlYceAurCfoUrV477p42RQ67YMMDZPJliskwwQNg1z4bFryqR/Vhd9z
BgLHtDYSOMtP0OIqS7Yj+my2OMcaszhj2HxsUsoB9qIcTTDkMaY1sHwRbHgZwTr5
FTvgSTLNyMAh7I2SErw76h8wlkUMEEMi6mr1CKjW86n+YUowlqJ2VEZNlxJrwoFv
mpcEmntlVn1beF+qeIHU1gCvH6QGfmLVZzoLfQV06pGuDQ8TDYuCx5rolGOWem0Q
ddGqDDIPr3Oyl+mFWjEl8D9b8D/OhrPQTIYm/DJ5FRbSmrq9cBusbexWHQxMfyaV
Mjb/A6AB4GPq0lPeHZX6Bccvnk46c3SmoJhoLSx4faq4psnD0e2EypEtB8OwIABX
LJrZqUD3nbRogCtWobdA2hgnMbLXx0b9mSNtz+2XpWRnbV2afHmldF5M80bdCOpn
aUsNAPdMDZ13zZpSvD1EQI0/wn8Tbp2bE+Tju/HVeYtsXHf/AYbpdrJODLxpqmDn
PcebEIECqlUGxmxRwdH/WkLshbQJOFSREWr+KXufaU1dMQpxE0+aXNYZcCQdkWjj
aYuTjGohJ00cnaWXGt0dw9ULCEKEk931dyhRvetWOySGrzyF7iqmqUNaQwLPZmNK
rPub6NAyFcSH6H4JpPXyZsJrk9iEbVFy52daeY1O7IY5ucU23mOdn7ynsBVI9Evd
X600DUjsvr4GPY2s0rL/HtDJ+nn9zBOCm8o56USXvs3EQX6O83nSTotQK4rU+jfL
IkQy/KLCRT987OF5aOFHmeaOeLaJW8kBvWE0QUEwxVC1RYRWPAuJf0rrXKGWRQkL
Zb4rtq2mMant00pmFxVMfnmdATD8aI8p6FQHqBgS9U7+/n5HAUExXG2kIRxPJhEw
rHyUEk029g2RP46+f7cL5QB9i23GMsidFeweG81VfngRwqi6yh38RPiaiEqQ8YCZ
mvt5SgErzuuDUu8VxhR1cO8wKcv5nOzv9NobrXT7PzPg5ti/sGfNJOHQ6OtwoeoB
0aYiP6HGEWx3viXhnnMQLC2NM1Mrcz138RXRYazmrt/Qh50rKIfXlpsLFG8RXyg3
o6Jsdbpd6IdsoK4D+KrvFnNN/soblM1hU9r2YF8vHxes1tLvft+mSo640jRedDTR
4YAURJ1ej/tengAbFJ3lJCIIyjYBCj0uJoOKSb1h2YaLGcUrt28/rQl73IpmyaMX
6CTwWq3rqtMVV27BXoyUWzbMNVhsAyz2CQFhZYC33uJkbbdAp25EvQZQ0O2uBJk5
O5wbQwm8W34KS4wY391AtN1eGWqp0d/beNpD9nWYytyum3phkIZkfZIeeFUOMd68
lAf3lV67Kxeh7parK+oJ8aR9/pPYVKzUhPw4FrxHlukOs9W9dYkgQxu0L+pws7Hp
pn6CGeS7NTmrwAEClw99R57MRftFw3lLUB05w8PjwvyRcJBL2S6Y0/pmcEvwcpJa
L0Dhf87Q+tWWXYHBTb/4K6VEMQWHPvaElHj4C/8J8IbH7WIEtVcXEJKYjfshrRU5
IHXutt7pLS6GQLXMCdZxkDqH3Q3eY/jTLMV9m8Xqnt0sylDdKLN/2lMc61tQigPO
NGGiSzoj8/j1Gu0kSOErjRoEszHkjPWCfXl6WLS/DsFETB8P9HmptCicNrNhCfyT
ce4NG3/rQFryHlE0zphEWfOBYqVw6Oa6eRhXgCzFUyLtRNzZFnV5bEDnY+svENHz
pIOvi0X+ejkyY25sDmccrcOq9ezPOTSG1skfOXpdsmm/jCTUAkBmzlSSe0Tzgw/K
GA4nqvCwRYTdXb/2xln+CdrNJXmDDiUjjC6A5yFrMVW224KvZggmnZ1o6lcHCphW
DOGsN0N+TIDFcenLgwCKhbFBocR0AFjLIeH7ag/kAZTvuuWb3xwIwSx/rVQK8VIQ
H7dIW6kg3DESlFM0MwGUE+oBtEbieutwRRwiZcGQ6wBjqrNPJ0wHr34bQTtBCva3
cyKfuOn2/LQ/SN/8X6iCrDEm0yVh0qFwdnsa8rNSKkilepDigr7XiPp2wf9edwRP
TFOnbRKwcTiqW/4/kvSFIm/9ioOY+CcZeP8wrImry0HaN2jg+RTfZ0y4hJG4xS1t
SwyjXgZ6TiyTfyw9tNDo7j33uYA/oHcPN4h6TweZRn0XBCxtlcdR0DGg8yYEEupA
O+VTCxaLAm7yrLFhFmlOido0iWx6aryQr0BrCEw6af4xMQ/rbVplF1ULIcsbuuV5
Uf93I4cz2H3tjmRfNZdfdFnnpsH7+qmWDo/2tRYmk9Q7RzN3r5g5zbAl4yiH6omm
wezXdrw7gMckVUidi+4THMygUPS/7wPi25vFpckwuVflN9TPmjGLPkFOMQ6rLAZ4
ATqmuI1++ytQH4SOFeWT2aXdtIJL4m0N6et87KFF+i1GVNg0hPSj2FTY58YfeIpM
pHrp/tScaNTSCp/ZJ6cFXNE7JwG5WNIz/CJsNA8Yx1dXZvwq5+V2DzO8PKR1hPhv
td+TfprKSKhrkZt6h8ZfeLgcsYoNG9ENq2NCI+87/417CJU9gdUinNJdHBeLRDsU
zQhineOnKjJSGjrv4dEPzo6XzBbxAIq0ML17hW7EXXXpvDuTScIRofHe5wuV7/7e
HHjwpjEf99ebRAErdN1Fwe7mQK4hZmO1k1+YBXYQ9ZHGLbyjgfyY4Y8haVBDre0K
xOwG1UmZ/AKuhA0IdV9jSY8oERZHF9EvOA+DV3jHP5JoYE2JYI4wiS1OB0kDFKr+
H4Z7g1eNEddV6fVDyAG3ukpWUS7C4O+2tDO1wifukrBc3rP1r0g3NyxlmLJK6O08
S2Xgi96RM78ILGCkuoaoDqwob0vpzgGPrn6zG1YvqMD1LfmqQdW8nrT4tWzugpM1
Hhk/GbnAoXd91SsPyMJgYxWd3GM3zZy8YbKpC+nhTitMjxr6VJZNbNh9eFs7nqn0
6/VSLoxBkg2ZsaLAQzSIxornFw3Pcm5m3i+7PzYIA3iWBSORtsY4/Ug1m9M9jBuj
VX89051GPyPJiPAK1c3tdejvZWTnPh+X6qntea90nwmuXC2AOw4AU/aOiKChtYE5
SZTw704TEnxbPrV/cGCLP+q2J5LI8o/BdEFGpe4xeFWGVydnR2k4y5cyj+VIQwtv
KLT+PQnrV0Xf9v/6yFwV4Ttd+cL5VHzX5uNB+dOeol922YU6cUDX3zhqfCykEoM+
amTQfqsnCsbkz/UAcuCSVtjAs5C4Z3EItlathCU2PqRPJ1dPbKw71L3YOBMQ9pdz
ITA0Ybh/w68ynn8tMuq6lgOxRc16N0TyQHGIHCvLiwDoy2q4Vqsmpr7iGtFGaYvV
qx0+MXFim4fIFHdKo2lpqBwDyiCEsjlDJ/6SbB3SHE2aOZhKt2U3huDP7TFJoZMm
ge+MGxF8YqABGDfrfBCPinSH7xvbMwv0j8X6CwkPyc8UXqo/+u+hFGk1AroAJ07v
H/HR9f1z9LTfnPvRHB8vlksEKid50ys2wxCAwSDQSiuS4mHHdvbCwKmWK5hmpu/P
PjlIuUYkoqEPLkN2awSLZSDLF2QytSYlmbEJtSJfT+PixD95UZo+faorxhyZlMd0
BWhA/2aGG855VIKe66fzqpj9zD1WvL2kMJzMtw9vwwbY+3tBUwgN1kidCylA47xK
pjucoi2T7cvJ6AxPg+10gvS63dOXDsdSvnrBsEfEBLOXFtyTbpHdtxTy6sFofdee
2X+iTxTaID/X14egJz9JtkYV2MtBtZysdsK0wSWLINK8SUov38uP7MDHfzSzSyo2
vqQVSf89QcjwmIf9HOrlRX2IldfxxQm4KPlGQfbhHhsqiTKhJnEGXdKNl5OeFJsV
zWvKsT3yPQeYkeaKCPP7KF2l9HuSlihbgO8pD5hvZuRIAGFDdDB3NMN7Y3MzmWgF
MNJXSW87HyBFJTHPwnCled3WbFL2qe8CbNTyQZ9TPLeD4MYOZYuEk3PRBnWwYuiW
lJwXG2YVY+l2Kya8iGKJ2I/VpTJN5JWM1qZcIT6SI+LE/FMVZuMhswyRQ9pspni9
m+9gwCMbuLfMZZM8PDF8JqfUTO6+1WQLtF0ZLGxOWkPjuGKqewPof2/VI98t5d1O
U4RE4o4PzJ0q5oTFm+u8Fln+mPIKtCsMqEYMSb394I7Obtc5D4/5HffnuzyReI7B
p6V7GYczt+SB+OiX27ETZJ3JKb00wXirGlpa0g9QgwSV34cKGecqLFFlXLR2XbfW
d11C83/A92aZFWp2kzG7EnHhXjTqZjZ4Ff6Vd5hy3acKB1RJI3gxYrMntepLVWq9
YgOspUxd5XjJlMtMaDPnlck7ODckouZSXFoA8ER77uwsxSiFdyHp1IsFggHGjYHw
ncnpYmQfDbUuNuMnOTuORgO98acH8ITMdSj8pgOkW6sIsplMEMeXrk6Pc+rhz8lL
nONq4IezzGThHfORpKmqwE8keFTRM3fRxLZ66MXZd34SbOg4+hcAFckXQ6Ox43sw
pjKCqj3kBLlEcJqfQAieKqhQENx9IDTItiY3gS5WD+qy2OIgnbQM4+Es0487uoKE
kdAVjoATl6T1qr4Ftajq42kR/WNN2R5RQCh0lBkSti9NEv6wQ7MKJ1nhLDv4nGTC
LaY8/rfUDKJO6HO2oQMDH85Ud5OfInOFjE6bSiEvBMKb3nM4YJwLz5MRiQ7Bsfzx
Zkoh0l4I+xEa4so2xXn6lDi74Q517JM28bpdd0KOHkeO+nwPBbKCCoxyMUJ4Fqqx
+aE2F7EO5FSEWN1u8jCm9y023Q9xznHSg4x9WNqsK/reHCIzoYw50l2sJxZZr1hy
o5WEogStDGKf5LF2albKY+JLkIWHyImpd5oLUidZNJIncb1lesb//jBvbi+OoW2Q
EOpMWstxYz60aW09bzwG7EiqtZxZAKrDZJ9zFCB3QkLQJz7GUhiywmw0zZUNWgwa
OLgPo9rGYO4rYpPKfYO9GJwFjnFtCl6PvFjbVd+o/pYs3EUyT01DSPbEylU24MpG
O4IYiN3iVYedLDSEtYRACbvbSkh6MwUXsCz0hLsWKMY45602lWs7683vYWNCRaZG
fPrrbBD+xb3jyMP5cop4Bmz3+FxBwnwAbM6s1GoSZNIs+llK/7bL+SZ3bc7F8CBu
tT7qiW6z5IYC8NT3od2wjWrPTMEdcVhis3i8+dfpoMY0bIdyy/8R66zLGHXHAXgg
rPC/vluvd+fiE1iYjtVj+k5YlysO5YCqpNWAuWLoNrz109gChGdCRW/20K7DiDkz
s8hngVqcfkpyhUVZ6GGvis49pbQMLHq7zXlGuyGIg09mjTz/jiNsKu8q+wK5x3aE
zS9o+VUSOZu+e4BVkAjjODMqrLIlG6iO0ZpXDpzFfiZ2H7UOZKLorwz0bjQsKCga
IqoWsut44tCzqUDLtOm85YmExixmw3g9Bm57iPr7IjphgOIm0XZDEu0b+xkhw/5g
jaUEIIHKC2wMk+wNnyuUq15h+h0o4Hmd5lqd46CHXUykUgTu+Ju0NDQjvbEZK188
gJVC/j3clMECb9aqU9N0DjM3fL4xypxRjfc6AxE9hmQVuJDCUo3XrlOXRLfEeIqu
/eNNqxkibpznKraK+5QMcdiT3H2G58zk9HrrgkBajzjYVBb6XGwYcjdeRlGTkiOB
KA7ihkOgaenH4Z47jeDuDLgjGM5EpU+RygXK+VzKxlkvFI0UuO+lHU6hKlwPqpYC
HG+T/2CQIyfvRXpN68agiXBV64sn9gpyJLmHY4ZxcgdV13Pj6q2ou/O84ZeeY0bg
UCCToOkvlFoUYgGL/LJ/IdOgOAvH8h+e40LdYdS0NnUiRcA2vDUcfIYtJAaaDJLn
83nQCgVwM6G/kXSpLqa39IoU6U0/r6HWz4TkhW4MkRhPSXlm5Y+Sam/PNUEvI95t
5/yh51W5caiBwyYbYy95d9gUMQNdJfwsFGYkh5zaqPQ9t+SbKrkAOYCRVnXZ84f7
vHOrOTZJpz25gwq2gF4BrI5wHE1JnIfGf0cGgRQHGLVeTlHnlKoLQoAp4hopYKOt
LlJrEnA+nILYmC/UUunOi9T8ePOD8mn25Ep1yjhROldpxy02592oO45sytp6ut74
pUh64A9+yNeEVjbcuuvmMm9It+bomviLK1BT47bDiLRzXUNaXBq7xu8ZZklPxhNh
ucdQxmV4h9gvqfByVKW4+rqQAsqbU//qhrndj5vcWDmm0ms+7zIsvScBWgvJD/kk
ZfpwIXlkuYxzLiUREPy3Y8cQO4y/uqsd0m2ZM/bCCi9FXuY4CvrO/PIuAJfOwRM+
mUE2HF8x36wzufmQ+Df2eQCqxyH/+akH+25vrkArrRFhFrpI7CEzYi0XPhiBFnHj
P84TV8cu66Q16sQKAnxFpTqZGiC4I0InBvzRUNnj8ozvjkUSEsLrV71o99MMYmMb
1NmfFsmhNfZ2paskmQ0a40WLJrVW+tzbn0UHnYC82gfL7AXljCLZN+skx3axUCMc
WrC8IKtPm0GsCPXR/9zzev7ML3STa+c2v8jnEpz2yWDEbHQ2rk6cnL934Uil7Iu5
ATdDPTcs8/yrwP331OuW0b0muoJrWs6TIJaDGNtVungvgRDuH+7YGDMCeI0/wMId
fMI4BuVrjylaW6Ki543ePe3U+gUQJaiir75c5CeWmF8/l8yFJReBaNax6A1v7atO
Mu4NYoDXQV6XqZZs4jbtkn2kGZ4lrSVnfOUuxR8KKWPtjQzWcrUCXuq4NoSL9c8q
7fFS+BZgRhgEPHgAJmWM+R74aePKOPNNfaG8HvRSy5m1i89Qc1g7vYUjSAaWzEbX
boqrshi3DzQ4TRdcRJy/CKOFk41J5FVFdUWEc9f7x8myxE3/rHJt1x7gt4No5Rri
cN5PV2/R7UuFza1gnKN7NY40pWCfIk6AOzyWw+gBtKqCSy43BohZHgWERWEb7wP9
oHy/ZpJW90ZQ6NDlyaQQkkXkLbk277n9SmTswpOgcRaOeXAHECK5WoJYU6SzcgIg
PBTZu0n+AdFw9PjGRB3E157nRfskYPjov1p6wr0jH0pJ0CpV1Bz8qGe7jFVQre/c
bXe/GDqyNLYvoYjqDIj3qKw/jQ31C/lMjfBJUID46Mvlwel+Fj1bDAR5X+2LpfuL
JMhFLEixGjWgfiT1akPGpg83k3kAIxDGXAN+wug0KydGeHHJgr/SD0Q6S43Nyl4Z
1pU6risL8iZmOccDPOprInNLC2zTZ8DfJ6BlY+CdZa/QHkwmHe3sOP0zA9YyFANB
p07M+y7CFXG3ddWLjFLLh3YtHsmR2Vv5Tx5iwz/cFLESNPliSeFSZb0I/mDZzxxG
BMf5SiKW8ebGNgcXJIRELWN5NDRZAA/yo3DmIRGRmqz2ukaoHStwEwvy7zTMCf7k
oEVMq1MMUrxxSdpiuFgCK3/vCBX+sOR+51P4gz0UrelAY0awxUolyhty9fRHebYs
Yv9CjL75VQuNWO0ieMXUQwVoJW9IL02rTsMub1yVHZq+t+pU7HmtvsSZQ4D5D6nW
4yLOUrYkqqMU5nfoOHigYZ2RghC5tlnHQISfF+CLsKYuYISK/7m9vIMvpzDu5O7R
WSCLqmWbrP/+s9H9KQPSmEEf3OjitMtkCQ2UQMkAsUj/MEs1Y1Zf01g3LxUJmHdv
elW3gPpsz/xTMWBVasv0cAdh+gjU+mquww0tlzpoQATJLVPVIisBS4cGk6YP5lho
Ve6kdimQm58/mpVDv8erDHKCJRsfKwUIRoNefltPx/8ioK/8Nm1pAZla66kLxPSg
RNZ59Uu84Y0PvshmRUmM7SkPMYhbyy8Up8GVwWbIK9ZsX6a9LFI7ymQs1UTxscCN
8F90TL0namyZGFqcANFhp6gtLmsdsBBLJCPcAxfSCDYtUZC0k2+IKC3W2le0OrnW
D7s58jdA/fbkN6YyANhioDF1j135Qoonxf+1JC10twxV30k+vaDfRPCEEkzQjs40
lECQ2QIZeVxKk5DWmoUnAmu8IJ3H8EkyfLU/RcHtjYOaSBr9DYWHupW3o5BRUBG2
+GPhl1VJHSMgT39PXBeFNT+SsFU8bcLGuCmGZ6Rr6UZXLc5nMMULFWYv4i8bpCXg
OYOzNxwYjVwWyOabD/hT4uUyF5LwWWDp+Cm9HS4aeQN0AruNfWzueSPEuxSPJ4/o
0e9EOCgx5qKN5T+6+0KVDyUQ4Fe1ushuKtzIpHwRGT26Mxv4urdDaldPl36YbaCk
AcRoFEai1nCEJ5dzz/eQMw9fTehTWpM61V2T9UP48tCiZz3r5SSyHEH0UyjnMIDs
dNgZWKhiiZBz6bb1X6eSMbuWnWmoHfHR5ohI49fUoYllq1Hd/sE7gJHq4o2agtSc
0ZhOq02Zq2WZhyz4vZWfg/fupFd+XbwrK7h9MczSWpofjNaGNcq4NzGy5OZIZ6c8
bwcmLJX9BJwt7SLydWuMSyyLUWlXLU7lvIxRhQxiJWhdZmXvjWrJ5CH+yakz6U89
EiMR59JrEo2myGgxSexX9MnjYDpqAek/VtzS3mADFTGjqsWDXVVD6uKQX+C/TSb+
WUg2WW0c7hKO6E4eavl1tezOlf23vOoG6F6zDlUHL4JuhFob8CyB/VcMIYJvOkEH
KsBudI/6e4fuRQgmnxxBHnwGHL5RiZQe10o3fTrU1/S7B3joVjo9grXgzSNsDs7X
g0VjIdrZgwfxCtXhHwAZnBtA97YtAwZCvNXP87Zqf/sOdbLXtdQk56MkmqP/YPyq
9kMllr1He5aJdcnvjELnzyQKz6f+7EDYhmPWuwMatJEYguquwt1wd7D0jHPF8rLs
pAUGMdE9JzZYmAGFT1yPlMXHnRBz0ju1rbEYmBxi2PBNEPoxdyCXBTnQ8B3bBgNH
mO8BguNvkOf6pOyz7/k/h/EmwMJHjJ8GQGdoJTpKmyBYE+nNw0aQO8/uxbKaz8fv
v4eWgbpN1QWo89Bxq0UgvSBCRCb132HD/zjvXdk9PfsFC0tJLxkEk5fNQ4RlPHdZ
zp1mMl0tRf9+bLeZkErXLwr7m8/SkC/ZreKzGkXh30Q5vtGBvyOXnXy8WcmCJxTt
QRZxg99gx4wqSCumbYT3jiP7Hqlzuz0OrO/5n6rTp7rn9wflb43583jSU03k4LpK
Ileo5Zb/w8n+mXVG8XeOWOzqgJcHRfQFm7Fov+pBCG8G9hd1O7fLV83hgYhb2NKN
JisYpURW2++mIFVkPSaiaAgZHAXrgjZloXvTcDLQQVYZUzABLqKQdaVr3YUQTnp6
kgqViU0HVToO02POoI4UGDW/GcrhQjHGa4o3MX4mojqZUm2l9SZ8lEc7w8QK1XeQ
m6F978Vmu/ui91tha+55YwQfsFfzGn4ICmlE4gG2aTX0ssXVh3CNWWY4iCrzfV4b
V/wutowh4/P9L2nIE4Ruqmb2siLCYK01NCYFF3Vvk6IwgwA6biCQLGuqU41eYSf/
Ac9UceZxleLiiIMNM7hPvhq9jEMT1GXf3WQB8aYulKX1CCaD4czrnJ2Qletd1Tfy
GZt6hOrkqK95HLYxWX0wNoectvY9iIERM2YETcrQ/8FSrcGcCK8AhsRgMiYFfLzp
GqxH0nZnKBpJ27cNk9f0JZ9vfWp4oMdQEKnvPMGE8N1+M4P9Fv8IHscNgFFmH2Rm
q9JMhrN3UHKFVa6pTcHGBRd7PHW0W6CNc42YWFcrhOJNDGKHhtIfluZMUTEvapbA
S9ZEsZjKxajAgmKWtC6gCoKDx2Ks3fT/tk5YbN9NEltRfx0tdVRGJzdSJzK288/Q
FKk3T3+bjIkgKLLq1yH6l84P3oaUb46HNlbKNfJHJZhUDH1yLeNgtX3lpKvEmkqS
r3ix8iXEb2iHd7QEeCFuoL5lFmoGqhlmS9dH6tYrqGgHUxU/hFfih5gOdn5mu5If
VMmXuzcKBvi3rjRBfVRIyG0LQP4z9Z6gCQA5T/F8wrkv5uIKDNbGKD6if2dZPd4m
DCoCns3nGoeIqIHrksuvEf00ujz8ml/xqnuvx6GSP5USmd4h6nctr04gaWiIwVEa
tu7NoBbDmOa/y1fG/elIr5crjX1GjeYmrRcbuTdBn9ykiBvVVsy8I0ak36iQejSl
idlTNIfXwdaFwv5FYbCfZLssdy/r8a6XysIbRjjSGcXbsAJtTPUnHW3c+BuZDLg5
gEud588/8vy+a5Di/QrA8OJ1807WwYwuXwNLgh3ghE1ZJTHRlftRoTIvz309FTls
a6regBSeTdYEvB76A7vz4yZkM7nyx45obydWKRPUTPaGiSCMfB/Hm58eOngB7ibW
/pgm7ulxwA6BSmzr70R6TPCIKOEe15ChYeJEVpYOnhPVPHIsVa0c9KqXMoMq3AnS
7ZeBQgabrc7Ilu5MU6ErfdsdoeIKFFervA6hCrpACh5zHuoriebIrOLxoZE2QvGb
WtGAcI1niHhlh2xbHUYSH3J2Du+d5XkH4H70JTOLD+ruOkyVP0qQCsjniQ1A7aJR
+++ZW2v6Q1wf/XYrpaF7WDONfEogUsnskHsQq6KsCm0x1k4rQx7q26A8S0tbZqGm
Bk3iPNMQzGJMXlw0PI2oMdAdxBjiwxid4HM5UbNoKxJow0XBt2/2VUHc/t5cpEMG
gbIIs9wUG3es+BlcPpd1eEXliF2XBgyz6JeYtRT4d7LwhBSU5aWdMTFAyY9PDZkj
pV+IBen90dQIRClSVVSVHrwbDqimhrV8aKfaMHYKd2TFKDKI/iZkcCh0FUEV6HYO
VU4MengCkw2s2dMeiap/RFdnt0E4QrDDQsW/1ZA8cNeC3WfTTTgjQ0/Eq9Bef1+T
c/VLMTm1McUdNxagnYVEiB3YmEaHrDUNLh5WcHv6lnQ56Wd9460/nVMNrTBZ6e9z
Gm+1LWrmCShSkSH/Hy/Y9gVN4FN7OdTKWX5+e9l+kq/mKABcVa/RHADSL0np2jw2
Mht4/4QKIxZAZ3mc6mmTWKZAUMjNNuc5xQ9JnLK4tEd67bXD0T5sZh8ysF14AKe+
AmPjRCBmu2X8GYkOW+J9XfXDqkRlRh1tV6ki2mNw9q1mrYHIKvx/3M1w1XnwSByc
oFq34CtS4B5SzNEYIZMQmmsd+/BFTcdvviPP4EXtlVbIeNYdgSLzac4Vfggu86N8
avMDw9r8aKgNFYWxwHjLLDXjXjSxislYRl4+xICL/EngegYKR7enou/eYU/R9zes
cJuF/SyvmfGJmmNieUWxdib68O6vWwjMIzAD1KRPkpin7bhl7Hu47mZBLqRC8eSH
+HBTG15kVCJgpNWp1sJy70uwrmV2jQh6+SA7sMIceBSzUMva71WsGXlYdc/sG2Xy
I88kw7R85TUTq7m2yPwigPBuVZRg/nNQX/UuHYQWWqbNa96MU+DhzKvBY/ZuhkU/
7XJJTLoQjmugt0SN5XfiOXY1RQNkOdbrHLTZTRipyNkthgNJP9R7hvMSLU0a/gOv
bpa84Sycr6X64Kc+nhO56VWWY17jLwT+hNugTMPOrtVvhq3G52FFPALqMiyGsfic
7cndcUE4V8vIsd623SB9RPMu5gJFIXLHQKNRdTmOnT62gH95fKfBne1aBg+24KW8
cbnViQbSTtOK0k4N0R41KYcVYzAiLVd+KcLZ83I+xqqE5JNi+I8KD0p7wwsaVkzV
uMN7JHJ8hYAi0AdXb4mx7KN6DNogQN+73AU/FqLyr+JzBGSvJVG6iud1kN+rzKy2
fGY+HRnxOpj6nSmySxg/L0akyGgbimXsxslnV1Drr3F8sjKTLhord7g0PZeynvht
le76eiCsmklCTU21V9zRXEQenF3L9FRAIn0DmqHyOtM2TH76p3ZhR30IDUhfXufe
SM8SslNuOD8QvNDTLgAzieWa/TwoEQYqcV3/Z4vVPQTUjZmnAhPb4IDxMlgRYOx2
/O1zJDm4M6BoXNFHykcZnAkI4ObF3FandTGlRPZy+esGtK+qhhg6eOBLYXMc+8Fy
YoORr0Ri1G6XxdJfCsh1uwa8jfMSx7K3YOEpiEpGN3Nwu7IfTYA65YgJYGYb/tsn
HkZ9oxTRybqPLClOey9DpCfYGHFK4Z3Rq2i1xQSkkS87v3Wrrj1JnZ8tmbKRMH8P
QXefwfaEnN6JJetrIA2tq8aWh7yszuyRf6tNZ5eqj0XXRGx1HTid01qAisGXUdiE
7cpysg3tdW0N/w0QG1zdokeCOoO1LYvFV4Z/50pcbMbKD2pPWlcZFk0MrBUB9EnV
/RXMdWlpa8KnksWEfhCoFAgOg30RufDjuYjsEyTx4zLhfHwcb9KQcoLEzUznIAUJ
7nL+gn1XFjADewl76QS67d6CCeGvX9AhfDmX3+pUihcXKcyZ+/r4nP2qM1gEte/u
UPSfibbwaUBEhsnGsOiKdJj3xPqd45IgMcthOEqqQbmTGcEPkUY5qDVMXTQCYaDi
rwijEQV+rUYFYTzrFV3x5y93GKF90lcenYUgTcCF96uMtogmHKOz3pLgTTUuwQuL
Irxedce1f90qx2Lyqi9ix7MFK6vytY6xsPkOFtPrzLrmtaD9RVM8oXoQfwjnrIx1
3NZVxsTPtdi0rWxkqb6/fgR+NIlqYKO2q4SK5PWHxgy6KdOnMe4pfvgOgcZOnhvT
W+lEzBRAnhlnRRXLRBPyA2K4V65j/gkK5WZZJ82GJni7ImGot7Dpl6vQSo1f968d
tIorw4TYSflY+MA/JihKWjqQBlzF1A0LljIqylW4dpwuV3pXXqsnDjn4uSg4MNb1
LosBRgLzw1JHt65yECUWS5MX2Ai8Gqbi4k/LBPIYb5uaY2y/1RkpbuIKpqwe0/F5
TzTBa2YIbEsM6av2UAjgws2dQntLwDRgAUVO7DRA9391oOUwp3cs69U1i+KvnA8v
B98j3saUxGEHjCu7/N3s3nEtQx8/fMp6bC2MzX/Rcpr8D1JTT37wQThwSieDrB2Q
/UBLBAFFgrXqRKKP6MSqY6htG24Bkk5iuIemsS/BXYKe9pxuoebU/mKZP1een7BH
PPBn5dOdTWThjB19Chpw/4CkuBIGEbY1tCnj5HGapD5CzdD+iubJdMaovHC2KSak
O6ftpF5V5gaSUmTymuqsKdeEwAiNaGSvfCUqKs5f6qISPpF31IqOEYjjCCxsVy4l
iwG6BIKKypjBGJGmZ7Z29fBJvhWzSN7/Hzs+jkiCYsE8wkkFLF+lX/BhHJ4fvITd
DjkvGQUbJrcarF/PGKYTt+4avWerBRJD9kiixEGNL3Ov26sEbm/Cx2zt6XvZtdyv
yOyCEIVdovrsXU6kBCvH7Ls/ngo4a3DP9mxv2aCCJVZPlvRrlllKjJV2TojCSu6U
6HExqWexoW+eUmc8LYq7JPjgDSIo+7imz7HWEH+DHhT55LPnH691n/IzgTAFheAz
14Agr1FFITv2jyPrulJlW4Ajx/CgLuKiij+PvogllzVaJvCT4t3nEJHvRQKqQQdN
GtZ1ApdSsH2DQWYYQF8UmR6QdkdG6Y/+73FB2vH9u07HQVGJpi95x53b0DlnTWMA
FqqWYYTRQmhD2CscCbpCY4PRdCqOtCRbp1kK5QWOyhJgnaxSh+jyLhTbE/+5WOs3
Q7qwbTvvi4VN7eHCDFsRbv+RZd4zv/LkbZzrdlujUteBTkLZXBxTEewwSfmaZdkT
tLoXbqjFNU+QZbMrQ2SDRsI5T4gDqehuKKeIrdEbauo3+rP6R4xVKO6JDQOVBCV9
DjOIt1qNNC9F2ACA3IDwlaS91BwZWuBPEN6pNkEmamS7RnaNRqY0AK93H7mODicN
K2wvcy6mOP3pn6Ulhym4ljrVRinSDs7mfkB+RI51mabY0JdpuFo3Xz+rSfiuon7m
pCEKzUpWfLfrk8VmQaoh9m6iTkEZTe0l1Pgt8xoUP399PXH2cQ9c0NU5F3bVaJNy
iFiuckn5cA7g5ORffBdfPnFeiftZHhSxy7Kse7iavO4OYve5jS9lp9Zc5s9CRR5L
2ON6jQNEnDpboAwfU23VyZrPg7PeUD6ra4AKeAYVh3ZxNS9pyNsbRaAiKJMLnDEf
yap3wkmYxPjDJOkzoTBy6MC7lkaf5C9MFQGwyCfCVVBdHmiSeo+s8kirLgawXxE0
DOB/an+VmZ7Js1nY3ZIeYSlJzDFj0de9wUjgI8GdRAJ0TGuIhozV9nvbyJz8IDep
XCrDv8q9wYsfkvRtbv7R9AiDIMrdiBMlvNhljtczsXv94Kyio/i5n/4fzn/6r2bY
vrhKNzfyZQN8uSpMF8AXa1ajy/RKgh9EroNwHeXXTpUDrbKOc+4Dtb+h/nQgN2LN
/sJrqladSkpUcxRpEC+KeRj38PvKPDb2lHhBwMvSgvx00vZ3Vxzj8tHJ9onhk7Vi
jBaK+mpj+1Uho7hPqAfjU7ymXz6wPjdt63CUD2C4n2A2wLkvUurHqejWw1o1Ojyd
QeLJ7Pr/XNE4kmQlyAtsVMMHctpNcuaCua9LGWotUato3Z5lEQthUOrNaAHq+cTG
B3abNSnskYHJNRiUPDx5MHy152sPpZZ9fh49yKxxUJICa4r3npe5akDohja4Koh6
ixzThtiPBApbtb8IZUfDilMC35nTJItRU5ByDEjpnyE7yM8U2VnDiv3fb62wt7D0
7IQkH2p+mRyqt+7y0BBRaoi/B+oIOp6Jm28kwlsyrFzEBj40a5cydy+horho8+uP
obeUOANHMZO5QMAHXCySfUnIIdAUOEHa6TaP7jpUQxJzTH7XdTOR+ym/p/CTFFRG
4tsD4vnImx38der5E3Mdf8dUWihH9R7QgP/DCLWC3zl8PeLDtpGPTADFDKXAMtkC
mHJ7HxrS//vSVuE4a5P9g5GcSpD9VM2anSy3ohgtyGMBvlFuB5cl8pWH8tIRfnWd
Az/HpZU9OpQF1b5ax3TBeA4t+GxrwR/PJsYcZlnyKSmwJARZpqTfdWsqFokcOt5N
cxnZPqvoaFizGyTfHb2Qm8uyZHjRr62TID3bc5FijN/jnrgSHpUiWqxq3UGLGQzZ
dOwDCGXz/y8G0rtp9D86DF6177uEi7AxXwUFUSLN6izhhOq3pARNIPKuCHIbWb2M
bXqBD1reW4s4TZxitHnhG9fYynmnlQk5nR1rTB1VWVp39AfoHpfQJghGv+r0MNPs
YHs27Z+rQa3Z7bERI0QemafKzFJHrPcDAmKEq4tX3DzMewzKsyMDROj7tis6V0vt
8qJGAYJG6XzBYKZjGDy8VW977MqQiIKxV8Nj5vWxGdZkZs42KOOtxPIkcuyi4X15
QbETAa5ydEpSGzPAbafy1SlVN+8HRuHf8vyLre75HyHi6l0NiRLzXHyOXXERxkgR
pti1fi19IlL5FyU1qWK6Zp5AucxmAo/P782XZ62HkjodB4vy0uqSSh/urKYG5eAE
NfwI8A1Em3tQnilmVBozGx+bLIHXUZu1O+qsIjCvC4ryV0noU4ez3TjbthAuEflV
FIBKQfmq93WA2K3i0jR/ulyEAmldiGgLBWFzooJ731SCH8abUASZsjKpX7S0bW1Y
lQhN7NvREdAd+Zg2Ilzt4Z8NXyv57rWhPS+cMCS/EXgb7W3/d0o46nSxfZa7KBi6
8zPy4ToKEDn7LJcF8l+7LAaBf68xPFeZslnQCbNiabLSDKev8dJDU8QvbmGzsAVq
53Q715g8mVQ8zh4TmPeQ9C7g2H3uWYljPK9RTEG0UFIIZzdnoBOe2rRN4TbW9k6f
YBsUemc7GllGE5B1aXcAf+2fhLOqRlhgxOshrGuBFA3PzHo9oNGLH/KmEtSceYNw
vod1pmzR65S3AZFsuP6N9pBqn/oq1K4dUn+vdI+ahg8i0keFQwGMrEr46zc51Jtt
bmnvTY94iB+ILlOX6OBlvl86SRAyoT77V1U8Qz2pTED9/gihHx+RugS6RbX26X9w
hGYuV5cEiQSlW98dw4WRPWon9r1AK9VhzidjyHKa5F3xYqBBdhBwxGH35dN2pDbj
2+XW6RJ9iCNrcV3LtYcGbyX7Fb/trNK6OlE1In8gYhjF+j/YZKO+npBqEwlnz81N
7JMGsH5lWs2WSsxxI+Cla1OJ8vM9SHg/81JxXC4TUYD2hCqsyDijH8p/8Ru8zr1N
mj8MtixsXFVDJ6/UyZ7LgCvzoRNiZlyrXSG7J2QVrlfdboDcRaH+pOqzRtKAnRrg
gF1KIFUcs3Wzt63Dd8jLOu8VwNAU/B3nyy+mZBIBeQg3XJd8Ic46KOu5Y5Ts9Qom
3IZAWJq5tY8LKyTVzvoJSbbdZ1pIwyUkMywMdrVQ8aONWMGgPVtwbVgHKOoiKOQz
K7X53qB/qZUG4jw0xKeetsD29wHJ4wUFIM4V4MZr3sVGwNqEz4U7i9llQ0Foh969
Py4CF1EYj99ZE5hcca1rw4FXTLGjICt0vJsxL3uXK0ngD3+AlIw7x7d2iOkCZURv
miyC8HY+MoDn3quSGa3U7hsV6EghhUpt1xqXbcNRCSVW1Mj2f+i970LiSELqJ5/l
37EyE+Cm+eqiDYkF50EnwoyoHZPk2OIeifL8etoPZ8Y9cIMvmNvLAdbFbP/BQFUn
5OGkIEAgP1EePGAcljwQ7NC2oyJ1WJrRBkv1fsk3I2plBh/RPnB4i2EvS5IqCIdk
uUEj5xHqSFD0zodA9EwlcNnDu3cKjxBA32uynjyFAy3zE6YxlvzbvvDepHOheQQc
Tw/CkzjGhzFHcpqWEpJ06F4EyTBcT+qHWApNpM261H0A89k9dphutgEySY/PErMi
7IMyVv0IpuBvDoqPtPU7c37d5Zon0vNsnavkPjQXS+fC+SzyKh2gyyDuxug0jyIK
gnxykkowgXC1vJXPrO0vmZMUxTPLwH9aKfagk9Qhl1bKwg0DwQrea2BHlD1g4xNR
kSAF0bL0p6EkaYi3wk5N3YljAhV5mFVnor9t9oSsoGd3n/sEj76anvGpAuxyhbrl
aE8tmtgzFSquJRn1GCGr+SMeQgIyD9VNxoJxgOV32LWhzGL9Pd7TViHs+Fk1W8Qt
nfH+oCpojYWzm84eOlarLDPpB0QGFxMeYsJf5NRygM9fKgpKNydJt7I6nM/Pxpwo
C4xDltvu8TiVp+hFowsre3nE7ZU21KN9VOlnPLUZk5jrI+xZvD5/4xLNhy3Wl5nw
+7vhAW+Z9WI/QOvLZn0pkuRETvKtVHWXRsThREYBO9Lqgr4gK76JAaZP8CdYcOto
58fe0mmle4yYITPmi++fcqFMwJ6aO1+cNgfojXEuero39rEGdLM1WuM3ppmnrk+f
Jmg0u9mBb7bZ6VoP23bWoB50vVqokr+DKDhH9mAq8t3rrMnzXS5p4XlkJzRNxbZi
FwvG0GCFu5OMiIE7HGipEWoP4x5XsIPlioxDs9v/rYscOYwxYt+tfVjy+6Ns/VDr
OY+qvtxoy0K2oUjPrMtjxoOHP6hUtoVOZS9eviBKpKtphpBUOdQKERGW581Acoyg
5LUPUpMkHbpXO8aNvgVjzHxofx77aa4MJhbvUtKFHxzOWL/ws59S6GF8xQWoEbnx
ZgPh95QQFejIxuqKsRayztHLihvSCzdiuwj6LFqIvh6jkLgw66OxBGF2qD/g/Yfw
7bRO3Vdz2gC96DxmiH4rRg5wQR/LrLn14D5CIAe7yrd4Y9q4R2nZNEsSiVRsiIsG
De/H8WUGPqI4YNfA+YN2cgE+NSnbdfhVnH8BVNjIDXZMnznzCnH+P6KrQ6Lua5C8
MInwAXVI2Is4hmLb/c4LMVI6dSMd8fqAXzpit8UQgdYNFTiaeIHTGoiKUftNju6G
akoFEQAGxeHjtisvFmehruZWDeyie/fT94nCBCI6vTsEwMZCe4HFj9CGb4WBS5ad
kPok8zg0k9LiqKJZ/es5JDBvj3Ytq54+RzcoJ9IKXm06yNCFlOBumTOVchRufyt6
doCjYEf0laZmNQfm7xJjFjYZGueEFi4Ws2gqqGyg76h7uQeOtuMCLKe1+GdsyZD8
mD5Ie/KsBdL2ovwQH+W6SGC0AIZczvGC5h+OCvsV6lkfON0cMa14CQnuAKS0z+VC
eztkoR8dehDer9KYPw24me5k5NK05VIT9ENZjh9U2XT+CFpRCaUrJIJI01BfSypL
8Wq0OoBB+VTaKySCM7+I2DuHXLfBY5BCGCwB9DabgFdaPtOb64lekuyweZ+blCXy
WJXvm/yoTh+CWQgjHXQzci5LsfAsRA3YtueafJsYfgou9wrw/tQiUOpY4X6pbMha
98ASOkMALOwDqyf7s2C/3vGOG67Hj0qWjAkUeVbzjvOExemkOhHHZTI4bQFrCAxX
RdH8NMWay052yBq7qOT0fC6XWVWUCdFkE0BCiUrSjCCE2zY5dKmvfHS/4ph6VqJ1
5zOTZldev75QVbE4K2VYJXOFgL9IINOo7TvTUX2dVqMao1cCFSk4hwN152wvwZ7C
ERmPXOtHbcaxLEELyIfHB4Iq0XgVNp1ZExeBnAR9xV8d1fZ0+m0PHzzli9jdTN3i
K4MtSVe+P7yz0GGj9ImFWo2e+0ugnkUB2BHT+q5TscLDsaBG/oM5VmIZ6bNWkA5D
Ru0ORmewf3A045YSzFE0c/cMQqA790HXM1e+zA9oYh+zcHbWhYFKxx67PW0fiisU
Iq0NIRL4W6qq3290exVOsRB1YeZvWNMuDPZsy/dVzF3OS2CSRR4B9Mp0Hhy3T8LJ
pqXjAzHyXJpA/ymjPuE03ag7iqdmMpw0w+JMGX0nKbGrVg3JZrNM7cu0FmSe0KS1
2UzvE9MMrc6r/kEwCxUkIctsFG8FVUskmddZJkwsBKmq5o8IgdG6BQHcJ1E7AqOH
8Sr1ruIEEVgtkMykm4EU3Dk4remGwSLuiTZ6k6Q+yJ8/5oCfdCByZQ3L5NCR/Ghf
pKEeyFe28SOubqYE/5Wc/h0s2Of921nfRkYJcjaed0n+HnaCQjb5+Uae9ygs+i5J
zfeXlh1yArFCk7tweoWnBgWP4zG3vch4VXPLlGfNSMVawWWAGizFSE91iivRTuHn
GAK6oAVls6dgORTo0LRAy9I6n2P9oAzgj55YECFgzt4aL8V9IiLpfUszk6SJuq1l
VB47gJWnE4oUsSint/9RxMN/N9TTlTCLEeT/ohpH50k5BQ+yNOVCfOIAEnyDSkoT
p3C33yBmSYd/NW9J2/lzlPva7SO4gS55I7wZV3psWUgBFbHoTjlx62b3U+on6F4r
5g7aG+MFroTbmVOy+qNdHXRrxaSZ/GWxPdHzL1C3lf+ho4RkKNBJPkBA2LWPTrkm
0VJ1G3edEHwYGl1bwQLU4B21ZLUUnHXhwBR7NHAkhR/A1j5nVCUKwPo4J5ONe9AK
NvhqezXGt3EU5pXl4KY4CzeSS5FUxDkAF4jMGVH4q2bCNJnYz3KsWynCR6gedwpg
lyUFOOjg1wuRhqHY4Cn7m/7/YtmlTAFZc3soRLq45jrp4aVhfUdl78kxJX+oJ/Qb
xesou9cjIKF6OL/rZbxkf7cRrdysn/pi2DyrRJvCj/ItxkmVmBjnVsTVZXph1uGU
+FYJdh3SbrT9KpxR1+781eWyP6Gsd314shE9juK9To2KxIPxGdeiSGYLzaoMIzXj
836y1AvpOpzbjB/fglQa3nUAHCwCq4J5CdgNeuVLS2fP2jckbmae85D7C4CSEX+L
W6jQG7oslya8OJptxz3pS9nioaYCfafwkwJV2B7qyBg7jq/sDyDyncB4IuQysXEp
zyMV7LkPL/nOWOQygywwqoLZIaFhG4lo2tJ9vL9hDBahrxUeO38ZjB6QoT5v0Srb
i41aS7ZYHmhUPL3B1rZH/pjUxuU7Z1P+vCQGieMuDvywzgJMlt7OOgHuVRVqAy5C
mTWViuE3DAA7lcA1SQmvesp6G06FD9xCW/kC4kzMhqW6VIxnRgraoVfMXHRubnQ0
30gsIAQiraWqjd1aR/gaq+cYtGSZbSoIsbBoQDV+wz3uRzPTLpO6HL+4BeVCBf7c
b2gqERLsQpwea1AjRd5l6kYvzd5/aLSKE9XBQdKsmlitIK4AeL5zBzS29Anvl/+z
aJ2mJ5SiB8j6FLUEE4piqdwdWUrUUI9qLCOIGWbT+3W0AVzMuT4RICxYJFbY2Ay5
QORBV0ijL/Beohxfj7ybJe0Mph+k2h2mYDSgrYwMeyimJRz/LXSJpxHkHkMhu72a
cmtCDL9xmULOavjnesnoLvGB+iO64AjUmdUOFmi0rpGkzkcHvalaNQS4qfuapE5K
G8vAU4dkawTVKxRLI3FnsWNVTbL53XUaCNVq4Ny2pnHWwvMMmQw7cB4sns335yPg
c8VBaybKdza+jmsdz6x4YXW1pJ3niA1cXI5ReQQNUqWCeX4B6RXdKQG+//NEy7BU
1KkRu2mT2jq5Qk/UIRswRCiVOsSE3excv+OozE5qg5xQiJ6qWLhYE05VZeipI0gH
uncpdKJv9PyzNdSGgWUZxczM+iqtuAhqvzdCHiQBPgWwmXrjf/et8wd+viDq7PK/
uYIru5BNRQN1s85zxAdgeT4NkR65KJGYZSXqWUBqzO1mB7tz3LBD93VDynX7zdV5
KQvI4gFnOAgzkxLFHYYflcjHwlYz3Lm/e6czo3RzTNFZ8Ox/SXKMJUbkKD/xRpRW
6VclrBNaH4K/suTjazRrbtTYSZFlEP+4gDsRXV2ONGEt590JUgh4y2uzNHaQtcmj
iM4uDRNh5+E7EfNIwoSy91kztZdu9ZKYGaU+hvdHXbygY7MNvhjd7g+XgQZSBZ0a
+SjQ1IA9VdFxtmvN+EH3xnJxeLk0aFwI+b1ClW7wraqNWqVjX9zIzI6yT2X5dapt
w2WxWH87b0QeguMqmbLEhsGwZrqW98h3jmCMK2/zqWo0QiiNY9ls/fpzHlFlUXJE
d+qOWstb7AHciz46ODakY1IBp8mUO8QAwxmqoZSl2gXWTIZUnkI4alPUH0NuHR5f
9RlUiO2Nq0uggLoekLo0CGIkpj35tcPirZiMJg9xf4jEzQFvimm1RFZ++QYnjntd
d3ldhUdVabnJoS1GQILTXJHfWWCXO+hRGUQl7hYNJNXNO8OETBpXJpjcU8i5v297
oQ8Trj3/hjhcH2feAITGREvKd4roOgLDiIMZnL1MzrsIm3hWLDcwVcQQhxfEc3aI
Qfr4rs4TyTOnBIRrFvsaiqF5T7XgB/HXm/43MrW3qe9hxJWJ8sWqn/jKEjfd/kaI
14zRCIfepIAGAoGWCpeZA+Y5utK1OByM9BnkCalZs3U71HTyN8lUPepO+UcxVbQp
r1dov+4qUiPsTdJQaXQS9VL5CfJsxV8yPrXhBiNThxTz1xCc7aUK1E5zvYlcNGzP
geuh6kzmq+srJZxDMEpHzm73SN34kh9cx5Pg0q6mmauN7xLniSWLHOHXBBACl3hx
l71A6oXEaAYTbrOyMugQq/DsOrpgm3NFgutJrijSNY8GpdR3ftvL6dWY5o6kxamY
SJ4/GOSQqhwmAFRAsxFxOMBkGKOEqMc7zHmhc+oDehyB4X3B4zBFeemPhfZeJ/xV
q+Y7AaMtNDsdwhYIqLEIDp4hDXz5KH5bbVTI8xtRcZxoVuxMdPbYtyd3RslDquJF
XYnjOptpGS8NnhVQ3c1m6yd+C+6R3/UUUKncY3qM93KWLZXwViuglBb17V+xd5tr
rc7o4Ics4WZl1CuRM+HptGFz//kW/ynJE98jhcO3P3qnZ64cBOjTEVCgfbuOAK8b
8x13tkcp9t4aX0NKnuKHdrXGm3P1CElzWiw5hAq0K9rKl8b6mpNeP9xosop7lpSO
SVXBJBD+1X9SeLti9t1ZDM1p6WT7imF8LYElkS3XpkSovYrd8y3MvyGcb7jy1DW+
LmKeUL9uSiZsmJhTWTVqkfwIPoGvSgJvNW6LZy4bW3Eo/eU+qoyRdVqcC0reYeSr
catv7/Umsy7kFyv4cfhtFcObaBXzR7U7UEx7SSvNzsfm7+4jBJujBM1mEDCblAZH
ymGnn3gNZO8NtOrWYYLD1jExUvLrDIy6OrBAWHVwji3adhbrc7nWruJe6Nvr86H+
1WJl0QeTref9lPp0wLLLs3OU+Z24LnetZC4wxqVOlBMtPaAaqzF+jFCSNC+xTUfa
heOhaoZU4dp+5GKZIJdjc3wY4boxYmNI1rYJ7VARjQMpuc/jtTAk1/O+sw4UPfXP
CRekVlunJ8mRDHr0TOZq1ghgYVc5wId6QyoTxTro9fQ+oE1XA76cmJBy23O5JRJX
/uDblOoVoS4TWJ6E2h5pgE5oDmOwPzCFTIIV8uMdez8nQzPgTFvSRdNnuxKzxJpk
YRuZ7w7E/zT4F8HUuHtSoi4jjmmUTtT1Npjt9qHotj68Jk5USPsKN4Sy6e67X7V5
Zzr4uG5jMc1oDf6INB30Rgpha6qMdOTUHHlUNlVlswmoMxwNcfK8LPI1ipTKkPhj
BeoOkQgEqu8nnDAvajD2lBctmRizo5KEHuANvhtUJebegy7cq4o4YIqMG+GG1hff
VnfBsWnkdW4GlobnKHCcxZVEkAe+1d4ZYPFZ4pAS8CFIhH/+I+c2iXGDfMRuwgu6
9dbvfSxGGhn+eFCcutaNa2BQjCrYI1dDX9t0mz/cixqI8jcoTFVI7Er+VkzgAoWS
IP0Op3q8GFtO6jVNfcM30S0XFaG9/vnZqReQom0XUn/iAXYt4aO/A3Nsf3aOnhCH
e90HNZMc99ZJ8/hexXJyFh0KnRMpfPjn0zftbngoU78+mc8yE8b26Obui0R4htCQ
4we8SGi2qqLyhWAtLyAk09ULC/ZkHds63pwn8TDVD3kT8/FchJp0+vPNugqtKRRd
L/hlq+NzemaeVInLlipwPjfUOs2js8dn1RdcWSc5/R6aCwRxm79A1/lcLWii/GXA
YuOxyQBQtNY5HYuwlQ1sEe0uaJ5qjDvpXUxCsqEamayhBtsG/FOXVVtw0H9T+3ad
flAmtUH2ATgLgeXYY2W+pXoYjExrcQz6DzmHc7pTkErH7EoKA9D9QVBsnOKQTqxy
IPIxp0CpahrDX00r91ntWZWXZMA+M+jlXbF371zhxTIPdL2nUGbNLOqmKNHKLYPi
uT5ekmd/oSResXBUlcE6T+T55uXKJSFxq1vi2V+c3G3xSXvU8dBDOEjGg1ZSvRNJ
TiUTDSoVg/zQAkn9clRlqdAYMAQ5XCFlAfNOO9ICO9aln1huSwDuL7UCbM3/9NzH
tRRwCatIdYjc4BSNAwD7NTaVnZ9l4iVRBPGCuVZO/9AevaYCpebWKEZCRMrHiSvy
/IA5oENqnF8BOrIhPnCBVLC9W5cOa+W9sIoRoq/TFxnCqBmRJGPcvaIs6nOYCght
+U4gSogu+xTcjSeJvtO9q8/P9+qcTwy2B96fa9bLsOIuTo16Xsq5W2XmSN2NkiUC
bIl559Kvu265lyvtaXebYijhiEoN/v9irRTrb00MZcciNyi+mhChIKIkrkWDy/bJ
7j8RiHI3kfB6DpsVss1MXHLgfm9kASJr8H0n8bozgotZe0tlyZMHGnsF44BiUQQ3
NJOcMXT8EIN1OTGl+2NFIpUdx7E1PqQ29G2jbHx9gIs9TZw23xfnElO5xDDjUPuq
X8C21ObYJcrXDK30NFTPhboldLGD9VYCkjs9/vdlU5omTWc6cW7JSIqeINWchDrD
X+QSfu7OJlgUVNcvKXbUKibHYuo+r+7v9f0NLcGqcg06gkC6JFrbURk2ADVDQB0W
NbDAejAqKPI93DELP8DATTSn6xc/6LtStvbcCvGxACTKCQWorSk8UE+itKtU0j6y
qDp2vOfk8UY54uMI6+CKWn27eTSuBMLDp/Fuy2t9v1gSmnkdnbm4iJjQjDdv3KaR
WTbnrs2hdWgVoRNO2haR7XU9nIYD0FUicZRetjJvce/P5SYW0awEGxVjMhlqESxZ
q+cnL6IrenO8/XMzHgTcxH+RSnQbXBr4vhqEAPPFvaABcsBBlAcTY5CzZFC2segG
aRp2RZkVA3e39r3uCHssS51F+sg6qoDf3aiS2NV5zQ//U0Ib45/ujgu8xIttEQcA
1h5IyOT+bP6AzTxKlfkO2kBkiJ3IzD4rDV6ydFjMKHmFbPwqeJIcjC6vJ8bcFxje
DXG3SIf1xNTWF8s73ClOn4jLOsaY/NnPwDrq6vYx2aookLLO4FWIisE4+HlS1chg
DOcEU/DAb5VjBDhVHwo1ur6ke0hOKgn4O9gsRfAXWmP0oyEjxqCwQxSQI6cS/mWa
iBQqHQySUVL9/0/KuWzeY1tH8GtU0Uzu4NhlN9M3pK3QXP13iyA9156OXTiV3/dH
kTRuz8Da1bWGEFI8AQF4NBm4IEvIerA/5dJCS9HHc8A6c/cWNbAHHDqMDxxJabK0
hGV/q2q2LjH3IYmcWVqK9piCngHHkqzH1usawqQrmUa0r4XD2IuIfmQaJCO2+zUT
vaZbwBQGlUNMkM7uI6fhArUIUtTFN7hmvsW9VaCnWOwUMErpqmCa2DjLte9i8KSS
hvi9+ngK9OwIV7r8ahNwduSIaNXE4kASMnibhNpp211LGZggbzqUeQj8Sptt4tFg
F9LTlbZjU1jbxMVA9PvEm2db3sqPh6qeBskVyDq0zLsb+/VJ+HWHyMiIZVmLRvcp
Iywm+/Y/d+JPi9B4bxLPZXhjWxDxNFJOZbB5KG3YcKWBBizqpZ319KDI5FcSVIj1
Cwimhe/fH2edYYAE/U8hDfka4z/zPYbgec+ND8bCyDS/7aBOQrIwgqObsz8VLJNm
6U7ReLjLZQyR5dl4LILEoQd1LBqrgljwSyzaK1hQgh4cS6R8BWN5Dfb4N6F1IALJ
dxqZ7Kr+DuJRfOyL1cpIyp6ru6sUXockPz8fLQl1XWM2ydRDoQiZNrA05FrNcel3
NYE3ddGZ3Dyv4mehYyON++fAJbfxQF145RUFHw6lvYBbT+lpfMhhxJIq2GGNeUpO
VctuPzdf34RZ295hCnXTm955+qBUUIlobaAHAE6S7kT4d7D20Bu6zGkTecqzbASl
6Ih84KBRKwcaDQ3blFbDT/M25mHMzL61vpbhFce4hYUXMGB0rafx2DAY14JSiXls
XdS/+5nIHiShMeIz6pjZGByhvF8CxN8Ytcyinx8GfyleTUSCn0btA4nPbqGWX2oI
Xir536vu2hyedSqc+W+3+csn9lRVDVaNVH0GHKW8AwYcnFNIfPhetoR8T75Yr649
gpzmONv4iEhtNM4t9mxrERkOvy+fZIsi9FKSnNvg+3wlU+kf9C8W3H/xVhVDDyUM
vfZ57cBDy95pGRf+I2NoU4F09LEqCzhPVCcGhmA6Hi/293i34OEjP8JxW4FdYmrP
DXvUqoP/InW0kX9ifR6bVEqyctjAH7U6MIXsNQKUzGFapMBEgRPN4QdDB/bRBKU2
hJU7ob5fLKeE+bcxUUxtqQiplQyRZqQwFGJKvOH2Rkefb5RNuq6v6sYIaXT5NWPC
DFVdaDWKJg1cZqNldq+QJuVHmuX6j1TvnFUWVYe61SPXPTTdqotIp7iV1tyPjDrR
ar8MFFuLKBdMmVoxKI4SNvFIyySuFNvZ1Nuv9TYchKAYOk9P8OIPsZbAIqP1QWhh
5oTkqqqkLeROzlGIeQL97tYnEtJ+naE9wnnm8Rj7cNhToIhX9Khib93KAq7Lpc+e
I35uXqrhVc4PvQafNCF7S69Jzqsn0CeXeibakRVHqKX/S7M405BAfiiH05hEZA1U
zsl0b/PHMUIP0qAjFj5JzoI4Jy8lQtC/OhXaZaaKPeR4aLQ/BsNTAbElzwt/kS19
0kuoxNvOVnExx0VpjVwb6mdyy7MZS0LqCNdIGnGwfKkLk0jV/XtLTtjkXNZpApUA
zTTMnZYaaVJG/Ww2uXricNGQWOcuXS8edYlyp7PhcjLq8d7/myzq2oTnLSAi+D//
hQ2H/5EXOF40Z27G4s+sttS/pGK6SVut9Cs+2s9EI0G4/I0BCA6vEwfWpqf35i47
S8vvY/gYDYQoRDv429fLb18m2+XB44uqfGvDKvkkA76xUMDEVQi9xj9I5eI56vNg
ZmV3/xXuaMbxmMr4CgPGBUMsnvUs8SrFObItUgd3w0yTA1ExOWm4X9IAaWWZqXL5
52XPL9jxUmssoSAjF1YuA3pPYPl/0ILhwpFQo9ZRpZYIGqxC8HVGa+7tBQecuOs0
CRtNs0uhkqeqy7r5OwfNZx/ddFMk7QV8JRiidjE6g4yaedp8r3oiOkZN4wlPyuSU
SyhtnP40ASR3mvxwUAnVt31S+cKG/hvoR3VnnomzexRC4CTAWEHaC0RoRQpRuPw/
CVX5O7W9A0Y2F8uB1aOLPPeO8yQ4suhcamckwQk4atAnlGy+QU53DGE3dIdrx3nO
GeyVHxTtt/lRnrMPixEPxS89innDQmqgDu2ybgZW3uJFGV8xQfNVEx37vz7Xb3b/
DSjczRC3ni7ntSmXwo90ElakE+O2DWbUgUh4I6qgADQNbhcESM5HzNEWLWrOTWin
dYo0m6S9pIm5zza8GqhacYyBMF00vtE7MggdyYacuu6HT0pYx4uOX+9IpsVW5hgs
3A6rU7o1x+W9IBGA4uKsWY0J6fOjxChqXViO0Wd1l7yFLNyOC/NISieI3NHPCpSb
DKOhqvW+acW/ubNcrxU4bO0Aj3ATjCffUqq8TJ7RKekqodnOVQglDgoX+Jvrmbe6
eU2ug9AK4tXmWsdfcyTUuEx/niPjkCPh4U02L7Jlkgb7i7MkHeDQ/TWU41nNNCev
b9XK/hR8a9kHnwkGL3kQgzizZTOoh9KuTY9eikxcyBwzIAF+yatMioq3u7wXCnPB
NAyl2m0VbUnu5z7Q3R0NQbT8pgX9x9tVmop+ATKTUHzUFRg4G1xh7woG1UUVA2t0
nPYgrxNqM3FLyIzFV4n1TOWtDMjZGbbcMi/3//ElBI/VOZEIU8KeK4yQ1zao/nTZ
6GvnALQ4HpcWtAV3K2Rl0Bc5m5EFExxkrfCTLLj/+PBS7h1yGHcZI4gj9efe1lJs
Ruhdv+soj+DyW2n090993vKjyCWQbiFHQv5Oikq2wV0f1c6vH6r/wl+BBzoS3UGL
lEiZGUs9VAJZLRFm2HccFZ1dG3UQQ+r9i8LIirhpTtPADF1tIjWgo02vxIQbGd8V
OgXMNu+SSttWvxaowQ8betF33YjPrksM3eN31aOgluvmO0xB9lgpUkbSNmpR0FNO
P09/HAI4GFzONNAyMjOp1GjUtopaLEYtERDx9dL8dWoDGFse4wRCnlo7zLgkTiDr
X4UoYJRJmpNbnpIr8Irrfns64bPSV7Rb7A7bIbR/j0zdZshnRC8xrHzvwz0HcgpV
Xm2cNPPNrPbwv2KBtJ7onf0baaI71dR2JoqObxEEkJFYWWrW3kmtzIlAxU30U4a9
UcSuWg6DKDV0MS0GlY0LMaRprf/V0JuFK58SmxvOn4eyyJG7wsDPVNzyzbr9dLCO
ZmmH+WedXzrZiZgGwefRZagFim0hAOSy4s7BmqTfVbgrJrkn+JSQFE0I26C8l7TE
mhnyCgNnvdsWYsycMNhl8aJ6FcgFUc+2G+9BOvXohx7dh4cL8DEdC4AJn40urjJV
JA58TQq6vyInezNE3Ou+Q4U3Lvv6Mv/XhQPiPW+qaqFteyRLUK/AYEe2qZQgyPG7
ud7VYpZvaxSYDzFV7sdApOmEfMXPUIVKdpIPBaalsAPq0VZWWngtguFmLf77c1QP
6XP+xCtKs6S/uw3f//vTGfoczv3PUOmf+bGPLDNOHRLOC550f//wW1YszwlnSmWP
Tg922UV+Jp/RPsb60pnhIBz/p9AixcL2cFq2JPo4L4RI2gyDV3kaFJu7VdVa5dN1
t12i4zzF8Nhq+IqCFZgrRInfEa940nfRPVUH91zZVWp6IFCuXQthvC1oU4m5xHYE
7X5LeWZNFQQyzwSE7fzT8YWRFrXH9VjCo7q47hAnjqZYHpWsdJGDEjsyeKHLh5F5
bgJ9fVkpgmBWKE+6kYi86v0Bq6sWdYPkHwpVFFKTnFDbmzgjU03XB1OfVCPFggAx
I9SXkRx+OnRRCY0Pd2GYsyuDm+LubgCWuElXZk/af2iI3GiaU/nJ/eioORmuPCaY
CTX1Rq0f3A+q1ayaJp9uZskL43Yp4Sktwu6n4IghZHvr1CQ7NFu9/DJhS9QDDH3v
0XpumBR9uE+LOnERESzG4+V5+JrSR7HfvzSnbnYjgy4rQoPze/PGhP8PremrK30p
eKxGabwzzv7pDOKrkXcU6MfxYRpuqqLSLdjBjXmrfB/DgoMfGwtt13WIbUm4hvEH
/NDhtirE1QFo/KRVVUhhZArGsiAYpXxgnmPWPlmX22uTDt0m07++uxscNm443X/0
0vvriMQSFbYwMd39cX+u4v/SoB/9YUftQdgoucuNQw90Ihy40FPl2Jn3mW1vEE79
KtSnuusRt0rTHJeIOP7eDZ28GNoPhJBLAJstYuGupgBiVvgFvGUnGMRSPx5jzT7D
neCNw4gJok1028FN2PJ5ZRbiU83RyMLNVlWCqYxqEOgAN+BvsOTfdLWUwP6/ba5v
kE26pU9RVG3OUJLAlEkB1wKxCMHHyY2YKmZk50/F+XTcaKbZWEVbxuvDFEyQA8Xh
OwhJpLF1eVzhXoIT+a7MkwIOcSPueKl0M8UciJbTnpADupbJIzLozqTBwEF4rsIs
tzV8/YhZHwailpzbDEmRXQ4jYTFtdERUCJaN8rKmsEzzSY9CVrTcWHRIkpWhoc9N
nG1Fo6KArgnWW/o5m2pb4N83wYrQR0Ztx7bFi5TJwz4OXK0L8+rHU5Cm5/kcqs6R
lSu0HJxMTBy2B9ytRVvkevamoMgtbLtjbKx3R8DDfv8hBysiNRDzohEwyo0WSwtX
GY6lZgPx9nASOauw/J0hKMLgI7MWSayzpvHhdUChGxDYwB6lo28Nrhd+k3YipA5b
R86AwbhY0Sr2qVQZufdrT87tV/8myYzdAxmfyA+9TCmETDAfm+xhtDedxxcs0RBN
OR7tabFeuaTcthPs4PIkkYROpFuBm51sgG8kMgwY4PoKCCpsrUIvcFJEcwPD9NpD
s05geIfLNgG4WZ+N2707qtKW2iWYaX579BwEPAUmMGJIgt99uC+CDhwexDuKOmiG
Q+FTRoMju49Moz4BddryfGA/MvpDWLaqt4yw4dPVmDzvfZ+TsG+SqyB+f0VYYK8S
PWW0imvaHwGa2g9BtRmdc3VBumlIVceSD3KLeut8VyWPWnafP69isEICK343aUsM
aROG7bGnYPsdbStubJqjpUkn0Njfbau9nYSVzF2tlS5QmAZTeZS4w65j3MRbEqKi
5mLH59bHjL7Rl2GBnnCk7w==

`pragma protect end_protected
