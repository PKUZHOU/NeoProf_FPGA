// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uvDF8lC7aMHepFtYhTmBlSmfBfbGOy2nyUNz4BH2hY5CBLKWmiCO/9oxThpW
19HiBAVi5PA41mEYsDqz+JsKOcHRzOPKmPnBWJW5wKacm5LADvOIda9n4cQo
hqOrrNplvx553Z/oxh1KtpgAFL4YWqG7ph6QdaHtQa4Rb0jaQhWH28L/+NRW
aUWQpRpBw0bs+BWk0t8bqM7dE45SNhTWatnrr+JJS1znlSokc3pvMVNrxTSu
2lgX/fBkjfLymAwfcozvHszUVRotlVuQI+6WIA2Di3UnmgudRAQ3L6RxE6Sz
p+l2sti+XDbNIEzh0N7ALfrznfS3UB7v7EnUopNCvQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UplHfuOp5x65PEGE/5VKbmzzf3TWbeEXBw/TcEqwp5+qno+N6JOJlTJXjWqS
NS0Bb7dbo9MITirXyS9Y4GjiaMvVGgyvYb1JJsDNnGDGbxLn1Mtrkg5P4tlW
A5JXq/lWNoFBVjFzVWdKUIfBBekOSot33tNirIUlcMIV2SYJOM0v0xOP3Epq
TVBzdTqeAly6m0PfwIj+ocfNhMhaCATFOsoSWtLNXrEGGV4tUPmqvY+nJc1e
BBVA16FsNWRs8vhi0iObqyvICSRfnoK1MsvdZw+rbSbSNSUmAwgg2gNgKLJU
jBSWXMU3Z13IdgztLrt9CUocd0IIq0RwcF96tQmz6g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Zor1EMb47NTFSP88tJ0F2XGqmCrbqLUjGRnXIIN22Arhnd3kS5Tcoqv65Vv7
DB55L3ss9QWrGfTjvpDxTq1zZPCpDiGM3tUgl/bRvb4yrqcVTDKLlh9c5BQN
G6Zm7FIBvbn1TNKuhT1uySMwCSDqs4M7OhehmvnI+8GNqZCC8Z5CkFweGvQW
THIQfLItFhAV1IV8kO2T0xecguIyh7qbKoD586fAByCkhyOazZeOXt/PvD5X
iwo7EHHnaGAatjj8uE5sAOLvmrl8vOqDgOB1fR/ncSxMr2JbTC6ULxuKtfew
LfwCMHvcZocQKJGXieIyJJ7+tjcte9zuKDhLWDjK/w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Teug2x3/B375AHeEU2eQ0NStSyj1b6N2CA0vRRDjKSSFRROGOpK902zF3GSj
ZNk+8yMDDIl2Yrop+C32c/4LRjkomWFNl2hT8BNLe5LS0DzLWZ7+C7Q4SpnJ
Va2Hdj7j9GZb/cTIRPVL9Bx4U1yAeCnXSLz9KabVvSsDDOghwbY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SGm5u/SzIdIAQxRcTd/zYaPPn0QFnYITZA+dp4rri5SnhcwUixvq8QpJ85Eo
r1IMNLA9/Rajd2dGgkfOqzsCOSbFwUdlxUxaB7i25/G/0VRYm8ipxxEehX6I
ExmIH0ybIDhw2AuUmZffn7o7h7b/vmn/9gzUX7RGmP+4GM7QK9duTIpQcboJ
BL0IXsDZOQGjQv5/xdOjH2/nYT9VP81MAK1nCNseMNWfCOFiW0Q/4Mk9TOrd
OJ89dDg7VmkSguaq2Q8iyj87ZyiTARL3HZA0LizCpfUYkDlMKWDIfLpUKjvQ
Rxzk/a58t+nE2zVxMuUqX9+Epm3S6VprjcM4BsZ24BPAmVD432/Ccv18WGLF
W+Zv2KWfiog3xIzzISRBgs1Kmduw78Fgd/pSUDYFdiMs3Si95pPQOo0qFo7a
bGPuWQOJZzEc1BdiP9pFvKl3pvJRAQGVA/Q840yMq0sSXcPSwwTPcARQ+leO
ZBh3JCcwJB60rqgRxVzESkui3lLa0h3w


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dmfWtgZLzRwUOacQtoV+3bYYrg+hMZGvVYk/jM2/N5fli3wMqRe6sDZCrhKv
MYkDfqxNFgBSS6yy4p7cEnRtcJ95vnTA7IWzknpGu1iqQmYjYyFwM9YX1tHo
AXq7PIdv75Kb/NT8N37k4Nj7k7WUf7g1mzO4Y841YijHo0BP/6Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hpcztpkHNm8a7Sf0sK76Fyiexvn9xEKEvyrI5CRoTSYdH9u8fWRW6/NobqOn
EHdwmnmIMkTx+6n3OAz8wvh45tmWyYG6trZg8TZZaguZlAJCHJDOFqX7Bx5Z
1yvzZQ5Y4HxLyjdQcAJkg6wzS9tl/Qga01rLKZx37O2A6G5otrI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 150944)
`pragma protect data_block
FlfRQyb3wTGsN72YNT9slVmLUKZvnNjD807LcjwSfPYxVoc52C6NOatcVo7F
mVsVAcxYzTitfO2JTG1w260RsrB07+6B0NMf7/D4FZdOtVT4bBQgSOnkqAIc
t0EhXPBQlBL/xs8vlplyV3+UASsPkwp+8UH5YT125ahBLBxS+Zy6Oe1hUgtN
6iXbJ1Lp7kMVb4jJZn08DPMvxrXgGW3vM6nABZxLoK5LycWEzD2mPuFL5tNn
/IrV/Ra+GOKivW/Ba2BO+64bL8rNdIexiv2qHnYI2qMYQkr46/cHsIduSHzR
O4L90yqvpJX9gAOLS9i6mc9OVEWtdWNyxEiQ+VdTWl/SF8UFC5MKM9eh8emt
47pS3wHnb6alSgDko/dG8ODj3vIjfI6U5BmCgfRqEk6ldOpHTKiRHyEVrtA7
w1DalHvmIdubWsPRTHKa2fLvf9JTO3EX2eOHu87TevInR5Tt3SUMLCB65Dco
DpABpP2UbQfY++qJbmuNBs0GybsEwvkAWEEsJCV1OIpG+6SLjPEsqi0hJb3S
FkXQqVO4J/7N/7S+t5emgsgJHOfYgRocuNDWhhfm+aP5vJChtNvg8pG2alvs
Jopzo29njegqsCD3IqMKKitCBwFOORU6uPKmVCHmcHT4rQCIIC0X8wMjb3eK
TA8IOcHQUC8vVCqG1Ndonc3bPiAFeE1CmrWhmWNiAdbh/DdzN3F/J9nzepN+
2nhY9zJvBE89L2cM5il5tJ98B6R1VWa9qgFVHHzlEh0vYc40RMZ3h6mY9cgj
ZOcBsIRfcwY699em45f1oidSBBogDZAsLAioserlknu+6A9PxwGX+IUVUePO
cEQV7+jDgMYITsB7LtsKvyLdkv4prXodMQ4dkUzD8hXFlAvParuEK5/6I9Pq
qMjfxzUi5Hj+BmIDYTXDwUEfV6phDteohkQzDMGcmhyynT0b28UD1H80TExb
w2eNnoJfR2LrZhGXI1sLdYXr/+oPAWW2SGh117NYduvUuwtcwleKO7dorrlZ
knrM/Ts6EohsPHGfL3U9DpYmcdcs9z409J2/bkFRwYRPJyElz0Im2SgNBDal
F4yZAeL+aF9U3pSLePmBQUYYBReez6RPnk6gkWU4PRvhk8BrYxRFlQX2/oW7
eS9QFlN0+SimISA44YEtue4UONXSs82Mo+rJ1Lfnrng3igAFz+mf/woi9aKB
yhAyIEgYJSMPxuZGwBty4XwqTP1y0iks7Ppdi50xcfq0AriZcEOcd+9tJ80Z
LYO8Ta1RDEc9rdkyQovxzp9RCzPQaaqVpmsQtyinQxGCwwzxnYGIol3ksILS
/Xae3v5If9bN//1/IyoJyaNiN7V8CNC5J60nt3lHmGJTCnrUy0qwTDYuAmbu
j7RCYGZXlDE4pUG2BwNtZj9VQfO7nxfQCmtiR47qKBj5W7Iq8lsvpuFFAbvB
xjFKVfLnsdEbpd+N8mLekeew3MyntXHcSxvlJLW1kKNi1uTxLRtXY40jAKoA
3krfUI/gC1O0Iz/rDr3HMocEUZSNuQF/9gt6NMUUn9+VVKdgmrQVu478zeqz
nc2TDq3OCYUX2A3zzmAj7rsMiW/ysMj0axPzzVxGoIIzPbXf5GTWCteCPyIs
Gev3Oa6yNjsuDmOJY1qptDBagMXgC0gUb+ymDUN2c7NsbpGs4VsOvtII6nmE
AitUtAWysPUVT8U4qmuBVIWc1tJkMr3noWOsf6zo6pu36z+CAb8bcTvv7MQ3
5NWh0clWf6aq5GidH5ZZ96127Je36JIQddiLZPpRn0Qfrpuq7QJFUF25kGaJ
2wAIMptUJb4VN0LwFn96VvqbiGLFO0Z+Otx3x1DQRnOPaQ7SlKijrlq94znn
LdQBngyM2ApqphGHRGVguCzX6O6a/8B3roU3il7pPGu3I7uGRReR9HzXD0R/
37bF2ktFS8jC4GPvI/cxi851bEWI0ZS8lqgo8L6uOrNCqMGwQnu8P8VFjX7h
GcBeejNhJ1HK/vniTu0jBSx8TO/RkUlyF+DJZDO4/LBqzYzxpn/6An1jhDuE
rehc4ykl68IxMh0MtDXCUf9Ye/f9YszRMKd65MRLWnjXE/uzTfYcE3QEZcBH
hDmDvQnRx5ho2PgtAcgVWNWNgXfbDGWGADx44EF0EDejpEZdazFIwJEm52p1
o2P+gDkvPyLWwMqTpchW8vsMMCs4R/EZXcU2QkQ9tfeL4mC0p27KQVBdZ2He
LL1QmP6FvKcgP4s45E0opctWtpLH3AEcerUcKYQls3q2ffNHNKkZsTlnHicD
oD4ktjSEPMYdYBam597uWAfmF9p5uHRXNnomF353X5d9QuCLz+NLmtTNb/lW
2ILM4H6GcvHprwB2alyM7C9kX/uz6RjgSv2qjuZLH/Pv3p9upr4RgDo5lm7/
CjCjdzJ1rRMeylRw1VMGMQNcvnrdziqL/U4vr0kqpVLsUrhKZoIPBt4bRbo2
CvHXaWTZGFo/O6DSakpQd142VKzpZV2h3/OSMfZRQFOZ6C7QdcCzPx1TbjGf
VLoeK54wNoJKDELFP8NEcee/6GcOw+cTemTuyyBbB19XCfVz0lRv6cVo4BTF
0/BrAC4tj5XsL/M6XjfC2ZT+Hk7UNtbUxWteqnOYM/VzQjob/l9YEAHNDJVR
awSP4a2wTeSf5jOJ0xaVagCRYMTTfXPyFp89q8ZtQ+UBVtl8QYw7I+IT1igF
QIcvzZgNn0YeKSZTNCA+fC4K4OmQ9HdQXLUn8mumnSygy42Q0VhNeTxsNH5e
EU3PANnaILP7MEAi+xZmEMZGnLM/Wcorvs9OW9rLOuRwN7//j6sU8x9czHh4
4eq5D9QaOUSnIufY7jsJADjagSqosz4mrCG54xIqLWY3tX7OfoHY9UT6wX1B
wLrZaynqq+asXiMIf0Qqi2nxf+/4IwQ8DE81wq2CieP00ngv44TKZOpe/Ap4
yiuAnJUH9eMTO1wtt+p6jy6+1YQBR5pXNOnyyyO5/RUnsfrCTX008Qwd0IL4
U69GPfP2UbkuW/eumG4AggCGsuQoNcae+HZY2BWV0U4NW1IzGtfCZ+0nhdvu
1rnxN90SnBlCknMUHZC5pNNXo33a/Hr9lspDWYFvII1h0vF7mKITfP/qmk1b
dWB8DMBlyOHHdNx9MSQWl2AnlOoicvbQoT6Hsqf3t0yDvfN90ebK1yuIavnQ
1zc9hYSIhmfOfjEGYxzj413LGOrdyOdm27ZpyBaYAhbZadrfHbh+5jvL+NWv
AmiQIiopCjbMoJG13b3oZzoYniutDfah7r2XGJfecJiGETZc8Behvxex7v9e
Fpw4mdh89mMKX96CurpN6P7wl11v3mZY6uegP8q3dnpeYZdUJRkntbq6lvZ/
WHUcZJ04+cGE4Bemgr2CqcuelrbsmMobnAwKB7nNPBVmTFd2ji1vvlVDkhzx
bcrRPCwdFWPqtE8ntFAC7+5NQwoprs2DPMp03isEYq6ukwTuql0yc419oeEa
DVNObBQu3lKLOmYlBnww8YzgRwb6tOK41UqjF/9ezLUc1qje6xXKMuYt5iNW
rw14y2m38fjk7DaVMnpAx2ZFQQ7Rqvj37pIdwAqCBkDUNe8JtLDU6hb2YRvU
xolB3rVZzONA2yFJ1xka3HRmBbtn+KQCXjAwsb9xOHi5nvjkF6GdQZ4hTgyk
ypQSnDja8f1AQ39aKabaejOnV0Gp634N0B5J5JdHyMYhW2WcEn/CrlOPeUwp
yyYNqB17GNuR9NGUciu4s98GCAovZttQpy5JI4M7RVb/SbQ1Qmp8DtNNFeeJ
cCHx9eYzxtC6fbGBPXfMUin90RA/3IpzdB98PsSJFEr+DVUdbayNlrJimG8c
IG5EKQs3vx+MtlBXZoi9834x7TpB76q9IaKuq6SRSXGZC88T45/miqrrp8u+
aVXAYQ329PVKWIPpXI5l50eXiXxr/lLK9XK4+dY5zwVZJyuM8kfm3FOHTi+E
e9CD0NDUFuUIRoGdSCpNpGSoCebqMrNehPLmSnERyht7VMlsgD+DBPEnLfe8
yw0wDBEt8D/tiok6bWPHcIZ7zg8IacTFR+k0I21Wrk4vN5cSlHomFACTAN8Q
R/2lhI0S/4Q0luyF4hIVGush/H7u4+NVZfP6mlJWw14a35Z+ywg2GJFt4oyf
mT2H+O1gpMXfZ3gd1ciBpitlsBVFUt3WLhky/fHGolJRYQ45R7xmrwsgyB94
ijyvGwGuWaDPzEP5avb39oEqGnyLNuzKHhRm12KnfGgRrpbfcQ2b2vatBJhW
YIFXGubSR+bI+TGFi6lPfoFtHs6hquAG8ev/A5L69No0wc5j3rKKHRsjDJUN
kzwzYwWlwDKeFXKCn02o6RBdmxvz5pJ4lHwEcYSbvt9eE5CPS63OFixDKj27
02tcRHzewhCKufpm1+bigB3R4en0xou3DPRKQt6AurpjPU9IfnhC/yaRloom
OuquaW9+EvQNt90n9mPE7JBt1dPtmfJJ+n2Yytfbim95qZ1Mi5rqOjwfDHtt
teTpN6Hp7BmKsvfoq7JZTwvBfoaUUfmFYtcHp7UZiLJ27+fi8XFaN84Y/l3o
PARFT/3kdwdgPx7T6PljcebXBoVmoPkyolUD/KWPaaSRJjjd4jM2Szn7Wpzy
uHys82MXO6uRiZm+tECndfiMxOAuzMVcHEOfIsCf6TaMybBmnlrGjW3arYq2
gfytp4Bu2L3T1cWEhvjDA4ZWcWVTQ4vSsEFoQDqdbwxNDb5bbxhAjcJ5susk
arfpH/ndIpI3hb3/D/rBP/LQ1LU89H3jOij0lsa2cJnb+4Bxr48g84gGPiB1
XHh9VyL3DoRnRtFgq+IXfTYYxdgysYQjTi8jIeZSdcC4fpOY72EJ5JfBLgiv
+8cp2u8mjKdW3+UfSRr6yDX8l61XGvu7a+ccZ+TDu8NgQ+cs/iJnexZOYC7v
PGU3XrBr8uggIWwk7xkKWgS+G9zgA+VoiM4NNGg2JszhtVvg8M8bFaBVWY6S
wdq9ANqSr3o0SNDkDbIHXbvoFwnRwaVIIZieR5b2Vm/1r/8teGfIkwDKLz9K
IiXt3InUc4bFDYeY5cc3ymC5os4axSos+vGZ/qOfuvOBNC4w726lz5DlerFg
O4KhnEZLZqxqJKAI+1DFCJosFd/JZ69+84DBKJINytwScAWxqQ/KQsGd6lKF
k3s1mRmz0zvNU+1Qr/72nNgCjQ9RsXq5JzmqnOXMdB11EED/J0K5hf4eAgWS
zyMp7VLKMtWJ6Kbf+coDvtkDEmnGPFqQeuRIHw4j0tYmscf4EmXf0TaKRgxh
MSnVzZhZp5mXHj9+eV6ATFesOc5H8xwlrOJnLwJQb6sOVxtWNrIrDYZ/bypJ
tHDJs+sLnjhQTydbckXh+07sejY5DS5gLR2gEzh9RnXUxkXRUqrcTj0ESgMS
mMjHQuAglXLsXkC3vu0uTfiWcAAsPrmp9UwtN3FZSdRxNZ8GJohv0kcVLqmx
oDwEoNwbsQnD4CCIEghOHH9W/V4G4LvCYqYH3DTVLCp0qyhvX5cqtN8DobYJ
Nm1WFWFq4ROf4s6CMNQESZdiIJrf9j/No7QOedKkmF6vf3FRcTJNLc9Cexah
UI2GkP15JR35cOCSNZ7La+dmhEOYnFy5OxUK4rO3mJk9LO2/m8/l8SPejDKg
Toe0r/sDd+IJhIshH3N+dB0713UtIeNw512Gy/tWQoG3ey5mfBtkGIBUA/j5
rY0LF7o4AmGwDgjHjTHBXVHUopIBa8teS39VnmMmwKBwo2gC7+Bsd3rXmVMh
VCbOcmkn02HHilwAzon8Lg7AiyiSyOGo8sM3oq8kc9YI6cqzZWHWCJRLzTb8
wXvVgsph+giqhSnETBu1sZWf9UrijBOuFxB5bR6op+XmJjCk+Wvp59Mxuuy6
CJvXEjBSNd71nUd1YN4nB6Oi/7DXvj8TvRuoH2wnY2dMry5+PAvN/tq6rNOW
ukViAxW0POCWglUxEM9qM31FD0gdKrCOySG7BL+WKf8PQVdWtjRXJfoECJXg
sE7Y1ut+uprCzATsE9jgxj7e8gxkxAp5RH1FDmZUr7xjGM5oErSxjBV9+k/4
sLRY6MzGCR1YI4IHqIWflItNwWnjsTy18VfzL5ppfAujCInDABHwK67OEkQ8
+jTBL/ZpWJFoXCtja8zFB8nBwCWshrMoDhF0bQFaXKeAH+Xfgo5Zk/NiXfxl
TUZvsyE74FzKC62Kh7eLkjJyCedrmEDobTcRZUhTmNGu5sbU0Anc1QjhyiTZ
yptdWmOkAn820OKLgPg1O8RpXlYekg64ytpIxEoIMDpHGUdaiDV+Ul4NtGM2
KEqtGX43MHIM54GvJrY1Cj1+5kdgWR+7I6pf1r/HGaKPjkW/fgJVaG119Rem
MtZ4lLV5hQEja4lEK6xACXhiQnxs7Q5t2lPFiTKTg2H2p+/6Z6pvAjSB/FaL
p6JXRYBX4twIPvNt+jmyit35bjsTxORaXq0KjigiaQUg7PZf/DtvnBoB5W24
ZEU1VJWoFr/MuZ8ef9WplwpNhN0OPigVWbx3FsPS29PGzoUTxz3Euwg0jl3O
h46hWFZZljvaE56spV8KLteqVvoEVWghy3/aIC2mT3sHj59gXnB72lkvK4CA
kseCYa9cXhOjvj4RYdeVpbvVZwJQgOkJZ4MYyGTeC4miUOp9fgR3RAQlLTsY
z1g8tSvDoFRn3s1rHlg06WLllLJ52f2nYv+zMdWAC/pC0Bl3o/RzNzCj6L8f
KwAGxA/Ursd7xMTTvoAeJMF/e/S8uDtzwY9Dj09f1zyspaH96NYHoO8XSAsw
Q4wNteFr4Ugr0x9cOzPbsDKimCvvtciJ5sAPW7wv0N+h5nGhqk6N6/BgWnBa
wJ+kKv3n2HyKw7aH4GM/XC9ouvU9vfMbomHqGVyv83InxEGoI02bNyt7vkcJ
stmEQnFaRb3tDf9YgYbDhOeT26ppBQMmEoMz2/oo784bUalNsVkJGmqW0LLb
I5Zcy1u8YYvpgdy5Pw0htVbo0kAYk2Wysmw0bwMF6mwQfYRtHicWfs6QbK9O
Ad2JKrNjFM9hEHG7i6BizPcCsW0PlixK2j2NDxpoBm1tKeUULpUrarbbu2ri
GELDMYwKUgtRZ9h/uCIMjqAIQISuD6jNJSWvdsrHmjK9+5Goxv+Yme6Drwke
m5BDUbUYNzOoV14q0fQvreREaoS5nG0lmWX8NSCVsnffP+lKMFNyn5B1IJVW
Ow0Q4SW4A0DFpcPvKgCxRjk6ze7776fS17G3EbLPNs7Kzj4gbnssHyWhV+Wm
30Gh2FCgIQVhxdPHoJlezcZjs8/UldJEzPZvn9Tf1JaFcfj8ofItLCSQqYDI
7P3rwshs9VYB6yQZ8DJG2De5JqSmZloG/OwvL5K8VAeNA6eSv68dM/anDpKw
BOavmVzpTVbBGUg5sUCaV7Bk0FNQl7IU67rh2Kd8/chwLhM6/oFfUZRhQ5ZY
pEGHyT7TZB3NYEYIsb4xyzwQRqf8ylBfiRTj1AFMxdbagSfcHakGgbDKx5+K
7IVau9RNeIYX4QPG85csX+mXyaMkHvJuy9Gzgv6fYb9h8+6GQpFvAyezzFGY
Wvfprm4z4v1xA+WQslnRmEay+VB0WJjjDJZQQNYyOLAr8NWrHtDS2dW3deT5
T5zTWhjT654kZdAvuOtDo/rn14p9johS/hyxRlpvdEeI9klGegxqDKUtKb/x
+KguKEhaYGZC4lMC17sJ2jtD/OGmVTiLf/0/f3yIECnOxl1l6EePmKWRrlgp
uIQ9ZPmb62eVgVGqDGwqHEcHyvkV8lJMK/bKTeNzHLf4E0XLTV+Y0uS1rz9d
F3NbEmnVQubZJqK1/oOnnMopBe4ePD4Z8Uvcu+YsumuYB7MvFjapqcSVi6kL
XxqalJQ2uaKfXNmhBR5UcENh5w7SM0xerfnsZYtQlvzIzIBo+lBpTwqFbx75
KBj6wPc60pCyg4TKg+uk9TIEIpuR6Lgg5DytCc3/l1kgRZM99Gxh3deCBg9f
Ca/S2bmMHGzDr2qkkDw7PouOHVNfY7w5x//BP7wlqc0qT0S/1n0MZOytc+z+
vlDfLTMeNv8JsMbzdxn9p/PZTZakIp2Ci8GEttobh+s7ytFwsCj2/ebZHKNW
Cvl8IFvjUThgs0KcKlA92wbyyqTNCj3HRGVq1Zv1Z6Z0N38+Ls0HwSV4Czuj
YI5AVkFp7J+Hd/uMOzVEd8cq5vjpT7WE6dSOXAynrzMljBjt8COlthIERYX2
l1tI+9taLclp6jhch43BBaTdbf3avo9OmSuQysWjgQMakgaR+2ibjx0rkClp
+OPQSbpNkVGKMavOg/16CVSO9eBIPe+qR+Sj9oJAqyDgGXT0SUcUtVwl7kqi
bkZChesUDiMXVD483Ov0xtUrci2k+3QG+aP9w5F/g31ry88ZtL1h8Dggtwz9
lC3AIa00rEmltwrHO4mUlgyP7fYROnYTJgMubvi7gQW7yeobh00wD/SU/5bh
iwBvKhfUjwo97ek8aLDGwzQvdIm3tiwIHVPTKyOdjt/GiEfrDo+q/AGC10Ix
Xv9R9L7lEwxh9tDojQmwWR+7Qo4jyA3blswOniTEhv4drqRMHydHZzmd9XlS
K0aZIZsiA+Pua5lBGDU5CI2FYOOpdt07B9sCMlzHPKzFydZ89g8ARKULPC6L
kAUEnzuqClmpG4JdQ+RUvg3z1DvvryuCh+Bw26cD4JEFYOJfShZjRjmgusGz
rFobZCyMmX3l51sg0FLRgrz0h7mxnD+/Vv4WrFAwvCjPem1BDSe+pSRByfn5
wKnBB07cLeJEYuzfdzMhnYBUodJGZTHtzXYNvnM11Td4J8yjwB1hZT3cvW5n
vBnVYp4wo6Y4BsN2ouyVIivsQpKNB3P6+ct9pXP4ucc4ZVjbsEwCIedLg9a4
G98EmIC6Oc5GauqTqOzldXtH2nhK27wUQi8ZVf5PTm1rL8MnpoT/OABB2CfY
krmlBowGjX/jQuWlQrb6HENEtW10laYlWopHhdu3y04vm5GLIdvd2Yq6UZTs
oX715JNdC8Ebk+t+LwFYTyzJOuO5EsSuY7wL8tv9KOSxV+r8g9chckg5TVTV
L5GmGxquoBvTYH6mjEWc72h/IiSxjsyh+qOdZb/EUhLsq2/iaTh4qEQttTf3
W0NrkaPEnJkOKuqoXsCgO/boILXV6iLIVEvST1q6VQJ9vMmsAKIShC/V5/Y1
q2f8xA1w3u+m7Nl0xMa+/y+Dt3UrD6l76NUdTqc1pXgys3eiQSkX2sY6404Z
0I7+HKmYNF6OWow0M2wd56cxOJTLxONjT1GyI2/r6EZvSNozjZ0vskk7fezU
fHsj3bFgQo6ktECpnN98dm6r2Mo+R5KX3q3DPGk869xpgBnnBDalEoaDgLtr
3WvfS4o+/OTjHvNCEKXXypzm9BLbrI/KXWhEG2xvp5e0PxPQp0bPEWR7NvJI
oY1zCIJ7YKHwpstlLvY7Gjc7mOcXAo2sJonBOgFNG13SsuvhvzCf3Q10MfRp
pYgJeSH34A9loP6WF9/Uv3SZ/B33au9CLTXk3KsJPpgXarEsFwPMtXs3tvG/
tQhZmo29RmqnUZpAD4nxs3/GDR0Di4neQWWOfFk6xfAUobclH4KWUsHsiE8R
qc3GE7SQtWo00J8JvY4kw4q69n+RI3sSp4tClBP/dJhUKRyFqcA1ATfvW9tA
2OQPYqdz1SA/kNhHx7P/dqgDv0SifG3jk+NUE+Ci2S28bbSlDtf/R/LLO+MX
k4/pRXcztLr5+69QOBGrrxmvYD54x1jvifWm7hMVrHqWMEq+FPrzqqZ2SIt+
HJwaekEFYkgA3ajGNLGePENL1dLRYrjb+0NBEcsCoGMH5/MH/Fucvm8xLDvU
UVrpaMrUVZu9uLVKCM6tDbAKoY321a2L7eAD6qLoyryPyihkWWoqjQYz7qio
7RY3sPbTfY7i41gPCqFPJsoTIOLymptYkICjaPMp3LKIxdWu8hMTMfbg0c7Q
HBimxqSBjkfID6ETI2gXMPaIqlmfL48kehdCGI4iFP+tfd8l5V/fvxY7HRaw
t6oYNibROuMCGHVR2InxuZgtG2g+VPgNtDdunufnadDrJzfGQi/XDxprnSbi
vFkMJjWUc3debNokvxJX7ZfLrZSFRoqkti3Y43LrheT1btW8FuMbFG+OffqF
+z4Obi/VSlfDyc6Q5sAd3EcXoQQVvUbQ/IeNReq4wR144jOu2QWK8R9zGvUj
OhtweyqncsONSX99qmEmv/gsIRQDe3zBr25qVsk2u9mLtNDdKgLuXSUFMpkN
eMp4NxVMNL1QVGFN3FoxJXPFzOmZzJzBaMxBnyBc+lcBY+NFIfYHzf/meWx4
rIoCIW6oF1RaUsV5DNVPCNbmHRwPaOx98/L3naaLWCZPlVyrQtHUQkIT7HXI
Ke0FnNVcILacGBY3GT91o1+ZXC7VelpY0PmJOzAzg4lid7VILh59d/4BHWhX
O+rpZ4fDHUuKzE8gm0VUPyAu8KfaBBKG1GK4W6iG/Cv3BmAZrsxkaIR/X/2I
cqSFNTFr5sFPMUpGjD8SgC4l8SZtyYdjE16MNeacXKD/9ZesYU2H3qdY3Du7
uoq/5zAeajwcllemeBYJQahVtUTYIYADBkdShACpSzh+bnZaBatDtNMYSr4e
zhlwIr0eRDeACBAeupD9GbQXIgunn0N+NvHp1rGwVOHRi1oJukpUSsJAxCk+
ng+otoFbljDyHcjhQSZvvBR2bA+zhi3cUMifIwPTf+jzAxxJt0Vr2y3boy95
yQMWKq/Sai4XFvsq/J5gVtoVVEJvF0fX1X2+prEZOscLA8ycdoPHoPdbul07
fFjxHlEY3mjvgRryhspnVLqKllx7aB9PE+BI9Ve4RYNB6I61qzuq4xD0mIed
HC4N2YiW1/YiTCbWyLEgXHcvjNKkF+gK6lQMSaAc939wXBhLL6aN2X+Vuy8/
plR9jtg2Xo83c/JJpjsRr99rI5UFs7kiBZhkm1saTGR4xgvReE3GVreUzYw0
Zs3OhIT3vzMpqCOC/ofpeLZnf5wOXQ9M5nfInHmUXZOJ3vV9nsCO5eLIeVbe
itpfma+k9FKAQF+/n56iOuJFUn+uEdrWsvf3ViZ5Ur/1EqPepGSsuzbuEqE9
bzlzOVk4SuRTuN8b669TsZ5Pn4q0JfdrWZginNcw7vGklDLwaF6F2e9CWGdp
4lMUmCBmyfUnZ9PXm4SNKYfBTU60DRYlETQmu4LljQXn9X2CAFVvpSRWa7Or
STBdjLI6C73n5fDYaRU8sz3xH9FdEZzT1Y1Nfy9lzBZ4IALl/IHSOQGSvDMe
wcDIvIjSbpQXpaHQSYZ0hW6Uww8wP+CHYRhROfPzollmp4wtVqWw052xn9vZ
jX83qDvhDUZDM8ueC+LwE0zzsn0PKr3OduNzPRrsS9MHoNUnf5px1+BxqRcy
FbQmIjiRIqdVrS0YB+pEa1lqtydEOxGMDxVEMDN/q5UnsRNz/exQ/VtZT482
fI/UjcmwVInTxPMq8ZD057oQTdvdFJmksd9+AK0aH0/fgzSpLghlCGvvaZfS
meltk/bubu5FDEMdKsYLZrilJDhalROSzwTN1STZ6CHwBnZxEqBZ8yAa6Ulh
cvtuegnB1hol+JYFQ9vTxggJftbVpVb04FYUNDvEEVIUyjMd7JX/wbDKdWUu
U8Lk7BEa6BvvTIdOVaXK/s30o9K4EAcRxFMkndIL70Ky2AJUHa1vPyNMXia5
8SGNNsmhV2AUSaJas3fLEBAKyBppmJp1EqqjrNU/T+g66UKGM6kQKsblMrj6
dsso7t/NYxjhnB4AgxqJxdN0o/OpR0ZjSVUgUeEtBMoHdsrg2pwfGE0DGbjB
/8i7pCigpRJTHWNUgir7sLu5Hwlfmb+MOPBqzAYwLO9BxfyhUPPubllMnakr
Yj131TGZU7dB2g2K+WAEc+EX5GG+wJy/miHcwAP4KZWESJAjNC/J7LZMZ9tv
Gyb6ih6eqxiC9oYsXpiKI4R+FC5XI67Dv3WhHMMMnOPDUWZ6HUN2kBosYYb6
n5l6LMDIQ5QkR3roWur4J2IV6du3va5qxOliSlA9f7eghucNhTT3HPwm160J
4BJP8uvvGHvK//0VWqVQ2W+wfn9JcHaKC4i5mbfoHXX4+GA1prfDGt4muchu
Rt38AYGxRdZNi5+2Jz9FbEvJbe/p1YPEtEHa+WQqd3yJ4ZnZfHzUaPgRDqoC
Q6yc6KmKW1D12JZHlpJ6q5AZ5ubO8HJcmMOFXTZgyy0rItWmriXEpXnGPkwV
BEVFklr5UrRvJXuG+C9Z2unclU6uxhIWGdY+lFgVMsq2Nnyy7czEqOjYcmuw
WyMR/ulgQsu4ZGUDI7Fct1wk2gkB4wgGapjrveYfIiA0W7Ohq6tcGUTp87lf
213t5HIZSVeDxc121S5XEWjWTMHFCj7KrkFQXBuGEkQ9zlguaZ0qAj+zRfVZ
w0+JvNGNIFaizIW50m+v4BfSVpQNgJ03c7XpOlWrdZKqCUK/vplg5le+mtb/
ozaxx8viDzADnt707Ss0aBo2O0pZq9KzYRxCJNF0Sszv4AxN79/kjgzg+tp/
ThsXCOvRk0MVit8jNPL3rxrqIO9d+UgV0nH6hLcFzgaYcbb3i/6eM3tTqGjl
z5sQmBtFQjrxTawBBJ1ko6wHmGeTH0ZKJlnZUb+Uw6ABB8hxGDMON0BcrDoq
dNY7QOH+uksKlBtKcbuEf0upJxl0FE7vo02BJpXsnLFMLB206MV21d4kXrWQ
hz0mwkU8J54o4+hDze0G9YS1hjWd7TH5iPG3WAsAdZrxLeTdwmTof6ObScpA
H+SwsijHHnTuwWaPBLzb2vhdxTw6Mu1ASbVSUT+QJF0aqcj/aEYKoynbpRpW
l4xYoiYDQycKvYP0z6J1ThJtQx3iayc6d52BuOtz5MNnbO/MfuF/QWCJdtf3
AmIus1i4DM09ntW3kcuXLBgWNvqQ4iN6hMSr5iTlh7MxPeFVZdKwYmYOCVAT
CZNATJZKLkjjYOysKuWr3/q09QYXS/PuSdv51zNDrHVFz5bunSoY/QZ4PolB
RdHZYYfKNPkQI4CrcmQaEddxfvmCIF25KQ/yq0BiUvOH3Zx3GBLj/ttnjXT9
mgZMih0XE7gZvP444ikUp01J2xc39KxxuqfOhAvAU/c+QhWWVyD5KY6/eskU
LbTy374HsC6sUA0F1AzGNyjxIlfAJ8ihBxu5kDyJWs+5gk7b3MQGVGaZ9q+7
TMbI80Ky1JonxJo0or740LXPi6VcZIcO628rqDH5RLwyUkgxSX8jpiumas55
HqU+gzpLtm3rcZ6N6VZu7xKAeOrAZLlyjl8Pz02jCJH5W73ycBZhyw8fk8nb
GvzojTIgcLhwavHWKPFguhwD+6PMU/4iQOdGxD5l0FvdxHSkGysIWJrmObg5
NUxY56ZdFTnbZXLc1GXzRGC+qnhLMrp5XBQZHBttM3ev9WUc38Ovb09WMddv
uUGxlXh6ZqH07vnQ1rhfDmFb+8vuqVcVfZIN4OP2g+Cit9CiE9D3QPpbTYmF
wYtcBINvbm5qbuluGHbHWWPDmZZkgNYGJ0cxdyHZex6qA1WIJwdBAd31w2UP
t+8xVc0e+oCYaMFmE/EYkg4V2PMeNpKDKxNJNLnCQBED/nW2T2zFRoNj4Crg
XG/iH13TM/tRhDWqEvjJatWcoZKbKyQRY0FzuYmc7P0G3/R1RbAma/bjjqk5
UybO3AFKGeBkeS9bZN2GodEaREG+tz6/GEswY8Z8BZdWkZd1MHotcqlUGp7n
GJqLmguD/kAw+t1gIwUOKCtFBnS7GBJsJXa7L9HgSJjmBDP7cgo4AosJbhUb
KW5cDvCDvJyZVHGNgC8XRad+l8kSoPlahyppYKxZ4R9opQw4Yu8OBSXUWyll
nWUR4ufX9WqLPEFGGYatT1Dlw/bDY41Uh8ZN3sfrOaRFEq2BeFFkd9gK3mq9
rEsT0TUBXzAJZPTseeJeEkb/Ox2rXY4jcrE/HTTs1fNxFuQLEAz13SUn8GhE
y2dXzLJSb7MNcbU3uKxXoKPYpe08z1Mcu4SfAoyHPfTrploXm/9m04YumTwk
UN4cgx2KLZMkfevhmJuiBl1N45/RZLnCGDWesbarHtviLzG5XgBruiVc8Az2
TiOjJVN7219E7hF7WtjOKtFWBmHVGuNQvjiaghn6h4uHc7um8v6FTws1PKud
ZTtpy4Sw0ei88dlSdKKMmXQi2V6zatMOauHGnip2wUKLqck8NwlPIkUJcQjj
5Yp0qly7pIoHZ5DDKKwFDHY8TeHidwZojb0GAU3VbyxEBdPLD5etdbikFxqi
2Igmp6zp3P7gpGMntpVkU38TXz4lQ+BuP3XrTv6/6/sndGD1edF3yLs3MMeX
Kp9GyLj/cYH0yqyLJxXA+VUZCYb5RWDautlrxQQjjrbqmPNKAtOZ0cRZGqWO
TBn4pESl8A7w08+pzqdgb1cuQQHdR2i/EjhBye0qXBNsKp+YyjTJNRTvtKef
zEG9t0JhB/YRy2/kH3L+eOgrCjJ01ie5zsbCAqF6Fk4JVtYOJwhRKiOUhijz
czT+1gXyOPuAt+gjvaVTGlZZNREuPDOE395WAFJ7gu6G/8uTZoD9G1cgJiF3
MA3+yM09kQqRuzVp8NFnu+AVsTuSLqanRCyaLdowdhhBnuzK/tJIy/R6gc8i
kyFWeiZff1VrDJKqMKrWp0+IInwLm6MmILXmTydQBK9yzY656sItOo99hVPk
Sv1/Wzg30kPxvmX5GhvaEybKg8XA0pnJJJqUd38tqH/jtlouaisUmWPSpjF4
1VQgLwsWD1/iONPGJmuC/xs7dZabSb9CY4sFYBFul0sI+0swNhyy5htpItRU
Rwh9EGce+Uyp/6XD9h0ltd4XNOlDI32vplcLYhWqaFtIWVqnuuYxp69M75Fv
YIZmgX6wB4pKNOwnnn2ylU+n62442isN0Hwat9tIKI4M1nmigxA1OEssBwOQ
/YY9xUJJbXiyjuBtyygJqfGn4PhCsPj5obnlhI0Y8/y5SZLn4/6vuD0SnUu2
RTghpEHhWMfqubXgx23/UhTaEu1eQ8XTSbqreljs6DHbd/md8/N8DxP2jePG
JKDvlX/rvdZ2pLT8OHX4Qz1uuF3lRFI4UOsOeHJFqQlYfIBJe8hL+euYWNEx
xtAN4W5EQcgcSrQqIR0FjhmQBZ7I4onWYvSykezRU/kn0MHDV7F7dOcbhbA/
buH29zLsnWGZc9V20xtEx5qq4ar/pMLKoD9J3T5zpJeQq1p6EhnyyXDCjA53
7oCx10pdOUDoq4EAY3bbWXNOhpOa1K617VRn7zYBS1ak1eiDTJlKI72677p1
u4eCgbFFfgYGO+wo46BoNfohCleVViA0LoMsJHigKBTa75fTjJbTUVB2CEhW
2biwH4texMB82N1PL+GAAnc9obcAQOUSixV1kYt6hmdJohSEBLY51i8qnZ59
co2XWNQGQnuv0U1lMHJddgBjwzdcGOrp+KnF1pULxqc3E5f5ZtJpTcr2fvnZ
X4qlX4ljKFkJqe5G5hM/bE8y3o+BEZWvD5mfD/JWVRolj3p3WFV8Y9WAt0Yo
Fxmw2mew56z/zfebX2YtsU24CkFty2lbXHuSuajNiwvE2ooBNk5zTHQ/zrV4
e8URZsad1+v2VTAA0LCved10J0fBSuKd6TZnW8Uu0tTkIlF3v/PDEKDhjkZn
bnWkxjZm84VkaxDncK9gjvwBFB6TCFEoHmz1mEf5+bdisDPHDjGPsKR0gjCg
AUyeaWvvzVOnJUySR6MeSoAw236PooTp3iXwYqSfU88cYMKLzJOLCOfD++tY
rny9sQd1XS7U0lmmDZxdf9h6bsgcaA+QxsKazSg2wAKScEMGTymQHdRCWpCa
Y5QLeO3wnv74afnDP/sIdiH1Loos6eNwd5jlovMG3D0NZDIkKNkKHkBS1oSF
RoJGf9obqo3RfmMFX5UjI14oCMPjYkU56MTq0ohQeUEudY558H+OFejogYeE
7G7Y06erh0FUjA/ImBW646fOKYjPUSh8Ii4U3C4B81luXW9z2c47dCsinHn9
o/iPjLm+/NHcn5+lCiVk8PoBc//mGSGHmeIxTHl/ko8WG099mVNgvfsdUW/y
kbiA44m/apkYFnjHjOg2RQSOY6JBHSRS4U4YUgrHWfxveyjIeBvl7CZ3fCXP
cJoj4kRUahu9rVYYH/DfkEy+aHO83taim1kzCCZwmPIXLY978QDZPrTpi6Gv
5xQ1GFcwJSC9oycPB4VzepEn9UNmR4XQJfuGNscuzdIHSS+DUo2dRlkd2afw
F6/LvjfgODbuWpLLNobQk8fa1i1tiEZVP34ozGIyh59WaDTqL2OtAa9oWPlv
7D7xiGQ+iz4m5DHzYz9Wnx2DGAr4TynZz6sXqAqNTSLBQ9kem2fZCKIqNK26
wDtisqCLxcfOa3IqJrPcs6wq2lT3vFXm0dHJwKWH3WbVxEfEijwtmW6LM3ig
lAH0gbyvmNneSlevGxO/r28f7j4FVHoOMSm7kThr1kKIDxVlUL824j6w6cjg
pPTfOnIq9fliUGFENOd3DjykBV+crE5bGcLn7fmNzUcdmOsUnx4Ziyen1ssZ
DZDwc/WOA2PMZTcO9zdOiqqnbYNyeSRx333TY5map8dYbSXgPmcFAQ84Guj+
SIXiTR7mQcwIvd134whzKWJ1Fc9chZF90k5v2yikVBU3TYChwG8UKzFDcdz9
caALbEvYHflXYJVs8SVkvAMaGUUYeHu/QdIhvsqGZdw4g7lVUS/DJVUjp3kb
GeOB33do1MFpd46yutTZJ6Q4Orh2xx3YA6mHLr/sdI7bzh4GKhodvqnb4jCS
rpUwiUUMLCaaJCO5NvUVyGCkZWCsa07zlBZ2idlgKFAJGUsL6kLGvdH4z0+P
cOB6gcOpyGZMNSlHxoZ2WRtNNlHr2lLPsGqe0mK7jP5eJy3rW5K91m+FljJ/
YJFg562CIf11sF+A8sdo1w6Jnmf/GNcsa/V3pF9neWPKNIMwwVWFHvNqSf/4
/MoYUU/9cXb6ch/pMYEBM5+jaxj8hh1YOKk8JuhTvRkrjWHNh3nl4tp+pcu1
b8cPRXyAexGXpFYBtNoxwmLEye8JkmloHh9H5XEF8yD1oorMJXamXV8TGDCC
sv9jTS3Ctn2Pjh4PWBvPo1VQp5c6wH+u0MTdpWz4hPy9zGzC85Eld4a6+YPu
2pv3QlM6kIYJxnl3dVTaZLn5j2thQKoK1uh3VrQzYsJkrYUsAs+4Zjf8sDef
y+7CDpFkf7pdv1oSyfqv0L+VDorHllkpp56C8IRXrZDPmbv6kQsIYY8TigAj
QOrYGluR0XXNoCsidmyiVgmj5C2LhTBniAPbXBTrzxH556Qb1H4kRz+P01xx
NPJgrjAVBnesyBej1yDesNgffEctu0fdEEYexGqQXXQabSRugGL0DjCRUAKw
lKWDH3cT0LNajJfHy9bOb0tjqi56vtMUoCX6C1S+4XzW1/Ydzz2TIkPO4DNM
W+SZ89pjF/hZ8adFvKiTSU6sn9JtcFUWDf2aBYVk0OPA6XDseyNzuNEU/YJh
ScdzpfX8/YfJWretApBh1QPHU/B7IWm3bBDNw0HmuCWucR2Hzg3jdkxTbith
o3VrBHNU6hWzak1J65roz3UW+WMLTohwIIU4FeVsjChe9rcQcLHxFOWaVTs3
DaAXcHC+SeyJwsQfgnjkyWln2V5/dTEdlbWUaBETaVauiEojy5PaDYA9R8HX
Pe9AXLf8Lqq+OhlEVT7j2lmZPjW0hme3VRYsQubwAckrrebE3J/kgyRo+wdB
oPsfYnsbALN0PnJm7WXP8/hMRvm7mZqIyc3T/HuK2/iTK5IpPgwlew3ewkd7
LWTmPEQq9P3n4k0DVhJSWGAqZN8WzmlcB39Le0SeT0LCBqABsmC8uhQQBzoB
3+eWopM5WvQtHP7j8Ay0LF2p0xn815vbi1bF8TZn0bkYXAzZrSCUaz3PUePI
oHCnROygyL1vup6Bc12ihrzK/zRnkhp8fuBMxB1ks0HmXrn+2e3x5K5b4cL+
UJAN9KFDQg70PjhKid1/gqkrNV8oKUM+Vti2tQUg6ZgoEE6K14XVUHySQKMS
dE/CeyRMW5Z1cVKDNEO6mBhxNg42V09AJzPO9xHuiS2vLolSDKBcugzVDpcT
Ok8LahEkQq1fHrP0LliAjDwapr3DFTWuuyqqyLG5M4tC6VavE/ZHpegoW9V1
UqZ5frJ57d3fOMQNhUVO3FphBefmd4pDYvmhZSapWKWhLpM004a9HM8W8c72
6FTuJFx+9bt1077qO1j9oPK80tCta4OzWRY0MyUyImbSuGsifXWc9WqDO07e
pF7Hto7c4QVPrgnUwry3WJg2CNTB5kw934a3xh79ZATX6H2tH9ctvVJ1eVJ7
tOqD/XX0yakzWgay0cjG2/2HSm/gCAQm9gWkaUUF+cmqWIFsAxXTn3Tyz+65
l2ZtLQl0yrKCFSNL/ya4R0AiMiydE5nvEY9mNb3jlpZz3Yhx5FahMyRqpyNc
Ft6L3PVWOd0RYZCTeXRcxSaVD2vqAyX/n8rQXIYl9gCs2/jFCjeU4aIhLoRI
5th3SyWbKl8uFhmVFH9n+8YPnPf6bPVANoawTZgy9CpKNfl2ih6H9sCcmIK4
1hOfacS03l9xej5PRrYabKYLmMCDLSFB16IehS2SEBR8a44kFqZnFsoGO3Yl
H+OCbmNQQuCJ3Txudv2a05sduJl9xdA/628MF8JMVMXTLBJrJ2U0VPPatnTb
kG/4ovrnbA1bj5vB8FgLC9Ypxji8xznz3Hzl+yJ1oxopp7nOwKI1OV/5FXMo
Bjf/uq38Efsjf2ZAOdH9NA60wzx+f3mfVHVdqDa7+7LVLp2o3x40CfkcCLOT
F9FZ5MJaInrDJD2Bm19bBT7qrfJ7t97/Yokb3+rmdysSSOdsXsVjbPoKZhuV
5TLQ+I8POYmq49AocxAB8wx7OgkCri8+EZkPUpkvSUuzP/9E7jaOuR4+TP5c
l54WZPyz3xcUGoL5al1E4V2LVSp98/SDjzMfDkYQ5D8HApzDn3/Qpakmx4dk
wCcC6vqwPaFwmhFX0Balyao1YazcmVAsN/cVd+FUVj5kFQxCKsTKo+u0Spib
I7khnUbVYCbrZHVXUWVkAJDgES5pg3qAObLEESP6boRnspUz06Ymd2/n8S4d
pmwIywmjgA+JUB5WaHuYOJ1LJa23je61540J8rDyPVJpdJuReD+4l9G5hl63
EzVSfFtOnwSds3dRDcqThIyfynlF+aJXn87TH5fWcxefOcv2NGQVh4ddb4us
9pQQd9YsQnrXs+mDbjybp3t58d6PCkI4K93nGPJzNfBycQcvXpRFta10mFhb
E8W+yHYvIHIsMfQXPM6YWwqvqMazivEOegDzX54NXgt+OZTjk9Zw8kglX5ts
FC0+2QplYxwQEMQa+BdF8EpKHvktINujKiaF9unvowgI4nUA91CTCVoQ01s1
yZD0Kv+7QGrEwSP3TBw+b8mEBRE7c2mRTramvsU1TeaLyBiIVdkuUQYNczL8
GxGP8RsAIHzSKRVwj38IK+YZUt451898ogLPrEIh9K9+XFHHhFZTK8U0+AFT
XTh+JCXm3dh88c354BQwtkuimo0OMq/TJdMSnYtyg851UYi2pBan+KR71qa8
PkNdmRPRQpUtzTpi1nevpI17zLAYHLDerz6/LzQlfDCP72GLegm8/9GmHDg8
8b0eF++lKF4mJRBi8k/n6TJJGoOFLD4I9b0/9Z9RyWNRldyC0L0EBxkBuHgM
vcLSNWV5l6EMu6ZS+5P2dwxewLq9zDBlGwr92e5sKzuN+f5KB7QKcB8kQ2I5
ubOh9QTZ6gSdpY9Lm+1IdqoSnvgjMtgM/TuRl9c1N6Im9T981zhOfUEvARRO
uh3Z9luH2xlrRu+2YVo+lrUZng+NMmlQKZ7k9TNtwJuVfIi1ZocNOXXKiIKZ
o21b2uJTxUn9d7/v2FqlT1fTsw/9uRtwVP60dwXA36NQV/lcIgxgIywj3q5e
4ROyTvXPJKnoAqJ+Exhz8Yl0D2bcBEXaictdcZ7dNLmxTjS/AOmZ7y76HThj
GpGnoOR0+XOdNydzjxKEUEFlkvZmz1QAwUJnxhnXKrOUI4GYUoojrHX8k4Mu
9T3PmFeWMrw0PeTsUIo3Yu6vPAmllmNPu0DPxmzVfRWSsoaSjOW07dmerg+g
x1QgAVShjaSQ+y6vJu5PrHJgMz7vPZudzqQjGGHKOC/DZof5MD98ZFEZRnHi
k+DQ+0RIxzN4kheVu5sBNvaDVNiP89LCD3E0M5b0n5hlKOkST5TgaYVUEnQE
5uQuzoJPVJO9tjPUC6wPdTu4rHTPtvGb8x0m91pkoxw2clufsoPqJopHMQZ9
EMR//YD2GYsSaLUeWOpBUSFR7UoaNqjcL8P735eS3WfgFurFZZX6ArLUf2eU
EEsAjNLc07WCOiuQB8PvvuyBE1HKiaYFQwcMuJolpWD6EOzCMfVAjDIwj/3r
BkJuI5K8DGG83EfXF7UzxJvRujBlh63AKONP9t5ChT4Xl4z3HPOJc9XJNSA6
rFql9fq293eZB5pZSfzN6NYmDyAjwQ7/6oqz23qlkg7Kle2+YlRHDvlny5X2
ovf/MTTvStTRMWsrMbhMJ7ZF9gh+VvGuZtk0NkYcVK+6SpCnRspqLLu5OTeH
jdpWLR7f2r9iNv1+KR7N6sVtBydWQSj9lKWbA9C1b6Wg+XXMNY8wCnbKfc1b
EPcwCi7u/hPsvABtZSncBSiI8kwocX5XkW9wNq375dsveGIdXfUDMS7mU6BR
nUk7Mwfnez9mIGiCmCV5svc/mV3NPXQ0VJar4CAn2fRLnhazEgB5roUyN1Dr
F/AhmIh+nXmqLBG70Y73MzYzzo+WkxXNxlMtPuEE/k2he2wsqd6jsGKIdfAw
VUm/ZbEEQdWVQcefGC6BGC5yPckRo+0fBWjcU8Rm+pOE+Wqu36g7ykVjJzqY
5F8ewrQXU/ObxIBNuDwvYErIRflMGSdbbBUS+N+BMRYpHhnZAcnZK8FbbvCS
EFTrC4LQ5mBXW5XYUlMKYQHWrJZKZQ201e3QqwAja4HDRnUScKRpuGWCiBJg
C17k8++CmIKWt3K8FSHc6iVqKTQ7pIolXqbnXgrkBC5gkGX7cNUCJQpNrBJk
4opYEr8dG/A0xYyA10JuuJ1tWqLUBYgPwK9SURzpY/L4M2drvQ2zUuCXXSx1
4DMO+kBxLsTI7SaNZGA2AV7fd7tpBpNHuyXHPOoeSDdhzWASQxt54GFFIoKM
VUP4f/THhKfy7TPYM4nrvLO1vB28CkZEeESmplGEx6GzpzUq5XAMxe05EYjn
GCHcmWuLQZBLU4FNYDjtG28vyriB0NP92CJ1jW9jc5d1z+RAVBTBOgh7ld6X
laxCZcsjbeEfhiEyvRDPmorJyuQ0cKNdiYFSICUQabtQKN94Sqeay1RQTEk/
Bh6IXIoIOHt2hlZruYzU9efA4ml3yaYN8PZGCfmKGR1U777yNjZDB9HuudAJ
VWMso6IwyZ5/QCG746q9ZMsTje8Vo2Kk2LnqAFh1mfcNfN0cNEw4nkCLN3Ar
B1C8BR+rW8xZXCB2WHxpnJus8iP5XAAqbQvlnsHwHQqiitqtKZFhtvzzz77h
olHMJpjeB2npkL9LdR9pHAH6KL6XQxFyKruftux9lAxwrrsihBO52mzu8AW/
dMeLaYR3BT8hoSLP+dMy1wxdISgzdNUF/EKtr7FEWYWogK/O6i5nI7gd3qzO
gXKkn1/Ye1pw4purH/jD122yWmLHQWxGadDsptdPpaCBJ3rw4Na9xeC9HjV5
+Cv03HJhn7g8P9F5fCYiGmChK/1+fVjeJBT8m/By+ab5wjKwjYzHd1hlGJny
Kh97MDftAGEQTGsBgqUonFR4blk1vr7nvcrwGHVANw2G2DQdSRBzLdfG6uzH
043sHSPdj5igFarxnotaQvjd9zE6E2S3V4OoH+onVXpfrE3tgl2sv+eZ7RB8
HKASnSR5JPckcvkNXN3SgsgX0TrlD+FL+MsWFMr57w9rBwkBnLeLt03kQkr9
go90hALf/GbcEMBQG8bfIsKkLArvlUtxCqKzIEBaI+y5sIbKhI56ittd4aJ7
lcfPEwFAVN6Lgq5Gy9qtBw9rhWo5S4TuyayRMGquLiHFTLdLkwMc3R+l7JZC
edzKEzK5yuBmkA1jDY50xY+qny2uV6D3+KHtSQQlSy08MBu+5UJ5jva2ipYG
Qpj1CG/cMejy17rKYRzWZNA22dGBXyoTz5nn7qRx7rs3ikMxiprqIIbn8W5L
tbIr6wrqzLtfBm5Cx4d956HiUr/Zd75T2blhcFjnw9X/8OrpTj5TUX/iMUGa
g6nHzvn7Q7X9UQJg6vJmSx86R69ij5bErg13i9KCO0AGv+nYJhg8PP2vhdpR
3P6Cq5R2E1EeyIFai3+4DVlh0xA1fyS/eyT6zkVPVmkrLt4SZ4iDo7DwVFTA
2sDniIPrsaekk4r5fde07YUUOkWHDOlQB9jqJlmGl7ycovW+EUsCcKDVDzF3
T6WhI3ki0joyiOMaiZI0Hz0BLB7GKyva7pzZJebmnp9qQMVhvI0yF8fuqHLc
Ym12f++2eYpBUZvFJfCXNnLUjN1YveEfZMCsZ/yOAKtBsqpd+yO2BxunLeHn
F+W/QLRjWbZWwNBqCuK5xr0TYYHTXK/GjE9rIKYK1C24BEuzUm4voTme9V/Y
2MuP4NvhTlyvsD6Cl6gBr/xY8dbRQtP3U02VMpub1+hqb4dGyfrirqrpEGSb
9uewuNBUvI+lPINcv9id+gveD1BsULlGl9EtHvArC1MNGPuE2Yn7T1ay3FeL
LGevxuBCu+S5lHXSi2CAi5KSVfv3rVntFFq5S4qkEkihnB7/LEc9VqaBpJ4t
YBndSmhbmlYxI+t25DgvEppRdgw4T+p7HF3nnjTNiT7ug4ZykTC5x+qZNqlT
tOAvU4C4LIb+c8bkEYntSICgnPlKhPvUWt4xmUjb8NjtGp/bHscxfN7vpTsi
sKn+bQSTEmAmdAB6cbCVJh6rpg7q0DhJSeSH8YFo8Ky+0k6dJy2RD95CEZJ8
4oEFU7DABWtdWPNn0tbQUMCwfdLJHs8dNmhTyhKppl34ATPlF5FGJ8Q8bLdE
/I6WsjSDNKyOxbuh3mGpQ/O0fhj+M2sRxYkeLIKWf9HGQVRDX1MzuyqMcVJS
/UF4mIcb2reeBWVgugjLd/A2oeWJlE0wtQHP2Kuwuu7bDqMV13gmMgR6xFJM
S0swMWoxOCksqinhlBNHjvsMfSj8v7GPPxmYTd92Sn34E5XvDFOrG0gjiO+n
uYahJVuoxoLdVH8vrLSgeTu21T5qdH9iA31Y2cbKGA+zQI8gfHBmCyV0BJx8
Y6bLdvl6vak0+NHqT4ZhgKE6PznZnin/94YiGRkWgrA7qy7IF8cCbtLz0FDl
uVMcJLgNOtwVN4UXjsjk45KXFhm3T7k3WM/ag5tIxiGys3qrVNjCScHvbKQ/
RnaGUtukNeLWUB6xrV6VyPavEK8Eyfoov+CsCjYtI+qmK3YrdNaKjDVh9Whm
j87dCt4FQe4ZZM2Po885/WIKIIzF/5pjLLR2/udA8uF4mMjDY2WbYT2ya5H3
JXVA+3uSLsFMi5c0VhDsETd8+Av56PL/iDabszgk/fC307XqLg8q/QW5/3yr
/IwxEH4AmONnWA2zAgKht86QNGwLZqn/o+uNclJAKbWw49cbZRGtNVs9RTij
PBmje00oobwI8WIpNxZI5+XLx1r/dkPkECNnOz8p45dvh/APZyXsiqwc532O
ZV8HztCW7lb5DEJNue/SPjQN6fn0u4o6oKPWI8owxwIquR/3zBb3NdqfbCxp
sPmp+/tse7gvmRgAuOEVgSHePhIaLz3DIjfub0d1xNjYDngXCZNfruS1X4dE
XuFbGUcsivTPyUnDprfg297Txn44c/yGyudO0k12gpN+6lnkYE7otXfkiwJ6
zRYaozqGtmUMHQm341c6HBApag6HOicObnrfxFU88g4Z+jYFPkGsnXlZmh0k
j6wBJW8b2j7AhKVjRP49BQ0Y5LIb3NH18xPxA4jqbZhHI3+vfqOOfaCThy9t
cz+qGDPP5tV0HIoSZ4gr2U6ngEaGiZiypfu+yxzb1pnzvOP6Z375AK2rOr3b
5RPLrKoOV5oScKEP3tRjZ9uw8wdKtKyEjpHQNsxmoG6oieJC3nEtV/+YL426
4hnvQLmllU4A7AZ35jTfGf24RYpidBbwfCy3V/pkPFa0/fxlXgksCYUgF4Ae
X+nkp4cw7PI1q7eZjrud4sPuFrOTHhx6mlQnvHeE+gJbymf0pXxOHw/YqkzP
MkJhegjBYLoKD1/d04JUQE3GihR9DaQqK21GSfrxODB1tDEIhN7z5O7NWC+S
i2B+pFxkbmkVi8+c6jq7WzxHNRjfsUxntVPZGu33DHfO3vn0YSAFc37EFMJD
t4YQkMICpK6JDlY83ahIO1uZG2c6FeaZ4lcgGDOjD+ty6j+tA1OA5jeNonHS
srAOlLOS4/eaBeuxLEUO4DbFhV8gYgZXXopJVSme65tTVlbktRr6kp+mMkrn
7gr/nvUHI5VfQl4E3eNhyLbu21+3G+Ptt3Ms6DskzYxEf4l7KcHEQMEmMcC+
Ho71T91I14pyvKrvzVlPpCOZcxWft+hDXuI8h9Hi2mfRzCJ5o6foVRuCbPzs
8VdAt74z/b8og1T3+bgwE6ifRWdhvRx+lgHKTG9eJnmg+1B2cOS3rVIbx/n2
xZexO9j7H//S0OHoPp0NAS437kFxwgQqkh/ECsG1rcL09nXxyaZiiA1vwzC4
G3DaSbdhMUkmRnQ1a/bQL2ovZVEFRWgfvExu+EK5MZisyPVxAzm1M4fzqK0U
CXRtcO9JBENBgfVb1r8gOoThbHTxG4DQNK3ksJy0k/1T+5RiZt5+SDX3ymlY
VWmefkevX0Q/zKVCqVq+vADD0NlZAWWAUJE7R8Dm/MTEhjm2/M9g01vkOWwU
donh/0EXQbd0m0wXvGzaKmyxAiDJkSD51+U1XT/BuE2y3YvC8zoRMpmTydcI
LvqUuXwFCRyD6WqtDir2CWvS0vi1GHhXsIM4n4bzTgE0oZF64CPf61F4QRB9
zOh4qZTr5gggO3GWRyy+ubH9JgTxt0RGCNnBbvtHxjDywmHx3uTy/2SKV5SH
EbgLgFdyEPrYdq0Hu/gk9QMorCZ7/bOiT5hbqGn1ZAj6eSjGxv218nG4vaJE
8Xu6nO60fsXmQJqVNqG1jeJFVUFe0PTLAYp22CmvcZdThUcKp3gR6SkSkkiY
NOK/KywJBTKpbwZ7cWEWy16vuMtwPc7NNZ2YBTd08V07yluHc/vBW/l16rGy
0BU+qFpUgoEifn6ihL/H+vN/62LkuMA7RonrpHj4zU2TfhnqCS7rpcEGAH0p
8r+ESuuzkGbqlSHo0KvRQoUFX2O6gujGVrefTkpt8Jk3OGYjYJ8U1MG4NS+5
5QsidfQaxJjgsJ9HzSRKaZt+b/mOn2W9nfytLl49/coCngo32ZvWSQp88NUi
tRFw2ey0na4qVuNU7+LdhQvaolr/P1cUynhnkLdPd0t5xaLVsD5Po+d3RH1s
382n5T4GMVi0vosaID5+8mwGITQBCuM6ybkPbVOkVRRUpBI6VvqiBck3DCV0
qvQL0XVMgvPh79tdqkokIHwLFcpPprH+5mmmFSp2DW/heskuQ8ecBQ5sEGKS
cpbluNxcnhCAS2SLjNc2dPz1EQfbgJUHPuIHuGgSiIvY8+YDW1v2IQOEcrpy
KhtgN1OvIOFddRQr7Kt8M8Mc8rlHow/wExOZhEyMwMLmYdnXFuoASGrKLOHi
o0gfk8HWyrZ9YEkpj6ZNV0VDIbriHZ+u7L0VdgpOFQQxlvPu7atWoK15ZIqb
834HxzZ4Zydp4h7IYo5zieEf4OcqvCeWxu1xSznzurmQv1JOqamnbmnG+dvc
pK6inoABDKUX/JYysMD3+pFtqTWQuGYaaxDJdztpZvWBwXC8LhUoyYV7jCHy
tDH3Y6UDJqSSyleDNv57kKMSlJDP8IvnudAWKtdemHTnrJyM0QcyM8G/DcZ2
xoo+ds7GuI3AEatqXydmldGNkZo3tzVnBwqzmDgTegxeJVzhy5tJkVO9gwUh
Zim9EBTX2EVl8N/UNe84SieOiONXiKO0rjv4q7e1HNwVIkvIRLYVJp3GdhGw
4zlvRckPqoDqYIJuyg1k9bZ+TtSpg5UyhPLfIUQaQ35tyRHLpCmE428Ukpsa
xhtrBjaHFv+Y9tetGJq+N2j8D3DYRTkAbFlFdCJyxuaNqCbs34c8Q5IyDjtZ
khSEHja0UYWhJtzEfPr0MO1qetxKx2kf+wwq63fCNnUpQ+1LKk4tGIArK/0Q
+qWplMvyT+GsI7Nlb2G6CFtJu54TvLNwmjBOZvoRGWzee1z05VyG0gH7U2C6
dnEM64pXk55WGSVHXX8wQdXRu0YpGVbR1Tf58Upo3jaWvBYn7nulgVYEraxW
khR5WDh/p5s4xeG98tzhbzuevLOdhlc8bNCnXQ98wy9r0yeFATFwPdDEw8B6
Gwooe8WypThTqrALe4FhGA1WXj/gAAHxtc92zgvjr2dPjUtrLVyd6HCbhYMO
CvAO56gyLijBmkF+qFTLEmUwcPnmgtzM5hHWUZybEv72X5DEi9jNzn4xonwV
84pel3zQU502DxBl27SFgKv9LS/eNy96+HcVyhI2yj+5DFNJOURzj/5cnn0l
kXoZelTcdRDUgYG4enxo518M0N/FyiRc5TvxMhw37hFd95JOCsd3nMwCvyd7
exgyvk2Dd5QrAyNjgLQtKtNxbaeEsNHdhMAAR+SVSm4DXzjegPQSUvag0nTY
5UXPpNLuye3ghKmp9oxGsYG0GD+isu2dowrrZ5KNTjGu1jWnT8fUGV7NPXkS
vJMoafRJXWJ+aGxd1FVePPTGgSovKiU2cZyFsgnlUzwcW8Jh6KutwSvcyLDj
8d5Hz1cTASegs0++/6ZrJPARaz+8PDGypq4V3yTso8RStKzH4BtONIr8e7dF
ScHI9hYas5W8YsCLMXQv43DCrtyGxdmkiC5QWTmF6nEDaOLGZi2OdLjWZ0BD
IyQs6dux853LKJEPaaJkHfuHMQeQ1Hr891o6YjauIakEcKhRboXBjsn/R5H9
bVGbvUHAOO+2byevwBpNHTfr/fvU8rvMSNlhkgatms7YYi3qFzOjYxjW8Q+s
DXwqHpr/3U1k4tqlF1xPsm2b79Z7PAb+SlaEHPFSBMrnV6oJkYSIQYDWhmli
iRGF/QsgXfC6v5VK8/oidDHUNCyNqf7oRsv+qVQMmQoDjRqkf/wdlUMXl0Dz
91rmkD2Q/fOLrxwf5gxUUYiGRxguQ57xIVYcNBQSk3tBKyFS44gpqK9NQP3r
a6C/EfiT4bqwNSDDIamxAUXvp9XLhXVABqkaszM5PCY0oSOfSaM7OwiXkFs7
A/h03+obYnpcBno8YjiIEc0CK5aYoO5s4osNC5Y9TmbKkeYiEE/IweZteCgR
qyYKiuHfgtLoz4eMVk1eSRqcnbbl0kqxfyrqkdGYYl1FaJBdDi8+mSuBeg+r
rtoTsnuCAneRKczxJiEOtJXXg6uMCQoDBqE3NglyV/VFIFPM6xX6Zvm8ZB2h
srPGatkXpSomxtvbl6y9QjRyp2KALq+a0Rjn3OUS4HM0rPkXsOAbtzWn5nT8
vSmGbZeK5dneWlFJQCvmT4syJ2jZiEIWBjVR0NrSOhhwy0yDzbqx4mPOazKs
wC2jPgjz3K1aAd6nynFLx3nZntosW+8oxemF+US4EYcekdidiofTXu08jNAp
4PM1TvIUAN7Grgn2so5mUNWghCwzfpgMK4ElPrlEh1Av3wf0ay1PDKg2ynME
+Z5XmLIAeD3S0CQ1Y5ScCF8xGWS6aeQLEO3MLXvU349FWaho8bYrGXMpelAp
dcxEwnZYi9SF9bIGYiwOnwQ2/I5RIbalsO9j908QE4GQIYKVe72T6es2AeWm
aAwaKiXxTsyBuQaZagMalKmU9LheQTryWMpOBm9x6nhn0E0MGwtgKQs/bDDa
krDujUL4C4FW5/NyMj0FN6OoKV66PHt8FYcW7XOc4CELOjD0ZOiUiTU9MKVG
kZ4Wi1WFFmZLzEf5XdOon7u6Qnx7U/Udtz2ANPgLFsSyTqtdWfvkiGGAmrQp
qcA4n5CfKNC0SMfaj1CXWFS+71pzNEJeNgltKhqApYJCKPQc7zxbiAFyPKga
KgtKnZflLPyRHPj20+wu/4W1zzQ0VjsB96raxTgK2AruVsyBAXCsjB/loE2Q
vswfs1WtJPGBEPbKMItFaaRB4uVwbeJLg2haA84PdrP+298HxAKi7r4UMBYb
/tntxBwZtKZeW3s7xqtmi+mBDTiUTY9McBBSzPkFZ2KzXwce/MEjbJnOASKK
pVr6GBGBjh5tntvjhZmsRGWIrhy1EkkDN4qhI2GHMa8tfqq2XV+Dl5FE54lR
EaVOp1TetGdgr4WRixs9hONt3/00JCcHwijImfTTBErt/GgY0XCqQ6DdvMVO
dN9DhJxQMzk8LzEpo6sTXpAPepxTJayCnIOjh3um38/ZjFYx5HgPqnkHUybu
d8X2ww8Fq3c93//0U/G6k4jai8P8DYlVCMnJXcKu2v/AE20XL93br3S97/ox
YHkKgUAsqWDtFJVyEkL+LeIgCXSgYOKXkaSWa2KTCWEOkmIurlNUCm2w9tq+
BujBYHm9Sny1ek6toSyQpGuWDYej5Eq6ZKGMJ257wDurVajmxfwLIqqhq3KH
TZVBwTz5weuIbnBOzeswSSEGZD3M89mPOD/9nOxdnOfSOh0YMkgJU3TscMz2
osHl2OFd3WBOgr1P7ykDcXVrfidjQGiEzT8JFVBUxaRk1AE3mlGtwcNqgdes
jVNUe1Xjlu+i20+R2vE+ddEVPfzcs98cs9HPr2M5xN0lcZJgwRoOaz4whOzl
juHffLar0USNBPFbEZ2zzmiKPA3k99VPSYTyrOpj4+WvhylssKgTrkE9eimi
Ou6obNxer+Kl5E90zyZQZdZ6wRDV7l5fs6TOJFpafdoSS+G/FU1bdTIpgs/z
QVTRgK4qdq+Ib9tckAoiPn9zclVOdWkWON5szZybKkYWTsOFwaHZCdva/8Fj
H5ZfxnTqgb5TtGH2GebP4rXjUEufXeWSzmQOSuSZyYjSc9w7iktcTFVyGBhI
89qdGsx9h3eH5vWcUv9hyohwgQU6AUGllgL1XkEtCgBjLfwlVddehLNM8LNf
eHAIqvBayd+eR6Ac+WU4SepOkOM96GQpqWE/OeOyGHO7c4NIW4wOKk9K8pLV
mIPKWXe68IkRlWQWO3uSC8VmDLrvN1thtioLHeIkLgoUTslqv8rqaF1Gavkv
8VcvFe238H4cbjKuHcT21JVB56dONJ85BLwmsCUNm3ZBmWDvMbzDlaxfOwqM
/xDWZ+1LtflxFuJXYJufwiLfJhwOW8OvPi+B1XOiPvKiZj+5wrxNu1GDxU7W
BnO1NXBY5qLO5DsFGyW/Ir9MrknyqM/9goG+qMy1WDla2KWuYC6n9seTBcLM
yl7IkuENHHfqpkjSJ5LjQdQP1STlGLfp5zSdEeTpK3V8BHjzIO6t5dNVt8wx
BUkpH1fQweqVxoyqe0+47XuRBKtwfTwf4MbxSdwoYGrFgA+oCl2oPAboC/k3
5DpDCqFxD6Quz3crgdijUCAgXdVpGI6s1nFd5akk7Tizgc5Zax4aLF0EkTGE
8h2mELQcjJ/H1/pUyZ4Cob1TTc2SlHz3fT9jWtRb/vvGH3JW50ieCOb5qGDH
mbQo9YJAfZaXARqYxx7GaE7euAJBw0alnQzbe14n0eiKyr+FVTbU53SxL8zG
9NMdF1MGJ5HoLpvD1ofrOwIwZrS8qC2y+uYejvPTX8u+GwgVSI3Zj58BW3Be
WOoCd5Iy7w4R0mYFFxMEeK5IURfIfZCdtEtVibSfFHBhemGU0g9anJr078Cy
y0tOMk8XXcLVXBHBSSxRwN8YtqopW7LqQ//vpHnT2ypf39B8XRFgiDyrTPKL
lkhdUJ3XKXVmcP4dP0g1e6UNHCUa8UOfMmhC9CHO10cZPe87nOa7SX4Gu079
y7ofzaryEs8Po71Ltql/D2uiJ4jir8zY1X22i6VXD4bonJiCkfQsZK7TlkyE
JLU+Ys7iRntl3uOf0H6QaqC6iqXVLIGB7SJ/yoBS1BX0R2eASvUfM9kTq3Io
dzdWDTgixWTsPbECdI0P/BUHnSKUPWK7/h20dbc+20ES1kAj3GYNfHO5cJEP
OIY2XWZHNzL6DzGjpxZWBN+Y4K6Dwk3uq0+uubkSt1ZR5xzzHruOC9p+1Lwf
F+nGX9PE+pSiJtwJX/v9FljSs7D8OwCLsqHn/Kpd655rNl7cwm+dn6lN5M+r
orLftiKIo61C4jNX2RseG55YnPfIalW0/64XhBc+G3aOvdeifieEWpdnzzwW
2e7cfariYt1KUEFLUQ+M2vhvDNpiN5DXM6Bc70Yl0JmkNOHfFt53xU16dgBl
J1jBf4I34fUOcePto3/nfk5GDJIkMQzpgt4onY41Vun6p4cWotNp19sIi6rZ
SqRH8gJ+FSRd9fg3xpFvwfbHVuOnkmIbkUjHPtC1zDnWEkwO21LqWZUC+QSm
KKyblf/QdbN8KUzhtwrWGG4LgDndqsjil6+ZmlqSI3/EeYdoLlI7EFljuxVN
6lK5BSNRHpMaBQg3IIxrqCfIILD961L//5G3Cx8KKSD4ZE3PctqW2ZIQEkvl
PsCH+MIDno4LrPkdlt0fOuI3tteET97nUXRXNRVamQ7qKpa/SpS3LNYyybrv
0m1YhKgKVcby5hn/pL3EIJoAclan1Vi4Fc6fZ2jFRYugcvFE1sddPuiAQe0v
fyPScl0bDZO9/cO9Bgo08HRuhVrHUrExzsaApU7GkTvTvCekQSSzNrRSnR9A
s20vv5g3gWxH6/D6/GAsH7+cx63UT+iZVExm7Tk8q4GjhT7901UenkBktQSp
/cLgfEGSLv1n5UxNlYVwOqnsuh20yMBcMZyy7nqnpFxH9lO+WRJIGjVTqGvi
Nzv11Js2E1jBuZlmWEyaZmLiLQDQW4yuS7/jBhE+CME0CMx5m7Iw315Qa6I3
w9pqyyVrJPfIaTvW+cEWTkJAJARwkTmjdJC7YAqn93VyMSjsr0qKlDg5kHTt
XzmGtZSzpLRS6spyCROVoFno+g/Zqq43b7j27cRcUMcVWLXuG9hBmYqwjttf
nJ3T7iAvQtJV0btZkShRe4Y+/0uRQwby5H4nVNmvefi/+R8vTXp1aX2gypM0
QDY38XtHGjkDHcciimbaSgFaHLxv431HxmIB01QuZLE45nWzWeSctGAZa+0M
81Gf4rzMlez1m1dl1AZuGE2Xx+ORbUo/ZNc/Ds12GOUW953F6aXW5NSig9Ll
QTVCl6YayTyw4o+34ek4ospoz25ZMLE1upKR9uzly4ephxJiejQ4170Ra7Zk
uz67wx/1Iz5nmoVu0ZRbjxyhkxnw4Ath8AAesSEp4kdr1O9wGJx5PW8lNF0v
E2Kq+NXiM0RogLnKQ1S4p0AP6CoOL7xhfg88MI+nwsjjqeNG5sf9uM9Bkmnb
mEjt3gBkzh4/GmmMPJw82kC5t92AHDpXfptVYUpcslUL3X92FSkgX7DUt20j
ASuoOePlDrTDBcsP5giHd2GS3jht41PaIpHkPkLt3qsF5aMJSKrln4RVaolr
RxrzQExxyIK9hdq8xAfU7cYw9Ls30/sBlzIc3VuQH5kWJVCdkr8vvukzgua7
diHdW6WgSRC8rwP1LSp8APVrQtGINSNZXRI1kHwF6iLzgHuAfjqLBeS4zMnd
g5OF4EqnnrbpRZ5jN8P6QnxYTIbyd8uIxLbZAUYZ1seowx9fMa05EWMGVJKF
71NHddqvoXomZomG/2Q/finDtGZvgZoV/jJMnUzkNVTZ3LBw132R9lpnWkPC
u9JC5EnGlpSBNxQh5OzkbouhKVJfMH+1ZubQlRe3ZgFhRmLK/v3M/aLi9f0w
V3PGgo/zcPZq6aPm60yZ5BuwWAOLtJc4m0kpfK7aT0SoMwyxswGOoBKyifiM
EMOv8i1hqeTBRQUKpSPVXuGjzd17bXqZ15uy8nw+KONboHun8nj4ycI305rh
sS7FqF2/vHo7N7d0yGVXdcAezUnbA38qxLNvSFtYfKmJUHmmHdkkGSN68nRO
9WvsP5VHRw4hC58iUqk0H2FJljavGRZn0U+19h4Gc7lDkSCHT6Wk/9tkPQoN
H/lboDs4S5gBnZe/JmRqAtfd9Xmwv1S8gYDYO6MbKGQi658IPiP6YbhElqVx
gMWKKfwdnXhIsKdryplPSb6udFllnlhXDCCjIszAkkZvTXPXu0up1UkAZxG7
1j3/TdctQJWMBc0hg3DTvTvW4VbyiyZt5QYQ8hFDm1s890EFJsE8POo9emW1
J9wrpPV3HjyQuSe/PP/mkVv/8OJwSg+YqfAcIb+9/Ufsx/GWSK3XBNM3/Z6x
xrXXXY6SPrIzg3ZyVsxTRSHgnhIIuqdBlshq8JgOFA6M4WL3P4f5e2m2D/Ud
dIAlHbUR3BrhWXd+GpoUnvwV+bliJ07cG6HunvjLzAItSDZTq4RkC3HTMYky
kLlp4Kq7/PpUzEP/qrw/P6a9GTw/upxC/8y25LANxm6hvKyZnsyX/aWYvDB4
B8epODQVxeAiFZ7SvAZp+/FYi5JBh0mgyo5rqQWNidrHfAsPMVGe7Npanvbl
lQym3jWG0ep7qobNWzP+HHK3Gwgz5j+ckU3G4aV7bRKUuRsp1i0FhfxXAsiC
2mgLgerKjI5GgC04zu5i5PZHZZoTXIgEN04i+J1vGmw+/4TutS5wmgrqkVG5
eWTb/gqMO4GP8EeKNfU1d+Mq7V2cWAXq1HoTMD7TyUDeGrC7n7JnlGZRWzPS
KXby+EoJ6uuMcS++GQRLenbp/UFrUBkXxVChUaJgvmxLdk69snx03pTtDaWJ
7qeR6IvebXoy3dOsqjsmkXNN9Q4asWty8GNJR00HyoZs2QQ3bMWFU2EQz/Ic
/ppMU9wmq+ZRXBS+KW6+NhrspnbaNlwpl5A0+HngflQntd4uzSJL42pYc8Gg
XP9T84x6IfCsvopQ7FYZAYUaciMVG/gBQXhtnlQsdiJSe+iR0gl2ehw6DmyC
Gq83z74reCzm3qfz4MjCFW4Hgx/QKOVMVwFRa0qjbms2VYF0cOlkcwyi0lcH
qIYm+ylHrkGAtZ19zGNXSA/tAesQ5pq5a1mcJKwtutv+Rlt2qZQM9gdzZkWK
MxS7vZOpYnJc03VtP9h1C8I9/u18fGYndrMySkVGDeZMAI8qDrpSDIP0Z6Ee
AEnCwzfkn60s5kAFBVg+CvTaZxNnMXaKc/aj0+j13+6JWzVYik5RB7iK8uYM
GD086Jmhl+5ajQOxJD7YIs/erRpLFC3TZ9PJVpnkInNF+oH4ew02MQKEwbt9
IvvRZ+Ny6D2T+YJxkTXkhI3559KBjraRVQyja1Dwehs7EiFrtP5tI/XUP97Q
bvUTib9ypNhAd4IfsQOKb0t+EfDcJyFY9sqnd0uX1bfSHWPAhdciRWVTgp5G
DMtZHOGF4Hhe0NismaCk8ChHLCS62+zOm4ErGsRikrRfJDaSlN8UorbUJnRN
felYQRKp71/gMvb/YfnQkxFBaLpTuEF3ISA7HgBGr/biO6sAWf7kqZowCXhv
vYgjJ076C/qK/+B+kLaWk9cVzFWd2b4VikqTgE9ts5+7Olnf6mNC0BBraP5h
hTmuEIUeMOoCsEgBMtbtcXmgTcAJ02Wbae81+CDSIbqcO7czXJ1WtqNQiR7t
27jCwdZpKpuuXaVklmF8V8PZKtITR7FSMlmXku8FqILVkDbOWYspvAw7c1SJ
zd0e4SQyF8PLw0rSNXbglE6WYOjhGXyLNG2d6rzfRm/jqBBZ/5VvVSjGbkbr
X5hAEZ1zVZLGKpgesMnUmjiJgOTejM2UuHTQeSPvxeogVQocgVB6LwMn8GrC
ISs4ZKmu6BQtvXbNIggPBwgTFkgZ7y27AQKhb9nhVQclpRjr5ROm/IHhldZO
BZaNoQYkiGdzBQnMjq9cIgf1EVJbmlaA9HbyixOv2sKKCgKCFMBVqV39+N0F
wigOVMT3KmlMSzPP76N2Hw0uQPYCp/iJoL6uFc3kcvrlIElOA9rHMthxASUg
HaZIzlJEfhSSGKkIgR0dQV/NbOxmTi7dGT8JW/AeS7F7Z/PfCMRpQBgYF4WB
7bGYJAAv+sztj1kKTXu2RnTsP7n7zJxEpGXm41V2meLbUTJMHfiODU/dOZUo
rofQHf22yMDr3tW7UHRf2VDW2UEf31snbJcebq44u5OLFXDSTcAv/DxWzRfP
ewV1wP9O1IfzRGNGT0wOnpXgRR6lq52zVMf8cKj7fFaxWHHMRoNFYyugtclr
4eG06PnM5rY3PyCLwlxQEBFwlSHRKRL3erXfhlkyCwq4ocQLP4N3nWgLsWFF
Rx2rxMRC16eqYtx1w6HsYusecIMG54UHuet3b6tfGIlx4xeqXwlTvGkJG61K
QU48zQa79EGytSN3wBdL3Q/hvkicLi/ddbRDcuyC0eDDqXgktW7ih8eseVAo
oGIOiRzPlbM/CY4eZna8DdRYkgKcdujeTGneArWICxvuz9REXt+MlsSyrf2d
6HKEIjMIw9ofCzEm0KFwPQopG0UzdfuVnrXMeBDZKW4vwtJY5to4slN5LzlG
Rr2Ovsbn1Ba7DYUblnEbghehXnJn2yZp4pMU0n0KQ9xqI0RKkAxrCavmKIMm
FEOeTcifh7N896nEcEfaSC096zXFybnDbLHDq+JEmJta3ike6RFWWssU1Zcy
lYMpKyNMN8PRab9ssrQsvm0E5Nnzk9RqODASMMjKzSTmg9GBfGyOoxwRygrp
uqvkACi+0t1CfjQ/x+6CE8+3KCHwIvsGJKsszi9yIYxC+C2uddukfPOxGClj
Lq34UaBPieQoOuAjK8nVjFX9T7152u+yeCrrL5VrNGLzKuT1iIQRwtcJJwVi
AXudULg/ur1IFJy7kdcEyj0q5yHvfw2OU4CKQ+pWHM3ZnvW9ePUgZoef5kON
2jilbO2RVws/n7FJsvxJGJ1ZtQ9h4YeZba/+y7OLbOrrvEfOOqCii07IGmJM
vfDL92XfJ75oBsw6Z5ImP+fCyUgK1E+B7S9XYoXqPIRFH3AcNL+EtVQHY351
wUCdCEeyGENZ8bMrO+VC+JMU9HzSewXQLbi7cs53ByGmp+V2LhPlbhc7UBBz
hbRMIhk3jMYlLniKToquR8uHJgfbr0PYtdkiSc60k0NW/gCdg+bUmOqEUxLn
IrNa+YzySRJFOd/vco47oBmnb4gHqgCJKAlQNGw1D5bSlj6BaIew2H7UdGjr
WYTkusHmJAYAy2b88zb2H6GQfYW1/TMbcwkCzLKC+V4Lmj89IPila9pFFafO
LRQpRY41kdWmWXwGFjZI21WGjgBZ0jkrDXFv6IQj5ti3xuKtMeTprGJ1fTqW
IvsXgOlHlYU6Cvua/qT9L3RkYO0KMQxKzrMFOj1G8Kd7iYsRQldj1V+utEbm
uFVW3lSBxOIQwvr4Bx5oKw66jDRAO5k//UIHCEXjjMsXRcHeL7Zqf19yLXX3
YpGD+ysXkXZgnJMYdr/qI+x7Sdwag/uroVaNSb9NmkDtqKnWEeQvi7aH0g0t
QqwZkeQU4ZODG7rgqdhGdrR6TI9TSCrNOkMNVe2GrzsUXcyl+9etrJxnnfW2
urgjNa3rtskJqBjKWww/K91d/9AZiFZ7Kw6L0kAae6POFswnEQcAk9v52HIn
GlL5zYTOPKHbRt7gEIRDfL8fxASMcJ+pMYBNISZR2qoS+gDylGJQNWnkwUrI
/fM89D9k3oP3CaHfw199ddLNrwlcdwlM/Gl8rfpT55oycVesjQsQOjQ25cNj
J/f1/2IUCNpNstBkYDa9peQ68M58hc9nqyEw1/FUgOnGKTed9D92kD2xr+Wm
JaoLsGQS4oiMK2BzE3v1vRUwXlRynPamKsFhG6s94Mzv0CiGB/0qh8I+tkIg
ju7rkTuDlik546EWd7WPa6L4PiPpe2HZn95viCbSfTn5/F3rN5XrdrKT5xov
UdeMEeH2XIgxdZLAiZ0Ykt/EjHOfkd16uxhiimfG25XyEOhr/S89x28ScN/E
WljxBRYVuNvk1BVOcWl6aJItcDH1BUMoMHKt2CzD2FPUcsn+rRGeYalW524L
aHf490uI3tSimMI0tiEGHoaMFf+D4bQsHvZXZ03zwPwFUpspu5hle6eRYMpy
r3MIuIBzyz0J1ZBDRLc7gzewa3OQstraEuSbOMh4UX7RzHyks2AoLbErrdLA
coqQMyxOdTRvgUVMGXWpAJDgP7p5o8jS/tHFS+5ADPPoELDxrAeV4r9epr+6
PX+zub2M+d+gLkHr4L6FmY1U0aQVCKERLF1hLs14hv9u0l1dPCYbYNv47uR/
hpy3Gr/h+rpt1BcLbaodt1kHYq/kYJ9tS4Fel2bghBtCwIKDdEqWAS73UT7y
8r2g3VRA59TwgJzDzMWtX43HhyKAuJJn/FsOYSS6U54Gk7suBwuJIjlsWMQ8
M2Da1guxI2v9/OeHhaxxoQYLuvHm2Bh0/lUa0uMmGWWVuWN6Lk5/A8WZi60W
TqQt5btOwCXbSiXHdwDcQHeR73s8xs/vDrB4Tx2NmvSguApL58UNPJBxMFQT
/rTtvBpW0HUBbtDqH3AMO8nDG/X/tAsqkVkvMlS3cFCqGoA9XUFqKsOIxf38
rSsdNzShDCxEJT7LxIlLSam5mbrfjI3A5NdTm2471KlD0IWBIHx34lZuKsRn
75KNQxbNlBsqKE1pflGT5SiIbtE5vm/wwapKysiiazIFEPy2N9YWcZ+oWztu
49jW72GrWKK0UIDCiLohkBE4np3lIJTDsDlAYZi+vdRzT8Sbr/cHL+oc5LLd
vWS20xfVLPm6xyLOPkg/yCADZKHI7CPdXEf0gTlY47ucMhfywJJswH/Ky2Zg
256duaSAxUtgVFKs28V+lE00nIsNWKH5Uz8yJlpA7pKUmWHeNJaW+JO31fqf
qIP2eTuJ2gB95KBId5blaXiyFB+GlAGmtSRd+5iQWsP5hmlybIdanJOcc39W
CJTLko1T9kDeoeRT7YzzW8WIdjUjT8clzlDwRPuVi+dOf3ldSDOs+W6Plk2v
cOyWPpcddccjes/nVXmYGpXuw2kQK+MpliacViemM6Ju+RyppKQbpyzj1QZ6
w4bL0a/glyBwFiX02dY3uicnImodqVjuLhBFT7J9f9A7VHCqbGmTqr+0XkgM
ypHY6d6rcAuHX2tA6+2hS9CmMKGh0DIc9O8mhakEMp23K0+itf56a9sHhTjK
weBXhyj+7BUFjTt1/Ivy6thrjLucDGY9Av56FOmlwoKQMzmJMNhM0qWYggwP
cOzTbv/MnWxz0SEjcBkYO05HS9fd/z054WcHDXWl4MO6rEWNCSkPDU8toac6
on5cR/aJ8lnHyp5yxKV5fldKzpvSs6Pxi2GgS0UllGCEGsvIrGYOrlhF771q
IDMKSoVp+kQb0RF8j22TnQUoW8/P4Dk27PD4vOJtVsNuSRN5BpqHRcsvtxZs
9Weez9XpnQrtKuc5zdtSrsubmhs8VV9J1BfUF5ZdhSTlTloMuVJcMRBBmnG4
Z4BeqfuwkQIWN6HCWgIrix6IxVruD4MyA37KkZyA+H4H6IOkv/JMkRN+Dq9B
RQsQDTNUu6+GxHRP6z8s79roa8jrN1nZV9RHV+kCp70G/MTRmDVHnOAwPA1b
TFaLH01rxoro9L7SaBEXaVMPy6qJyzaOH85zare3NkZVEQwy8xEw9NTBlhqi
NFGEXZrdcJOBihHN6f2aYCMz/rO6dNRwtlPz+LBB0ABCpQ2EoiIG8OJATrMu
5ZTFxlqer2F5yU9x2k6Lg9NFTi1sjVRPY2nl16IMswzDeGL2Wn8Ps+0L+6wT
+tuDcQRg/7H7xQTTK+YTUPRSGaNf75w8oASjmez0r+0a63oRyE6pKFnb6LwK
AeWU9RLMTR2NRCRTYPVClh3nBO4kWFWPK67dZs5Qd9I7YJByKSfHIwFWKVYR
JNdAXqZZw80VIwgGky3eFxlGTJ1shm3lktCw7B1fFNhCpSTCM90//pSEFn6F
IdCwBtV+smPXfxGpxVMr1pYQz/FTs0h2GXIgL1MY7MepVzqFGrAMfoSO3S+g
0B3/QP08Uyg4ZWjMP6XwhBstGQqEAtQPrLnnHbJ/tHZhDLzuRpUifBAH0ett
1b/XusZotAvBOZrkJAmFfFU35L5Qu68nn71TuW8W3XbGHMvsHxKBG2m/CbNl
jcqleai7s7Llm7cbXWw+IxrVRhpXaQZQSyIQg4BQ6ArgXDtwwxgIUQ8wU5lk
oawV50p8YvSRmnkFuRyhaHCRSkM1jLN7H0catfEyRTI//NI8UllIJfIYcLtJ
rM3wbEVsDO6+BHgTM6jzYw7m0S1qgrqMoOtz/pBE27DJHSmT6yCQrsInwyj/
iKJm2kHBinVpl5LNifimn27DjRcqCt6CCM3XZUGuefGpcMTwnvrIkVmyr0Or
ZriA3vA1Y4+u5El3p4RrDVhvQXp2iJFaYmTbL/K2Sopb2rN7Uum065ppWIte
NsZ6kZEg3V6d6v7jD7YtCPV2/452HVC4TNoKwnS+4OxxILG7JVgomBUtW5Bm
6pw77CogK2b1jvmqpTC+x2ToP+LrI05c6AJNGO0LluzuUKSx7O4BRw6T8twc
LHzEleXYa/fOIqVQSJ0kmHq0ImVZ/TwGaQaJQfjfN+rw3SCo9H8YED/IYFAE
KKk/V3dNPEJ4nCoUwq5Vui78bez0TN6cvpXCsb6r8lbO8FoF0VTlHGe1YbIt
mjuRgeZTjOHD68eo38THEdZTmBS2ugVtOLORUzxY9jMJTU6GtL1X92F2+4Ds
GV3kZPPBp3mYLjb6mp2bxbQ2bnqIBsOs7XTVqWsIEKLpiHSSrUGf5Vc+ynvK
IiEkWKPf0PjVz0RX0iN9KzxiNmypGRqpTWkMKvGiXRAbqC2+3SQOOtoU85mo
Ixouum3fZxXmMW34q15teYehO38BEl+PGYu1g2YP6WL0keNIg45Z7Oy+wML9
wf8IxDpaRm7Ooyy8N1zz5ras6nqVHlU5cGfiPNFXVB7aF6ivdMAxkq0OpKfg
PUtPRnsqtK5Fh5dSTSYwwPJOtQG2x08wll6KBl4MmYSjZVXkd9LrOondyxDU
fEU9bMmGAfDgiRCvkXKG+ZQsnWgQNFeZu91q1qhUrg9DMxY28KAfW9+DxpUg
zo6m7ifaZF2QB+3JXPDu5JVNlP7o7hpdRzl2w8fM6ACIqTQadkE9orUvknkf
ED113isIyJlbftigR3ck3D47NCIdXP/2SSUh9rIXtcWdG/j7DpeaXf9twjby
nv3XOW96wIcjZutU5DueyhC92S9TUJw7wBs0Yo2QakTxtLttp+bKJq9Gq8qm
bvyfe0BpLKzZZir/gZo0Vhlga3NIIQ3vUrqcImaAw/Fu9aJP/MZpIsJRc8QK
Bo2U2/OLQL7LJhVN/LjG3sY4uwz68H7sYlmU2HUW/0MmrVcaGSlcv7j1YR/E
7doXjCv87zAkudo97mqyWkEEZHtbJAp+YFjRTsXkfCCo5wGDBKirTKcjD5/1
Gc9Gn46ERHRasGSv2borRdRerPe1nCNEsP3/2SUuphctj5RUEYvKYzy0l/5g
GcSH0ouiZx9ubft15Te/5PULolCS3lPoYvanl9+a9zbDpP5wRx+SfU1e4WKN
zkKqvyytVKXewOl/no4bf5YH3VSSQb/gtBnPqhMA8X+wbeSwHSYXXvPa7TXi
RM9M8CZc5ZzUpZAPv4BXSr9z02mToQ5UtDNuldgmgIQJL6vSJeirVpiO8R0L
BHcfAVPcG9qusfil1MQH0SxmwmjGa3C3vECUgDmyZlNhcJTJ5OYFHCQ02GQd
mhC2cdGelHOJkT0WpionYYSxY/YFUJuIkVbP3illYSoyfEdcISIyERPYw3be
xQzY0rDAHGjlN/KMI8CsqNdbmBTBjva3v4W2alOps9k0Jxc9tMEKAFy9fU7R
ZLLoW30ostLZQKRhDtFRzo3RzFuEqDxaPmj+oxur52aZ5ZNPoLdbotLdu8af
zcEoiISpZmOn4QmE6ywbj9psDApKj1g1XhfnwdQDOV5yZ8I3yFp9LTr0nMZh
MjaLmcjCNiecDwinE6NS1MNyNs719gUDCXv5hIn2viiSmAOVq6AX8y+4eSKt
NROxfChZXvdrrKb1JtoMp9D0869m/1dVeoLIReoOJMsptpLuaVRgwkaL8Kh9
HqwBbLGW5HeE24+S2p1Ty5BXjbf8Cyk03rPOs8A3NJ7JFdihpAkdlzrSXXPX
cQn+RHkpJFtbrqD8Zgv6j1MtjlsF94+6Nl0FKhvJVL1Yw21OBGskxHZlCse7
xtX/W4DzNn+oBugMlRv10jS897GlF1OaB7HzIqwJLfqij2xzRFK4GJGHePDV
6QhGIY4qCx82b+P8QNt6GIDII5NeN6fzogCFA5t7mMuJB+nRVkJhrFt5oWrz
wRvD22LzaPxhkYENep7cayKIMJqrlsLbUCmOcucwgS3BPJEpIZnxC4+35X5X
xCH7mhZxcEHv+elSPL2TgcbOGsnaJG+srbe3EELvoq6E4rzQRVq42XcwsdAr
7ck0xCwpyM2pE4vbSrO1o08l+WxWaVqd4FYgemgGA/Sj6pBTBc3/udM+spMU
bFaWVVv3DfZFnBBk0IKiQIpCS2+D2aaZXMkgF2OsUAmzCDQ1iAIkFaU/tNBv
TeGdxxjvlQcNHf/yf1qv2ju/9moqXhL7uPbApq9NMfByKGEtSN0xv2ywnAQf
a08SdzxDmVGY+ctAcW3/7Gu/wZjLUXpWVCaiH+gFg2YFBBWJiE4HhmRjY45L
iWLtzKOR/HLJjoIx2hv+kVZBrkuZ0dVk4YEZsxkFnqi4eg4pYdYx17cflUv0
fpTps1rjUb3nXsNA8Z4InKID0ENnz6Xrt8YzPJGHC9NLUtgK307Hq5LTMSXS
YI5daibALZUH/+yvOqRCWeZNBWEVU3+pBHDc5TggsI8P+5RGVoiUm15y0E7F
QLS2mYuZTy7Dt/+YFqNZ6hwT+65sjSQ1P+ULX940BLaADd8ogXvuDaixcz1M
BVk/TpHf2PTpQdYzbMyV+YjDgspIe8/RvJH9BEGE8ZVPxlYjEZg4Y7dzdpfK
2DbnvAHWG3TbInYQ2XkgS8RLeMK6zY9fY8PDBJnwRxmSOkz8L47oIgDdOqEi
NmkUoAvxuj2gmlG5x9mMoS5g1ue+/RKjVhQ1s9B9I6NjdVMlSquqDr8ohAKl
/BDA0omEADhDCKCb5vHuH1iDUyc3iwhMBhyL2lXheHXE4r2jqvdruHxUZv2m
20U1COJy724QPiOFNbpfdFdFCqC0b+I4iHtPngiFBnPgw0MwXncK4iIvEyjF
KKd3Thl/cRSqenjk7R6IUfYlMjH9lNZ9rqWjVIPP3u4DpER8qc37kAfcrn+0
MjJpvtCoTsti1jVQV6hhEbq5/yfJNYN8RcWWGUmeWPyrlVZR1j+JTGYK8w3a
CwwAANu8T6+kG0f5FyIwSphVOgLJNeDTp9rKLp4BSaluQW3M09XJcHdpYASd
TcSCLtypCph3xPylBqj9TLdtmms/c9XeKBAdy5T2JfBQQ22mnwOmqzZoupc4
TSJblxepezl9R//ZaJXLKRaR31fdvDE7VzEOAR5xkDcR2xydeugQ5WfEM5bW
d5TapOemD+NYRVYgxNYkdsIS9tQb3LghxP+T73hiXdWNpNtCZ6PYJuDXSy0Y
M9z3HdoW8OXcPP3+XBKInaS/TDZ7TKID0Jq6AQcyJIDdu7mYUnEKPHhpIQ/1
JT8iAbVr31nYQTxtN0hlfBi5XRExdHVPebvXusHkXL6ptgr/x90M0+o6kjQO
W1K3/SkN2Nm92BhrxSVx6sOfLOOtxqOEuL5JfYw5AGLZw5WMuL8cmD/hCyog
sR157GN3Iaare60v220kjZc4biWuMeYevC8FzOSLz+ZxHU7Kw6sxys3OZlXc
DF5krWQq6ZsX9+xR2HJX1rtBLeyXnrRj/OEbbSAhN14zqVpig9CJ5J267m62
4LgkOiXkhr4hDvTF3/cIUCX698XA8D7l+hDTERLmVeL/Vh08A7HnDpzSeLGP
HhovyljVsllBt49zvwn+SewKv7ggnhth5tHLMsBkpPZgBBejY+yTmtiFYxKh
ljpzzqpL7v279ZDqJ3wJm4lVCxmBhCg6lDuw5NqX2cCl/PA0RnkEXRXE3OLU
XfiiMwFpyZZiSwRZ/8QcXKS+LhCK92pDbrZyfFbfvkyoK/CgtSGhg5EraT1X
5TR7uuFr7sEcp0ff4+9nQZEGr1CGj6/vbvrTaivneiZfs+UAsIKcVdqYfvms
QcH+RtVdtTLddxAPosjjvf9FSiftkvSNaKrS2N5eTjb7ohyqgrBwe3PCiZaP
Duy8aoAajARuioSzItJN3/AGXmfKDnT1NpR5kTaj7DmzYMxkZDpvNKIjJbdD
WIkLVblAWtQ1npx1T5XkAQ6pttBT2hyJgr24J8thFRP32t4rtN+syo69A/dZ
eBXijiymgEBlMC6J9mRdeJ/W7q8GUq9LKVtCYuiMqUZb0bXNVWn/iqvrQ4bl
vT8f2QEjZJ8hkXvHmCh721ThrlgYer83ZOajZx2amiDjHeYitGq4xeqRe0g3
5o5aHeM6G+jx1vxzw1/ZfE3G+JlPS7Byll2fjY1ci1RP89VUMMXaPrb4hIRH
ksMtYoLNeQf2D+DuKQeauaGRv7vAI7iP9q/98Qx0X7zktAOACgfk5qZrMxex
4fLoSkkkhG4h0IsOo9McVICEgRcL6Hwx0vjnmvxyDgJjGZz++2dtYu5gbsMn
+X35oIFXuA7SYM9bBIHp7Wd8LLGA8sPrQd3lh54pWlYNFXVM883mXb4l5MYW
vm2FHBziQaSRasb7mFkUGFNu8DdUR7QUdRtu9K7JJ0VZKeGn7m4OP/QP9KuX
H2r4n3Vk9/o/BOuT53eJD1xn/BHB8wi6I5/mjrKfVVbprlwark+CjLcSubO7
aXSF0wnXVA0LzUFa0VNG8QfID250pwfFHCMtygk5bTv0VLgxTZ25O6bgV2Y9
TZn85Un/D47PeCk2+8jf0KbnPhdUPAHqJ7W/qPMl6pXazsa4WEHq1XvBlcE6
+u6oj5Hfn7VHflLj8jddglcSKNI5+pcsj6p+TZ0Sq8ZLjALF1Rey2/ni17/v
KjjznGIrOIEOiAaYSr444pmY/un3KXxggSiCcpcGIogmSfQ66MSq0MhSUouA
2e86WyNMK/BNbFRGCRI/XNOoBl3uuaDaqlkg+wIh4h0yYGgHrEtXzgqq7AvG
bZo5evpOhGgQTQ8Ei3QmMD8eh2k/H7Kr0MlJ9HhdGh9zfMlHmAR8Xp9BZpf3
ze2TUhv8qPgm1za4/BlMroVoMEwxszseHyBM76I2ue3A7Hrx4TmaNWfe4GLv
GytlozNqOhI9r7AWskL0kne+IPDgEdcgSeXutA8+LKv2kqcmKDAelpUVsbL6
NC3aCUN/s4t/trNkwMUHrrAJ7ljYrKCpsZyGkeIo7lFeKZkhk+SIBoXBxQxU
MTg2lCXdIX+OkZnSzks9bRjXtrYLXwh3hdcXlLRe4fBi1ZhWvP77HaP83Ysm
VYV19KHe6nELXdpWT96l/emeEkMv1kM0+oK7v0PTGcJ07MKVs0TRZwzORK3v
f483op8A/BsFPBk4oM+K7aV4wrzAjPiBPfGUiqOdJH0owHB43+hZSYcP68fJ
lXQL7oJdoZqUSUVWWBgGsYJ7iysrdlJ06nHbQHe52cE2mDU/Hjcpd6qGPEBc
tuz+VdJ9MFJG3OctjcOm7LIUA2D6FqKgbbWc/lMJqyet59nA3l53CYcZTMGI
9K4KrC+JrMI+Wg/szMsAOdWSm65ntlp4LqWDbcMgjjr7O1EMrBhfTvbNCfAm
E0aAj4hgAUdUgOATFZHfCr5LF9zizTod6EYh1MsQrNNm4jfeTJ3yaZEGBHsF
UJXyu9F6Y/dq6c33XyU/ranay4MGdfTXoMPrtLuHptlCGRe6eSfah36//ZdZ
nL92uMZwlviuyW1118sEbfMOgcycnkswlRfqSiztRZXuw2k+uylBVNQpIg7i
lCvXWpAdnhCg6oREWk3Xny9RmRHIeGYSmLJsefChRIU7yakBxJMJEnOGZCQC
y52RmYZ8mkg1Gqzvi2c5eVWdpTtoJpQPjq3NqzWl1KX6pukgxRJPUlvd/Ryn
XqSrWuknY+ajYCTbp8eGVSte3TxnYrPZQuZjRHy3iTrCAHsSE5DhdkIsaiCX
EGLbBhBrjLT72BqJbZAGmZcl8SaILllE3kC+yPjO+8Y4E3USVr1apPQLINey
y5xWi6hCMZOsNCXNKjBt6KIYcPzDCMHZiKhogTa2h3eUWvN0wxT2HngBIe9b
mc6OIMusb4dWe3brQTxIeipL4lAIObP/vNh0TZDVOieGGZKgCKZ+Yyl5Acex
mjJmmlCfl9qsQr3gOgNq+lTRdrcHm15nVJt+KKnEWd+/yy+8iJ/tZiigz3me
FouWlNDyKup29CrymT94JAD4qpWqDqgWoeT3kR3h8LIZOiC4xow8Uj3JxkWI
XaSD65TbDGvGwFgvAOjgkrWPOQIRvttrvy1MAKjV5IXoPGGleH2boctg8SS7
CR6EfoWcO1KlRaZDx/I/zf7Lbl7ddgwdvu/5M5aD9tzG5d/OMYMQj7ha5ZHK
Tn0fZa0vnkQj7431kyGnA2PM5b0YWNhO8F0cK2CUBgyWod1xv1d4Prg10f+J
NF7C7W+TscSwYuA/93qJxvTyM58abso+OHj938qxCnGUaaGYRFXbjl2QM3//
Bt526uUIV7Cji2OfcJh5ILRXoKPdHVCC5g5pwHCL7jMTpXlxognQmxlYmI3c
9Ydja7uMKqNcZMzbCjiMzm0JIOidG/aQD8xhxb5qwSob+6EcOE/xBTxYVgps
SFvsM+EsLHiVxMhohvgVtl/DGaAXWqbLnA5nGkeBVm2olbiEs1mvq/pQLpGJ
+qGXHYNPXqMsdmn1oNlL1V5uKJ/5qIAj4BM2JfXb1HMbkrJ0rOan/5IKT+GR
KxYMTmhS8DxwPzzWFnfVaZCWDR5HhabbFGgIcAMk6JTLVT2kk7C7VSoCbR91
VLLEIcrrTsejm96h0jJLvwEnobldOqKd8Dsng29LLSlU8c3jrA3iGAn84Qpg
Kfw1fgmmLSe1SeI32VQ8WA8JOy+YzqqcODb7FujOAkdOqrGfYv7IoF6HUE6c
p97pwBJS4mVgKUdxNlAkrWp0vA85BS0KSqpP37464sMN44/KFASWQuFGKE7Q
1R4Lf3wlvEaRrKJyN4VJpk/oUq/EyVuyLetbsggS8iLySwr2N7WVdQt+JU+o
4FhfagoY8mDt0uyahlmqiguqUDNDgzb70RCy30eUZDV7OIDuZ+XCy421CnFB
+f+XmUi5zcx6bCtJYlshJdz1rQ/fLwmue6D8uqWFTUU9+YmF0SVB21LCIf8X
iEcHcQka7Nd8koH0l5B2lAvk+AwH15EdHsWiZ2BeWMjFzznxmtz3BrKgy0Vk
mZBp5R/+emu7hgmdmqmIRl3zuqJGiPRVT586aCJ4HiQ5z9GfB6vCVl8K8xmd
9Smw2yyfeFIfjhNvFdWbDO7/5bXwfLy8WWrW9PcTYN6qk31Zl2uf4hXd0/at
4A9k2atQNn+D9LVDxoXEkMf0zjF/dTXdo0Pea+11IqkhoGKv/HwLGUM3yK6q
MMmR9aN2lhnoYwRLvzURp/oLCZVaDXipL9tmORZkyvx2JVpjPHBLS49aIOYr
Dwybc+Nbr4HhqlAf53DavOy1/XWhftgYbuz3KZ97irOzz/RvBZzom1AGZClY
cielQST4pAKONKgl5H6MSrf9bYrZZkYPB04DSX3WknW2OEa9HYyFCQZBsHpe
0Z7mpFGxXPFCdX8JY3jaqu0e4wQxaSIU2PtIoAGvRjW7SO87nETkH3hVrXdW
y83ZAL5Q2nCcM4GVDGhyVjO1Jc9iwtYhVfDgrPLAIbU2TGzURTL6tF8F8Hcr
Lw76ihzwsaEr5Q77eShq7RQ5+zKo83pD2kPiSlIeIgM7kD3A0WFGps1FP91B
yKz1KMTdsvLAWQGO6dld4/BnbGLM2wpqgVL0/+TszL6V7BswbWeIzbgpraOH
h2Vifoc4WoRDJHy16rP/bt7XAHLzVvkztfHztcZgZ4iLe1TE+aKfOVH86cbJ
dAxl5+YdWDmO0ABJYgDiniJyzr0/VTsBgfQEokisa08N8HoCC+IXhRnGpbYY
rJz1roZ19z6lWyymSI2BSJp2lNIW2sjBD9Y0D0nh8cg6sfbZrHOL0AYk9lyG
VIhuoSSHkMC4kgRMrt8aWE93GUr+chYFeUX4F/hoVVXlBIj92gXg09TwDjAp
pKIxKx2f+WfewqC7BFT2wCAXh2Bl+YmdnzekZkfEZU+XUaS/s9470tmKfh4T
TjD+ypnxWrRVIqVXvzK+cPesEbjhrC4njZlkW6XtXw8q5dBL0f1g1HGw3iOx
1gbURYsySX4wn774X7Fs809qY/DIQX1R40nWi6qOx2Kz2+4Mhoh4knjhDZSV
thBfyFG9g90x681JWwoq1y/R6NaWv4vWoUH2ftT5JdBQO5zZ9+2mR8F89PHu
pdDN+P8LPpjYw9nL2cDxaI6nZP7vtZfwFYzYsHosZhd/2fj4j/tnHvXdgbiH
dgst/39xviNau1/sT3Q9IgHx8i9NmScMcphYokWQhp6uhti2kI0NnMdsPev+
EiExLWgtVBIKAr/1fwu3V0ro3U9VfQ9vjJmfXW6WMGJFdKlVl5d1or9Micfq
QHaBuo4VcJBsmWKswGx0GXwokIwzDLdaq4ph5ep5nJna2kUZIv0MJhmTxChs
VjLpP/aEA7qlDSAcaQH81XCAliSN86n4K+VMiagVBHrmsmRighXpZusce/9O
3//SMqjuUzFuQcypolKYt5637e0MlFmLTcOLGtv+Bv3RJCunIswqzeBIyh/l
8oO/A3NdspiTdsAKJkhxlXCgmoD2PeoZ1fxGvY/M3PjrjdKXRC84StYCHe1g
i+DeA97s7WmLigV60QUfolR0o8eLllSozCTgkr1cP1AhdsDzpFhNTZFKgT4v
yJcmCoqHjfCtpfoUUh0glwBbeCxJXSpzJ7t9ilsLicRhxEP9pTK99HBk9isO
6n1zXs91KvlAo0CGMeARjzJAHiKO2I8MNwzXdV9iRtlvYTL6G6totRC5FdRx
AECOk5qtvN1ugTRjt2m3KWC2w7MDbrQE1Rn/GxnzINca7Eqw8znGMLDaCoTZ
qETgmXpQosqxrySDyZfV7o5XhXQ1ATq9OOsRng/kCkufi6Bcj2wQzvdJDOD8
yw+l1w6KsVIYshjKbm7QbcsngKWRVkK9cKRNvftgaMfu/d3svxWJjC0klRe3
wZGObyJvRlt5i5AZy12lJohK+oRo5ISKbQFj1/In5l6j+T6bLXIG/Py9+IF6
JwGpb32di4Y6p1ML4PLAyflyzKbqRt2HTXG0Qo5rNYeD9bEiC48glj4jBt+H
bCqdj1+39BE137GGw5ExNzN1Siakv+LhICUkOQTty05UVDh7L11PdgHIjoTX
rdR6ciYtQNXgVftk7gvYK5eprTcdoX8pT6rpCkXAsFjMr20xX3l81NKXl29q
DAmbALHdxDFKj7kZ6mVaq6qYLgVBj+zyyqRI3Z8WEn0Cg0uejQ5n0aWf7wbq
BIdWoUpzln9JR6y8D81yn7qJCCs/pC+GmtMKTgOurhomGcU49KgX0hJ7E93Z
Q7pz8DLdMA5zajjsWFyB9MqKxCzC8sA7dG3dft34zjf07y//conEByGhMDSh
bfvvx+ESDOwgnjI6Qd7jD4QRPdTLIlJI34Z5U4zjKcgA9GC7pRiBUbSpEDQO
g2saOifqs7yD6/IjZerFm1W1nI21dpHurHOS9sBs3D7WudCsUjrLQyCLLPuT
i/bW4ZzOl+zloNNWwWlZwd1aUCOPKuuyzLMYkacdYtxlD3bZEAgUBQFPjRtw
h0nCQ+4JoI4iZeQzqM+HgTs3FvrxbJ9/gdcNdp/CrAceLqbeVYnjgmzbrp9X
aXSuPKPs36OMwBiBgaXRUhwx+fwIUlInfAec4PvGZg3NhK1z57RnbCjU4etF
luddPy4SLZTRCC1lXzjKYEE2HCk1ISv8tuag9V+TjQgr83BpjNmtXt6FGu/v
JCgvKj6W0dVCSjbNndbSMphSyH5IeUXZre1t+Mt8ekilfU6/u1GAASHuCcH4
wFHnmzpNnbpS/szQFVPMVXllt9BLSDTFDS+kBkilkJ5OY126e1Q1f/4Pcso8
AG2nshc83SHjTQK1NE+2dfg+u5pYPOhpmozlNToG4wmsEGyffGOH3uGx3uqw
VPrIZIWGInObE2HxbIGk1Z4TYgXsGN4TddF+YRHhOnpqzSRNfzgPqlnZRw8t
HUTfdO6TPdt8ujbNDfDBRFYY3dWuC9fHJOa6kxIaJj55Aq4yAc/4T2C3hYpU
PqYFb2/Wvi5nV+krvp/738ZJZIHiNugPzhyqTN6fBVGWL7oz82nz6AqNW4oi
l0eh4cmqDo9SMy9jsIMSm1cNLZE2QNzwmCt10xEOjRJTmKmqu+vixFvjmk1n
08H8jqjiE/v8+5VeIRFF1Qril1kR3y9dG19I7587rINsuwwF0z7HTe/vSuTm
9dZDX1+P4B0s8Ktczcj4ZvW85LWMpuHbcdTmnfQKcKarOxPwThYagKQUqvwY
JgHCMtpkPbyHTnQ/F2fGjsTMZ9OjsDNEnAUKClJCDXMNsAbR8Jp66e4zsjvY
P2Z6PJ3A/ZFNBV0iq9onmnoaXKVUjRNSYMSXz/LICHF1V32zwD2TPBDbXymN
SN8hc+NsUmt+TN1rlvAmQ0UXO5zL97Vih4trpFZFzPrX3ReOf5nFpwcpvV7f
X3N9fnuEaMaBseBpopGb9mkKu80irXMAbmg7gIWwwgQ1LeNLNeZUCe5jz28B
zNJI75xutY2OsmTIo5zy/hEvEEeusOuHqj+jobihWz3cV0cnR2JAuhGrERaa
9jDYrDLQkYXwgH67uT6gnV57IQwCuCniUiCSDIDNz2eVqSqf2JlESW+irNU1
DDLnYWQZv1EE3N82AOqgVsk66UjQtbSiUeMK1wvh62t1KxGJsEjA3gTqWcc/
H3hHhDdm3btx84lenXiYMiyFYbqApcZTVvApXQX1lRuNC7ct/FCmfA2z5aod
1f4hYhWCHu5ZTA8pD4DXk2qHxN2UqeCsrVjSZlS9nr7LCIU1xFRG2u4Pn/50
voPtieWjJTspwuUw3Rb+jkXTSvbzZDlV0VlfzgvhMOBUwLlh5kFvwXgsd8eb
6CGKqJ08eV0gaMl5ktW6hfg59WZhIA19/fjO/3y3GfFGwXulqirWX8J3ZBlw
x9UJeeL4yz5iBSRdJXDBhD/hR06DYqZEfGWMlUx2ZSBEefYnnP2Y8OcYhv49
n/18/UvMerD67ABmjk3716/nHG2RY9Wpep/AlAFdl/CB2B/aO1s1OuJekjzo
Qw9m6xpkt2iZ0+fmWkperXhAAGsK/ZJYczpUGx4EixXr+QwPZcHTpbxFsXDS
xrk/rbNMlsFzU1cN7kqc2r3kK5SqyLVdtLrSal/+h3qDzdZw9B6S3A5OJ8Un
SnL52Aw/5jiLSutix9uogzWaAe0SkMcuKh3zyQ1XXEdBTW1HkxgukQJLpSOn
8Bl0+gNGozUZ5PyoqOhs56zU193jMjBHul3/hawteGOL6BGI1FuRwKToGRCT
vZyEq7alCvBQo/w+d7fj0dDZ5TQKNVLEOAKQom7GZbmKaJlJqTdJ7hyXWv5Z
N6vKXkTH5PcNbCLbxCUjxeLAcCVg72F3g7hQ/Z6XWTxbcRiEnwlzeOO6aw7O
siVMIdJU3UHICruB96XiosEPc1sZ64fUHdgGsgajACLBRekoyncgr0WmBy/l
Y6GUc6IpUV4RXl7cbkSoJOYlI/F2yu61qf+DuTPh/IYeRqjy7xzCgs/aSsMT
gX+kQU3NU3yyENbDW3qDCPS8Rz8Nn1I//csymNpa6ncH9SF2UITk548kGhh4
B/TMubjE9DYGwTo6cG3+IlFu+arbIEdkA981JcMfP87DDf2blcb9EcXvTn36
333CMnXl55PKwX2khAt+eOKXCB0tJTYcMxSNQm8t5bqiibZtva72uKTExbyy
wqO6zSz45JqidU9+/9DLirNaAp1GN8Kl2/+Wxdmgga/1EitUpza4P2qHD/NV
Wv8IEwiusnbw0Y/ZJ510bchwOwSdVl1V8ZwjSud23Ht6G8GVxlu2+tU0qqxA
c2RPN68uU3XD2J4jEcM9jcwwXPsWpv49ad0oRwcb8JyA/POJjhnC/Kp7ZL9x
r9DwskSopfzZH4CPTobUvnmz7lwk96LkaK8iocOIx/BOEAalqtcxczrHfrU+
whY4NSDCUu3Vta0b0LhnDVmBv1U4g3lqFYsJg2ohlRzQd8a0qZXSjA10aO5D
n+2dfeYtBEj2UlmqQfCiAY+jiU8K1gC7nmR0QbMUOHS6Orxp+VDt/aLjMW//
9XmkYLcQTNW7kHHPQPyqJGVphW358tL4KU1kbEaYnvJ9K9q+8i2+gqIpY7b4
9I6BHklWAx7lk+tpTSUx2sw8MdSmM6H4CcIcgjVZnCAtzs1Auu8rKAntzDFV
tFgvTZGAbBZJr9PaQl6NArsKHB8gZlLezKnotWBGeMd2tUMCZsrsBDV4SB6z
mG+oCs8hYrhhL8cbjCiwsjbfFPnFeNucvpv3qnBKQBX1/SavyrI3nxvvlekG
LbJESZ0ud3XOflxydKjw9jrmdwCbM2SRFFC/geYdxpo1EjIcfP2M4vvQLEKK
yoWTrtnXrux/1P7Tj/JfkGIBZmytbgP+ls2eURV9JZ5pymetrnhzf2IL7W8I
+ZDXiVtzzdrm8kohTNTkFHWucIcoNBNwvhc6HGOpSJ0QlTI1lNolxs1cLo2S
4vzvarvnHzDP207mnXwk2XsjtFV5qEuBedOtw3rRDt3q8Cxf6NyrYyOZYFKL
GFeOfvsPoRzBCAYGlB8c4/hpruDOozPG7R3A50AH5GjPWUVZ10T4qJdFTxvh
KBpokYENCvZS+btjCmHVDXw4TShIpaRFNTpOq1q4wDtMnlSVBYyBRHrgDetO
ZbDWLUktymNQFqSNljbVneBgV3yG7muNampWcDdsPsLdxoVEHNwBv4wuK/I4
UGrPBga10u6CivT2QeWkvOU+JkxITrcyh2KBbP2MYS1wVuMKxvhZqzwgMVGW
zLXl3G/BZLI7InSP7NEDSsDGLPgg+CKhJ4Qw0zrEEZPQeypXoiV7lrXp8s9y
55b/SNWDlmtUL4/9xdelgHwbDy466xjuW/m5J6/62ut+wV6Z+LC1Re3utffA
W7KUOTrCHqmSCj78gc5EXYqJt2PVWRKajhm4p9mbsEX7IEl3kLWzyOmnhgyw
FdgQQxg8JjfTFA8eUHCo8vLZU9YTL6ZbeGKWPAIA9t+1gnmmF8RKEYxxEMFH
iHv3Os3JZwI4ayO4D2i5lDQoAsbaViwnesos5HlkhEIJQHHl3PmFiiURbblG
VGywj+HKcE62EiRsG0PWedOezi6E4T5FQHeG5+s6/aO9TF19yOqNnikSz4S8
/iAAjxo21jpp28H5aYt3R/A/qumMt7tVQr6aRWLycB/qT974Q+4N94KMo+ri
GK9tHZ7qOWaHnMSVAioi37UA8StuorSxVVh2ti6jkqiNHJlrAA1k3W+55txf
aQYtEFwEMnNhA6MxXfhCZAAhelkwAua6vNeQr9SMDdiWeEbbcEvRXzjRseiP
8FMJmqq4Rj+GYYlO9+WETEJqOSIZF36LwofqAR9EZxIlubK+C/lVaiVvjOA6
PQIEwlA0eiLdOeX/OTmdWKV64nmSP74B4irdPnTkr2rgkAhjs+p/gJkvjLWi
QScFpZpYUdKdNNZ3Q9swiKKVoaj9cJ/dVEj9d/vqNIFl5TGLui2C2DBdHmdh
lDkpUSsgmME4d61nR3jRehoaV/7m4Z+Gl116iOeAHTEcU4q33ZQUzDMuM9Wb
yhy1rYz9Xe+xw9zJNiZGpMZYwLMkBBhm4yPLKEpLVWVB5M+ru9+IAOwiSDJy
VBW9wxAxO50WnO5GrzJJWNfGKjm4qaDRcPZyrFwT883lCp6uW5Xm9M6dBzdv
z1SRb7kVqo21tGWHU6ZftOUS2IkMO/caY29w/8/l+igkr+7JECSbPk9zFc3B
hfKbtL6VjqpH01Y6xNtdozcJUHurYzVF/Ga4InRwvX9zjFoZPP1thgAWSJTo
cBh35+o1KyzO/bzUhpP5fnu40RAv6Y1Q4ZkdSeHT1avtahiQFZFuRtwvcFu6
NxSMl4mmS90jYAzaMzZLllqAQJp06zb376zQEnMVW7XoRuGJJUHRaQz2fs2J
7MuuxgcVItobhuGe8ZvuPn+nn6g7lSkYB7tY+E4K8uKFY6bV9oZKLbLn0fXs
kMogwjb2HyRwsJDzp0g0ol8CXKv4QP9O4k1RLqpDond4ki0qCLxnbnfS8Itc
QB13mSn1UneySggL46mm44SqbgLQUCj3YqOSB52VEmuFUn5PU96lzKwCBJYW
5SxHnDfszCqgsTI4zEv+ufT6sUi/TVQGYAwjGpcYmq98cKaLHETCSILyeFoa
KwIxrSz1pRKts9A4cxHfDGCB+ndTgM8746Trw1LU/G7XBi7vAam/QoA39RTT
dKKWDN+Qzw6yqgsj5cosvsRrmodYj3XkSlij4S5dzgNfI2+yiQLzDPtz2zqc
xrkwP+an3nQDjO5m9gy0iwiAFT/M5+cDkBYdk7ryfC7fsAcAqc5to4K4+pdQ
n66i6tPoUFGT4V19IJER7z2OuqzOyqdH/c6Ljse0px1me+Zflq6RERjcuRJQ
Qgr0JOB3dlIG6trbgJd26TMfrzQqdi9MG6XDpnDvgn6zKtTXisAVS62AAiud
xe6UVRob3I8JjKYKlCKmc9QC7hHTg/BqxbvI4UrgxpPegriDKvlzlEmnEtJq
ARDBabVTjIFufBVz2qp0MfVJtWnKwpBbWsBIjCOPPmYZ6zlwJZIzzlztpUuu
46pzVb+Oqtz1B9PRQvXhfg96tJ3eJSdCjK8pVi0TYJlFFgEXd2Jkv/BFuQcD
YEkvivjb1WgGMkURbutNS++OXSpK2vT9FCFJ7XDUJ9vb7hL/q49wF9koQl/y
dXpe3YIAgchIg61OjaO8ZhAwsUnII25s/BMKNwR8O70ds3wL4g+ewZeMhDgy
Wt/MizNFH5E2720M1p3v5YAUT40Db1YpLmdbbBf8bAhsmzaGR3IbPWs79y4k
bf7fej1yo2AiGSiSyrtbXKw1sqAe7Wt3tYZGvgWtl36wWqMf9qLRt3+vqrsk
3aQxrcE4B46VeyuyflzdG+OonbpsIPa6cwIBfxleB9AngJ0dWvGjBjjgVxeY
VIwurLbDdo6ldgwsr5ID2qDKum72OOTbZm+7yss1NImURhNlPILPIA/OipDM
voPSuvuvk4IymPID+/hJWSgcKqxb35Ga8qrsdXd4wLm2tc7XAVtwj3vMtvsF
8hkHIbj0Bl+EcrqII7ikeYBtVVYeuTk4FEvrptlJf7+hgBVaEmCrEVuc0O4f
tY92HYJAHH2Gcxy7qzMuBVdJYBUazOmty2zLBoZobWxOEV/l1WZN9rzeLvZP
mtA+S1rUnsNqIRq33+XwU1eE70Y3imXu8T2OgcIVVQF9guYH7LTy+oCfGc15
rLw7nnKOuC5cbs2tH10dQP5iAXnsjiO7QWJdHvCD0rzrHOCZkmA+Z6KjkWie
CN6amWYbgN2GNamIJincSHuKmlhLFB2LDGDM/TCu1at4YO9gIhFIf4SLnEA8
gWpfaRQrOQ/umm4np0PkDG4oDZYicrcVvznFJin9Dx/M1312eJEQduK4uHEF
52o7QPQg5EwPMdGZ48KMT7/qooAIc26QOQjlTnoZ5HawCRbTf1PSggUi1PvX
5E8ljmGe2K2v5eZ7h3Ue7xnZew5+m14DpvjYzJqXY27x8qqgu365wpeZa3Xf
voCEW1UN3sqwAo8J5jKzGBOy+WKiLbeXfR5UT6xhMidiDGZGYRgC6xc3kzjF
ZVJwNE7RuNIYrqqs3/6fCb4ZfKF5rOceVzwjPi7vqFeKrJksXTQCDhYqQyXw
mrFbMDC4/2h75Fy2e+nTC0bVShVS+hXlZZD4RbFbELTL8EDGEbWDTaxBcXIL
CXyEUEE81S/0uJ218dwE09zv32Vb+Y7slEEeJZYluxlzk8dcZTWYeyKTCzg2
vfossc80wOvr05ctrqBNAkeeGPicJP04MxY0Kx/KIN5/9cid0DVG/giIP4wc
8k0Z3B1lBnbB9Y+wetVsoEM+w9+uKGM1VfaFRsu2QvE4z4FH6lgRDuqw5do2
1QshavSWBUtEt8ecLaizC9JuhhMiON9nkOG9baeZS/pt2YAMY1dVlSBmrGTo
y3RXmSORZ57qCL8m2Z8FjolWC/PJIDDxFm/dlmOBw0HyQVANGncRoCbt1YnX
E3/yOHXsQgSaur3Q4rdbLUEzlXCBnrZ3kDxMAeygiRNKauPZYLbZYEGalL/z
SO9mNwP1BTJIB5neel1zr1fTGaRocXvuyq0h5qLr3CG1RHNyemhz6Ngtn6Sy
mmRJ6JT/f8vJRHbBTsAen05c+mldAqFeo0DI+Dcwnb9kGIW7D0U5LMDp9USn
rvv4f3sbbVGZDl1d8xSUPuuTcB/DXQBCxiO3qBXxwNNUA455+NJahpNQgUx0
OywHL6SLEHa8sMsu7QKEPv6nRtSQAoJpK5Mmfyes6fD1Xg2kV21/oQu4PLpr
36+OLd4ur7R3y141Gl3peb/Cs5zate7FGsIKx5aatuegjVApcn1HgQ6GxSw/
69BC70AAwCX86S59uqFEhcqZrXTbTWSpusLcrmqMe2o+iqJNvZNlO870kTRT
9bci7DFzThMTPP3XVPrPx0zafVWD9TRgMeCy8aS7RtiQJxA7jDm+olF1TIil
19axXLUWKPf5qOXOPt9xIBEqi1SmJc7eIi8huHfuvj9Se+edetJ1J4EDCX49
os2nRtCxNcNrB6E8Ge4yravDqZIOW5KQPGoYcbN9VZpIocxhuel6fld892XC
AYlgYQpOTmIhGSkOgv2j9d7XzrgXY6vQY3ipN5/wQqjDN8GXNqkFtRf/vF/Z
aejf4W8aiHRcqqvHug1vyYeDHSJ7ykUegKPEWJlDgWH1kNWrwBfRMKNYXFqt
c6CWImFGCuT/+dQXIP7nIqnfEKs/xzyECknUQogLyMGzSeXU4iulYOgKXF9B
3ya9RmJuYhcBSoCfnRUGSwQ+BK70K5rzKaIJEL4XtWjoNeOowXg3Iz/aQUaI
UhxT/H845Z+ZZsieqcyNG4LLQP4wfORerovI7Cr+ALKGm8islUuwWfgR1fX+
ORkZ72a2zIgiCu6vt2yHDb/h4UDXCN5XuM86DADRGVrXHFv+9DrSAIT57oKZ
HeyPyizqA2qNm/Z+cWgFt0caCLJl0XMd3mHkYFKHufTa1ABoKzfFX78XdJsC
dv6bqZt8vzQ943taM4Imi8gl5xo4yapd5M73O20PuaCcZj6Q+p2CZZWe43Le
rpKD4OzL40VczRMIqYyurYc2fNHnht4aztcmZrLTfqB1Rof6pRJE2+fGY6UL
pq0Od78z4t51QUjnxBuQuWzT0izkqYjtJ7QKT5waO/jOCej+kNdS3s4N7TcC
FCPeCe05LzfEaEpA4MQ+c0mJ4owj6Y6YNoTq7dqaTl1sjCv5HrsgSUdq8Vpk
sTavWLjM13dW8YeoB6wsf2MzRrApswfCowocKZY+QPEwN9h+u+G178Y60PEu
JHq5nmmdX1o50PrXz5NL+OOlxRiYOYZNwZW86RM8iCd/b/qQkRPZM3fUopq0
tvB7CHX97BG/hrLrK/adeeQP8UvaDQ+gbZgRf0oglNt5Z5WgzZXIXmJQU2GE
S+B6/Cal5kB3ZU50T6fa55lXtipH/xV2aPFS2qe5cG6Z8otHRabdwpiEfqnX
LALPSjSVBij/vyr7EJtpFGGWl0nWGfeO6X1+WeohiYcGtvvikKkgBZw3E7uL
GLPjUf6VVQAcXuBQV8mVSnS6e3RDQgKxPQWveXjU61jbtfvm+xqGLkNVSqQT
4gJ0xl9E6eFjeEJPrq6gQbZkmgFibJaHGoHQ6PcZ9qsLSBCNKX/YHpDxxZbG
/TcO+njCJGeS4ELvf+AtgQp1Dzgjbh8sA8qRenO/39nQi3+23VUlWP0tXLbD
0+47G5eFG+g9kj7H7knwAoxQO/MyW7krGYuDioRBpg9zPFKbECTNS1Y8fNeH
k3LwU28BTTL+hR57wjmN8I9xIWwHLQPBNZzvepfS2HCRZY4622MwbpFB50Uy
wFzNGscOe6M4CMrfFR1AKVW862qCcHmD1zQP4k0glc4UT3OMSs9Q62BVEPwY
XeBeY0JWfXLlohxtGYeMncYDwd9jDL9dzIu/PlVG2TFJgH3wUbEB6qoiSRJJ
3MrXfA4Wt4dV8nFodgFFlHbrVqkoZHCnx9Wws0Zu++JM/J6fc4ZSGUYu2dIu
IBrvnWI1LHtTOy9yLWVA8pqSY7pxufjwQfMERisa6CvqoDQxpBmK+Yi9JBPD
PaFGMU9Hn7OLDip7QZ8gU+x1YbpNRxa/QJOKZo+1IWcyJH6H/QS/UNKFTzT2
mfTa1G7lShhhOdEy+MsvTt450SMI4X8LN1Temv8LZS/jlItmjsgd58Url8jF
kwq1Bn/FmE6q4vxoOLtoEmRn10FDqpnd1/0dLYNYByzl0RHwoflDLGKBvX9o
6Vaylwckb/6+acIoKkUQ1BUf0GDnEr//XwTuAKWGNlSmCqvqg8E5umiecpkI
4DmmxP21/lbmaNmY+K0QirRP69uVAIn4L2QDNOKtv35n1nVgb5bbOxvrKp/g
C4h9wvQCtZSbnXFV8Xfr5dv7FB4vfUFb7VW6AhvuRgLo6bdkX5GWnHS0tb1J
I2RYF9jmzPHsqgIzUYQ0CB3Q7fzFanXW+suTTXeb109bQ4ahF7RIUL/1cvhk
F+oRDirctYmxXMK9fCIvHzMUAebxJBG4NRtXYURWjDKhRXKxDLUUYiV+ztZP
Qi6dUqNChfUWVQm+uKaP9LV/P9WdxpN0qJOK0gRLTh1Ey9Ki1YH4NagVivTT
2xCb5NHfjgu8Wuuh+kqGc+h5bcSNnH+dmzhy4Zptygh2HOcOQa1sytk+/eo2
vOOe+VMC6avNSHs9UF37xXNlTB9k244HzGt9ApMIJAlxKVYwDRWwg1mTLJrt
ToSsiq5ftFjNce5CwDr2f67i1TpT424V18E54lzf+oVsgyPxBuXC0mIc5vD9
tg514xfC3Z3kb4++sxRlpBWxg+FWN9ZeUlKznW/20VwGpl2e843LCWfEVaef
SDiQhxDagAamVPxohSqgq8sTraLREnGEPptkPosogNv8HlRQkdf/d0RmVhx6
EUJQRbPI4a6bJsUcyZ9mWa6UoItRKJ535F4FiyGkgpO3qdm/RB9nf04nUZGM
JQ5F8kZzOooWIZkP+LrDELeVWB8XVkPJzPWoBzVHAlJALy8+K0IIBAUar1aN
XOCBDFXBvp3JAK3LUluWZ8VH8MIkzQ5jrTg/W4XH0eSvkEfdJ2LBlRo3qWaT
Lq340no7a0Yp8IViCknCvRyDaT8w5BxrSkESqjVxWkSSSK1Y0h0Ty5tnPT/G
bRhkn9Jn+pEFbMn23Oewx0Xu+t0ce7BWXkBAD8wAoeA2bgAX6M/4N55iEE77
5A+aCXFN7gwd56aY++746sVBoZlOllBDuLU19TRywxr0ePb3m/7rfDrSQ/Tm
DERhAr5zHIJ7wHsTv3g2Jt45BBGObOZ0rZuTRsdb5gvj/2CGBRIaGvb9URKN
P6oJEpBfQQZILdjieiLldJUdL7FDRHXpYqlnxwB7oyMLFliC46bC3CoCb0fe
0SzTO0zxPJ7AGrJ+Sf6c2V1ltv9/36RbNZhGpF8bjJIH85I+oTQXkKaEW2ag
Tmoy7J9tjkwHvhEwgXpww2jfg69YUszTSS1SctuJrKtnE0u7I1buCP0jf1iJ
wz3/vFSttiMfFNxQpdVJx68Lj640a5tysgkCUjpf7iIufHcP+Y6xXxWPmFtt
BexQr2pND59KsT9ZmLRK6ENQzgGa/GCbbJqwVWaE7BDUC3/hTr3cLs8Vn64t
pd63iKm4vL1la+Upe48vY+kMjlcoflesDEbUHZQMQ/72IuituA8p237s3CBf
dfCS+9/YiQJfRa/S5wPhrvvofU/iVUEpYq5djsBtNvyHy46CiM4CZpKHrlx4
K3ZWA8IMVC34c3PTAp6gMA1nQ1clBf/9kuyPTh/LnD8QQ1lCzPq6SKBiMgdr
4lH5DBh1gWmShzlWDEEQHS90xfAJ1frvat/waT3WoFDLSZDLwH7QRJupo7Ua
s21F9CzwwRuiI7G4/rjYaKlgTHMY5ccdjIzRBKdktwc5gqPg5gDOGmUYRSPn
KX4dFCdRuvqFk5I94aQfbrizmMJ+yaDaJWIV8DsqgNPe6FGtP3NajBU5ca7T
VJNhaWeEnx1zyQCb/nja83Osq0ZWUXv+/aRiTPASGcc4cUOz9w68W5VMBiYx
QauA6/LA30f4EIRxnlKifKOCcpTJvkil+vWsZPL0YfAaG6b6hBilHJse9b2y
b8+yAMTxKzSfr3ph7IPpomD4x9XLxKAXMSmDy/f3Iww8/SWL4hJPq+9O7rbJ
w5vVwD6uFQ5gBTxZu9MxmsC9/iW6u65HPtVVa8GPG6zMIGsbDp6WkJT9v954
AcvEvqTficg++4ghlEopWkpIHFYmsnVDjMoYmsOjPqC2175zbYb27LzFLJTB
6uYEEdCGODeelJ4lP+LHL56CaPlsuyLw5k3IA6bnUSWO3CJHJcBduNKiBXnn
ZJ2nyXXHs6CCO3U/ez0YLb6N92J/29ZFl5UPPw6XzC8MKQy68gDDJ0ihju/I
zhIaGc0pmnlw0RHRVMEGi9YO1oxBo8TLwv59EykVbadeIcBbvpeg9sG7pa95
0Thcb+5oyZjA9gQGr5/XNdXGOfuFwX7183Dm9z1PlgpTVrx35AAVzt47f9eI
h7TenEMt2HR6fK3S9+vGVBeKFiNDeBrEsCY526tBVtYWUznNVr5TZDkjW6bh
t3T2f3SHJvjf5c4kRh3ueivUXSTU7jFW2lSTN/Y6HVhyim8YGj9zDoVqkLyQ
NxVLbsn/NMPCrIOaoO5gNg/651UzlcGw2KnwiiKnsbKJPNqwd4G1k3xe4fTz
OqbQaL5O2ZIr0dZ2Bjg0sYcFu4JmbojFuTXOroY10msuLOED2j8I+8dbKNq9
61Q9ddfjBmBSESI8AnJXCHjK0JZv2SN7xD9bEtoVCxFgNmOqHFc63inrtuZk
9DQb2WprYgO6I7DBBLjzww5kQiv1fFdF8xSchN5JfmeEI2tIpVWa9/Fxd2Uv
RlMXBjdW1PukoXHhGnroHFVvgrwEw9uFGio5kqbFCpE4nwh5qYQOTJYJ+QwL
mHYQIc1xUxCfSoEbPtN4FnvK6TvLjX+9/Df6GLdnxisEzK3sP3W7azkpFrFU
cteDxA6/6bramGF9IGapINBAmdbsDJ5T4zjzbEl/3B9zYg93CmSYcfX+G5vM
aSniRexCGzaGgaqxXZDQcqlKi8R3AKd8UVTpxsLE2lqy/0zaNEOlxc7D/iB6
BCyGBEiuAXiib2B2O5x2q8cVpwgMyqreGd6Da49uLxpla+GuW2A71PrOE3zb
5sxcZg3Rtpib9OTNTBn2RDuFp56NhGh+hwSbCIblaJnBHjoegKtbfbP/erZy
whs76T0aKLqlM7ey9xHuCw+ihlEmyMNmWumiVtV0hEmxzK25N6d/DRFACGEy
uCttjSCrpGHaX015z9/WmBzPvcaJpIRBdTM9LGSOr5oLZNqottUT23uFQR7+
9wvST47Rw7480liPVKYTKPlQF0nOOqdVV7HRPnX2R4W9RqkUFngs+sO+hqHe
gSeeCyDfYJRxj1qVqT1h6PCB+toqDv+lTU2qw7T1Rn+0V243FNaBeLOhuBVU
3CFEYbEPuJD255HFrKdfhMG/7E9VLerYYXopB/RHsluQfWP6oMQasvOcFaHj
DB8Pr0UCi2NV7FJ2vLUOzf5c0u0/J5LrYwjt6rczQwDzrS3I5+mfupWJsdFz
1yri5MQZpsz3WBL3AQmavyZI2Nwzc00Gi9AKRefV+hotD87ofdFYac/gXk66
xK9S3PzvZo7SvGhGAz8SoZ/0r8M9iTCi7Xw7TnvKafyEZfxiHhuWrbGl8zzG
zYn+XYVtfoKld8Sy/Jf1fm2mSmNlRq1my1g4QgymdQ9h0JqjVZX98heHDZ6F
oYOqqHfUiD4b4Kj2tF6CYA8IQ6xe/05DVxnjYJfxc1IVaNnWVyAE8At1eQ6p
kSGPia2Owo834ywvcLe/hoW9aHZWK3k/7G6K49BDN0h5GYFYoGzbkg0i3RAa
AxBcwOPxxLdoKCJm1REj5RbjT9Jqog29Ujtw53kYvKUGgUpT+/BAozoHSiWr
eUqpp9yb2eTnfuRIs/mWW0Isgpyqtu101GO812k38+WR+uNTMtV1ufRkmaOS
fk3CjEtuLG0chmh5af3hIWMF5MQhEtEvxAouXsxi17UopyhFiEtnxPAtP/aM
Ekwat+/7WovtoYIhRDAFyAmm4R6rYdbJ7Dg5kDsQFMN5oYt1q0cu/tpFxvXB
vKQwKyCPWlJM/RQW+tRhawxFsJrB30wCjsBmIImZfA678Uj+jde7aerLV9RA
miurubFY2Ivyox91biM+LsH3zsp4AbdYeuCe+9CXKc8bSekPkB6WZ2YBI5cJ
bhstlmUq1IB/6YIfUH+YcesUbtPEyfrO4Valx9MayPRbRKsG5UUJWGRwzw5w
DwIeqjy13YaKQGIRN38giySZYf1GV/WKVW1QxG22VDGJ/bWAitMVbasHP3Ee
leQEfiH9oljY916iUhSy8Nsd+nteyROdwxuCLAb0IFPyg+er9nElIWqZqgmc
QWqeGvhWuCCv3fM6g0s7lYpa0flmxfEJDubcmVBjObgQsVF4FsFT2lXj22wm
+11S9/GytMVQ/LiOUshewFP925Fll3t6UQccKTwvRTTyGDrE65A2qkLJhlUy
8ws+RjJm+5LD19yHG/GtgupW4Wo8cGxvyCkL0GwZfGGE5LvX2rfZNjyS/bw0
nzZor4WO1c4M/21JpZNTWKdUC0BBjUCKCVqaUwNLEZ+gi/tkANOIPsgSKG0I
WEEe8aMnWpuUZNB9lFevok8cnNI2uJSGGfD8WECRLf+9QKQpRyq5jamPnrqK
haYePOmvGwEltTx5STsunErgHcaGd0P3DU4Y3IGquFW0rXEME1z+KlY5rrmT
sTvD5Sk+EDnUjYEWgUbGbi5cxOtHN4Ap6dYQuBb0GRljq0z7MrAoovoOqz/M
6XcxS47SuFZlkJgqHgCV1YxegEJErCnnowp4SKWHbcKI1Kjy+Q08GgnuLiDo
TkyWQ1EDhw4Xt4vPK3E3hLYMJ3J+9iuFBcwhnGvu02McdU3L+q32bB6pQ4Fo
Mc4i74zi3wcSWSrw5Yf4RrkxIgYHhyUgE5FOBr87injUHo168iUQThcHWe4f
54nQufP4aKH7bmuujH3+VJ9gcEaCC3ZfTTfTX7AEbPaXVpPFhbg21wESHk+8
xfcxnQy7AVqGKB22SFfPwQZoTe9cpLFLJNpMekmD9Uts4HhrmfIZQfknnLIS
o4PVprHXRQW8v/q/TxhoGN9Fg9fSlOo0HxaI2JmNana3neFC4qTufpyfioaa
PCwSl+nIgseOrzY6rIAFAD3oVPH87IYrLMTiT5MPRTBal3utb9OyuCc4VmAU
aMXppXhlEVhySMW/488d9ZCSlIkNqWztuM1hlbvI0qgZwQ2zM6Y/bE5KAre5
O460TYQgUR3AkPyQfdOKb6LubIbZmzWYbPNNm9dd8PdDuJ6dp6dMKKMl4iPR
jtyFNucfm75YmlHo9hb3AYfseXnvEUdbXGlWOCCv0L2s/s/ZeZMVuNcVa0rS
9a9MoNUE6kS8mpc4sQPEoReVoLKcDTk4LMdxafMQUspYk1nEemSHRLhEjNd3
0FJdtFVg801/i7trE22vpUgSlfBuiM43cr6fviWM9CRx5vo8FSV62blBl6pl
rzjfBRwYFYQgM5VbebKO8nE5AgzVFhf8RYPwLUOq2OEbOhY2Pld4rMw/C5BX
v+V2ufLWLGatuMvWBSA3BqFr9mlXYs8dMpIInHKZLCRS/NSrzyAJ/wtsmfNY
5FUOJhKfrQkVwhrEEI96AyCV6ttx0W5AwH0ODx9VCkswNgpH0AQgUtyzxZ9F
nYcxmqDfDnpQpxx1L/UeI4LP3qc0x172fSXIJXBk7tbOi7AEqvBUm/1DBl4j
WdCGxTHeKLQp+zKA6hB46JLytkEpOu5ID7lKvEdxJJRSVce7sGaNvSsX42Tv
JipAy8PfqgWkdHaksTtdMjuvnia0UBjiYF/AvRqFq7miII6xZ8d5FZHmzIpV
Ddo8SMkdUCpPyK0h2z2F+j4Z4vEwLOyzdNZOvJEAqEQV2tXlA/Z+W8H2GpZG
93w97LflkCxIo1zKFnJ5nUPmjsfYYW1ndF4y7rHzqqKTS4zgIw6mSS576shR
QoUblPkWeAM4IrbxIJAkaRWgDo7lC4noPGWqSR51/TVSMVl1m8VzKimFllb4
neFFnbRFuvMpM/UliF9Rcb29jkIg7I9y5UB+/C3E6s+yrHHxs+fTVkjigRnI
pf02q0g/hd3GB9VdcMKkT/ZMSRxxRJcLUZ5N8YkfnHE5U/uta0JFlvJ+b0UH
q0oGTcS0avT0pBdC1LZawjKACjBTp7u+xh4aDNaDDKzlWXgNkQB5fyn6fH5c
+zWzq1Bidou67zzjjlZQ7PAX5iMslffaequZZFfCRzE2FJpEbspxR1bTnEJX
LEr7Nx+upei802k3TJ+eNBgSHv06uM8pv8nhvxtPwUt9G6LqFWBK0rwq6Nf2
WGBYmsysIjYqRaTIVbNdrdFT7evZ7m/N0NKg0dSvsNCdCSNZMpac5S3xGyvI
hp9zJ+rIVT5J1h73ID20Y0ZSOTje8nMRnJrhrUuO142feSrQu2Yk9xacYRBt
LVW6M+h8T382IVJdvj7dbFYpY2vvwmE7PwjXdtuJRo8V/JyE0LbSIvNwnoQV
NeLy4aJ2sAE3sVmksj3LwtL2LfidXah3GAFw9pIvBqBKWnJ8FMzSCBdxxEvv
6ORBcbfrJ85zvY3LB3n8k5UzO/z1cUpdvsIXwYEfJCPvi55RsnziUBja9pkP
kMbZmKDAW4DmrWlPU2KuXtAklR9trq42ojX2NHcwoMna2EoepVDuu5fg6TmG
Au85+YNLCd7HzpMsNKPHjozXHKRdtQn8OX9TJV9Pfl44kIkFfjQtI9y6C3El
eoLhuYTyxFZXz078c7XbunlSdaaUqehAVwaxsnrPAiaXWqa2RadeVZaXUHhX
8M8P7RUO8yRfVpWt5k6QPty0lSuVJTmR7Dj6tsN3i01RISrmU1yZUn2UkQ2S
jvYDnzyqeL+pI3YmTydhaLtC8kWYbo/jFrGZHtfiGkFd/oAS59x9i2puE4Nv
xgnTbggEKWBYzIRkAwRsMu4gs2k63Q52iMHvKJ6bsCLJh3nG71RyRcuYHUBW
36R5YznbdLkA9pjQHzL/CG9r9cqo/xDSA7YYZ8ooITn7m44GXKozIgZ7fXmH
rb0aO1cf+xjpnb+qlSaYuSEtsQXccEAteElUHmveoK7CfFg9DIg74clUkydQ
/BlyTsIQYvRNr5EgNidgT29BUV7Evl9gAUz/UnDtLR5H8Ye0IY+SnRybuksk
bLMAwk65f4dV2d7RSxfJ0B1eMG/Djeup9jbBohtbsGuJqmq+aTtsCjiWE0WO
vrel+Ml4npy19AHnJBzsdrTG8W5Q+BGNUmR2JlCGnY5gLw+2fvxEK007OrYN
28M78K+sEf8Y5rXPgu9mRtFzQp5iihH9RbgADUDyGFgdYzIl1hVp+gltP/ZO
ck8XQW9RbyVzHqLpfXsK/59hB4kyNQMH7+yyL1Pz6iLKcBQ2ApVJv1KY055L
pTMgYEjhiciYtJ997FC3Glg9oomkzMUz4HhUYvnOZkzqRf7ziQdJ5cwtpXiS
O7xflZjg4IZ474lJkr11jguUmMTgBOUX6XDi+F2obt9mGAkWIo9c4PrNSH1n
aNfz4ycCXVmBOEb2W9lpGo9yprAeN7IqHl3ujOEA0NdOp8mbAn6lGYHfpIbN
F9TPAMmBIuL41hSrhUEjgYQ0w3uXF/dahZMSOfip42xNq0mBqVXGnSI1L9C+
fN3yZrGoawU2UJG8AhhOnuOFMzSq/TkZ62KQyjmsJ/98svym8OJ3ZKlYCEiF
rXzG5NwJ7YQegUNdXL3HESps2EzEx7OxcOtz3aG+poNqaqarXHLkC3iIMOSA
kOaMZvw8gRwkZ3Roqyl4I8mIzwX/wLuwHoaXsiggiMg92MNT5X9D/ZGATDIU
YyznTyCzTvAYdeJqigGdKLsQmDMi5xuHm2P0ZyPUhKgjbecY6u8rv0rbnDl3
YWwyFQ/+8+xGSZuxXW1ovNpewBypZrnOfobl4ykuIJOtNOTnajomPqsL+z1z
qwKCTBZB/5h8BfZ8WwBhK4piiBvW3FecYkqChuGAfQjhqYefDAn+eOGApX43
KMD6Orpl5CWXII0J3XykHVnFjnR3i6ODiUCyxIYPXQ490zngJvI51uGiwbsg
DPZeVXcrq/8pgPHngcxa1n2Yw8SPg0keCZ3dahDqj1WehyI7m+Fb0HuNSuu3
Tob32HpGw2Sa5nk6SpUSukxDt1yUe02DtIbldQK2LfuQYCvtW284Zbew9RvD
jYQtleH6/0AMjEXZn249EYHnD5TFWhx5/6xGwR35uGav1xfFdQWEzXVGvbLs
qADF+Bkq6EGidqx46PXdw6uoSeUCP/isndBodi2qk0uElujaW6fLy4rWG7YM
CZMtmzeYv5HPUkExFAf7DEBqAPKgej/zNAxZFiPbG8PHUjvcuEAqOLCNBOn0
mAIHHQND8mdHod6IE5JA8RSxqQ/ojLflH7U16hiMi2PllH+3i5/Z4QbgQGKg
7OTtBf8euWVjkESorB449NDbTviG3VamxiBOXajGypKtffLfKhb9PAlyzD7t
1R7N2WBoz7AjXFml+GRYyOGNS5TYmPjUD14zYINcDkVIidrn9UgMr9Jofu5k
HLHBq5IzMRzLlewchSWn0H46J7Tc6ucY2xmIj7USiioaJH2NkenrUeMvPcmQ
QIcW6lJeRY2cDb+NLUg6LPgFiJLXn60IJaWg0jVTY0uoAh6dAlhTUw4M4kXS
eOCkUcmBFhGOQ7VrEG41eENTsPeCgZUkVEljwm/NopUxmsvO3uEaRNGV9K39
eLZiNeblRw1rqU9UrWpsMAPbc9gF0TY8aKd9dneBhNYf7Y1OgFoMf3hi6wu5
QAEhTzvc+xa0SLAGwx8IC9QSZ+HQW2l51wFzB5krq1DK03YSU33p2BynR8Th
ulyb9AG0EaFy34gZFVI0DkkWiKWkwWC/DSieJiDt9Vvu/dimLigLnPnWTVSm
9zsT9593kSt0Gz8186U1b4JZp79CT59eDiCKk7Zz9JjxBQZZRMPlgOSjUgIN
SyEIzJA5QzMpSeHQX+heSbnBq0ChhFwjABI0b8wLcDzXlCSfSUNQLnhKi8mw
9oM7TQ6+eEajwaO7JxHsi6rjSlc/k7Bdaf534SD3cPkhveKjgo+a2hrRkt45
fN85erOH8h9sDBqw31wcJfyU7UgM42a9JD9IVb0MU/3knGSfwTPKOeiLDC/C
rrKoGgYRXweCWN512BZaJgKzK/RRphR1WVK3kynawCncME1byEI10neovDPo
HOZNN/i07A9F5M+NhybRnddGUxOHe04jMoDDjeHJp9TrRZWyr0P0Np7SaM9f
BfE9uxck+Kwpf5CTcFUE1VMxqy/C5GCY3miMyVkjqkTZyZAnJtkQbc/Hwr6Q
s5dx2uVORghY8axFp2cr+KznAA8m8p5rHSxYCnwCJoEOEJgpA3Wz2Ou24n9N
nkXa5YniO7iqOaC3s7szXPKYlZNN4DHAgBzNNnQCDPOxI5gPbZaW/xYBhv2Z
zTU8uEr8vCEiT2SrjN+CX3LqDZ55ZAtr1L49tCz/TmYHbyamrbkqsRTQWaFv
7yik+ebS1LatTqsKCS3b2/cVDWDeKxNqyY5XGtLvgtjDmNceHWohyeefIu7i
pSn5CaOVlWL4dq8U+hCM5y6RCQD/BgI/O+3WWrzi6V2DDQxzUQ0kKhWdRuCK
ieCAPghLq5NUEldVOlS3nX0s/x0OTcimJwlSGufZWvV3i7NIY2D2NF4QZDLw
6PhYX3Cx/isS4tlr80WseiGmhQSVfUQUPck2EWT50N2ETR1FuNmIQwk9CqKl
UKmOWVIKdgNsjKT9SzNL+3l3R+bNADh2iuCnXCQToZIthUPJVxscaa60YUbq
CThiyidgcNIriigLmxNyLaOl5hGusS5snZ3EawiE/qs4YrH8OgC5mMj0EWk/
9N1Wya7scmVegSdktSSZ4UymfMW0P17womCf4xlI6V+hSY5VMkDKbicXABXw
+BV96j0ylmGSzjJd0XY6OKWzbYDC4iBlA2TTYk3SGucwjSBLKfQsQ5JWQpbY
k45XSlC74yRdGjar9OmbFzPoG4KkThPSt16c3YyfmmVkFwsQYcK153NHqVEE
vdbK3Euic58mIo6vQtrXbGMvV8Bp01vZKTNm+iiUSSM65eGdImGROWa2mCYJ
gKCRjMriVjZ3QZuh8781NgIyr+yqTIJS5pwfVIpHbgNlMTv4Xikd/gYnNS9U
n5EX349JCisuxDTUgJY4FgGnMylUOxfI96zJZ306CGGLTJFfL4cG7SOM+Rco
/L3NwbNv16oAOXhFJmXpKV47VnyafoLjAlrJdiFe5Ywkgs4QiGA+xsQ4w457
uJe/L6DJxK19xotDMQ20LE5PanxSyOZjIHoQtud/Pvl9awENyY4YwdZ8NOoU
LoCzoA4hxRAToVPTfLNiycCz9UIo+LuiuRsytp2QFWeZ6PeLI/yS7fj7SJAf
xWwLqgzO+qyVboWiD93vHUQXVESqHJqIn4tCmxn4iQli5caoaJX5lZ+En275
4enhjxf0+4OfQnWRTMwmrz+mTBGNq+J7noWNcKS8eFqQtGWNVAGIyt+PFlh7
nj7yOGkM9DHOHRdjXAFHlu6+MAtp55AS9WLm4Y+ZM9gVzhmotExWYEHruwSp
w0HcYsMriiNVCkVX8VQwDkoTKhzS4cDTl0L7E8k8LMinqUheqJpmPE5VrT3y
SVMLNXPi79L7YrmhoYrT7smdAEUJENrsvsBhMzYYyNZlmERTZphjUVwQXB7y
G/1zF0W8TOIIUVfCfPO4Y5jHw20mj2BCLTULQ9d0FsnwvGxCpeMAza4VuYPX
QiummONjzmF5mZ6lA4RmwbhKFKALN4vmoBV7q6Bhkk5nGlxhfhC6CqPeDkTo
9Y76exeH3i5yVdJ/fmsR+yDd+G0NWolsPzZVN8v3r3+XYWHbeBC0oCSuuRb1
IT/xez10VQ7AnyV1UK7DZPw07qHdiJqakSEpVpIUkhkp94SLLed0tilh7nHW
Ac6QvVP1gL0BWPm7GUaIhStmwZwZ+6ibQTC2iUPu9BuUrx6Spa110wL3N1vH
DSb3h+f1ZWzae05n0RVEwfRlOU6atlteMSgyMbOttTu/NSPz1Hm7oNGY6/fL
3GjYjmvHEqy8sGtv8RfyTQbbEekFSZCeFVEeJeVyo9uq8NX/sD0njwUEczJ0
GDb9UZZuFEJL1K6HHYG4CgwQhUORdAOh+Rt8jBKRYjx8neC82WYXRlbzWON3
UVrvQALO2bopaWENNTXoVmCiwuZoiQO3MqHePzfEH2a037+fDcl1GO4W5BZm
2s1dbN5Dq5UJI2evW1mru0hS4dkcqVxnKN5P+KU3fSKxPrPtuL/w4tCEQ8sQ
1OCzy6DgHRr2hkQBJJ2ek5nZSCuCfCWXsRurnSNCbgOTiNY18JOQR7iLsOIQ
zEfltUpfimKCNhLJ0mXXXEOhz+qD5KT3Ke/T7GYzXRcFmo8NhaP14evbwz+m
keq9kkfeHTsjSWJtYcnH5FITp3K5xlLkv+wJ12nkZX1R1FAo90mBDyg3KH4W
7CQsI3s8xg4BmDg18RTuTiYpKSxNH61JzEU8wO7IVd8iUt6D3Br/w92+IYqZ
R8k2IcBmK1B77UwJTiWlBc3l8EzXpvi1b6EST8Gc9LAL4k8WH7pmRUzJfxS3
tyT8hEeGGYgp6ev+J6vCHeVAnGvP0d7gUov8rcK40PuGkY7uHlPdL1snxcsz
gMAhutpPzspMUCuXWdatr+LZs+qKIOevNI9C0UOtHPrPHJiNF21QVJDf0LG5
taWVAfdegV4TklCPV8OOXVbfDi8xGFCWXDPSn5pwHbHqo5eH5qU1j+VQ2hsb
Gdi2QAhB2cQSthcXKjzpsMErn/A5WYVHeQXOqmJLI7x/4Mlq6ObA/v6/8tVr
r1ro7MtGEjoHIUwK+CNVa4HY0KN8pWBtfJLaRdlB+hOOgkmF9+RQkgwPGVYj
7eobmNYB84wkgXbMB6f2va8NiErrLNUs7paSO3qyxtMkn9w4G3jdWg0qO9oK
KhblZW0LQwxNvhp9lRlnQ4+mxX+4zRZV9SBU+EOkO7LPqPJkCXzpO6tyBkVc
KW/GKpGDUiW7kWmkefROV7ZpkCKg/M59ZAR0vIXaqhPvv/hj/IeSULsl1uzj
xP85D1n93aScncIhK+q/jwpNbITqkDPokjmxneXyFd3+pv+kSQWrrpqJu7jc
kwJnFZGgKktGy38ZNfLSyLxLoy6LwenQ6PPeYVsesniuthrGsAXaOWqGph2M
TZ0m/dabW6XVd4VOlGKZdAp3uuFDFjCNGHl6rAsMZ6OmxOZvUbawYpip+Sur
n4PdyEqzmm0SPnpmlJQElTnPld380ItoTfcarFKgGXtAKBz6s5g2bEjfFXLH
wbADmiQVJxNcF3x5YRxny8SfLCvxSdaKPvnAc/mSm6ZYO//QR8NoANyVz6dV
e16VFmkY1w28Yon6OL6LRlMpewX6o3a4TyzewePV3IpocTRRVvABkag8lFg8
ILiY0rznCVphQZe1hhD9SQK0J1/Hk00Iyno683Zj0tQz5xI1WsWDlsVHqqIJ
aQe8RgFWh3jILBX9n3/xkxx/CR8Hr908Q+9BniV91yZ+YjrgFObSaFUqgqwT
R8NMCLJxyTofMP88PBMfaOPlPhy0SJewNIhb5JI6NiZGmws5Kapk8PtntZ8X
jf+zo47Ceh0FeeolON913F9wHMVwXBP84csBwGF7NZlr5vtXUgIpsp3ZcjeE
oP8O14D6cawqtd14Dyr46svjBEU6/c/kV9NKj5zpbe8KBk3wXrXrxdOCGCEX
ZxIZLxizOJv38Ri/UFG61gMewYYoa/PMsdS/HLVkT1uXdQ7W4zGWlpFW95WZ
dTYEoieiF7bae0vmoNw0jymqc82jtWW7FqPaZIr1FFyBsfrg745S8e/TRxxC
rtiiBfj1FELS0Y/2RjILVVmots36zHQ92ikTdS0PS71pbSBn5r0eYE6pHoqt
bN2LYoLE2GDId+nKJisFZmdFBy8XRadDj6fVnHhHCMM4/9ilaPSYwIE4L6uy
KVNGBxBo93Qr3SUhX7UcftQfGUxRArW0hINxN8PafuCVD47plMP2kA2m6oqL
jE8yVMsigvq44BiibMSDD7b5337H4eM0xoq2rgzIyOdYF4vcX5sDMT8H5EUZ
J5KHOk22S8xhPGGILW4tTtYFYvQRh+dD18UWA5RkL/rK4c2iroy/rKgft4Bx
maeCjQB0hES22QTqQSX/s3e9VCgtaAXNci+bSQg6vusfFpBDibBy+/tJBHlW
iwdhXA5Hz9e37zTU29bpPCI0nRfHFMCazoBrpjFFXmsgsOkwXDaSyFwOsc3X
sCjehtxltlghcgsGjAIGBytHyECUpgC25YoUK2APLXI5piLByMSlXaUpJ6st
P3yRf4sQNTpLrNF21nr2HE7v1IK2KV7I7EaNcsm92IUfDEPdi6mNQLeROqMF
ZALOHZ6CpYZMl0to+6n8h+Szb9qgqJAjCxG3LP2ORxmoBtg7GNyP76Ucw80c
34g05xXk9ck99kXCRsklAsQO6gZmEi884VIX1RhVucjOQOwxtxgJBH1i+3Co
i5Gb3jK4JlykKvAp7NhBQIGR6sTcuvMB6HQzSvPD4DGbfFj2Ri5HNv8ddpy5
JBY3uk0ciQnCo4EpQa5JbarV5XDOPjIZJTIl22/NDzqilwSzXb4h2qB35kLW
NW2c50YpYNNeonEppT+ojpCjmbnwzsuUMJak3KcniDxO6WjaOADDaG8OxOpY
TAzEjrTaPOBEO96G3uRhQOpKZeOHEqna/9WoFwwI8DzrPLKCg7oNqL0TqlX2
M1sW8xlO/B+Jr0L8qdoX0YQppHj3sLFtrSJiN1DzlhdAWe2kcNruOEOdr7KX
Li8rIYWq+3UmYfEjDiM/hN5nY/shgFyfmQETVMU73iXM1i11nHx7ESDfsqXm
VDdOYu5dKnLn4cfEmiTUv+00L9lQfaI0rpkuoZASaTYwazmlTN89bCWFAGwz
lz9jlTBGKkhuJWCo95eqhXhq9tasULGzxqqbI3mi0hta3Ug6yxTtCNAB48Wi
6sb559PH5LK+0oWi/cxhwf7tM4xU+kseG4kVW4vjnTuITHRfNfjk/6028wiB
gFspcZqdL2QvwoEtm1GflHZrLBzFSjcHSTPwx7XEvTRk/dHJt/Nqq+8+IrB0
qPfwxCbF/GpKwj11NhFuNhPFwybVJUuOs6Bko1yIdco+V8T+3A0gd2xpudqe
Sc/d3wK4eCHhWdpQsw4euaDZMuRwPKPvJnqQKuPcO6NChDJkweBSv6Virk/I
ksqafg9NGpFF7pfBvbIgDJaOfoqvwxUdzANE6LeCGwfO6LMJBd3wTGmPqA39
rX/envetJdWhPnYLPKitmeiMlAPjQZ5CNixGO3DGnaa2rgL54q5Eag22Nc0d
XuNrIcNKZaX1g1fnxjl8scQcTH3A22IkWdMaatQscKtnnndCl1a77CCHig0z
+Rol1vX0PtDf0mL5uIJNKeK0ZjgN+X4SSLwJqpkOVDE7hjC+KjgTztR6HAfU
JJFch24WjbY97yCnTnnZWxPIRIUWtwfkeKOTx95MYCmFmze/jm2p9kS0MHiI
lfV7JOy3Nzlfh6gUEdS2eOI4bgenfTeIhIJooHpPwwMChlXbPOTkTiTrmESY
PdKzQlIxWkTi8Bm2LrlzJy8i5SPLxQz7DYEliT1NfFqTiFE0uwEFxJ/IaRwu
o9vEjIXTaQSgkApWDWsTkgPxXopYZ9YJYGapse5Fa0XtqppBofKKwi9IAcK1
6wJS0xkZS5N816ubkdWsZbv6Hk1STWvM2ZWv6L0kaoIrIof3ket112jiTFBa
J4GhWpU/n853AJBvGWpRLIXVXZBUvCvldkyAHmBdL3yBIRr61fmidlVbxiFc
74lVR8Nrx/HoAEBq9yklOGfrGSv41kKKo9mVkank4ygMJkagJVCrzFX9k6wE
7k6h+c7xvaDYA2FgIWW0TNAsTzaWfqQLNQKax9ReuzB/h8sIpev/IK7JJCED
M42hGC5ueUN2HnQVy2pHLiNtL/j9WK4pHWgxaKHZN4bABk8qYJknivbcvh94
gM3l7UPuXf8uwYlRpXGeVDv8/QwamjZRNer8JfP30QjI32hq8fV3YeIGCU12
r2leejEkCx3TQSNaw9MJBSbxeZFmX4GkQjGQaXIZWhXcrCW3hZWv5PKKWWkd
2t+6tlAzURW7WY7XhxSvX4Fm/B5pM5/C9ywd3h6tRt73Mt3F+vwevTquNY6+
cgFhoSeJEH2cPc9+8taEMLh7S8Ug2767mShRg84ZYGWOJtI0iH0NvhcCZQDO
8d1XhZfU+JCyQnHlb5WiVPLrdtlpw+R9SgdCuEVMqIDBQ7gc81BzNsrfZiW6
qx9agRxafQMwq/VGV6PPQX+FRVpjl8SlP9PZ6uTfz4VQJDMNXW6JKZHx+hUH
zCcV1IoS+0fOQPiRBHvAh+gupFyD0JJ1jiBvY2PqAuJsc8OrjKtgbEnOmLkx
mKqXZj0tGlSQ51PIVZ7kqrcBz3CqkGlvSYrbNHviXLVfNV2VzP/HbqomcScL
QnhnPQBuCZQjOcAb7eEflDpYrePIOOweMsTyhDmj+jQO9ODW/mw7oM+k0UmP
jJkEf6AaZsd2t0Q7uyur3fM4iggYCox9ydq0GrtvYBSMM6xSmvsoPZjXM4cW
/tt8fIhyqJ7sHHFD6qm6NstS/iBxTTipVQSe6DfK8t/BUpy4dkphW6hQDYnt
ARwzj/aa1pb6t3SXMJMLwYseyHwGwEfydC3Ltw2vi7WzwIkmG7/2uiU4ARka
ukoiZnSqKN9nch5ZZx5W1S9ZxlH2lx8nManglzKjcSdoICHFVXGKcqmiC/cF
u1UZIl7NkiMPvefwuVS/s+rrgHlY+T8D///fOmTkwl5ZeBsqtHMymTgg9SC+
tmmu7ODIA83gpOXHcbj2c1HL8uLNtYMA3kxeSNhP5iTBXfKsYInN1O2wsaEy
L2sOj0o4KdKZambSAokU1aQCT05zwLwRPk5Rn60xBDwZKMikCKH7/e85Tk90
fKW5TBctvKtK1RotHNral8V5kt60z6mdmPucYF+0fViqV7dKMXS2qxoLDfbF
tXAhMt6t3QY6tRlDZx/tyXDm6nLY4+TvHZbpJtfrcmMg9bGGfVP0ixCZ2xeZ
MxWTiMEb3vCbYHNzDku7BFMTooe1AOct6l+h7NPWfHJMRxYrfiZC1TLEokI4
u8rAsSTXBNTAHhZVXj6FKm1Qv8ZwIwWBcHyPexznDJIkf/pBGsJesJbOmi0c
x+kYUfD/avfO+VZqYjwxBsEOHT5uzRp3sq20e1IpoTyQddxSaiurHG2kPJqg
UoC2vxYJFdMC/hvMOzGionnkH5JgWCepK1pmhwt8i2FZBvjNKDWwxLCKmoIJ
lFPkcc2D+F8DpmIx1xHozzVXUArvgV9OWGOsP5y+c1VfM53WeMoMLQVguUq+
qlBoMT+ZS6mIUcwobDm08pyNC+vz8BsfO7aKnk9crx9UYuT29L4ZFr5v7TKr
KADaOJ3YLqxXCK+haRCqtsHrXVK2oCft8guPqgaFLvREkqSc8wpnyDgQTcN8
XeTsHF5K4z13nBbY8z9H5RzNXVBLqOy4AQ9wBehebbe/fxb2o/drxH0xyf0N
zFF7xd35dfN7r0HS7nLURhYhsio44SfoWFx8yREpfjf1S3/A9KPxwiLrfH2k
+wsVoynJjvARBg+/NTmlKPkfQhsDkPV7rQE8s8+ObwAAB2aQx6cer2rHcNDc
hbE3A8EkTaZxzMRIejbAm6h0IzXFWnEqBywqbzpjOuLUsfYNelv+2KvV1USC
HP7UPvhdCKFJfmbOJWUnpP3SZv76VrvZYmRiJdMDjtSq/Zecud1U2BhqMKXY
bAA1Zhjx8Hq9m1w6PJ+GenIxiWQJP1HW3C8BT01DpDdnnsJrEPim7BGSGP+L
ifjeDjFCNjQxGrgymeqgMBcNlRu1sBOJZd5ISDRQxgG7eDaHk9+v0Lncm+lD
oDIGoORP0T+8nKsne8C8RyFamBb8ttBkw8SpMGAY4fDeIRqcAqlx/kJ2okK6
aY2eIX5n7bDQ5lunEtf2HdyUKiVhMQPEnaV01T70dBeeAOY50GS3iH3B9mJ1
hA1P1nWjGH7Gs88R1qkilnERxrAiFR6kD1kLkMa+QTzdzAYm/ByKFj4+INS5
G7C0P7nbqZv8dQARJ9DPNryENQg/02csZhjViIZU0Aj6PYLkszPMkwk3mjJn
FfJbdQjMVrqVzACzMRmssbGf4WWmLDZ4dRWbTKqes6tyyrUCJUW6orssXe6s
KtWLDAFJvXcSHp19aVZtmIWN7gt5OByFeJQqPDHH6faBS3BIkt+0mdb7qQCJ
/aK5Tt9eFEidIIA8T/e1CD3YfHNJkvF/AJPWo5ysrTqJP2jlKilo57jucF3Z
QoBHvcv+r1aDBj8Q3Avlab9eNbifqXRCakOyXF0r7Djmm1tYvz0+dR1ReBPo
sbvMW1sGTqyB1ymlYktajLY49WVAmgZhVSewnoKjZLl70MfE417D9hKku57P
KZB2Eqoh0riKbZpBT80ZQtnXqQiLXho5abxc0RDgivYZiJw1z8S5sHaTp6nM
4/OvRW5V9IYsJrS9prqNPVaUZ0d0ZJ80Z+E//GoqlXhqn77J4/H0fLf9a/Wu
hDHJypWcktrLJcWJFbj0CrUBmvP/3GEYYol39msQ0UiHNF98KYLOD7+QoDHk
SFkncv9pgHrDo89xmN+SCrwxIKCdYnCErjYfRnA17ejVMFqRSwQNy5BIMxqd
5noDyNm4DK1uKF5THXm5d/kpKot2/kyF43P69IuUBmlBgOU1wRsethe5lwUE
eygByRifdOdAwfSTlJhxMruEAktaekngETPBDYVO0ybmBp6I0wg0mrdXym3c
zjO7MoLSHLnhjPZvV+7xemZyQOEl97KlmXcU+o6pxoeb/LeRu9HcuugVxtHI
IWcI3TGPZUd3YHiHy6ZzXLsOq9XbUqf+OZr3/mwpl6KSqkBS8FAFwmUQ6o0c
/9Qwu/QYWgNo+DexUFKYRImhrBuJHc/DpKryfRglCgysDnDr7wPKyHLaf8Lm
CXy7Carj4BvSSM2EK+J7/HJJws1dDc3tnQ9SM5g7OSZsewV66bzGAnWylBEb
YiKYZg2y3TU0h9+G0hj4G2dY/8+DuyX0TFnVxcqCFaSfZDkWWxTOydhythtt
koWjwlDK4k0MYnckPcdDFgEKOHqQxWFeNUdtmNPGGtwmiwB/Rvf5YmIM/lEM
aDbhstw3n0yBxKeLJ2NQOXp8QjIgI4kzqN+IE2+W33b3V20u5bxCC4sqv1JX
T70BzL7CzdkSrnnoR9rRKOYUkf5D3HIc4/Vag6bA1Z2tFCEpiCLt2/SniMVW
vlp/a/vPe5G4wQxwe5JsJgVKDu1nXPvmwli2zZVV0QxMLEhvBf2ocqJGn0Lw
uqu57dP+toX6vkolKjbKVo/ymPq+lkVQ4CmDdlHGs5yhwmpiMvefvTsbZPYK
OE14YiDcYHoqTW82z0jDhe5g0+RECBP3IrYkOw9oCXv4em8nGMw051lwUQTs
Qedd0NwTWHqrKF3mOyZ/K+6VmRtazgcp91Q8KzhaTrwl/5GyVnP0f/exJtuv
7n+UyYJKTG4UG4AW7h8F6IeGVboGEIkQm4P5up10n6Q/c2agrarnYsrmdm3N
vgrt9AtTtn/zHWZlEWS7u5EWVjKBDz9HKRL3dDwNeCx2GeSYLyjaphYSGzJz
8wED84BOti6zhGK5R5oMvVOtKZCd+MzeNEAMNaRO6o3qSJGfjPD7eLT9ZtjZ
LvCahxLWdeZZUV8mw8kKISm6mhYAC61DQ5TVhsYzaERM51VebsLI4C6OGdih
fj5KziHjEJjBMQtOIfRteK6ijWpUyXvUS5o7mRAA0k4NXHRkIPteK5ZDpW3c
G5n3FWp5yEoIFb5vasU71kkdtkpal9lbwjQkjp3wpL5s0xcec/ipFLquL7Mr
CmlUesi5d/PmIO0on84D7GY4gvjzHyRKy0+7RFy2U9CW24ZRR1tnVeuB7SdU
HaINZbsrZYGTihmHfxd/4GLuwKA0RTM2T27rcWe1rgfysgyFwtfYAQk/kvLI
Ad65ykbFZUmdYgx5QbE6CBghsdL2VGckb/QgY+al9ksb9223IIgeOZKwWvqo
a3cBq3EDTfqsARYyeg65Ch0QCaI3W+1UvSPe8eCMipHRAIsJ/7SpCI7RnAKH
/MxcKHOBM4g21ff51hYtKOnA7BzKaKE0382x6FKzI/J9Z8clPrh9lr65q/iy
/9tPjG0c0BCFXgM6wqWACgiAN9AaD+yha7PbK9fdn9beabsfPdjssFb7ME77
S6ihqRZwN+7eKDl6g1UqALLhbyBMeloi6pwOhOy+TKC+IRWWwMKNGHNb9J5G
jsnggtyBz0HL5lXmlYUXCDjZ2nypK+zcTgDqc3vUyKtHYEZL1/bOLoRoettB
KiGnK3m45VYX0uUctcJBATWRmZChXnOuCB3V4Pgv15BLgzy1bYQqUp/EyXeh
FVp6I6DpMdnb6AuYwziIFjcDvijZ5wt4sM6P7EGwH8uJT9OQbGcN4AODORx9
ywfg5WjQhUQDS6M41WEuJVL59DwyB0k3GBWdBoE5ZjoyxrlR6CbHmSiy8tpM
8NNGcSYx5/7NqO7MeZBkT3pwin7dQtkA/3eCe4CMpZZd4kdfF123tKHhqxkc
yM958ojUEwJGQyl5UeVE6acf/Xdj/vYebgZuMujtXEiFo7jug+bWmSC3vTat
818RB6wnqXBaC5NIcALzvSXaqebtkKtm3HnMnocr5WvYzMoFaPSvc1kge1iB
RztfzSkUQe4DtaMAf6CZj6nHUg2QavPi3Sz8Xga9viP5FKnYvjrzz/Gdc4Op
yqSTDI3wbRZYZnAjdDt1ZwUK7mDwwJH0K/NkW25DNGV3zTLc261x8ptwjvWg
/qfDJdq0x73byHhnvpkU8CansippON+5gp9UDfdzW/nZl0tiAAnZy9GSej+b
cZVpyOHXjJfAW81c8XWelb7M5WYbSPeNSPZggN4e1DkpblY22HQt/THCFOQG
CYz9xRnGzH13Kjyi+7ZNpufq68ictAU4P5rKmFsmYA0J/xmPAdTyBHnSDpOm
D1377WOkVqAnKUa6I5NospPmLTg4XA5GwiHsjMc4lyOv5QPoYhkg3vOK2s/I
BYCaAgjqdWN7hAmU2iZ8stJhFmyQONug1oFvFNYshDDY7gJmVNTs5PviC+i7
OJWn+fU5ViQZAGOp+Suy7pLT2gmUyRoHq59uieYznmDPaLsZ5AG8BKVxuwJU
x7F7p1NUDRtUNMqd6yoT4Ga4OLNy1PAvYQRWjF1dvELouSgdqXEXc+cHkMvQ
6OYGfKCbxEhR5h6mMxkYNr1JlReQ1LB8ssc5EagO10Py0/yJTKW420Ia+gVp
j8FNamVp6chjRFQLCaKgnvbGC47yKzvwo4Z60JfFopQwisEISbEbK3aRJfCT
Tm+WEb7cUDJ93L1geCHeVanTzz+ULiwH7Y5zWTapRKtdGRCmjJZUofCFzxPv
nwLQb+zwNnTWhQXaSa/XEu8okZrG+TuBB2J9IlVTWyvvjQOm+x2S4mu5NQ+z
hJaVyPvCYQn2SKsFM2uYbXxvlhNDYPimFkoBnrGM+t6IcdrQgfbzdi2X/I98
hjmSbYlBX7GJHj+ISVPyzx9o2LXYZk4mjbQLx0cMbUcZWMY1/8VIV7T3xXV7
s7AgUo/sPdL0PoggPcVE5cnOE4RiLthnjhN1A03epr4ah5RvBPSG7pxj4bsf
1qoTWG9c3PbRBeHPARLS0kCjwUm7EKSpOc4KizfFGg5T5UPPY9IFhEk9EsBE
DxQ+T6uVUs10Pyqb46TVhezfQQlK8JbllJNWB0F7KAdnXDYxoM2mGdkn0GIr
Q+pVF3Cn5kbSWt0/OZjz5YemU26UHidtFXjfHHc5mUeotQexVGVBiaNBh6Dl
BbnouxqlzvMfumV4ht9+2oLFrPOBRXnQCjC9UQgs2v98fLiEpBI+54/BdgNb
EBlMLpydPhu9uLBO9LYqEb35Gfw7L6z0myv7bMSTpPvQCHqGXW66iZ6kBQb5
UxVuOZdEnIfa3CosyxXTBOcjoc2JzhtXPbd0B7pp9v3DgO97gNCz3fs6ORAp
UFh0kNDDEzj5SUz7cNb5fFp1FN1W454W0IQheX7xKbtlxaKo3vnE2wtkxS8Z
Nb0uj+ypw4eTJ0Okzk9nTvSlRHUMdPvEat794cc073LyDfcd4yKwSdEqtexK
9O8jL+nYqula1gt+xn/sMfp9xsqAz5lrymT5kyez7F5ut82X4YH/vGz5lGf2
lIPhyZDuRN0Djxec2DJOJm82dyLNZzg2LOIqwPehYkPG+r2W9jc6t/f6ygdk
W7GSiRJQNNcXxU8TFbRbkcsYpWRwaLqXtDxIDZc4muAs+Xy5Dfh1hhBpbxMi
AVe3YKzad9o/f2Jn8DK0/F9jflSUn74bVLONFViKWnUjpTkfIqqTNNPt8RZM
sYa7u2Q2AaZPHRb0TB1eQKl1KhRQqokPrwMa5T9Pryyd7IEP95td5ClSysIh
AAiUFVWAr0suR9nj1QH7M1LtHd8j/osEyBJNrMH1htB4w3XpPZ+cb+fsw/Fc
NWp092C32pYnH+tOMgc3i2HY+YZGf1q79ZRVNFNhMQFuwpgWGsuj+tivG2Kq
kRiEe27jIkBz8RUPGGmpBre+R+ypdp3VHfBMiqTDM4LG+fCkIR7tOeGmi8BZ
ZEO5BiMTiiIE1t1TTj4Vw/SCLvuhEwyElOyqzR0EmvVyauhgyisgW3ubtb1g
LXcLTmUhDP036dZGgBAwEYcL865TXLMV5qhuFIhYo+wAFjekBEIt9lXrNbkQ
qYQgQiyVIRbLV7v5Cn/cpfoyiVJoRd+U2C0GeJaOGmZgkMKFxqoABm03m5Fv
vAjQmX/XqrrI4khA5iQM9OXbTI6zEFQ67bu/9R8dYRLYYab5WnS9hkfryqEe
fV/QLcQYZ4GqMInbixfDI6fedzIWCYdwtDu+c95ztv2E3ctUshFaWRuFWhoU
199fUWa6gbAIxEVSb6zTh1SBD7vGo2PeJlMyg+NTiCnwfToYczHby2+UsAKG
Jtb6jdXuJFfvnUKZsZ+qMCYSkZY/0SnjrVybe3rYzqk/R1crp50qe3fUKqAw
CRhhdOJK0WcLFAUCPtvXmXM2j0Jne+69d7lLpKLtXgIYgyPv1zB2uWkomphY
WkGeVJ3Os6OnwZliXRdD2U5kwA7bfIzyuPUH9hykgHGkuyruAtvnXPnLDM4B
ZBrz+hYTamyRRk+ZgXKw9UnNqT4tdfHZGvxfthJ3OF72AqUo8St/x52/hY4u
Cl5uIa0tvdlVmnzT2G5Q0RnDeAKmTo+RQFAPGL4ARkvpf6Uw4ENs2urXimGi
ZEuc4ZmNZFEa8wBynWsEWYTh6p2QBlLdOU9nSJPwBLoFYlpFD8w2M7UpToeR
qOrXkzeaBqygYXMpImT2tiFim3cBaM3GPT7qVF82KclLVkucj1W1E5jw4ZcS
A+dHUqqIpuNxhfWhWvKaQYpPkoWvF9plD7FSPXreRDE4OgE09nNNBBuRAvU1
0fUDj93ps8DkPaS9qq8/bRtZdMDpchtfzSfm4Oo0PD6eXtWUuB3wnN/xyZ4V
ibhgZw+4RKATCHgQak31egt2QvQT/NsFf9UE+UW0choU+U2TFK91rh/E2J6M
74m+0CFmRNZz4pCs5J/g3AwdnXxPUAtwnek68XU1UMUvVV7JN7N1U7Pt68GQ
ZhITfR6l/vKGI3oFzGsOF2z/HXM40nReZB06JOkKquKO1f1FYTAM5tk2jhiG
sva57ILFXYxMLyum7v5ERCoB/VrhFWtqt6z8wHRGBKorPoO79cxPGdPQrDe0
o98BmEjjCK1ZzblUIW48L9AeF9pKgdKZ5WxvwgIkiUTj4lFW+Mi7afEjUW3X
aZ6hxwB0jPQWha9S+YFiVouJu4uXtSQb9ryRovOzEuhPl+7S55y97QkQRVPf
Wvg5Ks03vPNVt/e1hG2zYiOpVB/EqbcubqdejCCYNK8OEym7YwCaGLim9UHD
EfF5gF0flNYUQ/IxVBNO/TS9NcDoIvrQ+PCJMGR1WlHvCBs8P8JSmO95Pu+l
JOOFFD9xmtl+qheeU+JyROD8pdeJhG4H3zwBDlSDW9T0fNpFrKAVFw80VG6P
7c+oqGvOhAGcngH3r8iJyYfW/WgFsD+7zYsVwNEVQiLBFZHRns6njUaO2rKj
a+lp/Bd2fom7SibkHAfBGSfIxNwX4ehUi7D4RrNXqXKQp8RA1HFJjAYF9aGz
QnhP2PWkTRW2abo3UJrf3X2jBG7vjgGcmZx+HG+oubZDavLEW3VkqaG/EGTN
GWA9iUPr4ViivdAjbzKVwuAxqf0Zw/bocUxK4WfxtjfMnQqzNXQCMF6wuH+a
aGwwCRyL0CoUO3GLfCuwpq3cWhftb+Cl56ew99EXSyQBKal9/edHAOgixUvK
35qMvGtPjTyXcnw2fHfGtH0lQXCEF37xrgHyEddpWxpRejhD+EZu8SJJxIAO
PV3RcNORsWIWt+uI7xlW0g7oulM81/UGN9qL0X+/9aymq3Tm90ZypzEKCbQ7
jVXTN0IYUUX3qd08u6LzFYLDJ6edXzBAangcGooTxNFREyMoNWiY8wpOQZLI
BdPuqdZ/7tA8PVSjua5opO5vaJbwDcNEnVU5cQSmBPYd4UVKtJzoN7/397vk
mYTnoGPb/3KRlq4FDhbCwkJJy/Q9YbEacaL78vVaABrY/p0bywJzFln7JkG7
pTWv9s21OkL8Lbfat7ShckO1RjI/K2RutjutV5nO7LTPqS35qHSkVouuMxRB
3pJTAuG1F1sQ2s06TvLCGQMnLxQJf9he/QhwVcnv5ANRNX8OvwrDLggSlxcW
IEb/y1vnNub2+Pm53zYmKIRfTibsPFYwMoU8xQfYjNEuPWX66ZU8d7vEfyn4
xdQ/Lgf1yQZHuWAXAUGVpUoEpDGC2ti8MoCjsLJITs5Z8QcbJQkX5qjJ+GSJ
fYbTNPXcreRIrEFDxSknAoaERNjt2GueVggBw7ar9RNpfnhgxIum+VGDADny
cfStapToOVJXN0PzELlsRX6hBwAvvqClJmsbokZQM3pLeOK7cLebXK4WN3Yd
DCX08mNcRFjomiveNXUEB4DBDzbd0Yh9RS2yGpXQ6Ok/5ud8hMdjDTPNW2x4
77rWiGESEzfkehjkEtyPJGDsVimiEEH0UMrR51hV6cjcsLsnqp0lcC69nE/1
3HSAxOo04VfHUZN1umgXL3bkTNSyxlwKl/CMWvUoQjFGIZUcVaq8j4E05Nkp
jSNPa28NmDmR7pJZAkLAtnpAwwbq7x3C74mwzQskr7P5cmSoINdufjXpARqH
KD3HafqiXpM6NnK9dj0qIizvYaOyrVq8r17P6dgP15TC+AvhwZFJQX+ENMXJ
jW3b5wOhr+9sn2fLttjy1MinSNbk1UMyDHABrof7yZ4OHe8ZDSqM0oub87m0
ogMX6Rgyj3cK64OUGJ8bsDZEY7IHWiABVM7KBXVdLdbE59m/p//obkfLZHqd
+ltdbdeWCFABIsphU+hdrVIgTNTGeIJvAUB65KHwRrnFV/8hvjQWCdRDzt+4
kqhyLOPApeSY7xYSHnIUG64lyEnswCJR3jU3/16uR+0DBnRUj+t2NwtD1PiD
6JaP3kbXqp+q6xCenDTCGttNfH0rq2KieHT0o00GSS3VSCfZoE9YrIgipBeT
P95G8FwDfTviyCCCmvSDS/SijU6HUTAJLK5AAI0Q788KUrOoMJLCqZJoKZ6h
4oHsjVQdenKGRZFqNHBebEcL/2JyhLvmCFNUh+Va7F+Qj4rWcjDDRpRRV/+x
Gdye528d+yn1vypd/Wy041lgWWMZuI3vS7UC24Sn5RpBx4EolPGCkUDBQuQr
ApeDPoa7rcQ4otem7Lc1a6sEsNFsZJRTPY//boUUEDliIdmNgnlCflRZiO9r
V3CTSGPaa0SftYteafjl1OtDvwBcfU+wWclBfI/cgNnYuKdSgPfas27LShcD
Q3Td20hFK8iRCnP/LscfeT+jqz5ckzh920cVHPyVv3QZqqegQZN3y2zJjdJs
uWrEs7uza8Dd34+dIAIgNxWX2KGHcWM+Yh7JQ8yA3n9tOFp/HwKukQStkPef
afgETCwSt8WcX6InSRxqVpMssJsRsCcOiZVYmSux5mY9RHkgKDHxmm2yVKUn
4tmSQr+Dj/apy143fetHI8v+2WqV5e3GR8ZasBqEdrfdsLt4CYWPc+lZa6uD
8yXw1kxpoFXBjG3RmZ26T2oBfg/Kj6iBiAEhQg7llg5M54MvQdoS+r2J8+e7
0a8+zm8W+/5By5BoXTSy3Imiw4gszuIB89YX+2FplH1x17zB3ExnYve2lZ0T
TXZUsprUa8K/zYoTuWCyxtSNsuusWS2LK1CDW+pEseR7qKueBTMb0tMXejpe
bCN0Gf4GXZOyDMLOgS0qgdCS/2lP9rIa2lvLD+dtwEB83XbVB5L+zdyyxJBr
iGCbr2jv+Y27lTTiTLxCYm387Yrq2M6chwvSlkqwyqA0lKiWNoVfNfvSzD91
9ZivBMKGtHAFV3jDdh3UHOpvXXVFQjq9bViX3hcbvRizc4KHpHldCafVAwkL
W4HZJKfEF6Ey3nh7Pr99Ulmk3cKJ6K1hj1OxlrHybG82A6xq+dxBC1nzuzDo
WyxYjUOqEijK5BcHMsI4fnjqUEbsDnB/EICX+a09F8GwhMphGSEfDBirmAxi
A7v4ayOjUoGz7vR3wSgWreDvsEZs2ZyNoXk9PFpQmbDhL9sb1UkPfgfGIK/7
ZCut26+kEEnOf0IGgob9UbxiW/4YLg6M4sg11Q76hhxbH9zZSKKoB7KVRaSO
3rcSs6dCRJatzB6prawyOZ/Wh0R94WHyXlU6vWlMlfmAsFnfTS7y2jvePQzs
vH/I8ec+dwNK0usf6uZTQppNpt0mfQSX4j+lPEaJwv4GPfOT2nSm+dBHlfiB
LURvck5Eewot6U/ZYnhGAxV0dUcJPacr8qspSEhXMOStL/kD8CAoBRTlVleL
E7Z5tN2GRqdyD+zMiVLpWKhUivQfCr+wgGklRR8pNqJI7NPbCSFyc9xCbfkY
V723GVuWgZ6Oyeja9jWp9kD6wAEaD1lxJDQj2b83/b1TCN/SBpHdssFN8Y1f
EsrbT5qmpwGR0oKhe2r5GWMyA0RtzAC+1dVuYgmFq3hvQrAf/VOtp9P+mbgf
N3gL7u/fsS58ty7HiVOm5EwT0UEHNNVszguU90exHkIkk/ufEHKdIwPOzlex
N6OhV4iA80YJNeBLl6k+XmVDzl6KazFT1vqNoY0AWGP0mo756xNiyn51ZisL
rjXOV8Z0iveiFE+KI/v4J3Lj2IHp9tgfvSofFzuAWDdWE79fX3IrXen8a6hB
EB2DxIgV21RdmqDATqDp6LB8QLA+E97q/lqSo+BITuYeaIXtaiQSwtJI1buH
ozf03sL2vPtlFYhppMN5dTjH2O3JZgngveDV30uF2DpC9aN1UcKLpEL7X8T0
SL0uAVRELCHbE8l5dVMpLK/hngh3XpUI7KmDeZfsjYJVItPtQeeGdMfq45kU
sq9afDgj0dJYLPsFBw1NdELiWicKNNFx5aSjFWlz8umN5Iue153mPOfp/D5j
eevTvBY6Gugw0F9XL+hO9qk7mE7r6OLFtqw+n9jcUwF/NOAEUD0gfaK5iSie
2hq3UD9l8KEpG/5Vd0ZnJ886oz1N6zWm2kI4ijMQXFi7DLJ2JwZIMHJI0h3N
wli+BAulw4x0HEF4KgE8V7at4+UMc/rILQiGAU2q1jbh1nbwO7Rkuue+XGXP
pq/nkSXjBk3mn0+e/1V1WJETLqJCXeEdE9uYSBLZoHB+y57r0tbaF3XaJAjr
tKsdo7NHRDYuY3ar0XwmgtGDCCoV42n4W9GPkf3XEgl5dIHq5F95I3ctAAxd
Azy44gxPhvNhcCzLRbnW1BqCqo2XOZSCJojcrt7FYZsgu6WyiW1V6Km3Q0ye
7eI3E9+F48hsEv9EtC+X7mxQ9Voi7wdRiTHHNjb1BCnpzA8RMf3PZ6BL7Ygn
WZYvDNSpxvbmSsaBtt/WdNwNF9u3S+5YCphR50s+kQbDubkgMghMzeoVbtpi
Z2mKjKsvbOWyZf6V1r4dQZuU22Nk4ZXA1GF6ubzbdfWVRVeU+P8UpUBZYSTJ
7G8MRCnXwHzfi5WO4MbpSqvCjrox8oHkbanpBZRkKNnuu7lDmKuavwN4H5OA
8C8dHDZYUmXlXMVGXE06tPpMFirRr95tuXX/tnImaN7Z2dCTZ3m09OwcY4zK
JPJo3qZjBELvd9XjAtrxy/F8eBp7xrekVu6UV8gPgr5sQmE7tx1qzZXX1qpm
tEwSzS4qynKzp6r3dD8mmzX2PUv25YNAcUA5RHxOlVWOAwM5lnsgPNKRtnYa
zXMURsJbGP4cMrknErxBeL2/fikgYFAl7UVqv/m6oGF92SepFC+oosIIZKUr
fYfUB+RZJ17PWRxdUPDyAnQaH+2EmuvzkfITQkBHr379jNEZoYTaGaSedjAx
OZ5kkIpKCbGM0Be2W5nTqXhgH/N89ofT41SBsMK9LFQOBEdLc+yUaIvCP1/t
fzeoNxw4nPjegLYdYVQupjC0BYsUus06TB8TRyrk+wyVySgy9ruPnEkQmlBk
IsPJwfy6QizubVA5WuXDS4dhEEJDR6AT5vXgtc4Ji+ZHfYcgGwYpmoIXs7dX
w53TYp+bvwEM2bs6n7PoWs4QG0CuBp+sN2ga9dR2xJleyrExO8JOyN6Y5c7u
uvkBF0Whon4YFrgYv+EnVFTifxCtTo8/KB8a0q4zGwDhM+J+xmMeCkKYRq7Z
OiOd1Sr/wQ87JkV2e5D9iS4zb7w73ULmeFYd8VLJUr0aYcBeXmGNUgy4a+b6
gCCUC/xe2jgAMISdfYsa0L+DEAtynIeG56rN+1zTtOZTbxE2AalgDp+x/aDb
agvv0dbLIX531leZP7xCcXa1nCNC+IOxg+XofCq4denfawlPMln3L70hNqSA
l67UIBXqTAizNljH6ff+3XwFjrU0LDQ2X0wQ1KrnwOYEBuyK2ngFgn50Qkh4
C+CsLedVwCSdDACrUqbEptFOx1z54qWDZRX16wLjstLItMvot8NAYJuDR7Gu
IAZxblDqc828EDFah/RTevLLoMdFxTpPO/EI0N8OTwsA/i7qcTspxDWAQJvz
/AXGfxEB+ZTK/RPmZRWgJaqEQOAFs/1hhPlMVehkhOzvm7EaOTfiRoSwAGjp
2pb7+oeO9DvjGjxQP8g7oEwWZGyQYYXgK5wfk5AVTvVMX/p+0dqy9bMAb0xL
vhiEHNlKVrGyjfnKdkO5/ES5b4RBeo6plLsRidy+fX5Sw8mE3ECmqhdcGW4+
q3Fw/ZMuvrMqRNMAYtMacVIDTAnAzbu87Ak+DHF0YodUHN52J38HYNFcK367
11BpbUJBmJqsnVA6ncFvBs5kjduF8agvpZCRABT/MLXq1Xs716srMHpuyBtk
MrjGxHQX/qetysZxgTxwkZxuoAO0dtDKtbFld8fpERMTBfPwnrdDglZ7M6ws
r/D5fpFJvnhVHJ2UwtOFxvON6rHKOmPZFqqrmIlKwSeZMTo4eRvXPiWJmAA9
GxZiuqro1zC4zI5DUdALbNmkaUBMqbt8gRfhFt8GJy9V/T2Q/R7/A+Gk9adT
HnptwoyKtxPJZqitSub0ei2UBKZUOVtoWKRYiQ2N1ahQCf7OOiL89jacGjwh
WQuiWRdvS1AyY3BLLuupwShXziSoToR8nwdXFTPvmzrpI7HfEYZPSeCB6FPY
spZ2zOIEI3gANasZhKjqch6kanrDSmB2WbtkSyEu/9siTRCAqJ9aoe445Mx6
PKRa3OVwK3viIwIxRHgPLKc8tHAOexsB2Zap+BWzRfSYf1WxKyZkasQukYVm
iY0RVYqseHDvbHs/LmAZ7NdhmBtW3qWej7KPSYh5ns8TLdTYXK/P8629LWjD
G84mb0XIuVSSkBQ1o3RMAu2rKPoSZM5DA2w9ASvrT8qFk0icsAqIRYL84kVM
M6s1ld4pI2b58CFh1KC6js3159wED19bjjhfHzv7aGz/oi9jpegNfl8G4dIi
QOGlOCHL2wnTi7X0Kx5poCHnysnmVSYM1OpX+i/x7ZLzgJO0q1ltyhee/5XK
o3ao1skiz4r7MsqkKRZMyvtMqv/gzpodp4VaLmnb3Sb71kUyijgwWfAQZiAy
pKr6DngN5YvbBDgmAV2Bz1lH5pqv2H2OzJOc3lpE8uuCiicm8nW1/c0pNzvz
DhPUesAxe5nhejqzZlMibjIMN+GmtA/ovyL2Y1xUPBi+LllMdY7t0QrPTqt+
tgObbv3TVSRCEN1G0NTUOOVyx1auHzjDfV0ywvOehYrBflQxjM4XEhMfKP0i
klbZcL1AoxCNelGO1miWCnHPWI6Th1tfedpg5hRCulIDcjsDkJjmt313pEJM
IbXwGtKceKK4NI68FBe375kXMH0aB/EWrL7YXoI1eFFHtjuVxXOJsUQX35LT
42QauAHShxgnLiywmmQ02/GnGqgWqzGD9J5NZNpsrLzqvlD0YAPkVbnVkjXi
6VbHmB0YlBAeElogSg4dNupo7L81wJEoH9ClFVtrtGXmCwFRBL7eNIgHp09G
ubq0eiT9JF7FSPe5XToOaOrqRJPWYq5qYhsaOZA8g3l/8ojOyel4jzfowKBi
Fb9Tb1foNyYzIghAVXTNi1MtAHsDEpNcubrH6+vHkFd6DmKF0Oo58FNVs2Vx
vk/Z+AuzF/g7eTMW5dRm03Y59tkNe4D4U+T1CXzJcqPJ1LWlhIof17UW2QCs
EE/1qs9qCks7mM0G0hW3VM+EWUotUnAzRKheDKtoUX0yUWQvPuaSOUOvLYJW
HtsHH9VRmzhQ45WWNi3NKtXI07pfCVPapMh9DjJgZOPTaQV0lgATe+uYA2EV
zfaouf5uaKggli3/7/NdypmMwXNE3aztnFvyKJOlexih5+UzYLrTWlC5Fa3/
rcuuWrEB+94ta/izGSEGA5oH26o32bAqYl4xCOySN4UuJ1CxqIl7Anc9jfVa
v9pgEpxFOvfgcaQ/jboofohNM9m7jzH0lyTT4QThAlm6v2BZzOeSLFVz2FWD
06uJdA/QlvdKNEQo8PMy3d0BJrOuHPj4ANDsf5G6Xqeyu18TUokIOKyhzCDM
8GvMrWvdLloeoJbLDwNnAArn0YisPvd0cCfzw0nY+NdFg9KJRx7p1oPpPzt6
G3BMlZZhgfY0puEFz8ZjlhILJztg5kJU5n0NG2DgZ+Y24iAD+M/O00viFiEx
o3KTghloNdF2C89NLRIA66BBZpMhH+KdycJqB8EAPqBWhxDwzgBl/TXd78iD
dyWaBBSNpyx3rKkpaPGuyQ0lLKtjM0igK2IUcP56KerI9zie8q3iUqBLm0TK
Em9JCYOoJbzKNcHDxRQDsqxYoI58yW5mgknwMkJJW+H/nKl75MlBTJLLcHgK
8C1ApHapzPJV5+g4nLuR1UvE+KS3zDfUIaU7nYvYaRL4k0TInE0NAItiG+yW
QfGbh7naPM2CvbPznnIVNGxeOS1V9Bxi7JcPfgADhZkUKVR/TAW5HwwFGIYb
Et4JbkwHdCKNI9oSeeGCxE9qKIBL+fdYhxJmA9isdt106a4HywIVaTs/WcdL
WdYWkUvtOYbI7LfkcMq0oAO3jjmFNgqnrAMEdMq39QwY+H9jJeoX0Ycr+oxX
W7fxgVkFusjTLueUZTNS8ZvCpLpzOLAXFabZdNfEXWZyAqPu4BYuPeleKTpi
QYEoR0HExlgwtHcwOFlV+SR0EgGq0vwPiqp1WSHnp0pbr2IoGmP4yIIgPMJm
2Usm/0rAN1JjxR1LC5FPrKNW3V4yte2hvGqD2rECK0FJxC/anFhyb7HG/yea
+PoC9eq/63Q8xIpqv/ggUKll3/OoSGcK5wx2N5nHeNolZ6vBn7cff1m3Xk11
exS+AEnTYR6UixByza+Qkko3r+DnaRIaL2SJdWtwQuVX5maYoeMdQgTt7CZd
7l7k4eExs4PNvqd8SDxcst1U7yQGhoaBxtx3Wl7W9C37TqODLTXrwqiJys6i
OKA5J/S/sWiCDDoiprC1f37kSO7he6+RlCvReZDr55AnUDWFgqfv7KU0AqV6
jJFUosK3J5u15QipWe60RzpPwqgVm8WGeQ/3NFrypASiFdTKVvFe2XOGKlBe
Md9llc7Q4dvlD7YxYVP69HQQt1EvcIuJuZ9VG+Db73C5wt1aG1g3V4fB6GG4
Cg7LYv066yW+7mbKjE79Pdas6on5E9eq/B0TwfAx2dvQ88WnuEqIdAoMRn9I
i377SfGpKJf8fgzFqJbdeFmIWGn/pGb9wYAzCEdqWrxWcHt+QY0ZSUJAA1cu
cd+zZKJDdpCCyRERezIAGYplzfAbDXuXPbvuyH3c8qhjErv8sEYQ/YN+DfT8
3li8GNV4eTqCNVxeZ8xRuMTC+MeCEvj0tFUe3meToRgAA3YFxobu+Tfe2UxF
W+DdiK8XHmEu5yCOqizB9GdKVHQ/4JQOH0b3IhKYv/lJVxDDMhvYe0YvkCum
1XEZ39H/WNkAOGaJci0DrRDcj4Ro0JZERjaqsF8Vc2w0IDmLGWNs69qOjjQP
n+84/VqlYloqvjbTEbJP14zJ+JZrkFR3pbNFttFNXJiDenNKht3ampkVYbLs
PwIUshl3ws819EnEsm9390FXxpg6HjLG0BVHOX2W4w5DZZDBI2Szzz7bYY7W
Fghy0TSs0E2ZSzRAIg0+MJ0Gaxhrx9bkxSjKkp9ZPq4eoHKrIT45pH0YnGnK
HkbwnaTngLmKFH0Qyakx0sZ86fTbpNAnYFn5lOy7hidmDnB/5fcxMAqwXGUZ
Qhs2NZ0z+JSIyPb4/N9BN9MdBOD310OMLvTwaycAtxUhltxfJbSAHrdbG5hO
J0IOOxbghJ4TFUsFR3UKj/DfHKMxiLxSjbLIpHltX3FBwprJvddbtKyFakfJ
SBnH71MF+XQOuHaHXOGgBlo6tsDbCvk1FlMUADhpUIKZmNA7kHXxNPgVkRGP
5onWFpjPe6CFgI1pnZjjyEYBgoczlXExwEzFUhSd+bl3lmgYGk3SQ/M9Bpth
Q5tnLtDJoF4nCHC/MurGTfCnmeE2XrGiIdEaDEzba9hO9QZuFpNZdUmGJREt
wm8OBgRectcC4G1iKwxNcyIsmM3AlVTc7+ST75iqzpc4KA/zSGl3Q5CRypNm
W0IDgX/oXL233kdCWZRQrY6RxK/UVAkNmoTWp7ALpGi+lvl662/0+UllyQLQ
sGvBpyXXK+zZPC7IBL9HFC3D79WZCTHFBbjz/X2B/JiElrw2EKoipdW62tMf
AG+5617bRMXXrtNHChsCEu6m7Nhv54VSgZ6HAH05/maAmov+mgYzVuxjO/lq
Blc118abCWfOS7UUcn3HOworIMGM99FvrO72n+EsSopFF1Mb0fiQc7qyHVmn
xmo9jcK6ZN6AlOuTLKPnB8SWhsBdGrsJ9s3y13ZCLs5/8+RaV5Um52bklYx9
L0hCBb6cVprUD6lkq/76baBIxwG35NButdTY2w6JZb32H30ZONeunB13iBZn
1wj8xjmGVJceMSFFK0G7UZBRQy0JY8SCGs22gY7Gm7M2a+gnd3zihD8ILgKO
x06B3rcBKSpe0O7f3g5LdDJw8ZnsyyJJ+xqhzleL7I0y0KSshx3x952r/6uP
gyRbAHHTA/JY+zXXnh5IsxWOqO9QOawnr06CriC+M725YdVa6TLYUzyhZFgC
HixlSaiZdQzeJ1oy3SkID50uvcNSQRlIbRp7+1lJ93wphux4jvRAbd9nWTH7
yQ/h92pcKT4jUXSD2Z33tLU0zMy2BkJ9IZsHKXjhxpdDs4cDmRHxtnvavkRF
qKOqzghMTIWDQi/3+tXsaIWdZpou7JhdW/D2Z/faPS896zQxdwxFeAfga3fs
wFyJ7xsgSpP6Hcnwu4ikS6mC27PBTcznmUSIgJtrRRCZpGdLB8S4SeMfxCl5
5PLk9WqpvuP+UdaXs02JXDry1ZZtYctXlIi4SZbbqi0BWVI/W9dDDprbG/a5
dx/oCJAUBBphmGvgQr6+nuoWRKhH93RWU13RfxQiKnCuT379HYJoa7R3X5bN
5T0QZQtFQPIEfVjWnavW+S4z+atwAsiafbZkc33qtBYXq08O0DE0A73fLdPY
HBM2q4cvnIAaoiQGwk2UcmSzZtxALpNTWMBNowUoIFooKVCqnDyjl/xQu6/z
UinWQEly2P8hnavKjaImlrPdBwTHTwp1oW9PQ7ngXtV06e+1LxRq0o9DHH6a
+F4OXVFP3uEn9rqdvIrwAyPsk0DN2ww5hM1mSugzfk72jJTFfY9ffXNgEUwU
vwA9hqW8bLljjP/bKNuSZ2ZxxvtUp81sRD8T7JFQBks61EhMAFS8wqQ9J0/t
RM3xFsYbXnvZCVwwfVB76SdpbVQ+fdaGSXDt8OLP9+ziAsokJTt4uIT8j/px
DJOohSMCd3t7lwUFki63VqZdNQzTWdL/k/j/CyBUlxclv1ZY1t+6o6TJ6D6R
wBpklfo2vZPobZS9eeSGPDj+e1Y8GW4Hs0XUG+PoKaNgZPq0PYvTSd++q0zh
xvLvFwTLHt+dYEliK/ozy+mgfNwwu/vqIwyjR4M2CyRFhlAKPLGO7Aa8Adqa
86W2LElTD8pCloP9CKwefFvtWgdvaTXIKshCEzkeM+3xKuJvEOxmdI7ZJhqX
O9JMXLASBwXFa8ws+pIg9/d+fAQ9Pu6sG21+3EShxzFQPzmZsPVi7oO7ig4L
JGFE3KfX0dXmcNjloax9wcw2cfZ7YhypYO0BAOy34/PaS1XwIP3EztoCoeRv
d6j7bC6jWuFg9zfrngyYPzDMHTE5lL85OdNMnuW868MaJxhOTjXCd97ZUmZI
jc8uFybHKebP07ysZaFKc3QyFlC1reNUW0IKDrmZGsq2PdJ7Ri8l9Ti+thr3
gn8LF12X8V1I25kckpT+jjWSqc26s3Ir6cP8Y2Cb5po3Rgwp/sXN5Xx8Q1HJ
AfWm1z1ie8YCxSZjsl24ttoXrFi8CRtezXAxRfFe4bx52fLLarlwJd9/PDgL
NDEgcXnpV6Y15TOFNUNC6HdpSm+Ur8d3OhHbp5qwGkYY4qIlL6S7NHg2i59n
fJKnu/3gAf3jnd1lKLNlY32oGdoRxdU+lH5d8M5fqd4aM+Kk2J8/PRidHV1N
KOk1qhIgDtjWl6DhiwoicMmQ/zd1LfgXV+Iq6HEKrKHJ9ae7YLj8VfJrySvw
Qv6aosYuHSoGN8NlUU3vAt5/nrrf7r8qpMGG9hIpMW1zNMf25oKYLQ4aL5aN
9Y1E95i7hcMt9xcNFasuvxHfLI7NNY0lFtZCfq+UwmtMaJibFrjYaLcOQRyM
+WuZHWZh1M9pfHpMeVt3mhdH+wHVOtC2k28ty8JUIIsMWAtKVkfzcYMHW9lo
rC0gHdeiFmdENPrZvgQnvp5bXXkr0PN0ZidCMlYZt6HE6iNKKJwVn8KJbyMH
rQL48jvNf8/OOxtxGKlcW6C/Qchr7xI/+mC3Ain5/UvDMSXnjzA1NZmBzEND
LAkURNWr8UN2tsrTzxNF//Uxu+NDyzFatJdW4M6aouDscKJvg4bvmoABEDQG
/2aGKl58EoPCx13ZVcFOX6LFTasnh0XmMIIgw8RfF2l2ijHC9sSICt9s3cfB
DgkwcjWRnNvUWBoYF8nAf+vku2hW6YO+yER/Jbt7j1hrS5mEHZW+R8ZYqdPp
Ro07XAWg2Z01SO+mRHkh3gPRu/oA6pWQK7Uwmsc+IgXMMHiXazEwIfmEt0Kv
SObIpyJQoJb/01YccSxXr+oSW6PnGptOLxWOBy7rUL4tP/n8XxsL/r6Aqdis
ZA4s/5x0UQafuPVz4z00aHAzaHJA2Z6DqeqC8fIYqwqDbmeZJisxxLMHal52
zXTi2ee4XvPT50/N2LT1n3TvEccqod2gQDPi402UI159PTqS4krt5OcaZtDb
JfL1wDSoaYtST9VWgaldUQYLUABGYVZd6ZyzjYD+hA7GZ/z0i3zJUgPQNnqr
S8Z0fT6lvcvjre4wy+FIlHSNJnGYyn3e0csiQLhqQtH7tqXlI+xQN4WBxY58
zJiKCScZSscCxkWBjsOSGXVkTg/ZNLuS7A+JLzLOlC1/yE6tL+JDCP1d/E0v
IAxbNf3QcWOitSP/eVWxZhTlKve4MJFpE4pElEwqRALW9ausu59Of6LSstWf
XK1PscyY07tn+BYpTEjPEEXTV7izPBXSkkyWHSa1mq96oneVUDkSsZzWNaiH
ytc1CkFn0o2GTohQQg8F9vy3zYl+Wn/rsXGT6H8FxeisR1qLt3dKZNgMTo6l
hUqgXwtbVQ4MtojWK0+VXF3plLh+xkPA6IX2FfGBzkGsR51R+0+N5fZ3BxHC
0ZA1jEoKpMupSECkRLi31QYy0FIPeGvcn2kqDAqyp2K8rgUEMHACS3G7sZFv
HkU6TN5xmL3Eq7itAEFqNR4wvHbistd3tobJj6JFNypIEEkcHY9B9rt2W8g2
9jZxCuN0dHd4Sph7KtRIWDdw8CF87BKCHh9/XipEs8rtcFKFocamQ1pikrUo
qcKxWKMLd9VVXcm95HdFw5+ZA04xFbrgcE1CUMsdllp5yrJv6F01kvmsaUpO
I9Kjt3Bv+oV4KTY7o0nj+5cMgcmpwKW+5dwb03M+N/5Yz1URshOx3MDeWvZU
UZE5Q152VDRDmuUnvFv3GiuqEz8y/Ar4HjmFR7HkkycEcZAzesMhh1DOA7U2
2QsVy/QmzoIQl9B1M9CQ5SV49xv+TCN17aYISK9nhTZsriHLs5SB6fv89RQ0
4X5CyCQm42xZ5UJjl01mPHKzbq8lLV00+MhyLGURGPeusaVESPt5tq+xJA1H
FmwWI0GIpTT0n1RrySLf/JCwuNDJX+xAB6gbjPwENVBm+TPjYsUzUjsuqv6k
WzuSSEauntu1psZc2K8kTe7OzglB3ZZbHeAGjbYCqnWmu7VPRPdHsYyZohBw
3ISpRRMc1DYVenCRNBVsOp4GfmJv3+EDGhqF4qpFq3UuYRhBtQl4V8PiP/jr
mXjuDoq3TosRTid/Dv6IsU37P7RNK56rZA0Hj/mkaq7IFehqfDzcXKAOGr61
Bu1OalCrXdKQ+o99iszgb02CEJ6bu2Vk9hB/Vls/h/VysktgEG+ANR2wxLuD
ul7GHvMPIZzSiE8mx3d3Otd4UV3VbR+3r5y9GHuDdnIFaGZ7f3FfJoVy2x6Y
SK2UmY3zH8yaS6swcMop2LUR9NfKUDzOckvrqh2+/HYohQbFuhxiwBY0EyQ/
+jTlg7scGGR6v/WaeXw1pZmByBDTfnVWBM09jVq7zSVNDdKtprvQR4sxT5M+
pcJ2NFo1zxdrlbPgCzv2lEDxaCsU17iaFJga2+jRvhXY+qQ0W+YEr2klwnuD
09aqTfD1AjKlWwIOSMM1buuJdPK66tQCBv6uHA9mi63W2p9CWZQWPzE0lW7f
ru3w3PJscAfv5EcHRUAKYCNA5q2/4HTRgIrEZfWSQGlfAugSOJo4uRQoOjLd
mPqxFhaWbdV+3JxoEWNrJmS+xhj3qqpQi0apuDekBNUy8i22RTn5GuCxhKz/
QdDmFfzvcbNlrxhZGTlJXeBDMVGA4K+uny/fHaD/iX/0m0MvnDArMffg6iPI
SJ43mXKaaWbDkepy9W+tMOFZzA2TbJO21tCewmWI7RpB780NBfAsRjRxUrPq
QwdHI6/zB2prZ3ETh6DsBkqopC7xHHmr/RGW03MTKBZdS3jWQathcWUA2KlL
mzuJGz48x15BUJfg7FDrk1vfQgf3SmV9ykNX3WeFY8noW+OaWOhtkcyGL74L
A6gqmLT0WJgj0ic7goesRmLukv5kNxwwlbXdj5Dz6WUsWNch3vyC3mkwt3PW
p2ISd8l3Vj8osZvSR9k6GcCEaO4xEJSYuCX1BnYX3s4VsYl7v5j9VJv/zqpQ
iu2L8SwNwphZOSNfknw6R+BZloFH3IEUOaHZlJhPH+u84/MI49JNO2DCHSiq
0PKtEMr3kKM7N+qFOSQ0uLcbdylDXK4UJsRmFEhDyjPhQQ7GfL3emjsR2mmL
WEZpI/iSd9OULCPKX0d0USbL1YRjwqjgXq7+sgpZpcTOFyCRVdXhwwJ0wake
ASbVB0xkOHMs23lZJ35xwS3tP6KPIUeqzZJTzsdF28sNOJsu14Uzpmak8Soi
/YRU5O+TElAcGkDHIHhrR39OCRIax/+/erJko0muSClUzs5Lq/Xpz9AzeYef
ZksvLzjViYB3CWe3FcV1XG39/3GVeihIvt1PUInVrKgUIJs9aCHFnhYNFi5U
CFNK1AxGPfdJBZmsEcPCwPDww4Vse+p+tUNES2gpspcs2wlt27nlcgcfp8jb
2wqHfDLHmqCfBpO85LbN+s8UtNRIfkHWJhUrbkTuIn1I2VMp8/Zo6gW2j8EX
AAltogSyH6cEIXxtrbxLF56NtR/f1r14RFGyeVtO2C9opq770ZeM8oJcz/v1
qUK8AUA7yfna1tGc2C1q9Yems+PTUqTDqhkn+FTnPqg7zR+1kTx0SGoMJurI
Kocd5kmHZ5bC1U6kKUtzIyFfMY2WH3IO0OONpkTn9uXRjZ25LZvN4Scl+agO
16J+NsFAMV3GeqPns4LGEpMkIQpAxwSK34SHXWROMO1JzIKksAK6X4Zbn1EL
OQzXy6lnfUlfE7/XwC/nGWzsoKyq9fNmxwK68mi1Yq+1FgQnTe3YmUvITYnL
s1J7MlcVAF6vvpN8okUjezSDYP12g0F8vwSSuQE28J3pEQsgFatDfs5Tzizk
e/SSWjUTI2vck955cvf2ARrlI5zrfFpk/zOXJnj9l1YxO0R118oWLHxDNhmS
EYYR3NZ0V2lw/Gf8BSFcMZw8DPYLMTVsamsfB4nBPXlNuZ+DlN4B2vI+sHwc
45SsdPEHbFGUe8nh3qB6wXdaau/tfXvgQynqpP3VP9satyE1F6YkS5QjgnkH
IRDpibs8chFe0pYIMHPd9umYlPcE/BH2+9BZoQ7+NDidPUq3lHWFLkZ1JB9r
5QCY5016oX+Qbg7PNa6HCry3epAdDAFQcl1BKiUGYmgvNn1z9nJJzWg5pthZ
sNttVSFul2fm35bNYRderGhV6QTfxr8siH0+QoAjgWW6kL50fgqsG7cxaoX0
Y9l+VRwXdpUl1wz9vvCJ5zKg2xSPOIA7rZv8jJkZD457d0xSdkC0Oq6gUAdM
LipxyK2JK6KYOCU2dJTPH3/HVdpMGRxQgUbcr4aSwd7HDaqm1gu7az5LJ+eI
ibH7gUEcP/sfl5kYQ03Mbl3TlzvQxJL21oOaewEZ6GJSUeoUI6a2uGeqZlWT
VTGTO3tXs7ToPaUIkEoaw1ImFUTWFwCLtVZkteJb3DkgcjMwcw8zL6j5nw4N
XAtGlr2F+MoJ6npz2LrFkTst2jDy8XL9OsmlYHSb4GrbUGAFC8EqHwMknuS8
ntTGNB1B+o9MuNW9wIe8xiWFX68yWWZMRNARPq+tOYao4g+0ISgQ8QqgTXoH
Mwn18QvSYa19QLWHvQduWnB6pX/v/3Af9ojDABFaYXgMxJvqZ9fwC3yqapYm
AbnBo9NcEajRjJmwdx6UsSqX2yfu9hndcqK8O0i+Sba0x1p9Qxeb9BJjbCXB
O/NxppIxS4NsI4YDKo+qm6gToZt0O1K9iV/zJoPtPkRgow0Zb+aSnPaAyylg
iKiYDZUd+RSWdrwrtyrVP1r/g7HYY3NlMKlbdDVN7tpfbTeUcitD+n5ZBjQw
hyhAxI5EJHcYUqa2SQlNawo8PHswlgBkq5K2hDTpu7OWzJSXB+0hWIUlRWnD
gxvjQ45NrIzC65LJ/f3o7Q0drUhi+djKewekX8GAJLrbrJNuKLEF2Y4jky3j
yA0bt8nPaG2aBX/Pb9MBBKvC5JpHc+fcwABwBchZldzIIJBF2Afn2J5JRdF/
Hi/EY6yg/oW0en6ua9mufUz1oCLkQ5s9i36GkzKivyEDQJosQ7ylz18tbkzu
umEple/COkY/cRGHbeeWwpUFfozahZQ+CxcoEdJGnLVU4WH3Yf3PW3ozkGES
Dv1LQQf3Qzn19Ug2m2yvhq8UEgdnBFmUHhj8zeY63FHddyGkHh+Z95+3D318
IKE0XDMr5zCdf7chHEAha31qp/tMpGRjs/pQ6cy+wOkZYJRH7DfkSl4fCL9P
NfoY/zkqKOns19wGLkTeeG9CMjYJCLIcXXNNI3VvflogRknuDm0ZSSjQtAhY
HPt72GJ7rKYY6FXFMZmszuhBGWhRRigCjmy/K3ZWz1hun31tuVsDiFrrBnm4
67DDCICBytjWyaz4v+e9r8NiWIaW7BxQ9BTeUOMDcn1VaJbweqMgtqQxQ9xV
3fDF1N6vh3dsRSPfPv2+SL9wEhANCmh6pOXtKiy1tCQYFubazT7dKeCCV1Yk
iYdKank8BclzP2OQqvv/6/+88y+X95FukprIleJs4LFdH+xdB5LZ/jw5SO2W
IVENawaKyjp+AU6SmFai8AAgsZDgc6z5QLRQYPM9Lf9La7ksfCl52XLsMYGK
GYFU0J3WO5Lk8Zm5BvpXri3nQEzEJg3j5pLhGUQkgPdXUqoKoeBQ02p19MkY
UjpLiiy2OINw6Ti28VGPqOrCTKkb0tUou6/K1vdHmdNLviHdo72TQtfK9yvK
RXUy4uBq2tYozULB92UEpKTrsVnSG6eRZ8BKmsq0SectBsbxUDmVVw7pxmBr
xm1pOySBHFSBKhSFrza+6WOZtSeK9ot0firqi7wmtssFaHiiXgqq7PiorTLm
+kPiEO2OCZRMtE2MK2sCSc1fWPrKzWW2KN7GHAjtGk/YZqvVLPoiLirzfROh
mKG2twGkYuhBELH936P8GxExmrP6M+twhwdi2B3j1mtbGFc53/qGkJwqtgK7
mxcYDlMb01k5uSHwgHiUCpQU085OXDMj+5EpEMvSoR4x7X+GcLXRSlWNoyjX
4vlDzuQcpToKsNmvIzr0tE3FN8C7m3oExiN97VZVb6XXzf+ea07r5cmbyecL
wY2/kJkJzzmJFVf4qGPvgM10U1WAy9SQxM23cXAP/oaIbl0Opre3O2+rneiI
TqqEjzDUsKuUGXy/JKSTACW/OL76I6Y+vkndJlzLwJ6QOyhk0ZVCaiMl2/Uv
u8N9VmW/DMTMrUf5/cjfgtaj1BmM/J/dIzmyWwXTk6KUYJcXkDjftomAye9o
fTp16f1VjXEqSXDy0HtoxMc12gAkqKazcHrCtVTMaeWJhMrZ0DptZn8EZQPJ
y1PyC761qo1a8qxAgRJ1kEoXJOJeARKeQeAX5FYYx85OrSBOrfn3mjfcP2q9
zMQf94vFWpVIIwYpO/JTbQXfskKqU3DaegKAsBvI/ffRZZuomzQVyVgLq6Sj
ckbOlTCLOKr4TOxYrC6FmknErZLXE8V83fwVjK58Lz8LdosLBc80zzA200OG
ZUpbppIceJsd+7unkFG8wluT2EK8RmbjF2sFHjEPB82pW+12ss6mL4TRbU5L
oUvhSVCOahNZ/xsKdI5x8aIvpM//QLSjIHivYgntcUDx9pSXT7NMSLubMvVA
9d26OzoKcKr1H4G1M+WJOxLFuePuIDrMSPXOn/pq2kNQk4/cElOJDaBgH7f5
tGu5QOiQJHSy92j3a2pUt5mcCxJPmFuUYZwbjBKfK3fisNGAaAyehnH/vh5U
vnusPA6gJ5m5Px0gioaUhDhRcH5xJuAKVHb6/lHmd7tdsI5+fiYc4KRSDHZ6
IYIiXz2mjQhTGJ6lo5gKkZDEV2c/hRDpWtyL2xTm13WHYIBebPqzmtcM3xTN
n3k0bIfi6DEu8mQI9vARoQM/HJP92oQatymUZQBVxpMiCqpSSEZtXbdXDzVK
fn6cJ8/4Ni4Ex3mPELntZqzDTq6gSKRI8fOUScbLpvVlhM5Bso37q5jaa4Q0
YUVMgG2PcmivZK79e/KbzYfaW3MUIotnAOKfnaVMHzbszcV5TeQHCxKVxtgq
25Ty+uW2dwNnqek4UewUs6+CR7HKydSVBH2KXZhlmV/HgRltoP+9pxpEZ5vj
y3RrFC4m0Hm2Bk+VFFH8LR0cd0bw5QmecGe04f/JdIzHxnN5Xc9gNsEitfT3
6OMLf3oDuYecJJqNWF+HO5WXygHRyMeu3ug+Gk37OsyO+JOlXzRBdMXYqk8L
CBlhmb0mBQkSIkh5SGItCq/FOszg8/eqsIjzv9K1ZFaBaSIaUC0y/NWO8nxT
Zlf9dESJQ8fa46S2PJu+tFbeEwcMl40CvH1Wg7/nGN11aZ4h/uza/JLO9xlX
t5eo6DLDeJD2T585BvJPWtLQcDI3UlHhkB4JfwDdvvHfDqtN7Qy9yW/Ioeku
TlakkPAWlPftehtwlWVfXfDNWFDpiBhEUgf7LgCKBX0x2uGtsvtfhW1xjFxj
2Z61YpcVe6+PPMp5XJJ5AR9CoOSZd6vNEz9aBF3NBUGQG8MaymmnkiNVFGA1
SxwlrS4X64THCGlflTlpBBX5J2suXoHtFWZM4x2I7fTkRMbi1tJyBuwChHu4
DerhHfOKheTjC554CSim/u63Z7iLy9pK3ObEKWeCZ6QpipzOZ+p26ityRbRY
FGHUS7RTZdIyhQgCAgActBWXWWEj2AEldPg9QeJS65opKmoVmlcWSMROvQmw
f5aYcj7VtGrsrw0HjnFL8LZrbKbW4FasJI2bLMptCw4Ywj5S/uBFXqCL391D
sZmxpoUn9rHIguXkdnkWs4zg7aRnPSF4RQg5jWlkdrffjFgKP3QQhAiBoYzH
QfPBWINAazZqcT6LR5MAtCR7fuyhQPhbYdIiCi1AXaoCFzZuTNvBBX9QX3QK
8gr1lIPg6+AmEZGf58Y6B8vJ//WfJaCVgm4yV7FipprlQfef0i93egnw2s0h
DWG98eX/oPpJzH7ZZOGSOZORs94fEyI5BGRmXScLhXl1CyfckuiePxPk5B2n
QKprRhXAvTn92PrIwlVJtKC74tiuLS0xfxdBtbUWIcSykot/xddQAGlGlGLR
c9a3lbekQgC22WDhtnWoRBCKtsDrIwEDxS5RXWbjudz8UHWPTDBpPZngRFy2
3GALcoAi3T6GNtZ8NqNaz/oUzrA2RCq98rqBs1ZTR7pXRcMbMRmMRN6rd8qc
FutHzFeHtG0irGuza9SwwLuegWCPvqdAG2g5S6ri7PxvoCebzyV0XYnf2NBE
8hhEBmsAKpYnfCTA9U83r9WZuC1CiiSEVHIMPUoo//heQwpCzHbDlKiWimH8
XbdxT0l1UPsRlU2gCk48DDNPOBRTMv1jNL1G+JIj3EeH/sqSG0q7qC19UjaK
UFljoXebIgLU/Nm4/b2eiJ8rq+nWLBBtL4HUywYxdtrI+A5SnZqeoo3sQWa7
bR3L3C5NyTsZFc+PDHsgUuyV4bfXvRe5n0F5KYnD7y8VYmH61EnFOUlk8S7D
Pp2NYDIGZvME3fHUG5G1Kfg2wT/M0geGDKauAAdStHMKAr7wfMMlvm6UOupa
JEKQqTshXOK4Otp+EG+bDQb0GGGQfmQ0qF60+cIeDTza/dSo741sdszMSYki
QMVLTDogk9egsekbjyABoUnevh7sNkzDvwfC7B5tO1l3ZnUoP8KYfmsc48i8
/3RCrh0Z0ltnw2Md7GuXx5LcBfzvTaOVrw+tF+qIwemQgTJDxzHl+Q0Fo6js
IhuREvC4tX2xqcO55IJEr5MuRNLLL17mKLT5iHF2AtbF/YWoSpZb2QrVvbQ2
geLOj+MZhgNAoQ95543yTMfpBMJllWJnNKhwqWNWoKL2Mzz8wj4WQRmjrwo+
Hgvj9Mq+JDV20rUy7puaGPifK8hJNa5ExkOc3oQjwtCAUQBYqJDoDQVh3mKW
YabscOWxp8UawxFaNhFHAt7Z22yXOvKVfsdTG5XQnkAcLXR0HQ+L9/jbkoqe
LeajpjGet5zAK1TqTSVR1xD35NjD2ARF7qYRULY5uUVfO2KviX5paGAx8fMd
ys1nU3Nc6QFBPLgDO3SXVtWnffs5ndEGUmrrJl2xVQ1wdCx9fOx8ku4dDBwC
Lfi+/L1Sx04zPMxBcmLLqmd5Uf9XUpSDgKHI2UnO17D+JbcQaVpRC7fENwTL
siXNYFmZngnqCbsy1k/vDicKPBYtkKNdLwdQTWyHlzLRhvitS/6ipfpZyisI
HTbpTWQcnkU1Ndg0hLzypNxB2sTU2us20WpPOCTxD2kSQI4xS+/MQcn80jIw
fUWwxWSOMrDP7/0Jil5ylbqefnHS+LZhp7sDTE16yAMJaL/JcfhKguNrnVtJ
zFENdTsXcPZMdNZCOxKXOe2eqaWueRx0eaCKPWgrH0yRUSjJMm6ujuRR3fNN
pgDmoWTTDDptqc199KGgmqK47w8QM3lRrAO1rykFQVknhVoDznIx7IIF2QY7
VymysYrlS3iLONVjqw0cZg/qn82i2ZxrvssG95Q7rShhri5CJc10KGgOvNPQ
Npdq3CecRbB3Ysi73JgJ2LYUHNTNNuB3XNh/w2afR0h1O7KuoVegFvEhoR0I
9tRW+jqfITZEKnoeFTrsFbC+X1/28HVZJPYiVhyoWFh5jQSjTk1xjZpUYDPE
A1ZH4xmsdiGF5lHSUrOn9r+sf6FIHlSqERVJDaI5RTzxveN6K8iVtYWsUQce
SaB4Ak/o31umdwkQSzxHnrdGbjOTSIOlgQhA1utqN06OtFBM8JPgBfArKdvM
XQ6elOSZuo4bGoGs9CwjEixnUPllH2EP4dc/iUqOj7TluNZGPvNwtwm6thc1
zKfxV4A6QQ2cyJdhyU6UbfIDrS5ndmj63SkRRYos7OxNVXPHmoQaZ1jZ7AJ7
QMGcODEGkbGq49Giy66LjmJHESSVOQK0GniB1PZFZa9eJVnNcEZ4d1bN4zvj
l2vZ7VBmMu3pNSk5LPQ08YLlaV6GmjqUA0ZfSWfaAulE0gWqqvwELWF+33FB
kUCSKbcIuo92ZH1S+IIrbc51Dh0FokCPlux/8G3LPE2zuH7eH6pt3BVunkXx
JUkQKa2U9xl6bDgU/afdAF+wdHZRTX1ilUCP+KVa6j78q103E65M+2L83WcJ
pQ6q+SM77mLIBDMZf/GPXVeWvbofteJvdKEa2xbP8LpohKXCcV3VoarWOxSp
MPsIno8elEtt9mmXpfxHzVeP/9Rq4oL8ebDYED1l9z4y1YpDcBCp+J9RlRY3
W5fBlRpCtNpsanqafO/gaBb5uwBpGw7dg2yf9qaQczgsKvvwdxdWbM/IxJq6
qMZdTTlJWO1z1fqVoMNaslg8JpocuX4s5JaJShlnSe6lKBuwBIHtLwosXpwz
m12FrAhhSHgR3VFhoSfhnal2VSeZfMH4053vTlLDZ0aUwWpWoFnvFlGAfTyo
czqJV5UjXBdex6pg6tqxc4HmW68mlfD5Rt4XvFBqjwAi3xrdqzf7SSNOYMc2
riJLDoSUgvdFvMn5JSkS6Sq2ITDQKoawMdcc+wUb7K0wWQSVYWMh/haa8v5d
lQWYKlhiUMRLH/RHbvDp6RIBUMMPTY0kA/SqZ3cUHcFB2Nz/iVqpCUJhHTHd
drPZramYD1c4oNSm1xIzoLdNSosqFB+A/6L9gqhPmza0pPOPZkQ/GRB1Yffm
yd0+NYn1XKm6F1l0CdNnSZqhV1jB8VXp//d9t0Jh2LLMv48brGA40yWWPkMQ
etEZwhUxl3iiM3uD/5FL3XPrl54fC+6rJXVYPulXGifZGE0k5epMmaLJs96c
Q4zuI5pcalkOVjbjSWVcVkdzSVTjjSThXGvPofKpvMQa1UdWHaSY1pxsyEfC
xD4zv3toA3Us2k4hBHdoHKW/6eflWN52/Cus0WaSwCtphjqsA8IlpxUt0Z/5
heMEls6jd9NjFNqvmw1u4vMF5slKSEaATi+a5HRc9Kkg32NYx57hx7fk1wcA
9EKR/b6i3CoFaR5DKaepyws95t5514jnRSuQ+GfRQn3fJayhQICDuClb6w6b
eeNet3mLTU0laXIKLvhPPG4krW6QDbvHNQhNlbLyGHkqP6YtTpetvpmMT7FF
wbBy7XM3Phu5KwXGxTvu4zuwEEiP2QEBOFeNWvpRlKFAz0OS1ASK8OcEzbRk
QiN7/9AvpRQqM1wEOJiotZVJC3dM54aao0DdkxoOazQXfMyOG+rOsfnNCUwb
gM1cv7u7qfYO+2g2u3D+FDthoeA4ATMZAOImwRgJ5Hq/ierzDwryDc/egQZL
dFDEQiKX190J4CiadziShpPBdWR9wvG1/Sc7njQauKlbUAAf/ys+ttLIcrv7
kTVPRVDzcZG7k95fki8BJnuTy+1W+tWnRAJ1Rkwpq7yoZabegO7aoiqR4YNo
pV1jdLFpx9kJGnVtrnDD1OVjwALXED0ird/xjRnXE9bG799RRwPuP0+a1BZa
Zp/z7LnC7FAzNJZOrs+hh+Jk839bSWqNYWCQX0qg6WGc2D1ezzJllJkkFVlQ
h/6qdiK+rLhJJlwUIv15Fr+LOXAyj4/klU3X90nfJV+uklg74nXOMyEib/sZ
Q1+0IO48wU65gi6/cqLQxkXHaJHzVVYbuQL6HoU9SNkmC8ADdD+OxgfhP1H6
rlIYJPjGv8i4wX9znPcC8k2uLPaU9Ng+azL3OAQCOZ/mgW7t6u6qINL4KgnZ
fuBMnRjaB/x9YQnDql/q0RYPvm8rXITdbsr4Sqvznjb9CgKSP0SsffdDzZQA
0HT3KW0W+yEPBxs9H6HyIAChXs8oav7MCsYYP76iENzVu+kvUT6eMZqYoyxY
Cm2YkG/HGZKv7e/0GaTBt3tykT4S+T8bL6b6jrZaHh5pfx2GoQjGKTU8dlSC
2jZxJ9F3tKoUjPy2fKxoTA7lkhVtEuBGYKIqzFq7W7zSwhzpc4EORaWx5vta
gQTx2xOLCaf9nj6UGg/aT6IW7RqNQGsQDea7nSpBZVR+AiJ6bT/f7/g9tmAT
xNsW109MWggxTKBJeVn0jqx7PbMGBMW3pbls272pi30nu8YIompKlhE+Wghw
wIFMSK+AwOT2ZuiV8oOWCjHxyOLsFEaHzkq4jUUlu5EATmEqbzdMFcjpvu3v
qEsDF4PfaHfaR7XAhzPj0zE0ZjXMll76u10nwLz6BfiBinJioe4neRJ4xh1V
Zv0/ImEsHZJwwshKq9GnTKTxVu6enK3I3hOLjFFme5BV4TNixxJbW6OeMfV1
QWbKt2hMIGsezIcPAnWUJx1p/6sEHVYLrntPw4Kbmcpn4Csdad/BpWDM91/f
1iRpufuXDXgI1FJ5EANzmjyv5uH5oZCdNgN/sSb9gvjdc3cxv80386iVf3KU
4hRF6Yms/6LhvI93bFtIaVikLUxMu4CiGo37ywYJXSTzf8wScQo84m5D29op
UUrGy10uhN3HqdyxXp2quJMUz/Y1kdfV6O+TL2ld3FnOthJgW5xF9w8snIpo
tJBqWjpEFGKbW9oRyeaoijqD6RZpumAkvku2eO1BU+ztLeOpU3FQ3oHw/bq4
1Jg98b+0TVsxYS4j9lF+pzH2v7rFz5POl8HLwFdmiubVraH2KVlIFzDlYEDV
dFTNirUOj/A2iNlxHV+jo5dtPXd+vmVe6gQLCpho8Xw2d6LsGVklEZrNXa3d
olh+i/u6U6cUuHaUDcR7pKF2Yn1sxakcJzuFxPozyoxBVJZZ4YeyOJUqOGg6
Fx1d41sfD9tL5rrwykGv7nXN/cRz8uTiEz9ZxnF7Kv6qCTD1q6bCNSLDrtOp
KXC5xpz5g/Saky3oE1Q730oQACeSAJ+zRNFVUZELU05auqijjh3TEJUEyMZA
PbZQcTnbeI8JzRVSWnveGsWnaKqr/+cqmceCxoBwa4Y17lq5szbnxqPf2JjV
L4SUjmNJVvpWFKEjknzZ8qmvuc3cEeNq4SvqgWJewnozybr/c3EUsjoTVTIm
+Le9jlMZ82Bhz6S4wrSn5mt4lYFs0nUWjV+1+aMXzv0yam1GmIyIryowSmDf
jEEh8AfDuKENM1uYslh4+hNFr86o9GuE323Vb03OLTXjs8Lc2Z+7PU2kEmW4
E8L2kDhtDvd6ZsaXu7/o6+rsTCtczSu55BAS3AxQD4BZHSakj/Zlfl2ooa2w
r0eiJ2PIyqci9b4Lz1Q8SsXOkIlBaPtQstslZiiYanJGLcy1I75V9OltMTnc
mUPVIrjSEbclKYsVkw3A3YoPTDJFn3CoanYhUnM2g4tsA2GCev/qNX5eESRB
uJ8Opv67AJy5rbVcImEWW4mXVeApyQIAipa2MjU783AEMZdUY0y8C4nXiW2/
hunZ5DoaXfkKxWiiPkKafFhLhThtC3sB4Y1m9Je2fM0igi2tQ8QmNC+VsVka
ZknEs3TY5+vr/EodrN17OT5dpz4GlieVJmi/52JWZIVEQJGXF1OsL2V72d9Y
LfsfmNTVEuk1H97C+V9r0/S/KRFSs3ostLt6eybB5Q5kgilZ5fxYYoLicNmm
Gyh1C6Dq3Y5JXwV6CkhcLBZfMFkgIAG6DsjPg5oVXcSVXMDda9ktPyVDde2Z
fLlkiJrxLm4tgUNcwh0g1SXSoZaRE9AzpshiExp1RqEVDmQFLEvEhIj2Y8Ri
exYbPhqtaz2pS0jR6wG5AO3oJXG4j8ev5jHowXv/Ly916H/damNyY8XYtV0q
/yAkk5JsX4xCyzy5GFC6Mlu3ODbQ4CygItcSJzipAHNYdwKOxnVCKONV8jxx
g2PYY7vXXXmN+eE0loKKs3JYocZod+CMGU++svJ8itKSjg5j3NLbmhvdk9CU
wqX39rN8/k7/+9yikAq7KtOU4T+uF7duFSkTkTJoi5rYoTFi3Q9p4PS/8kC7
T65kJWVKN5OHPZrk2WDrjEAoiggheeTs3qMDVgS8tvnnoBXH5nMicSBxMcpn
/TsMTzhh3ZSCgFAAToxwqWhe2eCvhBhMsVILYb8drDKlI5moOlkNbpV+WMtS
ZM1Z93WO7nj9kVzIIViriYW3JMrBMc9WosvsiP+s1W3yPezkh87HPBque4Nk
2RPrdBJlNh/ndLnw1/vt4xcPyJWU41R524iu+ca32uEmuBOu1yMGjTTTZkTa
nevRuw79WA9zUMjCcCrIrt78G09tvjHe9mo1d1LxmJQ7K4r0CWgU7/KlmF7r
D56caCnrrqMXXbFL/gTNJsQnnz0BaAUNmB6Wjwt1racvaGyhoXZonrKTHmJc
LomUvXA1AP3BCkDmYtTPjS4h0e+REuwhIujcsW7uKkLwwg01HdXyD2tbG8Hr
BuRqtm7kZN/9r+u/dmeNVaRPPYTKR+lLSS/k//m6t8eehIvj4rqAX8pKPTvh
gBJemif9tmOCLRRrRwlHilLyQcfCern5LAYw1c9uPCbkbEGN8miRhWzCKA0I
8kqNkAAQrgFjDLvqbor7Do/mShcyK8tF58UKfahU87QeiHd5IaFN332BGhEY
c2rcehVx1brwz5Os5/PJSCb6CdNJKI7JAvBWVfa8N2o40CwnmOlOxiDjToeu
XFOr+AknrE+1O3UcLHe0Q1JvsHyC85w7ACM+HzGt/xeTj/Huspi7buwBQDKF
5s4fW3G5f+lvu+0GZc+98zERMRNlgXbLkYk0aTvp5gfi/tyfkEKJzI7qdc2m
kkSrrLn1SzSy2vNruDPudcSFwGssmeZEKKYpY1onf7vkz3xvcRRMLXCFXIZq
ON9UJ62NSJjNGo36T4ht1YL0jOmSHbgneTkPSfCUPksXRSeDsXwg/GyLRdo1
GC2cbn1hgXs+zEnRtHKi7pfvrDxDI9eadG6KeKkPD0s1OQOM6qbTGeBfLZKM
BBdvc1vwDJ/39RJkAmoPu90ASJm/7KAhfMnmWvPM5ME6M1xaWyX+uN/WeQmY
k4Y96Dc5pYdvyGQ7oikyagTZcTHb8tahJBRl6U0wX6EzxBm9+c10O4iwctwV
wn1dNamXKI4qfuhSS+BCHZ712tIz6TitiQ0zkQSQbljKK1rhvYt61jF/cYIq
A0QsdYTKbVas5DN3JhajCZNeW7KqyQOYmiuJqrN5VzQxCShol25rbsLiqJ08
9At2op8YsIV2TBGQqWu4x7NH2GteBE6eIkugkVDZ5go1908KYXVZ+Qje/RmP
u06CYB6r9nQ/ppuv10lpzl0z/X+zQ9QjFJyb8T5NWkCH5Vv2wxHt/fDxqQP3
2wHXLLFlUtQ1AGY3u+W0aL7JwJvpLhVZYoirjHWdC7eP0fHtNuPCDCwSSsnK
grOLLNOCuUH4cc6j555f/aaw0pF0JnKZycpieaUubnHzya09hp7pA7niWa8P
ppOZlpDn8fVLTZDx2mv2Lp9SK/R376vxJ+pBxqMj1/lEF4/Hi4ZjvHbLiugT
HiMrVBcXk0qKSTtrQKQbqWpTbgA5bd5uHh8z2y1bHuQePAaIwN4oHrFrqkLq
HIxamEesOo1Jbnw7a+K3W94ClTqa7TSmkHr8IWjnTBSbSNAVpMJCY07E2H+K
pU7p4sHW/ckGOsY+uyfJA1Ze8vNkbQnZ7Bxg5233gFqqcw1J2dvfYWwPLHjs
4/pRu6cogwXC6f88yxFg8cwR6WAC/qQbDB5tPSpGhFS2XC3hdprnXLLVIh7E
4hNPwjm4kbhC8EkopS5CywQTzhgMlWqurRcSChqWdWGK2dPhhsvhqasHSN28
jTa1ZoMhtL+7HS9g5ZqF3jGx9zwOaICc165bxrTEw74+m8jhihQ8Y55Z6ZZ5
ao9l+bRqkeUZlQfL8j/jC8x6wYFNciCBXOKIv7YDN23dp3dpDCnkuNDtEpX+
N++AXH0OWJMMS1YClKoFt9+/VuRp7vXonKMjhf0zr9ePC8lBktxJ3gKuujB+
m70oQ0OmjjkqmcfQo6/LAWBEpWZoP/sb2Xmsh1M8soi1gtS/qNpUqJIk9e6t
wdjOA2Kblq/eUmJ872aapm2fgjiQy6tLCdMaYzfMh5+ZUtAMl2nfv9wrPI9s
V9f8eg7WYpokVJe8+VXe/EeENmVpWymCiyFeIkVr1oIDkxxaQiHileLa8hKc
HJ8O0wKTxy1jJTBt+7jr48alN39/kmNMbpPrE8p+wDCEC0ikZVb5uep/yPEO
44N8mjML1Feo40vknQ1/mQ+dsGBQGQ9tA9WvTBXkCA4dtVC0ON5TkKY6B++A
5slXJtpjLnKehouLIT8FOMUyuv3cG78M0t8jcJBZ3pXv4AUWOI+RIR4MBU3O
Cvb0W2F9m/WFOpOo8SVzVBW6AXeRnIZ7GgoqST7bsBvYLfjwy2KRRecTDWQ4
r4LIji2VLk6g60q6zcZfq86Z4YNsXb+bKentuhIGeCe8PK6+2QJEsLqciawv
ZbEXB/mHrx1XUgfxnqu8uK1VgbU938OQyT0I2d2vROFXYH0McfV3mZd5JbDM
lGdx+rj6bTLXtq5TjjTC9EE6r5jSbAEXV6LLB1GVFYf0LKcgTJTeZjBC7Wf6
m5pMXfBL+K6L/kJw8AgxFpVDo+X+RpFn79X26ntiyba2N9X5jPthUHxC5gMh
rYudFHuf7diqyTpM9ALi9NUqxY30xWtj8qE27QmJBZvJh2xNunBON79tvB9o
7TNBKdEO/jGAuR4Jltl4LdpcIc/rn/YBG8sIR5dxjfOPHvQn+NyXcjOfIUOi
NIJU9d5vFLsoTk7lM7en4x+6oc8OZe9RIP4NA/4s+R04EuPQumEphten+ae+
gIKUgLnCrcMsvCQ3dhpE/nf5DB1nTUcTh1nuezMRQ1BSKaEo/MoL+J1DweBR
xoiyySA3at+D+jniuRtHflkeHPdGNzI+vbY4Bmo1EVzqJ+ZOepkptXybxRGN
oh3Osy91/A4VFQc4JQ1wWpZjJ8bGeZoZ96fH9jPDCUQxbRF90PgdeYaf0WU3
M+nVYMynFDjib3MdoWgcP8ws3N8w9WoJoEllPi4NVRhGrbkZp7VoNK5b+RZp
iUFCIh8lyIR/T5ayQzLD8k17/zg3sShto2OdU2w9HziFmuni43hE/flT1/AJ
O+ilU2E3GNAtgmjodnCSEpKhZiVSFk+wAnkKnqNRnaxh7CbvUJiGHWDsp8Zg
QN2AghcbAaAiKPHJslBDGiN92EcAYKhsomicNJFWiMFnL80j/YxyOJBOK4zv
dOGFFPqNoZXAaTx3gOmGyx9KVpzp8uRB07RNG1KhY729c86X7e71GOL0rnz2
s9rkWom7B3BC47JgeRnk4qQpm17GB6ri4Mviv23vZ6G1m3Anb1u0c1GkeCaX
mvv+E3R1/JbxK3jMb9oHmXhX4cXvnI865da21fxetiYEv0kK8RcI3zPFUwA8
ZTFVgWavPqbrWhDUcaxaR5wdrd77CatuipefgLM6AoaFB9nxZNu4RoweEBH7
tn18sy+XdslA6p8bfHDahDtlvL2O4Nx4zbTn6bdMtHWDIu79wN/nwlTVcMee
qvSoZ3hsHhaJzF+QHylSXbehjgE1eQ0KHcD1BEmn5fGho21ah1xRzixE6rV9
iTig3MS7OOwSIdy10LWhWGbB6UJIBvBxs7IwCqC7mE17y4hHr88ZT82qXCUh
KLZa+6hllSGWzZA6U/zkAH2k8WNilybp7WfOLnaGZZH5Uz35rT1gnxefdpAn
i5GB96YjmR8bb97XkdTZw4zM9UmlrEGoXElULKQNevgiDIRsE6XMPetaa/jH
lvVhwKpfPM69m/B/IV86ooH4DpiI81HycK+pncJqh7Be4I0N4mggR931fGFA
W5759cdFOmBXnmsnMRaFY+XmBKG4I4oWb7XeOjwdHudeeMY9p34pFgIRF0Ge
lINq1uqjh9hd0GoglA3S/BJd2+0I+V+keEhM+AZvCJt5toCWg13jNjxjgys6
eoj4ld7PhKF3L2VueSyYJ9iBKtyfmlpiCiMaOxNAqT2J/4FUboOTKb+HIPlH
uDgm3fKtNTTcV1Ppkeh65Sq1XUzOQhBhNlY99gYtRmjDd6vrQ0OhgrZhu7Xw
fsfKjtfa69ZBn8d9iTwNe5PCbBhB1u/5Imyb9DmVoggntzT3+ldWrwI0dqf/
TobGjSfXDNcnFUac8CYcdhSQDXJmvGjtKOpdmLLQAfUREIpxXgCtallg8oJO
28gq0/UYIgcnT3eBPTQQ3rXMWALDVma/2+uG1VWnqnQ0lm5vIumMSDu1CGNb
e9ZouOZ1X5yCYCccArnNrhnniHKp2kKztPD1L5gR4O7ROG1kT4bkHGjU6RcY
wbCuitw8M4JAL1KIF491YaWR291waIgKswQWKMrL7WGlQ60aWqOmBgBwM7Pv
0ESh9vN6gtnfwG6F546/LnIMoz0UsOKgYWAYWE5C1t9jcoHh18Da7dtiyVKy
+qHZ/az8ux7KL68CFLQe1S4swuZypTx0FkydNYCYDhso3dG9iGZ0/1Zgpk96
CyeRSFoqDR0JM2BPkPzF6ARpW0ktf+Fun1PKEnuoWhoPwVnEqTncZlaHVSYZ
em81nAsgBiBlOUeu6JuCYU4sMrHlTtPtTArypSpt1kXWyJWEmW6YYdQSgCjq
hUMpy+JiytSdC+Oqq3ZIlc+S4bjveSpjUFSsJudXs4iP1jefKFGkqvTy1kFb
LA9qP4k0qElykt5+Izx5uNI8hfYdtc0+wn6vaVahTYoYPUIqypQeEWmSWSds
0z6ryvRPwt8Enm7ICoteC7H5C/JlIFSpug41LEaeFikEsOzgmtA956HJQ/O6
oLArZPtzquhmdxrJmfJg3/1Ulm/cAzbIH5oXywwpoCCV8RTrJatgJ2rbQccw
XOy/lczEBj9NnuQyTVdj89Xt1WLpNNC8sqBUi5Oed7A6bmOa4pE/IGLX8FM8
CdWMfmudMa6+9cFRpe6u0jCmRV10o8ebYKzFrzGAFjzVe5H9po8OoUDFLXnR
qR5p0XcITOfYrS6BBEoLnsU5JqWLYRBZyN1RszB0O0JOM6JwnQc/D7q7JJG0
jYdjIaszuEwhI6h7edhkQ7oxr5ntv645NIRndU9N/16LYQ8pQ+9dWVOi2MUa
81RNK77UL4N8y98OegxKyX8HlTdXtK7yJTmTT2Kwhr9sOif6wDNn+0eeKhCL
Pg1tLJu9DavhWriAGVwglHYm8K9AbsKqY15c0Mzrt4XN34eFyUuaYqdg2pi5
F9jbskxPEI71xdZg/2YmiBkHln/U8GVIHECDjUzJHWMxuhlXtV0yKQISLMfB
aCNUWAi8HOn+finZzTMIEUky3sV/Uf7FG2FXX1uwHvsU3+X8Cj719KD0jyAR
FBMntnL6NmOmpZEh+6K3QzWCD+OnB3S4QCsM/l8Dcx4WWaDzkas8LiztMtP1
vzQXwb1utUKGlSYz2auXnqixM6lpuc4uwHpllccnXDymehGnAZ+Mm2K8ztMQ
HwGEeSHGG9vG6Mq4e/E1NrpLAmmWfpYWnqLdCMDEfOP0wR5TWq+TszafEu7b
PFLVDtYvGqz5e6DAHwXet39a3Sc0/9+mxAnTKpY+3taxvKyfIBtZwNeYSXTA
hAJGX51e/u6qlB9+Pu0mcntMflEKTxFQxhSbGvSUK5pFH8kUzV/rZnf3yBKY
EaxuaOUgJXIPlcv6QHRwZPDJrowOqMyPlFXeym34tmC4nCLIPiPOzmkvGXxm
vV3XkIt9bt47TkG6yENLY7rPW3TPsVRpf56YpyZ0BQSYCUppn8uVNFJKCt1z
1TlLYC6lr8266sj1E0CDL9zSra03Vf1MgaIE7IVImQ7bUtRmdxe8E9JUi+bR
nFYlsAlM9NYDdw1mLwzaZwzT+hbiStK8VSpHZD3BP4+2A26zgTVEhQQvQtDM
K29u9itBbcGS0Ri5Pdy+DbqVOlWJu6hoSWnY0e0CT2dCmLUlxnVjXPy8EM8W
BQ/YPhMFZjpirVxKlXjCm7vqWeSa/lZFHNta85Y2GvoBKcgMk8ZZlpGFq4Gv
MgPRiV4biZ/2YHSrs6rc8wwIs2Mcd7IhK822f+6EgzGx4DTH73xVrd+GTFET
2ebtBNngMNtUP4NLwbl1efQYuIgH1USh5Vz3ePwKUICY7RUDiRw3nkky982Z
ONedHpPny4rMdBXmmEsya3OyQZ1ILBjhkh5VFP8shUvCAJwCz8Y79Ii1axo0
QgOU4xOYaP6Mh64XpaeYRxd7+UciC3MtqQtrmdDo2jO7u8o8Mkcs6TKfXTWT
swEuNk7eTAGfiaWIbpaVtr2bpeF83L3a+3xKT5zcMRHWD7Lao5WQp+Pc+Xat
2uOTOdQdsgO3hFPZWIgo5wkUdkdj6USRoddakWYZAQ+nKq73JkitheZ63Rbe
7oB6mNYb1AtHZsBaFB3sV2VhKdCjq/uoJMOQ/CyPi2maxyjl68RhlrYyUCfo
4h1L382VZ+GRJ/4GH8bEuAzerNv07z40SfZ4NYMn7NCusOu+rORW8iH8F+qW
0T6dfuunKRQtysjHuIoSaBBOVgEGyvB7jC28Z2/biTlq1x+r+euBCHqfu+d/
M7ATkzLr4+IzxarX7VIlhqpeB3bAvKutR6I5sLYsEZqs+FHRsJNQs+0D4/ze
KiPTfmEdvQ98IPnMKA9gNSqeLo2AIPp5UVbSUtVq/sgPYTA7VIGFbLExiv8v
xOhXaFnNu5r9oVBqdzBNRlKIe/Z8Dnpt0Vi4/pvv/v3AhgmRzn7cvBPHZvRC
dqz1HHFeeW2sWtybSjuWYnWUDpbg42PJ///ohsQ4XzFQ5Xfey2PZ+NIjytSm
TbPhbXLQvE9onsu1sRwW8dUxFoHi0609GbbXzsoIrx5FxtR0y4h71/bbLx+U
WYFYhkMHQM0JEUxHUBvwoUgAdPt3h+6anVypKuXD7w2jY6vobd69CSZRI7Az
XgpJ4SvlP0vQ7ni1er6aiKWmlFZ0iyBM7OiRb0EQZsXvLG2pRzD3GFG6E4a+
00tjDJAIrw6l4aRcaWLjcxjZ/rgfdhFJZVAT0dmwFF+aco06MkCJ3gANrPrC
c4SDUf3f14D1ilm60p98mzYPyIV7cc6etdWcFId+LyKKkIIDmiviTzzZ+xri
FS4oNo/9Zn2tVdWfW4soFOOjHr1S21T8fbSr+EkGQNbN+AYooolqS7Vlvt7O
M75WbQ7QPlwrAhL6mT7DKCqLN4ORLCVtTMhzhg/EaHgIKkL8h7sxcnRXa84y
6Uoy2I1v62QhvvwgW93wi0qiwyQxH0EHb0ugLhATwYS+lvE0mnO3i5nmJEDm
iMhw9RsbsXhi+I1ZXUPef1jiwSGwBTy9GNe/+p+yOGT4JuerJa9xZnrBEhCN
2/Y6gH90wUeBkJfgWsuK5/xiIw46pA1rVHVXfXOdZ7ws3GuYzkJ4YHSi6PlG
PnSGxeBMt8CrPsTqs4BSETwS91FzSKMoTabKqkrCEDIy2A0PcAyCAmhduFHs
bI1fEuyZw7YbmN4B85dmUitOdFQoDbpDOzaW6LSVQAUlqk2T4KOGVQzWLb24
PPrkgVcQ9bM1rhu4ydbmMoSuREto234e/CD4aij+tDfjzOWrFCOp2ceyqJYp
sU/Md9iRka7GbpYz5uT6+hHDBbHla1oVmoWU85FHY9qEeIPbjiEcKz70r8AH
OYzikTWGFTBegyYAx7lpe3m7aLvZXPQcMukrr5sfFoEUk7g6orAGcAkZCoNr
3mtwjtExPYSaXRj2hrVUXZ0q/pJqMyblUUX/NuU/J3CFhPdNPJAdvBqzrvtP
0KU+ewjarVgmsRn5RYJ9JkWJc18ihz1zU5x43GaRDFEtn2XkMCRGaw26lCX0
lgJSxlUzxwyeVl0xBAA6dY6G1UahwB5Jdm+7onEQOIX/4qpEb/OWfSzdxBBf
8DUvrYVnA9t0RxhCVMaropQFWC4z3w3/D5lpCutuax9pzfE/HYV7xb5sgmht
RpId0jv5vY0DGrtNC/KXlKJ/bQJy48+aRdKFl9S1tHajhdZRXL7//9T4skVs
klaJPVCTt0ENGXz1BKYG4GF8OLaGJ2dLkwiHvB4HqhxwH5bHqDfeSH2ds2Wj
8fclTKq/eUFzY1BnucC+Vv4FhufF+GavXiq3dzpKTpaSBR24pv1cOhtfiGup
5O8QCX72PdNdBe6DTa5O2y92nx4cRFKdk0SSBb2dLquOHKuKCTrcBUecs1tI
YFuwqnhLwATOjYj3V+SR5xOY9XFZzkBqpBcQfvmgxIt349c8qbWXEInWlNvj
nmbxt7gY0Lufi3YO4g8voRgM2zeyNAXe3QYjKKuIUNMSEREeMfxeOJ+2cFNo
kKB8kiQ07d4flYit9w6pWK7lZnTBvqWiGDXTpkolGQO8xUaMxdHqb1BsHf1o
BETCRyYr4C0ct5q3AXDwsnGZ2qEouXd15RZ7NJ33LgGi6vxmmPH8QZF0gRAK
9jx0NRRgkU9J1xydzag32O46etRWqbmLCWXV1+G3XU50SOu0pPW9hgsZrGfJ
bx0j6jFxkpdo8xkkQSPnVTk3OuUYiVvHFC957wglOydxfeqhvGyaapgg24CG
hz41RwuEPUCE2ulQvydnC11HkYF/gvKDU3Yg87nlaSRBZaPDzoJLf4JjMrqf
rOQCPmx97gJdolZZ5zbtcUnvHLVFVzio/KacuqToU9EPMJXOIjF5Jt6yT2Xz
uSVxf21jcrk0RF2p8K8zVStoWLqn+WOkdwVpmefMst13N7gPb4BH+t0jhOc0
FVqRX21V0N+RvD9za8W0Hh+pwBugYiSF7b6hYg2V5C7T2kX1nWBOCEk2ONvL
S30FlUJR/lGwowOt5x1wMa0G8CKO74dsngC+sF/1RlNw77etTVyrw6//ErDm
mZ0ke4bLDNehbnWg7qENWJGYa6qE9pe7pa19VMVSY1gmeZwOXF3iDLt8Nbrj
Rkum/fa0vQbdnfahFlVsppGyd8UVqfPz3aZjvHFbij4jVt1TIoLKRxLeL1Oh
r9Xb57MKuU/ub2hGvsfj/SAtUo0FUzb8fBU9whtneYXaZLYx7zlKdtVvAMCN
8MZm0pFJGdEwjPvltCU6BMibZS7DlpPXSoAaA9u3vE3jjEjfD1Wo23KSKJBP
bTSN+y8F9vM8/3k3ut0geSPuBQDAf2V9b5dSyG+VGmEJegyeq3nJmXKsLxT7
rQhL1bjvhdeRcAg9EDozhdrDhtu7DUAUP2d7jqTCpTlxSf4X6LizZihTBjWu
4mz5IAA5M4H8vBtk8XvyBa5Qn9dMfyur0zbyUI98FXfXbGYgjhgWp6tOStml
OICRbodVVZloS/bsrNSXqM7NJiaUKB1vocPudOLuCUgHxHgDEphGHBCrlaKb
TBzkK3kvpNe14AVemzDarFdzKFGrPxbaCS4M0wPVme/L7IlHy4rrfMGh5QhW
RMA1F/2IBFbLlguQj/kFT9IA6VB+OxQ8b0Ugnl7pBDXE7AM5O+2ruHBsBYUp
CfrnYD82URhWwk0RfrL8GocjsbKWNOB69lbS0vUdZ6JkyUzWddORY8jleKM9
b42BR+ZdF32t9eYQt0T0W4fJpNJY3Wc+cunr0X6NQz1CgRl6d4ndKW2/fiau
iIuYWEk8hY2VjuSH9Ufn8GctHhm6bC7uZs430Snq1bJsFaqgirLiRsAKTtnh
dckomOLVqqVcIp8uos4D74VyT1g+YloTfhpI0SfdZOkUI2a5edMXvPVSDEpU
UHV2shWtHy52V6ZsIMq22UdAHO1CI0UpyxXd7UUBu/6vIHfKtbMBWgg54FAy
og5BDXqFuPvpsYycleWbbJfVAkt98q5Bxi1EGf2b+usCEl80wkw4vbY4u1jm
sW3Wb2K2Dlt1w0JUchD8DS5EzqgJeZUrwOl1LNF66LDaGd4gVndug69Q+xxT
GEZsaGmEMralM0eB+pgx8iaQ2dL5yWDgdAFwbn17OmT3PiSYLBvQqGlHrBJZ
kVReuKac6mVySkgJ2bfxzvD1IcBGhD7MpZHz0o+FSKOAqHnYH0qI7fJ/J//4
0Eke2TiojrAlUNGFnFviWhBBDrg4AGFbBMC0UYHlq7iD4IqMNmCHrTQyuo3E
7PfqIZrE+Zeh/hnCqsumfN8we6K+7seCsMHlD76W3TI7yMtVVXrbUww8UUAs
xVl1mK2ioguahFXIivHYbe3wPCk3oWK5AEKJwe+B/+oUuRxPayo8aJhsBLgz
eVxlD/IS+KSRxyHZ5EQzcWj85xUQ0CsP5vzdvdE1kN+Uk3wmj4TNCRpjNfXG
TrHrc41hjncqB8tlMz4zzk7X0DzI8yPBxArvYEwUBghDWY2NorW1O6Nr2WWJ
GGCKFoODDyefG1RzWEZh9lWGmsticaBlFgM5turDxZe82tXGQJ9s60FyCQfZ
abApFZUJlPEHFxPIWtGeRTi6BUdR83HZYFnFQdeEiujdCz0+3OqnOTBm1NVE
Cqhmg0E9hs7TBc5WbfNvqJFPDd/3QWYMBfAWUsULF8gUUuztsM/ktVg8/ucr
Mf9NrvXMFWQaGwtvK5Xoz9flsyZxGdlA7R5i48peqfmFUe2fetEuGz0j8dk3
kGHdilaL8mLsEFkjaw5ocFpVAia5sZFkueTpHzRqLQipiVP+Mf1v1v36NB2M
GywDJsiBvfW85wYxa04ay2wg3rRtkXlDGOIT26Rq3EP/SpPR81IBskNAkKDP
ueHQdU2ZaEjxrLn3MENX8/HXSM4AUSR1y06gHDuiw0abrQUPkukbl9fgXVUA
1DQKX16+gBO9ypF3pMzayRVbeSQ0m9SpBBrE/PO0w0g1EjaB4Y4qro4JZI44
K+1enZ4GRH9xhe+Dks2BLkOyM+SvWvVDFwwU1zH3hYZiJ2R2sC8cMc20WrrP
KOu2mvnUxy8zjaKz+t66cEd265yIil/hmtoFcBtpOmzglb1ELXo3g5tUs4n2
Z0wfEwsLtgJ2r89zkhBxByFjH9Ks+WDV1u6m8EfHv2enyGQ/oXrxLKKinmam
/iUD55YhE5liKaD5ucHhG4Wm4B0r2/GatsHV4BVlxF6gopgldM688+MYK3En
LkT75vwkhyfshBqFlrNMaY4ddGxn2XtJnWPo4oDHQNsT7XsaDHQBkckH/bdx
fDtzj9tZJKDQSNzF52UZHgLE8QZDj9/IL589hG2wi5rUh9oWEEnsMI0B/EeE
8pfPwBP50URQgkW4W6O6m/jDAt+FSIsLkMBkzGn9TKi8S9s5S53G4El1AP0E
lN59TSNX6Bfl+mqMeikb8vpHVUolOY1l83401U6gXmvf1CrglMqwMAfEAiVV
p1rsInF+RoxHmU+nUKfyRBMzHPgvpkBpotQoULOJd6ZnTM6fL5+Wb7CiC82J
uDNSRzZQjirR7uNjND2eTPD0j+NVfrQn5BZc0t97OIfrsGV8Am0zI7DjpSsg
vLrnKJ1UdcDgCXb2UB9b3U6HuFMFyd36ix1h2j0cxQ13KEL9FI/dkXwEAeBZ
zbHQWQ3iCaXbnlb8r9c/MgQaNzur493l6ex81IHChwEonpbC/JTvHoeD89ZV
4+C0+8MSkVYIqeRWJVDIuStJSsCivU5RfoVXAXVWj6JEO9S0hXShOC/7Jsox
UO4uJf7WT95NNN4T/yEpqyWPvNTYbxLKaLMCOsmGiqVjouhMHcmTR7KaiUa8
Vp8SkKE7rd+kouWZXPtcz8Yg5dzXPA/+m/SHsXcPuc5FG0ySl/wDI1c9LCk1
Pp0jashLFKf9gTeD35QM402n1pP+dLgBsziIJZrFzlHhO8jYCIocTo6dBAeL
HsL2Oqa3LJAtiJqW2fnvWRLs2U+Ecx2TeZu0xOo3/Ujw5nhB2JVhec4dkAUw
EDwGBsE0hUKOHc0jMxdYZg/Qdfe+sicJ7xJo+Tm6BvVlCIAJsndt5C2WP6Ct
gG8KkkgPTuK8Uy5/ssP8pGDO9SBZ8cOtaK3Lsc2Jcnk0BUMfNYJMBEDBI5X2
MRDmxcBaoT3yxoz9ctUcI5BJ/iFamlf1HjfYrX6cEZ8YbWLNd72UwqV/4OiA
EnSYQrRON/0ukLef9e2fcvFthXU1DO2trErwurNO2GfMSmZBOCQijtt5DiEZ
G99MOi2kgB7Bqb7aTnYOs9niRIYLzPpFpZRGZl7j9LdXg5hSSeGk3xV/UQGd
45SZico6s8KYBGKPfAYCtcNBIdfOPHt0fj9vmFP7ezRlTFFfCGoJ2uGJqHm7
cm29jFxMfglRGooN72zI+kzZXJkU1XtxAHdfaulf1WoHaGMlELY+SiqL/woJ
ItS9mREJx7aV4dbEaTeNhcVsPvGFyLOw96jXQdsGM5C9WXGLz7U2IU/6oHuZ
2Hd9S5ZjzrKRk5K7qUmlcoT6NUe5dKTkTcIRr9xtllUssnCBewqb4RiFauU0
nVp3rVJg8QCQM6ZHZPB2DoOIzsMy/0DXzVYLeqiiAIVCkEC9bqI9wqAO8odL
KUQx2EMdNjGPSn+drqJ0XDu7y3t0+5K1nFzThC0D2ClXXEvMgAK43pfn76xr
QpnUv+KJ4UQc0abOdsdQxtZlmLo0WCEC+jVYvnQLyxm214xl79QCpp0RyKGU
El525em04HbZN5Lxsm8kQjtMZ+SVbtzdJsG8n5nTEjYp1QJv3vMMgb3/xHFg
Cp99jgfSBuzZxokK1iksAWOyW/F6Q/x8Wc0qj9gc9sZHfttqyJEUjwSIsmWR
xpmFAbGo6CoFbU/CFOeGqKh5U6c+fz+M+VGJUiw82LpnPB9Doia8PMRWnvtt
C9R7Qis12sjyMwdbruvIyw6+rzTSa0X3RUo9K6RLSaUx1MxDAF5Ars5UGMIp
sKvXA7N1/gE18yq4bhpIXHNb2olwMmORQvzeL7NPKUOP2bCxXcicTFO93cT6
v86banWTs16BXMt4WT6snD4mZ4Sxo9HKcPf+35sQ8YAoYyHRcatgas67A4Ix
7A8b0OHYiFSSRE45FJ/IDgWf9PhrQttFljZ7DOVUux6kLlnuu0mqK1udYIxt
YNmfhsZ//aVHcvFQJH6IA2AjuN9ArReT2kW++k5q68+bOPxL5fD7z/cwbD6X
CjZMeHyH4WbdlSbvmZ2ur3RNHqwVbUaQe0Fb3tcNK+CTOb1xxfdIclmyHRYV
aoEFG/tkJ8qTfMlFWTExTaMYPYZqR9NKtsg1lZhFUVzOKwVkDWtKgAESTuWe
gmPay2l9Ax7BLdg38Hq08qj6wvTtEX16EQu/WpEm43ya/xcWZTjs+qMSyRrF
nnWu50KYESGGSkGxMfvknmaWlQ6uCgvmGuK+enzEHMkBMQ98ChoCmTVY81to
UUSXfqZCpWg8Adw+UWLiSkWZH7DpOaa+sDX6A3HkSncDAEEfVQK4L9b2RleF
Vu6SFJXft59XscLrNaI6MFlRwOZR6T+BkwGH0zXLejSUE07ECEYojfe55Clz
J73ePikc8zhuOhWfWOmDuEhahzJW9QOBRv9613OQ5zz3SoKVedlx3wqtUDHE
oxtqT6I8rUgKWQ1FAbyq3wpDu+lnITxlfkZ9inn9MlVUKUHuz4zM5QkEG2E9
vkn/9kwNKWTETYaxP15JcCdR+bxYLkUIPwjqoh35rdL+hdSv46PQ20MqQsDw
V19MYTPiojoMG9V4U+m8Uigyg+35FdCQ+UWPKbrt3sdfQCSjLSBuGnLfYAn2
8E5Ff+P0QirGRulmwUo/ebxH+YqSjdLCO/RZfnF8otQ4tVQCffwsbjahJaxO
Gq3gU+uTRAyWHprUOV/HMAxLrKhhgdP+I+L0ZAd462xq+5jiWIT/Ot2XFGIr
idyoa5cVR3RFaFF/G+L2iQJ0n/VhDBfplBDDa8tSjxTL6cMe54ZTsUKtUm/3
4YgYigMA6kvlnv0n2u4akrtGA0/WKeBhsi9pMZLiqkwaPEbr+c2P8cqs4VsC
eU9un9LKECbiD078OW1hm5l2UqvaU5+Jq8KYi+GQ6wcc/WYfa0vAYgWMIJY3
6hNxkZO/k9SNc+PFyVPJtmC5wGtb6j2BgCxAqdA4wgHPqF+kq1ZC2g4srpgd
TejKiLLa1Gc+Q6j9cRVVZuyYJbevUJpaD7VYv7tSK+eJFrcfTNWdQl5JayO9
OdtHkdKWer5fduAZomQ7LAM4bYZ3bjg04znIccJFGHwbjnCc66B1GZss55Z3
YXki8piBCmPi2qkcIZLtESiCa+9weLly1uVfzXhKzNb/sdjTEKCsir/zz51l
7md6ofoz5FT/qLdLl0GdqN6iFkf9s27UvSR8knCyq6CzuFges1Bo9y8QN3Yp
AjUHwO3FkRNNbyn6HiR69kzosoHa9jEdpE+wD9LGpC34+N0o8PD/sIezpVcJ
Lfo4ubQ2IaaYbA78bcmRpz6MyJZAQvJc67HS/Tfst5o3gWHsFjnSkLCQC3Lp
ds/EWGYK2rRsv8Fz75IC2iiAqjbjLa1c6gCEiCu2C48UpmZYJ95KLDPrOHeg
HX9Iapxk47L2v+oEWWleDiQnHiAtfZQ8FgAVmxbz5HiOZ/UnoP1SZ6oFdevu
MJxagI3Satw0H+T2ee46xQbVlD89/GJcQQ6lFh1BYKKQmORoYlPC2gmBSMqt
LUNo91QYP8sLKE2KtTOAMqzVXQvNHJKzJeoe99u7p7Y/Mrp49CZ9HfAIa1oy
wvB2AhQjcN5z2EdyQ1OFdAfAbV/5eiVECGetfcKfagLqgrdXvs8R/EY4JpuG
RcYNBxbRgf2ht6cWzKxKDmgvVjlWCPABCMaCNpHr17RLbmOPuxq+AhP5pRvk
2hrUErRd6bllKYmg+a4vhMXm48CzeI/HXhrhGJuqOap/FhX1kOhzGePie0j/
eift83Bln/mnsxHLVFQHr2gy1XFVIxMQ/YoV68e9193O5U6LltYeMdfJd1Gy
6Wzj5qNi1OsKxzKKeIoZO4xfOeoDRvLmjKf+/WqCDoHQT36ZzJ6+tV+UuFkm
WL1imcaWVSNbF5zfkc4LmmjOGB5ZuIT3muTMWk+pDTJVyvosbbPisJLdCFsl
V9rCiQoqiss803gJc6p/YjRYAm4QLpynUkGk1MAMkFsFTzIQEVINLaU2oRlT
WbwcsNa51SeuNCILiswGy9WWPT2PkEPJ5d/k80H0kkGeriuXaZ2moo4Lo/bb
5Bt/uG0Nrv6dUAkl7AFZOBzGzKrXwQ0+d4R9nE8oArNSZ3tx3aBjzfP6MpD6
wCjKnMjbiQNRjNnEb6i8QezzYWFzy+HkvP/oByR0FPPBW0UU8hmXvQj8ga7M
9M6RQpdQWFu62Wwc3OLuoW0fSW+6Umdi1f274XZdhdNnNKBPZv5cXOGtfvQQ
EnnAEWWFlZ2Tz2gQp4Xoovt8SjJv+L8KtD3yG5znbLQpMOwzAo7i0zfBwJK+
KOLBV03VdC+cxJwJAf8e9udWx7aM87EFJIp8PLE27oo4xWX8lTSQj4kzJeh5
aZzLGtIGVdPcpOnuB8SzHv84sVPhLxDZ/F6Zh9QRW0QAWWSa1pWiHr/3pe9a
M/SR6yr4NTBGRp6846KxGkRvBcKeVxLbBQwH++Regl1Ek54k5jahwMll14Ls
hnF4T/OIM12QZdAEuFyBGDo/zP6/p11iYWTM0DAZeU2LMnVNIrJtAwKh2QuH
i+yPVGhYhW6i2UpB76ZhddnTm+VQ9iQSLpk9P/+ZQFgwzZbJ5g80HFN3DIHu
KEVNlLRASsQBN8cuJFRASKNFy5vD8/LiJW3fH9RIAQB9brD4pQrum4tAK38c
n8JZD0dQxlXb6sW1WfK2LzUjx9WMrMv21x98dCPo/3gI+tjUfE+CwV9PY7g4
BGCUVnx7U9wPOO1g7Z1qdbLMaIFkWjcHsKfVNPZMiV7fFlp5LPCdkhqA7kDo
2DzkeWnRwvygaAaSpwoGNJlra90zpWQ4BaoGEJCa9lDmQjaIOQcBzayuq9x9
8Vzq1VgZpbG9qGN7SI2eOo6JV7Bd0npbD8xJDFdrDMPRcypcABBTzzqSNbQf
kr/ciUpuBkmZH17UY2b4BfjIsqbGfuJoqGFgcbZxVQHpKkGuyriJTewbRTqw
I0YszGGD/8I/K8EWQplWDtLn9yMnUwnOaWTeXPwknfNeXbz1l8RBtEN7+GYn
bIhJH16iy3xuc+K2Rr1I2rY3e9whl9KVqJPFqB2hcpLczIkz2GHbsV6Sxiu1
GYdCmCnA0Gqb6CzYZpTOJ6xQzUgY3lXILtCK/Gl0jxl3xnp2iiFdqLcFgtNY
rH5TFJr494MPUkLNtka9T4QzWl2zVz7AF+2lW7RCDvE40dYbbjSV4aTzoBqa
dqRehyXrhAhNYfKxTsAL4DlXNkU5srTDKYsUxV3GDQPvGF/xCcMqNSVF0eQX
XLglY7372SsvAHIJdCpa2IQ5tdnn1jnpN1Pig/ODKq2ldNKPdx/dVbmC12S+
S71MaPxluJOuyb/ZMywesGSfH7gA8wSsP73MmL67NbjE4kakh2G3Sd6GhhJ2
A9Int8GxU9UAM/NBtvKMoCisvwPhYQdHmnSYGzizaH8FlBDR60S/yhUPTS0r
4la1RF5LmHef/lE6SDhaJNodThCEBKFsGrAOogUZFWQI2fBOv9BCCDM2zQA4
B7g8Z2rlj6wJ+/tAlp1TNfDB6cUMlX/J4LCTGLHZAdOLkEWDw7QTj496KWR0
XP6u+OWQcD4UDAu3IzHBE/iInqFl+wChBZn51b/FobRnh5iZP9fCf235+5RA
Zl/vlPbjJJwsiaxNsqlKp6yUVEEkDX7CshfZTdRtSxbyDdyF0xfK8mJKiWuv
Rj7j41Wl2MeNdJ+/fZyCoMxUdcFQrQXnJLjG8ayQibK1SRGO1wfaKqvHczAH
snJl0/FxQKQDuY0lHQRjuFpoL7ref1oudfX3bjeDvjZ3LNyAgMk17nrY1oTm
Wvm5XYBlmFn0A6J2GJAOx9at6g61x7ZIgpgBiI55ebGYHZ5c817KM8doKoX6
4lL35Ui6H6pzAceuQZGHTtIb9SsUtcoxXGue8Aj6AcouSgYRXnVnYIIGpyWI
BUvOSBIAsckw/OiCumGSViWKFCZxKgD3yMDG7/3sPl5jbkD+Kfl93Xw94tiZ
3wW1Htnkmx99OXACTJnBrJFxylSycxhWm4yVMZxWM1fHIlz56C04+rbJE9B3
UFCGTwb6e3Z1imyUD2TbXNgszR5IiePpMkYSxWoM+Kdu2Pf64jcKMkFzoaaH
P863F0/oZUvI3QKLdOXiZ4Rchj5kfbHhUgA3gP6jwqrULQer6mXMsXzaG98J
pU/PLyxUsTAsDllYNAB/xqg7ntXIcVwDXEy8iddC3aViRqBsv+IF2m5vzVDi
UH6JU2y7+2rYoj0ekxEkbG4JoqALILmcsIkEen+m79odNQfDhuwYdRv1ui/G
LnTUuhnJU8Ffsn9FAAGka1sD2BoMpp1TDVWczJbM14BZiSuiMhJM6uTKeWJh
DDH8W2Yx89O5jQ3w41lCJDXWo04hX4VmO/P0LeoSlZq9zdMG5aax7jN4FvSJ
ZLH+fV1lWWuHczjy1/T7h03nzw9EMjh3aVvmTCItBA1pDVhHbHBaaJSGuKrK
1OhAtaj+rkOoD6RuQQDjRJgA1ELg+Jr1OtBXcjA72UMewiTj1rY5pi9XSLoB
z8Mw0ypypkxJd4xLcnbCkD9iqFs/TzPDcweitPg6jUuZaA1ci1SzEIEQOpSz
nJ5X4ksHvCAhfYZ+4ZtBGlDHyUU5YP7+/HSGSzrqVzNGpPFx+3cLtqqNfT52
mJeOuF9FTsu/dYhJpp7Vtvla/p479jG7kx87plc8B5O1nBp9uwd2TzmX0jO1
txMIae0odSePKd8mGs/K7nUeG7pibpvH7p81XUGDdQtck/joHnqCDtlgfaT1
BiPsruTkSLI2ozFRnm4W67DAku2DHjBOhKXVUWqA1zNQ5wCWXzvJRpSAJszF
NQpjLqrjkecN//9efuhKOQIsXjh+V3dovSmpckctZll14QhVNHBgd9Iwb6e4
ReJmHs/eCoQxg+jTQN/8FdGiE5UEkGXRbqZ0U498LSl5F5RoHKNNfXVt/ua/
I7dSYq+RW2yxEa8LBp6kBDFgtt24q502m6E5NvrLF8k68DvgnRQxUwtsv/g8
X8ERcAyxw8ImVMPJz7BRHNkKY2Fg3i96RDHDyKY7L+tz54HDZPtMiKnFMVSk
6xnUVoR0y021prGxGUbagR+5n7dbmZyct9cj5T7Y3d2p1c3TQVgooIlhHwos
3XqWXie7+BjN52lwlRYQw9F9IFfc0/SrciZ7JtXlMNg5viT+mTz0dF2p1hxx
ljRIDKZztUfqD3r+FF1v/MINqS1iJiSnPJJYYMZ/JnpIHk3S+VA9ye8iYFpn
iIFuDry74zqvK/XeffF/QlQ0SqeAY9WYl3rfbA5uNBRXQZj0OK+e3dRqwi3I
OOubhGV119hU4P4QR6y/eyzDFmRq5RZti4dKlp/IzXwqAOr0WIMHaW5axJyE
VGT3KCv2Hwx2tZNQhKO7mtFNDqt1JEih5i7eoFRBag6RlO1eFoNUYvMVBeTS
0e9ANBQhPbep97WWAzc/LkT3Br90BMqFtSXId8DfZumpN2pV1op5DU8w6rXl
KfcIQX07uVlFYflFD+eINvn6n0zuksVop6lMJ8oi8klDdPIu/gpRk+9WBzSb
bDgGVE8zp2ASOXd6OabasoBDof6a1uesvFe5DMCfH+ngV1GXOQGkVS9iJaJs
y+giZX7GP7Ge4WMnR5co34T0lzTPjCZ89ScX06TDm1INDZh7p+CjK2IV1qLE
mxgJx4r08QwzgjGApEaf4PmalXRbyx9kCFU+jkPSNtzdp78dqfls9bciciS3
JRsv/tMd7Fck936xhvgOJmz9KBVjeUT2ORLhDnb2WfmV/82WPi4ulk8JmjMJ
aJNMx0OUyZx01aRIRZBZP//q2qOZ3omrqqbn3a9fEi3kzsbiZWUOvEpIDTYU
PAsOGPAYV1E87zg7rPP/zfvRhdcdGixDoiZOWzJHvJRuPYBzmjN46HV5Jpse
2Ky/bc2KdOU9Ljv5osWOtV9UZv6YwRsUXeZuUS4tDSqzm7tJtTWW26SQKIs/
1CaYPHo4ETXg6V8rHpH8hbHWp/0KLkIvxQt/e4OKyI0T5ix6FTlX6RUjhVMZ
5cnD1pnkJqG+KiIrsiq7Ft0r1OepUgIr/kNtmC8N14qFt3DI1U3F49lCuR9Q
DW4cIzUsh01plbXn3PmbC+W2TT5UDuO31kmIeEVhnmpIyjSz/tCoEIaGBEfs
q/AoFI2HyWz8oWDqM+FqMppl5ZnJTwG+3bkuhWb2RnGsDZdCXo3m/bLEpcGN
ZkC1Y3GKqMwKMROdUnvj2HMjAeZXw5qtXfFFCCnKcWTZWyyogUBRJWSrhI5Q
BPnnsY/itoUPQwv7YNx7yRoPoynNbTWYZpNJs3MCmwm697aeByiGWz475Xqi
jSwzeyQWoH/XN0V7ed1b14ubiUPLYA9zKVOiT0lb67/5oXdSxnCtR6JzrjJC
qImMua3kCuxVKbFtmB20riGlKcBuM/XotAqVK6W3ECMfjU5JDsqy/EPHHthL
aWCCNyvAcf004CwKKRxLdiDyDWIt+kBUzmrpv5qM5RtZIMKD2dsYc1wzD3Cl
MYERlYPi0cjFvu/CiQNjlaWCUiWQEg7Pu6X5JEH5ITOpNlXRPKPgbiO7az1L
ftgEqmyY8+R9hmulhMlYl6FJvRIDyXJZNzYSULalGapbrQESoV0JU8KUC/Ei
f4k2vwNY1M80B9L0pSpzC4rlYcMzhbH7ZdAdfgBAQU5CdlnsO5rb6xlGx9KD
uYBLibXHOX1RIfzm3CJGZzIJzo0rT38pFv/i8WyDQcqC3KLnIdJ/yG6Bvk4a
EJpyNzF8SgGTZL1eF6D6gd8gXm+iGRlzoW/7FurcooXV+T9nRLyODqbPCJHm
LD5W0IU8SRwDG873LY2cRybYPJQCWb/CMqKx269yjP1H168ZtbRaB5qbVjL2
MbBRQnRtVLRjcsr87WscQO5R6pZB/BlvTgsbgBwB58WidsEl40/AyRvpO0b8
289zmEhpuEE63DZUAPCXTj4wAXQ03zaxkje/mc/X9RV3Fq7uGoHw6jEdQXFt
LssNfNUV1JtJQR+M+q37nTvAqfaUyZkttol7ZHNy4yNW/mswREp8GBkskUSv
jgqDLKvmxtD2/ybEZ3FvEYoqEk1+AdRaGolleGd1DNQs8qzLJrzd3/RJcwPm
8blsjm+/s2WSkfsr83AUS8zIHeKY88ctzWyi01EI9Ka8YjelutbKbRAocpyx
0XpqwNVQ6AiAAw7AxuFE/90naXlv14Yq1blqqeTPA0qbflo94/BDhTZp8yF0
tU/YOTWLjo52uNjOroCuriIOhHqpvkcw3LIsfNmxZT/zTLxqx9JkEwNRRBxK
jrovkUxyyfstKG2/HM4glhms8OaUvZw6Y7dOswLRIDhzgLqqZ4VtuubeJgED
uiHGwbBu9OyuS+qwXmlO590/3rkBSqEvLXVARwroU4U6BesLqCu5WFriGvoz
ydKMdrg84r3Bm7HxLtIYx4jcVq6Sjctp8L2+DxQKYBo47qcQKAlOSPor/ZDk
+MaqLLrhYIFix/VB1R4PiGwitWWcIW6/4B0+xHKtbxDVMhNO85t1BilPhCZM
xDlHXyaxHUtn/Qa7nB3SAfG7RtWlecx0yoc9kU8h8c70FsS0F7BusoimOSQE
iOMZLpEuaho6n7dKA/rULT8T/Bzyao/h7sSnYzeLOTLqw8BXBRhG7FupkyC8
dhLzLMYv2hyFzI6aPkHFQ31K/hhpBpz+cnv1FQOGhFi3spd208f2/0czGEn+
6+nX2j7kP3+1mTFA9o3dX8/91ajd4kBPvGB8bwTJgwB4y3/PRxyqQPt1oEhN
vjHKU+MlGynuwb3uKLDZExaFKETYx2O3V/4gKY72xnkwXsS5sQFFeaCm717E
EWVn6th7BVeopT2RMIm0NtqNN+6PAnVHae/wdbZoedbeQsYt8joNbNrWMwxx
ooMYku7CAlJTSvuil84bPxEfPvDHhqwbobBz+FfyctAUgumy7YNEuddAK91v
mfMq6vi+IXSqjUoHPzlEdV7yWUuRtz0VYaA86FbzdpPKjenPx/ONyMU4QTAD
fQWtKI/sX35t8aupe5L6F+0JyPD3VMh31/ygwEJA22HLHEyeo+cOVqE8Y414
87Gl/2E7Zl3z02gQlcksdV4/7V9uTAibWFHFyZKHiHU6BhWbKtJ5xSsIDIbC
ECspg3y9bkILGNANXrwAKJ8V5l+rchP54jNtsrePqFt43Jm+3Yys0aFAcr8j
FnCTILiVMm48rm8ubojmCI6gpfeohwHyN6fPWBWj74sxr4ZtBLrBAjxIXgwG
6/WRaxph9LGUSzh1nP45+QKK/4hzKy4KOhydLqWVVKZ3xYImXGYBiC+uadlm
wRfNJeH7FFqKiw9CZbeL0nG4CRAaLpTcGkjLjWXV/lhtwtYpz20FnDghzKjF
vIi0FbRKgmAg8veuF0RITuX/Yb3qM+HuhXwflvcTi+Iz/Yay4xfMsJy3D2Uj
AsI+BY20Q4COpU46EZ2SIYJ8aHPiaYoCVWxv31IKRW1nhAn4q6gSE4O0VvXT
0TJJ8WyOKhEAY/MoS2lVyIut9IXvbYdN1wtbvHWm1VRCHHGtrdVQl+XnPmJq
HFY76FBoJ/mrU5fZcHmQ9ecsKFGlycv1m54/3oyGYBQ+NyuQ/Xgr8hmqiBp+
qyGwbZyVGldmIYseoMf/wnRcSePTCOnwWtJLrmkw7hmvUmOZcDqKn7dzbC+b
v46/zKJYWDLFptEpD9n4iadzXcgXMwun/REtcP93nnzplbQELdWAXzxiqp+e
2f/TMAay6JPCQcZf4U0zd6v91095/pdiVdvUXyYV6zeARi7mHKg+XMzIYl1S
yXmt6m0MX4A7UEA0MBamzhtvpU/4ZbQjf5qmRcHcG4A8UDEDnij4k9xN1foE
r8jiL8ohIclsZhrIhrWvGNFr4OrxHf2TJXAXZpWTUTqnIMq4pvrdIqLJERd2
0VXreMpeRi4LApNlhrt+uciW0ekf0qATapgCKDu5ZpGVPsXUg5E5Htbx2qb+
qTtEodsIU7Yp9xTxJHf+kdrZDKumymH5PfMcsl33GN0pakCJu71VeJVrvYgd
RlwXDKyVG6DHWgmHqupTiGq7lQ2l0g9Pj3Dzi8GCxHSLmfByPHwu/SGW/+5I
m03yk+WmoyT7W3xYLpV1Dy1AxQg+q4+ybUM3704tspS9PN9XwReN39k4ZHc2
Gp+vIo26O/47fLzYq0EQJgyKaIYltva/L4yFMsyKNs2AN29Rnro3mitNJPzF
xYusnNXHLx8epFhLgOV/XiXugcidLt6oongHOYvYPZBGmwOVluoH9564b3hc
n1Ngz5zjZ8jKFJPfx2pwub/U6Vq3kF+O1O/H32hlTn+yp9QBpKlKEjuRTJ4p
UH5ksGpd0NuI7gC68afPDsSFQYiZQVIPTMGC5BQzDGV/rXOpA3LjauWOPugL
4LXhFTKjVuYDrJLfpk36a0wUM5H9IXLPKvJ9A8gXiMn4QGYKHfy/x/y1faqS
jPO8R9/tTMMDw+IX5AgRJL0CofYXSnCe0H/oLhSQU3ULUmyikc4+dY17x/eU
PsTVBAZCtCbAMFSZ1N3HJZOapa/FrOqWriMVo5TqA+ExxOi7t3H4bklaWPy7
Rj4ZvAeh1NESth2NZ5WB0zmdXIeoehzGa36bZHbAp08i9eiUzKHgHGYF7DGt
SEb1icFqHhrI0xWyhLJ8YyXzpEa6Xa9M23n+xw05+Ca+B7frC3eYFBHk25Qm
NxCZa1yX9oNBVBwc6N9wi/DdJNXvhpY2lxcbWTHRujbxLqZtscS+jgIcD9vy
t7xeAizTq1MdAnG5vU80fgDGmp6vBsYtQnWlxilhZeoD9XCv2CtZ4D44gAFC
S+0ZHvqKhpyeG1ZEfOn78IAqwc52uSHPXKcQ6pLcWVIqVv1HdNe0QwvMIUCS
whIME995E2cpNPeIcrIAjGQ3jdz17MNpw/O4s5qKpZuhjhYn9bPa8aVIuhBu
73FiTbkscdpF2J5E58EfGWhFAXjrwW+Jyzag/CyTgmV4XWfmNvid/PwmGweZ
zobRjxtb31CEmPJOKFkmo/thWTFwNfKEgdtSnVPunKownuaosOR92CFdK7dE
b0YAaDFKgSrKMfylbGmWTR5wGLH8LJjY4H/pFnOOpsBy/9ZIIUQrQO0dI5k1
4zT4UpfbngIBmpJLHM0Ln2O+8pzjjYdEJOaMVU0BFZgtd3xDiAaXr+Wu4GBG
ST1ajCa8m7K5VhRHpepo2K0WTP9zJ5pNJXD+2nkVZ9X+pk2Mb7EOq2buzevI
BNE2gDSoi+k8XFNmmyW68uR8kB2L+ly/wJLAZVjGXFZbDjaeKmq7WXCZML66
LQQtfdytExVtS/wWsSpi0tSdaPNqzKUgR+RCKc6D0XcZQX6f58VfwKUvSe/F
5eOBzjYU1k6UhL9rhO5CIMBAZQIHP/TF65WP1anGlo1+Rmf96Lk7Hg1dys59
ETpiwbndBXUiKdn9j70odriH5EmAHU4G265ZpiyoM7YBh0blDiDpnLx5QXDs
W2fKjTrab6xDfid1ge4svbRRxaHtmvSY/VrK4tbnJAgojlCYKcz2w6llndW6
iC3JBxy8xAJuH7PR4TH4MOIuOvbVQ+O4KAg6EybR4chQJesZ+Bup3M1kQD2y
fxFZtIwVrQOPGC1UCMT6JWC+EEXmFoL2iM9A7aLUg63HPIoxNapbhiT7UwkR
wt3+6BMkTn6yR6HMAbRsWfgS0C1QXiJjPbYkgpq+iXqEK4KgMd18OYrKXFnC
Ne5fm6/qJXLWhO4sOwpTw2QRa+8nPDlscj11Nxv5sSWmVk2tSX50/bLDvqlm
L5DizY4Bzw8olTvzM9JH763gIZT5H42MyleJAk77XukMH+Ppw5xrDhuXLZXA
UeWoZR1iiYAtvfjS51t1n/Jz6dkd3PIZhtr6SFbHGxRYdQZdg4xZqab830jz
viqB8ptNy2drEcB4nmJSbS2I1aTFFIQsFAOTC8pJYmjOSEOu38t5QO0gq78J
oeCfkAo2IJUIWP+dzgaLNfDEAKkhGLZux0qMqCMiWlhTtG92L4wBOz8j7FpH
HN/X0yrEC6iIgNkhURk7iH71tHrUyZsS+STwu/DFZk5g7pu7lnzqQFGWVNHk
o3DnwILrThQfJn1ZfgqVlalayH6r+i272D5x0qSJJ+QzoSr0hk+d2hZI4Qbh
qxxRFauqwetXfyTiaHmTNpO+NbKp7f8jzsHpZu9MmhaHwe9HTMpLkTEdYMIQ
yOGj6lM0r2ytzK3nz0JaDcO59G5FHn5iipv3dzJ7VLRdWOkMV1jlT3MRLtTr
yN5610eRRVJu/YgWjeiPfjRRu9XmJM7bSGyI84+kPDxcFVThW1k6HeE8OZXy
JxwdQpEElMCzmDwrkzbStmxzOavCbo7NTpCqsk+FdazKaJ2njFaDTzO6+PM3
5Eco/q2LBz4qO0juIMNkVIG+pTuGbARIZpHA9toW8DYDGL4qLgHRH+Ggcd5i
8wLWmL2HkxHeBj7et1e3onHh0Z1SNbA5H93X56W22wotDCUKZw63bdi2TC/p
VC8AI2AV5SihrpO+ojDJ2cbzpFABGb70jKRS64RWDaSOLc3m2DOH0ZFOVakW
N9niiziXTemq+mQJKBKUMoMKKmkpyrnIylrBMY1KGjItYdJwPTPCjfh6rcHq
0IJ+uvPQtISk7KNHkNw2yi/Jd5YL29XXrHxvWGrkvvpEWWnZSplKTduIe3mQ
iqcuFzxbEUbWbsvjTG50T08rwu+eqBJatfRSgvHHdHecP3UzXVdNDr0uJxul
D46/gVKT7HKcHDywKJJ1K1GEu6de6JVWzTBRFEPeyrtWTqG9DLORaMWEZ3j4
1ar42oovkhZHs08BsoxM0OK9dZt8CPFDZVaymOKpClfyuWvVDtMEBPkAWfJF
ftIMPpgZLcJDKyuXVi0xj+Bp8KTVRdDJFpTeZz7pP9y6A1/OjGbsICrCD72p
JoZ4hoLdjHn6EFSz34wL77b+RmDYz/ZcoUHn7T7/46ckttza9j2ewggF6eBg
WrTOyTTcNR02tEGpTww9/1GKe3ovpkbWKZpzcx5+0VWAL+6XNRZpmPkeEGeT
SQiq7A+/JdSHqFFMzJRQtxbmIqsJmQItFdt6XJkG6BO+DCifXRTWLR0fhzkk
A0aKmYKRTigGexb2IECcSsT7nkADA6bNzLW/r8Li4DyknHxW7aAbA0TxC8Kd
3kjH9eI1ZcxRXK+scYyADHZc3UFw7RorixUdtDc/h9cMHEKmK28XnQTQ7R2Z
TGaFnqDPbnOdUZYiwXyejH7+Ye85MwEnlJ4m1pmKbibM6w1hrHDGaSe2rRp5
7VrMvwnixRpxlIlrYhV/4HD+JjP0tgrGpEhDidFFOnT7TV/zIxJMni6EJddF
m7LAmEwBrZ9/i2uUX5KKk+hNmiQy6PXyPwZ2IFltsTNM6JJAg97NgJERf5R0
Co5PB5ckf5wOI8CeCTnJmukmCBsGR0PLk8Ct4TF/y/gWhYvIA3HlA/vOkRKl
RwCNWu9y7TmCVefi7H1wmdOyY1/lkm85CFNIMTBYo7YpH5XI9WfGEKVKbTp9
scinRcLjvkLIC6jR6Neu7CUca3CNPGoIYRx8XrO/oVxNC709UV8xFVxfFS6T
vwWLlGRM0C8z94jzTAvdrHwzg3Bh0M4dKdZSRsWvmQs2PyVwYHonaEae0Xnd
zwD5H9CUbNBecq3lIn6CsMJeunY5QCqMapBlFX8m3IhLEFGX1mqt0uHCeacW
sOK4tQd73linAYhnF+oMYeG5B84OX+6HYUnEiJJPu3PpfBhCqMdMHhGvhi3O
q16qg7SXgqTiZqCPbbGw48/RVM+JuZg0NERXvuKn8g6rYBRqZ8bg9w3H/gAu
JHTR0b6zXB7nj9yB2Y9WggmN/gkBErkdNCbTGcX5B/fTkGZgkTAXnaZJL8ft
Ymvkt2soxZbdcc/s6Ro6b0Qtu4CGLxilo26MgPGpMF0SLGGH8MMlX282DNJQ
ZHlOSshT3lSilzouYzxVVaUz3sTgGlbB9V1vYBW3VMvjHe/T6xMsdxBP0Grr
ssoxJB+S33ENbk/+/mxY2YeBVYBvGwff7BgY5LyQbwA3x9qUgGOZTvUn1nnj
ap/TJO6i1Y3Rou51HfddigR2odBrVxFwvfLpDVXl3UfWw5uApiJxyFMi5Ubl
POjVpMFRsUDq0k8YJvOVqF+qk5AYgo7d1DN/SeeZEC0oBlxxVk3doTeOLEOA
YmlSKxt3sksGa/V/JRseC+V1t8kxMVCgkzPB9wseXIT6qoBSuiW9tKrnmo+W
nKmPqNhbCrntIXtlyrtILnMaM6vWcdwc7aQ8yX3fPDFwEVhyDSTlKyt7waYV
keFnYf/Vc3VfRHYOzUstUvxUqgxwoxuMnSJYqaHo9ptUJm1IbTUeyeGbSGLd
C9NQM1dSMmaPgKmmCzVXCuk6p++0vhzN7ilL134go7MPEmxyeOIhLOgXmxvd
5CDzTDJMk90fKiJIpWNI4dx+2FDTYZV7llfs9rGlu8hfqCo/uezLT+atuQB9
jTa7mTsHFQCzSrxOeOC4kajRc8rbTeTHUPl8rIuooeGVMVJKCVkNAVuXoRN2
hq8Ld9YLNKtK/tKx/2xE5mS2dpsDNVZHEHmDOjF56gmd/2UJBrK4Iz2Kw3iU
SEpFrCPDPBwrLfJ3JSvt0KDaw2H4kHew21JlyHSSV9A3NLYR6ZUofR2vL+fV
JxrWSwm+qne3FMM2TkNmFvxDw/SS9VUPSEiPBX7mK4uqau7jUdAIt94c0+D1
GOn3P6Uj74K2oo8Nb1hgFWRm5GpsCzMldD2soTNO6HySXhT6i2pnFshcb/+q
wPpA3z0xotlDVAdvWokJxnzw6hQyUoXBn38IXYUC6Nl84ZRt7RV7hib6A1xk
AL7td2GB5Tog1WxIAlLadJvdG1tHJRTaw5wutL1jt7rf+4Nj8CUAiuUpPo93
tPiqRpxcAgCH95NHt3gd8cr2cJ4aUnvrqa+L8Xk0Tm7ejHo4XsRfjZwosfb4
9XbHIP+teuxu1RCXTKC3vcdRSNsYJ3e+m3rPadpPf38foK0dZw6GBNVLqTKU
u47otEAYvPaas3DI3eimO8EypsKZC5yA7hsoM9G76mo2hTU8WMl6oGrr0NiH
OWxBOA3U13+H2t8ciKmhUwu2+SAZarHOzOD9Rv9bSXdUkHpylaU7+yWHZtfR
Ix4Vf8xwbDHLJ2f87bCAzCZsmAh9zAfrMsoB1HheGoZj/k6BwEkKgOUDd9lI
6s+Wy0EKmxa4yP2Kwio3HC+qRzo3zst4TdPdCl35SEWBfGq+8ZPV5g0jnFSc
dQgz2QOY861ZoJwiUwTmfJjGNSvvLGmLxFFKe6BMTza2kqoRkRGQFSQceMBZ
127AIxrwdOTA3KM26LzM6PYtmyZD+7jp7k6nePxqW6RbEd8h4KbFGgmA5mOc
qMFPwsCST6qAX3dlESbxoruznHjFM/aRC1RnhuWP3oO4qgMjNDpgCSo/WcWl
H1zesEZbyxgZspHZX9M6MMODxwTJNRVMqD+vCSfGaSvqv7FfMFQGFv70H7De
r2cRi4xawZ9v+EhYiIKpjpfY4+HvqvCLbrqueOsEiehKL/ASoZhyMdQOKZo+
QCXuZ9ewfgPP8tr+ItFX28DNdWWryI7bYTZsgaAuhJzzoyr5AeLdV0CR+yoD
7uqeZBcGUCE/W58PGdUFhil4fUv5UmQmLq0SIaa4sMjfvJhlDDZpSQC487Tf
hA/XWPzCgn3pWq25ViI9pXnAdqvkZHtUXYJFXzbquzNBrt7UcKPctrjmg+Nt
zdJNk09Gzwq8+5QoRheFMuPj0nw9/lBoriG5IKTDt4gyfhCcm+T6FGmWZatl
hkII6f3yAgi9Bkmqy+rFalZMpGlc016Xx1yQ+dZTn0gKlEnhMqCtwqkP3erN
EC34WC6k2BZtAJAUXfkI6suq0yBVLGdbbOjpPb0x42bRd/8r+wh24sh77QyG
dquC3gtdYiu7PyOsX8+pm96FXoFzd24AmeMDf793XPEjh1MIuanh4dLd6TcN
kuZJpnyKrcAwQRhlV3h+jHKDMzSnpNWNJ/MtT6Gtv1bPJX1Or1347skPVvUP
N34hp45t4e2vBJmj18t7IhFqbl6TpwsIb6GioqBAJo/oDU/NSGk0oh6lO+sj
DMD/BjfBU6e7uISnFDymwAtRmz2NwspXAsdBhz3/rbPMRX7zR8Fblclozp+R
ak79uJayBvRjHKa3V5X9iutgT6X7L5XSyrfhbPzVPROWVyX3BpmjmeHZjeCz
ns7zfsLSSHcYFNVPvmfiH3YbVTydBiqnj/MaEwrHeEDlOwjLoe+4GrbzEz89
tanKKscxvbJTaLe1lRCrmdMSbD9amoQSWwhRLjSGKJS6tR3yzkzcx8Xc6jRr
K79To2iphGwV5qou+NoK7DFgkRr6w9+E7eByjjWCp0pHaZml0IGbVoo3XsKx
DYQh7XGEqZW+AoIN/g4Eba+OS1ixEHmYS3H+/61gOb1zWmUFrXSnhcSoYqJQ
HvG1/k8Z6HTtiUPBE6QxYQ346AqObQAmNP2dS/74uIoVDPKu0Ksi9t3ZIsq3
DsgnHoCjZIZhKXPIxL1vxtRWSeOT13AzKpOLml1xcQjgB7JW1dicnVWQFaBM
jqV6CFPuy4bwFXHvK9R0y8pxaWV5a93h4AoKlRyvnXuV57tK9AlmVCH0a5cd
ZDzEKUWwQhOA2+knLzsVaSNqIE18uiBHb00+M0Gqlpwowh/jY4CwvcwRLLYY
RICXr8wYlvvgUz4ts7iPzOVIFqlluao3qVoEiwsVeO6Oyh272PPiXQMi+bGZ
jPf8PgHDT/PK8HLUOGvxYkvM/dCJeo7CvxIYkSSadRPf+uSbYmIcyOkktvJM
szXYURzhmY45dUp5HgDYodEfBD0WBHSRuKzTixsD2sOEt4BXBsX6qB5e3zpZ
FpZOh1saH2r9alVEZW17IvUKthric9vvPUmjdwZGFdHpCz11YGuYFnMpJj+M
1aFpnYt5IB+KNQRgSBHpp1o/pxCVdGcwKFDsayTcBUPgqZOZz1DIvKqWNu6E
KlbbssAFTjY7MhtMMwQ1v2PZlylryMyOq71UQ7CE6ETSzWPyoftRQqk1hNO3
GzgS9PfUybrt6j3KZpgxPpymCVL4XhN4YGDr/FsRghtEKtaF6RbMRXx1ji/g
iEFJNupjk4s51fyh0DkIsSBM+vOrhCiw/on3/nVo336NBKXvPplKgrWZlymH
PpSNd7QXlnZGFsaI0UEUwl6BZl7nTCHdEzYroxD+B+kzJrofzU87EHOjVw9+
EuYO3EJS5vtygYE+kwVr2xYI8JAYjnBydNk3zf4XbiLaNsN/S1wOQcjFaNjo
VAfOjB0JWPgmmB8HkvKR6TDpP10cXHt2IL9bCrcTyeIklkBIFYygbhIvOAn5
ZmxJjClmszUbjDCnGlAI2tJqKTPviPB8erVZxyB3arX1YCgF2YjhZjpara3g
J+ZaYRJChQ0V6mcuiH3xgLVLCrw4enLMKN9OHLzKYVlLNZcFO50shyG6E+eb
X4sSDF2ZUki2jD1qQXmniJPrB20v94WgX7z2Reza6Ps7765gZ33CiYIRRkuM
hlzEJkM8dBJuwlnAtjsPLWdG2DmDUpJvEMwOPXosAht1UqIjnfOdwsQ1L3pb
86i4vpIX1b3QQMvlHBELgFkkBO7Jh4Dxo8kDtdy4rZYHZEAT6VMBxRDm0lgm
AceFTn8JzejmCAfkzOb1RyHs4Bfe5LuCaX41Zu1Q1hgKk46fUOgA0Q6He6TJ
AICUU//OPdzYwRmO7Bw2eeO0qmu7fnSknQh4ah3HJVNeJkJol9VjaaZ9kgHc
BiMZojT0wfNza32ctFAUbLZcQq8yiTo5X5vy9eogGGpNZ5F2JLYE5kFK8CMw
C9D5CicR7Sj3Nn8yZhSAWyUyxJcNfTASF3G8P1YSinWPYfwjaWvm5Q4FHGhs
5igGNG4xoa5TJ+nhCrug/QwDh0ghs04f6/GZKf7zRLm0Ho0zfQm2s/z+w292
u1wQ8kKmRD1ThrnIHrZpwtqPa8LcRiYjJlZUylsfqH2OqxuAcIVtu4w6gy3D
PzftUFoV24nMMkmysU0QiXFiuHkaS76P1QaFzyraTSdyGJskbFVelVj19cpd
tR8mHgWSJF+JLh+7/KWGcYgTeZfH2Lwbq04akpZI/8i2g+SGBh0Vv7nCNPSJ
wEn/aLFEodOJ6VP4IThBNK3V4YgZ3VY0GIwHIIhLM5cuYC2zZQNnSqY0qJWV
VFlxC+NQNJVDse+YS666YWsITdurgqPaUWLAZc85e19PqVL/mjuYRp5+qnek
uh5Q+05YX3Pir7Deu4Bmqp2qv4QigiVHdn4KP1PfgWpJTsMEP1ie6kjxZYkD
KYcQbgu3RIYm7fQkqGvo+PCfUqKiWPrCOj7yUmpmhE1AUoRwDhJSSZc8iA/L
ga+zY6tPlkAIXruz/0a95WTLt43JAaXY7yrv0kNtJidV0RnHkJE3/Cmv14TN
+pM+iPcSKJqjWUuV0W+uAkjw2z1bl5UIAcSSjXpFqlV4QFNNV51U4/ZRC3uf
Yh8zdAjPtXtXDPHpi5MkyhFuHdyzOpnNaAqhUW0QOp1JfujgXdeDMzFrU4sI
fTXUkpL8F2OsCDre8Wn1eQIjZVT+x2tTObs/jyZ0etWcDlKkxX62gz20UtSV
fZzA+VUkzjlz26Ir3OTuRsFL9ddnQTBtm5+05czB0IsITJ0egt3O3WfKXkno
g81J4oDFWp87oJTaNmATrbVfrY7R3IuHb8Y/SYJJgjrZjhZyY9Usds/MPepf
/CWGqt96mhf/F4V13/OQqI/z9llm4mrFYmC97RepNN8bZHz5cFLyur52N+7F
ROXf0rIEQ6O6iA/jcpV9fF7HZo9T7rQZ4HWXRch4zwrj7zcCL9S3Xx1p01Tc
UteCwHhge2d30T+RwjxKo0GT1kJ87xtmMYg21RCLqzq97fE7qI6+GRufXRvh
0uo1MlT4kkLdt8KffCBj8e/2hdt966A/j4GRYW5QRkfxTxUL6e3vW0iBZFGv
mWO3pghvq1FZu8FYu7/YT5DAnpDN9VaxGFv2uHJ3vJYOmiYsb8rbaSUWCF36
EFW5RdFXUxhQZnZWl5WSI2QHtdY5v3EiafW3rYbM+SBYNBSqLldg8bCIyyxM
qpJB8J9fqq5vhyuijIZi/41oX0WdqLcse6S/EL/DmSziNuPUh2t0pNbEzthT
RzClYflXv/Pqxfsj9YSxu/z6ylk8TTPLOv5swMSjW8JDDT8/V86PyRadhLmP
bTU7XfWIV7+ivdBJYuOBzIw6IchwIR6ocDOw6RkyYDw4LO7iTYqTLMM59F2n
kM+eX3BEnfePA0k9l4rof9obQ7+pGxOFNfdawMaBmQ+71ShgadKnROnfvu6C
p4C1xBcFThd2a/VQJonwioNIYdtIddqa1L7leZzU6VVqeytnYKOjWQnq7+Cq
FCTt1tkYbUXWLdIebxJEXcwE7cpki0eZUBr51qr0CyFpvZDXPlntYgSg99OI
IO0WhapEFpJBTzU0j9NUkK/VffZKkxghwFzJ5PH5bFuVBufqbd/fSvoCLhZC
7hQKMlGpeToyTTXW8PoJNn9GKwcKbYtezEs8Lrt6Ro+LJ3UF6Bg8UWT9xjzQ
/GfVgXHbIOyN38JRkCMOUypJJP3bN3Ty3+EnASDj31OUUv8vtFyRbiaBhmnI
kf4uwZtGTs6fnl1YvPz2BA4SKW9Tu2bm0A+xl/fyV8TzTaf/fl8Xp/FK9pP8
WDD061ogUcJ2QoiI7+hPnXaFJqqrhVrcuhSIMkir3Vp+Jk/mcS+972xGK8c6
1vrWKscf7dxd428XuyNJQGQws49TzUXbjJ7ACMLKeXYO01Qu52tET0ZVYqIv
FZM9jLnOXlO8f8hQhdEJymnUENas4OpxOhXyw0jfHz1jE99c6ZEozfDWuRaz
eff5XkJrYR/j+GSr1ue5PVKf6W2hpVyAC3QsLA91F5U9Avejh+bv8tlGg3uR
l0ORpokU040dTPbi0NJ4SbP/aIO5EyG0kjavWb/D8xparQ5App4jhGNtGHQ5
wHmE6y/RbFa1qZhVHTMgZMRS/oRjWyEObifJkI7l7a/udBzVa1OrTQfao2Io
Qp3pv1hIHlqEEaFj4nwlaLxff9sVuVv1Thb23XajP4OczVyohQFnab4DK5Jg
QF9/8xU/4wGRwkW4Fm8e2l9wXc70OVTTxSAGO4+mkVnsQuc4aLAQKkzRkBOl
AXpp3j3eXUPDKZHT/2UyI5F28aWF15IyBRAtwACI/lFix6Nj5Cq64AGBxGYQ
LmsctFg8IOvN3I9p9RJ8iGJ4Rh31r4XHjWjE3jgL/iZqhPfdGoqoSJOzlOjD
D5KjsGgGMX+j2Ayf35xCq83G2BfEXPJeTx0vT/ZaTomfkvIdaS9RThJiDYgF
KQo9QMN3y54Q3A+NygUFrrqvjNZwkymYZmgMEd6IAPbLnwhOUN9BP+8cQRYE
asxBdzjRcPBXLV892DLlqnHVTEQeiUnD9DjS1av2mm7nobrdrObUA1eY4Kqu
cGmgoRkFvDHc20Hhg/TOxJ1bWx5qhd19rtORFkZ0mSIjYwThBT6NwY8DU7dd
AfV/oqsJrhGrW8BdT/OIeYEsWTpOtcx5ww9dTDlpjSOHmjj5zRJ18qBEFPID
3Kgkz915MiSoQe3jAZFZrhbaJzcClDIJaaTEnb2tVs4buO4vJzY7+RQfdHWJ
r6Mbq6RucGOyvUI3+svpieeLkieSXDU7Vhfl/edeN3zsGBsyvdOkNLVQzAIs
ceQbZroX3/hwmS2Pi9qBkIRi+LQS22PT8pOSX1iN5rw4dKv5aVVWfOridnmI
y8ZErrkHRFbVuzZE4WEew3w+taK5fktmpaRX27/ba1VU7YkVavjVv8UpE1HY
aRuDotdE34pmw+IGfJfaqjEQishMPYSM46r2p1bwZOOs/rjxYk+ZjTOj/JFi
3upuiv7ouxv5VFeB1UQsmYFSpE8qBXmEO1PmLbMqBPXFEB7C2hiehc0Ie5ge
qLXKPXl+oGetgAQR3RQg/rHzzjCwWdWPZl+ZbzziLDC6pc8UWVQEymHeoe8v
zRxEUjn3QFNrvREJSI0HiZDqKbcYnsSO+giyFVsIAl95j/TINZhw8lNcf9Zt
+CN/vIlyUXu2EzMRpFEtC+88jwUtV3rDhmkLu6M+CG6goNnboiLEzY5JqeEK
yA2dz8gAMqv8QELr5mC/ddOCiNFxWAJz1MR6Ot9RClS9gUVuKxiM3bLTWiLA
CTEf4LfA2866QtNd4EBSCS8Fme/vh/gLaVsE8jGCDRjSJ89UvKj84XIoFpay
LmeUJQemuF2gIHrMvJzWgoxdO4vjUChOyzDJ+eHyIAMxCtxM0z1MOEvCjtNz
7owCLMD/HW+Z0XvuTjOt1LGuysBD1HXk2AGUZkAYApPrB1FQohUxRK/+vTrC
vHcWRZlq0MNtDnj3JIyl5dYOr8QloH3h9Qd09O5zdMe7JLFrNyp1L7Qq1dpL
wUx2wBwYO/b8iRfB5UUxnDK/h6EmKMUjMYM5N9jrAyqG2Wainkekyr1866vp
auymbmvDA+wpNVQNYUQjOE0ZtMoHaimR6OZ20tlUucCRHJ6c/tAUWsp1CoYR
x+FaamAioZ33tUvO6blNagmFPLnVHChLiKQ2Gmy4Y3Ocfm1tXx3ROSUB3kw0
OJhBMORDJCGvdcwTwS60mVAzqLXuVGR5iT7AVvxhqrRrasTA2GBCW47d9lKZ
6aq7vId4z3LjMkcmc/LWUPi1DKMCMQ1SDHOs5Ct/sZREFXtcLTKPyDg9egam
1LtWbw4kRNTI9FjGvoUUmVMG0lpX09t8JWI3A1WQN9hDy+bU5PI5R/lNNzpA
ysH/5owZaQzsVPafSqt0sQ5EWRwHbVjSqWeCB7bnmw/LHuyKqjHgIDX78p2+
7Y4mGExs8yDG+01bmMAW9/Wv2mWTjJiCgOahoHyaxgFueYEYJI82XrpQQjOo
3nRy3VEiqZSUuuWVWF7cTe3x0OiZS3gom/e57jUy0LNdtdc/s6yCAWCDORzv
dZSEjE3Matq7oNIbSKUGGh5Q5Z45bbpHi0C1BFarhTeA4jqM8P/vsBXsfHR3
gCaJ37H21HNS62YNDnupHDO1FptqzE2OTSH1wA/U3iiMEGtgV5lwSWmD1YcR
EvitDte6aTWGBZhWU2uupGXO5ufAPKZ/uzVeustaManlEiGwThTsAMO0yZDW
6gCYY2CFFx2DI5bkf/bgRrm1pJbBppKwFq+V08G290lyJHhv6AWtv4bm89nA
kF+mHjexdm3P+GPXAAS/9/BqUSP1F2a3GOsScJQNLehqCzbg1H5Vwh5v1TRz
atf4WMk2PkSD6pX1a1K4r7uqJufYjrcTFu60JNjG1iuiiaQRXWDvB1HDfc86
DrFF1f6Se4WqEqLNBGS+XvVvt2jR7oKEdwa4iM1Ish6jsrb1uX0NRowfwCSy
w1bo13OVKwlOttAYhWr5v2htJIwrWYFBVt3bsCkWi/w92z2PojZEnsFia0t4
lDDSMi90Dy1SRcY7upfF0y6mzeI1JrzXL8/bJ/c07GziiGMmyju7I3/CVmsG
kfGsfr/zeSffTnDYqZKgHOT86SMwdRl4IjatOLAqPEyy0JdzeUeFANkYzDOF
RBBZaj4A/8ruRyN6h10BGcPklB8krqX44m81UdZH8ETpDKh51jxAOYpahLVf
64ZexlawZ11hvSDaPyMPhcUhHJMY6PwJ1tFDhuGjiiuIz26egMITvpz99VyS
viP9CfOKfzxHmMWeoEy2qZMBI+fmlgIkd5kQA+7EsJUSNmRXORGUbAGRMcpf
Dy1gDRAQIfWuGm0E1oUz7qFEO24YEHoQCdzWqWi7xPGQzUS5k2QJ1dml3RY6
EBrQAE36XaOsDYk5VDtUo6Jp9883cfVUGB/2puB9f21gdqHXIPgtWPQYx8yC
rHrWK2AtnUafeOgqKb9tmfeH9KKH1DEa8gj48ymqfe7ccjlVgUPPa8tMKsQF
t1XzAWBWRbzE9bIp8o0Xnqr6zU0pnn/HHDUgy7bNwnAlcZN3etySj6MtFhc7
vaa+tD/NyR3pRYr1HXthymRnkbrZC7b7CDKke6FNe5MCTWOlYbSyr2ss4l+B
gTFjoOHMaEh1CjMEqRn1n4VY0WYX1xhSmZl3Qw42DDcRGODstdBHkqXXgccl
xz8z5Bo/QP3nd9Ahligwkg6uQOLo+jh8R6nllOh/9AR7EoXpYpaC7XclrzWe
QOP9IlNuKB49P3DqKc8TH+mhS3wYwg4stYdEOTSQANV2ztXY12twnb1IwO/O
HKT5Fr9iYoGg84RSxtqBAo5q9K6aA8TFFfvrkZkaLpJdh16qpd/TZhhLCPGI
PocwqxBXDy1ktpp2QBT1JT2+gb2SydADYxzWHXzPbJC1ZIVoo/S9VbIFWh2z
eI5FNkgIQYjRMbimz7ZKtqdBukAfyTam4AeswhFlsiMh+5Ke5q9M0p861IZY
gfPDucF/EISqHxaaArZ5wIPuKm7zxC1oMzuR0wmC9TUJ8AaosRhJanvlA5rF
v59WADRsX5dvelJ+TMTHALkf3IaeMYdhXqom7C+fgtL/M1mjkiIJbzTYqh5g
7Tin1NekB3Uahy320LD2+CXxl5MJM+JUFF6hVx8yPvQVWTUFDf7btt26v0SU
lptDPBmHu7rT5LV3jxukCwnUPntEUnI7/7DO8/mR0J4spzVGyTUARNbdsKlZ
XMN3T3pFSdwmhku7kLvYTyBrU9i46fU5G2dlSsPXe6NLqt4789DRhPFuO//m
CbJwXCT9A8bH3gyogz8AE8PNhwp/OSr/E/hKFdPE8Bb9/8TcMczVItcUWcBU
wxdnoLJMd+R/2fl5tlxz2yAz4OQkHRZqjpfKwNPsHSy/GoqilBWeBY+fxmwx
uKSiL8v7n+51vsC3Pcr9GpCGu9kOinDxYFBoHYcjHGVPRFJ5OUIJMBk8yQbr
EozoKwV+yQthdyztam0If8RjbL1mCluqUwlq9vm9ZkDd5cMl/R82daL0RFBy
7s7nljmyuWpgWD7rhbtduM8+py9QPnWVvveQbcAN0DSm8T25GubwjwENdGdb
XkRqv6JjCbWGs2tFtoYw+HGEOZlmsK052mhpSc8Lmx5gI1aWEf9d7xXqjZdR
leN+jFCDNc0uGz+qcIWTBCv2/47VUBx73VjNRDF7nFXhy4kHGW+3J1MlWRmm
Mf3SVwNL7u2+LCKNUgrqvej51SHPpXK7urpJw9CsttOlKKz3CFz+NNCyldSs
Fv1dRcTZzCmnL1SKTXEJKJ6FepqCPM+pC+nhsC0WQAbRsWbkm/8EwvbX0VrN
FheqzXTLBINrWp35PlyTGHUqEGY8LrONxkwSxQqAEKf04YAVkVF5yT1JetzD
va+/SIJPhhAfN5DGJDR0BU68rYadGKujikGjJma2NyfstT9hjPEpr0tIZex5
rzDBBI8qKGb8aRNaPH8s8BJsWZORIPosToxr5zHa/hKrQSMXWtBw/TtGET/3
X3wuAT9e5KNrPA/943s2yTOCUqQ4Pvxnjdf5vQZj6sjOHycFCXwExf0SLg9q
3IlywWNTsPYBsVjALM9ux2bki67ZuJ/V9t/VOMJpbEx9N5KMqHB5bTl6dv9d
/Sm+Zm+w9r0vV1TlIIhEOxrOXgoejKrlnOiCkFxeVxQw/pd86yAa5spdF05z
cM11alXhUSmEufzX12L2c4pvi4r6IVzbpeQTI6ywWN/3EUTDAL1u8P9wEFZX
QaGXrK5BgUJY3V/L/dlrX6wHZvxSk25vzYs7n5hq6cnWAvXuK+aZVGXoVbWw
uXXOrtlv9yymoc6wDyd2D5wzkkgdixxw/wv/OOx/t0GsG+3FaH9QQTnkAyi7
VhCtZE8xUA4XMRVQ0trLch7dMNizQYWfNLKTnDPmvpijpaCmcEkmtRzy1fDq
tL1ckrlrqFBRCXla3nPs2tIJ8zCIMH5KyKvFswvjwtCfM0c/VO6Wi59Ng0ef
GQihezxhGF4Zj+OOPNOn7/NAIlgkZU6cuvdjpTGqsy2wpHmb1rJgafuSinoq
q7dMplnbypAc8rBNT4qjH18KTnkdPnzC228ClGO5giTYv8EEOJvUTNdEFdMM
XF2tu44eEmw1ZzJ3S6HnfmrfIgo+iyHo8SP2DG+wMjgYgbLtWQAF94gIciu9
3CMjuX5Cy/yzF838MT+6zKLh7/nMSV9QfacvispNs+n/PKTuUoSQImQIZrdJ
l68UMrCQIokbYepg9LLI33lT0L9yDjl66oB94e9d+VDkWSx2vmKRl3wZ5L7c
R3eJFWSKOChCxdLU5gCnpQuNDJJajC9OGjCUoCClXz/v7NJEUxWM8N6DIf76
r8AjUhN3owhrynRglO7pMb3UozbupOXe/pGXfrnnlx1h47ntrLjUEIYjtJgI
bJ4DSB0YHCXLFPsXeUbDOIevQburUYzMy4qhSTm4FbdK+Bj3LxdXd0pWuNNX
yxILGYHFJNZc/IE6AKJc/vX9SfW4BgbTkSMMnNTAaRUTGZRm9OXX9vX49r9I
ikvE94Rw5jAviMskKCRv6tuQVViyUiMEK5NFUzfB7TjiKrz0YglcXpOMtuU4
inP3t94NIxAzvGMydDePvnlT31CiPlNmymWSCU6+8Tnxb/qrDEBdndTsuaIb
aOEQqwlJjGJniqTyWREkQIV+3Gq0qmoOnL5sreUHtVyjAti3wo84TiNfJAiK
svMIPfkcDvCXbFdXc/I+G/xE9qAvhssrSNugBGKjcY37goKAKH54z9ckqr12
mtErRXE8U7TSN4wuJvycqcupRYfSzyrTWX+sMRLE3N7ZtoHVl4BwmZkasiL+
bBPFvL8B4Q0+z7XDIdXh6PibpPLKRPsZUQpL43r2TBz6DWL8JJhx+c+GhnmF
b+YN+V2SgrTiNKCSRWX4hs8NssnqneYEx3A2MEcUEk9huEy68nnq3L3kL9aV
OgukC4tBbfzMXF9Tjw7YMdCnC+U3cULnnyTcVEVVc7wdp6x4eOjnWs38UpHp
5/8w3MXnEmw6MxxDN/heKtlxSSqxPm/a4v3wmHjIMEcWOtiGhKsiC6GDi7oD
S6WQVeakqQuPC8yBjD2THRLxglTKw+Zmuo0moqJz+cdhGM+oLF32J2zBEPpb
ya+On4E5zTuoPKFHgh97pl0l6FesX2aNhiqLwrSyyCUNOxXLrY67sy1Usa/v
lrNCfxafTLybj7HHug4H5VJB0XhzU1ROcBruml/Lv93iylXKUAVcxRdykD4H
duiHVJ5Q3b/GRn32P9fd2oxFMlk5VGXfkOnF369CettfTr5GBs3kBsuo484c
95ejBRPXfPhw3A88MWkVd3CmCZ7UQe+bzejhixFaJp4Gz5kwDMCQjXAIAN0u
l6m4t6QaKSOjB4ABZjnkW0lzmzvM1tSMVocjIyNl9YjwCkeNhgnCdAAkIMqE
qkQDoGGXhkkpPVBttDPcd1phMu7dhkWmngBZLItugfGge1b6CHMekyoETnnI
iUsQ+8UsLZmck+o3eqRzr1QLRNvss+DcTqENkit4dOGx4IQAc6PirzHYaVx6
Fn7SOJp7ovYP/46JbgxFXuoQL6ijmX08fQJtgHA1HYNKHkiqaVikAih92HIX
LH0aLSdf3FbWoE1EmUQzY7bwtkjkna8etXgf4rXLK5ty6TR5IADK7Ajejxy9
oD5bM6Zm7IzS/0EggOrlKQ5RHrgLoBTLcCAuDF1yT0pUF5cWqrPzsBmKsIE2
MTItKtP+kHsr4z++xUY2Zy700pE1lOcK/hOAlNSwWvbikBBSTjpOP24YtF2P
TlmAjJiwTpSDuP8lLfbol/DjB5fih0VtZ+W7An0uEum4Iw0nmHcyVW66phKw
4kG2RJX4e3vaeFtAUOiAgay0KWq/nOjewYAIbLVU0wkcBB3STg17tNvXrcFp
I6tYsJzo4k+SkkQFvTdjNA4G2A3BzPaKqyQ99EHwy5nNgbOUzIejFmD/eoQa
+BzSjOns33Q/8/SVbnM/b/Um2qCf6RF5jjmXzL5tLY+MY+L5X8nZiUuAYnaJ
oPEDLejaoCTuMzkpV4nsS8Ybp6YEyzZkiipAETKi2JI3YWYL/cKFe75bOpOD
6OAm0ssqX/KImqONF+b0ysOQC7Kr9mQs4QtcN56yWMVHLvNc3AAJkeK77sn4
cDXqaV+QQiLOkWHPwqQUQ6Ki5fn5dAo+yNA3NhaWniz+QiQV3j5V9rWSEiZ/
1cQWrK+f0/k5NgnWRjTK8pH6l5nmtvG3zFt0nkmckR0cR0b8yR1MWYe+go8Y
dhxq0407xvg/F8mBAi/0BS5G8xbKwwJ8zzyeON+a2lGOJrJ6Jji3RyEqj67c
GjXlvILx0Mmy8W/tthi9SIEN7GQ4DfXkhQBqxWu1NtAzlg2irAZFirqJ91wj
LSS99M6WgLPTbVcOD7UUAdAgeVDwCBgjo5DOFMu+wo7I94vRsKQEAe2eCt8V
f7IiIX1tB8rz8QfEUKICAX/2oNn3lr/qgj/BMzrIN3fpzCRKWatjtXswrXos
qeJ2nq01t8c29iZGFalkqKKH4TrHotdcbRo3Z6I0tRyOIeKhBvWZ1ZeWQRi3
2S6b82Ezj5PW7f6IRGjTJzyzWOTNX/jiQaSBGGjIfq7JKnUb/a96MnfXvdD3
fnzrzBpGKeSnfbyuf+2dEclh/UIgFCrmQu4MG7Y9MZ4/EV4mWni06kNuNaHp
PYrOB7NUAYznC7YaNxeP3+jt2oR/DhXLTy+HE58iWXkbIqGa1gR3yS1y70kl
fwloJVofSfaxboN+Zxc/nb/Or3WiEJwsmpvKuggkzeIEUeo6VXsYqdN6VzNK
Xa1UdZ3OqwZrEk5wFhMlUwfJE6EufTd4NNahBG0j7+tRaslWXkaT/H7b6+Ac
eVgLQ9LGPBWQUdx5q5yvQR71h++5lkJ+bVpMka7eDRtpdkGKYaTIqot63sMG
7+CqstP8AJl1DwO3NXg+pTJwHjx/DTD/wPkKBpO7eccJo44NtjAQnF1mte01
RuCWzy3v3WTwZAk8m+1tcAaB5oGgQvUt7H1IIaIgbwlRThsUG5WR0P2TzXH1
tNtMpdiM6QIfXhSmuYq7b/Rlur4d4nOf4vpUkeroHDPrR7MhSoKNK6li/ev2
0n+30o/9jsZQtvGFk/ILHEt/xOFJpSWcf1n4wIUI3jOAXaRLYnuA0HBg20Kh
wiPivtazSO4KL7MRUxQuwOhnlTvJKfVTbAjchrQ3LMnWoYI21qoVVAx4eEYS
hmXRvKWrWquSv+D74aWhllQLAm0GtSc5zk7DFW+xLAG4X5RL0hCIk2w8QX6Q
DdkamwdreMABOm7ZMKk5YdjdoikT1aV4h5QwYILQjh+swwa5koG66jSq7bOn
ys7hy4inFMQ6duyHaY+daB5Hyh8MNRMS8zhN+g++hms8oBGypTbmQJ+BjLQd
hbn4XYV9RrVLYQTmZopozkhLnZAZ4DZzarjqEvYs/TXZfFJoo2ycAoSikwUu
3xLQl5zVX+pVeXOzi11/D4/2CfpyGY36fUSheeUrmbsQoThcYn2Xp4v8PvtL
5etIFmHYaD2c8Vkrx3WAcNZZk80cklUlrtF5z0mh0lAR7H2YwLZN9dG9JzMC
l8lJHyg637LPf0Xgv9BioXS/1QSrSYn8vhqHe8RZxguzi1Mux5S5Io5IA3jg
489SPqSy6exZi0oTe+4Ud7aU/1OTUrHkR+Xya6hiNN3N0GZtAptb/fyZawU8
rg3evQP+zTGbYaZEVqnv0thN/AHFYr7JEWL+ZYrjZdgvsqSN959bQl77rWpP
v9cf6o05Q4KgvEZ6LklkVECeaD/onyRdUuB3igpdYZles9x24Kp0agHN9bpa
oqeuSIDZJ9z8rFPJ7WWhxuCRcr1AKkcabiwfcsGzvYBXgbQ9clb/YuTg3rZm
sOOwnbEgqPrpwGEUubEDbJPJxiCHZeEwyAue2JHz6Fvy8UWHslxf3uZQmYNs
G1WajW7wPylvS6L+llkVnJbtQSY56MAT1mM6ePu8DhZrcQLOHi8B0+BIsgF7
gE9ul7o6olQLFKXpJZBqf+JpncqylIl9NDDWgHsUM5uVEDc/DJuAai5NlFrx
nfpNvNLU6mqT2T69qgHH4m4qkJ75zE38OV1LosHY0MRR3UZU8crExLSdnS1u
UHK9LQAybOtBaosqLo4WYTu2BiZ+6YPPCSWzIP0/FSBRDryxKOyfkHn59E4+
TtTErOuYIF62pgU68ysASiFcRB2xRHD5jcnS1BedPzlGB+19KRdQ3L3g8CS/
zjjCUft43ubKHy3sTsjQ7yydu9oBUngiSziKVUngFrLyZlnDkKYT/qRLqxsN
P6TB6OVblnsBoWTZ7FAVfCYpnuIUsV7Y8IHpcWDwCm7QUmhiKG0ktMYfVHdg
mwSnZ0lLRUmqR72yXtBxjuMBhMcIREQN9otC5+cZ9yEcro7/Ff8n3IeU8kUE
d0ygVWL3j+FR2OTh1obKJD9UW3uG0SDQjwaCcatM6CG/ImfEcYCzCQgpfqth
n2NJXue94bU2Roz/zM29iURj5wmVm0h9nJOeKkDxw91BK9CEMmjgD1D6gy0I
DHzm29tYaNCWM9VClIfoxi518UhiVW1AB8ZwH9AxZLmNcvsRd0wBVJbP5Z1d
wi8CT5xx6IEdeCbp7LoewOnQRZQhHKT1ktNNBUFaY4tqxWqY3+SCqkMtKAZm
NuO0oZmc3bBSNqGqWOwe7UdFb/hC7oler/xuyxIGEjpdL9QtREFqEjC3/HWY
brEjmjPl+44GrVJMihhbP3AjObo7rZxVQbWk3THefsyb1TElNpSDOSfwOAVv
ANDO2SFFgujFPAdZy9VUQHxcQKWQ6d2B1nUnhKEkOfLA20v+jmYklZzv5ar3
lk0gMPJa7x5yJdc1UNbimAu2Is+h+tIyH6NPN8r6ikcsT7Py6cd4ZX+cx1es
wCl/lj8jQW75rCrrQyAIrbpClAzblkUmFbP5StOsLLaCftBnTL1buIZV18Tp
2PI1Ekd35yRLmITUK//D0LyVYSE1eABVWJAdsq1TQt2SRZtYsGjx7rgbn7vD
3mud7S10TRcIg/J9edbiNNUrnh00sO9pYFN7p9QfhXEmoNdCSgtjFKlYn873
1npmbFQtdX/FlIp67kCzgxorAZUfJFFp7618oFxdMPrVmzCATZphmsfaMVnZ
G02tICgAzuxiwz0R9zWYAN5AF7toVGSmJKpZq4VM/Lf/l2SlDadO9+zj6k/K
hrFSlD9aLzbb5xBullI3IvTAEO9ClNf3ns172VVlJikEI0K1blSoCq4i1pHt
t5GKtZotCwFdvy/P5x84X1wSy46FGjhlcx0M/fH4SQoBrQ3K9NZ7Z9XVbOIX
8xu3Mqr2/+uukqjeVfC/Fl+4R83NU0ChrLCvVq0NjJqAv+lTUZjgVRjrMU2G
2wrNl45Uwd8QFYleV0sLoOvCpTi2vTZ67JrrjfaQwH6uVrKXFf3wXnN1uc3x
R2Vm7jWtP1ESNghSnTPY7CtgswBfTMcuMKa8NIaZzxQGLK/mywag944uw1kc
rClGFsPRELutPTsIJyEXgKrkebQvVQXvUy8+6GHFIEIbYXpQ0YCmhNXEikC/
XDMoMKCmkyjN53w4ODjTY6aSf/XyuNonKpnx7zs7D2Kq2tF1At/+loJsRIcB
bHWoQERurVoPjmZXG6R2+hY+0HwFABS95XlIAGdZMkQlapppedQlXa7DYO6g
MDz7hfKaxPuhMDws8ahrkJwM9H9eV65ZBAnM313caXfu/S6oL8Fs0UV0X5rb
Z7a8fxryV5H/qM/Ty4oOWXGUuPZv7gWOYjTB20smCDF9IwYpaBg1ZQPJwh87
fidyH9d/eDIWvV3+XCBEN3pCLU0XRlLM/pNRGMd2qIgTBVcLMqwLi2RuLa5E
ve7G9NBJuVeLCtbfoQLtRU4Rew4b0D9i5Egk+b0Da7rP5f8aR4sT59zCaNZs
pXJdWJM5RxJOesi3sdRH6/CT5q2TepsTEDBNit9yks1y8fpusmopciSG6sxq
T+a2a1nWck1LvkD+GG+jboUcwRfuKvbgA3vKECDj/mlkLaQUf3g8h1wyo25a
gBenVVX6Jx0HtVOQV6wt7mzunFcwatATeJanBlcg6v2MADVbOaiZLTAScA4Y
9/V5B+E9nqyPFe1pWXIqYByCDXrhaD3+2kp+Yyg1UhdIDcTGEYbos1VKJtfF
wucGBu1hGIfhTu96CeLn4/u5tqe3XFb6qUJE9qiVT0qyQ0qwHPcVdxHk4kF4
vS+bNHLuWNFSdN8E1JeGCE68dP11KVBSWW2Ceg/YEIr7T3zqG1uFXNeb4w3I
kS9HkmLIS0LaInClgo5GnYDTsx4b3+2T55LAjlLsFQISCg9tQVgJy1mRsELw
eYTSYVieNij001HlULfdanvNUZbNdyg/Fxxu04bJT/XMNx0rB7a14nlew9uK
kMDT0q5+RiTjn5Jvkgug40+MLHwB84MP4n/H9NwpmbNejyqx8iNXkapcGLuU
arxyqUNE58Y87y4mxinkdC8YSkw7ugpjBLs17bUsSpTp0t6xKI3vhKg+YnGP
kHgFLdGU4YExo7hWTgHxZaeb8/TIiv/wX8qZwl+brtIRiqzfmA1eyEoorMmc
G2NYKog9GisIjAcviW+rLaDnguqsZfoqQ+2MGnancMbf2fl21ggE8sbu/nDI
qteO2lIclhYa6kmGsscftWcv/nqe2sgxDKXvblWC519ecSajMUsNRq+VbYQi
CaTj1CnMl4wtsET+RgVD+kyMKT9ceI3fvvn+5iq0mZ18epsDxoG5LNc39Dpj
83jjUUjNt/XibIVBoEH2RQVjPdVDDU1AQG8MyLep82VqHuj7UIB1LW8JWJo7
56mtFwhZ8Roavbl4/LyHFFpn1G5poTiBY6U3e3LGdbdQaMQ/QJ7vip3sDXsm
vhGJxB9slKlR52phWNB4iYd59QwQsKI3pAAq2ji6LdmuVLsbH+CxfK0GjHI4
AsrP7ZNv5JM9FKeOi+/sxXbEFld8AqQmP8KykVabESoiKGw0+gXN/WGELOg3
xAJWd8YVcrO38RsbSfXGHOmcxImDlWoRyOJFkwXGnzD20ZyBf+U1IxMSytlz
BgtzSONXpA4R9kMVi4V+L+2uybXOn06ZuNg0ilOqS3USJc24N8l2qlVjz4MK
X7X2gRv7SY93cHG4D2iHudnUlvOKaUVSUs3U7HX6ZwmM++Q3CdHBxG+aDOWG
nT7A7xdfHmjuivOCEzeMVYWukNkm8qXTCAe2B6JMXfUineCyQN5qdxTKWRZs
sqOLb0N7kiG0BOR9ny9PwpVkDeShzIOt6VX7yEUp590abZPSELaE9YCqWerQ
JDRHt7/+ef+V3neY6/eBgqCzwAZDpoy/kDjqbGsjKPtq2KwfBLEV1UMxagaw
ygJ89ri9jrZNG2dGNr22VdDNCTv80Yt6Ct5htrUR+v7z+CQWUKkXnkwnovv4
ApQbcoGEKCHDu+rAhfCOCFYzhIvUqXAB0UpFVb6WYEYo8KEGTr7M7eedP1eH
O/jY+de3iZnb7EEhndo5zVNUmuf4m5aZDr0FJvgaLu6mTjeWCMcwEUMZ90cv
hqf3q08hRU9hVRZIGnUF5zy3/JiLatlO6TU5sVB99KoW5O6uJAtePGIcnJ3p
Scvkxza4uTZp6E+RwZ9ObnETZ7zcbcCiwV70fVeaegwJUyAdY953crH4u0g3
bGUMrqYSyNMzn7BIsqjovkEnV2kpnwk+Gz9hU3+I+q3aPXvqoqJ/n22Jy1zl
fWOUe2O9AT/+X+tDCtUNS+WwoO7pRxIvz9GHPxUGXhyDCrLqh5Z6rTSgqJAm
hQ9wWSm5iEdwmurM5O1CldcMEvUxpJZfSfPOuJstHoFPIRXY4OcU9yZ8hctV
t9FYBQdQ0qo1o/af1ueT7U0s7loF4SSRubetQfyFmVm/nbr3OJiOV68stgux
7FOWhGxrNhDbIXSSV9f1PSuCrtvs5Bt2wABODLI9ZXVZvnTdI2YsZEcXQKg3
3SoME5A2R3yyLnHuIxABOPqLMc2of9XaYqrar6X7wyOeFOL0oENwVS2o1fu5
XqI41CKwSuo+SES6Cibcq72SioDsNbmxtxjvMme4PdXRj49MtU1odnAEgI5R
nvw8gfdfLrJ+Bn4yEytfWaNB9pHYHnqJ1KmT7QgYO/3WW+9mIseVJn6frnUg
vRYI9hS5+BrqIAANn0dQczDsCn2Ir+dBHrYh0IPsAKx5gfPu2doGOCemDMHy
u/ldB5axigkiKaeP3Av9FSgPAjPkRGmRqLvRsNogiZOq8cvQndzrqmMGEyFw
42LIyM+D7lGQuhMiPkaXWIYdk7ogPsyQyIeD2K+7hYnLVn5/VOTHNdh7xjek
W6NqkNY5JPZqU2McetgnygsS36XXm+RW7W2mVJKNfuikZznOeuv53Ac1KDr5
IqyuOwmCywdqKs27CDWSVx4oJ7M2bOkJBll5e5WYpPJpRD3fvt5uAUnnAA5C
NEb9rPntsZUI82SRznrIIYrlMZ3iMtFl9cbnnaaLIpit0anicc7XUBT78zwd
UPv5iFk30/xwlVCD8p/aDOouOmrQlfzOHXbbAciw0gkUBqApYSjHU2+TVBGH
zo87oXPcw8QRjP/FTBRJnitbw7HJ4+mHixwcN8zac/9tIR5AZ58DryK4VgIA
idiQ2YXrwS0VKQD7LYd/t6XsGg7rUiZN+qZ6oTg5aZ2BOlHs4L+ASRcb2lhJ
MBcb/yiXQQcODsKEdVY7YMRoPJ3vC2lkKt06fSZUS/2Es6QP1ecKdLNH4vfz
dQW4madw/kIKkxXHY8jn15GYBn+0CiE+0VHMQrvND5v2OMISiJA1QqcS2KCa
bcq0/Yaka1ls2MmCfJANaNL4a0FvPCxKyMYPo2eeUcji+LeUfWzEBXS7oy9+
XfwXYUd23pEbWf5fryacxfHUttCeso+8xeBM5PF1Mycg7Ea9CoRDI4bwJDgO
UlgrIIt6PaLO3QKi4VutJwMo1/Ka6y2B3xnEFU2q5jII2ZQV4PiG4NGYRnK6
omg04XqB7edRvthOQlWHsXOMXqCXkn5Xsl8dvP+QSm0QtH9iMq41WTP5QN+5
riurxQxDmxIgYtrYFlpLxTCpFF/3PFFim2mGPkj6MsoE0dwwFqDxj2mQ9IxC
hdgdB8gSHcFJJLD86QtzZIw+Rpmn1KqQW2zintYR1AwD2p+GRQEAwh0osZvi
q03pNc7tfWAdVKZNHbdKs6fE43beyUvjFvGCmtP4Aogx02aLamscCUfqiRuL
71GXFUWFMHR2wKXU0/LpxJ8bySWSPk3cDYtJHtYNY6F7mbHGDF29WgQFXmA2
3hgbbjaWv/MrBPGnqHLITbdeVei2h+HbtWEy+grNnqXBDBVa3ubih8r8hVdL
Y4Mqn0eiVHLJaB/+t4PpCSRd6Ug0dBb63Gqids/XekISQIa/B7l4TgAmCiyg
VK2t+nP2iYPzh/LqGM7EG4yjG7SgL5XqK4KV+8kYrYIXXHxxFU5b7rASZx4v
Gc9TO1xOg4S6fwmc2/eG0OaARjPSB3n+8ML+LSLBlXJXz7YUHaT/OSYoC7Fk
Nh601KS4iQodmtvU4r1QWJSF+lgwq9fTKmEyBWTnxZ8eS+CIA5FI69w6i7IJ
AJf8B5bONDedvwS9MdnY0besBsf3j4Bhig3ur6rXvUzjRUAiGj+Zr89nCMZp
RTXQglzcNRK0fnTMJPSlEdVeftO2BmBsFdmwzSVK53LjvTTUdmADQnCpYHIf
XHXQSVbhrUHT9ZTmmrJbQNmGLFegEmlohgV4LMuJ1dLF9jutMd63GxSjnRuo
QVJoRmbOgOlWTNKLWd78NnHI6Tdm0JYfjkZq+GaFAvvRIdo2XFbKPnRt45z0
jZByLhtcsD2FEbuT+cfFt0nCqVZCZXsdpak/eDlce6tdxL1MtVxKSOaRPzXT
cixqqejp3AdQ+AAFaCHLD4vlALvkO84DwE3P/bVj7HIzZTOst08SLmjfEQIu
4YMXw9CzVjSJeJ7Z52MM54yCL+Vsvksv1D3AOe29grAhdjZZsOMNnvDf1oSI
/AdHXhzqYZsqsRNUGuvo/y175jTRI4XBQ/Hdg1231JucHEjGOg3DLGoS/27I
n2u8PpmnBE2MDjbEzHUDYoCR/hct2xE5EcaAjyS2iOPOK+yssovTm0mmhS4d
dW8xS7jngDEcPAnIUb1m9dYDt7GBcCVu3J/vBXmZ18NgviqzNSA/cJKcWHCz
4uB2zvjHPkIcLUW15ng885j5PQ+J1afmWExz7JWD5hK0I84YA1AvMwp4hq9R
469cvVWVa63St0IJJnq/o4tf938p9bAKlV6eUbZgh34nfLhcL9eFVfwMqOE9
IfDgia3a2WiKfCIQNa44WXGtFF533iJSwKs4NE+InMTTxpky5tH208SkZl8A
WXwN0EJaWkMOrCWLq5d8sAkz4DPyx51WRqer+l5uK9FxmJ2kVmtL8gHQH1Nm
WtCTl7HM55Org2Dw4MkNE5ggKqPaU6eqhHQ9Y8qlzFQAOi+/HsumX79PID2V
GIOxAGkxGrdUdnKz9iRamSZWhU0sTyf8zL3d4K3e2Z+PBYFrnTwXmrX4TbUk
HccBTVecnGMoaV/YPg5WbUFOvffQBLGLezgjCw4f5RUsDNoJCKX/M042PcqE
wo82eIO3srvq2066+ErmNbbPpcrk1vzwbx2XqO4+dPmCOcermdlagJx1PwRV
Lp3tNjdsi1kUd6u+mjpfNRtM6TEgG9Jrcyf2J6u5qvq603lrHJOY5GJquLCh
lxUueqT2RkawufAG3mHop7hVPyG/nFTFDCXqoAffdN7j8g6tErgN7jqQzBLy
g+lGvD+zbGjCssoBThRkzCbVqC7ULGmopzqaYmCllM3g6by55q2YNDcbojo6
3+q2T0RSzAzksH/3HZ1jMTokCXLXUNPWa87zKkgWmhXR5pGvgXEeRz7MshQ5
LMaI7/ux9/IgBs/YIgsg+7NYDXfEtHMBQ5lo1C0a+AKBEAXGuCjN7rkKYEmi
Xki1YWrztF5XucQBYS554Invf5wUlQpfshKq3gjGpr/yXAkE9koZ7uYj6KWI
begWXJaGZ602p0qXmIE8J9Zu7p9BWL2KtCQk1LqvSIqb3WtIC9ACiG8fGK1w
BrMngAtWdlgHb4T9i+xnqVjm45AmxPmKhzrWXEJmQFkSNECR5j8tDq+C+8Ug
APvkuiUVjP9rziSDy6T15XasmYNf9vD6GikpCwtvyPJykfjw0DsNoozGLWP2
nLGcZupdqH/IIxtTTXAwMHj2AkvWdOPORZhHhfYaa3IY2Pb/4t3rYf1/3YLD
ARgMDc5NYxI8NOIPa+SXTX2llf2ehbx3Hxlh8f3mMwVIqk20CTB5y1SzTBav
VPefawa0bt2wVa5vgJ+DI9enPKgi4njuvlyLMd1vl/3E4Sxgk2hh/Lij8wve
QLWCIfJHuNLWzyUFTWugGWwRL+R/vVoBrT1oLerhYd0zJMAXIjOkqPrg/3f7
NKiPW3zVbHfHgbxwBZmV3AiZ4DFuKcevkcnhd7UiFFRbNnFP/0j0hBgSlDnz
rymN4SnZsvrkqEAAhakHOCPXVT65I56WbrSmbFEgbS2OvgCnpjlXv/knRm4k
TMoWyUKfRKcHH+L/orgceKBVacsvmu75aZHp1nIpBgs2YqkuTfvcQqLDptXV
MEqIb69xjX0RIvABclQMhAlQP+ECmDF0rgCfZM8dpZkFppuUNbjbIOCyezLs
sgMwI01tuFkDsWUSbiZPW9LsCGmskmREmT7SWJ5LlQh5INIsP7lyRvq4NfW/
/JSPXPwy4LGrlnA77oOPXcg1VRwCzI7hbwYsdtiFbXZCf7NCPPVnmyvlH4VN
+fzoifeNuzv+VWSVyw6oSN4qigd8dUmMvWjP2bhhIJyLpNQIF/LWInjC2Prm
jmgwYsuDupt2m+2gr+u5BQ5BUzELn+iQpsYq6901B1O5bMeUefpIArJ541UQ
P7IKTKLQ4ckCfUcJmW3YaX16kO95WIQEgLG9gCvVw3rK8EcKSA5vnT65mLnJ
O+NEDkpUO3NjFa9ZjegOirGvMOTmLKym37aT2p/J/Cb5l9QY5Ps5bPYBNXv1
VMO7c3WV6lEzpjLEiTnzy6GwtrGvc34Gpcd3WTdNputgs+91ecGwFzE+fEj5
omVsfbZvIzEkqe8yDEY5rHyDaNjgRKNogmmqPHAM6piNqkYNckZrQAIOS9qo
7jOORxqdhIglJEBrJyoQdnbD1n19Gr0trN7OKS/m6VHLlvce78Q0WDzRSEmw
hC/P/LCcOjepEvoxHt137mH14mXh5/TB4CqQM61g/I8c0D2bv/82VZi8kEAi
dyWKnYpNJsA/ArO5ICFIPWFflA9jzX7e92bPn1OKScV7IcC53OGCrUgH0Kww
szFvWgsFSj7jTu8cHHxi8JqFeLyb0C3wmAikGCa9dvp7QcWpJwEnkanHjBWd
Tvx78QFCcbdQaOvo8/ONpKwPaQDJthhpuv9Y9JE/xTyThQ46O+xNteup8iz1
rgaiCho2qwVDedfHtNjZmEAhXGsB26wJthZU9F2aSvoDYsbWhx2rDc6J3w3v
dZhjmTBFNmuOMomXDAVtyC8ZTDtTeTd/6dc/lx0LFRxKaEC4CFRY7GoxrKp8
lupGPqz4EaDBFuIXNIsztEvV/9kkhRO8/44yMNeNxWwgWcUslhUeFSakQ170
MsXDMXh0mXO7O6VEgDcp8Ulj8L7x3ZJ1OetdqbXaPiuSMPEHSBKvP3umHAex
2gFph5oBrGWrlwfVjDQ50IvsXlIxapwgiSoe8uoLlcFEMcWA6XWBTzFwmQR3
/Y5L/j5RsJPWRKoHfnclmS8xXIn+0LqGuIu2yYtQxT5kFxATco3uGD6sTWRU
HZxoAXvI22FUvuXkSaoDVWvYEBzQEOad4esStEJ40av0tgDJrSlB4wf7bExr
KAyZRW82AIgsdASkUKPHI2YM9ImwoH5u5kYaEgAXoBwDrdjAUkQD0S0gynvC
cfNWBD5epFwC4o8vElBM38F+jBYRYYUXs4I/RQXUrsOKSWcH3iLv+IBvlRjd
nXiW1SiALPMXzYPKhC6veKoQCI8aghxFtHDfv3jGAtCRIFJ+SjE4dnu1CvBd
m3woLthwilFd49xFJRNIglnTOfkhlap490+RbBCzeihGAizHPOVwubFUpaIk
2fPSsllhebIG7UrJeTFNyaLUDWZ3V3nVVWJPTuwiSwvxuUo/jnHWgdUGgud1
r3nTtjjmaRkP9fDj+Z4mwF326t9qflrZe+yJi7rcoqySAbNO5ZSrHfQLN/R/
S/qtqdpcpk+tHM++K2H5B/zey5kvgqpLldOjjiSHAmeZdHI+/9oiejGMssY+
44GBQneKYNUHTdF4kSbdBPzwFDmsXTPniTv9ZG+v0InIPyRiPJpWHQw2g43g
1rV9hYozL+Iubut3IvAnpfHmSMR8n89eGkEY5pA1jZvZOGhfoVV4O9Qopkmc
DWtE6jk1DbZOwaq0U0SYIiXVlLlJBNMSqxvzN25UJmfHcuxkj6aT7u3cKs6G
KETNDcutpAFeZfzd4eVD4eEHja13FAikUXoEcl2+0ndOs9zHn0A9agjst/An
gF9qwx/nhOqcMrrW9RKHDPC9whQQHuqj2MUL8aLiYMgmfrSunZs4VeEyX2ob
qje7M4Cc1PGCvBSVhrRTyMXezZURn+p957TvOL78NOvSfUH95e6anxTmzxah
yWOTT9AOv3+KB4KbiELOoYMM0ufaTmiKvMHDg0F5JsnJgagWq2kMvaIkx6dU
E/PLXioBgcqo4ug+gBLAaF7THAZocye5YFSbcTk+F2j2U4zcxV5OJvs7HGNl
0wgmdOiDdlsEjzUm7YFIBB868s7yPxuoOnwDDrWrXsuJkSkBS29V63cB6bY9
ij0zGCKKa56iy76JpUvmTs2JbpXfYvi3zUjLmH8/z2dEsHSi5pBl43RHEkF5
7BFNDtADLkWRPvhEvmXi+blfjw0rFlAc9MCjgm8ivQsMYkJziMqURaVU8Z5a
RBQwqV26HrjpoSB9U7erTSqGg2TYS94cz4eZMWdikemh6gzSUkUDOcqj296T
vTNco//RKgwXprBbNdEOMyhmLM8GEwgdBQxpOYgaXNsGH3Y1fIxQNMlct9kI
Jk8qxLMXFehTiIzoxVdQcHOpCn6aeCqIRNM2GWOWGiHNZnmCOEpZ19UfK4GX
2UqFEVgQCzEuC0q+QDSLGG0sbU7v5baMITnqwmJcBXRLODbyyVJC3lTs+2gx
i9h5CZbgme5i7hiPKdm//DssEob66S0qBW3NVaGfq6xKc+evfquqOR0p0s6Z
phRnoLHam/u99qj7jyicoeJ8CjZljfXqb7dWPMjgwzfuOyNdpsz3cu3iYBxg
kbhN+13PKoKmffV88aFjnnGQ1+fcrxxFLgP7WtQcMv+pHKnkE45mhPGfQMkD
RavdDIAVoUxn4crsGjDpnDibUqx9VgXwJRj4srkWKl3CSjjEPSOh5xMmE3SN
He3m9AWqtRjdUQbfqPnymcnsczqpG0zlUPJUw5Sx3WFhh3cHIWpPqliG8qa0
KEA+rc5ZPOQrw1QAGfIa9IteJCCT8V4aLwP/e1Vfb4R5zL4Niq1Q/mwfQK8f
+C/2W6S65qwc3y70E/wRr8ARABMFU4a9RnNRsMK9gzM6dnMUMijVaXWnRvqJ
GkBJdD4/IfwFHKCtKia95vH4Eoh3M24woEEoWJ66NkfB3Jf2ri3+b78l5jIO
Mp8wn3elOiCYGAPGEHGmNIXyXobzfxZ+2O8jFgwM1FL0vLkDfAwoh9A1q8EI
lHDATlCxnRvh1eLXws1ec+YmUGS2s44Agw0fWGTA9K/2aO/9xt6YwZRxkR/Y
6/9PG5+s3xlBdgTLBmNsSkk/5GhtzZ5pjXTmm7KMgnLV5xvey/tVE/+WFKe7
Z26J/yn5+RzBTyeFa0HYTbfxL7xC2S5uPQjJiyjdHEjhY123Pm5LamKugAtH
PM+zMsP7nymqxh9+5RMNtROU+sBWMfut03aKSM+LbRozgQEJxlZB2A37gc5B
4tZoNL9rfF5zA5ITc2FGFbTC7j7hq3/v9T24mQarfS3blnCD2YBaFcmfewUk
SHry5b4E6ffcm5m6vRZi7x2SDnYdlPrXmwKEb2pXXLbKxQGFuHBJkjLq9Y1+
1cJ+MsXz1xP7Bj5+WBhmj5hVgg1t13YSfwveQh2AU7O/8SOtFazcI2OPrmjy
Y0e2QpJlB+7vnj+vy1Y6mMSkh5PC4K0KYE73WngPnFL/79I7suszsGa+h25t
KYoKv1TY1lBLpoBSLFuTFaTwrRM9veoJ0F43WD4amg2fKzZFkEgglK/aM6+o
ffTrO8gPgzEYRsp0oPMQP6EwJglQQUEcjM8G4Rz3rojkhUCPyJ4N6X7T254w
TYY1CGH2mDOhnHcxRJ5z6LhzCkxsoFl46Md/3Joh/lhIwKBTLmvQyXreSjUR
Ru9fFf9kuc552AivA1VVNycHd/VGkQCQ3uU4VbiJFIjapFXkMbHemAvgSNNW
4oKPLGagvBo3OoN5gOXJqJOD3XHHEj4dIGh7DNYvYmFFkZnByyEOCC5UWT21
rHdfdhkT3TrzeeTdXl6ldktqAJczV6ZIV+rL+c7LwTbVTWbKntGLYn7MYhcS
wEUG5qUXPoPgMKVIICsThDf8gLouXA5tJ3u1fQgGkgzfFkcDwOOchKkSKj6D
O1St9OL63EWd44/4UqvXMwlDyj5Dec6AvOf7ihRzf3Cok0BJSrEr2y+Xg9q0
W4d40tvUWSkZNVeE/HNq0EeN93tayysoMto00vyzEvIxb0flm6oR8/Nf7fvx
0aITx/P12OoeKw5WARYdENAXFVlELaJtA5ChPmn2veSiSMN4sq0jFfp3HN6M
ID3Q1FoqP/xGHPFQoGlYuVu2lHXYE2L+LeD9U8lmR7TcqYoZ1T7z2O4wEM1O
8EKKMDD5sT24gay02H3w4IkWdZ8FprWc6vv31Xqshm/9fmKQn4zJLoo9YfDC
Bn+KMwdmaE7KChx/NivdbqzEknB751voHH++C0o/Kw2R8CZct9ImyQcKU972
aqLRfJ6PpM2SVXa2buI9Jj53jz3Nm78A8+lG9ZZZNYbbN8bI7P1M5mFIGw+m
pMtOONWepI1KlhnieGTk794yfR9eHFJHNI3/plJ3HutZ/nCQYSB5eOiG6PCs
G9g6mJQUVoOqYR91hUD9QuYKsHHyXONX36b5ia1gClFVmLVCAR0YCLA0CFFN
rvbcTfPjOczag9LjuQ8HuXwSz+RNKlB6POnj+RmwQ+G6RtK4IZtXReSRHgdn
s0Nsr9t5yHEcRyTZyfGrYItJzsBVd/KfbQmd/F5Lag8KJlNxKGl20I0xWviD
jzYmo6RzbAzU15Hxqr69x+TIUU43sg3oqtmcxEZRFAQXzPV8fNJ14PthhTRt
e2tv7GFTSFtwWgmTqtrClgd6lNNshecXu+0v0dNuc2xOZGyYk/9cN8GvSBqJ
Oe54j2oxZIQni5il9UNoSRFmTJLFkwRy9SGvaRKsiQKwDDH6+x0K/XFDMXKY
5dpT8c0rxAtpmHAqirJcY7YVDZJ1F5AiQixffg0nfi1EtYBXwoV4hvdf6HEn
61ftRo5D/Y6LOap2aV50dHKQoOkPIpUWpTrQP+s6PAUM0whk5Pi75s+Jc24z
Pbv/uNI8KSrs37Ch/RulmvZU7CGXHjNjetnuM55TQ2zWOQ6deXwBEm3819p6
tN838uBthOf3LeHcloYxKVCv3OMFO3nsCCT3dR9S9wTjEM5w8/QnamQ4ja8v
poSWJ+b56gJDN77v4jOiGtsUNW2EdTfoigMHA0qw0+toYAkVlsS572jzv1En
JaHj3i/yVa7xhPNYTDzlaTSeYiIfXO/L5MtYiNpdXKKeFR39Du49YpnNqBGH
EM0h7CzI066yyFg/4NX/M3ezKCi4uZYAxUwHJMgwi6ms+WcovC3eBbdU9pnE
McP7L0ou8uwEt38xMe9+KwnHTqXVGQr5PpPV73CAx4WAFWLCjFQcC94bvD0a
dyoX9ymLaoqrcNaRoc3ivW9EVPYkOa/8BQ7I9GRf1VWN6M7nOvH4zSO4joj3
zhE6ZayiVlEqsmqZ7QFeBukq8lZija+M9OeO7JtdqcoW2ySZlTV0E4lYIelm
GJgWxwixUMyBbY2wAhFTYMUAJOozRCp/xdq64Y1axHsEHGpX1I6vS/felPo3
RINZDqNQk6j/hw6PbOo0Fmql0oQLt+qbHHsCWcyl04eCm2BpHjpW4yZWknBA
jBwfTYm7twmEtsB78PBjJ7OJKrcxdsh2flkFxmQQbLCI7mtqi6BrapfRr5hR
WXdHQR4Uq4z5gWjDdr0Vw32WXu2yKjx6XdHwu3FTD8Thy9ghlyFiO2XUFMvv
k370JTYoLrfpRLPIU2+OcaXeCRa9J9wV5hz14om46J+SKfDnVgYSf+3HG5zP
1GpS/219HPLx8EXGhB441o5G0vMVzY5pJTREK/l21boNkkzVoMMUhCJdzYoh
qEAZiIUH7E7lrbwB9/uNLpxnIrImg7tjzmZb3OF/by715i2S66ewEvtBLplK
tAeq1SPAXokYw5ySRIVIPDGQ6drOLMwRKEphsdM/MFOSQ8tabyf4pg920dMc
RFT9+dKvldNkKQwE39a/BEPYlgbA6divYsaePHWZfoBiFnJsDD1VWrIi6+N6
ObH4ZhvxsmA2ey0VjSmXVaKTXQJzLweLjAqmNL6rgVFPKOaqbhEFUpV5Synd
pE0G1LuCn2ptq7FDGGuu9KWUw+l2lXoDIHThcPUB2356B/8g726Bjv5Sy8Uh
b/8Rl6OHPRlm9uCIdVDDArqAbyDTEGdMQI0RRlISM5tkD8LzFuq5y/Be6DHw
dVOqhv2AhkooyYAWkQBnO7mYZ9xSNgfEbJ/HTRLikfNXxlYlxKnKQYkHoMJU
56lFWThgRqTijU+w+agd0SU0BBAKCw27V1ZdO7VSYVPABqmcRiEWgZmzfP7P
nF4HdCD0/Z5Zuhu4Y20n/8E+xeAwoHvjenLEj0GT6HEJwi2HOYB4SxoPROBC
JeWxdLYiT31RdveHf3vgMsggXcXo3VHnPKkNzb6SaV8m5+/pvaeWbGl2TCfb
JreSkgLpSkkcoS6pdzM8fzAXpKiXI7Gyz86vfP1d/1QKQdiRdVFJiFpKA36r
8gKVUPNcYTxeMCBewuAqiJNwx9iiy5n5vbKt3TZ8Wqu+UhIWBpZMT4slweMQ
wybDnaJykPl3xGuTx/OV/BbO3AURKIgw+VZ9ZsaXZvdewksh0ScX+uhnQe5L
Ci3nVzqXQj7ifjVrFndxgl1caN531Lwp6eeCKJajQYFmU4D++yVFp7xK/N/L
OHwiLh3BDynrLsmhsbHo1VJaqq6EsDSDs5He3bunWJu3Ap3b9DK3NJAHlxGb
rJQZx3AQ9O7gE13Ah57/pRuca1yHxMDkUBClCh0JvdFTIh/rEOZAf4sFW+JM
FD0Hmnr7DDJoJ4T3srbw6ygAuyZzokxcHUsBQ2oHm8+TZtwEgmTeQbKTx/FW
i92wgacH0uSkfhW+5s5XFMgFAIWffFSCrBWtceGUdsQSHJfuVh+TLgDjQIsv
C+SfmFjt8K0uheopylCd8NRdVd+Ei+wk6f7OIoQnJC/FfRIeRLfNt/04R6MJ
WIxXmzmc33zvTaA2IGpYz6RnN2CFKx2yQ7mmnSzeIyOFYDcPMpy7pMVMEpl1
hcvNb1rwjvXCVh85iexdBLtpIYIg2cFQo/jWiZWR63+OMn+c8cPub8aN80wX
/TiW7mgWlHXoSDlWVkCb3dUdCSnhEuGXnQqaYt/iA/nWQjRWeFUS1iYVZQDG
Ce2V7JnPMio1fa5g9tlDAlikslu/q/pO0rkTSdS3IBvxZ7I7FGXWq085i4VQ
X33DOO2cMTkJL6PMAWSBwJXWr3vXLxjgvsaWzxruZwk9W9ZEU5gPquRNvlZL
BFDdqiJHXk0CIDYqnVT8+aVPfxt/ntD9EMjnOp7FE2/+Z+PEF5hInmOF0pAd
heQTRiPheK450QPUT9tuV72ZBZlIkuSjE9pVEF9ATFr6z4ICLyJML9UzTlqO
H9lZd8u3SQNSPXbch4EmGUEKBsQChRFNPS5GXNgJOjem7mQreBzG0hN9U1Zq
E6Kn/18qq5qI4vDicKdXYYyX9toXNTAhHZObbFiq7IKOQpHFTd2UsNB5F7wm
nkPIJm82EQIsHqgmFon1gMuN7VKnaWRq4ASpcbjaPwB7pNuCW8LyCVmjC+Bl
FhKmmo1BeBjEdhcm3lOpMoRSPbMxhj1/DNB1mWHnTn7MyahG/XhFYZjiNyol
t+doKL/oY4U3U1YrgWszzAkk56hQlVXKJlgnBDUo71gg5NVAfCEHwaxkl3bj
xbpsDwwkcGaGb0ove7riyMhAULzTbm4lrLAYkaaKiB3FiwhnaBpbr0g4QWPR
E5RY0krAv/nFrja5w7nGTqJJ5aOB4lnlJw4cTINOL77A1DLOfi8sYK7CjSI2
bmCVihayNTIUU8gZEJag/eqB+xcQVgd3E0v+wjGC/oYUfNn1fBqAh2jc+R7J
SpRJ2XmlnKFWgRBXo4vKFkWTCaOXExGiMX85nSUVc0zmVMcLHXynMU0yDZt4
0r0jLw3BYBFyMJ6yxb5hfIWkfk4bemO7vgk/E89ATQTEccwTXEhajOpZ9PFN
nCQkw928Vamap+1SQZaxF11wD0wlAvbaZVbNH5aaMtxXrANKYPnjW1ia2Tdx
Q13B0CHl632S8imjZ2t5TOpEx81T+HfisTTY17yBpbgLmR7TQaNzoUOCzNo/
bQPXdl+KOMvzy1dQrg2vp2PZ0wcC7RKP+fPSQdMMl15sXfnFzcPrY5LFIOWC
fWYDqutu/mbhbtYBixMpL0IY2vxZYP7TWz5BG6Fu4yle+oV/LW64w9HO5vZq
DRYheKjh0qGZwSeF+aYJ3Caz7ymikSDohp5e/TK1J+W5iVHpEe3UtbY3uLUy
mJlW5lGilofudkspcX+QK0zgBkNIRHMecWZsAvuRtSEsBT8iGoJPHmJ8T47/
/M/LtfPg8vpIWtioZUZNpT/9AQrAYiDySfMAQVHV18ls+1YVpE+it+sged7P
QnVl1s2s+ppxItu5V0PCC7utD10V/Uh5a/UG7tIaxNwO7Kg0svCkjl+SLh2T
eNY7cvMzH92uejKGkkqRGntNtG4gLLG65XGayRagt2NgHcyGh7AIcOtSg4r5
SWcEkKTNDcEnQjSKy2BLt7wFx9t3DpHRQYF5LeiygH1HGjSx1qGiSWg79bBg
KXm1LHVdVKzh5YhunkK+qhpCIweQeEU4ZT3COQplGjI7YMYCHT3I2mX5aVMF
8Xg3r9L3JEOjUarumIYLJySPkYmorPUbgcdgrodZ3KuJ05m3RmpJ0dd0fk6j
H75cPQvxaqsb1WCXz6VUB2E2CgEJln0hSes1GhVtfjQM/eKYoqcOHdin2QjB
963MGBGpx8WQ1DAsIA7EI2MDY8/bsmkYys13A7SX6SRsAy6UErPKP9m0lwOm
c+dqJ1bcVKdKny3WjeWxLROO0i3hJVha9Z66ziJDWlaODavypwCeAE7YJHQO
Kyibw23tXMecP2j68MRYbuEfUZ4e7BkOSkSpb16t99p7fVN9Zdaxtw7aATJi
euiB+5xvo6IeCkPEw0mJa0ydl5QHFKx462p/g0DoFuFpuzjF0nqUiNg3GLeg
QvjD18bIUXMjxxkDos39D5u0p5LCoTvH2DEdrFss/5ZyBj9eyQ5NObSpBu1c
72Lowc0w19Py3FzLEsWhlT3XTjbKYntC/qZMgAGck8i+UflaltdryIAW/+mV
n0R5j5WISI+hGJ3X8apyqbMruwR/sU1M/VjUugNRRbKQmtcuC8+47uVMcKF0
+VpcSGf2j/K8qjL/SntORcgVPWyeov53TrxHuHcIqmMG89INHNGjCUyukwi2
KAP7ezuzhNj35aFo4K0akIZ8Wq5hcrwL8Q6MN7mQNa53eyQU7Jyac+O4GNNy
4rQ5Tbtcb8zIqPiIyBhA79F7Qj+8zgcX+51DSCnGvlAi8OKIRX5HBmxAjNo0
xIgPZSxF7/MFA7LCQCmzimzed2jQyqFnXhxhBIPR3Mm8d6FCe5LhXqWALOPj
LG2v7W2oexa9dSBu3txSMT+mW2rWtjFz8HGCOu+p91EUqWoU8VA1OmXUf5Ez
UPfioIHWhqRIRGF3qF9qpx0hw9nUCp8PU9hX7/x3Yz9XInL41qWomUOKg9pk
fBQO5Hg9oyfjA3uUO9aQ8GeCmbcmUlu5wtJ7hf83DE1laYjQ9YnaL2Uw71sU
E0O2ibzsZiP2tO8ePE/HE7ZAB2VgLnoneOGihqgXuwWfS7FpUscW+9Tz6MKl
3mp5BY4JVoPMglNqAgxv7q4K08Qx1juaDs/H/Izr61U8ckVaw2aF5IiKfuIr
fSVmwuFjND9ypHZXMddmoVpcCfLdCEaVQ1CIHCU0Urtk80+igwDxXNrko6Hb
mumHjmGDQVoGW0LXrxpkLJA4M57RehoHuHWpxbQ1C4u3Gis4zZbZv+D1a1kJ
H8MUk/FQ5b5E/7i32WJrEqIuitFJgWwXmS3iZ68ew4YORecmd0KM1QEuRH8C
NvkF/3F3MFKvGtzInVl5xAqsDwct1cclV4aZNgi202fJOn2XvqWrslsbyed3
vaQGegjCsTXW33fzAyv8yS6XGIzutjtYCCO9CTFGXdxI1rKxj7lp3ynKHanw
VcH4v7XKmZc2YzIY5QrE3UthtQ/9UEcXxlieuYzzS+u1cCADetiCUC83zgnG
MOaoCAqTt/WihhFs8SFbHvkj4Wk1ELJWwq7EE5nmAuF3arymF4ArYsaShAas
m/dp8QLJolVaCuOpa97QK7LmLtUDdacIeyULiNnQL6W7vhw7Bf6K1O0zGtdM
4epKitKmdsZZFOXBWSE/6Xoc55bKqQuuKUSQBhLsknHeDcOGxAsHuXquZrIs
BMdxwavYCxenv5icuTr2Poh8/i1pvHCGZR35x8w7TWq2oM9e1amSP2q+LvMq
RqpaqFWi6JsIaO4l1tRhZSpOC4HBXXRTN5dHP5Kegyw63urmHEqnG613Zqbj
XYylkw3AAE/ZaOEH5BV19p4wRKmqZN9ufKo4S77rJ3RG2r0npV/corEuIFfp
JyF2+w9RiY/w9YqEZRdhq7BenzbEh97BzZ0wTsNzprBU6qc2lREfejMYp6n4
HIz/5O23RWYbmdo79sTdRfvbXRJxhmn9z2bjbt+IZ3u/DiHonkbR+IV868Jk
PYIdnkD+mvgE7ETveENa7x5zL2+rMe6Uf3pyBphO6nIfcHttL1TnAMnlsssm
jYDEfXhcsrA4s9HtKQ2idSuy5l0ZetbFMzPrROOw2XgrU3d4aGlRLCO2/Jp6
KwBQO6KmM7PZNT/7PbilyNVQodLSXTJlk+6rluJr8T5RLBbykmWVcqlXVN9g
CNfb7Zi4bm7kWtrZJSdwOc4rCutKpo9IRYkc42x6ftNoLVsLA3N/M03Smoh7
D9Gslk6bL3NchOED9+3EaFx3Fpdm6hGH/y0jtajPafruNwMdj+b/0VvlghLf
8kW3+b8+3p1JXyIbrcBvET8q/Vdw7vWdVxkUiaG+rF0jTqMB9Y1j+k3qPNF3
AfYL1c8DpuvnNQL11e95ijTqHfBHZgDqYoS/D5J4tsEDF+DGLdBhMVir3/+L
MyW5AUyXLSDi683alKouGQju6FPEFfnA6J0UoHhuQIbKf1+HyQsBN/SepV3K
gmtp363yJ28T/i3ca6QqXn7opcgmd1KZJZDNC7DFU18dV5zbS2bFtn9VQKqG
COq8fivfiITqVZWGfCWWzwoW3ad0tCNSemafek6UxGVZj02ExsyxNd2TkQFP
+zTMnVJfvasxnCKUG0EtnWeyWO7cdGWJExMt72Fx9gX3MZHWCFbRfgJuyzCB
0coOy3HyrasQG03Dc8DKRzdv+O5t04E191cx53ZaO5Ir9aYfSeAxMolx50Vj
+/7jMiQvULfOkGPVVveAs8uk6xNQ1jnJfYXl92trDSm0dRGIKacaicsUvAgr
zxpgD7IByYXq2clQt+Kdh2SDfuP6LPM7SZKtWbS7goYqANKqmO18CM2xiMFx
OocgrFm+efWv44rLz7IGGQTmrAF+hHU0kbCsf1Q6hWraXTnP8drt8Ow6biCH
wfKIRmwmE1B7IrVlRjlvzuNMqY6hoiGV+VHUu+fXt8SzxxRz38utVOPimfGX
EEe2MlBClI8LY8CZrBszJiUirOPs/g2/JecttF3pDwW86qs94EN8pNkZoAJI
J8m/6Y4MiyiMNW4jWAZlMv5ed7Poe+1nvN5EEt/6D4E8MqFToWHPhhqGSaUV
oM8qQzAuFkY/5OVmssI/7Xi/W0ZArO0R5fMyIL0wd7oDSaOUJd/QkCQCtm5p
eloO16i6QVyyyD3dQg0GXDAfU0IVnRXzMRyUKn4P8F+dvYJWUjx6wU9d5uu1
SC6ARTLxx8YV+TUKycS+fVluwVAB/eWM6pCiNAbV0QDPAeXBXP5E4fje8EG2
4YsOmOUK7RDUZiV0iNbwCWMCJ4tYrY9cVBwOoeA3I/s8qP1D0B7Lpmr/70cr
mQlKh5P6/AYGTPi/NGtY2FZOlrv/4g7UWp+gehd8m7e8TopnnQQq4ssbgxkg
FD2oKaumYyIroLIis1F51iVqnX1z88SFL/oCu9XWfHwErHLx+CPKOasK7Sp0
Ce1q4p/wHbEgqAS1L0XOnFoTFe7nZ/5juDPYDKqb9O59lTM2Un2CjWZYDz/Q
RQ4LS57dkC4u3YiwGwA3U2v0X/bY+1WK15kU6+inup3sRjCLtWtIDlMH8hjL
DqHX7ZZQXYdj1g34IoUK1TyfF9J+p0RHR/JVR+taajvjCwCyQfhNpsmKrUaG
qJWyGwh2Zl9Frk+Kv+3uFeDlwD61+o0TTrYXjpCXZAFtA2k6XgDVAaqpT891
KKOHW0wWcQmdqD+OglBuXir1MsV8Jo0cPrKQ9YG80e6hR6OB5tQYht3xUw8Y
+xSD5eEkbWcrFSv6SdhTG8ioW0aq96ze9mCv/asxrR057uzrydpps3X3SADc
YTSn5BAIFR5eh47xdcuf9yB2lsJLd26rQk1ye1szPFjHj1kM0MKmBgn9BSlM
hCbqmoJyH7WBW2DCOC2Q7C6Y+kTQK26X2xHGjRWkH9IB0qgRPBEoYfrhg+O6
QuIII0Y1eFf5FrbMymlBXYQlb3fkYrRXNSXEE0TTsjeJXDfOHBfXDOblWUmR
O1tbn2Xp331SZW3qChPsMjYA+buj8HaveK10kcNUwEc51HuUYXvhSep3eo7V
eL43esuSjkNfPExXx75LnsE0myMVB5UvsxQM7EjLOUaIGvV/c18w0+2ayRim
/t8IbWeOpveniYceXOAYTO8CWCzaCpzF7KsMnX0m7jytBW1Ywd3Bf76Q/7Zj
a+8xQl5De6CX38fQIDzUuacG3Xbk478K2XYy9F87qHbqs1BLmC0p/eiA4rcG
Xq2TZBpMSnt3OLJQga+Dq8Rd6dRixKDkYa2sBMmk5YqaatOqy3VekU65kZ+Y
LhX16V9NjR5Plr2U51f5GEopII2xs4wLs+M108oJrA8K2DWQQXxmjDwc3OoT
LyahhiP7bPHaa+CnD6XIeO3zlGEo9hjSrTcPNZb6CA/+5SWZN6w+Nb1pyad9
Rj8cJYbTHtVBO9vpH3RRNoPEqjde8RcdKG1cF3VzJU0zfBpMsP3THy+YG1QP
R+bCTiVP5ajSgtnsxpSAIPzFHKQPu9r1sCfXtawDM2TM+2l9I1W46fxKhKZo
BymTB1eqZEsnYsW1PgX+AN1yAsbhHlDLJDZXWoaRU3sf8qG4Sy6iQ/x/lh+D
1Hu5g9gwmOA2+VLGhZ22ws3JTk1Rbjcnypk1yNfC+AnMG/GZ4YaqHlIFmjLB
6jBROfjLIXX2WmpsEH3cFYU6L+3+j4EH5XFR2qX467GlZfeEJZyjM9x0V9iX
14X+qanErHzLLf4lf/2Cn9RoGgTSP+xQG4feMctGRVuqUM+ELMocFzgxqwp1
mRBUpsDTIlg4kax/pnCfDHG1hvVfAtEEQ6lZJZEh4fxpy1Fc3qoAqbt0aFv4
9ihRBJHgnb4cP8bbc3hSSOS0m76ToV5NQz0H8wgvz1XaHsmG0cWtb4EzpM0c
XxFdyzT3JKVLrZRLhxDLrEvWfEVDd5uHdDup0CaG5UVwtN2Fz82vuufjMVuQ
8cZ4mhDxIoOsE+d1u+Wmofp4H/CAok5Fbkuk352q2PbjICzK9mwegi1plWr4
3hdLtQri1eAqEgwl+jG4DJmcTddSE0wAG+6I5xY+0Z5DikmuXBUcj8zsHAqF
Ho+LGVVUeVNJyvFUR02v2LjupTUFr0Uhxfm+4LpkxVcMXIW3b1OOMb8Ojc3y
8fAEottezmvajaA7gmbkYDR1KtvwKcJWzwO0LzekiYo5EUK/I7jPyHY58ZSV
2CcX1qPScqL10XNny4fJViJc+Yc2vCR2h2Dmgv0/4VNZZzl7DSk7YsDswpw/
IJLsVAUfvm8zo5CSuRDGl+hE5t52daDK0ItESoZ5cWhWbXoYHlNq6QC/bG4y
QAasXYaYJY8AoBP1W2hq77SyJOcgfb2mxCK38xnU4lbwcIsqMnr6ejDZC5ky
phnMYM54w4obrA0xnhUX1aiYdaMR5PU8Zo5xd5CWyvLAazgRxpNgDwCHqfZB
3wkWoyNlaMuw97Ax32iVMeL482swC5tVHsf2lygYbdDs3VIkhD89UCgX7dYO
BY4Ssjl1UNHQkV6KB9DbuP3PPgtDAa9tyYFH//Jsa0pLSGqEoXe5+y6tXL+7
3bBJP/Eee5UdaPEe25lbAiIYCIXLSou21e8IJk8rFqe71IfYBZ5jNxHCxg7Z
iw2xJ18eAK5eKkn9HZImsc9mmcN7qlvOJA2etv+R4H9rv47zmIui/l5ekICU
/cZJF5yqdoojD/Ez7tymUkaFcwGUg68HUZwftA7ggtKZ1RLWkl/YVmpx6pWw
CsuuqkugfpsN1uVWGzmytOrev6Cn8m1XHO9nH78LlgQ0KR734AvPijAD5xa5
rzqAKVUdCijgm/gRTzERioemCS+zE/2Aq6yZxoFrlOkndLRPSODe9DNW7bqe
ZcyAJFY1XjmhTKsI3mTQz2SSmNH8pPyNyuJkzc5dFQKCb6Wyq/oRnmHTxvUx
HUv2AvxMn/sibVR8V8S93Kn7t8GZ51tkslg8oURWM9cPwHbknyaD1rfZjPss
sHMZ8UmxEbFGuqQb1+QZPPqZWNSbV83an9KTfQzV6UlfA5pMgsDEB8UawmBn
DPd1R4xf1rI691EUEW281I9Kb2p+yuV27ee9KZm+TYlOV66SK8QsRsN/AFiH
lY+p8Hs3HnROlGSntYgW5HJJHkM0/qsYKSy7jeTSXlQxS2EjtYbcjfSN56Oc
W9Kk0vk55HfeDW4dEVqN9Wzn4ifb3bVdFgJxnPe8cH1bHJ4JD1pIuEmGHd6y
0ZAsMmTMw7KMoEQSHS8aDFVejrMuZkggl0Ah9dMZKoY2m0+3WYWc/W9TKy8D
7Q8p5RqnQRogvnCdSOr+4fzi/Vt4Ahjrcj99Yji2aEQFcHHC7+pXZcoeeFm5
tif57NBTMBiNRzH2IFm2P8EhxgxqqtCHY+cHZjB37OY9kSgIUV38LFwALQtY
xB/j1c5MCKlYbqT2VMTYABbiLabaRorZctC8DjjSIBrX+iue8GGxf4lY8hH/
+poG/2bP4P4zpDOz+WoyKJtFSkbH7nrA00OLK1ZSgZSP6VHDbubhhm2rPDcx
ggXciiefc2wt7hzFDIYSg4ljtqqh0GSOWeGdMMMH7BL5cnWbQNZtjsvHsfEZ
4aQBFJHkgv/X95myQSck9/km6/eiNF+w17lHbwdqprp8Paex0HuNQot3Dk5p
zDkWt4oHLh148JLYyyspY0+ULBJNkukltR60e8NSf2q3eEAxP3Hhoia1oY3x
kC8b2lqvn/V7HfDHtZBas5VxXnUTNWpjEZYETOA7Jxx2jYyAHAOLxeLr7ieW
HYx7ROiFGqJuPf8OGAFlFN6TL+kXrSToAYm0WKdP2cjLwOMcLpkXEy4xX3Xv
0QrSTZ1gLNylafVuoVtMYE6X/2xFvtlSqw58OLufrZ99Q2FCb3Dar7kHNNPi
NH1b/sP7JavO81fUjXDoXoBMH7YMmKAPQ37glY5Uc3Ntispz5xrssvflyxjy
ynN6fOiqamKJKvNqxF+FTUGyoCm9e48k3vH8SeukEISteH8vYjUNcUxmeqSX
NMdiGLD3/W+hmhCLhNowW6AnIrHL0+e3i7mowSqX9BVE3M7F44L++YRQk786
vZzRdPc014/ASCM7UmGS+aiJiIu2BUzuIFeGoTlniTVMYw9DX36+f8zT7PlP
EaOTLc4ZgxQEp/ddwuM4yvWBaDlOoZ4qf9BWC1/qzp6OguHJP+EFVGQYjAw9
snoVu+kkc75neoyPFogJbb0w2grY+RUelFwq5/LUU5uC6EI0jlwiRcVXlrQz
TjXxbgfjQgAHxFg+zdneJHZ7NM/5ojQDCk2ECnsrOsD0QPAlTR7SBzBfQv4a
SRzbQVpyFXo6N3RM9f074bWtmHiHykfj68B0Fdu1UlWM0bmHYxJC4sJ+GvoP
U9N09juQKGpKWmtcE4vEC2+sTxGQ8eHtLi6ewslfuLOomQYsihK4sr82NrY8
69ZViS4lAKmA9RG7/ociL6ggZ6jZHsBe3vxLPkBodSKZsRKqJMl8lVOVIdPB
geLawgSMM1tp+4NRZHZb2sbCxIhPB1b+9LVBUs6S4M0J1c/YQT9bIThZrFyk
oKKKLTALSRggBrB2OZqAP2v+aPeKu+GoE3JwQUa41Ru2G+gW+X5AP7Y/sTQx
VPuEA19E+b8PscrGAhFhhhTP5vNq88iqkLqIQZi4a1ajSMS8+OvSNMyBxKg5
1KVS7Z3JLJGwfnNwo6yB6kz8klbn2UNfag1ZBo+1nD3N7f6D+O1jeQ1W9uJG
/oB2we3qsbCA01dU4/dzoJoRaq5x230FysInGKNMWtyz7I/iePXSlmz5dxCm
1yrT+rO2ZHMZNXcVa4yScBXSaQGFTT2+2j2LFygUyDTfgZQLenPvqhspQuda
vB4lQrp81onkUzuJNz6g/SA1Um11QCi/JNYMweczHSqDsrXfF9IjYgawg/yi
/xLA11bk3grqQCoXBZxbYOH0AZHDCv4a07wZvcA+nUZAJKH/C21gS08uwSXO
YgOPL3AdZIZqeCcmfc7Y/NHY8E9zOzupZE7f6HQZbwrCA5IWiYrmDZ0TjaaB
0ye8NEqB9b8fn96c9R5UpBSC5IGfl6gZSqg7K8tQu/4lquRBbDyVGPZR2Hww
KOVou+EHNhIsy4MkbhViXm14DaPurelkVAFK43v6q2CTgnoqMHoWMvk87hJN
tzUJKRARjBa5pduxwFHyOIoW9UlxYujLphuqZXyW2mk4tLcxD9bSWwFh+DRM
RVcDp0/AAoLplcQN/oy13k8dY3d2xsZg+3y4NXDrqL5W0PtB6luL/NdZNiLF
M+B5rBidU3MQWuD3Q/lcZZvrycaL+580EFZZJgrSbVwEl/jXO5AyMEoz28ke
K3PxNRQVy3IYTlTqLiH2q9cs6z5HFfwRJiPFWlmXottoqoEDEPO/LxBb1cPt
L2hl3M2L78/RnTiBzh2Ilp/vuipxYzYIy19W0onvGQYRf6EhnzCS0ZtFIzlP
xy9LW1MmKfbiVrjhO0+ZzEpTmfvDq8thT4clOkRp8CtdLi+SWXN4FXTaeOyR
D2mRTSlACcoURtPkaaOv4t09KV4eTP9Sj5BnNNFz9ubfsOomAxxyQUAR7vfB
MFbwJljU3rqdvE8R/1PlUU4z+N+6zyK69+hXH6SqBLEBiys1rtI1lmIEktDv
O81/Eapublj1D2OQ5G22m+ULHcx4QQ2aD5I6XZxrhTZwLAcpjc+gWXzJO/QV
YlVHz/8aegHZweUCby4tA2SRbosOHzFyQftlfHIiopXqUdxvyqjp72FrqoTF
mmFWnU21BAv9iXVHB6SfPDAlsgDaqFiKXjM1xGzhYbynE9xfjAJx9wfawzPV
6cvwE80xDSYLbzQOM1ZnmRbE9A1JXfLPD5uur3Zbzdd1Jd+kmenK5PLXPmtt
UTeihGIvtnATdYB1tXGlwayN3T37WBAV7SGozrPVAaKr12B/jhKUlAF8pmMH
fpC6CXYCat0Y197ulE6T+yjF4RKgzt0WZ6yHXm5dSQRhqp+/PoXsVmQi7PC9
pfVmjiRN0AktT4YiwQsIOHsm7o3x1oviAM7Tf/8omlQljBEjrGPWfKxVDCsq
+OzhPpTVUPmFFdif2fgNkTbgOnNVJoeF1p2OWgAeve6aYsM0wvMkeqPXDdp8
v3iZO8xh0opjf7EpzJkYHa4TjJZ8XrUvXzQ//E40F7XwP/GsF/eqRKX8d+rL
zBEjUhp0sSZq8hYs64WAf03BO+i5lUgRXfDEVNgzmY/oniQ4rT6ftBCoFvbS
1w5g0hoZNWCvlCuF3dlK29DpBzTHwXN599uxd87dM2hGHvMZifPdLgglACL+
Hfe9+CXFIke6N85x9eDgdxxHSnMx0MuImU1IuzsUVD/yqh8dkEumb5IojEtX
qIBrHdwyxbg7Xt6/8hYT7+EmH9tA4MfrrWJkB9oUGtYQbZPvJfvA/8HOQ2NT
yNYUnoWeruZh1nZseBKJrt6uxOtjBKdqkZAyltdDB/BH+pX0uCm/hsTV1PVh
MeIjEuYP2EcRLw1VQlMJoIkHz7LsZ+ryT8KaKkTb6n0UqiBD6v/WLEp60su1
dTxauFs4hNZCTCH+OXx2enMZI2HcT3M5qC+m+7raHrkMUeQNIxiDkNkMUvqW
rCCmBRQMbVeWwqkdtBUJTrIbAcW89/piiMdSsmxEBPnfUZu/PvPRQg8nXQjy
O9ke8gpVd5IRNwa583Ryd9TRBJLhOpuaeSNmRAN5GhiqOjoTyWYYn5OJn+BZ
8emy10AOTxd8SYaFxWrtNonrtH6eU3w7b3PosmXWRAVlGgDUJmNurKwNg3Mz
2y72SRLM/Co+6z+KNEq4O06XfjPZrMfNRE4EI70IqcdypFJ8+B8fJjBlIBYR
M9Y+tksXIHWYjiwPrmK4Z50XGqnt4j5Wkz7M5ijphIU9VrFyMcpyrvhWxJRt
GM0fZkyWmrRCO3VdjuP+E/L6f4E1kAHrry9bX1KVnm3khuOL09MmLVyXNlGR
xBl2e6iG4LY4r2eqOy0o1Gd6Af96ljbcBq7DVD3p33FClMkZHYnig9i4QoNC
vZeLYKAs6/IkWNBIdZ/9lKCYwT0+n42cbu2KNj8uR+YoonA4Y8QuE9yo0kiR
64gGO1atDrQcjusNdmlN2vaQGwE6oS6E9W22gl+221o9HlFSV/CAyz+sPlvH
LjiCIFSk6HFTZhdMmoP4wl0LPajhSQZNU7tG+BmFtTpt8ADgI5yuoB8jcM38
oX/HTPzUBvBNYK7jyxh2SJJONRBfA82xcLmks/6ETLVNvcp8/BRPt3wgQAUM
8m1/O/RwaGANO1DOI1zspqT+7mMDmz8r/nN97F5JY7yZR0TnzcI5sz9ZzyCB
8peVKaDl/Z8kG1MpAYMikuFyMdvgfLt5ICB15c4aIkIM1uyt5RRmMNiXJCfy
iaVl8WhnSc4AYitt0LGdmvyCxdtpORkcvYxn7n/fmFA+uRHQ74UaZa0X7qWN
D0SRm9FjqmYs8HVzTrLGmADB4MJgxpIsZYu0nNE7o4uOYeDEh8VVWnt4vbDL
8MJBp3CiUziTD3N/lV46tgq06qohqTeo7yjf60se6v8g210N/Xa0YEPbjDKP
ZuHFenRlmeMiBkswVjPniHm3tacWfd5aQeiS1XTxT5G0dwLIhtWhe0KWwFCt
x3NqqN9S8622Dq6eAtDzZkE8LECHqtKcP2G6p8+2RuhcMdw0M6ib0yyYBz96
SASCp9VxizxP2ORS5cuyj4WlSgIFyJo818hmtvUU5iTxb1yewi/VA/VM5oou
/qIfIURLdj2ZV6u1CZ2izHpgeCI7hXUTjH7QBETaqOBk2aWVR7H1z0y3X96J
6C0VTIlOkPAWTpyb46OYcGUbM3xO86sWQP4VEB0gG0gk+GHFMfixZPbi29Py
1ds9NrQSSH/u057tyqHwHRgFDBP5k5W0Jx0Kifl4TJudPqWoitkASTftNkiz
4czUwK2CkPASVPkqNjYhRFpfcR3qN1yeESapZ2mkjqGPm5wuOi/0JNWP0iT6
joATP/fVxGZswy3fbbuj5/CQCI76rEsK2cA1BFSduZl3tOI+kDIyW/lwo/yW
frhoRxQdU0JgA/i+T0orAcngPeaKKxrtGlVlGGQyv7Sk2vB8IwJxXYXHu70i
1ul/G4HF96GAavjduj1Gwxyke+sA4RYhUGwne2kDeGRtQqZVeVNDHwuoveue
r1Bz3vVuX7+PcQVu9ozp70Vt+tU4l1/QVDq5bgnxTdZy9j9vdQ3udzsmgH3w
abosCPJOOVfRVN2MRv6m2LBGQdZSk0fF0PDToSvMj5ecMqY4nIeJuTttHk35
t7mfbD2mAH4CWJVjSx2hjBMHSgVYDvxGm+QPkj8MMQPUuiRzEhcbDFg6w0L3
7jwEetmCnto0iV6zTLK0W0HcBqwI0ibBVDd1wg5XDGvRRsELGJl/Ss+gjAye
YdEtT3j2EQZgg1rLcZOQ47nVSeZXiuw/kS81syXOqI2Rl8dOVwOFmPMUQ2lr
BX0q7hE+dX++KJf1pM3qesfGr1mut2fTdIcuw9iTgm8mnZwu1Z1Y/w/QEgKs
u4QCOwWYg6IjJr+OZHvbTb/41M4ikeVv0RETZKp1ubzXVv5XqgnwskHX1q5v
/FB9TfMsEfLHi7lSyqr7DgLgED65DfJuBJx2ePXjpzEoAv3Qn8+75BK/AbZx
/UW5DgG2a1dxYSmTqbUhhSR6mrw33larrEbcc2po16MfMvy05O0Ksei+19b7
JylZfaRfdvL7Py7ibC6BTZsuQTfIOljfK+AnNnOi85khk7wMw4sw8tjXTexG
oPZIpiKSUEJhL0ttf6W7btERVYTClTNY1FwIGFZE/CSA2bKhv6IwNA4AAieo
5Wzj/T1OKLw19AR+852DpH3xVOceyouW66dZGYjp4yl4kSEONQCOvJQRdAyC
2xDyhGrQ9BVAceLMw4ANUXniHbAtBa6Tzi34aBCc2ETSaiqdl+8r4SNTAGHk
IrjqdSAvyvQOLS/NRZv5UL1Lc8JaPD+zvXP3lUBj8u96DYxMo0Lqq9t0drcd
Y/llw7PrjCWJNDQP8GGc+8m4Ey1okeljxuekP0PUqsOQzbPK7kZ8R76j8qTU
WbFiz/5dAsDu1O9stI4DJBZiG8OZGo8lFrMbzCUYpMrP0hbiAyyfuP3+GLAX
+0Ju+43P7BvxPDrSyUFkS8Nx5RFlMeY5p6dKwzmtAgHwtjKzqlKL6pgp26aj
TWcGCk7Hm/U8ccl3qd+x7Z/llJvxbQNuPdQzhLQ4Dp+ahCUjz+n7LZgClFY2
0aHK9NeXv7X3OB50IkJNtzWsrzwPjPP5lohaYC+0wVsav5Eq5C2l6Ql01f/2
CrEMPhnKn92VlG5pAoNQ7PxPK3R0EGyE01ZuZjtELEAwDVf3tTM1sHkvVvYA
B5KyZT+/PEduZUGs8Uj2PEs1AWehl7bRh0zqGEyTcsKr12YxxpUqWwMKFFz7
53QrL3nawqR3d8QGLcv4WooIj0gqJExlvgTx2BAuQKqj6Ni8dlE+myXb/K12
fDFU5N+DkG5q3p01So1YSbf7A/LjQayUiQtGFfJycMBIIHygFFhBHOyAk9e9
PtX/x9PbpZz3EkMFItLXjkIzPB/Zhq0InbGuMEUFGwjJyVutjODffJHtRYaD
Y9Rii2rp0SDAJZmdbpwfA7+7/Dl3JcddDIjM4aYLdOzah8zHaXbYsJfUy1OU
u7yCwclZnEO+MxLnmyBjxipjUn/8HiiDGgu2UT9O02lod1eHKhgGu4sWFeT/
raSsRfSufQu8fsCsLmBNt+s5Vz2g1nTVbYQ/pD3bjw1XLKJJEio6psoPYMty
jj0DaVW8mXzyiJcry/dzXEhKpCvta1syPHBEX8V104zUVrbVTHegcnAG7t7/
T8jqxRyRVQNSc0iDU5iJfk2hWqwQu7sB5ZN2s6b5R0V8dGQBPrNq8iC5OXo5
Nb97G/IMIJLzwP3SbtBkbI80tqqBSjmKM/fg3XCchXupqL46K3ZQNLbZZmZT
SgRvad6LbX93p5k1RPDsG1CR/KTtz1eSVpZNz67dk7Ok4rtFcn6ayeY+WbcF
O24yW8+7VlZT/xnqGxuqQCKarGhVCgV7Nx0PquyZW0BXwkFTScZuWU+sBw/m
KaqlueM72Iv5P2cwUdlMqSfPv0Vujlcm4llc7Aofn5oLsn7l5CsPNm0M0P0w
QTHbid6YKJOZXOkIqd0IxK25n1/m2o4fu/hyz7O85nGKJB6ZiSz722zwuRcy
xOYc+O5mOE5ofC+U/wpwFX5fep8DowFR7M1RhFvm4NpOFneBdENCyWBxm7bK
k0dqvA0yxOBvFPfKjfb9V/HXBBufy/i1R/OtJOLlJOKqLzlDKLZZqA5QCnAe
6PDM22KY12Bh4RWL5H1FYKVrFLc8V9HtuRPbnDOn4VGXleDSG4aGWVLd9K6E
QX05loIGfYnnCPggIYDchDNsRz1b5LkDHdMEwGjncW32FXQ+JWuvN71DseO9
gKGdKEl/gFePHlAkCiYzxpIe8z6dktPuplvNWkWxTKXcTpPWYbCdZuvkTFzQ
n/BV2N/lHPxM83lQfUIcMi60o74p2vsWrcJ/9wOIodqKD4TroRmz3Ku9fy4t
TUtPJi760Vr2dn1qfs2a53XjCMk8RnP1Vs1hFLUgj89pbrdxSLBORrWzzmXI
Aj6dVArW1YBs3fjP2g5I8LkEesmQwBCS6Lg64/jKJqL1eD6aEFFm+8GPNyyD
2Nxa6xPZXFhSIVeKCkDs49S+9bcAxae0N5QzIO9BCnexcxrCroTDKBe4jv6T
WhgSPSNPXm1YUJDjRKQIMqdzkh8Rxovcy4ljkzCLnfQSmdDVeDPqwF3qdjyf
te0eEarx4H2LLkmzXs0fc9GegsmaKz0OQJ46hPpDnIv08w66WqSq3jKTsW6S
EQMK12xyOgLcnxeZo4E5UpRd/Zv8i4uCEfeIyBrJ77KTrQqhUq7/rLh+VYS8
Dyj2sTvMgL9/nddrmu2vWvvZLObWfHst0z+wU5eo/3RHO6BZ577Qc3nI5oFi
J2qMGVvVVBOfqHf0feKGGFrMmBjvJiX/Cj+7yYjswMmEWwlhNujwHdlp2OiD
/mVYBOniXjwozuOB9LJrC4pbVus04uk1xeSF/Y5p7gWn+QPwyWx+OwQyJIIJ
zwwLizKox11R4coIFtNP5KNue2+Sj5wfybSzVSsvs8PLFSMoWiHLekPr0VaW
/fgyy0uq+dpDhBi99YFykOa/+5BfkrSWw7ENmJ82Czs9RnfXlyjPACM8kBsI
dy8eZwlhrp84l6UhryFaa7MymoZop/JqpYXywVMuNVKiWk1zbvXPQakjddWS
mNZQwP6jX/RRW+1296LjKXLTXRByaX44LJ7WkV8gzEYhtyzHPk/FEd9Btv6H
mofOTyJyjAtoqpqozB2ljSYLlOlqBB4zsZ6E0FWZuQaZWO7vBgxuqm6IhBGd
50YT5YekxoI2/WrhIFxbmObCu3Eh4eJQeofSR8QUNOS3t7v6x4/M7eX1c1Wx
gDeyh+X76BvkK/rAV6a/okbQnxZo2+tM4Tu8V5o7381luicfMk4mpLrazNER
WaAEsdSgNCrqrnyqw0ASlDx6wuO8YtgTWEZY3jg/fk5b6V6VDzqf4NCuIdSQ
F3PnmxP2/PaDT9NDA5MJjCiTAC1OQxwqPwmbnFgV+DTml3ZuuhK30ddK1y3n
73LhRjpqaTT7595nBrKnqBi50YHUNXRPUEE+kPeQJu/jXfZKiVMaOshjLbsg
w2O0AH4NQ4REYqnO5fo3MiYbg/rHQspND80ru+5K1AzJwFzAQOuGGlRFkKbg
uSm6slTmQE1JPrVHxs/9KK/SUIAV1fMge6oYtHUdYFqm8jlE+jWwt3A+dt2F
q6aCh06H+sOICYSvfiHGpLGluhrKQM8BOnweBHF4JT9lba9TXAlfX5PgUBG8
/GDgU3MfpCVOwLWuoXLElZcCTI8ozX34Pc+bYKTcp7crwY4nX3RDgLcGWYl9
tXROIFdDigHIAZ+LHLdVCp5wjUq9YOWuokB8PagDhD7YMPwbPM549En6o3Ax
49eTeit/xIVQjlSzbYRZBwZwkOxcIB45aLkTf/+lR4GyJ4YS3j1ggGe3NO/+
623C0IX8gINqACyx/5KBxHbOI+YZhB8ivPqe8+ufvz8Y10N/Nw8WwA9Xpexm
Oxwl0Ta/MGBdJJBfJftcTJ/d9dGtIxxwCq3NGzPK9ZFOSFGrf9UKCltrzkJc
APuQkVMuuBVkeKAARHaOSkPszMwkd2KH/WaL61XXnyylAJV8a/9c+pmB709M
24YKN8GyzPZtxE5c9qLrN7hkAp0rxdazJw5pS2tSl8f9NWGYZSzXSMQ9VYuk
V9SusMdYxZ1ynnj3jtclJfv2xkqp2XlhqVJvAKtbGBJHOp47R24xYTn3OO92
6ZfkgNA8RcYnJxKJrD9uFS4IaLlVH1baXFTxMi2nx172qdQBq7DyiXEGbQDr
FsqIjcOdxZcIcnUd7q0MC4ZQc6H9hVmsU8wYdjtSODQ6zmx3Yh2dGMfQQpUR
ISQ99ZNV2PYqwjkd7L+wqNKwFUQUoKA6xjbgjBdtrTW9lJvNbjQsX0pDpmhy
d9couznF9+s9Tn4n7mRSdQQKWYfyG521c4/onhIGs0FL1MiXRCEI1a+0zv0g
co5oiPBCb905myruSF12QOTDOPodR/1R1eHBEc8mz8U3jmuTRAEB0xdXUJY6
GTTDVzZALnwq7XJxpXBjkdcJLC0EZLXEjgUEt9eL6e4X2AlgKiqbkChAOdde
Bxx+T8mYcbYHVLQYXZFIqEXwRdTtaz1gC9WkLXoPOereK+Ymq/DYuhUpqfyF
Z4dkrsDQinITLt6HzYBaHkBfQokhY+Dc+PcvT/Mj3lkNN0YjueF0UoYiOHtT
KV2R6ixH/vRztKt7t1GC4OnQNFcEf1pAT2a6jQK8nT3lLGN5QMPjnpcUEK2J
M/weCik4p3nVnHpAm/45ms72jM1KeFD5vbJq2HMM5I1upD003HO1NeOjl+uL
4A9s0YOU3gq5184vIYPpQYwyVVAy67n6vckmbX2OQpmt6rB6FPlocffaCHNR
EqmUDqeTK84SBG4hRBeOG25CSMYUo2fBwPmqSm+vAi4DVERl7wI2pZUJ+IQZ
A3BZ+/Qc1gyp6llPqZJ4tTSAepGQMipzC+mMNNJ+StvfySUgJ/Z4rpEaWRd8
L3/LrNCme5U/xY9W2x0cJOLEpb9KZmEGwEi8nBRXeEGPaSuLuhPPMpocaY9I
ickTNiL/i0Xit0RxJXeNVyKU/QSyVY+lw72qCQLfXC8ufI+DLMpK+nAd53MR
1BgKh+w5NZc/8BlhSWKaPDcCuws8GeZd8lL6OWaObm9SLmpVittGpxfNdqbf
v8b5UssU42KOfN+87Rl20LbDhfXNBpDBjg/uPabWTiTvwoVHydKykVT6GZ5w
/cSh0TTdCZAYk8Zedl7RGBiDvOXwKiJ7+FraDsT0RpuX26BGhfILZ2d6iASb
qYxJKF/hNVXBR1VIqwpOMrH2GQNI3nd2sFSGc+64oKwOu+93bq8dzrcHaJIt
kzEo0R2FfkBKTZG+FUhYfEMV4lj6VsewSurIGX5iI0c4EzOfSgyTkhpfQc5P
qZ2pVpAS9+r+QDI3gX2GYkuVtzSrHLxh4V5BW73sVr9Tsmh15pW26qqfxJ3I
9+8Ok6g0xUp13oKzMYtLsO9UNe47AOuFSHtMq9iOZrrWgDJLQuCUZyQNf5ay
LgE5i+fely2wPpe8h1ACJdpC0zA55hfYfTX2FApCsu2orfU//hUMiD+wMBMC
rlN8MWWWMsBvU/PkzDwnbf4YuHiHYhlPHQnYXZsbTn1ZTfd1CpYrsQc29hNr
o/Yn5gVb6FgTK8pfJeMdb9GxUwsSVKCiGDRJYcNvGxAfLVqT96/x9JgYM3G2
pw7Ocnh3b1RY1pKfaqibD2CTCvEMmZvPypuvJS10eL5v8oBd0C2tVDTn+5zh
bgbU4YLo5AOVotg2zcL2ERdyXSI8H65aamdPsvoHqs3fd7MjaXENY8q72e7z
q2ptcwH41VgmuOia8bg1AiQEDIcZIhG4pwNdlbDwq9hapeVEzcsotb/DOiaa
VcWqY63YSVPvU1lfX93OLl/bp8e5ZsxXMi7HYV0djpH2+wO2+hIVuo8ZLa67
eGbMwD7afYe6QCLirvZ/xJ6F6/bJjrQaukhO70V49cA4/MLEaL6v4d9/M0m+
0Z9eUK1Jkp78NauQ74Ya9rKHJcubLz9C9Di9NsKa1v/L24m4j9v/ALpL2wa/
3xI45DL1Y7E/Z8L5+aXpYCvenFS4VGpIsa6YKNOC1oDWgpF8M5F26SFQqwnY
xGxvrxPMvbyjtWRI7noaylTRPdPuxx6pqS0KMTNIqxJwuGAjqz3K6dMzZWP2
MT0CktkI/5t1RWy5t2becWZWSf1xQZeU89JYmRozOhCwwDu/WuhSMAdAuIMk
D+JnK4BqTzA31eq1rpxdD1u2diDutdmLEN0MUsPnTOKEyO7CED0H/4642zKS
HMPOA9pOA84W1cBFH31d++xJlNGLtBOFIRZJiuCqw4OuVHH13H7tsq9LoHYg
ZWe/ugP/mqNc0Q6AV1u3/jxnrAAiEt36TEPSnyqRdcB04oXHspMl8gcLJB7S
9VdL9a+NQA/r1Bozs/BpZnRhhxRHZHF9zxwsFc00tSJpK6tOVuhDTfZEruLb
zcTEOIWTnFO3Nffk2Pl+OfO32vItUOfWiXhXXzWgz+yeuRZPfxmxEXXZqVeA
FWxSJqZy+4GNOyVsItJ2lLrwjZKmImR8UYT6gPQ3Y0NvpyvupeJrr0kJg0LZ
hLmw9ktgRNGXCPplewLI430HZCztV6dEufi5hA0qTg3fhJNeYW8OYC6wg/bV
KRhr99nyrFn3pLuaZoQYxMj6uODDhWav3ZTS2ZL6VMybE+Wm36ltl8E496Oz
Fi3gms3vNd/g57043SQ1p0jXFG5E6zDD04M2fQ9DFIVXcNIZO4rMcT6sQhy4
uN4LZHW1+PS3E81IK1z2g4zEEuhyLiTfHemvqxvikgpnR1g+VWP/hKl7xX1f
XueAzkKJ1561/SeB9QvLDl6vZxHUb2QvmejusHAoNzNG5miPDPcTmNEUzEWn
y0OCBWrPvhiypAunwAll6HId7VGOekpocf+w/cT19s242Uy03LSMHth47oQv
L7hpWWYM8ccQw1zZVRDw37EDnjb7jcZ/DQa4/7TACJwudXmXnN9vh8yYs2kX
2qoQ14+DLs8ug7dnhyD73eKIgXuIJPCruAQyRRreH148YMm8LR3vovDArFLH
X1panUC19JdZWLWN82Qz7UQ8Beze5sF850tyJROrUXikUtl4DSDKKTlMGf0c
1/3RTRXilvR4o8OLSv13d5MasKGcQXypoJnJSFWFLU24vWXzG4jTjljoEL45
gd6R7GWEXf00b5eh+e1z4jl9kI4HhaqKtBsDOnTlVnXqxjV+SiClB1v3alFA
Mm9/8dhVR5femWXUepgX8a+sGLGG+GQNlGhNyf3PyOL5h1W50N063xLrEyu+
ijTf9mDdZudjp0/zScenV3eoToxaIZDhkBwJffkUdgPKxfCn/nfsKL4toUnA
u9j5diE3Ri2T5hluK0Fn9bShrPLThdqChDrT6om+MJDiE0ntjgyZMu+W3NG1
+P9GQmsuUm9+IEOSlkEeCFtELpTAYyBS3heXuRwDLh/A8dXkcsyBhTazONk0
DBpQKDHBzbkZq4DnLrlcUdnW1nXefQTc3U21Yrj46q3GbZVQw9KJCXV/Ltqa
/2LBShDbPx0v50Zyrww1W5MyM0z/uKI5vVH+heEbn6h7ehrHFKcTxQiOaagk
UaH5jvR+bQYg9ZnNQja0YwJfs8cVZ1YIKdtWrXcioY3QCn6I59mPB2rpH1nA
oQPNbsJgcdS0gNoSnhe5xTOxU28xzpDShyNmyy0HxA1VWanUmTZq4t5otUbX
1Eb65gS40b74cnSZzjyrnu+y7Ti5NytjAqYXh0Y8tp3z/rqxmrItoFAaaOOf
igOktuKNrK0UNba22BUSRDMmtBoeiJLnm61v2y9oQKOKEa6phrgKzohhsibF
lPN4lTJ8PN5uDgafWC/z6urRJradxZVP/exBco7o7hTPWOmNB9czQh/Kj05+
Mq5MtXoBOBSUCW5EX3A5m8fJhd2jC88uMKXFuV63nmcWPTV69Zl/96unMDfW
JFtZrsVsXICAbGqo/SZkbshY4WcqD8p60rtTm9vnSERjEj9e6ICWsT2Hrkh9
jDmwfeN99j7394IO3adJ1/MQcTzYZ0UmKvvWqg7dfRB1dCa3SCqG8y2XLIU9
DzGQhZLeT/xoM7YCH4wgO7dsz4jJaduJlgmZqrfowcvnWwhS/dERgx1i1Y25
L3GOP33Od+54MBAMdlAUeyRoZ1YiKp6OwCijkz+RwLBo4sdDpFSARqxrtony
n5xMuiDPwK1WLYn/XimtQDDVlx1HP4FASWv7lvCz7h98KE/KI6vh2JYyhf5k
ehPbHJrau1AFuk8XEjSd38caRCC1zKBFGBMToR2yRrwQgjszGKowp7xGwdZb
cA4GZqTStRxHyj8znxZWwbtafkSvkGOYLwtrCdaMZ5vy9doPWq1GDwNtBQ8K
dFGzTt8r2K1T0nZ6nNPSN6YOP6eU3LNeSHEJH2vp0P2W13xViZ0vnsvkD0ez
FuxRHKTbCIUOJLjRYtQuj1P9zNyw2AxqPIrDCP1Z70xq3fYKU+S34P3xdSJW
RqRvtRgN0TsgQbdmz7f3Q1d8Wh96SG5+Jh6mJOj42tKo84QjexGGfqnTk6u5
mI9VfW5lprxmxKsvs4XeecDyypqBasFh8yPzm6mpQoUUBgs68n4PspJbOYs5
kG7tMT6AWsJOsh0aDljoCeBBdSo23/KJ6A8o09EsINgwaaEk1Gyk27Ri8WY7
BCNki8sXz3v9KlVIWP7oDqwa16OZbY9W51CVADJHzrgMyjVf77ZjcBkxkhRR
Q66L64jbHlE301JVe075tA7fNxGMF2ix6Gxl2jZrNT5lDCQGo3UwxchjEwvT
dSUIr4QKtYxfHDAzV6P0RffqxLgt76v31QNhPN2gdYdyO1DdLWaCKdW2Wcum
vQFlz3sw+HHl1EksnKwi/fi3rQmM1pdlfNtph4PeX4UDs8/U1oBlaflD0thW
CIaDNGGUK6n7LU04jELuEAws25a+jYPypaoKgmt78L8O3oWwBgqZSWWOq78r
JaTAKxjhG4Gsves5KehDa3XqKdYDLp7jf1qoCVFYXYrm/Wf+HxfSmbiKEyRY
/T3adqVgeCjBwwswbbQzmPc92PsSk6aKsZzrYydAy/tRsHy7UF39SzFdCAbr
IihuClECSBlDaq2078UsKOBw95JB3nOZ5COc9B8sruiVVpcsPnmC8yPIerAC
NfoqqNWn+jf7kxb1nnng7G19BjBj/ghRqwoexlLwWCbVkpMGpl56U1+ZiW7n
qpyWOAcUUbxN+vsPbnBUT4EDnQJD9OtmOTQg92lgAX4R8CucUZCRNOpr8ymq
m6DW5lLIF0TBHQjmB0LnbpQhwZZytgwRVY9gS9gXx6jNCh4toAp3XdjfuyAV
Gjy995/bS5FP+hVowKMEDtUVujaKrJ+w90ZAdcsgMkV5oQJemeCym624tGv2
p1RLHIY0/mgCT196JGwC4HR5EbcYtAVoE/WcYHn+IflsOqMeiu4KlaxRYW53
0QD9UBTLn9c/sLImipGKK6snV8TBJPvEzpqY2Jyufu50pTv4pGOVJ+dDuPsY
kSJ17g65SezAHClo4c0CXTxTOGcNVYNi7eHKVDlJYAj71N+KjQNYInKgIrBW
wYj5gs99TZ/DYLDxW7ihA2CluTETJdDOiSw+HJJZxX4LJ3IWDkmTinD/O48L
TX2/I8kS+But7b+dM0nqsUVJzH+lJfr/yfskRlXl16QrUTr9WHWAuJYydhXU
FfK9C6QjhsZ7k10m/OHlXiCLOn23H0hrQMb7dFcxsVD1Rafkfz90F1F1p89v
F4DvxWcJSRQ2jLE9Sz3HcCWgIV8EP2tVz5JkdRF5LrQF6U2JYkU6i3SH1OGK
ik7+b+fixsOesnykfwvo/qcckeFuykth1o3zKX9+92AY84nF0t2qhOLaMQpf
i85ns7kuIzngFDk6KZib4zNGBjawV4HMCL2y9GTRaBYy83M3MjCOHgJW3gLs
NElsaM4gyTisLQFUORzFK2bqnbSN4rPV5Vi88x1F4A6PYe2VyA3QeYY8vYgm
vxxUamTlvRCEH68v+VlY3HDfQmVE1M/D1Vpjb7/+9eAHhVhS6Gl4gxxmHBg2
BWmyfzIhqpXGpu7qGoDQvLGqMVgsdmVDZmKqobvF9FQlYVt2QxMmdMj3TmdS
io4I+ceTG1UayQ/pkNXDrvG81jicMbovy7z3trTN8dTCZSVfp2/CpBtM8kvn
m/TkDl25tTcSO3bi16dTmQppa1UjlAg777zDjTNMmasf3l/fY/7ayorw+Rdn
TMz1U30DWwKMX77j8TbMVmv9/YwyaxM9y7beWmXrDfhOyfHPR1O5ycr9kUpA
GBxJglaAQIUzrJp+dTahCRo/6n8vZHqWP83Esx4LVgWGIcH4YYQGI/rL+oCf
IBhctwq2x5BIO/ECrbG3YQcc1CMgrmdYa73H5fQdB3OJzljIoE1zAUcEA0BR
/YsjHA+9+yOkmRQQWmtGGAV1ej3BlmyVPy5QyxQOBaVqH6JwFYbsnJezExYQ
pxEFx7Z69bbg1Fbt0E6ozzaU+KB/1Z+gA4EvMH0Fgj1kUxKTwcxLOFLo/2eN
6VKeoRhKsu9pcK/jQQcGVZonIZEmG/8Ha2kwwS0jOY0AdfGKNNi66Fo7kT7P
WLDDRcqrqWR/rHhEdtQ6Knf56lCL4z+5amK1KjelS3/mviAo1jgzxqX7v4CX
xdzf1FrPvJWI3bcpw+C1cfHxNh9Rx9MdH/wJq+JSkQMjy25gzjlgva9JrcxW
1jdI/rB8cSSFRd6hSuzMLdp1X3P2ok5VV4FeZl086UoNC2QhB516JcxuyZ7A
bmW1i+0OE+rYl9casODJSdYSpt+q5hy1oGyrA68rPGY/zpDaqJaFIYd/ZbnG
n6b0CVZUahqYcKNX0n8yKgZuRAFHdLfGz2KDZN0KNroJk2MzCKwF21EfJ/v7
PwtWTd1oGLGhTuzIyQqn+w1+wMYRt18jqAoZ/y1wMF7J4XfbCLyWaIRVbFw+
3JNilwJQA46QkSPFa5ocDf39drZ/iPXyuKbN2svylWlQhBOcLMX5b9G8DDqR
TcQrVm+C5hQsiKCfMNyuhK+Vlq+h5ZsDucJG6O4wYDQVhZOv9Nm2i/OIIyGx
COYFdDOPEJvlidWU0q9KFueklWnhnDllsgHBC9pMELXmqKDNtlK2iaJk9LOA
0FnKyBKf0V6+DrFwyPziUi6j2YKNY6TJ9tiM9OEruo+q7E/0xXVkYo1dOQDE
mtrg6WXz8LERrq2W6JgnkkQTOOjNQQoxycJWUNI0+m3DP84eXNnBtNu/6yqM
47z17MeE181oTrcxZGKAm2sUjVTLOQHEz1veFJciFN3EPEl7EeOkQw47qXv7
kqqkjLPqcxgnFYpIW+a/yL1S2REIEsO3VMQZkzJP7PkUGS965Kj2hUgLxi+4
R9piNHTLdGSSiqKtaCTLagCEgZbXKYeCQEWYwFsr9SxdnnZPRpO6xRDCxEFn
AwxlStiYgHAYwswohmXaYfU8GymCpYzB9ERSikdhABRcf8q63CTlk+aYtd/k
KsqHzNMjQo+WhGuv8+K5wH9ReZqNSxeiPPJdD+xBCbnPmQ6b8kmQeAvimpFQ
5870diwmnWJWKg2MlA0+Flrz9e+IXUsQSBW5XA+7/ZdzKb9WoifWfRrXeozx
urJ1/OgQdXLPMT2sjPRc5EwaNwLPH6zgsVlMProgStuAuQuxxmHTikzGt2rO
sCaQpBcUIR1hRg2tCOuxBNUxP5dkmxL23Vh40BkIPqzjIvco4THAGbaaxUTx
2uoHA2xHy6Xx1f9CzCTQkgwmSwQB/y9/+hDJpoT9DYqgu5dipxFu/VaTL+NM
nYP4tta7NP/KvTrzBWWD6Oz1W3DMhBCZKIXtMNJcKmoNjdw59axMCqbOsdPW
G2/YHykg0tHre4DCbVOiJ/xQijhbf8KHs4sKkWRt1IUTCwMMmKHw8taxJu9o
tMC0uos7liVldv/mwoEwsSIKPEck8OOGiDoaU78sYIjsKzrsTD05VaoagzCH
A5lIbaVvRULJYSjvf6ucpsf/LLzD6KZ6J3go0kBHQMGEgQCk0grT+xSNyBfW
zK9jyoX/hDeZEyR2UXyiU+ZN9lvOQaoEnu1pqHQOUNQtf1VkkFvpa1Ii5yn4
1WLjXWDaukiHC1FobZ4MEyy9xOnH0PHE6pJdpWKJSQtxEZ4hWNSHKdeSDBTW
DlzR6HOgBxdgQnnKj5k4MrSH+mU89M05XSGiUpaprB67l2tVc/dxiZ4Dm0+r
ZwNHNjDW3tDlGBx4DQQmBEyIHJs25krBwyAiPteY8zPqSdu2BN+JG3AsvCx3
/M4ga5UtwLkqbD4+N/lKii3O+Vx8VahdMLSFEm0xQqkfDNyA11CaEGSPLgLP
BlOXztEpIrkiTAJClBCypDt1EGfPNduYs5ml1H9e0rpqc9It7sUpjqYxymfM
ZIi0qopW+jPdqjea5TwNZfDHExV03BTNFOcksjP49AOUhgH8NqIO52rxkjHb
X4GVbcmOhV4QMWyL3zvcdUQ8OxLT4zm61QwFuWhV7w0HXS1re+rxlWbdnbsJ
cB1FZZiEUPnGtRlpjdCpyKcP5a/Y8kzvU2KCBMxUykptvt8f4Jc9DZd6/SrR
qZkwamSN7DwKmJYSrRuep07cty7l+6R25LAY2UAQ8LbE+eTfvfD0lfrkLizC
UEGmE8RtMFjoj29q7LVYhrx+ViuEJLVlxuOVoBIPa+9dO2/5HBZj4n4SCl9J
z0cdO2/gZV1RTEQVfWazSBeynCBjs3WOliYCskNB21WJcygZeRqp7VE7IMGX
vN0qL7AwckmECnyVPmlVYoaI+QQ6L7VMpM3+ZYCA88DqQf+8ViW8e3zPh20I
ukCL9Qv2ehGcwLMKxXlEvS7+E6DDE18Y1sFmNE1cwHFpI38Ns7oWnrGffQb5
TV19uLAMBrimXpkHyG1L4DxdWSg/0jGgKN+ckJvW8iDWm1L+nC/kV7dTcd6c
ODnolWp43qCj5v1XJ3kVTJTevjBTwWKsPhwY1Wn8KwYPfcVWPYhyQjcqsux9
+zgk6PoDF/tJAkfc6CTGxa2Rlf4RfjOSwme7ilBFpkeiFihOGAmvYuFAe4ra
Eyig3qEl4xBdkM0axhWUe5IElcVeBF6wrcyC9QMM/GnFhU02u1nKPqNB4gFu
AIPdUgZEG+LJoyZCKpx0oR7pUwIf63MgrTtKHTZvMEcVoUuQBWacWN9BMUlg
dX1ZshXTosrzgvhuLP2G7lZNpC1vLdrHumfFKMwK/9bIJZl8wmYpmTnAOE/Z
kJxsqTrCzNhr0+Xrqn3tzULTXC5N7eBzQM55yhekZzRxzdTJAPIwxOBCrSSx
JCbpD85IHGgcg693YiyVT4o5r6plg8qdwP0F29gqvaf1f/3u4K2gzQ4l0QkS
kwlI5Ua/13XClRR0VC+35stoWPydgvNSAWWPDyTdJeMGF6lrEt0slGTWYe8M
0oGo8Wwbkq/Flofg7cSO5fRZI0fhnChz4mv+slO9XLhW2E++fu/HsgUKooKu
Is68Rhvt60gM0tXINl2JMKCm/yMZJCA7ZKbsr60WqYzQ8D3OICs6UI+1uWWY
MvsgafpvoDHLkfVnz91HjUwOFhC68v2UJbp4+Cfq7swi88ULgVCBpudC2gPG
x6HrLEgG8kRhw3s2vDhHktXawDvcpeh+CoUaSUMiFebzrsj9ErA9lki4ISHH
UqK5pOfCRJr6xWNNM5xoJdBYYoI9L9zFMDZXG/6ZEljc0FUYKFaf7f5slQmx
b8QtT930yPtHB0nUIifFmKIdSv3wTzNNEEuDkN9RGgRd9tVZMNvQSJBByECx
NSOVoIF1mzHpY04EeWuAPc9uzK83MTYPcPbVtT+sXq5BRqPlSy/VSaTC355/
mrJ5KUW4ptHnIAcLzSvtXJxtIqMkTVQJI+mypq+3Xe80GAtgYVJ53FpRA7Wq
hUC43buxDQCP5tn9NnbRASAOdfQR9/wElAPriWqOcRjYuvYJ3ZR/LXnN+WhN
PctshNSekN6MEAwhxfPurSgNjpcfXiqOqfvDZzYt74PkRAMUW+EKSMjk/HK+
DT6l7M2ym34mJgPP+kPPE020eDRz7Os54tL3TZB/B5Zfsj+I413xOwg88WeJ
NQGURInqDok/F+yS2iITsD3NLBVKzFiQOoaduoh3SJEidWGPsl1zkDvnCFGy
KMxzl8ybO3tgPHne9L9MDa49BayKDVxqnlJIbtVvD+/OlroCX5xqroXXcRcO
edJ3phnz1HVkvNzBEsp1nsEjmNVVaeFGYB8R6akLOkWiV4Pyqw+vNvj+ztEz
JOw0TQO6DH5cKEmhZ2YFqsI41gS+26I0SkrVNDaVaobnbqhoZ2fnSrt5ct0i
DNzcObqUVEargzqqamTl4ioxORtqrT/M6bVew8c4s7I+3TI1utAMqH/DKcNP
jMRnCnRFPgyNhl+ZalOoBTuUiLObIuwDumUcNGb8jLn7ok7GS5ge+4oaKYmc
Cvgee3d2FPel40iEy4H7gOAO9ROL/cFhrQKzG1h11+Qq5+GliF0FpsjANXoL
3aSRKQ/U7DHAJq2sry2FATsyO149M8citlModhQPZVs/PkMc9oGzjmGSiR+6
SDmIEUiGsyWQf/nAhky5DIJCzPqpV5ptc2324KYp7Wdp4+964B29efNWsnLW
4teeDhG6qAnm7bz9e2tYTSTENi3YUTXURW3JitZNt1/4f1SjwHUnDZWoUzvb
pg02PAYT+V755jCZ0HLYIZrLNI0GpN1XfQmXqvLvb3rSjiXeKv7LH5543JwA
T1yfvBbDfbKd8gGj8wfkH1EJ6/quiETM+0Fv74O+uVHAHXcr9++RrxvDCMqZ
uBuVEWkD7OokA5nDGmqJcD5vgUZh3fA1NpCYwoOlE2rnQ2Ijmp1kr8m5/X+g
HeqXcnGGstTGDTfbC4QIPrX7ZsQ/7KfwTt0K0Vhh+b25gzTJgyZM1QF/zq3a
PFQLmAWqGpLZ93pMfFT++1yjvjm642H3Hk62wlcKqxiuVFEib84F1tXnl/4I
s8q/nuHcXoy16kzNHabsdmhtAz5Y51dUo4b378sVB/u/GTvG4hsZU98SgYW8
NYR8XSDd8s5l+PqnpPsODi2aYOoGEHDMg4m++ciWRFzXTWNlYWudy8suYe0i
UJfPEUhriRIjWJzCWPTvu6YjeZ/siSQUZLtO3fqD4J9z1Wb0kCs5nWXP+HIj
rZsgWzKpsFmM7CRtkVYB3d67oGW79SH2iHMoFI+yncYrZWJsxf+UWXxvp/1V
R2i4iNw6S70q2nFzGQUMGQQYDLfhQCjdd/X3CFkttHQDAV3dbyjBDn6DnQXS
mAIYyejCm27lPHTxZBvpctYnKH9WUoiXpnpboIMO3welojDzlEsd3/fAC6os
HOjSrQN0OkiRqxQj+1BGD91lHL9kw3AVzVovnCJWrbyS+r1AQ2ose2rIvIxh
iQarbZHAAr4XyWQjUVzB98CrLpEhcq2OGXZFV50bRcLnX0BxANO11cuFPm+3
jt2G05ItTjsIW3qsgmFRbPmUPqW+hMOm6PGYSD5BjR4km33x7XwIyc/T+TNM
1EGq/sjbCmn/6X/M2dE8zEwAbBaQViYR4vCj8R7CQJ0OEiKUZXDjwL+vKNe6
Rm2+tUc7euPGVc6Xt1+1zDxvQRKneQO2CZgyXyR/rZ/ahWFku3u2ww8veyYj
a0WqT7z1R8a6ccz3bF8lnkTTvfa3zQGlKJx4bt2MmIvy0OJ6GFZlPYR0mXHZ
YZ3v4e69qfTz2Mgip16fiRU5pzHkFQsOfn7gLZ/YYG4GqZdw4PS9N24mW7fu
SCqsYGxaCuaVVnMiq3w/aqcrhgdixCLV6wKUgnKfGlY/TswxakjVREw5J0QP
S3Mqx+rhu4O5yjZGMfeDX/HAgUjjwKAVNkwOaxqwOILVZZFKOAW7fnd7m+B1
eDAIDuOUyhLzHWT2xWBpfLQh+g/cXNyi7L0bD7kTsMQUxTbIE1N95/9/hEAQ
HyuJYy/6O53eXegF6PP1jyj09yxmBsUuZP65H20qh3MXMVE9q5dYcYMu78nm
2QSzlfFfMGUKH7HL+/L01vZkUiWuhS8FGAvhZnWVBEFzmgE79omVXH4ek3IN
kNdpIpgLqzKB/mKCc1XHmfHY6a4Ul6K0XaddlWn+ubqKpMMIO+wdoQaFkydo
PsXaJ25rY4STb4P/0I7+ukU4Il0y/b/40MSby/M5ZtG7fhO1kHpGgBRiIPOL
6Gt6stdcjVLWAWlxFR7s1oQwmsFQEeeJ5fdq6XuNaI3+GlXua7MSTsWX3RCi
jc1n/oTwCIMQ1zuZkGngxmeRNLZj5pxLnwfLbIHXUpq7fkiNrz3livi7ja9L
yisp5amrjz6CeIGdFF96Aml6qZ/cvjoki21S4TbspzwbsvU19Lv2CDXE4hUn
msX+jinlOKrrcCgzrqKzcoaYHHFZrRcKFayIRJwPsawcxndZvGVMz3zkQelD
VxeoOlJmLwq9f8Ur6PiWf+2VZSetZf124O4y3EAopNP81zBZdfkSJdyQ0z4d
K1iUPYDi08gQznpD1sltGm57siEn7lI2ua3S6AfCi/OZQMtpJ10fXZE48ko3
eWgdDuaRK+t0l8TcbqCApWFlTHjzTr01SE6rZZq9v+jTPiaGGBHEWtAV9YfJ
5FwPJRNyG0vJjvsqeoX0TqqZpRjSgnoY2o5BwJCv5oawud0VihlPRpSmfH7N
QjDFkqpCV40x9WETOxfCW1BwIXQAEbNH5pk1J+2V2OVodPrGkzWPlpnOpI4v
82iVpPVt23z//ZaJ4Fb1LF+hYYUSZPSEut9gnFwNB1NhVovFPFfXEodp247e
xo3zMI8qTMasJU6mJjkVi3NnZraCvS5nRW4k+vC5fEEevKLS4xUGjpGKt1jB
NjHdPZopaiMGFSVQucoNS4SfDJO2FlDCmz6VV2UFen2hh/XJQ9TiEvkfxlnm
Z6ahbqJsl8J57jnhO4O3xGtosbVrJSoQemdvhDo4Sh4ebtg/omYTfdb0vcvL
ejGtNwt+0uvLYez5ODv4PxAfHPtr7/TH4Rv9bQyQcCbaRcrWJvVHO1FBdJes
6ScKwxQHm71mczGHNfTQ6CtWWTnf/N81Vzwe8Uun5/HuypRJ/FO0AiQjmy/r
nwkOyVN5pp3LkO7kO6MfY+S62sn1RTRR5XjwQ54ITAubRdU3AQOrZFkiqaiK
L45nuxMhYGwgXq1vWwBjpHbZU+68AZ6/mAKjgYe8Qb4vLvG8iYL84nBwP8WT
IzNRByUNb9rGXW28lqm7/HQmrz+XoITx51UPccInu08652wgmpqBMP5F5vVl
K2/L3UNGMFVB2HJzfm8BbXpzZ/a3k+q12Gecu/SScEQFkMfOSuPvImOt02Pb
3YqSY5INAbG2T0NQfRvD3RzZvNZHMiCYgA5oqfYm2lX2eIf5drI5+1k10hpM
92AXfHom1ugMBlMatjspfiR9nGs6vjwblp7x3gKnpJvthcUqNdw56eVGlPhQ
BU1gsyfyDCSR85AdhJ6IJ86xo7HeHjmdKh++zOSzebnBVJuF5mdyXemXHtrf
q8vMLNwEPhLTrUik2lw5k8vOqKqhS/qSbherULs07CXW/eLhanHWzRsIwgXC
etZjPJOkkgJCQO+fQzI4Ow+IskJn1CbbN8MtTN8nuiICH47AjkpSL0RjEyHZ
Wscv+C0YZ8x1fA/x3Yv/ZYHAlHCQzREchFtYe9pukgVk1M1hAONJCK+jiBhe
1+ck4dpKHrRv9iahUrnF3IIyHrHyOP5pXOsMjJ0pXnsvkvCtkCviONM5PHqm
ABbgtiCzf3icZqiJK/t90TH5/gf5Oxz/VXMJSXe2g3h3Af9IMi13//5wwY/d
cVbVpFa7oTSiscCcRPwureqi2Jf9AJ7sv/QDcO5n6VvuNVX0+7+N1rLdIS4J
ZZfBpN/xdTATAMtjY+V/quX7CVLRs1AlV+o2ewlhHNfokyulYdHZsowt7otm
78uPS2Ublj8RAg26OM8UOg7aITsjTArVUrBEvQbpw8ijPw9WQadUNCiP35jk
W/9ZwQRtbNwM/AchPNJusNiR2vXN6FN0nsd3ZqygD5hOSC3XLrhBfGDFoKO+
PZg3D7jUGsfms4NT5gfODKcijyJmIFnFWIDiswTSAaJnQiQgc3pu2+EAsOXP
Ti2Au0+FHmVyzRyCW6DWEPTux7V3ibXxDNigAsEmdSBGxn9hphG8QILcHrk/
f353kXid6ou+7OaVSAjHnCKGysio+IZxSOXgOdkm1yOCE9D7i80QzmVXAWw0
zj8hvbbYcy2xoRCps1uzdvynWK4NRSS6xbVgKLSQbsKLwGaqPKVgwxBat8VN
9bRJtj0z7Ef9IOxkhVYOP+ExRrg6ETezREku/RJIJa4WzO6kwHfDlBMO9CdJ
49lgPUj4s5uClnGokdkZv9fm9Rrz/A0/cVbq5qD6qymRxcg7COB4iSOBJMAe
L+z4NV91jZiQ8tUexWaxbOfagYAU/Dj1SFy0zmOOvollfnKMv/9tgVtJy1Ba
xJgq92qytcHYTni6FWZNJf+RBUcNQUdKu5sZhNP8wcIYPvY+sw6SMBOlsVxg
Zpi+VjOk2j1A3XlopB2cva6wYewB6UgjJ2rIdXaqbyBrwbd9XoLosmY7rAqg
CyHLq6qJ4/fIc9w652JGRpPOkWKTVmY4ZlYpfXznuy6Mbuo9JO5Fc5ccCUh9
67rjSX2F90GUqSI5rNWk4g3ElXzEezn3O186Ck41xbJLnT9p3V5J05VTNFwx
ahD7PSQQtYlidVkUvsFt7yIgOxx/KQrrZBsM5Kl2ub69sWpEwXkoch9/InJv
vM3JPJ5NOtq/I9Nm4Rk2QZdPxZCJqcBHFJ73tyVsCfCbDWCfMvpQ+KGnGz3J
1f6IUXzF2tJ3aHvV+47/qUgermbtnYEmaPGdNnwSKD3LmVlPpmEQ40mPxglW
AVALMejaFWwtxZR0IqSswMDah6fmbT6Hq2IRTEziYUpGAs0vFk/1CVTrRYTn
fDtHvwXYqA8k39b8wQBTEAPJJR+IzHp0D9P3o0i64O69SudebSeJUyefweYB
wGea5LQJnkfRH3K8gmtA4ZC6d+z/ROa+a8XjdqpBSqlE3adP/maZpqbBF3cU
/gu6XT4OoeNj2VsRGmuRQwojj/DaKdlunGq8jhVmj62W5zEgHXQvKIv/VkXY
J4UeVY3/mMn+/UwDM5M5ZpiOUDW9iGVsm2/EoKOLwmLjUBoL57FUa7sPC26J
JFMVAzpDwtRA8bNX82AEH8aA3lpRUpX1mblxIeq+WUzMXE9gvf9QG/upRjJZ
p+nKe3aSo+pEg67Wle8abbdJSrUNDuxhB52SCZ7b/6zPqGKhqwT4D89bFq6A
/JRhcCV1YJ9TvsePRs4rtxxRMIJI7t21xrB3FIavhJBhauKeiS/ZI08jD1Hh
eB7syUerm1wAeRG8ekGe0RcraK3OqDpXROw/apshWch0n/lsBr6rFe+sVOPa
T2zwdIJrOivaJZlj1YTOknhv9TFtxSaOcC6FTRbSMJ6kvrVd2P8QHrXQqEi3
9Af6ERMc8Kyr2/z6XcIR0e+GQ7tNWDQ15mQbrVWKNgRvGDWI5+nr9IP73I77
btutieEemQJuhbH9v/qbpya5wtLVeIXOyq7jmF1IvEmFsn4EIQjDA1jr3p1g
wwqrNKhOqWk6TS8Foc+KGs5cUOMXo6e0FrmdUG1ye0FL5CbfVfDSORstjdP6
zIr8LghnbK1Zki5lUND3vy2COVzqhDxHQIv0aQAmR731IpouduTMh1uElTd4
Yjkcbi8o1kC3n5+MU0ISg4PSAb15OzITbBd6Qnchy53LIL2IOege3klYLvCG
m8N5In32jyXBoCrlhNBiuLrHcT5FZI+O9Dbev3BEmbYaockOoJwJ2eokpamB
Q2vb9EtwvAwIR15TKx+NOWwZ0BRWxXZO3MRPtTJpz45GAqLD4/0ZwFvYv/1w
iwSVgAgSE2Ig9dw9XcMld+ZBHsZzVX3uz/Fvpy4G6Gqr1sG8jQhFuiNaZNmN
OCBYpb8coyTeFUueuB9QQUgVeBlJ9buRe7XyAscpf6kYnnK5aJTmiAfW4UtV
QtFdtish7EYoRasb9yK62ZalSAyRT5i1J6P6aOi2k3Xd0LCm9Ya2FPkHKWqX
RhYHzSzktrue7dqjath95xsubo50T4zft2HfMdX5szPuyy/w151/MyG8zSA1
ndXxCM8m5czwVbmL6leOReZVMVtm04AwkkXiDsSrDbjIYFEbNaRFyZpzXrZ7
JWoMxPqBUpTgSjHY1hwC//Q5hZ+lVg09NCrGNsYNP4JsrlKQbTBnTyLkzm1r
VlxgoPeeogQI05ZqRy6PfWgrcjwEzWTIt5U5ctnCRlkyY5kc0otnywS8tZ8+
k7lLHLT4najDx+08ly2xzSOmakx3FrjCfgjlgAaSZk1F6Ot4mSxJ3fDzWfYH
xdPK0RYEIVlM0e0v2+Td/AQk5kjCWw02IEnLCenrPgw+tFSd8H2pHa/qr+o4
90uOz7euDw+ZNyPRKwWRatYnxfPSy9fFwz7rDbCvMrOvggwWrVxEZPUFGXf0
7Z8v/8RLc/AZhLMvQmUMJrpAjH7lXgCSupG3q782nMQZ+5JzaAiMozBZksBE
38ZFCuVVxp4/JVIPaoQ01/92LdesNusRv4XyBe6genn0Ane+bHh0YXl65cEp
37B14hV0VJWOOEsSy+/2wc/ix3m/AxJFCK1n2AEjbtyZSGqna/MLMtHWEbTW
A4A3CmAcxJGF4st6Zb4uBB5AqQgyJOKPapLaloM/NkmYE5A9c1PUbZPc07jj
jOPZW2iuZ7HYN8ESb7WWWWOn2pxM+ACNf5vl4b5WjGxnMcMZiIeHq7pgM86S
5uNpgKMmwRWMDXYE4D3qKYeL28bQ8/RlcddokixV3VuKCT7aOfcYdtbs7qo2
mHStJM6bYt4wV47TfwIZvx1LFcRkgVe5hjr0WtlCLCd4q0Dw0Gu//q6Wusnz
/wQqESnNHwa0DHf06Gft+NUIZJn4nwpa5lVS2U26zViNWVq8kcVpeqd2yIay
eWhFlqNw01CI8y2DuaASYAuM7/CJjr5WYZWWaA7VvcaP1X75rLurvURDc7mC
ppe52rij3Tz40tlne8/cdEpKfq58CJd6FiMPU0dUEfgBCoU1+Z6wNgbqYtjQ
h7zsPO2P6xs5rpX+qsBzsWOPj9RY1QbexFgqGKnO0qM6qz4ySaXOPdwMKlQi
0MsrCAia9DlriFly4YSHZb2NuXCbxxp28mnuW/IBh0kP+hGoWuW/yJXs/tDT
5aracSD3TvMLwAnFjLRkBPySUAEXj/wroMum7SXou/RzYTOtRTKhJfzyH0Ps
+4kfCybLchiKXRXonlp+9883539VMKRlQImgSFQS0IheSsUTUDGTDmEG7ypo
GmibjkTuNxBoxM8WYzkd2FwJkj+VImK07m77rXbl7AA5JbiFar07J82Eh6GY
otQ8PulXlB6I+hETHtp/4v5XQNNi2KfzcBCjmrIJJD6n9m3sOtsNcYYOw8MQ
n9fL28qj8xzcsldWJANH2o+jaRBCFFOw8P0p2Ln+4DgxcIofM3CMEG/HY+0R
f/SejVbncOEo47w7UxPh8svXpzxX/Y4QGjxTErd9V5CYyy7EtqpJV8qLGkT+
VY+ZiLhCFA0lfrBKjW0v63fhi6nvLvamO37tRTEnXdUEosLayDmMn0nPhTPR
LBhr8KljiqUQ0jmTa529vjRQxZZn+Zp2lmAkyMMhTg27aOPv/ZhkED1u/ula
5cLuUkKyNFw9mx0CJRBeTJ2cES8cm9Mn3rZoGJUH9CvX1Jd2d63fVy6syf6w
mNyzlHKdditogxtYeIHdwXV6d4W8MY5RuldHi7wJ2SCYlbDM0wNW5Qz7lHq9
s2vjrCQk2pVyKY3vpYI/KIAbc1RmEuZMx1dFcjHh7mncRcHYobNOcp/EWCln
ezQntlyOqkB7Wk0ZGlbkvKWcVD8ztS/zlExSdfDluGeGe9RGLyP6Obk5oD/K
qqbqg6j8z4G14g0ifvkagGAQsZnfB3en1COgYJr+6OvjdYtHrz6xMSvb0aqj
7oSppy/DBrBOXdlpYvXOeP0JI9MiQ5JRI70XioD+iVkODCTtbAlmfJ197GB5
yD8v8RBlNp9dvIEjTgJxFAsQ459yk0r/6m6MVMAJDMJf0R5f7XBaQoJtP3ZW
EDoMw6peuMMXsEe16YTEwB7DcJ69Vo7M4AOZgUqe9lhP4MSCrKljPoXqNkbP
7q816HHu1Eg6oCBgFG5SCmSWrDNDH51FidNur76EmiAFWYYBlsyUnuVXcz5O
XN82JC1jvjzy4fqFaB7Jcx83I061VnHUBsKq55YpzJmZdtYieoJ+nSsoCrtA
QI1s4OLpHJFBYs3rUU56jFKlienXy9C0/rBWhW52ibUhRliuWizASoaVEjcb
3lOfB+Yepd4ZJhLnZ6WoCue1J2M67cEXYLkHgZq2EfAhKvin4Zp5/vDFN3qw
+ocM/BVxuM2vUEY7E0YBSZgyGl7+7WmDq2o7XdPfKKIdUdkoTwkGmKnSidRD
3h20CIt5tJ/xj6tiCIqlu52BiuQPYf6wQAxwIwXjWF3Dcxz7lStC79XjgUjP
FVbTLMXbWoarS0Ny+zROJ2kaLd3I2dau3e17W+JRknzbQvAWTPW/1C5hiloo
h/bSTT70F/ok9EfjStl8m7g8Rg9D1/puvM9tDLs94E86XYJpZI3yXi+WOb3U
P8hHL55o8M1Oe2Y3yE7I5g3EzZ9lk7yHOCbdzFDqx731iaxL/0EJYp8CSG4a
Tgl+jQ2mnsFPcDY8A8JYwk0KMXHtZd++9qIrcx2a7szP4f3WcgZoKfyceGav
CWd1iXnl4W7bhytQcrknqhuDFzsYe3sy2PoBSv/iycsri11qDsE79TAOzvIp
nPIKseHBU2PzZ7CP5IWmOJaKYZeqYWj6TlWnc4UEje9LmfkHXdGAbN3kEa/0
G7mMYlNj0W9yzFRolpkj3/5XcUKWpu4cUWzXrGRpbqoPSW3/BvVvj7octgHF
EWmmzuIxYlShJACrGN01ATi5iH0MhDHgz0qMq8McKDtKGaZTnzBaMWFQDXm1
BZg2CFh0N9fUjoEOqbtUr/Yt1Eia6/U+OMJMQ2JZzF/OcRV3mD5CzjVeCnv0
LI1cds/t4+BDdZgJdO2WOH1/J5qUNHQydKLzQKmYXPaXFq1i9vOHI6znhYzr
7m8V4Blz/ZwecxEKT4F9neo5vOYm5THyEUNtFWd87yzmRxUbZhRkOdMZsy81
3uEvgNo7zvrkv/Zpb8aZqbyCsQovj3oxLMUeWiqwWijMkFlEJpzK7e05K0Xo
AIDlOXXUsRCldCBzm2ETOkz+rceCZWqwi9yu+HEp1L2OlOUA31S9lCORHSvd
UFZEH+HqrU0bt9OC/LMi8naRg5wjB6u4IO8dOPMh8fbtCNt/62J+4+/UlUl7
EnXzC3U8SgHwtx1PLsySMOWGZf2JTGrSZ4HdJtmain6NC1CIyzGGd7mY/50f
Ax+NqYpJ+dTgV7JmZHGEaNnJds0Bfk0ZsEJ6e+4aj2Jxngu4/NSG6VtJbJLe
SmdPuPM4m4stWU0RWIhuGobRezZzMsSbAxIkQlM7JGtKWmjPOP1vKlRVOJs9
s6rLyV7LDoLK9SXhM9xrpPo137GQaBuhy7DzyReLAT4CweZvQ8pKf9/z3bIX
sTDd8W+tQreXaMaxEDTJdNStR64zWm8ObqRsgWwH13G69eiqDUoB93h9q6xj
ld4uixm0408bFY+gb7a+hIPnsZCQWs/DdmpRBqLPuGl6GsqfloIkK0FP4P7G
Fb7EhNy6A55pQROCqCjc6mg9YcZS2ScK+/Zm//RVHOkYxp7B9s7mJRLiMJoh
ZM+i60MucgeoVH4r0viA6pfZUAY24XkuyXT/nCCxVvnPN3sKVnnBpJ+HhEqK
0nB5D08H+wwGRAVG36bs/oNfP3OKk/V1/Vf3+IW2uUgToTcOhbuxt+3RLeBT
Aa3WuUAGjIdO5M+nR6CvIw46PEh1zoZ8k067RxDtn7Vg14SnthXh4qnnpuvn
CncQOwDcX8OofJzCz0i3eBTT2BT77OGCk60LwqvtdRpff4zy28ivDFYeems0
WL+vkPbZ5wGDvW6g1JQCZnoATS9r8FeBD07gSSXXkEH8q3Ibcd+LUDmcYhzj
97CWAb4bK+DfcodnN8whmOxCBLgrQZ9g3cqQ86zGnJ/lnmEcxcTm9VDorzac
gZkfj/qmswtrhBPrwA9imV17wkPnEyNIDPvpgz5X5yKhL54erVeSNu+W9Go/
q8i7kskrm1bQAAIeXdY9tqaZr8qhkgPgCqrtI3hUEjxMtC6c3rElrwlvNVGC
98zLg6/VyDhvPMb+8Km3dnVYEK4vxoaYXi1sfZDRRYAsykE2BKDk+ZVQI6Ko
QY1g1akDx0isOTdflZulZMlDvyHYfFGz9X6lHgnTNE8dj/okJxlzkeZ1Xjva
wcx1H7Mi1B0ePGFo+NGREoCACp62836gKVtShoP7jJ4dcrKFSxJwFOButygO
v/Wug/oNRP/XQkQCmSvGwbwlSYl8xy7Qt0vmnoRnpxX7pztazzUJjn9aktmz
FucqvHBa175g9yBuegVZmZ9zhI83cDk6z2X6gUKMfJIpxM3aP4YXaTL8ODlW
dURr39768Ptpd66sTNrWo8g3nJ0MwDwPRFKrclFR9nG4cMCT5lU5MmS3GziV
vhAq2wWJBEfhCN8HsWrnADOLml4md7HSD9MN113np1O7t4KPBqsJKoGiXldF
e1VZeOFOOw8MmeIffQjy0NFjF4sXiIYz7CCGlD+JG6qHBdkfGqm5iOvTF+Fo
p46UNsGKkWbb8CZ25LkkwMSwxTcOdmTOc0lFIo3txzzcgMp/ZzSW+3cJ6WcE
ix3ur+iY885VLXm0uKaHHfhxePJ5tnwjps3yInK3+W2FQbaPVO8cQUDFUoK7
/A34i7OuCfeXMtiZuOLvR0jtUv12fVqrYRLiOr/61s2MmGChmlWrgLHvP2q+
hLBw69dqDVdGSQgH8Vx5nUWLbpqrRo8z3L6rK5nxomGayuAg3Da3FlwLfl/B
yVwZogMLAAKbqkK+xFoW1/uBqEZeIx56jrqMECjceJ4FLqPXMHrwJIiF4bns
ym6FcSTGhKViIWN8hiIo+gBT3RP2iEVc0ki3LjaBqrJ2oqGb5+T4hg0ujNaa
Ui04xA6ffgyeddhd+k/48d/ypR7C1GBiM+xJtINOfx9Ri1NheARvCl4DqoVO
9fn+4YOkaq6xryIpMGR9bsYd6NFcbY83WtFFK7xIL8CdkKlYHlfFeQNEECvQ
Dfse+2sVryDcPiBkG9LZck8GvjN7FKmECWHqhIk5g4+3ivCfGujrlm/M7er/
7ZQ9u2UU6DMA1GPHFwCjSRgwX4VfbC1F89se5QBmNHqFK9XVUKo3wTEZo6lz
8OjBOMHyoc9f7idE3/v9pN+noeq1BeVa7SkEysyaL0j2qgOIOVRlDY9MrF1H
rNM8EbZWygRBlpPVWm4L/zKx+8iJZPYsmQpQbnK7xqBmzoDqPvVj/+3nSDHL
8jlhuupT7DsUY/OlOzIxITM9/W+WwuKEoTqBw3Rj2KQ620r8LpT2WM04nka/
iFY+q/T5/M/0Ds951/3jtbjU9e7qny0Yr/Rt6r2KUDXA2/zogo9ZmFjfsE7E
sWTr96Unz1zIU4zIDdk370MKKUmkmiD0dOncepLkUxPEaukFVJR47O9k/Uly
JbJjSEQR3D5vthruAQZ+rZTsqenhP2OkDs5iZehg7/yqkjIqvZ6adb4mNSDM
l0RnDY5MNYsR9pMhdTiT1AuhupOyJ8x4QCuE6h+BOcZiO8pFjqqKW77mVwi0
XB0/W9iATw3avJd19o1Ct4wVzRtWzzUT94X0rnF+n0uf6VAxhAD1wH6Q7cka
HihmRtNCRkOHNFF6un6GyWiz8M7uA80dVWTshPjlotAdY48QP3N9jiueNteK
AFHGOy9mUmkDuFVkEkk0K8aoN3yhcwUrumLLV8iwMhHQVeJp3Mh219PNW+Mo
IML3DVQv7EZg+DR9udk166znkl/YTwqjCoSHs0Orjp5ZxQJltl7aEhArWTW8
9UK77mJAYHlzacDgQkXhAW3iHGOTdSkJpBzUcgly6QfuMNeYq8p/FjbdFYye
vG56DlbPRXbPYNVdmBTVIP29bGz/6MLnv/6kmc11EJNZY98fRxtS7a5q4z8s
VnE69Sbm+vsqFbMLjLL2UAaE5ZQEivaiV1mPa1Dpfv/Hp2SnP3oXxlKqEbql
pQDCJa+U55bwfVkZN+B8bIY7JRhk1B/dBnirEP/U6RhnVVubyVhj16gCJ4BV
lrwfXeEALdDWCrr2OyXu/BUhOzxAEuV5h7TzWe2vXPbVePPVc5rx5m9oZHDR
NmAK9/nDqULXI+64RuSlkNsg+6geqZBFPmYicGmobARwqPRXhhQaj/dFjAeg
HyZ2Drm8qC/kBZt6fsosxQjZKS/JQEg6pX0Z/pnC3hNw4GL/uKFHpl9unyaI
vpCRw2P3eUfqk2tUzvo61mCPXaIjrpgRYHWIqXPsd8dJbj683uIIjbDFu4X+
dXgi2lDv66iML+eIP0Yasn0uaEUOkizT67GbxN/buGK01tTGJjiGLVw8YStC
u0irSlzlAc5k+Lu+J7fwBK8v6VS+9sJpFp8ygHgmHhqbOyqlKbQrOpT7jbQY
1oePG7AbVPlCIIh2hheoVrI2j/eUm8oZ9dEDzvWpXUOKT2yttD9GZwgXEANB
bcKdLfTNQlJEOmKXnHHuUfuLkvDMTaenBcuqyafGEkWCwVlxvNrF9ensp9ah
ks9Wky+mPKapxYcnvJ/ydsgM0VwHMUVlbDP1gtmXIBbzuJcNykrmWLbZkDCH
kdccFeUkqA1K02V8nqmKJKHtTr0KSiI2gE3jd6MLsMHREj1uKUKyC2SiPVhR
nGX6lzMrIRM6epDmMzWrQfh3c2ZZSuY6rkjgSDWyZ/g1Dpj979cExT9iTytZ
2T8RHGD7rxz5uEsV2rOet6syke73WKWoKAiYQbdWnGJph3RWDb4Gv9+W3W1n
gR4eNRrl0z7V2HpIghvimeqkUbHlJ0RSBwTlZV5t42h4xrRMHAKHN2kau9LP
Bj3WtFRs0AadnFOND5HIfnrvaIOcUHyXJiOM5mAxR57llzn7G3LdYk+xtgwY
iW4DTkl5Dcwl8XyGK/F4yyYBmOe0cjRhPxkiiu5116i/HIxgFOowB1ZHGVtj
d4fc48b/gR37+JoNJQWpVfTalueM0cuMNBtqndb3bz2gDQ6JoOYedIUibPSg
DbL2MSt1p+E/yUStXqE8xYf8o63QiPp/6qen/OIfR3RvBSfgbe1W9iuex9aK
+YbPa6va89QgjUA2ymjQe+bwyUFEFCfRuTuLNIqmxbFZCsRlhOXXXlvUSJzj
W9ev86I7T9Eii3thjpaDckqffb1B+xngmlWPDyDaWJ/6N4H3JKTcn15X6Hp7
KZCbkaXowU8afnO2SRaEUWVlfa+wMqgKyEVV4tO6iur0H+AV/hveRPiTFn7d
neRGZ3eT0xj0yHEZ0D1lu5tWWpWkTOXxlE7rT+u9cC1GElYboxun9DmKgN6L
py9wuWqKDsqsCrM1zKKSIB2tcN43UL82xyXKvz4SFK98IE4UPvvsPKRTxH2h
cctsyBqDHXe04wyEGCnPNKeb2T3wAVWXn2CtEhtjMvRXrnoQRXvLeSCuQpNt
CDl5VnZCPwk9cz+G3OlRJw8kj8JkLLh/XiiotnjNkSMRqYWwcP7SKCRMPedc
SKsj+lVQ1iYQWuuD723EgdH2/Oq4n+A821xMAfQzsyvu0Q5QhkMwhOCoUyEM
TnWMWFxDm1d7lpBuSIfB+uGzZsDwu7958WnRRLEKUDUkke2M1nrnJMRkU1YR
Op2+euztDE/Yqyo8nLg0nQ09NR0ziVGTw6dieNGr/Io0/jT6IijMdLSJvwuX
UK0v24fd1fl3/66MEnopaA8VZAedWVxVDjF/RBLTfwYkNhyCo7d9AuEXdhEl
QIo90glipVDhtXMf+zybIyPmBjWvJVDdfi3QeB23ccYMAo/i2j44V6GrGVUo
n+BVXXcPE96jiRTGW33h+zKPcOZFmeJbSZsgqnzrqj9jkocNWD+s2NF/61bT
kDc8weu+inAR9SSReRK+EHIHPviBsZvNNEtvM5skclP6XA5D3xeSTa/q8PLU
pLE/BN6EEFHTH8JufLckFIpibusdkVllyMzheXvXpUp01M7foWRpPNp9eESn
hFVeX6iAg/EH08MUEUSZqr1jCJa0Br/hLre6mnvlIIxox9R8BY2tCDZwQcsE
ZAsN7q2FxOs7RlDIIyl2JGxgH19h2d7xJj5keJCrjLLFBDZ4SelKs504Y/UV
dH//HCvLPNE2dfhsX7nlhe9YZsCbSaf+3dW/ISMbqLiLSS0JA/EsIHqPT1wo
jS0Uc3godbf21MGyQyeBBEtuqGD5qevmoUoZTdHpSiV7R2XmoollwvbtzuH1
5rqPLbYm4G9mzB7hA2Td774YZkXS6B9KEMqsMdkOFuN/qHafuc4DircqoJyF
jY7A4spqaR1MFpA1I2ZRn7fsmA1vuwnGkQoz9+SvoF7YIszVJUZXTMsI6hjI
mUOTNSApw3shCu06bz7Dav1lTxETi4PAWEf7mMmU+/axepPXuOan8XUO5v6o
YMzvk8YLZ7qrOuQR/44GYiepI8+pBmHMbFTVkzLGxfaILfWH39DiOUBI1gc/
RGdltAdteLpeHL3ptnNwDPbvzioelBkHWEOfW1Bn3cYpUY7+1jE1vliMq4Y9
1ofTzSr8ZALzJs6RXqM=

`pragma protect end_protected
