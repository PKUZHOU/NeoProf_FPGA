// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
GDcHGhUy54aWeXOIvHEcKxjMGtR1gEApaTlb2n6L5wB9oQqxSaBh3Awg5Xj2ytWX
fOUWyDY+uiBLzItxHADYuH6wovEC0DLc8GlX7e3XixnVnpFydpip1tRcWn013EsZ
q4I4Up0v0b4QxxPeEYmbV/PQZpjQd7noqbwmDNh4KZFDAPEJSG/kJQ==
//pragma protect end_key_block
//pragma protect digest_block
yaoS97E4SxMxTaSNK6OlD9cfNww=
//pragma protect end_digest_block
//pragma protect data_block
VugCl4aXz8Ywryoh2SQN16j8yXE9pBh7Vou5SkiZ39O8Ld+6EwBnJjbHA9QeqIg+
jkzcMtbpafvrq1kZfX1grAvUIopPNYrTl8DVc0nIHvo2NVKhiAWT9OG4iQxPgH+p
CnxhmbLq0s6k4kSgvI3YifUVffEKJBCzQZKspd/zwtE6nCOlRi9jvjIHLQWsTKLI
0kHPZ0M50/Avv+ABpbOEb7t5uqtRyU46C6hN2oSCr/OYhIYpzdmrvIJkbXyYVRbA
W/fpwB8we+Q0j9iqrz3AoHT2PE5GLA5893K0f5ysFDvJvZtGxJYJPmwUQp20Tpki
hKXhWpK6F7KNZIAhcS0fpl+4MJTGUWSC7Dt9ivSz6LHtEMzCkZzW4fLpKjS8Sz+Y
L7GkXQCZicqP76xh4A2t4anJKVqbuMnrjxxr5SQTEN9PlQfquOi30GwSuvbK/uQ4
/1ZW6shsbhOiqQCN7pl0Cbxthvag4Az9+ZwyN1Rc0QzYH7cY5U6TXVkvT8qI0s6w
A+26zH4HHGv27UiEll8GlTo3q5FEks4ahYYEqIpnrnQU8m3gqLGXUmF1o0HYKp5c
qfLsrqB2tq0/SDVrnDjMETyUIFDGPHb+RaHpmwn8CIP79S2RFyU6NFvevrygNHhm
IjPsHglP7aKpUz61jEVUJvEIsqeKcaPYgu6QrZXFTgn7tCEyAGaK/jpn1w9MwBbj
TAVtyhwDNt95o7/hjbnavQXxoiFSboZcEH8W1BCbIxe4vhGMwTO/btiJn1v24G+G
OzG+WlLlnDQMpipJmL/lvqxZs4NEovMIldHXjACA3W7RU62c6sOApymyR4eD2jRd
YHk0n7nq9WhY0xJAGE+J7XB4CJNnpBtn/xFjzgtWV21sr8CJHmbxrJexp4xML6nW
q8hKhsSnOCIo5OIaqTOjJCjTBbfR2GuB9moZWce0xLDEuOtoErlwAQHjrL89/TEL
BPfS78kWoOAF9HAkCc85vxN/w4yiA8mu59jiJ73q9nTiPIo9JjaQ93zegKeIIe3i
qWUUHD3HH9FbPkMVglwuHML/bw1m9mkmAzZMKcWSSSjlSEAYoD+jZgk+9ysobnlv
9Ymo3ucx4nZBWSnQdj87Y0mRRNYU/KmJQJZg9dNZQYjQYNNaAjuRVbbttTLMbEEZ
F/JFIEFHAZC/PaMzzhjSdGTTNvbr2zFrLgS8lmzBRW8m7eB/eexBIe+onSY0MNw8
B/YG5F8g0cIJff6gGqU13znKbhvjGoyjL9mZ0jKiu9MXsymapR18fkaraHfRMjcZ
i25NjZIUxXgtqn0iec6jLogSTub6nxwUn75fcfqo1+em33fAIxe8J8gnJyWU5XcJ
9FgWTLtdGzaVOeoqbI6FecZQKDDEMWgvUIasFmUgp58mawsuMCe3IB+mSM3a5S36
IkhIwDqfM94fTQt7xdwVJ6eWTmhuUhKaybE4L9Q5TRhpoMdPSO1IJGbs0Hfaf6D0
yloB5ulZJ+S/ma1Htb7awTfUhP4qYir2BGvcmrZA8pHIslZVjU7R3aJHZtnCZqzq
voCh9MccP6ASFcX0um0c58QmchYkDjNOoxXdSnTNV9pCxY7qXfNSdebULoXQhSAJ
HJTEY3ZLW5bg1wUIfOnuorTzXAjUj830gfxmCb+BUCcmoVRucogxKkHCw8hsF4yB
jD3WzX525Mnx9jscEuL9HFCMzERdPkP9JTI/UxZy1CypYZJF7lOXPbf7PD3AuAaB
QUSx8SXEJ6We54jzvtRsqjqwztwGMmuflAKe6IJiMotjezzVtMrp3qXWSvUvmBi7
MXRxlpJYYIJ5XyCOiSWgfeVdnO2pzCkFL5bit9NcS2BkOnF06ahfm/ATW6Kp0tvH
i8RKl9TPckeNNPGRDuVIf1aBgRZlyXfI6czAUHb/zYITOYMOinP/XYI8wGrOFHWr
a+MSf7Oq+7UJGee5JJFsPLzbnNq4VuFBs0yKDccKPyKqEhaMS8OXltIk6r6ND3cn
/opPbO2cK7XCyk+Vmi5tofHrtbTdnOaaYtySBTUI65JYMOMHfk9eUQ3OltPVBpTu
Nwen2Yafsc981QCo4Hbp48RqCfu4zmk9zY9S05p1eiWSiuTglqn9QZtR0VJJpLbh
v1OusGyjRSs9MWpQavvmsuUH4Lo3B3a0V+OEuEL+faMUyzoX1/Qb3c2Kt6tsfOwt
D7iCh73y/9Y+coYZuSPkPlShTejYAv5Uh3RTHmW6ISKYXQq7los1nBBvDUoUep8u
f4gY5wzPQvgNS/mH8PAG4gAwFcZtc+X2SfsVoWntTmm29hgl6sOCQG5eLv1AhTHq
83cZpN10cyvQCPta9nRg+ikB+AYxzMbi7MxmJJzDZCm5Oi1TKOBpa5J5QqmRlvLl
97wqEZRC50DJYg6EVV1QHSvj9dh7XSVKVDpOZgrbmOeEulKlqfsSQA6EpFVqGrkU
h0DrivQb4AuJe5EbfilSFMUz3OM6PWdTx/IAVKEHtzzrMFtT97+rtvb9haDg3bbH
q9CpZcWSHimoEJSWB0fvLM+fG5magtqXHkd8UTZ+d63obeY2Vv+KkEFjJvwx0v3+
TwRB1XkmZ0FhwyofBDg/E4e2aK0sMvZE7U0kUxRCZ0kM6m9QamkybbWDMGBLaP7c
fDzhhYJ0LY9c2nmEsYKSJHaTXZWRVtfZ77iX6rrHaH7/eax+hICwr+nYH/J14vSu
J9qr5xjGD2pIwGzxgUKGWRmGLqSGXqSScHuqMiU6fY4mab7vT0vdGwahLiSvutVi
IfHYi3MhBeD3GC0ajBkFMn+LcltWj37xbV5RDMDofISD4oXYtoq1iuxS8R6wf7je
Gfmom/HE4Zwem3FsAALwQT27zsde8/JFiljlXTTgBQWWBXJCS7c8l1psUs3lmXZ8
6ZcFIN8OHG1amHAAf107W5qlq6NOHWiUdlDbB4MLtEhbjljDUxE12EYE4fwq8NHQ
Kknlqui61Lqt40GBdJAhjxk4+2Qc2BDrRko1L5RIytR4xVHye96EWIOu08ZxgF+9
FTbjnAnkrpH9H+MFx2EyRrxfn5wB4HmzG7iuRo08cILGeq+gdaS9LbA2U0mfV8eN
iyDBkPhZr/bEwCmGLU9Dj+ExH8JnBoO7siRM9X5BBiRXlkeqfT9B1TuqZk8qAU+5
NtXzMSCbgGKHan4JO0+WEyancDnRoKZMxfila8JHHJf3YFs2JD2hQq3qVOZ2UQEQ
v2FyEi4kKkBq7nyURJqzYoiRMMx3Zp/XYTaIIIyWhdaQNewL9/u+YlnJwTbQWihh
tyo6C9xZifZbGhM8lUSId7gXq6o1O4pqoU8ngHnhJj7n3gJmiODQ9m+amqCI09kq
E7YjwQaA8rqKAqt+xFTKbpblHrVWOll/oY0XLwHhbvip92S1vJER7dMLuEnD509q
UyV3tu3C3QQkcI5ouFNaVqLYejwg74RD0ugJVzj2P68YtEM3mNOYMSRPPJFrVSpt
7rpiBdhH+evscJJPcFJu2cLJGu+CWYmgV7bHaPOsHzYUfdjhExMk8gmsng0RjPLA
pZje4BvfUzu5TQ2PBNwcN6dGnZX9SmoXLNJv1b4EH1jGYgdF9ZKxbSu2Q+9jDZXz
6M8uoCK2BxliwUZ5GSrQuf2o3Jo8CjLcPeuKHu8mGP59Mb5LvZzBmVVgv2o9cjfo
fzUmzKElyWZ0GFuuwPVFXsAVA/qR/cXYzrUSsXpSFZ+03Qr0745dKiYrSC34gYm3
a8fdSNy/jOIuhWmTlh+AXdL451bhmHy4SIsbOWZt3ZLh8qcnpKZ5WVNAiAwrTg6p
1h+Csk1ZpNDEMMJiMA1WzNwoEg5XU3jSL24htrgy1xGR6rhUiwAfCk/ATyStum1J
0mKXRTWNJkg6RmFH9tRZjEF+C4lnx6fEwjR4rszXvGbaCO1cYMvQSwUkhuCv4Otr
p6J2cJXZIIoE3ToyTmQ+Oap21ZiZicxZ+8BOFvHArVO+9FjT41nxV1wrBh4dpmL6
Nn0xfrLyR18z55+3HpmDMgRSEqBT3425nakoUbJ5HY6g5r1SdMpWMECcAkC7c+w8
LkEcSg74bg2N5e255n6ZoLY+nE/XQdY/4vjvWRcOwhkUuLGDcb7HyOLUBSh9NmM/
lfQ4/udxbTwXNsAd2Kdjf4heL1u85nwN+OODwe7BAL6N3y0TbeuPd9zDjYc/bvDT
mFS0SIwrK7+pofJGAKuG+wxS0R74OE23oyI8WLzgbKKXto2vSnn6D8JI53knd+kv
NOTpoj1vHI9E3oAWrOQyX6pvv4ecPm0S5QfkjLlqKuvCAezViCXqOTM1A2J/b01w
YJ1ljavmB3sa6xLSYpJ7JlQoGpzQmKD76kZLaU0bTtOHp5fz6wOa5z4KIEnA5oMr
DRFoDb/F7G6mWKj7nJmwTjv7TTswWsKprwyZFbXvzkOxg8vEpfUPGRQ96q1+p9kL
BHw58WaWJWepnnuLbv8OW+5FJlhDTxywRFyMYGoSp4Rherd6YoFER7c5GaRfipvK
YIi1Y+8osx52FbAmnMsqXO+xEzvugYlh5BnEmovCymbrgnbA12KRW5mtK3FwQNP1
Bk+ncU0Nr2al9rPtsD89J0QSELXEbOj/u8jH9gCyk9kbVoW+n6YyWVmstjSIHByB
7GUrCi3xAj7dYjhlvAakJOPL0KyhOi/WMKps8hawzOHkZgWgN6YCnsR3jgQXWBMM
k2N5mifzkPWUemavqtuaneMvo8Th4z6YiYvP92HBeK8JEi64OaFwq4b5ub2Xydx1
QWBsMMMLv2Vy/yUTnvCgIUfw9qD7ABWdxWjM5raYYVpR2DmgvW+S6gFOmrFV3kWz
9O8C5M61PQPaWWlg9Aha8rh3Ma7UNLYiZ9Ow4b742h5g/sm4+A5yrdZx9FfsBLX0
jWBMyeLSQEXdetwzKN8/FboMAFIfWMrk7RXMD31mrTvAM9t5mFV42DOsmrLRmv3k
tVOXVtYvCDPQpSbyln3ndn/K5J1Q0XX4rrC3m+Lkt4etnjDcUQenctUwKfz3adRO
tqeXJF1Oi1s+P78Ps2TlI5p4Q9N8Pf+BNfD3US2Jf/xqvlsH7CZkJP27NFIhba1B
xgoOGEj2XBGheYG1fYBCqUVH4Lteegn8Pg5N0vM1XTM0aAOvQZ8CYJ9Ys9SM+JVV
zTH8AGCk787sKHVltlUd5GGM8K0dJ6vGZEPzlDyYsQq6pWPx8eo3Ljol7hDKzHtX
R8d+HecZtEny8Eh1oNWCtu3K2aLQH2HKzRAZ9Vr2Vl4AGihsdCPEr4uOd2RDNK8D
rJDR1FaMKDZfVwsUTOaCiP11W9XeyUEdXphNW7ZnV1jM0S3Z28zc8bDncoxO5zAt
OfPoVJ3W/PVluXuY+STKvkt8UApRrRCtvnsfw+6+6HwjRCrulrzLjSgUG5+bnJoE
qr2xCTkFsGWw6Ds8WC0s/DDa5lZah36jRcfwCZ9FB2L/000cz+jntNwiuH7Ny1EM
fW0Z8UJs2dilOTi330Owymtr3xeAqghgaJL6m0kFi/dfhV/SGXhzbD137lsPEuvZ
WA/CMpmXMa+h1oDx1EU68eSt2jjzjU5rNHlzTRHh/HkExhm+xIBz5I+eOcrEN/hs
mi033w1OdximjWMiJC6XJO+PaCykgqdLVUEKO7iCz4CYDV89kDpAG2SJD3m2tbBG
gGQ/Un3pzd2G63z/3WxvmryXisypdrQa8gbEj/hjIR2xb6V+r3HPWdIA/X5COP3L
tNOGDSMDQf69N4cmpwHZYRBBWcjEJRccZwvstGU0PK8KEUCef/eBNijwfVRmZo6c
9waNWVHzpsrtatE6hCdyMw5JKxUXF7hJkQu3/dfQuz4aa3pByHL9U9E+yX2DAHmT
Op1YuOL8U0i1k52RsZPcirT8VuQvS2/8WcAQK0oZoWCg5h0/VI54iatczpNe6rcp
bycuPoPo0qniPv6OBUZMJc/KMuE9meUAaABU4x2o4voRusFOKRf2QJmMXZq9Ze7F
dWXHlApVSfCVUb0idSgu8Svjat6e8dnTWsJhYieaIiQsJQu9vHvutSi7XS1gYJVM
brCHChJ3XgSPJIHYZMVpGFVGxxMDcEMO30JtTaiO9MBUH+U6suJJhw0TG/luQE1U
IAF8Bxb36FSxSOiPzrgH/u9BviW2SWpAYk3XV3Pg5/NQsKfSRRJKnp+dlldwgM2T
5ZZM/fWpTjRx86K0xU6PkzR7REKPu7dwUQzQ6FLZzYCDCUCCQTxjh2+l7mdCxRV8
WHeyhB4fDwqa9eigd3PDt7SI1Fb1Dwzphrh4ldHpEL/9k+LXrFO4cV7Lf7tkVnJ6
nkfeZG9LwFI9UZ6pU3ZxHp0XJgmVYpxsWstqoS/QbjydIoU+Uu6iNyqJ0K/Vp8/I
IH3VZpRvIoA+dJMOUojRB9+dASsMrf2anudXC1tmHxlvG2f2s/GznMmtawaBKrNJ
jJdxyVjhilMqG66foV/wXqNeRg25rQVq1O1B3c0bCenjc/BtnilqZpxPMfGUP87W
kPYudKoABnBTVYKXgYpbCuhpytzsuNyJtCQ38tgEydaf2RNv7kEA1v3NCOyxqLDk
SQehx1CWQdojXEr1JdrhFIgsK2sLySawzJqO0DX2G6X+0fz/h2Wts1n8BiXrF1yO
TQmcfX/d3tyKAt8BPd4c9Wb0iSCEgJCkzfpPpfAeuxK/dAdJJe9+tAiHQruSjNGx
W2A33+7c3MFmj6xMbRWknc9RndmlnJ1jYj/yPDzk0FyPaV1M8YVTRlrXLvnXstjU
+0yp8DhLFPXvzsTmkrNio/PMupuJk1XL2pt8cxz1HPbqKoWgSR/N8bva7qXS3zcD
NoRY7nbBys0IBHJJq6cIWyNgGI6fzzEdo/E0WOYy1KU51ARMhrca20WNNhTtO9ry
BN2gpT7w6MpDhmVZ/rFnjoKdyALA1bRGmU56llmLJtBEnWQbzXUpljGvaMlaB6NO
aiJZsh7sv7JxpEObNSpTl8Kizupc3BheiGejsM3yk8i49baa8m17KevsUz71es1c
mHyg0jcaRq9ibwHC4+OcspVqKtPAYlt/q5lopPoomPNXf53H0bqgo8RjS9iHRhow
1lpCYmmuo/o+gBY8PFWwh+UDJB0sHMC6YG/Dxf8kMvQzPzKtpvpP3+ABNSKQ/Olf
80WbHQ7ZvFueBVnedgb3ClueUSjnLZwv+cFFIdnBCyHI/CJ0eAsI1vavcp7kzX78
QCrS2sk7Je/E9ztymK/WVx73s0V3IToCijTDJFcdg0GhVCceQ8INZLFYSUfASBJX
WfzWf05waYxn7lCWzamHqfPgMLgoQjl2ZXkdfaa6Y7b7PwFbldYLAK9f+ZF7eEG5
iYdRaXvwOaNgFhjKygAGjk47teiQuTYA+cea2DTsSu0Gk+UwcN/C5IUfsjQ61ZFi
aWDK+kEfghsATy82LfmNJuhhNgUOe0DyFof9BdMsJ52X3WDLZhOtBPkLNwig7jDe
TI8tIpzB6aa7ZFip/LvdKaeEbi8Ov0z74TUKdYTMkXngdoPzDNWJb2SCUs/2t0vQ
kUNyl22A+blwCDT+m+pU3QHi9d8ysJ3ByFo77Q2mk2aCqwUb93GjC3F/hrq4RIba
LDTJ9v98PoXNX0YtKNtDCAejtPjdvjHhyXdoIUwCWajuRtGZzJ03qbMnJDI+6I3v
clXeO8cepofcmqhanS7CK9gqWNaskdn9u3PpqUUN0DFn4HdyBjgHQbx6hvhQTfYH
qJTNrOiVrnDjAeQ9lXqRdLmOnhJ+/JRpupTshWZqKpxK5QsQAJrZYozrvUvr++2R
9LMG8aSxeRUz0e/siaZ9ssZ5Zv/WsvWuml2nX6zlFTvHKu1zgm0JRDZevStvzD0u
buYa3RFL0AVt4MApKIwkKH1SnVAnsQsee2+DIt8HebhV2+qyou4NvkMzLsXUqdMg
R59jHRq9PCcxXSobM3aOY/x9YZv9dqHfDuDC5UpRLFjVnesIvfuZUUBsbSUMx2iz
8k8yynFHQtNaQXlXcKFNhlnngEoTFX9Tdf0RqpUvqhi0K3v557jA9lK4mPZtS5KE
JR+F5+oNTDjoJB2vjD09K4eUZAzl3g7U5gIsj1wu28m2S6X/uwfzsu3XYqkC6Dsb
8WcYpds3Dss+MwZe2JGVMWQPGGTf2u0akRmmYC9AjjT/lj+Ahl5bOWys+eZ26+cW
AZpCwvwu4vn0DWP9ACfZAPPlNKMM2TgYS46D3aMBSwOX6JHhzQ2ozdhwrTxzpbkq
s/LroMnt0mmziWzAmAlUMrB5LIl795g3Ksl6BgW+mbxCoVqi/Oc8mJWm96jOrPCO
YtmdKUQtj2PWXOF92coEYn1ZZKd6Ha4/EbIHE/M4LUlK7YWeUcyaBxIa4OgT3NMZ
3Cue1ZvRT7+CUmGQj/KNC54H6qURfw4zxGCa9/nEfCjK8v9LdpCI7JESvMrvA4+B
jfoUd6qmyXcocdV0dyTHl7Z8noryihY5KRXMbh2NY2DP/g10YAU/ce//siuSNyEi
myt7Su1FEt7+r2RZkwXKRjwFjAeTnhnJj9QilMw9TM9kSR3SJ83QV6DodVfbPmMi
61l9vc9r8cE1kglSMW/2V1zUt6rn8CzMIoEuCQzMaOlIdew9vay/32CLCmRC8g9J
ralPvHvgM1LC8jI7+PmkjBP4iNLMislLMwThCibVJwSnf1135pPkf0FFQdxsB2dJ
rfFxSp2RsmVC2NWGBuTlre9zHTL1ONozljC/JwicMjVuwaZL5xXtUxKSz6R4zCDt
f3hXk/G//4iQ3OX9qiCa3G65XDHvMS0CmlY4OYZLRYkEv/iRcyhSM/RhwVICyGIw
mRyqJo4DeSHhsVr9b8THucxJsWB3akictFn1OyaT6SfXfoi+eU2rbXEdzPoXksnL
dNI30eX1SESEydKK6CYhqab9h2L9fwVOjDdFQ7k846MRnSNOAwPnM9PNOfi4Ywzt
zoU7DJCZruoH/eJ+D0KLDO64MkkpNGiomSXxbrVD8R7mOWTAZT3sqSJ2SzE5ArPT
+bsMTu38wEPYpG8IGxWtmo5KKUDrxcHDlgcSFHDrJuRHDMjQIpYllITdeuJo3qX8
ru86lVdT7cBnqkoepISS3MVUMPwUbMopDLggmwwalEwYNqm5wLcNtd1TgGqLqZH5
C0eTTNHXuNN2JDxkIll1jxFpQRW9mt08xBKgOLUqqV00fGkmUpwgmO77+q7jnwcv
k4RtZWTfZqPYafPEXVMjdlLaPDlL3TZGAdxVatVOnOVliJ5JV2fCAVFKeenfdMEA
RIbOP1+u52Jnh6zSExoXk6TVhVHIaLhLw+YM+DJc1KqxyT5hDPy0YEzfCPKDaZqr
yLaECn3BwuMT0EGiYTyzAxBCTym45+4FupAxPTDyiT+TEbbC2HQBCYCurCMdIIlG
NDQ4dddAYTjMaq5q/sm3QkFMEReL7ukcvOVCdxBOIjUH41BleKE06Fj6v/cmLvDJ
lXoyBVkerYIwDWPegFy76Wd/rO4wK1Q3ZjVkw9KqvDeQO42mBmumUzALA1DXfjZH
J3loFYcPPp2qx4QXxQrfFI535qjIsQNhRoMEKGUKBDjuUNzteplnB6397lKKUfjY
LJpIpe3M5zyNZDyMBQzWNd19RofkpZICtPWVgqBSKjaeHZlyyRY1cMQUPuECcFb8
phUQuQe2r+e15V0QAPTzyfEEfaMMVgQdQhuAf8Nm6JG7CrntbwfjhdRhrDL8NH0b
V014xpc9E9j/06tITkfCkSBIKYNX6kG/f7AFd95bfrpxWGB7YjISx2ITXwcgPFs9
ICX36GghBVMc2AGRzzY//qUvPERRDjgc6zsGug2GrhVkcJVpTCi9WtLtYkc08572
LM2Q++zlbjKM34CaaxjPlNu4u7uO1hcDDagM+cMUoZJgNPwp4jt0/zsTrPRyO9O6
5pUXbVwRMYGuzmIhXu7U/DE3PFhJW/bos352WHgC3ThlNQ5R55Y+EAIeeLn9DoDP
WnjaPyDtXHsy4p2UcmwoABuoiQ1L/JNx18TSamvZQ/NIes0giR1OICS+UiM5SaYg
m5bD3kwcCxtIZJDk3hxb1Z7bvXHSSyJQ+YNOJ28OV0jJkwOgYwAQe/3EhuQmn0xy
SWL9iNMkAHPEmI1REBFCjKpVmgspDrSuBQO7QHHqFFWWqOKRpbeUzeEUO6GGsOnf
rfeLIU8yCAdRWcVmhNDv21CKd6Udc2MSDzI2+8Xpp2ar4V8LdelnGLL7MuKY3qwU
6cazmpVk1do/acJ9hD1ZpIAdCwoD0lSTKvLZ7loSkHFAAlioPuABN8J0rh0QiN9A
7ZVy+HvG0sdtdQcTnge9I2fMGTyO092OiBqixASs5svyNoSjPPZm0/hM2e8sZKk8
7qHEoScdIbYdDaLIatV1syWOlkegxFbsV8Y9jIUWmQWEoShVLWERTRmLHCwQF5nB
VIxaqNeramgtM6KPg0+O/rXkx+mVVwbNfQUgtc7eq/xzqnvzYsOeYU9G7JnIQuXO
1ptIi4gR5XT5iQTKoJl1bfGMFI059fLnwnqhflijjSQ0bN7U06ewi+5TyK1EMNDB
ztenqB8esG3NaiA0T3dRsSHpxT7Lu+718tpb7a3zfO9EK4QSUW0n96E568hVkAA8
VfIC7s7CTTDZFzSF7xlRoVuqHo923VJiSFsYNbtvmQXHbvl40ID/GSMdBfdUiOrh
3fynDB+9KWOaxjr09O4gb4AXDKeFPBAuhBk/0YYEdfEhz0qF0hFHrieFsDsJqBh/
S+HdbEPMSJ8G4JIPLElPiZza/JpWu+66MXiAPzU4ftXEaGo3jDnmEmgDAoGZMUPw
SVpZ4yeP/m2YllCv5zg1aqeroaK0y/bbeLQsbNerUA0Uxs8EjpuBmUDDYOicT9Tt
ezZMqtCOfqtS1OQiTHfMqcQ6XXQ/7h/c7NgiqyjRQOhKS6e16re7nGMjIBrWG+4U
VLTNT54LuG03ug/yvtdeBos0BtPSecuHp5GXVbS4QtU/PbiDFgp4uAVD3uQnXV7I
h8Oaf0iJiuwuwX+lmZd38zzMJMDFumUC9XhpwlTsTrbAkdl0hhLPP9q3ZJB5WR2C
AZl5qWgb5qmo7+cCZuADQx4uH3DqS6HNIHa5EdcidLemF2slcJekiTsSTWZstDS5
R7tDcE8AAN9pQs5mZa4EjnG8K96PwtHib4MJc9JT2pqD9jqj+dEdcLuqsvMsPklk
34wsY0v0gSSeCm8RTeDJ/gZCUzr2gyvbXK8XJYyt/428Idi6Je7FNn/Nr4NheY9m
jF9zi8DEJMGAqPeYA2fiW3h+QYeveIc4PjNcJpUUxsiK7XvQNwgrf4AaYW3lgeBw
vm42yg0cPqJK54siF3sey3cB9m/PMIccvnLx0bmSgBR5YBDfoQQzMvjI47qGPfrj
GRTkIoNyhvsHN4HptMt3/li41iyqr/tJq1omE7Gd4DDzsTjzLHkUP66lguFTAugK
/Eu/o/VMnBtPHtF8ohgoElNQSDdkWxEA9Npzu+B6q9hUPz4kzw0XgVpYQcC0BmH+
sz5MZ4HhErOO6RgwhKvgtlfc7DQ/n1xKGvGelE4pQ2sIReGGukBckmvfZYiaPqwn
0Wen/srNb+O08XpZkuWslcMqXkoggvnJKEEVJxCQYud/gNaUgEbCA5PXvzbwWKT8
GGHsWkeAPMkZ7FqJNz32HYyz4RxBA8R9eb7wu/6cPHqbeY9Yrp33OZ5mxzCnKHew
uElXBJpR3p+y+ZeYiPv4t8Dyv8BoZ52+tDHrECw4wnq4ipFiePZ91AWihIyPmVMP
tiGmt3etvE2dq5ZIv1I2fJyAMkQRgBopU27Gd2XqwBLnZCgsdwTUwZtbAemoGnTR
Wsj0EvTzmg0waElRbG/dU5v7UhOLdhEK2cX/kjT8mQCx4rYXSrvGxMBVQq+WjkVw
OkE27Sl/2dGJKeiDj9YLkDBsKcYMSaNGC7mPp21yuVXU94RF9fIltrUWNJz1+pTs
qTP77fTXqcXtUzq9uPWI/bRA+0lMpkbXD+9V/wWnIAqKuQctEypxzA8JgmUpJrLv
ImsMVerdHdAErylOEexuPfEtaVHiZxhT5B5287x34WSlMWo/szebymGAZ/Y09x2M
mM85SW807AAFQPkfBGiH7rBLsQS/3S1TpBs7ZZRVTrQRNvlPBsHg7X17BL57fhSj
S0VRkBglrNyoN0hkBmTiTIjSAjHm981+P6D4/r363Z6wq+9pUpKSPIUm4cL8SGGU
yUtML7ARRvECCSB8GS4MLNTenw+pkQPoOQ0QnW+nl5LCWAP7RSpbTMrN7VFL667K
2SlngkfGeWbO84XILxBd+EIAZ0NPCiCGT4qeOmyb/dawdTmJ8ZPfsjlReqwYuhjy
moKtFkRqvoYnDGIC/+QFOG8UQZ3B/TzO+2xxclsl+tBumqlgubrxSqoB9L3t6IyY
QLN2oTghiArsBp3GddmntZU8Hg/xv6TEPQHmha+krcfDnq380mWouUw6oEMJ0Kuv
89EhrgMhfBLsRSUph53AVpyrj+ZxwyvlqlO4gln2lAMWSPsiLyZih/0lnxg+uISk
01KCyAtGEL6SXjfxGyMLtOvrudgUVdeTItRnnJiByEp+SJ4EVqyU8wXpzo9FO2QI
xW0LOsXpd6CKEDGvbKb784um1qjw+1Z1esFQ9rVIX2E/KLh+fAkKe02Vjyl7kswQ
hQgJaDBQGz2l4fpMcOynE1cxF8fG9wDWbyR4CEwdrks1EKd+OflbRyC6EjcbiIFY
WnoBW84TuV66P0MVQ9j/NyH3X/Amd8BXhMs+vQP9ACytuFlMnOzLXbNkAuoPkJVR
zfOoUiQ3uO00n8XC4EbHCRjlSAWUVB0TjReaWTIgc3yjvRL6W3YJDEYnjkEwtMOQ
C2QBKwK2K4Euz/3nVHl9ZXttKHhDiif1kxJx2wfpI7l5SXDEr0uLahpn490oPc5e
PAadoYUWAAIyZ0fwSqvtMWlJB2pMJ0RMI4+hLe9ihRGAUTgyiTrH1C0/fks7DeHS
CgnGS7bJj64oG4vrKkJgAIUTfxD2qxHl0Lu8kU/JrIDslUKjm9kyrWQdaMo/mXZf
5g7jAatt+sOWBVRJPPRfEQuCicTsIcmQc9DfRoikLEMUJL05wZwE5SKbyXZUEjs9
kedG5A10yksQMgJ1AW3ZmuKruKAy7ulTsph7rb10gC8k9zpBQbLPZKpbgy8WIBe6
B6fz+7GRl3qedxOGgWaa2CC4AtIUvjhpk3DDTXSHY3lwdschbmkZoczZIqRST+UR
neObrs4uf00MVV8Eig/LQC1rX6J69CAUBEvZ48Y5Q/l/ylD/8yfrcR14ZqPA37B4
WQMzuamTu8aWpfV4GIUFRE9EITy6eeVh/bSd9pjgbQgCeJg2zkWOHKCLBKYtdowd
l+o1HdntZKz9m7j9Rt3ycmu367Vm382suditWwlR3vf3V4/i2xqnvYB+8zLFGuR8
WizZZFrKrQlyzyUIkBrC2KZfPkkw/Vmr+5xutmKjRvKvAZqfQSO1IYMlOBBKNG8+
Yz01ytGxQVsMst8J1Q2YHDRgmqCcjSxQUkXNA9DFg/jsVaSi9Y/LAfrpJHjxhV9b
Jjpfu7RC6lQ05MQ18Fp3XzdYnwc/Vxlm9a22sHQIfMyqOeP/9zkoFSoncyJDb5Qa
0sKLJi3RNAw8N19JKirU/9nuIjNy9diNkgVGz5LWZd5sV1kGrRHawBnwArX0TSoA
1CiDPKN+YREu9pk4T7yjVS8lm4Y8cg/upUhZz88lF2DT3YRlCxTYDV7XixWkBORb
TSXzVjpqzh7oeQxdYMLwPjJtZ2TDzonF85EwrDYWEyOvwt5ebo0qTO3AmOcUhuxb
VikjGG+6b6IWxgPmUrrazQcWWc8SbAbn842j3uddtRUK/lJfex7Jq4AT09dmYdK+
bo9B1ZYT6OZMVMLodTJxiDngByMsd1ro96tRT3NLKebPx2d4wMgcewM6gZPTJzPU
Pi1JAc/OdlaNBjaBftC96zBzEEcYyTwlbm3Gezj8sSbpShArcbCgiK4MOXxFhEz+
oeOIo0hUhK0INsGSbjB4sNpY5zjZ/KM7D3OmF10U6t8euaYQJC5CH9XCedt5haA3
+MiZLyU6tPRiteTcplXH4QeCxW7ObV2jCh4A8l13odNLAYSYc2r+EhPH9x6bKhgO
59dwhvJZiUL53iY8/f9QcvMPGAW4ZnRMFsoXLDJDrm8yOTnAxpSND+L2SoT2NcfE
VhCge8AY3LYbdDwu6tVo23hxv1FpxHHY5WqXqp76hhpG/SQ4F3erK9xjI1KgB2Dg
6j3u+IYSz+C9ZSNlQkjI5+3n7QIsNXFGuQdjnI5LeoGIXj5Bia2K8Ai8YWPflbkH
NgzmXAXghyGcAjLV5L5CIkFEXxEvHmKDLE0Z4NWglLdNEyD0O5qOJZo/XCEwl52U
QuRrxzS6DhtLap6B4zW8bY1DhbWGMqbyQiPWBG1a7ezbZoSef2jrI4ffR6feeEmF
162AK4HaO0xNRQlmPZa7HtqmEb+MtVpRGimG83GxGaGgyG4zjHhqkmUOHzxL00rC
d2aGzvN2440k09KeRbwsupqcgWXsNRE9qA5EBsGS4O0ZgQr6w3qD7EvzZRe0EQLn
oMj+kPP1W27Fuc2WadMNyFLKxaqVI2LnRDqvLfjr9hBRlOrj6Pl/IHJV+taHIIxf
ewn+6w8jE0JHemzYTiaKd4oQToW+kq3aVoAPfyj+8fDvaOiOGtaQYJ+vuPl5mt5T
Wwj/xeFwcVapPXetLWBSFMGdvfaEJWD4hU5hsKC+HKv5KxUpO4q/W3uJYtg2uNx1
4dwQ3QMmrUr2eRrYh/hTC3rFQr2++MNQi0fSWOQ2lMu0iQI0xlfby5YbRaye+caD
vmjclTK+7xyzpAlCRerCaENigOCLnQfgstaMw4hAsY/XS8RbYtm0wrmiN3NrdQ1P
CRq//yGeMPWQnaMSekZ2YvX+L9pz7OujkFzDnvwvKqwCrzIGNUSfoLQ8F3SY0zRR
73FpvcnUZ5FALSeggdcFqNPNVTcOSqcm3Lk1kFrpdpOpz+3a5Zmp89pyTpTUfJZA
8ekfEvH8LxHidrzbfCnccUSAVJHmtMIUMU+ATSlD0Kv9pjmt7MXktDzQn7Hr9nlF
VXavoqVVrLXOpNOVCTTr53LeUPjE715OZIOj/kMpQ4FFvwuBuu0YmVmZBYSLCJFW
9WMJrJOMAXSPnTn1Pjo79m9BGIQcxhhxlCpNqnuyCF1WB18yVoef3CJ3VjixPUqL
6KTE+yXfJhV1UWOKIBWGXzKTxyvSHSwjCZZouwzhvil2adlQAzPV23gXWXnrUOjA
PSYYKIlW1M4A0Nf3YQuElvsPLdFLlz0tZwT3od714+BqMNWje+lq+MRVPATlvktI
SrtB8z9kCQKoBSNPGYaMfvDh3svRykHYsaBeevuiZhw+1bmLbaNxfsFqHOAhSZW/
zD4hy93+dBcFi360LttCZiuKsaXXjcjyttJ7HUgj2oG4byW3ZXSNOr/IlwEEbMC4
IGTgG0oyiHTK+rH2rlEYTPc32f7hbANNnko+IvIttygvZIh6SGfGoxWJmbvUDDCN
5rfR2AU5a8mxmaRUPIu5T1w4fNLh4WYGIHe0p37mPFoMH7hvnCdNEBtplSvBVH+2
74/J+6ZmEYpF3K0pIOxO7ak2myTZYyXQx1iElwNnFUhErQYOLCzcDoQXPCJ6QiFx
u4ir2TyiIs7BG8cEwZyevue13ZgNbAlTEz+Ct8bUSWqrER7LYvr0sHQZBWeoVh7k
oS1S24Xg7cLaERhwCfDuJMJiDQHAJ7h+yzhxNIxwOElwmYAUG3B6DCJvzwS89YLu
+7e9kd3mDYGTYRLmFIAOzCRbdK2iKaGXwjsHVbkMypr37e1biqG+Y+uqHMaqJ23k
jAKXyDthJ2iWc822JFZWciMsJUIA4ku3GMDMMLQnRXE+MtyGZFftqeaLHO7g2uCp
timO1Zjd65b4bUQW9cuKMGFhqqS3we67hZNIrfl/mX1iLN4sNxf9bB4hIUHKURrN
sPBBVpOcZAtA0y828e+z+zN3fF9EvDF4+9nQFBDhv3ooxU+ZWC8p28v8+mBMcBEf
/iIe3ERK8SwGN47+q/d9iak9zzTIF33F9g/Ty3cAI4O85ePNJexPt1TsjPkGHyRc
db7vEcgUWtjxAXvS4cv5MB2vvredS2KBYNYnEwa6GlsG4MBT6aiyp9bGoTFPdPT6
K11t6TxbYxqJcbOvWt3CNwvwc/dfalo9F3faRD2Qxdrq7d4mNKnQhOyzAFg8w6qC
umn7AhJkejIXV0qx5srnUx+D1QcZjQJpwi6jHK6XE8C5DDPc/pV3u0K9lE/mSxEW
CX18qNRzK5PCAiAsvtoYPnTSzpxwlTwnvpaEFJzfZeXnTXfTBMdY7258Af/k1elg
KdCbo89rT72CVNE7aWsGUrZdUDSJpt8BFaXfJd0tPrjGq0ukm516AMfEzARUNB30
t8BrEcTKYfLFjrOnMgDVlCtyZfJSxOAMa1G2s6tZeRVzbOwYaw9OlVPz68Gww+yp
w79K+XZo2B6JazNS2XghfuT7uHcoPr/W21cyMpoEu5zprzskFjdIm55MOTt+oqGG
z0ukP5HOxX5AfMVVVoW4HolzWLX6V6TQ6B4SAJNhXq4ahOywUMRM6ghSqKBpT+6f
RC/ZA54YKxoZiw7FF1GauTE9nD+EhoD+QV4fCbvc4av2uGtJnv4XSZ+11q71vu5g
CwKtE4czXG1gsDls3pyd2GWSs25fGuVvKIYt/ro7NPfHUR7lZIqvBd0oh2itrJhv
J4RUukVIM6hfg54V0p/E/reJa8N9Utrcj6iLx1gzHzb3Petk3+1w/I1Q5aCasikL
iP74cdeQSc5EfyhpBkuzorJ/NQmru2Ryrr+7mjXMRt0eqmnQxfbQ4Z9gWdFqe19C
Stq1v4quYB96fXstDIsQ3XMswNXXxbVy9QEKuiNII5jeJ7N2HbsKPt7Q1dTPtjDD
Cy6mrF8y77iuywBlpTAPpQrfW0bb+kROVqt+EKD8cwndKikl9ZqnESDWiCMqtgnx
T37hxpQgPkfTigMMiupKcgogpVYwvOxKXvJ2ivaA8NqIJMEQhc8aDF5MmEspRG9r
FJiePsPaCdxnNoTlBE+LHgK2sbbFBnxHqBg/sVtjgsjnq+c4XEtVZXLBmv/4Z9mO
YcZpBW2bzZmgmy/Bhy92wD/Je5kv3wyzACa8nps2MYCZx1Z3EtnOJrSEy14wfT4n
pI5BaAA5AkfX/3T9aawFe8Dwze28kh44g9MKwfU4aAGqnxNMhUl1H71SYiDGEBj3
PMSjMH7IH1MSAa+w8NB04H/gVQvVGoDJM0mrccyAdVlZRYi3oenzhIzYKF3QRo19
T77u8XwdnY+efzS7+HAj8K0yUVmI1zuPhxq58XNWUNfUpjLv38hO8ujRKJFyVkKp
27muY3VXrzUDSdRpClJRIKa0fvw+SRBQYNis0JFYjElbEqyEmtmo7gzPtGWsWWTQ
HevFSpYbWK/fs+Lr3OzJHDmnaf/f55rEItnGg2VyQkdKbuieHHq3KiwqP/cZkfVA
axQJ4F6ehGBecfz3S3lF+1gmAMIwiR3jGttWrbediEAqyP51Bzp5SfcJOe6FkBJi
VOzeSk0vwSFfKSaveiIg8wD+ejjbGSr4iv//kBuiA45rguJypFxiuqOWhPWfYAEU
1RRdCD04tfcf8a6QzIRKAToYziUtp+eF6ZkjKePQ9tsMD1oinN5exeKZPOzzG0w1
CHlM5VARxG3LiH5yz1QNPQKw1MC/CbdFye17dwpFL/2kFNOFh+VWtylYE4MOBGwA
GPD9AgYtokR6Ki+/H5hQ0E7pRgV/MTKtk+rAdJymDE8Llr2E2J0P5ChuDS9FR5Yx
PgZgvZlKbMOddmfxw6nUb6x6UOfS+RQcnVJYDBfnalKBAT79T+S0perRU3pYgUFv
sj/vl8rSfPfeHz6zA0V633OdRCZgJHtoRmO0/pqEF5OKwF+mlzsgNJehmQQK4DaR
dFJqWFM/2dK/Fc50fTWiubcdFhQCL6ysZ6lf9oNZMptmMeOadZFp17KTa6QlyXlu
bl+hiQ6TxI4oYf4UeBIMwCQdUz5mCVUs9C/dGa9vVwL2crvbw35ydwM7Htf4BoH9
YIijNkrUS029idIrqdKTO5v3uiZNrPLBGqH3Tv5EiVZHttUq9p439Udbx6PEJ79P
RU8HX1xzHNsikZUQeMG+a8z4aVAta1t15EioC4Lp8D3aVeBNOoPHVjodgitzR8Re
vMrI/vFGGmJwbk0IRqOxzRuAj5xOqwz7WZCCRKlhbB78Dmb/vTXZQPPoc1na0rkp
34laXCMr9Qp9YMrnoKfZBcXrQ1PSxfHTS9Y5d5eRSkS973eTIAZhafJ+qHBwukel
I7rkLJNrsHGM04q7r+4BUSaZeCwG8u4TnE2hChNLM6bB+H8nxRYkk4RSG29xKZC4
Y3MhSEi4hBmZfen1FB43LsySb4LN9KaaAIlV0+haxNBF4sI1cw/BGfDt0NTCpmsg
MShSJ+mpbvaEMbFJdx4/7AhTAC2Z4iNVHS0FBiYx6kfZomabqC8DBYGEr8Jr+Oc/
M7mXeqznRArY1/S4Zkwja/jlkFh4N1BFAspgg5sPzFhaO77oiRtvzsyNYnOCmL3F
qzWvm7MSXfX1vsSnqpLL4waLz7cxnwxUSJOtVxmjylOM/ALKzZ1208u5ujrz8wUi
8b8krzDXTRP+bTYQFLDfWEmlAcoJUnnSxtf/Pya+KW28agcbUK4obrWwOCPp+6dC
w1rrPkoa+v0PcEx/x+xp75WQti1ewM4RQxJAewcQmZdsk0Yn+qOkhitiRrglHVCj
DbuLbzoXwMQSJAAXX1Ty5d/Hg7hbOsErnQdk9OmKHrRYfyeAS5xgv+moLkyB4Q92
aa85MPmZHDlHbbxvY56irm1aQRNNTomItk4f1ODzkQWPDyeorIy4zjKE0yzJsK5v
wuPy0GE3w9t3tpo2G5h4QDK06yrh8bj1Ywqq5OBnhtkvUsO/twDAMWgCsYXmetbW
fAlXFZ7b46mcFmMtjnL1pV4e5Z4GRyBCFcumscMrSoSR+MXzlB0JpaUqU1PJdrYK
3Lj3dGQd7YN9FucXvCSQkext5TCjyRdaatS4QIsbaD06axaCGnWJA9sfWEfk762B
TZMwyfXcJYpFtgH4QK37pVVkZMJVtHGO7L1T86kihZoRScoHBDT0xjS//h2oof5H
GoJZ7Eq71PeXWDyFxN3maRO0xU2A/0gthOFo5yJk0oKGM+iGcPMhA/O4rghkox8C
RXDfUvcODLlzDVdekPHkN+GI143QEqUkufiHqvDDQ0LSuf8awRPYgu78HYxvkgm+
7aCDn+stgP4OunB7hgoFbl8YYWMyMqZyW5G/FNrHqxu7PFgCjjc5m22QIEnsnb76
Is6POA4xXStehSUmY+/HDJrIiP6SeD6u6Z+Yr+VboObmKbNZ6eAeafRsM9sFk2oj
Z1S8Og3TxQzVPLjrX7QnvFGp08vkPLZsX1jBYAE38cK7f3p1qJxBJZhW1gkJ8xUC
GNXpqJ3ec8YVW5rujwMjfFlKlJJNVgS/hDAk6TaOwcM594ANyBdCtCzMgr4eL/1o
EVu277kVeEXrOCkRNdR4zP50uS2r3H7FUHp4eCNuRCRDsAwsb/G36I0qze6JYptI
Mztc6mYgUbTIMf7rYaolSBKzJ4q8L6poCiVPXNORPvSAGn+FKndxlLkKqkipFqtG
L04mEBlWEP5u+AGGKOE50riP3EK7KhoeTokRrEzE7iZk7MhguAQy62t9qAehXRd1
ghSkekUjTxzRL0X/cjNZG/2QNVmMMqZjMA9u1Smg6KvzGgDwjU5pyYyrc0atMdZV
f8Q6+I1uku0aA3HK13hEOB2KRTBxpjUYKQjDyVIni5YPGZwse5ISRQTAmS6rRbor
bk8TWHZ4zBpPCk8FDswsULSd04/gckZNki3MeqX2DZ2EZxvJaejjSCcVQNP0hX/c
dr3Cj36gmRjoXcQyHsnAR0FraHKq9ns09xNJdD7M2ELEDqQwwvL+4EaIRmONklQZ
6o19epdaBnrmRNaHKxE6FiN5Nv0nzLvXKDgNIvPWJmla9WZcGNZXJD6T/FupxoHZ
OS8X2apSbTjVOKOcL/DxNqlMkf36jR/JmXSSW5D2Najd53f9oM10yEYs2ASNhzrJ
MNnabfOxqupQts16ekMJbwq+M5rGWvgvG5e8bZs19QlcUkxLKZa1QXb4x5NUwapU
/Ut+UO9nVA5XUQF7Cc8Q+ClCEX/jDPoqxmKLwtZ7a5kHFAYrByfumxinGUzvG/1q
gIUN9k+YRVjDS5qNS7fs+djjaoywH6Q2nXW8lIEO2yNY5h7C2Bf6qUMBV30HHOLX
pjTGiWnBE7BqjrdRCi9sHJnCVf4shyeCE1oIl3yIjos01SDUn0nxO/3wAssANQ1U
t+kN/wdHrOp3ZdGTaJNj7veeoJKAAMMKShT0LdgsBSR9Ij3eI64M1Q3A94NPmy+L
WQ7/mVgUTzVXjDhdxsdn0bEFC0Jge46CUoAOxgEGoSomKMz/qflkHgWxFGNGU+qD
omQ3QEaVNrSLwFk0HnM5G3wa6Aa5mFoYcjd97XUd8hYF1VwO0FboH9oBq8/qcOUd
a0txjQMuVF2ChQWQ5tztk47UrFMHx5dLnyfulT2wAeoWEgjSgnoiAhzDp/4yPxCz
CwKViTG1zc4VC8q8dD4pfqgYuiqFgKgZfEAZq6vnCVtE0wsuYJN6Spp5zFioaC/L
AdXZwb8Qww71xLdC/Y8BM5EtSPB/Ay7hBPFrG6/pUOvPhnhhGGqItX9XIMghpfQZ
pOV6/w6iPcGG9WcOCceSO7gRG3vva7NQ2sYeNZMp/RxgAIsxxETaiqnc3HRKTVHg
Ahz1qbj9a73gvlNM3W5gorUMXg1ky1Ln16yoaZifY1rNz9HazYNW1VB6DOLsGxLM
xwr9w+xMyU1+ln/mfGs8uWELpz1JaWo9Yb6IK5vjBDc0U4vwr4P5bZfSMKCL/hm4
1O6H5ln4uVETQ88R5xdZHKQIZlcoBjTR4yPrShTs+BrSbKdmAhnZU4r8zPLrWpRw
Q5JebnBjDj7ce16IrBgPdsZ21r6AsalilN92mKT+IEdjIB+wYxEhKz5C9FWJc/BR
a4fSyymiVVS4QNIvYEzxhU/rhVg51I1975vZqtopqMmuZp18BElER5ZlpooVxk3O
T2/ALL19sa+nmbTvuTFQUZIHM5CCZm+zZkWVudCRIHxvbcXYiYk4PQGr/amThQq0
S7q2KLu5gU/loCay2tZiKy9AT1KVdyfE92UcIdu9n30uogCKAgXQob/S/EEClFsn
PbaVQ/MhjA2hjPNP8hvYBh5tNhpY+cykEMY5MBMXmzS/zk4agGG8VeC74tlya2CT
piEhWOhzg5X/szG6DolE/pb85QuIPti/GOJvopF0onTRAwAULXHn1R67z1bhM3ai
1876E/yk6wStdfP4GMk2W3lSuCOvQb6M9Wpim/CrrVu4CV3mQtNTwjO+fvkTWARB
JrCRmDO72D/r6pi76QBVxROJfH/CAFlcghqiaUYLOqkmeABIGfA79ic7OVxwVxus
C3tzHMACrpWPjSd9M21gkeiib+N4P4xngLESghgjesdpqsfMbB1x5Hj6Y+T2WS/T
LEPrvJmBeAUyu4fzS83k+tHqlLr6ONPU/a3XODt9dxW9fIvdzi3J03uVZ7OZ3z8s
LX2F7WmcsLBxJhFj55dHn5cJ8si8CcPNXRa+oKc4CuWCUJ7DOhpqiwmcjSw05xX9
R5j6yfUvOEhQPf95t/VWaiDJz95hykaJTZxBqwuxEmPVzpHI/i2TPpAapUgH9g7R
GKdN2l/yrsmDSM8Zrb7HzWt7PUH9BLQDEL64I0k/NVGVHduFlkF7qxiChkGMLrpR
WRqRyojvO9EWLJkvUv/RlDrqmJVAkzldrsXI5B03yznud0KnNDjNhne0ptefrgCC
HFEPiBtJKJSXojyd0rSSwdhTR8Rtvs5/6ISsywm7YonP5fryXxBCtHzkmqGWpQMN
Xwd9RGswRpXIvrpvS6hhmIbxsc9lvz0gVfyFjk97ahLshzakHTtopAvPbrHzWC9F
R92aRIk6CDkN0Scy9oEPYncHAASdVtEEzwPc1AbX9M8LkukZkxlnjIgd65nC+UbD
PQH9rYxEn5gATFsACF0EBMVrb6oUkXbW0rJOoAKSbRkKA0yvp3ElYV9vvk/b6tOS
qZMDd2dFZXW/kOmQgSGUvmhdNP1gOaiB9mkzYsYBZjaKcOcFvLpn5pY0f1Fl8ied
GiUVaGYDT2kaaSx8JN6N7tnDX1EXVKfHXaws943lYYBLJHnstD7ScrnB520oXVa6
PLNvUh6+a6s5AqGViuITTgjhnLXT6vsPPcH9bddwmUf2wi1oiojpgczo4kK6e0d/
VY2w95nrrKSUVJM5TGWKb44625zQ4ioTNQq5CVSiLbRpGojXr6ezFVtUcOsju/sn
IR+7yDUuRnct5i5Qo2Jivy9BL/ZH4ynasm8xiRTyFsaD2zoQe2lwyuMAHTfGV+oj
Um6GQXF5BZgRWQpXe9Nm1/aIRdhyzpoe7d+pXk5BN5LvujghNsIjvniUbCfYTT6q
n8uCrNqrHmJr/FaYjBrVZOnnrf2GyaPZ9BkJVLvPUdvGEQdo/QueKgfWMlUg6+/1
7so8zOwy5VY298KNW630bXVQvG2paqobiZdTR2RVEBtOMrHXDWMsgpooR5+/ri43
P/zn+2xqFpxRnqjTWmkCOpIqhd7P+AeJLa7ACRXT3DxVCt70idwKn35mHBvtWd7I
tHRZgNXVfqcdBJb+PZL6dSGPoJnvQFaBgpgGu8ZQy2ImjpnNwxhFnkLS137RujwY
x00vZ76Ntj1Y57BDD3nUQ1Dtnm44N8aQQ05DdL4nVkHoLeyU9iDpeaa0d4CHdo6o
kZ8B9qvc7HSk0nPt7xu61j9sipVR2//QI1XzsTmR3e9Fkn9TRFfOJwM0onu7TZAM
3EOGWOh8hpfkp7hNaeRLJAvf0BC9YniLiVZWdg3soxu+r8cjtJ+sW3R9wXqGr8He
WYOfbNwdpmpx0snG4keu+NTnvc3VUIA8OvLHxP2sQGW49HofUUfTkfT/yNgJaTBZ
qUpTkn6rvEa3O0QFn5uPfroLvrHru2rXKb2DatG0innQSX76XXbPs0VKchZntxSK
tw62wKb9EQxiJwCOpzhvHRzDcjL8x9aTxhHiixua1R6eIlz7SpSrZWfdg2O1avIu
IsgBQW15BHiqt89tvc+njzUwJeP7MkzxOr6nWOnqvn3/2gbDMTRAlTa065bWoCjB
GNMR9LwB65YZsGOZfXqc6V7uFaAIlshV2OFWgamQSnouh3ug4pH0mZmEARWgKoVg
DdsdqUegazsVjA6w82wEc6CyCWvbTTWeoiciiwoRqn9Xtc3UlAmU4Nqgb3xYktSZ
dPG9OQ/AsT4kG2OB60uj+r8KqWf1Cshb69ZiFVgELzvQOiJIOqT2zgbWvHzOiDPO
NdroOiEC07LqRzJRC3L3JsERq8dvK1/O6Cb4FsnKE9auwSS/7dyEEssy9J4jcOgb
n4dQmoD0MQOON4WFmmCrvymJOP4ww+P7ajkU4pFEgmwm6yxxukbAt9hEpQJ28oid
wnI58zzinI8+wOUrlkBGwWI/oMskHWf6pcA2/13qegtHXGuNCpYPFgDv6FPJzpmG
C0z5yLi1M9KtqFUpVMuP7GRz+QMYotSphEJvERz+KhxYjISz7dV5mhSfKIIJjGiV
E79VQuLO1u5+9GvT9Hz/T8iF76+AJZ4XAkJ725ynZWWJ3hsd7rZSkJks47XXXiyb
IE2QQuNfuXCzHN4f1kehGQm08dPaK6BQj5KmMBwSmJkpeMEGaOqb0SaqKowdfAxo
UOCcVAeK3bVCvhN6RSzuho6h735on9wutfp9+ROwbBX93KOOc/dN/OnwJc6wCcOh
6T/1LHbopCwGc8ppsLhKwPKzafjLTG0O+k4agnDRS5Qh7XiZF0xlXJFaQ3xPXCX4
YZgjhfTEM9ShRg9d7JMroCBCFHyoM8yyEZS5VEFxPb5F6c3jVxaP+z4X++vGB7AH
sQxth3RklFAjKZq5VVhgumkEAYfz4O0lrWoXaz7/upM7Pd0PfnQMEBCJ9udHXamZ
Oo1brcsAap9hEsn8rEE1ozWuj95oFfZMNGYpTPyL98bQRgxps1dAq30+hvj2skC7
DDVZjmR9lo3UpsTLBtXiJSGMx4e9ODCKmrj8yeqZx1MCZhP2Zg03P4Xvr/cSxeVR
zkY5GfCDhzu/yhJr9vhQYG6/8PoTTVeyTHoZm8cGVVVeV6fkyxlDFqDnLMpg5iHf
lZ+8wtEzq0cQ/06muD9Y7T0/66xOzy7q77YX9jsZrUaCAZagT7hHJihmZJlkeiGz
16RZ4j41C4JS6GJg0CEj4hYpyDHIF4HVnMDbYxyBdMap7gSc0Wd9Nsn5tn8iM2rO
mE5+Qpw03ACEORyukBtE0mRAytMopdSK8CzCBs4s0aI4C9gEj+jEb154ViFgZctY
vI3W6DVmhubB1sbNJ7mSS/ODThXmVneDl5XXr39c6PiZJAm2Ik1AcBKdjsM1hIn9
R1BhqdW0PMSNzUqPPsBZN0hvZdVHYSKLb975IkajfRhBDtdD8FWvn76SuLOzTjmp
oM35af+jYGqQ8SNEf1zrvLMoRiGchfKP3TBzCvvuWtSGnRByIJ6emnDC2tL/GaeG
bsRde4dd0L4mf8E9ccir/P1gkwyLJlHYCdVOr3J1YWDd6jCks3dk8/6HDi6Dn2AM
wh0tRfTcXbPSaN/Q+ulQwezx6RN746Yl5NV8zfCpGZt2MqrI2JsZi2y4hUIfkJ6x
7c/FB5lJiRav+y3DpG6JUf/wL/tJPd+41Gh4VodEVM3fr7YHwHjlwYnHYZU0ztug
8O3ym/6cFrZHsoiO2kNMhrHm0QpkL7iodkt3be5jn6T853sVsXFzbQnLlWCIRIbl
5n8FnXXKJN5iKbW9FvvlLvytDa94WF1mH/cgvX6q8aY/XTFGNU8foh/gBy7RoPjm
Msqyh7+++M1SIi0I9IQOey3UvPDO2SPlMvwN/p9U9/OsRQ6pe7EtkIJw0+y7ddoA
hp03o2JFimhodUOM/7R2i5XZyqfdbZS+AdrqQR/0W8Abiv7Y5gyrTWGzboa5A1hO
qqC4s+8q9lXXAD0ghnIAHs6nG2GZPiFoH4A7QyxL9R1dfBCAa0AoFOByen9AwKiC
0ecnXa30IsllUHbs/K8dJf0acGZoCYiuP+amGbVpNn04a+VLg5hSRtxwtHXSXX0A
0adDs5hBmQJob3lQ2KdyEACb+y+fouTuerNFjbzoeQ/HEmMzKv+QWaOLv5u9HmyN
v+Nk4DBbKXQ25Hm6BQABsJ/i5Y8qRa0Z1NEO0VbX2jFr/MiRUN/+4eSKAYElUVHt
InJvC+VODqRHIf9l4hC+S39ar2qf3RrTI1G87VBjSVeHMgOjQ9RQ5+nH0hC23X3O
DEByvq410AV6gxMp7LvsYcNsyCGoeI1oVjITaMS2b9uzNYmyqub7gZODnoWKA8y4
0E9Nz5xfE5djvsQKtkNDOASriK+aISQr/ElBC0jCy0RkT19otRKGhg1GsjRiyTKq
9JQ0lC4CkWQL5qFOP6D59Lxd6n/Hq5YEU8CP488mEbeTriWeGvXqpw5oY3388mlA
zrVo0ycdRmYonMiCom8ghSdIsZdDvrePFiSvCpgyO/8fcZszaLv1g7KAkd0h55qp
pDTkSTigwsqCEz49YCEFAoCIj8CIjeg/ZgVKNf3Iih5Uqvfp0LgffNfGcLOSepMr
pWGTI6+ls6V2Ffh+xO6snFfdCyIAHW63CEg2/fOWT5gBQjE0vea7AK/ESXlZesBW
9z64ykft0jisnnVVHTJxL9n3vD4ZTury8zPAkT9RXNy5604BbX8c+cYfw5kPQF7k
Ti09UOdOHXbn4wwSOzv9Tx/eiHq1hbvkH9OGJPfm8SY1RlP/T7LfTeiGPfGeuO5z
TsL2fqoy4qUo01vcIXTN+YNVxfBwCq01HFyfsQolUe9WsVYe1mEb3h22P3/jBcFV
dpxvQXYqdxiHn3IhcLVl3y8XKqQmHEMG4ZDBlgnE2pmuLk/8d+NMaX1uQuJ1ZMdH
igggakRiUUUVuf686c+imryCjn/4r5X8s8U9uCXkjQcvrQyFIYklng9wXp6/nQzS
lAvQ472C96HGAAxZA3awv/2gb8B/Unt+MM7ELwNCqviIM5MIuKD/XeFwebqIebs4
+DuB/IzIgCUtdN9HAsvwoK6xA+VhlbkOdwHdQjYTCvrPCRODvr0ffx/DkG8FsMyg
qEgWNu8gH5K6040IdPhC/TwS6fXVSG/fXJip+HzsLeM6ZunA2vJEEWSR6KQCpmFC
+Pw1gffyqhRZV0IHusyLKKpmnunhLz8qVie+Hp119KclPqHaLyqfOMl2J6CWnYOX
+C2GIMsFEm48qVC7IH9S97ursirvj+PkAdR+N7NPbDs6OU9kP7kSkV5mKBpFO7nt
SG+9vX6/y/zLy5RslnW4vjackjDVCsFJK2C3CTahmdv2d5aKk1Dzhddf3ppw054P
Fb5tBr3M2vmlHUpOc7toXt+GTTEmYo0kds27pprO2j4fICOvghkRz/dKIHEhRg6+
WpdOWoS3OW+5nRnFiwjuJWZEKHnMRJOeXN/RQf8Iy0gFIoOHhSgDiJtOyXNmFS4E
RkjGozBwpjLRhxbtYU/oE+N3fSB5KU0rO0kGKDePw7qG2ips22mP5EuPV8ZgqWui
kBWX/vL7AmgXAy2yHsUlRIKxmE/53TIWNSLsv9aeudNmLaXYbdB4cqQvAddDMbzP
NqRjhxI8uZFXUzXWyu2DZVZRyUliOwZ7lzrfrAfOfWDGstlVhjvIgeOQyABM1NFU
Z1/B+yoPPwf75J96YsZAOzDIvMjwUTGc9Pp/szsqA2mb778JmE5O1WjwPGdYB8kr
YhxMzV3yYLmgObq1yT22WQdKYsJuLmkbukfBm0m0WN44GbMHc3EanD5vMhsjRZfe
tLqnVxPpd+OxwWK5mX0+B+kTTWbNOZUErgI1LbiFb5+mipW+TsZMIWM8g956sPg+
IQryz9ZsBUyfbyh5JYOxSXE7PjS3FMwiHypQUCsWybdVBTjgUp+xpJFAh6i11g5I
lW4wnkk01tUL1IMK5jN8MuZ42cuM+l5i7XTd8bMdcASOJhp1IqoywbXnq8FsrMpc
Tfb0XnD+UCPfbo9nTIHMx3Zrgy/E7R+sM9xcw9HhwXfdPCZkn1OusNU6/ZBcx84X
0eMbDc9DGFZ6Zfojc00nPb19FMk2UYtczZGnrKlAKEIBOax02ADqjX/XngW7rI0i
q6KxrF4rJy6IlgYvCCvzZQ/2tTg2j+bTw9/cuvB72079GHnaSx/K8HTKUe09vhht
6AZdEjICFUIlwvpFtez4m42bBNghkNd1+U2WhNmDBqmPBxgB8yk1QWW9NP8qx6Ld
FVJAgQ1AvfqsUGuugob1E9h6/XWoHHnnRu/fH2Bhh1szBdGjBpVP+JPW4KBpja1R
ScoeCkatVQR4/UtBLFMyLqOjXeDmhHJIh8Ro9LyIoDcUXxr+uPr8FcwFKUneH+Gr
wREca8ZHTVqK24fAxupS5/jHxhjOUDWKUNhpEk6usJlxgJC5iWzKQniMtrTdfaQ2
LES5+qKHrPs3u0wdmMikIgeJBQfboLfpRB3swE3AL3gQMK2eGB40Q4x8kATyOedl
98amzeQsr0eDGr8aZm6c58zAVHAZQEwwduZICoN+x4cCqzUnE5TtylNmLUrFXBd8
xfU+dnNiru3K4llrY6ccKmYimDdlBgquk3kxDUJ0FdFVQGeMn6oaCc3ssBiXbeUK
d9+iy+Rk9O/WX1+yofSTcFljVm4XYJi/ELjAgu8j9araDhNPuyVCXa/rkLTeVuLp
jODiKDbMd3VJUOi0gKE4yrqu8avBPL6j8yNq8S2yGs1K5eLNYaw5ONPHg+Bkpyzl
yLpWzkSSjRii5aBFFmnleN6JSs7yy/bVWiUXAXfaPiupZRr5vSBynu/JwFvdM0oy
DFvkeNAef3NDpk5EYIm6liUQrDF8tW/Zz4lSlWJcJi8h9BxYt/pdQcKzUcve/rUr
+GwsBWuB51H8XCN9Ona+IPbhNl+xxRaPW+pkBFziI9d58lpObqB2a01roPt0kaXc
QKvk2uZuT28RBkvuvXxqGoP45SKKT3tgKTcr5sdInEMqRP/jcCIKkhYGTnjN8vrn
YaqPC1ZIERqsj0RGbpZ438lPuKZf3PpoeMDQQgozQOlKf4r4Iq92fRGul8/VA0zF
3K/THxjPdWhczgDsKWCcCw0rGGTLBVFPWnpaO8oaH+QRrPL/iHoP3dlNfuTjXO5A
CwiE6B6ott+g6Bgg5Zaf4AUCBpCwtDA9Z2Fjtrmja3tSzjO+dKquP6koWXdYvL27
+xQdwGuc13HbkIBAnJPqIGPnKb1gZ1rs88EWGDhKCeD/bIwN9l040nO48oUcPJUM
Yyb+2+ky2FUTmpdP83FFFaXXZT4sMeUVJ4iR6mBcfI2oP99Fo+CluwBLSZYeb45W
a+AK2YSpdxN5tUaUMz+gnk/HSmwq3985OnQtZ/W4gzhbunqGv056XTYiPQ1trqXz
P/E2VWlGL7A2fHKBuCRfhB0nRd3+oKX3a5m4LEVwDI7mji+N1RZtKUTtTlakmQGH
OP6mfYU3xpyLdpU6EnkrAey7APy1CkIvbrujr3PYWSFaKjAEFg0iidD1ofruIvPc
SfQ4w9DLnivtFq4AbEZRF/+JwOD/+35R3H4QEiNWyCT7wEhTg+Fl/3r6PGSmh3Iz
oWwFZA6sJszvCqfOWT+J23aCJatSfOcEYWY+WteDNQYX2SBpGmzSOiWRPP9atAHf
1CK6TzdKFX1qGIkWD1TwG6z3/6dIn4UVXo8QB+vaNAAdROsGKzcKJpqJCl10RAPc
X3Z4gOZpWhfpzZzyQ07Qq2cTx9809pYW5A3Jx4pRHyDFd+xxUbXI6SMAyP8supnu
bUSFQ1kS1IQYo4rwYAB6SwzxgJH3aIOX921sulJmIpZbECehaIfDTAC8UXq5MQMk
qYUhjyUXR/DRIaRDycI5aMrNPHFNpxEre69zDa/2hd1e9guBfCFsW+/V0OY9aX3g
GBj/Wge2iEWvJ7pxnSJb8wjMkZDAYeWkNSsiLfgqa0k94B2V5q8TSMoqZjRY9iXs
qNTOh/bBStSyhoWfn7KWn76FG/MRpCqExw8jyLpQRVy8hrji5RVNR7H/SWSTcCS9
6mTmBd8hR2YrUrZ6A9W5gT0m3i6mukF3cvi5/+gULhEWmfefR1BWGf9dsCByHhps
OAcA3ljgzVDUVm6prrIuPNtbnP9io3rEwLrOKGfFtqV8sZGOTtYnsrgDuCoV+D9E
zTwIZkwDH3nm1vodDLdGFuaJyfjPN12plMH6v31Q8b4SHR2D2WX+JAPeYMCQ8/7d
xdaT+wNfZ0K2UoPtw75VFgAYjwEBtC4XCgQM39oCTnHjIAM4u5UCq8J3pUbc+Pea
i9Ksw4l6HZc/Hyv6P9Ut5qPrd1MPozdU8fk9BlCv7NllXzLT6wB5W0VIaNRDJrOV
Fcx4L7IZkFmpkklbMHYsy5159omrDEa/z0bGvS8GRVfv6mXf3oMQxA0xM/5tve6n
yZX/Yy6rYnvQxctIQsnTHpFe9O1nUvxTXxckKZwH9002t4eZOgRd8enA7H90H42Y
bTbhu4Kn1p2v0/lGlKtDdpvklKcshYjWAzIcYC2Y7ZhtqNiQwZhw2VghgDrVpQP9
u6QE3Gypr+pb9Ie8LsFIoMDvtq1NG6QHwayNF9Mreq5M+bblxh21M2b5QnTPr1JW
FhYQQf+rOVz8OyfvgqTwrE7iaNEbw/j55WyaODC3QzkpRFojtKglkoQheD4fGMBq
kJ8MbQ1KwrwCdD/sg9ezGvMA5/TMILi6/nCJqqTteBLoN1767WoUMBhHwjdoBm+N
PhN3eKGIz8wjKkyFDpGCYRbLF4AL52/H1mmLzXDLshmBARr+6eg6MAJ1iVFY5EVu
WRZtsBlxsMhPHD3JVjNY9Mq0DrNeDtMTL2wXudGAV+MiOild0+12nMNs+ZduEupV
bFkMMS5MFtrD90uXXUB/MZTDpdAZSxtB8me1OeuegXVeQB3dlMxeulpb8bLX7WSs
dc0qYdfSGa9AeBiGJi/Gfe/EYWQDDx+5UD6Q0EJotLOBHuZWnn51zx36K3UpW9e8
LN4EqMqO+tGyJV+Y3xNd+iVtUT/o9QfduWcAXLs5pTwi0LenScPM9EjMmYCnjCQu
nFkIDahpKfkkdKWVa5vmREiDeagONEGm1q1ieoAoboD0+9FQvQCJuo/bRV7gApfy
nwFLYFBJa1AS3PWutdmiIqBeZFpwBlYWiuLXW5VU1KPhLTJfnbtSYaCrl+dhwdWP
QtXy+vIp0ZnhQOHgIasgMqoNDzxGbfpifiWl2ZUAphcigHRdzkLhXJPPTc1OWbzk
OCv6RHFY0YR+iFOZbVR8F0U6lrWId0pFIUuWPg5jpxbQdJA0ZFl6wDc+PO4jblvd
bDCeIy8J+HxYCtPhAxZRjhP6afRaxyzSU16gt5Xe9Hi7BxvhnxgVZFI1SA3Rq12Q
y4OcxBZ96afh8/F7eDfeuys4lSqyfx3yFSs4S2bzQ7k/q9pU0393G0WBjDpCklGb
BQf/b3Zh8+US6olw9Q2vIhIorIobeLkuP4Cxvj2FqD5/nFiM1l0e6Ht7teTtiYud
zKvVsgHQYytYYcESkn0fza1FSTKFoFhUEWcMcIyUYC4XdBJvrKUNKhf1rpz5xWXC
t76JKgz9tyC0UZvbHplmlmVgamVZlcPFg5PUW3iTk9uuLQ7xWjU24F0Go0Or9Dxk
OVbJ5LE78yF76S6NfsVJ3j8buQOuOyjWWhqNerpJX40tUVgp71ZMUUsEe+1KVoG5
i/x6NsbQFg7ELWoJF3lO7rGtBj4HnFCEi8RAaTb7P/x+cIaEfJWZt0oXH2rVgxFp
w5wPhVjoe+GW/031K+rVO40pyDACMl4Xsyrnw5VB25ooj02RYkNO98lfUW1zY2hp
9EHY5+GgKZM34Hap+l1jxqRUowQTgFRL4ywDfMNKhDZ73hzrOW7kUyP13jHwTwiW
xGCVBDSc62ijhf+4tszFikDXrTc9n3hvXV0lxe5nDBB3zwlkEXbDMtRM+l65cEB1
vg7BY400r/i9TYb9xsznfC4JeuixHjrhoVo2yXQSNukVviYKsKcHd4vJUCmBCaEl
90AazEInmen//TFPeELpjYVPaBXi7L6R9QRiYF6NafISS2gkl5Bt3yJzr3gTZYTd
dnHEaPEkEK384gDWOROD+MANcgdrJ4rwbIukrKGGLPGowj7sc1MR9Y98jUkMIDLz
4RydYGFm6/e5OwS3vAo7I24UKRqHpmcc6cULOjyTyr/RnJT/6sWAHgvOkRQ+Z0EF
2aBrLZEfAJ+ZyTdbst3MO0Y7lnFdDPJoXprnnllux+3sCHMpm4yMX09Thx2Mx3ap
ipRTmbSQYKx9wU4kTYbwUOl+grTBUrueHhoOZeMBcpvOlRDwMKw7MWoBvUDckwEN
1qNxRbo6gfdVc2+gNGPYTTfbEiTgrjpUPYijGh+lR9yNDXitkkj8lHql24qgSiKt
v+PsK0rW/XGfvIKExX34Fx83sRs8nnEklfMjiFoaeAIaNLkE4vuxQ8WA3BCPYO43
oA3uGNwpMRLrWfDgE7pJAOPnQ2B48SsN9y2r7frF/AHQmy3KgvjtjuKnJyh6qfg5
EpvjH4W6DlhHJ6HA5lWW66ZMv7yR3YoNKP+QJfXIS58BNVvZYJfox6XV1ZiZB+Nz
+N/pD96fOQe2Q+XHvJZseesUdexfXCDdRCbRJEMuP4k+oply2OXmhaUqJIN5PLkh
EWx6YIgLe0QfsalvqAMKkfKwKsX1asFPnw2hE/7USm5uxNY1VgaflJDFRgaPZDwg
yC2OQj99pUDweERGMubCZiGZBXZlljfhDsxaIj6xANv5RbhihCcaAhZW/w/QKvM6
M4uze2ZSId99LPoFa4NH9+bn6dH/svooGLNZ1CFAbpGRm3lL5lVEa55X1vZjL+NA
G/2WHo5HnDFenNdYMU+7Sd/UfiviN6K9KYBZlgIsH6i8EkUTt8LtjX6AN0tSmsdX
lIYiknwWitGE+ZNglwqoVHsRWK1CArMaYexO89kzQVsPim1Xc0AHyPiZ7pIoDch9
gOOuFPtdATPb1dUFullCYaEvK8VN6011cQgynMRgiVsh6EeBQEZ1DvFp12qYpPdb
N+y82HnEh+YTfeEpfDCM/W3SXWZF5S8EaJLgyxj7T4KQI1OQwsWDP61BLUrjutHp
4HVy7y3TRKz0B6Z3Yt9MNx3vYhOKyTlEhU4ArPyjad6hf7kwWufDyzOC+31mX48S
IXbtjN04lIj4tG1BfBQCk9DoBatllNY9WyYbkZXel5E0we9DlAWfSBbpU41JttNm
U53DkU0X3RVJBeknQJauBngd7uhZPSgJ4OQo4LZeTDJR4OYwE98yJK4YE2V9N6Bf
cKvsDyyENFWtSbgstV/S3A1HPVLDCxfXs6w+gNH5MbfKY7am/HjWfeoc9Oltejkn
sRzWL0eEwtetJnSB3B6GdWngNUX1SG8lK1rylzr3oWcghXKUuDnBa5bXf6CzfdOY
HDIMXG7p0CiMs8o+WfleDk8/UulxuX6f7i6BP/lXxKnl6D91wwIt7942GCkJGr1m
PYnpLA6MnoaumOg4P44kxHF5gARtZ1G3yl/8j/dZN6SdcNQxwn4sWcACUDwSjW34
Nb/OXKKehNECjQ7J8bt5DV9mevMOyTnpumLsmNIoOv1DPaeoBXhsqjgEkvopD1vl
+mbZjG3ifDvbPG2jWg104eDrUnc8EZU1F5qa8zFD2pbyF9s9rYao3qxopQMYr6SW
NZdBeOKHmEOUJ3+WPl7itOu1cAp7H2cKw8y8Pvg5Wqp+XsBJqYxLYt6r4JIKlhdi
RqEgg+E9TkOO/aN5Gc0oHIz70bu/Me9DAOvvTa4PmzS+ddKvJuVyIaA9kxnhb1EK
zcp4HuGgd4fuzw1RAGku7mQ5bzEQo9n7Hxk+JweTa6G71D+MiIjXf2QmJZcoy3Ly
uEhoiXuiLxhP1YXndNyEAkNDRG4qduWkBCB+j9qvVQBG505gvtAqBADzFRppJ9FX
R0TBs+S9oZOnJblP2oxObRfnhY4IrTp8lKcKPURfPWfC55JWXMbq8UO4ePWtMvlU
fPafFf+2hPoSC0dYkPvGWdxqo5M+PmH1GBWO2xDlBivsy3jDn50ZbZtKfdilCTjU
jCbOdb2YmUFDPNDM7pj7QTXAanmjrQPu/B8HS9yD1lqcSRXEGawcf6VEeKvPw546
LHNjr+dX88nZC3gKhdtHUazs3NOhp/nSjcJeoZhmeyR7YgwWbSqD2NVL6R3EQSPn
ffrGiHo0NPuOlSqDAqfnR0aeQErCpQ9PbF22nMzkd98yHcaWWawLoeyb6+ddOUwI
WPMLhkZYCLWeAkMdmMdXa+X2AaHGL4Ydgb9/lQVhpOhwVtKf6sW4MsCiD7ZNCHlU
bDOM28Z9mzhcG3VmXZkQpyVjjl+qcJOH3mVSHoeI+bNarqs2OESyLiHTRE0fPnI7
iV32D/o8XPIEAMNuj7lpL1ZW/i8N96BJ5KitEVBz1zCdQR2akJds2eVG8WqDgJcv
0EdcOqUEmYuWifg8IsUTJ4HWSlqHAj0WUEAPnLV/XlvR6qaq6rbvH8Y2/PWw0fyE
1HgqjPUV6Ac50LjVh55JDPBE7EvaTPRtG3RquEbax3CWrn3ZlN71FRk/yjb17+9h
WaNz+9oYwngqn32uzq/DFbYJu30oZB9ASXU4O9e1UU9d05uIORMZs9kuwSuO4Kx5
HhtdOQhQtaer7nYWXVNYbQ945fFuRETj71rJuWlfyt99IUJ8J/My9elu0zOt065p
ReNLPquXrX/pdbzUvL7qZ7Kt70gwAInTywm3TomgEseDw5V9CNcUWIlVPS3QM9B2
YP2yHfg9Gf86Cz8NQChzqoS5sz7BTkvM+WP1NZe9Habi/rQKK++NW5bR4seNM2CV
bXpI9E79g/g2ujxPzzdtY7WwHfKlEBS4tkeAFDP+ivQOU/Do50ohUg50OlDHRsrm
NZmZeG7Lu4eD3O4CZDcHg6Ipi6kp0LJSOkUNdkMF5OX/DWZ85J6hF4vVwtbA3Jnf
OCUTEGM8vKqvqMF03eGsenIFp2FtNP/zs65mk0U00URT9n9DqNpp8oGhb4vO/wGg
pjyl4pJAm5uXHYKRTXdeomfsS9bBjdqB89mcp1uOAJbAZc2owUYth842UFpix+Xo
HWbFnnQuhZP+fOn49b8WHitTUUdEWt3Z6EejHm1RMhVx4qU1cmdme6+koXaRI+pr
8F8d94bh0n8Qc7Sm2XqKBsdO6WoXtHi+lSBfVEeaIihDmNWu9DMzE3lOxGRFyudK
gR6Y3fcmAv/DIDlAE/7MYto47AIP5+DfdJ59ilyz2ItdvOmgdo/ZbP1G3Vthw1b2
YRpMtjP/A7o9mufve420etv2w4fjuySa0SbQR6qXqh7htB4qgYIHJKr5PUesoJme
7Z2nY/k+rgTJfLT4JVBh5GH7C/Gbxf0mznprBe2IW53KVy0vzESRhdsfC1JUXqCJ
MBADl2zOB1ucNFuC7mSRncfrquSHC+vUN7a0pXugx/oJkhfaZNpm0DEGlmQ/qMX3
pFhA+0euFOmyJPgsmdfWDFh/JF4c6Q6MPZyptp9ueVo5kUEK8kvjg9hHTR0fxRqB
qoMger/HfpHKf+p16PXBV8pNm1YMltyuVv+Rt1ra7XAF8DI4u61zX5N11Ipq0rSt
r9mBLDY444jDT01jlnhly9rUHXYeXJ/YFiySCPWHjeZYUsJVWmuXliB9SMmJpz78
Bryq9OylReEivxVM0rUQLA+eRstgQoIFKYO2wT3jlALWl4ARFbSVvQ/GY6eCHnY9
OFHSFijicNRPQ/QlzR1TdtLFLklCZWrhLisDsf890LhU42rcSNB0q9y46yNQes1q
okj4J2w9JSzfhB9D0g912rheqBilH1Vukh70+vHgPH3nvm+ZJaR5lzxSyvelN0NF
Er91YQeS+i91pYY64tamzyRUhT+GRG33wJSNjXTDgY+iGOG7k75WTciGP4Q4kzSn
o8ICR8DnDnQznYtubLInJlTwHKxRJJpIbd+q6ZwS7Oc/1elvaLdQFjr5TGw9bQcF
5Sryr25kVagee+vo94DLNJayWf7ZJJA030W0aResNSaWBgBoM1Q7f+S8vcCYDJBD
EFRrXSr8SmH7rk0PihXEJSsYiv9TkAJpbX7rfBNTZxzDBxVQZ3ILMPt+mzCQgnZH
IuQ6wVygyRyG2bHn0xsQITof//RVDSkzBldSKhmD9Etl6+X4zROBUhFpXd+LYUs0
Vke3G/KaBli2G01sCwmVS8UnTiffcnMyIIJ/lL5JDNdgpay5iFLUSQpGfQUSKi0r
pYpXyIKaszsmDZXckv2DMka99ae1u3I8xiyBFonszn8eHpnseqpiZPMZzA7cAFVI
pVU+Vb9/8ulo3mZJ2g5PLesrZ5f3a0B8RBY6Zg9/frBQBtRhxbqMAsUwrTrtWVlO
oBTV/Z5lU459N6iOs7OPan+q1A+nSijQAd9HAYEzHZqRP4WqG5kVkZkXusrQz5pJ
8FlSYi7VWoXzYDjXq5avj5SIk2AgcfX7Fxo/iGTS62xeQ581aT2me3eN47SXwa87
SxbMaAhJLo0AC2VwbyuR4VbAtKRvdb6rmqzKxFBPElf1rLlQyw4wTW7ug64a8sg2
j4dwFnwbdNsu4Prvc62XloUPHJYFhzzVNU7D4vjoRtHqAuO6ayHZEPlEJIvRWbhg
o/HuUA3C6794FlDS8J/cyHk5Wz2h3R5vM/mzQjNRnzkh3xYGJKtrXKMcpWh7lbOO
GODwnur4Cckz9TIwq60z08fPjiZxJgdPCq5ekXixkmLmcNwmPD2pG+I6eNH7DfEm
vNH0S2fAKmhO6LKRjw1Q7G9ZJnG4oHJzMYOeI0Cyjat/B0F//nE+RpgkOkB1KvzB
Ym1nmgWqh6oqsHHOMG6PGQxpl/slGNOLX0Y0o0c2hrBvw9TqMYhbqKuzFK42bb1D
0/AAhGsVkiEmUlM7pWhxHirInIBJZMrsPS5LZFgsKR4BcQKDIOcmekFAWPX7HgAR
DMJi8CiowSbVJDs6FRFtLkkwOXDlKK2untPc9OtJzdeFIBJSskdzMGdr56VIgh/R
kmq95XZVujn7+aSNTVTuv6v31FpuAfjH2YGfZgy5u89kf83H0U6/Wfw7miHhD24E
/D8a9rUOzCjGrhuCCtynWeiJOKnobruVxG1Kg2pvtUXh2wuPyHH9d8d69PCxxADu
jROmaa+mxIf8iD4EJjC+9Y0IiVYj2k88w5QdoeFmoCvNKB+PHvfsHAZzSE8XRKgv
0F3/pnLqpDmKoDFnr5iRG6UHD0pOa26gvawhZWrcQaXxSLXYGBLYZImXAHvF8eIw
TK7HL2s7kQa1L9LUmazXcbo0o0XSteCo6VusU3K16syYaa/l22Wgz5sqABfdj5Go
/YTLE0Zg4Cx4H39WIfclYoHF3h1sUsUyr7pjsiCdHDBFq6dyUYb3GF1V3cMkh8S4
+drTOQjFo5hE0LZEeh4r03J+mOhQm4PSSiWFAmlhKNgzud13bZOudVO53eyQ3oid
KB+UwM7SI/vuTAuyfDFkVuKZm6L9dX2nr7HdZcOYoYMeR/8J403k00ydYPjqSq98
lXf+SYiHzCucD3YsofOi9+rs39MvLiWx/IhJhb4FJYdQjwbVROhmnEBn4u/rxh7Z
/SzVbEQ5TqibsDEz214qJ+6NvoX5rqRY0go6CECoCexPh6xShJsEo4/wmcBkh3Qb
NAXWZJSnM1tThW8prvJdg834USs6caNjqZGLq/3Iq7Lh2M0MNQb/pSkoBmG5BpBO
ZnFvzZ3iRpR2wn/HzIUiouKTeIK8AO4UAfCOcz/fNVPn/QGG6YjMQo9CUmtB9jDN
qIo0IvELwmJC83sEV6s+TL9WJLF5bniDCC9u7B+if8Umwu3jA9YjR/oEokL+4x1V
U84FPYwoLnsBP/DBrr6zxu06apOD2OsAO4I+kYTnBebNoAVJG+TlZdiIumwhxdoS
4mhLnwdU0aFrlNgoeL+6NLhYiipDaCUAt3TaV0OkBjowwT+yxsqqi15FMnMPirrk
4p+9tJng4X7CFPdml86R0Azeo+J1yPoh6y7om5WUj+l4EIUg5BnQxH6dnqzXubeL
MlRM0fP/oZfSobJksTbqfACAIiXvYbNbWJJVTNNc+Dgbwt7+QoPqfUNJkheo8pd0
ln+HFn7rTp7twZ6+DmDiVEg3cA0Eo2vWKYa5CDrJiuJ118zaDAb800Gmrd8MUN2W
6gCG5L+yprajN9i2RfxDQOVQ4xs/IsdO7V/AtxVtVZ11i5hd9H01iKIVCqSH5+TX
9Iy8reyGO0qvp9nW+fmaQJXXDCKpwExT2yYciuokaeLz5cGR1F14Bb7UAUpiCEqV
PcJT2ukrCVBqcQRmeRMdKcBDBMikJCjMqEdFi388Lj6H4Mqs0N9Vp6TcyDk0WHVP
13WBFnJVK8zAvSI75WDFLAECzKwXDD1YrOmHJ4ursC2UmHSeTeiUS5VqQIMCLNo4
5ac38L3NRCIqbPo8Eqjwdog8a4LXEdU7oEjA2/CccxOp5Z6yqkfjMlgADdRE4FZU
mI8+bw7kTOx0Mydp14pippNOi0rH6M3FAw5Wkk6RAlLEMq5jYNrrJtIhcb+EdwPd
q640vIZSrL3kEduSTJ/jQoZSI8gCh4L3YFi8Ls4PfBjKq17EHiczBqwbG5X+ivpd
kFl/qI/VCWN9iLQ1O8ONGMn6hqWv68SU6xNNZ2L9aFYJ2L6JuPicwuVFy1W7YgVJ
5WIbIztM7VRWMM1Pz82kXqAsRaEOZMMHv6tgBc3O8MFYIH4Mqh54UWd/74HwmR9R
bT5VjBMC+RB0qbWDz2qs3ZPFP7ptaSdzqs6GkXU0EYvAKKg+FJyPzdmEa3Tbc4rf
UxVpSSt30XAbiHXF/kwG3YMd1WcXFMeM6s9zN44SfWkNSiMpfnNX9XvNp7b0h0Re
nLqYLrDx0yOxJnemQtHEsImzyj+/bSYUEudrRbISzBrG03UB7xmC9dOw+EB/ICSK
dMbbEoWZvVqg06tH7njwwUDynqGkXtjHEEIQqVjMuoNMF3MJ9f4VK+U1P72UYmBj
qPq2m5Cqi2qmO9nhL4XwTyioQGvmznA9jbR5hkGlw8jM5fRdVyVwkE0X8RMkXRNM
WPNCRxAm0FBeRt4qxgVCYENntwAi5qs+q8NLzZ+lPzbc0nXL6LGVzBNFH7kwRZdp
ggDiGlfabW/VekZORTTNB4E394DVGwW5jnHY1Gdq6gAb5cae5SpFR92yXx2EFXaT
XTK/iseG8Z74u79eAC59JmxCIVl+fifwqLLPMy/vi+gS5mayxKaF6gWPMLbRBxeK
2HSIVUofEQ29Y/JOeJtQaucAQUq7oz3rZZyuBG40hWP+hBMGV5QmWx6RjQc2EcUI
pFL8FGHAuuFvSY5u7/3yT91Y3IX3VDCtX1QvL15bkCmtah7pUqA1rLu8kdLy33WT
xUzIU+92OoowLJrqo11ikoOhvmDP0gAYMQjPkw9KUKrFbKey4L+br+BPRFmjC0Ww
JfBmVCS9bxHU/U+B1efrxaqdhVE/qCWNBBx5LXm2FO8iFwRzjrwUJE24UbJU8q7i
BsRFeXGhG4BU+riqX5/n5eUdHwqPreeTyaKeqJ0Gs59B+VcGhY/qx6Q07HQ8JAU8
BsoZa/ic4923TZn7c04mIyHkl0oiZKQsLOSBTj+l0KBAmTfjJWsYkkGmU0hVOrWp
feh7J4CFtVsXN0uWfbVfhSpO1kUC1eJ9mUCchtIJoBrys4t2Su7sEjg1uSRQOgWB
GIH7GaFUBA1poINrcdKFjA9g2QxoRx8Xb99e8Da9g9BLuJQi2kACaS0UUGQ42XdU
n5k9vxMY3HPPFq2HTd/RnojTtOBU0zes5iEA9LgZxdT8RI0DgV8NBOusZHG7DMd4
AUHPeCQktEDZw2E13l5vUJoITjNq9A5g0pmlNJSmW9ir96xuhgZVsY/PFN+DL4Jf
4WGZkGOCqqVqKBzHrgiXEgqLqUsaMUlNTWTxxRBGPbbikvRufgrJSidWhfg/pLHG
HXQdXPQ0bx4p7VpsYwxamTojmVSLaO+qWk6xYNygoZYppbTNu27ku7Ew/G0JUg05
v6Y8VjCzJ2tF1fXCV2UGtd5v03c5mKAyerq2vB5HhiYBj63jG101Zs5mnVI8LlM3
ba93zHqd7exfMH8iVo5dWfGrSY+jKXK5f5RvhgUVQt9f+XLeDdhZMjQN0Yb73GPD
fMeuOqeAztUsLi4e553cJr/69T7kflanxt5Wu1FfmaPmgdfqF59mjiU9/yX65xNO
q8JaigZAturrjKkYac4bN0Ingk+QYasFjjHIZ5isiGFqNW58ACAfBQVgUTjZbNNT
zC9Jn5N6UCehI7vEJi/uvblH9H7PSuvTKT4GyyfNsae368vrVSm7PZIpR9Fy9jOB
LLEqexLuwuN6rru1bx+JhFNiAdQx1Xz0WP7cmnBsdLmVfTUCSTl0zgv/Sn6ajiOJ
dGNVYSzTvNZkIb4T1mq7iaXtlq00l5JK9cPNEFypi8bZPuwTTZinF8NdB//SiTzW
WOdKXUWosHlBMcKaeRjgqWvNciuPYZ5a0ntC/iNJNEt1qroRP2wl7uDpLkxVTrxg
YyKeww4/xJzkrpytQ745698IL7CCU6RPkSA6D0PQesB7tqGU3V6mSM7I/s/+LQ9G
B30X/OABeUjHGQB26Tphqe35HuQctRBe7uHqBmdMEqN1P2w6yezh3R3yNAfyeIF8
LQvu5s7AI+D+ElXaCfDMBUToXQ8QIbC+ktj1REyGOfUwz2KZvGUToqqJOwoMX6VG
YYO7BcwZdFPm30uxUVxNlMK3l419cF/5G4vPryaNHimPe7sPPUPN2cldT0ZRcDJM
N9MJtihCf3qT8y0gBN5njK/hMMZGePjbfk79eeUDvpee355chL+NlibnxUigq7Ol
+4r4RP65dqdCBTaInwl7Le7yQ3LZKuSp8Sur4COJkwppU0FTL0P/bRb24Y589Ok5
ColUCupZSMhSDKh+oIASAFzU73I0yalt3UqjL1tPRKv5TaEXr2nSSCpdM/5x+xbp
2NBcgsPYmKmrrstAatbkM9ZCJQJMOr8L0a2MNGsvLE3NAk4nJ5PpCw2dHHeTflD2
CmTty6ldTNvZtnLfDkoAw5f9ZInRNNyd12MpXTE7IrNn++T8zauvE1lf99ttlxjd
FG5I+2rRXUTtjab3B2EfBYWG8yzdnxdNPDgOUccyB5knQUVV81Pt8o/dI26Xinkl
uFwucUrK0loI33N7LglkRlK/KydoEFOFDzBt3xAB1BJNfqE/+l0Y4JfzcuC+Ehy8
Rb/177eVKFrjVo0y6goYzlIIcYGpgLNkMhOLa8TDl7BTjVoIKsiBd92g6M8J6/gl
K6p3VZJO04uB3gmo3fOS5FlUIv7BCtLAYf+Ee8wNn2KMT1j9kt/ZYo3W8fqCDlTF
IIBvS2yBmCwISzZjJ6lEjjb08ee4/4osphd2/ZkeT6e/o/w3M17NBXqVxnAyvade
cOg2yNs+dCFzNGMPCwGeyoghZZcc3pCso+rL900tmCV2Dwv05QQxfzE+P4mehqH5
0WbBYi8mnwFUQipcwn+rcFUUCsMXyFB8kLjzFdbOUbMPfQdsh4gxuvtdxwLMnDTu
cjzzcnl/Sil4FsTwqG/Zh+ts/GV5wZ+kFPgkt61IWCMHoUQLtMe621wUApD3KOLt
xPVbyS0EEIWzv4bDL5IDbLveGVZzo7dU3MEh3GyjfU2XAhuJ9TDugEw7X8ehG971
8n0mqc/9PpC1znnYXQxMxcCzU6unVdUqbxsWa+Mgav6G2cMcqKOXKl5ZAq4NDVHi
t6BVnRFdgvkCv2LFgdLS6VjM17KozOxZYusT0CpLQoIMsY9XODmAtBeifs1+ccr1
x2jzHxwV+DS69CbduiyzRx3LwbkGyOEp1g4F9OYYpvk0UCRUHuE7BYv20YEZanCg
v4PQdVlHLVCSq2feBG79trmK4TyuccJHcwKXxIwlyp+Y+tYRRfGhpTHLj6+3nPGN
7s2kep6zy+GAFMBVGwcnN3WBq7uAOltvshNQP5BuSW1o440emlUyRblakoraU3hg
BQpQPIliP6kDm7Q1gJV1m8cQWgEcAwZIPR5Uxkw3kU7SnoZmFFwBB1qUtjNDva2N
LOz9oYq58cFWxucTQAmzbu9lGN810XQAHnY1G+EYMtFTnyu2rS7O9UhyZPdvTxtE
ZU3qyN0TjAqCWvKZKWDbPQEE63kMi10WuTZSydjPdS4EwUHsgcRSN6uGHVqwREwF
dOep+MxbqieaqVOTFIPIHBrrWb3U8cLNhOEjTicuWZC0VPDo0dVu7ZVqZBqoLT0F
T4xuVB2SPNSNLHZMTunNGxEIOIOWea2rsBosrUiZ8SmEg6o+TrOZd+VfhEtt8T4c
d5Q/sUDvzY4btTZVKa0pXTA9ptEJH6wEYxYWGkHP1pMsarB9F9K0Cu2a2Qos/BJI
YRn6lUs78n1nhwwmuWf6hdpkhwd2o7TYyxUnQs1dhlgPyJunvRmEB0beNxm3WddV
qt5K4WqqbmpHbbHEIEwhNQ2tOkUFyshhiq4H25Gh4kMs+SwVk2OaD3fjgL0rWlkF
3zJLfj/LVH2ZPujnZFff0GTz7sUHRlgPZUBkVHiun0lczMlK1Gnzxvn0b2OCeaK+
aP/f4ieL4TnZoda2OgYXjfA/Nxt5UqBPlA8mSDu8EDIX9NOrHU3J2eZ24yoreAv+
FklxdW5G3bZjdz8iY22nzv1ISaPfxT+DV7JXtuyQSrkcrYK0Bh+UqM0THMKQxY1W
JJnOPxZmHXARX9r8xRJYKOoF463mo+PA3jzGoL33ESvE9HLkMdnq1qRW1hQ872YC
F4Y1+4dR3mMRcf0qLo1Bm2ZvF6ATQh/ztQHo/8mp8jhv//F/5HCpQ540dyhy7CoP
xtvubpRmOG+P6eyhOWK99RpRLV2EzHWWaRkdCZ/fhE4yE1Pv3X5y/gtev7Fgf4+5
P1190bj1Xp/ctDeQAonNYQFUjTpse48JV3pdXswTR1oZIVsXTQUQNBV8bwc4MMvn
T0GfLVTPpF+0UXLnS1QSyTmhwnf76oH0XxuiPaVtWKQyyqjnlpnFn8KWlD5U5SNs
pNOmi9zwia+xpSIOQA1t31EDNWE68TSN3MiRR4/tNsKNrMz/FvPEwnUSYP6PMdYj
sYjlkLUzaHFeZM4SqotR1MKD9zqC54pC232vv2RbLVqqEcaaUoOWF68SWMUa1mZn
OVwX+aiQ+etfuBGeSIyY4tTy0ziq0uS9axz0pXBJfEvOuwVJLFZcqZQkTxlHzx32
45rB6AkGrY6q8MXUT1MnM/phkif6IIbYRmKntIAcLhypnEfauMMnkHYPbReJPWIG
HMFLWrwVNj+cUoq4+GEneRxYb+R9VsNGr1xtTCP8/hLXkEhuzgAKnGf1WpBn+bOK
wfRdC/aIdmne//WiPhH4Fy7gYctspkOwpWo8MNs+4DQOkwnO8uWoQ8XA7GZ3BylS
lw9GTOak18+8jiYehQqI3ScsobzDC2Lwpmka7mv4IM5yK9ov0sstFuV6CPF7gPd8
MPm9MgF9rmGLvRht4RoaBlUyrZD55HTnIHhQlOXDEW77OoKYxfSPQnVlLwWWMDA4
thA52pgKBCJ3GeRdDbZxt2MHm7hq6qcRa9osTJ7qU03LQ/BuYaxuCg3a4zcyn1Mo
HZxMg8iOdrEheHLZtynBTrWKqKTj5WmVXbfG0UOj9aPzwscmCvH/9smGqty/9SpR
p2kzZyICZQ/aFUTfFgIB9TA8kEc4bQ06OCV0apc+Jw6EwB2GN5lLbbOqjvfdhzWF
x2iXSmk8s7Ds/BBlQEaKtt0DogQtk9ErtaGZUcOg4PuupTQJSscsKIxD/jro/F2P
MtCsJgbPn/pAbsRIAmaOBgxbp5UwVU6S93qfSRDejIm4el45cdqYWjSbsWanmziK
aQIb0K7QQBP8aKlmA2vpzjD2tNcefU+EAi0TjhRoLXscnjF+15B8GvWcuzK20ex9
m9dwwbQltdGfiSweusmv4f5PVeOwe8YGiDOCTdYl9Y/zJ/H2lwuJEt9OSc1svgY1
ukmAlGap/oojqWSxNFJQeEX05dHLLWU7IRjAmKasGzcRAmBiYH2xWDJLminWi7N/
Psb48Ki7N0w616N71Q2NhDIiEbnXfpMapXl0JjkSxpdLvcT48lfb4Oo+/WemO237
EqPZFK0dAFtLPZpsVH61aSG5X63S058sHJ8+D0zzCelDlYEUM4+ACP63DkAeanVb
0JAALYFix8HB9vg95Da8QQnlaxvQQuLb2VDbeRZiR3y51qUfixlumlm0Isgc65/W
I2F3VRjrrltAwpSow0dEwwIKtmD1ccdZD/JKn3fS3840/fwSxn+k0nkAjsfOfO6F
fmGgtfCzJZ9qFvIjkBV6IbYFngUGw3KFgtuUPKWhBo1p05DOrwtpg2QiuVu4e+IB
Le6EVMW/q8DZKSyzEfUHrt7wPQDCAy12jPhazdQwxsYCyoHfx0heuJcD8vrxyVw1
Bxl4rBgYEhhntVV1HheBKoDQ+Yg4ezrFDSnqiRHKhApLrlZ9kgaRvBRTzTmF0ihK
8Xm7pPTF2h8xhe7vfdDx9ozVA5qZ6UGd3vOYK2E23tJkei8yeiqCP4+AAlH9H6qe
EUWLkg6Mv59y46CreBkhjSGEsNsh+oW8mG1fzDobnjDmKezRnYxpW/RWd5xLn7Zk
vI8MoSIfzFZqYe6V5KColgKuNgrd2ghwji6RoqFtrmaUbTbZriGx97XJOqc6ULre
Uzfg0vkcnnuygR7J6bAjQrtwkBr0sOfPsgErf2WikeT44t6ivbiB/L6QZGWGWYL/
/uWCWA4cmIwDNAJlJOfDvddduj8RNY2OanimIB/8tt4V4RF43VUmPXOQEI8z8Dp3
nFaLCiF21+X+XbwfJ5gvmURuqgPWkVGog66yjvIy3+UOySRPAaWFNnybMR5IoF0+
mDPnRMsdzeZ0kO5pn2jZPzfhKtykCwjJaaVitG0IK1lbNkjydq81ew/1pV9SxmLF
6kHN7TTN7ravFO82lCz/bYVOR7o9Erg5UzHTtkrJz+to52AnWEF4Su+0aszVVzBu
94chicJQt0Ccz//xdrgk34OFGggjR6tFzv5gahilY9hBWHyHKgAH7qSj/nBL827p
XuUG+5a916pNoHht7z7neXo7XTxoQyjV+Jh2bVU4shuIj5oEqD8v7er/z7itpoIU
rfeluUrLJDf80syyvT4gxmK8r2mmLI030xY27/pgopCAXNvbjdQPOd7PhokWSX7L
I67RwIl5CSwVovGHpK6VLGPi3AaEpXmeRKoEakRlWv+bIh/tEJr58WileNbk33ao
ebXZ+md9QKfNZGmA3sLJy5J5b+JukKOoUfXVsHlXREq1gaD3bwB7lErQ5qmXIHe9
bDhHqboEcyk71Gibqs6RsK7EZGFkE8T1ZIJXa2UP5FIaeRjp55kH9BKHWhi21+av
77oE0m/jqHYtET5d/1Os5biHNR9y+ziaihsP2socac4oRowszALqMtJVwdxlOyXK
P0a7nDOUTPctSWXjC5rZ2wgOAfOAiExf8ilEBhdS2fg4MXyqgzy3m/6+sepUnrLB
OIrKHTp6ZHRqMiKbaKaWsAM2Il3XD4vFTD4tT+0l9VRwoB35Jy/DgXRxkrb1BQgX
0/ZwBaNCBPxcTE7+XfQ8rPKd4RPrqqyLkfRpwMermMF2nyqjmLVYFILSjEitTekz
VxX/aGse37zgVHvLDz3FZYHGNr6W7Q6TXruTsHSocs25/rKkIIiTWy2WV56NqrVJ
/DOkeK7ZzNOJZU36mQCDmKV24Qmqxk/ARWQkPRoxdJjJOAholksgN4hRIVJ2B8xF
9pTKHpZI2P1cRtEHiAiQBoefeKmP2D5sLb+IE++nJ66BMU01WRwaBmUbqMARQdIP
f3RAbWfL8UW3KXX3xe6apPJrjBctqklNzJ6cNSMYXvMwThfeh0RFC52yixXVqxFK
s+gtL+usE0wCAJ+6tt9qAhAJO8vbz7XCs51V5g5H2gOAFUDPgMxy6qod7K6Ho4Ky
plwwqy9OYTZnHSzMxU6aG2/cPT4Gg+/ZBj4rKIsoq4Wbc9APWeMsReATOc/7Ihvs
M/AQUXOQOHLI2n7PyaXi4Aty+5gjABCegwsM9tePj+l7XDqrCfPIPP6NHG3sc1OI
Oj2aOaLL9C8cSDLPHBNrVJvpIyc/DzrmfWHuVonm3PPvF38DXOPmr98QvWHxIYFB
1bDNgLZXgqL3uvkia/yV88WwfaX45/8pi8AovdBlvjUZJTOsrjKLF+/hDQA+A2/x
jqM+MISjR9UlFjfBzzlOjExjxUUlVa9cZJQUo7A9KCDTtlDpRdPwIAmShXnoA6Mu
shTt4PcO+ID5n8P0mLSMefoUJPuOzp6M9w+NPz9fCizjAKoYQWAztqjKM0CCGasV
bwv8c5y42zZig53tHQpsj3+fvs04KdyDxsGJ2NoRn0wj/M9QplhuCiV1TdRkxaVJ
27zqG+9ZPRJO7GYjDqze8Nsn22EZzDJZV7zgWM4WnC/EeSHFTBsKZ2zf29D4Ragz
2v/5TOY/W6CMRzN3wVCXaHJgcOGJF02Kuq86+OHp9Vu6RsHsZY+XEvb5wuM6rhq2
2X/+7+2X+7ruq2Nw9E/MfBQ1z31uFGYg2bWqwoTM9YCLvGkBazMQfG85y6C7J0QK
xuog6AzmMwi58pCuITgVTS0ZFDWi0FFdT5F9JsAaoXd6Hh7WifFWHi0baSFYFnYp
v+IJX2g+WEvee5UXGWnmJOrbp+Su+3InHezOL/heDfVa8b4SrDpcIWsUWmLhG5lD
1Xi3ivsWg/wIMv8tkNTG1ju136yNZkdRHzjllpvXnm11l9vd2BY/a7+zZP4qmPvK
jXOl+Bdx7smOvNwjSsaL8rsvTuh6nhGVumhowa5EBoKUC9Lsy6Z/OlteK0PcEGbR
is9xRQmZnJxYLF3xjxoonrmmWJiMbJk9WJUCeNC0fBv9E1TvK7GV5wojoP+xEeFi
ohriZx2sqFy5c3yj5UHsiVARWP8LO47AxRZRekGMVINzbVdS8djyCcn0Pn1qQ5D2
cq+v+bJWsDGOIqS7+cyUMy8sg3/wzlgMxx8iLrbgbpufU5DFuD+/NRsBDF1YvLHI
ogD3Pa7u7eF1aenFexcxCRBDSZ2DC2GR8QYH+0pDmQnLvKv9FIFkfGQBHVrM7ZE0
0r1hCgGq/FQAlv66kfPwgD0WFRmJUtu+4PHwoWFkUXeSlhnk3D7zbHuB3TemVi1H
Mh0syF9VUaY9oWd00/y4JrwoyK0b61kRQWiw0qktit2rso5fGQH08oA42S09Oxbt
XFcl86BHhSfQYxU2Y5Tvn53r/gwzoAPO7gLk4pZt8BinSmyIxMxODCTkNBLfXzE7
36TWI/9bhZf+xeXyyv9tpLiA8FZ0/I+okwO+v4eWFcsXf2kE2nHSVgGIHD2lRhRQ
Plyj1cSF0fJi8MA/g/YNngtbOpKyTqzfYEs5RHSh+VTDOJnLjuC+BmJdj/e4yBoP
UZLPBTbCktZeVemrIOmaQspNdeEsg+bMRSpiD+vGapjx+qrrskxlPVbWdW6TJBQa
fOB+N8sdD6HsQH2TJCPaa6BPfavdAqYm4LHSmfekvjElWWaIutwFygWH1F3DSnRv
/+OKl+c+ZqVxDRAsunx4gIS/aV6I1hPrtR5Elcgt2+A7Ak6gb1zgrG8YcExEEnbr
CnSLCno7JMWbfOGWQJXP5lQTm6i/TT49s91eNnpMv8XRsSIo/nUB6fynN84xZ1tb
9BSl63J1VcDh03f4Mr+l/b3u4SGDH5hnMH0UTGBuv5Ly316tIKavtkTjns9FPWS1
HsC5PkN1/tIWBYOa7vo1FW8CKYDaSZ+InaoZBcIm6MD4B/tq3skqB+e5saLtylye
PWSvoK0KzS+8N8hIy50uhe7KB6WUcM6yHYq/vCduh1Iwhh9u6TX64DX+0Is5yCo7
YVBtbzZGeBI35QaHCnRVwWrT20zOxz6a1B85ZA8PZC/OelXPhWL4npFQtWXdp2ZX
hTazMFnrGHhpfnZp8Ai6/5JBB3f64rvCCiAYhlAP4AsgbrsPFSsgKb7D5lsGSRJe
09dcirai/oSrtF9237HRXEUYAOS/S31Gj4GaSGJsTxWGXys8UUKGEicrhCsFfHMi
3Rh88K7xAD7VGXQt4F8scldPPYxjxDpFE+pbWdHySzcPWdgR7Faf9qsKjXVjkXuB
NGmYEzcc7vKwpKTMGUFyOk3EgKw9dQimfMLZKtt6Z2QLmE1tRpBeo/ExF30BZ8/1
lfmm0rKQokATsX9LJqRjyVxjq801PahxEqM4FhETsHqt6nm0bFK1W+XtWclREHNL
u7X+Nyl3elTk3LOe534VGzvJ+uv16nu8C5v0arTiAZEUa8LVO5qYEz74b8k1T3wF
hcWj1VOnytZK9U0x52+eSGfSrPCuYXu0ZKcVVITxVgXtMW2gnMk+lXcc9HrtXlrD
tMkm6tQrfPsXuewOzVZklbnYEXKNB1oNnu/mkaYZpAALiuxIdOcK9tK507Pn7bsv
yr9HfR9qZvRWTwU9qSnvibytIdponfkA7pS9yVPx8SDyzhu1exUEA+5rxfxzsRgr
GtV/RIPjRUOYMCA961IbKdY3DaBLO0Sh3btRjory29cHMPmPsZ6A/6gwaHkhzHNe
zlCIlBCwkkIBaMyWuEjM2eKisrgiHerh2gRjSC7rTmZGPPnNuqkqz3Uq8a/YxiYv
G7rIf6YiajBE+J7KdjKhdnGTi0vcKMM9c3lw8hh0ONpZ3berW1feBtMu7dDB9L71
vMDFyl6XA+50kMBVPVWEzykmbq7eD9U43KbDqAKY7CipLmzPwH2Tz9UUPBQ4zqv4
/rtoUmmSuuOL6CvdeNrztyvPvS+EIeAltroUj2pAi8t+olfZedPhfcESkdiFUlUw
4800CJK5zHnFaiutQPCHgnjqW/IvvF5ZLXETIVzqcxxuzw0jHxzVc9bzdC9uQQ/N
O6sQcQW6sy0FfV7AkY93cq+qjUZfFKJr0mTg33P0y4eZFzLkuu5KO/ueeuQqTacG
J7DcodRpipYA9wOZAdo9aqwWsPZ8RkKhrs/XMLtlHct2NlRUbOaakn9TD/JAneuA
eSZIa0I833/xbQFF5BSJYDuCmrot9kjzjIduRm9EJkrUVVGHGibFo2G+pinuXuJj
W9uUE8/+8nkcDhAS/mbzoFt7IUatjdaI9qDzVyvKAH7XC8uAdKdU3yvbREz7jyfu
1HgZat9PhZQRWXSpFVXQq780DySy6vze6dggu+OZOnE/Hi3irG9kkzd2Z9p0eQs6
tjVXDQO7ehhpCb4IdTYtH400tPCFUt6FmXsHcAsD+mjV6AbMh4PgTLr714ciViDn
+dFcfXHusk8gjO/ob1euxrY0QZ9x6L/qgiHX6fxO1BA6MCHXmDp2Hmr4gaTayDQ/
U8Tg/+WKWZyNL/QUxwGUnkfX9Nf5u4dhV206I+tbYMZ3Z1Hj99rXwDfjMVDKG1Ym
ntap5RbjNJCvaTP+7uI6Kui6zWOmaYB1M+UD7P5IgY/W5ceLOMlegeTpFBKW/6Eg
SuY5j60R1rBsrcagC7SDsd2SZGqcwlIanVL28t0jaOxeUD5bKMAsA/fTpdMu2EQV
9X/QJMkhcD+lsMG9sq8gTG8tNJc1l0fK3p6IxiBAkMpV4M3eyt1p01QJ1LvWr8HB
9ULq9TmnLFTcgN1ZTXjUx1/4L4BCeBnAjWTIUyJq9Puxmo7w7kPXtFvE60UYrT68
wSP6S726LJsvkUu6oH00zmyL8ogGZPLEJQCQOQZKZIM14t0eX7ygNixUUHQ/ufRn
/jcp7SNhJT+6oFw5UerKD6prHxR6bcv/NorbjlHIacFRAZEgnxkvHH5tkL4SAI/Z
yQKNaOfRd+SpMyC7hah7w2wQQYVU78ZH/59z0vn59XSizM9hrck59e+bcn+DuEFF
kgxBlN0bIhbBunWCw3C7SVb7Pcp2pxVHuXMaRIEEZ4ksAvFQ2ejL9jrwSaZRE0+D
2dKRnuUkc/OJEx/0pUoaYEMNeC8jswyIkg4MDa/h4Xvf2ZRlQjBAdE1dKWdXx9FH
rjJWshYNWd/MbQw4yVPUn4dBLzydEFGjN6+rq7kBQrg/vBqzVGUn95xiwV/Ti+93
fp1hCmIVl5tom4A7vLrOngLsIiaTfQpeuyA/9zcnuP61BRkqgsU2DrK/Z0ZpzwEl
LLa0++TiWNIHO0NbCqs5gUt/aernT5dWXWFN2lO2GbFIKfyiDO0wiEYOW2pNDlGR
PEYU/LGe4/HSeF9av16mIJ4bx12KJcCfaKvM6/K71MIxI7G7/j333GG7gWIsvSXN
fGU3HA+a0Q3exTHkuIbZzNUdKQEC/l9s520UxuyKvEaKDZxCIDiFqeTppVrorE4P
HO8CksqR5Iumrenio7fUTL93LS+LQaj+rJKyD9ed60z8bctksF6nV5KAhbqp4gfw
7ko4n3HXDaf5tUNAYzsZQb5M13umy/5uJ+nh27jEefHtx1V/L7Ql+9c/17sH24RA
3CGUGp95s8hBj2C9mPEDrIV8Sw557oBN7Ed2XDrQIK/NOMj+0QY6OfYcidCKv7BA
pANEZ8H7fPooYZcg8WFZ8tBoSsKCimqZ8PXTMzINs7ofsrZsDfB6GvGlsS3RKXbX
8WOL1Rk/Pye+L1riSdpkK7n09D2ptA9oXyk9ER1ALKa1K/2OyZTzU4uQ0aXZg0lr
8jhFgGYtZd0Oxzh5eyd7KSk4RT8riqzijb4+Y+rn8l1Be9eTwtCM+111CC1fCAxj
CkPVnsLPuYgbk68l+jc6W3aV58q3hZeTtBy26ChExAcrUhGwNg3bsy9BtdEjRaLt
4uKSpu8xlK6B0PSqaGBr5dkNXOLVquYQ5CRxngYzztatAr/RHeVmvj5faDpu+myj
dIikspqdpRIhNJK3jprcUvkmeiOg8yD1okf8otD+GBLl05in1VRs/KB2XUOTQRtK
bQ6k12+PRzWdLJM8+u/xLSgblVIZ1oQ+6DE4f0IIrofYZItGuxqCOAbRCp1fXB51
cf6+D1hDJUWr3RoboE4xomu9XfUgON/tQAFgTKdropv3BFmIZFVaKr+0JLoV58Ba
JG/8LxwpEJ0/hySJR7QD02d1bd0pDABbw6gpFWslMD/eJ3ei+dZ29d4DMVhfC4Zj
Xo1vo/qJWwG+j3PGt4U1XFVFI7STxzaqdkAO3vdX78uoTB0hBw/uyD5lYfG6XU0f
8zNk0Fi9nOpMrkdtmjZID4WlnofQUcESpJjuSJ0cZQ3xh1DuN2e0H7rzYz8TnDFC
KF4QWoOPYsaiJpCba1yq6MzHCKCSmZtDDeuNkPe09Yvdd2e6x5LcX28OroEmmNCt
g4UkqG7bl4z56ckxB8+UeH2ECg1bil9T1y/VSuCwFIH29zH1R9P+D9L1WEqrQO7e
puH/zG/yJPd8IQ3feBAULp/lMBkloEIrkruLwKhU/2sXApr1vaUm5fXKsi+dOz6l
WC0NJDzKHmyjg2DPtA2Re7dykdMPegMfhg4jXtTxwKRaszBTlBX5dYTaMA7amaMe
pwo0o4Plb8DaEVv93YenvS+VsenumlTnY87pSPMg/RMpxgEP5Bo8gAlrDiNJlRkW
NkkpmXqo4NVuaixDtTfUG4zHhq0eeKTHOgEOhfQ+mmkoNX6WcDijxSLPL7Yz5PP2
4gacFm1D5VGVRDokJhOBTAm76Dt3XnGQfE3N9b23COpB2skIxGmLIu3ptxdQdN1q
8376miK+rmjG4Fjss9j5lqnmlNrNcQjjbKEwgjZOktAaYnptIilbvdnj37Op/QZ0
tHpw3jYajWhru0fDFfCpoeH+YT4RJCVfI6qkRbydeE5kK0T2020lgiqN2AGvaXJv
1a++pohBn5O/C3AmAQmqBmg+JEic+Lr3DJm+wa44D/t24pGMX16Gah/EoDOcHfVz
QSInHWX0kI/fl8oc0nbwHmQTWu7rszUnVXnCkfPqCYsM3hrIZHM4CSEHlAA/4OyJ
ecQrxFpgIoVNr36TmZJE6WLITYrjfz9vOUJcNel1B2R83VQ2u2oNs+SA0YUrT+uM
s1qidHg+XzmiN77bZSp+2Pf4HsrW0KShvc82VgaghquCft9EvK8pd0DL6menIBs8
bm21pSMsloZD0XSauyvZA/sc9V0uUCtY0OR8Apcj8mJc8duIBqPhe+lKmzh7ngGt
BCgZ7cizaQ8/P+B84M6JR3uUu+b4vRbDYVJtkRpt9Tvd/UYHhkg8863NlkSmO8Vp
ND/WcxWba1M6dUSA35afwHYN3A7TVYCQS65V4jXL3y8669epGMEL1aE7rUrqN9BZ
HU5cEU7a2OMAWtCCHVlToah81Ns6Bg9MVPyvAfGAVT5u0iF3AwDzD8uRo00YEvqw
/aBSKGxvihiFtJH2Zdf5AAJFQZSUVF5WxFzcM9WbySLLkuS4l1dFcs8RJcU+bdgo
VjBxcBzcF5/Y09gAc3h096rBGmTNdxXn1iR6aFTAJBU8k17HtGBTWKiw+WQFLJVX
xxxWkFe1H7WJ2nOVhuFl7nObYDS5JO3ggY5eFNg1/TslXmPW6eJRrL5ycmjmraa8
08qu3gNQ5mUNtfbTjHLOx+31FTBDvRKLqUJDst79WlVYAAIAymILkJSXzZy2CpWP
+ZHOAYCt9FOjNBIbyP25LbkC5GyqZig3TUOzKNlUscRd4QJDCSHkksZJhtViJ4JY
QFeqTIYUpzOGrDR3J32mFPAUlZlU4es/Lv6c+gCyO/BcEHbjfQvlxFhrH70AuBUJ
5rSpv4nL3fWZpeCwlWv6sAli8Z7J09gKfjec72nY4RyynECWOo5ja+j/6TkfsbSF
wMF2T2KSZAGruRiIvrK25eFpBksw+Mqc9VkgK/xPKCb+AT4okLUMLvAj7GelKXl+
WQopxaPNq5aM8hd46fYH03XUvOBXZ6LTvYUaxv4+EsWb7GWJW12fos1i1lyttOi1
AwsI1li8UvxMquisZ3P0/sefMteSN75yvmNg+UwBiYEga0seHvWgbBM8dkjrkRWe
ZxdCR8BRH0DG0YUpMw3J721x7PqqHMQzfVeqKnxyH/EFZrwA2ocdtJV6Swt6K3Fk
Mcptbwlr4TZvgQQ4lfb7rWAyNcSwvE4Y+gsd/ghBd5YMGcA2iFt4h22IG2xyq0K7
tgZb5zG03KsZ+6rr4d3bBEWdK58bmv/YF5SbZMg2tMMmYet/M1VdHGEKbQs6mbWk
y86I1/VsWoYo4IrKxbd3DrqAebMjMLqclLUMc7lHBgS8knE8LN5S66y5L7xFkqbd
D9R2BPfnh7US7x2tMoWzz35hXlzM9jOEYRJFZU33MD5RBP8IUhWhF7vac6rn+iJI
MmHHVr2NrBmaKy8FFDViFUDrwYRzy7oO1vKG7fCbhVWJlzly5XxHJWNKGbydio64
mGKQc3fmoN+29PMe+/hTmVY6LXyX2EBCbrnRgJtM/ufFLmEdjlBL5+EpjBtjn3VD
iB6OPQp68r2qjUZ7NTax8jmoVeG5YYxOUaNUsYJHKxK0vFCGNg4nUr9TG+oawQXE
txBUPacexqLUxEf4x4ifPm5x4EwV8uABf3ccH5/uDsNNMv3I+cKFKD+UYrpbN8H3
3qS77iNKw6S67LWDvszj1mSYUodyhTL1ylV/oDirrSzq9ZaZ1e3ZBUl9J9wcDruY
PFRTs4hhdJPhs7iV65/EvG3Rd3Z/Az2YYsQ2gVUFAHkNvkrcFoAsPAozEWXFK/uK
/zPGN+h76nxMUZOF628nRb9LNRM/B0E+Y94zh/axX5wMxmzIckhbdzwWbkXu5JYe
3qb3q7erCU2qfSmLA9KKwvRBQU8tux05Wf5DyLx2lKXWI66MvdchYpP/iMfseMv7
8RCRHWhFaa+KlWufrk2y2ETnM994pB0iwx3u5KVpj8aHnGf2Bf4qEUCDXxjYWFKm
ZB3m57rsojWPjMX8JpmgWJmcAs/LFrgFmAygrddrCUKKvGLBJw/3JwelxBrwFfgx
f7iype/Th3OT6xc+8N1kvdZDL+gLxiklcksMU/RI3djikvB8vYHplARYHRn9//0L
UOc/HtIr8vn8qG9PqbZgKeBLcsjn7y6b51fBC9hoE96CWgJY5vndgYFW9hUyCEFT
RJq+ofQXquYQ+1IeWhw8i4+6cWU5SPQrN12YyZTrKD9KVHe1Dr6g8PkAVI3cm2Qm
AXq4H9QYBmG6EDPmWfy/ARGkfsJTiOkrfPRiKkwvaT/wPwrAahkCnbNv1UoPpcud
eD7JpG8/023STUT12W6lksmKYFevL1eqRCvlfvKOK5Kk8Dxxq93LneJmKca28xGu
c76hFrM7HXKHYVpZ3+qzCutM6BLs5h7b6zY87ASH3aVXN9I3jWF3d6FUTR1kXTRx
vEvN/8fNDDzMZd4rLQU6Mh85u9Zk66CNNVnpiK9FxCn5+R9R4u63QMJKobezWP80
XoaHHaLjNOeo7vnLh8uSxMfTviPA2Kpumzdh+cAz6XBf4JDUdioouQ1m+i+MPCiG
GUfb2CwjuC43wNrp88aCEVvdHD9bKlxSRBzTJx9Al83TIHKGwj4uLUFBOzdUreAL
dWiQZKr2+zGS+BEdMcGEFkqBi7JWFWRZ9OCxFXqjKoIMH3v4Ry9B89pqQQZhzSqu
3LaQrQrrD1AUuHDMO5I4QR1DtMQgKdg7tSTAk6UVVLa01nft96alNuDQkumiM/kw
/Ie7N65OTF4dHIccM3q8+GIoAkONCwXCjZTEk16uySaaXLb14AJPSmN3OMHzkYsD
qlfYF2JtNNNJQ+okMkFZDSHsWQMBlQndzOudvtfF/cRVR1jEFALSSRwRwy7i3YYD
/wW+wmKaVbpUnWv3isUfByPrP+k6riSPGey7vd+ZTSdek79heqlrqQ4xMqgbSpig
KfVuz8UNolY72lZ+Q1jT8aDwlAGA+2jFL+rbZKu88T3/LZWHg+HhQFoIsVtuw56P
0r5cORCL3VjVne6ZQd5p4c9aMsarSRoijdUp31EV7CD8/RQQKzHMnx2G9nmrmSkz
PGleDXsmUzQ35edb8xBCTQ7iuKFmrptHQvNYWOtsLFKO0hcW9OvThSMt5UkSgxAU
FmQmqzJJo5ycE3a9WPihqZhKdBP32ijnai3IP+E+QuMwKVXtsw5DGelsJMBLoi/R
EM2aPIKMXDZDsJryjUzeb/jH/mJnOvOZ0R9pmeMvgzmeeqkqVdLtyorLeXSxT4ua
LvcYEwHB/YpNi4iujaxewApWnTa6jxBksiZsQmxyBPAPXKNRfLcGbI5ALBo5aRAo
W/CXVBLf8hjiXDvc8CinMAV3YTjAfXHEU4cKsPci3Iu833cd10YZr8yG+J7gsI+m
hm7oBzFBeJMvnJwT6KxIpZd/SEfapOtPPm5wwczPwwrLp7G0tayP4arh+CG0WV9j
mYH5CQymLrSVmqX3NFAAuwXKuZHM/RiGBolYG4IOrOfBP9iOqn9eEshzTBWdIP7M
musKNna/f2JbuFjOwwLDbw+LZytj2NQHbGwNUT4u4vpWkTIrOkZi/O9AXXAaUxbN
LmEBTJvoULQFbnVBoZSsqRPwDOLnNXCVjVd/CiolSrFbYLJzoTZfzqjGmH0Fkrhj
E9dnlV1eIspOkhQMvSsSwMBryh7m9HUoY0yvF25Gh1J4rbFWqhRtx9EOPh9/vtlm
z4LTu8NqJC8OP90dOVHFZKfFOZmSmPKNlOV9kRns1Q2axoWsnXoT27H0toVIc8m5
PwDYTxn0i5820QZbEGlARtG2HlUxikxV68dIfVnpdWe76sVmUSlYUXcIernDLqGt
oYS/v/S4lt7faTISDhXDgUZCCiEsvd5tjb7O/ZvFS6i6cTk+duxGXs4IdqRgmWLZ
t7k0DAX9iiKFLj63syLr0aUaz1b7lzxoClXlaMhbIpnJBlbtaF/oxfVjmz9OROF2
yE8cxHdQxaxm44SpMVjMBsXgV1c7jljUykmylEbKab6Gra1jTJvyQPXDfWSsurBI
so7JaihvDEWXUJiOJACDWUxpzvhzhYkyRWmw9MlWdCw8AG09eT1jN8UaJ1iH22im
s8f6/yhNT0xXqsIvfpja4TfVCDNDhrW6q8pmQWBVMULrUIlWtTZNeNc2SbjSZQiI
Z4hG6BFFuYO1i1hpE97UCD5YE92ICbtN7B8RGNYU0YYvhguO77kiAFnHzPKqD3DB
a7hSlnAkVvkiYQ9I2bkus9e4T5WJy//8K6rPz14LokiL1+g0OB2cccVeJOCkjhIN
/HBNuWr6zdRW8tqMsid1+Up7kwkVXqCsbQScQuE1DNS1fKFsY7TyCLF0kgeTdzz2
kvqpGE3cipxMLH4hDi9D5yqU8QTy7nORxilr5zZrBYSRcUdLGRc4SKU/O2sztm7I
JQiingnPIpazXQCYlfvnRhHUkd9L8ef8PnjPwqZsZfX2f97ocoOFpWfu1okDgKA1
I0YL19IH5tfccmhzAcIBWVTzvcRSmN4ux/rljtTNsyzlG412eX+WF7HgR8mBxEAN
/ZEL6DkF4lp601nn9/knSpEu0r4kPPLa8KwbZ/DoOaSB9OLWiEjKBBM9K7prwAMV
IuqX7Jsfzr9z4gNhdrGlWapZ0dP8u1RxXK0OhLQ8MoL3KSRfYoGs+A40yKxceaSJ
X0hPPcv8ni5xkSMSV2V3tdRiqTnRGgHFDwUzKxvMagkOl6mcaJbMpOc9AlXwZJT0
0XzgBIQOTq+U9oZT8QQiY4mimD3i3hYvQy+no78A88g3Xbyl1qWBzPOzb/GRhGlD
wA4um9DUqQd/nM7zetz3DrSL9gEcLf+dph1XmIBFdSv5HExspT7oVdYJAnZPDCgl
RKZB9MrtfYFqpdgHJC83lXVArdWSGiH1ge8GjBJK5OOFEi7eOzmm3/TMwIgip/P8
0aTPr/h93ev54aEnvshWkYWwdydvegp5jcKxVhfDaeCna4Qh93NBZYtDSubyOS3m
gdb1Yr/sZ8qjY27p4LvCOMwkhDephPE3SrYfTPC9XIhd8l0nlBp6GqJUKeyN7jbk
JXXSKM0xJ/k1HVWe7b0WTRgA9nR3AL127EInIzA8uRHSy0rSgp/+ez1C2UXjsV2U
vhl9ZmgQEaimAvUb1Ij6HxTon22WOoFPg8ZbUaArYuavWa34yOMVsMqluc3KYpMR
c0t2vi4zrsY6ykFMKKl6/27tuEBMXzOGgAw/I+y36c2XGt/SiP9edX6omf/X970k
ew1S0W9y4h1Fs7Mwt/kEEVHMw0kZnlmlRfbDWLzPOfeBjqApYiWMmRjQqVnyL1GF
SBCVh/kv+1R/i1PAg7IWGWt2oB0jA03BwPAR8zyGg8RYpMU25nC0B+CzlITW1Vos
u2L5rKDv+H+iFiO5ZPTkplDUPzZcX+1HMb3NIm5xVvbw4fIzokSulDLEtZkO6owX
4MnaVCJnypuN1bGln7gIGAZX7RK1iSvYNsmStYFZgVMjioaYft+X1TWfnsts3HGO
WMZzVahFjsxBons7EMYtc5Y08yP4CITdFpGW4jPmDn0KHEdLSpJLXUfMVmrK+7eO
YxybZz4rhJPhYmrArae4a2kK6UI7oUM5KnjnZBcoXB9xIKMXp1OEEE6XZfTuxbjy
iQTNFQnsBXXlOMHKkPbgwa8Xvr9RniWxlOdGtfIATgU8CVVcI1oqU3ZFWDrsPlfB
KN6L2+spRaFb7Mjb134w8kpBRATNfCddMx3A12Qo0QQ+A6E9EbxzLuFhfQy56DKM
gkNmZmTrG6EqTucRY+dmB0AIVqDXSzlyVXadIe2h5XhpfvMs8NMZgGRt4CJtq6Cj
FY6bDY3G6gcE4bzQ4ZbSSv2POVSX5C1cCABH+crHkMezm55avUh0k7YIIlItvdlz
pAoO/FkAmnq1VCvHy5TTuT2MNZjX1wTfubX94+MfZDt3yWfbBFhfnY41NJrHft3p
8hql267ZB7ec0kXRjzvl3PR5HSOfuPxAEmL24YOtpdzmXZL1bNjjVyIrWwbR8XdC
aQBDhNx2QgrZjjMfERHZ9fmc3xzSRKkqz8eE5tBPzBx24fMs99jjDWs6O4Qvx2N3
2xKcsNtCV83OA80ye4+Vyq+jDst1xGIWqSgZi26A0ht5puXl4SwxeJn64oQqu58z
UYnk5ogrE3AWDUJQiSirnTxfULtZyRdduVQvN49wkigPvE4lNMidSmte8cLFFGil
dqtLS3Bmy0qTbe4Y6+zfMLdKbQEMqQ1veV5JWs8L3E+cBQioIZr6DVe6SSgr4OMa
Z9TDO+5edqDepjlziz5Jm4Jb3jpQLFDqkIPtP5WaA56tZN5EEPFvursbd9jDAnKA
nLliKlXGj1MvLBa0Xlzygip6ofV/9GCEpsS4nuv6TcQFSBxePYpgsCVUE3a53h7v
JhL6YIP80g7Rj5XEPFPhawDd19vVUJbXAhUNgbC6Svb+l9L1EN7GBYl8VuCfzEEJ
Ywxbm/hB8AVfSl5sMfy1cjX8ELPZSBcd9GI9bNqwnqCBzHdyApwog8FqvUKt+1lZ
wcOs83TOH2RO+5XUiwjWc9b7BCTq2sxtnc+1+3kotT42WnRIA23sVCRlC1WhaLIs
Y8Qh4UmSyA7h/16JUhMHxPPJro1igjhmcCytrA6nSJxf/skSTh8Q2C8KX86HgMFk
o9XsJYhZqOkudhSvAx7lxgxQdUQlA6weAF/C6g+ceF+B5CVJ4ktroAD+Qaqv2Fmz
JKW0yThUsl6YyYoYHtmDkcgpidDFoqG8nmxiWSoaGqvhF2CjfsYNLM0DFSdxm9DY
o02CCmqgU6XPvrK6+IPOSftMbSIQu3eSsVrjoStb13KUGdzTmlVCkiflDjQuRCQo
vqfgFc93XM/Ryf8QBdMrnbv4mbH0ng4vFk1GM1g2B8uwAlG0ae1qP3sZCizin7WC
IpQFT3NmDXiEqKbLuD/ilMk+MXG6Ui4FQBYMqgnGrnCT0BHh0VpuaU0vT1t9ZZm5
oZUFmsrqB27SyDkHac4FARgez/R4RVDbM40U3hkmHKvFVaRKKR/s0uoMhmYiKBxK
fPZ0pD57s7RJ06UKK3n3QWK2RSyMF/6oWclbg2jEakeCDnVASd3RQ9+9lr65L3Ec
iyw3dMQYAPttgXjqje6DgX4+FqtoyK8b/ohobagjFOpiTVFS4y3F4xH0oFe8HOsH
+8oYQqWEc06Xu12XN8cn8fY9xsojB+h4hOpn/w9PCUjmTZ6Wu8U0EziFXYIG1bQf
jvGVjJlvG/ntUP2nTFj5kRkGqWWbC/iNLeUccOM3q5MaDHFYpbEZ0o2VHIwYu2uA
/PrXzKcEfg0xL+lFPGvFZ+DKukMsJBrel7zzBlo8C6rQEenzKmM+o2m6yMKnYPEH
JyY3o7OzQ0iFbnqwrZtVYln00nqjdYGvV85vAsdjIJKlWROLsLok3GByGiGS5t8r
RvoHCTxlMMTX2JVVGx+UR3HmpTj3+/HgdVS2Y7wtdXO+i9ZTjBgOwwrGIRiYEt/2
6s1PLk4ACqNqsEreCko7wBt2DBG23dSVF8AS7caWReohgPa67IIPGN5c5GLFl/fz
sPHg7jJ73VKsnd3spWY4GAjcINwy1oAeVy8BDuO3KFTPh254k7qd6qvsveAaSoYf
ry1rKcYYICTMmf433s0sSYQ0idpdtQFtHDsS+m/lqHmNbOEzpJYFlfL+YtgFPD5F
eSDDFnBwV42yTDwcWo/E9ZAMlYJ8wbgD0t3q6gLOvd6fwgdeX4kUOBvceImAKeuw
t2jO98uYQAiVJoLlLgqFtFiYcKu3KRckwptpVo5jCNi9GI/DzCqtpYNukCYvJAEY
zPPxJGEimrGbclK3rpdtvBbpnPojJiU3ic4sHJ0wbAbjASxuKijHw/SbuLX4pOqs
nrJM7gr+yBqVIGS3SbKwXz6vGdssSAgrU7Fo3Q103nZqsjkKIZTYKqEP3xZhIuBq
FZ/xOdv1t4K6YPPSbo8NjUi9qgeEpCN2svBEn4HRWRid6G8izsT/1vvm4FwKof6R
9foafBIGgivkJVlTxuQcAz86Fulj6BuyGkuEpFvqnWyOT/zoih6k3ySEputwm4i5
ttkBWoQbt4DhhJ1dN6mWhR2Gl8pf1lhDtb82E+i0uWly7M18rC1ozqYFFxjg10zv
AhQds0d97yoIfWvVSrLD5pX8dIxVG6bjYRxAplmjmx0q0JNkwe8oFzqftYKo1TzC
HMbd3TXhsD1kAIqRHhRciNXG2Sw9L9rawpUuMpIHt4ftntns1+Ql57IhuMBUA9Xg
cLARvyWaHkHHuy+YG9vjy97uLuJF9e87ZGsjnaoYD9stgjTBiitaZXbP5h3chNWH
5PGta7ESD474uBIDy25JsfgR41preZ2hTpd8gvt9ZTyJc2FIzLUr73JjnvB6QM9i
rYBomSh9hHkJBik6BFN2sFtdJv3jnAEClt6KGgNuwJOQupys457BeReQNrHjusiI
xpoPPKRx+mH8Tc1MwdMU9IS1mDtiuhWQ4QVIWbnUL6RmUCra5ub1ZoI1R/+e9Xnr
j5tZoe1bu25EQw1U38e6MShPaFQN0eJ5x71ycj/q7UI9cF58dcpjh4EijYBrLQuz
H1Zo8/9luFMrgZ023sTN7OK939GUOkB4VZOZbxLgQ33B92uRadyLjlIeQw2TLJt5
MezlHx10aKUy/sjf3dMifpuQ7S6mwekL2hkyWkeB04ty1g/hLdkpHBLPJnNoVUpS
flmssRXCFpDLT/Bp3G8FVVgXJ4YzVW697EdNL1FosnmK4DlLm5WrpqNHNun/n1hq
UA1vBFouggwfhOHtHp5WuT+bOIfkRZM1hw880EgF9s185y3g4XSJZc+SIX9YLBRQ
N/diX9QAx0GyTGDWIr53M1k9+NbWMJm6YUXIpVOYcQcMuo02OjN4nkzL0Mtd1hw9
9FqCa+Dq0/yhn9ccuIO9LwyL1u9+dNaqisPO4lT0Q8moaAWM6KY47WZ4vPtlaxkt
UUo4LaEzZNtPEt2pTKdbV/qNASNgisGrPugv4u255dvIYUjJrm6JNHiZdd7SP/Ty
7d0oCbKokNMOtRUHq9PE0OjH03N3uXJ+S6nUYgJHrXNxcQt2tXRH28CVfOVFlcyN
lxZ0p5N1ShKEvy0w8DBIDBWaRM0E5Ie+IYi5vkmLnPecPK81l3n1QJOZZy742Unk
aPTPnbceeXgYxVi1PN3C3rQia/4XJBibPjuxqaMBHgbXPbYIZtFCr8BAi8CqDU3/
1w9x15SBpya4x2jOKvT3upiSDdvNYLEsyeF7zjfgqpMHeOd+DkXV48TnEAoFoRn8
scsdWL8JK3TbnG+rFyJj79xMB2M9xtzBdDYT4ztGcS2GvDm4IY6Tgj7s+RSovZd9
KZr42yCgVUYCdAT8XF9IrKjNbaIokgRU8PcRfx/EXRVEoABq1TCxNqz6q2f0rU8p
Stmjnx8aJ0HNzlpiAKcSyvC/GrkalZMrc8pmLsNMeA/RwiWdF5hbTNDt5ZdDf5Fm
Qh9qKIAcathd0H1AEE21Lg+wZUmJACo2om51geI/CKUl93pp2uot0w89Ipf/ShgE
mZAu7k4yow8UJML5smbB0/xive5scbrX4BJDKEEhOVXAIWjkvVwbCSYEg9Dm0RtB
JLbxgZkkzLYzTxlW6K938K7krQfBfE28KdeTOY9LeWGRvs1xx1lOsJEf0SF1zC8l
PeyHYcv5XRzmA6uHN+2tfa0ukK9ww22DJ01QPECHEHWmREFcCPSG20o8S8HJT/A+
3nQZdaOjfejr3VVtGjGtMKzugibV9sOwib51284opJsFneh/1Qf9wc2VNP0V9ogq
OMP70b+YvdLi01UdIIhm+bjtf4MzOjzwD95jegke9s3KWuFkzWxlGz5/AzWGR4SN
iNCIuLa3HbbJwFjYjYVZRP26YdVlaZeXSO57iSu5Gaj09rJSL936VoqZb/yCvsx7
lkIxbwr9bsigdnqBF/OGz0tGPxhVquyW0tD5Uvn0QK66Jv+3mKR5Y5p6UcY3zkl0
SPAgRmYYCqFnZZBbnP1PEWafCIRDRqyqjaXaDDpeT30S/w6bCT7uzhV/e7WOM4Lh
GhzcYF8YYqq1qnfAPioU16ax/V414YVZDPb1xZh0z1wIpUetnx5itLjHxQn/9QoH
HVD4dZ91f9IPaPFfb84ZDjJjgKFwIgQ+3dWKyDNZgH6AoZwgl3QDGKROZ0ZvdHC+
Q3+SEqvARZQ+Xw2kYIb1O2gAkMaISAnHl0Rh0Kvsn2o3B1L7OW08aFNxpoWQg5YT
NlkLtZ50NkeoepjBG2AcL5omClelQbJJYfdx28tI4r33CJaQQRLodpqk9Su9V80b
b1EjiPPUu+nzdzo5f/S5BiUxaPQhIe2ILUQo9OuJAdXf8DlzfDCG/9rgp9Ia4xV/
G5/8kYVqg1hzHdgTo9pbt0XJuzz6qaqsF1CLC6JtNznQ9fSmyYdMI9tVWgGsI/b1
iGgqYE2lwtbyLu2GXwzNcFIJNkc1CFCUQtrquF1xU01sW5gyL0VTBxjfQ8BjHZ2Z
udAKVvFgoW3CVFalEFAqo6MDwsV+HHojYftmsJxqw/bknhxbyLbv5qRDhqfFt++W
95MLLbDo+0Xxc1oVffUjeofD0I5Py/wnd/OcbFuxdB482BFBbBk9KuPxfJHoH1Sk
5Sl/w6tXsJkF3rjIcO7o8NTr/Lp9UGP+dzMSnPif/rPaIsbenerOPAc918+AOB48
O1KS+ji89quM5+3+7OJDsv/QhoGONaTnV6ZfVCMjYf1biuGAMQZ3ei4FFf3mWVWv
4NDCgYeylDKQLvWYt5RUfrjOkio5zjTqMOOJKfljKp+bQ0vg1Rig5KKjJBBKfTbK
FtMbAkzBXPIaH03bBS0Z+0WsTp7DCjsMPSqagAOY2S+CbwGk3YjylbeM84J4FuC+
W0jxvJtBQIs+JXxnxCnV2i6qI2MKgRJJsGIOxlSiIGdD8hRM3VZHcDRYGzXH0MXO
8u6khidQ3he28AVVxsFbmvf8rI7JNCJIu6ql1kAjZqWS9z1wTWw6n+w73epEGsg+
OqzFzvbCH3Uvha1KNw1np91xmc6mP0eO0HqL9WFKJ4SNvnaaQG4mEpVPKoWraYtD
8eQcu1w71X3uB7u9shWRMpJTqWjHGrPUDZTzbzzOKKPNSRAK+tyxnvUu7yrvowWY
DPxL9vYjvr6fO491wll4rBAVCy2a1wIhmpoxlDegQXTw5HbMsn+w1DmQy7hCqf1l
9nV64Qb7HfMybPN8v07qN85un7MRZgyPDjAbAzdRe0wdLH57yt/WXJN30ajHL4N0
zRW8u6MZDj01GXcA/mv6gx6TUbCsxtZ87S1aKrJi8Z5KRdT9y8AVixviiA3q/XOK
nWnEEY/2LGgjg+kNl7zgS69HRGXtOnbKEHptTIwcqlaxrGDh8Trt1lHCz0dH1dTU
RTRL5Yi8ntZWzjHplShcamXNi1/NpeaXov2t6tQhv0RhzsgHpMjP61cxgDcz+YkA
Rcc7jKSCa0jY6jTkt/AnkSbfkWpxL1T62CGUJC2VDwhzMhuf47In8UYUsfu5ki4F
EqETtCHh0A8SMIfVqQRGUXAVG18dTFkPDmTB7HTU22XDBd838uL18xXXgBdrgrnq
49owP0rfB7m9IoT5qCQqsbw092LB6voiBo5vr3IHeCIVOn088C557FBix7+PHuIX
SSF80nt/bt/ISsnB8Q7+tu7p4+o7rW5zG26dFMTzAYedEsldLLY0GO/2kfz2K0fj
0gTS4dJBH/ejoPUqY2S9g+YjKxUcFUxjo5wyQ+6uXrQW1x5hcQJg2wgEEJxkGvrG
Nzd48KUNyRIueFKacQkoWOXQrjoLjBwJxKG+xzvNpNGqtxc1K+hmIiy7974tsdim
A5B5c+wnRa/gR4xX4hAHls39Xt6k4iYkN88/xiNIvFvSNAebMYvlrz7OAsif//8w
/nI5tcqdlfPeQlb0kGnCNZJSoJvhAR720bdw8XAdXa+4yA3HgCCKiEe3UyJbBQCs
nvU202pMFdqMWA8WAYgYyQvfnrj3BYDo78z6xQL8/ZTWO/1yEoqPv4B0PEHxoaaP
V1ecTMQW9U+BAWUjQxO87i9n+PBRNgedpmTpnd+d9C9/Azz44CTLQoMMGaNDTi5I
CGn92tINm2sueETGyxN2ohVpNzRGqAMTCCip6c9AtNBDHVdZO7JnA/FD2xGLUVxH
HaQLmFvr9SopUCHALEjFMSKhVJ7xtY94rU//f3WHthbvQcv2YP2xb7cmZW8LkaNC
i1Qps2FwJHMD6BVD2yiFO1V98CCf7zsWILDN787a6U43wvFRGijxNavjjT9cJE26
mqMK4qQBtK/2zH8Pj6WdhPt4w/YG1d4otZkXp98v2qzyLzpSlbtwgvw12PiZsnmb
H30F0PrNgxifiaSAMxMkDcAXRcZheS+d2HQ/3V3gAWkw1RL3wGbvlouHiqabnauT
UAu0xvXrGAcLlg5sl7FSgpR5smOR4xgInKEBHt0Lc2TadpSB5cJP6V9Q/xAly64Z
WkAjlTER9nRKK/ObPfOuJncYmP4aNc098yLdNlpogeiv1Wej6ZnNxmIgPAoooWb/
3hwNrxOQMm3e8WbbV1yNxEnT/ChQp2SNg+rOm+ja7PobXxVnfp/7pPFnu0uff9IX
XVxpf6JpxXpkHMofYrnPLBltoeQp74zBy+5EJLk+nbvgxJ09L5AGa8p9EbzYFnRw
mYZ4mZF4B5bDjz120rHTmPSacFs/1Ayx9IjCxagW8W5a1cZNm3XvB2sr7rui2Ayo
fEizxMe3c36QYmoJ51gMVMvwNEo/hiV+YJRPJaTFVzFma5fkLoS8nPme6CvcaDtx
nG8uSurSpyacsTtxRaXrjxHl+28PQUH6ykdZzAmdtJomQtW58+U3NVXWSlUrTEFZ
1kYQnN40txbz3gJOuwADHUC8wjVP7faQMnczUuz4XBqGXJc7HyfuT1OCYnA/M7by
cQ6lN9vlHW4FhonpcVgwxnzBuksnXZaMHZmepQuLs8cdV01HSF373tMgo/Ykgr3h
SkBcbupapRXaOJEJv59VmpX3Hb8voU4ALI3QQMh3BawcCqjVTXwYr1X/85t5sfwn
H8otiNlIkvt9GNiOeDygMOCUhrhEPtuc018KZk/l1n/yjx/hI1UafVVK6oWn4IkY
hs/Keoxxfo7l/UVHHDmTV0Ozvtz79NvkP13HblH63wS+VaXxoI4Gv+cSLaP4Ihi0
s3BiJLQDLmMFdftGNZHjmF9lh0oMdQWj1px86wmGiMCBHK8BxQt/5kVKH9tybIV7
y2SDmwLcW9kb0td/6yGZj/VxCPrU2JV78Mpx0SRKBgiHf3Ggd9QFJqo//c1dgfPn
WVGeDTqvLUs7btnWayYXJAS7Mxh7NqMuST8m5+SK7t8s2TrywLDzBdTgkrb1DUqf
OBFYcvHFj7VmK8nTGdCV0FxruYkojmKLs7R7ltr9yPSaOiFjtqeSGv14HT/d/1Yu
Xo8tmUtpm0av5EtqnIc4sC77aAj6R0h3j3HBa66BhPfUOuXhkaGztpqe/JsY560H
EiStCjTdyfABe0J0mmprjJ3grbNrEil2dZjO2xf3QOFFfBkoWAybMJhXzd5ACerM
sF01AClaFPyXFt3xbZsLiMJ+kbQRRUzXUONWTGw5qOqClNjuAB3XFDfxwKGHxLgt
0+qLFBh8PLio+lwbvMx3qT8aCqW78rmabbZaMaTfcCYoSWYFHqAij4eC0kigf8tB
EFMWxyE/FWshTQdeblfNDygKWT+/snp8Dn5oBZOixTZ1N9Oh6X8q8IgazFwHmKQq
jg55NHNId78PvGnwh+4KPApozsoj1DS7cxXmL8n5917oklhvTGAj+gaYAQjdbLka
I+2rm8ISWye9k5N0R4amGUBoZl8oXYE/lfYjr/z4qXjUMgOMNe381lLmI0eptF7o
g5ewvVMlaltH9mH18ZbCfEuewmulqguic0QWyJF9pN3RwR8hGPFg01YNeA2Wi6lD
M06/aChrsBEOJ9qLLpiAWdomvmiVht+2TfY9HqYRlsysLR2grmN7MGQHb1zBJN4W
h7664GuFc5PnM2UUInN7YKPEDPwOWmXZVy67eoLRJJ9GQ4RsdQc2xBce9590HBlw
p8Gh4cG1PtizKUzAcZ4bilXFQf/GLkpx0AJJrZuV5H4yqWdfi0psOjIpB53SEEnh
9NnpK2KXb5R1fPRJX3/gaB8/oX7VNMIw1QeL5TRRMcKv9C3A+mPpzuxNwHHx9Vu0
FvM/nj6LPt78c6DUKLOX9uUH6b++vg5hfdiH9T4rjyiXnQz5aLb9N2e+3A1EmnLg
BA3BmfGFczbnK4egkAVo2PPSI1UdF64mIzdo/2IQ3FeLkQZFFbUmKIljkQtCTNts
LMvfCAtn8NM3i/lxj4vBs55q1JjGDabumZe/uUJvPeLmPFwt8xo1/heYs36ECUhq
5kRoaPehez3z186C0UI/SUQ28KHjN/qJsHTIDUXmLcemkJFPDNOURSirPFzfDGr2
EBEmgZN0hGaeYxWD2ivR8gvMTrVCdiSiCaGuVCj1w8WqEERLqeE/2TrdGos4JsVc
t9flg80aYmBGVpibKzz76ckK96bForNQLVoJ70JVMbNeZXrWkN2rbI9QgwI9SICk
MP1Fflx+ZhCr/AIV+p3WPafp19m6JLmBfL1fytKUluSbMUM0B6C3it4mP3VhY9Xq
HUujKVIPsLd15lrGYhVH5ev+4rkBAQ/Y+VtSFawmn8ZpM68f64/gNP3HZ/iSHsd3
JjiZhKJA+dVo2aJwzde0EAlOzijqh5uvjPIkvjzeu9S2UeYR/YMfyPsPnoZCIfUk
s3FivH47AJ3DshuWqyahinrGjCVDNpoPcKH+cVAczoFn0sB2E4nMeMNcLXgh0bBt
RcQigNsTJ4Wk7RllItxL9x32HN50NaODFJ9mQ5j37X5/ekb0O3s94NhYxzBZLJ1v
EhK8SFu5Pybs0wZOlpdrlRNbx54cFR64EYlyDOr/VeoDQA81KAV1TapQpIYxnnPZ
KekbKGlaCtTS7VZRVPBjLPD9ZL9lIQ/5B5r4oN6QQAxBTEwdDF9f6pIWrkiyAnyi
50Dr8zCys7iSfJmhX4O3KKSZSpWRt4CCBu/Y8upITlMLlKHzt9Lu00qSazow44Uo
vpCCS1i2to/CAgtnyV0z00BejYwPRIlxO/awIvXd+rexcVmv1Xrw1VIRUUmawObm
gK8N5oYB0l/BMaCGQ3XfMWnbXWuK7l/IYuW1cRnumN09jUpjBKExgF9AZwFcEvQq
PAEG/0M3q3V0US4oc4KM76VYfRI566EhlklwlpwfmWYHs/uWQWtgRjkJl65NCY1o
CZ9/GKTapJSZmPGQNqcvHTiAY+NAgZCBZkzcC9H/Wl59Qb2Y6c0/urNdulnEw0UF
WeVHsWpaGD+de1WKwa1MMRH4Zj1qC54v9ZH8nOhke9d4apIuDXp7DEC/cJNZEyfm
YpV7m6/lTpRkdISCYMgFL6B1Jf6pdRANR6AAGyg5Oztpd2bKT9zNwccQhasOwPSm
frvL6d0aNv1dbOLniNu9BpQ3GPT/OOuxlbjOxVGfRVe+yBfkReW8D/HR8T2v7MEi
Re/bsu5fTPbata5lgQ+9vmzJFoikEajl8mJshXeP9wp7C3/yVJlexzVkswbWoVXD
plid7iNXqP9LHwworoZz16B3Hz4zbQ0S+2pvGhiDbibiJC+i+Z+ZUyYGr0UVvsqB
RAotq8jmQT9PWCPxmpvqLK3mz4Kz7m7MDPov975cCtgAmmlmv4H7hbWdAByVafVG
IU+rtvMWYAKDuSZwNMGpV/K2K4CNdO6pV/HPC8+bdt+gEXOc9Wv+aCcs3X7SlAmg
k/M4sJ3mzXj8gjfpz3Qz/+yYyXtV3xiyC6oFteXwJ8yLuqWKYAA5esKn8EfAqOBu
AWueOD9Fu3ZBTCO+XEDov4ApA6/68PHAHKKM0ca0cF2Ri6JDJ5/lNTQ8CHzKeLLn
qnQ0NoE+baW7Hw3+NdKDhyiX+khjOm1ePBgi/OyFBa1Y0wOd+0M2WbafSFzTqGEY
tQm/dCiZcAP09oJNd6EXJzY0PfO75pY7AmlLXCcyILbS4bvkgiOV4JChnjaP4RwE
KRavO/xsGbchs9k82VEnQWxBWIvO7WKw4bEX9XeL9Bi4aAdX0mlzrRqAnu/pj9+u
TJ4fTTf7VRrTAkOMTdi8y53PCtTAnrCFNfMBTSaNjc7+pFNtd69qimNemYv0GEkG
hl8dUGXgctu9k2qzR3PfC2fQvqGhrY5x9z0oY7NEEXTgtYe5FIKtbjdvXB4RbxR7
VFAWH4GZypDLN1a5CjO2vTuyCJ0zwkEE2AAzaaYtOpFpgfD9rEJMginl9dLRPvap
UQUVBOBNdOfTE3KIMrD++LzsEyx+Qm19f0uzXQUTsuVrjF3vhjoslO/qBjBaUtUe
7dd8O1Q1AEUIacwp+7wYaAfgRlGGihlKapEi4n3m7ssh3hYF5NGc3PzNbO6j+Agr
+KfqJ6c5YFFfu5tOo0j9smAuFSg0EE9W6Z+RdTConnSId/Cu5dPocC27/JMjSi5S
KIgpCVMqA2ouv3mXVLqxSqShzr8RBIF6WUF1GtZzEYXtWKl/1UfPNFUQPCSafCG+
PpNRZld/JMI1FxvpRgXU+moBf8HO7u1vug6NwfyLPMCbjLNCORbAPnXvM18MIQWe
jfINsevA6DsiQsvltjMGeVJERl36NwPvax0v5t5SOL+TjQZK0Df9jHcpxA+UcpUd
o75vEY/+Yv0ww6NFhF7SMzAqFJgS4lzw5uMBWxCVDmCo0Tjd1IJtllVjNcnNv89W
0wfBdjM0XPacNC5/gOt1Jnkf+xtZPta4x1HnGx0MW0JZp7Tpdr1HLggX7k/5pbzU
eD4CL0XGsAf15xgoqJhQ1bNimXCLYhaCKfWUvxeBHkqXwzjYgi1rseWxVa2PPfar
dK267LlXe949BI0Cqay0o8KAlbkiZbNrv5quw9irzwvGVMMezbjaHfTMRcjMiNsT
0gDvxUOMpUpsQmHwyJXlexTz8AYNMsFvPhOUUFSQTKIEsU/OEd+tOuIfYxg1r0RC
4+IY3UXNz34gPE6W8x2NMMlGypRivg3KP+KoNAZpST8pcEom5TkpdDHNV9cj1geF
O6tLLOczDKLBsIKz8aakodjb/ZHkJULQYBKSC/apiVkgQI2tH1jOSfONnRjZ6UhD
ikedcPtikHXkmt3jL/OLu3Yn9XNx5dZR8Ug0NMtrCyC5QE4o0wHqBSRKYheOnfer
8lWBWe2Z1MkoIgY8LNM4qPSvb4PWwUtZagXi+eeOy/hz/B9kD/JvIqVWZc7qYdG5
ujfSutOHK34wzGgT9aCkvaHDy+b3KvAkhgLrfi7Q0Y/IrlZ+B1G85Y5U5rWDLiro
zqF7xn2yOpgTZ9+1IraTe9kguNDiz+9n62LN9WxRrv4tfV5bfA6Mo1Z6d8Wom/Pb
8YVHM6cOyktv2VMUyedPHBdifr2p5bMqH5ussNNNBFYDoegEAUh4aVvQMvZw+F7K
QHNk40Y5yhP+xltRZlrE6jNO0bniujEhz7j7qPNqFpq9Moj5nUN7mns6IjuE+ObM
FhSSH2tj54q4I/twj49QZaTzBz2O2vcTnZzCD5cPwQWhi1uOwGlr1+IsCLkrHarL
P7GfZbyay8QH1zOf7mzQ7os0h4M91rvt41Sx42uNK1fQ8e7AtZjkmVYvqWYSeRsO
RA/7FnJI3Rdc/K5TMD0RxAN83RTwG9ZZPpr8FLNf7UWOw4q6L1CVH05OxRFydvRQ
vpCfpbpvtQ887unOdkxxf+N6954fEAmvOpaAwNM4mrmHIeMSjHl5n/NSrdFd/OU/
Y5/iuif35vbel+ts+9G53MOE7r+CANFoPYRZDbRkRFZtEaMCR7FHTLy+eRdd0MDr
LQiNpMQBbRp5XpO9Fua+Jbghcn9Cu7qEzGQwWqL8OlQWbYJBFSIagzV0Q5ZeOvVR
VieYhM1WuyehM2I/3NcG34YbGktXIvZOQ4m8PCpu8D1nOM8Mn0pOMT4H4pa1U6zo
bNTNELwgHdJ6s0HlepVgECEQTclpEJy+CfjIsvDp4cpecLYMr8pjmxh7DcwCuKT8
wTXiydbyHauZTRpY5GyMgMQeLN2zPrRI+qS6zocgJwxDTQXT7DtjNA1PDtJ6RwvU
LLLg5TKtVKE5ktufEwxa/gR22TF4kJKQALbk6iQQ69L/l7R1aE/6uIAc7sWRgOBs
0c5lIwlMbHtWkKIC7MO773W1I+swOTAU2faEFImloQLatjVR5naOZQowoIlbx6Nk
nqvNBgStv+c0I24WK4HmBr7awUmSHIqUiGCVDLmTUYc6kVzoDy7BSxcQbJtUFwiO
c8VaiALVJ6zC1QZyMSTwqTXcz+PZNWLeYai+58UFstn2cUBMpE+OE7I8ocnMMhTt
1XUFUjW3cGhF40qED4XHlDQAVu6UvsdRdkLTvPp6uvMM1DHbEXzStyKL/l5JG9iy
01ZIlyKSOmDPK78NlUrQiiJXhtOnLFmEcB8omhfIbuOXsyp45O48YucYhotKNaty
twahOlY/eU2SMN0kM4Px/f+uyL2fFxonBy+3XMSOa8mmvLAzVWqyAKrFc5i0jPFm
pFGMlbhaghnmOpZ/8MxopCQ86AbSq4AgFfYryZY+kJW001jiLs/ucILvou8UNVrU
TSC8TKI/BgSwOStAHGJVrERMgsALrONTZhGhIN+4TelOfW/6rHi4Stow93LK2C44
S2ph34o9oMO3LYRN9sf+Q2DSnPGEJ2XDXSSTfvdELArcpXgf7io/pCUnyMGmKAJM
TyxjG6yYFwZ65CyE+tFgS12wA87P9uF3qzZekVNbxJlF73w3O4redG7Gz04xGvvp
MJdq0iijl1DCbwp2DRiMj48hUHg5cJhDWdPQWLnhGA/BMM30/CX8jNlH5Zvj9F5E
aaf4IbawWyVNO+nAIx4UvnmoAwHkNR4HK6gB3L06RBT6YAtbFIUrbCDxxj1e/pCU
xQfLbCWyFr6f7LyqhScnO0n9QEIz7ftCbDyRFEt8xPPqBw2VKg5kpW4/BOmoQ4dn
0JqsxeedHtyC9DXcen/EF4GF6UbrVAjsf8XHH3uFc105gKT6RncUlD+GvhSXlVXf
b0DXwPEKoG53J4SRa7K8OXV1a5INzr4aZO9id1U9YJAmWZKrN2rFq8LkzHYObQIH
3aXZMASR4vLIa++H1BZvS+j7v/1Lqv6evgGOHAEbjzYdAhi6unbVPRm1PBZwJaIN
gluK/8tA2wPn/guIu6RBI17lMYrKK+kcpT233vMNf1CvlgLCl33F+W9DHORpbVlG
Z7Ra3U0hcunH3CS8yt28/yMyGPhR8C+KvNqMQGcVYv02EKeg/XFGegCYRW4KlYvP
Ik4kp+O3YxJDERuR5Mc4/Y3hHz0ASVQBxiN+AooQ2WHnfyhj79jz0AAq3TV0VODx
3A/8pEG+lYbYOpT8QZajbNxtXgHJjDMaXAAgRxWaA4zUt17OUN+LShrDOx9ykGyM
JJvLFZJxzemcGZd0TQvwDgNbBP2X5hYOlDggJXRODvjCIpxJw+y32aRZCJNmjPDG
zpmuq3Kwm3NmFhI0zHcX78RC+yk1dEUUO68Uc7oemuI8NKgBcRkkWZ2FDpsjCWJU
yn6XKfl7J6tu14RI4jPx+seIsGcQafdxPUb2r08UZFjJpXKinof+DVKbv8xEGRxw
j2aYNDrszaKJr/iFWrkNBhkS/cwiBh4q5hxwj2qJPnPAiAV3ziuRcY652JeAGqc3
AZx+BbyREdFAXrPl0nU4C0GfLJqUox7x+CwvJcXeZuHBpeKR6vfKPLp4mQfks2OQ
Iziks7PdLZaru/VLLv0grNiH6yxBNx9LHps5y7p+BVnddBPd+t1ojAlNr+zjEeYA
wG8fmtzkJQfc9UNOBk/F1jdMRQJ2PFvUTxoMi832YQdEPFSXpOE2ytHFZMC6iGeO
8+GqoGvbX1rJl1oYET9hf2T7rLyVE8M9FJ9CUNHvq6O7R5JUgDjfljmhj+auf1R3
FjdRz9z5+WXN2/wLyKPRvh9jANJJfnvSS93bt5U5m4vk1fGJjJIb0/tzD1U6j3S8
38Z5qzvoKpphLNy5XhxMCbR5S5V9QucGlrSGX6tC80EqU7otSGZE980YVsrr7CuS
AM+BBp4d/B+PKSUcJty9LsGPGgmm3dMIjtGeuwurW8++5c6tWFVeVh/s2181GM0v
zyZE7pF2rw0reG0UvPMewuogcC7rNubeIEZlIVb15EJG6NlGITSRd1/X5Zd+F6Lk
agLvd17ZoyF/+TnC5aDQ3qMcd69mpE1fjH4aq+X0hxoK3SjpjL36oakyxdgw1AgB
HoRN5+VHTox8dxczgtd5yNglG6HjVTb8xvXkwkgLWstfm9k/+mLvbQT4wF7+IA8j
deLH1vatD2WvK0iUa+JEgjfu20cHqCCJ+PaSETZvovGFTbApHOiOzFHLeDqFq3z0
O007S8grat7AQnQwRGYP7TSpj2DvDpwsxaxkSuSrkr27w7LotyRKVMrSRtrJ5ne/
Swjfpe2T8pnPlRZN/+L/wtZ8urQly+2tojfgVlV9ZSj6zOEc/F/bnWOHPrD6vSvs
p6ZK1+KdJ7IhhWrXbGstOuqiyg/mAXfHRZN7jyP9LFDsutvqJK9EGZkOYMhtRgUz
0uDxeywwz4OEVor+ffyvN3DNgGRgv6bsAV5+idJVSisuOtxbSDy2VZdpwOVqPbl/
8JhAB928JDQ21sotLbnFDLgVbRs6ssoY+vw2yUG8d/UjNyoafVzcLoMQMsjGAsdq
g8cG9xgUeq4qAuck2yFFj6lL+Tp1eZkomgz2bC/ltBy08up06vhvM+cj8tgv2Nrt
i5DZd4z21tCrilbzBRA1lOhBOETFVdkcQvrWicSbYScuMD3VIQekt+jhYJAufp62
34uRHWvdrybJpdzFoJC5ELQC9+SXMWDueSSZsHEAuCHpoWdbJw8WsmC23RC2KFnr
hi021wxQZuZ9fKqz+qvEW6REQqblR4pbcR1sfGVssre5kSNtVCpA2ybVD3tXNWvL
vgmN0OWpiW3hV7CoflDjwGXXEIosfEIu9/D2hoKMv7EMS9QiWtG7wHcdycZUdmJk
JFauGfODIYWd0Mq6NfKIiEruxKvWUNwehohgHDRrSRWriGZr8L1a8/2p+MKjw5HU
lNqP51Fv3gTdomKxzshsi6p5b9rQ2+qXEyB+QVKZ4oJbQAVH2dNg7aq2kQoRqBnR
TCNFmtuFswijIab7NUEOKDcXRZqVkX3cBRotKoGdwF+jqDPL922lvhK06Yhbq+Ce
+eHPrPYfdm0FciR97yqHz7iO5VbcMSvX0blq2onk55r+JmLdZYhFj1hPqa5hnz4W
/L6HN5hZ21W301tYFgmyMd3m7O/Dfo/GGbMTc5BzBaUB3OkUzHy/R+Go3MqEUHM7
2lDrTc1ZltTLhuQkpaSc4wtKk+sKPnI4IYNxyD3jFCHqSr8slU6rpLu2iNGmlztu
7N4Uz+JgegHumapBtusGHUXLlD06NhM4hlpx4e3ckNg219Z4SEXRfTEJm3/OqV23
8PPPZd+N6z9p8LRpxgDEwKSqOPC1KR001ys3EkqSvmkPRD65aqkEVmaspsy9+2E3
ZtKKCNdBZX0U1glPduaWZ8xh31AS2QYk2ueHgA2eC1XtGsUvrNPN6Ss6JW1hamQW
dhrDN+FE94N+3Yc+0vfUHyvLprH//c9T6C5eZ2HypqvLhPO16ryP2WySJAq5TEMq
gQP+5fnFQnX+AJhfeRz7pyjKUD8aODexT4A/hAkqaoG0NP/upcm2Fahb8CR6yurm
VY2/xLvgvudulH0WM8z8kk2t0BEyKI5eng2uq5YYTuaNGQZ9kfCO5ySgRg2JPAVf
bQozCCqzMny5YcEpgEG39NyZSlpJgAMFNKkPzrpYGu6tzt/jMAG+U3Q8iSKN9QXX
zyCziQP+c+f82wljDlhFh0SdApq5aADVScTrTqyy586CeB0C935g35Kf4ah90Z4a
EJV+/SorHHccJ7FwGLzsIlwCzOsCZaDx258guGaJKLZHl0i0Eg6uBHZZbOmvZwgm
yfltVaYfMIf/WxANY0kkaPfC/jWZlNHZcbnYE5/6MW+/81rhrd7OKojE5pARpZOY
q9pKdJPitBsoY7MJR4bdYf4DMULbhcukHv3Zsv+QZDCa3M6o0ehmCLpKEws+hcey
96D1C/VPcQLLt+fKtF8T4citRYuX+5PNg5qigZ1bGRnxfQvIrQkkwkNxCmC32AVL
lpeWxCKLlhzVv+Qygg9CKODoOl//WHsuzRfnVhlzQLuly170D79SH/dLY6oruRYo
c2P6yLxXocMn3f5OJqFXMqtvBM1n9laSU6kOOEkrr9no7l7wI5IeB9mm/VwyULpZ
jAycBP862tqNnFJCuNL8i820aUepMQ641QB+Z3+KZaKR8dlJ4AXRTSuGIHwWaWoN
NpdUEAVne7a5VmZECDlXsIG3UhQzfpkacK5xQTlGjWLWLRcBjpeKT5VevLIL5O2Y
HxzPJNFACFspKuMclDgsDvifiz2m6VGlG0OtHMGEW65+frm8xZEUJfbntLkNDFzo
eb7Rs3F5JU8iKDdPHqRlHijbvrLX6MwQo2uWLxaLUpRyGXu07oTvHqeGGC84Nv8R
lrGu5neGSXWD2OsIwdHNXYeXXcFX7lpF5QkrubKArOg2MJshKBo0jB+wf5NLHbEI
yadz1u/sb6UzV0xDRMgRP7q58pORWZnGHx9VB2my7xc/3VhioiOBmVColdedIabp
FoGuQv3wxQvYysQ7XEg1cuepNWfl3q37fRfuZxZMj3Wn3KotqBVzec3E0FPE1jWD
XweU4zvQVdR4PYnxAY2eL+ZY1nanpuAo02hOzq8UHjxjfeDuspqfs8OepoRCykiL
BrE8gTpW7hNbIOmbAcuFsSJnEowzkqGRRyj4DgVSyKwKi8N1DzrxeYhN/iE4+obh
nz19ENt4RT6Ld8VBFij1FxwyQ6dAzWyD8FQNY5pVCQCsIhk0e51lzGOfi3mQ4xer
ZEhvc6+B5lsUxqYBd/pWLFxTH1hWsB2f6EP1zfy7yN7UUHoW/KOxOmUQeGDAgo0E
fExEjWrAiHBPMQxOebCFXj12x9bCMzz6Xc+Fjc2JJY04cgWIjTHOCFiIYi1/5KhZ
ahkkhj3/jAHL6YbvUEI6o0McbAcXhKK2/ivaeOZTsGMwEEuT1j4qTaTDA8zbxGiy
SCdF3MaFo5cAJInGQy0cu+Der0wOBsqGrLiv4OXgHyio2TBefjaQqGJ3LlqbFrBH
ASjdl4/ZDIiZJUrDggOqRELIF7QXHaT4SCl2VyNUm7LOnBaA0nUx4rqZJX93+CbJ
vbmMsYaVDO6EByEAewGdCdn9IXEu2aS53tF8M7Jve+ynGlwcBctb09aj63JiEJME
moy2HKZ1HEwII9hR3NpMAlIA+EuxBr1xXEx9vZ1xe5SfoqPMJr6Om0GeIGUcapDi
fhi2M0wsO5RltKGPa5VZAxdPJpuJNf3d8cQVMPYkq+TAuzOYPr1pjpSdzwnvkNjQ
J/KbMbz/JY/PucXo2xl+6AWUCBLiAPQQeeNCe1WGrMf7F/WRoW6VR/rQEMjlliCM
+ItDESfX6o6pCPWtqPg6tNwWelf/tQveBRSdcD/82bjz/3RSr5EJVHg8rSsx1WkE
9dEFeSh2cSbEN/9N5/14ry/h4aU9BWF1394xipy1uxH/Ag9/C+Es1pIAJW2P5bTy
FYPkodx1xrsRQKwChdyIC7CWbE3i+ZiNZwNkMP/HWujeDDz/p/nhEi/BVS4PlD1A
hBJcsfxX7nRlLNNDf4fo9ZL6qr8hanK+D1ZQSQS2gAsS3gso3VCkM5IN4MUTEvCh
jiQU1Zsd5Z38Sjxkgx8fxAAKP2onAGa2Rrzzs2gVJzT5oI8qyoDFcKmjnsXTOo5I
GsC0P0kk0rImms9Qx8+if6iffUf3h6nSE9cL0Y7Z3n/wNqNs5sbL5yBMwR2hAyND
uMK1k5XVyAuRMOFiQFDvFDv7IXHrhbF+H8DaMcYUDEqKWHmFt+GiGE4Vh27iaU+6
0QlWrUsznzKrmZszCJRxcwdtTv0SkWi4dJP0Qu3YvzdJvfrhXCBh4SQQv9LoogI3
p1We6N4mFPv6+0EvhCvN5krTzYMve3LT6iKPQ/+GzEgWzjZWs5zlclJ5oGrfDJQ6
N4amoN6kFaXpEKkfVZOawU/FCxi+4u7rwntdkHPVAs41Uy+BVZYocmLD/MYuzOe0
e7jQyx6fbbQV/fR1E4qRiuKYRO4THYKIORG3T7yFCBZPkJHmIvdaTl5FKUCaUxUJ
SzhzotMgTFnx7Ih2aLpR5RkPDmLAA1JL54XsH7BVnN/7rKNsuTnjFUdV2nVMf1O9
A21IGnFPOwWVcFhFFRInEXUuiQ8Suuq3SOa6/i+mYEKJvgiYDpXiqRz+JjH9JPjF
58dU3xt7dioe4QRhPqMMqBoboKL+Nas09Vak9H1Nfur5XTSG0HH90H+sOgLBzuWY
5cV5HYbxdtJMr6ts+6O64xpD+pCtgZibjWRT1xPLzvnKVCXvZ5DK4v4U5OXzrowt
XlurCooMW5h9LkYuXaR2TTnVEprcPNhOxmh9WMeqiwq7rMYA2l7fI77AYsbYhQ6Y
EH3UmVKpQA8yCnlp3N8BARCt8WCrdpPjqzstjuIrSEXQzieXxULp6iQWyGD9V2FC
zLq+8afVQWv6h6dwIzc49muSt49o3FSxpHTQEY20o4YMEbYZi6mFW4RmugyAazzn
VgOS+dbMlHuv51MWeEDsFYUIdRsZ5yCycPbt0coEt7tpBdW8je0vVmsM5Sza8I4y
pfvmVWxp6vetLoK+KzvN5UNMC+8iKQqQTA//7qeUWxK5IOHiX0VI6M1RPtF9TBQA
ZLouR1HvwISE7DZv9N/gwGlfyzqm2NKafHcHA9iNq3ZavPIhf1Maklszn6re/t1S
mcD35P4Vq4zFOZRooUFZogDEjbVb3bCEgF9wuYiiUNssgEDvAHEB5OxajBlQfun7
RPAjoWqSyZpJ91jZ1ScjfUNkhgGsBwQNWSG13zKElxUob5zI2JWEymcpw76YA39U
uKaO6MsZRk0rSf+VtL0ZeiwtjpvlCBf8HTeO0yfLuY82fA8DgjMEBSDWK7r+wYHt
N8zhGWEy5juGM8ETH5fE3D9KjgRhI78MB4O70nD0tapNrNaWd6nffwUyEE5fowfH
+n8lMVkLIEBXGo0zw4pQQK1926VqBDK6f+5Ns5BDWaiT3B49e1ZqqOWC7Mq74hHT
soaYJrnDDTRsAAsk6RujMWK/NSSH4CxlXXO+kmEqfbQZmO0R4sKeMaKlq9+s/mcG
nAAoXu/+CTJabxRV2kYP8dGrRPmikbwR59Ut9pwNBjcyBW6SP2IeztUnoHccnRQU
36wt3nCiM+30zESXyTBF7D0I5LZoAQ7FQTJXHXywnOgDixu0a8yGvCc5Rq4TJD/+
9mQi6C1HFbYpQujG8qR4hd9OtiUwrbDSRQoVZLlDxzkvxjtNRg1qSM/D5bElZGNf
mTwLTP1v4Qlk82IKPOnXIKGvWyy2OF8/ROEUGFkV1/3tgiuMMxMRSb3QeTC6Spd7
R7DcTvWm7XAXpEQJBkBA7W0kDcJCi/d+eAtnE4ODtuXyA1AstZTj+wcwN0Iantps
s/Q6d1++9CSWEL3KfeWJORnqAIxM+n6ymq3bV2cvf5F+eMsXA7RtjNWVu3l2zYAw
MFkR/xZ6ByI956iy8Mu5XTUJnnd0a13ud5DUXsoT8V2o74ccdTwWvgZafpekweLz
nOfMKPBQpHF0GoOsSRGymOc7nmXF74fCgFoudDOr6HoGKuetCocXNkd+cyPHE//h
2N4P+YZACFdA265wqAOewY+TAHACkZRq0SZYMwiq1Ks625TcKitZDVWz5Pu7cT9M
UCx0KU1f7Bciq8iZuVAW8jY1NUqFtnvxmf4h0C1tHCuHaipx2Q1wx8hlHJA9Ouhr
n4EZaGWMxumjZ6xSItf9IUPdW7cDbZzWAolMpiXOvS66TJzR2+8ok8V09qTP0vhf
zpCQfj0sKkwhfUAf0Mg+sfDEJGwMbAJQHyNpY6NxtEvWZhICnjhUGo7bR1/CgSF5
si9Una6bSgxZabdSe+FZeRZy4ocl+s27q7yXvD+MUL3bSGrqYLpPgCcA5uymG325
EethwVPEdBq4E/VwDiBGEOQ6Q2uj1nmQBMrBO8xfCGbmkkaE6s25KpuY+/KSAhTi
i+NbvMir0XlnHDBAdN515GGcNqcmM0xVZ81jGeAkZKdozYBHnj1C9y/9cwXxtQTy
Z8ZfpNVcj0RUGQAjvkjl8Vv0lvTQ1zyCZh9D65Vwv+0U4wTJi6eAvCimzQcbu9Ks
To/wQZ78SmvaJLpfPI1DgPreXYbX72zC9iial1DGxbCdUb4iTOtue9xao7Z+EfYC
dgNMWwOvJMLbWN+5HO/2o6q0j0bmX4fNgSWigL7kOE43TK7LZWREOOx4Zdrjfu4l
5eRCMKJoK53+VNJSnlYWhRtG7xA3i6YQ1rj74+RS2J9z72o7UeX01Z9T5ndUsoBX
CgOZ1hCvKeySFkpPT7Jv7jr8T/O1SXoHNsMmYOg55MC9DfrdTnbF47xjuqNhLs99
kt7CrbG5PbC1NiTHTeHKhX1ips9ehm/8xhXjHDPxFo9fVO3FoMNtc5FMCgU574hQ
ri96hkIwsGUZvztKOQRGl7vjWlBC+E2VnksaUIx+cVuCVqhjYVD9h1zi0MjkbbmH
Zcda774qOMCeE/HAXuEnyRkbtjJmZWnkxsQvQTVSMV+miVwGxOXv/btNr5bZKC5w
fOoSqdnBCFPws81fwviPJMpXgTU/cxxroD7sfa40ewoeCuAQL6joV0yRMQKuCgjv
72zMyWnM2RgRADQjz0dUKxIXSEgB3F5V0qtJ0VKiyylJM/RB9LTZC0j0c26CCX7X
vBBn/vHp+oPonQ5vyOYpEQqsMCPImBILjjJoAr/93qmnsdsXnuhDSO5JeWg39Zwh
4BHzFkKq8TnLCd6eyvZzak0r1POofIXJzTmKBQLrf+zzd+Jt2wefx8DKaw+gZSpg
K6ceZCDfplTLDsKEttbEbHCQD4je+gwXRVh2UDCpe4btYvWR25LKb/VXGY+v49O/
/gAxPp9+OOkjNAw657O0WNTUGYCrFvpeGFAMZfD7GBREr/e/eXqwaNEyInWwfNjv
OWrF46gXO8fDVQ5fpvY7yVXt/c2ORL2NAhgFRBrxbdwNqtWY2nDemQ6oR0FjVJCF
hwcBMLCskZGSwHyr9x+xj0h1irodUaZR5FIXOyjFdszOCxoi4KaPovd4H+eP/lEL
dBQwRZAmG50a67U5NdQvsRySpExWNunUJu64U1IJ+RuGK7qkPtpG3hTPLEap9PJa
GXuwHYQj8/dHgt+4Dpg/JH59kDXQ6gElZMycb8QoRcuIUH1de30cIYNTGdkWL7Zy
+lgMZbXhW1dVzUVRgqiHQ48+fFZXVScbLB9e9mqFOwbYEw7QiWXTxxakjA7eXHs3
ctKGgxSuFFhwsFQWIUHzlgmYewfd5ykAlquP0XxV4gc11xmLhbmySNarFE5wn+8x
xlOVDngdDcEb/TUKAxTmoxZDIT+J97nTCkoPzQZ8mJrangZCwH43z9/Z+yy+yn7G
nMqUTKGduIUUaHceoQjQp0fPYVNFDlMZxppjJzbN8xkdgIG0D7kkNmZdZZgltUdW
dQzeSdeXLZ4lR69VhyfJTMViFX8rT1xMyxRAHBbgwmwq26FLVZonJr34InNuXXQ+
d4lJLoJaub5ad42rNohXUE4/q8HyxaiNTQGcqtLd8lhPg4J9XpiMSHhtUxn/CaBF
UcHklNokWfECfAraKBxlbdBV1vcTTYBWJW6WM1jUfoFyLxT0yXNGQix8U4lUbsbk
Tvy/wXAPe9qzjHfdBpfFFU56IPlOFTNvVDPKM+IUlwUaMEK5gK3MbeOcn0trrxjU
hiZFOmYL/4ccnbIUBOVn1CwlVyeTsi8hd/Z1H8rtSYbRMnY8BUoSazaq4itBi5hK
lo1ksz0iTaKBLoz90enAKmbIrsrQmsuPmdJqo7uAXf6xLZWGuL1qAKLFq1Vo5OZD
XuwDBkjmhOEJVI2azphvWBWx1a3EDv90HL6JLrGBDj3P9FcBG4SXnJjYYu5sY3un
ysf1zJNexK/V69Yd9mTmDamk1X/tDNBe1xybZiqTg32aayZ5Y3Fs37y0At3X8XqG
PxYBX1Nn6yGgSjAPHvw3N7FlYNfnscTN314WlHLR9OYgGLxIQm/fChU5vmbma9tx
yWm5e0/VHSjYOU46Ks/3BPnOig8nX44LTC7BNDnUmHnRbuPPeEcs4cVPMScHyxLq
blZpljQ9/uEsjp7KEvBehD7vYSh1e2fTNne+YOwSM+4ovLlXt9IW8OWlpfuRuE9K
I5IJ1MHImsTmPTok27ve6Eo/k9BtGR8VltKFpCM4NDX/JfQ12PU/wNnDvIG8HgS/
8I1VM9hiWvGiyfmD+LsJI0P/2XUbvmF8gzSGAAz5VFCboRbCF93LOYRI2Jbgw2A5
4Z/4BPIlsEud8cZFPVVogC38N+9dogElPsufcs02QZLMUpPazEyPrBFvu7vQnOf+
2x77VsXzYnrJ/zL+nIycyfOhRjiNj7jf+zarbkD6yY3wWt+3asMzWsdfYEJ+nX/t
jwd/BLCg6s83OYBVJHsUySKbsr9qkqw1FEVteYpIZE+yRZyG3dFfCDaaQa1uW9iH
P3NpS5oB5pio5EefYnWCfJhGARA0PDilOkJfxpKmYnuRV8NClP0CPaQM6CySvXUW
pQ4O65gXt3Iq6OB3m2sNvz1yZD59+Y7itEM4E9gWNlJLa0wm1OBhmOCgpXDeygC5
cdCVVKf4xZPSQ06vE2tBG5DQYXQzIOxN+CxdkUBOr4Cw1KQvbbVw01HMZ9h5Sxnz
4W6Qi1Vdr0OgTphNzxvCwJblW1r966idjPsuEAg3b5sh8I+b6qWY32hQPbFUrvou
xojKi+O//ijR67O081KQ52uEgGzYniZ2982dXruPtme+425k/dD09SH9OjTERKW7
0U8wdN0IGNqVPod8BYhAnZ6hl/UkZKrKgbggRvrCssLa8bFEW0YOesaA06gIxBgO
Att0qzCu2r96pys/dijd9yH2MgTXk43wNM0FfHakP62o+B8eiDjlow7KexgD8UUh
TJxTPfzNVPcjcIC2YkvfsgBVISbbHNOEMu+taHmVLrR81uFwrSs7KgV1RrOEieEy
12krSqrHKthqTgFb71edRGGqVWbQ4Ojctf8ZePFcxoXWvSuyCWZ/4hbQkACPxUKW
c+Bl82p5DOifs/AhQkMHUavN6bntFKkCTvMc9D1rLvknAAhAU5MGlmFTCQDq2R04
wyDSyWhKxtsnce+FR4OcfjcEsdTvahWDKN2gGE+Vb5EQKa2glhVBc5pz3m1+4GwN
zzA5wViuhz/Q4SWXA/CJBDlfHirxbKw6AlZU09Z08VRNs+G/7RntH3FoK9I0DHqb
mLe+83mrZb/cABUxduN+I8zI+rjAf91wji+7n5LqP5F/XUGepc1AYVNmwivIQHz8
Ry/tA7rzq72Oab67tKn/go+3HhQMHt7QAkSLbmiNjJ4DOTB4OvtS73MLvZHY2qYA
LUqi0xuyXLhTpNE5vJTgyehNPWLL/USa98phBBOwdu/RVXlrWVEAGcY6PanxI43u
TBsvI2sXO2ndLUl3eV70V1QxbXp9hplFFEp51wGXw5z9LqQuJxVCbJNLon4IOx2D
rI0ZWn36Nrod/4cqiCaULTWYiusYYQ3B0n47xH6/h0QBKcwFvE9SBKQQ44jgIIzZ
uPtFLgLGpM5vj133CthxEu0RjTr1TGHGTistCLkuzlCBOoB9XYXQ8ybd3XKARbYH
nVtS24stI2PQP9ch5ruP9s4YckGfqJkfb2prFxfg8V/YcmEI2vHqTD8A3Ye1oydA
dMBJIo2+OXKTRbf7IJZR/FHL+qP5aF+DgSzFYUF8cOHkAV8o7LDkFR6vIhsBYzwD
Hjo6s2rMNepFkL+EilSp+4vh7FXcsfOpTEytxTIwlGcLg31GTGPXO8yWewi6lZbX
U+m0PAR5MaOsO8dsb2cvhkU4hROisF9FRJ09OAO44c6oyh0nX+dknb/FK4zONYqp
kllrFb9lVRgMIb6rGYwELkABXKBJyiyu2QRORKyJYBX82hGaQx8EeyF2h1ocee/A
6gtSCprDQKM15hRRU0o9jAxrFtlCQMP+J799j2txnSTpIQFanTrKOfYNvsNLVNO+
1VKmwswqeNcaDIozqOic5IIzCosi0t3UTpe51jx566QocGC3E0i3cgM20g1nnMog
rwSsLZoD6Ck7zt71hY7OKcP7/U2AzlD78/4quiZLSCrfdUuPdVqg8a2D04XpiNOI
o4sEEWoqi9F2oLXGm9HHZBLxqSlXkkxKceR8eb2kQn2+4nC6ZehEtjRuYsSMlFgg
H6sPuD7EAX2nEK5wEU2sESKDFK8I+oMDI+q7iEPr9WZdelaz2RGtQsLnEDyiuDx8
oRtuJm9uaIg9T1NQRqarI+pEqjhz+ksnMYc//6XSU4NZ2iz9y94/Iy+b3TjztK+G
+OLalFDuxqWOLCpYWQODYrWMFwf2R+PqqUBHhCbdMuimAMTM35pnU4w77q9t6Q0K
a9ydyh7c4El5M34+set3KSBEm++s5ybWSW8o7Hur4xH26RZWQi/zVSKZ+BSt0X5/
/uOBdPMLc/vf+/Cmx63z5hIBcrpKloFKxrwKppvBpYHuZM/OmbLGFNMheFjHYrxM
sRgwLg7U1lAv4MslpHXUXnkKcjZMqDdIK/5kgrV31mZd7AEM/22360To6VmiPAqb
jt/+XpUJwz/K6h8dAxBh+dndrtBiXsA7gzLRvHati+uniIVKUDaGm0aiYhjisZ09
cgdex6lL5uY/aUnQ7/mxlmS+cujNI7cgjqtNbVnH0MBtTKfTr3cHjkKvTyvMwhHn
lsQb9vlc//qCY98dug3J9MWxC7f3PXAatENP4h/K6FlSmkDfMbJfpFLZVnAKHXcG
GKPocK8YNZaqV1bZmA2kJhPSAwaxJp9TxDiSg4IbxXF9ZCUyj9ihqFMpxls0ckMJ
EblL3NkTa/aFInl7VUqqY18rgDFzvFXiUdX1If2BSL/hsltjsl0iU+Kc1MpgDG86
YmBuunzdhQOmMg2vNWsSCuKs79hYPg27B5KbUoFg2+sfgfXMhKWb7d0H4TUUqGiX
vz1d9o2hUq2+psGCGkxuw1++rzWiLlGA8rxbFEK5kn1R5BRcSgFJrvV2nFHSGjft
5LuE9PfhxXfRrfbLXkMk9C+TwXiZWwVi2PPNy2Yu5DiAn7TqBU726saYfKjZTS2j
UqTlCThab+5X4sjABabGDODeqAXOPFnN6BrEb59djWuhIHu6UW4yTl6tHyKnZN/+
8dZJe3H8FfVtQulzdm+q4bDdhwL27vWmAtrv1sIeUzYFeBnX4EwNhoiucJD4I3AG
a1ez2xUf+9ChEI/G12HShPSNLEz7afRZq8xi7nyUmIhJlKpWLtQR9TzMXF9xmA6i
tnbtDyVrvJQho0A8tyM3WsdsYXnwWCBD75j9dOpB0HWTyLiE5xSKu+2kNEzQ4xCW
hLrk8B6XXKBoxMNyS6osslkCnheXtGoeuG/Xdtc5LyM2IeSEPAiCxfJyvKAqAArd
z9b8wvXZ7WE1aC3eY2OCoqjccoHVS94/q+XCI7asF/jv3/mwsTdV4effCS1UM/Ku
jEhuPvlb9pf86/Dia6HNkXSH1t9Ka79h+7+pmA6aJcwNr8XXp7NIL7maS43o5mLu
Bf/Ou1ztCFaoUWO9iYag2LOVqUB5RouQFcFm4rJw6Du27nMp1TOey9eWnScCCmHt
awwfaTyVxzekolYaHHFMgG/NIVkRuAGQJ2Off4H3FNrng72TVI/NvcQtj7et4cqI
/VnW70Txrva5liRuotbq4CIongEsnQB76rd8Iz3PvwfFdy8DmznOJKd62hC08hl4
Um+SESLge44APMXt7S+H8bbx61+cpiK0aQaVDvtNSt/ME3yEOlp2R+djG4FjddVt
vVKi9cD2goi3ctl4uXfhgCW0YQJUbtOMjczE+XXi5GSCWb9EW6Vjn/wfFoMQGNxA
f41lis8cB9GCkl9ZIlp2vcssHRnd/MaPv9Au8mg3KOZDlY/OPeDyTo0x3XO2OZg8
vXd+P7YQy8+u0Rjs36YJNRy4G6S+x+Axlykjllc+EXGv1tLQeBAeMQ5tQHCyqbCS
5n5ABTiy5905nWxMR2VXD3QLUAUJ4KQUWJRRF8mF6qxd75qc9gnsSBGTYUs4eMV7
xSblp8XPMKtH3izr5U5GK8hNgwlW4bGIHXjODHfdxpZ0geVUkY0WaC9XD/I4oJOL
pQrXpZ2Ea5UllqQbP5pQzbrI0WQAeXKhqfLMWUzZjb8aKiWeTs8y2pyExYBX/8cc
IOrNJan4Cba2FdSvZiTWtVaKtmCbVj+cDtYTwBAaJ3sIxQb3yh93gBeauc88K/rn
HP3HQNQzyx6jmrRqi+mpmt51a4fjj68wXzgN8SRbOPSMmgCm+62QoJNvyCE1hWM/
6fKuKYnE9Fvq+zviahoQUPQDfGBaGYAtNu2KZaaIa0Ypb0ssHpCjkGFIot1+STYt
tp0uOXvyK9FkKV6W1hqeLSqWp2VC2EBmnDw8yQQoL1I0BZgn+5snSeB2/MRezIPi
jG9MAwp1DAGp4ys59EHVJ0uwgmrNt9Lnk6CSKAI981L+cRwuSyjcWExtdZokUVHl
Hgm/oz+8637K62LNh2AxBiTRWMVt5btfvf45LEs/SM/wXEEl0gkMlaRwm4l7goKD
IaPtdOQgxTbJMPiGjCJMUGVTZJ+5MmeKOHYQI91nxKkBC5tgXS/1x+AgmWkIH0v1
dvFnjyhdMGAjlPIlBwfFcF4A6MYIqZP0vNNB8plnUCZc+fKDzo2KTVeFMILI6i39
Xpp9zQmPwzzk4fvl9Khtk0KnNvfcPGmbeP26+ady1pcwfCkOzilXl1a+wX6WUTGN
/GwgfNv9zroDPqSA84OBbn4XpbAEvUJ3kmRjsQSykn/WxNSFzAHo6iU6ulAaX9V4
bBn6g1TDoKv3mddC9tYiJI+rhM2pYbvtnj28VPA0PwsSyW3ilmI3Vnei4cScqXVe
1m5sNDBqWJIcQFR9BJTAXf4+nMRtKWa/3aVYwqzR2bUiZE+dk6gGJXYL+Z4+fPit
LSfBycguqnERZ5AcbVB/QZKF+9za3zhWcFKpg8FrPRiUuVzdqfrQKTlJVD34/SmJ
3czd1BcFHONlNVmTVF4kjO2VLWgbY5L+9kN0RKY7pZGWeq+piUweeBjM1f1scEa0
9Fz/kCk9OHxTEiW+pJdB9xekpdjq9FMhDuZ1FiaRUojDmdXvfxcKKVuJU1IKRY4d
Nm0m0e9DZhiPzD3+vp7zRLyPDp/Rt/+cIF0VI8d5JZNKrNa0meyWWjr9RijtGl5x
fcQgc7fhEtaM644M1grAat/STlVB39hctOy1kFEkhYMUhZYXAGYx+tAF5u5RXosz
alaIio+4Q4Y2HD7bXkeGhPK7KyAkO2XkYal9W9owq5wC/7LbksNTilBUSoWHUxgz
e7sR4Dp0jvp311dG5kmuADeI8GrJMbjzA3sy9NtFqiHklGtxMLd+VJGs0uL/25mJ
KBIV0ecqxoaQ5KeMIj64Lkc60mzHFq8AxyNnpzp5k5eswJpOyGr+VGznd2u0QKY/
msHfliLvodhfiG0henV6zB6F9GAY+dhKBaMvb0K74CT2a+VxqjI0g7gi+eH3+Khz
eqmCWcaooL+twWGOgsPj5+ioRQnD5BFAQeuO+pnPCTp6b9Jrk4uOZEdR/L1JOHL0
A0gML4tLJgJs5/8dRQpuwZp0hlQMbdxHNniXy343Ot25FPvDtp7/whCExWRMnjLy
4gVIFDtTUYyCBcpb+DRA326NqGF1aGSB83ZSOFnB3aXmIiX8t92tXb+SJHUzeGPR
7G8RbnMslcSzjzBo2y2gfgH8pR0miUCYTN70bncidgN7jSyAs/3RazQnV0kOFe4X
3mg6AwuVT6ZmHF5lTxJcCx0zo4V4siMaX9z8lpgWq3R+nkWWrbnnvoAUorqmPuBf
/KQG2hSZD4lia7096wv0SuXthMr5OZpz6c9dfZV12gP5nzIQb+LgDwQHf6mBEcH0
5R/CSA0bjSjo9k+y9ssFXJtLu1H84Rw1gEUD7ySiA6PljlrmceArLmn6AbybPtM2
BjRu5PYkJAZDIAZz7lRcaTFR9XzJ2au3G7AamlygTknc5Q+9M3L/VYVb+/RvWIp8
ghAow1l3j2BCBPIA395VOB6ePd2aehA4KcHYi9Xx02m8Xvw/HNdUo/ujtmyR/WZ9
oy6vAhmcCJCs68jczS27ApZQ5ayvXiDIRlOGHJ030NDpRTuKcVZMFWmhWRCT1SVu
//zsT7sFpYK8sR5f/OWKCHzJoheZ4Fv3nqlXRUd25jsWN2jKzvVEnDrijaBmnPX9
9xYhDq9rN2b+mgCXgcJ/yOHdsPeXMifxuVxqVHUJvzaI6UbkWBMyapvKSH7h7sUg
Twy1fOKR6qfXyDIXHrUorTQXIcux6bmrqqZwg2NKRYZlOhTe0Ie0/Fy4eocEyYeX
iVBI5dBpQRpkdPjJWwzD7H/n8oFNJJIdF2I+5rgyry+85GvsdWLUKxpSN9DgcK20
TaGy4CfJEOdYmllso3Vz7vo/CRHauAirhlAxwgJgdcP/AqD8VwZP+ljW8Z+CBVpU
6nbJ/zp7Dycrmgj/y5OxONn8fGPpCyWETVbSjR5aPBg+yvRCm40TSHOyqoPaFnmj
O1kCdu39m6332GsUGppHabgENP+b6wXMaTo3G80WDHt5j1//ws4uGfMnVSzEuKJU
mbb+/h0KpbU6rT11TKxtwzecQrE2qobcox2uoh0R1Qcew10Sn+8B9KN6JuIft3cS
y8lFwfZNmlxAee6UsfNLL5U8T3wIQ+dEB54nlKFzOAwKVm77r0vOP2+C8c5l9Mnd
/p7xr05FlQzO75sUKCz/Fg3J4NlLj6YnbaLqUYEEaFUSSSR9Axg/yWHiseHAa6Yn
bp6A4wCR672RjqZkhdhOesZ+a5zcVkv9k9kHsrJjWGJVd+XxcJNdZT/jwiwI6TsV
tcSaRTCBixk73/wZ5x+x7KX3Wd7CXVJ1ULiZW3gKCROt5yfSCl2hZJs6MC5isgME
/9/i9rUkWDz1MFuMwHfPShaTy6jSJ6RJxaZZCIA1V2IUq2bcd5csBmmUNOmoXb0j
mXyYofRTmAA2XRYzywU37Fa0/6JlUmL318cMTJyij1y5BzoTWnXh6eghjaQmESv6
LgANAgTrfl1cb4vN00DDvJy+89EzTpgTJORSnDRgtNxB0TkcIcrEUKz8RlfnCyNs
l2eeXFYHJcis9CCObtkD0PKCEI/j4ZcaoUxWF12erPE1PvLFvZk5I87pW+HV0+nO
PhJNJrycvEs5MekO6iYM+JMvbGejeSWtCleei5UYrWGCIgp4FYyt62RmeJBKSHGl
nl3O+8Zijc0lzzNNYYzNz6Sr+yMI1vr19Hv7hgDdhLxNFUvq0KMXuo271QMpeklu
jYKsm/fxysEh4ZptNXxN+RuiqAW8sSpjVTBznjwSV0vxujOrVUJqwIPesCGjZYnA
a5ykYb6KZt0perk1dDkNBLWHURghv1CtSiEvTGs4mDBxfJrP2/WMFdHtvARbA5N+
+BjDHwsVboWdteQ4UST7+7tkZzEbRdQbd9YETGHzMo7pBXefrCA1GIpc1vPlD8Ev
MtahzoQErTA4ljE17dKcIeZrewGhErKyKQO2qWqL4Hi+SYRT37TNP/HeNArwisOa
IS5LH+2J1QWhkeo9JMZP6QH5RAO53+DfBX1gPCY0U1g9PsydbJAhPGzkYRpAr5Gv
rRX8iyFc1AYI/xUE+wE7rkakGbrL4CDpOLujRh7lmIe/rHSfWyMpLwHqb+5yyKZn
MnyAKMkbTD4sIzY8FVm+sW4NsCk6TdDKkgSVlu4XGxvOqQAgg6FU2UcUzuSd20eu
0OuUq5SyHXCieJE/WV5Nfiqh1pBpz5Hy5Nwxl/6t7+A+ANVJNk/PiyUXS3ld/t+N
+Zmw39ytq1S/PPOa1rxq1sEk7DhB41lC+SreuIeBRiYFgCa3QI37T1ipxkVcd91f
fraCmy3IUbfIDJIGmH1QpJT5syHYyyOnD1riSIp1wYQPdrHuhE92pT+mQnqBd9Qt
vo2K93K2FEX4Qs6FRyIIqvuqcKVpR079iPhiI5mTqlz2pVYr9X77jS6+9KNEpi6b
qXcTJTkTV0y9gv3zOqq0x7miAQnYAuJjkGRjoQidIsJdSzdNep7bqeNqhfk6tT3t
KZPVjQO9jfEYua/Z86T8cMiJCp4qteSf8VIGTe784H0j2kI4dqDiYn2+2KycJvDU
ZmIgY+6PpJfgMDqLvVlxWRoLU1AbQ2wLzoJeGxAh/k0nPxfmXXpstwYfOBlmx/YH
OLYDG1LLo/pc2P8kZcfIPHEeTJD1SxeO0/Ij01grsq4ETlWK5SDOGVaSLsGpSI76
azYzzclRWrhV6+SK95ouP81VGz9d8FwrOjGpOhQL/1NVY39S1W+oiSI8YiuKjuQj
Udtg5FICKT20m3sh/BuKp/oXjKqvXZOvEbHVQoOx+Edi+vgtjHcVE0svY2deGOT+
KUTUwRMaOfIh2FyvJyz5e2DBpV9OHz4SgR0wpBrUfcU/f6vu42gdPCeqbqWply0Q
t1Dg86iQgKDXlaeIBO5zS//6haOuEYWWMQnL0Gq0RBUgNJuBgP7hLn5p0w9KRfn8
gat7D4S0STZwUhaBTnrTIyro0OpKF5GtMBX2Ym1Nbej4FDuuB8No0oxk8orXQXhT
74jDIx/DulKBzpnbDO61y+wMEYhoXambgZOLrtORT6dCLCI9TmIjgqk4YrDp/Iw+
LrYkC8LHXEvNjCc6drGR6TPiiSQ7sr7iv6v4HzGHaKetO6IWfFBqwMifQ0OU6gox
enyX26JOMqRY6R87+wLKmVP44fkTDKYkrWxqcSTCwHOvbhsqnOgnOjjkOTdK2fSU
NMtC9cB5bRUQDPRGhDref5Zc5u5qqd5UU5gT2n6gFPsSpfrRJ1dmqYR66v65zl7C
qUFKEpm9P0kzZkaLE0EKhr9IQAB4LGkWat9HzDrKRQhjNiAXzptrjupEywvu6dbA
ba4xWvUNBTcg3hJgkozE4bu/clzAtxh4//PIRl5YbQJtjsVs27gAfBGNDWcvsqEa
zHQKLzqa9oFmN2yY1mTMpP1rqSAJWWdDVj0Rvwfbo63ZP/+ybFvf6Xe7SYgi30Cz
/T1yKFf469QD7ey5DJ3AjIfrDQQtTCHRSHPNTnXmrXK7XThqoLB7CXL2034xunDB
ECzIBY6gJxdh6wb9FdUCRyDpfKbumCNUy2TNWSeywOvoHP37+xkpQCPThHyjx1g/
xE6DK1UeZ1fVPW7mbHd8SBRY/EBDvq8/S1GXkWyxDz8o5Qc9v34SH/GL0ydLN+w+
0z5ESIyhaAob2nJQzidAv2ezuf4mgYOv+QlaYDUggMg4KAXXrBdV9+YahAw2jYmU
s5BcUjifxHhXvquFuRpQLdlueo2eNqXuXBMcTg6IvtQPh4TmFBO7jo71Z9yP/FCj
S9NgwTJA5Xn3vC10vPd4pGCxQ57auQ+TV0ZQm0QeKxSzmlaNB3H16UlW8XqwhnLK
aDcRlqbkrPwx0CK2FdlSIXCxh1FkM+91Jj9BoAcMZyHe8VTAt23WTggOlnhd17MU
R16wytoKgE1xYusnPLTyLIm8XrhqScEp6L3U7Lg4pMvE63qSYHb0jgtRoq0/+RUW
siFqtH3I2Phe5V1FZR99yCMZv5pX1ijuVA+7SoqsrmCQjcUYq2eM43w77YoG7Ewm
gUzoGMX+XhUovaPm9iH2NKXmqGIz5gHE/y1OVet7Ara3mTtrwh9jmH3DHmV/K3lG
2F6nIPMliqNRsdAuORfj6ivtjJJpsPySmU5Xbbl7OY1GjQ6orI/4RtCoUJ3sgoa6
+otu8IJQfilecsGf/kN+7Mki1eI3c6hC4iyTM7L6Nv+juh42QaRtVNS6tS7tzM3B
Y/iwvj4GJbtO4fCHGy5Orrj3syr5qr3sDDapT7R687BmBBK6OaxKswUxjOTC+c9d
4BpgJwVISX5W48zJMol3f6c5FT+aVcI83WcNobu/Fck38wdOAgSGXyYq//yk+0ak
NzKd4w50EYIxDr9sWqwJ9IkYSBp6gccdCGWfcBJLxQvHqH+RUvnpKg9jOG6+LJ56
m53e1yOTbjlxq2efF3IRkn5fbx7XXOJ+MQzL4osyjxy3+PV0UoBl17HnxN+vrQat
O3FVSEccGib+1nod+dve/wBhw8Y1W92HCJDX8PNv0yutI0llxYG5jw61UcOVtsiz
NvkVX9jd/dDUFX0+wqEmYspTGCRykiWFN7y4NKxJZ/hHeSluWjynhnXrF3iK0Plp
cKV/Y81FS+FtLXpJR1dZCA0ZwOq2q+Sm9DabAT46gl+QgMkHp1sd8sew1w2p/TJU
9kq0jsw4bqrVJK36F0hhez50jte1STbUmfViotDc8hRcwv9DpSpw9aJ3/ItRIb2A
QWDJRlUC6MjwG41BeWiV6MEzR6DndhL8HPckXcQq7bwQwhbqIGgl2EHfbEmzo3jO
eN0CEs54fY0jalMPT67Rc9ishxEuH0o/y6mOM52naXNcx7EjpWpSN+KD4VirxYhu
GA0BitY+EBDa7Jl0inkKHwr7kJ00mvpNvX/RgRMTXB5o6a+1f7NWK4epqOntkuoG
tCw/6slRM8Nx5Py8GbB/SeCameLHOjRH6/OnJTjzV8hNXxSOImlh39XlwktvOcJc
1OXe05SvqJKX20QG7262yKC3t6PzAKeLGCttcmhWlFW55KXQqMeRDQtID/tp2Zty
HYQWL6qtK2emSXCTZi++3XxY4QfenbzLRORhkDMbEDBslie+pIkvqCUhVuo8SKsD
gIy+trW6Ueq5qKXScAa8wCkD5/zDseF2TXFL6myuR7aOd8UquhkrDsNZhdvTC1Nu
aQsJjVF0tLfxUb3t70SjH8rX8/530k1zwt7+vUXp8Uw98iNrZJ5eVe+L324HvvFP
CWhLRSXD9xrRCDItQIbXTm3GKwMObKYDWSrxd4MbnWHaeoGN3y2b4v+O7V5Fp1+P
pErnk3/z1vlmBCYRR7DcxNRiRQVT5zt8guzIOUpO+rL4ruWAMcySfVyb4BW4kUxb
Jc2ByDHL7bfcmvecCR8n8zItjJqwSYYhbkJ4pA0CHKhp+VUZoGNlfef1jQgPbdrH
GDVDbk/nL9jY/HEs/oUcaotW7zGUz9C5uPVvBaQwpFKyD9JJJ6kQAIybUGqpl87R
7HDW2IiJ1h0UqyscUnqO3EamKDqQHYUXwKxSnOD3b+bK7scYWoW8fqBVEDC8S/Bi
IY6wWR/EHAjopyX7buiNcZ2uomxeG1wKpT+sT5wByJe7A9NhMDuSA0VIEt2jP7Y3
c4f61i+aXFL7Pk2ks63OcmQ5CmwiFz42dHfbdUqphWlq0KzOk11IxmhBfrE7Mbec
wUHKh4AVDKYACfmTTsD+SKbcj2ouR04XpROcPXi12Kd21sK4uXS5GoJtr0PFuMZU
/T6JkNSouV6wzAEvoqJE6VyQlN8uZZQxrvIYuvup2r4o7Oj3hsMbsnDL2DoQ6j7n
Eyn8qMAqFHQHKmv9n9RuuLu1ZbiRZDcCd9bFrqFu/B65jhh8HN5wU8w6hE2gB5yi
Uy1ZFtbvJNuIBiu+FsmxYxQ+VPHolUWMgLCSX9MpUYyPgL0WcsslY0tvqb7sMAhT
hwHVu9kHCuD9d4WmjcxCVwrXHGAlS8mW47PLQcKceZRFf2PCtA7fCmgezGoei53/
dp6xu2qXA/eXeYbcLbcNPLRDvQuC4Jqv3PU8zESasBal3coyQl6qn4nKCbDjyjq3
8I/xP1jCwu94fo+RzXu/8rLDFLTza0H9BkWLGu+IQ/2hvsABBadOiwbYGbrPt6L5
U9kt5aR3vSTzCnuDsQG9E5EQbMzpOwB7n+x/6vayh2gwVnI+qnT8MN4wher2PBPx
3r8rDhvmooDhI9GLCCePQRBRDDlK6IbNBpGXPorZ4gA+7mwlSYnmgvKMV5zEdxWP
GsF4W4TtM1IyurA2yavPnG9pkDvaeAvZjLH6ZTm7Hvxh79ZPrbrepfa8NwCjfq0T
W6H4UmHxPr+AVSW9hROJHTeC81wPUG553+pvuxwOfuXr0mae9NpYFWea/tyJOP4Z
QbDStINOd6H+gEB43xPISR8sOp6McT6y5WOnS9EfW1ifikfio8laaMyD/tBUoyz9
UTWf/igcauozcLuGbj5XIM0B+bL1Qnk0YZPYICnOT1T7dD9WM8oB0f5Ln89D6nDC
GzFmDtaj951HgKeCQ7VBs4lMAmKUuLH4qpsQ8H/r/Mt4h9CCQ9FeiIGOMFnCv9Os
IvN1dqHlRvNPxlDhtl1GPC8cJjiUalNPjLl55VkokDwgv23bozYmrZSHUIkQkNeH
G8r9geIZXNN9PfFKxP4CIw0BXg+WcznnyfK2Z+T4kj6OcWEV4MC78oInps0z4duZ
aGU4CtbknQpbr2t+BxwsMsHT070rF66dfA+TKRX25S2pqObf/uKNR3Imtm+Wd/2G
/COxASlWTug6yYWKa7rlkPsYBSwwq7eNlqV8qmIz2RfjTl8b2iwlpmWefSSThqVo
VN1YZEdWKxZmp7Z9+th3S99YwEjj2D2bul/v0BL1xSKztBHuVxmiJFfPs99LsuHr
G8XMN1aIJHIhmRgAJGP2gtudU+YiN7dfGPw/0uuwGIVcU6b4Y5b2eTmgnG7TkllV
hkFGhmNGwmE6pdHAb148g++72mZ4g8Us8eykLbusIZIFK/co2g5gh6MuqMAlWEQm
xMgJIz1l4ntTCT2da2C6oNMczOvZxkRmm+1+l+nFgSVRyX2kq0aQQqqWAsLvbjeI
Ss/YIpqWluXFNYkSSHT2PrbXk/ROcrUtJOuXGakTRFYrEiHoFSuT/6/mH3jYekED
PSgIZ40Jvv8xY3OrWmb3SmoRO7oes4iSLBz4xmIR6DH5HP9jIabh7KymjvYMLAhs
rikYQOcUfj4dy4Ju1lJIpZvr7COLW6JdtynbY691lm2oWxHx3IJCgDV7hymKNG+K
0E8XnrKtqYx3I5xgZyCZkXkdyIwuZWSqJ86u3Hk4rL71AjXA3RBdX/B1H5Qr6bid
nWHFwikZMGVbQHynfuiCcfQ/Suj2HvO4PEteE7uc1LE+5ftkY3KcJCelpVQbWQNL
Fb6oO0ul8RAsnY2hUkek2xtriKOM1604dLdhzEviaNGnLSB894ifGlI31NmzOyPe
IsyKPBCcwYB5qJeMfaqhJrOnkG3QtyPJL9Hsy2Ds++ArEWTeLXVP2KfJ6Evc3qhu
Xorzi1fuqCphgW2Hez3D1ZR7rTVLjAdpKY+Z6R7xkUVcXa1SG6vGw8BMH/V16ty1
qaTVB3H49cIajkE6dqBhHKwgZ33IazVxn1QMFNuV96q0hrgG0sAxXrLqIm2epFOx
QGKhs8XebQCet6mPJQCd5OyseJqcx51jwD+AgEDtjPN0gKbNsZ3F3XXOBiwZMXR/
nEL0VUk2gQ5cRPxXDQsQXs2hJcoqZ6en+Y5Qr2A/rVgWaab9hZIjeOgByPVBB+qf
FaCubK9poPJSDTMPwSaagFp7t3QjokQPZqTEKjqqIq3PClISA7SdqJ+74XoZO6sA
fjZtrK+Sa8LaxZWNhcT6b2kmXKazPQenF39aLLm0fwU2yHGvV1v8JDqLCaKoAYQC
+hSXE5TXLf4hkdLcAaZVhBaH0UmIp0ztHmlbbcvXe7nzYEg74HIv43ZqCDANDpFB
VdG9wL4wis6EVLGh5kuSNfLJVyYy/2HzHw7zmA31CD8KPL1qwI2CCAAOSHEFarEL
3tQHzSaUjrhSvbay9PxveS4WDRstKSabjB/6ugmTOlICi/jvjsY00pun+qznaYLJ
X/FJKMwjLPSJ59oeVhufxF9w7heoka2e2YusRT9nvpykYWg54wDqlcdmW2WFVntJ
giLPj5kyB7RzgWT8fxlzS91dAqwhy75z4GyP1/LaoyAB4taJC6RQA3pAWmzf2P87
ZYj4DbcS/jVD8VInbWFgbuEAyQkZ8Wsmjse+5E3//lL8s5kGV6aPTU0q0w5xw91G
3ufORHrfjAqv0KfFfK5zDgCi8pVrd0nBuUaBeWf9DpYA/FF0QQ8ud93ZN3wEjOQp
LxreNqjHb+oE+5PYjAAEwDj2dvex3G7zuC30+m0fm81rQJlIkapvzIeOShcdaWKw
UhtLCou5PisvHAForfiGB565OTuOElCTxUwzCqO7/aOyOaCQY2px0kDRQ9XvwawG
Zs3rKSKRTZulGDQ7ununJOonLX4fgBwpVU2EqkN+9H4luiNz0qd5JoXb/oAdiCKm
etT3xe1trFtjU/RS1M2b2CYBiQjriTi6iXOcm+8fqUuHZimjneP17HtolL0NTWw/
Ojb0zz6PPjx+naPlAoaPS8BFIQzKJhiXaJZlNaouqP6XPLoWXJ+SgWko6Q1QBdEN
EoWMNPtPwBygH5d0Ui7K7O+Pqj7OXEfFfiMLkAYaqKusDrYMJ/nrUZXsCplnTomN
TAGAamNZWpg5yYUOVWWWfWzr8WttsaAFSpuyJHquEBggF6yRsJq0mZ28p4Y3869Y
7/0AvBFMei8mVADLQ8/RCVnNebqNUcBcr92V6+3+dpu8EYBC7nBbLfkcVAz6x3d/
8K90UEpvIa1bqBpJyWMokY8aru4OEWZheMjOSrzoOvfyK5FSWQqC7GeQo9QHbNkS
aycYXC52cPSM18BWgxfK3Fb6FXIKJ9X1f8vGJsFPmdw0+YGUuDU3IM+KNn3Q7Ttu
5hO/s+fGeXOL+zmra5G46NNSow/+EFlIb5iHy4Q9Yi0jmjCfMRH9atIe0GQCnKXD
li7oc7F6oyxEYSzYW1GPjGGLqewquitstOYx1b14mlCmDJ1yl9b9r037xDUTlFpb
cDMxTbs5TIHDQRVZVZrA7lNlbxnOkV87CCRPK/6E0N2TIGDSVcc/3j+xh2HKIwm2
Dyj0E5nhhTo94a0c1zqOFXSW6UO+HPindz3r6Q6sXvivWP85OVD+20X9FUxp530j
HePwook9XmxWgwzGj8D9wj0dFMGVi1B3tMbUNXtwq/QEexgRKIgDOiOtXRIpVe8v
O83kW/wF0t2iogpU6k+6kizQzTZMfJ7oxIZXe0IgwwCJH9n3khc0+IQ8AJh+wAMn
EesH2bZPvxru+U9q07ZWqyPffCgMnsTrusz8hWU7Iii9uGYgJlV/8XFPd8NDykbr
pKvJHe2FVakEpPM7McF6VvRAow3/dNHgc4Mp+NmU0uev+m3wyqVjMVBK8tvsJyze
uGgbBJkqElT8NWD2JWJU3w6iYkO3CM2r7sOCABS1yo3CJDZGKqIErAgI8iuhHUSN
ivAngbg/mf8n2ltoOjG+9IPqFzD8eOz4H6LdjBqzz5mtjTs0w0cCxQgxs2uP0qkJ
3iM3VQWv6SvTXbyLzUCXbrm+OTRKspOEWGyzyUbgaZHycOwf3L8eHsGFqSAhAVfw
7RN8H5BX/8hkP8XS3y/a3q1l46mmAnByV70NUc6KWegCJtvnEGIAZ20uMHf7zTDx
s37EPnXEKknGqFzbDvJhVzUIdqIgk+z7jwL/+EwUBzM/2XwuZJbjIbHPIPBU2mA6
T9gSVKFHq+78TkcxODLqFJnDA1rKxcsODMkJbL3J6P9IOxa1l8504F0lyzenxCXk
RAaDED931gTw2IeSZx03RhOWKHOtjUsG+N7vDDypMScHpXx1tk3HcZo1NwZRD7sg
oGn9mva/Lb3Dyt0LkAvjS7opGXs7ZYpYi0nJDZIGWazBCmlRhGz4emPGdu+nehXV
2qZ8Fl/kuXYWD4Y3NKh8juqgiNfyufaNnPpjXIskwPwMjrYN/3XAv4TqcYyIUJvh
EwbMs7gRVqfOQvtaupuixJCEnElMRfTdIGcnLDpykXgsmHEVNCZ+YUXC2Cccjwld
Forazs2ldDF8ZxkusP8PWQPljQUEUOSEDTXAS2HMiXmgLP437IHSOxAiXfqk9q1/
Ip0H4h8JKzkJ5HpF94z2AFOAI5JFQS4n43fuJ4ULO+jf2teLFRZfexi7qMmA1yVp
UMalDN9yf5idSwbI0IC6vkjhGfVqtZ1M0CPhUtnI7P2Yi3MqXZg+7igeyHp+o7/B
A6byCjiooKdR4tcdG06M1sXPXH5ckHfOempDrl/tcw28nWWl0NjYj6P61K2xCxMt
hYJQHhAzWKTIf+BxoH5636J8EGuQqheK9+qxX6yEN+zI0AGTerOCOOumqq+balt0
lxDpfjm+1U0t9TOLN8pjt8+hvAGKVe7rxJ6tsQZn2MOF9nooBdMcEXi4wfCGsf3M
8P6QT2mTjzjZ31jCshZV/6SQMLWzDrffW9Ou/K/rj6pOBazCKys1BRCnFeZkiRSe
zdRzyonol9ew2Ql/j1L3cfFqLA4b7p8/IeYH//6ZcCh2RTcOVm3qlA1EKOToYuxZ
0rU87tYIh8G0PsDXNFkRuK6qll6hRPvpzRHtSGH6gQ22LZGsr/Ai4frbK8gL97r+
nvh8Moge35hqlTzsVxBzvnbS5D+dDMU3IQuMV892NyzzQKNl5BHjcExQeTpUgyJC
WbAaVejfI2WPCY4vHohwRq94TTa117bJoccozpVae/iKaYSPUfx8lfQ5DkcsObd6
rKMenv9ydMEooqmVtM7f5A5FVbUqw+5fOZBZVxN8kjDyH4c1H1FVE1xydXj25lCE
GvcNilWrVZlAsDUJgptGYgg0UOcWpOsHxX8/lwUqSqj97gKHFIb7GHXHnnFw3o02
TSHDAo4VLO7e+uxByaKs5ul8pQS11GcxbASVgJUdzsukyQ4eIpvsrK1KICEL9p9Q
2xBE7WsCjh6Gt8RNkhJj8/BStVTtG0vnzG1GTzcwIlRsaAd8NHBCi4aoX2ATHqKs
GTFmGiqDSb7OqeNCEXafXd/O8c5dewpTrEKUZVRKRXeMvUfqjziPXPQLIOXTjtxn
PfZptykstjPhT0aGB2YhrNLNG77Qw7eOIxHZhjNiUvt4Lomj6Ppsy2hv9MSt1sEv
kaisv2LhXrLUDuPE7EMGFr1+rFbF2wewB47lAAPSIBOt7APJUooUDwh7I0N2Stbd
yvyypDyFicrY9mEbLd170xGuyJCihGM3TgZfXoTXbzoZ2krQrNWMn4IXZM/THs/g
MWjUK9aZy0e0WSRN7f3QFr/r1VOKdOp24mMxjYmPHxUqOR1rZkT/30urwzKj5WYX
4u+BfpOHgCVqUAA9seW2Xx7WXIdV/w8qXh+OfYMAdooqToxc7LXmNGAq4E0TLyn2
q3dmYikmk5cPXL5Q2veMIs5URziW6CGfsug9T+bvU2IhG0M9rHrOJH5rWovPZTzs
qZrKplgPImfCFFC7KOMyAm0ug3n6mEmYPZP7hrn+xNkEg50BsSoRKTadqxui8z8i
VcIMm5Wyt4EVpQf4axfD9IeuQQgbP3ALn/jFmJxZ8aFJCwQumze8W9TnF6mnNVfa
A+pSN1BSAQhAm3dKBRLzfXbBOdDpTmS6B/gA+jW4QvqAqiwtiw+OMpyN67SH1fU7
1sLxCF81ErK/P1Vn5Iw8jD6zEC1GwqfnkN00FSncQodqlXF2Qj5HgCJ90MVNMWPL
taEZeJ1YK7SfscTMgs+3dZHDxkT2RkvryclxgTtAmhmqs88+ueJ9YSeShgqrjV3C
Ty4XX2z7WNzoKiLwtfpSpPK3MPq8vD3yyX36Yl56EWWr2HIR4dDzSwgJ1tQuMHZv
gDhA0A2cQe86HYQE0rR2jRMOImcdwAT6h0YSqwh6RgOH7dqZIueaiO95KU1h6AS+
Jo7OkQp70NZJ+uKJDzNI0numO6hnKcdIjnU1LQSWzWktAg93afDfo6QRTd3svf+W
/ZU17mrSaL9vG/ZXPMcCsYdYQuhyEuwFp1y+ryicTM7VAOocKj8Sb4ziQ84E/B8A
3eTg/6p07nJF27I3yEsa2DnhG8sImmmH+Ek2HR0AXI7qE4a5saa2EXEUWnCy+Skd
3Y5E+N98UBHI6obUnpDGglvK1BENHkbtCtVLHfudK/XL0+IPLnYb7PcKwAoL/wy8
f8glyysky5IrdE9RouO6OP+ChCkBTBxVwK8wUyTUJ+6b6iT55k3p9Y7bLPMzBVDL
532t3V2b9CA+mB2NfO6DPSIcF1VRfyifYscdQqpd0xNSBA+eYNhT58o4+Kjgv6xC
mPr+xWbZXhemTtTw0PRtS5jJREGOnaUoc5w2nzscmQSzISfDOQh/9HsP7N2He3xi
gAT7bDsFxOeqPLkpF84pFJSljedhXit7y1pZTi634+RKLmf1nj+UcH69jdVdXy02
TW1qVwiKM/GYZcYr9N1DoVT57xUMteX08Q+rP9JSOxBf+Fx4W/lq+zDzs1nQ7dks
EZzOxfwDfHltKkL16DVMb3w9pVSEc5BMSutAlIr0deBBjiH+qghVNVw9JYknhMua
hUzsmNQk8Rn1w/c0jU+2sNKqrTAfOlCFuFMSR+ldW6LNIbKBW50KzhmBoYwGEOpd
PbvVnXIUaLwlY/Sow5sQnYdD0tsoAJO1mnPHA3xh6byEXkuDW2qp43bXkyFkCF6i
N8PoR87uUiHPTbKhqGroamdd4TCGcpCdQJAtHYtIteXKrw6N0dwcS97SPMK7bqPG
QTO3CGuAcTclWZgyuEbGZJzxH3+lhQLAtEVMnpa3iL0HZ5vlpCTt1ajtZKBKX2B0
kmt05PUuU5rZBZeh8pWi5H5EdwcufIsWLgi2fLgAOotlloGPr2LFswA/FVCU6S0b
rbhluVabeTtziXWsquj9lefHqTt0VMjAeT5+aFhlZR3inIMLAZjTVPmdUlAfKujz
uv+W+nhrFyNm8nu5bEv25/TqtqCtqF7ejW35t8aBRusrihrtFkDN2NivP/k8vyGP
+rROaDcybkJ4GEyzwt7xsHMl/9v5oc7rkWtLOlf26MKgxFViAIMR6dznNJhrzaV0
BneH0XR4izEHettyO7J3I8dVUOtPTcQCiI6A+Q5APSZ9de13MqYH2CNiwUyE2Isi
cHQQ0B1SmWGifyhM4Y9fywGrcms0EloCVLrA97ocqCxjrJ8IneyYEgrBhVs06GyM
xIByPNQwJfxsINDeHIsvHS7yXPsqum+UaEcgBRkH20YMNYR3xRwS1mc76e7R0myQ
Bn6RvTBdzJTNdf62x1eAr8JLL15wLWeG4Q2Ad0w30ohE/IoRVqpPlPRM+Jw4MKeF
7UbUscwzEEoCPHqiJ+Xe79buaZaCcHL6qxvjU3g1wTsFCQca52aCp3gZf3uYq0sl
jnGTGX3T0TbjUgHmOaWB86B6AdxbOYNfNj7h/HR5TKpoaWDkN4pbKb6yxxjePQnR
qmwmdFW014ZWNdTjDP/+GUP15iLlvwuO5a4YH40OXB7au+3nnrpyalbXQt0EMb8Z
n6POxszE+9pRnBdMxIdpPS3hrHu0JWRSSxPdAdj3lMjZ7pC2kW5L1m3u8RlLXuQV
6G8dh5x6Oocpur13g+Abt+HUdSeYrjJ0koMTDG07ifWT1h0WKky1YQ5KuZnIew69
a5bESRSxYOdXZjfMtIjUzuLd/WetVH3RH9f0MzPWPkeQCPFEjEKAWek9XQ71wBL8
93il2Fe6ATq5vGTdginOk+cVj63ssr0ntzuhTTg9MKGeKGzPSlMOZ5+OFFBlbDnl
3SFTxpKERbV6bX0JkP6lpD4nr//cIDGriChL26cdPJVbgPz5y4sARPZPXPCqmcg0
o8TrOE2cEdgFZhmqu6/X8xE8aTfW3Fdz1lX1DSmWOhmvvsWkqWaKVHeBmtB4Xwh7
6F6V761MA/paPTDhvIm3mwAJcpEb8Oof+xrPweLKa7AzHjlUt3nxw43Wwuj1iu4Q
rf7OlCKw0cL9A83wLrgTQ4Y18lDk58jiXDj89z0E1mhVBrebrEElSzFtaigBmHPA
cHKiT812WkEf21rYMDtEWYtkn6iE1HVlJ3dwtGI/Egjlw4UkNfneRgWPswZtHw1b
VFSiYfkziJ+QsdIInFLcGu2exW5BmVGs6bY4JFCnqVu49sMk83PmgijlVZmU0RTy
bRin8n8WyaDMEFMFMvZEQR5ITORb/Mt4WTfPqWxxTUnPE53KNf2O/sKoRihekvyo
w5XRCczCjx+2/MgjI0IC573Tf1GNgVYETx2CZBhH/5J+NtglmzwNiHg2/BRQpiUs
+F7NSH2m0Caf0vGQbST9wQCRGoEdHtOEviFmKmO8jBMAmxQ6U6+bbbvg38mMnYUO
wb/Mz6EAQn3CgjhQeQx/19rzSCV+36YCfMe2Kyo2/Rka7DP8XSUdj36f7ERpeZ1Q
udi/CpCQHAojIfYQScST6YotHSIagBH0CCv/9Y8pEpJVmyYAEIkiDJlYkc5Zk0NZ
7cp4Y1zhebs6MI9NyUwsy9dPZXFahXiP1wDNLcmkb7hAYPrbywJzfIq3VLFFRATh
GjrzjuvUgSCBDVq01g+X/+o/zYMyoybYDT/Dw51LB5R0XVe7dsgdqr/KfkdyCO3E
0oT8iAJiWdJ3ZKiGZzMbpju3E1YF798wUO19sp49ojYIf2sNRRZODGhOq6oSNWR8
1WqwQvazmyKJPhAWzsoW6HtPPxsF7t6l7P6hmlP3lsXYywm19w8XCKJppM4Hh+Yd
4sy543+kKi59LAjLLQdSJbI/hF5awOEukbc+RgMS2kznT+osd+YMH2fsXbqyenl2
1Eei4t+HsRTQQG8ZpSgCBeyPrKLZusOQFsZVxQjT5I0WfAeVztZuyyEsJq80VqbV
30nEbmtw5yqZBHwkK+8XYfpiI/kQFlZ1RPTaZqRbCrQD1ASXiNB/hQBGTuhBZ7nu
p5s1Wm68uSqIbciH/d4uglJAsXqYEtacMQDBdlc+AU37WFDbnPhTZSx941H4j9D7
9EzThzAK1LRdlyzuD0wMGS/bl5UAUJ6wx0AfLS3TZ+JKcS6NAhIeaCmB8lRg90uT
AIXNDokvIhUJEogVJkAgtUtAGXzLi6XgLU14EJj+hRMcaM3OJ0xFqkeNk1hX6pq3
FRDfmlZitAXXFHn6vqlFtsIzgG1z9a3HBJVdkylevBUfWJXgOKu6Fy+O14DJqLgv
tKzffLa7UbUcqF0xP+fyqFzXJMq/sfDyAoTLf2rxU5ByZIFGzlmF8YZlbAg1Iha+
12KXLA5wUTXpwP6+6Lvt5q8UEmtkK8e1zBYv1J+MbZg7DUp4VMqFfs7oTJEp/NQA
XgbxbeMUNeQ7FEjNbYSuf7kie81HfEdual9mZ15lx7IgfgLmL4c9umeIRIDV8hHt
h15rUPwgHoz6lU7uAhMCaZ6OW9MSgu2jY83qTB4pkr1hKrGRI8GReaL+jhSfZgh8
p6mFkl2prOtGDdAfbdOQmZqGFAAzPyMfkP2oV112DwbmP0knzAj/zLEnVH8rbd3X
3DJUlgnGQPnTpN1NpyBDDzz65BiHLBqra7G5f3bJrd5Pv4cU4dldNPr88bnx2F5u
lz89lZJVATDBlXnDMHENrhwcKxBXUnpeR3AlWC2fiE86BHo5i3pmBr+PPwUB+ri8
3z0hyeYrZXd5oWvoC+nDwNPHQYSp3IYola/ZWfEXUvAsojEvstyfDdFekEljcli5
7cg6TSmxW6s89Txyyh05XJA4ZsjuPfViaFoHkpr5ISFo2g9lQbJqEs7WtJtwgK0l
5sFBGd4Kg8afd1ny9sdJi5ittyjKabumOtKI/XrdYy2BOdDAfuKMv6vpkqoHXfIq
rQcDUsMhGWYpJT6It+lKDZkFClSGAqp9lWV22iAAy6x2uxyQKtwsp77KxaeHMfCd
kOQsU/xoQT87ykW9mb6dt6XiOC/cs9lQguI/9/aj5E8GmkC4jWGgHdS2N0QuRSY4
NeVnUi8VtdlpxnanRxcnYKjJpfe1opY3NKWfKPcFHS7W9D6rhQzNamXfvD1cxBw0
klMag25poXephu3OIi+XDX+ZC/taOb5zsTUH82hc2o+jX7JM4bvMIQ44qbXzM2ia
Vtp6jrLJYtjHxqrzILFd+/J7UI6+c5jWQzch4vHqSqelH8OKKetvmjthx96XElGI
kwv6Y9Q4ZpEvYJ42nyjs+uLQ4C5j64olVZzJLcAye/FmDtLOqX2GGkhN8YcoUq9C
1x5haX0fBJfiN0hEQBqnr/2t5z0bdvexyPWdjIN0WnBPNjcbKSMWFWetE/YPb18g
g7d5+dlrIzCRJnn7N4BjTX9yPr4AWRkpKu5nN12VS4n1V2zHwL1/cq8zwzG3YgRQ
d9Eac0N7ZK2auCcu3k8dSX9CTd3mIukMaxCSfCT4r6hQX/DzmbqdQ9oH+UBVEMgM
SyJipIGSi5j3mPOlYF7PyH5RpHHP4p/46iIaXwA/NveADP4Yep4NDOeidSGAn9Qc
p0GRAywumWXoA/DTvqUGn4kbpxQI1EftF1VUC2Xe3Z+jJ3An0uYit7x9YeRhH7tA
SJtAPK18auTwtVld/ZmA9aMgNf2C2bt7C1C0I3omf736FMqMMm9b7PF2U0Gp9azD
D2InOE+/X15vyj6JRlRsgv+HUNbLSQNXPOle7T6N9XBSqCZ7AzMp3thludAPn0wZ
prP1G8ddsK6e9f5Av9t3iFqi3X2S83+Kd49Gbxo/LBrI2t0oIVdrprvHhXCpSta4
PUmXOVmpgEJRcGb30fMYEjKyRYALwZ4u4nveMoYUAMyK0LWHIAH09hlZaBiwDMt0
Jcb/rdzwVbg0r4spg1rSNlO66ynYPkZmi/aSp8SxV/w9jEPvg+jOj/EiLpDanctH
DssANza947QJ0FEzPosR3Jk7SKrftZOXc50yKiPv6shrR9fzvpwzLpfH0HZR8XU3
o5//8OLDcmAEUUyXY3RAf1BtqNQAUP9DA3cWy4GkKgz6iHWoXtW5LFN+kZBMw/sf
f82TdgchOh+2jZJLiYY143pZmV8Lv/j+uHPcTaATxSR72LRrk3diqCQGZxTswAv6
VxcM5duW3CDsFX4BqxZKQ/3EWn+AY9rCP+eG2mKXe6JPqZviPdOXpfklKKJBYdLe
iuOnjE1HaCCl9gxGGtt1wiD9vEHA7Ea8lDpePgBuJneQVRYgTA+/JhnrBzYBECIu
ybAZhCRse8s4EGfeVsRWtz/jhYgi9fCdHHCweU+IKEkqGQqumvisvC5GkBmy66jW
ULxU/qaPdWLSMF4AjkYigVFbmRkpU/NNvz2nICoFy9GxPoBz1Q3D+3zjCIOyiBpP
o4DhHnpk0LLuS0qugFFbXh7gmmLQXxhmynEUQTnZl3CCHQVPa7jhJb//jwuVA+WV
iWwVaq1uAH3+XDFdWrfWjsRnXATL6ZzXW6O6lN7PD8szmDbdMG9T0uOYK0jj7i2D
ocl0TOlest9Ky4bmsvmWUyCf+bfM3AdCPPmGXqXgBUPBde9PhMCpKz7itB8UNoA6
N86SlhuUVu1mVKg/HTaM+b+FzDXZ03u2PZ8uMIwaX5BUJKHdSCpMO7dGNVRcPs4B
1SkjZdoDsoCszsbBtMQh3qG2eRuJEq3OQFSkq6AB4IpILBOvKIBMhz0pmDj6/Ug4
QLksm2ZH4wV4oeRAACyiTVQMuTl8bZpf/s2NZZVR9TvOHtBe2KCFMUjZuvTDBUFY
U3yptfdgyHFFPW2pSQl3bUauJGMch8OdUqyzwidDkAnBE+UJXGF2zXm6DP1MqMRb
prw3RiqkIxGYXxmX67Z5UxWfv6zuro/wO4ovldMql83NcTvtHHECKVEuSZRCs7QE
FYVaDAisMm483IJOs5+j2oVD66mnMOFWgQ2szDVEgGwvlPnfHeMk7jJpUGVrUsvz
FLdiKBStW4yaoK1B5HzsBGA9aFXQbMYHesX5Y86WgqI=
//pragma protect end_data_block
//pragma protect digest_block
HbWP86HKzTmKKJPXFdTcg1sfcig=
//pragma protect end_digest_block
//pragma protect end_protected
