// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
vZczFd652f3PnaEPG8iLBLBD0x0nRm24u24F/Y28bB+3aRNp4AVWhVhfen59
Uzi5sKMiu+6KDvWh+qNwDHWUxV/cwnb3wYNNRCY6BsCriu+48BHzSniCMYES
ToH8bLViFrULrlaLlTgUUYHghq2/PFAgEVB9s3t8coEOHZedBzFZ+RQKWp0E
DpUkqUWDFZD1hiFhbx67KbQfuPs1OIaug9CiCBm/aukXFEZlAptQfKzK7xrp
wM08Rom5B54zQYSYOq10dOg6fFgqHQF+JlLCylE4X5YasgzWd6rI4GTwi3Xi
jbFPvUia1sugmvK3OmcnfxdSmxmLLumPUU5KCocypQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gLAgPuI5dk/zirnMeHxoWEdmmWcbUGAFcH+XFembGUuH0PBQeaW39M1USoMj
Ngt8A67rpYWhqbEq4doCPGal5duNniOLkUwJUYqn2iKW7FX2Ll0MLVtDnX4R
KOVpHxXlfJXJ8rGklmX7CGq5hGaeQ4BgjBmk3a4agSBcWh92xy58Vi1Ub9w9
tQ81bxHlwaDQV9jn0015HomnQdOCdlkmilAYXmOgXQ5prh0ylp5If605J4de
nIJ34dnnlB4Ul9P6xTtFfEw4cSyS4n4drwA5XtVYRqeDkyxcsVuTXg0gv4IL
TKhwpn4Hmj3KVA26xL4B3e2Ll1Xztk9xoaodOzxd7A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kuG9/eHwPBuNA8H80mFUJtp6CncnqPBqV3tp0fePyL7G9QJhACg3syKX3Ke0
PwtW3IusMJUHoiXGC9U5JMTf/f3ruRAtJ5bpsqh9N1hMgwW+02BvxlErJEwB
pdRPAABjZ/WfaH4eG+2AZc0/lNegWqn6muabuYVbiZL2qfYhUUtKX4D6aI6A
wbXIF/UHSyTjhD6LgIPBQq+O1jxsm6MK3DEi7hOGlpzD6C0suj4/vwTDJNGg
rj8PeVZ+qP7oOZMnNYNzuRSW9DBnEjhH7aJ15yTsnIzB+hf4cnph3M3ioymF
kdjkDjjoFV5qTtGIYwblOWfGO4BbGfKq8F7lfgCx1w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UXn0i8TCO7n1haNVyVUx+8NZlWXa/Xl5bFxLnxAqgStGsA+hs/TlTEP0sgk0
AYdTH3h1aaBhXxHsQdsBJAFbFtoCYD5BPHE2PeE4afOmmx0zliwu0OwtuJGj
nPjSgwHdMUUshXOBm/307xBlSbsbHd9heKUpOn/zpwZv3khr6HM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mtm5dmIl/bHJI9nvVmmGoIg3sfrBrPR7CsJ/qs17x+TktQrlCBW7Xpszm/8p
QDgy25qd5AHrmQ5VzLUJw14dsL+F+WFw2/wy3Hv44j/MKZwbZpNr9jNbZRtl
55OsJp8eGbgUuhGn51XMDpMvAHX2b7fyYIWUxR5B2c0WuXv9bWOcZKZHYexY
i2EoUAaUDtr3hAwpQWoQ2vHXHRUUfx2asQf52UL0eRndJ2EJufBnxq0uxN8k
iW3AOkE1Pksx/WpA3TWSPB7veEz6EbWy1z5WFB4wn35qHBiCYPwK2aIXxGlJ
QFibuUM4/sL8c0L845TLCJu40+d1ZR22ZBwxOwep/bXVy2Zmg7ABCaE0VhSz
TPcsfaV7G/XwwKl1uRxCQOiNRUjyyYcEArWLmCq/DYhM2yHkOnrAHR2jw4sy
93B5bGkHquU9z688cRQ/NrgLPkd/DO25AhXN80ki51VsD3XOBCJo613Q/DFO
uSfWY+3fR0F6eKIzpggWJ9ObGQNQAiCo


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pnzftb9+n+nxHXCF1vZSnQg0BygAiddmiTbY6s3aE2udi2LRqMpLB1QVJTvf
iG8qWFo+aBHFIeoIvmepCmkEyqJoISJmwdYpefofbYRjknNWpb7aC8davhs0
HeJsaa/uhz56Mm6DsUlHeS6tKeeY/iBNxPGf7sSFviSZ26WGQx8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YhlpkoNiFu0Jz7GW7ae1xLzhtjz1wcGKVAKkFsMuuQleJlI2j1B1WRinZTM6
nl9uFsaDc6jSqpyk9Oz5R0U7CDMjC9OTXGzX7SXEptjWTHLLfk/kj4SQBhzi
XC4VfajWw2kYfJj2ukWF27bbu5/nlxfyH/T7JPeZtSFeCHj3O7E=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 91632)
`pragma protect data_block
2mYwnc0vBESlE4oCQuRt9WrCwyzebaCXkmgxNHa9z9IKBs0I0DTEK5kMZHxE
CeSLpfE7kGRtDhE1bbr++cqb8OHOw9T2ndlacnLCuAeLy/o2hAsUyFPBPdkG
RmN27wpIcfjSbrDPxgnzWql7YQyK7KU0NGHsrbcoGI3PHRUEEdoA2nP4ZUzU
6mY1ERynYXtSDk5zRsqCxZuPIYl3eWSo5mGYq0gd2ioNWOYU3zJStrlgNCjW
gCoqvnG0g1SppZ6/ih94FNMa4GUpIGU2Xa6x2JY+K9S5I5i/lgnSf3nKCs4I
iRIQ28WhQxf5Jbme5igmBPlg33d9lhmOD9oSm5JMH+ZeVSfZASyJnAzIfq2R
4k8PiXkULGi6AxP8jANL20Ogx3kczSdGXEvtg8ND0Dahk+C6lTjsjhI3aSl6
0ieYXQ5NloWySmjpuwf00oyHfRbbIGV9YcBvTPnJ0bQ8XRdJdO5G8HykUIWk
1YYco446a4tnruSpCW0Gt5VWN1+qE/EaNZoZbYWzH1VxdJl5sXZAeD+4N/YG
C/bm7P842IIvoKFORAPMNuZD+el22ZS8RXQV5yHRyx9fCtfOUTJWb5kqJSi3
1eIoSYh+JYO7NJ6AgDPifNTrFnLJ4ZxaF4ZVFBZni1OEelEU6pFqrIkhrbfN
ADbc1i5yrIekuf9YvC7DDqythuLxr6nrM9netqqdORqAYWYEt2kzlvnhK6By
NZJL3bqmG50XgX82gEjBPKqrBvSgPlUd09zIJuWtVqzEebOWTufw/u0ZqRbW
MgpPkZhfVxJtf54IFSymDifchcjdRPGFIubsgXWX1auLHn7DDhRRCJlkUvqN
Jupr5vAC9D2D+YeivgPv6Z+0dUY7szd6vH5MsoH9bDPnEiFRZdCsd97cjN3X
tzXQ2OD7ZQb4EnomUfbpQR42nBGvz0uN6h0q6bqeq4ET8Zu20pLGwrTWk2DG
FCgtIiD/+x1n0vDiWkwKk9saB0pohbI3hk7ofOwTH8BdBMqFdWk0yCVrffBH
Jx+LA1sVsEDUWZNuvCQB9zfotEKBAuz6+i4dOj8s4yJq85IVfcQfD9okzXXv
YvV7Nh1an5Y0d7TEeVd/NS0qWKJw5IIDdN1mk55SyA1S4YlwRKpmQfF53nZw
3br0gFQ5zpdR3K3it9Uk2Q1q+Q06s16hsMhs0VUg5nx+ozmzG6KBRYH3r+ou
Q/uvvQwiycakn7+VJIbecb6MFS7xTK7MEjF9knr58HQrbN2IvPOF8uWb3O6H
V4AhDrwPfq/Rc3w/86U7tocEJUT1S4tQkswfvBaW6uwP/LL5JJcyS9Glj+cE
I2FkNdC+ZPQ5FoSjp34TdxEFLZJl9aCwY5lRT5MKEJgiYyq3dgVfys3424J7
uuh1NssVN7JPD/95JVVafNrvzChmWmmQjkvoL9mQHTGWrPrxTpC9w30U9YaU
HHSN1FgC7+PUiYEEiqaG8qhB5fLJl69CBufZRxsfItoQr6jb2p5O85z2ix3e
aSi9N+B9/hQcGoqf5hdCEMIsDQZAL72aURuhQnV5kVOaFV/ZRfzbfG8l7naf
jx/DJIRsr46HBQvyeutJwjmrif+h8r1yOv7d/tVPlNxOqcazaeZAyS2FPEms
n53rAGsrFeLNFP32H0eQEPdiiSc1bBMCBi9lujqX68GykPNfy/gnaT69wo2P
Bv0EkfdvN63DoqGdvRSPwbso7k1xz3aqxcu44/zO+4pwWXbh/MOOzoQJkh/8
+YxkF259Y/WMc2uDwbGtgQS0MqjMgXYBVDLbK8LLrBHJ89BGFdzK3KtGndko
BwPAU6D20OvoencSZXGmE77tkGWZeawVuxLMNVAb7xYGnPCSL5kS6D8TMvNf
lInZ/3DSu4KlSdU/Lpi9g1XVgMzKIgJeHcO71N24NGAEEEMM8uZ/rFRslLXB
eoxXcV84S9LaYocrnWqav8slL9IsCT7jEh3XPpQeSb9BAHrdPoIR7u9xKcLS
KywmprNaoktwxiPzHRcmALSYdGvpYSZphAvXKUYbWyPUEdGCfEFeRZEMh7WD
/mqPmORtDUhwoBiXPzq4fT1mkfIjP/DCt4s3RLsgdefA0lMflN/MiMSNC0rF
rXqw1qdwAImMTnEprEG7Jg2qyDJoUQc+OUSHT8cXwAaI+WmVeIKJEKwzbEF8
TBaj70wfSVsfRh8vwAH/NrcIY8mnoEs8BxITJ8egrxn9BTu9SFgYFngHDLuc
1pbnVCdrLsR+uWaXSJaMIbd01HaItdsK6Tg6EWQ0sl83CUMYHuXh3QmyFfBV
tYOBBtg2K5KioDyoh1B0cltptNg/abcy+8+w2g7yUHgA38zqc0hLL1A8+3xq
2oBqVDW+LyG80Tg+spWFIswSNpbmHcxHmyUBS5Rf6OoQo6YbnytEc6opChvY
b/G9+07SYTsyMfXGxK+p7RnQsRq/apbrhwMDSxi+qrHlUTxfYjj2cicGlcJB
KePi7jfPPrnQJPEkbJKffvDWR3H6lugpNmAfvzO5vUrQycW2SCPMTqMqr0/B
oXV/tqUy3tO8HujaLEneoxLs0R8eZHAySinc3n8F3ata0DsnnJtU6H4LinA6
bgjaHzZ7e2S7G3PTPxDvlbJUH5LzWbYSsr0NjUd68/olc1g2TqDtbZhix2mh
/3doxpvlY4LzahCCy/MInNY84hoa7UQ7aGHko3sa9IrNmEVsfI3ebqPkoP/u
0PQdVkKW8/o8zjELl8TwIDHf7nWu/fDhioBTt1HZvwhenKS0a0QQZmJa/Q/O
InxhiRwQ7lbIPpHQDG2hEVQ/tfybGFF6n/0T80FQ7anrRJX5U92oFue7hHCs
r1GidZTbrwRjVGKjukD3/C/gMjPqeEM71GY3iewUG1/HGPv6x6qgeEhTSZZX
qITng/oSyTXPKOy0cfFOwTjnzIXGz7Kj9UB0zhaTGkZgyB9f8A4nlJfJvCu1
ZflMlmuQy7GubM7qVQUsJ8p0j72PMyY2LhmoFT1UyuaxoIdy7A/RzUywl2ff
RFv+oRK1ErnQQp/TyLiX/cBIMTDnk5ihll2zrX7Zenrlcgu84iswiieIKKAj
clKq1I4C3CNAtA8DSiFUE2RJqX/fs9WcWLPlC7RZSaWfvIt9zAuCF0RsuLK6
9ufpRaRstXThajEQjoViWU5Gvmcbh06rn3FY/wHWAjWQCBu6/H+rDE+GgOEO
b5x33l2p2iOItLsW/eQojpmyLzrN8wl14S1tPny0+wPjLtahYx6sQ0A0mhOT
yK3osPbwPjp2iSjYA5hHcDdrZDVTR0AttIGH6jLOCI7b2cDW2nGtn0tI7T99
eoO6mPQyjxCCRsVnLmZBEIiYRnOSi0Qs/6KhGAJn8EMbnwK+ae4lhIDdyOXQ
qNKL+lFWVYnE4b+vCwhF24y3G1kjqVaCcbSZf6RsI7unHWhJX1iZ3fNbiKLB
4M5F5oOOB2VwO8gFjZBDwi0UOHFWMylf5BwpP3xAEUacujZvFdBBAs25/YkW
m121zJmHTzfvugYdszsB52XBFosxoZFyqlYzcXjbf4obaoOf4ZUkgfveEU/K
rW0RIZ2rwDZFwuaDafEUg0pkhfucceFya9He0krH4g+aliT7d0jNCqvQL08/
tTeFNCZGzcC2iYhczbxha18r4NboPmwofDqh1SO07GayFxt++PWjYEKhZvau
adKioaXY3SFEHMDd+ZjYDTG6c98Cji4ODVlWbxUMLA2YLHLlboo3W7p9NWU5
zQLyOPv3kSGkheNIeowAITfcBKS8jkav9xgPqQiEEXkwiDI5coWlTrYDY1/l
YnPsVTLa9YcHIlTOgH8EVR6GtPlXqJrDzcMcUURZ1OuKtug3/JFS1hgGzS/x
rvGZDvrS1FcxVKnvEXzjzKXwCAYwqwWiXcsh0wb4M3DLnQCCWf/cIV1wK6N0
XSXh6mbg9UCQEf7d4YrOfVKNX1x9+D3eiKAY0FBxxVZT6I1mRICfXbs82Rfz
AwICjtEAe35Srg3fCunDUg5syz58dHmOtIjya+m1L33RdSKhthawKyZ7wCYU
zDSCFGupKcehNARwD8325miK9JLRvAtdWuwzpBXF1vPLYToyMbp4RN0Lm/ai
bjRo22tqgTm9zkKMR3XrqCCPHZjOMaXNIsyUbDi/23OMjqK1ozNUD9kOgV4F
hDWYtXoVEXezHPk+2Eajr+KoKtJd1ksiTkOfza5g8cK08yRwJ8WBM9loBoZs
7ZuNIv1j+UYWYoQD+OkIQ2Iy384MLyxDNraiz16FM1yIK4u3Jn9F7cfs/iOe
HjdAXWIbcIoCRNeg1yXGUO25mx/YcOnAoFvr7+YjWeE0qZ2F4k2qfyPVAQvI
mMk99sNDVOVNloIe3uwcIBmrGw/OpQxb/pDPZ1kswJJsy5wBtdX73zXnisEo
u6HK2fnl/JmkpjmOhXt4qyhXf/8JgjjEdjN+yFKU0HAUHEokx3CGlYMnZ6VI
w0oTAgC/QLse2nd6HhOFDn6UANHa632nWEqGWOauprOWZErudmJiRtEK7/SI
VH2Va+ReT8lTuR857zN63vcR+zXqseJZfqGWR7oWo7u24MtG78S6mzKt2Ie5
cGvjlsfIM7+8LTJI1HjaO5SgW7CCNgwlsBS412e695oiuOEKTPY2MuUdB6zn
ZyRKP/1RDYxSuabtVUtFZx0DD8UKlWDY8uYKuqVtfAiODUQro6/FYzRuiaDf
bvX4e8kuw7fo5ZwaBx5EgPY76cNh+37wiqeT80XaH5FGDtorV1Q8ZqFmA5DF
LNm9r81qKUE2mgMts+eQyWd7B6w1w/aT4QF7sOXTEZC5wQRqjhPBhyjkcTnG
Cc+rNu563DpbTxJ9aHnXZ4cZtb5XVhgODS+7mHLJ8OuPUhPxhQmL/SlC3tRG
OUciDndjR0fL0Pp2avpn4OcDjMh+MJyak1ReY2TgmGRKTGxGqXUMbQxxf0Lx
ts6sSvAFKz4zIY1Ietm+HTUSq8nnWwbBi5iSLBd6otyEJ6jFiVIjeCwnI1E3
XLE1Phf1q0YIEnDNizi5u2edpbeDAHv8tAy62oTNXIjnMXJKIx7Lig8WI8R/
Ftd5DN8vsqB9JPd0SjHRYIg6/nzrBJ3al8i+F6/bl44fNhTxUwG76ChP/yiB
DTWuh7YpLI9OBgDXH5UanzF96jMQAmbURLc1qDKARIpnLnQqhM2ySKdkFJ/G
Y1oM/kW4A6R6uSTlQx3RJT8oI1abNUvqQQ8gs1xCoxQrOtiQ18IC2TXkWjwW
3kEq7kOOtDCVoKgY3uuo5eTzNXc/Tc/l1RVSUnaGSePBTRjgGHUsIVRElDkJ
MXMh8Z9bJgGW9W+AkLXoXyLoD4vhHMEg1a2+LLE6vTvBdmOF4G01L1zdNcZU
Lwq4OhLVtAIsQAqcRmrYENSYEL+aQtomQ0i7LXMTFXj9m462bzdBkgTlUOzR
a9wnOfrRMW1MK8ZtHXxrltHGyHdYvWBSmg7LtOzkV5p+vKuT/sSXxPTVKk67
fA3vkshYhnrTkL2JngsxLhRrQ+0d1yw0ZIIOXmaqw0GXNBQuYjX866woJEwZ
g/PzIY6Nir7PzKUG8yZFT/aRTHjYbgHxl9UeXC7q9OjfzqfXDPKPUnLSh9ts
M4rKEtEiORkRiGdygtb7LZn/3+LLobyvq6RRDhb5v9KAmjuTFlI/bVYIHCHt
MMS4Hz8iZdGYFfHPhKb2tzR3JJ01L/RvhAEJm2JwFdisM2ZCqWzCwicDsjjC
Wga3cQzqvF5MGeohfG4SoJ4GqGv9C1VnOWP6QoY+KIW//k9jOy85c2gGoMCO
+eYX0SRc+OhYPruOI6lZE13+C0YW62VyptOhusUpoILcL+KoX3HEeghncdEJ
glGxW2mts+H1Ndd4IVb08Zfj7c+vJ8IvKRxgo6Aep83rwFPIQVmmIvx2f5f6
CSVcrlfu7/XbHJllFzOHTFJs4MlcPhLk2UZmD0yQLuqXB7if9CdWw+Y+QSGQ
fYkY+c+RYnd9uH8uw2uaasyYbvtQcepQqkOCUI2IE7FzOXgqawAa6d+BsGNG
S5ldy2A0AxhDgZTRoKOsnDRWXu4PNNcVsVc39L0cVYBInWzcQsqg6TH0QOLc
cbJtKHGuEdcS1t2OQKWCKUsUs0/ByOALs62zSoPr1ODQqQ6ZNVQcUukL5tvd
iGV3DE12S8DMflVbFywuWlZjTSUybhFoVWtoHniVmvyKM+EcTroV3NjRzA+C
TaQNkRQm5wMSw/YT+pFWL/J83xCQwmImakY5Itf6DXOF4rRdDTtZicZKDhF8
gPZQczf9oBSbrvJV1We0mUSID/yT3okClmybKu4grogRtQ+GVHMqsHo6ii6N
bEG53+cAy+lyj5Xf9T1hzCnO0D1/9ruw66Kw+DBsbc3vMmMWvg9JKJFubi1Y
FWPAurQMobMn0elyjJ8+S5RFB7OOKrGvH/PioKE+x6f6LimTfa/RXeFe+pLa
PFVPj8aH75t6Sr6+eCsHuoR8ScLc4rj0skzn/EpnXdofwUDy669q0/O1PKAb
e++J0pretgkeK+zJzjeCKLt89x0Lqpu8/cVv7cySN5CmbIMLftgUqJixC6jC
ysYNj/pBCE6DnK56+fKwID05qrLU94m9fq9vCaVaFyu+UQRHGQ6ZgBMnT+ZJ
I4R5Bx4DibV91P4pqrmKBZ/agiZsQCBK60/AjLUTHNnEiM1FXCDhjwgIfnWS
HvUg0owoAfu+IzI3lJOHA3xOr1yM/PXRClzLWfMYmxVx1BARSz0fyS4Q3Clw
9+NyAhbIiKHtYHibr6XtMvsAxKmjXK7p3muBd1r5TepnQR2eIPy0FutTDxHc
ab4cYc7HoOEHlFvjzdUUGWjp2/d9kPPmYE6pU5UTkaNlkkUETCabWT6aLE5i
MlpNWOXtgPXM6mF8G88xwnfRleuFLAtZslfF7fyaerRJUQ2ZYtoCRwzvT17r
OKamV6fE49kmeYrpK9huhDxAiJ5F0jdgzjRHGKpncBgQ+x/nms6TW4a9y+ws
OhSHzyTk0vbHGCaMfcvK6W3hkzrZV7nHJ1pgpPAt/Q5NryyO3C0PRpAPEDF2
H0M/+Rs4MMdzm98Re7Ia1a9TaW5BP0huIfn4gq6FjdLcr170xsPmDkB8KYlh
62EzrSKu4uDGlvETJ2vtUVkvPJNEqaXOaSM7QS7QSRO/YznJjhblNItSGPy7
XsZlWKU8OM/9dSsI96qr8gRPCmBevBadWkf8MnkefNtMFRGNx2nbVGZZpKJe
Fj2e35u2mSZRtMDIe65379f30aXzSR146uDxxr20mHHDX96uBSMbtlC9PIKh
jf4d8Wh03dgZsBjdfskoiQINis1f0lPmkBnwWwsycE+hDBB4az8xpYokEucM
pQTfTpTUqbOcs6Hdd7qw4ff4a7MKy+H81n1nYEGjCet5DRqjA08tPbZhDYNR
EXNlqTSb7ULlGB9GqBSWmSVRhT2NJ41VuxQ+GqcO5CkSx63eVTD/DkIP04dL
4/7DMxA9YmXw/ZIXoaEmUopGdu4eCoCQZ71gAd1S7Jc3/QeLIqE8m6mhxyQu
qb1KciQ84n/mqiJFhE9OlO4MsVpjxjZqL6WWUQeYxdZ7FvgakWhms5D0qMcP
cekKOpF1Xje5uxuRwferyboecFAdK/7xjLiBczxPQTU6RMPE+DZuHSpaBAOJ
MVxoqYae+A4DM1/AQ2Scy/AaL1pwxHVLiNMcDtz9Ztarrv8HenzbOPoy1T/I
fnoziWCjfuPsJzfpD2RjRj5vq0FO5x8wrbxLbz0mgJVR3A/isT0wLA4w5Czg
WM8sKCBoAyjKEHUNuch6Qjgakr9MJfFtoQ+BdvoiPt14Oyvpih2yp1P1kRlo
nrXTbtPtIaNjJ49HCSKnIQf/Yefz2rRGhpQSnrVfazVaPN0zANUhEPM68QGY
K0Tw11YXrlEOIziYb8kbXNNTDaC0DJsxNM8/9271C9CYhYMlmXZbyLw9ii2X
RCvFwjbL4H9dV6SXJVc9BZ4tkJlxrR4f0V3yx8uCrvKebu/yd4uZAl5N5hjE
NFkurYnJXvZEMaerIn3ShCx/DYpNpcUReHJHhNLinaam3ki34PdR2EkVJQNF
c8ZbN42gqaPtqmhdez2noAXuNqXVY2MiIwrp1DTAYYMyvEG+ti1/30CZtvVc
dCdfNNdddxlNq0CRYurw7HYyYC0XX7lxKYT7PbkE92CHDeUhzTkOFQH5Vyqa
sCiPPLs3K4uy/+/RwGkivd5WiLZr80+esEx7kp2IJHWoJAE03C2kWFmok/Hv
APCJqvxv4cjxGDW71v3M7C9qCxYd/xQqUB4dlh5v3NGIV6yFausPiLhIcNUv
dLNXdDqtta08GPCQIH6jIxLsQax2wopggz7U+P2re1HdlZVaq1GqYQbIb6Kc
s78bO+6cKTa0i1MPvwZrmZEFpedHZ+1s0AUVElMNkyqBAbA5FSQDf23uY4vL
rO2KAU0UdSy5QKshBmkMZKMFmkGHTA/bbzCTRHyZzu8NH8ph1FbJqapzuygH
i9EkgGXwz9C7DkOMdZxYxkliQHX6Mqg9kUM+1alor3yMWKyUjlp0K0c/x+sH
Lq9t/vLIMeZaBxXzf8/OvYzwP/wM6dEE3O8ZAzzxLw8cNS89b34Vz3aIiUA+
gF9k7CRNSe1w3VFoH99Kal5Qsmv6lTETe+wi2azl8nUAoszWwWoidIUG6w9A
/nJFXTophOA8vXDp+LUU34e3UdlY8fAeUityFO5FsTsC+gzElQukeBWNXKCo
YXtpqU0Ki+U9KbNbn7UhZO+8PYj4T9A2P67vltIFmBt/lhgBPdd7f8LuE76i
XlLyZD5Nin5pS1HeVKPr18W+LytKh5WrFd3HZ7/Jq4DEzXM+i4+79WMN87RN
lmcEeVKA1LI3nfMcnanjnIYRCrShOIfnPuiRx5hFnEZmOytu2+luhzOv0s+Q
4HU/0Y2IRn7D+hkcA5CA7xGxltYvJBMWev4Eq5NxJjjQl6p4NKcaawnQIxYm
KmSg6V1mgWncop7Q5+xzeE8Oc7GqpmdpUlUUVOZLNGsX3Y32PLOieEd5R+Fk
sr5g8nZUEhW96+4C6ZV1ltl+w7JjRJe5cYcGe1ldC8HMKU2SUvUze0FrbAQP
ClpYQFxmD8Uf8SL6m0qD1mH8FISmdPi0fprZ66UI3+CUxCf1X1geeO8Cl2b9
oGBV3XbD633D4jZRDkC+5aDtF75xy+GI01bqPsVXyUidOQYBPT52WG0K5o+k
I8LkQedhqtAQx/IHNLNoc1dzsghM3cd6ZwfE76BSu8bY78JUSVu+zaA7DkmF
FIYbzlOXFIOp6EeBfSAOubnThuS2Ydv6PT/305JLIqUnxFGemsV0ycUIkRw3
lrkCsJUY0s1JtbNAHA7a8OtoO9oxaB1UD+Ivryb61JwcX5916mbvTf0jDER1
UecbIRB0w10UTWIRtkvCFceksYgosLqeeESXDsWlG7/cvBmRzQj2J2xthSpL
w/1+TgWfvkBYJZb5sFs7B2MlX/qeVA89VE/OjmE5ldijBl4TWfKrPkUS7som
i8HcqQ5gQmK4vvYWxdmPJ53SMtJ1qecz0Pzv5BrtqgCxffMlGOhy6qPg22IO
3o11xlXv/dFUYLf+LUTvfZOLGX5dGGnkdLxMC3UvwUmGOLlUk/VHWFDUAcNm
CmZyEdWCDzIZ3icSwXSBMUnKri1/vNn86adHxmhkABX7E5BbIGBDhTbWghZx
A0R1+ciabmlAPlM55yBr1r4fHhrD236Fs9oZHQh4JzjX096Y1OPMV5IqFc5l
J8Mp07xH0XBJ565QG07ycH1oEth9uGnhHhgi4oW0r2fS7fvc4sjNA56rviuS
10EfGnoidJ+7QwKXnFImiMda6wVT9X6A5AO0jSjBEbMfqp4gyRhDPKUIIhvE
JLYnKAmynBAqrk1UPthts+MkJWGUCrxU4mM00wh6N7I11JIacjhoyJgVKFRs
l6oljHFhfOjcC3n97wJE30Q1PORSKR4ScSSZgW+NuNWK4MWWF3KxSEa1z53g
cZNtC4esZqh2TP+N3DBVA+CIwE6wGYDb3D+VUxnafgrD4qrvmm5waxyb4qgm
IJMHCw2KWmSapbdf90rzRSoN0vbj27zIaNf2RcYziO9h1Bb/OHjLZ5cE3XFE
TjlE1DbGLIf6fJHLC/PhqNAii30VUhXmmGw57BrTQ/WND5lLMTpjI6hLdGJi
oh5sKgv6Q9hKOleWTSN0IjS373R+9MJqtGTyvJq9ZmK9YnGLZOx+ENienO7J
/MDTU/Lexy/gFqdKf5k1vfVlai32LBtVT5KoMRuzgS9rp/CNXSnPT8AzHxhc
RR22x78RfmZ70RTGo+2mpcj6x1E6fE14CyAfdyA56iMl4jDkq4ZT/8byjVLr
c+eYoCCKE/JF2woMqlahv0VQwHHZpc/fQ6xrdcEEKEfZQs4nGParJ5L3b6As
oI6+10wywuTbNmUMObpe1PzAa5FAQnElui+cwnmpuzul/Pu+NRSS1lOLLuDu
evAw1lfbokEVk7ToMP1ycsr7f/pCJ08XoqXsVgeairs64C0RqR9iCIFdPiiC
D78sPFsxsah7azp2h4LKbUJA/b2MJvvryht8YAU7/g5sOjdOUH0+EdhWcsQW
hKdeoEyNZ7bkEYMAIxle2qj4wr2aKy5PpbysNqD7HAUCQw5SAixB75We0MXH
5DqWttNWP85vkGpbulehrnI6VB7DKPRCWqrsvbKLoyQAT1MWma6uopLK+MHm
ZEHfcN3ytPG0blLK3kcWBOlukf7nnIHWf3rdggLY0v32bMLSi1cXcJRkAWAb
MU7qrA6Ajw5SWdFwup5H2g1VVuPUdobfW4UBrmniqo6SFl1pALSR9YI8S/ar
T9/HvMDkN3DzB63X069jb+mN9+0HtjhOe5uH7IdimIbG2maJOXz3eaWOkir2
wPBd4TqioYz2dpWZm75E922BsHMpGpyDQLzK4LpSDun3s84zzyGbReaojUAO
L5/rX4hVngxGSkO225lpTqfRo65+glXJtuYQ4dQY7tZPnI48msgBnM0BvNcw
x8sp4c6AP7PJTpT9BARXfKtUWM4SXwL8PlasE6aidkOzOM9Z2ocdL6GSmD0u
3CkzA9lVej1+OGHpw0lJmzCgm92Me4jLDvh7iRi9klMWaDeR7VTTCazl7WYB
PTBsco/58a8+AtQMLAs0ca82jQGoj9wFFjqPe/O1quuQ4D/3WVAAu0YwchE7
LTRDnRpJuFsRXWAJzfBQ9+z8IRL2Nq/pZQJLipkKm3HgUasDQiyleLWulEqJ
snx1y4O666kIodCle5XvhTTkl+mdWXf9jO4SYLGV5Cas2EZhzrn9Hzya0KZy
yMiHKAx/9hN8tHi1SCgTtDYynQ6L6wlhZtZjKpKt/9ExkgPpfUE9DFo2C7xL
vJOe+kra+eapB52aJTjZ/5LPpnEw4LvHRY+6hDVqpARL/+YdzcqxSJLindW8
RET82o3Iv00Bt9DR9QzINkaE26KfEQpZg8q6eM8yXOyRzO+xjyOf68FTlxxW
QKFWfLNUwQBg7I9wavNMDMKdZ1nm0EaiC2TtuRefmHqaz7RLRo/c/tmj5XVN
okMPXRucJLeaAlMZURBaorkOa+kNOXQyKlit3bPO1W7X8iDf6rEquEoVbDNG
4WpbezVKCvwNkrZAnPKRA6TuWQEy1/O2odo2iQ2Jhd0uShXmdjxEVxfrybJe
29RDeF1D6/rzVxM0dLHW3XBXHrlpd5eI1f+Vi9uEM/dNv8+ktAeCEP8bPmVn
u6RSiOqEP63q+iWN1YUK547iH/WBd4LR07AfNX3xP/KT02AVB1bmFbF2d/jx
HPCppFRYdJV20MIEbB1i9ia+KfZfuAF36uojv65KW8k+agFbCxxPIRVFv1B5
WXpjeki+jwAazyO1hqB4nGH0gpfqvOqsJ81cs5UnHFDDIW1tz7ytuExqKpXs
mBYLTZJwaK+PVvsO+wZdbJx1uCjh02/vydqOLAH5T3F2tMK7PICKrVeKo84t
vyhvuMbs06ZFstMldIQtv4wuBpInJrzKz51CDJj1+xdroNOU/rKCEzQ3oiFS
zkJTKfC75QhDHIFajlAwEbrjAufoHyn0RXNXQLXQQvUnjCwEyf0oORY6Wku6
NsM+1GY9GdTCzsCf78MlwxYj9Uw6ApgREmVnYUK5yZYibcVg4MGCG5z1ucXJ
1pH1R1gIb2UQ6f/YUi4d6gsEmQtfWArZKFxZCG3IeEGOuRTbXyw1jVyu1Xgi
Clrq6tRlY6vNQrxzlt6uchpdmoE7sWMlbzZp1NIl2urv3OvcStTL9raqUSTl
HMAkkWZ5RIxRfd+yb3k3jVrClmN3MI+0VhiXWaZFDZuXxnTGFS2mF4zNg3d7
UPhDGspsZAaRMOKQTBKcZOVH7EVajeTE4alBl73GqxW0Db0fyxacYfbLs90J
z98R0oSOQTCCGXkwP9MCK+DijMYwL+ZE5uj6XwFJ9PGYrYZ3QLzZ0q0zpkzH
mWl+nZg5KNiTaM5tgOoQX4CJ3r8Nn90OjLkFKHGvRUhFr3z9iRSwA5tiRsRT
/2AJ5gecyZ6u/MHb5lcy7KKRozVwMLeIIIr8vKjok4olOg3dN1cetVTDeUJb
J61n4LfAoVp5fHVi9DMdIt0A3+r5X6U/xRFOltmVMxxXqChejIePBHAZRGfs
YLecdeDkS2MlbK2P5t42PF6F2Jv7ZLHlFPpyePAb9h15PxsDWFyW7lsbZqjb
PFJJ4fhn3k6BdRd4SsQx1VYwKwFOb4Np8qkSihHVAo1XXrf2SQHE+EB5bUT5
qx4XRnBszqRHVl8GBFTjhn7RH24jQu7omTnJ2DpRmsVa65CQ5G4t8OywtYbh
4rP51NyAEs0qAYXVOqrE9PcbvqU0hU2qCktEzm+QJoCboKEI3UZWki/9BAxF
i93bqgMkWFl3c1bedRAXIpIP5bRIp7tlCsn+3FNkOWIc9G0+OWFBzwfSNXVL
oMZLD3BWcLlta3TED23+J4IRCvsIxJvlvTLsGIYL0ESjzl31jbUPu/gzks5U
VZ7Fpi8L4I7u4Dkn8+cM9W3hQTM8mCyP21aiU/rET5M8717cZ/wA4nAvkxq9
yQ+z2JDiG7yzdbI0nC2ttDaPSUh/Tdr1mdHBQdFjGIHJt9VaEh5wIAjROH+J
GozdmzD3WNq+WwkasmVQbfdMq7XLiBiKOqTZrDLHHKXRrnFDzvIT/inl8a7m
cQ8D1mWadU120AzfElUcgNik1G38ht2uWeItLWKGMTmuwu0SxadeeAH21cMF
N+cnAi0BpmBEoIieMCxAdfHhhinFHe7DzLqb8EfZt4hmK2QLCQ0wF3/Lcwkl
9k+VbvNyB1T0PuZ0Vz92QxNnJ56qFDF9KcBul107yC2dPJpxxI9stb3vVaHN
qFulLwl0gVi79fedoTXxiOrpoEnBM7kSxxjAO10DitXT5uCQ6b7HP1zx2WET
0z6QTcbemYOldKtqMjyN5wLzaRWe8NrSbpuE7wsmpIoXSjGwxBcBsvS8JJq6
aNW2dpRPkD9LEAGvOIi83ksEWL0aJpOn/I6g6c6KlrZpJIpehI5ZfLsjyjXb
wBTJ0Wf7NwDH8SHrDxtK+vHRR/GhilZ5vqKhG4HVLLTWUTSMKLuE11kd0VmO
wI6G5verGDHmnOHz7k/nZdUSwFv01JELrl/lmb0bs8Y/gLVuaYhKNpbZqkzg
w1oOjvK4NwdiG2HS7z61ypYEWcOe14lqFmLFK0s2cY5QKEt56Twznge/IK6X
hvUUVo8lF4RxB0lh43zdNecoYhHSJ6iMg76dpOboUTsGTiwbYOhMpsyZPFgc
3YpoRrCuDjV8vn0ZhRre7Q6sQfWbs4kR7jwsCQ4egmplCDp1shJKCUxZCxZl
JTUOlrXYq0vPR4y6wU5vp6RbDm9AILl9bPSPN6Vm7TYXoUQpREzZ2SoB9TqX
VGPliEPkxj2AA79Wam9xGpNlg28P03QfNb9SXKjkCvfpUIcK3z1f+qT9M88Q
GisyBSth7W7d2t68y4d63vZvRxXjJF6nKvt8k2uQgl1LJcCuMTf+awHoFNcv
nZH7EYD58SrR1rgsHV/2/q7DdLkBovTxRl1mtL6LKdvHLb2bDlj7EEuVu3gh
28ELOpe/xhmlN6VtJD42rnHkYOtjCK5WPRqyBBnK46tu+eHc3uCbt4d8DZDe
667Se0ZMbr8vgtzDBnBKcvKRVNBAySRI+xVZx0WWYcHpk0Z3KpXt7kZRWpFK
1NGWhmRLsmMfgWNhtbOK0sAwG27g0IDW0lvMI11M7WfU5IIQiIhtaPGfxMrf
IxZCwfU2u8eZl5MhiaEq4yuYJUxI1XiGUeOXATDs/ab+d8vvYI+5OaB74Jmt
68HxTJKqoxtrxICQ4FITl5PSaglVx22ZkqDzpO6FYMYN+q1yU/0/gqtvVAR0
J95lnY8NS0VUvgv2534nbgfIQaVLEzc/ogh1BUVWz8gbcjOUrdszz58sKcV+
pCrbmuAsnfEY5SWDG4f7wmZUBpmey8uGN7WB0lLRVaFx4idl8i00hvfjPulu
SDjVi0p47qZD655ZspcRvopm5tzc1BpZCaBvdT7s/iTON3IwHMGmIJyZrfur
vVD+myVgQFcPws8lbbT4j6dD5Em3WbN0YnlGHgtG5B3fIAkvtfikQX0TLGbb
77sqhobaJNVaqlvSq3nKcPtQ3uPdPL9vU3gw10jHQV66FWZRfQaeAtqafo2B
4a3hNOf0gKibYOd5KYY/FPuAjzVephxvX6U9PYstPwbeN3m2+q7znF11ELhL
b/FOsM/H6r8QssqGHhSpz1kSsR6N3Z2qTcTclxBG1axp7sPTlkhfWAvKK7vW
3iwm9vatAbATCz5QV0oyZIYaXY9EjnBMazXOr6+f3XrYTYB2UnJMtBG9A1G8
nuaeFmSkBX/SEzSo19HYFoPIyQm6NugxmONiteeaIA+VxctIGfB+7NPcNk2b
PqKAKhEIUyVrvh/V6vhMIVGw5aookjzJXWNM3MdcxoHswqlFaaVkij5ptgri
Y7rURCpL4VlquuZNCQUTmOXsAn3IJI8g0kl0KdySytMGFs0fq7lEiNUWAVcC
95q8D5pDNrRvbJNLnzMSMZn9nh9i8UnJkXVbWWxQU284OkHw98Opo17k76MP
yYe/8CVOj02KG//b8eTUfsyeT5OnNqzX6uII6mk+yyQFDQ1M1VZ0d5XlTGeu
baN2wmHwVnDCuDWonWDF5aAaaa2+HchECK1M0L6YQrfYRRHXy8OK4l9Hk8A+
HAnKQR+gxn4/bwnGE0mvX4RkrcF5Top9XLTAbBC1RG+rWUjxOe2PeaVB0OKJ
jj/+xherWGrIX2YbZKKGnVt/ZTuDMI2oVpUBEafoZWNh3OgET68lqKmRwwNo
AaUgwrlEv63epyVtkFbzgo/SGerRLXiGm1cV7cWoT0nvhMy2Xnxp3F6o0qZo
IBSnq1qk1g+Hj9Yrf0IoJc9cvaft6XQkV7ysRdMZ30Tci3F8XKeQXaoMmyZv
JBUU7jTUzsZyHo72uNe31vEslKf3YJBB5lLveezRwwTWIe/mvQYDaP9fZaQX
PL+KHcl/vSQoklthDw5joqsGVVFW5I8bEkp36uU552E4bToZMEYzBSMv0SxD
RVHoT4LWclAdZZXfdBg8Ey1TP18PfukHf0rfNbd7qs4LvqRo7HaJTsqKQqPq
bInBWL5hl5SQ458vQtyaHiABrcsJ5HlGd6i2grtDn6vYqw7bGZzlNRkf1xm4
/jVqVq28ToH98h3AsMuntELP62BuPqvo7Q1M9XqVSPp/gAB0B6BGSI84hN0f
ZQLtCOKrGpENRxhob7XthGD/rff8eEZ81RZBsFKZ2Eh6DGOObMCPCPvyLhDd
8vkKVgsrSEVkykJOfc2nAsLmDyjFhNEaWYQ6MFuX7Me2ydreiKqdNitn/WEz
RgM9k6N2oxIUj+F5fdhyaOEvua0xJjIln8eatL/O6cw/169TbfRq2yxTHleI
oqD5OMr2Uv77dR4O/1TDHGKkfFrrpFdRbI4R9GKoVaRtH7/IYURn1QE8myI4
tCsrBSpWx4yi3LBpk1eNqW9SPgC2L73fQQJA4pO7kF89QRrZX1UBR1DcpjFX
KxXR2JOgYk+tJXFGDrvMZajJzjoPwfpVSszRtzt2lrJa2kLm+lsSgEm57b9y
oYLoY/z2WLnqsbyLvS0yhWVRb+4sqhmLHd+g5/Srk2NZlK/x/bj2DMLKKmJz
vNvywGJUDQXjStXTAJxbaucSjmUDgpUwUFUYW875Am0o5k0xNc8vCOSqCz2g
PkiAo2YQEV9/5DOggHxfuIh2lhY8ab7++44+YIJrmcTpn5G1yBxRHdE8NrPp
kotSp96t+fKtA7q9GrR72f46TOvGEuxSTmhplLVT8zxMs49IY22cAL7h5lUb
dqWz4jQxhbJgbrM2xR93bTNPP+M+x1SUvm6Iw8Yayua/viHJ+OSARAmJ894z
wjkYXCCeHPAu4VkXQZ9RiAryZgCDzTGHsSVvlMIsJ0WKO1U45f+5NA0qYBmq
+gXZyFerh0YfllLLAiPKdMmzaI2k2CJgECF9kOVCOVrwv635yBv2pIxqSibc
v23eW2tHeGzfq1JuxPabIXGmXknW+ZtExk/J0VtFuSWmWASXTRZ6ifmVeC7A
4Z/tX7J/+RhL7ewRYU/QzrHaFdB+EgNJBUNZ3XRLBVxz2pd4qjf54kvaTJ1Y
DSO3VjJv7hSpHHxAAgBgRDD5zp/qMD4kwqRL6nI3f8oMqRRxvENg2e6O6P/C
FmxTjgJCU+VW7NrQ4JUoxZ7J+dInwKXDtpUSSXcJ+NLOYBdC2Xmur3NNPNBA
JYpYFzXUPDbRR8786Q32Px2CeocZOxeCcgXkqBgoURr4ZEJsdXyqC6sMg+Q/
667etS0omPmY5n9IivUWYVt5rjNLYqQWwnUDG4U7ofDsPHmldWzAPF6Cy7WR
CeCqwXL1JsHacFX9xsqWVFZHuszeyN6dSAWoABTn9OTOQeBmkMWPEkUlS60h
tks3Bjo/wbw54W9xvSWFmwO9uC7ZgCxD0hY0aO0X8C7FuBuy/XAN4eSYD8/1
qKgfcBxQ8wSewAMlsSJraeMO+qhTX/x605BU4BCG8sfQbRhwmJ50vPWlqsvT
emFJlfVzXvxWXWKdhxWfWffdCHsL5N8vX+sy/1VVzGtwDSR7hw2Ff+bJnekz
0BJXCSFtPr30fdACnFTf0NIh72exa/Pl1J+pZxE5eZvaHHoLuc/LKPsv+goa
cPhLDGLnlr78vG1bUyHX2EdZTtLOV5fM7kpHKsyYMsvHGw9XOvn8i3xXCs8a
9NT7iuMm8Q6+B+x/G/MUM25HXsqSDAzN9xdOo+4BmPhxIyv9/IaE7In6wi8L
Un+TkUGeiHTzRiWhczeedV1/0eLBDwFmNLeWe01flh2ySR042VsFmj7u/oN1
OC75jHBAZYRQDnahflESlYPXUnK0me+641aatwGm7dP4Q16KmeSc/VbK/4Fd
5m0QH9wpTAgpFVJYoQlMsnaB1tA9zdj3orI04kaKvhkr7OcVGNoqvbSFLWTf
ouDDP+QR7SmG0YA3zLOe661qtsMbp2aHqSrET5yysYnoUdOoAdVxvzrt59G7
66rWVdae0rBpWu/NJOsIf9l+sK1lgA4jqjcDEuHcJKj9jf/CMQ3M4RzjdrJ0
8CGefP2keZAKz5T/RpqlTKKpMFZUpp/HA5wFRPVXHbvLeFWQrqgrLrS1v/WT
1NAh7TWvDIpbIAWHwGGIotFCmE88zirilZVg9kIqa/DyKJSTE48CwKIK/JYs
3yFaD2WTg73tP/J+oQLlQdP7LBlfu4oQ0f2iC274y5GCX1VILCzsKZh4UwWn
x8N3nNgR/DOhtrmmnGT5xM+FawJ5QYSOgRW/+t+erzDkhhl0YBVXOCQxUW1A
IuWdY01o5xb+/cufvijz+rK8lddihoFW0kebGA5VFaLtU0l0YRbaN93Dzc7V
uzrxZU/g0DYCnUSdBuj/g7tHiF862HWaqJVhZHBKT7XOvJ0QUdBcYLlI7FLV
6SKeG1Z+oKDw7EO2EWXGwzncLrKMHjUuJeacyc7ITvD+PnSqzjMHNV35KaNF
o9g5Iu+zDeZMu2M0duNnUnCbYroawieCOBbNcMwIRmWbVDtlbGPEvb7UiaC+
WdU7oqBOJH5ksZD1/5Uv5D3l+N9LlEKWmhyCgrPHCvz8dSxh5PK6h1ErFuE9
Pc83wJXryO9JHmV/Sp1rQcfIyz9AFv3knc4JNOdcE2eftJ4LxLisTKT7Huqf
3RBZ+XHlxxGSmX4GtnpbxN7TdH9P/shCxtJpTqeBADWcmi23jNraRoPcqmXk
BlGH+A4jHcR7Q2iK4/gysMpqVdU1yvSJFTMfW0UAaD8crOu8d1U3kyb12aWf
qr45MZRbfIXVRnMlBBDAr2qbjHBw/85dzmD43aRoqTKtJ/osxhLKJePjOiE0
3pYBMBievtKwTGwIqSG0EcQ1jGbcEu5rAkG4UlMEbKzHqrK5NmpRolmquZAn
fGXhnCx8LDpa1Mpk3rbDKU4IQYMwKWYWZ3XiLXeOndKicrwme8kaQmXXcnyP
qn1wGgd1pi63qQ7SVczyBi9FP10m53IkRFvYhs/n7d9HSJezDKkYCdt3KJ5Z
jrsHpTbIaAfxur1tfw9/PdsmzySh6OlKmCS0UgHmqh1C9flMeDl+UHsQlcLO
Bi67QMwGwPpIFNaAHBuZsSIQmMKOEOg70iPwkMXJ/Yx8Z6aqurFulaUxEmMq
3a96GvLJlXdzia00vgJy/Eo2r1dFcFqTE1p/prtHG5k3dLJR6H1NnB9Ej7HY
9Im25VY/NT6a08LmEowa4Dl3zk7V8qx7m+GwCMJwX9XJDnGcLA/O/ireF12z
J85sTrT9oNICtBzMOtDIKjRrIZxHz2BdXy+RYgzTcNQyNxwBM9JQiwCfLqwb
RHNEfgG21K6fcYeLhEAvkffCSjIU3KA+h++GJsu6fXE9X17FrvKPQzb+T5yt
nQX5fWwu2hHIquUpcMq3rGZbRVeHkvp9aKjbLQgVAOlEhRp3f3TUlb+ZLBGD
yMFTXOH8dbipdUwThVTKxIJD4MecUos5CCJBjY005pzo1hLiKxh91FR+GJJ4
HWyfK4DATVS1WSoEghudje1qsqKi//zLfl3gkDeQa0WlTOdOMJqp0+w/jTMM
OQiJFQPhftJ87us4LBk+U0XFv8onmwnTad+XI3r5G8v3UQ5iOa9H3G7ZYVRU
pkFBgP60e2IG7M4a5x4gotThe+fv7RDb9M1iaIcuP3CNghvD9qPIfW0lbuHX
BSzE88WuGUJbzEzsSJOrQaDtRPbKlvcAfAG8S2Ylt880aMTko7WdcKBvEiKV
UceVMATicgNWpZRAehLyeZze3cNblluvCkKEKHmUhdFpxuph4KEsF3/UQOQJ
4P8omgRLRcHF/pV91R/DBJ69vfNxoYQmwIq3Vk/YCiedDD7tNyjn2/h8Pr3P
wUG0sM6aN9jbY1C/MUgljp7UnYBQ1UwZLvNIYiIxnOBIGYs7u+4le4+b0k1d
A8mSd9RFDIB5Y+egl8JIrcMVmZW2waMpKMKdVdMjZ2AHoEl1oooDQZ/h8Po+
5z45Arne2OwR5NRZ3SLkt15bMKuP8Ykx9ToyrhiOlCyK9xGK1v9VZudooTWV
nvsogFfvx6ESeCPxmJWbV4W4JfSbfb0JprpCiKgEle59yog+JXDmRuORguJ2
ZAQCATraDxIwoXSA+6M9UDfGDggdoIelR2+xx3CBiig3w+oEV1K0tw2VCTge
8ACIL7kGyEcEmjjMBfj1HU+rsLPvffunmEVgSwUKGHN7M592HNKgBNCnZHM/
EhYNjcmjYyIyAmfZce1IZu5GNSkb3qUXGMBS3Fomtw6QWQn/h1ESLF5A5i7h
+llFW/lrKX52sZd1qCT/sMpTY7F/nIOU5eUQFFs3JZdhkPBWrgVvyfkjOf8D
XQylU7JY+Qu2s5Z2aDD3X9aBNeZ5XjlUGAOyv4TMChXvgQk+TY+ikUJMFhV1
OPsP7r9+vH9/1VkyAnXJEhBDnTlOuVcN2VGJmNfoBe5YCfB2ZaHcHPeFt8TJ
Zx2q34Q4hy44TM8Mbj3oEWablgKWMx6gSenTXEu0rZ9CDFMQoz99kVW6Nat3
xDsq6ymTNhuqJkXFzElKhvaVuIbP9UDd2Owffdhiq2qQqJJBmON1u/CDmOjy
BvmCqvt4uaBLIZ80yPRsYCyvDZD3IfdveLTfxjR9gXNrUuIcrQn4BLOyB0cE
3zYFhwGyJuq/kt9BAZ/1f00LwkOgtVwPJZHpOpEzRDG/uI9pwcEzH1IXH79T
KG4r2LxmvaYeEDPfoyIVV7Yex+PYfl4dlxgwb/jB/i22eoRyh7G0NliCBROK
qdc3oli4swkvmAtsq2ftZ+QmMyZISc7oGbHYvWgryPEvFqDOVKCpc2QF1XL8
ykFqhBbEkT6H7erQco6USbxWv7tEdrHl/EKKmceLfmShJgK4habqqEkJ+Nyn
JI9lTdWnQr+KUITs3qKehGbLTdHrOOriPMPwsIgoOpEUACEiFctyKOHfXT7f
de8pQUbI2I45SjrKAuoQrXgdhqicx8sOSZnZczzeG7U1/3NFPbtrZ2/7+BS3
/SVdKY3CCxe9iSdS1ZnCIjIQCl0p26hINi+9xqZHfKWdbXFCWyT+OlV3HhBH
aCbx8lwS4gfuKCToUoxsV71zsyEhrv6SgEpn74y5eJg5b3pRlaK7u08E4pUU
k3OsohQSLHkeWYOWJKNJaX0cx4jFGKaLp2ZM17Q9CaIsLYP+5qe9k5AkCLwp
qXANkHn3qCb25fA3JL1NT4hIo/myOIEt1hWD/2vauNPaWx6ocNTJwNPqS0yv
lk8DlASW8Ubwa3WrriPeW0/pm/Sw3lRb6zyhBhbEhvY3ZV5tMeZEM/Eq3jDd
Jj7o1/i125PEeSLFdnGRluLhDsJYEGZt2WJLaGEgq07g66Ri1iwfRqk/oo9x
prg/OKJNtAPwLO9mLp7qrXP3+VyuI9EgEty3xrcsniwkG/mx+cKA86cjfYk/
02olUTXLnueTbzG7Z2p05tOWHKx6owIP4abq7dxc84WNzGymOZsfOBJPeHPD
8QX2Zf9GiMzpSMbrPvjiWYEzhlXspJM6x96DRB8OCYMIvfbzBQt+tRkUTy7a
UmXDWXckth0aPWgSXWY8aA5vvT3W3NzyJLPfSumHJwxCgIwhPo2EoDaZAxFX
UEv3sXjoLttxhZNZN+ub1MFNgHfBx6eGbr1mSbtLo7CzVqLVWGQ3PxmZgO3A
CVtz5yuhpgJ5n2g6kRX6eJuYaIcINqFKJrf/w+jyQxpdEYRLjP0qQsby4GJr
7v7pBO/XgEX7a+Vp2WC5uBkj245JwrdqL/IiEhjPPl+j1dbyF7/oMpx5nHX7
aUeqOJ63d5Q+IKgMBmiGPHSzlJUeI3+Px10b8qIVjjBojeMQ0C5/8YaYmZpG
LffQ1QKwXZjoKeApF5k4fOYh2vPiiWn7xx7mQ0LUIXskAWoDK/Rp81d4gI3V
3DP5acldWwjpgZuSXDI11tlCdcu+Yop9Q5ngLcTtgVEjGDGOlyDaOIlBpaj3
JidKA/P1OTmIWrT6o286tfabUFF8H7+1mIWIERcGJpzKQHV5s7iLshhpy0CC
IVnKC14CV79tLGIWMNij84FA+YKrSNMVKfOyZG6fir4lQJypH5iF0FH4cghy
NyXeawLTn00F1wpVNK9bA2rReDVAzaZBPUraQoHWaOhgHZLVfgzY8XaiCkR8
VXOgetF+AxQdftExw2/X7EhbElSypD36Zk5XE3ebtBoMQtQYwmAn9OqFHH3h
mP6vRg7mPUrATv7qfRpczw1gh/SvRt+GuCdGW+YWkXeJBobK6MuF4vSy0rbE
Jhu2vfpWezlEi+XH97nEpZJFx3LZNmZKBNPxX9qIksaqzJdCPTBMbHdgstYW
9F7p1Y8N+pngMzT61Xmn3x5utChsV9hkwBon9BbQHXVQ2/x7a3S3Cwy3JJMa
w3n3weWTwZR5LYfAcFMeFDfstIVc0vvDrgX4QjK1MDaqEiWh00U9gxB7xVTX
PEId8MMRapiVWA/PAWPAtsOS7HupSOYd0cKPF0Fdqj+K4kfbupIvBc8h+3g3
eJ4c4M3yXACtBwvmsxzKR/wra1W98dJMDRvo3xC5HtbVRyRy5umUorCarkog
BjE2ZS/RfLcl8AWfHq0vuycCUtxMKC2NRyLQqbP7WoI2d2oPvyhZ7HTG9cWC
zce0lw+CTCRXgy0Yrd82+mYEk294YVWtF1z/+m/IT+vm6w9ymJ/6edjFVndY
CN56mPbrz20F14/zgERIrb6HeEwpi/sBBouzwtvoDbIVo1rvG4fntxc7ylRf
siUN4x1oDljWGuGm4w5WhobEbk+m0oCGyCbzlb7Swf+4ww64U/eYcdyrYjlC
3mpugCyjdwU4Zo/sI2M9rh4pr0eY5BwhNjm/htXz3U06Nd/9OYEpEI9snyRg
XCyZ9Y3vlIpEU572RR4PdIxWR3aGLfv7IZI35e1oPGn0EE3h0gS3885Je4GC
edZm2kl/kKNTswMHGG1PCKF9BkTjWzI76dse1i+LaeWlBGL4Bl7W+kBSxn/y
4esJR0RovIET/XCC3k24Xk+7B7yM0AZousyRO4uPGtH0ZMsnAdQajiBv/c1y
ZjXH8GPE54N3jFjAvEIC+9YsdgaNTC9UwFj1wEFzl2e74p0diB5wTltosU2l
5E/B/l2DKejBoRA/joV4EmridPiTPgUSGkt4YTYptzgZJ9VO6fZpUF+dALh+
oimeBQFmKPxYRGxIvVasypZicZqFwJ4odiFkPL4YedKaj26eQnAeEbRDgYXg
RFimzawbTgPB4WHmayWHuUiTR5K8hSsdkmDG8ArMrOBfgz6PmfRcOjwiVUQt
e41BOe3OBW1czl21W75P4ap9HmktGqg3x4rLvgBLV6+3qtPhqUOlfjxyUf7e
Vp4tGx0fL2vVc4trGJgf++oaBdB6GwfV+FKnmWbl8iAVHKECKQJ+aJRl3GzH
M3EdoxiF37k/w4pz4fDTuJsQwtQ3cBwM2sETM2HSqHXSw3rifRm0fMa7JeZs
3hE/E45O2uzciL8+UkpIUzdps2n/P9NtcBNV55Adzg8gMhRYV84iXzNlsW+j
r26peRnNm/JUVcVPJgO+UHXm81VOnMBFQBhDzQm3kuSD7/S68rcN7MlagJOr
dbadMDMA3KqjHK0JOIxn0N9ho8QOx88c0J5q6i2WTmqkE6kmW9P5rHYxE51E
8exuHC8W4Ete8x1iWup+eb52PIqk6Jzn1FSLGz4oaj6iV5Jp0EsQufhVb5xR
OPXXW08Zs3YsGPmKJgGZoaChVj/KJGRGf2dPJDiHiMaEfKmU0EaB7ldCoJUV
tN35miMaq5Gg7+CgQ6xL6kYj91hIulvv+65kLsDstS6+WZvA/b94whG4f8GW
87Do7DmBteD+B41RuZAjnIjSiCC347EUXlgjxOhNi2FcSG2lsDepwELpxiln
hGxjCy428fdaNZWpCFVzkKU16DgRqxn4b1fGiqh4SND9UgeuUYHKLQUztuMi
VehfSCVwZnjpCLsJe++fmkn/n4eFV4hpPJ5rny83C+bRQAtEHR2kqrNeebsH
oTK92KyOlj3q2iMRWru7pdBqE8qDmafr4seYw8nXQRjH24M7R1cPUApb432P
j6Rs50/l3r6BnBEHR4wT6jR61TbLsHovY11PQyTa4gAFwwDdV96Y78HFlPpK
E6L/dSZmD9Zk2JZ0AVcRdS9JFLpYnY+iXgBbxtMIgLdgbxQNky1idQ83Wrm2
BZyshtf6p4x5I1545wn2bGWlGiXPvCO7R8aiDzKtgVuO16FCoHpVCM13I0sQ
UpUU9VinWXOiMxhRVztZfPLSLWybkbxZvNxROm6dkszRtQNiWiJUyUfqhrCP
NTbpzq4nF63EooRhRUJDGDH1leeCoyt9WUgGdOP7NPyKaBCdGxJ2DaxDCVGK
gIE7cNjKQhLSODhrXK6nQpmDCPtfv1+RGvYVHAtkpgZJj93CAKRdhoOSFZGn
dO4CT2jpbE4M+XCQlHghheMOjA+DqaoZWX37rzCmW0sD/O60RwZHCMjze57W
Qg9KlZ62K6LmOedoALlMlSa/46rps+K3rT3B3aZgvRCXdDINux6/IWcrQKie
Jd4ylRH22Tcj9/0Gu/UYQsrmhfWzZX+ZAz3bDPTuY7dA4f1zLBpToKKOOQYW
oAP7Otiu4fl7Obm4mFQoRajfdk2cPBWJ/Ash3LYzeZYZLmQ0IzGFpAGSUFcT
WhCqvDCLjjUnyymxJxo7qa3SiDoQC1+vgG8ks4eD5DOKYVAEaOrGYQe7tEWZ
jdMIek5+8YEOr7pmGQ2P4XH8hQMbLMnIhyGgTLd2A5IM/NaT/tS/+6/QO5m+
b6OLGmX8rGHTcAxEdmocNC2qsEKqQU0Gn/0iHoa9L2yMbpAP3fDFG6bE53zU
Ph5qFF3nNgZiX+o+cHSp8cUblnJBzTH+t5+DcS/4S0oeN0bca0MMm2DmdDrD
qek3gv8pZOMAWXQhwwcWt8eKQ/4J9iSo8G756w6WySGGNM3VdrgKjwriiaL5
PxP1/4a6G/E7UGvpJF96+LTM2d2c7LJszTDQlXX0pJAleBLVdPY0yQ6bTgun
InS84TAWs5ndj4nsz1YxVGu/U1rNQYTI8cehU5lSWj+xao1fRymRJFphSjZF
Wwq57JoAgxGf2iBP8Gv83/7276b0BVgFW9Rk/qF/HwPlAyPeF4bxKm5aSoTa
eFXjaH9siDBTkmYARbkjtTrYHYsUgo/18/28xZMEyPwFExNLsPkBSftePtUX
wKPEhlMz7czGJv92E1L34ogV5P/DAD4SgZLvyYxDovdtbhM66GL03+SFwvbz
LBCtbiAmXFP5yzKP2ccFOLA8jigNJUPlSU4QtqzPii6VQPFBaouENGIQs5XC
M2+UcBMxaEP2h/kJ8voddDRTSBDMRB/mhsk3l3vxhWyouJqKKs5mLglWhv26
XlQCt3p21TZD3K4dJJtcbjnQ4yUOnHmlfUq6ICqKosevtHFO4IC28xFUH1mE
HI/2x7/vHrKl1shK2wXn9A8MdRKpYBL6r37ierjUW0xd+F4Hn16FYrg2PO+/
V7RuC8sEb9m9Fq9howkaRy8YO9ndFlk6qikyHElsc0ttMqarnFnx/2j1xYsc
lDIokk2Z0IF4iE7Z/8E/ush9WrXXQNDWHP1ZvbXhvSAf53VwlwsAfqG9DZrE
1ohsbwSa3KGl2jNeYA0eeuNnbyrnjenAipqWSwPr2HR7lA6T0YWhQvh4yot5
IQ1Ot2JlQ0N+F/07WJyVo4lMr5vaW/SGCSfeFEdGNU8lr/gr7PJhqC7TCSGs
C7ymS0hD+o7QdBU6ZzyjMnKoOkVTULTM787Y52xe9yGKCOSUTd1Utyx+COBd
TdDkcwaM1j9A034saKb0j1RlinmU448d0JTjuHeC1GRIx1oPSlxJgVwP7lSe
lmqqwk0mhWVAlkpAP7TE8E6S6XoOrNXoVZzcCD8GTrtzEdBDJDZ1GQE0cJz3
7RLYrpEAFExuvoozx2houV3ORk2kZqsQIZE1DmdUqFrrP5xL0qIeHIJJc2Z+
zd+KiPb5YzHbp7t6OpYOA2KHBbbclebONSgb25117KZNMnEearPng+FgyQF1
EweMzpTT40oUjYF6NziY+X72FR1QGI/rSyZvOkcwzztUbIJ2K1Rf9pivY3Fy
Sk+fBbOlmAP06khTmhnEQdGEaa1b2kQJaSk9M1jZWlxkfIxGSYOg3oBNo9Eh
Wx5hGGreDfdneRMqe2Dm4T+Qz+IWcB0tUl0ue1JZ87+GkqpigfkqGdnyt98D
IcTj62RTloDRY0XVq34OV4ibKI8fR843BsMKVDfrhgpRED5mGyOKwkdFNl6Z
ib7P++OlJRHPfHsk/a2/GQFQMJa9zfD6pJbNEdAD++AZGQM7pYQGl5yLFL+b
LqX0NdMAoLkwWGvpDB1d60QR7syt9v18Vl8swNHNEyLzD4eCVgbsXLaDJ/T1
AaFXnJokMdhS6Rj2F6s1wX5AM28ZFCN4CLZ45fPKZuztXNzj+VdFjn9vQcNj
27jQa8xkZ1epP1vu8tiZS5KZ9S2xE4rInGAb53G/sncqe2MYtjT+/iGAXVPs
L4NGJ/kbZ1Dd/ouvRnetkdJgOivqTiHFLcwLEGNcxP422+A4nSbhoEAQtzUV
ZufoRn3u87OcrHW2SflM0QE6SvKvCdAObghd+gImDmWk1m6dxOdH6daOehns
gDpJN/Lj+A7iQGd7uTxG8r/QTuw/wZdzISbFjUo7xsCQ6e8gbw11N4esqYJq
PhExCOly80Wbznonrwu15kjmM6f/6gHF8zS6YEmeW5KtAr2ZeSw/wdQuMAvq
MatPt9b7UUUhJF94dlvWFsQoNxeWrJoiHoT2HL82tggE3NX/v+HskBzQrT6j
qtXFz9+7NzzaRMTFdCFlo2vQVxnc8F0BSfHcMWfA1OE1r4OCtlQy5fee4HUd
pRHS5eSkHztkaj6ZvNO0Y7AUiS+OMTg61REF6gkxanlZM3v/PhOgllcdciVB
tF7Lep+HkTxrtyEzMU9pg9BNz9QxOE02OXbZRMjUEKno7BfO6bjQ/kP2rk8q
m+HKIluemyHQP+8hvdx+Lf/D6GR3c1fEL2k/0ZdDMZG7C3iztXX156er9/up
O/rNSogiYi/S2dawQMoIjtovIzgeVkXtz8qUD0/wzdGf/lAA06Wweq5wE0Wg
H4z+ekvGd13B+ZqPBJci0nRNG+UvtmNtSa8MELYtOAdxZ5f6214uxYXoOk0C
afdyqnTLMAHYD8XU7LZOUlRVz2UStS5XHo2FJuoiWyoFQ/9yMXF/3Vd2OT8U
sJDpQ5Lw66ASjnYn7OrHdS4y7jMuANypwPdV9JgpmlajwgokzcYqaOboE0y/
Ro9vOXZvnZ5T52tfJB3AIdP82qdY7AWvds/D10IfliWP9DmHXXLeBB02JPxO
obzbjS4cPdFvNzU0Wv7Bkzj3M9JeQKpMdiYD8dvL1Zl1ysn+o62bMhgh8HwD
hu1VfWsZyuSjMZnGmtYO62IhgITqyFYAW1jxLv0crAp0P4fhJLAAeZgNMYQU
rdRhvAxmosK8QoBPMy4Y2+hkm9gdKfMgF/uOMTXxa/D82A25MUAkPyLHTtMn
YfqIXXyOTiwyl9Tw/3njgzVdK45egHZCnCp3V4wpgXfz2wB2eQTDo5UJEUfB
e1/WS227vSf3NlwVkgkdhS6a3NaGSBao89vJF4JXzqDs7+F4k8xtA6sQBaBW
XQX8/qLV8+6JON22Z6PLDpoMoqEPSrsHQYIcMj2gm+7XErRWkwXZtAOY0gpz
2zoKU5q+b01ZpizJ85VaWALUScTBNzCtRgPXO0Rm3M8qZN2he2rzwamIiAGG
MIAWXUXZVx6MaQmfkyR6c+OQIj4II58PjBQ6U3mFTaaJJJfx8BlkGeTnKFVY
+CxluiEnvVKyHpACarBelcIcggghOo/YUPhHbxdQZIBR0xsARJiuup+UGozX
l68R/HYnQRBcHNkqS3i6Lvux6oAM6u0fL/2UbbDyZFziTWHuQYp453bavugS
0fI7SbbP1cdhiBs78X0NmXxWrNSt+s77A6PNlXrZ+vKSgm7WGdW7PdP9ooz2
8SSRJGmBktg6mGKZQUW5Q4wrcA2K/WCtYdzCmaSDYwG4Z+zS+ZfYMZGg5c5D
bH4Szm+TWidArPgW17gU/ot4n67+SjGO0IYykhwpVWMgdxIf/eX1+jej7sn8
ZqXHDSXf1uLow3uxiMyqBhKIVyyoc+nuvmIhWTm1XrDn9vIles90Cs1BLFsh
Ccx/V4SVeag/h6EpSvM0gQQSl+lhQqlpVWB+b6mqME3VXmellMs4sxnrDEfX
O0VB9vt/8/OqiPTowtSWZEErB6KTgF6a4EtPq1KxzUSINbkC4UjzP1UOsIG1
aZXTB54M9a/ouTIlHI8wjc9za/zZDUsgyvsMHg8X/06aZhBdiOFNBLELQsxa
NRIXoWGzqYOuo/rldMBqV2l2j0NitHs6Ojg2CZsCh+r6FgOvvo3DRujxBHT2
U9E5/+keANHfXHXFbwAiXFFpod/yEkJCzf/CiSJlpuAPAyiLl2x36hxPpjet
BdJAtI/uKwBXgAvBFXu40poBFh1LbVrALHP7YTaUOZfOo0c2x/Qd/pJX5z4J
YFcE9o3eMjaXdC2Tv8wDp0QviD3Y6nNWsMKr874+GFC07XZJ59H1TotTMkDs
gUU3B8/2aKaRHqCrCQ6InF4GgI6bLe3ufLhFnNq4A3ShZzHIbvfZ9Hy+assP
xWmpdoIV6qfNmAN1xhPV/YtZ9K54uzZwHHISfdqs4pk//Q6kEOBN80vQSYrl
tQPQOvlcL5zMoJWfSyhpJA0/PBZPTH4XXfxBljkAOtcAznQ613da8LosYXXi
TZWDXB6fB6qK32DvNWuNqOHByoLiXa1ll69TJ/wiv/zZL7IwkU2qLez+IebO
95MUEubvcZOK4AaVW0gDYe27Z9Qy57FcXNtNl2kV3wyeJBZPQ2dBBa8lrYcc
Yn/61Im7Tjo32jFYCLe4fja776gl211xsTKTkkjxDE+Dns5TaBaDhYWPJfP2
ELyzShyjzkfSMZCIBVfgCPW7aqXRknVdN4oELoRWrepoN6t1gjT3o8Q+hFZI
g2eSd+76SbbVti06LFvLZP7yImk33ekRcK8lRRNexYAevgvZJnPeIHvv8VO9
F5BF++i6gizhgEMiMNAoS9niDp4BU7GT4BSE5leX7+Im3qtk6hzeTHNsDIHq
b4yMpGKOxqS6DyJq7LBJ3DzAdVSMCBpmNLWWbEGOkGlBr9duz0C4QRIZD/Nq
Xf7idsFzD/XtOPYyck3PBnNignhBNK56ie6EYou+6QK5PphcXqEcPVquNvBd
dYTa8G2q74sP9T6pbiPr/pUeSNDUTLqrWCu3qv+lIWk4uJbmEgNDXdK20OzY
yWpH4w5qFLcbkTlM9AsLtoi+sqQecNQnjTalDr9Zyt8l9HMzLdIp5nKjmqq3
sN7ec/7hrDpN6fMyUJ3qQVq/jqoAabmC2iN1wCp1sKXmpkkMZ3APLmWeN5cX
Kgcx9QOlYmrY4qDBv0GFIRrzl19acvmq0uPd682B4Clwg1AY633X9OBnllIN
QoUHsVbW4qWlnqjc5j2gP6EjWQH1e8iYJeFy8oaEJe1/Agko6dfwQ1SlVkgm
+zqKEbAcmwOK8q7wS0e48DPbYC5JyfvyWL2oJPmdr/0d1um3nQuoBk3dbjrL
RWR2hi/3svxbvoU/hDz+pZ0BEEtRSLyxJxE8ouKZf9syQHIgJrYvdohkWDs5
MglmrbqdQ4cm7FW8WsPQgcqKtBiqBh+SAJDSL76LoZYWl76QZ4s6mZG8As/8
jZtYwzp6TlOG4RiOJVcH4y1SvZ2YLNkXCjcNuT1NlW1xP1lxxUcNcX8JHEss
BVraHKIOX5y0WSgHOQtMe4XJgnV2Bp5i5o4kVQiAdBYIZHidLZ+so63CRFhj
ZguH+Xryu+rqSbA4uAZkiZIHfZBb7QblnH4W5Il65u7jWolE9uKG/6GXRDlT
8fZ3zSCc77tEzEu8rlkjMSTkn64dkLvlVxk3FHP1ew3NHDem7Rq11CMlJKo1
pA5aSoxKLddSj+kaginsxy0qpZpsXMijYok2yt71rzKOnDqTTrkGHyPZCu6E
AdNmMlZ2WLMqs0LwgDQG/cUi4ioNqlACOH9c860GNjPe2wECQTkTA5Hnus/Y
nBGsBxL4fcoPIuIGZx7SG0/xAN0Koj23HSzJDQ2xgFnqRzcs3Y1GzJZWPE2v
s7g5SWq5ITZBHH/OTAd1/44DZ8ecFF6JVI9r+f0PyS4bdEEMqzMw6K2iTijy
9xgATQtHg3MgJfNwc0TMhXUyjDb9CaKWCwfb5+Ca2BAPybtVTzvoCiGISjwe
OjXVFO7U0MkLtX8kEeDu1U7ugFhT5xP0+0Bgy9nDqTwAMGDYjaA5v7mDLSVm
XQS3wuvhkA0drhC0dQCW/SO0mPg1kGcccGOIJikOupZy5RSvUMs3JNB4FUmp
aS+Reh9ygA1sYeIyWq+Jg+XRF2y1wgM5wP6JZkHijQEZRJ1enpJIBijlVBcu
jFieZFu1JwWUxVxL7ptTu28t+p57LI0gfu6K0kHRNjbMbU+QS+c+GsZtcY1N
hhH7aQLq9uSqnSfaNH9XjjhdCluHVXmmbxiC6qRVThFf6R7Sf6h/vgIGGFaP
uNnqSp9AZm2FiXw5+XUsNdnt2iiIevzJLasHaw832U/w0u9s82KFuUHtJLbx
3SqgFhr/b57zokCD/hCvLZaF90MnogyUSi+mPJ0ReiyMr0DG0DZzY1xeUf0y
R6W05Lko629ugNDGZejOk4DNK4WvZjtzz4l8EHfB1/UxIYHBJJ2jkAObs+/c
DsHzq4iU7C4SyegNOVhPWxdbcUKnm3cvAII0cIl/njMF6YKh7+/MntC51wuA
UWdVQ8FdxJ3e7WwE7fg2f5eteUCQ7ZSAlVy3H67CUShUI6QN7PcpJb02wKdM
EYXSmf4wltjAvTEdYDp1fMEhb6hNYDZ+nkojb2Nk545ZuaCxPjhKGkBVRsEI
XA3wRjOedMpPiG4pb+hLHlM5Tp0JUl2VQ7QQ/gz4/WELFba9/qbGEpYjzy0M
6qdcL9hncN2lDhHYXe+cmZPnTJPZUPz2u0FH0Yn+YAbTFtdL6j5V5VxFSDa6
IGTKXenL7dC6/1G//p8SMTZA44gP4HaWdL82M7IXyDL/F+mZo+6aLmGli2bR
ccxefc2u0QSUWsXbCm7+1lFJdT9B9V7jogVZSkmhU3QmJAzxF3BswYLlSlnL
NEdnRDUeeddaHAehLwFeWRkFs257EXX7k5iE5euLlNaLJwChs2gt9La7mKJj
uxMrlpAcNeeaSli35Z0XE+oShsOt975kZPnemIhhao2WDcTll4MW/Ts5ZRo9
wKH4Ck2IJjakV1ZC1LvxrGvmT/9l9k8gf00OEvPY07ms22KoP8ACPTRiMck6
PaoTqkl83ALkzbQHXn60KrRnxo0wXCt8imkaXO24YxEkVGlHhzS9ognRS7sk
5jrWlgwc/K8yQ1g8gfQQnn0yahhmq8NUywwJuGeFuyAkJPJ1BQLJcmeECmLQ
fp/KoObiMJaBfeGMGMM91PBSuRiOjPua4FtdcT4ss9jKSr8skY0whi0+0Bmp
HyhOvfMlpu2opWpnY2v0fjYmcNOPyBQfWTiLjDvJ9yPvCu8Rv9/NRT0fHqjy
W85+NDuvzGR7fk2tu8iwPMTwczEudno/KFWn30XPMe0anjkNRocL7hWYFBOz
bknWOmMsHtmsSLSx3ENFeDUambvdr4LRuNIBK7sfzJ4//iR1Kbzy9VoV3r6y
I2eW6ePaiPscgzVLF79kp7Z1jjzKTjanzGUmZ03yIxV2fntFW8zhQwVUvQP6
BGhTJwRpWLWiduApDbfdl2t8QdZk7WgO5APo+nuC+4cknp6oLF+aqjfdjU+c
WOXXXxNSV4QwZo+PLpN17kE4wG7J4cOzRQ7/eRbmt3q2FahAcpl5XP0UwVnq
Z8/tnx/Y/q2aQCZvhI9UYCJd2oBtgrp9keXZWB5P/drAhGsynhJAdUrPc8SQ
1950xcLE9okKIRkkhZb8cyAO//u26ZfBumAiCe7lb4R9y2s6Att5wYZjDV27
I6inHe1vriLpWYoGrcIkSbKjCkivr7sU+dzHVurO4IN9vbADeMqUT6YxW0RE
sc2kZuBzC9VXQEjafQBnlabq6RNqacoc170ElVjJDvM2SuhoYWAnc2UTtcZT
159JL+1QjmVocOunQ41ztTxjmc+ix5IUl/BY+Pp/tpDpUMtnrtvDD4q8HLA1
jFSHo/O9LpRAo+g+IhyEmEehpLV74FnRGoQeD04oxHqqecHE5JFweAnK//8D
aY42IkOb3f8RkTzcdfDf6YRLuZmlcJjFoUIRr48VPVSSJnr3WS4LPizNwNJd
lz1YI5q+OtGB4ZxKyUTW6T8Xv9F/v9qu+BJkvjbacY0DhNtGMwv7fOaqio3P
ZekmhdI9M52d2KYax38StN2si47wwZVPtBXe2nBznM3zRh7zpdH/4fFeKaiN
7R47YeEYi0MZkFNzryQIV5WfoNMIKO65N+jGrN+7P2/Q1Son2tgBpVyxCtpc
6+MbvzNEBcjMD30dy+F5CLs8V8vJXJGxH+0edUGYlbDCUW/DWXOhjviACAQd
t5Dw6QJ5jMeEcsH0IajoR7+5xHZJbDeLqwS5keu8dV+PIGfwzw7JfeuALmcc
wiB8XW5EJeaSvPXEjZEXorqFnl6KKLL2gPb4p3huHNn/zBZT5XoPFxJJ3ehI
kpkkyQ/4FIutV4cJ2LXXoBPMndHAO2ej8BCWLdgb4gNGplnZzBvtXZcxm6PB
hLyeZMVle9uIslY9nZtWogLafc5fQHpgQ3euW0VtSP7xk+ymKN65VG6lFaQf
IG7oNFFLdm726aBJRevpt7x1ggViyeSkz9n7VyxZQHVRKyEzN5Z1uYI3EVj9
rXr+DHwbcKRX2dcjzhyyAzauimzYCIboX7895ghP8HC4ArgS/K6RLUHxK1Zo
HOFSAt7hXc9QU73pMZ7lk3ZJUju++qHx7AoJqeWQwTfh2kgzqPZ7V1Hx0v7k
eGlK4HuX0WmU1E03jKAMMaIpAYyGRDeTt3fE0ZM34POTEN5SN9hPTGQZpD9x
6c1fAGMrVfM6kFfal0wdGA19puAzK9eGChN7iC2nb8fdKsuQblFUwO6GNoO0
bBhBeh0B2Sj0BXJfy4spn45QXD/MGvt8kSEkCTiTP70ZtAwAYvc6m+rLLikV
DzCF6vdfM8EW+EF3Gc/DW6SVf/+jJboL39SP0iq6ypZPnYd9j1dUHdaYFo/C
NRdmMxwbE0TYYwSkfi1BqXE765JFPhTpSAGHgLyUACPi0Y0oollSbmPc2P2P
S15xFuwTAouJ92RePlClTAsBPWSYSMl3+8NGhJ7+0Oz87EJgGG2juhxr8h0f
GjGDFr0kNBuKNeLJHFuip7EcdtH8sv6QPkxzMMEgJ5lUMZJy+E1C0RFCrlQa
jaxY+glZB2VuWZm2+1ut1x6Y8G64LnnFDbnVNhO9+F88JIEmO/881+FD0PK2
rZJW7RyMgl3L3Niekql7uYDYi2ZbY5lPXgeRxbIUbqZl1zoxZ7ENtbiKpU8q
2NY9dLJyD2fP+efnQTtYehA3DPIQvDrfc0i/FYweSSHneuckqp/9l39Dat9m
+i9DC1OeQSII+0qSmpEcQZ68hucp3YzzzAf91m4ou7YAHLoRtpm2PrEC1m2y
EO5njB8ER2AelJ5C6NN3a1ToYpIFV1ZkSAmr522/Gx4yvRVTy8k0PDtb07is
mtlOgfjB91qnhlpWfdxlYY2bshVWdoamuHB7neqWoRKFDL8RVkbIkL3t9DNq
iApcBDv6acvJbSY/NNddAoTjrlzEqWAxDEggm8cSGmc0QKf3m1xhecPTzRJz
Bevwj/0Fx3+jG6PPU+lh7fWisfpPu84bJH86c2j4b7vsUfL+7ZuCX4tbAQ3v
Z8tGRmfST/8g1sR6tWa/sdoSg4xQkO3Kv5PtHNlG4J/sUiVXXvKuEZjkv0jk
/fpHDXt5PuCYrINQtp0MEwqmYGZwrAMf0IC26a+DuVys2g0w133eaBeXh73n
Bsf2QOHlOaVaV5gMXkKMRSrUnX/E3PfA9RjqOZGW7++22k1IVvVh4fnP3Lcz
5oTJmC1VZ8jQ2CzC5rfdnh3PSAtytyoq2zOgIGSseKtAhJiscZkqIUJComA6
8deKcnJTlfbEG5TsFet4wLSMHTXWDXuA2rwzNTZAvuYa031b9owV1CcW1gXQ
hFECIiC2ltCw7NKMUIiQupBx4UJAotw4U8CGSLjqzb8k7QGlTVVKNDX+cNzC
iF2AAqitK6JltxQhrxaXyxs2t2TVNw25jz9M9Ypn9h+JHiAo5ldcu6K+ALBI
/+zq4oKY5FZwK48YsQ3TIUG/4o69nY1s0q47ZprliBQT0sIV05S9+FzWbk/U
gdsNun1OKU5XUJJTtfDNtS1ySa+Id87QxW9wxcYPt1SsUtdYhaRKvJn54mY8
v/IQG53NR1IjkMuVReJ4Npr+czcp6zGTroPBeUMP6BmbLm7aLiS3MzoadsOu
TEttjOVEWxKdF2jm3UgWNQtfMI+dVGUiY7maAxI+woIgmf7DD70JXZsy4cNN
lpZMkokjHVyjAQk6+pd0u/O1kFj4oJFc8GGtdoh91D8NUbGkkvNRa7ami6qE
FMd/C2YTpYEU4VzJjzdwSP77OZMkGkGie197uIXDmlOFJcGQJe5Hv0he6LUN
BqB0kSEjO7aIWUZj+IIOWCWwAhHqpDGkVEkjE2D+k1wtpyCjV691xyjIQx7J
JxA7Hahrg7Y8b5QutpT4xXFfdNvjhr/Plk+b9ktgZthdkLoywdFoaezNlJ7/
+hHAYHj1xfbSpMyjY9tYflQKHNlvBpfGPaYcHm8ty5Mm0EFW12z9kxbgz1ep
dvI0hV55d9e8FeAERKmPfuhPsz3+ToakpViUF+lPATGuYntNuVDZQIheHiif
6G+Q2KFewh6llNN0I2HCfM2jt/kMrk9EvdSa8EQpTpqvBZIgAjlLK5G4XHjH
2JKR4TQuM9zVkPSKCYbBYn+6zIUpXGa79BqlPY9dV+LFHBKffSzAR2mFRbiM
N942s6zr1v8xQ5uSi2n34MinKSPZXv8T8PALxg7OHtNR94KTGK6fypxMndhO
+SV115j+yfChgx/XuIx7a43XHmiLkel/QYlltzEYidc+JL1qZqOj95CTWCDL
DSzHSkvtVYnM+BvrsrYcwRnMRPxlVVoSFmWbmbsdLdxhnwnEhXYkMh5YY2hJ
6fjnykbAqjPzYeGwKDy9C8Nuvmhru2PL15K0fg9ND9pJ24XAc48U1OGsmHjN
sGVOPkrWMFTd3lIHrnzQktqFgF/hCkOW7KlCwL6X8J9yhtNR9qDALkRTgAla
hHo4Ld+CMAnMv+vvfc33RpeH1xVoWFt1ukJ5p8vM5vhzbhreMfrihIS1frc6
Mg1dyC+EemsoRA7DOWh3rj1oSJ5yAAuYTz9TYU440Lnkz3UGrsk7U+I2EJzc
i6C72ZrYqiCNNcbQjGpno9JtvGVUR2U2scYTAWNjSmFcTRPbruvxvJTH9kp1
/etbqv8w1HMvUxdBIKXAf/94qdyKvADeIFSdz3XSK7GiJCqJl4KP5kbSzU3J
VlFTAf2FDEop0rAkvMR34OFyULXhtLbj39nCHRQBGpBg0W4OYqOHt++opSWc
JLhfTWNuIl6IY6VJkF7LvRINTz9ethh3SUjnzQ5CWmdIBDMpfROC0SqNClaN
Xza+xRwAfjdT1jB3bPiNaEq+/DAtL/ybyUChpy8ceiavwJPy8iKfIbIYIyoj
TBv5tLj/UeEPqJ5qxx+2MkdvWgASoCXN2zzsjmrBsR7OEdtXWNCHrYkgge/O
+DKg7NHWE1jhkeXyfa8ul/1bFjR2TEHLwMUuCozGBtCMcF8A8WUMqspBq4ej
g0eUorJgTJtuP+8eV6Hj4xQFDJ7IRXRMNEMN1TZpME4boh9HjLBrwWvq8ZqP
EEhd6JwCPFJnkgiDPwiCG28GXgO1dSaxTkxHP6pAXZ5XNQuSC0cO4CP9Ttie
Oia5V03af/SbqZGqzHF+SkctwlbqO7Dp9qh0Zhi7/k5dwsdoI2QQjn1nD5SG
DDKtG9uC1GFzRhmwDyUcI2QcNAtn0tmVcWDHyc5X3QlIFuc0LJu2BFkJEJXA
CM8CfdSunNzP+V/83BUyb1SoFAeuPQYfckT7BadIAQBthdgmOD4s+wV5mO0W
3i9sFMspwy8m9irB3o2m8nXaOO5VxWlZfbP4tWSYiyQ5x5pqeb2qr5s2GqnT
01Zc5adUgNH/YIN5L60pvFcmyaExnII3HIPZT4e6rHNNM3PTiiyx/fS34ksz
u6RGTDIgm+lBRdGPuEezGCAbd4BGtuTZYSj4opCM7AC+EZoMOXCwWU7CnILI
Xcv8wQxzkaU2nam0zSZ3PcDKPYhSQZPJ+dLxw7btETAlZjBRkEUWPzrkXn8B
Fupqr8zi+I6kAAA8SDIH25b592rjlkH5s47oQ2oeCqMUdBoFuLdsVUWwcadg
UiqGHjvMw9PgFOYG7tmYNuVlFuXUy4RNk8Bf0QNh1pw5JTAojgWpBpHnmnty
YSEXe5InC9BtlCPzCtDezilaDpU/4QtAYWF7PYLBy6tgMV5K3lfLCB1mZrNQ
/FFYYEIifEEjTKgSzrBEQoyj/XV+cHD2K4bH55oVUg0fgnz2tDYiij+XcuQ4
jQdrHJXsSZkHAuuuz872I+Oe6LlPCMSROeEZpcXdmphzKL0YY9enmMo+g5vx
t31fGaqzu7e2mYDcWHdNYma72qNx6NIEOBvwt6d33jy+u2lwiJK6UfnT5KLK
B1SuwZdVGsZ/loBqy9x8mEnw7jO1aXLLoRMIV28VsXY1wtzZBaJX2IbblSex
OIk7a2lIrMXoq8vZOlB88iu8lJyxQ1At2q516n1s+w+LZt+o6WEZLRQP1b6I
4aaon6LNIHUb9pyH+YrRtbO7PqeVjGT26zA4KsrjPCRkdgwX4ctWmbRLyiuw
O5nVetwQuWnP0hdrcWXgg7nI0YA/qVQE32e1hTkZtGqFUW9gqf3Rgx7PpQ31
v8DMdedwmzB/jn0Uvxh7HkSIRRn/vmLnL4w71wN1GvTIWVH2AKs2g6cp205K
2M5bBnF/yAiL9funNyBKqgjNpCi4nX9LiqBfYMKzUabltgoYiGf9RfJEpj6c
WZknKXSLdv80kJGxyWQSOZVeJ1LBf2GoHVSzkYweFeiBrtSLzPBPcwkCDl0N
K7rFDs7tkup0+/Di0HtaJjgPV5+rNhvyEOJxSGX39p4ABCFDs5yIpQL2WJgc
y1opa7CE/JyfePMQTJe579D6RV6G05HaCSEp+qZiBqosz3Fo2B7224j3bG5s
LP34DI66vykW/2MwRTs1QsjdrXOsFIV1qB9xLU8cOj4+XeG1MjlfgQcYPw7K
ZB1kb/wWOT26hW6h1zgBJvRAsxesAH6gvYi9lLT2CqwXYfe63qCh0Z0JiofN
mX8ovb633hSstOkCurbfqq1+s0lHvdbhh1uTwyYg5rMDx6DDJ2E/rh8fUKri
dBt71+wszbHHYd3rVIu5y5X3VGtxWf4a46kqWRFJxGY3c/UUVCCBBE6Oh565
FwtICj/bDmD/EbhLA1Y8N6D7l9pSpmJB2EwR+3aeDq/IZmUVOC4qwwKtn+En
HhSGddpUU0JsihmuLQH75BMT99KXYX5H8FGlXnx4nkB8HuWU0pFBpZZhM2zh
zz6WN0dwtMMYBmGuIFNCCFVPtVf4C3FnETurYWH0M8S0Xzu0FQTH43AvaYeJ
QKbr7MDecsQZlFjavgsLzcspehLZOXCa5R9N6xk+7IhTKvqW1LVzBg3gwWxf
n/Krm+Uf9JFURwWsS+ocWWxZNFWmUGRJqmbwWTGQi/HuUHPUB11baccIKthB
usom47f9TzDc1wOyrXndWMWH784SJR1tv6W9fndOZqGeEWfiVnfuBsyjNua6
o2aBEt+NyEw8fH0/VnOcYWQ+gCLOYBOo1YP7lBKbigLY2RgPh20tTM+5o+Em
ismM6tksodiunhrnOY5ftVoICKeJNztbjZDAMZgOySG1e8Y/j6TOsnXMdLpk
kJX4U1cx8vqwWb5g8tfPjOg0WZ1IIdtEaY3qlvdKggAIuPAPdl3ilODW44R2
dVN6/F7dYkz00xo2Ry2U8RETPCC4ee2zujxO+UZXP0OwwdtzUGv/ct0Z+HTU
DsfCqrx1Hi58bTOH3dvoAjOJAmagGNVws8Svd7psLqo45owy4Lno9RV/8uk0
GjP9cjGEU0tdRfzPKwrBDNoc8jaYbvJTZOiJ9mTz4v8QHDyCgP5egPS/yhLP
OM6XkN0SsVP6IaAL2NZZaZZBiYN5dxorJ2k68GlY7Yxr5rGFhriJqjjqoVvP
2WbZRISQrMW0DVln8u124Lzo4vxtb6N5iADYc5wbVs4nFUK8m8kr3NPr2qvC
G2moAiKIFR/2d3rzSdNRXwWuNzICAzCP1Kyqzn7yZELaRBc9jy7R1CSDqz5u
EcrNFzQbO1OYlENYJm8dnkaZNtqhgloco2B9DzEN+XX6KcNpr049lFFDfYi9
nDTwDuolz9h730wLZJrxTZcySE1vRQgRi7mmtGpYt4FkD+ExLi99pcoX4IeH
uO0tvXMXkuwFIGe/t+MoopDHnv8H0xhVCwpc+tc3/D/Hkg0s4xz8Ds963o6S
octZupT1C+IlDy2vmXY7IYPvi6mhlgKR9IBYAhvQVh9XjDGkDGSl+LLeYMMj
XjtI0ukkWpE4YQamM2mWwDCmPOZW1XT+CC3RgoH3nWuYAYELQ0dbhx/wHcOy
TkF+HcrBqYcJ7WDARFNIWbx+TCdaWEhS5yHpMsiHnK/zrKrX1MblRwE/WWtN
Ez6KEM5olVG12G571qCGPOF0RGiNcnkqwSQjLGWl4SGdncCy4kEZlRO4e5eh
U7g0pOJ1qwWJaq55LIR8zlNRIZT/Qrq93m1jEVG0C+draIgv9G/a0O+8bsVs
X1t1s1gTNzJHizQrU6NfrKNjsUDj2ngLCNWTY7sz7k4mubRsfJXzicQAxgbb
WF8IRrWaqywgaDaUBF0Om7JtxNZqsn0bPN46JLdlZTTB1CK/AEfW/0pHZHTw
nAp3EcvzFHF60c3Oml7TsfEmD/QSYdt4G4eKN9w4TYLuSOZj9O0y2IcWgfW4
2ZcgQ5CTnMwQ6r8I2O3K/mtMYg790VHQh5qk2mZcfBMAwpDahVYIFafZem4m
yQy6CCxC9Ty6scpIOVTQDP131HwYqvC0PnikEHyWUpxgnKbOUlIzIKuLdcru
XgT3mZifFjNXtzO0NgP0EFNIo0f4+OeU9jLDFBF/KVt9OfGWNkRgYlZOZBFP
VQZX0xCjtxLHKXeZf7rMSrYJ2qiTt/1+CZJRAO2n28pxFSMiyU9VVqjEpwPj
ObDVGfhhvwsiyImEqpf3D63FgmqFpC3knyhd1byQP1CekTbfokdxmUtY0qz6
SIfmpXje99qOVZTAcDkJ2VQwn+N2ccIYH8Uq6Hl2EZ7V8D+cxNyaqe7EkdQe
UN+iVGap8pqQ49VtscJQ8ryJog+hMH/ww871zz1dNI8h5/r8VgBooKfol/WQ
Mt52Q4Y6dhFucqtd9YMaG/WLwXwA8eNmoCFJ5fefrIP3q0A5jZijQUkea3Mm
ej7ofiEKpTdg4Bam+1Xu13rLzc1wM+OtZSB9+75wxfZsTNNZdlkvVxKJbLOx
nWsV7THE+kaOcLTehNpOSUBclqjGoWq5MsaUi5moB/ZUPWmxQb6uwPbYV8df
aaj5ZjVeVtuuzvd5ArOIUALoJxeZFHf2yOAIz0zlz0a+ztByjWyi20DdcjF4
ZaLV3oUB61whAZo1jQaAx1yIDqcl0LHak/Nqg5gLj4vPJtLwmnazDf3TMvy2
hNZGD7jPXXhIlzPgY3si1X68v7o/OaEsOQ21f3mQxyZY/tsUgpIhkAOJFV/Q
TX4BFLP3l2Se57fTxj2CH8idse8/jDNz5Zfwk0+6XPPHFyPpGepnu+ny+Kap
gJv32ag2oV5hyK8nc6vGm2c9QUEhau3CxLXgEr2KbdvMAtAizWV8x6/jyRio
mL7mVKcWyP4miQpUctsf9TKD5TKV+fE5aiYUcEVO5FGxkH3c/VwxJh0EEREu
M5geX0wvzbKLi1XpVNTcA3c45hBzPqyevwVALADswUE6NgO/6a/02deZCBFm
AGK2+Ce5+5hq/Ty02/GzR32cp7wvwvBkLdKqk5v+zaRjusvQJr3nWZtNgNNj
mqlQAHKSMrqYr49niHiX5aLPF/WTRKXbrtuRDsHSgyV3XNiZm2uaxrOGVI38
mhD0jLnbJsSANi8s9WHzVeJkV054Si9rW89v92aXP9kR3OHm3mrYRxEvZxD8
hGb7ZOaMxRINJlVcMT8J7GDfAvnmh/ZdKS2v0MliSyC7+MK24vyxXbF1J2Ps
7LuVAUrdrZ3/cN0OIkdxN0XyNK6k7f2tIVTEK2ZDjVFhTPKdH3GHhRIsUsmE
ON3bQj1WVyfjamp4L9I5NVsJafseRJniqRngIKSV+/G4iOHTuLl/B9jLY6wc
JySaDYCjp7F4/giUZ7Cwf3cAlgpvcRGD9zrLw0qNDPIQvskv8z7srb30YFKI
AY3bA7gh/DdNWsgiqY+6oRMlOPGBQq8vibV1B9oCeUPIzb40iruHxZQBzjz9
iJkyHBfbo04fEpGPSqX+NDm4Y2IwVlt/9TYnE9nYEY8GWryFrmyJhWofhvay
oiikWEShw6/FpQ+LkLO28b3a7aQYFTYCHJ7RGGeUI7c6eJ+QHW2gDQ296gXR
dEoZB1zP9kLIcus2QjzKQtNchmolw/X2OKlYQ4iy8/EiHjz0KbF2w1DZAavL
zVF4ybEgWWv1Faum0XOTH2gLzEpyINJlIi7Xtt/gURgRd5lWrF//gk5KvNgA
TOBQxN0xnV/D2Pyd2rsk3TbK/NKVpucxK6x7103ue5j6Lfec8KmDe4kpPCmx
YL6F05SjIp5G3ShitHu2YhQI6Eckf4X8W2Emrux3n++qtdm8qItaaO4Phwee
79wMCfNPa+evJ8zJkhX2gIz0U4jWzrLKHMPsqKYyDu4gT+IsFo2cjZyXO6TU
1icV7U3atPOurti4TdtBDXShRgSIWDHCX9B3T5u6b03qtJvIGo8iiDxLegt9
Do8ZX+OjVT+4GIihd+GPF/RxFIhgCuxM45q8g6PH/x7wivFREgPvLy9goEe7
mlAdE3hiTMloW0YqIDUXze4lYw678GDMIRpJOiQuRwsAXswzdlAnrBWz75Xo
lSRpcS/W2OLvrdULOx0qVuHjYGgoX/mg+tViI3Pm1TRslxTWsF8xJDm8+wev
SJRPD1kXb1QHp5S1UORVJh1JyRMAphx4BATi007CuT3oK/4m5S279P4FKJl4
42lhVFpdTzYZ04kxUxSD9vRCjZ3s91xiA3vQQDDQRe+/+iampeEDMDn5wO4R
v/1sVT2GYYoeY7c7744OSv35zD5ne9Jdt17rqoZTOi651N2oS0eUmEHxTw/c
vqvFYRsdShSNipaV8HPUW/SEaXotzTZq4fQCFnmSLVXvHA3cXb8OIj+U/pBk
7DOMRo29IIdBCZrEeZagoYIbB3r6dmIUeXoYZ1/OaNh5R9ScZ5Q+CsUJTnDy
1/0eOxnZxEIGpH/IB0S/xM+8xzieBuEgwQM567XrMkoLB37Lpu1UHZb4diaZ
lJj3Bvl5wMQG26n/eCkF+34NoUVA7+5dnmL9ya1yvpr0PZTTM7eyOqzAoGAG
vUhqjKLNdDd4w6mgeh14VWbl2Mh/8spYvLkziApewq2gDnRfXtuxsRSqX7nx
Mjsf+e8itp7c4l4hvPDR0OdUWB9P8cissXo1GyfvqcX+ES0T1MGt+FXQLzBg
OVXJ1bFIJxiYjz5WNJ1q9Y6AQGSVB8WdH17r+ds5fVCitG/Elkm9Mb60g+VL
1MsM9FaBoOsGdycn4yaWVwBnTbyAe04/VufbVqhSZO8EofHxPaGjOxgDkjV2
PE5Plu01Vv7wEwtQPH2/jBgWqpcP23R7+QSMZF6sHn1FvhhqJPlrfuskpbpi
KGtSpw7ElNnHPCD9YH/qex5hAZjvjrQAQ0zeA/6tO/U/zxPAvrO/QT7wfKtE
Ws/fmxFEXkB4cofC5HFbmwYTHKVUOOtXxOYL0j2wPfCBOPrdUK03/4qIH9sA
HzrO6qfWUuKz3p7eELUpVf/83pX4xcg1xejuRqLy3qGBg5IAR0+VwxQKYDrw
7uniPeSSc57mpDyDXH03mEObLnazogaNkPs7+U0ubtHqQ3DtcGSghfLiMAgW
v4N2Lqv4UerhBClNUyCzuuj1XKCqtmsz1g/0mBPgklQjpO0ED9uR8ovCufnC
Qac6bxYIoojhdK5ZDzLFsBJgJOM7aPj6cXzUL/2lJVGcAMsAFPm+thzc2liB
INcIyYo02rBf/WyCA0oNzz0uSdwZGdoUF1M263oW/pR0zlHLbQSh3icrr0pL
JoYVTC6cD3WqSUd2u8ajLtzo7PoGIaRUyKVGmIQ6XkNZ9fA+rLu3PAVodCFB
hpzSolYNgiGugDmE1Ipc8tRISy7k4vbLyXlJMHY8/yYTS3juZWUxOetXsvyO
jxO1q8LYeUFHDiqRcfX6llpcjW1irQuMkpaWihVTm+NxlPeGJfPtM1kW6j09
jSCuRDqM3vGc2p2kUu30EqTyfu+z0N7enY3xcm8hKH3wEcgVYr7mLmWc09AA
2ym354+i98NBxM3ZqKqrTtNXgWBLCd/OInrSL4mAZyUrnsEqt/yc+Xw6qnwn
XQSp6WT1ooLo8bMc6ZE7o/+Ht30TXYMqVpHDjb11IJdJ74d91vWsvRaPyZbJ
4k7s9lKDJpzt/5ndZ101D8JkhsPa1Kk9o2zQHYeGO9KTiLaYLB13WiN4pULZ
OdlyFWhOV4vfR+aYPOTlpYV8YFyavuBbX9n/Pfu++ZMHa5eyNeqQX8ULMTRT
BQHFk6x9lRGwSbpDNB/N/+MTTKwK+t6yAW+9nbn/QWJ1K2A73Pjjd92iONj4
1l5LRM3G5m3iz+ca3ljbIKGh+Gy5xoTLf5SDDjv9MkkhYT2EQax/5VcnQsZD
RlmLWZTjyQzwQmZAZ1RzVWHAiTA4BIqYhOp9fNjDq3iwGqi3V5Fxj0nk47wd
BBg8R3FYVpdcJS2Lb1erBeaPXi6k6nD3/2VR4yQKyCOpzNRQB55tF3TfVZq2
PJXWr0O99kjIsCePLma8uYlA86H84f0KWgH4xk5O2ZVvKgRkOeG0jowWljtQ
chBRLRAHmj0T1836zYfQMJxRU10Sis4KZdiBtSnDIL9ONtBHwVGJ7ky65UqW
HM5h8rXA1Axo6HNkvHNFfD5jPTYi3F9BycEmOC56lUEF3R0d3G5v8UIJU9c8
jD2lcZn9Mebq3jnLTUrjE0i6DWQD88fCs+q4GBiu4JqfTow9WwrDil+SpBmI
hs+u6N1IyYTiPzvqTLqAvfsjaI4z+h5ZX+HNCgfLeEmNc6VczAUTpEtizSP3
x6C6Ql9/GDQ0wjNGNCa8DpAxyOAQOZ4scXSUfraj+AGcpaoLeYvlnkHDiy1O
mWdWfisWNlKL1fL/b4q5hd4Lo+k2vt3Dy3HGwonH66yMgEjDOInc/ODbQtX6
3C/Tw8/3ATbhNPeqjG+IKPD2SQ6nbesrRzn5cyHDVK/IEJjFtIgW9iQT2EGP
Nrrgx5sDsUrNKuAwmKxYI7V4tI850xzKoUoVskHeoSz3tQDQRWXUo/7VrhiM
0UZCKXCrndZrEwANdGsGRtjPdhbZVQQgIq1X2LvvF/CEdPauhDUtl5C1xHo/
JirdAqQ78IDC6zeNFuZDKhtTiuEuCNkkpDPY4Jmz18gyKizSuqrfoE2nzbSN
OfVoOM3qAvzv28fC386h+J2b1jzENFf1g3hKR/O1U4FJ6IhFBkz8XDz0lmDf
A2C6WUMRvfNHkjbVFR16M23+r3JZ6RQ56ZW5aS6+lFYGZe9qtaEHiWuJOKhQ
WQcPU8igOi0pUaAhFDE1YeK3a5lhzaU11aRMmb6L7HWoMCMRB2THFw6IFdR0
1fkIqtIBqcHkfG6ukNtMcSXKhOvR5dgVxGNea3wHn5sn3u1p7C1Ril7jmWcc
jms9rS1xSwki2LgZVACE3bwx/2VZpHS5BdK5uTfctheRMO63v6SX+KtH1tzN
j0fh1bc43T0tVoSpanCV6QI6U03trS/pcTV3JpMkDe8pfPUMIgIFOUD+cyez
fZgRSsZthOaC1tBzCLkul29A8EV5wDUTG/sqLC0Ui94hE2OLIT8uQtj9i7Dp
kycodAJk9CFkh2P3Jx5FlcyacRgDvgcL1CG6f1xX3508TEo1W68WQ6H4VuT/
GRTWXKBedOcHYSPykDdS1KXiZjYL04K58rLmB2lV9YH2LWb+XfrT6RXPxSwW
SITQClttnsIJH5QzP2aCwcVuxEEgpj75aguFd30nqA7Jl5aMCsVHmFBqCc3c
WP9N25HxBnKMP0R6MlX8ZdhLTW1BQZC3lllQNV3iT5uJl4TbID94D5WHkS4K
2vZxK+G6Ed/kCUjEO1ESUdC3QhGzBuiU/27/kVCR8wUpMoxXTuxzUC4vIqPd
2ZkWrHHhJ21HB/eb6FgDmU4WfTPzU/vrxJLjo9MBvBDnGgeOoXgyf2eP/d5N
UD0U8DdaAzget/0KxVODk8jxpD59SoKSqEDwkRI3zwekXlJeZ5qhqK8B0U0p
YlqHn55oKY2BOwxUUNJiZZBfHVUbcPhfl55nQCvuq9rQHVf8O/pE03NGRlpK
Dr9Kxfc3ouXW9xoiFwumaVTkGqRgxtcuT4DdzHkyxwxTwxxcIG4JLiPRtY0b
qNVC3McESieroGYzW7XGAM/yBFn8SJ2QDP4/r6cHiAu4+kmN+suwfYJ1gs17
47wRZj/tl1yrqOyWP1Vm7bF8iiSRN0RqkzQfHpbyD3YqBcTMHljs2hwCqs92
G0ynzj1jkdiPlJ+irKNfUYfYeyOFhj+bG7eqlH93Hcu+WZ9q3TUcQtBXkLrR
0bl8+Mv0lp6zEETpPM+Yje2PXBGCCYxht3cDwI4/uCNrzC84jdS5nUr9mtJx
tBP433auQuRs4dXCN5MhUrj3yZZH39SgUctJEf7jx2cek34XNnHjcEr6gEi9
UPTlQ+lVYA3HY25ZnzyB+25LlWxIgtp8+n/gqHsQJkRczusmV5ZNZbxaCHuM
Ogb96fAI2IlD58T1VmEfAkP17IKYUwGPS8xm5WKQ65VPGD0ir7mWBiLS7LOg
1dbSiC2CI2NH3NmKCymvgxTY3As98XikIJLomYabrIeKWLLQrO3a2tb/Sqre
gAEggQ3MHG1qwEDIJdxVI7zu7Q041WAJzqZOWXR+penCK3Iw41GyfNv47YsI
O38gZVrJl79VB22X7q1yU4jMBJIm9jZhTf0MYMIbmtOmXRVFZLyRNYOirdzT
+/iEGMPIYUzNYEX5sr/FiMcfnloEi2HWQWbr+yzf1s/9pSC4yi6gBQl8fCag
RfITIRUK8KIMFAz44xgO/EvRyi/R2+J/b3gVB/5dZHPueq5Cfwhd6pcwpS1y
xMXK/+F0BW4WonzGgbkIXNk3B2W+IrhItKrRGIR+f3WDvZajD5EvcuZUE5Oj
bFENhTvkxmIP2zb1QX/6jSWwjdslWK9zE1nFZoU2CfzBf4feupIgjFdr/QRc
S7dB0tr7VxvzCMsyxjnprYPA76XinJpu+KgDV67rFXIlUcWyW33lgdbI45hH
lrR2RBXOTC1cLG2SyPvfzWWWC9kF9oRDQBfDMM+MwiKJ2wJNSRU8gggta/8k
WWBT94+xz2j4vyfLBmnujSx01Z98sRGNBdn4Egi90N2UyBZxne6kLDCDr0+u
a6fIeJmrC4H1q1EKbzc+BOrSE/spKGyxTQu7bDJi8B0qHncVvrTjAHGbWnct
e16yzYYUZnFAdl1Q4Wf4Kcxn9ueSB8WY+izT76a3THCGzCTFFVY5EAMrRulI
3ZkouCfGrj9hPFQxSt41CFJ+kZPpog0YDx9K/q+LNdeRhlOvEQ+SngApuCnG
cXBX0681sQRFbULHoCe3C7xnd8jeuDeGUMvgRux+WVrn7UMDP1+WaS67Bdr3
WbiY3b93CCHkm6XD/pEWwa59CSwsT4cpo1phK5yD3PHl52xNdtl1ptAWqa+P
GLPLYLz1F6D5SAmND84ADaVpkcNjlbLQKUz4mKM1eKT/JcIFMxjACskEdHZK
RTlZnmzaJE2m56xN7AlyrvQfD9R1/FEaC8y61OV79vF2GhgOiIXFiM9KTMa3
8fxShNmpSdRP8XHX3bi8Dpd5MkjqWc01b8FWF7/3J6q9kZF2EKhd3gBUc2Uy
vwxjyF2Qt7gu2JbLQQU74XWEEiEwHUSI8g61FPg3sr1YHoB7Lg7zW506i5na
W4LeBFl+6uGIfppxhHs85dLSlGPvwpBoS8LrB3z0B9/BLeI3fNjhP+1GKKCQ
aWF1HkNNPJBTfDqXGSo94E8o5p48k9TZ3lb7euHePXkP2v0FefyXW9JC2OVV
iIPy7KjquYwQcO8ukKBqW8IwYD8btll8onBIOnTMKjODIJJTGBD6TLQMY6tu
OHdnLztue2nrOvQATm07rvS6eIc3yvOZPx356Wkb0yDZrnskGBG3m6DSPfM4
Cj6Ljw73TaCU4Y2qSwu26Tvn7BnfdeHolZWsv9fVN+oxFsDPo80PCLsgJgEw
k1zTTqceR0WZPKEWvqtTuwuNyh+yZpzkG4V4kpjY46ELvoBeGT9sL3arajaz
JZszq8/50DYcHaMngIjiyVIpcWQzh+hU5uKdCg8sieODHYlRoATPj0Khv4re
SCAJVAiKYRcol/aEu1ssKqnbocQum24gOCYEOKl2DXHK/hanxxH0Yk1GGA61
pDTovfdQ2ojplLS1QI04OO6/mp54otTO/GuNs9RQlw1qI/1AotuaOmM04/1M
fs+UmLVftu7bj9L3EFy5EErWNCrOM6turR3mUxKutbLE7Z31iwwcP1t1dD8C
OnxkDbK1Do1hJrLwA8R85xpX1Pjt5r7aLo7a6ObBNBEZ7AZalzr3l05HPPR+
6WpK6BJYBfD4SiLKeUewC6f5wNXoJlmdXHoVk6iee7NZ4JPrJlAAYzEXrBcj
IZqJTyCja7aSDznoEjHwtU1imxSSNPZjGdvRNSNhEZCcoj3ingMfhDSSunOF
Rn8QdUay5V3hs0oIABRhSWErYItUVyROInC67+Q5OjXCTyDUMlmV3eAOEDss
F072ZyrsMg+gfUSoaf6rKHCsw1r+6fVSpSuzc/XhB0/eeCKZ6vGqoKTNlOZq
v+23o4Dip4TiPcdFjr07ranY3z8NUiqFh7lq+GxDrJHzIIXRUCNtGvucydMt
Ccporfdel5CF3Ce+5MkFudAMSl0A0x765RmkIfw8IlOLQDa3WasO6baZle4o
QZ0LLSzcky0hzoa0LZJYYz0Q92Nr7G9vDzjdIcqVcgWAOTYh3Um/mr5cdKhz
CGKzcGyg8xSDxdcheqJojMNLcMijS0O9i/9Y6P4IHmvb+PJbZ1nsGK+H1LiH
HV5IvYWE2byie9E//4NZacusrZjuXdISGKEuZKi5HTqdMEUiG54avb+JogUU
lPaiPVLeF12HhqRhjB3MMNEdKH3ssAY7Hx59MMkKrDe5gH+Wlwug1jvI9Ogu
8AA22WDPHcpK8cEMj+zvHuYAVlAy6Q+BtyfkDeTfQ1/JO8lDxI1V9rXW+bUd
3HfDoeWrSrySWBwL5AsQRCuz1UkBpH4FyVK2oeABDgyup78FtOUTlS1dGwlP
dOZbGgRj8K4+oDGptvPPa9nV6WbVxOnUL72riCRH6LCG5IWs1wY+ZeZvSWuq
HPlbEZ7olKlC9f7ASsmbBm6vLn1+dzTlyT/V8bKlIRrt4WOkDzLi/MaVrDtn
d6My1kYNxcgO+iVaWc3+sj1GHwz4wNDm0WC82/Au7Jt3/26wW3hymsTsUWga
bh46aKw1op1v4hcXahmnF1batGS8atKs3AOGdNj11Gxc7hlztNbliQ4x6DXO
I+S5suFx5EzybqfIu5xuaSvvC+9CCH9TSVFdpLnfuTXNDOE/Y9O5BhQZdu+s
sirYNMMIpXypPi2SkL7/P/rnxG7sHcVvlREEhzU+EqiPdvD1Aa0SW6yQA0Yw
t1Denka/UvWDkO/VrDoMjaEDEUmZKl95uUK9eCz/EkgRE3iwqELkF6Ijj4io
s+CT3131xZuCj9kalJscNZH1IRh5L7V4HbZ1En3lngRbi+4GoUBI9deU20EL
FFLTeKWhV4Ljmswx7X8m6WznvfatY0/oMkaRGbXh51zTcIdv1WgkxNv/LqkR
C4ycql2Nys1oQmQ66XunRwIjtUXGhn9VHLLGpQKIpEVEyQt+l24Jq/nVF2hd
8rZI45YBZN200Ny0wo+fOiJ4h7bMnLrpJ09VpCoH1AAAFZD4iPuJNzOPf4YU
XesMQlOS7tsb3tLjDFX/R765tju0vBEwaIvFMYIXUPVCGGB7s0symCQc1BgU
GLr/7kmqeOXODFY5Ez/yYwshALz3EYI7gnJEbJpekWN9qBpyBmBz+68mwTrf
roaIi0kJ5dxVcnmAWTyW3LZQq8HWycu/113khesQIKzqqNk+6fS5hS1fmqKF
GfXOzOuz6VpdF66Ze/kkcYmOBMQBEx5WRmDJbDrIrYfZxmUZx2LiSGVnrhGQ
rbja3yqQuR5+5zvtZTPnRpawTNdiWMR2cJinnh00tXe3CyGnfBrhqVNpeAmy
D7qb5JF9gXIrrCNdhcV1gIF1gYgJFBTZFNffbPfuLcE9FmZsDEAl/NIXU3Vd
iVRQq1RX+oE1ulUXOu95nNVKpZA7g/N5cacIaS7g5ecpImBdi9f8034LgF/C
EWEBoaxUHtuSkHYRi47U9UZYdXMcmGM6DOVafAY6jCsLb0xN0zvjqKpCnn2s
35Qy9wVhHrLCCDy07TeqHxeHn8mvOuSDTTlMysABUeCtdXlugubrEOW7dnVf
uth48J+nAoQ850cB/nTvi2FCqK/ZsQs0fH0vDh6QDCSg40VikNFGpqYXKswr
SAONu2ZAUWUuIgUlYaBhEBJlxdoqm1lk9kUa6gXMgwfYww+a3rzz9Kn2ovu0
vebYInVJBxijMFfw5NAQCSSrvto8QLg8fZN924jvuIB5QCees020kPJfTAZC
9Qj9pw1Zwo823J5Q6+GGhiKbKZcVMvZvoz+RAM1EJ3gIgKZ08vQsN03F0K1m
Z7Gb5+R1zQL6g6sYZGxE2P1wDr+dy1DUFxXQ49f2wgaDkx84Ie5RyBc4i+tQ
NawLURBpkmxdEe5Z8f/sx27mmIjCggT+F23FGM7higVrvPQCG9epvWeqZzTF
a/erkLblQHFEh9plzSvMumtzSStd+4CBfJhj0Ii0dN4vmBuGZnv6qybWKUMd
+/+vBxaKFHH5n+ftjyd3K/gZAj72CRXvkfYceua0nq4HiQju+trX/KfS1Og6
TuBhi3mKnvYmc8J28V+CKKfBXCHcbJhhqFa7foiJaUom7vO3HP+vapKAiEnW
sa1+Dck25gLSM/jRXGF/0+nwB5ODHvUGTcP8JDQDFX3sUrrgVgl+65DBX8M1
dprPw3OF+PJGqjNlNgnY0W4cl8klqaDFWrZ2OKmt8vaV0vCprYVSEITlTTLH
bY72pnTGdomx7rhU1mLNnaumnmU+cshedXdzKc1qc/am0NMU0Uvl8nOHgpDM
jpRUpC+4X1sZHegV8diMhTb53KnsS1+GOYtwvLYAinLO6iiO+ZPJPm2JVSqp
UfZBru9fLA4pgRzQG9VrKiRxbaK3LAvdA71+iBS1lcwGEBdT15cqRUzflR/a
tZ9EWhOq2BZGWWX73USFYWMnXgavc56PS8bJWlkYkHj5WgH34mEg5Z3Re8QV
FNLdlPK9EZdoMcWpE+GWkgcBt76orapqlC6xWmtGohl4mDlggQ0nXW2Zx5AH
0biL5zs5tvehWzqATaOd9Bsb3pXFReVcU8WV6Oa9d3tI2ZxWKcUP8U9Now+P
Y+hLiruRsF3qvcylddsEwBVBAzEmzG0wkb8sKl4aH5MR114+Wsq2dtVjD3Rt
TTDqp6QJPbBUB1Ei3Wqw7sxTUkSgBDIaAVtkXXc4yJDdDUGDfePpr0YExUyF
oo7yNGYX3rPHYrtfgO1i/OxuLf/9kdjy/sdVrtzWgDBPxCMWJfMokfyoRqJA
cfOZg1uV4NacgfkJprQEYrgyH0A227Olr25akVUFVvTaR7IFoz9akRsxFHs7
U9HzVnnWzrmKsZNL9Un552XEVJWO1SD9QrbsrGjpQBa3Mu2ljhvKgMKW6toR
KJ5PmkXuNWusgGY1e748V/8heEEup3I14y2+MpHN+gKQIa1OBlY4KtMch3F/
bw6HAFEWcdSmu4hAOgbmBxsU843fATrvedgRIB+Nroo6RjIvsSt0oDENTh6j
6JeyKOIjRXAYy9gEjgmUn2ar9aWb8Cfooy+U1UGRfDLU4UTGKbZNgnK5MSrt
uPG9TU3hbw2ZlegSEI3DKVqScF1O/jGSS1ZIr8bOsJn75pubKEaGz6Oi59Zw
TxU5V2Q0ae8RoGGxeFyE9Iv+iL6yLTz25TwElMxSpwkK4cQBC3W0V8mJ9n4y
DFXuebK9hMVswzYxeQJdP6skfuIKQSzqFtYhNBF/jtUAGtBHFY9h3QHvKnee
ciofF982dzbt7kijSvdg/gEopPovrHJgJU386djmWkeCZywpRcH3qJ5Tmdkg
klD/+3qkxQPwtL35cxsPbMAc4URfB3JBBpznEULEw3Kp2C5Krh5cBD4u/HyL
Zq/JY9J+yrL83WG69H5tHA8Xpa82gI/4dY9vPxIKCRTUAOl9tzT533p81nvW
8b/BaiC/q1ewEahinf9CZZAk/5eXhqdQaHkyDENP7MlnsyLkkk3dWwLFsXLR
d/POWeFBKbiRXHqXjsjU34tSHt2jMmdWu7rgB/A7COCx/ED464HxRhKD0MYG
bZ1Mu64jNAQVo5oR7UaaNmm7ejGzXSwgFTdoAz1r/wqrrN9Z7fBgb3EXWkES
MQrNlDpqNOHg//5gbHpBmCEDs8qbm3afnm7d84qgJ7qqXUbkSQ9f8HvBq16N
ejD2uOfbqDRp0pbm54nu0W9DhTJcuBuHPygW2s7DCKhgObpj//OaQBHndn6u
IZmQmyRma5j+ur6R5qA36DIQqBMEEXzVqLKeHlzTHsL+HLTLrBLrPGk6PndC
oa+fJAlpFjTv6bD19qPRAJZtQ5UqYw+RUi1MBpHSHGEvzb8TQN/+hN5rYYus
CMkbndFltlg8Vt6IZh5qkjcvrkoz6ra7FKnfWiVrGWy8u8BLBzpiPwH+XZSt
RAn0XwD3MEjlkpbv0Ma5spXwxoOMLUaAVr2zsSWI1ow8t44z/RBPuJeoSnMy
FZtT3lwmvaj26BRXiyqKI2KWAaXQjXCZCHmRDxzsucbWwTej520ewF5viryd
PmeXHOdgJQ5CNeJK0SQtBspo+LV2IG9xciltDJhBGz+2jj68f2aYIuFzWmmM
WR/itsIoSljo+eKBz7hYgbXQGdhrjPE1qSGNDMrnHJhOhuUGncTf8+dJc9qF
e75o6cZnapb7mkBDL9QgJAnyobK+x1rFTLM47enU5Qtmi0fo5mRRDyCLHtqL
/Kxl8xGXLPYkwXMj+ijI8SKINPihebmMvAkp/woyHS4gjflYWchbNxFA0rFO
gWdYX/12NSOCNW+VOuDBJ34U2aleNUsgGDVLSrhMYGe9OuR/07ooGWHNxcT0
T4N0KI2eepMjA/zqZlQB6/3q9G8RzsIVodt/vwPW+x/rd58j9HGTmgHktGNX
hqSz3tmJL8gU7/68AgyeTDRDxXLMA9V6GKh5H3H0AITVWBARzEMjhrEfgZFw
rlesF5QgCwwZmgqz7pNPdXe83YgoNUbE/tfhisSKu6VeLXx7+lTrnx2S8jMg
AzrbYBqCCYUEa41If1aZGJn7UJDacw9tjX+EURISr8a/9mzxfl0UaEeVXkaa
Nej3Ottp2qohL9OqAgQVFM9fU5aURxvP5t/1oiGp1aVqlJb3VSF1ntTbO8BE
h6y+Y6V0Nd/41np6gHc1YZtWSw1uVFqZPaD6WJcOyQM2XZyUQSWred43Kiz+
HvDe8Mfo7FGoONRayQqo9wHV0ezn4kPQh6bWVvd9NDZFL/nwi/K6F7Mw5x9g
pBlVnVySx7cLPfLKrEyxouJfNoFkRYYUPdruv4ahb2OTGXYzGPHvmACjHkKj
ohJYxuOGlXeBX4kijw4l5A6mzqcbBMTItmvXi6KYkJo+h72rxMQaJV5cLMmP
6LN8DchdDPL2hBtpRk3JcogHQj6kKYlxCv4ZMcyR8qcAiavX6TuF1/8J+eAz
+VqPy4KBZe10EEoOSE9lTP1VKGC0fDgVasmw2SOH4no5UKKNVz85uDwDvu2A
Jplhqu2OCRxA+jO+8KL8md0QTsGm4T/B84EmGeE8PxtQVqCVwp/4l+EzKXmi
E5j+hR8QW6GdAuaImc3OQESk/aZxvLqzaan5NTMsr14VYUhWdEb5PiiYorkC
eA6W7KCy14plhvf1TsC0YEWHZxVYf0WHKAyruduJ4XoVB1Hgw8JHY6n8+DSg
CrtDPr3K5cKOAa9JYV9y/ZFbeidVfvStY5sZ2LOGhl0ySqeALsQkYSANMTpG
qslCTPHYRrLn8I/zGG67/m77dwqieQq7qc+XoNvcmCng20Td/YIC+H4Jrc3a
I8E9xDKeNpcyzrYF3IqV1A3JM/X+dHJakRREh7CALkT7Ze/iOEgz+XbUx9it
tejoqzWe0JRczKcl69k0B2stBAq/8RKnhEaqnuq7gsEy1fXEVrsprOzbumXn
PRtBUP2tUDScEvmZ/yiItulsyFX+p6dPb7h58G3fxwz9eMq1hGpMY6h64H+C
RmFyhapp/3HQzTcABbd7c5Z64+O1aL9Q4uyaZypaGQBmB4+9Tp3ULEVihMik
+c54fxzh4DAnGY4rfLVtlwPv1syWUKPDBUe4OXocZgqor5v/ECPuiaKFjmJT
JnIVdgHFt9ZBaxtYpzGF2g+wDg5xM1b79qv9sKEGI7SjNJeljgQDc7BTSAJN
yo5bE4MT0vztQGUoZ+Rkh02VY0AKrVCF48yEiph37+kzs8unjw7hgcO20cXV
FbooJTnHC480ueO6x0sc+Y8EQg5Sy60As+tP2O3aYczPnzrQunttG0ELkKEL
Zet0BRFVq/iXgbCbrRirsBg5qEqdjGcpKzBPt7UTnvp3TitZQz8Aa4aLtw2V
d+Ul/eYCcXoXOPhq2JVMl9XLDqVzjbkiZ7IU/Ql37GCg4RUqZ4bR7qRyejJZ
iyU7k96+/QmQvXQZ96quySlVKBfyLPkQkw7Xlsm4VvjxPa4c7T0vxy1Ep/QZ
vXB4WoTQB43CsRK+uuzXFVZqlb+Wjj814qVUZmpYTEmX5IZjPohPawU9HFal
vxEspj3PHqtQ5bn1Q+DN+YcXZNt00WhZRxwlw9eNMwQqgraeXEG1q133BW4i
H9+QboE6T1sN89ko1FQrYZllseQC0NrYkrA1cnDQ/jDXLeOnNh+w4n2U8ZWv
w4upLk7Q9L5TqXEEf30VH6S7yslLtkkVAwr+m7lJiaGEAAXrNxWUhL1IZ2xK
nwqKIKUrrshs0R3jIMg+6o7c8lLdLHPS5aqBWnt8eycBxIxdO+X3ZlaTz93p
gWLUMYOaluNvzSe0UD3jErucsR14Q3yGxsPdTdeSMUdgYg2ipFdqtlxSTMuW
4wAv4oO2nAzVrDeGuF9k53pYDMqVB8FhOW0bh9FCIGRVFjMJPWUQno2GZ5Zm
+jYWeDesSYBYWBTe1Y8xONDc+c9g8ZXdoO16rmIdsbz1LcsYbNLzql+zYFyc
5vfHQvSuh7Eh0G5S2HEEsIVIaooMnvf1xLp0F1nPo0SFBWqSeXQwVRKltHPY
qSwB+5JpUn9wG9YUMhqut1QKstdCqvh3u4d4wo9Aafy/BsWpKa/U8TQW0eUm
g+6HkdUq+8knMoso89i8/ZUgpqCi8l619q7LoCxYxj29WZwPYhBdl1wLGnHU
4tKWVVErzil4gva8qBjDwXVE1bGesS60jwih92DmEGtrLZKoxzMKbi7DR6YR
Nxe8o0ZmqlsSMzYHrveOlICffmstaH9PKnhwBfnVQg0QupL5kagXbraqWCPI
jfyMkiTDDSh+YpPL86+G+d6Ilcls4w2k9Ak5ppjQf5Ag8bP442+K5XhEP0KG
+XWfmOwI6f8LY3jzgH/LcIJSZp8XLdctQOi2uTZ596De+UzBOiA6fODV5D+1
R20yfbHYZawV/kqZ55BB68eajU01nCR7a+vNZehLQRGa9LemLNFQr+TapbV2
kdAwjmdvPPmG0G1c2AJHXL8G4IKykRn/MVF1jHDQknHZwz1Racu49KE02rnj
sOFg6dPF67KbFERa4D39C+3iQtdJgFpIxM7Vh5u+PZt1yodLKlCqawuQTBhu
byHedtGCaN/4XhO0or7I5vzd3tcBchIW64D1PG0jeFLDbO/QTdxLYhrNCjTA
wQu4pW7IiWonDZQz807aeoFhTjNLH41VvIlZIf7mLXBwWIGxgqpSfUyApojc
EFv9biayKJT4wdTkt71wACgGucOHw46vXFSz8Mv5HguQWm1uxLuW2x7c5WzV
0bGZlhYWcVnsoyr3/wkaAuMjUBENkKvBTy/BeriHGR8v8jZ5pP6EDZmJ0hOM
lW41XPIxhxfB96x/axJD3AabfnayW+J/SbVV/0NeZ1hzlZ05ViRX0TzRW1px
H6B7w7TwmhqnvZpahBZXjVRwMQ65L2Gex9qdXAObTRtb2FpBUvnSy8nLd99C
FGSDks9ACy8bGosNq2GXQCoauqcz6a4pS7ntQO2vMLWs5fMixeFSJceAJc7C
dOR55gH8LOSDcm0sszsIBJfNcu7wQ+X7PlaZCPnb6fsJm3UlVjaHxpvzS2Op
T17jTY67NA+uWDv/t6B2Qcanst/N/7yvqgAm5WQ2LmxR7pDAuAXv0foY179v
1U0/pjmHsxvUC4bBaxW/4NnVDBPq42RYOidWf+C2sAX1cE28fLROg1ha0qCa
wuligYUKRJ8uHmuxCsobzUu51FEaYLAXwlmS3DPjgy5ZNtFw+XzOndLO8LKf
AobEsfYOjgvHpBeuToCbYlhG3Nt7cJutdLQ3gsgVQ/Tha6GXMjE1WHwEGFAu
K2zEaESunad7R1tx+FV7nARTgTznwGLMZJEDlqkGP6hA3vBjw2zIO1hiX2JS
qDsynQQeA2/zfwPAzbZ+W+tFOHzYxzkAZDLG52EdoUpvRKdKrowjiKGwKOuH
jS5COAJs1n+oXw4PfYG0AEP36AGjXyxHa5wp2VlYxM/V/6F6fATUwrRdzRF1
cLQZARvOsryq8lmnVOiGD920i6acFu6uAOtCtSRuhvKMCT/QRIsMmHwhb954
G7fNQmRIFM0IKZRt5hD+1ULyxgafEcgQbOMvxWRHNkzHs+irOQsNx0g7tFSx
dGXa2YpdQnWSnjyZ42sbjoFw3iGJvAW1sFi6BZqpFRdRvlF8DB1M3Zm6Bluz
AFRXAI8H86ie7870KzCwRO7LPSUJSZiyqt5seQObhM4iy4fMZ5d40MHBAAbi
It7ey3SJU+202cok5j3RriePHww4KCGzXhFd7xa5bqUr/QhVfzDTamxSV+l+
IaawslPJuFsg4xT1mOlA9CHOfK4iaGfpNbro+MEimMHlbeXun63oIKku2Exl
YWO48QOOvDe2b+pROHXJZxwg21weYSFPI3ccAaEaaVNO5mzIHfVcWAwpRfe2
MX+KU4sjD4rJDdPJeg81729auMyXCrUL9xOjT8r8Rta35BPgu0MFYsPuclOY
1f67maTB25OfflkwdYy5qa9HPxuBxGGQzgW4uN3e3FirQ8rmQV/xVuAh3vUF
wOBc2jc7WiYVlnJjSUBMjl52DZk059m1FtItFQfdRtPRVH9E5b1dSKG+Ft2g
pO/DPq77UhBtAh1qOVy1+gRWP8s7vzNQNiNKdG01TndbM0UNKgrYVjeEJIX2
EF7VTTitU40wo11rs5r5mGC2NXPj3BAhfZ9ilt9s3I4Ev1Hbxa88ltOc/7IT
nd/l1KRL7Aa2xHiQPtfXMAU+KU/3e3kLic/zkY+fxXamL+tYNhd81UFsS4jY
c7HNsXraaNwEoChAAuIdm1DW1TRnHL+0UPyzi1si/I0pG0Ro2SPqhtyEmkDE
rjNeovMBq+cQjfiPCKz0sUZt6jS3YmpVESLmlY00gqBTQVkn6RirMGXCyDyB
WuP1ukeMUU3JXocmVnRQpTzLIBxNj41R66xOJb3KOQLDZj3gyDQHxa/zeisJ
ZL56yNkYTLT+aiwRvhq68C9QjfLjcznjNUtPtYQb++nbMEXPbsPruOdqL/VB
I+4OpfFPt1ASXXD8Iz7EIdr9gBnQBzwzM/iBbL27P9qrc0TmhXN4Xt3Kjsnd
hPiixRFsu6W69WvF7rW/I/nE5wMIXyoKWNpXVomYKQ44wyMrQb/LHiAH7019
qsj+95iqVa3tZ9ojJlkkBY3sWZtbCXD6k/fQlQjGBHhyOJMhckHb0Y8Pd+R0
4pUclphl4GGEq0gayAqj0O0sd6XS0RT89q2u0Jtbm4hj2y+P7u4kSZfuiVMR
d43ijezxXGWsYTMkys0vl9juN/lzF2lRSsSz3u67jdSXV06LI0kZbkduAw4L
4vsHBPYtK29RMjnEgeD34XxJq2RF8dgersp1OQb2lieybzZnZp2ZBW6gd5Ce
yaXqFO44nXLTKy17dPe6nC4KrJDr9oRQagVTTy7UhjItFTETfqxRLOhBYPK9
GPD4yjEpZWEVIdU1OboVCccw26Vs8kjDrGJyExSH0ndXjBYtTM1dcQ/WoHOs
cja6e6Td9Xw3J6xRN4U+FL7eptt571jjUJ/gRAsW0pwNSSp9FFUZGhx9fF7Z
kwSgHKWUEfFkd+7uO085rVZVjwGxgwFYcwAg63D852GqCpJ39lHkQikHUu2W
WtjlYQrBFiGzH70YHiNCYSm2cjftMA45583ao6AbXMFy/UxDiGARBv7qcglq
dDyjjg15Z9W2j5XUkxta65ndj7TAVae8UEboi5V9UF5nZTOf01FVMRbUjfMp
wspPbva4ZmdBcCtYIBgcZ4K8vIFIyGYQqL5b44Glesk8NgyvLxP/6nyKOb4y
n0Z+2Kyc1fEkb3Zz4bzwvD7X9bEo96rwUtTWMRI56Rmv3hpQj3Zp+Upygj4H
q9WHiIcza65OPw6Dog6PVQpk3cl90XN4c/K2PSIpFYIO5Fj6oYFgnRHHdyia
+tI4WlG47/DU+oSrvfvn5QuX7R06MGh2epu3myPFctpbnQvi2GdqT1qlrNHL
IqNk1RIznild4MoaSYFmCrMe6rkNMLfMuMmbxi13Qh3O+yuWQNRWCYCNiyrZ
5vPb9sfH3CCX4jgUCwI0tF5lw/t/yV9MmrVTZGQZLeyBzo69uqMA1f2x+zNA
MbCvVm8P7q5XlpjEmhWIUNqLLIrsjGgm0JqBRHiYyS1z+H5lFwLEw4pe32hY
4Q7ZOGZrKc+JGueEvvZsBO+ucrVmSskT0Xp6E0rzzC4GRIAIz3dRlWJGO8Vs
ANFEQpWvyFmKUir3GqE6NnGhTHZacfjchLtvExxGezKJCmcsf72lCkX6Xt/s
lGPqShVhe5dWJGkXYmxY7tvZAOfuDFoUunyn3YsB9D2sv9sVfYgdo736GVdW
rtUgYL8KbCno+dOgdn8UgLL1pr34nyaVX12pBxRFwEbf66GDtn61S4bE0iYG
rIt8KNVaY8RGnmWbOKTiisc1LEYZyA0h96RlbbnM2+NhITZ90GIo5XtJSt6c
hyMVQ03ccDZ1fBKG5VknPtEvldCQthtB4hhsC+SKnsexc2YgFxlM5aPBY11g
S3+zUPUvsAdb5a7uP9PpzCZac4MSKigoFUeOQQfMTma2W+7zyz/0b6tAKSid
81CCt4zcT+UwF2oiWidPtq5c2jTONj+e/fKilXXqPzjEiBHbteizntAMdXLE
etHV6k1I7K84IZMuzDdt1Ov/wztG/PZQwLcrmlvjxtEyau4WOXUlNenV+7dg
dcmooOkMkYS9gHoe41EmJQ0qTSxVYU4vxfAoODh/Xm9xujSYgH6kI+ha/sRe
a1vADjSxiJ9ckL2ucGx3bYKHLHTYJEUSZyo6WEVoeftjaDxKmQjcgUKJMd7m
ZBCemRBCBysJ/teqydVugSYMZwVyb+OyPbRs6zFR1BI+CLX8M/URgx5yTq9p
EH/Q6yx/RN8aCWHeHOFQgFyxxj2tf63G9s/tmOLz+SxZQeMp5Q1wGv4OZ/uf
xRKIy+io4i41G57/xuqw8ql+RvHi9MK1t6NsEDSmhy6DELrq6VDiAC9yGDiW
rJXqlmEjsIMD7n2DAbjcCEifqIggKNEUI3iVmTga+0syU+i25whUD9TRe+2G
boCQHzJh2veMDzzW8Z964EGBqhsYMNJEB7t2+4zOeJJYvIznlVz03Z6yMCFZ
vgPOd2J///8N6pnBSL2YUGVFD4xHEQHYuQ5m97AP7TvIg3OzMbalpvIhGDn9
rXVzqjm9xYRv7/KOqAocKz2ivMd0YYk7xoKn77Z9ujisfYSd/EYguBbZc8k8
QUqjYLldmRENlJM3KuA25C4M1uelG5fiSW5GZ+if7epZlF+ReeZXrzKK4HOq
6Q7RMmHmzVypOuX65vMiwdGRwrPNTgDG3UHTF8y2hSA1KZ3xm8sWYZ6gGodn
nAiUK0rvPBOcnEfiPR4pqfy9yIsjY/uuyTELbscWA2nMG+qmx8yIwBPISdee
jSjAgIcFY4rVue+POj/Gx7CnMPgCXQyJQS6R1rpBmeUAB6sc/vI8DfovWugQ
NvDI0GoL6KYJF7JxjuSPQY7smdVBaG4biCQxeaanNE5HDZ8UqzcK4o6MasjV
YqKeyCBKVEKzR6/e+Jf+w9rz2B6ZN9SG/VuC0zVyh/aBlvD3w97W60clhFiG
cjPb42WPPMYPcNiPzA4rdEjwcBxE1x4hPDQBa37MDJQQCvZ+UoMIvwNpgW8w
01uV5PWxxFm9I1UF8EFBN7LUYCbOcYuaOksisdgp90R46TnRz06sAeCQWrld
BjOheta6HUXykA/DeCIC4Jp9HGo/cvAAdwC4X22nhwZIo9ILu0tvF/I2lKC8
u34xpLJYxeDxwxHTgkIGoKKBTr9PSiqQoWOtu2kwoVo5Mc0cqShzmg48pQJv
Yo5Xx3LO43OgICDmgnSm/oBtsMHApprm/kewbP7J+WVXDIJwdChNn8a2xlHB
a9i9j/zEbTnLnn9vi+p9CCJWcm9YuftRImz4r6HG3i4hkPUMWiaGSKTyR702
kbd55iZie3PtiyUVPNN5XYZDeEGfx2nNKZtYNBbaLlECD/KMODFwnH+Yo68R
kSWYpqqSvglyhFCR7tsCzCk9gptWBbQR1ZtT2ZHDb8vH01RusQHI3D72r4JI
oiXfErSkeLFQ9QrrQHgDK42mrjkVgSH4IDUQFIEwhXFEHS0gE4BsmK8Elw7i
Tx8S44WO4cKR0P1Dn4zq4jZjX3PScPOe7Wnvs1IVdXM7ICo6upGqtP4IY9K9
yT1JLvYB0URpq0yvE/YW5MakLOKs5Ccy8eAZxF1KdzAyMqfab0TNNZ1NrB5u
mlkUaj2x4CKT9+ifMgPxDCLvLYUWG+SdOfHPEGxdjSRNymJ5lDuym9oqr5il
5BvoKsmRuxdUMqWtuiEsrasq3sX+9WSbdZNz0DWB0lRjsGZQbEvfW2vZOzey
7dlTQQ2dTS7DaqvQ+U3I4Xtd5QT958SVOIb4UKbQ9KV8jJiwNCMobZJcFYGP
lPfUgrEeR9VLytEvP9GBVVJ2sTCHi/yRdeR2jC6vwnkmHGn/uD3TqjclYq7y
cm5GR733d/98ZT5gVB7G1tm7xMUzTTYnPPdrRVqr0LiL2qeTtqxT7x+odeMH
CBu1ajRoIY/wqPrZNglEmiY3gWtk6PT/QwxFtWO6c7Kp+2iKnT1BMFMhbGLp
wLr3Tg0qDggfs8ARxmiWBt10ol5joWhg/A+LM+ZSshPMGp9GgwE+P3Dm+NO9
7bA74rELXyzklX/CdgclZhZLd74s+EcGbBXICZgEhmbNuR+F8+scGf6a/gNP
ivaQx3AOcOkoHhzYKstWkaZQHb15KyNNQQj1lrdN0Et/cwPemrydXDA9NEOw
hQ+Y6X6l45EBO5zVqS7wgfbDNGpd93yr7wrbFhvlYlS+0M8Z2gIybXruF21n
A6MMGtjUY+3IjUp3Hv7DuuI0v+0Sp3Frl3ewezb+FuKDfFTTfHLzRLO8TzXt
x+wfFYCRyytJDLu76TP2xe6mDAR9DGZG6Rw66WBuQxrRfm2rLD0Ds8uHABro
z1tLQa3wfZ2yvg6iqEOve1NzeB/tAVzMz0158676uyVazwHtv1MTWzPEG/bk
aJDP4oc1/6zmHCdm3xa3D2nfUNFtiK2hH9+PA9PBd0qyHQ1GyHzG5v0zSDdB
cjgwkK+sAJbkrOzI4CyF/K16OeLUIeTR8LqquAi67+j/3Umyov/bgD3HrDK2
nyMayKtuwh8EiVwRLufRpidvTRJarkBiH13lZOYaxY4x4OqrKhxJhPCroaIi
X8DbEFI/HQxCxBRsqvC7WwYCQNDxSobFr62xnfDZ0lGAQR8lyQQJQa2GdTF0
1mLEqPygw4OCG65SnxtgvY4OoV6mSnlT+ckqy3lRV1RTyKKX2P/0n0qfL9/N
UvonbTN40P7klS3xOsgR6+iYjMwIZ6Xptbt3mVVQFeVAsK60zihidIFakU4U
4B1GjXW/QOp0RVoP2Y5WFhlSVIyMncy9dsv1rLFtHQiT5KNxnzqRJkbGhE7E
uFPlaSXOlP4h/iqhbAIa+f4HSEnktIJxq74XIArKbzRIAOsWsxkeO1EBtUoI
F347CzsYgMKtVVv+PKrWsBEuu5qNzJh8DOSh5QnfNRWFaM9Vn2X0FbcJ/vQH
iVBR971l7FGd2lPh1Iiz2QB9J3idjZftWQfloFraSJlQY78Lt3o1k3LD8KhM
MNwT65tbHf0Ha5Hxh9CmgTUe06YHvaIghrWZkD1xtbiVM1jgk+84nb5z5F5o
Vfw4ZYPQmhq4oGSFflGjbIY4+7+8Gw4ysG1ZYZoGx/RVVmMvvLCu6yatnynd
fty4BPi1rWrlXAnN1Ikxh2PyClPZCgtq41m1K9j7Z4OFoSM3wEBWijdZ0Olj
duCIXKgYBFwHyhl2gGJJg8UXPTh/Xbs6RfMH+UVyjXz43BsiaINmeCvhneCR
0T+sGeee5rU/Au3DU8YW3GWfsibX/ozc9kq0xoxpezRbQ+uhQijeNummKb19
Q47YiF8XqPJaZCQksDz2gmslV+At257YVpkwSL+qvSCaHhoryCi1jOMpdk7b
U2SsfpZEcEwjRfaY2iVSNlf8yq29tmIR2WI4GzKg95LqCbU6rOkZlrTH1lRK
J8ErtZbCwcGb3NZ4OYQz0HtWvWvhkHv0Ifb8J+NXFQwakmZD9tU29TO7o2h0
BheMOUuKToz9czeeqFNNMRwNouGRZf0gcmRr3zj1FJaLpPBiUirHgusV2Vvo
F8qB71OB2Q/okT9FA72+hoYU8OZ9AeM40Vxm967UmrslmyTGq5Le5C4LYl/7
HVrNUUoVD4ADjgXH0NXDrHmmLu8sVa1gOtxwhSqskWGRYJORBzbrJK3561cP
A8sj0Afwl1BIO4AF+lLdkeaRvyBGIXoc1Q0xfm0s3MWJB6E3fwHoh9LCdQ+G
AC/56uqiSVdMhYN/JTpesqZCZS/rIwGyO5ICDEuSTdvpql0qbWc+1nO2vrq6
ZvtNSv05XU+nuu3oIAYGdfPZKOW+CrVXJE8orSVM6WBfI6PVC3DfqocShZku
CdYcq5wjbR6v0Itwa2Z/orMe1wfhcRtOKoe84hmN/iAUOhCUvTkGZH8t3NgJ
OksCisytvkJgcciNt8cGCoXIL/qwIEosqpuTmv8Y+5zbo6U04/BY1/XLunSD
CNStyIybSXVZG/qlfHNsvT5hokEreRhpYylKLe1V8p/hf/MhO/8GfLmRKfx4
wUz0//1OsrvIkcNQqV+WybiasCiBNxWY6WsFCbCJlCIWmv5HFQPDId1Gt06K
+6qMKkCCJ+iqL9DcnW5W93dZBbYgv6PP+PhmcSO4V1yys+drOOybamk5NHhv
pATkFqRAQm73s8dGFlZg3KXPydzFBwud0LGwh6rSwh9scgIFGxyZYjU81W5N
Jf0KhvxIPPU2VvGXpxtYLn0URqxoXPewfajKZvSqn0deq7tjAg+DcyT7asSZ
i8wOHZZJY1g+u2/XUezlXhzghIGzN2P65S65gK+YN0bBbbcnYRTWVZTDHAFE
XdRHnijQg67aeHML3L+eI8+CeW8/I2Rwz0ozJRrpvjicJWJ1775m1Sj/rvR4
EbhmZkCouHtlMVe9bBHkhTqAbtQRY/9C6leGfvPiz2KIRsOaq7mSASpXZ7Vs
4IT5zzfMar6NlFufRLEiS59ok00CcN6ZqzyvpKSu5fCvO1SAnMEo4LX/8vJ5
ZF06FRyYvAfpCv6gREYM+dwdeEgA9x1rtvHiLAzyg/StkhdpJKOqJhs3SALX
nIW7+N+u2aLsFSqUuST9eejGslXB9BBBDq3F7QMOHnMY6ZRCBrvWPrGlt7fY
TiyiMO/+W8UMR0ZUH84Dd3Z0/IXLHcopzapNYHkhoFabkUgLo5qoVmEI9q1D
+T2sKtiXmbWgqbLVYrjnd0Keo6rag8912kg/KiQBbVwRwBzY1aHaQYW4t/KW
Q+L9COghP5oud1Dgzxv57AenKv9llp32VAzlcDC9us7Jf+h04YqPzvIf6nZj
4sqjg51Rpz+uuf4ngfseLlsOdCF4k/c2KOv5cGu5HHZQya13igOig5nX+h8g
Hsgz3AX2BihhMo9KQimPzNlYPLYSGvCfMxyvD9drPveCZh1X9+NTuaiaS+E9
4Kfor1reLfCOJLpH4PUYPKkxTkZ95JTX4BgitHfFy+nYxtKk8LGl408I31Q9
jyOpU7Tc5CkYq05h0WyK8sE0QjjZBAu1BuB4brP6KVbf/dTU1xDRVEdkatUB
wsZf8TkXN3v272Dx9qrJbAYiGm+HXdXKPAj5thBheFP9h4zkitgjicMkV6co
Gomu0GamELZMuXQkUN0TK+1ztfrZSfNb9MRDvoOQaZzy8kmyMPEILSx8HlHF
iNaxNATLT0U6lxTA5Ukf+VIc5oBVAFKxK5Fb4YP0Y4sInMrR9gZzLMBa50/+
yJ+6OmxSxAv/2U4RSU+kT7acNqzg8wIrYEzP/tAiNQza37WfDnUJk0f6c/Mb
znJVbYp62qHWDQX7tlUuzRHiJ6wGUDf8jEVVsNuzgWV2AQ7DRrnZX+V7FKn3
tRt8j1sLV50MlivYcJ0gP0rEWl8Hxs8p248Z4uw1dL4FlwiQEcWfZgoOaPD8
P4tUGb1K5SyWPpGS6pu6h7Qpk8nSDbMq+OvAcxd9eA363y1/t3ZwsmjWyKRh
dLDQMxajmqRNXC9NyCFa0Gcln49MVdiwIzdbC4XRfiVQkslp/b88Z3BCRi9p
jGD5DdCZEgwAsMX8PohZqGlH3HnbMfI7jeaN5dF6JqIKulYbsZLnnDB1pXkr
NIfinaxwO/SoQ7JzAh3q3UdcbJMdl4ao0M5zGyJECuno/zHB7jfIp/mPsU/4
IEi0W2xb+8QAxoRaD+z32lUY/h44YrREYFiZ/Abn6JWDHqblYayWJenEBJ3e
SoFzgIMq/dGkiwD3hJSONZWrHHc47WU2fgqeJJrnVVh2sdT7HXDNw6UdXbxs
aPYGTqJwaTB84uBPEqSDHlmCSwgRQy0chMy1FFkIPk4b+qN2cyH5QgvgRNCJ
tHl4TTeK2XsXoazwzhM/OIHE5NRRL19RI3LS4v7a4+xd7Ux2nA7ywwQhukd4
VGYqNyBKYACko9V419S9kmOGweJLK8SaOuMdEQv0UQey90vAMdOB07hsDzV/
IN9KTVmmnosK/AdIjw3X1QGN1ecvaJkCZKZzPYEanjCXY19zd44GcUGOTSh2
VNIxGbI8Houd3oAD2ue+lDvNZiKGKPVWVo2mqYLPbSnXgRsBCjSfNvLYLj2v
ik5w2GYT5N+HrlFIUAoJAS1RZvloLYnu4+lj4W40LkOnY5vnC1O51E/ex1F1
sHQvdJ7dwsvVumMscAzeJK09nNZ9QzauJhB/irImNNUhAWy7DGJKQEDhm5i4
38ODKbipz8WtcHjR+nFKSUlXewsFEVo+ErhR2vtCoTrYILU4N4H16Kho5nTW
9IhNx9ETytpXeEDzxvFH9A3Cci/VGN2iGgzT/4GUMe7I/myd79StObTE1jdc
PuQJIqzSJwSB4yaNnRiRS7PJWlnBMmd8wBD3BytSyp8ikFv3POD4Ops/era1
p7nUBTVPt66sGmvtc26gzae0cm0X5uOVnhY1f48xX9O3IRtqjpgW1gx1fWxn
EYjWLHsrfd0w76lrG/LV528jiL4fEvvtPsZCSAcAi1mgPV2RloCzEJDu+ap+
5tAWu8FQnbYU6rs7TLvVFq4Bla6jRAQrKdsZDdGS6aiLRNhgjAbGr/54un9f
ie4GmDxw7t0kOfqvvWiZHs1h7Lmf98TTEVP+32gQb3JnB0Tpm/ThFwrPMM8Q
BE1yfOWYpc0+wcGbUQi6yckRogQy+i6TWLXsC4E1/ElazETZK74dmN8NYy05
s+Zs4PzPQZfxYVybYI6Cv2yeZar+68JDD3h3h4ZD9wfFRKa+qw8bedT3Ld86
WrUCo91aS0dkiqiiBsRa4do3mSoV08sQKj7YwfE2dIyGxrgSd2DhUgde4ntR
K3SzQ8D37gg0K8lFuy3fEKQRMYw8SxcU9MHiDd7eZYWUVg9rACuDY26cjbyv
o5l+LmY0RgLT6MrqU9wdOBtXC3WrIu0UGKy6N6knpqGU5NXl3xS4XRiFyOsx
bNlCcHBg0qofOFe1RXLDLp/sIah5kCUSqTzJ3aPFOUiBPaoFx+qCsOG+fmKn
6Gi4y/0Su4J51YLXWR4Q6EObdH1wy03O4LvT3W9ryQoWDwNtDl9WiQD8lsHq
6E6Sq5e6hhPrw0WIpl931W+fj0M0uFEZmDk81uFbfzJvl4M11FWT7AJmcYXm
GjXbNyPkzQOACVBP/krZEKvrcEqqw8wON7RlSXIkPXAiYFeepDPDykppgZWT
9mNmTxc7oKRr4eRq/OsWDzWLs3Saur0iz9D4znRJeJYrRWGC6FBFGfG8Vqfi
6hherOW2NeIbMvlIJGtsV+QbWnrjRs4b1dTJKmurJQZOqgLHLFLLi2EX65qS
yJqe//TGko/9FznNmn1WkejnZyobUl0pBn3hPXmo9dI2jQ6v27ekz4h9gWJ6
DGFWk300GXHCCPwgVSZPE7UVb5nsGGCeBW3r+Q6ts8rzvyXJSziDjwRZJHOe
7Ot8s7hp9WaLRzb6OKwvO1UwjDMUQ3z91MFiiD8SgS9Lc67d4oB8FATB+yXf
zUk8grWKPypWoSLmXU0hXR4m7fQm2gwfRUKSi1+FKph3hnPqowQcJV7b0GyI
0Z/2i9+6SN0RNCFpqllSu3Qz2RfWRuDALSNx3d8d2zXAwzyZaJM6Xzp0+Hpy
HxfYCjLjdHvavpfUJAnbpkVte6+TC0DZ7ul0xImKx0TEL4m9kVeH0osGZcYz
kk8U7vqOsksyvtYc/gfGFfePH/pntHe0A2zMNRepNE8yXQ0KFAUNPZsy7GBJ
NicBvX0iMQmLbGF92y9xc45XPLna/7VviHiG9euBJAMPl53s6rfmJLAr7uIF
tsHdLIC748fTz0fE77hxy33ASu+1TSD7T4Q3E5mrm4y5MVEwc+MG4bxfBdZp
Lair106wOVlbX05DbscJDdpyxTiDnzUinx4zoh97SG+0kClbKN2nptcEb7Qf
Gy8DWmIttAclV7+95OkRtxnzBUrcb/haBtVWnElIXwz7dUM2bbByY35X3WOM
zZ/O26jbkUbR7khAwO1026WYNIl3dhz6SDh6fFaz3ANvfR4o0CMMlIWE7E3s
7sb/TQ3e9eM9kqnnFjZ8JBq1IMLdxIOPK45biJ3xrQ1CQnJqfttlDiIR6DlZ
a0DitJKxUW0LK+J4GkqUICwh3Nm0oiJwUeKmL/b+sPzKjo30YfRBX4ofMN7h
q0LUr+lxy+J1nfZ4OFIfrhSP1mp0usWImpHY9DYFYgqS/WikoyU7pBamvbVN
yhwrvG6jVattaIdNPKP1Mi/pmE8PuXJ31tUa/sRSx6f0fywYj+ZYqd2IVHHn
z4ORwLKBVFUmjOLD3mVwZSiV2sitWFJ/bs1ygvw3jsiCB2BiljcPOHKw4uoF
dqHAxCEopK2hT1fluko9EdQfuEVmu8MqB7k18tucgnxiD+1c672nQFnxSWVb
SVztV2il9t3FPVbjPvkEPPoWZi1mzj8THCMLvydsl3LyVVM9S4INqkkTUHAW
/Mr7j1pQnDCcN7fSNO70lDn5WCVFxPz3QM8ZqZ4wGVR6kyS8bEn9t/ksZSIn
cE09CznM1vF2nixFuEaeTv3J8A9TKIcDciOPnwvWchljbLgkLaCNsdol3+UW
4jbnlHJKAG4BlaCDIQBPD4cYcksSnWH8qltOh1rRA8xxmu3anfuiP50G9qMx
DWmvXYvS3ErSLUQa02vZN27NBG3rpN5r0iESo14t9QYBhtjMSCyqpvZKgi9P
01xRSOdDvKcobA4XjaYISmvv+bDfqjmZtcGivUQgieIWj9i1Uw0ZnP9c2isR
3DuC0GgahGHIEvmoYCrIotQbBg3vtctHVeDUrMJGhry2puNM0QNxjfiZ+dR9
BDmJVuDkf+I35uAqmI9Pw3+5Vu5qgRDokvPH6CnE2HgAE1yMMVqHhfLiSDLA
b1OkiHtzqKBYiy7Yl1/i//EKER5Zf1bA2n4FcGhoS2XoyN7jFOYywyKzlWRQ
qhakOYZsdt2TtjCQk/mZG+XEAY45se4/MpluLRwQT65hJl6IwFzg5FX4mvB9
pXPGUkB1SuVy10SECHY5onwCrynfaXgR11Lwqu3HtS5D4nkt4sRI0diwEiss
buQ6dhM1VkU6xFDdJehLYwe44KTi0lLgIMhjusC9lQlxS/+f4FW1zmucTLor
m2yntzHnhwxP4/T8+J6UqRzOWDlZfyKamo2LqWO1N6EJiYdxnDpbriF7yIqY
l6jfQqNEUgNiSW5ai1PQztbI2CwZzeMKQspqj0IojfSmbCFXfDZYh/xI2wF7
yP0i1hEUwxi0aIIUXtSP+8UtyzrzX3W3e2O9Wg857oWAqURReZF/DdSSpT/c
t7dXetCTbayjfljgY267NXWZTvwib2g3m3K2R2EMsSF1/lsFMnEel92hxEs1
4dgQUibs4gUc28R2q9N2YFKr9OhrypZVS6waSrLuCxyEfEEUjNSGBejeriwH
GaqMdr5yr1brliR5fFwjHs5IvLTOQrD6+rII5xcRHEtq8eGs64i5k4BmWm9r
n2YmPv30L027UU2HEhjeWRrnOSXuvrDEZvmwJNA2XlfjIqlu8IPKrTOeaxS7
ssfAJydoyIOVNMWmdKUHnJirZloTjpVf6qeZIBZLv+cuY6HUilVy/qcM0K52
1W5qLW7Qf7dgeAT8eke1M5bjsmBPfITtbZ/dAhdpSke3fe+DTdx5U6+Hh1z+
qSZaQEcLOipHTa9IwOm67jXpslRthNgzXleTHhKwnkSzpIhwROVu1zs5cfKv
eFjMLERKeMfuCkRUGYawjmzMXrgwf1UivPUKP/ospt9S9rnQr6p+28Y8s27R
htBx29HUX3a6kCWDWGc5Xu2WfDfqElTdgvLjraEB/DIP/aPjX7f6yZ1fBk9S
sDPyh5/yW7OmvU7ZC9ACizhhhdjvbTWYlAmDTDR00Q3GrsHaqdHfLLFDCsjo
9jBIVSL9CzP1CPw0CmfgttwODhlyRcLBe8AtWehwAPPhN3BSgK+fX7ylzy2Y
bNMwn/z+GTWzy1JqVs1H4ogzRVpf77ieWuj2dlxJrmOnJiXfwGQz9VdYDWN/
cF8xNAinwBeIkzeg0a1N1FOMqKv/Y2jVlJO22+LqZmsfWbLOXTk/CvIFd225
4YqAh12+q1rkYGaTBCv0GsK5GkwRjnhdfMg9hrgxthXPZThGsNiR3CKnDiG1
H0M14y6GPpalbCc9NTKYsm3Tz1s5Zc7xjfFCkthXQxc53YZKA+5SlOY8lBuU
R3XTRb+DcmPmwZoG7cZZuge7w2P8Iu5tuaPzXLtufI7jh0bJ8grc4LDrkoBJ
pj8W5TZ72OutW2cAbEFRhTdwxQIyXjYlZSv4jBkwnjqGw3bm2UZ6nirSt7aX
3o87lvjyrwtM0sG+qK2cxCr4NcPiBuEA8hBRp4uPQNLQhiL/uifGGdiD4K6A
HBYBbP4HX65c9WVZTHBSWlSR1gvBvfoLvpn1s1fZUlraYmXW3YtxWIM0KQGU
Idz0rXDpCtXZ85RhtMKoQ6SjQ1ViNom6dZUIrCSvNeuX7/U+w9fUfGQtKOXf
WrQcuSgfFCRenQrU7NrkgSbWjqznF06fTpKlaDrxucHKGEQ5BZ9G6+YGJLu4
xMjyi0mKbaIhvbfX/tPkQH/Nk1b4yRnmyNKO/WcC3v3ZbwsvUTdHskX/nVeG
2Sgyz3Ae+cowji7Gu5iiGXInxBZ5+qc62gGAw8suH4el9Oo+/PtxNxCindvR
DxZCd/aPUIkCayBIMRBtpXmKtImWYjLOBz5SAFGLLJQa50cjK4Tjy0hvwSk/
5hj8ngGUSoKM+cS+4plPEJt9+rwX2d+y9bcB2VGyA5arw7r2iPVlbqRMirEr
czehpDBTeoy5n/y32ofuzHvuZTCc13fyrLkp7pqgbGVPzOEez/rR2vObqiGP
t/hWsDpeJCYGr5R9z8C/gaxmU5L76qavz7cCD1MyA4N/Sjntxzt783uBL5U9
2GZg/26mSNZBiM8tVLKLyrWkFBmNhNUNJubYgurAv04A/Wc4O3gK277dHwf+
jhcHI/WdH2IjVxEPIgITOLgR02CFryuAlW+dRSd338FeZeFsO0ipUHade5du
vZ1AQek2HRLY/9zsatMLaOoGJlF3bmYLYxSdKDF2Bxx/SC0tLO+oyXORMndp
JypZxrIBVi6Y80+xO0egowu3BkzqRrRrVdi2EMDlPd4dl4+jJnJEETqqHPhg
eQ3cq46NE146tWlOA+aAZ7t8E/N0jHYmSMr2UuD0l+6PnG8pbmDewukoIZB/
QpQQBs4IDxBfsKGp9thPl9jojZpwt7I0QluggjmH2KG7ClwL7vg2UtPJWraD
Yp/HjN2YCgVDQwXDGE8oDmJTUiqqSLRXERqRF2kaCA5iZfWUatsRyj/SdFg2
+QZ8NPJhwk119oBB4gd/gBkv7NUb69UNq5teAaO5+sypjlFPqX5BJebNXuqp
JWAUm0UiwPNCDsk97K1qoOhrhZWNofIgmnpJxNuse6h2D9VwkPsJj0bx+iYv
YegcnHt8ZGY+FYig8H6pDLLfAbQ8y6TBanSVku7NMJqJYi8pI2jik81eJpIU
XsjisNLtc7zmbfpF/3QP8X5aPHg7MB3vADnuv5rV6d7upk7NQAwD88BpdQ5M
1UU+J7TCswX49PtZDqKiv6Igy4ojfnc7ha8aIWeV95n5mIhdHVfy7jbiNbXv
Zr0BuE1Mif9XCjQCwuatGUhXlB4Pugdt1ZpRyotkeU+NTwR9NCyfml4uFmas
qx7ve+TkYc0/j74repa9U4RmdRquFTB/qldepvYPOIxFr0tKJaUzC376eshE
3dttH0KiTz56U4j6alNReSoH2lK7DSxPcErG3ReJpGoXoCsz1HwPfIvaWX6M
3svkS+YFdHAo26D+gpBKAFf1UyxysPduc6f5wKHtqJiB6EeR08DTj4DatUIo
csJuveSKp8/3vOjrqfPzeSuFjdSFKUyaea+qa19kWHOPnlYrxZPWD4bCu0kk
//nwsBq4bxoJgdMu0+Suwfa4MalpzVQwe6kE6Tyk/aqm7yGeGMG8J1kEgEKL
I1HeAhoL6II0qS1vYuPG3DxbURoYOOXSnomOyD+4rzqPYL1G7Fn9uFy9Uigg
g/hbZZMoFJWJcITRRER+iC96AnMHfSQMkQYj2T7fs432fYJXMH1ZCVAY/ju6
7AHYB7v0LDQ/9udeAznMJGm3rynyJ5fACNwADwhyeTAmLOOuULuwGB4V+9he
KwxOiac1K4lB7ZVpEE51QIiIT/6tzlTM9W+9gzsK4YZn0r5z2b8TXyQOkcJn
YfRRvve+NM+RIoMMYR/6f9nemon2BPUhPwQtF7yColmhyiqQtuSOXzprs//A
YcdUYW6aYPEkSuOodSEjZEMUQ1a/9YzBbe5QtoU3mI0nfBc5cfd60LLwG0SL
1hHvwHm0kjgNm04xg11+iuapqBIrKdUr5JBZDF9BzTtpmufQ8RFgPu27jbK5
iw2a7fL1suec+1fLNHLx42j4Mk27hpJo2yum4Q0ANh+GQHffAGNLPHhGGO92
bGedQOoIPMGTHzoAMFyYF7NFbqrs16uhVwZiDUHJ35QGcluawWqIT7HmsR0j
683eart7gQtztU1E2fc4MfUSKk4dCWmgITJPzBJJwR+r9n4hfitzRgnfv0Kf
9R3V+g04VJX80/d1BY4euslgCHoRN5WiKIaaY+k4Z5ih8fGL8bLd0lwwd0HO
p48IXJQCkZqnYB9d8RDQTgchaqz7GBhStLhcjiFEszuJ18viuoYdyEN0+K3f
30F2DHsujXLvAGetBXPVuU4xWSnFvfAtU99qTZjb85C1JdmxxtlJ4eWsaVSF
lw+e7P6V3bWWqly9hbjPmHW9Av9mdUbmLY4OuIBBxW8KCYeyo4ic0ZT23tVR
3NVvUD0+HyG2fF7Equrhdlz4qF3O7rlypCpXKUURldBRPc7C+JN1oTIN+NfT
Byfwy54qlSwLPozhfWuHsI8UGqQDBuAT+8FXBimsRz9YnqsT8SXQLpdcMsB7
rZ3rP848d0LBiFjwVJxJhaRnCECtoHQdqV/JLSc7OZFt16kcjIl+9eLeXIFD
OO13clsu6RzAnFNMqkIceCYh648ys7Hkgj1zGeOscVhmXbFYX/oOfeJtq74j
rlWz+qLwYgxts8zIdZnzOA94/4Yvn6Ao9CwlOkJWRU532qY+icu1r3Jcw4Y9
eed9ZTAGISgFZkr2++wcDJDDkZulCsusFkgVa2a97O6D7FNbhgV3qVuhMVX+
tk0JV1DAkznXB8Yy4xe6h2hQnv/maOzWXHfCTfVc5Z/eICE+aASlhl1UOXw0
dnvqZVJzVzIVaKEcKgHyYO95oBjFQhBM43BtN7lgeP9wcCrZfZs7auZxeejZ
P0qQczc/Mgyo7nA0SbfHmwUelT6VbKuHxWrNCSDIQ4mKrYIKM8lXTmhmgNUn
Du30gxfRybH9quFsHq5pMa3/SXklcaKV24yPBbxhHlE+Bynk9NKLOjaXqLBi
tped/WLQNXh86qcMdaNFpQjA58PHRSjlyPqfscFzSQWiLOagpVFxX9+2FK3T
mCgbBSh+oByUPOHb9agUfHo7OhtXw278g16WV+WwbVaMOx2rjwFruicaUt53
I1mVcL0i6tFLLCXdmRyniulkWhjFwJb+unvNbAKfPe5t6QI3N0Mb4lHLNZ5M
ofHnNH0AJ+B5ItsFeJe7D/ztSNIM2QqQQ/dd+Rc43krRhNFV6CXgtMCvm60x
DiHf/TTK+HKFQeRh68UvU5bWP51BZHOeCoEi1UQinOJlp8CdSRIb5/nkEf5P
KW6ofzr/NndSMpj9TmCLBhRe/mGEpI0pFEsMZO/Hdz43Q+9XRIFXWhE3Irbc
ixSPR0paFpfjkUVZOJ8pMpqIwhywIbicrKr3ulc3fAf7lSgy5X4F2znRIOWj
iF83BES5RardxXZpMkim2IGy03hcBZ6i41teh0e3cpCAPKTAzaWSueF+jjiI
6XeDhjmv/0d/l6/UOgoWFMu2n1XZI+WKSPXl7RclSZ+D1HdnN+Lyulo3SjWD
Z0BI7ghjCLU4uFBJVQ90vl4fHlrAoBPuDCjKjDxfhkcaULnNeWYlOEqkdnvA
V26KXKtWp7HmfJEu2MChNypWbo7Y6m94GnXd+Y0Yo3SL03fmg+go5DU0TKgs
sVwuCL0JOUUutO6P1iIvD6AexN3HPPevgWdkwTxKF6tNGRwEHbn2yKMPeHrb
ELhoJMJFvDm8ypsWC6rQN5iuvrvWri4OiO+M87H8ODfgoQC94eQiBBcnU3fW
PNrmY8a6UhSOCQs7l8dJK4IKkDRTEdzVlD4KZCqm2+t5IWzUetQAMxtIkN0Y
9m3P6jbLpdcE1dmatFDbMZmJ8yDpWMVPGcjXauh9O8rr402NbWXUAXror+b3
ZaVKWWw1EWf5jQaYOVAKrImNBfavcVNDz6ApNNwQH5uqoAtQNgRs9lTgVgiU
KCYEDDsvlylwAZR5AmSBYGZuQi7ZkEI6MJPSm4Wg432l4FqUfwXPtSqb7jDb
LFmLcEVPHqUr8RWppfuIMBN2hrBCTSV9UzFR+28rLtCRuhp2p7MjKjskNvAm
nwGvRiUpROFL+EToMQ3P6uEDOlkp2gIGL3whYZ7bR/FaK9iv0Tmz9+L4oRdz
/xP8vXJAeZRoMYxplyC0XRsoG+/7N4Lz4rI+QOZcE5S5ikQOjem6xWbhDoc7
5XM/Ccs3xf1mCW5G2SiKp1x/dqF5Wim4U808wZKIw+0iaKpHLK3KHm2B54dI
xeFBP0OgkDrM/y1LAok9+cM4xoh8rOWZwWZVzTn9vmMHIodiEtTD+NhiEbm4
hsqmONl3uyQCCfhmjdi/eSV1Kcvn3pgfLp0o+Tymi0q2NkwyCwYB0AtVwfwQ
OR0UnIpPp6pmolidJhm9h2LnVFiGKADhdjfY6BI7pUNc6kKdZ0IsLbX7C2E3
Rvga7hSdaRd/pR6e0XjH7qEFqFPBY9D1GJkhyNi+E79bUvzWYxPyWLJL+OhZ
g/DMT75t5F7fdab1vmDXJokf0ZbHiJBitOB56Fu2EIbQeYosLnKd7ZZSvumG
HynIyMgRuicYjNBTdKwtHhv8mX+OyD54GIc+sq2UpdzDj6ux+mY5Xkg5SuCd
xnza6QgB9gxheQG+CysFIeNsQXVMkCqFCfhGe4PFuFiK4rc6Xt75MX6H+FIW
OZHErBw4szJjniW7EuA5NigGtaQTdBk4Nmw0h8rDZSm7Bjky5jws7PqfdisY
64E5e2WUGtn2A4hksOiRvQBjBzP1oe6Cy9XL+gAB0/zqmdCJVxjnkNkCQuG5
BKBTcUlFmz2iaPeOhjo0pHZ8yaAlWt0aCqNu4n4ZTu8fyjI4P0sfoTqZcOBr
cKszjejdV7Dp8KDvhe2ZbyY+Q++4gCoyvVhzi5mR4GqpF/VcaEaK2FZblRb6
Lw9yU+eBUV7iXnzXq/HPirtGiQBBoAlT/GBqWb9twarwyyZjQZjJTpdnacla
6MLbJhBE+onqcutb0ViZlYJKt51bxC9WJpWOSvTSNrq4zsMGxK8yfSVpBGO1
0yUEF7HvWHb048f5ppt0DTeUFpa1vI8oaapySTssn0zoPvKuXI6ltWtVjnJW
KO6+b8yPIfr7p0QHQBYyT6ucOlVS9t9zrEKO4awb9TSNWauvR4X5d47yTkhm
KWpbK8/NwWl7vGZ7uRlPt3SeZVPPGYTl/LRNLlwwuL2km6jij+NeWA4+aJdJ
o4IPAuScZkwLJ4mO7vK4xxqmYr8m6JS3+BUKzibzUeIO7rKkEggFpwiDrHyP
U+AjXcMczQgGMYp2nFAMwto95A6P/uReRqHg2ZgJqGpeBdvnddBDLLZOuRa/
dk3Ibo++ggzFYm7+NT1TYb2RtyP8XmyczsgnqhIkbIRi4B4YT6y5h31L6fQ8
cG0ZaeI20ra/MiWIVQ3Er1qNwEWEnTZtlLvj61qWwcftc+60qJunF5+IyRVd
nKHeQ5RckyfjFDVsxCbSS7IYLz1ASJ8YDVvFHdHGi6sbg4IGZZR0lXIJey0W
WnLM44/2P+Oddo4LtdpXcYuPTQVyDiurNOFs8ndwkaPAM9U5hHT3E+LeZsIg
ziI3h2xSTF97PKL41I7w53IXbvWaxPSBYPJrsM8/aILQHgxZQ74QRlCPFysq
6aVV8VVNSRqEUalSl75J2FR1YOHSqp+MCWgXLt8FhVEsOBSzZCe508JhkBme
G6/M+9snMrVbB09TZMrhMOmY7hfr2c4qmK6Ta0MC8Ve1X3Z/LZXEpJWkHbJK
f3tUwHgvOdHmY9rfRm1PTUVUl4B0rKFkccjsMGF0vJzX1kdwOTEy7W8erbmd
7eXqxpuQ2zZUIR4gg/38ANGclABfwYdv8Yy10FwjPqmueTKmSVms7Mq3cmvL
uoKE4jLUzRxpOjCxoFMeo3iiW9sgqT1k8FtSYu3qMXh6cxXik/Gr/Y+TOehn
grZyLwlaaaG2pKYnarFc8R1klWLwNoVrwwzV46wceuylhUrSvIsN07VRfw4q
t+C/gjg8BMyVc4b6uayJIlThK+I4++MN8nkoxMa8IECG3P1J4rH4U1Kc98W8
mizdVi/Yn1QF5jQS+IHthrjec47v7kkvcXwPfIYzINrn8yR+hZS1dW/io7kf
i2eWyvgQy0m0tbH/yhjvpMSbTCJDLDW6BQWN7mVF+I7/Wqf4lnSKaeykX+rE
j/bCazh6mn6d7NOaQyJYEeD15hCweyjD5IeaK12LRcrfGK5qAIqtHWcLg2F+
j5qc8NRkYYGs+EEwQ0cvhnD2LkeexFIh6CppBYyKHqz2SNGqxi3+BdygtBms
zaGIqpEimVfWIFyH/nj5f5A3rqJUM/j5vRqm2jQ64Yy5hYhRIuQ3WVAuXsUe
+FWzt56urZyXQqkV7XlureL1tCdmTLpaf9HS/JfDJZHal/iqwJh/TUNe35jr
P2ozKH0RwP3mA+4bCTtJOj2Pw6VBKOFgtt+J+vCCTHx936kiX5MUcG/J3TYX
Dhio4ludcY4KfglqisDUWa/fwq3/xvTsZ5eLqPjQ0wrNfW+pPgxi/96clH9U
vbHsmHbLDeQP81bSpceBre7LKoXPA/PSxuMSAoh+SkCjDWXXgcjdGhjYjVU5
e4em9h3n6uoC+PsMgffqo5E9jvHJ+Vd27wAhSksgyedGbetWgif0BsDT++Ue
KhpIVaoWmfTJVGId/uV1426WlTY7m6a6IicyRP+tn4XPtpPOcNCnPF5AD+oe
PWJ16ggIgbJZA/Cx8j3kq5FqUa+P2zulUW6xYXdBkWDur54suMnvM+TSkD4M
erLRIo7IvzrJlCmG2Zo1M3DOb+tPbLlPUY00A5GBDdxzr66/5qQ/0lFHA6t/
mLhH8RG8UxXI6ay5JTqEmSCRq+i8WM/MWZmoyDUD+aobNu9MahPN97i//NtI
uTESQ4FVUaPjuU4GP7BkKL1MPitVfcWz12vuYjcNVX5wkiXrCSLyS6yhaGjY
LrGpOL0+PBwg7dyZ8gHWLdS7EqKAgZuBR9WU4FkbCKfXIghVifoNh9qyuCKV
MWiUShN3iiImGkrWb2lFd6yWWgha4ooDWxb1HsM09Jlk9yWv8U7jTaMQ1Yn9
MdPTMZ+wshPZ6wl5ZOGrP7bCGoCQqzNyi8V6fUb98pVRnbF02LRyt1Kru9Gw
7BVgtBuytEYsAfnaw7gIOPAlCvaIMxJ8kR8w9ciUkWtQbLDTuW861P9IsPO0
KEFSswg90BsDVTeZwt2QCkqDwY1jd4kJdeMuwIiNUaoPTSXAOK+UlswhKBO/
DCmXp9dBEEeCCagZgoxayygBJd+HznZjDqGy7jUug6kR7NkVhRywgrbGXL0l
vnkJvu8nfKEgPYEj3gfOxRkp8Dg5I37bYS5+MXakY0yz8StKGyTS73ByZrCD
DKYoCbsTmOFziDy3RA4dKSlRkwC3HEu7pbvkhxt27SpGjUlfXJtgPbRjplSZ
GrdbjM9xEusR7wfjNKQm4eH4ujmucJVmk0Ox1H5xCpxNwaG3DZsZEraXVauw
N2nb7Lz969FzQ2rUjCK6oZCx9a8FT1cejX/T/G0/Kbgxaw/JQCjnbfWm1hos
3VQXXqiGD/TfJt4LFye5+ko4pSwe7K3yaMyJnlrC0I/VDHOC3BE+NK/tB0lj
Ne1C9dMWyx3ra6jwjiVhhYV1vDdn5IV6+0z2NE4pbMt9qejDKK/TbomWSHwA
nsrcBw6NM83mByZL6CsuFNo5xiRzAwocmmN0echTEYe66gj+HK13zuWSi9vi
qBL/09S3hq3ckSKpMWqJYiPEtidkxgdQb54Hst3F5ljGQgm5yFa0Sy5qBOwl
qaIMvSQDvJiw+UuME20aQQ5ynR1JfSGyRhFb+iyDQnd8Tc027fL/GY3496Dv
hrt7g2acXxcw8+AN8yq6tfxwnMnjfBWQAPoFP1JS1EgofQ+JXz4XPzqVQUZe
NlEsqiEhqsybU5YVy5tYYbuQv05q0B1atCLexeg/seRCbq4TmF7h71eV5TOk
Di8wtzevPY0ozeqPIBz/gwkxs5pnVMHBiim2owfbeEtdBHk+miTvd/bnGgxl
aEOFw51LWzvtOFhmPn0gqe5+/zSPaRXOdE59rKyv1m6Xx++R8p/kmiQ5Tn9g
jI59QcEQRTFwdjPyvyLKC8n26/nPkYbrx99zHkoZT3SRIZW8pJTm2i8PXZuU
/REeKbt6V0YDr47M7pbjtqZeQ678Z1ecJ6Qs0l7zXxp1znnT9DRy1yGfR8Tx
JItAhQDigvBV4/2O5Q3WBydkhWtUZ1zs4M6r3uSn2QQVjEWM6V8SdRNHqhJv
Ur4f7xeIihnXZHyPvUbHKO4hwXc/MPNaFY+Xq/9/D/F0kzXTOtnNNDekEHVH
kUwmQkBIb7AftaywwZALCtfi30n7QvXYiCVDoNEI1a/MJMdo2nTeYnzgPs6B
1rYDom/bfbn4mjLtEEe6KFUA4YB3YhOdL45oUNBRgDSuy1ueYYboec0sCPjx
O1EMTC8mZNWIGgbkDD7SLPYcNSsm85qbmUUdHYVHwQO2j3zwqHG7vj4JSXp8
OyyUY/ri2cBxqw5aPlS/+Nxqg9ZRh5ZzR2PZ9ckfPMmNUF1F4b2SUVvz77xb
VhzSdKH1lq9V3y7fnp+HUMhrF81d5fkVvwpODFg153rGcYEJxgX3tNF2ngti
1DPMOmuA9ED6/Stgx4Ibk3bEuCBAH11+8nr8947t+AeToRaIHpph60YgaGnR
KM/ArqT6gnnVbmF1AP+s7syDAbMqABQ9ub7YQHDx7kLm+iNKym8y7w3c4cEK
ClCBhYDMvU+JXNy4zHJIauqU6k7s233SkgNBPML/bGC9zx1zlvz8qPb+gZHY
W3yr9eYAPBmRnAWzT1kyUQR1w4oQRJG6BXKu3fpbNh3ygOI8YjDPwTYQr/53
GqAo88QUDqfbMHjvw5Pr3Bu7oexFmSOUsUWaiVsCWELflHxndXg+nryj1+5H
szVJaUQvelgEMzpFKWGGG7KiL5yJrocDIq/7LiwhgGiCfaxzPB45flvXM33s
R1oPfN45z2pVk/Kepcu8cWZf0mUbWlHlRJjapAX8gMV7DtsOna8ePKVJaIL+
qgzMXBd1gxbEC/7izmYQARZhTq+CNdNxi4hJ0JAtkyPxuA/gCZ/HUnZwxZzS
xYy9r46lUDVdEH1YAALr4S8UIGcP5pqVIFV8eLY8TFliXyPQOCYo8EkbrP1f
VMie8wGhT/zep/D+lGV43xPszcT41JFapR2Zzo4PDNdw0guFevtLdo4f1H1q
4FSFMU/mK/Uc5XPB5IK7qEXzIaMD0QHoZy5fBHN6sq5y1HldNyNtqCAnXOMN
8CkOEyM/O4pqVtJfMqecwLkL6pDUzvtSGdhYZTYvMN2csK0H2Pr/9jziDBSF
CV5ETl0/eBl9JsgsvIZwX93O5YqrrC02xKHxHIbC7YxYVBI2JRl9UsW4HXUj
XgLlybyfQ2Ntq31kBQL9C9/AFQb7hd1CRqA7QH6j+U+AasGhwda3JFm40qPK
mMVxhx3uWkOsAASBR+WCt78EjgcNM64wmTi9XN8uqUMcauK6Cv7YaJMpAoGl
7GxU5YRsvZLuK2PjwoKAWJssglHu6quSlDwmhja1lIof8in1LgNXk0xC4pJ7
YRnTftemBL2+BV3vLI/oT7hglAspLpZPTIbrYZixIja8JeXBkoyuoY8XQXu8
RiWS8djWEIkZsafTrNI43L9r4TVXQ1sRZZd46ybV5Skisdvh2gR2N21I+e38
ZI45hSptkgmJw2WxiN3ThVyhUkVkqjQF7LMdu3XABQYS+bmfvKs9OWPZIFM/
llbflpdiu6ty9eTNkKsuRvqLhRWGMn/+CGc7v4DGmE4LVwwDtnvtfymwvmlv
Jq8/S3G8VD15Icv0M7Arc6gDora1cnkIAxkXyPcsQLos5u0SJAPxdfuJDcOR
Kvm/Ih8FUgJ6IgUzeugPtdWCQY9tvnvcweIWIHW5ljNN1ssvJLXGoDmQGokU
lUxGSgJUvAXhjzpkcNztLOBARLMn/3clWuwnxKHndl8E6XwcLICK1EqeFKfe
ftC/t45LED1cGcK9lCwXW8+hNvOP/ChDA66Ue/rSIbVcinm+hB0auwiFKL8z
afpJmNZ9sMArk1DpMa7xafja7CAKby6w2ob0luJm9JxYcHujtn/q1P56BSt5
ZJMw8L8gSRnW92HgvXOdr+PsxiKv7yB6osjj1mKoeaIPvu4JKaRxkIzLi5qQ
YYSk8oUrjZ7WjEKIRnakjiAPblIzNxaaLz8wb/IlnS5qZfECGt+Bys8eQ1oH
ddAyWbFDEcEWPDDleNrNebcpUD3ckSbB4U8zoX6W4Nhr8RPaXLFtp/jRfX+G
e5fi4Q6NkQvY4d27Ydt/0vXNG+/riI/cwHnrpzmtqa3qB4PtALWZbx+txdPZ
S+6neWjM6PgykKk1SMKoHGe2RZ9QZhhz4Om1M/ImzIOi3Qm3QsFQavYA1oqj
r4Knukd2zbZcx/Ct2RvbjIsDKcXtWnTVl2pXrH7fMFP6u/qSm6Ypwi2GCpzC
zVB/qU7J5ck2FgeqcTt641nYyUhroXCX0yDtvskQwv/gvNGTecM4EUkVmSIP
IsBPnVz9/BAWd7684UncV/98Z2VEHf3pEi+eqE/yK6+GQL1Ls10G03uis4it
Q7u/sw8m4MizPbF5QGpEdQt+bhowXswEJ/XNr7zTF1RHKOnzGwGqt2R3Z4TF
Ayj3I1fLhwZHfkOsHpJzjwyMf1lnkEXNsAkjaMr5BEJGynX3j2OxOceYRVaB
3juwrVZ3zRRUiLbklqJ1a8R++EiC7GqkqnPxrxxT/DAQ/a8Rc2Ey2e3lU5cN
dgzmYju69Qr5E+txCrgtnQHKmc/5rTDjo2+WaVfeqnB92ZCz2LxEQC4OdQ7U
KrWf5QW0m9W9ta3Cn0Nq4evp0pWhAOwwqE0crDRJw1+v1I9fEokMPx+vQwdW
m+ESepvqvdixhSHgev75xCRV8402lJRROGRhmO1NksxH7X0hMCdA///EHzvc
6+M32RFBoGowb54n+pg2lcxTjC0hGWKIHHt5DVQqVk4p8a95LD09dEM/fh7Y
4hwPaCfjNOxA33p94Qua4Nv+LB4323gWb9mpODgm5HbKZpKF/WigkSHyjXnZ
tXWhGQhtAweUP6e8yrlgmSJ+dokShk/989kaWzfSFgRzKdTGkkLmTO4LF03y
7iPRe85iC8oFRmqxl5eTpSJSEnFEEEEkITeuy7EOzf26A5neK6BOHBxR09/I
evz0C5+Z6iqdRknRiuCBTCkNIqnrKHjhLCqrg9XoI/m2LqIU21uDaAcXZNWE
1+IqutS6lg6dQWRIHDRQPbNZ7atNOTHhPemya+dgn0Z2GCKQAQaCGrCQjYP4
/Ys7tb2TdCkN07AA+jEOjk35UzMGUyen6fxIZYpaJNSo6rF9z4UTU5ewBnsu
yAXOzKyeklfqdhGcRh+rkY1w3/ao2UVG1guRvgQ+77v160J48n5kubfM9kuI
qkWeKVf6+nQFffARkZWW2+RaF2d1CvMVwfpJSQeG2aqqmDRcEsGXJPZbKxyr
OpfGqlYFoCf8/e8qRF8443kDPF4EYE7EUOXN8XpDYXxvu7Tr5pf9raiIQs9P
cMKk4KhwDWdHkw/zMadrbcSqMsuQdquPBsZgLdMXgog++vpA9E6/freytfRi
UJ2kyc9F+9cSMmGkTXvsgYBkEFKMWLpN9aO7MPQHzLg3Yz/jEfNoVd8HZcqA
Z+l7e74sUstpaxVWZfmnlWxq0lyIZ8LjVjGlMy8D827oItpwZvT6qX5PcoAF
JnswTzUURxegb+8WTvCg3KX9WD2NTbmGUP404MynT9lRhQq0A8X/73I8GoS2
HkcYkH9GRxciYn56sJZ2fyW7eblmFUIKJ1Dn3aaBuRnKebUEOgYr9sXZxMt9
VP7jWraE1ohtc/76AllIkejBv+VS2vLs2Axfzgxy9n6If8whh0JZ4QGhp2XI
CXPO/RErGMur9pvsalRxWEOkCfwhLDCvgePXq8+C9YfzDUZLW5F7EweX3KsS
wIQFFTOzuOpLzbpFpZkCytxz5VkNyBUlcPkRoAcowmlY057pU0A6bCjXNnKA
3/mBX0tSW3lsTII1U4HeJNpXTVGQvqxN0ELwP32nEgelXXa9W01qzQB2MygM
8UF5u+6q5JRYJBsuSIJzT5e0vFhZEFmgJyff/U1WL2VkCqH9rjRmFgqs2BwR
IcKlgXjGAo7Lby1zOAJG7OBnM2BMU6qhDlArCQSql1OhyvJzAWIR2Nju6vuL
N8oank54EERAtIVI1U29N+2yewGJFqch2sokeRxnNCnBePmdSubkthUwZIju
cky9ohN1NGwHqZghKQ15IsVNoMxnDv/1HsJNW9WMV1HkSMgWrn9HBptjJjXx
ZCNC/Wm8maSWKljmWR5PTDhE3wlHMQnnCdbV1CzsZBVz3x1o0gBeaaWOgW/B
BThAgck0/uN6Ltd7O4xwLS5ei/ZgVN9X1uiLgeBG9GDkLPsPJ1lJrszQeLQF
0hfV5bcMSfrQb0vGI2uFVzmqk+6PnyyW9aG6lNB4SdneyjUwu2mShbVpl1Vb
4r0akLjQ8efkpvR4w9wZOLL3USP+3ZBntTzR28SSyHJ/ciBEOpb6BskYCWiy
1cCqTUTw0KlzZuF8JTX905WqUPP8xvOvCRxG9KQa0gjvmOLzBCmXrljNrxtq
HjpQgMrLJad47M0cTuUYuPfZUNBWcbPkbEeVJNudC930s+vtp9Zljxxpg3pQ
egFNLYxSYmqs8jqpp39RcF5qCkNoDa/UfqrWcEO3lX+PLTJd1yj7cmy0/iww
wm/4LFn5kZLJXXpxG/mBjvCE1cirMjb9yHmpmcYjraft9NYoGWVVHVV4SXDH
OdeATShIqy4yPra7dYymkKo9aMp5y3RNApbFPgKRLjJS9/wGYVW+hJ7zgcua
uNyZBVt3euiF+H48l8vc8iksitVA4H78TCYniu/Ms0wFi4s7TAL8VemXxM6R
qEooTw80fq011VAkw++LoAD6vntLQ9dyQhGada+Tiy2POkOt9+4n7FFtsl8x
i/eBfI6+yT7ozoQ6PaiuUstn5wIjqdRggdJswxe9PT14ShDSiWdHUrNAC5Hx
skOWMDcfd5iHTf8C3sVBQ9Sp0U63lTPfXvnOq1jmL7jzIFsHFS+vhj6xhk3e
MucBR6yOpKw1Op/YyZJuPo6gOWuTGaz+QiN3lJ49zQqfMmOwbIsnfkJpJjJk
m6thGVYjdk9fvWSq3Xqaps6th+uJthm4j2+idIKZ2rjYftOHHxYNM9p2nR5k
Yp0g6pcUhO1nIIcb4c9AYu4pwKS94VGQI95NsmwPtCiToBMR09WI+9ZJxRgx
lpXZT9ywFqfioEDSutFcOleZ9KPYc8gvAf7GnQNsWD5k5zpvsy3dW5CQlTBI
Oa225RGRLQ3DChYbpcM9ayWHofERrFKEHGSvL6QGWDgGKJMY1HFbNoeZ/Pfa
xsMbK2X4wcbgOQVprh539R1bRTX/NH4GxdVD4ZVm8M4kxTC7u+0cwc31EhDU
YnihwLL5d23CdSY2PLxTIZLzgxn3NCMTx2Oa4gVvnS8qFgO2pcaKy9QQ7dkB
FhI5m0DhfnPoNdFjv6kcPRIEGpJelxgh85FHkLI+VOxM4M6BbYSQ/WhQZO8X
hwZU34LGYytVuVNVIjKzc2N2zBqdyCrcCm7Z3MEtRjIfkfiXbUWATwZdP1CB
SgkpYra/vooVYcRYyRGtffG3T+zYJkZlWngohOifpOjgBb5J++0LdOrRfPao
w2bPs7sZkRHAmrKIt1PGe+wDN0a0LexQwRGrlhc5nogU4zbUMb+HIMekLExc
nSQSK7aTk+/cbpZg4WgRPsIRd2LnwAQWUjEQSCtBGQa7PYoh3TRupLa01yvF
erhWzl5EuircCydfoucGUOK5v34knI7A5AV44QSxvCg7hSuDDBoZI3NzT0xI
NqnYWyIWT00P7EGToKTX6dBNnkFNbqqytf2jNdQCSgYTiV0zpbnMjG1YOjnB
6emlKduo1ulMFWVsaUcXfehRai2wTEJ+42epw2cvqR3mnLERTgzUQ0n5Ta3k
laF1O8XT1xdLUKowWeQYfERgs8Pb88/Y81xkFYWVaNEgoRFvCeAZExokr1M4
hTQVhV4s7zuzJqtdFbh8XR4Uoe3DAHmEfR7NhqjZEMYMSXvvHNFqqV79nwjI
n3MjznO8I7fS1ZaxLEVdQfYLsW8c5EDDVscqgT20WVD/SRMuUQFx4Al+Cy1t
hgi13Z4KlhkT77Jd1SpjrFEYi/sx/7svnViFdKTy0LZUkGzIlwa82C1SZr8c
UqmevhXjtNE+NEXnt45pWmLMvZpJhaaflabX6l6/zVJiDSsEI2JgfJnC+KW6
xzxa+Xgb3++ALENPKsGMsDwCMCoRE+9iZNNDNFAhR6iH7k32pWsOFasQtyrj
8/a98Nfjae/CcPRC3da5puDQcvPbLGSvpMh3KYnUvvRvsJS09ZPoYqVrDW9R
wgwEFWoQZa1DJnajwMnMaOkVRKL+fSLGAUXLvB1TChDA3gVsJa8mjjsbiZJ4
MXYOYA2mR4Pob4Zx/4ImmW48EzCfEqQsgfMyDIPEWeqh3tZ5GSQ8kEf5d/TW
bJ8A5PeVvUmcDaJlH4z1SpR/yzMHFTQaVSLtb65Fff+H5A+upEJ2bhEulHjV
PyUV84ZWikCOulFZBB1DBl5w+u5a8jLKcgMaReWG7L0JylgG3Ns0HzGWlfgu
MeOioXVueyUD+mkbRz0C/H8Nkx5BBda8cf+MY/dRzPGEbvKdX7gIpGQTzASx
OLM4qClRjRFZRZ3r4VrN2UWs+gCTp8tJRuJkPiTcSXUGED7TMK68sfQQ/HZn
DxEbGoLpwNnFYwPSoQWdKatVkz1Vdc+1drDTQndNVCMO4wEQ1zjiVZmMusEC
GbSisNo2pNBB1GdKrbhG4vISfkD7X27+kdjrPulL87Ib6hjNgoGB9iNU0F/R
Rx927Td7i2K55WLoYxAlhQYfqq8RncIGqYdFELIP+Mabq0bXcyyJmHJQCBoW
NblJTnEN1w4iuFuVQVddgcZ/wptcpBuZR+JJgWyQisEKRKwaDvi7t7MyD69V
sYaitM/82jO62MqXhXHCQCYFOPX6Dz1F+rI2Cvzf4wPku052VOLzZwwHJhM5
Yy+6z37olvxbjKmHGdeHIsp12OvBHzY7ErNV6sy1eqAzj4uCokx49u6whBlB
MJ4bHX5UKszCsJzMYNGxyrD4vwPuEVjsVucyabSW+NXerW42Rz+EEEtVj1Cv
PUtVtVluE1yQdYV/WARt83VIgb+/UDdFdOgDSSShDqk6fMYopePi2qTGegFY
NgGNpSqzbEvyG/UeZuSjqkvsbmgCjXm1QKSS3kanikpovwnQkA4YAdkiPvGv
wFBuNXwGuVsBdXtEAEvICrTuB0P7p2Fo2+mMvt0Kb2alAVpM8tiPDcSJU9Pp
qHhob/tZ46evZEAeGZFBL0GPNiwQzGCDtyA2VIir4ByyI9gu2lp5Pcj4uV1E
pvmZyQxVj3S4OrTu1EycFtRkYBs21xe/g6+nSdRUOBvuW46U9RTFEZZTa5DL
tIeaKRpS19cqNi2qnSXubI5Ncvi3E+WnRPpF0MA84pGBdybA8McBztdXj1Ta
JP6eBy1Mdct8trfjoB0PPEKi2GYOWczTFwa3rZr1q5m5jAIaDEYMnMWFaRUH
s7dWQIxW/R4/EUFmwDzFP8GxMHU8G4I61WNIdzMzJc3UH3SmI75j6FdrW0mq
ylXbsYhbNLHP7Pn1Ie5fFXXtd33lghBNsJk66fIvxEFrAsppiQNfr1fPVDfs
TWvCIrez59A8c190dhiAi8+zid6zHbrOEIe7xjRcRm7shX+E6GbdCZDSuZvb
dUxO8oiNvGEIIRbBZRvZWljoqPSZszjYSjPZJZtwXBQmqksOzUfh8EW4xayL
2i79hHoH3gCwbc6TPcfFiuZh+j9gd6wtE9KwLuuIp2Dh3C0VNA+tpRpcJnpf
GxEKHyMXFFPY8+x+5ZcOxyuzBvU9g31TRx6uBGZaijXHULgcD9jA05/O7Fi7
IQ0aLr148ZO1LFwHvQaemuEXOMFJYqFEixdTG2abXOq/02kZ+N5P3jEgiWKn
Bdc2wQ47SOaqB1+WeibfqfmN7RUFRZTUE7b+xTscdjb5V+uEXyWul4J9rBwC
stDSphHP95bnUf/hxGmXp+15ZJrOR42DeseT5Mc/+J0qBsxZsDZ000apMU+i
mm94FzDEo7Y6u7c6wromKthGWkbtZhkJC9tG+mnpPLZ4PFh1h78uMAWwJTLS
IkJg+aNygXH9fI4JKiVpsB02ipI407FuyOyu0Hhi3dTEq5K+imBI8zpsnTA7
o87DQKzevreMJGmSA7Q9h1NTZPa85Y0BJksmBTxmvdCXVHKmIOTtJRsZibgE
R89h2VBO7DZcE7iXxS1sYYdunxqne4lxs7RxI6lvg2VbLBJuP6wtjnHCZCMr
kzKhFH4mR1MI/xMEWNm8TRFSV6VJa4lF2bAa0vUuDi+GM7n+J0ek8V+z8/gV
c+ltTaLROLq166m372iPdk1vD1ZXFc4fVNBab+Z7323w2MbemF/0xc1ASjPF
+ZnANR5p6lV2J3OUqGdpncdwCQzvFuLaxQGp+LAZhQP/ZUf/SSq9cn2clir6
z5LXmdFSiYs8mdTH1QSFllyiNKwYMmpy1cimt1FFQXKtpvrQUwqfClemoq/V
yNzbs+4onkG9FBsgpJrs58WTprip/nLhGMQePT+o296Z2llsZqQKV/lUq9+b
BrA5vmow/QimmkJhUxBESLA5ZS7s4a+7PAu/QEmfMrW9DdD0AVzdFagU6/fF
5xnLPFpdlfMFTaxpb+i1fOI+8HPkvTf3xLML7/nezCLkwPFeLU7lCqkNeE+H
FKeKH/L5RwPzSTLpScwSK/GBRcIwK/Yve7VrgJAnj3p8i+BXVgr8AKkPYRoD
5cyFyFsqKuiP5mUT8O7R0eMdySzwt0IVnsB/LqUu//Ezi7k5zhcNczZKPaz9
FFRyVUfFJsPabPYWndxOSZX4ivRnnD/P7DRowdoqB2Mu82lcIHhqtb1CWtUy
lgF8RzEXOUbAe4lgK2Q6FS8HDqa+7SKFFUu6hk4+55+51qaOCtmNT549otMF
VhJu/Lmf6A2FLQ4QEDYBG6pYbEhCWL3H6ZKoAAaTeZRj3mb5XMbusC3N061r
Ir14W4rJoMn4Bq/9y3WP2hzUGwO/DOEHbWCDg9nKX/HlFFXe0zac+/ND+sER
3NDLwvVF0qL4m1AqeC+9y3uS9b1Vt0PrHqjN+Yqhn8sXKx+ixXXSETaxVXCB
IWGKRgqo2Obz43xQ90RbzOla5X9GmcHfZfUyaqn/kTE+/O+wQ0y8kbdrYtno
lf9vEX9JIO+GX5wHCSqs1+RVgaPFIsNUQEKLbQompQ+G2VBMtsbaazPZzT45
pnQzDWnTVA4SFTYbwU4Mh8iMra8bmNxEs+Qn/eUsBWqyAzFdh0g1J/c2FKZ9
6c7mLND/fI1o7zTP8LbqJn8OJGBOawYigZgoAnXM4Tk5MIkMTA2PFrPUQpan
0tV8PWka97M2Nzc+6D4Cs4k50cZgBEb6T65iShpHYswFebyNryP5W4R9Bs+N
nRWDRrvdBMgOrqfQsAi/SBCwIXrPXcvHU7fjt8UyNXoaG67EIfB4YfQ2mHbc
etub4g1T3L9pFXwutASS98y0glUsYI1hmJ2xtAKES6YvzZ+fcq1AsUTtShE3
IQYtxfF+T5r6VHu58+Ak7BI9tiP2D6JjvwgeMWBasIcc+7Mj5717bM0Z4GKF
e1k309PisXIYOH3HSYt2+OuNDMSdDoBQG90u1hWTapiGg2LhUOLHNSK+c3/3
s2q1DshkHwhUiT7eCjl1QC0xZLRPqXCVz3zSkrnBSorUd5ee54baMGxW+Ad5
cHZy3MQHjxj+gEb0MP9aWMZGVTfYSC1uKlHdVkcZuiym9JvrSHwlOQJFbUCR
R94WRnHEvTUqIoDkARLBGHVAZRNwb6SsK6vkvSXW9apOxcCt9plkjVJbHsjp
cxKJd87nXZUBEwvTFnz4rEW5KKYTVv+wcMctV9JyvwWCYDiQ9cxpf6OBEEqk
20ViMv4EG15/h8m6rsye5L+nJYu9BamssLWl6d/JgKlPlxxX244zWt4Wwh6d
Zvzodv/How5mZtWzK55gSEVSZ+wctltIN7IgRvx8k6yvNCCgqzNtYTO2EA+M
cyLEl6ItEvquOh5onBlZ9G38GnwNgSadgjKnH/OQS9zv8XZOJouoIxhoPa1c
Zhc7xSy9WvXom4zU3KOApw4hCIU4klRTQ/VXJxWNl1tm6Tg5qYtXnuFSyHbk
Yi4dzL7rehOVGoCPEJ8qD/V5+5ykYqFk5zdWpZQ5whlNs5ru4eSROGqfry7q
mql/t+UmryS/Lazkj2iQBRzFwWwLnTzNDvcnvOeQI35CSWa5lKqGyqI+jKXD
losJ0EnXqVf1MISDF7WJgNOFy/BWN4SjgkfWbhpzfgzRaFsSRRplXRBb6ltN
3mpijZh9eHsiKMSUJSqOHmPwLj7qMFnTwZZzCwTiHVKnFRJdAhS3KqAyV/pH
35TnY5f5maA8fdG0Ampur9cwZlUA2hIcGW/aXBrTMwySslRuTYO8sSUNGCas
Di0BWpLb5mcYtBa4Y6ls0K89j3qQR9ziKzX3zdxHYlljo72gYOaKa5OX7kss
CsROofyOjUTGOScPIUeiJhz58NoK/sHI3jfE09rU/mYZi9J3bcVVDv+96QIT
nP4eQqye+5R32NnuXiRI+58FKRm1EGoT4T7td3/3HR2rxKb5VXjflxZA3lfB
kVBT8Dw6b8RGCsbeGFDDGfvZp1ZhAwpX4Vh8itUgYZfY9cJpX7RuPso7nPhO
txcVoju0UkhmrqI44ly2S+aPFFSNy4om8ZLDjTuiqyJ73Bmk7bwMdAGXDgxX
djJZ7kVSKGxr6uSKFtu26gIfKab3cuZmijQOjKtasd/iwQZ0mqLzl8NNrOB0
MfWB66iC0c9nfxD/enMJMPBOz/EeqdmKAfsudZlB/ovvrLgXMOv7NjCQcjsw
5n/TWlLUGpdZzqeJpq2whtNGm4jz2zoPn18P3yvezjq7HZuej2XuyJKVHkNo
Vfds7hirm9XHONmxFx+At8SJk8cXGltjPB1BfWq51jgGAy8zgSLuI3WYM96r
B+yHXHfqsOH7sXXQXvkwEX0NnLR3IJzAjSpj86bubU+US9RcsQTKrnXQKmr7
7zQwM5NrkH3Q+zxlgEiYatWSVLZGeaAs5bpfwESKS9GVJ6oHzEpxHZyblOf3
DmFyCrtVSaHKg9sWVcaGGD8hBrv0u8NjcMZvofAC+K4xKiSZrinpAcyW1JcY
ZDlBUflwXo00wRS+4UdSD7F4qBpfjwLHi+j0Bi1mZtxnRiWx4CuOY/C291In
tmY6jCOjpBUoxe6a4qRqEfWuYbX7tzDvgMKTc91t6WJdcXJb9nVd17C+FXiN
WBBwii76UMQwm5/35t4cJTYyJ7XaAkvnRzPQfW6RpUFeDeMKIQIip+T/iNx6
1PKyuAC7oSEnR46Hr8/KUKRfXgprWB2gCRjG9chnaYl7oRNiwHlSybrd3V23
bCR75Rci0wAPX/vPpMCH/PPT1/6vb5cn3P8qFKwiJTfAoIswMolOU2F1XWXw
tLC9gtdNztH4sPUIZdpazwJH3PJgwJGLRxfkI+g5jx8REEmJOJCtOdlvfeSa
OheYz5Jzk9NQF6jGIdX6B5+rR5eip1QhOp7IkvdmepOVHwUBNeLmNbfoMk8i
Zs8XVIotFsTASynv655E34BEH1wHwiP0A/3rFItavvT3kHjGkrB0t7fjVaOH
PEfYUhNo4hmmvQh9eIL7Gg2ZjNwJu2DVT+jXdDa6MaFPU5L3hlR1KJohIv2Z
33qtJEUTxB3sR2OQV9ne5IkeN36TTwLv+Rl7+V+oVwYFzNZbCcV3mRCDl75r
+MTgVF0GT4oPey1HZ8Ld5p1WhbjDW/2QihpLqEUS/hzsLiH7sB7NtJkGcYBr
t+wPMXg74b9AWyO/TzmrkuibRTxKCjsZwO+pN87wmhcyC8iO72IleSkvwp8h
6amBUZlBUEylshwkqXkfyJfFPmRASgyoHk5kelj4vRYIwEgg7kdvuKhTGoOX
txdTr9iiskgimUdqqZVEjL5vCaDZwd70VZgYXBfzLrFakjdCH+vQAbWSEyLQ
58xykZWHjciTQyxxBHPfksCy3B6KepPeSrar8DkpoOG5xuX8+Z8zMnLsRMwC
qJpB9MW7vWjcw/6/olMbNw0+iBnZRl/vhLZs8e37ikgIqzqrbZx8q/c9xRVb
4NyaJPTIZLFbDUx44pjVMmnNuIhfl5AuUH4+mRp1rG0ojO9S+hpIHUIGyXoR
0Q7DQkvDqwyR4i88MXK48RX2CY6H6mSkeSmlXF99TvaCbGjUwNtmH8Yu6non
CrPIWrT0saU7kSRUCcjtGERGz//7CQCSxi3tjnYPLULbiRS4D3rLDchnIaSd
2t1ZXYllhr3NhzNQ52ssx3CV8QOFarJkyLuIE8RqyBHyfPA3fAFZwGEmxEMT
6Sj6/7LRUqndHeJVRLy58w8/Tv/aF3Pda6GelMB1CNoS8BhZpPwHRTaN1ST/
43H4/K+d06L6VnnKgn32/5CgP9KVXBuzd1iQ641F1pXYBZk1pQE+jTrZ/wt2
FXErQbRLf68UmT/fdRQtpNtpVwDZGcsJkqLqsU2+/9VO2XgpR13G7e2BHmLt
pWa/FazNKiDersgU1g6VpIh5PBGdSk2E9VlQ2szWxqxhnFQ14QY9OeRwP6uN
O0sHjNTWHSbCZD/bM4Rk7t0w2zrH+i0sw4Lz75Yr7kq9RisIuRNLKkgw00IO
llDPAGkrx4L9At5fTWmdxGZxBFq1elDcVYp8OVqbOkPsbtlibwfsRwrsK2PL
hzO4I8u63+rajzYJaPr9TM3tB/OwNToSF2eqhQmqoWC6IWk5GK02avcNfUDr
I8YS0pn8o0cWc6Hb9XoSNDDOt0XzaTy01yZM0K7YEAM8k2XooGpxXu4eWG4Y
XntmXlmjuWP8t7DMT2DgS67Asm7WMePve+zYn2C3GPgQ6iBWd2RvBhJgzSGI
WRlvuR4zHV4xMFvKs7wNibHAcKdrNFCEI7ca3LoxIfrh0OEl0vatAOhtTPc2
256KZz5fLk0JMoYJCGkiLixFHJZX2i93byAQGzLKbD9i/WeMJozdXPpbLQow
+1EoKgInNQl1xugNWJSOBNzipmnRFMlJGaSW3wLsSCHf622EdK0hEKLHBCEk
FU50p/U47PPgKa01kOy/H/wiJpT8IzUZJH63yx53twbUoHpVBzSTL+D2bHIS
g+zxkkHyA1eXVTtGKzWTtglxFS6pZct6ukmMDRV3RN5GQDdHkB9u8OA2lS7d
wbNUdp4Mu18tv2009jftGbVArr05vdGdZJTRlahu509DG6lnymZw1fzUs+V7
LYaQnfiehFLVzp1bxzHV3C82qaJPfZvWHP6jhSFV+GG55iyzGHTYbHK53L88
BPswi/3uw1LrfaBt1rTe7JVg+AUdGVUbJJRESd+aZgBcUggGr0cCX9YtNwvJ
7TwHKHi3apeIGM8kTV/03CzeR1sR34RMheR/JLkwW8VhY8hWJuRw0vdsddmq
gy/DkpndbXLe7dKFpEHi7yXJszP/Fqd6YlG6w9rbIcT2sqGiCWuO/mmZ8Hwc
gXSu32Rq406PTScx5BnnXnP3GmFJQUfddAx+po3yK2KPww1kOAdATC2cxBIo
AybODN8+Y0DSowbNXduRQqNtW98FixUWxnP0jNrlhOJvVvbiODB2s4kjA/3y
vLgzuJiLzJyrJ/IEksYaIUcKg5bYQDAx86p8hA0SUMquQ1JdwflwPr9zbobm
J8xenSiiK6G5yWM9wSGbcDqJhaVGfpcOFgtcvD/YGPJFuiacPRzGU4W/ooV0
fJ1UIVV8pY4hD+MaIpGPhxq0P7Cb39eXdjUzi3W/Diq1WG3+Oh2ZENVe2Fzg
Vx93tKvIjHDlEjbrm5b9AgDVNTdEo4tyYEOI2/V0700vZmqINYNAV9ioSXLp
v8S9xA98xwV1q7jLoCMFIGTaw0tTTJFLX3syhlWB1BNALgkj1TImSwe4fheP
EoeAc+3JX2MzAaEMddwgo2galHL9/oO3Z5vGzz1NyGC/miPql0Wxzb3hWoPh
QdLfLKNOf9utJXmYTYTsCbu4FNS5EsqXFxFuqQH+Shi2Zn3Dz8YxuuBYLqxU
0GZBe+XN7dMqflrsv5+1bWbiWsOPDkAYGZ1LaXvIuS95zx6XnK2x1aRHmEWn
TZOHteDe3mIDYokuHPdyeKqlnGsezchVh3BL4lGcv+6SUWZnPTNmCkvpMr+w
qP1xh1tXTIcNGNaYx+6A4gC/V8ETCfYjMYHRStyHsuBo6Jq1N1s3/PCFPtjs
sLZZ+EHOKwO6cYxZD+LAIKydXuIkFUB664C6u+JjiIBL56MleZHG4YzI5b6w
PTmDzknM+RkuLnJ5NB40BER7fF3B0Top1xIq0hMnmaqaajRM6mYJtlp+ynL+
aiDckm33LeqmDM940ps814Q0SssZ9md9BGETjr3QtTvzdBHsSxCTg7go/f/Y
E+9VbJ+i/L3bsLtywwDrzZcDf1UmtbRmAlXbQLjIt8tSOEoJsMD/RtE2E7Eb
85Pp/OLliZ7nekRwvtqeUs2Quw1FP3WhG3PnlBtJ9ZYhwa5ftlPmR8YSihDp
5jltGiYztOfGaAYMIDASrGiTBQQmpyiAooj5QvZo6vHC0rFZQiE7ABP4ZJwO
54zYbiaSkM3nwbxxVKse/PHdx18UgrcB74wW7oiFyXe0mmtaiudvtu+kmG58
dJluSjQu7inuloYbMm4LVXUOg9w4YuaF4RTwKKtV82stC3xZKc3K9oUOzTij
6ev5N2tsVZAfr8u6AJy6BzoTx4onjeRLZDwHmGGcjldIIzYKQ8QVoHzFqxTy
D4o1Tag4i0c+wK9TYgg4UQvETjGCpyIiaojM3iyQLHS21W6U6izo3mJ0Aozt
KMi7E4LQJUVkfJjtmJ7fggX9yamRzLTonzxfEErlSKnefA/EfI/uDkQqiUnV
aZpWmQUbTIMEHbmzDNhVcFsFuNvlNrJDXvYW5BPbYpvnt7Xwjr0wKoWBwl2q
kpjUD17mT7neknyEV8mUvz4sBqz3W2H3izGZpLuliADFtBAvCeW+Rf4B84w3
s0qmvJWQS5BgNsOaZtJLic/RQShE13Gjo7BKSWzT7cFwQMO0PstNK1FJcL2g
rv8eVDKKd/kG5pvL+y2196o1wewefrhlEyQZNnYai/+3B9XKMbyvAfU67YZp
KxlbjBLN7dYdyeYU5DAWpD/n1wdIzJCuL+2ameUvEyjU0D/HIiMy5LA3XEOv
yDvqay7E9E43OSaI6o1u+NeH3av/71GbRWmDtYAtKf5VQUMb/PNmKbkbH12G
5ldKuMkRZANichotX5P7e+QRQo4TaOdBM+vL40RAdpytHtU81VSgmK9NVQqb
CbZjoyWb4zkML5vdhZdCdzdsHZlSuIe+z47zTdV3CzWyTsfNJp2KxAQuv2dH
fbP1vG/e2dm3Zy6U7EEFO4rwGZie3wVc3OQ94Sjqd/kj5ScvGTLxOnjyh1yl
uSXocPwjBHpLpqmax0mt1GL+Di7FX2UVdr5yYvqQQsQz3HrwM69fSGkbfP1l
vBB1Tw3NVcvxI3mtoLUXMDmmOVcWKe7DTvPp+6YfGxwp7e3JlfrH3GafNd5I
Tat5j1K5peWz6Y9KKf7QyDyQLzdjzZOnJN5+czdqLhO/3tTjbNnQGfFFr2Qm
8q7BrUk3CF6ywGE1r3AmfmiC2z9N3cLjcV01q187Isv0kg7i1LtpmhWJZuMx
JISwhK3UsRZf3aEc2cQ5ctpobOGvzoB+nRhmAPmPW2yftc8ltRYPWNpqn0zP
sCKOdETA/3OrDt80qu2pnSbU3nzY+d9lDb1bhBwZOPuDBI03ziBFKaB/H/mb
GRy8bT6NhzVwMmdQ+eu0yPiVP6p+kze2erDOGkIilfHuoamWG7cmo0doyUlw
+2qWSc6omvyYbWxJn3KFGC2Zm+JPzUc7bzmgo+pTVOvBRecWT5k4zK6lOIqU
TQPiKUp4pmIloMTQsWvh5lRvmsliCR/8ECPNUBE/REiZdXezIWOLYBIHQs6n
UeRRZAbcrMxLUU8APq/m/4oQzawk2bezQpuQhEPuyFWUXDoSfl5Bv8ogv1OA
5ohvL6A55tcadTnnSCQotcrU41nn2MhuR+4bV7x2iI4gLgWZH+IJU+Cyq56a
l9jnYB2SbuJCV0HgOqaqy3akma9D8+VbvPck1Ywi6BqaPHfC15ztO8zvEL9H
EK3nq+4D78gAWG+6Cwxeqy6PL8G2gSg6OeFvTwmR9m2TccaiSwRjOerIc12h
OW6Y7WdBEWNLgAHrVhylnJ2wVCLoEmSjHkS1ALkCtrtmNZV2j34pmm10dYBx
npAjwDms3DKhtQMlhStMsFsLLv+vFQY4DYCxXmNtF6JPH6Q9ZkJxEeL+Ixbx
zX3hthJGXA2qIWHSS1n/bGLytHt5Eak14uS4tID779ro0cSf0xzF8Zg2y0ad
bGRI0GEsHNG73jwLP3sJFbs5lemIp4WDLT8aMQXpsp9f0OEcuTJ4EtQWTBrU
yBv3Dnl3GEB5lUMpTeutFlJ8q3A0f6NpSstEG4H4hTPDvUW+w3ekXmxb0enp
5MMsHFjrGcEy6fzeUonpxpbJaHRRHjkMU5g34OILkpX9EZpsjiWzIk6iUXvX
t5OvVupFO5B2FxFRPkr2H2XxEUmWueVXxwBPpzQ5SZHSRy3Z1kx21n/Xjsim
BU+WYbtJ4bLT8rpBpplyOrCsnaNbrJ9NoGlJGZUDHVRpxaSEa0rW8+dyG2pT
XeaRalKLSfOALsLLXjnJssSJaGtYLQSjtTFoxGsVi632FQfJd1JwmYUismCo
SjtCX7ZSn5CYQ6kAcUeWeCHEyYYkb1e/zSAPemLYsQGCYYB9qdGrDI+pEoq5
oyOK9tL8/d8KRnMSFdzK0/Hz+AmCA2WGBKMbMx/gqN33ATmz+nE5XjTP0MNZ
0FyElb4kEejpo24sRegRv3kudXdfVZSSlhDsvQHoUs/vCGXgvCVm1kuofBJt
TALdQeEPlkJw4dU6oA+2M1/Yu7uP2/ieCJe8boIxmm0q+6ERPch+mNGY1vjz
CVIV578wOZJVZfUgDcx0vwEYvanxbowLZAVs+J2z13DUFf+J6Z04Uk/TO3rf
kBCto2yYIqxPwUcF9Wv28pdECXpGH1Adq4bBB34etVq4U351Po5/EKAZpyeI
eiraKsEWlWNKZyxWRmI5+pCdt1/nx7AxvHtA8WTQTU1cHVeWuJmB4FPGrgBL
GM8J3SUD1CmMBPZXyC2MW6DdzxEQKm9Ao/2AVg0TpydeDRZ8Rm394hsEsnDh
UVNwYbVWHiLeNFqNMNcpBTGHaNJZkm7jW6EqPnh9JdWQfKFpr8etS9u3q+MP
4kF11C+KNh93yKrFaSJy1BFERjqLDOloM4eHTlgK3dQ/29FlulqYCf4lIgCW
/SiG4iFY/PkrIfXULeuiNMQG2jW1OSMyaNCxID+3dZS7uVrr1c75zMKY//WB
NWcV4LFgnfNDS39kQNcIQsFGm6JgJUwTZ5P2sN4tEvMRcfIcRGmDPARIPeKz
HBkfbVd2EQJEVfOG8HQcySeFMZW42EmOAyypri6ChXEZHnoi38GVYRjHBEPD
CjAmeMxqwqYFDNE/JXgROx0V223zdHDzrRj+veahR+ol7j8CQC5MFC/XFZbA
JAsaK8jay8HYXtpE1HRkpXiQDRIxIY87vKZjr5dBazTJd1TKoEQlE/iIy8NZ
OguS99BC2EOeqay8oR7llIwr5MbrnBCK8mFEjQGlYXl+JSWxYD8IlHP9Zt4l
BiOu8d5hEJsuAA8FFb6fxjnVlPQbOdfYimEjwHqSMun4Q/cIK1cTRfAncNds
roYYK2DgC/dXyaKfrKZJY98wZ40G4ZFIT8Q0F+5/fGrDKo9zVeMV/rW6wWsz
fKJYbGxvlVC9e43cHHRHJFKYJe3Dv7ZDFe+8MkjqwdoDeoy6zZNuVnSrtSPD
/FVtDS1dv0haJtPTXmlHMqfhrwZjaKBqChGSScOhGTzV6865iLXr1ywKw2O2
NUuquilaPbG5BWdfOzpqujM2p88TclDcLbwQS7aJNj3mP0v4OVgi0DFp3Mv1
pqkWCQuSQ2PdMI5HzL6SPHzlYgccZaUO+2x0JwuqjzajNJJrGelZyLjnV5Zl
3HpNl56UIQ3052mQCiEEp2bbs2+zEYWyGqQAiijB/eKMwslh4BsDoCyc81b3
gE8WgVZ5d5MfWBpmsALik5hH/sfH5cD7JEEWYzlQE7ITyyby/9Wwlp+cYyJ5
46GykvedrOemVAjJM27UuKB0qO06nWgv8lX4bMms0H0Xy9xSwzK3ZyQAyRbH
DQmrzx2BgxQyOMnjOzeup3NFI9ymJBJ+TNjXT/9nGGiNlFZG80cCGy+E5dPL
l25SSdEPtyZMvW6gei3Rbb/oG8ucMBvWUKgbzAGZOfNqhRBQOrhxwoXNvNyX
S+LkXS8feR8iNVLC2RkeUw9XZPkftb/QZsXcl7EDZL0cdq8rS0pnSprNrXJc
CsrYBt+yJUGciZgdigu9NS6FyCG3HdJRJ/nL21AraFbcAph+WOIetmUIvboI
VIeeOy3Hw+iRGZoUzebr1MQISuUZPYOuwmCir3oBG4CsqyC46+pKNqppczm2
Dhzpd7ehXtJfFePYpAvH3S/uopiswPxt2G4aYSFMiaLP0uJWihHEQHYsnha6
bnlC0yF3KbzJXvWY8ynhAkuQVMc0wPOZbxIogj5eD7m0bS6KLNt9ZyP8u5J4
8ry4I0NFvpTchQgxtxGfoj6XU3TzMh67Tephz1+1GciPzvvBt0U9DKfJzlpK
rM0yeg3Kysi+5wWlNP0F5VXCAly+u9Ai5jJysUDbgHHBqv0ob0x3Ohnfagyk
CIyIjs2RcGGxT3Jvn6YoslIdGQRcu4zXjyg+yEBeRWgPfAoTwihQRmwOelOk
JhZS3MFdCmyqf53cYc48PuX1Vqy8IZc7v1kX+OQgyWT36rHg6d4MfepIGFc3
A9YVDZoGgyc7woSMMXEcutn3QvteyBbL4y5Rs4aHCVRkz5P85d+L3tgqggRk
ivSOIDkHJqlVesmtOu8XirCL5IZGPCKbBfT0jfYglBDZijMA+ohQWE60NDD/
vE9TAcdIAoqAZvCp2c/O87xjlLOuBCQSsKMw92PmA2xtb+xSmAzSt8eC0tpG
0SbeDaz4EuHHZNg+v+ZAiYS5XszKTYXGHg6lQiIIOpPAGroWX8cJXf5qZZ+u
6Y5+Usvmk2a1RQ9mC7ya2sVJ4xcmnv7OZKXcYpTp4cyMBRPSvOjZSALN7Oru
fJTGXNa2XPQVdxRYI6SPEX/f1QLmGhC444ApijqhD5nTS6nGD0759cNaojf2
hTC5xRaTzUqy9eNikIWYXg1c5R8b3Qx/jbTWOsAwcxXK2MMYUNC+zJAcCc0M
p5yKz3NEEzjKULQ/vQ26hQa55UNKD2bprsyjkP93jDwKbWDEyupFn6n4Jb+u
VzGKhMoqReWeuhiogVnl6MCHFm6oSY2R39BznNR5G7jdpMjR/aww8Y+V9I86
ato87xgI+qCUBTfooxfAQmxiOyrlsBtJYZUSblP5z4XgcEEyFVbx7U5nF3Y1
io1O8uFwr7q08SidBQ0oVNoh70bbfkCmB8iJfSxc+nNEcqTb6me0cSaTUUzC
UMirWGDYHDKzCpGk4dmngyaDbkdufSQcvSvKRFQPRXdzTNYlXtaGYhCQVJCN
X4oCwUIMzRosrTmzrEWAKFVfYk2zBPVM/4+iDkJj2g1YTIflCRJVmarPG2Up
xl7wwhOyNF83KoriYlQAsKxcjeL+bgYjL/5y4ZzzJkU9ktIp6/sHd2z1W1wO
KQ0xSWUQcXNSmoM2mTRpk2TzwmEJNfQS7u3ZwgcrMgAPwPElfyciWRFR1omg
LgUAfXW4wv3tCqPAfrnjVXF0L+FdERbIbWmegKsec17UykXqUQLApDcasevM
Dsumv7FRwIwFlT2meEt2yKOBkG4dkM3L/mpPO0Tf0VJHtJk+EV84M2rTiOK9
2oFEAeBPAEFnqTg08iX4SHOBUM1CNNmzNVzHPMRmM4ZVXZex40V87D0Z/ynm
IJoRBbOqS9OWdAmcqXdNr91HJvVmEFGMvaHDXSEghhuqN1JOG49LX+nDHYOF
CWFpY6xtP/aK8tuqIEWhsthZfAxMirAxQIOSeWHu3kYXVAes/zZE49pWHtLV
qLtmcY+rboM2pJYhpBKrjBSoxEC6QG7VXGFUO6RcOyP7VBjoa1STGAszcysS
9oRarqy67BICr6uiXWwf3n9e4+6Q3FRF0AXRwmxv4Ei5bWobXNfD2wEA7Soo
fWX0SUBtZbauAAUD8GqCKhjwPMZ/p8MX6Md0i8fTQJWHWtafSMGOhnY4bLYy
aIr/OvBQbbopqu9KRLoIg3Bztlt58dTLpTVBnNaom5Pto/5nLw5ymnFvQ5LN
im1UNZ48so8nJ+qkh1jjBe1zKCRyHICo5q2clKDXrCwLMqN3soeBWlx9XWAT
F+v0ij8aIkaomNk7ucSOmBXIJ9C8PksZbKU7/jd6eeRMIrpLKI3+WQUTI9JJ
rf9bw6+yt8juamNTBANgRejnyyQTnjQpw+eL2Fo8cQ2kPEfF1H+WBwtobZKa
vxWRxlKjA34GWl8HZWDciQ3V7TfpFQ6pa6MEXFIBgKEYOtWKd9PApuANdlyW
R4unwqyL7FooG+hYslIaC/O3yBfQfV+kgEQQaxo1DnyINsmyNWquO7bxxIap
FWNDNLQPHh8/CuX6e8zocVT6pKf+d32Z5RCqKi2bQ6WGcctjuKDRJjSEIXj3
NEBc6+ziHd238NdID7I9g6y0psM6H6zulX8cnJtGUdGCV65eaMP25BAnKJd3
3MUaoVoPOAPQGIXESkZXyolcP5zxHVod8i+aFy4hnIq7q6JeEG0lTbsDP5UA
MHGOB/uTcXqAtrm80KAOGSHcVCnFamEwZYQM1Nn1VxQOyEjrRfCkkwlAP/gz
glt+gAXXxvdR7xx/6o+Y3junWoZjnalSFV0rxtDDAnLXX3cnrH6oxS+Pk9Ww
RbHWm/xD9YIjTzuIVFxnvyAhO6eUO7d8HHFCl/r708CvO0n/8dxYvvmEYmaH
wXooU2kOvDJs4Ou24ZHxPiZ5St5TWpaWMfS12Hq4FV4rHyZVD+FI/BUqTkgt
2frl3teBD4b1EnP1Pa+G/oeZLBYUHY6oTozQdE3naMDocPGi8C/JAq0VLDxK
RFecLxwCm9fzE/QK9Os6T4/65/1rcGnubjrcg8okdj/EgJlRQ1NXJs/9hsqc
FCsINbx7SnBEY5qOalGTXAXbb/0+pGPBFB0rmhHiVBWiJHnWL04ijjj+HzTI
PRjB0jBeiyXs08ytqhfx7r+KgRD7W9itE42e56FeETfTeyMqrYJ9ZKVrB63F
9hTay+GAGkhgEvJsPrieUYtPdmtDhz5mtMBIUPRifTfNe9J/frJWf7Ir+yEr
tw2PXo/Npcg4N8aIiGpw11yTOOqMefeI1ng7DguFBnvjhlWgLbIA3GTclw04
WwYrEMMCU9m7gZrghqpPD4OEow5ms2OiOALSKZcUPeAB2BZUzyHIGoUJLEys
EJiSvS14Ih8vjLejrlHK8KsQSmN/cBliGbcUv/8RZ2JSo6503R0cmyId/1Hh
1fK1KXom2zsnnBsiUj3xPcnWRr6DrxHv1zjx7MEFJfsiN1vHm+rybqwWiZH1
aT4ij+QxzTjE6XC0tg41qBNfd1VsYNjawCP0+f9zYcA5gtDrPasV7ueiXLJA
TOuINl5PYF/TkCxK2s2+Al4Q3AUyu2na8iVLRATaf/NsHtIZ55GeWCu3AWjQ
i9OkWk3ND6A1qplFIVRaz3WU+hjxX4DSTEFRCLpzjPD+QCT1t1aCBfNyFUcS
gxlXqcM1dnoegGAoy+fx3BuAyfot/FOKYKjQ9fY6bRblilHgAG1I0eODNASn
ioifpN955boaXSse1okSLC13ZH/F59ftcwKMF4qZLZGPNbHPxPQPMh3g2bgX
9cGx0bzypaaXyWuNqaNpfO4IRNQpbkBuko9syeO6pbTKS2BB67HbJ8kSi3Fh
VLmRSM5wpZs+E7N2K6OI3xZWjwC2WFRLAFU5Y6sV/4c5tgPHehKNX8mNpvuw
x28GWP5Ts7q2txQ6S7VUjEVWjufoBgu4KUEaZfAEahanS8k5lAXm+SQVZgSU
DIuO4nF1j6wZBKmukwG9nSiPBzvouLxFyAlutytRoZUkL6qxg6wWiBgvNGOG
wseCYTzSbZe1yNCe+qABct9+lB7EVV5aNBwURnRsff+FgIipPqyEff45hLE+
VQc+522T6oaTjTHIR7KeF7ll+eCSoFnQ6PBqj+5sxG+L9ms9pQQG19N58ojf
0OGhoxPcZI5iv22EezKC2ZKqoVqwQR07R7q8kwGmYdN4XkQ6wd0nJ2I3Fsdd
iDuVqPW35F1MizUNed/kfYDjn4BHHQN5XKfJ8DFDgWHepNF96fjHglxRYhbH
d5qFMYOn3iyDUWu2B5Z8TmBebzEM08n3i73PYa7M+8yzxrgXUbk759Zf6EwX
KHKYgomZ2/ZL5CuiK60m47k35MR9FTt2VDfXIXTVUBM20pACfU6ACWWcMWG9
FS64PLpE27t2xVsTUICcxWz/cT72X/DxyZTjrp1rHSQGrZKhTdD/KzvZQTu2
Fqoi8GfQgmmYmakUys+KKBMgiyKrLsdpnZkTvbyM9Gg1vRgEZ3SgEPDRJEgi
gYUQ+IikBfgg3jc0ldOCS2dz2xdh0aE73vtyZ6AxxGplrvt+ntvGuG5NVqNe
DxRGk2MLjqGzMStkOC6lNCIRPfvXwDf2YjCgQLO75ZwwNfSlGi/e4FPc4tFQ
oXabkDh7AVNACobt51Q/xQiqstGAAvyN9kIUcEYDxZ3aZA5+p3DmMSPdBui6
zI4lGY6yYmr4HkHW5KG9Sk1B2nrTgG4XhxpY/9hqqR4iu4RmEJDagvXrNB3P
vAV9zCWZbtvyKYGy4LQLjhgZVmHL3EIEwtjW2yCgnAthFdUSWmAtFyDnHYQK
944FSDQ6G4uG1kmwRKwkR+yA+4Ft9I8T/2/Zk5mAK2AXmZqwAFZw91K/dw27
SnNzUISY3LCrHBwzBau6AkySsdGy5nWrbzT/35dwZRy38V6OTTHaDz+8YPyS
dgybQ0Jw9hPd0KMUc+c0RtvOJ+sqPmXgsWG8FnnRcp7U3hZTCeuzFdjMsi96
oHHF74npEznq/T19U8P8H2MZl26BE2lR+27u6u/0KALD55AAlAJf1ykh3F7I
Gjy6J0RCLLhfarKSo4OqJstHTpgA9jnOzvUPaLfveJrTmkFza62QdILs7K0U
jlDVHP1UapnrpxlXweIGG0YaDFr3H4phrXTRjTtcToO4veSbre5j3TKKRal1
bWgIAHfn5+c3BjifU6YT+dMuTpAli/c7WLHL3mAGM6vnPMa2TzeTIY0YIIZ3
h9TBYf3tKSWipsQatzZQAqe0BMG9CZaxL+7Gyi05PKpWkY05FvnTR69bo86Y
+F5+8unsQuOxk+cQ32Jm119y32oXCkU+boyShTIsEWWmcLkRpMbvKyHPCIa3
o9QSBLfcjBbmJ3iUfSuBFOmm28btAlOovO1UC648Zc2aYJfzI+bpwlv3KyoZ
jqPwLaQVesrV/CdgICOPCtRPzXPBa2kxajyNTqXX8wZp87ROK2KU2Io7WYO7
J/iTAZJrkOzBhSfCodBd9fPj0n0VV01LQYsSzixZ3Cg0SiLB2SIS8Rhoh+qj
QWq0M1jIcxY3g2LILdb7lGM09K3C5IyOpiWCsDN44OSOBkClRM7hl9mThR0U
Hhx9JbpQ2mRY12Gcz/lDiydfNly6qHbF0bU4Vwx5fOnieyY9tqeKXh7T9hZ+
dSdq9FZOP25v63k4YF4akMkaZgE95rLmmwfnE6Ip+9EgklT9j4yM6hytDCjG
M8I3Zc9SqzrrbFojV/sE3pkEgfGq4W6M/nhs6AdfeiQGyG4otYdqrFHr7oIn
bW/QbFEc9QSYLCQtkYS6EVTZ9WUpiCungKCmi4NtRwqytY2D5ttIUQJGlLF1
Ng0FjBjCC8do52EjvYn3y2yw/CHEen5BTbNKRoqTTJ/xXaWK3ESp8W9A9AwL
p+QD4xZN6YR3HbI1EJxdt1KXK8NyRzTqBlGVxOnRK8x4YvuJnJoB0N9OczAq
K+oc8QSa+dE3dGvW0BY+1KzbDt9yzQCjP6BVl90OwurlxB2IHOoJ5AzjljVn
/E03vBtNeB6biv6Rz/caWa+fVUJmv+kCVWgqb/KNJMDkBljht6lE7wNHWhSp
FBnHB8vCGoNuYw6Zm+7B/4NxNuzDjjRyA1447wcFanJrdq/N7/6bCvsyrmIr
quz6kJMTfzUiTjpaybOVZsGivd2yQ88oZvd7AvLybhhiwDn2P2/creDSj/jO
omLP4BET4+Sz0kY70BRX2fpCAN8ikEddqbPDKeh6466qRx6e100yThUbwPSL
UvI9fcI1uI+08gVwWpEjPyLsvqn4Hs+z+ahll1lWd5jzY3QhgUhOd+ily/Kr
tTCm/nF5mE9NWKdK6yPySSXA133ugj8gkV7vVcTq2zUp2JsUJxDSzt06RZ3D
YE2yKwMqSztG8n0S0RPjJIUvs1rQIA5HzyGMR7ZvNTxme92xAAeECxeqDJws
akdRLTZUk7UzCYvbXdAm1Nmow9UUZlUDJ2E/6oC099uboWM+93R4hsAP7IJ6
GLsazKMu7kYdEKJwvOlHYE+6aCGdK8lLdZAevtqrS7ikiQX5HcYPuf9lmUyN
dLRHYWNlAx/5DNIyFB7CtuDJh35SWJVq6wG4oiWp6eu4lTZaE2y43wabUrsg
XEOBB4UvmyZhZG193FSdk5xTgC0be/nmGoh9pk8VBnMkrEMcCCMfj9pxW8oy
7Dg2KuOF//kx5BkPi3Uabj6vWcbNyIULKrRtsxHV0WY3uhHBv2QVM1Y5bwN3
GCfGTTwdjW5KahvXDVJ03PsPZv4Ws4N9mD8akgPlxl3Xt7zNC78Nf7uPnaYk
AxeEqXnFuD573pUFcZnRyS4qrHt8ekgRwuJihzO/n8Gmkbm4yJKQsm2awicj
DrUNlkK7GYDeDpajxpCSpf0LEV7eGO0tLy14EvYhXGP+t6DQkWKNzaoh0XZL
5y+enP4YUtTkAQmjdE3rXdYA0jB9QIwbS2VsxDGiLemdHRgw9W3QkXI976tG
e1vtJrRlPS7bcxVj05gSWd5dOfht8xHI9IFIgCB8/OikoWCmbMpl6u2XhyOi
MNYAELWdLxtXg26fFeN0tHgVKLRNI0Bu+Ha1kLuBZns7/bX0aPNWcKaFTaVq
yeiyRmBGxqc1RzjxQJM1z6GV/r1HNZyrQikusi6ac9QEQxNgu5hFABDj6NJv
j+wXIIX/cWCjl95D0ALV7TkI6OIoeukV0GTId076E+njVCAT06iDonCUEY5O
X1Vhfa6i3yb0R9mURSRTDf7O1q1dy3KVG2RXEaxaojd40rwjtKljRGIyYo0N
wzvNOlFm1tHeoxfdkw9dymLB6NXvCupeGVin1SqXSzDiDPfpb+shtbjCXNas
JntoAqLkngaF3mjFh8vB6Rs6rwjuGY98wMghsBS5tghpwreu023vt2kZFHla
uOtJL99ck1ChB4shRT1WavZa0nfsWDEpDesYTn2RqyMgL6mT2gmDToxKGeLn
hh+X37fnM3FHUUhiALBMhaS9H1NpKssT8Iq4DiuJ5vi+kk1vTikiBKqRlzrD
RQglf9qCKD0z9iwyLyJlfISH96+zwmwQgxH8pqxKI/0bBg9xT8VRXUWhRSFj
1xKr6nQMRY2lkTisgPaasOL3DJaGVh1JyqsilfhMzLiGK6OwwgO/nbGXFF9o
zUcna+6oRgAJhHjm2ZaT6UZ4oIEUq0/nnm6J9DNq9HXzx2yeO3+vLlQ2gYf4
Ny/uiqHWK77XQ0/jw4xnwewQl6LsiwLO5OPvP5UuqNYhenyCpyyfgaUqRedU
aqBKfZSKtksYAqKpKKGGStGQQz5rR68IxrXl+gBtXJAy4jBTudo8Vp9nRzUj
4wyQPfLc1r4xoQBTCccRBSRlouQnWTvWt2ecyhSwRbz/RJlr7ioOfzn2fuNr
5wL7tFQrBe140KhmURE2T/Xbw9kuvnzK+hMgVzl4+j0ybjtI5a09HP/cQS/K
aaCqxVeuLZ2L/os+vtT1TrNH8aksPipie6v0kA9OszZDEAt9lc6340STWlil
HfeaupMtGX7lOaqnQ+MbgyOUN0NzKEs6ebhk5Bfp/n7SCYbEgz96ZUS30SJH
5IebZrvkT6vYA7JLcMTb7Vea2MSuLcz0dVgxEmG/Ar0NBvqLer5r3um2SDoS
cU1zny4XvS6/n2aeObg8WVkPs5XNu9WdaKdX2HJxzj6++99LJHw356W7RmOy
0kSntUwz3pRrGcfa/vBO0PwiHnMybBHOND4Ctc4Z0QL7ThwTMLDTyLFm7mlO
BpllmB2CBMKSxIqzhqK1XolEoUE7QMwEFRtYAu7+j5AXBCo71Q977oicBypo
NHxKdvArTZ+CaL9nEmZMtaciDy8nWG7+zMZL7uCfj/tLarYm7EXrX/RYgqoP
KaR2zBEVHxJ4RzmaWOPfLAiG9zVp4nzqMcD/yfdWAE2wLpWEP7oc28+xuqPw
VHYgJwYHeCimrc1wEmg5GbZiaziYFJw/6eRGe6Zi8TxLCZHRp6EdE4EIGI4L
j/o3nJcm1YnApTy2f0IXSv7RUWMcLcx8Y5N3+kb/9OActWKVhZf63eU/aYOy
3/ToThbUyOxuupRzSR//FOejJ4ISJUwMKts+dpZjHp3+W4Kxp6HEVw46m+/X
xYLjlpcnOA6DlWljvI3Wi5vl8ahuy4D7k/+E+hKnCoSHPwFbiWBQzXLTb8K6
IZ0B9NEe3uKXLy6I+9bj/zk85xPFQr8xjvuYNv2GBe2RS3toU3SkxO1zFopZ
fZb/UfgmSe19bS/bFbFl0z2H+Om9K6TbpQyI3qz8MAp6oglICkAlIIxEB0Rv
j3P1gtJcn95SpySTBCgjOcIVUwoeUvn31BpQd606lQgAEGk56Rbe2Jcraekm
exg7VGXEX77Z82q5nhyChNzlHUrMs60DZsINyTkO0XVR2iTt5q0FwZ0uAJJ3
6ay47Q/3rLUJsQpSLRuCPWR9a0AdGelD8dbIihQIAli+q+egs7vBNNmXYaPc
TCVRNpFzT6pKkWmLQLQ0IU1WJgPmsSbhWsvk+oC1ROuz9R1FEEkU9xMb4aOk
wEzr5j4JD0t8C6QS3esWTx6ZQCyjIw2wwz99AGX2QZUKT7hO5z8mJXNQlTWY
cFjGD8qpPPJoBaKh71wFMNSZm8tjYETw1UbRMHDHNjEd+qjOgt6McvGWJhEe
D/4ilFzH0SwMD2GnL+arvA/qN9ttfUNiaxD1vJuu+gDS+5QxPmCDn1QbnXaR
k7q6O/oyeHxfpsF304GpeE+cNQH4ekQ6Fw2CUoleUMBUHnSfVFO4emLXb4kg
L7ByG8L5nAtekf95R5u9OBzqszfxlomUhlfFezSLI1/E7jqmuTFW/5v/2iVh
c6arhcEn2qsNmJiK9I8PJUM1RbHzmCKT4yNFbCYT1g8QONvPwavv/lZLk5GK
VpaQMHsXVpldHZj6fQ5P5hS278tv+OVhEMKeNxhI1tgkLOixCzV9pv5YAAgw
8F/fuCjTgJUOw0sR1KKqD8pQ+gMi0UHieb+iF/Tbv5vepLcwXEDJ04icsCxa
vVSFNqJ4hu1DX8KXRYt3JYjB4bn5wZ7aKA6KfXdSCDaflMIdAhzGZyg6v0eb
udO1XcrFosD3q6/VEMboHdPLHwEtnZQJ1RpzQmONd/46EVAha/pHh3nymm34
feiQjlbhr00S8A52HWhRTqVUDPWSzE18gVb0jFye3hZ8HKen4naYRibVSPSU
6jnVa4Lky9k2OMh7w6rPxArbSTbxYHwMvJoePbkIR9L/LYuJ9bniFh1RFKnz
kiprIyofO4Jt7EQITJh0KrBivh636k9K3WyZgidlxz/Drn2SBB6GH9nSgLOM
2h642GvTGXS/PQFBKCZ0BCc5nVNZLUGdwY4+IJBZwIaHM734Vq9+lbmGxHmq
etQjMmSLfFlhJwz9Xi5M0TeNE2lg7NTOfRzJ+bVFWahxF071lXM6busL7Mw7
xlOwd4zCJCQnIbODOn0qEUZsblz+84QURBYOrKMjSVKYNBlO7ApTkpHc23WU
SYoT6aVHSJJlFvMxUX+X/s0zsuMFBRKfxie4mAQpzeKim821P795J58FOE8F
KPW8dND6OaZ6Rfm8a8fo5PKhUpkcKuVsXr+95mCfZeATE9Wi0bvCT/DJJ1x7
vWxhdGP+pEPmMChZja2v+Z0h0IddVQWTCjsam0FRadEQt432q1ou3ym8esWy
1HE7obYTlSxtQ2tbN8ntPU/MqRSwbtwGCzLIE9xsMGgpA2oK4zEyYrp+adv5
2UZtU8KLhjgf3nrwvuMN9VAtYk5lQ3aDPpgOtVcn4hjboSqyOYjPFI+/55IQ
nYyA3SiWH1HShRmMaPeOqzp90PB1FCdus7ERqerAssCdyn2crp67p0jnCsQI
VOFaKd+CUV4ZloWxhtCuUvNvBaodPosg5X+edFbVIlKLVpf8g7GYoLWGzKFa
0MaD1hcV+EThVqtdzC3aSyRKf92CHe7EB3kzBBwpRPmZcGKQDI/JD5L1AITy
GyyO86WiVPfjiddixZTpZBcNfE4D2zPauKss5Pz+bz2d2Yn1tbqDpdlrfmpa
Py/vLwl9HRrbNf6Ex3zMeKPOAzIQzDJ/3pku92ihcqKyfHXhdSOswhpou6QO
S+EAlj0FX0adfPXTVivQOwdtv/2mYfw0ANmHQNNkAOWmLFqctB2Amrd6hstW
pSS0SRPKYo4HXIfIndFUUsM3Zvc6iFtdhHVkrN1/ciow2gln6jGNC7N4h7Tc
VHS8xb5z1BmmwBB2UPQ0qWncWgm4n2lcSiwBFtBGYZbXWUE6nzJDOFhx0G+/
RnbwysEw5k2p0xhHcGRoPbnisZNR9Uaawygte/YslJjYk7xDyi4TTNIsoGE3
sR4SfZDuq+Dtla5VtpwbzcEN6o27I+9Wm/DSF5et7JqoKS4KqQrdnuCeyXL8
vuGKjNH4n2AAPccttMzZBT7nHh+7SGAOhsOf7h+ISFc0UT77Pvl/fK7aa3A4
dxueGAd6/jRrPwLez2GkIP2/NltYudXuEPa2pV5XwQ2PoVyh2pFj6HdBrF+P
1vOv6/rbRIJMfctb/KS6xlsO5QNrJU0034xhv2FKOriT1rmFSV8LbHtwRHHq
vL/Uz2xNYg01OrduZhdaPwCbcFBBl1r9JLc1BimS6j8t3E+gezADgFjiXTU9
/pRuvxS3wQvv8BkeCZROvEVYjrHmg1R41aNUInlCElaXNXx4TMpjykHuXIgJ
oSba0gGYB3/uS52fixL8OTlRITqsdv7Ty27rG/I5On2YpEVYrv++nfILGSzm
Izk1uUPzjstV3px14pg0PJCBycMvfAQLRBUuuHijOHIbcCqBnlWbTchHkHXi
Fn9ZPnuXvB+4VlMTe9qaZkPstn4piBWw2vlstdC/f9adteoehob9H8ZKeMRk
WHtpBWwuuYnqNNkxjC093OCZUjdxSgteJeY+pPyejCJa9ImJYq9LxyKq5yEu
k7VQSP43D35tHMCXPLXtPrdRYgRC2hZr6pG7D60LkLxhTr+Lx921FOn1kYqR
oP00f/Rte5ZTsFYa7RUrWPKsQmQKCW/u4XMidEHYn0FaZWxc7Fy+K+4JZZef
fQT+y7onRjQRKe1D1zo4gRwLKThJFnMHf1OtFPploq6XS27yRFd4uF5WUnsP
4IfVD1TLu+4FV4LSzlCld94g2edeNs4HfItVyYOWsECPwIACV8bGYUWf9Nxb
Z9qhPRZITxHvFCuLh5dVuhj5wvZO1Dd/MLeknhSzutFktB0vgxOnwFTyu8D9
UuX/EATZwxHLpmKYX4HnGuXSnOGrdkWyZLv9W7Q/SHr4w85BsQ7PZpsvXAUK
yLlMeilPOq1Nlx7THmg7s792ehOb5cSzZ8Rri9lJ7YQBzboHFw1CzFaX6ddL
jLk2iz5Fn7NWejt69Zkr0xHeVXgCMmy8f8P7bnlsNWjqgv++ClTqsz+KlXKt
0cQ8mc54hlaia5B5KB5u5UtHndDc4eG0IStju3hSNNsz121Ac5nljS1lpIUA
/cpt9Pw3lzG7aEmRuEoFgZN31EUD5Szya0Fgxh7dBI/hG+9KhtYGLWIHfxDN
rQjr90DC8lSj+EJ3MEe0RRMh+TMpPi+2KjTkMUSA5NmefSi+TOLLcx9Fgoh5
1Rv+mY34uqXv7Ki9xDThbePboOYG8SSOf27ouycBqepDfZ6ZVWTYeGTFq1pG
Wg71FjlKp793Pr3DVZgUvUFfE9Eho1YdY+GTUV5k/8agreyrGdlXY0US/ziV
PzMy9d5hEjmaHgLeDwOqsw2OQpdEVqJaELXJ5v8bA4JlrNv/URGPW9TCsAOT
n/ZAuLBDsZ5hFPm6+gaSvBXJdZbPebMIzr7WJMg5Wu7LQZILze4+NioYGQO0
GwZx+UEuQj2bFfrAZ+ctFmqp9p2RMrdibacxD9fOShoTbFp3agZf4MlURbov
oQqlXWKmWKG2kL12P0ooMTZsHbBA0cDafZGu4ugyd+7K2mTkIxK9T1X9W+Hi
hQuPK3ykHPvzic25MOQqpeR0YBaTJKiIOQPTIbkjtW+Lwcr3cWwJT1BeVAPF
ZlyRJCAoe4xVAAQQWwwcmGf6C/nppyYS88hVN48IzlrzA8zCAtOWJMUV28HE
BSoRT2ZwTntEdUXS8KXuoLskRZeRlk8vVgCKu0Jh84TY3MjF34xBontHcKOS
dk6qefIwZgy0jXq7/p/lVWW1J1Inqjb6SZNKf8fxFNwJTOJlB/i9foTjMrEh
UbgsD8n0jfzZ67ud6fdUH0AKSdblWDkbS3XreiTHQs+OjZmNB/863kr/Rzcg
GBvr9XzAoHI1FF8z6VwlLvs2seYQ617rCch1AyRzE9J40eR9Tn8KUNkczvmu
R+ZNF2T2dlXCGNWiC+b60UkE30Q8/au+utKu/Lpry7JxWUF5Rcz4ZVj1NLEV
5/Wga7ji3dZ55LpibUbflyyrHucRkxz1B2lXnXgRfI0W0HQQvoEWwSrw5OK0
g0S+E/3NwLCuOwCDh2IhdavsYAyVQz0S3qLRQye5u0qARfWOewzXhG2ZkPvg
K5/NQMekW0zZkZ6UD8pnn1cqBowuI8PpO4wV5pjzcSb8J2rr8JfUBqgeVy+Y
Q8kSJGmJpthonZD+zV5JY5A+RD6myOEqWmR+w3J/H9wVn0y4FiLCB4sQVi+g
cFuJv1hSb/IbUov7AR5x0E+hVO6xPjA4ong5LOIXyUQAsNARkrLYq20ruPgJ
yiNIcuAO0mEm8Gc7jYxesNHrcbsI4HF+j+Hh0AodUhcCq19VHsygf0xlgYJ/
+Rvr+X9qZg7n8n2bX6x1mBl2ruCvST8r1mRVTy5ym/wDF8yTcyiGt1AD0GLY
CccGPh+kt0RsBBTkh9Siw6fyOZv6NC1zDr1xEUDS9QYcADHPnY8RNuk2mOJL
uItWHOSc78O9A2vnJAzbOu2+NmDz18ZZuETA9vrF/zxYonx3Dca3hfj8TgfU
hsBjHPSKj0Po4f7lBba4KcrRKmqgQSbhGWpaUaU07n/28VKeS0ZUf5dVp5xK
S2c0iwDQBRQbRx+CfCslfewknsW+aHfpyT+Sf2EJERGbwh9NMZolvX3N1rSV
GuPPRgyaHXmTyxZD/E/oeAZV8jxX1atwW9GDQRYVu49OgdMR0S12o5TnhNef
hxWeVREZr4uTucYmqSfZpRLaTcuiWnAvzOZQzybIouGpczUVSeZ4qp8DUYGf
IrvMMuYgPdQHZyW83GZj+LGOgHa5YBquV5Xi960QYzOG0YZqRqDre6jcYnLF
veCGPohNOSgUkPsX/07LsqenkbttAFdezAwSro5T3IC2iBa6YWxzM7CamqE7
uFsLEg+I5sXJ+yzUOYTAZ1825bjKOO03br2B12l+y36fiSEckoacgukd5hUq
3HlLhOyiEctlNRGAy/lxQGz9ujBNUUR0WFcVEZjUncpqB7hMcG5BN9dVIG4t
s3ZHt8p3it7SPfOCWeQMz/3QGVR1qMdKDXjMO+UZ0mir+i+D9S8g5uKGN8l3
Rb9IdbmBdWYubXQ47livm+iRzyd+8IXLWwRKpXbOWDKk3+nwXzDMtu8BR+BJ
x9CKh4Jccd5VtLGX7lVBGyPHzPrjjwVilujgjRTGmNR0iu3QJ5uTJv7XI1yO
w5GAMHMLlXh0ig7dzdpzPDjQe4UvPjz1fsgkwG/SJfM3nvFBsi2YJG7Z7e+M
3bFXSoJuZcXPQVGLkEBXXLlATyqQjJSfB4qYLQBGI5UXLbVDrKZAAy6d9Ueo
fMXeOUPADDbTBAntW56icoTSKRgnvnI/tHCOV566kOySdo3jtijsYMY6re9j
CgxCqbvvozSnDAB03N8ei7yCLclJK5dGi0dwEfY4hIeEF282T9rnfd0q2omm
JK4war8Q0x1X0MjmKLRoj/ZTxiy41hN5bZK53uGC+8aTBgB06/+R1Wz9hyvy
Prft4HDSEBDlLyNx6fIrsaDluadQl6PUQmTN0eGszHiPqGaoKJxuR04QAj+H
qhTKzACbdWlduRRw72pI3flxtEMbpgU1bM0kUzEhizTh5ufQzz5snecjY9HI
5xJAZLivs3ZHbVfnhkBqH1CK56GiYCF2iHT0V0SAvxMGneJ2hZhuYJCrRlKW
CNI37QVUBVjcjwUNPsOy62pYf7icLezbCdkjtUsJS9PuxGydtjZaeislmUDD
/T/fYVRQyR0ZZVIiz9CN7sBZ34oV9W3OOU38ZQTaJg6NOV/KRlzZpIJ8mrlM
SqzvRLJ7qS9E/Jy+FzGMaSsYrd56QPsGpjQfl/5ts1zcJWNuYZ3OpkYwlRJG
payJ0EItbpiGb++LpUa2Z2RHITWzJHiLBsznYXM5JEdQZW7/yItmjKVij3YZ
WS5MKVvaXwaVPX6iUQtjhrIDmCyE7QdXl5E8nEFk45WFmc5x7BrR8oemeCdn
508QzUNOd+Ldviibxnp63uVjrbaWqUt76JJVv9kQfgaRyC9kAPf/TXt24Fri
5+uQFlJoEG85vu306tTzQi/olAUu1hz9tBqPuSka3Ddm4ZbJ01OvPmTxb+iF
sF6crm8myz0NYIuCBkCVl8O6ctQelKJRwYzVH87tN4AjGYFXLSCbrHfldx8F
qIgkPOOJnaZi5DwfElxSt8vS402sdeFJYWsVwqxahDnb4r0uYagKWt9B0hqA
HNDmQ993hXUEuKBnMiS3Z/daAOsDVA8uCx8VsMcwz/BxNtjHPL1BK50Og3kQ
eztLsf2pZSzBBLjmxd9xVpgn+KrueWg+R3s7daJwvTDwJfEBqbTpBOubGQsQ
IcFJbAYhioHIPR/FPLHUpeTiLaeHuS6cqwDp20BNpbu5QUPe+9nhoE262cOC
7u0rIxUCXuCK5VnxHz+S56nkTYlCvImPjoq8ttj0BDpG9Df4QKAcKteA6sKX
dVfCU/ussjVxfVsrevq59vjCn8Hk4V8Z5Uv35gLDC3ts2DJ5qm+VtJrNYHJH
Y5mbWFPqk3PHJz/+6Y0CehLmWHxS3pggux7oEj6fr9D0eXU09SQfdiRhvCdI
yPFR/2JIdaPJ02qdF54CijuKDDO1+HvzYccJUbJz+5FLCz/PDmRMsBe+Z9XT
5aKgKczh4Pg+CeFm1WH1BeAh8f244AjCtMU1DPU3gWN9fyzK6kwmf+5MDEaK
1wguBvcZd0TPyPnx0sFvNBMrMUBVovxL5h72d4YamLtYWAtkUmtC0N0RXejK
0KwSFLgzHNXFthNDopBKYo7g7Yv9F4xDslSR7dfYo3gkYT8pKcM168VPMaz3
hS8brZ7FblgQLqou0j+iYUHibiY/Q8Pk2MZO7krTlh2/zoVMG62xWXZfnnUj
P5z4mPWgDrwkWWkX0mhGoz1X6T6+hOGLm2DxtPPPBJKsP2bQI10JonnvsMG5
Bb0eyEnkEb2UuInjQApp5pkwG1XGKMEYNzwwCoxhSi1x2WQda5WmfONVWIg1
VkgKc+ar6fsyLpF+sNR4aYW4zY2uT3gDRyK0ZSTbUF35uafFibd25eMvS3xb
0nNPtEWHxwgnw5ha83K7QD6M278bs1Fmpz02xwPpoSQor8TzaYjW9UjDrQ7+
C3bSXSOmzW5/JCNnCus6rIOlIPV6hTYI1xncwV0uhB8fEiERPaiPM+4XG5Yb
spPhjDzGibd52lM0SSkqeVN1ws3rpb1oQZ/9g2h8iwM3Y/Mx6W9tJ9zbmo91
s0t/wcix81K9jFbXxx2VuqCZdSjdycKYJWW0LCt3LEr+EuDpsQckEHzHxcKj
RjA+00u6xyNWgFdPk0DwBsbv+ZpwXgEVMFB3+p6FqWXp1ZP7lp+wwfIN3P1c
RL039QiqwhZHsYQOC3kN4dcpw4KI8dD2BpDyDxVJ/nB1CYY3jSi5z+VW1bXE
HtQfy2sMFYzDzF9aOXG8FKup9lSGhe1f5CZf5TEnfju0X+54eI3Ys0OUYP7g
BjlqTvcYyq7Xa78rNLCAzke8iVkW7zTuZ8jGp0/jTyVDC824fXhnjPBrlEp9
sLxrRndjEfzvQdT0W5ve6WPZqEPA1QWMQf8QZVM38DcBJZnGYs0kYE5ZVcJq
aYJT8lw3/m6L0DAaHEii44IZOiY/dfpTtRvxKIyOhOibLQkHF7lJFYMehkFn
MEawh7WViJ9F2a6vWD7yU6lOKmXfmLsBQJ5hPFasPB5BWFpdqmlwrZ7TypWX
7NOW8aBZLjkj1+ueT1GbU93LKnxFzQZyKT4KxxnbLeLY4t4fcbYsAaim+EFw
UQS9fEXhBBc3OBA1aPGwY7vQzt+qoaJrAjRc/xDlIYq+IBNYk/MMEMOLnMqh
TwIyu4w7zUq21Is6crBdE/mdK30C6Wyu3duJxM69URUFPvWJiRQMqDsFhNCu
tvm7dY5QCf5dlImYVzxGQzsj+yv7RFBj/uFB2Ea+MVzXeckPXorkMaBMXofz
MRm8C9svzqlAIcmv43AjdLuE0Qt5jveyolG9RXWviPlgPVBBB4lK5+Lt51rY
brN0kFDdFoOQa/ho945tChWvu1EoOARdmT5rdJ/MoVSR7rbxBu/uvbo/AOLy
FsDtX5EQKInLgqwzUxl+lqUaA5ksk7qANclW4vTexk/WA9H4Cvs0AIeOL9u0
hK1BWuYQQ7o281Qre+in3+OZngCqLaWwgS2XG/ShlNdKzC+skVl6FKhrA4Ex
G3FEAlj7FwBDKCWkbKLsSRcvkcLQQ7H8JvAsjuhjd0HK1HGQFj+9meXwR+rS
teOnHOsrhbviY27UmAcSpyVGgFZRI/s7/Fy8VTDp0TwkzYpay5pCbKubXLkU
chdTPKukV5O5pIqEvoOLg1lTuPi25ftcjsCUeUnlMcv/yGoScpi0rLbh6TGG
XlykmXeUF44EOk3sNKJKVQKb8azH8+ncfpyM2zrs/Vy8iI5iKIdjvDvs9xUb
DOrxqlfBj7A7dsBnykA5mxJ0tDbZ0Dp0zqKpkcWwprnx46f8jeA0gtXr/5bz
9CmAS2AYG3zb2I0gnkntOQj/tAbVIdpp+gm2DwEpVJiMfIfiDyEK+1SXP1c8
AEY6coevWmjej06sn35k+ZLJ2TnPB2Gdx+XsLWCNgptTgfsB91IQYiqgN5az
GuHvhVfGM31UVG0aWD83biZB1nArrMVkGMsPyNG+0HEtuLeAowuxazfq39vw
rCLsmQC/zXQa1s0um2PSjMdVV8Dvlmhf2Q2MibOX5XY32DYf7FvswVKJQ+Nb
QeMQFJRnKAMaHUG9wfKreWjnvMMJ5RLI7zo2Vv+eX3HEKpGbR19NXlzHVVyb
vI/2zIXRCX+5Kby8yXrUHOUKkXXcyceX9IZW5+GhTHF38ojrDLziP9Ty7k/N
IDXX05KY+xi46YOGGRqJd0+xT4sU2sXj5FgbxPGBQIwP3MNy6+btuEVeFEH1
Kqo6DtJa7nPojOmiuL6UhEAmrzCSxxhgIQtsexKm2FJe9ir8e6Ss0xDxK7Hn
XBaZi+lf6fWdd3isNOQc4kwn8575Nwqz2X+CH28V6DfRMUdahDRypQ9wV72I
69aZk55OsNvo5Kx2MyvCMOlemdiJ+/Balik5t3ZB7LrNDuNNmXDm7lukVSTb
y/62MUhspZsjXUei2X8BdhwnNiNhDDeSVWIHBHMCtyl/gzELD10QsiZqs/HX
J6vwMjdkLZjo+NfkqSt3a3dCju6BFzmbqiwIa7Lp40pgBZrn8l/ofT0yCwdo
ks7yA6s7j3e/Z3eVtcbOIOWWhq9mzKEOVRV45/cej18EeroX3zAfPTRnDQDr
XWhX0aQYgs7XapEvRY1UU8RiyUCHpHvQ/wiDC8HNKQBlxS/KqYPWQ/Ys/PPh
jHF+qP74mA+7zp590YX1aNrr8nsU2h9B8Cxr7xrjQk1RCb39PZ3cs1ns6bgH
E26CFACMJXMQvoGv2K+Sy1eUcwDK4v/oGv2xIKluIavkxYH00QyUHti3gHPx
7/zSUuMPB0WRUnUrAd5cFCVFt+kjMf7UkLBjhBItHbakNIMeAMVyDTS8h9ph
clUZjleP+2UypUWSoRq7h6VWy7/HAuWeVPQiJRdaCSv/5y2rfz0gPqaJFe/s
RxNrT5I9p10BcfbTWb7tZVn7Svu3RvyfZAD41HeF28aI9F0JYMTk+X6nvIWv
/2Lwxqj/chrLta6eRtvhosriTeJ+ya70eS9Lf/EABiDeCw6tcxSQNE6NZuCO
bIbgEq63V2IRHOzkSWOJXOv+NEGYHvmJqoKreaN/pNagKX9Mt20RNTrLA6Ln
FtoDuy4CBEBhXQUFuwSrUjJ3uDUfczkeUNYQpDnWaV9eVyQyMPSvYkJuD6y2
9tqwP7Xh+iDm1u7d31gH20elG7GXRKjizBT0t1SoayjJOtfi3gCYuPrGJiqk
1ffsroX3ixwOISYFzWmG+1/0fupKwp96S/B9mdjkrZvv+zJ12gMFyRwmOrzB
pHEJeRD1ezxGZjCe/zXmuI+Uqv+SiPvkGsU9575iNPq7iPl77iJorbEz78BY
yCcLiUkJLmJInNfiFBORO1q9Dc9z/2ZoyOdGXCRcCoqUYgPfzwRVOMdG2YKJ
WIfjHsqM0j8EuQ5+EqgH9byswilzsncu9dMyO7uQnPt7p10c7SZSmjZCu9k3
IDb9D9bM9++Qfsu7+CBI6MwFasnhCHmQMugDD5epgqmTDYrJy3fYzIQDuu84
FtzzRy3o+VIO3tORuN1JLzKW6htVOuNfltPAfvmc/hIMTyWq6Sh3T+loFG8w
65/2gzFhvBDNsrlDNPx4IRd69Q8J9dd+GbL/r+rcNeY4IycxyBelV0T/s9By
Wch/EptQmMMGBPaaxPVgOoKAnH/smSKxeDI/hEyOvkoFDWNUeMAziLT10EUx
k96B+DhHgMRjlyrwVGPyM33uTztHNzEdzQgNz7FZMdy8tfCY6DA60KGCOqZ5
VtynCKN6rKxslJjoxS5Lk1kh80mPIRWswEqrNGJsjku6yabYfGi2s9ttKVgB
AkfV/EDqjAdIKjc948PYKk5UPBiAxNB66FeZmfwNYLRVEdtXEzUDBRwV9VVT
9y3iDOs9IZQAcGLtJgkgcWxkO65EjphKAtdEQMKXGknNGakWBNqqV6dJ2vDJ
yjzFvTVyN2XQeuOBHkuavMkfB8x6/WzuvnvpalIj0CzRmigehl1aH8OatBhb
SkeDas8NvHL+7z3nwIacV6cNkM3hgNzYzmS+ujWnsRdVnBySA5yqjC4lxSyb
Z2WR6GJJxSSc4BGToKChIi0jENQOm6MzoXURB9s64AYF7SpCVm+BYK1zULKB
PucbbdHVElvpROzFXeqD8crKXUOUx7xM6NMZ6AgAfDkC31bv8aLQm7VAl4dz
nDyOjLZchFmhiRyHnUkOm1Kq1cq9nqQeH3vwNpDGTyGzeJD/Uv287idoj2xH
FODYpw9eXVWSYIBdyqV3bpAYY/j9czzZMc5cYwZl0yBDr7FYaPs7F0qj/Kxa
9bGhLQIysg0igjrzjjg1nVfehdwz175NZRdOmdM1xVxMglLmuebfPKiSImQj
aTWTJsuj0JDGZinF0Q4XZQC1G6RjEDxvIVTc+v1AWJFCym05w02zjNCx+SEY
iXs/aLMrgcUjpn/o3pPfvauwANLLAzhPcRUdUn/DhfYRyrFqnWpTdY4LzCr0
THHHCCtrbShqBGpiv+G8jIZgexwjqQd0K7L3aLGotBfJNrqOT8rGOvBwdLga
QZrm7jUdo1U3apsk4xr+1BuTwdXL877u3MfT5QXd4gNFFLyAr+SM4cEJ/+RX
o5jwwpKVKSZ9e+mqsALhfKnPr4Bk1W+IknNlnIofc6wYw6kjcqCJ8nk8jo5Q
Vf0qokJIhnJueK48C7sqd2jpROXsy4MlZS2SiJtbPkndIv0fl7SxWBc5VntA
xd1dldZacBmba872ozJCjeuF1kPelI2NPfhaONt8u0QzI5UGUvdsAEiZN0UP
QAEJ2lcJS4kj4r3REItzP8mOKYMlNcaknrPyFT+lyNjntKT1fpJfyDyYLBgR
zqykbxBUy/nNIADDBYHxTdOO9pkEYM9aJPkbhsjuJzBquYocc/T2o5fd4YlQ
bPvxzktLVBswgHYKpoddWPR3wdXg5TptCyELClRduCmAg/vE8lKiqE/7wXW7
wBuqexa9fk+Fm//4duHp+JTmAi9XNdcuDX/q26tOd1TRaMRZkXxZJNzZ6zwV
xpnrV3BEPpXrLyO3hsla7tmT86SXlNWgIcJzVVZa24bm6ybH+ZkZX8QpBASu
QPp/wmf2SwG0oUHG2JHc+TMexRZEtkYoslj0y45p+FNTBR83QD+FJPD2v5vM
vqmqeWvhIzGQ0Eb9B6NQwPLwx/hogsz8VTsYwWcU2Mj4wYDmnpAgzBxu4GuW
wHZe/iz5BWvoXBaJiVgKJ0H4q5k3J2um9IrTKuTTcjsb8CktYku5PrfH66Cm
519oD6Vq6VIiMRiLJK5bHd5CeR+uSZlangVu9bO803QB++OUUC1bYNYiUCL+
WMuncz46pqfM0VUyWVJfqrdYC43Q6hvS3gOnhajhnnkfQCj2IeMUaKwXWXiD
eQiqGxXLdCcr2WyLwYfDEBozVCRk3h55jciDIgh/kEFOsXtX+/dzHHFnrw0t
2YUCjlNQa3/3XIqDzzKelOM/4LWt4tQVWkDEyuRjXA9jTfcpYaijW5Kt2D7e
UYpYokKIE0JznRv+rrFu4iQXyOH/zxv55PkvkDpT2sM4M6VtChX3VCsDY4a6
dQltU2mmaNBYB8lvUrGG3qmlWlhzStxYbeoqq3RNjViulxCc04OKDvUj8gP4
lkhGjyOjHSyMZP/ElcZQtz8AiqWRo7Nyy/moAVr4pgG2TuOQfHro9vMVStk5
L5ihdfggI5G4/hoaXtLU5daqC0rGtRlU4p5BzQkYnOC4rEDaYMZxa3BQLQXN
bxTR0pR5OYKxIRagfOsrYKchxzoqmf+ZY1Rltjkf+48lOJeOeF9LQR1Dbw1a
zTYCSyuJB+edIQ9k43xprg0VPDvgFtzFUb85tuWAmxddX7NWs0KlmblMe1Yo
gxF/eYra2ZjVRIwWhfV0J4t8zdeQf+6xuPe+vV749+SLXO9S7SzZR1wsuMD0
I+0FsFkmWWZzdqhXO3OSrsnMxdwVXGgaSwY6vDP5I226hHZMMsQNF2D0cQTd
mMH3/MO1jD0yKn7f9eCbwZP7zsK6JTLD2U0/Pxmq7i1qDPc/vRsW1MIUL0Mm
+Zpqdr3FrZ+CKuPBwXXucqu6/SNJHh8LFxl+CZL5txBwHY0LeREZTuyeIx8w
6nUFh/pXcU/cXYX21eLbjDmnLJJ88SAxf0doGXB0S/NTqxyZ8qOVpMf7kwTC
aWQs+cGHNcRN5BL/Wmp3kPhtm76hSO2B+hiMaPmF8iPnayu1FWe9NYSiPNqS
S0OK1YFTX4HbtC8MgW/RG3DD65rxFUoy2e7vw5pLoGuftOmTc1VS0yz0z7yc
Ub0oK8Lnem/wGpb87u/7cOK8JHRQwkr2OYT9G0ZrwkjaQA43fDpqK4+z4QiL
2+nydWlXEBc3IC9Tf/LL3pGnODVk3yhM+FLNsIbonu8CpE5PN14SZDx2BzyQ
knYt3GRWRoNmYitMDeG1EQC3hhEUSXVmPJhSikXMwGKjDVvv4DJaWAZGm7+v
psrjQ9Uyj4/0Bj5u7qw5uOTVRvl1Ms/gumK1U73/7QLDI9udpW1xc0ALsFKk
kVNbSLtEFLGb8EcH1RSbL7DDBtuPEro0zy4hzQVP4jhC+ncl/LbWLHvzEkKy
aQ0l2hfbxK5CYsLUMCjgxsZNbjxPwPCdqCgAhtyqM3nKiCULL3NpQpt+U6Rs
pPo3tnotWOTq8aDhSGkK8XsCkSmNjmel4dXPV8A7/jPz65sAYFjmmxc6BbnI
cKZYeH5neMDCFMfaQ4hDsH5JANmGe0iNJAdJH8y399REPLOt5bVbYNm2ylxr
c8kCKlTfJf1dahe2X57PGeeN4ZPpiIjTy9Yatc3mdj3f7GLhg43l+wRSu+Km
5yI74YapoKoj74Z50Cvp4QdK90A2kn08pGOt2BGenKEL89MZYmeKRJW5u+va
1evj2apSFfW4Cl2b9bR3K3RoIeZQomq0iJOx8iUrXCMoGz9miCiDTa0uMEZc
/yHq7DayEEIuxrWot+NpMsA9VBBkFAxHdkB5I2kslJzu1QmerLKaxZcMsGhg
Rmp0VSlkaqpjisGFQcgnmcuV45psKuxxB3IA9R7cCeeuCug/AdIBmTO/sJk6
pKkMqn26CSgNPGunRXVOie59E+Cx3q63BOJKvJryA5/U0KL5Tp7L1cQeTHBA
/aYZ6QQ9I9pJrzlNAmJoplJ2noR+W+jY+wBfcnNDdFlKuxpvQ9mXdJoNYDaR
YLWrD35/0hxmwoxgqmyU+tJfU2ocn2nRffVVZHHjGZzAMGq5oRDEO/gWyuYd
f18/SWw7XaB7V3mkWDRXQhkOOiUkrnC/LnTbtORzSpfsv6KIneH8cvfi7T8W
1BP2V2dDODX7rCHOACFMZ9qNk8NtjyE5SqptSxc/ga9nS3JmWujNEGu4of1b
EOlVks5nsd9TNDTqMaH/tQDKpLARxouRm5FD2ZsFnOnlSsKH1reRnwxqBVU9
BWGnaADV8bnmCvsU0PmwgI2cpXCewcr6utiDqnPFvasVRo03HrGw2DOR4Tss
uA+62e9lNQcuziVoLaInxsEPom/cyd+p5YYeen1uDSSEBMfw/u/MYGvzJujR
Q/NO7qzEVVPEroLUk+cxtcaOljjfdqS7isGgCmlPHwBZFV3apxg95gzro8EH
Go/9rKkVHMOTkT1saRqDlRLtK8pWfx+d3YlUWXn6/Uns0kNstRxnfrH3VeP6
jHfPOmCPMzUUd9Evj7cGmZWrg+4O+8AuPymu62siH2oy6RMCi5NiakN1C7oT
2+B7EMZkNTOsvJPNynTnuZV28rE3kFKSL2m+0FFGGMbGUl0xL8HWHMqM9J9D
MfCKUgCwAoy8TkASpbUV4dweRaGMgsQ8IB2OhyRQJkcPoKiMxRFkrSpbg3Bm
f668CnXJ+Iv0ZI0l54+ikpy/RThpPpnU+eQoIq32IaDwZ3g0O9zNmSXn5Kf3
mnsXvOIgt5sTlYLR2r5/z6aaqrHuoLFfJpKHAwO5oSt5lSzrFX4yyrXf9m4x
HW3UYC82lMV03jml5/MuUBmE8cvhcbV0DZM8ryLmnrWoMgIgMwg9leyC2NZk
4fuz9A2ie+rqb4t/rWh/UNySlMzym9GTD4nyIBkWNv9RnWO2BD/cjOz+Lk71
CXtsVhtU0AXUt0fb8c8a5KjcAZHzwjNSNgYHgEtLITGCGemKGniIs/IihnyR
NMTvicABEeSSKedm0ktzi/FdMeYytcacoBQB1/3txmohgCBdYzwwS3xODPHZ
uZBZ2/R2DxECR9OtTHW/YhumkJ0p7kFITPiE1ELJxtI6zAD/+oKYsIde8TIo
QndeEXwcrTh7TxK56F6XJFjvD8GVTLlpTyvpYgUJatisfBTNEWm+n4WWg9Rz
i0oXIVZemhRMvhPR6M5tWcaaHzeq7CjoAW98eK6XpyYRodVNdfUgRN1Efz27
0f0Cwrl9ujfE9CCa3F7vnD+hms/w1p1yVY4kIDTLrfba4lwJnUdA9gLxjUHH
n3pYjVEznh9EW2ynzU1UmFsqtlhaz+Lv+X+w45iJ+gJStVMU23BSDe6oQ2p5
BQtaw//S71kDQE4BO4qSgjkbUC6d9Vh18PlogoYyH4FybunL+SQyWiNbhtnx
FQzzi8dMOSfuSjCwjndZaESa4q32dGuEw9c3FA8Lx5HEGUQ/+/BDYGGz5AQn
xkaNE3kv4kCT/KOfsjzbla2C4y3nmxnq7UBzyG+tIMDbGQVY/CC9e5gZslOU
U2B4cWZg3Wcd9P6uWBbXViY2gJk6Eo6E8d5Rt80RsaCvFoyYmmp8ft/bzivb
+rafHDj/tPFEC2/uk36KFxooGhEvggKZFCvBZVbGVFspJQBLu6kZuJ2JR2D2
H/diVVfEPBSvPlkqAqJqdRv3onny3heekcJuff8BdThdIrMhWwwe6khwDP38
r7EH5FzXxDp/KWVCRrk5Zdr7MkjV3PU+s2lan0paVCcGKRhr/JA/Fl+72OoZ
Vox0sz8U2bzySYgmGman7c1qz4/0tGBnRqAT17rAj1jC/d8NVYDCHxvjb44U
arxJjdjpnsad8pwwREyfsToC0NLY2ZvRm8YAP2wDCtUFPq/WG5OvCdwWNjSU
pdFA54a7x32xtI/SJSoqss2R5Cy6ylMVvfMK9iP1XK4LVOk0PGgeUywGMLyJ
GdCq3rgEltzebXnwymyGfnoXYAhapl6TDZ4XCzGOsIJFAUxLdch0QBejDNX+
X/UortTkR+Q/mLx16bO57MWP7Mvm5NnIhGuMACYHl9Fm9t/UZ7voq6fuAk1F
O5WDV/H7HEebDQM3vYEMZwx/ETCuRCj9mCW8y4ShaeslbT6TPkvRTZU/mnew
26JWdRb0BUfU1S5HtvZPg3F9/NA+sgK09B3P0VaOuNlInAhFit5VfkNkr9en
inG40la0cHsu7jsW9mBjo00K6/kq1nRBWLv6i/d5ucehBWWrp0bELCt/LP6p
P2Ju8MXvahWwptp/2S70u9lbgTeSiKD8Wsqo/u69tiQ509Fa07rHDB3alR7e
j/wPzrjEVi6yvateJ19Js7fuvSlgegZqTKYWPg9b1swTThYiJFFI88eikNPt
tUaQatMhsoPFxYw9gZtxszmli7wcOdNYXAVU6rdvrQaOSnyCVBsjtVPbMX/f
1ovQciTjs68Fbg4pE/jVRj2eGa5G8v6f/pzysHRB5knVMODnHNJ48DUNmi+h
M4JCQH//iXKCAC7ONZQVGYltmkbDfq06HpWOqclVTbDT6jLZtCwl+6uG7HFG
UxPVXqwT//CoaGgWuKlgCGpnbRp7RJp5gkOQW9duwIAHGSL2UPNJPPJJ/dBG
8arcw+olYSMrBd+HrYZcXSMmwJ9N/30FFh8KoHVE+W/wxgIihXVtOpuudjra
2nvRK6P1dWlAHj0opFipXFkqDiMvPMcfbf0SW6r0xr23BfEhqSf2xuYxTvE2
L6zRaQ1Ixp8FhYXCOc2yzbTgb2VAxm03+f1Jfclv/D9dGhbUW3kKzvEvaTc3
Iz48QXd19AfTl/ZMYH1g22w6qpFOwVDGx4DDBQaYw34NN1CRaDACs5ckMOwX
KjQ2ZE/hU5GGGts5/iKAIhy/NBqSxF6jr9832WnujO+Nmh1KJQcyEvizJadb
rMKfF38U7+Dv/DhzpnSeXvHYcDFI1SWuV7ROxl8KZUq4h1eDPWbLbzjfiro4
7NuYvvryAbcQXCHcltt1YeeiEVd9s9kq29bQRRFownpjiubSjLh5F4nsbmw8
6nLzoVCHg3/lSCmhOlF7CAaI85uSE90jSFIwVfMikKdE6uMXebFVxPVj4T5N
rxD6tL3OGEoZR7xq5d36Ou1E8moMzOZSLR4Y0xt/4ez9NSw3bNnDOJhRBmc1
mUJddiMxhdnhjKvFgqZflLS5YYKd3teILQjyaJzYJ1xMhvb11xBsyqVjhOI7
gUEDVNIsuksyxRF4dxacK0k1mYaxTM50tRSybCcMopkb/v7wbCWTNLe7zBwk
Xcl9rLevR7HSJ5DZV1D4bylutzOlCTuDwNlWQh3lmjKTYv3O4lcMZzYdVSg1
kaDXzUQmgzpc4dh+ostjBZfnZIn9iUFub8kTdu5Pcz44oDCmp4u6QyY49Baj
L5vFAz7CiM2kXY5MGWYEIjH+9/s9qjxHjFPkeeGXPgNhElrkyfzSw9B4O0qf
df/pkIqecl0fS0PzS8RfTY12VkAnZX6C7g/jRTFmnqaSXRmYP95GECJBMx6r
h0Cdihx1UAYIk6PcXvwHNL5e7e92brqCFc3vfb/eAhUzEJIsk39UF2kTqiui
tCvzUPek7Fsxt2bAbtcD69qv7+5Chq02k4mT3+NIoHeolI5VJcXDDn1o6JLh
aFJPb+9WB1BeKufK75KEoaewCHp4+aSaXytgIPsuvDMKcFKLu7JRrmy/V1hs
+PLHi4ABowgLasLA4T3dpYxCPIH9zdifapdKww7emrViiTKgZjk5ZuKDLb3J
MzWDT0HfkfFSkd1wcEe8Lh04ZowWozcNXONwF2GJxRpWWsGNJxJut163ipi9
k73IABUN9oIRD1E6GWARUzmFMHZCbH8wSNHbxFru4sazz2FQsz2CFxKo1d2s
QVSjoxU0IL0LYECGc/id4GVrW2O44i/+YIhL9UxmKSdhr1a6HRKJJ7IxuQ6U
n9SNmAK7rpgoYMFSZZsWbObACHGGZFsvEEVFPX0eP1SI7CK79G9iEh3MPI1R
+y/lBzZFY2YL18+pJnR3JQH6E+HDRLiATx7QDK+IxB0iQ2LCPcwTcVLVETZd
dSGaKNvQ/98TRvJvX/YZQGdmIcCLqs+iCHvYjtoR/0f3clZKI9GzHvbjzosW
PL+6qHi3uvgSSLf9HRinNF3GioxUD58lmnRUMwD7pWYzz6EppZl6pH1LITJQ
HA2jIuizKa/yb+vA3ElE8qeBsTbA0xuwu6hmv14vO8PJ5725/Src4mTsRwCP
FqQN1om3Pa8CoOhUmop2Vt5s3VuGwY6jBOxblOCOaZkPVtEOtEDkPCygmoSt
DpSNCF+MMDeT4SK2dNIdPmzMieqTTY72yyKjZlW9IBuCBD4sgLeAPEGhyTSr
3dqy9cBaNcuHJS7sKA+MieVbdyuR1rtJotgv0iBmmdrm7YFwXHgY7mKoayer
xV+Ul43MVVSlIeyvDZCTBtWNny/HeqxmBIVkdGNG/BmyaIC57nwlE88ti4/w
hC8Jup+OA4vS8EekAZURvjlkIrSB/icqw1P6Hs+RpgaZu9tTdpTNAGYnvP/5
g/DhKfDkTsPXEMUOP0dPwsUoFlAazM/jYHumu3Y2xV/nnVcZV0eUyhpEoBux
kRbl+tmBSdNLtXTurncdSI9lP/R/xHocpSIDwX6VqeeR4+vnqNBMHVL/+g7T
TuyXyr5VG552uh2cxYJ1fy/areYWSJ09eGekFD+h4OVk5KoTLECipre6AggG
6jmZgVIFysoJL30VhlueSe+bnYAcUUEl+KUXq96w/TVYCVdNXpgSDs5sQlar
NKWMVulnItxaFiHwuqLOZKmc35//NeK4Ndep1ktnyypm6BUdJuf693r8KQz/
jYVxOxKyAj7X0pyZyKJRERXKklA8ziTDYdoNC4m1Cx/SF5BAO2AQAs2+QzYs
NJZoE14dv8epBrg1u8jRviNf80lR/9GNDFZ8avcoQ13yeiYsJJA/WU4tPllq
qAiURACGxqipsANMi5Dt8m8rX5D1LujgAygNt8uTjyvSTj/bDMduMerrbaam
M0YcDSePhx4Eb7F39wszPOyETeBkqxEguKTEtcAtQY//5f3rZ1ACE9OfhEZj
CYPAXrcCSSV6CjOzpJhrMIRtI6ofEGm7eFg6uxBetzzNgicf9OHH7yx15450
R/WvuNteWmVkbh08DpK2q5cBUTJ9asq0uASKhEu5/XPgPJbSSUMFaliwkfVL
KGn63nUa6kB8qF7QIiQ0kfpXSXGeBVPz6abwqrsCSe5ZoUq6RQt0AlOaEfuT
h+TcL+OOyAS9Yz2PlafNdRMVTzIXOzLYcwjR/3yseTBr/oQvIgU1unMEI7AO
LqYBVxutmY6FsuoogpOC8ZAjf+m7JnktYjxfabL/LVFQcZFw4R9c2lqM1eiX
yPoSpTqpnx8uAXSYOaLINJr6lOWfEYO7txs7ntFFh/C+6frs7+lldStf5BfG
FWV45K/E6/UE6F3E

`pragma protect end_protected
