`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
O9hn735AVDUnsFnlyQBYY0+6XIysb5EkqyhjxoPb3UuCebMlw8CnHX1vW9FCVcEM
CFrPXDGY95CGExu3nANxXvftTdmEelKCIFNn9Fd7Je3sN9tc36FG3PIb/l7gugC3
ZsR8HWl5aqzYVk7uAk6/lnvWpTHCXJoU3EpYxaHR0QM=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 32368), data_block
ILOkpf+Com8hSK6TYQg9o1yYagdQRIp9i6x/457uhqTv/86OaWIlpBU6RoJTeP+0
F8NswTxb9YEYfK68q1W8dlhKfjZCVoDHoFSbt7K/+UusrRjyo41slJtMl4ZgGyCF
u8nuhDyrackhu+zu5sSCpU1YcDPVX83+hDom/x+qhbRv0ANrl4hpblNdMBB4zbA1
+fJIP4/w/4P8GvhQDgc1qoUWreAvOeDv3rP49onMzDuLiltGZb/s+PAuM1O2LpNP
LfyhJtkkpVPe4Vi2iJTSgchpkiegrQ3JuNmADh7khAEj7u0b7b3sWfvbRds2+XGO
wYCBWyueTJfxYFTkUzAkcdzzn1avhg7dP691SHIPywUOaFireuRh5Q4he1ymIeHw
nSDIWmaalYbPotilY9PsASaqQ1we5QQqPRF2XqxJ3qgkF0W3UqX0Ji4Xhd72Nnk/
hea97dk362x+bf0OFe05Udd6PMQzye5vEM27g9KIyZ9UF099wpjet+i5BaUYKN4y
Lhmp21+uvnW4aay36Axc93cbJ1uSX6sRTrAr93QxRWp5isScswGSJ5yp+rq0XJ0r
TpjQkCw/JZTG0kAF5f9CPdxJUeIo3XCO7NJMbG94hENZ9oiPNxuum0TegwqTqUUg
nNQtr01SefKergJ7hmQwCnujExk9vnHCx8qpE99pTgthZ+r2AN0jahsMowZioZDO
fNl/dZJ7uUYaabebkk06qIdqHMO0JgA7bAA4q+1q5CPFjPMkY3d9amVsd/yg+C9q
O5D/spnfAA+wDBUCbFERG1YkISjFXVGYMRHXMR7r5si7m7gDAqaFTfkqeHTbm52c
qNPlxW7N7kJWGd6epymfhtcDrv7G1TXbDNfFWo4kEUPhwzEHGh9KAN56FMRpLYzd
uyMLlGSRZMulWGEiML6tfNnYUtogg7S8eErUF3STg1opKeuXDrycdrInymbWcNfH
scvkGeS6w8XKE+Xx2M5EX7K46Bt/pGVkW+TaOOV6G8ZsQpne2kHXbII+0JQ2VwhM
Sis7qOhNdaKCEw23bvLejiDNL67R6b1WvO8XD9E4uU4ITU7cRIqs1K1PFOXobPmr
GWAnRXmE0TkwhxhMLjWfjFzCOqjEWU9J44rdH7scMIvBkOASOn8RfoRp4cUsrLtU
dnHQNHNvsIxM0STvAKxDrcHnbRguUUulz0dSzjVoFGuuVOR6lEkdP+NzdPqfAvyr
rADsibtpJyUyD7S8ljjJzSbi4Z0qjPY/dLPVanFSm28FUd0nQOOmSHxSWjAENWug
AtxdC9vtjntFZHVv+/yAQtkQNG/WApPoYkaSsHSlB8pHo5aDNESfBsUCdFkZDWhQ
7j372yex8rwGwVgxhZkPQOR6cu7ACz/DsLCXLRL1PaGp5cD5x5Q8u1In2loZFGIb
oG3WLtvsFiEfvXcWTh3Sxpki60Z1GcD51LXrhpUtQf8LxfDYVTYHN8XhrtyXcxm+
TXhWEYyQnrtRc+OT5oDuRqCDKRdEPhGQZsf4k3NkEiB1azKf+I/Zb7P1t98FuWSv
pOqDjC/GjJiPUu4C4q2w5eUtjbDp2nxOPEQiXoDwHkZeIQOQIChvkOR3DG1KrynU
10tno5R4S5W8E8HjAfUnUOeMQ4Z866+KptBFjqlF7scAv0qLjg4MQnPnCfSQB4hS
HRuhP9mzOMeSLrIss/4Q1VqKGliJMCivBZsJxozOsCwQ3v2o+6a1jVwiVVHdcJSz
J8jYTw2MNetF1OQeuOKFTgAsXYPK+2U0xdjrIZqlnII5wpDNUh1OPNOmHmixZ1G8
UBi/YESCymQtITFQNWKWXXmFcDoahl3gYdKNQuceVEc+3i+bRdapXi/LHx57wZx4
TvDop6kOiwdHG3b+NpqbmRTCIACUUNEQMcrokRYepRf6HqxQP8QdLx1rFAb0+ppy
C12vryNzNeGbKG6/g7tsBVUVDlm+xi+HJHcL2vbSjBZU0Dxt0b5yig9CIXo4ToRs
2R3D3ifv9eIWZxsxmnBSLEnRsO/BgsKTAe4NQYGGvakNPblLFDgol2dQO6NavYXf
xJdxceQ/I2epy2mcEbupHgY96Vjl67BKY58eL9tzv4KIj205k35YZZmOLvM8Vb9A
O1Bobjs9O6xx8B3QN3JtHAa4R4xXii3QdUVowhMqmtDkoMMqdS/tUPR4kKHptT57
lFF0YBYnzwnHCAV/VmYTLNNdcjhVVbb3QBb7TBVimhmgjGYGWD+pQxVpxaNzs4M/
80Wj5/nsV6fPnQWuzI+AgVoK8oNt1sW1MgPLI2pZcrbb4v3Z0qlbnFXaBD/P0L8i
7W9dRwlZtF67w3oOHMbgs9W0lhcquzgE3xlx4sMzU8qUP5gNp18vo7XRM0Lo5ZbL
UfGIVYBqqOr8QvtUMEhdBqjfu893zxsDvIxZ4IXzYpoe+ugqXpxEMgoQvgq3hCo2
D2blR7/ZzDMd/+WU6rtQy2J8lXk37tDTaF1fw0otTI5EIXWUbs3trWqVFXQEMyU6
/p3B84XvX8Tpg5/aKSobf9jQJOft3s/NIjmkn2/nuXp44TAZC9rqcjnj+64OzvAu
OPLDcTLOY+M+iXiWnvgNFyB+cREejZwOur5ZBMIeQvo5aUDF4X82h3ivONtHmO7E
KT8HfeJV61bsPaE+9ETi0Dqeoa7EEKE4kj2sua5zIPJDl7f7/g4eW7fTZ1eEh0lK
uzUfNcKOPMVWe31dDK5t/sb8FUO8zOJhjbnw9tzzDrSYLfinIYjx0c7evYwTRHic
sA73Q007xrPRaf5r1ezQOYyLZAtmoAJoKQ5/IdYB9zo0QXkUClUYtW6z/PkrBMMJ
ccl7woPKmkepNbO8fKGAadOaQzBpyDHNIeIpJ56rMva3MQNLw4vlwcf+Eivcjs6G
aYXsqGWKikBpEa6fcoRB9LMkdpqc3Lh8kaaMeT6jcCUaW7FP0LQXFPFrcr9wrq8e
pD3s6IppeH8Yb1QrVYIPqCz6S/rAKq6AP4pFRGkHIHZ4Fc/QCzgKktmZ7dg7tM9a
2J4Ko++1ZHHn9W9BYS+K3ClV2qsPhbHpQ3bd/SOYZAkvQ8PNX4YcLAT0vYg0ZU39
z+vc6fQt8zLe/JhrCIxZiBd12mlh+IO4R4PTquTgiY44oXllJPEsGi3JP0plQizp
gCnBQnEoywdByUbbrDuIyyBCgopgNTXZsu5JzzGV5BAvVQ3ykoXL0rhO+SJrd99a
URX39bxkUe5Q4xHcNT8tCbbu/6TIzefK3ZJtosaZ0sBy8Jl3WtT8skljW3ZxTqxA
FBzQB8GJPxlqqQfVSii3j30UJKJx/bNID4FrBiErAFhaSgWDeNk38kWvvJ88yKrI
YXjTTolVZyoN0wQwlrOt8Ulw+UB/tTmlVtts2cPM3fEDg6cgaBwIlo0EZnNr6Di/
/UFre11p6XRWX9pf479Jm8WUTUsUEei/n2yj0sQ4BuMOevLVRWQ4LRbxz/NDMYkH
w7g4Xs9gG6AbY5t56hgkRIlS8QQxDMc5XkLnbUB3KdRrPJrn1R2vwNHx8j+4wXmM
WmRBKnuRwELbZ/c71yJxRFx9GE0VBpUD7Vtz1jEp6fPHy83iyDqNxeyCoHhFTw5+
HldrWg5N4XQfWngrnCxsyQuAcTyx4Li5jApH3cLXs+Cyz0PqAnrmgUTqj7rzTXxw
EaIH5c2XylzlH+DCjq/+qZWuhlEgaIbbKAlH9bBGrNxgrygP1GlLq5KWSSc85UbY
6Tvif3xO9meqiApxQs7eBR81dYr1Pn/tYzKLsndLF0GpvTdkPjp4m2Vu2LbGhvKK
CwyyTS53sjxYuaxg2VX5hC0diHfnu7avLZaYGYvr1kTylb9F89Jmp+8iP8rFjSj7
sg9Q93RJSXGTYqCd809imuyxLEOAXOPGFKHvZlPU9UYBFo5ft7ZN1AAN2zwb2qhu
vSB9D40JJlWgyz99K97N3GgGMKqYo0bbGnfSCej4TJYjV6Yoy1WCautiQmUBVj90
4WUlnnEgHbdtd7QuNxJ4r+DbTVot2uyZRD2QV5luV/hPXVhRcYskwbh0DIW3lw+G
dFEmMjlYVYEpHcxT/BpKPMWKEpCskn0zkpeTW7/JKC8v/OV1t0CpuUlaoARSFStd
t+ABcDagz6GP5wNusejXD0ccDRyaF4vxnloVNLSAB5wviV0bybnNxau527rFHLZd
/UKz63pqtN+dyFzRXiZJ27NxZ8WcCGzDn3idaFzDL+OxcpCF9qtgyT/e7PWLWRFM
IMZCvucXJqhPXnw4CBYEfGN6WFd4NsZzhry2LrBC09eC1uY9GfDaqa/eFWVCCtIm
EPAFJKNBBZfJ5Q0yJ+1b76bnmBMGY8Di/XqJ4TmdNbI28LffFRRwzkt72xndPQdG
Mi5vFOv31u0CQQIlFbbEXuFzUjtoH/aNIRwR7S1Gu3iSuGeyqQdcjYFThyfmA62R
UJcOncUc83USaUOJKPHTZOrN536eIuTl3qhyw1uvhh+3t+OQNST8JYe/oGO3GW04
J9o4LL2+WxZv5zWphjnO9lgYwPEE6XktSHCAD4XfWFTF4NCHZ7o2bLWK9gKqs1qJ
qjFg87MvhPi53WtC9+gI+jsMcnQKaW7snX5polKYYaUuAjlU7VPPUINRjgLj7ky/
LsIK0wBi4bUVZeFjYdYP5sz0HzkB9GjEd9yReWW7aY/taBgECe/3Rt7hg6ypDsVe
4ZgeEpApMAaVRA48kRTpdsV7MZzGrIx+q6icnp3jAWZHOgC9jsQ5wp8lVXkRaHHw
BuZ2T4PUerBjj+54S2Tv3ZWvc7k4/G+OlcI8JR7QTA7t5PUtv32o0cPjCC4U+FAQ
1nBfXrvCd2bz+fOQDBYqVoB7+lLaLoCeCYnWGIzQRDyt4VGJq/TJooolCIYVD8O0
jjkoIB8WqyLZFWXGjfOPKvwPxgaQAAlcCF3GKONFNX+AFfxiPQiFPqQdNfsjIOJh
Yu/dakkMRDMkwZucVVvD2qrd+US3zwTa+Od7fDVolHmPcA/Wole0RBtYv6JO5Xci
qHDhuoDGAVHW3DJcf3Mu2tGYmOYiwgzUYDow7JECe7ZOUIDOU7dCAVaJ+wapyQu5
NZD6L94B2keWLaBZ7tfv3DJvtxfYCp+KPBLtkIsp5VxcgoFP7PWnmytBuMwl8i1i
+BVAQF5lKjpPCBD8Cz7vFEYMWhMyltGCDEYqi91RcQ35IQoaT6EvQHhZDSR0MStk
O2pj0NlLm94cLBmH0ZsmLSxjVmXuYmibMP2UGgqhaTDX0On84OXFdzghVdhsw8cK
TWWVhLzBL1pMFEsqiV/6vFTykH77BT3Qm+FJbMkWudYySfpCuVK69ypA9pv1gLP8
UtQ1Sk24GYIw+Tghs4u2oiEhif//87Fh4AHFD9C5morppOFkLYAOVLqxxQlo2Tu2
9cmkKbcOqI2glf0B+qDf3A/idM+NzG8hnvcEUzxGNykDaPY5Dq5/iKgkVyGP50Nl
xrlkSGHljugIEgtq+TSeNmXEr2ZGdwx+xXkqEFjdw5kYP5bltFWHocTid15cUBgn
zDJFv+GFSMXVkI0DQyJtOUxSV2EOqngaLww8rnSry1WI8fgdm7P4TZLBpiNSyaCj
Ugu9Wp6/0aSMSb8860bIG4QhP76CqA5hFnnA7WWebbayeip1fkEA9IZxeA8wd5OP
AjQCFOMyqBmi+Sc67pc2Jppa6dVOoHZpRnhjoexSlY4If46bQ2LzHlwmpgJ+5muG
a8WnNP4KdS0VhDTw+4wdag6PUbIPSWmiEoxW1aRl8hCxSX6wcpBBFH5oe50Mjwew
LfQKpNzqwdLQ3AABwW3aIUQ8QULIps/FAchNvx5DVSNENWCUAGorP+0F2TL5KJbQ
lOn7e8ZWNafq8/2a888blj/+THbZsJvp0d2/5PS+vtlQ6nebOs+K/sNSTCCDrsXz
ggmt3q3ckJhqakCp9sJEq8hOzgfIGv2TT7SEuv87DmtrKloMLdldnOiTcsq63MmI
XPHTrwZnfYI5MrWcAzfKrhOqhk0DNv/ani8ptAugI7w7gNCJ/jodSuElmo41HeVB
W+hLMS/YRTSAT/0y2iySPJOFByNQwkKV2bXX+7R+Vanp2qzVb0SpgJsabwC0Q9rq
GZvbChS9fYOnCNa5D2Vsc6zY+aiPdzpMme9aHJ1V2+MNoLDsQcZCBJCfDTOTdwfM
pn7bYHV4Fjw18HnOsMT1oLkql7CkBjTBUQQx5f8Eh5u/U9HUxdnLFevBVaTW3B8y
OosYgXH3wKesCe4DfPPJn5VbC0DkbYQjdBLGjwZXhiz0ryCvSGk7KsY2vGjLdlzx
UDPb0o1Wq24N5WzgjJbuqOKOP+rozsB9h+d1+crBY5Ykpn+OYypdcXQe5ztZ/AIY
csv2337wppcKCI04WlgulX2yEtMGgB/xrEK4JoL0RYx7ZAk6ekpaoPlBe84iF5Mf
/edNBKyXr7nLmGcJFQPoRjb5K+8U/PmFGcY2v0rmi8cG6C1swA9/SB1PgIm2D0G3
R53ZvW2jMa6/LjuQKvArA/kW4AXuKF+VL7Spw3hfbGdsHo03eB90GG2p93DAZ/FI
cReu8uylz8up1qPSq4sYlpT5JvdNlnYx2dJzZ7Bpt/5Ogqdo6AVj6xLeBuCVvWeV
CbQl5g9/Rl/MJ36pNFVkKGlseJCDF6zjcrB0aUOR3gRLXfVwzUDQhHfGR780W8ML
nL/7AVXizK8EAxIgQ2nlx4NrafkOjwkNC3lkNjB9HoiHnYMMybb+VqgR4iUoLZC3
oFZRoj9hwWDXL8tODHGNE5fuxziw5Dr0YnENF8MzgSvMSQoo0CTon/PbSHRjgTsR
h494Oa7rsp3zTmj90MIfdaSrwCfTOW5wUSpXOc7PrqZzxuCVwgBnZewqFWC/2Ib5
CFP6l0/mD2RbvpxqVBBsoqy3ux3l78KR0efp03X79xF3JcheTrmXnoVfG9LEtmnA
zPqUBTuc3ZvKMkJXGGVMEs0R5DEpYHXLqsPykilCz4GdgsmtdH4yBF+wD4JXh/Um
lRDnsggfc/QADBoKIsbRMEwxOdMesWdAu9ZMngKbZeLLGVsf7OHgs99g3jgKFItf
U19A6JmnSLB2AZe6qgv3Qxg+w2BQnctpZ0XLaaG4DttBgNBMpu7ECd+dsr3r2BUA
/c0RiZAeT//a3i4svyBNJR0kq6rDIT1kypzwA6nA0B/4TmekdGcKWaqNs8WCwGfJ
B8UnnADdEJQ8nsQWYTQyfG10pf7k9bS5fg5Wg0bjCB3fUvkbB18+jTdvTRh8UtB2
QzScSQbUazBvK9eCCImqIoJMxdBon/FXxm8JKduGS6KrniGzUUH9v7DM9zIEbsqC
85vJrdkw5uUpOfbl5S3ihpm0gKRbaUFoyYEyYm5Sg0vfsZU9W7OqSp0OtaCKqhfo
UTf+WHfKoOQ0LzPQPD5xd/tueTAD/gSZ0Vk/Inahq6pRbzMLZhnFdQOCTc8t337x
a71xsK1u7DUYasSbjl3lDOcLm/Ta91fYah2At+X7RgUtmIHEjQBc7lYxMl+bO2fw
TgvNJBGYGN6HtGWEqsRRVTA/rZtOwvh5jLbclOJnx1PrHzF8k1p9qz+JWSXa2j+N
aiATQFF8E8bNIldjWsjDZ3oq1GrDdOX/rpFp4VtgCFZd6Bk5AYcIqu33KhHQslnK
XuOntHJPC6rSa/feiDA/xPXFKHnfjhuDxRpzJbRg5iMceYHlDjwy9mbFf+J63VoN
OeZ5kWTL+/YpphAZW832fkc5EokqIe0VeWoHiTDWWHOaResaoAPu4plzN8yVj5TY
xiO5RfBoxOn9zUhRs6zWpr6Kwj9ZFWcbT6DV9THBmaVHNQfGn6mm3bgm/8EpL2lf
1GVnb/iWHKyZHFNcVFFLwrxiUMHDOYHmbern4agJ/2NlmH+lwnnE3yn9Obzu+ctW
stNaxvz8tdVgZrN7UrL2JatSwe+QWT2jsIPBfnYC4ifQ9JhigIBBwJQ/sZ3EG2hW
uhtFc1DueZKIft1pcqCY70PobpdbCQLyyMf7Tp6TYWwPStbl7yyOgHtkGZWLEA3i
ILj547lzQcTwuiJkEpU5kR3RGbufX2U271NvtFsMK4zHAJA9P9fOLZFR6Ugw4vFI
SuAckzuRl1ctcPUaCr7F58e9mW6Sfq8+nNnRQoWn0kKwJ42yGR+uAa4GPr0q9SH7
QpKVsIWGHQ4CApAWlEPS2znxM2HzQi/7H0DbKE+SYE/xc8ATYWaZTtToOVSX4Cp4
p8CehvZSlVH2lfEwBs+wb7OmAtZIXfRyv2KqSiHfZtDyD8+u50n3tVCW2j6ONbZD
qi6vxKEWM1QnKAGYGx4lrIp9wTJXgmryVdQJju3GN3TMYXOYq3qe+uRIgj6AcX8u
I+HsIBVXjBEoiLJ/g4n97UmPfZT2O0qhIbCa3Mxfq5+/mOLjQStuzDhA/u1Rwe/g
Xf2+NX85CombGEnSBfnuN/n2Nu38w9XpHzo7pWA8BaNxJ+iy9sBk8ACTG+DUWFMJ
DtHc9WBbVbRo6XIurYRd5+dwcsOEkMVOtnpXd8jF/cecRtmEr73MVY3cZZX3Nb1i
e9uMuUa9I4Dutx1B7jd1e7ROvYC6ORaTPXVR6Vpd1dLSSNysFgN7F43lfLHYtbH1
tpziHmzpjtgI8bUKXcoWf1Ubx1/AwK+UqkjUn8aJU106df3Tfz3JrBwd/91E5xkX
9sn7OwuuGD15XLmLDj/WtxFcoTvSw78Z80PXiExc1c1n+9a1MSwPlx2ilSF3pUXK
acui63GVokzFpkwDHgMHgy5xj+SPPMIJkEbY1lKcy0Fr1OTJ6eIKWERp8GDO7FlI
w8m3k3DMqbJqs3hmuwLkoG+/4MZAfnF8qjc0bzAUgjohbjKw4Xo7Rb8oZldtb9Rs
/fCodUM8JVVglFKq0kjJ1p63cWFYDNpwhtw5yZ1KX1P9crmliHYJMUCU+fVwAyYI
hfP3tdCSiPnbFDH3oExsp71YEn7uyVYEF/f17cloPLLC133kEYiVAiEwmm/I0Ook
0NsMyPdve5JCBucxIdQxtvgBdHxQgnYl+o6zodbPBMmAZPGD1F6sL8y66NWcRqou
D/sHDdaNEDOwKEXdRVptk++sKSk1zOUZxpXzh1NAlrSJcMtTNykeQMOMkmja/wBN
YiXvbggFTb+jrP/9gMQQbaxanTRPLGx09O0odo9HO6X9gmVfbKW8pOQvv3glyfS/
BQ5241qMZ0IW3VxXuw7+L+0LfMMFIT8wRGHs9ifPeCygFXPNlmCAWQUdN8e7XD98
7wk22jmtgFzBo8v14Tb8lvUJogrbm/kTQHWoA/EeIHYCMxgn9qQIVlKMnmRerAPk
es12MqEv3uXaKaukfY1F6w38ypELZsZPsYdEwJmyfK3q++wjGj97aohCfEHuHNXM
Zuotyt//PW0d8kPaGKFIrgmhPg1dWeXXxiFoLQRcB9gmnQEvbZtuzlW1PEwzdeF/
taiSbBfh26paGcMIWjbqRF6WRa3qgmVWrcZznIwbLuCQRbOQuYMjTmvgGIZ2dTw0
UASKobic1xz+lMh3iVuvxjjJ2WbZA7AaGmShTxDs0v3JXiyQvd3WnQPSgjir1NYa
vk1Irz6HxaAFnwzu/UOxECwPQf6nX60OjodgbAKZmPLN5fwMbKE6Urp9BaaKPEMi
Iw1vCisMB5nJ5k67OC3Rl/ezMU800gBR+OrlOmSp++NiJKXHG1Bl2C9r3JRAwYjh
oI4BGQv1EePSgDgrrcXqJUjIMjSvmI+C096YDKBTvwFiavQNPOekG+tOTVzabsIK
RQI+sGEruGNhCLfYlSC08O0oJD350pZWfnBU/wEr+hf71ZczA/qWamvue3LIGtOI
JT3BMPjgWQ3hpszMbGiYKR7zw2VlGfP9MzhHMySqMvLRqpppnn4v1WtmA69u1VW+
npd+zKxe6Igji0aIT2CsARBS35GvLY2ZDqDoxcZ1kMp/p73OdW8Ua1MLPFb/Kas/
IVYvdRWNkii0+55TJskvFKcLP0smSKFzIeFNjvhJ6dVTRQQDyyD/R4FKsT0Ykglq
b/P59HLMn6KXkvyyCPtmvjHeKW/x9jMUVzd+T2Ti2thd6+mjHW1zIvNdO7BGTuJO
H8bsnLZuFuONau/0ixJT7h5HiyKkEo+x5tQzY/fhLZmqWYx3BsErqkssKhgwxP7n
yamEfP+rIdEWQwwN7uGad2ogopa1jaEwjN98GaEEDSpcJxsbopn7j/fwPSNDRpNO
PnwN8gZI5Rd/LSucew/asihPjMLcFWXKx2L9Oau1qYmV+GxCmWF/Gry9gzCamCEU
yi3ANbJySHiKehevtsfsbMNyy6r0eWyRMPzcuUwEijczgFo2SzTwlaSF/Byn33HN
fSDI008S6YrTy3zVz8wqhY1+Db5bsuTa6RgwiraJgnIE83EzIegLGk32QDSMCX8y
4/5R3owmZyr1L5cgbzTaiYE19f2zci9J+AHLEH7wb1nvf/NTI6HVYdGkVmD3pv9E
2p4lZmDRreuwf8mVyOlAGgglViqBQLyRYjOzk0yVroYJB04ztgB/tdj/n5CoV0u6
XsRxxgLIzFggIyJGMRdPnx/V1Hu+qnAUNx3ZgpJ4A+nyUOpA9qqUvccxCZPIlzWW
Y/aujmgeb8jOJ5hebnOre7Zrju0Iyg1d0Dnj+iPwF/kb2ULKK5/uSmRqO3moyywo
2xbf7eofaku2zYW//YFPw481GlevOcVahi1czM/OeQQNTp6rHAffSEUKtPvpBNGu
HTPovxb2z5jzZ5ZL1VEFuqxiO4Teg61LTRdavrBaOmMrKDFfK5xgiqWMzOztHhsQ
F2GFTVeoQ4SwpjJ1eRiTXplq3g4bNXdkQt6nkpPVYYQFCzUn78dWWX/bLSLJdSY6
8lyBhg0ZJ6lKszbLPjS1d2oIen+cK2H0Y81Um0FJyKEw7Zw3W9PPA0ly3l47oRtb
cTXaWgJi6JeF6JeXxhaAmjaee7BUwhpO2WSowqVAtpR6oBu7RVvdGgLKMe3jaxHo
VG8uUQuQ5yf+CnhOmR5X/e+EBLVrvKyJtUszoo4/LTYKGZIVbikbAyPZT84QXPlP
PT7PmI9UBjSoCX0Agm+GVSOKgpnqiTBc7Aq66d3hpMxHROfCY69BUTXazCxAGYXc
EDuSgvrE66nuMyMB6W2q6XB03/4CDZCxJFzxYSr2Jhb7eKGFC0oI6PeN5HZXk4iC
63xAVIj/QclHNeaY552YDtMUxA8Yb4CuUCAd9+GIJuNWPZ65lCP4914KgHQzyKw+
3sVhVxRhBjyGjug3l970/z1XdVDPLEPN2p3g7Ibo178vwhy27EvOSbp5aOMbHvE/
a62TNUBUSy1UiequxnJ3NJorG96f7HNIKJ9WgnvY7A8G6oxAa5ntJFfFPSgLlA64
nf5lWm/SLd8dSQ7T9LljP/03u2zrHaGctJoahkLVPXm6Dc2Y0CgPnzCo0lx9dHuB
59oBsuYIIRdrr5AnAapSvq451XbLGTcMuHZT2s2isb+hBIO/jEJpVTDdmuSvq1AP
lUOllIUw9O2nfGvMoPGaPZk4uTnxv2JjnyWTK6ell7kFxrtMeHHDrF5W5TulFIqg
7jewm/H/Gvy3dSvSvqbn2GRYLCnKaFx1Z3HcDpXWDApNgR/OaFQX0cLwLV+VOZMz
o/vc9xHCCvzm1w7Gt7k0nVE4ybP214l/2R7ZGwkBEY22hrCj1vhC/zYzhCOxnIQb
pwSsdN/2BDclcfpMr1ZCiqVCTUAp1Jx9iSPn2MGN8KAcgy1PbFQfQKAUbCBbez2m
BLA0rMNdmwdIQujJRf0fbz8ymDKHMkonWAZhVkKCduQeCHpo44ZwXwaL6CkNoUiE
iWUDDlDwfdg/zEPgJzONW5Uk05Ikqc0E4U5npNHHBV5wijaqjtUhA9pDgqwJWBgp
2GWRvn/OO15xeKbRj+1lfVPXOKz8DmnKPWRJ5397nkcp16EWBckViv3WL1sPmG03
vJXTxDRd1ByMkdzhweqq1F0l6FJ88jGoLWnL5jkgikjT2z8/VyFsQOz9OZYhd3IU
9qECg7EIu/cC0eHA5GRBtPH+XTewKksO17bXzjYYYqA7Vvp0sY89cT2HJgb308bx
p7ARYLat4eT0rsGIAK3rfMX+ODBNxOjGebYVUe9oQ/EIglL8Ogz2Ilf4qVf5Uj/+
9de2d9cHxOuRoIqDJd13hwxprmpMS4te+QOu9IT91ZnBMLT+1KINsU7nK44jmxIx
TBRJ/+HJrd8fMqOCR4cuAWRFv19VU2vCeBUsli7UMRkvooSFeitXF+ZaUK53NmXH
r8TIP2R7KsM8K/aa7OJEQtHI5BtN9mkwRJ3o0nWZHln7vnyDGHPogJG22X7eCQHu
t0SPOi8VDd3QiOoauI5gyHCcsZHviOq+7fFS/j5C+amzIA4gMtQXterB2i4+Y9g1
bpuJP1DLDEa6Dv59JuYgBeWB8sv+OWid8sEoVqFh2ozEtwRIFqlZkGEU475oBGax
Qf7Xp7SVJQSTxLtLIZkBpZ0qYYMtgB5Cq2omQ0JcJUX5ecrs7x44nN0UQmTtkCR2
+R/efJK/prB2zzHvNAMV/Lr9wR3s2oekZevmFt7awKHtW7FEyWJn/v+JNKSC/Y2O
5/8gMt5awr41fYyIGd4ogYlVL35Ps30z04jhwuYPnVIGfG/FFsgm3vWh8t4dnUwd
BcNaRZWhPl5a6ykUOn9UhnrEWcnfzKpholQN4eCkF+afMH0J0b4oXU6hHnL7CUxJ
YBixFsH3YtiqhgdkgeHlMoQwbFcGUyYFLd2PxbpaKNsryivcsxHgFdPYf8DjTosV
OTJheK5tlrFVuGvvy2gesnWivjnXCLPy40yO5cQgUf2+o6tGD8SHW72ue12nuGYh
3Y6rQy9gJP5lxZy++GIbAGLB47b1JylN0AgZRSlC3hTFG6PvR7wm6onV6o5D6SJs
gZZzMaPI8esdhn9r1KzMPVJ/atGAOZ0WXS2oxaRp8v0ow2EBU2s3XNlaM/J3RbwI
6W2pDOuYQS3DYGdQhJKcOex7qW0RyGJipuCF5kLsYUVKbpa4qgLEw8r+E1QpOzsL
8N+J0LgO8rwlGeyEv5RmazK5A+vM+vZzQdMJjfhUoUHzSJ01BgcXW9O7sI0LxmA6
sGXOcw/neLCVBjJPM7Xj4QX5PvxcdeudRHgNj4trx5rQnp/ZHLJ3xOJlfTXF+yk4
1fpOREaOMx6x/1bmG6dyq0r1WJS8lz/hiE9L+DhT6ECorrruTbNq2OpxJyKOLjt7
rAbCPhMRoqbeh5pQkfXi/Qk48JbA2UCx6s62sHjdJ7I62n3psqKyeJrXenXaJ75x
7SpJrX5Ze2I8e9JaNTlxDGc6fYwiKdkwLRGwdY/lxurUgwSDNgMseh0OWmdrn1Lz
UtJt+gvD1TRKU6MPZmMdyL3+N95VOLYGSpIDE96uR0ZqImKBMbqppZEWC9CmD+vr
ueU/nYQ5b1SOBlE/z/OiD9vPEAhnRdqm6FLcXpZwWqbDh75MONBLG68MQWWlA6Xq
9pNKk7latMu0DUaaJH6NX4VY1VHTBjICbvQvfD2L6h///hLPtCUotoZEwDZ0xkej
UywKE6TV/SABCmkQHacdx3rnQlXJhxPvnpBQyCXt685xkGxpAv10Z7jywnqvJcNN
2KFy9Ql4FR8Dxje0eaumCneyR5JT9OSq1K0NZqhM9coOzZtq9WgZ6dAM3yeMMQm2
4ldnO9y7lTpeGMoRpqwgwocAd49LogjcdXYnBfGOzvhIHhzPS6eki3w74M8GLI7F
wJ5ra7ysA9VmFG5xJpYAyUGVwEARkMuu3NYc1xulRFpIPNgj52Jd0T9NLAhEHOQT
7yx9f+hJMFVTd2jT7afUFhiD8g/Rl5MJXu4XkGegvHQhZaCfqggDyCOBZznf3s+1
ALLazJ1aY0JBVlssnVbCMfZ0rYL84vSgK/GUZmKIP0aBV23oW2zY6jR8hCjuxnST
OklMrZoTDM0dPieXQahQPZcYtZh6GXKmiUSnZwFkGm4tVFd8fWp0R9LUKDTgmGLt
i2PpxqW4ThJpmo9ebvRxHKT/gWNwP8IIEJaPXwsu+QDwMbEIiGFJRvicbBPb4MKB
vPazFo+aOhQkwErvPA1MPWxx/ViHvOG9viea4DFUjwgfvSpbMlEcLbyIZ8vFe66n
UbOfl5jIivBRWBK33MIkHnOfr+uOSQBdup7jpejmzem+FITDNaa4h4Snhus/jOPg
qRHTrEB9j9cI7Q4eCRbsr6khf3jFzPZtBPZf7Ulx4MqZ5nzM9cyhdw4G1jYbzB9u
6VMW85x0HIYocuSG3xhRYgc6bHf0xn5MJ0d7mOENpJpTI7O617IZ/XFXW6XimPA5
YTIrQLVk+STDqqqjC3GNOgYXTUeqxbmq1JmPwzNDeo8pFeEXbgzvTmLkiDuLAJoN
LCIPt/lk/N2YFp0s0JDfTngy3as1Nmdmu/rolHYdscGbqcROcV+by/SYqxzgeFYh
M8r7fa0B9SXOCua9hl1anlpVzsI3eNp6j7buuBo7ydLBdU4nVHFyxOOGaTfhW7Vd
iKmmIXkTS7SaXvC0mS0Q/4gRCTTzTV4y6q1ERlt2TzNUixGG77VcNqH3cdZBd4pU
RIQpvyxnYOIGiVK4o3X5tTa0UiqIfvZe4TNn9Q9fdP3qKK9WK2hGBR1LWNvwTqUn
EQ7eJ68tHDAmLmhIIaex4H7abeilGlHRaUHa6pgfT3AnLRXkdJf+BgfzGvg3A1d1
owcSeANi7F+kYWJRLbcQYYL0FE/4XdJeP8bjLBT+tVo9pwUo+gOJZJc7/r8BEOw8
dSruisT9+n1TWnouFEqPnezPutavVaOnKnc+WtHyW+QxVmRagqHI3rrrmnLbQNGB
HMQT0Sc5W+Pj0muMw2ogG9i22pwMsLoAC5VuOg6dd7bkjg9yLHTan+874gDgm+Ok
N3Sn3aHjXNmxht5Egx8rBSH4noL5zow0b7jpKbTrZKqoCfNtwRXt+7mx+oJwNyHQ
ucFQpLIzna2duxaKqUU+slEPEOCWf/SUWeABFoeB6K5pa1JVcE3bTa4VLbr9I3qi
zUoFZoNzxQnIYlZCUBCUJ09vfzqMCGpl1cMpobceltuEco0xihX7gTG0NsnspOmt
0FiHreNogecd7SrudlZjjIdm98fz1E1cwBoMt5JkKh+tpfOJ4KpoR72aw65605ri
P97ZRoVlwyecLakF2ame9nQQv2qzduEMopyg8jbMmRBHUj0YCayKYJPv6z0UHLwN
/2zGBkRGge/yOnKPHnOoG9D8tZJ8vGYgrn49uZ9njryyEDjv8P7f5X5JoPKmHyUy
8tk5EHbirRH0fCJgdUkD6/GohvwlXNiDV65DFnG94upl17IlYi7U51OveQQsGlfn
lCy+LUDjYFI8kiEcBq+2YPS6n7khfsDRw7D26UlBb0WwA44PSXM52+EdrU8nf6X6
fm+a6+ayQqvcZR1S9Hio6x75dcbl2jMdZgESho809fwreqycixTc8cN9KdzjJnL/
gBEszONy5OviW0XxTcNxWnLA35sIGGOw6BFSXQtSWD7zKuQDzhJ/1+LtypjLUTLa
vfQ/QNP7wBhd9TjVfnd20dYgHwht78uukkbqw6k8lwgJPQcD78cdiGA3Pqq+McZc
OYS7Tr09U+U60PV/6PHB1R+g3LEQJ5U5KSVhV9HNByO0CMDAY9VH4pZEaMp3a5sq
SB92x2rGMU9DHX47FJh2fx4vn9+g+X/5pRHuar6ZEta9AauHDdxJaDlUu/wtFt5d
gvkSJuINddt2/sU7D6hH3OrK3wj+0oaAzxoglHEaS0LymPIr6968xHP5fR1CLr51
3slFAXn2TTPdBJ92f5d45wCppd4GMWP/1U9wJQPUSnvH15dUbGsLoFatJMPcZchq
gDWauHnLJTiFcEYk+J4PiHwguDywljUNkjdo4lGnTJwzPXKUYrl3riHiVpAX5P0t
YWhii/sw/hv9X3VOtAwN40XUdXF/X2cHRiEPNdpYlLaM5mQ6BlXhjnauHeX/l1Mm
PLMpbPrvxgfW78wUmb6NYHJVvpzkK7cGWKBBwvpBC+NJhQcIPgQR0DUBByVx6+Cd
39jG3TyMzAfgfvj0/M/9/9ootMO704cGaGHTM81sFISNlP1dHf3FHonvNgUg1t0U
pv35fX1rYJa07f/AB/19+TnpeQybDYz0BJMgYSLmACtO0HezQdjLFUJBn5yUPfi8
c82WomkQU6jfLBs0eBm2PLjddvYzjjQFIbyZF6gG0r+0MEn1GyxOV3HO+QaoAoMh
3vYxtZT+Kb1ijGr5pE1K4dY/U2yhDXLQC4vvXlrq+AR9rrTbHY7Penu6VbPgrC03
sy7B7XbissHILm+OObURp/U4cI5aspYnFtofQ3LT1tYXGnPTUj/7Z9nln/v/qMQH
qTaOCs0bho/XVZGe5TY+FMaMh04i0Df9lD6lHuO555R+GWKLSEzMNasYXx4sxZI1
BwuqJYEviMyFf/TOihlZgd3ZItR3r8EOX/vCi0anXvsNAXSQbQZsfUQvg0lp03Dr
f57X+SuTAbwBG1iNmzvsFKc0hzG0/eW8Vmr43063BPfwbXRPYGvOym4MzmPDXo4+
vi7MDXMmkJJd3OQgneST+EhyUfY04WebZT43ZJF3DNHNdApELPNwVKiwb1visRxq
1iJBfCzu/51nwYdpL5ocmKCZ92abH5LFsCu7FKgH8CLL8/zJ6ABuYolQHf8rEy/f
lKxDYmx8roAVi1oNsHq33vW+PcJCV2rXDjUNyVOgM3Wgaiu+YO2YbvUj+1uoOLPc
IHWVGfsHu8Sb5bquoTiGCWVPimPBcuUoAeTjnwFfluPEjf3Dda3UTv4nrYqPsVag
Y0ro64grbFgguyNGw/30YdKBnC9R8OLu+5vUcCFc9Db/4l/LYG04sGjQxSZ8iAz+
AiGf4N5CvNTWfVD1z9bFI9U86txCK5ffKi3Q0Vwbhp8ltpdcR+E0VM8cdXMqco3p
r/yNENIKb3K2tN9yf48AFo6KW5zHMouwLfgNnEDiwgbxFvQ8w4xOk5J45wviotA1
l8qSR1ZKvMyU2VCJOAUFOd+Keh7zlTSfJuuY9lh3fVVUJxbyDdnoi9udg+8mUo8v
djlJQZub49kfp4bRJ1XLctnbKQPoIGoJl4GsZL4zU+F/JcldrFtEa4x8UDQP242l
H1WeeoU6V1T8gsFBPoRq++R3Kyz4GPm2F9OwZXQO/OWbQvqCpW8uWsB6aXhRcnS0
IOkepPBfDY0rRWwfyy88lvhs6ylCDYoh2M1yy+m83TCaJVPrQ5BfsagjqRV37Uy/
rcjrNngRVQrn7dyyYE58139ER0IdzsFl+16USPnhjKud5j+sSIuyCvcfo3jXcJKg
sSJHfo8t/ObISNzYL3Y7II6PHdDvM95t7nY6CiFe39U10gd61uXeqjPBChKhwGTz
MY29lhXwkNig/KbGX0ZkhMoDtW0mH3nTFDrkEE4DOZbck6bPYbfQ7IzVXhAdzini
NI3Uo1LPFfEgJ4ti0xBWZqx4+UOpZ6M5BE2bW7YbCQ4Zdr6XoXg/dP+uLdoLDZI/
VgzaR2KRNnmCfvR0i/lgl7HttC+QsZy6J3p6XLzAhuU/o3WogNxJalETShZ3zr33
CvY8vVY8CnROBzyJKhl1s1+kzoD7g0r/f2KRCgrgss3/HdZk7zYis8Ug/tEL6T0t
ADVscrT+95fUShMh+22IYN/RUHbf2iaBJmlfNVl6jyxLEceMp1nYXPcUyfbURxbX
yFZQ90oy8nARkHE/6we33RnNmvRFoseDsiqjgtaBHZGO6AH/RyQhml9nF1pW51jx
3pkNOH7Oe/33e59mhiMdYurqkRgT3UyqJxDhmC91yeKbfI0w2hVxu5p2CfAlyNT0
DIOhVgcbtfDFXkcRLUWHFVGRvh/sa5n3DRXP9/EcEz/H6J52JjZiinOaxwKToVOE
AWulSWk8t8bXV6J1oIqb3d6RVbw4J2OAIUUpXAbeYlykxmZ+ZYs2vDvClZlnNvRp
pFcZInDngVVESnpXy9f2jH/LibDzVEIt6cpNi6lQPEbGRhy0ISH7JWTDUy+B/UwU
nO58760kPjcLOjN9nevZwZI/2FRX00gAUHimWVxyWPVYWtukL9cuC7vr6qbX0lGt
O+I4WC2CZOY1hvbmXp8p3IslrUjZnlJWb5YnT2x/YBHflh/mdDs33KjsN4G1R07F
2xSO8ggxMudYZKV4/W08PQeBg8kG9qVfMbhhsAgKwjcLcHCTUovNl3ytDE6nuzrk
j99yjj9aYtNuHlS74wvYLfbuU0l6ZlxEeoLCnYy1lU43SK4kFZ5Fm2pk1C15y/pU
1Ew+P6q14+zp708Gn4vdX83rA3IyPlNWtnxmcPzYOi00Bk9r8gK89AODa3/WoZfj
hw7Ys1dUG3TFKk5zO6ST770pie6le8oIFu3GsGiJOzjGZxCwcz/yR2XeGOp8jT96
I8DSa8l3pQNFITFcDK73JigCzyLxIPhb7BnkoO9S6yP8L1vdG3l+edzYc/CzArt2
/m0oxWKKhMjbHuncrnyTMcs3m6VgMZ5QHIzkWQvPPkxxAfbEZovkNxCIQzIIwC8R
6t4IHYlZXGU+ZWPcbikLmeFjYW0fiYYqJqIQmaotF6XZK+W95sVpzqt/iWxvtkH/
tUzL9MdM4SdRXWonzYmUe7wlAE8s+BUdpCVENmG0FkPzkBGh8XSVxjXqmDm+Rj37
C6AjsKo8WiksXFKFabme0MBJqpXzTDzaDwN9dxzgnmVr4BiNZNeFl3PJQc0MBmkC
IrYWRoSsDFLgSdkYCLQaf0nocElRsQCwSNycNme7efpf62c2AnkHXv94TOwKoJ8Y
iRcesp6BAxc/iAZjtGNhvUzS0HAhlH+2JaiV9i5FhS7nleyw1rWGLvIe2MQ5kPI2
n0igErbAUOZDQR8S0gRcSyDwa+vxAljgMsowIpIcikGyZTIxzCKpUd1KLxe+PALs
3K7Jv9fBjsReFyNFlU8JWwDmN3/LPVVl+ZelaDCaeE1ET0lMXz7Rk9hXyymO8+ic
7s2GD7brCZe/9xfnmMziPYnMRv/HbBMXwAr6E56XVewCDtMlINRAdkcC21f6op2Y
C9EDfZ72FosafZe5O2+qcBqCmOK7pFdcTo8QLmMJqBycU4ajZMOZaCpKPldVI9r/
QeTi0Ah59rBcX1MPm4PLGeQtrLZqfrx1Twj4U1hIlDs067yFJNcuZHKGz1aw80+O
y1ZHNwv5P3H0MSkDuXlfHfrbVXy/mY7ywQR5wKnaNMZN/5g5+LLhCsSS7z29//sk
hf3jJ7FaMM+78xK2Vk3E3qtjfTPCvdDJK7dMvYxgocOxcEBcFA8nba1c+86vh59U
CkNohyeOYtqFEI+lCqoyY04mA5AXES015WgjUEvh2Pn006SOPQbL7FOxSA8HbJL1
sP12REMIVQVmSQM2ClXUCGis2vEiGZAf8zrWnZhVTp1psZyjfQSEcp5ykLq9qc8y
ioQM7nfI8kG/TfHJDqOrdoIgW+81hVhx41+b0b2nJqfpPqDkkBkHs2lGZIRaLO6r
Y/a+TFPwoaUB9Lrm7/HSCJs1TN6QEMZGydCkeyVJFS+JmMdJglUhjODglC+DHVHN
lfp0EYNw48Do0x4PPOMu7vrcL9/HZbW8rlA9q36+6w2U0IfpN8VhR76vd4MywY6v
pxLvdkrximLHTVpIE7kJgwjqqU0RQZ3bMoeKO/vBbybGvYnS0dqpqY6SBkR1Z8f/
54ZPC1PKYOPZ/NUyCvy7zENa2VdLS69sYnKuMzb62Kz0MPfIvcsVoTffnjWqLlsi
sZzPoo7sxY5jPx1ACO0uy4S4rvwnvIm8G5WY6q2HoV1Sx4dg/DO/mhsLGseEHc8U
20t8cwcRlqr9lc1i+aghyBAV7eKeMtsOJtnpVSPQ+FLG9Qsresa/vO5e3tb1stem
uz9gSqiORdixGa61MmYu93eyRy8/8a+g5sem7dk1nVVuEDyl+zbPR7Phh/rChPzl
WViehL/kV9abgslePjoMYUwtozP/v6mepKLg7rrNpa0olQIxfR1Wt4Pc294U9hAD
1IOswHE8PgPCMvnA9JN0IWSGwE/lnxgL7pou651bwmRN8eVqF0cll0yp3GJ7iJTG
ag97FNk8se8ug/bMnxDXp7lZbw7RFB5ImTiM2wPoeQP6KbPxCfcKq+iLmro4sE6S
fZ1Es3TRMy3EsBxcC9d7xxROWI0im8TKRJVIgIIKtj5Jm7I7vdgrjz4yUDglfNdm
OjClDWrMCnJlVL68Z4cLSswOzqZe3IiVtTn4PfwXKKjDcCH0o36iiVeDRlrUXeE+
3PS6+xCvZl38NycdclZIj/a1bUM0rH9HM2MDOVSWap6IbftBd5+kLF0FKECdtfuE
ud+ayHOLvMxEjyaepjZ0zn9nsVwJYm4aEMFzvUU1g3tzF11uo290PNcbYqqV617I
CBpF5cE6tl0dQth57mFulpSDeZ7DMii09s2iTcoOLf1QUYczO4w9OkV6njr4tScV
jkfGJfasxaTC4OP6vZv4yABlkL9QU30ZljQZPD7J+/G/OCQqM8VzSqvUapq8p0OW
eMBZSISQPaOcS6R9kHEywCVynh3mQ17ZNdCPZMzz5mQ0FRSDpU/QvTpCzC9PWT+/
bOulHOwkwIBfSDNX9L6nWh0Sr+DeUvlmInUJM162MD26jbnawDlyz19yjxvYpXIs
FJUex3H4RBH1Oz0H9V+5bROnEvOUgsn4wIk23+rszfiMiUDVvAgV0hyd9N+bEDIw
7KUOqDdejjxbMuBt7PV5g/5yk32aTxGHY7uzlIx9GF3zI1ei9iOHL8xgnWlp9YOM
l5iG2MMw3l34wRgWxyqjgpGawz69Lj6sz1RnSU75YNduaretta5hIx5tsn/qp4W7
nacx5Zt4NQO+yOKE4YvY28ZAfpXgrXNBO1Thxe4HoYPvD03BPqrjajSRFJ3MuZKB
GGMTF039Muvs5c6mt/g/HJX0m+VcbPO8ZwatxG8eyBlJts+It2Q5qc2oM0pP8ENE
I3qqYxznLGhKOuV4c6pPTgF3n6miGko9BimqrfJHyokrhi5yMLCBnoTwPfX4An6R
FevLtsXpmCrJeQCE9fzKr+5QweQdK63D224r7J1yttIM5o6jjpCpoqVJSghs6uOv
5L6ju0q8nTVlGahsv+bzIL85BGNlqx/tj/wH3ii1LaHNUCUs4efPlVKzWlqRQaid
aR41LdwSxTa3CsWhGlrouugcPpTjZh60UHEh6hjxi815frbiLdf+vQA6idNc9LKv
SRhEBo5ZcjSFCOLXzyNxZevxaeqN1GrFlITxcktWW59Eb/FkCk9BsBFJ2CLpr6jK
I0DKTx1gzNIGWBSxmp0c3Oay68hsAFe1HW9zFptHIIf5Xiyl9qjyjCq1NMPPf+QK
xxVHarvkWCAD8AsVkcxSJBP0a+jYgUCbj2mJWyzjFGcapoa8P+ViAyQk6DKwdgw0
gfsda130cCIy0lJNHyz4KpUNM+TuCCmqUWVgtY3wuiIADHJMHAKQPMwd/ppI33h+
vasrttVonomdO1EZ+7ghyi4QRAoG9Uy7qR3c0YGlahxyVsjs0R2gd226knJyrxkF
LKg5snJsWBriYbLGpYKvZ1ev8Fn+aYWo9i42ZfvQHWYvjPyKUIxsxBAmfCTnKBcs
ulw913CFqpYlul3C+aOrgWk0rtZI2JffltFX0XI7bHbWgRt5eWOGFvZuRfjH12k+
H2NLOJ2+fbM3gaHOaRdecK8nt6WmEmim7UGGjcjroe9IT7hy19EA3SbV+j3idN4T
ok+g962AgfHVt41Sqt5mrvpn9VWZTNtTDElYr0Q2sV7Hb/tZ9I0gTRXVcFwF0iOU
9gFSoDUygcMpbM+xBbcbZM+uYxHeW8zIGgtwsme5fRVTygqDfTzb800vmc1T00JT
8TSD5t38C1xPiLkw+pNECuvvg3vTLh40k6ZlsKE+rJO9RGkIJeaH4aS8+UkPMrV3
USme9o1/XdZUQQs7d3WC+agHsF2Jx+vxVD4iI32l+bgmjIoLRbl/P4qQK1uW7+6t
LKqPqYdfJgCdloSYnB5hwac9cJR5MctOyHYYg+/oWP1PDGuhkoMTmmYRFeIx+gGu
nXJgcVrzuT2qSQ0zUqfdVVQlh3ElXHTEO6Fwmk/aP6/ErMFh/PzIPDujbJB2VQvQ
O3NvRLyhFY78qbj4aOyphAbaX4EmQhqfA2+cavCbgZtCjT6uoS5Qf8E0SpAJoWPf
8kb7+xo5XtlBhGWlvHJjBkBI9RbvbVhAzg2wbyGoYUnFxbZEpYbluaSTYcub6Ycu
Up6/TpkM/f5Ddr9WyMByGCcJ7RyjTZvw53Oa1ChnojTISL4SEu9HzlTMJHomn4bL
6cy8U5S1w6KsFdCoK3GLuFQzw9PFAFd0jO9A/Tp9o/wO6HV1sEj9QQ3JfI4PZWuF
KM7oOa/uYKIm6tHYxwsK+UvPFEcR0t1lfq0gm8TKqj5ZnS6F6N4iCgtkbZ3l+PVh
raAJTb5bgokLBovyKOk2zG+XpwPOMutPfhTto3c8cRuZtCsq+FDxRnTI1n5ZiBt1
QjCP8mHJw36pX2Q66jsY3sPB3otUb5k42docq0x3bfbfuHqsQJ2tuJgRnJrnci72
1Im7+4TZ29K0ToBD5wGJGfedv7Ah6CeZWxrcFKxf8NyUKVaI/HT7O8yJNP2whdZE
rHPto72dZQDzdBIHB8+Y1PCXHrKn4y8OpdX6u3dok6l5PcmNwjIF+MShlC+fP4qN
tKYt7Mj+joqE6jAGeD6tHayopwJQ9kaS3EUexvho5womRTyF4IPvuBZkuEnfCp2f
7ro7Ca9F47lTG3rnzq82L9BbkkpnFsebxi+g2tNR5PmyZ1tdTiXsvF1RNcqoWyOM
0NZue+NQzPZQuiR4o/Xfn/M6eWAtkaHq9bBhk0UL27G5y0UY9to8z/m4z0chpSxq
XYMe07mdMRxzX0ULJk52s5Z0Nob0lSjHhE2Y01G6HU1WmzAU/iThn1DO1nK4R2Em
TP44kjkkxtRXcczabSYFR65tRG6AdCms+ky1/HxsJ0zO+yVw0VTV5NEzWH1ubzyD
AXsgydWExYQZuCrnMvnfRjQOuvWgoiA1ZKsX4Lcm1zokc08OT5NfiG+aON80ZH3y
1aKgtKCWMcxDx4VxqYKbtXvL1VJXCmIRAEvNz0o3BBGeQaAHzSSqOSvIqW082UqO
I9pCnyUxL3I4gx72lvB4ZIfe08gWzRQ5X3P9zKH3m5rKhD4b8Wf/kIg5D5nzs4Ad
9mC5+yT3Rv9ssKi5X8Q/n6luE8FgkIM04p9yZLinkeZimgDunhDxg4sA3IECo6+c
WLS1/a+qZBvhooO8Ops8kIcQWiJdcBx/zzMJrX5t7RxAwgWfbdHRkHw4G9S7Rj2Q
lXHOvoiKcwhZ98KmwEvqTx5AdK+SNn1vhtE9gJymXO1ALgF2ZNzDz3G4cZYN8Izz
2vSdTAtsZd1JPf0iyIW1hiRgN1snCTOFtolj4/B0P+C44rg5Z3rWywZ1Y+SSE90d
iA/nq5gQhKOiBlh8Qk+IdWHH+eOB9lPpLyYXOkj8SH8SQUSVtyj4rJ5ki+J4Cvs/
PEmHWOwzhYivz+iXH39p9TWCIkfykh6fWOsLm7+gyvRG5u8lckArK809bBt61mu/
UheDVMzXIbGDawFR00hlARYoUlW1XwmtzRov5eCym2VI0QAoMMikaVii1fAq8WrV
CXuAi2tKu3ExaKR9Lx39hgAlW6jLMaYuEmK8bTuXzECHgy6Yvvr1PQ4lu0hM2pQt
s2G8oQHyXNvIv/hF2sQOFU1Pj6FXj1HZ1JFeGAW2Cb+Blv73Ej160wQ2jNPC2pko
64C30hQcGBoMOvawmuzT5AXq5mj27J0Dxhy4bUoIuazPU7Zb47mQnVJnbDWovMyf
g9Y+gx29K8ojo2RM6sIhOE8AQJcUk1PcQGkKg6h8zLs0yZtCZOrD5oi5E+AsledY
yZTNALkdc2sNzWMn2Uh+9EgG+nuGkxW2HnJocReZT/wfKmv8rvNxfqukNuruOptV
QN5ARQYQ4lSN594AERG+a2BtZkLSBYE+PNAzA9apxhUsPot7HncXl4vPXn3y8T+s
n22tm6uVJ5z7FxTFeSscMTaAtVrwBWNQgi+LY+EOb5gvi95fKMpx7vkpf4bNAPOe
/GYY11JttPOTeO1hUlSWeQeIV6MaTepcF58jFUyh4EQoQhYMLUYdKqpBozNVvR5T
ZD070fgXLB5YEetitPZEil6f1Dm37OPuT+DUeNxhLIpn/R3MH1k1vIBFfcfMlQat
wVreigbxFDCR3CVuZxYgAXsxTHSNO79TeYM4+dIi+J9UXU0ht6ssBDkdoAnRkccP
4RFXBKgRuTNRp5zMqyYL8B/3AKdAmzakr8GdkFZWKym4zHP/RTPx8FblTK9gBOnZ
XPo1UceQaCIzfFR9FFVhx8sKg+75vqEcNG5FV0xa1bjtmNpb/Uixif/pLLJWvGwr
EJSQnagWADOUf1GqrNCFqmK6Qb8pXVnibhI5+nqmCdsn/BjbQBLtAYIDhRA+4u0a
zvYa9jxOvgduj/uAnE1sLWw6HGq78BaGF6E7pX4fXkQkWFPGtS0ZlyL/N0Gr+09A
iu7ZUUPzAB85ONx6/UVjjeax3eVM6hfPCz2crrYTxl2Y2o4stE+jbDoB/CTBB9BL
eI9W26UMss+SGHw5JLC2COQRYu8Dgx8YghtIDMGigbBr39aGPWuPR1p5BByyQFu9
IZltAKdnI8MloYjeQD4qtOr+PVBJhNbHxGHTo4gp2wHKQMVwYIvAoBS/K1HmAXZ1
sA88o9iVnbCgG/EmhJddzeKwd9jxVh4kBybW+LNPPiWlSYjSl9u7R8HyIhktQST/
Zhv4gAUbZnAMSMuDYKjabjlgSCuUYcLnX1KV3z+NhRDZeFHIcc15gZMO416JZRTV
3f7zH3Fc6pvehuQ1Qwnwn55YMc0T4rP2QJYuQc5T+78e6PAX44mI+airPoLpb492
vef+gvatIKyc0YQ6u1anxQxHwFNXPmbRO1eZ9WOxseWsFTAkPODJ7Kc/Noeitxz/
swT5stK07/G9mEdJe3huDblVcUpnkqknWPX3UzoYHrRvgkCHxhDUN5pY5nlEuR8z
4HmsbtkU00td1fc5Qzxclwsn6dEy02kQBvIo7UOfe6vCXW7R/1eRJ1R2hh8DV6jN
xLulV0QxXByPRCuL/aNIvLmmz0cUKi5thG5pGMefXRWy68euqnJPmCG4pKnK6iHb
sqmSQ+8hM4gnCTsdhw+mVvdtbQPD0xOHYnXRfZzvd/ZPWqpp7+BbNFYYUuGnzo60
z2ysun/WL0jUfzYGqb9nf1VlP5g4ErS3C7jPUQT15I+ZIpyPwFVvOZ/Wf84TxZk4
Jn3/xmy3+At41lJL3GXpR0T87x4FdHkMZbPhVBKQhoWPxIa15pKWnoPbHNBQBdhd
cVE17CVEkmV6MgVz/Ia6srRAxtZH3y7e5djqqj13s+z3CAytLsCCbBNNisfmNyBR
yN2kORuVd7Xxfg5OH/zqnyHQmlYGs4A7altqKqNpkkZebw9g9A6ivUVFieYZXjdb
djZd7F7SJY76uT7JkcX0Ym7nBDEhglRVUGpXIQ2DECuEN1a6BJYAlGsCB6UBphHV
ahnMMPaon3htpzObARXv9m2BZYZrgmuipr93ikXjUKHUj1Wyh8bETr2WSVaYCz3y
UobD9mK2byGXzOw0dKJ9AIf58xMlJZFgRVt+++RMNsfHyiVc+bjmu2XhTYgGjChY
HuzJN5x82sD7/E/Sa7K0w/ppSlmWOmbBnw00HLG7oxGqb9vKqzdXZi97Lw0OQfVg
z47n2yhWsnkqgamm3tbWNHLdFlEVo4Ue+sQOGuuJLW+4NPPoHWbX2c6tNqVtzDZv
Nqju7s/9TFPIoSkit/mnt98RxXeMQooAhFqrD3opQsQZKuQ3TmzgPkEmrE8726dN
Y1uq41BkMNlq2QXx11bC5ovw8aUgWEmRAFZwBtgHtn2ug1zTcRXZXBSpMn6Rp/tM
jHPwuhLNOa93zyzjAn9MyYQ6Fn+jNbWvCOGITtHSwrZ5gXwxVkU9naoB4DSeaCeZ
uFvuZEDj/irJYanuy5OFJFfWCmzKt5xV8sKfilfciciYzgNtjjXEuVWAf90R9F97
pRqusX52BAHbWbj0wWgtohS35Ct8Z9RBXvYT3u2t89tLUfaKumCZdqcYPJXXtQyS
hdv7XYI40vXaxF7s2ay/jZkbKpjvp0s2lLOCOmcOtbrgvKTHPfCNnvBC1Wr02WJG
8YB7HR44ATopY2poO6su0jXaZHgfFQWqP2NNs1wayorMCzpSCiWeF8XBldX0CgM5
FadDlwPuqOkh8kEFLQ8Q00v+HASIQH6WkGzPXMm2F06ZeTRJzoAwzUIw7HgRxBJE
ZSHAU+lMzR0bj2jgRvdBocNVDQyD4DVnEubiRpX25v6eqm8Z2IqYMQ8b0qhdLj9L
QF5X+E95CPuLPBopuRhXAnAVVfXT/0HQUNpQcAULbpKxF7E8u2DJOn2jMBCzN4mb
STHKM6VkhHDKnGuBEixQ+cwfuvxfGm/tQOTE5+ICS2f/rMf0bD6GxDQcemlHviit
lH8g9NeupclPHIK2ttdW948HpQsGiisOJsLL1jTN6FUNnNA4Bn/RVEZwKJd73Jf3
mC51Ab31/xfxPaPYCwcexGBinwOZcvLnWBrj7G4aWLFO2gRjJ3Ts5hoeZgJ+RZUz
C2tm2EQHJq3TCsh4T6NzEr74KP8NxU2qSjpW9OeJ+AsLVKxDcj9H3+SlEf2yZWqT
klvEnzMMThUZeurPFdKzPkJaB2BrhXm1VrL4rH1iAOgJy3Tmtc4gL7IuVAthWqKN
kYvFyMyAf5e8zMCOVZ1jVMIR3F0aEL7g1l52GZzWZaM5SgATM1X/ZHjMQ0hfSbXg
8I68Aft05AixDmWbm9F9ND0b85j6dKCVU/LnXdB8bqkAK/F46V0xbYqKfHYQ5Y5Y
iSyflZk8ZRCJuQw5JQQ3rRzqu/f/xVzD/M8/1Y5FCiIhM8pdgWtBG15QWk+zJVdp
yWXw94oICa5lIgEichqdF5ztO2NL+pzQ9qkYDMaD9weYcy7QCx4avOVsE/7R+e46
kBnY/pQ7C5qezs0rvVNFq6owK/2pT9WZoqdDi7nls104UuK3Q0P6EkDEBtZhKQ1a
Ia2hAX89kk8Pni3ChAt0WAQ7tCc2OQiTpUi1gbEEzQN8iDOIJpC2EoJUdnwEcsWr
5pFIWOaRq62/S5EnPXkcJabUzpURVOqhH2m/0QzqkQ98wPwyQB27gLbgnUs+IJAt
5S2vWruIgQEo+10XHhodm1oKjOiUGYSwmMr6pUX6vLzbtQ9jnhZOMSGV8XV33dqz
6fNikIh1lBbEd8fE0L8qpO4mb5N3+XQiFfAT3uo1Qoruu2f1ap0rcZ/hIdjZtUeR
LN53CmVTdw9GlQ9ILPzAl6VhOnjGN24jQnMw71T/gKo4s97TJe27P2oWK6EcUSmH
TaPWfYwB+lLz6l/9BgFcRPHbAp7Y3ek4TdwnD1Dr4qmd/pqDbH05WC5rHFm/OUl7
e3IkklJgzIvkBeWqN4CGv+qtvg7r0ax9PlxThmYpqWnb6SieUla7JztvokhLm+aJ
2WmoOfn3mVr9UzFqrVzF+mnos5vrxrdiusr5YH0d1YqNEc2KnOpFdQBzY6t9MGQm
/ger8mqQFEHWXzwYUgpUcFGZUrntZ/CDiw1h/x+fA+PDpG416x4ghaMthB64lkO7
RLgAEs6B4ya4hD0R0+R3moO7HVZV1fog9LxrwERkw4PFIL8VF3XZY+WAkzb31epH
k3D6B4YVjVwr81qyuSFHoTPfxfEY1XsC6UqkNw8mn9KLim+pZN+d6gbonVPJ/Vrj
LcmNjM9kEYJRKKTFq5jWqj1ohNhxiqDevPxTzXHgbSnjBhJG9+5X5i7urGmp37lT
5AAmVXKyCcFbphzgi6jX7X4ib1blBfmpflx+Fswpded7l6RlSelelKRChhtbgkPF
pBQXjjmri5qQLw9KnLZpo3GZ9w64H9uLXHbsByYsKhC0KXGbnIujEO96ejxMNTGm
iasPbwQ2EEdV9nzvMehmUXT6ERAzvRQ4cK5g7DPXpF+rbh9tfLRLileXslOXGFAZ
9/OdhBoJ5RwA8O7Q95cL5UcPXkvVm9KJqkgHY7TphfenchOOGQfExxv60TQccnvZ
OYdWeiQZ8uZItRMkiRrSH/3B2cuAvPErY3VgTk88gSVY+1h4wS4NuEPGDCGOYK4+
UiW6sF7s+VmjePDh8u0bLTq1QmKzQEyQrf8R+2tlqhuT+e2fMsLHXrET31Y4OBe1
CT2N41hUeNG8nlnW+g9wNPbDSJKQ3f+vggcePOQjh6xuQX/9Z+to8MNTPMN57yL1
GarJFtM9J+0hsFyDTzi4XzpaDgv0YbCOrDRv+19x4Vr0c6I3JmoxL7DQbt4aWwbG
bYMaTUKSTfU61JMWemobjgqVroGAUbschc1rBCcQw05BC9fheSEJePoRE88Dv6Df
L5ZTaVSQFhEW4yqjDHHvFpeSbeMDTmfkLc/UVcdXhJqirZRGj142gRX5HEqpFF/5
27TcMRKLbWQoCo4ybKbtaft4Y91CSL4Ou4uBTFGg24cDoZ5FL54pBO5Q8M8J+jvv
rZgGAX4fq6oxL9537NoAAPhAyw1EaJcTdyVDAA6FawRh8gqhXmdX2GwRJn9kZ/Bo
5sq2/y5iohcxACWef8R4BmraQ9Vn34G9S9QnlP6eyShW/0gY7NMtdZxLC8My+S28
tkkpXTm85j5MYm1a7xfKS2vD1NFWwDKpv5uX76F/LhG2TqI5IvoAEU1BJpi1/z/m
6DYLdULYmuucc11XYmMx0P4B0/HASsfrWELJDvwfqIZ8b/svBTJ4gX9OvgwZgf9S
NatdQU63WNNiDBpjwfgwcQKo53T6/bjXro7Rk8aHVjq/PQnPQzADIYw/CNdYI9NQ
oUUfzYVQXLniY2GPpSuGcq2jUsNdYDjvgehrl6d7vnwIvnmSzuQhLBO1SNlelJw0
gXyCWUy7zNLkz8dr4Pu0mYcM7ErZzE796Tg/hCsPN8WsziX+pE/DyLC7/lrtvSuK
NdQAk+SFtOoR7Dskro8vV2AAkIiwc99a8QWPNpD9XDmLhwAAbHsjv4xLMxaaH4hX
h6cCDtMdL3bDKL/54QQoSz+0eZnSbYrBE/VwspowQKaPU8dw3jKPxikLel3oYt8t
nUDnbMI72S4rHTOvu2i/HvWlcN2fiZbUyPm7Y5fj8yXXrLMPJcpXs6sMMojxqPTq
3NHgdJyNeNxNZJ1QJmp4KXx99/g/C0oded/Kt/Mvu4n2lxa5fIx6zpMMnBSZfibk
hmuIHNeVgFpO4H+NSn92E5XbwMHkM7FeQ1pPvkYiNidonT3KCyyxB830BVVcKOv+
XDbNmiUUugAGVeDIBfbanT2qC0q1MLx8Icsrs8DXKbqv4RrcB4danLQp49csmxW/
BGVJG945CWoVvbSxHVqGFgAKZVEZvZY8R5ICs2Qt0GYnZsSP/AKVj9G1HUV2qP2h
ypLD2PiK2BJyhBs0TqR5A6jpHxssPljrwjY7YdYqxKnyZjTJmKZW3NWnTygUsXhK
tq8oUoIkOcuL5t9aVckYgcNkAqPVSgIWeLYagw03RevVHSGQmktjEYjTceyxH77/
W5uGX50yllGgiZsFH4EFMPWjDt5w0CPosB9+3WEVWj2/9j43ot9x5cVAuhHgTcHz
T1RNK+9ZDUb8eOc+T7MqdwTbUD5BrQ3XTpqPJOhPD2HiZ0/Cp3r1cftQ0j1pZ4I9
wlArZC+mP1izwmVGXR6tePdR8Uyv47eiIddQT9Am8mrHq6XQbSDD/HfGbHALgb4b
oEo+TWiJidwaIwlpd2glneGIJxudVuUw5iHVrydggUWs6nWMyQzJzi/iz+kwAALs
aXc9HMXS4F//T/nz4GbSfwr9hjcUO4w1a3QjtyqV973mbwWNg7LBNR6SF2nVWQJx
s8WPFonQSI+BvoDWunfjPgeHTUwapYbUxjlHMElLgJDCmN8v1NO+/fpeFo4bgX4P
55plLuaLKvWsAQUv42yFW9buzaOiuT7z5jHAs0yO0vc0JQ0fldFqrO1F3N88DEm9
YQd4SkuIahdeAXLJxczfej/Md840sY2O3KXPyVCxML/rb8L1IjawCo97XrKksMt5
qKQ4BdjdjnRCbgPRJa6wEK9hAIe/EDMiwGfP9A3wJhcUR8OeNvPgV7zbgM4Rsrtx
GgXbgfFv3i+Uj7hQ9PLYZC1cOkQ5ftCGdXKXmdtwWJ8E5dBVV55gkUIbSbnX56Wy
CAO2XxusSntE4GWS7eky7KakRxFVkJ0iDJ/htMkmxzrv+Z7dbjP2zfPADhn4/o99
Y3J1qI8oZ7lrTMrhO5Ewzo86zjq/7Ma0TOUAR4nNpLvOm4Eqoact5l4wzhhZrXVP
fDfLdKGRGoA/VENap28BHDFNmtTqg9ZJkr61g1qiQ58UjCCwINB1GeMW0IOUbYTn
7/nqJ0Esl1M0r/XhJuOwSu5DcCGx9SKH20dEVnWa++w/VcS7nRxOr765n/WR9Di0
vtIreTCK0jAnkn2j8rQg6Id0sp5ZIYLtncKAh8kehaohfox0Gm5frzzNpn/J+yGb
KhP4LNDW/TFxKjI8jzgrLGU2lzthStx7hJp8eheMq9404NkVUT7r6vqLaNGvxwoh
yLyMKduYttmfTg4Mw6JlSqtOgqtxOJwcEejP7XqBJcdKa2vgR0L1pTv/DsbJKjll
pgO5kidv+wdTjVXCA/XZ3oJfAug+rgU/679peOyY1GWZh1zsoFscTXFu6Y2UH40Q
lk3ohnTWsOzSctVGRu89DINk1g6VsPthhAV8u/AJKW2u1lSgKz7iXVVAdlIa2K5k
hcJWUNLf0D+TQBLYiv8JRNBDu8k23OkufvqWu2OpVaQHcU3YsSbxIy+F6p+NJUlk
A+79sHvUyNipSj+blgEHt+h6+QtmkQcvTpu7Gf5nczFm54xfW2WQOKsohXDMF+23
3A8i6WHwjvBN9mQZJ60bsBFxzrG4ftX20JuD33N2jO7BBhiPbA0jXz+PFRXpgWPB
zd/KoQaTPKo/QcrypjGBkRenMGWA80LYrXoiLPZYOtaNFXXN2fDeCaA+nLQVSlS0
Dle81y22gYrxVpy88kM6KMdJy4Ndhy6bXW2fnrX8RZHIuLf5jhd5RazZlHgeOd8m
23PCr/KUgg2S9S7LDg0MieH5qonDTBDyXMJEzUpsiie9wA6Aar0nHqVeCQK1xvuj
hJ9TB/8jemvbzTmMq0lOuKEoGJRL1IwDXLLhCcI4fyFpyCvdLokaBMkvhAR+rMBs
XXKpJbScUAg4xt2iMsJBBxtiSwfHUbRmcJeFg/whtLPHDb5g7634h5DvKf5sYc2N
JQHx7xasDM/XyCqF3gJYvSByCuGwteMz3mkJkV40M9mlRBM6qrnQgAGmj2tohW+N
EGAVvgvq0iBhpzG49og6Idb4+GZAZ4BqRqX/hLUeK23RI/11lM0nbeGPkIKYNnrQ
77CzkzAvztKPQ3XxQJskhA8klV096J06G8+umyMZ4jqjGpgGmGDnrwNj4R8OD71H
YMmS/eYNLh0EU0/Jy+gTYzmm50vnvCmFirhm7nR+M0tfTsKS2yYKuaNnCkXbUX84
/98nh2wb6go/wuxWQhgXjFBVqLQ/rsNdglQnD2uZL4chlez6XwntlQsMXZkEtV4d
OYI1Oeg3Cz5eKEcGarJVIoBuYLwsE9307LFfoq7JO+vTMGcmqyMcO+54jQZ9XT02
O+8JgoJBo3PMyhWM5mGkF4RfDOR6qBoDdd4tNZjk/N6nPKinZFo+nvPXZJ7BfMgn
revNeqfTatAkUFD+2CTYLk3HUMs7zyBa3wsEDNSsjuIkhsWEv3M0FdUrzHLyu6UN
UfrYf0CayqF9JH/oMIhA3gfPm0sdkR8cALcBlY/IkhoeyTCXmg+uA9NTfsb5FirY
PKfPrvizxHxhApAWaPeQcEnbXFhGO9QXUZZTaZankUg8Yqu82ngmih0eugffHIpL
dB2nCS53vkrNxjjpbL6AXT5lotw2+yGRL+DKuDzaL3qB0AXY44VuDDjLCZs0LDEQ
9m7OVEdbpgw8Xwu4pLg6F92gR0Jh8fyEdTkiTHYpgDznoOnqIoHQUPTBiI+UL6Vv
vRSEb2MuDrWbwmKj1w6Rl4NP2h0/XIU+F6x8Z5mpscgFqcdH6RCPEO4928g0C70K
NyFsq0GHCDqfDflzgxWtoxQ8TnlDXSschBMSSSMdKqh/5TUCDN6VZUPKvuCq7rOG
CbBMgCiCRCarGXWD6BbvmBCJ4HNCIeT/rxbvBIQZmBTNaYeS9xa4Lx2cRU/ZSZV5
lg8Aynilg6ESUFLiPSy0PvcB6kyKrOMEco8xKax9WQCJo/mZScM/Y/cePKU/lGaa
KLiclljFNvHoK4np1ataHWHZEBKMb7fFP+esJ6S3HBqJBuTn8hsbnweoiI3RxXts
eBshtPvVY0p9kktOA9eqrYkPxoCisU+gf1KLMp4eX0JVORl2FuoRm1y8Q8fNEZnI
Qx6qrDcjl4Vcov7w31yX+PukU0boskpxaooqcOXf3SnAGRqIqUwV+myhb4O496DX
fhA/F68LWANy2JnAGDmYiXtnAMbY/TZlAsVAzXS9zJvgVHenTVzfs7DsH4d5R+qj
C61JUPaWhTJ7SutTZrvM6QO/aezQOJUZirFZJYKhkjAkWNjJ+jdH5Gqjv6DkLVMm
W+lyNJCwt+NLpyyOPdEVkbDvbTGQ4bjOVJxDg8UED8STWWgtAPlWLxbFuA4XGthk
mt+UkbXlel3yaUGwsP4/nqhcunYpX+HmnV+QD9DUyvfZjVzdBhozBHeHHgcgM3Lt
JSRVdDfN9UIv5W4V4ailQJcJ3d1V27/EZJZEAB/ApkpXp8trx0OXMAbs4ospLCRF
Ue3GJW5pHFbX+pisDJ6KgJpVHvVJ2K7Y1c43NrJKu0tMuf9qkWY+A8HDTCxPTBXb
sYbbRPDOOdQ8YY5Z7pgTjyd7rt7/zOhOzyS1k39ORgxk8kfTNk49YE8TcBk79g6Z
ixaxJBC3IKAV3PzVD9fNy+BD/zkOlCZV/Ba0gljnT1TvC889bPstPA+UuLPKzcQo
BAA+k+22rgIFPrA+ISenCVd0Y5hyH/pRcF/AaJ0M1n+PC1AkWGV+lbmDdSVWRgxL
2Z0byd3Qfztssc42fPl+c/xK3/SWBBxEsJlWiPbpsXyhvFvC9gWnGwFUe8ecZymU
U3mi2V5Mh5E8GHJaYx9+Oi9qbKbFqti/lREg4AddMIAEAu45dzahfiamIfWF2DTl
2snmc5jYrmC+W5kxeHVQ1oTKv4mz4Krk4Wnag62NKm6x7WCAT0JFy4rTNyoIzvMj
GkgJ1OeThULd+4+oNrUnDIrCiuVF3ZXxv/CFB2n9Ok0D929u11FvuCiZQqOqNrQN
kJ2BVTEfnUaFcxNipaG/TOIi4CdYi/BTfQkLV6x+ZFBvyy16GdZ5NY8p7BnBcA2D
QWcT8gdRvMUxe4VX9uC3gHLbpLCYL6xA2vtGIlG4TQQyu1zXfA9VZ3XEbvhwElay
IpE4bk2p8t2eMUeBn8ecbgbq8cs+TJVu5psAszAF8RpQo92bdlUEAaMhogshWmdV
bnzEg4gXurt4xpSEi3Hcj7Ms7RziyGF3xj9PncYs3Y0GUIfL2Z4jacoQeOk0H1HI
hQrKFdOXqVCvsg/irQaZl9v4B98HXW/CAmEPQ+cke4N4n23eeMzglRWnejTSIhhl
dzW6IaMtWVDb9b9z6vJ8nva7HBUFprxTp3ZVtaxRptLcLsatHFYv9xZa+4pOtTuB
2m0OlCoMua6kvZHpADfiezZRF1vaJF0MZ1K96JgFlpwyv49AWECbbCpp9aTj78bq
Tpg2E8l8KE/mnP3Q8pvoz2x4SY87h+kiNVT/UB8Fh6FSW2YY1Lo7VkGdue9GmnRc
dxUFAKh2XL0V5KytODaIhkEn71muKg3x0qaCy+gLNnnmzxcf7lAR+0415b2UL7gl
XWZw7kfLfK5hC7jldTQZeJjEKoCYfhG3nqJoalEz49zulIjPVLOYSXkxwGJFNonk
7SLNJxNdW5tB7J02k920m+RpDuC+xuI+ZMXu/1ymt5kt6b6i0V9FnvpE2du/m3fI
EpLrCiOQIKkbCmRumbwIeG9DXE1UlpVWPUQ19FlT3WLhFSZOx+M9IjLt6tEvZ7A9
RuqJwIdzwaFEbwyRm1Z+5wALxW5mUt0qLJgC96zZWXI706QDkCheof54SZ28Az1U
P8vXRPpeSYfV4nL+E49/RtbDORXXHRbvCmDzwhIAX5zNZQVnNh/ZlSsExXdE/xFi
2GrdpIIrHp6jveOHUrh2DrOOlJFRhLpczNkvekwH+7KtLg6XXId9NVYB8xPjN9dh
KKbCaOQ2NZJsc5iFp3if1/v8FJNhBKxjsSNczq1sGJqgyjBXtcsPXIArZ66uBqkz
L69+DnL8onvk6li6ZHIOLrYeUx6G5rKbEwMHOr3rDNF3lKPBIvGbgQIClyIER17m
MEYC22ttUKYZBG7ncggVUQKcn8lvTegqfNmnOVt6K/RwDBXA+7VSZXWhu+ZgQCwj
y8WcQoCvR2BLTIPm4Srgpn8R5uPCWADxFPLbv37HLT1A0HHp4CCjDyljiPlycVwu
t5ozEiHgwwyo4oEG4NeQrG/jcTdC7obsXIqo/TA8EOG9X7eid0U9V0HnqUCZkYKJ
v9JrReLtleus5gs/flZB1DQ5z5ZJpC1E0xh9X3PC9mEkpJX7fOHkztoB5EvgIMCp
yUuZ1mel+BX/HiZe3X9N2KTr16Sr7EYxNVZYQcSTA8c17l6Rp+8NjyjZWJs4ZWFx
wDDShF1ysRjPu7Vy9FkTgKTneYsSnvQHkeFF1FE5sUXfR78ZewsgpFwjpjGOBHzX
EcFCiPdKFsCNOk+QKvJZpyWFiIDUFHlcBxBlxq3POdJM1newcCpDJlNW83CZhXNq
h/ihPMjbzZoEILeXzkZ4cLHYuMw+AbxQxW2IGiatNaS0PpdYnfMHklFMhpgQWM8t
0qx1pNFQqdqr0Z/DWZQvGmHUTpVR6srwDWzLj+RUqfl/2YNvIcv7AT8YrQN7PQXE
VA5933nrOKmIjx0O/9ebZdA6MsQO+am+bTGVYNfWldxXEEVcMTtkMOFJnsHDS1n1
/jYFOeaywgbkzKvsgaljosjlTaznZuOc/U7iRnGwvMQ8sn7K+M96KYa4jWkle5CF
VJmFrAVJMAkQ4gFjjDqCYa8GAVzfE38YS48g2meIkRpzdSdqvB4FQsqC17OTEt1Y
2tFk/OvU1iJwjoHLp0msiDveds4Uz2lAcEUUQ0bu6xCQJO02Nv26TM67ytSBAMCF
Vw0xbsc3BmKoThd0ouXgPxHWZslzsrezAY07VrVxNcVZz4hYB0lkDXF2C1GyPLqD
rAlqlXQRNXUgA+JBOHwCUYzAyOXRvN63VvFeq5cDtFmXrNDtby09uJyJauT9tsy7
LkaqsUB3NbUbcvMurt4fsHY2DWkgSiT95rTMpNHC/0Lj9Kyu/NblpX7jJ6lqkR91
1ldQeCjC8EKoohxgiuXiAzl6/2664trpiXZx7JNU2tavnFN3iR//lFby4Y39jVHP
sTIhs4FPIzI6nPZM9Ro0xBHCaiRLplZocyMxqqfO/1+fSxyFgGk8s0/x4ZJeQ/43
xD1N4Qtj7Io4u8vRgYK8n8eUQkMdHVl1AtEqlCYWC+TfJKTkPCnUzUBJ3sqx9HM9
sK8tTn6FCersRTMnO52QcmTcKkiEQfEhC2E9MKy2ez/P5sZ/1BOkBc6OezdWFP23
O6jMdlv1vRhfOs9qRnr4GkoRvwjj7SbXJ93vuWhP7Gr6Oa6lltemyDc+SW9mmJ5+
4MubAeaRBQHOuoimegBOpRaHuaw7ihDdY7yJWpRYE/r5koTjtThLhvzyLkWaooJ0
vjahSBjdY0+M8ZuYKC2omGA93J8z0GUPz1lTRFtVwA+nA9VPg9XDQMdS8CiMJs9I
No6LQMjvvZgEdQb/vJs2VCiLis1xZndEwo908TQojmdK4pP4MYRi4mUK85XA9E5z
FyfZw6p2uQItBv/rb4LsbnEhti2R4tZYUQW7kdZYOQbV80q0h/Rj5Q1GH22FA9KQ
NuvAVuqVLpIXo/Kil/nZd4U6xEqFQFAPsiWmvYYp6Hu19zQveYehGNb8J+Fv5v/7
aH5i3rJlo2gMH7P1UHVjJzHXtx+SqKVTAYAi7lKGOIEHdsFUs+wZB23iOBArJJsc
wuul1fIBeSZOnUHoVtMunaJoBPZgisrT72bkW30A1rnBxlefLZoO4SZekj2QYhSX
jeF8afiSkUq3znPhoiWww4ai5c4KDOd1IYRA2aTVuJYquZvTMqfyXekYvq0nmLcN
C0pCe7tV2KVg+BVDKdDoEQbeCXsuQnRkQj2qnMYAIvagSrwj5/5y+mdtkzZP5P4P
BmqjrAwyW7EmoWyBTTbIW3jmTqGuGEx6Mwea/VPGd4yzXzUM0Hdn/f/uJ381WTIA
xXc2uX3pSscC8ykZnTaoFYHmMmzKXeuufb5E1I+cZfiF3rjh4YO12jlxXNAC6ttY
mlb3COn1yfh6o4LBbrlVNCLOx/KvQS1KH/fCH9+cD/rIQQQP9SJyYwwRUc2VPf57
IK7lj6HiAHb/lOAByZNBVepOqCVXn67HeVJnMag1MfEGa6RAQEC64QONQzQrzipS
tcjg2wSNLvKhPakPc8c5SVQd5ZCgjhMa1stzKeGCycRHs45IRGTvzfkBrgzEdZ9X
/x9Y0CPlFz5CEPn+dtsHcjYak63SCTZNyyQLCkVUamNw2n+9+ovvBxdBQwoNRwBw
5uZA5u+JgqxtHLPpltI5/KR9eeOK++2FkRC9g70Pk7pyJ9/u3aE7VJrpvJrKkiXG
O067BIndXP2TKr4kitX7yPsJiCe5iROBh+1JLLIZnQO78WTsKU4sDMABzYz5ZkN5
Y+0hsqx/wReVDAWME95w7oWBvs4sXEiV6+icsAQe2vNjqQDD/T90AheFlTr34z9S
u86PZIhL4Sbn8Gttr4hf48HmxHS/WuRB+nBhFhR9T7w1vFjqV75Tn6YlxsQIXyLq
QI4OPb4nqF8eZil+f0ymC9wpUq95oM5V2xOC2ysThxUzPKR8aE8kIgKqaK8K9CAn
s37azJ8GZtjdZUsHA0EDVsyNeEi0r6k9PjvIRE87i1UvFpxGowZSjjRFXCq9ddoX
eOSokWTGkVFHgOF2Xk/NNnHkZOWflxS89SDEaL6nrg1pi4B+Np1K+MSGyRuC5EJs
QcPBxAG8EaAtdJBktkdcGl1xlbNajjqM79f7HbbeBxAMvAcT9DPWwJKuUM97dVJp
tkhrwZ/cEFM4Gcsi8JtjnueWh7LMdhVuY2NKVo+4X/XsMqZFr8rgeuyxf8ZdQRkT
zYHMKE63UWb7P1kQLzSSLz762Fqxp9MVFtWW9kSfUqIMwI2ftROHUHUTO437BRXR
DiUomtdaQQXOST/dYnoD8P44gTTri8xevfbHZBTkDs6i05Gmo6+DmaMTr2g77G6D
kOhPSlLqP1p/MRwkKf2/jI0vqqHaiFnhCA3DzfWNECAyxIKQ41dcxfuO0Y4xmZDq
g/fGmPliGvqY2KbZzuyOis5foVe8i4M+qB1prouNrnI7AbyZQ2ZWl0dW0BufqZLh
mNB4d06JHK5Sm4SC32dJqfXYVGoYAycGeSDUDw5RqYn56TAMUKmlbtCwL2pebRfk
WRyCThhWLem2VZ7CsWV+1qSVIzGgYWn3iNmvgDaAoD7bnjCBGKmGedpGXTkmkgh2
Euu5w3J9iTViCYijHbItPSZdBKOa1Bc0dHR7DLadG2Dtssd0FQvlcYaMW2Thi7iv
eWEPbumtDfbwSVwZOrLUpb/ZU4Y9+EXVv+QmS7LF3VygxmTRlHLSXKzsuTq6VSKy
avby+vvDCbbOW2MFs4AQKkayuk0YSzAmD6ZtuQIb6bJ7ur6irYuWkA8aHB1ruRfj
uGpWkEd9Jrzo3wDB69pgMj15R+Pi8DVs/7F3VwADWMbQEPSJnEjwrKcaeD24acwc
AJdDC2ZeNik2o5NmEdC0aiERMVXxsIfxVskuDAUvl+ADYwAGacEPiQ9az5qMMHQ4
GQ3NDgCBJeXUrQy/1Ho8tHuAub953NKF22QGi+0w8IkxUqef4GQ+NsKJomupBnvP
3d23RSNjdgT1XSo/LBKdJS2G+o6TOxwCG1gxl0OnpRe8zABum8NNlj2BIzh74GOj
k9xzrWyFmkPj/AKqAhu5KPvJfEvtJESX8PVjVL+SiMWzSdXOkFHaEZVjuLYeCZt5
nVOj9Mp6RTmUVo22TJ2KchwJyk/rFLr1tQnTAowcQi6GciNwSBQwpNxJE7Vur5nM
mnfIwRyQybupbCb/LmyxEbA4NebXSBDPmmbqjShixxV6hmn+x0pKmEcfsq/12Ddt
1qN02xE57vuzBP1MhSifgtKogYq43LUKabT6eEyWihVZBWcsxD6XwjgtvW/zAEr/
o4VPYZ9PZUKfCwo6h4lK0Gv0mW5bczAvJmt2c2ox56RAJaNY1fdYyL1n1tchKjYL
HXgssvx7MJuOz28gf7qunMR9F9F8OQqmHARHohX9ggNOOf308bySVAkXkmw4Ztez
nE7ymdZcNP9P6fYN6UXbcnCcpOhhmzj250wd0MP7DXhMw6rX4nR8Y++KcgN0H4Jx
MBIWAFjzXqmR42I5ZYt8ElHHmwT0lAN/U0p0RNQwuVQT9K3faUBOFKHlpZjw1/gB
YH/JWpOptgosAnJZsZBDuJf4Qx7M3PTkugObjkcsc9UnDKQZrSJXipH7ywgGqi+B
o72p8dT3sogK1tXZwSjqy/iYMYPvO2PxCLA2l0WvkltJuWrwBmAj/F2ER+9aEOsh
u4tQEb+xFrLCs+/KAvskYOYZrL3GjWKBGOYkgNkZYVno79FlTjS/PLjofGx/4K84
5vh7GXdOLiTRCz8XjNvpUNikdEUFenCpoy/yaXFIR8tozLRIxXw6kMFbpionoldt
zq62ODPLFvq9SQNViajW8HUKk9A2HnID0z194iEfyeoL98MPBZZwGd6vzi1heKIh
87sILgx7YIM0au+tHDD4ZJ03X4qLWr08sgxZSxmuam0NTyzwAnLr4xzQ6eG+qenF
Mgv4ItxHlrMC29GxB+lMVJhWbs4L+6sefyT8mnP1jiE6kbMgvmWUXfhDV4iIrkq6
KvOWrWgdU2/PZEyB6j9zx7LbnM+hO023Y+AUd9urvfRsUzxJ4grcgxZ3YYkP12f3
ADiL+UYLJK5qzX/LbsWFr3Lsx2BXOWTZKPVJdYrw/XdHil3A26Dr+Ht1oaBvcgwO
yJUawZU9nzQO91Vfsrf/clqlM1pcTqPd/IktgFnJ/9+vVqakOuFuUMkyUBw8/ZR2
u4mC9ZT9TPrijoVMBpBWVJa0gJ4yDc4Hqy2Bv1VWvjIDXA7D7j6cK1y8nuj4K0zM
Umyo5ujLcixTU3aCR6xHMEIq/8JLvGMUmj1IFrnTk4cNp7/qq8+F5vRNHHx8MSOG
KOpI9cy9Wo4lpgkcJT68pO/pN0G5pm8762S/ZkOUlnT8FcKqssa0Il6XPh8HcO9I
SiunjYlgYaFgwY/OoiIFE+K1YdiASfdZVpshHik0PB0XcHy5tWZB2D17cSfBnso8
Nn9CEYXiH4GyGWmHaxs7SJaaLoUXXiPTahRL6jW0zXLnHbs/qQO7erBSNoyjzdgH
V9wm1CUrEPMB7sylvUfrMomVt1bZrvwPojCY8bFFkthG/Mfm+tJEPUGjJWItdywh
Xn1tlcwZAzL4BI7EJYV8SRk7hJ/i9sChNGBF2pHgfG1y/woBlhplb1IEupi7eRhH
VA+7IVNIewLOcd08LGMGYCESIKHFWTt/X1Xmis83D3XiN0f8MEjc9Wxh8upK0Git
burzpUC165e4AFTwKTKPbH/WgZvUarwJnf+NvwiHK+SKKK6Zy62LcxyZI94Vg58i
5/Zc6bb+DkenE5DkdwUfiKJ5yeZ+Fo2hupYh2qzPfN4Br2b+aHCOoY1Bh1F7Kd0B
Sji0NzdHrbI02Bq2y8nJ9TIMhVxh9xvful3a9e3/P3hJPJ8SmDy86mY+B6i+V4eU
JTy5GbNEwkgrvOpPzCWOfLaAX6VFQ+KzCPjxSTZfi07LkZw9kOVO0w6zuehvMjVx
0F4PuXs9CFZLyXKjcbUZYW2Bm+lhmIZVjSnok5V/3Hda9QymNcAa6ysV1hcE8nEc
JnS68r7BLYrX1R4wiGhAQXeoxNVslgILGJsioVnT89M742Ky3BVkJiBW4OXG3P7I
kcYZB9UdnMHXy5+xA8nE+KcTSZT8LcRh/DBntrF0hrBEJPwqxbaOZLDVAsTwGSoL
VaPtV9fHf4O0/9VWGgiaDJu9BfDGIHq8A0fskaGFL1jyVKANjgJcloOzKMKW3KlO
ac9vkNTFDBT4RSdcF4Xc2Bc1q5SO03Et9sYHgvRkBFZ+iqEzeZzioVexSS8fu5Yq
5nw6f0Vu1svYBMTby7RWry4WkLbGTjCvuUZVz6+OyRRd0W43COty7DGbxnDIDOBW
j+KpzipGNl25Bs2acbbVjTES8MpKvKLFgTYnXLgLvMo2iCVylkIfZpMjqgPXGgkd
o/IoWcgtAUUT6YkDz3r2sOeGkuR2UEc/ftevKjyB2iQEPkbrafiLx9kOmbsAaLd0
mpV6yJMzrM00T3+arVRe2W9fvqitlkfKLrhHZz4Epv9OKTcaUqCDCohU2+bcIcxy
siPuEwJBc1PBRzUZsIbqdfry/YmdU4FklMshuYAkWMbiVGzy5MwjBDX9EWMKXtik
lIhz8jej2CV+H47M8piY9llyMkOSLk4F6dcBoiQ47oNASxYPCgVt1jLBmxesAJID
UeLLCw/Cv0t7zKmrKiNdO0q1NgjiIiXYAeqm6eHk3471quBl6WXnv9dZSt+2N+RI
V/g20WQxUDY4rUPjxafnjHSoHt0OP/t5WW1WKtwOMTUChH0hKumW8WTHpwotloCP
Q5Et7jBTEW3SUAEfeWACrC8UmXJpEfYV3uvtNmHexRtGU55bAFjioA0r5kq/WKYk
NlE+oODkNMGdJrgA+2GTLezTU2FowBVfLr51LQKDzihdZAiDWh0VVZSmSjkyQ9ni
UUYEkFtLUEihvZ9XFl4Be7YLwceLwX+ZIKomUGAaujcGFFjvYZjdtLuLVF91NarO
DDnc7zhPRuSYYJnqW6VUKvh+z04TC5ZKDyVzq0KDZo5rwGJZU9/qh7uNf7dN8fP2
cm42K91AwwUMaztp53uc+uZFOMFfuVelBeTaY40oxakYzmMAIkivuTr1Tj8VlDxe
P7qKdfarH6Nx9YAdybHik/QCUtt/5IfjHz7ulUL2d9ruwIHb5z34NWfZwHE44jZx
fT+ag0QBscFDO12JdG32TNh6aH5LXG36ssrWN9BBc9cr2RTfFhuDuNCLZrG+/7pe
l7/A2LTeli5NK1qYNe31x7Z87CzhKcZvmOq/xcRIXzOy75PHLdRDGGal9jqdN77G
ncwervPMGBUe71C6FjHChcLQ7AtbPVlinQOTXUsKP0JbBFe+OuW18VqZafoQ3x9k
+lFauxp2TplXlDbAG2xLgeZe0GJlrY3vfWXFMbJKyy6JzJjYa7+7wIMwyddlIEmV
+ZF5vgiz/7dOGrpdVcV5cWjBedLuf9rb4r8h/UX8sekgMQuon/Kr/nkbFFNwKKAu
q566iFZV0zvfmVdCALKZJ9R5uCMci2461I6nKnohWFo2mLeIP6DdrLyXc8/4OJ0D
HCsJNZjCFaaWxQYbEZD5xa+eX+sogqmg8fk+4Syjn9I20GfcENGr7NvVYalrcEdG
7Y2LWLtoqRrFra4/rSHBAz8lfPHQTQhNg/DgpqE76QB6zN+8NUURN26VTanCdSal
ttRT0OXGBOdkEOGyzXzA3k5VPoiq7negUce82DXmXXs5/uHvu7VZVFDlTPjBfnR8
g1pLlsnggCAJftj/tpTCuwlod9pf0NH0TR0Rrih4R+NPFyLxzvOyicXaQC6dKRln
p2h7755HR1RpgZu4l9CGDc9rSLt3qCKRD+m00m1mp7pGsDgv2c7R60Cijqse0B80
AS5LjQ4/Y+yNROlkzO5kNVayaujmpm0bk/N0i3S2qPIOMS8V2w1dontU0taqoKNX
5eAayUQ3eGm/uWUPtkF6bHBMSfmQ72zi4qRZ2fGtLlylZgJEo5xHjEtUlh8K/Xpj
PA6I1aTwDXvVoCA1wcHb7Arm3vvV+G0pOtpFKKuAxqgdZvCBR72ijfnmnqKgjG/J
a3y8AwZAVRg3wX+tpsfjT1aG6PogJhvgqy1sGeH0c1PsFY+xOG0ZGpA5G0FSVaER
2KDfVkLdNKQv/iOaRnyJxsofejHsHzDFv2auQKT/AjPzWX1kgn7NGbIZbcHasCPx
5P7ATPqSpOQyRsL45Aem5ingRI9+fwRuI1Lurb30jA/UryTsC0rzNlfM3CmfprwU
QleCguEFezfnWL8wFmm7Ygp04H8WM468rhL9HTVNA+Gz3UN2aZtxXBnkAknDy9mE
NVOpVJEdUo8vrMKGoqOtAUUUCiqEyAn6NTkq31nHsniWDt7VCDzwE9fFzrqcmLDm
mO4EgjY+AL6QChQfeLvxZ7Tyi2ptJVUMK8tRRKkcbCHIgYqooqYFCsnKkMQ2ae+4
z0Dwe5kN7cpR6YzPt76U1/UVAFm7qbnyOmrxBNaawsQKN6gPgbDUnzTTVdauLkIp
qXL2iJvePLFdJyJCyN8fNLxOYTsZUlGpiWLFWF9uK6aJ2Csy3b27l+Kx9o7BZlSY
gOElIaKd1UE5YoEV49vU4BTWwiz1QexMr4vRjIX11qoxJeA9QLxeWEdgsnLqI6fn
t26KQT2Nnb8geAsPWEJrEXjerhDv1AmdVcCURL37Dd/u7i7Xek2SifftxY2jAgQo
ZdcWFwmuLtsyHfKDdfCxabZ0zKrnI67148usKPjf3GeAxUzN48aI5q1pot4afBgA
4JbrcG4DW192caw/HEbQeuSeqGf3QGx2lpYkyAyshDOn8DL1w9go55Rwpdx0/hdQ
tTXJCqeHEzQajOSsI2d+ZP70j8sojReGJ7g2+ejk001rM/YdJ+pYV6XgCf4Tknpc
9MZZNGEBQ33XUPK61HZ5jUNlHIuNHe9nBgFkXqzGd0JZQpRiaVv/BN0IjuZBI+5R
szTxqzWh5gsDVXnmbV2fO5H56lRY8hZ8deksQCYLB+twYdlLHINEYPbgvkze98/v
Q65BJAI/GKxlTFiAgCcyQg==
`pragma protect end_protected
