// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
CEitw3Ny6weTJWiY+JqTvxkMMQsBZQvaTMyTx3nXSy6xyElHwsnB0RHfJv2xE1hB
x1f3nXUydhlCRnVh8+fc+H5brHNwRK0XYcWLh2ddSXZ9Cf5xB4d/+v/X6yjAssqm
4RAhkecmRQx1UJ4Ff5hQ5QrfYyxhA3Kphkt9HtPqrlow3OLzoJvlGA==
//pragma protect end_key_block
//pragma protect digest_block
JBVCkSCN8+jggOCbj8Wj0r5Lbu8=
//pragma protect end_digest_block
//pragma protect data_block
FEMQc4RKN7imMbAcMr/KXYf2Itn1CSbersPFRSnAHwKXdEHJLhxPbF+cMIJHTlsi
UfiTYnmqDChfFNKmuKELVUWYlZ8K49nSB5pAJDz2tEQXw9sf7qz3hvPstsVaMzLH
w1wz7VUFxEOaIXHwbxmG/OFjPp3XJvxpLYWWkLX9dE5yCssh4l+YJCCTmG75lgwe
W4dU0UvetV8bbzdWkBP6jQCTKV8UPRdRvxDPg03ZDUD8Tncf/qBG1Q4Zqg8ByYmX
oBTsY+m4iN5w8MuskXC/6mIb/K3PUPy39U6mPqnmTfPo8X3SrmAiTgP7ntWQ12Un
y70VXA9sHxy/ojQyw4CaSKG8+Se/WV/tRA/+ekOghfftEyadAeNPi+9cCrAasK2B
mSSjLC2L1Ezs9RHSMaLl4vvfmXtOO1pAT+UnpFdw0xP3Hb/nBS8Fm21OqSDDmBcU
i7xqjCBJdtkWdFC04TjcrP38Ag7ajfHGV3LTGhWiufsJB9/BbBaKfC6KIUg+rvDR
kabDqRDnjLAL4AQ9urbRopVheHEJBNnfuEuwGzzkpbxF8ilVc+9g8xm0HW8MI2/s
wcUFco5vp5UMyf5fwEr13enQ5hmeqmI+jGmHuXYoo05VHmbktmar9UrmbiTiP7dT
K9MFfrg6jSfbNsnG2H8OSN4fqiluhfjOrgJIxb9wfIjn3O9meUNlh39S7TOduCJA
qw05K6d8h99zbh3Z00EPFMJ/MqDIJWSjWFWtS8wCjVXG7H8uO2qHPs3NM9tDCeiU
7+Q8OKKw8R+FydnDgKgphluma8uM1TVUGMyhNXrBNz0RsCTGm2U/666Q9RQz9BAH
Gla97BriaC3jBzZvk2FnZuX7qhGkgk7kcRdjitB+6t8psLdoAaGN9jtG/5bKzlD4
e41wfw4O6bdmHGFgBKP0g9NL9q1srYBr3uFZHt/wZ5n5G0hPioOZQS1gD1lVVWky
f11Jgujany3FuKkUtf10uS/fh4huVQY8oJVM0n983mDEnL/xBCYcjKnqqqRsUsQS
z8hV/6VwSar0LcI9fC8cxuVDr/CAs1qQtzQTI2Ww6/c6qfAYZPmHlGCZ61RmdSEE
WKC65s1Qi3/l5zsc6dXyqlOW0/Si7V9loMBymk5PcBIT8qjprz1nnZpA7To052ra
uTSPsTontf5NqF6V9oRO7MEZ7lQc7jabnuknyzyx3gLSQmDaXbbFQAb/M7o6THA+
zBk5mjcCYUXrdXmFnJ9hWgnqVCp6z9YZ4DdEQPml3rlX9D5h3Vd5FBWC6nIc359n
XxVLuYufikaNdzhjAMGfifBPqnx7PM0KOAYWCDOd91iPQjtqB9OgH0/7I2VBRjc9
MycDKzA99UDRicyUh7/M4P+o6JwqkbMRJ0bmj/fQU3lvCLUFcxwhDcn8MuL/Nnjs
O1xDmOL+MFQa+RTtPGMsvuvxsZmFcHtaKFfZJHqvoeOEgpV1ozQ9GnFJQybfjIoQ
JSaRs5FvnpKJaFcsRWS9Z+j+ZvplthDTaURGQhVoF/5pB2FMTFCFWJndFkrg6yyI
2YOZRckHqMbJlAoN77lNFGkEu7IjYuPp1hkWE2j8cYkUwQtRJ3MichtFoSQt8q9v
LiQGP5EAYaDyiri9NqsDfjZqkWJFl1YRLmlTLO+58GwGZrGhSnknWSM6eZc/awV2
i7wOGgWni/en+Sx2l8kkRz4XFBJncgDoWVI+YMTXlRXewobGC1SbxvtjCvFVu0Sv
vS5KzOviZU99onDdEYG5qUdN3DbFmngc6Lf5OuBZSZ/O7A3/wqjMnqjNdUex+J7F
ldSws04+e/eucvOj+BV1ifCjEhjtLYpX3e+WNK7jDv90QNJV7LKKU/NUqc84doLA
f4n4BVoyqA+jg3lTC61/qfAmz3zO3yyavDZfwVnExu/mo7dbch7HFAY68hm8V6sh
kjvbh6aKafzc3IsQI4T6MfYap+paWDJoKw6gIp3SFCu5DVC682CYhWg7qx0WB5d3
TN6jPjff9artRsUt5KQ18+I5sOSlAmqJo+zud+qXcynbfSFZ5t0+4DnJXhnll2xG
F8aTC5iWKZZvS4KhVASapHyu5Td7oh5DEYPVHLsqUm9vF4+ycOb0RfIc9u6nlsMw
cAsUMle3VpjfnFYn/iREGC+Mc0iultkHhpPNpPUU6jNmP3o9XzbXM5OB6w7dn1kc
83RNkU8Pc2Dwn6mDXGEfLyqhGigKFFBqz7aNT6CNhWlH/XHucA8tIzJxK+aQNuAY
17zzzttv8HUnUpT/sLearKcVI3JluBjotkYx/UWolkP+7yc7l7YNn8XBTghZ9FYl
B4W73E9mQ79GSvOrkKsd4nJeZItmYS3wuK3WwXRFupdFA9bBC6LKsLNaYoRvYNn9
bdcwYN4rqKCqEWp7IojmC77RM8Kou1+ZjZ+RHajfpKMNkvZixy5KqmqVcsas1vsZ
ByoHCHxUTPi2x5m3OIW0kMGKvMVBxQO7yJGWfI1V+SxwZEb56XWqBEcx43Fa1Lsj
8FZopCqADR90eGOJ4/zrwr1/tBCh8WAGhoT3FlnWuNJHx88Yn5E+B4kYUqIEoiYy
hOxl5gp++0g4Jn2o7ObiiYtNzIvfg6x1xyb7dQekgW/CzukKXNTlacZosECbf+lu
Tnf8ljZup0/yxf1SvTlXSY2rAgDggo0SEbUk15xgtOaFVftVJDD6jnD7T+F1ML9Y
tE6jv8ApOFI6rYIaWL4ZySOQW2jKXIb6E3YTBRl/dJlAvYEXzo1EKw4dLH0nHbf7
P9ZIaM72v468lkmGpM5DGf7R5oIrWhqfo7rz9xek3IXr7qESvA2tO5s6YSj4b+UE
6cCc8jGoZlshhJVQ0iRqGMb38dFmcVJKyfCHQsxiiWih4dIEMk1NScS9CxBvfd+1
u05aCU63UsJZhVxYENO6/5nqf9oz7OlEEVQKJi7h5WPLzLYrV7fKbo8UTgeQl0qa
qvHhMq8xiUCS7IszQwsIigy682tJScSgHzkvZcNxPwkCkVXBj2Jrx1PhONAEqByJ
l1wfoA3KJFwuJEYCEVcQazS5DF2PYgG+Z6jUatIOMTvoCY++yD2XjQxG2Orty+rM
PWpAW03sgWT/USxWgcGtqSeViNNHpMjst1FzbAUrevqaQDLgS4NM5cReiWsAv3dC
VcRCVCjRfs1itNJuNbkDW8jWvWgQMX4jx79k9un1Unq+DKNdljuTbvFSnhivvLId
3RE782r3OfgwYurjJiWu+0d6qnP6SKP1K+sVICEwoOLyQntm5IQreSdp63Kv4rot
R+w+oRdqiBaLI4E6aqhc0VBcyUD090ZmWkQAeEqTxkV+3UotVzn8ybrQW6sXP7aH
BY9mBvBAYf0zVOixrw7lVtwaRY9c087YeS+I0B4O3PGEAZB8LV9GrJycqyievGsE
Bs7VORcKrLTclPPiwLGuAkBzGgtKOiKUEaQ2N+Sr/jmTXcVnkUHioeQC6MsTiAfl
AFUtSFKb9dQOEjLDOpHe2jKL51vIv4phSsWY3M5Qg4pF2cl5NqR/BbY1v4JFVsd+
z125bVYirWRJvA81FtGQVJZtg+WwuxIVrcjo1QTM/+ug3ErqeORD5hJxJh8cvHmP
d5/oQjsLDvYzzxMxD3G4FDgvuUdW6ebrJqiQVr+ulbQLdaqtmRfCOpX3/GLEJS75
0Y0xOccFQPpjQv02DYHhgENVfVdAu5auf4y6wcCm4KqJyNFm5Qq1wMkN2vnIdt1B
P/qsexxApkbswwAymKWRsjdA4b9o+Db116+QSRKIB06nzYWDGHRF/oTwEX66upUX
f2pS8hExB3nuVl7ilzNM+AWFzBTxq26sRsoNPUVZJPb7Jz9GQRV0nCj8gnhsF7iU
RT6LVDfabDTWlWIK6Gi+HvyrZ3apSLC6PhBTw16STmV3L9iOhOd1Wb9A/HwDwZlo
KL+jxNi4++V9biTkYretrScgx9AMWAbCqJlbZ8aqHAGECApdTb5V/6cd7fzCTeMi
HjtPqGcTQsmHpX15ZsBAkuFe7v7QBqvC2MYwitjVe8a8pOVB3Afm8lJz9FXCt/xi
bI6hBQUqrjbzSJ1/qfxYiFvDc01Kkhslb81UxuTaW/zxmZ7HyueoK082GcmNY0J5
mCRr5g+MXti8ZZ5yd1U6xBo7+OfpamyUW7pHew2bJnznPKnPswDW7xyn4wetdrM3
y5sWoMWmeYs47nhm40N9vN3BvDCEYu6H3LUQ8WaMWBNtnNKGnaLa05nWqg3fJH7q
if0WK3gKS0HuT8eW3vKBmjzcdB+vdAhCkHKFaVd/uJsLqMUcFFKzBxTDFDg5yOYJ
H/YCjYDs694Xd+Zu8/XQKZcjCErar5HjNdyVtSOwY3PVZ/ORixIIcwjaipfd9HdV
UXQS1inJDJ2HNp/GN9QqTpGFEa7wFlw4Z6bYggVNnqsfW7uiXKW/rlnaEeyn7jdF
BDqAgR/TyEl6Vlk/j0Nu0haMH+1fkZZx+vyWpx7xstWlbUgUqVJ1gzyr/GpiFsr7
BOlxYEgTfiWPqR7P5ifFG3tnPpRgVSain79S38gS4j+Z/4wJyQEeXAV7WIL7B/SH
fxQaY3G39eIj4wqcq5IoqdfDZwvqVq5PCEuyNuLVml6EVdPEaa/XnBk8v33HF8yQ
KqvQL/LHuR4t81DRASnNXX0ri7JTs6gWSRUzHSRcDs0xTuYbODbL0ssCFMVSEsY5
XloIaHDfYk4O8z/nqLVD4ebOjzvky3C64kfMLmMdfBpxJKlGmAid85r9lsyZk5r+
9CsglmyhDlGN99mwQaurhIGw7JY8y2rqekZksqsXvZ4K0OZbiG5OQZFq6KtdPvCs
cCyMLiXcco3AyP+kNwTs5F9aaSTCr8sQP/meBarHvI3mvRHWs0Bx9y+BBwdljENY
bizkMo1DCWYRFb3AHDDmBHYw/J6tmM4wVHzx2S/mK5utaVyn22elMV8sz9FAuPGp
LZpOO6+3tM2eFqLE1Xv4ZiBj8Z/lc1XsWcCcCQn0MrkEm/5ixjvn7XUGNc1BnJDy
fiAO55piwh5qz2QxaidIWmaSSi3gOmNQXdL3nSTu9/nDWVzNUhVu0Qb3XifY3HET
0r/R7R54fLb1O/Bx8MKNBJg8UVsKFIYcodP+WO9P7Ed/YqWUtfAyxV6n1NcAFq6c
sMD+RVY1kymCAH92j3ZT9bHHk3mn0ieSY6UdRQtJ9HFJ1SEeJcYlkgWE6IHYBO57
wXUtBp6tz4eElK40tP9GnN+3C84WRlH4omrm7yhbXQniCm+P64OJvskvNyVkxXeH
fB+KZTaFRgWcHueBAPGa53dUWoS+fUHWlvPcHlE+ox8N3fP7mzILWQ/cOUvSf6Ab
OcQMkPWuBz+VxNdfmHyfj5qPpR9XuyAy7t1+7yjV1jbwV63gNVHxWO2Rwam70svQ
eGRlztvsJnSJHp3uTPha2osYTBfExPCK1rTCk2B175blpF3uEKtzM5ojU2mH6dzm
GR9X/K0EcO+5do7CyVFA976Szcr5dDqs/HF2AYRfBB3CIG7ftIvNQG6C65Yy5khR
E2K+cOyWig+JZwkIUgfwbtTiIZJVWcw6N6R35WYSxplkpYL/lbnRuQWTx7TMfsw4
Li+iqrsG1opOViFVmFzmlvQuJx0ls0V3L6W/iulSzZjEUDWbVU1s6D8zq68vXyn0
DdMvgJzjLBNmpso++FQFKpA5atYU/plISQp9c/w4r/d11YBVH7Q1YwO3ZeTuFr88
CK74GYK3T0bJGWlgwBKfHEH8/Iy6SrrkufF9i8O/jZosxhoRZ4T7uUm5A/wpKNFC
h6fEouP6yBsi8nayFRahpD6hYjqj4zdHkbN0AQAOeSCmT5/YMd2TH+cVR/RB1w9T
erVBmLMv6aSTwDCaOfZWmg9ALYKQY5/5bYGnebQWqQkUpcBB7etE/NTUyhJvx0Yr
rtDM57wDY86r1599wNYtYGYOtYxzMsiPWYxYayHu9jc+bVqJs50iThkHCUIRdnYN
MCvzSUb/Jaj9R/fdNO0yC0LqlsCW1H81SZPuYYNOwc7mJ8JxPHwNuA4VfEjTgDtg
LDFfrAySAXWjtMfhrEa5pDDDHjhhD+N/phEAhcbHWyssnMyTxbJJgx68jdwjobWz
yEcLcjMwBX3qLZfCM0KlBCbURlBPu8CEgbwMR7UOzqbLS0WaM0R1csY1EwUJ3L+p
94lSDqYyNRyjw/gyEdEEE6qzzkz8CaULXs6dpXhNVPODuBj1YcCf514f8V0XlfOQ
aIgLwVtQkIpegj42hHMxACZ5hDvrhFme87wUkbeTbvRbxLVxlWZgHad6Jup487kX
XKzvtdKSUU9KIZ+M/4gfcGodVHSO+JVCmo9oPKPrMDrhUY/2avboYzjPYibaFYdQ
LmryN8KTTQ3DBGJ8jZYHZ53MzrbHH5lkXbOzgjg2ierVzWdz7vn6GmcxHKJrqCKY
al8ibYgl0lH3UiOgcWngBejtZrrKr+eOJamYPK+QXJp5gEjeY5jZ/zXqY318PYkJ
nvM9kL7nNktuc1RjhRUY/DVBFjyRQGPR8IHT+vjAruCt1XOiA/SHA94AC9nbj4Kp
NW4qc2xuwNO/kpwcPHcPXR9NlYT9vlliOrpa8HY1aJVC2xA1QNVM8vxRIphuaLob
bw2mS3I5zeSggrUOwDwc/Oxuh9FyAvd0PkWEvYLDqOfbqNwh/hzXSLmbZzdcUaZs
KQNU7TC3ouXkGZxKpxTjQUphx77fWvNiDvIBudkOCoMzpki2cdWuSK9uuZAiCaJv
OQMy2lCpooj2SMlVOfzVWF1qL5U+0zrUPThhVVdoUltagKQJRMd3EZyLzTZuPI++
xLcbu5VsGtR01iQTZ/6LvSqLNRzmW6azsiq2DYbmIJoSeJDzWTgsykLbEcVX0ZcW
pxGs7cxJk9bWRpXfAkm5xumeLFvDPfyxIUYYsbFJR4KYWHTdkgDdQYchx37WdRaS
CKe7Y+LbVNXHPxS3e8irjMwP1NAT1ywC0VVpWTMcaKFb/VRLmwBJmww9zcsn5zS3
Q74MrqQ5+dxpvTXgOHGklqt9qp5fGjRuD4ttbB4hUC9wVZJg2oZgS7N1Ue1ADTcZ
rbioxDAEyQHVhIGrUqvS8I4mogkajG2SyMQsJPKE12D2zt7sllz9K/gV1XvC/Ik6
+alM/E9KSkWl7+m/3snrKMD/gkLRkM8ja8nHtMkNynuvNbFecF8JDIZ5SUlgbwLz
BNwpyvvSH4uA4aDOKufkPx2xBh7wvszjHDqltmO5Bu2gz464kZ/i7c1TGFpOdMZL
0OMv5318XngbSSUl1aO9jMg8YNn4lPjyXD5ynoIk2MHmRtMQeHFo0CJuVqHXscAP
Il+4T576ZDy2VXT7jUyWiZMR9i6+hXduzYy6JO5DMfawiO8oUL5zD3Un37T8K6gu
N1QBL5nJ788ZI36tUQiOHSeayGrSOq5dwrTT+z5CEW0EvqTYQmcPQ4Ek5dSJJDNm
yEPoRbMFcZgN2WppzPFdgrOP4COvijqC95mxUHVEoFSNIVE8L4BVigLtyQUcfgvP
4JfvC7FrgPuawDiidwtoI0FfTtf42itDIsLr5NE9e2y2HJUvfIehK8De/l8f6h5D
Ey/FvoxY9tsPM/Efzdf6a9XCOYhjkzffusV/liHKfaJuLT8VOIc1/jw+H4DBp9dz
7q5bQsbypWQ0a4foxaeVnrdyfDJN+h5JgYjJfzgu0oZU7Trz/cvTnIJDkAfdSZuN
CoeInEV5mAWMHBrxl+aN1I+6grzW4MahL2n8st5MiDHlwW7ex4t8+peUO59bjCy7
9gV+KoW1sQ9DIUE8RYnYIRssfQ25ldOPGD/L0k4iMkW1bGeJFwXzN4lqMu4bCeUj
/x1c3TPwrvE57fodWCSFD4KuZipF1MIniG5suqnC+gfvPAZDQy4ZIAfZ1Qe8qPsW
40O1i927PIqtNM0ux7v0xy8SGxi221262yrTfoiSHIg2w8asnwLQzjgtLKajtAl/
JF3nR1ZDyc0R8ffthaWpMiZsKZHyE2QVmcncXsOw2T1OHew9ipQ06oDhIq9JO4Pz
1nNPncjFVbRZ0zxYvF+rH5tNfQ7OFgupcKSvzXm7SYXyTLKboCdaBBmRV0NtRPp5
wMCpcHXyDnn4X5ZRGYBjQYgCqxEV72maK64XAWFCUTjgcFWYytsXAM+I5HftOqCu
jz0zoclOSEP8M3mfL8AVaGegny55E3aD3+uHiOp5PpomW6oH3AOayA1LCDgLnpcA
F26DGstkEQ/rwv41RG5O8RjBKWBoi2hx6XQp6/3ehtysleKf/9exKR4lllAc9vgI
fA7U9y/Cbmw3558Kl2A7e5ofTthW5RcqXAZ6kRI1qqZc+fnAAf8CnvaIPbWd36mb
Iv8egDEtLoCuYjxBUyX1da8AXz1/S129VEDvQI/7SaOZOzI8E+G5Ak2f4RX/gbLU
rFTbrlQTkycK7Ualf9zERhogCJRY9WaZHCSc/sa8uNuSRlwFsaPnh1i8/eAXMd+e
Cpw4lwzzla07E1QyPC8WWxj8jiqiLosQPQW5H3ofIrPBK+2C5QdMItq63PtOUoWO
p/JkSAJtXkH4lwNIP1AHOy1BIPa0CeFpmlVhzFdKurDmbDN3HVFQqGxz6AWH7D9a
9uhimXC9QGJk+92ic17oXmRZV9HbpUz8gdlKRQ3iOMk6bYFOwdEQK2Fh7fxVdGB9
+OI3Ojgpuj08+Eg+cyJKdYYVCWN73bnzATsEsSq03UhwOdGdhtT62YVULDJfNnzI
MMdMIHeJgYTziT+1l2OE43uvhxTnn+HmFPtrUxsR0vhmI94tN1h7/xmQLmMolMLc
Q5n0S0VdyoIAX6n91pjawXl2IwpERLYH+6OYNtASEIvjFQm0EKoeNy37Uuzlewwp
IPEBRnlHc0CBFT/p/RgMuearssFwYhkHpFB4GQYA02WkDF3PZ8wrpySZnSFucZM1
OT7TmxKnUX5h6G8CsnEahIpJ9u6qZQWVYmVhShLU6GkHMFUJYslxCCihWcUM6DR4
a6lZFtOg3Sytc1BygDokDbeSiGWDxbuK9x95nmTnzdzIhAQTO0LN6aOpRnzw2Vwg
jRBP5spaXk9Ohu3Hu7FTej8rUcEJ/x1ZZvdnK2ve7QOTgGjT1fSaDGYxVKQkfz9w
bPZ3hQmKqwJb/Mu8ItdXA6uOp7dl4Q+43Z5LQKfy3HUNj4aDlOLndfCNXPjvRVDT
iW0bqasj3gzya4yWaTTAm2GCc/n5Av23CrfEnwRembSlD2T5336/nzdnvrhmtyKl
YGcrc+HlgLh7s7a5npJXM8vRLueISDkG+fM4dfXmeTaz0ahA2OeuOs7/Vu2LLLYj
Q7AqXDJFFM9+bRuK6ihiimXiMZ4eEBO4mokyF3+fRmjaUF48QqcKiD1P5WFp7Yp3
xOh9teF0v2ANNu+Htgf7E1CFuDSiAQLVkQ+PqBLGTqPz72BAW3GY1ECLb96f9ttu
/I0mgrxz8H/RucRov1rAOIvT2fjc+Q2WQAHTSJjqpO8PhhmZWW+uTsLyhtV7ngb4
oO83rScb3PME4TirrbgzFrs1jlVHCUJJZX5z/hJWchnIuunM95NB+E3C8PwnHAzK
vLK3F2+WnDhMuBBev/YPiT8jOie7P4y19joV/9G+GlnUONcT+3nGbP2nXNpQb1FM
S1/SuL81iEgdItTp4obWpvm4kj1TpL3OItTvqkEHd0y83CtbMVbDbwIT0tyGMimK
P5O7K7JmhlN+W1daP5chax0Yq7FAJEnpSInDywKgQlccoXedBG61YdrGThSh1UOM
NthSf5vDTb/ydXt/7QsuOFQ4MkiYIHQdkuUHkzTVmEahXXF/PzRVk0uqmezDWZjK
V3V4uXTZ8DESqN6Zv51aTnYKL3VYa9kUkjzSDZvD1QaorWWqutzxwqYwp44q0gSu
I4y1MDWJvkF6WF++D0jIc5XKlA3xlZ0LqIgPWsNz8VhCUSkUk9o4X4mcWJ7Pkisw
CAqYTr7l1sGWnu9d0+RcPNsitHV5DuFe9ExkCgjeReknBi7F0Xv3YkPnAnGR41Tn
yJy0fH/CgbWqM+/PsfCcrJCNXY7cfeFtUEcOUHkJMudeoLnh6VdYgKsC7MeOdQBA
RwncbCAyi/10wpjh+C/MA3i9iP2ZxNGrMgL5OCZks5nspQQ+4EVUma+Lw+6fxidk
72iCI5RO72uD7TPB5TGyy96SdkDozuVAvaLH37HkOHU4Li46qqDryhMEISV1JcbG
HGpLuf/glDt/Anl5zimziQ==
//pragma protect end_data_block
//pragma protect digest_block
lfbTVYKMl1AAWlLNmuFtKBN09qw=
//pragma protect end_digest_block
//pragma protect end_protected
