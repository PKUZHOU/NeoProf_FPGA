`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
kg4r5v3XLwVGm3XsVse3bziVnDCY9o7kny2sKRK1l/9FDaZZxAJvMJidG1mk4iQE
aVT1T3XWc/eRFPCHpJrA/V7CErQQC25TOt7yyrm2B1dGj3NNx1FGL5K0W+2h1v3D
Fkem53QXNR7LNFVrWzN4jcjs5NExztJXYoLgupYqf2A=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4144), data_block
e6qi9zdvlRjJ/IyHtO2ltt+dr9zbm/bL50VJ+Gd4Yn6UCCBtaV0c4Pu8QF23NgiV
qxLTVb8NgibJ/bylDLUpThSKKw9evG27+rQDpNDPiWfqtYecfGr+mAUTGpTsgUN4
kf6M596w0hlU+Od5yUiY2DqpXDdi0tq/nZ8R/9rIOyah6dWsiavf/Bb/o+dvMNyo
bH04U85sYy3UdHceXeqs2Hm+6q3cfqQquBGvRdxRXmFaXevIdw31xSxAKp5HyifW
hw72Ahb33qDrNVXWrhkYoXojDeJT2NmzszOEXw/3ENAZIUXdxFIf2pBDmfOQiTN6
FxDP5xrMhbHEGrfIXdKD0t5fm+4nfnbY2b7lzgS9zEXzv+eXjzQ7ioaw9/DRPiTF
WWuzKUm9rvwdPTwLFdGo0Axt1YjCEmsUnoMQWlyUQcPY63xqFUd4zBuoo9P3Fp6a
/3A4LeXT/00W/BV63TsSrKp71FeUMLwvcVTsCQQpJvalcM1PkrwxhAF9SAa8T1jY
3gmepi2M/nwUyVT/1Y83nE/TiZwAzzewKJ2A1ybuHsFy/OcN+dmTC2Fspq+tRjIc
ZDlxNNDjLKA+2byeESD+0sZfi/HfgTzO9LNLyfq4XneLeBzD3FYBFnujoiS0JDW5
z3kmCBIX9R3f7XRdxI2SBvY8MnPRA1NyQmNdv51MOFFw4haKpCV35Q50lhRVUBkH
9uW0u0dNoz/PZWfKiD10Pbo2Nfa/1PZOvIhpbnGiJfXItPb1YRhu8j44cUN0cMZ9
4KyFiArRx+E0iGew6BLwqo2kSRgsQu93HFLLf5QKFGZagx5ksx4IEp4JCL8Vm/Hw
o3RU1TEfzml40KE+eooMWC3CtdhUOGQK3f3lrOrAo6OIICMwQCLh4eHOP4rmed20
maLgiVgdvpqTktHNsNpLku1OfpY2h3yborC19AW8pCdXpvHTn0gUWH/uh0Omj17x
x5vSNpm6iKqwO+71xKvy5W0PeH9P1ErUMpPKu4tegkfW2Q5SyJazLlgZLdOjGmuu
fZKmKNy7jPdRWYNPPnjgo2MGldyGzN6Km+ZICt95II9NK9DhUudM5AQKlRrZ8fH0
lAYuAaNLsZpNxgKo6LVSrNPEoubM3/9LkxVg3uLZ/6zGqppEGrWMvSjwTIaF6c2r
tMx4IKh4DSZ6zklVW2atl3knILakoPn26P0VRECoyASWzTl7lJCNemxYY1dH64bA
5VF43KScTW3KieWUeThPr6tAzFUe6CvXXstCtUixqVs1QVDGcMj8GdSnzMMvthoF
tSiSocLlDViUNJqagSXlvY4QxPtX996uXKxilB+L2nz/+s2LD2MvOXAjIGwHI4ZR
XXDheCeiOinflsisGPYkUKJH4oaFPSaOB0w0WwVrsgs7ajuUVvBGR+5lGZaMdbj2
4lvisIlGcQSugOeBe17OWLSu1gjygF/z3/Hs1K8WckNRTGRPdvFSjaBC6gSQswOr
IoLv7pYR8Ag1F9u/VsNMB1k1jH7d+ZC11CTKssM8r3Lk4ss6lqJ1Ew3H6Xm76IZD
Limzx7K3J5PTpoMGOiv6zx7gmyfDgSOd9t67Xrtoh0qq1BbSU/pLgV82r2hz16fq
T+ov3hNO53YjhDkQhPjgsGPQ/aesZCZWPzax69Co6zKajDaWxkrF/OcAqogK9w1R
XToOc4OtZOHSkQYQ4VBHWUZ+81nYxkhFW0OjJl7EMMi0PUoPDERFTsoF7NPLv40F
QIvrR0dMVj76mNhXVKOOf4tEv0Q8MkUbpMc1blnHdReWDBFHc51AsMXC+SCbxlE4
auN7DtAVeCyDC5YPo+vPhGdQ3pnPpSFw6SmdziNWdaDtJiKCm9p8rKYTlc0s914P
fOshVTsGh4gPElgLnuc0IcWd83ZSp+oPq9FuNegfnsX3heloQNXWmP8ohzVOD9R2
hi9xbe1Q+Kks3NLTDQh02uyT0A4qxvTBGwCwSRDJUBmvL7PItxuS/7znhd2+wP0f
JZJNVCjd0vFTKOmh9k8UBockYsAgWSVqcx5xq5+O/wUfd8xk5GeRdBV0DZOusOgM
8dM6PGeZ3BqlMIN6xqWuIs97EllNH/F6h5+CSM9QR05hygKbn9FtaYHRMzORo2E4
kGQ7zIJNto4/9aZKJ/e/VVCCW+0trFLcDs/I0+WQL/p7kWhYz2yo3XAbsPPGBLpL
+b6huGWTjw/PsFjkI45CbMpFJR6PZ82N1YLoKcpPQ1SUVAFWRA3DS71SBLASrE3V
eP7ocw12aJB5OsfUqb4TH3OcYpuP85h7pUOFLbzNmdNdbUMk+1PqG1D/F7pQNjln
9llkgQgB/8S6mR18R+fHqd0Xfiu9FB51EXL8hGMK8/ZDgR4dOiSU5cI3VnX1afmx
ClhPgoaz43DWBI8Uhs8vN0ZKLo8N4V9KWhjq3F9NaVayLYRRWl9df5E8AAvUFG1f
PzVazseHncJF85/yNSRUbKLT5sPptKTnv8O2pIkrD9fY5b3MOYBlRHPnpxDXWtnp
LZD/Zsd9tQuCoNxUc2o/FqLMYld/gDNnbGg+RTWAYM7UkqRXCXMi2STMzWroA9rX
Lmi4ZZ5MN5AFfV9DBRqb/zWDngjKExetgYK7a5XVvK+tLuI4cX/nSpReh74D7RUM
QDOmuzG3brO8Znks1V338+UmzxkJ/dF1JoQoniXTV3MgxeQKDrRdm2HfCzfvpB4p
pZ9UJR58c/4Pcfiq8NDI6c1MEIAOItcC+anzkAk5Fkvsnn94FgF3OeoAF/1hcbZq
NCz9aETqEj0UYq/PDbugCMD+/aXCO3xTcflCTGE8NfBJRA8ZVL50gbSkcnfUZ/Xd
s/K6fxbW3z4NU/Pf4sBcgvNfxZT8DL/dtWib4oU/SM6Sc/PsnUz6BR/ZGcQWMtDF
g+uGkVN9/sgLnco0X6g5yH2lV/AmouwJUylzV+R+VfiRKKK//u3/9VCxXFqV5VuR
sIqkFs1C1af0V5p4GMbXsiDtbFjvGAkkx67OF42WIJT3gP0qsgClvVd6Wmw/mJ1a
/k0Pj4DeKfymkIGAGb/f6n5nOewGOLhgjX+A/IzODDFBnhWDv9m9aYqd1JOikCqp
q8tOoYbiwuX9MuCFc7BA/8paS473WdlAI+pPCkpfntxvo2NvPuvWiivsdwdLFWmJ
1smilVDsh/ooJr9AhIfITLahNGFN+BegIF0vpHFfQiC8ag4frLAkD8bxSZhfeB7L
f8hJRQ3JqGAwxoL+0mY7WFRRsZ8Lhw2+1Sko7GP5QImVEx4Uk1cO5kIQC7Ao8qVn
vLC7PHwBGIQ4SZ2MtLV+zducGETWsJqUwn+96e8eKUdCUI8bb6YL/YZvsgPOnlh2
+GlP5ayRX4z76TjNWadYsbf5OmggtCyX/S6zIDv5pZRyfbUFTDDA+118UuOrjGTq
E/2z70rnOvtCShrqD4xDhWAi66/nZ8m+HpIJMFX6iQ36sNM6TGINWFEn4TDeClAg
34wYwe+MbgtdIDZnr9G1SNBCqsyY0DsWgGTqMtTkS3Y1axZgzmrxZqMrBZPWnGBY
/C6wDseid5r8YLgWr+ixxYpXYj6FhFzTBktKYAfdbIIjzYVyVJD7NhZONdqaO+dO
8kMxIbXYEXChQ9X4V7z7ixQBAo+UIuT5aHz8jloSkkxn9B62Knx/MyOr/tYXusSH
1reYDqIbv62loKsv4GMy8QDR6gGuRh0v58rRBnlz1529+iTEPH59N38lVO13pMtV
YVY7h/qcESHDBdIfNCbXASDpg87bY5N3/JNW3P15uKU6VJLHAJuFZlxyHa+jHmWG
kiERGWoHb4b+RDg9VpwgDiEbLLIbvQWP8llJeyNWAW5Z1fv31tq5NqFyOA9hR7Cd
eJSPMD5jHtyTrDYPvxsvYyU1d9mQ4oHL4EqoSvpIJ5/5znKVPRBldFMw2FkpakHE
dDgS9Zi8ZIHqLejbNGqhPpQfFutCNLxTWRbLGS+ytFHHG2ElqNSM12B/VR9uDL21
Inb5w/opsTvoRBRQJR/0z1fCeGQwJSad3PywWjelBj69eLjBX/41qaqqJ/WrCoh2
clG+qgr9j9nN+qQ207nA96UKnVoPXkSguiRHa9AaTkWFW2/BNVcMvoCJ9dXuH612
KkSAO1ylOMWN3YTvnkacr1TsF8rm+qQaITMi18cHJ/Ur8gU/eNeOSYgGt2aVgc9X
izdzDQ/Jv2CVwfDvd1+dakG5m7n8PQfIvyR89wlhPThfFFS0jP10mM/2HMOSryW7
7OyKZ6VED6OplYjnK82TWD2poWsnYpQuLOMO42jtjiEHXrgWX3tGER3KfUKeE4+R
z/CgavgVmuit62JCh9XHo8DJrCgT/zcuVyNHZNfU/hZF8Q5ilOnRX2MfjxrHu0V5
Ey5+PFWWyRKFH2aRrxUnvVpxl5REsB6Nl6W2jPh7WAbLE4plSANSEH0LyReEEs4G
bIBsLJdoJc1lWvIBsG+Yw35i9ZN/kBi0hO4KRYM0PEUJMfH4OSEqVj54+zsTeSD3
vL8RJYsiTnc1YlVy02TEs6McTnd5U1PbwxkC4OqL6FrSP8YhdVVvKUpRdufkf7sf
A0F6y0mulWx9bElK0yAm9dpsUCyUN/EOV2SaDnDFgiqZNmbFJhLNVMDLWFPdK567
7ptJm4OjskBEm+RHB8nDCMxErmSCvfOY3S0nFO7+Kft3kilrH0mFBnQeteeMF6cl
9W+10CD2ZSWNkNwG90KouKReROiyk0FZs9D0450YVLuEsmMZG7qzBpEWSEOE9T5P
wBWOvhoUVude4/s4QA0N6et1bOuoePnMmuXT8D+0gf41mlFQF/4fWL4JG29dxqNp
2uj4hqT/4D7Fqlwq9IKffqgA6+5Tu87wshIg4R78zujKyX0WM/QH0xNSFSihfdnR
RzrJm6s5WFUreME0+lhZXjCtqhD4DGpU4wQTeKu3RbZf58/gKpDZCdX0I/RKC+th
O7NvttzvhhmteR4V1L8N9C4KTh/Bvd+9Yjrmd82v5V2PpNKlvzHkW/P1bsOavIT8
y+2WOA9mYxNBqg20G5f7S4xhZck4O9WWQsLzVjJw52Coin1FiRpqubvT3LDfB1gN
2SweLTfY7RoHhtij8XLTCzlkJ7fo/xPNhi1Tm9a4nTvgiMgUCMCViDU/fMKxknT2
/YEqfSsYAbywSdia07GFwr0A5avoQzESn/r95w0ScA0T06YsjozwU8NXaAx7aJ7V
2yrDnN6XMbrMLvOJrM+cmlY//gMt1E35wnT9rqQ/bAmHgKqAgwctATKIU6Iw+SsV
7tas7tgy/kJlXLxg7R2zOZLn+JyOWJrvJwabJclh/C+2JL1pvoeQ6BwzYd6hYj58
EomXQ4GPwUG+25dxDSVNhoxZ486ajAc9JWhmQSRbL8lyw3kjwu/hx1+WoNR+6dg6
S7VqhElnXJx1Sr7E+gK6b5kFkpceJsZ+8dcqjeuJxqzIC43ZJ8tdvgor0Cl3vayY
8bRXW/+aQBHVzGy6q6XFjdET7OgCspxpODs0Zvx2hjzoHe7yHTurb2WRznnamHLQ
+uWT6N/zP4E3BWaGigRHzg==
`pragma protect end_protected
