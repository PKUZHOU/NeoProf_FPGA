// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Dcte9ot3JrkunWqYxtwaAH+T2GJCpejsAGrFSlWbgoutgY1aLakRsVrwZaxlPd4n
GRzMaVjTJQfUvV+BQiK6aI4HYH3KXHnja+4yUYfHTznQdyOuZwOpZGUWozMIrEb/
cLKW4bS9U+FfthZd+xSGRShiwbGH85ERdRyzpqZ471Y=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 11008 )
`pragma protect data_block
IsSnCPiz81mR1shxW/6sTdcAk6IJ9jr1Fp7tocyN0EGkazgzftKffM5BO0O6d5mF
q8YJC0yA9d2BXq5GxD40JWAkFoukx2WsaVTo9fEmvCXLKXvAm/CFov3ayCFmP4Qm
apaKM7dlVpMIwXpXnWze/ePLtB6V+j7NggY3jpax9Mt7EwoJFtCFv9ImM30fG4v8
JkOEA+BPCsfUYJ6KLt/y7Iger1JtK8mIAx6yt9D8AzEaEqdtPZeN8AIEKEM10yig
AQnhzIE9yvVv2AtvpFVeMGttezZB0qhMKkj8SqwnvO4Ff8XAw7UbUTcEKdVzTUXj
NZd4qLNoMZ3DUEyxCoszmAS0aVP2H/jHb7hShknSHOEF2gQvuhxtHcuhH4Knx3qe
ljbPHYFuIo+v5YV0m4vfxs13V8hnYyrDSHQyc6TJhsvYjHz7hqSmYsktO+OjCNkU
kVB5hctFYfx/lY1AJZpU51yT+9Wx37omrcpja58vB1HK9RFwH355xwgvRIV7C5kf
N88NqFVC3DXAjmA9PdkxJ4DMPV5vD6qHYQpzP1+HF8cJV2zbrQN/zf1wblcAIBaX
n9YqdzLwG4Z96fOKursUi0/cSDO8LJ5bIr23So5cbd7snsLbFJ6MKOjaw2yyTx/c
z7aesJfuoW7QZ2SMSeLNbx96cxv2sVrsYFP2ELb+zAecEraN1ggJ9If3N/rE7Rxz
QxRw8pE019LzSgUalh261u0+pzeOTRlcE6d+LrrwjNlSESw3U9vikDa4+CoUj/P3
tiXaGPOXyK+mezeD1ZqVZmEqzbGTfRrJAR5Fbl6s34jaQzS7AGY3qCOAAcYVPC8n
iYTX9yLM+0rMNMCn7qE9JUtfXo/6viXKmzdOrmeipQ5GTwg7Q68N6fypr7NZ8WMM
8Bi/dSF0b+dNTS9TeN6FTCBsvxU8vlYpbQQgA5mn6raqsIZT8qQ3zKnBO/lPIpdv
NYQtw8cuYABWnTpZbgsnA1UsA9hbigKKfhiX40JGP7V/jMs29gPz9KBG+iNEz2W1
luBaZIUC6RqDV63OPgyKKqb88YrtXm432MO3WbIrPsupm9C8ivRkL9ZfBB/j7PPI
WtbibPeXDcMtkjY/shVU+gFiFjhamLvMFVzVoe+MCYEvekdXm+/6VIh8KCH/o2vT
HniDLmGaZvzqHPw2kaqXypPQWvzdhoXFpEalu9Ws0rEF3QfgbEWvbYlYqwPhQADp
Hj3AwkVzubVFITVjoyIOmXUQxdl57f1C/ZZLM4OX9TOI0I88DuxbeYsOH/QPXPlN
gPozHriDUs17Iun08wrGsNLkDpUgmKnTl/hdNPpCnRcmF++q+73u/xMWD4GZ36Xn
sKNEPAFj0Iksx7HkJqmyvwuAWRzLjX/9R7/3tL9lwIKFZdxjZcWglDZVw6pmIruN
G9dTG3cEvP45KxtpS9hkUK3yZ1tJsCSZa75hpElgmmejGZIHQcJ/siyBQQqS1JlC
xHgc+KAtoRfuAFjLFhXgpyo+RllsE0skUn8tpwqs+hzXu141tMt46HCXgBkS5zaW
Z19+bZ/D2ezEULHCi8UsSGEG2CW3lq1UW9LaVEVUL91NUMMpWzDdhI8N4NW/sAq0
ljEuCH2U1vAveNL7yhx6QSkkqifu6e5PWqLf/W2mOptrY+ozu7Nlqk7HfviEX482
6SK5aBNN/kBLM41LvY9ziCn/DbT6/kifArPYnQfVhErhhdc+4Be9JxkyklVZFOBJ
+Ch+bDjEYuTJYpZRC/qz9moOhWwzlP+tu7/4FRE9Sc4scQUYaz/Xtj1W/uQ+e6Z2
Wq/8Ka+rpBryrHfwRD3357itTx8p0TMvOnhs87Y4ew6OQ6SCdoiDvfOHtbT5ejXL
LCf3R1E0JznntAOofq2gIxMYWOe2xKEXLhrTEEDye2liCZEzqW9OguKa2PuyP8Mi
NBA2njihUFlfk8JIzVP0XL0sNo30D/BGpviPprgSMODlFiNNJWY6OS3EkyWmUPXT
YX5a0TNlMEqX26itgXoG0QyGR2yJcPrpZOmxuIOc3gg1sjETgnRHh084S/al7lG1
j8sSD2zw9bq71GtWFizWKBnvAEy60qJxQjHyGErSdaN6iqgNIb2Mp+q2ag9Cyvnc
4jMditfxi3Powe/6JdYhNDNhetRFbPpU/NBvXVAL6VFrTfTNkxTIWS1zhNn+6qu/
L1SGtDCdI3bOz1BXv3Qa/rxkoKTd7rQTDXl/XbkkNHhGp1hE7d/UYhBOeo3t7G4D
johcScFJ3PzZsF25YsPWfLVaERTrz2mobfQFv8+8sbmrS29u5cTuPpi/FA4Yul+n
aWklUQ3cPPsYkQyp6QFIMb2dnQh61Wv+F4cT0mmuwdupHuHz2Z0azKzcLrujt+lr
EyXfdRdcslYieAROEDui3BizrEXjyntPi3uTM/i3PcUK1DvTEJLfYfCIHVqe86s5
Vm1iwx3FiqUEimJZsHNSFC5kiIijNeeeUIkkB+y2LfZYri6d+k+H3S8Knpuu9fAf
0Ycj3QM/7rJ783lU/S2IDp7ZNYZRoO1LXZiKd0EAz9VG9T3kYQEGsGjBZsohRcYu
hLkPmX9Wbsokz4JGicXhERIF14e6ESGUkir+iiW0xX10VYpa7eOcYFmFfdncLHob
NG5iPc6AU6o1wAem80+C5/BFOVONSCcPQZ65bNoiVTerESdScDnsHRAAgYLTLcbL
NcogoWUSgFB+mYzhzQM9uMFzufcDajTcO9n/W6Knl2YwAgTP1Eoh23jqnMybc4Oq
pusYhegkyOU50t+DmOm80UWB50miedVL15rF6rKRIg5T382IY1Mu0pv9empeptDU
g7d14h9CMgWrBo0O9SxLgAa452EdI4K2bp1BNXRNnwhpgzCog07hiCdxojjw8Way
BqsulMJ9BWUAcerPhKjRc20/iQxQHgr8pkuYQxaBua5UsainSlCccIGwT+olNFCV
/fuzC2UExz6sCMG7NerHHtBzke6Kkty9P3a+0nnIrmP6btAz7kFHhUf7uQp10skw
w2D3ZR7ks2lls6halcosLEKsPhuvk/1bemuBaienrKONQHZ38arBefsFVXxGZWby
uQzKLuP+bmqOEu50hXWRGWrAnHbBT3H5sO4WkW6w8vKBCrUj+xvPjkRv8hGHA9lb
wpGjGWfhxazm4silORj1cRNAlfjta6zBv99L5jBRhqqnwbX+6BZch1+nivKfjK/S
QvHg1I6mrxsf31TtpdB6FwT4WjyIi7oVcegd87ixxqB2QdVOmQF027yA19Z6OUNr
Wk3zoWKWk+4tN0Wr0T4WYmb5WiD2tB3h+Sqn8s6BzZNeviosaxJOXa0ILR/7f0SG
mRx2ESH4kX5FFrysoN7q0ePBIGixUeFnMqQQsZKZ6c9YI8FogGwnnm/2slJmbwJj
oP4JG51iwkJHLGyForWChGTFypyJUVrn2bpCt1GpBhfThmRGzCBDhtaPaEezTM9I
WFWo6vQSqOBKBR4G0VmY7DXIkiMKNG/Smv1nWp+BG16dAlxsomITIQb3+svbhMCM
YY7KigzO6gIM/RLIUTbnR6hkKgzfCzlIWFbl6IIt5EY4rpnSaGL6WrSQwUArwHNr
ogij8gJNqG+w2pmIiObFZ/yidr6suGO2EPzLawoM5Tt3Gnt4oaDtWN9yacUzOwO0
MauYdBRPU6g083uF54F4wHdGxwMJaklIKfgLGCypCw/C7LrgVMigW6dFfMDfaJQ4
JfQDFQC+rhtaGYhUavjY84+MgYQSACV3zeVJUWf69oOtsUyJrOVs7BWspj/Q9tq+
F91C2lIFmqNWApT1Gb+dQZKySiP+rXVGzHMNvFiPw/+PknmEnVxKoEgjcGl0hu63
+sdLUxS30yS7YzagM05lgx0lgDZJWvWSlX3flpshSsIqyypYNq3fJOHlN8bUAE79
8TaQ9KYFoOdfwzST8JlHd51WoYUKHinAAiWIoF9FloPkRctLeFmDCxk8JXfFduw8
GAP11mc4ukxwWS/L6uQAsY1xQvOnMR6hQxpg8a9lGZwx5IMObGET/9MB7ANN5Pts
9F9WQ5xRQEajNPOjiKy6eA3Js8m+IZw5fp8jDtqRgvugdHIdyjSB4hiqQ5Jcvn7n
oE1jDcsn+wGjawPx2/V/XATcJl+sCykwSOg/TgA7g0ek7ZerLOFWO6qX2Aa3/vbI
q6sQ//nGvbXaAPMlMK1UHE3scFeIzqP+7IJaUY7jPS0+Ka5yyALjs0G2CWcbYeMv
gRsEB6cvGoAID7jvXyeasLolpewK45rOEM+lL5Yyl5Zwm3pvJpWrt7hUre/5sSfQ
JxzBBZt58htpDo6iC+C6nwhDd20Y02AwYUlZDHHNCYmSpHZGnBBxJgOqDADxz7br
mokkTBkialt04P3SOIa+nn8weoUdivARC4IufCsrAO1dBg4zpcksGsJJSZQTC9Un
Gt2z2oLKqc3wRbE3NTu+NaO7xs57GnRr9GmVPPJ7dGqCiLf3er88unsRu3cV3Kdg
3DlW0I/lplICpYB0eEg56WObokS7FUPtIY+ZhPg/vzmY9KBu855amioI/VblXEdW
ylbXoIdr/O5VSdVwFq2uNCibX38TQv246vBsIASOQyhwuqo8rT5RiQ/jdbn1Ex1/
DkfMRgnYThDrQ7kZox/cav+1SIc6PWg3RDxaFjMy5x35ASBeKdY5VUj1SFbIWqCq
GJiSeLn2vKZ4Bztlo4FJTtTi2tz9HnABTuZAxM6mf61CS3UxWxv2hmAegzxJNt2L
DDbOOCdCqBUdXpaaWeu/+n3b+ajVP4nCeDskFwPwr5kPENRU+HeZls+shyV4dv6N
MdSHcXqfJn+q0zr2PfMSJN82LMpniqNyurzDKx8f9CCbrA+Vyfr2kCfoljLiBUVv
qO83SmjNGX+snJATalFJnAd42mqUzjovu4CDJR+6WnTAqYtVnKqWtC/z1MXlMUUD
Ue/H10CYNrqS7skYhWR4tIUDMjtxh4NVZfQAGB9/WLeBgrVZ8Nj19o6ZfMC5C7+y
1P6zTIetEl2fiSy7c6bdGJCaD4Yj57HjKtmZeYyV3rPlxzwGtCuhcnb/TjYCB4EL
6I/Uelnkfnh5s3Yp38sePdUe75fKcSYK9iMmjg+dTTWOhQux8+1jmuO5l/W5swgN
qzanDIu7z4ehc4Lo9dJl0pztTnAvKZW5j+8arSGrOjK+VkAYMYQeLKIpbNmT7HWU
WfO55K4Guv6LBRq1YngGv1BMBeu2l4Ydz4bMhm/q3aseS8nNsNpS4GUC1viwcKVs
JG61+Wdz9eH2Ebrvp60qiVPIU/TBoKUfwZ3aJzhJwnSRUB4gAAn3fQ9lQNhWaHcN
Hjq+uphXP4/GpDlH8RPHcGVLnFnsvBLCeq4guYxzTwzVUDYovvlq7RIc8B+h+Uyp
ETfMyQh8mIWUA/zyj0tmE0VkAOeUbRSLBNmcit+V+O1KbS0jLoIEIpQ6ekocGalB
0AM5g29Pn+IxxX9Qy0BwE3KybofNA/B6O8umzbEV8aVq9wm9loDoB5s4EuqLqNWB
cAhGSnDzURFCpi36jfIr+UXGXSH5RcCDYg6xH4W6GtUdt/J7dhLH518FxwO21JJQ
bFxu3+yy4RrjvzREg9ZkCB8s+sklCGjmtTm/fPpClyH38BvinmvnI5HOCJBlPCvQ
DpgX9G7GAOy5n++11oPeBTAv7xtv/jAWzQpwnX/o9g5dIuHCTL+dlMnEKx92PVUF
5rXe0KL531CjI0qeRalfLxcarijQ+DgDMOsuVFosrd9UTclml44XROmKU8Q7riWP
9igByqSCf07Uh5ckrCknrcEdMtOrIljXIyIwnDmS5RXZCl2bPO4BpcQT8shXIVNp
xT+iEvWLm0xWNBLH/E9z4JsScF6qdff6v0aFucEL9bE6Bpz+isX8FUZVFTud17XF
uG6c7EQPZCCGbwywnvJ45YRobXAXCjNLHEPpSdV5l9AtOXxI+gFQwmJEh+o2/SvT
WZFGiwFlGNKO/rHdtGiABu9ZdpOVMEecoDQxAD+Mt/xWLWYZ9EJXCqrspV7a9HVZ
HZfJp4/QvrT397YZfJwLcJ1fUPpq4v/KPMynESm1VKfPhQN5oZCJL+xK1J/ixWiK
36lgaH5Agl3HvmOCQ0y+6rMbbIIkvQUHvdvw8aODnwVE2sx1HYcPygwztn207b07
UPvlBEJ96oFBu6RWJuCJ+dl64NT6tj0h4+dFKAEWwn7Q9n9vt/a6cOmLLkmVBGxv
qiANU7eX5BFHU5nLqhdqxrRqtY5cz4WQMMJ3g6jt7Nzubl11k4xyaexfwS8ZmYUI
sYBYGPKbj8zlsFC9KEPaB76ZUhX3FT9rQnxocTXrsxL8GbuZG5gVZxxIc/uzMQXI
/TTy8gEgvgfPPDvPM+c10TfbWYu3Rb6ngV3N0wjpAogxteTtwDz9Rq+6vSIdEKdg
xuLVDVAFCX+d1izqdnP0X1Euo04iaiAMo01a4uJN3RMwKxk9Y426KsO4/aA7MDqq
4A7J0aEl2cQnZnXYu7H7SLIYOJguyyhJfHXmAGBdV/UTiJrd3YuaNwlPuo23axBe
w2+ZgglzzgKlSp5FlC3pDRYiclEXX+q98LGtSZaL8R3A1zbPNv2qzOAWY9Lxyzen
yHNjb6VNLbtvAlLkuZOidVsmaL4EhXHH2ue2hKZ6ZIhKLOleCiQL/kMRGDRaRJkq
1pE+hjSdqN4acjG6PG6VTS4Suz1tbN4gQOa2077eYRi3TyXTk1rTxsExV2Nhp3Pf
fQ/hDpBeajsnosEqAf/g9uce2eTqD6pBaOLmqdoWiGelNL1PIaCwF2NyWx/i0AQ8
jGf4zbi1tKd133PnlrUE8grqu/WhY9LZSxEh5jhjei9vKgsOCv3oLuL0qNWSG2lG
tAur+UVpP+AAkKEPVPsDsNu3HT+QLjp6SihWSsJEhdHUP6YF6RZaUY3cuJFluQz4
e3L9ATIezbqbqT3BUphY2W7W31hEa0rlQTmyxCWQTj7UkcrkKwyd1vMRszWgR+6g
SIQNWRklfolJgs6JsCrkzSiFaQEH/yEB+S4PnFZupJnNT8dqL4L9kKxa6xm75QOw
1U35Bp2n9W4MLowZPnRHPPKmvxbXIzQjxuA1W6sZucWKqvE7injzEuFC61klHA+s
qO+TfaNF42rh1TtVW8y4DyYhUxkqiOuvULoUlNTGn7CEtew//bNxLD4psYQEHkWY
ZzU990vEw7uWZdEvpRgGmPuw7owZCdAVw/dqP6iwJHSYztG8ByqaQvi8OqU86WI2
mmEePJvqpC1LsGvgPsdz2n4d3ZN3lcu3JGEhI0m0AgeZfiZP87Cmg9fugZZ4mIhd
btS3lLDq3v+UfPOoeJZ4DxQntpnijKjgSD74RvFtxMXWRViXPwhY/YqG3ObGoNMX
KlbAnWRcVeYJAMvMS+FBMlFL/zy1R0IVDsMsa0j3mJngsNi6mJkwqMhTuCgkGAMX
LiOezibbGqJc8+CwfxwkCJq2kt1aiH3/PSFa/IYLh+sR0Gp+y5Q+XGURMabGqdrl
0iKQ0yUS/AmU23e+x3B7yNQCrsxbonX54qCjluurpaZabkS95EvQ6+DOBjqo4MGo
e44iL/bfTSDV65xiqGaxvLnvBUib0fW/SeUS0brLAI5QiLERkpigKe5p04FykV8n
2iPcPnqPvJpWvZGUK04tD3+s7V1Mm1WZfTz872WaClXzSG0V4nGUtC8xdVhrErgK
1kBlASl3fRb/KsujxNZPJiSfpi0fJCl6UJpRfCFS4Tb346rkOOteK8XbrhoKihu9
z6IwOdMDjcgdf/678ukVUoM3Jbjmli4E8XUGuSgym19B4bvRbpJ2iKY6wyYR54DS
HVV2JtvdZffZ6Ufi1ZKuxoaDx7jFsAKHevOyaeMHQJzGjmKTaAfNKAKSKkPjeY5U
AWCl2CwPHGkBDe/k0Hihtw2wA1YrmlRYrRqW76clvYT3rWuZtR6CiELmQxglF5B9
YUGciIb6WxcN5flnzsSToVfmqnjx4G8+ISw6pWM6NxWVNsNjul+bLjQ1SYzs4yun
+fd6Qm8WNUyXj8GntHuAQBbaJx24BPRpIbBdXAc0myQNoGm/LOkbNraB3jUgjCTb
kGeoqkB5x0KgxPewUoNitTnhA/x97OsiqNMlE7puhBzZwH6Shyl8qVHxD7in9WRQ
jlkL/lEreWCz7dWnIswPFhWyDb3YG3VV5rfM6eKT1hWcrY8ZfHryHPM9LhVqp9X3
5QEoRb6gPQ92OiO9HnYC0eX+tKhShdCtY/dRfpAmMj0OUBWu/U8hc7U+2XFwfLIc
VjaQGWR81m+iqD7wbl9oEUhUB4T3UVqqu2GxBzaegRhDj2aY6kgK+bNQNw2zq+LK
L7TVj2mR1Psqkg448VmNU3dS7oMGEuYN84Oc5QYsWjnqqg5zUG/5ST4HplU/IEgV
RXWo91jvHEvZ/CU769Is1DabYiiHJl+4OvIwD+pV3ibTGhCafGknmg3Fdu1kqB7A
1bwPRlHcKtYl6JGbA367Gr8WbIdPzsESP25z7yCjKqtP7DVquoRONus1GTfaX7E8
+587fptMDSUq4fQLB6qZe6kd6jspVv9OYVYYhqBe1CA+IMtf2SnDk//jgYf2jtuC
h1fX4ZHy1+Fh01YMPuyPpM8+U0iONriYNwV3McBkNm+WfUpaU8bNcjEhEOKjIB3k
KojMU7NkElwtwQSuJ2XQA0eb181XsOuk4K3b8wGPMlT07c98knZLt9vtntAB3cqs
7pi/AbXEwW9cJ5zqxEjBGvNAUHyfvRUv4AO8nNkV5AugqFSYMBxQ9rTyzWhiNKFZ
UXpNpxoWTas56yoBxxsKgiGxmTvV9Ue7kVAPYpJszIDfa8EjsCpIfBfEBASOjBYc
pRkWptcq6ondF8FbvD8dzreNCNBk4mTrPatxGrZXFxIkku6tqzK1F6TLYgaUrtNq
z5m7bigh3OHoVxr7HumH1QmvjaE2OS8/WOvOqt4Ak+JwNNtlI/vJj2ECW0zAW5r8
swaNQnIGlZW/7Wx74TarkjSxVoxslxaaf/l96bwDe+xneaO0cqZqoK2wX8AVY/f1
n89N4KA3fQkbXxC0WFeuIr7/T4koYpSvwNl4dOV+eSBm84xZp9Qlrgn9ycYA2cLX
FyiWvroqtOyfYR4VMFtqMLRJw0Trqx8an9vmJKjpowdLIV6sf8cInFCx9DyQIBy/
+3Xm+H7fr10r3uyu6y9rsF9LvJFh1ZdHUuBcnjKkm5NQIT9FyfNqMFY6vQNNXEco
JOjxL/Pa7QAfUXKux/dS4eOZ53AK1s/hpbi3ArcYOkarDsQno2hiFharfwvAVIqj
pOvOUrqIbZgU3+pjHl+GbUAwEce/kak5GhUiImNxyohHXIYSanXFxYkLIcBc5VPK
KEMk1G2ehum6/7jXo8WOKtZNM4C5AJ3jfQXt3RoCFnBQ6raZAS1tEDoPxa+RHZoV
fLTGA95nPpyOWYXY6sL+D2yluLqMMzapVFV5OsvDlFHtd4Rfor4W0awwAJbr2J9F
aUQ+JBWHBI8XO+X8PkFvNOPntNG3AOm05YgOQGUb4fIU2WMpuUO3bKhN6paDGXgc
VFV+YI7+ksFHsHeeFkCAlX/6jS9qkitTAeqKMnZz0vKb+mDWU+rrt/HcDhP+RrJ9
o8YaF+GFfNc18byvTo6GiGhTkbYCwKPMpQVxJaov/RidmXqP5YH0XKG38VMag10I
N9dOJbPqmX3ZPNJxuR3b/vdWSXt+vX+RI4zLnbbetG4nVYim/quv7xIFtj55UMfx
JQE8favKu9tyZj2ns5Nxl3gUkpLV4z+wFzWWtPKhUF5WCdxl4jFf5ApNRCDUBc5u
ZJFvELkwy8AZ7BM/eWWkqk0ETOV6KNJDUEF+XdQ2pNqpmUFr1SbLclnqqe9cuFh/
Y9xvrHRCYrsiKDCV7NvJuwHJhz9qc1JWX94bPsprXatG+o0RI7/+jzCtoffGLh3V
9nfYCYRAxdGVSBlbT6n0Yzj+ibJfh/q96ge8iSw7QuI7Zt9pRp/P0w5iCHmFsnhV
CF+/okhenQV9/vrCQ3SSvA2RHhAzr66n6/yuth4B4SheI1cfNoPH0fRYhjXJtPZ2
JTyW4T0Kn51mS923pIIj6/Al3l7ivZg33TaAeFahDjEm6OhjNXeWLUgZ1G79NByW
b5N6Qes8lRNOEsV7Ngaz2WU8cfnAD7lwmPGYP6h0wH1aDjNzfdkb2/oXCynU/l7Q
/T657TfXg6xcHMSFYrjNbwcSi3LvHjwPw0BmJlhPRgIo4GMvoIlUnobYXhKWytfP
9zujZgqCLZvIVBg/aLH4FUclNaO6n9N7Ga19b2Jg5vt7QcSW8vD+3UngZnUn+ZXk
uUFGfUlnuXyGN5qjQr829xYorqLy2oryOCrhY7WKQsbYtFWNqQV3vpxmYQIbyZrL
+T9bzmPvep5Y9W5xZXOCATfD7bYkB2H5de3Uuj8GuxjJB0V9ug8n0A2nENBeNRLz
IFM05LJJwhQSeshvH6h51qme/C9MbBV6gZn5WnnQGn7WIWupGu1Q9dOnoPoBOBrj
tlUqExf5DL/tO8CM43Ixgdo/a8pByqUUysNBznDpy6ocBZatj03am9NAi18Ibt54
CTrEtc8jbzocb/j0Qk9H3ucaliV0nCyF2A513ON0WHIuXukPb7aPRPoiAH7jYUR8
51eWoeBhy5BkgAPY3xajjAVoWPVir0a4H8pSrOIFwyp//S30dhajIbsfODHLqset
GOY23Izn3SmP1bwZpvwwuGV6sg4uw5qoFQoVdrDP05GdKu7nRj/rfnHq4C9sEpBz
vaW6Da2/VzRzExh6Pq12goGcDqHBJL/yeRawy8E0RxCg93mG23Z4gaQK3CkuA2QW
v4uA6GeVjDvwhtsiyGLGNmgtomaPx3pRC83Mxf7hVp01wJi/KoXg0bmB2NskmMpg
ROs54/iiIBuZjp40Wu6s3wxUk44gX1XqyOum05LMs135h6GZQjG8Q5AJoKZD3/J2
7eJ4HUh3Fvj9FscmZuZ6tYRb2M0ZQ9NcjPcSXT7nzNh6EdHqnZqqHFHdjf36EFbw
GHKyKyhesbA+j6swWs+zg6WYBca/EEkPmuPmFYcZWNdMGMxYwmOUyMgLt1UkUBT8
3gniGWP8ayVgSFEzjgAlSLtAWz6C6dqgTQvoolhMup1U7bkIf/aphpz9oeweh/bp
PMxopkoTvIzoiYiPBoBjPU19rd9xvVSFm9Z4ckXZmThaqJEWmDvE11BfpYw29Cuk
706o7HipLYGk9DFheVs7C+/HW86ZR7Nb1+T6uU0egycIhUD4FOopgj7uJ7GJCMRs
ORCvc/e7ZnAY9MMmlHigydcCPLoc4AjpseZl7f5rb3mpI/BpISVBCS1435EyF60t
BaDH7K4zZ+y7oegTQYQwy7L1ueKxsGBk3i2ciZOB0YEdSJoblSXvaaBp3UtV7ycV
hdUgZrdNvruKODahSAloX2f7600zfIx4KG1tqLZokFWKxH2scPETSoaIXtsxROUS
UhDaxYemqz5FxAGbHIJl1dHASQ8bDGFCcxH17m9jFGKfaX7mwGBegUQbu5i3k/NR
WAZ/k/yHfj8wPt4BdSeY9JMxFfxgUdS3fCLhN5fgJY/uj/eVDKib3oXGELhRppIH
fiSMfKCuwTeNQ7DW79j9GO1vdPCkDgAji38l1VQws72v4NTvX09PNQm2xKZ6DqBM
9krwp7E9pUCWaJIYCczGWSfq5okPaeE3QhRUzdC8Q997dCCXppitnqIdAU2DRvSl
L5YaRxsTY2muKpDlE99lX1diS3In7ryBbkiYasIvMTi/hgZtXTPe3sjNEP7MkLrv
/D6dAxbovNcDqWtD4LqRuR8IerAtuUZrhrMjd9qHm4tE7LGuK872qP5MnQmf/ba4
mOa8qmLSyzzcTgXlMqt7k+6JyeVtLX21BbklJ/GDCG+kYj53rN1Z4ogioHKkzqHY
GZ8ykx5OOS3dXOp1TLj0wmvbAVeZUsrJIXsyKylDN1E81tUsxmYDPehpYfA4PAq/
d8mpn1Ht8juWL6t/20RQl/NzuIKRXX79Dtx9UJIEqQTHUKz6bocw/+dHmYGCxN5m
ra/mev9GBqsho3qw1uWJzx1BACChPRGTMZfMLIqQ2zu1MSnUprohkSA43f5rAEdq
q2YQPXLQp/vVcPVy0hTkTiLHODTn/shFdBTmU2joj/BpMlDopqQBV1n+fTq/u3Pz
tQcVkOeOnydftbMNKu15RosWRbhXoq5omQjZxqakCsL9Lx/R1ALmLQkest99X8Zp
sPEBbLZggfG4RTLAAcSwAl36CLasd8/xdEVJuwJJdm9Oc48HgiuOeSbzRmU57rGa
fSytODv3cSZfiFBefLWfxVKXg3QbpnkTgYpOi7Ne/Z/vbx4cQm4nk31Kk8MBR3U8
T4yLXdZQvMqPyO1BY3trwzYU3XYUgIiU8KgxWiOBDq1NVip5llztOhGO18RI2S9t
U76DvAqXigqi85M5yVZ5ugyFTHD00nD2x88xbbiu+kyESlLOJMdVa9io3ZltG/di
c2qXIYmu8oorc5ophu3H//UkSjX+h4urk4sYZULTQk8NVwKeToTaDLQnXNaHZvr7
cLmdorKHgz0hvnptLeVRikHbNMm3IEpk+qd08vd+iuHreXRM8HSbA97rNa3/Ogkj
PoWLfHmjq7ji3a9m6x2nM3mzoT/5CNWIcs750WWHAHUMJ8Q9yAE5nxBLWDICVZMP
BLnCN+iF2uoNog/2DVakUI9JFToYfvEP8JA8b1VkLbMcsKgaTbbb2QMLAISfs7M+
SVM0xKGpGmeOXhk2iNLu+dV95GvjDK/TfrByo1R4isO51DZZdKO36iyVrtlTdXRe
C7ygHatjSUx7QOJODbt+7s8qzrEkOGpmsHBC1CAciRyL8h42L8eUovmphnoJgDvj
LsDUj4B4rqva7VTlYqTn8/3RCyQwW9MmKoHCOr0X2pSKWpsc51IGjy1SuzYc70EV
dDchnJiscATS1sa1PnGQdSPoMsgQPFv22mFxdcgwDuqtP8IYz42r/3gedv+LqYbv
o8bPFzthKiLZ42uMulPpNbXYnK7Vtegy5WMGs5TSvYrQGXW2ootJsCdvGw+tMe5c
sSjAXEJAY/aA8nk3yVfhj85ak3Yf38lFJ6k84Ws4jDBU67AJln3D5VM/p7jyBX7p
oP17+QqlUw6bEumUVbWMkofs5t9LkN2u8bO7zUZmUCBGQlE635DlPk5y7+1oiI91
F1vcCLcmXwVlV61uRTHuMgley/ODxPZ4J1NI4XFiFMP9XxHUBV1eZkE3tybwFaHr
/qZh5TPehK8BVjwHM1iC7UaO7TCZttrgjjM59h3rK9UkkitH2oix12ICI4C0fAPA
73BQsM20eP9yfMNfyU1HpvYNJIKi1AIwsl+kGfvimz9hjs8YPMmehBhMqOqPwK/T
uqth/sKKyA/KuTSZgog+mY6laJ6632rMd2hicK7NQY4lJZ8AXVY47rAchvHGWPej
ZNSDyeQgWGnrrrc1e6+1v2fcWCmbTkGYzIfkppA5CpIL2ToACnkmdURI/vqLSm/x
mtgstmg/7QYIST9zD6SIBI89MBVz6JbxxTBGIhzJiEdloQugYQ9jSpXvYI0f82pJ
D0ydzYVlppvMgRU23AZifWtpZ46nHg/IfZ7bJ0sJsvZRSWNmTOijib5PlTyeK+So
FVAvAyGoN3YtT+cfYsTveyn8/Ce+aM9INkP+xdSc7v/RkAkH3X3G+AvMNmDfvneQ
8PIqm5PnKXSP1gbBW8Dack/gw2UChIRTPYyenhsiymaR2mZRBKGOMe4ij4oq4Gi2
lypmynLGhh7I0LIzrCJxGn9uvmpW+qh1rXtMJJOcZi6Bg0vM/s//l2z3ZtGMn02X
pdWRuP7z9THSSoYJH0OZCxE2E/LAatVftVi1XzzbZD2+vV4GhORRTvc3TBUwbbgP
BnxRe0T2Plx6xyE1aaxIPO8UyJOYwdLfyUQvT6ooMsw+0GgsudLiprLtpUZHc3iT
2zaKkaV9OxckfnDImIvIeDUiYezQKErIIoDky6hRNNs9sprd8Dir9dai9RHyGPa0
Ld+Rh0nzFb6q2On2ax+YbFbSo8oVKJ6hCjiOzcyoKwjCzK14ygSEvY5NFvadhbj8
FSSbyYy6RDbd37aWk2hjDP/yBm2Yz0/rX7YaOZILuU96MVws5hVWf6yJsOaY5dPu
huHIRGBCuTbygQ//2FOcVT+z2f8Oq+vRz78X5CL+KPMR36BM7o4Ju1d2oXjJZb7u
YfIxtlWolIRTYXIrNN/4+/F+Io+nsulfArry0uslVpTpj8aJVK9hutd1nRORNcND
eiU67XIk0eLz2I3/vzimlGq9jwgothWJMlR2NgK/ZEj8H5sYuhFBB0KzySC20pvV
I4rp0CDMDvw7449z7nB4AnseORJiidpyTU9OWzvB4ip5K9/XvU0whVutqGupa5wn
aLiHnasEAKY0mZgQnIaJjY8DOG4uigMKfYw9IQcuWb5Cn4NS0Z7/W/SRbglcOcdH
Gzx+dKQrs36h7kxtHBnwItFlTE0Yp/nG1myHtqVU1RbtOgNKqDrRXnJ2f2eFIk2F
vwLCQ2u4wX7y8vXTN+TvKrSSGtFkZ77xPgU6NpT0Jtvuk6GFVRpzw0LTw3Yzu0vP
ueTalZD/dwp5kE1kjA4GA6gF6p7EeUfvcZsr1e53cQzf1cZGFIi0TLQzeO29dVP2
q+lYsklX+E+UxCQB3RTmig==

`pragma protect end_protected
