// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
OELnjnhAzQG6uK61WMhR+lrlLnIhJliGFfRiYUZoZvxAaG2EYxPmjhWYpX7lleL/
m5pKW3jhaT368RZuCC+UPRe3dSBX+C7ZwvXQ9FslBeX9yMjTlHt2OPbDyB2H0bJP
nRGBmZ6LFAwW+bwDptrpkSulNe1yOn8Y8Kp0YXya6vO0il4CItZtLA==
//pragma protect end_key_block
//pragma protect digest_block
O+RthcCYn9CBHSZKeacOcEgPnto=
//pragma protect end_digest_block
//pragma protect data_block
KFzsj/i3myDs5aAguu8BMHcsStcUhHZL7mmn89HwNjcAxHUZ1HQwPX2B3TIkmYPD
mPin9rN8MMPWxodq+2lHn8ho+EMY5IJMkqJ2pTH8FcOk6tcqinrReN5jCuYA/YFy
rwsSDNavdhgIVWHXoSn+UKvwWgT5jenY2TLnpT02ShGY/+DO8EBwuMRRbFnyIfBL
pWJ+Tx3UcPnab0pGppM8SL7Z/BD6TNi5bP+O/HrGrVV2DH/hfpFtBxuvZSQrA0II
tSMpgiQ3dc3+RPdbDT0w5tNuwzrnA8BPSY97qccKcO6zYyNh9uUDdcpHlcxfm7SK
Zvi7tppZyAUIW+6fZx873QUKdhzIJd9K1k4jCpEej6iJrda6++qptdxTPGrPWzUC
5CiErc+/saZ+0zutHFqdYHfYgHr5r5xX9RRO1Qs/06gPkAiR0gX7lDqcv+gvtmGm
yzKUAprfhV0BgrdnCiJYDjXnkLxvLN/XKh8w/rctCM4IzTJj8k8V6qjmwU2nhWsF
eIQ76pbYVaw6FdP1BffPlR5G8zVX5Z/WnRamlbQiZkJRFOQOd4cyKNWn7T4L64KE
hk4TB4XHW6NpUrQ4qrvd88ZSyg/254adZOy9QyKB3oildV3ibUOfhkg92bqNbN8n
OePGBs1f3Wst5hm+2HJGfWemjLIquZjvO0O5zC79Nmub+T/3XtxkuG1fx6TPJM2q
cR+nQ7Kzl9pfshOXEBvrCABDLexkCiutOx7XApeMiyVTJqVfbWqkRyhiVleNJMl3
MvlfyFdNjzdLEg0j096V3YONuSEAlyGXdLB4BHBvWw5NSz4UJJG5NBSlGxxviwOh
LUAtzb+4yNAu/kbbxy7RgRgXe8hQu2t2pILcp3fAuIR4Wddlj9ba+X1Mr2ZbDtgs
2QnelCtlzxKmei30zB+8JYA3BapDKTEv++Kar8+QsgKQzJNycQc+u8qIAWv0yFPS
pxHSfPYsTcV+5P1JZIXzje6DHz7E+u7xnX/GgAhDGlXwmvDj2ZQu2TCjQdAKbRUE
IqSTBn9VHG0C7jAv04OmTyju/ZVJrdEiIv3AlzodF8UEDQx45+e5grPtQ8QIzImd
JDltpLGpz8I8ol7R789Ui/rUOPpNX36jYpSkIEM4IspZOTROPqAIxROerhuQKpKl
RVlWs57eP1fevkWhUiZs8IGSF/bPNXE4cHHPeWd0qV8cDW7yeuSpFV2/PshjMhs7
r8tHCk/o6bszNAL/ceM6neyI1q2b8Gr6WCaXBAyrUY1Eyxnbda0gW3eNgnQWRP7U
/44+sjWEOQ6MHv9NxNLJ/cv49wTQ+YShUbfSRTVeY99jbaZ5tv6C9AryJnD7+TGP
pV5Qxqlnx6Spebkxd/Pd8Fc6fbsV8sg+aLB2yVWuFkvkQNITWoUqTXs4BUMwlt0H
8Yj39SUSl1MMkqRC3H//Cpd1A0NyVdNMnKIhtKnHc58abf/bP+RI16bZd7O2XFmp
3uALVrUnWPdQK7492Hgn4iihKrCPOa7PjwadGzOfoiqebvVyso5RhK/6kMtt/a07
r+tv6qFRNJG/5BaCtUcMZBJrCPeS2fT22Eev8B8gOIjK11V5pzTKGuZPYTYVzgEC
rOOh03Dez2Q5jMliTcxCZCqML6m3sUUK+xjV8YdPvPZYTiy2iObhwN+52k4lrbZj
jKb3GceLo5eWVXDXw6WjZSsiHULyGKyHvckfiFUqNBDJ2Cs7SmxwFH0XwfgEPGNx
iHTp4RTvLOaPyr97Xrc1rHQwcLNqIbdu3WuaCpJCeTn5bpn3OoIqZf89T2NdcCcF
YSX2wB+Klapq+XMCF6eb8pKwvvVmoQg5ZSyxFM0XVv1K32hB2bE1BTKb1gcWVUDr
3N2jGAE6aJi5SnDw8/SWmn98/aW+ZyoOCUcIOOn81HZ+4pjMhh+wVNLxybCsxtAG
dP+LntlF+yYaHrkSarvruJMyb7GwiXyLw/0zkP+3Dl3hhIx8U4jUsy/y2cdWZdmB
/yBwBtDs4EkcrQXZ6p09Dc7vrv+5RaVIWk5IOfK2SRhWRqCiP+peh5wH88KrWlee
v+LoBz+4DVi9rZZdgVuUo/mKR03m4oRAo4j2gUlIbW4P4mwoBmpPLQ/LYKdgxMQs
Os8KjZBEGX8P5hbw93fCth9ErmPELuruDftHZuCSSsidd6LZVu5Yyk8aLlQUwAZz
wnySMrpG+2UiN4fZAlFfx0YkuE6yHjlvEZg9hcZVK3oBp95wq2DSUBjbR5N1U0Bp
NQsLtJatojKFO2w6SscjTNu9qkoct8QsIdAv1BDc3YWWRW05ptyhhhi9uFkl/fkJ
rzVhsPMx6pGqySpfpNeh0ps8Bdu5SZIKa+SyOovJteHRQOlT+ocsly/VMOwhzOuT
htTSp7t49IGq5bPLiYOYqr98EkRXqvkSpNdbZeaIAO6hphl1s8rE6A/d+EEwWBpH
PLGQt7GBwhEKyo6FHvaIQ34QU08hCSDFq2Ju8nyokn60iZc1YFe8yJFZVhlUNMXl
mYhBCxE3Nrsu6kIGCFGB7ezFRJGJtp6/FeG1OWJYgJpxhdEQYRcz8wsU22mDbieX
kQVNdZBu7KeiCZmAtpnPQwNAce4ULTbjYg/PHUe3LuEh6B3Z8RnQ28l0jiujPUmI
XmWT7o+ARrqwvFBz3SrMOYJXS1QZ0pATvSq54xFR23AUQ4N44/s3Ez44vZeqdMLp
wvoJwGC+/WzMGdgXO4AmBAdKFRjclS0nAeLBQPQu+oSSXTR1SxcIvBbe5gkbMpcj
h5XRHvAkWXe4n1cXKz9T/QaBlAUt+7NR2+F5g63+JavmjB/FSOnyimPYPER6y7Nf
mb8GQtyhCByMXOgKRS2FqyYsK/pcL987cGfhjaEbSR33BvUbkYBpghJkrTP8+4RM
TrRrmkbvQgCXQ+FEzwOTHOnCq5Mgj/5cjwXT1h/Lh84yATL+qOyVMGKi1Arx8ZGD
fNO8gk6A5sf6mkCDtlGM/+kwl2GOi8K9ifNVh/ok/PQTA8GLqA0DbjrfU4z99nL9
Bx/aYZlaFDbMfY0cAYUvUtjsbpx0Bs+Y7Agie2xBPVxXPo/Vi8gCNed/IKHcJgI/
EpRU2U4qo8t3Xitr2IlYhuk24ktvUKS0WksP6mXbdZeSkz5rjMZi3YxoTAsph/R2
hFDwwtZiEJ3eNkyIlLl1YErtqBqRP8oCQg9GMZbpZMiObRm389zbavYuE9amx9gr
OlLbq+TOm4S1Vd1hiOs5QTF9qv8RxzNTJyowbriC/IobllsARkh+eyWJ6ZN7b4a3
7uLvXH42hTj1YmPn6BW8eOy5jJt1yirGii5/vSB6WHIbkKLgZiQF9jgeKkAW8SqI
5/0LVJZHfAx/cuWnvNu8oTKX0qfYlFnyAXsVL5llqt15e+LhXB3wwn+JE0qHLgvE
p51xywdQBHGxzHIZGX24tjW/tEBJ0uc+x0vxn4kq/ckb+vq60kbZw+59fQtfFJ1Y
6wZuUKEA3Sehd1N8NZ/1u5m4jnFdUjZ/1QjAfxl762kB9QtXidfdZ7F+Lzi7cGzD
8exJCZ4hweBqFzhtWZ6jK38rikUw32idOQ7jS6APuVla13IBvvQ5nIS95TDDSqJ8
w5uYPAx4fO2533AO8mUCBT38wIW9qMrGPjNs82aXof5CfzB4TCYL0hKoWtVDNGGe
Fi0043YDAaIWLKUL7Qh690+w+q5tLdCZFPKXuvzr9BdJfZzvTZvIZnLSwy8dejwt
u01Kfrep30Wn1VCttwXo/qsWNe9yQ87/tDA7zUOY2biZr55HoOOPz9cFkWiJ54Rc
M4Wxckna+yL2LP7mYe4NbZjblqwqLHHwhbiDM5gyQA/ZN5U0SxeGiepBuIv7wdrA
/e7T+13v2QdZoJ+1rTWzJ3D/LO1BRiGAONymBGZ13jqZGwD+N+HfD72ZWpr+kP+3
AkjJTSWN7b+Fxqpl5rHdTstTn62lEEnZ20pOVgjRREzVAtOzkEnVVhnbWDyUhIZn
FmB7LUAg+dUYz/bUpyJOyHwkUmd8QQOWy9/qEbJndLdzzXy6eIumxFZ+4vJwxu/F
FQmpIK+ijCLW8aHvh4l3O+Do4/Dw8BpDLvsU2gSj9zQ8nHiAeaoYoOxBPXKVDMdh
6FqdOKwIW49j8bgIXIuhkB4n3NcF2Ee4U0MlG0q7KUMQo2I/Pdmm7w+EOAm6AHri
DcgHfoiWRAT3n21MLC14LmB8x2apAmwMTWCvVTNCAOmE9bVWwqQ8opyCWJjRPVhZ
FNDU29gZZ5AfaLrBH+TuUJ7j1GjZgdVfuO/k9dtsUHy6VMPI9A9924h5pT6rq5t3
ZAtBu4LpZ0q77Gd9w80eNKYrTOxMBXnrUKBRRqZPie1W5nsJugGjqc/SASS3dDJu
GgnKR+1MNcDmfDz/yqATeEhJyacFCuIzMPYsYeZ44Vo0xTxc9d2obBsKYdILM0VB
GuipZuSxQmuetitqBhCVOA8PcglYZJ7bTABAboyGUcQk5gQGy8NpFC20P52rlGvy
A3TbNuT49eshYY87y4U+MC1azJU0k8xtFfPI9HS/Aq126EEChdQwHuNMe6xqYjlu
PPSyHpCJbFqIjMJ1fK4Aswg8rK15K02GLU/vGZ9fH84Uemn3MDwEaIjq1S0Lm0w0
LryI6Lzce4Ao3iPAkeXR0AHQnTlOiv/MajQ48GpMuYIKnXowbrtwLTl7gDHFOyJL
K/h9Z5e0PYzsc3xxsMHUGeTx81Pg7PWyVWYrF2/ph9SXmHrsEXTIRAF1oSYWjm95
OEMi2dMpyFNvOCO8r8p8I1Vt7TGJggRyXGH86CjrWaecBURI4eROlVhanK8541GI
Q0j7os8kCHujNT52/nJNP6BQGl3XmMjcKuVkv32U1GmR65jQfMtkIeEBmp1y77LJ
5O2+dRiEZtnEUksC2L+dn/DHiUCYAuw4r2ZvsCxT53GuvM7QFmVk4hMdkktTZRU3
q2/qn/R4dE8BT4tHC5T9h4/wH1TeBa4e3+aKa0J9KDqMzFM5Nsr202/H3Jfj8tMW
IvcNvv0l2GrUZqcIUZ7Eu+dWwY00TneRqubfO9xgxJkdwWVAeVdoVbmZuXa4rGpn
Vdnny5+384IBwZsp2nGOXcqP3P85JMaYByHo5t5bhEPz77xqaV4du0pQdbGK+5Nr
y1DQ+WX9F5W5aJI4HRUGj7a6V5I3ptX7ibpch/hS+oE2n92YQ/AyBYjBULpV/Ttk
rj2R05bxtLCk+LXpYdpUfJZ9GPXbKFKeIpD51LQ7bUS3rB1EyWyHRICS/KjmMcMI
Td5OMEeWr+FbcZLlXqa7sgNTv0DROj/IgrI+pKbWAyrOqGZOxKKE1NaJVuYhSsPv
BX9CHsYHQjTDeV16wolKOXhwbqZcnVa00jpS0UWu56zrjLed7rMZBcETVybPv4rs
V09S20wsGQRkDy/E29glZ1YjVCdKGZEHnavPwCAi/luOIUKBwVp9IqbIRB2TXXju
INnNNE+8H0fj1Egzn20VznQzAgv5mQ2McPKF83GSLFSFhpo64Cv3iyMVnbQvfBOi
zjgNnzJi2ucJw1CzY+4op56LvAPWLBO8msu6L5zy+HsnoO3R8iQF3sQ7gSOrn5OQ
tp3ais+T1NsOyx+pkpGWHsvrg9z4xUq48+qDz1FfqQz43igJawjSR8Zf9CIpKlGX
7/1PgAEZn5QOJfGTyNTOQYp4WOYvMTpcwskwdhUEQrTVh92fssaUokLiPtb9ao0O
hRQ6+5y/iCRsn6F+HopV2VhXzUZaC+MeqW6mJkma7rVvHQBczgk3qIf1ueV2c3QX
QhvUL5f/v6rphJs53vSiAMA257/7jb4jUIUfKzSq+GVf/W/qirjPxeIDjU1VX65H
OWaZ1nlHwoyEwChgKr24wFzSIP8eduqXgqw30PGVxuFqRelw9YOVzv6H4GuvlHM+
rGTa1qTglNtPU4qjAB81fim00hooENhYNcojGpdyKFqmiMR4IV/f/MWDA8iXDsBc
rBREwZP9Sy8nngLnsgMp5EshLP8G1lmtttn+Tc/so63aU9zVGq1UCvB98nDYqr2Q
UHk319iN64JjoPbNAYps5T/UpbSmKSxPWTSOlK44tMqtofk3eDLQ9xwYsAlunNs/
O8njIhJhWw+UaDN7Tk7Hku80bEitkC3tJJ4NSfkXeMHQvkvHqAG8GkbKs6966LsL
Th0iyISyKc9D81ZmInOxu4ou7oYwAZeZQA1Rvs6x0xh330XuER55IBs4u7Wtr0Yn
iJ4aI1NDgYU1Vzmbgl1pnQhu2hVWhqJtU8Cl3UjwiGy++bBYOzkr3o6Rv0UDOtrJ
O8w2qEnWilwyhwjh7HJ9OHfcSV7EjuC66KEMz1hZqVMS9mvUlfV6I1ZZjkcl3JJZ
CvJhN4IO/ybahPpwbVLmhhaFmKPKjzFTKybquuuHxZGPNttxv0J2DEIkPq+4cX08
uXIlnUZYqX/XgQIttO3cXKS3aOg5EG1BSLbKYwCGLExBPyMLfkgWTgvG/npfWMRx
+qNDFry3wdeUXuBTitsE3pfbqfjnsofs0dx5IRU0yhKPwH5BpPMp+GWpCzGLwVBz
5hFeeuEiXTfWs7Q8V3wTh3d1xf9Q6J8+uJPPgl764TU+zU33935DTu68k7ZOO5DF
ZjbJrK7Y1IyW92DYb7lXamAP7OrnarUDqKTWQijRisJHD7Zr1rg5YFhVtaZEPIKc
Pklfq1Gq0JOyxriyLacpA4+mK9hHvK3/BShaXQ9F7LKZtmUI3QjN3dfuLB6hmbPz
iWt5YhX/NsR8lZvMFr2di3XjehYRsthJGfTKVJvN6Vf5Nh5iOFVRavDK+3oWf7b+
LmwvFTnqgFrgGd0UI9Fm6rubg7TBGRrjf/0/ash+YjCI6+x1UTmYBdBuZ6d1hmj2
3pH3vpIr50doriPb5EdzekSK7r3SO+LMEbKUaO7sQgEupvHwMkDJ28CdtSTRh/nj
dn5lhj4d+lQ8KIc1Gzw9G9AD4DX3quMHy/yLXoTN4ud+kk51FrjgIf7waYiRGc4e
yirWdL/9X0OZeGGm3Y2CbB28rJmTvHLZ/UiwDuwdYzHVdlI44GmeEcUArOG52JDV
r0O9bquXKsBJLBvef36kdiZ1tvKT8Vjc473eiZwwiCwfZqyt4BFFma8UuypzmkE2
dPpJTnaMH+z343Lof+m3ji6TbjoziINga/jgsYOnnJD6Y1pkjTI++ggnEAWGpOa2
/9/1hVWftPCEBF0vYeuy77VhfCaGH9HJm10yRL8ihnjadmyMTbfu6V8q9FK+Inix
A/JpN1XgW2Ip0vUX5IF1Ut//NyZnp+pzg905dgk6e5GgAOBZGLIGOCj4zPbk3jb9
eY1PrpdAr+9VbYimJzxtfiLa3VeeDpJAy6zvNY02Jxtpj7R7W5E3/2e4IqNGmhai
vJ09fuFiNuwVtX8l+uNmCikEqgS0KMHLDFKJsFXE7SyqfIZAW1HaoNHAzfx33qrW
YhWvLvW0NtkP7kmsD+Cg6lwcE2K8VJuoSM3ArsAWWiDIRY1QYOX1V2/JKcePswb/
hjQMccVqJHtvvpx+9Y5T2tQ0y9xLEy27QTjBHbw9m5rbxaK69jecYY3Kfo8zHG97
cW5POO6KJfY8Tq4BEU3APto2D4IkAOsppJn2I4/Pd0+3m09ntFM/3UNZwQjoisXC
P0NdqNG5GCitpjDZfrpr0OP7FNMehqr8IHA9WNCHHyrqqJ7ea4I9jQDnLry5lk7v
Y7jQPkC5VA6mEBbp3P3dwsxkmFe3lU213nk6rJklLqFcVKmOGzHRgK9YraB2o5Ek
xMlrcYyVeFE3cPILldVRIRVPXQC61UzKo8ne7rf8tb1GpgAvKw/2DABVkbEnI5hw
jcmtFHsDcB1q1QSDM3EBFGGl11HkpK1X85kUgwTiCGIANXJJSzuxVqLbGtWKsRF9
X8TCRm0uHy5qq/Jyh4QWuYbeD1o1WDARZwuhpfC79fuGsIAOzhD/8fkyq/ipPj0m
K9rHgl6hsNimuKsbEybI4VTZGxwtc7KVce68PJ3Js/EQ9yun54u8bLgbQSHGNxeN
fxyGTjyulMgcJIAiIfJwSuIqoYKPq8/himJCCasPsh6DicuiAjW/v9VuXJDuWANC
KPsQHCtYRFLdMGTNFpGECGS8weRYdu+Xg89JLsaBKt0tmmK55ZRL9QTp8pPqF80U
zCDlAyL/cmady2eOqrodHpYTl/GCo0wZMoHZ0lgAIXUib/yijp/zjIsx9AOwCQol
zMMS7f27uIq+guYHhG4ACQ==
//pragma protect end_data_block
//pragma protect digest_block
dGzwmMA1qrmH0BjvX43VHGXN7R8=
//pragma protect end_digest_block
//pragma protect end_protected
