`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
VeGbhIcAwafpvsESWcbRQnZGiq0LzONdtZqbpbUXumY1n9qN28jnqREY2a6grlyJ
el6U0XTMt5N2lHiwj+EwL+eljpVWLPWY3yt9PQSuLpVe35U4QaC9J2o65d7h50jz
qo4QJWJnWvhCbu2+bTQ2xk3tZYMSv9O6xZx0vZ8vnsU=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 99888), data_block
vI+gEWqAKuyrC5lmxbCyd1FnrEs8pB44q72qZCQ8WeXkCQdp6bg6q4T12WGwE1tL
XEQLa9afD9bpPM7y6dyZF8iLM90uSOuULVxnn5IZ8PxkYT9BwU9C5DTTS5E3HZWg
mSJKf3IFZMD9XvV/R+HcMYdFYamCLNBnAtuuSGlwTkj017K90fxnrk/H3iJZF+Cs
N641El7igJo7P2omvUpQAxG9WLkOooWVfC8m9pKi0/GWuucgTMDBxrd4dTM18s2p
DDS0Sq7cBa0g3QWgY5fselHlHE1bPmK+s7BUCIb8ZOZ4ZRPcffAx0nHWYt9rqVZc
znHapPgoBZ4+UYw7Vg7IxLaPyHDXJ33nO6txUU/WHe19/RllpfjU/731omP2o94j
TGY5iMgKiKdJRmgM5KElM0YkHjMmy8FrRZOiS2DT1F31WWdmvy8v3dIxSnB/hbwV
x+BR/IeWqt+cGdGW0c93puOv39uSaTshoDJzFsBNDFSGJyQHPlnpBzJqtN63K3im
TLQKDNuFbOwMihp00O5PJT1DKhi54LLsFNemjmL4Et8kSJDO6qBH4wjyUUsGhqCA
1UOwlORpZTIg155UjDmjJNyqDv95G263Nw1NbVwG/g3bmCtjHO2103kpyKJY4dNi
USnwROusnDx2kxFumh9dPRXaJCs4zMuABmqKe/haiv0sffFGoQbt3+7O9GrxmEnX
IgrJoIZW7USSLUiNQ1VCQoEnLiX80+pSLEfUKZ6B6AM5OzbuLYX+em3p7jIRWs4e
0fxTvJCuTKF0KwqV9P6dnD7Y/6dtPhDSxZL21C0j8Kfs4gNuFKkK61YsJhbDTfCx
KG1+hBky94/+5MPUSDFO/gkpDDgkx4QXx8jFkTFsSbBMJMziT8LF3DB4pnY/nznk
FOpYMJXFq+QwhIbv3mFbcGWpuGPSGWfjLC4TF1C/RoIUoJi7IkBigCk1hTBYLVXy
ZFY2Kf5SHZZ7zmlxVrmBjmCFHauCXu821m721IihERvDX8LHKP25pGf1NWyZ88JW
mquZ389eDGVFdVLGIVO7QtyftnfgSwUkK7ynebZtDZ1oc++Ut1Lt5vqUBKtBpj2o
jzORWotcgA/IlMN2xvT+CqgU4a0USkzdQCA0flmJCS3Ik33B6HLGPcxlBuencdym
NeyRCPre0bqx7ER4yXCAvx0ihcZ+NkGbi6MiRl2MrVK26Omev64KJEGhSzb2gFhD
yD+jCWw83ni7yOkVZSqVUtmg/wW3fxAq3g3ZHlJsiZl9E2TDFr2mscBU0TIf7K34
7CG8Aj8XbiITxcM5uIe5Ag2IF2iukozHN0do16cRa7XeZuNFEkRKMXndJZ6Sy1JB
em4qts1/6kM5raWyoaNtDmXMdrhzadye+3Vp6K0/XYSKOFPIB2tj9kxOTWIZBjDB
DLLP2OjRxbUULeUO4tt3dOOU1jSzEKhZP0+HCUk+rxj1UZ/yJki4NWTigRNO5Rqj
FbZe7EXKCvaonqDpsA4O2ZUbbSQ0mrwp8wZqqW1JQ8NQfWM7k5YfDhyipI7GRnfV
nm4OosHji9XLT1EG0rSv9sDxyfwpYPC+q+2oLwJzrZrLAr6hf34yEjHNPCb/9MMy
5CB26TSmRj6ryj8iD1SEUKPAJyK9f9pujLogmftl3agVU6tRQ9dzwN5n6uXaiWPf
0BnnIxpg8Cf+2LnYLtQWtCmW1g1iG/Xm9SdiEox0zzmcf1dE1M7Gch9dFwHq1Cjw
B9nEil9YZ90gmowjmsYPkVwRJw3Ysvw3KlJqlmOJe8oSB2wMA74YFRQbN3UjHhm9
rrm1GL+HghtkND/4ly8ByjY7mbf6oJxMdbDqD0fIC5i6qRlzUDyrmCXEzyPWLXeT
rLTjYiREMQWLL7LXz61Ev6VqZ64XexkcK8gDhTi+/YTGkdIoafVQPIcnNQNzdV54
L1OIHRe1C8qWk6DCx0bZr8r/FHhxnFRyQbKsNmXTCRhXbTdp+TTR45vYs9QpLWir
txfqjJiZE+73uyWU7Eu+WTIyL74u+0upAZ+sjofpvrO6yEyFgVwUEqbIc+GBbUl0
tf5oAGsAs24KW8s1XbkggRAf+bjNDpV9GGEleRy3iHhs/d+ARzODSarhFVBkV1do
zxxsEZU4RZu43VPhHyvbZqVZ4POn86KRrvKLgrK/FEppL4MFzqWL7LJYsLp7uYpj
sR/vDGdgZm1Xcu40/Rzc6gS1dFWbL3s9df8L5pWA6j+WmCvU3P9AdNAwGVy9Oq9r
dq66tFt9YcPw3yUsBhwZkwmKV/xhADRKOKFkYscq7NgXAAlUlV3VKGf/m38z210/
178/wo/apWASftXmkQp1fte5/8vYaMjxMwIY9TfP61JBHaAVjJZR4yAlKbfeuwgv
GFyIfIxD6fyz6x+hKZqMp3VnleTcYxg6U7OfpFq2y9++Qlys87dD01cF6fYd62J4
c6p4cufAbcGg6TQ/5MCuk8ibFmZZpN+vziqzB8PzgiesIIYVeU2C7/ZXoDtX/j37
4oeI5JE7JbXNxwRLSAtXFhAa+iCW6lM6xm0kWCTaE1HDmXKsK5Byu+jGKFU1vCU2
WmPz8r1drpwwLjR1jopUOipGBULCSsUDf52ZaepJxZbHgMcy9w1P97ylou5rme1v
8MrYVP0aanYuEvqkUfl5olT5Rl2gBrb8+PApdEMp/9Q/CCnD9G3yewMfeh60J7TB
zVsYJ088DMVJSgaqkq75PXA/fad2kGmUxYI+DK32+mdHdrn5u0duPiBbX5YqAKN5
t0eoCFqbXKwD5yaMaAOnHOCf74mMmX08kGw4RMZFSs+qcU0DMvwZ8zqrdv99CFZT
y/CtbF3an4w6Eg8sEm5fGhw1DZbd1tFyECVafRksb3YW34slO+rF3zBzbA3qVbFW
PhqwU2BC5kLHfs0xvRN76/quRlXzroG4zqjOnSPZcB0Pq5aO5F8M9L5GN8GNZAwD
LbpdEEfLMYpGnIZbuPTAKRn4zQCliSWBUWksjNz5QWo7RwaqqzQ3NE9xP8F3uoyG
Fyh81qeIIrKnEVcgwVLrxHvGZZpIQxzriBKJho8Ioy2ft6WPE9bSQqu6PNL3Wtp+
NQp+pdTztWd3Za8aEIS5Lwi9v4PJOy8dOg070/DgHdM9QAzKTLx9sPGXh1hTDLk6
fpIkCxi2P8ppOymuPyvZA5VsGJOn6ePTtmzZbbwRT4/b+GnsrotW7BKfD6RTmY0J
rjA9+2PMzrarCbXldr0DRcZlYOibXMJM/H4a+JIUU810eYrwcjq14R2sYT4lWZZR
A1LvvJMPjE6w1nPGG2i6NuCMdO4/A3tIff1Xg3oDoxIGb/hi0BsUVxLFhB/DaYC6
kbcU39f3apBbn1KHdJoNf3hXX5GG5CwSz+4THQQ7YZ6t3Ygua8N4DDJ4d3V9nESH
49XJBIrQNKhJ1NMISzeVh+zTvNBdmKkHNYc/EWphjztx5SVY/p4LeZArtURkggXO
OjaD2bsoDiffu9aGdAVxyM9wLjUFMZw4vM8ePUSUWH7oUXMhZpSoHbQBrPpwaw68
0IPG+xZm+Ptj4fNbnycaJ8GTpwfu0u42F+7hUJfh2x74AQnsRstj15W0S80khKJA
4+BXY3QhhkkiESf/jEsuzmRExg+eEOaws+BfoEt+ZAyGHBbNn+SuSfrO9iyU04Wn
HhuhYsj7fh2NvuOrUBRMMOQ/RXFtdU2JBZPjWKVLWJh2bEdsaDGOQAUFWBmQKKIN
uwON6syl5SMEYP5DgfQ2FMVglKjknZAkKfFooF92IxkP4cFOBItBX6LN/im9lyhJ
1kQqHIkgslE4g0DaxonHehnQTHTWB1yUYQQ5lbmhQ/Xzk5tpdRJQYqOBD4ND+yHA
ljaB4W00xmvCot+PEm9iWs23Cb5xJ18a39RpVKaCjSz9nx8zmrLSJLIZ4CUokhCy
qwZObMBdHFv7Z8aEPLX734CZfobOJ2cYIuctsdB8RIV3eWnVtEBvImPL9hMMym9i
JeNwLNcjELyi10ZVaoBFYr8yq3k6LofYsXSiLKHcBQg/qZSdlbgzcYXZHZ4AfiJz
qDkv8kH6f7YllZPeNB/aebuiaCTEe8KTM56M7+irgkXqdhLfiT3RQH1fyvUGbdmS
KJKFNElabGMJAjM6TAUlEhUyIKBIgPBy5sQ4ReKI+UAVp7V+UtWOlW/4Vf+j4cqe
0ZT9ODcVH8obZonwoZY3pr9fcIhGhefxSof2zz7+J6Zz0S3tsufi42bP61+dMPw+
tuQSbE2AX4TuhoKK6FNYKYA+AzfWNAOVf0iTo3uYeF5GNuDV//19ma9c3k/Z5req
hbfSltXxXo5HSB8Rwx8+kPWEuqXokK8Nv4Tt7lBFU2WuuSzXzn8GMbWoLFi0oJFI
axOSU7eWxCw1DWHupjD0XiSptum4Yw0xBtzL402x+vklCgGvA3XjhO6A4e6R76Y4
cnLy2wtbRQ1CwcnHZ6RvmXput5CUuAvlrWnKnYK7z/Py/W20lu8qeYFQLmt1183k
pJvNOqjdC5vEhEngOSZ4T3BgbPg84yEQZqs85MQA9zNwDO4CBLR2gHjGtEGGpvN+
S59n5xXRHKvPaiT4aPXiVYWF5dZNK/UVIalxwlZZmI6K1/PnUVodkUjH5NDCILa3
xhbqdfgre+N2X157kiQYp+JtmawX47EiZH8Nlh1LgjxLJAlD16SjOr3sFek9l3MY
dfn9xbTCAG+SNS97BJ4jqCTqhnL1p6qNvhkypdM+zO5k5TLlHTtNIN0LidlKcHXH
oxA4vwS8N/r6oumr/3JXP2nmVWGXPF6xpzBv/vmIDAE1QmF/HuAc+bpTiiWGb7t2
+8+XtMsDJ8cN43BmepH5F8FO+smRV8aSYZv6lv6HkyOY0z9NVroGNyMiEkWplj4m
KY22Vn6us7sVJPABs4Vb180sLGfteDIotGVWijkt/5TxcMjY7b59D4QlwfGc5OaL
GT9N0q4Xm8tlgLX1MsZkYZxKoOqkp3yPPqIP0HwD6NP2LzEpUbqa8PjjxrXmp8aK
D/ywK+D75AGnkHoNaeDoT8iSYlEQko9S7Ot0KC1UPuWy4abBZE892pwhc8AvVCH0
+wA+FoM0ohwwcEQKoJHoE8Z9nARdynipfPwZ5XGRbF93tfO7hg+X661fmUB1gY5I
mOxtysl9r0WqFxWfqfyLonk5x0UoVY85e9QpJ50qtUmoAFP9lZujLvq2e3OpQBe3
ZZ937l6qZH6/rDjYqD+DDvuGT5FBcC5F7JFSsOoOUuyl3qoN1v25dDKeEqO4uikq
ed9k7y9JqNP1wdmVyolxygtDwfUTurlrCs7pfaJqpvDNfz5EvANkGRNTUxhjN0vw
yOJCeNgZDIIVo+AWY+iElvu/VenYB57CqbCgVznfkAUBHgC8nDq4+rIUEtH/dJoC
eEsyyKPc2I6INtVK7ukG6gi7Q/zC7rqgSY2GjupXYfxhOl8c+mNJQ8WlDrM1Y8jP
ZlJEYPL118ErAzRZ+u173QKUJDjyieravBglz65ZW210PCXgt9XoyqIG9ctOUXR/
zU0zZ0tcIRFIrvrbDo4ApDQjMXahRe2rZCSeV5XO3/5zTs0IAgLuyh8DbZcm+/Gt
lpFbA5BQl0xwHD6qaLUq0vFouEAqq/FsK9DJK0z4kBMJh11iMeJyAwpPQCj8ouiQ
PsIP1yQx1TcCidvo7oZjPrMRF+s0+0DYOJlLoBjgPjcV9hwMpUmKLXJpYSZGmoEL
FIbdWA+mC75rThgW+9rmVYjNiCvOzgJTzHIQ9HKPrJbVZjqQgaLmZWdu16VfBmtf
dLSpuieTcAlh3lQcIBiP/LUAjo7H7UwdgMAn4JJgK30hO/mm7ZjBR4Eg4J8jH8Xa
/f7de+nz6mMb82gC6S+JzqTG7meUv7lkuUk6m4vaX5wFDgG+7QjoT7iki3AfN9OZ
v/HOUrBtQKSxWz+mKqpENwmyQF7qG1ygeuA1IK7awpxfUdxXxWwZq2H1YhxLt3ep
lF2En+yyZPk7LL0Park6rcIbhlU7REr6+zTkRDjbsgX0XCPnEp/yZ/lutqUu2VrZ
fzSH7p/py3f5tx277BsylPPvJrhow6CHnDnTzLeyviIkeMJmc4Dn0XAct+hqw9yW
CUphUVRA/hiT5n3QshbXE0RhhqE5MFwanBpsBYdg3eIxeIjnxCVmpCY29uriYCUf
1MbT1dk1+FG4n0oQtyz7RFu0zCyQgBJFn1Bp3eyxv5muhb7MTZgnYoGWIN3mH3oX
gQrtmnjZbcbo/tPxEJoAEdoPFFS2TvqoP5ECL3vqnARjfsBf1L7ny5+gbiT0vYqR
KP4i4ZusSOKvgn4fBgyjI2UPGtSKLFkiNvs1XNxV+bb2CGXUoYQByLGuRB7s9Ix7
TAA0c0vj5ayjeBWO8FtL99xg3V7X3FyNYCsOg+DYrk9ZP1T0ZG1OghtOGJ36LUn0
LsXwDNy3Opa/mnxl2QdW0kTHvgCMTNnJoFQjLLvx33/JP/wP1FyvEnn5U9VyWUq7
iAIcI1b6PoVh7BdfImUPU+KLxAd09JHXFw9nDAOLilKJnkaVRie0rDlilR0XK0Kn
lNxwfGBCBuGyVY3w7Dd+f2d11yZIg8eEBthVUVcXn3/WMzI4oB6qmxtH/13hO7GF
5pVcINdvjB4tD0Q9zNq01+E7Dow1rkII5lyM//XeLdjaokXLVeu5K51TE/ssvCGY
jyZbNkLcnSzyYZ//7XqBJ6F7Lwxsza/ZCnOF9aJ/DLzLpILixi/OaIFJ6V+lyeOP
cGq39PxG15VmOHbfzPLsHf0m3d2n80SReNceVD9hQFToKl5BJOko9MF2f1n/ufW6
mF15Qv2Mk7Uro9HlU6NNgDw1xjykOvCuL1ZRk9AhF4LJ71kDtWhB2KDQj+o5ll6g
ynYGRn2wRspB2Lieiw9C1YOkkj/xFmBXLGqlKdBRS6tC/ccD8FcoSDYrPbvYwv9u
QF8x9h0DmM929BBmvoIqEfEkiu/bpeLBKkuZ8+F9ALvVmV1hiMtrT6ZUigTeFmOq
TL4yQerOyfVvXYMBHg9dsUzKvPp7qP0fKGM8ZGsx8BXxZfl9cGWtmlXiFOp2RmEn
DdlPUCOaNEDt6Y4KUE8CxrhwjCSAt1p1Kb18hnCEYekJxE1JNg71JJyMpTzMWbRs
V5r/CzdeC5g7kU9zrqDPuc+458IXJdTv+acpZQ3Jp0I6QcJlx0YCm45cpoeo7AdA
K+QRenuEEq6bVXb2r0ZzAQaP7+yZ4F82eCVSYbOF9rOzXnbQzE/0upvhLhBrYig6
LwAzeRXMLJE1+2TwIUgRjLCEx4JuuwOOemR1eAK99Bv2WpjpiJuyLv18XbMGkbL/
q55Ra3NTXr+xddHergWdWqR051p5lCKyD6IjqR2AC/BIYHFRJIrAliPc+9fyhkyT
3W0UFQy/QieID+NswEdjtNwuBetF7j3raWJ0fhotoGyUVH5FZuMD3qD2Cg4kpN7L
39XmpFdHGxrECuP74gKa98QC7vI/CHuIhjjE8/FHg+ejVZAmk8/b9DyCf5xrZr0D
CV1zGmKLyD9Fud64UGpN+VqBFtR3uMxq4xytbg2FclOL2Uh2P317c9azjJGg5M9J
CN3hf4m4FV09UbpPFdUzmOf9gWy+A9UMyyK1TZ5cuqDyJnQurQCj5AlFr4an9swV
81IEZcTvvVm5xe5WkwebpXhW8bP4NedcESbmuynfzCJP94DLQ4OhgpWO7jYc29dd
jQd7Qx619UhVzruAWytHKqmBxw3CR7JPmCG5NEDdv7GgtEj7g2w5ifl44y5w8WHK
uV1C+Xz4OA5+5lISY4GwKgEhQMHppTwAIEElZhZA3HoN2ihdWjNbNxZD4o3Fr1Zv
KKuVC8nycj1PjapMUQ1dE0GgCz6IkQDUQKq4NG+v3pwbmCrKce7X8NhFhe77Bab5
01AF+0K5dlf++AYNSYm51QOjwcD+oaaUe5oEC4gmFI65fkH/JUdB4dii4HEQuJY7
dc6ExqLFSCWgaI+C16BOdAz9rk38DlfuUGBWBVuXB++zlXCYzGQN36rMXhjtGiWX
cJ7o9sF71lDM4x3ML1rmSXJS/XznpR74/Zi/v+JmoUdeLAcwimLLf4moxRl2/Nvc
J+sB/MstxDpO5CSqK++YliPOJ305nHp1DLE8k3Df9WqsUarANJwLn1te+rJBsDmD
fj6AD8Lpg9NtcsZleDc5k2rOmo8tt7qc3Ijvea3H8P/ua/NF//NnMb3lrcEUGJxE
t0G/lyqKdzUq5N/2iYJv4quLODwK2gu9xfKnPKYE33+VIGTGb8CBdEuZl2FSgk52
yaJ7XqG56hNGvHSXc89yZa8RqGLVqhRVs9CgrzMmCcY7pYAQ2JSAYutUYILp5ju6
KbLEAeHDHXl5PSlJyDOHMWPgAc8dyeRh78oeHR7istSevWP1LxoskM1IMpnoV9MW
2cCJXqZUGBJDiPG8lsmQbDwVvaP9xx/ObwAfSx9Asqhpi+u3qxLNplcg1t2xu1qS
fD+pJnG3pw6uVRXDK7hBKPfAjoSC/02roIrGGT+/6v5R00FebJCx1yhmrL0w2+to
pqEfzQ4SC9XUC//30mdl1a4XA1O4r/DhL/vewJ7o3cuuwiR/r5TewRN9y8fYdNbJ
vpCpvlnN5k3d2PCcVeXcuhtChOLm/WKyRjdKo03ZixonR8HlNoaBWKPNQfQLJj1h
qt9vIQaO7hbaozdKmNjNKGxAkL5edw5PJmaAjs4X+w+geaZ5/fBSjpeVx8Opv13n
Xc/SR432qYI3szFNv6FXcgCP+/HbSAafxsWHAmKOUicvzMaia5+6fTKsHKlOyTaI
MTZVvYiSw/mKYGGnYFjpWL4H9Wn/MVv9EgeOrQuIXDhv0nXLhmM9Urq0Eiqay4ew
9AZgu38scb5+ogG2Eb9VptQpWgke7LTdyPNx+EJT45We/5HZoyaRA7Q2S5jxb8te
acv8mcQ4vOr7/ILrbTophtXgWvk3Q+TE2ozUK2SL7/RZ1cKJIHomdEycwAtVxr3E
2GrJOdwIcXrFqNNuCaih2rUUH+TtB+m4H+OZYjZRHiJB8F9PWrIZIDz6eM9Xkwhr
0ZHjizC4a/pwN5tNRJB1XqBKZVspmc40AjV60LpXggj7nZQMvSqSRbEAVvmKJXEb
wjhn70/LuBAa6qLyLagHPv3ENHomCV8HRPe+lpaOomsBqgU6bRhyTHq1iz8ln9wa
m3RowC0Y/Vhpey+lODVvN8tS7WL4rfxozyjlt3mEtyhsbOVZT06YzuIXMa5RITv9
XQ4HTvmyVxm2ts/04o2rKrH1L19rVMUfrPsdyIhYVppPwL8+hej9J4TM0HVHjCQJ
v1K9xPVehiK1R4r0A6kTC2tGIGEEkOf42jUQS8mVUMQM7X0XyTWFJhz4XGrHe1cJ
MHa4zws9wbtWAZOszwVDxPuDTgY4rlWHUjaE+/i7lEXXbEVjEqHJQs7Uf++6yDic
SRdzgxcYn2aoMu/u8y3TXG9sOA36m8BRifIZtiC0/p9h79ZD5+p0bdIsEOXEP0/Y
4tUf+c2f5RreUfQ2jOgoLr8wk6l1C4NtajBu7Rlv3tfwzXeMkL3ta95n5OcMS+Qt
d2CjoJIF/m1MxK0EjoInxnRqgNpTuIgigptdz/osJzqTpvO5mGn0IlDueKUBl7Xg
ex6ff1TQs0KQ8/FZykviaFFpVeA34l7UOBgoepTBhb6o19SOlQOrfPn8BU24sY7a
WMgyV1jKuCqQM4CAnatWcm1OSlQrEp1nmviPtllNTvM1vBQdg9nSEFcDOuAiLq9Z
AnVX2vc73WF+iVEvjWnaKywP6ezR+PbXEUOn8WOAnuca9pXs8hAbmEb5/v3qpNT7
J/R/9Md6l3NZKdzmOT/d7GkeqQUmotJHGme3dduBqX/UhH5XEzSEEVgTZFJhCat9
0HSyyKoeVc3hq8wcqDYuKgYeEosxohnTTT/GqL/JySFHMRcTAwwitkmqb2Tug37r
9pUJcbH8QKdc7XfSYEoXkMvoIEQUGkTzvsbqF46n373lP9M9cn+DemAm1VPuWnT8
ELchE9QTwpYtdBnyNipBY89tZc2tedCAXi0Fts2FnnSiQcdG8MHufZu6NCrzN9il
yX7qsuSbTDZMpI3YUuQkiS1P7wvZTVhAlYqM/Jh3fQIKmksA06X4wDrzc3n9hyxM
MXdnHL+K/Fzeq/69OxY9Vm2YAwARhF/m5VNqapHtj2hT9XmGlsz+4OTMuEop0ns2
DN3Z0SfIiG0kiPK4S5fY0bgv0erpxPXCPtrKu1GDa2iO7wUndFCMfhzW73hf5FJS
Zu+l8AXbBP/QPN8AupJM+wSUBCPJCFDXBKGNfsuMH1qgXJnJ7pnbNVmFZRWJsxQ2
QZgtjw4JdszoVDZXdmAohOsCTnLShmfy6P+qCAVTrw39K8/WblRc5v0LghNwssju
/106PxzNXbBoUljRsRSqdGTT3vENm6Z0CMzi3imptAkUgBY0Kk1hrAJEc3FnkhCE
KeJ3Z3iGMPDrUWpYOppo/qZ07JGsYudBKa9bPXt2HodF41E7bEdZyanfYdr2nkmV
mOwX22l0tpkXIsI1z8CCvzgWM7nShmwJoc1K+aTnVFkzHWUS4yQuifhb3pDnZQfo
qzJfwcqliZHrSvE0HnOifs7ktRoAs0wGCFGu0jxHL6kg7QwSQl98z4kPdhOsF9wN
bIiMrlWPw3TgEKfYeQmjHRZqFG8UDGVwIFrLdsNfA2F+Z4YdVRpwapcGBtNOYshJ
BtXfgEFCWpYyiSSr6Q6/JzvRUD5Q05gve4CD9FtAcxFslka1UBa/O9XwyOmLUf2u
6hG9zH6qWNYP7DXtmbXpcfXKSXJoWEE1gxFkKoxyXZYTc2CI8O4cnsqbrWQkDbVN
k5Z24nI9amAaSKvXthQbGt0CmSbN/zjCoNSUY52kMYqyavK0oQsdutt7gKJ5TdFV
gJ8m4ISk+SAOncbJ/hAqWyGYNCsueTRL9Vj/ag9yiKUrAGaB/qlPgFKUlBKCmFMF
JtIN1yl2NV5rhBPO38xmVWSZOvzHEV8b9jfN0r8IEP1Ba9O3z6nweJNCAjmGCEJR
yFAXO73e+f+Zlcezzn/ZbOKc9BNf0J3OGirJ74LzVAiw1F9x+PaZYxm1UXTp9Vir
8csS6rDZJNaVmndAXszJ/bsGnjK/P5pxVyFpgoNGPMygHa9Gkf7/ZOKK/MyKsDGl
QkZvX+gW8xdWkDp2AkYfLNvCA/dPZPKJMY+9JS0x6rMlJIwiX/wmn2hlNWs9WaOG
KfEuWUWwWIEpMyd75jlyjHJeKHGb+wpTqjtiRVAM6dixo0r65VhahEK60l+NjUZt
A/9pxc3uDqXi0Q4MF9J+Yj4r8oUgXvIbqb6sdYCzkmfCQ91E5A8y7YpwE7SqU5O5
1EXev2Bb7+DIJhnguvx3MIrCpbwXBpsodN58C42vt2LIxGNiE7PBZzuOfCEU1LV+
mhQ70cdxjtlRvmiEdzJpkqE6LKjrYBPh2qndCD1wZv6rh9tEi9u2+w6zg1DsKFDn
UBMo1segB44OZ+4USWpS/JrhWFfkwHhS/lpiuqf1nFRnSlCX2/9Y1/vDCtxrjCd0
NwH6H2IVcZSfnNdyT5IBudSP/iXd9C0Z6QKs9ezvpb4PffdBWEX7FnL/eM40rD+m
aFCbNZKKhdvRJYuowZl7zmMHmjwmQN9H6VGX2baRxbDo+Sc6uIB+NH1EmZuoMi0J
CE369blAvaw9cduxn+MK7xZk/vOpDu77yZuF9r5Bxe3ZAiNWWzkh2abmTJ7IetXj
Z4GXVYKrBHwz31T4l1DE5IkaoYK+dcSCI+oB1LDJRUGFthml3vXycYAGR1pL3bda
388TdXYX8Xq3GSaRfSCDeCUst3BsFIk1VeRaZwEd8zcONYLwtnIZfdMMiHWvO7nl
4g3rqSaTScRGsWRodmelJOEJQCFYQxvEy2wXHLydihJrDHwSLPTrcE9HmamvF4lo
oxGAtkACIKgSg2f5FZS/sO6iNgaSgsYx2beUBm/aNeD79R93J0/xY6fo+Z4omLEb
bll8OnMIl7ysBF+ZXRijThwlKikl84yujid7AhSz7VADOG9t3s7/8UXWrXxzDMQz
pa9ALw04NZjPObWjOsux2QPgNWeRALlnwBZ1SScWX8US7+7m9LE5yl7qwIqsqqMI
iL8ScDtipmGcS7uzhnOi+V+nBXcdQRaPX9IaHZ8tATrB8KtvXXVPvko1aP750HhJ
60/+4gwXfRp2aruIstNJiIiX26eNDN4O43gA9zNO5UmhwIMU7sPByjSOrV+D59qC
55vscBsR0hxAQDM7FPTuuE+KygnmQzm+y/YHh+DJJVekNFNYAyI+jlJESn/YTd+c
ldZ0lRRD2qHd07eaInTKcCkLSbBWaS4Wd4rZYaChy9gG8IlD7H4LeXb4p/0N6DgV
W/Lgi/r/S0JmmcUDUlLtZhGezHoNR3vhob5l3kwijhYL7+FuCJt/wdpgEnteaVA1
9UC6YFIc0kYutuFpidK9f13FhemcQIxc+jwmSvH3KR0ZROsE3husDdPHFxDTPFAX
e8lgkMy+YVxjfq5RhxeRNtCJl8eyBz+RxONrYabCRNVbZHljWKVn3SE9u4buy97D
Xw1Ux30VHhayH/yhsG1jhH1T92T5ql3WmY1nf5OyyoYxDN5lXJqL9mZkGPXD1m8p
C0T/c4kVI2pezEzL9Wtn2auLAxDZc0JORsuAEYaU32thhOq/wSJB2HRejP6dxB7F
5ZfZ3JrAIAoouWhj725x52qpB6QpwFDyndLz5IZ8K0l9ZkSFkbwYee5qBGv9miwu
y+M0RrD0uj51Xkkt2yTIdsUDkCfAZygXGVuk0tl/p6kSkHcspocan5xpSFLix3gI
cG13ky/plIEBNMeXuTzcC7gmZ+EpBvHaLcmQqkJftb1qufAr4ZHskgiaptkY6YyQ
D9mQ6QTxlN6aFtI243tnQ+FpTce0hSna4Qy+pe+o27Ecx+zdh48qwUQlCnn4hidr
yyT1va8JG7CC3QdWci6yT7JMSDwE3/VY29c0A423+Ru2EYNN9qt2xjEKuXxElu3H
Fg3hRY5aU/5FWMhYuCs4U5eRAwDN+fiIZK4Mzntv46uBPv3x6rKCNRNC2PYKbK3Z
wlme6pR5PXr96vU4hn8ZY1dGevSAJagy/fAkZJ1vgJMu8cx8Mul4vwVO8LCQroTq
xVVs3z3/tBXc5wqx4Jk9Xn8DDAVpQCrIh191xwuM5JYTLClCoWPF6gQdy05/wPgg
coIYwost3VA0CldOlEkKvTBsiSUo/XEWI8pzjwlnjVPJt6a8I+5ltN8aeG1BE2nY
6+q8FESWQg/2RvfFjLvykrfYht/nkJC4epd32tJtyF9lMTXwUmJnEPUxUnq/9Qg3
RkeRAbCjyPwvaG8jFk3BprBV7Jix7oU5mwToGZlDQVAG2NufivQac2kdwScFjk8X
x2e79io5KFiVbBRnjkfd//EVr63oOagF9E9r7JclJ3alQwe69Ik1X067s+N5TbuJ
PJ1DS4J4Gl9pfAHDQhKV7iSQQM7eU/p+TYgvd+qWKTXxEovFwk+zWmaZccpeSsTG
O1zpeEPQTgf7XdYXLLhb1KdfS8hCnds+BT0tKwNkDbjR9biqgyLe3/kX97KEXpDb
zdYvK4A1zXJx5xXjyNsNlC8lnBiuLRWNqTxWwvqY5VgSBBle55l+Ph/KtVxWvJHF
w9muCVIPL9NY+Ql+uTIubHegKIX3okIet41kmaAcwqvWiqOPlwf9BqUSoaAxp8/n
Xpc/S+G0dRjsoVjW6SlNLafiTtwfI97P9z6gv7NN6eZVTkHUz3biiASM4tmB0naM
9/pb7Q3Iajf/pmGZPnTKFmax+NN8eBeb3apLeIfDRVR7Q2bDmqLbRpRBNljEV5jl
AGJJnFBBQQsbbiK+3PC4U3jG3lns4h/3XLfyHtVH0WDFII3Ry2QWrULti/vzbRaO
spGgbUAlKFu3HDJi+c6toUwESxXolmbURw8JMXnZ0VmhTtZqF6Sz6rzfxs69ZO7H
V5s0UIK2Nu3t3RPSkddtvkNmoU9vPxdmv/MeJt2JHRJ9cVJ/UBVo6x+lyLExZWQ7
O8O4rgi2h+4kmZis8fECQECAjAkrdlOegdtpr7JQk7DdsYv9o4sczZQ/0DfTNnfz
kYdfuHJlwgcFvZkMBdJ53d7kPzHRqojRl94tQKbF3yejAAhy7/M5g/7OnIPXrRa5
i6mLDiR1fIBeGUewT/g0UhHFvKMmvm7gSv79V+TTMaE8sqRn8THu5pN4V2wJ4Ahn
VLlFaQChXd5Ag7fRU4vKtrcQAYeia9ulwyrtj/LCvI2Aj1FRvSEs4wE34lGmsH8/
GBCOJBScvrKtrNJhfHqE5DcGqXnkIamK/l09kDRZczcsPpyRBgX69lRQyut07wns
MzMNAaZXYxNL6yFui/m/XLmsK2oUHr1NlRkGJ+7KCbhUJUIrDtmxkM6du8Bja0v3
/IWpwVErOTsj9pIanizF3YIObZ+t0CCXiBBnTVfKfBwtJVibmNlbAsD4xwIkaubG
kiyaMrXxhos0o3sxjYoU94u1r09wctTypqyiNkd4x2o/sYoF1ykvqbKeR2q62th5
8QEF7TVrJPBthJYmh/zovKgxUk64csbJxnBUbsmWQKRzqpXAV13oTI+MsVhDFVgn
V5m+K+qn4c+wdjuGRKyOnLIuotR/GSBLiv30tFwlCmJVTGlYCjT3bvMjJiasxfWF
mE96d0Q0ac/lkCxqunCusLE/q87UWX45B49Tcgjw9fNoz/eQ7KKcDtYrLMquwRgs
ju3L6EIwOc0cyq8H7ATHLNlsmSy4RHLGyxEzOTZQjnh8O2jFPzb2Lm3VXdGqGnbU
yKG6a2Zdr1mHd6Nx5eBbrJ7+MU+tEpHoRtGJu9RmK/vfda/pn9awYZUz6ERqrq0w
hkjQx19jv6LSsbwiO2l/IS7FnaZsX0CpG/jf7Z1AQDGuk0RevM6Ug4DwMfFwqmra
6gtAR4wQ5jyfeSehOGPSPXTSYJP7s7lhtggWsd0Ib4WXtxsXxx6T+3cLQkCxt2Kw
guXZcbsTG9/E+yaxa+XwmIAAK14rDcK83M0cwhKX9qGQLe2Z1FRfozB+WW+JKzeE
A+oYMhjETrtjYti1AJYVubattTbzk6Gxx/bo2bPGw723PXxyeJ4K9B4vOXbeQ6PT
MiCMcxRKuJSn0Jt6l7jR/wCueAdtsXS+WBHbHlw506hrSK7xoFtGiXiLFcTz1UXZ
+qvFsMuf612CYNyZ6/cTecfcKXd48kd5Vz6JmnxAw+gihe8W5jkYpy3gvPUMq1SY
bmeiDDkC+bQi5xW3eQ17npKPrSixXWGW5MSVLXsrjKi7iTNjSB7ypYDtNWazV5yo
TxoPr4BBVxHPDN0jJ5fGS4WBzCUpnX0jA+8i//COEqjgzvsjZJlkdwW5CGWfa5Qw
hOmR08vdwIEPlrZhyFI/Hb39h0vnv+8N1kBuaICHsMRornNE+sBwOKaIdCi3EDw+
rbFrdbKscmRoljbwL7w0z5Tj3kgY+AstNyIyi6IEoYwrmxRwMNhejetxHmN7Zc/n
d4SdBZ8oBrVWu0wOSvf13kFpfoqJnNHcEOy28icIC6kdR9Qerw5eIFFB9xNKgZKX
62TR4MzJtSOcvItu48utkoW7GqfQE9j3AFnrd2EX93ba8zv6CDulOwRU1yBAsMXk
MOA3nVrhLCmKk5XHkh9pMtWcWdiycwr9H0WG4dtHfX55BDI0GTG1/N1M54yRpbM4
HUy1a0U5VSdg1IBUNl3OFZKG7fzD9GSvjdse1dY8FPv6774QXOcycJVaZ3zm3CmP
9VpVm5yyGLtC/vtjQ1c1S4rGGX61Rh/sNcCQ7hYNcgX/TvICF6h/uFa5a9vl6dXA
sRrVndAbwp6WTZX32VpQzRKYpuYzAwPqP2nRBbNMc96vA5se+ghiO7D315W0qiQi
4HWGacaCzs9lb3Y8wwJB80Od5XoxfImYSPO1Iwvnqa9x+/uHISh973V9ewJKv3jy
4bTWgeZ0jzBSxm2E7zFgMaKVLnqkLuUkFkPnq0SeYp7eexzvHb2odF7vDuOY8hhP
BhM9NPHEpeNFS1G2FaIk8DZkysF/8ivvSt4xRN4gzILLYBuaoAGbAGigK1ffbjX1
PNFoip+nfBJhj7P+PCqM3f29CszN4qytZjbzZHg44SGqX1T0qTwMnVQa4MBht9TH
4e7cJGWBNQxfgae1yI8m8clmNPx3TRZoZACGrerK/li0mhTDShGLN/TqiBymuYFl
26UY8/k79M2048ElVttHDHde72wULY1G7TfGOfGAlCrc3AaBQpHd6BUV2bD08OPa
UNCNBZwEybSKouzTU7QEbNj9HjT4VAuTNJ7e8oeQBEd+g6F8IR1jz3MMwwE61Vza
9oKpuVkRcGpx9tJYDMZQANMVXjVque/8AahIf1jQOR8QhK6XgWtBH7NVT3jL7NKm
UXX67QG6sdH/yAu1qZ61iv4HeaJcRMqYr0b2OVhEMpt2h62UZ9INcKrXA0tdwNWZ
Ci1oqDYQ0YIZry/EbkEA9DK1pFUg+DuHEMKZVd0KEk45S6G2v0GmhgDS0n5OEq+/
aq9SOsRjt/SRESMEB/hpGNmhp+tBSVGM/oc4qYueibTnsSHypC+cbqefjZfopg2t
Vju5v4ZNOBoiQ+gWeLxoM3b627pixDE+nFHZyw9RGMH5P5maDA3Y/OUWFM1O5pC6
zXJIZPT4jeCJpvuA0P6y9pvcbgTAZgKlUhZLStRHDO1tge7+tFTsOZXXS/9SyvYB
1TqhqMGBYCVfGDwQ67kXFOkhOmK4vCRT72KMb+18eZV7NfgGnQXLP6wIJsneX+TP
17Ri3oKAqFceohsaOWG+wdktGPfYqsMHs3O9CfU6PVFoSuB3nc1U4yoAJ3acBGka
3C3Dr4pRbF4gStdqJnBB+PSCRH4GRTecco0XlYfRautztoEOfqOeJRlXYxU3PGbL
HxE7JSpKKcWmZfBgaECNL1tE0ouRicug8BjiTaIcfG7SJZf80+xlyl+z8eacqM4B
a9LKF6WlaykjVd9jDNwfD/yV/GpHvhLpZTkjZ62W9FiysKKh1Sh3YmGmIgQ4gxKk
ECPIot0TmzrMHvK9RpQrMdfDY5+idsPozjvEZrrGVxT7q0llyadS3GL2tGTa9039
Xpfr83kfcX04x7wwb8IzGoIUzdcRGbAvMzsLwP/HqUlTw9Rr+8bbNtOcyrRg3h9o
hlSLra38Jg+6yNLrvngH7Rz0eMPVMfLn4+MAPOlcVH0JvlJ8U1I6JlaDrZ4SmgqJ
TzWX6eKcKrYKMzmzVVzTa+1aACYNCFoL4ZrBKNjvBS95BCjjUKtDhVhEDzPTTz3n
8lLNz1QFD8q57hFg9VxJXpgSKYZvFIW7ZzB2hp80iQeUHS75q3TWo81zz/ckANhR
Jai77ZCt7IbDmdRJAxtzU1cDHjue4EE1Sb/BUeKS/d988sojNxasVEN/VbA20PYI
ISQkZN5JlEgsskeAN8J48CgK1Oj7cJNrMEm/KQGudNPwltPGNxZmqH6osAhpCLyv
dKL5OovLnfnoYAPAG0qrZzcq9nGTnS3zkJ6AqM+PlWwCk3H6Wl6YssbiFB4vmRH7
vDccN5KSXCMbIINtex2TMer8/pK4SjTBZrg3Fktb6rGZASpQmBfseD8pENlvswhw
mc2sZCSDwiZVQk3eDY686IYiym9VDQRxoCoN8PZziqoWvVyK5f/t6vWRovsU1MSe
f66m7lobcH1p02t1v/yAOav41Y4Tt/WhsdQQt0gDRnhdIeVGmnkeZkjpFQ+qtI7G
B/Gmo+JfllW4FJrTqRV2HcqYXHJOeU8v8QxvWHvJd07PI9ntOqM2Zu/55YNnVzFs
iNkzGz6Pt8USRnlxUr/BnKc5weY49qPCcZciTe2kYi3WBTLWiK+cBGlfP6gQ0rMn
wm2NZjtel88sG+DHt4P/krv3j4ez22PFbCN3DA7NvDncImewFyVtSFDTYh0ZbWFe
4TOUHzhvoxdSCrdS3Qy99sX5NMpC7ixd9UySl9AHwJHtaWdbQzUkt+gC+0TSJvUb
oJhvdwTV7Rg7tzRBKiboYCegAlOFHZNPINUm71tvmaxCKwtbwyfvh3ZFH11uzV2y
xPFsy7CXDdl20bP0QR/At2HGMPxne2rEQYLFI0ZLGS01KpLTtfmAUPzhqIXxTFcx
6WFeBD8futJ73BDme3qtwR+bfTUCTVy7naiWRSqNluHc3SRDnIsbyEVmL6z8usVQ
r9oDDvS6M47G0rqAN3Sxn5bRK13XEXRH2st/FzxsPZoaH51Nw/kGd6Z49mh3zYxl
tjWlB+gOz9DrqtcDNYEGv3JWTNxTDbWZdO2tpO5Y9Fntw26K3a1YHNfkdtpF6Em0
LvxEwpuTVwGALH1wrUgqyncSCkMMqMj60M2J8CEKEn5yPjVG6AigFa88RsrvsyS5
AXoF24Uxn1naCF2RdyOHlT0I57PqaCt6eeiXJWLhAuzkkjKnegI7Y5H564qWevtu
8YXUFYRnUaF4aQ/cR1uiQy+0X7HgLdUtPwwHxFT9PsXjPBPxrRMFF2/7bp/a0FUt
s5wel2FPBL/t+YBFyaq5WKj7+vhkI1WAVHwZijNnxBg2ln62P2CDW9oHNtWqQmA5
92zh7drM33QP6u2ChyzTbO2y8U6ha6ieES3L0eOK2EiCBC9tDsLINRtaVIx5QO03
9n/vAUaEcPzl9vNdHLFupko76kUWhKkIiGHNnSduiLfu8M0Ga/qAk2jsT+CceQUW
m/N5PnZyqR6qv+yjqIjHQUUv8MAZjSIOKkRKJWHILxabx5eF4h4l+HAFnvIFuaSb
Ewt21hfWlvqTq0h43Nb0ZAB+quMYCHFtWgxNyUXpwwleZ7Y1mslWgL0aAU67+T2x
D7i/Vulm9b9j2Ye6T2r/GjnaH7crw0vl2ayapKrJvlWDUgjjF+aD5aOso4PX3B/f
tQgeRiVCxJd5MjQk5dVrp3r+aNRBwRGGnVzUKpDwb4HBxuoWyghDXTHJR2tmXmGv
dMzMlDy5fPYMhX4Vyy1kA3zmCiyFD7V6XK20JIkIagHrH4bcryrvqCSB8ZrKYKn+
OGIayBrF0RxG5bldwUZuugry1RQ432uEoYj0LmYzp5ZokEE6WTFarH1vB91Xw6k/
SNIiU5r4AQ2yNYMlQrpFVKpeSACnu9exVstKozCBWJRepoWhPiupGwyMzxtIRPiy
xIHTbpvm7vg/4U08GzKbfeBJtPIRFkDEV9bKb6ETOFYDbbeoHnljiytpMHnpwo5S
nuZrXwllabXtgxuwJGQ9C5t4KOZDZ1R+MSgAyb/nA0JnMb3E/dEepmFmtrjOdGlF
ukaKy/Ouiebd0c13FwKeIRgIPtgs9nYfJqQmkFlq2wO5vn8sw2jts+XlO/hFQ4rv
46HaETXqs2e5FAu++GVI6HVc70u+YnV24PkQpBP6EXYbv73r2qZvHVsOOU7j2MkN
qkwLucZuJOqHNojP/XKFvLAfD8bYtKmhZFp43LA9lx4T9pISA+xWvUxNb93BDiDx
O5Zw0KemGuLfsHO/Te6lfj9oa+q/ngjtplBXrnag3qBof+A1FRXieAwIWbbqRhMk
dZdPFFF/aakLHMnxdKOXQsDf46ieqWyT1Zexlk5bxAfv6npaztizLAheaJS0EmKI
MZB0fUPnbXII8xoPxn6dBTXQCP5pLWJRw7ktmgHnnyp4OXSOrvXsfNauKlBD4Pha
2V8zCnLWFVpXMLCrcn/PuLZMapkPrnWrkyNIXj40HfkX+8sZRiz0iVxtqXz/TaA4
XcToHF5lGp+QyloA5VSibF5jBpKW2aeHqH4P3jKI7fVRoY20V906cr6fVnr3rgAu
AWsYBx3/N7pn5I3qnzbwXToRo+PqHt756wdxLWy6tHv5ZB48C/unpyrdJlnotp1J
r3ZZXgVH/SRMawdTclOyfPJadKVfPBu6uwbDyOS3s2McO5w3XbOmNm1pdlL+VR6F
k1kB6pYTeZCOwRWXlzNlrlo4KjLE0f0MynK94R1+oP2Q+okwKwZfotbjI+MxhxPB
LfJSSA++1aFgboefVkCAMC6l2PDtX6eNlWSgx7qudsjUN2xT9/uAIdpW9xSC+QYI
S4FnSUS7r8MJdzMY7Dgj3IS7c1TsvyTOf7OOS9dL/T/Ohm10lR000rlpxtYhrtaY
0qQPW9punQ875PhaMTOUQ5h2V/Rwam0m97jSsYsStg6kNLKO+PrX/CS92J9Tglik
Jpte8KFodrEgnp1LeXzms5gwHLec0aXqTqBwezU2dWRoAtN4yWpFk/Gm1eFgMSD7
+vYx+78RS+L6siferknQo1SZVJbuDnosDA79jMTm7pG/ZnmTdQ7SeKabCwpLbmqA
c4o+1KMcyVPQXaFEMA4eoR74LQXlBkG6ohqSkLpzyKwOT1WRMKHTS7AJvVlT9pL3
HLr7i7Z6JbOR8hHJN+VXiKoiVKeQSRUrzEuCHLeUGEMyioSfthjFVVqlLBExkekK
/cglN3AfmQRdDeqPCVNKvjAX8ABFz0ZGcYHY3241AXAT8v1ty+vl6DzwHGMLyZiw
FdFt1vELiUyKKbNraRBny/vvr1ExU3lU0u5l2a3Zw/6cxbnNxyNrigGAgngT4l3n
N5H4Or8+4+ef5IxDn2A+7vN6B87Y1Fvvo/HdUQhyvhgFg8TGsOFxlTzmul/6bkP2
uAEjpChQ64tjlrkfF/YE5Nh2dDYMNiAyATCe0MeckU2uG/bEugttkUjUrTQHk5bv
NuFs02rqRB1FTIJhIdUG56VJ9CZ4EXCOi5hocLYhh3xana2++dLEon5l+F5RW2BY
p74jguSk3se/0LRsD5OBxqBfbX67IRQnMTIW6iWyZbDw10iMPnWpmGvBDXLgr8Ny
Ew3BsXMad8WjgzIHg9onzRj2ZMsKE3uaDdaQzIRzezTkB4Uof3QRTK9mM/S5HBFT
wJrsKDg7tqecfeswJ2OQog05yhvywHMEOcy7tnlJde46s+AifNRPNHITH5ziPNQo
EgUL4I2dKYEUE7uMIUwBDGidNrL/PRiqDNiITcWy7pKKbc10VTjkl/4oxaKf3uDR
n1IhbjrE5/i83hDxHlKF5sLGEa/OcJy7mapmd2Zb323AtEF71CSINlReZKeXPgXU
XVv9nz35LgM6ZmNPob542SMmodXTuae6crFxTohRdCy8xWhUPJ7tBM3D7gWSp24x
rJd0EA/TVSCB1OwHEAYRQ+10ZYD+u+Rd3B13x0q02VBGIX9pa/iEXBY/c52H9Et5
S1pGTSi3pWZ1rSRtpW56HhjmEIj2T8HnJYeXtUd2n7+4YSCu/FSGlMFbMdysj0Id
iIerHM4NLFWvvlIwMyMt1wbJzJ0fJjrEqhQeRI6EVuRcyXTPMWaFfg259MmBaUIr
k2plZdNZVLSiiXyl8MKGqn3Zak9V7Eu6WV5uiVLs3DU/7bWX5AtPJV1fjCu4ZYA5
A7rShsZLVkMnLfcEq8bC/Xt+4zY0bPe+ALm/1VHmzf1qIe2ZIlOVlVFV7mAmJgU6
ILnlhfw/TE278AbJ/AJpJr7c9xv1Nkt8D6jSEf/F6WPj1AF/l8EKuHtIt8GVrxrl
nlyY6hMzMG0zI2/m59h6V1svz5M046r8ry0h+DIi+M0QBs30Oi+Jo1cSBiDyz4IJ
sRP9fwXXbuODbQLo8L8cbq8U62GkJ6wMMPFr+YgJ3AYTyEiPadvqiRBj0IiPmbJU
533br1haiqmNF7kY9ortDvcHVQPbQS+DJ5ohsdzK0hybqAwSq7MYjO6RP+dPGZjB
C/Uey15KvWAgQPdk+xLGTH1j9+c3NBv1INnVB83V/8dr5HcIz5+UmPB94Ohdm0vl
pDa5gYYeJdMvi9pZ7DEUWXrklzh18WtX2+Kdj9gMxotKppOAOHZuOo4CSsuvTl8A
tGS1AeIw1oZ3R7DYlb+tvUsT31rh8G/ovaphECLI+b/R3gMLV1IqBevSFcSelaF5
kBp2wtG8BjluScNJeEbMq/5WHAXEzCPcCWG5Z9yJ+0OG4B0LNpXfkMpojRCaFNmX
Z2rsRoa+kf+XrI+QSBr4RQAQvP31kZuO/VJcdxWUc4ChC1vpx0Qk6ro0W8C+IFLj
xZkG4gn8Ym9E9aILv/R4D8O5W5sPsHs5IDCGcoeyjPm5fS68qN5gaTTzuosziShr
ioUknSlsy0aLzviZj/zLJkhP/Ew8+mP3Af32QBuchXBrfVB+g+GaptwMcVYh9N5T
iiJQX15Ui0fQgtNoFE7SSHgBIssph1+vXXe7iUzo9p1Cob/fphFqnIAJ6xvzUZiY
QO6efAyS/nSqEGRhd+h9HkiT7xurmDnZEv99+S+CTygueKnMowAQhgwAetdjBXw3
v9OkNfzlQjEFlhBwdhvuzCz8nf8+BaSOLIY/nv+ydg8Hrb1wTi9rXg6CVZuhJT/K
QfjcGJrUQeQHgDZz9F+yyNRK5g3hy1Ww6TWnkaB4ToYj3f73pDERX6wxyBCSeDUe
zlV6/e5jC1h8ltiEwysxM6W/RVrnaLDT/WY5/HgHijfOu8x1E4+NfHNB4Gqrqoi3
5TYfrWv4PMtWK/G7cSd0CdCKn/RO4hYudaZMuyVGnSsrqu7qaHf9BITCJeRCeGZu
IbZHveujpTiiilqnERFJryNVOeFAQfhrkd42deGRLfBncoILSb3GDoXXfL2Xp1La
uAbKv8l8lJJqyuXFgY10Q5qpSV0EzlheCDKpKtcC58X7Tn3nMHNh2MCkiTuY0zJK
URO2HxgSe7g68PMK2wfAui6z+h6JEE+FPBmKMvhDHDlU//17WQ9JGnQJ7t2ym0pM
FMkFQOtI2u31/DpQm1+9ZGjI7v2xLD0DXjzYHQGNDoscrDeuKpCR7f1Q236vnx1B
yNSwQmBZsd3BJ36rTE3OPdFJTS3lxoZG5+zhYIBcbhEC2KxmX073T+WFdoc1/BkF
4Ta0amsvkQQ7yc3PQzMw6f+KcXXpfIotvP2bShWbEjwtP73dLEvamqgHHCjvDS/6
uUV05aRYHJQZ/walJXdPt1+kj63EdR0o+h0w1cbwH9A1vra6GBblrE2rlalsYAF7
tkDPKZr8JwdsvIBM2dr2rjtdrSJ0r888BNbkbXj5Q0vFD7gs0dGKB6u96rWvwcWb
3q48FvfumivLy0sBP3MtfKxKQ8O82e25AnYibFMV2SKBrB4/rcI1OjQl9m1/Gjzi
F4j7V8nYnIggjJT4Jit/zty3A9U4kkYPY2MSroRAzZe9oTH7MaNc+6tLiKyvaqfW
td4NKHyxuqRsUa8dLGLaDlfuvibdJifzI0rHw22rOOo9UR2BhOzccAuaUnYhv7es
81kENIHZUU3A/O+PgbgvPCtWKpVKrZslld7dmqcM9Xip5ddZgTPoxuHSWDWdgYVV
u3lIx/qH2U58Gs2YqITvo+aEtOkAfDqP9Hqd7h0SfdGQWYdqvDgR9ubGek62UcqH
C5YbAGfZmqab9eQ3oBHWa2fAjsamEQa1p1q+HisKqqbqTBxiFOauBCiQcwwnt+Q9
BZ0irR5XfU9X23WtlZvlj6dHM1k0XIEHpp2FnHwwc5Au98eZBEfBqnCDLttMy22B
KDxt4v8yp97i8FMN2q/TnmGREQUg5u/1pE+1IMJTXbGl4ULjb7/fhFHFzqUpeoHH
Lta2/K+0oZNQ8Q+oYR5AtTIQuGUrVZhatrKqoz/OE0I2Pjp1z7g/K8vl1gYaHRxx
wqdRyt+xaFMxUJ3wWTAqhfskica/6IGQYZFmU3+90+XAtkUoXp2OvWIxPwA6FUsn
blwhLvu8r0F201wZJxSuHBTWkMJq9loXYMVYemFe3XrUtz4yK/ELLQR78AZVp1sR
dY4E1zaR2evOcrcFbRsvJvuq0WoQKqN7N+4UXdAMHWJA5pcV3+NgSokwl4EjjUDJ
r5HZBKm1I3etKe78ZughbtVLY3YaPUqz5+0fY0Sk4IWremhJ2ZaOa0DDVtGG5o0v
m8Osa//YDsEldCeoqLTBAO0Qy/pvhfLEOql8o03J0Nz+b4s/7E77vmJ5aYHqV258
Gp9NYFhgAkM1MpHsIUnwq20qqRyfW/fBUxSAqHdnYgYECtPIAkUqN45fWFpPjgNp
87jPMePMqrwd5h2xIwNf93+NttTSIzAtRJjEl4IhZuxz10Wu5/SQ4Jh6kKS4hNWN
JW65DO0KOpiSIsAkDrjCayVG2utrmikskxA97TKoZdEdSDlulgN6jzZhD+MInK3l
o7WYf9Q00ZVtcGLIEuBRGO12r2ietws0gexavVkqgNtTegn+KXnO7X3ReTZ3ShNV
2qKKRdqP8uwN62jWzCZMgiw41x1HbvsLXnegQO84wne0OjLLdSJZ1yMXcyviQ86C
w+W6ZiZUuUGlpOVsMR/rUfzXsGNM1XT/V4Gp1o2p2JncAeCrUtYO5pACXK/Jomca
NHqjKFHf6EGJG4En8zmhTqNnYnacHSen6widaaOjexcfHjREmmQ6L5mSFzdIUeN9
PJW4VsYsdkkZy9kziK1ZDGAbIfI2q8JD3+cYI1M4xmAzfTCPGYDUcqugTyDJ/km3
deiPyk8ptuu79WODxjBO5ISAg+e6XUK+hrbZ/yoTr/9dQl224D/v07NCS+aQYZfV
znyut6JSYewqLQmvGaWuOEHJtT9/EHr9hjXDq2CuhwV4JdgdqtL/rT+QnibNql/W
r5GacLXPfgyjL0KHNLqZ2CfjpFwQAU7l0Fp7VlU5shKyz4BpzSt2zrDSnzJvOHhy
QkIExiGBXJMdkO8WhWdC11fobJYERQX2DqCbD0cdl6z7fJgg6fiswGkye2k5y0zN
JKPzbaYSJ+Jn2wrLFYHm76Ow/j8Mbuh0rm4P1B0ozV7PiSPrd2Vg56zc8psGCwnX
ObhhDHqwdfSxaH1lXirLIWuvE+yMVTRnwOZcm+hFlNRWmIOUi++j4H03SzFDDzPM
3RCFodPwOeHfZm5yoUWwNRgLQglPJJibYAhtsrhkrnf0SiEx4soZty1T+vm3iNo5
iPW7DvI/T3PlTBnTcBe1aanno1WldjfWuWryB63kp1jMse1I7v6neQT9rETV0cjD
46AFkVWf7a7O41t6Ne4HaMbe63Qe/HL0VD1VsX1oTQFi4B7vSsk4+ZDIWDGrymdV
qERBFopaM3wL7En1fU0FeYhPKKmxvqmrdl9iDs0Uzae9Bp1PDYCSycVIfgHdfhWE
QLCnsFM3PSxWvjGPso+bW93KAIVvvadEtwohBgv24VO3dJmX0FUdDNy0WdocDtjI
fV1a6rVshaTZqITIYsSNJdsPIDCBzVCbfF9sS/3bFomaqTCPpCXyT5qN81Frh1rj
Vpf9zYBFUYvdKQkzm8590R0+89z5Lz+ZFqOwJZA8hJVCglC0nzzHCY3LDoHZ1VL6
x5Xz6lnPlT3gQlx5Qf/rj0ieHnsKPH0boPX5I2Aa7P+/3m0U54edHi6F1Yp82iLQ
Nd+D1dfBewbRzFm9KOQgiXoVwUtprobQvMw+ruqgJrdqeLc9Vak57wPZsQH2CCyZ
I2U7SVdJvERi8ld6cgTZPWi7TgyslB3g1Lm5w5xLNXOr23TJEPfWYOG/JP87f9Oo
EpjwBjS+d1DTJl7tla5VWubrtRGZ/N7h+IMUWPIv7RufE0GqWxoDnsHFwIUq4E+l
yECp4sH9SBg5wCRozQeWpYZt/Y+UKvb1lET2sb369Xd7C7A3/jEohwBPhWskKj1J
LzA+5VQlPs77uJkpzwr28q95MUjtNalZoP3P3F303KgqCk8ouMambU4VvsQbOFKe
VYqmOp4aZtN89MKuQMJ6ykmzhCebyeNZZijqehEYgHmETteZlnwxJLOWnIc13bw9
MQFPVG1RYgqlfl3lMfaOGB+88dkUT8nK3t1X5CTMcxIvf07sH9eqZ1Iadvoq+Nuh
WoeQ5SbgChk65QyHcNsKIvnKJWu6m+FyQbijQCnvpD4bPe/VDTbLYPdpzDKmF/Iw
n9stXwq+N+8ZzrURj6QHr1121kMR+CkD3aE2vJvsJkxi1PR7fpuy+gSOpJjQh1ao
tLKeLVXXSVNhCzGZdXS3f/8K6NgDWO8BwpD5u09TcBbzN3w34sKowNwYLaTpgGuU
zXECi43iRIcvgorMfVvw1b/BccRKeHIijSANIN+A0IMDtNVE/YQbHd6GeeRbVGMk
rc1wVP/57hGswUHsBnDCL0X/+9QAhOQl1il4lH8s8wWudgaqfU/XPEBP8W6qKDdf
4oa9CH3vwWk2N2f5GL8DGzJhqNUalfaM1Ef801bUTcrfOOGJWu75it6QgPhu6Nio
spXhhdL5iBfz2Zxe5JDeqbA6rOPmyr7CwB0mCYW4bb9VW2wO+WYBKyVA17TSUpfM
mPXuFKoU2oKI0HwG1XM6efhTk82OoyStrwvZynFZBXS97YE2mljKRrg2DQsWmrHR
7ozB3+LJWZGJ6Ldp28Wweby7cwJL/0Q2fGmbChl5nNUrtHFII2CLrulATbDcpdBW
Z6PPRGGNYdl4vHwdKfU4iF1ssODkvTnl8qBJEu05cUiu8HnmGFKFNImQlx7HayfJ
aJ+jwXbAZKrp7TOSbFDisxlnUUJ4xVDAZ6Zm3Edt9BQIVepQcV8+TNDZ68pnwU2O
3uGUk02DvqgXl3d6q2wEfa6N3bnAYHfMGEW2UDdAdRtrRenDZsbRHSn+j/B9gSJ+
MZIIBjBeelX7KcmmzDyHXhcgOGrGsMCCR1IdgA5IgrJkBZh/RE13sL+2gkAzVSyI
cIWJHXi+mhIFn6VMgO8YoWapUAELLPvt30OODKm+tBCFgQv5L4Np8pPBIz0EW2U0
D49SeFpAlbNHnblqBEqjAsaFuBqPc7tAHYgnLAVsSjJmYEIbTk8BzrWHHgFZLe0K
uoTYeQ8saTaGDd8XhcaAiP7iLP29IkuYFELbzoFS5nUi40mj7WC0LDhdROakRd/h
8qrp88XUq4curLeRMiwTPW+qhWbpbjYxHhgo7tEqaBwL74gDcNpaIcwPMW0sTtUd
A5Rwa+kwQvKnSiJH8mL2orX1/a8ayV3JC+wOOXYVGKJefhFQorX1HwvJ3RcfpQgZ
348vU/9q8DjNLR7z9XXDXelsuRWBarvI3Rx8EB524uigJrDsvxMsmrK6fqxVGWgn
MKnR8PM5kaceiozQ6gn12qvWxDBpavuWyKfwBB+d1Uh5Ftca9RT/QrLp34mdM0J0
jIhzn69+tNxbCrv9hVOaoLsyVViJJ+OMUE3TvF4IfnMOyF5zG8CDNl+4Pkn6dYNW
/yxbii0/lmFjwGOgwqqoKn1atgcsRxEx/Q1Jtq0mVtgWt6cjGoJa+wNEMieSasF4
DbGxpbJZsy0S0brGeppMZMyBJRzlD6wWFb5cMWcJm6eVMSJjJR2SUSVItptWc6Zi
Qgc1oax/OaTErbBVUuEiAOVcxNWpPDCPE5jSLUBVvmEdSSlWQDB4UTELnpv8t+hS
SuST1aM5pA/KTt7mbpQzL0mc2sOA1xmN+IEHl3q+/mb0bCNketBiRWaiHNaqbnzg
LJo0BAPZ8w9IV7U2yjmioyc94GnY7CY+mIvRFnr48AQdTJZwuR7DR/sHrmlzzmUP
Lg2PH1QWstZHP1szrLkUPjo/SugQrGhc6Qmlz2nHuFhpV/EVvW1vkqEff0oIK70w
SO9kqcjKwJAB/g3NJFwACd0cUh7/fqZPB80SA1fFklfC0RQrdUiWjOMu3CMyIWog
tY7lCnnv7lhzDtUQ67UtQqkUGDE4pfXgaywxB9xIL5a9RLmyk4moLRpWPuwV0Kyz
dAYdbTP0jcQQLJlAG3bO7LOFMvagJEqlXXcUoYlKq+lo91Hl2EJDqYtYcq44Osxx
p/fRo+6d3YKB93cn8vWycowa6DFNzH+P3kuH3vAUC+GEDBziBDOlhNEpywkW5pa3
xyPSlrDuUNxJ6B2A2mIQ6M6WM7lJfdJe9qRyriIHyXs2t+znAUg5C6hpL/ayGfKm
JwCikKPzdyXR2gz9nCnAIvi5LOgWyO+s7sDNVua/ojtFcFM85spVpavAeyvTlhcY
XYz0M6mjYRK72TVwLnz3qxt/aQOQ9J+8kHLylItneRohSZZ3BykWTQqkgTQSnxag
R2bq06wtet4KaB6rc2EMZwl6vP43I+6pUvSOssy+RylulbfSMUHk1FwcFgGyg6eW
Oqn9Lpl/G/6KoqP4j2TDue5n+I+71iLwX2j5GQOgf3hiUfF6z1sPSXK78YuDFG75
xflAJMIEJ0QuJbYUWYxMABCXXgo025+hxyLr3B8mqkPSX4PG9kn6F2GBtRv95YAt
Lp7lelNm3rJMZ/NxIA1DHw11eCizTZYkI5Rl/P8cJW521NrLkTOxIAWfYNnrY7m5
uBYIqfdZZRmeY8Z4kqrqsgE623k3yYIcoKbvafwXSgeyNFhQYS0zUHYaQLQsySCu
VM4NatEiujOWuaAatbV/D/g6Vj98hDjWwfTqigfyb2D07xoAFD9ZYjilDvlFGilV
uM9r7G+Qmc9W5m3cWPVAMqE/4kBwtYzZ2BgtbLdvW6pwt0DouMgPqdEjY/P6WXwI
OfxxBDeRvQZaecR7jfqmmv6nq8sdLYF0VG/MLBVaVUr9DJH2xGIYyM2kZGN+JB+6
JuAHPy492/iz2vrxRDfeKu+POvTkshvIKN7MgsifKiu65hfJgjvqvIfF5zhzvxtJ
N2MQ95/fSU9ie+bGpKq+g6RLg/YVUS9zC4WFNawmRV9tprdfwg0GbSYbdjQuJ/3y
50W0A156AW/DbL0TW4QT9p5l/+5Ff1/Rz7p/vwetLiwJgIWoLNzic1b5i5DrQDum
wTelQkhmecB6MDUdxu+PJPegJ1LF9yAb8c45IHzYOElb4qAkdP6ji6+mh/BWC1DE
B4NqtI5W91UR2yA7VoJ0BbzU0y9jDuoX65qcQdiM79aX1evcYV3ED1WdPxMcYSar
1H3wNo1xl/OGX8+z9GqZvhC+TUseXNLwKZ30UcpCABfIMKL//Ywf72K4Fs+v1hk+
wkRJG379DJi6GVzzkqu+o7YoVFkiBkR257VfwAIVxLVrWqq1jssVCTaOiMquylQ9
KgK35Ke5ZCI/Zb5tVmzcxn6bCLQDm7CFYUf8/AquZeh3sA82zwUgpMWIba6Hopd0
6YFqmR6UlIjnhZYxzGb9FFDCUd8bgI+RqTI586hGwIx5+bCnQX0AT4ntIqBqpwcg
p/2Cf2W+gu9TpDyVn10U14xNvOxamHPerGOOsyhtnmNP7+07jaAd6fieasTI5D/2
8QzdoMhYXiX42J6tn0Au6o1BSCwYPmNydFvAuhCvOdIasjJcRX3ROtKBQyTY9FKM
HOrG4KU7+UIVM1HbLqCIcazfkGn+QuBIeC3hCfzukjXlRUDGi+ar7F8cOXrbuwha
j+bcaMtyY3f9BdTUD2Z9Cuv+BL0EkFvMuz1e+y1sk3qPbn4wDkAd3cQ7VSN5GyFL
4u8G2KpGtU65SnlF6SLiuX+PdVpbB0rOBG8OKaTHoF/ER/1g802AGD0N+5lde0o4
xLdVNDk8JuuT4t2veKt95/vITJqc/PiM30K5n/xzWBcmxndOtcphWHorYi52t9dX
/T6dSSYvfw6jmWLLW2FFUki/mZVj0JUtX+J1w7i91B42ClEqmDc6YUh9Z9t1k7cp
wid7fZKHgEHKYJwBcV9W8jhvp1q70mQX/KOqI/hd/UK9TgYCIFKcnVeijMSdX897
Rz6cPXNsjtMxQQuKvdAt3/MTpdNrfiiIqICjlcIG3Kd7lR/3PaI0HH6jZQxX5DsK
sm/+LFl+3eLdscVm0TRZCYred9cRZ8sL2Mw8bfmURglx5YM4gyv4gbevCJVqqGtm
klv1tE/zUtbk0jTiZEws5099UDH3wNSe8sioMbHtNJP3OScUcKNm9Ag7IF/Pyy8R
3+jSzABVDl+vUh035Te08Uhcu/4L9+aKCJjGPaACZG0TmA5KgHdVSR8URTeuuWwc
RVp2Tckxtt0xFQpCC1WRo/H9sT5QVomyTakGNVtvuyhMvdwiatHDCMq8MciNmtlY
SLpToLPlmz6ddAzB5wOg6LM1X6z4zNB0AaHQr18eejTMfJJgrMn21aFZQc4gG7xq
tD7abDbZG/Asw7WrvbgACZHGIIYWiyya6gu5Fi2fhvITToiUFaaRlXwpHkIXgP2E
crUgHLJSMCkyS15+9NgwJCVjb9pTwHSnj1t+uZ04bM4uFvND5Ue+OW/dAclc8Lly
lmgyzOk/cYejDL5An+qO1tL29ba+3ZDXlmzyhg75PEJx2S30ZdhOMDw2MX/F4mwk
Om2xHLLCJxrAifArMWl6devEoNV9ei/TdSzDk7gNTmSS41TzjZxcHf3MLHwM6ejf
nNmuGeX7bp29f3+3E/fH54CT7uW1+kvUgRRB7rHULlvPyQ8XBXzXeGWr0hOG2NGy
nzHPluwpoxINp4iT2E9Tbyccj/Xq1AiqKJfNYa0fJvF5F4PTlyPJjwDriTIosF3q
puQSZaiDRT4GvO+wnMpt3EvmxNzwE7/FMEdE/QLQ8JZuoz1JUFFqL1VwqXhRPCm5
905ff3NG7un4AhK6qkwjonXJoOR1uHpWQ8+QLhPLKZKK/506GOpyFMA4p5GsRNvz
pEtFGs/IS4qkQup34iUkTOtxa5DNZ14gf+/mb0FA6BbkrNe9HsgdwE/ogD7XEvmi
O0rCnheJpitGY6CpyZUantPjn0X7kc2F54iWtbvqWl8lxPPK7l0s6maqrUNHtlgv
hza+ANgMjIoSRJE7FcJvGfvp2ir4zhHWvWOEhqtrgTK2xySMC41lOSHCBW9TUvWW
9WhEO0o/QkeLQD9WTvpjVYHSPtF+h2uIQOfuRsLIrlf5AX9RN0yCmYW062rddyUM
T8BMJEAt5kRxoB7gRkAShzgaSUBL4ZHqBsze3+kHeyNqu38TCoVgF0cIvqT2La3J
UNbWyk9MG+h4hrdGcG8258iC8u4Sk0zCQqZY6Wee/nMcEPfMUTFzEyqD7QsxSCqO
YxAM8cHFr0ezipESmKpgGo8JJEdfs0upqsi2nTIN1yVEtaIlVC+ojoIn/7XR6qoG
LQ0NTvKXyfGf9kGuAelw2DxpTvJTAbbDelEGh4gqJ65iHLuReiSpQd7SURkQccu3
tW7yvADNo4hhLgzmmwy87/oha8L3NN6IMfRlPXFW2BaK3EghqFfGog/R33CoXZ+z
N4q5gJXjMJT5eAekhUSJCSuJz2XqtDmHEOn/Hh4N9+s93w2f3IJ2ZuOD+8LJj1HT
9w+0SMCfgbFKaeut27aqSzhw6vOKexYM8bT/m/yPnTcRGC8zw9+RHSTe2srQzQQ8
kEuGrSn3rL/ouG37zUU6ZJ+y8Uu+qwcPWpdvuygPdSiPr9bFwU7CrJJkNIDjOr9J
tEFQ/sIHoqLhO2VO0ptMASboYaDS4iCIO1bkee4zvagiFytaorLCxIGzzwiUqXpc
6+5d1g64a80ftUamRkisDBflcMGXymk72UqWwhXD+O3Rtqs1xn9w/V6x4y5vMfNN
vldFR+KUUiFgUdxlTmv/d2q4XVNH6G1V2KPgXmt06blIXPFh07+rUOrqlmXWMroz
icf+P08nsc+5LLOzwSUzvbuW/CKb3GxwjFpXQwBSN8WODMjYZ4h49Kv/4Q5fdu8U
rDoRo2sTbR1tziryu5X/Gsn7/H6PsKobFsz3oXXnDXFr89L7jkjcHDQXeFjO/L8e
ADBxmwV3ZeZetcs6wo/iEgXeee7RkU5urL5Kq5uIfxH9UNNnGv9voMFYKCFZ/wwZ
EdLpt1raFCi/Z2hxQVTKAv5+P9EjhC0HYscqFunrJCwUQW6xXpomJX8+CMoJKISV
8H47D1N9LGHzBNJ2p7vSdDh2KosWKIYTDWI9a/S8u2psQ0Pu4pScET9f8+ZsjbSY
/6TfVKngSK5ivAWZIFLFpCy5NYyOA8mRxR80LSQawr0TQ1JVjfIsj29yyBioNPqV
X1JbJt3eZQuIeooLJug0K6tExxClIoVV5HkVtaUJmFcAdSRixx2NAPfwdHmWw606
Oj53vxX35QLKwlWaJth51Pr8hk93hC2E8RpLZ+mL6Uszd9StBeI+cAexMtbwezyA
TxpMqJpTnfjOSlPTwaE8OU1ewUkniDrRWiirxsI0/o7r+Xs4GPP2HXZD+oFrq2E+
+C4ZzjVj8xp/UyAlWgwx3tIOE6R3Zt3vDprNSfpfsRJl/XP9j2RqI0M1FrT4o8Da
W8Qwp2tI06Gg7Khq9hMDrlWDckwOUkh9uXIEkaba2yaIEvJdV62QOAP4tXxowLlH
1LPKqcm5++YmTvjE3M2lNR9hYYNkVw5ACxzQ4JNQeLIKwrJvjGwyBp6p0i6KFjH6
Csy9PScSsuq6115UN1NiL8i8Wo6EzZ1Mj+6g9v21vVR1ON3SivJg4aQ0SdgaqPJS
JjcpH4W3Bm0MzfzI3iWDpNYBDSIOdSfMHNRWs6TwoG27JcqUTIZch+TR4U1qyOZk
FBNKnpkZfSmZorHiWhnacEm6ouU9h9SATs67Vwac79Ljs/ELqeKMVsjGu2eEHm3R
vT5GKa/OyqHcaW9ysQu0M0dsjzA5jSQq5TAyGboM08eklfklmrZ2tqFDuG1dI084
MumGcsIUXA5U3CeG9Ajnx0Vuu8sjInVUfocZS0n2WlNs6tW2RqWNoyOQqQ9lvdhk
ebcWt2XMskBFp0vUEoMR2EMbtZvGPSOqWlG7a3ng4AKiunIw1qFpnbTluuyUKs+S
Am9UJZBd8EFYLn4yvwlugPY32ggPiQ2N6S//TZInCeYT/+GTdtNrmpf7HkD3yrZ7
8tvKV85DZFgbPZVr3NCqw754/TcOGJq41QxUZ5vWaI5RoD2PLGiCu5rFIS6c9ZeC
7Y/1JYOxpIP9k8f8Ngxss6DZn0eo6KYH0++fQXd23k4c2JL0ElrUZ4W1Pzrk8IJE
4YSRkhvnXbmGnYo94/Xvlao7ru9fLPjbeiIH4lFpVhgm5uNhqgsF4I9xk0sgyEUG
HizjEGnOudOY0RYtZZ6zZAXJFfnrhbOEwIRIVdTawU1XofzV8ALSMdltYaWb6hsE
eWrsLDuRAWN5Nr7SNChQJyqP/dtV+6cxQkl8pLRASdGfnBCJ+W0dV/ddFZdl7G8o
G0GEFdIKUqiaOm7xGduU3Ebeji6Oi1iiwmUk1WcwL+bP31/nvjebd3BEsvztvsih
Ta8VGgvXx6dRlRTp8U9ZUzmTLjo+ukUq9w4qJDdgGkL3AyWTXACrWORuXL+rMKhg
UpHQyFQgLE0xYrTb2wUH2hsMxfsdOatHtb5A2alQVd4qhbeq87sZM5KvhPxHwH1B
rcUiMwu3ufTqHicbMS4CJjy/23UWKoRs+BiNa3gR25wVvB1EvbEbRm/icfRnKa7B
bGzY7rDtloSMYGCtEyOOnAQ6Ge0t9S8dhiPweiDWUQG4iztWXLLDOWhlQrKTi8FI
ZwZBlrJOouqQ50slDPqlG3QqgXS52PA0BWuyFKhwO7ZTHZeS2yfT9NCdSLJL6IDS
2zXjGIp2pcfaHdDFCJXapb/rq5uQDoZRchHphu0ZJzJ/tn8uEbQUQzN8wN0d/me4
0KeZf1aybe2aTM27yvwVc+oZMAQbOmHItTPELnJ0CDrWcpoKBmT3wDT0delShN0/
NUXvHLvuzi5MvtABT8LvymuyiPMr6xnEf+KCso0SQwl5Tp2j/4NjyPkt73YrblpD
NTx41T/9DNfGvj+sqvOY20OsohSKlY+hA6NRuN7dhdMk0RArMF6zxttmjeK0u6z0
TmWMQyVBFOtwvt1rOKe5uCHK/590rQEdqTPsFevrUGlxdbduRVlt1P+DHeXqwT7e
dX4pbLw65vpWXVQ/ttUp3PAfUnzCPjfLXOl6ZRTesLl2EiAuwj38S1hy0oV18bOB
3pFYG9hgPNNqFV47nPvDWlnTeK15rZLpUP6AXD1bRx+09MhEOVTopBsdEcbu8PRA
PAydz72LzHfu2AxSu3DdSG5SQPdKPzwyuYVWe+lZ8kJjvNIF7H0Qk8lwZaKTtR7V
NhQoHFrF0dHythY1EPJlB4Nn2FDFl49X8ayPorYTMsmjJ7GICq7+z3NzCmoLSrjM
nxbv/Qb+Lxy/Bf0nErAU+RYUc3fB72rvEnJaRh6tIiKsvHnc5UWkaAXwmk0IpKcd
fDaq4pIzuvGX53ZdmPw41RCvyayo86Tn34wInybAbFLZBugwQ0hGJihK27f2a9U/
HUKfZI8cdCKJQtQXj3Lm+uxYH8pAwovETYxFhtGE9OJMOOHTo7yhpTBtrqJ+TG0k
hdMAmSlRgeDJ+TdlRlwDMiqzCThKxZOvL+gXXsPvC31EKFJT3BdV/W/kaJ+3zAbk
+4DlDk8mbnvBZES7D+K0+KWFWzSsHPqxXcxzGbKWvtMDhsSp33NP8TacuL0Zoo2U
uWFCJ6l/sP/lajSvP16BoZ+gBmT9fgFd2zR/rtVpWH9YnHY0LloiiWdB1ESQMXhE
eediS2rVxUMvptApkyyQ/H8JgfQWAhaLVZ8wsu9CFzZuQp2dAaNPj45bGZXO6+fA
Dtto4Mipdf5rhPavRm2NE1Az7AZhRtIWzpJNVlrUthsTGmWT9ETtCQ3279DMcwN7
mrCCRFe6jNyxpMxbzei2OVP+Odtoax2v5RiaJVxag1q1f9kf/SaNfrIYOFvWmOn0
L+03wPpENDyw6CJGZ1k2HzMxAtTemrijpGZxl9PZ57cqbMLNs++YtwvhcdGzrLBT
a9qMp+NwpIv7XJeg2mMLgm8LmPCeQGtJHD9oY/VATgclwvrH8Gl/t3nC2LM5b/Cf
IQ9EWA3eytQc/bZVDT8hCx+S4WwaDX33R74S657eo1bc2aBg4bZKfBBooguolFTV
pn+2ls0wqssV0fbX1NuhZxYT2uPqkVD6coW7ElDxEjSx1q6fCVM4Mjo7QSzpaekV
IVysNxjh9uS39vtcwgPsGZA6NcZdawBVFp5hDkyptuZi4Dbn6A5LBM8j6nJkFOAj
RGUqOT05zzgyySYQemUNC/ehfESfBIYnXPw+Cb6GFeXnKutq3ZiDhl7BbaSZrQzG
pXcdayYB7U0dE48Re58JVT3dUDNuUc8j0TJqnWd/rx8DhIwooLEbsJhN3mDO1Dn3
CCmIRobhbAv4rWRTr/SbW8Sp21au1p7CA94xSmucHo3Wnul/znJOrERnODjQn0NA
Dwh7nypp6sAzbyBZqUDbTwhjLDNJkitVKYCIH7qRjEzj+FmRVRR3c0QF9MqSDVZw
tVGaGKjUH/BHDajGSJUz7Y7gDyJldKoA85933kPrbx6hNw3G1ftZ4Am3kmGf+JV0
PIMGAsYyeqRegtp/xha/j5Ci0RWCFoTTxAMWu6xdXUwp4ryZkW+dljlilHeN71/x
C3RVbLN8RqiY7A09qZj36n5PFIwelSG1xVDSEbRa4svLc6mGKH8MIrX18otlSJ0U
rP+hf/e4Q78HS2jSUmBaEy0IVpU+CKVFG5RT5eKG9lixgK74v/QCr+H+r2KcXYda
zwf14ABMjjyw0fuPcKd4NfjsFetqLSG3ymH3T2D0I4uyU2DCDE9fOZeGP1L0GmNK
UnUbZ/2jigquBUsswh3dtLgHQTpdSrVa1BkzOcTvfNoerKHK5S6pzefV8BELJ9hK
S5otehZ10YGFiiRphBWd4Kd73Gb/VcKEBug3dyiPAb4z4v5XfyBKqgT0eTHfnTPU
1WtRwkuI1RqHs/MY1/Rfr400yvU3EkdMFqBrbLwu3fgdZ+YnU5dPNITpqc1yWLA3
/BBKVlSuLFDRFJsm8XbvGV2VSFxIh16Sd/e2g4BMCW77j7jM6RBNvIStqz6HIg+X
sBPSJr4L5qTXg/C3Dni8ci5d8khbt5hlwuyCCoOd+0s1bt0/jz3+qq4JiGq5hE+S
kYML3rJWNIue9613U9jMkrHvazXNnLYZqc0FoQydh2ga5uDcqUWg9XrpzSmbeC6/
t9SHZj0BT3FbsKqashIXf1dBS32jwbAlId87Rcl2cc8UCEowcz4loxGi+XbLiFWT
Tap7i6WvldzBmMqjOQA/6mrHapG4xSNTvLBY2fULjsp5WUWMbG/31ZjG8VSgdF/p
jire6qjlcPWkP17QaO3eDFxz76guKdQwLS0qQR3V6nnG9sHmyYm4dpzOwWxdCKr3
2ISI2SsvLvyCJe5ZquQXpeEcS3zZAVjLcMithWpo2SNLW9k2IspE0xs3GGJ8xmv1
gqKzZB9sjmDjvdsUT9EkkB8vJR7+yWqJgp/R+i69Wf5aMxr/0dbm4R37EtsqeOqT
Sk0FLx4VroqDmMK4OdvzW7JnLWqpx17A4N8Q9C1idqCvcuGpKXZnCiLxsYSOGprb
xGGTc21Vvdqc5kBmFMS+6a2lGat2nE2QTsenoGF9DF4EA/VKFKra3vLcXZyRnGdR
aVLwJAWWcpIWtAR1zc+BJgY0DenJEkJK0Q1qWs4kBZYX9BI9zIcM/HwEN3IAVp+G
IQWrwWZ+z71wpRzBGU4NvFdLNjt8nyjtsYkG3XVI+hai1eT6EzWlWpnlOJn7JTYh
2Qi+0bmLPWf/1vqDsevJyhKiyru7jF1Vdp+lgEfYT1s4Q+sAsEdMYnjjmNHyu0xC
y96kx9pi1A3hhSBLw+iDVHF9dc7xBNgDMnQQfY8KeVnAQpNBfL/Yh09NW4uOdwOJ
rj3g1h7tfWHcUZ/ujz0OCTf0ilGN5sem2c2gx3ZkwPHhlObyimPktXM3lC92OjuJ
M06ZgbzooRifsZ+qU/EGcKdLTXXLTurPvJ0Sigyl9XTTNNmG3QvgqQ2ClV/H7arT
kVhB+VfEmn3scMKxfWydt7A+5JFH4Jk8SFxzRZxglh40RnLmnelDnIF1mUluTEPp
v0xY56Z7gjjyEqbnDrCKWY+CJiMUHwt1LLKlWoviFRVZC606fnlBQwOnLa9kAJL1
25pWJVRGzmyLQCi3DYaARw1tUKwUoELZZwzTAUWzPR6l30B0PLtnPusAK6WMZRsu
VbfSMDv4XxzuNV+lnkOoHGqWoemqa0r5wPkUS9NuBK0uAytvvw7LFaO1zT10ZhYA
dFl+pmFojQ7eesfl9r3SGHjVebdXs8kXUj/TAUTI9uF5fzBrXgjhXO4AAeAL2p7J
dY4XcyjfBgFyzCpAH3DRVvQIV3F8MzLvDyMrxZ3KsFn0nRGLUkROdIgGgfPY8uIQ
nioo57tsEVbnW83jY1sO4icA1KbK6hMMFZ6aWzqBmOBEoM9zKu+qd3BqVood5Ord
DXgod5YTnYbKXzY8BygWYXP+LHVH2anRmvr3pa5Np2QZmH0GhkAJUk5lPXU4jAut
NtQGKo4SdHNg2xD8V4Wz7NM3ow0qThewWICOuz9Fq1B4a1rr1nr+5VKKgmiA3AQT
nv+DPHInGyS1+rR+LXS1fv6XBZaLc+vzfyv414oNfQoy7iFTXkESfSjFo6vNtVMj
N8mqlX+bJNtCjV8DpqogiqvHJIjk5xw6usV+L6JjPQfLDq+esL90tMbuj51FaoAp
R+DLeolxr3aEW0f9+N2nZ+eAloRNoxJFtx7oJ0WqH+sI9JxLuxZ1cVB7KbCvlWmq
VTUVu9idcDnrCfAPe6ykO8kC1nDd99mrKPlGfY6hcRfbDs0T1aJlRxjYbn4LoQqD
SId3/PZ8sckClVAReyvxTFczj2BisvxL0wfubdmk8lEeeGZU7AferVo08kRyv6cV
1ta0M+8YiQLMuCswfzOxpIsjXunc70ChOwDU5yeTUwW6tb4GQtfpcna9EzOVzNUy
HAyY4KajyxlBxLvTMrlMUgei1tH45R83MRvroBCfYQL0MX1uhh4IFNju/hcZqP5o
pOfNoGn+eGuu37mkMJN+TgRZxy76RexmrvVzbY02YrA6mywX2D5eJhA7Pj07/Owv
303tMeHh9l+1/c1tq9NlW5co8PHoPTFP1NowVE0AoITK5pbetC9lIzsi1apLhvG8
9/jTs68lT/y70Kq/HqVa6FCAFBLith9TTAZV6fSlNlAz1p6tR3ptCu+UKciUCDhL
o1D/GgC1EKzAw3ZrPot9Op+z90AzOuLi4Hqm19KBcUv3FwZoDC2PcqCqKXanCBtp
onZREm7wgX78SePl3zUIcyy6biGkzAAi68mpdd++b+wX2UnhYFzRxoKZgmYSPoiX
bzHTVc2G9wjm+GVlIiINYDnBw+F6GHZSTcKMJWdp3nrpDXVQPxlEG00GZUdmBwfA
yrXMSdJEaqFavl4hkjY08CNfglMH750VQACqOORoEXiZvB9xUhGNQhv6sDaT1tMT
j6L/Tme5kVjxz1jx0g6FNEkfkyzhxeXZIUeAOGGF3hXEGokwcqUp3lsTahI5D6/l
S/5MacYHkwmSBTNAXjvBJguRZ6Iu73kxge/Sigpkmi5KBaLtSE6akfAPmOFhaJQf
GCfRnpZFl89fF1FqMCfsx7cowA5kKslZ5je81KNPxFLfKFxEkuFczovqRa1MGfVR
g3/FWJaFCE2mZTdxBdFYz9z4srXkpdp7xty6sKLPsK9duLYDEI6UbLo2H35B027H
kMradwR/0fBdt6yrwIsm0b/kCfzfwPjMsMHubYTCX0tavLU96zdRJrrPcRPtfK65
uYTiFkFsuR2i23bDhzba+wSqD7PsosdxnKCXLFeiSjw22dJgQLKQSXbx2zA9tZZc
mbGf2lPN09SMjHHVWOBCZ0fqChWXLoO2i5MW2Dj3hENd9AjeJcxDNm9U0p1THUlK
CIdQcFPZ6rtHXo6UqOAGKtbAlejIuBFWxuT5b6kAQ8qwyqIIuI6SFtitzMWJpD9F
plM4E1qe80t8I+tpjXhO/8GTXrBsGkwydeHkYUgAaiNMVxfsqv8CeX5SYHbDx8si
MzsrD3Kdb2x7A67pohSZ8w3IqGF281ptwAp/ZCmi9CtbsDtycOIs/9tpQMPpM6Qx
nX6uR6Gl8FLb2FZR5MdcCxJKTqF/3ZjRTdixB8rdNjJpzC1cOEFoOD0jcjCnUf01
dQM/n4/RhG6qKYnIKvXW7w5YVEU9WpTcPCL3kTFIKjQjbxoDWKaxeh7D+HvRcjA6
wjvcr/Puh7qD9zqHIgJkPdrgq2RUMaGXZjwFrKuWElbnQDyKzhn1er+gNgAweIa4
bVyYtlu7UJ4mZz/lzbqWXe+xd3AxMPqU9uyo2x8IpGNVA+GWVcoqvIhoX5QsbrQi
r1EPJxOXD66Uh4jqzsIa8/CxzM1Fq1n6nZ3fATKqQEeajkDJZxMMtBbaHBvgWkwq
2lT8PbsT0uFsBjZC5OaNEu1xzZvwHvVHAgVl+Eqv4kGCWJLxp0Y8xDsWm3FlKbU8
5zhHADFF3EV67Rsm4yi/RKUWKXex5DYHNr2iI393KMaV+4k0vchIaGlOWJ4qyw+r
/TxpMzTyKaze4tzDhLl8FsjLvd0djT0e5v3jkl3yNNaqJZCRABnkoLbkS19oMsS7
K601x4Jxn5pM2n7axwKWk9XDyU54WXSN5rCYSTSE2z4Rf8CqtsiaW2pVSfkDulsy
8MQ3vxp+z0jwp/8Zp83d/WUQ44YpppKYP2Tfya+YbNopp+1kLGWPF5AKKbokjdJW
01Oe5uHfHu9KaxNRbZJfMWSOkX+80bOE7lLZcSSfV8WSLw/pu4Et5Pzfzyxjcrwq
utAUWvtJB7VUWliGO7j6IOnVskDptktXyR2poLrmz26v4Wk10kLOPEG8bo+0VWs5
7UmI84G0EFAB+MQDvEsrLwGJ0g0LSydwLS5ntxzYAVPWmj8syuA46qCJ9n8u2X1M
kq0Ub0vqWFCNluX82iM7vjxi2XcMw8faJVzDz9hWJ/UksM7vsJDg7j48q4stT9oE
DcQkbw603rGKXuqQdLqn/heqMdJQpcTvKCcpJK/rc+VoagX5os6P9nL+7Lyu9Eq+
Uh7sshjJ1nJPVrhYuBmevnODgYaLSm8rpbxxaijQ6DEzJyMA0Ska2+Y1ol+OESyt
edcz2M3P6nDjUKCn8sYotpQajVwqjgh93MuqhtUY4Jp4LbWPTq63zXTWFvDSJpzb
4WzsdJMiQEI7W27Y+wES9YLEFhSEM8d1T0wQ4wp4r+G/VAyQ75saEA4LA8uCV21x
Lx+blINunZWHrcciS0eYUWrDfS+KdDL+yvxA9yGNaG+9O5wBOVm0bn83ka4y+v1E
q65igon9enriLQtcjtjvhNE4LoQKZQ02EvFoP6daOy4ZBtSH9GvIEy07UEFKsbJm
JfJ6lzqq026ccvN2aeCmKwm1J4lpILR1nNw52hAyQLBhgt2zJutsBrjAYhPvc0CU
gb1IfzRwhbijGapAN+nQPeUhAEmcUv8nS4pfHxO+yNIF0vsVCnfjrvTpfAXyBdVz
dnvx2OoWJJx1BnaWi2Z1qONav20bn4p0WE7hoLyyyhBIbQzLYOwd4H56scxek27Z
qMq1iji+xtgK6c13uA7PEjoPrigy759cJqdfhU0VbcWpRt+eRAbGfm9W3BB804wv
Mp9FcKy5f9dYDml4PesFP5ctAJW7pU5wqUBTDvM7L76rlXCcaF0sXOPj+GbDdMXd
AnENkpVPKhLipWhKt3LFvpuReDP7CbYj4LKLsW445JmQs2dNpk/w5oKCxx6nDhxJ
HVKQ24JwaJX/0rQtUZCZqq6uvLzKVLAxaICoTFFqn+St/II7TAG5uqJYS13UlRnx
K0UPQou06b45PIKkdLEIgMc/kFq+kpkPu8wGlOXwYaAWNe5gqcnIH63Zg/btctHZ
yJXGnYcBj1W4Re4tug6tTmgLelubbq5TLQbD7koA56V63fe3W+4xoQIyzEPsG8Wh
Yvo8ugK73Xsq8S+mJ54ECOATsOLoQg8lWCgRkZ4rISlzkquln7eEzx46oZ/LnY1V
MV5xBiNzTgTQWF5ZX24ppOfk0mdKsmYyHpp9FW1HxZkrT/0cToA6QxMl8kr5k/Tn
+l6l9w0gDJJlqTnnDfsmVsqpF/OULsvxHMWQuULx/+YJqodOyVxNdmU46AmZBlD/
ICTUzx/cAdWWW05jGKsHQPQgvbcdquToLNWZew3SU+0zc5EmkdLEI923XjQYkeNx
6rf2mSQeDb9zP9dVP5uykQRffBOWOhFiaCm97aDcltCwOhZdehl8fkWGxjK2hDa/
55hhEoTUwZ044hPm6QNfgcKH90GKZWbzDxDX2n1IR4t7YXPW1hF1vJNDbusX3d6F
XXpbCP04YnLBEcCed6DARjNB0BmSvS/dpKJsEMi4JZHUceBkwxNhPWb3e6HCLW+F
cuopr7z28o1EgMenQuYXHxrplYEQ1miG9LjY7ViB9DibYtbtA82LK0eXGYQfyx/8
uow9YLhIIx6b9oD+IWay95GOK2WAZTZ+CZ6nZDrTyodsey7K0PLD9AwGV4j6XjW1
01UFEAImpcr3Gs6Rpht3MrKEdIhQo37JYajmaUa32cpvqwiGpyTRxlo9FFk+L5L5
Wv/8YhxaDPeP7ZhM5okWWp5GzgqKBZ/k9+pbiN54bJj5UrtGinCogeEyD8gS3NbX
6bpHPTbaA5EaDUDDS1aRkMY/vF5KwyE+2VcrbHYcFLLhwJOUfWv8F8TxbkFOTTS4
Eif/XRYnUzZ+OCV+cbKHRFf9naQVhwKm4lVpS21F8Krn2i+Y1W1jhkuq40wY1Nvv
Y1vHLAMRS6q2mvgI1F7LoJAYcsyjIUYemBjCNtXhRDQkCWQYLP+SKsusQ2grh+7b
npH3jxCmbjgvATxNUSE3NaOCrqOT5j14yBTZt1HMickVqbtjQVWKsJBMkg01HSt3
mUi1z2D3yKsIw3TNCE0lCBKRndTj5l2XLeYEHmgv6798gZThTSFILGdl/u/9KoXK
HoSrE2LDIhbJXGMWkeEjzCOoWy8pOUHPsOng5rUiZT8n1MRGxR5JTYNYzkH4Picd
KZFCvYRe/a5xTfe9eZFdTs5rCU95gY/BrwnuI703NnJirGDZXEjGp15BJK7J9cw2
V0ssFb6J7d/GDu1HmDv4KCTmB5FCE0X6NrByWk5iA5cmeHNUITY9PzPiCq/VCwtW
YLN/pG52GszAq2whkYefm43cWLXJKckckJqlOqgVBRgHJnhOyXbcCrNI7FS8YBuB
cljJGiumcLLKf9fDQcqi31hNHUGjEEfH1X0d6knnK9BSS3Roc6QswmsLLDilbVzx
UC3wVsQ3YsMvpR50xcBil69RMdA+QdH92e46AKb17/X7vikwY/eUT+dsVz/8XKE4
nbIpVZff552kbUsFblBK3Gs6uaSiZqkthnnpBPnUcWyplMhY0BHvUMAN2n+0vugy
Us3LyPYAvmYpJbcurRPA0Ho0mOrqubSrt0i4yZ23Jd98mwdT+I5Go6R5nWP0ws6B
paNkg1KEajQsW2b3F7MgKDonfucJ/m5PiCqsSlsjVRIxgoOImJUVGh1Q0+ym53UA
WroFFngm/Ixp1H6NxBROrv3KRE3gum02Wa1VIryMBJGYYG/jE+XkHTYuksdhMZTL
jEzcsN221xXP5r9CD6RprLK8gHh062nZOPMA0dYK0a4kddOZ6O5XHmBpnsg95KSG
TNRu3AOBJ/fuRSwLkzf9DjKZBMCQhuoclVuQQk7PQAlN2/V4Ba972OPII3B+lUja
7CQr2YlNjijaryLIdxQDMogwshFBeZDaWV4xhAUe3KJEbR7XHtDCXWkLwDbDD9+t
TVTAFCXgOwxXbObwMYHnMNROGOHKdMOkpv8bqKBvEabvtP5m2c39YeIZTlEmNo2W
rUdS4kHRfEBdZ1y4NobLTQIc6wqtiKkLKzFcaIdFR7qblRy3TapP68ciZf6hrqWS
p+QZ+NaqT+fGuKfRL8VUeX8exL9Z3bHuUBqCMNLZaq3zsTz+OrUy5LwJFI3L6fud
QQBNlvlbXOPo/FwuKtDQh/v0OgElWzvGk7VU02SQ0ULAUfOoDh/01+Dkhth9yvjt
yCS7gR35crEGiU55GztJVtvV4+GDiFQcIV/Nf/2Q62Epg6H8HqUB3+ZHljW3R8F0
bNCINVCqmiVydTgjbj9QvK3kGpexpIKRsFCDsVzIq6lbqGPKlZc2noW+u7CUCirm
joocTDKE3DACHFnrTL3GtmjpxeDR68NnMVdv/9+lZA/o78Q/GXVzC2u73SkrVbbE
DwlyHv0lNPLFrMOAPysUg9lAVk6sebKCFl8L/akHLfC9cZt7V14TIo0zIUHejSSj
fGEDgLI7A6OdqkBLupdq0wVQbv5gsLez/oFVMQn0KU1VwdOo80xOq1RFkw3wahyL
qhDA9ekbEPzAsdmMtfoDVVH5L9PGrOkxMkN/VSmSPgX8jC0qkMqPlih4b/f2qL/6
qcHgXsBrsOFIHmENqQTOedxW2lYF/R8o/ofv5QY5LimR1yyMk44YvRA94p24vWOW
2LiFpjDd5ehbfDPQ0SJNFWN//nZZsYHbBxZq3wsUad3D3DLLWvoxC8IwwsDWKDoV
5vI5VhRptUZMrg7PuJafKrPO4v7e1mgptvBQQOttVIj1+CrKdD8Zz/mEcoimfzSZ
oDEpdFrl/M48rK5N7/m+JJcq5jfCuTKkv+zclRallXj9Pn8IAlQFInMB2Egn1/4G
MofMPms2gTcNO07UBb2WySLK6jXwmapcm0YHyeS8l3egGB6L0isVM9adg2g3hAhn
N0RMfnpNJaw1t8w6cle2fHHlnkfQRn8bxmFiQUs1Ivi7oQjRYXodO8shXsexHBy8
ep+emot7xpUWBw3TY7jShHMYynjG3SK0AIcQ5RIy6FdWtERBe24d/DfC71asGtY2
X3I7zQQ63IDYU/FN4WsyQcWFfjdqVKV6v2rXnZkT5EKImzEeoysgnUiaviSO+J1X
ztwdX6GVYyabtrhvhkqnY1XFXgkE7wdY8tv5TMYZ2eep2lgHoi4saGvEgkUnR0rg
yPg7zQuco7vIkJ6K5JmjSFQXFtLZHfMkQG/Er0UwHaQR31k2L0cbrW+GwS4bwnNz
W2sKgZuewU2Z3v59iVDK2v6jLEYWF+nFWIKy/t6Kq+pDSE5ZQRA1eEs0pdS1IBnk
LxPD+kFqQti7a3yJTB2szLmfoI40WazRyrstRP02cF4wGTxZgZP/DJAL6m1cje4N
daGRk9uOZgyEoFspO9uSdb48N7I+vA4bA6e7tCeWrGc4N+oahvYxjv8VaDOEgll1
FO6xQ1Au9bgjR24UpjM4skyVOKz1vP1I3p8jow3XvQ83gk4U7/jGZ8Bk3nrphYb/
aoOpctToxJs56F9DfGWQvJKnO3Zm3DHLFd7SxHdUD8joWNqDdWhd43TzkhLRopcE
ngAC3+OYwg2qD5NDP31MCDStIJtuUKOluw6Jrvro9cYFXshPppIXjmBN8mPNxJ8q
6O2Cv9WXe0rppxZN1GGfuYv/zYziCsyVGhffOVEWOTRoF4p/SyYUMiuLCFfzJQrj
9lvQjaxf8ODO6Ttj/Jz2zuv8KCSxV/zizeBL2+Tr1WgnG1KStmhp9Zsw3EM644U/
bBW6rb8XQ1hMihNqFCogfWegPfxw9sgcmkGOUwkBYOTuKK58xbrFBJgMsdJIdH9i
Ge5PCkMrBYqCYIk98T3bwbFjtlvEdm3KcyHTpGsNKcLBsWQ3MRIjac+h90VszRJZ
YbFNzigXSq6QWhm/Zm67t+rCQaGtWgmzOciLq35YcECjqe4C41R23d/6Gbh04tqQ
093b0Grq7d3pul4tNkCVAzEEOnYVHOZRPvwk5tkW9RgBlDR7jmPMqbdzdvmwUhIX
f7S8YEOCN3bhw58b4UTDjyRfW2/HaJGGGXpUJYbYpyeXMDcl124iHGZ28gHOS2wf
HrVJduO2jqQ3sQCazcNmEKKzjACFMduHyAheCsNIIqG5giv4BHpq1tE0NoH7Gzs2
BS875zE/psm/M3vtdxqLI/1ri0j+bENjfIuzBJek40KmPlqXAlhnVIn8PL47Jl+b
0m+j9mJEvx7vS/1uEellU68t6N3gYTeZ+gQpXSWUyJTtOKCUJkGiuL9DgkC5pXoK
abA2AjeICu0gM4rNF9EF1BE/hP1XQIL4kU1gsDpGbBeh6cBMq/p7z9ElERzCqKm6
Ol2/tkk/HTxheQJiTGRUyCUmIEt4abNQ8Pus9+2nSB/pbDLJtVa3N6x1tK72IF0E
1g56DyLgddqoDMg9dLBjiJSYJ1jpvjiPJyUWp6VvDJ4Gl08OzbotyIP2zRoHOz9o
6gsLS2nLucK0916PSV/aU903pO7kCFuJO4D+5zfZyJqGAiNQxpeR538bac4nCpCg
tJZNBOlsqgONGHvI5Bg+OEpi7SNlxmGoTrjNS8eSFZSTx1vIxyq4j24GH4xZe+RB
Q9kjh4G927vp6DbEH8LnpB11jqRJYd/AlvVcRAskxHRVZ4UIlp5KNQgAYKkwtTX0
hWSUOtpoFKX3NMK9D/FJIyu+m2QGg/lk6vqBsg4HZZ3XutLcR4emWZ1hHY43M69k
6IhY89gJ1n7s+/1Bfo5X0QYtDax+NnOnuJc12gz5bKSXEdQgDFeTHq/4e1tGUvPD
59zA9wOKTaNREnvaDRnlypu3Apoz0IJrU72x9mgmVXmQKoqDiA7+FLCKodnj0lMH
Dsfzwy0pa4hMB03QiJFWMSRvB7VxDJY/3x2g/O3DPq5oADOF8kfy9DFfu1DUfdx6
vqOmtsm+UG5GffpiHgn/kkIJnOlsj0XnsnescvjtHF2elP58mZi1B6XHTMKDqi4x
CWq2SiWr35PQf6lCm3IM0Ynw1yCWiPl1lCfGJaaCS9eAOC/6tmp9M6eEvR7mx0zJ
G1m8R7bCmfSnW2H66thT+0tQf5FpIjGMBT6OMNwv0fktPQNNtK43wt68flE15/Vp
qPB80zzkBlw+F4Dn7+9LpiIQM8Vc6LIur2Cs1UuwEwqVC9pPaCD0IFvppnxXZbDQ
fLa8qV7Mlzjb6PiMF0wZrOwkF/L9nVoLjXqihw+xzilhhoR4bEjNQI9Wf8NlrMLy
I++reZiEpjeVrKVah26hM9ljsUW6aXf7UGKkdBeOvBQghRsDUF6npnLzkTFk5vQf
30ukWt6ibzbtL/+GdUyf+ey1bF2VgNJgWkSTSsnr4I3aDLhZ7yrdR2UWI16jNM9X
qGDjsflBBPFwYAZQIEOAMTBKMlsuRtUczcr5Wf6B0ME+g6+WyhHAer+AMbkyTsMK
eWavxS0BybBOdozF1FwEbabyWOfxjMUpbxGfbcN9pl/5UIzoIbMjSAbC2u45g4G3
OpCC1cMSZzZAlrDwCKtDhqbQUGJivluxVya1YiixUizuqiJl34v4psxaIf56vNGU
YLmaDjTdyrnx/KU74gX1XJC8Xlz9rpnMfKoJhyk+xGfduXGWLgu7LKkaGcSrShz5
9av3GQt48i4vnNPh0S7Ig+aq2j3+XdP6ovp2zRI7yRFY1ofK8b4x6SxVPnLP8p9Z
knJSy6fILDnGNqmcyK7p//uZEFWxoJSMIqfvcfMBhB9byoQGfg6feXq0xAuK8OyI
WGLDXc9QgA3OooaSqDaZ6bt69Ec6TGDF6wWGUNnDjFyZ7v/WAODkLAuBapdH38u0
RSamYJTFl9+xMciLxONZBfTjnFQM8eUSXhlmJAuLB2mOpGqRRAkZ+gEfBdE7nR5v
8j/vlZ7dFbzKRUMRrST/qTu/SRALucsgOyLJf7bsv/QQcKdyylfdJKX8q8EvuJ47
/9Iub4RMXpKRVfbh7MB2iQs/dGcohGyJemBwBYuB62afAxKkWJXGkMEZ0wV7gSbk
7c8PeorgSqppH4Y3t0vLQ0ldfFQHnzyhQq3iASoVRpb1LLNVtDHrqLuoeYl6LbsO
5o+o1w1icIpBO9GuCKi30lP4e3bSvUhbQwXSBZL5PSoG7DSGdHZp2MrtHRhexFFG
Yel3on9QK5hm4ndp2skTUpImd3vnpql/4UfDFoyliQWnzAhoPAZJvaYnVEODHXqm
K0/ITxoY8cEjOD0CaNPMJUtdAsMS4Q8OfZ7jX1Cg+2jbzdd+mC8xVMXOhEEE4NSu
ipmnlWHKauhW6aU6P+M0w2XsVHNMd1M6Og9QE0T3ZSIONPSUJAyoN3mrQNnm1RxC
azwv73Fvhzi+/BvDh733Jbtr5CGssnOhFyXipFMrQmtJWGOzXytxoPRLgy1n+JDu
xcfblsAlWXm3/dKFmVbsNz8ZWlam9WW0kWYjldvFu4P3eC+jCHjmlUaiexK+lrWR
5idPm8VhvDCAGuw6AmV6YiHCykUR5Q6GHYeStc8RLeLeayKKl80cC1xiTbPw3N0w
LKagCEtawUbRF34f/Ks87qG1YeDSryz3dq+DeRrRSpgm3HHBXcLMkI/n3tKA5XPQ
qMwlrzCD8Al9QCslO0fOMALnjPvkOxioSYLBt0w64z0PcNB9z1vXvuk8M3Z7UHyC
wgvNxpaPdPjjSDWgeYxRO598C+6CF8048NE5jmyByk3hbrRakz2WdSxuEstwzlD2
JUMFCtay9u7x2iHminWX8OIJ38t5rwXMaKENwBcRaGWxLAWslY7dCqvv8FnuFniM
tZeCO4OwQQ6ZUyWPzkQntgrtlfgaqQOW7VejmmPkfl4hB5D7CqTN8D9c1BoIY1dm
YXfQ9ctzEnSG5IHUcdyeil9/LrhhbFbU5NzSQxE+jUXvY31hIpaGOof5D58hJlKB
MSX4BrdUy4YedV+GEGFW+ly7ZxSRTn/YpzUmcsbaCbkip68mPgDlPbVkBCuiSI6O
3g/IsYG4YvFwqxgyt6BocELw1kR+23OU5txbMAKeilaSZK/s7nN0DOxlmEaHYb0P
jj0xvM+HvQhcK+56KzJ1MEyEmOhjih2RGsrdRzGMt/W8svRjrVffIipl1sVFTIc/
RR3BLX9ANOlrkD1NhJiimrAzx5REgCFNesrM1IxmgTgyL7XkB4c5HpAUvJU6ly4n
3mkd7uMUbdL4PRecZkO54y4vFZKZgzDLv6KHFdMiU0ZXw7Gi7Zi3ci9YVbDJApYC
pLCBZIKQvLS/Ow31vncLK82a1oL2FGUZgRQvBhd6wSEVm33nRN0yt1lyXIXmh31L
uk1c0aRW6xT1O4fdAkONWmRdgZ7QKMOgeCJqqKCcEwAw+MRbi44xUQJy66wk0t1f
HPyPDksUnsIAqWD+5un5CZt9WQQ07crVXgmIfZC+mENF9gAVdFDkedDKF6HObq/3
eqhWvLRs8zatOxg2/TxyB8zONWe/vEmHPq1ttQD2kQGGp5TdO5CY5piJ17z37Dzb
5tfPQRX/2Y0XCTJpkQXoWj8FBIndTTokihY4+SS6QquTxScaL0hBUOJkgtKhrfTW
a3XESHjC6lYmiGgvc7Qr4jKZsZ1cEjkfycecnE5+8hd7GyBYupABh0uewiL4+5Vj
ATKlG2ku10ggV5GmvbyMpIy45U2fFQ/fLkZXhzfIgUTqL0UOSongl5CfAKZXz5Yh
06roK+MdkpDLvH4VZVaCukyxsfM36gEDS0qJtyend6Px+YC7608DqpMST5KIsbUQ
cPgqKmVYDsoMfwa9jgMfdrlNG8nwgogK/d1BHsUGpSALeikNIHeq7SmfgMXy0URq
6coe7KMHrErh1pvLvMVRd0d4XeG89Sb9XdGYZLBYhwmnEybIhOijfzNWJDEr0Ac/
qzsbUODStSvxwlJUIaBeBmyHuHrVOP2kS2O6YwNeKXyg8aXT/uXVjfVq6uWc0jtH
99xstSjgyHhjJ2/56Q5Sj5/4xGuzgcWsBs90XsTjTkKWJVvyxVUzm9uly0br4fdj
dVLpIWaTXG/RTSM1fpg1aK1Ptmr1eNBSWc+VPwW/m8Dzt48y0wXh8dM2aNQpKnO6
dQJ+pFTq+fAG48sajSdDIXjBaR6ZQFVl29mI8VWyynDAL3WGZ9k8kwY5+NpHSN6V
M428yG6NwwxD3LCvVrXhwLZTmRdKnkz6dCONOYttdjFPbwuf37omgi2Ic74nyETt
4JxxW0MNA3WzUXZp68V1+nQ30ZSJUAStR4K1zyENa7qB73QRSdsU6kxWY4fQhlbX
2Ihe5yAGm0NKsJmoM/tGOr8NlDyVMB6qHH8gRCV78DBWbK/gaualq+vV0k/vcKOA
h1yJwyt9dSzZRROOokWb3a2TR/CZgaC6NyUotZWmA5ug1QuZ0LqX6XDOYXlIPALS
fogHQ2uLBm7BtzG1Bi4Nd7/qXaEp0gEWQSBj3jbdX3NywQ+wqDulhWZNDxx0pFwc
K9iKgxg15u6DpoybuNtexqNnJkw2qerNsFeMxbY/yjd/zZMjs0h+jDi6WSROD/mO
EhmISzlLEqb0ufTLEcQKDbhoy2xPkt/9nVTfORBAwVwDNfYppJUvL3w/gh2CgU23
v/0eRNhI9XdODUyIDj1nbTATmN4vnusngOGa6N6OR3vqFTZJVZ8QOE2siNGiA9m6
hgKUS3nBgw42wbgKKEx0dB+paaZM4T64V86dh2olE+4V607pq1IZ9iS6uug9CJyQ
ZslFQK6SAZYhhM0oNunXsP804Z4FvzRSAJYePHrRULxkf8XHML6/CORGmd/2FlWW
9PEAzaQVNDTnmQSbeqqF0/UZUPPEh9YAS4U0WAfSAxVuHpq4G3AhgsnwQlsJz5dq
JIVyBZh4FDOVJKNu+6cOb6ofnnuHGfZkvzAsmIfFa04bDia3Kxln06CYBYFJG+Gz
zOI+IJ8e23KcHyM+fxWil3FVR4C68mRGChGsIHVO+pTnezpkoDSnNaeE9B7XKrEq
yymzKJfn1LSDzoPY/4JPPlGsCi5sUbPVnumTFgC9k4eOMBViL9uz44BdRJt+mIa4
1QBSIkPsaZfQ5OjbvDqFMNSv3n7pWiuaQ36FoFO6AlqQW4ICq/QuOx9QwJCqGGI7
Xlh92oruyW5Wh5NysFvk9nX+tB2Z185C8hftex0i0wWcz/l1Sv2wKLQH/CklfxPr
Rw+ztQPZXk6hpRknhSZhvc26AlCby/wXNO9SFkLZadro1UrQwLYKNDjOiZigUDCT
zQhP65296x1HmLgFDNDPuGnOAQBfWvDnUJX8blgu/UgOuTlrRw86xRhTEgo29vu1
ocEBgWtmPpNI92pfBs/JDszI1F7LvY5w2Zyl0JgUZCs22UeGq32dnrMIZSRuR8XI
XgbuGZ8DrjjSw8eja5io+POGxj49FMLD/kMYQp/tBcGqBKCLMpX/mbn+hpn5yEzR
uDdZux8CCmVsxbVvO3ov5AYOk4NQ5LifFEoeBh0RNfh0DCM39pNDsaTNHiJVOBdk
aqUIpdXeVAqm/QTXzTMHIeipsk3kUTqdWyAzgis6BfpIaD+pxp4FPWwaqEaHPKW/
TBnUrX5OHGYgRZfTLnEKvO5MEDMoxIZT5tNuKpEvj/DUIUelPT16F1kZWYB3oDz7
xgWdPH/xQMgLhuCd793lNBSuu0TEA27gupMWukNX75r9xTnT7g9aOj9cuIhuJeO/
l5NQzZFe/aIY4/nm5PQuqcX+QbNi/O5ur1w1GQZlxrDFfsTw2W2LRRJC/wv28wV4
j/2JcjriGp45Vw7NS+24LWbHVn3i+9Md3RMvfubHCWRugCiFlRqfxygfnar7HOe6
y5wCnkLFbHlawKNSD8AnFCylD/FCqcPmKwWw8diVqmIj6HeSwqHaW+F3kTZYOeoC
WFjSoZmiOh6103JGIQY1qCQTVzO7f/EhYtDn3N/CsF0ohXqWpUbfQY2yF4HMhhld
04+j01rQRqaZY6tUtBDbKb4DJNJnC5oDO2F37tZsLM8xvKBFanG9XoPzEQNE9vJv
nIQK5Gen8YBpiaqxQO3bfUG5uflZSUa9a/UxhpG5HXZexd+Ve5P1sMhOVoQlcARk
7acg5GlosLVNTVk3q1nlZPPEK6CKM1tCzSjUbzS9sRamMyODTbG7xFb05zv/gq3i
4YjV9yehVzoNqvysLd5JnpJH4RiTLsJLIoE5kqi0vEVx92C5mA0YZV90jHezCA7O
jbqwb8YS8BHbSA5UHlXBG4FTRpnxcqDetBojOQV2HdC3KC2qU5+SOfpsPe9aKANe
9bb6xgyCAAmk5y14gEDQL17C3SH16rroC9YbykrBsUgAq3yRbs6TlCZ3xeX9qh4b
wUNjroRXFLFPhBkCqmixvDhwP/3oCr2MA6OrFmREarQh/VEvme3m+3HDfLSzq3en
ie7eY/ozL5DCHihgJ+HdDYrlDvQP3oVyWdOXY/T0dF+yAoAxg749FSiIuEf4USCq
d0xdop3TwjzAdEkrT5dN4wVq9QvpAN4XYd7xZwvL/9nqtBIyfcWBlhhE1D4Yb2Rc
kyyZFuDqyUZMNLcSs0nj2flAVd/kHmi6hdsmH3gP9uTD4/yMgFeelV2G3UnVpOb3
vl9wlnjI4ZH4T1YMa0+oAA2Lgy2Iods7bqK+f6l9j3PrH1u068mjwDtXQ5Fho8Jo
Vgc+MoINraK2DKlVdznbaS7lvrlo7zHwOOUpsntH7XBH9BUDehykRASP2hryaILl
f/Y9piMcg9x+BbO9b9XeKqQmwttFTo0lyM9ymX94YxyjHzvp6natmafQz0sMKjBc
7ejbCs+n+7XcuhKabjHLU1oFH1Mwx82YrWZ9zEVXUeZy7oeHl8Ao42UoOEaNVANu
RHRsL6DyY0P4DRoDowHGNz6EITO/QgNKh892CGY17xlA+yFhsHJjn2DEEMiN1kDw
8Vi5p6J0L3ccDjzmrTSAwr43TQlfFcP90fVAIQgJLYbfkXPlSU5VQGq3+Z9KsZjO
896wjRzEWKVvalHxtfnPQ+zmbbnGX+uIa/UgdLoauKX+Nii4cuAuq+WEHMQG2NXz
plF3FyZjDUkx5zl+sYUA9s7uueXHiSz19EYzHwpkVCYHY5C1iI7sjbh9tCfHnNd3
yUd2gVdePSdSSVa7Ftx513nGUUIq3yj2VBKZEl/YBCfeO2FRiN8Jws/U0QmJpZE/
Z6S0SJSKahL6X6FH3lujpb6F8D0LeG0DtcnXhLrdxcljSUUACHibrB+sudB5YTNr
ynRRK5pxqixvvgh3oXtXIzLdXRrEmFX6Z5sh436JRt4CszAdy+pfEhTslT9jVEfv
T+NAZc2q9m5QNzahvesPBbiO5+6mOGDhZw0PEnh5oyyGnPEaATJv9MbbJ77bjpam
jT/M/0trL01vMC2iPsjfCmlja1ZVAmbW/SdggKlpAK2w4ikhwoMDSxkru+mTkYeO
o+5XxGsQezL6sjXkY6mAo6I+b8pmBm87MX9+BFAtCSBeBMOiVK+c9I5LNY5lieBV
t/isC3Tj2MCLNYBW7phvABsWTe9hRsgTrr7BVtZyRY6IkQt5QSjDA46WoSu5VI4V
imRfgu6YfgXP1YBBoxrT60PgS9xQQlvXfICpp7K0OrildF4eQzs9Iyt14PUzETv3
7u+vUd7haGJw28SIKyOqyc6ZXsL8U00+FEXVpIIj5sXPGBM4lnC+rFdC9JtfogW5
qpHSqpm9O7uPmsrjPtNNguWvSMgNAo4SOljU9f45NKyxU0niac4zRhSOUXtSK08z
yQWbhZidLFagk95KP1jEWEKgnSrDY18DW3OybqWmVwss9aDGI6R9BnI30zWRUZeP
lXe/t/ju2bYBao2YvoTY7eUNUU/ugUxssv8orSJ+hou47mFaHMT9oXzG3tIV82yI
T1fhr6aY6zDaTX+SvKNZCJpN6+YXOTJ3w8nktHejVu3vX5Zl5MUTVBv+W7UO506r
1hSSQYfsugozqiFs6wWHAzJvFymf1OiDzwx4AZSd4Mtt5AtwadDOP3Jf4gmfzjA1
iXBWs/+lIYPdI3jo83W9WlhaZkkHJEMCSbN/lRleChNrus4XTUxqjSCXrk19CJ+Z
7nvbVt3PCEIK5r6Vh95Ea5AH6RId+EcbT7OiW2E+Hfg1elTSCXo6bKKXmBJmwEeE
FwEqi3hC98SwE8qEvF9C/Xsqs7J71fTxHRU5AV+mbih5VDCKR7QHXa+0x3ag65y0
rBsROTEORAjui1DVwJSW2AdIeJf3JRkSUs4FYEkKNX560fe3bbv8GsxH8oPAUYxl
NieaHBywr3DaBpUkhFSbwkzfVfM/XjSFey9LmqaAGsqH2nlGS2QiRVKGgQitb6K3
omlFk03lGnGqdGT6yrIBVcoM3RQhu/CH4iCdWYmqOHb1Vd41afMLxSwLMJPE1S1H
rUpa8zQohPwD0aFmilyg1bXG7/uyEsAc6/tVjjhsJwxdaje8CE7yRhw+0F3BWpOX
662IWIhN4dOUYyQzKgs7qqgT2KQ+K9r6ZMxu0NZRiA4IC91BAbCVZb3FcOOHRL42
/HKp5IuX+sjemPTa5c/uJxMfR3tYz7U1KIPnAj30QSKQK9n9B5TEM5+rUSl6zlZB
LxR02tbT/QQ8qoSAxZV443m704+6VOBKxQTMS7ab3ZWW9CbNDCjes7PtgCZQ1txJ
h5d1ShEcmHil6+0c5tlLLFqv06/6bi2MKigjO79GjvJE3nQwiWEpwaipi+EiuJcc
VILKXWcXPpymu31ODlF8Vi6+rr2ULl17Elrnxxw1AjnBm0kXqUYCmYta2qW6UUAk
2zD02YM8N6XcP4NPwABpMKMxFAEsQJoyM08ORBwJEu/Nf0e48OfGiSq3t0g71ZIO
XORNdAlZnluoY7S40WXMZ5O3QPtmRr8IlQI1r66SzmpoksvDfk8/ckQDXzRUmWlX
PEuyBDK2xLStS3Tpubfq9w1zO08mLnGDwCSVX8XvQGUnNC91hDj0RtZnS7hR25e5
sDxRcOVnKjhZ5pYjAwvUtEHkpFxhTZAoVQLFMsFAHWYPa6zLqkNRgVFNrcWHOgtO
nphaxzhpfMe8q8rVBKPNxb5L6EzZGIsERUBAFsGrQ3xKL6s5Gd/wnzchQztvPqC7
9uY3yKDo533zBc2dJHxsiOYl+OCdZjLq3Hq5AjskBaw/sWicp1DbT44eDS6ZL18h
4tC2PBw10z7tbLtGvoJ+GQ1UTmNhsvpIJgax2KyicaNZD/BNfSKnD3A2Cjl5Bi4U
YD+SNnuDXgL/3ezGZoYYGUVP1X/nryU85JFKGEcP+miWvsgc8tj0aJ2220wceKL5
eopoP2+hz599YMmYypznLYXg3DdsaAUaB9oC9eB5h5uZ9V7SWa4oIce2Vxe3IzlT
4p763M2jRjfQkckmoE4Pe4SOvu8YhStzP1/7WPdWBhK6NZ8bQl4RUEnBkrC4QCDG
PcgpCBJsHxA5iekregsejoH48LY1wl4JJh2UCYlZgbkg6VCGes6uX8s1S4GomuHs
oQ8POtDspnrN6ApFSHiVOvAx1KBfrvjVEvnWOykxNYdCA2U+SoHV5L/7TJ9h5/1H
ckvD0CoGKbIazL8VbdS/K03uTZoXkuHUIRTIY1Atp50lc94tVBF2JsB/R+gBf+M6
bUDBsRm0KXHnVYIinPFyjDahBDJ48R3EhgESir8J9P4ct0uOrNJXsDuppu8CbCvi
Dt1yWo0/s0GdJfiKbCA4EZtueq0x6KYp/xH2aBA5s2b6QeHgwcHATj4K46jl/3zu
0F7V0SBqhGqaYboMeftP90LT57G7g7Y+aesZ3fdWG4V6+cZy/vOnWO2RqPOEMsIY
v4DsVEVZBKOP3Kr6iIx6Nfk1HxLH43/bPAG5MxpcuZj7FFcBYOnk3EwgOiYBbzKG
8FTsHO/qpaqxZrXT1Bad+YnzdXVqlEYlYAH+a/2A8+r9zpotqGzUO8pne1n63AZN
SPc58alLkLMN1xXbZA4NVagQ45uDPqu6VHUVnstLZdKpJL/8pUFVKn0e5xHU/knr
MjP8A1coRvoawHf1PgIGfXEiTazbN4cXSAqr0slumvyUrS3cpf71cuTrzl9P8A68
hxe95WOKVt2hkDz9nCUjFoLQKNbSkuB9TZH0C8c967GjTYpEWNHLKpZk5hSiFqur
T4AxT3AMw5Gj++i6UDxXYyccvrDrjhp/GTj/8U2SQEwvv8wIRkURA8otFJ+xt9aP
sENMTsCfdTR5e1IeBVyFOV84G90soHcMSHKdvbQvpDUhYFWvzj3RDbG8KVaanki3
UB91spijwGS8dMiwL1ZysObis9f1wf5dAAx+4r01AWM7IAkDKXtWvjS2VhqGwnJj
cdus4nFGk4rDUEhdQnBbJg8kFtxKiTDNCZbmWEv9rVbrKHMSkEErok0WejkiGX8k
0RLEFF5oz3Gij0Kds73A0U5+Kt0GUl9Y/oxYZLxttS5EIBn1KiSs1gMGkOcpzJOg
hwN+c96HGeHjfn2WfH5/T+VbtntJFDW/ixnICDHxSqXYwW4zpFmBXcxGgnc0lx76
23YYlTxtJLWgIQ1sXGj3celUolsCoOdMjWcYm+Rb0pjG0/q3Sx+fHwN+TQ+PsYrn
V4+RejwBnm8onh/cECNb3vcH/c53SvIleCho4lytjXLZl9ZZqaTZRiNspLphEyMd
37H5FcdLRzdF02UdqC6gNZlWPiRLl4B6mpTb669RdXs6A5bTvTF2TCC86y7iayL0
JpugmxmZ5KiqSAQKyHZwdayDqvrw8VwpG59k8w7p7u4DBWy97hzEJBSbaW8vkBue
o7zeWsk+8ZmPEjOST/xTvY0HHOEh+gNEcSzeCNmYZVqOPy8e6ltpKxhaUeV5ZWMu
5yQwO2lfFhgirhH0oNfk+/ovP4wFu/UFo9KGMCnAp9vmRM0OLvX5AJTL/dZApovi
A++lUGFIpEL+hERsOhvJL/0i9mKhsTpGMvPKrsxhdkPC3VDlRQUy52H2dcObM4UL
ZB7wFOtE5sbDeh61TGvbTJTY9EOEeRpyvGv9gJJjjd1aVCpUJt1/iLHpZi34C5m6
jDaj8T/YowoYQ9z6ubg57602n/k6WyATEtFCAvx21VlfsHkQlfltEV7SB39I8TYl
thd7pV2ybfiHkeAWMbEBE4mW3LWymOsiTsLHK3w1ktUVRAcSCXfkMxehOA7kQBxR
CExsAHVBVNrpIKurXEDjimR2rciSDUuJHtHKiGwaQaIwrZwVC6zOVGPTc17uwQ+T
ynDCq7shlPOGkOwiOG9Oa+okDFkcBJsDeOJdn2axgSsTsboDwHfgEOlbyluTPsUJ
zuWEEzk72LookUUaOhB7dOZuPbkz57VHMlkO1oVtWANGO0M+TQyZC/TljNdc+t7G
m/ncTrHtDaJnlnngUAoq4Zfs14/AIRVD7J5/wP0nJNsSsmdNKmddq65KXsoOIYKo
s1CEmnlKJ6sskyALyPzmszSd1uIRf+gsvg/uBIu7JtwpS8Xm8c8Wn+bqHOW/nc2L
ntgMBwTHcmU9Csqz30jipuUdZqT1jGuC6CC08fA6F3E4mYCkWHOAQdnIoPVHpVel
cBMqnW+XBUN+PZwmLA0L/0OFSIDDhloDYZZOZYajHyHZ0Ek8oNdo0IsnYx3KKBc5
Z05nKqg5jpAFhVxPg2JrGB2RjRLre+U6FAEp09WgnRacKHVdZa8KigvBZexJNT2W
Tr/h2BaccDZcYlk3P8sjC0UKBfgbaw1fCuYY6SvSrgMm2u476+g4KqClqve5iZxy
B7IBX/uUpIz9YiklhFIM8AHmb+eXTPlLvXUOHWR3kexf7WtzvuA4TcTWFk2oDQRJ
uPBGLqn7BfZYvwX7kPBbVRGDJZgB12gQKeNQHqcdCZ4ZRc0r1etBZbqwpome3Y4O
DVycXoTNA1GSqflakA60Bp0GAQlXDA+cSNDvXuliJKeQx3YJGvZj8ASi30tLsLmz
7nYlVYSjZ9OBxM0wB653QR6JLUtF5TqWUhencxT1Qc6BDOmfgzNSZt1E/a/jY7Zh
isAlasRX+rAG6dseJ18s9DD5AcmUM2Y4bCVg2JE43rlsCt3h0aw/t0/V/r1I15hp
QmGM/8VcoTz4g/MU2gxoaWQn1tFH1JUhqGSAUqXrw1QoV5mvgtBm3Tj+q+nsgYKL
bZEX79EAXz1IMpUAuHdXo7E00x2thAczIQ8IAiU2h0mW3+kUmnPeiMpNQvjPA76L
UoXncz1ImEY4EYBTRZ1Mk4CurVSB78rW4eqZv4O38bfe+H9vFf/YeYSrPYw6pKOy
JXJgmu1nnr9+Qz+La6WljBJ38LiUlTGpADfZYD65rlW/yBc0pNvlMChV8RwmyW6N
Ez64T6HkXep+EFy+aFQ666Q2INU2KdFQeTu4b/UHX6mcdG3oVBmpBRxwuvEiNiQ2
LN8Hhx4NaPt/6NlKTNT8rrX/htDYidyFn6ngqJcvMjgs3JXFAi8xdzREIBU5dmwr
kPkef5J6RxTe9rGAuritP64kZSN6Sp6LwPdABJKKLfRhn1x8O+ZoEqF7f0WDX/eO
lcT1PdN7Fa30sFGFqrlEDHPRYCfuZfmHS+N6RcdDdeqR/953jdTkZLtO2yyP0pPY
u3plVqJuK7ndK3nmgbdLSN04+DaK3MRmZ4AcMUx3LS+g1PuwcUSne55NGy6/+pAO
Rult52hEbjsjoHPhPqFw823Zt/RzC0ZQviBAvg4pdBL5rTeAn9UORGf5p2AxGU32
gqC3Yw6lEgxuxE9u1GweiPrkeYbMSk1S8TYKOU9DdnUed//7wDVg1D9nDzUOW0XB
1fvV0iFKff4f4I4tPnqxEp5tt/a9zHuBEhhnTnMW5sBKF0K+qBCUPafMLppQG4Nv
ntl8MYGhGOwFbQor2GmZePXWqzRlnI4J4pJTL2Zy8joBNafX87MfFwveaYX+qlpn
oP9Snz4Qt6IXuSj4+ggIXDt21EwoQ0zaNIFRoXE3r4QKT9PWr+yEM8dwDv0j7F8g
twxvDobgc3c17XDp9bNvLH7GTeqQ4CO7QboTl6Ag24ZegXD3hLaIzyleOL0++RQL
5uc/QVu8u5YwNJLslBuqQxZPKANsfBu1G3vtR7KWHaCLlXPSgdfglaKyQSE8axhF
3nL3yAALBFjVozgfN4fbAIgnlUfFv9iKuVaYbDU7OJIMkmtAIz086aUYlBUKeDiR
qIpX2oMA+5r/DpvMoD9GmpNG3UebCS+/5da3Tzf5iQr4xit55jmLr/ccZbXgygWX
jkQYWdjTm2LIPyfqj8cw4OIsV5rCVofLIxlwoVazEqaWmzcAn50ddrDQ4Fg7fvWF
OPJoBV3Ej9vFWYJsLNWWDI+WKMy8nCaCqUQzOw4g4nvpsouTkpdtCYHX7mQcHeXu
IBs2yBAxSKzM/7u7dLofM4ev6agxKjKeUc0Fu32072wCwXJhMx25oNuIWHdfGhN3
t6F/xotVlg18iu8/SIaGt8TonDaSpCRgQYZBqtVSaUITLdcxkjjYitq3xbWfTBL+
4W1NSJ4KROdfv0AzndsGgO0+A5XQkyTSQhKhwBzmuGX8XsXaEA3bcI08hkYZchPC
A9OZQCjQytYvlua/qvSsXBCb9792O2e3pK/A1BAInPMM0+jBjkvwX/NauW/UiZL8
cjcGvkK8zG+BrZ0kM0vNEBiNz77aSPjX2lPN9ne5hrRA8Z+IQAQefMHs5Rc6T/5F
8nQ/oNXbDSgaR4JbVcJNwc9ckdV6RbRHEQq/FhIwzvSkKb36sUD2eRGepgH7Aqra
7L5kQuF2ClL2w4vOmPIWmJEwUP7n2y6UDrPYe8U5AFLylsyTamcvsY+b8umEPOk8
hZV7kuSWfDXucbF5ijBHA6d+/cJRwD9wvepyiX/sU1A813eQc7drVhMSAYgrluGF
bFKVJGO47F99xKup8wW1jdzSeal/Fli206OKIhOZnTCjCtXhvblzRjxkSZx6oQsE
x8TUFj2fmeQWgXmoGZ2ohPyYuREkKxW/yu3+UNCoVAJGLn93hlZTuaege+JUNJFB
jY+P2mEfKAqeVBrS0vl255SmA2uR++mu/t/XeVdJthx1AKPfMl64hudRPQAnhE06
uDRC97ou79+i/m3MQL7qWUBQkafoKvWxySDdUMgFbjcWHcHZLKxyBxPoBgJhXY1V
8+dcvD0TmaYY3zV8Exu/uEgnh1Nk7W3et6Zm5yhCPJ2S0TJyqPBh5fev7nDjsiND
SK2J5UYTZFNSLNEz7YqPMB5gxEjx/3j3HMkbTqMui0OYb8tfCTMgJi0q4l6xbpHC
DrZdEfziFgJt4It5GuOYq6EyErQX3NKodsmoJx10iPS507faQbQrikuA6q99fUNv
yXefIuQLQst/Jv/mFy2H23SIA58NWY/OUkNj0TBdX6zmpLEqoS8xrGsOSPX3Vpv+
T0NFg+UzCrdNIDj38WF7z67qcBzLwIakmp6/Q9Qg+g06cQGPNGvFko1VuA5ZmsDe
rn2svgaWsS0sH6r/40ymx14eKODJnDHTJ/hcwqz4AwTfBOrN7W6E/CrDjWsA9DHl
3iko9GislqH4eDY/Ngwfvpe8W38XiLD6diH9hQS9mJnQcPaKLD2zKiAQYgSbIg++
WVY0meC9L1FNEDdzbyKZxvY2haGh71NLH/5okGloQ6ebuVFBXM1xyZEoNFkRrEAi
lD91M21hKmzii9dbbgrPxadtfOcMuLhRGXL5hd4II5FDMXu5P/YmxCgcPV+ssgOc
TZI/n//AgQvx6urxiBm6WpfXhkFos1fym9IB6m755ygf3prZJpHZicue9JvEYeA6
fPRGRORb2yYQ0veDUzBoUc/ojWFiG1O8Lj+vsKpjDDM8MAHuBXnl7npKIxDrfTLC
WfRmCIYrsWDZckPz+1d8kjY09P2uBeDOuIQUxg6GbscIMG8O3heLhSLhSdV5/Nvr
nk+qCP/ecgrtorz9DEoOW2Uzk9UVP/yjdx4TIe/9fviPZN5SZmizrauDA29JIiJK
la9+PYsAeOWSoDKqGpABJPAQD7kwJ7QIM7wLBnZIrrNudCDAKaoM0yIIRb0EkOcB
wDHdbJbWtjDCLLsjecZBbztoxL/lB35etWl3AKzGKFBKol+j+dyFvoDC0RD6Nrsk
ernSSBb31cbZUqtLmwyb1kdYVMtWpUjSgWyAVtmZUT3ncTGorlKfYh8HW4lWXCIH
Egod7igzlXYcbN8jyDeBo1Hr3Avcx4a3PLaTj3Yes+2g8sYtYDIUynE98Kpai8zp
piJUhhoj/UXDpHNhrNGCt0XxQ4YoBCEQMCbSo7qCD9QDbYx74MhtTBXsePjNP6z2
nbF0+UeERCfBT0LFQDv0wzYQdsHmFEryDqCHn6rZMs6ZB5/O9QthgrTEoLXkT0iG
wu8weY6vWJWgzS79mX8oFRzox+Hu6XEJQdVAmEVipL8L6+CUvnfEz3TNxhN9BBFN
EOIXReGBxENkz2AhYGyhmwEtDApxetbg+ElyAy4UpdElkh1BGiAD6RkNKicG+XdH
ax1E68DfFlLX5CZAAbD36R3ctbBvMPwKr1d6p+6PeUDY6APrZ9CtJwdQqT9rR2K0
s8H2Uwkjc/XN9nTTHRg0a5pU9Tdy8T6ZwUYENu3qrzEOkIL5TdR5Bcbx3Fw8DwV6
e+JUaEZ5Ns/g2AW9tmNYn8ONsgP4hiI5TP/bab7CUeDCCkbY5uBj+6ChH24O5A1u
G8MhS0BKDTpl3ajFCuYOkEuFYdxnyyIFw91qxiJM49N3XlXilhyt4gTzhm7vU42A
fwgdgh5F4BCIybQI4bjFcolxWnOE2FuN2iWIkiOqo6IY79EM1Gf0HOa9kQ99jMdS
zbYX03LAw+s0UZkhMFhwQ2djtqFUlwar3QBMwIRkr3gLGJyidtqXvV/VQVIVAUEH
jtXQ+dl5vsYCdly39g/6sTFwpkxa/v8bR8v1mZqZcNs3z0YID15PMavf/fAX5+Yg
mS425hkNg6dHHqoGs23On6hrqgZ0Yp+/JniZYs3Y/0YLQCHHo+hBTiXvZ7ZB7GXq
UNjpPw/+JniL8tyxW9nwNFXd7DKMgnnOopIXbJaHcvO7/rInouqgqdf+DgBpKvH9
CbJgFrX1MZUndE73AlEk2zDTUuLErL44XRHTuzFNd99qR4XouzOirll5pi/XLHJT
9VMmkoGB9NK1PlnmYiwEZNfys5uexHoxnZE2M2oKV+mfx/DemcepWwkyysVnqrPu
I//JvccmQTe25U6uJKcn4M6Kz+T+HPRg1AoHZVRX1XawKKzDsSw7qKrn8n29Xl9n
V1M1LZwj0LjaV97omUjWxTsq+QPb8bln+JAfacHeOgwyz29rE/CD5KnWQqM8PTCG
HcX5ojkVMASReB7RKk+ToMowj/BvpK+z+xvzs8t7Y2YLQDQ/PiVejuzjyCB7MmOR
QBxcfwnuvCP+7n9f0XTSg25VXQg3jW38uVWeGx8YgT3wZBRyyzOVFmbjmvkryKDJ
cX/FF4FjPRPJHhCAOH8bmcc/CEJVFHFXFfgxDVdtIXICfFI2A1wxxtSmdjszsesx
TShlHlkpZKBu+imb+b4t/ycc6EES9hZWQFqV9K8gi5U2VionEm9gZ3SaUAOImAQr
Zbvi+LIereb6AyFJdov4mtXHPI2zyliFckmygzR2dnBaOdAryn4eK9/upDp4KOkK
N2ErJUfza35Jkl4Q20pqu5mNfUTz6RSAknHoCIuY8NVmPEmxv7JLO9LBXI4ygLjN
j7y4lecS1kBZgji42yguRaJR4srfHb+QFSTWHLtkcHz5/LHJ4tv70GpJCOANF2ke
L2xnPVsVbrkK5sciVM70S0NpKdbyyjBq7+o1Zat+SezBznNUx/BgL4MFu8UHdmGK
fnHKcBeitYE3vbgwk9TZMidLFrNNWyHK72x2UGB8BGXfmHptQNiHr81UJsV8p26s
iV8niQYpMIR+bQWLDtPVT+1z1z+EX0Uhy3MdR1+hAu75WFJ91lcdY+uA4UTySUdj
ZRvJbdG/3Le3nS27YSToPq5yCIbxW/u0yNOUeITjL/n2Shj88+tXiiJR5l8IGgBY
ZVULcpZzlcK2KqxQqzmXpcKwhU0Nc2WyaJgl2aGMKbZGoitzAW7YO7aT+Az3S72H
dAL6piBxNNc4ui9tv2CuTB+zVtIWXhg3gb9eGl8aPAoNkJs1eBs7wUvYI6eHsdzN
8vkdq/Nfgr0JolbT3+DDqVuRdjTb+yq+OstXNWd9K3rpQWulVYAIYZYbqHsGOZVy
R3mGsVZhtVIGudLBL5WZCx7EjC3lpSFMdChznrsgjpq6I1fqGhIjvwLYzHIXA6JG
pao7BzMBk4LQOUqFTmraS/m1BhdXc8pGFy29Kyk8iMY1LWzobN0HEatG5kTo0xtq
ErnVz3T0Q3TPZTLyqX0VFVX9XhnwxXH+glSx1AdCxGSl3ZynworxwUqTexUSj9zC
j4mZfk+B1+5m3bVAmeqE606u/PSiIEa+N2TdH/dVoOVXpSVvlHVUWdv6y1s2o/P8
ihU8sv60F2ZwLSD6nNh8z507maLaWNmAyWC43OVLXIMTqAbFQanZ4cZP20sesKcb
LDinVbLL2NtdqSC/HR/6f+DIUI8nBIPO0YYT5f4VlCMhOtDtpLFvk3b5t43mxFYB
36l+1Ziit5zTMTiuxYEZnu5HH7aiU4zbgaysBs3UfSsRRCyQ7+Y/R/6b8bTQJwKE
pYJBGQYR3YvqaYp/dn1il0RGCsJYhz/5hqGeG5zLR6UDW6D3LENB8+yUd1OtTHcX
XdDO1r99+GBTkgfoWhfh0HCMwecUU1zJUJYVA6UjqpAFuExD1jT6dvCaapiQUyDc
PlHOdOs7W0hax6lqL3s4+W9O4Qf9CwA3B6jRIMHF/zSwYv1fooB+Ovtzv1/3W/PK
G8Qz/J5YrzOOYwonB21W9E3t/67E03urcB2n1n+BUB0eQtdZlnbGPhq9so1Hg5f3
POmp53CbpPXwTN5mQFNwEveZKcPodRn+7cJ98vu3sgIaCNkrG+lra0GWYeGDNqTi
y2w79Yvpn08PONSRIC0U7G9nNoNh3KkBC1w09So0gX5A3oi6IIm0Zv7kSthqUteJ
vkr3v35csT3kfKV52AnEksdrRmMdsyo2d7spE+VU+Tw63sJ1rtDn4PJ9TaeIyG8E
58gYGDjhe5OLbCYgmzM4tQyNuco8MLGsT4fyg8iG4MDNzdvRGjU+n4EgP9+LpuId
VNTjyoAoagBEIm+m6Hnk9yZLnWJwxZK9SiV+2uM0f5a2kQilAtvsxsd3Q5Rnrg/1
2rens1COfTviHal5wU9Gt6+3Q8Pp8M/0HYk67i48DkdDOUQHtJf86zCUYGWFmeSv
/j3fOfB1C6FrMvsCLdbjiJK9RAksz/wzlXvLmg+ncx0ps7Z969kSMPJC8XSyEkP7
E3W85se5gv2Rs8ZeIf6RM2U+xhJABlVTfUqGDOYfe0jgPjCFi/PZMERgsxzzbVNe
Vd280trqL4A9vJtLpshi8vUeKM6DvBKyPWy6+AUsRaC+dPqAOHSKZiliVyLfSGit
2lQW+giXEFQJ2pnqCAo1AZ77Clk43GgPprr1yFOodiOHc5+WWSyPRQB4aFvvGffp
wjQQfYFKTg9PoCTZnNxHFzDQm090hl58upvPVGDY7kAhhwQ43p6DDdiN4CofoD56
KajiS3+n7craUviLNSt0wtKp/new3uQhi4tfmm9L2RuBf5IX9lmkTWmivfKgRZWW
CXNJMG36Qp8RsfNYtF4gD1QibyBrNaGSlm81+lqDI4TmLCU2Y9t56t0Cjxqj1aau
TZMvSoEshwFtt641p+P+U1iNCUSh8P3GXcaFOU+AY+XBifaqg9AyqoNo4dWP6h35
ilON/bQ3k8uX0ZJsPpNi/4T+xzsZgGi64u2zMOWwAP9ECkvkEVJ9qmdQNaaIcz0o
sFwu/sHxVZMjH26+CWts3UjfZmDGqWzc+Qja7mB0e9w81ctsX36By9TvZ7xXqvZg
tzrQ9ZyR41ViI32H/2aNLzKUUqNM6uu8HPxOuUVEK2tPZZzrjgCdDIQRC/EqUGaF
bJzgAPDzTzqk2nru31S5jSEi3pWe/jLsv79GZI4czRu3QQAuasYhytalayzjvAdV
Aeu1divNH6kOkXYfhnBzfUZUU5EGlYOIToixa5B8FP/KX1SMCinedc/uXRY1mEcS
8knVUq+O4Dj5tGZ8isUm+s1i0UVCKx6Abc1Q690bAo0LclENb/UnM8ZsKxaHVJW1
pAPD4wM8ZLPwjQbebc2eft3jRNLLdxxvGOk4v77DpFbMZZ59TpHOIssr7ElCYF7q
rnNoyinskxUkVZBZGN6RgKHOAZW4xEzhB0EB2TUfkknpuTkGQs6AjHPHdc2lkZUp
YkMxbQe8QXLzO3f7Wlds7uitxHMPBrfjHNCufMl9RxoEKlM0G//7CqSJVjErrp6k
sNJITB12Kiayjm2hgYQdGQmXuP4swlnaT0q3ShKOpW+AIPAa0adJZLRJOQx9FPuM
vmSd7u5nw5YVDZsoY9b12bRTEi4FPYaRUYWejmiwVxquZMy7SJf9E0bi7K63v6df
kAkuPuRRQj8i2XtGzzeB8ofg1tFeG04Jn1XHdLOlyeb26unnPRp1EEGeOTPjgpzB
ukFC9poMN1rOhrSfP2wnmwW6JkihAKVqCrGWMjkhPf467ekIQc8N8QTOzoLUfvzb
D2eWP8zrspJoWcDXaWztbJh2QcIlR1sunptAk9p9QqCa6C+tkxCHxGsje2pw3H9H
X7tJPC6xaiGqCj03WRU5ICJv84UzOmEQkFqkmZl32qSnUPWjdksKHtHtvZpJ1Ahp
V4SxaEj0NCEHZOp5qNH6Mm4oSqqasbIovrLC6/Bxn3HGF8HR0zeqDm33urSxHltt
cv4C76hBATiBvHE7hpuOof+7W48h8Wzteie7hC9uyHnCyInmKYdfjOC+NBb9o+5t
jaqx7ZY1F/gnv2PXTudqwbqDJhlqubsnt5nfWChIPUb4oM4SzU6dRq+9dMI6Tljh
3QSkGGdUSFWxqqKLdo3XMxz1SIS0jNklurlS1xCff2s/IVCCVmo2LC5OxAjL3VKG
lGISr1MhU65EjemHcUywPKEjDlekcqry+C+tZKYLRayc63Crh2y/VuohBaQDreBq
pfJx7ixm7Z5EqOeG7zVp0XuUJWL8sPEyozzFgkEVmZDfhRbFy4ZGqpinX26pzeO7
x4q380GC3flcp+BUy5wYMZTa3uHOfS3KqlWWQkPoAtKzvqYl7Ae3v4L6qeQ3uPS+
Oe7fKuguJB5eFiEBELbWm/oPF3pKVkW8aGT4Ayp8IsF28MFZug3zypF3jDRq1Hr/
07Ysphnq2BIc7EOTvjSmdxWEyRHM46uA/NVdxvS6ER6XiP91OAn9ATZVNCsDwtwR
1gvQrjUnoZZrWp494D4Xr9Vihun5TfhWPXTF4vKQt5WbPNM1ZU1V3TvUh17omQnU
cpVk8dPgC9xtIxnoiF+uHdOi8RBNgQuWL2/W9d4PCIINL/wPogirctBO7jF7n1RM
NCov/6i1VoQ5G3Au0O9rrZ935l5oYqf2U3V2YrYSYC15L6BcQnxtZgV5A1dR0yti
Ka6Td6/uEAiC9ukegjyb6R4JdB6O6KqAmyj9P6kPKQXQjWRZJHndQwPYPEc5CIIR
dAYKugUgt3+SmX+tcxxOcyPaLRbcoReKANCfofLUGJXkA2Xui5HYJilUJTY9Z9rp
Gv6MUrtXBXmE429i1DDAEhKpwDUjVbM3ANTT0l3dOkIMZkp9ldXc2xKaSv9Te/CC
oJCFFeR3vahVJokB8AzmxV0Biim9SeNymP8YjDYmTSnI7ticxuF+meKuS1Nej1K9
jelz70+zRuarvvrF0tZezOdWukot3j+FkdD9isXBg9HrruSOU8KMJXcLPkN//8pX
CBumloao1pVa0icBduOQLSZy8LfEO52tUtUQV+XCugBNorhvsWgL4RnJujk7TMFa
yTebdq1DkLbmWLWZ6pLldFsQvXOUhtcOHI+1JTGlNC8DkVdsFQoyCFQT175yLjWV
iNjj6TQcYqtBx/P4TkmYuJodp30AewEni+Q6/7oQ3naCjbsQDQRVuErAWIfYrUc8
Lp8V2UA0dvMambfGqmQQlgjL6GWFY9samm/egBf2isdrHnwvZZ61BGK6RgBWQxun
vlnPq6QCIVreIPzY+GiAJ/6w9IyEClzN5agM1JfB3IL3PCrcR0Rips+vumMlAKNb
hYmtM0JlcA7BWzk4Q1XNlqin9cAtz4e/WFOQApDtL+50x3xzU3fZAvykzM3VylLD
jBXfEAkThegvehEXV9QU0M2j+P01FqNF3Of1IFxl6sjOB/RK/I7EB8TBh1zFq1lD
OP+oCh4aRYGSV5a5NAb2Jy0oRK07ReTNUDNrLaBmKo20zxM1eVdVsmRJIaPrIZT0
Eq1M+WjlBHkdFrUQ984xjNdBzJPKKU81HwESbU7S0z9mu6hk1zhKoq1a6FMKeDac
H0MWNkl2JsRS5qrQ8T904O9fnl/PHYOCx+J+y0Xa8XzUmAlP+uvuLXG7irvYCwgH
0vy3nlFAktVhrB8OxoJtdfsixbrOAQqIaNN7XwD3f3fSznYbX+kAJ5LZW85ao7BP
sIwx7PMeQuk7PUT/eLdQ278X9cM+WKkj+yyq/PWIUyHcJjg1hpewjsqcGQr9sNed
/m+h5d/3MehYeTi5xo7Xs5VcqlWcJvLrAuxfU692ewPUbfgS5fJ+OfNB73WZ549N
vjPLsyt4GKEP9cNSH/pNMjAZYVu8otZ1F+ruWLTLAyriUdJn52MHpmWNjzLVT+jK
OtMQKxM0iYjinV7uKyOR2wvUuy8ObDLpFy9i+2Jaw37nVXivLK5xDI7tPAAfq68U
I2r1a0VN5jWLpg2WRjZ86Rfd3lbxdsAaRB+HWBoMPJH5XxVxsXIMJ5q2Lg/SfsDi
NmGqzE6Eb7pKXBhLTOYdmLPeXhyL20geqky1h28i++9uxxRh5yQgcOJhPa/8XATM
dmIO2CUL+gVI54F27iTYszTgqnltxvUnTxQMww2Bqjc4sejwPnTTP5hiyaq/XKea
x4L1mXEfe8qdQUmwlCV/9VrKL01/upDtyLkJ9h8fE5v5d6vYcXk8CkuQ04HCpqeu
IEMkMMJVrIz7czTf4y+oqyyonkchtCUNonpu+TFV1W/vPbxcEL//GLFU2D8+Bhbs
Xj0bPhmFhfnfAuCKENfoU7TTNUSomjR5Jr5NwmLvL1mDL0wMDTS3ZXqK6fWcJYzF
79yXBayEg/3otnFBQSNvYBRpYvuhQ+K/X/F8qfHmMqz21iVIN0EaZDopHhj9Vxvh
DWBxcFfAJP3Im13CnsNxhf3HmCPRS7ng8NWMDWf3muGeY5oY+yHJdZGspkf6pNgU
wRyXwN3ZJqE7cMVc7tzR8LdpeLq0FulwOzr8dflWC1P0WjEKN1jLZx9i/jQpS5GG
6J7HM//XkqwKMs+XlT7g9iRhUT3MnGkQb/7BsEIMAZnAdsQnTi2ZSJpZhebwiDew
QFmXLSXBTYnEkiE8fzIq02oUb12drgAx6IgMmbZ8STg1DmWAXNTcGZCzHBzCVlyd
DzBz3TqSdQMdxYJEvh3phlRl07t7RX+KlHYfOrnYprsxT3yOcxNg99Z5SoJSiVFH
BquHQKvmtcyrMiy28T7MdYClBngcH8WR4x0HAlqKvM+4HqF2iVCnFjwnmmwkeOVi
qXYhcwuvBMebGVopAKv9AiAF9IE3+qXZj24Gq7/QZSvhruqi0jG7LZAcRR55ZYTN
AItglQdXXGoIs5PYkj/r3q3ytK2O7pexcSAZHQzrb28Aa9Vp7ZghGl2FGilPaKtz
OkcudKacBLTjhzJf6YOfmwrGiM8F+cjkDGhr2B8CuqGmpHkfRUykoghbDLr5swoS
y0mdTVGco+funYogF3EuKDIHzPXoqLRFfjw1efnufknoMsT7So0dTB1Rq+GC+SIC
xuGHPkiK6N+XfyFCGIg2MFOiOsxHrlvYA0C5Ro/tZ7jhsi6B9e6KA+9sH6AQ84RM
4juYhDe8x/0gogZp9Aeyb4cCLUVw7jgtWsPrDp79jzPPNG27CDXpCdGEV9ECxEHb
14KOr90Kck9v1vlgLsEGDeymt0VqlIYiJcsw2HlUeqMqHEf0f2rmiLruNWQrPKkD
ldblK7Lcn0kz5biDOgMNsgegB+7EjqUjINDhXn9CXqo0er0Jad/FCdSZzaFm3AN9
zX49KZbix30i705HSjG2ROU7RmfDysGy/ZwESPP4HAleHONyDnGF6F7Fr3K0fp4m
94MH2IuOg1b2lE05QHFa+NGwkVcaitrJojTEILoqHHXDZbEw2E2HoYfB0Kp2SEHI
6Gk5TSUUOzSIvwyRbliTZvFeJ1Sk9yCeC2gZirf07ikHEy8Ou6Q1eUfKemNUpOTB
AwBP+KDLO/cQwnfZuVZl9drqZk8NFZhKUYJ4mELKEQzha7is+oyQpgwxWn3ORWGz
0aOnCMS3Kw05jULaXBowFpBwW/kNWcmF/CmLdN6cX1V+vlnLwJxSGmswjaLo8o22
qeh4EI/5wEA1RSssUSYCbU+PqG7JHoLfRac4Vq7a0SJdAtkIWhBHbw9JHZ2O3jLv
Dqsoewcc5Qapuy3PDW1RRbT4ffTqYSzTdz+kcL33m3c/uxXcEs30TohcSAoZ/xPx
3oyohRz/2xHgna83gp1rcIwqnoXqbsL39APAKJlgFdlKVAUS6UDl8cBkgbINOtbY
bwNbulh/4SCndklb0UcDBTp8oxyOBA49WIcLukDUAC/eelS5Hk71mK3c4numIo7U
IOytN2i/CQgnMz0O30UkeutAwY22cYVZd/nOrUk9fN6PmjDyszf/Ya/DhX23ZU/4
9TWWbS+kuB9fOiGd+G7l4VZFBS/0SuA1ZGBcMgXXX3zKOXPx7MXBvDRvnCuWCF2B
bKWxBoO6weOEYoAiPOXCnC3+Q3IeVl2R8s/p9ESyHki8b2LYAt+IS93o0Z++BS/s
yG0fGb608vl0cHMEz0+OxCOK97oXyDVLHl9OwaocTSBfkMaiKcW13TQ+0503eCOx
YzXlewvCjlIazDlTfbi/uoo0x/PmRdGqYy/UC4d6YKHWLamhosnjlH5RRWcuAL4f
MU5DCoPQW5uK9a/zk9DSm1QlHyiPOBZOyLDHm+q4tTmsLa0Z1b8CcxblRJftTqR1
AVNk8q97L5j+LeC4ThfaMT7kUX6lK+etkt0oIQFn9ARWrm2C18U0Ewr+Y66SS9a+
zNqNCVzAaTMGRSZCESLEM6QkW6AxJAu3B1aByqiF65hIpmaVcMFa+rJceYOSiLi/
oZKuYTvh8aLS+vJbhMK48r1XsiucxanyYxRkNU8r6/cF9LadjGAOJtaG9e5o6Bkl
gCE1QzwH21Nn6qLLYH+kYNxqAD9CJa4sDej9/+9p3RklgMOmT5puk4Jq6pQ7xuAQ
uqoGmyOmQqAh+wV/VAp4k6gwfCT5xnuSJODni1LRfkZpJ4LijVL6oJhGeIrsXOdB
H7oAXVfSxWMYT0uwyccI8y5VOnYyyUjdQ70SBhzDrw4wYC89eZXeCAqSMo+sL3eC
28bAlqgLZhvmIwJbKKKPkb3Nj3TB/uMDh25L6WpLT2oP9JUMW4SCQ1/0O/uxIKQe
2H/zYuC4QtOvh0dEh/ATrfoKYIpBBRON3daxFL/YAB/X/nxKsKtDlShTFFc2+zZs
JxE8qIJIqRMbn8YWHGzr6u+SQdF+TWJ9M0/nMeC8QjniVFL1fkl8Dlm4fVJBIcnC
uzsDPxHnss7CvRL2u6F5hLJepVBDcC0byfQZYLyybmtK/KHYhfzInJBf/0X63i5E
ZSvqns0AmKlnC+jOlDWGaAJhweVfSvmrLAY3nKTTdosk0BNV/sNsdnbI4nIF/jj1
BchzhHpo8zkiIjWyIYPsyMzye0O/R3bz6I5ZTri6UVs7HRX1QFBA6m6IF5iCpeXx
KXPS2KHHiPd9f7vE4CZucD3O6QDk+//DsgaXBbePafgiQ9KNsE90xIPv1iI0JycL
q03vegXx9xWrghoKrRNhc7rTmoWZy9x3Mij0avU4whyodt3d+ju7gLLP/m7VkR+P
Q+zfmtQ/dicfhKx8/T2Mqulvy1OkjLW2BHAITZDf5EzUh3Jw2pG4prLiWxDNGQmW
+z9RyM44hoHOLnJZ66mKJ6dc7jwn1U8oaOs+GBfdFxnFJT5fTlkZ2UUZTxsq828b
+nGvSWspORc5wVtaJCc7+tvGQWW6QfsRCyx1kxCv3XZqX43J09PWKzNY6MR7mmWs
UhqECJNc1ePE+Rb/eYpIdKgyLwpg4t2zrYK8G4dXjeq5kNBdSBldlGO2khL6BbzG
bj/bqYS+VZatiCjKCH2LNNgJcu8STv7Ie1r9h4fsN+2WLHdxx83Z+j+51NSbMACs
Ef8fXp4Naobi98vPll0+MWWJQXeigAnsWHFNeNjiPKnAChYz71wuRc4vm7YAwmQP
MGCW2BfwDSFZWASP2UKtHHy5ibXU5odNCgF4WA7OPjxsZEHY1Y1QW3zEBiOtBAW7
owM0EwycgC+5Kq8k+ZF6SRGEHgWLxZQbhcC3FVq9AkDw+XksgqwaIo+WS2rsIwxw
F9NIH65IBrrVLvQ+ei4P/x4ycfPGvstuoBRJCirbHM1aLtfyI64lwaY8EXVz3NzY
leWpLJcu+xWagCyhdBJ1rldNzVQwYJ6paGwwijewt67a1JfW0AA0fv0TtrMfOdhY
gguLAa3YH1jwi/N1nc7diT282uLJQhEjz0QJEts2WtvEcOhwk1wyk33BBeG6n8Vh
eEVXumduxwmXgQnW16HYJcAAGdJ1Lc77sBxrJEiZAbp6KIkt85mJFZf82Px7yzlM
U0O4BqFt5XghIuF9Hy76Rx3H2hq2sL2XVJsrKQTIp3d64w2mz5/h/P3ZmJGiCH7g
uLlDe6H1yRWDsVsAqV18PIhbcTGvVK85uimUS7cXazbshnN0IP0xuN1iwBbEDJoC
xRDFJyVwPrzGf5xF7rKV2q69VEqw4dDBlV4brBomEnm8lbVVp3b3tmgSnUFX1ClN
FCMZXOGRoDCtgTEZ9ia1x/UmZ3BQXQMxd/zD86frczl07U0+ITrJK1vrY4TdiwEr
hxHkBVKdoG4o55O5WN+3pXyxdq/CeKWF9sLskJ0iPRwkNphv1ATr2Efwm29fKSLi
0Wx5AjDjjnga+yNx7U/63VPSQIvIfVaXtbYK2DyupH0n1MV4q+ceZXSGuJXCttIH
wAw+PJGQbhjviL3QtMbUIthVQAi+NWNweKPBjPBaspSUcbQiZVRgoGmwEguBwFIc
hzaB5AxH/KIocAk4uz6sGtf6sFJnUPjL3qAELXbeTlfD+DuNHVhCmPTUu/y1E6UT
ZID9rAm/vlEMw86VAer0o45SbaXsYCKjST0ZctoimSwAc+IHK06v4fF5+C16MUM1
hxSq65VPKkzlZOZc45gaVZ850Qtsbc7QOPKSI4ldIvGMZ7pYRWzzXYxGs+2MN+jk
RQStOqe2n2VRjhISrbis47wJqbne2XlBImbBNck9xk7i2v0+YOh8EIaVWdzNHxb0
LXPbLXw5X/WQFwg0XcYhK8GBWeVTCegJ1vU44hb/CQFbRI8Zw6j4APjM6x2YXMe7
4dhLDSl0cC550ypFK1caT8pe3hB/oZN0Ofnpl2TIZ2G2pYrOgN/D6JRXEB/Unscc
/tSnZ5e3SNXoDSVoTb/i9TCz8YDeNyS6nvmRF4z3XIWJJU7yEgmdtjA5HWiKwuEB
cXpYnkM7smgxIyGkHSwkj39aXFDsk0ZafLb2+RX6Cq+sj5Oo7Z63Y/++6BK0LZUB
HimXHkWOKsq/yj4/0u+p5zhoYTW5qLIds6FaJgok/1EI5gzc6o24SADzAXG0lO+M
qs5Bqy2jCVg1pQ2beAA0Ve4thDWLL1Ovwl1qXZ1Y2k3l4XbUP7CxCEozMCV1fYAH
ysFow5t9oWS0oBfMUgYxiGF9z88WTqVHIUcWq4/JBc7y0m371hr+5gbfjflSbOg/
yu/ClJ2HXhzh5XpScmOXw2zFFfS+wLq37gA6LqZVI8vyGwCGuFl1OpuVKsnlL6j1
IMib/TTj7Hr9nvmWfnz6P2oUJ96WZ81Fj1HQY3lOU4jPO/nDjBvXWjCy/Acq1pnP
23as0ccaEaGXUvt98UrhYuLCtWyWoPwL5xQlIs1pVdhSe1tcwbiiPDVD2bqFdzWn
qcSTwVvKruA2GI5FVC8OmfYBzqjeWzSDkPdfGEVrKqvntE6WoHeAx2v956diRyFu
awjS9hLzV8KGolPLxV+e07Kdi42CwaLmlVow29C/5hv5U44o+subyejv3lGTaVaU
uyKlU+mKTpZnE+KN98tTtfYE/4bHYb3L2Yq7tojCqxijBQ4iVXe0lj+00Ms16U2h
Ci/uxR/hftb1ITjXVPfF0yNNyfUY3I1hgGpMYpY+dH7L+NvKYDoLVwU0+S6yfXFC
K6ChTW7tsv8woiGlwm5K3H3hQZhuL9M5t8HhOfRhPy9fdf8oSQztRqeDs+byjEeH
Cia2zTndR/ma4ilKsl2CBeF/vV7yy3/mQgmGvJYWDY82do2+HOKdLgFmCJN5omdy
NS/9yHJXoYeNd0v57TIORRrqO8o8VqMlOMh8Hwntjv1VhSCE/2K+WFh470ZNHH9h
ihAlm8ohsTdhi5puKgMabiqRAQH1c4iKCqNRTfy/F/2Ecdsu4hWg26gZq4qKmoLK
FDtV5Oa3HadM4srK4dV66EAbKVvtzBG5v5W1Ba4xsNSeV9ivPAJIVWgF/E2vPPbc
GiwlHimi0wPOI4OowHKKs7AmcdFvgbESklfAgmv4jkxXPBSb4I0oWsyHW8ygmiU/
Xp/dGZJx8Gnf+lB8f4Q/pV6C+lULfEG8wGiIti+JuLAD8QRZBfi+V7SuHNTXxgZU
wGDjJ/MBDW0ZuRBAOoG6ACopag+pQB9Op/JpEfKfR01AHIEiTvnkSvlGgHI0+IYg
yMLbCUA/RaPekUzALt+LR6ZwQyxKSt/SzecwxLCSNPuAma4/76jhdhlOEzMlTr61
VUKF0P6yJwv3wVHgkTWhyWtensD65k7qvcTVCqD9NXE1sb9rgNOlxHDGvk67jVCr
rbO/s6FVmO4EmzYl+TdbRUqwWHKojfIfHonO0iJTVaXmtVe6Tc2WQ/8CWcs3h81q
KF0EFOG6bMbUdvhCoCvMcrnDpDGMyHDUpRglAfoOCAcgCFCcUbP9Fk2z+ooB48Ho
Y0LqlDXcQ/7TsnS/BYrLJb/YRLM1+v50Ftc88nUwXjFDv+08AtVLONFnQstVVP0v
C7F4rpCaLZKTJs7FQeX+gHWc+gI5bMbBWVV9N3wBfKxRi4kHJQO34mzevK/noo6Z
a9QKcVu25rJp4YXOsiu3GaJkTAFhsYmUNYLm6Tq2UujcRtbnUvPpA/K6xRdOH2Mk
eJg2jqlYeI3v3j7uYTOd4L6x8i96vCU0VcLwWHmZsAeZDor7uPwNBQPTxvjxj35h
3yx3SmSUELb1hh2pxx3oJ8ZtU4a5gu6wtVsPPn64k7lXB9zPLnWdw0W/TLuVQaEn
4pIGSvFdmKfmhluqVEOBBF9GQ5SVhLUjFPqMcUm+Znx4Vxyr+Y1gh9A1ExVIkQ7M
jXA6h+1zunn0TegYtbby3EhzDHBmWQ5AjS8pp5TN1VUT2Ie2NiU57aaoI0CK7y6t
Q+yUJXcw0Iyngq01BlgrCWqzN+cTq7ggR9Ipjs7IZNkXJORtCr2QeHbl/Ab9FtTT
JBZjVSgY9PHWefbFS7bAMPRLyN3mQtub4UV2QepVL705WSKfwMzmyLo9sCOd2VET
Ow45LDRFgyoxpzdMycupNAxY2dwrKOHhhHLQjyne8CaQXtEkVqSAKVn8NJcMVpav
QNZwm1JdrmUTRQdEb1Gb5WNc3pG0+SGibEC98g+gVVC3Isktk0afmxFsXjwqmrA0
ATp5wMXoLYVMC8kBg5Vo35DB+Vw/boWdQQyTpEihb96RWOaI3xC5oKaOxFRx2ORm
w64jCNY0Sxyd7/yrcPdiHOYfhBuKuEsf/iXQ0gTPdmtvusM0bxwFyvT/vqX53pIk
qfgg01lym+Gf0PzTRx6Md9qNv0q3zkb6GNoZu8IDZXiCvJKiVN3/OaCSpLZ12UKn
bkxQGMng0nIx40Kyde6hRwfnrU3TNPqa+kUCf4hKG0hq55N65Vs8Z4MYUi394fcC
wTB49IQwMDseJz2ERPCyYSVkcZ+t7vU/Em1JKeiz7rZei65hS4/zJXUfkAG2gz6a
mHoKaTqi2gDCpWLbbBNlQRyVz41yaTDjkjpAKoqddX2eZank/1e7EKMxV4QzgdcH
oY7hrn7x1t4gOcCsb6zINE0BDbZCsz2bva7W9Uzs3C0H96tPgFcQQiENR32kn4rL
Ubotjx9xdIQdOHFJs7/D684idU0u6c87Xh7KhLIXOHGzdlnRCULQ0qBf4tNnBzmn
iHVKNBpp0rLHePjK7FgG8eBBkNDcx9XwRJi/2REDLJnkugc6LIifob9bMVHU8sgY
NneqL6o+hyJuw7kZMfiMaRYFF61cq9+Zbb/Y0CM7MA3tKtowX1TSxujzFbO2h8ks
5xbBx7IwZIr0gPiTrwzGS8sUrRb9F53pH3SHMyAGMdm5TzImM6Rpl105/8ujBNsQ
y8twG8B7rWOBrjPPz7hwrdcXbOT7Raak2gKNW8Wwv9+6sun6QdJw3dkgX0TjysOi
gTwaW8TN+rAfi8Lx1bsiMx6BDI0kMQQ9dUBxK6Pa3PykQqeujJXpOVqY0LP452Mc
XXlIP2l5bd1wYCA1gQRTWYcZnbzpLV8wXrNws2QEcjgRaos+Q+3w/XEuKqA/7aN5
9+S6F09ZjRDl9BRAjkqMIjbW6Ty7/P5OO3c74Nlbz/YtoEqEc3N/4KKV4okpNUsg
EHOFJd6WvtrCSG/ZXMI1jGZtBDa6rBeexQ32z4zIijg6K36hkpRD/ns5FfNaqOad
Su43v6T9QTm2Rjnc8Qz5yRqgDZjEEcjvzZUQnd+RWqsTNV0zgBr113ibo8aEctxV
HE5RwYJSLShqecpBttik2AM2/wV9qn6NyiVSrkgAy5ZQFgjVmfWsQ6HbyOxl1D4P
fTRYqn12a2TtJsfKl4jr5lKjxTm9MoMszkzYq0EcB7P0/sS6GDNd8sdzrQaa63vM
qvMZI+AEXWlq5Kbd4Auufz1TMYFs51nSPk/HZTfpFFw50OiiBX1c3p371Vb6adZw
bMlHFQdO8T7WrSPMoXfl+Xkq2SlYHAvYEYxgMmLvY1B23s1YKce1oRUiSmcyVtBB
mHCbtqe39d6X5i6y+SRB4QYgB1vC+f1JS+zpVhmoFGlV2PQ8AS2itA8FkJTxvDAv
qgHNI/cQDyxBXO+GGbFdYZebx/YF/PbWgSpDPP6Oex4uIRlvwU1/WAgJnIS3FNgE
KCiEbVl3hyuvNn3WjBCjUEJGYWdskHkSSoctTmWv7jm5J3mdcFV+UHgXRG8E/hCA
oljMZvIux/SVt5AoZ7XFHdiHRm1KhCVXVO1fdFBvVOVE64p+JWX2KkRbn7M92ER4
kOP/e4MWDNKIwlsFOEaTUpSrhWOLEyzOFdFbMhXEjpKa4yKHtOnLb6mCG0eTNy8z
jVFNNHauJXkYCIjMccVOtmA8PByHjpnWjm18dfSovV2jH6AUxTzwp28mKKmb6x//
lMHhRNAbrG8bcwxT0cCcjA/OLhDNSlwiv7lJCVoY/FCiZvOGdpoJh0/rkaAC81pE
h/Ipq6SnYLz3cWvoN54sJLee5ZkVoXCAslpeoEHnMBYXpcVak/8q7jzJJn32Xc3n
vBl+TkRv8Iz6fxx06op9GdJjZIuWtGf9iWXHMR3OGyNPta6+GXan5sr/aaMbje6f
Yju4u3mRm7Es1ChNy7tuE2cw4yqGwC4Hlfleldrs6fQXqOR/h+Fsx6jHR34WgGKX
1+AzwXL35INPX/Priw+NTvsPIAPwnKn/mB1NBEPuljW+qQsArBwX2hOu/yF/XS8u
t+6jV79oWMh8MPSJXHSPaUJlVmjuuMQaUl3GDQZ0vuhamsyCCpqvEKnf6qesFIYv
pMEYXHti4pv1XVPksdJcPMQLqSheBGVYBjisZuhxVGLPOnHEeY2/Zw3y73SdrNyc
yzkaH86s6R3bYKYGbQKQ3YD2l8x7QDz484BSpwd3/dR0QzbwS7jDz7WYfjOJipS7
C64h1i8v6v4eEejVuKVJrTHxyUYs4uW+d7wDjYH2u2v4w3wL0py4Lkvtwi4bEd4h
Om548J9SYvxElSHvTfD6qh+FfmPPtSHNrXimiUdPgjCkEiHezTlvopWdFD7vqui0
WCz5O8mOnzmx0gAfOiE/fxGdeATYqM4y1qXvVCP1+fEnTsvmB5YDtNAgXHecaXl4
ZpkCTFft9yg63ip/jQ/n6oQN+k8LrTBnU7MF+s0IQk2PMem8aRxCc5pGjGUKOhtg
nq854+IqLa3WmIL4QcS3JnjOAgCHiLcq9Pp6Zvy7RueuDAUgq8is+Bwi31j3dpJW
KLg74krNOhWgMjnIwuq84pgGReJ37zm/yzAPACSd5n0LgaA2PL+qNrLajsDcxC8l
8rhQVwXaxkiA7FIUmrKmS6deJzZte6rt4uDpQ/CoCEuQPSZ+hNbLZCsB5zGwz7bf
7p4BvYyBwjHzBT5+1srPEcXXlc/IiorgUyEo8HD4Y1DfJ9niqSwetiPNQtZNCyDu
Ewuxzs34aXeN1wLtsAQqVdk0NoBx+2LBmemWOUqblWyDff/rgAQF0SB0fojGoHCl
Hv/5FsNR0CCcgGGb8a0cK4hQea5evJKNSRjgqVOzRw3qx9dTGMwQDDl0mGP5NjJB
w88rDvY8LsLBq+potHkZB6TtfImI3icXl7+Jclg0kXmdzJLo+UbOqlvfMJycwHdV
euGENowlqXNl2HFVIWTo7RKjO+SE7mog6hbmMuSfbfu6+YOo+CiyHGcTBZ0MFFnC
EqpOoO1jGqcZkYUYckkVH621mHaCytH3ak6l8M/kFa0J2ItM8N2lCMx5PTN2SDbb
8SlsqZ/1KpxHYo9UgoyATHc39G5UDsGmFxraeo6ssQeB6JIauCUXS5SEMbcnRDwo
JaQOBs44QgZaRw08YfzmUHQWjhCs/zwleAhAoRMe5CmDJMLLpFjsPNKDrchfJWZj
QVeHT1026jrCx+m60XV9o7S3glzdGIckztjRNH6nbUuJOjITpledk5qL8zOtWwel
xuU0YQoWgzDuzygshD0Km4DjGqmo16wsRSjGQTTiMSdebR5JH5qVV7jImxcgtkXt
vuJcXFt1DgNFinSAUFX/DaalfUAn4w1Z73+AuACeob4CvjzyqZq0e++tFPTPJNVl
Ru4r1X001XxACKkC7W8uhkZOE6GRe1zs2yHgPC704yuL+Vml4BXdt0VQkg7emhIn
+7x0CIWXDF+bLmdQ3vtZjeMY2xz08k7Ckgj5g/ZP9CFxvAYzOvEeJrOKfnZLp8+t
m1z1eqmNoj7FZOmR6yoywXdtRzAqHC0ao4O/PIa4eXaFR/79fF33Gzr6tkFsMjTX
RXKLMBRL6QpRl9aC9GtxYQ/AHj9r5KUWUcbN86Qmg/TD8FpajR+FNeJi87rJyiz/
xIxcEMhPqHmnm5wCH7tkxfuC//7IrWaI/uG1WORmJIj+7JM8IuzUXG6HaD0Io1xS
hClrNSkmvtnJijcm0QuJ6W2r1AzObHHvmrez/yb/OkJLbeOvAsF3OIxeZOW+doCg
ETeOd4qtDHiXvWmUR4Frjtym6gS0iYf31xImBvH1PnkKH9R6c2liNypoaWLlYP/5
Az1QxcQ7BarK48uEwkakXI0Pzxax6UY2t1jq3Yi8fCbn69UIcpexMPdg5JD4Q8k7
auaTtiDfmza69FNp0bvMdzCR5W73r54SB+GEqmSs0X/qKlNFX7Tzfuj0WYEOzBJC
ArcbQxuEukdAia6x8xeIuqzTNlltAr52jChO0j2KzZpGxD8U79JIY1cRwQHJubow
xnjG6M0JlIatKdSXOqaZzusV90CmFTsAEMlk8V7T2gbG/lNMuf2o2gSUX8WhvXNI
qv5lXxt8sMIrl3hin5B0+VyQBrMr1IzAwOQ0Pwbs6Xu6qumGV6CrYJ8snss+sijl
8S0WNXRZMg8sYF3HbXYgDlD8OCWON8m8OxsY9IHuHAJtZ0B7IzX6CkuYkk9fhCdg
/I1pmogmWyqKZDKaJ3k5u3BIegNO8NX9x66c5Wv/jUp+bjXHC9vMlcNkhl9mNIII
MevP0PtUjNYbwrb0cc1Qnyf+mO/h/iO3GrXxKPPSl8wnOFl2a1u8ZU2RLZiaJp3b
rRHqwhrUldTu2pg4DCNRIxKQSNUhp+IFoLBrwaqyKXiYokGdgQqcG/XhlRZaAAqq
q+aISzxP8CvIn8pxVkjfhNFlZTrL9jCsLEqC5d46ScxrTIkuZCR/gH2BgruB4k9k
TAhw+4+MmSqE3iAE9z11cNnST9dCMyaSXvxBJ0N2dWs0VcyxI/yiig5E/xhtLymE
VMvh/L4+PLWYUu7llYV+wIn0myA+iTt3N2WsoY0fPpgE5jLW7MHIo0KSBHiZI+Tx
ut9LG9Es1/v6zjcUo3iaMX3RHFLtfb4RWhW2Fygu89SMp7oTyc3+RpEyUnIPgWVB
gj0bNKMtwMRpHPeNRLO04wZbzYHydiGoY+68kos5OwSKkeKHowUEpOXM1PB8UKdD
1eWAsqTG+Hz3gbbCh2dTpDIxQWWGt4pB9MOM88gaqkq3FILUzUx5M00I3/Nl+pht
jkJ/JpTDxDk5qt4Puiv3QnRbtk0AbDvOUAajz1qTAu1Jrs+mza43Yn1Z5QXG8ZkA
VAFBKferyJ9f6i9CK0K8TLLidIWFkI4797S+I+ketrXTrsfj8cuTlntfLrycqW4x
uXyG2P15Kny32JHcPDjuTBVJKHFLMx/mZTltft/c1dDvgD8/SUnoSAecH/wzFatQ
jqyBbYlEnOL63/CDVr/ocVhFxSooF1SLVCuAt/k0WsvlneX/LSQHnmeW1t/g2SCY
Il6oNnMaYHkBYAUXYqayf15a65WRnSIYyjxaVoQehoJpIG6eEEaWemLrfpQejR3S
ZWOYKZOCYrAm/yaHqokLG76M6IupI0Lj7DKKYt5Y4eZ/DrSf28u+PFiJ0r5GaVrs
odEHSFK7ivP3lhRDvCdWeig9CcbT0moEh3UUREsQim4VjQcBxGTiXf2cDW8votnU
dyd2dlRQZ68+coJw7i3AQVqZM5ZcLWOWXGj2n8NIf2dsYZIb3hYZgy5W4vnODCQ9
cE5zp+qi97eZcP5f7KfBr8ycrPQmRCgcGqhTzMcBaLnCnfaPnXj1FeseJnaCZjIN
FVwbCgjPm0OCcq3m2l4cY2+eq7811Ln2FYSxji5Ssk6bgqccC18muoI1HlxNu3gw
JJyoqq+9tSg0ta6D+zTkjiEO3arWmijX+XZ6B1wi2KEoUF7tAzPbkmqgrhyKd35y
3YtnBv1B0Yfv1cvnb79fzZIgQc6JJl351FiG3mC+feu3Gj4RNAmRRGLebzMPo4Zb
zBC9dtgtsK0jz5mXQnZKFsdgH1hE3/TH496TdrPzF0MR10LBPqoqVYdER1wlOPhW
ApdHxRjIy0qKnCFeP0qJsU/ZpQ2PNIsjDRxN0lNmS9rk3IVZN3p+K5YF/pCNfHOH
Jq6WF1PLSjSiOcGf1S/foJtmb7gQU3a+1MRV4eEIH7fpdugvvNsf/zLAAlb/ILfi
+eTGwoCYjFDK1fP1rUhzI7YsQZYOIIB6ZsgIuK0UIBTwko51ImZDml25RAviaA6Z
QV8B7GzH11Zz0hw8L4WBZiFtZYDWYoGvAnNMO53OaVvOCiEZ9hUnxySuKC/KgsH6
tsRqpw5v7ZqY0LQmQGfQP4yFOl+nLnfysa4mwg/bb4FGq9TS7CBlP78VQXqC+bCw
0KqmC8PfdXgSVnsZ9hGbMLPp4ixhThU7KQEfP5R8n3Gxr8+HkoXXycjK0ZFvPsN+
M4Eq4OrPIoemYLfLq7vy/2DEwrhzoiksyLFE9d4bQBIaD1dBXRUo3SbK1r22icM+
P7AQh3lVNIL3fN/aj2cqLEwIXB8qPf7a9BBlAKH/3HVyDo12uiXJFKABgJKC8Q3F
ce+OJPqC8nwSSvYuexGPK7jIhgRq1++/Dr5KgoB99Wj+BJeNPnmH8CpjxYoMqTEX
p4GJKoorLfbX6qB4ETlQuOPecfpCsq+T8cxBq//E6CUy+lKmW0ew4Ldq1xyRlS0L
6uQbW90gNmxdJXpZtkGTzhypN9/eLGpusrvVy57ymj012l3lY+Fn9XBowOANLeAi
+Z21oJUSwDefMMoX30yUHjATcLfebn2bY+JWmRuerlG/Z8G6RpzLY1dfdUl5h6vJ
OxGNOGt6DlDCTUuZ1F38AJ2j6RDqPIzCR5563vuRPRVsfdnnAd2c0ipMVpSewwro
466FFZrs78JNYtTrN8sR7LiCrxRPjT34r9mj+Q7gwZcweHRdHa40PzJjxfTRt5HI
tvYunUy6TL5HN51FCxlg4kQ1ccoes/5QfWpQp3/40M42/PiiOXJ0orHD8SAq8AOp
HHauyU72QWOeyBiojKjbnN9I86gZ8hzUTuQpHmCO64ghDSacSkfzQkwmUIfatqI5
zTAwoPhOb0kYnACDkmbop+QmW7RuX0rRhDXDUR78IP9PFM+w/vQettAkPvkSgUOF
tkcmrh+N9r2cCkkoc7mOGEo33IY2kDJ/VEUEXZDJXjH26rMp079wA6oKvjLISFQm
mwXARe69WEv/Tggqi1ZIyBhDSUNcahvk9/2gTMQPou00aZgSZjId9o3qFg80VueD
409WgTUOV6d+29TiMHrAjn56GXIgHFLvqkR7MRDIRdUoKqWPqS/WAJERRJ7Ge4/L
/AmN3xhaqPxAR1eUz0TV4NNzSWyAfBqKWKOUlqNCtXEcnlaJ8cXhoCQl0nJqI5/X
g3TJAcvQQjUyToLxLBpnQ3QKl5zjOKGwr+mgiFIIw/yStuWXfs8xOFevDWfn8vnT
JWKrU82gvFlG7/n8w/Iyrg9BNPKPr3wq++Q+bhciASEeZYNhCivYU60bljFHnRMe
glCRlVDiDQPc5zrxY1GCBuuJbRkaSVOcNuJkXOGw+y63X9CUMfPD0Efg14DNRC43
PRU03XDkzK51116H2Y2zBDACwHTZYoiut7ROeuwd5fCbVwvQx7VnCE4PyaC7M/c3
n0C85LggM9tzgM9DvSpQ8Mxkq9MLy/Iahd1yXKVoo6hyrqeqQFvXdFs3Z+nfuJCY
xzvHBV1JmGi8GrfV7uxoSBMWWyh1dsweAlrb92x9AT4PJTcjaNQaHAVc0cNINMYN
3AsgWKcv+pTkbhXvkslhwMvVORU3j07BgacMfQvH3WHWHV6mrijewURauRs0XRZt
7wzbe7ffENMejAkYvpnzNLeTytOO6ZGQL2ghUekaf6Q6xsoFkBUEfwXUHAdCy46G
Xpd+ymCa7vOBbRhh0qngNLCibYJt0vvu1ZpIDewqtErsscldg9ed3Oi7p5UXeLm9
aNd7n459Gpjx78K95ge0KGmitKiJFbrMB3xENq/Q+VLIaiYgEbdlU83/lC8e5vei
Wg4PPDNfo+HYUMZ3LxqK7A+y3Ua7L6vUCM+EslZGtMh3P9JXmyYcYhbmik0FTuib
3fd7lMVgQu7QvW3gUKx6gp3dlar0gu639UdHs2++e4YSElcYklffzSX1FxHR2faJ
pNrsPgOks6HA22odvjS992rF8LBSPChb5+mV5rpIuVMmjR0hZf3MN2rRE+OoXoFl
L4LaPAEIvFjfY0q08s6Zqkf5ooMuU2K29azxQPotxgdurq5bW3uYfbiHvUjJ/nqK
+dNuzPe1nEzuG+WqPj49GpCXDqeixTxJZ2KsnyCfe7TdcAsJxHLsNhCi+zy9otlG
6LxJMpS3bp9KsdlidxoT9PvZf7aCDFZUtUxHuSP7wposVgrxXXQBiVWEPvIstSDa
fELnbPv8pf2XjD+hER471cRqOAIs0qM6OLjYzspZC9DiTD0YRGp9Sw3hn7lXi872
iqvj+n1w80oLD3iIjcc/7Tygrk+t9STZi8Ir3iTHSjZs6Iej10MiGK9ISEx8oKzZ
ss4sy5HfSPsaQR15tFdoQJW6hwatKzB+S9QoprEZK0ibdhS/ecG1ZyCzxhDDFc4V
XceDC/QTjue9lkKETHRG7E/GnKkQDDOD1fa5y3wHbvY8EagULM7kQDv0Iut4IPwQ
SVEU9q0wu7zn9aW5fQ2kfLQWbdrzpUw/ZesLiBwKv0DIxRzezjGOoRU5oL4/I1om
hXrPf7tTWpn1JCqQsujB3yev6AS2Bs10MyZcOMeDVnRv71qmpWhV8dFJ0kH3/SgC
zx4pK81R7/EAHkLEfb5Von0X9NSWwW7hNnVYGni8BdijadCCUZRkkrFc2Bk4dLpI
hRZE/zdD335B2seOgufXjCyngWh4YDXLRuTdmDChBIPhUs3wcYJcLWFr4cpGL2e+
MviYC3kIaRrZ5/17+u3EcF/nfZtGQj+z7nRLejFGXzXcvDF9jvtju1rpniVGfHT8
eJnQC+tuSxPUWTtvuA442BiFYUGsIsODxgLaRqzWm0XXf26gtJdRd60fhM6lQy0p
DppJW/J8m8VXY0Y61rWd1zVIK/cKqLWAKpwEcc4lDQ2m0vL/meAZACj+I83ntWYn
6spohhufE9RrwjA1puDvzGn/tUbEfwpmeCYZpaqApgcXXk5Z54G8wiv3XpWr5SFs
oyuu/Gau+IYYHtmOdo5qGN/yznGgVXMKV03DK85ediw2wLghMZu439W9lV9iW29J
cjnslnZa/aEmm3DCQI9QpmzQY+gEk/KBT9y8R4mO/QKQGpuEddw3x9aD7u/zbFmy
8JFfW/OrkMUA5K+5a3jrogRkV1wAmgyLi+COpoErfOqlLKHL+OTWToZ70EwwRbpZ
jtMdUmZEzmkVLPofC+D1J3uk4WyzTOn+rsZ/bPi50wgFjWavfVyNuNpWjUWSOEm0
aNQOXlpS15lySAn8OKbRtWzvRYNB+FmFmYsqL6cGRZBP8RGi1ZlV5toCUffwurVJ
fgMt8r05d7PH6PFximrR6JFq3OJLUSU9VyLqNGMYnlSeq46q84aDR5R2p9yY0Xfe
TrHcZUiJ/kkV1+Ydt4BWVKYK8RS6bPSuGS49k+VkEFsjJ+ohNF2i2iMxmO9TbsqO
xVgojT3jZbdZepsokvpDqW5gUxPSzSEq1LG42iXyhtnozNHfD/+hXl/fkkN8ZT4j
mLalBnc9mz8yy6A3FmUnWeoj81e7mRGz89h6HdDre4QzYISywe1mkQZpYYhx9wUA
PJt4G8ErHArJbGqFSHd4EJu0Y7YT2rCmrtaIxp8VzakbzTwQF5b1yGw793SqXoWV
44TQDhzul3sFjrtPTaCWelefp1U6c1NtUCN8ULSCIlj/9bAt9hKH7XTczQF/U6fR
rkoHAJ/+39m+kD7bL7k9/RRfi+0Juh9TuC/X9yAEXS6synRIf6Z6tZkX6p1CuJUY
lvVirJAgj46ogYSLaI5qZ6x1VikmMgxL6AQLdFmIgP6u+apys+/nrHV7x1pw+Mgk
0ImxNm4uVMy2KdOsioW3OX4STqjOgNBNMbZF0KCm8PZ7TG/tbd0R80IiOHikbRin
eopV2thhuX9dVFPIdL4wAU6jzo8LFafr30ebqH5Pf63w4vLoj0R3VwjHv9A55GV+
JniTcksGPPurTqyPniNekvEKN1Wi17iRjOtHsBi5gelCUnHmsb/N6GwZ1XR7uCNK
wF87q8vnHacEcgjGh8fracl/puMljIfCjcrPfNiBJ/F0HntiLwAqQM5G9fUDCjoC
T64VDDca4ZIPFNjNL1KKuMxw/y/5f7rwkLALoD/gTinYobCOQwclF2pB/nC3nPhi
OGvon0K6LfzCEP6HnGuQ1WLdlKuJ4SkxjBayJMEcyI0zqdSw7r4TEPj7dNgaqJtp
bLW9iiwmHzBNKVWhT2KSZ/rDGJD6ONEbteyFedw0G2zwsK7DwzvhLKUybmfRMhd5
VllE4FditUGttqcJxgCWhC79sGUfvMMsaAzzLlTIjGNAFg+uh6C/YvnvIeQAWY/b
hKuQyENEsC6pjjtUB1FKvO7vLZdl6V+9EtTYMSi0STEtNYgFdHaippmgID/Rl/5z
rt0LgRsxFjz3mGLFIUHGsMvdkZR+7TU9R3I8MhIXTujS0usBJVYN3RKf+c5jeHLG
Kh5qfEjl7b0a7wNNolJqM84xvxsg9Ul+HsEp4l5yw1DFfxwf73Aogl9QDBEUk2d6
AlB/JcAWbzK9IRW9L60uH1zhaDLnoMQBgfawXMfFQkd8FO3elNvpehZwVPDCzFLp
zeGPyr7u9Psd5g4npoMUUf1GCpP6QvsTIt4Su95VRXl68pDyQRkMX7BSiitycjR0
MMpgsdQkoboRFjvK/5xiGTaDB1j63dS3bWeLeWN/TvTqfWQ3AkbAX/m3wzF1gEiv
vwm0EAA2Q2a2UUSeS02IkwQkLJi2ryy0Oc1U+gsYuxXPTAj/GshTFhYbx7K+JQAO
QsXVaX1tSnCJQUDuHL+VPa54JYs9U2hHbTM6bRVYiGAbXX+LFyGi7Cr93SDXEY7j
bcIS63tVeUvf+11mJzrkPw8rs0qZsrwWLQjdbxzZpmy9rbRAZFFrtPmp92FwpYBQ
ydAykTRYuoCIg9i6aGSTEYVRM8ZnqAUqmdqnACsVm46X7RzMAIQh9ffp6/ixmzsK
I9uA/jY0n+tdnnTaOHONhkodoH365zN3qArvBNHvFP49VNrVrwNhyPgHp4lDKA9T
piWMYEuKJ1BAbHsIVXO4GSp+On2qNfbZ7mm60cWH4eElSf2slCcsZ9+t5LqyMONe
eEamHz9RM3Evkgy3jy8ayO0i9wkR/hxkj+S9Awjp0nHLzAUsJKLyTDJJqJD4+DMk
xpYieeMIHSyLgYZvEIRjWY7zYYVcpcieQlCRBzODZrU5XxmyfVsa/EmQ/9wDOaqc
LcShld9PVckFtur3vWFuCmjWfmeWWy5Lee2o0ahsXCytF1ZnpUTrGhM8WvhWTHig
3FB6ufqxyXWy6OcCqysFS9KkLbvkbuPQsKbYzLLYYgi8R6+Gra+SAT0wBp1tat3k
sqvqyGK6dM+d8ywwuObWUIILUeURWtZgacoZOfhShxFPCGB7E6iXfV1Q4aS6vr6A
SVtZ9QvkiggskR+7CqpK2nFqhM+gqM6cdZGGqj8jR7JIovUg4cTX+npNaKAsn2x+
7FU5eX5IqHOYOomhiSQXSF3RQP1T6ggI5fzFNYLdDZ106cgbFOHKRkXc0YnntjJc
g7w/yRCWkSV2iHJ4akelF6LzWMLUFKrjtMw6OlUKYPGbsJn3LzYkwG6cINPi7DvP
/31cbaRuQoBTzlewmgLSb10OeARtr4X3YYj9i7iJU80HWJAW201Wace/hEiRzAgG
f1hI5BXNfAOPJCmdNB/s8Z/RapN2bjeO6op7Xue/e191KpcuocdvRquVHwVH1PtV
iSxymZu4aFKInixmuy7UtHW2VJhfZuLR4CMstBwXCCifpHFtx7Cw+pfiJ6h/jRZF
QptSB9eV3rgdQ1e8I95paJ9/N9xuLyT11f36NT/JTWDPurdKy4KI/3XnUpimZLKg
qIWhdbdozqxF4GdXJE+kqfwfFhkSHjx0yDzHmnaylL4BSHk+aFrw0wH1yAVoQWAd
GB5Kx2LmDjBydBP32iH5wW/AN9QiB1zZbcJ7I4kMzGi0LSwyKR3lJaxQqaegQPAF
jdmwTW9IqMZOWrqCtgyGrjtaJNRtrCH/xxe9vJ3/zalEUd7euh8GpVWPTR0AS3L+
WySk9usxoA4P++v0RwbNQTFRbMYZ8d+9bWUXqIatHQk7ngrhcsFwIegWitTjZe0N
ruye0bkvopHk2TZAEsa5C+ZmzKWXmIaz/dKSd/QbQu8tdMo1MYkDJ77Y33Ct3VVv
1XoniyU7+YiCm4Gi7VtT83SkY7V4XxCyiU2MiBAqAbCiiuUsEBVozorBj+H/5Jtt
84BCfoOXDU2lmFQHBDTSmlUJZKTjYVmm7/c+RGx6APqws1kzKjoql9Xs0jCqt/MD
4Fh0kxaqCSLgZDgG3FSYbZQVDRxPctlYuGt45lgU06vblL4sDOWkvD3o1PgI4jWA
X6cTE/UgHzv0wwtROU/kTwhhd0SoffKelovSCcVYWsUGAx06AyYzgsEMQEIfrWxO
lBlduPrwh8vsBp8FQGZSCD8ns1X27KMP2Z59xtW0GAMXzsXn5UU/Prhmcf9ASzHr
ZTesgJJX7yBsfcO3sYjZPkA1Vp7qfprxaY039eGMzkdgOz8TaJNjdpvv9u33qjrd
OMJOqLJsjke4Oa7Ipr+8qZSKy2qCjLrpds01Pf0lkzEuJJU3JrrAupm+SbOb+dIf
Gla6tfGmC0+WHpnzFUFw04XdCTeGDscBsc6qjLAuFTZCqIIXt+wfujDgfHInrO1T
RSxnoMZWGLhBwmfSF107bzMeUf9Jke1LGDcrm2JoLj/pD5aVf9eFG3dzIQ6eFjtQ
EwabLaAeXv9QOhSaxB9W+od3RCNvzjFgJLuhxe6kfZhtJGDFJ9y6uKTfpxZVE7We
6bh53e1sbapvGe4aI8W85wFxjXf78lBaNWOJnDcIVm/LIjSQBF/fmhJkduBk2xiw
uYxgqje2Al1+IsyvX2OimtL3VQ2Km63DIJ1/fyqQzW32E0lVTRtRIJyd18q1aIw/
v4orNoo0hTOKrI6LQ3RVdrBBVhMWw3FWSpBvyo31xyC68h7O2Qq+oG5KYHGhjNDo
ncRRQ7xQbd+MXTCaL7T65GWaW4gVEep+LFft1EtU3+ro+jmpK/+0gRJyx5ANPyUt
3wIq7XNFShBrgUi37Hnfj5hDc+SAjtJWy2AYagUZX8a/y9950DQguN+Dp2jFecK/
8yCuj9KMk+3gkoVrsbwfDrlRXp9PZmRZgoWIwbufnoEU4j/uo5l6OS4AFHiefYCz
m6NKDi+9iZj3qJRoaAfYznNkbIBFt7MwhgGFLZXD/wEbhie6/WJ+D4cuAo7SMXTU
yBLwdznxNVJfRLqHs3j4fO5LmAkkZDnFdHVZ7oWTFQelQ/SVnDPMRWNWfrJTXPi0
UHZCkyAwjl1soJtJlpQXFYFxXtb05s7kfvbFAjwC/Mt3G8ykoXjDHTu08G2L9Nek
/9abztNGp/ldeIK+w+6VnTpoQJdNTLktO4s9gS9d9855XIARz4aox85TboRipPWL
LtLPCgqxGWMDCTirLq9Q2xq+2qXJ6pTHTmI0T3TIdsLKu5abess6y4QnCyz4uk+h
RBZMbTbq8URUJnUXQdbOwX0X+Z9Yn5PnUVISSZUEEXxqXd9mv+U/xDtTs+KKrfzG
1oMNJ1kqf71/zNi1bK731VtwXPzscu4EMGJx+TfDSofqGqa0r/p6vY7Jro0bV4Ls
LKf59tquGdUOff6gXHNbQ6GcgWutUtF0IC/4lCuZMaXFPFgXIiJ0XGY6Z9J4EES1
G2hqXTr0LQ+01P4cVHpqKa58gccINcqpSJ5GSxcKlo2HrA5OMPomWzQi+aXU3vMx
kclwAfzMVt9LCJ61tH6lXyD98PVCJfa8k8ymXVQentkehB7ZONCx8wHlv0l031Im
zANlChFp/Hv5tADba03DFlmOphQpUqpM8aUzjAgQLQzIixCJM3aPEo/UGUzU50ZP
LdemXrMWGNKdYNgTy+BAJOkeHOfEzxlmW8FRER+KEU43iUAKEOjFt1IAhnBLkk2z
kkTr7pAoE5cB3TQMQOKrFrEMvDGuvOTNS1B83HWX+rRVgfndG6fJHWnavhGjwKey
ogIEr5rIu5InndXvtrFpAGm8BCaI3ppnBfqstC5f9SPP8h69rSbncUEbh5LEjCH9
G37whRRU91rTjgmUlRLT4L+kMoBKYx5PJ8QSsRpPFHGJ4mnjI8scZSuir903YH1x
iFD04f3AfcL14FpPbtXxPBjrc9oA/+x3nUS+BdJUJdBuj8/CrUUMY7UVCfGr20eQ
1vYukaX4rOaJDXY140dwA2wTrZK/vzrO9wPTkI+2/HANNh08qH8Q4QWzNMUSCXhq
ESUzxwxUNAjuYwmNwZhqSkvdJm/wY//yUMobKmcTkrLhBQTvy/PIc388fP/+JFGT
QKDd6HAb/DjmMiXuE5llCnV1kdrHljDx29e8aXh8qHje7S+Maq8jk8i5PlmXkWp+
sHVbbpaonKuFSIFTQwVqpPt5QZFE+qfdajqu5S80M89r6YsYsMPaoIWhdNgIkE08
CfmO0Arn4MamebL8BXoqHdg2t1ZpyzzXwlCnGXBOgzD8OaiWGT7udKe6rAAxGt8h
tYXFzrC2wLqCBU41p6J3u3v1QIlxaRikvHols5EZX5rpIMnEjF9EPmAVzAWn9veJ
/WoWANW/Yn0jqDy0ubNqtHFXPy974qe4P8Iod0q/fK5ZfkYUh/673eRzhWw/AeSL
QLhhKPcQzKFO/qvQ1GwKMkYfA4vPU99bfOCEKXW6xKTXwPoHuoqxUAuPXkidXqB7
8hu/8jYXrYFpLQ3Kp96FXa4g7e8GKE3G+UXX2YONyEDaA6anKjK+TjoQyuSvKSCA
vVRw9OcJjOYNM6N7gx4A1xAVQqqkKfzwPC5F/gpdePJDLv2mhoKAl+FKlcABWoas
92yU3hxOmOsZzUZG0Y3OyCjNe6KU9oSdnF0ScYnbUud97l5z2pMFlhrVmzi2dtE9
RjaSg7tuWPdsVV0jeC7DA+jpFrN4Qv8ginmGULXwKE1kyeuDoKaKA2BeCjVW0wH4
2uJ/LQ+JPJ9Yy62e7ACRbyXG96h6Xj84LkEqK6K9o7x/72XY/rqkNnzDXroTeMTa
HqjPGSiqnFuvlEgz63xrlS9Co1Jyy6qCWvgIkg0c1fvIHWzCi28L6zAGY37QVFLi
q2tbRx8giYrfMjkCE2REj+xNO13vVchATp125Kz9F3rblePuEzQm73MI4F13qTu9
hFty05+dtNdSHWWY3l1an7jDCDLVC25j5Fh9fVXcLwhzOGlTKrjnxjaOyEvTjMEA
IXGimxBtxF92OIl07tQetV7lvJsPF8hqAvH55TFVeJGfSHEgua1lmgbjiBbofxtK
NkvuD+6DTz45eCf/+Ua3qWDguwrZ/gaXotZNYUSoHNeZmMUgCshZbD1C/QfEslKM
O8Qi6i7xT9QBjJ9La608zcV/KK5IAgfxW74I+wFbQQO50l7R6cDa2fk6ktgBnr2C
miB1UGmhknWTLQmEd5zEKKoniN/SC99Ak0YE9i12pBOzpTwwL5/iD/2UotjdJYeM
NB7DlPlJeJBj8UK/l8tI5dQTEgxuKRqFbn6MXe5rIz9Us0hZHiduz2bIHHN9a8/N
K26NhuQ+ZlqeiEjn8jxmXgrXGi5NgYj46mPKmrTPnenptxtqzkRhwod+BdEt60YJ
A/A+WuexRsqdmUqTYq2tMqHnfaX0TNmvdjPCvNFU6+iH/wiXWNNC4ELcUwTlLcDp
MRLDCYVv8/IplLFMOVEf+ZIaUo3w/6aQ+6OHb9D8hHqUdCQrbECvNiExRLh+oqGx
qc2M2vbIh+5bTKpGGSHrY2Fl7Y6E9o5rZSHl8c1cdg/scKKSo9BqeUUxmpxVk3wZ
CpZPppEJarrnherRjrN2Ov3KIZLOuYrvcS+UMDK/5dam71HwECKMC6ABrvgx2k7s
MdzGLqrY9xx1mtchua6c6WzNMFloYOZI2kLa9MBWQmc4k8mgHpTh3GMVgOfp/d14
N7z1jInDlQ+sFH2WsCHsWPNcww4eJXI8DoIcj3g4z9DMOd6zSq+9c1/Y9F4nMCtN
Ln/Nv3WAoQS4+L/QPNpi/1eCau7Rj5TGdu7IkJ1jjrAqI4V9KlKfnH0A8ix8W5tH
uLT0ebYSyveYEdUVfOU26cw1U3aoOZXPTzrYiUaSnyR/ox679tK7F+c6NWa0s2xw
BiZTa/Y6duuMq3Wz5/0T2GXQSwLI1HDUT7+1qpBercDrlYCucXnSEGYNXCkQkUUJ
XcvZ7MGf7/VpuvrkHl8Bit4xGwZFxN8oSAg6GOhw4T31sYBBeIlTaPr8OoZbD57Z
qxUfsIoii+aCZcO5afUa3l/1JSJ+RsbQV7aOctQ+cZ1hJex15JpP3O1LO3anB+WA
an4rymPdbaXdCoREi2uAeobhfCPI1IKzAQ+fQ1XRyHlf9EKkAdhkz4EdQ2Tqii3Y
bbSTjh9n7JDo3QdJf57c9aZwNXedjqDHZrb2jay/wPNrJjL8jE579RePUacE4bJu
LETBfnSLcxqcgXngGXqdAFkGm4MXsU36ZNVDG//SBglaKJuGjrPfXLoRnwaEqbxj
4OC5gqsKwKLdQ5b+pPZFt039Znq5Ilxt67ZuB0v9ECbYpz8aTD0+XBWW57Cp/+/j
JTZmoVHzAEMeCyhHyoMuViL8vCp/vXhUcw8elh8TiKmV+dxp24ZKJQtPxPLAR0+X
B5ygXknvCG5krqdXxZoqasyQh7kfbjFpHlnU1UixLu3we5ozU+gynYt+Sq1ms3Bs
AGzmSa4psE6MwpFXlIsn5cg90IgsQ1ZiVtnTkMqGubVeHj/YhiGYYTN7yoX0tyWU
hEPnOT3Vw3LMqedJyhamxSSAqvxJOEbH6o7KmPAww02T3czoxdQKMOgdJ4ejdo7G
5bcRIK+2mDK22PlkYnu3v/1CviQfzo1mUUyspQaKVp+Legj1otF4u/UOoPIT3oSs
rbuxrGszVH+JHWy0O7Oj9pRgs6SelUsZnBvig/bX+y2JnHrobxAVzQfyEDmTo2Jt
dsFCHftjF5WS46a2v2t2iktio4PpcgO4hfxTILioMqWAopXWdXiI5OmYd/8RVXn4
TvPCKsBJ0hIo4YKYQHkFaIji9kxqAlY7oAM1hVa7na92LwH1MCJhXgBRzKqDb540
EcRTcwBf9n95ctNgIMDMSL5Y2RB3z90kIUqf+kREk7D+Tc6X2Z64yHoGnqnUq7WP
rCSTFemCOykYrJNHXzhIn8CvXF0ncsW0/FmkZ91mIZyKSpZTPOhJrGtNd9R/TVZM
hWk4+/jVGCKCFlXlHp/uiZa7zzYHS9UBUkYGpX4aWVMdjniDfQQQaLAQeyFTLw4f
QntJY2853b4+SfKNadfeNWUN7ofQE6zDkn+56NjDfIo6bOiHJNT2O2mhzOIA9oGC
sbRqWH94/iR8MVOcddeHNQvePjiY8nnEqUDAloNcuXawHU5cl7N7l18m0UwemMqc
sUeoEK3xEo5cXXPyuMgHZDzeKxNngQZ6AfrpeuaRYjgN4tfzRkRqXW8lmx4Ua/LK
evU06+183iSXCkhLMbs9v8skyx69AnGhQYBprEvJW0LaJsAxvHj9ZnjUqwd32JCB
kFjgL+UCigeOV9OapSjyjQgjCdcFwmXSEI8pdC4viIf4f9rrxFCyKEYVx2221Pj4
FwP8QoN6jtQjez2fAGDVp5T078s+khp+0MvevrATvbx+Lehg3PvEvjEvMUe+GekB
VZef87x6/Dr2PLIsZCPsrLfUvihBl7pp+ltnjcZKorgwNXHE4T/qG747CmaUJmRV
1Q7zZJpTBIF1Vy2Ao/KdtnLboYUc/ckBDOrh4hLtsK7Sb71Vl1NQB4xOSUx5AWL4
zB88WeDxhv4MoYvWNfPhk9IoYnJnuKv6g5OCVMgdZ4rSnQGKIcVQr6dOSHjQDW72
+gjroC66DeIoTVJqUuxefthoDXute/2zfwksbj0YU/i0n9VwDhywXWuq3//0wBLP
QIxEHDNcqBLNoD2DInH5cIAAT5TdVCFXlkNDGT35YfeRgeEpiT9vCUMpeYvDtRDw
9MtlIOXvFOz7PV4TFs5imOKVOAghSyX2ZCRFp909d6PcNKd32m/LDNPExqBC7Zw0
Yw2tjC5DUbiFjMRgLdT0VmDsRa7ttyBDu8TIUrfOZmMCE+fBvkG8td++SuJt9MPv
aPvPGEqZxMLFm9Kreue+ut+6AvMlF984WvJYoLU1eY6N83EHS91i0B/jcLPtH7qV
DefJyzQU0BuiSsmuaDXD5sBCjfcoihXHsmgjeoMZyRSydrv1Glle9ZBFYh3Q27lR
L1O0Pml3Db/T6UJtn0CrCd/UCaDvy7h2H+DFeNxlpYZL2Tt+OEz4mq3YgzH8vQ8z
sZm75CvGQhY6hnu3M+QyCKVZQxH46tR4wyzbfifZm81xIBkX1W6KZKr7qZygnyn9
BolYCSLskAN6E5Y+ygAAvbxCmKaAgMzKUFAug9D85nsmrpFkVPxZNog75pf1WHY+
+wGJF4X7S82oVqZ3xZmk5OEXSdlXxALI5lr3ID+SEyo7cquDU5T1H6LCK6xW1Tyl
dPQbBr+MlB5u5LWVmeKyZ0wsK6if5EvJvgC3VvjIKIE6kyD3c2BC9V6AKnBzOQTZ
btMUuVYHN2ATJHLinIELegYAzQdYAwsg+l2yvk0CGjZPuTk0k0Sl53KiGH4a9EkU
cH5CBRfXn/iyBH9qPYoeObwQhbsTWhVcRTF6/hpNXoTFmBrER2XiRIlZnh3EgVmO
woqQ4soafYDrk2ucTf0F+ssfqlqY/RRfeuThMT8Ta+6kttWYB5/PObt0aKWzqdFE
iyfGQjmbDvOpFcWcJfaFWJptDLHigOe4REMf52iU/TNLL/SaM6BFOFwLfNZQtd2N
HF7/ZzMhC8tVn3VrgdREp6+D4aOyYX/ivmzz6iM1/tFn7NJl7oRH1DJoBERc8zDB
CT21IJ9jKOpP5aEbs2qCfkY33JvPMASLdkVFDyYOrH+b4iMLZFJcWCYtx6G/7IGF
oGu5gByqBpm4vt4uT3yhpEpB/XnpxQyxmjwte0FDUHh0BqUmQtu4pPSlfTfdGdgp
aocP/OdNx84x9kGIDTDFiVHzoXsoxHxJkHQpkYgwDdcWPBzRt+QJbP+7lBmCstBU
feHfRFFtvN+OGpLOkf7rxmGC9EbQG00lSzKEiZk1ZmGijWoHFC/ASfga1zsWR6yr
5Vtqi4hYPinlSTucZ7TY52pQUYAmGmGVE4K92YAlJ6rsR5Gm7Yd55wsczItm4x4K
qbULQzpPEz/F9+dHAV2Q/0rciALOPZaQ80ag2HNKqu9vYfpPo5+++wYVlSy/yEJr
wrT0+nUn5CFlAJdN117fwnQm9H6sLzN0UCndw8aLuXoMWwBWKpXTjtG/jDaeD9XJ
Bqqvy+B+YHDJxA9qVwNi0wg2A+oUIVSOFF5/dBTtnWx8UD/bQGu5CIbjwwClW9zw
THMVAWlVSkA8iRPSJlHI8yS51M+MHgOMPbxwCGh+jrGJt1GK4sG9tHIiR/NJnzzH
FvAPqd4f3DjkrQREKrVv3TkCc8iEdQBlTqeGzkTW7jhZeXHYA8/AXWZBXSQ9PdQr
4sEG2F/lrarbWvf8jEB3Yqz5hJSYXEOF+LpHru+P90QsyB25EJCJm+MMpj29mF9p
6bEVvoHnY7K9Lx4wMTpTzpzbgZUDbZ0U7TtsjstB6awlmM6xqEg975zJ5GWM9gaO
0YQxagN73sYIjkv2Kvwda3J+H6y3nKWNkFh/pZk80B5TeYavX9m5Q1Nc8h+faVnP
V/fxJQa0+nzBByKv+qGE0xKuRlaORkkN8WxYDT4LnteSMRFn2TXTTPtVZ4KwmMop
1MIrj47Xt4GN0cK8JyF/xm3/gmhseSr+8p5q+akvEaMeWnu5XlppIv+93mc/6dz2
t7ds73jD0zGP2icntOerbQOUS+/o/YtxMRc9ujJH0DhgN8Y1RpI6GRq8As1rhP23
8bfoX6AtwqQqOtXYafzqpJsBIF3kX6un4lxucX4P+0NrwWWjtaQgnY1pZyVIlSqb
Tf64ShgcIBUENGpKvqCIWFhje0mNWJEbcoDt+61I6Msai2WC2dekAaU/QNcStqzh
J/ZoUVB+3ydH8DN51xr5C5vba7WD0sbINBtKjH7p/INP+wNlIrYVy+5G4HUwe44M
e3nt1jLNUk59pnxkHG9LMW/N+lx3HmiOw5f9kR0/7+2U3twg/uCE87rO4wBOVLOP
3fhcVDvUEC3wHSlOoddiiVRnk3RlSwQwGgcAJVb3k3ue7x4E9SSfSFW9n/JqHm2/
0gV3WzNKDO4iDnQPr4Xh/+Rbu/3o7dRwiTmo4K7wTEWQ/MvML76WH3dpv9FQ0fjX
/Sgfi5AGt+swKL9k4tD3+Pe3Da2Z8cetx9RYUghjA5Gk8mXIZTIfZOKqBjhimxIZ
trQXawvAKRLt0oeo8BczdCYK0yhLipVz5g3Cw8xhfm+FtFQK3gLISFVi77ZCiNUl
nhoqXmMgOPZ49KLwv+ZocqE39qMwB8Noq/QY3nP0S48tCWDNeGhCEif4jMW+tkjm
g4BWK5on8ioTwvGd/G4iv7xSvPeNmsRnffC/+yPd5Z16qfXfuRxzfl4wWKUnznC4
6+91D1wpJq00SFAP1gZj/JcKlmijE95FndgnM+w/dcLe0f+9VktVoIijKcFExb2m
G0rk5k/aLnFy2gJpjdvuEk742JEfdeVdBiZpCiAK2osNdMoVDWqFZoRXsqgJ4jA0
ZYO/CAFMFeFPaW8HC6H/hTD+q4MQD3S/rEVY54kRNFmmO+K7MUpeno7oocecLU/s
LsNH16y5K7Bg3+oFoM7La4YONAmNaVQzxNjcue9yCwCxOVawZsm9DQVpc/oxMjJk
SFblN0Num+z0QjJkFutFbWxu10FlIP6c+cENrxdPevdHZbMIWxR5GsXEhBhim0Ms
c1W8Ud7XS90BTtB0P4gssUx4x8h0ifh+j5hEiSZlvctL+4Ys/HcAfNDOjGRBdmE8
7Jjy50hi4/BVD9F5f62fkbXwigu8uZPteWoZlg4ff2vfGzvM14ksxb0l6reUbm6W
uo0aBZNcdvPG9UpT4RJYbWgrRJvRRLXOboZ+Eaavepwx42KLueb3XqHGCMkarI7e
jIblzru9C3ZV8ycOJ0p5/+QnIMVZCnZDf0lZJeTKThklBMwWl3X6+11w1ZALOuXi
1p1Dfyx+Z3WYLmIpNxSfe+n1mLOZajqaMGx208NilPSt4ICom8Aj+35XVVZYJREY
EiczVLQp5A9Fkh97x4ygj7nd7Ch31R/iTuz0CGc7wO6Ib+bCwOIc5g5yCFMG4jIf
rBYWJVLhYC/7wAeoUbIt7l9XqXqbTZ2X8isasATMuOnImxdOE93QJD4rEkK6w8Sa
XLlljNVRpoBIeGdLdjyELeP+hl5aU00px/LsKN1Ifm6f+Q0IufK9NJ7t7QC8frU1
rm+XB7jq/70RBTCTzqDJua1fMkrCB3O0VaR2jQR634ZXctdcTNA0KuO1WwQIObJb
Gc859xRXNiLwA8CXoCUwixfTZ7Gjn+vvKcucQTGOBTQe5+oBDHQ3wRIwQSfWc+IF
znxVihB2T5D7/CQCmuiubVYF2fPspBnl2KiW2afUv/de+gdz0HJtbKpxMAroNhlt
jh6PMJeUmpKd1g3L0+3EohUT5J/4+t+Hurs8QJ0Buvvp2wLuiBNO65oo2YV3GAJQ
MsV8qHY3bX+C/J2KS0uHnpd5yGO4qWSw6CqYFL9yndJG0NRudshmiIFgWpjKTfSF
WNyK3TsLvwTS0Y0ZMtRL789jl6ebGOpPSjknE7ACJduJ08qxU1w/6rXax5YJNiCw
3RSIrA2MHjNoI51W3LVhuNz085KSf+xrR852p4KjlDC2rEIgUS47vbTUFjWXVlQA
7svSPLEYO4ZKIlo04sBmeU7ccASUKBFbvtHVzHkqRLq0rVWU4R7LxwDLfJL2YNow
03fijBX8bxP5ve1ItosvSdYDOdczpSUSVlP4ptU0RMvii53ptdLeqfx0tJ1JUWJa
UfLTY7ldBPvjXFItJ0y3ifzraSE28AvixC4xGOTtNlODfpqIjB8CkuB4ZkyU15Of
c83VF+ltw6G1JF+npLXLpctbDdVvC/ChIssfSuZVBhNAp8rc3JyIFvDjugrtuN1P
z/2cIPZFyz+gpuK8z/ZTBtrAvWR1jm61KsJIPwh9Ng1dg6pC1WuEFkrObexMDrFG
NKGVp9z9ltI/gm8fE42YTO5CWaPNQZikdZWts8q0m028OM74z3fSWuKgSrj2cavy
A8U1weWAauqLq6AMUAj/f/p+QQ7LAYdlOWiJyLetLiGWtBitSDRugf2ytGmbHVpM
ZDBV1ULOy9JeM+Z7QXO7MXJYs3j2H5bDA2/OmlOk2wNn3u2mV09BJRl4Nm52vvpT
72e8GBpEZTuTc8dlP8UOUht/4BUZ9YqctrFQUbgClv/X1MlvVMtRou+WOY4EYkD7
UkhrFeNqjo6W+Qc5ish8cSIrxGwdU03spW4/pjMs0Nh19ye4IsyxS/DscGxZSRCT
jTp+WF9G8eNmq915VE2gLJU7TTN9ahGnE5aha5r0QFt6ADWjMEChoQRm5giNlsju
hH8TcVy7gE0cXfpDox9WnNggRKAK2iJ5zmgmI48vlMNB0EIN4R79jVzfoBDLhhf2
+f5VaHolyOq9UgxBV7M3ZM2n4Nhil9CKxygqRayZzzeuFO/AYUy422XYYvO0X/aB
RZd97PsGdvyxKrDebI9btQ+LIivroUDocnEsSNgtzISotQsxUSFqdd0ZxtA4Jwot
rXsF4D9gVuvciIe6mEhdwanmomFmqKYV1ha/eOObk5R1nLaj5U94e2bT0iseRRlQ
/MzSHOZ7Rl586dfUKoidgMj2KE9Hc6eiitfdI/GY7QuTnAyon9dtWgQhWeRm1Evf
EYFX0SmdIwMQFHrGlOQIF36ESQoitEi5eL5It9xTknuD8kto7+azcXMU1ceO+1Ol
v8RVVWJZAMz2Jfe2nm00/ixPIe334rj1KlAvqvzd1VS568yiUr23925A7eHaxrVf
d2k35YYKTUELiQNIv8FAYTq3DpQ578UnxwjqLfl05BmiYLY97G0DGiG2Fgyc8OdU
Z8L17Od2wD0h6maAEU5oOT3cfY35q2aRgsBwMZA6kiGKg57Mh/MbZlfcGJqReQQR
kfCoXhz2J2cdzFY0MhBLYdWEgfQoTB1WkoutyN1+O0DZ2ncVKQ77Oov+d8DkGl7U
/sGZfdRqYnrVIMsE/2MCir5pQrj0RfAn81MGSfT8nEIPjq5+PWOcUQLUPqdEhRod
fWU+vZQxuwTuIg6dikilBWxQE9kCN6Sovdc9xx2sn1Azwg9U2qqChKktIBfngARl
YrUUfhTABl3uzU9omQbqMxzXoDCH4zlB0XDH1eGo0CeEV64xQ+EAki6qYQpKsMzR
voIf4I30yZGQUkBzBYq+ppfjcP8t6aB8XsP2kxr+THwsL3+1WaQeg3slgeacWMlP
5huGHQrzmLIMWO/L/VcVldZ1uoBihWYNYKWfzfaR1xiI+xIfCEngpD6HCQMRojWW
aOG6pfWb4VM2Fxd/Tn+OvpqpttBQbISCODrDb9oaCeDEzKVQXCo5ROG3VHkwpFAB
/8iC6cb5Co+o4mqC6cDSGPGhX9h38LM4pjtqKvHQ+ueNuy0KDXzGD2FV5O484jFR
09iYV9q/egZKCR8NRrHJa5FRFoIErHivkJOCqXDSb1bDYyVlnBUf9MIlVHlVsCc6
iM/YGfSjAbEtUqIH1WtGCcFR0Ff+NjIN7jO3A6iTruNqJ+jZQ6Jk10WwR5w7f5nr
Rc2S4YZLusmRvgRBIf1GskQNZ3kGgeNhUxis1EPvsfeyQrsb+qr3Mj5FyvD9rUcM
xPkukXTu5mwXHQSMc/FCd5YEB67U8mMXbXnEhXemnRL58Jp9RfXI/JFN7ZaejMOJ
6tgJ0gdNcylG5qO/EucJzI3EnLgcPYCQIaUPknfl7wQAWTilK1CUxvRupNUTyxvt
pLtThpPFV71wUGL5/ajetzcfhEFjcK6z6TFBSVb5ZJTYZ3i7xXZpacm9cWZQIe5r
kDtYJzXTRjceC87Jlu4z+NkZRgfJ07rCitubzFRnYc6Be0+pktoiMJDu66wvP3E7
5HrUPVCSctQf2lD5I5+QQcnVbxVJVV5QOoqo7enDMjMncrvyT2jVW4KxrHuz6Ppr
HH/wyqcdUaj1J/kCS3ovQ2KMiEmU4muzvoaIcESfS5lsnM1hhbhemYhtGuAXzfnP
ze49rN/tkqeN46+LB/+lTGLrSfqcOWlff//wLdSs/HKZFE70BiCYlXTHG1hIBrca
9S5nxCGIZCHZV3L3d5RGIMNh66GBqsV3VfpE4RuC1n7pjcZ/Utw5MasmjyKoSDfR
MRhcuhADbDrV80/vt3bZf78xF8sfTySHQlL/gW1nBr2e5RFBgGIN1qRiM5/2e67o
/+qFHrD44f3c0G6VQhORgOWVHjAnTIf8RyRFpc7gRbMFr+FkB5uKJbRcHxLq2bi9
sYkSQt9dXfMszI/Wo15JQGzohMM2gBY5GSOqsd3Qa68wpPGccHR7f89m4mCQgLx/
2/6iVUbDKzXlzTE7ZYUJ/YqjtyZ+PeEKMWv9WXVtiihoSlbmb23BSYBYmtJ2FyIq
FX3kIEx00Z7xracn/4QBKazlHV1b1b3eQRGft5YfL8AstUrRgYQwhlEVPeZpDJ4F
MrzASrtwujJ6ri/A7nuZ7ZfwFjQwDfPwn+9c0VOnMTBAgVogJ7UoRWdLYLmQx249
7kdvBK8jDWYj8Xkx+I6wsS8VP26Z6VBfo1R6ItJX55nl/muXIm7+a10WtKvFnGTQ
1WzSHOOWPnuSVRRzqnnCM+AvXjBUgDTJ4bFiQ/BJ9CE5fjlOD0HTDM6VbUC8ATcy
M35nVWFDmULQrsOUeOIwdwhaGzw4wY+uMulpqXVjHwg2h2S8tjl3TQiXJTU12CX/
Ao8WbUKESKhpzFI3P7dOzVropTyv+Gk0puMXJ9xzKHVLCcbyGfid03LcNuGGPhlt
HKttoD6XANM5C8YXiPLCUini/HSrAuu8ir5S2pMOdKyaLumKt8r2oQha3q1rmfl7
9aOWewwdq9wv1yn1Zrj1tWMAKqe1KqXHKcpoUzqFuPExwy3zELyaCFYAgTiYwaDz
0/y4JWJZt6qdIVT53TZuo4kS8F0PVRxGsuUQNsOIgw8IzTwneGgoC1U11/dX0ZfT
KZBR843fMUyBnXKFjye8HMs8cMk2ABii7R3i8WZ+S+Mnukywa5UXpKBVKRm6/pHg
ZMA0qSZojHx0ruLkSSGSwfVJNLqCJ84YNgLYz80/ZsfDHzTenvyq4EsRgbKm7duC
LuSzTpFL+fTUqIqWXVMQQMenjDYTJdn2BlZ7rAEFQgCvh4pNndiGDXtF1i12r4BC
0eeTUJed0n+zPyf6ClyOO/D6OWITfJrHlNoiAGCDXEyXJohsjqpJcuSVL24uaNeg
anYyuRNhqK9E3wc7Vv4A04rjTEmpdGyq18fTdx5OQL6Z6+4qs+ZQWhntF7X40nwl
xSEgfko6MWnd09UdPcwAdJZdLjhCuVsGBTCuirZzX16Rd0kYnr6retUnpQmgmnO2
Q9jRO1bSbDb6gM6s6nEadrJi51ofhS8H8uWkozNKg+brtdp6WmNvrwZUYiF0iTMV
y1zo7iZ2PWMtZ5a9hYbpZ1GzmtSuYI4zJNs12LKobL45FuZw6YYW5YIs9D6uWXHr
vDDpVAalzH/rznXmwVBO0/JJD9kGmSWcSHOJGN3lKT4JCBK99o31KLws8UdDNfSK
YcXdPiv6cf/jCulP+1zuhOgtZd5Ici+3ip03C1OzwGkSaR2Qfgi+FTiN3FfF/SGn
UuTT/+NeDH390TEFkmzUk8GNYpa+2CWyrInbVAwoMIJfXhgdY7rPui8O2Ez9Nc6q
5BiYtBzDV5C9MN6+yiH+nL+FgK4nA9wwELLwE3cAs9rTz/6OgDF6GJN8EE/1LE0J
lsakxFPjxzDpAfJTEPzKTKljDOFgHugLynGeGGZVjAuBnqUl8KmHN7ZJsWBMzl5O
Jn3IRbTpV5Zz+uq5D3KbNppJWHO/oBI3FVsqKHiVUox7OajI2+Wh+B7iR/DOnKv7
j77rHm7caKwSLSYjJjY1Hao+lHh8M3tbUOehl/WOa5YizkpnESWJUL8qKimqlFFs
4svxjPJMssnBFBY3A0tFs85RXdu+u2aMvPC6MjkT8God31kze7KpzGvdzEiDNEq2
RxuaGSVYRDzv4BGhBosR70Z1yKvUmxEuk6Mc8o/sHwMmvlLhejRECNFB2xLDy1Kv
h1yEdG++GCv/nUDjGeSBv2sPY7qPFzMsO6+wLa+vNxFAqMOcstmTjQw0VKzDzl+Y
83gOHi/QLFaoO3fn9EjmAYIL8XXF3EmJdPVDKKD8aSawLHnj7aIB7NbB2muTosce
qqLfS0hlpTrV3EX3LUCsTxNS077QMYYc1RZxiRj61N6gsAmAZflQiWb39BA0VJLS
Ya0NgSZIeT4rc9pcFq0eN1U/1i1iOv75N62AR0e7Zh7y6uK0DowiFhphG0zmXQg0
vKJvM92K6w66sLoAf0bSRtrPRugbjMkrxMJR8MAeEt/+tx6hgtVO8Fn6dmld8Vr6
yzmGbbFF/FI9ds8MaVNWX+80a/aHgh7tIVYNlEas5FepSKt/pnnloxtZDudmF3Fa
vCw8RpZQnjk3IGCMm2poMq4bTHL0Cupgg8qboq3zlIc725hyo1IR+bK6JWZNlA+v
MoATdQvSoItRi17fS55v3QFIDrQyThyBCYuFe30BdZA2yhDkyu1nudz69Dfq8aFb
tVnnuCknF4QJ6VE3uHLwhek61K4S1IFqRyV07jKsB088/crJ2urRagHeyU+pobzr
iVh82a108OVOS16GNFToORJI6tHIXdt+DsryRcKF+9+TWy65OwRWFLxomHa7dBC7
dbnjedIarFJWz5eM+kRO9H9pKuQyfG9FGPlwnDChJPf+K3yBZE91Z0r7p1KvZBJw
sihec4XkghsodWCXL6+il4V+MbvBHSPNLgzrSpFyYaJXCfIy2ZLIR1SSWi0r5hEg
C453iZ8y/dzEd2IlcA7UqZdCiPCRR2PhcwdWi7gWQGXbGLnJfd+60QKikDamBIex
JSdj8KyZhXgXKIG3qncJic66ygYScb76hqg/gN9PmR2YcRCqAwe6u+4uZHbSKjU0
j2SONr4Z06i+DAcxXyPJhC+FgTEX91SI1w4ev8MgqEtnB6fxJzENC0ET72nJn1hV
vie6NfH4ot89RCN0791Ph5uPDJOELqCMPTFArcEC+e1WzgV+LzCnuDejzPpDqXxf
O7MYJu8zYtu4AfCSnsxssQ1LYNLtk3f5+4amPUcP6BV/UygonOUJgAnOW4KkQfXZ
SoFBbwg8BspGyNHkmJYxbpBsFepjsWVTm8N456VHlug7Kyc7OzGtNzFKvb+OF3aI
w2uUAUvUk1BGY6risUgKZjctKi5p3tNXaOawNfNwtu0PchLGKGpgcsZ5B5e7pSno
T29BWiynDtnez2KUGdu/AUCwPNZHqxkhxzTihigYvaE7jkvmEJbdLSzROH7pvAkT
dh/OONTSm+B5NXtk2OcOUCwSsPvo9BtohFR4jgPfaHpATzroznu4x/QK+426Nl4E
v7FCheoYdlUdtWH6tFw68O2oFWyvzTm5HRfOuK4u2PSanHQE5acwTKkrfHNQjfle
nBmElhHMFxDuX24htqWlDije6pAVAtumOVgE9tdx2tIg5ijIm2HGJHKR8UU+Xkyn
LlXJXo6unR0rBIeis5JmOBRArm/r/7HnDaDG0XyxiHdZPp91JzfRpv1wgpVjGMq2
MtYugJDSht+t3STDqCrz6aRoMzjqGCmuUpfSYoYDNlb/BrRD0OsZWrzbibSXGOcU
0yVWYmPj293LYO/QLEnTbcfHlpb9HNSrO0guuhHhOOAeQ78CUy+SXtgiMNmlq/6M
wX20K8JNPP2VUfVnDG+IFcIGmdGP2eK/rTNtN45gKHHn/RA5sim9MUnKvdsg1lj0
ZFLHjafnhtxs06VUsMRVqCDezPrfxeIzyXQtEP8CZrwOs+YIGXch7kyozynUG95p
pYHSJ8h0htjVYVTAVzyD/kaMdco2rnFzYnAe6Dq2UT4WiRqfM/glfDXH84HSqGHF
AbkIn2sXb7UJpNrIwCHOXlbRqRUCwKKhuB4iev4s8dBvcWxOj+eQcSAFq+zo8pVl
O2SwsBFmIyIYdlbeB8cFEIj3Qe2dgzdytSLXPPDKcbCFDqqotnPABHr7JS7Zufoh
PlHdhKKBoMXZ8SrJ7BXV+9gWPBwQCvQp9GuePtVOdDUwnkr8t2oQudiI+8h+3tHw
ChYAqqyHdTeq1xVMJNMsaQA6hrr4oG/ey75TqpY8qY60dkcuswbwvwlvj22s+Yo3
3E4dzF6R/IszJsbnFHpJqpl17pVT8C91ws0wMXC8nKEEMTdOVd4XeGD4v6fXda7h
jfRaeFuxIA7jSduJ6dtcAvY4d9sO69q2ILP0nZWwNRAkF9LP6Af8Zcxk3u2+U55+
hPFIJIN0CwveLY0kcDDRPHp4B6SBH9qfx6qDs3CGW7sHl9aRwaViDKdMH0KarHgO
y1GmLI18AfD1aCHwcMpdZQ7pRW4uFprFTbqPW8mGBJ1OFvQcskgdRBaidIsz6BcU
/YqYrccXHP9b+o+mpZNzPoK/TxKLkl2Ah1tFFYpc5h7GINUPcTGoXDeZtJnZSSN7
8L1m5WQ4Z4Upp1qWnfW27yat4mZPT7NYPMbrPTO4HdIdYwRlXU2QAs0ds0+zk+++
7khiYKYTse8vP2OrXAIp01cngh2u9UqA8pRQlWwdtyh4cbQ1OEQqE2my8991BQeZ
iTFIYHX5XzkDXsn9tRnzLxxg7CxLZDWs8qHi1kfWCdm2O1zE8Vh1VqvSfNAlRGFM
Kdm97FfwaeBLI5pcUtxXyrPnZ71W4ZpTZrVn/bHSPv6yvRztPyX60+CebooVWtpG
95KUxUa2cPom9zsYQBMUBb+9hoBhEWbHAas5o3EW24yUn7QNCklGWbR2S8m6cVfT
Xcban6TTzBotUVPP0TFwpe0xRZSZZUxVic0O4cIHwLdLLhgR8DpiZlbR8u16JAC9
vST1liyR/TFmbu6ZZZ8/3b91epyA9G+qwDwdWGDxOUSTiVGLFsYTWcq1z6I6e3e3
m9adbhxSEUPuYjvdE9KCC0/PQnnr6vTcPkMPd+kMMfmQ9QJxSKTZBGopuP5tE/Bs
u4dxNaGoTC4E08H54vWolHKfWsCN85mTO+uKuh0o5ToF/E+AN2HahJSpxwSoUwvy
p/zTrqiZ5A4Gbgb23JA7oKBpbHzItJPBr1PbUDrLyk0me8UKk4TAqBYRUbj12qAN
5cNFqN4Eb1PvkJFmdMkTRlOF1dYjgdOoy/wxNf1EIMBCd+UelscqKGDX4f0B5ue0
o99+7dEMuHqjNZX2SwwyvjoUqxatrjnOz7zzAGoLIaaKw7uVAnliOHzPRCQQWTIa
Ywn5w6a6ZqG//4pMl3JHRU2G8OtToqNYy9RFtlFoo2f3GrOQzkHdtti4Y0HdH9PP
2wd228AiSoNBNu2wDjiCkVLo4XPavMSgi8UhMuoPpIFIQfTsJPuB2E+vqIhYywc4
3DmrNVcT/qv584yOMENX2TN5x5fj4cgcfPEHxAF8DwuyfxTBFwRLGzVY4q2TnIAh
VFXqZibAtyLn78+vXo0xmhpuM7YdjwXloVAtg4HnaHftzQmTnyKJQCmSuHewVbjp
Nrmu7mrfhqHrEygRtcjwcyzLjyg1tf64b42/tOqLobUyQ6GPZf/1dUpsdGUyp4jF
TjAoNesmkModWr+Zk1wbsgFdr3g1uYGpE8NoCX2+cwODxUYvw3bNXXgVMP1K+RVS
VcWEL4bGc2C6ftaD2bD2wSIstKmA2SWS5gJM4WAD4zTGhVyapQRdBmIXLu36bZu4
dyEuu/8UGg+9LWTT0zWOEwuAINX+V8DAgzRSytHQhHoqW+1TQEsrcVZwDsg8/MCK
Ziilnap1fLYwg9f4Jp3e7jbBgDD7QPIruABSvDlTFYPuHdfzYjj6VlyoQ/vPzPFt
zH7H2JycB3cO8nV5TbHQtvNtBsAokM3xCpsX2+uh2Jv7Ab1MnfW1kljiWHjmUm/l
wRCPNbKE3w/4HsYF4rxpWJ2ZzxpEVXi5lK348uHz43bduWJ3QDdJwsfqV255v+4A
e7S5n/T899Vur8Fyo+eOglLB9njDQAG2X6OQhYLhaOC+UWYTCSyZLRr5PIDI04SV
aW5iQpLKmQfbFP1soiFXwvsR2tw2d64hAkWDKQsryoj5oh9k+bwcj4O0tcDfc9Yc
t8mDYuGSkTwoti0b3z7yjmpBPSgAkAUrUIQtFQjIsG7wAu/dmXuAcscZbw+3rKZr
/fFE6qSWfFHejK+gr/heff1aB43xyyUNxOTDFrh3PvMWjDKG5t/pWFqYlla304F9
ptOuMKux72txGpONcWYWpR5hYFbIyhUsv18Qmi4WuiyVeQkuzE+DPU+Y1SMLImTQ
vAPiEBAGgQiihgH0JZe5FeuyOnwd9r8qdQFj4dSKK5IR5hoDh0OsUD29Yf+nomm3
c0Rlb+JVzfOip5gYs+e+eWGf5dvOkHPd6xx2nZzKJCNxdzLjVdwew2vD60GGHt2b
yh4jZ2kJ1L+AvhLWWT7PxJlu9yvn4eBzLkjGVnDprxK3Arjmhcwtq8RAZctfK8HD
czsriEp9UhT6oq5mLR0VCBjvF7pESvaAmdJsiS2EX2vY+vINPHLkXWcS+I/0T+sO
ijpnoRgsPLvZb7+ySKCEWUqbW647n6wy5aLHN4HqR6xB7XgZom9/jIeIqDTvLKpI
4a3yx3vU+1MUmBZS0upKKF0yPxYzxDOkxmmTKzRRB0jSYyl0GgjQ1yNM8pgJjSEt
ZUOFVyC4EiaympDeju229j6YvCwd3c6JXBmxhtCCwym+wfQiDV468F6NYaVFWIhX
lGYXRJVuB/djbKgwHIWMWpZcbCJhiySKo/Q5uWWYsdigIq63h8nr3VPo0YWzBGkI
HuAhqkn30tr9j0uwl9hAREqYA62pSDapIYyS1bw9KOYz+JwwWHy6KvdPIAPZslyg
j4cyldMGO8e46M9pgRjK2FvNd+ZCCZDNHj6g3TRR+aWv0Ff210VCgtjiY7g6pdgq
CJMm8KIx+26f5oWsmQwVKiKr3f+9qrWaLnyc0pR4d8ytNA+gKoUA0poxKb7zWBE2
jCi+fJaoALsPyLpulYNIzdkkLJnd1a7RM/2Ya0E1Uoki9MEeQXab30zS6/mbeDm2
nqFjaxgt6uEDBSr2/ao8XD4sD4dRLH+K7YHYaEAIqey/8gcs2vHfE2MHb7bUkEXr
5DLC/kQ6OQ1VsrM0kuMAOkfGIXCdMtIh0+dlUIaW29zqXINqTLyYUW15zZmPoOTd
mvxQx+YFpT9JLv3DnsmnhSORR+/XN6odgN1p1kFiHC+8o7DVGiFTYHP/aMK8LF6p
X8ZZC0qQV0MBCxFHnYpk5jGx7aY/7HIl9o9Vlkc0NZ7xFGKFpK4HJafVT6WMYvGa
a/8DGZ+YYG4WfDd5kAz9bt94eXsTepuhjm/OzH1yzK1dg0DoS7nyjmNLkJ2K2An2
vz1dL5oj6Z5GU8hKLpB2EJgaVsHrNRow1ZDsuzLI0Kk9iE2wpmmXaQD8J/GMVqvh
PlXIQorkOh+xDTSh9KzIRlegcEOCopJtc+yH91nINhiTIsftA4qYv66gzThTeNNy
bVSc5CRbCENqme3v/Dz3RtoTs09QDkhPVXaFkj3IN8csFdnfPKgr4C8BpQyWm+9/
cpz5RgPTc2o72NXoQS9d5DW4EAlX26UjYPARo3Fk7axuTt5+1KDo/XX/+2SnmpoI
ds/jvA6Yhih31cQehqskcHSAWbZTSoDVen36V6DZHfPeeETAiEriURQHureCtpSt
keDz5mIToQuzSRPorCoJry+LimspH06fgdb+gC00pG/SKkJsDVb6j4rVyjMm3aaL
CMeb7xqB0n9Zo+sDw/0B6QQmmBWw9dnNRxSEs0lcdPjJJLNMrdjxXp6z8OF6MDx7
LBo4V4zvQgMS/MiHzIweXjLoOsiYqvLV7D57qZqG4B4v5713dEjxgAba8N1RW87v
jRbMSBJSjiJBjaiePLWNvsqYknerqYQ9MyQYSpELkICWb6HWilgqpW2WXbcJyQ61
Eg4l07F7E7vV+4BpawIiEYgn/VrCeNObpqXBInWO/GLZYRDpQbm00cwCuUKrlA+W
kEM1dXiDOsww9EteH9N4l5AsBAHUub+KH+tIIUzjScfsswoLglYGNxRVe2M0QKFX
47pVWRAzSEmO6XgaezG7vgEsA1JSxKEfgPGofL3PvCG7TBxtOkYim9CarAqrNu8U
mfmdzOWiU76gHCeMnJLlUrxD87ZGwFCx6Qkm7YSbDAFOCnkvK7sPiIUZGf395sc/
HyimRxD+QDQMyz0LPDfhvyX0pWqE5h0dQCIYNDD+80GPsAnpDG6ELDNym6OVrmX2
a1Pv0iLQtNtTLOl1Q37mT0Y66mDikAvqc8UU4JGO5kQ/VHdBT1d5xY+nDgFY0kQp
m1xm4MMf6FK7RYTSGp0PKbxHob7+P24SYVviQE+o+qrLYeHE5Yxr6Euax21O4KkN
FFM8F4yFUd5aFz4z8O8G6545CU0hyVthZOREgcwPW28fefJ+GsCI7m9ZZWJNatx5
zFaUA5w/qUFEtpOW0/LifKjhZg2zZTMHoFSvNZDDYW4mxeUFC/JLtlzbKQbN8Oci
ErAngG6kvxHIfdWKDH2NUs9quvVmLj5OmZKpzp9McX8KQqhE25tJ61dEVTsYW/K4
PLfF/fyPbRrQyI0/CxzGBLv7yMpeIEzy3d+okOzi90mUJd5G+fPoHJxYn5LGjr+7
m7QRgKwhXI5cFk9ecsfnW9cRiQvxUjk0WqrYEmXHWXH7+geF6Hp0OYDIM+OYKFQ7
6Vfx+NtOKSPkoHYcrdo+L53EyeJbNofq+PeNfnD9nNSYOevKbFZBPm59exrnxRqR
NPDqRmaTtBvUHgTV5P6JoSS51B1KF1wBm5NhZOhUyBZJxT7Sqst8XLT5p6ruBZSe
Jyoaw9+2ciHLS3jQb2zaIXx27ClISZdtNzMym4Dl0B/xB0eTcfopaJnpb7gMcmsv
ZzVpd75MGq+jXvzbVS0Y+lFZzE/ESvqwMt0RkCsKfZKBRdxE6N3O+5Luuh9GmY2S
x3NCbhU6qtDTzG9K52M47AXoQIPJpw1oVNbmph4EZbClP/SGxZuWUP03OR6c4X3a
7KqSChkHznaA3yv1TlWsKKeGTuIWDfSyXtgrFUHcUBx3voeqiZlZXtyrKUiMIXnU
L5BNkOHsRznJhOqdi8M3tDlg215iCw4Vua1d4auUHUeQaxWSteJf7slNXQuTri83
/WAbTQzPwwa1qqGlHT/B8HWOA3McfkPxzxjNKa8b1snOeho/9tg0pj+ppAa8YGf2
jKbgRTZQcnUEpXW/05Gx49rbDr/YDLwAY1hbjzxTdd7wH8gJ0oM3r7m5dZ0Wvk4H
53H8bsGesijMFm3FSmOff/h8FtasUtBZ/dBdg8APEPFPIQeQvG7kWYLLV5FVH/Vz
mZoH40ogc9ceU+skOJTL1tHiBS1tlz5Mkd1I0/eNS7kVqIWj+S8egsVVgQMSC791
DsSegp38DbSIcxW/INkfo0zNHYSGDR5p+RotvkC988v2pnqoPWeztLSp95wKNbGz
e0YxAv6JqXAsQvtSz6ubkZ3cA1DOrZf6XQyUtbVDCO49OC1StTS2+YBnSqIqXLhI
dCscM+bfaWA5WFoxXQd7eqqig69XInNkIXqr4sUbS8JDkLKhq4EBlKOPZU3nzW+Q
9XXJ2o7G6JGW64m1UgJjHyCOO+5H3dAF8fRr2g9M+6/a0yKuH6JR55rN/epwuW3k
2JgA73IBeEsJYghPEBoihh+Gm6Tusj2Nm4L18utQLyTQsn5X0069Su+ph3DenHZ8
iH5LATKK5btGLcWzd6P2Jq8bL7JYGILDbcsR+qrVXqAd8yAIDhaH2U8yUvg8LgOm
ucf42MRhrnqQDX84jMlWJzQnOA7wuAtZ5f0RwAr1rfDy8Ptl9sVhdrm2bYbnALP3
2HYpWJgXHVx21Nf5GvDjNpMXJ6q6UxybpwnQd9yehpBOlK0/ZwZfKoh3vcGDuA6D
K0crFlkHFrykfIbY8wLCuXg+7Hejh4pleomMv8THpQZGwWYugxDI9SlYP5/KNk18
kGIiUjB1ZXFAeEr6aya9Xefm/4bF4d84g+EcKUEASHdQ0bmGwi1n8rZGkN+QUv0A
QrhVyy+VlT1jxAzggfbAQbNlyaU0t6bcUA3JzPPNGwg6daK3C6VwnGXdQtKMChmP
3AQqtJf4HgipSdyfFhI/2vC+Ib/gEzwjmjDl4pQ54U3bXDFkUQKN4xwrEqxlXHNd
a6IlZdaRtAJh93Tj1cXHtIWFIgnkhIdRxabhe50L3qh5lcpGjbRv0qrNKNkAnui5
Mvc8eqTjzgOY3FD26JjG9SkXQZyNgDvjF7pVm9ooMSWmEqBMa2PQ9DHaemxercxs
/E4G3ZKjX390se9nr4pofcNFRFRgxuJ6YBGPeSH/1Jr4bihm9h5ckfiSKjXYWBO+
4Sc8MY0gTN/b0gS3FXBVmVV2CHDdUf6D0TlD2SYjuQDSU9cb2QX5qcFC6HQofw1I
BF0IyU56EdqJdrG0LeW7s0aAv5JIpGOwEBsIMFZnhJwPnK517FW9KLHB/wv6xAEG
ovtoXmZK6scNP8hfUxj1FuZaBfqx72GiVdf5xB84rUrOmb7nyagMEIVCL8pUgsrX
7FoxTW0aH50zU22QaCzLwYxn+vp8CY/+8VAvTlGSFBqtOAFYl2ohdyJlCVGH35Rx
7wJVeXKFfPARyx1OVLbJ3LSEVbh6N2OhQl0AEo55qEWFS31eLeguMTtgyp1nKhV5
l+VuOVWtBTmooQJlkNuMKDW6PlUH0BDtXqOnKZJhN0X5WQF8h8KnHMVxN2AsL/Sz
SzoYRLljxS4XxgToglIz+yEQ6XmTqF+qur03D0Y6UHQyiOxhQ0ZS3pLTDFEbrN8q
1akE6xFKN6GXW6QoX/un+JG2FKWSHVGc2m0USKiMAEKg9yyiQZ9UvVCQUlWFcbua
pC1v6E3IcfxBWna5Y0pwi3omz/E10ON7ius06eBtqBNILJfkjU7HZkZTaReIIM7s
D5rt/RT98ITaakNCjZ9PONC+Bt0XSSc7QE3rk0Zm6b3gM3Y5/Gnf1j3kz8hm/GZ6
GGma/zoKE39Hwg0l4hL7CEz3nO1wDsyaa6omLkbjibRtKAYyj0PF/Db1fUTWR6a2
YJj76RxzJy8Q0ByuCkRRxydN6jZnFSAPoinGU2vc375bLx2otZnKF6vdTf+8Ajb0
2e6oBqblRHbg56v6sfrQUXwA9UafejeA4ItYoa9ErZcrtpLOI6eZRgh9wFMrmh9M
5dH70bdOgeURiTXYRdFvUA1nRcKW7Ggk6l0KSi1xGzfz05/+kqc/EFW7W3BfjLis
9i2M/ncPj3o2H/3A40CjQ/PErSlqAR31d+nGr0EbYDl/tPd9RLQ9HJJZ70v+Rlar
xCu3uzSWWiTJZxaK25SSo0wo6a5VgHqit/TiRBVUUUxtfIQBw6w439k6j6JO3ItP
VR5A6aKIxRyBi0xvzJy/zN23a6ZBMGkQ96yXXMuf6mG87BNUg/zTWewcHIq5IkIc
rvGVtJw/GjXpCXjoveksq61JDk9i6B3Dx9p1fCrHwKo0BCUJTP14a5n5g5ZOkXlr
/zGDW4608Pf0Ed28x3VN/rf+lFebdMZyg5ptRTuXnxFAJpdqDcExFOvCqM8gmOPV
8w0jBoB89eAe0+7/+tAJ+E+OpKI1syqfplbundC1bBFY99oumBWB++W/NQ34EZ3O
syrdhdhXPxqnnbMB9dezSTpOBsLS5KzAHok2GqYhuL+7Cdgvckk1EVNU3sUv96RN
7MPE1UZjuCtiUjrKxhfQHB9zDv+2xoAyAjHlYA+wJEA5adtPbPp+zM2eox9GAoas
dQucwxMaVt3b1j6vCmCSjCme466sCRxu6DCiibf9wCGUpUqF1U1SF9wIGtJt5+po
q7MFBIFNG6zTzoxyjwBodjEf3ehcaz7o0RanLsclVYZnZry0uACxp2IR4ezXdC9y
4GXoVre3kUnDmjJXT3GSk1XOKyOcKzIdgldttBdsAOk1eycHAOLwm+i5fPxdJPbk
A0iVSOCOmThrsIa4+LGYOsVgv9k2G5pDSvxGj5/4I1MZw+MPK9Xg7NYMzYyC/fgE
SZVC2KXKAAIqZpzTVD/K52LhEfMbZ1FZtfz3SWnmNfG9WYuq+rliWSExHRXNiSrC
fuyQWw24scBGJMwn4XN6awbSB03MaiI8PUOvzsgudm9h430VEXs1F+aCX0zAxTMu
jJHUmQNp5+KV6VOio1Bq/Jt7tHyBoWEQtxtJGlPs2Ws4tRekZlaSmerZ+vzCghBV
FG5nSF3I1EmD25AJYyHZRjh5FfJkepaPNMh7UymR9jH/F5Q44lqhpfKyrygHJeRN
oi/FXoPZx558blNGNu++d511mYIk+b5Ft4SqACmrD4GpJzu3QjNInhK5XdGX7JhX
xkTiGPY23LJRNCOXNKUP2ARpwQtycy3V8uzweYZ9MuyiWYxWsiUifMcCeYLhq3Aj
0s2ubSsJCd1D89TJPRjhYgrFe2FmFmPuing5ExkgeYYlx/QkBR0X7yNCNLCCd6jk
EkO5BMCvX1Ciyouw8q1f77qqa+Zr8QGbKWsTolIY6QqzWMOqTi7xj+siDoCVBqjq
63S15UuIfh3TYWMvznLczUQWn5/F7rnQZM1APdTh6NKoiTd6u/7Zs1wOnv0yNePi
huWRikJVGs7QPJOCEPMM6bvtzi0g7M3HcQzvNoatj30i94QY8duMri8yITGiNjse
WTfKcVESsg5HIM5wD2kr78zE1G9RTFdp8aMqBWbaJwEiS0GntISEDt4h7IrjZtei
Eqi+a7e/ur/uookmxuAKzqE5um1sD79TCIYFIixU104N4KUiNm0bPNmo9I+myfxU
tY+s3kJYPDH+viyCAxQa/kWY/DFYhiIoSv/4qNh0WnblNC0X8a7xgjASjHEcN8Sa
hTbtKVr6RYKnleyyN9icrc7tcDCt8I3CQ+yv/tIVS+vphHFuugb9KJxv1fyTNnGz
v42QTKRnk1T+OPodkfmE80w+gNSurRefrzkHDN+BklTGbsv3266Qz3/oV6doRvYC
5aRqmmiHYVkKnKNsf+ACRn3Bz/odYJVD8LKqXnR2JorBt+MCu1gWT4xVFYZiywb8
XESkXPut2D0BOyRueBi7AaoKJEp3RHCDM7bRyJC+/tB4ZGcurmSpCNqQEVAOWQgP
e8SFdkyjwBgBx0eYtC9yPqM0OdpgpvtgJhxxdGBfQNcWdimD1isufbIDgpqwACSe
FWRjXkjpCkhw/8pKp8MtP13u8ex8nDUaL9TMwf1q1a4+AcbdAU9VZWzuF4jjDIv7
8FwV7L6uASLvrMpAHVf40tGy6e6ymuWkbpS964ywF/9FNHQRCuJ4oAy9hg0SHNrJ
AEJ4t+qOWOnPHlTN+jMz3E6AhXw3oDYu+2d2A7TJg5R9tYPOmrVuSSnaijEpvggC
3m92djX6iiZJ5UKZvM2arfNAg2ZrsIJsa/Yg7p5IZWmGy8DIziOQm4cH1c8jEGOJ
xVtCQbWXvb2aRl+u4cneL7Vtow66fB4lLdSicrpKu2N59XqHn/5SWAwXsRXZFFXm
MAukQCDXVUbsabOKSmpWjpCPsNjJaV8bCPklApdG964GQefAQrDByZbhgMRdaieD
fIIKHouaCH4tI7FV5fvcl+9BACelp5nx+7303gFkRNNu2YSdzqkzBK9DmqxhGcNQ
JcQie00gx5WG53KMDfxEx0pFQaig3JxtBw6SOZvZvIeezrihTfRMyY8v5FjaX6Sd
/ZG+vOIBCBz6Ww4zBWF+IC/Sith9qayY7R1kJqm3Ze4I+GPtniQ65kljycqBjG+L
CqPc4BQ9tEnwsR4lyzK+nhYcPPLCiTBkyN4BvTQgcUST/xQJ9KhQA8qZ9rEG2TvH
2lL/N1GPJZFahqWshBaM7/GdfSYEzt8xE1ZUUot3QuKU5X5CoN4XsEz/2PztP4kb
p8VMI4wHoly1lCRmdNgtP83gUWBmtC5LGinV0xD3OBtWBgVieC3if9ENjEFf0Izc
o3HoMc9oq8egIM9iKZrPv5ZQ8y4v2lkNuMoDX/mHRA+yW/lcQbFnSe4HArD9KtUc
jpcA5yc8odBRrMSwGmAaQav5yb6iWoOhav8OqfOY3iMuPl5Q7uglE1hUlpOk5oro
ObZ2jVZQNXGXEn+rMz7spZRrr6V6PO7aL+efs527yK3hw7G3/s6jw1LP1DqRe+aC
FDUqnVl4r+1tu1WBimCR00Rw3WwRClRKiX3l8rSKnOAsqU7YEXmDaT5CAqlWZOh1
BmARqHfflV9uB5jbDDGrZIK+4Y8fwt/I997I0aOnDgnmgrvWJQlvwU8X0PndMja0
t6WZuF/fWkK1XB6wVSdKFtxQV/rfoS0dK7QLcviWtxVrvNzkNCg7dRaGNOl9Gb/h
J1BWz+otAkmNicH2J5sYtMhgrxFDGbqPEQCBTZKd3YSurP1oI735/jMVmBrsc8gr
aC4t2r91Qh6O07AO/1Usy35fcMFGjHY98+wxflusEzJo+qFRjWUpXd+3zliMrpyV
JUSjQoe37tIx7CkM7AhydGTUGQ/EvA976eYTTnVAibOTy5HcK1eWUo4RmdlEtqt5
ifCXcFp95lR3jpjBbJwA5wYkp/xck7wXcnzS7+yi5vRfAbZBYEDDVEJEYJW1C37C
ZlZveKd6pudiXS0GxQPpYw7jxShd4FvhMshInMnyXv8cVjwElw0O1YMcqcdBFARg
MaiCCq1L2YbZkUwB0tCSaRxMKb4UWNiaj+nVjTdBeubfEB90ST8GGvvUamAfvGGW
UHY5R1My0eoxlhyiyLtKeWzNP0NpoWwChnP7HC4OtDhkyi9g2Erxyf9x7hZ8K+Wg
SmwPsvdvAeMqIrbJ2q9iXPAhtyCZYlibBCnOJXUkk5yigAkLz94XtMPpZvJdOoCA
F0cg81Y3RQ16fzyLQTl4WAXg/hDq8pGRDY+0qZcQHg/cBqdQOK8z9G+Q3ST9lcyY
LV4IVb9QJwcUHwoR+ZEGQE2HF3FIRWWXOISPOY+qWQl7FCtDwqwdXtYE/MgkOtYf
yYzmHZXbUFKOx0BLxcXZpzWv4XtsLWNB3PXRrTdTHfbZlNbEYe4YzvAeuPXBrNkq
h1PldhAV6bYAU7D69pMtbc4k9r/0DvXkSCLKech+0g20JBo3athALFxMVZucVzuz
3JMpcodN7TQAvu3m6juS2tEY+iVrpMRtHR5oMobUGohYOlfFJv59yO1FVSGXHM/h
Gkw0e9apk6ODoJUisYGrAshKscc1eR/EqgcmvUrYpBjvIS5JucjccpPk10beCXMN
pWEIqZgN4n3SvQmfbEUxosF8GbIMfbx8JqloWe1O0NeGVPkvIJ171aPO5iGxSUeq
bzDn3pocsbv+N2GCTvFotWz4EA5l0lk3HqPr9e2/AtLwSOaUJr7C2JULluWe2FPm
/gfAzPu2kz+C2chhiXbEx3MnP/fbBZ17I35GFNt+JZz/D8SjPxUVAmq/Jig19O3h
dgNQ6azGFq8/BWoO0VMY/UlV4q+QWhcdEE7Zlt2uYbNWOIe9iHLs8Ui0jVs23tgb
GZ1D0Lz4SPJBwAS8nlwOLtGD20iZf0VIWfopOY8TdJzkJKj18fpZQ4D5OUYcS+3U
NHykp8e/r3oe7sz/z78B+Hoxb84kwfG3M3xBf53Ltx2uWWUWPJTVNLIip8SxBPgd
YUiengELeF0YYM3n/2FZ5Lo3kjGChK9KJZJolMsfPX+n854au0dCyFt2SDx2tBDO
YnyrN26kTSeFGrQxzMWYzBRFnGlqvKF792sn+BwyxgP0ddPE9KJdUKtXO0NoxJ9k
Y0H0uSpSMy+sh+O+hhL+3iQG3WtnCJXUySKgI7Z+Aq/2SDl9K9f8KX4rcd/Eylrz
d4JWg+r5Ow/fikXIgo1FSd0c0w87YAu3prPbGHiAaqzRoiZY/WoRJUxfJbQ7fk4b
9mX+IUAI0qDNmkaqwERVBgZOcKCDBbkud8HuM+ZBP9CQRCyTT69B4yf4LDVXzUAL
4BKp381DMNoC7A56btUGMl/BvxbbH7Qy4L0knEj0U3gNI11Ibm59v0f9U/yINXLW
tJl2Tvceiu2jWmT/zUXxj170MHIWhXufPMYYrs9LlEDKj+iUirU8AjOZHR5mcc5p
k1MHlpLmzxKttqu5//76HSgJa+7e9seHI5fh1Pw9Qpxm65qv9nxVzXQO6TPYxU9P
/MKNPD1oWD9h2jiv8LS6SlvOkjxVWeL7Thex2ZK24z3ZvVdxFXtUpPIvvdoz0cFT
VOni2W/veHMSBGwoXykXHIt4BCLwnkcQDHzDOMGP6KZ2ePxxs+sqxobt3Tf0RkLX
eWTIyGs0P1UTZP+j+wuW7JJ3CG86Z3zb7QGJO+WGYt1L9oRwk6aDYz+c2uv+d7mj
77rAiJ6ZNrNQXVyIIFACjbvl7BhfvTcGuPavT1JkAnfViTIYBJhKyc5uAknkXYO3
/IBRvLZr8ESwycn1smunUp9v8m2v+QDDy579RN4MvxLcZT9Xxzcn0mCJ61V76QxZ
J5BNQjm31JwxvB+mSKj7lZzF2Tj/I409D1D2RAw9nxEwzT2XwI5ZGcFCsLH7JufK
OEUpEP6WvFmCVmSIwIefDVJlLEAh3oP2wfnTLAs4zO6tAVHetAY6kUi0E0WoYFqd
w8tvDDcsKGyn84248pnF9zP0Buq8akhw94UT4xfStdwD5K3BTI77UffQsDcqhKA4
gKUjXHYvJNhsRBJXW53EVwYkG6yzubiJTzVHxD2fQ21U0yhj48E6UAxKdW5RoZDj
S+B0Gq0Joc3RjhkJm+uVFrop+T2angvBRCFW/aC/rKV+X5OeFH89V/wYbRbE39Tn
cer+diQmjUi6Bj+pw6z24bwjpGkV6FW5bdsTRFeB5jbICimzGRBl8WkzguNhcVmt
0clxAIESEwXAMCKkh5GrUoOVXgYmzAV+uZdu3kczmS2HVttL4JrP/PusaKkgR58d
Igm/wpwnUyh7EQf9i+SMZRRjuIFk9tXiyOccmocLKh0aPkenPd5DRQs5gjBh6Xua
PNt1h+5FUtSJ8Dj5mzv6+FF9miW5noMCV5puLQdOM+GtqlLNULOYvWIQDe/R8uLi
eTkvA7VGSRWYwpaVkwR8AH55n6tqWvRdHdVndjquEUrRff+CO2KcUI1xelcRb569
bUkx2K+bt5Bioz2sjdtmqQKJkQ7fWHoqChbnqEEK0zhujpg7kdV36gcFDbpEf1pU
aYmSsm/oWk/ZyWxat2doNR1Rar6K5MjGkCDkzjCyeCAf05WccR11kcvGN4htHeuu
fBl78/HTOTiaTikQf/q3MxQ5pmToOY4NPTnjVohD3uVb1/pYaV7W058E7XwuwcBi
Xijkv97T8/rp9pG2Y1X7WdtwJlDz/qEZ0fdRU/FDu5ohcJLsLC42sMaftGjD3JhM
Xg6psJIzWYhVBcO504THUNXPsxDHyl4QJJoQgCGPXqw5K4Oy5kWJDbkrA091NDgU
ZIwKdDsG1FNIfeZcEoq7M3r54e/1EzIi3nbHG+5fpHcBCfRfORxIjTeF32/B9eFn
E1odoWDRonfMOsVhROMPbrj9YUXl2l/7/v1DGzhDtKOfJXSXARtd9uXAH2xK4WH6
A0kfbcKwsxlX2i5VUNKXbgXkkXToX9cvx2mfIxWoeLuOrNLJoCGu2/cI0eL2goZQ
9s35gcYUIIUikgNsyw6KcAhUmV0yF7g7yDVvyDN5Q+EvU6gVpsWX35dCCIGnh1h1
lMDHBMRxLqV2WeC8uQHiN43rDqeJCvnFtAiRGH1LLyRkJCACdQVtzLLdJgkdIXx7
kNMuRk/7Casix/tgyM8ZpaOQV50vFEf7uTtpvOYt4gp3CLPOxxW1kqHv6HYlETUf
SaslBIRzbbMPhohhRvm8kH0Vuc8+JNmbZKX2L1264UUChpQ4fjkeIzyP5/BeM2/b
QdJPwxN5dbONXyRsJCKl2TPDTSRQ0TLUYCKN3WxTnTs8q9Ue/1MpJ9McZm4DDjaA
1EeSsvUVo3SjzXKiMSfwcH1ysOqkKGqK+Ny5Dh9HPxNCPzNksBLMpZMMjQL8fj4t
bbCL23KWJUZEdXCA0gfJqPlyCi0+3VbRB3/QSNggd+BZkN+fjsGoFmgxS+FdFRaD
0XcAY+Maa5JhyE/+/FlyCUvcWx/Iijj/bsLH+cbo4WGicUrRTqPE+q5CKFUgrTG2
/3lDxgDS8OCLmnAXxYrLjMXx+99w8SmKRu7kN7YwHgMS//rxnd4Kh3p7Bg/QrY6z
+rm8U6LsNfull4NhZVO9CVAAKidQ7aKteSJ1YKcR2FdvH+Y7dvveQtpUrQX6S7ZU
TlhYXD0hzzACx2/E6B+I8h+EmhrqrcM5LfRBQmJzxMCC+1HFdfaTaa92GwvCw79g
SYvk7yBfKm5jTWlxNT/Ni4/O3to7AJE2sjOG/es8cO8I/GHaC877ydDbB2lXYWVB
8J/Hk9nD3BC+5NfJZ0p2bJpopa9QFgRIvnMpJpQjNz3ugb5wxv5HbAmaa3pvnw3E
EotYy3EG9udW465pSOG3CKJH9toajZsq6IqdhfBw4+Aps07njLNXldkOBGiPzFsU
tJXLIQ6JSNQeiX6Mh0kv5dVgj4OrVGUoW67LxM68/d7wYwvvjbTI4u7FrfZnBFod
ogGdWC5T5qxXmbworsG8UJS8WeakJLrEIOMh2sRlsX3/6/vUDxSjQcFkmBTKhEX9
nhzUasFbPm4qDQOi1x7rAaGOg9VMUD7vFG9OGWS4I2bw3b9EWRLifcnCUp3GFVJe
MZ3gYxdkl1UyeEfxhiNwZwdK36pHKDGQy9cG1x5PHwxWosBvO7c9Wut3dy9fUyPw
K0QeowzvcXuoLnsc1MW4PHuCcbsxAuVwriLQVGpOZYV0msBjQsYfX8uuyhyiT5VX
i65atDIJ/KQovXWCSkXDaa7mApmUzxVM8+eqSnd0uQk+VDSzTxN37EKv2rV/hASk
liK1YNWj0rQMBIVkcOZgq7Yc3F6ozPQTUQBKICd571hjcE11HMG3By8XanKUv6yo
Ct0bPHGg5v7Jz8HXax2YDkwjJZ9+3bYT3v0ns2neqlUdPow9clqmYx76Ohm+DnTa
gLke667It5Xt7ujbg72bYtIbv15+ncGdYBJCanb7t8t3fdlOOIHM986KXiwB6tQ9
ohUsDk5LUq3h62tIYrVkobM3TdNBCuunJhAnN+Jg8dLB4+PwIL8kGaPNlZYlID4P
qD8JLbrVMq8iAKFCBcRxZrWMeuiKGpUz3bzvFVCAlA4lyinKSQyTEkmyGRKSGpCE
7WKjsW/a2gy+RuLUXeGuIe/5AKgzCSgV9x/VRAPTUEG5OkhCZawdAZkLnzIKMq//
gnvV61MoqA1Dl7CZFT4P3x9fxI4eaGIXva9KHOgw58No988POTutIoptagyOJdFF
URE3pilvAgkdafLZCq0aHpFfohOHSvL+jQqFsHkryr49NO16T3+UEJw6YVyrjHG3
YitVDjE6nMt8AJ2VzdfjR3ThWV4hwRl+7+YJqha0kNF5murLJMhCuaRAzVvBs6SV
8AjFKZkATNWSiNk1gKxUXlhAVocND7XfRtk+bFmpmkQYcingQ/Urdt/BMVVQ7Y10
SKHuWn20GhwpYXoTqvh056QbaRizEoY842Ir8v80TqaD3X5j65QHNHfQ5mEfhI2d
DhfYpAoJbqvoiT9RLgIvuOgn5AEF0NVdIAwSuEpbBcM1v15XSF3JWnFWcKwHA9Tk
OtiAM9gnuHDmjiQ4OZfBZy7b2K1O7myzQf+gi8G7wCSIXkwQxKsbTzuO6LLB5HqA
byOvfia2z1fQHmPNtuOkHzfEiKuxCmfTi7/+3uAtyleY1JlVn7T/5UfuZ2u/8lD6
N4AcIrHYPn1GcsVe86zbR+A7q0FINyw8/mvEDQIS0b+Gbu94NJGYhwuAARGccMMh
HYzaB9W2VbSp5l1N7xE40ckProFvKOTWshjTdDZHLu7Oxa28IeB18+Mp89Apbelt
/ZQHkGd3l+oOkvzi6ugyIxicbWQQmOWaBv4dMaD/tk2RF/2Nioivotah6yREvtuJ
UAxO3otNmIVWtoH9/ogoJayXST3kugFwc1aJdilWO6j89ptZ703+hGvTIWEBB/st
2Hmsvv1rni1Ee5LbxHEFXR/282bOlDx2Pb6cx+lKK9ay/kYZl9s0uMx91kzYkkFD
5JIGIWjrHBPzMprw9TFaB21yfl9yB3uu+EY56yRK0VFaWv/fhW8TdtR6RY0wwZyz
mdTKzsqlwlXbOGKOwCsZT/B1JL/GlalpOIcPd/fQ42UNiqtvZTTb1juhS5L5V2wX
FpcRd4UkgENSZOf52hludPGg1alm/qm1+aChW6sT0c5Gd8hj6x95zytLN8NF4kxX
s9BxEpD/Y9pblm9wWL9D6vOWFM3LPBz6DFYoohG4ap8mPUm7H84wxKcp5wPtUsPR
xyIqxsXyHh8MVIXHrxCWao2u0xC/tGUP93uk5rA7t0dl+eeVlP/CHgrLVl7dCJmn
eZou26mcVHpdd3nDoodL7wRVcdQU8JzDEKSKjycevTJ8XzVSXJjYeAxCCjLHTW+A
6fLH2WdMnAM9FVHJSMEUxyZqRqoI0Hg42IRfX5WWeBb83lk4rSKZPQTC0nRFsnzI
SAPq2tJtqrI06fGtAgh/oXmEkRKtLoQJtWsrOjT0FJEbg3xiCTFRw13ZrplJUrgX
GUTycj3qc4QhUtj1agJK3giFNWU6XzkifmltqVrSsxwxaSfsBWz43FKji5r94s66
VfBbSLyELuPz05mrjKxyqrRtXOR9bsKjUxv1gx4KJCa98RBGw5KhDqTZ81QPgrl9
msA/jJFUmp2BT6jC3rqq56+TYagkbAGvJi9syCO2dwl/9qFDwNtJF1geX/1tfaf3
YCKUp1s6pAbRKPErYtN/rgT8+cxqTjiHgAQZt0k1HAHawEpRAfkK8plkx1TprcsP
eLSsVrbxfjBmSKgk69OpZxo/HF7bv9m/B46QZQKrhbnfsXCOfZJKgldKyrD9SBE3
Et6MUrcSnr9oQdoKIR51DVcks26PQ11lIIwHrs8SDfBuoIh6cZ9tmy+sC/4M+Jb5
DaWKKhrL+AdwHHIB17QuOmB9eT4QGlfzmIWTd8OqtL6U+pDuKRkpu03ACfP5hjDY
lcEkbUO2/BnOrsWZ03/ohpek3L6r/2NRKveyJ7dB8ZgtYfoXczedJcdBIYeObeki
PAqnGTYITjbd+KxZ4gpHHB01nyKJ7GPsVRo3gs6mWheSyuPlV1MEoQuu1LDc4/sd
UxIDkDZmc0uUclPf87+76HtdAZ/SJrvWufUnyjV4c5iEVcvn7iRUnatmP4X7VsbD
TA9dYj5nYtiJyffEv/WxeuPf58khkT0NPIWWZeLTImDqqlbHtqjTCHkg9L/v/PPX
80GZ+XzmGW5ivc/aWjkSXJMijzb/Wv/UPxQNakgEXUMRxKamlM91SJDBtFZ3Ejw0
KxROmjmhLZznHZmha5YRDGIA7//ZqF4uYZ27fnJbLU6VMx6eOnIKkFO8B9KT1Se6
kCT69Yel3W7pCDYbEPoRI02bkBjzayAQcLdZoHQ+5pw02qHyjDn8ktEkB3AcWgrM
yTC69C6f55BFKeSMCHtgQyXF2FB6zgs+VuOQPywCCiIunhueH3HnoviiOjQGLFdj
aPhCuZy65uVNqNT+ZJSVN15hNZtGin4c9XiMTPxkXlmGJ/kkthaaTk8zsPDej/7k
/6TSQbcak2fm6sdGcAM3tyzjSJ+hm77HauKqDfri9nDks/a1zJrqpXdOK9k+iVgd
rmS3rN4xvJ7NjUZ9CWWB2LL80slBkQoa0lUctykZQYxBsnpv7Vo9UDLb6q5bDfc5
pvS7uhKgvqG49aJk3mCxErk1/5IveybzZZ5EUZil43Gbe+FnQvmagU/nQYMRNyJd
lrUx1jWWUj/DKr/LVo3k3K3tMdvt1qrD50KRmrRKKbP/oU+0CO/WhySwko4xxNew
1IN5FY49gJ4VGl7Rimp2qZUU9rcwsx4kfxyUW7Th1tGxlv6lQ9usGw5xjTwPEg0T
cNxaOv3EW57iebakU2+EL4EjH4a4dPvdZEmMRcHV7BMSpBUHZnyd6tZdVpB2YH/L
bxWoAEoAzTQI36fnTw0wVTaYGEG0YEktni5Gb3twUDgYHZU5hmTRBzLlz/NoVoFM
l8vKsEWI7TUiMQjHzf8dtcUy+I5aoZaYUGDrJJl0te7WYWvQgwMnem0nti6TTlN1
MDUrOM3PWiimNKKMl9h37yyvwjOuTiCNX515QojxkP5/OTp55srgYTKmpUsAPHoe
JO2f1a3izCPFeryFh0SF+25eWjnyYe4sLWTETB+Mh8SpYP+yOSO5wK86NoNmkicB
J56YxwEXrDPCpBvO3ZlO9bt/LAcxlZdCSC+xACozInfKCROT1smnA8rRhEMJ2DHG
co0e3EExyAyQUQwiMX2Z/8Oc0mkUSd/EiFvuAxrvViakUS9bOB28N9pmDoQ43Tcb
3qXz6AbALqReJdxJesM0f4w5dLQJ3RJmSpiJnlAAhZXxyJJwx/eduxx4ReXsDpxe
x5dF2dqkYRrtLwpB2UciOt2bj2b7vtq92W84RVtZkTxKuzFpMot3ywjPwiD0dxF0
2wOH73p25bfsXmClVW0EwbVfRTzbnYcSDvLv2XAlmtd6YWIF2N7rQIlOapG1BxSn
zT2wN3rvQXNoPGZnux396pvIgWscmBrXWST/BnXosdFxDZJEci+kNxTGb+kmGnZG
JZfo3jMvjFL1ntWqSEh6nOSunbZ9j3S2EsT9EvKaP0rRMIQUfkphodS2grS6d1oY
vTSr0RQcEID5MEFCyXRkePwfZ9nIfTgOuURCTx7xnf+2mvmIjbTuOkfKtBBYunyH
YmaXsO4xj0ewEFilixK8z/GuT5TpE1HErO9Q/lr5mJFYkuzCZt/+c41WHmDxbevV
+WYOPO8X3RJ2Y1Eeeb0HwQQBgJDDo12Z2UoWOeciTGgXz/+8X3b8zhiAryTvIfSx
n1f/TkP/59pcOkzyNyZBpFXOAV+5s0RUbVqkMwet7oW88lNU5LdYuO2zTDguSc7w
WNiZzAaQhA4Qhzke3MhptKh7qojE2KBPkzOnXgcTNwKQoPDtM8ZbH5nFSLMeNIb9
LUk1zaQpZx4y2FkydivWXTbg+PH1qoLCGmkVckBBFcDTlQgeEIbGiuOip8hwr5V1
XM2rwBCeB1sYT6ZCQ6WEa2K+YhAp5cuB8EsyCD8/9QLdOss/PYnoega1EPza2/Vm
G7hICJAVWNuN4COAZbV4L7BI4ZPntjKSaXSFADGT94a3acUYzaYpslQH8itBDaYk
dPQ9lWwSAobBymqmjez6Fk4jk+NZtdByxIPBfWxGDp250c5a/VHC3SOodSLCIHPO
vadd5POKLn75eXihMfaGgmBxdxvWCH5WB6k8YuFqeYGLcQKsGZpP7mMPlwl98/M+
jkJhu1u3ghnNCGF5x15LuJ3v4yJOwi8cx4NTYdHnxlgEkRrBjn40JQp4MFDkDOUs
G9CZx7kqzsoFbGMpBBb2bAvSY+fPm5/4FgZRaV8FrVYu90aLGZfvBwu6Nqr/TWYX
zv7/2KRmYz2Wrpi7jp7LBTjHTuf3jrR6ftsL9ubK3ir9rMi8so17BUSg+gZAttnU
1kntbqzDPr5svov5AsWGqpGDm5octHIjJgSaQP55KXZ5W1fn1o5+HcccHox7PmPt
nFsNlQ91Ca1b/q0OhNkg39CE4I6j0/szz9CajVQO3jwh+92Uozywj1/GVQlKL275
3ghCYnUwEjTYWujfLG9G0F3q++fVC4mFXD6VZWxrJ0Id2Y9esFL82iAqMoH9gzFV
AhUF+LYhA2pdlg3QKhswg5VLXqV90UVzNkI8gB7SqhOcPcMyx6hzuKpHrV2XSIEk
AKN5nAXxJ/MZ2HeZWMIBLJAr2X60EikebE2EBH/LCap5SPP3ffwQMB6ueEVmd1R+
F2L5svURjQKJzVgq2pJpX4G4DZ5Xflqnrzvjq6EtOkvL4QxPHYTXx5xFQRkayKsr
u6jLFeOHJ55B0zGar4wp0B3gK5Eru4/WbELGYFCzSFLmLrrwVc8UEcPdWDXMrTnv
ShGiYC962sELKpjKYnpHHNez7GIdIsEQyh0wMk4yEKRsFRlR4IqzQIXNpdSWv5em
Z2XS/1CTsr4RzXF8HIHMKQ5IZO79AD4f1piBwRFaiQ+S+hnkGjNAcfmmqWPGzJjj
ktxbX5VudGfTb+XmNXCh+I1f05/7H0sPMlFQJxInraMC9TuIdAfaF8W7RER5IvIL
S34UN9z/Xkh7wXxJPvpKAGiQHsex0SbL6TVuzPO7lipV/TiUKYcwknyoLVFNmByp
N0Elr0NTQOuQ3XGqhweGYWype2uQAClF+IY29S+1q6p2sz2aAkwSyl/64EnkbNR/
Os5RnjlNHVDXN2TPyRWhCJvBn4XYl3J08DISSYhVPGNdgqC55CVOGIuWjl++L3xk
uMnfXWMq2cZOR97Z2bVtH97nLFitRlBUFbf1PnJbTs2UKLSvCngpQAMp7Dh5R7nw
1UqoSYSm2PMmugJ3Tdw+VXSD/9FWt7oDdnbzG9ajMGxQ8t/C6L+fLggHJSUxk2YS
lRr6MQ00Wb3Ke74y17/w4uLzLOcglh3c4+PoL6v36+kCrUSejccxGWdHMcoi4Wgk
QACEc9dydZfZ+7CjauRJ+LwuMVzymLdTShhePhlgcAk8m//WiFUK5XyQHkCx2xA4
pcqqyiJCz6GjFCguVvS2tdPKZ8V548x89K18f9wmThBJ7Xvesk9/ukQxCf1etou2
8G0Xxb7OSyQOV0oP3AxLehLzs54HUCa+DrM0r+9MG6p4haL+PYk2vFpeqcQG30Y1
IqraifzttGKR8zwYDmspyfLC/8xWOHqGvlt9+PEgk+Idm6cruPHGdm6OH8T1V/XK
EH7Dm/KZqD5Z9JC0AVdJGcZMcZmNfA6NVxK6SA5RLvKP7Yrf6aw4dbxfqdSlaBCZ
mOet+ijV9seDPxGI1gSwgmZYudVRoYzGJxQT2Qwzz3kKnt74Ro94D61288shHyR6
yAPvb1jNveOyyjw2cuef5qGYZmVkxTUUeJJG5jhN0g6kN2pNlHcJKzkfbcv2yZOx
iGgFpLWC/e6yBw69xIUNpNUr7GO98llpiUkttX2Y/7INYD/nnLgzd9dWC1lasUBI
5PHgFv0BQH/zZx9AkWzfPHO0ssTjiJwAMeoF5TTlIHv0dAT62sLqWqzEXZm2e+YW
2MIapVF+/DeaHSav3WEq29Ga8BOS48+DbI187PPx36CmuBrYFzJUOxAl+E7n7Ckx
fyxzDGvGNryO3TXzzWZfcx3ng2pvsfsL4NJw6Q2pZQ50cRVQFnzCoRIiMWjVEYDw
9HFVE/ViPeevB9vEpZrCuFIlMW1I+v57hbRahEj9x79vhlpGFeiIVxAezllG2xnD
K6dhJfirSDN4zMTMcPCcOiO6eB4YX41Fz/63xTDYnDA3sPmNwFDyZGpRKfE6ruxW
7CfrU6t6iPxQVAf46jo3rdjyRD3iRkjuY9Z29gcxnS3/ndxPTMoRljSDoqVY1wrU
0TpUc7WcNYOkXMm9BPCkYuqInMlRktHim7tOaeaBN9qq0Icapeg+fUmk4HY6HJDw
Z01leirz5lGRVVrqTPsL/41vAI7j/bUUDOlhh6UKDCEQs6Ma1DQXKHxEuY8GDrzV
9Ab/L9nP5lVqpUkK2pf10YLRcg2WQSpA7SR5etHRhu+qoVpLuhDz5kz7LXGZFWci
kNmVEW89i4lvIN0s/GGSBUOZwUsm72S9M50xQ21e0HQi/Zm15FgQNiT8V2bb4xio
HfL1K4/E76Hzyoc+PHqAHbziFIy+vQRCH9gd5gSkL/k0iXYagFGCj/zDej6yYrAX
CMLUP9VQaWOIb2ETDGozzxm6XXdti+VZsixur1CuFVNGEWpYgCJ5fh85WOe8oTGc
tD4C05VTUfSAJb44ndtOkYjm4UrfauVVmnGTQG9MjzwXq9k193hyUD50TO/BysMC
P46IAcBmCAUtb6j16Y2jSC9rDKUR3tXtwLe4dCwBqtTg7HoLhGBJpdSlidUVlDRU
Y4/hDH5ewK9yCT/A6V5cA2TPs0JQ4Bs5IOq3M0p3R7SXk9Llc3e7nMe9UTZUD5u6
Ou/qN/gSSjqMb5b/Rh/2eqtXDHLMw/ZOGcbJ7is5DPjBqRDhEZuxLM9yTLaVWRAO
ddPgxVUCZ0babLb9hJrsucNOmF8qZUmyhR+ouT209x2++ArYP4O+ZWNsl7KlCk2P
fy0HFfGv3LL/l3tVLdeDCYGCMWFAADGauPKLWOaBaidcBobQzqOJw7acrKhSmo3Y
kEOzLeuanB76Lh9uuRlB6zfTw87SFziiOMrPFIBQ5+EggFsLMq6x+AYyO3OCVo40
wW/FHfYA3xEBlV8ny/9E/BsFCxLErwPeI8Z3kABl+/xs9/iKXhZSgJ/38MpLfezr
MyJCfSh3d6xM0BinDnfZD2X1WmHOuRTMfCx6HJ8D3wxu7n1h3T2MiCRI3EEBUS/m
Txm82I6wgDei1xSvuLE9adCr4tkTSihuq0LeEV5TBauwE86p7lPmMRIQtr24wJCa
JRasUWurkrjnCC5Y1bfpCtMfHAhONp1sRUbS3jtJc5OdTPf9/BKb4uCtA5Uocmyo
0/kj0T7nTLYCZINwTopu+nuuADzJEEd0F6hmOlpza2dBgz9LsGKrsCZehD0QOf7D
IHQgqZJF9wiD8pmTZugVs4VewepWMF2bkNqI4zJ48q38enMJr8m3XzyrGdcbrhFr
N03Ov6QEDTDaOdxF/YxTchrpgMLN1ZKJiSGV8W1Vxkis0NqLhuK9SzEFDx+2nH2b
UowPUjaRV3amJ5KVzfvGHDU6/7dQQQx29uUTnMS/pg5E9NN2B/UcUZBK/UBBgYcp
U9PHkAhE1gE01NTTnqm0S5KUsy47rNoZrfjjRd/+D0w+DzJF4JOh3hZGqVrUfGNf
S3gYVRaRFn6Tq3pB4s9QlHVF4uZ3XOJ0gqzbCKa38vFJUW0A39HfhlDVfOJsuKbX
nkVp2xUTmLzuTWzZBjTPYaTKHyPY6J4wk+ux7IwwlEqLo0gvQg84JqYoogdjkalk
u+sKujGz1n/AcWm91ImILy6PaaD+nMaFqvk5JB7/sXBsSFYX2cJ65swILa1fX8AK
gMBdoww8DR7WqGCejuPUv+IfAVdtUs6KdmXtdAhfCdKKS5iNAscadiNXlMXK4C1m
dNXuOWzUW5cLMkVQJdmNgUFI52m301vJHcoAC2Q9f65uNPVX1kuuB0XBClfHJVYB
K7Tv5XTHZrTeSyOB1IeLbNhdchnSHnr8hrPsJK8EuMdJBX1cj3kgVxsrjZlYIha4
YI+IYYoBPimjLXB8c0sLQ25mj1EEFnwKsCxnPTChSjQJDqCMwNKGOrtCmybtt83w
lG38qLTsUSTVjQ85lLFw5BDXYjUCYwMzMFRkSxDowQs5KJD5sR1dWNCbJBnO6DdT
KYJrp+AgPIn5LPhZmzy89oUIrpRVvpoUU8O+mwzgcSLXkAEyQl/598B138IQiK8w
J3RfxwRy62CgsgLubXidReTEbtA9qwBo24xsE+wZ/WzDRpkFqkyBowyq02sHW2X9
ZK9hmFfzkLpym6kSAXyrf8F/fxp0BECbA5Rvv3c3KTa6IiMNY9Y+5XPXNpHaBcbG
8uAN98ow1gIejHG7VWE/36yBNd1xURdzc0ru09GbOmcBMCudGAcPFC2wVlvfDWez
5KXxd2nXP1yXg9mUTmXeU5w1z+n0iRDEzmG/uspuoCq4w4OlCCFYULHRJPWbCvQj
22IIhQbyd2fXUFYE2bXVsdrv4PyPL94ATrmXXSEbMxPiGG6WIuHMgI5oWNoWYW1F
7tC8DisDP8XbztiRMOoHkQeF6e9lnjCUbmzpHJ3jSoM43jypQJIs8ty4DrTW2Fqx
JKpn1iMWbQf3XN0mDPYuACGG0HdgHXdfFEA6C/qwXZ1UE0CM7s63/5Tdz3EV9CUK
PxkH+NcTCghRpmGXudCC4EkoBciv3dkBvj4RSestJfxnsAIO410wNQOintABPL5e
6B+hgQ4hlzTis+gJB6bx5eLBa1s+334gho/8eCSQngyKtEh8v/GCpCIozDjncPuA
8HZ3kNJnNUvgarA00zjwAH7wmMtae2rKQYgyr1LfXjZy9YNKvDHOX8//yWWxnXDs
y5djSU27xUUH0pTcVtHeRkwYaNK9oVNLCArBEa2iG2lXUTTjmKiZEUM/mrSPKWcV
PjcYaQ8zL83p8HtOH6nyjYyWzqdeSqcWoK3XH28ESJBJNuxYoiTkS9w5lTdPXiMD
tLCo9k1gxNk2mIx+hdIAE9hS/BQrkkpfhWMSG1xLmELC2cjlEddUAjxSJO6RiWI+
omhNlLFJiPU05sxa0bmxc2a0v+5XD2top6PysdjtWXd7f2fMWBD5oO/IFAPcSA5I
kYfazfv1q8y+JlY5EHiZND060zKynh/gB9ZuPPnPoRTLnFSDUTEk6OlORRRJV66J
43V3lLi928X91OyENOnrvMpnd34IIjF5JuIJs2dO0645fovu0FBptk+pntUh97mg
eJuaWCfwLMXftjnK68VwbY8dgHlkPFvKyX2/MTCtef1hWbyntumb2WWSSUg4moct
V3n16raTmjUqVM1+fjr5wopOMmY9e01BshbELafxtBji60JuKeaS+0vX/EywbpcI
+xEjCwrJC4gMco4J92A2LfkvA9D5e/Wmy7fyp9I3h0+Yzcl2UiJaefVq6ksP1pHM
xowSPdmMDP6aKy13keO0bkSLF0deRIqqL9pZCtmWXVgAKpjtAmYlrBdUoIBcTY31
RRWDmhhYw1VoqWYnJkGZ+ujEcg87LZPGVaz21jd6rbZ/k5QMCvQUd0mhlGHDTGx0
XNFTe2KljSvbxx2yDebPv/IKbXLFYGQKqYDdmKxTQPevvu44SktDUT0W+48M6BUJ
cJacGqwlP3nGpgr/zLPC4TQiqfz3L0TtFlg0E0AnDungIC4TktPoMOCGl3a3ANzM
9LviDQqjFt7BYVetmzSm+xBGlG1dsKcJ5WNxxsseopox05DvN46Bt82t5hYJQNyB
6oPsQvCCq283xyphBM+3Qmbq1Xvi7VmKluawUNOW366Rv8zWuIPC4x9zb6mrXPQv
BqF4ujQH57Fp9zNaP0IEsNfDmX8mvYw/DQkzOPDR+YaUEyTged6ElJp7SNX8BjK6
tjtUofQo2lBvGnrrICzBNazzsorS3e+g10T9rlqa5DQMXGfN0ZafZ1RJeBrulneW
UZuEoV3l/+36yLYIgJbmIjhoQXqoFmCrD7E1iLdFXLSzBONeZtZ8PrP8G9dlZ0pZ
pwALlqmh1n2vaKoQ0a4m1zyH4NAuQlQ0U0dpzJn2cuC8/EcYAEFrHrOQ2K+hy6ng
v/bkCv4FCH2CQm8WmyJk2A0EbFV8YH9MNmtp80NZ1lVywcU8989TIhRGIqywYLEO
nB1GtPu4HTm80lXsgULWb++yE8EQbdki8812ILIC+hGDrPxoqjq9Q9tiYTOf5P9R
h/ujI4wTVzoxxuE4mMiKItmZiT7QeHnXLUWeZoPCcbHbmmcpdGL7qDfghg3481Ck
0Rezrf2T5Y9WweW7cbltWBKeP4a1Svpmm4LG2sIiU91AP5ztJJfgHZvg9Zgj+K8e
Hyd+aGFZpiQFbXhhEhKPDpN2c/IuiZ6mEWInyDmx5oxbF9eW9ywZmCls9RTGRrAG
X+zrl6QFomxbJMxi/kHNta6+plc6MZ8qhvrHpS8avQ/L4l0aDQXnKuRPLkeb6DHP
qodahuiGtHBu4ucONKkqIN+K2f7BjIMCnIKj+Mpsa228ZxtxAjDttbWa6YueFsM5
AzBX07z0vVgWgHapQKwRC8yoaS39MAp6JsP82NPphNxBYAC0ZOUDoRxRbBkDkNzQ
L8CrZyjmQi98L2lZv6Ceae0UqBKdkLzpqLe91DvSm0Eu1qPCgadt3gXEqTfAR5++
FyW9HifoZjOhE+7GoXPvkt72zBpeAJrL5La74QthISZNFZzq5tyKPYMdQvuu0EQ/
wxQfnEXHq2SP9XlluH0TNpQCjxHQBnVRPWjU+mlX+iDYl+5S0qXNfSY7K+5R7dK0
BBxUHw/XDjZaqGnXdqPClgHhj/3fy2YfGbdA5qmsBAAygdwhlPzkg0080Lo7jOIO
1ZxsawFH4tGdd48qa/Zo4wcaSr1ydjQ8NhwvB+zWIjbgQK52AbNUpUMk3jRQPhpY
T0NsSN0XvfkeJlK5KN7+wxBO5pG3lDGYEcmvrl8eXZQMydjHowS7MXbXozV7KiCu
l0TRYZBBCWnI+civG5uYkzJMrTjzAzFXnOb8shS/nMzgNj5Vdo21j2rnY1ceoEh6
JLSDJzjigOSgnjRNZREX83pNrlEtUGA8RTjCST9LWEFj7OtCz5yPX+od8v29ghOw
OYESmizk14EALgDkwseK32l9RnIo6yFS3f9R2/heNmOpucXxiccA80q7KQd769cn
EKH+WSGVeX2+g1dJwQ/kBOWOqbWNUu67HCbhkUA8inWIZGeneD4C/4PG6tRCabpX
3TFrg5rxGBXDnqJIwX7y5eQX+vCdrCvnHsLR6covtyS8Z8611J6Pxb56lrZrQeoU
XHP4ffN3npjqTfVzzCKNYBkpNBdR/SrPJp4zrUnbEuSjza98pBuj6wKljTs7Wr+P
4eqypVE/v9YeIgVINpDISNqrL7twlUj4KigTWcHiCk6gu/vmsww/U305FjOa0kvV
pA7kF0O79pDCdmO5CP0Ty08drLwFNjEiscyE94CVUW02cOkxB9z62IzCGJziGMQy
I/nwBvUjLjdzKCmbHQLDZ2P94wdTMd2e5HlsnnnbbH+xgHEsADxr0kGDKvBxkLbt
/8cQz4ejuzEO0MJxO0V/JDxL3hu7kCkKqbEu92IKnWxyrYa9vH9UHecGCX5yjUZu
73Ud3Q1Ew1BYYf96NX35qAzJiVygXcKjFlLWFOpQHACgf85wDjjdad73ZEOvyukh
gkeFtFyaPo46p6SA4tJS+qMl5daviJjfq7YLN3VA5uEV/4axdTgIhwSc+8b42XUx
dnljwYIZ5M9a74GPn1tOZxr2kEhlS91FgN1xj9WrzTUhQslB4McznKvqqDJFXHl5
XIoHafOTlsvIdUFr6LxiIpYZmLl0kHWJY5JWpY8oGcHM/StSvWsj724Atk1y7L4b
beYTGwjVboA/OEBpZK3O53dLzD3jqBePInZYoHovrRCPGoznLMrWqrS8nYQLHqt8
kvTtM63be74x6PLz59C+GsEP6i0rWZITCJW5Ln8bdnTZzSnVNGwa2xob4rvdhCm+
t3L6H52eRT9vyXwun6HG8mLBPWHglVQ9bDe9aoJYVTeLEBRZtNXFogZYXr8+HA3u
EOX0nQwE7nS2ss/Ud3aUSl+uvIFXLV9Sbcvl0WJ2SLCEVK6KiK6fN4MqdG+Bqquz
pkPmSMtujE+cWXMiJ0aotg9J2waEcCeEZ0pfLjg6+we3rpHJcptxhdVo+TwwZHv7
z9qafDrPcEBkLhaDZkznZY0GnZVHpc4MGerYDaj7RuTKsYqXtclNcMgv4lPreOmD
4vYQrPrAUkBhWf9IdMe//ziWIhwsXSCdFsbjvkzTcqP19an8AGbpMhnSmhy3Sove
kuNhHwFFAgL5tnjpXk0eDtDt9oUKZYpdKSIUQ0ivuXfLnES1Mn75v00UCcIYkqlU
9XEwX100Z6n/9XL3dDW8Xc/lXcX9b8k5QUh7MZo41UNSNzX9Ut2Bn9qXEN3Y68bS
n3nDawV0UNO+M8C7ICYBkGYTUOiNDY1/4yGn6CUsUgm76I5c81doqiPcemt5ehvK
Os2U1RLJIeh433MifTtIq3clAjDZ7LQI9FA2A6NZtJ2XuYzzw+0fq3aNb3jcqfzv
TXkSrHKTvCy11EKSQSPhXJKftVdWNTTqwwJmhcKWOpaelL94SZhCIFveUoihL1S5
iDbqBAiPy9EMU1oH97JsDeRq3hcBSVUeNViupOo3ZW8oAenS5vx7lb154/aY7OZU
S5vPENC109mS9d+i59QVLRT2EqCNfVX7okmiwy1z5pEUmpePxccayIkw3ovv179O
ADmBoOhqCOP7v+OXTZqIk3LcXMW6tJqb+9J0fFcWEGK/x4caXuI+uqGmRuU3fF8q
t/bfXga1XZQIJD0oPx5UuAKMXf+uUeEkBfhuGDysd8cjUxR/TtTKqfTDvu77Trlp
qXEI1lL8mfmFl2vXDatfHncOubMuGB6hsabHNKdB4L944DZRpddCTT4+fiyLWTrj
VSE+qoj+4PmECP5QtEqdL8lasUH05oPHxTgjO1l/vysjRtq6nCcTZTcdP7kOUwT7
H32Jjg6bQkfwimZSHHYHWKxTKo16Tkvh2M7AkwTU56aE+sY/v4ao7WCm6jF6SH66
9LW2hW+wmEGOM3Ne+CNpyku/21Zx50xiUHP9JefWPKM6VavUKpFCF+TrdO3Uufc0
GoStI8lXZY8+SjgvH0bl01H/Dk5rNwo8XK0AqJXTjfXeJkty2POEnMQjD9B2qtop
8h4Qws+wdBa9hxZk9xtHQQR3wYrCHrGIEUJq3sSx38H2XMwDmSO4MXUsx7lwANvT
o6JmVPZ3fYy4R4HCWn5EQ/UqSOg3Qrzb7FvfXCzoa2pdSHGea6tvNIcjq3seDxS6
BhVwmCJyOK9ZBtA071ExxvUoi8zPiYEVazLeD2/eL+rGA9GzuvelCpvBz9qrXLSo
i4i9+0J8kh0ERJxY02sg8vsuG/lZ0gtuiK/2YsoUOiiX6ULtwKIpzrjeKh8YO/7B
P8GowN3EhTNDqACuF5LuJa7JMFs04DZgeRVI0CpFJJwjXsX9DHLF0WhTjVGCkKSE
GEe0Cwgx8shPhg0BhXkQu/4XRMO2ed7o7o3iq/BI/MUhB+hdEOSWDg2Gjs7aWm1V
SbgJMBfMk0uDCOFckbS0pPJU+vNGiKlAOl6QNh1s2FY3q/oIcdx/TI3zp+5eYVb3
QGG2dZ17NOQLRLslNMrDfwtbJVoRIIvqakpD2UY+Iq/Eov4sdNjhs0R8FONRJ1w9
aVijUwzHY0Uaj8HxbUFVcqlk5gCs1wy6ZlRKeD7OXo983NBTtSuJJMTaeOq9cKa8
iePuZeQpia0LPwaopobv5Hv4aXDVd11jTEIN08KjnjTA1PEYZOVf0OXLrsUm1hkT
QRp2ySVXmxn8kzx07gkjj1t5lACi9N6P2WInYVgTpEeRbN6QhauNCQAeLTTJC3JF
Ssx5UeaynVNUOJ66HGTXvr4SoKK8YLeUARQFOrQor7xGjyo5rC+nroC7C1pvr/PB
zeSUXBQZiZoBUqX/kanZtBoDYp1pm5fvKOMLaeiCSsxJyFvNWVmo+94stxGz3iqG
z+xUYhfIOYXUZqs+JWSYLXcmjudeVB+4/9WkcFgbw8C1/Ne4k0htPFTNhCPrgC4N
t8bCdPvwR56ZmHx4JCad2TZKuvlFyeOYr1CI91xXmwk3G2nLqHLhVzQ68ZAMshwM
WBTbTmmDZlAFNQ+D4Loal3gR5jZI4UGbqGRWsYycAhK3yY9nDGz3TD/0ARWSLckU
C35BdrMfkqMkTghT2+MbsadKq8pCD2Jnai0gBsmnpf+Lg9nVdwmclIqFngIcDDaq
o8Gwwu9kMTd3/smCpoeDb345eX9SZ7d19GPIo92x/NEb3RqKt52iUxW3FStbTNCs
MwtVgcLliiZCNaVd5wNgZ1rQcOUvXh6jWZSLZ6S4eLcC9mespo45oGwSxkujaj5K
ka1Eqp648ze/eSIRDTkbwss5jy6beD0boAjh0aX8y5/adW5uFX7061WZqsCvSdMJ
l0RylHiWJPMvlQfWLBirAkmhFiV7VTUa/z8NY3xc14M9L5apQx+zF668CR0bcW5x
3NLS//SiVtUmlOgSvbYPfs2++TBe8u0Fu61I0h7iI0Fmel+CiWAur+ah6yi4ZGM1
XVS9PTO4gl1+CUuyjcoWXoRevQ0S2mUZosOXmziPAYXZicn4NXjPaBkJtBW3nrJU
QamH8XhRlRDfi/UG8Jd8chCkpO/283O9Yp/MorXTpdj3Vl1cWh5PY5c5LWLHZQ/h
SbV3KLBV3AeSnfP7AQB0m0J/2mpMAdkjbeWGOTZUQGljOyi0+reYZXZoMvwNV+gw
fUd1+trd8EOa9vzvoccd+zPc2fiZ9P1j4esdi85mS+LwkJZHFgq2XK7jCeRc9Qou
6lyAuTi2gW6s8HL1uhSwogXpMtxQNsx4Mp6T0q6/EIcuM3TltdFyx5e4vwME4WHd
lh2RiFPSwu3/DNz8zM7jijLTzxx5x5ztZMcjZS+VC424MuvVkAg8xzbG4mM6XBm1
b0TK2miL7QckAdVcI8bNoRKWjwfLxAI4bxR8ufkmlyhhv+jEzCg7oq58cYBwAnib
IxK0WudcoDIgjL4IpkrjtA2iwMnI1xdKwFkH7mcUQBj67YMivIXd+5cheCnxS3vt
gm/EKGpYQ1ptizO3gEyalkVv/+RtjDVVtkYD1Hz44GIn+cckoZpS88i0pppKlfzV
bdd4kMlqnk02Nt+YD9IibvnOL9z/vJH5kSD8Le8UhnyTBKjKCpV50TlNZP6QTdkQ
a5U5aLCWd+fVjSZiVI386bXMG4mtj2uDrxYuSbu2vHe3IwbZtUsfyWSxtHvkADMF
lLdSlXNYdTUEmsWiLb2R2fJw4XtuZhWgKmypwb+7sagfL7JyDzRUi7t4n2nZ4AmE
5u/Lhc6uDk1JinSv884iJx0TxsWBr1hDWk0azJHGkMRvqNXP+NzcC/YmwjDtGAWm
RVhCslDlpOliJPk5RSLBG60+GyWjWfQkPJlibHj7swBQRswLe+WOR9wqsErpHJBt
QGZs0ZC22+nTFsTbXmx4u7Ft/HpHUZYalRqaA0O1jJQ82ZK9It3Xt5L0hfrZ6e2Y
up6F+qeri1P2PUUffol3Zpy7jOzYajyXzLyG2KItKxirxfcOiWvqBaQwy5C4yTNh
7cFqmdqBPZX3ZtM34ppWNh/QpJ2axTFAASnWpXAEGxKuZ5n00grMXjH2jtKqvk3+
3mxWGbtOFH1zDdHJfE+fOAKhTi31CpwzgfHo4POOQfc2fnyjkah7x5lO9uAEFt5b
Tr2oHXrdHCOjxpM3ev3eZH50zM4aJAM6f0j+hZhHRFz24HkrQY8jwUr1tQk9GE/D
GzIDw8XGGy4QI/vW5BDWZSSabcOIZNDdSVvgakAqEQe0MdyPmFtCOrC1MFhCvfuo
xkp1XpxzPLU6AvWcDvbuzMmlqLhQlMRXua+kbvd6Kmtbjl+qW6J47xAwdpZ3PP7F
nQUTgC7BS+o+os/MwGl7HSIbr/QvO6zgMC/vOjRz2Kb+ez5eDQ2JePLgYz8gyeDh
2TXyGho7kfB+xiO9lN5RDaFeWz9fProEIlFVKYCedWKR5lUYE1H2mBAWsFVJINj7
f8niae0Og/UOcre2CcmZ1Rqx55ZNOy/CfD+HDV3JTKqvdhDrui6JjceflzETi/3z
Rqqe7jxuemV9s4+pQBqZ6QHoVchGJenu7Nw6hc0+KdLR6Rk+tclurGCTJ2+RjqBX
pOuvl4lS7jTRBY+nzr3vYp8dgSkMYiZldPxz76zxQLcMQX9vXZ7ulJ1eQE5LZdca
/vEumNBe7vC4SzlCqwEx+iLTK6JzrydcY5PvQjKsT1EwAe3DymyP9EaUY7bL3POc
3q/NA7AlBmAmkI8PG/nGnkRh+uj84zUL7TyMmFKsjS/2AvLdPnpWzDztvCIurDY7
sClZraBAbCQE5mdLjSpfIKND4osS8S91sgdt1gMCWYtXMBhRjNFJKW1v/svyDE9A
dVOoo6z0Y+bVCXu8/7hVH1RJEQ1QQD0B2+KWghUsT54vV9qL+s9fbtpHYhUpTOZj
wrprQmni2ypwF2lXpzfqzf6R3t/hI0iJkrkU8e4AvLodmkzTxs+rX2cfe6V8+iep
cy1GtUTZaz31z7sungNUcziRL2N9SSHDxcQI1nZgmvkFRZ3Qq7y+vQPg0TTInomq
/qFDaNChsYBtwadvVUv4MjOo3zScYyAzVvQK2IStmKQsr71WRX+J7We6e62vcOkO
`pragma protect end_protected
