`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
ciOc0PYQJTIXPLe39cbXGN5kkiada5S2GsSjCYR2PFiKiM5LZW/TOpdHlV8IIEFs
J/vRIlXrfLkYW4j/p+tVCtr2urHKYEYWpMPgReorzsy/Icm/6UjmPPVi8wKT+R6v
qKjJA8vPTj0Gz7eJhXZc6F5zBpzHaDpxrd3Ra4bVrSY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 14912), data_block
7RkF8wjOl/T9sDYE0KTESTaSuyzuLJ4PlqaZcQmLLuDu8ECZQRwZg4HKuUf/pZPR
0zd9sPxzkUxhNod0UNVpvQJbycBDdWaZJRUORK9rD9tATIPB9uz3uiX5AOby/5GL
AOVBHHWTHJ8VWCzPSupu9OQ6A6niZaWYqZah1ePWlGPprhaAmRYgvSkYhVcC5627
t4iWYzmUCelDDZ0d6xvP3vKGijZh2uA2fACa197wAQdOVt5uoxxb0jUR0BQWyj1Q
JgbcrO38buvkUGw+vvoyamHImg91lgOIwWVJA/zGVNrAVZ6RPJ/K5i6mCyXlWcuL
hpU4QLbGMWWQXNLO5G9dvDWsxiVGoGhfIrj0ZrZo67LQTclXOqxbZ1ZbfO7bCkYC
+6DIDlSL1/sOyPlFMW5J5aIhMFv9Csl19h+3sTVPKhWku6BTEKShkdz81o97pYEh
g5TPbf3P4BY9stYjZIQKbZb5m6Kum4X5zCgV/8+qMwPJzD0T8RFZgp/wXC6zPqem
0w2OUjfLo/UrRBMpsmKo7PM10TIAvmrZUW6jNhkS3qCQ30yNsvTO0qqm7xFwvH99
su/gc7vZXIIZYirB/yHyVXI/H4qsG2h0c7iKe/O+mIbvRMnmRsaqc3gbmG08LES1
8GlDcktyLybfQGYK5oVhCs6nUDspD7YkPcgA9pTrMWIBVVlbN6IEWAUB9EYCEzHA
pf+gLoJW9BYHrBTZaMvyIFvbpBZTREvUhZJ46awWoFRp0iKOdpeE2tqytsxQJiQL
kv+AC9XeAC6RIU06lF1mEITD/Wp2Sw87BQ364aznKFrUf8IFf1ZgfRIpfEeffM9s
YNYvOY0mPAxqSin4fsF8JR2xvxUSQFS1ZVbOGLFhSgF8Msc0S9ZNYG750kxUSwEH
TvjD+N8DJpNuWYfn8x3yridvU6oiT4bv225krwZm+EASgjvi57NetwqbmVu0woSV
H13kmNYq7NWs99lyC+M4XAs5W7j3t0QmHtM8j4TXr3hFccPNKDhZ7pPkSOHG+1Sl
7QrtwitNrTFHX+6YM22nIhv8zZ25veDcWc+V8glEwxTO4cCyVY2QVG2psiCvFaVo
QJm5srwUKmBz86oEW5kDhzBWcqAwvfUiZnJWAcvAPWImvXXoPh1KWELVOR5rFl8D
4hEOiFg7fwMIL+wBHUOXIapAHuMRkjV/wq52XZjzs9Isigd9BLt/6tevfyRWk+0v
gDv2UgWlDQaN/K/ft2x0Xn2Jp0EKD5inmz3oWCtDx0d75NBMJzb0T0nNdSZBBz41
BgEkxj3hDE+XYy47Unvz7PkFZzCSibCArgSX/dDnM1vHnwsYQaEepRASVJ76huBX
bdygTLotpZaHir6kye/exQ6+jhtqifw7z4EJEwM8FH58Qck80F5Q6524Mp0k6kS/
pOPNqT/4q+aH4AF6HSeiLWbVCMqXNeysA91UaHCLm/12ok7J8nx4tTQJFRND7wus
ehiFdWiZZccKrDighD7IgdmT/hifVlKu0vy7KgZF/IP90ztNowy6Db0aGXKYn7VB
ArOR7uh0wTg0TFBeE2gy3Hj/C9Ds1BaWK2rTGcJcSTcBgCEM1BnPi7NxuXVqpx/N
hxQwYvAty0fmqaOaYpxjWWnIqVwgTnrj8DL1H759H2x7oq0egQj3VV5Nbj1MdTxH
xh2WRm0nOH/GVUb5+1lh82cwKG8HtaGbn+U5ykQDxcVmDvA0GWIFVR6PYZrb3S9z
ZFdfblpnEiAXoCGziPdLgJrZUwMdNYRDdiJFPxCcTEqz0FxAiDo2z5dx2C3ctLla
9fxvXkqsrsQoY7rmIH1VASlMTxHJPWeo7r0BPYU9tfyLI9qsEGVLGM2/JmBknCL7
Jky9G4AZtvhWxqerSXqT7YDw5gP9UoPCkIa3IMWZqxMB0k6S3DcN8rHCrxg2/Bsg
5NvsRUNZTiXE8aLiI2FNdS/1OeyyIYmqMlbicsugqloO+9jhbGK+o8SlsRSX1QFv
hsr1XHkXLSw6nmrnLnScAH3LskizI4j6nXZQFCIEwnrNQ9d4ce68bXPaCAx89Mnu
uyagDtC8+okSavKprGSOhRobq4XNjt0X41Zoerg974fXqvx1WLb6IGlfWakz+JDs
c7spOYU8FPy8TG6Y1Xrc4RbIx98MPejqQ+QpPpStRUNVOPneImW1HvMknePzg0b+
Xk7eUks1OfOvvQg0IqtE8wcF5B8HOZfec370y/jpM2EQwP3lvURm3+mOPqGQ9JFu
zatjjnbnmkupNGXfwwqiIfxFuAJrK6t7OTaZfsCrGhVznjm912wYvEpUBxkE3qqU
puDtgweaP5IgPH8w1/7RmJFR4LAhF5p5/bNNq+aSRkTwy/baD28K88+DQZyfaJNM
TnH0/N5W/LIjHFdtXfoiIqK62mEJiEREVM7DWAsNli4m+XyPxVOLuDut1abIxzsf
W8HVyZgkshbNSTcsYmrLprQJm8ui92GDSM84SYHl/VEct59MWCES5HzyymmcftjJ
xCTMsDx6YJ6sGq92xWQE6Zqyylzl1MMZGMwmKzqEsmscjHw0dT8tkBiDIHv/PtI3
AW8FI0mOVGJyhf5ZtowCXpErdwnqHM82cH/PXnOvdK6jDT/DUOvq1XVlO500gOYL
93O2D3h1tJrRYmxJksrf97d+CmwRkXQhTjOkr2YnSQk/RkF08DeCoN+ukBiQFOle
tQjQ/bJO32NrmqpWfazgV/2UTAdxPOa+0JXg23g4xuA5+s74rbOaC6IZrcePiMXg
WPGpsZw83k+GIXJLsb3t1GWnzIq/upfOHmjqAnP5QJKl+Oq2ZE+4ekJ6UP9/HEo2
LqCzj4ZxEmmdwgOEEmTkp2I6nt9dEFQQiseTN+1VB6jNi9pv5XGxEts2AniMqNU5
6GFiwjk5RJViPqxKkPQPiUDn1vbr3KJ4Eq/UU+PwTWlFc3PebtLY92/RRkAuNG5A
cy/6hTBQNyI8aXkNabwFdGunWMoMtTe2U8MT3BogAmgwNqBFVfYdWj+T1Q2XwUvk
denJClMPqhqF0r0g70S/3uTJ/C5y9aKdRJ2eFMX11j4im1J9VyTLDd7Af/aGU8mn
ngSSFP9bmnEwKspHoMlYDbfI2+H8JcLSlmG7IEIRfL+NM/2s592HTNUWGsmB0OVD
6IGSqJXixoh4/akuhEP4ya5Iqn7TunPr/EpMGS5cH/F/Yh0066KjfpZu2TbtU+7m
gvggeZwJlvtr7VGRpVnl8kigjiTC6CGdeIF5gTLbPU3RVZnSYzVWdtv0SM1mUov5
C/XDRHN2+wN/dJZBeaHAu2LLHewoXvjd6wY3zbNM6mj2esDqMraNyG1n9Q0emGRw
e6c2qGg3twl4aD3zBX8RKcQkgWUEQVCxA6B30tFL5W0XJcfGVbdcnr0F/lHmE3fc
GdObT0uHMGuLx2zO2Qq9nED1B5j2BevX86TqpAoPshvd+rYp3a9Hs/bpUhaKmfFo
Se5kbcfEEbj0hoyRhVSEN6HC4XS9K0Tur4B+tEfbBGwkvZucJDHHvSl0ZPfnFFb1
gJo+tQIyyu0S5HcSrbr9pxDhM4PieAR49I+WultEkC6K+g/+iAHjQcJNNTpoiEgD
cnw6zUu2eOobLjesTbUo66DgyP6BleFdRdsMAr70LEjDbvbJMWWCFq1iBCrL+0eT
vSaY1Up5UeJQ0SdyrE1YoFrqibI9BuFR+eAXErfKmNi8y1YWcr16FQU2tPNJhMhF
pPLADnVLpxSVV0QUzcPHjqLMuAhghMF2p2CmuF977QJoD0FQ2joUO2bpzCt1ZB1x
EfojplFz6x7t3qD+atkBGLsYTO6RIpmxYVpdjCZCBxQxS0taKuN9K+6L7x8Jj0hk
//cz9qhMV7c+zpddadu2SwcIWEpNM1ijE48N49PV9IzsV2cpC9ycbc7Ou6zEtVoc
Z9nPhXbNxTfwduvwh5GXw05cC/zwk8CvYCUgJN7MGw8rimSNq8yJgs6L5m1/rBk9
tPGi5pyePu1Up+jSfMFbok2ujmi8FDpBRmUYcbXKdDOwCofcdW/WfjW+YBy1KOhA
acirvk7+b9zpG0+nbdJebFuboVlucoHOIQi1A6ul89fbbhmfaFon4T4iBShc32qB
WACEWhI2GmWT0AZ4bz41UgPA0vSU83Fv28VQevT4lLI645xh3uM3NPujQWeHe1rO
4F879AJkuw2kjxxkCHqX0Ejn3VaRonb4byalZOP/UruZdQnbGLJ1/iOlsN9P+mf3
tdHp+PD1ghcHefVIv14Wffb/azk7vMsCsaNa3oKF0uXDl5BANLm5snZPA86L/qyy
bF+nyZtgt/zggwv19BvcecHzitaZ1wx847wb9kKgeJ42elN45C7dGPkgKa3OmP8v
QNAxOf9sAVn7UaCvNUEcVh1AvK4cyhqOn+85ZCqtifiFtXSa058JL+WUJPuXj2n9
OTmJCsu7Otyr/tWWtE6K30jZ04psxkpE3uqoPmtCAKjG6tG2AfpPAdB9zf9/tCzZ
l4vfMhWXqd1gTgANl5LVqy+sEmwAe+xw52UD4o9e0TbLiL7h5wU5+oL0HPa7xMSg
Q/5w4wJBppdNf4i3/2Kvi1xi2lmyeB2JiFcnmeT14xa/v+0/nt9ZruhN50s3fj46
Uk3DSrtZfrS5hfa5MHsMjgNP1bmiNj3+pGOwXg4luOofRypFzVhvr6IAa38nFVCO
WwvqhhBtVMOD0KLigISDmxGnw5k3zLC4eH+yui5OBGooDoF5KIdQifW+xMFnUfTD
f9iyHPaPrclW3T6rzpVRWNB2EkHrP0Ft1UfWvllcLs9bhH+04vBr2aJQwXmKWt9w
u/b9UgtZArKJTfYwW1oM9E3HLUNo0pZuf0KoUYBuIRNXyxrpwYNeY0430BUHbDnR
DUw20YzXHHR0jroY7NAnfLliFv70jGnkyS0ps3D6LsmHimnVfyyS2m4CfqL+1ECc
aSoQ73mk8c5aKYG9CkIGDngPBo/sK5jzjqdokpvFHOM1mYG04C6N9gwlQwLxB/HQ
cSZ90ZQyzHXQsnsenl5Vou4KHo6Kt74w3jaV494TI+FKxxbtkIIU5beMbYQsNTBf
M7wr5QP9eYOl3jUXZ7waQ8M/K8OuREgXy885A/CoL+cSf9cAbq41BCL3s+iv1Rpn
UhrU6mDemAZFI9CbaT3ZJSkFPsuiqaXfZ1GkoudkbWI4zB2nBknsujLJWlbH0DvV
0zgm6D75BDahg1c81yqybiIKAccbSny3IpR+LyPCnAwx+87LxhNAfh8R6rK7Q8VL
rPQjBrMLrIN1X3nHCYFXvEJG5BEzryYlECWBBacR8BoqOtdfEPiJyDtA+PvMysrw
bV48WFQ2bopZRLlY4Jgdh8+bjfgBqXy1LrPQBqz4XudM3wiHhbIJnHSsr/XUacx0
Og1qSlcIaBeFBXlzwAbbXc75nsAgw+NvoIg5BWBNnXrutrOYVcyCDuGF3aYEQrtx
R7M5gpdf0yrf/Ee7PmGuuNs/qCNoFb3o2i3dgEhjHn/uR3IUX1P6Q9cklyj8jukG
e9SA+eUir/PYElW7IUOI6fwvLoxWOBAtpZKcxdcJLtMWcuzqKFftgUaoYaqEGUVs
n9UXkhEgdWqVaGWAKStEE2roq8hRKOaBj/VK8FRdDwU9zQkdHBZjAdFI9JDbvADo
eyYNDi8qvh9K6QC/kIG+hxoJESLxj40dGLEVTjpaQJOpbkaeXLuQHTZdyFWWEDR9
SSUIOYKYWLXJ8WkthmD+7s0wz1bXLKNVhhgUE8+mppvDMj7gNY3b2brsSqc24glR
bQsYhRkJP6RlvN+uVJGSWw287lkr6k51/F/zOCBnVletwvaD/pYPl1YynEC7NVGp
UopTqKJrlH+6/yVlV/vzwC940gcdCsFOf5VdTaQEjnGeNWgXLZzTeP+03wW6Xvig
IPBr+Yh7/c0r0Rn2qnmUuzfQs90PqC9qLf4XpeenRvhciOzehFGHkUnjs+PHSsDr
XxDDljFyBBPkshjtm2qQSf3m23f7E37Mx6qKtKUCtkejCPuV7S3VviwUWZFGx5yl
Yzhfh+yrMDsk0Yg/Ak0E9cPsVRpg2UsFTsBtf8L95X/NbwnSITTzqp7PB0jcinaW
O5QnAU+uCSXNVk8VO+WM0F17j5MXBz89YhA7yHMCD7qReh5WkVYz8t+qDeFBYk09
tx6oB8vTaPkbtghdDVAcKBUEneZayvKFZcbtW8GIJvPNA475EL8EReTwi5XqEbVL
X012dxcGpAa1/b2A8FPo3W2vGEWncH8fZV7zxVEYbPtIBUMxfiid4KTbNR/rd4tJ
+sG9S1HUrvkSAehCYQ2emMAP1C2G4ZvRSUpCSyzKfXDsdZ7iFCLB9qWg+Yu4Aul6
8NUqgZH8pZjRvjWuLPXYZVlabLSmBr9Xz63r4ip0VP6rqUj7PPiAtI33UBtgp7PB
MUnlqOL5R1penupA1UsrKuFSdZriCP8IXuNol8o+ivhZQg6KcR1EAeQmSVkn/X+5
vCrezU9C0MWkbG3hEYZlVlUYKNAWoozEQeHEKSVv+doPu2EUER9D7/hHqTQXcICK
gAwUNksshqdIsXlibtSuOK51qdD87qMwA3RrWAbnb3CuU6U5UYzp3lDNZeqtoQH0
/vcEi5Bv0EKSNzxZC+g2YnoLJ1SkHlTvtUFGtNdtoinS4v3OdMnTxKbcM0xhh7Ak
of97XlPCXWOdDOL+hInC6kga2IoAy42zCg8Uz8CYtz4NSRGTagoJXCvRyHqRJKzk
u1CVXnrxc+q6uA168k3YLZGbGwGvdLN0o6fEA0lVILyorndpW5VW8ArtzlxTC8Rl
gZiJTXa7TttEjAkqoAR14WZf9SVJsW+f9L7fLk82sL/iHr55RuhoX16m7YyvDmXr
yJKtfi94AmeH2FR8JPa4+ms+0IXWAU5EeBT37zLOAq/04fuShSPcvncs/AL57Owc
ywkf2oaF9eb2UNdmETYaddTAeHpyiSC2dhuPCjHjsEBKhXaX6ZZBo0hH/6ZqiBxH
9mjm1nv2Inv66QVpHnDBCdmN983cvP/ywLUPodWLGQ6tVw7ewJZStXDfku8Jo/5H
a0/c/+QWK7+nHdeAOprm0szHX5BCRoXicjdlGscngLeKVXbhoC2S+1H+Nyhdseeo
Q40nNFnVk1/4aJYpcQzpPSkS6PKmrRSIUatRcgdJBQCp4NA5N7m8mkOeK/7nuRvv
Gj36kEaau7iEwvHSwU1hX6c198qcFeELkFuNvanQBVp6YA3Y0UpxiIPkqxx1NBJA
avWEmCf+6CDZ/QL/PIdigo+QDdpzv1B6SQCPM2OK46JtYu2cdAjieLvQbv8XLNld
mGiKbOpXZnnJ4hEYaa2wHJRl1qfPShRa0QppZoZjqSepZijSntJpeSNZb+dUAojP
vPeg+JzmUfW/AYXQQ2ILDdDep9Ed3i7xkf2C9hF93KaxaKGnUU9fqCRR/z0sBWP8
4yFuu95DUrnoVJl/sGbcfYs8w6QRQf3bGz5h9gRh37uQhbXVHqUlNhq2SPn0Nbzk
2UvqJEMciFjBmhVHKw4lX3vaFkRo08toaDFA4+VQeupZ3hBewqUNtK3knYvtjCdm
2f3itbxtbtVqL7OGLx7M8hmc2kSAmYJZ8Mj6je9MmXTFtS8HoNMPy9BzqRR3vJFU
/tZHiPn8B6qkTzR9ON/OmBszvFha9x8MbqhX2gzQ+TA0eheo0dzl3ebYLLfLmcmf
HAlwImWhfVMn55pLKhLuSHpd+W+hU0qssbmAVmi5/mjLXh1FIwB9vyubS2YFguy9
GuhLGOKHksldXCSGb94aZ5RH9d2qAfMniv0DsGvQW8aJtu4G56HVPnnY7hwrUAK2
+fJiyCwfnt7RYrOicimzUTvJKf7JBqq6/92FwNYoc2Jab6Mj9kF3HAx6fvEuLped
nEhlKy26wMlulFvpjVodk8rniJMfjY5gGv9yjAcPMqaZ91ZOWVkbn2b52gt/jF7v
ueih7lqDQP5LqOyE0KRcGVRWvpTVtsjA0cwudqERCxCezjwcL+HA0VwuXgiOoL+R
yXxOb5BkEVRCoXjTwYxsdDsm2ZtP4k0/foVuLBr019hfOcqF1Culk3NTohKHrKiH
vID4TP6YGPAWJ/Tjp2U2X46KB2AjBcHPemg/CR5whsHcnCAd31hHIye0we2PHPkT
eYJjhrUSKO6BvQ3gTQbTJiUvpv1NAfs/wTUCBRzElIWYJAvrWiB/CWsMtb791iU/
Aib7lGRg/dLfJW/hgTST5ywrrpyrnG347ChZsfK0uPZPuUsFMLu3cvMM9CO3NJFY
kb4Js6CokIgkz/xvSSQyXK+c2Mp0OCka3IvYhFUX3EhnUPHZK0ll8g6f2fMSYzIL
AzjcWROlZGQpbWbNUw9ZPYLUC9DFJfyvxTvUNJk7YAy25fi09Y3UEy5+TWDr36O9
A5S0FrbKL6ElKRM8EhvqFOHv1A7YOsZFVfy9TWM7wAdudzvdNABsPvlbbDRjnkU/
Qtzs9ciBS0b7fnMesgHSeFvGXxoSV9myYYW2ykvXViADnv1PeH0gXLK4o1RgX7Aw
TuRNqTXqYllbaYopo56lc/7zeDY6xh5nmi2LLjImtK9oyt0xzIBE51r1H6EGN7JE
7a3HdMILad/ihluaoper0scra8p0C667x2+onmUUciv/mijWkNhRPBVcl0RDO6zs
RGRJ09/qDcoLHWEsv6kWoKHeCzEIVMmT1IDbBWYjH5Rm3uxoYl5jirU6xuYwIMEy
OIpke3NJdZBPYopFU2NDN8YtKXSxzu1O7b10Yah+ViJ0d0UGHikWCdBf8KSpl+Fj
CCVguI0rQlTsRmPRK4KSgHVJc6iTHNBjOHYxvPwfDzjT6q7XjibqiTpc+THpoP7z
TZQdKVA3bRLMTpQqWvO7SobIcavb7p4LxyQkMEEzJflVwHJV/MkbN8ac2mOD5a1f
x4hQG+AehDUD3ktcYBxmqv5USWe9FgPGS4wgZ9vfCEW8vRtxXYCBydz6mQLZAi/L
aK/uxt6tJmAVmIF/kSPHBTl/eeRbk9sCKMwUWyRXUI6KgwimwQg8wKKasSe25i7f
ZDXVPI3Vrj7vux/slvaOytHK1ctWpvX0biwHwyX0shdV3Zprbgbg70KxT6+H5Z92
75sT/6hBi5wpOXqnXcL8LHAQpRbei/JayweZ1knw+zLwN5j0A2s6ryHzlLmJBMWv
M8jrGMWYZtEnGO4ywLym/2nocnGjDCXPcT/2I/5wm1GOML7Mnu6k3+j4C4ATcDGh
6x+648aut8nkmTnDHZshIFH8ZzLr7Ol8aquni0oNUBc/QvxRxPuYnyGkMA7y8Gz/
xtvSxe/OeLbB6Yim4+chjHjMTbW2iJr8xcrRuqZ5S5F4d75cjujxkqm0ZKFfvBW5
vOL2bMUMPdkUrlBycuCbR05X9IQTi87cxhsTu7DCvK2xflTKhqkA7ThAYTrIWRyt
z9pwrsMtP7ign6ExFRcAkEO1FD/HerZH+qsxl/+Lrw3yFggEXnuVh5hTxINBbXdS
qvP0ST1b2iMrKbUN3NkaXfxBXsU0BhWxP9kv6pef6ai5uSENBQsZ3G6qsRk4vHcR
L9L97DJBWyLERPo05vOvA9JHc9St1FnUISA/Cp+uQUtso/D3SAqFeb6bfSE9Xz9K
42MtWJsZMpBDbSN8/WSk2shmKVhQ8CevUOfhy1f8uhGV3t01MoJxrPpJwkHzlEY+
odBbHgYCnEBHSp/VfVxIBAqayG09EQlsAMGziyt8Fe/i3MkzAynCnc9vz+Fkbsep
sCSTUypqANY0mSZHZLIZWw70MWLLYb+fWJo4QDNd74gC/7fj5t9/k3ZIdtYbvhzb
x/Lx0QL27xZdxa/OemVtYnFpGLdSZV8GoVcFzIrj2g7UdoZGcK2g+oFbl4BFP8D0
XzwM+rDOUHumHjOT44ucuNqn7t4O28TW83hTOv1r/7lyJ3iLAV3l9tyNcP+UPIe4
/rBeiecuxYQJXWJUZRRlZgptQfW5JbvT19oKLE5anvS2VSAM+a5foUmdncZSETfj
PAgs1T8ntIth3yU46j3CsW5ohsaebWUZpFGEoOxQ7yW3pcQwyr71TwzoeVC5694N
vzBSqChSMCD60wBu9cKGp89fSNDnxGk6UJNQ/NeO1h5HShkGzJ8IRkCEKd7UEk1I
KVxb3x4/X8JKFCmHWyuLlFibmFeXJvYKtwSdmmG8miGG87S/ai7b1P0MX473NiEz
ERKFXIxymynmeGvNQJh2OxFylNusyhC0KT7zZKAo4DwVABsMBcJ1rNQkglnZax2L
0IAecyxBVYlF3KOxJgIKUn8HRVgHsH3jGbw9ktwy/HP3IqznT9l9GqlwtTXJ/jfk
xHFWBTtgt5uPDGQgq1weotD88g3YCcnkTWOKl3tpMdzuegT+UcoCLqMhANzwtH8k
ySurDQhvprUq66uOv9MEBGsl3TxTq3P0axtoGuT9ZjdFahwQZ6dGCpoQudZEWyqE
ipTv4Hhb96y5u+xilLAIGZU0nFxyY9/FXfsPr/XgbUH+ei5s1CWskAGuGcLFZ55a
Cv3jF0mFNOEx0bdOETK+ceHGVZPk4BOXJ738RfNfimkHpNvgbzDYuyciuiSau5cI
+5iiozxURMkbd82bfA/7Ci8xvIS/drQDqzap22/nvTIFGngwf3Je7gWnXHMDu1kE
lj8muQDGym3MKHQw/PTqazQtpY8wDfUoOBL03YmExAdS5yDZa1Vsn65Ho/A4x5x5
i0LT/dGUI/lY8CGp/VwJdI8ugiqUwRyzA1soOifMH20NBeRBCeBF2rbh7iU0QwkR
+p0K58tbiird4Qh/lNuel9SkqOpRtGPxXjAYSC7PWFhgNFawMuXvr+Fd/jwufvzH
9el3H+dIdHSDkg3Dun/ofh87+5uzYum7e/Q8VW8BoFPNuLGfSbTSBXkm+Ct9SP7v
5NjHcOQkETIhvr/WPUiv5XxXg/gas/T8VtZ320Z08jVajaHQPlQI5ZPGmJ2yDY/k
DlSxa4nKZfy37ZQdyqvcl8XCxpS2nEXriK6byn0BpjS0tAGSuYgS7M+OMWgjtZRA
13vs/dWPFR2SRLkcEPSsinFNABttD6Fc1s7V89gsVYwZokVLPC/J/U3UCGmvJLxw
G1h5vRrIMj7neuwBJFQJ3pQIRqimaHdT6WDelIBtEio/vPcKrMg3ysZllVyIZCgR
EThmcf3IFRsjj0SDICQtaUWxNikv53uWUFr547zTNtBXusgOcTUTnd3RRX9VdUKG
z4g4lVdvxVcpNPYqozmYsfr47aR0XDSZDCkCj3mwgnxv/HM+PBnXn8EFOnQSAMVm
rH1rH+WeIUYKHAZCTIctCRCy3rMkL7puIanKg9gWiuG6DyfQo9lN+pI5P40mpM+c
nqw301WTQKsCwVWsh6oOTMb3jZHvjxKkP8BuOCkAc7qCsNtQ0SdsrKhziBiW3BLf
lS6W4GcbNxDdWF2Fef4jMYD656x2z3ocVeuPDBDwpOytUztmOWZpW6FuAxObdVtX
ogauIWJOauuO0smEiuR6D/RzFVt/eNDsoXExPJNBR/WL58px0oC8LHLVQQytwonI
RfcaoK5BhIH5rvSSfzsEtuXHyHWYZTlNgHyd8aXM+tIaLablCc7MrC7mNaX3x2CX
jqDPZfRdP3w+Vei1ma6rxyMMYl7kTsFg+dM5ZiBqwiJRdUIkSwQ1vEmizkNf3DO+
mwRRsyBW3PRSyA5zW1mAoF2gA2ca8x7jO1riaxlv+hfE5llJ0NJNQ+0pH1uxgFw/
R+Z+A7WN/UVpZobCBQLwC1G062klSHXeTUAIu/NVSfcH1loeIefJzH8urAkNfwod
TgyC7tErJBLCR20QcAP7/jOV0LKeTMxSM1M0D4UxhEGvFnwvMShtxMwQ9mRyIZ/i
+v35fxOAjzwL+pds1nWuMkTJGEJQjr6WamXrJbAHepU3VaXBP+gFhibd8x/bC+Bj
8cHr8OVfefE1tW4gHpbDtpVOyflrs6ckOEk7ASyu67yFE/s+slzhKQZjxSmkiDij
V4VBBEHwXPNxE6NqJ3wdBFId6JX3lmdDAEFyLDjbubNgXsKoP4ruFY/5001OMMb6
Stv6KSTWeOrnd8bun9j2z2zKK8lta+fetFhIOf+4RrSSEMpDQSiEgQZ+8ZN/ll62
w6zcIPkzASEOQlbjLMnJDl7Y+3VP6QFP9X1hcIHhcvEma3RMSmYlfF2mmSSZ95XZ
lqSJuyaim0jHbrDDGgABsK019nC7J9GTznXfjTdYPRbhheqbpccs1BRp26h2vF1q
KdTn96UQNvbCqMACG/a19LvZ1aWCa1QIHiorSj7xQB54XmJ8dKBSUYctvDWVMnvb
W6KfIEnhWHg4Wakk8dWYuksOlmFgu0XvqJYFz0ck5Tc/EDPpSMTx2mDZiknxRFpG
K27brC+FH2PlX6J3ahDNPnAIatitRdtLS88vbJ2+DOCulb8ife7Gsw+BW3qGGAOV
zdVOQl5cE+CznO7h8I2se4zKe4hSLxE4/nOaOqUbmU9/SYvaqEKZaJI84Tpxrv72
2DhdOZgM/oaWM2H/1p8tktPZhLdh5fba16f7L6HpQtHzpxYLu4wZZ0cvVuHGw0yX
wL9MeZnEsSg9f8UYCtyB982wXx3Mnd3eRBAjK9ApR4si4bwwcNObovxAvbQ2izVm
FSqC5MUa4ImeaPl6/4k9W00eTajr2crr3AeolGB1Bu860O910fij5U75SKAkmgRJ
a9OWFDU6kIl1PwBHXx+S2RIoCs2Cev56YfTpb+NIKKei1/CFtDWZeXaO9u+ZIUq+
sqs2KssE2euO0/QOfFz+X6WvQjfIl3uZFDaBfWGi11XQo6wRVmKd1Io9C7Iysncb
7ywBwXtt/AJrZZ5w/VH5tA8jzVMizzQBllsauMz/MZxNwPzbHIm5557yCUjDJb80
TJSy9ST5V74ctnUUbwVhsfclTiYlO0oZHoOol046fixgt5lk16e4jqWzp4mqvhwK
IKI9/LZUXBqo+RWDUweO3s3uw/WbQUCYPurppicjhlF2L9DragRmQ97V5TQjKxTr
vN3DNZwdMlwCwwj7N/+42MtAtT8IJuIriB4KS2p4pxHPhzKKFgb59YgyHXK/cHRZ
8M3vy2xS65U7DrHCfIII9/pnYjR5jQAJrwYLpxr6ngNIoSgFgretSPDqLVqe8g9S
fjtePt/WI/mpjMoUzBunJtJDt79Sa8u10Em/WDzmsjH0rMePeiz+VKiqN4oqih7l
UT6HJ+JGAa3LyaV31r16T63uMpC0kUZZVjgd5bRNpj5rrWm2kpYP9zFeT5sF3Ydd
7BK7mzY+7JwTv5EsL84uA9lMpfAqmjt6HgxfqurSAd8kpQgJ9tRcvDuaorND5W15
rLVOQt/92cXuvmRk8LLMF/Skb5uxaNEtgYZIMMBJDp42AHmVqbybSVUR55w6MSjd
Bjmuovk511iPY7taKuq3ANUCrO7aU3hIP2hW9O+LrCLYDIPWiOFddikikQPuG9V7
97g3PWtW1JHEh/d9dl5d8U3I8/FuhaDZfHiyXXe+sLui/Ais0AMymrb+3/dn+BHB
KrSvvhdO5H6IfwYIGC+dCm7ViXlUQy6y1SzT5VFsk9fr8tRvsyJmxG8rDE8Or4uu
SbY1acrngWsNt1ldyJy0DEKvlruxeFQvQPGuElX8587xhQGRieO7DgxATSl/RAH6
Y2lM0RYdjLM+OAHBJGR0Zgmg33+GbmsTgvbubWj8686uWefiEWQFbVSQ3qratqu6
HWhMnggiUIC9L2gUP6s2wEpBExDX1t38QmBNexrnZPd6dttRmKUGKVbp9P4lQ3Y9
pa+nHFmLT4Sp8jdlYR97mZjIiJT9O8dGAPxGWldZ5g245wOt5UF3oBOR+hUFohQL
jIhsJuEaOtixuXBE6SlkHmKhRUDmpDh14r+2snXMgTh9pSNr0HDQ4Sp7/hzSZVBD
YWbGml/VcOzYYgkiZIFJadvTVf/EUgFHCrveDu73qzLG5MWQUeLAha9S+Z99RTKT
BNTaf+yo1fk/UfYxHNd6+ArUFpLZv2Q3MUAIM2bGLnqVDGIBrJwtqKX67iheZ3cW
nL0QrFeC7Ncn91yPJk7I+/gk4f4KkYLMojBg8ylvKKlEj5J88dAIQDRwYm0K9Jrc
LfMpFVIcGIh0ssvTM2Wd4XeT6hI0eIY5uPWD3NAhAyLXEynaEPrfjQiGOoG01CR6
VYwYaS44daatEhgBW5EIqnEU3wBfVYi4klU30WmbJCqyBovNsmf8+50CPYZuJ87N
MbT40Na6OHrNtuM77VdImCkOEDPdxY39PHwfXZqorNX28DC07y/oCtK7xUQTCKCI
TZ0fpPgFkTSNSvjrtKHNm+5czlGUDOlWeiMNFzNu46pFdsip1yw3YhQdHE8H39hj
xeXZ4TsaJmevL6opcvpUeWb5uRjxiAqiQeTnfmtIKXQzcf+MG55RpP3AIzD9E92a
2W9FBZuxwyjFpoeZ6V/Yf1ltzAZNTclUEQkwp18d22g+ISZzpsr5zhNnEBNzGB6R
ltoW/pC0BfRJhtXzKeN50wuntoXm+uAzEHL/J7HYEDHs0ih/RercwIAfuH2kI/Ms
GQI4MgqRJAlTQJ4Xsq2cu1HpTmDSmMVextD+q5K+2ChzrRlr0MhT20ZV3uI0/r+y
T8LShIrPiGarWEdMO8x3/GP6mYj/Oo2ZO/4CG3oQklaBYlUkmfpXlLBVbZTN8KTL
LD2CBoUpnU2sIbIwpzzR83+fv3la1biaHP2jgvBn/3edWhHgobo9sSmLu7A5hjCO
ntsE1gWTvefHyOwVoHMub3FFyKlgAtH82oE8vkoKEVGEgXcjhgSFjnbXzxz5Czpp
AsC9pBvRjJxFvHYSGCtarTtXQDNHU+/jZmeQ6D3i3fUQ8JyqjNLwthd0lDd+NYBX
Cw0xbxBTxbUslVO+HZpSZLo7M2QnncAv80jh4wBC6Tfat+yQTMMr9RKYYTjEuYKv
+DcHKcetP1Ezo1XtZ+4z7WwCJuQIlf4eR6qJo3SIRkIHT66Whoornbi1NU3d2GrF
c6WRFRBJz/DjBnnfFdJ+qYQji638jerIQGgHCyK6/81Pc9N1if9c4rE8lbQ3zxmL
hVu+MG4rVwzg2aWD//JmiMdl2nFX9dOHOzkrfioTzMt0PoG4Qxu0B0HB7yGmreZN
z7fnRSp8Lgjv2IqEzkCcHrzFRgVKS88E/27VGyhWzpWZ8YcYUx2hZY2L05VS8g2j
CWNc/CkBenTb80yORXDdPGKOBC0SmBw9O1hayTTyvqYO2Wf6BSvwfPRgBOdwmFgZ
pScDE7qT8AYpxOfw7t2WvWqAWSaE6u1ZRX6B7FGglA93B89L+juEG3fE1O/QUOyA
Z+9GPxvBIph8BwZqMfVDjGGK1ldS69UoVdX1xSnf0m7c6k6Ye4vtEHZVncCGosBw
PhntsKGZV5YAL+3jZoFgo/dwwSjKYM3VaDzq1M62p23gQn5cs9BQOr8MvWsrAxaq
cY5aD9RLScTq+7Okjn3pKOHlH7sZmDo+8nPf//MUCUeceKM04KbiXB70un8n5gvx
cPjxehZfv4n1PGV0qv/JP4rDQGHb4mYu+3tbN5n1f+qg5zBZY3vEIMPFFjftOgL9
CBwhcCbsikRR8H3jTjOLZC0gsxE9ikS+CeA89ANB2vEgXjVIOM6D/u8HcQFQNBiH
vItxdyafVT2DqUFkXiLeavgsZ4KwQzJtCBGop36SDaIHaFSbp+qRbAlKdHN9pYSU
DdOMWw+mWoeJbazL2sylrJWCJH+ggHkCjrrWsSyul5nNxtrkwrUIyeKks+sU/BSU
9pDL+WT6/UfFnubdCrNriSTn04X0SDkaDrYgWRgfp6FcmURRUwA9AG1QBPaPqpn2
pbzoLPl6hU2z7qJVgzCVYRjabLo8aZaFEMw9Bn3VHSZPClB2Vf/vELqQ7uLpD7yQ
bANTPUy1ad20txzycdX/mRJx+We6ngiau8TulDn5Z0c5ReL7YVAeJgxGPAUWyqTm
TRYMr0k2jrVH/qJ3cMHcq2GNgu663MB9jVc3C3KZxmra39/FUa3D06ZocUNdrOux
8K1UPL4LrhNIk+p2oBe36YJ+4HkoUehrw3DvzbcD/TA4lsXDUyptr5BdMvMn6kwZ
ihCnEmuGZbrhJsHkotL1+MGKiWt86zj0v6JjObLO+84aNFepsLQ9XpMkfBVhB6hM
RLtWY7etDuienE8cTgiZHe191vHSaLvGwwErk0kfKPcg2gD+RQB0+IRAkICDxemz
fSyk4EkdfJv98NEQA6FmbaD+1WHCqZ8NKfSkdVw/yuD1UFzNi/j3LWRD/by9b819
Ta2ezIRsKoSMNoteUqfVAKkcAK+SsqTtVRuNCfLtK7S6tER96DtWJAh2UQfoNHCL
dpiISLQtR7020MC2xKiiLA3xXW9NNVQCKsJsiGejE/aBFis4shyJ/WLC7xdnexkV
prWwe0oroA1uC1fs3+JQdz+MxB+F1LcKxq0qor0V0tXEcy6pWtJJAyRBNU/6J3D1
1oEKK2ubUnUw+XA14UJ4aunKL30uMWLxg1Bubh2lnDg3tG8h7b6hbEFRvrP3Agvr
N3pogjSkbLY6h+dwyoLD5Z5UrLg3i+Z4+q3n6wbOVFV1ySdpF4jNEOvKzpn1kuO4
9jETmSERncpXoocsQSu72TV1kMp4oSIV60eh085i9tNxvqQ0+hTzKYZmgRFsZ+3k
iMURieOBKNeMDOmse2W7GQ1YFj7tZcBMMxPlRbhjJL82dT8/6COeK4+6QLt0uE/V
fBAh0uPUM8o7d/2YwQD6EiWB1gA75d1ZNJoA9JVmn8MtangJplFMSLvreTertsbh
KS2QkLMWiUiBzR8bhDcAFO379LyOZBxfxBLmlZ1ENHPMGPRtAHi3SI4M3B2+Y7Dp
6NEOu5KZbkUCYwX9m2bNHG8uU2DhlJzpBwb4Cf9wN4vU33HsLA1XI71eprcFQMEK
mSr7mYsbDFEdUZu92foWmPmnSx7gEz9/5hQy8e5AxFhv/mie3Oj7HziOEDYbbnvm
o/ZpGiy5eGrKcshClcFpAebl4V2SYsGyymKghpkfvYBfewpSyeuoAGsEV0pAJHwo
lljlp/LuFnoTHm+jlf3yWZ+LA817PPQTCIo5XRV/bpNqyA5h7INLr3oLaPo0GBU8
o2rHDose/Z2I2lhugocjfEyK2MFsDuz+zt08F8EcBPbYWIzUSRnvdQVBJPxb3tHO
m4p/gVSff6T1X5xxieNA7o822sw/PWXIISiGeAN/Hi1li3UdtDgUn2wRRvkNOXe9
ngS46Wk7oQRkteC/zTXKWGev6++K+83egCnW0Z5mSLRBsrywrpsv5WVsT8AsvAIp
wr2B6NynzS7Rq4HEcpGtfukvmv4ooOGTr1OQCx4kh6pJg49pDicAZ5wvhhv80Wul
lHKpLcfm9JMdJiy7blYiQHirNiw5efFQgbJTMJ13O1kFRdIC6sQgsV5kwAjRrTwc
GoHnfRubObWsTh3cMCFEyu5Ys9mswRDddM8Jb9usdkjs8yC+Uqz74aknLccOtm1R
GlgKsKmQKojDJ0+SffKon1OjKziVyTsqhoH/7f0zkiCihBMt6BoRb+d6u62fQMNi
V8HPAP27bPRftGZZN3M9RfqIs5PySt5rMboz40/MlVtNfnwFajxeVKy0oOUDxNI9
IsRizqluUauI0eajHPiOitKjt1+BI577pvL/Kpt+5D6CybG8pqqPJBcPktqOv35+
xO5LdJioHDvWqCqI6uljNJc4X6FY1sbwuMDpJWyLY6bCdu6kvcYKCA5hhQlQUnV5
CQC/ZWEC4q2XyAFCciH3xQxmpj5yZ8Cv3xZeiCEfRG7YanH/VLsWkD0lqb3SV6tL
KUHxUn51cfw7yp5U32QBfXYEtpG1ovqgAygVvAvHfSbHXvef15D2YITz/n6gV5Ep
rlwyNKgoTKEiZwdUq95xYhyPFm4nPBCZ6FA+XCRhm39uyVpXJouDnlJk86Ogvojn
c5i+md+PvLUkfbTfqY1R3ztOQZ4C+oeu1Xnz55TXcAkWPijELMHs9EPPap6E3UL5
1PYBF27eVTWnfemdjrlq3rZ+LiydVKVmguH7yJBBYRe0SXYLPe2RZhDdmCMBzIbx
RrioBylZ9YMfuk17GEm6XEuRV3DSC4CSYZ47AH0vrXNOEDkh2RmWVvfKKzgapN13
685en/MGPnZbpI4BC/UpxcW1hLFQUEqJ2tJWym2nGV3P2crWjechvl8iMdkFX71O
mmk6ubmega1ArTyIPCLK26QPvAC14brnxNTZ5TJtajZ56qqvMcsNcRO2OBoCdck7
9hnZlzCq4bFFZ1zPMof1B8JyLiVNYnz/wraG8FdCaP0qiLZ52o9P1+tuThvtcRnY
INoul/EytOHM4/Qt5TfIgbE3uec83uNBkv2IC5IehDaH/55WgN4K3ZdHVbCc2FrL
b8FoLboZ0yEVDllWozXAN6iuIVdhNj4J3iqMYwP7CC1vEsw3S/sGf21CU7E1j4IY
/AOfp+lObMk1y5W1LlJ1/wa7/YLO290UHbcQNcrTHqK4DX4fLdyBjIETiaDK4HQg
yCJ7jdNKnDYI+sH98lQdQkBN80+qwKQDk1j8r5Rf0yl6dPzfD0nMT7rjdLBvMRNu
3/WX8hO6s7839XnsUnkHjVzsxjZSR2BTQCcqLkn39BIdI65MvpWijkfwjM5N0uDc
D+c62PfFaO2GFJM8WWewDPSnzT3bFo0SKvefBYzBI/xqSnDP90coKgXH1bqAf6VF
SutLXaZVF+aJ10NFc+g/NCcvzLpOR2Jl9Tidu77ApR1bAPy8AZ0bawpABNJocj4d
DbJHBqH0UDCOReF2Q5u5ZNg/YutEhWy0q1lk0eA0md2GgQ9cmxat2Jpx4qAjBDBU
gk9kan01YCFOiZ0M+LWxsduBFxuwT8AgbjxYwIy9nFcOrDxK5QeIuNLWXFQ3K14o
+V32BKvbRAUqjl733g5tlHF4eSIg9XIROcIr8hZj/+oFriY3jS/+h18uWGgNk7IC
AGnoe0K3rXau+LSkkJn7Z/vm6/AfX1PyrrRgAbwPG3toIkpye+kBs8zaDhOHEej2
L0aPJ+OQrgMdXfl5fenvHCNFSB35jsJZKwK4TC/22IK+PrM8m4L53f7/zq0AaFyP
v5J519QoJaM06THKndtoaMllN317z+LT0B0IuXiKiyNVsLIlWHZjFqeXIjvyg04g
yMjXQRRIbBF+s69h/UluET93/I/qBsrO6CBTZ51sA2yv2SjOn/a7TyB1c/3aJDlL
Ay3cEvvwKV+SWRcE404NgJIomqDfHL5h9yHb4m/MTtGaeIfUvZSYJ3HUipKmskr1
hGmq5Y9m52Sp/WsO6/iKyXOXJSfU3sxPIgn//TWfpsju83Oovw/Ia1JXtlBr0COc
w92BDx7W60u7SIvAzkqq0ZIWE5RdRA7im9agC7VCIrQmkzY9aKfh3/IYrINOy3bM
mnUNiG4LvCQBwFYR5NOemKYLbKRsCVsaI8SDO5FoqT8+ogDaIlvZqvldeuzvIQSE
7T+Jn855vgRIl25kETztW5pmcfJ4gFfpbExmABSbRwJBsCvvhPZMKLxuz/0M0+0J
cFrBe7AzvhDXvXmtZZXGJiLPxxSKMxafNqn05izdA52ercT5jNBTyPzGkKAlK3mt
XVnkD9N8yX4ax5vyF/HqVI28PE0S/ObGtB7YQlCT1f4EWhFn97NFtGb3B4NP64RW
7KwmiqKQZ0Rh+N1UA+iXm/FMlyEzM5PUIRIMqpL7t6ApASlHQbU1y0YIxNYAZijI
q5hfHU2chHm1gxj6H+Siego3tYV+ev0hfkLQVIxuXrvQbT7GmxCzjR+31wB46eOD
48K44yZXeXHD5obi2d8z0pYt/n91m05XteGF6bPpjSWPsuW/LXmg6cvubGZXFP2Z
O6CVzLteLcwo/peKqqZhRo/xdKTYh5JV5VeWnfJFxIM=
`pragma protect end_protected
