`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
KFEXxSR6T38M8S9AgpH9EzKwaBIiEK1SCoQso/SSr5rwyeltKpNeBogOewQIeqiX
PAUwaEd4BMGLpvoXOG384nlybhR6NjyvH0yC9gL4OgxYwxooscQgwKDGLncD88Lt
rY3J7ERybFnReHwcbub9G9dyrQUXFxKz8rm3InPC9xw=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
MEM5K0uGR8lrBxA2YTl9thvSVPtgvHkSt0rFmbbsQrJU2TCfQxwIGqNXzMBXOW3H
ZYOwEwQXXqIDuTtqCg8YWdrrQ0QfX2o9oa5XQBTDlxVzSX4/2hPkks7vvSaqUExW
ZPGQsZvLkh6ecD3F/wtuzSzsLjTv8pElY2D64WhbrBiaHL2U5KHau/DTWDzlC6Ml
vz9fOHYFtM1MWjDsnkvQgLqyb/xZQgdiZxD5B85qmUR+dsN1hrK/BFMBOQ1yERR2
xgvrbLL56KfKg5ErLgRyOV2B3rmlWNDku5oX62guxl+Min5P3yQ4OMoRf4kfnG20
15UMKUxxD2hCw0PXWbe2hxxx2xAAVyjc462ObDPD7vc/tEISP9F0PUZhGVl/n9/Z
v2SpWgYoL1UDT83LfEJ12t9aWFq6AlMN/By6TYuUU23pzmHVqNkxVmRWtG6u1Tm4
9ukI376Zg639lfmQeYIR6rrWtJKmIwDRLHbpW3Ok8TMwBXQVee6Fehp6t8lYfOs3
lnlKJU3oAg77hLt0sTGWvPhXPzzpVfBcqoT484Ok89KHvBRQ02u217uAXBGYJm11
4VbN2bG3fmYiE85h0zohb3rqR26NaymOXddP3qWps1weqBq/rYPFvGkBnIsKvE3E
2rp0Y2rICtOQ5Q7l8gNRdcIpIOZs9uoXfLKtm+XGB27YLLgk9duJ8oswEuhvJTNi
W5BWz6qPdtaiQBYRxZsyGqRNXnZrAM2zrgCYaVItVT3c8H7znLw4Oy9zWdcUSAQa
pOBNscIQI9eElClrFsCaYVZzR3MkI5s4/RR05LVK3hWVKlWnj/YYypZGvBkOXokK
mnMBQ6xUqr+ObuUq5G7OGqtbIVRwUOSU7pt29I/djfy03AisRjGm2DUAdnhKrJak
vj/P7tm9TrBHI8m81nFFAuKgRgPQqy6VUx79N8bpSbI/HEayfBWPfb6y+foyKt2T
ql3jb2jD5Cpn7MA3WafZiF56n/+Q3vHJPPw7D7GBcAJzhUwJOIXADM/tzdXaBYO1
nWwf8kiLAHqTxhn8KJgYeqEgqdS+4IdbH50wTn8KTsnAc5RMNqakSItUnv8KLnZS
ZqP5kbGZc1JSXJ/k+gOnk6A9sNHzAkNcd0MOTn9c+q+Mfcey2fPloDRkum/hk3nd
nDCOTxKQZrB6+foxD3cVHhXRli0DwuIfT9WPCrJ+ru4ycs37n8Wl1UFZgYORRLo7
a7V0h6Uz9f0lb2o/j51VAxbN22F73uQoymo2ErG5Y0cpeV3k1/GnR/1EdCNKFBQr
BhiVbFI3nHSB/9uPfaWBvjIpadXZ97ebiOP7VpaP6SIAVsv16yjnMdIi9oqfoQ6u
+Wrs4Gq52vzGFjUtuKsXik4gVM2tLmm1hSHL42Y9NP9wZJ7uGj1QHRyHh2r+Pxq2
wSt9dHwRuL7mg5OsLhX5vGBnT9fjKoz3wEpKyz1dnbIv6GvpToUFJXjU+nZfRY45
Ofx4DEORCl7GcxjvZmlTq1SMrizQyht/FeVH18dBRRBWkMIM441qqqLIignCpW0H
7UJ2f1NgMhR7Zf8vASIfzLD7sSG0ZY5gGix4XHRGNdQFGiRnOaibaK+0QFXue1hx
uco2AxhxGYQDt3RRMdozC2rQXD4a7B/8vjvr6FuFyPZulpUZdV4qMKHJgc0p56nR
5i1id+3yFbe6E9u6oZijgx3ydT216pCc1pRrG+aUtFj5pbZzEXjcvHzDyJUJAxE7
FqDwfaADXHhCCqkm7Y9u4jqQ13+ZeFACzYpjRDwXPu9h61uKQy10G88AWslp40CY
5MSQbbRwrP0XytddbclRBX0taT4ZsMg7EAJU8NSbxAXLi/JsWxr4YnWNCKKZZN7l
fReDcTmwKLUN5jP9ZLUfo8yQ7f/mG2hA8cWer0mF7HTEgczPm3tlqITykWTblHiI
PFZG9vwnPB1l+1HyOveDHF73d2MH6vzBJzEzkIJFwgPtvn0yiPmHryNWFz7lZzDb
zlzi91l+hfTyj4uKxDq8h0LZ8j4wWLpRJR5h0w7p2CVVeRrjXdKpFJIEdkvMIHLa
dRES7S18J35g+AU5Ja72fBt5W4SCSLOSez2+onujuSh7AKnHOMWdfBIO0Ehv/pYv
SC2R0LWWF0e8byzLRVZMLed89f3MoNhEoyzJEzhFjxrpsMQ78cy4KuA/k7kX7Cr5
u4L4A5igdMye+c4ZksyrZc8c1DGmExV57RgzQea8QHKVeamtKQdYvLmq4C6yRBRZ
xq4Wcj4VMVp1LMT3HyI+SjIDyQN4ptsIQr2WBNycilJtpzJ3CWfUxOYK8BeaOk1T
A1WdUJ0toxb9N/NZjtbIzY8hTAqTwAYcjZpiXK0K9l8CsLxsKRM/x74UibGvK1iY
tRyayKuYVfojk7JJJSG0IIb2r/GIPyZ9SMFibX67PETVWR/SmI8wRnyCo/F4v35S
St97QYWtQ/a7IhgRtTR7ENumb73+n7ul3v3MhdOfxwUox6BZH6HRc5tvSEs6qcBg
yheuJCEnaqXQo55+2+5qWQecJhq6aYh9IYbK1TBCOaMie5LwXz5DaTXfWbBKIwTr
snMy9593JXim0muL0cTZAK3ASGRxeLm33+Leh+X1MPV55eNhuWs6iTDI1bCwXON3
oSv5JKKmaNIET0e42L+FlRw87ILhek3f1bk2SczFx2HYXIztMKkix1Yjex7FUFoj
5sdNPmFCTjYBz/Ltva6IcAXE14RWtCC47+9Ofa980Me85j4r15mKj8mHovGlUZNa
19m41kB/DRoRbZu47K/fX84/MlCr3INNEJ/XZBEGEYFrQBvlitRFaT8K6aUcOw4b
5Ordb0hY+aF75oVqcWvuCuc6ltTn6d+KQjtyQvBJ4eNAVK6z6NriqFDjadL6UBMh
mu0IGZr9N7LXNIVlm5iTYeQV0HGH8HXiZ46HCNWoN9aT6TP1h1mwTy/R7+Nvlhzy
3Yqdm6/lL8TI9HkU1UKaeCZUEaPBpYfgl5JjGALo/p/5oAr4tiZpDb00ljvHmuCc
fdcINU+AeCrxnfV9zpMpiYHkT9z+5nTC52E1dYKY5C60mMm5hrZugdNhyFHEDKu/
N1BGV93M5L3Rkz2fX2ubDCcNhCiOu1Hcg/kPnlqd5PAAbiPhPJJPfNWj22QQDH7N
hNyqFPHaWArWb7sCIY+n3T3pUFlXj0qKQ0ljBuOQUaMe+qxfd2AV0uq3rIKjWGqX
ZXPx/lxSmzW5KR5ZU7V568BFWn9vjgSDh5tUU3WPBPYPVUvKVpiwFib9oT5I0kFz
znS3g6uDcziY8rHOozoxSK5eTQ/mVvXV1FTAnKLecaXiD6/DM84lt4hB1Bng/KiH
8KspuZGHF6dnunOhKJNKeHbxqhxYbNf0a0IeangvyKuRPP37QfjSASjDrfsr+ZJM
/+EyHBCrmGMeBgItaGTifODq9EhtpgwC+z9NEHL5z8cAXf01kz0FJrNHzjJmcggR
6bsMgXqaPIxhEUOoBvbXb4omYXp7v0sD7+SIuH7hGf4L3OfJIkeuxjzVEFDj246K
bOKNTcMBXk7zjOJkh7yMAtQ14AwDnLfbSQs0WWXbTGB0TPFz4yvjqk6cH3EhSunX
Kx7/5KVhP9ey5j57xnLi6jpf6VjH/mTQdy8pAe5+GZIwCze51GtGihlTp2RWfsGA
LeTb3mmQ7vpvPAJdWeibbUbF/u5Bz9gjwwGhJYv58M/VB5rN9Xmkc8l4obyaDnfH
t/BxFymQUnPq1it/CuWftt/stv6a7qkMGSZWAZu4T076GoWViGHV5T59qJLfrLHy
NjPjcLVHcbGW4MA2mwc8DkIAXsg1A5VfzIDdqOa4LwtI+ZFSEhzkfkjFxWU0yM1o
0JFvDqjD/31MUbJ+7sMyTDeiPON+nMBK2UyFVUPeFp6l8bLI8MwlfQPzxaze6m5f
6nixSevJDBIPnQC4I1EYt5KMKwtZ3YrZ/j3E7C6hurn9HUqjwJD2FcizgHKz2eoS
fQeHjtmAUpQeADo6PLf0L7MWkf7LQ3/Zqf/+ItC7RR81+sPUvPAXapXyvPXMapPe
wckJl7MCvLdm6tXLFCeJTRg8QzeH/a6RV+mpM+AMvUt/b8hMzaPaPYjNG6PefYI6
YPzrgGd6HZnL7hF8+6SW8kZ7m7xHyXB7dtmJlgtzkmdClGOMuhc3ZsB5QYGRZPrx
XYGiwfj1iZ9Kf4KWflvmX3DcIfjXjjxN7YbiQsLG14iQwuJRUCK6kon1dG8PCWc4
GQ5VhPLE+XrUeg3ucUIHtRYAhcH8nS/m9agEfX25zaEfP10wPh+r4PWYm2FBqUHJ
igj8LdCWjfEB2t9qK01Sbv7t9aaoO7eMDRrhD9H7skZmWsezcNXy8WX1DfaOj0e4
t5wB0GkwyogUqFDXhbkQgQ0dT4U2tO9y2TOSibHwsZi4xchdYu7Q9slFbRSXvXnk
1+CCBtENZRlnP6sL8wb2UUKA2lLALxXZhvhQ0bm5jaOaPxMEpQlNhOUblYByuMgI
R/yEgkFM0EV04rZghgr38uAwS/dAEfUd1a3MlYM8KV1Ky7PXmJsUjkayzmfgo1SM
1wboUoAJEg1k0bg2v16caPgOSIVYB4HIT4OvPs7rdpFQaCieWze4bJBioJAgoDbX
JLpNIF+lXWl5xWyQYXWzflC8Oc2hHFQeVqpIswEi2xFPk8YJHSCwdNSlHPDGmSbl
t1Nwk+RIxZKJFxmb8H2sIRB5SxhphLSktWz/XsOzNlQiyGSPeLBThHCRDENsYRS4
t9wbhufa6XbausL6/DA8tddTJbHk8tMV2WxFIvtgbEjv6+8mdvgWipV9eHJhLesx
Z692VR/qyaJNBoQCWBVXpOTWKKkA1dMN4hc6DBsEJQLJKeND3GlxIagQymssmbk7
6+EoquRITcOf7QmRhRNk2qaiZLenCh2PxLaotj0g3lxFTueuH5GHVJwMSp6ENFMV
uIMWBHtyvCvoJ2lDaoB0zSK7AEMa8JFXnLDsxqWErY+zEFiAntxtijkU5OYBx+bc
avoNWvAfHuKFfmKma5Lx5rVXFN2/6gHp3ft/CaaNKEzumQq75gYHTXmVocoBUnpr
VmgWFFZdfY4FyuTY5v51xNnmhOEAQD7oQ3W8k+nJE3krvgxjOzOwER/nrpYqPm6p
4OVygDZzv2tdXz6d9RBi5hKdyvRJWcz2hqywJaPxqf4/VuWPgO5hCkUZwQqvUUeh
cpfTKUhKRFqi7FBZohan+rLbCd3iKFujagZ/ml8vQaghor+qiHxkzpgFYu09u+Ff
8h3mgiNkAIGZuAeqqRNHUlC5pK6JQuTdyGJphoCAfoqx89s0ZDu/RhIr8/7Xr9Et
j2KbWY7lRH0JvtVO3/NpmFhHhipZRkjAiEr2y4PQvzE4CRifm6kl6njj+Wm9FUkY
kpF+k4oQJSrsUrZige8U45f6YzMqzpjl4DtFvQAkjR9Y9LQO5TJyYCoir4fJnM42
kw+mWrh1eWCqV8roIVA1yIiihSvxoKEZypouc77kn1jzmF+UoNxeYuYbP3bd0jUA
UuYEDoiXwJ5JOXfgepdWymCAN4XY4m+a/0xLrJ/HgppB+YXmKQgKG3hTsBtu4p3z
CK6RgeHIbXD0rbODU9aNJNyMENUNfYLy4vP2JsU8qUqtFyanWZr2AaFhPXsEcuaj
LBNNLciImeuhFHjqbsxpVCXHWHQ9ryRzAAVvMDk1H4BZcxrtZpJgQ0poB/wYa/x5
UcpmeFvvRvxi72duFNyJAMJyPuyo+xPEUStLJ+BRFJD2FtD3V+jRMQ40Pfe0RoP2
lFmfJKQGmAT6++0Ke5nmKm/zD++B5Rjdv49PBeAYFMfReg6exLw7bjws1y7zcxGl
nQzc4EKV5ARPwb7fVR+hsCFohZ4E5fT2hKpfkI+C7i6BhrQgiRmOS9ZLO8JCBEWc
ln9n6i+ocxR2AOoNDhnWEGxEUAEZzWBp4fyDY6uj1bqByPV8I4N7AQ2nqtw+FQr8
ZjdNdSqGoE5sLC79/BNUcjVlbojRAWcS8kS/7GRKoVp5ZYtV3l9F6fU2gfsa0gEt
31vWave0YZXxjBciXAtoBHr85qr4Hx+CcUzA58I9hSfhRnEEtxIM5ixe0c8eCEoo
xbPRilpfnqyCc5PODlCJkz1ev6x4IjyIUOiu2CODN1KcslfrsXqLWxklW5f9vfs9
K0NzxUvGrxNXpwWZ4g4YCLOZR3bYelcRuprdIHm4wuVbv/ld0mYsmR3oOXZR1Icw
MyabYKKxZAl4t1+/VaFibFwzUkmu5jElU9ZB5TBcyG2nTKvdNCc+egNkDG2fV9/I
YR1o/Yq6AICzlR6N4Z5uHeVgEnVGTsDIzfBCWB6r/0WkEqEDR3BDKxaig6Qk2C+P
ki/KeMEUp+gY6EuD1urpOVuCslGGe3E/wjtzwYNZrb8osuMqx4BrNr7y6hMHEgAp
g2PvSgpTi7bkawIOpMDx1CP5RxWSHNqZ9dTJlJqU2J/SgfH2cLsBXatKxYPXfXwz
0kor1mN33NU1941M2J7D2+0RLMXT4VCXwBe51hBrXRG4uNo6TqeqtbB8xwnFB23n
PLE8aAIjL+O7lUpQdT/6DEtibagYIzN5tb8MAStYe9JeCTsC/24XyJNvSTkVMxnK
OrzaT+7pscrWtmG2p7VYiKnP5nrtr8lFEIFzZ4sOwQXh7m3rd2wv/8rU5iM2k+Od
yy+3mWgo1i0GOhbSfOKun/4VmSyyFlUbUvnSdX+YoCbRJUVdTFk+ITTKpFIph8/G
D9zuTXXHWB2huoeh4kp5Nicl9yp5aAKPRW4Xxi92EiocJeae4jjBN1WsDqybKGQH
zBqnUBb6YYXRTuO1xqS1fpOkyryxsb4GJEl+GX9Jvp0nuc6eLYg7GHTeR6s5wfl7
PLZA42vP+LUtimhQvQY86uHV0KnY9O66zGTDlA19GYReJtNpNY23IQJb/E8ZpSXu
6FC85UjdWwnCpWSSt3uar0rRnwWIBsn06kjn3lilF1RAaF7gnizsXxpZLYBgN/1U
2/6vFyTLKFci9dQn8++ryYEwhuV1ypXCLtrt+NJLxTQ6Erdf+9LouVaYY/Ob8Jw1
k1SD2d1L8i5FXVkuguwWLTiE6yh68XAtyRLByVwDHUygWtxHlxW863sSavE+/i47
36xoP+WYD2snzmZCR2AmAvhkX19Q4sHcYCv/yv2JNlbtYCsQatJvE2F5GjiIqoeN
uDrItc8+TqHIihEOXV95/yMQr3PHlsS4Ub+G+0WN144p1ezedvpLeyUUKJ8Wpbxf
4s1Pfr6+UcGmAcgOibE+2C32I6wZjswCRYEofWv4GBoFUviJQDa1fzt1ckT782Oh
xKvfyfol3wy0zBXTuvtsUWcVwUYu0XVTX0ZXxGFGD8jhRWNFyojTBw0sYgGWkxCV
TkIl299/Nkl1kadEnCxuS2xKE8u2T2OBNDFLb+C8FXCgf/IHaWG62aVUgLwFUmFj
e3EAzqeK6JYVFXounoKbXURqkcPRhU1/RYpyoWVteDgU/yG2XnA+X7NaR3+L97Yf
8kbfLUAICFZIeuYpg85sVspWA6twTWkboimKQK6+QOn4TzIE/7k3Jpr/lm+f8xz+
7BxO3GLB5pnvpKe6WY9aBHBOWyEKga+nABrMEs9RoDf8XK87mke2S/+d7pxQ2/Tj
FM5AV5QCy5EntAfL0uiNaF6CgbNNZGL1Q/IYkaLoSNwj5T58LPNeIIySCXdQeLnh
ctEMv/uAIpZ/bB9f+ZQeduNDBht+ygnFeFtNyDsIVxBvb0/derjuXtG/jsPRKCuO
JuA3QRafwRqm2URGHM1pGVPdjX5UIl/M2n4htIYItlX0ZDDt5bx5M1zM3ilTkOvM
wsbysgc919F0yI0xG/JqXVtPrK/1eTbw81FVG/Ga+DrUNO4u3h0MToQe5PcKLdB7
+cDKStuDKQUdSStvaUUbhp2XXWCF6u9EFks0wrCBfYUymKGk5235vDGXFFNCLd8+
vyTviWZAX9+1yxPIiXkI/dvfQMcZDyfqcz/cdAzOBdjTxE2g9cTRvUowD+DVwnVz
wD9RdHwYcgXcs5p+oEamuu1z1U36KE6NeWm+OEhM4pUuicTYRuEkvEJ+rZUgZ9rE
Xa2NBG/zTDmnk/NItub6Vx9aMY6btgQfkNcjXY664fphM6zRJm+beQd4MEruAFn3
8nsJKAsHZczwxqJgecOdoGMa44J0gJCEwua9Yu/wcir2QWMkIOlezXghtbM6a35e
i7ajqsyBfBkwYz58cEFAERNYfZnNTvR6LHVtBbhPA3jwii1W+qKSQ4TCbCftfRWu
eyhLVx+S0iT/hI3vnNka8AOMnZ26btG0Vjfu6cVkQ+WheB0/JI9UngHn480cbfEm
cbvfIShAsmXECgNA7os3kQjU2iMsyrdJmrsAaLjKt+iWVKkUwWcU+xGcGtZRogSP
rOy98pP1ExAnN2qLS/Lk/SK5GT78ku6Z6EAPf3boSetFB5QSGHjaIjgCbG21/3AJ
YPMSUHhcMPOyRoZS9cml+qzM+JQF95O+lvgwqPypyQ0W+Ogd8uA2uFgE1hplT8cK
1RqdVbc1YybaaIKxcYT4K9cE7R1bzeMlzSiZWe/9AC5//0DmRpvJUjIdxZUlp0eU
ibv7hQ4ND0WCwZXa3PrXna2/DG2j8jZ6AKTQkVEzkJJuMRHg5JF28lWDaaONJU/N
vnG+MGtxQRl7Y/IgkNeAeqQ7KtR2bcE1Nt5WO30P05vQemBg3E4fuIqNYXQfR1tE
32TvdMwGRM0lLJ1TMl88s/f9HfGUFri+tyn2l9/hdOF5sh3bqyyn0KS9ZwfxwxAu
71fusJa963niEC29PEtPvDtlMBheW/8WMD7W7GkbMefjK5+xxxkJl//OAgAd5dXq
1VQdpk5WDlEGQHp7MPQFzHx56smxbIJOJuCZm5yEkAfU44PuwZv1BRro5DvtEPTZ
ckEj79+RUgwapMDYGOqGDc2yNo/co+aYWpWXZaMQzc85/gDq0G91GyQzj6GvDC2o
pmGATBnIxDPUwjrYcQb+NBMjfssFwii6mWk+RHOI4J1z3Mm/Sxh2g5WE0sZJE5GB
n11nVxOPxR9kAg77C1iHY8mDI+bbe3LbvpUiaBqN8pw5zXsKGdompkWvTRmjGybM
wAoMKqJUCtviOnWIbw7ouyfrOx0XFNo2UWaqpKH+zNxCXugI+JjDcthPfBjJVc1q
V9i1fvx3fvh7IuPw9Sc+tYYF3eAnV8lEaCi5UbR1ZPYovmxEwbBjDCm22y+IzXQ5
1MGpTj+r95sgIhz8h+rj6giD0WZrZu6e9DbEhDlq6mVSrKLzrCPjjkKcQlsmVG/W
5WxGEaY7V3Kn0ZTrmik//Uwark1LyGCWMDMVyp/RH6zxZxcesDaQ+A92fcv2GdNK
H/EmOG8JhCYppoa+n1fImkSNzXOAvghubWNOe2cc3zcN6Adi+mn0ma+gvp8Uva2z
WTHva3rvoQeKeAgc3sShEJQhBxMdT6H1ZgaEEpYh6pejcz9cKc8MOjAp2BJFNCNx
W+N47GbEilil+AfjodVXZTMrrVUI81CD5uboifGznhu7qio04ip9BWAmzFtnftvs
Rp4PirEyrBi0lsBMPbWQKLQGlx4Ih5EyuKxvx3Ivz2lafuVSzYH9bdqtE7YUIENl
y/Ip/T6+sIDGs7SGbL1qKP4KI5R8KpEliSmF7EZ99Zx9z7YVDO7iGAMkg0x/bHUr
VHSqKJ2kxzuiuEjpDEEWX/ghwd73ZihCFdkYapxCtLe1X0XRylZVRXfY+GpSJI1L
o3l+uDTp41oJQyGJFkDiJYWp2317g3cMd7wT/fFRRrP2DwTmvc1ixEmQ2FaCD0h/
XbVAiwUsIJ23zi97QkuYPkHyrC8ALqG286skwOTqzuVDHZTHqzqazRHh3d+0d2Q8
llk4+xZfXTtRh2nRw1pUjdC15j8BEyJoY+FJTEfNfm0EAnTeJQGWfHHcZf7acYgc
opx3wcoHsoaVjoSLP+b/W6bU5m9LwHKZ1PvjcUXdkxqchMzP21iqhB8VETkNRtIv
5FDB7EL9dgHYLEfvyEQlp4PSbwo2xCgQFKDAcwCohMuiz4Tl3x4nkII219Wr0Xnn
Hv2fuDZo3/F16BqwXkAo1MNo6Q2OMkk9RVkdV7dRcPteaHmBf6WpkcVOpt8O88dL
r/ou6fdYnsnU3SP5RmiqzJoE4/NPsLXSnw1cWnsL9+og37K3XhYoCRvwsluayfed
Si+zRr8NTlWdkZkwbQ2qZdjmtbcLm67p35RcB7z8eO9obOEQMnt5Ql3dbu/d3rZU
TOH3o7g9jsczn9EjnSZBMEUi4vmxJeLVu1eINbGRBggm1mc3pCi0/ZfyrtjhGga1
/ABvXhaNUq58M1RbuqwbWffxTwUj5q75b1APh6VZEbfYvewM/pgdQ4ucti344Yau
9ocqntntWwLxHsKVukXZwmNGp6l2iRArJiUXNmoNJ7ojSguBDtrcOV8T5d48GtQb
nohX+a4r6El4moDeNJrN/GE9qULkUX3yaO+uUgFjrZJ3Fp51UDJ8xq01/q0aru0V
D4vkXt06TEY4lmmkCJc+ZSL1oo8vL9gHMq0/Q3r61kISLCcX4Vhfb3DNkOgliJgB
vl7NOU/NQLlELszs3dDLeA1IpJKihC+gwwe2Ur3ETiQFh0Mf5PqiJkpB9V0eRisx
wCmUa53DGCp76rQXULzuY45ddDTmaH6PrOL8TDVySCbfQ1Evt0eEZrD+1lVavwXR
621QPlZtjtcVUk0kHNsTS+rzGa38bSom4zYQ6bpXyfMzlyBtbjeWHQdpxdOXs2hb
pZdDhs/EWPfGVyYKzUSlwAaUGwdg9lu+qpaKwH4Ld7djP9TGbMNOaCV3NLFeob6h
jSOo1ppw6aj5+fRY4hjDxyt8eiDGnXp8/kOV2E08/NnY9WcwNxMVDN5Me7yLJdY8
G7/woJl205BYudCuKK3sBqwMIxypB7vvoueL6vVvevD5MhrKtCjmBG42BgOo+C0O
5SkgVxf6jWPScNTdWeev+fFvD86IbMtVUtkaj+Mwc49MmdQht872hjtSobiasMrN
JnEEoAfuJOWSQEKiYfP2f+UBK+MMQsohjUDTrZ/tCtpIwYNELXx2QPa1hAs3nUI9
lQg5w7kOLeQQ7Pog1OgvTOO/pc9+nkt9yuuxqJ2q+JmYcNf0PHivrbUafzpd8S4R
j41FPe/sXTv+Z1AizpOTDco53BYatJW0XRqpdYqubWXonjsXKBkqlDFIrJES5pJb
QTlzpilSeBke2e22a0kAYrL7azFyxuFTJHj2mOalXr+NTvX8NfRMrBV7ke5Wjo4+
8qGxuZJt3aHWt+NY8s+2RH7X9BeXzBg0qpzTLQjVPheT+6hITy5b0Q/WRguJB391
4MKLKU40qoPH6nbijyHe0zHJygltp00GCntImkn2Z9wq9ukJFypqteMUMh3cQTbx
7CqQi97GHpKYiSNWxZZyKntvxiaf2BDzKi5+nnDlYhY=
`pragma protect end_protected
