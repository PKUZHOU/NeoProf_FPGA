// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
UiE0Xueb36RW/2dmMt3ZbuvEe0m+wz5tyTkeDZZbtouya5oZUW6jrBLOwcfcCKRJ
Frok+DABqdgytQDW7bjT/YQzkoah0nT7fFC8hBacjROBBq/SCSFNdUGgv5cXHDqw
u9Ib4eVUQJDIUFY2afFiTEY66WdjTkF1OJ18T5K3L1U=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 25728 )
`pragma protect data_block
fVHZkZWigxD+iJCHftmNJJZWE1zrTGUed0eO2OEvBIXOEL5olwNEBTAYcW0U038k
0wCOjl6Uk3vEP90XKoshjcg0ppbTySsdkMdhx+nGeTD5Ty4kU9fYtV07+Pkv8wbv
Cz4p8qByCOMRSSUlTI5tEmNmpwU1vWFxyaYEHUgiOeIrDIVI5l1kJfAg8KD0gb6+
x0hXYIHCYVFr9b0acLmP8pL0wjMxjDZ8+CJdQxKESkjUsAO60IAPO5EVH7oDiaaF
VpeebLDWfCRJBAa0o8/RjYSSLBL5qVfQ9SL6ULc3RBH6h71PTinZnIWxP2UrDRUQ
tU7np3E4iXX6hU050YwWAwefPya3IWjXOT+W7kpBaB5mcX/Pb+l40xeUv9qhV9p2
ftT6bqPXIeGv7w6AjYwcn4vWzbZQ7IpO0391ZKrg5WLdDn07LgPvKvc3yMTihymq
9kUfRkdGlq9Ud0fCHRmbJj7LwEUbVKdUFt89B6JC0Hcm4axRnvjqHgcXFgZ8Qr/W
WvbBQtq+yMP5ozDknVQebJHiTYKBHRmtlU3hTihgQrVEfDkAkboed3+hM28HYDRV
6xWN8+Wzo45/bHNDdfK7UYmk4s4rGemYpJzJw7y1JvlLhziJXu2S+ICNz8giARNO
KFWWAgXZeCesmIxHNH4DjM55DzIheaSittkQfbcYek785gPdBER49ChfiMIdbtMF
NFpTRI5RU5qJQVRO9V69zqzvlzYDE3XGXulUzMJHtzDmsmpCLt9lhIZt/LRViDeI
+ZQywlh3jF8UR/L69TGJeo06+r5WUwu6QkwtDUeebPD7Znx0a6XfpyBRyGi2surZ
WF+80XuLewojsgQmsQiSGlv8dzNCfuzhIM1gWVHPxuqGAHPSz6rwq6/FWnk4IPIL
Qpue4dltBFsxc8zCXTU0NW6G204kO4AfxrdVZuviaZb0Mg3gJEYdg0EZw6sO/5tL
OV2CQDaS+o/Bn05SNhlDAI7QeGJuzRg9GaF1xRJ0yZ1iGSmIavXvpuwN3mOe/rOf
NTqjxvsLhywIvFqjKuReWpfX/kv4yZgNsrDEppzd0V+dlr8s0MLvK23Vot3i/Z6k
S+yJeOs7PBF3E7Bd39nFWIkUo8atLCD5YMx8eg0WCgecB8Hwa/MIP8VYkRNMOaTv
+ZfdkvZzyDmkTu+Bah3Jw41x3paNywirq+acyrGTfMQqrMI0BzKKM1/nb0ZHRqZ9
vmX+qGI2lo0GGohW9RHro+wXnSIeAQW7nC7qZaKEh73ZT67B2JUET7Is0hxkf5KY
CKqzdw63yT4Rn+2dwvn5toKLrVYx1URuH9++bhlFwADsUBBpu+COj4VGUwn1TD2/
8tCdLOhu1VoLxNWsYxAPlYOVpuMlmqh6YNilqPCiHKPZBujFBJyrJAdwOSVLjlPM
CkxQ4YOW6TzWY47Pn3GKNrp1Uq2GTT+qDp4dRbYXmdiH65vLDr6cCXkyK70TkcyX
ECNy7X5RH4/eAxTYVd9ODTU0HWgUysBgDrzxgCArlMCOtO0sDaze4eciaELEn1Ly
FOsiG4izAVyrbgeh8ZGPAF+Lo6f4y/YhZrP1E0XsRv56R+zxZz+1XbCubBre6jnc
2y4G8JahYrdR5Qe1m0RqQ55gRApNUQJ/hzh8QWeGtyL1wiJJBbDWtQSku8Xxak7v
RPHlRoh8ZxZQ7Wgb8ZBTOUsjEyoeI140tc9ZZlGqWVujlNGSCKXO2BRdiyiNGl+u
srsQVO/ayLnMdL9qDPgHgER3YqBkDMWa7r9MVJxPaE/iLTUJVPDmjuBTNTPZMTnH
Cwzf/tqOHXOmNktMqQ2ukluUhlv+fGvePkjvRy4AeKcNMRHSnxlDxCuDHGzt7MiV
ghHIlcc7qNwxKE7kPh9tFo7BzQIi8Kw3CaSdirw8uZ3/BwK9cEeklvry8HK0+tp/
qI8v9oE/cN+GrDez9UvAuyuNYky21xI9vEXJ+0qIw4tYq11lkhmuSibu795ukhp5
3ibx6x9GM2HEMO02oqKJINHuHgVO+1w9+caGBXp63F+Xa1u1mMtXe2N5zAwVMBtn
84n+H2yYDWReP9cWP9c+Ya/iz50f5eC6mmUifF6z+B8Ts7qeMH1qNZf2wW225VYi
vSTQzWH0i0vpIJ3ewCbpmbacgOCX+K6HoJOL3GOPoJol+Yn3B9cJkHK2Q1WcT46y
AzLC89tx/Y/JuLWRZfUipTp38M1RlchXnHqFAXOv1elQwy3U+MlpBch4aXyNSoBE
osq43JGw0r2/jzKyIOwYGBiVUZ3pdX9UppWs9BOj5MAuV05phG/TA+KSFySPAe9q
nUkAbg1LKXYYZPkpE4hc+3sdAzRGrRAkAsYXQlrq39XokV/Q56ljEJKCWdRLuwLQ
puXxF3sBjhcpQ1sBVBHcpZnNNDGBxR/nohoY3E2Kol+jqYZ23/cNQXW0RWCXjIU7
XMhdSYxPSgLA12LXBFvIv9LzSum8OVrdo3x5xte/bRq9lxyPsnVr08wGOIVtEXn1
eZQkpykIY6DQm6LbKfNpceBV3Wcxjrxqs9uDO1YIOcAvVk89ft+7ngWrdhIrT1KQ
UTFN/YxpHFQPjwTtIOq7wJ0bd1zK9uaz/T7uYe1FwWZgIcxbQU1bwbnnXt9NELpK
b374VLcKW4iL3W1Iq/7iwH89/cvgDlIt8nk5fKzI3ZY6i97EHGbOvM+j6n73O0zf
9ZSorOdeBXtEiIaKBtGMqBLj/AljXsACQ8RjrjmQrzHYvYmbFFRTpWxEdYxVPwsM
xauXeG/hwgcRFMNb1wekxZ4/qFtnoiWMlL2YCxyZcf8Iwf4wAb/6O7tPE+pIu2pC
bQc/hKl7X09mcMbzYpCdP8P/zMVGJla+Ihvr6U2L3irqKaZz07XiacbqTxKsHmOS
yMi9iGj9qnNyz95RessMCa9tvs/Xf8PEiiuAgGoaSO1sf+fFCGYYpPBimrhwxDkr
2GRkkciwivlUjT9mnqfNv1W/fso5OO0GYAn+5/xI2lzBklixAq/Q0SKUIyUR29m+
7OUSaDvNL3KFfEOjVtPlKuU0kDA/O7/e5J5Kk5va1qVe4K08fzYBuW8nu4oD/3iJ
H5NjZfx+wazAtdAw1N3pae7Tr4jxHNfYpBlZ3nbEwmh2nRHwePORbepZGdymj//p
dsx1eS1HJNRt5zUWKKGlSIEwy9ZPpmLPDAJOVFoHxcM8dyZbQUdRI80J4BYvyGst
vK9xRj920x3HQoQV794E+pZXTDRjumN0l2vNGHGTM4pjS2xTDBk7DvMJHDksDZyO
F5Jp3SMypW6OavkocQdrYiu2ttNP6VARtC9QoeI4cFk77WrsBJUdyETAQXwyJSwo
5ZicF8QOWKpwPCLbzFOgKai4mD8ckRIr8nYuPyOMKaM2iLnSsVGUcuPX0u+gKW8w
vvjxakNnNEamj0HWp9lqZO2+QnYqejh8k4LIoiWvzpkCIwVIBoCT/EjjLmvBYd/+
9REMqFIbo2LM2gc08OLaYv6qInTKgvBPuKVJ2S35uN18Zh4vhCIYD+j0SKWKDhAk
ehlpwmLmy/HZrA0tpFOay3jvIxa1ez5QEHz10Cyqn8Aiyr5BUjPtzFamt3A7n4jH
A//HXOAgdTrMv91g5B/uCzDFO3gE4TAAvncNcBKxSJxKmRSkSVBfH+2A50bDfKc9
pfZ/d2a+0SFl0cped+19BC/4lzUTi2wEXl7Y8QNHCREJpFx0f2JW41xaDvNGnrxF
Q09ubZKwYBsLR8AEh3/efp7MjKRQA5QeLkB/zBJGfpNxtmhzWjNW/k9YsG4uP4V/
ydTHg8k5P7Ev9UC79Afg4HYtbxQy+TS0H3+eqF1zW2L/tFk6KxDMCJE9ANtmAjav
3UvfMHfy3w9YeTvSYUiDGOngMkHSnCk0jjdVpSsynhp+XYNqFjL1MonKb7Z+j8Z8
PeZONK8ZiQnQ3D2ycxWJnKOmWqbvesKZuQrOsNMjI4U6Oo2ZkAgkPOe2JebtsB3M
bbNcYqpnEeVGWuRwFuOJInufsWMhndv8Fi6YJgLvzI0bFu7C9aB+b1ClBjPWVK4P
9dAmzKCv5vAWg1VQGktYjGIAlaq/Em48LKZklkhQjVWBjAoj6V9pvfsgeraVY+wq
cuP5TamkfyCc4WjYnzssY3yP5MI+UgrEgp7qiPTwU+mzKgW+jD+O4+ee6jWbEAE8
OSAYqZpQlVYuEmSweMriZbkZH5+8tKjbZksAXa4Tkx/ftGcDqEUu3An0l9nxG2+s
Iz2vBZ2nOVRaDASY/je091gkAYUKlWU9s2BCuMGRmWB6Y71BmmuMWgC697Jy8uY2
X2g8ZMfGiFWkSDcWwU/DMgoV2b8lxu2D8OGc0r8d5B2Fxi9l+R90qnI46C5g5hhi
nhD8Y0kZguoeKoaWgwS/7juhaHUDerd2G1VudgCPUHjAYPUpVhPoIkxptdLCF6GJ
SSfAFVu/SfWQX3EXHIPWf7aqR2lVasb0J+NCHLHqSCztuXa7tXeH7VJo2+1FgHAk
z7AnU6ikbM6/BMmw4P17GqGVQ5d7aZhUy/6QuTX76BgO8ymllGE1mKBfm33GtoOf
ImIKLz2ZQDarSgTe7UQ8dk9Tbpxl/ApJES9Tx50RDX+oVClYv9GB+Qm0iC0hGEY+
GUA734poaAyf6WyPmCkzpe2/pnZMz9zjuvRx+70eJkgdQm/fuQFO0ddQ2sVypHXb
N6SJrXM9zXKXekpwYUBHUzVMy+YbyzP/cDr2RTSz7qaQpJbAvCc3LcMi9tIsmim4
Smap9CuEMsq9kfe5V8JObujgIYSUgySM4tbHT6f6lMZQQqIyNNdiZimzYVkXxurk
Nh4BhxF+wpnp6gX1v+t1NvvOhaKO9wnx6jcpJA8C/UN/dCJysaL8zP7GFtnwEtft
Q02hYHGk4X0R3Z5+FOd8ZTFF6lurMrq6ABIocjkcUNwgf5BIxqyW6x0nSOgZvZap
l6NnW2bG0cqbEzhVYtdS9BuE4hKCrIUnkpsly4Z+QSKWRjMo3njyPCrCHvzDjWFy
MI4Ac9YQ78cEr5ia0c+pArsLg4ioje9s8MreEcCznowoXacG1m39qeYrb+E9+mpv
rPXZUn1aLOx0wnpzs7gRQY+GpScEA7CYwORNt8gYNAr+9QwyqWVPfrtIvYzvyV9W
zIP5zghxPTedJsKnRTBEeQNtnvEcLGVQxBci7b9T5qz+njhWb3++CJvFv5m1Qg8k
LHdJmfaZqwsSlPhWFxtJtQqIjWEtg8UhHfuB58n6YIU19j81h1SnUD6VeSr85303
uPZ34uIMq92gdTU3CenA1ThKCUKolOgQpNNVz6TH+GlQt9hzyeC8ei7OkVfJdHDR
W5Fs3vp9ulchE0V/nERHQvvLC2oxnj8d7fLNdO8hOop4t1U5DBuoqbvdY0x8W/On
ebCyJhokUmVxadFR3NnweQRC44b9zD0Y2Yy+oeRZB6g2nHCbWiELOzcFsYXF7xhw
SiWfMGouDlfWfYAisqBiaSPItgQO2aS6+Ids3+IGtwTHPl8FdNZj46L66kgoHXMy
8QObVWRZkWE3ku7XNIF9pZTA5G5NTM8ZskTObmJNrkE4FdJx8zjL1Y1u5lJ1tG4i
lUclB7ulJ9EOtSQviFtyyAqrOJ/FmyOezQAm4Y3pqwVl9fxstccH3bodTl1Zb61L
5bmrH+USniiwgbqWbL2gXsoDD8MhEdejlrNHCVb8jMkUVFU0gpR97/r1oHh6x4s6
TLv3FgX/sltr1bZN2ArVTeS/jj1ClL4LyPj3RhhlJfSdT8LUp6BT59w5uvIYOMaw
8D6UTW7bOynA2XObi7gFdPLbSugcir/PAonlrqeb25Kzz8APDew+ZrE7BGQFbxJV
/ZEif9Es+TuqGknKC8bSaUI79hrfF3Z54MlB5TFZjsTeABIvT7DmhKQbwSnJOI3x
XqMx+Xa0bambk+yT0ZG/Dd6AIz1ENjxqG1YO8RS5IPiNpZbU3D1P+11P3p7iEBBk
KkQ7HsFJYKwIpR0eCEHASmJXVmMR7LQidOx1wIlNWkEC0vW+RoNfxN8g2EFBLJGW
EIX/ZUJ1kQyj4VHC5s2Jo+49h4qdJfa2Rb6JHdVxaD6ErQKYRO8P5J2LfkWjovTg
BAdAXsO4y6+1kOfYMkjlOnIau46ERPH2iFaTBOqVSpx79oxG+uHL3uclwOG6htgg
gj46oQfO439JrkcTOYgaSa61xC2COtuPX1ZZpJKzxhW1hs9vOvQ85JFeg43Qqqt+
URS1LZTXP4mIdIb6aofUppCx3Dte7IoYuEYilj2CE9YoH4XAO7mupSFeQrOs072a
IrKebt1HM/Rl778ijPtbhyXLspq+4ACs94XWdRs/nMLp5l5RVPBK4v/O4tSRwLXe
UX0uQgJ0rKGgLSilHf7wuMEG+9yPTSVQavEpblMOEMxq9wWcl7jJ6tmgrzk55aj8
+80nSn522rlHHolv9FvOgJVTHFnjBSLQStgIcDbaPjRBsPluhGMHeiUj7kDyd/qK
6V7NU/Dk590U/2A7Ko3it73E0Obw/yZYuugLbMx8HumCGul5XHKh3S4KvMpoRb/w
3WSC8V4+HZ1chyAWuMFEiR3GdE0nPmaw+uMf2HIfgmDIzqKyJLqnZEa/JGD458Sb
ziXGVTXSGWLqIf8ICPYF3ThuATTbW6euQhWP4B3tRec1W+dJsQVc/W5Ks262k7n3
MQEZSW2UyzDgHz64r1A0nJ88kYI2uNEVwVB50zBD0rzoEaU0pgOmrJGG2vqW8orS
PX2dBiJBj/5oHoEAm25SyjsTOHQDCkvmCANXyHmwSsIXZzdbBPUF0HhgoGFRGkSX
j7l3p5cuVm9jXWeW8AN62z0yJn0/49Idu5EA5Od+d5Z+SI45X+kNYuAgAGVgqHzb
HSJkmFnLFbF30F4VqUy4+6zJ3nzqRbyvQDtSxC2yPbaX5Qv0pKKrj0yg3Va257Nw
AxruEOSr1Vr7yLPChvxrb+Z2LNEF++HzktR29Zqag/NNG9fSWrlgdww7Gn1Os3A9
vo8W0Gt4lIc/MpeB/5+APUbvQHLvkTXFtiEub9ugS/V7CIe6HlXd1PdYXuXDiMx1
EDKB+jKSEUsPYlVGH2BTetmSjxaRTsxxTRRUV9e/PRoo+zK2EH/wUffURzO1yivq
L9lfWZ9+cgr9kkpMk49/pueDwl7OXDYzcTHvLEkMn7Up9HPqCbBtgIDxJRm3NjaC
0XPbyIwje96T3ppNBsjH8+EnB3gGGkYmNydJyJv7soTZOJZIjctqMzSiLdeSm0dE
C1GVcMJ0ZEStskkVpmAD31lf/jGFiP029MVqxVNQe/aSzrEs7vwhLSTFam++9s80
T4n9HZcxHzKxsuzpB/dAWgVMr5H68RoPRJaCE4ZT3ObXITw+9c/fIPh2AvXpl+Qi
tEmgG3pwtdVMn000IEIkAMcjryG7Iku3+zDT5WynWtitVSwCLPsYERIDezBShSVH
+seJ29sbjtTJd3DbO6fwisjieneUCkIUp8Wnz52KNOWpbx3xF0BL30vgqDM7Jxrv
HAAmleyRNmIMUTslccnkd+sVskcPtoWecUVQnssr/lnLW+38wAedMBxBwlc6dX62
YWw08+dmAjssrRs3+BEKgUjbWcAwyCRAgPE6vUxodt9jHv1IVxPPfkcKeJCGy1RK
SvF6FcrY7dJmaXJNHr67I/j03Fz3edsgF39fGNVC2KJUp/WHptH+YGncr9sg9GIN
DL72XEzenDOhD7Irh26F5Ev3UMa03L482CK9D0K6gYtZpUR4inJRrqy0lRaUvesV
AXJSNXHlo5w5QdYGq4PDOP/8TddAfCWgXPuyU6PY9wAC/ur1MO3JQDLhFvy9aULx
2FMoA8YTGatcpf54CKv+mR2pdzF7R9pukewyJrXQz1Z/qJ15nUCsTwvBAhV04ojO
0/5YIW5mB+Zs/q35syUxrtVyU3pA6Cl9YbhcS13/0nZ7O6KH6bwPMaH+vW47ckG+
LnLri6TPyhHpSn34O/glzWB+fUfeDfPLpoF92ttu4cIDwUPJ3RFAPwoBNbkobYnd
2HxOrEbes8OACQsMVcOj0P/3m49eHsIBIof5w7QrlKQ5RaK/lhMcsLymN8sSHZwj
6G1oihBhebJZKQmJ/IOIiSdS1Gy5PZGDOpi/0uyX/2+I8y1ZtQPEn9gisR1J/EQ+
d4NADrFeFcbBeDfUL4GX2vl0s/gmBAeBCh5geRsjv9lGc+OLkHkwi0+2Jd/Zg859
ImGREkg3703vzph7KKpFU2jrs4VbSTjs8CwOIbJqIFM77MW8hJoTc2xCsciAx69e
wJuQ4t+OLO+qhhk+L3WnJ6w4amJ9LoKEQM6VL2YSm3KPNYKrtUaxMti6fObXbonw
JQqIX8ltX+px19z04v4YbWrudp0zDyH3lCbBPDw7YeCPTnEGrkj7dhvCIjcLoEUX
SgHZtCKcNvZfujZtQOBCNVz+SlbYay8s4+umbYMdWGP/u6/dioE033fLVU8tDdwD
ISn1/qvIPUFjpoGO4WCPHPlo+TkcrKFCOmYkLRff3yEP0YbrP8MirKouZca+JS6I
mw7dO0Pe79AIrgsbdYlRlD4YCPkuKzKR/nV8wCrcjWXUmvXeu+8H2wLhlzqs3L+b
xKqWmvNgWsAXf5+kPU5TI4Ii4hV/qadX4YDaLB2mBajjsjaQrY+7NxfDrwt1X89m
4U5Uj8hnpT/w3g7SS39OTAN5rOrPReYi6jIm8hcdd8UMcQgy06vgJqjsFyp0snQi
dquCWKOiLtw3uPaTzXtpJPrk98UNLfmNTfAWJHclMRnYG/YwNx8eQSxJjXSmxh9h
ynFgVJ3BV2HZYv8x+t/vQg0yqsqE6ErvC74Lsopf0+ej1nhkhuTANITDXhLNJ0t2
JDPbpCDyZTVu1wQoDel+ek5WBo3bdMTkdQzWgXV6UGCcsooRYRmWwb1dQy1daYyT
t2Ka0Gaz8GXnj+V2igxDJDGZWZly67m/93zV7fPiQB+NG5QcPjKyPOnRG7ZEqdzp
3fi/OVNDvZDGkSu2NkQ/J5euAOfbv/HCbnk37H6jYt7eAniJMkgfPXjoUorEYGYU
WAK9wKWHCe+9RF6ivB3VExcP+jEALqHiFbnwCLhx6Xo0CkVgx9YMV2O2GWbm4K41
JRN9iVHNr9A2uuPd8ytPaVYdzOYhSoGnQzHlo2vNfca3u6iRM4AkgmzfEJEECbUD
cJgXbraViyxuRIBT2D6P0y3y0Ls6zeqXD3nYDb1EVGZyCvzsm9mvD2L16egywtsC
LUAPAeH1N268/JdKi+lTD/d4Q+3X8nlX81uG2IjlxQfPfJRlM/YZipWhSvS7RchB
ciK1zwnROrzK1uImEvDkVQo0hR/Ch9sI3lKo41Setsl70lT0Ca5FqRKBd9E+LfCZ
RwN/jLU/zcwYjf1AYecljv7sn9up7Bwx9/4CRaOWVACvJgGUzRCSwH3Cpxc9a6PC
Qw9NAchQyBshbSyqHCBmtN4vh6kxgYJddNV9w8CnIGbxd2E4lGIy3437l4J/F68F
/bsyJ482BmpwVrdLZQG4ozKTGgvqokFrn/ABv8V5BxceZGFmcnb6nbLSRs0jWvCJ
W66Z1i8PNsM9PDvNLgqoqlMdG9rG7QnHxLZxHdvugIpxiK64FBLxpsDQY40h7Vqd
q1L/TDC6NMaw8q5cmcmz80Q1fXyWpqx6iC1opV+wme9VKhDIeC1ElqfvkrEgd6JJ
1h+1luNqKE+efd+p2oFanzqEXti+nqEJPvnO24itvAyHisgr6UIYahJB/gK93YD9
Z5qy4YX/gHGHvKSKMrjOO9+HIsSmC/KD5MxC/sbKUE3pZBGgDCwZgqUZRKTOS/qA
4FxSCKQiilr6IELVHJ51EFpNkN3G2EkcOzmVa9kSFVRUF0nIExSPfNl0P2OmVng1
sNMxgxPVbg/CSSlVuk5kWtxY7AijvOSGXpr9joFEXhhU6M1OfvkjF3okLuB1yuge
LCidNzVqhhdj0ALmtamExxPd2xM4f2H6IO6TLzzfVg8j5ToZN4fVo3/QKhetukEy
4bvktEc8TKZM4F6hM80uk8calDfHTs60NTbDcSHmrU1jkW7FOsVS9nILjBaY6Gta
PAt1mLeiejmM8jRtuvp2LuPHtq7bfcfUwNO7BpCCuQ1DOtm4VP/V+XsN8t9JD5xh
xjHTl3hSr/e6t2rGKEUvpp73dd2ASR+172ptVGHol5KbEQk/ium/IIvnrFECR3SS
Fk0Lk9cGlejvDmSRhWR0drlZIn0ZRyrQKuUSiX1DReRexRaXXZ2DZUtjPvObWGGL
F5kWZMly8t8SFQxmEkmEmtfn8sSYl7Vq8i+RbIeu4LD+tFo2ASX/l7I6kkzhjODf
3FqCA1xVpO0qV4bLNXd7AhKBt+BuJseRCpdDo+KHhKjSaqGRDE5EtQAll33af0HI
AKcjcb9+Q1Q324joR+UPxXYVmPXEqBjJjrtbo87sPotveC4Y9qYw4DHyP2lCTJhr
jVGB1r/lCnZxuynz/8QFkGkm7prdCnJWq4m/KM5lYvqgXlJvKSQ8P0b54rQSwVoe
iewhXkrLozz+NktyKw2sCp8Cd1N1AK/iVz8mDahZ/GrP29I051A2wW6gZLJxBURP
45+iPmUy9LwK6h1GqoD8xvnDtBLvV+BjLViLo/EIMwVjWK/2hqwe6HFLinGjs/0S
lZtirvZHHDTvluyGUYmtSC4h8Tf72E4cwdeidlXc45W/f2amRHgGBWJ291UVvWXU
sXosse68hBQKZBdFkGhLOs3rRss2fYFXD9EhQTdbZkTwtSOwc7MKO3WEQ8aCG47Q
jQauZ580mFQAR8HiI9bABs3DeZMM1PzDefu+yA53KOP/heonny8xwQ/1nrPp1PuQ
4VtfiLueIRUZpMfQHeyd4GdmX6u6D2wL5CcvRfF8U/MTycpvHhR4xbR2Fd7DZpuE
rbQTXvzcUiwy7/WZp0EtAbpZcrhUnZtvt5D5RlYw1C1JPCjM3+ha7HNDN1te71rC
o5EEm9r1EGBdVe+BEp5n+vCC5RV4IjeJixDPTkE2Yz8nEdu7J4/3Nd+kzVrePGcK
oPByRWt6Lcw41caCs1gew2tN6lgt6JnH4PFPkalNby24Xuni0SRrmSBSIjFSX2l5
fmqTV/TWNfvRZt/+ajV7imnb0lL+eRdvV6rfTGpfYmg11TtcGKs+fTlkyB4U5vLY
ArRZ4c3CIVOxiLCWOlPzb/uUSaDXROFyJs1fXrEqyozp+cbGYYXejZ84FsWffv3y
OnrG7G6nO+gYivxwR4qBHpK2hiW6Vbj22j5cUuyBJWzQbr7Vu2axb1Ekm4DrgM8O
mqAZ7DWGcOHLKY+2ZP5plmAPlJ20JC+V3jVpdWG7L39rqQvHCIr5PO80tE8p+wGf
ZkE8tZuPOzqc/Z53w8Pb66XCGpjrUvBY3TixVPpRFf14tSdo4q2/HoA1V5O2Zq0P
nFv5Ha6zj2V7RzoCOUZ7O1q1mYjuXkWX6OR0MAivYrKugH8Z+DceEdYxd9xXiSvq
odcRoitYM4iLCHa2MeSkRTzmUyc+r13qJmVU/xp0EQxctW0rLejoFr3YYSZhW+n1
jsPRd4pydm72A+YsrOVvEnYE2pBnjWIW56cFQFjxWKqUSK1kg9+bBWPWRl36R+zN
AgPM/xER6njbC1dfr9IjVxz7eoZ0y+ZmfSKv2mDr8BQn8A0SU4LldE7PchEgrZo0
J2gu9OwTOxsToh7vDzXg+1UopuyspX7nEgsMaw4U//ayiWPspQjqzVoUQIuDM3We
2zCGvUH78esIVivRbTnttoXxvdVuifLh+7oTVowNZZi7GCFGPUfvPWAOBbC2iLeT
b+6hf2TH5BmRD6Xn6HrVmuVAbuN1XtaTF0s6jm3OpWM7MfYXC/HP7VfqSJAF7Wz6
MWwy0DhS38eRtiYhM8m1vnI83MQA4iY7DyYeCrEkDr7QEDcDZ/KFwWPPveoU90dj
gjVZExiRqlHrFDsI39Z5HRIMrOe/ad2zVAel9maArz3EuA6Wuc9f0tQCp9/7YldM
/7T32cTZdQ/e4QBsY1KbsbgUzmVvIVYwMCtIoLNIbR/1dsJsTKVerIey7oK3KPEO
rgmqsrfpxXZnx6UOyFXGCTxaJjadjm423mesZgBXjsJL7ilOerAAepEgtisXhRIz
5rYnFiUxP5oe4xiiaiuG2MSwKaFQaZ0D6/1Um0tVD57oEQ8ae1XAsw7A5+d1LvhY
Squ4qrQIK9r0iw+Qvn7ufLTqUyKsWGREpBfAE0QgckNVJ7j/ZDef+6Eenc+5Habu
aJXUtsz8rFX7UQgg94wo4ia20a+OaMRtRYjr7bdIqFFNZd5jyjAVkk0aG6cO+KtU
nyYpquske/2AxAYrWEomXOhp39eutvjbHQ8UrDJP/pAB4Xz5gjpOyWAvKwVNKk+d
F1ywuiCuFD5fD47zPxSelSGzcSoPMl8cgtEM7GsengQYPqJcNFHqyuPB7CVZGa4q
Fx/d4RU6Q/zmmHgSbCxfVpGpVAfUJWwKCiXIazYLRUeVzDVVectGlFYdEyyYm/5h
khCpZxL4wug0jBZLBHUN8DrTH4AP94Up46xcZv5rqNCg3gEuIlfPSwa4clYJ7P3w
+SW9X3pinXgqLHpM6h2h/Go9T99kZafIGRiCLyaDQjakGHHLLFDj68jsh2ZorS7K
0cHBpHmkSHJ5Z5eb1mJ9a9iRv3McQ6vr6V4sWZK9V2JffDDC8qhBbtFvVgGbLvk/
dv8lP3oL5BOJcw/k5sfH6CvfAPdFxdL2CInid/PF0b+1I9mFy02/1pus6ICzbvwY
1GpXTdcsXa+uQmwp00VaI9AQ3spor3JbkabmFs0pMTwJqfifzbMh4/P1veDAvfed
QbZoMxl7aK72igUhkjuRO03PMSLk//0hRf+WN4VHFfTvHf/3cBOm64DnNLL77bHq
Ye81L7ekvqL8bLBGAbU3D+3asNrlQk2Ljeu0hmyDz18BXSao5T58oZktj3NisA73
rqwBAaR7biPhx050fKJ9hd4Qj/xYtzDcl0GMX/5gge7qh9uWPq7oXcoFtEdAX6mS
yccDw3nr8chZUv8P9top6SIigkgN+LE4On+yyKrFUdYULYaID8qEeWT9UCCpZshL
wMLiJNVOAkaoOIBCcdn42wz5XLp1l6C6uLW8ZzICg2dJY8yJN3Go/mRkA9lx7z7A
kpHzpZ4dthyZtIDXtQYz9QFMpHxhzNmPW2mRi2QirVTtYaCKFIFqP8+2y58hk9es
+AL9CDgACDivmGudDGPCiZxB+gdxRRkdabmzXAII9RLBFQjTw8I0xmcRJf6+JJho
OJub0Uhb8Dx7+ZwgxlvUcmdRb2vFCp+aTvSchyAZ9F24J5yt2JQ9hIvxeO5V5weq
qI0YdOLiJAILuGIj+iZMwSrCTN3Lbx+Cj6Kx0EaBptdh4CNNKgURMzBTEFvS770I
mHMEc+3IUt2ByZxExJP3kX0x31tOci3ajBwxwvc4p9fVVJYmy2GldvfWWoSnkRBT
5df2KdHPgE9xp3vRhh5Axnx/Sekw/qBfc8CTwJOmTH61QyULBotLtk4KB8k3ooge
u3P3tIweKZruQZEYuReuvNc99EGIe2hCwbecb9KdIyRi/F8tHhbteozD1ch9V8sm
eHGrU/gxymzhyN3KzxfZGZcZPA/Nd7UB005apP1cP9I/SvJO5/4mSJLpS9dPmBIO
37NwbQfpamfzWulJo66eOSBMYcfyt37yMfrTd5CNg3PZQU8EBk3IQTW2bYnNhlzB
hSix9uzvKFpQQJi5FMX9ehtE43kzueKiviRL6O/a4vOj57dryDyHCSb5/n3q3g/K
cwiiIG1Dyld0dVmmhANH/ONm7kVGZ0asT89okw8O21k60zEpH8cNasNOqRnu34Bo
BzXcIcwIOwBjHrQCDtvliQdfDvITazA3nlkVJUrwKQJ8vlyume9C9oudC5vUePOJ
HQIYJgtTYw7ClNfMCSonZ16qNK7ZkU5T3lbT5lASQiE0o2hwwOc3bcsUEGJ6V4Qz
/S0tv1Lai/wUyR5hnkURX/s8fPA3Q8bR9Wu8qNn/iNPK9E1wH9ikOysyHBQbKb6D
De1ujphBmwcqlBnCeRJ99p/ninefs9Omnoq0R40BtuD6pdlX69uJIcMDdlXNS/IU
B0Pijh42EhJpU41ytx/7o2NRtPcp87idZ2hdcbvO9DzqzOgvOgj6o2lArgqT33uC
GSw6iF84G1jmRt3XyRfOnQDTmfzOMYca3JrtI64/mmPA1owQEH4NE0QYpiMASesj
CC204Eb62RxQA2o0nbvwrEz3Z3GuXv9/LWRsmTepsr1KxQ6COhNJUqjAA/OTzL68
fNxgQkBsAsfUt+yWiUSwbt2znNwdqgvAVrVPUSdxrAAS6i947tqTDsGW0z8ifZF3
bsbtsfrnWAi/NlAgx9CVx8g2LHYTpfTy+M7J1LgXI1BIdMNDfiNpVbP0l3uL3vem
frh/IBCeqE4BB/7NhEj/ETSIRpkfekJSh67koM2Gdl/pwsLVR49Bzf3C4YME2+0t
hJD1KJp2exAUCcewgjUT4ZVunCw90taB8bM5u1e614PE5aXw7Xng0BF6UE84Jjn7
qbDcNxcPDvg9OBa5t6TWA2zxipdBJaJF6Y+FwpY+JqJEegH1dz/SA/WnVvoIOJ+J
sTgIBGpfqonJRDocmgGNVuHRkpfEEUKlHFsXRcJZxBcX4EXyVREvwYqa4d1ZV/gf
H618FiLWKt9ScMDsK9ISQMNAS01H3YsanWNRqM7q2LQZH+IBLB/IfISiJYadlIHh
n0N+9Nko7Vpu8LIPTCLWlyWsZlY8ZFZpiB1bo3Zi3IkinJMC/V83p+zN4VRFYRT2
71T8rG7NSmGUx+9QJQxRXhDutRtkC/5mS8h1j4k6lYV2UzzbFYDTxZLkFT3nMTIa
N4HTj/RQ/8cey66VS5krMNKiwkC75q+Whkg/ND9OElY+rjrsBqCKIXdiJOUqPAIH
0s04tq1QuGXfsQkxXxi0CxOIV+ObVtrji9VtXjiAz4zJLFDMImhmscz57YTc6QtL
yqRphFYIQtGaFCEH7w8/8UsboL54ebRciqO8fVA9rNbybZlw5kdMpRBdeCCglcAL
u4x/7LEEqHD2rGic7cfj2JZRGg/Z/Bgi9EiIPzAbOZBHAFpQoCE1+XSp0sKlzQEV
j1Esvxtle0Bv5Ctw+gcr7olkpWmNaBXcK+VaRqzdpjFvFSxpAyCkFHcfU9dbGyCF
pK9a34S2KNPDoOCIuRC/vC6DiuEyyUriQXUhAwrWTRybHlQODX1x4QjqADHOLVof
QV3UB0gD2iXFUuTCvt0ZvcuRMt0S7caS04cKZ4RbVpTel0LtaWIoY1W7DcMdNyS5
LRvOTy1IeA4H4ezktTvl9AFfYcSk54keXk+Miy0woHUWW9xYB0D6QC1rtRR4i/Tw
iS8tg+E+4iD7QUi8dEIkcvmC38f9hNfFHXvk8vDCOac3UX+pnsl3d1vGxAY6wPVG
OYCgCFd95y7NZC8/9OeMNgTso//Z6PW5udRCWQB1H31TyP/FMMdoz1N4/tKXiotJ
jAiGGOB/iq9yuQLcA18uBraFOd58VOm/NdjWLUpTC3nhLHiBh3muVZzs/TK7CwVs
h/wAb1qET+bEcsqWoUQFa56RjPr82WmB0IC2mI7QtrKkQfwQpG6TOwq0KstpDU1u
4HmE2Ul5IlqM/nyIHmD2Jf7b7qBRReIAn34yg3DFfYGZ3qil7rFqADBIqsIWEQZZ
YONS3vdF5d9rmCV5nqLcvY93MvOO1vSEAHaG39XWFOQowCoqe13g1l0lmBRTRLG1
r/bBPUA34kfkriHRcB9IVmkhM+AH2VyvCXWGkH/6jA+47wkJRuWrOuw2PPE+tOyJ
icBsG1MPjxIBflxffk02znEmTQnxd+8GbH7xVJ8X/nGO/RWybHWfTuvhroyPpW+v
w4z3rEV8ChAESqaymOjXlQy+T5ZQt7HJqkPrNqfJQTe11rc8Gy/anbmKt43riBW3
ys78tu6vw820cLj1t3D6/pToXfwV71cukJ9LIGtcEdbBqyJwoYGunb9G3hdH6tUL
BRSQlFdWi6SLvOTNgAQp1IIZCHTJc/lli13UtbgNGGNF1jS2nc2tBSMjDWqdCsuD
dU5X+Ti3Ft8IzouAkv5pm/EG7L2hEapajc4XiQTIrWOcsN82lyt5IotADGIIgugd
jHfsGYklgHgs5RkEX1IPw/jOnHv5Q38XS32Tgb8G/rnI7LVyKT68Kz7syWi0rcsP
yZq4g5rgYXf8Wc3iesF5LiN+s+AtbNhWf4FGCowjLyC9pdxBT0/AOeUHoZt2ALuh
kR2y4tpczx5tYgaK9oWXkllKwox1aKEKn4W6ZrhdAXyv9/no+v2HgbIhlPOARkZH
A28Sn1ChlJHelEQhOZxYYORY1+cKKuwkM6Jq8y4XY5FK0bvp2lcDA1QNc9aj1JRw
5h3paa3iSop2NAsePJZ8WrgloG9ihfMPSGmEvyN8mKCLq39pSlNa6k4yVCfrL/ff
lcQdJLFgcJ17XMMd68AUX99AfE8WA+jffkTqw0lMvHNdDUOpWWDWwDUHk49x7Exn
AtEABjURnq8R3WTMF+/jjlUalVAQ5r5NxTpojp7mTVemdddLE25sOx/DDB++v5gs
DsBrBVa6PqaZdAtMGbMb3uZy4N3HbB2IbTHCvX5LwCBbvWLRigpTLCBZH4NparvU
hnvmtNfK9mxKJmJ7K9A669+Sv7T37Cdbu6+zzrTpAhVupnpI+us3jcGf17Bjgalu
OURvn7Y5ePHXsW6vfAMqm4PbroYQVxyvy9v1uTSVTvLG8Nmgkk+R2FKDJbLmp0fz
wstnTtFvewsINu9gAOBu/xSJ3HLYZoPkfTCMr4jGN6ZlpvVChyl/T8qEvxz1psDN
xP4Ax4+JOtPjQSoIFlNw7ullubXvmRh3hELtOQE5VIH4QxzKS2MnczP8raM1Z0HT
xCns2VY9sBXskf9KECu3yDI+qd9MHRyfYJVPVFuX+PNFxEo8gIDf5HcgcaHwd+K/
kZzLG9i8QHXIOK7IDl4EQNNWmK7uBiPSM33hgRvk1OGvNy3AlfpvLHMgqoFcXZSt
7Fxt/kes4vF7hemnV0Go68Row1ArMyF9d9ZZ1b7PRA5Kk4qpGk0biFB0C3wuVkvx
dj4EFB66M4dg1dtNGInm02AtKFQri9/w/kk8M/OVJNq1knkVsAMa1O/xZTS6UPe/
WDQZXPYwCLsvyDhEUL3Ptbtx3z6qDmrfNbW2gqC0fbqlr6DHqe8q2073XthotMqW
Wq+EcSW2vJenS+GGIkHJ1Rnvle11IXYUM/CIub5CSVEqu6QqJLXymn7CSEgzQVD4
zjjjxolyjckSJSZFfsrObY2EaslttexPcoonnAQL7R3UPLcey4DZSmJ7yLPF2+uG
7PlNJNhCMugi7dyRsXedMNa9ddDoU+rLdRd7UrxRlYaZImWqce9QqXpQyUjUz/1F
TZAilGqhS/TKCebx/YKCAjF9PZ8KpEkzFYUdL0hQPuerxP9XIgcadrKwo1/m5e/I
9nvBOmC7ZvpL+OM6XjMclGQ5/+eh+fMs9+vYcc1yf1eghcK8tgZYs8bqd4R5jO/H
lC/5Z1eJ+jXdX6RG1xh2EEd5QQoAOgfvR0Sj8K3mNX9UQfhDqxYxNRUIQ7vkoBn1
BQ4u7+zDhxKF+8+yYX4ENwwjGQzulA0Btx/p8sqTDS4lchhwi7PiFJXOobzJViWc
Y6K2332P7LHLA3DQf7quS9eHk7fFSg53s4qX2/P9gInrBTEJnKMQp11QMrvpi3xS
V+MycY4DHQAY7wRIlHy6ivvKf/mphqfGXWNUGqkia+F+I14l6iW/Wcp1H/efC6Jo
VKO8dANbO6eKY8adEOMSrfXExqvGnDVvkkAE0RMDaBxIK4cP+hB3b1ARhVO/wXU6
N6WgNYJMh7gqjyAp5ju5o1PYMEMXoUAxjouFvWrzbNmTPDV4ifqf9axgwIXBdwP7
UUSKcdtxTZpCNxC/+oZxABDQySvC1kGRFzp0qNFcYEcu6mWFprs15t3VuVg9fqsY
m5d8lwxrKn8bfp+rDTmQTSrhR0mj6lJtxhbiQ+K6/QhFpN2G20V5wsTo8rBtQZZW
hUHWu22kzGBaNQrcRwz0+iKI8KlP3xLJUl08Zur+3F6mbFeOvlbBMRGPJRemz+fM
mT+NdPqTNNsSNLpJcsgqZ0cnp1k+n1oZiXyeJ8cQYUo8LBs3IOZN71fIB1J+PhwT
OpeQac/j7WGg46RhxOc8HqPUddc+QBL0UR5coFQ1xKOCPnS0iqwdSJMJGAozl3d+
5sAnDNozrEUn63IKH9TToy18k29Cq307nyMi6Uq2H4yQEk0m4VeFveVVgGJMa/sk
26snMybHRfD72uEWJkyWZDdkNoa+YLQCaDW1JvnAoYTzE+C92hl6kjAHQ6YxDzms
c/zooo+mHZACqoVUcAcIKuULCM7BzWbs+iZ1Gq8ycpi9cw31JMkvELckSwbH0rrm
MsPaLvmntnrZwls/GcIYBQasbkYJK2+2QiBcCeWO8AHwsojyUSiFN9USPGw7zrIE
RREQLIGMI9EMhRtY0aQTNs384bfPnISp0mTa431WWjH1BkHwFb2pRF9NqKJgvLCt
9VLnSdyPeBYxpB1eWJsMvMF7bDhHAUsU/lq5d+ikHV+9XfIAsmnyz4MK86/qLn6d
5ua9SG2kFufrpgPyjH/I8WZxtlMmfzwLrDOY/CYKyUf9rgaLSOz6KMuwwjnoncxB
sKS89LX9sIZiF+TwW7lb9vJ+vp537z8FseUGszIokicKNkAqS1+DLroWSN/g9aF2
1TksbewApkflhEq5X92rjXJYPWu/Db2KRsmmohwCT/D6K9N3R2r6zcb7U8XeOl0p
oY2uYzXhR/WMdZww3PEFdHO2TzCKCjhOYpS6DY9gCpzSIdofQRoAYNZ0kgN4xR05
Au60yakvuZLem4yFE6YRDhEtqq7ZZY5PpZIUa7KkYAkBCkRfB1IhrBKbKxzvrGjy
o0wZp9mzmPs9vsgs1BYIYJJE1JJN6HOA7fh41ITf+TAYlixdt5IQ+UvTcNklZn3G
xDF97hOZ8QVHqCjqzZ0AI97hxyFNl2IvRpck/j78jZHNiaWUVhs4nnI2uVtZ7pIK
7oNXf/0i84RbPNrmWSpr0OA/G29oJBsoNI29xdIgxzeYkk0evFq7cmX0OU9G9bV1
U0qDT7w6BA/cNGcmTm6krWYKxdyqkoFE/GkPlq+gjZChj5eG4ozunij0C1BCv4E6
cOsAojmfzy0ArPbPS3Ut/eJmLDQ6z2n3x9T5O5UhOWBoZ2sh5A4PgZNzjTB505Bg
J1PjNvEexUucHnLMQBLozIqOmAl+gq6303kdiCRDwzauVs/J1w0kXgA9PRszgwj9
7tdahie9TDyaDKAgfaMWK+SnS0CdeiOyEH8zrS62Ci0h7HVuoRfyMybO+DaRVwzk
/5EFp1MUMUc72tV8b2DPQQlgq/vmFcGI0B60RbUjYKSMLh308IKNjbnijndP3DZc
Umh5okATSj/EdZz7iEdF+1OKdI7tNcjq34ePdifU7ihl2Rhgcvt7J1kCZh05TuK7
vLD/ucxvyvYGD7QbW2REQp1USDn5zb6it+1zKceA++C/Se8UH40qSv4GMCVLHw+e
yH1zJDx2LT+3S6h/kpy4aQCDli4x7pWstGC/DTtKXQ0bUGmkse9gwTjPxSNIBk5e
+XRQmd9Jq5jBvRtElmSuH+GMg6rdIV8c61m40967fNZfMWD8aVyRmkKUb7vurK6V
b0SAZUYn0gOUbCq++ZtXtt2T7Z1+E7IVFj70LtRyVSqTG+38hpXQVGZqtNqPwwrW
mza3MrYJwRuU2vHL6xo78VtIYWvuqkFVL5dIrGJ9f3PpNnhYk/n9dZLSgTu8d9GT
I5QI9bXyr5oHVGxl1Oo/hHp+GYFM5zTAhUf0rpsI6ggnMdR/yUipFSZJDi2tUYoe
Xgj5pgOrqswPOMZkQC0vyd1qONV1oPGryuW8Afozqwr4Z2DTg2iGAyETlS9rD6ei
/w6sRf3Op4Bw5Cw0z8GU2aCEpVp2hcuSJMtGUgVSwFbv4qdvePM6cZ6fXqvPCA0C
R9oEG/g2IQMwimag8oKS8nsnwWbGAMEIFZqjm92fTRVR1MIypa4Y4WBzbWAYaBgq
WCVq+WT7uQfJrb4lSzipOPArq3aqpJVc6HbycqIi2M/82hqEYAFqLXyzKtrCuygD
zoDnnTo3yeIHchDf0iaMcb8D7M4c5QnOuCpnuGiTsppBrYLOFbIpBHqpen/BfdaW
1YSFk6ZJY4ye8yLkcrLFbzNQ/Plw3mSET+sG4MS3LYJnSxrIKTgWoMbWF5VMW9A3
2TN/B6X8Ro5sNWNOcAf1gD9b85xWIAyuhq8MVKVxxyMe/qjWBmNkRc/1vso1fBfy
sj0y1qvAvHQhd2kkE6UIzQ8UEgS2lIdiqRujiJ2OtgFZwG94X+GNIGxEUJ31Ga8G
0AR5XCls+NwjA8rBbjcUe7AlyGLEp+QdvM6DObrVVxT9nK7+3U29J90G7TJboqLk
WD90HO2CwxHqMHlwTT2EZmk2X9t/MOl7eJp3Owh3e3yUSUKJeyssza+X0FKWqGKQ
CDRCCPeiBYwfIt7B7GLYQ/kCEXyNeN0EgAtTcJlhUSo5LgcZm91xVM68CVnLTZkN
pBz19vqYQd2/Gw/BOurXcNHzMf0DiB+qLatEVLNUOdOBgc2wd6/FDLkyJHUIElgs
E/UAnir6+FXMKYR7qodyH/ZCbP3D27iCKnGRYE/lHmd2dAQGgGrw1c8rbAs4hdXp
NTalg6xBtWuw3hSZ0ENaLeiR4QpTKjFsvwfOxaKffsb8tcOIdOkSOUQZJY0wmBwR
rkCUF1n9rVoFV8lMS+7s8F3K6He6+76eFBo51K4xxJPbiq5OLEk+xHSnbHgN7HC3
GBZ7DytM9M67A0NXo1tqGASe5nd53gCNQAXO3RaFIEt8oViIw8n3rGPx6BYPId/6
dfZvd4pHCR+3DnU5MvKqCF+DJXcio2bF5h9+pXqYUxVAJSAiy8Gbs5B6vVsRi16W
Fikv9kX2xRrp+8Y+WkKfuSBPq4Kaoke4WVxlw9l0O7hALWOlBp9mMD+Sw6nC1ThH
wjHAFoaYUVCfZLI+ET7FtlqSEiL/FNRaeOW52kig07WxxGLfIAjQ4WRUoTOArt90
LUHtDzGdEj6XRZSpI0JavESgK5/U18g6cV8qq7ezsJuXftio4haRfF6WpLH+ekcF
TVk4yjlggI0cxCAuHVCsHFIPFHjE5DcT5n4i8ZIzKJGGQqXBlLCR5k52/0WbPcT8
vRxR146EJhqPpMCve6INfudT5bJQVN78KT5Yli2wk8gpZF4ezF1xymTznZaT0yKe
+W7xdKZR5b2XsmDNOxfQxwlo/CN8MzExY9NrJfLE6JtQtVuYueeOP5myeaZpqYa4
OFCEusUrgAsdn7tzQptVfCt7FIh2M2XFQfUp6FvmHb5G9nK+gv5KlB2qHNAS1Tq1
R14TQfmF0PuF/CPBE61crygz8+oceMi6On+yWNforSp3UohApy2qSTBYs/BMm0H4
WsPF/RHebzxYfLWxVqdqsOiNSRlvOVlOJ6jib6+X08f94zS+dF1V/kc2x1MVUQCv
VcaOXqE31t6yY+t80O5fGhj1RtzRCUKi6EI7t8RF0trdnl9RxXxMy5uQZcaR5rq5
I+4i6ExkAh6CIIyr6OMQMb+eX7xc1S4L0EfviwWSt29wgZBZG6hQH53Oq8d16eo+
At3kyL0DFBIQhouK969a8QOvgs7x+P+QJkzh9fOzVOAOCbAhAHh0/R7HV3Lhgvvl
eLN2Eol/NqPmn5nYGb87sFzUO+KboW2L+J2dM0JJI/nSHsOG8LOWctOEQVTjylYT
4faQF2jCykLLnEU6LQXdVGrda72azevcDlGcpxx77gyoGCDe3RK76tQJniQZgL8u
vnaFyB8SNvO+S2wsaP+8BvQcUyTIZ5O5MEgook6Wp4g2hagBwTPuksyMrvZyropK
nMMDZpMVYRyVL7b9qQgEaV+4ulpNYLIGIVUZ7p0D9ctkpNnctiZB3rDorJFsD4FG
zBcwmmFp/tjzEv36WAUIVkn6w5K000CdDkfrQ8+7Sw+K1LIgJsHOSxeiggf9zdjK
eAoZmqML7uqdeP9XxleIP4kRjDxPRUgYzCvJuqqNfco2xtoyPcqikHLXjyMUErcb
NOASKJgZEJAQ3EeO4pFcmP+dJFacXAVkQ9Oc40ylTfIC+R+AyjiEZmjRP4d8WRIv
ud38QbYEAV0NFCT3mmOSzOsO2rwfna0GIj7/e+qdid96aYR+N9/urACxzRVLwKDm
Z/CIm1VGGBE9Ra6sCmmnNcGglFdA6GBB3Uu0IB+AoZpaikiTYBuBoYkZCuxVloXz
EXCkAwqJMYd/S8NGsPewqE965RcapB4f0poJ33dSEEnBVNZIxZouC9hNde8xYbrj
vQ3mgPJqDx19gBsJioeg/Ew/L8iLZ4GMPKu1SrVsFR1uyBoIOuTLkdvtzLtIVymB
K71o4Uysb//VGnrahw7wIOw6jW6mTP+bSKOIId0MA5cUNVJk+dYHa8Ryji5cLTWd
m3ZLZQAgXbboZar7t8gj8C5RXyX8nhLkyvaKMsH7kuRRzxLmZ3Whn49zigm2V73r
N/Vn8B/CXu36z8xFSK0e6ATrxtXMUKIg+Y+rIN09H+K/sPf71uuqm2Ytvd8Qfs6H
enXPaILYRkE2658dQGm0o3UA6LOvfofQsCMVINoSzUztLY0g8HLpa0hLvvpq4kl/
yLzEsqgFlwIG0+5lS+NWNY9EChoeIH+mFZ3iGFomlc7NJ65EYFdO80eYE95SM8oh
VB8hMQUVVe37RwIvD2c1kEb+OnCxaqK2iOBrR2RPBVmwHgzcyfiF7h2KHSqFHQp0
BsB5vzBwoPq7OOvVWt/E+CP4pi6/7XCDpjq5V6+A1tEQnnz8kcdvq2QrxWLzA38N
x5PdjJjcF+Q9NqLTkAPRzDNyvDLbpvxIMnVjXj+HkH4SJGoxbu/S2L46wA0HpkIP
zEHq731OJgpN0pbF7JrKMOIFYJVaBplPfPs9SAmntJKCQaj9yTcmFF6OOOFiysgi
7QEIgGPVTRD0R5YeNFHw3e9h+JruDZ1gLYhtqixegEYab0BQxhlrf+4wPu3D2c73
YYV4xZEL3RsWdHQo3Y1P6JCnsQ/xnk3BVLLjchjxsKBwPzD/z6pN/wKRRi/jj4rv
HqPvRqXbtEUah5M4w8w7A4OgWSdRtIlY1LCeUppJ9COAAjUm/593Os38zhqsiL3u
/WL2Hls5ARYvSbYbgt/KvWEtmu3Al0UL2iX6K5PM2/47w1I9UxKbXyt9xRmYs3LT
s2iJDRAsNUI0K40++A9AdfpA3OVKielHI//1B669VuCP7sHGeQAL7g5JWxz3++Sr
X5pSOw+lvtLXaJ3lHkc/BaWNo8UactlzEu5KE2sk3/EL9SfIxy/nWJF+B34StcRw
Y6QbeBeWqTUbo6mWGZ2zRdzI/XmpNUfVcwaBn44RRz0nU7ElDGoKLf9jHb9IuF5b
cbl5bf96I0Eu1/9dVKCxLEm1H8DiT3JbvGIg6vXznmAUIY7bfjwanvPny9xJCLF7
YBMuF86nlUKmkS/mS+/0jNale8VrxQ3sipLSHIuuTSqVbgCPy3mOv4ryrE8Pc7Ru
HBFvc6eBe0TLa5A32C+dtDZcSB7muQNsXSrwJ1OHW0NnTb3fbscfWq3jnjh9aTfi
4mz2cmMyH9fc6+B7/IrfkWqhkvH3GDjqPPXoEwxjIlwAJi/dlry4sSNKBGjsqRmQ
QquevWgZPsxDk29iogeaxuOGnvEIz4auZHWB242q3JZ/Kh2xf9/c573lP+qvsTI+
iBod6BL4JO5zdCbQTr/Eemkp0KN/epPdyHtoUrj0RiYm/PgJPXCea0X9Y9Knlxm3
We4EKqcdW3uUsdifaTEnXvMfEfFCMuBNvQLxmj463t42NgkgFpPFHTML3HJzTrI6
UdmgF5GNxlsr/jFv744jFCgumfaPjjxTTiL86jda/7i3nfHzhinzI2AHrqvDNXda
JX+K2P76jchqxTcNmwrbvep8IzyMBLEWEDvI5SxtPwsz32UI2Kbo/i6y/yLzSAZN
lSVjIPhvj90XZDld/ljFJTN7hEu1SYurJcovbcJtNG9kcZsy1qF/WxLl95xzLdpL
t3HjTsPgFBT79n2ccnXVKKUIicxzFe2oV6QWDVGQHc4B7+SE5Py2LA3s917+ZHlw
PNYsANyUhRiVRK5c+t7w/I5i4Tnbj00kpW4diOv6NPaW7Mg+wqjRlFq9aitVXQec
ZN1q1bOW7lxjw8+wZIKgis7UBA+xi4kpz2cL+L9hRrzJHleK7q5mXmEUqytO9Ay4
f6Sp287fDmsHB4n7OKC3MTeApKMj69HGuznFPBAO2UYBgqxsf+/jG7EUHsd/aCzx
bnO8brigMMYY2hnal8JTwWbwIOrHd8NfRGRCSSfNqTkg9BgA2P3Q08TLDvKH/8zM
MUpA5xGobJa92HztfTY6RqA3z3uijEjgmWwVm01rL9HMEyECLHfkp1x9DjcemjkW
9wTqUVZxS9RjRVQbrEFMTwcJWPj4OZ1qqrobMmtwA1tDb4/+raQhv6DSWY3yLYvC
4MVAsnf3o9HsUNJfOGIVPCkZ/yvT3YVepLfAkPTANd0Iip0guuYXyl87sMAmJDXT
PKQyKXhIoy8S0r/oZLGm67ZQ7z4YmeDlYAVqlhNQbkj5WA04MI5AqA+oNR/QhujK
6rWWt86aIC8VSlDxF2XB9T/Q8qNSXa4CCoSH4TuK+F2MKSsq9RCsODa+FdgZUajr
8YawEsQl8VKJJx8pQ5fONfaRi7y7H3asY5zT96GhIngINlVF0cyn703q4NvOEHzp
pf2Woy2f5UgZdFOZoxE8G8R9NjkqiZxJLuPoLmMRxEXHOc3EB/m3T3v4ZssvFAXP
mF3W6dreQBs6z3fGMwyMyDGVdo9lqr6DS/YbN3lyEedN9vA5kqdBZ4uah/1+K1tR
kmZRo1DWNWoGtf9Qk+dC/QPDJoH3DgPF6vCVAkzW126F7oREUH1Q/8J99WZv7hXm
aqQe56mpco0FyGYPSyIG74rveFYfhYAJlcUUOJcOtlwD3jqrn/1/NgojPQSTwbna
H0sSbWAhzSaPm8gF+gSNp57wj4pwHfaEBAqeFPRSFqp9Fk+2zA34Efw5hKLGttY1
FOVRXiIPMl29xl3i3MwDwphnT8Pzt5+KJCJ3AU362tTUiFhU0OmK2t2OALEAcRyX
xAQrllG5WaY5FYrdTgU3JwQ12mI8k76czYMfJKaXnC9R2XH97GrFsPrVqPRwLnqB
JituVZEHAxM76IQWbNIR++VhWZsUDOy5CzP+6vvFZdZBgUisaIgh1xHSvdvvyYhY
xt83aSAzlp04OqqVoYzq9ABwsNNJFGhKA/qWO9wCF+uIJEKJRSe2Ef372jshq0eM
d18GGzmJ0qYkcFOzmpU0gyUsuFq3Fvq6m/z8411lj1Q5w9DNIxN4fpt1xCDwKAif
6yrTWF2QwCBO/Ct+4yl8pP0zg8r2T0MPzJvZ61fAHRF3cY9attkozo9t7cw4nTcN
E8Nm6wfHSWLQMix23+iI1i38hIT5iiZEHDGgY2g37pGrHiU7wegRrrkLLNy0r4Vi
ttVT8G06+OcsPYYTPrDuNYuSbhXFAdM/e9X6/RUtcL7FG7twNYJV1GJ4smtXLN+k
M7CtI3TSlKwYn3tRWqlfDJ0o0O+6wvzf7neUHsw+VFjNHPkEgv7wknog7+SNAa96
sj6Uuug8MSVyiICdpSP3HhNlzX28QOEg9QNkqyTXUDk7AZIkdpQp/UYRcmGWmYsF
YUBt9Bi3xl/rKdy2o97zQNXC7GHxtbK9rnippiu+t4dfPJoguAU35/iV9loaoFhf
UKdDsWXiwrZs6Tkrh9PxNAK2ZWKZJbS0i73CHMV+i3R9YDmr6pIXUNnWl3RU1/VB
vqFhenO9aV9fjnyqGo7bBljjSIABqO1vt6O5XyiHjk+/lCKr27Ni5F+M9uChGuIt
vLfvI3YNcTDz4jKX1ks0ZcH9xC5vKyM9u46ZsrQFPDKK+u+T4GgaThMC1Y+awKK8
rsIZ9RhZaF4CI/w3xuDCJv/9Rq7LnDorODriJh29ShXLkDTFym5HQt8RdT3xSAGj
XplHtvxs8XupJzmTFn4HfvKdCghU9ZgdYAloa0mko2GdtRKIDTJ6LIDlGcovVlVS
L8j0A69mwcPgIh/wKzlxA4iUa0eN8tqz30pz/eD3+VxCywBH3lWIsNty8f0AU+0s
kuxFSAiYTljasu+dVmdWXLtExQtdeLqbipZmY/poDsn5DpqSre1LwN9ujnHfQHSS
Vhlnr9i6cPT1oXSned9wPWcrkfHrzW6tvIL/cOTRoSlmkXEPJ8x3PLFdonOIXjXz
m72WuIUpIfGdyq3SG1Wlw7G5/W5r5ufPf2pIrAkTYgtwjudY0/dfKxDxAwHp5S5O
SOrKWFGBgCUDwTyXTBMnzIldkDodyMg+P6XvbahMw3l+XLdAg0BFEKa8QqAup7J5
/UVS7u8qdsqsp5C47A+tPg9pTvr4uBRWaC6Pdhq1sFD37RsR0FVrT0ET1EARNt6b
sf2wZrKRh80k7uTUjpHaEF4b+GupUOQMtbu9KRp9JQ1MWcS9dWajLJEq6nanRrLJ
CkxPwefp0bqNj6GCGRd9QXiGTPgrUp7i+TwTdf034dMSKLld9fA2TawBJ119zFyu
OkdGN8QawPB0jKqFg6fbimMNsYX5xRdD1xr8ftSMBRxGh8021VEw4MpVnPXQKQsV
L6rVmzraTwcedp7H4lVsDFW03haSms4iVslt1coTE4rjwzHhLQNOotbPU4pMlaxj
MWPSPQpdbZHxxeWPYkfrjMS2OIKHNY+U0eiwNMg03WcnUOTQF0NSmS2Sn1jg4TA7
+w+03sIwiysnbd3b+HgTkAEBu0gBm5RSPYQOvJvNv8XjBBtUSZSNbfEAm5Vg6MV2
Ja7UXHJoHU9NYg+5KxdD3nciOmV5+xz98teMCaCNMTYwBSbJQ4fzEcu4LomBMlGy
1GOFPuN40exrktWFqjbi+Yo0llIzJWyjJHuVzo7mdTzc9TVBQvtkVQSUFzymZZPl
bU+PYCv15gyzoeg/fl3X72awg6idi+gopGam0llvbMjYgHzx+MqaGstyU0omv3Xf
N/WGKgi/JimJae/XboL1mYQ4BGUtptUQL1paHSdHb40KJxwfK0/IdVh8RVaPS7ND
Ct68BVsePowigpLhy9AC3JL9beNdlCqG1TN6FTGwdZkxj6RJQ6Dc0yU5dmaSmfMf
FeYnLbFtgiNzKvE5cSdxApIRhGHkzRyJj5RFSk5PL0I4x/UZcyuqw4NVGYMIy3gb
RpdiJw+rUAXbVRHtdLsRlCuMZNz903VZAdNoi7I4D+cso4khe45INRK52mhJXA5e
So3iVtxOe3Icm0tb6gLUZA9H3V+TZ2tJ4SnhkKExDQp0VjLKtrgTWSsuhl+tN8M8
GrzEZkUV8tMaXpcYcqo1pOUHGrK4lW0qcfWDWNJ+9CMPzrNnDqJnRlUzTlh/CpMa
BzyOMiu4HBpKsfo3YJdQ5/98ZXORlE8yUdOtvgMH6bcFW/Vh90lscOJjtDaH5rg9
jtFhOyjK+GWkF8vKLiOF93Wp7PCSCyr1YcrgUK8cgBVh5g1Ci3eHH29jKYpZ/JnY
ij15j58/PwI3YdnZc0jw8CGHm57kbCT/MseR7QJu3Gu9o0ux7avY0sZ3KUdc8P/z
uAliKbqX+LawItkDlWDjD356jFVUaPfo4Xq++5FOMI0hnlzVFCTdaWhwmOVWeYZY
dWN8uxaX93RppClghmuHCAFHsoVC696B0T7HxxU5sUEEHiwDkAdGCdVcrXTAA8yP
8kRjMvdvlRlcyWGV6QMASaBHmrXi0O64CtuTNdG1cZsj2HXIG2gnT9JidkLhQcic
9vgCWEv7v6L8GJz2muz5X0xN47zUeSN870mEnYhngcYNIxOCGU8+U1v6LxOFSa+A
rYbn21G9kiX07K50I9QmLbpawtwgV+7gJ6YqrnxsY/UnjtsqWBDXoYB7ebXNaFMo
quY3Zx/xcJqa/ESl/a+r9kCYtQ4lbzUifNsmZ1vRXgJpbWvAIixdE8UftNMtiWXk
CwQ5FlhFOlgHjGsq7zL9cWEQDZOi7MqwMaFT6JiLM6ND5mZDor5vr5GUPH07g3+R
359v4aOka716UPedr/FY/zQ9LJtJ3LK3BdJFFZDwWvDfhhB7RU6QmSvy6Jeiccfd
MrRj4oHiZzTVdHhWLtL/p9GNQ5SjgXr2b6wdQBD5RcxzYgsX+0fgCT91n7yu6ymK
UQ0MZpZc6qOzRidUiPsr6mdjUeh/FMlEn2ln6cIzGSGOkmSryOm49HhgJBhvYt5x
Q+hZPhCcGslXV0HuIFz0wjGdoz61qA90RszLZhIUHMLnIUKIAmqI03IKtqqXjujL
n3eEXgVGiMiSMrAmMYB23qkw4LCfzDkTlhuaGd8++0+oSxlQUYhR1uFKSKrltrCn
vCRs3PqtT7/PJQXJXLVHgC1fMxoCYcmxDY3vHwRPlS3TdroWebtc9eAJSBK0ZYv/
krCwBSrp6WaqcsugX7una6Rg7Ov0XNZd0+ZTIY+XEc6I4I8hMBY6f1kmMz2t7gY8
FfPO3hu5qeKrn4iWx1X5jMA4hsGXN0+4XpvJn8qkBFExJKZIgZ1KtrWDkMH0EXJc
dj9FruO1OnnEdO+sEGKW+QlSDLaDz0yu9eseDsy4WlfZbl8xMbl6BTmBvN1DHefs
UJzJcsHefZHxb6aeLw4HwRr/itTntSRUZBiQ4faJvhOHK+l68ie+mggBeTdn3U5O
SgVhXOn/BVGYiGKdLdnll4UYuvIWfruZRe97qKg9id6MvMS7IKTFaYA9X8je6vT6
vA3pGl0pTYX6vERx6APEBULFnJgX91iLDZSmmaOptuYFj/75J/3TvY+TYwHfR9oZ
DueOiyY9O1E9fHb2YR5lxlqhv8xNENBydSEzWD2Yz76D2b3StUMS0N9RTXzdNJs1
WrB3rhS3ivvAv7ZoI6CA6hwwmmKlwCJwrhrFi3yIrIhJ/KPDJ18Rb5TB6XpepbqY
eTrM+5O+z2gCOJuL73ZHA+uCWpiVVtot/ogSmcD+29Oxg6tGVtgv+GZAoCpi2dLW
nEK/yPcV349D6FDgUUyS5HisVVo2wgXa9PF/39nJ8yPxpccm+WYtTEZzt6dj8cVp
r9Bov4SGxor25/1a0d1nwUfBrR11c0bKMtQfjD/o64B/yqg8PlkZWs4qZWAlLRlX
o01kQ5ZIJ0pc7kPDgs4wY+mtO8L+KC6kuxMNblxMgqKe8/0W8Owh7ohaDQcrKS+H
DsyzdnI5IQJu8gYmJhFnnR0kpCpcgRawKX1mWxLv90b43XO8pbTmD2jv6k4rdPOT
FmVsnGOezHd7hQRX5KhzeHRPQlOyPrpGP+4Q+Qsx98w/Uu0Ut0PwvQ4/p2bOXOpo
Aau+Iy1/cD8vMV6TQo4IHjsRTyDney8RGYEEIjsizTI4tFxLLjEwQqhq72GBy8EZ
UnG1UWmlsJ5IkAG6PjbmJehLyS7dXexwExzuGQZSBlI/Skd8LL412me9YxvSsZN/
iNMUD9Bj6ORnYnBHM060VkX90WL2ry6I/tzWQPrgvERUf//8L9WMZaxlzdcJsO76
O2fayFxqa3BcRcxSp6TZIF4spoxB8wYy/JSY+YPwtjARmiFyQ5MQLW8trkQ03B+Y
zTrqW1KmjMrvo04dwWsX/YDw4mOP5N6M6W2CnVPPtRi+bg7ywSvSEJ0wjfB1JG/7
INH7rdRljgmK/LeQk9W3G0yYIIijfFA5wFt8tvCj6tNcjKdqT9az9Gt4PAp4MAb+
A+IuzgtYwrdjS5v96k08OxdVJq4Itji3LpmhEeqCESlatYCY/qxXf3SndDabC6ox
wkQ6NXuxtdRbFKWFcqnuU11+JteyZrWO8eoeyggoxlLIwY/kBGRGtO6vzVYJe4UQ
iZQfzUQNriQWhiJST8UHodgs6xnCaryQqSkSdhJWfhNspnp6dKp9Ep53gTRKcQsn
mTplSqnXln9FGEqGWkxoPbsI33eaqbcba75aZ8JDgVxMtIHWRCPjAaycUXP90eg8
xAQwI8/Qtom2AJRoX4E9J2ki2piltTXjnkkd1Q3wvWXx6gmynMPpThze6Rbcuo9j
rOh652VPle7OBznNfUhZ0Uh0sjC8+pB3Jd7oJL0k3OYIQN6d0rxKETYYbkc29hAs
sIrNi8dA8EK2SMeNpDIvGl7qMP8QBTfLsGwoboyi/UfAI2KBfD7gGyGrvvAqFtEz
5gT9VStiqNDmyDAjWrbyo3D/v+VJ8A2iLXsEw3NwmfrypYOZUqLN9qcLOjL4qXU8
lh4ZpeadRMcSPc0951P0Q0qsaZmKnbGBMhavP0BnxuHgVj9TTcbHxVVvu/+UQH0t
aNEnCUwBwmbngDEDNwIF0Nou+rDxxt/nRBRfvKZVvLfugvTyMnU5QTiUfEdg1vLZ
Vb1nKuFXFkYTgsmk6gzrObKNewCS87rk88Dpd3YfXonljrWyIZX7Yw3RpqF4nrnF
KCaQ/IfNfTefK1prPHfWKdJc3yFwYGoEZqhmfQIJNecGWuqv0IiPMCfphMxAxPhT
fGJMs+MeQWQYAAdpyDorGadvSlp4FmfXBUJ6iQAN6YioKtbNMqQerTmwoRT8eShn
E6J9+Ed62LMy7yQ1aTijDkfVmOsKIcoT0NKLPemNTs5oOmx0pmgLgAsyuBlihf7/
3ID2KgsoeybMO8LGUpOWORuuM+pM8aWVP2aqE65c0F09PvwsFrokDoTwVvj8Tybr
1oj5kMU99CA6eyagn2kunHVzM2MdbcuIA6j7PxatF5K89XcfMMz4aMYO51wxM6Wm
9ufmFbIvWNMMxvVSfMlvQOuGCbh3weyV+Sri5FNm5Bfcol/At2w5Ecl1YS3cYgK4
9hd2wTsdNVc7J2NMNhCGgEp6eIlSBtNBys0kBFQRJcmlku5SxTD0ePxQgJjDWSB3
0Bnc2MGOSu0MPwHjEmRm+ofDMQ3k5Yka6YEkhctonka/WnUmx8Pxqdrxn58mvIiK
23oSp/XELU4OoUdez4rZ+u3hKdDYxdk2eV5Q6Xa0rOuJ7CMOtTlBkbXDcKf9xaPq
cVqPE7iDkRqppDKzUIOmNHvM5mAubRVG0HRyCox6awpY5V5i2nMzfGKuus6iudbO
5eWC5JK9NHYe3d1npOHp/4j8PW7AduDEUM59COJFMfy2ImV1ZK3B1B1ttgPMK/aa
sAo7Qws8RJ2YvUu/qBjKJbBk3zI25AAtK98MWjZhsWdJTbZdZfD0gB8zJn8aguxx
UU41P7faBQUY66uOgEltrXED+bb76mS4MMechkxf7GDghAuJe59qlrIG/dODMCsS
hkuKI0bztPBzGdMEI+IMrGmkCEWXmiZb9dfCiZEqQhzmkzm3CVXspZMAYhCqfhtA
PhUQO3lToK+hFr4mAtB4YbDcN+xms8JOOA7/3MImFxUMc2OX0yn8Bg2uP0a5QiDX
MMGhoIsofD9h7pntGMkyDAMGL8HG/wT0o6bBk3juXGdybZ88n+5jehEVQ4rKnBNZ
yfSzQaGZqTEoXjZKx56NHnAnTRRdd1l2qyaN5pfAMjylcSV7uJ58Di9SCaaKMfuo
3stMWrdyghjdx9LnMAQ1KjpRGA3A39uJmL8GCikw0eaH0SjS/gmBQ3DPod9QBRG1
cwN12OWMijQaeDnIQetCoxSA9x9ffgHbnZFe44XsZevf6kfAilt8l5VT1borgeGR
c6ftJLZwc+nKoJTlFCdjwHr3Yx2K4JlqeB0cpmttXKJnxe0rhi0/a46XeZQf8BUQ
MFIjybV4SppV1B5sjcG1vue848zNuP8pTqh5k/If87FBvbBQI1zjCS8GitwdwQRu
AJv6KCaWc6gWfVGwd45u1sWE+xmPWaesJE8QGJfrQKpVNOg5V1Ok/VfKTbOL//A1
wxwiIUtSYbHaARhxSmlO6cP+181C9E/PWPpUvdp7GSVyJOXR+qlXxnq02gWSlkDz
3fjjWpmw8XTdXU4onmeagtrtsRh9KM292jbl3sYPjWLEdJCAFyfZfKZ25Ju1gnBO
6shWWhB8j6CFeqKi9YAXEsfkbsiU3ChiVWasKdKsXTn0JXj1IwocH5Z13LK/ddS4
b+OnJ5VoOuL2XSkLE+N+QCC9We1xjVeSMBwB+fX2ItiwuLcOLNDY4E2vi3sfYgBm
4QtMzuCTv1/KmB3ecNfZtTupA3xZ6NQfm5cw1CocOs//5i/pENLAHXr9Lk11pS3v
jpPv3Utl6W3cN1rKh0A+WRGS6zI+dV3M5ibx1a4UDRewHx8stcdesO/AQfBJTMEN
+5P3f8KcGAz7rLqZUlZbaV1uU0/WoGPTbk+ZD6Qd4vemnu9BVmo2aZ1owcUBmoD0
86unzkKp5n4vgrUa4G/g6xdZnnjPmJkuBdSrk4LJ9qV14qpMlXza8Qemmac+QxK1
qNQCh1nQnwBa0p4B2D2Tojtjzhu+OD7wVqn72LqIjmFEvTiHwkwMBUjb96sDElzS
SF2WV6QV4HqI1dTe1PpD5yx5xjw1jR0758OAo1nO5phW9uZ4UNEmtooBAverizs5
llW+xxVjvbqzDm/UVc4ZFzg9lTZ80GuPi9zNwAWzwKXpOIXxz+432E+/Kp5Oy/0f
FTw0mbPnOEQBSzq985HrJJj+foep+YGsnANf0aMiKSccgiH1zB+ltKYLIenFLttK
WHAwm1sIPXb9O3lOReaTWfg+LPcO8i7MKPWMG3NPAaXMldoUnGF5gdw0GZIHIkf2
D3jBU7Y6bFP9GkVBAdNoWPIrg1oF426IMzGVXULllS/2KAfziydjCVLGBtEbXjbE
DxTK5n30XnRykQTsnwIAyeCoYv0RSqmGC8VUSj7srfCCyjjVpM5KPPjflHxUM/bo
bpcDUzb1dY/2FwOw6arcdJZeL6NBvb8tKQQ82tQff8aerodMmpqMGwLlZAsMesU8
Lcfrvo2kDwOb47BX6xAywB7c64s8eXqWU9KL1tmkFzV+fNH4fzsl1zXiIGzJDjTR
p3wkizIZlovkRgpdebdmWHvHLyR+EuWUvZGR63aStbZ7Ou2DhozY2B9ujj4rBc5q
sR384W0I93oJWppzIc3WsQNa39kPYcpm+d0gsfwYIllQaAtiUPSIl+lZNUjl23w7
gtIUAAkwCDe4idWGTPcI+gRw3GdrUswasMOT2RWaeQ4XVujAdgmwFxrNplshY9LX
LmFbtTMNJK2oaCMqbfi8gjsDWIqFQup/vpaKMh+RyEeoNnj/XjHbmX0vwHgb01RV
7O6g6MRKwDQdid6gkZRsORNNXqba90pv5C5Rxyo0dsc/awFxZk+LqbUIbJ7zEGkA
kvdffxLp5D4saaSUbQqbnCgk8ZwWJl0DsOR7/L5/6dYYibmdkBa5gbAgpKAY6aRN
7ROKFQ6uf+KzI60gLrUUZNymVicmQutZLSHcVZN97fa9GIWiZbXICt2RPvz9qUQE
bBKRynbxUKzSq0yzCmDUOXdgy0zjOcI3dTASYDS14Buwx7+FVklkxoCcKLGv4Nf7
E3FAfriQB3SYM4wctG4qDVzHub0duAid6YKrocYWu6z8Q1pglX1InhjNunm2NPAP
GGBrBD1PpygF2zoXLnXryhIwem1oPOYk0CXY7ad6jrFqIaAt8v+lzgptcVmgEmaK
abjl89+3Ombm3gzV+qkYvfU2QoSzJyTrpY5JMlSivsOwPfQlfGuah9tFkLUXPISz
oDpoVWhDYkxIFXy+ve36f7pNm40d8ZJ4wPaU16ihdVyKarnb6nDgjGdwB5Bt2Q2m
llnC4oIfuiF0X+PLnBgWU9yaDG7rFuBUTEqgR/NTzU9jxxls+jZ6sM6YaiVi4Jxg
K6YxzjvqW8j94t6UL67fhi61vAnHykZI/kfqbjjxTM6B1ARjNuoSJexMrYvgtsXV
UCUawsX/QaqiAS7PVtasyyZr8WaKU/+epBs9v+RZI87xpHPsMJ4ZjMxyRlJwKKDy
xSfRcnpiV3rupjwm4SNLMcyeskauQe+jsPcm5+k7zsZPRoxOfpP69O4GDVktaQYY
4ezNsBP/SCpRjK24Cc0t5GysftZVrhdHRLDmUbJQN2KZiCYTwjGLN2UnnAnfIC1Z
fKvU6b4CS2tEYGm6Ncm2ZQf4NN50GnXUyGzavr52RH1qmg6bxXdo5coIe2MqA7UZ
C7ja32AjOCHKq3KrESr8uAdzSFu+L+sIVA5jXpwL9zdljDPfMOYHv6qWjWRWFR4R
11nIrebuftoCVPDM4O7176XsySba4L3TcvNvLCDPQV/h04BbK9HGSibFja8lQA9Q

`pragma protect end_protected
