`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
gueMR/J1TQVjMLKS/u/V/AO+bX2pdSHHEFJUGC4jHQXiu8gbhwCqNK8IqkHWlyY4
HC8eUW58R1O2pvHeZiNJnsIh0xhw+9qPdiqE5mqaPE+3/nZURqMUh0fxye9n9uqN
Nvp7BCCpCltNbC0JWaMKdFDrgdmhDQzFFY5opkWK8aE=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10736), data_block
G8y7AlR8Un391KY9LuaRwFFbMPn+5iNffKzzgAfyj59OZk/+77qfcd8todaR0FIp
AlDV4pLRi3HIgJ+/V3EMZAxnHO9fVozfyDxiYCHLVZsFb5y5x36F1le20tSht5xv
U5ef9/9DGNxaX5xVXdAU08LLLqMdNl1ZstHQGhhbpYp0nFLjxiAxxo4rnNLs9UWn
1V5yPydXsORBEQD6TFbQCZitE+d09m9+sDHpTW5EgoBoqO/V9DoVQbx2CE70LDk+
lKYkorA9CfWWIt/NmoKLsRxkd1DwucU/RgToRRtFYfCGcwiQ54VVZj9IvKdBvtIz
lYz6rMMdesJclDQ00lSsUnGX5ebDbrAHBPxlNXn7iM4aa2teecdwCdILFcK4r9lH
WHwQ4f3Q57kHNQQT+OVWTKTHis8rH+ZxKfngm7E9BLYlv9BBK1T5RfWQ3VlklMsq
mgD3JmhFU6FTPSz2yNHWypV9fbkAaXzs+2GDKBc1JeW18uH9sNd6I7KFC7rYKHhY
1XPJeMbLbREjNetPz1WqHtMfhVDZaXtSrRTo55SAVxhHpCWgUDyXZd/iQuQzmcB1
8WkybCMbY3jSflbjEgBSlRJE3zmSAF6tWhl1pkpJve2pKEAjtcV7QhTD3MN2bpDn
dmRvI9uVB/NWRgcWvjk52tdKftOVnz9PN3tCtYFcnPJESYU6pkSXfbtJstPzy16q
y8YK/iBFRqSWVMJIsa7rHyWKx5B9UQU/ACLs7ZzYAPa+jJm1dnNF4p4FuX7pJJhU
YzsgufcmylFZZvjign792vEpqxGiTtioGgyucqeAulEldbIJ4MS+IW2w0+3OUpuo
UtnsfoEsYIEp6Q5Jm1L8BZsMl0uQ7Clb8aUfPAKyN2CCBfPzSaV+IEYp+WoX5oAk
K0zM0TKHXZ8H00VrJNXHYxUSjhPShIGKHMd9VdCFxvCFHaSYP+VrvWarUTM4b0O1
bwVVlkIViKN/lZwP7qvRZnYL/fPfjlozIwSoqZ0QZkhZYsxnXu4o/cwBC9GwCFGv
I7MkfWRRBB7FD0YkXR6UT1PTDL3KiOLrKzfXWcZSmuzQYM3MFP4IKmgtazLf0LpV
zo7nQXPXWGnv9skQB4tbnfDTvc4tMbnrL+d4aTWNQ4NPOuGAbt6qW1S+1GF4BEOo
DWULjZN02ze7t0RS6tOh+sgyeN8yxvFDDoc0eGi8kfmNXrNQIdanj8B9kvFSP8sM
vsc0ER0BZnzRkrKK41kp1RO9mITllr0217hkyo5CZJZORq/fDNst0fjafi3iuC4D
eOHRDFIqNt0rxTzvPhJK0vkmp7A08ov1vfQrfxYHCAYeohOcGluBqc7UF/k8PcJ0
686AjZS9wG8SiL5KkwdxXQhx2YC40oyQ6guWh8PNEyXehYFoGH6OrbOoro3+PSs0
0ujaH0xsQCg/8hLUOGl3Bj4l242oFPp1viZfZNR7d9n2/O6gwvdEallMCjuJ4+IF
zIeXNUJNEgNWEhBfx0ilrm5/vtiTKF87dNx+tGbGMx67XZttMJWFKC4mjuEHkKHg
Y4bZqjZ2j8YDRS8O+2eb87Uooy7DgbLUYbVy8B7er+4KrK0e1XDT0v9A87BmlfRR
fwCb9CydDyhKrjAoPD5wNUFA+Wqh3Ahjhpn7IRggQ4bfrzi2yNDg6rSi7eXsArxd
gBvz0pmes5M2/iyS8Z/ZYqyql67IMXm4b36x70u5dfg5xlanuLfGXJFMts4zoQpP
yeM/cX19+z2sBBtz21ZA5dCpgiZpHYQZu1Am/YfGu0AHNJJrJF1Ja8j1rJN/NIfa
Q7NvcVFM+IkObTVuAYo+RYMBEv7k/F1uo/ok0OfKnCRGvqc8FHsmDQWbza5K0lFf
rIaOXDVlryAROHgqtbZNItcEh1TMNotOYYv+Rk7nD5TaW6pVAbf46BViB6HXOHe9
UkIjb8Uqu2a9URuuTHBrDUr0lqLQ4ExP2YazOtaLqaymaDGMKvNfhwM8JHPiDue7
D+yfEFVNWlYfvhYtn5IQrehmyEg1pYS8JfZc8d8BL4PNdJQf1D4aWIA6ZOljsbrD
0BXVa31nErjpsZeC4ClWmHqfOdSp0hJ9zJffV6mHzjHbqvJfIROhwrCqOk6c7lPh
ETX/EYmC6D19YwFe/eMM8r0WbO1XoWwNnyViygl4Bi+btfJOEU8R+i6Ww5RVTWyA
X/OShfE3JzSFxakm0STNuSaVSzbxxg+7JukOcMk5oaCBdOiSsnYgxpDdIwTBq7VO
MES6qVQnKJT7H2DnEed9oce0/CT4upYdbGxZzKzSjCLkb/5995YLg7CgIOKeDpaM
eGKeAUol0mpM/AT5k+MubFN/ZK3k6mM9s+Gv5J7avyFE5NsjYAUpIZ/6rkiy1v61
Arvi0W/cm3/lo88O8AF91WjfGftPwCgRkQjsPQ/Bq6HAt+UveID+v2gynnKdRcfz
Jia6Amsv84fpadpe8KbHikXIkCUXFGnw3WVmmGFJHQvYa/yAC562ZQHk0lhFDmFG
uq4ZHz4qt4NeTbWs0ybMJAjl+dkLw5bg0uQ6TYtZVQo2+Odan/A6Z/pnhGuM+vhM
1WOjqJd6AI29PrOluD4TQMD0Y+DdoFb60YAaWXNbwhvB/5nkmiCm38S1/Nj1wYFm
vX6p97FH+jxQeO55YUQMSyPir9v7ZMVkjxE/xv4+11kL/26M4SxZExK4Kg+Gsm34
VblDoyGAte5FAueo/XXs11nY8P/KJYSqoj3B/Zvtgf516zeVaGul9Bux1Uk12wFZ
5TYwUZvCR6SB/k55ko8msPRawWS/RT+NGLH/oWBfZFy2bKSHLIbuICav0iYTCRi6
tZXS61rdkHeUIoUMbrzDXIMYbhHtjj/5s3BEbOh8VS/ToJvE/KJ7I1dHpI8CgviS
Bfdf/1vXnGCkGYonY9D7moIagnf64MVtPXEAmmSnAAYswI952uhxoKIb2KPqkAX/
yJLCTsjX+e7qsosd2tdgjR0CFCbEU31rRnRFNuwP9dJ77GkKHFRYdQ9u7lXP7xWq
WVcG1JeP5tx9uUK4FfTW2n2DZ+CA4+d/Z9xj1g37FcGaLimc2z22QC+6pHWQ8hY2
j1Dg7Zb9p2nRw1nkOqxmrON44BaYOq0bhHaniq1QBPEbzZuqBdDAJYCvTB3jGFPg
K6Jh2lxbUmBqSVHQGpNS+dC9+39yiy8JGodiRmpeqrw3vp84bxNsFSBv8SMiDlt0
oDuUaMr11vhOBjsYvvzJAb27WKqCwcizJLuQNzc15GqogAiA6AO6JKmolxAxdR2V
q+U+e+zQHiLLbmvdT/REKi5MfPmJcYQbwGN3O65rdD7F/oVa6b2kwOc0JYbVgdQm
1xCwxlSwbQY5UJex4imgNldwMrR8+iGDK8fz1uc/MMOLLqNXN5c95KuVpmTIdkIW
/+zeCf7ZHzJeo3GghSPv5teEZ1PrkV4taTz80X1jKy/yoTdJ3wfkx9l5OWhdneG/
xJ753XyZPNgv9lNpTu8sC0RLvsnBJDLvKAj+EPtcMQxENMqe/bBTPzGd5CFmUrCb
R5+FeBRBhjyp+KoOu9pu1srrSjP/G+ModkwCg8BOl5SSalz4kYNVNtepZnpvWzqJ
IPgdz7DEzJ484fzN1dj0mH/nxmHq4BeB5f710FinbqvARYU4CKJbyFxovlsIcOVX
OCH3cfEUFOmzfw0IcRYY3pIrHR/oEJvvsF9f3JJt4B+LTRpL8pRFvE0XdqhsEb7Y
lMgx4ugviv7oTxJUexgXYq4lzap0Y/c6+EOUMZ9DyHAqEsvPlzSgLrCvWNFJm4Yl
gJFDZ4dw/dQdilJRzHYDuJZYyV6QSLBjrGPI2M+bjPf9t0iH8U45u9mDf7jMPBq0
ae6IJ+JbSmYz4OZ/XlUE3CLJxJZ5HPGluzpFTi9lcjYBF080HpHwivhdcRWdmHtf
OWCiHGZZ3UWpwL9Vu12ytdfxlrSHdsQM2OhB17DH+XeUWeSujKqEgvltDpzcUt73
Y3RAOnNZvVqZxIY7msGNHEkMHfZEyh+DRa/cXYezd78lOE2pGr4qJm8spXspiqsV
N7RgeAacK45Yj6xcgokJlb+nPI71SEC2/m6RbpB79IBIUQ4IXwNZAemKoQUvTUGw
WLoQOhFJlkMcODqic2AQDZkSCLWJeMa7bi7EwmXUT+Sd5yjsnC/8u0H2COmLVflt
nhN2gQ/OoNOplpHsXsk4SvxR1l581IKN0xvf2Bblt9sxefp1xf1cOTS35fezf5/N
/KCadsnPDE5ZUJYouJ8tMmSpUE4XSKTcWP+tIBegnBaZ1KWIYGX82Ozj00Lp9/WZ
EX1LmGYs/E8n8nogMGWWLvIWmtVVjuvJ3givX1DywxzNMr4ByBZ/CDBPobbH+L5o
7LyhoumS/urPGxb+5d90j6WF5FDzuhJfPn5Sklu8AUKSkYOf+qEwka0Ed5sWhwVr
3tT7td8LMDWe9SwtrBafpEeX1JDVn93f2v1NwfMzfM1qjaQkYu/iGvofKwODzNj/
4U7q+pkH/LNCa5V3ISg6OlMoWYRQibgKbYtAHiJb60Rpw3JuHNBd+JIW1bPyiZ/E
ZHg8pdvOT2q+r51JLizEcnI0GJSjAnoqNeLlPxciOI5MWSV4memHnVFOxZQdSa/E
fLDbutPOruU5PJAcO5FPouWcZNPjINSEckNbv26RCH5zK3jnrER9UW4MSuR8/YHw
NCn7YUbRM2QjMWog98eHXvk46zUaYK3iKESpCYCVMdXAyMCgWDIm3dLH47nUxEOx
F6D994BlhKGZhhCQD68IHeLW3ZOcnmLjIi/CclQa8nq87Hsy2G2uJvX5Y83FBJpL
Kp6K0J8HYmIo4oe74qfthW+ZTnD1+CVE/3SbznFZf0PPCIDg9b2jdi9lzwKFE3F8
6gjFu4QW6P01Ayl68PpGY06W87e/HpvPIxwuHvjiQcB75taAOCOGHqF59GnJo1jF
EMhWI1v72hUG5hVxO3N44V7koKjFNdat2JOm9sgr25cOaUR5D/E6kxWBXQwrQRtL
IthVP4ibrz+XjHWaH35I7Imk/sU0589qKebO2N2icZOY1pJfpFIHWXybu/3cYhec
DljUK4B2M+MUp27IF13UP20hBK/azjpOcLut2SufU4pwTQ1mNBqDDNDO/nXyKoLS
jDueGL3QPmBdomah/Pa4jK20poUXwKu4j39hlnfN4Px8MsmoN8zMqIbjra61M4kK
kgrVjH3Lyj7lZW2AVs0DTwHHE1VW4RWNNkocag6H95yjPLQP3TJbqbjZUdf7icJ5
O5Mie5l2Mffme5N/Iy/9TnGEuuaAGh77aRjMl5BFNVNS91UQ8/KGD/SfyPrcI/pF
3TdFHDZ5fpi7QHwVfKyHkMbCDXYcBlHurpKrignrC5J3CpxjWnJO/TtbikTJnDu0
rI/FNyHcnR5OuXGoxR/wabLpCu1u+tG4W681tZLxxw00jH3sLEUfj8FxPFcHBytM
MOwC9liUUD/vX5QZR/d1AN0Cpi8IdLa8XdZSaoFwD9NqJHK7dmS544mc3mCMIiUe
WJVur/W7F+T53YQ1C35tu15SH4Nh06PBLBtKe5kLrsNGp/I7q4vaeqOeli6cGkeQ
iLzPPyhoAA9d7KK6IC/+0u3l4stvJ4HSK9RbaQYRc1b3H6+57eT6e/iALQG4ckrQ
HM9g8R0y/mIgMYA06eAMd/X5LEeXbHB8/F1xsIhBZHy79Ul/Hsg2whtNKK0NBwS5
3vWSP0KXrRPUpgPwg8Jr8l54HGX6nWD2c2jntGhUrBP6XsLkwCHxBwerhDta26Jw
PgFOx29O/8oSUZCB9eINHijpAUy9fcNtvIuCatIz+KnbUkkXvaxmNp22Bi2VQNXi
Xh18r8BU3Tv0h84gIirT8TrrkEEqD1a7mcRq+OD0favjiIVQl9Gfm5oabP/jB0sF
8BGUmZpVTZ6lWnLqfbTIv5bTszIgPNL2tBsCMffr2ErSu3dTN0xSRV0Nal85pr7g
xE1JGXT9TKXxkFcp8dW7/4VRDlIstF2x9PKViQcGdqAo2GDZ8Y1j+G+Maii1y0uq
RJlDc/ko4azILKm8vfM1mt0iptRmlskspvR8zVI/OBB9cGmibLFFLwXDctuCgLlr
AXY3fuNnCsGEbtx+4VlSIIx8Lt+ZyGv6wtxeHFbt9QYOn0e7AOpJXb309bePfMv9
SZCqdBRG8Agr5cJfmqlGwHC3PR9uINP0j27Q2X5koXC945V8dbsqcHJboG+J6z2+
AZuNaBOR4fQXA/p/lciG0VaeAOxEYUskkM9Aq26TEhX6x1cXN4QseyEZYlALHdke
nZtDTSem++Ufuj1aFODnV+IQj08G6nL5BIXJH6mOABrXVrJPWN1rtAgBTkx1UEuf
ZgsZnkp5oQeqm3RW/J+jpqHJU2AR7nmFDj/WPJOHOGfcQ0utGHx7nnxxujangezt
8jo8bQ6ZIjZ8VAGifFyjMY8njssMwM5mlWpyf+MgKL3F7feMpp/js0yI32vb8i9P
qWgPmDAwhshy4zeJiVv8Tjep/9o1clMZwlyRWJpTrbLMVxQ2BPx54FUj4jHjpHue
BUEYS80RCiyT3pnpu8Auj1RNTlIExLeanUXkMB/ZFZKU3gunqcaS7dj53YUDffRm
61V6VobOdm5RDQEQyuLhfTZN4omP+sIslhetpiqbI+qL4IRE9LSVMdLN8eVLBD+z
jh7HjU8cSMbNb9oFfJXBvpBZT0Dqu7UqFRMqSBoDvFMqZhsokbIvoF4utWs2yMO9
rlPghtS4eYXqKhSzMZLpzz5ahZUcvOw7rhi9mS10FYiHhLVNBR3bxuHcSCtWrO+N
H6JAlFPTvRlOFJhiDSZNFR4C1lQabc/LZNIhM5VcVPgKm2NvtsLE4t4GPlWWXW7i
jsGt/Hr4JIVmTPH276gA/xT+Nt3/g9W+iEKMRufaPNMDOwhi9DMHWw0oSji7BfTF
BQFKT8MzIIBAL+OC5CqJdAuKYJydNd4/ialOezKT0su6mx5otTUFYjPadgTeJVeJ
BBEjI3eSjZV1P7tOoYFtLnm0tKMa+m6VIBQUgGKHskCxykdRcybMMngpezlC/cTi
Sd+gXlMBZJbf8AZ+2tth/ZvcLSTU+L/NSzNGpXogZT3L8wSKNUhcHeIQMnKDx1LX
nzXQ11bCEIXUhMFhODbtV2d72/3e/viIRKN68j46PwwhByFm6SntOJJKlSKB8bOD
PQJafzWmCt7wmCh5qRXd+b81vgNhm9UaQ6GBCM0fkCRzKHWWyKTl/xIoBrzD2eTj
oeeOy3pUVoQuWUgbH7TfUpWDgjTCs8dfHE19+Xr0JCEzqqHKBxlk/Lf06d03MLBs
ELnjkyamg+XtQV+W4Ne7criyqFqaPHT1AzQnIe09Lz/tX/47DImz04muAutF4x/7
2sDdFSJwnehlcIFMxN+Sgl4/+07UXfhoPzmdJGHwwICNokg5qnSulA8IchT1IWMb
0M+U3Kgy5XZxEKW/4MO268olKyJo1Mqt4qKxLF0AYlNzjY+l1YsxmwzYzlT3pCu2
XbqOUcL088iG7wWZUK149aG0y8VM8JQ6/veu7k/OkeRDdc9NHIc05QwwFwDcpFXP
DsqqOKg5nyDciEo+VufDZ2hPDjKLGH28/3PnqLwQqy3j02bH7c5Mv2H//hreuLhB
kvu5mw8b/B2+u28SIELmKq27CX+djDuJhcM2LUtsA9BvrNfIFrH1+uwlH0QNbYRd
L4PoXG6t5Hqdh642+cxvL+U1KdloQ2IuDUmksCPklSnM1jwrPkDTl9Vheh44oBSG
CJfuxzueNugVbyM30haIaqycRY1cNEEwzYinyqKXhxeapZknHLBG6oBkeL3m7/O5
rUV4xe7kcNwBoIqpWmc0hErxMo5SY4L8vJnNUQbMni3vwDG3UO+1c/O3xXVBSPX2
faWPohl2SBHk6bV+u2VO8Dzxb0oR4L63hOIUUOhNvsRL+QjLsH0HVijcx8jqh4ZD
lqXuCX00NGXCUa4PSyVtui2OiFq9gOmERty4pXVYjfpA5Hqb8SBuYLFKjHKgi0FJ
byZatDQqU+QBLmOwA71mRRBUaU/jr+0S7aPKU40mFKuQgo/iJVl7rCWQQR/L9ImZ
8YIsjdoZzva4ur+4IHHRmnroSjnZ49Cl1pjuxzG2Or8gi5RfJCiv3GMUwr+xRJm/
87VQUUmu1sS+bJ1o/foFHE+lRSw3Aj1vjYFYWQSdnunuzUetn5AQuCW4eNKb4yGM
vmoGgf/H/Xh/kvF2YyL/fKpPNDaomtYs3xqd0RQzptIVJFPkZtkh/d6y8Rym78Xj
RgCe8bj7Y3iuJqsds4ZZXntFdI0iX4id4nTIqJSaaPwJxlJ4UEfTWzYelBRDWPTR
9G8JeWD2ezSfBHG7NL4idEV+AoUaYWgyhDYmgytg6Q6BSmjuXesJtUSfuIMTZO5v
tFH/82sOX3679xuwbrlMpKjxsK9VNwFYS3J9mIYi2zhjn8fqo3TCqXlNBxXxoGpr
GWipTaQu5t/P7FrNUsvj/EwLuSB/Jj/Ir75xiXBgFEHLqQMoYxHiUqu/QnkUmduX
xv0Aq7i8UDZksIBU8OSgsUOxrmL9m0Nob8hHHM9Fz6xCrhS+d9cXs6jUNg5utqF1
7nU2bPD/dzDJ9dLUIiYVA/pVT/VAkmkwz4ieK/Nb9+OiecSOI61DqyFBP4cvajre
JzS7VRx7Ns11/zYWd9krL7sqf/qkKLicyOfdFGoHExsbJfKcTFPIu/7xlM3qeCrO
47yuvYy/Mf7D+v1axUIaXBTP2q8d/HlZV7kKrk0VLsNJV2LVmsNxkCeeIcfZ0I7C
JsaPdWL2nXaiNzJkHAN0ywYPAe4Uj6Tgo9lYAFBCUCfG/29PrtnApJJ0ZzRycHjC
BjTMPkS3WX7wHvh1NwpAK8yXv+XOf9G4v27q9UB6gak5JtYobVRHhyzkZasJ74+P
bSRwCmQitoGBPUX+lWOh6LVUZ/dayJnsX7PdUG/+B50b2mnj5Pn7wckn1+ZIjEex
GZTbaNcwUsaVxVH6mdaUDwNtwqdOCaRmn8adOVT1GVZi13IZXmkhpd673jEZgAnF
OuyjMWwAZYOMtWQchwX+PLDRQxqTm96F8rNru2pbTbG0IvqbD9y4ONwRePVgAKGR
nagKTMrqaNMfdxzCY7hQXsGIS+0jXoKEY7iAGNUAGwmgeH/a20izzqYMrgCR/tu4
fC+8I8we3CWIPbQH+gSZqzv/vyd/uWTfUTm5CE159w1rw8ChJYwYyJn1KyB81/ZS
f/zsBLXru4ZD9nT+xknzXbI0jKMFlr1MfmblxKM7Y9MwvCvVG4JAyGKVCtfs4jFs
3cv1a9Q/IogGpTrh5jZYhkegmFJRq+j7ERrZwLxyAJLjshyGFlQmQeXuQsvtdn0o
8/zNxq2sDIR0AqlyJQWWfR8VHYVTl8WWQhozbUSOkihr+0nxFzBR5qcM1iqN3RLY
Kko5b8X5NeRESscfWG9sES/zoJW2Y7XAGWNsgflKkxeRqjv+6cWi4LpUTfVOOwgi
yPRuwC0kOx3lRJzTzFWhInU2M+FLqbqgqLMcPOshmaoZERFKWncZBJHn5POhOKER
sF04NNo3/RwQcxLO3yEuZRYSIqvhRDmD7P35HSa/gz59nu5+B/x7jhsJgeqJSsAj
wFgpty9cdE4gSUCapI2Vx/PVEXT/JXJS6rN4k4x9S1XT9N5emQjL7FwrgSgFLgOG
MHhQDgC1XSaYvv9UnCmRbM806gGRyXxk3vTsqIbbgaNkUl++Alqk74gC79UtZMPr
5w+UUPVzCbBYRnAsHR1P9leZItmEgdGd5kOtisDNo4yIMsG+NV/InHpr2+1jlmkc
Bjor6dmdne8ZFx13UAFlYonmYKAB3vgq5XN3nnrsBsSHiBfziuN7N9uSG5qcEsiI
bVt6glPV01XCuiEQaQkgizT9rvJ1I/mm0AsUnuuvoPL7VOND7gaWwPkabnF24MPw
mi8S3Jsi9g2Rn2yD7wwSXRnrESWDsxEGGpqmJt8yYZeLhqYSvNwhK3Xd+SbTIAtS
EVg0gmKoyrIX5589zkFrlTWtkcZAcDcRfOFZR9aAT99cypx+y+TZsNmKEqp+0Dns
w1LSzQR46NcloDdIibxPhfWKDxqre7cduEq2ymMFtktAkn2WA9WyKtF8oSuZ+742
GNHbOzg6bm66YUIEy0/GCpmPeCK3nDSfxXRZY2QHskemfZyYuuzrn8eiWfTf8qxL
dgPakU5RROlrhlVhoYCGDFhYMdbcen8ylR/zJsZjlMx3Gk5WXoSDXSz5DVXJEWUh
4+5c5mhyneXlzYW4k5fqn3i7r7lB1kJmK9frDEkeU2Uv1/gKjQk5iafzHpCJsgtp
hKdis7ZYNY7cXyi0ZikB93/7F/I3MYe+Pm0PZ99zIVM31AOAFXzvnS/P8nLug9ZL
9P5WCdrtPx5VE7Id6ZLbaizLlnHmxjXza1+vvxr95b+1c9re98wAg1EfE71w2qwi
zYOFb5xWkmDtCvloYOSskkdyZb6HSbQdhFrxGZPqpryllT/FLATWA9zZCxXW/6v+
wbrLmw59S28P37u6KXFapKMz0G/J5L8TjSoEMsv7RPmUbVh018hthyrNgiJ8av67
EW0ZcE2jnD50t4AgQn9hKJTAzIkSwM4ZJKarqsNK01usDtzQ6Vgs6CLiLRDcQRpx
1z3Z6E6qb6u72U+wHIZq9IwgtTUntneIXn2hS9Nzl0MnlOA8zjyHQoG5AG+rCTLc
Hq32FUs1OE9aIIn61b+r6Ocic8AVIajD9b2SFYnN0qqmVZCDtBCxfvwKktsYeBwy
l6STedO1nYi9/XfWeFMEqI25uwCgiLASPvkPg1nLqv8edXDhpjDjw0xfJe+9Wq+0
JHjx3DaQZCnRxRy9uVXI+AdaF14NBJQuNc2c7CFnP9r9AToey82cyJapoI3vgawC
lZKMuKd2O2xpc6YM7TcjkDniHqskePk3HXkuzaZpPTRfhDjjdFFVSUlG+rt5rXTk
Rb5xBQCerdPPUUFy/fscdZUeb0kOsTEI86t5oYJ1EQMPp7PL+zkg2H7/PGSeV5GC
Guab1VJOmXndJSaghqSnMIXZRWUmT+/9unqQPwz3IX7TtXQei0ohIWe3HU5HwA5i
6zaDfIglQtf8OKQFQh3OIm4Q5YZGMZ+tf1uqLC7GcJcsNmnwXOiRVKpO5fBi0Hfp
pbOUQWM8tVwQdZtqg5PvNy8NW42YYQeJdT6ufQgiAxVYgIOh/TAHEO5hSlC+aM3q
1pB6FfpyJcfcOxVZb9FLAmmLm56tMkjD5begT/V/bDiFXdH0PxylykaaY1DGskeN
+d28wmporfjqwfsHbm7n/YBOrQM6+iugh+DtIUatn/5285dkTeZnLxX75+3y04M3
ZAPrjdTMkCOH9V8CZkeYd6jVTqhui1hq3UhFhGK9poOElkkBDE2lj+gINcYXmXDP
BiSMfilsYn6yNnCznn8ju8lHw4kRSAkB70fcrPFWhtu0O77DlrqHV7dM/RvO1shP
4AnQIibRfMbi6TATZXsZhEkHKVzWHTlU8lzbvuw57D5NYt7CriGeLEHl2urLXWAM
n7fMeck6jT61PAgwTgoCOXcXYGKOATfWaLdRwrNHAFeNeZaOyCp48zRfgY+nkjfd
oarTA8ppYURrEc2tZXLQ4BtKuHPJ9jySQpqEb3ATQuZxCk1zzDNoAaDO77DmCnZZ
0jg1hUg1lElOouolW/e8yg1Z6hyZudLKyUqsI0RCtYxx56pZZPnsKnRvQ3BF6gOp
I2eO8LVbY8hqG9L/JKgZ45P87PmdIIZyemHma4dIx0av3q8wxQ4MPDqbsYmqS/ff
4HyjCNOm491u+F+fmegWNplKQVlnTYjQsaR5rvcWAs42p28iMwlcULrD8VV99Jk9
zGBhQUPB7xzzWEz6q35/sW8Ym/MQQD7HWOF7q9RrrkfDNtzId6YWADUJ2t47TRu7
nI4gPL4RgPF2sHf95TL8OFipTZYKU/YcsQAEwvmmmjMe+bCnDF/fmR+xYQfyvJBe
aorJLCZzDA1YjXVKfkjyoMr8p0qF3u3QTIZOmdHkpFNGTPHeXzdQ6splhvRHpRre
GeTxBy9kWh/29r5HwNpx0sAIgRSCGA08D9esaMJiimmdaTzc7xmMhgUxsWPO9fT3
1IGHvfmc73fPQbrWr23eURMslNyPNjU/Xl3MVESQQr9yjFlz8Q48DEpqrxb6omMl
0v/fSD/enF7wrSmQkorJNXbhdD4Bowc2ef6KEHACC0zwyErft1IDJlpqtY4q/E6L
/ssqEkG6MQcsYnLjXAyqBBZdUITeNP7S0XbIHHrd3WZZs5GpFMqpkPW+EjC+yvDv
BPKUhOP2M3t0M6GQwWLsYPOTnWHnCC1mIIi4cM+WELyARlMMEkN39y2zHBPdGe0Z
NCbJGrXw2pkcUaQinZQpynOS3cpwAgkt+pgQLNlU5KUiOSxnVD7H2uyxioNh9ka/
hSEOpVLSaddpaFM2F0hH9guwLfyb/MHLomT8nAtOzSsvTXaooGHWAKPgOpTk2MAy
b6Kv3t5MiepZDGOwbKPH7WwXIyPxxOyqXXl3kqJe1DZ6JdXb9OqcCChXKNF4uyr0
D0gR80GZVQv71HQEcS7zHpORz3r2nDY5zN6YQDsmURaGckq7TeTJZcTG3UG+f3J6
uMF2AmjWKAGy2Xhve1kLcpmtdKuG21aqLcUTmdpuzAie9eld05jhmfDftc34iN5a
Ydu39nXyOBoo/gwor1ClrcahraP7l4IaYscmLC3Hfm9M5tdB9NqTdX2enstiK+r/
Zxf5N5G3kazKN5hRUC8Kc0sMLcW58xmLmPa9Dfw9mD1OCM1iEnHd7zql4M2qGVdX
C7axsRwaZRB6BeFjxXqliHL6Tu6tMJsUFauUqGCYtwiDlPfaNdo4Cm5NtEBGmHb1
IVHSroEoQWtHBSTEHD7oqLeel0MUspOxZr5b9f9U8qYlMJ3WMj1RuZ2eOvmbbu9j
maRv41kcYyDytoyZJXN/NYRzA3pSGHSbLZgTtx7k5U/BRGSgey10PpElxmwG1Pup
cyycaLL6e33UJHshxKjO9G4ilgo0UvZyFsKUS3ZVD+Apxm6uRxwKmaC5krSmJSZW
3ErHoEphD9JvM6NWe0sYFkab+leoaga1kZXEJX0+xjUgPQ67Rp4w6OA8hsfj+G7d
1tJRm/91CBlDKAxLJMRKVBA9lJlEHqDG8WRkcciD3MDNQMEFnmVBy6a7Xd/jqB9Y
F1+6AAwvQOJSLN0FPduXYkYc4uWyNZO+sD2FSKbJXXn8VrvzkMLy3ERB9/ufkt+u
pPjFWA1/aqmHof2ijM1VcTBFZ+vCmqoEMN8C1Xh43ozin9mpLJZc2O77j7ZCcu7H
31Ib9DxYNN32csS/LW8TtnBWCZwVR0pyXkHtECpBxfNi855qfTH0dNzVtK7+2eQQ
9nCmHOU0qBtpBcfrgObbQBK40OtIOP+iKmUOHcDKOpceSeJ09fEWxXWqOjhTXGb9
Brfy23ikD16Fhxmwqa0wGLw4SjbNvScdA2yH1QbKIPOjzQzZc8sb/TsADRILB2V1
fZnWavt1v4n/RwfaJ/4pZE8e/cw90qRs7uFNOi9jnX4AT/KvV+1v38akMumvlJ3Q
/08cUsV0vlrzSCg8Fo/Ce6U5/ucCZuyOqsiFxV1Ji6GyA+doajASHn0qp6O0GfGe
XWtil/sqiIQ6SqBYQtp+yEK6bixiGjdkiUFXjYV61seTz1GRFl3GlnhDRd2GcYRN
NkPuNvcPnIqQfUJnosENzo/3s7/+gA4haFcZ4mkMQdTclQ3Mk3MJolttmvQro0ic
oyuU4o6n4zkwn0r93hLbaaooYruqn7G4Sr0BDChs2qc38VdUQQBtMU1q+2iIC8GU
XYTAlhnErQErJkgZBvJ6Oa7Z6DLD5BJmPvzNx7TwKwZLnZuHqqdIsMm4dMoBM29u
h3ugnTMl5VRsI4pr/MgW9ABCy5UKTXRB8m/IruJOlyDN/udF7G7k5QPEPfzsgcTL
sXLNDNjTewzYFdtxSvOtGZMBNhc1bsaS9gH17pfasm7JiErgEV3xjB2nwyDNSxAw
Hhk6A9hi9tKCH6ndvuWXUxgHjSzC0/Iv4asKrTw8tERQoTEpHypbIVX59w4g7Iv4
YGYyNPDTPWSEazXRR3RNZV+8QHLXkyDEcl8JZp6/YcMWvvFjtfJRpkjdcycvL66e
fLKiSBZ921qZodqUhAV+em8VtSxldyHU6kmyuPmgyJBifVXMN0TGSmjWYXKWsQZu
3Ph24dvh8g6xC8LwWkb8g7B7h7i6dzW/QijaOP3WPQWtoZA7DJQlqZ0fnNCcKI+J
bsHh9M0Dhhdsjj7+0WXa3sfyNZ9rCqrhM2Sz5GNFLIY=
`pragma protect end_protected
