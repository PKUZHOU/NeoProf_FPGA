// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
e6mlivdmVVLQv5J+qtNmqm4+e2I/KcU2ocl23JNNYbwuHldmeyukbkVizWeKfZDk
vaumj1EViaftpEpCPp3mJk70/4aYsje1DByCclyRrQ+hy5jQZX5f8GlG6Z3rJ+z0
9QTTyJwvNQZBrQjvouW5Xu5TZGgjJTnrGy4IM1aJMl6BLd0dWqxQAg==
//pragma protect end_key_block
//pragma protect digest_block
eB7CvRitsrBaRBd9eRWCFm7DAWE=
//pragma protect end_digest_block
//pragma protect data_block
bRjw6wZtqi8O340Mdhv7Y/suchVcumeOP87Xz0HcBiELBZ2ExypPKPm8Jn2G7Pw0
8PndIXiwppK0VRd8M5z3c1zL6ZmnnTnK46zMJnspT+ODMHIzASyrHtF5x3sqaZL8
RrhHzTkbg9n1xo3qggur9FDxM4L30xWukL5o9opvtCUtxU5suIBj8uHgYdrFR3K8
TUhOtXNeCCIk/DeQzFecSao1msD24igzYj8MewnG+5oSRonMYYN5SdxYeZ8smgfF
fHqKgw7+1xKXVgAnPHJF2MuRxGhqH1BKjGc+Kcf6gb1lj2G9EGzXDfMZYGWyRuUt
QmjUnqHUq4596GFp8C9yMmV0EgRv45qeCcbCUmCvS4Iyj0Y6fEYdxgErvs5jPTwJ
koxoLNB1pus8i2AM7K185ntzHPuDqZnTyTJPb/A6Ik8caEJksurvrTw29XW9xoG8
kp/1pda6VTZpEq5j+mF/CQ5yqayz5sh7n2KuXtSjd/FGfPiv2BMWdXJVusaKrKRs
AOb8hXWiBxQKP6o1TNIhfuflnAaAqsWxQuzcQdCMnsDvJcbrxq7m7p37Tz3owu5Q
KJs0YbTdMuWxQfSOJ52FcjyPWuGkJh9h/58GgvZn4SKaQJw1cz7a65cuckk/l0Xp
eO0UPDglQeopBZ4iE+wxC6rd5jeo/DkC/3OrSHnLAXsWev4QkY9CPFSJCes9VD0Y
9x2RHpVtqzvfUGZ63zMhl8GTbzHbBOVWPUZkt80hT2FhuKHU0HMIY1R2umGGuPIf
VpZxeiHIvvXmzwWW5BhtI+JBkwI/6lU0PtTVB2x2e/Z5LEIx8rT6ez/4zXDi5YP0
uouqQ5IM6pqh8hiWguzmvOu+2ftFfNPSGqduTe5CgxMYAgz9Y3rHK6v8mDMXRN7P
0jTheA1qPqNR8haLvUrEgGi8atvo0Dd8RxXt1TIw/kbllvsdJlvEcCQKN4SlTg/9
XLauK9/hHS9dBWMNsB8RQTeN29sBIX/qbmPjl0k+FhRJfCSj7Bu65exPqSOzYXzK
Sq3bmNNhSKwY7lL9Olb5G6izjMmwRAV8+fdiLPcx7gPoFNFoQSHTi2ASa/19hH09
jPZ8imK8EOJFOrRzdnRNaIs1CFT4XFoQhmD6ZGIWdnexL7CrgbASkGcle3rVzjin
d5aFecpkggsNj8ycs5fHvohNLmMU3sJBhkYHrCuA1O7vSahZRSmEPzyQFh82hvp9
Jbit6x63CDWjn6QfetRkvSHPsv+irucie1EspGwAy4Zv6krQMjmXpBC4bAinLEx5
d3fxsex2vmS7qN9+ySNGyw45HSiS52rKC2s7bVmHYUiI6cs3d9cO8nGwxa6WzxGv
6mdinJ6alaT2rdzeG6jrbcjMwV6uujwfcsG2fL6EuvAqq0/QhsdhwZceqv02p+dx
zxl1fbDUbPBwK9VNQowbrUrQ6au6Nm2tqVMHsZ7bW/uOeh8i+hOxP3FrrQEf+Ghy
jrDY7Uo0goficyEOQCPR4A7k9CFIQ7rgDNp42LMCjm+9vHOG4MwuevVDHVrGKXnv
K/EWRATvAmOxPbjEUCKNYkrvf4l9zTaAVU5cCZbyf69FNVFAplUlDa6hAPF8Y02T
u549KdXayjJUXtcCHn7srz5vxQCHq9349EKQtpmh6W1XHO1z4Vz8BYDU7RDT/e0y
Z16oBzfAobUNbZASXIhGhDI1BEmIp8juKt47WMDCSA3AfCGSpnicMZA7GPIMQNNv
nM6Mvd1IFHSibuqm+bhAhRrS5Y+L2VVDQeL5oQQHPcWo6i4AwUuTqfPTvy7gPPP5
pu9oI919HM45jIMnLEEjbVeFLRRJkDwn/6koUXBozt6WlegeLboElhF/BYwfYyxl
ZyEmAz0JInKal51kRN5Hv4W+zZkRSGUldSm3O6//NZOli6zItJ6KWoOYwDPL7uHi
iFiSMQKFeca7Tom6guADJ92BdHbOVCD9o1PnkZaWbibsZ0wjJdqtAA+YTL6bxZT2
lUX74bNWYrNSANjfydvLUQRFWZg893SolCVi2VTYNIdoqr7ASHssZM1XusZpDVIF
X4QlFasXXcjAubE69Yx9NyvrsKaXhHk9WcGztNq6oRdRJYxvFmz0rSbU2mK1WAnl
dXCr61ZK1h8dRXvUfsrwSv7tEZcxs0ItKdcNjapEkraSpg7jjl/jZL9C71KwUwvV
OBBCn8TZcDvIbHjSujdZyrazQrK7OYDY91zVjSfs2F07/WHcXXUW//nd3ebPXwsE
qbR0GtZ5QMvmu0yuql9/SrUhnS6851G5z/ca/VkyChfbSl5qrwoMjp/3Y7rioJqy
yqwaVw7AMtyIhQ19NgnvUsfNFEWNwpNW/D5YWJQkdv/z1kgudip3Wk2HswqnkRHk
fiZGkdMhudX2fXmcOgz/B3akmY3uqZgtvfHYafXR6UUznbY+L8+m3DpCbiXD9dB3
LRFzEboTKccaUO8G5mpgT04XT1MqCLaPqQZNcNpozEK/11hufojmOfmlkAZMeQrt
nZ9atxNH8CP6NX+gfKq7ZudLtUrNLXdnukO2OR0FNOVh4z+X1UlE02hcMsz3DonQ
NUNNKA61HInZsEWquyH9D3VyvS1C5FGiDn1CKml9WFQKlhWYHwpWK8A7JK80ZY3l
COQhSJXnzOGuEya5NDAa1w0B2Rv79k74xcR9QA8x4M/ePw2vwMvhF876uJ80lkUI
4mN7OOPff0ceBLMIuBr2tt1VxcahnVriRVIG67oTupiPAibKPYACZrrqb4FWykah
OKG8vzdjYleHDCeigaELBG/mb+kNsjqzr71AsdGDV29iOA8nQ10Ag/0JllatQ6Us
8l1yKA2dKbAsgEOO6N0j7o3gNRmviM5vQ65yaswRxfJX+omSuDwIjE8+PonWGbD7
QEerK5UalMPUjwBz3MCBTgopLUWhQYLz8A38EN+s8idPrNAKXJrean/7sgvAjauo
0mFVD3zchJoS8ApRMnnbBTl6KOFt2o2WY28MObWciegdvzjn1TCTEUiQn1yuvYhE
hNhw7VAxCNFYvvwyg9KFFx0zaMn5EAfhHgZd2Mvo3bU4jZ7J0vL+Kskk7QiFO1E7
WJAiQv0Gx09yTotkhQXuuIEGh+aocCaXFaCm9rXHOv5wO6k40kvvmaGnjYf0p9e1
seuoxjpI5JtzfHYt7fXekHdPbSuNAUEtKMKNWGAx68YR/wheiqPeAK4KqzGeZN9u
TgBJO5QvKj/30MVBXhilwW9aAcXCbNVNGd1pFP5rmMkdJhbZGjI1s3A8ShigHkJf
+U4jTDuHUDGLARMqpS3oTtg7lWnFlDhoRnC8giy4q3nJ8pHDoTlw8wFmGz4DnzS9
GFaX2m/l9geyctofkHv5Cwt2RLBsyDBUrJuiD8OEhMoXETjZoRtz9QpYzgGjbizD
IOlt12Ic14M3vuFd72ZMV7fF0b5fIAkY3Fux6tCOiHwvqpvnExtwd1B5JrMpY43M
8IEfl8dS57PlRjIFSyksf32+wAGpbMOm5BDyPSngsJl3QPoXqSuFQIjK8Rq8YW9Z
kTsMX+j2DzTrUXxESNJGQQljwM6Y9lu2xsKEMphfIMFsXsH1FDon4Tgw3UrRDVV2
05ePUbevaKIF7ZGfSt7euquLK5uGKTY58vIJl5BsaoKwBN1hABiSOn3TUU+Jo3eN
u3ZXKthTGXaSjshPsWorT/3NroCKtAH8qkVslKroiWI+EK6nNJSs9oPXKC3flZkS
Bn5xxHMa9YMKHMFmHc3i5zayhdyfylhwzxSK28KlO9gkU1b4D5xYyPWy4hLS5xSZ
e8f2rF+bm2JkHlYKDgXcPKSrsU+mrAJGhgPLs0NWyADSltha+BEiGB72CCx8y1h4
U/A5FOmV/EcYc0dfxSrKbW7DxKG2xzjTh2cI00B7VpME7Ij0tSYfuXihR1c5AsBB
ei1nEW3sgUMmQFYZCCDN+FIPpcteOkXykekh17iny6R1k3tuU6uBwCDhQzWuS8VK
eic6d+x0KmtUDd4mjMuPAA7gBid2Jh/V8JaPQ1KbPl8jkR1GLES/l5pmYm4bMnB3
Xma5XK0OxMA9WaVatcJGgU5mFjU+/UpBAH3RzIniT7QfiTQCXzeKlcnqi8szlE4F
OH8olnLXzkLWSiU4ei2OM9TwqTzXGoyGS2NqsLi8bgV1o7O9NR0hATQ8KVDusLWb
LV80fP9Tr+5Hbc2rwOY5iF4ugjKyBrNKqyj/OXkI//ru32vYgwPxtXx2hbGamAja
DKgTAMNicJE6hQC97eYaewWf2gycm2iXkqJbXrUcc/o+afLHXNHhQDS0JN0X9Kw0
Rm++TWi7y+LaM+eUuFIrEQypq5BTXvC6aBRN/IqFtj3cxaKvtQer1PL6Nbn9i7Tu
ETDEUfFOjhTge78tw3gVM3MjmwfsatrccHLS0osy5XNEvX2jCw3EMUcmUIzn8k8z
lNT5EZYJhyVlLRB2jiIYJm2MntlCrjAgR2LDls3Ir0C+O10NyzF21TYtuptNeMud
vui1oD7H9UbPx5PVxiQMqgT5dTl2tjk04sFRvX2rZfM6b8GwTYbiRp+0B9Euxccw
0AvDf6xcULoPlyTpfnkIhAH50hUwfHpHhLskIJuVsoosa7/RGbetsky8Lnu7t629
DinNOxdqQa0XxD/JFyFZubqZqa3aQ3E1n0l+uT/YmjvGnkGOIvZH659L2y6rEdkp
/IaBnLIC/Nu8O6k1LusimNs8kx+OmgTX8DXh3gDdM7DHIgXfNhNv9be90t3njxRb
dreeY2BzWTlMH4rpc+aoeHhXh6O2Byx2uROJXOjFt1u6HwHq5Q9xH1x8FMuUM+nR
DniaSV5PNtP/gU0I+5bE2Vid+dsdzeJnXL/UnCXpT0v/GVC+mXwxcoxGuVEY2Vlh
fI5i8BtfRU/9YcvRjCOlz4kDaBkAnQuJ+dfvojF2rGxLma+YWA7hY6tpq/fKlKWL
RQ+/LW0T7VISm9x3lTaBoC2roMA2GlNzFLoXHXOnrFJ9UPdF+/Q6okHUMvm8O0w0
7CVGSho6ZYB+6PVctfsDpPVhEu1pDLazpidQvZWdgVIjJB2LFF1i/pnU39SX0yKl
3Bu8HVBH7Xi7OrYg8a8lMuc5zKn74Yxp8bp0G7gkvLHpI1hlg7d5sa/iYiohovmt
CDDNNnuxWnS0TR0ggFyBj31wo7+9TIq608xpLr5tfbKyomrAYQP6HGhAu3u5uUXL
q4hUrYS6bxhxfgE/+pP3o4tAve4Q5cADVo2wQEUqadrQfldkTOxdHn4qbIplHjXZ
212OV20+lmQ6++QXcRMerbDYzu9Y9BVdtKv3venB5wzNFwZ4SnhpKDYpt6lkkxeq
PCOY4uXagkzsza/mBwIc1TfLOniXO3iHDkymCZMptjpASWN+jPCcTj/SREyDnOGn
O1Em45gcr+veDqcX9uJ7Q7P87AObwKszFXWQ4R5cT1pjR0V5jAFu4i/i7WkhMUtT
dpLJslZB4x9LuP6QCOzVzqjz0Z7Y9yxyVe8pLxJ6F8qXbnOO9WkYtt+8VNjhp2tv
xhVyjVVHoDqrT67xJ34Y3qqJr4t44RFdAML7tvDzmcg+jdFCGXKJfUN6xVHC8oNb
89OVo43RvsoW435CNesBz6vTudPafeWbf605v6T+MJm8XrijqkIgC+Ea7VbRqnRt
01p5NO8yDNdUZkPyPHbZP7bIMa1fVe/BvkF3TWZujE2KJEbt+lCFphvWjxO1wlvQ
7VvR6lSFjm2mTNconS9NDBruZk+G3/qL0ZS/89cwqG7ePEV3IBIZvQarK3XDYPpp
NTr047H/7AYQzAxvQsHwwCRlQUihEJAgE+mnoWbGvC4+S5AxSpt4MvaNbspKdeZC
hsfy2XfPWeD5MaePxIU3wsp2TRMtCjF6uT2VZ83aQXkdw4gyv5BFQVoIE+lqv0qe
kPsfCwpnrRWKhj/3EPXYipOz5A/31eGcZfUwC64fCUU8GuMwGPnQnPTyr3RyK7+x
tf/XrT0SWv7P4a+mNJfry4jYp02Zbhw5Q0et9nmPyDuVimnsigBQm+F8B9Macdi/
Zri3UhnImN8j26FvfmsWK1Pp5r9xeo2adIwPOYkt05gpyWHgfXMNrR+hSZvhI93/
TFYgqriccKtXxJBqPw2wa7tFgArIl3e7Twb8MSDTf0hI9UkJxJb14Gn8hlXwbgzK
XnGtFX4Kq8wTSraXvm5VC9n6z/g6toe6xz3ZknjAWkod+9GYSMhSuWgjd4O2GJy1
nJPArMswO1HYuKxWxTCv8GJK01BkyE0sQooIsZj886uX8Ymwe7kpzhJm0+FAOIpJ
yzKulexxhRKi1pW1ww1gLw0zpotMLYYd/ScwoynkTE3dsOrl9RUnmJFLL+78qkFc
LAYRxaaH3/butsApCa+f54aY8oUHKhtsFmzTRnE6CdOuCvRBV7qolgE9uy3fNGSU
k7G1LMN/07HgUhE+z79/9ZaujEGXfO/aQibNQUYRLh4vD3Plecnuf1ZB6B86nft6
XIeBWmdopFZjJQu1RBflTLWk68OIlwFL5Kd2ns8qODyCDiOScu+mQzaPIxF7HuCE
4pXiZrhFse6aqkgGo+qNJrE61J0EcR8vmzip/lyFu00nUzjQ14B7GYmGybNj/ykW
RiyrDYNR8BvbZHTyt9gNd3cWW4AkI5HyoNbBWxTnfELYHJF+SsAiIwUnC89g1eFZ
1dnfDSAPnn+PeYsWuiLCQQTzGOIc3OG0Sh3VLsL2yJ1kuIMgpwyNdvmrgE/8H+GF
8QiC264Gc6bA0k226dnaoscbeLNMR8xj8A/zmKYiINTq29Jg6D5flRvh7N1A8sWk
eXbH/KTeTHCFwPagwvaj/KweriGuZ/3F4UK1354abZyQ20P5yjK5o7S5eFh6lQ4j
La6mCc0KKGdcS++LjXWt2X9mBZl64BCggIK1GCPhUKB+8HU+gcnJTH6imDDwQy46
lx513NHvyhr6lmWJ/OxMuJQql4lNpYfuvt+46buM5uOUmO0tFs9Qgk1hRpHnd3JX
L2WBR4AO7aARaV4xPicOJVkJObJOXYCr8cuYBD/UsfqNtByeSZrTWD9EwGbnMTzi
/7UkfwBGm3utmXbAn740XoyRt9WpP4IwDHvzsyYwHlMiLzEBm8GXH4nvWxId5rIw
DoW06CkFq5SaeYSo1OVWI8RMiTNoc6BMuywbQiY4HghedLTXh6cViW91uGq+jgSX
zKtEmRUbTpuUu9TCMrz0swwq2lgPOXrXkgAqbS8vd8vftbOJ9J9UdY7+G4CnVcK0
UiOfiK5mupk28x08ipetJD+vv68s1aD12iDPlWMr2VZnlE8VCPqDrDiMp+XTUEJG
kSi8I9/JMSXWURIuHWSJoN9YpUaIRNBJh8yhzIznZuI/MKIrAubrK1BR/C0YBTji
RSWmZgkLQmdzDWg5oRbDbEf/vy0WNYZmwwmI9dktK96it66sSbLROHEQCw/MwU1l
utMpCTFNLO3WTPt744NpfQ3ZdX/np+2iMp7eU9yqnq4He0REWnkw0R6Qiz3OvC5z
w4IZ7uQfn5wFsCGivXnN/iVlW3clltzRAi2/Xc8mwb0gxYLyq+O8ZgwYsYcqEoqR
s+hT8A2R1+NZs3XWGBC1N57jEJ9Pzy3yG+neg8wHiWy/2bF8yTZglljaWJDZ39Ir
nMa9X+gVCsJ6yr2oHZB7wCSWcEO1xdpX9KuoVCk8SSW4uYrk3YN9+jHllxaAAZ+q
Y42lH8p+TdWCVA04D5j16eT7AR9S63IlxrnLoT+E8jZUqS/ua70OQKP5V4+wzai9
JMo+y0xrdlTdxK4nApmf3URKKrJU0pymRSnrrzqZMvoMmrWrFB2Xp39dJIZbrlBh
S47k2KBp9luineZUgkHhwETVntsRRfYKFF8CaOwXcvh9Yg9FDAVp1ySLdRpHSJI1
EQrWjaJoXKzhsoCieojceZLXj1gooFcVzeQArNNDQBunOAkpTK4fHqgxfkzp3PDA
ybIxhSU9hfoeDYkxS+aBTdJAYA3QVTNeLJMXJ/mgtyXBQicAKsLNfSYvLahj7g0a
uycxQXpjwo60b/hTZ1BLH+YCtQ81nuPkzPPS14nZ8ozg4Czwar+Zgtfy0ZfhnxqI
Z9oZ4TGdWhPDtXDwuj3DqGNLpMJ5loCJl0Acqe2BkvWiGyxR/qdQSm90bPvWIApT
NvL/zbp+ckrSQA7KI+oMcKo5loYagsxL5FI2N+y0qUFsA/0lpta1RhjHzlPr3xBA
bm1AD/E+MEqzWMG/8eVwtsNE03gP7K5acMXSS9OBUof7o0BWNCrKXvWvSrWNfvw2
jrgbC/SxN1JpDSDX3+8vWevE+f+GvoPmhXbMqgV9tF6A4ZL9BDjM571BtJE/FA1B
SdYq2ISLQELiQXHUOqHULESQhFxCjEHAySoVno+RO/heIJ7BfHZBTUhdlFECAAYd
QzWz7CHvsBtdL+4nMJAbO8M55Af9eFgtMOYjpUxc+W7HE1Wm+W3KrMCAgTclSBcw
2apv2xNX2EnmU5IHpKV/4iuNncK+VVRUuJu39J81wQ5mh19XanB/PWvOpQYlxe+u
2aW/l8Xpy8mvX6a4nwmx4ZqRIsIA6Wt8tff2WW82KFCeM/8EDr+1i/W26z2GgcUu
YwOGUBEbGzsnCEH/D5gDCOSSBv1x+lZ14hH2exRAIu3HIAiZo2LemvUlDp8mnEHP
pbbgOo5/uyYQoJb7O9d5Hms0/CkXJ8qMofd9MXdsPrtkcdUHBEuosNtG5L0q/yae
bIoM2YWL/WSSMQ2t85+LYk/G2qM01G188QsGBmAB67EYxqiNL3S2/6sQpuBqDskw
ArDMXwEz+PUSGhXhha4Rxea8PB1+MrQs0AMo50gj2NPxxaFR6f/7BrcFM6Eo0/Zu
ZjjPNwojSI9ocrZKJMCbq9X/l5Pi9MD27RSYFuXVtQb6X1U0lxc71fOFY2VIxv8r
zQa81WlRzF+VcjGqAYgq67e4YME2uCxs75z1/bBML5NqQh4a+zOOfFxururV++3B
aZcDFUTWcr5hVOoOa/ag2CFOtiPmKCAbEdGJcRabpyi5z6fMaVTTVq0ZDOVOFFgi
Q+CqK7F/enciOScR7wQuLNppZ9pa+v5C2PxOv8dNZw7lpd4Jmu9/6GOKFyHlPrbJ
HL3+oKQRaDbkpyzzyZp7TNqC+HlvFsPl+q297gsqb2nX9uVcJRW/qHvOZ/I1Dqin
2kYW1ryNw8ap27alj0J3I7s3xZDiWFd9cjT8XcVEoeoveLeQFm8DMhwsYyHTRB8T
FIrq31sH0yO2o0xhb4bMHb+CC2EuohWo5fRi/ZjEp+gDSL+fGiRgJfHekgPfdokG
tFLyoCsO9kX7L4PDcPwhP1y1ObLt1z1ca4GVabCCMhaxZ8ztVornci581j6s2zxb
Q/eJ0R2UcOGM4VcBMogUXTpKk5WEf+xea5FTZzFMp2AsRp7DcDAfiCUBUsC494uS
cmVxIl9acX6B82LrWJAcEGBYSdWwUzKmjmRgdUxGAQpyyFIONS0o3AQ25k4QLMuM
Ao5ZUqNQo2oFHYJexMKIbhtYLkwgNNrdELQ862TOW1mz54lmiRXQDpCCC16tvs2a
7CNGvAusHVa05cvgMHkZ61ZgkrxjvL5DcwjU7v96R7OqizGW13rTqgKUxbjk0MQr
ghxT9nqAdYnn79u+kqVlyrLgWbNRcC9UonoSC91BSru0JOwAPTXmniafQefDyji9
eLtDeid8cRXaAraPBimWMdKCkQvKhkwmQooEu3LbA9br/3cD50CleqgksLju3Ey7
ge/kOwwWx2WmWzSVxS4hwn7b+qua4dmPWnbJXAAbZxTV6ywNGHSCQoTxWsoyXyiq
r9Hk8kiBrNrbwhQdtl/q5ABdMK3EVQBtyFExDHP7uaQ2RV+MNmaUyUKLvDFJLxS3
vM8yp3zIVhOCUXuVJFIZ8PW1a+hrpfzDUksvxY0uKK97jBZF72aDbkIGUpZPE8+A
/68aBEy5esRmme9aE0z79lDzCCu9I7SXGKwiemKYzOlKse47bn/wCzihknnixUwN
WWg6d8Lfr3wt0ZEstSSBx03vnwhAUJK2PAQ3QiXvh8NK3Z3IE7shASbeO6oyLTQb
T085eLfxDQ8pnsyI+17hUl35tBspJNsr4gufIqkTU1I9fTmM04AmQ7QmfETlXgoX
oHOtCenXKE/fLTgB0E5ciC08DVEY3uImJ+ocyy/J7wQFhUmGLyw/0Y+rVSFPnwUe
MKKcI7rEpO4KqPnwqZksYJCG5NtcLlnKcc/HOrZBTc4u/M2enp8wwbNs8xASMoal
17WHWETXs8ubZoG7wT07Z9AgdopQM5W/At3qp0PnSLYnXTb/TNwKhwDTWjAmrk+9
Fd3wp/vnyj1ZBh94fKzNxIrsqmpHDTcLtFiLPepa0edq18ZScvJKb31cPfS1RL6b
s/FCVv8EHG78pThLgnJZZlKK9OzG7W758DgaFseXyle/mI/LXgeQg96OSd/IVilB
ejHSpqCXlcEWLuqsl0crI2jK3C9vG2nZZaZQik5wSfFpGTn0xz1MXwkWZaPHWssi
ov23PiECBSWL3eteaa2nsTxchM91htJzsbYrzmx3JhXBfw2zq4PPSGyH760QqK5v
jcs0p9yKqcWLc4FDQv9mWaGbyuvA/yEdn3d2tLJ5AyKNTaeuj9C9N7RGTFN3v7CA
ywkj8F8nn6yFnjL7zuhKav4IL02RzwVWjXw1JZsOUmvP9UxnPLDnVj1jp1lP2WcK
SyJ/x9/0HRdaYUrm+iC8Jkbyss+28eVO+Xa7nNjMt9nSgTxdYAxMIPvo4b1Go6eg
Rdf9O3cxOUbNUE4HdHV7Ksx5v6m7vzKdyZrTB1Rc6REJawJQTuCjucDekcxsCe8N
ndK5J8SMy9PFwRlkMUsxHQ4IWleD1+fRqMaI/8OBegg1Bdb5WYdaNZynq9v/FIHT
PWPv3+MxYCQovf284WeBgCKmq7KFHB2oyOnEjPbptYsd9Rjd5VEDPZHZcL2dE/3i
zVC8uERLEzxc7jg1PK00cqblCYrgYbmeLnAvkEk1SpIEmkgLSb9bw3GN+KOS+rbO
oubgAQdgPG101LFUH5yTfLqOXIHaPh+SybAz/lPqX6Q0cVQJ66FuiYHlMf4BVtSN
9ZBIszanZQZ4xNLsC5mX+F6cRiAu5t9TUe98+8rn2EaUcyLf+uxGVoIvTp+KSqj8
4B5fUuAvBBGYgFZqxP0EAlGaQNcLqqQqsXDaus8YABm45RoMwyWXd7279oCVw0HF
HIYaQtjmMzlY0E0IvHF7UDSnxpO5ie2qTxbsrN9rLDZz+JV3aHSaGDIGqGgcX6wf
sp0ufhDo+SM9offeC67vb0bqjjfSQTi31+SgK7noOV+VxfTkABTHMYxip8oo6x6D
eDmD0vEk/Lo0olrJzWjQbv0/+Q6hfSF6mUArhscv/cM/xipaqC5Y0ERLMGO2vsQE
UoJoaZA8y+H/u93u5qNRrPLKtOqEQ1UKPUDfIaypcvxSHF/oxHYSx4WvunkTYckN
sWqe31ZUL2pVenkazk0ifDdOYWfGdOJ7Vrsh04hXLZaIQbQrp+Ak3jYOAmIqHrMg
XerNLiZBQr/Aom5bM1JUrwLCwMNoBQXRa5zafeZvq+zPLE9zPwuo+owXpv6t3lsh
t3btyeB12cbRKlgqEDaEOt3W/JinmiT9fbWLKtYZPGbfwDGjSZw22VIwBiFggU5c

//pragma protect end_data_block
//pragma protect digest_block
X47buFHGdAvgRe6JkrxUgawaE9I=
//pragma protect end_digest_block
//pragma protect end_protected
