// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
TelzYDK6AThdMqADFqUzXfxV/6waq5DVqa92897l3TCXZAQwPqIcaJ0MZav79mbM
jbNHPxEOzUfwE9JapIjmmdG9KSUR92tpax08wcw7NML0jpHG0WvL0g1uelUmMrNi
eDZOmybH0NVGn8IIfjr9sqL79sLvOdNBAwOigAG+1IxJ6u0beYmh9g==
//pragma protect end_key_block
//pragma protect digest_block
n8C5E6Ups3UFLr3dPth3TAwmghs=
//pragma protect end_digest_block
//pragma protect data_block
MW8xbMiySYga4QNAHBomAxi/L5FjVqr/4E4emhwijV6BG1QhlQJ6a/DUSprKGIsD
q71WCqe6xRFg+7v7WnGkK4Lxgl2NFJ5SfODvmFYjRZunbd1MoVbxHfF9dn3eLFUk
xgxM+2G4GwPu9Kh6jb8c6Das9o3UEXwUP3Xq+oZU38TDk7NmRWkrpUgGRa7Na4zW
xpEOQ1jBxYxtWiqnT71MyxjXZzO3BZZO9kpv7ytwc643ZkrGyfI4kRbrVHUwm6qN
h8y2uIbOYGQ/XT9Gf5SrUa7pK8ZRq6j6//H1wi1BYCe75bKUoWBCkxt/j+USNJZ6
6123GxHUOVH5i4U1o+/AcH0g8HZZUvo54TJ6aOdM9tpWIhrhGXBCZe/J2uUpDdYc
em1eBzm/g7E7GV05H0i0g6WF8WG20CHwwap4bkXQ0opGtBr/5CxewxKOfMiW0Z9s
xVRzq5gkMpDsdCr6hSP1qO9uJrL/NMJoWXrK11Eh96dUm1zj540CPzZXfL0eZ6gB
HwSH3zMDUUDaxa088wgUubikQH+qcTDMCDGL3/V+4lMZyaq2Lk+EwBU2jnMcjKy6
40tclKj2AnJee117ypC2p79S63MLO1dbhRj341NJtrKBIlxLH80cYsgJNiO/w3u/
p2/btOZ8KxsD0+rGC5uMUf8pZNej2DKdzss356KoGL/trPeSXucM4LCbmH+ZrJef
8m6sbXnA39pPBFxfKICx5j1mI23ikMCxY/fF0eeLQgMrgjjkRJqC/SaSf9m3vWGE
Or1uqiIrcA/IVYX35C8pkEqxXKyn6h2lYQe2EoyJjwXb4m7xtMie4u0RCkko1hGe
RmMzFTWOxjmBni4kjWAEMSo2SPLbPfGQU7nRxEXY1iHT2dnmAhvH4TAl/32Xn602
ixf/y2oyq4fBxswe0mE4ujVxRqv6tzLk38R5qaiKn9zI//OX7JbklcFI8WUa7eMk
Nd3g1cIjdn8QfS5rbc32/jSMo2Zj0PI2flJPonGbedYrQjQ2tJ59z4OoCDZbHePa
jtCsHf6Dcvg0K5LOCYkRpgPwzXORs+GjS2oLrlnuhSHMksmpjg+Rme8uXgNffppy
T0Q60lgt0gVv1dO0ags3G+YhvPlCh7KcxUxgBBaMpU1ue/59aW2TNSiUPtuB4RuX
8wJU+5RDmHedTaNR2EoUC10tJYd6IfNYQtJevU5l+cnNYwJxE2l+O3L39D9cW3+8
UqARTDJ2IiMNN8ICZYvZoCUscj1XpJ3M818SSwqXGbewbF4Gid/c45+YSzuAFN3Z
C9a3YDQz4Fthxyi2aDkYsscZodLOp+nnppvwEkog2Ols2/E2q82CC4eRm4qhPMmd
Jycge3Opv6tqSMvTHk6IEwTUuWgM5TJ4urNnAo22WNdpoul8cJHEacIF5eB9Amx6
qBFekpnrSk4BgV0xRgXNMqWJyxucPyFdWFxZVHlKDUv0PEiWykB+F0cXgwsEC0rp
5Vgw+dQ/qAnNqDyYoJ/w8M5Eih3nxvl+oBCz/FmGJ9uJh2kgPx9UrYRK9EH4w2w8
wql9CBtkY5SU2MBBokiy2BlfBcD5slCN2ru8VtNlHM5Kq0JZqu4nyYx+S8wshqtY
3v1vtGNPk8cxPr+XlwZM756/ruQLXxeLfaVYb2bgnwl4UE0iH/JUoGI8Ljf7TVk8
a0PzGT47DSw1i3WnaOdvGNCz7oYjTPPzdoj80ElN/zV+zXA0BmtZ0y4wTnz2ciCe
xdLQjz9XLqi5/PqQdIZGvK1ooAl7XLvk8oigPSRQFsmC4/0DY5zndDKjW2xl3M6E
mwfa8LDRpT3necwbTqeH1No9cfcBJynSW082bceTKlBxMfvzjaH+oCI+TpQgc5l5
4YqQY7D/SkyfuPgFhn0ph2y1x1JfmWSc8HZyPXla9K4yEiKq/p8DfKrJJc8ZKOA0
zCeQN5UdCZ49BzkjnMEjkxu3j3n/y8pWcSxeobzhyBR+HmHl56mi2AAs4X2nq1H4
qTKj8lgtODr31SfMu61F7jc1VA3Nlhj5F1GAOB5LmYhDKebmgcxhvtre34PZgCYW
9oxF9ui82zW4fdVt3+9mY7i/Zi91FUFqqN1KnBIotHUwQ156dVGyc6I5UrK+f8W7
R04hM6eAr+5KedypYXy6TaCxDrntCG3PNnU/PEQdY22WdSkH41zMIyRG7dZZTyLy
msuXwIcZBA8SKYjvg456/OPUOCQ2oB41bvmqph6qgbUyB9mSAkWEHCRno/b+STrg
EFUD+ljGK+vI0dQe1Kn/o3gmMp33S0knNghaq7yWhocCw6UorRAkKePPYO8NR2N+
Iigdl5wP4BOlBl/lgbp/DoiEPGEgjPtkCzDgE9tga0C+kcKOuF+iyjPBhMiC9kxy
z0zfsICTRZIxv8g8YlXBf1pVMkfZPCS3W7G5S8S74h3O/6Bat4sH5Lpyhhm/02ch
278u7rRHJ4SmA7VhDgnkVDzr/CVPh5ErK1jIdTQUwzggCNdsQq/SOMXMGC6Sxsku
/yTQr5aWCw+tqgisBVwwTNFnQ7WgK3zp98xeuMgH/ON1Mf0D+vmDfMiACZHlL+DN
HPAKAHRW8HQR8Okuadt4rztPe6qRFc7OX82mIENjwg9RJ7xZ5CRjboQTqsn5YnuX
vRYCGcEZPVlukZYyI+hiKQB9tCJ6rbLGdDt++/AS2jqep040NoTxYmeZ6rKAS6Op
BoFfCZe6IffVQSRwaIyIrneSPTrnNOpunajhjUyhJpSqrCwUKkIAZaRNFpJT+uam
ZCErTEPuglOpqC75f0sIsbWLJSRx9dB7+3QgXh2hNt1SK2mYUPzBf3ZWCrh4HSkc
KLabGqLN7bWrD/ZPfasmLdyL5c5iqAYFXUb6ilLpSwDiTX6QTaGxV+c+VMQITvJl
Mz9Rvf1pFFGYIdJI0J3ZuKvXen7jDZro5KYZUtsNCsxOt6UHFuuJyOlgiX4he5xR
JnfZVX75en4upwzsFDWcYGZAiU0M3NQM18MHAxA34+nEwiCEi5yg3PkJA1Q9ArGS
4IA40VYm7hAZ7hA4C5ooCRnRg80vqqKXYmyUQqw9tZEXNtKo/dUtPY0o6+UH8Ry4
I1W1Y58WlNep6ViVNZJLrQ5ClPoF5rJIwXjdbjonCZSnzzbGeIgO9bn7o7OW017y
C2lxEm2BuwsLPIKfWZUDya9183dvIpJ41Tv7+Rsb67Qmc7oGGJripDB7GqZAyyBZ
ZP4+34B5IvMvpCEpEysjbt/U8EnD/t42vK/d3ejs9E5mcvqzBDrWKWdhzrF3HIWt
qiTDUi3PDsq/5/zHP83W3dSID4sRZtGSyJhZjEHmBLodFSDqXBAJghww2sGWcLdn
+Phbs4PvzVks8uqaSv+ikZ+Np13oyWQcs/0plpK72kHtoO4VZMc7o7XKd1AKMB29
BP28/wjuNfOrbUtRezYNcG5hC/af/HWYeOTgNVgJIfFQkS//qWuXNET76SSJbU+g
wa2s6lTx66dqKsg17i4AlN/H5cPQ/zwZLFB5L1cVHlanN+cw9Fy4ESCd4zjjXJRk
Af2+S8zT92f4TGq+bMxfwBYumBbJ727DkEODKpscgsOL/QJzndyU0KUMWN9cyo8j
jqbtkAdTqHJfGGM2uRmpYS48dnHiUtRhCsGndng9C9FE41oiuct+lBWHpdH42tHv
3t8kgKZ7xOoVztAXLHVsam5ugcMLgFm+rHogkM7Bvoj3Irr4RHYtuW34AU9CNxVw
EojAI/mxBesM3X2PYs+ePRlVvSxNAq6GF4EsE0Ay7fXvPhdAEqXIO3sOR/gROBG2
7ZJSyqNmMW3SHpX7iehlmkU11sYihq/uXjOB8IRpN9tdUC9SQSYxLGHqACDJbSTE
MpNTBzgGUY4/67veaBsG+/H1zIPZ95qNLJQrz7LI9mm5FWE7/GWyyEaDdPGER70i
ntL58dRNvtE0yvoowQ8NwuSA8rXUoH2CNjeiHv3krC/jwWpRLjRzdUU3hKL9huxM
pS7WOCkC99AJ3JU0LcM5RzURxQk9Y962fM80Pyyh/4+fLYjZOIK8lRpgynOhsS5e
UJ1/UxzYOIR5Ynclhh01u08RpWbekE6+QbriCV92AS89NNRuOASgsD2EqQawdllu
1oCm6kiAQcQGQ26OK8lGBdLvoXWXQWxEzPC7yq6bJWSc0xXg4ea1ofKKon+AYW2j
9UD7UCFj8z/Rm3HaipJ35jEr4lUGzJ2oszntFZuyvDFIPSown2ZdT1VXbXT4v3cY
QWVBuf48kOFMEA0xxaDkvvxZ4Z/IFf75ooPDnzYn4uBUS5gRT++YdGFpPrW1n/Hf
G7NODl5g7kQmnb8coqtgM9US4O//i7+HaQ+VJegJAFLT15svQoOPW3c7qZjjpNBr
Rz5pn7AJYvf1p1qI8HxGu6Uvto6hYrifAmYKyj36/vkkaG+9R/0vKeshj8cYx+Ln
zv0dHRf2pTG1BUA72r8ICY67kDgSlA2bO+0BsbPez/gkV/LPQ7WovRGLHOb74lET
65CbvbA3O/s8f7t+X4MURSj91ASgI+gk+tWK3lb2FTLci580Ff6f+F+0uiMttppr
I7iTmluO7l0MrUGPwvkxUSCVwHrea99PVk1mK3vVLoujfcKor6OyMRg0wV/FNyqc
kFwExXSIgwSy0NctQd8aJoGl1avsYf7eJlDf62H/AKUh2COargQmplEnoIGntNV6
J+hUNvuD+Gqm9HnWlDEoBgJLB0xnhY6B7kCEMPKMot2Pez5+WwxuZ7yhobvliMx6
mKVzYONoyl/vAiG0MyWqRAxFzZEhx2NKY8oofS3lJz6lW43l+ldbbndzbbY83hQd
5ejVpKvGN3CjT/hFZLgOqeWPb/QvxUh3Up0MP5opzqrBpODopNR75EgTCi0EPWtb
2qvK7BoG+zrjhIBpj4Cj3mFRp+6q/mYBiTlBe+wEOVKNfbCelChRStPfG1RaPmAY
1FiSKw7k7LotdS7FjtLLsBabn6ozwBQAtcG/A1pewfAI5TvBlHe8bcvcGjCep0Eu
2QcrNGmx2oSefmWTRlNI9SmT78CNU8luMXMHRhs45LieD+u7dPctSivSMtzFV3v2
qDCSyUSWu/c4+VfytWuists6YvhZ03MX5vxHwkjz2StNSZgRQcbf7UL7u9ekF/Up
6hlHGyP6qeKPcIXoRgV4kyY35DN7ZeR/ZpIVlaLc+w4kS7I9aA78UTbZyeHBArpv
SsMN8CwXbeiYycvMuaDFX3MRMFfUGUXAa/iT85TvHB5psCeWRDpGzf7cxZG/XoJA
sD/hdJCb0bcZD64wMe4xDbkM0DoK1AzrlSJsrkt2gdyZFJB+EeHr3co/ywfqW+BL
6Qg4dHqCil3DY9AoVzv8/0l5UCcfGpSft8sYMBauLPeWRou8aKc9X3U5VtoVH7Z1
jG84TdrN+JqnhiAwsu8Ud+erhRiu+d81Z7tSJfPCvgathmzy1/W+5g4kBlENYHNU
Bko84aK/vrmpnltch9Hro1DRvLTpEWFP86AKN/bsg0MXcPIAMC1bKzMMoY4YMupB
5FUtaUuKvM6A7R3stcsdkkRjMnotIt6roKIKXNBuXiDMjmiye41H4BBr+JcBxknO
Ag2Rtgs+KpOAVOSaIDlJOI2YYXWrBBhquMjtOs9/WyshueH4gYs69mPFA8oETC5t
VBnnTofav01irt3Dz8MWYdAjnWkpndOreMlBMj8YEN+41HwH90ms1Eup28JhAws4
O93Y+F/zd7EUA+Eh1xxSYeCPuhOUmsql6TfCs6+s6jab4hhyXbAmZnfJtUQ/lxwj
M52RGUTviXieJu0rUTkkCF/o3xhWyxA3E8LF+IZ5qsbXsX5jvGLwqcuAFcZ4YCIX
UINmnqd5BMMcriZL1UM0Mo2WigeGZHBxVW31brFQ219E4MZcZ5oUOcaQWUXXcrUx
vevYi+0fUcoQTu7j1HqJ0bObscORNxfcJTGHsIZHj6BocBGpLGv2FNStV4UD6yXD
sYu8x4BxW0ib/QmAvBQJNTEz/7uuuOE7rEpJa/EB0T5MScQQ7pTgO4tiArlsqM4R
7HRgcUo6p3IOwu2Oo2tWu6Wm9mjwHhA7wFjyH/hxsD4T/WfmHwZUdV+f91plRKes
O24cx1pfhncDpPtB6YGPs6Xg3rlMEcxd3Wig/eB7Eot3l98ni//vzICaQJZperVK
DLJCiByqH0rGSWl+J2i7OBip6QSh1Zm/JjvXW2BwGT0Rg0DiA7IfrzIpWlEs43+L
RTxsu0OGefnOtoglx+4lfOjry2yxY8d+gT35FRh7tzcrk1Ll/BWygH9PQ+KR2Afb
aV6cfjttKZkLlti+pdpmS5kyVULpVe17oP2TgpALXOYPNnDsVEgn+6TaYhyEpmYA
gzHleSduBNizceyCYFyyWCNnwjvfSja+2g2a1RrUuMMoElWp8hZIJcTPyIPSZBh+
m46jXK7GqEZaKukYuzSjH7EgoBdjUupkq9WvK6Bud6bAoFx4mHHsIvfX/y60uSlu
qV2N59QJrzCPZp6JSrUT9DAm37RtZdsymtiTCt5qoPqKLeSJPzsPhWZ5VrBXn6fI
Y9OuFUdhGECxYgYDokKM7sc3c7QN3+ezfDHPi3J7jouOgldVUYO+scYRh2nc6rWd
HNt94wtJFYF82ANFa0q4XzsBGUM4BTUNX6jVdOxLOUyPHK91Q+3o/5VeguiG/iOC
XtOra547w0YV58kCTLXRL49iDx4vcHRyNxWs7XBbMPbcLb7ujhT5OfDuH19LEyQe
pEow5ce6NwGa/ZRWuXJ/ZIIQnMzQHiF0C25iYlJjhamv+HPUAJqwRO3iLA6pi4Gw
bfEHoreLomSgQ6DyA4ue1hqy026SLEhBLhaAUgLqc/KoB+H3vGmoA3xVYa0Qcphy
jzCLvLSlgtoJWv2ExUHjNc3b7AdQceGgWe/sdoIKLdOoB0H55DnmuUDeDvE1Vvpf
NQFCV48u7nLHM/71qG6rDPRtGGcWf1HaPP6RvTTsn3yRIsA9wbVQwx2DwMp1CYpQ
YaXIP/R8trGwbP0LIMT8nFcbQzR+Rs9+K0ClDhXxcnZ6c0zBvP4KcR2LkOvk0v1e
9QvzCKeq5dCwOxzVJUpimgpySaL0k9r//UdcB8KAJnlfy8Fe9oxHTjPE6NQezcE1
auzRLRo4UkMS/T1Y5jewDEs4o6zpsKBgTgCVr+TImWpxmgWU5BnbeiCHF2uPCAj/
fb8RRBLFhbZG3mBlJl4iohxVgfrCnmu2R4bt1BPBb1Ml88Dx/Slym8zvYcKktmQ6
Gqvd/46HHEoV08rqI1Rt+5C66hR46OUkc7hAKw7CdhT2jyZxtzxkcbaymw8Xm0MP
cfOnzXiH1qGrEM9aqwEzKW+pTxkdaGds5TH8e/ecOb+ZSFhZRjUHI7lDqUMFlyoh
zW9ChJeq1O9ektHRIOKaa1NCMdj+u8CIsTIxqSMrsYhLyoD9g8CQmSMR9q64F342
/EzWarLYo1u+cGQMpX+8FOLz44kA7ikU+1VKd87RjjsXahRZXTER4I64n4qeadd7
Z1n5L8KM52slrbIEj8U/yrMV/+bI7Xi/+ZISC7HMhdQGgb3QqHcmdXyIP8LRcSR+
/ZMi3rdbxRJ1fqWq1YWYBtY4SWeSnkLAhoTduP20i/Rjm8Dx9wXnqBIFN21IyCmR
riE1k2FogYEU3QchZMaqLLdgdALfrJexXnFHXqlHUTti+PDVDnmwP02dZdMBEipJ
lqPoGgl7oc+SqmcEYPVrIxjd/VPluOSZ+o/SJq0Hn7E/X+ZqOQSk7iJj0lD00U9X
nlOdCxEIkk7knsj+4LImxAHDJeTRXPOfRA/3JkZaLCupM3Us9wQGs6RqJ2yFQbor
hHoqRLS0XlJBKb3UJP+hFCtns77JohGKDhMW4+/ekO3OYdV/ZkaFKrmQ09eeJdKK
WZpR+rUmyZdw24A3rTl0BdVDcUcqZjOblp8AFYH1IbKEKzcJPd39WWNpnuMoX8uA
T0pI3M8ZdaX9VmrLlkp2iGfi4OksnQhkkW3i9RdtbrlXP3h4qLrr24GbcIA1hG7p
O9p7H/Z2LqHOHujNKpPzIPIgMRZWFN6cZGEGbtfXEbtQD0b3aZtK4g0KQEzuQrpF
PwGJqR5AkDgg62bLlOwGfVmhj0Hpxe/Rc6lI1SESLVV/cfQ0KuMLA2gHRGbjyGrW
7K9BPLu2TFjK2p04pELhHBuoJBemXO0T+R/FnC7AkxEp0qXyHyBOV6qvC8IYhRjE
XwI6jffVOdRfscb1T0/t9l95cxlI1xLET0QQ6sfNyRlyXBFE2xS1/2z91rWHlp1j
XLWYFRvo19b6o2rz3szIHAUGIIKNMPIGA4wx9pA6sBoej07VL7nmhHAm8kmTS/kz
NCgQkWhSLtrTu5eirwr+Lr+wi4ak/NIpnPj9qTJZsTNtnKoVLgN4ZgHbNuDChRan
nWPmgdCOUuBlwJAk47xxApUeTE6H9JemFdP8uaLp81U2Zdl6k7ESRavrFrvZrCm0
XwuVNkJHPj2ZtXk8PRrFJkiNpegSbn68kgSU5Pghbfb2CLaMU2OeyRf3f1vVCzbe
Lhm6MCywNP4C94UcllR3yIBVysuG/Zt6WWN7EEneAFShDIiJRDwzyok83wI0nmjL
40QDW1gvYCtOwYjlYnt5S7pMfmFc2xJKVPahNo/BrHtamnZP8Tjm17abHnT7eJNG
+hs41OmNRUxNUPeMWwE77sYUz13ulYMRKjfGBmnjhuCiFFZ4kIf7kkc55sjy0Ds/
I0I1vDm/CSIZo/xKELlaVeFpOo+QBTbyoPV21nMPH58XNDn5UBkjwpGdItSZBT5X
pcdMB/QdvZor1A0FKclegT7kuXnTZQG13h/YgN3Ueqdrmjha00CROQ4Nym5szuF6
ozHjm2naMtD4wbaUpsKYMsS5nOJZ4xzs4HeuQtYOoV4bif6aXsBeLC/T1ZiP0sjR
KzmUy/rrN+r4MXEwCxNOeuWGxa8S/RMWuPpFFN6MJrNk32efE0HUlqu8s1c65ZDy
VN0coWE91t4shrJynlf0hMhHR5vvqcncr8sAWfdd0U11aN7RT1/OmakD4QJSLVmm
j8hzKFVwQAEksOw6E7UFAonztMxx5Yxk/BRFbzzKxu5C/ybMMlOaIX0bARsfzUNs
AG7vnrGT4wHVgdqavks8eYuuv0JquVxA9wOptt+isV01yCvfNDeIz5vbV7QN69iz
0pSo8NKt0Wr7BHyvjVno/Pqc47VoGqCmhAGXIt4cILDionPYaPsexYT5++zE05lB
JR8nVrBHjl0T13bzPeo8im1HEZnenYPQKz8NzL6NHfi9Uttwg9CK2quI3qESzGri
3oHS29EgyZ6qm00Ipjz6rq0MQHUp6x5b2yKkzuUgh0ILDuenwVhLSAo+97JfeKTc
ZtLD005g/DOhjk3Z5kl+Ocif4YGyUw9Mk0/EeLxXmp55SybEzA7RnCafdumOWTHU
s2ickJmDiIkDAA7dOxBVTMv3mKjVr8qYVrSMv6Nm7+AlYUe5mweJVdMb2UB/g5nc
wJ8h3BkzrNse+2Gk4dCyGyXKHYIgdGfr3D2amHddM3S54NuNxhJbABn0g3HZ1KSS
jiwvIVQFP34DK6dQpIzkn7RtJay9Zy69hEAM24F2+dmxJKUx+6S3lyFWmve6d1uF
JfHOB2HMDVDveZ96ClpeOqdA/DXNF29+j88VxdGMD/7/kn9DCcZQyPNcbjJQ9OCq
fElnWzgwBtoHX3t3Bq1m3+yfTRuUbsc1uoaB77biEjYL3DJu3SRuPfWvihcBBCKG
eOHXGa9JnGrwYEBG7lVoSiYoxrDSLyis/BImsBn7dRmcoPTgqVy8JIt0opVt1182
YG+tuvOHCoJz58Z2cPLpxs77Tfqj+OfUkl4OBSZQ+B750GxHkpYftr+KlC2FKzt3
+kYucO6tarbEp8z4l2CWzfJ3laE0/1ThYfZUuWRfPq1Rs+5OmQbF4OUukbkjx4tM
UD07/Or5j2vxYHJG/Ml3+WzP+/DdDVD3FBU5flXe+mA13/RDhOHPXNV9fKjaJSgV
zWm3OqX9SAcC1NsEGwCw8LzNuJ81S/h9g5upSgVEoJwfwPjBEuHAxjkNok+yD4cj
8oHudc91jTe6gMYWgbgUShNAqHkkTZmQB/khcSDH27YCQvsMQihByl8PSOxdJtWj
peVKquBFMPAoXW/f9mgxwVzQLpPzvhQh+iHhco1zyfL79BKUQXh/jGObHIJ7Ic2a
31dlYMQr6B102nOUXxeWx0YMOsQ1AUWbcB1I/KSAPV5i6iWx3oneejKcGpJskQgN
7VdAe3vUvBh3OulioaG5gcb7LH/7SIz/JM16DycY5P/KovHrQxcVMhOk0Cc5B/Ig
/L7iZ0L1fqJ6CL7kRGqcoqMRL19pAC39FkkH7uCgGzCXKq5T0RXe6k2sOLc4f+x0
QvnMmZpzDGpGD1QiQdAmdQ4vk/p8XMsFyv66Wrp6TArcXW7Lx1RD2JyytkbomJ4J
bbwzTJAP/x/hUZuX/euIqocI1eBTz3a9VuJMQYi+5DD7uoZQx1C286szN6xF21Cv
hlxpOULeQpAtUTppsTtrUEzUi9ShpRVfjeHuLYXbkR8n8NrzwGsoz9ZlrBk8iccF
Toq/3bJ3COHZlmcAc5CJOJ8w6enSPrtvwWxaFnHV7SA6HxmBpvdZf83UpTO0x0MS
y5jljgw/+VABb7gCho6a0h+Izv9kjmWA8ZvcRSnEco3OPyhMOAm2YQ19NBCVczWY
CNObFpLUsnpMrxD4/AegMClBV0SQvHRD/4DJ0aMgjjYqOLr6JuZXKjcVtjikgVAj
f89I86AzBVWGXD9+Hted7O1MkFsnB3lwjm1Jb7CFPX72v117axWI9ImdO8MhsHOb
MOPNprvCRth2dJ8yIL5YdKmU4Sjee22TJ5WhY8hfSid/Lbo7CRFrxueQUqp4OMmG
ck4BOqG//4/MMrr0C5+Evl00JY9Zo0Wup0H6nfky2a37tLUQZ6vTOlt2zbIH5zxd
zeZ0OSIplYmrht589oO+CPp90KOlqdCfJPNESamVZDVMT/YR/UvJPE6dQdZxN39C
yqrhsdiS6n95JIK1jwJWg9sdYUu/hHj4RDuWxjvtbYbKZNDMR4qIjd5XiN3HhIed
RHvtRiXb02l4GrPpcMBaYFC0pq5z/j80+3NULNp4p6saY8ON9ilX7OQVWLI6Y9t8
SbSWtLgbRZj/8aIwCy++np+oHdT/z/g5NgPQdbch7TxnZzyK4bgw4DLUrYExhQyn
W9h05+WUhGrHh+9G+eaYoc21SJ2wwVvFfgBClXPtiAW6X1ezV6qM50W1p5WdPI4k
qoMpshpg5xqe3/S3RQNuTSmgQH5GDypQlCySN5uIMQQ9xJR7BWclnBHtKRwamRB9
9NCUEZ2H++qJ2Oat7PL/jbDRK+arqyNP03aa6XBPAO7+fKHDA121PcbkBOdFz0kJ
LMyNXI6DYPw605MkG+y/eW9f9AKtt501kj7wB1HrOCVA1TPWV3WQwBVzMGNxjV25
sVVDqMwN73fcfAD/zZo1dSaNSIxqd3N8NzRAwbNNdqpaAOFHU3n+jEkQzNi3pydO
ZH3ODxdx5OxTYj5e9tkuieGmmn4nLytx6wP7LLir8qUfBxnArHaTdHQviRLXneHR
2E0OUBGzZM7cElMZ390l4pnwtrXzBMWCCchzyXzv8iAMwjOMcx0mBdBt2VRLbpZk
rV12U8566d+ndjrhjHATWsXrY6+LrSwzdPH4/ygM7CCty/9SLCOynNjy8igBtraP
2y3a8hEB0BqKfC3ibr3IE4tTTkFYifi1GoAgnXle9N89qn0KCduu5GOTD0cfRzrS
pHiPBRiieGIiBMzOhJflZiY96GAG7x4oQa6mZoRk9vdWwt4VYICRXPBy37Xx7TGI
7K78Hs7bNzGh2rDNFLoozXALxy8m9Mlz8EzBhWNdzmSOwW2JS1+hieC+j0lab78m
5cmJ88FCOSbICBk/kZvp8Gls+Chg7RiPeAHts+5FJUb80VXumP6puomc69j3AhR4
sDMIjl80F5eR51YqW1NLWiMbUJFY7EpD9UOOCMDSBe20c37B4NNyHVhCatR6ADsv
nN7d8VyEg5P/hhRwNSZ4nqmCjvRswSxxBeX75MHV5sh7yqxBcyTDg+pZAGGGEzya
6vt22hpq97YdfwNr25iUpgi9vhtO2diwcu934HGPji0gZjB/vQdX4u7XWTPf9UcL
4rYDY+4xqbTbz64G6pmuygMV7iFX3aNFxIBBOHakhuBaDHZj84tQ6xylFkmcrEab
7JNGyF+FUsCmy1ELxvwFJgcOpPAFUBFex6wzvhOTqetKexaGHD2d5NigMAeSd10l
VARnM+2siR5ym3sQ7eWG+VGsjpNUSbE8RyU2G6kSnJZxgHUZgBT/hhZ3AvIHb3lv
5htwR27YckPJ6s58wvtPiegGKiGmGD9P0U9Qlr0oayT9+UKR55usiwpXLe1SFCKp
x6CT2GwEyn1iafnkaezkvosHv97HhfPaamSL4e8ogHFzGL8SXi/5MryTd/DzmuQ9
TREXbnHd04+KDRCC/yCAvkrNbV5O1g/CVioxP9p/NEGfjy+fuq8BsFCgzZJ/GJgb
4hrXYGvAww2kr/B17P0WdF0FGlidGMvkLPKYxE0HsmK3QZT6p0Q6TW6ldjo7lt21
w5VZlfHwbsD9qsjURguIzdQizEf8AAdMNWmRBp4RkFQ/t9f4GPFPSRs0BAqq3dn3
yQcKCwIAkowJub20QAFvVW7wQhoUa9SvDQBsQpx6PjXKXVizMaL7ijcEx6mOILhB
KwnDnB3s3Z3VYBjt873cLnWd8vQwvqnM2eZP+rR3GNdPtv/o/sBMp6X9jHtx21lD
PjUEJt0i4QJsF+WdIA9sixhPkaEa04UmZvHS3DfjDPk9qaPjcBoQGHpP1eAc84dv
imiCUwgvHOCRYnPYdaCMEbeKMmTwxfZNDwTF7/9wTNN/Dtjum54rpkL6jX44wSTc
GRUtdZz5jIKJ2RiDzpiR6a+hq8DYHMJaKMn5pS3eoKBuxHRz2t4wDzyPDRlM2Iel
zvQuKYmLPfPDWSUG2apIHhBDlgyfZ/yWehL9V0RnKT1rAFUbjKByFxU9zJ0i8926
YCzWn0mhQFVcfzhES0mVImPSRINagTk3UzIWcZpP7LBPQAPlXlvEj2rlRMtYknoq
TxXgdubsDXloLteismP0hujW1L3CrIIrGlEYtcKFc2XsbZQtGx9E9nOsnYslBbJ8
K/maW2A8yzdHFYVTnWR4GSe7ProhEkUEc7JYxKdQOQdvRndWXhbzo9Ln0tD9rC42
qpZtlBKyXVsl/ZEewDGVj0AN4p0tnPw8iv5d8mXKf2GjzN4qIY3Q0S7tY0Ub+FHQ
B9PDO/mBKzgE6YET9RmICYjLUQx9MEDLbZRtL7GfY4CN8iV2VuIuVCdBLZGSbvPz
o9kEQAUIgtocTAcvNefvOcmBdANaT0CuFiUxlar4VPLlT0S27mGvCXCaO9k3kGFI
SdgBYAPEyWZzAwkge5k2u30f5cEbHyRrTo2D/BSIaQooPlO1ycHJ124x8lFFZ4fG
65PRb5xxmsO/kVXzhjxAzxoQtM/f2TwxgrSkVS0WinvmucRJCR2jewW4rmjYBrN9
sGd8aT9cIVOnH370MdYSPAE88TyvzCmbp4uxUWgY++dpXQ1VE3Zu970f0cvA8gtV
rvJ+i/M0vNiOwBXKlS27vdobQReA8HF9uBEC1QYZPg6ZbpknuBHvkWfzt+sBxk+o
tvCBB8VfVNOXpdg37L2SkzfqyyOV22sxaXWVkjYI6/mThzbeyWuLMrSi8EWDl5Gq
3G7hngv2KlLlFG+CbBUsSYzW9SrN6+iB3BgbDg/PkPSN4neVdztBcZiDeeBN+cr+
yhe+szW6Zyf0gNiNeRA2jMq8FVxsTk5khsRGteUPWMLggW3Sh1akLd4c/arXzIdO
no1zo8Y6+poEmUOi2mNngMDhpwGAKRdxsuKWTzZ17akZ8eNoEhpStDsMB4We1D1c
l5rtqNm4booOOJmvDWlAEYQvLtA7ke+GoWqh08aaUawP9SBqDIon1gPJ4avDGees
5q1BTsCAzDTwoSOhE5emhDlKtFaWtIxpKGTc60AQqhL7j+0W6gHTc1SnTCLP5767
txhJqhZyDDMDqESQHaiQoD+56dniqvpD//3N91AVrqXeDOIxGmANDWGAoH62o177
0Nb2Znfaeb3aAjLbUuzJpUs+M60wyAIiEAaBw2GdZkpiGOLhrkX9pN5J3P6joe1Z
xnOouA69d7LtgXwdOez29hgszFbejenwDrCBVMIPuV9lGMVtZ8gPBC4ixhUcwWY5
0CKCATcApMGLAdcEI9aCotzn9AIYglNzcefw4iKEEXBM5QAZJMOAel2+hCrVVtsC
itK9RNEqlcUDyklwJasfoB1mTD6Hwn0HRwkUVLgltbCtXEVX+PVVypxh01vkdhxZ
K6d3jVfpQBhsQwrHY4yT0b3mQk0/kPT4Wrdshnl2zy/Tn+FyqDF1FwL1kNrSWjWv
kqNKnepoc2pUPiNMx0b5UIeejbFooJ8OQFcvxqASskK208dE0cTkcScF3yioWOTp
s65Ff5Dl4dqK/tnL4DmXS/4sES7nSLbxXGKDiPzlpBLHRlZ8sWgUR2KlpSGRIWjg
68AIRxPe/5t/xEGTLItizuIFZuOPONQu8ExePp4KhrZps5p3lKRaQyLsNBogF79l
GpQIK2niTpsae+G/7cnLl2TBnH2TOGwcZEEcBhPAACK0TZGEqxtlAxBDpAmFQ6jZ
cTLLEAQUYiz6PtX5NFOCJ08dQ+GZE9ZDB3GPGMlofg45k2qozUt0nTIEKVMHrOJ5
3M1yLBcopPDjwKHfhw0AOHpzUrBwRGQS+wH/x5zcLIsksRtJDnupS2flBazL/M7S
FsNlKK/RRLoPy64vv61sVfSCOo3Qsy9iJRzOsUGKFtwUvSoAYnpN5lvFrOvd8cUx
ReBrFYEObKYVo2zvZxgBD3NYqA70GrD1GaIm4N7RlkV26TXRaNQ+MYOB/B+grNpj
48XoY+akobkHA+ZwR8+ONNmhLNqb66KwMa/NKejKkvZbNDP/mAdTl6cjkCigaUMM
rHYIGQBRen70Wt6o8cRBAw2X7HfmV2uLq6vQsMUJaRJFc8w6592Qy8hV8W+SRgJG
NIr3Oq9RKfO/0ifYqI0XxmSCW2e2NFPjTac0o2jfVdMyAwp0iX61t5zWabQcqHCc
TqxDyMv+795Rg9mJRzoSLpap8cSa+EYd4c65e19fUmu9U/9UEkPhVfhcfqPMkriy
b4Naq3Puxl87KYEjmr0RdOLvVDD57SDkd0eW8kQHIl5N/Y0AC583xFzFADc9IpMZ
oiNn4zptqQDPkxZyrzHn6zXkF4JFlyvuBaQwwefoocKMrT2q45UyOr+uhsS6Rt+D
jsPth27thDfpy+AQO1WqVgE1GkiutMxgi639XtFE3SxWZpA/NDsxLbLyu2F2muO7
c/6pPK0c3fZuRkuFbTZf2JjHcj+YFm/OezIgniCylIB9VRwpURREVjmK8YcfHNnS
Rp+6JD6UiDgCvO+PfKDVRp11kisStyPz3IOCTR789WTPingH2hlVga2jnpEGNZ9F
pS9yhACb/tNNMdMqKlscA2eSKUEVZSg+32rJwzYqgwP4XH5Pd5+26Cg8hcJ5BLAj
YMyubSOXCB0qc6KW/mfRCcj119P8S8PSjE57pIRlCRcG+fLxRndgxLInpq7oCBWc
y2nRagoET7XSSiQ93hqbSz16BMvGhw+UcLwvjW0yjvrKN8V1CLYvyfE2qLeX8yrd
qBNrK72FLX21yS2gYDJUSzrC1GCmS0bx7w2FyfT0HpqPyrTdSx0PtmF73oqxoNhf
EjCzIt1lD33COz0cMimDW+Q6S+vaZHifuDJi0B1Z5dKWafvVTOPNDyhrH9p1S2mp
aejMalG9BOCMoatgFLueybMlO+7U/SAoifT48INOOykAthiJM50qr8qj6C1vtcaz
4dRV8RQSCCVhe0IfUHmM6JA1uXU8G1S6tPiGh05yZIb/aYd3Vov+mXVeKpCNxf+L
piUK4I+ijuP/4ecc4vzLbU8oLyx7uosK/wnSQKztDvJrNvsIv2KoUhKBz9KSrgEQ
B06Xi3+p6ZH4uzmaJQsWoHMxCkxNu4LmnC+uBC5Ioezp6KL4QU3MYuGumyoG2SYq
Unf0QsLW5842k5jov2gj4vadyZR3Wa0mY+HQlp223yUyC02atGIoP3/3IBBZj5w0
mXeLlF0dcWu9sCJ+gwjqUUXXs9PmbC1bvkApFkZwZHYCvGMobsMzSlN/cJUMHcAh
s2KpMc32rNlRVNusNm+vT0IqDbOsXDuz8qzVyo4ieqFss7PZrhExrI2yfT+dHMbN
VE+5fwerE9ra56apBQPqpXtKmJbnoWBRzI4BhZbCxoqx/mg2wwnZaKoQYUAW8fya
pkZvFIXEziAbRczlfK98Z5RdJraT3rcL6my4XX3EUBx/IUHq7e0VupBpzxOKjxfx
l6mDyDcc72Lj4HgJ5SC33U0C2mh5F/RPVXs9KsGLdaaS6OoiQlrygPqNYFN9CUqO
tVN+AEdh3eGGTfismCp5wsiBQz1aUDLEBg7gSgLuIhDeuWJzomjXCVtvPByZci4d
EBskhmaiOQmwKvnfPKDpODKIi+Me6wCjHtY8SC6lmn1amFzIkjwcs+0aQUv6+7dD
7Ekm1ye9hC4udhztaGSNlxb0ulfBsw6oF9/0XXLfWJpYEz2L+HV2RoZsr1HAJICV
u86TYeKX07dCmOP83UYVXJDuJiwSzC8onX8NLCZ6HUwO3srVRYEKQ9ebRxLCncfx
IPIfPRMse963zO7DbTFC6MHpsEHJ0JVYJlsXiWthonlXUybs/3Oc2TFLMm1d/4wJ
4NGMLxaGXzfQxAFCkGTSB2I7ARfhcovS+k6HoGzPD97/TLF0XCSE5U7kaRXFCx88
YUJDSAIJpvfoDae/0yRaOHU0sv9aH4mZqmqlG0CTwZNQHHAkoSDPOGc/6UcTv2OM
4KRAJ+xADL+mACfcOV30sqeHcCvwCNL1g460bxPSVGqW9S9DtqOhguxIn8ueKSqc
BW8dr03jHlemY681dIABPWLW9FHONtVX6jc6tL7htdO+rSWZ/ZK7CTK2fqn/e8OD
nFXaVpholQpFMVi44VIKX5SE/aNR3dVgjVAryPn/3HY2wjwF0q+DTtlRq5qU7a7q
ezO3ot5NnizmSOXRO9XNrRMbXYxva3mLljprsDYF9PEiNtSApMWD8trxR5EPYlmg
LRSn1vyjQDz3ETwPTHq2hV1eAADN1CzYOxV/Sq29fMFPP94SLViylGQzPPiPs/fA
c6qY5IjmsY6w5XnhX1uR96+kT8rpRWWTRkeIAqrnWqy3nVUcyNsvr1StPNKNkUTl
8MkyM9nPLbIY5G8yhAg36ZnyRfYf9/LJ6DfJgJ+89DrSHSC6aCAJ4ffhvLWhyiDs
F1Z+d5Ze3wLVLWPvPjlthimMI86MUAxrkjIBKVYfMuvyJbN35du21gXJ/wsB0SEz
sP9yTdIoGJQEGq4Dn47DAv4odGJWy/vcasAklpxHtXwn1aIxd6o+RUgZt/7Ddmxa
OKGyXZOFmlGf8MCZFb70mx4Uloo3N/XTEvej3cdKNzJqLTz9Jk+u472yAk8LGm/1
w9UUPVgRKwAQ65w/GkrGn1dtyc+vnsjaABxB6yWJc2VD4EtzJfnd82yo5YZ08EYI
4Eab42zx7Trn7tGHzuDsfbxVfT7GXxoml1UXhehT+NDk3vSmj2pklTYSt8Xk1Azu
AnTdz2sgebJBkrVvOQAQq05N2M3sc+uMh5N916qe6fG7J4xjfluxfZiSe8THlQv8
YOc3fISKqF1AuokYxDxUTqDB1yRuxoH64W20k0mmampC3Rk5wrGm2NQNpjXmy/oc
WEDRcgnOA21J/Dok2sMk+3Wun4Vns1byCJ7L9IDw2iXognQ/XF4v3/ziN5q3T9vE
TA+UYLanBzrkpmjmalqrD4WPqsnHDwudBG3DlGD/6ZvLV1pTfdOCmpIv45GS9/Xq
gQtUZqe8j2u6eK7HNJotQWD0XhuztFMQ0wMT/nwZ7SYlsawClm8g5hOyQZJW0EGp
8TDC1WkC2pYhNguc1YmktPRJQ76xzjaENq13J6ZTg9ZAPHVvb/eT/Rr7OHmgUyR0
WmaZOLwDG3bYnOpyrmAEum0JviekAYwVpXqI+deE0OqPTbn/mtfK4XP4+V4gWfOB
IOONLl0VK9b+H/sbRNJl8rQT/UKbR3T+YnG7FkgXpdPk+g9gqUoKqPgcIMDqKtZB
pbrVBOtklgPLZWinZRQjt/YzQG7O1h2S3/vWB+EWBfeWVZW+34PRUEx1GlfrOkaX
twhcPlrfch8tJZ4oB73YHKIDkrac6IFynMMx/fXsVn1GfDRUgdayluZyRRcxngR6
Sitc+bbM/BaxSExHREHptl8YIWspAs5DBZ5s/oCl7e8kUMnnClEjO/JcCGEyemN8
KPQb+tY8GJj0Y9hbcKphgQQmxFikv6POEGh+uaFUR59QDT5+00gz/OjZpeICB+O1
f7JYxsP37rwOro8ySo7jRlKy5f8cUVNVYn1Dm/lwh2ihpFADNrSmxhu3vTDMNpTk
WX8zsGyYDtm7NJC3wO5kvOd/w5jlvfgg5EJVv8/fau3n1/liWQwXXpHSEm+DTcZR
bj4wKIGoi6S25YSsPSW3yLxzzGeyTEA5K7u3BMkexMNLSxWV39jx/cUq4ip/xDyw
bLykLmfcKYbPcCeoKxy2KLo2co9xYmclHWnYpLU+bTjo63VUTBLDfoRj82PsiWRJ
fpQ06PEykWeRRo/tz4uIS2V7Mu8EbP2HILrdQ85ZEYfjy2UpZgzMoJo0MvGXgs9y
AK+vhl/NY9dkKWWiFmu5PQxSpvQR/KUAj1uz6GRl9KDLF8tGyUl+hxwAJPMBm4hm
D8WOnCn34XCSK31JFm+DQbMjl8uorbol0GzXdmIg6+Z1eMYfZVZRT97jXWVWERTF
ZDO/2JBFYtJHRlqGMvSvihLmOCsSPz7S0Yz9SVl5Fbp7GoVxdjUluaR2oxb+vRbx
8QV0CxOWR6O3pcNfgNJ2MqLPG+LJ/en5U0fJYALyQXj3u4kR3WclW6jUIi/qKQZC
+aHRTn+ZwUO1KuT6ftdNnD3rwjpGfzWzT9AA2sy8LdPjzoFsOSKHKkdElaoHf8PZ
4hwpCe8NZJq2FNdqHqTHPyNcj7aNjB87zbFYVZ9ffr8piz0adgHwIRXT1WAHimYW
iC10DjpBdynUH1TIX7p3mWZjIhXULqOP0XcDEa4Gb8PMDsG8SvxYq5Sma/tRB/zs
x6+9dxbKvjCQWtf6JRDsY7KTSICcNzGd4B4O2Gfe2YRUS4gVp/O2CDjkviRHpDHc
hCvv9AiPYp1Oq2afRwczKxvsgxJtm4CQWV/n74t9NIQgXoEKHYcMdPm1loZQIGe8
DgBYmvvpb7ViyvFnLY34pFacoZFtTCd7xEjWK8EVP/aJZbfwKlrIv/+dQjlsh1ik
Qp9TzWQ6vkYPvbw4CcqquEiAjW/TtbS4Qq7SmkpSgugmMeYAU8f2GZ//rSEPuixu
m3iEOBgck3tlRMKqUdBJpFLihrhZSoH4ht75AdQX8zNbqA/feUERlgV8k4xB5KSd
UZG3IHVlAKL73yMZu4LpUUnv+f/IL5D5XDNlbGKfjJDslDcRy5nPGXCWJedQvND8
+I3X/+50C24aj1WqlAi1nOY1ciXvQdDuWmcerIUN4ddIfangn2rAhkHgXUObe2p2
QZNRTho4UYcVrCQqGg4gZPODQkLOWwOEcO/QuVuvsaq5hYk1/Umu1+8iU14Z9I7s
d3nI8Is2qfNjnEqracMLW4lStu1guAc9iD/pn8oiMmd1oQjpwA6iDu+MyLeb1dHL
mvAqNgTlzWk5ewO1ceIWHNtAZJVsBDQCW+tsaHAHAYuZzgijjpzHz4sLm1fTce/D
JDsfTrnn8rG6/K0zRV+Cn6dh4sdhJvmev0tLoyzZ0w5uc6wY/SLBfe2YKTuIsJGC
Yih4oGjOITJh38enQ/Fb2hbs/Ioj3GM6Nh3Vh//kAxdpL/6lOn5+TaQXA0oyLWAy
nteJp3z8gVmNw+QZeQGLfb8yp3LmsQq/z50IjwSI10zXk4vhjGy3+6NZ+ZEin7bU
6qHNZta61lFU7WzX/6Gh5AvZZNvseE7jm4IkTQC58L6SOsebbki/IoIS+DJDE4Lf
HDQTOAIvnOAoImKRaRONeaDeka1zO46xHy3gICWX4LyXXhg9TvfVXPG8T5z5Bime
OtQ4BmhsnjWkG3aiOO8k4y8ZZN0jd6+Hu40DMyPGxGYOlQcM4useMngO08zszP7W
Za6wAsNBJVX5Is999Q0xs+GRnk8lkeWZnOhmdT383VfPC+6a5SquZ4ChfLdVXqOR
4DZPJqdS/Rghq1dy/pGkGbCEfO0qJxp40Z7M9cLFUQF1Qx5FLa2T5fzVPaZ+0Kjl
HjUdlyGcQiErm+9QndZkuDDofkGjcKAXM7JDDTp+kECyM/fzDwwRJkAtTBP7HFHO
MFAG7K9M80mM8AX0369HIJ3ayTAlHrdM2XMQYA6TnegVe27hihPW8B9tjXc6fLev
Yt1c1+InGvaPcbuucSK8nk7C9gTQPSgMcfgQhmKOjzHT9yqt6mzsd3XBzkymj7li
+QjYYE7ZnkaP5f0KsA70bUTq8EvQK3E5Ebbnx63gXPksiePBBqutx/43GoimtjLR
4eyDfzMltk+LVxVX9EJEA/S5zH1pcD5f6fLpPb4vrFGrsa56x27nJypkA50vqfPN
hrvdw625/Hp2szBm7XTCpZ0H/ZtbYqMioIVrLOa5H74rOtx43ezfCt+a6SePHiX5
uvetB4vmeZd1euyAWM1WGBe06brxJzyXwWCMvQYymptHHadSLqV8MhMA0XjQOmXs
PpyfgNGndseS68bfmjfVRzkdjnr4vzAQFGkcZvkpgtMHQZb64ADq3vaRXDMb40dU
tq4exA2YhQJJglqrpffQ/5d+LBPmWHJYyAFgKm/aI2BVhx2ijnGXoH1WF3k1zIHP
SiPqBUYktYa/yco7Nf3vOKhSKElacg5MeqXosRvJh7AelMbHDCj/G1SqSBXSbGL4
wIs0h8/2223KUYNL06seAe2cFUUNTXkCrfiJ0kgIRYtdYk7Hx4LK3SKI0tM8Qu5J
cWfrP0ZQZ4iJ1gkJ7Eoaaq9OwA+ZiNJbhNj5Nl848VNujqsH+AtRJf3k0eBlJv4C
Q5dNWS/C2BN6I/sbqUJzs/SGFkpPmPQWqR6pf5Y7xC4tAF3VdjpXKaxmlZiSBZCm
vUuMf93Kiccm6xCGpM/hm8Ub4QaRlOifJ/viJ7T081bVsyJ0fDgJLgh8OSzGPnW8
iJgNEwbCiHLeoBrKSrgYyReGl5BeQaJGTRxFM+o4PrBAi8D27XZZNC7GwNKfop+/
YDBk38gM/eW/bCXJzy8kwsvRJ6vB8cQlStaYl6jzTrESs1oWhvOGYMItH9wdjK9z
lMuHDNtqSl0LwanqLXan3D43mW+iY53s1dQ7U//yzX976G1Xq/oKnYYZ3Z62oNxQ
qjh6Z8LbvB0lz7/bZCf3sNXaihFhrN65hrxYiuEQdghOfyHBOEMup8qVb29I/snZ
3UfltppfwHzbJidlX0gJfPXox530piLelkdZX+jcCRJBsCfjr9w6NGmRk4UGv4W2
qUEwCwpwwNd8bgGZbqfDqA5RRUsLLR1Fj23ehfw1mMY0HRe33gPQva4Yp+/STEK3
U6Rx3oPCow1PNXpPrtZn5IbanOKPf22kzYIq1jtXxseEG0b77N7KlHz+eD7e59uV
qJax252CU/eNzYLBcH/jD+SqFfTPjXjvBE+GevYLDw8IgOPfZBQnbW0vU7QAHhDs
7aRQhYHAA/xgu5fl3OlXxSwdDG5ZcLGloXJ/AsyLwvR3RducTadGxt37kPY74Qdr
G9/Y4dp+JKvxSABmL5Vn0tANSaM/W9ZzWrn3zYeLolrxroaa7ybwz5cCe6JitOwQ
GmREch1t8l2Q9rz0jVssR+U9p6fHBDSCw/IHfYp4D0FluPQQb5MixlM19WinprIi
EB3SnaH+38crzDjC6TM0VEayi8Zi+J8MlJErsE4349ku4eyFM+La/qehwHpl4Mkb
gP/8r6t2yIAfFOOani+wANh4VZDIlj2FfNhdmrqDtRCllRJ50QshAUTd1hHtChTA
B3KBxxEF9hKTq+ZUoYB77TNiTS4Mi5AxjDCdeFyR1OoKMx/bHPCvb8PU6SDpvwAJ
MgcZmZhg2W7N9X8B/s8g65pZoFb/QR2E0N6dYjjkvFZ8slJyupeSAw1wT0hSGKRA
RGHLuJA7w/QcdVsqihyrUlxkpFMLMmpm3Xk/Ev3PYHa02lWnCRrmNZS5VbwbhUFL
dc6266sBt0LwH/b4PbPW4DW69o1uvcHsoKt3gsL8e/gPXQQByNTNe5kRAqv/s0wi
8W3yUFe4gk1Yg05/IqQ3V/oNxX/cazNvyG3xB4LidJYJ7cfr5rdodcwvG+m3kLtp
beIL6NldZlA3osQivj1CpgpuwZrIQRL92HHywjMGicHWaGBJ4qkTGzwXP091s8+b
3AqJtvqpHeJnz8HTdZG+xiLys4Ns+LVK5DAe1NDZWpk1WmF6qC8u38QoY1aYJAcG
OBb4IkFonrxqu+nyC/lkQjzSVNl6escyOVPN/oYNgrJcTP7EZ4uxXlBZWd0YhEVS
IILplCuyP1y9LchGpQ1CPw1MVQ2TZ/PA0zNBpk+GgmsjmcOpWajhi5McAnVHzEBI
ONBx8aO9EZo5ARvQGV/6DILHQxgtdwgXNJdvhN1hrljmyiUi3k07l3Qv2twhYsPV
zoZLwrrpsM5QXfbRBKOCK+S8apSCzt4xsW1B4tLv30KWbp15rHC76N+c1VoI1v2t
3oX9DG8a5fOBBPgNS2LXBNNlyWX3zuaot0onQQdnpdY4yrcHhVJCGNDYXjATsWF8
BSLBS6ILw1j/o/qhBnTZj4+wYgPmmDlAu6fjS2X4i2Q7taN8qSp+1F11TUiAvNfI
qWajSbej5RnyhVTnOfuJsQtiAaBoEfz1R8+jYLYmtboGk1vYaDORdVYq6gS5mXue
ir24Y4i0ZPf1LPg+CVtk6urc+FDONHjwILbDfk31LIPgCZLmiV5aIQ0z/6UPMlNc
h2pi425mDG6wpPjVWAl3B0EeNsmFKCip6s2vAF5PF0eus4Jib7IYOA5+tDy1/nW1
xz+Qw93AmYmTC8V+6sC4H3Jc8BPteqv0sUMUVHhj8wbSbeSN745ZD+4kUUrgUKqN
jABWaY/0rUOyXrW4sbmiJTP5we6tfObnTuPNGvRHkeS+v24NHiXN9vYnJlwKRVyX
ntgTnGVyenlDjZ7UX1M94w3H4djTs0RkdrJBnNXrC07VQfAWUc0QycZS856sP3Ak
IsT52dXd++wF8JoiDSBnkeNasopufRRLpBigN9wMWKuMvV/ApBwHBMhlTEwLBBSK
9/XyOYBHmzP2Sk7q9u+g04uH8R2zDqPQ3WQ/qry0gjZYW7Qj6Yl06zB8QUfRXU8s
FGeAVjjh8tnBEBqEjyzBi/V1cH8jb3TQTS/fdgCxEiIyE/ae0+cf7//Pqpwv+U2k
I9EftZCyTeUJ2dUpP1R21VV4RVB0PxKdQwmJZxFL9YyhofwX0jRGSIDs+IZKHWra
FrQBdYBfLiEEtq6eKs9iodrO3jGMpEOCS6LXMZWTLKUnm/ES9ecY2XnE2ThsNJyB
t1CKgu0slv53zZGeijQQUb9ZEEl3UBXzyMWV9J3j/AmToZnUmNLs/MG8Z/I21PkB
KWOynaHrzV2PCfhAnOdox6NCmApk3wcaHbyubdGiL3UAuUSRlLTufEdZd1j4AYX4
fnpgToX2e+y115oA9x2VqwPViz+K6NvWkaCPA5fQExkS6vikkTCOnBZz1VXnjrW+
P29vAytX8i3SkERB1OO4u1GPomlLYq5yBv9qhwA+Daj/FywXdrm0lhD7aH7bW78b
N+RSF8yn9tnsifo2p47y9EKIIWCR5xWwfGv3o0k/Sm17mH4I6Y4W/U9myHcj5mZB
PavCoSBVFosS8vvgEJH8QDXsXiUCZdi+VhbAVzv0CRGYUolqt/JfUqTRcIQrSLbz
JI1O5rRh1IG8+EXDo5KWsdygu2x6KxG2mVQdSs36Pr3mlRZWlpSurmGXR0jdUvZy
fcO75GWOgWJNIHPfJtNaNYOzZZ2+KxBDHStCxpuYU9gX5GCOv01E9DuXo7mA7Ung
cbBwv7Z2IHlV3zuuw7OTPIICa6/VKxSbSkQPW4txCw/Ji/+kDyNMbIvTWHxjOgng
7UDkGwiVtoh3xKdiPPY/NapoCj90CfBkJrjg1R4ZM2FjOIIJ0c+7BwspN54n+rMQ
8mcfNNQJ5lNuJ/y6ChPciHydCxv9rHljudnioOK5FkJowbWWc+E11Uf9MUBZkMBF
iETcFW4P+5lCoCTyzssbr33prbZzgRa3a1sQjDvgVpxdft7TpBqU+pYAzxyDKgFC
Y8nCjsMkYhIMq/5dK9RUR3E5GpBfomHRMSe/bPIZUvLdV0G9um/VPkFo8Lg/u9KA
PjLPNiW51xjrB5XWYmZlU0BlbmgTOLdDQeeuJdx1e715infjtIli4L6YV2Hh7Ny1
AXfFnQBrBKAhjzH4/WKZr3UxyGqeIHxrEzkf54RSBslyn5qcDkX9kdYbIW0ZJktr
6ypxQW+a/uAPqFOpqm9KAssODGD2j8zjpe/mNVLMOz1XPNz9uJ1mYg/hRKboQB+F
2zxudVKAPnc7FY7a/pj4nQZf+pt4FCjGo/s8YhoUvC4kDbKe7x7xZECRafbHT6bu
Zbufp0LM89wcYP+yTAu2M8tGMHpbVFiynInXz6/e0NwxzoBRRAF2dnBeBree9q05
aIiifKpjhZVDTzCVfE/lPdDGCxQOGqccWR12h0ZkSBajUqFMXVXtkkhYhqARJY5S
tAGbJq/6uO2vo/ki8Hb48ht+HfUag3AUTtGPQw0neNNtdSlNIdXsPpoZc7LN582P
hyrFiRnpU1yVgsn2GsM3hS5l9jVRdOcC4A+Ywu9mTIduC6lnRG1PvydFf0BOtYif
c8f/VfNjKzxeZ/ThujCxqdA3nczJIDZ1ttRcXvg5u1ISW6bsplhS63VFf3fpujDF
Pt9SyPKDxOOTOuHQeXYOiDYKEzNCUIL/YNmKseN595jcVpEht5joqvtqR3EAtQvr
k3uvtLqRYmb3aXOPm5yz2dTb5xyaQ/Xk8HoPFERFNOM72Qe56fwW1WLv2TCjyIgv
j9Sm0RrzIk6pEUUlrDgGjadoje2hn5NGyfd3NuAEjM3+KsHQ0XaXooPoBd9cEAvq
MA+nJ+6349KglnkikgH+rwchJdLgVzImkfwZv3nTzoI5/CBAoZUETUhE+kpRKNXF
UtwU1R3r6zFiGwQV8T56sYIxVRWdKMdNXKFurccpyVg/5WvBc6dV1KSz1yp6d7fB
cdi3hoFfNXfsT20B5tZehsoElq/rEHeiyoL3gl1RHHs8W1R4n2D/UYlf2FSQO0jG
IXr2C9Vn6qiw3BnzKlf/AyIKGcbAc1GKlRIQB6wDzrv6ElQ8wXuG935GNNRJAAY/
6/tPuk3HAg/Rf/bsWCfiE9u6M9xVVyFFAIxsdJdkUqzzgLGReePij0XntnPs5/yS
rSGg9BvKknLEJLIg5GrNwAOPZ/kb66KeKkpDIZLP17OIzz7MzXI8+LrWc1u6yBaS
OgEO4gTpltxxLV7w3/3/LYIw0KhsHdG+MZ8n/yOAR/r79blMkWGp4xsL4jt+BnSf
8vGnj7kC2GTWnV83suYlqrkQkq+Biyv1bmbEPC55HkV8V5ymt8HPmmO3aDz4Fm8E
cO5bEv0iPANtXt1GhW4FYj2Y/0pwYafD5FEHgjnMHF/gbXqyxERZSABJbphcSaM5
NH80GQMsoSD7Y0EbAFHILg92M4eUGDUoeJlOnNM+uDBckxOBTua1BDBhRrsQ5M14
LJzbUTf0gl2SJwSmiz+I0HQX31Onxz+TXHcYnzJxyP1FUgASC9rpmpIBsiMJh9/T
eYLB/gOiEtizI1OcE20Bn5de1WUinhvzeYGetX89nYcW4Ve1HSDRb2gi8VOYStxc
qC1GbIs8/hE2S7yr2VQbwlajDwHW9lm/TOa9gc5R1fkK6aJF+z2bt5+FWmJ3fH+v
N4syLfC6aMIHqw+epb8ccutqAniH1IblYNTKRa98do0FxXKQulU9A6KSEdlhKGgH
u3zAE1J87JYVP9YRgezuKbFHEEz0oQgdG8LQA4J6gcr9oGk3hValV+RbhYvY1Xcj
qQWlU72YMWGnFP5i+1vyHbrujTdKRfJTs7c6zzQt+ct90ahoedGodvOXdEl4ZGjn
hLSMiUDop1GruRBJ8CwsHn/kkUhHKvma/IyyrK1o8bKMEjdYSgLFfespUqvU11GK
UN2Acxm+pS2iaLrJjOVaMKrQHSeMYEM6j1zEQX999ZCt1rapYxrv2G0xPMNfZ10K
KCGbB1m6cmpqhvaJdLpjPSbcAyhjSwjgdBpHKn1UJqbdT6WgHQ5v24gO/rrSnZ2V
P2AD9AgBL6N8JU+jVpIRBJt1/f4FZSji3IJBt0VzfQKDW1U88+evsMASVS9tSqcY
c8b5TWWKuNhQ5tFFmAlItsjjc+hgtzeBpOxQwZDrJZeg3TlccFbTjk+BVhR3d8xg
Qmic3bCxWetoKPQCXJrsic05HkQZpxdGVwtvt987MMm2yPQOMpidR9GJuncY0l8F
lYDUFjw723LYMjjMRuX8l2jCurxkwYD8UH140PQYzPiME3U9ErgLRh5keoOXXvHh
px0GA3/PeJgc7/amg65tybDDBeGAVZCDAPTXWfqsqikVbq3SaDIwY2rwmb0Qm4+n
sfgJ8n1IRXd87G8tK57XcVAEXXBGZM6+ZVoBIVRV8c212BFlYlb+zVG9luPhH9kV
0iAb6+W7R7U3va7/s3TaXrNUS33xbFGRWAbYSYLtgNoJKiMGjpyvPnFHpuK54SB8
ruk7Wz4ltExQI/XT4x7zDB1tSogT/HJIQK0G5JVpVjp3uiQkXCIkyUAsKTURyzL6
v5ml+qcBgO/MYsaiN62gPnCHmUkIiQ9ZOt8eLsL4GbmxTc91SRlcJzAvVU1J+H0b
rw6+uaMMXtA0VKBgHc/6NRVj4TIKsSrtuQGESdxrRe4XcoSvcyxuSKCW14y6syK8
aQDm4+C6qoFhFW+Q/ehmkznU2EK0Z/dU5VjudbA6ZsAnzNmIBORcKVm2EtDi6pmN
qADCdzE+wHhwNbqxS6Zg8KgS5QwbNHNmJ7CsCtY+CU/e+8PyrTnyv9zgpRJmeJTD
Qnb+NYfjMhfhgM8x1VrQuujEDa2a3uLF5vbLNQ9PC0uYvMfbwUCtmDAhTQW1Ts7m
hrYXk5UP07vqatXcAZ3jXke9lbE/eRGgYI9NAibMC/2loL56Nr5Igt8m2di/SfMW
jB+oxdQ1QF7JD3qhbMav3HN/5MbQGyf+8p+9L1hx1wQ6pr6b3Yj6czG3flFgDMox
8COTIqD4O8LnKp1nsGF7LJlokLV5ZMp5CO036dUp7HQacmTk9ZI+VEYJyVzjz28r
xQ6XYB8N9X/iYU/Yfw6PbWTkziMksl8k+DAKR4dsaUb7NzCpjDl6hKEptUdd/QRE
PAi2jWZelKyg98afM7bR4aJr5EtZsNXF2X3TpUQgeoehTUZSgYy3ojT9GMCnS4bR
K6Km0K4d4nCBMYgVQE8jk+rt0QCH29FNLXto6AizxcpHqg3ARPaltxp8ZE3dyozZ
ZHiOU2xcmrCZvEeWRH7Iim/jm/aHqVMFdAtEiNQ8CbUnl9S1vZc/WFlBD0DND6zK
gk3cxsqnkAZkvZT/Lz7m684z8cb/JPmIPFSlDXY0ECkC7AYpcQAPJ5pk5YEEZc82
ZttPDY76ep937u1VPBWwm8v3wQvW7ylJNaMX94Sj1jcNhyjx7WkMKURgkdy8VAvu
b2PuHt7e9gArh6TVnRLWbxqJp+U2Yz0VgLaZ192/AHIZ01y4aqy/2c45ZpAu+7IZ
D4t2qI5XBOg0ikD1Wj6nE8s+eqYXuUzMicDCS8K4Oo5UCjQzt5G4OLe1SfFIq//t
kCp/gup6lMz3JPOzNjWOrPNDulv/FuHns2oFLnXLT46q4I/FvTyO2LQI/P6QxbgA
QL2rqu9nmad4qtweXuF9x+zAEqKmoWAHCgNGPXIvWbCDJUnigK9IFymrRyLoMgpi
OlNDkMVIXaNx+MJik2rcnfVMbvFrE6BtaTGRnSJmkMiUEXUsVD8QyngKHM1QIOqw
LjDXwAn4V3TmRxIx0Vdxl4fpDMB1fIvTNix0jjaPgASxpgr7GPxhPnsTEfKu95uY
OzjQT0q0bIvaGNujieS1MXQAqjrJhxpHI0RSGIPGKJecdWrae6qf42JG8R3Sj8qR
H96X0dmqaaq2dkj1Bl1z/tE/YT0QwaZ8RKxiHKyRSCiWGnYT0L+oQZOJ6x/uJsOi
w3i1GMXrf8J7oU02gIM/8FrBEE3mOA9z71l1EpC5jU4ji5tw+kzUDJNuEekTW7BG
do6o5wqkhoHaOtmbqug4iXxY66b86ABlvBKxOX4es891xPNXshmJZxa6/XdE5/UT
WjeFWRahqNr3K2vUJLkxD6covCewrj/hl12goih+M9Ft0xRopt+QzqhQuC0th3I5
a+/dwgX4Hz9hrDve/lzCQi8LIRJOE0S3pYScKihPwm7TatLd/Gwv1d6yA9qWUNC1
UXtr+MhRJusQfJUuXwko2MtZNkh3K4S4uPHpVctDuNKIwMELuwKYTcHZtwusUQTd
JuWYM031LyazdhkH6JNUwCJ4IXurpHPPGmNlJBvj6MLqbs9ph1jFBab4/mxLo9le
rhTuTaGYyh9geTUkCLH7nAzj01jieKUESf17Be/xsOCXjyzgTiiV7WWv/YLDAbTI
L8Sa7ijr9VLBaEpgtpzuw8qut7T1bApHA7NeqwlCwVKY5ixaZE3ebtMXOBX3A2Rr
tVNpKk86Sc//0lmT6aPinxncKB+q+AMg2A1GZUuuHoPc0n3vvcKvGUSoP+NdmaaM
FL7f90Qg472oWfv19Ct3TiTFI6vYpwzpr8hQcsrQNGHLnE7uwVAZCctCJvAdpKEG
IXT/fZ6dBreexE6L3K8QZvfqVBy7Dc4N1ItuwSULpl3ezLhlTyIiKLFWmCEWFk+K
Xo0muz1D3HLz9M0ZKluUlbjyCT9UZtjPMXkucpOdwiMKi6l0Yn1rCRx5tv//QwOz
y3qPr/6BI9qbicfSU+eAjub5OyS5UNUyYf76d+yhwCEqnExGJhgvScAZ6sp7zvif
B5IN2zFjuZfbh5TqEy1TRxbBf85ZR9glYlfaxy7gyRGo9CRBbFwNtksuPmSszPi5
XDeAdOyu7nQTudjWXgvFjnalQ6mXkTHpjU3WvJbo30cDUyPPxBjSaPeW2jQDVaAs
NhOJGYOFS+6q+0NCJ7TqPNRBDTf4Q7X342LNYxCRguWdazyV2TSr3ZqoGeLBAzmZ
oJsazTp4fnXs3D7eq8V0CuZOfLs0PKODqicHA31dxUfr04cLpslKSv8NBme0cl2e
xw5xb5StUg7db+h/doNtftMTWsQsMLt946RqVd4q5C+kCI+QZlZGnyNDazOZsQZ3
Zaecfi6c6jYJwZdkkysumcxsFwzTmfwYzeRcH+bZJzerrZ74Q3TaXgOjaWE2BwiR
Xkc7LhUvJBq8fhcGKNGdpz4x11wTb2Z7aJBmhj2OQrlFHmO+9FJ9tPDfmTZR36Db
0nj5p8UVkO/hoMOaDJWYzoo9IXlRX6p94Hiw8Lr1Rz4TcOm/jYzSIVnRcbIsWfOB
/AlBPWBS9ndYx9/HK9Xv5RMa80ufwT8fD+onxq3UpvFZDUbfKBkHqAgOI5GEyqNn
xs13WuuW0/Bf1mM9+oMRVGtZFxl42S1ANU7AT+AZ6G9ZENp8a6FcMXJXjyz6bKrL
BqMEmLDbF45122JTvyLJhH8qsR+HHy5kwBMAWzNBpKSYaEtuzz1+fZ9psSF+9hfM
eaIGF9R8fcLj3FmRwtWxK97nrWxtH2iJSB3gppp9t54du5GymRShTHordEdrosZC
5r0WJeOrL4dgPT+03Z01G3wbXeYmi/wR6SDjHwZ46loIIAhlGY3NBwSzAR0Vxkr4
XIAbBdAf/OeY+ID3/1x01lSlCGdAyioh5gmcPAvb145q8HprjNMxafWPY4nT4gsb
Hq/UYNoRl3VQ4rjVT78/dQK+EsBFMs+8dExo4K3u95xuc195h8GjdbLvNGvIWVXT
ieCjqXObFKTayUgJNU8M1D5eI0EAzuciiRovh9+v4ereCZrv3M37SkNYDXhqamCw
SbBT4T6C7FaCzJ+IXlqJc8J+X7Zk0uKlBKN3ysPZKdGuw4SdS4Jy+nfCggIttksY
lvlGJkciaYoj+iD+l6vLa/61fGf1JIWw215bAZQ5fIMwg2dfB9oJtHBFbs/gN760
yduy0d9JhC7PmJFnQk3SPKyMxNs7gB1sGQN9C4fD9wVY1FqxRaybpaXBIEOG9YkU
KOW69isXN3yvWxqcDygmZcN5EBms73gE5OgygPjo+xTY+tr+ji40/phZ2p5RkaBB
zYwTJTKXp/4eL8n0uzUT0I5H+RScNs8Ci2mYxKHveJ2kwyQdv/b1cG6z2O/71gxI
o6l0aLXBEattwkaJp3rWeffUZzCqmiGWiEGzQoGgDNrgFBPN3IviNgh5sWMa1Crt
OiEQolEUylEvrPV47RrTr/bhvMK4n8hrVxSLLLnV+GNRMhJhPLQR68F+mw/G16lO
/tT11vKmcYdStq7gkzpC8fYJSdpgkUR8jy03do9P/kHBjQtxoeSt0LflcPfHGC5S
jTD2lOdk+ev4ulZummEkSEZpoY7AFgbZwzsNKxeIHTDtvCp3NHGw5hP0/Uvqf7ek
7bcvY2DsscoiTut7jGvwe305/VvBySV4nxkuLvAXx4iXSgl96jVksh3bZ7Fp6q9S
k/qpzZn9+6XN0MJYcNu8Hv32T/8GlQKicjmruS155eFMVpbFOMFIwhChGBRfTF61
SoPGf++H8OJZ5pnBYRfiQHbH0gB/uXrFMcVvbClc65YMkvDJZwfELshkqP6kwnPA
EfQKyMchM84aFml3G2Aqn+24uSDaZrqnu0WNWc0GoHVG7tf2L5WcIPR6cg1OQCZg
gOGV2+AUwc6wI1RBs0wwVnnZlUmLx33sy36M2Okk7a0BuQoKBttZ9WLZWgYyXD3i
BmVgy771gmq1jmrkGpwk7a6d0otGg/HRw7L7kheJ7RGdnAH44HZ+PP90HNpZgbj1
7p7ZjHSOflkMbALxn6J/wkxp3njRhytTeG2bx1g16pw8Q0C1Yr6KeVMmpEbbHgdp
X0kMKJUMdFsTwr6+cqVbs2tL4h0pwyaG2uuRRaZ54vhLl/LbBmsH4hl/G8DsYU/J
Be0O2XvugUvU2pzncbyprE56Vmg85lcHB4t9APeVijplWiCtI/WXanq6Lp43AXsS
EgqsJLRZmLrkqIPVbrt9ehTWb3qokBz0XF4vwaMNJ/qEUsiLqi+dIrfgQ3bjy9Hn
t/+99ASexGP5xeLUz2I/3URlrgMfX/uPA0kXAEpKASiJy8mJOHPTJGBmqr5YU694
O8/qgpqJ3R7/VpORT1/woklqsh9CkrvTxxR22ITjk+/CFAZqWMYpu5DNHx9ypwWs
oLW6hEpCCsdDRK8rziXjvvHecaTuEc+ZBjOlXx5sZzpnq5g1nL898rW+g7og5DCp
jMv2CKd48naQiU3K2K1edjVueieMEJIHXK9Fly8ivYmdP5NODEZeZ86/L9kLUGKK
DaEUDpBLWxV/B7Nar2znT/TEgX8VVfKTyjaUG9dSb9s/sBaki3ZnzOdmwHhpRqdl
nn4CMWm2CP37xAh3QMlbSIZUEP3erFWjq0NiQbExfuzCK6DoTJo0IVZSUmmDQ8yK
78VBYmmKTds45HHsaG4YzkCwLaqLtc3HxTc+2VgL4a/0kLxpM1/HzsbdkJYNylBB
3B8F2u1nttlC97wpRZUhag/1cBMfMVdK6XUz4eEPW5upTsRffotZ+75jaf/79jTL
1bjOYyd+805+R8y04lWSc/ANjWIy1okgUZrFnsV8+0+CW8zirQWyd295DPagC78t
f0Vm3jfXK+iItXPgt/3e43p0PbODFIC12RczY33GjStPWpdey0E2Iyn/g20Ea1jW
Xlli8unhfG8yJE07fvpyhZFRO48+WXvmZxd+IRXUs8N+wpjt4kCY+pQSaFpjFZMg
/sVN4OHPgnK+25cT6FvFYBwYQpEB38BTIdbk96Pcv5mjONbnAdCb949v2XzryNVu
fXhCQMJOdR09wTxJp8u4lwoLzlkR3HHeYNN9jteTeGomVPo3xMMdyeonig7hSgmx
fiSSMo8jCXoeRujXAUGTGsLEvaPB/+71ccTdqwGX2x9Rs0K50gpWTdPvi2fXvcIl
aitbVT3nc4hF+ZWvJRh/NL4XF7h3FU8B+VnqtTyo1QtFpLOJXRwJrfLRA9tCyv8j
EroY3tEHSxGL8euER0Dn6/qS3CIP/9BsZ13KBIyEJy3whzi83BOQesO8qIk/bPBJ
1lq0rU5Il4q6qdSGk6g7fRzIRjqVluG5yzoHSJl/fe2R8M9jSS43AtdD0y22ZB0E
OeNLmPOSvVGTSundnJZD5XTDv1veKgtI63w5jdfXu7x+73AfEvn1VyH6wQRLmicV
/i00hPE7MCdxFeouk3RjZrx1rTvsaBjj0JO7sQdTCpvdoDywKgXR4IT9jin66knK
h/zz5nBC6RHOrZ0VbTK6YRIv30Bw9FPJdCXke7usLx2ARioPCq+zRus+kflYV2QU
vcqSUNv+nA0y3XQF334O/cHekk8bPYDnlsgTrOfRPjGczQ77VTJeHSPACPjtuy5n
aEgjv/kPzXDC0sSiWAM0OMO1ulS+ui346XAkBNr+t18UduvXTZw1YuJGO3YRbx+E
gw+RqWkn+EZrr5YuKXMBrlNNZjLaqg6N74qhsv3itUqrOVvKblShGlig5TlTf0o7
kKR1Weuud/p4cVf9mpRrI4J8XEt5EJZwttrXVx65jP9qnDhzoPzX1e3Wygmx43nq
AvASl5WWCdTOZ6WoiuMdKEHb2kdyif1nZNsM3CsN9m8Jw1PdZWKrcS+wLnrB4ssX
P/fuDTLv3lqikxk+ctKgQnKUqYnebUD15qhAfkmPSgRYvcnbsiRnzTowpEBVBTeh
x4cYmfeAzFbzwPb7K28LAPpEMxeMW5BroK2kfC1pAozcdx1VSXfeNfxZgc0LLfgR
vhRfcNvkYbRnKuZhQJ95qLtNNheoHsmq4fMAFxAAvAcVqvU6dpGpTASH/iUy6TVL
YeMhWiWoeqkXttUzEQZPc7Vs4smoif2WiECTjHCxUvPCnVgx/IMPxQU47bRVliSA
tskHSInQyThg60pRYo8K5/k/3Xwh8w9x+AQ4f85xf/hcJAD2NLxyRId+McqDyRVR
3KIRazigTzKvgm4tN15xToTRZUyaPRn0vKKc/j+XzMo/vWuls09vyKTiRWkuM/vu
LA6lr0cyx9Cjr4H9MNfUxuULHoQkH/i2aEk/0vEkXq8AMyob4G5Pj72WH5DMPr00
BPtDfLHiyc382lKgR5t/3LvY+BHqY445T2Ia7lcfTsAxhGHoqWfMyaORdGLlTxZM
BOoIXFCyHQN9gr46DT0gN1xhDAm7c2jhSXvJw9qAWm8WdwKKgUHfsusTevH3i9Rq
giB0E6LWijTYA3gbQZeovMXfVH7LIhO4KTZy/tOwwO0fm3ZYAW99VlQ4gmCJ80Ft
YkR7HtoNJbGNeuarc5k50A2A4e0kWKli/hZHBdxHN5lcT2N+oQ41Zf4+lBOQ9yqv
PTO5MuB/0bWGxJGLiZRBULrbu37p0sMT9xFBqu6ewTtS3+fhXeXfF99zWKIgRC/z
DbyGouQ0C89DHIBm9PTFwZtZkHdejRI4TZ9oXW7uc85Z6gsdJy1h7eUwLqNmD0jl
icyfxMb9lQmUtVg12ZRfTRdZu/eyaT25DCaYQRJksSqA3v3vNbvaN0jO4IZziXbs
5v3DjX5Y7FGt2qnQc6BH8bhqhVcdqAI5sYUTcZ+E1G4MzQEAhid5Owq3KAUPteLj
EsF4HrMEGZRfSJfQGoFMni0wrODetS0odx1GvipcjJX9EoHm29j2zr76NJtuL4Bu
Yy/tdXubyaVg6hFmif/pYpwZbnurZi5N2BWmPkBY5g/hLpNuWDIneOrugTXqQ6My
46OVuTyKv/lmB21Yr8tykaxKOj5LFsNarXs3uFGGHrqB4tvAS6knsO5M0biQ6bJQ
QKYyLJbtAIdMRqx4thFFkc2pSPCJx/Es+8iukaQepUs9dGxcyJ8qr5fsZdpSbRrg
mTx9KfBbqWACUkUL1GBp1FTi8v5X8rK9RvhZqBZNoD+AJxhD2nvD6zzCezZqK/Fi
RAgZJQD3I3YIBJUw0nzOupF+r7RdUVqVlN8rakBKcr6qnIBBEIdVU/erpC72UkbN
Fc+mev5GOte0Y2JitN3wVzzAEsC9gBGxb9oKehLpDpLcNKNYM4T4pdRVCU5uBlxx
MHoc1lkwB7IoDOYRF5Y+A6vqbm/IssjUsbC0H0mkRKul+6yxrSN3QlMKpUF34Bbo
uT9VT1j1l3jhNxYRVZjwubxAMS8l6WVXWWzA2s3lXsCYe63w+d2LQHUt7ZhEcWLL
Yo8/UijycauOtjHDC9ZOCA+fAX2WY80CM10DHj+iaOdEX7EmlOm+JldutYWWpf92
ug2NoIIJZhoY5jQMv0C70mqLammD4dHqI5ng/b9SYGcZ3dG5E54QWgheclXsJ4T3
9GJC7UGe9seAO7q2C+VHbL4otVEurT9U7yIrJCSlWzu/P9CJ3qMRoGl5nEYfo8Nk
B7RNE5vNxB5+Jpk3kN8jCVjrADAD1u6tx/7HF8muNyf+SDXlpytxijdMbq48BDlM
9d+4CCJAKUUtFetjv69B+/O8V9G6jO4NVRDIRgDTINRduxqNWqoQqJ9cWbL+ZUdZ
lPZ+8aKsJNlzwBEJLa5FmsQmpc0xLIRjWPUelzj3DqEUv+mckGx+J3aE/1or9iFo
adRXio8g5IkgWySfujEirT6bhuiBbDL2syOr+O9IqXoS5T7oWTa7TDG+RvZU62jK
wIJEdOS1QoQI3T0z6Uz3KsidijkQAJBi9FxJeM6dlf+LmYmuVOgYUrJkX6ivJQZw
ViUU2kcxN4AgTV4K1vBQgon2WBWeZa7O0SEIySb2mbUQtmtuux5S2FYogamgGNbH
p7l8lfiXiN0A+aDagOpN4c0yGPn3f4fNXPTOdudexndE4U1QtOr5QTP1rBCJM+S9
fsUT2PxtkXaZ8aj1bDeO9EiJAYDn1r2wPERDNqVs6EdkyFHuSTh6QLpGIPCifKZb
wkbT30ABI6ziQvbRAdQR2lWF4bzrab/5lK/EjwI+ZnfRZnUAkam2nh4TCHUDbiW4
eYowshaSAgVgC/MdcR1KDEnu/XkQXRp/AcNwHeQTAd78fi+MP9NlcFZicPT2gazI
GJmu4GYiNghiZaRVGT0aufQBO9Sdi0TvuhIyoLqoDunlihjDzVKPOg2JYyUtDMCI
Nkr1Jf7eDKSC5vZ8yPXwZ+rKOu89a75RpGlvLnOo5771P9n5ivxbPLubLOMprULl
4c8VkjKK3ho51RFa+OU7fgDr1WN2ibwfi5ke3EgNVlIKo0wDipjBwM03xFhJoPm7
86BzHuY28k8xwljNgYFDyhzIYU3dabP9TcuD1WV9aLtfEJae/tJ9qgMe+/N6AKZD
2gUcghhjvz0dBqh9umCCESDCsY1XOGcIDVxDga/GTyKhKVz0UyLYEptW+ia1ZUnn
WX/ALpZNXH1sgB7UGClztgxGjP+S7CZc0FC97DvjZ0Dmx8lvuyQYcUhuGINMoJ2P
yK5Lgdgn/NobZRnR++Nehu1B8fIdFnnV4bn2EvErprM5j/DkvVfTyje83gyqZWae
0MilOahzEjmZAn7a8zCPspGsDdxmqLw/F/8NAwi3wd+eB3jObdDszmN8U/ql+pdX
qlEVqsXkgBqMpRYJIaWDisyVZCq7fuQyfDXjMj+8hqdf4MZ1qryfqtIh20PTZQKu
njf/467q2b5I2t8nk+xKoFGRng0mAz2eF1wZdYOSjya5G6xIDKxUNd8LcBuacQG2
r9T1OBpGRe7c6wMpNfnf3XVJB52ifrdRMV+1Fb5m6bu+YkxCvrNBgDvOp80j3LJA
TY1cjcHGc/ojArUR6BCBtWjk3BJ001h+qJccNSNhH/u3dWFB9puDvu4BdgeQk6P5
NxyGsxfHnceubWY86suBC7omcqkCphnNmgvWPWQse/MLx7J9BnYrT22ZswxydbuW
izxJxnkwHgr4dtIpiOGV4IASG7LQC8+JHJMDLSreR3tzm4VTSTMunSwjRThhQ4GY
Dc6iRhneO4NhQK/nRW1WUw8d6w4akAarK12OKe4xJpSfhy/NNZnNAgcxlXkZ8nzY
0sXLv5khO4z4XsaK77cKSaOT2V9rfp88h/H2pht5MmvKwmogu64GpO4/Z9t5TOrh
S7KYjpEfjOM47G5tuXDG/EqHkdVGrF1gdoL6KTTBgQcV3bSeHlv65luLwE7Abj+P
wKxD0CslFh5YuTORfW/pCyRKeK9nt1ADGI19mtgjJLDnLqq4CiMSQwX1KYlrSkfz
COySWIfz0IuORURCa7b4bzVzChjJmQl29MX7/K1pVVo63Ry/o5AxkbZm+72E9OnS
wLnYffCzBnkNZn0x1IxrYlZT6dLc8AwRniDZs8jnC9SJOjlBJRziXnljBmrptZg4
Z1RsXK5na6e49OF7oklyP1VW9mDhEoQ88YPiD7oztO9hIzrZ/RUAV/Z6lAfRup0m
UStslnocU24UNbwktw1sywFZX7dHhNqGeVP4caW2me/82E3f8kNxTyI+f9SSfxJC
JL8+0WygAJCijVaVgxSlWud0BCwyuIkrPxe2GRiKgNvE8KOUL6BcJBlfC6kHei5o
i1B4VtsSS31V3gzX5B5gVeOT0QM3x3P3eXOqlCRg9c38eTNco7jPg+putSOA13rM
84K+a2HifEt/anCU0d4WAvjSG9rKZHwGdrsgKrKODlFt+c4WK3Vduq+xpuyDkFpI
tDKopdF2eY3Cc3GTjqz6z56xsMlAIl8E5+Q1mvAxRQWVBa7gV3tWoFEoDanEmFzg
ImCKv5b7Cqr5Cgv0pqmFFv3WJCqQykLShmstCDh6rMfJevbu5uaZu6OWmhf1TL62
/HIuoQQzHOyqUfkLHK3RsZSwFFYnUAfIiNucQpD9uqAEP5fuTL5ZWR9bSPozQfWB
A1bCbTtkfof2BHtoY6ZMu0g/UFpKFXw+FinBYs3szb9tPx/aX4jiAm8nBaravAbN
dq4GKaYyb37evyMZ9i0C8QolqptFXvIHdYfv/Sw3KXMmJ87vobR1hhYbEM2SSv1X
ut2H+0FbmycXdEsuuAgakESH0n6Nf82C6WvvYpxZ1gx8j74Q0IDW/ceRtbDY2zcT
GLAcEu+6Ia9wcclTAXskf05YUsnRoZsfbpWXn/BG7AxBTYSPqnVgmFHYWTN6Waoq
ybMgl8vff+hRuxH1riMO3Qp3IYntWwlUm8RsYRq1sLlILrFTeKqgad/1gyoRlW13
hcJzCRJSdXRx2AKSa5hI+baVdi0DP3z10qAFYxQfogRuvfAAIZ9gGETAgsMaIq5k
RSa6BKlBXMj8qHVmzVWQeR/9MdLoOrizbDzNZda1x+qFFto/mUBPHVXIubxGl6EM
lRfw5bMmamyAxLembv5LH3+Wse4NrNkxO3xn2VtHIXnd4w6L8ixaH2JO4EgkFaTL
6o2wwIBfYe6Ga37o/mzn9f0Rvk4wEsiVHTc9RtbkkfZYezJIqiKja8pEm+cg+l9Z
qalfrplwdRDmOHA6EB0mZUNWFGxkriaGFCbfpOh77J5wiuz6riFuo3qGmFo5wqSh
+hpz6PnzfdQJ7jwyoMkL8CLNtQP2INLQQBbZ0Ug9ebNcwt1DhCCP5eMXbpxcYeBw
q2TibBBKB0vWWO9BcKk9Pm6IK1Bgvqsoyn9R3uenjGWVerHbw3zq2kjrf/5AXEFj
pH8MNbbEsrKqViWI56R41eCUKK5e810Q38qd9RPVFqPiLA5C2Tb6QfATHjZdQrza
NebAucdAD/eoX/DUqAoXgYfqDEYkip6LeZ6gDQ3pwD9M8CdmztUC6x2vb+zvUMGE
h2dclnxh0MHiktnsa48S7NA1EoUPBp5tE6AhHn9J6i+FKs1td41sdVKVOSBjxaCH
Em5BE718Pbkn7aFj9z+4XUnIsn1U2wmPyI+J5Or8FJOmVqBO7ZsC3R4p2DhO+o1T
iVCVyuKtZ3Kgi8/9muwZpcb+YNS/Cclq/qQ/gLThOBfowknne3qQZ8OIeKcIfltv
dAvXEtVvjKspUSQ5kfrDXwqQwI+7ihyqH2Vkch9KJilCUt4turEi017/O87I7ozi
h7QRqNqhXyhNHxBmRN5RmHXdcpKFtT2Kx2SCCGBc096daFgNIQKmoWOF4xBCZ7JB
/NB4aqCOQjRALdTF10FImfXLCPOXRwFvQGjX+Rrrxq+1YZF8D5XHhsA/N5qRym+w
WROzSI5IgSWtmxIKKgGnTTpGu1YGeInxZ6HTQKi3GId659eH5E6rNv7IO0S5GNEl
aHdu1i4kF9+t0mDJGZARv/Td1Dug6TOFgtIi5UPS+2N7TTJ8L9jOeJsJxvqVrtzm
eNYnTrqsMTTKYocb60w1y0bXiZYvI8EERPI9I7PxcLTm2BQGRgiIlw/MrsLGY5zC
2BtImPAVXNmaRTTnxaIrpOtP3xYn5TqcAfkWOx9tDPmvp+Ri8H/fVI1N6BKOlQKX
osIXvYPT3N1AZiJmadIesrAl0y/56uQfiZyPdZhVVWHWtiaL7QvrnnFdeMHG2NgW
VqvDjjMlmn7brmvHxqZbrVm7exgXHcHfijwtpWR0ZYZiztOrIq/76LMZ94RlI72D
arnwiv2nLuNp0Bxqwc6IQFS9YRNFT4yRQzumOOBTZp2/otO8SvxaAT+OWQWtpTlX
ywf76vxyzzc2TQWI9FlcEo2bnnbNaORYAqWbWIZypilAZ1SoYL3ePWzu1T3g20w9
TM0e/+XLF4JTZ3AnxdGXtR9q0PWmoh2czhcWxtG0tNc56yIbJUnQUspKaIufeSvo
9SICah76rBDStJaCPz8S9Nt/bp6mUez/0hSe+OnUeHuEcW/Mn82ryLi6NK9aNU0J
GRuKYNiIw6/yeKGK68gjISJw/9KHwZ+ThjW645SauIYo6Y6qdMusfzwnoi+C9JLv
8XzkCQ2QwSlUJPWSGYLWYd1BAOkmpDVW1X+XI+i5xT3UjAuGkpWrkUj1YmAz4ADF
UHe3WhRfUkIS4C2PtXU1uPC8XPhkL54g7YfuuPgbDFTy8KuqLUjpS/RpACRklbkQ
YvuIbZdCtZ1dlRblKTBWiYxsSv7/HymUG94n//vOhvtEZP/kt9dcX8xj0saxzYJ3
Cc0BHUuSzDXlQ/IqirYffb8h3P8L/VU+Y8fc5FF4oO7Rvh+HhD2B3c6yubzZjXy4
rWq2kYfX8pNW3ip07RJtTL2tEBrGgfuXBc0fMpvwBV9RUE+6cX+rIclSjEh8x6nl
1Qxv2xRJ7dpjrwgjPbHyNOW+UnQBxRAKvCLnWBgKSaqD9OseZeKLIiR6vu1O3rz4
81U/5PPBECTimdyS/lRkiTUkfx4Mizwrczmw8jmXhxCfu1BqhznnKpRymIekItFP
6jimpj00pju2p7Ip6zWqmrDkZqtTYj7MQvDAGTdFSUaaIHNrwPbdovYVNpfZQZ9s
omatnuSkR/UzdacAlzcAJAuc3L9nevAPyZCeaGYETgKk7MW5zrP172bP4bPi1ozy
Fz95y5zKePVG3oxDsRUSCWaWsKZjfVLEMjc64K3Km5/QPxthWf081/8iECtMQ0ZC
OSMNcqAlhUqOxksi0SoSTsNHsx5ZNIefDEn5fyD6F9tSgE5Y3xHdn2rh+nYLs9qS
vf8JPdoCmooy6oRW/Ti8n2pvi/07yjoOTJ8JhgjU10bOuOmlTBKvs8W2pR2GsisL
nrdZMwSL5ThtvhuMjrOQL9+9M8Qv3CClCWtO65QLHb/Ko1wnQ4J9th9BOThn2Pdw
JkkxB2OiIOPv0/qcgQn7v5SPT351K/iQI3erWxc0yN3s0+QEaDY19N4+QjR0eIEf
QkKjO+CmwCjK5tPTdXmZjEthZP75Z7DVTrBf79MOVgfJb0wZ7iEXdV9nv7DTlk6i
CBsiiAO0KvK9DipRt9z/C2tLYvoGcoy4rpeGPM4uGb6RNeYDPaTEjmsyK7GojI+r
amvmv0kKAIH+Sxg2BXKY0JAn673pQhTTX+ryni9bW8NZAk4+Qiatc0C0S81fqkuq
m+CkMrt2Ayf2X4WIWa4k1IiU62Su5IEZQaalLTKSMOMUOTLd9rfkbonrMgx9jyrx
Qe18JN1HcacvCXAo2Fq/V5mxr4L0GQLSBuWwjf0LXlQnZJ1bTiN/KTfYD9X1QX9h
UFJnVR8i67/hyMyj9IuybMPWemfDQAPSFNfPh9E3gQhWDFGZSKK1sKYLEPpjf7iG
IJNaWrxoE1Zl9TR87cpYwwS4jCpQfP0bvHVA0HMhXW6WZEfmKCS7nm+1XjS2a4VG
7whZyosh3w59iFjZDEiPW+LqYqFXjpnmnysbXCHIqn5TdHZgt9TCwrdE+rP/sJOL
emqpNeTdMr9Yt6iTrzj5AOUx3yX4wo4/o/bJDcyrRh841VIC5thn1IP6XqNHOVT9
f6LWcWEtteftxJNp5LXGt48IPh9kVGPe+dYJ+C/voMHBoIdEWfoUrj6D7rN2qIv5
TOkVWYBHyHqthnQu5g5ipdrFVSLeEAfYsxjaIMpMRQu9BC9n+2ZGQkys7w233rIs
Zf6Ik0i70PbLegDeBbCEzyLs74yuZN3Fb1cPEc4zzIEGcTAlE8utBksZFwrC6NM+
zw4FI+gmmamKgQ1a+2FR3zs3akcwYBiWioqDmnZfWss8Xcm15WtEYqT8DjCTiPAP
SKBlFA26q+F0Bsdl51ts9u2FgdbKkJ9qqFgj8/pFtrcOZTYtHL0OuQgseemq8yIi
74yxMIxrhP8XLBBOWfOHoA9amak5DbCnja1jOYNMZ2TewqGc5tQEzhStnQV9e3qg
4apIM/hTtNhhckYmYdufXaX7uTjfQuJPTLyu4OVRNkgnHaU9QtwnZUukGbY4QuJ0
UDyCF31FcdOXV7mHvaZ5WZfI9OuPX/nwsHC6ndgDF0irqXfMvh5FbuZyDjAQI8I9
MqXoKDM+0BphBsOUFwWo+2n/FPQUVUK3ZQdsscww9YE81lxHN3M5H3SUVbCxt/2N
GJK5+I4/IU6+neH/b5V9Em/EPucZUdW2aq4KAqBPKStpjTSKfokpsqtoRZeAH8wx
zH4dKKtYGu4Q2lyhpstLyf0KgGj2Jxd0OhCyLPI0tOm037eLNzkj1nQfkBevA+hi
HDZMTtVhmYsq/D/G56d1HujkhsZg/CLBejAYnEsngVD48s8HWrBNPHRU/PKsxOgw
bljcSkra97e3b9KF1y1oc0L815AgIRWjS1aZVQVfGpi/mJqG2dWLcEektulXR5FX
XiwpSRzmfLk/sasacemUXLRVbQFxs8qJW5JLsqJe7/3GpxWGOcUCoZZjERIK/dvC
WjG9zN0VCGiTGnwjV6YjiKc9NCfQCibmtqgcsEf9+yo00WxeZXZYgjDLps+ubm+1
Chwws7CjvgonYNaDpQ/ofVjeIODd3mtqNkXf3b49wLVqXyWF8U0IkFlYmL+Akszi
pTD3civ6parn4qNwbjLJSUb77YTJ9CB+8+MNEhJH0J5BoY+jockvaMObfAr4iVsX
q8XEpXoY/Ed3ycLV/v7wjlWonQgOXaa9J+8330LYF2ZVe3030EOLsI1u1x3pR7av
w4nBvh9fIoulz2aHWaEfqRn7UHYRxOA9cxov4yBfw5faIID7+/wQQ3gozpTrv77F
M8wMrdKnjnRVR1Kse6rtc2nN0hi6UqOJ29Po5B0J6NOPdEBuDJRBG3tV2r6rJ/UU
e/15uM6+WQrHXHZVWJctdPwVk+ueNFSCSZYOMTvIVjTP5O/p1xHNqbqDCjCtUR+3
4fv9jbNFpghi5dsa6v6XsRiYFcYPdsrqKlIFL9QRgQJsvOe3K6lKhbi+av3OxkH1
XyBiU9TChMIqkr3ZPtCz/80YVEqCHSH/M6a9H8WcR5s9qNf8DMgOVu5diJwqSqGS

//pragma protect end_data_block
//pragma protect digest_block
esReK4ITYx9K+PQnUyba+j81AQw=
//pragma protect end_digest_block
//pragma protect end_protected
