// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
J2MkBTDuDdfdXFAwtn80uQH6eDFFpLPfH/yEslgOPqTSqIiFA6q6h73u41LitHPI
sXgz2vs7LK7I99JdBJsw387S9GbIDbQUV/mF7EPPkTl9SaL+mIo63Xn4dLGHiZNW
Kyt0gdzZON6E2dGkMce5ahiYZESMdMqr4WeA7y5c5TM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 14832 )
`pragma protect data_block
pkFVeSbOLYS1+sDGsIfvoRmF2D3agtCjZNvuydFauD15sKw96UM/Gd2kZM9fYr1x
kYYuJxB4oOaItBiqir1RDYHTT67/yz/Cwg6P1HVHT/b3dlpx5+6rkSHNQX2ynaQX
8+MmhpunwPUZ8xaMtZ0nR8pSnvmlTNmT4F0Nhh4CCHw1pTq4xAs0YSqGXfoK35xM
TmH01dr6KZmPC8DclKJ95LH2zQ7ZfgxFWZ8l2FEdf8W6iMuCx4jYvPuHfv3WSdxr
GO4YcpBD7szT8X3N28GtM4d2RlQtN95ZVe84v3k0OlOq9RgizBbqN0m2pIWbmhH0
Mr/XVTYqL/Ad36WnzEa+en56SZuxEnQFO4lILpLX45UfL5xbOTcQwBgLHdVpSdnd
l2YMBX71zd3Z+BVgSftJu0p8R5vLtNB92cDFqanD2ElLxrkxHHxLhYN6/XHNuzRc
+EwbR2kFMv3tOQhaVq9vCu6Ra9MbNWVDZUlqSQG5xC7nqCwvxjonlXw7hr4YqVhu
Y5zIcwogI7Umbr7yxAxg1JhYFi/WKWO4yOiKFxZywLVj9RpxphvyuPKiRMjhN8rR
a24Q8iViIiNRxA17OMWPedMi1Gf3mX7XeEOKB1YvVR4dVRkEJANehKHA88maQuM0
B/AIEbnsisjO1T0ojHHl0FJF6lRChHlMjRpGZZiTz7fKvM9JlIYSG7lW0EvKfxtI
cpg5FTy2Ocz91ehPTdeJaYF/uQMo8Pnfybz1tMiKdIMBLakjLEDS5CEDyM5E5Qkc
3//FTf1CRkse+ZjCHRcrUP/cOq7lgrbasLXR/F4EMR8ss5CS80J4S/DLI7W2BoK5
1aADOLW1kEVztsZFfHwak4obD4OjhH5MCzsqKruBkJbG1+o02Oop7jIfWcCBMxLz
Od5eMNgotfr910hH7UMyWzwQsdZiRVl9+QQmAjR+DiiX1ZdjLAf/yKFXZFus19X7
SuFDm2x4/qz+d+eTOG6h3gf9f+4dPe4bPa9a9eYe9khqqWY2UqYVIuDDvMNSt+Q2
1tT3NTa7f0hfutpASANc7WTjRrCIUC6KY0Vhb8EudopqtnICqdR35LRQvqcIaUgr
DwBnOt63w/rO98agN/T+Opo2T+givSsFVZ0Xh9xYGPWT6RbVxe0qBBpo8tlSdWAr
QOuA6iaJ5MtvmC0JRF+O1XkZnHEsjWzApz+nkseFy/A3D6+l7j057thl7o5bvR9+
wToNxUv7K+iXihoCTm7X6Q4OrmrGsIcU/eYZlX6Ou7+Vv1TGDeP4QPzEzgffuBU3
ADNcZ/vP4FyrCS7F1kIVFvLstE6byG2TyZX6QHy4GLFKWGmqzs7BomRTBqwhRfqs
LS2ynKPoK0xk0l2z4frcIyt8KbvGNNTTP/EI6DtotHqGtU8+udnpb+tamectRaHj
B56hfy7hpBpviNE+BhkqXXqDfICiDQKtDgS4KOOJBKSnVVQj31HREUc719vZd4jl
rh3OXuLoBtFosvahbo0FmSvoxEB0PX8W/D1MPhSwCQfoD78e/jM6OMczSfif7mza
Ywc7u16M0h06yS85d8OVFsrokUbOddubEEMipxu6fh8zIbAsJ0FslWZNkl1KWMYk
8aOpSKkkdobarlsjji7DWfQkn79NGIh4HruhtkehdjTRkMDJn/cma38pDHXyFbIr
gNYjl5acFWPdfLEGp5dyD0YxXDJcbGYNY9Lpm1Mhu+5xmETRMcupXnszbX4Z171E
rQeADs0T5Bmrwn0g4LRmlMqE5mdrI4mfknYpy3I3EMvZhWrm3V6ikNpP34PwBvoy
/0XUJI6mcg02cTuckc+KxPvGSZxD/ubXdVp/krMk87b3lYcCmPHocStBxzEIWtbB
rf8ZW/nZwIk7alkNn2K/zxhkOEbL+twNVB8LOxdoS2n4aLgQPOlCEefZFK01Cht/
b57219jEM9tNwuKI/s5mHxvJNWBavXWxDVc/rzM8KuMFZeprIBhAJi5XPPctvFno
M8uyhQ2axZK2KY3/KIo4pdwoNeFTM/mbcXVr/oGk+Q0qUwac5i0dl6hNGwpVGqN/
C1xhmyaMiX2h0Tsut8u5/EwrMmwwMogUYOqnOPkSP2SL2sDeN/5nhBEMy4Bj8FNa
3sPZnCjTBtJJHZt9YMHcA99OrTkivumqlWLf2HWq12b2L3pfOzrsOLOBhltYZ1Zi
V9uLP7rl9ypsLaB/EsGlF0KkKEgDqAWI8tLoG+b4VuZETY8oxh2pM07L/al7O0cB
KeoLlwO48VM1FBaSkYgkHEThZMS2GN30sJ+RfEPcZNo6w8RD++HjAIylRVSg+G6m
HUP+xsDG/zmxMpznksCyYLGG6DC/YGeZhpXhxw6V6SnzbbmvKsDkuBDi6DGKKA6B
/c+NyYi3PYvVyPTfQDn/4FlyXVK/z4BgduWl5nyINZtonh1vdzJYHEUVyzccApXG
Ph6ywItsXlGA0vyKF7nPSnqDE1uL8MX5MRkcXvksjp9Rh9MU/0YYYJesakypzHdl
Y7EP02gqqLQisg/b0XLoSvWWYkJ7yaWLh3bRHI1OYnxmdfw6/gDLmjt85LlV+5/u
I82pu/UVK5b1rNdMQWxmTMKtVGrlqpObB8JYmLufpkBKl59HDulIQLBYHJjeUrC7
cb3OjKVyVqq4jyTkmCzaJihXwWqNXVkpTm588ZdVcfjzCNd7qtW+oi3+jmYhItER
nES6cEutkXLtnii9btUI0xfoxLv9MFV+c039igW2Q8E7BucIkNJv4ZMEqYdYYHpy
TBnlcvnIt51JrN/eiDwadErgn8Vz51X4oIaLxIR3u+oQ5Vk38c4B3JsFcelkR65T
mXDE0cnRVSh1FDNtz7a0PJBiYvDfTnjj8TBprylGQCtDKLVqyMbUPVIuYi+j+LXp
RE7W97Kbs/MS1yezpdoMvK0EW7sMdrgZIPFEH0JrBoLvZ7GgiQj6bMucPVfhGgIO
XbFYzWmPd6epOGaDKW3asqlSK6UYbKXvBmNxbzVyGh0twag65OvHMH3eOmJWRoVj
4FU3O/svyR4qsiBzvaIOrO5ljZa3F5qP0Fsx1qVUskom6W8uWzIPbw4WZpeeccTM
TX2jYBH3ghC57MtLGc6XDCG6Zvo8t6nme30E8Tpxjg/s+RVpZvf565ulLUKtAHju
EGC+Q27041RGK3QpYjFZgqr8bHE15XEeW1qzxqepOixPYznf7lW5yS9dV04+MmNN
q3izkor8waRouK6wkGu+peR4fUiErqsTD1UVPoUtxYqk5VRId3dwhWEvgpTCfZF0
t8YaZZIhcyePQJe/WujNH9uVYfSdcOMm6WyA3LGXO/sTqmgi7W1/M/8UxWAfrOMG
P+SE5HHHQKQLKCKwM8T4JoU/1CkbPw1pFQZsAOWBVRJSu9rYRDl/fwnuAH5JZLub
Ylx3VGQlnMIjZffFDQEIQTMxkP3QIrrGYojNzCIxqOFrQ1fOQl4pLZa+jSGvsOkE
TengzxV2i9W31eslj9R+UVY6Az6ynwAnrTa7XJdjrMywsgzeTMWZD3vKpkzE2yvH
JFdaqeE6uGxN2HneJvch08XT2hqL8utI2ZrD1qwvqsAfRaJ9iqDzdRYrRuwvlBtp
Y6YpARKeaDYt6LLLBcrL14/iLXvhUmk2j0xk5p3gfjZiBdZdAK7ahEUbifmSwjh8
yYj+4wr3N4KGu1A7LCqp2woBhSUpL2XsL7REF7xTPW77YVcUN7IsPfwzpPdZlnKw
TMUUF5y1hUXZ5uHO4Xd1DL75V8rxBtE3CUrAYa+e1qlVTmDCBHffY4nUpWATHNTY
twKe7oEj8FNU006RnnddvdvJO6Xl8X1txVFuKUGhkESYp6M4i7cdutI1ooyiDtd7
uUTczaoufvrtMQsUrfJ3cFuqp2r0HjkX0dmrgBRPt5zl0Nk6QRlizduV5tyAx4QR
666dY180Bbm5kQIw8c8nR3njZsAFC2/3tOyUgbUZXFa4Wu4rqhx2u65nAbS9h6Xm
KETN0V160BZ8EZPGX8Rbd1NjLBAouPA1sanGZQrTrN6YvOq5rpgcRMj5k7Ss9iZb
53Qc4DS3MNePJ9MVwQt0MLGeQoTCyOWo9N4vQrGo4HEjA5g56a5xrL1I4dqwFCkV
aq3Z8uHRhY1tNIYLTl62+t4AzzeY5sJ2CiMipn61nj9wD0SqMcmDaUTceffy/pET
7t4BTVNCPC4OZr6BpB9t+JLsWfXj8iAoDLGkpRN+NTnfZtiNFLWehG+UNjIWSZOC
CtIw1050Xe8W6KFz/mO8A1D5xurKg183l8dTSVDWj16o0PuVUos3LeuOVDwEedhb
hHUe9XHAgzFhGUl89m6RuR4v3PFd91/vF0AMyuNwPLjvn3bOsI+MHLAxVXWln2ry
DrNHLY+IiM7Dw/mFtYIJUDWHpAgbv8aiminbQc5ekbb//9x5ke1PnjINsx8cnUCP
IhKRmEUEtw3bNxWSNKx5eFIjDhMi4TmDx8+i2jjiMf9i1CF3u1pz2cRobMYnoLRu
ovmLsS9i1RNj6OFge6lPPsraERlbQymuxeysXnOX7EAPEqo9zQfWG8BFdreBy/VB
eIEw/qToAxhu5lAHr3QS/BsObH67fSrBV3yOeuAeVM0yERCchswhXV5CqWaNBOBW
2qtOCXOkmOA+XMcwrPuB4ykF6TZB4Tn0N4IWBL1jbDo4bTWK0RPh+SwQbcTg9SKt
7izAD0zS+CQD5pUDP7geVWlgkfEKr+A7n3AHuPJ44k8qiEwCkZTccXuVCmKEOJaS
n1ATG6xhd2OBQuALVSMgeNOSR6jZm2pw+elRZd3s86UcTwiGfyL9gI6P6IoDNBXQ
DP7YNgRysogrHc3zunk1cdeTW/oarmkHs8tgFlDcbgwBewJDioADtJ1S949Llts7
MlJRgzoXvpRqi5C2BN2p3XTXyFya1OJTVI3jSUS6heCcZuNL2o8iaVVw011QQenD
JaqgWFiStXq2ahJWGwADkvjFCaUWRWLjQlo0vO+Fl0aa92x/IM/42Zr90VR/zxs6
w/ZlEwdfGNY/NsTt6RGetQkluRs4YaAaYDosdVVEL+bIDf/V+HIu7uhtU88S+Hvb
ENXEsltfbJaFEx43LOiLX0aib/NC2pDo0QwYQNU8S14W6BGwYJsLlpvlUWxgfvnU
tZ37axARfSrhzK92EqBCk6VUYbFqVuAtB3LrV/P93OZhncx4nrnn404IqcuBpHIo
wDlOJBpuZLwEYqrrftYkhlSKSIsAcALDGquNLV8UbAmbRNt9ho4dXW50+iVAIM/7
a4MfLaU/5iKGb0fDb1fTPVYJIw/FxgIkwRrSuXdKufp0qmYMh0PxbPJ/K6ZoR4EC
ySBcfCytW4HmVFNZYKrEs4IdmbnzIpDaovXc23Ca81Cthc0STJ9c4CCVa3RLHyr/
iDrUdrnxBB+QQJiNqbt+dCv8nzgMIVPAA1rsZirBKVxHTYrMr1U6M9ncf3fZi2MN
13EMOCxqZ3+rbtGk20PS62SrXdXRw1+cJhLsggFDO6ux1gkns9RnPPMuZjVf42o6
LwULb4XUZkxYXd/EN1fOyWkRp1b6dnoEpffafSu6yw2EaJlFsnNMTkFz4OfyfykW
YV2iOxpL37TSRK8CpTRrZHEYXnj5T94Ad3tdWC7Bb84gUMvtfK4MApKjjYsW1ORe
KCASGM8e6zf64AzkqTRKvlvIKRIe0/Mg64uzXMhVFzLNoDoSRU85Um/1d7EhnpYC
Tw5S7uUr8PpiK6Vk6rKw69xMz4gMPxMliq9Ps7N6ciHW4xm9RddmeaA53ymtpIEc
jkEtLm5/qC6OWSxbfnWo0mK2Ae6UIpLQ0klhBPKIz2nCcM3Jmr6MFcTBgxaFz49A
c8WZ/WfdABLjnoBQqBiGyZLkMY3hX7gNgf+4fObfBPZJy7IMCJphNWjd8fGhXnr/
75ATaW5h6lnDNPXG7FSvSELNg/cG7jKbLu0FCqMNp+MdVtVF/XgulrSa5DIE3KBI
nWSLjLkZC5696M7pM4LR0oVdVaNRBFgRIzsmSyorPzJdyaXB9yc2XbCqQ8lkmMMd
AtbMB31Lgy2EvnK+OIodbFcDSeIS6SM3bjenWhY6nXrAZ5viMvYSEqjyctLzOX4i
5vX7JzHHBCAd9IHfSFXRjEf3TkdWBu8om0Z/0iGiEAs7M48XIUB/xtvQPW0Yk6dX
gG7VbUPVBqdg4kuXQuT5E8LY0CUrMWebpJHA1IfyYmek2oqosz1ZpV4zPPx/QpVr
+I/4b1f7FVaWx7Ip5jxpclc942x3MXi9JBE8q5Wjc78TIL6zqdPUKVX6mqlF/gqj
dV77vsw5HbD1zLFDFbLV4vWPgIwi620Izao8BHUaanS30m/l9w1jcYIWP/XSXT67
zra7nGQs1BGA+CmryqGilIP/7c2qH8OsKsCKRZGx368551p4Kg1qa/gUwaAISRKQ
VS31zNPYB2AkJQbgCcTncczQriDxWKkqWGk9rkW5C+ZBzyDK3GegfWgaf0VJzVdc
oYjzGqgizl9zutAKt+BiFRlo/FxpD/z4+C4Ds+CLZ9OTqd7a9pr98iKyn3kFCT1y
IEVp4/DfnPLNSEDyfaMdyKnDOs5DTF98f3mulZRbPwTtStqYmWD14m8L9D/wrUpL
IGShFf2ZGPqgO3rcwhOBeEMWIQDcY5EdWzPeMGa9LLL2HPL7RLczHNBnEaEPL6i0
ehlYg37nDPFBxJpWJbVAtug2hclh7EEwWGIyKLA8m+sSh9tCGGd/+BNwoDY0vzSV
JuZuMWUhFGLjGSpGi8CNPlDd9OFmoJsUDD1KxXlMD/HFmz4XNr/FiFSqEjssupmC
nrUyX6hjLHorkBv5OKy/5xJvAWmmNrSzj5uJgLIQ4EljeYVQAcyH9Uzp4MitQyZ9
XdMLuGNpXud7FBFjAdKr/NW2nqpozFZgHAlG40gFLnntiPf/adNEtxaZymSFYBBY
25MZoK4ATuaEiNcRulZJ5ZOpho+05vwnOiw6TuJ0H2IpoK2Uz9F3LhLI4yyh9f7M
sETo9VPZ4Xlu9IImp3ukLXNnq7L10kd9E2cko1Oc7f2XjwBqwDvgKPUPtI9N+2ki
jOxJYBeF3X2dP10IiWPxU+n1dpiI4AoJZGShNbLc5/MXr/rxI9J7nJIFLyAORius
d+cQP82hs2jah3TQxFDU6ly0GK+Pl0UIBS77FY/YZm62E7chWDglA/xiuCgmNL3u
W2EY2+o0o5qGiHgfP1U1tbC9k3e09a5qF9+m6mI3Ii86UC5g3ZIQItdCjuUIPBh4
5+iSDwIyF8hAK2eYSLFDdc20kZ9nlPl5QjHTcCBZ/jnbdh8rxMimWTqXk++4p1uk
rnd0CtTSw6OP/380AiVaZEQV4K4n5fqQJmuBpoB6fC1h17kpu51yUHSMWnzEEWgB
3I+WRqslu3dg46OhStJb0/bsxc1X4arxevqJLAjQIB59Wf6iKHYOq1vqPQ92qzzb
JjqRexQPQNwvQw8mmpajq8ImCWCQFlJCVy5jVDCKsoW6usU/UvS69pScg7OzxDmK
0eYxVoSeda8hbTX4hd0BbCgvKXxYkKC8dRjt0CG0H56+qMfWnOz8NhAtikecZPWx
yg1KZLn7wzyJoYFgFiTAgprbQZ3x0CnSgOSRHOl5f6eLZBakpyafNw/dyb4gdoYg
ucihME+hNKum5qnpx5RbEtRktWTXepcU73obmDu/RoxPpSJHsPX/FoerF8cNVUvu
HxbNfDibRhVo6Uk3v7L7ohqsR2ySNotRWBYnCy3YiPCH7pX1h0NC2LSGKXdoibBo
kq/c+7/S78aVcYKKKxPgGZpoTkJCaN9euszVtI4jsjVMUQ6V+U5yoLy1HCMBrGVL
gZVoVMHmdIGl2JjPtC+MK1gKToiI599yQnVJuGmclQqEhSV6UgTpqo79kKHQDWi+
d/tn58LNRiANg6DDb5qFACIn9CO/dsD+0JKw0CusNVukljuyTuvaXyndmsVoBKWS
E1A0UAPxk0oSIS6pYOlQyvH6DPWmQj4xT7sxQEvqg7zhJkeLKUYE0ErAjYAa1Bn8
C6XBuCJSMi38kNs1+qnd3OThvwbU90KuZk5DzgjgQBtBHBhVnjYZovoVL7TkM+Mn
wGu7MvbJvepylT8zD3vV1o5Y7mibkLIYzII5lGdi6zouXjOTkm9GQy3WbeVLbhzb
1QEPID6swnZeFYaQcHLeudouo4Zz8MH9DcoWW9ZdzS/86feM5mUed/yxh7lNCUIR
aYGIdmZCfSa2+SyMYGdqIMBsqR7aZKINiDyT1q5zBNcOH+frnox4lxMhdGKsaBT9
AEsRHhQFSdcbYWwvEaxL5VBtf4R6dEjdGHYPIwrNcWa1IYnFGgHHhnfFcb3EMUGy
CQw8AlkmSssylMpiHhbl/0pa8DZ0PRHLKvVJgIS7T+88RQh0OKwgmP088EkVKuUY
PkpMmc5KfRqHjZMKNie17DJUCGPUjUHbEt7IvcLXM6fJoLZWWVuJq94x8vStFGO8
5/KM7KYGD59iaRE4ZdYrjxGwHPf7yyFkKDEEvUqln7T+Vn4BhQ4+jD2azKvXy7UM
VYZhsW+ZTmG5b7uKcQ2UKHsOogg8oq7flpARfRIQGatLU93pBzOHH4jB3DXOdVu6
N+RFXrVh7kqw162Sed5I+Xx3nagmFPXvMzpyJBoyzjuAbDvDW6xs1Yqm+TBYdlLk
WZT0eoKxhavSc2LuqiNOdtPiMfPi+xc9eBRoKIeZ7Vs7S48RkzJ6zhWRWe1RN0gg
/m9t7Pu2bwCeXoSL5BimrqMfsOVDBCIYHzs6HuL/xXybEYst9gx9MY54zN0U6Yj8
UjNVU1KBVEBSx4y89RZCFlUkF2Uji3iHfNug+Slmt7Pft7a3D+kCE823E8XDM2pg
8eEP+ekyfRFNVqQ73tKsE249CQUUwjBIUuKVMSwS56dRTeY72A63MxRfU4w6wJP4
Lt5F4llvWZzmJ0iohtvKAwUeN7lrzkg+FuUXGZbrOL3ATliZlYXjLQdylg+eDTP3
t3R8HFs2yjIYrr698Mezxuopq6N43igsQWk6aT3JB2c+vd88T5p2O5OzZ7Nm9mH2
n0kS7Asw3JxSM6GRJ6pE2ucGoC3j1RLaNB1tBMxcJXYx+i+fRcYHCVJjH1+zYV8w
pHq6dUZ3o4I7qnMANAXnj6WpVt3IP85jxTRwv5Jrn7r9HwvArEgdqkwVW4laC+an
z9WI8p0cZRcjx80m8bSRr/4MVCHQtklP/5FNZSZ8YEUdbK8ATFeeXxXQOvBn4vs0
Qf0+z3AeFbLO3E3BkbLcgdcfRBAUAZMX3r4Su7wICpj4sajQBOLTvFlqKfPKTm22
f/bwdCnqS6/iiQsSWCi//ZHZVmc3xdhrbVysOJ5NWMFdQaYvMq8UKmNAdUv7nGTq
X30NqtacVCF7AzoBF97lSqC8Wke/VnitIOCbY+ls2cKbzzFWST5kemm+YzCqrbcf
l+P09pvcy710gGx/3jZ5U80NVfzwSzBXlh4zg3qDS+by0z32B3GhsDQP0qDewJ6H
TvASCVJVgQKPBeXNO4dxu00+aEqyGnG5wUCqbYrKyY1kpwzOoG5IiD/r6dFaUkwJ
HcUxAyrUlqoCfdD9Z2tXh+ZAaVCrtBggpBaXFHjttAYLvo8w7gYkTlVKz79FLBsv
py4wYxQaXXn2iw5NE8H7qeisDiRRfEobYzqAFcySrYpb2S94MFbg99sI5oToJnHO
5SJ6jUp07+Xa1VkE2LFdzOH0UmPJB9nbla4gfZg2WOVJQco/Jl9OKhUOp0mlfTXn
0oYD3rDfgYkSYu3uYHW+BMAOmD3Plqrch9RktSFV6Hd/8PWjSInQ6kdcvYc7rv+Q
eEDIqWhW5hXhjXSxoeOo9pwYfVMNiSoQCwxszsZCZnIOYt/wXUOo70CVVu2PBwEk
wrah7LtdIaq/E/iOliOGA6sP0To6K/RpCwUNl4vpCzkETFII18cyY5uX1wuf5SsD
akLSVf1CE0fHzcDdeX23h0XJZe9Ay3QNPb696fHR6ChRST0knRR8KyNMGVyhlTtE
LVgQeOwaf0wzZJofGZ5wRvpuuVlcP0yDpNlDtoc3Z5KAlEQ0rsh1uVQESvVMagXJ
p0wT/tWWXSecd1IFNAzK5dqxkF1kgbVQJvw2eHpkoxROPhlE5YgMQB/Ge8SE/uT/
bHGoM3iBDKWDSI82EzH2cn2Qf92Eo6o11FvH2B6WImq6l65G5HH0uZhY6Kbmh4cU
Trny2ArpcH//hoQPcN6qgtAhtwC7hVjTHZwZ9PpKVPX8sGMnh/Na1Wmtr1pifue4
oVuF3wdi19hXeaxjhnvvNYsFsToUVWlJcA1+jjUC5lIDYwVqLh1EvRC0UGosjjOk
0yoZay6tGoXl6z9PILL8bN7RdbaGS5KSSGdkGHnLAkxCKbsLfOiHQ2kjzoqPGk1T
ucO8ygb8pObAajUQAXAaYccJvT1E8JSL//tp+mRT02Kp6ROTDpHz8mwK6vSL4eEz
/ebnQpiPeYAeidWbbjkg4bJ4ldRMBNTNL49rXGjV/BUJg9e0HyUxOvYv1mqek/3P
4WA9w4HunTN/f6nHBvwopS6e8hrB5QuBMAw8xjMqb3//E9TJE71xR+m5kLzl1Quy
ysPK1r+Q1AKGwyIFGWCpsfyRQXVo+vIOW2Ko8DTnnYFl64fC0YCk9dIgIuMehXR5
Tz3U+b8jWYYoCA0rBfRtgkhSUIPenEv8gneEFY5XSRhnsY+aExUI7hPd2owRabYt
b5QQEMaGcOATP4/F4bMfad2shjJvReTvpLfFNC5LgMdt+j0QBXxf/2y4F8T6nyne
Px1Tuo6Yx6hezT7MZHZ8C1uQNbfEegM5CmBzbjys0mLRNFk35ti5QCaChsc/2RiV
sBgRZd5v+7r/jkBWqpQ50FBBqkSFGZMRA+BKxRltfTvYQZaH9tLKnVtt29bSOl3z
W89A2yfQ5GE0na2XNzjHLkxmBNvPyB5bHF2KxcrRg1V+YOWrUQ2SLtqTIgE9zfS4
NtLpQLte7Aulj+zYB1VAPA1UhLZUPrKRavAvDX1Jd02xRiBUSPSmfOqXT2Q7pbD8
obUpZL6onCFn+zbfhJYUh1HwjAICfjavrgZbLeeUs0GDbcA+LYNsv+8ZniOjgXaM
lX7Lw0uh8isKgUwlHZUv/rNG5c8QzdDufwDV7j96HNWeME5XFFcqXivPK5XwBgak
diPPsteBcTY9NK+Y5pLwDHLuDhRBOlD0uY147FOYLfB60mQcF5tUS2epcwELTCmA
m/oPzfJrWpQ28PWswW5ICCY59m7qTQnDKSlcvaKDFR9k/1Hcd3DvN+ynZUpnKv2y
hryAPFIDDs4dD/b5K2DQa/lZNxJnMKM0Vi8OnQxBQ0Md7r1aotUP41AggTZ7YOyV
0C2qXCjyEgKjfrNtW8wcltWPwVv4pTDFCU5zL47Fas07WHjmBND8fVmf3fbGGcy8
Cd0sj5Ie/+7lXDpqFrLNsSVw1moyxpLWP59ahGrnS7ZSZzbGPEucw8g0Lm7g2EEp
mI9bHoROCcTbn8zAdJ8bwiYxYQN1zCwes3S1nhZGtCipb83xSY7K7RMRq+f/21c4
6ZygsnacT8XXkRYM7aRHGqUniwzUf51OrzF2Chn0wiCD3c6iuELL3AFcrZK+81ck
LWNl2AIz3v0Mkve16NXFUqRgFlMBuq+iTd7jGLi/q6Coj5jhi5vIG9RUhCUw2XDz
wUkonBDqab14eJFC1n/2P4ipEEeMPnIlZ2TfmZfOMgGRp05y9B0y403zAcUREvTq
rhcSWx7oJfSo6KMTXEF6FGIYPAHpldx+h29BXbZpGDS0nof0bld884ETLLijrXW9
s9n4CwqI7DMjOlBDokUPp33/ANje2kkPVWT9X2IJktCT3i2qpc/KsxYwZ5lKPKwP
cxlmGAAZsBPtwcGmG7pzB4SjAXNeZcO0tUnecQC7rjihYSamB3B2See7oEjgo+P+
hou3NFmkLUk0ZbDQV8jyf8lEOZv6RSYz4Cvof0kyBB5smFua3vKaNOI1CY3B+RPL
eiccdo8d8GF6G87xvh7IQMFihq8VEAE6LroyF55XlQWFOI6BCgdgKIagXoWsIvxg
rQxBtPrkNdlj5yFRHgWYz9qNDZR+GRIT+BFbdFT/wQlfQl1qO3JlzAYBW5rr7yJo
gk25iIx648551cxOrFRU2M0XeI3vJ3QRGP8h5AXrAOtBfDLyTlR9FUJIguLP6AC0
3Jmr3rgaCO/MLGzHtQy3oWnTF968vTq+XG9Kv9Z8PKMxIroRIUKpNgBXHXjrtvdV
dFAmkBbUZwAONqg8nAW51SzMz340OtlS8mZJyiZH+jvGCf7vCo2CeoG6unBbiRkt
yr1TAG8NBmc5IIIGL5zlNN2VoWcPfaB4mvRF/SuZcb77GYKmhdnBKvUmWPm0EiwL
ZvdHvKs2FV5OeD8jkT4z7ons/udg1775O1BRS6niDXhJaZzTnee5bC2nH9CWBsH9
qioASBYYzT7s2B3IJmSwyCVZFKDugDLPYO/pRtsbL6hf+48HgcVYXfWUN76cxX6b
NYdFWa6isi+TuQMomu62eP8ZxNXA3SzqUv60LV8cvlpIEPH1dDcyL5Ra06tMCSjb
I0Z1/PUit9APdwajIpMdsOL+ab5WX27H67DbKgp+uHym6YocWPq6D2+agYue1QeY
jVLaiXEqyd0z5HiIuU2TB3mpZwa8h6SqWuHPa2VQ5DwhKi7j9V7akPIeXGz4/FE5
+HbKl8z4pLS0RTW6nPyV6U2V4zOnK53r2MrmYS8HRlcm5zIZA0FYu8G6YnrhQAi+
nLZF0T43EXtzcXNxhl3GtRHgtydELLy1TaiLt/rYlUwMMKfuZ20I0JMd/jXyjGnj
72+pJe6gJPFLDeFHRmns1aikpr7kly4ZP0oTtxeRCLt0vlIUu2H7FyVR2gErtFNe
0xJbFrb8sxA9/7Oo/P7f+BxGfpKZ/ylGeUwpgsibN7MxylJdGtcuz9zgvfny985I
Jb1gqsuBX8QCAkmebojgFoqi6wJePc6tETSTMwmousZFWXLfsSejhUXbKXSOxblr
xG5JnVs6acvGY3ZUHI+NbSri2wFDlzsC3WC3IYb8ZOWjfDfl627gMdASETXXLWHk
eWiIcdAvhMsL3C0YRnyHb7KoYywUMVuJDTbHn5JPIfOOECHzKUy1PtHTzIgV/dn0
zohZ9udJrLR/+63yhqAjpEXCN9rWWLEXu2nMu1qS4B7iT26S2F9m9LVdMVnzgNTa
AeyewMCvjnsGGZLocSrbgE03z/ZYQ6FOtZB88/tt6WTQyoGVcQrJNBvf0e5O+EI3
r7EXoZYE7yvLyDKYDsqyzKpHehIFiDTTclODrKPU6f9ahv9Bt38Dg20/b0rRoO2Z
/nHw8sLzMK1kGNlEQ05vgQFiqNXKoQZ4c88Bf+k2I2OwWFT9nSm0Li9fJOTpuqex
f006W9Rf1hbWom9YG7QQZQF2h0i4GHBFrB6smQBzHdRhaeAL8asoS1khUKnFXEdY
Qcvsghu+kpwBYPLmk0YI3bglbBu2gZ76rfOZWGFrtwNFQpbWOKynq1oAFNlM4tA0
H7mWps3TVzCleL5yXppHkMvJc7uW7j/hckDnSSoX0yiQmDaYNNYBBDFtFoeN6Fkl
LErLePNauNettff59V5b8C8rZ3FxtJyIbfNf5BG5AezUacIf0TwJNE7DahRjV6MC
rEoieYKdKWDP4Voazua7p9QNtNl6R9eyLPeWpEqluOzbkz36InDLbWVy/QJTiFTx
alNsLpfjrHOC2YYcJaGHek8UxurwEgQkyg1Z0Zor8M2QLm3pm5+VhVYwH8PS6m1Z
2SX3xsUE+iwgwhbwW+SchYhgbyiq1nSoWFPAHm8EpBiHA0gq6O/8PcXEGrxtesMm
XZi4Wtd0hF95PKJU9eD3EhZiyxwVQNLShPGCgJ7m/HMsQZPl0SFFfoVtFKhTvH68
W/M1lk6p2ovnwAVHURcho9hC1dLJsLGQNZ3GKsGYkEWLahBvKo9ef8RsRcK/xpxT
YLz/Iqfc/yKgjtwv7+38AQ6kuGQZKw2l55wDFLCcVwfnEQcjFlOA+C19EGzM7Pc8
E8AHaNgUzuNaW3hf6GErSDdKboL+bx+hX2+X38JIsKdIhfznzzw9hNN5e3PRBT5l
WY9KFs6q7ZWWzS4ECKQOm7VBEEa9nbWnWk2TylATmYXXYXNV3Dbd8NtSkxanWTCG
18cQ64n6ZQ/V40YqkznmjDDvjgao/l/oMWMcIR7b01vau3Y2CyM2RzhTNR7jWYfz
6AnyNk7xo6yC/FneVm1iwyJLn1hIBeTQev8kTZa7q0M1FncKx5t4E6F7vTU0GHXe
YXLEJ3oRR7tL6qv3IaICYeukb2Th+plPDFmXxAehjRyGvrRJQslsywMPacRD1gT1
a1yLGPvCrV6/BTEVWn/IpAv8cQ+zJWNfrk3805Ss1NYe2gZC0lDyI43RyV6G1+bA
Qo3QOb9Z7N9EswFb8nss35I2z9nXlO9m8cqK79ueZm6DdYWqH51jAACNKRv/tdZr
+k7Gebc2RaDk0K3rm1DEeMAGUw2RpygWbQUwCfoY1L7C11cvDcceU1S/d9cB2mc+
VXugRWnT5/q8YC+Xldnf4Crh5NO1lOBaJtWXqua0Z58B59s405LyijJAm+8NRKP9
vedyAvJlU/p7zY3W2m8qPkI8JRKl5W5aciFFkX1487PHDcqw7o+IuixHUEmXJ0jN
Uj3nZqgZsrzHK43vvA3pukUjU9Kn2SZjjZMoW5lYf+dZukc87baH/Ey0Dsmvn3vE
yAe1/W5Jm7+2tI54l65eN9EhYA1+WYMU5yi30iBXSnttMZRNJpJmbDvbb2YEMhhp
qhIKpOCKZd8HiZ+XmL1verEGru43mRTkXypqiFcfP/945mv6is6tsM1Ol+STYVYU
eTAxYU76oSRqFyNxBYF9E2hwfFDC9/FvIKFDOETvGWrdcme1NybyzJ+D6LE2QhaM
HcJq10fVVDTkmMIHMJgXAHbGA3Nswjfk+qFZgRZedxj8063LhwDmO2ayFkz/RW17
euiV++lOCrNWtUk6574Xd/5db3Bhn2xwSmyILrQEffDHoSEJD9acDMwUkaeieRNE
ET7vKdSvY6y/aLqJf/TGnzzs4Guca68Wvwt8nSRWUTlUYcHWqg22jiwxBA9mQOw2
3kesDkCOX0OMe1/MZt9GQ54jvUs0lq7MOciM25XM5RshyrkfNNiRMVsBQALWL6Ne
JUq27CXrCWry0osVtfQwmcMkHqsGm1n0CkHj8gzCx7DG50n4mKgtrynkoR+OFa0v
SCs7/4HkmV02Evc9LFMBglnYvu+at+qXo2qaE2n4VMSRO52sIZEkKLKyThd/tizo
xlXNE152xMfuRIe9qNpZiic8Oh7JlKp2LHKkrxA4sRSU3X9XGbP90osAK1lTOTaK
5xPMMTRlFIRR4C1ZZL4lxGdgzRg3uDUCIadP9AGbq0iEMzaC73a9xSaGyG2LyXzb
UE1syyV2nWTy2k992CndOUAzRSQf/it8kALvbhIBRChcbFCxHDEBtjCB/kVguyEH
kOBLLumw4D5J7kYIqeVXjwQdrjFkTW4lilhonOGyZxqQV+0nuEONVuYC4frBHx1t
gBZewV/zeArlD82ib/94phJXYQw5xOQHFU08flEGmhF1BOxxGItFL1CpGkwMCuj6
kKMTFcrTT91NpNuAjiWKjxOt+PcdhFSjTOhTHJJPvsGdwauLFTDW0X4nvYUI8GV1
fC48Ecu/dm294x3p8IwcE37K+34fknFHH0BrccE1nXold9B3ltBFxsEbqN1gETUi
p0ycO6SuvoCSO5pJpFHveXnkGa3KaSBOszBIpDE7EmSR+DIqA8G5XfX0IQuOdTsX
k24Eiw3ky6ezAmrSqiSxBvWry+Ig2Q7gG6OJaGjLj9qVABZzBtGgbAePRWDrjDHn
4X4Wc24c9DdKWayTxrO5IHJ+JX/VmEBL6nt7iTfWxy+ddA9mWi8o1aLuzbIgQAWN
AHcU4Cc+6/EU91aATLPT9B+hydHhWbrGpoQPId+xgaKjUrXfrs0DwWvSqPbe19W5
fvsf9p1QjzzGeNaHxKb/6FN7tKS5KAQZm/2ysTfS8WWq5S1Hq2XUgSAWLq30nyBQ
D5Z0Ss4cC70++SmEdoFOE/ubO7rUITWFDpX28L09sZXEQYHXbpCNH2w0Z2cSE+Sn
H7EglAoJDmFrjebfIclrjJeR0CtSPrrxaqM+iv9bh1MMvsE4qk2MSxCW5wXBP2gQ
smK87shklLjlrUViyOdPCOGYCaOGttO/PZAaOIs4i+c06id/tbr13LfdbVBQKc8A
Cjjd6qhvYB6U4GN1vZS8PvGXYOw55a4kSOWFjwQw7QNlsneDBkf7TGy168WG9uA1
z+CzMl6aVIv5CojeT29dk4xSrn+iZjSzR9wnXe6UqK8UfBl8KlhxMHfFH+szv3m4
VsgsFpXe4hXN+s37H5tRr7mrp/WXLYI07afqByqq86onQWBlpQD4GristOzyuTmh
zLiSoBpW+JVw8uZA96qUlkvZ1ZWWaxDt1vZrAfakjkXbblcPUypDm4P0MBboL2di
jVJmUJVae1oi9eQ3oGcaE8YfEYbYQ3C13p73x2Pbu4iu4hgnuvNfCbSJNGkQ7jtF
QiDTn4xRt9JD/WH9J1+xoPgqN5y7hAXKgRTBEr4kSHN3EzEMWwwoqADJ572KtuHF
KC/N3qbwC+wkfXUnt1wnUKUUKSilbuz/mnR8cHiXdLB07XdBEoRT8TP/nHgQvSWS
BlpF2zyaCY2VGV2SJPJdXLeoKSIhK8Zoce1Z7xVhOk6cQo7WqaHKt2QZUBimgFuw
rEu0Dbi5ZhopGy5SPjRtLVShfcHJo/CF6Z7q8Prh0GL8c4WU9XV+B5VxAaQeIoMU
BHtwRqmFC/l+ehBedIUDokyupmJp3kzx+e4hVveTweMjBuClBUQfAAxuMqBzWouU
YecCWLRzJ5gtI6QcDxUxwh3mi88DoiDeJepiXpQLn5nwJeoSgDZHwSPOeTa2mktU
mx65iY2c3VGcEWgL9B6yGli29fjIio2xwgu1dP2jg2TiB6P5a6qwnsi9LwLgmRVv
ArUyD4TV2hcdZptpgSVY+xbk2hU+uzjrHUlR68FQqHhZTtDAjPkXaPuOm7a59R82
IoUj5BnTsV17L4O0i/b4VpSNn+mIu7hQrFoknkpwPLcROTaTtZQoIXrJnnSssNZ1
Eii/FvRmmI524GShRsT0xvecHVXSdeWk+iu/v82vmyPXDjQgeLY1KB4s2+0SUHvW
2EnoJHf/K4due+0Lxpz60uIfDgbsCFx0A4njkHTwFiJv54UetS3lYf8Ar4lE0Bjb
3t7yxiEh0J4Y7NVZu7QpRT4jWSuyxprH5ql+2QiszcGZXs0bpDEeTNwCdJ6dCXex
IJE1931IrZIzwEKkWIf399c6gsfg6HZkfDtPrXzpKCIFLR0lGg4VORZdeFqM2+XQ
1dhS0Kr5itc+addcF+0wrSk5MxLKPVpoDgDQzmL7j5jgiLfuwOTd5GZA/OE/WTo2
3W3HuD3AtA4ALjyhbFywdIo2nj8KieJ58qVz0i4gB4Modq1TRuG1kRTDdxVQFjuX
/AJ2c//dOTC0hDMfHZYLa2TN7avQX4nEhbJr8O6AOED8bBoMSfAP7/BxRuckNgyb
Q0S2uMixfnR+Kn0Iw7hpOYhTPOFOS5BEN/WxFTubmG5e5dZIQSV0jzIJVuFC7e50
hijgq4O5mWIGULp5sQPat7BSdGMGciLZZI9vRSi2sxfRxYw2TK0YY3x4Q9dDrLXy
fG9BqMSF+oNrApz0JeRWfFeXBFQGJGhIndk8kyhtRJzvX1iJDtDN+UnIlG/5Ayfw
gLalt8JieU7h+XzAdSTf0x6nhjnplubkA0uSZDSx4NrEmcKECo5b8GcwCU3ik2aU
VpXAQt4Ddhr1QJvLOrhasqv2DZn8sTLG2eaT9dWYGSml3DgCNuQs97OQaYs5z3G/
0PqxoShcYuivN3Tb8g4xYjGYKCvbBNRTvP6rksfA+vPd8aHynTzFFnGOO1NZQfkG
jE/pGWiYHQrKXD6rAdXrwvVrLQSbsBM6aZU4dV+J4t/+QaXOFmPSTaZr/mkRM8us
0BAunew9qOl/OTm6EVCfXONivdAEgUayGEo7iaYa/FK1C2H07js19LetnAA6NSHb
3BARqzVz2o7qKV0ULjR8piphl+s+5W78hE0DmIYe6qcPs+R5oP1TqxObFxakDyU+
WNGX18w8ikOo7lcs1k3WJoJbJu02MzdyoqESVeSUTQWDDEEEGpTaB52zfkQ9/yO5
FRRF3fEWMYY6quP0IkAsjK6/zbanF8YYWZEHviz0BJ+J4gd+yVjO6Jv58qUudAsk
wfB/zEfr0CLpD6DMinuE7ONEun2wnEk8OsikvW7YfqJu9QD3Bwtm9TRcGjZbKUUa
GZzKn9kpQ4RUW35AU45UIL1r6NH5glllTpgRWxzCEoOqpifxtvYVajbIX6U77LF8
GqumW5owR4i8dqIS87cmmTgDt00u17FrIyRLyz9zN/GWxwbTe3/cZT6ckAUM65Jn
Hs1mIOwCuJEOfkjMKJpj8KrdfjDb2KZRHg6+kZOowpbhWgewWr0UokGryS/YkyOg
08rm3Ychz3yHcXHFkF3B3d41APBxRzfChnSWxkKA+1ySifJeGGwkBdSnfcZy29/J
0gep70FvTOXxp7QjaNuSRxD5uiReROgiKdVPswOOoM37eNreoHPXnqpjGhyGV/Dh
k/6vktePmCy3jIRbnoxFC13XF5Qo0pE3pasrH4OgkHa5nMgedTw6fBzd7yVSqYtc
rEAZiroCVIMoGWOv+Sjffi8L7ESW48ZLh+i5tNeZzEzewqGH8pacqTRV3ptOO21I
tgj3WwWwR9EUNb1cahfeu4U8gBovke9xQ6mawtkQ7br2rChnOmy3KbvKPj8ZW+S8
1ZwEzPw8FnbZ31jQqbNAnhIatzALbXxAOJZ1Hnl7rlNMNH0ZZ+rjRpAEQ8EudESA
GFYRTL/Jl5zd7t2794uvZPZTiiGQVUh3UFpfolYDsb7Y28x9oHqx/hh8BbIDhvoF
+WL7v85lcBXbSH6UtdjOqSDWLGxR4bQm/iFZA7EbptPZ5y5iORsoXkj9cYtPuulf
U5UOuKzTnoYG3VQ2+T2qpNnLXYrcAU7D8pHywVEIthl1DtceYWyhfcP+5YeuAa9h
k9Fe3aQiTjtok6kaMlFFDsHSIkqUSOgB0HOZ6lPlhneeZNUTUdjxMaUjA18w0d6i
J+lgP0GVXtBS08wL6RlJSuDMyNbkBPpaE5NyH1qE2xmSAFNrdYpUK5N7xl6RY3a4
GgaRoMa9Mau1pN24jJpSexiztM8nZqjv7bKJwFJ02hCjzjWRpASkjf3ILxs4U0HX
32fxUCHcLQWJJWcOMNzch8TLe6M44wT3UFVb48MQOpWKZ9Ccrx3a57Dabs06Sxy6
VaPwcmVuEk6ZDXD9iLpxlDWAFB6pTOWS+aAQeLhoJWmDzvXhagd40BstphEAyvfy
2zokk+nLLmfiSLv4g/toTxgMklSFBLdRyrh5mNgxkjcii+xIJKdymOmhkeGDHull
Ww2Q8mrFpLPbO8cfui5kw/AhDlML8PSecZrUJ1+hWtHpy+hKs9Oymu/eXunfOM66
YOOindQ2cv6ceUgdoIzgh7nF4Rpm07S9zgAOFQXSXfrGSO9uGvyjWGwR/fKplfc7
IdVZKuZFtrqSeOJAzUn8q0swxV31PiXzNAMEZwcamsMhpzye5JkCMx8zTRYzwot0
oCo2yoXjfw5JXXW4576sU7KWMlk4AttId6TRFkK27ncaE1TVUJ96O3ennAzQ6SeT

`pragma protect end_protected
