// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
l0cwpYTnFbx/liMhiSH6HSR+YQqJIzBVIL8x9iS6WZ/qCSHnpo92CK+qzGbalNCx
8RTZyCpw8VB0ppp5ACumg+qySniv7CdbWbm71vtXotTe6scCySsk71GDtKVEXg+G
cXhLtXmwGJG6AkYBFHPxgMPOwMCUypmIDZDe9fxU8Lo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6144 )
`pragma protect data_block
CocM7E18biFk3/7DmFGY7BK/Xh8vVg7Zna40ZZkCLXs2KYuNTZfj/YMUxe1JkpGP
5i6ccMgRt1YSZufN9VOdat4sa26t8ZMvVyJJXIj0sdTBRhmbGjK/L97Thbw4rffe
uhug8z6LyQLqScsRaQ9EhFXC7CtNqz3f5GRYsZ/LmoqBWFftokzVmTmpvRUCHhbA
payCONXGBZ8JN3ppaGzQgutkgJu5P6fcgo/4dJERuVI6FFa4cVx3VeahrRr8gAzQ
ocOk11LD/1NVBN189JKbxIzm/2HUeoAyjJJJJn33CldTyyPhz9ZIzxTquNy2HuX5
9rdJULtLCkhU+oSBFAjm1r9TmfbbJsC+FZrk8UIo0FNZXFdvQQeu5eTcAmTp1mvA
s4Fm6+QHzKYWV663JTUYxf6vURN1s/5ic/EIem0wdaFPEJQzPt1kGxkVsVPSZ41w
TBbqGyvpZnn0Dbf16OLGWEU1VluIrfgrU0FQ1KtagpPLhsxfhon7VpLfRwteebRe
EQVp0juTmAVTFtElhPE1N3yB+G6UT1yu/xH9hHGfx6/6+e6D56j++1yO/A0R0BaN
DB5JYywIwTPIZk2CY+juwSATeh6AzfI++srnB1YUOSVBSyRM5h5nDEbkdTgtJy0+
QjWRjEYk/Rk9A5C4Oe9uW3Rv2R7GP6nVaSEzZjgOGLPztSJxiydHWf1xSvE0Vz9K
pjfiFtvbAOYeIxUANXlknRSzsV2GAvCt8Vh4Fd0nyTgZVmMVCetZ6T/2S4ngaACH
iPhfE8wedGJTOFD7BxcWWWDXJPvCIXMu3z0DVHOAuYfYFQBkyQpUPLq3+U6Vv/cv
DmWjJUyqxV1KSLiym1etC3IfDq2jiotKgY5aLWSN3llAavJUVg+TtbKy6+XRxkHl
e7iqe45gjxeeaXK7g9anEIzJWEK6Q9/KoIVvn5sRntw/KQPuBnbJpGT6Gq0nvNnn
tZsoIDEO+n/iwcnRQpRIlVtA5YAkI1uLinb57H79SlX2xFhmU2fYPP/PR6E5zXBm
OSGMyrKUB6cg4KXibpFydl4detUQJt22ndxMLYkptx6BitsmSKHYjq7HHOhRS6rt
ySYyWQ9NNWL6omXm7YFCyslq/BqJGDN3fpSXd2agx0xTmPKOI3+M+g9EBxIJfL0r
EuUd/pFN2N5zbTI1JJ1TiiSYc9nu3ZBl3iSeeU6uuPcIOXy7FQ6CKSLKzb36dEVQ
sBIFKEvHqgCfhiypBjvJ9hUNgSGjTcAlR1TTHlp3UQU3lOD2+BUfJgTbTkElB5I5
sl9lHqJPz/G3yDFvGPx8YmBnTtPL/bIbArZl3amjCNcQXbkzzBdDZE3kgXYBGesp
QkUfvazX0jMbHg8bqh06uMPW9pj/VrSEFu61PamaE7ef0o5MIQJ0a10WlokZPTLh
j4FkQlZB2K+VZWf8GnYDqou13wqorcPABNiNEeIQFeoc1BAoXXNE+nwgFnqVvFdN
2axS1+jya6hx9JsN0NNt1cbG82YFXBhLbPM8bYXGbhyohanfZl2qNoFkC3X8B5Uh
ZN/b3nane2taBFhle0hxq/66btTFxsVec7wtJvxLUl3nERTtWufPAHaf12ddb+Af
SikM4EPyMn9ojPT+ifeuziXOadFfWfL84Nb/rL0vg/cqLWqdivcERJIKccaiBYlK
GEWgpfC2Up12LbxbTuSG0AydcSwQCbASEwmlrWmo+/MoDbxCNJwG7qdLXcEAL6cX
Js+hT40qHEGRL7To/91Vxg0Pk3+0nRBd1lDO+hyUHSMCOl26SDfEH+Q86hbxj4KA
/F24d20+ccjcLF7gyYymcn11Utj8Z/MgL0Wnj48hP6V9/oZqQzIT4dD4pKgDO66f
tfng8BgI3SW/qve7di4UlNKCfoJu+H9EAHDxxGR1Of5ygKvEvYNw50tJHvDUig68
USijf/pNxXUiV+c6iemGm1Duc8YKC7tgn2z8vgrW7Z9wbs8t/1LO5awd9ObIzb4X
hXYQZ7hj5gMZCLfqqQZUGC1Wd8dy+3/ejbqLN80d7a4i+arQJZbXymidIc7icG1K
35OZDiKNgePFoeXXGD2TCEkCPvQYiCVMGkOwlNbW+vGpVsZBST2K2UNku7ApZBzP
gbcAAfpGsxSJkmZnqiGZXAkYz4W7LlEVlPQOF70CgzEtjX1HHB8SLBfG+fWCW7Qo
Delh+CJhmzxYxUpSQJg79H4dwkPZlbdk+NmE4/N766weeOB2r6ZXHMo2NEPrDhgC
0H6jSi0RS01gYVzEoL6R+2lJzv6VWsts91aTXliVjHrRH07uxfzociyRBy7IviNt
TldYJV+e0JQmyCxZP6OAc2SD5R/CSQ0vELKVkz5KZ6ENDFhhD7lxBbhWVcrNrzKM
9Q1TjdyXibwCgU/KmrYag1Pkfo7X7agz3AK6fSSBXigYwDjEy4EPWZAUCJYhzAHm
LRMNfODI23DVw6itT+nRd8vdIbkbAmIFW1u1bbFgXHlL79K+pIkif/6LsmljT5VA
TC+FPcd2shW1HCyvRjXcAu9PBP3//FYR7EXzYNpjE4PpCj8gMhiG4JfpDKeEsUzl
RMhl9aDD7hx4zYUBJQEM5Gta8hFoOIZa3fZcGKLpa4rK4n/JH0C4fhLJvNcjgC3v
UxxomYzSRoPdRTgPoJbVQHJs9H56smbTogucEyrgNyQbjiWCulbdz3F/QRLrMmuJ
LkRVA5Acqyl6W9TwIl3LRleHi0ba/J1vR6k4HQMUrpYDeU6UoXUJdxdDIPOLQt6i
VssGF2PZwktuIJVRR7P82VdhvVbeb5lkabHIBkQMjndB5Sb/eQe1ik4g5X8OUIwr
NqERmKqjDoow2ZhjUoEtmF2ViE/SiSTQuZJHMgLV997s5d9yWA/EhOpb7mWHakSg
VOnJ/S0Cww5a5bFS/0gGysiaPGStVDJbcTdjbXx3tXdpxXu8CcHPO3vljo/HGvQb
IPXAb/mr2p/IrDOmBXDljVsf5eAV9blM8h3b5GYCLQ8iRz0SlzRf3GhmRpNGAxA6
eIo6IONxaLMlYSmhBVIgoOQbscKT3KvXwXj9HgvX+DeJKZ6ocmmYdIkSjB4U12wK
mTL9yP2UAKzM3od0lyG/gTJwZhnkjm/GWNWiIJqmlzP6UogvdAly1McZm1ckYYrJ
joP4xYyEefyTBWNI2OYnfzimcPdpRMHglbwYAMV8+HQE4AecOfZUZp9DB3Nan4G8
aXMkEyaYHNd8vQvoJEfU/pv510rEMHoEtgfjF0gfGLlA3/SrwhTFMw7zCGIf1baV
twE3a6IAtH15QQpmqbdKuXLXYgzq9pbGZS4oPjxenDbV+wadvwvDHKMnySHzeUWH
ULw/2Ka6wBdOrpdElN8MUgATkmadAyAWmCKVjQ7FSRw6TJTyhRy9Tgrv1aBfdtPs
qLFe2F627YpoWcZPlE4nrnr2pztqzlpt6BJbH6M6zugbu2jI8o3q5XmoO/c7LYuu
OzsuB+OsfVfsXuxqZMenhfL2QzW0zU0JZDi4msZp825GKuznQXBbfYO48Cl7MrT5
JdRIFfyFYAQK1tU8DVc310VQxWPRe5XBmgYsIQ4uAJBSbwpboAWWFPz7DCSkrZJM
/1KyrT5GqPMHKwER11BZdgB2unFKtD07i6LCl39EUMqyajANsY88VFTebEIVFn9I
um+lGBG7P2PECa65JAKL8c5I9q6H6Mpcu8LbAJcOCONlP+HXMufh9y7Wd9ttOb/1
ubpcAerF0Huq8uXIoj2Kkit/ipVj+ig3LXZD4ZKhx9u3qkGOOi18bk1UI1EQvnL4
v0Be/f7ZvjTgYB+HDJ+dv1wXnAFgxO2RU5NcS0JDOX4Ar9hVhxv0xz4TDzP5JdOw
FYaDTWaGA1KCPyWDK192qkw86VHy5Kxelpv4Ased5OTtlLe7o3q8yqu+uGZHgGON
fKVPX1PAlVL6754lmuNztTJ0QYpHQ+i/a8eT/zUGS99ZKofi7xFvOZaOjdKzW2rx
D1Fxbvod8h3Wk31XD5T1/bB5WKIslLrXj1Eu3+TtN9Mmdot3XPK9W+odtBcDvKBs
kBPb0sbkZABpc9thl6kWHeKKXq8hmjBEKBNKhdg7d9FebmjEVFf+/Z8G80HLGWlc
yHByCr99KBLDDuRO53V1EtukCHjYgAjqwFWp74c12LTJ58OjguvEELArsLX5epaV
/UWy2HhTVLtcmbdnhuFHmTyw5jrn6JIzwNyWDwM7Mv6bHv3C+d/eHeJNwOSG4k5u
uvsYW1dXMhoi0sKjjjL+HDHAA+cKKFCtEUJeEvmVKEEp2qeq/Yvb2AR92mwv0v59
cxKoEy+BPUiaIs0Z2mgxm5yG1PhYZngHY4XDZNSNMtTVXK44T1ynRd2VbVupiNey
epcPbE8GEe4rDHfpUAY9GD9TkplGbrlH0yNPzbcwc9g4sXE0Ko85ZGFbEZZOvTkm
v+tBuAD7vNnr7iEeD3FWrX1NXML5FN7TTT2OzveZfTbyVuuSGjKLdqGzhs6ypF4+
LeiYHCsUy4sp3f5ZhvuwCbc7kJtGvajBHszoJno8eQUOSpEN8v5aDLcAWhGt5fip
wbSAWvF+WJLpDyO0ZLQx8iEHgUv8oJWeOtBfI8D99qjrF+1d0P2NKFMS1thJnSD5
fb7LgG8O1mkM6JGkr/9JQssqViVmo3MPzJCxK03LJNTNLr6y57b0V4saTI5ljS5c
n73b59OScuvxQu0qW1yynfZwTZB1hMEAt45qVcAhD0JUmuI31E4R3walFrH0IXK3
LxUBqIHuLLok3zb2wtE5Tj8fgBZF8kS4wZ7oRbN40a+9nZwXnTQjjvn94yvuU5df
hicDX/XQDqVvf1Rkxe87NghwSFG+zW01epxeLgP6+pp9ie4r4I3C71+fOKJdJc27
v5auE7kfsCPygwamov63AmviE9Alqu/7riMht+HDPszMJ+Vq++CTJV1Ea/D3eppb
sKGUGZ/I8EoOQKvn3Do8nrLnwQgFxuOJyIFClnsrP3/7qiGWqu1PyWwFu+EisQ8v
qvyG4ATJ2uPDPgEy+TPwdGfxIiyutp32jKjKFlcvFrmalA7xFSWyBhZc2IjlVg0h
sPHXfwn5nIs3Z0kq+0Sxveud9LqBs3N5vHgWz5wkz8pnvYLoKuLvmK3f21vVwmpl
18dTzl2hI1gvxGsK3P69j0ww26JKuP58QrghY/1M4QQMa81K1+g83v7YoBl8S3Jm
qCgg0F5aTrgcOMhWjbzsD84ALIPLfT7nnAhCeqqAaMKonWoQ46aSDMREvmyYMaPT
V+5ZUrVraLgpVAtHZ2syMSmeogFaTWFRqQS5sfNKTQ6QVqn0bUcsVFUBB5KRVMIb
RfmOD9oMUVq14WKyrfASwkDp+LbYMa1XnDI6zs0KVPKUsEvON/TMLvXZNeD5URRF
94waJubai47Rp808ZeFmZ5KksUmV93HBjlDAY8WlLejj++uh5R8D8dlMlGJKj9Sj
vf+0GkzvwG6thBGQ6wx7kzOt2Ef0dr1DBkirBpmIl0r0IipM/1+NBPczQl4R6vq1
uxQyi0Ss3je0mHEmXGunnlKmDMJ+mVloWAfcYnXZ8pDEP5Ce3/i5bKI7F6773hBN
P8f6siQtfxVXgp2JCrleTPKRzPSLjShKfWoKa1m7nWjQ3U2pBQqtGUsr/AcfrmmY
LxiF56rD3eDIuC121GOvzLtcmKSpp3muXDbfMhr5mvRYeL9qH7a6r+T+rmomo9VV
QU5RvvQ64rCiZJZu42C6Bq0llWbZDPMPYAyXziAUQd3QDRstBMa7uJRu8Xt+ZLg3
WSv1iuBQzEmWO4xiinwM0n26gixvWCzV72S5VXkNAwcgOimUjb/kJLdJ85wDbRie
q3vg42DHoOn2hiUKPnarn5XMSfuCpima12EKE4aCgXHg3Pq7cF4h9k7BjopYTc3k
UTEnRMDiinoFYpm2Lu3aU6KfLJQ42u2o0q+P0DHEbQTx/ayGLzbm8tq6gqf/9hGc
F14cgS/XC+JtS81dm1KtBCSSeD7qOCepOy154MJMKISsy4SSps21xEX7lfouXsib
duk9pty+7ocDMerxl9FVCf3M3tcyuqL3HZ0IokYRgBa/Vyymx1YpLDZtchgsA40D
8mcWB2ndpE9tNNnYmP1eezT9gTa3gQO3mwAuTIsuNm21tKf0VbhawI23sXMrL0Yu
z7uBy1Mt/UI208pKKVXn/izbEPsO0Jo90TPIZpyWLZjBIlP78EenV+uyJs4JZcoX
a+8RqdoEZleS3CGYCqIFkPvvd5ZHAvsowV23Hf2QH3CjseTa36PCSUWAGO4Nwjmw
CwHDAkv0jrSkGTOsgcRb0VG/Gv+BbugHbxjFKWb0BjwEX7fF2+piwSFhTmbQ0XEq
sEtP/p7hffMd//q0x+nCyNeYNjyws6SZgrOuT2VWj2l4Wqix7or64QW8qX7B3bds
Aq0KL+AMq1Mz/lJ+uG0xcEfevZmUiMFSrRkWiMtrr+tnLsTiZpbnYhEg+dU9aLC0
x/wF9UruIsR0FK5BvdLyiPkKkvUjzxgINQd0ASsTrO0O+XjlQyNyAjxjEpOP4Vw7
PjYLvy4IPrmLQhNUd5C1yGODkDTlohIZ/8WTUz1eTsp22rQPpyR3VR0Uk8CqziNH
A38B1C5+UNZnmYhHXyjwalbGXdVNtOIab8TFvfDVlvi/KARnaHxnHeoqwEt+FnO8
cn7cPCj37SBYR9gdGvMxp/ANzO/PjhM4T8HkaR1AQB/bQupWa15FOSNU+d/vb+2F
B1/QTXJmV1ZSSENPUUfLFwIfs7RBmVBsvxyrBVUIE0OhsnlQOMu83sFwS0uWebXm
Z/zapA8OyNkMz2jLKXaXTk5DSpPtmpX5zeBz+FNQavwwpCszQWzHr+YjEsKLzXKK
tSicXKmg4+op0J8bAqMe9lt5AilezxhqQfgb35TVEG9zOXr6mAlcYfU+HYCJdXAe
YsI3tnarItzZGNI+hDHMqPjg1PdkodEytZ7QeqsU0MvZt0CSTDAnV72qX4yiuJzL
VVXjrVEFT54WfUDU3P7QUKuPV/cZxTnXe4PGZLjcDx3goSlxgAldl887DZWT+CR7
0UIAQ8IiB3tqvPh3T26dh4zPr/zcDBcbeOlBo1MivGCnPXl9XXMG2AA3LTxPLuLl
nBA8DSWRUOeQg+jC1GH6dajxLWlxy5V/pPb+59NpauyT1cirrYJVpsb+x2JikJJq
lKkfeLi4qJeMhyU5wixpaTnxfCi8upl+Wuan4ZAPYF01pg2LTNaf6nifbKgj6V5h
m8TebRG23US8ghMM45ZS8jWZNVtJx1Ra5p7V52cB+n/HdD1BNORLQJSpRsaW/Bos
QDQi46hJ0xOR2vavMNrTLCI/rL94CoUi7YMeCj9TURbHe3Lr/4WYgWop+aKg/8uB
NUp/ge5AUcWYC7MBpUyCLTHnMfnSkIVCpJ7mZ75ueIhL932X9ULDvobqHNWp646h
+U3L9sh574SOOulpiLtw9iIVzbFt32rwlkW0u06NoP8kz1Fc9R89kdPTQsXLvKV3
0CTQ+66JnGetzMAxGFoMdKghwsLkqGChkrdeZh7KL1zK+681AeIykQ6zdTzmWjJv
Q3S2NVt2IbyDMe5oQ1YyOKq9w927fYNiIe/Jr87Yla2cJpcz0m/SgUadqUtV0Fg+
hXX3KZt85p7NN3jcZfWlJDUrdWpFAqN9bcfwK0wLEc7ajfrWiN2FNOJHSkUV3hS+
aLdiq3GVYTDfS3sKuJc8DTIMmg6Y304nUue4cw8CTTgcgiYCTIU8I2+01y+mZU7t
Y/lya1dGTmd+H/wONcMp5dm/fqesNggt/AGCttGMfaU8WOJCyWifv/JRoLqrJ/tG
MUk4OHvQbrhGVJBWQeWEl6/qAXwnzpcYcWdv8EG3Qidmu736Chue5Kb/mTdeNB+G
eOVZXkj7m6smMNSsOZPyoPEKAEKEPoQSvbCEResB6ODQgduM7WiYOelrBtd6LGnA
mvSOMirqQ5RXWHsQNOLMXT/kAkOakMkzVjsQKOyhSo/Oy8ojb31wQwisI3suGZIa
/hHyhp2wEO9ltTX/WZYMSDvhiKFKvGgPXiXOxgUiP49xjevn4PBk0Zg5B4tRiQpp
SPvLl7qLtIUF6QshhZ8LfsEbx6YxAc7Q4IgLM1dmkzxUbMCCx5VyCEip++ruvc2+
Js8MZA01I3JP3DDPSBp2bm7odZMBp+LEScQ2VSKt+b82NICNjz0L0Nn5mGdhBwRZ

`pragma protect end_protected
