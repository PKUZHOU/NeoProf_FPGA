// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MJCzXSPDh39L8XM1OFbRYoEs+OuXLDAFmD9a27MqgU33tc3OscRvhqG/qC2d
nUcrpKpD8p/cHz4+Ojba1pQTUofHpvqkO2pOaSjukE6KWLjxqxhW88WzUFJv
dbymX8fQYZZqKKg8Xv1XzECoiZwbsKU7xOQZFNEioFwpUgfAbx08L/z7qchq
gi42wkdnADk7ef5hqylJCTxf22mIgIBSz6dVSNJjyEMie6fwHsvhrygrOEqo
urr+sBNOLHvWVOPqL9HF98QHXdvUBrYtEwzgVgXBEtM2L6ZTviJlCEJJ57tP
1RlJIwQFuiKOmgqq8jeXcIBcm80Fp8Fi+FIwB/5GmQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
caOXAXxlwLcTXqPQZ/XHE2g/DzNppxmrOqOmJKSyYt/q8oFgpxjZdR1wu6Y+
wo8FpxHCw9l0Cj2XXyF5xqmlizvIExwE2ZveHhHqMeck0J7OgNwrJzt1GSGg
elaeO0IHrhmPraRxBY6GhNm6FBROc9vw0BVXrjK7px3dZs+GD3swg4sV0mf/
+vvrv2JW4kgfQQYjUlPI7EmHdOPmSEhL1h5Wwvyz050p0CBb790hJikjsaQ0
0O1/+vALiVMcwGpUIm63dYNVJGLVvylcUF4L9VZf0RcTwW+Cw0dwzMAOAMeC
ot8Yhu8pAp3URk0CYrt8TM3O1fKoZvdV7dsxSu7GSw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VNiNB8IWs1toEd3JwlndP7z4TMJ42x9Dm20HNpSwc60PvyY3Mko+iEIVl8/Q
XQLhYYwt5bEb5dNRv+fHNTVJboeO2kIb984jBoOknlq9aSp1Yp67KkYhT5P8
2tiattDI2AUoCGzKUk2mOtW9KMgjGXmENG5IzC1TEPLAZdfE2/C3BF267J8r
rczSL9pAwwoEu4iHUQkAorr6MzzaYSa18Fq0y9lnxDpvDwRWSzC2BvpgjeLU
w6ZQCno9gzylFTZTNCNoQV3qDQM06ZGiBerx0Jrrsh+nCk6R9ULaGY1TdPWW
v3CNfOgpsINDtKWJyOqQWbYSo8KqS6dmq4BUzGkTkQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XJ7gEh+I8n8GBuqOHiAU0bR7bV4T+rsq8PsXqx6MsoHm1UNgQALSMrjvVukn
1rwvOsg9zoK7t4YTeBWoOhNC5JgtCuFM/lvNYuIHvBoof6PKg8qWub+vtqrm
Fld5yW9qAJn60svwsKvZ7oprdV/5RSN3h7euh/j+PW4se+MmKtU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
AhcD1Ds/z0iPyDpIKu32gI1esBtOs2ehmGTbNJ6aJ4PyUQCWb5yg3piGjB0F
R9Y9Hkl+pxaP+dyzCMo3Dx1x5fDdNkZ4620u3rxNll5+grNt1a2CTvkRm5VS
6hgjhCEJYLzlcwsHbERFXr2WTeRkoNWPRyCycfHLGzoazKIaF64rRIhUZ8T5
O619U95/5uFEH01OQ1vXApgPdcYu/zKSZjRmY1Ur3pdrruP6QdZOLNFHQI6H
2yw7HfoWLSkTuKWrUWZ2YIQu6HAoV1KxO58FJFAzcxwC3V1+nB8fixjhwT9Y
kQwTVm1J8MhnU+wZoPYwwi6dzFlZ24Eb086DN5aGLD/T5BG5/hkGlVBZsEt+
lXiw3aPBQiMFzVuTCWnw4u1wicHi+8uLFO1xeBPjO3T7BS7LVdum4iWZAfrM
Jiu3gTjiXgakI8gStguWikD/y/Q0SQJgyTT1k7g2rZK0uNdNzlQ/d23kSFqG
yOxON77PWqfOnfEsGsbEQkoT06x3ljWq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pL2hmLbS0BTEGAO05wWqHowke/nRqMKV1cRgtMbo+Ta8mYB2cqAGXlzFI0sP
weFwAhMRt+R+pDcSUwh1hxGqWOVzZCaYl2QQngCf88ILH1/KCdyQlLt6c5LO
pr6ZbIL2sjky2s47pTFiOSOIFy4fpxus/brPPfO5xrfLClw464Y=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pNcfAA53nVWUuiwgjWVZl6qPvp7bpqschUUgyajjqRWgFOrT14WY3bLfkeiz
RogmLAWtxXp6KQSaQvwQFJ6cYymxljoCZACJBsMzWyb8Pg8tzL/RklkW1/g1
Ss72xI5uA3BZjjtWaPWkrsfIvfL7KZcBHHc8fUkCNopmg1RFp9M=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 106272)
`pragma protect data_block
dwWd1byr1omuh07lEPbpGgAQdAm53hDBBGy1Bd6cbqBkbaJpAeJexGh7qOJD
daycR/0U9WJLpXfCR7bMj60uplcHSv2DwHbOutAbU5x6pBnh8+cTXi7Pfj8H
HO0aVQDZlFOJOcAJtFFtWxNgVr/dkzXKVb1rzqA4dHw0pBXEnyOyyd2gBIV9
HphIiBYxOf9Dbba2y82Ca5P2ASyLblXx/4aZpRJg5/Iib6/BB1jYuEmSxzM7
oDCCnjWDCqOtYyuUt72BkCMQSu948OMQNsVc2jdsULF9E/TdJqQFI7UGLMmo
RRN0wdQxIf7VDm33pbjfnCJtYk0MWkYH895FmhimV161oS9y2dfyc4nrZ/aK
h6g3meel9PFa0pM+MuUwLC68/Pcxd49ypSzHUVFebxbRYRf5obBIu91dfYkY
PHsNVWWG20L7bsAO8e+A90pbb7oRq4KQBorit+w4E7iKksjteNHFTWIO1n4d
xUhkIwZRzkdYu87bjtxdcFmcRHm9b5bJCOZqErCBYAjMKNOY4TKekF9uAMzN
0C9/tfm+yD4fzfBVfdLbNeI8pou8voXwXj5cYXiTQLaJEn861skp1Y8OtzXF
1nysB30pwEcRE131BGbjGhFhQFr0jszC5D0SxngYDSjiFgrzuBXRMaVDD8la
DpbMpPjLx0kAwMAjvfNTFytSkb3MJvg65KO+Usg1ddU6YamE7Cmt2mAJXLlR
/cN3wUR1rl1HOpM6U23Rv+I4RixuZoLnzFCeqQUJhFczAYoV635RWJ0YBV7G
+3AmbaZ/FtuYB7oWLp5PvzfYtnB2pnQ5oRQEuL5Eey6nVG1vuyvU4We1Rv72
4JYS7EkQsEiydx6f/uaoHI27n7fr23ftudOZzHm1PO6oOOdOyMHjW2+0LOJf
0U6fDOOYYC6KrW0icoEq7C1hh2chbMEyqE3ji125NbEMyZ0Mh5i953XObjH3
Ggey34l707M5pIoBE32HVlcIJr3pOlXXhPGvqz0Tr6ST4G+1JRES5g2vB3W4
fsGROsjGuoup865Yz35BI+OogTJmJePvzw8ZYlVmL35DZTBXC1cvbIquVRm8
V7Y1fRMke0vS58nMccUGJt9I80VmpHcjusRJhkUtpapA+XU8l+N7Ga7ygdZ1
8Oqv6BgJnrtEzHgKWQWZBYuOAtq0aD08M6QSIWMtIfRt9RAUN9pI94l+MeLY
PA18UiamrrPh3aGNA/lfS6oE+kBuLaJvDxwHnLq5LkUas3VHGcg/sDKswwdN
OGi9q9TbuyIBRnVZgBhZB4OlMYsakPrFFaz/B8kNvVSeqUiV63+WmDgPFBbs
m2iEvIeaRSQOJQVF2s2vwAkz28pIwLRfFGJnezivIplyvs7m0j6oUrTO4HKh
w7beCidVYyEEQXt5jHlRpiQZ64dQz1v6T+EvD6Rwr/phpOQCBBTFaiy8879F
FSMd9cXWgnYNL/dQi0uoqS5JfjIWpXw9jsnwmkyAKPHV7/+pIDvKaOrtOLwb
NuMBnRRV20XKvnijwpAvP32EkDrQlfhkYrqhQG3w3jocBTI9XOop/m0oC6tO
99uvpShXlcNZZTlHzh3O/VwIzwcz+kbXU+00PYsXTioadu48mIFR3iNOOdck
m//XQasYAvuMS9SFCbuPUEr8ncCUFfHjGtVIaJ62EbX3jizhws09oLGcsq95
DbVJOKkSExcmOVEu4Ki/nBeQcpXuY0IBLP41aAAJKxFKUqKCg0mL/A9p1IdY
iBQEpri4xdByBaESBUtISR/qud4bm+tmYz3VDRZji8vXpQt19HXt//MASaap
FbMU82hRptoVuP5AeAWzAqxnZLPqF2vYpu7OXb7WUq1xJ5Xtpl71owdzUuMl
lzvjVBPCfBDqs7ir6NxXlhDPt0UBTUzW2ScrcU/U+yqoGb6ugPz/y32O57og
DqF5hLXOG+HTVp2RR2oJC/FENqALOHLtCmoSlzzOtrqHqIcJobrBJb4SnVen
HZonAR1WEELR3zkDcJlo4mxqpr6BzdrGk+8msMx6EhHC3JLSuo/F2zu7J3JO
XiByljUwKxgRh6MeI6FMaZyWPEqGmz/6Ev6aLANvxYXVnlLXMqZ+nl8ovsly
KW2f43QGbiWLrCBlrVFDBpBC9PeazxuG/UJS/+dSpwrMa/YYSq4Tz7eLg4j9
q6iQQA5MYkyl3bnGmOAdNIf+xS0ZfEl3LsU9nD3m0HpyfPzCCIk9Xufw+Nhh
lFeeMhF21/K9CEF8eerlwx64GWqgD31pG6YIUPVi9y1TO4ta5k3P9gcRPQkh
cTgf9JYFKaYgAiz+RSZ+uIOGGaosovqlHVF8iD1IZbjgkZ3Z9PB7WNEV4Y2g
dC/NRxUos16J7M5BQc/aG/T60rZgoT8rc2whk48TejXrHHYpLYafaztCg4M+
i5O7/YgKLUqtQs00fGz119SI8u3BPMF5k7b27rTqcxh3BjkuJCFwiqudx5cI
G3S8ggnQIin5xJ9L6bguMqJJCQedaaGwUw9Uw+yRvocXtpLOdI703Q4XXmN1
mTqqViAs+UIdEfZU26UZbae0lZnnZyb6hoB2OP522XIo1oLLJ2xmNej6x5Et
D3tCPWWzBUrBVZkqG+OpujeCV0SvgTOLrIaJEOTqmDU5Two7kYTVwuGUc+CY
O2J51670p7RNFR+fLoHH9M0TOHe1qgdI0yG1WHcID3RFjUJPVb2RJ7FRCkcD
ghyxgAeXw0mioblVjG9gUFe+WqZFwCiE7t2TNpPPkZZcDfUt3wLlKxK98VYA
6n7Z7w3uzrHzFoVAsENm2L3o2NkVAP8c5Y0wMJQhwgY/xYkTHbTWxFBdhn08
d9bsmsU5vCRvEVKBCrw2ePRxHi5fqF0CTQMcV3smAu1A3BeQocTrQwUatQnF
KXf2n2ONNohlYFy5e7rEwdJBJ4wUP2D5+oHCmwkTg/FCfZkqDaZzjt4KstdJ
Q3SgoJiRXXDwxnUXEHn/sAAxxPqVd/yF8FceFRL2zvWYaVQW2m0K/51iM/0j
xIMPPSPoEHv57tUp+zJShg28nc6Yz9ja6s+Zunmaoc2wEki/cuGPltTB3QNh
oICalwZKxh7ae6Xlux49vgrab+zJOtrrG7vElhpNUor8Z3jplND93f5c9HuD
nj89gYa0qavx4HCxo3ZWd3gRBiFVV/FeZ+3raO8jzSbt8UmOXlGMrj8M6BJO
fhTaFKarb1z/b9XVq0/amg9peb4A5HQf55OskJDYQAzbFmMoXhqThxUvvtp5
KoztdfdvGuwMChWRIMvwFkqFw9u/KBNanhXB5N43OTawxCdR+U/2qIhNf5Gc
LhfWT9NOHzR6CZbkbw9ffo40d2THMjx1221FfS7O7GC/IM+gcyIpt3coeuyk
0KdNjR3lh+2ppYPwe74iGTieEyFKnIF1yAB6LVmoXg9PFv4zrxMKt+/qpLpV
FMuExvMX4P6ZkX66OFDcQ6fzwuEpw5estBIl8uehgAdddRXuUZpkOdWYOfu2
bJqkCesy3Oxa/ryPtrv8CJjBj3cJConVh7GfcbrZkqcZ9VVyPiqLB1du0UrW
vuxP4jh9Z2pO44YGMhRKHWlxqMFdFXrQ66E2Udjh6Rjx3puDmv/xC/JHunWJ
8Xm6aJaLzjNhvibMoEhcKtwhPWkmYY1UmF+iQBa1xqVm1jI1j3zB7qTHhi5l
JRxb4JPxmsiYEm65pemzC713EKbD5q7ET1ov5/GqEZl4n2FyLOZVk2P/YCEG
B6dB2Ap1FZCZkqI5mqrpfpP1gWyuL/Q9UQQv/GZVLrLSekOZce53LRnQdPKD
LX8Dljx6W8kqQZ+pZjKYgcVRfzsNl5Zj4upsYspOSizqQfzIRrHlVQMD/Gol
ISQpKU7G0GMTxMhciHcv4a5/uCV+kca0zvBZ07FAGGjFkZvQYewT565O/cMZ
dvVXHJCY5D4RctrtfkUFmzFamHbiBCbPnpG00tHCp9SxTYw+BIHIS0bB/dZh
S/tkXluzTLigOM+61J5KdJsZIi0CYzAZbaLn58phYVBshbK61Jco9zClRvrJ
pE39pn7vfk66Ijkkzglarc8MLEc+R4Xrtjh362rtVf8d4x7gCusBY4Fk6JSh
dNo1i8ilLKGlTm2fCipFyX3Q7bYQLgYTDtUxzOTbcBEdjNL4OR+CwKfkaieI
DIGlkKb4cxi7JczpyeOlMy4pXEqKJZxHSMIimiMyWimtlcwo8Sm1GPYu7zGs
KdlmHBPfhcL5/axEHrchrbzGAfEgYngK57UrNV/+6/hPhhL37wnJy06ovGHk
05aUf4mc5kMv63uopG0HJDeVUT2hDOiXIQGakBsLh6v5eybUjXDuUbipv0Ch
g8oQrxLw/0QqQRLlvhxnDOQZwy4FBOoDmhTV+HZYDyhVrQuzANLNjTMav7hn
GqSXi9JWgg9PmGAG61IbncXa1k8/2t7HLwaQD0BroYNV2YsWGJ1RChYDL6pb
h7JHcxV32++kvwPHW9GRDowAZRFOAErZgttZ0ZlfMs8LczEuzlwOO5ry+wdU
+LsMAQNKkNImAuPBzhmrF7n2HT8V0VFPX6oWlTsgLljTmuIAXrOsvofSlN3X
NLHhQaKEv5h4TqM4WAKa9WnL4Y1z+IIVWfrFswCiG9Mve4/cHcMPrT0uGUQs
LSFv6jLMtydc2dd/FO6ctx09WfrZQhRZIUfNYBYDWt45dM/mD2JFDrLv3A7j
6iPvG8+vlfaBgJn3vlt5QZOwjj1NGsUP++JDkaTt89PKusylJhxrJdlG5DCx
1LHr+8pcp5e18ngIjQBY61PBlmaPHqe8tZXkHTd/PCKxMoZT5oLcATTCxoKz
rKFfOXKEPjCoWSn50z8aqgsfVG5p03aHAfO/aGf01ikM+p3asHyAA7HKCvlt
TnMDCP7hGY8dmm+RUw+zMc24IiRg1Q4gEELoZcHJX1nlm+2aKF9obc83UPQO
mYDccpUQo1kpJQoc1hX7kXniPIQgBYQLJB/WK9D6mIM8b22zi7tbiTIlatUZ
qTBmDEHohosOtG4VC1ecoUGz0qCdBtnytfedB55KLy27jAEtG7EFf/y7xUEh
b/B2s3KT7he4ylHqwl1OMedJc0JdpDuuDTct+QqmHk85k5BtSVRGRPogkpri
xxj0C1Jcf6UIDO054Mex+cm2+6CGToHE9g39h6glbJoK3uAcEH7D4dh/Be5y
npFzOLsKiu2Ehp9WKYnTMXtcRlJJK4DfWXtttmCKKOfFaLyuCUZA/TF1jvHD
PMMjo2cdsJ1jO/lMlkVxcGlXWmSd86p7peoDNIt+0wMz3PZWL+e7UwPwSV7e
mRVJ8Gb4TuMD/J0KXtF0I4HtX0jtOWuZ5AXkW0yJlpY+xgJtjAicJvHFxKlV
Gf+lqoxbfdnelhfuefxj879y6Br3JooBZ/ui8LSBmUkKkV6GHyS2Kmlj61un
3VD7IPVWlH9O/9D933UWpLDlb0FUFsJSnV9ZmW746Ej2gznNbtTrQBYIRPWH
FG68UWW0zDOdmfGbdOGPTlcq0oNYNpmbfYMHEnQ3a4nmOISmPEGxLQTwQhgO
4Minlbu7FMa8Isi3O1/9fF0ab7pUMgbShNYTNMvDDnfwRbipHhYu9e2u/xtb
phVsJXUYcFoHepo6CE/LSCVixsVS0rjJS7ijlQ7CQHcW0W3lxoX0RBIrj2+7
Pgx3ABmGo36Nt9WHBuJqlmF2T15Sm0kQCgl9JXStXxoryIK57WC78L6rZa0l
sC24Yl2VPLBKXWL3dtJdQkkagjuCMxBjz0DIu8pcvRBjTS8BUe3ZgvKYbkOI
x7/zv8j9PU3tREBUnmImnOBPvxeVoBgT1qz7WehMrCYGMoJAN9Q2R7fjbpHY
l8ISWwXhRV1/QtmPVF95wLfQ2Eb/zvF0QTeiRA3qP88HJA0yRLD+2MaAoQ99
UT/Q4cTIYVCXgJpfcGX6j5cNxsdGxPenP+C4z3+yiJcKBxN6tHZ5/wq25RZI
13Ss8HAzLGIyJI+5oqNsMfGdvOhUHFOxgeeq/stoM0ajPlHeMnVpnNM1RN8u
XEGZR2+0pansXAnfuuPEOzMpT3KovjHNlQEEmCGWsn8J6mWXoH9KKpDOKDVs
ys5JEJURK6E91TFFZL0LD5n2n9j5P2/sc6/6Uynl8FhFEKCtkRVmDdtRNAls
dK9yhKu0alm3o36o1Lz0gB4uJ4dPlyuGjtYWSyGhKpF4R2e7JWTVFvuN1D1f
NIT8OOmXd9zmU+hKkRjc/dzjo1ksZ0uS++oie32Gd2Y4b8ZNCzoFe+XLSIFr
O4PXxFTQxlBXTvOhVB91Q13+incJZ1USsr/U2W7IWUYnWFlBvz0oEE6+rdaP
21lcNymvjjfvCTMAXmdO3Uma+HmbRguOo57/taO128c2+D8XOz26hQ/oGfYk
SgsGJppjJ7ljas883wgScaBUw1NN6IAuVsd0QrZ2KY4ccMigGzwLItld43zh
D5VNT7wNwXRYESGldQpXuijPoL8uPOr8PiH0W4hbBYaknRoMrAc4wJn3NPPb
F6xCI74JLYOcXYurFckb7xjZK856xr+nw8gvlfWbsO/b7n50pW/VlDDE2kXf
J6tEGrPkc5NHYlpIxMSV1FMN+C1F3dJbYHFlYsWsovVI2Q7rWNcZw4RSCF0c
26HWnQkQWR1kK3YyZRrn7wm+8BdIpDoxKOiEuF8UQvVo8PmlHC03YcJPTOba
hlftjg6/QGhMG+BG55THEIoNvaqtNw4mULWNk+S4aqpmtdE5xrBeXW2/HvWQ
KwZS+g7Nb3Zrp4iiuIVKy9ESQS2qCPgU7FqNttXQDWPkypP5FO5NQY2dxA8c
J7AdUmXQgK14Vi4K8KgYAlPn3HmPXXL+K4RHVvehHwWpDVmXWhOhoKgWkC85
9dEin5AKeQil2/sySn9Ce3iHuoM34wq29kucvLO2jsUTUaNMYJru6Cek+tSj
quHUQQw+O9X5wTXxPeuyGbH37vZdw0oHIeWSNpY6XmbKLqZGzupdeLn+CxMN
dvUZcwQPp4argDe0LtgOpCoYcY+JeBdtXddpgB3fjeLErb4CVYxBL8s9Esgj
0sdNd9qY/2HkwPo6fUi9Tv3M7EIN0iGADch71TcbhRwRI9h4ydBbNZWI/xMS
R+i5BKMY9pfvI/0rqs0yJfovCWXlfd6oAJjIjvYr9nPRfkCkD6g3C//+rOAF
DfxDohmLin2/BEgEkq0INXGpj9RW8CUigiDrRCU2UCJOu67s/1oBiRnixNBt
mhpMuEQHIBqSYJLYY4D56zccrDWKN6SLjr8clcY+/ehY+KtHW5j/mNzy/cFG
x4V1oLashqI1tObjSOUcEi3K4iRIWKZHj/E4++quRj2NGNj01DRrCL+FpzJ+
aK5Sl31GM3F2bIX4jk+Ppu2l16HaDdT91ueSRd7Gpflf1gtATIs2qq0yMcWN
iou1dUSTwBaUN+If9MUTvb077biLFQIy65FNEZq7kXVbn2fd/J9dCK75ZZAg
PrBOKDQwh6mNlIAEp2F5aoAO5ymV1GdWxWPxUIKBTGKNmO/0YnpkmZTw1RQO
E45lYnFuwO/BE1XVBqdTyzf545Cv8y0gFAG1hSsbNk7wfWzuhxpCrBX9Rr3r
UPsEUk3mwPuvfbR/9i/JjfXICvRkVc5bN2dS/4Upxcpj8qBCU4R1Z1uIFppI
MJkwVC2hijSjrvH/zS1EUXbshXS2KJ5Qkg6wM2ahel3y/Ul4ojgfoEiREedz
hke6csUkqwJvZfKGMBAAI0Zh4CMz1M8dijn+EVWivgFFzRwKQrFHPAo4DIn7
6HMTSK1pr8quZONoAQ2Cv47JQGgLF0jT9VtbV62H/9tV24tmP3FBx6B5iUPH
S3dUw/Q9tfoHm3cM0viPNzm/nFlcQj6QqEfGYsblgVTPwobmiCAmFECR22NZ
qjKFEJHvHUhWbdMw0IqUqmRGR8tsIx8SBI8i+qcC220DbFunPolSXXzUS/QF
wY0u4W2fwovBZtokCM3dz9hKTdPHRSG2opaorc8wEvqnyce/ic4hDJZ7kDdy
YUrcdMYziC5z+/1UKjj+E3HDHAjgYY52Wyh+BI58LKED6IymO7WZafAdEPrV
yGbbtBal20/UpwVOE+5GMq3Olju5xeYiKq1t2f6+NL8z3myfhDQiUeB3oao0
+/lz2QWa1/LcC7QDEaQtUMb/7YntJB31LfFRKQNyuRQI7c4d6CTonXrbeqYx
hdSBxC3myavXQH//TnX9QRN/4GqFkAe3Ly0tP6LOxPhht63dwJQn7dTcCl5o
JdbCb6O2HZyLthFg94bZ18DiLYAstfnI9aQ0OPrO4D7URMgq+QhZmILrY/aZ
58IQje0eJghHbnIDA+hNRR3xEzwjY85VoYkTUBcXJ4xWYqWLdZYx/RDcwLVy
TSzuT7MjtRUuUwdEeuVQ2/al8zEMyY2XqY5JrmNaOuGohAcTeASm+RPPvW3D
CGDoXNWt0+nSHGHSULkujFkGZC8eDZbCWdGSgSi11s06RFJy2pphnFZ76aht
FRjhxgczGY+2UWXjA76nTZVZghe5dPrqu94FcuIX1i1M9la+wqkh1JW7ejb0
tdzU66Cfx0CuKeGcbV3ja6CWnuTTwWfjLIXzwMbBb2SEBwWCQjPjdoDsj3LA
rdYPzFuEmKtYB95zTUdxPpQjU3w3Wg3OcaQXQplYwHHSYOGMyy5D44qhxS8a
+vbZphDn3T57Z1azFLugFug++E0nsumZs3ZB+eo9FK00+4TofcGIw9ZewXzl
F/k4Z4JV1IVuaCJhRydiOfhwZOpB9sVjMppvmtM1l9tPM853olKRy5dGEsbA
GA5Zk3/n55mUtHzWdTKOePftWzQkNsPNfOQGEYD1zEyzJoLMlRdMp2wFHB6V
VO3NRaD1wjbPsdXh8gGs+M84+Ze2rx8nZLE14PcooTyzZdFEJE+gwiPXRUWI
juTN8Shd7Dsb3ys7SmkvmDGXt2/wilzgcwDFCj/HCFFkOlJtUAZZQc2xGwxw
jIIvaO9T6jPup2RkYq5YjxGtqw+fk3q4YMtdHKkgwqy9xgWe7sYsOZN15Xtg
ysTsUdnkjgedNLiG6A0vY9fRWbQ+8kkeg1naVpfmZJjw0mF2NAB/yFIe0WOu
7csm/02veqsLvv4GjvpIqccrc7x6mdr9k7Z5q0IxDiUnTfv8pATzXoq+DPUO
xPULGyPRfK3gsjPJvLharBkqegVFHSBi1nOdL8UCx+bDeRC3Hw7nW0S72Zaa
3O5rwH9PORHo7frL0Zf1JU8rIHjwe/bICir1w3DHTFyXszg5liqCY7dfKY/p
h+n4HCRzEMG+uKNEBwCx1k9YOZgNkobcuIT9Q6baP8+bOlhcRNcTfw+VifnJ
EcHkvLoy2AOg4Jhj7ksG6yaTjFXrF0FyO9pchJ9sk4AAlH6vs5RruhrH5I6Z
2c4yohB03vqJH/pnUO4PxlGK4QtTfxvzeBchXPXUeZmckPIvb3rVAO8NrMn9
Q2sv2WAgzS3LRbJR6Gmui/Hxwv7Sih5n/nogccwfRHWde+VmFQBjtSti5J6q
FGQ574TL2yAKCizvPbZjrIW4u0uoZPcnr/1lTAelrOAqowWYi2tQ+eyGX7Q8
MiyHBY4T6sm31RPIEfBDWLwOyMBRhH56L44DAWy3Ibkv/8JhxtgPT+iPiCch
GzCZSbuE9MgNEul/1YA3uSoeC8gjf57EMcCUGoXeJt+bH+uG+SJwUdxebGGE
oOoTAFM65oFkyX3+xWDHr0tAxpNXAuKa+TiMWPg1YAI8dKTgfhR2NTpC2DG9
HpsA1aPFsKyeeE24SbtN2bUGhgmujhtI3hf9pMv5EiPMhaV4qgFZ4clvfhKz
/92iC10AKVnXVk8c+yIt1nb654jU6YeETm02VhAepfQ4t13hS/T3QHozwil+
eI3X08fA3TyS6rafei4nso9CdlQ4RIy0/1+FQS5n360p/HAxnhIYdYukZxu5
DliB/XubiS0BHbCHUQzxGnhvryt55qxwqNUCPASphCgwTp7XhjNWz6ETnzh4
TZNpE1/AjF17sMURMnmEdv0yDIY6lgFAuIrA3CHgM6sFNCwqoblQNiGN3mHW
wMgHo4DqvNFNm05RX2ogEyK3p85l+gB2YJe/remvSFevTlVq0N9UyzTBXZSY
27Vvic79n1Sb5hz8Kj2YatvoaD05EvK46zs2QIZiubBzNqc2wAvMoOwEoEP2
lj7bF9/4C3CaIrtz7qeGrfxwC1KHyihHYZGan9/yrzWxJ9pUV3NTzYwzk6Un
G9yz7nrsSLQDOc/SOv5WRojVSC+Vq08LTGMXQoVpSbMrNxQ20Wr3gQCnfAEk
sk275LxPjuZP2EWh/1GFmwCsou5wwLJvSIeagDZ67J/U344sM9qoLHdEZ8yk
0A6erdDlukXWX94+ziH7EguRRalyILDYWSvmlKa1GcDIyNP58TnECPJr0YsB
gD194pLqdWnC/BdPHQGvkKAmiCcWbQNf85RJowyn9qlSPBDjrM/ISYIKj70q
BvO0UTfroAcbU19Fol9S3a2rj8AkyyLB7xgICh2nUkyGHhWq1Pu/sy3f3LCa
gQskRYmRqw8+fDivzQocBg/7y7DJTlBCjKjvRzsnxMjz/xuB8wr+mxGbcAKW
UoUpg9f8hsMRBPpTvkMPsp++8/gS6bEvWyNX+7vxoyAuSeyejdbVC8SjT1o/
6Zlf/HfqVG05RaQw3riuqAYFDiFTeMN3CYlOhGsFECDGGsf3uozbyzcKdhYg
HtKh8dTGNTBNluXP4GMyChxCHgULykA3Z5Xam3aDENSyfn2ViAx1aSHWGJbJ
1w/IMiEMaP0Jd11nakV3k/d19Tumgyc2eqjIntFS0Kfs8wLqD6keuUEBXvxg
5ZBGA4XkxZWbs5vLMRPS5WASgyt6P/C+VM4gsWHmd4qUuBrwF86uV453aHJu
69/No1nsWF9PRC2UIhFBNmdr5Fci9PZ5j9TqLuU64ygfzB+1sbr8ocB23Z7u
7KYsCM9ECgwVnzURvP0t+Wu3zBY8k2h3RkMaJQrXCm81pdr5ROd/IjfqCJa8
mUVHxq1rW05jh1aEKlVTDSFNb55kGVir3w+htNf1NXIFfQwIfstg3d2TgA62
spN3lMrwXuizLK6zUjDiozK9haQxgb531aBpeIWrctUVrpibawyR5q6E0Byi
nDcxo5GzhH+fTINju3Rr/EhvCtHqnPKz1zXkbOk4TIk3eScR1D++Vw7TaYSV
wIm0+UQJ/1A1sribwfuhBCtsUPjyYVnS1peJB2sbC3Nyxpq4zlVic8Tir4tR
MnIsdD8XTDZw4Ii4ab1aqwXmU0wHiRnRbszTA/sBqfClfouCppJy9Ed9SJUr
uMlHf2h9UusMiYSjRkV93N1oL/vsG1CF6xSNDwsCnkU9tfTwrGlEjs13eDJN
yrRLtxNP5sX3zD3O0KzbogLs1jB1yfhXjiRzyxaqDHHNfN0+oeya9ShYzxEA
DTLbfVaMDCVTkKg0rAnJ/pw7kSLqA8ANqcUG9GB+xKDZYZDRXSw2k7t6PZDf
+G22+44L5CgDqO+PfserOTl0s9FGKs+K6uLPwAYUj3CY8I86coLcRooV7BoU
Pq5GLlchbk+hTZ8c3L+n9LpT3scTDtqDigrK2GLXCrxGtrUgUKWECWNnrCZ9
rLGL/ZHGbV/SVsVTPEbfigO8QCRsd30UaAiiAri17BCRh5E/dgth8uVTWSwa
QrEj71dyZbKv+u+/Ol8n6QO5GNgvOuiS5Ggke4D9ZjOcqUBLdSDxtHZJjfof
qGteiEsRdh22Dwcq0RltL9EFvcgSkmdTunPICTeYUCaXIbwcHLlS5wzHFQ4c
KCnWj9bLNpB5REzxJfHEgXVDSYRWUBNVI9GQioLNnKNgCxNb0ptXhxl2pSP/
HaZOJmZyi3IbLCdSl50PlSFkKKFVp19uTqO/6qdYzOUJgstvvB0imDgT0lCn
UpaeYqkRc7u2PoM9ENLydPa4M75Pq6VwIRVKiA8Nh8hEBMvs/2FzuYZLdaD6
hi+3oWUlmJupEygtNyYlHuG4VUp5QTrUWDzLW+RLq9iRnXHpvXIl6PharkfU
NuPIj8ub90U3egr//tTdzIKm/B6kY5OABv0OV9EnIZpacqE8Wjqeg59Z5vLV
es+f2sGsrfkjIjGoe/59mMH2dCkOhdRRYdHzKwNTb7gSuynb9zMSmFRRH5K+
Wr/2vUjJbKl2JAyVuo+J+V+AH2XCmv9RdHxgUTMgB/3nqZTQLZg5KqZuUSYP
zIxsZBQhlx40YZ8s1sUn4xBAQduPSWHXTOzwSe1HOfOxXhPmv0UswW0hgG3W
l5l9g5BGrZKbwXFth5cRqbryso8HbxMQFhm8Pk94tI4VKJHk4R2yr2+uVvQL
HiJI5hoGjsqRPLyWHwNIJWy2Es16w5+xZsDEiliAh+kucaAion2yZDMAoHDx
5SRqZSrQm8einFJThAF2LuSyxqo1SYkE6SWTDnhuKAWTM+2ckSmQE5rdJEeA
Tl3XsDk94EoQwGup6lHn2KYQtnczfmDn+24ychQcu2EIUN7v/USUXaNqR0qz
sNXJ9Isuf9NxkT0U11W+MAtjdUX6O8FkCrKu47gm/KEEDkkhNJtWJ23nEuP0
11mLKBnIMny7YreXuBqdTUN6OCWI8iab0OoiArwQqfXPNn8Flm5zOentmaiY
gPOyMPFxgYz0jyTWl6b13TyLov7vxOU66ECIbdcBbSp4s4JbBQEymtifQRij
ypa3ARN4//buqfn9UeG2fW6FKAXxbcyHWA8doLzuC4PeWhFgPB4sDDLbqueJ
XGfTDBQEcmaU4HThN7Nzggquu7oHgoOK+YCkxSq56hoiEJ0orp/KACGAyRuU
6g6QQetIJWFdcg0PM2zMQ240rc6aYwaxHpLgE9pOQeP3AlXlkUgqtcsa8VXb
B6xG4nyd4eoKj9s2S4FyVNW1gzfPnd8p2ZR0bNsVjVC7Zeo7VAmbNLVtZhGj
46X6cMUFmENgY0Ac5gFWqkIsw+fa+sxfs5xxYPLiBsCozSw4gBGmjYSAnyRM
zcC64UWS9K4xQq9YF6EE76nxDMnzizZXh7a8BnbRmEaYLtZ2RF3etARQA7Q5
hYwVBtLPPZNHySrKRgXYXpCGquqQfpixBb40U9qdVjt4F6IJ1gd8EPwLNN01
VmOKqSBi1uLMUB8X7ZWUzWRR7W6eiXFtcEc6ZTokZgTcQ8Xq89gYMvJ3lGBl
ptGMhFiDwU7EHylgheq2bzNaDRip4F75S+t/xHCjPwe80a5qcxyLpbPniT8N
OT0VDG/MOZZZQz+TgKH4uBR8H6Fup3Lr3MEY0Vxnm0WDfmM623jo19ndrojz
MDjaPJnB7YOukhoulpawv/WnnakHSZmjT4R/lXnveWNbPFYtHsFzy+47taLb
MhUeUa+pLupV6dJ+pPcc6JF7YTduzEskrWHpxir95kbcVj0vOD2DkN5FA+dr
GNBpaFrUnZVEDre0yFAt1xVNpCGPZduO6prPvBnS71IxwTWJAjQf/xDNC4EG
IUR72cA8wm7H9NA7z98nACEpkTXonDMeFvgXLToPoJjMCjtqdNBGM/el7o6o
X2NM99mHXpixkGxMU0jTToCtPQgxMG1PrjEkvV+KjBcAMn9fJ+o8x/4iso/j
/+gE7YEm0JGn1GdPepWo7ttuTR4/Yu2dxfx5OU4Jjftsim5v4sF4MbVgaF2X
y8Xmj2+QDM7gY5wSh1DEIHdfJmjdXz3qPt5K71wmLMnGtAe05yeAFpBp1qLM
0JBT8ktRudkrXSnv/GNHGgIaR87nMVp3fkBx6M/J0ZBl428PJi7/JawHzBIN
uWOluCgPwwhSxkdqb6gKW+Urx8K0p4kruRd1QGnUrA+SY4QO8tXHQFDRv5pX
cs104kPuUoNK4tei7WqPAUcQIYO6d7Zs2qFxYG7MKKlYggl6Ws2lEUDv6Mm4
Kk+eXohlki9sjA6NAWcHuKWkyfutg4H7VNl1zfqrN7ZBTeWkTWOM9G9SvjyC
Kl3XNx5e8JRCNApxtP/JoXXNmS/789BI9bw1qC/wp0QVmSyVaZRBnE5mnZEa
nOE4kMCW2zfum5lb4OJ16ZJPn0lrnnNmS20raR4hai2tjyhEXNNEXELHJYQ+
Qwimu2HF2ZltebZ4ozN7Bo6C/UEbsAo+A+bVaO/L9uvIraftv7SD7H9F1e5n
HCdcMhRbPP0JenvikEDiGku2hBPvhQPYZlJkF6WafMrZCQ2ur+peBipTeYTX
Gzn0Z1F82C9KvAMfcuEWUDK6jIa3XKUiLjiPwzWBifkdp7oXmslTV8fQFbwm
RwfwUy47BHVzrS1jABAto6rfbKY01x8LwrZFx+RhNJ9mNms5InbyBO4vW3oK
/yV+qyyDVAgy1dE08c/oWai2564bNOvY8vzaV7TpLTJLLHu99aThDt35IuNW
G5QNmPMQzKXh3vO+xVoGTIbnCsxEwntlHcCYepRj75+gIglnbxvrzwrhImXm
NSuiHI50WAXcz99eCSlN5VJJTT4LnQgSSQ1xGT1CfezYtxR5qN0goSjEHx9+
zyYhvu9qRPAOHmEMcKjCD1ZLGWnGYMH1gOggH5S2FuIf0Bfw7SWRfxZRLljp
/UzXaOBYlvDY1DT/xR3pcLuNZ/jgL6XtkJ/0WiYal8+5gxnNSpr6r2ZGeT40
uxphmvokyDTzKlzAATgbz2exXgDWxY1Ou68gEewZg3+bzhn6FYVI0RNeUCYZ
LzKYHkuRDoJyayXeTTBmrLkNi72RuPSZEIOSSEBAzWKLiCq5xifb9UBphO93
FmrglAOhKV+oX5ALsM0uT0uaEGFyri/tSQzPLbmtJCjLAWGF7DJ4RUgarZPI
osddPdTCrciTrQnK0SfeW2MkKX0/W7U76YPok6pDLLKSK2BdDwzzfg8gvxpB
ucewLeJHG7DKLrepg415e86dPEamiNVRUwXLULamLZNTQPfjJM/87IfvCQup
QOcskcJ9mJm0j9qXv5SqHAUW7Qof3yEGs3CYvVezRdkzJggBRK1SBV+c1fC5
HiZeIzf0eWyk9dCNzsofDtTwIdllfyMSP4H+z5Y3vsiNDVVT5+qSaFd0X6Bn
H5mQTWstZbT3N+MYvhWnHU3N3uh4on78arBqhEbODmWXSXXPMErcs9zpecFn
SMyTEKiXwxLobaqdOcorY/j/gYerQ/YUz0th0eA40wNw8fxJA8MaRzXkZbc4
LTQFBU531ih0kgm2LGQDkEwSWgjq3zIFAkh2BM8hY02RgX1uaqe9PzCPCg9h
uW0dJ+957kcJI9Autak1tZspppo2Bpy7XcKyiX4looJfdo+tMK9n+JtH7OFf
aG7hwklQa3ddedAceswic1fvt1laVoJL3CRMtpzblKUe9ANaJCveDgKLQu0M
xpTA4IOJsOk7h+hunwn0w9b3OeE04BRHPOOWHqzp7brOyY5z7q/VhZaOavoF
IqEohx2Y/snscDGQXjuw6nsHQoxGd5NWtONvPGHvy09wlpS9VXWRKua6ajQk
KNGDFAIQXAEldnbWxhfaTgXsln0pS7TQP9LkNGavxFsvt4FeELfQr+Newvdi
BBONptTCQAeyl7MlaKDBbd80DF/z2sH+F435azJYl1bF8anFkHDsPusWjfY0
d8m6qh6Q3Vp5NTcqjLHn+zzqbfcW75aUztSJMH+tbDNmusK9HtTop5w8oA+s
80VdY93WpjmShta7LS/OajRI3ntSUHOsv4Zcb4kdGF21kGuaNISxY575dgLL
g9CrfEYqciPyWjjHbKIglnz53FVW9LZPvP0XaCEKxo9zt7cPF2OsqkzAQpF5
S2H/+Irk23MwjyofutxoDnKEOKJ6QfyRhwAQCnZIttd2VA5hTOhMIDaymXIZ
b37dyN8HIIFpaTCikcpg9v/+mHTMNwFTqbqPI/dIAekufm3jQI1uNEq8RgKJ
ogTuXnYkUXCKRiEAhQrAQeP3hTeXXULYI9caovuGOzJx4OFtI2zRUcD4dOiE
Wvudj/sPDI9+8pkpnBFaAHq3jD3ZFx5F4FnTCHE3zJFGrVWZ8pe1geDVCyl9
ia4BPuq9iu2TmcHzuFDfwf5HegR8iJKloeLO5ApeYLJMOd2oZ3qOJsB36+pV
zBBxUVCO9xpEtVep75HUNMe2iCDJF5D5Wj2039tmjmMBPh96S3BXGeQqHM6r
eU6Gn9so2Kl3+XORYxZhWvVKoTxSol7K6vupZAV9NkfEKL90CnSjVtlvYzxH
V+Mu/6SRDAV6XUySdoSZw3+YRa1WTJgiRzMWQROiogWvwPo/R+d5IFnH2i7m
uTxYGhLd/IL2zGJUjZvbBSZkmJ9MICWkk5E4UayTksPvH6yvhmo0zY0PVmMk
2PHMdz2cLJdTQ+sIAnor69JRciFDtJOv9y6lbaqptZUP4doiZAeWA7y2PWf/
IDWQd7HHmEPtNBKqSKMclFipTMrGto0Gdu9j1AOb2UDGp/gtOqwd1nzl9/Y+
Gh1ofnmvcCBpK48fpCwZ/G2zccW8z88caUEo/ZFQAuTSE2EHVikg/Gu3d6jU
LzRk5zKY690ZCzGWphzVBXnOSQIVlXVILk9cEnbfG1ZkQUXYV5/ZOVHp8lEh
vI8tO6D52ypYKRdaKyjBadsHhWbv05mLSlcU5i2KouNeFTtGRjh+K/0ks4aT
fzGoZTVo64vKlRFxc/qcxIgsBuCm5ByQHAQ8Tgduzb5E1tAgP0Yi2+IKktC/
B6G31MehgAtfukMRNZtTTnDTLH9XhlErEpPNTJIb2uJf1VodN0UDuSCpusAJ
g0d4CnbI/IADZPo39b/2u3VyrPSg2o12FWlkLHYudngXL43SrzPPjTylD3gZ
QKVy45h2sP12zWQaV2ORGKYDYKYE0LGCatUNLl/WsTtgumF945hpuaza6dMF
vD7HViH45qb1YZr0OCzfZ/hMc17pvfHgxtLjjTaBgalYaSnDZg+i0xhxt4lV
f1wop5dXPpahwR+9nSPecDLVWkFVHVd1WgIlKFFA35A+Zy7IDCU/aHMxYEId
bExp6hSccGZ5dHlRQBLNrhRLVkCWD5jF+IXZEh3cIoXove5NoiFZkvASCaPE
L1uTXNwvSEVLGdqkhEz0DbTSDA7wBWY5R7ClNdRAbbNLpKwFLBsUxfAR3Xyf
S60hnQXK8PpU2TugeNKfvI8Yqi3siGyO12jLrANUID9w+K/Tb/xcFB2tFdBn
/EI1WL+sasod6sQlRwmw3aswAylk2+F24zaP+Uuv788QkW1Pweq5jQQGVZbe
6MFglG10jceLVlsHR56KRVPt+IAKvQzJ6osZLlwrxHog0BhRKB6W4xtU3Pxp
p4MRI4/5c8criSrKuL4YpDoeRnCBR8886is32z9LGM5t8Vm4j0vUshHLW5A+
MZLVBUJU2A5o2sjS8Xa6jTzqn3oTuxd00GWQjR/PAsEE9TquJDTmncxb6/lz
1bfgWi4W4ar94itSknBNfbsLqC88nIvaKoJ/UmytyDDJd8t0Vdx1ljI5a89g
sXDrct342FRhOueDxML6mZ3L8A7Ta3dytxmsYNV9o0W7ItS8Fhs9U1dWW2A6
3jjwUESUxUZcFGJxOYdrQ/e9gPfZ40wg5Eysp5W2DwhEh9rO2m3o+2P2tseM
w9S7ps11ZyrgT4dFXYTwlVm9U+6WInpogCR0TtAavHMpMoZlm9ea2C9LCZx6
ctRjihq1YqqiFXl3TV9gHlHBmvoUwAu0LsWPTTypbJFNpnL2QQWrLsKZNC4V
aLItBBvdCdAQSCgKscOD7DjYqfOABHks/evCX0Zat9rMt7olbUM6IaXhnHFe
4tTv0j/pDaNhyqq82eDmXdXfrlLxxARVYxjpwJuvFFQMTXja1PbX+jnqMkzi
SEKhkq97I4YllJTVCacudVsFVFHB2TuZ7Qu2ADSQCgQiopxDr6kxWWAwnp4k
2mMGgAn2R/inX/9Hqn5LnJvJpdKibataD/A1JOgKAJ1PzcvxhylttRhB82+F
oqFPAxD2lcZRdqJOlx+fblVh8TBo0ybr4nqIXieLlaqh39uhQfONZFMzOet+
n03KQ+Q5yi1CoiuVxzQB7WwoR6Qy7L4InL1t7yY4USau7hNvTalPe+NMJulr
h7FAwZvX6tfAxO1MvahDRsxndUp8D7t+wujxGw6icBP466dvoz9NyfndV7P3
RtvOx8KyJn5k+2njZCbSrdBqe5IiNoHmvwVdbEIkolMdDjre61JkzWOAEW/M
eYHVsmNPlzwl3x6rPPnZoixY+9lvbhJeVdnumjwyi6vGe5pYlH1+Zeb2hSpf
hDqlPslnaD0bZNvnlDO8Q0LSQOfW7UBacHo/sCqdzyINfHll0pD3zg5pZyBG
qp/CAJPtVuTPBrkap+BB6Nqpw8j560kPW8rATJt8WirpXkbCMP/Fsuy3wOUU
GUp2GNdtZAUOPq1/VVW6den3uQvD/JNnQU3zfPTC++0uf1hzbUwos5W82huP
80cztvGavfQxpn5MsKSj0TzI2xZGK1wdt8DsudktnR/6NUe9X/YkJwguCZg5
zzOk/8NR2Vg5b598or0J+4IO79XcLo1aTVW8xOvXqTU+JMCYLVhFHbA/t3nS
uh3hcFRn7dmu4gy+aV7qLz+4t6ERmBod0wnlc3pZPPR/FNuiqm+OZRsmNuzX
Ne3muekEU4OZvD1vDHt+K3+A7nBdpTIJTpJ/jv4kd3si6u9Z975YeHtlZWoO
usXV8BvKnAg261vCrfIWk5AVS7xQ3Hj/JGS7ISYowc6Al+VueRbo2L2MJUUf
EQAfu+HaJ+JdsL4wlGkKpyIpYWNdrM5BEnVWVtPqY8HpVAO5evHjfPank2Zq
CQmSS4udZs40daQ5RFpUUJUmmE4HwPL5NttnSxgyTcJlJeLq3Cb9eO/N9gQt
9f2a5EyDwraB5sah808gLO5MRShbz9rkKtTIdDBa4kQA3d2nbHaXgQlOvQFG
2nmL2AU8FBTWV0tciE09NHosFcss1LXLr5imWIEl4GC4Az0JU17IpmCloCBS
2GlttcHqc0HOmeJAG1b6pzH+dH1WBPh5Cn2yJn7EUEUDehaEXLbtvdo+8Jp9
Ah3rj3ZHrpoLiGhJ4yvRzcRommZF13BmqcTOkyjfScLl8gjxpPL92mgcJtL/
FiqvSutmLB/H6u7oPuHVAQp0VZmtJIAkXz409/353PEIhEoqLg4XWfoxDqU9
wdeVJJyRcwoLOyYtgXQULtsXaB2QWdCDiLMrlxsaqvjINwNftWyCmv/UNxce
7HeRJzlFiVb4u5psgjgyA2In94mRwkSE60KVuN5L3SG3BZI2kHNSe4mXoV4Z
TYdwZGsWndo7D+X9ziDS10j7oLuhMXgtzy3sCdTh7SBEWGEOcUv7aLyaUbMq
HdvfJBb9R/OyiK7IcH20a9h801xKx0sUlIsPO5/fUmm9dU4K5fejWQM1Ez6C
8az1b87l4euo8q/mh2Deqn8jBftDeUEinDnmBN2K5zYJsQHg7s6578g4T/Dm
/PLoVMnPU4OpmEeWPYXSzI5PYDaHVOTChYEg/Xpp3grGFi7tVYg3h282xESv
e0sAfiiwnba7X40eKpFkUFr+1UCUJwkteEQjdGTqwUEhflQj1U0xyLBkUhql
Y+vPDp/GrG/mbjGXsB9DOhwyILAU3U/Ph8REh4ZyvBPW+Zr2CHuSPwQ5qm71
ar4SJfPNVX6IvdicArylEOSznNS2es4SFytxDNjpuT3z2CXq5WCduYlnMtcS
r9eOsKlhhfVih3iR8b+JpjGEeMpB9KndYK7P4FyausGueKaQFwIiwB6c2SjJ
e+3W9TqvWsfO6gX+/Xl1xo8zCL4uxwRhoaOGLMqHuKZscEXjsygG6cd2ttln
VTIh4/VMMqMzezi+JbhrvBov2E8lnk+cQ/NXFjY6Jmk3g1Xs5NjI4Oe0q8zc
Y/DURWkiUbL5uBLm9QuHr5VtpIaQiWgobG/N46CUO13Q0qDUwLo1PyYq5U0l
X0hFaZuPu6s5cPuGhZDEKM+EVcgwLrt0QE0HJsnBkhn43kjlo5f/0lKSzkUD
sUu6JlDTSx6yrqWxzLsOOUlLC2WIfGNmvvJQJLOnvP7YYEV0c4sKF1u3PljJ
/lXFlzx9NXs27AUO51QAiToaLBDrin7RWqdW8Ml95vY/j/ajgWJN39xJlmyJ
rYPARpmNihb4xbXZmM4L4bQMS6siLEQW05RGc1ud38Aod5DPDRZXJzdZmKAr
fkB1HBbGRf/lU5M7iL25WYMIN8phODeM7A/eoDFNN14P8NE9RPOBcdeYfnqC
dxjYQ5mh1U0Cy1Vmn63MXhsQwDYpR4wSbbmkbOwWD3HH/R3glMIzuHvqSNkx
4HCGSnUWdkuMHJogCZdVkDtK06N7tho4Ri9T45LIBsc++m/fixMIEMmeNhc4
pcJZvvHAkH5JKAm6AW6JVVTGz7JMnFS9L/jtTrlrrlacO6USZOSf2zY/WTiG
m2LenXFLy/MkhxQ9cdWUWx927Be1M6lq+kOebmrOWnp/sVtQ1q81q4PjNISy
bW8yoq9xBwEqgcSuS/GRL4H7Q5ynz+c+O61gMG0PxRvIYdBmvhGDB7Wqgl0a
3I1t+j9vMGYLJcEBB91I7eyWMm4KDnCJpY7m9iBJ0CAwkaIexqS9xLbQ37pg
X5leEvHkjYPi8yES6ZHtq7E2Y7ASs4o2XJrMLf7cZgG2H4Nn11OLhaE1gisE
+t58KXnISu6U5jC8YG3WHhSsKtmcxAyCY9R3mvFunQA/NvjyJ0uIvXoTFsTo
bd6CTrru0SX2I11Fk5c4QLW2+HaX+keC2IWFeK8w17YrKG2+zTKJSPBSobs1
QE1xdKFVxRtYHU8Ff+sx/M28Ir9Fp0Hr0n8sUivyRtFWQ2+14TaMw+CVFw+b
msYbbc8tXMzDFrEKZQz1XprxCNhi6EayOX+1atflsNN0sJF0QpjL2pzn8Yj5
wszWntxKX2ZtKha8d29kwDaAqiMTTQH6djtoloJroFEHeKDiQuyIwtdg1CY9
WcT2OZ7gG0GcVErRaKqGy6KgMJMjDrQjOHstU3JO5S/jYV64kZo414NVbXfM
nb7P7on5F6i4K5VOf//WbzlzI5YD8H8AN0plJzqtN3mwn+h8ZoHhbknGfeH2
YUi117C9r4xhJ/7m0hnF0PEBESq9qhFxN9TRdNwqYhCzD1t5v5UqflFpbHZ0
YGqpMw0WYjw5jyWFZJsg0MoxxeMljuFgNwZ/KrkiGhiZl8s1Ab+6KLFa9P3a
3JvBIVU8owN+hcAeoHXc8F3tpO8Lw02blIaBDKDbcQ/DDLTnosuKFsR+Nua6
zIX8aS9AXUriLPRWBLqzWnp7hzv1/EjZ9IKiyD+0OvkZu4e2HPTyTxl80AUE
FhTYCEJRRkWGCgKQoMk2BkYjCHfVi1bSce2Ji2lDixSeOPUuuGi9/HC+Kjlk
7w/T4D5DQ4//gCoJc9ZGXsBSjwxHEuxll/e33vd6MSS6VoSSDI9CEO+jVueL
zNwWhbhAqNbHe9VxXWl+SBqWgMIsv99zYktcKy+8tu7AcbgfGGYXSk2J+bz3
mZe5jHry0G1bHgYWYqH4LMr4rk6iMFhNJt1Fwn9N7mRaq4mjtRV4McyvKvRT
G+8pVUB7TZ1NOEv/R4FyVKTOO1Rfunul4+/Qo03icC2Ol4AQvnAG+jWuMv6D
0dj/8qOO/9sldXkmcsH3SqktRRRs/td+eKqdhDrhALS96+bUO3O0rCAwGlOB
P4HjO+7JOj5QnZ5aw4y5i4oIBKwb877bgUtmhyAGDtYyO/j5oZkRZxcgg2aa
g41SNtzsKxWKE68W6Ww2IzFMrSYoHnHkbT9O4V4Oc08p5jHvXWN7GoB9qaeJ
NU2JL2fRfp4FMlBjkZXEuN5Hbh6Z5ZEP59L9Kx2qBmuO2JdSIbCVO1k9ehs9
oVlRdl5pbFAKAKQQvvYJBeYP0fnGYdIaIXV1JRPdw2/6bcchg5aniAKb64Gi
RLTzZtddMfH1P3a0PEpelFRfaABdc3Tmz+wfi8tHvpnioEtQl43k/pTBbb9v
Ev2FHyGIIsMeMvtahtJ+0PbCgceJSmtnEcVfl9My9bDXVxAzm6cYo+Rdtz5g
mfOn5bwkY1EDp62wnKEd4BIRKj2dibs58cwIfDnj8fRAouOQ5UxIolC4fups
NLkldCh6MOEv0KZHl3+VJ44zj41ONa/E2X2DMn8fLkEBqpFAo8vlMhQHxavC
IoYDpbKwyBHNRZC3CBVQGMYTFS4vnYs4cKHuvyvSIMDiLLFNPpSQyBr0KafF
B23ER4fUv4xIrXh7DWKM7u0AO1tXAjOa5nn0WVAd0tYzhuIqu6CULeMzJ5hm
3YsdX9VWA4BdgQZbGLIRkfRbaEd6Bvs8sKFdj0lFW5ay040KUtuyRHRmJ7Cw
CH1dZV6cdC9xk2qAw4tUWNOm2diqGRomtTFS8ZgYrPLN512k6nlrqLC//3vb
FuokIfjQLw++GPt3KN8yL3Wmyl+weNwNgJrW0yWu9fjy1aVtf7zO43zaPMxg
ztd/fhLJQSl2eCuKRjOmyTJHMnYuh+nwjZve6xZ6ScL5kNtpa8La8yLUoT8t
Za3YCKFbhATD5ThJ+r64ZTeR5PA4w/pFoRaI7V35y9ZkxGCnt9xCFs1uAS28
GCwk0ZRnu9aE9Kt/A9kPWEuwCEvzT0RfQ9uSLD3MDzP/6z2hrzH/0m9JXkOo
1s+lenjm/w71gXbDEcnrJWvaoBZrnM52q+wzm6Wbr4+IcURCNDOhXinE6T+B
2BwuQyc04y+MuKWuNI2UzVCmd/2kRknfIoSaVzeZHW/rz0Mx/xkg6vLVpPpt
gUEsCgPF5PyQTPqP1wq8pfqmCxL4g1W8+Ae6x/HIaeWcfH3snHDUp3/8xY8J
e6h29Egtu5ULmwgIE9yflYsdfpk//sN166uKiamiy18CgYJm56WhccBMc9T5
undaz40Ak2bdQnjH1gFf8GwgNes4kqgXSin4tYByBwYwY30ZDABZjW1b3aYU
s0TP1encr6S0QT+wfx9Nn78kquk+31V3uI+yeRsQvC9XeMkblTZVszr6uKQq
/5Ss5z0fnYTLl0DOtR97NRACtItBU/TuQQClVD/Ia7ZHARzdMYbiZVUQVDLU
0xOYXORDJeMZ416NJLQ2u9mXxQkR+jSGs0KH2RvGswvSWTFhl+gHJHiYSDb8
9+EfNZ/3kiVDvHsWZ//92FoZnFrOUM+UA+nqLQYGe6BiBCCB5upQBok8yy6m
slTewag65kOffpitBO195FuPffDiiTJ3jRc7YLL8+M/QtMNwAiUPrGKnlwRW
NRoFMJglGWHT8dtvIqDYwg0ouQ79c7AZw+9UWzjOotvAeXZaumeMDHPN5IBs
Cwpj8eLNVJAGNXdY7dYFXNGoAyur512S+KRdr6p5ZR5YMQspt2heWAXcSvbx
gUjY379kfb551EUM31Gnx+J05uBe2yk4RioBcrviSzxtzmJ6HsWNtsZqQfiu
2tsIWJRpTC3syNvOF3IKMhQGf5BcSLwRC+svqeH6i00QZ3jcLD3erI0iiaf0
FhPBqGQn/1b0co183uMxLsYSGUPyIw94pwQb2/PC3KcCHCm2NEHjzTTiVSg4
l7BudnoYBWDXUaOYeLuIYEMhJ2xL/FNy+57m/i0BAek5eNqAOM+g7DSjtGRR
5rv7/YMa+TZGsMQVGB/om9TAtYf6RbaW/rY+vYeparCRAQW7ZLUqrGoM7Lve
34hUZFi2Qh+kx5pCj1zTgJCd02JaNqhfU2k/50j9v6YJyFCOvcVhVR8GhfXP
/Rs6Aw4Sp6TNH12z7hXJtgQlCArrv+KL9iHc8KP/f7RBLjJd83pDFD19r+56
e3G3p1/Edl4rfFbrXoiPHfS9LtiueLktgZdSrM4+/QMv590t6ptxN/99OlDP
sy6PRCa1fI53bPSsvg2jueGbeU6IhM4Vf0vqfoFd5bHugQlfQj10dC3Hl9oG
cWaWFkKXdnhe/32sHEpeK8Am2B/oSpOZoKPqX6FjF4EuDiOb+P/4XQhX6HAD
1iUk408Qx2B5XPIimi5qCjAMxhcjnGBXdzf+NuJoTkgb1pvPK2CJnjFZwiUW
xN8PVMcy28BWoVEvp7dkMGR/Z6doTUWFDvSD6BDCCXjpBZnXvim98nYHeeCF
JbJuDZ8ka/FmkX/HsBpo5eLlApZ001p8rsAhHBjoEczFxS33grCEEqstMo0j
VUSL7zqakiqlaDSRs8VtqAOqXAAsRgL7nRAlctHDZk8zqk195PRCyEl9V7Nj
PUUSiL2+1+43Z2DgFKy0gi3ls23gA10ZTb6LlRFumVZeXkRsmyXqiMloz/g6
vDdMvaWF9+h1MW9pSULFslk8j11fxxnE+1+4d8soVvowUKRaFy7mhAKnUNd6
ZpfksNGBY5jeRa/6eMXUR+oEn8d2JBX3OdBkK6lpLi4qBL78zwJwpjJdcV4C
CGRbeJnqP8RRUpNTJdacs/wlmxBThe5nOw5P14/04Pf90kM8WXsjoU04EGT0
KC0HdBq3SPbPw031Q6qWU5UkafYqmy4xRRX/yKLlOCu8pc04FnUD3vumgEH5
u8BBCxAxkKzQDDAlnxd7nUmoLCi8HDEYKtNv7uDhbt13oMIKvpbnFIB38KIF
LfkqmZrWpfyVRz7jWHaAYAPwmrAYAyzB3IWk/pUd66UUoyrXBox1cWxbPfAB
1M6pAU2dci57M8+bI1g8rFASzX6UILw2n98MZbjbfrE27a7nKVCRC1xJfz6U
dmEn97Yqqf6k/93XMW+8NDi03dnFOYQmGL+ciFu7CngfCgcrhKouHza75m4A
z0R9UwFGEqj3TAlPJ9qpn9lNWzR9DEzhNW+BbD4q51vS22eh9bYI+hAmsC+R
O5/3gytK5iP0UOSTuDl2sbl+l98HTA34F9nhev3UutckBEUke6P8yOenGQB3
hfTjbpM4MyJxvT68iP0KDOKoeAQ1FEr8sNCnisgYOfCZmWfvh7jIOQHJ8SB3
4cn+FjPKPuu6KlWqJt5P8G0brBClKGAyIgTSlL0jnECI3jU+bQCwCTWreq6I
UiUKsPfPiu6KfmC+W49xgEm163ai629yVMPZuJ/p1qCQ4kMWYdbwmsW3FGuO
JGtWVjvbtcQejFd5OrEg/kxn6XBvU8KX4DhtooS1W/aBawzHvmGTQsDlCC1q
+zCbioT0j94wF4B+Qs/w5zqCotz6ApWriFV0zWvGQwzvKbwvR4tN55U6mvpD
F8CpPJt3T/TMMbKGB86qMcrz8gw07/HXHBz3TF1YzyRpnMndBo+nPqO4Dxgj
sAFIO3I2sYZoMnhWxEmLMU1Qof7ThYHB6EBAIMiSw30zB4D87cOO6/COJ9It
4ljTV0Po+j9Pfq2NcZRg0CR6BqVV6fWRGKSOIm+O/cZ/6xCkROhe7sboKgdw
uyDt3Cqt+5BHka475dS+YCdWRKztQwwKi45+pgjjI5G+hEMtHswkstpQAuug
ABTwRV/h7PEzUTsgbpFZCaLShAQFcw7ngNwGQBrp8QJqi6PYbm7vmoVTS4WU
76ybNGhUBchMGzuEBZGWg0P8UnouTuEQM1ycCT7ICckTYehFBe5BR7PNxjG3
HdglxFQJdvA3DT5BMPN9eu13p4Ub9zxH6YViUyDKCVX2qA0uLkp7aj/LuTy0
tAvn22BzR9wdrSOvY8+eUrBW5GX5xRFcxNoMWOj/YW4aLb3yu+Jnp7ZdxBHW
4IygxUuVSAMQoiZFCLnZuZTCcaUpr2bX3PHZVrUieEvZ5yI18RfUxL0rjKC4
Hz1bUow9GBUXm5hguns4MzaGs8EvWxDgZCUDYoIUfH97PQykTRPVjVqptJvS
jlcYdWS05VvIpUT1l6ytw9FMYYaNemztmY2Acj+zT00vYG4TmOqC1/wdbbf0
LUR/VndNcFjz//HBm7b5xKJ8roNSaKer2hCudE940i5UuQgkMKRVtwQi3Vmd
yJET0A4GL+njzQa0IZlzvVsNI4NwSb4Eh+r/hh4fTlSAOtVt37tI1QibTW4K
+zyRMaWG9GFWCuDE4kZf79PGpBI/4ZOMVzLjEDxQvduO5qJmqRHrg4GUb3ID
KrXYFt/lAPLCD5oLY/Smx3jNRocLSwQlgJ8NoNzhtmZLGX2xBdFlUZqPQptM
0jFzm6ULrBUpniuBLSxaYgHBS96GrMv+DGlkB37xJ7H1PQVL4vmVmVYPaciI
BxcJMjBV/wbenmMyJr6NH8T5tAB9D+5j/ek5Ld0r6k8xRkwdlEHpUkckGu8k
d6Z4kracFDCsI+lHWgUKJXedRTDLSdBhf8ptlDgxWs7hLiEplkJHmvWYfTgQ
ItRiJT+Qoj32dqoKOT6YmdeBZxn39sMdk7CWPecEe3Dcw1F+TQWLtmNwO/wC
BbLEG4pwlkNJGWK+IBIzGOCK41IQh9D448SLJ+Bgg7ISsTwR+NFmjclfF9da
Fh7GviRsTpCFgQROz83KQNMNw52or2ocxm5+E9Lv47rVsP6KRvJG5CATmI3j
fgNK4UBFUVzGX0Wy6PpFEohrXw0ro46gKjmbILdYrQ99/DF6+8x4p+ExJQUT
tlJGw030qDNwGYvfXPdnSjjrX7ueNw7F8ERNdwo9RCUmG30lcdqW1kyPZ0Ya
w9Uk/Y/3Nor0RT+hQv90mHzrJWGiFyVmt5SObEX64YqdWWyiyWbJ/qAYP0Rs
E6wHPMtJe6gHbVxw0QCEcB6mn7lgXXyDwxhD0LdOwCY5L9QXVuVYRVYlZ9Y0
6SLsLM8k4Y44+PGY9dovuLYaJduXi9PYpEFNPJY/SO0Yc42m/cDHZk7uenky
fbuBKILaTOK7PXYXOAxoi4hCmBpwVmLw+uztpV/Cjxd/t5kgvWiba/+lxfm7
N0O18PPrceABFMW38dxOR+S0NXzvC+OaW8ziOjrygHzWJ2htLDG/2fu2TqNS
OYRli8vzo+7shHipcRHDviwsOdMNNAE6v2fd8CK6hjVxPR6IVQ/sBZtoMB1P
RrodlUcUyZjgdjecdjgg8ILsl4T2KyDqbc2kxsiB7eCd+jjrLDQKRRmlNUy6
hHc0VsUeXGv4kJ70x3JcTkTMDYja8vIzg3Y8IdW4KpT3qn7/J03ezdL/J5Gu
kOI9AeVXvn1AQnWji7rJOqKrAtJzTrg1YG8LWWLodNi6WRrrM4ZCyHGabnqe
1fUgGkyn+D1OxRCawKHsOoB0uvzhMl4aGnILefPYbzS8xUY8lp8Kd0ybqwD0
1kWGvznyuCcbaSkK1xuhhh23idbz25lRwUCVhPE/ZihdPTzkFP/SbF7/r73e
ctDEV20BOcLflo6BhQJw8hGExpxBzUSO1L3br7gbcQi7EhYX3OHPbjQhXm07
flVP6VK51y34Y/d7qp8sLWx06TgOTnVRAPD0oGgyBN4eBuaEeJPfzib2GUe5
0naJVH/j0E4IRgySfqjxAW/zefla8eIx4iwKBjbs0zW/7N8Xbh1v4n1xqgvH
Ygw00ZnK7j/Ei6Q8A7u0bWfMid5dl9mMcO6qO0ZVdSh2fqCoo/iITwL78X5Y
rEfspIbZ8A+jYmGOcmNjTEr2W9LIpY47hYE3GNP8yKPZ+Z1E0zcFuMdYIaAQ
inhpVEHH2gdENlu7Edi8NFHNejCNPiuZERn+jJ0UoWPvDoLD3558lTGGIcW4
q+nDzk2XIdjWG8hn2KzRZsg1M+3hZOtsiV1xHnM0FpiD79lLaPMV6sjtifVx
8NTqrbrsirE5d78cBmTg7E3FPxmMzXH/8OrAC7YiHoQViHuFkSyliUstNSGL
SOsk8bZQWpQWMvAiMs0vWk7YTzIbFbMmjOxxAe4Guc3xbiYoHluWEf+RyzTT
bR9/dLQD3il+JN0wyVa9huU8xRcPgW7M6e/4Ka9oqS/vqs5rcqy6ule7K22o
xCWw16vFjtDX/SdpBQ5UCAvKzp1jovVUAyhkYD9LnSioUX+bLgVlyr5L4Z3c
AKtO8tMGmFTAbXQEq9txYBN7lA4mH3gCynTLF11M0bMJZ0msIAkFcHgYYIke
byTPy2mHfEzN6C0bPdI6+3XTuQkL0gGtZ6vgudq4RVNsXt3S+luw4SRiW984
tPS/KXI2LKp+W7rNTYuQXPqHp3GD5t76hFnfzcJTCyq0o2/7E8McVMpN4vVw
Dh/suUMF305wuJTTW08qUKBK/kK1WYnK8+SRXxIH7Yz8AxHYh2fmtgnW/28L
VwXd6qbOHZWm8Rl3QcSZe/HHBZG0Y5oHh+ot1CwyTDuW+AqweMVTpZ87gxm8
H0TG2wfHU4uwhwnFQUEAc08tuTgDN/YzBkwRW6kDT+PYVGziz1RW5igrrA0L
qpBoq+PDJGes037j2L43+PoTGZLnin+IpeFvhvgBr7ddcgss6pmymU5S8JjE
oNJ5FEvlF1lVUpEUzOx5H9CNt7Dl9jQ5Kt2EQBPHIW6ZOYXnwPc2rhAtK5MG
M53PKM63xQb3EtymfZIHVYCKn6I9mwfBHmHpY2PIUn2bMAsj3rYgXvv/XKMx
oFAxVM7BRpyI7apF1lC4LRvyKzUZSmMKgaAdh6cJU1v+I28MyT20bgOKX8qO
guRai9en3oAqV2+GJpu07N0fcTeJczVEig1cgyZhvCe+Pkt/hPZTKreIVlmr
iBdSsq24aZ9srZu1KEl8+AQ4xksrMseT/v8dHoZhr76JjLdCGGUIdaR/8mfS
IEntvMYndYHT6sQRZ8myNh3ccBxoS9+A1ZKEsHaO8GVEtHakiUqEpYsNquCF
bM+4mIim8ThPIldSZEvo/scTMH33HcMoDCjZLHCVZeSnz57KgQrErC3GpBOz
xbJHnrOuKCh71Qh6gO/YPTxa9/X1n8gNwGwk6MwH5OOZBXZuiikZZ7v3dpJL
JpsMCPXumdXGUQO8sS77SRK+nYYCiIOv3t6lXAhsigM7kwjQPqUtWTtP6ixQ
JHnVff8gFRHbKjF2Dpa4/O4+OTHn6gNrUsEekLNQXGSd8Qinul47RnVisojK
cIlVseEvs6K7Y81DSKMGQ+YIRX/A3bw+BQs2uk+vUKWWnQMfhGUlgrNbX7Wi
vDiEO3A3RL2p5BcC+GOKci15JBggkJbB7eSWEdONH0j1XYN5TZHG3P0SxmJr
A/zFHucg11qXS1MmuHKDY3oNGPdCzU80TzFN3q8DfY0VZ4UgFFLtxTPbcsYU
KI29NmICmsuFWgsCMTALGpiQImDI2pelWvoVsZdeuA/hXYPqzY30LDWDOVM4
a/8lF90yWzmdMwzdDWKXCZs6VOncUBiorUzIlODISI3AkMxPvcxv6zjmdNtc
36orK4Yc65feCgsMLTWGdCv2pgxpjUb382rEIBcN1rw8rgdGMPLoCvPeS0hT
NsNMYSyBQ8i3+7E1HGyh9qmapdyxw86fbMbYD03qWDa0QwiHMy0X+RwgR+jn
psER9MbQfmMbTLjHyk1xjVJJPIbY4nLlHlClCU9jwyfBEL58a3PDcoN04v2r
sMfWeLvRZyFLeMiN3jJf1I+rb2JGDbkvLpGhkSryzMkB1oh4XzBuw46dpsRN
sJZ6rhDOv5bnIzrR8S2ZlBa1OorcnxrGdvhixS4w+AfqmrizC4e78Rrnkrp3
toa8NYHGHcV6wR8++YLQrFGkiZ6t7TjSkoCWIS5biH8G14EZo9MPv3XtjsGO
1jh9MaaFun1DQENfzwkzUz8xR5f/4QUkEoTm1j2FaJsYHmZDjpTo8gImNjRz
o47+Nd3Jnv0H1gzeG6/DgQ/BuZcCiAsJAZblp0+hgeGDlfadIR7xZSi3MpVj
/9lZ387qS6aYdp1tSIqRQe+ziiQN0fMiG6X9VQZRnCDloDZGaljhAThCGiO4
x/bZEeLZF+lbqnkxwAUi9LhxR0lg+o+Ef2ETY1Q7khRR5YFjJlGrvCVDkrIx
Q5eo138Kcq8TMEGd9QDdyZUdZE1bZjuzHq0mScrp4Q9B8VPDbsEJevbs2znH
lg5+/Az1QYwplhAxA7DmS76AXrM0XSvZURg2/twUJrNHMhAov5dZa4u+q1UT
WcSLlR0YUkl+r3v4byaOzHSG7/CBufY5RCshXWN7GBfo/eaIvCS9wNscvcV/
imLVrB+zy8PH98aqy2QeekX+WpL5Ow5CzqcvUvx2TFxoHqiE5RyvjkzeY8ro
0feLKbHWGlzUF/CmwNdbvl8Ehs1vIsaHzxwUmHR7yrJWV0Vpp0BqyNXl4mcL
l5Lh6azIv9wV0qp4RBUfEx8CmOyd9fIpzyuLQdYFHSSYgmvlJfYY/psg3ttr
RBl7/MCdn83WzetNhQmTkoSZJLdwlvxrrUk7CANhIEr+xkCpUq32q4T3UquO
a1natOyl3+m410SFVC3Tbvf9IY5RUrFGzd4YpfwrETqoA221di00jYWr/8qd
VlUUpUhZq2t4L6eBxkOPLKol2Bx2sUlRCVhGgNtDHC/rAxl/dBt5+GJPPXSL
kEwvzFK9PVu0evM/2BX40iqGng3mgRSavNY/o8vMhLavBbN5Y48wgxfrLdks
GFpLyBtYEOuAtiQOm+WCOL/qGh8Ki4GgxfAtocFH2u4zUy6ZHuUCF4fuIEe3
3ef0NgINqlurg/m9axM/189W/mC2sxeD8NV0lNbQiwRBTqHWHpCv/dtpTwsm
s9atDO+yr8I3h0FBMg5hgrcLYnVaBYpd53sYSX4nfz19r1XVVQ+uRQNwnftz
pjhIguKwHtoCtehX+AllH04zvessu2S+utAEcmsihl39Tw/nK7Z01lBvZ9aO
K25+S6Hh5qseTTxl+aUtyOE0GQHOaYMkbl9j9jaYR7vOFiY914zzQmKP6VDA
Fe9gTcKH26QdEoocN52XBd3spToySA/jTupmJqZj7O/raxKQu/Ba+VEjNrrU
xQsHMVeNL09SujIppmkjQhvA8JXEi8BbsVyn1fhv2HRmcznWKWsqd+2Pvm3e
C1R9PFUK3aG/m0G8TVXUjXxYtznZq+tuqm+BA1vUz6KZzERraBTEYEVUuic0
WvuYR83rARpqOQCn3qU5rYCrYgNLrPFvt9Blep6hIP4acU/PvLC/XKp6OcA6
zHVh449PgVYb1fIRluFjiU+62sjrABAoX4M6ZjsfBrTYhawaDuCyEhCghjGM
ameCT4NzgQeFmP5sGN3npHZRl82ncDwJdISSzI4+azdFrDKxfCQZStRuHCKK
jAmQ/TCqPQO21quOOJgMX1X73ljKr7Ym0gK/q9LNgdpKRUXlJG8SrCid9rjp
TbKFn30xMX6V0IOb31m8YFY0HOHSx/XhcXBmssRhRa6vUE0HayHa87YLzdI3
nuUFEnICd3j9x/Q41ISGWgAu5B9US53+9W2H5iIrG3OFYmBcBCxRX+VYCKNk
qJMU/riL/DftYzy2WHy5MbbsOD26dtehhUgmPKf86zlMeMtrKgKaYmDhjW8t
rWrQvMnMjpEBkWCV36NbGpgxxW9/MQG3oXVYHcgcuZIcc0/jQ7ssfhac8bT5
FtBYzWdMLccUqogbFFqgOAYnBpJ+rPn4F4rlrkoGpdBeowz1VxX5ic0w+xMK
BJmWAxmwMW3PmJDHiE792IDjKP2R49ioYR1CmpB6cDpEch3nT+CzKlECL8Nc
IFe55CyIOIYSKuIZ5AzMtKMvmof91Bug4BF+9obJxyFKHoHQ15oEd3U++zPU
7MLCCvnFkE2fD3pAnEbqLzGoyy2jw/Ij81nqyOdj/vZ9GuVtyt/UJTZWYzjZ
ZvJZT49LWxaEGXB5X0nHpIurMSQFoBUzf5tmftvsnR5hPwb+RysHwjN7Esya
W4xUCHerMb1fSrW6o49EqOd9YaRqJa1YPDNMuzHKXU425hYUkznx5twJ3fje
kxRYem2Oa6XhNNdFLhcZnGLDx39LuwXmKuLQJuqkslQWhpqAMLXKk4swyjV6
F++kBrGerpwt0wLky72x4mI+EX/QCv2KZVamdNpOuNrhNGM5o26UI3LEetJL
oktmsDBMHvacZ+ZgPG70e2z80Ae7PHyKW/X/uRGJBuuMoAwzTHiAlRfz0cyW
BIeOsj8ZZ+GZO+lZ9JqVmJIKsrFdycUhJwHbh2FTkni5pI7ozbXBo//Ydgiq
ZpKRacSVMG2NSeiOtUXxRf/gdAwJpIzYcPbxV6O3FF/rTPpWea+FevenAFvq
30sDftWElDGihdQwIXptfNE/HAneJWIPKDajmw+LJSKgmKaeducS0XVWVmGD
Twvy2S7V3koT5zsq40cKHTZczd0lcCC9Z4MjKa5XKsyc0qMHHlqoUGgWP20z
yCkLBHfJ796AMlZisHk36FLNyiO47g/2xr1cxHxCjWLrF5nkLOYr4WNn8Rh9
pVWKIjQwiRznjXocsA16+XbpZd9eD6Ak1Is1aATgitRyEcji4PeB4+E3OJSz
w/4mQ2Cfd+HXKbB1BqaD7/iqYoCSJfozclpm5mn6YuO/VDQ64Z42UvzJPYsW
MpCxK7nzWf0chBcP8w4jhCcM+9botj/ebNn451KwJtvUF6Mw5FaZTI+O532f
1lDp2SmxQp7ACme/cMDMXH/DAjTXjl9jtQ7pGwtMoOeNWNRgaEKMNTeOnXc1
cai5nCBpCNCm1kk6ZCaID/iWgsBynIwVTxIiJp1hlwykskHzvgA/KbUO7pxu
HJjzaLQRttMvMH/8FbkTFJ18onLddU1v91efL4iudUfa1dBh4sljMertFSt+
Q4p4c1fUy+pSPY84BcluD5GjGMTgk7TXFo5wWHDkLpeahv9jZG7wg+4Vhpka
6B532FHmpbY0fD8QP0wC39rG6Hu++zZDyhcBHid174cOfSvXeSchM0CjGffG
ufUvCKqxVH7rWBWKXfqJltRrwWNko1EsbgKrQH9EV542F87eLy710TEDM8/H
ckXjl1oxzNrFje66o/h5ZjXgjcUi8F0g8A+Mxlb6uYI4amdJ1lghTqXAYsaQ
DXMJ0v8P1u/DnllHg5/CxeX9/HdEm46ACxgpZYFLwGCKwimK/Ktmq+3nPZBg
ZaP76oVXFpXXccxzOq9DWQN3EXnOSLwslyUrkajRlRh4Q2kHiDA9E1wBZNcY
gYCisWD0R4KzMUuU0rvxiXIsFJyhUBxaoaHjw1QSqcqLz+kuWjpsOMA0uVjI
wMBaOCr8XYYh4iJf6mMG5o1lB8x1C/RhcZo+Ds1dST0qC7RcMkXkEewc+2/v
3WUTKerTOqj89g6FJ/rFHleuOJ0NaenfBAzIhe/WpgHQeyObB2jCG96gdxJi
2r/jebKtt0WPMANu5ar19mASZbGcHGmOcD7hKuZukBxJtVb635pscNK+rmoJ
twiyFDY81jCamw+GzCkxuwP67U8rZ+dE8GUEtFYTRGiZ5C+FPR7oATOYyEQ2
S62hIM2Cu7dcgqkc5rC8zrrib8ckEG4JjGJgQQ19UMD+2zXMdR6t8Ap9WesF
DH2TOvDudnCHuUDsf9kWVG59AVxlw7XfQErdDnuovrqjkA4qy5bju5gVdvAi
EEmpeINHT9tf2da1Jux+xzgHdJgdbP8QEWLA8dyxbmknPiTEvu+UFOwNiDZ4
ARzeRjYAKcVzvmwpscPA82rsdPPPKnRyhjTqz2SQyjW8Zo2C6nzNnAls+45D
owSgI6ckT6eal9FGgfSG226Sc8kz9keiOcCzbXKzEMTrrUGrpnJlZ7BQhZaT
HmYRHtV+uAZfYRCjVKVmXiiPRjsC9Tp0uTrLGZZQPR32JS2cM7WuZxyHKe0t
PLANtlMsLmDcdVcRU316pk+HGgNfPhVEqgxyJ9M272SNs1e8Ui6VNOXzsjPj
sPCZpNxmTdfa7dnrBaPqnAqdHe7GnjddQ9fXrtbtOyRqR3cqEqpTKBxQHfpE
70RmdWWxN12AZbB9DPBPm5DwLxRL60AtJVqeIqCVBaPBfH0mbULEVLMI0POF
f2EvN+x/ORNXubuyKH4QWuRr5qooPyywrccpGYFPfTKgy/UiG0Vd3PI7STmd
g3rMnzIENy7p/WjFz+I1PwpDFqBxKCFkdntdTw5vhiuvBYLJr8+7tQh7jj5u
bEIshNK2hVnfYCix+oONyefHqXpKs+kb440J/3GXMQMtfo/WSLrW92oWMgwf
nzr/fUZj/LcPWIPGMg4Mob8TSGyqfZVYQYjQMq6RzLNITQeNe4utgRbJhQ5c
5mF2M7+jsCY0alI8DWANfw2A9/j9xtjj1r8LsAItc3GbfrQ9N/VU+ZE3Emsl
zAAVBPAAnlcU6H6IJt0R+t6qVHSf80FBviNghyZ6LsOnBXKdnA6gsTG9EX0A
il9PNESmySnpsOExgkv16y8Fq4jwGg443FWSXr5pLdIMRg2wSz9xBKY+cQXK
jtUKI05s6S0ufzu5W6c5GSWuYxEl4BgNtgBJFORpv5ino0GWY6OGTmPy/aY7
hUSurBNjvFefKENG+5rOtiHmKtJfCkfXoBCjsLRXrWWv3CECsZuxd29n0RV8
NO7/fl4vGlanCObAfG/2XXAGkZU1rF6fzwfBczieb859UXwO09cO15r3Idli
mFTtMEaZvXY17NinsHjUcYBN4tonOE+yzqIqD7pJBfv7NPr7CaaHUKKdA9kS
KvOfI4DHIESDsyeyx6iQPqYc1vltALVDWy+k5YHBrcpRbLNu24DE/Rri0OCY
xU0WgLfanPQs6KU00CajRWy/MUaS9/8hc+nKlttGorIPHIExtMX2mD9MS8Ar
nJVpBh2V1iAG4DmI/Ct1FVWI7fe3LShmEil5Whys4Rf/2UN6E4H7EA9bHzv8
NAXf46BwQGkmPM3wlvjJvMcacQuaIgTePX0zVnEM/PKe5vOaLj3qLZoz8Fdo
HrNwRtqcKL7joQ5g7r9qjmDTivcoKNJKP7s58w1pzoAXcWidQLDCZXEzvQ9k
TZt59Z87PpKPpkONDBHj0V+J3PW3EMS1t/DdCwndu9M2/uv47pz5/t955ipJ
+l8HdDcCc1GtYVbpP5PP4wWazGEPNXqRK2o1PtsoYi7CttIhe7ITtPxLbsHH
SmJdwAwlArN7fEr5muWs2T+cUpoIqMf+nC69K+UyFo1rV+H6YOShXCPD9/cx
gYybZTUxd6S1djvOPO6AbBlejF3QwsMLWagp1IHEVlndKoTE8F8ojno5dSRZ
AGQJKSW/UqpaZ2xaCvQKTQ0luEKKFeYILi37Ehbt1/4xAoAdcdg/AowWdU8s
uRku+kLaIN9Gsm68jVvYdEJ3vLSsZcO0uVza3TajROBWNWEymCl+7bhf3jmp
e4kBUHE23o3nWLAzRdVmNS3MlTeIsa3n8DWA1TkSpXijXtHXNmrmmQriDih6
8fq58C8m5QDg8yic9ovSlUKnjJq5DdXrn9FU+Ar9Vn7y8+YrQ4xHJ8aWRs4Y
/gV6DtTv7sGJ/F84mldfxe7NDdBnMh2VomP/o6dB4GuKzaz1wLEh1qnfJAvd
RpHZoZoR2KhqaiUtM/aevVg5Sqh5TlK9E9kYrmywtnFByo28vwUliHoVVpZ4
go8tEKPbkfkgUkX1ve56LnqcXazas2iA5aLzv4arzap9KJx760u7ayRTEYDp
lLFr/GMeugs5+QOY+ZHCavGxwmtM/eK2sEbDh/EY9mSVo1UOBjiq6QHizAkO
vmlKqKGqXitDxNi1SEG+7rXosye79aDLCqQNSospb/f337iRb6tdwwHmccqy
Ap1WioqRCGyBKsie5j86Sf8Ty8tNHvWZ4mwCKj44BGMrH/5jGC8WCl0GHhxe
qiL5fZuyGJsTdmx1xS5J0np1geLjL9XtogI/dXurPU6/zp5C5KyRRMh3KDvl
HDLCGsZ/bWtSTZPdqM21AGM5d0rrVny8J67caGLm8ubiDpDSvtXZVwExIKdN
Os/Odv+tSA2n6/351cnG15VomfVMrJtE0zKVvjFtu0YIFIP2gpQ0/55nDTO+
yoAZPv9+9m/3rnV/FDfdom/LsPJpiOodHItdOociMd0C6EoIJ7fW3Good/XM
aDx5TmQb1ThwblKWFSGQoqqe7B0sGEloSSLftjckfuevzd99IoOL/U6P4hkv
b/9MENGYiseFOL8Be3csPrXwAxTITjkRXkBGjMsTexEYs/M78lSENPiw4Smm
OsTjJfyC5N0lWUxQhVpLliH9TZGzkyc16kKTtxbx8tAePyE0F1mH7af3Ml0k
aN1fvqkfxNlNX+r8bm4eGPSNLoSrti8xGJCYTbXd0ktTGeIKVA/+ofuhBTVY
qc2xUS+qm+PbiwidoTmnTIeZ0a0ITlRZeZ9i/269CUhHLo4MYSnalDfnntFW
0LBD2wSfWzTQvztpS9HbYUeALvqyIjlZqoWE/XSOXd9Ad7iS9xceppseR62l
BJXqiCZcaUhW6yprM3IA/nRF1xdBOWSrenV3Lr4+dfp8ZfLOMCy+tpJmqwcF
zAapQhe71Szh5Kx9kpTKtzOTPjsZ2ScDRv0gKsUIBaBJ2U48nVZwCiAOjJbq
yXYLmiJblNZ4ySM/Rr1KS7VgntQLu0qa/Y/pmuPKuACq6ecZ3bKdH9Q1NUNf
6PU7luNUgbuTvOasWUQh2AubHGq6KGXow+OwrAszAr2zpMlJ8uqFHY08Poib
7UrzlmUfH0KeJsEIAOwIF2q9tKN+zrjTrM47F2FBFB8iMrx3wLG/EzrHtMq/
SFukYERv9bopmIpynQM265G88hL9z2hI5BF7zcGoLSyztudRYH1VqA68yHUS
8wKeUlf5O30EgE9QnqRGtpCElXEztTUjsj1c0xpmNO17ga+RKhkKypvF6KQO
DEYoMPUbUPNsP9sE9voMqA4wBJgAG3zhE+SI+437dTwzkBUHBJgcnqnYeFGb
XPdz1pYtChqmgXXarR/R5fhSeP+yT0BKT1ZDSRsGXVhlUW4zqIlhvoY0qGSN
9HM/FABDVl+0GjowFT0jv2X0+mv7dji2/Ug/lZQdfzaHlJkyCeyk7nqPKiVY
JLt+ncKVjwcXHUb6HH9O7Lq3KdjwZfxx3VJKUN6VGH6uszekJ7gGfLK1WOZr
JyCarfjilvs43tzGBise7JRF/d5zpRHf4LajPGFW1ZxH3SujLbBfYTJfgvhh
icJgYoDjxdewQFpcLhLtG69Lf64AdJ3VGtvWaLuQ8JgDAB1shEXMJPJ/Invk
3xFuJv3wkOu7FLkKuZLjSBn0iy32y+SOtVynvMZzjW7hXIqEWss0dcbra63N
HvEF3jcVW9ofjqcmLaBug/u9QG1z34bgqprDcLuaTDS5w2y/0HEo3tz3punu
NylSffoTqtclTJU6SuTenz5YgZzYr53UDRfhjlufH+fNYSNJH9TrxIbcoFBT
bRnwnOW+2wy8ZxmlLp4Cl/+wwAPBJihXfzDbP7W+ZBvhoiViy53m8sxHYc3b
x/KXlAJbuhCH83c+tAXKDUlcaGmcf++92NMFOD34mVtWTWMy7y7ocvnr/WCb
+TMZrQcfHpLvvU/m7viHxnVcuOujyftY1RVBjI07hgIXNw9rHJ9Pa83fZoIT
lggWcniefI18r79nU5R+s9v3MKz3v5elA2dqJwrjHX598gq0dcKXvDlXJ4EF
rPuCSJUYYl49r8TIf21vAjhCsw+kjq69w1fdJt2uY6KlZ+B8zQbX5JkwQeLI
rzcl8GvVlMvymLMFniCAZNBBI8d03mG7GGYMzYGoV+D9ecwy2ZGY2NoJpOcK
tb59kzIktaK7nxOFM2+A3BG66VyBCizj6za5GPmkr/9pjJEe25cUrBt6IPMA
TE9CeenjQ7/HHz0yZ6zvj2HKWk9HjG5TV8p0un7vqUcH/ACpIQakoMoCpZGR
q7k3a7tjwnxkCJa4bMiKYKPbY8QXD87ioumq68qEgv/9JQWgfQtykklIxeRO
HlD2c7AgXCFf1wOyz2SKcytH/L0oEHhCxtWZDndRxrFWhyCds/3uB2cK2CgG
oO223cohW31WWOuubprTpJu42y92xvYMm0+hwxR+UzvvQbNgjSqc0hLCMTZI
yyFa3fPp1KTFXiMrvANHgROTO8LGdBwQgY6kuLENFGoDyWQCCwtGmm9qq6lo
iHhemtlsHC8ug4fuHrTbuDdorHw3l1uIGH4NxA5brati2/f363WpCPw/q6+P
cp1vZ4nEIsNk/HHUYEGyuOW0zXSKBTIVe0dyyEXZ8U1AzGSYKzoI11f+4DRa
UJ127biazrAfuToQAKUi2Lf7kfrIyuKds8ob8gV8wMphy5igJNl9g0QRURpI
bo2WWII14Sq9bzSBfP1z4ukVlEW1f+8Pa/DAkw6T1ZImNL9FlCCq/wUcoD2a
GWdL3xoAsaJ/oLrWfnIE4C6jFQvgItaZ8uIPCI4cT+Pgsp1lxm1bHCTw3ue6
dCHVqh6Cozu1BuqilnolRqJ5g9pGCf5URbi7Sv/Bmtr14zh2tjw0tAWQ/ys6
1gsi8ebG4hOP9RdmlrgGebmJJpebt9NmSwzJgsXmgT0Xu1lcE736m5sXYHvg
BqO4SSnUaF93tNIIZhQGdn2caI7EkegBcylD613o/MxD3nHxsBQS/11TJyJ2
q0OHke9DfXkF3fpeEw285JFzN9FNjou/v2GkqVU3Id2l3ntT2/OMkz0mU5Vh
4P+QM60D7PAeOtze0rBcIYBka61qnHprQ5mHWyHFSGTMEC8n21NmQ7cIGtkF
4AOwW8FZagSdYJUXKbetjAg1LfLslvXDRjTW6fdu4Cgavi6ZdKlHuvT5dLs5
l26mkRZ2eJ+UE9cWOa/9e9SrCoYVr5D4/R/jjX2J9Bnz/PS7DeOE2SAxns8w
Bv+fLjLQ0GvZ7OK7bvYHkYRvE/urznmTa/SJX7iEci6mv7GDT30tTsQR8Hf2
ORDGoRrw+0f4Fr/+phu2jiwWUVrpjgdf+4qovvverZr0tbSi8J23Msys0OWE
EY/crwHQQCPUU9fGbPTTnDNF04HqZnLdzE8aNYpTyi1VucqLiUgtS96SPSzK
1CeJYhLBLaHhGGUsI2dUjbS+R7bYAS/WfJJmHpUewmBv+EcwgcnJBb3wbXya
SBQ6b0urtrW8jfVVg6i2OaI5XfMMedRYFeH4bksmsaNsm6ZNjsNP+HuFowYw
DJ1ryMTtVSdpMtGKgWRza63AdlKG/uACE3r5lJv75rF9+qvq9P2UiNqtcCYs
CskYbR0rY3oqyN7sflVkOxMGgsOJQe6/4bInEcZVvrwAGpdt3gdQWkCd7eb3
QOkj3mYa7l9I2vG9RPyeDao7lPs1rkD5+XM1F04UeY5p7v5pTuRXhBUHjM9w
6Ld34lZmKU7KYJoYFFiLC9Y94SmtrTBfk7w51EvN0gqzwY97FavpjFSshJPS
IeHZFd7NH3XZc9aP6ewZK+hzesZJaZaRYL2ZMlHfKf8c6trg/pHWUWuzmDkm
+/zVrnmX/0PwA+p4eYT1mSLFKecBrJryOPgIeUd/NqdEHDLOvQBQXkAROO57
OKVoegcK6iiEJJEsSBNVyUG2477RilIPj6Qls8COSPXd+D4ZdlKcmvjzOf5j
VLLouQNJkyuFK3ioeEnHwCXBuY9MIHqA7tQBqsqUPy+5sTKgUDOyPml/5h3u
Jhb8Yf28776IHvYHKKKtZc/y43b03mqmwBTJbVLqSfugtSNjv1bET/sN8zMq
8JSiiX+ZNa3oQwoPaNvVic5bwQOCVIuMmUXOVlsrgsVLqduLx53ZUdZknnDm
cS2nzkfPMIs5zrQLPGngpRM1Y+/aDvHGmv2k1nxeOHiKEw4jqcdHgRchOhmW
K4bgVEtXwTECqF7rVbTp0wuXXUh5FEOq8ycv1itub64tFF3m9poELE3I7goF
c2c2eRzFdf4xwoNhumVx2YS2KVjC2SyCC5FQ3Pckbnv3mqoMPztl9V8CWHSI
wCRVKjHHJXxiwwkaRFOHWpNw0Q2GMRsJwgV1xb29qnQTI2Kb4UwwN6fA4810
ysZQX5BNo6zCPUYJMSLLq23zCEOfghrLVC5sCPdMFCvejfA6GrdxWzr9sB2z
0SU/bqgL7Pxzzkqlf+xkSWRRH7DOFs64J1pN4u3q4C44lo+/Z8Dq4jDvOfzh
zqhKH1B1mrL/iPgJFzT1BkExruLCntDeuJ2EAffksVIOEWJK7d13EtFLKfka
LD917N8TRgwDWff9jLSh1qS2eZzB1hzoGWZAjkMxa7zJ+irhfkEGZP+Z3ZG1
m4PQM5ksHz6sv5Xq5ba4OROGUmThHB0Pp3kY2ejMZdobMHliIV+pagA2O1nR
z/HVNjt3B3myOZMCk/O3Kiokls0cC683mL6c2i0pznAzUgIBEuF85ruWWlXv
SeYN5/DqWXS8jngJTHMITCwWebI5uCBT7gh+FFBHzxSye6LIP+tCHiMcczfV
Fhbv3VJ57mas6j50YdxoQB9uI/3TomaA1uA0V1YziXCWzjtwHS7uunYSnU5Z
wfnsm9pSU+yvlqecaq/XNLkD6ihKDNxGiPnEeEJKtGcFv9c/tfIpWPjXDJhv
zyETzrysv6dh+G9orAa2cnlW4G1gMVb8vhk8Hw4zqsyppcMlvCZZp52yqcLQ
OhGcZ3o7Ml7iG4IZVIYCZoDjbNI/hiTpr1313e+QCgMATfgv9oiR1Hi1NPt9
4g2Q7FULP5guAEzN5K1ra65NrnQXyORIf6CxrPRSKoN++dGawx7PM46AyCUI
QQLBQv5kgnEXIl7Xktde9JIjuxwbIpZ2I2y8Oj86rIowic5tAcvVzftAGiUh
79SQ9pojbU2LIJAjyMg+xrTOycCKCsekywFx+AOFI4HM3x8n5xVE3cOOR9r2
4czW5Qjx5ctu0aA1hkWA6CmEmtIS/9896IyeT5abggnfPUNe4s9QfrOPFaMl
RGxq+xG7HExBvSg+sbR5bi+UKchA+bal8oibl37VzUv8LSZwjpMjJD4BwJvr
e8Q/m4Xf/7AfQUhHdhovY/Iy7fBlFdFyIy3nFvV6vYkbZDvpsSZKQ3i6aH7k
hvtj9LQz5lxHTQ6mtxBasgBAA0WLd/GdndcuS6NliEjXKHM7F9y/Ua5mqVi1
eSayF4F1DaEHujPo4YC0WbNRLboxJBKcS0JBk0VANt+AtzLds1TxoPe0qkjS
pMQDc9TP8DxzoR7hMADJt47to2wLeunBS6zEWSrhZ1Z/nBRcpRmfTY8RA8Bn
UyZTLcvs4vdhp3Se7VvNwSvGG5CRMNFsvNswuHylbwFsiutr7A0zG9qePsjn
4F2rzpgQofAmRT+eavdIvXhjzLzobCa7iAmnsAS30hwIilu0qSp6NI73TL3B
zbAg2QJ633PbTe62vwcfx6aQNwhwhzWzTZx8wVeh+VAQAGiZ3V7s6U8zScFv
5n4Lc+qeczlmH6sx9pGUDJMB+oiZec1JzqfWi7iw/vKoaCKofyC4XsfAVzxg
t7d+AD2mXOvbeToGzq1r2EEeoakmxfpxSQ1HzHEx9cKue0jCY72oECx8CYhL
6IMEhk4RXmQ9+JhY86od51bOTG7yQmsT6M/gWQJTAwGi9xbUcmmhznel8ulo
19PSVpIqSKMPqxlRo5c9EJG/IJpeG2tTB8bMl1og+4W2nfi/unm8dAVk2x3f
qmAL0UIcJZDzzk7ma1xO93DKMZNj3uJp721ErOvUAsDPd5mMUdsiDBuyYrtH
FAdv3chysJRXrahCkVll7U+/hLDKAUfzcJ/jvRtJXDoA/7CgRa0iw3esBswB
scd4NtKKPeZuwkfVuxLbk3J6MiqVoPPvSUYHFpY8ju6RiqkSUhj6CmS7+aDV
LqbEHbBw0FOWHwlf0Ds6eYb2vSHE6Cvpc0gNLPY/MekUH3LjntY2rAOGQffJ
2BA2o93hV54iQsw0fKovDIahoVJ21zgvAfgF0uF1+bxBbwiB63tvH3gP9/gs
pU0flytbeaS0F2VM4OXV14DF+wxk5Ju4k6SQDgxDvZWvIVxJ7CHWR8trwtbg
ak5RHv8qOnJ1+jV4bNWLCUgL+1jkVkDV9qWTt9hzaewqv6VGwN0CPnwy7He9
eqbq9+HAPwLN6Vl4Y6pi3vONuiofoNX+WEIQkldB39mplV1wKRB/iSHo+vr6
imjT0qCGSgvK3Bhi2fSxSp1Rv4V5FoDXNHD1ltJiHf5sfmdxCulmhPeV2zRZ
Ruqar+F/4B61a6XSw3EiuLHMb1PaINVoChiQBEuL0s7ov2YBlmSy9JsMxP8+
C/Dn9hk4JTdoAPTagGc4J7pZwJwQOpXuPIZqSpHYUEel9GlTZVxK4dn/DmSt
c81q+BdFUwv7esZ8reFPcHMKvLcCp7Iv/zOTAyCbCjTOD47N31H8r57DOm6F
xkmqN0GEDSH1E2/nNB24UTn6ci1gnfC5M6YggmD1T5j1156clBcTQXJK0U15
tTd062bomfTHmBxfmHzQpwyyli+IfeYfluwzV7XLOLs6l12yv0BUbW9Q3Uxy
7FKSb6Ot5+/tdqHhn0LA1UaIre9uYOgAFipzFQjsaZ7Ey40LIcOaOKAWvZhG
1ad4/+FC3VK7DRjlrFE09yP+orEZ9zYwo1E0kotZim+j6V0brPlwot+Cse2G
IjnaZLSSI6blFvySzusE/hR75v0Zl/MkR6FB4CGu5y8qwTM07jvrRKC5wMmN
y0BTEZ/YX2aEbpTCdVahEF2BlQ2M5btJ0HuYdKRKh6l6AAESb1zWbzwtB1MO
nnpC/MUl1lFoU2hQ9l3xiUG+P63ckIHfg81kiW5FoWQOQRwAJQ4gME3sqgm7
uyWgdVBACw3rLmVzIh8PZxB0M2gHkKfmnNTYu0Wkp3RLFJnYyCOGHYYCYtZx
K60/gvrkcRdt0VLjx3P0CFrHgIojUjsCUuwJ52pmIXsedwTczkeU9PQaWKCn
C9QUlQIGAdG2HDYK0HY05WzRfiIeDrjImg928D9aNRU2I1oiFT2HDf7y5YQ+
8BGYnKwnX1eisyf//TIz4uO1qgX0tCote20fSB2bVgXGFWBhV22uAstuRDXu
9QHTfGJ/J2iCA18H2zwcV20p7/mwicJlCn4tZWrZ19/eyCXQQhwwoFakElAy
ObNgWtSqxXcZ+bPwRl6unm8Ti3sZ0WeLlqFAZo5lCqzzm4arOf1eexNk3A8j
I3WQaHzuNrrgAxGxNN0+Y2QYa7YaKJ59FaQMr1+HyxaPaH9F7g1bGruxQVCG
dgHfXPFGI1AWsIz5qv9Pu8y/KtFzkSkInGISFkpRGTQD4dX4aWK8X8xvQn58
asuc8KeDB3TMj41oKJ3wEaWq0ffyCOy0TxdO4D0aKils5BTFZ9qzoyDmjEOO
YWgQlfulCcgxj+nkS5kzvwMrrwPevbSE2NnmPLPShBpDZya9opyo7TszPyOu
706q9peXDqz6sREZhBR1MoEzaBp9FCSxD9HVRt7ndL6ViFTV/z2fgqRlDNly
eezu+Dh7DISxp509+yEc9b0mVscrKjrww7FYaFaT0CVCnKekjzdbkikqFEiv
81irvLQb2CdhjhYYomLFI5WthUnwHpuU/P00qIlncXKS6xlUDyOlyvFWmaXx
+7TUOkvlKp/EvFA0vlIYythj3NYKhaTyK/q+zK0GjHa5F0ObtP1q3ror+mlg
Bb0ZV2Oz9za00aR//yLnCIHGsDigf3xGWjhBLju1t+ZR1KFnAWVpj6W5Nn/8
E6lSug/ScgR2KokuUBYqUaW+IKiZ/C3N02UShujg5L5qhhU82t6obZYncNg8
ZJOYYKIYfxarI84VnOSophkY63hfaixy/jesYJEyY7zcQ6mkzYSY9yR1ob9L
ZJaNIKjRy7JfBW8sMXAkHy0YuTiu/MQdFFa3OSCTOxs4to5GG851x0SkB3fJ
xEUEfOqKX/57JH2obOz3WAxjDD0k31GxyiOVGAvLBA2aAmZUgAOyY45EXvQu
EAbaKWj9SmvkfqSpv+dsRpWWzX/4G0hKeCWykNtaV+HMwKRuvqO8e34JDanK
9FXLUipDZw/ayYle2vNKRkcpU2Twc3rWNRQTg9Nv2w1L9+ENAXm2q7dZj6Mn
vL3UIOGU62QRV5EIO1V8uotfoxS0lX9dAeAe5TJ4U8ed3ssI8j0IF5+ikEG7
kb76+dH1vZKuX3GMEP6Xgz1zCKa19f5zCp0PkKpjvzzxUs/lpCpKTHEsag8z
aMfn766bnVEBtfwGCVtyGD8HH8UB4AsSI9u2oPjKoqNFi6gB5Nc+mqNEjlsl
ckKnngffdkYEDQmhJR0cpx0/cWRaJd44ucI16jbiHjTFeQW72zPKsAPRNm25
YVDu02nIY3DiDeH2rl5vrAsX+6wXD4UdvcZ6qOkCNZAV2v+5uZHT1+HSN1vo
nl5oVOt7JDZppoHx6XsST3B57ZWuN9g8wdf7ODayhJNFj+mzrYlJMyN78/HT
iUssbjx3BtjAIpED7h/wgqxfkWTvJgmN80qIvk3bvmt8UCVE7MDB+UglPpgZ
QB2bqbPstG0zmAvLMm/O/yhyofyGGpEF2Pb+nOQbc/C0f1udKYeXO4SXase1
TbG0eYsW7Ybo3evmurZ6W2CVdfNVVsVDCt8Qf54Xb+JgD7GlRv/DlJ7lft6Z
WyDZez89aX+ZOk0MbLVqGMO69xIGjTnbRYys+Cb8NyNU3eoXlQ1mQG0tRQbY
LM52KmJD3dngN8TGEkAqJq+HPhDNuGUWs6MKLqMLLnSjnA6SVhG5k5XBRJgm
wdWHwSDt1Adw4lWBkSZlyTSWN50lBCb0bhkW07WYrADhFjE9yXQtzQk4lYG7
NNEZitTuy5LZDUckiCEDowjNFxbmEWdfNczku6Uz0CTrXyUBAE4x0lzvg6UK
J+5RSOpfWmdsv/RCzHhuk0GfYIdzGFGDFrUoCj58Cr2dtG8oYjfac48ft8EG
WH/JJZi4PXvfvGFdz2cDZmb0CS1eJS0/+7zGm4WkTaEAnLVo2gbd5IWcKVtM
mGCyl9uvZQuwHBTSia54ihGkP071WMGOpgsak70VO4iKy0B9uufRJywZCh5y
82gmNs+xF2az+GJDD9pGq0Qj4Dm4WTfVvcJofFDW6G+vddeYoO4hrGMj0iqX
6su8cQN2/BmtMAVrD5nriIl7ESBNO1XY0Vq1y1nJXXKfmMOEpJqULSwwRS2w
UemRHtjcsvcLpzj0PVrPlqtFHD/pdmK+nsPsIqbzVtI7cDuEJRr6zhSZgJMC
NsLlsSrgptynzOBtQX0QXXcK5RjVe7Mw+Br8GVvLMNq/eQKqhsu9EbaEcuwp
jl+SynTzAbdZnJlHXntp4c+ZM77v+CavXwJ6kRMlJ6qfBSTdwMfESuXCbtcV
KK89yzIP13+1MZZY7l+y/YVvqNX52wJPZWwCQmj0xjVumAEHdqModGtqhTBL
q3GX0kyb8tVqMdQmB3iuWTlhvdLGfHRDzxDD9siL/xNarIgicmpKEh5pS+XP
Vn6YInvJEygHTDxibTQHeo0APlolHJ+SGvqtW1KniQfn1Y+vTGliT9s+Dt/Z
98u7xgK/YUx6vdrEds3+9ZZ7JipgnhY76mrppTaXMJDaH4qtI7uDjiWS8e29
Izfn9BzIRxFaq4AbRBhgc7ey7pyAfys2K9VuHzVtkTj/Xnr7VeepmgsztseP
pi+CUQr+7gdY6l/uUssARbBKqi0XtGXWwZEaExUUe3prj+EFfRd4vfNmVOBu
9RftumOqzObiDuB/XC7QlbUA21mAaW/LIrj4kx5Iez68MB5RZJh3UpReuaGt
hN/gW0QCCXuqbMmPnD/eYovKdIZR+bSHGpqv3I8iuqlo8PKxYPaJ/N1T9GCr
AIi8kUp2dXjTSmlG+vVTiwLaSeArDNbOpVEXisVwvSNR8Sx0wdHL3dbDOFT8
+/CqJK1lJKS9h1+CLdWK2bY5pgDGkzMqMAfyK/UZ61POEihjI5ixuDcjju7i
+AmhyOk8RnnNUzGU0BF/zu89xmViuiJt9aFzDfHOotxD4X8WuegLjhS8m91T
q8XR+/67YgiIK72oCxPdgccnNNh6CFsejAIyFbrGbaieK8xpoE3HPuUeqTi/
+ND8EKhtllo8nAWJO17M+Tsff7jsOXRhVlrh6F/PB8fxwNiNsvDAphGoO1hL
FEueIKqMs7aWr7YGECtF20Uwbg6abC3T8R6E7XeJrxp+rtBK56o+PZV6jtdq
EGCsR6w61onFhMq0x4TBmMgblE6954dMYmn3rd3sVLXokfl/lol20x7zeYXt
CsS9d1/nkoq9k/7i4Q5qlnmC010rbZwgFSS5X6U5+EBytmNzXn61kq7+ra9w
aMZvIOnL7SvVdfUWvCX2fmU+Io8SerwIHrf61PJNlaGrv50v9IS57msOVSKi
G973LfF6GI7ITM9Cun6QDAxxZGJXufM6CDGaijifbLk3ntw3n4obU35ayiL8
ZFZKJ5U5CutgESXxOZ4pvrmQ08VlCpJBFIZnEUW/4CtJHY365mr3YZOmM8Fp
6zhUORnY2G7aIfFUxBL/RSCXqRqkKcSFtEQEGV54zAWCzTv7MhC6ekqD3ttK
l1dAQULC6IfrWaLu4scUCmAIyzjPVABvm/XVx1PfSmtziI8Lji0Kdpq2eK9y
Rndqbl25abgKGmkQzVyEzd4yylpL6WIDUad/DdvMteDYvoQOUWg8fXEEagvj
sXbfimRhUH2qioqa4OHwQx+AAz2Y0Q/6ZHxRn4R/QH37Hm4N+DT0pR9TesF+
vL31c981wPVkcUc1WeIPsE8A238Fpvm+qmpSpMDF2QH1oiUuv+div9+qoIBG
YB/4dS2I8l/La33lkVdh/8LWawt/Hh68Tm7oE0LCzwDpG27gWEYco+mcZ2tl
qG0BOhY9wUycuOJhGqjhAu8LIlQ+W1zkmVInAicqdHx/OVhpUGZi1hRPzfsh
mWTQpEpVslzu85szJILKgJ1Z60bs/4njCobS2ISJmPJ5kJ1sXHFwMasueVoZ
plVFkr9tF/L7lxemcHBrQjRifWCllvFOyq9wKX2TGy8+KpQBLeqkZsgkIQU8
P28FODUY9INobf2VU6UwenHWpU0wVQ17fT5Cq9KrdbmqZkZAurWfBqTClibr
qLq11QvCgyKH6Qjj2t2sIF+hLmjPvY3lRUKXsYPkmpTDLWQO0yHICWhD3rRf
vSHQEL6lR0exwqtVcsMvVVEgZQF+mvrlxht9q5hyB0m0ZMG6oLTBbafRExl3
iKhfmmaA3rruJl8/yy2hI4WYFljJF/1QpulI5Q5Q5MSVpbFAZC4MX0QOZMr1
d+0STwVLRtbswPreVj2ZllpyLUpqknXH6pHL74L7WbiqSFkCPjhn3i7jtW7F
vGWh0YegyFW9vLw3tJfefyUMDBnwVjgB4uo/Nxx+8R4CmnPp5JXKtPF3XSCO
tWR0b42SVJMRMaScnYa8j+UMBUrG87xKML0Nt6NA+jSMBzvwMlzu4vAztYml
+lu1c5AJs8hWMMLSAPjOQF3FSvbB3Xb7d/F8/XDPhCimTdoh0YXxRasrKZGH
GLwTdo5kFHhAMZRaOKPoeBAGPtRCWm5NXWUTwTAXIFdmRRDuLxzJ2Llq/ghW
joqcQUQpsVojsmd3Vl/qBZpvrR9k1P56k4WIxnenNTg6tu1zwsd3/7i42/ZX
5VV9/CSAl+P+KbAMehkGDIVYWi1XIGpCXCXssHi3wI/YpbGPTtXt3G9vG9Qy
CbFWTQihLs46+JrV+e2ZtEVLprMLQmERcJXPjoaCP1M//UBdt+jZ65VvgzZp
ZNG76CrVW603w3CYw9cYwHUyEW2kEW3ty46OoSamLX/0SVHrL4btYvVlN2zV
3aQXUHdIkmv8hbRo9alC1V7jNtSgZE3snachp3EDmerYJ9VkgKQxui+YZ5Fs
x8DUbZ4ZG87L4c40PsUCQNXfZVSstRzbBQ+0hXanY8hDday4KLpcteWrQZNb
Kz3zOXeTfzCQGWbn0i7cyL+wWdsxXqDF2po1qhb8XMYUzutBFDFk5PC68vKs
edsDYsum9QMz2MseHJKIz0AAn5+7Smsi4REcKfwy75eAz0QZ3+wUqx/ae8Gt
pFQZNc4KOzepVcrnkcwGFNnwYYXtfwEmJHTdeBYgIgTTjWDfMScgYIhN1vri
F1Dfn98kERMETXLmwASULVDdrjWvjt8FgRbZFGa67JziPhCiVMld2LoySEdU
uibCtAdeHTAw1aYLnbL7JK0ENhxRNwE9gvnYHK9mvGlyf3sfLIjCUq1lSn7l
S67riaHp8u6kuUDvo78/BR5PRT6jZyMvOTBwZkjjOc6bo/CtqQ14VZ8qpekz
JsJDYnRoXkaR5mpy70J9fJ+VjhPXTXB/BaoyHAHuCV5bGqubSuj0qs0Liyzx
nYVNBkWnUKR/bht/fgq9L9Wbguzdq04kmmqDB1v19QBEU37xTCcf+fY4qvmV
PpRN5665KYtValtsrbvOD/MbwvD7/wY4khXVi4TQBSL7Qz9Nurx7abM/BE70
s1mrw2Od0ZhD78By3mUgapiT+eQ1YASSVns5jM+FLcLXYYTc3xKFRLNcmJLO
FJtRVGtOTxcuk3yY15vHCfNAbRsh4GizXJvO3wAaTMJD7kFoNEI+rJ/vs5ji
JtaUMa/1gQvMk7TD5YJtkvQwSLGIgS9VwhwV7ItR5PEp/DIYnpVeQ02KMzXv
hOH3R9bT8TSb/GXR6ivQKCQ5VD8yi0GkYsdaMGRBPLCC10wwiwWp+veD7iqx
M2Io6EXCEUUP0WVcdrz9vWgsDiTpADqW9Y1XBx8EpwbhDlYaVIuA37Ig4SCh
gFHLvyKaE3hor2rgfhapf712WTSZOAkSIGQv8Q2NvcP7YT3Gy71XZbHUUIJf
ifA+4V3jrQRQChfhSqJkcpJTRk7EQ84Y1uWFZluK0VQwrQ9EbxoCnrGMS3Bm
NHYdVwSHOkmT4ZLIT3yLQu+JyuaV6RUl8ZvLvER5hc4nFKjGPOslYbxa7JIR
90m8OeuxQVVHcK9U5bsv/x9xoDOqIKFjRrCl42bSx3i/PAg3objWAeiBzE/b
qgYK4zU0hNvVpB/2EGBwnrt0AhwJuu5FUT2ooRvC2+rb9LnuQNCHIKnE5Ow5
YhJjXU7/h4XcKJPThJbCrXJlwuandcmdE84+AapNU7FpgtsBpF1AwoTAMDPU
vbfKIJdsY5piSR1wA9iQGGup0AwkwJw6VzlvMLO1dqzSvDipUwEzVW6C8F7o
oCXTVsXFS+u1mWeWpzCOiemwhpNoCrsbrrKdGH0EkqREYjtlWTj+iy7F/Plj
ehVTy4ZgoPcqg6OOEES0weEsED3MtkZpmeJv2wZh840r8IAXL5c5HDSh7gnM
XvlHpFCg0VytScSC+c52g2ANQiyK7txnU/4+rS8xmBlE1PuAZDiy9D0Kk/+u
7XSD8HYROCkvSyA0UCQbfI7Phbj3o0djTITQP3nKnMJIL1BPSB4n8mmcKwPz
WMtXMyiUrtInzN0229NRTgfNnMQiSzy8jamZFbDuQuMAjEfNR7oZriF8kXr6
Sisv6qjOj67JBzry/S9hwVdBuQ/1xkvPG0Y/sqc01Llqky5LH40sCwUZU7V2
BlGq+6DJHV/GH/xTiDSHHJpjK/2a/xOdHNnenfSzGRetN0PP3qLAe+oewdxp
6IYsjif+Mlm/EJuQfODNTMigK6KQC1BoqUdldrFPHaa+e8R2SzrgSHM6vaqM
rCs8gX/ddVzQ4/zHAIAAYo6l54PYgYZoGOZkvtKiIEJ+1iq07XjtzlRqAgG3
vUvc8EWWOA0wDskcqs4hoeeSRxMJ7/Gv5sdrvJSCGS4HREJoUlrEh7IlnY3W
9ZegIra7r6vV7qyazuKr5e8bIRULvEEjusrTdE5/OLKoZAvMh6SKKAcbq1SG
Do60kNMm/wRBQY/5qkEYJxSKcrClwbNViuuBdXRIP2phYW9oPeCMeF+x4uFU
l4YE++mos+qbWxjQJciMH3weqnvbZcxxRJsacn1nmSFzfb0x0JxHKG1v1ZIb
8GXCmuB4kzmYymdy+QI6Z9KLDemK479eKsIQNFqb4AuOSlffluxbMvtR0VCt
O8Y89pI1C5Pmmw4OFcrNowO5dBkzM6//1IUpExYC/0Sp8J4n18dyN88mt4AW
Y9oqchTjDHV0IsA6iQWxGjFhHm7qh/9YFIeyxDvPi5zPkgubSzgE7WhFmjzT
iUPw1lzy3sdQOtofw+8MKkbX3BWjOGBeVY1jFpGsQ8gwbL7pT61Ozre+gUsV
BBLDxlH4pGKRUCqea4Pd57qCYssfgIBaRH/B04gn9XpJYJlrvndc0uxuToit
4IhGIdZIJHlThnKGKTPEf/0Wd9DvgXplqt7gkY+LLFXK1CPNcWKI8jCyjkoj
7xHWabhLwG7bS7V52XnHLlTBDX+zz+9lq2ivzc7clzng7nJsSirx4sOyX82a
hjVk21Xfd/NFq1NQxxwxK/XWoH+hOmyX7uK1P3l2akmPYyQ0cSvHx7viJ7XI
9o33LcznAummKw5kH4tNKoRPvzst8XhRUnPPlzquJMD6fAQbcwK20PenkEuo
vzJBJoW9339+s2+U2TuAvMTFnc6ipFRry/BbGCdhnFo5P4HyNUQp2S8pJqa0
yMEolRHuT0q2cVE6TPp2q4rwvy00dA5xeiJG9JAfnzhZog+fBH0hTmcHsjnj
rzqVQeCAyPMg4JXFTv5MA/+O6gX5DA3qlQ6s2DxuWBBqc2cLe5Wg6v2IMF+a
Qf6vGSqj8iseGBGygGE3QAlfrbZd7+jo8aGAYGa+t8hjcc+YbHLu2Lvtp/tM
gThXt9p4QQ2Pz8qQ8xhTQZdVa5hjXC4Euxo1AH4ZZb+GRXBNSu4JKTCJZRhI
lCW13IZuFLz5bY+lR6qhukDwuQUHmiqmKPWQmbRjQu9w5yy0avl/X4wCJinv
D5YrPIXZ1mKqBW1m4BTc3hHlKyYiluUB7IOdguexk0vy/PTae9EQq7k+E25j
L4DiE5hEU7sUNyMwJO91nQrsE+kEWKXHyT36VsLf0R/Jj0t62nni89rRTH5Y
9exTOAD+2WbkUoMPoMBjfnPN9YGyBFzFd+BD1nCiHfIiyZ/3uU0PkT/CMY69
gzUB5uCfqv6TO5sv2Hven/phF5aMuiQWbfAgagJRkTYNn2bMwo0d2rCz9F3t
SeTSYOQhQimoJ8q7LS1mbIAFedIw1EpNhgJVI1v4EKl6hJI9x9NKb3greZNF
enBbDh1sYrBaYNwh5qLhk7FjS9adFmYu7XQAceC6J46fuhikA4ZDb3WBe7Y6
gUknUfTj4rhwLiFzcycEdKhpc5AQUrk22PC94Wr3LTElHkoIvdSIh15eU2mR
Aeov9sjpWrECk29v9WTuhUzkkX7IoKrk4nnUG+CokZcAHa05JXRc19FE8RVs
bp9oAoRQqOksY7lO/oNhoSJpLRKEEEVJBo94ATCz9YXaHgZNLqsk8YSwrV1X
HMMWCuFpvD4xKXSNUKj3GorpuiX5oNMbZSwEAywaPqcI4gEuX3i55Va+2yVB
nWAuWCmHmN46oh9s5HHuAA74LOsj2WpxkkeYe6Tbnb2ZVGyKcDqq6NpX9AMf
X+mkVt4hxIQdrGiIVvzeIeer8rLMehBwXYbAqMWXJizfUK23swRwpIIgQ4Wa
REm7JFpeRo4ql0A6oTYbjSvFOOpvV66RZkdppq0eLMw+JBXwFlI6tkB9vyMm
u4H+A5DfX+5QXnLhkYI818ukOUXyOWHq7Ejg+iUeOpJI33ZpzblbYULKn9Eu
c5SISkG7HmVrn8VtfGDfUaw5dzfdkDZtWzX6bucIopj/4j7nSR1iJM44zhOt
XxExyXHscwEVibU0QKEugYUo8NViJ/fwLd1v0XQzuLx2mITbxG/NIvrGBiVS
ev2TwfOE7g0bn6nQuiA7WER5kz2AMljfU0aqvlgdPzyg0cBwahUN9Ps+ssmh
TcFLk4xoePtOH4wjhESMppctfE9gBkPVsQ/nRuuCp2/QAV9J4O23Hel+yBS5
BV5Vflz736u3ph1x5k0M3XJqbwH4ZKObXg82gdDpR+DnJmvvKZssDrmDZy3L
S7hd3U+x+He4M6TTzotxSDSd4sYDVxnT6MDEbQJ48kOU+wt9duATe4Hpm7pX
KsZYqThL1nDlcvNNci6RO8gMiiz4/fUtoKBEr5LNQ4HaQg65KiBY1CfA7IRO
+HuYtDp4BJbfTxreGRErOl9YqZTm/IOVFlKCASPA7FAb2v6Ohsg0wWuLx3t8
7BCiaqFh/vcybRI2d27zITvHYYKO7qxLIA1FXalzRw/IILhiD8b+29nEBf9l
fRGZvEnm5jyED63CrLraQCLDoK+h4hKQN+RniqQQz/hde/6DIG5O71Pzskfb
FwwHAhj9BhxGUDpr+yoh8QQw7Y/pmYPtd7HOAkXv6e5uTmZv1znDDIWXbb6D
ijiEpKZ/F9omYQcb5mejVmHpkBXRCsf6aVtvSlJXJuwQD93daPPeI3hlB/E2
9HLllShfMHJU7Pbdn7AGczmm2lsrguM8aewZ2P8/qmIMV4+SrddqieLgJG2f
/zU7TX7R2aH++Y1KmZ5MU++UgcS2r+vSE9F99uUY0aju5IHd71aTlsccSYuj
TPppdLPIufvwpDjFon8SlEShu2u6DOAjxucUy9EN2/6l0EbX3ISkbV7rafOA
KF53Y9oM7bgUOUNqRfWbKRwnZ/nj05jKDzBwOJ9ET4Ajif0u13ixDdZeP/nt
5WH+88h9hPY42FomAexhLply+4A7x/i5o+JK/eWKs6MjXO8ndxMsEQtiev77
69DzJb4TD7ABX25GC/mXAl9CBNoEz33sFNn1jJ7WoFYnVcjH5hXO5BQRbMZT
Q3/b8aqJW1HoKz6X2MLTezOSJ50PwGJdHtzsmlKE50Sm0XtfhsgB4tU8LuHj
c055F9jL09SIjuW3Bx4qrm2GuS367adEk1Sz5RTjQDdF/wz2dGTyDXEzzBJH
Sb+OirpKJxDBGeo+LEAQuUJ6UW8zVT6FgQhMY+HoEFtYKeyJD4vpyyLOquL7
Zx7NnJvWDFpTytGpyvkterYdZdMAIzabDivQF8r3Jdt/ZGvNnMGYjbcLFjXW
YXLdwSC8P85s64geVS5TcptFCD559sHynbdelK1Naig2sIGz1Jizwx2rb/Nq
jXNSeXs5QfXr7w06C9FmWdR+krqP0GZDdduyUBlqpfkYDGzCq7rn3/QuEznA
ETDI+zmi5I8WVFgQsYKu9oHvHuvpYRGTBGGrMvHt3xBwmpGUU4zFyeC5WH0v
PzbYpS9FR9Eo04GNTUpkFjMj9QMfqusyN/8RWzNXb4V+EZ9zKGWSJxiv7mU/
4hlq97Lhn8VhHcPWscjtyuPradkftM4PRD5NRL0stqoIgm0y2glYa0kdEd+/
WofNq6/MkSPwQoTPIOEi/TZhpm98JjwEdKNd3ChmEGCh3qb5Wak8l0RDXl68
8YxvNc+sICUP8mAwW6aDeGc6oIghMLuKGOjiVYQ9YZwIs4AwiD481nvWd15x
NtXZWD651O0KBrTr0cPiGu78R9dIvIZovYgZ0T1zGMY/YfWEoxiK6hDEB+KP
Y2txHOpMZnPfwoDoO0iq0jDEbzWY4lt867UddIsnRbA4KcWl6yhV8MTLxyQ7
QOEG4dzR/9QWJAS9zHZ5a4L5jMl8AJMi1/h3fYBXotpVPMRGmeSdcrxeXwxc
nPtVpMs/eWIgGugKspcZAf50E8TW0bhROFmns88/496hsS0P4x2BWVQDbBi5
Gm3BS8G8XP0wddYF5iEOwhu2AoldqnMErEkxlSgG8Gx9SqO3c3qLVgDRJBtF
b4X/rj6K9ceOl3DmGrMGaR8qOHZsuhzsoKS83Bv3IYMPM3t2odusyuh9s2iS
6PDsYducyjA3uaP3KTDX5R87YFx3ppVs4sAfKaFRSwfQzB96IehnLk9DqQhW
/7rMGDNKGCTzJYwvQDYFUufrvrg/I0yXo7u5Vq7VSGH2+tFMhulb3XyWp9BK
hAxBAHYZcA2LoaifZvujrIuc6g+u5P/m3OpVXLt3ECCmVtepM5kT9n2UUj9q
+jT5dE6y5ImPmEqxAIz8zbw0azqeHfMf6ot9hslBgCDg8J3/FiDMXIg4Qr29
m2w7IYb33dA20fJQHUwhTinT5fsfx2mTr5dqOoX5rB6XeBjQwnUm2WFkJN8x
nocFk6WJInIyn1msK/mDOAziVLbeDVWgBLFzp4cW9E371auONjdDscK4WHXM
ffXIJBWnqDFnH9j7VkviFmRq188xoCGr77htP+JDZ24rplz5xmaIJWUp4cTe
6eeWYpCjXaScjcjv9x1mGvV5OscOr+3iHCmrXx58zsxWkQ68eraiSxxSLHF+
UKqi9+HPUX3XluAKGVutjfzI54DwukVidGrJetaA+pL85CSthMNS+S5/SmzS
MYAuGPXju/MAvFNE6Oa95e7U0E0hYRYcOaxYpnRWy2nPtaSAMy6PKGaRuvv5
zj0KHfRP5KCIjslLyss3VtM/SAAWJypPU4ZeubFup3R+SQzhBkEVvHm/8pkm
RtRUuUZAUXGOpISZONREZQWzHpBH+jHbOlHK0ueNq1jbE0vrou9Ebj9kMCXo
X5Cod/OyH+ueYumvYeJXUHGobbqrtAxxDsYeHbhTwZoYqFJHcIUAuoDRCdMo
qmpFT0gdWDGgT6ELDxBqeuaV2qB8YZ7wYMEwL09yfADYKhzlZS5+1Ze2oAZW
ezohJz63l/sYbSGmFSuTqr0iupqdEYDuRFEqwjnGp4ymDzYs2XCfD64R6g2+
7VYhXsaNQZ/yXXe81kB69yGBrSd0FUyJFzZ12YJZPrH0gTywdZgBMwfOzYT4
uA9FuvrNRFZc9/uvWX/yYFKFY4sfcNhYl3m7/KRa9ECpTpaAlofpl/dxUsyN
drSzNgoaNeSTd5tRY/CYgKGBxTtq8n35jvBr+ycoiWApQ/h9afxQeoYBb/a9
mtZ6G3vgXVm59PSUTJ1g+MBjFae03N26OQL9VOe+qRS5wjQkVmhH6acrfizk
TQ28PuPZ7ZAFLjGo3nRrjY3a9Ll5dcGky9kLnV8leE3FgaVbd26ahAxORycO
D+MFucJmqrurlsGbIwiM6s9rwMy821EdU9OcCRf9gfXkJMIaVpc1G1QtfSzD
4iRLDDaUJMVNPUzEmq9znLzhzon3WTilvC/bWyT2ctc41mERT6leMFk81RFI
VqdzknmQ1QT6z0R74qySWeWvuMPKJyCp8ufr0Q3uIx86vd+pjCrC97GVflDw
cgi4tSuAlK2UBQa5rmbPZwXwNsSem76gqss4quik4mxfotmgHDkTSCNpXTqy
v9Lm5U/jBuhvAjN/ccnTEEPRfqIf7+zG5cO02XBNnHXzGvJDFb2kLGg0ZPMY
cRIeMj24iDnMG4tD832uhnxP1lrwzFUEzhHQSFy4PWBq5B9nOy6BHu6CaI+u
zpx2s72WLF0WdRXffM2a/JFhy5ejDjRuh5yw7PmBSq9GJiGD5T+I6I6W8sRr
tMCcpLBPPvEA+6rkIyfVRiV4qDx7z8Yt1msLx9EVYOxIQi5BNllUxlDsgYOZ
JOUq9BCm6AGEHH6e3rUobXdi+D9AAjg9/PggG5Gq/VGN/814lmipj5Q7ObgE
57XZvlQctmCMvgsSvXDamas1d/Y9OrAO3Kt7AVZfgqHjWFa7verimNux7U11
XgqgLqheBBy6f9TU/ZUpQA/7guD1pzbFc4vwzSTfjh3rRwAxmZZMvdM4LxoM
7lAwEGP9uJtowFxQzaTTlYfRjSGc8lhTNTFHITJAYK/nLY3vpBZ8+/zC1PLQ
ycAx5pZ0Asl6mXfqm8t63NtdJx1jMeXiIe64gX1ElHExSGBcud1bos7o9RMJ
tYNT8qX7+YcqJ/GhSMJdsbJEmU8u2a91Y/PCO8tB+KYXWjxM2ahexz43TrdU
crBZl/SrRSomaN7gUHwxKuCmekxv/PFtC9SeK77hha0BkPK0+0ggEVzQ0G5M
o3vaNNhsiNOlTj9x8o6X8pW7Ba+J6Utz2g1uV4YGVFZ2vhY0diQKJNu3flII
W5LJ3C/yCAVTEXlpnkfn3bUyMpfHKnagd4fbKHJgYFi2LVPyzbqx9y0e1+NA
b8DSNn7EqDjP0NuM0PpF3I55cEFo8WIdPS5e6s4+thLUNSWocapDi06zq+kf
px2EpfiEffRAhOec8YWBWypnh/amXNpAeYLBpVtfwPI7lH1EtkBdgu3jJE/L
721jDfjxRmKkBUEI+/2D8sE2McUuSt/CQlioeX43N/TbVpiDfVHLdO+U/NZV
abzY94UpKvQBQMi+sXunVakCtoQiMOijjlrZ9gPOrbV6pGf+IzEmMOxXK9G1
S5hphpjeoEL9v2i4Ex/QhIeKGRXAoXRvC9jQfBfb52HZenZcaEdM4EntNpJq
6c2mJfgQWdPy98yhLRoi86g5eWxikaeZEFyDgD7bFPq+5bGoUc2yXHwNrP5E
N3XOQSuwb6Rzvogso63AlMibEEOgJUKOgbQMYdhnt04wTIFOGw7ccJrbpax3
MAijrSbOgEuLiELjYXwEZpK6DjCGH3ZJmOr1i1yxvahN1H5EFFYmRVqNd78E
UdoPI8rPHQPRIVwEicDWp5F/mAYIqBOCcDs8e88MEGGBzG1jukr/ZQs1DVy4
G5qQ6djwpKxeDuLt13LtgzZMQISMp7ryB2lYe3VDkwam5Lt5ZzwQikrWN9NJ
6mVuzXABUmCIw9f2gocJ/pvF+9XU/uQvDzDumZ5i1O8ON3pvgH78xEm2GJeZ
WTajnGpb87D1YFvSWaMW0jxgvkBxJNlSL3BiqaNR65RkbYCOzDnQ+/WJj5Vs
obkK6Kd0sMG1JLNtPH7EGgZwWJP+BH9YPhio3PjMK1YJR0dXT+nUjf8vVfT7
B8mMytA929cCvHfTbbCyl/zyN7J3CWSUUSktqE/rD4PofHSBELBDCNUdv+Ty
lGKxIAuZ3APEsqwLgxC6nFblqHJnbhmpVGRhIZjismEc0cy0hkVsR8cH1u9a
nfd6Ho9efxqxmVaFWFtny/qd1Vj5YI1cSI1Dd/U0NCXnYJgLppWJbjEfOMF1
DHdd5IA4H+NQGXuihpFeVs44FFyOJYpf5pLMHPc1gaGYPD4SS+8i8LhJGyMn
gocKBvMa4L5dlbQ/N2OoVB4rMOH7Kyotr6chsioacM3sBblNBxV+PdzEFFKX
qqS2m45qeRES45fwIRIXFdWDjgy1N5z3sLkLhXCixWt5m7JSQeX8v6hwVSoP
oT62QocFLqPeH3cKrJt7VIcVuXnBFd8txXYo8+GEgHVyDxXSOZjoyAMI/7Zf
OcHnf69bvn9PyTmkjygWQuazh7zgoV4eBvCSZEfdvo2sFUBuVOmxn4wKxtsA
prWyB3e/aBQ2zoRDZduZiB0U3z22S7GfUXMsBOf71tt7I5HPxkkvp26iFaGx
BXH3Gihx/87vowQaDkhFB/OAuuy96sERLhnq/zeVZG5NwiDvUJaMKR2VjEYR
aVcNFCWnqqCIXaR93eqr8istsbloFHsPk3tiGqgEiMpy4dJDsS3+5oAaIfpW
VwRbccbx7Eg420+JGl2OgssXKcmhlE6X+SS90OMJvI57mlJ77J7Osz5bjpDF
w0TrRDVahj4L7dyIcEUfoHeMvvpUUD7XD5txZxCvIL3FGHBPabZjHZH58bZr
YT9TT1hiWa2zLpF65QZ2ojrQ1s7mtgclvFpZ7PXZsyBQVn+6GNX9K2rZLlOo
ftkud3/dch+syKFjWVu0QUKtJV1Nroy8qQmAOJqvw438kqlLTIT4FEw7e1AZ
zLFYS+cjeorgDD7uAmjum6psm0ub9mQckRn78VijedcoYCGQQQpMAzqnVLVZ
OVu95hlQHR0L40zOjlpA0IsWNG4soI1gg1z55lfhhLQphl+TB0IgdiN7aP/e
U/8DlGDaARJbxe/UK3v0CSkwPwRSinQDMBWcNBghv9lczs0qytz7z5zBhsmh
tm5fIJy3HRCPZJHjquXZa+ge9ET0+NDlzFFcLpztk1k0k/9kVyvM+Li5AIbG
IN79s1G1gIyheLruRqZn3MmID8CoicI1K1pWGUosSb8/CY8uSNM4sj2fxIIF
oyR7Q4rgoqpyCXuWxkVzp5Vmzrfa+v9JJzKlh74JP14lUWM4sqN8Tl1oEFJ9
efVlbYfjlZH1athJXYi7t32FdYd5fDo5LVa6VykODPDWM+ROQVh9Yq3NyKYw
ItLUaxVhV+5J9wb+reZQOhIdVBD1/Ou6ontYRvnb6PND7Ag3aE0AMfrWwGmW
fZ4AFqm4hhFXG10baH9hbv9aABBChUs+B7MjL+cI5M/iVwY8rD7thkEQvBHj
0mnDd/PPaCAHluJ3vTubPKZSPWwSuNJ8xhuVkNVFPcothPUuKhjkqwCIrE1o
BQnAcbElZ3n2mXB8BOKqs47x9nZtEdWq2WjgtDf1WmQZi+kCo5xc/OmWmEgf
zJ0YnAhVqKFY9SlPmufeCFvWro+ugl+lb79/ooubgc3peLYBae0pJK7qg9ym
FZxxzPBX0AThsTRT+F+5xIfKSZycT444u82dzQAtxU0YgohidNpcp+08Rb69
mwu/X12a++tPoEawsC57H4l5z8yPQ8u1Cf+T/WOGs7J21MZeburJt9c7iwKg
zRvsVkJ2+ZOddibaC1PeA3JuytpqpXnO6vnUOvtU7lumIwGE7F1MtJyCQZs4
IQoFd7Fa0cLBdvAddW1wC968I2W4YcAUUg0TvHUv1gFTTKjmDGI+bREjTm/C
yzwzDgd3cHc/R+9om1Wc/eH9tjjAO2ohhUE3eQL8VsHtuVPZBO6udtGaBfpJ
rXVvhml4Y+BUbKUQ/kAOfaHusA/t2y618tIqZqKOxTm9yYMGiHZdTIkj01bt
d4v++3eMlAPivC1o6eK7ExpK3eiQEIRylqMKzgx2jk6UILfN+Xi/yaiA6SGi
c3z1Nk2UiYdyKIN0JZl7o8C8x1j8dojgSXpVAIOWhwqvOgROEGJWzVA6zrCY
TwdFTJoSfSmHrD+09UzUett1RBVKxcrvNeh+A8nXZnJ+G/WAJIVea/Q1ApQ8
Bw5r8OPTki64DJhMI9VT/lHhp8uSqADB6XwR5+kk6BcFwn60zIlAI5iDoMNk
rs4gfuAzdvs69nJWj0JPLQaTisfcunkncEco6NaH5wqwsLSjEcqfmM408hg/
gWRv/TPcQ6y3WoechAxeaQQP68lACR7H7SrSVSM9cQzm8G6ZwW3MZe4IBnih
iqc/HiGtt4tH7pxao4R3E3pGVteQYKPWOz+TlDXcj9jwMa7G/GZOj0B0WP/a
jL7UIkb4/oKssL3ndQjGttR2nosQGe4SsObrEhxM/o6YHBB56Jw/z7/oJqRR
e5HDHHB23VnxxNJy31XkgjUw7ZLyZtq/PW9R7gh+F1KpQz7b1LybEUhy7lLT
J2EWBjxo39TzSjX0z2gOt4A6I+OQ7VH7d6P5SWnrn+AMI1ypnsnqFQkghkUi
8lqGBi4+YrvYuOqmyU2l+S1vNmYoPh+Pmg0aKHUVzkxXbj9f8BHHWWPiylZh
9P1tHqaw0FL2GfD3j4M4EFwygry0ulEJVIpysTEpDLqJYAmfhtLozU7hBa3i
j4Pwg9fBBhYBI1psU3Vv1P+Fh1Drf36J8F6FTPCAZeX2ISIWcV8WitFL1+4S
o8Rh6pCLCQmrxR5dxqv4fiFmM38V+VVO7ZRGttYaFAQ8NY89ShIt4ATVzSWV
Db8kiVQNlI8bqtzdmiVy2K9Sh7blD+S9Ek5TMRL+3MP+Ps5ljb3TV0RVEc/h
RhcGYoRD+7TvrBEmrHicT6Mn77v4MB8YbYXelIXTHcUl9TXq6g2HuDGkBci+
R3MH4P+FDfgdJollo9a8rKQpF/JH+gpm2FAn8m7l8Q1X5oy6F6w2qT/TNZb4
sevaYrwNqWnJPCrbW+N3HjPPairHDPxU4/8iTmP9CMMTgKHw4E3M7qhUWEpq
j1HHeIGDwiWIXORDAZX3w9FO9OV5DaGE9WsHJmiaAytSi9oIjsfNMJyfhqKq
gJxaYDhsFo4d57X6oUR4WD00NEOpudA78gAhAzLsZP73AYGcoZwdtEUuA02k
f7vOZ6EZkzZViQDlaDJdwnaLv7zeBD4kRoz0DVZTbtYM0PzzMYcwvf0OuofS
SMTe19ZGPaVMHqnltPVyBJa0LYhtSfuo90VL5tfpQLd58v15nn2Imi/pgQI/
xiy/+39p7T+pIxAFsF4bmtUhJGBztDgepboMzMyMvLBo+7oP91xwquuTl68s
NoXgtCzOoc9bQTuHI29XGCUgrj9pT6fhxbXA+AJTyYlX+hhhcAkfzucuFZUL
gzDBGOpiQ5r0CRprMgdrZzDVznbBR3eDGHxYcbXfGDa5uRXp5D1tEoPRKcXa
EGF5Bx0BXznME0ieS0EXPlFM2xs7vCLP4HuWxybUo/ssAdBTM7tbynedP8Y7
THLOKTC4BZFws3ZVKzzvJkuvpA3rJMiDnof8v8eZXr2bnzZXRGsffoPMCRNV
Kd/NempCT3LfVM8hkhF46otJ5Uv+NEmVd4VyU79lmCxYx5XXBaCQkAtsv5Dm
NTe+LM++3OfKRQBILRnPFN7dTCtT0xZn9ltj3HX1urh9TEO4WR7wgkhkvTMd
KvINTgKRpm4zbpTXz2BxBJdFZaLC3sYVvy0CqwCr8IZZjyG/GxopsEHDJrQz
4cHLLmpsy7/G28X/LpvN4b5HNltvlPOp8G31hFgb9i3WMqO+ut/nHfQeuAJw
2546p9orwzKJ6ZuzB+dDYfcVXrsB5WN7DpIZAHbNR94Pw9qu0mKfYYsvFVCt
S2LR8/OJxXv4FcNSn0zXJP1KdigeZPDFZ47f+gI1lyRRPweLL5t5CGSsjdrO
6tILUUd+AJrqZdmrAJOIJZ2Uh2kL5xW5AFttOF0FIx3/tybf0z0o6snFiTow
N5ZSHNgEUruZQNiW/pvXSqjFBqVHPgz7qDNO1AMoQGaoO8SZO8+G53EudIJ+
rnZDIR8fU/mmN4mjWss2NTyaWRL12T9Xp7/sdjit+YZpZbY4Y8y5mgYCCaDz
Zcso7gRDCZ23luHyXTlzCTw4TVGCCDnGYmuInZ0BNyfH+oBQNUox7Fgl4Z5E
7yxCxECCowhA9w/XFGLpb4JY9bDL6GQaiBqk/ypx7xJxm4/sdp1Hux/vBhty
Bmyc9/9Q/JVcGauPQQljPRya7x3m0sqGR0SJ17WdshXD7maRJJiOrfGywxOE
GPJQh1Vp4e8Cf6GuLZAeKhinmY81DzgxfPZlCKR4D2yTQSWRjjlZq+uhBRgq
ilFMmMjTCGAGEGzVX2t0889qycBkya9i3fj/YwZiC3fKhENy6SPxxCK5SlQy
jEzfHIVkBCJfuMGD144hDQHIm0ST6lbh6nXu9J/2QItsxo+Uc2GQcQtsJdnX
cm0kKtNr9/4GrcKF15KAIos8h5XZfZo1tmgf4cETmNcVzw4dJNsrUYxfqZJh
Ogs7JxALQd54pQVAMFPL6h37ylfneMlUf/lMORrBAal9dRo5BStKEPEu5giB
scEJ8Zh4gsRtey6gQUT8WuWPk6hJsswVFukz683oQkE0CxkkA0mGprhc9UGn
B8vlEuVbpHxkKjUJpqbLyoGPjmsy3JS8oajvPEXOwFaGixf81agmjpgYTm8M
4EtqCcriO9WJ7azu+kg6LljPFxLOKqg00+slVyOq2D/nteKiqe2rAFS+OeqZ
hYa9CUhtIfE008N5SbRtCPIPkFdsLsZc3tUbyz7vrk2wwHaEJ7O+o6yCeGCS
ywTMdyTZVPGfErRVwQ7uu05Be0GV3buE8f8EST/gSWH9sSjFb7dhFXfSsB1w
hi1k7fksjMsV4WWmRkI3c+6W3enCJrsRg3TDGdFJwMpYBcPxerZ4TY23LAG6
MuF2PEltkiHzf0mXpn9ooZGpCLnxV+KougNrrn96weOMibTnhpb+iiwvXaQA
msOfSQISZnWvwWbeHDRwL0SVyrEz/SdnkVswx0In+c8M7kOsNjEYYaSWyEfa
O1AuZsx5GDaCfDJYRc7n3uq/rKngjXbuKoqbMuxlV2XvOsugvwAUtbPOJEW3
R6Hg4HtQGH38deHcfRPH2G49/bitjj9t1psdMp/EOjF83lnkLyzlaNu1Ld8I
FW6q/8hzf0pBaiaBa+sa+HMOFBu2SWvxiQ+AA4qYc56UVxnmsQbpJxDMH6Ml
jM7e3g0PK5nFnnifwyTzshg7u7uDDAyiMLN2+WWWf/i9G/QrgQg2GQX8/CdH
8/XIHu+io4wc0HJASLK1U3d1slpeBdzvzhNAMTDUFlGdPespBU/XrsHXFyg0
HCic6fGnhXyhkhlOlue4cL6JyqhCnHHD7zVrJ6iOtQnjOqV8z5QrhhKJh3d5
oald/BxKDLU/3fjWujN/STbqUQ0fYBFBESxZWwuSXJbfrXqdg2UW6R1brwHh
JqJIcJ3308Go9Av+HSKdsnfCW7uK+lUpTmf/MWWQTQjpEux0H7O2UJtV77Ax
LFk/iz9a1DdWGRfA4oj2Q1DxlB5GKUjKp6PrqsouoqnzaDZTzMGNOTTqGPFt
qaWOLJE3GdG+5SmCroC395LQ//ymSLwDC9cq6pi6UMO/UKollIqQXnObgN0f
WqNIv+Pfl5qqNk+qAkCETDGa7JEtekE7+vSlttE06B5Hlm3NFjlj+tlT3EkY
Hwtv5f4lEtRowkwZUONhQbjfFe+Jq4q8bCBdPv6qNswqIvNDnl56hJ2afUop
bzYiM3cUrjqlpXoXaXQc2sEy+XSA/O4G1f/P+sCZpmbO/AA8yYQlICLJWA4B
WxpD/qAcNhpqMyJPp8YIn1auyLiJ4hs0tJIX5+OqW/P9UN9H+trAJ9K8S0mR
iy04FgykJ9AuLLjmwUS5dA3aJ0iIPIopbnf8S56PhlBTdsLaOzrymjIZDQhJ
XGJ6m2NutHOSjo8GpeXPCuTigJocBRYhevqUTb3nsoYIsvJqw5ToKRywD6pD
hAeWxmDirJJeKcKT39JR7jNyo4Cpkk1vJtcDWMrLjU14d2dW86P5GovXWsJ+
jJQ/n0UBqm/aiy+FZFx6TDN59Um1QyYAbOwg65WZFC2QzeOr2akFK/nduyAc
VckEZ34ryWjJMdrWcdFj54H/OofDBpzfR5Z23jMWTYFlZ/kRvkj88YLHI4AB
JyLf7xIHF0Rh2HwxaqQkKLpGf4pFZ/ddDRoCy8RVixcFlXEkmsbh6PH4NROM
XM/4YKo0Sr7wziiepboYgD0hTfTOcBbub167DQSFd6QGkT5wegikyPAISypG
jbAFfz0a8sUr2OJjBOMtPTVap1GsFyM2LzzAZQPumWYNocz0pSzbzrMQDc7S
CuEDI/w8j9o+naSe+tvZwZJRmRN8ZBg+ysAyowbr4galxucVPeVqhAFZz+xB
B7g4IV7bzORmCRGtiBafx6pworbmJpyfzc12UheqdvBzM/SItEtS5QrVyzYr
1PN+jSQYBGTrL0ZnWy87vvZZPDmT2/sj3c1ESSihGkuHmF+08zqw7RdvZi0Y
+Ew6RXMgh2/5BNx+lgSm9XJMavifOsH9Q9rcP2BJX6Ip4O3VLk6iGERyjv8u
KYGA4d3mlqRwDRDIZ2iBOVhvDuR0blRAOr6Sgju4Beq6kHr8q7wzXVmxoPEW
2BK2rpBe6v789mww9jH8vg1aorxTV6MknxozNzH6mVWOf64rssleB9Z6eaQg
a5Gk0iCv6TbfMCwvu5Yb259PggEjOvTtNjoWrZ3sgdgUCARIFofjFYNEL0Oi
KodCt9kwcYbxfQ+y7AiIz+3ByeJ3wTWuy+mgIBIfUnGOmMYBPI5CRnVCO7Ex
zdngcqiTxrL1gz6BB6piTLgdUT5coNENps8rC1+Sr5gFQ9NCAi5decck/nbJ
blqWqobuT+xslIZV5wCbu5Pqa1UHXaiUHvRp158EI6DNEl6z7Mr3VQuuANFX
YsoyDEV2bnZXKF2lzVO9l22Eev0AVWrCZHR2fmp7ySbT093cNDQMhky5nfGm
8PB1FWVKPPxsJhkwNDHsVKL7jxFPPz7p8eTpk0V8n/kINMUxJkE2pXmESiFI
MOG4oWxhtVHXjK5zZEEUm9PeDkPxW2OIuDTQbabj0JXHKWXDCbTrLnKubDQP
nncAigSE+n4jAZsw52cwo4XTAnqSNlqfSkQbEboDyLNrySoZj3QTW0tNQxds
wBG2JEzc2+x4tmReHasMUYrJ0iIs1uQynTGn3YTz2kcKNxlGSIpwKBj6nYzB
bwQ+yGEeljc/5dnkqjlAfCtCKmF0cktABBhKYaH8SfVjZ3s/LRiDcAkFGH3S
W+/+mMjCCZtb3eUerJOTllmJ6sK7zXKJIp0VMp34mxcISyDdC4RI+D+swOQN
MQfIMal6yM92zPXvmjduhYpQzjO3ArQoUAVykKUKgxWF6Z9xoBB8++HhOjVn
wZkAkuyWz5i9Ui1yX1JByEaf7iAUPqoXt/70ujq4Pup7fdEfiuGmL7ae/6j8
jMf5AsZQSfC+gr6P2o11zfkvYuzeAy+bO8phtaDVX+YgAEjXjhURDPVEGoj1
A+8+EVGZAfvhPjTaaiGWgpY26kX+LI3yP0RpPoKdYB1geuEN7g/QU3kg5gNU
mcduXPkINe2TLO3uKXlOG482g2O2V5kOrcW+ik3h98n4PnvlPVpjfO0tFsbF
FjY62Cj23hgLb13RRPVbWbGsxeeuksxFn7FuicZuStUM/KTR7uZvwdyxKYbK
UR8TL86eyePYHGpSscM1hvgihh1qfH0/70kCDjUmEphQ72Ir7voQ5UUJAmpO
N5SrRmP0yU9XCmKs6As6fL91VoiRg/RDum8YntlG14tXybj57RTiiGsyEtWx
LOw8cYWjsSPS8qoFVCUimCT84+NXqXH8ebCU4pWo/MNfNgCsjM6o8Ny+UsVj
AeBjtYQdWaeE8tf9HltSRO+Mairkv+KpDomDERoVjBhn4pquxRcVaMnOhL4V
SCcLHbOUHfd060+rhCFdSesfsoa3g1X1EwPSevfKqdG3C+sElrBfieTkggQC
vlB/6/F2JUijOwL7WtodNaCWXNMELvTKU+nmbgEm0L6KIGHivvclsGKJ8mML
VWI8CY5PDGegiHWzzS3gX4SYpRoA286xOuWQodazxEhQnh3LjsDFKxBnqbXp
uLDd5K/cqKX+foKgvcYR9QvL2Aql976mqaIfL3/0mb1NRL5LPO+5hhgKJWT1
52hjt49epPwUg2bcA3Ief0WYOpdeAFhg1c7+NVfXSqqoe3VbmkQydq4Ncl27
HDGq52RsR8ka9FY6AJdX90SshZ5KGdNOTiPnfh5O3bDai/HiP+vLOP3+XsGJ
xZsjX4ppTkC4/9T17wZnPhjo0z0q+VWj2zUG9Hp5OmK9A6E4INmvZn3ACBdA
2yy3KwQiZ/OZFjQOImyfKMUJTkkr4j6ZGGMbd8pkE9mifydL0RPhuIy5eO4M
n/RrW7sCEX32RIFr9v2jyWBhi8SaqBQ7PPQGysZP7uM/7ioQ/lpU4nYXrjGq
D+/k3XP+pb2jkLxpD6CSXDMALxw7qz8oBtB458TpIC388uwYFH59CKdzx3vV
w7TXEmXBjuJOrdBLtOmY8u5yVr4HgKTk3gZUuYupxYb2NEuUK7o+fpfBUjsn
x1xLjCiAp7Ei513hF16ix+urOKjrvGsfqkPRHEKjFWHJHMLmx2E+RLvbbCc6
HCwu0A27YX/fnTn43nUg02DYTS/WGUCaf+QZ9tfg6Sj5M8o8AbG53lZv4Ezz
E/Z5eUtapwjW5kdKcVsFEIzdNNS+soOXc3zWeK7XI6D2ZvLUqW5xgXZETjea
QqdkzxLDSt2Zwjq61PeXe1QP8Y100/uWMfXsDMTRjWWDzipjIGyQnQi88apA
KG1FddzxmxNmCOgLB1zI0aZVWJs600SP4KHNvtt2acysKk+nXf6FWOoM2mXz
ibtdr5xfFA93wjfWWgKQVLlOS/vJ5g6P4d4+7bJXanty670XOJL4TzqcBob4
2h1tUBmRzIMNcCcx1Yq0xnGkSTxquvR/7UkVfzbdy9tF5t6xfNDtOwvpitVP
batUbmeSyeArTyDCAPJD35tXt1+nB9sqE+1ODyzdPK3QUP9MT39iliKQodhG
cxvVYqH4Z8F3NI01HKtBMLZCBicgUuTl6/aaOIyL+Jcs5af4/2+kOOCpLrK5
DhdCL68Cx6JwVrbjQY0soRYR7tS8/Z7RiojHPuQQfMbgvzdasiLc2H3/Id8+
m+keT5hCB6UaA1zmWSgupFB6HzTcCZ6wlCl4gkA/VMumbEV78sX1eRKidrGU
EBO6A9KVDLa+LkzFdSd/zI/bH0L6MTVJQrI/2aiuDpQBNGVqSKg+a7sgFZpu
LTB3lMZ9sifePQbNCsLxTfpvMsffvZh9+igMLRXV9pA4bcEwAadOdg1eGajh
dIY9rc0C/9CeqZNn11T9psIWS/L/suh7UkQduFTS9ODJUvvQXCeyzt9eTNCE
sY7N1ssJ81sBR60FKo0vwR9AGSuts5I1Y4hf8F82d7yIWOlYxuMLbSpnX5Mx
ZmgsyrJCdTheJOROv2qiNwRE0GJgkMSa6OtNcSVdkqpbiOUikforvClj/5dv
S6TPhIqH0FSWB42vljrXNy1viEfI6nT9yhwK7gb0wn+PDy2wkn+GGc/k75l4
fjzZymkOBryu35xSFDpK2PVSJ+Qw531XIKNeBR2+1ZgFPAZkmHGDW/4oCh4c
wO/B8/DNfAXxr7U/D80XDdL6oYsnHrLPNvH1Bz2JbpvkhMgoLi8Vrp2m8I7J
N0dKGnOqA2gXK6CAln8+hYg4SvznvJPaAFcVFjjC9BG/OedOGwgL0Fw8WSC0
sFYDS6JXFD0NMGI0dJb7ewoTyPpXC05lUlf5IjQI3+Jo2b5L2v98Z1huUHQd
uqMVWt+b3oDSYfc8we0OhJgk4QH4m3lp4Rykf8hMsN/WjVQnf103JAO//uok
YipILuBisYPRfY0ZbdFaKWkfo19zOx33Kb6Zt6nI2Bu7yqNAg79yHEhafOWR
bLAdhpC81upW+M929WMwtbP0UsixY7xr4SFQU3dk4KHTrxcrJedZvX/iGy3V
2q+xBdYdQ2IwpA2z1OjMvisojYm4OiQ9eObMjqe7fbB4KtOuYd+eTor137HH
IdF0ItoFtnBnGxDg2EPZzMVI+M0TTl0f9NQ4RcVdNXe9SYuE3Ie054B5yDcW
mMMM7T04RERIrklR5mAVeDvsKHepvfPEHsLl/r8lubcOCKbEgxz0qRdWvjCp
+OPzPVpnwTMxX6PJns4FbKgf5rbAyjUQxsYlS7dX9j9uuPGX0IqaeaVJfZSU
+W/N11qAnpg7Z8iYobkQJMWr7EVdZJi1WpuhVcVegLPop3NbTSwIb9G9LP60
LRUdNcmSPxIs3MR1uz3B0Enf7Cd3HO93w87zxaU9ZjigaZa15A3xvdCnMKIp
PILKpIcFf16bGhRUu5o/bGvANHkIT2OqFtVqguxJsjrixNzlAcix4e4AOSg3
EYAT3D5kBYHzeuD+2JYUN4s5CM9k7I6IAzBB9qz7CuIk6fN7MjSF5eW6BOPY
v0RP1/bpJ6ZsKgFsSqKLgUKrxIxAHl2eYOTh5PBBCw5lt3G88ez2y3rY1JAW
TQNw/t7PrBZZVOeNrqgTNKSARmHTIlzQU9nJhZt7PuNF6o1pFS3cxt6tTS7S
EzqC+r9f6VMoDMEvgU/G1YeE0/pWDTx54DE+1OuwR/Da8nH1fDoreR7E1V+b
x8+ZTxCpnlfl0wQO1gw3lqM5kXJhNluCei3INObekzZEHrrroXvYfg2eA+Pc
SoNj8F5oKgBcbKYFYSpzAT74jl7te8HV55FqWh07fe8Bn8i1THk/h5ic9zKx
G3Dr1WaFfwD4R9lEa8xv57c7Cpj3WfIqoroafiRXtednISNhLUDA882tembk
VMP7teyH3YDqcv3uyikVqIEeJFpgskTOVWm2GuX8ZvemA1+pM+BU4XVKe2Uq
j1hK4Qerdkrwvu0I9NBbwY9kx1CI1slkOWIBUOiUqvQbmE5aFjsUOO993yCE
eThQQYx0PgfXlQrbhgKGB9/vkmK6Fd5QiL6x2FaUh7JLnXVFb42+sMU8b3t+
3XmC0buebWqKmh4vCbY+3mr8aE6zFxOkDfd0K5ywDYChP0U+EeDy4NCWGHrZ
FJgugbRTyN0BIuBn6k741xPAFKfYO+q5PBsMbvl/+DuVw24gMADGZn0tAMCY
8opZEOYUeKhJmgex3iXt038L4U697t8/28icxkS/DKIlyZczOJLbrM0RG0hS
q2isnVt7/s+6tLMU+1CWSeaOouEjlhVvxB47EwcJJ91QzBinEmsS7A2PfpE0
AfgVKYjfF0VG3Z8s2Ab6kY/ipRqDglW9aMLcOZRATVCeQ3eDBctgDvXmH/CT
F8lNbibgM+OSkiyO0qG2+UOqdLQpFLyKgA7JYHgpyIxOhuHI0yQnYc35Gszd
nCtQd2uQYDn460EseHJSSGlCGv4qugeg9tvFpqNhv7K42ejLi0T+g3RGTJt4
qj1zyBO7sk3KRQv0YX4asUc+haX6DfNdNA+XgxSRKN68EPDqxxoEaRFIIaNO
EGJRfEn6BKAAOKKbnMtbbT7tMCK9zh2FunZw2FLrd/ecwc3e+xx0pqZwJyqu
2cVIcMa9GQb/XxNmi+UWDKDCR1a5+UPntE92hvCS45VMqY7cGZt/pCyaxxVx
mGgWe73Lpd3q4MuLUa4Bzitl5UmJb4BZbSY6LMk9t+3fAVI7A+Hj1P++JCpD
LIu/QrTzT04UisqFusdXnTCnFvpqqhrX/8PMO6FtAxkkJWSxBdGZ3lI8UY+m
73HsVs+zQG5H2SPD4XqnI+loJf/QwWDI1rAULzpzKiv5LJGWsJ+2MXh7pT9u
TbB1YhRbBIZBeOoIwb7u5lJP/a8leVzlf0Y3H27h+eHmgncvkNPlTKh7eX3D
WGeFBWNacX7AOckSo2nrq0XPSQvh36VEvJNdv8t/+/cJPUcc565vS0CE4Thk
U5hwdMuEDsKn/LQp2dRS0DJj6I5OXU/uD/EZJ4ceCAiEOzegzwGYyFuZYl5r
CDfaVp0Obc/Eym2RbQRXRRxaQjVKkeW8SqE6MtiqOzA88UI8Ck7shRXT6upX
pQ91IwIUi6CcUeNPJg0BWEAPm8lh1HM0ixKD92Ar7Iybu1VLzoaUN7Mt/k/j
lOuYGtFtuJMhU508hx4NdDjqWk4snS1OqnbblSI9LXxPGulPzIlu1ppH2uCW
1B42fnhC/HjA0ZCyLPUM611U3tNgza37TGE1lnm7ZVoE7xPtO5nU9S0f2EBT
Nw1ZKbPAb9z+E2Ismv+GfSur/YWl9+MiG8TLclU/KOo+gENYxOJ4j4oiDFJZ
faZitXLucbp2JCKzG9mli52DEu/ITI+JmSX1cZgoFlFuVvJTbLuVIZzyAY/z
MTr7ZtJn2xSBu4KovzrmvyHaY/tsnieYKkIZQgNI8u0h+T4/Hsw0r+3vzQLG
KUlfIoMOyDLVMZpd6mwQhGFxuaviyPXUTNlokIMJCCtsv8e9WK66nS4JyoOd
k4C4wsDQfsdtkUYrrDOda2Cs/fTopfqHrrWK7lwoDBmV3CKx7QHB6cIkhASi
TkI/AszPVxxj3FlLgDo1PAgeydEvlQ14H0VjV5GsK4Y78HbbNeR7iEn9NKZL
+I5/uFxhhzZ4uJ4XDW5/+joFWHGNa+09GJ+nHu1r/iqNOWgiQ2M8xEwMEhJT
98t6XEChqBJgHvgLbjXuf+sJcxov4W8vA7Fd8A56ypTJ/4vZ8vZrDow5wGBE
usF0egcSImaVCXxljOXz996ZSCudCe+FOP/1ykyRQRq2e9OxXMKfFwTO3/rW
C1eQyAvs8A6bLV0LZ2xGAGpDRADpExGWk0lrapEOJmUBlRPOkH6AvcLXtRaN
s4znoO6r2+X7cIc94BnQ5NX4qghAwMFqq0+2VaOu+l5rs6eWJMq9Yw5gk8yR
e8RTY8khxhSnk69x8++nDJOUOJrlMYZAAFORbsVbePUYhWxYIEr21IV1Bf6/
0HK6evypqateKn/iVi22dP66MCy0MZG/JjjI37j8WjG3FiDLpcyoG9O6aoXH
/XFwysx9YWoPU4ooU2BVqM+KGCK1XfvKXpqFEyYjkFzuCIhDv9l5Sk2TRp7T
OshrGOn1imJjgWSid57/DsX7T/kUfJn/DSYIlpZQDser/VFabVrsStIpF0ra
PiDFSt8n1X6D+fryetB8qVvHYEF6dEQUp86e+JBPhuJdizMnJqDWo5ZnAtdl
RmU2TWWRnyX3vFjTk9cM8CBUEEiRV+9F5x+TCHBDJynJKVt9COnhHLGEDtpO
FF3aYRiF5OubtSxu8kPtrPMKNkiM1lSm31PExhtOIomMw8q/PcX9YcK75+j9
xqszfb19//wH0U4VrGtBokpmuE+wT+vaX6FVR63Q4DErrjZQVi24hXmn/fma
KaPhTVgngZa7KiF7tDu+N9N4azEWdanyzZt6YENGYwUF9cxeUNUDTlt3ry2d
jcZ+OyMPZinM8GWSvxcIAFlRfto8xD7HvGnrp8oz1KwHana3Fe9CD2c/DLu2
N2XIABzhxwUxQMLRX8SrS5no78naFxPD5JriJUeeYRPnOur2s/XplQPKltb2
Vliu6Tpc7UGJv1nkLyWuO0FkH1Dxot5mHel7JkNytfdLvR/HRZNYfFX298Fz
eQquyI67Hm7PHEwS8ujBzLRWg0XkEemGGj2Rpcomue8ygwtcsmFNMP4nlDCl
90bTuLc0ClxXmVjkNN1dOOdYmTZSJJH5cfztXrGXXdiJq8/4VLh4Olij891a
mi5sMeJ/EkB9egnq0sOUdS7Ij3LBi4r0Zp4I8k94NFt+kxMdt5tkiCic2G5+
SAvSHKT08BmE/2aNzK3/L1uroo/7oWmOflAcnpaOKGI8dBNZ5bYpXlmVGYGq
uuD+q7UKccic4xmaxeewrVNdAQE8yZOkLSE3FgYHmM7nV3pg7uSzdwB2KtDR
Sh04ipbruA0+EbTh744LPx6mBwhvvK3Pzfb7OstkpLJwAGivumrDYjrAvP3n
cd72Cq1RnM3s3+GwOx0M6l7HSMDPAqNEOIoH6tH9+ZxHdbTIYHavt95gFTGo
TvhEmC8cXl6gYTIamyWDAFTO5B6IFLZrf3yVlNEqmayaTDIDLFRXTk4RmMni
BxUph8HCgL1axoUMIMVX7t1kJd/E/t12MJEJMTjqr5doiNxjv6jkmGoElSTY
XqsgR6nX6aEZ2/TvQiDzSgwCaQak+BD4qpFfYTvjskNRly3EMhKM2Jf1omPI
cNopjxJjNI9Ive+SL5QLr4MFCUfWuJB8IV7eU2/kVT4YXtD7/oJdfmrjLScN
zuZnKz9uDpI2A1vw7NoKyLLKb0TgkQIRz8LwXVnr+IkjfNLty/STC1P70Uri
xCNUegsE1Drvn14+ouJVL/Gce0LES4FVJ8BRddIwvp4LRz7WuExcScaaivAK
wH00KrspZ81lYCRfDerrS/j74+Ydq/XiRYmVV6tWGnvjCebRoSdEG2LOOyzh
m6jOBaQr803vSugs34NCqalMmPFtHFP29kub1sMxTMtT6b61zQsXuy3Mqm1F
nntQW+LVtKsuoAGRZWugNzIQpEMgOVS5CN4pJ8bXgAKUEtN++noxEbdId6/n
SjqbKUbJLgpwcMhzRTShxrGLkYD78QZMegVirsU7onPO+h4tI/SL/2Y4p8JK
Y6oUUjgfevcEu/sr8LtX1KgGq2O6iW8eZXM9EP9TUzttZe6mSLzedN50pIqo
ZBNch2t9E0rixNpVJbGmlHS+bAEFzO1QQs9ppz2WA+ZPS/ghJ0vwwt1vgWbi
e8zqs/a7REJtoBgpEFI8hLqL23Anp6/mAOh35CaGLTa35cJEJjjcKc7smzBC
XlKI2nMlrO5fXJtvzCfDCb21ecYaD7AA8ubU6F9sYgQfXcILxoJhfa+aOH69
+RdyU3DQvMi53gDhu28TOWKvryJoS3Qot+z3K1I7giFOnpKAfz/LVTtD+Q0c
+Zh0uE4ZT7X8Au75NEoX5HdEuwh9odkZ420C/sjiy/tit3fLgD4TIJUbQS/A
qYgg6+G56ofPIB/+l0cqd0JyKj3h72ZPBao+T/OkNZsO60KjU0jm9JO1qHgf
E6O/fh8Lg6kQ6UCGyBkWQUz0gc+AvZVL0GOz0hwtDqCcevb2EKx1z+pn4Uor
jfu3vTBKw8weuTaOIBlrd3VXB//eQXvI2yPhF//ay5wo9s53qEdMtRk46RqN
qNdabECesm2e0nqjDRz1VQGMvh4Jh+GXT1FLKK8Npt8SPQmYoQeKDtwWfBat
PzweUDK1Ca9PsVpaPEwfeHhhef3r+yHqpBY1MzRqw05LQhwJWOq0ycIwpUaA
pccO8oQUXUkiHel/v9ZTv6d6XVZzyMhcy4ueMBNd97kyQS2AKkBK0bRycvhn
xTRWbjVukHnE+pR8jE0VHQ2wOXe+4FeWqK9d8nVtq1xeucemZcnB9yubitmX
bt/Ntvefkk9YzvyccLyiXGQRtMhaFVpig/N8V9N44Ak6aJ11OJ5/5XIKrB9t
kEWVLV08nI4VBBKS26SHoxq/cNYUTt9ct34IgYpqS9HctCApW77lyUn/SN3t
fmXej/NjzFHoeuUC2m65XCib64q6iHyUXtCwPGr1SPWtUVTC7wb9tesbavye
BrwW4JxO+aTH6910/n9e9yhq4Hq6jYOOzQm/1dSVyMSaYIuKYkvNODDE5vAX
qrDoJ/cAUOVBbIL2slHQpmMvJVJfVhXIEcZDN0bSYUtBHDlWPxFMCdQnzbEm
2L18oO0nof0nnAsfUQ5V5e0DTesCdLo5EYAfC8EiDqWunmhqzQSUJ5RSN4UB
JpeiAH0xj17S1edeiYuPCnAsbEiM3UHrIBz6ihsJiH2tnsf1GgOvTER1NxZC
KTqHUK9glOIKg7ZgSNH3TWr8e5tF+JXXR+0NgNtyj9X2sbg5LVU1Z1+G4/WB
ccmruKEpTYw9HFtW1rrmVpk8pz8v82yCyeA5yojhDZ86DqHbx/aQvLiJp68D
JMz9dX03n66jkEiCvtxnX2TL2vOEGXlcg9ws39gLyzc8Xi+PmS5Wvs3Dgb1f
Lq4mzCQ8nz8jnJVjDFRblGsFe1/ceY2DMS+clnzi+dy/NB0cN3PMbMxtt4b0
7l7ay8nD//OgFe+Y37yacJCU8XQl/5e1y06MhgbIm9Xyf6Z8h1YPZI29I7ZV
16fBjn73ZzOs7U9mxgrVTyKho9IQ/u9rh9p/CE/CfT+wj/htoFSzqs2w7K6R
7MveEJVP9XqL6Sipe+O9ZCJwM+ToHUD/nj9tUa90QkUDM+8dIoNRPofz2ixR
JPcd1bw9SINUZk5UrFvSVrFtgIsk18eewoa0cavxWptoxx6uNA9yaOl7Sema
PhRO4eWsaoDbO9NTC34ZLi9x+lQeHZ9myGMoT6ar/LuhJe9mABDSH6W8nCUS
JbePqlQeIHH64p7KhFyEYlw/1gjYHTkYbw8ayt4L9/0M7mexgaSTfd10AcKC
VCWdNVAtZpSPKT7gHJy/hJi/d3P6i6E6AlIw7FtJB0uukKsZvTwnEBSD1Q82
riZllHbGaa0ushLturLQ3yVeZTA3DrSWLqgeLidigMQIg33PumOguQDn/QsT
NaN/bNYDPX2hStM/2pD3OTqT8Y/mdLLtSLjZLpsoG5R/ChN1oJQmud4hOCsa
s4ADzT5bGBD8SelSMxOrhBNI2KwwITk15c4C9nnSvhQ8F/tiaTTczQa+ZODh
2X0zwK4x4hO3BPuD/rSFjyJ92YNtQBE+CChvoKsyAWaLdFC0Kj3IPfNc3G/r
3hwNOFdWoY2fqSf1xRVvuKV0CZhNPiAYlhjLsHKri5fM+GHwo0UqE1ARpw6v
9GD9wC+DWeWOl/9VVp9abTCBWg7UDRqZTVFro+pGJAPFHerjMVbJkIdlRVeU
EYPsZfQ/PIWuXbaC+Obp57graLsAPMJnKAsuykk2lKz6SIjBmrFyTLzSKxHb
eyiUUGVb9LbGFcZRbTXhM5DiRYWH3Sd+xwTz0lW9CBZqQjXtWOaF1PHDNqn5
goGzH6H0T1K5ZLz8oPgfRvkPjrC8cLawlinSS27kA7IItyu3RMSBwsZ0+DET
38LDBYL699syDvXVoKPKwVPEDXACU7c9vTAKeVKD2jkeFyp/yHI1VAYTpxaI
vP4IHaHWVLfmiYoLd3GqpiIM7I1Dvfrfq9BKyB+PP+Lz9FBdek/4RjaLBgUk
tTQVsI7hBMqoBrv1RzziBvAZw1Nex0FFJiPlXiwP4X44rv+yyw+FKWjo3+FJ
7cZlXis5xl84zYRBsXwQ1dzQIOpsGxMD2VDQnBVEYZN8bbYyg0/tRzAYxg6l
KWmxSvYfLAtGKI3WRWYFOa4gd6lUEUd5CIkoZ/PFgUpFRenVJ0G6TknHlGWf
F8BpdfegbUdboyHOOqBXSSP6WLYHVCKRRXiKN1VKd0FzorDwMIWnz2ZVnfNZ
E2RZak0ZRob0ooUoT6ihbDD6qLESBHieonPpg0586L9Bwc0l8Mz4w3q8bcEF
Tf8p+5PVpynm8dZ79dsT5skx9zwlMJYuYdTLTx+hXN0qWaNKP+ByjwqQWhKv
Uzx26GdgAovHlYJlgl+AYI71AauU7Yc/YCtADS/4jfuSxRPDSW1TK+PP+Bl2
yk5anB+6IPc+FECRDOfxo91bTlCxlI0v3WnxPr0fD0JhmxrGHyHd6HjIjiWc
DQPoS+GsaO3RJMaNGfKL6JYEGowdqnMBy8y+MMbgAf5c56PGNG0/qNBdyS4J
BvIk89/7+MzHCpmg5UNWHZlW8HxU4k383YuUOd9rC29kRXBkMOrZTpBycuot
P70KjifmeMR95G95gbNvPOwIA8f4Z71bnB02vscoI0fn3J67Wv2eAPM/9Uku
IWtuF2sM1QiNZAa9YNPOF3vo3SxSy2qSIu6F8vOEwvplFnvKnubsTn9R11BO
11gbWzwYgi9eY+6YmETgl/w/RhAwQqr25T9x6sOF3hnBWicT9zzf61/Zf0YF
UVdZP0BbdXdCTA3QMNNJ6luQdyMzUap+R8bkkjdl/xn4MGzEAqvTyprULfyp
7VQKWEFRejkxLcQO8EF6WlxpGYSRui3SslZ99EAiZSFrEVw1fLFqCslc4ZzF
38pT0F8eae/WksOl+k7bHTQXyeet8gXD8+IDWqRs9XKdgg4cw4F/G3rJDdma
884BrNrZiolxpZmAs47vMgJ/efpNRb5lcxBuiAimvH1MiO8i/oYXR7KOK1Ey
rQ/bS9CLig1EsIssHCN7/FZvLia7OAGB9EdsBoqaQ7aUbEGcOt6sRMsEwLNU
snJiBUB+KPxidq4U9iFCw6E371cSIfKkCnn9Bym9w+frUlSf/K4nGTlURrjp
5Snm1M/sv0FhhbwMG/I1iPKb3jxferVOOTzYWu1QSc8jGhTs1uM/HLvG4E01
rHvbY9tWCgCttZKjYiuHsibizWGcz2K1uZU43Zt5+5MxpYt57gFaB8eWrNZ3
eOhAV1ZpDHkihzul7J5MhrA9aKTWz/RohRThTp+T7nFe8ZbmZHob57MFNDjT
g+1oNbH/bbx5uxANLaLbZ6ix3tnm3MX/2ZfgE1uvGmn0k75syHOhG2hD9SVH
ZJ77eQ6ZWAZqEM/E1hs/Ka3ISWXV6DEE1lf4HU0kkR74JSBDY6lraXmP3B6d
nVFwRIy3ODOCIP85xRFM3oOFLhNybKMahVtuem1bYB5nX/GoWS8x1GJrHzL/
SK2l13r28ZEeCHaBfQOI0JOGu792yuHVvfcw1sf+TdMfH6vnzFvuPolTn6NS
8AKbpYBvkQwT2SFcgy+UuNdmcTavwIiMqRyKzf9C+ZDG8H4gkzFY/tpzgvfU
sLCbY9qNGiWLn/K2/gKIxNAR6gnJf7yW20b9MCqKJykj8M1OzSe5NMJBNC6s
vnEBYJPTgvSEzHBNyOIO7kutYh0OR6Vj4QS/j43UlT8TNLLXlK95+u0UH0IX
gCrV1PoG3cxJZZH0lNNKDWVKgy6HlOBiIbKWVpAvDRwcCxo7B45bFes6XAuR
jgyVz927QkMGmpPzjfZ8whLgGEXoTVvrr43odDMYoBmEaGKADODL9d7Wd7NC
gxK+0pdPrmGLcAm2Lr063cSYXK+eZ4eeeKhNbSxZ16M7/hHdRD4ogVLZGuF0
McIYY82Aq1O0ngR6S6z+fuwZQ87lcrtvdN0ddiz75+T9r3edCEuSYeI3783y
tEFj9gT3Hnf4NRXVtC0xfNCIZ91wxcGUn+4vYss4hR4UTq/6JBAGJk6GrpVb
oZiDFwyjsLhwoBUBpRd6Ksn/uRF55VZpgXvg+vqrtSWpcou8vB9twc2yC2LI
JpdiZrbo2RppSJ9zcpcoe6GRkQ8Fza4sN4Mc0AYCDYoiO8sD0sQNa7arkJOo
Xb4uEWgjlBQq6xIb9RrDHwmZLejVrpsXILQ6boMvNIaaHsOhZFNsUot1XAtF
T4DPkyto+0sxTh/jEqqs+481hSnteHYLG05QdvbDOpLrJe2bYnDDt9Itf7GQ
rlUkTk6LKoxlz/2C/jLU6NfJ6Ete6rh4j+FGHKWjGybMy3sTruZDZsTRH0cL
V6qnLcNxcMywzbCE7dgdjPn68Eoucd8aDMOQXtNHvNGPtvWfvZj8gnutjmK1
O0Zoi3EDn23MeAzIda/fsbviDzGX/EP6xUofQdKmkJWEvBYJDrXrWFbZYi4f
m+e0kTFg6se0G7jxjBG75GNIgkqh12ZU2ttHPDfDJsLQM9OjTKQQqK0pqyYK
P66EJ22B/quSoZbASuIKjgcFGm2ceQdNrTFK0+HsdfwosbslFGZWetmXvQZ3
yFvtOULakTaxzeyuJRv0lcNuu90S84/JjDK/DWHbXUAeokoaKbEd0nrfSEPQ
k4HZSom4XSzwsp2kavuUKYMDLjv2SVNn/sginaeP/afIFD2O17vFzrbaj/DX
P+UmWxYiiSxPwkm28zrGzjB5kA+hcCngvNk/iliHT1cYvvd0fg58snawPHXs
rFQxEhbqq6cC0ErFQ8gmVlsYldoMUslfUp8JEJDUukoVyrepXe7RrrWXKlvY
nzhi7Z4KK0NnWY34dAxqbXczn4tJ49HuTFHL0OfV2KsDeEpOfgRYtTr6jHAZ
5qvyNWxB6V9jl+A/V9tH/grsadntZtRRT3S+3id7/o5a2jCOsv9Wp5l1QCGI
9p/TNf5DrW7EEA/iFJ7RDOkYE2ZIlKinRA2MytvZZHIN+Rxkj0v1U6PlgX2d
M6B1YTTNvKcduWNYK223vYFSTIGD6TpiptowWdmQWzCDcP1dBGia+19VGAW0
euRqGAwNOKFztz2tZOvsvlMygXbLjJ+Os5WQV/z92PLrcNvP9eQxHltPtW87
NTKJfAM2PbMUJaiLBs5cpUHosEswCPZQxW9XS8aFUeAcjP2l4pv8tVof453g
mIO+Bq2H49R4pnWB2tLou8+89s54K1VJW8SXB63NQmu4qu0lTgGi+Ypp1m/o
cQjn8GuCO3CkyZlfwCy/0u6bNluWWSh0XAn/AWsIzXi+8Bx/thEaogkFYG6T
mXuE7I4PKuVrKKMDB6ly3mEj9RCdKW4hyG9APoML3G8KD/f7bh9Xn3QKAAYk
LRiqHIkHj3owlBUHmzb06tjb1rhBhx9KLqHTluMii87ZFlVhzlT4X5BYCbvT
Y00YqP3XBZoaP00SAekLb9snOHjsn01FIRT4TmRu3RhjZ/DwJLJRprJuF2NZ
/NZT4mohJuyJe1JNqurBYktqM5YorJtKl1qHJvMKgJ54L6xv4fT8pxpMZ8P1
XVLQEirXtl8+g/SfnbopNsJ/MrA8t7nr8xhYHp1Q4zMPQTJ0Zl7B/hnaxMb6
KIaxDxMRkQqKk7s/0zgYgVLowDPD3eYoHK3cA0Ks+1w2QsVJqcWa9yP/E3Xg
MxRDQOXl1MRDdJn62MhUxFI0uZwNNRKxct1qE3a54PC/AUDBqel//RS7XMeV
uEE6kJZhfwSi9FqrXArODVYiKGvPJP1oDWefvm6KEkRaAKkF5IHFxKWj29Cb
/6fqGuUo9es4DiFOSQOV3Ivxq0HvT9c7mfILr5mU6ElZwtucEbyV5pdfmnlg
jc5frG/yFd3c6iYa6OIQ0am4y5eQrpxvVn8aDg2KQEOOVItaQZCGXtj9NcOF
LvArBvu06zAB8mnvx/TuqHqdcbpEZy7MiUSKZQmI+UqYmtVZsKdJAn665ZUj
lSx4xyl8TGVzP5pRTOi2UZt1Wr+X9q0yoJY0Ir2jSIO1U+nB5hBWlRUybt/3
y8dQruxAcSztQg16v9vZob+S+OrfvweHCIFt8i2WurwUbWRFieA95iVauP3p
WOVTicjsF7JXWp+z6n2nqhgA62j2dZr8iPFhJnnx69zyjBDkutQ2sxvwbZ5V
sVV2s4eIo2S4EFoZmKN3Agmfy6vCFmd5oqdx7xDzGI9/Grxhc20GV7RsMmi6
NtUlTs2t8zijdWsLZZfTskkL61Wm5uUNt8+ExSZTTJzo6GwbyMFKQ3sdh8sT
Yo0nNcpmPuwdJUnOf9/NFU6Mlg8agTFhtzmaSDYm86lEYMKaCDk+5OqwjHfy
uKQBzesvWAMVY7/y/nNiSOrOOXauj7M0AK2ldAtx5zYJpDnreuh5KmDreHYG
bGySjlaYDQzokIrEngPJ1c4NphC8qivhGN0eKb7Qr4VLXk/TjEiox9IXJC5K
o8QslvXQpbEp1r1G84Dgb0mCPbd95LFmTZXPocpswtVdfy2i+omzgNuO1jXw
iDEkMR4+x5g0+RiR6Mw3rMAQBsV+My1WZUZUxXdms+81tNUNdvUoQso47PFd
oZ1qiMdicJNubWwJYFy5py9/Yh3BfYFpQ1TEhsgol9eJGf4XjQ7+Sb6ntFst
Ohrl+/vIR+nE0qs0qTkSv7BZF9M8CoA8Ine9RfjoLF5gd2nbEO7TB+zZcjN6
bRLUsSaz1yBSDQD4O66ZgmY9JahR4IMAsHqLddhMfMUSXsxEghoxXb33dbmx
8rPjW06uFX9n7VvrJG7nPoZsLfOvGFZgl5fDDKwhfHhvUK8V8vNUhsSGIBOG
/pcf4sYtwFGPDcpafo+dJL+PFL+kjcRpBxjsQpW6nNLSHYac6P8t6ai46bIz
lF3U7lIyjHfg2hTQH96eK9qZ8FlYVLu3+tghUQFiLMeA7a8FJ4c+4IoVMosO
DPFizPK875cHIsFyC/BAPgv8i1qVlDb2yEQlg+r5ttnpnII3vlT731P8QnBn
Ld47WEz29TpuAoWAepJhFQNbOvLM1k097bYi1w9zO83jtw5ca7U2qYG/Zzxw
FwUoK6er9GUMo3WZLZaMM5pXsSZFHzhQljD3qRGO6GJk+X7+99JCv6BYcNdM
PBDHt0dB+Qe0vjVpC1QBD7yUJoWE0nN8/nkhXuybc8HnDyuPpU7gF5oFm/HA
+GRCewLyAdzjy89DLdUoEAxpBEPCmdNHR3uLE6Qoh0S73etonDJJWE375+Ge
V58mjGRsH5vOUJP+K7/GFhUx2f5i1oJFbPU68c8QYs/d4tAToWU4X2DUa6J1
8wwT7SByMlR/b5swTxAB3B9+T6MpL+zwk7lNIiBfvWN/j05IOtbBfV1cMKtW
9quSsNezqdohNWPMM+juXPEsxfVwY8zzDsjyjfJyFbgrviATOKrtTUidtcXR
SBvioXmBXz8qnUa1UuRY7l7LQnk+UINfYFePnDsK1r+zZII6BrrxYKMcBasx
W2gIruuEz9daqNNGvQzikg7VnHJF5HkCzKrFYxk8Q3CnAC+uwnXo36K0srxu
9OFUbmmv51gbu4EuOQPOl8xkZArq+jpOaI8pbLGEVXAYiUD7gWXM/YlPBHE5
I3aK23KeSluVX89d2U0xbrhVwMnP74VWy2gWDspkvVZE3LbBYsmJMg6yC0L+
o7ktv/PVbfecNEnw1tR2kjomAWfPi0voRLJ3MMFtCfI1QcveMsEtSOyAc4m3
HV9Svjad2WUmeQo5bppUrwx5Uex7D8vyyTttdJ5zyQcANr5qpuqNCav0+N/9
uhj7voFh4cdarK300s5iGOrXcH0rlJ03HjUxFoafHh7/3J0CLseJCLiM+A9n
qPVaoNqagRKtE9k0xpm51/uoH0klBB1jN1mHz+gq6ulxsGi9GhHRHa0sXm0k
r2yNvAvBZtTqoMEV5gczgBVtA41vsQygcl3d3UZasPl2hGlFRRoI1Rx8coIF
6gvZVP09YAP8FSE77ewA0T488uVQs0ko1oGIx9LI4U0hRmO6cdrkFhxdpTrG
G4YrGUmDddy2KYoQIsn6kDSd1P1nP6tvjSbT6f7VbhBbEn/f/xxVn1ESPxWu
UYXKTADJq/dmxXxQ0z65+qUhhHMYQtjhMGla+54/vzilA6birHITSnLCAtD3
6s580kbr7P8epfgd7AslrSEQnZVh6X5/t9Wzdkt1gN+wB57BIgjKtiidhPN5
tRu3PhLwecD6fdUjQ5Pwk/nnCkfjNfaooiqumZQV5RdKvF54brxB3+GNJ9NE
F88mXNQ4DYSbQiBMM+Qb3BwjMt/STQqTFix2XL0nidF+WuOrGf70lz9K0/nn
f+g4dUl1zd2R3VR2diVmDmFkysadHxYlh6azaKbZIxhpxLNjrEvnTMwhbUOE
dFNryco9KmuWu8GCCi9e/3jgR34ia9JFy0mCMJEWgHpLVnZLiY9dDVIzH9Hl
mhTUIiOJJ6E6qNtS35nOXWFRo9QGUwKxIOifo0OWgGzhFSvR3NWHVQPQZwzU
sgp02fLMMkBp+y9FdNKr8ASlZM3zohnsWmUOcE2FJiM4SDo0DujdooK4q9n+
QyKheY9CjNd5II6c/NOsgvC0gV4dBz0l9lFJ/RJ2jsqPJ0RRDzkf0XiB3xt8
35qoUa8TttylgbsRkzG164cOxRVjy2mzOwcL2wykWrW3e6gzh6qfuWghQ9lm
kyojOkUo/GcasS248NFeC2xp41RD49gAisF5YbpE8XXXe9NKdEeiUM1A2vsx
ift3twWlmZPjESblQ4ESRgmwUf7DhSWgzmhh9Ij3rKA9+7hwhFG3L6+i2k7W
cFnT0z8NB67qkJ+uDApJUjVHsECeJycNO54DTo6s9MqdacElwm3F0nPtSulc
STZgIfEZaaysv2JO8b6NxMGV0/FiFO48nstuzDdfhWSTZoee6bZJCEVDW1/V
7GC1DfSjNt1A5/PLzRsZCTeTUXyN4R/8r71qC0Srt1dPJhIoqJZ6G91NJ4cQ
h6osqo373O2e5YjlxY2JJK+tMyLtwgbHd+R7fYkHuxNuqVsjTMewBZfK7P/z
WNxj2jUl8+eEbxZjtgL2gNFAexoCg7eMyHu9w2b7cGZjnhGq2sfLce7sq1ab
RcBp6DdbmUzR58937p9WzVF1zDr+g4g3Yah/2S+hE5Q1ubxBlXPDzxxWlf2Z
K+LTfSKVBJD+D9IFLTqmyIkKlSzqo/nOc0JsdPLM9Ng6/lUaBLrBbHvc6qLP
KiY92JVMdcMGgfL2SgtsPEmkUqml/5NJ0tQXxQei7I98FWQQBy515oqQ8lxx
SJTQ3ccmhnhKEW2817xICAdrbAoU8+H/uvBmyFDZ6PNY0xDa2T0gRmvH3HeD
P5WPEdeV8+wMKDdKQfIvY6Q20+g3HoW2ct87GQcg2/1FCxbDvcMxuGb9bOzy
b6WVGQre9+P6W1AyWGppTly/dVm/hFa+tqrgXOuQc60O2tKXZmoTEootcmHN
6ORfz8EfFrX/IbJtRFAMJqgeVvrzGhpQCYGYqJQUxYwSEUSFYT9vQuYni0dc
iTrBzb1pBXYJL+wdyPeR9tqheIG0c0SSztvlOKun2wHH0d1/qgO2ENroDEff
pODXc7lU2ZRrmM4AFc+pwEm34ZIWfdsd0DkRHb6iI+gKKaqiYzWrgwB9juxF
goiAIk+tgFaP+d7ygjVJOAWRgO6AtdwWY/JqZNXK2XxlWaitX2YBqW3w0dVe
qGyd+TfEnZnYkiemslPtu1abHfi3gm6PHMG6VoND9i6LjVmlPcllqTdXP3J4
2tdh9PDBnw5CO4dGmuD+6hG2oq3by1EWlUNbfKWuAxnJILKeKeLQHk/liGjk
0qePhJ53YW8iwgLiB1Tm1yI5Z0A3Vz2uO/++efKfwJ0ge00YbG8bQALkt1lM
0W2WLOPVAva17kizY1yUVrqqDs0af26NkjEoySJz23wAFzFX9+16pTYrTp75
6KYRuTVO8oI30r2ww9okvrASms5GClTan8k/R/Qa8xSb0hpUhyl0zj5lHWUj
wnfbmWJRsJ1q+wUGre7UPziem4/7bcJgZxBc3FhxrhNIurrYDYIRsr7zGjid
yh9VhhWF9Hf1C5IUnt/Gifde4wNfG+wxpNhsTBffR6SIB0KIoX3+IAbdCkd9
8eJPd1J2Al3An9pQGO+lprwq5VYlYBZbogOz3FJqh91RDozug7mtEsnuxJl0
WZu0aqEk4BngpespMXQRnKjEi3iOWyNGTBGYCZhZwB40jKf/+N2iwCrwinc8
ZfeieKUnxSOmqYgKPi28yQsCfhZS43zQdcG0Z1E7rWKkH30/zfRngIfdH7Jg
+WdA1+ZXF1ZeLXMNHcVa98bsGZf+fZn7CZ2kCxy32dZ9I07Pp+OitSaCNWQI
aGMqM2Ap+SpezVsm0iwuiUTnjSFN0ucGCikBY9abUJCfZwocoGUwwZr5LA57
5vVlBF164kIDEhNA1ov8G5d/1TiFvSU03w5boQ7FNHMuhvZFPY4o7/oN/gqC
AdHLodjlOc9QNS5B4ro+RIOm7ZiLglTUZb7wYPDfFyWtIXPyQTEIBhpf7GRG
9zqzxp58V2ZKf4TRI5ITRKeO20X3HJwEGwRMC8MQB2TkMoImdZpBX/02TDzU
RL7RoCKIY60ShusWSFJOHUPkr1Zge4QziF3IcK49AYboMccG/57u4rjs58uq
JmCo1rpG0+qjB8LeBucWEXskBMdRd/o1lgux3vyRO47WWBHsOAaXVVTU1lfR
vo5WTK0FUZWJDT8ppB6MjRB+rD22l/8/dEBtH4zmhqXJUGZVcDszChjiAHGw
CWXTAJFJzT1/vxoFy5Mm+LaFWb3TaNkQIykY4aZpezDR3OeXcAvqKGFX8A9W
XrplPaSIkfH0TA+N27y0ly3FNNITgUon5eU48CiWCJFn6MFBf7clqbhjKdW9
lMFAQpAwHB197J4j1dgOCsijFMYsxlKteR9szgzi931XOyblC62552KZV7//
mXlGpuIRwwn3qV1iM84WOuomSmyLyf6zWoi1fadzxVFTowowMws4N2tqOZba
N3Mrv2gJtfJXxs+8WPRsDHA2LDsIEfzP0Xla27Q2XfCcpizCaVCzY5p+h4Ic
OQuXy4/7riOVp33KJdvhQJtdG95VZpv1oryz30jy6ynJM7rPrWWHUW0QB9mG
c7SE3LNjMx1ClZHE7ZPDITmsgncoaNKZDdFhDCjSqdGPqT6yJV/XwHdsLXgP
vNL2N/sC1PU3DVAitWnYFIiqKkHWZkImlw7/6th/wkhdLmZMGLB3e+cqCwNW
JZpNA9rR0LLsaJWCflG+Q/jBflMyOTh6mhnGZYc/+CbN+UgoVCexyqHisJUO
dhZojMwV15WQCgEXdltDXRJ5Yo1TCfN5E3nhkSo2QqExSsIXsUh+/nk9Sqd7
6iFnHUtRnAT/3/yI/qI9ZS0AIMkfqKS1UsXGssL5zwqI9lezijs+UglEQjmH
wYxDpWQrJCTsRkoN53lNXvOqn6bkuH8Q3twEcaGzZ0zir/3RQKVWwI2oRp2p
VDi0J8rCFE0dO091AF/aaBTfsn3JIl31PvQvgrz9W7cYklUj/n+hbtS+TTtc
OILHWlPS+y42uko4uh5cApjS9jlYA7tpiWSUjN7SOZmpIZ1awqle/dWhIwUr
T4KvqOjWhrHSjW+YzDUjaiZouubdwVVLF/7E21UC+ShryP69/HCppW3uQ7MU
IbsvJMCNz3MGIKF8Dk3g302fVDiYl9Hrrq+iXMtATNZ+efGVPUkvTgRxwcHL
/5SNPoGNUsxxMHvjPYz51KJIxCkA4jBuvnDlespNJ2DmgdFjfdolXPNx/2Ty
X3F6p2UU56HHGf/m9HeHD5uvWPGeG54WHktVqzjJzNDQtsbLAZQH7Bn/gwKw
cT2ROPIMT36me966O0uLYCqXFDQEVLx//IyPo8Nfch4ORUs6hEeS7oKhCmOP
9TS7vt4A2e690YdREdpyu6b36RN+UO7STpP/wiAYM2WI/rSUheoPpIrn0ZWp
8MFLsmQsq/dc4+bigQ0I9Rv/p+63KSMczD4zxaXhhSx6q/Ljo0L3Kzg07m9N
/RJtAGfwoaW9CxCN4WMFDgm1u2DgqzKDS7WehyG9DSit7sQk30ZVE4/Bnxwi
V/GOYH6TBCquEp2Q6PZAAe3ZvInsQpuGRWXckN9N30teelOoSzuAup7Xjs7b
01FK1GH5gK8hYylBqLR+efMa9GxJ5FV7Kwmq9V7nubywwXqhVlzXQHlxEA+d
AaU6gRp72VsSIYo9EkNZK/R/eeDBZsLxChKhhEK9+mDo6X20pc9PWF/caxXk
MiUj7WZvqFDFHG5rl2RMNhm+1DTwRhWsIo6ItwE9e2HQ1pKARsT82zjtSEVA
1CupVeJZhiNPOIXyYVO3kJw1geA/Oqb9XjiWt45iFbfnJntU3nqLdIPpyGgN
xo0al5NJ6FML6Z2An18O4qbPUm9SQEZKdmaVzmTFRWgM73rrNjkwYjesDszl
Xt9/sO1Dk+oCqdk1jP2rzcUuvnIJ9FYAIRdMXhfRNxfYYx0Brqeyg2MHIJhl
3v+yUr6JNPTTDZcvQIsvxpcN/AZ0hzrONdAJ/zMFURMDDHL6cnzg/ox+orqj
Fwb/RMOjQNNHNiKFEEsyuN6/yqqPk1lgFmWAmBwJtzkGbjiPpQQPmmwQ/gg1
x3i5h4uismRejm5k/djF6amNG7LMKZB4mvJEd8YwFTfr6KbmXlOboS1gFDE2
PQNdLBTeparr4BIBOIDNmgxVjUYcUd0d/iiXZfbbwYfKnn1juD7YadBXd+CL
U50cHYyzAkoXGkSDL2IXkK88ibNmjphK6Q/z8t2jiiNkpGQqW01dTmjspgOA
fhB+Vrgc8CTGaJOyDKf3oyR2gelwU++C5RuHmhEY1EeyDpI9cJISML7hqLBG
HlC8EWPtFkJidCAfpSZgX8wK5FZLkRCc6xEkDwP80pP1X0IkN+S4t7m27e7b
Yq/K7iDvqRvyIVNTL7sl8lXfC0jPx3UkZZzcMLoFMTtIMu7R7vmE62MxH6Fe
nQY8Y5iR47Zzo1B05LZhEDmWoAwwKZTipyyoEXJqhryz3ZdZqB/70t+EhvoO
i1CNLWbZYE7t78P022pKpLzzO1l5Sc53y81on5HdRn0CrudTJ+3u58jeMKnf
u1Xp+urBRtsKMKmgPEnCM+A4mSoOKCPezgTWyBmbBW3J+XzCQ7xAQzE3CxAk
4ZJmfeKHa5SxsyKd8tvMaJNkv3PVe2gkfhSt+HCveqKwbmMw/+XDqP/o9N5f
gA+2OGXKJXHnReJNsrV1hKUW9VvFFR6OASSW4n7yDXnEVKSuIVBXbulsSZDw
AseO78m6hMdZ35FteyAG3Wwqi7+IHUHZn/KHaIUkKVGJKOBj+2tenfOvxNke
46Mh2k1dm8mJxyQKTWm6qCptQaGex/3GJj2W+RVWJ6s6IGIU0s6WZYJbZurf
jBrE1xqu0p10gQiJj72h7M8+6cTm6iyW+gqIjVZhgn7B52TXQd34xz3M4Kpb
OmqPrWVQpUi/PFACMSBLLPbsaU2AX+K6ysRtiqQZ27vpkuX4TVzD04Y+jNQR
hDt7HMC1FFihP/qYvG/sb4Cxb17gcfrP0BAXL3tDEcw0lHsq+IhFuCDo9U3X
7IqOkpqqvJfKcpI7oD5Yx+gQZ9yv32YyYEfwFT0GmP2vmCx+w0tlB6g74i64
7scZXE0JLpTDWvi2BE3+vCGz0OjQmTh4QqnPAzKKYSm4gDy6kxgoezbd3PtQ
XZfgNW/SfuNpU4BCEIke6Qq+AOtfIVNj6naoEKWi8Y12zYONUIeyaJ67Nq7b
ZIqaUJ4lvqfImkikdMkaaKg3Dz916qb6oaxzfq4luUp6L9XlhcDaTvZZerRw
WiF81DbPuTv53RVaTKSUjYsHqPkXy/xPQLAye40tJBaDTfbmOCECJGcHND/5
9IDF67UdCDkkhiRunsxc4LAwBlT9YJojM/SJo9KaGTQrG4Ew431axRBjqH+M
3RTxDU9c498Df4Si8uxhvYNQ0gYl6pg7MQ7CcbHK7hwHiZK0Mk6+W6dffhIA
83fgUCY+4Q7s9peWzXBTX2LFCkoLSFYFALYLODfhY8b9fDSk1lQ4fd9zpKQj
G9W3Yxe4DBqPqloiCNfsALR7lxnPGryanSAd8kbsXqip+K0mK2n3VSXQErGJ
088JE0319FI0OEKq0DAaLTqOAMnDubooTykdaFeb8og4yxvzdCMeqOQaHHiI
elRp78fzBYC7I8W0c90hO2rIthZ7EWx5TnxLHr2I9rn/uPr1WLkyayi0tPan
1cNHP2e931NZ5rGilhVzdcr89UP/yDVO7szGy5czMQ7WPazC5AqO2f0uiGBs
211WTYjuy/tAZ3hZIqm0YU6YjInIdvDn2fWx/85xsoLKXAM3Tf+6qp9GfNLy
ivMkOD8tX9tZW+i3UA9RZHfOPHSf9finGDdNmtjHx2/8ZGTeaISP02a9L6Kw
aPZ5+Ll/i77irryBX5von+DYQo3syDdEC+mvtyP5TJdNzFbWSQ5e2d/h3cOK
5THBCJdbsKEMwgXkz7tCfF29gK20l3qagYt0GJUmMeRw6rACSvbnzw82m1fk
DDN9xidNBy2ylbk5z2SW9HONzzXJdc3LuD3Sw7hJep3iiunYWNnIFY3opCPb
UxRFM9bHRPNQrtzrBA1bL7LSU+9HdiPhV3J7knwxA8wQqa5KL5o2X59FiIyM
S4Lx5Q+zf5KhDiuaGYFn0oBgv5N1N3ie7vJP6qA9c9wdYaZwpshsg7Pk9ouE
jWsT7wuc/noLNv7GR+Etp/d7n+6oGw6zB8/iSytI2tpur5P2q+CK9tdBSqr8
Xn5MCeo3CNDZKXBklMYcKK/NrGHulpRp958bBfHcQyVgqeUKybAoHT2OrX9B
EWP2pnPztbaVmwVo3/K8+SCzvudEwQjJzx5IYaaxC8aW6lBHnLGvQBfkklkr
so3lW4VasWD6aoJJdgcvdHU0yaS3B74LvovOVSHmJ9YSg8h0QIpHk4rOobe+
Tpgw/b1KnNvr6Ew2U62NxtZ0/BfOnLq+UFR6/c89XncZoPCjXFCXAoidm3Kc
CZBILhKEbNGy0RiZ5Rxfu25u4EmKPQi8pyc1Xo2L2wJRvo5X1rlqT3zwwd1v
NSW0TBuhkoclGoOQduQABrKslGh8vbi2qZTOAxr7m1/Tn9SUxh05AIlIkU2v
Q9eZwXr3C+wIA4GkP6rfv1qwsjQYspJabVB2DJq+J6UYxm44vDksfTd/LS7C
VkvhcjnGoxFmc++pLBF9geoCummElJWCooKrAF7+dJne0Yq/FQxfZTFbRxOi
pYqS/1agDIdNVDwLoG0Rla1YCADz6aAeRkZ6i40CXdwDmRzwh02wGKlnnyD/
jHp14TCi2IMI9v6DUfoNUyZqzeF+IUwKGQwDLVnez0HUQOypKcH372IFsXXv
61Xqf0u1wC1dG5Bz9y22HNUDd/65gsldHaLwOf6CG6m2E+QsRk6lJquNKoxo
LG0uxgmCIurn70q4QDlVWH0O6jXL8Lrns8OP2shNdiA9H1NTUaaWQIvtryPP
QgnwQr9U5/ksjjx8Sop8cAgRy4ZwYQytMkRPMIFgCEN73Gi63LdIj4FHk1n1
VlOOhXcWk0BqFL4NxVddBnPLo7OsMSHLgXUMFjAP6XuSvsqLoNRS84e3atNY
Fir2wfMti0aw/EtdMngE6nKOHA7xL1Mev6V5YfkcEqsz1hw/oH9b7f91DyHf
tTGZyF4ZGZf45xXuDISSuUYc+D7HdrcK3FvvVkVcvWi3GP4TcJ/0+fa/HZt/
glL/FjLdk+x9MuaBogXAePufx68OjW0HrRToFCzdA8uSnuRlv9RrUrVIS70o
S4fKhwkA/Ez2aF3GEYRxh6zuGz2Rwm7qPDHFD8de+ojAAB/9N/7IuOYaDOeO
RhqsqsInb/bXoTabB1Mcl78mCK2cm5Dlo67BFRbpiUVrkpdtdL03fYZwm6pC
Zvd+4cRXzqdGraMu9H/Zfm/pZV1zFo0p8WW8w+Xq8Mc5i8J8ZgCY5CRp0OGH
aZ21rHOUdxpxuXjAWCoWv4LU/2JLPuKgOl8SXvrJ81EcC8O7033WFQMOwQPJ
KGBsvxiVSK+KYte/Tp5Bcgl/dC6uR9vrwwI7tuntwobWVkrHlFTdBdE2hIVR
/YHh8IoMxri6G+3hXiYSzWAiVgCIt0EISDeEGTrW9wmXl5M6gp8lStTz/huF
bGnHQAQVFSrSZrxGbXjvFb+ICaulAqD7Gu+wAu6+h5ZeTHfdgaIY+AsdzhpW
DIg6xO12zaOPtGIFyB2L+hzmR5ccpantpR+q0LmojpTboVBRHxCU6j7li7UK
VMd2wRqU6eSbDbHONXeHPlsQNvK+bdSFmvaM7GQkpYcLyCGSe7ezsP4HYITH
Sp4dWxPMNJQlcKDRp8Yb98bhG+MTtcWnNn+DhaWCnQBGSEsakxcPKEXmox61
n+S7s93FcewlTJ/bgwG9Iak5RMVDnMzVtktD2fRUAXb9EyCSqFkpwbHgGJid
g5B6yrHDhKQNMph+IJhwN2Uvxcls6kKjvpdD34LArO/Iez2ttPDJGUSlYly0
X6oPV5BsFt48Re0tNvQnOWHo/lXV5h1sKjh3FBcSOYKBdBVl4ijLSQgk7/QQ
g9HWufXipos0viSVi+Dspm05Gd4lGQFR+M7csZhGkYq2f8JNRDH3ydPWrgqZ
LXHd40VCAtFQWScJrGnSUYwnn/XOBz+JyG4F0CRxiUjxF5/HwSlU/9cOaBjQ
RCe//sqKmiQlrUssO+VcAn9KaU92JD/IfJVYbqrFhKJQDHnsulphDycQpRGd
nzbVR4NQXDOrrnXs+rHQl/eIHmU0iwPaQVs+5ThGha7EuqjmVhlwkjQS69/D
/4FBh9tdeQuPUCLQLBj6rYWbBYmiR4CvUJTZv408bJm5of9LKodcO72leyxa
4AzzO31mltVG8nucxJkQFy0TWxcnGsbiYBfk2Dzf8ReCtQza2kcwKhbTnf+r
jW7C3jizP2JLLep9iS8GGLYsw9bQN90jmhNkSwaro8l9uFJRkdQFZ1GUaIe5
/7kM3CoRHIhIQDz7JoqPZSb2E+bHlEs7eqKW2g1PLF6+D2Bpg/xsYYCKdJUe
i1QfGBaFpCZZW/oW2jYXaV+G8yZV3xPWw9jUBSWydvrkK8YSqNd+2qOlPRI4
daFMQoJsPiIFnZcV1oABm5dCnc++dYSJdMCrOseh9jAxVznXD0RozRB200PY
Vv3Ypdd9HFuiYe7ThzS/PKEnRIMFVjxjdDDqrhZFjr46u2eq3voekrKcgVEQ
3ZBlLngJCCMeYZ7fBG6pzstFT2bEZUlF/LxE9phsvA/KuSY5LoMhY8Y4Psnj
KGtCe/6BFAKfaujcbK7UiGVRc4E6g05xioYELiYNsqrurNZ/DCLAriNXhsR6
lTH0JBvksQ39n/EkF/qTsvWgDfVLfijT/l7UM93RKw2NrRh/RZ96bIQPm2Gm
97OvI76n0JcrsWCSH7ZGWCv6mvH6mA7EN4jShYHBtJjuI3TIGoJtI8NMzFnv
rJhHvwNNs4gnXR609vxLVF41699X4x+AsSjMqY9JKeE+aUQy4IUbIJOWdcIu
lW81ciMV7yQBhVBhk8N6ovSbrrRw0pXjqwI272hsphcNuuD+Qxh+6HHzAA5r
ly/arPCFjqx1Rn7MjyVHpQC6Wb3WCkXcm9KTNf3OxvQ7bdmFsanMih38iKxw
7l/cXQCYtHvI79Zbsuj7nFMRioLHBEkMIqV5D8ykupHMRhw59/h4V2V68PmY
xVYuMZE82y1gDHiZQ269RCGn1PJ4abYJjvNkuH+ceB3jWvmwAFsC1CzBpYr2
axrUEH6lAluV/bP0O4ol/O+mjhM3rCegl4IipKHDR9CWRvUnvmeoXVfxx4RC
m9byFf7nQtLpUlpuHFIfaMSLuIDH8HJX4tIlOeX9GkIegS9oDP5vC8Zl4QCG
g+eb5yAItf/3djpUxF5m+MhWpPcDOrIs+H38anbcI9RIGYEZnUYTpME9gGJw
cpxZz+wh4+MIZFI0XKZMgcO/ryuby/SDU7uP2yp1oGyE3EVwx7zbni3AM1xA
eLE2RYMupLJGGHnXOoHatYkI8xJyal7tlX6vUVEgvHIbZo/k2wgB5Zb93ASp
DWjWqFT38BH+u8jdHesMY3LS923Wwl729arkFaWLb6gpJ9XFkvx5llK1d0v2
nQ2H8GjFHLzKbnDn/250Zwk5+NdFjCaofScsCeB1Iqyu1HRAk923PT+/Jy/U
m1wdKSZfuveRDKoPzhYb8gl/N6PI2vw02o3RZdJGW/u5ef61O6U0YKNMkJfP
k0Nuq8LQ1CcQIEimdDYLuufu1kQLhLlJPeGGSaiJu/yi7rHt7MYYZy/FPAau
XwvKJqq8GM8L9JvD49thNPaa2OcwnluLQQY8b/gbuwbEaz7sxweeFLCUggee
jKWwAjqEqj0v2MO+7Dpofrg8istNDFDdYce2DJpmcHpJIoY/K7GgdmX0aTdM
hc5HSoyTO0+sMxFCp+y23TK+iQCqjzK+lhcjlb6cbPk2GK8OzrhaNI5KApKo
3M3Y9em8BQjaPwmbsBdjF9yqra2E+K8Hqll4AVPMCHriCtQ89VhZEiXMDkC8
Mbpqn+SCn6Tu2jPe/FQIsYZOoO55Fq1G+VzZEu25OgVaQioj3ScK4gFg+SBv
A/RWZ/Vt7GSFfiR4jFWxWwb9X7LEOg0o4NIWezA74PMFNer6FqcYyzockmbH
CdrGmrurJg2XqdlYSKXKfa9+yMuSvkupJJn3HyRJqyD9UX9LUagiDKLYB+Rx
xx/5nJglTz8Cw0aCbiSixpHPxjOveYYeFbN7Qy1KzgSC1jpvBkATJhhUVEZs
R0e+PiDQjx2cG9O1ho6KFwUHEv41r1UGiGOEbvyKGZuPz8mosTmhg6as3Z+5
TaUGet0QLRkqpBQdlFYajWZBYseaRbgoA/0mmbPQ4AglPFMV+yer1VLvD1N7
dlQU83mauLfkbXeSKV6etad00OIASzO9klgrXleG+Z2AeJgj080RW5D9/JNK
+ruIFu5KNBnMODpLKFMq4h329UXblw9bSc2SMfWAp+9/tIagkif8NK/aOdlG
+R5JkYRGmrlg7DIvb5c3sMfsHIjG2gNxVJRjiJbO3hfNtOb4Rma5EDIvjG25
H/68WgT90weP4wJGKIAOR/uUR0KLpEUI1m3LfEGqAqGypoPmr7319ktPeNec
SntgAZSDLIrqUuRB1oXI1tcna/hjNNWpxBTDfWSLSsrsVOWCNTwpPGP5ImvL
0JQWYogjdSoR4nZMNOjnokyB2ji57OC7AzJFel64EM0+yBeAxJE1qH+i+bKw
RritaEq3PItwh4Ob6y2lPPgMYPipklOo2znzAhxd4qXk1DtKlCQ9ZnwNYjTX
xBYC4blxSN7nCurMNReeL63R8uksr/SVEHDYg9gs/Eg1AMt5TXX5IcQ8QpVH
uYeZX4V0ux6rsGTmwttx5UTKexm60BBCXAt6evVWMAoeEwk0BFDC2aeHKogU
OXzzJbG3EBwk2f+VTF95WEnKMXP451rfy/sn/lbIJlWTPWTSssv8U4qFXVfN
CefdsqnXHzan2cs//c7dF10CttkrjZGZ0FTAWGrJlKWoXwyK1Ij+chhkcKmg
6ytGHzdqpfqvsDL5qeWISCtd2YYnN9tRIxZ1IcrCR9d9MfpicbysdO/3FkTN
01ROHQvD4PFrR1+Q9arVch54HxD+mJEnFXIqSqtrV2fMwiuC3YKE9enDGJFY
SgszpDOEu4MTu+OU987ix0L2AgKB0+WLHc+sIkaYRs+FgpgZ7dT4LKuPUqku
SfujDOHFOFuQN68iVFhtvztHGSwMaPDeE2WovonasKsFLU6eija/d7dOeMGY
pJL5+HA1F2wH6V89Si1Cqm6sbxtiKizwwa9OQtAES9OBGE1m+GjKwL3TvB3/
A4V2exsQXawSBj4f5Xw71eykLCfqiU43185ZsEBKRHpYcIoJBimrtu7/KAmp
eIN0Z2q/Soo97wl9QLuqXo3KLPHjomrjuDCTu8GZytjeVjF8Nifoj3t42GM8
nFoBe0unIAZw9HlkF/v7orXnnvkIHod3jjxUrKs8QBjTEZFpoOJtzMIQkkin
Xfe3sYEMd6WdNAmF2o7EWW/V8idNgjS/KSxDrO3IV7DWtFsIT2KigqHvg9I5
sWlt2Dsw/S6PAZSkWqBLW96H9c1EVuIk09UYNSgdUDR6FDnTvPmx/UZJLToC
iH98NtSbDCuVkDt2+m3WtVipxQe6YMdKH4us1xqtqm2WZziIU64bCehwomH+
6KGSRM+a7jelsOjTXyizyXHm6Ro1i62hCygiDlIC6EyL6w0Lj6rqyLXF4BXr
luL2SLxrAxGR3iBAN7TYHWSQ5TGJf50yODQHIsvJ4z/p3sfdp+FJgxQqOAdz
D081XIwUnIxx+Rr6TpmFtuVen1QqmMGg8SW3uSa917gHUkXaKHsfPyLZeD8T
kOsrrtpiUeh6zWWz10Xb1ffDGYRSgU9JyG0LqCtO5QKUth8TP4qrv0Hw9m/0
4lriEGqieBaAePluDjrFLutRN94va1eLNfl1IflDsFsG8YXUEyLnuLGaZtTR
VzKJfpJlt1b71RR4PAfWOmRS19gtyc9rb8HpBJwbYWQmZp6/Pc6rYR1fRvai
tbDov+m2E7ZFo/tRxA+CyHbOcMV+NlGWx+/jnStSLdU4+8OXECHCOLUn0j71
uktLjO8KZmGA7xdCZNVsRQfRi6NlZhnx6Pn+g/rvyO2uVEJf3XX+3Nl0L2on
OozrxOqhc897ZzX3GsQ3JrfAUO+qeG5cki1zXCnY4p6TAW+sUuxgOAyqOZvT
YVdMhoOgCw5FbtgOpVIAwfGBg31hfc3Sn2ycOj9xVkGVL9ZXsrRkZA+tPYBU
AmlQRih6v0kwWtVTMWy25O5Pc/f1CcSoixa4y268H2dnmYgU0YBEYAtFV97l
SgTx+NpT+bP9X7IVICw5YiSKwetRdEo9htB2u0fv2nA/h1XC023O8wVOzpnJ
qi1JuFexcB5DNzaqJHDI6JQP8TyvZ6ex12eWm/QNYpcuMRMlkKBxZLO8Rsek
W9LGcEQ7YMK+7oVX0Zr7lYZq6C2e+xmwJRCmXngRHIUN/bO8g930RC2cybvd
xip5Yfu1Zo0uS49lyUvYRmm2TydeAAqE1W/Lblsh9hSjZeRONIKBX9pZoSzk
ZnAAKs6pzHrAyCe0OMtGeZw5fOr4ZCbF8y1L0/e4LZixGzpwZ/eX1F+GrOoL
v1b/hZnNf+Ls/dgDobU4e6W2PbOu8sC/juu0XKlxw56hsX2eb3bFLfpiIgYk
8YECMJJgaoWFWgzET44c8hc9WHJ6Cjm2hyRAcpxd58WO3OekdP0M0eT9Qvz4
FmMZuN5lqte57iGV4KTsYsp0x7B1lug48nVYebBF6Lkvl9n9SjeVM8c29j9A
xSbDpVwKA1RRmS8J08gXAXBk9w9lZqGF4+lbipDFdTrRvL89b/NtE8/0w7Jc
MC6PVLogfvsh6NPWtTaHxrFOlHZIb7PVW71TM1ovziVBO1QUaSVz+gGL9fqK
4f5SPef7BngPEiBQEcWmxhnI58VF+KmqVnV2NFW9rQPo9Seg8l59eo0s8bXZ
EekHFgzJaCrsjhSbC1pRjAU5DJtY4qh1dsG/qlw6IOLIIlW6KXiawSJ8lTvf
iN/iVVk22mZU0tewVf8HVSUsHqZ2vvPmHag5fgb6Ql+9mYWf0pXm35ysyjJ9
Q+qQ+bQ10BvskdmUCgoQ61LJI+GDDt4DYX7rrZRdNElgh1puYEN3FIZt1Hpg
6vKH2W9p3Cc8ayOaEL28mSvupXrzvMGRNUnaihxnIkgndaaxnIH7j0ZlGhip
WRw45NYf1sDCt13tb2ZSUfgyrFbL0pHe1BKC6w1MU6yYGmyV0UxyAWkGO0ZR
X3nzjbDmzgaHoJViOIFPaUTRTGNRYeL6gB2I/HM3Z1DQytwUGykNzjB1Oo8j
tQrfn8ngDkJy2DkraWmTCoHwHrMbJW+8aWxZa6GFhhq01FWyo+SRzewshV5z
1ZVNgrABPjSfLxJqTXImIhUoE6GdFaFgr/VsMbESCy5ZCRo7WYLEF7CsekjH
VzRMy2r7GvW/mvM4uQJzXPc7eesCjBMZz4lx8OKtGsuChIpVaOVmwbB9qxjr
DvHbwjjzdQkprrWdC3LRZ6UIaJI8mk3/l/AanhBLfM6SzucxN9zdHPanZRiz
9q6xVC8Mwo4fY4M1q3NXFfRUJMHSAUgKVezrctVC2mAwYlg41SFMMSf92/lq
gKAxeEAYv760kqkt4lHZCLZD9UbFv78nn5GZg4Y4ItR9nMzT93Cw4oszediS
/mIb0ZQeik/VdLKKVkUmzDtjBEXjzjpskFkWk8VL0+FheVAtjmFzmCDs4UdD
TS6wrHuLWvSLjG0mYTfUKawerU+iSlzbgDKex42fnpDK+w19cm3l1KlELiX0
UopMSeOeRYwS2gKIW+OsEyH2FZbYqktGyq2bUt8UNNEYFfr9p9CpRtIBxMF8
4zAbJLUSVKWbLLrzTMEOv/ILsxQh4G/IiV8/BBAXYAomuIAWLMnU8oeosF/w
YiMR+Q9Owsioh60BjhOA6PtrjMbnKQov7Ax4YfKrfxGKPWUMUFeSYNQI69pH
u14fZkVMd/idneNDPc3aRGgbp0SSsR8jR4XqV6EYAg+iCehwRlgzge+TlIh7
MkPWSqn8K/zN0c1SjE/xzrpe3Gfnt5A3SbgiKneXi4jh9WOTkHreDMX/ffVo
6ddT+VGNWxJFtjNs8sYjSS+yU+88lxGICq2vOuskBg7Ph50pYQFIbhrZlsY3
GuM2YHcq2Lp/pTFyH2sKVKSINN7F28h/dWmrf1qOQQnqdbmyIz5nufqh5fr1
3R5jGJe6dWLKrfnupbZOd7C7O/dnJXwDZ3HvbK0D+5cBJy2wwWJ9+Rnc1jV3
yLFx7h8PgRwD3kZKi5HS+/x5z98BbSp8yDpNoVe2R3ak9yfR3TPsedfyfpIu
WUFQzkgPpVvtMSwan+YqOxjAWLfW18JBOabUc0/N7nCck9sPbWlaRK0hUcEQ
KXSsxMj7sTw6ZrmFTl6saiEwzuf/mR/Qg/HS++CiGzSHbhSo5TZHq5Yn/9Ly
EzqDKBvRN00E5qQhzlM0XSYrbDwPTYIq2cpEWIqAqkXQ/BaQLbghbYOa4GvF
VTWlsaqx0acD9h+TsXhXXtYUUyPzVavyi/d3OAClSn2vhFGAAFCwinnhBYuU
PwKA8LdzCeqso6wGYUSRxy/G0J6LVWawovN3JnQ5/PD3F4qsyX1yXvoI8ZZA
Q1gT46gus1R87t8xuM9cvr4+pd3qwD7V+WkOllJl15Nr58hCZHrxSMPbogaU
sKtQYuv+mtQa1vFt7HfCqKBGDz3ckoZkByLHKhZFggx1Nywn15EO/vV72MX6
LzuIawDSSnT5CpD8hNHLPnWrpUDm2ZQZpMWbvcSjQxfgMQIClkWp+1ZFE+bc
lOFQwTbHYDirAULmpToVq/DzG664kHuRxInYt4qYlJNUiFR3s+yq0OyDMZUz
acXhPvcQoJJJfwgrktcrseHFGtuv+/Ma2xAmYeiTbDGhUFgUNOmtoRWCz2Pc
5WKqzDAZN+Cw9baOKxMTTNXnEdn9n5XyqIZdpp2NutnZBneHEnE00AECqGjv
w+12jBQvBLrASR3UFkC6/D2Gn0H6O2wrCyiKAv5QvKlmqD0ZlmULZUZS33yf
sPk1klAYtJNLg0ZMoR1I6uo4aLAFz4YSJvHyjy7OnbUibsZ3MKSAfIWY+yKg
cGnKG8YaMjRru+Qn05TnvmSewauzDPugxrgmUcxXdzaOEHIjekka0KJIMMqG
9073XGNmVdrCnTlylLd69z/jEQrs21/HKOv7FZUqY8M3b6CcQAl6fUfhr5zF
qtlbk0q6z/xy70+dx/ZnTtj4TchiWlCzRUUfv7dMST6XDRK+TgEBrXE+g1KY
9MSkL7UkHc6Yv8eGAkO7x8yPI/QGr78m86hajfEHTWaGSz2z7jMwEhbbr0PS
5KhUYZ5jyfp8M0cjLYRaAHYdwJbJZUQhm6+DzihzgK/dXSWTPFDRMtzwx7+U
W/XAFAknBs5zTSYtt2Etb+8nPCGygQAwuMmQaSyV0GgisoM6ZKekTEz5e418
VZnRSmbuoh5oz7Z0aefL4rPaRrhpi7Mp+piBWpXBC415X39dZrMFXCCoTQgi
pjeJvOJVOxIxXcf9lS7rAX8eeo5Ooc1vECxBsUy27PphbFCniVZyJteOODNo
Cn/TG8O3APpaWBHqUpbnaDhDGerFjAtTtC8nGQRCLwrHdfKMuw3JgXlOrRUU
kWj27P/qNKu2xpKuOFkIH823bjoNPkiQoJfcEeQhkfTtldSscByB+5umDej+
/GlYlaErEpEQhxVTSxd+2vLNl1eONhppjyLcRMfpsyKbE07d1aHLukK8JTmA
QWLSyIj2wrsDTnv99Eg+seghE1kOr9ny/gqV7cf9nuWy2F1fU39OpusLZ1RB
HC58uYJDVQyVaFhUtzIjVwELackDe6xnBY4GcB2FJEYaJ+tK48hLO6LaotNK
cUYQWahUg/IiO8Hun/JXLqTVbSyGR39IqhvGKRgdJJTj9uLZ6cTpj73jbsGX
DcVSSMGWqPK2/feDdgymBLyctXtxJjoXnTn4XXOMhlbY93lIMmr/WevJYHSu
h4kgGRLC86yOfymjVuKS4DOpxyF5aMYpPunRwQyPCGZZi46DM6uI254n7gyZ
SIGLRMJmDx/RcL4O3m05JSGbdYCOGsOCDWDh4qSKvp+4CbGfh8/1YUQL14J9
jBjoa9strdtwTIZthNMu1qmupIDLaLZNPnmVKS3dlheH9E3/sw2GiS7FKJU3
wVMaeS5RQJqQKZAUyoAsZmOzKKEl5sq2nO0cLLCfXMqBcp1ANw2hZpmFxBNS
uYozmOHXVpvWauwL2OSI0I46S/KojzedQFk4jtL+7LPh7kRQccT3JAPbw5Jv
UlQXk5iBEJcFG/yg4GBCx8A4OeyNQRjOcbO9GBDxhRd+8/8dVwdU/QCkw9Fj
l5gO5SeVM72FWDGyZNwql1n99XB/oS4NNajyeu+Ik83cKtmkRJZQvkwsWHak
odOtMdXw0Ch83eJnUTTXPGyuWcHFm5ru2k4yY/Dye/HxXh0yVlcs0lUQebFv
3WNqpOOXOMj98zWUbpzd6GRS9c68hWxu2MKjfRNoDDtMslYa+C3avf3D6yTy
dluL9iAgMFRKJJ739m2bhaQelRdHESOWqWFWr7pIq788Y+x3tXTzzHdl5PZf
4YGzbA6a53//zJJakBOjnYNr86WAUJTzJRXsRo8MVBkkIs3ECvmLHG8oI5/q
/AVkNdq29a51W3S8E7MT6KOuvfpQEkiohcPVXlAVa9bppiuP7OGJXPp+5TTt
PLX3P86I/1Af7PycRAOPYsOwnbZwfZXfYFO1d4eEVbfQbityvI73qOPtW0L6
YHpg+bhAHuNLJuG39PbYH2PzdEOu+F7u847U0TzB/EINgQsTcGL4azgni8j0
wXt4G+M0b6jlhbO6Mx5WBSLdzY4xPlJzHvb4J52/YrVqAzszl0qhFuKXx1fA
uf6i0YT+Wjry+lG/lfLk+GU3Qt/qJFlCkZld+txXFz4howiF7ZSt4nmKt5/c
v5pxM+5ZUKGYwiSlkWclrNs6l6YDGhABpuUxxm9Re+/Mb2FKNs4QcWuWURb4
fDcIvTV2mH09yj6wyF1tw6JPhp46rA29LGW/U1avYmgyfVuYA/neu385ULHL
I5A2+SsEqszmr9Cs0hNy2kcm7mWJsWa7UZLbZp1pQVQERhQJOCsxsqwRQosN
ISwrWN6gBduLgwOO5KbTtNTFoWNHoAD0/BMPxD5Hz2iMZ8hfzqAvepEaWOqk
Tno1O5ZFceZcXuKdxwLFvpUYaHhxbD927SWf1/WXMiHBcoxzaJCB6OXrgJR4
hdLPBhTkIk7hEzxr+NM6EG3+fkbSv7KTadnow3vEKLDRNjxaqqDCSLbQhsme
tMmH0ufg41lHUXpqe04gVFk2moXzuhijBvJ7r2ixsgONR0glaE7AN/7qaiwp
RvXeGAMxSERnMrKbF3Xn3rw4ieiIgWgunaACWFJ+cF6JVa4pAzG1eoiPQkh/
pZAHATZlS3utcoIz+ZVajyiynPb0oELRNqVgeQHlUyR4OuDqn1IpaSuCBifu
S9ailHCoodld/vlk7o2T03I+4qBItCaymWYQOhu7h179wYXpfYPANZPDYb3w
tbXOSbparsXzKnaZb/9G4gT1y0KrsHCIChbcZGyvP9xELSNJQS32ix+LfgeY
/ybw6tL2RCfGVipc+GJNJWhpWmbSMMZt5lerLM9h9Pzn0enH3HvMP5yZWPmr
scT3FirLoNLgr5GuRYPY85RNnSoZZVZ14N0CxUjA0eT/TqFG/LQIlJ5IPGU/
P70wr1L9Dz+TszltT9PWiA4UTxO2E2Y5QqS3nrDho9/OsTU94gZCL5wHYfM4
pjJvpOcC9ISDlJjkhtzh1hxoiT9X6cxVscwj0yZStnCCzIDfymFvY10JnzJ+
yJih1OvyDtBKkkc/zJQDULlIH+0S3/TYnoYjXTvoRks/2hrbLzLQEFuXBbNF
mN6muoEQSkQHYmesfgBdzQU7GTet1yjsjGhuCBAHRDgnEpfVInwNmMUHjndu
rlDMTXu/Bi28xpXbQ2GDOdB07ecX/klPsk4cvjMOOoP1miePJ0RvybipjOT0
pc4w7lqYBYwudXAEglf/8Erjr3JzdgvThhH5SrVPPbPQ0nOA6JmkG/OCiFY/
qHI8PUR+Rc/3OJGF8/yPVVQp1u4ifckv15K4aKlOeqtNI15EwdD/saB1I4EJ
U69ipjMQIWd/rjfcEe62pZdB0lG9i4WuoVlQB9NgZCCIHpxZFHb7fy3ivvhI
9Chq2Omwafx+hQLiaZusGiqGt7tiFWH4unG5u5M+LjSHuiGX9blAzV84dsKo
81lqHlQulmht5vq9rvSa/wRfEIIps3kqUk3AWdGve/18BP7TZS1lErPERi8q
Abt/mm2uapZk2Xw6r2SAEGOtYTnkUrCztqAJmwxCwOl+Y7ibiIO7j0ncaIM6
Pv24EdO9jHTTyqzQfrvvkZR2tAz4YMMfMeDHyicf2WVy19QROZOiZO4iWcHX
uMNzGsulceuv0bTM3J4KSbbdlU5RG4yzSF1HEmFUtd85RsOdFQyPzkdVXwcU
SHEQM6PHMKRmqAapdwEg0yOTpTEoPvAn/MVBg3Q4oUvWATAhOO2Lr0J2GwdT
3lvHrmoF/Q+CdOpRMsGll238mP9t5urDGTGHo0B7R6rc+h9ckn9F0JTw3Yvc
bH9yjTtJajhLPhaUrpXWFusXc3cRTCi7fh2geRMLMsZaVj5d6ZvhbH1M9nE2
eQpPVN7PiUE+ZH04GOgYxnd9D7MtPQEEX4GaB1ll88sdXJkycJBBgSIDWSx+
I67GrgLPVFID8m6IJE5YPO0xfcV2wUcr4iOajcr5X0QK6x6W1BsNokF6d/aI
XTZ1wf/R7ymhNSKVuEWxPFVJSidxKVkEjGHCb7JmOMjiMV3OXcf6wj9dlOkO
y0dPoC/1Rr2wyh8pVCKqp9y2PkVxoA0R0sYcKPUmkZe5XnU3oMSEtfW2Ofl2
h2Cz7J4acloWyjAYBavzEzuyuiZFH8RHU1oW+IUGsPWae+C2bnU+RB+nqoD/
t5SHRF6iE3vA37227uwDngSpB755VEwVuBz0lzj0TecZPzmrk+QasRv8j5e0
3MPfgI75SjGQy2RCBFXXt7ghlFQTWEJYNQJIYW+VfE1/Vsbs+kes5yVCPvhe
W1uB8wmhgDJNQH8TNb5Vb9BpNln/vE23GDWrhi5LUYh+RXn9PVR2/h/JGGZD
oBMHAxZVz6gv+zByRo1Vh3/dIEs2uXy/rvSq/crmMgWxY7fEhKj9LBIojS/H
7O9uEswZLVvKc39bF9xo7CiYKAocsaGDvT5J/fGrMIU97SJNrBQJ4y5xJlEa
Vn/huh/RAZJruLtkatha0eh/LeREdTOHU1ASXsHNO8a/jaxUriQZSBui1tCr
VD15hx8NG8u2HFfxGVlgfQCt9ZBM39xB5F/QG1F8eHl0s/Kfbe9Ed2kIDYMq
V8eJ+sLj0CWCrtFuyLcZ/7ZaEUuT2lgrI6EPv9LvgXL4hUC15GXZmV7+1UWU
IFNOw2Cc5enxcFx94l2jSVNUCS6Uy9bY8Pc0kEYXiP3T2vz8jWjY0uL3/sJL
Gste3L34oGuiVBd9E7zhgQlb0MOdGdx6OsKBrC5OOjA8JevAnToSYW5/tuHv
CoiSO6Pavr3m8dmA7ILzUPAav5jc8yLcJ+wSUB+NAhzXOAHYD3C6EDGR4//T
+riUDDRXOVFMDoXSOSYCEnQ0BRVvFDvO7Rq+pxoUZSWYwWBhhninDAPSpbMI
AuMedPG2eit98bMkalhY3tUBWyCtA2vPr/2i/inJZGPVx/CVsk49CXksJDgD
/RbslisvlAe/143owdelCQOigmXJCGAR9bz4JQoyRImXzUeq20rYFkNm2Q+I
tdWqwL0g8eOYwxrD9cOsaFE1UAQkGaRddBVo8a/0yoS1BXqa2baC3O7k3Z5y
BNFC8MRIIGOjaei9kouGgrtGIp6ZnjCI8NaJMNZYvTovD44ar0GjJOqE/h9t
H1xC3ffLh0raFjdeN565h36UQBg2txQmIu8yDsuzbG4GKUc6z26WNsNbfmBo
41o4u0t3uHjEu1+3XHk1DzgF94nRYUN298C8v2Wy62f+fuX5Rnpi4755jQXL
huSD6ILWQv+tXe0IGdS5aF7C5YPFUkxEWDv/U2ukzwGgyUaC9eBwrfN4Gafu
YDl+x5x1zo5XqIWm0UXVBwzsXTElTKi02Bo8hZ9jOuS+JmHgXJFSLnDdNMBx
MhZs78+gAz3JnPUAqKAHsQUvnMSRfekRjw/EYUAVgb8qC6YmWlXvW5H6LL5A
yDAmoP90Ztps4eyYuIMxt1LEHTQpfkJtCbscfdgrYsKcHRM3M2bJeIfd8XeM
HLmGzsw932zNyCX+w4c57qez0ULltU0zEN8nkq8t+JRT4dTRkTGtTO6xFvv2
vV766fZQ6gN/i2tzdDcVsMD9+N9FkCliWD8d/w7dJSw5mZskzonY7RZKeSEe
kqSmW46fAQKC7Z28NR4d2Oqv6mo3XjVyX+JedtZrM6tSQRO9sMH9a6nOQDgu
7oZHDtP6gFhaOw1NQYtDLIxAEvMXA2mYqOL0U3dHOp2aE63FaiN2Lbm7gM/7
aefIsYft2ENnm26PtxppKuyLZl0TtzbdDwa6baxBgvhTOUHpRk/3H3nU8ZhN
S4AGxTngPFYfk4dX+s5hzP8+yD0+bY8wJilWh9a/42GABXR7SL7AUkmduV+v
ej08q8+/NOnS8bohVH3Y9Hi2tqyLAVROQLPvjFS166UjuXyz8dUm6esQWqQg
lNKuKl5MTkyzdE8XmcVJiYdpBDyAUJqsR/vUmxj9YAZGiLYR+ppnn/yDQlYr
VgDL5lUpwlxsmBgjHJOaL1cQk2foRKePcEGVWHp2/qyvF8IJvZ2IHSoy4AOj
kvZEGCijr0OUDA0MbXgctJWscXJx2y1tqT9JsWKf2LM5oQVJAjF1bifrHPnJ
wZyC0aXRolG0xB/YF9N2+noCPj1b9vCmddebz1nNMLQkyyiD9Y3yzjmh+Mzw
OEBmbNZLF5HZUm3NfGmItKDsAbGSMbvcw3SMIgSjN8KjF/W/+hQV4QTFqEmW
I2+hlJzUfs9yIXvgfDK3R9gG2triTI5dNr2VC4R2yCxSg+cg+hinyNS7dfkQ
8xjlSS6psBD8NdqEIb0jC2p+Xzs2vApGjun1s2xCD6yCmWCHkA2Mvc6tO8jf
nBUCDJSB786Sd3bJlOFDrGoiC+0sumRAHgbut/k9MayUQcXOWGv0Pq7xfaK5
ZJ7ywUmhwWFJdYMOpTMtM5Py2WHgjgeis6yfVd+UgQQ+bM/pz4X/H8HPncZa
kV3Dwj9or1RJDegkXhalYWxBhWtI+j0BtFWoIVL308X8MEbwaqt1iQFjKd00
VU/cjLgUlKtLl+kaHtIQsRy5JrkADkd3S/6f88QGlKA1s//qKSO0K64fSA04
fGMYJ9ySC3ZbKQQW/RZti+h3wGeTMSwvat64ayeY8fcVTVLxcK48Zm116P8M
66dSMnYjR4fTuIzECHMH9dShnNa2UtRNzJ0/4TFEiqTc9WY9SnN1uOt7IL62
GB9b9G78ziF4kxKUBs/yle8tOWACkic61VslRmPyC2uAfZdnvoKCG3ET5U4g
FD9Fyl/GrP0ZubZqIX/Ff79OAXmx6Jv2vXtFgPqVxI8ZaEtTJXOImE5EwlFG
lvScMvyC0bWjC4SXuyMKTJiOOMuBK2SpIZMwNQJi28g8R0gin/yCYHgbMRAy
cl4obncAujXsk3zrh/kSOlYI9Qc9xIcbq/Gj1o4BIK6rMxGqZ7yQyIwAygEA
oNmNx2rfsoKgJeAdYafBBG5AE/3IN9HTQ5Exs9WtpbdsCiaJLyc/NWPlrRw0
clW53ZpU401cSpxSruebkl/NHwkbxLDEI/VGQGN2vqPA7TDWsCzs6FppvEr7
V8zF6RrQ+jRvrYxqr3UP4Am0iBBt4lYwWKJVt7ZqTTIlsjfvrl32WWNxscHe
tWDbxxn3G9VyQhr6MZnLr47xAq4HoiyDzmmIxYkTfU1Q3fuBbsRgvdt0thRe
TgiamQws5iHafB8M6k1YkppjGqEBwJQ8u7qKAkuGNcTE64Dsq6uYqT0vSer+
54RGEXW1BOSujlyoS7i3MohoH0duXT1d1WvyU762wcBcCTQY4QKMipvI4iTF
A63CX6a3TmxlErzXi5ftL+tJpG/uNYbWW1Tzpt+q0vfO8dGOJ/y1z3q/TbEj
eXCmCbVVR8RmgXu6ar9N9kSkcLzXhbciKmgfV33MkpYFEkc3V7HxJfkBBgZJ
JqywocvipScGfsFhN8TOfeVcNZmFgGD0IN/H4AfbgGBYeRff5SnT7j66Rw9N
tIE6xXzYzQyszYQhSL8iOm+YcxD3JpS/jlCEvoT5I9YwBabPpXvin2ENARxI
2mWzXSbILPH+kwdWJFnXAU1z7Z6xMv2CRHN2M7djUU2yH8eplMBR9IgaxzIY
xnhpUeKWHPy9hboqab53K1Y7/mW4atUZyiiLNFo66pg6QamRWlT6u+Kv9GR+
g/FGWzUsDYh2qPDhZVVI09glUSYzWsuBKnX1dUC0411Xkome5X7rLPqt8s4b
KTcxOptxoqVf6yPV7GniqpUjUK6MxiCACujg8Dt/zHMiNBT8slna1HZz3rOz
iOuIDRq30a76l7yU0GOXrFR3i22uJD4DGhCqD0N5PBBgvb2OejFHDTIkymwK
lpDXSTjBzz0AGfNmHF5LHqJFxuC+PIM+XL89UafRQAEVuUkn77gB4YA5bV2M
nK0BiUGx9OmdOSd3ffqY2l9q0KaAsLb0cBVbu0T/bFarvo78CNl4fB10Uw33
8BmlUHrhwTeaFeS/ZKK3lD1lL/tmlhh7V57FSPQY4UCTZVl3OsViLLtvIukn
DyAi+7a+CzaXiCP0mjUK7ykK8g/7n+1uAeZ+XcrrDR4kVKPOC92MADVyQ1R0
tKA921RuqeY8fV/Fibzc7fVouFS7Ojll0FWzmFd5CPFjA9cxAZFs4xp3yRMl
W6TblcEn1TE+80xE8Mol0Tg11oRCwUHDQvOBaiGt1ZwH+9XUJPa6TN9ks/aZ
2a1rDORdoH6O3kQ+ADXaozHVLeYjXno/I/TyD3iAc5l90ZNo8p8YI++WeJcH
pV1TUhRFiOEhAC5C0Awl09KiJDg2tCfbprg5YO+idRECXaZXMQvbg2L7dZGz
+oWgBP3Ra2ip57byXXqYE0khBkNQgOH966EP3UWRp7q3d/snInK+Jxw2zFqp
z8LuBIOcnTFwuafPqPFHu0osF2yLUUmvYCJ37QoUWrKJjY4j1vT4iZH6O8bL
77BXQERPyVRDGrrBZnWC0v9qKQsny3k1VyD7YUSltwgThwaGnfatWBSyAmw7
1XqgXyNMX6ev311IkWLsvVlt/BuC2sE+r6nJ0Mj4Wy3G2zjg5c/9pe8+aXIS
YyzHwUDM9dFzJQAbyVjGCc01zTqd7rOVIWc4ImK6W1ZbIzx6nZ1Npl7wKpYH
jnBkDDN8V440tg9lTB5Cm/IYZR2GVQQh7vrXd1mtcsRuUUs6dJP9mR9fWQmj
o82vLyCeoVfyGxxAceFPycESQX0zWwv4Vb+7sXAvtUx3LbE2J6xurelecX13
+1xEid3CIjn9cGIXtvaosSy503bT/X/DPEXp900zy44u3QmUxs2NJNN0giks
cyakGWWzCEe6+n9AbmRxwSvTL+8VqLbAHvoSLtpAkMBHSGL7jkLwNkjRUafS
65LpEuQrFRe0suaGVZJqSd504PxFZ3ktfegaM9BSQdLFgI8j/M6cJUgm0sZO
TkGtgAOQlMO8M3478nJyiEUGIs1x6ikfNJ12jVwMGhnZvjKG9bU5lr7OvdBH
+GeHF+BVX5Xs53W28lbU5zx45NoNLexTrWx+SjJbEGptqmhC6wVvz0kGDShJ
pwFb6xZMWbvaHoJlRdJUmNZvmMIzHE2hhCIUG1DCOl3VIHYe1K2fPJnBF8oZ
H8rpd87ojMb+CaczFbGbWulQ62hAjcq7YBLzLRLFW72brcEK23mfpgAY8EnW
OUhYyDIKHAcBUBHs3sEbl8ZpJ0z6rHfvbM7JTxaE/qVDd0+iJn57WZJs/kZw
aFJz7PDIjfA6+eTvEpdqtQiSEdsU4ZswdNqRXXmpqPXrw3Ey77csGYD0B/n8
8VE5lt/wv138BUNGRYonv5GgKgvkQFCIrZQDD59moqrAtrppXP+Ma3U5Ut59
nlvFiQamCA2M+RRncyK/xv0kLAErzgQADcECoNopQsBJ5XVQElsA9+1NbDiD
7TW/qGxeEw585RDN0q5GaqdAtCsHQaWi55xH9lJWcy+XE+aZZMtzEb+eW4P6
sg8zkt3LS3vuR+p9ybtQTwELK+p7hIAPnphrX9TM3+Iy/CT2loeNTRR8NmLC
32CL21y9BAFFO88erIZkC+C78GiP7+nM2a990RYg1STOrSg88y5tfQA26h21
iFZ7/1n9cYNrsDa/iqMLKfJq65Ra9xS7ygFOEqJb6N2+gpHCWTKeOlunROID
DH9uRoaoxHcNEhs6dq7oOoGIeIwn3oh//xW9AN/noihunRKvryNUp1OSmT3r
cqYJRHM+iSSoo99cm9VNyv0tBiFuaNUeSapclifo4zYMoAV4Flp7u9jjqfQP
ZDcUwU+M+2WLIz62yqySUiQQL+fwHJ7bQhttZyxq1notomDcNpfwoRBJ9L2z
qrF4HdeFbVLQAiEcPZrJsxm8jtVfOeFOErvPLUUzZIuQgnEX6RTOywlmvSx/
cQraSCq2HrHHAKxvw9xZX+VP4cfA8crNL7xKocWZAGSy3qA2dFTSfPgRPOKU
v+DurNH1cCIC9DLLjsFnHaRQZ+qh4wHS5+FanA2H70FlsvSbVrJ0OreXOpMu
akYn2lRo4dbPQFL9HGbVk1mfq0MQqKnVs5ndlVSQK/c9ByUSAUDlQpFrYf0g
Lp/qI/YGeug8nPP8hYQAPUf3i2dyQ0KC9NPKak5/Q4+vif9VxS/OJ0E8waoU
KqTr79o27OZaW2yuW/t9fkQ9UoyWFXNbRXjftLvbSswPWkdcyCoYMfuIu8ez
3vTWGW3dJu/sA5sz6wC/qZCJS6v6eJYDsk2CSigaFVOaGFH96XlzaBihPhMY
u8mH4suzfN3Gz+6HOthruFijop+nswtvyT15UH7jq8FZL4qQz/o5LSmRmLRi
QwrLYOLqW4Gl9DaZcQ2wd6sq4qC9NLNy2Oz8kKmoAGyyzw2SORKhix368DBx
r0YiZ73DjD9/yC9Hzuedd+v2LDT9DZE6H8P8rVNiRjevTv5ryw4Vtvrv3tTt
Zu7Ryob3zC4mQfCLlhafRctoNYAjqXBgdzfx4kvf4d/Cebvt61OHXn44rFMh
yiO2V1AzISCSQiHBy05qNrtZ2afcg8COcLiAx4q5QZTcOtykSBFozHD2teiQ
7a6KnYO+1xpJi6Gr25X4uhyJMe5qiTMKVZWJcosxRhdjNJ9n3Fc7/1z75PFJ
oaIxtAJwgBhs+Z7fLTol4w6mjd0/Qa+M5ry2ecyCAvgjaV8mnM4BFtqsU31t
+3rC+85MZK0X1iqQXctUX1LK8o6P3wBrc/fOqVDIrmUaP2qBeoXATSqltBOQ
W66UfTU+pf1VYREEkrv16HObBfdCWJIumkX70GJ/cBtP7CfsNEEUw/tVi5EI
hRV5cfQH88Zip13oxf/kPmS8wZTL1jlHkdfxz6uuvyucRlIByqhmOUej5TSn
5Z8iaMUW9Nngagoj1eb4QxuUASezUiivIaQtvGivr7JsYug9PlJ9chqgtEpq
G5KcY0Vqf+URwlPr9gX2XB8SbwAqyvubNzucccGD/DddVLnf/zE9LT8h+K2g
ViYSaKaHexH2UhihP/6VsMPBFcfIBz/Do0+Nk+GPw1XSPPh5y+Qhm40iFt0X
aQzOOtb5U/idK45Biwbgahu4WzV5d5o3P9zXKLxoWJbmJkE0BoC1C/OtWjZ+
yX1pcwCcSPYll+iau/KdvNUFz6iYLWo72aiEyIhXAMYdwSLEQkb7ImN9PmZv
wqrJPYmzO00wJ8C5g4zxPhukIu3ldD8TWFoJQH5L9/+bz99pTtYH8ZUScsnN
Db04TdgYCfFxdKtduSHzJg75MYLDaSHwTS9rWzUupisnKR0fGQYFlxp/Q9sp
qJ270YvFrcLn5Nm9PfOrBQGA7w7ZjxdLGPsZw0q6ryGMw1agG1CAzpzQVYqX
8A+IYMxd2VrPKm6bG46wjc3iT9oFG4pkFvxLoCdmuKhMR6hzSDPJ8KSfjssP
zYjHP+VrMMHWpZfl6PxD3+nt88fwRzeVG5ZDqTynZ7jOXK254ByuALP8rBhz
/fhs5OcjJ4bLeplq+bE3RGKNQhYJgyqV00VdzxegPrSXc6AP81bPew041sdp
N3M1Hy/45CNwTh8t3WlxeMdNkELRAutfefiYW85OZ2zwtq3pGDBsx8VN1Ejd
8ydY7ZYmJqrmtNUCbCvAulQXauar3EAt6b/DJ12OJy+T0WIUzkYpHiFkmbOb
kgslQ/6YntNTM8SdeJxxxAQfGgJwYaPxJw549uhsDeQ8KJN6mLAPCwV5RPjD
heeCz2ynQDA+0jFyXyukewy+MYvcvWUJRnYlbGJ4jhO8vzZ1Gui5sbeFJu1G
X87r+zMI/MxAtg+Calag4I3H9qqHvhq3HjGE8M/dpiI2BYMbcgsksEIC8EZu
Vhpy1tPIgId5shqbqBdyJr08DOFLYQ3pLc2NkP2Aq8qK7eyTGiGKP9jrJbfr
5Tradlt6z7J6ToonlfEtmUGToaSyob3VX5iB/Ta7pPJVBIJD6icxpJFlHiwe
CVslNIGAUj3Bewu2Pz7Ixyfl6U5Fql3OwXZuvKI61LEWPKVUZnbjgphla6bt
kSxVpF79RZb1AuPbVtGUUDq/hHp6sLNIwulPafMQ+Qk2lQtqbbXua5IsL97X
fhaEmwPzSiFyyZ0smDh66sZiQuKTcJ2H5uF1vumIPkqqogcG5vbioF1C5JEr
d8NJpyDPCQZ5YwCpYUOEThhLZi4F43BIn5x2RyualRi1C3eXbGHJyFqvKZrv
nJPX7GBfA8klJzRxeGgfcClAbFNan8pGJT8j5oE5XX3MLPwO8HvbLeCSUjZ/
md4qdX2o4dI7k4FzeQWqUGhGGcUzgcPFVqYwa967e04OkOM7Jndwzdf/xNkN
Ibuy+cQSaf2wl7HH2o4hPDYXh8TgjXvZkcDMI9qVTJFzmsGw2+fgjSfmGlR/
hLXCx4FOr1HiloaEsSZm9tvCIWsEi8t+gPTK6dzKKY8CIP1lGm0OMHPtCuis
6w/qyP596gMDhuo0bJqozd2Y7vanCJnnqJJ5Z2kM053Pbx4DrhwtxD0MNdrM
er9FqhKPqalx+wEQrSeErM8kaHbVbRyOXThwQeRK3Q7WEIRG9U/c9LKDlHF0
kZ80CrNZebBTo8QQT+/LvwkbZ5vG8nVdPdABpzlikk3x1+VQ8j+ZeQLcaglI
hwenuZJT7iK659GD2B5Nm4R4VC8FG4nE+KLa4joqbRKOm5iruwZjx4BAXHQ3
9Vags3kMtXidz/2lw6lqkte3Y6eP6hzFGPrnWZmCNKZfD9VAyoSRuQIbbMek
+X2GfGj8A9rCcyfZsr6rABxCElZ2V7u2O8LGgeUERmZMXFKUxMhvcCZEE/zd
RvCrg/zt3IqWh9wNy68IJv8bmw5Tx04zkmicbf66rEnTcIgyN7M7k0HIpkRE
mdWHBQ5zGZJXyktVEkuHe4T8zf/x14twJbF94xytJu2v/REqTIjQgg2gWZGc
pZx5VPEQoPVtRFLj1iyguR8TCAXu72sEn++prrTGxVQzO1wrEDdW758cSJ/V
fXt714iGm6VxcQnl0G9cHGiNXb6wVy9BUWxPdSh2Mir1whuVqy5nPeq5ymZG
SMjkVAs7C4cAOmpa41hsXSuM1EdyxOpIsmsNVhRdzWaFOSXj0JWKqHBE0KVX
zWTbuZlCJZhUlGC8yDIW5nRQjxfiJwv7V2KDrns/xrSsRLPDwYRYe4Gn+LVT
gY+TDHH35Pz60mPicuhQay/DNueWiQsfA71BVpbQdr4CL4Vwmu/D7SdNnoXW
LjnREyNSqYxop3BqS3LeLcYCHCpiurA9oTSS4aQlTERrIE1LI+X5676+YGuB
YRi1oFheQYe1RQG3zzE1e3LfIB4jhgyAUEG8Qj72sdQsfBCm3/Vl+uH4Va8P
OlGHYCCyn68LZFN6v5kQMYYdXHcjLjlKMH8SsCheCxUKjyBxRLGk9bPEGtEj
bbr/Gu0svcA6XXd98FsA2JlTeQznPOOziLjIsMGgfRxAfsUdbOWsKJyeV0uS
lgRTU6o7RlFWHdmLx7yLV+QCXib7pX8B7+bt0xs9UDPtXLQlW4SQBAGow5Ex
TRQMgUD6yc4TdaCBZOWQPpNEqzMVmfsVw3k3cYDxG4reJSY4D0lzmD742zXg
r2AvXR6GLOXDsqMVZkDVjy4UYVUpTjf3yPIUP3Yj8SxvfGaPy5jYXYPywMn2
0Mmt3M4IMyUVsl7jX3s+iuCq3KLKxLx1rC43iv+Jco9U1MEp1zyg7kwT6OMk
GJQcfzz3jLqkh99bCSdK4AZGszS8QDII7GfEmvQK+rxnd3vQzT917/BlqnoN
wt6yDXsYyCzcAHYKFlu1zBfkOiamfT/ZhSbAYQsIoNSf4QFV8aKAw2Ecm/Wk
d5XoJQViEioo05VUUTufA763BtoD5oIZiBsa1Lrz+dm8Q/aaM8SMk/a5NVbF
pgWc0EBt9rI+DKyK+OQ4IwJLJWxvheHbU23Kr41+ZnF37jwUY9hpqt6uW/ha
w/CaR8G0DnEZUV1Py23DysNL3DI/w0qpypuQSUmbKNA4T/E4+w8SZZGbkocB
RaZGNcmIkYH5G7M4k91znub2SrLr2YiGB0+n90UfoeItEJqrIT1UW7Cv2rhx
qyPoEqa/zIG2CntROgNNKQHemE4ePbGsx1D26x+TQc1YWgQI1xh2pQzr5FS+
CeG2W3Zo0aA3kGNJAw3/33E5AuHX4PpWMe2I6VWxdMH33iJRkXaLHaHQHDYm
QVBhzt8NEhE0GQ0clZUQKA8hBFsQ8abx329a2y8epinE0SybC8aV9ZsvmBMF
F55ywMVCmGN6tXkGTiy48HBpxz8tmcHWoAV9fU1hLYDnw6J9eGkaeVA/HjHc
GaRkcJWFmzUJ7YT+OLYscVOYmKX2kWsl2lTu7BN6y/Pq7tDlWrFq7kAVUZhK
QExIJgKJaYIarmyv/40IMMlGoCiVwV1WFfXZ31rJiL/wwqeti/6sS4+zlO4h
lMpn0cYMCcxDgozbcc2I2nuM9j8XD7WUzyv/o1Ytg4z/BxEUX2A/g2lG/M2E
MV4V0y1NW7S6+1E/NggFxB4opRZdeD/bwq3zVjuK54s3utB80k0cj3/ZiZlM
GQs1cVwLGESkf4dt4+MQk5ZqBViZNLOJ0u7va+Re8ETUgvDxM/t5aSoB1CSU
RUwKTBUbQjdMudn2eZDN8FSg4UNISWw6JkWVUylKIDFlE3w76MZgjsMxIXtv
shd+uLKsn4IOFPiTQzhUlPml0Q5plP6FYQk9fB01LAlpghJ1MKelGN63Xnej
dad5gHFaD3Z7IZSdblBKeIMkSEGE7v8ASByecfCfjxhyt1eMp5oI8xAKHc5P
p7aLPkYDLoAe88GIvnjzHeQJVWqdcsSENf8aYi3Q9YZIJ/DAAtKwBfzTsUJq
UsOOrCmOs9lMj0QhxZSnXh0iJrQA7nIqRMj47zSYWjJC6Pc0oL17Nob4WTbb
yFcnZsRjUG/moBXRV2IZ7irwL158qVIdekAsb1CGy/9YBmPFD4OuzOTphXni
MttRA7nVNIvgA5FatSGl5K6bfBD/BO7FnnoROIBeUNRa2fNDjcvebeMTBVuT
sGaNTKfJ+k2BccEh5bDnGWJK/4Ht2+8YF1tWff9kcGrPL1SAjiRLV6YI45Rc
z9XW9GaZR4yFJjCXFbXNcZeiXflEcHqRVIwp+L8VZ4Gnei9UfV0Rm733q6nb
uBm/ecTUmRvbDPFDJiIyc0xXrUEb2KzLzvfN4Iy184QyluUuW1ivXjpoYOir
F1ptpZ75aq8/F4YfhmTOuaBin98ah8DVveZtUVNBu/wq9EXNfLroDaKwXGv2
+t4ORGDYKNfNZMxpMuwVpBckv/a8sMj7+UPW8aDQNXHcXgWc9zhd8aOfyds5
L65weqpJ8CQ6sGiwGM1zzvSh8NBfJagGvb0W/Q0XTcrkVC3I2rUZ8mipqj1j
LrbNV0debVk9AE1k2sCYTUNC3if3wD6Tch1H26EnLYAcfY9XLWNilJmkQUnR
dDadAP8C6Cr7Se7eDYMFeDs+LFeEgvczKoePDvB+gdEEakFjJACm3Q7MwtjT
etwBsyka5tHAdksHLDVokcX3RkqxsaN17PhKKtRrOHBYupUB+g7p1x1szsbt
a71igcZBY2vWVsNO6zHipywL4Dl21WNzujUtf1zZ6qUKzWodhx2Sb0VFtTB1
0i1PYtAyAj+uZjDXV49bvAsODts5imIxdn6yVRWiqltyG9brxox4Rfew/RD0
JywcvTF1djNQfznzNaLq5DGhol6U/PonsLNumEInYTSG/u+tBnUfoNCDuFni
bbmCGTf+AbnNtzl/+BTKhtJ3JRu0EZB87FMODvNc3Udab5QajpWvmojb9cU0
BpDx7jZNy05U0B4KpFmiskjtO0/PZ5o6ltuvPIiYGtycMRD5twkqBebsF12n
iyR+1FIjqxSb2kGwQRohtHcZWv1jPY5Ns8qFbqBa8h81X++2PThXzgf6PxVG
ZrKb67ZK983W9uCtjSCv5ar4FoOM2+aI5UG6MhmZv+brfJYwws/BDS6L/ni3
HNtHLZkt1Eq/YsRR2GwShmMEfjpg8iqO41UGvm0oB4iZ1L51CfS9nQfdHawT
88p/tBS+JWB/C7KhgQW9zcU+rzA8cEzcldyPvCHyheE8+XfgZIMaJsn8jZhc
8r+qdUkmwofTp8FVHMrYinIW/q6SgeDIO1UoKnveu0cQdg9ddoA0JRx4UUek
apIThaxu1hrQfaFLYIncraYBHOJryLoTQNyRgVmtI5TJZb/S4OzFbYjmG3un
7uHvJ7WuNw//AO3x6JOo75SRrwwygkMrq6hahX22xY+ovRtJYeecKYPWjGHp
9ElHgEYF96yq090a+jszRA0zKb98ra1rVBfm0GlR8zQIQibMKtt8OpGXVTTI
vyH8JIK/1VByrumjnv9+1J5bwmu+eYc+BR5p4TkLGnQ8MDm/cM5DbQGYJc2P
UJ0NKK6FGY4hTg5uqYIXlkSCdHmy+1r6uOLdeZR98fKG8A7v4cFWJoxx3CJu
+hZlEq3BE1MHI9zFlsP3Lm8IBTt/kpJtw4cZL/ezeacUQx81Fa6XpBRc0J2w
mHO3RaIM5P9zu8DF8LP96wjUPn1WwtYd/VbCwBugtY4Ee9R23kD/4ouNCJor
QOcQSPISJpPp/ubqlMXQ04YlQqyoeOEM8WlhDgsXKiNdD3AYbv3rr5c+/m8n
0C4vsxci8Lp2Q0wmGpjTxXL/UjGwekUWuQBP1gCLnQ9EVrmkCtOJD0Yivlle
0PNGkRv/ASPVQbVe3zZdf9b5ezXxyT1xEfCeJrSG/gIi9tVL1OpMsL3jXGxT
vuxTgnLoNyxq1Xkjm7jqw9XpLu1jROumBBO+bYW3q0LAuLL4NTbASkUipz+V
KM3wjXQVnfVfSuTMplG9eH9tq3KsVQvIFlD6KomuwvrEA26qzbx9MKr4BBsf
bndN7MjiWvLPqKyOPc/wwuo0HbrsASW6jJWcD7ws/SgPRINlTrebDGM2qL0h
tyrD+U+5zAkR8/Vtbo6UlkInN4hsT1AXtlJpU1XhOfqdqY1OL+YBM/sgs11y
7LqAj0qRZz9tU2E0oejE83FMPd+gbBa1Yot+heC2IrjXCEoaKI/C7ucaDjf6
HNJG1eBYExbuRGn7JYfhFlH/mUws2QJCC292QllytSCGDywLhot0BNdY0H3X
j7eCtC6zUV2xTpQbgoBHswbjm1RXSh0sPLSYvF7EFXjupalDt4JKU+5lfyJW
OI7EewVtiZ95Nyn1RWli2N8YcGK9P1RfmYl2DHBxWubzhQl6qnyKoY/jLjdk
/oKbihR09qWO+wjKunKA6AVn9KJto90TcCS2mZnHsis2MIW4p5ftKBRIavvO
3MsTNqrhLwqjKqFSWDhVphb05YVxzzz6Y9JKL0CG87e3nua2+C/GDRq4Ik2s
VHdYMiyYMAfgm9wqqogEZgBTIbqQ0DZKxYlklB07qvsQVE5x2WojK7dBgJym
AtXUx3+HDdbtcp9CkDZle5J38O/94srvEIl06hYqrmTDobDTogM2cZJ6XIWD
4FfHSV820ccKZ0loW/1D1b6JhKzZbl3lNIoAj7lAtD7wSnB07IiLDdWzrSiR
B8T/yCbC+jW7gM52MsUxKZv690vFr96S/Mff6P0w56yutqAeUMGDOlEwP0In
35/psO/Ir0ju8thnl9DtsSsFQs3NMMzuan6NJQKEs94pINV36IruN0Pzd2ud
cA/rl/E41h6pFyFIJEAdfQVQIKR66a4qjkGyV0zbQQgTLg6ewg6+Uj5htH+c
AnevE2GuPpgmV+2PpsNL6ac/cltrTo8CnOQXLofqOBtB/TEne//vOhF41P6F
0wyBug6JgIWMu9pWknFzloPe4ufOlBR9NYQQ0IF2MJXAlAL3bLE3uyT5lbPZ
wgtMQvseM4XVBd6lB+D8IYxOucmuTsJ+7X0FNgKQ58cIKEH2v3/qXvr4EWFI
ES5bq1TsxFXwkPUvdv1JiXYR8QVH9dvJENDrrU1PiezLcJADNVoSfmYXDx8t
sgh0gAS0QsO8zi3cdevJkrEIhT7KnilvUzvVup0PKlJF2DBI50G7u7Q009cZ
NlAkJqtwYNxMrfnel79uVUGLKepoa0pMeI4L7dox8vXdgfPQELFq3o5eAt4G
yWungJoW7nxuRxbeH1gYqVV/53CYxi8t+tK21xMarwAhvcYxCNRKnRGQ8ecd
jmYy1HdkUcK4B1l2/40Y8ilglyr+5KN+BiBHIfV28xJnLrWFCz1avsUd6uii
8CRo4NE7R/JHg4X4dOFtivujbonBKn4X7MLZ24oerCDxb9kZbaAY3lNRmDl+
etZGmRLFfzKbC41VAMl+v4HKBVHZqzCRO231fYXSSlUFFo7hBBvh8OgMFFwN
m/FL6VXu0EZm3GpVqvei1mamQ1zbK5tfsPPNOBHCQoCE9z0/NB7GZhJBL/XY
niUGA1Thw8j5Si9knZIHQ5HibFF1NQ7JzkoO1tGa+z0GbQsMIqRDE/CxGLVz
/pOi2IqiwsNmx/q5gde7nzXz6WRYEddRAQ2F98O7PGQw6s2Jk/9Tu+4Alw5d
hO994vlgkZZ2ci+KRWI3X/E6hKiqfGMoW8wjYHmagad/J95lvBTaS8eG8MfG
4BVgYlG0cYyz3G4hn1P5pEgyo62xecWBiavOHJIcuulytoBgsBDz3TM0ioAS
scw8Xn6NvFp7ACUy8SFVvmIt9vLk5MRWZ+sPTic+13LzLMoiYHb7kWUinWiE
szzLWh6mwL2cFJvoJuYYHygpj0ee4uQv4TayK2EFMGMaXwUXu/pOaVxiwZBR
NPp0cx+yCAlIg8hV9itIjhPlDennAf0qlTIC90j4Q6ioHfGSz7uQ5ZhJKnwF
tzkU0FFTvsLavU5Lq148YJvn37UOlofDsHnAFqMxeOf17Y6sIPLgTfEwC/y9
Wjy/Y8cfczJQq5CweV+34h7qKCd+RawBUwRClwTD++cnjS5IcO4fG6AIVq0B
fDfhuuHFMPJtLGfN9WjySmB9zsZDCVa9U+/qamMniHwiUG2IN5Pl65cTTs9W
pw/U6J4QVlc9amtQ+sYXz5H5efxEeBVCQSF5b5gqBFnP3pLg6ExVaoC40rx3
Z9Mev4ml4SGTrqTqE0e7MLLdd3Q3/yAlZTAE2ZCgn5p7+ZN9viIILYTAb89I
Kwujti9JIxVs6ZBiU9ONqDzS0YV84mSJQKJEalTnn1r7eoE64UYreZjoCCtU
5ZJpOV+h2vDbKvHNuNWbwqPyeu3Xf8r9l23aBSKowT+w4vHP/0iSm2i3rKO2
MCCHowdRSd/jUT99+v28t6vlIqwW6oVHZUCyWSDk3G/PoXipPC5COf2HJ5Tt
gZTrFvOdZk+7nv0dBPFjwP6OD2lJxSG2AGmq6fnhsMELJxr7hpATjNcK2Pc5
MmDFWMitkV4hfGexACBQ/7f8c3McZ+MAKgMmlL91aKP1F3h8jlQY9lQoal6K
tivHbXNfAVsHchy1uZjHKhQFVxbfWrcrFcWsTG7qfWLbuyd1yLwMaCUULAQZ
z1nJ6PW5WluBgKtLwZTgUSkvl4J8JBL+PSO02W/djXF641SIwyDTwoOOQ8Tt
p6+GxcVJfDZLRsUH7g7EQfYeUzyLqAnclAjrGXLMYANL9RE59wHgvmdzTkzl
8yFKj5kmy0dEdKu0yU7iboWcP2JYuDAjAReVRzTOYbTG43HmIabmiMqerTqG
JEvodURz/kMX73jS18+KqfM3WAqtRwdZxsep2tDobxVIjdvCq9y5bGCrynx4
JUV7qgQ63U9zPmIInozz0X4LKYoBqXozG0FWX1OaVsyvgjwOgJiVyIC0n53o
gIATzlv6MJIMLIud/Dr8gvaTukrR2Qy0D+muoEd2c+O0b3NVJ89mMFBXrUUQ
nX/GxI8fJFxeSWw7wt0+B4qrM/tAmQ3Zz34dROveaBceM3yfiu6CcCJtD8l+
ghZZ77cpD+YJkBcwq953HXhJVgdg7t2bmVcFhsA0+AqwyXgK0faBHjnIZbPA
uf+LPs4/ymzqw3wDi/CkndD6AfRRJyw6sbpV6jaJxk3dXBFFJlO/netKRGAC
llUT+SdHCQQnEFDUcfO+EoFlpqxz5W87z7/4JLuXjL9R7zcgisnqQtYwQV+a
F18HNKSTMJApk58WA/nfgVfZ8nqgxX+3YILUgGIT7Ud/fxrFg1ZxfA0M+/Ck
BXTw+711BRBtFJGg1v9ExawcueDNXih/L02TND+m/izAd0XHE49RU0jvh1jr
MNCTLw83jIj3oFrMXjozlZ9skTSTzysY0pWInTvPFOjRAr7fCqYUjyxxp+Wr
ouNiawMzB+U4ibCKACiZeRd35sUJrmlPndpMx2b3gjWe8iAntPfVT80IVt9f
BSLK/2UXNGZLNpa8ggGLVDMV8bmijKXP6cVQ6s3obo0vVMPAigvedBM6CiRI
IoOg8W1qbIeBRG4/6HLRWcha8KD2Rk5Cjit5MsP/mZuCZU+J8tTYcVUbRwIh
5bSpRC8RLVb3Za+Y/B/UXDXDPw6isxv1I39xjaZexSN8Beu2fQKQTK6jFt0+
jmtPGPYmvSxGWJxYYpGlEhlePAlB16gblFNg2FbZQP03Cn95QCF1LNh+7Y1S
b4I8e3E/eiAYrdr8pDgtCrgHreL7heCX/EtsrazTkv3uyZdwC0MS6uk19Jej
utCnMqn33pDbmfWFJ8px/j7f7zPGVZh1bkGvLmtQHigfWCLZHO15lVdra2Qs
Py8DZuZfmaGBjvgTC0MWeOCrqv2VUBqRy1+CziSnMaIQ9T+t/8lCR97770R8
famIm2UT1SWPUmBY/1V9iMBo1Q6vni6O5auV8LnFQEKGnv5l0ZyeyE0WF+9S
OF1OUltxzF0tNxXEjfLGenATfnMXmkBDhgpnFTrPq6WXzDGJQWA7+x00JTpt
mCdiFiSOmPhCpDrhppJxwntCYeuTVD+KoJQa+uts/2JA8dz0lWuTZ/DJCXrY
YHJP0dc1qDrKQ3reejM15LEgWII8AqoAvzfZqq50XSELYRnFi1tT5F7s65uI
wkecWPTuaYJCjIlKHCznpYW+9EfOZoIW6mBXfVzkkJTghcaVwaSImnl9BNsk
KO3FJwYw/zWg70ec2DcKCNUb9u1UjpE9BJc296atic3KZkmA+ldqVrRhi/5n
aEitJIrrT7UcK8XpR9blBV9stFWPc4uUdHcrthWFEl/6Z+v66VPJuRse1QRQ
MrQbGIzUlk1sQSs/nIgkHCgO3FxPBXjZYFDnfWGzjjbBdFfBJz/kCoPkj8Or
thlFYjIhpy6gRsOD7EGCTWHeyQSxxYiTKB/FC4JW3rnXsxVa141CWZMOUY7c
4ijKMamG96anO1k7Y3xG3+2EOBZF1cKqCj8PSTFMXjacAxBITstLUYlrY+IU
5cOsMDJfIn4oVbjC8v3ht5ovMZx1zy3TO9jPyMV5mU9UeDDJJTXq6+7oFvP7
cUUGmzWoaV5qaPANWUJeDavwKSKTTcUjugFomZGGEov4vaaDdNtuE7rHHbzk
CKXn4pz2LhaDasW3QjHOE7pua139eCRLGpP7PNJ5wN+zQItLPLrYV/TtuR+b
bARsKRLXvPRFx1Y1EGC2nSwnWo0Uo8m2kOMavrP2UbUfhGsF8fL/dHPSGlyO
OZFIZpuNC0WDcmE7ixw63jj0YG36rILeRy3S3HsKH3Zoc+9vDtH2e05R/45/
YKe9/Rl52t01+b20hEtdaU8NvxClOmop0GwXvXSiZvrJZJmdsnqti8tTTbh1
E6WTfo5zQWSL2pVbiuBvMk3dKTuP28AM8RDetUo5ynncGjb29jefONaup324
Lc+7kYlpooO8ZwfmLbeBN0Nd5ZevNbYmqEKoCIF9hPuajZ4LPXd/9Ydkto/k
8iuX8PLk+Og5sDread4pJGprotQ3qyMofUIiG9LJ+2yi8w9AuOX2W0PVw4VI
v0mzvAHHGKv53wS2uoXT9VdiWv19QgBAm8n5EgwyGCpjAXY03r475IZHOxnz
nrGFFle6DSFTUr7+WxroKC2ery1W0Bqzc9Xe6k3enRpkar4pyZzNHoQrRVnQ
HA8ZBqVvHSUrQub/DMGbh5m0BpHszzX/GfbsZ/mQOJrcmv4tiFnmkA3FhfKP
8QkpCyWsZHw3VfdfFpAvO2G4H9E0FTk3Qq+cDr4X4LbOBesZOdyEpqaMZOjg
NEElN4eDJvfo2rxgTK4sQHtvHpUoKHLxqoX1entf7Te0DJscV5UTDcrwxz8m
bgNs8ZRatpPPUYYgUYAn/Ak+EhOeN6VI1IxEAL86K2FrFMglI72mtmbbCHbQ
e2Vfy/7sX5DbU0FnDXDoxqHRNDP8jv2GvbhamOxBEZ7zFkxY9x4m0I8PgPEv
HkFGf9VexcpecbKlPUEAjbi1QqqSQ2BZdc6vIR59z8fPQXZzUnChv0eYZhEJ
CML6rcjx7xOdy/B2QHzZfuUoU+OaTokAKF0jnRu2KZDu44dOng6Jt4ron4BW
KTQkwLGIGpqcA/chbcVUW1h/BvPqoCPXzhgiKtKNdBd6SUsY6vk5+UmW4H3K
bt5BBGbE59i8Pv/A1cebCWzNVr/Xe9O+etxBk9Ing0ifZOT8U6rZzcABhKCY
S23OCZ9ApEl+kB7vM2mm54yDVQT4AkLbfJGTsoawrags/tE9pgNo6SKP7JEP
FGUe2zN41hpQUYlhWt+I0tc1BdRj4TGes0oGW8c89kwchoWTeyT/Yz/SVvlw
p8LEwz84aGBwUIoD7tLa5h/JLcpuJtc/hUCOLZlruUySdFFfiKV2GV0aOp9Z
GcoCRquBklTSGQ+q6hdzBB2HdMl2D98m4imKD0zcPLHYZ2YTH9sWEC3ObdXj
fWMcfx/ORaSf5mohzikJ3UNrUxcLAgbZyWHJdDQ4jYpLhTqO+W+mzYQZ3uyu
awsSlpQ3qZKp6hR/Eyek+ZNV3CIyjw/1KLAYXIvXp8/ZaoIyg/inTkIfrJf/
yTFu+tQe5xwOf2xg+UFFQUlglgdfePp9sJldg/ZVXpYUmCpeW2RpFqVWccmD
ru+g4wOoEiC+kRJ2nleR76/Sq8Tg4bFzX7oGMYdD/x+kSrBWbQokGsyMFDeI
493JbJqhiPR/zKIoMq2SlxVPHQhUOIDOZ3iYoThsye2qEL8XUQapZ33Y5+kN
4jsWVcQ/qZpQl1ln8cy1pos0H37wof7WZoNDcACZ/D/+4hul3TVtNHbZqT4j
UVdDJGa4iOcbAC3hm44gwYJW5IVrF5CUVeX9nW6he2EyndiER1OXZAkHl4wd
V5vof4XM06rHSIvAQFWi2B7+c/beDRiM17EZoe05oSUIod8hWwRblDzpU9P1
e99OmHMxOB+asypU0kaGWe3hflGgghorONfratYJNk/tzb6AWCzFzO0elhUM
DO8oQ6JxzHylUOPc5/21VOGxAEWa0tvtxFnVq/m6quDFmIeIVB/mYext+UUK
F74EuX5jLn8RVQiNOBEUUQ1cvC8azyS7v+RvCPP5rZ1QnrM/Rp3dAB+I+/ia
+9I/oFAuNkgojpAQU/W/XF42pixIGaPLWfL5/WqVAYOwJnAe6YljCTUwNJnv
UoN/cC/7Damou2/XMoov4zL4dUPjzXpE9Zzo2sOB4LcgdZ5IukPUJ6qb0l6e
SfSjItWBM4NXwMAKyT16kcq3CVZrbq7L5ozTQk765uBiAPwSuyXVkBf7jq9O
323An0Zuvc1stp6SQBjFkWTiOKF/ed4FwZUpVZEdcFgegL0wsvKiO6tlANBD
YWdd7FrJxnxpSeXUBBY6V7gNOG32xkn/ZWjzHK82mPYKGHRyzor/JiuKhJoW
v1XFu+T2QaJwG1h8WdeOeE+QYxJtNJi+QkdnqtvlegNLh434ItEKQiKVI7Ub
vhwujx57BEElB3wPQPi4U5y3Cqs/9XpacW/Qxvx/xH98vZE9wAdNHAms4HWZ
Yn4G5jN3oS1W67GustyvcWOeKdAmgrUnRyXGAnbXjhfWfb846DAAuPZOerD+
uNW81zaq+KdUkAZ+V7E4LRzIcqNMYNv2946wEBIuyIbUMfS+lRlYNoBv+02z
z3wxZTFzHqplMbAVSoMGbHFTq/xZY39dGEiv1l/SY2AHj3E2cslN2MtOiPiq
onn6w8JN1ccVeiYgMd3rdKn6xoYT25kDXhHvLC/XmJuHKVdAfmvndsjNP3OS
xspgx156eAraDnR8gvt/1bJhu3DTnIFs3bpyOmnD140ZNsFEJV7xDHIrT0CT
boNMJ7X3tSG0RB67HAUj1UpWJ+Ndbqi3+/n3pMabQ8P2EiZ19NBGcf9yS/6X
z/gNKhJ7FeIeqzWC5wGgtnEaFtS39LRtwEwbcNWyF4TvsZ9kDZOPCLh3jLDN
v4tKazWc3AWJV3ouUZY8wJorvXoB2FTC82iQ/ogSv4/MrEWlz0Zq8bE+o4d8
rjfKHyPiaLNWS+3dkw/tX8yRMlGct4afZZjQgp8n9CPHs7Wrl9rZBHZKES7N
m4uxw+wC6/5oRbW24r9Bw9eJCLxxRiPuCFWWNPXit6xWwZOhf0qaV8ilY9Le
JIQtxGze79FlW8peinukIFlGS/MKXiZfU8N2oyueilOSG42ek+CCh3XOBnTS
QgE8gW458EpoupkBGk+U5pKzG/gq/0ugaDHlxJabVY8vEvxSYA2qWiB7i6rs
+51yzOzOCzjP3jUaRQ5nuydGEoMDU3oNU9PZqA2/HjmQ+YtJOMqzkx27HxUb
wXVOQGtNXFrd5dMMbtodOr9rdu7yv/EnyB7oYhmY+vPjg33vlv8zcUDmAX01
Y/1eHZIxkCROmeFlFhxdzGSLgoj+SVCQ9tg4gvnepudWiPhF159iWV82pNUu
GTWUw76eJts/2IARpXlziTb79kNSsFen4QvrGQBZPxRm8es3Wwf9b4DdOM60
d0jfE0lIVQD0SCWjdyi7C4H3tDIoqLlyFY4ngV78NZHprjCKK1HQsmXtMwkb
VjbYnKm0W2EbBMQ2WHUvV5GqlKy0imcB6LP4NQwvzVQfXi9JY9HCh2Y89V+I
Ix/JzU6YZipK19xZJWCMltZSHixL9DSqVNboJ//EIfEymdp3/tqG3r23ffNa
USvqAYuXzVr+/BmGg759aRGIVQ5Lnk7Vb0e6eSw9FcFVl25CaKSgt3Fy9aas
H4V3c1t0uSc2uEE/IiStbZ7Q6ASrqL/R3zKAXtZBmIJavMRwsBzEw+wmPo84
fAeCaKqOCdIYvCWnhj2JUBXHeNem4YPMpkm/sQsfNfN8LUeVAbuqANczqfeo
EO0HtdnPWZwyHZerWS+nUy4WER+edkKuSgy5XuC6VKVW6aXtYSL2wBJ3ZM7/
jm6/kAQLWRqM/i90rwga0/zP/UDkt1//eVaY5M0vjSBeXPo4ek5MtkC34OE4
TAtnVqlMsKpHf6jqXdJg4sXZBpEtVIHl3L4W/6iUsqqb7nsgJ5nuow6/o8x3
y5R13W+iA7FYW4CqtdX4r2yVZT4Mbz2/UcpcJPJpGwXXzcCNGjHcEWW+eGCR
BajM7M3YI90zjXf3LU3wfXXMbfIWQGcMBwiLRbXf90TQFKxqkL/nbLy8jzFZ
s4tIMvtCASMX0POlpjD6gtHzIVWmavA+IzTiPbYNguJNlHbpNKYa4X14+/45
DVw1QOZJdpMXtLt9mGG0PNUAt7mHwXdYG1PJPA77Fjj6NXrFzj+a9q+Qmso4
lStYU8uI1gpyP2fIZb4NTacSYd/tybS8u4vhhiWShjD7J2x1JOO2H5yfU8uL
zbyhjCQ2XkA6HVWZT6SE878OC6uqaeV7HPhE0+G6MvXZUG3Cr+SYXJwHGdMl
LrkNTn3azkYZ98ynRj+XYVDo8Ddk7yFG4FO1wyRp4GY+VNdKWs47q9d9HyLt
l49tm5+Xtcj1Wr+Ziig+E379OM7mEM2evydaX98RQgegcKRT8M0WF60jA1Mj
z0+dSJY1TeXvfqiZ9SGtJudj0S3Ca9z+IQdLBzOFF+n1qo2mbQor7mBXHr35
GQRsxfLt67ceB/Z4/9OxnYQfckneMmW+d4zcXTVvlcotliA0PC08jrXERRjZ
Wunr4usSmhlvlkuekk2UfHuDNJG+Jd5NfZUFLWPOZpJNZTw5d6IU40R44wkY
KbPGHzWaXXFu2S7YmO7AJlIXu1XosL4JMXOKF0Ho+61FzhkXn3qV0dFwFPmp
1+Q5eXSazbBzNxVOE/4l29tKJLS5OMLSDdsSwH0xWYRvs5xljURky8R96J96
RTxW43gYfdsFmTcz4G/ZyIO1KRGuT1unf+z5PsKRqlfLJM9agFeLNDY7FDMw
iIKo9qZ5vpxOMy7lzDtjeTgrhcW8uxwnF5L2x5KWG1HPvt1zqGwRLkcbkbCi
PweduenYjUNqH5IisSIXtU1/cAT2QqMay1gtTzLmEZ0wOeRBATyn7Bopyvpp
j2UR7dBELMXgdzimhNXElO5rJzrmsTIypgNYbSwgPHyAiFFNaHFCyz4AWo9o
HRdS5arcUZ1jfYsU9uRYQ1MnjwlNyyq9hYOF9t9eODs9lO88mYfkj+WPB5mN
ZIGVadmD7sBXl4JK9eRcwuzPDsXXTEzbZ6PWhCyhUYff6yRV2P29bwVWuOuM
U7Yh27ezHhu1NYjXXR739aCIv9su7Fk/UB0H6X/FSyQxcFNGJK0IySyqT0Au
UCD+522EaoyaeHu96p+7PaxSGvrYtVSMp5eqs4ILO5bbwCdSODVHlKMmr6hl
i2QJTUJhPYtgJSKNQq4lPbrVQHvip77ZJw4mGbgF9/kqU7OFMqsYxK1wTdyY
+jEmBPmG9panueedXAXEdypzqjp6xIYhdQhO5KGpthSK4v8UylpBRFN+NC1J
lA4gkS6Wf1tutesPWyOUYqOtH+m/KMouqwfbpsqlRiOL+C3g8Li4K3s3rBZD
lAaBy4hqKqulYiM4JEGExUSdeu7sSOxRbJjGS47+ynpZBbCL19GKdLgJyfwH
P71fMo1FRdt9hvAHDchx1femelzHOLFagyMbFm2T4Hb8CmZfZsIHyjGCP4rx
mPoeXeCz0eyCXDl0oR6mQymWK55kV+f/pOiFAF+B1+pM48kEriwoUp9Q9acT
pXnooFlDwgcreXHpnR/NN9I8U/gjwvxlhNMOYyCh5UzgH7HCmUvJesPViKtt
rp/KvITJke5JwMxbSPYT9QBKK0ActanD3OfC2FdZE4W9F6VseAc8tG/wobcr
1Mn/TAxqB9JLVpahY8/s/AyVg7dcv/ahhNs3Yyh7g535793eWOvF5oHsDg0J
O8y2NsvQdkSQfqMHxHzEwGF57PpStSsg63XEh2bQ/VEI8Hi3D291bQo0lq6k
pz/bD4Jh760xKc86X3cIe5IHXlCTWtkpehv4CokLfsnMCnrp3VVzZWssUYVO
uDrR3K8dtPwHLknJq6f37+0RlF9G5yth8N6bKNhHBdCchRmp1fH2M41LjbOx
UXpVme6kDctGcE2DBgdi8NbAZLJaCvK3e6kwEo8pJHLC6qNpjdt1l7FzsOBK
PWrW1pOScqkyi3HZuAIUVTv/4QOqiOEJvu4kho6CiA8oQkCicOpSohmLYJFa
equyS/NeNiZ8NFNb72qV1PKqKDMzOxSnrB0Iht0r7QksudN7YwXAY2ZIVWiK
wmQXbxbwDyDIohQuJxTSy9MXunpxR7i+yr7DdxhWRdME6nNyl7kfqeshNrXk
p8mb5Fozh1a2yVD3m12PVksjoz7SGV1PiMRZSsnPRyxvaLZSQxVXqrHbEFpt
zpIY/KiXt1SKmWmfKim6fUAmaKOymFICfWPnlo0EE0y2KFio6LT94+6SnMfN
lvUgXk67K9JZJikTOOx2eVGBdZc9PJv7jt15JAWQxIqjC5JZlbg/vChlG1HM
ncnziKKOYRw1tbpqIaMzCJsyC8jLKD2+M7gmwfdmSeJKl23YvkV70IkDCJ5/
9Z1EzO8U5H7rFycJ7hVnSJeIk0nZ8V7lhm3/pvPz8lcEAjj0rtbD6mMO3KXN
tDcDZ7dJTGkwNu4TUTqDCuGzhHBs5i5ZGyClZDhIYfHVYiVRGhR7DyA8anQs
Vwk4b/Lu3QubTXv5sKeOitKsRs1HtLr113rMJTKAtvQSmOIGNYqAeoKoMSdi
hrAr5uDciKWugG6w/ciWua/SX+V/O2HwRUAoD6hUyO7AeNg0YixwlEcxZ3eJ
ttWkELFB2FqhldRIbKKa6td1p3fnnYrtYP8tWxtFSqhBzs6GAIfu315kFNyS
L00FXr6Xe5OTrFW8pjHWgiR4/FBEeyNdPlSfRpL5FyTnJ8GIsAamRID8T7nk
bE/rv5XYacr4ilpEL1GPz+AfAnaaUtZah7Tb52/DB2IvKkPZXCpwI1OtaVPp
iXVYBofiRyMl2D405KFCAy5AhZuLFd2lbIKI3en5DuXs/9EGMnfZdE44GuDB
uXK4aOgHbtqaZAR5CrcufURupV6QGPtiejFCnmrTV61RjKrJdjbkQsmT/Z2N
x0qDdC0MXJoF/yd6pyrpkR6eywqziXRMPXALiuqelCpMY5fHNCeuEI2sPGWx
VZPmmQsJ3FxGHTmCO3KCt6lg6kIjPKYBaLDHB2/XKHFJKB0BH+ZG+RTNMvnB
yo/OquLMe6JNT1csM8KcQzNbTsoDjZMwy7rRw+8y6g6O2ultTxLjHd6f8A/U
RZVOPVEvb4l6L28kRHd9cEvfBEpOsjt5My/f7YLwPi7b9T+bRT476BsRiCg9
2kfILRpBRV4ZPuCeOJWpWSrK9X0CtCKTzTwf8RG38S72ZF7eNisoRJUVDQGq
67x1dwFh179DWkVaRu0QRYA3G3tnXHDlmcOi5YNpoEGmbhOQRIZMYeNyexYX
0Fq1hljQlZuf+X5gLR1r9BnfidE9QXrDe2iZFf+bu8NfCFM9GU407cAn8Ztv
wUt4v6k6EXg71QImxa8f6DrdElTRFvYbSLdlBwY3r2m96WVnkoXlffICKWX4
iXBhuFgBB0tnDUEfrLSIH18TJi+/phh0sTi73ZMTKPQajHkPgv2l7MBtjWyH
bvN8xLA40AJUihpSrdoFlYoXHC2EaSJ4h+N9cRH/HXR5YL07dZ70vto4buXv
QfReDQWwoAPvPU9ALj0JHhRDn1BG4oi3sr5Y4S6jVKNXYjWbWFUsPDqo53vO
BvTUez0VMjbMzvkEK58ylYto6JrL/CtnYT+NYRKWz/fnQDL1u7QHQqQUrwYH
PJGC2Qg/NKiB9oFnpHwIPMGxanvabPEHvcYZwb/JG2R5Y+X+XTlg/jQvsP/5
S2nDAnHPuSEUz6qHZT+79kFyN9jhX4WS4PQjI7WI6l+8FCpzwGIq9v9Loy8r
76mSgMBuxzLah1tF98ma4kFLZITxi9vEISHUFu9U9zwip0smO0uMHSYbH8rg
FbfemUAZgmJUim6m2VRiYzGqzjVbGtNM5/MTmNSayhivcGcVRCne1Ybkr4Hj
DDzQnqz/uWi8ni+T1j5tN/hSz9EP+RO4hAT20UpshWW6xG0orRzfnA//s1b+
DZ6+SzJFc6NjuRTyvE3RSpBcxpbEajyZpRqoKJy9fjoUZih3a+CWxofKcLrN
cXXVS3YBJhgscHnRf9HWDRZbGQmoUr5TORuMnNIp7YFanGL9TVmtl0+s3fkD
LfHOD2+OOK3J/vULK7ALlst82h/UyIeBR7XSwf+jNglTXBsknz9jeNXjCZ/D
dKU1/0sfZC3sBXYiqUKC4klzi3R/OolV8feUClyhZrTyLG5wyXHFMLyPjeXY
eLvhHE44rLew4p3iXBCZUnGRgFFNxDj0hPh4jcyRic9exnw7iFIZC5nW/z7c
mtdhpjNtTMdQnw2b0TuU+mldIVyGr5n41sRyl7zbTX31dktQ7+RCA9zV66aE
JLMEwklLm1tgZxv8367cyJzktkCRBG/MUok/6IdpPA7u6DTFJ3BU3JdXK/sR
yaG3QJ6b8NjdQCEMrJy1GGuq/gSEuSK8VbpUt3jtBTibOF1HmBDjUKxfHswr
tnB/lparzq0jBYiAXO9TzcW3R7q41isPGFkxDzXeD6rdBOs4n2M0QxG8dJHB
dLj+hKWWE/1QDFN342H4rVFa6fYq3O1mSyIHPQhc2d9CZTx1uNzITCGgT194
Vd3CT6ScvusP7iY75wLc/HRXwfNvD9IRkVPJKr766xsEqCtcCKJDdLQjYY5Z
3lI5B2cRnQWQBUq+ylZDMTlvzA4x9w2y2UI5w0MHsWC64sj1ncV3GY6Eco8S
O/8hXa2C17XMe0/1CvlQz6+eW2aIAe4R/7i632BeDTfI5igbZpPSsOv+cF4d
JjnuP0uHXlE++xvJvHKxtJB2X5l5+BWJk1rs/rT3ZeBW4GBQcfQjkc1uKtfI
xC1pT0PTIf9JyfbBIbw1h1B4SDZhMPUx6dwNjhDSzbX1KNF8aDO9KYf12O+e
NUWkxr/uPMP1wNgRFkm6TTKwVZUKCvDp9rPN+GHg+lgNvaj/TFAmoQXvcZUR
+4LWeQusTAOE+HIl4b0rAjRiT0yvw2Kj1p3tbDilqIpClcu37XdUhSAFjTYT
M+PCbZbmN0Vc0vxp/G6OwIO/IkBMG50c7y8z+gxeoVOocnK6htpzwWs3MZBJ
UOhTUEZkA3zF8lEmrvijqqwiXrJilyEAgoFIMlnbkL64wgIWiDIFZvIy7kzr
8/YiK4dT2Tt2/GkSHYCY2D4PdYpvKmVl8HpPh9ZBmR0GoVzuSC/FYV2XUfZh
uy/C4tJ2MjFuUZ/VmlHMMbPWegWTEifKqoBz+K0+/+DgIg0JCdzkeo+HTQqC
m0eicotstJL8+om491/OOHSl309j4m5UT5ZEpN0DabFrYmkAwhjWC7IxH/Ha
K/pN4Agyeao+a36W9bJnWSFh7fAs/W50THzg13nvuWvsU5W9Yr834QAS9NoP
pEuGddeQNv2iIvAbLXuXA9yUBrz3JeNrX/bEhqt4dip27zC9E//2DZDMcNL2
3pFk3q8Wmkevt5FL6BmT7xbdejUu7cgoioWRajV+QIvSh287ayDYEUqQ0rIG
3HXFzmgOFogvbx8D2UkzMRricNKFS2CLYhDm801eognI3wg4d2BnX2XazgZ7
Ue3p+veWtXNnx2vRoiqA9Ma9szkacIQhrDiLJH/GymEcpgCOhQ3+wMvxKm7D
hVgC2g3ldfjlc3lobjXSi1jPj2st3AdF5lkSqPgfVek6jAMZvYuZt5ECzbDP
gqvauOqBsD0iYhVQjrd1JHMo0Ciwh0dHA0Ql8hkmxN1rQtHI7FBscqRZUXx4
b19eiic6UW9TqGzoeIAUYADXNqYx/zkwLOHGtGv9g4MlQwwy3dO/VH06Z8zo
pUaNgBQqWjQCV0G5fWWd899z9cFfjXLaCv+1nB82DawL6jPSqpEYxl/tnes8
IudXekZoHeB8jeH/4IEKwNf1AV4c+iMrZbVPC3HwyMw/n3oFbn+L/Z/WdYxR
ByXK1qlGuPfAc8AFyCWE/lDkkvdhQ/qBsoMWuL0fnVz99qr/dDvk6GXL/fAI
8lekwpw0KJltUbrADx+Ejig4tmIY75akuCnx2LOhlOsj0+nfLMery82+0Ftt
fGepVPvBypfa9473KNf0WYHv5r29TFW5Tc9KYNB0ZX3eWfDoRPc2rWZ7OLOo
H576HvuhjwWZr3DtKOMZkt8HNRvIB6lHsG5YZnsi5avCZKCRCqh/t00qM9+f
hDI3ALQVe0Wu+LXrCeRblxfYg0ZKd2K1l5LP5vbs4e1uXVAc1JI/Nof4XNE2
iM8V0Lwd9bOOozBSHs8xa58Mv0QiI32Q6iha7HMg8ylNXj38BTqhFdFq3eVJ
iFCY7LWcdBe8aJxe4QfEBmP9k2hmljlTpJMagin9w3VBRyVrAjIlPEeLKzUR
gLWLLGBV2vvvzDl5oMoNNIEF2l1ALSWemUgbyz1/MIAEDYDwgxnBp/jdDBfG
EzyCzyI3VOgxhVQlPV37l6gV+c4TFdcaf/P3U71xeY89i55u5tiOXhFbyzcd
rmRfdkZLEOgQ/W8X2mVPCweIqSMsUewzv1YJi1N/s0CjTOfX9EDsHBFxRiGl
1hvW17uj/N9/6tyktsAwSqcuCfkqvxgdmztejcIUedPhP/SHW44AogpgUrZJ
23r/wMFXqAsjyC9hWC2OMeZ7I4WpHUekuzlrHnt46hnhdOIcz5Wqqpo3uGeK
55vOPvXXKqg1QTM02cRcgoTSiM9VeGx+dx+ve0AUdPdNUEYilqccXrVPimdu
P3LJZ08mWSjRJ0NmsXx1YVOsELVDhM/waydEh7VNQTHLNeZWSZpQ5D4M5aeW
W1C+/6goRCccjHPv86WPTiIOjNz1kWb9t/om6/LkXOMEqQRqs3WBKPhK1t6N
xhNwzDURf9L9vcRU8PtI0INHHn80pJjPBiw0kM99h+qWNDmrDz3yCp+6qTFN
FYUGply+VxGDpEQwnXNY38vSX4Lx9zQOch8FUL1h7R+DMxKL8QJJKvUg4jJF
+epSM/7lrEcQ65Pl/IB+4zfJ6PvGvO7ruHSCWHq56/mtRhxI7P5vHNzGTsEU
JaQYOGMMt6VwnRKxwAqBzx2N+NIMy9ZhPwIjIG8evNGn5LjUp8BhtpGSKb7Z
EF8RdVZkg+pksafH+3tJrsUJcpAIglvQK6HtoBg9D8W4BdoGpsCwT5Bef7Xb
97cQuCLh7OsmfymNoZ3Tx/qcaGOzQZrb6FpopEu35hSUi6e0yCBPtOGrCG0+
DWjnbGM77x0VgBmmu7MQwS374+B74GJB+lOufOgLQ/c0uGNrOQoImtRbKbnm
WcPvUbMa1xMhvOMvaCEEFnN5kww21tIdSzqz4ymU3FxzMF/XnJwcGZKwAMUh
N8NG/PoVn73CUOtOko98HA9Pn7IWTpdqhU7Tf/da70pk68OaUZvYL1CRyQl9
bUVdebJyJFUe3sPw6DAuqMhWOJ/0mYaiZ3Q7YQ7JdwvZAZyK+rkVKKaUILin
SE0faUE50a0zNjqeJ3Wz9DtYY90dcyiBTiN/EQjfrTPMxVO4zZEO1r1CyfkK
IXU3MftX+CNxIX8/AM9IFca0HpjBB/kYtT0Ah7M83GmQP5r2BYM8XTuudWH6
nJoD2oIXTOmlXoX57Nat3YBTEK/4lYd17zL4rzeUltXeY3ZS3Eqget+6HjJG
kDVPAZH1PHyQ/4GJDLEOzWSqyt3DRt/WJB5FYeOiFlmfmIqIhV43WpMwMxWd
9Pt02L8vixWZHUSqwQg3cbWXwYpLrh0l4hD2VGJ40KvdPdsfw7pS/ej4OGUY
VrsCqcRm2KOQceav+Edm9PFnQux4nPRt6/5m/8OGzw7VjyRFmMC/eQccaDcI
frAde0vPvBjgvoIen08dqV7AG+74v8GeH/CClvS1HH6UKDDk7TnL5XzaEwAl
+VdSF8uPXqTINRXhJACLye6C9tuOE6cIyFtEbiUZ0jBR+U+xSV9K7klIO67O
Jt4mXoZJZ6L7PK79eCUUZk4P+y8n0efft0aVzUIRm5PgnWDyv71LebTmPP1j
7x5T59Oemiu+vcJTBBxXWhDS87RTGSAoOVg89zlmVgQ366QRetGmwkAdr2B3
5cLj/bHOgZOEe8bwxWfdsWiu1X9GVe/KqFuG+u09bGgu7irgYfaIauV/KhvR
bSfm6dlrnuFHDwyQkG+LwkxnFuaRFb92qvILLsxApwSEURL0Yda/XWjw2yPn
kPJ4TmKD+oSObwj7UgkpJVlbopF1ISRvIwr7Alv8IuWZ2Jssj1DmyYbuhpb7
BIdS34zb9LX+77LgKIdv3Ivlp84DV0C8wdKzYgLUSg520B/1CVnvL3hU3Ic/
/hMwj/YM9K0A0DpIpjDV8eR2QskiE9HVvPMuK+He7XgcOzf7CBEk17kRQ0lJ
IJ4HsAZAXK2s4NpjLDJHnrYFqMMrdecXGLBUuzdEElU9dnJ2xtSgoRHoVuQl
Tx7bjjBmx1E2ABkEOoG67tzm4TfceVLH1smCSEuP+vXwlHAHV82uqXCggRso
8uvM0uzGJFcEsu1ShWmzSb1dhCf7kFTl7C6cr6GLSReA8WZYgc/qNGQij3B3
Aqhlq2TZ7jzKK8DwdSVp/hM+fdhiQZEu0rxHXYutao81HJbLX4l6paBoApz1
g0ESJ1FbyoHlFm/Tuh5j99sDElEPzxFfZyfVtb+BT3TSo3NjM0olum2IdxyW
3ksdwgTbTsfjEmHj0LwpHhd3yNNj5nzWa2ADX3wb4ZMkASoJiPYHquIlf62L
bN3PLHTVQ5szB+mW3YD9ZjaQKRb8Fxu1huakoiWcew1I/KeCGqeB7Ezrf135
l3oDFh+8ojbBBNitroxYMIMvvHSc0wcTzbOSNC6GPKQA08QpcglQJsslZzIW
KAcgxRfu0xOjmVs/K3z/vhH4lfztU7fxMmZvz8NXv1UCgpFvZf4wDwGiV6u6
Iq2yyPTDjuFCMbhsu4eFsbT33lIHrbLt5A/vATLlAyVPtjBlL9930ofKCthw
Y+KJO39AOaSY4/YhhVHkr+5ho0eLjh78Z6q8ZAfawhjz7aeNnke2uWiXAnQ6
GRGOyQtXDh9MSwK/G97kfD7XojmQILZZwOWpEdTvIujYntHk5qK6mUygVNp7
Ee5trTmFzlFjVSp2pU/eMRPSEA5htmixPoJMdEfWQlfISquKGtSGukh9vuVO
9pwtdJKtIkpABEl73PkLNCpRRXawNCCs2mw9Rean0FM3I6RaXn+MwkAI/CMr
VxhEvrIPPlEnAp/nI5ubdSWxQDAy92GJW9zv6eV9aON2WqYOQmRzD/Lewz34
EakDtAurLqzUIAaFKXd76tWDU20KbGUj1TxUWPMkDfAk/hyzXHTgGULsUHhB
0M/7Y+ctpUXDDzJ2E28NJv8eoFf1S1h5SOWvcyWY3W3Pmu7DzyFNYHVq5AI3
Y0c193nB+cgADMNn85JFIKttN5+wfYQ9NzbKDLdeiNyLoeWWH0HJF7tve1xN
ds7PE4KNDuFB2OIIkPwZGY5BFnq9VaurBTmE06XyLC/iOaJUnNmVsusW9TRh
18rWhWEPSQn1yZIssGT5gwesjJbD1/8IkzTuhJZbhTIzDP2Nu9lhg+mlwmfg
eul97BZ9RXInDVify3sGjD/ZiK8xf6fhACyVx+zTEf3/qEs+EU1/NB1/oCbo
zeoW93wzQpBURz48/nOqiyBOJVCYhm7xsvmEoMzS3MKiV5GNEbbI5pgv8F7G
0vzUMXOtYv1w9jLnIhyi31GOef4zFSs611rrb2ecYQrb3bHGgpznJlTEHrcw
mPj5HnUXOOG2mR1olp3K2hAHjKjqusWNwo2VqobzkJPbJJxWG3hRh9i7aO09
+aTiP8UAw9Kxqs4y2xawsOdb1cU6kmP0H9H/d/inkcsSyIFEbtVKSkNL+rbV
UpSp1ZSXLbIXlpFIZHIcT9gl6AUcYKTlDDaHZ/29rHDX3Gv0l8i4vAtLCTLS
/jovLTqsX/+cJhFet57lkG755vX0YjGSANjk6wNBlHJHZvCMWf4nwpdhp6YM
hMzZyesizuT+69+uWtsDr5tMaVkPigA+mgSRTkuj+WjSQn9M0vMmO4z9YAtt
tPzBLLKuQEE3gxO2BLRQJirT0WUYzTqITLUyG7BMMPtEGS26+A19h6/6Lxzr
P7a/KYY/xdtj/ySrkZdf6u46lby5DozdHlM+2TGQ9RBVDO/QIlk4YZW4CpfO
UckhRpVy5tL/evckYkIaGU2X/YmBytPU2UX8GoJ4zioseVitOrP46TTsk+Pm
/pPWlCSYGXBfbiNotSRBmysd2lIUloK7771htpS45wl02ggX2Pi80U6bC9mo
SNhq7wNvabIGzqot26K/MgFWfkHujl+vNkPk7krsXWqktdJDvGx2msr6d/YF
rDrqyO3xqP65cL1TRquJV8ifnNtpSHi4hC4ZE0qo60L8t5bQkVr/Xzjrn2Y0
G7okuRQMsQmJHHbWYJHAFGGNiTh1tsZ53fMh2aJdq8/c/Y8ZG7hPbpl+JfB1
mVcby7cC7J2St8/XYDUH+/ZU/G/O0WJlaIHLaEv1BqynnvcEuyoUDmmbhW7F
2xc5U/jbzy2REjqmrAZinKWv+O0ny41/3M5R4X/kVo9UW34mRUQmSBZivoI2
uMeJDaybKXemgMjGaYaqrl0DSTZN0R9+HgL9AdKm2RQULHwHcDkhaGT9lEg7
hzcqI3oUKz3/EGT1NaLGA/ejdPVnxlLGVU2DD/BmQrcEZyp15wmbcbF2a788
5bHNCNeP6wmBdQAqI0H4Z8lCHjdftYkZxFZeLAdh45U0OYxYs30OUDDC9LES
7lbVZtnXC3sFuDxDfSOza5r1X/Sh7rVGiJt5tBJKK/l68cTyaDrkRnplan5X
k/udQCtO627QB7WRM93e7rf3X2NVXsfWd+HBOD5PHdXKPcrq4O8lEi2Ma/rh
tGpjMAzWsG47XMuBXRSiKwoWpuTR1nlnTRusOP/Kt83EQQ3+AOit99/ArImO
mE3a50URX4fC8ThXjbWv0ds17k4pQv3OqBfEZ8yUgnkDkLJfMnI66xX5SQvi
Z9jb5XCd3XjYe23PGnLn59zdS2MSgMLi4ePWQKzFrc4gzLMkhjwbW/y4ESpW
mUkVA+jV8Wk/lHQy7p9KD4pyfxrNm55X6ZEeMixby6mZCg9ErJCvHshsnTV2
k4Z1iczyI0OUSkZVkK2b4KWAe7NuR1Fm3FRoCtsv/e7yIyHzYn3x2yIO6n0c
/QACdBFK7WOCU2a4589EeBXHeIyXgJI0lLFHvVMDboxnKagQoScbc6e5q6W7
mB/HWohXdyLBXBm8hywXf5BgN4X8p7zrEeLAjLf/hOEQUVXCJn+fABU0bLhp
SVh6EfKS4ocOkOeiVKYUhdSC00p+Lplg1cXovUyQRY3Yl/3MS6yM1YOUJlJA
J5/gw5ikw4Fj2f+QdDVt9bGOZN+cpDiahjXZWQc86uwak4V+iGIfbHMtNBT1
QskMOpoNJzxib7flkWtIBIDP7MAU5T7imqHCK4YmeeF3tkYIAVWPvwEVJDa7
ssOrSjdoIdLglSru6/II2Zs7dX+AIH0HFM0dPW4afFN67z/fNidmUYbswZVQ
aZln2xSHlefcs36dPaQSawgLhryRnA0PPswd2Qcca+57naE7idmxHv6LWlHP
bBrquQszixUK0ecrZluGuQPTDrOT7ca6z4ptXT4JbmxckTc7iFMLK5aEbIXO
/q6naeg7TPL1zry/ZZOf7xa9ntAfaJBVzjIG9244O3X9ea6ULSoj3KX4rg0V
ZwaE6bqYJOj95jGEEhOCfOcPJpZJamjJ8cyGmnYXW/hT4MkdPKNlPX2yzGrI
cT/4TFAbfroZAlNYLVORPB01ONtcr3j+wm80fNgRjb0wGJA5U+rEKP9V14IP
y56eFHk3O9tY0U9GsfNOEd1KLwEenZjoliTL+R8mn5CsAzVHeB1D8HXVSWam
Qvcw6wGGPS3sZeaerQhg/bg7nE5kCZfeVU69YPc5NLsojZbWxJhNR55JrNYI
tO0vexqKMx0wBnUz9X41nNrISN/52BJjY8pkHU+yiy+CzO68M88N8BhfPtSA
m0ForBVP0NA448RpwMdA1FHUDn3YVJmNKG9D0lkOitNQYdmbWofXuoRCG7n2
btyGBHxVBGwlfUcIA1//jGuEzyly3F6YaI9ynWhOKy9HzLinTj+Pz74Wr3iY
lsUyQh60PCwYgcXRAqr32KQd+eFmWOZQ/b72I6U+3dkc3jZth0mjZxWJnfkZ
SSPGc/Kgi1fx5H5sQ2o09iNV+BB5NiLwFv76T3tXjW/Q6CaPCw7RsRNYgSpJ
hgRdrzeZURwuEyTYydUzUmfWQMuENKGIlV1GXMLnt/FB0VhlFAa6iRNbU3Qv
7UA6/R+gsuvA+KYGnZyBxHdTDW5cWPHBZLa2kmI/SUH1+hJlwqgZBdndS3M4
Ffsa6OC0Um0ntAPXxL+BqhIM4pv6bBV9PpcOUNNzuHV51rYJIq+hkNrdn4in
bfod4V+9UZBOcjgrmLlJj9e8ozPgXDPxoiee1yYT9yLBNfm8MKQBkaslXY4j
UvmuosN93nVJqleRMcAys9jU8WlvXMzOUvYxB19yayG/HnWXWzyUDqtqEmMh
pRuLLLW6YNQa5pgKBB0wot6yl+EToNCp26rj0lQvvJLyVBO6xbZY+snjFuTm
AVuPmFUTcT5HM7dTyIbHOezyq5XV6fI86MCB9I4EQfyB+JzLWLUFuNhAqITG
jIePJ5572RExtq3hsc985CAp0+vba26hgFMp4Z1UWTZtrJgC8g1P1J84BI7L
uLNaUvVxD7KtWqKo1pgZ9whmVVVZw3uh5IyWERw2gETK327rAT5MCQq7pSTo
WvVlB3WaWFVJcHVnulUN6SpzxaUfWNCAcI2CIaQpSPX7Lvku5JYML3xWUr30
fJRmBPhbFobPZpw31c7HDw8wtzfvYXRzUX0au00eC4RoJzYWyXYTkB1O4FyB
1P050PKEoEqQfmRLQmzrv+3PGmCxSyQZCDDBFun7CfosIwWEbfvpWHxTPmDA
d1zQEkfD6JeBsbcy5UT3PISGaCaYizocAl3ZSYf914lRElLPRxJMY70yMbg9
UQ0pkmx7qLhWqq93irMFoKQQAjAJTh5GibUqfR8A68zQOD7n4BBC39bkxyVf
jJznpfrz96qBBNa7pHDQjI0QTprJ/wGZIMfQpLBa5n6nJlxY5EEgSTQe7Tp4
ZdHhRwyIB3U898hMNpgllX7iHFBimUONlz2keq9fcAyJdWyVIERq2NZ3S6Q3
RhzTnYXBTfwIME6sty50t3UfZpLgTyN4FAzIC9cLzHEpUDgvh6PJeJ1OdgL3
AOg/CLbsAcihwpUDnMun65CUAXC1YUZMN5coCHYB0WfUWDkWYR/kULqW7Kcz
TSvoXJvrE+49m0rty2aDalORsjBSDjBBxHbQCtJGwM4V7qAvd7JhhLFnM2r9
Hk1aopTjPZYCOa2NCSTGQ+vCv7ZlRhoLpICGiWvmIjVqa3eRBMExZkgEp5hN
MQL1b+jtpzQimUD28wu4rC6cRym9+TkKsjPerE4zDQ1cwgA5qVJM0R5ISTSk
XNqpMY4uDB6yETkJzX4jxO10gWWQuFOCzy58+DLI7zgvpMdVKGQrVTWCSStA
X4Krnp/9ykM9x7BTPVzkHeqbgSPHt5mkQiTxLAuulomp3EuiMiRlf27IJw/o
UoF1Uw2msqGq/MiO3JKc0podk1FkOJTbxA2oUAmVh0vgQoHNpkE2prWiE2CU
B31nE8pg4yaefm54RZLZDpeE4BKHFur9IdoamPPpXn8yw6StRC6s9KP4K40d
BFLpc3fFae/O4jjGLAZ9QawFHnCJnlOmNsGFLe6pSJJgsSZuICRoGyeofwqP
6yR2lMAYIcj6AGorY/9AsH3aPrrCmnVzsE+iTPpS+q/6MNsCq3F7Ke6aGUw1
SBH9yUsaztWF9f+bJUfk1txi/KPHzk85EXd8H/KAtIrC19oqvQpowJp5sst3
L/mhXdxgpGXEoR3PgPKaiApxuBWi6SpClYElVQPtQ7VwJTiOWLRnR0n5/iH7
4L/vR2msRR7AyjHoVWS7IULtBs5X55fjRz+7zRiFncYPI2dZKGPIkyWdj+kw
3zNT4suF2YTP4KhYAu6zYo/+r1nJo1Nephmx5kDcaef/QU7GpOdn9LyN0qgs
kZc+EZtzQ7BGHlfVu7ciVbgLxrhHQy2DATaLFDmLLw4Hfrsun2dy+6PTlcJ+
aGW1w6iypktpfRQCpECMtmUyNJTq56X66zkSCs+ozrCqQcbGfroKnlVRgNCu
DYHGpLoq8ByzA7fFXejRnGvsnkpswFD8CWufWcimM0SJh33+kJgOCv4hmOiA
rO66MfvZ3k4LMo7ZbdaZ5V5wKHGtAAfGdNYwqHMnFrU3nhNO7QEcKpjSrB1g
RjVygkMb+6VJnLGdLtz9sh8EY805OpmAFON4tKJBoK3txw1b5lW7PoH0A1fP
i5K+j2Af2cIV2WbP1+2tx8sghvxGuwuftOWNyCBddkmJ1gKXdt3H3QtlEdE0
sYptw6drxlXNPvDAi+39CC/M0+73RTy5uuxbmav6gjxkRpQr6GY32I+sPMuc
U9NJqfvm666JRf8qZHKW4/em4fvPiGlRKeXOQboZIZXOMhdE4e/eUAckLfZd
RYzrvpaSa9yR83f0skqwdvrsy1Eej7ADbBkCt6Vu5mSY/gpBLg3gaRjMuTpc
ks8ZmkfWOOZZmGpV0sxOFu1/lno5285XP4BJPVszr3ll1OTQwUwyjvcsd402
bBDQo6ino7Bak/CSV80x89vUQPfWubJsIqEJpvRSXn6m5t7KKUaQ5uy1ZueO
rhSjv2zgsiJhWnFrv6VJYnxfRsbxa4U1+g6F81Fmz70mUVHslj0dPVAEX4Ck
7KJ0Gwr4MK9iJn+banePPFt0UZRaKMXcAkBmo2vKukpeDbdt2UEI01pmu1gf
cJaoM2qE6LtxQNrb8VAaXB43kkobGQQB6ay2ts1xNYDlwaP4+ByAAuKyRmJk
8UEdtq96LNfHVe0ZXeEE6joMJuQbRTK8+QuNC3gUpvQUYsXmzhM9CAiPKe/m
rDGdhLiBaB1He0VnY95i+GwmVWNml/lll15vrcxtuuBHKC1o0zPsPmsVGKVn
u4xiOde7fTZUL5fnVCqEv7xQhc6GW96Ky16S5FUz0u1DUfe1luiFn3Uc3eGm
Xj5z2mdE0N+iV9GHS+R4L8xqgpd9Q41lDTjbojWJg9OSUiACH6KhhJzX0e2K
788g6iNW11YZz3a5LHBCJIqwicEvNYJMY+M4gF4klkp3L89JUysGUvvShoPw
1GYCo6S72bGL2x8UYDmweROmRhwQxlDqpdheogn08kWqbnSVO4fePI8jrJYC
1CR8DROmu0QHVD0zjaPEhlaqc3esR9+Tx4aKrfWhPuK82NatA+mmwRYlCKT/
PJDuM5If4ySQHk1XX3BKgIWlGALtQWqmS/AItPDsEUZWE+K284PWp4KNFcxW
jCA9oqw4GEZLOgUg5aOSLm6e3QFkeOj7R0BsBloVDXxnrI255mLh6SFYh4hi
wllGAuBhPwtcKceH4xXh0QnyC7yiOzGn/MH3vKlWAIRQKH+vnek9PRHgX8Dt
H2bCN9KVOfvIMaujywhYU81+HMuXQYMRtzRqC97LY2cTkMb75or9G39hiIOh
Tg0HsXPwpLzza0kMq2Z7868KNiW6Bm/7/+wWeIttOL+e30Y6CsroiS0YO0yb
c30iASWcXqv7MfPIm67NIM/shENicNI35ljSDKHa+GAYXTl/Xxw8auM/GNYr
cLNtfTrU2O6mxNNQdQQg3dyko6gRNgnIXfgGO0o7NCyNydL0NBiIajTNeY4X
mJbDFJ2P0VWzslR9L6Fto9PFsoce77a5E94OgdHHh+KXNlm6d1jxIMeC/jbV
26ECA6Cxhfuur48QdOd6gDoEWqIlmHn1PQyVXn8xI2bY94gGeGTYZ0FRutkk
7m4x8qkNj39iWP9dPA0pDfgU+LCr/qAar7qs36mxRid8LOvJkOwvQSkm6Hn1
SsZjqQDJMWzIb5mhull70QO2p1yj/wZ7tWIjmA00I5qVC6VdEk7xcNWbj4Ws
zRcYDBlKBSutvsKFk16N3qNGnk4M61smHlD+lbeM1swrbSheUd1xlBf+CFBB
dLdHC7wMwjc0QMmr9kWkebUqzibPv9pbhYqFJylxAUANTaKDG4SS/pTFFIJe
CQfvqoZpyX85hFO8tsM4WiVBn8b2CKy7uF1IVEYFS/EIFV8CBOm6S7dxUW/Z
dF9lo+P+GAnbcGNSdPVj0aDoBeOUKT7mlmVKqibPv2keylexCEJ2wJYUWr+B
CDfmGAjunonQN0ciUw+OB8bV+EaUaAvqEcaOSuRgiWh19H+bvbF2s2LGuQj5
VcnnDHVkTlufdl/toxmO2EpKt3LmVGiJiYwIhqhiUmS1C4EAgnF44TyjLtgV
3cMv1LX2MkrPVWI6knT3oEiuAnSzuOOClUXtVLF78f5c9vdEcZdNiopcXdFh
I9x3Bul0lqhm8MQHQ+0nnOe5kKplvGTx0SfOpbOyPCh+XpHJG4F4PhtIR//5
r0uTjJl1I0LFjwu3vWCz8/osXFd/7pf5OTrSeUhHUsPVDECK5A4iX92F8g2Q
wWaSBxwc/8E+NxDRr+UVZMTn1DlIyJhsDjnFWP+VW5YnmBHf6M0WkELWDhiu
boPH5Xh6o4ZQB7vEY2Lhcob00c+CobrKmWpaDZOiU9SOHlHBUI+sX73XdQzI
by9fjdl7YhvAXpyyRoCKETQH+zJf/TuoEgFeWCE7VD1wubhZr9zOke9k0RVv
50x//hWJg0J0ByZ+eEsnk9r8B/jHTMOMPD1cyc5vAObJt/QDr2s/84Oj6Pol
rWsGnShoBy3PNQ4nb9AH2n0PNNC5e2uAWIMHonaLAmH16kKTN9yZ8sI3l5Dy
OA6BIjK8Cm5CqOukQa0odnfUt8jHSEiMoW7FDi2uzWvJ8YDYJypoXWaKW7DV
dMggcR+R99VzVbzuiptf6sTS2YqibUG/FflZkiJFO3IOyDIz437XMYwkbqtD
+VE+1oF+vgg831HKoAw4WwUKaGnqSR7TqbvxvYTvVnT9d5u2S5UzJHt1PQfK
0fooKenqXHrL/N/4FXEjZZw2rxBA65FIJSbgdN41pEoDB9xCAOLMOyjJMgbA
09PkwjrAZpjRIYBcjz+r74rsHrD4BDXyMrmMjEdgsakcVz0DtLBZ8/6hte4f
zJvRAEtlHbr2T3NaB9UeeljPA/XHu3SJxIHTgPCBipqTU9QZWwoj4IijIqmr
ZMcbyxG9tS556NdL2jEcP0ZG4XoMqRRYvmkp0lqcr6VfcV2wlkFpwJtA57Rx
VR0JiWa23U+w2JqXSvoOSYblSW4gtIOmt7cyVrZJV+ovR4QuuX/qHKoQa9as
DajmvzqwbCAdFMDg0v4qJ1CdNboTj0u5V4/6SK8dOjqazTVB5+YPhA1h3Mkt
pbTWY+GGT7KxofQQ76k/C5t2kKJ5zkt7ZQfPzlVZqEB0rqeeas8tuuh8EIBQ
CfJclD/dbfDz60/fWJt4R1z5oX/Uxmyo0ZTSDaHn3OXfLMs5gMbNUC/TcIG3
ghInLPptrbLy1ueC3kcssQLWCp1KQ6Se4rvHIw2BMWOidKy8zQW9u52cBqFu
2bu+SkXG8nhFUJHwEyuID/CfWpfFkkriq4hBOoPFubPgpA3v8NXEkAmX4FPb
i0cRyoFuKBXd81JTWK0hKVhfFM+ejKHCCM3ZyCVHsqvUb2oYNSAxJUiWI9VT
2rgBEEWAJBoM1b619qSu4FWn4fDc0QDgIodMkOb3Z5B94sbIgEq0ngNQTHsn
SMqyJzdySUGLun3E8atB/tu5sFrm1h/HGu6wK0wxageJgOg2s5zYhPmGOqMJ
T6SCr8c/oXarQP8o7Fjzsmh8ESWw9ce7Yms6fhm8umaKp1emunQieWjFM19k
V51mLaUvYpjTfIcK7NYMoP/yIESB6DkyAiCoY31nPqta4BL3GCzWgpR3Cu9r
QrD86PGyzZd+Nlfm1oFQJ3Ua+3Fmtx2uxdBShWJM8bGip6sWXNU5NUle6ytx
scnRFF7I+IS8s81OcRvHmqhvOA1DUjekIyM2Kx7c3rPErO9obiEZi1tkPZfG
OkG2LBtgBCbxkY+bPZJVBctn2nI+OrdCSmoglTivqQIifk9O3Pa3pIu2QEQA
8dzg4Q5JpYgi+dOniCE9koJzTWo+rd9G7kBpg960mZ11B/AdFvDRMdpr6fIH
lTHkXSTRqt6uj3m6d83815KSxsBWuLh2w/F4SyePeaz5AUqPBAlz59BR8HTt
h3gU9lz2zU/CTe1Ab6tWs6sPWIVsBgCFKFLnQkRJI3DikTpt9jwNI+htg9MW
TwFO3rvIggMDNOMCvSrYG7G88QjzsOc4xIwfD4c+nxsvoaPPw/6H7bbOTP/G
EMfOjkPQSf9QfdU+b04kCzbYeLuw2mEZhjsP0HRiiP+AONWlREv058M2G9UG
E/2kxfIG9Yoaooma6jSigs8USgmXVDecoaz983KMlbByb8FDU8pf5CuNxxC1
BKN50w6cUp+8vskT6kmh2rqZKpQ14SyEP8Ygj2zaYlaIMfB+TdSl2siKKlDR
k9MSd+WcbsWFenyJSlLbx8KL9/0pOMYA2TTR+23d/M5Zf2bMaOoQFNnjFae3
bqioJ8L1QLbVSbKeo7f3UVReRVx14oilxKdHgDmhDDoV+4ZGE7+YhKZTjFy4
rCBX//l/8aqijR1wnxQQe1NLMudgKpU2DTDjrNwsZOHwFMy2LBN/JCWIOERe
u/5eJa0OnhKKjzxpQ2kOEdducF4X3ESpI7FxoF9Y8gXgoVraxbm39xJnQK6x
bhkyWgYB5sGZh/uQJDf+UFKODA+0E+Dl/ChyeSBdK3yOWWiz3Oc3UOJLK4nh
mPjzoMqFBnK0VAgpjXBXC9efav9DtwL/kTTh6/0R/M8XvGmTpvlJ+7/5ZFlV
cmwLi5RA16yAoSiyLyyHHdz6vFP+SpsW983I0X8tWboKGeHV58Xpw2vsKtM3
/UDXvCA+rKN/OYg+1TGWSXJYtyZKVOLfE7a+LvbwaDi9qoi/hleC5cqAafPu
C6COtG+1omTiIgkMT+Kyz+quwjnyTDNPZmZOIdGO39S2OQ3e/C1RTRnzcoex
fPm8qRp/6lCVt93WuoKJZ4OwnA62EVhUQclEegMoORgsp76hgB8Msf9ohQgT
wu4hFPFWlTA194+TDl5Y87LyqGCv0ko+DLE6ktuIJ/OQYQjyZoAIKpxB8uV1
gfMSx4HX9eaoSmfVuxbNBLvuZxvhebbG0qGhHQYLoyE4BdwjrY8XTXcMwxvx
khDcNZtA3nsvkR/YK+Kapbhfr30AkBqPfgdJ/Fn6xhqhM4ViOnSJuCMVKDrQ
MNcW2W3rqse0CSIunUCuuCra/CpOgyAdcd5ampL3vJJqp/rjC1rWTL1UtnmC
qpSfdcwzplFw7uYXKuAMtLlVxD7tgBG6W11gZXhwddzecWPthIymNBjoe112
5RKAQBw554N/0vRE93mC36h0yQetWhKO9VdefROfH5p/9XfOSa/0XE1q930E
vHUYZbhPR8/QAsxviyspvxZdISwEkDjH3eUS5muN0B8vC3svmC143bQK+AVE
KqUY172RvA9FamqnEtD378kcW1n9TRPpbt/uFlM3IT1jxFMdxA3yBzcMbSlG
oWVoe7x6JjpGvbx6A91BbhueXe3flx01JCi/LFMgyMpoeF7N92yt+08b7jTj
rkIFnorCbDicurlRYtIICpczaMreIvQJBhqyS1B3ZQS4WJMU5L3HyBc2cN5B
3UmDrBTLlIwK8BucV1/Jukj1ugj6W768OKujQLl5kDb9CHHMKQcQNkmmSEo8
1I8tRPN13uwKBvH4FdMdKaLyfuyZqccoao6Ok+L47x+D1P9KXxeHcC9ZV9cx
rYDbctkBEd3UjPkhGiYMIVu7O1naDY3UddhPKdritMtmw5qL71JoxVl8BKHr
/YqUaZAmK4/1u9AJOGVocTIeNljWylUvLOSn6I3KFa5DcMJtUPtaMU/FXkAI
byoUDURbHyn7N4ZRVMADAit9LLlHH9FbV6xifZ0keHjvPU350h8anbvmsg1H
eC5MvotyFxs4n7LbO4/vitHxf/5rHrYl3YGE0MdUMDrq+2lI5oD/tbRtVTW+
+LNDDS0WSYUITCWOzvkI3TxqUapKdRfhE5BMmed3AnggkyXjSALXI5L9iLvn
L/ur3ISZx8vXCuPfQ6QFjS7HizaFXiD4f99iEI7CdlIu/ykR5uzUxYo7Z6WM
kkkzY5zNAAjMhLzodzaqrOre6ADwP8TCQEv9x332qT98mxq0HN74l6wV6UB6
C8UYQ+DbwI/1zYN/RSGl1TjJtX/Hx3bGCrEcVmCShCnkq+Ut1EG2GxA88FnS
EDnKxd+rj8imwHPppgbfP6uUd0I/797foi/i7cu8o0pF17gRZ9/1bqYK9Vhx
D+NpH1HgtqSXOLOUpdQnOKrUHcuDqaGb3Jvm8LgvPEJKbYQZkgWvw1iMm1pn
6lsFxYkp2u/WE+vRnXOC0jckVDJFgEIHa4cbuJM8BEkF5ya/dRrVcjoLH3WR
WgWTwva59uC6l/lEhHtJdKtXyxnDxVtwu57iMwOdxpXOyP2iukCsmFnNkSXW
VF+MUnO/E9RnGL2LlWR27pBXNYdqcRoUK3X0WCSIZMPxyiEIwXXesX4flkjF
+dc0+1enyy/+T7PNiBQrMR+oTCaMfCMAnyREnrMg945h6zACvbo/JW0pfq1e
jCPcD93P8VOHa8kAYWdxFaC71nUYg8aD7W9JVQz5ff8+SskgXj+qC9vL4Srh
GgSWvzuYLglr3PMjYIz+DXdt+tPyow2Dlu8UVRf+FPrzTEuWCyZizmZxuoYr
t+NGM81XrNhLRv43S0ja03Z90IlP2zvi/REpHnl71dpQ4m2J2UrcGmaQPF99
NzyouVPSsYzsVbRSLb0nu82CY/Dfg+lC3Si1GCZrc6RglKQX0lGj0GOBavTb
O9NOa16IHOQMSM7tx4uAaF2bnnfwHY4QtNT9H2sL/cgQDXYyqGSeOe/sgCkI
tA7bAWvgmZ3fQklAIniAuixqKEtwEOW/qHwsy1ypRMcHZi9j0UT7u3jBC58Y
fdrqqXNC4kb6sFpqYxiawyeR4/lsn9pldvMSHWtoVBE020Q4hn1mxpaK4i/T
e2SPGbZdRn4X89sNBLIUZBntj/2IeG5y9y4xKd7hSk8RG00SlSoIOHmd9gqD
pwc/SicWbP4YaSj+yvHc612u2KbiVG2Ji59VMFVGX8HcjWomMm4vP7OAlGpD
dqCqhC/eY0LBtHnJE32x0OgAtiOuKvM5lZvY+zLcURDouMjLBRO9CMPPkJGH
r0xiayPobB2peymQ4NDuoIK3wX4HAovxD0A1

`pragma protect end_protected
