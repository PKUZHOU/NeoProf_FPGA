// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OtC12Tko3HVeHdyoAmE2+sxjiF8XJJSY7SEtw06uWR714XWMT8hTQUsCGdmV
3ZgWSWRKswgti2CmHlZbrenwqPcJMSDjxEolJRZZGx7Bi7SmZ2CdXCj2kugy
ZYm0cC/01/sYbThMbco3bdG3IKnYEYwNs7LzoxVhuNO9CapZZ+ToJu0bM37C
W0/2rTAsO7Hl1y3hbGZcAsjp0mgRLzqygnPiA2aSpv01+67xCIafaAsr62rL
kwZhkH7Q6WpPBa9QRjkvtJkutJM4xLgswBo9MqEhtwWX2HbGg32HHJ+WtHvJ
qHZ/mznKdID2/Aq4Huk0KxgiPDogB072S4Z1KvQaRw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OdoYLNbyyO6I9pQj9v2Vda0dTlH2Boj5tQu7Rk9xZQd7e+iJUB7bP9KUmYKj
0J+MtYzUEoQ07dxtC25BqdNewvxskkKXiAPO0OsG/EHx6+f/tpjaS459Vn5C
oKAzLtUUT7PP06MBGNrPuJdyG6hqSeiYxXBp5GW10AqAkxzQWLKc+dl24OiO
YnowAVGzwaGOL2SVmfMv+SM4WPo1yEKucFz5fWDqvlmObDgtxbul7IMx7Xq9
Hutxi95jcZH1rNgg/DePoOuQJVxTtgoo3QnCMIX0KOpbdnhoQyH8p++aT8VA
UJQUjXIi8f7B6PfHDMnKMm+tATShwhzhJc+Ls0wD7w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qBjONb9vhxPdV9N7kOIOjNqm9OhvLMennU2rusBtfy1tMbaJ5mJfqTyW4H1s
s+pCd6wFcOB+xkgucH7t0UvLPHJ3tsSp2gXzbTWNEHHgPE+AvPDSLXiVOBLW
m70QDb/CW2PgZQmIp0otBAmI7/rcOMagLFqveTIG3FyYTV2L4ZqFHTHEiAGF
bPkI0HTLATo7/zLOn9G9dAqhhyaAcXqJUBzqT+eglikDjDgZ9ug2AcM1/A2+
NWbRNd8KQqcFs9crA835n4W1lcGBLweT5jmYcZYR8n8yAU3ZZ1N7pJQcfo+3
7MuWoaK2dEMoutLYBb1DD/e9DxYM34ZxaHGvPoni7w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rh9plfV7c45bmpoP1SK8bGdu0VhO75QErbOdurUhZdnrv5ZfGCAk6cNnOM8l
lu9K3rcSaBYz2H4IuNOg8UOWKThoB4gmRN8SM+A92BYI1DdiFCDLYE7pDiw1
/Mf5Q8abKIkp28fPgm+PkC489C2SdhcUQqRVmud9elwrx3HY3NQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
dDorl+FjMXPjzy4nM4ALwpNusbkMx+qtjhuWjhqXR1cOc3hDN1lyExvEjvim
PKwlM6UkO7/HFG6yY0qvlGiaq5X8xSsnFphxi18rmzd4AEDYyVoma6c9s14e
fDqDPZylt5GjGsP9qPuPEPpCu7Z/mbzUrTFKefWQrM4v+m1jMbNDtDzVoNE4
gC7G1W6S07KyYilUEF0yOfmiKE9nXvD6TTOR/Bb/WKzcxTY43Lk/6xf1ahsm
X1YaQmn/g7+HrcXaRNru3/cuqUiiBW/FkDTZOLlF7tUdA+uDW1zJydnTU5se
02yQ6B4702UJhg/NemTlquTfOz3aUD2wPSaEo6JA/VHyiaYKyiOM6d/J4Nlm
cE35r6n0bLTzWMg1ZPZ1cHpBmrJPQMYlLKDOfJytP1nzmkV9s2nBstxbqZaP
bDmI0eBZJ+vSLCQ1EN2SQXbxPyvbhfxLIxIcV+dLI/bneAKpE4DxxPG5W1dN
5bHpPGPHNRMxuIc0NsW+369Z/nLgN3yd


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nwHDqxDnUERvm7bMUNRCtCRL3xnBdH4+IiiSDhiVTOSgQo0kopsBqCSRDwbE
e80znVj+KVuYojLPv/eCs1AQUiHvGHm+nD6EbrweBfeui8wj1tHKvchrfXM3
gctwrd4W5dMoTpPMN5OT5nWAcYH1Vym3bN0djO1tguEMSLZ4MkM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YZPbe96MdjFcggwE5LUosuQ85gvW/qQGabkNHoVYeWCMj5wkbDazHuiKN62m
ZxYfb9piA9ImINwXwvHr5X6pI7XwZ/TahC7qPJIIU/YOCzdeTf8jryxedI5C
qOU3QcUFSj1HGPqmhUn2M566htlpBbd3+YKHRlEB56ScG7hjVzo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 188432)
`pragma protect data_block
5DzC2Gk7J8uYXQj4ZHzAFQk+u19W0ylgqChwKsR91lRlbGUdQ0vSa+Zg3WBh
uBssOXVa2cT75AputNqRV2Cq7eCJ4Ca7WB2q7rmeavrRfFNA0qIxXE/YoEn6
VzVucTZam7UzFxPEaLokWyXhSKJ4lbfOpSusz+swPhQOAWRbRFuNZolo15VN
ySbSr1eiILkhx+4GchxhtLzHzTClg7rTdbp1eUSDyT3Z6gxFgvvumO/LhgZF
J5DvzMJOTQhhPv4oEoDyIxfUxfRtwXHd8VBK3Pp3v+dn2KNCKrj21PO37j6b
bga8DXXWXg2A3wqKK95qZh/zrPTA5uAoKktKCDAyRnchqlvbXcAfPHtCrrun
FaOH9L1/uZFOaODa/hK6SyExhB4bH46/NQ68VnL/EjD0AhmfxHmHuIjwD29G
BI58sZL/ygTxx7W/sWRgZvYwwyiRMrjdjLP4HqPOFytMaytfU6dG+KkWDgkG
m4P9G6KLVAYMvEPWbn5pxAtEHu5Pthpo8dZxnnkLONq2Hd3pLclRTpJw+Lqa
dsUcMINsZK8IDDQ2BYSuhkL2m1s+iY9sTemTSPMALekFXrJshVJ33ENmuGXk
amwlAFppeiSgj5pv5DxV6TxdTAwAjwcICga6wJAkxIDvouyGjQmJf4/uriSC
wVnNzJ8O37evrziAbhExaZgPMTj9gSu10uCszocetHImErWND23FUXV5ecBe
kggCE/kntsdVShIvMeNJQm6X/VJb5MXQkYIwOVEgMq14tw5pSBM/iWQK2isN
3rA5TEA8WTBVS/BIM2FQCxJvsuk6j8wJdAYA+7tzWuYevdDfrIx/ddgo96/u
315jErWg3bbJW1r5mFeyW1mJo3cpWsTUQN2K+Ka92hAgPA2p8TD93InQdvpW
fYFueh1EVgeYami4ZZbgFxgJrsZCo21icBp/n8XFfl5RWr5kTHnpMdAvfJbv
8fem7tqE1hvaUJjBC5yaC3LWgKtx5WqQ2B/7m1RYOVE5NQ+KGiIqp6yI+zF5
XHjiSiPw7IU3P1La52Bh3+lV53R1wWxiAHWGZhZJ0z61efF+GhLPide1MvY5
BcbcI+tCsadtBiFUuHOGRLZffol3H7ozXSsbkJhTaXPaXeuK8pFLAf44SZB6
K3ClX14gfAqxFxcmTLR5fLv6mHKz/ptKQ/lJeX97yPyVDFVpoT9VJYrNYAIB
k95o1U1Sr/2bwqupS7GjVKTXqGsmO4rjTOkbmrMrkckFO6MZeveyCW/oTgO2
4ym3ncCvSw7KVqgM6QpxRnnAzjeVi/D8znGxQXeV+K2LXr0PlhzhP311F4cR
AlEk4VU7OnD+UigkG63bvsm55i5kIMa2civXn8WbVh0hrRF6qIJCT3ohK9aA
rvXP+HdzcgrJiRVh0eL3MPiPHpjBGyoLXulfydrHXDad6jt8lxQrmRq1Eru1
KGjqnsY/eiFsz2sI/s0VqXK6j6zOBPzDobv2AyEW1OVMlVL3BCRmK8Gepdm/
WOTER78kPtadfv1ztTZnh9mG52dRxD7iEGA8pd4lFBuWAmbXfVnAk0E/WjRS
FjpExwNY6ytYq2wOwjNJFEhGaJLPncCNYIYnxJczB8THiy/kzXnT5plh1ERG
K/Ao2ia7n35yKZQQrE/mHUQkhqoTqVrhuNh153OFlT0gxHk/4rDkjfdqt9fc
70SzGmTOyD2yAyoFm8l8Ihqxdm4JvWLgE4BV8zbyR7tPIfrtKDg78RTlNBS1
X0JCvxIDr7Qt0mmMJWXI3zDIKawXJjetdrkeKHhmgtbOSCTwtSoPWbhKsMa7
K9ykxJSNSHWjLTkh5LFlGNppziglWgznB2UUywxMpZbQLT3+IHbRIjIWUv5c
u353ipsVQY18DpE+LCjVd7q2xXHMfN5Qca5skI1v9m4z40uEyyrIFHSlFo9V
YJO8w8znHJDLggWKWproW9s7vTMmRwaLTfEae8JaaYGooyPJHx07K9OLitKp
ySLriLHCvHcnaJie/MdeO/07oHUNbcUHNSuIoOt9Wm+YWHiYdxwmbp+WkqLg
QIvNxK+k9WU43QApGdTnxBfiYjK1lQAuox692CLOXFx976PU7tqqMH9Tg6Ga
7hqDz3v88EU6UxaeSvZulQNVbwfgJN6GueX4nti5ndogPxrvqGNQEdgol8Vq
IMz3ub0Y1LnswQEqB4bKF8p2zqtcOE8WttrkWoEMFZVpr279sxvTlUUF5nsi
VIaetMdDjI254ub445gyVO/P9Fbt9BD4BefGgDyAv01nQ0bvz+vUWVneczE3
OEQeADXsuHXGApAdHkmF+9p4Czsl3Ug5V+ua3+CjAfSNv2as3qZrOgnwQXfs
b+weogtu5zJZe/OQivC/anZU7B4SMn3f0HgWvqiTzXyH+hf5qxVgTY8FZqha
1wHGJVMD9kJQwmI4rug/dn+pq0fKvT74H+kTjL0zyWYvscBRvPl6bFs+qpX/
Z6DsBaAbalMMQco32VQHXm/0XSuJw8+d8AO+iXzv79PBa0cfcF0xZTAxenHd
cV/Fv+xO/p40gYXvSDPnMw3nUKP8+v3NwHUSx6S0NpboHU05e1TyMsYLGrEJ
+AMD+w/ZWcd77fibJcSZntDYXW9qKy9nLVk6qrZ/ZNQtPNur18+3G5UL+E10
ntkYE4EGlxu2VJE+lRwcKHbfuVHjEFQpstvzf/HqfZbHmM5N5nKGv2kP/RG+
A/DxRS5p74v5+wqCjqDAcgLEn3jQfugkfr9cRW42O4BvCL9GUz9U7aZ/k1s6
7mNrMsnlYIudUJOfKxnQQeNn2au9z1G+B3ET6X1gCYo600vZpJuOg3AMvvjX
/8l+jrNltgmHat2ILxhITR2dt5M0OzbliSbc9MRhdwjwk6tXI4S3xLO8hTja
zwe6DPPTj6zkkJr6WVWrjpOlg4hoykNPx66i93c6VfsUoxCrMkZ2Ns7mtKe6
fSOMws5R6vPUgp7FizrDbuWZY8D07sNcpEpbPHw5ElbjTXR56BlkSyJNP2DV
HaTca8EeSm5TPSlz2pOWF2r8Fa50AZ8C6RsJZbv2StV6XIRuOI4CWx8mP9qU
Lmaboz3XLERIUYvHRX15OAL22uNDZw8tWeZm45nser0k2uv4MWiCUD0s2FHu
PL3dge5kc92EWUMtzp7gynu9JHRRYZPvaiWuDxbGJGIEREWT7N3zXbwkpubH
htyFWhtwNyPIRIXd0YyCrlxJZcFurRL4/cPj74nl6EVObcg6asjJGBKL+pZN
1I2lM7XygAS174dy8Oa1L3aDmMpk0TZAzbG+sWl2nWq3JguYDSrEp5QOt3eI
D1bUklOR2SGPzAcnru/0WOsDF5TmaZsuZDKUdKRaCQvod1veyyFtocG1wT3d
BvfSP6LQ+MdgJDlOm41t7Ei4UL+fAnYZAg60yy/CQVW6ixfGVIq9254BlaU3
50bGFxhgY65aFIkBHrHbGwVPyQXoMZoBqDxS6F2bctkSI4LEynlqtsDtFcZT
RG1I2uiImUYIaowNphqIXO8b7fFu3sQf2dVTNhhI2SmCBseVpeJi+JfePhG0
56LSQ3iSrZzQuqh1LvUGxVacRGJEBWg1aw+hA8r56F2xK7Xk4Xf3V9LggYpJ
0yZE4RE0uFkpFYLke1lVxxZFbxyh//aGnEweGvOdcp3WTIgqTg8zNLSlcmM5
p7sKsqCpgGyAQWQ7scMePMAnROXmlyniT4Z8wOjbAeG7vYzVaU5yF286zhnc
1rqUYi60/x42hmBuDYhsYLlbQDFSg4Y+/7MMVs3/nzZdS/MhCzBQEjvLNyOO
zzDuG+4WQPw6siv7O64gYGUbmatj7dE0k7Yoy5b5KMjZ1Jc5BGGFf4DaVimc
o+I3PgD05irYv2Y2FfTVD0waGeml9vui0a0c+DIpL/CnqyljdmvVK3mK9FtN
6KMAjMapHTvc7748jwXIkpqWX/GWCZSnOWb+dfMnsHpmMl3sxQjmG+ENFGy0
ARe2yh84xPshE6BjH+/b12fcwok38Ls/hwvYAUOjW4mM5H1DOxYjjSGrg7+1
cRQIPNaitkw8yoC5ElPnxIMpidFIUkaYpzqdTZvAejFwEbpUlKSb5CH6K9/9
IEEVL6DdcLPzuXfiIOOh9p/rKtyi3w4k3LTWge5fJd/XZGMSlNQHJFI58tGR
WSr4QeCFOPsu2xWt42koZqksPSJDz+gKBiuqSnCXd0qWfs77LHVfJlkDsE/2
kqvKW7NmEAVIgMzHGfuJI4CoaNg3Q8qbbCGkYzr33sQro4BR/uhTp7zGFlIn
Y8NrURyZi6LUThYOZhU+k4jih4SHWFdBxYxr5OyLX9DVYAlTZpSwtn6f3NXX
w+b7Xg6XxryUB93ILNyyT6jXlZfbzeR0MSv909gfxlA/Y5lfEMg00+SJcJog
vu9Tjp5nFQDImT0wMTm+A+9cEtW7M9OJA7f82MFeAtCaFZe8ZHwyDNpTDQfn
WqeIN6QkiatjxCsAC5to7T5120yJzhiS4X6waicQXE85Tb5lOQPwvg5zxSjy
altzNtIdfRSUrVOuixfWH6KvC1LU3n4AEev8joNWhZmPNVSkRbnbPASKwFMo
O0Mlfo8ExlgDKtdgjNdjU13vJZwRak/tWStO3buBHiiCTBxuzcvufffAt1GN
78z01qy9fcnf2ZcIuEgMryq5CLVU4ZVtcug+vcRWW6Ihin4hA+W5hcDs1ECQ
w7/8y+37oSfB2UTJBYUfrOMu0bGltgBLaCN0EIF79YxHAPevwjCKhr5y5OlP
9XmEFEqOiON48fjMYRW3w3mnt55Wq7kPE7375A5B9YRmZGYx9KCYAsGKDhgB
SLHLqFS/NlvL1cKtIMCPOea5nHzPWH3v7Bm6cuI879VGnYiuSp9VaJ5s6oGy
mNPF3FRiCx8n6K9zTTaqLx85WWEJns+rfQS327GK4KJqxV9AWU9eEJCPsaho
SfFOFStKwU5YvUbd5ueyl/DsGtMF84tcK7q1+LzzGe42lJtxmvQbWvWCSzts
XxXzGP+y2D8vgsVkRzKzU+qsECOymPVJSUCdLiA2at3KDLN0DVAjXVq5Fhj0
VL+ilCkvKf7nfQlsyvykYd9n+byK57V34U6auRYB3bR9KeuzLjWuW9hwxoPq
QoWu1qKXzzRIyaTB0L9X3Rw8OOtyuN6+bXoZeVRH5pIdwBmagnY+rvJfaTOE
a5ouyq63Dr20EzCI+JYJSppRaInnO8xPMSt1dRo0jtnyrfxaMlLD9DskZXa+
6fpZLNSD11JXD09fxcNiBNMtjIrqGCmMidL22XY/irYqkCbmM8Fh3XB+Tw8q
IV438E666xkOB9/o4TvQDZsYy9cyQrkFUDYytJvjb8cA6uCDRNw5F2J1rIrE
pi4AHbGcjyik8ASyso05ET3rijC5wpTW1eGPon27eXKmqxEyFsVLQBQKXTpu
NsZ5Jh6AWeowIK4zC4JRIJKn69GqSxGQcmqRYAmYZTRU6Ut6aN42Vmtijr9D
q3vpbYAXkH7hSzavj47KrQlLeY58DdU/XiJSIncGIm+5EzpRfYLUcsZnlnar
5yiv8p4vO3/8TzHKy6I1BjljIHnrFfsiC6UA/2pWsEOPsnAirRUKYhPHKgtC
WEk19evkGAyzjYa6zNfWxWZE8fDYorTcZzauW4mAJ6H41XzGK6dML77ItyJT
ksjTsjElVRvbAIC6crCxMq63J3mL9qtJg8Es9i//lg36YGxDyQBNPs5YBf+4
pzzRxZlPzTXrQRscrVGTrXb7Jso9mvHoo5I7gSlDhlikfNY9MBJJjiR4Ddez
qxWYJxDoLyZOaPEPBX0W789jkiwaYnk32rlHjnIXKzH/020LR94JItcokwwK
LqALuzkkGk1Ya8glIFFKiOFzMPO4D4vUZgyH2WneAUNfbgW3RVczC2bPY1VW
Ckzs6sCLLXaxxIcxcw8FVdGcuiKaeri/sm9ZOClYaVbJGK7zk16bVnw4ErtR
L0l31OQFcjFiKcuZQhhx8PDsI7R2FO2soFElOfR1jhgZh9tkBbGYE7qnktZt
rmt8IuA/sRvdGveSWjgO6ul22BsWZKOo3r7a462sxDVotS3T5BPF9dxR1c1C
Q9+MSnU8o3k0s9hGm5sBjLubT5xw4bC6Hchvv6gfy7/8Hki8jXHvsGEsef4l
Vgo2CidBdz/he+16y23dtzwGdcAWB/caJQH0pZsuMDVBK1HC7FRvU95S4Ggt
47PlyqWFo9AwNgm6n3bL2vG8awcpHIHoZMfo6uy7zFQ9UuhGA1zetE04xGyL
2YUYuIglDkMiiM0wYPROFxYEn7U1fy3eqJsun9gBrKiOBj3oY9xS4oz5c50n
hmc3Cc0DImGFG3moeL1XKj0sNH6GhcmyEDhGVKHGq4QNbKMIUabwMIptwX5f
RAZdueGDVChBONpM8IAHoSekkFYHMEhGMmLyI/buwX1zk8ISzqj541nz0rJX
R6/7m9lPWEjiav9f3nbT9z14kleZe32lx2bLLPsUs5StQY2tlwLiFkFe24N4
OnctgDrmrrTzQUZ0T/jMRixDFeGev8f3y/ostyr7rnmB/gNyNZoKO1ojGo/k
5L/Q/dWN/xrL1qCobnZuXNeSVea9/4c+fM5yXlKtfp4j7tLyDYs3IUNiXhKx
Zk2qAr/+jFJzWNEn7F4oBKNo/p4xDSiNE9GcBJpZ7TRpSXPtLVDmRqvCnTnx
MuLV0FJR8uQNLsTp+JMauy6H1i19FIH+7Q7fyHu9mSZebI4YOEY/sbLjOt7d
pQ1LeJdrK5P2TMQWBbTR95rEG9ay1Mo1Otws+Xt+A6YYHW2QG7WHbWYaMBAK
JVOlMtyxvN0lDVxphnd8bNsd+a0WLUaltc/EgT5BFd01O6G2lFVrkebm6dnp
7AWz+Dqv7osrWu3GPhGg0tr8ShNFX1HuwhPWPR6aTB/gvg/IJ0AW8B/Ss6x/
wKw1+UsQUU7SWIyESKJVRL6JHgHg3L5MOwDdSTqpb0wfqT0/ulb5pBBbMmiZ
pf5aWipNPM1AZeWJz2lztAhN5EFQTHJ4+CA1zgVscKOkEFljhDY0//Vd4HiO
2rtNI/O4AjMBS2bYaWgM9AlVtguHGAcpjltzhy9KJLL9Q/XX24NuPwAREJOX
rONW3xEMw45A5r2p55OJjcuDRMukRiFHoHpnU3FZMyf3HfdqI/yAO8T4BDpQ
v9HQnnUGTp7jIEnm66iIRfBsk+pNGHllRi4o7xfmSpMK9ejqGmZUA3qnqD2X
2hhis3OiQA8sIlKoUjUzX6xGewXMyiNc3YWYcD4s+MjIrsV5d504e4fCCPBZ
U6KxaFS4+XFkV7+uOhd8e0k55hgvmL9YjVx/O8kZUevhUzZwnVtSCfjTyMHK
/I9hWe9mvzgf2JrH+yFO23RbndK1DzswmwLgMjxCW8LrQOt1KgsPsy/3M2Ze
H4/z7+DdI1EG+oiLCtQInM5x+ooqW1BC8Ee3wO917UaSIcRS7VhKU/66LKZ8
rnObzF6/hHteTJrZW0sPNDxXNCM0WwdCNFWw8hapGH2EluxoMDN1NQPZDMYV
grMWLwOqDJIaIoKhx4J1hLPINgzCPB9jXmI1y92lQnxCd16YcQ/RGP6yH4+y
EycZ2lHfZixeNPMu4fo/DGwTJ73xzqDFeNWsKMy+ASpcYb2O6+USGk3ZHuHp
v3JjOWaZd/UxGsOzbkk3DPnSfUjW/w94lMJGYes0x5WAmOeWlyvu71KQL7UP
n30glWKCXy2VMUjdL6jn0aW4EwBEJXpzIokFhBQKu3OAGLST9jt4QmnazhwO
0IrQijIKPXOSGpDy7VB0qIf5JGfUVwbPLplfuBYTUTnBwtssqlytL1DMJiW4
Y6IQmnPlXOQN3Uyb3jL4vQy/Fn/DIsvAVJJQPt/UIuKL2rNYiOJcoLdWJ8VR
G9X93Ta7Yeip6RLNfqhei3LMsTmrPc54M9Y0kxnBIUpcHTsSwz5faBMWgEMK
7ImX9NH/yPpglpDZseORhO2CmBv5SRBGx5vCxioM39SGey3oAk1MvEsS2qrk
QtdayDww6fHTQ6flTTmKawK7n47rZv52m1EOAXOud16dL4Mj1CPqK63HC4Ov
/2DpBaHh/tnaWTrGh/QzUDlcD4y0G70TJ3nzZdZs1fR2LMtQGvB4XvDrAHnM
npRZqQaOvX9KqL/6KA7nPPYs1ZF+lffo9Zg82eZH3Hr9ZNd58EXv/B3GWWkL
OnjPuhVL3VeZG/uUfi+46YRadG8fWJbRHMAhtTwXRsAKKOK1yOIsijjbSHKm
AWnX7FW+zTIPTvDDtqUQ4MxWrzD60e1YRQR1E1++uYxGkUzGM4hCjqYTkw/X
JsQWhzNZebqiZ5665dq/pJUvzK+T07D2CILl9L0lDa1OeYanl6VcOjwsqg9t
v1QZFGqaUJ6Hov8G2EfGYhUICNVC49nDz8S2Zk//JBcT1VXpwBfAuD/xx1lm
tnpLdZlmXhs70BpX6himE6WXXMa+2MIDOLJvLj0QYVB0fbONeV/U023jOPrc
GlETWKTpcgaoGPxunwx5M/SUjcB9A3bSXNJdIEkQtISsdtN3rOL2mapNHonX
5sBFeB3WUH+Vsl+j6nL8XkpSUk05Rw+pNDofyHdZJoA2GzswSJASZ6NMidlf
vBoiBrePCMsgP5ZbSGhwj02r3e2wCyawbugsXBd9dx7z9zZajMP7OSzptH6W
kI6IBVXNw93bquWS1SknQswDtS8mnv65hXGuTq1HAg1x+3Mvtp8wmaw0tWN2
hwCwjoTsMCqcqXXHqergfBl8yRsneU1Ukz1FYVz7BjRK7ACxxmgHw+zVIcPr
tQ0WTo+zkHVjL+DI2vA9qOa1w9Po2fIN41OAcxAy9nLnX1dRMFbXnN9rlVd5
WU4MxDYzjDoHXFE7SVATPSmA/8J3wSiGse7nvFzDk9xHwBMpV1L2BvUbDqmZ
YgspwMRPo8B7YByiVkpYzjE23qbgautBoLqZJLZumcTAG1OT86ncCqod09Uv
H2CcsnO+9JBrXvs4hOjnqF97r6CQepcEosT7Yv0/nR4lAzh6LknRBhjLsvUd
O21nTyVw9oWCzVq7ccuYC0XloGtxeA8wvR8z3D7BuBUzYHTo4YdUshWMhRpG
HPpsNcFZxzZTa01txLJI/YX6fzOhHY4pj32r1RreFBo+nNZTwwHg14SoCxiZ
rzepfaRQhRWEq/g0JrsNQwkkWhhI6qLg++LN3MRaavtvNVAvVrS7O7CfQPRI
RWzowBqgTM1ALKiAAo8Dy8XaW3ZIDv4KP8yXn6J5TZF4KRML4pFKqYv1gKnJ
h6blVc3LH8dvAqisG+ZkHh1h8Jnuk1I05gyYE9MerrxWrmXVmDVvAn3LjGnu
JeqR4LFM0p5eth2TSxDk5APsRlt8Yj0Mhp90tvxj9q1V9flAl2btOLiPZUOl
RepjtQJJ8BnBG4FuejaCw+2sRBXLyZzte1jbU5+ZIWSqWg0ofDqDp5IDzT69
ryW/sXzZ4/RiInhLJOeLvEpL0TcY8oMomomvpGn1E7F87UAaXhOtcU3BWqaF
w04bWoXklHJ68CBjFgfOjCiHY9jPH3h807tdPxyp6T1ttju4A+hjskSiK3EX
Nbm5cTv54jngRNZ/dIxbk/SC+IcDivd1nar4MQgvRVvF+jNnYf8P7UhW3nDG
eX1urGKO2HWk2EtnskmX9XDkUY1RThs7BMEVVHJueR0hLlTNOZq1pusQ+YqV
FxTrI7Cpdyauzd7S2t6FguJkxvrgM6xmUddgPQC14we3AZhigX7bY2v6Xhl1
loR1bZLFf/ISp/985xt2Gr9HZ6Wb3MlaSElJKE7K/4aImxx5xYB+ry7uasnx
Dj5yyoojM9nrMPiPcZAcfH9o66wxWsaB4ANTs6aEv2dEf6K1ZJc9gWBJsaqo
vnHbtr5KIpLQVHCA1S7Itawyzp6GOfg18ymPk+7jA31j3oSMKtMFYk0Skcq6
/kmW+PSAi3V9+u/rzfuSunqIeadZVGZ8Zyl8d183rPGNFOwT6mgEq1aN2B77
1AL0GGNi/6viOqSqg/PIUegq6DJioRbRlj7P5wa85Iyx6fivriMCdnDfCXXE
hKyfXSMRUt5V1J9aYOIcf09dKUQoPjGWZEEB72sqQ8pikyPUYByMSY1vcUAp
0KEXa2JRW6MQA5dylZCiPw4hf8/9HVl3FnkXI3OlkTT4dVenPOI9IPlaEo8L
221zEUtAYBdsXRKANhVUWV1jzyvMp0QSm8By6ZB7LLbpGR9bLrxq4mLmNuz0
fvatqUg0qcDXVMBbBwvfgwO6qLAIvNymVcqQXbZuhkhztK2IyzOihNFlD315
sPV9EmuQ2wTHmjTs4FlQISC8Fz3Zdj051SgoHocnpMhc5818HScwGaOuH5C0
1ibdZXjnUQjxzCEbeYGN7fsZMGrzeymSx/U1ppsgyR7YcF8+MlPzn606D7Ax
evzxH5QKg8DPlcUNURV4hkU5qfVC9jxgGcCAzwefpCoCQuM81HnBgCY6qPJm
YMg56HqGPPhi0PBVrTYw/Md5UGBf+jcIwOfTlAQoNzB3ppWHU92nRxHBH6Ky
xw/9XAl0MoGPRi5vc3nP38tvUGQA2ziaes90LyJOuuRtD1m3/LuSsuk9nP34
45EEgL3X17iKSiC7Nv0XPh7YWHEEqYHC/3KE8wvEnaF6pUa6IZaBgW5VDUL+
LAL+BLFHyFBKOSmi4LQpD1Hs9FUxjs6K68g8xYy2fDl9Rxlr6teHA5ainYws
DPz5mp+eKoXfgB84SkJuKUpIn/bIojITMbXPgd1xv/dW5Ii7OWJeQXsGn+4L
7BSFHpb9PsQ7NjBhi+w/Ctp1WGn7XM/HB8cpPI/mYWs7yS9Gudyw97Vu/I68
9hBrz/u0wAPJ3RMQVE+rcVBUDLVwMHxK9Vz16+oYPUIxaRCOUrDmklqeuqN+
a/Oktkj/ptdUXBCBkkLP0ChWgxMpfjCbuAfMXXTKnz0CL+r2N7lBl9QqNyER
uUR0LiNstI39PRtF9x8Lfs/C4L4wNg28gJeRBQjiZoj9UbVuMn+VI2TC1Tgn
5Ks6xdUDrr+x7y59AQWIpl6H7k16PawNd7MD724DDo01nej8VXu68NWji50c
AYHEe9RioyifiJOtIe7tCL/ZDvA2VsGWkaYMgcjzSxRbax5Nr7b3HqoQMO5W
5hqAiKGvjMkO2XlM0GmAJ4puebPVEq76h3kWiziluDKNnheq+K/UY9wDA/Mm
Ubw+ktGzCbD480dTe2pRPqnqtjk/gDZTx7I44RXqn0jixriDqHsb3DgCb27M
7LRVNLb/PESI1muvUzwKlWBpU+EDgq5JsbWs1a8kxxlUTnGicORuW1Dvvi0F
J4DuHd7DyRrmNnCbUU2j3QIGJ+EbAsRuavxhDbchC7TcLD0t0X3d4x4MNLVe
xr7RDso9d+7vgA0JXoH+jcUNHBzlHo3scakIc3TLKF1x7+aZP1+6WWzuq0Gb
eFJOgg43AeXKqc9CCgFuN40UD02LpobR/ZUZZJ5SHvGQV7x7SoWc1uixH/Te
UhWLoVDRrBrBYSuizvt8O+r5+BwekCGiKAM4QyyEYePllr17O/MI/7hBzYo4
LZhZoamaYrFlp/CYdaOQVoILyDPebAkwbkdhgf4iUi9oDl/CMVSbDC+P92tQ
BtDASaMhL8dTusAIcJFazG7i9OvWKPMXlvqGCNA6HmJZcKMANITejGd4irb8
7+ouHpIoQsgvlPXnBk2iZI0204JJe7Bn5LjXtY+2Q0B1aQ6A4ee6wkVgFFHV
fLpxGN9+2a+N6EW/GcxWcBKOERlM/VcMR1hHSgOZrseXNtWpFcYpqzMj4wWc
KxLlrxkRAYmIdzZbOAYK2BcgjifDYm5+utCb90Pl3e4dIGh55ufPksiEC0DK
ltPc3pJFS1m47QjPZcHw9I3oEsR0rRbodIrWn6WidKxwMXnl6OiQWONrYdkk
56ySR1MgLpuSRjYurG3hVFz7wthFqC6NGR6lLSLnnCW2g17Pb6QUuk7fsJXK
jgh8ytkzAO/tlvQjpNA71HdQre4Ka5s4wt+bno5i4nwaeUqSs43JL0esEoFM
VAlQjvlc4y+9ZrO7Novl0Qvq/ITk05w4/H8cOIG1b8Xg8eqwoA805tR4vkPe
HdHkNDDfipmZPqNs9kmJ9ECzuFc5km6x1iSZvENYFcjcm3tfU1RPDajy3txn
WLcqKsI+WZeCG05H4MkXGK9Gp9WMzm9nORB3BayVsUvLD1UTs7x0sFin/aZu
M9xIwCO/5eLd/NpTZHg0x9ilrVvK49FdhUYk4shEYocirLKUo1qUkQRztEmQ
gvmehG0OXzD8NFYExgKWbI5OHiPlQBjGmMTuaOTBtmxXFnlQJy3CM11Fqo2+
HK5g7JkBMWv8lBEJu0r82eNnu/F9lMrO94B9Q6RlkHz10S2RG/sk+JdiHMA7
+1436+TyPAD5wXCMo/9jgZAA80JJgHTQMg8WgkmcK0jWc6cjzVqAB5JijqoV
i4HUYQU4dwAcAV4dUkPocvf6tOQSdiBWLURQkHPaII2QaDkG740Um1J8p6qV
SVLqaGjccwFEeiOpDMLlKQ9J0aPVQZb8VbdPmPJqK7kWVbJuxu7MP+AW16le
sg2EtCLS67tRMc97L9lwHEbQCSD9/XiZhLDkaQT2pEpE/WZq9MPkVa7u56Qp
rb7Pc6g+6o62BRlIx6TA79cqwayECjVVKRtW+GVZWaPHY5m9CkNsG8S2eU0d
DOfx3Emtvw2oIEVq9gB369CI3signzEnsnU7+6qbypFMg+YuRzm/+Nt1f+Ig
gLUJ7c5wKffBM1+Ndnxz7gwnfCEZUAwBh1SPnf7BGz+15Z0/MrPGCaIEctUT
nDzfTqOt/lf5Q9+QKrJu80/qRu22BxHUHzKXbOsu0Kt1uysEbj3qHnS3INJ1
NmaMIBWBQwjtu3t+IYPXBSmboXv43DPdOxuwxWt5jitKr3gDJVhDm4QYO3ZB
BllcPEQozvfexq75ttxW0MKdXVBiOBkG9HjngSQM8LIyUGbHFjC7sjhd2CHH
pU65RYy12TB0Av+smkIIT/ebCHhcIzQyauHO9lWcNJd1i2X1V2tA+w4WBBsx
xSdkg4mDWdWfVt3bk0ycfWt8exHBufq8xT5WU5P14fFsbfKCjqPYcehl6O75
4vBWCfRjQ0dWyRuvy7JZdblEQUqoD/EbCqFXjZtCRHE2w1EhFA9YLz/YP4SP
wZqhozByUuky9f7vz85dwBGWzEJuEp8zqainsIFJVwaZnBfwWaA+V05ItXI2
bj7CWHG+46wJDYWacunQgS/R5jqpqOdobD3sRGcqDSv1nZvqXJYbyl1UN0Tv
EP94I1TDgdNN9zDmGeridghZVeVAG94m7v66q+jgt58RojkqanWKKVMEjkOy
e87K6yQfVp+VdfS+6rx2H5IKufEyHDVVLEy7G9idWYVdZp9wDq7PrmTu2LfQ
2qd1wksyMgz9uwhLokMwfyUA9X4EhbTIHoxvMbLbQfQBPyDdpdPDTUuWi31V
y2KV37Sy2e2UAKRt3SlEb/EZ+9EvSmfC5gpJ/RDRFIWKH3A1xmZRI5FOZwcZ
ZVTQZu0XvhslG93l1+Da28j/+NeVN2u5aHNE6M457qSjidBbjzwu+Uw79KGD
nED4g8ZF4a2UXSqWSd5cdNyCtZrhn5nfqpO2+IKW/kBrsK4hIj+uJnwTQv+K
bgjYLYqsWySDcP/ZM4j+Goc9OsKwVjs1/chthiE4zHFPIeuvbFWlbv5Bcjar
Q0sC+YGeFpKTXdU+YUH/BSckGBzBbISsffXRmW6dAYpiI4f9/aXOuNW+FksC
4tVhTT2/2LR6XnE4/jxTYh40C5VnUyE7rBTU2Lowz1xCVYtArFsC6W/Xjaq5
WWM2tkxpNkPel+iJfV4Er7aCBkw8jilRCui5HjMtL5dEBLTi0SIG0+U0bjf+
+Pg4sKdPXsYszOgJN4r1mJiPkhr1BB9vHvWokTF03E1PJWhvC1lgw61Pt27y
26jsacTip+L0k77KmuZm50jCsf2zWE4IMjtRAhnE90LC3G8LVp028vczCSZB
szGQsSx995NvdxmOp11C82EOCzuDCjt0hR5t9tTES/j43SHLx2Byh6DmqF5V
4cfREkqpcPh3DvHBKv6nlhBj0N0K1o4S5TSbj2K7vgQMd/Bx2+QtVKiTk7M/
VaOdhDyfOzEVvUcVUD65EkxJJXAkasMIjtEzOrkHWicHtWZrzMlvC0b8yBKQ
YE5jOJ61IINdlyIl0B0asM9YoQLRRnXGkC0zeMcu2iGnW6Ern+gzJKF+FGQy
ys2KsU5bWAt+iinID33/CF/9tX+7oWa1qRVQtAZ4/UdLxNwrTvIg9JE/SkRs
VXRlcuadGiZN3CR4tCaNWuFXS7A92QUDPn4qGF4jS/3EjG3C3/18ZPqYdfU1
j5ndkf850RYmNbQnHY6b673wSHGxFPln3OrOqiqhOyBhBwxC7f59zkxMh0eK
MvmXRGRqiqtFCYwZahYKztLL3xi5ilxgQmmrzixJ950uvwl9LBcVZY8sjGL1
X4l0uY8ndkOjlfpIWS7SZUj+wP3DDpbqsKLA7dK1+0qMaGIRL74ovkI+OrUd
5yuKvjYgceKm10ZVZbblZN4AzQkS67H4lRo4BV9e6A0iQoUJmQmkIoP3Tqvy
AQ5WuISXBjvNv6Ubg+dFuFm+TlN2/AJmE+x+gMp7TTkzncwvC/8flYy6uc7D
awYtDtyPSoFZWJFR77+gfhl7zoaV+eMRTRcjmH5PsxI8hDMb7yW+juIn4ead
BDoxpK5uCmzTAENNxim1vJxNdfNITNJZRtIwrdmDGm/WUmd6P1NguX95KxUp
WSEmwRdCqDwIEtlEj0G2vovhnH0gvEE1YiW+eP00ye5WkVs2fhdYk9Vbx68W
LyjQnGplSNXFR1Z1RCIAjJ679MGc+0cdswM/1HrHzANr3w2w+iwHbvI1BnhG
tNM111ATJQMni+qv/RAaCrEnCoL2KtZ+mG9sNn2lO2I2v++4eibuE0/p7/jV
Q96LKSLOsWMX0PwmJbFI7tCyS9OOhdwq2fJ0J5oxXdIlfB7CAO3zc4xPoZm8
W9s4L6TuqalCfwrHHQMAOcjc2Xl5saxQb3TlvR3JqzLMjzsWKHD7o/WOPNs/
lTOZ4T6Ahcm0Z3HfwvYsJIB+tqVs2ahn81oZCEADTpgCUlCmdlT4MXh9n6jl
hgz3vwPYIOdEGRctJvIhpNUkQ6eoO/+Z5re/WhpuWhKT9uscKxryJSlN0qdT
rHJYumaNb9TATQEKOwTSsmFpTpdcBqYsEMfyjO0SvjuQyqT729CPk4dwAEt1
BOo0GV1Dn6ybfhdIfJ2ruPbV4/Y0LQcEl3e6GKIHjI74IXU0dbv71XEMSFpg
O+hw82WlBXyTQjnAoGUhBx7kw6idBwUSrBh7Tl7qV8qxfog2HUEPRBqL7NXP
2cIWR4GNQPfA92Z1AbsXjwpnmBpDgue+wqRT665FVusRk8CWRgVwPv+j4sTE
R9ijpbchQMkhtStFX42yt3LKj3iJnHHyAelEcdKp6fiFrgb9bc3lgxr9fAVw
vE18sJ61jRdbLSD/npVGg1A5rv37Mye9BKC9E/Lt/lxdmyWrHP1w2AoGwS5t
77pLKy+PHzoJaoUElMpYlek6NYt3VhtV+MzT0IvQe8kq9/nHgltEgRgZ6WGQ
Bx9+Hk3jiiq5dOxCpbmfCaRkI4HyaJVlv+NMJ5WbvFZCBl3qk66rwmLlD09q
XzvwkhR0CihYvX1dPZaieWf4byqb1EeBS94TbPRy8BVumd8Y9W2QTTQFYQbd
8B1tq6V2aW+lTK7wCBdgILnYfRuk6L4qv6h7WDttfsIKrtN1k5Za8Un4/R8G
QS+qfAoYkUBiHulfz2444eaUA0OheQRCM49QKX94Y5mMzuTE2xgJQmn43X48
+TDm+NC6nk/bQXoA8jTfNilVFRFccpHbITXe83EGFqlFagKII2QsoKuH/PeE
DsIMwpvC/IBn45NX917FSDsEnj7A4BMWN6fj+apLjMBQdVdC/dhIXfZAnptR
Ce87OzBItdms0AWh4r4cuKmd0z01xzxmu/0xdCH7Wjc1RE3Wk9v9UtA5favb
kCEcLJV3+nz32MnL49Of8InT50Tg8hcZBurFeIvKu8Xx8POkUcWxs3URtTLM
Wqpcnu4qnl8oMJ3udebgV06qrICg7qT/tvqmll6MKTm49PQ7+0/O5Stz+2jC
5o0aBGF3PQhLzAWenbrHTtPDv1XH7JEazwq1icdk/Obqb4WeIzG/zWZ1680c
79S1takO0i/5H09xOrw0OtTfMK+A9p00hEkpccRsIw/0UX5Xrf4xPFECu9zc
xS0OWbScuSvhCcExux75YRW63btsTl6Daj4OLor/a4C5Jo9ulMVF7zG16HnB
WSJDcUmk7DZUtsTULXkx3Wl4ePNDV/QeN0bZ0+C42/R7+1hQuYL8ulCSnmJY
Io1P0QiYlSmwpyiKeYvyPpNWz7rOxzUOGmsWj4HvszxEJWdHV3fEg7j1BsN6
/F6Z0V9dUkbEjkPBnAtMAmw3ogWXDDuvrZvXFqIGVnykM47wPuDCzdDt2Ra9
1/C7n06XPadClcPqw+lg8hwqEF7NRQaIgBE30WuOYFW5Sg9wduxZkjzWK2Gm
5f735GF5vz6TBzmsqL6HmBBFx2aAlIi8piMLHXmaMmKiGsecTG/BiIhOOxEN
vFf/wbNDI0BGFyBN0K5WEe1eQXbL8ZnGR6LOcSmxDKAYTeTjLMIuD1FLAswk
6ZSHcDOSAuVICPthBK7q6Z1sMN+jbJ1CoI9T0K0K+fy8FtgFqx+bZbuwViGF
hU4Z/zcRezaAI1MXopUoE/dxV7PLR/0BrwvAdfMnLaVtem90yNvLqoLil4Ae
VVwDehlpDZwVKzq8tiyYEgOuTZMo/zYx7YqCSZP42G+T+aCK+J4jTecgSpCY
Lq0TPbkU+WPzq/9J3hmQBERW2ZIP/AbA0awbE+Knl15O4dQ2U+l2Id9kfCTj
weI9bvZmNS7ub8cvnolysDCFLDg4NC3hGnQG10YqW2Gk6R5fM9JVzwpPqQyl
1cOGP5Z3QONRN4JKlNEyXv9MzAg8A0Xu/PJSGr7o752cbWhV65O4ikPqx+vv
GVqHzOnX3Yk+MpL8g5gZDOWnBIIhcliiekL1PCZ0zprISxCECWuqM12Xgvgx
EH5+bQr7iYcuPaldGwR3IxJtyxpI3UmubGz8sEkO+aJXnFOit9brDwG4dnkw
Vdz2izpZII2tO219rSV5GUwvjBrVccxkZnr0MfOZ1eijgvnGBhUIMJqCd5/c
buwSkdn8X/KFLdd/OBn0FzHDaW7BBVrXUS1c9vJ9JgYOfc3cnvBAoH1ROzxN
rimMqTQbdEbwQKtts+dx67ulHu3TdcvflvWOydgRIcWFxArtzI4YR7YY4/Qk
KUGsI7sKrFvrsdLeVaAA44MKdg4ndWaNNyKNsYS+aFeJzHxF3OH7dNHo1bv9
NGnFWtYWxNP3hbYqfLYhZjUoqSiSE/Obm5TxcLMHMxL4D2u1F2vcUU1ZaUM+
itI0K0CynrsE5Vy9APbRXuStFIJdU75zFyU7AosgH3ceUOwmX2DVXRDMeMeR
rBfernappyKX9UoBP2T+PfXmKT4ZrgY+AdHzLe1AZ/YVDRF85YVFZEWW6PmI
zF+/3mfn79qLKL/4ONMP//by28R+eCpIH3DCQ1jlbz5505K7Mj6WE9SjApdX
6A8fLbh2i42zzdYI3n2xe1xWts9o5pn999xJdKzlcWEQKGe5mSq+EAVs4Pov
pqDbL35IWFhYx5vruOyXJERTyav15kN2eZ7A4L9uHGGhy8UF5mBrIAv2yr90
KTREqmV+N2PRSZr7sqWm86JGToZVjQ74jTDGud5G7KjVfOA6W1Nsn7tSQyiQ
yEikysyKSFy0M57fwxlYi6+CCSYmOXbvzEv01fGSve4y5p0nSMm+cM3AkcR/
9QAhyxter9tyPtzTgulTm08ROrs6jluJssCBYVKpjC8aFrjuifXlZfjsaQMR
7MwxAdLydu5ohJRRkc6Q0SBdPU3ZpTt+78UydaLeBSZCYKP/5Z1bMq1/w7Tn
71Dixn9vaWoOP8jjUm8aRVIsQL9AybXi8P4l9/ysYa5uyAW4xY6Ge+/RP1TH
qnABZcgiuWiseOoKmuTU6DLcMvYrntbBp5uVROPqYuW/mPnll5gT3okKL8/F
/xyEBbtpCESXdJodE3N7KdOhlNcytkpMiVrHx1VbNHukKv1Y6REuLZmFthwS
mYFfnAJCaYUj4xu8buDk/5wlJlZ5z3sPUsQJhs2n7dWDhcLI3uwNyIabaEfY
nrB56TC1D7neJarIxq+bOit77WsBCMhenLBTMm33G/1w285M6RP3a5Ze/lm6
9nkz6cv6WlHPkEi1HUzeHzrRSs/Nf2qvqlkBVelgie8dLRpOvLqKK2opIuMA
9LLq22NEr740uxfDsU5IWFvPtqWqoGuAvxSSZ49STw1Ht1Kq28lEv1P131lh
6d0tKkKbQn/CmyFZF1z/A55ZSOecjKiaFF7ZFBGIFnLvWLGYxElwovb/tiFv
pj7GB1onJqh/fnxMqDhqWy365Tv2xPDuIMelXow+pmnedTqaXUNNH7OzLnIo
/6r2xNmvL8L19g9T1IuY62JugIG04Vr8IlK7v+1E2e5bNrdD2rO62MgbjdxU
VYKJGysLUUYVn0ddBRArQLiWsKI8UM7U9kJUWLdMUATunMbjo9LXHZ3UVExD
Qmymc+emAssUfvkN4LthzyFqhl7K0kyGPLuM3von+zN1WJDETKH1VhrauWuj
fMV3PJ35IUtFdkelRxRTXNTa1AIRdUyXeGm4u0Rwgx68NFG3rWTw46TxBgIN
+AD9nX/sXnJVgfTI/QjKE6W30JG7Gzedv/c38cLIPkZMMlIJNPkkQAbU4Xi1
yIbvlU2zXwuATqqoRFkxPDNZF7y+v9CdkXrBQT25Tx+duGQ00PYJ/tCoTHZq
CWeU1k4FHWa7Q3+g6ZiczI246OlpGLDgKl7wftt+Hl2J+rjWa2oaKkhIQGJp
8GSokbzR09Www9Tj0IQW70G/jBO15BrdqdlpICtmnM7Q2iqg/3bFNIGYe5VC
5739YnfGWisEMb87atiFE4VcE5O5Fn4usTBGwhEyasLd2TQSgiYRCOs4dgDq
bUbSqJuDkXHqMpg9VhVo3Xluabri/B0FnimY6Zo7tfIBnO89E0lM21eFgzWd
fZjjAm3jqQ9RNn/f9pnYYwIQrY/dBcpO2CCK365VCGeJsTucVxATPjUi8wWq
5+T+ll1oWwMsKx4pvDSBSDAKXd1K0FPZiWD5hznMFQ44XKr7x/nrRz8jLypy
imXE99MJPS629coT4Jgyyw1sTcaHlxJAxAPU73BAgs5JVBXwNKb18DHiMuAF
TnFwQiCNIxpThMa4Q2lrHEFGwy/iKLkMu0ti79E/xXqQ1Fb5XsYI6YZOB/8S
6LqXK/iTWPNsAzTXG6c6DPDpLGPtCrEgenqCWVx63PRo2niW7VO4VqVjM1ZF
3VtP6H+zzQDgrZQuu+tIAJFcaG/KGDpYgSPQ+tXBDcJpSs3FGRkNvhg2+vxw
8q2LAimytgE4wUaSsV02ZQ1H84Y/BTrne90O1jTq5/4usHBuAHBVvVZ48kli
dcibMjMwz/PH7/O4QN5VbjVLqgyb38h1Gc+k2of8ZjeBV+0KCN57gzcQyH7y
rf229xhUt7XGi254Fca3n6amQcM0xLVWqxGOTRqbQxLpr8RG0ZD0rmPazKI4
5acKrifubO3xW9Fec2nesBO9Axt9BfWWeLZ2sN2UCHHN76TXAuli1lTYVSol
/2NUehsPY2M2Gc1fSffUSKrVlK9DyMJ4J6TSQzmDdFBKIXXrnoXNh6NDPrN+
zdQQTN0qAYCoRiaUqUQnrBs+4sqBmDGeiAOGPjunwkW7NcuSqEIw9poxglvP
YRGA67KAuiKCq8OqQjDCrXRO4i9/GvbHYkDktsm1SmBnP1WXrr4fP3u1dDV7
9KzrHLs9lx7R3mKDD0Q6KwpkX8L4V7mqtpqe2Mo5bxTXkgp2O6CIJaFs9A36
CpGU3vTsBZVflKNcnjXxlGb4EA/QlfJxkRNLzstqA5n8TXyCkixMU3sSzfaN
spMKZrN/bGOtfNbQh4u8fEXNBXBwLxeyLoT6hr48Lis1LQ9kwphC453Pxc0c
SSVBhRVv6sE8C93Pyg54h1SfifBwJaQl8gJoNa+czMqi+Kd9wMhGNZE3SX1q
JiNox6HC5mrb5S6lmf6pM92lW4eSh3dEsUIXw2oftwOY3SUc95dgomwze8yz
8Z/vEAj5bFp19htM3oRQ3XZu5TgvcoOzkN7q3yAU2R/zGvOsMGoF8PArwi2h
Fvy1cR0RoZSfnBQ6TtwpOK2BavzHc8fOV1OP9QqUqIZC+4K9L/yoUIE8JQWI
vFWQ1A6DPDbEqswxsTMHFHfX/YcjDgdbe8OjU4Na5L6jutTqyuLNuLUrN3N2
h2V+sa0tM8Ank37IrNOpnkSUkgi7byvZaQLY9Ejuf4LlpMMHmtYtyRf4M8Gw
UNG4oGs0DrFHgSJLAjorpWOe+g9UKdCLOMFnDDQTq/OMH/v0rImabf1cSyNP
Dr5DOsMxTxrBqjVRuOuJQ21nPrSkUueamFASvWxtkQxJzpeT9pH4JSM6+vKN
fo7aobynNnvtlaIjt9Z3AfDpNWN0h2lFRuMAZ0Y/NS/NkmYJdgDZOIKyNlQP
yCVsbJDdCCEC7smi27FRH4N/rBQAgl7KxW2Y935GqCYoU6tF2ugkhvETXy/9
IUAQ9hNvcicEIcdLxNevMZSg3TXqfhlURwTF8yN7ntsKZnWqveG7wLEiYabP
8WpiOdssh6X8dgK89BhGHK4FwNePAiL/+opDzoUdwUze7wxm68K6+ppQ7Sfr
/Nq275I+6Sg9Nvj1z7LGAQArgq67GpeZia+Y3t1He2BoIlGI30Tc5qCJZBx2
ZiYEIt1ma+pyD58jcjk4I6c+2Al1rulDAPdhuZzxwfcX+MTM8Y9XNcnaGhlb
mZJHFTI4J0MF0UXKQER4TJnWOZTGU1LYL/QvlLrpBttkxndjyMEKAw1UqniS
Zs2wExHYBE2Y99ySYEQ0jl6AegK1FefvSk9a4WLW/OF8D81zmS7msNmCSbMx
JfqjbJB0t0Meg2cYpMie/+M6Dh/eqZ+A52w6FE0SBRBmrviZpqbje5H2G9+T
0pt2ZK3rNlmJiU1ZEVVBtQZ+z2dRhHr8YtKRf1K8qqtg6eWCSVkAcw6en6xY
Ud3YH7YyvA+wPUaaJfefdUgjV8FwHYgBmUASiKI5Egtf9XKlidWpb/ELevGQ
I3ciwcJ2U+p7KFxPGDiwE2cA2evc5aOM//eOcs/LUkMDgqZOl1kKnroA6F2/
EcyN3L4dyg66yJ3oiofN1putP/pP1v7rfJXXd22wCbjuz4teVuwhgsLWMqb6
UnxPSKgRgngf6YUGlvndP3fsM4xPgZe7yO/Zwwp9o+LpcQXx4pMrpetYLDQL
I7w1ap6RAlITrvRtTe1U1YbBclj2DcGVoofivZLDreyjZn6SI5sylt8g6F3h
82RaMPb/Bs45hWti37dINbLXF1zwSkOydzN/iJIyPJcPqNwOZ9vS3b6PJHmv
tOVMwCgGCwiRliHkE5/DYH48e9AgCavQuDBl8nXwoxrR19toZwuptakCPdyv
f4rEsInQaExnfJAQjEwfCeLqpw9IoG9tK4AK+BgR0lipKwhHZeY9bDud5+4G
liO+bRuuqDxjGD8vqUuWwQ3ibd/ySrzXz8X9g8DK08YHozdVpze/pO5hyMxn
PNsLwHAgxrjuXY+S/A94HEVXvgtbXKW2lhhMfweh3cx1mkRshzLaAuJN6JTF
EP5hPHc5kfcEusFSGvbAiejd1ExMiHayJPOuKHDTOf3aEdVsEVjYGNv94j2r
T/cQAiCV+x71RGSvmn9AxDGAIKhTngfsuOGg3v66MtQjZhxUPwGL5F3AhZgP
vSaL6cVe7dOMzQRh4hNcnoFfmbPggg/Q/nbi0Lc+bj99H5CcCgHHstmHcYN4
F0XTClMdUbu4KSITnqfb74bggqWPELrpdGZjPT/xTh2gKsLxHkY/FieUH51u
hKPyaGa1HZISa+nkZkpFBssS0C7nLxqfSHbfY1Ye8UXhk/mll9vk6bcVgfQJ
Gc3jPbUN302kSZVWJhR71DuiByv4YUCgIPBkruuQlQhznVLRMn/n44mIBKtg
BKUaiY4bXj7dctST1w10Kfznzbx5QTxHRAbGdWBShMZFYCQ5h8sYkcmGCEOL
1m1kk0OexvuFRmrGVFbzFWxnfunDStufKJ9NRXGzkmqfaw70CV6i1BLeqJsX
iUv1uEcnzFmTDZlYILjo7PGGNWrq0q/1PxgzMoeLBnFbtIMRXEMtMOEt8aJu
/f/zUEzMxH/uWqefNeWGuPH4whrCSS6KfSo+Hx0KpVfZLemI9qBJLkHqsH3G
SBBEBX+w5pBFX81aV1/63MQfaipFRQ0LLLUy3hQe0fX740zIpLQH/zZ1lUu/
XZLaCCYnpocB9AyQ3rXwEwlcKfhf/3kTR3FuIiaI/eytiMNrAH09cyAbzOCf
c3P9oaDzsAVYH3h7cqAe74yCltzcVeA4jC4EP0t86PiJpfLojSkRZFllnuaa
TpoN2AyhnnpivoB2mLHXGzxwf7cRkTctza5Op5VbI1rlOR4ACGZkxdH927gS
liWkOKQG3Wt7qbOVvE86QdxvbLrpDX5KXKN1LRm2AT9L3nFTogXgCJyVTT7w
viUQLGDEzQv7NOliY8UAsxcsOhFTUVAOHcRYZKbJZw2+q3w/MNeUFdolzM7i
synLO8ApYRupwzDU9v3jYYCdUfFO17mwq+DNlIt/N3ukrEdwy/M+ZaJt4ljx
Cl1fBXNjNnmV5cGfJpx7IikMQ+xiRotPdgYqHFnl5XawLhFTMc8yiZ91rCH4
7LvZs7c9kYIQMo7oXH7aec21bplB2YLYRnguzzuETwiN1Jpg93Xy7XOlLuSO
yauxgflh0G0Z/XA/UIh9FtwJyea75/203RhHPchyrvKgQrWcP5VJ1a5NbGW9
ef3cvn69Wk9E4pQcEe7WRjQLck2nces3YPdYzENxV5d7xFY+wRMDFnA0Zc4M
+CP7jPzuVS4GP/jnlKQdaWEe1sbLoGOCW+PPaBZK0Ftn9tv7enQoObA3XNmA
K/zPE6Q5oJs9Za1r/Cl4XFJ++ZVhFUa6mrbPHEo9nLNvzIHIaft6AON2OPz0
mnHjlMv6+niaKnyuZ/tRA7q0ggK4MIheZiJ/FA2Y8vovEXTJjZidd9QwzgC0
41HLiPIfLXsz4nZXw6a1jn1n5ANfvMBhxk8FDxZjk7NoPlhujPpLljZvIP4n
aM5fBZHUQB8vsH1QMMIP9MZimhyFsRZMlVUAZRjSsmW8I8C2ns/EAZw/C72s
YCm1sxw0+a+ya0Hs941QEPfAdBpRkmdW4x2k5sR8bmPVf/+Be5HoVW8ArvnY
eqjwWl0RMbpxUIcq5zvQOJdIEg5+H78mfrsKGMsK84Svu57gE8JnIgG+EBxS
rqEPZDp5X/4+TS66taeRmqC5w0xzKSPs/HP4Ft4PwKr6INPM5+zc9tx4tzWI
pwkJ4iI9zGphaJGyUJyxLdqo+/Aax/9ikD3rEon2CcolL2JjOyStkySbVkQW
hJL39TZXvpXz2citKCV6dwSXWE/cWhB5e1fYf6h5lq34nn7jm9POe1k0ZgaU
vNgMfcK91sRSorX7g/Lp2eiGhRLG3rgjM7VVaP+e09a/lxwYIyc/g+izDYcp
iUGVEA15gzVBlMqlNLlCDcQONuLszsJec4odP9fKwsAENm01AVgaA33DJ5mT
MsLYK1u2RsHPTXTX/0L6lh/4jIBZyGYivNN0jO4qO0Pu0Y4eMYVRZxtBo5m7
jYjjxfmFc3Lgl+MkOxoIjTmTdWhHQeDr2cR78mrG+XGPEefB84dl/YGQXJP+
sCyUQJlFyM4DzJni6HNwvzmn3I/I2nuFxV9xwDfJl7LDinUCU/io865OaR3c
9Wuc/djgY69E6WVr4vKcePuGBm+VyBbLKpxjjg+v7xQmrY7tEfbQvGAiTvvV
O4IxGeziFztf2wV69fHnezeNDLXQqrj9bujNnw5qDedfS0Gk1+QrplGkK0K5
h6KUTHNOkMzXvlpZMVlRo2sHit63If7Llxw1NXg1lrKH48lyt5zfnTY1XlQw
2sNCHMjRXEuCq2gWqFnEyN3bcU9iy//LCxqJQnhoDuDGqIRzQ/jFf932FKRo
cMz2txEV4vDT2MqHIb6v+GXQbu18rI8UHSy1OSbn6P33Uf05C8I8V6tMAMgB
HOfyJsoWNBY9BIplrVMN0PlB7r58MqCiUhsredWeQMP23uUA4w5dM8o7opBA
B/dKmDiIgM3m706hANZuFH6gi4+cUQJ6pmRbLdLeKrs59BqdTGwDEn9TDmlf
O8UAWs55IiIzVzo/4AAxnaUgEITF5YMfRW8kNJ4jXcXmvmgrqome8nSVvj2m
LnyvJALwOMEVAcyKlkXj38Ii0KVoOJXo8x7XdnYp7wSZuCaZBYx2xdy3u33r
yaB/jBfGWbqicgbA7orMz+f1iVZYZx+NgeKNpXLnvbAPRK7eoftowmx96f1G
ufhM1sOB9NaG9cwPd5CkE/TnXxqk6PKEMIOLMZbzOWJDv5CQebGkEjxpurBb
oAuliF93ObeM8cowckgdlVSwWYIZswi5V3pBSt35NxIql5O3U/0IfENFUXBL
W0v1oKqVHaPOSU2iC4S7MQYIB8wjNMS9snRUMHm2FlmT4YFOJ0Qgc1voE+/C
bQGDvToG8k3sf9LrrBEXNqm8Q7I5nCDhg4Jh6fFIe5boeXYLmvf25EAAWJoH
nKyHqjgZlTXxxQQAPrZCVe79cW/WxlICeuTsnoPcSuPd5RLx5S+3WoLEIDBL
vpz56x2DyUGtpbHOay+i+vVlM/f+kYZSYr4yMcGvBtgNpZFUXuibGGsJRjX6
ZlSDPH0tg5JWyfjgHb450R+Vbutzvxyt6ScStgb5gmF/Im/hkmTIWpG590/u
1Wlw0LnzkoOt2dYGPFsOFjKIGTyYtmWlnUDcx0PiHaCYIjSvTsOEsFeezhTz
NU8fLaLDZ3yHVXWY3Bnrv7VP8lTKn67WILIXNPHCIyotRvfHe2F0YNPLNHif
JtaKLFWrkSrgDfuyA4eENhASvOKdyo9drOvbsvx0RCbxX2gGQR7rranVKR3i
LUVpGbkBUtGh9VI5FZXYLmdeVjXWFwb8d9H5MOzJUAbpAo5R4swFjoAWRT9F
py9RgRJ5TudWDdMCSD60if5+YrhFoTsERJu206KbA7lFEqTIFFmpqFZFo3G2
tJVgytIff3COCpkYc+sTnLpyYODa6FSeySOZuFCCsWMZBfV5pCLq161xk0re
m0lENXzrwO4ptPLfQvV4ACbyVUw4U5LeYZeD7lhNtBg5X9jtzav3FuNu9/20
pw7ZP/awWzuxGrsJqrtHq/ETbwAthmnMTBhgI4pKi2AzZZf3FPRvnCTtXc6m
NmB2pbyhH3bkbna7EJaW1BxsLnTCBBI62fIGr2TGDy6lK/Id/3pBxlWwaS/v
6EIC9qNL7Io70KDbqEfVSojuQP/pI/+gtaQCjcwqAyrDMlxAw5trmXq6SGj4
by6ry98zTau6IUx63v1UZG3d5pEbI1f6OBNIOBMpamOhKxZvoikJD0YKjjvv
k85e5j0m6/wHIGq0hQcxYRd6tX6ef5UDx5cQKkh6T5DGuUIPRMRhckhL5TYS
9Ugb+SfVZPkFCHrPzL4Gx9ZUQrCZJpnezJFcG5ffl8DF3uLVaNVSlBJnZ/3F
znCY8nLUBycWYOWI+cXrV1CnPeHzHCuOwGklz0qwaldYbxGXeTVqVaVocbwo
mA2GUETEfu07OAUTcTUvj/K559wSIDCflAO2py934fpNQmOTGkkpfqVKVx+O
PHst3R2SRWw2CTINnRs5W1Jf3D6a0aS/7RFliSlD/39dbJo9Jbyc++yrTLrq
aig42qRU5Ab5Ht1LERg68RFKzvZZkPEhyxxcCfASdFHq8ZRP0X41CjiYZ+Lb
ysg9WYkdVm57LZR/qfWcPLdxBeMpozU2auLSjHpwZHoPnUx2TW4QZE2Wi286
UTw+gHtB0XEQ5zI4yJvux1R4uJHAnIMWEYy1oAtmUpBMQZshqrqLyGfuwmvZ
XbaOhnQk8iPp/BiZtm7Z2KMDniwXamNPEKKPtzLVLkjHv01sQ6AC+XMocVWU
DkLsYKg+1sLAXdq1Ss61+T4CTF94cOWy0BLbQV+fbZgI2jtYsNmO1efy/fMH
xcZgzD0Kw6m6eYcNApCENbmwsLFY929caosfr+VYFAU+C8EEdFzQB2z5Ehgw
FvHgfmNBu4FYlzaYVdhY7ofzAgjzuLT67AkO+p7rMpJCcVVQT0ffl4nQMmu2
pGEn5QQHbrVSNhYY+8CYO/kPxHpdCQA+Ppqe4LHzVtvVyBXROdAFxT+F7u8X
C97nJr+Z5mDCpygK0v/wZLnltod6ZsH6q9xNZTA2g04F71Ur/2Xdcc9nxlgo
BtHMit1RZC0wpEMhGbwtaHCYGoQe53gJCNimlvqm79KuQdX3K+KJ9H/HTnor
cNLMggRGYFGp5LBIITWuRurfMqigX1G3UFNy/PJEajY+s0USygSXx3Nbp0wc
KtmQfDRBqj93+P6IVSIWrR70J5LJKzIVHJF6Hu5aAb3gSd22PSSRAnFD1YRU
61V7sv0JjMTk5RXgSTgCG2S62Vn7HMExmnfBHeWSm6oELvd/GFFTMdbxVsoS
GJhOwizhGhW/pjQRVawiFhzNRWmvhVsS6oTOZ9AVVRLje6XKDs0qm6XIxTPK
2Nxc9PGJXPEY1gpCoKIofByFHZ7phlddEmeW/GoO0iDKO4vsYVZhFLdmnzZc
cyDeDbDm1MXE785HtyYTBCrAU6X1u8XuLKV/2ZIOzMBjiG7JfTRHMIDlG/cK
aMRzMYMoFlszmMSBbw1gQpuIU7rFfT0+YzUHkagRk+DFXaJ+aAHI5GOXPbo/
5YGX50xUAgHwB41xB6rH4uOReri764uwPLuQ5s/QuxEpM/CHM0yc7IntdpwK
0d3fhhyjUz3S9lFSYL5mxIZgp5SytuBswGW4zIp6P8iFfipf1D98Gd86dE0+
SBUgtnqMEe4fnK80+0/k3ixo9kF1TNVfk8TtM8e8e7KCQbrJ9DNySh7JMGlu
LqXgXgCs2ftyk3leaXDjzGTYcGENZ5Nf7RV1t5QxhrEdrUh051Vma0x6mzZr
wjYpcvrQMBTUiEcNxwVk7iOEc+KnXqEGDgrgf70UZekIU0Gpq682o+85xQV6
7265X714rd6nsUU0b1dtJ+AkYYUHqczRZFTi1nFU2EJ64g/vRKu1nlp08FLW
NaJf2XeOvy3DysaYXqaI74YkQZlKBdOpVGosU5BfBQroinS3N3OcmaV1AlzC
VNXdU8YnmYgjC4oaRsXfSIOWsXq2C6l4ebC1bVlE9zsntg2clY36kzKEKKRe
rsFb+nKtUtwaumk+rapwE7HvIOuo3+27YTxbO8yxiTTTsXWmqOC1pouWmixO
DqTEXQDnOu8ALuzS5KS/LJfUNqibFPKVew2RXMoGZeUh8xja3WMTl4jaupOp
PdLkcFXlY2djgWoKy6/GqsNKiVYynTiJ7uliYdiUdeWH75HosdrRSLk/IVwA
2b6MAQu+2HMiUzlaOmw/MBuBGvquqQyWhgG5FplN4U+EYNu9zUEFYb2xy7kz
3GFDbHgV9+K9RKQOW9d3DnSUZorqwnU8azvK0foc/zdH8eIF8K8CJb0b4Apt
ZpfPZtU0OGfYzXDkEnhzpCGpbQYQKWA7g9+O+0AUZ2IFUHjNibBmt3GACETJ
9RteF5oNyMYMqPqK4rjFj0pLpAxSQuG5sJBlAII95/zst6VvgPOpFvq/ONX+
9bAUX05mYnkV7X/mHj7EL81fxYurUY016FD5J5QJBI26ZgtxJVaXfozO+lIX
zHxHQ7tnfSI9EaPITi8cpFSj7tnIsvfrhIDyFDlwDZWK6ABTDcMcShMzCAyV
effRwslMvCrdfBsR51H+qSAY4+LZF0FuXb5yOnnBQDGeJYhcofIM7ZsJeXZ9
HAVqyE1zsxAGfa8vycDWkYbsYhtvwwbPBQnIj1a43M+V8ooHZW+e4XDYOd9Y
Klx6VRXT5I0+vDAHB7lDps77a2+KbGJCWEw4YqAV6OFW6CelgRWYWbqBJrqq
V6Nvr4JOe48wOyIZB3hIFdwQioWDmakV9V/o50KYFMw44W90EcHYolymVDNk
Shk818iHGBBVxiD2+pT831CIX2TEVjqi6xzf9pSlE0GYgHJ+n8V4MtZtI6kT
x602GOzvMBDy2thJDJVFFki5xaPLdnhEi1QcKNE/VkD+Y2Z1H8DXLx4R2n0m
zmmEGpCzLUkPDkpbCrPrQVV4WOcYOCDhEAv1424e6s+y6R608eT6vtsOs9jg
u0R+THk2WDlWtTR9EpjwXhnr27PEobOj74FDstnO3qL2paSG7NY8dAjWAcX5
wkt4XZKfpKRXkM+PzXKggh2yOqgGKOiqQ+qW2Bgx4VV3oJSDMSwAf7ZKwvn5
sb69FSPSZtWFKQVkvrOfCeJzC6lhqoIh+ck9OAcwi3XKFTdkxVnNBeU4QabB
gRHtardWxPNCeus830z4pIviih8bGVKf4GyXvgNyqIqN/PhOapVooDp264gr
i57HYHBHl9b48Dm8DHjkDYRC6FOCDmujUYhiS+QtpEXzA9yZu4FWNyrOFUtK
rPZd2Fecm0JUiqKGp4lGm0k8PXl3ZOb6sYnAg3ibfxj421P5VFS0WsT/gTqU
1bDTLccB9qImHTEUvGLKFlVwOyUkEWj4YNZukViBHYnxvna8UmeVKda+/mtO
fwl4KCEox6R+hooZxNQNge6fuhiKtCZPxOvlUBQd4s7B9yEsO9IdqQ2lMjVD
aM3HwZUNrZiWAkrTseQxqjse6ijZ4X1CJ4nppFbjdPDGN77g24E7lZz8KMbf
k+oYOS/4fBY+UHS+PZQXISOKNJjiZTuUDLdUBJ4+56DFmjk9dN73dD9XSeLZ
e1Fvhk0wqBgfPfGMAdq+WQCKDJcWNb6jrs3RrVdD16kdma/Hj8Qg1a1zhAO2
IaqM4WbAYc7+LcTqHpQpX1a/1RRz58VkQyrXyywm4K+aMABtybB2CYkJK37Z
lRwsbmzRVURNWcN1rW46IHb9MlS0n9DW8eeVDr1fx8D8IMwOvt4R3CptpZZX
+VrpsIAStxokxMqJ/DW4rJ0CkA4A+nZ/OYGyJOQT8ZBbw36Okzy4oPbqzv1G
GlIwW6Svs36SoV+lelEOgWXEqQr0C1jNg+k/eFHFWdC7+soXuAkWdS4UV7qS
6COMVNWht0ZUSlxAC+DCHFOKI0ygXP0OTHP/vJVuYScJj5lgcuF7ggMmqI0z
YqMnowNDF7JcEmyIis3CPX1INEw3Z2r8Tr/n/lJWjtXm3HjfDyxZEKsrRfX0
kpEy0hY+c6tMwr7s52jK8j59LOwHS6C3ZZgypa6+mgZCI0oVzp+o2cXXokkg
aWIHl4MIKmWSXMBLVPN+60XSVKuEH68gHQ9QvI++WOjzRqBkpZBY8fC40NYd
OJKl1zROHVjGBqKpAnOLI4Y+IZ+iYakobxa8ckuhow5yAQQhAdS2hTwEbfg5
GjLMYqDg0smp6jfBxphsjQepBQOVrfjdc1Mo8tB7r2s6WWFbsEBLE2MiEbnS
0khMY+GqpY+op49ADPsXeT0AhQJYRKMW40X0VF7oUceOuiBsWV/rCFi0QkRm
KgWexlmBOvic86Xo3nAiVBOOeVgh58hiv6yESeE4lrrNNLuKBWeTdheiUG99
Nzejmn3o7cc9HYJCcs91O58Zg3ekJ9CeA7J0i9zq1CR6AzF966SvM6iBFO69
kSE+h18411amO/GifU4Qiooq74LKip/d+Gw//+b/0GahP3eSotoJdAV555gU
jvRS8iqQiLtpfniNEDMZPJ2DvuaLKyoKPQgxWrXpp8qjXepDBGcCoZKJ2NBO
1/mu6Aq05VbMqwZG7GISFml8TztWFKtIAsbp5KytifFoBPSGvM2XqOVrYmQx
+N+WD9CEMn/wZaSrRQTtc//buQbM60/qNhl5Kfa/2+44O/fVl4oYK9mGt1oN
VxUNv7M6c7PgsXEGPCsfuistt+xBqteFEOyw8uaj193l9IsVWqH/6y7BP+vf
KM5eLii5kTdG4+EZSHcAyZKQz81YqhqBK6+aY4xv4rXlYntf/EAAfA5qoJrh
Lqsr+0Ug5Bk8s819kI9+PVcb6LJASfoHZi4AZYY8wy/AxdgO/e3QDCIchbZ+
7C1dYxS/gS0CN7K+g76w5fzH5Wqaf2E8ajM4uTdpEEiTWZ48A/1KYB9EEzrJ
gpfeyeP7XhErBxENgOer1LM2mN6+ZC0w/7O+txIFrC67K4cbOEZRPah5GP3c
r9l2RUMHFfj/tBCliRjBpLXDWXkqnJoZgptplT6EENYZ8meAnbqxrFGv96Ow
Ys2JyZCuqrhENjii3Wi2QmL3qsbK5U95+5V522Y+8aRo2uq6n4kSGd4LS4LF
WaooKMYGXN1cHbmYOcUBpmO1qgl8lxILGlzED+hqQUu33MQZxpNVVOC2yUSX
c4SdQNiP5hrgzwX5HNZicdrNIn9Gmn5xNm2WYWeDsaQYhrLKb43+kdEA+nFd
RW4a+fGZSrP2gYeUbSM3Iytck5qvoHkSMKi8g//3PWw5E8sZLjHykV3PnI2y
ChcsW4dfr2vUjm5T/zyCZCqqC0y5jH04rfvDNB7IX+vDhP36o8DGN52NzGhJ
y51KDJs+I3pwvyP6+z5fA5vt4LAQsuE1EmnvXigMTr3FHBJ8jMiqIzMlN7zd
7uWdaQPzrW7h0lcVXeQjt+jnKaVfT49hAb9UzNQSnaHh2XrB+c/uEvHpp3DZ
+gg/fGlJq7uRuCp2I3Aq4pXry33oELXPgOkeMlgcNE+JA2eTW0ipeRuZw0Xp
e9CsdO1gYmCEi8GOAy9V/lJnU6C9u9EcKYlI8BNGnPdPl/8GyxRsX79m+kkZ
CionD5IugdUmU0hTbRP6xegqkIb/NGj9UCqeymlGRD0dvKanqTzQG3vOWPTb
WJcjgi+mYd3n8xTWUWBfJgqXAPDfYYThI9WUD6f0QNfOIF2Neh9tk9mvpJF2
iExBO0Z/Xnd5VXYgJZH8Z1IcuQ6wuIMp5jCOugh7204VJ2c82YTK3X32ghv4
gCeXI+418AG7hB7fh/y2u7X4UU1fmL4N3qQmkXeu/A30QW0aGVC/WOue4534
updw2QP60XQzi31ka0CIAX3jYrgzYHr0ej4mPJhyBQthXLmNqnpCZK515XjQ
S60BX6xcxgPhYRmU40pPlWhzHjLwA2S/p8zmKkIII8unS3nN1vn0jHRYsDEe
ztgJmsnNPXkIh1k0sRVncq260HgFKhxMP0+QwpYpOKK6hAd4lVjurrgkv5UM
2NUyFxJTklHLktyjogxDIdLlKi6CX9Zdc1xEzJdP90CMHUSp4WGJpxA8WkSY
FqFnOeMZTcTOkpW65lT7byoOulrl+vlMpEtBTfUtMUSzstaKz6fBYQlQzrWW
PhFxMtm5Fd/nGJYPnSigQCwF6YaW0fjPBbW6StXFxrQ6mE/nacvncg2p5Z1S
c0AqyF680llEaI5B76pv/+Xn8gVCk0+KszRS1lnM9A6Hb/4bORS6fW1FNJQo
iq/bhSr6XyBtcHtqsubDZghqFi5gLVbllxpAE3XRZXFjAJp5ukwCxKP2zuFc
FRNfhDGKBh4ADOshJH74KfPrXGX25IiUZMC+GV8Y9V8ysZgTRdIKCTbNSQSS
71VUz9xuXujcwo9CdqpKv9AvYE1rFYX0Q8ffRLXTOpPfiLAmwXFcRRgwMuYj
EPylLu528+zdu/Cf5VHb+7lw9kNmF7F3tj9AL3cW5fzf0EAvPzPtQQJMaBvm
md2n5O4Vzk0TICUxwh050YHk98OM8/kPgWqy0ZSjZcMP/DDFXXPDgjgke2XA
Zis+13dsiCvOP7Ma2JoaPT5DHbOzuZMX68PNLvmggG1DurRjJCPn9FBKAbN6
k+waz31whBEQoY9ijy62wXCmE0KHalkV2p0WC+vUm4/AUjD3ldRZDUzLTMGD
wZtLNaOXVTVIjlxhEZQn0ACxbvFW9gfWoZwoYlw8milEiSszLowEO80RlcFn
/bGaiigw43f8+W20wa/q6wsgU++wPpMswSdoyPlH2csyhXNk+p26+KlLGR1j
RRkXP4Ccqp30dhttLESnYvXmUrwJLu3w/W+SoSJky36GyLa0txAbw4aUUbCI
2KDVVIYLpaA6/JqX8juACCVdmHk9XlzNLoe180c5VymK9hVdBkeb+3z6K4fQ
O77cm2FQXlWBoeqRjHZgpj5O51RilgVVAB297Hfn9M2YyiDoqthY6+3UryPA
QOhKZ4difO3rdWQAxqGlGz+L3KqM3Nwjnl9VslEQ2Svyx91y03a8UrKKAoXh
yW0xLt9b3uJMNu47A/u4/nPie4Xbw/VDlRFt3je7JuWPrJXxV9wGfEhLdEGs
dMThMDZWhZ96GoKGkwM9FKkMFCBuntkb+UIYr7NjVcSY425RTi64YDlFWzwh
PMv0WnVhmDwra1SB22JEBIt8v6p8Fp6NoCTcTPVdJrrLx3m4QULfWzucRd0u
LR+1i9D/rsJ8jP5OuVOhb+pNstSu1b1b+bS9TiqcL+MbEc5IGsspuvslc9QX
WTbXn1zL2QAEt8gQfs8qjEKskbRYkLU7NKbDn/HbfKxGIlyEFjbiEbVrcdoN
HNpfuqYrEuPQ7+mKmVOXF60kO0M8y2E9oJBsv1sp8MwY6KQBjkvsGJzxi2BC
kRZ1G5Xuhg7gVPM7xeyKiVRbor619/U8HdicDYn3pcj2vdAXK6TYKU7wrpCX
soacKq4E3mMCBrcfZG6sOrVlZ1uMDYSSY+phepsUXSYTNV1aE3hFKSb8iNCr
KqLFLmJjMUsHl02vMFmL9UnwIryNdprpMtqI36CPD77q2eWwVqzifaApHwGm
gxgWv5L1bHLDg09CQ47WVQUnx/hM6tERW3/bXZkQYgFSwjNj8kd9qtq+MpA3
pHj7L5wAq7U3WYwUHM4YhB/tmAJCicRC0OoG0jjXv1Zi5489yO78BIxbCqU1
wKtbotAoT4mxWNwQ7p0pRgfzCpDTrQouQ9EG9idNdo7zTOG4zuD2xuFNfohu
ysf8ej6BJX7PngCvCOFjCK/xKFGJfeVqMT6JbDJxALCMRpdmaLClNaDCusWX
CiE8jkjkCBwo1UDR+HR8tp71i81JIIvM4inhLJ9V/ntpJhJSq8qspXlEmGJf
nasVzhpITsPP6Mv9GIHLfTPs8JwDHME1K+D8YeW6d7dTF7yaiH6s95JIVmiP
shFtsHGEXrtwAoXEHqGTxaz4zERf6tmAgIoAqdJNvD+JBERWqr55SS1YGRAu
sG5iComrfuc8W3DFuOhTfieoOJqeBl4++m/8TZoBHSzyULzG4RFRO/ypHlCc
+FK5iW64l47leod7l9PqAknbkDtgCUecM4ZaTN8YeKJ6Dy7xPoaUI+GohWEB
PeZ1gjP+wa42YPjwbOqLQjr0TTJb6Bx+HOd30tp5AHjfWrfiIcAUyM0WMajd
p51L+apiSKikUAU9FuPbb575ZNc8GZc7FyXOLXsvqxzMGbNUdB4CyiChBoQY
kSzolcmtTxPHqvpKqNvSUw8ncLalscr35vh56KAW8L+2waTU2YltPjOfHDgF
T0QGjsFBDfnaFOHImxhowiJr7UWLq4u8/lNrc9M0GfJT0w7y2YznPk5FPWdp
qmAmTm1bWY7NLsre/EztoJhyNlJ5x+qoZvuUQRV+IOXwSAsMAvaxwJkmQLWD
tDr922p/2RSBr+k64bSRPbVFANZPCCj9nBwsCLuPzREIQ82WMv1RmwWa60Yt
HAsxRZtSW//gaMm+ptO6P49jiufFnrQdbyBZ/ZpQcN2nCFf8EnrOCSzk9Ox6
hB39SvzQN+OKia/hqqsdWQIQA+bDJr2FOAwOs2XqvbM8FdAlmaQxATq7iOYi
O1xAa4kMpVD79gWWoulzR1LiR7qlBQE4W97K91jCPQbB14Q38zr4LaMdlk39
ukwWw5bvDGMHIK4JlXy3tVU3r3kIbcPXVwfzFQbtxf1qw5Ah8w/LbjT0fYrp
DUV0WOalFsSSXqZ9kG0LtfIE5CdRpQKGouxzPYr4WGqV6oynXqfOAFa6aLDl
1UWogUM3y32p+l+9+kpA3IEYMbRClUqUX4PuDMi9hY06SOKowAZSbplks8xz
UAo5vq6hkxPkMXg5dMs7fsjGF5KykZK4d20OIHzeiDOVd3ta6Ee5K6ZLDPpW
2MMo5ycf5mObW16LHmS9dHPizd+bAnkYr0jakPKkhtbcJoSPj52Lj+6OpyIc
n5JRtCeq3o1pQfyHCuxKIXXKvbsBRbvE7265gLzATsR1Lqc3kOqt4i9Fo2I7
jGr/LljYXf2InV9kJzaJafvFwEv8paXISckVInAnax7RQ5qzhqrRIJOUYOqS
W/QMhi/0eINgdHCTmPinp2kq1AcdDrSpEzNiYlXIQpx+wQt7JTsJF2C4SV0T
b+xvbDzn4jeUBCXGI3kNlgshF9XXgtlnr3VtHLFfZ3ZSccJO8A70RSGq81PG
5etp+wPAjvpUSBJmJMzNxXIow3dS8f9a54cz2suh07sY+1Xv8+Yl3wHV/FZl
luWkZYvpROlpoScsGWc6Yt5nNW9UtL1o4RiXziDhp02v1/dm9y23O2J8al8q
6BbuMF+Rtc1FqebnyyYrzzeQamSJA5kWZtCO3S1qN8cVYxsfdFjzYZN1eA+V
2eHVQYmyBB37mXgX1ax5V2q3UcMjjurhWzpwq9v1lce0RzzMFV8fsNoCvb7X
ZBvLl5YYEmlwiKBAgwXc95iOJkfW+xxlKANTY64qM9FbwWJ8jq3/0YCZteVe
4kco4Nr+YY3Oy8yACVGXBHYME6RDlna+YVCAy2WUUhOBtOgAjixRqHZURIYG
qE+c5i7MDjAYjN3iBn6iMFGITCK0hIq8Vxa+eovweo0A4USah6Yl7cYP7qpr
4uFRenOP0Vp6zIXZE2owIZ93aXPRvruzXRooCJUh0zqg23Ld+7VelBYt+Uqv
pxM48hCFZRnjeDuONFC/KB82w6TttiZlvC8KeflWprrNr+12Zz9bgYCPrrro
8mdsMn2KCND1nPEyNsyLEKP0wo7/HN3G5qNFT0rhCrJgKbzx5ZexUFnOOWlq
hzn1CYxXSaXAW0Xksp/Dky5PeUecXqIkmBn3RmvDLqdLP9q/DGkl/AIeQvOE
SIInMYzG5pTEumE4eKzkJkEn9j5v9FPlaFlwfeGBAyt3LkkgKq4oPctrIv0b
IWDzsmbjBMluPPGquipECyWLbYJ8A2c1lovUHaHWo7GeNqwIsIKMHZYNNzC8
7OcNqgf6OG89n8BhlLj4XcIuIQ1OW25iV4O0422lTR0EHahBnmILPYXURVOS
WnApOsZ1YFQjxMJkpvrONoldgu/UibGOUcwnQzMVhn3kjtKphh2t9hbPH8eQ
qaUlOmtJSIxggTeAFoYbLOQbVSHCVNk4XbqAdiO+o5F20jMECi6SQ/0EcJ9g
IlJ2btzfN010PwWtWgbIPCRuM3Sro+HjKQEa7F0J1vZhMBVp58x+p5nIxpCK
iWSNeLWZrSSHUEXgne7gYfVAGRfJyzsX/JzJQfFFnBUJtDX3MjpNq3YxI0i/
V3JAgrmgA3xpAupFTtcYVTPPY7dxbIfOF0Tn7cIlYxEsa/KXnYWHKcsOvls1
yL8C1iHco3TFEj4FWvNHhbpaMkWO7zbTtjMguYjDoO7FVH7gD1g+2l75zR7Z
EEL34lT+UwrtAsDRQ1ILH2nMN1JcCfy7ApGEhFqa4IXJ5YyV5Uf24PuqXb68
1S66cjJvKbYywtaxn8xVOsQZNppzu1W/JVI3204Iu2ItTLwPLwG4KjTet+No
IiqyObVt0Bd4UhJY8FehteC6MZb4PeYGtddsg5zHJWDh6dLbwCRJUVWOD0O7
mcEcBf0yMAxnApvy0vmltF6JwNHaPvFuDqiGnXd32Iz4VDP9xZ7MI3lECi4a
if2ixqy3klWCg9v05e9SIsP87s9kVRe3/PMVFb2k6jsqTpxbDO+A6PLhFU/H
5tgFgrR//PQ4gPYD4hX9wX2XPjLhgQfHwnGFMyO70iprTJ+bgi8P+rILCCLq
kZI882vQBGTKK3o6/gjypuR1B6TO9CFNR8YDTKMPjVWTRhGBQkFgWOg3rKxl
QBXyhD5qeRmTdIo7vj7aNwk8xfOg5BIFn9FeNPaLbkgtEX1BLpnifnM2tVyC
PuXqxGfVZhM7hYuXQVjky9qywfzVGfJl3ffE3Kavc+Ys+Ab0QZXVMNSuAjAz
Ye3SETouHxxE1v/0utdq01KsyIxoqQT7mP1igJ3TEE3bUJ9qzYpcDAUW6JHY
HvjdYHFhOQVRVV5dX7CSIGFNbfX3MhcVoMCUHRKGUGlHw442sAOFL9P5w7L+
dkS/x2EiDtUh2lvmGKWKtib/yICIOyh9QvySXZskeDmxpzVRSbOFt8vHiGpn
EzdfR040latcJRHXW5pfWVgV7Ns9GF+NIpGhRfh23YvpapWomdbvZ0x3KzHZ
v8xl/CT9okFUWLAkMGW0uJRObx6ZDxbyj9oeRCvuFDT6dP3C4NhL9Uwhgrlf
ID7wn/TNU4TDe2w84NPyGQIdh7VPNSQLsmJ2Qxr/KXgPLpT35aGo7R37wyVf
tOo4fJWcACWtDWiKUetv0DE4TsfmxabEI3FSCJdvaUtNHlEQ1tTRRg2vHSmH
h6ozpuPBGIcZFVbZcZzo2IV01XgGtCZfV4MeVf1NbCKNz+BaCLQR7giEsk2z
VEeKJ20XclDMnYCEVXcadgyYMd1pmiGBujZgM4CjcC44dCTQ5FA0+/wABlGa
M/rd2v3GNqMbFle5jr2QbKMGCPAzEVRFHTInmP7O3AEK7Uh6nUzRbrP1fKfu
i7Kl6cxkqpmJdGNVHfsKk5aJxyFf3D2U37faRJgQTncGntyAUMlGP54U/kMd
rmjmRPGhbJZgJJtyfc9TWAjXPq1mPQQp66H/+56jNhrDhNzhREp8EGGKKfb7
Od7tBUnnXWf46DzD6NkQjDy6Q7YqLMTOZWMrxsT5LN0elkoCczd6ded42nqZ
aksj7eg0GcMvvhshwsMYohmJcKAVUnJA+TvRpnlSs0OuFeqt0I7zovmWNEyd
19CJRwz01mpH+7eG6yq8Q6MwOadkNJpkSyIg2EHfSOwzfZeKryekwSYRecvb
XFZcHlo1UdN6uQ2Ijzlq3PZkqqy02SkO8DtLReyrbX1tWInlgDWIVSCwQoyk
7j+LYCK/VjP7Ca0QTiVMd7U5WJnEt/U0bAiDLhOxY8qUDPGatbq8dMAf+qHa
tq4BSHlPbFbmZ9CQIsIqpfpqI2/aUzdBHDPCpdTzbQKCfHT8PeU8UfYRm1pb
Ufwlidv1iLm/4hjm7s3dgxEzs9ELqpQR1dLJe4FXcfvyxdy8kyW9nswvzP44
sVqY+8OfEQsbqRLh3iV+Ry+cxaDEyMDxdlEBZdmxj4CRvF+/M6E4XWNP3NYS
I3PIRpC0ETmPBOlkijW1/u5amidvAAGHZxMxwLHipevYUc3wwwdAyxU0iLac
Y06yALMPaj29RFXU9rklH2dX1MVcCbP1F1a+GHPv0W38pc8TxMq5Fyjd8E7d
3Wrz/VE/XrBVdV1CbwE2DP2WcD0zLEQEmzuL+JAy1Nc63yk3FK6aoDcv7jIp
jCLdVhdM0CZSz7lDRW1YVWriF5SOJ+ugdugp2QdS1hILtr3h0muzLd2WIDwv
5UB7FQKaZUfnWYcn9Dj+B+KQEj1ZGMzsMfEQ+dTh2idcHfdyizbBvWR4nqMF
GUalP34YJuowPmGUtWbKsX1Rx/qg0QQVShzNcnM7dBQiXR4P7F6C8E8zbvKW
n6wvW2PmEs/DGCAe4sTGKVbUgMeE1ns6OI1LrMZMrdCfqpKX4/bfkiK7GAEi
4YHE7oOEMpbCVh10QYqnHSQNf/66X7AABn217tDKACI2J1jHGGZgl96UHKY2
s5vTamW03Ncwlb7XlR+aTdp+rgOMWRM9tsivSurxtdWxTeKhdYHwZ0P6Ufdz
2UN4iH3YI1qR+cAW+GP/LC07nZYVDget0VOfsqmkuR7gqjiXLMpbcfR+AMXI
e7tZ8dAbJT5YSKbOw4pGYgqaW6x0TwZhMpXQ4pVhplJSI+TW4y3d34UqEecE
/o5J55/IMXEL0Nt9xOcgU57RFSo5rG/PkxTJBohOK+SF3KcUiIYiW/JudDfo
9xpfUQK+5PeagqI1bkdI8JpI7RpRh6kzZYxy2LaXg3NPoTsp8wPkO5xAYRYH
PdEwZVbm16jXL0Vs79ku8lc+tfo2SjH12AfBfXy8goDH56aBKfLfzwz8Afjg
SwjKfm/MixvaW/pD7hlssJfePF+G4v+HBecTIuBEnD3rzgJWrWPrt0oyQ2gB
Y0jZhocr0XhMTxmCElV88+Wzia3O9CVeY1YU4B+/KJufibn+cBx7v2wlbd9Z
9mje05/W5PJTn5dvgKuC81fYp4dFh5kM+xzS3+pmp0lvClj8P2lLg+/KCnBJ
tr2I6ALyARWvD/tql1iDiHDfiLt1XOGgxBUVyrLDgMUQuK9qS5AZlk5hV37k
S5c6J2r4kVCYwdKgg1I4GY/Jl51Q2ySgxTzTfIucVFL71o9Lyw9zw06fdXeA
3iVNwfDeVckkaWYbut543z62F4R42W1anUBghu0j444IjlZg9fwOmueT58H0
Bukj5Lw31ObcG38+JOyUT9EU9R+zJpYoLBK9CF7eHOykbptPsWvOkt0GQKWt
Tg5klS/ZN6RfGdApr9OVUO63vK535QI7tOdmwOEVZHFSBceaVpWma9c/fFQZ
QxzQZcg05n6mjC6Xq3kawb55YKM9K5HiAneR63JQ0fUjN/0ii6oWxy6HRYlD
RD7zJch3FC2IXgZTX0wS7Hbb4yLUUpxhroRIB4sowaS7Ap2mOQPcPjXAL4Sy
hK1H482aP2xdx64wdAYFbKPjhPoXq1YqudY8OiqKIjzTJrzx/2yfC+udix8w
3iurTeGOkoN2MtxsKxlYQVZnrQMgeSzr846sEhDHeeerZsSGz89a6sm9s3tw
EHIGL3E+LLRf4qGuvBT0uS5OL7ZsPSgYWW+YTY5r1fxVfv41cCE/T0qwbbhe
NRHWjreyBq0rN3pz440ZFoC6Pj+zMbYEOvcY2QwtoU0uQ7jlbbUvqrqqFNCW
uPRDy8KXu335N3EtKmI3JL8+J57fR1i66IBDOhb5JNo6BKf19n6+NAJfI25S
zx7XcBH9tRxjYFfqb83L4Pjh7jILSSpYicreDQIxtLC2/w9OpSVoq+MNkakb
Jyc2uyDKr/0KB6UYHnrQBojEUEgjBmd4+Y5vM2pORAss6HVqMEf6sngWVf86
YSHYt0kG0jXjx6HhLvLRxAZHYBf7/cNLLaGhEY2CleKjrMuqEzUHtRFHSezv
9DYu5kZ6XlF3RdLOWWLFHUCYPRul0zl0zN8MXUCysNDLTE5f9TiJBQxPoj6+
tz3J23+IwJKEJSI28ey2F3FUbCFK741XmJWl+rA/Jpj6lIqjt9YUBRd5I6VL
aA1MKh5eolq0+Q16nw2ivqHn9R2TK7Cq5TSDIu/2qZJsGIvRZd1yQC57PWLm
glQq7gq/wibwoB/tJZhZ+od1xbwqo8f5/e4RfzoLv++CfgfdgDt21SQCpXHf
jU9QU7E8hUlq/Qaedg8POvhWMDcDID59IiChyBQbBiGM7oFZVz0oMVPD/DIE
MJUndsLV5qEPALMQ87J7H3JG/MG4yd5A7LiYPEvo9BRjUlqUKTYxwFXnfofm
9KTjHL7/Z0j0/GNQ3KXTNxWr3Sw5b5pwS7DjiB0ScBrNxbjfNrvK9BI149Bo
eU3AHsdwF/9hlD4SSEBaynTIGmR/UYTe/lp7wRs6dtS/+5S6IFpcJPMJGWuv
Y+uJgamttgaimaF/EeiDKFVzf2/emzVeHtI9ESqu5g1YXtP3/Ccr7bL/mL/y
KdCFy+6rKgVClAq8dY3FkjaWCqTo6AKHcGWxdSkOQoBTQQPxKSOKcUKFXNsR
FqxcEGhJ3oTGbFs9NkePaGb/r4gk1IwfbOrVgnypSjAb6EfKqMTXRbeg/EeD
++z2TwHJSebaykzO0NwcklZbgR85BQXDF7y5jRmwyR+YuIF1ZRew+rbc3TqZ
9uyhG0vTo+cHhJ2DvKHZSaE8TPvBKmGJVjPcJnHVcDZAV/puV+cP3rEkZuDU
T09930FxaIz9g04K8Zvh6A5HkSazh4NfJWqNeKNE1vumuuQklyte5Or1Pnal
JlXWEmeuu6fG0LkJDKnN0oMeQuGXTl1BsIqGzi/IWTRceMjlmX0DQB6zRNaF
dTGbDC5QspNV5aPxwZrEynLtMhi67/Upy+CfFlp6WBrcJrxUjlQKMjhzxylF
PBCoNZZM04oZOlhonwAZHDUITSy/5uGh6AbcUcNBIiG0ysSXX1upx9n7k1Zf
Xazpk7TbDRcIl7b5lJLLZ0l0tSThVyxNyepkodrfcZW1V7bFB+MQTbRZCtyp
CssGwKGRKio6p4ff2eQum310is1OL4AeKRlrmzPE3pcmmzFi7dOAa+IHFZ16
+mRL1SCHNajzmoGHyzdztOy91YIBoXwVSi0nr8hTR8VoPgPgjZa/fXKDm6HC
K8ZBarYCDlCXfMlCtUz9+YOlcOBVy6jyh62pgZZJGnhHvpIV8wzCECjn9tVi
rn8VjK4Cbwca5Lnf9Au9rGYYR2e1YUucaDUTMxQqGDuB9Cahrn+JuXFCZO9c
FWrwqBN7sHf3sRxorGiBBp5jKWsrb0tSnEI8PZMnZFx78BwJ+sQ+Vjn41Zwb
lJ0je3omlzpih2sXT1ilrGNeDLwXteNccr3G62auKuuP89iki6a8aTDEKykp
mjxxLK2ash6s/8QypSzmSVHGneWMTsNnU8C/BdBKIt1G9GILfkbcj8rA9ZwX
2TZwnAtoFiN/0fThYtRzGtskmaDG5bu2eDdWATP19ihBoeadc/MubSco+fLt
PdnriwuW+rwXwud6WuC7VfzMpBAgdqs2MQaV70003yrLfc4ef2g7xrY9uDC9
rsgfxjuS5tOaLqYAmX3+bRsEZpUrdbPc/JV+FwDqt9RipUhnusd8jBie1mM1
TEGwirE+jGSAr4Hotx5BaIqscu6KaGJuYgDIDKQwJhuaXQ9FascV4Q5pDXfe
zpdNrzEIyqjxzLCx03kqwmGGxzXgZJkoYbVXM4lwoTpc+HnX3BqgFeeNLIQX
7EGJQKbdgATNGiVHPeq8gIoZnmNFVbmE6AhCGspsh3URH8HCC7ox0NVIhyiA
jIRYTUJxfxdlBjHEZpmUioLML308HN5mgOw1FJzwClJddfd+O4apkMMbc6T4
/FovLhQWX5ZmKaKsz4xPHf2z/iDsIoTP+yPTmTt5lUedcNm6kPm92AdyyT7p
c6QGFlUP1EfLUdvl8wPHnWADu/2mYSc7ZPm0Q7ndTSVk++V/JBmhllk2dez5
Np6+97Q7JCjKenalRT9/8QmvIOMrmIvnVH/p3WBi78VHTsknqip8Y3gRoVph
n7UcUUQR+rOJn7GSX8+DO8/E9BlgAZKDqJ+h0Yrq91ww9g3hxi3dmhVBmvY4
589xHdT65KCboF21KGRVGl6zSL2Tgp9wPEB7RfyV+VepuTSFj0eqvHar0GNY
FbGw9D2nvOclD2dD3Tj6CIj7RdbWYQ1fP+Y9hJXywtX/Rcsykp/h3HIwUvSq
fgb4EtzTdG8emM1b/o5qFmdz2RPvUVfybN/7pGv74UtKJ6Fc24+7PyvbJRso
Y/Y7XM6wIt6/+/FBFUgV28vRJPn33fnzATIat9xoHJQ3rdvZz2ynmVkvdeJD
Cs3B+F6ytW9HBfDMEuQB3dy+ijUl2IL1L8ZT1bYnOxHa0/X/tAMSspuod85Z
FCIzerFmwxkAJ2kTy9rcz31DTJLTL9HMoVZtcMe1t/TN87PVLF2kbN9WOjcJ
ridBMiYKhbWGVA2O65I1rQvZoUtA7i8lRJ9HAY/oCroOotfQwOVKnw9sIMsj
LFmu1EbSVb/9+15Cm2jttBQubnNeBRBxcAIBaTrUuFivHB23FzgOfrZ0rK4L
1TSEEWKjweg6m7d2FoJCzUUcSC1rblfIPj+XNAZpyd6agZTKdhwaq8eNct/c
QcCCuouAqJqWt8ys/VR6HDTAAwSpgdRZ6fLqf2c5H89zQengooO4aVRjRZrr
NzjutHqT97D+aX3buv0LpUa6dveKVmeWpAcaEniUEtZyKw/ppKfi3/Xofp31
d18DcmdqyMn75oXaZTSas/IWnoEy1dYP5mKxL5/GqkDCBEpFonQ6lOf6DcLi
TwJaKTbuEBoi4RGZ5V/1HKpjUAzOKqDgySDFEyHaiY78rtr4EGD7v2gOdI2I
NRJqqiY08whUAPDbaU73pMSm63Q/yKzUfvvemEHCg8jwUgHtqZeqf75IO4v4
Ln2hQJskRGdomgJzjSlsNQI1mnDsVBZCptyOP2hy5onvP2bb/o+LJYkmMgiC
3XOlq3GCfOCzCTOeJpudeuhNDuDK0c213cvTuM7LsidE+XcMcXZKP9QLa54i
Dgp8eFxBYOzf5AM9eYK5Kd7EDN/n1Es6Zc4L/5LtqUOIKvYS9yZ5uU7rzFu3
ulGSbTt1+fyDB1A6vDAiJimbDu2Suc05mHxWfT6UdRVTI87X6AjKyBk3MpAP
aiVMU/XUi+9EX6uP+T6UyuzsKtVWngThNBPwdXYWTL2wlyRJBZgPc+iQP9FC
XABBnx8BN+3UaxiWFanMshWznxlH8CREa+1IRBtCRfOvKOVtBCnh3dtdtkdP
i6ccQXAOsnmpHzWaRVaUQaSO9VMX7L0+jMsKUk3pTL+i4moV3xd0bvuhRlj0
xA4KwwtkOgTfIUBUYfkhCPBHZa0cmpTutjcT7fUUt/2Aeb5/74wn6M1rakvJ
WPaNjorp5zsVO64KiWUJQkxnEgKzZjpGZibivU78eeIPE6Wgqp5WQLwPr+5f
SdSXYeGZKmX1MgabtQ6ha9iuNopUzvQN1dhoctFgXTP+eJh/SV/28xjpbzoK
xnSVYUYgAhkT79yON8WejiI9l79Od1O8O81Xvv2fSsG9h2HUnjy6bQK5Qcdq
+/GwkTEgRLsmIvVnLSrLVVnG1x3lbayqu6O4X7a04/16UoZ6nHR6t844se0R
m+uIXTcVQZ0senc2nZmZzpTjIoyeKu2sw4EqV/QIMay+EvNf8HbDMvjrI3Gq
BnjMNY/Bxlevw46ACFHmfgpMSSIdxNIHFG5xBJwto2vdy8WI+U9z5yJf+J24
o9vKT7ZW5aIQLJIgPtdlofZIfDYsjecB+zTS2xD3F5wEjvG2hTCTLkYZ/szB
fRDtT8yBqHaPd/pffvECrv1JHaSxmhkr+XcmOfXuhldy8MFot7+5DBJSTlKO
IMKwBunqm16M72838UeIFWUyt7C0Ah5C3AkK75OBlpSbcvEp8tbvrJy93qxo
c69obm3l9qj+K2S4n5qnegOiEDwdCq8HMQeHMPZTDMCpLiSjcdSj7WQJc9JR
cnyUdI8ImnMp4Ra4MEMDoNDISbsVLQeLcCSTOq7iZaOkqiL2j4mlSJZhB8D2
5YQAH6HG3skwKNXycAHotBMtXdd007hi/GCHiyhFsYvW0a/Cd6pyLiekBY3f
eaI3+W9uLeS2bpCaqpYxYrpaHrv6qisVwMVuOe0ItExWKuh4zUMxm+FGXx2E
cXoInB1QMjYxhLpgae7iztS0IhcfjMhNBJSjjV8+p+MKppS9pxJRKqTiEdfR
5NwmhGXwdkfLo8zlvGj5eJnfa9AL/+V2gsefYA39SsgxoaWZg7ghgesCFBVN
7dCaB1EhE8K1dKmKXOLx2XrFNOkFy/EMy6oxaW2FyTFgzK+kvLC6ENu7mQPM
0EEWp6hp13xsFXd4SrSUguD7uYUulNlfEqoIg+ZkHroxRBLD5JVkTrwNC9Kl
kkQOr89K75sKhd4HiFeY1XWLJb2+jeb0FS9ryOuZU6Tt+b+l2gn8Kclr7DGS
JIA5xGeHKSjIioJ7qXmC9TjFDqvtHttiA6925DQzgZS414Zrzq0NDBoVOO4I
KWremc8j0hNXbiAnsQnbMhEg3SuQdf333msjr82OkPJ61HIJ2T5XhOozFpZ8
w/6K3sr9kKEsjU9XaRMlpd/KgAjcTs1msTJwCMBI6fSReYGeUP/hwn8Y73ei
pEzMFiq13O2N4qnFY7X8yNeWjZiNrKCW1QAslfkwkCl3eR7UqhRQJeQ+2B4o
jOBh1K5q6qGyDUfDrAj+w3nYfexgMZspRdtu2okj41I4dV5xKFS7c6Q29WPv
R6Y4MC604o5LH8YUy49DUuHSvZkKIWG/XDDH/Q/gMnEVoO7i41HmvC06EHhO
kn6kXSkphhGzS4Cz4pVBl7W0t8YOwPX18YbpKoO8rvgYeWgPEf1Lijb3DbAz
aOfY6QgHjywk2qed8MIBUP4Bnb4/xEHVMkCFkob6yG1+qPr7zDczAzQh09I+
bIQg5lDij4GHDU/IqbBdd4LAIPBKjixdKWF/Xd77wDylEl7dtnaxaHP6YS8Q
aFHc+q08Xqmz51HPCOxft/BdpyWMBHv65CE4KHoAhc+UXapNdD4f6dvtZIj7
b1fcwMCfoRzqMu/9GsNqRHyiewDqJ1xpfl2ubY2X3vtQkju+u2HXrKeJDkkT
FXvXIy2GI9VikH6yXoXzIdQV343IHiy5fw5yCnHh68tDtz2uAYgc3xYC+9j5
eIxpVVcYAq5fXetUDLxwYwA15mOTxsDI2db0OMyTos1FdSYdyC0o0mHA445g
JlRFoXFrVF0ZvEQ5ZE5IJuvjy0tzannTLCHMYaNw5Kr0DWFW1ES7R1k7URSU
iJWi3B9FfKwv/PHydKvYYII0f8O/rmYB1q5AjcH17jZQ+5jBL7XUueZF1O2k
4kdc1gAMHNvBSEgBk16+7e3d2vkmJYtf1JhNiI6CIAVRUZCwi25sqP84u+WT
0O+ZytDU5TyVnePl56CwCHWTHfpAiy8dJVQax2W4S1ILkF2OJWZ80+gEOebl
xf7K4JxJZPQtqnkMUKDb04gdhN7F316JWH1NGp0XxcwqQPpmI9PdrlQ20UoV
gvNLXrMgomhskvQ+u66vWRfA/HWiHy0sMp8280TJIRatLb7hfriYTRXpk4KO
oOjSXYhR+rVWw2ulIiym5KzAv34kaNaPKm8m28TuCRT96pu7jJblHWmyQdsq
CbhZa+skgVC8uITcMIfLO5rHzOKHdEWyi20QfZY4H3mwu8VI7z/TqdoK4csu
mQvMyMTsoUYXUMR7Bv4ljbmVaP62Vyn6aigvze7XGcnUURJEd52zKZQLDP60
88S1j/3A1Prri5lBS9SDl/Md/8HpmRid7pWD7rXK/SvuC8WdRIazkVJkB0+i
N8788EQdtX1mTDsyaKOpCMTnD3eFDv0fwoEqONM9RmDo8xwA2K0IxJm1su9a
+1ZvpOQlZc1PPnX5FVyrGqB+HruQEEnpIdC1mEwxtbYJEB6rcHXYDmoFDuhn
mSQnz4G4N2MnxOpXgWKRWnN5nysd769r1/pphoOVxklCQ9kELtkjO2jIWLlX
itVHtZFMXxt35JA1UaH1TPX1a1/pWWnfsPCcXkkL1upLBiVqGVGgJCUSG12k
dciBVswKbxyxteBDv4DySOJgYDjVV01MMthUaRDDzRGIZQgkRPBa5ZgLeYtK
zx0/ILdPyGXlw6P7Dagcm3jTSFTD2YVijA2gOubhZPhProo1458Hl5XgPQPg
UM7XeAkZsu3qcScIRHm9grqAxZF7Xz2Gp/heA4Ub9oZ74Tte4a+F7IGoJsWm
IdVjUGZCjulY6EfwSjqduhQP+p2yZ/j3lqV4z/lwDyAT/2vnwjr6rL3iMpJa
/WGa8clkYQkans4viTuwA6VJThiV/cJCWSP82kOsEo8YKzCHah2z7o74S4G6
ZmmPM4dwZRHaXxWe1AXNLleddTjouDKLANL7WuYo2+kNHlcCzoq31d1ijDd3
4dpFeb7DAg91d9MxHrYqnlt4UXxrRqklGskVuvRHsZRgG2xcxffsrEpMBYbI
BiEs9UhJspMkcBxCUgK/fPVoh6ChhV7f0inXkpEILISMI2+wjf0cwlGsN17F
Fe8UR2FpABkHanZ8RZtrQg7SkMl6jU1vaZ/PpcAAwJLTSk3QEfhc8da2pq11
Y06/VOaAferoq4xTzJGkgQOxH8NIWrlqFFt6cIW6vafzHV2HO3Po5LMTppds
j81uewZDk84iqHHTXALiwj74di1KRXx98jModQduvGIJdv+PZg3gNmatnLY+
T3Xz2EqJqG+tVPgx0mm+yD+RU9vXXkO2US6dPa7jxkGVmprc44toCHLc7Wm3
9AD7gzW77RX2ZMUpexV4annlrzIerTOjBUSgTf2lbg2H0T119PpZwc0vAm5V
PKFFllDKLs1KGni2TtpkRwiGQSveRahzTAh0lgSJgV2df8HwX02g0yJAXdmE
a33b8WmIr7kdMlILWCTGO989MjgRBhF3iZ0NAisB20Y63X6axw/QIcso8DSl
mezxkIaMfMDcEynvQ5AQzYImP+ltdwsjAA1sMOXjAI+zvpOF9VqVpaw3Ml1A
pV4zoQ34H6QSfESwSsIGpf1xAO1Pu3dpeCdiwdPwviYu9Ba4CqYHeDDyz0hJ
znX/4TMQKdreBQrRouNyTogJKJiImoLKN+3fIWTA2rFGf7ihq73QrAhQJPeL
H6Sy6JXKGkGgNmSSQCGIl2xo/y9IQC79PurcBGzmTozDv2lDTDjspZzZYGQc
Zn52uB3UcY6VBD2Js6YRtdf917QCk/BzJBbyK9v90ssSUMRMUUIK9stH+rPV
B9jfcRwCMSgImkrzVqSaHM0cPRY9Eo2Z5+FHJqDU82fs5Jr1nl5ETsO9Lo0u
EumtlPEJJo8yy91yx8c1dea/+xjYTmkZgdsT3DNZNeoWnT7sHXvvc3sks4V/
4rbvqpff/Cc+z7UkGIRRhX6PI23fQCXNs3xSCs5jgEXVlFYvzS7O6o7Ym92X
XpFJNO1USKRu1E9Fwcw2/5qY6z3eqy9f0+L38L90mq0amf1Iv8FYd3xWgCaJ
e7vYoR8IlJWwUXAtNQ47VbAMlU0WYlgnvGkklYFDn24ty18TU5OJWa2u/Xp+
r25odj9+ZS6IPwWwzu+x8kfOxXn8A8+dh3mpkq0wAUoVz7vNxMqau5039G8k
Ac8kXMjbWxRIlai/j4wFsySZrq1k85N4x/3A5TkeOcKE9pV6YKcyVGz/hDde
stzO1sT0/sxQvfSAD2y0yi3qo6Ixf7lNp7AOLKqdGMCeaWRo42SKyhJU2bAf
5Scxf3kXqvotOry+hCwqHzQ6IWyYNeEvk5RfzWQBmO41ao5w03/0u5fzfLxM
EtQ5bHBn3B+jGqdSeug32mF7KKCPjveC+gkdK+0BJ2xTSYJgK4nMSxqFevC0
k2U6BgvrcIHKwIdn2UaeEKURu8K05LuuAsbtcQP84sfaILNoB5ARxp1RExGQ
2tMfqPf0rXgKGpqjq+QRatOWG77dQu5aECJvepZZkinFfXi64g3OyRAmYsKZ
fh5DOgxEm429w7wJoi1SC+aSq2q0y7G5OfkyOzzv8G70gCYAlUGWrXzORj2r
qnoLwIeIE6vaRENt+XsXfIuUoruFStQZit3c3y+pSLtHM3JZIReFnfBZYzrf
z3kNJM3ny5p7bqhxqupnXjuLesVumbVo2GM2u3T29Ql0yGWLl2yf3OSGqN2m
FupbGdPBlMzPceA18HBMGySZRjRzEKlIa9FU3c+gvut/2X+WKBjG+oo+AjJK
JPeFQBcdrPy5cYtg7Zu3zba4SGiNyk7iWLYEwcN4oUQxtCsenK+ikQHcJuIK
0BbAkaOJW8ymsYK+4IwVqsmChMva7Lm4uDnF8xZmclN+Sfo0yNDqCL9jBE2R
Immyh814WW9wHnW1YzmCWQ8i7FvYgdRzIpwBAK2U05noQPYvVbgm4pTVczDd
bkwbO2aFrhR+QxMTK/rTotgO+jPch8kIeB7EPSFWBE1jBGbLZsf5oVZ5Y/Mf
lJvGXWqPOvTGGkL86uvan5Bvuw42Mp26Rw9uRQLkAKVEX91ba3IYDNgBAd15
AVh+2RZYmC/bl+Ogmvxd12mSDNdWtA2N+bf3YalfxBMU1F8yJMYDww/OsPSQ
DpazHXhJV1E9sDpnizZHgWunwyeusSxCT7xzbZQQgs6xm9NBKB6sFCauuc/U
dhuztGRPvmroAV+ac9DJyGwCKy5kajg9FWxJaeprfiKDQaIPpWp7FIeDFSIu
pR19v/43dq9TwyUbmVVxHdfCPiYOO3id0MhYYc6xkvGAgjIayCJfIEn54AMV
Z98+igZfOz8VQFv7T9FZZqXh0fa9FkaQYJi6FIhyf7eEzFFMYl+FddT9610D
CFR0FTi90ddQZZlyx7Tll7oJ0kyeHd9NNF8Dp2NIZwYaC3jGNsf6OZsgYG3V
1idLlkzJU5rR/mH2P294EMvmUY0wo8uScqoqt+YMwNdAFuzd9KvHOSNe7uSW
X9wxOZPqMoHLPTX2UFPLCMSNNOxdzlNNolBnhocLkVUR+wOC8d60XN0IUe9q
LDTSF0ZKr/K0z4WKNYQEDDwtWWmPwTS7lbVsVTifoxXv4myIGp2L0wEPHbb5
zOi5RLwZd6jqO5v+/TJaLd2zOovig4OxVAwxzUESxa2+jffkUte+sVCI4KVC
16osfQWyFED2Hu3zPSV4LzROxeoSTfqWl5cqrUYxohMfqG4is2u8yn+GtKwV
uwheSUXcJEZA2dOJAUD80v3dXkayUwYNWqY2OKz9RCYgUn1muSV4n3c2JUxj
N0bMiB3yLxJUh00YJCKo4DbLd9po4kfUC4f/8TZkOnRI5zC6sm7J20Goqyby
7L/y2cQiYroutiuYUZGAdkjfFW0wgbGHUgWHjWJUEPer24G7yCZu6vsY60Eo
7nyLydVNieEr4uYfEABYlg/eSPTb0KLtqfy9v3SesLw0UfEkiJmcpKGyUTAS
ckwmMz1D5T3+8LKJ6ASWTg7TUrMlleHABpLE+jam2Plb2rik/2ppRnLIIHjl
bXOkoYYKPG4Gj5YJ+h2GJDT5UNOxXcGEweACa1sKECkPAngu5HyvqC1EOru4
6ZNcvANTBEAxz14w5xyZ4mpV2Mdl4jJJ8oA9nVOVMeVAdf97MauQlvXVCu/r
oOa4iIMVwRIitxoh8iHuuOp45gTrxJ2a52NyQ7TnAEja7iH619V+GZUcUeM8
R0aJcYuETltbCItwWH5EmLWM6pWdKe5aX5lIBI0f4JOxg83d3kTZf+AkwugS
sbUEQocwhIijCG2N+UH/diptsyVwEZIXCWngklWti0GYhdEDlEZ4zTjJ44Gc
ihxRCSK8Sqc1D4uZi3zp/mb1WW5JpWLkwzxGYCoyAKHfYZapAECdHNH/An/c
pEo62RYpRZmQOqOwLEd7AHQi/JvIvAws6iE+LRDOxpwnR2d0/8IUP4u0g1gc
9hDQlCllquIZyxfClJhPXGvcLtC3nR9leo8L+UnIhLZOlVk43fF/27e1cNmt
KhSO5eOOE+9hgsRskaaf7mIdQd/Yk2ixPB4udfjxZfCKGH0TJwflTqQEqAP4
Vw9jU7hAwHAuWvAGsUYK/GRA3gfxcPByF+l9fffSQQfp+9IdP43IMu3szbgh
HA3a73UybT/GpK4+OS8np3+tMtqjOQMXwDqZVk3S9WSK7YK4o/4KdyxWKsM4
XomJ379hRdZur//7sIOtqa6y8ubMkY3WMwvfcO+EXh4Unf4XwLwfSnvflvJS
n2aRZASmCWtiL61QacoflArbzkevyyv87BzbP7DEt3VbLc/PV5p8Gx65yQ6E
RikWnNlWlxLDG4PNihcHCktjTSIe3N4Rd5dqlRsSO/9MdMA08R/oS/mRLJIF
YgGN3DM+zrcb/hVotUP6E1m+t1FdnC20NlGHwxUa5jjAedesa3sAEF9JrvK+
K3o/rqWtFg0rs1ZIU9Xsh2CNp1hKz7SCLUNHNbTc4E3WmRTfaKapoiBcWypz
KiDNEAer2OOVmMvjzeH9TT3ig1n5LP3kGCKtPaX0QI/c1R5MDSKM2A1Du9r4
i5EcQ/GyFa5oojGZtAHGx6oiD7icothszs0WYZZN0MrAAB7Gphjvta3vGB2E
/sQclX/ZPnluDi6DHmAx7E86tWiFfy3FCkKm8ieZPVtfMOltuPrMd574gkzu
wM9pvLVIZAwRoXtDkPm9RK5K+RC2x2O0S+mUhiFKf5/6qnSjIlOpimBaWVtd
p/9BCkQCzQslorbfqJwAJrsSgaditNIkST4h22iHmt2rBr4NWmQIDhdcJVrb
fWQXLp19LzgKWyMrg0z/pYWGbLbK7t4Hl4befipr53sGTLhFKJyZ2hpzVSH7
NRlxIj4WygU3XlzXoJzJUJ6i6EElatzUFYvmfzKjQ3McvAzIn0GQA/wt01DH
h9r5pw5vUUAwYdcCIKBbeWNRQ7irFUtQJsz7jsZO48aC41M2E7AkrXwIrkj9
jIr/nNNNZYONC7qgCGdlC8EZvf+J6OGKyO0z4doTSTqKoFDsfnWdfbdSbNR4
unhozAAghiwuEoB1m/L1ondO082kN75b5Wb8SROTX6DsRZsvg5+3K4Rq12Lc
9PO3zg09iCdZJDG5+Ripnyx6Kg6wv9/oGrM/Mm1RbQ4t8h7SD4ZFeN4oqfGt
AuAaFYw1gRaRr+KJLXAcOZTxZ53WkYViJFKDGmxfKmAfnhOlzrbBgK1aQ+0g
ZXeYYGMSKsVj8MXlSs4IM48LeV8vCDrDhQJS9jzF87BrEv5pvXbDNbKPA6nu
atOsdwYAY6E3wKn8bPyFHA2zSdj89RYjbfT+yrzzyIDbhG52L+M79cq/Re7F
4EWip7aHqqoEYH3FCNVAWIW/Nfo7FW/3ev1pqaZnc+3gBzVfqSCu7r8nLaJ8
CynwF818+D5h7So6wOhRqAdN7Umu4PQxdQ8uVWMiFgnu72XRuGxUJ3/1p5Wc
JJrZrqtLSWFS7KkBN6H507RmoF37rRkGm0yEsg+sngD9SNowedNFaHl7PNM6
3XbixRT8/94QUzAYe2bgFgbOohiUWisIIG1rdWJq+7owCPLNjg+Vvz0uFUmD
Z04mQnvhZKaBdbHtfniVrhOqRJH3ckjpSPYtLMy710lI0PDeBQB5/r02vQ82
NRzzYLIbiLJxj6b+ZC/vkg89h9DtJJv60hnTHYppCR5dNWdndLiJz+X5MHdc
/h+UwE4z0g7IQkae5sbs+xCr+LWKul9vYtOsgEzfMMhmmUyw1qvTbSvvtIAm
H7XkJWAnLDUrm8tP3TLMLwfoFI87nRdhtPniXbFtacexRH6sb1NG0VMCo8hk
gmbVL18WuEeKCTjJha8ZnEzlBlBwbsvAmozaj/PiKT4DQaVomZyvlp7qCVJj
bO5VIoIyo8Og5VmUqfEg46LTjrZ+5EOM/GrcfHxLLm03fsNjgB69C/jo+tLN
pZkgaakp4op/0j1dD4EMdpRPody9+2hd6zI7ElxYGt1TfogV558cddTBGMhI
UreM5zZqn8jZ040W4qqEJhfLqhvFfJ+K2iwl7R1aMB+3XAYVxTErLnbrgV9T
umxJcVg8yVcNSBUD19H48yyjF9lYIbLPZcqiaSmTYhQW1hwb+3y2BpC4rmtV
fUbwUbcA5lzZfoH1IaOJVPOCHpOdVUEox/6mNJUd2m9iYAQu/ejKe4GvHLQ1
99OB2Ukxc03WqQgcyUyf6/XyI6vaZcIUfFTOhNgBaa6qCfg4+afJX3883Xtn
oF6DLQaZ26M4XE3vfV2hublQEtkZbXeZaiA+IGxWVAWor+MKi9hWoV6xvIWF
az7phUogBCOqxXOLCxw5ZVMZH+E7KgGW9i8WZFtSUJLQrkbovjwGxcvweUHU
7E4GNm6z5Z3Bv7aMwxlFomPAWSXw34nFlP0mqYzO48LU/z9mX1fA6InqTWKB
9+7vEQEvIIthiJX8iSGAQpxzyRv33PGh4ReE/gEifUy/MEZ3+zlEns5d17mt
E11dUQfl2LJ3TyJaLCQ9Kw5gtLyW4DYNYH7jnVwTnhWXCh2GAkEQwurzn/jZ
UE4u4VsjK4h1TKx/n5HyTUih+RvAz6Wi3tcGP6MNcHN1a0eMSSj/DsJnEA9U
ueH9zFuJOH3/RoenDBX1XMFxnDok1ARzSP9Qw2iySSMDNwzWk9IaXiEIFPR9
hQH2/T/oj/D0kMjRhzWRJZNISFdq/omcIG2/Kk1OdYtPIom3FDbJX1K1nODF
URF149JdjIUIeSREg+FWvzQmr4gJx6p9U/lDejvKywbkOh2hpHJ8GnwVP5Fi
OO/Maw1PrJRN2vPDVSjsptyPF6qmi/dR1xjbCtr9os7iyIlIJg7w7SiTgzPW
vRyyA4cQq9NmsxnvDyf1ydP4LdIgveT57uXo59FqsjoyVouWICljiGBntaq9
16K111lRyBeBv+URkeIW1ztj9F6Doxb15qQBNR6Qy3JeWkZ4UsObM7oae8UL
kXmh2vdNWwmKI/UYKjmnKWHIPmOFK3OjbaVqc9IIVKVrVWD8RBXGBWupNntY
gISmtPA6DmIM59K+5YURitIFKSenZaMrPB36/v5ycjF11AeMqf6sB0/LUNwR
Rmwme20qVQ3/PgxA9lp5tdi9DSVqxswEDL0+rfKuoVifUp7dZL/Ej7rUvny1
ekaUNFUM4Bm43S75TyXZZB+FP7zCfBFNMtxg8LZiXVbfBgxSmKdw0r6zmoM7
LcZ2aDp4cAVozjywtuLtzOo52q3spK/J9PPKM0Zjf6g6A3R7JMHupLpsmk/B
mhJ9J739ae0YTRM1TjKI9E8idF3BBvli54QHHQiM2SAZqlZK1U7fLHhXyhcn
dMm7w57RZZVdTBDPz9uQo4zMdrpsh6fKZyqAltoljrCgDrP/W2WY0Df3fM9P
22elRLgLrh7TINcOeJ0PDSoD13Un4R5Fn2uctdyskR7glO5IKTQz7zJfydFP
0+oxlMSGE61zGa4Ia8wviJ9L+ne6d8L5P1Vin4c465IMgKRCGrqZ2y1ZWlbC
SdUvXIg103rRTW0/LG17llzS5/M8zN0Wv5vglBVrunn7PlgM0fGC6oghFb/K
6euVyFTdWC4XtHQnW+irBkitW6fYRSaUMUI9pr14VFEM9Svo/hHDs184sHxO
3P4kLv+mUUNTAn0q/aF1kXgl+4gfe0KfGU+wWXazzMK8E17QNNGd6WSgjflN
c+2b+bCBmWNR/dxXRSe0Yc6EAv1eliChxcd60HVQkvKVwiqpj8zQ2IIO20nK
7gQKdZP8JZd4eXlt9m2N1byDTmkfGU23D+ifKJ91Q8qvuDeLnhnTZLvh7z06
iMN7LIv47AiFIS2GPPRrnT51uLtFDs9v2s2kSgL7M5b1AF0jE/S/TLG5yQVH
sGJ4X0TtZbGCsKMfvHFPszIUM6vdUyqECE9bqpLAwm3DGg88z8f/UJgGBKtc
/slLSJyK0kCkPv6nxNak//tBevvWvQq0Rn0PupUejWQ4yP67dZMIpvM4YeN9
UOB/yFGljPznsNvucs2F8XwzWLucM/xsxi99di435lzrRTkrIIQgp3k7NVcR
oAkLc8HAiuTr5PaaaJrZXDXyXH0UBhw2ooFPflaYp6K5c90PkENtoVVaTyqg
uTUlhrVI0TT0PlNy8e/ofqgo0aWJD3f45iaaOy7rALCWCmq0WDxpPH3jGaEH
nuuNqQJXWwM+B4rp1+EVlqh2v+3rBl1m8xO8s/51vP0nwCZo9L/dJ68OQqf0
gUW2jLGG5+teX+pAx7rTSj7d4Ns4ClhkL9M6Emkz9F55MjBL/xqWDNc8Vlm8
tRyqSHf6vnRio1oXKFapXTQ0VYTxwkr4CTXruITdwEFvGvZe5tVXCe7I5/R3
fFW4M/7q1Gr2cMMznkWyKjOlWIdRloaQS76ENjPSvjwf1rbERSjxEYLRM0s9
N7o78gG63hA2eOUqtUBLvapAXOL6DlEiHlmdTg9Hw1Y94un3P0ejLEfv5pfx
sCDuiRb+ysHuig5xeXE2RJht/0N7EXAHqrxv33GpYasPtAg4cKFk7kN62k4u
G4jWGu4fdBrbLAyg96iDKQbK7Ed9sGkWmX6VYfK+b6S2yRPMcGJi2NbybWIv
JQr3WzV78QyA1D2kJsOh1jm6lqObOpdNbvyh+gVwlRZWwKs+iiExP/i4Ut/M
o4RMsoIirC/s2tt7E484yEyvoG6k52OV6uNzhpr+m4sEvClgIzJgWzNI4Tam
XtRTB5D4iWL3GgiHdaj+l9Dx5vuMY4vCoqeR5nMwlsSE2pdQ5zpjRGUUnWAE
9B4JxM+SY7cOak4F4Q+T3cIoQnr3FK/guYCG5EMPF6W0h6KkojMSBR6Av3jD
nTyVT2Mdnn6Out83NItG122ZfyaSVr3+ORbQvtCmJlYEtveImCTeYbSQ5TaR
QrMwpt2N6K1jZNeglVDujC+zQNRafGAy6O/TjC1rHMIV4Eg8aPHPD8WOO/dx
8MLzZft505COdI09+CuqDj0iDEhEuRrkawI4DlFepUqP3fyAjchHsNwjk8yU
22A060ulJUgSWsZqtdP+96HSrIfmjWwIrZu9r/m0gE0a59Zetytgvyfl0ja1
32PVrfFzwvZX+4zb/SW+X8p4RgRlhVMEppo6EmShUronf8ORlJ4apg+Ia/9/
xKyEuMdnQwH9St/uYZFl7SzioTMIDcps91rYw5ZASauoaVKhZo+B+jamqHQN
LEaT8iAZJCKr1gs/YJGzSShih0spbdn0LvPB+HsoW9YFbLPJkKz82o0k28nK
rHZSIW925fJiDk67hxRKwrQ/ELwEl8wEcRQH8mtatJhE+0ncp2ef6efEl+cn
pWed5Kci/zp/zKWf9H/fTT5VNy79q7f9qI3cA6Nxi1IIEQ77his6e8K0j5IB
4Hmo9y9Dy+mRmaGXFOMWDlGIi+oqBqcEnEuxFnsXEJdA6U523s48LePrJibo
Xfyj8AaaIIbwySlsbLxLsOWvwDtvd1v9NeCzFmtvPBGrsScPROC2xodvA2lC
1euXTmj7MOeOvtTaEx1XLZYBeDi5Odsv+P4WB+/SuW/9q1vlstV8jAiWrG9A
8r4Kfbt6aCAOqdbUC1Au1BgSkqy3+P0afVctRwSHl5l9kL44uaHbag4iSIxL
qFpcspuinV5NOmv3Lp0We8wGpkOk9y+JL7EpLzrbDvAgXLXRLWX2xE+fOxuY
sNem+Mn6WTDUdMZgjB2jyIK32gjY6wMYypbBJvV+oKcLmMZkMG+Ydm7cXUCa
FEn7dEY+nud2Lz8v1+JpWJty3EVF4n3y6c/qFaAnC1Ksfdit5fB5zcnn36uk
jOPKYJtrh9BChDtNKCiPrKVMN+WXbC64ilwhduttA/ZLwxbaze13pCMREkhm
WC7vurXBOymcIeedDvkID6yxb6t63MzU2HbRrXRSN599iMBcd56zS05UkGYc
Je3r4QoTD8E1L9fUGjcx8jA1TBl/xTbJ6wujXwI3VJc+DNHm3hzhUp9pxwhf
7WTLGIMGJqjbS8g5A11122g2pKyqV9rmMU8Z+2D5Xp3Lsxew5ZONfFROj5MU
bCniKxYisbe4Soje3pujSIWW9U2XT9Tfew1E9Iq5aXiiLUPS0YKw+xg43lwA
+GWyum12u4umbX+cX0DrCiTLLrNIiO0ly8z09jxP+21B3+6jsGD8a35RK2Y2
s/IbYMq3mPolfUBrdCdzL7wFb2RCziAJyuM36w5V4dtK1d+ZndFJRiIlb+6d
Yv3gs/0jiz6pDTEN00x2hpoR2b7HEuK+X0jQjqOZMQGT2HUXzfJdNROHinMZ
/qX6/5NpGI616j0J/WqJAe/neVIkV3awwupyJXFC9sFLc6SXLK58uSYQvec3
YA6R+pye5FhWOok2L/rlAerwJXTZ6FjUoQc3H9C+rW4KGzw0JVz7TfKijrDD
Oz6PWf7M/CiHZ6YBUOzOSArZtnaIadKM8L5hza9Cy5WwF5++B/Ye1AqUaiUA
bQ8Pe6v7RabNP3P31vUEnt0HnCPp+TMkQX4TBTdWWTWTAej8xE9lnIZ2JMkX
sFXf2iT9AgVezmzs3tSBHCyiakCZbBTPIMw8ll/mKMBkpfSPatukK/NLCN0d
8TlTShMmFHRTuMCO7+Nk/pzRdxkjnlZJj0Qi0qkG5fzA+JtB8WtqYCPs3rVf
uEVryzprrdieBv3Cxz4erS3d6+EY30Z+MkB6UWwytL6LazDOB5ZgnuJ3+rmO
73W6K3cybSAXTLjIHCrNU2XQ7lpfngSQiIO8CdiFcagSfGwgyFkhi5HvFJUG
5/amriONcBKRLSTJbWwPp0WJICxgAebPTztNtOLU51ymwr1JNYikXEb5W4Qu
aRCp2TtNn2kxgRWDT0yefAMpLoZzlU2bWJ0hogIX5PmXcr9GfVNvwH/pbuAj
ZmOn995P68dbYJoGO0BjdK+WsRa4HiBevPxgNILHygtjnabpzx1Rry4nQYqZ
0BHU5SAjh8peByfDaLsrAyXQaz6uuMdGcgPKntPNr1qM4EWJDpKBU1p9KJue
5Eq9ZJqLt/2LZSjQG8YIMVYr46DWrGhGFZBsfUdFV0SIwwTJNkRCHeJH4/dE
ueC1IHCQ9TDKn48ExNY6oHCR905/5UCGtKNYYmtk677xCvVJNlZaPfIJ1Hv0
2qfSk/2J478r6W5a7AO0g2+rogtZYxT1n+fwtzwzbo3hfBEVcsDxfDS4e2A8
A2ENIklWcB4PXQD85wuGipTLr/c25hwWOiMJj3iE7tQuMnLtvWyp5g8yXdmX
SWK4E2ATqOAf2Kj2H+BNVYoPvd31U+7TCdd7sCQA1nSsDjBZHmn2jdeId7h5
rF9FhFI7whHFe11RNlhsaejctZ/u3KFrtOYtL8uuLSgGTvOlGcsJwfODvHmi
D5fgwFHPPdPAo1UbRfLdrK+HELIP5OwLgkISc/920ZMtBpFG10ihyNu2kh0W
/1beXVHBl4ooDWRwS+Yg4GAPygcTSgZAQX1vdgaSY0FQF1Gz4Io1N5ZZwQLy
hdoibm4E3B/3UO75Xixu2hIfqfb/QnIDsu7dX0QCEVJVHyX63oHPKbnKfQuO
fGapJx5EGslIWwF0p2SpblFUgL6JR8kVU9S3W2oBtpJ8seS20tmLdKHPGn8/
nCihvMF+veaVrlrHDxfJJPGdA7cnvzIy1z6sAOMEKR518i/FjX8BTWLUSr6e
OMFyeVJ46pGu1yDKthKee3qOQsZx9tsTIunLzzf4udjm70iFDyk6LBHlzw+7
gF4OLLgDfpYk67uihSUjZ/0VMN5MpjcYOBYKv/AXGOgFw1NYM1zNKXwy3NOQ
9a1+xlFYubwTiC7kYf1CFjs2e3UzONEvmXAfvpuybGnJtW+4SkhHdsD+O9K7
ruZmTFl1b48vLL0ONO+7Ogd8BUqTm36OqpNCdUsGItWJX/5brq0kWO/UKXlq
R4BMaLLH5hv1zrBj1BfWp/Z0WbWwqRCToCpS8L9i46gfTS/hO7M1VT2sch3Z
0ptcpYRMylSNjLDc6L/GDRXKsxrQ8GWpYZumZT6btHIy8rmfKrLeq1GGksaS
7nQi++frxbGICyFAp7yI3rfMR4zP82L45ll9sJQWDJgZiSE/CctCpMPALlgs
PVS4xJ2x3PAez/tBxLVmP2pewabcWrpggXMXRSvz88o3DqUpLd7or/xO4GG3
gOVp4Jwjx5kjVqzus3+PoSTbRk/gK8/b61lce++sK/FpL/1/tJ4D0gzjWNeQ
z9P//YkVMeRcDMxQQtSvnJPYfJwdOgfAqJuRmFB+gljtvIwpLgJuexeY8DN2
LzgJVypFKFIJUbeE3WgBroXdNjSNm29/wlKLksiN0002NB5+JadUhfNpGnKc
Gqcdb8mX816iEFXN4Oth4uz2LH2gQvOpaDrgvG+Jm3m11Kqo9TY4fzpXVWz4
iSpOZf9rzTuYhF5ee8BH05Sp8aiarZPHXFLvlQ8JAMjzNBMaOE0+KyOdDAnz
ypzEwgGKioydg2UFhpiV5ZwqB3n1ikxax/hqBcAgQ+jiNtYvMRkOFOhrcirN
kGipnSx6VakuosRbgZzAfzW00KuDX8gO2yCPeNqkg8LzUYBhHsLQOSaVu00x
ywyoROYlMrdxcVznDpORgCU+CljPHjlCdCJbK0yo7VtrhD/coMEmZf1D5NpU
SUBsgUkUqC/J6lf5V0XzjME8YySt1xI1d0fPFdc7q/G0VmYUdG4OngqfbejM
mRkR2ut8dgyVLO+++2du5BMsJVENSt+X7JHWJ3KSnKXmFRkW4cszhj5rX5en
GFNGFyo17LhaClAWmYD2+/li5QqsxfJ+cWLIQVN/Gyz2DIbxA81utpVrTUeN
M9CcBHr/MABj/DA9Qs9E2rCkba05FQ23eBpeIPqfnIZYRn0j4DG22mJyVLVZ
cS3xrtihIpbB2MMJwCFk9jGOghfwDKByQ3YRQlHkzbqViqdNLPVWZlTD/1nK
trgSohsGuM2pVBBSGU/fnedJnGvm6urr+oig7wxFUGTA93J/FaKfZAzsAvLQ
OPLh8QftRshlJIeKCnNtmX5X7FvZONClUz+zqTZ5mTLYa+7dcRFL1QQ3NmtM
c9lEQzAP1pKoq80JcXoN4TnSTf7dYNHH+bslXjUi0ObuXWgxuY1JX7Zzg4Xr
HDa7WMpqk5mTJnKSbqy3eYD/R1ZCqr5s65KnOW5yYBikW0JexJLzOK1zfKhf
/Aea/G0WNZ9+o3dyRwgxDhtcDaFzHCnnLutg392dySw57z0uR6TVAYsjOtdV
Jt9N7PsQ6ZD/lInhhFhIBT0Aafb2gb6j20EqrXWTF4S5iJCqcWqn0zUBXtqg
C+e3yaEH6XyeLIumHWPS9l22xtYlPC+gO3GHZ2+JUa9rUtxc10+9LAc3SLJw
YQvy2mGT9D2QDtVKaoq5z0N3BVUvxZSKY7QbQz3zQWhNT5+bArWLNZRmJWmH
eF+HoEuszIc9R56e6SJFNOTsvNxsu4np13jf3KY60RVOI3pdcsPCrrclq2VO
OdD42WHeqxHLMm8PutXaHrKV+WuV/ijzH6hNHbAYU4lvUI+TYgyZXkz3OIE9
KVvfYue1sztl4IEW7fvBn7I0f1hCzigtuE3OxjLB2pwY5mBho05Se/2VbyUH
xaPCFleolwbz8lDEtaCdB5q7ru3uno9zxCRE2/QB89PSIcItgFZ4t/4/abNk
mvm1NPRvZa3hblZvWurVO3kASfoiudmf0AF4DnSNJLePzgNYT8x1Qlkbyhnj
Donhoqj6XdY1UwPQvg0KY6K1aeDnwzG0KK3GG1JQDzF1J4lsQYY29USErt92
Qbs8NAwF63muxkP9T++A64Z9CaxFdt/OwcLDrpXNJkvpSt3hct1C6ykgvTv3
fnqMHII9FC3oCfhHs4VTUQKhl7ud9gxJSTpKRxMHdqL3qzObD6x+9ofaYTwF
Bi9miDlxDp/nCLMppLBtSsvy5nsuI7Q+wzoFc6PLkKAYi3OiwuX4HN+4jB2v
DE5DaXrA2IfBauXcosUxyW19dY5mcU14JB5JB5tv03+TqzwiVSEQfxuM9g9Q
0xu9T/T8wg8SqPR7h5zuCUoj2SRiyeTH1pJ3egJcnW00MeNRbIjrDdEO1LmK
Hl4JN/kXI+6XJQpxioHgH7kkqFtoZZuFNeiCohT/HtRqaCHXszVahwgKDSpT
aR8TXGqE8PPLFs/MUZ0K/dpBLdJwblQ9brvW+L9rWTjxtk1nsD35uorWRQZ+
8RyWr+om6FTF6NvAQ4WifONSdZSqUAO17KqRKAcJj9CS3M31XrpsafsU8rmL
M5mgG8l4PoQ0EzZ2U4usXFolqR+ZNO0St90hJt52wC/e0OUineHgOR6sTswa
7wpZ5UMagQqGsPjQcW6ak7YY7F2ccOO+08xlZcztqfIgQkE6IrmQE49DfZlh
VJ8RnGXwSSxQ6Sd71kgQNzMzK8x6gY/W2CJgNDPDg6QH1oxp+9fAHliNe1ZC
JqS+Mh/d3Ij/OgIrURPqldaTSsNte+53kOGxe4JqzMErYrZf6eWKP6/bBs1H
CI/6ZABXRom8jmIUv7j2qqZfaz1v4jHmS006K/4CuShcjOvNdPrjYT6enxfQ
FJeeNRD8+655pO2asyG1UQ1I5d60wwxLBe67RBNYFzf3IuGO2ZSiInJzr2kC
rXAf9MYhlmr4OW0UCdM0ThOKle2qHFvk9q8Y6OgrdOhKVFW/lmRC6Po49Gqz
o4aFASaYSGb+2x46jFfhu1znTdTHhuGBpx/3NismiVtyKZIUXL2LM0uU20S5
URx+s+OHrW54ID6aFSjezyBpPBRWZXaV/19oDejMr1cGwc6WjWWGvgyFvx/P
rdONZqMg5ba5XAnkCYbOCKPS7iD9SJXbU5WXJoaTK9rGgC8bfTdZLjO8QS4a
F0gBVwj3n4SDg0guomNpOAf8LwOs3F5rJ2npt0P0MafSH2e3VWiT2BM+aiHz
6YbATYy/wq6EL7URLWT5kyv0oUz0MJ0Aych0hCWdBHdzPE4uolMJf5z7sO6r
bAsvqtADt0X6yPZGTwfXLRSP2b1V/d1whMSLvBpnyWmPDVoKGeJjVUhsTXiF
lZmccCeS0pm4/zPcWlkwbpYzRJTgC0bXzBoreVm2X7iv51PLSHtSXs5G3kLi
SsyKpUtzytbKLZc7cr0yqETxPgzQZFz7W2RvnDfdkVhPGtzZPVjV3fynUf7t
xCkreEoV8fBBfsu4mleloWMAa+41QzydcI2UVsIz9+Xpvj3HZ7yuomaMD56h
G5t6j+V06j6MOu06/43lQrVXOV2GFCBiPo05MohrDu8NXFSmc9v1GzNBuXd6
Sh3icKO7lUfH4nUgdHcixgQs44Bh975JHBLDjQuJlMUSblpULsECxAVdQN+p
5ivSBp7Sb6Bxi7l9lXeuFCbNp3jxL+t5fIyovGZaVmIgfhFD30xlpXmsZZFF
YiDmEAe4vjWKhA1cWlcLqwoonHIk141ikJs0HXqu8xHLpdGiBqmevah31GWW
Mm7OOCmVxe2sYza3YgKsVqUAT8hNxZfu8FqS4QV3zceLojrUO1e45Cw/f238
kYf258HJUWYJRSmFpvPc7g3oRcD2Gglu4aN+38T1tcCEqDWxkDQhdjIURtu6
SUzCFThUy1kQxlOlQujcAp5qnQMvi7lHfG3tFoX6NycigpIGdlIxMi2FTNMw
RJtR80ImK9vAZu6w+DZBR7GaorUVD76PWoBPAd9kDjZfi+NNPPBVD689ADKe
nH232Nm7A+w7Zy1ZZ2RiP6cGT18TN9/dgeXyfk8jot81/mjh4s9G/MdRKp+A
diiT1VDEUtF26chEkEob9+X1nO9o5+urkF9h3MzP7aJ3THahgLmkiHCyFOg2
e7udTnStyOjKq8dwrKCggic/dtXmsqtxJCMQdrFV8U87PjEGT4h4APIpEqde
NhmjEmQjuMgkvdjndDMvAQ54jpiST1isfTicwKWDAC7bSQGhhIUx9yzAMm7Q
C3sMKQRKs8Uh0tGZItnlGbx1DrUyz7umusPdgAdJ9LzrDC/MhGMRkfbVfap1
4AH2GNN5syVzdDzx9/b2B1I6WovTmkq/BC3Nq5xcE3rF7ndvDLmgtBjK2pDg
QAZSGrAcKVs4CGu41wZTZUUzIXwrFAVXxlHVs2RUX2h0IqHHDWA2lZBmvijY
gx1jq39u7Gu0vXWllmxoD687TgdBCsKDKFmcDAx3pz+1KgeyPFk7Tlbzsncq
5/tvNCbW9jlVMTFz1w1EFyokJI+TfrTS6F04mDrpu++iZgBQdmJT8IENYP2p
B4/jD84habXc9hlvpZx9emaTB3cPjZNkJEkPAq0K8KYEUFvPhcKCHjqeFT8Z
EmwAq59zFPkc8Uvvm6evaE4rjuGJTb5WuV6F+F+2Gd5oBa9Prn4GpG8bc7gp
Uy77GJCxSTN1VQDA4Mgsb86LJpIiX3JezUQ1m71w9SN7PAwiEy4/x31zF9G9
CSAK+w8jSJ/fKnzGj3jqM/XyP+oxutgQnLo3wE7YOJ9BhERpD9RDtK7jPGES
SDOi+Fv6LZF66HgGYgdn2fHb34giyVbyh1c4kd7w/g13Nu2RoUDC8iLgWGrP
lJ/73xKG0lpPbyiAKj+9vNWKngegZLJivnzk9WoJs0ookp9EcywQlwx5CExz
9nBKAj0LIviCEmlSdqcqelRPYQ8kNlIHU/yqBn7QvHeeWPKD2VYx5xtxe5kt
r9Bs1bOstLXsPfMtRUopMcFY/yKX4NyoCGNbUW1g1beuWdJl9vNF4j2/0dFN
sSEvsuNaPnn9TJxz/gmrTzpR9UWh4J7IIMxOZBVMLVdYjHZemdEb4Z2Hb3sp
Mm/0sJZ8POh9ooxIscnz8ivmyiCWMdDPIgL34hLi5K9zu1fR4FD3uO4AO0IQ
GlErLSPPvFDA0jRMKSu0rZ58qIbqE4Th+7NlXumclm/QFnXL5H+mK29TKxvc
VfugW44B9Xo67XFP064i08WWt800VOeI8OuGk0vqjUqpc9XhtA2tcZU8bNYk
uMNfAbAjHTAHLXlIbJdMA0x8+qAiIBCrampZuG/4520rA5jSaZvq4tbC9+sX
wkeKw5cm7WRv+P5+jlE5vsvhyB8KqGdIEiHoUS0lG94T/+QJyDxxJRK1E3C3
zNGhFB2lXhF/YQ6XjsXmOZSfsSQxqtQ3CJ2N0zPQkAMfAL0SDhJe8lojzTCh
3k0Hlt/D60AaPk8hXMToJ8eXH/piDdi2uORx4p3LHexyCd62GJmBSW2053Y/
5ldBtPJBhK37TeqcjyszfJYex5eLASZWm2ZSIMhf2HDSDy0KsySLBIkS+eqw
Aen1nNd6CuAu8dB62qRjfcBY8KPbELNljEHO17ZBB7KoSdgfPhY/ddBSA5AS
315XfWkMbiOKHfMRLbMvOMnYl7oiuvLAZj2/STcTOklDTQ8ivYP/sJq2PUwu
I6Ff6/+unIvtLzNRunQLPbJ52Vycn4/XZmLYKnpRMttcZavXEp3eVLG7OEN8
MHJN90DXAYyPCXPCdWobxo4JhiXYYb9g3vZIE0cJOs2GFrlhAkYqg0sWwKLa
HW4Aygx1Y4plrepFD0BAZfXZPzMdYJE46I3v2txq2F/Xpo5Tbj+6dTuNVD2F
9Cwh2Jd7WDdxXwJeyMHsFMRhC/fS6+0mXTqXonfdUscx11alQ0fsPJrbKS/b
wAkDrAmnk3ozblsysGwpvzxHuU23cn154n6m8LNawwZbVkfZPwy/Xe0NthSE
W5IovtWBZt8US+A7y2pfrKkLSpxVgXKEsAS9ZxIugw/luKd7fzKucbrgBMue
om01OTe3qerbK4gsXBx+VitCgbMyROWyrFLiK4ZKn7DJITXtPDcAS9qCQOj5
BQzF05V/4Iolycuysy4sUIVv2sq19NsYZUNUeoRn6zEAzgqOLa+SR1XRHA7F
juwnin5S7aiyMHgLH9i3KmMU+ool3smgYI64nARt4DbarkQIfgCwM+1hUwqd
R80W4unkFEVp5vW9Di1XImvPvOLY41qqXedJuRk09U/aI3Z8DXuCyKQet8aD
nf0KIaaeyqrlA0FYdhZCTeBntY2FtTIboAZI8TQMAqHpLNzLrz/OT4eGYn7b
A+TktmSnFrroGNnn0T/JTmnj2NWFz9sRMGYOYRe1Zrw7GaOCk1HCpm74GbQz
i+rv/lpYzbegOMIUgmVFVsRI7TbODn/AnLfHD/OJ2imkc2P2nHpo2QGBnHxR
j+rbJp29gsCUKsd25oZkgzWvc/jfsv43AUgaJ/3gcB6wz+xwQcZya6fs2s1V
EmY25OEBTcQl2Xa6ugtigkZL0RqBAJGagIJyq8frn2ebn0B73PZK2XntGu2U
fsuqxwnvsWPqSwdbljrqf4zPXbw7NOp5NduZYhOAjsfUCEBv4u4l1jPX4qjH
L8Uv4wzKc0gMvCczuIc4jqcv6zZwioFmc7Gb0efL1haBseXdDv2xTZx4lssR
lGAKto27fHLac515ckJFRCPQ+F8E0sj+0BO/hCxWKx958LlgdgB3htghrAo9
FjPQFpiU/gbsrr+z6U6GsexQEUTm4/47AYx4qZEYUFyw4aiy3a1rGJz8+qsG
dnGZfBZmovFQiW7MNrmsK+v78ZWikbdA1bMlsnmYGn6zOoay65OK3zBx3nuT
ahL+C35SYWvSNdHPvUZIaOXZw5vJWwjhZr0Nt0oYuUoKKuXjOzv2tb0lMz+O
VR+LflLwyuI7TrHruFwVvL+w9iEw9hRw0lxsHYE1TAuacNjdYT/ace/8Kewl
lr1YU4l1jyE9I5J/n5Yg3buvvFrdxUeVTeGrun15RUk8tX/9NfQ78TfXOVar
dQLcMPibgIG213IxeymHU3Sz4TzwRraJAHQzGIQW5w4R0a/qgujuUwE5N8if
SwuM5KNPd60SHRGS/p39FOyTcyd/hMWYfSlAIL25LS47037MXPsBc8DF7LPK
SnhJoTdl1FQcuChtJN6Z17m2s7kJYvJdX61t+R+vaxoi3sy+Avn40PFgnKI1
aunqi96Ov6HJlb+o5o3tiMobYJSPuILL291TKVTOsX6GtWwGArpEhHo9GPlI
bp/8HPN0kIrndl4LnE56rYbLS3zY2DtSOTnCJcPFB5Oyv/JYtv2kL0CEU8dM
+W3ixb8nU3kUkhFdoveUuvKbw20lM+fCjpxgowMzPo8tYf5I1F/TG3v1qMP2
qloSeRXn15fLXBE3Y2k1oX3w6iLbgPmQLuj2Tn5d2sisW4Y2+MQtGyJg8OXy
inujL2F0tLNGnsF8bRVKOtYd24VulQhuypQzfQOc7t0abu2+/of+TJ5irex7
u6qRmKgfCkeRfliEduV8a9YNPWJ0hksN9ttkPA99XnLXlRXH0S2TTuBr4hjC
p3W6oKQ385Mmgv7eCTKPygJXi9BO5XiTLWC13kLq8LkBVgmBkvhc2FPuQhKN
jsglZh4tJWXnt3eS82E/2R7yo9inMmHu6WiFOll1WOynTUUNlXILydFMZKXQ
b76yQD79SAAj4/+AN8eaf8kNJHjdnwd3j4AhOh4+SkkGFQCAsCa92jAdvohl
z21/mu+SyYYvDQabTHSxHMQpQ3ryhSyh8XsB5AW9Dt2PVoXqr16+2eB5FNwF
bm2OXg1vN5h9B+R0nZwdwmyfjODRCufPilxysD4rcENn+iGiRnyizhdiJz9o
TeJYTJ+HLU1F5Ff/tqiSLF9vWm16aBLQVOAO4C5Rqu9QVnDEg1C72Kj6Yg7C
VucrqbF30G5zhcMQkkK68npM+vdekZlCfSmq05j86MEgWiDPQxnvSHhVhZgE
CzEdjYrx2pMBf5wbwqRvVLypPMwkvrBWU0SCiNFhZdNQBukvwXb8AGmeVqbg
JjbKmNK/vYdCRABkEjpOk1ioFB58waOYAbBq85YSRCN3pTJgC6TrUpEEIgJd
cnpJ3LN2MKqLU3VEHW4IFKhYBfp3ygYTf5Qa7fHy3UQ6WrG+tmugIQ1Y6Gr+
asXrOa5wdMmZTqdlsC8nzp2HCHj/Z75J/vdypJ47BjzWiMRHaX7LAb3v7LIb
6yE4mQSb+VtNZJGi4Xxwjq/AFcd0KjmSn0I0pzIm5KViw3tY8TctYvp5u7Ql
qH/VrI2yZcplzvKcr6fdCPyqX34USYTRrbinJnqZZ5TXbwF007Y9cJjbxhN6
DYIxEZpZx1E2s8PZtcB+4Y0fM3+ayAx9TMYGcfSZoBLyDnd13eQzLZ97K9By
yUHUu8HmBAXFUP5N9RpBPXiHRf2cvVU05cEjakQoktS6GSifBcVLy2wUVIh+
t45tQsizOF0iNMCLRI3aytEy84xp85O1eMxSEfFoCU/ycvMBqWeChh0Wodc3
Kktf0KZHvUZindrF5N4CfGb+7+fkke9nMLkP2rIMEX3WaDIoHzDZ44/mCd24
a6LRFNFp73siWDNCf0jmwUs5sIFvyotwodmItKqHiBeEgFCsjn9wNFld6/54
oQj+DFJalXIimaLGSAWS9KTxUocArUe04qSYFgTGjVx9dnDMtAqhIWJ2sfYA
7D3SB4sQDIwuLoJlqvqPWD8Ir3PNbhvYTBtWNXkPX2OApgg98I+nahkcxEJQ
HIhs+BSpxFcZC93p4i8WCHiCqznDfHZpOtyRUJOiCEiisXbZXfMVcJ9eiDlM
zkwCN+KKtddr4Ofqemad0k9mpGPf58xWsd2IPWeKaKxsbqdiWk01T/VPhFrn
OOaZHaMJD5L9AYw6OrpOvn6H71qkKTKrNfD0SApyM/Y7QQ6gW9wqo7otNIYh
r4+cnDA5PBY5dGI3w3r72hnUavM4OLvy5smaRnM7b6myRuZNHjL/OCQlQnHl
1+vMRulBcohnDG5eR1ha3tku/D9dbrTqIK59W5eIV1Lqsdm8MIlFiGrB7N89
geSLYrVPFkf/afQo5JyAW0F9Zoigb89nKYjjndMbNCLWr0l7TtMeDdwZp/uS
16SvF3Fg0IGSlqefWSuwMhXKTtEiVbRLdZakhp3RNelHk6ZMuE4X8AbP8Sw6
fLFVyx6Z4eg9Yeo6WCJy2NTDlhOLozoE0eSCZPbXKTAtzz7yBQdMEhYHyV83
q1vklajX0bc+ERsGpd63glU7abkwL4uvLW9cSa/wEAxNqqxyywtHUP5C3NGt
txuR3UiqttgJ4I4KpvpGRn5ZSvJVrgvr+9flaKcG7M6P6NCEnQYoWIDa+ZYK
ank/HWQObXN/XooJRGueoTwGIIbVZw8IRb1cPJv64vN3ePYgh+7YhESvJkqR
SLfE6ykf7Y4tVD+cqz5S5hTSxr3vUy07Trnz5hLTbb4aorfH3VkMIKXUl1ik
K8G68vlQFsN8nyNErDBAMEaIkOAFwB59hPW64+0EMm0RiNN6qHLoGJRYkNBD
u1xEjjHyJMdZRFjDk9L8ub8Wk1YkW46JfrVcRseuNE5IRMJ72w8CHina4cNt
X4fpLXZageNAtrNVCh2RfI/qVn86BDlK3t2Hk9RsIMRl8f6y30S5Yjrgj14S
G3qpyu8c9cIJ9klDHBAbMznM4/6tkubQx7Dqr7HdQlnlQ3y3z+wCzt2nEprY
7hUscogWgIgPons3E8KlL3ZlplMuMzkv50MNDhgRBHP1JKP7hbBY5yk3qaGf
jyFuFrNul+9QqrZMmxAEmBqRJD3moRbOSJDK/maqtSBEaPWe1U0PBOIOdZ2e
INHmBcOxuEOOfUyWFIWUZXCQG9VvvqWr/v+KVjqkfJ+s0F255N/hvo3uefBG
jZ6Ythk1pSOCevsEOVS98KQXxzFU3OZ4K9lZrnDNjYpXZpZrOhxjSSj3vR66
eQ+huXjbnZ8v0jp004aQqiqU2Ow/K60n7TkFh5fPM+EOR8rB8VdLm4kLyrrB
VJ1163/DwOh8X0LGlnYcdA1nZW7+Zl77i+WlhLN+DG1ub1GtLV67UH3xEKP6
1O6458HqidtotMsu8C9jzMmMLcKHPYDmHsEcmWdKK8FGz7jaGiiucIjDzOb+
HmMJabPg6sashdCciHQ2XgTKv4n5MNUTPZYH6NGNN1cfxU7mlv2LPGBw2xtc
IHuh4lWaoP3kcncU76JzvcgpIGdiHyc2qol0cx7ZLpcN2ry1J4Yi0AC+1f7l
8PhyDonQnMugbsiR6DzvBb4is//zgw10+FmVoXoSwBpOXHDR+Bvq3tgCnOqE
Ns0GM+UAQox0W+zCMv+H7tB8+MZ5TZuqyiIp1EieZZOAQVSVpJgqiMDmYC5O
gw8oSrlcIr8AUIDmuRm+NlAOUuLQwvUXGxnv7WXPxN5yk3TLVmp6MYGTTbSE
q9sIuGDdhMVoiTW0iYUFoIQS94bI8mCSLeDq/ypl3SiSUmRSeuxaQ+kfSRIL
yYUlxYydqNIoTdoNpRU1T7tJTujgtQk6odKYYGtGpsLYEGB4v/C4suZ/6JjA
sviglbyqmRAInYa3CmmZ6DWuuXKANdVxVKuXFWMnlOwxS2t4ieFs46XvVT65
ZzM+gly6RVGZejxLisLVzs6VPeltLpxBfOLLrFjZc00n3hrvh2TE+Xy2XMBc
4lhrwZ1rU+IUyxqFU+PYqEEEaIKlso8iLLmgpu78+J4U9LsSIGmA7F5aVkdv
ytNPEpv+BWBNOX0E1G1T8kgTbqpu+hiAHB76yb7IPD1s+F+arDq16zfttRVj
W1WTDby/PLrZf5gFHBedYAzgnEATUuWcOlDLP2e2R12GFIKiqaVTWnW2Gk1K
zkKShAOmbpW0/aoDSydACueQGJyarSoU01C48vKvKWbQYOAm9S9liH3daW6G
NOxP+aX9g3Ovk4qifAUvT9PnWB6+l4/IVbohRIICyP/M/MbBa6NeCf0/MyjC
SJwBczKym+VDDwOq+O4piASoa+9sR3u8Ld47zclzQRlFfgNUckwpfw8P6HXA
hFMOJbMGXzJgMIYzUcbrkQ5Do/JO9l1LVdqkrGPJDmatG72zu+ZZIC/o3z1u
t+rO/9cZchWzGcuZP0zXXpFA5dE+zLPwfQqSyd0IzORvvGiQd3lrNds8lpwH
aMuQypYBTP5fRuhqokOKsZrZ5A/baN/hGXbH9q1oqAHxsrX7b08ARANCFcqh
Uz7OQAzTNwuOdf0SDMclHQnPct0TRzbxrURVOlTMtpxzsZcj93AL1Ah9FzPq
0PQZ91K3TMKA6MDpRNWRqtewyHmW0zdugVYQ+U7tvAIwX4G0OoZ6ipXIfG3D
1fMDJ/q0o+qf4D+Ses06GrBSP3bFT/kXEaTcxs+rXZVyop25lSc6YA/Id5ld
1yS81cPHg21Q5bFiG+XcC1VAwoMx7a8Wf4HmKiXnKF3o+8YoZvG+1q5tU8dv
gMMN+i4vdPN5A9DCzVfLiFGdeX+GaigbS+BReZoQSIRV17bzpnbxUvU/2kZG
dx8pzm2AnpKOozLwb/x6wPAA9LoBvsEBqQCMt092DShxOLd6JkOEg+ujvsna
cyGet3Gz51cHZXNeA7nZ1y2Vx9/LksMc1NenYQxmwWfgDEJXJKc/BX86FM17
r/jYJZ2rbsEY3FRRqRC2T/YmOxc8XbSTX21fG+FR2GjGlOabEoLwZFsJ25ZV
LJIJ5NRJZUh78tb9DmjTR84lJiIJQoE8USbjAbxlxe4l3A6QrkbbWm/xBIdj
IUM7xzRqvHyUIGg1ESTRQbfu8okl0sEhw2aL9yiVZWwnxHXVdIyb6A1wcFnX
UZzRyADf3nz5M9O0Cdw9BB9eVxb4dBXVc8HVcnBXtscRaEjS1fmam3v+fjRV
Gr+ccrrzwAbWzdhJqVXwnVvoOL+sidkIKQCNR+FZOXwOI82Krm0uWVMXI8yC
TTRBR9FUN3B3MmdfqLISILZt+lLbJeVd+xOBai74RyjHwjccQb7pPUc9ZdOx
Jv7xR2+RGrPTH4FGgXWPQHk1G9MjzlpzlF8Vtekyv0z641Rz98L+mLC1PJrV
Uf+oJ4FsT7Ib+e+hfgGydPTxLVW3hv/cjYMGzh4IdizdmjxBlId9UrpwTxlc
U54myhjKsOSB6zPhcez4wmSPp6xLLPLsZb+Wgdo2s6kds7gTYEhj+lS4LEFF
zluXkToVAfff654aQPDgQcqyKgzpEjhxaQcVCTArNpWSvPqQLVwPgsrwSrKX
2Hu4OdpO+XFtDuWQYVPDJ4yxzRdYfUhHi9DWJ2N7fzxecjMwrAEWkT8Gq8ce
cvrwtMe5uHBfNEyzPP0ROwY72gobW7XFWH9ODi02WUQKbClpcucFfEwx4Pv2
nA9N9pMubpc6+bXljeuEILULrzk+RrU0cyQdD0s92o3ubqUfL+TwOmo/OUtU
mCQZ1g6w6JDhXQ1DW9H9uvcFRuFhb3Jy2/PWeYi6bwbx9CtysIdF3ZfSIeP3
Rj/w2oGrnCMTWT1TuHVy1qHwqlFMe/9NKY66Js89QySoWVQtVhboWeGXPHOM
ZoNxTCu9I2hsycS38dXcMULVQnKpRdu2TrElhhV1smZgnaJmeYBpgTYUjJWI
liQJM7mI/XsZmOxj0J6H5kFIp4IQxvtlpbATojprcyHiNGZ38xeOHa3evHqZ
euI3dAskgYqL1rv/mC2AxS18KwgDZTHHdVqDpeDDvKuYRJEQbsQVkmvkbxy4
lw/DqO9Wne1K2kpro8Qhhek791byGT4VrxdPHR294HbSA0veawTgKeivbdiB
BK1E49H0WJFKL/073vFgvspT7rvdhBEPM9BC2rEhIFQRjTM86mLBs16j0Zdf
xFbcrkA8Vw+fT26cLhT2A5FMKcH9QntUL512geBKzAumV2lf/O631G4ibwlB
PiGt3roC1C6YNks6XK8IrmnSLdUhywxFn7u2jLIlmW8Gdp9dH458Nx21/Dzt
GE4b6aV2uBVLn2n288nm2BOYP/ECBOyoWNWseFgVuexcaH+ORp43+iywE4U8
f0u4C4+Imh9NP088dHYtc5/nQVDoU7PAXqeaUSgudcWOjhXYWEcCqnT6Koaw
jAmcxEt4b1AvUZqOkm2NoSh4PxqSiNN11PfI/FlWF2OEccTNDgPVoQ89jwfQ
HO6nVzuavQaKqpbsrNlUoNfJKGcemz83LpkL7RNjkUrQ8Oq0yiFy4sMaab6O
B3MG7JnkzMGhH5a1zjHeKjOXf4Kv8csBTHy7V9YpyeKY/zgRSZSibe7lH5nU
QCtZ8oZZ+6owYFwKulS4fNhA2NAgxcXxf4fB0kemHc5OiTr5zXyjsr1nLH4D
53zsgwrls8ZAZ/1Ut/xuY2r9wQj4FZOg4RBYFYD8JethrdquC4Td8slpUeoH
JKQNgOOz8m9k9NETR7gVQp2SlX6i20DY/WHTDZkLJeDrBGgOSM3D0LzehVHa
2CbNq8Mrty6cfzN0CToUrEZ1dFxclTOcell9Xh+1IMrRrpbj4IXN05yFi6/0
f6FxlRvGQdDLk2IhHGd09GudHPPbtA+yAO85PF5V+EdxYG5wwB1gAQP2BwwM
FUCuhdhBpMCz3qErSbp4c1RcxSMj6YHmuyAqVwEV77l+bKvYl7KCa08jWrcc
vnz4VqzxNtD1/uCPnu6hmxOc2NJbYQBuYT62H6PRA7i5DmvL1yfpL++dpMj7
tfeDdEpT40ESFajgQCWdkjdmCJ6qJzAp1h6MNCP/edgFtTLgHLXtv+4wH76C
CoGMNpsB/yTkjzfFarzwqO/1Y3tzF5btG1VIF5lv5LavelBW9XJudsyjKeLD
14i5Q8bv6//LBWQ7DJ6mQo9NyAO+PTWoQnY/r9jV3ccsgcC5wAiqY0D0gga6
+uLCR5xdmbcTFl3bycVQmdy4w0MscUyNDvCb2RRKS/B5PJgPmJghdVX18zKd
4kP6+HaE6OLjD9dHynxPJm1QEt1eClhTqghMl/dIgpuJp+N/2Y+puVJW6HWA
KdXjWb8KafYSd82dCcTqMHih1TPbSVGKWqDsEvinHlpcNPUB5Pr13ZbcDqik
FUWrt3tNPslXTU35OWvMyfnC/OP9GwLu2UK19mQ1MsCAdf3GYynUhKpMrbOT
dEifa6cN7qpMl40DRecTB6fWudw7+yL5wapZIrwztKIjNXCkkgDpVnD07kdu
Eol2928NfqfRcGYX2CiZIGVoTAMz2m582S4kB1i/9qVYpJ1WNlEwADbkeJpO
b6IRYnokTjNx2dCf1Aj25y/H01iWlgKKF879LThho04Kkk6+x0VESSjPShtP
xy2ozznohrJL9VJiLw64adaD5dtFpQPnIcmyBHu0KVOYAZDMSHbwLad0jXja
0nebuiKmcKrLAblDvJ5DfNaIFZ0htCBd4R2U5UvM16T/rClYopgYviwyEliY
10bOpv6R/+QWMwhztEFB1ZzpOjUBzbenvCyxN8XeO97C7cxaxufLxYoc6tEw
z0dyJxMPpobG+3yIyPO33k4rnBU6q02q3eQwTaVyNu/OfD4ZI88/Aau2bM9k
ZW7hajPLufVQ3cBZhbKEi7NFrHOta+wL1Y+QswWSHPpWrwZfQL/y28tnUcEC
4swlL0Fiw72m7UbSMk5r1CJN8wlKmYsVZVAhEovNfJ4OUkreW7LC7QCwyYgD
Ini3/oNYPBf5KZN1Qg0h5iTkdIY8aIVFpCuzY6J3+JKoDVZJ/T6dDGV5Mxce
y4gb6ZaaJuFhjjvO6qTSyExZMImSPmzXaB++6Pp+qZR2yWuKAQ8+GSBweDl9
QJ/2QSpYudSeZiJWaf9te/4vJEpVmdGVoCK6HMhKRBHky9oPS4GXMd7bKH9G
0B06j93HrNf0KpYMaplMw9zuSJqaDWzTaaP383uVJVkxsU5bp0mxqe036et1
bb5F/B6sv24OUWSCVAYCFI/xbCVG11x+d/NJD03fP6jR3+X6sjofXshVnRK6
h0vBkLXRJqVhYZGNoKroJM3c1S6IMQorRcWJJY+KOFc3fiUAr5vdiBTJWkfE
8FZcE+PIkXl/EcTN79auqc2rO2aZnM85ccs71m7nmUiMyhA/Hlgt1YzLyXmx
w0g5pI4WoCQuArNj9uCUiSh/D0Hx/dZbFECIg8fxuKZ6xYegrQSkKo6H+cTk
mEXJjmvJ5PiiUDBevCXaXeUM7XfdbtoMbdtstBhuSFgW1DycfPo9Frhbp78M
ejr+ocZ4rQx1PHtunMYbcU3ASOCEZI9ncBqQ0G6EZXFnyq2NxOPGragwA8cl
70thhNjIGO1cQGiIXeZD796rdPEu177ty2bGLz9JmSWJRjgXPwTLicwwU/Gm
Zf7r2LRzyZd7/Rt843xFCuPvS9QwJWmAcn0YIYLETripNXABZGX+Yww6kT+F
bGxWxle6U+JzUrMrFXCYQQwPCYzrk798WfwqWDDnLxeR+pu3K4z4uHIr9XCQ
fCUsMqCgaTSp63IaxiUD7ikqcNUgWi+L8Yb5BbyIlsef+xyQzJ46IPFI26Wo
yLisxAAuKvUzB3WlAT17DyhvpBTxMqliR2epJh2uVPoroT/scObHYPDTiJv+
uCyFWowfAQaF3q17Lp+DC84ndt7jk+u5ugvAt5p2bK4zcTHfAiB21mXbM3YM
ISvCnVf8TScw53GbXLppNcDPAzAzeHU+tdvIkKXFpkHy4rJgWDjSggxWvwk5
rmHvK8OSimArztjC2CQT/f7GFe+deQw36v/By8fh6q7ra/F1IBlq8U1y6RxJ
YfQXIVIL5PEIsxPVOzaaQBKOGkBTbmGOiJZ6hxpm9eqEEvCVuWSUJpfqq3PG
D5IBpet8hf0obSd6ThLSqje66RUpdEjNm+p/w5d4A2XLgkEepNIqt30O1Xn6
XxEE3VnUT6Li5d6BsMI02u32CI8v6o+olXG2VBB3f9TTic5t5Z22oOgeOk/E
/f73r+86eu0Giq2x09qXZJE2e4/UsmIQ5w/76hbmTmNf72IFmZQLvzrd2sgb
AWQVSCKOv/+ssrAESmLTAo9CI2WHKy/NNwd3lM9PsKnLjnqGzA7Y2eFcCNRw
S+MJpJAqohrEfiFoXE+A3rZ8u6IAbY7QgUiQLggchVPzQ9T42YBGIuul2nqe
o3/VVAqrJVxrKiMoAwnfoMFeocMaT/IGeVz00Ryrv6fRJkxxROuFXbyFRdIy
V5gsWwutf8gksQSNqrAjb6Qo/yEyCwKCftoKEjCIzt8feh/T/V0VebLd1LlV
qd0qug5B7vP2P4YTlQdzOT2D7dwEOvA/XFyo2m8AZyFoTX6NeO7sOeAtxZLP
I/3Hfmbd2eQrldXJuxq75XfvOWXQUbvf7B43VPmyJ93ihNSRamDojrY+YAGC
vbK6Sf67JS2cHJLxSIV7VTKmoFhBa2rhM8LgFZhfD0UpiSv7TsDR66NbqhHq
lccu1GGJ4ZppgyUGVCUULMv2xtDWKZCcpum3WcoXUi3daQe7sikgicmCpnRg
4gkhFcvysmhz2ZzrQl419Jq8HwrXWHr5RB5YZR7zX53xOa6tvI6Mamo4ZnMA
4/320+vTNXFEu/9aMOb3mUMdgI8hMwgQgwV/Y7zbh+wW0ahApz/+43T9xJZg
WcPeurGxTwCInYeQdXgrjuxzuTX59KCV4OxVvL9F3nqhc/+p0b91aVdY+9h3
VqSDqOsEFks6/8FjtvkUo56no/lB5zWNhW7NTaylTzJEZ33w581SWmsJv0Qi
fTOSVKFNdmr39HDrDEQWviKNhaa+sa4wRVVr0S6FY84voiswOCXLOc0uJVG8
jxH1FnN/rzJcCjQ+gGZYIs2Kpve4ofLMtxPdW88LEzUs8SSsYqUNOefrSf6r
dtwyffM0N2rkt5Tq+my9nZGmixUotUVzkshyAV2eJKj5qL+jDxG38Dnr1Erf
wc+sQg3cVcyRciVO9zY/+bbynvndlOOwN8iPCPe3deL2aX+p5UwcSW7oSy71
troVWM7ETJWLmwxZ8cpKk6yiAhYsI+YVIju8O6VatWuLDqtB5W8xij9bPhvv
iGTTcKW39V5felarIwoSrWR6Z/9uHPlV6F6eZJnjgQ35/K9yXDS/3si53hoF
xEVQ+O1bheQ230cFc+k5NoV8GVcQ1DTeilgYMfg+p102iPX1o0ROHyYX43ea
ZbGArfxjxRPQC0dBuvpqsf6tTDHcR6pQv5j36edJEfGPG0wEQaKOsFf47kxv
XEhwfztt6lKTkE0TIX7gVbb5xvJxPNBaNx4ljrQzUgkctRckL8cpY8EIi0BG
5QGRTIboEgdNnYrkbdbVhG4K04brXO0YiBx2esiHEFbWtseFp4aXMYCjHP2T
2w03WTnZHT7stkZGljIJ0r0NDjwzdQDiAWfHoQa6Iaf7wKQxeCbvUEfXmcyU
Byta07e16pHDsLg/IRk7L0RUALuW5zoSzRyO30DSZM2Z4afs9t/UhMeNyCds
JZUUxWJ2hX58OvYHBgH7KxJRBQAI6OS3hbOiiSJZi6T0pgx0eagA0LTp2s++
nacBx7fdEhv5BR3zAupfzP9A1WpMeR69ZV+BZOp8KW10elQFKNmfTZbKK6aL
8xTssTo1aZduewO2tmKAKeqROhsOO41bBJyvuRQDbhw6+H/guvPRIDG372hE
8b6UCYAf7U0rjH1LuP499lYq2Y5CQhLVUwMlRTz3VGpRAASJoQiJ+miKNym7
uVoO3dDbY8PDaX5zAaPbjKusq2pro3ZiaZ+rg5xkc074oTuLUrPUZV7DSTmF
k4a9sZqTwK6hUKB3zT0wsEjBk2vOgoIDPdN/cyjIi5jYNz9WYUQFYwUiahuU
ovkZxMglbvWJM7zwV1gm5Z8Jb1B4CeToLsgaPo2bH+JX0XTxutq+1eYT7C0I
KN28imrcAVuyujx5dSNZlkOX09ahASUWeCPhXF/1VPfof05Uk2/tA4uG4RNl
1A9gA975NWdQZ36jJRFs9JPTeGLRjrcuLpSKjgu2iDhrDY2rxI52APje9wBL
Qo/j2N1orKjFqFBlaIkj5XGl36AOLGTcJWzWjq5NwKUuqgnr0PyAQIKos0Ca
RvDPetp169V7e3NyTDNK/BDYBD+Jn7vthQ1axV1yXtJrSaEWDc5pqRC/m/Ch
jL8PvSPMF/XHtGeTM+0EO3ncgsiGsyqj4wYdvRSy3S6NHH6Hi3uQ539aGz01
QQQIlOcwaUki9VnDPJYgM/gNhtcjNUL1+uIg1LPJBC6k+qE8bFH0vs71MPU0
KAvjV+8Ep286r8kDqAGOOJjKED7+UTx7RGYVKXD60Z6uwqPJibVydOP6ov2n
b/6e9B2TK5xLY7dFa10QDX/wbczzSS8vMOtul09lAGubOZKqgp2QrUTIOBE0
KLB6IDfYmUwmKquLMxGpg1hO16evmjUb1ICVfEnh8KZPpYhEGmuY3STMARLK
5X3TQFDV2O80XY9VHwx6lx9H9okJJvWKYRHCx3BXQs1CPrZ8j9e6EYimth+o
8v2dnipuz8YdB+zZrGdJcCgrOME4NnhjT3QHSiW1gsni/R1zUnhtLiDVKhA/
3yWONMyQ4pIRXq22ye61H6G4QXwckRm9mEjeAjakrBILHtJjEskoHlGHdd9o
1aVgU6kqY1UerR/VC64TIbKs3NmkEPOz9JzfwfthC1rbER/4KHWRECiW8klx
fVvscK5FPGhAYlsxitEffmshvm/x38qgd3rxhLke47z/OFJAmUrCeQAH8O5V
xY+DVew0oqv1BW+LZslLk3PEGmdoFoxf/u16YZ4ISsu8gFTmpQDf5zEYBZKJ
2XKF22XG8CCqt6MAs84/f04PoxeYUdF0BN898Hyzu7A8gS2R/N8kiN4L3YLs
6Vjm2DeulDoanhnYHXCBCBgLul7xj+BPDa98UYI4Sk7YujpwZ/wsGKQUSg1o
9MU0lP5u/2kar17kwMsNLB0a1U4syhZBEd5j5HmpveSaQMsqanqV0fW1xGM4
mgOPHDPGv2Va8sBepvKubffSHjmlsqWf2fD/CdaM1bNhgc/H8f8Wrurl/N08
PlsUHt82iiIXUSgQy39UCl7con3uFCMFBbtgQZ5RXTSdeNFjS4au3oEqmDgr
3/SXsyaAt7BSRK60ZmeQYOZfgB3rS7M0gxPzdbcLPKdo9+y2gTFvZhBEyCmc
4nqzgNv0FcUTCyaE16aSikZz9MF64p4k2zKmLMx8dR7FZZLGBJHbODXWG1Qb
ahxq6OXoozeeAsrasu+KQ9wpT3wtWk70VD1viwjaXRG3gg8gEmdIOBg0WS7b
mrKlzsMDY8T3iydfEFWFwC065GTWX74lfRBNZKpbBVbLgzWfpNj8A9Y6nUDP
EE0qmq9mQR4UWv2kufrWMOrM2vpS/ohv8b5Z1hAMdz6buYQN9NfEScRBTBSQ
moAhwaX4SLrY9nvyPZzSxPbl/FThfzL4eeScVZ9h4iuVX4c307/Iaqf+NVKg
IYAoBCCyVVTOVBGdufSa/xftWyH2hSb5a2IGeL7uTZuA1gocK/ulmCYNmxD3
INcKpKrlGsCCdEp0VS6lz6ZWUsD2rJkLUOmgRScXpzjZrak+/V/q5ugUr1zW
PvEu4NzGG71ah6Qlbwy/0dwqMRerAJ944C1s7gBR0QVIFbze4GarvrjTKchg
6B/gzsyzgXf8ZihSFTRXVTUjVbAp5DVPKLmEWM067SYeI2/0ULzf/AAyH8V/
sji9zLoBQd75Jj09JHmA5fm8JwdtUJ/fK/Df+4hhMMq+sDA+qb/Eoh5niHR+
zPWdImmGdTTtAuo4N8WOYz0/cBZpKRkpw+OKVKbzUSQlv1YQbudix09dwtji
Qz9Wmp+J8lohQGQUcRbVLzzAVQhdfdj8+uKo+arqQ/1jKooZVR75endWwkcm
8QFaZGVW8FjxCzBIgdeOI9GFMumk+KNTt9A6Qjjrnud1H69+JcIypcspX3PA
0VmyyuPPmgdqZ96Z0CtqgLx/jxaw6TsiRgJ3IasdOqQExo5b6vu1hZHDnxwL
rSn1JgMsxVebBP5WeuTImMNpysFcIQdsuQlptPyObN+Fuaf+PVVTy6znVPl0
1TOvBon6vFoGM4+rAU0Di68gc+oV/rSj/OrJBLWWwXj1rGe1pvNYHkBhg1uz
JhQezjf0QK2QKrGEEY1+xtr6BkojS3OP68CTfev7KaTK0cP0f/BLNeT7k+Z4
3Ga2GJKRLTAthwjyiQHU7ANxq1suP3lJrkY6PVLK463Sm+FA255TbCreoJ7G
M5L15TF2tByaKO4ewgHPTeP5d9WDTfsTyJLSYz1HEFEGVWlJrcYYA9LNaU9R
uBvpYnNnS6ZYhMPeflT3i5xOyfH+J4VukL8P8y6pRdjsWDO3eqrh6T0OSOg1
nqf7+UeZUPdfOUuHgTHWp//oHzNdusMhE5e6dBZDZKwdiXzfRDTzp1bhhLXD
EAjQeIqbIxJzINZDWGxbSmDUBDRURl0pceZifVdKb0s/QFUttl9bqVn4m6b8
qFdvlQwF5sjKxSwyNit6Sd+Et0ZpcluEq1p0KHeEYenU8poMZh5959nZgQP9
T5YOAc/KPAYkZU98QZMw6bTlATSWKDnopp8iJ/EyKMfoQxFVWbbW5z8zyXpE
SnZdT6c9aMIsskeehuYf0vMIIP09fJe/Nu7u/zO/3ok2NzdNpur8TrgnSdNU
IaQkUVpNxK8/uGqQeXkxNV8Uib+/KtBOH/rzAyStMJ0TwKbhAv4L78itaG6/
iEEP8Ms8z2cTwVK4BhkPEf0TdVmAaJSqz4U7JQVLSU956BB8DEa1lfVHzH8D
0/f6oISGflSuMNqAatqCt68kEFuDpmtRqyawqZurIj6qbQ3isGExpQWAvZc2
FFqwiii9PE4mVXJcuXDuAeEQeGYtwAnvt4BgHNOS9ivJWhdn3ew7/UhqIAP/
ekUwWLN/xT3NDWbsfd8/xHnfZ+Ls8+IwFwipEkA34dt56fPHRlXdVN4R/wJI
h9fbW+RcqTiisPo51iP4E4hVFsqE0UduCX9Zr87dV7FwMGShrtEND/aOB8wz
aH4q4DDLGXetmozvuNvnovZCWIIiM/o4RV7ZRcVS8XX3Eyo4cdpObzhWpANP
2ubqFc92tMb6X0OgSoiupXHVNf3FDpiVAZA/DnOPv8XSvSrw0zuEzjKSZOk9
IWQocU3J8xUfcPj5BTMa0xUxBtNjF47Mpv7iUMvfiuZrls7l/6NvSvrd6Axd
3g7uVrsz1tQnDBj2NHvagENuhKtAOgwXuXGBLBLdb2zQOecPZ6bSMFZy2Bya
XE1lwCJIQlXFtSBk9DpVE3KnidsGrG9ZRZiZinrBo9kIf2q4/AAdXfaHDTwI
pXLxIv45+HBraMcZUcwFhpyz2v0+yjCxRarh/7Z2KOD9l6TqtPQer2Y8DCSq
yXDxqIOnEJTup05IXZ968C9ppFa/hRasoItrGxMaJnFsZQwdWWTIj1q5winN
yViWLVaaBUJ1ds907cS4pqxNWTvZ0r4KiMK2bbvSmqbi3v29fHBbFffZ/uuK
Ts68bgGXWcCeWTTuTgAuMYcoA3IxynotoHPuM6cXqn9bOlqLQEKFw1MCUBk7
O9MoK/f3ykIRQFfNBS35qjXLKV5RmxGm9WJ+2704a/QpNV+sN3reSqRExBlG
/RF3TBLhZOPa2kvFG9ibwYHWJ308uEs228t8fXduH0fjcLe0/RMFpThwguoH
7pqu6F2XxhTSSZIyHbUEFKA16NydLP1O2r+QpTRBuIPLzIFYrcJ4KZDbeA/4
timdfef3qXxxF+WhZ+24WvckB8JdH7Iuwq30EM3qU99BMYUxTzInuwv/Uw1n
6kVQIVDLN1wOuVB3O8IjhXXVqsn1g13uRe4PFbnpmFKL2a0B/6LJcUfOvB6l
ISiXRN4PjwAt8NpPXYajFuvoh9xWcxs4MLYvFv8JqxtNkhZCt9USZdafIqAA
+7/TBnzOjOGayU+KH1xoZ3H60tZdLSWkfTqqQnqhDMF6wg0NDAFW0/mDCl1W
KfmfIw16lJDLxbjth/Zp2yJoEEpJFzfckNEptRsRF3eAstb0CUQaL0wRNyrs
sA+JIceGBci/I3uHkH78nUTHjIH7Spczs5w7evtxv6r51YrY8O6R4f9NgojK
fzKfkZO/S3EadVYMzvtqOWAzPNRHq4q9OpzdRrHJbdgXwZ7n9s10gYeVHCyL
7ASPRrm09XLcS6nBRZ3dqjwwE5Sxt4ILAuvr+wh2hUlacV+I1S2COdllp/oX
0odgIfSIlXnZXNs6jsTfNHlgy5a8kr9PSnkWwQ1VPYFroKgpGXmIx18Jyyrf
3QqvWp4JOeoCSq4DjrrINN4a0FZpazVT4hcll1Zk/JC6EqJ/teMlwxrnVMbZ
qcgkxli5AiQZyX1hEqVH42CB6nGj0wyuNC6sYibYWYb2qKdd0szCl89GWXL1
UYU//TNvYwRUb9/J8VAO3TutFpl8D38WDnS3qPhTcLw+aqqPUAPdaWAZMo7u
9OictREmG3Xt9MRTIao7L5zJYQuxdIwMbCURIUMdYzZj6hIaI9mCq99ybc8w
vjBC1mOVb3O1dECpvwFSOtE/BzQy5J04p0dUlUsb8ApxeowL6jwJ/ZGDcgre
lPGmYkLYlNYcPGsecQfD6KPUCAEFX5VDqziJ/BJBU3s76T09/12dTpkHtWqF
huwrXkp7DPif3LL/lv+EHGO11rZEw/637NHI/6Asle1ap6UYcXzBb6w3PScv
5s177b0lhXLykOFAq+u9o7pfAGLDGkb5gqldnerrqpslja9X7JEcYSIpZnQi
7+KhVLgF3CvqCwuMsCiGu7dn4KUn3wvUa7D2ZmZtg3/TYlFU8nsUE0fu3qqi
uRmP6yemOzZiwum+GSH5YUhzs2wWxbBaicgPF0Rx+vNcAViud37iY3688gmO
85sXhCP7rNKA+4BeA1iMsSoATrG1ALyqg5IaDLMcuNQ/qpvSOsMh6aOMBMh9
BOec5bphJzsAKLC183QzFGX9Wh1NU/kHfghHzc7sOYsmo4bYGZoGgFphIbDe
qSMa10jT2UCfk4eG5bnau29rwNqJwOx9GpyUYPRSwgbkU7uUvoe77WICajWo
WZZ0dwcpPOxRATlxUYMs+3YYaJ6ZFYYe5D3KelOqAhHALbv+NZ0aNWv1WwCd
Auk6z8tq8ZNPkvhAUtQ4uYP4iKNA0eJSqU1u6vdHNTrev/HHbezvL0+W2Waw
y7g3Rnd//FTDca0837KoGqSi4sobFbERDd7GKEdNfgJ0zA5RunRbkRhm6Ci7
iJI59lBMgP+F+BfM3ssJx3ydrPXmuzjdETTwcfmHvd8GusQ544Cef37lfogy
nNH6Kzyv02sbvFb4cf9TDpS4Hi7NTl3w8sZeJiRcBprCyNc03CTaD/60BIA4
fQtxHCDJt9LvLr/KT5noLZ3rHsTz46PAbnQqHiylCzskygkFLVOCl6VBwOCI
RaNFzX+3ZDtNN5+NqGMWbxIJYtOylxBRNZ698J0mgWmxKeL/GIOgZtbkBMBV
q07/CP9Q26iw9OTMYDPD0kVQoSaWJ8A4l42niAEL/UxYevu+OaOPq+B4ei4l
W1PJqFDMB6hLSlW4KB+iBbqVsYX23HLFDzEu5Lbloh5MszhP4Ig3ZnRXDuOK
LbLBwdF7Iq98hoiARnp4EM7Qv74L4pZBjm5L+Juj78O32rrr/8QC+2dH56pZ
5KJ226s/PMAxDs5KspTc9/D9TsJB0PGK83U2pp8eIwKu5jpD6DM+Sv6/fe+6
zF33tYO/FKwMK55fGr6UVSm94r/zARudFaEt3OwwCBoFZ4rrNNExIAfbk1X5
nbyD8IEU6kKNKfdtW5SC4IOQKCI5NCQdmGwnJ8A5Y7UXmpWWH8n7ZrnmXAa5
lHBegOZfy2Yye/lrbwkRZtiBoO6yovUDpFeweRLW7J1+utiv+JMWzDOcAeTu
6U1oyNLzpRCBa1R4AJ5Ezo+/bHD11t7iVB6V4uHHddLeGNY4t9gFl+Dshqhz
QUHynTFP7cEASTyrJX7eoKsftoTYONCyPjEe36vrHvpXmx2xDhf84QXbdvD/
Umt4k0ZsQzR15RRzRigo3NfJu9UjPz2tn2OQx0qsEhohQODqcIFPWvgDIhmK
aThlpHIl5+XP/X2Q733XqJTejv9gRhtPbx9jvCyHUx5+5pHFUCXapL2YoCVL
mjqxoJwal3ICv6OLPNLcwxC0DIKoCuFTmOItiGJCDD0A+UvWZer/bHka4+AZ
JUksxyA5aproRAuH2iPDKKtJuttrQZUyl4iN0T0YPUJxYKfs0hHxGZmzAoTQ
FHnQlRjAl32iAabR8GY3P9CzFb+hia7343JDXZCsjdk65c51lSlipjSAT8hQ
5yFsGsiVPKYC8ZS0yOIASAydEUmeGrFgwp6LsfjdHIglY5dWL1fiQhTU+Pie
9d1dMk1yhgehlXqXNvQitzXNQ6todO2aGjd+1SwoQxr4oBdakcirItfkSg6b
Z50b8Qu7cHa+v5wnEE6rHeahZXoJ7WUIeEH0UIJHB7xlNbwbYNU869gpuhfF
hCmgDQKgVQbjBLsangdik4RZD5KYKcDUED8NCA5OLrqswWwXhZNpaY/hAT3I
L56wcQhCklu0hYvlW6tdp3z6qazlmX6Rz66NIZSTHMQDrjNGjklYEv/1qeEg
+2nKKXCP4G7WrbHmLvuYRWa+iZvqKCIZ6R+er35mQtKobKB0fNW4HEgcHsSc
lZ+5CW87l/FzPhAv4vjCdJnRo8QwVHDRBOaH9fEuQ5NTjMmOpT5H7DxuqT1u
6MflcQR5HxekIM89PFzvZJflXRUOwbmYGtGfgRKH3EASf/RdBnfIoUiatekm
Evfjl20k/06A7CbGrWfCyJRaDf8ip3+OcgZd+PQV/Ws3vRD38GJstRNOdXx9
wZu4kr/4lRKxvgNTbrgkK2C+fvjCe/ie4Fb+dsyH01ZkU7+ALmfb/PEItYaG
xJnDnda2ZDWpEKX5XLF6V7IRGNGKd0CvXC0UpidWRToCt5H1oFau5ZfJZpZF
l1Y5KQwnJiKX0YTwd15fSlUREqMlBS7PgzN/enqTpqVG3Tuc4WosNrx7GgTu
2AV4KhglKgmiakXCzF+/aEEkD//EF8XmHwiz4rGOW+9Pe9lOIXZJLCxrytyO
o030nWBOPkRiKZAV8Prf8OudEkU2MCTq+f68USuS2y26S4+OA/6QIgDvFeNp
kkgziI+kHAR2CwilOGUoXraqyZWbtEY8/sepKbsISP1glCE8qn/QSwjCQTO1
EoFIXkF7Cz4k7CIb+uRdMyKz0+6EjpsP5DxzywfKPLd2+gWENoYemeraFTq8
/KS8sEpNpN9/6Amp3rmagCIEr8kVPmwyLWcwnoFGlMLWG+U2mzcqZt+cQdtf
dDv2Ea4DWUrLCGEtQVtZt7bkpQ9iW/Qg3QlCTsErhchZJZaSkHyW5Iq+uS44
nLGuyhMPZADvhpdO0JMqr1NLdxLU/1NSXx+3rMSyNYruColyUJbV3saEGKdj
3gVA+nvG7gu4Ozn9UBLULk5yHG0gSerloPOk4eni3UmOvna+NVFAe0aHOEux
kTetwawSNX4chw/ReuezM5XBcgfm72kJ+uvGh5Hxd8MfzqsWkubFkfDezDey
H84R5KEr9AWYAVVKytozcR+gm3F2Pm6D+dD+K2nZlh/jt16ZfmZwSHioNGPZ
2epbbjbPMRNmF8a4r6EKX/nOTi5VLFMjIXDKeLukQ4aCFAlFfsEhKb7OuiHf
JPpRGvGRmSnLLbTBPXdEAzvf+oL7Gx6JSbVTwkOhslTdm6oPNwb0lon9iajH
K4LzYnDXQUGfI24pgt2/4Q1P7C/xFP36PFE1NB607+y9PET9S41+2KBNoCmO
pe4y9wqw1ae0T7trwUDKLC1Na16VVG7N1opbnYFsFR35LeBE2MAWIvXdejBn
CZVPz38BQxOAJ9+0FHt3saeXgox7OU/QAdSUVMhqjqQK0EJzKhdYXaKuRNd1
lzTiFWyvQr94c2CTleJ9wnPvchf1RRSITIZo084BUfeaKs6rV87UP2OPavyJ
qjlbub8V1endMJsLtWX9XRoHgrBfGWnwD+dlqPGswXTwbP3JpqaHDwndc2R6
cTN/YtjEtKlCEhZ2/RDFKJZQPqfSsYkp+zIpkUD9h7P2JQhcw3HZ18ykxxMW
vR8c4ecooVC05Q11/AIZ4TWOkEO+OOii9epyLwsa5HjgcBEIEptMbqNBlrNI
kB8ywVv2iS/lJnAAj8t6eqxjOpxm/sT9fsC7JPJgF3Vex81AQvFeBeiPYEVw
YkcundyW55X5GbH+6UPhLrwOFCNcOdNTCQmpYOW+sdAok+wptZTfmzRnEHBx
JVkfQPbBlHdMiBxXBAjFSmbXQgnjEy85ckes70+oAbdb3tVuoXL6Yw/66EZt
xNgpXYXFcc/vIPU+5V1HlZgllSeFbuH6DjsPzSzIZb6JxEpg1MYw5UMtz8u5
sbsF3FZJszfTosJ1Qx2WR/JcuC4MLr6Rjtjq4fzinNedOnsnBui1cMnpJ5/L
TCsPMywxo5/ayy3q5l490dLy6SX2HwH7g4RcEccsWBrms2cTP3CwTJrUtTC8
rCynFn4C2pUgG3VEfjf0CZb4WvmjnwQjqrFrhsPETOE5lQ7oJbTNBoePyDsK
vvPXuwJMgXlvQ/Xo/pe+dSQ56f7VlxN7Xu6dmbYHcL0UAc7r/UGMLAqvmRIY
UwqEH6fBiDcJb6zU0MG4Nt2HpjqA7xQdiKUSVaOItBk+A3sbzA6lC93yCIgl
u50/muStzbSQNE3sMGh4d233MJ84p4+Pi/nUmmZIgBPEeg1Ts7o7IydoIHur
jd5t6KhvLxpcCZAze3/MvCZrV2xcCKkjoyyEHqDdTvw981iYQk/NeHU6j0ME
Dr/litS9fimFjJa342ecD68rQPloOjokcCMOlWYKPWDaNW2jA+NXuTvVtyP0
tpjG1Dqd8s5YahPVglTWqfacV3ZAyFEfC9D8DSiHywXn1IIHeLn4rYyxcuAQ
NqQom0ZdfbRYKHFxeO8+ME0vB4BwNqdjbyK0opJhNDKmPkGoYH2UL9+/lcg8
UyD02TqSoLrys1LZ0iOyXF5XfYdfhM1RAX5BGi52MqtUzp7itUfAN6PlbxzR
J+T7AUMuJBfJXhJEQeUTJ5U7CdnFhRi1bsh4NyfZMKJJzMe+5OQRldLWll8f
Xdf7h7lLKL7LEnia27359XHIBhja09tT7YZqN4O0gx9pK5S/8Peo+OOJM478
rwvHTYqre4/OP2lcsTrs2avZ9PwCkpTFxEWHBqLIEakaDIwTARJjByzwjU7q
aNUbUai+Nj+t3qwSpCXmqnhmH2niNY1CM8h34TlE44lpEShSd7FAlEgRcoHK
Hlq6u+ulF+kHPgIoaf/mU+iXyy/ReKyP7UtaeTa1uNAnd3FDkrnDZ6b2Y9wz
EVaiGw2ZDEZDHoqPXj0Ohm/aIrbRuPYZFTK7238+wq435boYEsRrSHNzzVtr
maGoH6ctwvEyvbAy/hygpcDPK3Y7/jRi8EExegcRTIe+Brdpt6njMPF2AXBZ
IWRhzd5LJcQPsY8sIqrYHPNx4xT5KKJOWI8FjWkv5Xv0SI0KQ2mR+VxqkwiO
dcQToghxiuI1oZ23XYYTGXwQYHWaxi6xBc860nrYrC+6DF9ubHbNuBQEfRHX
Md/HDzXvGIjvSaIqUwD8o8gmFJzWcbh/OObxrfcse+LZmFd1tid6UBXYIN/l
YPHPOJQ8rGRjl9zkM+skK9nKcLJemZBVbYxbyATbvI/3WbQMAsy9RWtPuxjV
7MrDBsIyjlmPoq5Zb3+i61E47UgTCn45TwcbK7BMrkNhdWCC0rjOUaAjbrwO
XwxM8qtgV2vTmz2z1KAARPr6vJ6kw6q3OlY4FZIw2BBNL15wEguD3I4tAPRc
6Yrk0HbIaT01RBzxPZRY4wk0ERw4em4tFu+wY94+GGDSCBACsnyMLsUG0K+R
kSv/yXiaS7zwlSlWq0LOAh+IQbrPVOz5oJo0173CqEgsR5tbenTMAGb6eXVu
LuGRRujUWB1lXjzyomScI0AOX6qUvPfGFAk9sEiEsG0WIi1qY5XOIXQ1FplC
NXWG7IJQBkOmInsR/5XCqHnI91AHXmbkJEAyGEBLIC0e1C+jOUaQoyCFm3U9
Hs7Ll3SWy/mJ9Myuogdr88v6bDki9X1TPQz5v/sgZeY+Yfrsqk2eg3rmXeG4
Yt1cg4VxTKM7Oi3QNyRY0JYt95rsMNQmlRCXvsI7RXyrCssW2VJuvTpNYyZO
otljm42PPJEKXn6674uR5ptWOkrWPeu1E37JZkgwUdeBvu/a6EMQsDHDq4tO
gGc/iWV9sOcgINapf7m3eRkBBhnwgS0h591xS4mceSgplmL2/bv+onBUVbqs
rBqdb7xwSlSElJ7bVS4XgTl5kDiB7hWL/IxFg1NVTpY81qV+WjdiYGQU21da
35QEMn7Dfws4uVkytV6sVc6fChAREsUVtcS0FC8ITV7f/8LaCjhlQWHROu6l
cv5rxeVduJUGfntJsir+F4ppG0bdt1GajmfRklQKVdkOucF4sT1HApZuoWv3
2JQSNyN3JGyKthoUKCVrDMibnzvCBk1EiXdwNW3D2VeKYT/U8A7ZRhqs+HOf
l1dDtAxZ7zwTnXwWIJsuJU+s4vhpY/E6MGGTbcLvdyyh3Ktcq5cIlzv1xTR5
6V7ZPWsL31ei7+iaqtDOKUkTfeW+7645FmR9GPzRyBF95UwvykxUcQyKozGu
uJgK93w7icaKQB5brqSfo7fM+sYn/D+skxxEZ2sAJC+Rw8TVMzrhHg3YHW0W
xt184cx/q3j8lBXBfW3xrprLaf8HqbXKcd0OM9adIreXdiVwAKIbynNpQN5O
pbBaPKt0EhvyIuTmDPBnlF1oUzMcs9yj5orehcMQuS81gnCeE7Ag+EPfS+IH
Yq9RwxWK8ov81snp5htJk1YV1d0497vqAHa4NB16vP/54TdMzKB375Xmb+sZ
QqtfzwN4oIryRrRz/uhSe/pPofDSPsLMmihngo5o02AWxBdiidDCzcj59nv1
0rHfBk9ZanhdAYz/JHvakecH4QloUlwJOtyVYw8QeZtNJvlRA9WxWbPwVqH9
a1bFQJ1OMtHbafZj90uO5f976psohQTCXfcu0Qv59QnnEuRPjvbVlZXiaSgf
m0uq7ZovmOPcB2o7IQzpjNyUIHj+YVKj+UGcRaJbE10ptbTNwr/U31jj7kDm
uQENVn5nysr15Xf74kdDlBDu295P2CWxiGUpwFnNLx+MeIXMTr6pfD8mjl5n
qjslYf0FVnxEZCW2Ip+UEMz70vZTni2QW7Kq4rQpGjsfSjoeMYc7rSSyjx3w
JmrT/ZTV3iNYM1W8kGXitBHFLbgZec9BCC2FuiTtXZsZiDVnFlvDiShfqQ20
/ObrqqIaUXnngnP31Cs/+pyR+RpWrDLBj+yNlS82ITTR+lBFpnU90fge0pgM
+cnZk0hsgEVHA4/Za9KMO8ViF2h6+6kanIyPaoYBxCmlpNqzkG7QwmchDrF1
ddO2aycDJNDwJg4E+0faHvRpR7eGUwGM8M0HXL8u+5ESGPhm6IUHtitFgC1K
aP5AyBDOL++9Iy2+JCEsKN0PHqcUodYu+R2FB6o/tljcXpofVmeq/QAeXJIi
JWWl80y8CGH4FQpPyAQJBV9o4vTUEVE4ew0bwiwALOj5wWY+WFxfnXZ7Zo+a
P0HNmbmTRb1v0iD7ao+/WRQu9GeMbBYm03ia7EPHcTwhZ6q7Wt5s1aInHlHR
9DF/sltDltJk2qwsmnEkhNaW34r44Yi3ToEt0e2PlW1ASdmTHKo0K3fHro4g
Au4U/0JttwNHK3nZTN28hIpIbY6U690ZHpHp2IFwAzzPC6XObufvLRa/WwFA
xpHYND0qYItNBVbx/Xd21uVPX9771TqcErm+1nkrLfgj8FsRAdXzKgnliOVM
3DhsxgySqtij3O5seZ0XWSGmty0UBqIK7mc9Y1wA3XNYVH5BeSuBSowz+LjA
fFpNol/B71QwvA1/gu4te+dv+ltlGUarmx/IHzwu1i29WgknX7qW+XlUt/wB
iYMgs1yRCADKu188G8WFg9zCK8ZS8VpzHhvWBtZDTcLOySaWZI/yCnLXNvbT
uFQ3g8jKmreNh3fhMN7RA67GO8khDZQwjp3JLm1vMtlNFeCReBb8lSIf/fK+
/5+a+DkFT/LmDRT5xKV+fB3UwQByfIO06B+oP5IpuxOfxpJv8cbnjvhPFZdL
Y/sHCU6Qh7tGs2GA8MnFB4opP28DRsUoFBrLDznMcOWEu6FudruW+an56mQP
p9KGX/Ul0mtGMNCVTesl7AdI+v2K8MKal3ccc5V/pSaoGB3uffPO+P1YnnJV
il/rR4BUeK7u5g1VtExvVILuUrpdU0FoD92yLvHrbFQVaWozkXz6yaKjuxFF
UmwhEaF8tezqaQBz97/GEWOsQdjMHnJhbl22/z2hcerON5V25I7Yy8MVELfk
VJhgsFeKUDd+M/1M0+/t6uGs1o2QhZL02VpZy5w5M097P/CovDdYmv2y7+kf
A2dc4GVAFP7v4t0nB8MSStrR3ocrc7jMYvObIFfyWhZ4L6rY5f0BUyW5w6oV
9RpPeo7Kgh5j2roAF7lxQqvspYe0GmmhzIMHBXFOg7yd2tBhsHjD/K2XImM5
ilnGun4MRDUarh2EDY7fMt3wlk/R8QEtaL0dPyRRMh7+wh8sbcoAqYt8XYr7
XIXQi3U8lW5JVoXJWR7W7jSBIoTvS1s5HX4XOAtUOJaYuhzVlvwrOw5b30yg
cSmyJzBayXhof7l64gBR1HtX44vkHgL2mFeFOdyrLz94Zjfhbym0uIDsz8tk
GAl03khtrskRm8GfhjxSdZuswTE0r26rS5bMeCVczRfNNOcgoiFlENzAOhiQ
nq+Im0VP+jwA9E7WZSfGHMZDaC3F0iYcMEkvPQo9fbvno+Wzjz08KL/Cu9WV
jUeXHGhGyt4gCjhLqNaRSTBoct5IF3R/ZCJWLiE/8v60AKrdQzrlveh/ix2u
xeWoPujj6BB1gDXMPfhj3Q9ELOyVfoA1uXhhz0jnDEFUOnjb7KbV7odywW5/
s/D3iU0Y2p974+K7tVP68DXtCfTTKbqORLbvq9nSILQ19XigaJAaiQuNfPyw
J4hE/gyQmPz/fsPxBSX8E1tU49Kqp/G1kAW8ycI9m7zpv8Phl9zlJxVhexe1
7tnvjzokmggZLLt/M4sTGnP6qtgoOO2av3DgG9dtDi9OD1PBQYiktTQt5mMy
QuM0UxligUjIdwa6zdzsyVUaNjpQSpw4cPGdPNjJb58wqMgnFY4CxNPnvluL
kA0ONgXn/Rp2uqqYU4l801cxkAM3vwk1lW2DXKrkBpApGydV1rylTRuAgZkA
ML+nFhCUsoXHcFriNlY3N5MPNtzXlx/GSQ74KwO78OY9YQkk8MPaUDxTM/V3
fSFdgHPswTWOE9gxd8H12fzqnACFlM2qvTUqSQTUkrjCmgpm94OnWVwvC6gR
BexxNyCMAfmKa0cLvFQpjFfQ9S93fCbPp/zCm8oDdjQM+Zu3c8jClADquotH
e78XnHHY6h8UbjFrCWGENdG3HnP0VdKS44zhG6ZFICDRg02zSZsw5bbdvWsR
T/ILFCn5KeGHooSIUibF2ETu8NkintL18S2xgbdfQ1X8IbYK4IHJghg6sbb0
wNOLmK1XD5fr1cd4QkBuVUtnLSNZF5IJ7uYGhHZ0fg90vrhXrDA78F2barUP
jL6nkB679rowU3/Xtfcw+d+uO50Sy6pGayNYcqJeofMk+AQtqxvP10AgQ7ON
0YyA6rKWiJJ0L3tRt38VQaGySqSPnozxd5snf+0ibI013DaSTpMTl4RdRocg
qlbrR0zJFxTCtWnrW7Ev8fhpi5ugZwPkSwG/TRq1sxtCY6kq1aYLXaA4XXpM
ksDy6JIZNsxQo9UGZfmRJ/4kTwEDwQX8Jh9udA/eDKgJxmxybRfewVsuNMXD
Y3hzWShQgwdoTl4O81E0RB2jGmsFOIBZlIiocsnSxAYcnXse3LAI/1GFCMat
VUmRGVfiZRukcZgeW/z4JmZS6EQp41TeBCKSrH/4UPA910f9tNIkh5USGfCZ
Wol7O/xDfxzlAF7BWVk0KIxGXkEcceaKUxYsmdQ5l6wUhX32Rr6jmLo4caQ7
ImgX1EfK3PiZ+Y3pLhYihQihDqjIFVLSuPLcKDJwH+2cJspfx8HWHPLVsnop
l6LOtaIGkT1FVEGo6BVItuFD7BKoKypeuEf03abSrBFt0V4rZRMZg0mnzn0f
7QnUnpoOpFM5n1iRSCV8H8TP5exfGB1ZlrjRNLVeAqWSJJCNsRRXNN276Xbg
9PgpQ2ku3QrOoj3tBIgz3ioU1e3+WwPgNvmrGo0dZaYC6aUgO7tXz/D1EFA2
XhzwOD3S5OIEDn4p3yHqNzdJELOxl/ZcwNY511GAwTZZSzzbC1gznUcEqnW7
ny5AyRiytu2/F3BCjkBEiYKEAhD9nA0jgKtC1VajyKMd6OyLmX+yNCqBNQdu
xRzIjn5BqCdnXMnWahMO3v9DfHKHY610rXAS2X7XPHrZA29JhW2D6V3toP9i
BCar2UiVlHz7KZMsl6qlyZYAKXU+aGjwGnd2s8FBYQ4pJZvgr5rHolaxN3gq
6FrBLvcBbmK1d1tlWLHklpaBzd6vLOrXzBltxfn8w/2+9De4meGFyM+EbebW
tuOD9m1Xh0et7g5l52tPsqJe4hF24tfPK9cezvi/sAK/wDXzeMUGQhsVDISV
zBvEKeljsJQ367kG1mC0HV8XJi/nP1fJxEL+5zbdSGI7vuAQKpB63HSQhDJl
oIJtaetjAlo2c/DHLTfvE1tcBAIiluhUeY9syhM8UXg0VbmY8OLDZcbSGh1/
tUYQDs9g22EQvwXoRg+ptVoP9JTUCRPFim6GiFuK+L50Q3gQeZChU0oiiC+Y
0m9g3oJOxwug1PmHimTiLvYDi0ASDfDWcAhrItz4oqYx87VqrR8F/qbpXxXy
uAiaQPxWZ7L/YMQxPvVp2M4O72hE7mhLdaEWPVipoZw2RI9Zle4PCgW4Ms3P
hua4uyO0dN83yoQB0UvtH5es6FAEKR+MVkNfGnnZjxXMRPmMKki+dEH1JSsy
P4JUjnHBWxpdUhx9oTiFNT0Ttme/70wDEoMl4MZsv4hdaKK5u1f4An5gwfFH
MjYpa+LQ4NKjV7zHkYKilvClkkuzobCfBZAUAGGazk/Gh1+1iE88xUaBdg78
3wskVJa2iDTg4yULHwiyv3leFY/X67pn7frbI3jaEED8OqqmBHPBdfMumzm1
1DdvP6WONwhOqUuYxRRtlcCssBWAk2j1Rc/9q9R4dIxZ9NIsTRiPr8vjfzhi
iLj0xwK0gMJMSVm112EeTRo3Dqf5GOY3B7lDC6MzHhsJpUeNGNGhwycT5WYk
Fsyj//tqTz4hDMWgvmkL/GKh5juygx6vWDAkwP5VEsGGm/U8qqwk/F6kaH6J
Nuksrr7FSNjdDDzp2WMljcDjJEzoMkzod11mYdEbDtUCxV3zAv6++J9+HPhN
NILMCSHYhzOLoZ9FN7VYEma9Yx3FvjErSI2nyYIJVoEhCMwfu/iC7C6E+hcr
Mz6XfLcjGcxBp4B8bUaRqZcnphgjDtwsDzC1B+b87ePEUpxtbh+JDoZShUdY
Z9q5+CcrSRWOLczwKHidmjHwdSARS9OwEYmYm2wRLSfXBoMJwR6inXv4TS0r
Xyzb6csbtmtAKy/ew744zxPjj2oB/RcEdb/i3wCfv76Top2lpe6d+T4GVbLw
iq1YmDESRqg79/DtBzcLCvOvZufB3MkKIHoLCkP6xYf6jMVmpVw3kLCNihld
8W78BaZWttAhonBWZPTxnuyC0Xd6+vzbA1/IPKqwxOyQ2YGuygT/kgdNWWKR
lZQ151ADPHRJ60WW/AI2cD/cCC7dSR65T/RsSSUquajUX75PfFNwhK25zsuP
uc8HCz2ENIGxuTCDiRKoAwUpT5cRF5k18PB4XfR8cWS5E3oXtknicMUAk+4m
/H++XYiiyDDbwQn5Dt4chXjG3OXwSAsFuLZjFXTIzWgxTrUH1dvqOke/Z6HF
+62xkR1gP6Su31XgoW07dfSJpZUPu9kxQe0qntJ7pmj0p/PELOQiD77HHPjQ
fOBSeBNtrttqtDdRMNV0eVShJ/OYk324EwvTjtoajn5k/dDF1oVYhA/OaRt4
LHF2lcnOhvtES3Jus9haAGh1mdagPTNdi3OFgQrOz9sm3gg0agOu4Bs3Cxf4
hN1oNtdzcjbZdB3dSAlHHbYudTL4CJHgghAz3C1rzurlqSegBHN1kgK5zc2W
bG+u/LuR0C18Gesx0TFleojMGxl+Uwz34UJCRA5qJgLk3QOlOfXleHd37ZSI
56M6E4dTw8QIWzFh8FZdcQwe6He4ej7ossGPLxRrXJTDo/HTq4fm35dN/E/f
4nKrpxHKSKcZzvIaa13SyM3x6UF0KU6JyHOsm4GaGCIj7Emm2RTp+uqQsnAQ
dSnaGU9FiXaX49c6PG+pZncLYC+sLys4siP6aKxV3kFPVli2pVWpABzCPbz3
AL76Tq3tLsuObGqjU3l1nvagm6REqf8uXiKaySDmybyCWD2Mv9uSrjx/TkH0
fhNiu1lqkWVgT+5waKHDuq3eaSyhzBkCeouA9Kul0xO0JEsMg+MA26lh2YyD
2LjvtDq3YVNazkhB4Ep/ArmG04isU9v6GmyH+XO/VXgYgbn1EdAJcloRLmx4
/ECaDHhtjgdS2lPgqyO+8/PfKVIyU1FYK9NHm1HgDqM8CeUdkyqWYQ9+4Z98
e5paQzvmGwGlY27SUB2OVeZe0zFvXp2EC6J5A98nclKu7NaRo6k3u3dmWoKU
Kbgm6fXLQAPnYBcHepDm023hZp7TUyp8V6m7EqlGAZgyzP0v5ls+lCW9o2rN
15J02Jf+qhzowgX5zLAOCB4FWaLUxVficoIcOpAvQx+1Z4R09q0ZDTdwe4Bc
VQmg7o+9+tpbguD0iisC9jeCEQP3MqlYB7k5dw6ygcBz+qPpDB/RDQCA9Tl/
Kh9zw5V//rTFny1lHLM2khII4SgLzuE8eEFYg8qlE8ZstZ4KNWrDrWWJXbEW
Oai0sJiWJflTHBxQVhKEr2W1sGYHoqJRQlCT/Vv3IyOQcAa1IN6kV5WuBnUM
zTpqcCKn/xd5uRxdWaH5kBO4za0owNjyu9dWvoMN6IjQCHXQOTy7874V63lh
bXq+U8PBNmcaoLZOtKvJj/7hVuc3uyJMth8Vgz1B04+f7/7Lmptzj2LbugDP
zgrfMxQENH0/L6Xk13mAzpsw92S8Zc5EunU2gMugxxW489rhzHs7dU912bMK
6tVuXDwxr8wkp2stAvBEETsJojpaKgeOVs03hIp9TAUKHEvEnGVksqcwYm0D
ItGybc2HQPe2iudxVaS4DykgtvSUvZDEAdUGBLi1hd7CgILZz14Fkop9faBM
hNpEwARuVAa6gGLjV8SdK3PD8+VpW7xEzZ05nNV4CXNqeM7BAlu/YJrSM3Ja
RIvcqHvCCkxx7Y1rdcdDAUXpk119myWL0BZts8MqvY4+W4dIALQRyA6EPfJG
qshveBe7Xghqsm0WjJ4M6HBLkG4Ll4qxOtlAwiu1dXl+wQFODcAfuVeFsRfi
dr2MMiyYJwYb3SX2AfnMDsuhHRNLXbrE+RwcC2sdrVYPhCtcUBOec6WxDAll
OzPd6k+Xye8taqk3vJTlfPDnVf7s6iXY7i4Qn6T9BZ0XN5d6rOFmw3T0oxiv
qDLIN6hMmJjwc6SPlBw42HVdHTlFn1gl+uzPuZ3nG0SjkxeOYrcZoOB+QUxB
nGqj2vMCwTsTYp3ZgsinOtBQOzXbmvH6iVrhNWZKDh6zrQ3P3g3Zt3hy+quB
MJguFUALxneP44RsDpHRT8Sj6U4qA5BM0gRhMDXHoRg+BPUIoVFJTxwXTqFa
7FgEL2K4k7FtdR9uLdUSxBwhjqPRgkFEMv58vodLnTSyB69UFJzwdU2GASkx
wbyuGictDekpETNIsysTevZ9mm8tFiN8q2oNRvamjqsY31fsmPMIlLvadQM0
wrauRP7yhWQGwUFGj1RmnyyUP7AH+63tWYfBuW0nzlIFGI6W1Zj9vzyABmii
5t4hs4Khz+ZLPo/KLmi0vVyRKVgvKeVZ0rbdoFa/Oi8AtiGWD/oysPA630w5
AyarT/LeTdoMdQCYG4htVPtiEAPfksiz6bohF9TKks630Yx/chV7Le0dycfR
AYfJNPcW2Ca41/3iJXS/htEXEwqw0KFh6EmDS6Nr3z5p8pw/TUH0h82YRpMo
tDDHNL5ODcENppNzDGm1rjGDY+dbizuwqxrWqf01E16ME1ZcJfqOMIH8Xeny
iUN+mJR5MB+iBwpoDng4yMP5VTgMl3V7CwSVRa4e4Y+Alfy9kQQYRT7GgmZR
+0miS/Kboijenu76ITM/OfIXtklA+EsCLNiz0GsoLiGGrv5tgmM76Jp44ZMY
upk9z7LJJqVX3egkk6dsCX82E0p+Oy+KoxhK3iMGvYRZZxbhzRSRbpaeRit/
HxWKbU3sxAz+AwUms2rRW0hsvznYJ99IbsNrejXgASHXA1wVjfUvbLgfYnGl
hmDbqg+z5+iHyXqV8E45rNk9UjG/3xmLor7gF9aeMTHldTEYwOdM4/Fs+ZD9
peMTEiBbLUx8kUOnxZBLobJKCL1Q51Ga/MlxsTKQRQQKOkbCKgBI1VupHyI7
iPNhZl2dCbYxxXim/EPNpciRnl3XUN1jXAOYBz7ZkBm7vdYxbmziQVgMC2ab
GQBNu7mM9w65ihc6Amz5fgNU95Hy+tjfN7gTxXRFbhUCS22jRshRNJrTH+Jm
f2CExdbhGrH01wb6syaA1bsY77hNlsIJpmj2VQGBWZodMQEVH0M+VSar409J
Ws83CfrbaYmia1D8ddXSf7l33+OAuNP8Ql16igPXggGm126CeZvhORf+eBmr
qKHaqAXqv32319JolFlLt/w+4eIUdaJNJKShZ2amSwcX8Vg6WocrA2xb5e0p
KWiU9iq3wV/Y/E6AL3iSRT5ji1sTJ4QlwJojy+FPZKI3RFqLhjnv2Wwjvszw
7s/Nfm2BS4bX9s63wn07+uzKElWOxj+9Je711Tf64+WcmxZ/odHPo33ZQQci
bICSP2OCajnbp+u0pIvPCz3u9l8DiTqVq7yKgJEp2V/vHKveu0LBsInOfl1Z
NZWUuiy8zF4/qDpCjIWk68nfarNa4/IqM+4Y/RUSRb4c1fgZXvK5uE6N3qB8
NShlh4cx0/3cg3b1WVeJuTQ0oVHdhI6ZlNR1saXrJoJ3vuXQgY3uxmhhv6Cq
JrOhrArn5JgY3c+JKmsu6WtnbfuIyGZfopuanzY0IW36lUehlG/H4LGIcKii
k5GiW2POml8pJHSBHz7L6kJmXmHPHST9Hk5eq7KJeb54Js65P080nJvsE65m
iJo0Fwmg1QoGC4bkHRCkk0gkY6d8zXJGMUuUGwSbCSNQq+JFLQKS9nCuLNHB
nObpRdWc1rAbVBAU+n3ys/EPd1APm0qRD/4os/7Ysn/mb0v+8DA8cdnOjgYt
XvsTgtmEZpLK+vtRjdUi1Ab2JcAqvg7wOzQkfkLmA5uP4NJkGbsvi1V1teJw
5W/TCwACvM8ckUfGek0ES10Ct+kXW/1B4pH06xiFxDX6avXRkf0ynXJbavo/
mA/xGGabS08/IumZSpUrg8IC0D2Y3ilp+yRq9tKqB/fa9h2OhUmQAuLcrqUN
dGaktuC5OW8p50GgcrO52RzdHUZv0v4lU/mlhqMCbYH1N2wS7Z1XcdJNPu64
Jq9hQaeWze0fxeTMeORm2RkT3EZ1JBgRKrWPEPGzHf4LnMgBFxKjz41HN/sS
JL2D9kKgoMeZHfVgshR15f2brUKjr1/rCkYnfWUNalfwZ0bm6/YFZf7J7WNZ
4kYVWEGyHEO1I1NWBNNnsBmV0Zjt4tgP4r/LvUkavVJcbkHeJyZwXWmbylMI
kG9VqsGmQBFSSV0v2ZTtfxZGSfw2DHFQudJoO2VZuHZOv7/LpwObfu0nkBJc
/B27C5S2nvfIVBIp3oCTgQX0W3sxotPXbSBPMAGornEo4kRgz1VhTh5W4dNi
UYCfss5o4pUcZFsvWAiP47cP79dabdLasaBNOioJcW46PAOPip6V1M4UKl+c
hnohjNXR0XSl6m/rnlEaHuxkJshjz2a3oIetCnzzLLSqSh/ZMhFwJ2BPNnX7
eu3yg1WCULsoE/eH0aM8ebmG7VGe65aZNijFEL+Qf6EHMbxrlJlPjIyZ54V2
d6oA66uXDQ72QC+CxFig3ja4XkCVKrCEr4lzMeqThwM/BTVuhdN+QYoCg8Xm
WIXne9eUHV6GF2sPfG0sNSE23cbHQaEpNkqylSM9Q45XpmY4KxIVqu3mMln6
OQMTCe2h0eu2oYNkT0QAGQsIaeDbe6WO7vdjBRtxxQBMFPqAtPrrlOsFLrQy
zQeBYYW1cgVemAlC0Kd4mVpigA7R+yVfgESEOc+XcbzNCke1VjNAPa2OzRB/
FwZVrHuhMpo4boWujhHqMpzlxJuAIr3qozyyv9iP/MDyB01GVd6vAegw/8oO
D8ltbR722oymz7xZSjh2LOYlRx05ARNwEsuZizmPDImWStChb6gtvgiuSau2
crtR/Mj9I1Ob1qLci+z0rH5VPsR11EKenSoyfWxOM83wQIsEdj7e02rJyOfF
IAns5/bG1bIGgV7P/7k0n1ZoZpp/mhk/ccHjhvJXhh2RMOfLhalHmo8zVnSo
hvcVDLKzcDvi36mbWhmQO+7COHDqQcY9SIloCtVydAL3vKeNkQ+FYIDzqjTN
hKjg00EIyHAoFNlWn2ed5j/+RlWY7pOKeGrmSoP9IjsuGID562Ul8uONTSgn
gsWzZVKZuEj38UruPigHz8RoSvgRicTcWH62zDpcJ7Ryfqc2niRE+A9tXmuw
mRbD56Xvr5WOBk6oglvYVayDN9NliHAQIHNKwXwa1004dY9f74VWKQbsI27Q
OkX5ieIIUpD9B05YnhxBImiNIEaUVLSwFL5ddOcHTLs5EWroelx1JQ8UDb2E
5SpY6nEetfLbHqeRQGw0HTRhH6io4uN2Y1BKBOSgYkk3druZblKeFlXZq74T
ilQcoo28Lnh5HB0PMFRX5RlX0txB0SgobWhj6ugfeH6Y8b6bWLRz2q238EQ4
IPnLrziRPoSbA6KPkdox08t9h4VQ7FKy3dNWPBFq7eEN6DlnARKUY48MzzgG
UC6lEgNO6CIupsh9qpC8Gw1VJB5gKkS7XcqqmykY0+/hGKsTsVLfw/qxNAWt
kHoGuOV4x0suoG2cPdJYUWTTzKefVFzFqXXF2X8QIJZiXknxiBjTVYxlZAx/
Bark4wEKB7etkrkQnWwP5FF7AoXeAXH4km+YQcBJ2CIe/eEACq8DUOO26fEC
wyVFQdhwClXtDFH3XEahpsXpr7/fWJZpL4MYTEFfCGbrSJ11tnOvk5pIPdPo
RfFdUGOWZZUOIM+3vbH8Izk9DT87pqaX3VlPHehyGe6sgJQA+61mHJLy3yND
LvdxYd4nUfXz6bmALuuZYJd2HGUEcc8JeTCiOeD5uQTcWmaoF+YxvnQTCDGO
3s6/h+27kCnabJnESgOqlZEjTdyeSfnD05sWlTep3X2zeZUd3vMUvy+VwstV
QlkkyPUyxnAjPWZQUdE9/RvD1Mfa++eSDgJ4HqABB1dlJ1YWKB7K012BCKQp
asMR6pWzCkaNow3tXVmWUVfRfRTTxxLUh7ssXRaWO5/DCY8T2Jph05L9y8qa
j/wc7Wv8y/gtoSDBlpXaZw2T0FvfYmhobwdqAg1YSWRvdCO/9GSMpoK82Z66
ksngQDuDyU1cHLc5+UP38t5MBeaXyhnPCnUXQlxJIh2/6Apb2LGYB+Q0H1L/
T+43CEF7P7tuqg+/FZ8QxPVkmOy2dcJy41w6o6D15RvB2Sm9TDTlS9cXgAMt
0c6awuPUb5LsZQc881rztXTEQs+r66s//jXSw6cPJSwHAQ0/p/0e/96hfrth
iZrtojULJph+O+6fs7rj3j9+ed4R7d41B2Ksh39KExH6MP4EgVGHAqClGB/W
1/h4iCimuOWci3HDg1uVMs27M04Hlctw1DDDlMK+h7f/N7cA8aMnZhpXGXRk
kT3NPAgqUhUF378yYqHIfl4E0e9C30gF1Zz1IGSpwkoCwuIGhhAtAn6SGsAG
OYkQ739ib4liniAT/k9Y+yX5beHZqIMvVV+RVpmI5eaXbQ0MAEDbdg3M8ksn
8/N+MmT5+yyWDIMq7AI/qm/uSttaPPebbNYqXfMeRR9jNRlKjC/CsVy6q3ia
kr4/FqQORk89JTRzj13MB5uLva7E2gFNh8LanjplVEXo8AHgMJ2fYeCxN3ok
/7kMvUjihe2YmZ6aMHH2beVXZRTLBXoRxzQbsxxyZbbR2cH+W8zUQD9jEN5p
R6j/R3I0WJ94VdkWjsEhyvD0HZ597fAfy+maNiN9t7ZAs4szqrw8+V5xUzM3
KFv0pexx3miBNIOsLcmdTxktRUFJzAp+VoVSZMDiKm3JvO9dT4oXx9UDwDWN
XMLEV0qzv6zM2bP0WDhM1wHZ9RhJj4+FCSxzYkvB7o/UsGut3afhBLHKHN6B
AF+ehywbgdi3fVjKQNqeNYvlE5TzAajVA94x6dZyuCsVmxDchhulDDSGeeK5
39yMVqpsAN7Th1taAaY6WFS8WzTXLoMji+VsHw55AoB//kXcjajldHQmmQ2y
urfnUEO97uOsIMnsRR79R/8FNrJofjnkNwI2ZqBNrApBeKY1GT93H7M0DmA/
PfgYNq8RxF+0ySBmLc9xbS53Ab239h4UCTTGxFt966Zen+m3fitbNSoxx79T
O51ZNogX8S7hTEeprpDTtLipL9wQDuEA60B5Zg11px4fEeKMPgz82VizuMtK
0xUnZOpkRjnoxeOKAj5ACDqEfCbKh1GZwvGCYajDFMknXPGJjK1/EAMJTZlg
CF11PsL9emL7hWr0VuD1Wm0kTYLc2HW3sGMJeDY1mzqnGsPEXU40VIOWz6Vz
YoapIAJnSo+3vGhmp12m72mB8HxXVHB0nLCqXs0n7LkHie+sXEXC2RD0Bzxf
jUvKwgnTMlEDX/CUseut6rCf0mkDVXzGV5ehFRmZ4RblD1YlbaXXRtWLE0Yq
Td+0nFw3eCsmCsDRHu5fwatbCSwuNXMqly4PPHWEKbQcdUg7JY5gp3xuy93b
87qwB0E49r6HYjLv3YCZ4nLinuZF5e3fGn7VNV1hW7gWx+ABCEpzhCBCqBjW
v/tGvu6ucMehwKhQTXqYHqO5T3AFjkMvmrkLa1b/Izc8TKw8GwmCj4keezft
Ome3Oygo9iylY90Ks54vVyNTaRw5tMExqrJDzO0z0RpGGqnAMafLc4Wx8+5F
A4jXhfS/zXwzZuH9A4lsGB1sULsSWSDUJi0ng7uG1brQzbnK/lLVn75pq8rE
8vb2oM5rbJqCvRNb+YJzUXNbhWzspBKpCULCL6T24vwc2RoSqFqT/6PsS58R
QXBw0XPkW+XNHkrC9rvLFWR5nYYlQKwVi1K1KmJ+pFD2gGABa5XKxw1mAlSH
mI1UD1NekDdAqIl9tEClZPwZ2zpmHvDUQcN07Z8PTRbh5wXhgjjZUZc4JySI
NJkkpCTcb/B9tZiEfjdt+H3JgmNC9JvZ21HC5giAoNb4aRzbC9LiGgZUVCtn
4xK30wE8b8S13id522YpdjUzcb8QGppJdApozj1OAC2VDoIhjCQeNji3IcES
gc5LqSWdq5RP7mt8HCfP4jgyrpZbVV42d9QMLjnsf0ReqWh0iGa/L1qI0yLR
UzaiD511FEpdoft2JOp9bY0dPvIAd/MpREQ8GPGneByMxNypdNg11/Fua3Ry
+Jo6TegGewCEe4i63Afwo8/SvCnR6jKQklI8W5ZqC/ERur/XLHGGoNtQ8Tag
YkjrWbY8U+mfSn89gEDUKst6dbbOYt9XnNbdnTf8aydAXqQChF5Xi8jYi1Dg
o94tRF7RNpAM+2/CdPAJ4UkRD6Ke0oaXLmBtjbLGay/X3+6V5t8JKRpV/C0J
uSswNVbZJSfqRVB9qtksvyJDXuA95SMRxIq03eugPY7t/osIL17Z4WezgxjR
7IIxamwa3Cs3wclz3nOH2DA3aqo+PVMbmXrHPb4ans52kFApUUG/rM3TyGKq
cX+u/KO0hsn/93POU5EVXJfSqBaYh+H3X7bC7YxVd43gnwTwauCnJbH2JCyz
y36v3he4cStWn3+Zd+oxXmzd2UAGiNtrjVM3yejXThqr9XYP/H4iTWxMs6Fm
Th4rf7T0hOsP70q8B5ZqANIhJc4FI2if2nUIyt8DjhEAMY5Jf16R9GLYyqrl
55jf3fKpsILKKsTrdi9trQDoB6X2TT9tu1a8YwLaTrnBWBKpQdJEyKbcOQRN
seojI5vp/ae5C6x4eMuQQ5BkuMXexM3arzhtfgcWqsiEM4Uld0AWkXn3+O7H
I/ymkpO3jTpCzY8b6ZAPaInLpZHzmRqUZ3J/tAZUB6wDAVVi6/kSX3cAh74c
Z4ISiyOUsA8ie75XUYrpNVg3U7t6/s1z1lWqUPdvULEWWh4/ioDaTp6W/zO/
OQ5t1slkApKav516OwpN7LFPqrMzVlj1Jo1fBDLwbLkfHS3DYREOL/ENq9Jw
biDONAijaXXCCsB7owaCa4Lo09wj2IHP/Bb0k3r+B4FidQgY56yrQsTtd9tp
gfCcJ+KI3PH+CSkWH5kQmSiZwt+YO2tYicPqMWLQbHueNIIOyLlrVuFSUhWZ
AsqxKC6P7HIqGaeiglPb83CAzECXQMOcFrbFqEN8NqKh+FDbco2Bl0aOW3Nv
oTIjtz5Lrie6AbkV8CyUTUv1DnE+kMlaFfXUulCssu51/Jug9TEDlw36EW3R
X/jbKTOdKZNwpgRQZie4H3QJKg0VkWX3B/xLL30PYkPFzojpdxIjdAXCnplE
wtrskq9fDo/TQprzc6j1mJaF6+WuJaOfBaQP8XM2BWP9cc9X/Yyuk2svpI9F
Hd5vLsB+feGapC5Y5j7vJNYZS4f67dSN7MP4VXMrG13PTut6snr3Mecvvcwl
vsQvDbjuuBPQV5tWmmNiavPKpHExTgGFtbVDZyvcBAwkkuiD5eBve/mA48Pf
kwJ4sw1Q+7QlwKQoPwEggCvIlLfa1OT5rZ93vpKqUVqSmrQoXdoS7RBhWtTR
+J0ToCKSZq6cmMBpZ4GIElQpg/A/nO6iZSNnWRghu0gOEIoOJv12BMlaYlTC
M0jmYoLjgNVb16sYpncZAqg5MooAMopEl3RRJdn9hxN0T2F4ZmeHRYfDzq+g
/TNbMFJFujiD+3C22dBQlxRotT/Gh1bI0vqdqFa7oxKrzzz+4TykRedGMzcV
2Mh2Q9k3YT9PgkNqyUq7BJsC5UkqUuH+1YqCJq7sqSXZsUdmGKSklt/u3k/G
Zq3yJ0dEANKTUcZIVbggQA6e/vmOgFR4iHVkwlxvf2/njhD4oCC8crRpXDqJ
826wL2psO/tijnvZB43wnIwyM9hQYoC7MAyKZwuELvrRI4S9CCZq5qsymUQj
+mxUKwVM0vYPgE0O4JhDCyF6Ln7tg78SA4wpIBlNabEhyTxLN0v4+vO9aN0k
8rP2wUBrDNFFL1UZ3U2r5fjLrfR5wrzS4s5VCDWwuRqxfxQwQxlFXXgJhwde
Z6yUC6ObMQUvAw0O8iC9ubefq61Ucyw1372tjsqrlmB55k/HQz6rJW4Y9/to
yZhu5iy9RJAmz0F9HoDNlYBm+mJuHgxutYg9ONajBI4ZEapd4fOVDWfE3BlY
Dw32OP8sdoNcBaEGZwddbC8K/x3/qAL9Evbg6EPxQjZ7trSeILfzocWrv/Kx
JJ+3BxW0GQXpQA0+XGUuxrLHErlfdwLVhowNLjA4oEXJVSjaohemBJKlZ1u/
mPS8ohXFAv2WDynLHUsQuHjnRvrP9AuF+pYZ9QJk+FS294vI8iNiPaTz0U+h
zHJGr5JFFmhuE1No5R+MJ8xzlV4zTIPK0NewLoIeUlJ9MA/jLWFuwwe8KHW9
fqbgUfdeDWrMKbjeAD2RF9U/iO5urm0aEDFpfjJHYXpJSFuLuFsM0L6SBK7h
3So6lrPQ5PQA9RmlxgrkWH6mgF+WKQ9HBMyXyiz8PIPvFP+UxXAbekyFo85V
Z+kgFh9d1WA7fUclnBfaRzm/6yKSEYERIG1EIQhZmglICODcUFOucLULsI9C
Cifv9Ok4lF/fCeFeDBs8dT0JxmJr1CEJFyIZuO0qIVel3KfQ1gJgREzGj9Rs
YkAi9icV/lYCpc7iADlMjM9wBYFYxvMrhoclnWeF3qvOb40EstEDmrfRvoG9
45dLHXSTr/ut5cisfNsxgd07EykgIKOcgTCQam2dHb+2OEPTxpAR/N3QCh1H
87i5iTgfmGVcE6Q+s+BT5tf1PuwBDZYlLdLeTDx7d+1ZGyjfivuLR1Dwm+jA
eC3ZrRlnjoOhwQaqgQ2B/3royhQiedCkAF4EP9JHiq5JMolVZGYzc4tOvYqN
QPPNli+66af8hhhWZL5w7cLpgUz2ROzNaNnCKg3D0aAJ7k/dZDTzffB1jqnf
gxA3rWLRrYqT/WPPhlSz8k/wOtK/QEz1mxvNbEIkUClcUWOMXJ0cn3O1+GXK
5Lkb7T++9RjqK63p6zhIInlPbnlCHlNXkwk736CGta52PDc3UVvYtNRqySB1
8Q4rUlW/+rmNcb7XRjVpRdUdd5IdKFhrC8lssZcPpiWwtMDuJhEFGwAd9c7C
L+L/MVW4MMkZnuXfCqqhgS0ldGoHxCuSKL5spFOdOzGYRnAFOLYq2NOUMKA/
tc4RCoaGAfGBYXXBLMOk+tYuj2I7dpwYwBEByfDNE4xu82sCJZ931Axiv4Qb
mhnP6r++stAshikKqQrUjenyAWs2P9mmBGYupIYB3jHZoP9XG7Q88SQZxPw1
Hfm0k1e5QRExGdRjaZBC9YMYH8+QU7M9kmFt0natiYPiVb06BO72apUU+/5S
F24KZQWWnIyYmWkiW+4fTDDZipil5z5DuBg+wmT3fmAZrCGoJpvrM990+UJn
d8ph8hcqgQz8GP6MoPD8ZFIiYTnthIo8usEu+w8Pft/BgBgH8o5hnqBY+CIt
Kl9TMWZ3bwwxAz26G9tx1NarkMtFSNIkRvCGzbFnWK4+Zv8fdRseTxd3Kh2U
RRRjp5MskMID9bf9ZaapshR5SIKVmwaQT+UY6IZxU6jJytrkZSeCFp7K1SYF
ljo9cVBCZCI0k6FG1V5+LFYOUXkH+Mzpk8yP/aLqrKRIRS4wb0Jk/Fz6B1h7
Jrcvy0yuVwS/7x+A8Ed2kgDegJeyFxBLVv0OLPae/ru6MskbRsMdPysC93aL
NM/imb3ViaOdKWPTzPrqE44BpfAutjr2mE4OCKYqNa7VSGDk2wVNs/hesuep
InnDPLjJ8w54nkGyr/slO5ZwIr+LGcH2QVhhRiv+rsCRipmnKvTl8b8MAPoV
uhki8FpI2lXVy/Pn4e06OUgOeohfeLkTtv1uZQDa3lGhZ/uhVYzB5JrfTAqL
OV5YBAt69aBoA6ZTSW7N77A42z9fJPegljmfa4EKS9yZAtoTNmwEEaa3OpDV
t4BW77zqJ5FuwSDEyXTfYyq+hgZ9KqwDaEv+j8XnX5KL6X32x9njz5wsTJ+u
5OQUBanmeunD9puRRGEII9hGeFgjzyzTd633dSN5BQ5wpt9acCxJYMuJv2OA
gX9hOVh0wPcSAZQ1QruPp+GXWDNNQncpl4k54jhOd5RzxpmvOMEgdxNGd8+f
ks2Tk+7HTRf8JllvrbCZEsno45LMIO2DJQ2E+UpLG0UZo5Hl2sDY7vMxXsvH
bg4JglTsg0sxvwfMoJVNo/mWzKKEqebFHgo3aXu3M/OD3BIcV2U7EZQSarMD
4VCbSutS3ukXDQH5+DNDHX5Yjx33SY+X2P0gyIU1Ge0kr7P1usxpv1pBIiF8
GHSQKyiT5gcJZsr6HUaYhG9HBFxccaFyniyKSD/QrZIxYwptF6KpsmD11hlg
hBt+S7YEVVeTBDlgPollPbM/AM+fxWpq910HJ4baY8R2t70doq6iu6TDzYSU
Ptxm2qbzh5SnEyZrIAc9g19eWLLFMn9gH2pt+p/MK37lYxMGGzVszCQYWhb7
e/8LO/RDDK9scph7kpZ+coB6O3MaSJ89/1YTjRuF0i6pTvchXJdCwSscsM3V
bTNePMyJaP2kvEQFm4pzF59nqvPTrV9bfQTLjgg7jiWPLdSl6Mhf+jHF2Y3Q
XFqWYeMoI5oNVpNQHUJa7IHQxZfI653dH/FE1/xgCe12WNvBl3cGVKlGn1eQ
385LvPb0mlg6LphlzMb+SA975BKLiEx2Xtjzag5/Mp62/H9Z7MFwXZvCJK8m
oFuegvQnhqBXCFAKbPGpwpWcxILNcF5e+1wtJOj2YMbu+3OpQKQnBMdnaxE9
OD7063RmfhWo1ct56/WxCWLnLDDnWvKXv3rEF8ynMOOtImBxfgsBOB7fmL9d
2jcJ9cg906d39yGEL8d7KmQt1LcgFstGpWglmFv04zcbAClx0797SSUsjSoZ
8haAjhZpDRWRryJ6ZzjiQD3ejoYKh8kjTN9PVG8Pb6Buq6q5qH9z3JdGH5XM
5yr3/5KBh959MjRpHaKikl6K6yCyvdH3Rk1fC9CzKIH/0CFTkVRHAo1m6Kxi
I6eAtAZ/eVVMsrtzhxtQNZKBIHBo+KcwLnhe173lsTeaAf6wttsTZADwhjLh
Ch0hEGSRpfSHLafFxM0YLoyF4Aq/qXi5rjW98LVjWLTgk0Osz3pp3ZsvcVRA
2LFftbYtxLDBXIMTlvDOWFHb4OPoAD/d+2xpxtU5u+gN3ITM+xZegk1zvEv6
4BNO9qfgNLaM9BCG1iC1GNMhbaw2vZcNkLM7Qnr1VdgsaCmzZknb4V92l3ba
8wDkbxLhu4tZKJYvFOFxvnpYyjQ5+ukF7HYPs8KEDyQDw9NHVCjmSPYtpRIo
XJ/eIQICXtxRyXSwxVfeHKIiMO1uh/7DOq0EZTuolYQtDOtcB+iiwzMN6qpJ
3rzPWwM9n6MbigkxnW9m0ArI4uzHdsgfbcQHWOIzWn94UNy40htWhxhb/cQ1
5+hMqxgcrXYME17F2pdxB0CIDZGzTKKt3Jy4eFsv38E4Nb5XCH384AT8Kens
d6V4SyjjxFCwg0rhHQKWElal3mhlh0y2JBNpM+74qX1Dc6z2jxqWkV6F1MgA
n7vU5NYoF5vvu8R8FuPAloeVqOxHoDag2xmKnYKvhA6zIusffDoppnxJcqgN
Zv6du923pBDsVSTLhjD3mLrvMSrQZknNDAqGwDAGaeSWAWDy8qMdhx1iFqHW
j5BMHzyNeOBjtKjadAeirrBbrIZi6Xzw2bpfgyvXWaFCdPqWwi7KmFkGF6m4
ezOeB9vuWI0jt5wZ01HZjZbTYzCBsG2vf6SixAki6nNmJCDOVigzUv0Yq0A/
P9rYRa81RWkj8LMxMHXH2gLFQT5FXrN82h3KiUuBzKwT5ttvO9c8mLPqGwit
klLFnmNdvggGz0IiT0f52NCQejVAKK2SbPEwIXFnuM0w4ZEOQh4Nnu30FzBs
ZCqx296uxkv4Ut3/2a0NozR7YrsGWO1vtqqeKn7NU1JorGUlHWqqWRxdWSuE
7ZC1G9Ba1kXOYOP8eYNibLxby3leuEwzXlTK0CW8rsZYGWx22aksgBhlnJmG
7Nr4yRKuJnjRyq97QkTUrTvNuVtYkMv1vvUP8JTfQCt8PZRRW2vMaULAOtHA
634cpYYBSUfsBFuFZPV4IykTbqnHyBM33phoaQkMLJiY1qzPn5voGOFCxgtK
HPYikATfDn8bugCH7mhV7Q0OzsLPuuCWv5jwoYw4ycsQki2aGqwru8cciCJE
uEdE135N912hGSO9dn/O4amhD4kFLNsVaVBwPfFHRRLnJquOexG6+UBJO9ZG
bq9jNVp/pdGhpg62GjfBNPJXOXsW+L1XHzM/RXYd1JqbzY326vK062Kj6toJ
OXwdNWIzyMUlijq0++Wt+8VG/etiFPDhXh6OscGyFTADWDBsT7k4L5hKDCAl
zGFYVBSUsTDpT9v7ai+5FJpp/Xf7gC+Ka8CSocWH8fhR9TKYhaAYNofS0g54
kjMIua9SeSaHLVzQeRUqIaF+17LUXdI03IAMoNjkn7p4C6Kn5HSVovql4n+y
LlFFg/WAYIgMkD3cI4rml2aWACZX4MJItKbgXdPytqzYxOzv9P++OCOWVNty
EvC7qZ5m5gEp5sycngp1Qq7P2h2xqnlTxbpNmEPoNGAZuxe/DkmBlHVW+xZY
0/XLdsGeiqQSfpl1oW5IhwyNINBIcUWopZsTIdn4DceSIKPIoWpgSlZ8X+0D
IYCBweCee7//A5aP790P8y/fMRHmWQcld4XTLgSadVQD31mvaMEYzNs9/Cxk
jgRQbxF1PqOOCJXmlm/14haeNE9lyJleL2CImDacH7pW9nzfFNyesqs9N/Ig
AuAXAHLqmRqFN20kg1rAg8MWSyRPzHej8dzTI37WkdWBVAnnk/Ln6/vOpb+2
VdNPoC1B24g6ndwkr7FKFVwA1nfReuz1SVrM9VByjaYbq78EUCHRwpxW1WId
lGt/FXw5m0GXMALbNZZ8EOWjLWRZXaA4JZ2d+ThVQMnEzqkPkMr7NvIWbNkA
fE8qtMqoQ+gVlWvJRFpi0Zf8O+GkVeeHEgI22FKBcuTQZre/ndGNdxW/uTP5
z/yMusfDlbxUwwQbfERhtSOQAkPYproekXuBbaAZzZWW8ljkqu6dPizJ3P1S
ux06JgjHtbhx5j0nqR4Gv+IjLD70k6+X73gRxUxulBDJf33xpd84yyjGgAiV
ar6yoNNx15GYiSpBWWNLBg6GUGIjcOwkbEqv9sjAzQNiOBb4QYt/jiUqEfGm
Km1yMZ2ZzDnnmiayME3NeiWiTxjXrhlkniOC/fUHQgAQpIgaHGz/4b/RVvBK
2DwnrfUD8Puh3pT3g4NXP6xP1KTynbDMnZVweZUL/6bO6F3tj/AqvH0U0g5K
SwWvxaBYBBPXHX8Wh7cG1Cljb4wX/jLDth6FFHOLLPwlYOClmApedPuKjpEv
PbOYEpnlNBpivIC4W692Ak2Nt7suetCVBURyAlMSY7BIxS7hTWqrp1akd4za
3/hAGmhuHBmVZTPbMoTG8tIqgRv2ew0g4k0mz0zmbB9iCp1Bmx9mZu+5dGVE
rj5PlI2qz3JTqIsAG/El+y9rHHgJzn/nIDP1ARG+jTIWSVzGXsb4ulhKndNX
7pU4GWEffCwT6iwoODQT67v2ivtQaXIJWiubx7pW7AQYNSvFaaKMIhRqREKT
oaxgZyRHVxvYX7o42IkISTN6E1qxXh1hF+8aJpUzA4dnR2UUOxC1hV8LJ/r3
CSRImVZCPqaKQ0dk02YuRYs+MFH5eQkowWJcA+2YdqlE6vzPkNIRjOUV3zzx
1QhtgJehBLbKLH3f3MdAk3QBr7Qi1ya4Zhcsry/hL0QVVtmSSZreGOy4svcq
5gf2h7laAgJQiw6fLMVsT6xvqzo7nAQgsUvdT9wbZe6KmJQfC28ZBt0ziRHB
aXhDjYDVKQCPG5kXsNKb/pTcHXwtFmQm62YKfNorPi8wRSdyng0ubfwcAiyO
YBiVeR4IO9iyyXmrmNN/3/6eIq9NudXkQyC5QYzjsst2AIbBK0Z6I+IVVbfq
1aPiKGAD/LiLwixOIIl2FKrnY+JBpbKd1UiXajlaO0JvbGFAYMOACs5jqnTk
AmbyWe7gDTptEpOQfwkUR42CnDBOAs+lfryJA95wEh3IFZBxBiaaU+RkdEsa
+fmnSwJBfhBKO0JU60b8PDGqrMHBw+H4sPbOl7Rrdeg6wA/X7if2C49Cnouu
1BuuSCmSxaxbd7PDY6CbtIXSCvgMe12ImoTwovn0m2Bcl4bPjtErIZsYpKFH
QwhUYeXzoV7tH7XIucEtXMpYMOEvVXa/P6zCua9Jq7B74u4ksVgU87zXzszh
bGu9lT+Q3Eecu35Kd6mxiok6x9YVNm8L2smKUumXrFar0jZ6czOUQXY4TpwU
v/dGYDRvubGYy9SaM06HS325P+tyFi8OaR9904ET4YzgLQbiaJEPIAYlYBUA
Bgq+MBQyNCGhw8XtDenj2yt8ZePtiQ6tt57U199vhvvjL/vj+K7Y8i1gcDX0
C6F8QqfxCN+m08gvfPDHAIr5Sikq3RgaLHYwdPQ8fjwhM5m1s1iQ5kQZZ4jU
NMGg51gTQXjuwm4K0OxPjMRv90PycRQBxCGDWXu32rxi+ZDvjK/NqMDEY19K
rRqOSrOQlktrqWcqk5ZKAelO1NCi9+JPfdcBkqLyNITrbW8T187rp4u/eeuQ
cExX0ybIeaIyeBu5n4y04BaKa/F/Ejvp/PoOwQ+Wc/Mxvnd5eKGNRtjBynrp
bPHS/Ti7TGsTKE5YuSvBeLTdpXmvxdY7PycN7A5+3GZ+H5pR9e7B6A0JhoIX
hHEaaY6nqQE2OuEupksTpR14afJjiWLXpZFtF6sLuDbwEPcg1Z136aA0dKav
pXmCrScvS3nc92aN0nPpiaGavQn59ORULZslSglqdYUwyZchEcoxMLAQuy/Z
oUzeN03ovIO230ZG0ca42qiRNHDq05Xcgp82TLrnX86ysXFB8yu9a474dv+h
3iQmY51Ny/m6H+yLORwCFcTabgX2dlLaPhydr2yZDpGXNrV3tdEyeN0LZdPs
fNqQ62oimjaMQnBijRfadPCdyJcTCyAabmdcDNjnMG5afppj1VCAWhsQGZiD
uiNvux+VZfl1LDyKhWHY5HGfIGpxdrtboprGzdaYIYdASsut7qTOGejEUoCA
aBuoNBsJye0zk8GJV8kJHqg3v9889JmxRZNLgT6N2b8W1Y17weDxIOs4c0bE
p9kSP0rHHK9e/Pwu1/xTqXtaXebMgJCFPw8C7TztM7qSXSb1jb1fcj8VMhln
bnLkthfGAWgYEwA6LTOu/oHfcpN/CnBV3vdRivn2hxapvsah2aab1M9QfpUT
ksiAZ+sT9RM+j5FssNUdJJd8AY7Tnjb7VqBr82j8h2+cNQqTzI+E75y2nZGm
bRecRVEGAzeGRlMYdjfXA+JQEYp+bsN6YCbaNqneOdBEKkMWYVJVuOonxvQR
PJkc9qGJiK2lcY9InqnUGVEMsRbu8hTpqFGRcf8xACm7Rjmgazpcf6MOApHO
wd/ASfTRD8Vhi855rZq9Vbgtuwi4/KN1HW4KkUwCk00GXc+baXstHc8B3M9V
VNl7xYBcgQUH2LOLEDtwFwAhIwe1xwLq+D5hzgjzVsRZ2QF3nOXoZ8gY7m1N
7p38kugTlP1PdleXjGTuAc+AUEq1i31eEBepBc5+60nwi8iIP7hZ2F5hPwQ0
0FO1M5POFcJJe/oLL3V5mitZdUdGLyP7OCBRv3Wj0qd2nZ2yPRou6oVweBFU
+B8/rth2FOXTA3/+oc/LBAVfHBBcwnWcylaGjwGpTtQyJgKL/XdX7DE+2BSW
+Zx9B7/ZySZXyejHs5xTi12Xb+eMCIlIxpDPCZG5OgfMO0Ces7tFloUMz6e/
aFTK1KvJiKo9I2SYJPEQDtwRYAtyL6alUG3L6I61hYQMXfM5Qb4GVJMxha6o
bQn10+3ydbk7kglRS9kxOCp/+CDwD2LsX8CAQnQFOwbfVa0s95EF//xEUEFs
vrosQIH5A/AUMnThAyJC0Uff+HxedjjnF1UzCyvoYpVXm5MIh1IfwsXaGugr
rFZCAer72adiq5m2rZ+lWW84Z/1RSWRlNeNfdJa+vNkYg+qsnjPP8nWRPr31
fAtLd3fGn5fT+VWOfX7VaHbfDmmRkKyrAt/K4ZlOE13JcHMWM+2U/UCu+GYF
Sohev6/4TErf0TUT6VLBt6KsTqo0WKFROtJopeZDlgj+PotkjgQ2oExfSbFG
Wn+zqP04uK8nH7Nw6ZCYRlWSbM7FIQyt3Q9desDOxPlzfslcZ2OBWqch/jCP
vkCKr42jJzFr/w8JfXEilofVPeBiNKzoHoJ/laXidnl9DyJtzdUlHbob/fWx
Tjj4k/0zqaF6gdwxrjLtfPB3Wb0Agq64+IahAsITnL/Iq9oby3pPOOZNV98E
U8ZFosEaP2S+UVpklLovc+9gp03WDmL3L4oO+UxJOR9BIffUN5Oxcera1v4z
eQx2TtutJcUgmNK0i5EUoUeUqjJ6KDb16ybLqpZEhFDeGq2xor6ur0lD7HHw
clCcJK7eiH7LUmjemezWMv9yM5dUhn4fyTf/FxQqObIrQ5KpLSuGHt56WXGR
9Shq4x4Xq0ea3SFkegoii/BuCejKVGSj2IJHvi6Ye+gJIL0d7h3CWwR8aCMd
ae/IrfRv8HJ3NFbkdqotgKQR22F6+OXKG5FI2TG6Gg7Mc11zoWRZ/cGl/PEN
+T8nR8kad9KStF0095m19XCoGO6u20CH9om4FGVGVKo0qYwnSM/Ku4tk8+YX
c1fgRLmj2MRylTmglvwgeqlVMwT6vJp3phjDfxQxWtlV6qBSTJOCxLjFEF5A
gD9UU1Pwfq+obJ9rW6TiJ5ylMMW66f4CLM+HmRN0E5eWYKWNO9CZlGFpep59
/7nA4SaPFMLxtfwL34cfbY9Zv6q/cFR942+ArQi9/jT6ArJDBaOu4czyjK4H
fRLQq/YdoYu1UDdz+yIe4d50QYrtpTKWIaompd/vUris2h7gImyVZzNUL+T1
75s0j3Txk6/CbsPPzzY0TjR6hg0ZAwy7EyS4wzLZbGnJFN4TZFdeq4IJwRjl
30clpuMyTi6GrCQSxmjb5uyfPn2KuJhyKBadcsWn6iRiL1+9z9pFSABsl68V
f282LalgdpNtN/kbEup6H7kfMAU0mAhugbAQ2cat+GT/2NqFje7Ov+mJBf1u
buC/eml9x7rchj3ah5h9Mq/QFBpbke0VW58o9lZPUF/RN7lOXrzAxxTZtKPb
sJi/UL2KpVzGfcp3+QjPcqCDg4lFO1WUjbaz57cRZrEJHCKNffrog4+5hghI
gIz9gmRp0SZ8YiwvnzkdpJZlp2rju5FSW2lIBfuSOnVyi1CNvN8Lafb3pS2J
673XeL44zrVWYDl6Kl7QkeUnklgTPIj7XRc3lRbqKdOVlaCbYunp4qsD9hdm
Rmq1XN0U1KlQGSNjBTsjlcYU6LRyg7nogFhxccMo6ofRqFLKIsYVbjeDrQ7B
ZGTNbmn3cH/OuthyOFOx/9ssqL/+V1aji63S2HtnLZ/KwFT6krUJv53THdR0
TtPhNWpukRkXfoE5qdnyhIb6NI5Bc1eUT3cA1LmtUQUEZQ2V8LXJssZatxqL
1iclq8p7cK8j884BJnlqImguxGpP8wXbbRiRhjxDfFaxBh6Zks5PtwYVSjIJ
PMERtZFvl6pW1m4cwdTKWvMV8ChccCLKRILyvMlXes7/gkpif8ALtsqECDcF
28WkLSf+ix0lW48AWgHNab1xZhqnLghVqn7IAkFWYNTqykGtKzSPbJ8pF6Zr
sPPiZQFTEdv7fkBTI5CJwtMB1FssYi1RuPnqjfF/KnKrmKYnN9i1ITXHBWzu
RCYsb2hb5hiykLbU6VwDkR0rDR7xhy6zf1dqdNidCa5PCa1IJix0qnf2yKJF
EGhN1lFlWNx5RTTSbUry9NFXmC3KbO/CHOohcN5g/f9RdHAoZT90xJb5fIz2
K254TzeYWytifXdSibYtn1b3wbovMZgYDNkoTWw4cWobqQbRUl9RE4qCzBXi
lvwwm48QuGguck0NrbpJWCtPstKQeZE5aCjVgpKc5TLeB+Fy5P8+IzJUtuwS
Ei6lgjAQxLVdo7iZuXER0aVDXmqIsXpYOJHzD5SDoAmOeTVNLy915wsAokOk
VBBuQPmBIHZeoU77+Ev0fPP5lcFxpaiM3uAqPID/dIr7N3Iz5A2+qIf+YvJG
VgUZaHlWZQR0bVlFliSIzDLz5D13ckdZhmijcJB4f84UJG8SZKaAT+0CY4Dg
sNMRKdmIDnVL8YTvF6NPv4ieb3Mf/bf4bLYPQ+m8HziDXyceet74Pb/cwenK
sv26hG+J0veDknn71DI+zyzOghIadpQUaznci0/2VDDxM9V52guXmfjIVBOs
+fGHBKl3/EyTmCyyur0YG2LqJrXuaQYWAntmnszKNVWRRmBxTFI0szMKqYwp
kgnGJJ3WRQIZZiEY2S8rVdhEZOjX/6gA0bhs2RIjvGOqZa7KLMJciV8kQDlB
mwjCgDJKBwKon47FPevfY0hinjvtXZOqi7sIWxl7H1wyyWzjE7lVnmvkM16n
Hq8gkINv1KHJzVZiUup8JtVlQWv89QWYxVQwjNLua7WzzoARPyudjZsTRdmO
7OUUbNK9uhEAQifHMPsmTPvQ/hgZFtnN3Itlt0JEm05h5anI/UliUyyHtiJW
OXAf4P360dyFrjbvK/9H9y2nXr3fMIqKXTP7xOxgiNV6tXrUo2E8htV3UV1V
fxfGnjdNqTDOjhG0MuRmQHauXeqW8iklArFNvy8kH1axZEaBV/gRRT/cYH1R
uHg4aglizdHiJQCOUduFjPXD89gVwYgp/Kxn9nn+kPBsELrcm+OTMQPV4d+G
b9cQZnFwAsgt1r+uVbJTkUOqFENaBzeAVyqJcMeJXzhtLfDGbycsH8f9fJ2R
BUj7OP1e/o0qn1NywSvAzQfdnGED9iGpOD1SA1budTJPWSdXGn1KU0QeFqJf
x0EjBecF+M82fRdfVYDq9U9Yjs0qX41CrSj4kXMZryOubp8Abm7hjJwsIhPt
oEMJSCLOgUtKwMpbVHl151dzd2CDRd/TQ7+VhFf5lDtBkF6PMuWtHiPlyW+y
yJ+vXtie8vVkA2+7XXVy3WbrLWC7vH4Tuo0lQ9FBrIT9zW49NUgLUVP8640C
1zUsA5JuNLN/8uVxKH3yeqxjaDIIIZiG6R7Rz09/cAjBiub7FpOl6a3KwT+1
6z3dSESOgSDxBhAvSJLAWQTTShqkTX+D3Cl/Uwab2Va5xwvxLs4A1f4hcrDY
4PfqehZ7ylIoMOUbIoezSp3N0UnvqEMt2D0No7f3ZbFtOt4JJ7zOwwKzz2h1
vDhRnWualKspYlr04s8qSgr7F5NhfCnRzz1995LWeA5zHUnNC9RsW18S/iqJ
C/hALE87Pizo06VesF4lyrEszh/pht2tRA1L7/kzHxB7MMj2WThVFHRM+Ry+
nW33D7NORS0nvstrotvYO3ZETSZC3x7dqRdyjuAYvN9d9MJo5G1XoJrOXvw7
VbmwrwysCPtK42h8Ltijq5t6BtitbDv90tchFeNWLFn+ZiTFkRyPtG7qao8D
sSZB6VyPm7/RlbneyKNvyzCqg8fWpfsEOCw0BslzU9fa23iXAJcTS8Ju65pq
J3OjwUWV6zicsLtcVj6Gl67HXIeVuZRjirm0a9RgLTvCnD/1svhvOKDBjYKD
0bKDEk/JcuwngO81p2Y5DFy0nO0lv1Tguoyub/ijIV6jOTVlODl2txuLZfP5
xvMJIez8pqAE0pt8Bw2BA8gdRcyljtnFd6am/eeC4xWbMJVi1PIAOv3LyT/x
DQXPA/Es4tFYf/CooeVtbVH66qXJyO5HmdTTJ135wjm41KqpA++48QISar6g
qOidag8FTYr+TshvOZz6zHJ7DThjizZEy7Ydt4bCJrBgKR7HoUmxx1kwPnz6
eVRQay/t8T1tUTM4W46ZhEtHYPtUv7UW4zNliilRhkVR554TdPwYsVeTyijz
wSo92Zh2eZFuETrGz9ETZ1mphObrP0yyetUcfQlXTVjEVkVfkLI22a1wxlRQ
pgpYu+/rwAxAUHtqIVAYB1yHAU2jJbr/GzpgM/S/OaPCJ4hLWnV8OV0QSXg8
L7ymM9TNd4JzlK3KF+PL65Idb9vdMN7MOvnIGThrdlCz26djJvpT9d4mpI5y
khFt1nk9Xzw4oaiuaZ5C2QGrJdXLzRYRkIWYh6bjP43CcE42ieWoMjGsyZB3
qfBzx3FbkWx7GJrvZHG6lfv5pGi7KUfuruijAAuQTXin/3YjrQgSBauBx+jK
Riy2KkOxKI3vyDNm5X6ptlzkxGzMndX1uLO5tDRC+qdCqsVOUQLf2nrVMnz3
PiV5J11CfmY21K8t3p2bUlyydO5/O3BYOqrz/rw4h8QIVUTATHLPbFB+9CgZ
PWibU/2l8uLNSumhqFtTO64oH//UtoNe8jMOgsNAk4KEdJ1VTOUexbq2HtOv
DDXnUqSWNZtu+xebutH7H9KoFeG1DJUAbPX2pmcUsILa/XbWUF3eNDzEigk+
kTSRlg/sHAasAAm4GfdzzSKo3SYTEezYMZbQ29f/lsBqcFC7rwjlz4+4rTH/
cjRdDoY/T6ktqux799UHO5NzPghd77Sk2bnpTikizJmScgdYI3+m9Jt46QEx
CHv8mJToTXXiAiJOISk4J4bdtUbESYRwRavJZZhuPuK2RHG8o25PPvqVi+HE
3neGQVGjOjOIZ7XMwyLGwX5ciyQu18GojhDwwa3XkvKRRP6q8RXoGdLbAP8V
iH+87CDfHZLN/qCu2YjMwvejYSqJ+tpqdycncRrkIKpxKxR0qagqT9GCfWmh
yhx+rXjRV5JmfhPvQAKZxiNBFZSC/o8w3Z/Dgh+i6PpRMaVvmzJ9nsuMqKPx
B11BuYdr2u05zmAGoQ8bevXXGN3VgMhEdBxuBh93LzLyFyprtivd/pnuZV7D
uRsD1VsmHboLMr15cNKY6Gf+J8dt/Dg9icuvbz6DogR/JlndcNgq0IuJ30bz
id4SRLwM6oDpAjcBORPxxIfJB5x+iqJZr50urkXmzvbbsywbFpmqxtStzkhs
IGK2qi5+EzG5jAmunMd0ggAnefYbNcH68icXPe7mXZc6fcdaadtyAynv4pn8
uVL9KOge+1u4RnNkAc7iM5CtWlDz2QpbT/O6lNRBKxbCaBQ+hpCmxuXiYWYF
Rb+TgScwbA04vrvseNp+6wY+vD2g3grjXPqxGT52Xjf+XKiKLP3Bu1ja+rjK
5hlO3st2Q462a7INN7oCjgvqTXFRHRhceb0mWX6zABBIyc3L2haKtkDuECxp
GTdz+cMaw9touAeodYaI/FZv1FMMTdCE/Owq8yzMtHaE1EGkA+ckJWTmDpoI
iPgiK0P7Fyp3KO8FJp0Tk846bocC3rUeQRjOkgXe9fpS+Lmhv5/WcP9D2hCj
Ueh6zlPaZPogHhb4zjmFHWkCMlN7KGnytzqiQ6/k6xjflc5R8biTbQT5o52C
MmtYUGv9FofhDvf3lly+sVqbeY+7Y8F283u1bahRAAJw+2d6BxFaLeY2S2h9
EMxxOu2dqmxCdF+e8afo/4XxhG3H/dLwViD9MVA+1vuPBs3TUvYnv9MKQ+Au
OMzgpBtib5Iui11J0JjD5xrgfBbuB0vHSwnuS5IPjOEMoHLJusRgHrzxzvcp
5DIYmy+oTgLIw559ENHnyUYExLB8uQzT1v/4s71PJG+31djT2ERJTtscnYBL
/5Ip6T2UJAzBpFQr6GTbmgoUZuJKx0qS3rFH/pUzHO3tr6t8yKsvNnfv8BoU
5DXkbX0cvEUVzT0ZuOIebq9vhjfSoYgk5/rz7bhgMSn66knkORsV4EMprWnF
bI7AFnsxRqc5K6+5HqbdJWx5BNAeQOQ7ae2G2sZXYuLNql2/8SKwJ+CP4AvH
ovXEG7qj722EDSjKoUgNf8f+c2pzIrpGaQ685FabH1zefN/FuvugyC2u98Zr
OiRlBXj1KhXooG5f/xj4RoEDaK15SZ5u4kaedEwyW4UT2z0yjmh/yNXgFN6X
Kg8kZYSUDgdBZ3ZOuzoMt1hGFYNS4AGBueNpwwoHHJFuONJTeyFeJDyj9ueY
BoeNX2JEhhGOmoNv4225+Tu7mNo+zumlzu7dWkVgujU10fkwH/6Z0vE5CsBJ
rbtES5aMhQJTHo03tcU2rEQ7trIWJX3pKZewF3/kQ5FKfM+uKBWpYkuhtCfQ
pMXVSV+AFu/PfCmM4WJNTG6Na3nzBxSknld9endEGrL0hcZQjlCxPrA0r3HX
qDl6YBBZSwH/N3Py/0JfpUegJ0OLxh7BjO3+JyDd5rVUZhpKWz6/SiECNHOo
C/8uEJZ6jChMCu7DKPtpf0Fqr+og6SE8gYdZ7S976wJ0Svh4N8y/QZkJ6WzR
esD7Z1al6UxMsp1Agm+Kdf7kvFOOLocXz2sdEtg8BRG0px0Yt8atu/V/fkUt
p9A1JDbwREkrZlhiTKgAXKYyQIQYKjT/0ZF8gV9WNlswQrypgAdm73Qx//b+
GIUT3u06ZEYRnPwVb4eaUq71OpUYPsHvOLJjXDZtd0UXhT/mTJQA6JQ49ZJs
l0jMhV94p2XeL5v5paG6vZUJlSKZlpGjtIYUdDtOOaYhw5knZWDGrQ2sfYVd
PaJtHpJS1hb0PNkbR+zNXMqDHpLmZelTpBW5GARl0YTJSiNjvP9Y5epw7loL
B2ehH28SHd8eo9r0mwuHzotA86n/axdP4qNYlT/+pDcZfF7dmNZCAuH/jvv6
x8aWywAxe9+hl0GbOiU7aB4EUJKO21j5QFaJzwhcm1VhOOGaSGYGtkt8tgo4
W51/6wy3K8qvsD8QuQqhfiOLYL6G10H9QZLmKkEuYzu6Eonp4+ZeTkYVmkBT
EoC+ivYqf69bFNHGdKrQSH44QIp55I65J8nIJ1EyNMYpf3bym3yc/z6ZVHWg
BgWfSHRUnV+6gbQGYJbUR5rsQsB6C6NouFOIv+TxIS29oKEgIDXNaG/B3lpN
ifP4qFQWFBAi000m5RezRuAVkT4YjKC4lldcVbV2Bycy8sMCO3hqnTGHlhKW
zJdONiGFngUdEYF9xkYv/9Gpd4y13GAT2PVYtXdKnp3fun3ZDsG/pGCkXOsD
b2nwmgc7nz2wYfcgD8YV5cC2zCdOIqbyXOrhAmXEP2npCiOvpiuMqdkvIj+J
BdKhIfC7tiMKCeKB/Xb9mltLDmXcBL8OiHgwMZK+D/aCvnwEelERgSFjzXBq
ixWAZiU74i+hnLkg65+XMwLdXzsD9n9uRgXNvi2zU4Hohxlq6ATstJzqFXJ7
aHEplbtByLdQ/CwY1EEmncGBtDuRYLL8IE1E6hIYzCQm5ZG0rJ6OgbZxulZw
rfe22R+wU/mFGgZpCgUG1L5WRKAKTDze7QdSjqqEmoNybJeJ7E7KMWI1EzPY
kkwBavLJNV+/4VNB7iVDbT/wYMUXOOPYKYt5Nxsl39uGlThoT2yvBY5c0m4K
3yLWNYTFZTMsLrRCRrAp3SvtX6JvYgOG3ilYGn9CppgthDy515MAjL+LdXIG
PCfVM3m7WlcUQwSAGe2bRyDu4swDE+zfWsSbHYrYoV0Y1C3U1Ui2cKJH1P3h
UvngKCCqaiVS8MG4SdWz6XEpUwYKmPMVkQFFmHGtduJCghsgHpa02vZT9tXq
7MAGolII15MnGNnhdTgsHmo5PQ+UkG1rSXryfQoe+lt9JvGrH7ytqA7m35yi
+vbZDnxeub30Wh45tyo77zOTF9JenKiqhuxUV0Mdmvep7B41VElLDV69vBhR
IrhMOZc68e+rWTg+3b4FJpyn1nOIh+KHhXfBqsW6qowFd66GdM7Mclv8eNV2
VanzwDsSw9Fbd9wdeINc+3Cq1XW7+hgkEJt0gFsBpy/43gC17wEGEAJfLlu5
VyQ19oJkG9FbZ/0Jb3tZWPwJWY+TAn6KlfnXJpHWENRVteimrxnIhcwydJQp
C+atwEPe5953YC3M5rveqDJil0E35ahH9WaYavZakJaM+ea0QmUDzWRBQ8wC
ouuvmX+NbRC5pI95d7/PXHiJMGn4HxtM1JYJGfSu/j4EI62zn+6pVG8MUAbu
N5RNbMDS2jo0jbkKxSQBF/mEY14dwy96UqITUKeXl7kKvz4McqV+rtwj+Xeb
m2y/TJzrkWF3B7UD+jZcP19lao99CaOBDEBdrCKIdcMgD0ZXb8eSe/86b1eq
TK8JzLBov6kN+Yk384Bf2/Df7qS5gv8E/rw9hmmX/ZbNt4jd69riX7DoBwmq
lkkcgZx+2fkDstusyMCZBQaB9VFBS2Qh9A5CWtFa/jmwpzJzWSC3c8KZYQrr
E1y8PP9+5L/G73hDPZv7jmTb2PCrpOGo8ttzkRbdzEmj9ZlrT9cIlwBQdT8G
3s0SIJJjbSkkSxp10RXoQ1VdAFYoaGsYIplIKXn7rWmJL1CK2z+fRVLbTvvl
lLdX1V4ZzVPNUAYvT+/ziZI1B5gBDVumWWyWIkDlrwLNE/weOlh6JawhL0Tm
MQMgrJgzfMppzWq5ozqQExTr3hMa6/tPHmKrlNmyZ3BwG2BLIQilieeO4v9A
1Mw0ZE9S9ySAdQfH6JmQLjrWvHajW1ty9wOVJdz+wP9tNGNM2AvbBUTIlkh0
QukZc77yXHbLJX8HNKM0aAlVzLznWUo+alcEwOEQ8U5pI+5MEoc1+zB7LrVY
kKA7Xc1bOIYcl/H0DmXITQOXxOL6PURDuvsYs9f1H7d9Wpq0gt5pIJMXF6Rt
+iR3gfpGxDQDDUTNPxsxcYMmDmmCb6L/FYLhy3Cbsdim53I5cpO2OTbCIqh4
oZxVTpirhVOQN00IyFpM+83LoKePb2vyC1mlzCNx4am0QWYH8wzjHrw76tRs
j2XwGWV5ZS9EzjyBxeWVoGkaS7IJF8Ll/4TStRfkonWPLVIhv9SUn8tej4O8
zQTsSBr9UwdBg+sVF60IGyju35kKAe5yVe8o8n8tN7LdI/xsbtxltMUxVoJf
8Ql64Bq7Uv07kXZNYFj8aKriW/Gjcn4e7szMI0VOrjz6uyCWCheDGFHtIQ/P
eg0QA5dQwYWO7uWld02cQCB9s13e4jP93LrrWSkH5AhX5vX4bV9hIe3YFlBy
bhvf545ylNK30WidkGO4b+SKqD5m1/8iiuY5hTav22gBAmRd1eiD5ndt2UL0
drSnaGW6xMC8Wq2PZGOC6HU9aFf8zDsRNpreq1DEQ1aRNGCn+euDiUIrYuqy
rX48PWSh56lJJsj0gUSPI11CgFC0pxI3ZulPB7beylt/LcciDEKtJDSovxWy
jlmAg/p2vZMeaoEdXWlmIM+pM30LSxKwzzaltFxoe7oJND+p+4n/aVgTUJot
Sq65h5XfQVk8UYE72Dg751qyX2uAd+AlCstQmufSmvDjRa9I3LP/iSUtSzaw
UO1RloEKTCHTE9atbfYgpQDKG4QuIXsqNuW+Jga08rVr/jjOF47sTXJdQbls
MNfgphmCnc6gK0xeow8lEQy4WfB8pFP3jFA3jfGmTUvEjSV68ZaYUuQ5vFG+
1Ui/OJSE8ewIufEPJmXm8H3OSqS5y4kUKwHV6JyQd+w3uNv3nLnB6BYhGfGD
N7tYD3Mf4uTlsSpQWSCJ5dktSb9hJbzjIDxhqNsIqgQn2C6PY4ldxG6CGxiO
VyHLkMEFb5NYePvRlUkX2cscD9CjG628Sb9QnrqhurOPZev77QJNT5AJ0tr+
tV7NipK7A3EQrcV/WAvq8Ug8IbV3AW9AQ/MQPwijMe8RAr4w3YvU05YOkl+B
aiQWU7TLvb/0GcnTQcW00Ooz12oFEHWjKzlNmTxWEwE0MKKlKJXNNkQnd2Vm
9fvtJQfX3TAMNj/GRq+/dIgpN1RYTDFQxH3FCvj0/xoovHWj5qroaqD2sVQD
1ZSBtJ4gygeVCrmK5oi2RjPl2O54a1MGfmJDH2As56kgZFFflScBN4JOuDWc
DubseZBMVlpFwOIKank9/kLEhgbzkYapGTltTwY+DnSrif4mIuMPYiMTfxUv
RqVdTQqn0vhcURbD96E58wsEIup61fVTL1nBZm373Qm7gpmqZcWAQC2s+CtG
4v4sfYhQn98CZMauB7NbtKN90/yvtR9NUGU/T7sNkAIhmA0Ht1GqcEE2I8+3
hhrM33pufndKtOiJs8a63uXy2wsQLTnfMH3n8cBgh5rv0EPq8T9Thmbe8WAo
IF+Kyo7owwlkk2gtUHCorv4xWtIQCp0EeHdE/MBtG2eQlaoSYOvqPO/WLYEl
QfGxazawpEi0yKbzloscxjKpmetdJ4OMhkIErkpUtYLABVHhvZ2RRDTPZCBk
j8oj8ptVtQbXQ2vc47O6okfMs2/hRbFj1acjeehfLuryi/I5eFpc1CJ+OC80
KXFWrLwBT/vj5YWIsdm+hLMBfjLs1AvxZLEJoE7kNLIKajGViFlyUY+zH7cL
Q4w4OpL5iwzMYEiUzTtYKsq3BGG+WDrQT9qckGH7I2NmStX/IurIIwndkySv
CJr7LCjxVHfeUpOZH4NolgEHhSa221RbpG6lmqhG8Br3cpMJ+nBEWRGTqzzX
dkHOw1m9B1BFB8BlZ1AePGGoHIMkCdZRgrArbQI5Qh1Mp9Cm4/dZ7rPpCB9e
SDTyAhviHEsD+Eu3Ag1WVDBmUsz/oHtG4jXZ3Mhr0tGllwFVjYZPxALOJ7a5
Oe5nb6b7qlaSR9NUS0/EwBLTC9djggdC1xWRrubC+Duxz2eXNFb/0yYiKlko
mQWoFegv50DStkNac5sO99psTpRrNtqT9QthZIGtqQKttFDBvqhgzh/yCOtR
hqFfxOAZ9v+QD+ycDcNPPwgHA9TtjoI9loj+iANe7p/BuUamMiX8DmsUibPb
0JCNQ7hjz9UVtv6yJ+iPrLT8ZYlhvFCWl8WzeECofbThiRcHcMqs9TUx2vN8
Nw+AEsFq5RPX8+JLclPr/4FD1bpkxEYpFZPU9I4DB0EP3ydIESRVx2df4Vn2
AcKcgBA90nXR8asDxqEXGizQAp50qHNZ/P+M4wmM50U42I9nxwPrBfyXNPpb
o2XITAj/9fsMwxE4iRTVekhxIAH2EIp8GVnC4QI3g/11bTPzpaj8iNqAeC7L
oHlp9OK4ytHYQLyh7i0buUSvxLnUQPzyUko5m4sYGjLj/kZrjW8R3RVjg7Zj
Rj5w0MkSSFLziP9+clDAEmfRV17rqtkB6Za1PHLwXACzD3WcrGks9h/Sd4Yl
abnKKKJfca0p2amkle1l0UxdiNvTm2a/oUCUiz6uH7rmK9EXtGaS0P8+ALXx
kMPeX/hLg9gp9V85krtIyLLHzkRksGyNvG+skvaaA29TeqEwzH1aU/7FnH+e
z8LPKAttXvDI1s4CM28NKhdCE/qIZWwuEFyTok5QJoSlP/S77ruZG0BzZo+f
jCRO1rzEwZnRkedyjHZg5WY7liGxC3b+qZZ6ZlA7SXZTZeO95uwAki4hhjzS
ahpdKh6AK1nd950M5higNLiX7aT4rLRTSi5Y/FXV89iTpJWbfKiCV1z6vjkH
u5R87NsrxOFxecI3VWSUgVEr/2pDJ7x7DFuk+Mgd3T9Jf7CMyml5PZE8AIcd
NclM1dr4bwZAnzMWNWac5aM6Hs7mOy1MRcXQiSGqH1Wf71QGNxtm29xhH1MU
IYeqCwrunQaAetujYsSUQBEsKAdHDXx49gDjr0qFVi1AcWP4mBlQ8fcjYQL3
YtTamwOQhyaiO94alrcM7E9ebN1nZ21MotSAJpZbwmaAhFx8prSMKla0p/V+
3uGK/bBtHXVwRVFOBMpdNmD/K5q6EBB5paI95eNuDg5VWDlFAeUNgr0+g0H3
XEvzvQdet70CsYAeqI7BTvzewbSeGFYpLuvFoH9PYeHhNswFFT0ciYd7evtG
TQYGc8QiyCsEV1D8sDHL+mfd757ru/jSQWFXdYjeOQWoqFOQB260SlYuJVU6
T0aOtlw9E2WJHH2Dl5R3ztpOodcyAwc6bAGMKxtWQ7tRlHyCZtDfwj2SxdfQ
MT6ZZW1J5HlMqfg6SdZ7Ie2ps8VEfObqgvj8fP1u+HQ7cb826oASLYU+mr2T
rStoo4zdBsP9xjteOL65Qo/yd8dMzQOvz7qPZnSAenxfqlXmuzcM9UqscS8S
kj8PgNTWkIEx3FDWafqO4jifDYd9F7Cw1GgcVEeWug36mZz7t2gTObdpJ3M8
TqDCHFnpe09B0AeDuGHH+f/HYvb02ytN6BtCrqz8UeMqu1NJOOxuoBGGRl6T
/9l8C8qia0TIleD73aouo5AfSWrT0KrDmYpwbLUarjlO6TMsmtbyssju70Ay
jnLPwq3686fsRkEYRxsZX6TJ8Ut/teJrbtjJ6KCB93D8b6XWFaEHGbOWA57n
b7XPHnW4DjKPDgAVtzf1Isf/2yN2GJhnpO6tOFrUPiVBKjtK8vtIpOTuC7kk
dNudC9jKF8OQsHRcbJ6cn+pCMK8aB4AGmakKM4sLKGp/GOXIcWc1ptOeEorf
E1aLA/92RrOSAbQmeeNoJeVa71uW7jpXfd4xXGC1yHv896tITTYgrVQ1diY1
f1J60xJD6ZbYnll512MH3bxQGEGV7u048NhOdFLMBWgB4yTinNZ2u3tGl4R/
pXFWhErpAxqVmrkPLOjvuWq4VhavOMHrKhkc5bj4QjwoFp1zSO82492/3ex3
fbR4Tu1XeypxRqZJ6/SP5zkdkqvw/Ch+V4XYx8M9ASy3Ia4W2zpqUo2qq+WN
HMWQw7xBFP3ByZv0AmhocRqVcQqH9dRDvXh61CNG2sFcNzLDBW2sv1lf9ZuM
jFoAqcIjlDBD4p1hkXQmTc8Td3xS30AaAvsG6CnPe8w3mxrnDawoo5Gi0b7w
FxSDKvP7NDpTAKG0o6JFWopjRx5RFJRUki661oqNEqWDyfU3IkfyLWYJNBlQ
V93oCedw3fCeN1Tf2uaIyomGzWQcsQGWpzi00E0CtEK2w8qpYEZs3WzvpuUR
HtOoM3waZWgkz0NyYNJzmp1f+2gOaEhQ4148F6nZL6QV+qYcSZlrKfsPsAkA
xdE1FkEhQXpb/XR24RN+Trj6ugFjP5O6qGQy2huzGHQXCIe6QqJAFoZGsfbX
G8SuPtlCgtxI4j91clv2VqnheTeHbYQ5ka9gt0q9E6vJw0tQFbFPOgIiCkQO
cnCcB7yqI5K3zsIq/ti8E/5lrUfNngVhw52Yv64eg3JHWuU7FFzwungPcUyf
1DUeMk/oYMemsr4NUWKV6E+19IesgCpSOmcLYREAyCeDHsY36WlLHQEzNW9Q
NKwKTJJeU/RfJBD4r7fTYzar7Srui/tLNiJpOo4P7gBR8QX6en3ppj4Fh9AR
DeycNdVDCsG2SfQpi1VsHSX2SXUo4MJ4ii/Z7/KX4SbqTFDUTOwTbj4oRH0c
yHzhnQr0Yh38IMToPJD3o/zd3JtF5kx5/eNR5o77TLw0cyo1UfAQm6TAbiRH
Djbc9g6mj+Sfwd5s7Vql7RbWNzujFoTLHWDNiyQ9H1IbzE5SrSVSqhib+rFk
148uiEyJ3mE5SvAXbak0XO3A2uXUy7kiavAxe/XY3NKcZSxlDEEVItjvWS1i
CPkbc4CeOreMMPEL58JZRt2kPXfsHaDixoNDtMmZZgGWWPX4XYxwh9DpyLcB
J+hhgwPkts7IAtEoWlV+0r2zNtrwM130RL5xass1qqfBJiJvSoYs9BueKaAR
7gRMO39/sBBHRVXAt/ZEhZiG7B2YjCenjH5MSwhfTtxqsyzHfbsas9YtesOq
tXiftUGxgb0vZZ6PXWYa3Mi8IEFWO97GIw2VwiUfkUSae+z7SKkfxqZ6zhf/
y6+41RPnmY/aq6/mfBegMoVcZ1jkasG8UiFtGqQ/KbPHs2yORA+U2L8HyI8x
il4ljVte1ylDvgEgzcky7ggDGBY/MGiO68mZ67KkhKHBcmVHJSkffDn9LDYu
jI24TbJwELhj9CfEsVVjNLnZqEodkjy68AYVISWJM74ilMgeCM3xjo5xc+Bo
0ibu+x+9hOAZVehN+E8KIN8BvP/VSKY5UwbMOcO8/m7Kil/xzykA3lL6Z32c
fgxUik3vsCMzZ6GHFcKEnjQRcvRszP7hGuVdYzgZqKeu7VyRYB1F+7r4pv4m
pc6X+5DATTvSHryk+WKlryzT5nrpAUgALmuVV2uB866XCNQ3o8PIf7fzzboH
9WUG+tuIAUjyyTIyp2eBGu+SSX3IxJLyvok3yLKC86xWBRqWQju90YtJ+Wa2
W+/ycoiaN7NkIE+oZ2QqgYXSWmCqIuOzbVWxHk068zbZJXt54YhefaGNmr32
wZKktLin+VBMYcxLfMaDo1Z28trtDEuryYMVoRUN1TQ1GPY6wWyuq5Jm/9fq
pPxuP1IbVjXbTjAUvrBFQ28f12lLXHOodagGT6yvQLLcN/JTeUMJTQ1N0mW2
DMKXv+DqRzwPswlxyXbL3qPXTI070EILom1KJlXN2zH1LYnQ62elbF8TRvOD
xx2jxY0y0/JW08JPTNvxOCumDbXytWMnYhTkOlKHb7jbn+Mu5WIIc5xP29hb
1bjm5g/dd1p9LjlX97Q1ePqBRY9b/1+w11Qu5eV4QqLLJe6eFd6tmnufAKP8
eJz9m3hXMYo+qIqyp4I5/++j9ER6p1xwEHuwi5KWG8QXYAr1vnrw8+iY02fO
k98nJZ/1+exU4EPn5TkEROY/2ETZTa8FNfiG2b7dmjOOt1Tfrcz3N993mvDF
vkuoSHTlO5yqqV7l+s1nzhhJN+uTwuF+ze3/LDBWA5iwVTzyrvNzwkTcR2w8
9XprZrWYXsRbdfr8MreZsVdCBu7QruVwrqCUZq0S+0kqasY3h/Vmasi7Xxuu
a4eRbBSPWldr1Bfi4OD919bRMpaQ1CoEBN8esFruieOtuJAqafrF9S2Ldkhl
RSZY8u3JttFhCuYxQdZgnf0vdSUUpnw8Qtsw++HGCzYf46ZYj4ZnfM7+XcFt
Kd/hvyNcEgAx+0UijMNaczzbbjnzKGj1kd6x6krPeANAnh8q97qNjUE7K/IR
IqYxPodWxHXIrr144C5JlkgeEJ8iZI+mlyuebpEmpoBEQ9q7f/bMBd/+2G9y
/Rki4g9uTct8A0pRDbRzDwDKgHdfU/CyRj7iKju5gxvq9EdJbkuDq7vh9suk
5q7yP6ds3uY4m0qJbBjsHeyB8PZC+LxpcwEpnv9++PzdC34Hwk6lduxJOB/B
CT16MTzFt8KPujTba+106F8Ym0C4IoxNx9nthGxAaUlHNxYtDGMyLgxaiuxp
QlUzFEOnUopbRcY13hOkhJHiRS6Q/C6ibUPIzEPyM+6Oz6L+iWh3DiSEwI7K
Tc7p/IoucHPdMPLBEFGdq0aK6T+muLc51wegmVTT94pk7LbxCxlSiHILVRri
cRrH1ujEgMKM1huxoTyHDev5bFD070vWIqJX8bXWx2LIJOJFROe+ufj/5C+9
TS36d9+aBTL5Eu8iekq45Hoyut8jaoQwy0DGwkHyjCrsZezq17qrzk/Lwpd+
Zah+0zbQ9SkQj+rzGBWfeF3i3b26Ax35gPOAD7YREmitzXpgQH7BeChgWDYH
HMJaoEhjr1QCsieGP83nqC2fSWWBY/AfjJF0VeZkylZOyjJLkcEm2rYgCuOw
ioTXDrEXyI0Uyjr+mtnqlWGd2SsDX/BAF7L/sOyCQ4wOE6NEKSgaitzoPlAn
ak+DHgiPIp9h3rKPAPRPlaZP3iLoSAnAR1UjAhrqQUf2xctZYZMdi8f2bq0X
qkvlpGIsayhWQb9W1y2CX3FTAgKrx40KT2M6MNDfbCo4FhBV9muNrqxVT2zj
HSpovX5jqiFmQ235CPTr8PPl8TqceLf/t0Ih4EugfllE6uiEtU6bf7v8d2Fo
TvpFdu4heSyrfqaowuyAZ6vfmUfhP6Qxf1GixyJWO+mLTw+pxfIl0WDYoLUm
eHLO6iCLy2mkq7JlvfUg3unhaAWMDCEq1kczCU+UQ8oAVDh3ZouwM6iG5ze4
RsPT/qLYtrnbzpQQvT5uHHbVIcYS+UexeTCReZetHtv+/hCP1zZFvAtYamsP
7bs1FJPtEgw+EAGnAnbWhf+yI08I1d1bIxWGpvsjBI0t5mf91PbuK3UPYCQ/
bot5qH+ln0B0VQot7QiQUlFC/DJpNz+Z7UhxrkXqAiuTG71O4YmASHRtUkvT
I4ZsP6aGzsVgY8E4FbSKVjYybBlL+C+arel5fDhrP/jC7yY98OrhfkRbUmlC
+BsPaVRZq2zoMj7D70eYxUr1/FvvVKFUfDqWG/R/FKpW3aB8u7oCQOTkhEx8
YfY254O+OpCTafGl68gfTjH5R1/W6m+xUjRwmHZnuxpJllDIfHM3nDUIvtSn
kjNu+6Q/05owAX+2YPeblylyb8/CYO1bHZOeNNeku8jqzT78dVR429l1jUR8
hRgRKj7rDQ0oVYhFVod4jfqUvirBy7u6oFFemIrOTyBss9sr0RKCGF6XoEha
lp3vIpU8d33o4h3Sjrkpl0SURltST+9eGq6Id/uEdPFnkFTQnna5b070OTgT
4H+fWjwS/Hp6SE9UgMY8I/N19u3YzYWSRUV7H/bl76wc1nW/mOWlSvPfKeeI
ooY/U3hFBstONcHbXlBhY4WB1wKIox/EPGbVdr0ARCypX54yWQn9tae/TbGw
Dt+9dIzJfsWqk+TJuIq55zaWseh20G3vxiuu+m4cgumZoPb9hsqY4FrCYHTE
n3o5swDZUr+tV5Vzl4kLtj0/oh9xb2qklEeT9zxKF53QdbOFZ5KBqo1RjbpX
A6qBz6+r8e71ldCC0pCr6b7dm2fTGiSnS9G9MJsFiMG3Fm/HGBVlegweQcSq
ZLMiBpe5Ct0+lPczZxqqleHMjdVhVs0T73yj1oawiVfPWQIVwWSeXvBGsFTc
FjlbxYBqBHzqqw6XaS7MNmeTjIACDaVsjgzKJLf46dccmDE8muPRA6XeblOp
oRLXZ1xOcXcpJR8Guqx91jPx9CBhMVRxEzmQ/K6HFZ1TalfLmxO0U8Wi2Zwk
Ts/HD1iNhXFP3Z4fMMY0fwos0IboXTIUxe+Lr/gP5ME4fl0FnP6cMZwPwG11
KBNGcvASySizL7LBSpkXfjuB/ttaRxPkQ6dKF19LZJokAcZE1aoEYfTVSM9t
GNq/ZGsmyj5qdvrwSLR2dHUJvY1XvW+sXdRaoUvqaea4m6rKK9ODiwwe2fzj
GtbxIAD9htGlZ2BfijyDDpmOivfYD/WcSrnvi9Wuh7u2aqR+tkF4Lc3haqgW
19vnAzOfCBUhGy/a03dcpPr4gD/tCgaPXkc4QqHwwuOVXFD3zR53M2vxrlmW
0RVvcS7effDzgthBJtjqi6x9u26CYpsuRIENQ5oNzhPu1wDInNwA2OOAMUro
SVvljI8iWEFBkgaqpczxNyGXiaaxVIHTvjaX6ae8zsUzyufbAkGXWgfkPvQk
RWWKyIrqKdqBp5VT/QqsJ8xHWs9NSddR6OMn+5640Y15nbcsXp0mql1pOGWW
zb0PzkDE1hcXLx1vrqYCGKMOIP52MSBhJ0Gk0h4ZBbi7MKc27eGDVR6D/vQ+
o+cQo1mSuJPuRWBnMlXNlSMgYCJOFJR45IctTJfwExteNO/BV7C72t/bcEC9
zKv+ypXiZM38j1cOnlr6T6TNP4e15l9+zYkXfmuu7Q2JrzHz84bMj/e7JFOR
1s85LEIsPrdMDdmiR+GaOWDUcbMZbEUAYEMUZzQoPHpVQgGrYSLUMhUHYtBr
Lh2hnC2Bp04C45XEwFIsps/iBld+oPgMxxoC2CP48SvOb2o2D8YvXekD4ivw
MnZLTyz33hWZXW/999RBv79EpfB64o+fvHsxvukwoBGJJsVqE7pHo/ikP2WJ
GnTztiEHOe92LYYK0JSt8kig7zQvMZEeuW8EsDIszzcwnUzQTSsvGR/zTzka
ifGPvXdHt4FRFUi5iyI96m6eXPpJgdne1R4mE9e1j34XHJvGuK8JVVECKrCY
pXHcuoK1xnMXLji0rBvXZbcWuVkW6iPtRy8s5KHy3ajwO/n+plvKC7uepRew
YVdFIFim903b6FQ9DrQnYorE2Rjk4wB7LGBV1+ZVmgMPW6IQB/bvbnivjFjd
e818rlEGWgW9AGqkbW/lH1I8+gFWyLMKWKd1+/odOQ5rIl8j/Cmgo3YH1/AD
VogXL32OlC+KtpNLa0WSNjE74tP4YZVmEpVaOGCD/IUXNVTGYK1QSQg9aERu
1/zqf2K0pnnO9wj1WJAswoEOddzX05Ano3Q9W5oa9nXiJMkSmqnU+o89IQ2c
VEm2Sss9ggkHW/WPiG8TLJ/iz6dGI4yRc38WLYJUGIgi39BjJiXAJrW4mF9f
DbLAVuWo54F95kpNF5vRISoJKOdXSFE2yUygbnn4Dz9OERben8U4fS4sBua8
ulOM1m1RPObAHCwnj2/XFbB0uvJo/A3eLLbdfByFvWVtW7Tj6LvCAa5RD+iK
OWPtdNM1a+3WcTsx7uQJ9y/Pvss41tRD6jM4jtm6PCXbAIilnbPj9hT25yEA
GPRWj7GUGXU/DT00PT0bpXNC8ln0p/1U7vhV9fDkFX62lfoJAGCKkpJfTxc2
AzAfQ1w072Jtg+cEytu73sNTRwnCb543HtikefMleLvsBkquNw+rjqgDS9aK
9MvkA1DNeRnRR/VKYlZeh1MH8G0cXO86unDmcjhJeC8ztP7gpugq53hzdTG8
L97TOMkGvvrASjNumt1zOqS3frkxIkf/UBBrM6MCtB5HVicIzSZdD70k5nQ/
RmBA1NhJ5iDEdLM3dtY99u4Ii1CTeEvdOJuDoiVOr0qO6E9wfDnz/XHr6+XQ
AXz+ZjAF5gcoUlKF3xb6XFkDHn6iacJAIX9e0LxTRhsZ1gUC1nYbDT//1J/M
Z7MCGIQDGp6MORQmaW2gd9mER4yx1guUDjcJUoj/IR05JOYipnC0JlMRpDCy
Ci7Twhu3FzApjvkBnLCdipsljc7MeQDx1mNLL7KaoJwvmXg6WUiVYu8AsIek
OTujxWZ2aVQx6atMtwd6y30l5bJ6ejibou51tQ+ogV8L34+NXthRCjLqtyjn
8xkW2atG5ZA4vX2fx7F7oVMYm42uPrY5hUKF4AMkefpiIA0/i1KeyoL/KOmO
MeKVB1DEslXhsQm6rUlDalSiKFTfsVx7YO/ZhON8MLMeGo6okq1f9MXgJwJi
W8vDZRYgBWdvowCZYwd5l49tesRBkFtey7Q22T3/+qRtDj6VKFJqR2PYdH+z
C2HDAbTNnRCNNLuZKyd9ciwzQCisX6uIPIkfmEoMJ2uxXbThmuaZRpQZqJCi
mSRriCUuixJcuCYCC+LEhMlwueA0qj/qC0sRBsvyjbH1gsFJPY8HvfyUvyl7
jrJGFsXnP76dU5c5vyIlFJdgiZ9w7jhBc7pEpoFHdNnz2n7KKg6hC47W/7SU
zn4xyayEjICeNDX5tHse/upWESBMH6y8w+Js9UQLqO55Py8zg1acMtO87v6I
cDUcZs+vh76jQXMY/CCxzMb6pXQXWvMas571/RVlYM744B3HbnSCvwXpEtC6
70xnNOP3v/KUpYnNE9AtxJJ7uhShmEZnrOwZdQmj4z+x8iGiomK6Eps+h8ZH
OohfZ1N2/TMcNXj6qoPfwGiq5BXx3/gHQpZa/5PpFNdJZD/gT0rPm/k4ykug
74kj9nd9+kVtXq+ehbUtjex1tfBDO/mZRaJvkKYdQsaIXIp/nQY70XIAsUfh
6uQ+BQ07ORWv9Z6pd058TzWWgGBkIgk8TKQESD4JBreya+8NLwMrTUaAzaOj
VimsmxN0TXo4+zQDp4Zx2mli970t9DVrfHyLZqohxj68zSMcyhUhgJYgBaWQ
VN/GlDyE0c4EJEPbemxR6txI3E4l2eCtjfppo8plnetLWEqk6wlW3U1ol16r
SWkprLplHCvywtxmlSyQkYAOk/XCwSVD/9rzqcziC+WuM9Ll/uDjBcdG75G3
E6VWBOdqEW9xR00aOX8sely98X7BLta1aj7PpKaqzrnLUS7aHDYFr8bHcd/T
JhCPUh/apVFX4dEaXEI8TBLIOuQaz4hS65SFUDzX33+duAdCgJmZrFYVj70d
QgZquu5l2yLDn6i9Yn0Tl/YTd7G5sHA6TY/jLwLwQ0o57+j51YKENLoKYCzX
nuifGN/uy9frjBTIHVtpvitsyv8slICBL/5F8RWD0Lj6TqJZ20x38cRtkIuR
t58sCSPApVVhPj8nhT/scegLKLDVAE+YwT0xJ3QNXAkdEWLHVnzHafcVyRN4
bamw6bTpWqCfLLfobzRQ756em0NyyPXeM2DRr8p8m4YvLcRuxSF0aDOd2Q7U
GTRiZla7iRqU76hH7gm3rOLgbvxEBiZvAIQKdI5X2UakN375sBt4ginTzZXX
8rOts+FPxN+kwbVOWysN1CFrbcrUOxPVTVKzaNCFciP9i0tDgtT49zbZOsge
eiyiEXK8iofwvwRvE+ZbDUCC9sD2F0nDBDFzL87QEHP2VOJS4oErMJHWgloL
A8WY725PkcI4wLvsdP8ivj2qgLpvCtMK7u5XDIPo0nPBUviuwGye2TIRtMxC
/z/fFwm0OhyB7e7CwgAOgxlT4zToCQ0bvq6uNP5VLRDG1+gI9PiaTsaSMuQM
3sgDX7ep0W5g1f3XlihdWOBguuLH92GHH1wlaRBfV+jGXsnYYhLs7z5BDrBx
yB/ifx4u3NiTbl986bNsP+UdZHIjLfzWUvSeJdkH75RT/m/4qdRm3xzqCRM9
jTv9n3bu2eH2CNXuj3zJHZrsEoJuUnZcKlkWS9FluPcLmKyqA2d92j12Tws+
aW02W822bvSBVnBUXGS9v8JMbq2LmyxC+6YW8/uIBvuy6JABxmNuVWmw9SoK
QaxOjg0nzksNVuUx58GOgR9LO2924UPLN39qubcQEq7evYUx+KikUliQAiXz
1fuZvL+D28rdwsGB3ShWuAzvqCxIwxjvRmt4F+rDF2u5fX+VLyGWDT4uSVF9
9aIBu5pSdKtnnJ6d4qXzUGS8+GqBrGXanSy7vzQGLciQGK6eC+yaii7mqpho
yFJk9JwjL5uHIEuxeH1PHjvkPg2C/GTPh4ep8BPg3mpBuWM3n1pKk03JiSBn
zYjWr5TzActh+hZE1eL5Y6PnKVrjTFWp+gHw0Hjv1apJBjcAXScwHGTtvL8D
CmlFdqRHDnUCiZVDuCEfJuLLnLBdGIQSSGp6YxybyeW3VNy2tLigqB342nbZ
lWPeqCDMAGZvglWhuxDsqUr56BLXI0uPnJvk52zEi1BIYyS0XVMpwRn6rh1Q
QVmK3BJLGhMvgJ6ewou+oNz7r8rFlJExe0so5eYAk4i//hPu78iOtqzgqvPW
e8myfV1Aq3FcB5J6Y/Qs6TED2o3P3cQXTGi8XF8EgZ6MKPAKqprBSVtEP0Ai
yTDpCrDyLt1+eYnnFGcNB89ZxniJDio7NzgIVmvGK+JLD5n0hOw6Phg/hhzq
YSIVizawlFDhHMty4HWXqzSUVjaMqRsPeRDdymzJzTnFK2pS3TVeEJcxiD0+
ffUFMyoMvpBTsD2j63GJFc9aIg19+OE4K5nd9C4Qjk35eGfstCJ1HSf/WE91
6rf4xayrN21H5CEUfmFb3xDU32rezeWJlYB3PEI+ut1Nl+ZHTGI4PN4fT9v4
MIgvKsfpwjPIWrYsDkSgF9GZT+JdrFyB65Tsu0UFhxg3moSOJZsA6FqN+zQf
KuGRri8WEAtbnTio8GT7KBrt6dH1XJwoyhSFs9t6vrp64JEfZpt0CnZI4kYL
UldngnriOvCwjPjeYp0ZJQEGJt5Kk+LbDktkVHi4GVmH+xmrAgehHzLqWhoL
sjsYJGLy22HlGO5Exvu6digAHjXVLoW2NGELt1sxI0Y8W28V/HZPu24bJ7AL
8QBx1nGtIrfhRJOPLotsqt5upw0OS7XoemLKN/J2k3+KSzV1l8J7HhrdOTOT
d86aBo/rDQgkrt/Kg9wA9PunHldd+D0dr5VuY39YLnlwnxmqGpz8cBe3vBcE
ARUkgBcKDVVkLkM1QKrVjxSz9n5ZM+AUx5ZV7VkF9nLKfQLNEBSl4bSIZ+z/
n32CaDMLw+qb4U8JeanRO5EqhtLAMsCJMMfu/xvHaMeyLOkKvAaz9QYH/MyJ
yDNwaEEawEq5Mw0AgA//+khY9thx2iU7vt2bJdAy67tuGZEQZZjRj39ZBfc+
1lJzo2+MFFrgI81hSmg0WzaWLf7ZaW1G0VKSXSqRWefVUPeV5GtUVldtitFe
BbzAwV+m+z1DZNXrD2eHsYoe2f4I7anWzlJDcVOvX2lwFuiZ/jwUr2/z0Eqq
+6q8deSoMbv3y7TwxZNjqgMJQ3S+caCIBfBIKd1KFlq/Yl/30Cik5+f8IHnW
69svtImB1r9CtMocicduRx5eYJWNmFq+xp8ohN9kW20UCcK1JuBGwe4pBu5k
iq15HoSfLq9lmf0solxDFT2Xgeez69XHpl9MPXy4MkRlJuDlBbEXUzLSYqyW
NtpzVS2LCF3ao46E/uuZCVx0ZGbNLkZTAeXPflZBdDim4Cs3GfN75zhgWLde
pKogAtT/pNUibhVKzmV28dkIkRv6h6LhNp10/G+YY/dzZb+RItcjdLz9xiCM
YMhqzA3/0G+P03XpLMHrQC1kF9N8eRiiVq7GmPc7RxDD/VGnWmE0ZhZcQ5u0
9yyfUGlEsbHnQwtvFVe/LVEC7S0NvVDOyqr3aQxK8cGk6KyM3DnBaauVAlWm
N4vvIFxpZYOEcIhbudR9TczTFMTky/ZPdQh4ClJBnp4XwhcRnJfCuiVjpShm
oBZ/8jFQYxilybjNP2iIOU/79mOxA7fS4woHCQGsMJFfct6eysztfBXjkwE1
hddZyBHQHNnUm3NHYgNJNSYiMliBGYApMZTXZx25hTgoqotRZS9+IQcZlsbB
0lytLR0iHSzlbA+yPuOIR9vC3oIvEzFaIZYqcQ6qLfM8g72faK8G1zte/Nl8
DeLZz9f0crOGeAFo8FDdi52BQ9ep9fAC2ad3Eg3jvGbCHtnzkrqBEsJ6ndre
0K8IgDo1hvCTZ0Pnv5nqXkxg5H7FblmWLrl19u0JQBk4lLgIWlS8TwxiXyYX
lCpYhB2LRpis3k0kenEf9d6Y6zG4Fc/uK1cDPckk+b3Dt7ZIcQyhmqR15l0f
pkDrGBKmqlswCCNcjFJAeaNdz3a2YzXsJy7m/HfkNROXcfSyTLUK79ib5CXj
aHYg6+4pp943DYmfe5aPiNaFH7wIVG/l4/EeBe+yC/yJOr5Ex5DBOEj0aWUk
gjL/IeEKDu4bhRGZb+1d6zTnvhVQWLGQZ4hlphZizHqQ9T1cFl26+LHOJQ7A
zzFmIgjQICUIYu+rLbs0VUrZxpMPFkIP8FnKxHg/5k8zAP1dOnO9sgwcPzZ7
me9OZwXEIYvWlXP8k/GkxMgdi8+7M902Zh+zdpM6c2EdrakyNmk0NC90guhB
VkBwqj8ODpT8F/nWv1ZjMMAHjcDSp/qBPDbIiXiGOcuQKmRnJDz7lQ4IX3yj
WdBPcRkODWENGkXY574XYUL3jDoxWxNJ3XQ5FQhaxXbFuG0Rs8yTBqUrKwZg
WcciUlGMtKtenJNLFGCqCAK2JD9FkH6jqcVuySq1EgUziV+rwm4PEWJiT4yr
z9kduMY1XOdpfI7uwAkZiSxLvx/Eiu8x91aTazoXiRS86wH04kyGPCfS+v17
aEmGNt+PX5R2Y/7NdfkihbYARYR/SCkO5FAZFDsD/lsBZbvPgNPWLy4hjLP4
DaA0UrV0WFFHN2baWHWrkJeG3ZYe/bTjWUK7Cg+0/PdtRClHQMKt9kz2ZqKS
R9c9Fl9UBGoWDVJIVIoKr8cG/KtapPgmF/gCWGyN0r/kHNepRLFGhLOsL2pn
Oznm6Du7kPhXrh1anVGq8UceGfT5raxC85pQfRrAUEyuZ+C3eUTwxi+L5KbP
dxu4ukVIZzqhkl7wqsFBcpADuKr6uXUGOprDEZp63la7Wzwzxqn88+NWcDEI
P8fPB+JZkC0choXM+W8ZZY+4ok/zcK2n1FZwDTy1DtBINwEEkaCpZcABcQfq
0cCcq7OC6KvqZByjEmELjzxFMNRkMYCKRo7uqLu69aS8qzK06lq2zrBrRDDy
N51gIjWfxH+w9ju55I/dI8Kv3h39AxT973Xm/fFDtuK2mK1Vl0XAjSpfv1ez
f6NSLE4KYxach8pCJrACCjgdSTsj5vwq1Ur8jXSdptpzl9KLjRsvUJqj8Z/x
desw8/A1GchwwRiPD/HMhdnzpLMnb8CUUZ0SfyKRcD1A6saBuBkxRwMTzNa0
FhwfWygiRLiN62KwqB2GsSngdD2AVVNw8VpOGrlmIzeGWGTH0agbwBQr9s01
Hq31wwfaeHsUcJB19mssygu5A5lhA5QCs8/pt4JOEiwGkhLZ1/cuhAXVf5SI
3jOFP9t5iyYHgdUy7z0B3SwGpi9UkM+Rm6loU4rXvc/f/3c+jezToItuUozs
9jEE+0nc0MgHMYlzMqdT+Nki5tIXXgTN42R2QohidehAGkssxxma6ss3ob/8
NiB/ysk9CExw85hRmwhBmTqOorZdWvYU0BE7xCurm9ykVbH1l5pdyLgiDNv/
aFcomv0+ra+F150UgmbY9UUbbR7ijg/nLRFPxHWrzgLH6EfPFhXv7dNVIT6E
KajXApn3jH+htZdtxPM5/EvSkC5Xg+ifdDVF7iJAIgpZmBOzf8RR0bu13MF3
a2wl7K//dQLP0tFnVxoatDa8dqSppAqYy/qF4y8XPeR1QXck88L/zEyMWcWE
lZLWsX7ey1oiTYUHfcCBOFyn8x/zEwSH5p/Cffft2ni7080ckGshCM20Y9rU
0t573jyGd9l0QsM57zRa43WNfC08Yvk8YXtN7lJmxKmTUD8p5LYQrFDFEv1a
rNn5JfjGyIXx3l9gc6cXX5iBgxQn4BC7uDz1/P4zAh1O/2ZEOssWEdkKWlwW
M/+GNU9TQKPozW9pCHSWAl7gi5Urr/4ou7lLObz3LNHbNmPtWIMpVZrQROqV
0LS968hb0PLj1XEWEXRPDuGEzLXcya7oc/OJ/vPosgwu6o0pAGkmgQSle4kE
J0AmHX1bk6V1avV5FeHlvvvR5wdZgtiJ19QvTkm72QvicqEyGZz08DSzoI1v
67oo4EpZ2xdhyQ+g5Zgtz83SWNY3SDhkmUwTdp9FaACNXk/CwqD6oM8i0xBX
aYxccMmaWL8yJ76vlvuiHLb52veLEmhmnOsynXTxBXEcQyoq2nW4p/9rht0z
rrMQn/zwSWeMYN7qnm1Kc0xJ3/OdUtP/gH97ey7KnfqUflubAhgwrG2FUOhj
VE14gruTNqno60jCaRJc/Dh3GgUkZm3ofJUa4JzhVqRUAtjtmEpsP/lqoL/b
LiQfcR4HRlHZ97Halu6g/N7jCVmxoshCmy9VAdXJoJ/7gjnQCbGmL8ZR5fc6
tf+b4S0GyxvO7saYC76Wl2HbbKwh2tOv0Vhg6qy0Vs8Y/0D9WCBGfBtIezCQ
cyu4NYrfBCv3XxhtoR1C3zs/0K0IKjlIe8VBPr8yCOEC7DE1LmFqI0McFzyD
nyV2IU+HyRuGdtIBMU7DoqI/Os/EqqkkSalpqcCtQmQR1jZhTJCR52a7w5jX
tQqcrFvxu/6qzKDljbo0hiAJ5/ztYxwLYT+vL6Jwvw1cPJJ8r1uhdUwpsGRR
sW7p/YlyIXcc8ianq5HaJLDik86SURrrWekpzIhSHPsWMSjEpHz/EwbqzN96
yDlFE+yrRtGQNpgJ4tq9/zfrX+3yQClDq9ZavrrYefrm+FWNye8+f5UNW7Zw
Zuiqz5sgr2z2dQl4J8MdQBQs/4cZwbcjjbwJKG07qqoZ9Oub2wLZZ89+CSHm
Itobwmqk0OS4/VL66y/NBA+qduGZE6Y0hLWshZFdXe9S5ZDIsBBuo6+i1Bcg
w80dxAX8OcrCjV+ry+Ei5QDMeztIRdMRVHaYxFs6QAJ4gxcbThTrzAN3N0ho
ICzu3aerMPe+gAT4ewS4Quqlvw37q+KxXf47pgIltgeYg30T4gK0AEuvOCCO
sCtnBPP1A5R2L2QcU/nJFvky1jXauI1k5Emm2n2jqQnpkUnkXvVgJanOMJhO
Kwm3lj14y7rKusxJ9q5zEdW2s8+BvvUecxkjRq9rw1lYnBvEaOzrFbXd49WC
bWLIPbBiMwEg9FlxS8+e4hG2N9GZadDbDLNGyyckxTZTRHWaCH6Vl6jWprRo
r3WYqT0JY5QeBDk5qmOC1hUoHSVANlxqtmmpM1wSdFRz38h3vPBuzyug0csu
7cysvWEjHIGZYWYmIQZhulS3/M825U+9hyTnZJAncQSrnZI7Fd+ICXuIVVyf
a4E0daqciKRXiTUfuSvErq0AsT8AF9WCBWlqczZA8nyadJw7+fUe25yjB6ZF
EB46I+IsQognhYBwXmkHuflWdMHcnEP3La5aEun29Acz8EqJ026/hsJaglUQ
RfLI7mbeNVgPFWqD6BLDE91G/0WFh0vltkKvg+GoaJL4DHm1cSBymeSPRA/d
+rSWeqGWA4ArVqaoBwypmS72oWejqf0y9XjXn9dbPig3OPzJWFR3eFZAix6L
uAfS5+zwgJ0o50Dg0Fwe+xolJxV6yen7wcAeB+23qS4B2c5Kcjet7SJj/0Pv
k5cXGdJMxGFOUhXIzGz/HquwzcqbJyyGyr+I21XhnItYwW5ZzaX7josF/wkZ
ID+6GrpygV+SH1ig2MJON51z5kPgkx41lfgStlemZkoIKOa/axTMsL2a/m1L
z0ivu2TsAQX8oZ4tUzB2TsA1M5bne/V1L99SO3qlgqGBvb52VopIkgEWqvDP
BB2MIbRxNVDP278UCkC1GZcYq7FSKiXEK6ljJK8BCBzXYxKc53XjZqHh2wg4
BtvUBjzsJombGwoL/LEp9dfsSQqBT3IoghYzWFoGgKJrC8WTz+SAnw+zYPPR
hnY7HgMTBdaT9LaIHIMVhfIJPauq2El38RdK/sxY89ehXVaglTaV6XrNXxz2
3AQ3Y3DrxoRcg/Ld6eYY6YXKe5wfLgaRfsP/D60gbEsUZ1jx0Tc8v4mkTir7
dp7IuzxXXchsRnNTP1c2lrxW4k/tqkRTXNICWL9TLK0fTvedIGZAyNd6mm7i
kJduiItUJsBe/6lnQKHDsW8329BRgdu/T3mxhGlWKU6UYGPskI0Y/wUeKZz4
itvToFE+NEqjMbMG9MNnVXptizd1X1XOeS7bPqZ9xkeTRN8n0AWKstzM1ex5
yDaNHd3B/A7698xsnZy7DR7dCnSUQXVUFjEtcI6oFmmHfOaCLEbyg/1f+jXn
yQtX2iCpp5OO01c+B0LH8PskGiAvrdgwehUtobwlLkNvGt/84u8nd7++F3OX
JipntRejqtsC5iuhxsaoDgAw/YL5x0vxkmHBG50DR5D3WskvagtpYjt36q8c
6xBsZnXBqCpbAOwK3YVKVK1y2CGnZ/1FGwsknmBrF7wq5Wfg9FqmyrfAN4iF
U0MiaV3wtbo2a2FWyKqbJ5V/J9ZWpGPMvWBMbZjEQUsVfgPt0Ky8e4Qg7Z75
EAA7uIUHt6IxT8VI2FcZf18quYUnLf/CIyyUMERdwSEr+Zf0go1z+q4ojlxL
/DdHBHmFaOF2TshNp4KXHyXxbGj5u0XQYRJHA25AYroWo2mpz+2E+3pighnO
f0hgXFSw1yi9AI6W3eZrFq63aPQpJhCM568TZ0TBW+FzPCkfNhz+yIpVJ2WN
J6aIUh/taemevb/THAUcIwURDo6xvH7fQ+vSfhFp//eCVs64ExTNMnwkZfcd
kPD9Imwn1az30STEsp8HT0KFVwTE6LCHxw5N9TL/TP943UfCR9jcfl0uz0vY
vjua78QTj38wC3+D4jE5T0SHlc084eJGFyj9CAPztc1oScf5eVCY3aKv5HiF
CK3y3skfQ3YgkF7w1QvlszKIoyzhSwf0PCSmsIdeLt127udepQjvcPNBcIsL
IfvcerxAINpHLwIw122+CX0US+rLnmDSRTeSF/vcdU6UhT3/wrC9hHSZjU8T
NOtcj95A8W07JqdFRwcREJjFhZR/WEUJkDM05q4O0LtZqBeXWVSvh9UESPs9
OULj+8PCDuGk4bqhftML2uA6xImBJmpING6e2vZ5rZ+WuAM11GUMtsJoQxqe
Zl23JPye3n3iLJAVCv5VqU0xPhHCKF2EMQYyII4JU+ISlEb5+bKkJI1pbP+t
s0i3hJy1yM+v6jyLp/lEP18t1r4ZKM+jwxuNrUCm2s0yQA9m97HwJkF9dgsF
JHilThs3Xd1mOc5x4aH8h7i7FsXV0bJaIguh2P4OwYoM+85nYyou76T57WpH
Az9iZ4S+zN1UdsohVUHzwJRv78wxOwcO9z9PFfjQ6Tr3aiey18fbtKwqCFDs
jXEXc7ODfPJIYBNFGI6skVjEtdDYShp2T82fsCvPrflNaZ7fKCTHGMG6mczB
CpZFfHZLKbTJi/YHOd04IoUuTluiM36bn6dsZ++R1YdzotpT5pcG2kU3v0wA
dD6uqbprc34Fe76f4sRSpSLLgcWtGzLr2MSktaHmmYcv8mLafI9KtyU5fV5P
2t+vWW5n8n4o3JfUzp9t3/zMjec6OYwPpiQlTnhhL7VtSirKTXLuNvK8AyBO
aVtGk9zL+vDWiDImYDXvUTU142nTWHaUaDatUq58joUIpPmvSmRwWDsih9lt
r/dG81cT4Lk3bxezICKnBUHRETgUubLckod2VYXxoJK2w561AjDscYuXHhYB
WhzH3VIdUj4+J757QEDY6ykBF4+fLEFKEcjig/mnfmo3jRfla2Zw3i1fp1p4
TgvZgKSFmrClYi7yeWwsRCPeWL8RsHhuUCaoGC1Wl+u8r9QOfd2EDewTWoTL
DvAMjFkhhPGfKUd/D9SwgRE5aF6vT/Rc0u3mRnOtQNnWe9avNZ+m3fPwvnaP
EpN6ahvZRfs41tPGVBrXbi8Oz0tMAV9tVbQct0IS3qC94USAtCt8fYvYAraU
5ufo4Ew77COGva5P2AfKUjuwcFiOGj7gxR2npyYkEqSbBXotJ81rHZJZUQZl
ZVxg1UghoH0f4DEinjE/cXAb3uoV4XCvKvPT6ZhOpcFNYRZphcsTHIJ0J6yF
Gfqj06jngBrh5fIZvCvJaLmCFfvfvtrJxuqSjMx83HJiAZSMPGiKOgbLfNlX
koytdSSncdDh2AK0tG+5k7U20wFKtaa4S1Hc4VA1PJFm9lfk//VIHxnkXfyx
hWo+ZK53vePBLXGCBO2lck9Tg+HN64+HfwyVwLbY4CKgCYzbrapxENI3hd1W
o62XkuXbryCPSunCdkv5mgwG2ze1cd3MBAcbr7MiIid6Akue2NI4UzzwQU7Q
VsE6iBXVYGb1aJYU4RWpQYC8sv0Qnp1WeFsNx1APn5v8GjuHnduMozNWBuAz
nRp3HDp9XGiHe8SBPk7dkLEaezrDSVVdXxo+mn4MWGqQvvFUWtTe3idzHtsT
VRJNC+ScjrEIVH2r7pl073JGeFLpsAXrHFZGofTBQnxOY/Br0CQCWagiVjuL
DWrjZvHLruP3A6MALb0xGLIlNQ1J8bhWxLj8L2yZ0ue6qHR46k3gwrGuisZT
xU3sSQbbsMPToyUeybpb8Mk59sN3+rHoarrpf8H1Oh6uYh2qjCOOizro/hFg
Uz//njHCILmGyzTZXsf7DTPxrNWeBcbnjbPT75sQwu+rpD3kpjtQ1sZPPGGu
rMqZEfOIJR9mVgcgbPGwYbn7tF/HjMBN96fqOplwBMtpami5/MMHpyoxrm4y
gpIivGOMwwXJvyMVP4fg0OfHe/XiynuivLRd3MHQBkdfCsvzn/GNZoaxChb1
medu/aIGcwuySXle/+/4Cj3OpDTu3j6YqTOGPGokpad0mhkGWMq8j4XbYlsb
z0hAnqjrCvUgb7vyDxnNqHlWJMrUP/D9NN7FYlP58R1E9kjj0yjMCwQ7RCzf
sSR5HBwUjJSWOzsML4MNlMTcb/5bXUmJU6vOs1DSxxHQm/iv1/N0mbo1SCTH
aVLdixe1y7rj028vfRKmX7uI34kk30Lewc3ldxwVMBjmmvFLP4pJzHg08ooL
M2LXuBeG3eN9cfB37PI1EWhMZL6F17HX+6czV11pEGGY5XF3h7+3hMcY+gRa
HoBEiFqECXY+U09TTs7q4QateoKuF+HYs7rHZRa9jUk1NchPT3yf6KkMrPpJ
0cW50fzU+XzH3M+u/VOLxnMng9/83HJj1kCm/TH8+sRiuL58dRcPMyEmtGf4
3/UpPAyhoGDeKJMNJzEgCSzbTNpKlmbtIC0LXX40+NSxyfkJuRnb8KdiU7KO
QA0x1iS8RT9vJhuLgm8esw67NkuSwRW9B3C5Dn5vvlpB6+BUri8cr395HT4X
xGVrzk4IDDaX1zU0sS+5h+Dp67uC4SErNh0z4Q37yQEART5K9cwLE33mo5dL
PmMROvL43onHapVPS79ZmSLGsIMWfYuCLqPXsP4ONXm90iVbYFt5n5fkSgvi
A1DHWMeUQaxaTxBOEyy/mMb8CFrRWmqZ/J48rl3Vnfnc0oJRVi47TSlMEV2o
S+IhGHa+Bc1xY6/VxedVm6zH5EHhpHbA6fEfF5jw0qNJrtcCmKnyPG7Kjkl1
JInVaAh96VFyP0BlhjpRyvgOVzZlYQda3zq2FRy9m53ABUKfsjyeA54fXYcf
ADhIMyidLEPILgEPKbTlIbr6mc04DeYGM/AfSc57Wg950bSdo76Lp+RWkfSw
0nCPBt5gazpx58tL+9biYQCVIQ6++vX0UjKTx+GOiAbiBUGpkYGK9Zq/z5cR
SpAnmi0FJVwK0O+JXzLF0z7xip8bjimtBU7XKuVX4NDPG4oopfHSQNseeC+0
nRFUA7y0g3DEtCC4Yyf/rLRio6Sca3A30pa520NsnTuJ6sb05CCAlJ6NQ6HQ
0PXlgh/L7jMPiuXlWjyleYBkHIONLgMcQXw2LuHPamxXTUcr13jMlP2Zl34a
397EA9wtAI648uJn1pnATO1/BSI2PWjNmE7r31DijhP/gcKL4BBt6dxbY6T9
pXc9hcThdFJQi8NzW65YVprjXp5JWjP+31lqWuve6OO1f0M1VjkLAsznxzio
BICmM4pZoaz5t4FAN+Hg8in671+SvvN01GCLn4tz49hyfIrSgohUt6V+Eqdr
qqecpZIi/mRRqIrvjVR5RW6U1MaDKfYjjJut50usdrZkayYSTrkXN9q3nTdq
nUkcPDioBAvyj/fTyJb+b52HZVT8M8LKT6YifwDI5Ze7eLsXmrStWcV3B17g
KW9s9yfte3odG/ml+JEXf5cDsIfrJ/PJcwWVO02uoAKPW6k2XxXJxHoZc8zg
iBk4xNI27ckw4lPrgkzAz6u+V9ZcchmaM8I1rhzIn9TW3ypIlCfHrbAwC1oz
cAkFE6s1FWWtnX2ZBpeJ2boj47wXu02JPYFSCytEOC8Igv+2JEs93ribK56Z
rtps+cXAsdK3Iw/7dWt3lnMFT6lz2lw/jHT618WsaYkK+vloyT4AodVOMrZ9
vzla8t4SAw1ahEVHFa+kQOpXVM7kRhWzQ3bQuWweAk/sfrs3PCLQDa5scbES
O2bVvA3/zq9G+gU8kk611qnRjNd4l82qz5POD/EtBEDuxe6JyKux/Yama/3l
a2CCz8ZdyTd1gtM8KmjKA9WfVuZOYzevPmyomu5INcMP7PVTHihQdhC1wrEg
/+WzQbbCRp5ktnocMyDY7w1C9rbP+Ytw1uAa714hjPS8NVawwL7eiqOaXRQU
P00EX6Ow5kF8Bt4/1bG811j/aULZdvCPJwDE6x0aBZj8NgxRkk1Auxc16QTC
xUnCpPJnDVNz/mQuZJqjB9wMzrCRIZ36soFd0hGV/4VcjiCI4Es+RgUYHrh1
KKBmJs45059NjBYSHq6WqqH4mt+IqBefm7BGpuQ5ZotlgaZBsyVz6oKK+T88
CE4KLPoziXyQlxdP8Xi7kp+3pgifA1JoTAjgTJFlXs4YHTvK5R4KUI5ir1Uq
oDDeahB6TnVYw0ulyetaa6znmX7mifFIRyAwQsHFmVk6aOWA7AOMizi4xWE+
Ap2gEntBTayZF2IPtUIA9c8Y8UC3eeGjUYHkWhU+M5oj4l1h2WyZcCWwWNlT
H30wo5omTJbfhWy86ra3KjQqLVCHfR5g03cL1YeGTNbkr5vpXHITrZKulwlk
AXBCVU9gf5k3DV+ZkAfrzYl9NSs9IQBxwv5Rpff9JxapmU0d1X0xdnRN9h1V
vPQPzC//ziCVDFIxo0ZN9V/Bgp+t30JPlU0Og5Xsbogcr1ySN/gAQbT9Axxi
waKuBYNvZhCzeHowwSDDIchQtOhNZTpekApxy37L0fUdZvPwtZZeZyJtRHch
87VPxF0pcjXXnRrG6YwPHvDzHzOBp5aRDvWgFsLrkKpCbiwnspfTc5lJUuMj
SYP/snudkqKCzePM4GVuQBNblxTQdLji8O23fTeKCCS+kEbhBo0PJhRD3CrY
Es2UJGhOEs3pR09R8U4/AsTzug+FFAsgpr3reJnc3VmVC8pJg8KWc/JztIDU
KBEqXWqVIUUrvOxgtSFZVpjzHzCrBP4YqKeoCilMN9/OKl4tntNpqavtrYew
c+S/M0SAhbd5ljg/P+vpVrOduXpCCRVzx4CHhZx3X1vMW8uCuRuSLm/WlirV
v8C41ZCPpXxHAiznFeK0jCi+vjDPRNY8xFoHzmYNSuaSn7IRTk8Lja2o2Fpp
n8N1Cwa1Xdh44QH8RXYqwQs4vwbsmmNuiVK9VrVHbgA5VaO5si2mOUYJmFt0
usBoYP34nX+pJ+32b5EFkemT7ZRLOYwbRked5gIrqngaZqzVHaX5G4kyEpJ6
u3rtbdN7ljlrthXZUbEMCA0QCm2pYxuHb9HkpzSgSHJG6tlGsnq2W4E8ch8U
1ZK7i/5MCezMfoEa/pko6Xjk5jw9X0g2fJ08ErvZss4iuZeEgGwZJ0mrSODx
wpOuwLrCIlxQlZBo4qL/+Cj0YHdlFFmzW9NPgjAOEFdoq75Fv3VQt/5dHwmY
bL7GoqfDQX4CVGrC4EsQZblKLCtlo+sRFKbI2kYXyiROy2kV7dSGIjAELx3O
JyXoHN4v6PdegksKRH/BMY3jW1bnkESUQr2pujE+fwLWuI9i6i+vQQGtUIqq
xyAAuYcpBAchyWeCWrU9Fwr45n6Li9vRMt/I53FL/iNzwRq7oHBp3Q8Yn6UN
ZOQbwJeeopKgBEKWAe4yWpr9w8ZHKvH6CPkPhtGt29b/8giW0QIviYnW1jZO
w59eDZxt+vfT7z3A6pfPu+4ooIKSWRplY1baQT0Z2XFiPNUElF2STopdRV/d
jwU/JuQPSqxtOTX/y4HRYDk7hlYJB/DtgvhWSPXLvQf2Cf9Wdh3lRxb7Jfas
kKWPER78XwLc08IINZLipb6xnXwdgdGODpmWsz3EFX0W+DYmkhMRUryOHFTg
0wq/+cSoLVaudab4+ryUTZvZNerEbeozE9ogRzqqS84t4aYWK75/po43rkan
SVmlYIj5zdT/4fmtEeWJu8l2olJ56+rkQuMqklOmurUq3eN+ZfpT5DiE6y85
vuPEbvxGRfSaXdCYf6TINfSltSm5ik+YyvyPT2Ni2O6eTiIVcrSdaf9BpNqf
e0TJ/XPYj1lsvi7LiXflT16O9a46fV6x0kNaAW8ceTK+wybX/V5sEtiMQat9
j6+BDdFY6LOh4fbHfNlv5H9Nt3lXxHKyR4k7pTVr25Lu2vdaEk6l6VqmzUUc
l5RdudNX5FhSLQUZosJmTdbCzZSRvdP+pkSFrXjMb0CvR77gUdxrUXAooDnt
S+zc8ro3xBSs8T55avXHtf2hF+6aBJwBAnsqNtbuiKlVlnIVzMgzJjJLngCE
rgeEKRGWsa1ozJQ1W0doZ6/Y4Vhloi5bMXUx8ZGUzA5ncTI3zSy0K8GDEbTo
IEVFpp4if76PY5a968lwlKRQ9WdRXtmC/1d6TWpoyzRduTqhypNbHGOy2bnW
W19/uK0B3iwmAHJ9e6yXIbE0z60Jf+5ssjC8YBg04YIZRRG3MJANkmsowjuJ
GvTp36R98GNIKfM7tCEN6CdFPkpoiNxqJQhtNyqNPSUkBrrnPYeJnV2iG0rF
lmA0CsXK1/RAC8Wg6pOTAyqbQro5btmPraV+csMNoPvtlyDNNEULfFL/4kPg
QnbqErVqawP3ss9ElvSauHn2NF94lCSHKk0/SeEO7S3yh/7g0qAqy3BnvuGW
gMsw9jO5bbZJD9WTHm78JmZlm0hG4DFVrmfC1zOz38q83//xNHXAJpIGIyYa
XMKW49yTL64ZkMwqNo3inv1qwNYQJL8lYgy/S+3be0z5x8VsuppDMpUsPv8e
fEsT+Hlt/DbWJOs9PxAiNVfl9eaKadP8ZsqDMfAVCOTG0vI7f2/zmis/cvCg
oei5rJok5G4eLw5pM/dukt8q+Y1aBq0IZGbhIfp9UFULLzWM43EjRs1AnW4q
pI/qHqxgsZYE5AJLFDo8nDpy8ZFIAkhpSfEPK0n+unP0Agxh/Uzv5UlMLOYV
esBE9RdH7613IK2rzaeEDUx0vvlq3RQcSTIdtfy3bAxudqBOhaWU4hvcuTNW
GmoKeQjWvspQMyZsw4MgJwIixmOxKLFdit5yv+RFjrxBsRdev8Ei+jS5GNxO
O3fB95UFdbpjv3ixRSGVlDrqkJJRxPtxXbMVEtB8BlLn4Vv8NpSCw3hHxiCh
1p9PeubUSC8vjfhK4U3f4uh69xZcfnQ7/vSdeOrDjrLhkWDkKK3YcsNJ5Dve
4IembM2zQBa/urll/YdZrEmRs7Y3Ka6eNzyEbeEXCuRZerHhcM15THSzoVls
2UaO1Kc1wud8jeP2jEWs9muxP/eHj7QPW5k854SidDXG2RiRoMBrBYO2v1qi
ofreYtsLr2qJs2Da0V0BHurX46EvscuJ7df1E/KjhVniUKvmI159hBHkQ3IS
Yv3L0x38Bw59EKYnLyzj0Hn7MVtPPARUnQRjLxOBsfHllVUK6t48IM4V7a79
yPkyidC2RNKx0GmRpzFDgyhbUGYseBCcGEp52VRB9cq8dtqaE1516jhyrs8U
gJDh+emO61kpoSz4dkklq0koRXPuH8N7Mby5CeInINykVyCBRmkY7K4xDsDL
i68ZRkppOmMCaSvLf+iztotScbTGobw5GvIRB7sAGyT3JVOdFt9ypLyc3KI3
jTDkaAe2H43r+z68uhr0anUgU6ZPt6SCP/dGt4wLqMPdEuJDnJ1sS3h7WXrn
iXj3/64iUCY+UUF6KQ6COHmEzq82x+zpOaO2sSpnyLjAaZAnCWIbap4l9m8L
0jlOUa7mMCj1yolzOU+EXD5oGGCHIYlMPRmYUUenofzOEHyVhZskbDSrOPM2
wh3QBpSoE8bUk6yPvyGguGPkw+iYXdbEH8n/f8HtO6zAPlNnSjkxQBubQs41
jkG/diU/edyBpaJDQovG7yD9OSG9GSBDk72CDtZnx7MXXpGw9WojhV/9Zvqv
XNjK2VFtQmCdwZW1vhnzLgyQhMLF2WJQk4CN4lJe3D1Jr3Zj5IeyAqaJxsyt
fkhEurGmcWtVOqR9qPyyRwfiPfRtDAhry66eS8z2qVj3XVNNuF4bnO0q3BeS
aTfE4+rlc21g+W2rPutyrGSbS1A/08b87QssG5ASWaDhBJdBGYXinjm1ZCmc
NqO6j3U4eOV+H9fP8pM9xfOxB4ggVVFYhWgktZuVyL1IiKcQNGOCv09BKkcu
ZuXaSuHC0KcVfvBjuxs2Osy5CeLdkpUqM42EanotGrcsTJwgkZldFcbK3w66
IlWLVyhb4l86G97GAcDB83z9JC2HR0YS68LIimgn5MNQ50GHQ20n+NoRD3UL
YPmeRRK676NC7aFnWrp1ybXnEPJiRDrxF83sHs4fGD8V+srZ1X2LewTDcQNt
3ktwtoKZp4r0vm0uYZrrVaHfkvzjj6BgRur+KT011j+Gxo5eqISOBrOVWxgW
Ws/+OyLfSXQwYLhZKasMyewEKJ0yKsWhKDIxreKPQkuy+H/xA3AQWi8BrxIi
EqNHxVHj+4rn3VxA4ph4pOJ0ISWDViolMaJly+Dr5vPUkd4kHIamp2a6xtZP
3nsmvMy9WX7EYMaRLIwlQr8oeu9Pwzt3RRK1gI9y8Mh68u5X7Y2HqkAggaGN
v5I/T6ETBJKfCL4OyAmFMj/aLpX9nGeXteHmcyDrx3vL9MsWHeeSpUOIp2HH
nnwnjhHrMWXKQNjvTtNXAtaAX0MSvJ8XIkHvoif0Y/gRShIgwCuOyn8xqrfg
ofQVtiWw3Y6IyfytUcQEGPcLVnJ+kNH+MevtdmMrjKd2z4DxY6ztRRBWvqfL
SgUX/qxZLZpvIj3e9krUq+JZgUh467nUNXGtpySQOeg0LfIxb+llg87xScxj
Ex2ZiobD1bH1pJC7dcA1XhaPhDBJH6wP1eWu+WjA1/qO7y+MfWVONPwOsWec
QNP883f8Jrr6DEUSpdBvV+ycQd8O2396TJUFDYZKAWSoiQ0pjjKG/b9UnR/9
lDwiSYwH+I6OajoxDAZDrTIL29b1awKxssyTsGYC345CL+/pwKZ4WlRMkUKq
VfCEUm3QkkFH1Ho2z+R6eRSML4J+dtzlUnqmnFjtTiOLdF2cy6zRb3sS5imK
+PlP+w51Ifq71zjy66IouYid/N65dI+y7w+l11USnbPMdJWvCxJeys42W/WT
ymkTNStc12u/BoR89nED9cvDsnzp5Vg/psUqkJJYno6lSLtruJs54P6tBzQ7
IrdOX37roFtbqLu3na/0aC3IIjKKONjglg2658BIf1XX5lxSty68iwk+KFD5
V19obHZMUHIy2Hf+86Bqsws1kWLv4peaoARU9fk9sJajVaQ7ecatJuY1GGmD
Jb8K69YwLuwhxJY4izT9UT/biZm0rZhIvynNX0YCe/53WaOY8I/2jV2+TDt2
rOBW+ac73wuWJCCnP61g8dOzy9F4+QyIRflRNlxGXkZ6G/wyGEeDzH9dxZCK
kkfNcaw5nVpzGfmYojjgfUTPbkzNIzJfdn52oJ9/RZtU7HjgR/8Ehk6lmrjf
qkXxS53E9wsdENXdFtJ/WLCdZtFiKdIMg57tF4Q8y5tKfyBNSHUGLaevb5i2
BN4ZzaZWQXMZZ3/9fEQvbAgibCeZMSFph6iEnqIEg+EP2I5QRkKTfjJKh6vW
aqJiXDLEabOUCxz5q1SauiRZabx56hXuKjRA7Kci4IyJuSrkj3PUUIbsSFz+
8Y8k09aGQJkLXmBBonJGJ2lGj0I4xiqUo3SwxOO/e5+2JIkDNy+Vvv1vfm9c
+jg/tSBek+K6HNeEb+cSwEtB6vjaoXcSUaKXmL7woY0eeNPn/Xd4012Wi1QH
09RfHGpzsyp3R5E1WbWZjpL09mKaxwdXVYLoDsTa3QCBXkC+MuhS37QVBlTH
80hZvUQMEH+cW7+h2svREkC9ARpyLm/sUjFd4DLwD48Kx/pu5jt0ALviPDS1
gUcne+XSDwmRNFXBuHsUyTvtE/owsln9XF5Athovu+BeYpLEoOLDzEyocGDb
KecOPleuCB11VQl23Ex6GzTZOfP32/voIoafL8gm3y2rmU/gh56sn3GzwaRX
GvS1lUcncFDEnddMC7INMoSvsH971WYOJMPDjG7Tp0Q+0o7kYhewQ9yo5zXp
AEJ9NfA1shoV0oDcSsVufc4hmEdQ0iCznaomaOlPJL3BeSkGWBLYO5yT2MRL
/R4nnuarb7KPj5/5KKnmqzGXOrDE40ZFewurN3Y5mxXswoc8LrDq16FEHyTQ
qaTTXZpIoqOYuXfdwhiH4OtKKW2amp8+dXcxZWIz23Ld3FcfRnBpl1GVzhiP
cWU3fbC3uB+DaiHv3JE+NLxTr/cMxhvLbPO+cXJC1zHABuXbLG5EquzpwtFA
wsi/v7LD0KR4BzxlwM4xlItXlqLjLWYtUh1KT4KEWrDU7aSwX/X0ZXWU4oEc
u0TfmQM2IXHhvkUlPfD5z2QnNBrLuzMcJg70YJf4YpaG2K2/UnjQWF+VOmUs
fPV6cCcq8g+wlbmu1zfJ48pwXZg+SdZlxnQ6GFtgCOpDXT2IjrvSr1pboOk0
NnijAksBw1YlpwJUb8/U+dRks8omhKXtvV0nlfdO9gyTwNjeAkggCkdzhWfO
f8ebfCHNxeLlDiONPVC+OKFFu9VwPaIKdTD1QWfxGzy+riyIa3RID4mllSiX
jsJ/lbTXnzZWbXvGKqFIcH0ppcQHLGBgu6+WBLxs6ARw34oTIs3Vu/XA/0Na
p15raXzBrQh445zZxMNOR5YXPDhkMhZ+qtuzAn1XC6Wz/VkbHPRGpu1DaDNv
SKgQRZ3lrBWADfvY/30A8EisxlAjQjNCya+yUVCf0mVq2fiE0ngdcMheklo5
bcMzYb7zxU90KFC5VZLiknTdKBZcoKmclBftrCU/JuCioNrWEb4Hm99SgrRd
ZtkmXegulPd8csDbznx1lGVFkrUdRrAG64wuagThrGNFSKEMUEmbU5/cBlpA
tEQ0u8zQQcmEBY+XnLkQwQVvZNlRRD3twNYGzehwWOKZO5nuBpsk2XZ4CsDw
b+xCQVwwffqs4gVRgCE9ifTNa+lFKVsoUK5am1M2QM1aN+M29xaIHaMgRZJ2
UKaDCjdflxqYD9TySvvHyBh3zAcosh2bjCuh2mo22GUdekTvl0HJVG/Ia1G/
zXaagg0dFurqEsx8uasP8k9eT4j9woo5KRz8xiU+TSR6r8uyREb3Ekg42ScH
0jg+jPJwC1vDjok+ker8Sf5OOEZ0u0veV3iOeORMO+vUCSnjGflDsfwKr2lg
lRREVcbuyThQrPPk7OHYVQqhUBh+do5U/i8Rpfy4YxwGbi2kM4m67SeIcO58
RoUt2kkzxKFcfh7CYyH2mvl4S1XYFcSzkT4j65j+1NxyHZfSMjLvcwVea6A7
gIes9g8miQWOWj5XRdm1pkPbqhADfT98ogVw2DYNejkq+fLjivc9xEHvA52X
Zaz0cp8uXptnXXB/j0EBaz6jxF2k/XQiMjzxdzouawJdil3msfFdFc64fNd3
mOy/t/xTu+HH1BQRfa5AfM1HLVOSWLTvqNZXQ+/OvpDUxX9Hw/NMthxDweFx
4L+TQTWthv8bpZg04KNdoN1JR/jJBNe6ugCt8Vqv5KcefSVTVaz77MwNM5Vk
eE5AGqiMdWSyrn6foEZEUBvmaDdU7q/hXdZDHwr25bGhvaWsCxd+p8Q0SPo+
swlByvilfUnO9djEPzREkIqgfa5JCj1lipIQuj1ans8XYX+gmOHvuEtv8mz2
imHkwbucG+8WyQ8tGO1d3qxkbg0qzFb+uQb6dwvfJbQlMAT8Db+0F2kEIhpE
ExaofFlzoMY94wKPjiku6LmVXQB71LvSN+1TU4HOfmXEtL70CLlXx7AatN15
iRSqegCcRUXpS/SEYMpX7FOZHjBIRfDa64z9uguqPjTC7a5E9O7paN+YNwu3
x1kGH3nt6TzI/Pwexw434wR1+0MHX1s4dCZdgeQRm8RWIguIe4tUVohJ6XOb
cFt8J+LoO3t++nx9e/xD5V/0BdSIZOsuk1nyAypM7shPO3V5U36BA6Tdc57B
HYEeYBSyiFC7lbEbB+oTh+MzALIdsYTjRm75TIrtQwdskLQS284ymBB/YrUy
AjQheFuNVdZtMyQB6Y/vcJF7NR3IqK0Od5135gSGt8hY9n0e5vI0lUfpWcYz
7+PoCnX60EFQRBEFIgLx5o4+kWUn8B34ub8XZdxRDC7YUMisJTxwH8ZSSTsj
4Fy25bKJJHUwrhATEstDmSC079k3aMSe0/RgrZL9Yh58Z2iKihM48GBhV8u0
KfQUViN6SyaVgOzg4/h0jsyu6tkgMbFibJO+DnVJXQbBvNCIHXhqzJP6/Kmh
xnodkNLvioBfT916T+AGB2eWEgPjQdbALAMsR02nFTjMjQtjz49ichnYu5hH
5rg+b/AKK8JjCQqrlb1PPprfc/6DAOjjM1LmjkB4w5TNrMJSaYA61UsIAAjA
OdMNhjMvXId1gCNkW45djg8286eM/CL2FxTAz664Bhk2xDXwSvrEnyxt/d1h
qnUVFoOpC8p7wC1YuML2+iTYdNEwtqnCG2q7gjyLv+OH0QCFoO/idKMA0nuF
2M35FaaEvKt0pxr2foP+njgewA9+Ikzc1zuKli+FdDUaA+yHONn8KKTMoh3c
nT0E/xdoh6mgMypngAVqSY219DD/JAgH+18UeEfqgL71kz7IvsQVPLanv8tq
17/prAucFha3ZGDMFVR+rV7iZ0h9mlPz3zarNCTLD35GTJ+ijEzgu4uIFUGX
XpV2+3MZRwjByFrRk9XR4sJN7KZUtwCb2j9fJQ3ZarRryWVOiDOMTRslC3Dw
mRDcSSWRznham6UAEVrU4H3Z9rOEj4pSbeNw8yMUV9hE5OXiwqN4CLjBXVM7
gBCGNcad0J6mSuS7hycpxwZZSj+IldV50gVcj4+GQJ8h0sI1+i79HGAC1nx2
2BCHfIOAHtIuLElGhdA05ED/oRWJhZDfaWyi9WJV8OSS2EuEoTa6N6EAK8HO
/DtnTMn1miq3GejexhvIW6bj2Rjh62uHN0IGufvjjkUPRzxeW7BOvkfGsyt6
R3s9iDmq9BlOexTRheaOCpOmHMxj+PzjNrsVZ6Q19eHwF7oct8cajDTN43gF
CPzuk8fge7a65BS491TgB23XNxGKVCB9cnuldM2Tfhsq4Wblg8sxMr/OhCdO
GEZLY57WeZSB/E9EICJnIgMUlUUqPenl0dqbYsZhWA11HEsK8/XmfsaBTqz6
hAbNIr3SqEzcxe4il3e5NUhUBrBo3auzCenvemv2EhAk++2uNKVihoMu5xkB
5HoGBeczMDSM3kpkOMQIzQfljsaC+4gaN1j0dKaRNsq8pMeA4Fx0M8S1Tctj
cJB8UQK3f8Yyn87a247Gt3dEOUpy8bcfM7G8RLzAC91mmP1qiDzR6LKbkWkW
5yvzOL2CZ3nmjKpyKqH5VYNPHZYzkOCkLaUc4W85YHJ/IhxgdLB7ChmtAdIi
btScmDE9UndVvncGgIQZ8urNsU9B9SQxQwS3DkY6mbhomsTbsKlrGRhyMKfj
3I/yjczxbvxQS+/k2zn0REf0C0EHBEK/F6G/DWjzLh+SAovkpMiw5oHDvEUy
f59RuawwmTX2zlLQQDrplCMZCbiGF6UCF2IBdhMhJRS6IZCewYojbyBOGwS6
q0NQVY2cltHJQwNwXaJUnWWHVT9kdXQvJjYTkmefPWHBiSgI+29VC8/1JPtc
bXg05jJr4o7ppnG2flfslwbzT/AV4TIGtVVYorBJ8SRjS+FRNbVHDLxQ2z6X
AY6JkpZ3OUA4yFxSgnocMr1jgFzHY05LotIL1R31mT53ya15yZ2CjNtddUGD
TNLYW4M3Y3AVND3oi2NvrFVqVyV4AbsqNw8+cBqyUEBGFZAjlBnprn4QC+3I
UDcP9oMwVo/7J95YlR1mlugISqL0W02hv5cPONzO4dJ9Kshu8GlK2NOQPlX8
LHb6BE4i8hocQlui/ay/e5iUCudKtpyj4WIyy/Jp9XC2XQQtxa/3N+/GgJfb
sG5D7dn78JrMHpOMnQo9ltGxndqwIezWztE9YemXcZWzPdy/E/FdNmZxddHe
/eUWjwM2saq+T3V3m0jBjgGWWaZxqOWMGYOiUr5szKazIP+kCJYpyINJt628
sgntx0sSfkLbSKXpc6u7zpyJ4XSmeOQUfhVG0lD6DQbcqNFgCNyLCTpRDz0f
wXQbYsLfqO0+S8gWXOceS2B2TRlNA0qtDtXMaeHKSKcFhOU9A2erSLWwG8Bk
dA1MP8k0zh0q0BQsnhICOx8gBJupt9a2F9UBH6Ecdg7qMrdaCsnRvfCoSWQO
kZOWQJEaG9gssVkZ3thLQMDYqAddRyBLUusF4tM/LwO39JLmQct+1nHbVzs4
uZYrIktp0oXiRBJm5IWbqHVq/Q2WpaWGxg3tEi/RPFuVN9JyKi48RLlFwzkE
7grT57UxUu9pZCNfROMWLlWZmIMOtwf4p7o058sPlALTbviZ2AJvb/AbbsJs
WAYREJ0X2Odq0WDFdGChtmL/drr3lTVF9WjDXgKC0JU4Ox3J6YpakXVcJkRc
d5YkGs+dORrQdwA0Am0sAeDKGmpAa2x2SovnznKsOKQa90vCooLuqwBuQNLq
/vTQXZrvfD2c9t5JIgt7I5LQx+0wxTrUQjPLBYZ6fwD5oAiYAOP/4gMzrXJr
CzUAeScrdVCq06xnzJ60dAp09nsejA/b4el5329gUKnMy5WzDeeoNp/hCo7H
hPYLAsvRVxTXZhlT4XJKspCDKPTf+WT+qkIoMIwjsWOwQJlpPRKbMdPiqQEC
UyPNU8y3zN0Xp5UeS7ThL1uX5C/1i8Wfn/t8/TBr8z5xxNO0ZoUPLTqkWZf9
RO20rfVC1YA0d3JInYu6vO3bYqSysvAD5P1fLn1URDSWVqIX8phlCD+r/Alb
wpLZ4nDoAqrmTRiG2FjXY01Etn2uZ/UYb2ZcEBYvdlLLBkEdN1467gvcEjIz
ht7IeKQ159UbiPM2V8pGqP1HBRfex8O+ysWdpV8PjJMrH02+8ghiRqNoUP7n
RjEM0nSl86D68JHNrZnQMaOGJYW6E9bfB160S36zNA03mczc2ye3zHCK610A
Lf11PrVT0YdjbnEhRGVskujL3juBU887Op+8fSOCgtg1zn1+GeyOFOzXH/rF
1Z1ZZDwNDQOVlr6cwVDz+ZeMmQOrIGjlb2Y1pRenPH/5ZSDT+19a+3yh1PbC
RyK49F9zeT3d0WtTCw95bguIzbek5rMcj4PvlSO4JSWGlHhZtaYGGk/PufpB
gcEcXqkcO6PfvLVbbul+qkubXOrmlkmT/vomhQO4cmYoeCkD3PrFuczfB9Ti
pUB4F0H3iGT2GIMzpGXk3kPDQ0mGdXCLCkF+lBXa0lkOxL16eEhUGT6gZfro
mtZ2XW/sYnjM87m0dMGd0UfCi6aDmTA/sC/qHHMFDMzQnVKbuCJa5Uty1ySH
gW/2uekf4RzRffzqQNnaleq2H1cTl8DPaNOx1I+B6Q0rZeA6b8TX4j3s2bxB
zAZdGJQFkzG2+NPyTp2KSiUjkXz/lWCKLr8VJaM279zSWZ9VwXONRaEdEis/
HELLsN9rm/UwhrfuqxZO2qcfBIF1rCJ/KbmUreVVXYQaeixKujCmqsFPHOYT
/rUS4OR6mO+2+7ik7pyh6Ti27A+7pTfqDm0ga7mQwwW4RKvnHV0i8Fl5q2X2
7fNzppdYlJm1s0XL2UnZUj94HfIMFOAViORNuZlgut0IMTpLHrGKXo/7MzJA
ckU4BtbjAOdC0kVHCkhgOBQ6jV5SIJG+PN8qhE72PvoJ+fIcL0YGEP1k47mv
ODJYWUk3wWwDINhevP38bstOAdoFTulqFd7T8z5SuiRfq9St0mv9lhLyogT0
9jMAKelqNeYh9mQJ29N81JOrx8yfqdTWwOtBlZ6n3eDfJfolRYOrp8jVhzat
nHNyPJgQlV8HmV/cz2zBlTvFAWtn5ouViw0lL80smieSO1ZxafIcYCAfJMyl
oBJ3qqRClXwL6OsYjrVAeqbjD9INGDKSlCl6Y51e16RRoFij5JlizLFcgpv/
Q1VXDKVfVPcO1c8nvnB/ATdtjXZF7W01B2DPhqq74yM77+K+UlofU87Valrt
rSRrWwRNFU/Q4V5O8sKok5V7lWTslZ/OZJnGdGfeh0RYbcOAwzc+z0jGmRNr
FjrX5QfaljrvxjT1CjI8PwQoYJSVy5tXnancLNCcDelSUjC9KF997kWHaSZt
EZvwuNPjdamwJCNN9v51SlZhuMlvSMT/0a2fCbv9Kr2PFoH/mmlRSZLA826m
zmxoSBqoYMzGQjfF/LTYnCfvThOmoDs7qGirtWVAF2Ab9qLuUSimVBuhSUkx
gxv5xo4UHdh2c78HCjYHW5AxrcReLE/h+dTncdMMdtSt0BPR9jLjgg70A6FV
7x4H3pAlcqRNxjJnMFU5iTLwk/A0w1kP8pwTa0xe0KvUGEKrmtNpGKFUPkAn
eIqAnW8lD232U0cdp5gaqnaIou/cKdiruectj4j/v3kTKTxSnhSrsof2KnX/
AJAyUWmqtO1RkBWQEk+Fl7h9RYaQmshHtUzp3DOCydLJN+IKTlptIYUB+nDf
vAs6ds5dU/6ZLHGBViDn6InLfAemlRRLG6Xb04sQcKwhGjvfu06Y1Cb5JdsZ
VQx9O1E/r6xJCCbyAJJ5EpZj6FpoMA8ATGozkAH9BsPrHg2cbxY9e2hexZIP
RFWPFlc8c6jY1pIoQI0w10hDxyfWmyzDIx5qJiGQp20VgJgV4S3vIZSWJofU
itRo4YGG2hGM5Yw59sCGWkEkAeAvTL3+FzQZPNKNGN83zR1TerWHDDbyML/m
4y/Vg4p08gvzpO5S+jAZWzEO/lBG1zoqvuQGQYiMDLxAHTgGGAS+eMgjIVvO
AmT3/IYAymsxFj3pqSJ99sbw5TiTlu8ac06pGkXfr8MUXA/JexELmcmrAwHn
uTedlUkzT30a3q/W+edx9nwCHZC/8J3KF/2q8y0o0EtXgLUVN/OmZttBio8L
yDjBM0pR2yWdRVlXdMFkT9isWfKwmhVOcBmNgneXBob582sFVt7xT1kGfgml
pgnWXpAOltoQ7h9vOUp2Qbpkj1Z3OyR/Zii+qW/rRjBB9rgXtkac22suyBoa
ClEJBR+SankdTdwM6WyrUrNHDTrxC0U1rADFkfO+xXWpPGPy7JiVzxaEs/c9
xdtgKJBj5TyvBZiXqII3itHWrw9ZY5Ep8bPmRx3pt767iz/b3Jybmtj6436x
4wsJ7Q/oPrGXdJkcKFQceuDIinEaNP4HlGpW20utslvUUCO7j+DAJAd3KcgG
3m3DM0XOvhNUHa+M+NJZny74aFANnc7evlTMZVhw1zM0oTIy9B7exQwetBIp
xek3VeXJXOr5tFTW6/FOJmS5DiPwXVN0fzgihUWRk/CK8E27+sX88VdNZ1ye
oiZXxOvCIUIYaI6gJDl5FJFbn4fwiiF2rFmxM5yCOIaFQsFTS9v0V4GfNrcJ
73q5TX5EKf9ovzbcBlYyao2muG/d6edzgpsQVj96Z4i8JIWO1hfpKqqEYbAF
tQm4g4iJm7j0Bd5ERLBY2BwiSdXRU0OY+VIPkahH8fL2nKU1KgwYIPHKJDhD
D7AhYFE+HJjamP+O45Rd4L1R8YSb6tD+zB5OsxRf3iovbkZKICO8k84+zVrX
Q19INZjRu0JaKwi3AFx+TsrkDlZQIYHdAwUM9cn9WBH8hBosXTAyfDBFptu8
SBXZuidceaXgocGSK8N0eDMkaiAtBDDJl0xYFcHECohI0meMnjNvMqtnlqxI
sXRHoqVQO7QUmdjmPaucti87mL8UdhTlzvsv6r3fEeFI16GV7c6qVrXz2QXX
qr+n7b9tAhoHgIuVJ7TdstE4nETqAbtIyb1MN1VEduPNkaPASWUWT6EfflAe
Ps7BsusBERpdyldMbIK7WKJ+HEycEkBR+FDxCrIjfYgqTY6BepzoL6A6UjYX
NRPsQhJsJ2Up5pmaxFZ+CHF9idw2a8HBzcO/cZKx39BjPPGtAcSrqLbB3Slj
2tgyn13Hsm7cm53JDHavpUzREUiN0cDhkpc6G4VjVG24vUvLkHfS5zbxRO9j
3dvjvbQXYnMBe3UQKRJcsOxx/hIeaXqIKacyr4pnt3BjFrH6ntBDL7oXnFl6
UYHPHTL7OeaSklBWb0A5qCFVMJZA21D6a4gBKV5rxCVdeV0/OG8G0O/HOto0
od4wSvoV9RSZBoeZGgb53dWeqlsnFdAcnaMENfAWokf2JPkLmoLjR+Be0M0M
KwD15c6be2IKhqtQXaiXfUHS3a3F06O4Vm26SbYCOKXwuAiHboDuiO1AaH4c
zvXxQamSSjogDHojP248ZaMWn8KxRA5AWGiD2Gv0gNch81ga42OcQ/Sk2GGD
6+sQbIoHX4VlOGJCfs+PBp9M2ZRQOWDc02VB+WgPXavnA4ql3LL23+S1Xmdn
B0W5truJGxM4XW8lLIe7GJIoMPCqiUN/KdX4q+an3t/I/DRswNdN2JmB6Ml0
ttZYrX0LGdipPd6ax1aNcJqmq/3PUD0T1ypWc9EhzmfFLnRqMH+XQKRRSm+I
bYFP5EO/3wI3jN33r1d0hXEuKvEEBreSbJxl1ofAtkctUQT0NIhCIc1sogqz
KJu33AGUB5Qff9nD0w+hNEfHgXChVtNX5y1rhGuwofgVYo7FzMuNRUGSe/Us
2sFAPzKlUoJRgIVhwe5AkNXn19lV0kqZtyl8akGOEpDnK6bD+Z/TEssMRYwc
qzSjgpb+kUv9nU4HS3D5rcRg/XeGtAuIlzmSKRR6QNDrim6oQEXkmigtGqIj
Kta1WnaJm45Qv4kpuFEzYqU3CDEvKQnS6DV8BZlnfyR236ymjAllOMNZ6AV9
asuiFMOuClB0VAAN/OIeHHQCg72/qXVu06zZphT7D9Iurusq7Z6vgWEMKovH
N6IgjoEDs8sEcKdSHoJPxWUIUvnUrTYN3SIhKuG8L6nF1tomPrZ9pviH7Cq8
caJ6w1Qk1cCcPEKiwg4sREb4UYrE/8mVVcGWR4Gd0QcguiOMY2s9Zb29C+vY
ZgGV740XAUxwqrFihXL0E6oYkLvYihpqV2YFQyL7UYZTziohUcKhuOi4uuLP
pjtlt61u6qt6NfOzyL6o3GgLYnX5H3jBNIK3vlN4hMKzQwamNjpZ7oAAt9ij
NUWkkc4GMMkFdh0fvHTBQUfFeq2IjKTsh9QoYoFflBijc5642AHHV48ZGyvV
O04NCQl1xz/qfpxbDI1Z76K9YSGRwoYUPe5XSfzbsxZG5uQvstarHEXUPP6G
06hBAIxvySDInV6VaSqwjrJX2w4BDcIjIFkTQU0v6Z2kV0cGMrJmvPTKOy7G
KSwGKyfoaI7uYL4bbfD6WnVPgnN9z5dzGnvw27ngWq93OhHaFv6i9pGvOZ2Z
XX3btdua7hBxlUOI+YqOCnHCW2YFxHQbfOc3DjXuIGzO6FI1VucFmBLnwZ1l
q4+JZq54rFc6clB7i0OwffJZJRxyM2+u73DZbYSZJgapdxKpVHFU6MtXMigH
7kdqXca0H+iz46ycQmxLTfwAEeij64IL96CcfEJ4Vi5lmbuAbGYHHFYduSw/
Ch8UGb2YeoCpNUWIrTEdX+m/DtcoXKiUDKLgLYlXjN5RR2KoBv5sNl9pj3J7
oXY7e3DT8y9BHTgbdnabcDNfqp9eDyC8Mf1dWw78d9FpLs7WGhmZ8t+mbEpl
zsZ1WMWfUooOJgaOPPzb8LFdb0cCe98vIC+Owh8RpE9euJwVVueOYhoBXx5G
GvUTR3IxWdBNKN3Qz859qVeR4fDCv09xVcvTfOwpJXI/ZocYrtT5QTjqijGz
xoabTW9pjm65hNHXO7ffqmu5W2/q6zZBptDoK6oQ3oWDl74Sq6OLHC71BfMs
z6Y8Vw9IY6DDyuXgLOgG8QEbAHF27nVijS4WDbcuprUgRJYF/XwUdf5J0U/m
tjAoDFYhNCljyci/MTQrhsq0H+5FBNaFeUafv4twbSDKnU8i78GMpOIykG5i
ci0Yo2YfIlHyMZ1pHUH7YYGJ/H8DV38oR7MjDn2NVxQaDfhJN0ahxwI1aXwW
8YwQCu+DDqH9KlwwHGwFNb3MqHZYZwP/2SKIMkZOApFaUcM3eoq/M6/zJAUG
t69my6sCaYrAGfU+VfGmgjlUE9OwtmLwfWYdL5pXchvtLCMF2IbTnTC67Vbj
RTSQ/PnDrixpHq9pb3VExhXdPHLckq/BC+DMXG717CVgo+A1kALCYL3F2FJd
SHDicq/b8gum1bhawgE46a1YRD0TCpoKBL8TXcpkPwquqj6D/gwA9bGCVpE5
oO5UeZkhlcHouCYTYHK1SgjEMSitrhee/rkZLeLkkhwksAlZvpMVdRSjBuOw
EIqUo83WrtFKDg12XaL/B0KfvSBU6U/X8XMaH1XwMQnZImbkwvhldqASM29h
DKsKj+tke9RCBWA9EcYBWcOzVSzJO5zVMIKslUby+QSF/na6pTcL1avlWHPo
GIHokcQcoTuiPPzw2ipg83HbPhpruJPDowpDJP6t6WCY3LgEHz+hd1UFyQ1t
J3+aLtwSugcSG7SNA3cYUIVBGr4RFALksbtN8nRk+MAoyn219iIUZ7YvsyVz
vGdT8D6juJafpo1E8+bE1NggiMALl0EIb3L4ZyA74qOQVf5yZn6zVJCR0AjP
BL1z0h0cpxx4MYVwtDpO9jI4DlycbE3L7qGJTqaGh3YL8cYYgaBTynpVQLPT
YHygDD5/BDaj9zvad+/0m5saElOs2zqzz8kT1MQ2oEs6d4gMqpwJW/PiVECl
6gx98zcn062UuRznxaLj/CUHzeOArUpo4hjZNGVX0ViADTwmTit+74AdmV8a
bEgWFBHEcq1Da0SDwNJkGhSN+2T0nnPRZvxsQxMQYuiOI3lJpHY1YzsP8dTz
TaZZM8BbdFUc8GKSOpeIB/y/WW1ptJbhnMiY6U87P8BcktbI9SKrSbKZMMGl
IcTsSf39tylPNhl48KocLr553lvofDXKc15TtDbjoT3M3nGH+d/6Zw19r2Wl
HzZolEAjPU9zAFnSuHoFMi9sRedVYndfgj4rk7fUdtUvC+Rw9kOlW5yGo/f6
rS6970pjT0R/WA5tSAM3Gn29oyx2DM9VTo7T55/JLLXlkt+lwvgYOYwmFW/9
H/YyCKWldywfqIUE6VwDX81txt8n++7VOjDRrdO/QJdw5p+2d/7tVFzSlxf5
eMW7FLjL5SDKgMPHz5BkgRMgdpsH6aLCSk929yCxDx9x+I3z57Rdj75HGcVS
1GX10zNOifJjSjF3wj8gC+8PoM2NiP4djkcNVbfXdu7Rv+4OQ2zQm0RqmIsi
pRyIA+CH17/TbAtvp4GqnQ7XtxSxN/kw93yizOI1vgUV1UC2gZRsuoLk6xuN
d1FbvnAXCtQ1VCMiJKNOFUyv0omI/fNqp5qHV1S9GZUXxAA57xR6u/otGR21
XCrGwzyfQL6OtCIHenB+WJowVqExhV4pgLHUobLZsAsByJxgwGXWS8NEGiJn
dfjAcfDgNy+DCM2RdHj5VKkxfakxUQTbjv2Lm08Oq3rKkg7ILXA53buvEKuv
hDgft9HIVj1p2kc4x+MNGheKea4jPwQcVykrrRWoXOAw1Y7F/6K6DDn/hW8/
ZSeIlM4hk0cUgbQ9k9KgFXCJHOhrhnIt3keBmdrehihRAoZ+nwaOMaNQnvAt
93HJdUrHjgzX8uH+Ycmim1ivh7kD6z0LAUJQSdlk7BlnM7PZdkQ6h76xkdW7
0V8d46zTL1s+Eu+aBiEG6jZESlZKz6q17T+fJyfER7N0A6b2jY6OuluRpP7c
aGk7Qy0iYD7xWYeBtkUWxdaanGKagOXzrDyMkvDwEoy0w+HosB4lRKGBlAzT
7GoUu/zyYFRYE184dlU4XPlA15uZtxRt32+PK64YSQX0CfSmxAHKw0Fm+7O2
PN13JQ1VH02KCjBPGQIf23PSALbZCUzAHnkOk4jScxyCYOSSqz1yMaDs+OeF
MgXq5TuiUUD1vh+ECk6IhyBjj7ld2gYyo2s/x4Td1gImBc/4sOZC4OWOuGbY
zHvb0Rt0UKVFFY3soN0+GtIFK7d1skX7i3wnXV+rylc9/CvsV774tAhwA8f2
RiGCr2WZqt1S9tmSw6BiQ2Iv+m1AOUFn92e9FjvbECVhANMnUFof9Bzl30QQ
AYgecsuwYtqxQUfW2+z1NsuRQl4VHDVHIvyQvdU8SCbJT3y8WDkHIf7lm7Lw
DJPf8sjlceki8wH9DQtxpOwl8W3guh5qX3BWiscIZeZVsuIByFjnkwiAPKez
4LrGI31+e3x1QOeJ/f/6OArFOK9EJlLtB7BzEA49dWd7Bq3hOE/wzIREhpJE
eiaEEbkClQQ1fcKAyllRqz3pVQ+Lx87kvAmZ7IGo3h+9jv5UuIkyWBcHdNPb
pKo2mm+6va9a63xjZ6NZV4XU/Q/K27EBOJcmVQJyaArCM/FC0Z+zgtDcLVlq
pyMWn0+RMvUb8IKKGLrAiFM8hb9tzPPoTn0erZeMw7ajcP0qHDleq7GXbw95
cMzlaIKs90eZgnit7DGFUjfAER/OHNy30gaQ+6LaJPkJMTPnhp97T4qeEr/r
ymiGXEuXuTNJGUYJ32JyfVjX91ifnrWKd1zJ0DxoytTyD799D3OSqv5g7v0v
Ykz/Bc5wpyvSaRSEClseMnE51mfB0wHNmWTrTSsDjvUcu8MhzIsVwxz7tNnx
Ws+qD0z/8GbX084yjzZE13IRIoykrLsirNYuBjM7n38hvs+pulzYA8AoeZFl
tP5tCgkxDApyJ3Q8AGJs1vxBUzAMFV3gxVlDOYiFngnJqtAD7Oo2K5kWA0F+
tpeqctCbzuWjmhatOb5WSnPL7IkxpLJmL9X6XuD65gm7dxz1Vl2Gw4bAWz10
4WP/HVkf/3EsfJZ8IyNSAgqJC2Maad7qlBlHG1+jsHVMpN+fFhlX9RCqWQjk
smVreVRWBXHivOw16j9elEcO5+c6/O4IFV3OBVOAdJIRRCZ0gChX4lDvBrlU
h0ZIKXEEDFv1ffVafA4Mdt8cojB3iOTPyWB0kFp4BGp34U91o1U3O9J112gb
WKV0ESEzl9v58qUmB8XnOwj5KJWZwUcQqMjwepoySgd3nqLP56461z93VHV0
M6U7m9D/subteDaIbVtESXE7r0AuznvXgxhdYAh1QWJywtCgKLY5lg1EZh3I
ymMe+DeyW/b8LgYTLI+y8MVABknblVyAy3CKipeLNP7jSscoTTJUEEoF17e8
ktnjkODm4lej7a7hx+uKYngLTc6Cbx+r+g2AlGom+FzB9fNNpe4YB5ElCK4m
tFpdDZ3f1NWhXlijaSbnaJnUZG/CErRDVmjGhUn6/KMh78/zCWIBrLdoaXuE
jiQRlNmQS1HDYgahgzKZcs4uGfStbKLGffhfRTJBdUF4Xqs45HtRenPy94ID
qU9mJzF6TWM5cwmh5DBElX1KWCto0TGrkVCnlcJDgL1u2unvoDgM0ZSJZl7Z
+gpKwogTCmz1Y7Q4r88fACVEwlbgq9lYoF1SsBPVQ2rvg0IUrT6OF89D7o71
UG+BmxPl2Jv4uWf+EANMRLfgChtJU3iHOMrCP5v02/ymDYhY3R5eYxM/EX1c
dV+7lGSXY1+phJ7EnIKQwGb5H5KzjWJ9b8prShpSR1bXfPOM4rHhSIWVIvIs
OrNMYHPuttxDL4/H3MIPrlVxsSVBPaL8qypO3jBXoqb2pG8SbCTF6ZDh0Fg2
ATdeEfnioo5e6dQBZXQKXDNbmImlxmiMuRkXXl29/0zQFkbRGwmUlfPvd2DV
2/33xYRhnJQb021++5cHNof/Y49dFSKAbv8FYqWMLud8t5T7Ky/4Ho87RIFG
jsgTsn/D0V94gbSk0peqzYueFWTWRFkYT77pnZtOZOt0izheHt4+o689QwhA
dKm4oC/7YzF3tEBhra4O+U5DkOlyBoSvEIRUCFjf3XFs2fWKqEz+0Ypu7Suf
229JM1WJjqlsJJqiKJb0yKybognhI+jCo0LcIJQAOLFI1z+ADKvjtbAWXpXc
jP0b788quI6SvUnQZ9XawVxtUs2G5ImGoTNV/xFJ5fbuJJx1o1u4Ww53YkGv
N9Xlf/ojS8Z/rLvIGwHxHEfnCTgu8BOATOsShxoTu0o/IWufnVzqbwW9uisO
bDVfAUUWyLmYoyPHQ/Am08Qvw1CkP0bU+4LTrDBLf5cTcuwh5kcwyR7JRP3g
gkMn1bebk774U5hbk+U3C48+ihd2TDMAni1kAODEagLTrCo4k75lNaK4hggN
BIH3QUME26ucDqMcymzlQT4vzHnUdZrNsphtgos2I/E/t60hyDPsVAtVCXsG
4IFLnw7nBjWw9lm45XWCs/tXXBpbxXo8CPrthpWybCUVPRZgvisAn2DuMsk/
eNt2cdL1o7j2eJdWalco08xaxoBsHHjkRZkm1H8BoFyawMDVrwf4DGR12xmL
Toacfum2XOADtveds+tZZZjOS/ACFxfZvUlSsIKIPg1SpMS//XLqjPSb4Msz
Eo0WK0f6V1ikZ93cElpbD2jirsaMiU6qZ8oKQVYpvKtLMccUcrm0v/3qPpN7
Tlcgci4LsNXrg6XGoH7Yxx85GkxYnNGT3CMe9iNqTj8DsZ5gywace/Kr+Nmf
ZnLb2EyhqGzMDwU9OlBormTUaiWZuFB73hSBl8UHOZ243ddpC97/OYoNMtAx
FfAk5AsCftGSdpT6MZki6XynvaNkLwRxKV5EcoDzqJtZJYfCKYhRj6M7EpMf
mc+jU04fZEcAy/CTfn+gLJMSsSB45yGrwj1kqswdd1aSgUPAiVvmgIIO+U8J
KFARnnt2FuqTbctP0mltq3bF5d86UZ5hJ7iUuUiFDFALaUo8KPUntMieidAk
3gaIKvlBndbKhF+Puj3FvX3yT7Sq8H1AEEpQEMSQjrnq5M78jHW0fBBYHc/2
+T6wZrsNB+MQuMMDw7jY3A/vSt+ghywchkqng5L38G499NqbZHa3tCUgzorX
mmPAEr873tZY/JTtHq1wGvIEU/v68/106ifzlH7l7jKVZaEink/OT871z1Sy
Ydd64H7PHf2DMG/XCQ6f4NS3T75jRNhIwTbywzp9npDkCtsqJrCgpDez9ze+
XMnbOqqSS5Xl9uRs+IRoNsxINjHG7IzAy46YCvJtcge9vChLWnTGhjZSeaY7
zcs9bzUZBXDdn9U5B0f+k0VHWbd/wQsrBt/XZWWX9vP7QAjlTGfyoYmxuE18
5DjMJpgo1KquJj8yZcN4PcXGFHgM9+/evK+YdaWS1E7Yr5glyMGVDxJDi4ZG
tstttrMSPbxOtpVK8C1TsNBISmOuJcu0/GX+pnDrwTVwXI/OTAvx4Cd3QeyC
4lYvHRY8ioHAn+392rJu/Bo5LNd4vcufyiPqkcSTaCkc+bQr2qSCNbJSMivD
Z2T8t9SviROSxYGMoElONZm6wi9bvpYw+d5nlM/hF7mmMakYLNfqTcGykxoS
7YpARXf6QtJcCpaByzec6KeTTGLutpDybwlAB59mQnUnDogocYWV4fcXmYlw
odaMIWWO+QUvlmht4pK3u1NkzojXZUvtKY9RP5rrRZVZI3HLHsdNwyciead8
ezRtbhkraob0KnpjD/OdcsOafyrby2zbvqX5I2svQJoYj2nPXLeA599ZW3wA
qtXor6vErctCGhmIX+T/f9ey8xBbG6NA59k/gJ8UvUPZWHHzQz0OLPs11UoU
qojJAFWDESS+4H2oylNshxR256nFZTRW9UV5K7ABRJirGwEmPDesT4I8vbp/
7rAJ+SKGoUS/DgLeDNLhdVZf8pddJ7O9ORinEcDAS8UsQ8Pv0zJClwKjn5g9
Cqi+UN9o28upljTdCLDTgR9Rr9sq6hvWjR7rP2AMPAYwf2tlNVHJx9Z57Wic
wtz9MfG+41pRvL8Um9i1SDSQU+2O5GU3A8Q9vxaWAzofIBs7NjTPs/dt3bqg
VwLQmxB5bJNq21Swj8RJE8AVwlqxUJceL2/2lZ5BTfATxHZBceirJGL1L6oz
EQIrMeVAlNOM7bQ5oKy4achFWuzWzZMo19NyZd5BawIMj5FOPTNfUqwZFIfw
xsA3rTkQN68o0VH6yhcieExN5Kk68nAcRRupxy8OTERekCYTLpG6vZFhCosg
W/VZkLGz1VY/MTMkCBWtMvICvzP9ws6s8zEdNuNcnmDijH/K9BuDW1yGQz5W
iII+XDYxVOfXvOSaLoEpxqzngYW4Sht+zVMoFOtWO1Qeu8//z7/nv+RVymB+
gE8x2XYPBTjat4a/X9/wjI2uJ1LXNdZepmTTjHpd2ZLydpkriSdRtXGe6/Mg
bci1y+lK6evNEyABB9Ys6DANXUd3yBzSBYqHJb4na9ESzKisxK5ghjk+31Vr
TcUDD3jvcvH7L/cHLaEu9cu3qxqBWCjK20Va0g/U603n+5nGWkKz+h7A2cg9
Buc5a13qtitgE+NRoe/thgHyYIFvkzJiWVV3122XPq7vS0dnzqs2zB5CM4WV
MqLutYCgpRi/gZy0Pk+9QyKIOfqoq3Dsd861MFlawB7VtUE8l01oIOlDFdKR
diSiOY7vK3Sv+64LVVkPfv/wfHY6Ky42Q5+oEXWBVg2fIdtQYKUzOyZTAnf0
sYL2jpQQZAplMdcijbjWmkuPMCZ9+t/q3GbcKDAHAyAEHrvNISxbm91Ouk6R
sYZFZ02x0ahGr7N/3owW5AEckOcSosQO+x7srV90lU6P2koSFeFKyVwVvbVk
r4hyH/pHpaFi09YSWcLzhgt0Ucn27PC9c+4fwuZQoMxehrfaQR+hKIe/kttV
DRokwJkj0p9AU8w72WEStgIuDhGa8+tKykkWmw+68j6OjtYw+fYAr+v+GIRI
lDk+LkKJtGFPt49q8EVLCwFUcbolfRzBTAetu87xAanVMQDGch3zmWVroXsk
tFaedYkt5FOTGr+06KUJEdIWmjKPDRtqwVOEegth9kXAplJ1IVfGG1lI06Y1
8/blciCUaBrikwXzHxLOskEpviZJUBsIN9oajKGqFxFwzoQjEC0J7vEr81Eh
baEAP/DuzF5cUY3UlhkQCjGOl1Dc6IM7QXjCTfRwx1Vzx3v9JCksL3W1M4kO
f3QpaPIGtNyT7kQHCS8r1UFWlObUxTfoBmXW8GKPWso648X6IoxBt8XoRmSc
JBKGmjMdhW+Nk81yVNVRkktkjW/1ToIIokDLMuFlUsIuVZawVAlbviAE13wc
WuooZBqu5pFcxJ5B3ScKL7ssxD/wsVbeaMEGPUy3Zj5ZFaU4LoQn7vUpjukW
aaB+6Ki8GRSCwDa3PT5RZ1bFDzI6znCC2pILdhX3nWsSPpTJ7wEQvQRySt75
H/8GYG9VFJsq31HZ3uALe4DvlYv7M1GkDMpehqW1H+X1HGFvYklrV830QJ0R
BDwPLrYSNRuCiq4LYdV6ehH9fwHeDTSFRme9BTPFAXRAbV52axju9eL63gnJ
ZD3PNOsepmFx2nTs7YjSFIKM++5AuRL5xH4BiVW8F6ExokBgWpF0fn5D3Iwz
v0fYH73HehanKREa8aojOSpzNTwc75nGZch+ZBC78+rc/kS3Q7/kCINP/DoJ
iliSJM8sdwRidldQgKYsiM8+iwhIkZr1Lo7LJ9ozUKKnoYcxl8TBmlH/tLYY
8rksgtxB4Tbr3yciSHetIG/CcxTp/4UzTNco5x9bmE7jQhX5Mlnlrvh3gSmB
qSHzoIbNc4wjfsTIvxvtTXnUuhKKuOdLwUq9XjOoqtJODo9UWnUFZehYywaW
c2hsrqCR+HaOG3yTVAML4wxXLM4HOzCfTI/Dd2iJM47zsIevdC6a8OIRr8TL
o+xiXLEjPd6KbwSsL1GfR7uCisa9v+YeSTPdwG+7pSAKDTZnbpL8/PRtjsi/
uDwIISaJvoCPVueh9Jr0Eox4FDfyCaYQEkxBW+bo+R5ouUl60ckYuohxC889
RujucghQuyYZ2Fkh/afx6R/EUpsjjJv1lMcoXbIQR9Q/YgDHFZ53WyOoRjW8
G2qwqLwBSAKcMIBRPjAshnsAb+/DQD792Pyfyj1Z8VEKKuLafWsxMukLbcKo
HHR7Mdq84oXg/DFbWEr1jK4vQUbeixt/3PNDzBYy2o/lpF+AVwd1TLDH6jGz
WAdLMTymcMrZPk4a6jRIA/42vFyeHwBb2z1+48mp5PNc5MK/jNG+1Y4WySOO
+/0jjS6GXoj7OrBabujb8YI4Xz2GIoINM6uWKbwVrxVzx+uLd2LgI4iKO/sp
0oORAed0N6VTRP5o84B+1cxhKx+StM+crKmPp42PTlVphTmGWMMefz2jNMEp
xnAgHfvCuUMVOMt7167lR+3Cg04ASGQs7Xewh/A9KL4LGNAa5Fduw2oB8S5g
HUxWbXPkycoKENn1HxMSD34bwWvzfX7msCcy9QAP7DGI1ETgZvXTadnbDsg0
8pt/OxBJyQ1ien5p4/ZKtQftMFPnqMQvAm57SCd6UkuWsQe3uHvpjVsWtVk9
eaGsXHoonCQQZo83WwPxiBV797O9SIvYyzA3fd3ihv0NiTtG3X6XWArqtnCi
B8dMDj/QjmBZax3/KsrNLQLA28DGNbieDZcs+HzRSHC76SQ2VPfVGv5Jm0KZ
Zn9IIYzyitsKD8j0aEyuH8dQoF5iZEjyr6UwI2GmIY4DdklmbOjVF4633DwE
ZWLcjgbsMdVHUFZlSgOwIY8iXK9oEOzuJ9sytkydU6U9zQ9SSRtkEhZVzn6V
CjJbODd/Acoix2NJkwK9CQDa06TLJyKXQZ14rcYJN/qgtOji5WeVaB6f3ge3
QRz8u4LD5p2kuzbQHGEIeg0HAsUMJ/i3WctHHPNHP/O9DR76Wvu9sd9aSmGB
gKdodQqByyksra7Q2CT89SnTQ8/jjIYhbp7szTZUEU40twf+HTdhVZxTPCAJ
2JbXc8UB9wIsH8/6i7LjxpaI1m1q26DnFCovYyUNbG7O+ZxvJJ9HKYN08ACD
3+U6urSWWmwjrFBnWKDre0GkXH4X7vuqT+5TJH0jNc6tklDMQIjXrTasoHDg
EqxDZQqpOG0mbLVbnXiBNfeJ+YWyxG6M3+KfRPu/Itkr8AzCOSovCvI6iZkX
wCzhlrfQry+B2g7YshqUytb3nIOaEggBngrZ7Um4el9lTQQk/CX+jRFUWceQ
m2YL66TczAhzhikDaPrvXoSQkFd6yRb1BEzcOpVmOLCtr0xvJBuBdEgVLqi0
Z76FNCsBiWCbsMnPypnjtCDRcVnIi6fX9f9pQouxmjWegKXKGr6U7W0VD7eV
ROMDjxy1yPIGxuhqUOCfomQlqCl/9/V0dZUpzJMf9sfwZhgI2/ppuAZ2/96N
KT79/4DeeV0T2DzqIm+J4ceP8zV7COsnRYAPJtTKRLtsqyVa7g8iZCWVlH4F
UDOdbLT1bmn0rCqIImv5Iu5+qHqFlEfm9aGY3SMLBrlCZ5RRoBKfMMf1KNhT
5yyCBoz4Ar8rdkCOsVH5JBEwYkUJgZVCtWGmeq1RnUokw954zkqtLNAvN8sz
kvg0sehTQOIEgynQiIQQrYDD0YEtQFT1CSTfVKDMqXZ/mn724z0biOSmu4Y4
ntA/faSB92bNRVE159aqEoozX4u6xE1zmWs3yOxNcYKXhIDIUVd71NjwYA6M
7LCCD1Q21a1q5KwCC6q4xPy8rOSG5+g+uq7Q7v5Zc4hBwq2GQ7zlaFhNFUGt
dIHsm+T2ow2DRkHwetr7todbxloIIeu5/r0aX0Lxge1GtC0luGN/8oTso2PQ
eyoYExUycu84dMdKzMvL4Orl33xd4s7jMa1HIGWdVdSED/B115Dns6AIPFM4
/TAbwIK3dsclM/xiW5QK2RqTHwyO8aVI14NvDN6ycxpRazcVyhkW87kzTQ5C
z0tm1jD+UaKGP+R9aX6Xm+6LqGnO/rtUCBIjBOAplVOq9QXzb3F4bQOn5PeN
9dC+3vhmzfX8SWYLShUjpq+c0Cjy1MThTa/J16ew8kg/ankwxE+aR03nDZnj
HmvKVmFPpOMTYsUDFEj66E72SYYaoCAtg+g6BXCJnf9lbtqJbz/idHn93dt8
Ig3wmvIj9vOVUzlwC8iKa7KZhFxmToOGXcpJHB8gZU3btK1vJKSj68Np96n4
JPCoUVhoLxfs1keqvc2p7rlIfc0Fs0rryqm+NOR1pmYzX0jGya4PVgvDHGEO
sA3UqzEHszfDHhupOTz0s0pzCsSs+4kZqYJAkKmxHicHfZ5Em0l6KD+/R47a
yrJqkgxO/pqLFYUkI+aKBrtjB3TVzXqN2Y7BXt+sAJatMNuPeglQQoripE8D
oXcAhcwKOeiylFQx/5r4iqe6FiByaW1yuNNIa/nWR+dUPA+OqIkJYnLK0Ciw
N+3Ds4KeTeiwUEx1bHHWXV32mEbQKkT3MCVsVl7kuudx5/ENCvXC2P3jNiYG
X9xdXugT/E6tDaM/bbruwmG9BcFXSlmrKX6etKH9We/IJ/M3X7JTlOMz3zqv
5E6XNutGlGqT6vALzU8ebtBhdAv7HpScmayY2Y+N6feXni4tCaZMVKeQkaf0
N799/vXqYR2FYqUC/bWOvaPfRzdQKebyuQt5XecOEo0VkA9MdqTU+ZmKNlbd
rM6x8rVruabTiZNZ/BnUdWu869jZr5ZJZiNoakc7O+CeB/MnCugfSI+eQoh9
+6oFduPtVy0H9p3KR9zAKkIn2Z1NO5d+oGuwnPffEmLer6jtNCMwEMqqmNE8
Fqmyu5BExuzTN9gL9DAp0jZxp6yuXaWRaNdWljcfqHlqiJXy6o0i4nMiMvuE
+3wTVlCfL51aOzNwMjRo+8eh4dLSA7aGsh6d5i0+N06F9aTh97StVGwx3LIN
jIU3anAfCyvJviHriWF/bA5lFQ85tOEQtxXyWhCeavSN8/dK/m8XkF7QeW+9
k1hYVyV+HtN5BqIxi2QdUv34wi5WqIX4FxtEV7e0chP7OxRO8pJjLSH36vZL
3Oj9DemfHX6K10coqRkjaUHog068l7BwvxYX0Tv6Rm5MW7x50MF5UR/fUAAw
kAbH4JLPlmMOdeVg9SLGMyyCVpZLBEbbHMGwMpKPpzo5PgMkZKR3mylooE4o
kkTUAov53ddEIPRCjQYCOvOQR/hqbpyzjVuUS9jJkR3J7/Gw42iT2Wnz6PDv
cn+3ozkilSzzoEwfPMBcCAja811REhGp0OrehieBYqcxuc+QIJ4duoxp1PLf
HbyOs1Nnsx8lBntxWelyceiu2yqKZiFZbt/nXZ7vbZ54ypMU2gQZtKXhZdrY
03dvS2Aj0YUMRf5RJJGFmhAztn3iZqOjTREVtnJT9L8yIEGu+wYPjHgTaUU6
gocxFjifl4yU+kNor8oj8rV6bt4eGZalqs+Ays2rr6wdb7SCzjhf/F6lt9GN
oRFPQyTisjDiPLo2Yefa/4XqWKQIhCWE66OA1o8D3bR3r0BLotNgP28InwmS
V0usV9PLgPe20BCPCeERPn8hssBdffrxcaVzGI95eouUKltx30LFxnLX+dYW
CyALWN6gAAc94eiYL+1A7T1BfJW9IKc5l/a4pEioXngrRk98tCpELIXVG/L6
H0WSUTDvsG9NnnOJNllm5y2T4tFQYWY7jvboLSk6qqZGBwF+MtBJL22i11OR
SU1XBjK7vY4mzPjeIJJGP8pVLJaBNM/zbdh43CyhnC7PiNteHSB+4QK2k6WX
I02BqEOYTnhYRk1H6rNYUWyeGvdblm5C79p3uDvyOIPaT9TT9EDuwrM1ZG/T
HEyytSuCTqm+bDmtITsEBW3ZHz4isQrCa927/h9OkAstSHdwIZMFyNgiN8A8
IyRezGZVasiVPFHNDGmzB9F5oVn7iTIwwdcg6M5rM1Neqh7yENXAybC9BWBx
GBPysLAn8NIzKDy01/+w6cIUePiTIWmMORyTfXflxVup/mDrnGjvOjrIlalA
+vAnHRZZaHqTIHksn2E67RgHyJWiEhc+ZcG+4rU7qlTy5tCjvTZvInKgfSAR
6JcGGuzpnml8jBtI/w7UKxTm5mnWmvuM3MmSDpQBwqZOAoWOma6X2Wltoexq
smhVXQze82pqqKwTXyVV4lkDS7cymQHKd2mNyLgM10xDbvFxSYj4pd5ECJXE
mmrQICtx/zxSMiRBxZDjp7h9vmlW/+0TR8eiOohzSStWzpBu3N9snkNDIGqF
wp1Ono3WVy4TZP99DpL+N+fQn6QPoMGF3p4FL+6gint98plyzXFZe0FuHzc7
fKuyGAOXfsy4I3DoRkbdeLCSorcXNuNlFMZLSRSL1WrtwmCQ85PIsge0jdai
K2mcHheG45C55Paykp9o42VWLlHjZ5wdgKy2qeMPiwMrkV3dHFSGR7VA8ChP
YHogePPofBamN7lF3Lsy+ocjEOEpSEetyvH4HQ873NGjC9ZwAVr9Yng3CvL1
Jzyv5ZGByltg6z5cqaUWbToGEfdES8YEvYtDwlkPW8RAd33Q5U58j/dXc4Jj
aipHkE8oKItDDamZQjy+5Fujr/fa2EtwDbh4nDKDlrdgS/TKQZ7sVedk+gCb
p23/EMfd/BUOFJFnFiVfioevfx9LZ8gnBOJwkVdrZR6p6vWFDoMjaZ0tixwG
Psmw9iOZEq+e/Plb5zEt0YgmBLcJacIyILZJYC7QMslvK6fH21Bmw9H1Prih
yrqqP0LkZe9LdDTeu7yFNeNmPC+7xsAFfKQCviBh1qYMi3fPk3nvW35qgZxL
2Dd1yl3HpjQ3th/K1/DW/BF+mMoxcLJqt31e02A8oX5T5wnX+FD/Vyb3LDcZ
VQwTC/Rozb3DUcs3BV2rwNSOqxLlU73bGoDcMMRBxOWyz7lI/1xknXwPMQuy
z6GmL9Quy6Bz2hzuZbM3D6OAzO0aXotUQfq3D8zmPrFermJNPqF0tBRaoFbv
WaNFD3Am8jUhT0uK3rm2OBPSM4WlhlCzKh53rCzlPUgfV25N1ScodjVCVGeW
bPuadDAQXLkDwh/dAs7gGz6zUH8Uw59vLxkLLXdgD94d7PHdu9doqRJejfbl
9BFLDeumJzI+wg6nhgn2aa1riGWMo5tZtYFuuZukL+r59zSy/5Up47xJKYo6
LsRF8bhF2J46Mx+uRFTYAdffx+5SKEtwDv8KUNvzW8FBHtqCDsjzlhiryQay
PXcOCK8dthm+IEr7zJijNMvHryUM+Hl5HITFkMW6v8LebNwf8lPDwSIt+Egd
iz0HC8SXOKMaahnllPckdg8MWkkfDuueQeMzJeK9QIZnLIS1Bl0IdtJSdeq6
4RcNzvOcxaUY8LEPfYnqUVGqnbv3LReDCkXleWJzLNb9YEJZRRSZ0LDxefL6
Zm4h+VGjBLp29SVOnoN85mwxug8qEjec3kFVJJYVE6j8cTzgZevu6pns/TSJ
XyJz/uVtWFIvhYIOUd+T7olWPzuf+4Br4CSOFx9CTwmxB1KgOMYq3Eceht0X
fXdHS8Hfgw9i2lZbDa75Y9gQ0EOipzwx24LvaqYgnOgeHceFn6u1CEBcf/TH
MLzZrRRv8bBRM3/YwmIetYK9uFVOi6pcIOnwAF7H+5L+Y15yNvn653jOou8G
a3j3y+GfT9aXYAldg5kWFpnvumdOEvS19NX9qd+u5H6Vtbc4XS6jNwmfKb3C
cUJsfgBBJNVPi5jXKYcIHXIn1fupz+JuwIFKTPAdqxF3S3ZVfiFk9kipHZqL
KWc+KVSVh1fiTWPK153R64/MLAYUmkPci/Bhh9HYXC5sE6cpyzEb3sf5+/qM
cHCumye6EJTNDlSTDqEe9QpOTRDsFBFIgatr0OhVB2hMTnT47YRwU0Owh6Oo
a9Q9huEwpvn96580CmnaY747aqjI57RNcuqYl14MMtFlcO5XG9G3MrLeaUmW
Ka/+BhcQ9FEPhSTf9awvkehsHo5NryrBSOtMhrKiZutsZGgKzkIAhs+oBqEV
aiHLdyV8iArWwKkiIUxf9cJ/mEnJUKymJu77yf/EIspVpJ8HlmCru/rk2bqr
V72YVwPiNWxsSPKH0fSsrrPzM1ayGb8xaFNApuY9bFl5YEwOjsObZCUs8qlD
OFAiBMc+S1ByJSP20lh6N6u+cc4SNNfFEmzQeyW58L3J/2tz1DxTFQrYtzpW
dckjjGIGcgRMFvCNnvbsPGMjJzJH2FIxcrGMmK1E0d0YgeoVEf41AocpfBFE
gCfGG/QH6pzaRxduJQ61rBs1YAem1DIrjrcntZ/zcYLdO3DMXbBVi4fmbPYM
0lCyDugD7SwS6wVHCAZBUt8HxfEiU85V1QLKwx5uwRXiUrz4dof2N6a5ACS6
ELyv1rqbG12XH7H8BDBobo6zA6/gYRjPmhdnG4N4FE5o76Mx5j0rgu4T3fc8
itry18yIW+cHXOUBceXL/kEK5hvgjcWd4ecqKcBkaJ8jd3TIg1UfrRsS1EPg
+zLcBIb+5XVlSYP3/cXA8pcVfTw1U4PWY41OoMAS3z/TuVGfO0/yNHWt/r0/
ZAZ2T1ctZsrbc7+fDRJLNimbt4UGCMpyYTuFoMB91ECpQzbZt/KeeJCsufpj
6CNiIsrjE9eza/YUnFuKHdvtGwoVIA946O+rxSje/NN6j0JHN55ipOhqdFou
AaPEN1WaB+wx87m+R8dV/lXJ/1h5S+dVlVtFD+vnTlNkvRTQ9Iw9TOlbvuox
l55P1K74rTmd9HBReAV6iHRQMdjk0k6i6pAkAPbfGKD8nSIYl6YBueI37Dm+
arzn4KuwGGiuBIh16OpdJpJyGX5gWqdEvCijC/znNmlL4vSbvjS8p1QWIUjK
qSM1XT+zfEPzVe9X3Objd9T6THgPEPujmcUYsNxobvfOd3mVeyTAJJCjjoWZ
f/5Dm/Nfg8P0cqn2t2Zpfyk/iFU/GNLLXIBTMaAtuQ9w129V0W/FzXUpGXo1
9pMaxrkqOVcl1vigfBKS09ZW0WXu7m76g2veHRw52NU8Lnu5BhYCOSAPqKhM
N8UiVSy7pZVS44+1re8yOzdTOlTKX+jGgZLhCAb/N6rpZkrzKjrzVnn5+AwP
4MOnt/BZ/BaWoYdEMUS4okFUzi1bnJISxB/klWp6Y/QsQwYk9FTqWAPANSgU
+8GZWlq97arYUMfY+RgEW19yfJXUIaRodK/meohnfxOGxi2hZpV21EWDIg4Q
/vBCZuNQMDINHY42yyBs8xr7/XEAVEFm0kKvgbfRBat1FiMgHYO++4la5lxb
/USbzha2VkJzEZDXXsPQwQy5xmXEXHA6FbiGBRIpilKWWFzqa+5YmA8kZcu3
jXMqczeh2vz+q8VxvRAF4UbNcBs0Z6cg+qJjaTcHDOv7e2G/2yL5bYiV5/7w
gga7h3N9JOCB62NLtYwpyuHIpigp9gInQMtAvHL8CxTHWPIC49inzsSGDBjX
Tr1kFdbm4UYgLW1DJCxr6M+6S5qLVsWtXDUeoiRnlnCZy9oERUKGmleqxivb
bL4lyTplKf+QcfZqyWjztCaPemWuMVoEgfCI1JwrNZLWl5jMjMMuRQgUNoI/
ojxeCfeaNP1S4LhRgk9HfHp54WGSYZVuI9gr5j7cllBWS59Knyi8MuBtXVKL
ESuRwVMvMh1ydplcuZMUULjxedHx40RnI8EM7nIidJhkojbcN97ykylxLXlU
ybXscCtRxjErvVg69M+XkgCQOtIzTbBOewbGxHbJupk8USERhGw+NytbAb+t
mR5nkoPT1o//wqLMzMBMQcViO5uBlW9HUhN4B43z5cFRxe01rsCJhi5tU3Jv
4TDq6ZaNtZYk3NqZ6ySYJau0uWSywAH9h4Xak9SJe0Yml+Gt57phKrLxlsTK
I6mMFKw+9eoqIyRlSg+OIu/FgbsKJvMOJ8JL8s3i/4cWnQydEhDwIPIS0scc
Bf7POBxFg0dPG1o8hZA82oJgk3eQjwn9fqQUklVyAHLZg8YdtoyRmOK1eADL
oIz//fK+KpQNNcLLF0MS0B2OXMFfKn1b9bkSqCwHooDSOg5rxMK266R8YS7I
OuS9v2I5YdSivRzeqO2Ht7Api0K3O6kUfE4qD58CZ37cAoXfyBiIf+yDG9a9
kBWELMSEL+T6nkpp4k3rVdhtSiqzvwZaJTsaNk0dzI9FM0GGKyWFA/uVdzQU
MMcu7xHqwo8bV4MaaMaY3OCfQSWreDW0L5v+67uVMCihONTMKV2ev6LWKekc
/nTPMPGwZqCJZblRVbuHcE/PUiK8F5jctHvRCNas/iEtSOCNDA4ySxFvc3z0
kiWmWr2bFW87MqL5tXVm+gAKuuClz3tcYdHE/qs2j93KSEYhEPlp8wNS0hcL
aFrw26EDEB6xkQe9LZq9f6MF5oCygIuudK2zPXv6jSCojN30JLpTQVvgSnIN
VUhIHnGg9rYJxD1gny3Dn2xawBnGRsIqVzU7371p6K4KBuqD2QO2wx+atSH6
dFr8bSMegAulT9q5urltBx1UjEZrLnFHcaWBTJDlMWH3RrBBZBGvxvJ3H6da
4Zm2DXbLOMxI9/blu6I7GOZ1ZqSXf7QSWvx4Nybatio4KcpTNyqTIj0QV7Ov
9zCvGeqtcAbyaLEdhQoaHETRkKuOK3i+Sjr7LLy+OM6+o6tp7zMHmd/Jo+7M
TBBlvo2jjSxmjJhFUGBKQ/lDrEHs3jRgdLQy4fiWvIozq8OKhNYt/Uggnssh
hGiPB0nRQ/oKZqws0fkuebvZE6P3kKW8shE2BxQH/92vSmcZJ38XgibQ7DNq
sd2KbGvcYJ03iZzaD0XwDDqW9/woLltrrePurOl1p1m0qTgBJRtxcm649XlF
ddtZQUZcRKzNd6oP6AJHvqoeD1BuWsvkvBllBcUpbvMuXiiO6p0sqY67I6KU
Jn9zHBaQTxCPlSR4uYeok2/lbofyZERyAMGm8CPICxeniYYsSFPbbK8JRNdB
DmwnL3oJZSZElOStizMyCw/kfWMx7+heJXbnnQ0Is/kWrWFHGCm7Q7Izwf5N
9mG4hTL71fxLiAjrLvGjWsOFFTveSrgqvskYx9sKAvNZz/fDTuRzmcOAoWLd
nDzg8XNld/5frk6qQe5VLxg1DgA/51Gz26lETTll7mVTpdfO2y8Kter7WGu+
388cgUVIB3RCxy11cpIw0+PMmAOdd//4tHQXVLWyRAzt0uXaaxfEgUw3wWsf
lCHsdOT7B12rqd1+iDKGnlEc5VHE3WPnN31qgu1VgPb/16uS/reoneFtIWkd
Lbbu9kMxENcFGwEXIkB+qWN7xab9b2Ha7C/jZM/VYXxihodMwPdX+p/QBHQB
vQoYb4lvnnrF9WJDfUbE0psA29wCLmGS+MNhT28zHi5TluznwXLv3u+OH20P
LTaWC84FVuxQCfKdbaVg0kG8op+GU7ao96Ji7rWCQZZPv9Jn0Ina8FVl/M9N
pORZHXBjwknttuZE7peZt+oeck6IdRZLe7LNs22UuBorcmPTjhntjezeu8O+
Prjl/8nwL+hWDB388+u6T+0ii5tyTIxEiT6jQn9MiS5vX5KXlFIM42rVBxKQ
354kCcE+qUfS5ZOibEKp/TIehegxLAH2re/5M10EyFFSNQHmBwlj3iLxvjBw
fN3snSLZUXf8bS94qE1SnsVZjfE+iBvcC4E6y/gwMO0SGIUJeRULR7zAhHr1
py0g66vFwwJn4DSEdfuw3+LwnDge30a4YMf2FsX+A++W/4aU2kY9UFpObQIy
1EGuxLZMDNJBxWbbHzQhYtgJxNLdZgFVU+s3BYtqOvzmYF54Hyu9Es1QE02u
Cffv8Ud4tp5QAXL2tNkEgLgE6qqza3oAyn2ByIsPo/bKMZEypjobXHxJlohZ
mEzahomXRW1TAvWT1WOKloeKFDAF8Q+UIwHRvykprQmgCxTriGn6Zfs0FMZE
Cx5jjQjDe7Xqg5qq4lm112YOWqB50Abg3+a+xQfe+daBEeFRLmK3QkRpnK/T
Pys+iK5uATn/OpQ2J+m1iK6FyBidtZjp7ByST4c4mkE1zE0EHQ8WwkkD/1Z+
o28GtKqsRNoicvdTl3HP9RorWPCfTv6vdv33pi8M/a8FOYGc5U+YrP1oTRAt
sPoYxJuAyoO46JleeRL4oFCMSXzqTvJMo/RlCLa/dtDDIR/Zm1lWrFkH7Jc0
J/k34TSagDr2qWGdiEUzD8ciLDLWk5luXJ3Yd2qmkh8EGAvwE/LlepOx4IJl
gtyHbGpkXwwSIq1kne/JvaA+RfOobf/+E9OW1p400l0wDUN+L4TE+lSXsWTe
lqJnZCeADH/A4B6y67iWGpjpkBgwzH9iu/tRfzQPPEaVrWwslCQL3Bw3vFze
G3JdsajoWU+mkAP8X/G7NJZG0lsSWdlW08v6Vpu0dLEI2VJ4NoZNiihQ2qT6
iuVa/cqneIrSJv/Uby0L2/g8/lCinuDpzljLBVDy59pTkxpKdnNomJA76FeX
pWhFd19fPlABnSpy5UbZSVWaMJkB7EiQtY+AtdwddUzz0O3WqgBx3tTaNYPF
qdSikN/LEifD7XcD9qwxR3uo9+bE7d78t9qakn1YHViWnhkHxQXc7D5joGYh
a3xjsoYFaYQ5ql0ugWVTzOSjXb8Yp3EPaR1rgK2Sz3xxsD3DH5tSojMxshVi
uef1UFzkGPyUScVsEwn7MyNC+WnMYlipplpTwCiE9UFf63sDo1FXhK6SH59f
JX11myS5+JvVuwvpvLDBDlhJ/pm8Mn0+y8Sk17dMOFNuXWenLfwKzSiZxmgn
aFnzqvvK9xx4Shi/CVic6NcidGzxiN6k1RNuKdamAi2UNwK1vUw+uAEDlS8Q
98RS7d7zeXcp6rWQphk1VcM9cXFdEULJlc0+HvcR2rWLmCpL1LudjT5rjfZg
cllix2C18ZtZdRU01E4WsmqOzOg3SqMmmp9pUzU5C1UvKDacgh5Yt1Eg1HEP
dkZo0qxmKHVwaOrAZyzYxz00nYgFG2JVPtqq4o49Fvt+rQW7EqJ15THG7YF7
MzUsuXq0OmN3EGpedQwOdX/YTrn3efCqHgJ8bhlcg3l3oIvF+lVgz4NIWz/2
nUIssXsNFCivXz/quHWlFjtnawdZ/Nu5dhmrkP3cSU5FcBY/j4yE6csVNQJ2
5m/IND90CJFwzl87M35kgzYkBxc9NdGkUqS4+ktlx9yRRJDTb9xlqRP60Af+
YrEgV0YqCc3judV5B+9+Q7SSW/ETGFRpY1LOZPFg8WU+R8Z+itnlI2BcH9FZ
0/YnPJ6bJhibsD33F3wroMR6aV7MmILAwsz4hQAh7rVgO0MTurwrfGQPUbqJ
DspjIxFDXblOMGV4Zg+ppX1o93Bv5QNMAHM2TQDiH4NWxN7taGNtkI1cos0x
u3/VTFHaiKbPZGOPgclzg8SRIBTd/fAE+sJgRHagepW2NQuuCLRraPMw50bi
3HJ9JYaOMbvrm/I9RqcNhB5a0DZh62vR5AGLcV2QOAy9fvHGoiyxXbCUnKG5
qBdy560S6M/0lrOKdy6XQJt2ZcDEIqQi8s5Vg12sJHKnCNxePHTML2dWw+rg
DOz6BCR+mtH/oHSsZyNGFfbj5gxGCczxLY27+/uLFUvl3PcfX8HaNNM8eoJt
k+qeOFYCQrZr/LxNZxKAaO4qmlMLvu8RcMYgJb8xBMBUur0G4Xwm3mTg38lI
iBcpjdHeHA2xsvjkEjmE/AY5uUNv36Lmyljp+zAY3Z3Ja4RTwivvTZ1kgNRv
W/dWYeZoTPz/kaXru5jpgm2vgwp/+xmmdV3+FUFlx3axteodSKeu3hG1OqDk
Mb/NXrQlPUfKq+QkkuBHK3mFXGK5V1fXDjk4k0TRsDhT9TbURxzUdWC/lQFk
3QI/mYwP/qsy/vJp5lRRhmMUwAhRn0ZHExqLgCvmKAsugAAblPo3AZTj4Oy/
uiHz94r0A4Qqg5mvTDN/8gBs8H2eoPKqlh4OJgP4IILO0PS+7p9IB6y6w5Uo
hcgqHzxXLOMov4Vjgs7HWapOSK3FySJmku/nJ0T0dA9BBReL/Gn7eYSfy9qf
JMSJ5GjfAUyLqrCYsQz1tqyhvhaWTnTMbQVc7D4T1zIe2WnMR6gOBXTOOh+x
SjTXeWxBvUex3kRjtFZRFcIz+V/rQbjEufmpDRKjk/+IxWylGDX3PcRMltzp
yK0thKLmKv9BeDecTQ2DyC+W7pSC6Z05jtksdMimMPF2BgLXgPXxCuhTYLLr
yfsBagbl1k/R/OzKRk7wXUcBc/9Jhy/F0+2mNW4HOi2y0o756dMoHfZjcOAN
uw+21Zeb6tX6qlWUfyKwJVPwMXbR57NlE4UUNQyIOyt99EDOREI9R2o/yEtr
DUqsWx870PUBAsQME8Kg5/sOgc8hwMK5GKFyaM+JYlfLoLhymrPqIQIrzvBq
XrC/zC6kzgJ57rftguRTkdLAQvzRds4iNFuSrppxEyiqZsUUyZvHNjgmL3A9
VFdmbSeyKFZnp5Ezefq37p/pZzQRc009kbaIG4vpiaCMXTcz/XdddjqB8fho
awn8DBOa4WsFuhB4pFkiF+dSQdrwzRkF7KkvkJDfbZXLZh8WLSlqOlT6gvnd
75VTwzG4hcQyJU8btcuZ8b2RA/4I4oJ2wmzeQENgi5GewUJ0BnIly48vSmO8
58r/DBDNByY5kf2rEQCtm7uYg1AIeuuhb99RuomtiLBfFI0NLa3FSQMJEaQ/
iwd3GmFJmdmb1L/RtHOkpWkONC3SAXKTtnm/hAgTUNo7eW5DLmxbZoG2EtDu
6uv/ikxNR/ffOZwijJ4cecIwv3vYX5iK5kRoGef9F+SKqxtNF3MdJ3mjB5WN
V4K061SHslq3IX8cl9eUBrETefYXs8NnqYzelw+Q/qNOCkhfd5ZhuyoGNyMW
3saeFF3rhkWPnaNCroiMW/I8dcTviLcQuMWRa0EkiyYLmVr2c4Ayx9cHtQEW
syqZyDigpSH69i7puDsz8U0Ftpw2DtKug82QI0fcHVwDTSx1CY5S19AGjH13
16yxkVoHwRTg2Fbdjbzk+pQBPc3AT8rw4u+ADg23kcu71xiTDgNZsWJI7gQm
Q4zSWvJdSeNgTrq6OEV+7WhfgfiQ8aWM2b0JZkzKumZH3WqJg7xOF8ZdVi0o
RK7RPSB+QrARrmTlym5Sfi4181eRqVSCRFkZ42srGQO+X8N3550E0ReC/JbB
71fJmUZ48mopCH3RICq7uE/KW6pYfLblNI21y81byUq+CXhCd2RLuZzFDIvD
5kdbUpmEt8d7mvarOAfxXDghSLWjXhwQMYpC2m1tysKbKhWCXVL9f23MZ+Co
MeU6jm2S8g3Llzv2VgO0cd9w0wincc3tSjawZVEjW0UAhwck/QepuvJNAyBt
QxW9kM3AV6Rd7cEeou+JJzRFqQbuxzPf6fKl1C/9val4yDU4GWUCWn09rxit
V/0CBpHzVWUHxVk9oVO/9H7CLhRLuq8SsncNmrvphxDDe455vDXouJRajS4p
zxTXjdH5dv+Q3KnimdNJX49inIXUjZTaZ7IRrEDqQquefidzMlQCswAhjYSt
FNZg20jJEL6XQzdsR20qH0NCfYY2b5rIJkdVG14wL0tsZMjGvbOG1L6DEvI5
buWcG18XnQUayb/ocmybw/iW5DSy3nFg6DdqOV3qPekT0myXroWU1w+O5qZU
59g0lzEFl9Dgu/28ZZ2v3Z/SA+lqE1sOFT2C428D5Ls9J+d9ENw8z0YaO3QK
mysmKOFvW2+stQwhOqFFyDAcmybjrMukVqgQybbA0RVewnLHbqE6sRTnc6QS
yoihMImwSVK3aN9qUM9nKACCzH+3/N91/cMRhq/R8wWP6CdW4xN31uEQUhxD
H8w2oZWOXWfeh8RQ8kGoespiQsjCR4twJeAgZOgbPcccurOCN2XR5dAKWinG
gGxWsX+qR3yE4av5QoqTgIJp8gZb1j0TjedMqG/pGuLXrmcm7FvaLiQcRs2G
KCPiGaa8MWZ7sjB5XtAPxN+9RyTDzfkUckdbWENvHqCQOBAt0qV1ixB62X4F
ODt+fTYRTSrefH6IH0pYiZUM5bHGHxbdTuoxdjG7JR2W2V0x0AyHv/94zO44
HYa1mQ2O2TEwHueK8xW7+wL1yKUI7EcFFz+x5ZrKSkZOMK1IiPRVVLTjM8fa
nOmB4PeZniziXsYixeejDnd7iUdWbzDf0QHdIYFTIDt1gaOagPQOw09knb9s
ocjZ1z3JbxAtZQUqYKj4kzRP0Gd/tVmrUKAtF0ccvm9kLXyhZHVOf1HwHBMG
vKjYsBPr133Zoan/GILc3OhI2oeREWSaawYNnpzHdqjBewUoXrnRNYkAmaRn
8YKv5FEwTJeuRorsSI41LVbe0rRr/uNBbzJ/KL/9S+4jFpLodDUNfNeABxjx
FhBv2SQGL8WUy9yfWP7PI5xIt3bgUEvHMp3ldyUwTeR+1416+6FiBE5y+vMi
B5wlf/3qoHeBeg1l6DbQ42OLrNuJfUtIfjfwBNlMISOtBgFE6KkzzuVYqESo
1hfWRnPYA4jSUimeZb6iOgs2n/Kx/yVYpXJE4lwzU37KWfJK4jzOMqIuIKYO
1Xzs3CzMYe3pEFISZNs3MnBTFpUJEM1ixxYNRcocodmglDLv46wcJao3Y4mG
s7Z9nOof1MaNlaoTzpnm0K3sO5gzqIgXEuZPCf1n/Hm/ktiS6ug4c0A+UUgD
31n5p6GSbyDLNUo3pbGI8OQmNWp+lqTNNrX+DIHgyqMlKlEFygJcrQZSzP9Q
RWVYes0gu3MJIB9/YiiYMdmeKGUZ5lUIyqrJSqDPMJ75oOcA5HnIdxjPUDbO
TlrRznkGq7I6qOLb7ioaisIoH8gRyfVSysI0EbRwSItPeMt2uWyqW0FN85Ov
GaeULNMMsh77nfsK1kXF/YgDntI4btFfUELJ1UKOuHyVOgWd8laUXyvd91Ah
w1BDssAMLxEYUKvY3zQwi8F3E8k8Nqa1y3iPRBj+YUthrNw1SxEhh0zMhZHS
zb7yHkpL/LLjYtUFsIOrkRlJ5j2UWEDYPiqgOOZEnHG95HM+JY5+PFWwYz6r
xFdGm/AEq/K46IYpRyLPnv6hfjXphBwvRirQrFc9vTK4UDefo0aYosAt3DNK
fa2d4OSle29HL/7j9Mg64YIF/niAVUZWhaX+yTI985IpJ+04IGkTVRToKike
GSIUwuI+C6cQcyogDAk7V5gi7sOu4OxBtwmSZmAxh96xIg74zYqSvcO1JibG
Hpu+EzvuxnA7rp2nzJIa9ECD01Kphcrt0RQJEEthDaIu9+sBXP07DOoXA3kA
Ofr5hE+teekvj0G6ipSI0RkMTmrPGG4YtSUu8kBNcXGWBkUIhQgR4y/ge2a+
JQ5HYyHBiGirjJH9SO+sPTqLEEo5aFDRvEfI3uaP5RtKmNut4qoF5X+VBanp
g+nHbErg70jkISq+dQvQ7nXUIBwmxwdhG6+KEBn5I56Wm/Q4FUEU7YYx4BgP
0m5eTjHkq23xkYx+41xRw/vqZnaBIucxhc7MCpmCzWt4sdsdvlldguI34N1s
oUHTxeLXkm9Pg1NuID9jlzrTywJV+NnYB+LViDSwUjtZ0mGIc1JUlZ+UqFjp
lJ6Chk+D2PqxkiayUqV9utQDBxQ/S4WPbymqfV8X8o9x/PEhqU+nfcjhSbI2
0GcXywLcU3Yp6IoJq7fVWlSM2TSW2Br3qMdAGPwz+5c436Glo9FGgTQzbwbO
P1gm6xcqXQSO1CvZIDKT5hMwMW0lBSn7bQg5EC798OkmM5HRUwiyWPo8Dnw9
PB62pPvuxMbLmwyUmeDlnZvbRP9+DR5Y1BBgHzWP/t15oZgLtcf8KyKZQPSt
aCzSaGH8CkGYUykRbtpdWXdXuO8Bw7Tj10qee57KG/WSqHxU+OQo2OnHBaFC
IakT6kaRTRkiTwGvwIdexjKwUEuPlPcOpXU6MdNmnRYszIvgq+qmexQGCZZ+
WIV8xtjfR4W4RtTtJksuHB7MhtXKPBhWOhdMjmvLLABDEKNMot8CWJwCIPeC
E2MuaLx/ecywXe75H7/Ak0ND4+HWdV4EesKvxiUjqpg7BR3lN036V72QRjh6
600lAKuNiM4MyB8t/Q95EOiG57lOc27zwroFqCu47J5miuVF4Xi5WHG6jTE3
3nDyCy9eHrnz5qB7mzvOXMUkLGI3U6Q6GX2td3SX0hIPQ3ZrXWVLQ4rCk1d3
8X2D7oCH9/PAW1pdpW2Z+qEHk0c3UEcXm3QnQhjVG9Ahm196vuEOBNI9dv2B
NpYeHLtZqlIS9JMIYJ7x/YoF6sVKc5yx4GBKEZZ5Y0I5aH8G6axz2TfsVkX1
xX3sMxAE7M0XmZkeN3cHgHCshXR9EssBl/pG9xXSG7nXVnvMOS6SBjv3D19w
9M+RRDo69A/tssqoiImGrfuc3LpsycaYxkX1DZvZJeNntL5Q4vl7Ld0KAE7b
yYCib6MNWKs5mbumvWsBrVRRABWjF11LyH+IXlVNSVHhLdoXvE7ZPo1f9NEx
0TvenD2VimPeRIra7W8v0CPkNn+NnaRwIFquoBVfWkgpZWWOa16oKQr/1Mbz
LoneSkUsclBtVCCI/LJHLe0kP9Mrlt4GxBOUsoDYwWi9hceUmf/cjtGEaBid
KH4dVprGIrN9+O8ntfxl76UHnP4ba2lsi70oMJQwsAvSgnfqp3MYbhgwy4v0
6nwcBpKebjMP6o/s0jTuxNVjBx2tQYiUZ1PrqC97bBZQPGnsdCw98U5b2tFt
snsTMvBIjjsACP0LMd1UAp1V1pVHAFE080ImOPmghqxN1W3gChYjwRZaO3Jl
EVaZLuMtrWTcPqYAfdYZWP1RbT2FeNquNvXyC0RnzAAX4efW971ap84f3fRC
PA327nAPThqUKi4tLmRbBaM1jjXH8saZP8SmlTrA4cN5N0cwRwDRIK8YTYlP
kk+YICdpB/t++95IaGLPP7mPRd/i8ZI2QACJjhfnpq3Fg2EfLeOeAzaFLykg
v4Kj4CHeYZ4nGiaFy1rnSJiT093g3cunhEWgHijIzLzr8T4oxksONOxwpE6I
g6/JkREdG2qPI/ikudSYUDoKJRB/u8LZrv014+QLIosiTXmjDbXAIrkLwRCR
D/O5ipB9qUgu4Se57/CXQcDkq3HmIICiOTgnw6f7hrT1PDg649OTUBPM4CjP
M1QR4Uw4hfThvxLLZg99TnWveZxQIjHJoRFvuL1NAGOKQTPkVqZqD0pKC452
9xrB35XoYupI/3mQpYozBFbJtfYlAnjrAHOowboLt/kFP82Rc4OJs9zYvZXK
R9rf3Hyi7hxe920BiUhpvkh9BVWSakjUEdyBDXk7D2FVlU+/H0l6AUtVNyA+
06q0HBP5yDplJqfY/yMDlsd+lzqA/ILQ1tOxWrAEfmbOn3lmX+YbSJqWgoUL
5sJHf9Ktn0Nxf2oIPAdl+MTDtcQbbryGpxfFxxmh/85MREYeaFFof/O1b/q7
oHtl1wXUDsBm6vLSiRAI+8ZkLlr8qiBX2bLnh99E8tKH8GTp5G0kIfa9RgdJ
yePXSj/SpTqul9PcGwLf3WEqb5/B4N6aYuvk9y61BvXJ+wtKzCk4HI782qvv
n1OJ+8eOf+N0VVAClsVPcxvA2JRxUp8UmPthaq+5uqgq3YfD14afUsmXjLTS
RwoP0QkwcW6pMB59LZgBXiX00hz1V8990FxtbfgAq7Ou3CmsPD445at+OqWo
Ly9cPsTq1M4uAHFRw43dWi2oy/kvA3bG0MF0QC+z12SWkCsxZPGUVVfKF4YZ
myE0lAE6aUvA7/PtDkoUj6wmiriGf07BL5w3+s1KYn3n/vZ9bm2Y9UAHK7pq
NM3jKBeedUgMnyG/7EYFqTWcN8/OPhmmjZUnpIf6csztpIqEsMm5uVX7hjrr
zxzDGNcEk/Tl+cbxT89X5qRBLZvIvXJvlRlQbEFcYMCvWwGLI9/xns+JPV7F
Wf6NP407ylCESf6U1KkPI4h+yNIZBTNQi6UtMyyrjsjHTYlOpQ3Jauf9g6FM
l9eCtMv0QzhDFNk0pG7GdCMxVcKlyltFSS+iTmx72Qi3bDr2rsE/PVPH7BdB
leQ9JCEOAu5G/8ga2hRteG4wFBmgXenBJCWHuZdHvUe5TK4E626Ca0a7JxTV
L+agsCeSQWvjYzPw6KyTbfm9qNRUb/HZSnA6fX4rU+0b/fJVJGPLljymysLS
YzMphY/ifeA1s/N+LdmzvPuFzb6Ez1EfN+Viu5e/vq6jFMm1yEl8WSHaaezF
wrjlfzo+QdOSKDTcDSPWmapTuvSNqnXPnYfmXp5tXYHN9yHMRgWmuMa5t4to
zj6xGLnwVKgci2rIZJlzU6c2vV075IXMBFLaLw+ScnnpM/zvYWQEa8m6GHN2
bMXnKxUeavZs9WWS5DrWl1ejhhgI/FczCoi8NEpxnOtA+IOxLa/QW85Z++rk
1wVcidr/fNW3R+H1k70L34rfX+XKGBa4/NvjBYq36o/Dz/tEU6M16vAu1Vm4
7Z1T8p01Nrhe+mLO08Tk6cgZvL9Fam/tvF49fCKzL3sgk/kBS+k9dSro4ad+
bTF8BxWjdVqeSFGbwWlA4ZhxzFyKAa7+i4k2ZWaqTTaJNS0QKSsIe9MBQCrf
KzhC+frRGNuOMDtmkAI4iNiVV3Nu1MbNGW8wT0ArIjLMnUSNOA5EBkl0Khwp
Cky0j1vZ/CNBbB7wAIfY1HwDSNmepr5Nw/NPgzoQ0QhDhJekncXGLNK5mTox
N8oWGlc2rRpF1pjYtyJWdhDP8ZlC6aTxOcGlEs+ZReQwePbbVNQX2zhORQSy
BuLH6kTpy9gToVYKcsLRTsMF7QnqY27faxrMhzeZpmRk1Qxi8Gl+blwtEoSW
OuFXQ2R1m1spGUh5ZzM5gH0yJuh1uoFiiNVFcVUybKPq1kwVicy3jAeLT4ic
NLQirzzPXpAbYRRVisU2JrEQqt3JDVh+m5WDvccZ0BCOhCT6WnftGUMBky5M
Ffl8zwpbK6OSaTWEHwr6t+3zJUptHxJcMZdgwuPOaMHjcUDNbwYu3bznpI1Y
KTPdCjpg40aGMmW0VkEf+6SkJTCoPe38/+hKFINi2Cw4CIcnKmHGU1W4ZRVU
eFRrUhOqOgQhXFyXPXUwGn5zOWmJz+ZW2iOPrn2O/dVN+JW+vs0Qw64FaTp9
/3DRJ+wNtTUice2KJiQRkYI98RHavAr2rr1pnFIgDzAmZeZtEL0NtFoL194b
aiBzUMhIRALpU5G++AtSDaF0vx/6Cfd7dWyFzNrD4CF68hn9NxuSTn95JKdx
kI7r7GECtrFCVyIajWMXes5tsmZ4hfqabAG3WoaZc1o3a+qmyMLzadEBxMuc
2H0zY2TDMBWQxf7cZqu/3m8NS2j3Byh7wkvN68yjTu6cSaAkrudfR2aVQ7cU
bYEnHG3gaL08jBd0zAgm5PEHaq3VBZOmwRTyv9f8Y1RepYVDsMs7ty+YzHS7
eAd987CkdvQuDzG+1MeP0QgV3RqsuEAewnDbmkf7slRnR7Prfu2WJ404UbGv
mLyqb7Gqag/Rb5G1Bouoto3559sSfWyGjx6Y6/YXWGSAvZXZ69mpQFh6iujy
NsewC6gMuH8d/cEjOKC/BkvIJLwRuy8dyi078S54wfTQXPYtYBYqQRfk4JE9
In35WnNvTRBE+7djiPcrUkFuuYV4IcFItZv5s3KFtLn5XNHX1Ij7j1DxtBSP
sUOjHSzVs3tglJEWYk1uK2EN9ub0p9+0JUCGo4am4BsrNJPYy2Kfh/QIOb3p
Ei/hUFN/O65cazjLJ/UDL4PZVMhcZSSg3wTmhVN6U66lglsAX7MxW7i1BGYZ
m7botzUOaMvYKGhjMMx27HHMzcSUFSJAP6C3nkfBsTQzaznF7am8T4Pg1vqx
Oe63DDLj+hEvidv3xTs02UFDEghrjeAzodm5u6RSAicf4NjJ5l+tuNd6uP1e
yRC4KaxIrZ0sx9gzM3se123aRzon0BQlxqgAjQOC8Lmu1pDl0EVfO6ptWpIE
oFzp5YxAF2WLrxEeyMH34h5RHhec4/iiLs68/VMv2jWj/CjiD9bn5V2qb4+t
YD87eH6s4UAWLW05VtLYptzjGKG1pY3c/buy8ZCB8TiAPu/41AEs6ltkk+Tt
Mgn6r4Mxva7ohX/ix/i+cF+yaFBvS0IQTCLwpU7v4TEp9VVx8Lz20dvfl9Tx
D007yetfJWQcpnUQT5+x/fhGAwmT29jSNc/FGOZ7i4jqCrOs6Ng7v8r7VA1t
mIG45qgiD7lUXFojOI2f4TpVyzzKr8Erk1xnLpkvd8n506mIR6pQX4Rt24Ci
fA9b4SXVXzRPC9jcSYhDQmnCkQ38whYWWsBuLddf39hNEDrUFhj3EFR4F8Gs
kEvIn3arZXJz2lBiEOHBmOW+GixylciAXQOTMIjDMwhVp0ULqecey4aXM3h3
9K/BB6c4jjGsaZBU2pMin6p5hTcx305ZRfZlsSb7eOTdnikVly5fO5KredBV
mNVoZX0Q2yUN8EwIT/5xRrymyUMdqBVQoUQCSxROfv+UjfnMLRaZEnZGBE2j
a8V72oyBznYIdc3LgSMW8q1Ry3Zrwd3Z0baVNcE9bv2CqXs/09cJsh51bV/O
vhpXic2w5XlH48wioZ2i9kKF7ppRitBHaRyuXS9AtO5LcFXrVA0tN4blIIvG
EyMOrvfb6cCP55lvdRUYvYtsnovnGNXYKwG01GgVWpRM+bbhSwuSSbbU1CSa
bfz5aewMlHQ75KYpjgGTo/Rmkx8Eos32jsxzJmbrQyzPEkH05CPdXi9n7sau
pC0z1PyI85j33Kyxjl24UkU2vcYZpnG8oZuUjrJrdQWzbBBdBOeojCejIEsL
ayZ1pteN+i2Sr6wkyfjTdE9cyQOGo2W2+z6Cys95DYB3iEoqBfYitf6+pLhB
32x0fmoW1lfJT9Jj7JPwsbds3Ixb9uMzHabVB5QxvL2V/j5LRnSzf5pOsTbS
ObhNpUgFh+kW1GcyiVTCI9Hv0ZMwKEEdAR4qvn+qSqSKdf49kOACeUGUmcgc
Bf9izXb9DKN5hwUFdDeFghAuisZSrHKIcQWsp1NtJ5kWrRgMOsGk1F9GbVBf
3WjQiYX43oKMy/XH1f2k/P359ITZHU1C5e7ugThedlG3I+KRwmITKtxnEDRs
OV6QDWpSvuyecEjNovcLRpVuU26zMTr3IzfNYJgDViDyGEx5TSsPKqKU5ANU
6NOwx85d5hmfnRAvIKIzLxBCucjGKvFdvPs6Zn18jXirUMz67DOJ9B3ZhlSw
EQh4g2uqxvHAMLMQmXIkC5MmNfk+Tbc96J58CLTDRpTjW8Pj+tQ6yv3QaAv/
ovXC05f2wYq6b8+ns+fQW+40nLW/x4RnLY/L74J8J6uuMWFhcrYfO/BAtStM
q6rBKYaRqJZczIVsuubj2LxFCzj4/zSRF6ibgqvlf15hPhfOB8UeSlSngw7Y
7CA1dgt/TBA5AMMl+T7b1oTT9+mop4TvAtwgigCRgeI57HGGM9/yMz7+9B+U
Ojq+j1QBNhPlvbUtg0FFBZKYDkuql3Iwmm39nTHl+GRuHrEHGEl+mhnZW9R7
ZP93e5PJdeHsG1VdVo3XKa8cGhF5VuOOqeNWuU2dRyeQTbjUmP/Zv3pWQq3P
5UyIuzz9TQOGkCAVwFY69+54AU2Ku8nVhO7nM0lA1N13+L+YrAaadfgSL1Vk
f24xEtcAazzJ/H/4n3FO2HUr22eFyp0wI0AhMh9NxAELQugdq7bdh6yUUM+4
iT8Rq/cbmkTkICik1IQLQpiI4wIwCXVXRwzFrjGO+OADpgwPOimyRvuDNIVe
QP5GD7xK1HZQrWiJkDS0IVzF/K80NareUMz6dGFKZs0tWzS8EL4QCWM3HK8/
OTANi/zexuEqqbWGxWuv298CSSg+e9+2J/RpzPH/eHlhfJ+7UFWHaNXS3QpV
Sg9piBIbTyWi2sDgvx3sZXeGlfrcbLxswYxQpcrNWNtDLDToSzt88QwIEqhr
jm5OkgmwvljX6J0EItg0UXzlsy+20VNGKF9+L74O8JdLx/SiQ7yc+tXqxMmO
Haykhe32lGxe540D5EweRdB6KMhTezxO4r2PME+M66HgnJrKxz3Kn1H6PkUR
1bAKWKx0abHobpkTOlWp3+jOBgiwhZDfcE7BAPTzzdy5WHpn55gZVKEEtLtX
doMYalQkUnDBqjhW3WVlgwj3bNtWbqS0dO7AA0R+e7Y2dnT0FnzS28oYWUw6
YqxG0mppgF/JDiVtexyGVrAYaVVJ/5txWo2wvHO05Kxuh3kUkk/qK87AZyCL
QgRH4PncDCVaYolyFo1/2tC+uUFHleJHcwQDe+hfnOONSbbYca/JLRLCyJf3
G0tsMOap2ml7w9Wx4G4Rjq09DhZZdbDJtxxbMZfXqEcqe4YBwlLLpVkjhaRD
GhO6q4b12mmQGG95DNl1JDTacG5Vqoz+Y8cDQ9DYJTF/MXxloLl7twD1wvew
7BhHgX2BkNssYSSEdQk4u8WcOKZdbompCPJ3OzTDuqKrq427TK2ARezgxdAR
sqWVEAgHMSQ5AUGT+CnWqDa78zajvdkVY6vlxHUq06Cdcx5O01DcEjGlUbTU
C0GxuQc8Av/IBJ4nIfYa/+iTcYMquyp4Loy4ZpdJuKz4cei53wdg/aWbk9Xt
BFw7QtWVrEf+VvZ+LnXXqPP+3Acpndv27mzQ8RrY8jpoIhoeeK47BVWFlkBS
00NigQwXDsohwqQe/wf9XJInHhHqTOmmRg333dHh0Ob1BOvtKXmcmtEcqGk+
hsW7C7MKQz02kn1Xbti3NXphRCXHGPre1j4vgeugdgwsIity1YcFdeJNZGmE
j3Ozoy3S2q75XACEVvhZEbm4Lh5H2wqfknGjqhsJlEoU/fChpS9+rWoJtvaK
4lnk7Cqh38Tao1ttBVnY8Bmhfd02QfzUMm4DClY8vTv4wUTvuLwJ1y9XnxDz
ItqJUbyHgz21TpU+Zmc3JWo5PoSWEWg/fdECpOctUOru5W4e6DRMb7tMxTev
ue4+h68MzBWjQwuW09yR5XqgWJUxPsxWAHPmr5fVKs0NNA79GxKB4YSAp0d7
ivSWF0Aepu6MFqWq65Uusv4sMbU/Lb2djT9rsQL3MZDIKQVSUdITHo4PfylV
oaokZkeh24lfzkqg1g1rQgfSls9P0I9q4qg73apgJcnT2YaVUb4BQKjD8lQK
a/Gvj/Xb5VIqk+7D55/ZtHndsEtejD5RXYouRnZ2DMJDZxCekc7GNgkoWwvr
8nbcBmFI/3REygOY57yD25ZId6JNcM+9moe0eMGaYdB0E0rb1ywS0UlsiBrL
3XhjgBK6tt5nGev27bj/j0RQ5yM8+UzrTkIG7YAqyR5yK3VwMIboquCfKUQ2
z7noJ52bMD2DZKKY6Eon9qjbxbaERtW2ixApgeSibo+iZwsrr3OG/kWTt3nG
NGWMcpZAMolE4TEc+Iaip/DOfD3nIDiogrDEN5e1i8CJb0k/x+SyeD3HbSwa
cfEyH5y7kwaELmOZtuE12zi4LlNnJwG4SZe/gE/akyjvODj9U5hN1XiDZ/nf
AHuMl/kP4SFyaGiVUzzadcoiJP9ljOwrZvH8UrhIleOAagyCkzfLQ79qEd1p
6s87p5wVeDTZba2n8/0iGCHi2fh6ZbQBqHsECpy2GceOcas3wH9B5JIFyCkF
UdcDfxSO96B62jLpTZSNINVKla6vlWT7X+FeIOJai/fV8G+Ts54E+L4Hcbnn
KjcfSJZtDjH4RYUrRKhVtkNvsvX/p+vh/d+rPFKU0SxZXpz4u3QwyfjnY2gP
ai2X4r/hGoLWUIxjxxp/F5knsAKi0ynpEq72MQscAZ8Yw7kLteVKuwFebhTb
R6fkdiwGhLQzSQW4Im/okd5ST08ZOW40SxF7430t9ymy8er10uJafqZsyLXr
eIIz4RO9KfTIGNOIgXZj1pzgubVJnKglWR9CNfSUakg3QEiqTrIAg0kvi6V3
MgJN+s971hLnAjSExj5KcNDQHROtJjpHHirrYa3GvN6aBILgwuRP7vJDJvuW
uQYV+MJrQhrpDCCO0jD1mDKpy0zJ20xnvorVKUbnM8Vn+B0Z05d5OHe5tdQE
kvTgJJ7PXdNTakWksVpGwtxnh7a/p82MA1U6APTluKH7N6SvKgyr3AdIiYre
w3iqaTs3LYIz7CsSuEUbjOiooJpPsi9SeA5fup36vY318mXhUsObqcDe2ndm
aBXOEX34tfHFDe54b9ZNxEu1nwpKatUTE0gXG6kiNBUwv7U1t7PqO0O3gkW8
7vdbYHgdyDWY0vyJVVKUxuEZsDN+uqGmmWGqzBFmx9dtZRFl/Y2w8vISU7pg
oO0WtAqKcxqqpQYy+z0qnmnffAF9VOFfJs+gs7lFIiN1lkfLID3Azx4UamSh
2ndHVW+FLV2mg5dbgAgjHmk0ZU+JbdkaHB6cTX+XF5eOBEpLmm1HxMZFisq+
l1O3Rd37cEhjYxJYWK7MMxxWG9Pvaziwbe1X6zmQFUCRhDLLKOwXAfTl6l7c
nohxnCXo1LCtO4mO1hEeEzKvRCCGhzQbtjLM1SfaWopzkyzTEOgB/Plp3Il5
Bjr+gB0hsNwF49DsK1RM7PhVhm/1AEQughJa2g/ePXERo6hH4lDZbfLr6Ib6
zhUwz7T2fXTzMeLm5udLL6zcSjw/uwa66SS0NfmvOWvinLGnkTax7cAKnRh4
XUi5sSxwsj7+iJh1f/Y2dX71praTmngH5iY8Ndro/MoysIsXErx4fCeFTx+r
zIu7qMiS91ixlNHBRgBDAeuMui+Y2WXyMKwEdoMMbCod0evvqMC5BQLdNVE4
pXF1Ia0aLvxLfTdnLziitGM+mL5h9JMQ+0NSxi6ueMaA9EATazkvfDjuQTYv
9q1FtxCE8R/p0KvvgDnya6P3uKiF19B2x3EFjGpIE1cx7ccWLl6kh5vU/cmZ
VELFo48jpgnfoIcWWpW2pun70fqQaBvAs08OLgqHm7pukZquOIhOoiYLTW2t
nGOvZyCIHm2Vmr41ENFfw1bP9nCcPMYRmwOhPZgvJu3Nm6K84LTBLnbqK+9z
zCcFrewbHWX//HktLnnw4UFdNc6rmWsAlP6SA7FfWvHEteOu/zkQod6Q4IOq
Yq3EhRlUKghrzvWIQ0fUxxsbBrhIatUtS8NYazej183aVldq05iAIJk6JbAD
5qK0QgNnrFdljIlQPjeBQ1Celxhsv/kcgTw8xquYRLtHQUXdGKKSYP6wk47H
+44rj08jPdo9Gz/lp98ShAq8Q6MIKOClv/ZgRwVB26ORgrmhO8prttj8urJ2
37icpIbLdRUK8WlWtq2EHGPRnZSHvQHaA3G5IqdrOWWfLTqDJbrtLfDK+Czg
BdsnEIMMca+ygKn4GcqAL9rI/ZeRsiHTE9Ws63qz238W0fM71U/GApDkHl2u
dfn0HikN8hgmWCmOIuaFeeJqT5ehrZzmKpKU52iIUpW4noN/bIbCC+U4x+U9
sOh7xMobDSSIjam1+M+O8lLAdFJKhzUibmKMZyc42mMw+muys9bcMCuBkUQx
3ffHKUgN+6Er1xm7KZ7/cYtFm+UGXytl762evIPIBt0JmtZJ/0/jv8Ni8JV+
5KuOh72AH9A+zgReb24ggr6Ku55ubn8p4wupojXvsrOEKsLXLZqUZm6/IAjX
lx/cgtC7zmYdzwD+MXlPlPz/6vQ+ISy9zy9i5O6Yv+TKILWeCMQBAqNibooR
rPw16epBBLKUuboVV72PnBfZ2mllQzlgO+2QBSgjIjvs+E3KLX0aw1rqoP7v
UOWkjJnLe9m5O7/1/xjqg7bICJE9AwpAjhKKjDNRiS6mwMDzk4hyEdXwYzg5
Qtqz4juhHQZhRex8LyRnekn2pfv3dHPeB531juRQzTY61Hc2pHR2zqTMGJHo
I2yPld3Ksk5x76Lt6s8VuAEXobQVB6VO6ewCTK01plUZUCCwPL++nENZqTJB
zNqo0yoQqQ0ATxkGA/lONqQXTv95oXAVHnQcRn4PX7vtuEnLd4S7ZzWrphLN
yHxiKyO8ucA/YGKZ2XQWQZ/E86ZfW+UOfLQuxd06AeRAlvbZ2+hM3BZRiGQT
EeSvRLfJv9oxNspZQbAdNZg4oKf+6rHQZ5DwE0YSbjjPNWRfpJMY4Oe2Jd4f
KMFfjSlAw+B4vnUnK1p4aT9tKINk1OLhH+pQgLS3Hygkj7gpq6pLEK6u7Gdj
m2bTkrWL9dxNE1Y5nHgh/pR3+o02Ctnu5fgLPyvl8Vb251EQ20eipS3aLuMh
flCrnLuT/AfGZ2Z6dFuOyT6tfdKaa3+8GWrHTNe/txjqMdy/58ItibFBoouP
G2WreX6GRCAPtY/0URnk7cg4fVb9hxvKKP3bV55AWY/gBRykZB6J0B3cLVkh
uDGFhbDkxlBItjNTcxcuUbljqsClmCBo8C7IPO9RcT9W4pt7q4D9I0p4JWAw
M3R6je2SI0MV58bG3pXDDeFcFa9aS37L4lGfkp4L7mT6YJRxg4B/oAWpNXQ2
cqybZ0lBLej+gfPxfwWjRed+HyWYqwCyQ7gU+X8/YUD+rNCCBWOX3hoU5haI
QDPeb5VLepXIzzExgKJObWvG7jYK4TUQa0J6QxYRkEXNL/zHU+qwaSGT/GGE
znaou0Wmaf3IzgB2P05fd4BRmN7oG7NQ8FrH05qRiyCNgWcbl1YBKkiE4t22
uulgQXZMvFPhb4QLcnuCC9L1qCSZRq/2HtvE5gnua1fryh/XJtSrlwLMVHkZ
9+U4THN9w7aYTB3i1rwKQ9WPxMqJPjR9CaGMbc+vNhIJT4dMSfZ+NdVanF4H
tgDuHkBrzbgNwFSOEznwyxWiZ8BtSg7Tl/V1n400+NZMa2iAiakEz+jHJ/YA
eAXZoTCc3TVRn1vARX2diG8nf6y8Oa6ssM7QnZCm/vl8nEO3eHYRWzCFgH1d
Dlr8NBNDHY/lge6OK3DHNtje3gd1JMbd09GzLYfpM4CykBUMviaWrYU/gzM1
9fOC6TbCRHQp+ldbscETkhMANMQB3ooUKy+4Ea1nOVWOmYUPhQfaGcgIQnbp
LfZJuQxV3JlyUPJ/275rHNcpVgMmQF3KEgEffvNiOh/301DrbzcJ9G7Pozx4
2rAZVI6Fu1VXRlHKmPOL98BsuGZrQqq1H+PcoXi5vvvdE60hTt6aqUAE90yN
oHN3NekOXbcxXzmZK8v3ae0W/W7KoKb5kl4YNWeL944EdDbw4brKaSz/Tuo1
jyNuBf7FKyF8d09jp81LQ6MfhyWx0LtUWv6l+5psCbrJJYKrACsKNXxAsh7o
rk9vIfPiYomMeiwy1z+mEnBpw5Ko5OdpwGb+UQFZqKk9YC16sR5AHnWh4E2P
EyZP2F6wTdV72ShmEn6YBdTsDGf7vGHxdocx51GOABKQfYMh88aOZGo38zFN
fmwoxi3bz2iemJm9hI/6vh3okvErGbEr+VC5GRxehlRIyMBJYg9iyFSWiSMP
h0Lsv5Cu8f7AdQWujMzNyDdKFaEGQh2vq+hbLG4ggFnxnvCtqXG+x8n4ETOQ
G7RWn1Ok12E3u9pGxZvVzQPmjcdbxjWyzzHWTz4xuOR8jTGODMt8n3pXiHb3
5Y2xh3q9AMHb74ApG1sqFYbt5mkCEuBSCxXOQECv8SRYt8BgNa5HiKgTzizJ
HgVzk6YniPitmO8uRMDqCJ1FJ4/A6ZWFSsTCMNjcP5LL/7LVoa5+KSwxDao6
5UxNSqNZKJ59dPN+kr7W6KFO7a2HsQcQni9iPBtYXHNoyhbzI4t6U8E1Gb1M
A7ZhpdfZ12UQCLxhKfbWY7LId+mdgXQ7AG9pUEKy/kahI5beZUn9CZ06THcv
Jwa/ProZ2HOguNhqFRFuRH1j5tgYNnWnGAgRiBx3ltzCC9Ercdxr3FhaqvSC
EnKk42or0HNa5S3LbfNkDgf9aBLNDhJPghkvJaZ3XBgrU11mgwDqGR2zu7Vr
nwCAYtlLtnwnULNU3vJG4huwtzLZ4IbBGqAJtPLs1tdN8k/VA6vxUuv4K939
sK1wI4DdMMaQ43FeaQotmmoUamgwo4IWUzj/nCfTqkOiIFSAebWrJX02eprF
u31Q4xPvU5+kxGDUZOxha7zAODT9BWJuPlk07GodWBkU6D0baxBnZ5E3WpSq
n7931utmPoui5h7iJU50hH7sxeHKepD8KRU2sYg1BaBoygMimN7w4AWWmmvh
Bw/ZEG0POcpZe4F2yuqOnPYZbfaBcw6EsEaNQvJKNGILfOJ4CC16dPvnIC+s
jfOU5XboO3bWV1KaYLOcTYO6dF6iq/vwpWSGOXbVCwDWVW53HGE0wBfABbvN
ZPD73CAS6rNsyd9RFH67tyRR7PDjQy/AvnXDBe/OE3dJ9nqc8QKL05VvgQMU
6V/g/oI/io0mBryD7rvXfvFLFnq+aXpUFd0RtRWRbSZfKctb8EVaMvp53YaA
ZyJDLaULDVOQap0Vt3n/NFJMn1cuOM5WsX8nT8tyUhhR5T/d/z6LUExZUbTk
Uz43hhqEz3MUvD4MRsqzXCPAmZKEHhslio0j8zkzqhWKEA4H+lDK6Kc64wE7
d854nha8h1wxpq+60nvHNNeVAcQ9IYnyEcdoZCFDpp4jbHIP1YfoY2kZwAjy
CbobZ+AGQkr7XCGqBRFVSRCWN7RWJUfqGE7l7f8rl/ZDVBvUF0jDqwACPXaj
xuJhTyuGi/mKy2p3LD86EOlMWKgxTa+dH0t/4e4okecXglWEzF7gSwYiJ7Yw
cVemQKuq25//t1Il8jff8NIviBlop6yV7Na3EZPuIyMK4eWVTuRprtCJS8Ob
2wP+N77iYnG92ukxBgrqk+qdEJnXgkiDBIERVFvmpUsWQqLth4kIKDwelbEk
F+C1pgfzHlVhDpBB04BdNySk3UNMf90NtPaCrgaqn9qObsGKSmVl0Wr0Qykp
6X3udFpKemcnTURIyqpxu1nUpYJARgoOkPOKn6UdlEz6sFAVU785z97xwJTV
tSEnJZBNbHRUt6jeLuJJ62hcOVpxdgKInPgRote03yxt4/Plk9mGXaPxTncw
RwYnYR4rU8Vu2wUEcO7Hr/QBLvJMsFWKUU7XsBb+CvbNspyCjX18bzlpQzIQ
vTQNvuwORiQPWAPk8rq79xAOGRSw8Chp41aFdfk9xo+OufSCda1YLL/UEKZn
e2iZ+ayj6Hn8mBsFZvGY9wCLVmn2qTkIvpF6kxDpGjUfZr2y/38sbcIlny+H
1P3bKgCztcD77bxImLiDOa3XxvXk/o8S1xNTR7g0yaklL7cDk4LbMlNSF69n
c8IM4ZE7XEpwKR//IYBKWFVSCXRGXsGlUBRYMZX63MDJSzEKbVZp+HEhPnb7
0umVISDz69KtLmtE4MFTkm7AA0eFRejlCeUcwi3xyTcmUp/emCvhf7Ux5rlg
tt8W5cxjSw5vveEUTtAvxKLCoXYJIynFB346UIIwNwhfVGRISS4Y7GT5p3i3
umlnWdd+sO64oIALhHmpEhKogotGdWZIXTzi+/Y53YxLe2gGD/D36DRI+fU4
27ZAMzTJM/pPtnzDGN8LJP02Ym5bJE9+8w8NKTipMJZxv6ByWgyXnI/QVyeU
XBCPp/4zmEpNMc5W1t1ixyqrCwuU04BQw/eBRan93dnzsd2I71XQR4jRT0lf
ziEuvTPpYCiHUnHBAGLOKxZT2XU31khcSMSVjAQcTyQqCorIUiOwg6EzK/bG
9r5YImBgCLT3XtZtuyTmK/DGi7ARRP/wMBx+lnt71kZdwgeYo3NWwH2bhXoi
Lr5Ir9YYHll9eTMbH94KsibdMOQl16C4miQc4WrcvNMPpDdOzwHRWXlv1Eko
AWp5peMJ2azjyA9VBU5Tzz8b1caqOvXlKjV1He17BYDXKdmsKXOeRirK8H7d
rPT/oef0VxLebU1pAxFFOCGXlwnGFCowxCoUH0NiV/LjWBF2UPWBwtLjW0ae
mw+eaw2D8f3QkrQSI8GzHeS87fg1azD//O9Cz7P7kUjB+VpcYymxlPiEoBIf
tmPgcD1+bs0H7t1MsMuUjefPpwAFrN4ylNMr3t4FwZqWCa/L5RVD7A+aEdFX
BVB97/jzSDwyviiQODIZky93WcV43BQiZh829rUOKl3eRd22SE1URLX1F5We
mlLADj8N81gxpdfbI16a/E+JTgNoAPLf9h0MY0rTq5sjvUi5h0uzHilGyQsy
TVKMrgsEko9l4Pj/m1XZbHy6oROUkYy3Fbd1DL/n5HNJCHQ/X2dEJCmPHZ/n
fMv+nU6laR0Zhr0OI3TEC/Vy/KrgzHZtqyNSiSfMNMsBPtKJfNU37GRjOWMY
bIGVJf9BNHWmPCpcRti7CEtjndHi7J381gYCF0NNMPK8R99AlmiQfEW9v+qL
OsHV8c9/MxWBDGXQJ29SEp08zQ+upD/bpWju0bt9Nqf3HP2nEMgCjFudyt6r
yflUSx3yEKgopzFCPNYHvTM+EjzgYs/I7WYPQANKVMm8ub9VrmnnZ1lHnVgB
/sdBRLKGRe3rBbWdWdDRgx33Bu0h03YcCVnq8fq/ASQ7k5FA5xLHwkhQR/py
OvUJvjE9k3lox6RGVK7W+XQfPRo15qIxlqZE9WeM2Y3KZv9WHYiosRKLgHHC
4oKSPF0oPx8nyqePwBaEVoF6Pf1Fat7UW0UGtiWk81f1jUCuyQMpdRVLs2XW
G2ZK5lCdUgXwyxQuJnbEMhyrBKtzCONQoXhzfTyoa0J8uHYMB2ZU5EzY/UzK
z2sRp3lk1b6aTBko+AABhDwSYHjrFZWZVbB32yfjpZC99tFp/IlM/m4Os6Tb
fXfSfTrWsgjO0vkqHXT7o3ZTJ11rZzxQ5KKf/YsIxmqt/SMU5TmuXY5IZSFS
4JpqTx4mKC0tjrGfABHjOCj15IYtQ5OszLUb7hCOZFx349Ept8T49sstCKNN
RRIyU5BfjsrvLvSxy1N78tAvf9aMl0F6lLs4kiJCYov4YzJMPG6wz7/fAWNI
qVvcpIFKbQdBp54YkNkyCcJZPmfAlIa9kCo/AjarYM0gNlKkOOy5hlWulAc9
ieOY1MG5X4WHOlH3w9TLQc4QIJz8/VaWfJzAqFnDQyOF5W8J2YfxrlYgfJ9i
oplblyuCyhEp/bK1+GzurVHO76QV5Gd0aaeNzz5OsmjooUsS/yZ/PysOL8I9
WdRDKY1gKLiDrB90YYRwnKMjU8nPOv09YoNNV+H5oTsZk5YAI1Sl9kOaPJEt
B0YPyh93ze1fIQ8PVJ03ECB7YR8w+MAM2rzV4JiWMxBlnoJGv7qVypvz61GL
iggThL9VGgd8CcXnFp50/hNd2aQRG4lwLg5S83Av5IzJNFar95dkcHM0cNC6
TOPT8E4QA6jEhmRc8rUBlWhdO2CQ1dU8FPnnrMkc0lcOlxLOFkQA8cobO1NR
42+wbuDKmJ+fqwbIt5YoKfuXiwMY7Wr0+lxzRN0gF2g8uYVaVFl9vTnGPHxn
zkH8j420e7/jIiU/tunFcNhTEeZyoIFkuvdL2xLpbWgVUVM8oiLIxFWDRy5r
jVnYUse4hHJLT7I3eBeTPFfb9hdoUPmpJ6Fsa/rQp3M4NL/whSquqR2HBoj7
cMUBqIMScbS5rnexIG5FGKqr2HQwml1v9CrzYg51v6zy7sLzQk9VguObh7Q/
ERDGC+llZ8bHRYVXIEnwW85vOBnCadiqrqr57xEcPMLl06+OPSpXnxvQy+Fg
30Zla2907Pcj+9d1xrnoVh51ves3H6XjP92KtQorn6mK5M+SWhK1WFvKJ7BB
F1yT3N6/VIc4q5q/+FJw264OZdDCH23KZi5XYRbC0+5QWHSxBsqRQ6AFajD5
k6Q+im8vf7Wie4ytzJgjLdG6gDH4FlhCEJLV8QhVZcfM0tXBNPrlZFjPxTRh
p3Vx0AbZEc34iLf3/s3Ir+qqlM5NBq8HsQ2bz1Q4Cm6OYnZuJudVGBOJSINX
Q4wHONmwGt3Z7waVBvriIO2D7ZGFhOheLsucwKlwG/d4j83484DVu47Dcx2k
oOMuvyZxcqj5qk/YbAhx8+6enclAE4ateGFRfZ+Ts3+p+m3XwOxBQk4gAlNG
YXkKx0vb/D8N29TZ/QUcA26DTmOQLr7k3YBKnXCM7ph/D57J3AZNzr7TjaVe
1CL+n30HqYsktxcpjZuabHtUHT6l7TtNxRJaE0+9M5SRpYAhYaEgmVYKpyqs
VJrZCAUgc2wvRBEM6wRVu469MM/pfZW5YiAB05cL4Z4A1xagzNS09cVHyiDd
8ouEYgvdzj6fghfg8jQY0WNYFKjXNOuXWOojFR8moj1x0O+m7SvvpMBCJ73C
4BLMeoWTzQzO9Y4psFyFwcCEwT+uKkLpTndV0autXOQSru9/KYTJuPAPqqHF
EV/soQQaIJfQD/4koUK48Iwx0m236unu1VPbHQ1zDGO78tO50Wgf0BL8qTDU
19oSOUG2vpI9Zno1YV+i+uYlPBA1cya9OHAIe+Efmr2c6z9/Qi7jORmx20S8
P04AI9agfA47cwypw9GI+/gq6CzbhqVNrVo3oyerp3yVr1nFdfSBxnT6HTqB
aM544bZF1O9Sb6Lj/fYC7V6c77B4Iak9uWXMmEgQdlXVMbzzwh1W4ka2IuX7
GGs22e5sUE6/xHuCN+R9txAwtPmq5iuN/M5/PcUooZ2HIsX4pM4Ay+my+N17
Rj3fTo6QFbx+x2HXG9KX1uPZG3Qbq/Va+XUgf8FygRIjDwHm/WIAn7EuYCCm
Hh3+9475spUfl3XTb/gxeYhaaLQs2scfamm3HxqiihulWny9z1EwEMN2vxW5
YhClUokN1C6PDma7uY7v0iB2DOfmNYo6eNmdWbug9iiy/U5oenc0hYL1U6E+
wIM4tD/cC+u1godhi8DdGAHVTahREC8OxB7PM19ZYT+Xb3ThxFcp2QTCDR3B
ACZtHsvofI3OF9RrnPwdKBjXCcAZiIDOql9ltFDRqodjk7t9EKX6PDTBEsdw
28QkSh1e0breWHJU65IyRQUWQTYK8i/4JyvJmAZNVJS0fS8mL74+pL+C7wR+
jsxQgfghPMS7D+IzIB8wKIy5qyHss5G8RSWsHWZPh8KMQ2HJu8x7SxqIi+Va
NIhh52S2QEyK5tPYZ2zv0GqS3qxv/TAeCr7uwhYZUL+0MGJZYGhd7uTJNiZF
AiOKuuEH2YI+C8S9m6qLZqaUMbhSpWj2i+nJbvZTsGmjITslgih8yEZY3B+k
urqkHw99emd1UZTuvkn63rZwqA04Q9RsahXhVLH3RGnWgBts+w18HLwjUOTf
xLwOBiE3k4ukQv81UiUdn6x8BgP2QNnkYYuACnK57ZS9sxVEPm7Z/Ocj38ue
f5Mg2lVq+VIvkEgAbMQXs3NsbbLoyTyK1nhtbN2KI7YeL418HatFytcw64Mt
S3KBE1H1dEDmIELv2+TGU8ewq8D9cVo4A6frbrTTXOEw3UbKkljcsa/JRLhX
vyOkNxE7BEdivMYSd5fx2fEU1MeS5jMeRJ8paJRQ1dMFC7HtL7VWuKpJK/tM
HMcseLubkSmMd6mCki6A0yakfoV6iJBOTVWX6ac4YfxTN4zKFpTmX/tBBpG2
9daBtj/Yrvfo+DrD5j+txX1IfIq77PvinAPRG2lXCQIodBOtyfyzG63WQ5BA
TOqOEVkXxmfnRMQsK/6VeKmR7sV7KoRiBj/rJOZDTVPB8SJqcrwZTULJlKtC
UUffQ8vhYyaASzbvPo9FMXw6k5XrhJn4OegCwhTNc/mANFIaHrVSrOs1Rji9
qX71ysWbDpiUEwVPcc/X+XGPoPkHx4JHiHBzcVhUCeS+QDYOv2AdC1Pm9LXS
He2Xh9anbCJELU2XA/PO1gxuxrurEnrRvV4vAIlGvACgJkncQxpEGbg45N6X
xrsiuxf+vBOEeHy9vyg59dBK4JYAm3kMxEPKX5kLk3F9y1eCqRMC7GT/m//7
9f0fwKVQ/aYTh3bubcxz04IsLca3hNHNFzCvJnF4OHXrKPLGNRaLaODZG6Cz
EA+zL/sX/m0+CWrs/JTSJSG/MxRyO5KJHC18KhOLm/wMtZslX9f//1lE5MlZ
iRuGnFDXcjGYE7heOUPkZJNZBCm9y0kth1eY7vtPEoEfHmdTy9R4Oa6poc7J
UOm4A/ZkC0kkoiIoCtsVT61eWZDK+TdARPve5iGQmqTi8E1V7a+2oUVQHDUz
cclsXEmd/PTdzkA6ufkoMYYjNPq4Bb9nsFRMSycZ/BP6uN/+UMtc8xDAQFGM
kx1b5Xa2jE/13eGWcDh2n70Vd8IYqf3Lwu3Hxr17cunNp/VVsmxKct/IiI1r
V67eHnCKEn3DugPqf2453i3sUvNT5v9AGt+wwYNvnrXAFmHuowrCHVmJCI0g
ZR4fWtuvLkcNA6CCYjegfmt4lYdjT8ibpR9dPjDkPTEZ4Xv29O0BdX/jdlau
hDBKaRNLN4OYo2d0oBg46Uaq93rsjMbSKpIGTMRZkIANwcNLxVU3sBfhnhKu
RLe9arKxSZIAixFFlZKfbChFnV9cTw9j8EMffMEmy7JTjeFJAGfdVMzmoPG+
5EwmcHLtG4P7lhZBgwEpHMT8BwESS6tG1nzxwULhjon1rd9vIyyxWWVGACKx
tGjd8F9530h78Bd5am24iIxdpAimzM32VZvTHlDslDgYa2BhUKbl8f+auztM
SECndocOBgkzewHv90Kz1Q6v6HW7CGXwQDoPFkWJ6HCEL/6sDXGHjHD9VQnZ
nuU0yv02tYtMkGB5mCBOKGLmZdIKP7j8tOmV1kguoYtrfEjkyWC+HVP/hDNf
2dBiHG5x8BBviAl8LjEzmFZaEB90EzMxTE0ivLmcfw8tOg+9mDuzyimxqXSg
dOsDBH0gFDKbMCc+VfhV9ZWyC5whrfzfWAeJBVXqHBYiBsZNGztrc0CUtu0E
AG8trknepCsJfoO+MxgRxXPIdB9cxKNF7Kp7lIoylsERs25DiBHoj7FG/5XU
5BBh6H8486bTwB0JVCRwrbOz55x6x5oPdH4iUQk/NjO8ZE0DCtg0M3oXwUln
bUKFkJTmYtru9tf2XqaEV+mw77XiJbvpGTrPqFXRt9aR4jcoO75/4aybWmgq
mUBOwxVJ+cccn/gzKgtRGBQWF0fAaFp3zsFft+MfCswcJ7duYvdpEZqQleiG
O6ALoVmDqWXJJUjffNkLuiuquHFba4xnE5Eqt+jv/CjLsOb6avbc/1MgQ2i9
ZastpY8iA3vsagP4r9Qzvipfk1BYr/FzFZyily19hqD18jrESUdIf7lnPF95
+0b5Tth4gxen9qLLPYOEwmvI27aiG9cXBRi0Su+BfSEZP/BNE7I11wGhJIEK
pysGYC/ykwHN3sdTBpEv+xS0qA0M9zLdxngZHS2hqDCBRYhctD7/FOBykMEE
CHj3/Nvsm7dnF/9uA9seMtm9b5qA6NvfUoCnUXW60oqrJJ8/yUM3TO9kRaeJ
nG2I9qh50b+skyQ3wFaQNAto27Ac8M4Ge1Kc9L530wvpyKzSERAAD1qTbG6y
xUCMtxKkci83+jEoWtxrkullsg8IfiHysN6L9xrbezN57VeTKC1+6vVyVjQH
tRbt3ve73Wso6hwRyCCOe979aowqq7qm8gktsEvScE0vwgXZoN2va6u18RMJ
Tbugky+i9weB1Gyop8nYHIPeHm9rZUuZIJUhVFQxseX+RVhkhWvbpkq3S+QJ
xC2ILj3gk7c7AnCN4QC7EBXfLSKzlyUXg8Bj6c8bOsqxcKSLSe4eM7z8Qqrr
lHtM22Bt9O8RBL+FiktS9rIFuR4hGKDGsauksiaeI0wS68Q+Ip8DhxbwSDrO
4FdQT9KHoCp5dDKSHaPD6PKP0Q9pwCDq8E5hqrThHwXGM90kojlC6Ru0JgN5
8kRxdm91vvcsff6VfvxMkKFHldBsWJBu8ykQezVaTcoWIeD5cjSclN/K9zfn
OVA564g2jMeVAyx9RPn5fdlNhaQB8ZxwZy0NVGtVSF0Jxxqnq77Uck7J94A8
N7j/PbUzix+xcUlMan+40YSR2BUNRbhxwlVUfp/OJU0ZCmNrp2NqOwrjVutd
M1cYIiOvzjZpqD8GKXSKv4+dmtIiiEEAlcEl4Khoi4EWA95fMmDCSlR9zm2z
HcNBk+pK2Hn0Z/8EMa5WThrOHe1dctdeUYBnWFzk/NC4IwOL37qNUBTBgfKZ
ft71R74MhDS1vIM+pbiRCkvTgyYhu0YPb/eJOP/jagZhk63+xJ8ke9Ye0uk0
YCPxuL5qs4KJM9/IKZWmckW9T1SI82mcqIZt1EbC2GLhJbK7TnbLyVEKcxj4
vBqPD4795llN9la0A5HvN4O9ajm6zanRpt2JXIJIRTZQvz+HMQJu5NpL+DZz
XE+7JDoVWgrOLoiNzTNGILDmS59Sf6mBzlT10ELV3gvkV+ITrUlmZoryyIlK
uKlC94YPMoUJMID1YHSHJ7uHexD0byr6t92BrMkFzRtGyetEosDZcM/13zJx
PKnp8YR7TCxj+zj07voa7W2xxCjm2wm7lxB6fySsuZ1g9Kcc8lNDiWIFW0nR
RHNvXJ0u/bSvSclRXSR1/bb2bPokCaCuIESLzlGl5A7/2qp4jP/9a0zNSYsK
Hg8JquYh598Qsp32DfeblaAmO2TnDmfK7pyewDarVfAL33l4GzTkBedDB3HR
wm2+LzjgYadt/fztQ83tb05QfTnLAEe87VPxRLM+zb+svVZwvgs/6tCFV1sg
AU3NkyOtq/zgN5APPRWywaBh/H2tKWOuhpKc3h43WIorIa/VbNfyrJRQUt2Y
flKTktp6w0+DYmyz9ucv7DMuNy+2ulVd14odSl3sgC1IsXyqLMaVdinKaRj1
6TSF/C3FjaKm0ZUT4GyIUaWx/H5E7skmQUp/Kq5Y2ne3ujRcabD964Fb9tY5
0hJhC+UQha3iF58yqLbc/x8udCQC1HOAB3V5dKE6LlfEOdv63EdojtEemLxV
FPVRcAmgXyYUfHLTKBLUdXsiIj0Ut9Xj5H2D4ijuuA/BEx2LCwvaU5DOZyz+
aBxWc2cixsoj61AnW8BTZNNTyf4LaLmnt8b4V6vZD0Lu8WMuuD6S3HXKagdf
hzgeBWIqWfkSdt4yllQ6yPTTRk40VfXu1mcw3NfiVlCcQyKRR57sk4iwln7G
bpe6ISZW1nfC2HXitjcOfqmXKvbRMWlggnwbFKfukCK+c1uS/K/dhSB0Vn6q
yifN7x1jpAPnCKIgYsH6TP/JFvfhe9scv+LGgxYKbPmE1N4ROBeuGUR0Swtp
OxqyV/VpJBetV7hE61d4TlZF7y/f2pnsmP5zRnOk7QJClZacuGYU/IBCdvgV
7mNbkkZcnPxE/LxM83WaJdCLWxFTSp13kyqacrU46brTal7E34wILIDFMFpD
DnEi3B0F7yuwOPwF6wawZQwXPC9kvqucJhFSRYCEStktzv612T2nJjam5/hU
g5Q7zf2M1T3A445UpRFI7Z7F+p4QVU5AAG7VqrPM/jxbjUd6Hj3Gzzb/sonm
I8KC3F3KsG/AGGwEQymLAMAs3yBlXtmNujPXKmcew5w9hOo3JdieGH31bm8N
UvyB48rvirdEj0ITG/z6wux/mP7pXB0KlFe7Px3VLDQ2LQ31XU573cYmpcJA
aTKkUXGUVdOb1UgYCfx0P4NiS48IqrNuoGZrdSLEAprCacVa+nK5J/FtECpB
76v3xwNdsxsGpc6bABPKcFess3QdM1gjQKpbgY8u1vWCt52uKFKvQouExqsT
7UFuJPBYGBmGcIJ/O+5aJNWUEEtDBK/HaJMeOai9NotriXVsn7hIvxvSXHgy
KfUE2LiHaEHi0YMbatB9EoEVn1sOlI042YshKljhvSmpoEHxDb4l3jN8S48u
TQbKG3YKdfJrXmMI4LP3c4EjK19D2cFbPWT4M/K4+038iftEShO/bfbz1ji6
rShhqARK2wLT1l5Mzi7DcXqo0o86Yrkq+xqDuuzqvPG9HhqgS5XoxxnOyq08
BKmyl5VapjgJ1FJpTIdZhO42387ARYfBrEWC1ucrD+CZO19QRGrlU+58XMte
RnaDf3hB8l2m0y0nlKSpDnIZ9QcKU3kL7e1CsuJK6v5Hz/oUttsHYK2yXU7v
VoTtgkHMnH+99S+hDfVJyR5UlhclM5K2MNvP2OgUlemNE/LaSDNgYmUDbpxT
K/ZgtY04bIEvngOPB3uxHuYh49m6wHim+VdfLXfp5aqAD8xOQIjsfaenfqG5
HkfBaEAmyRP3nf6mowy9YvAqyJ73dcm2u5qR9vIenuU5fwIdcJrLExI4ivah
AueOreoVv/mY5pY/YqkNe3FfkHiX57voo/asNXaoJ1WpP4cKzyPBEY7HyCCE
90KQloLDoTcJpKXd04t3x6lLDvstap4BY/GVbA3uCED4wyeLyKYD3cI9hinF
dQ4PDJT4NMUTXrAteeh/4L49n2izaMUxi2sHzrrp/XS3BcWssA0ffcHcbAOy
6OMsD3prv7lNKdsHppyhsSy/oZBWvuMEhLwTo8pVmGzpvbUNmCm5+Lgj8tgP
1SD3CSZ//gkdT1WL9rccPN5uz5d1Q0HslpsDQMarSt0rKH8txFRz7bkql8dG
PiAtZBk3dvAkKfu23KOaL71Ch+tl4BlnAdClUefeQbvqkpP0Lqv1xKmT68x1
Z2kz+dJKw9SOaFvmFFV3dJi+6rJsEsG/CzALhPs/IT/iM3gWyTgQGreEiurr
pLTy59LVHraR74ZgRBsH/rIms7ccvqPu6mWv0oD47Wh7sQHhZDsF0O6VOaEz
6Ew2gW5yivCPuAHsGd1nxNgfXbH4KUGT5X7pfGLqcJ48T9/Sbxda+dIswbss
xf0cUuaIqjmDnzR3m8KnE4tgol+aA04WJr77PDNdgz1HKSydIQUF2XE8Kqxz
NfM6WGkgpUUDFVVnvvRy5NAuxSOzwSWFACbd2QOf0ziUbKh8Emk7ocqk23rx
bDSSIgfkiGz8mEB/us0EqfcXwnwapE6ddhg5btBgDM1oQVof8HpWfJY/sF7C
uvEjGyOeRFxGOPjVWJbajVySriWOxINumoKv6XTAV/9Ayzp/Afue4F58wx/m
na5DsJD/w5gWLxLxJNvl+0eBQbd/t0OGINxPkQ8aoAPxDfCpvJOVI61dgR89
d57On/4Q5W2CGdSe15qMsAYkIBpIgMvjOBbHAKOdU3zSl/kuwMjidH1kljUq
z1UMxf1Cr0v0YibEGdP0yiZBZYCLTbWL+FGD8Ae0/Guu4hHoE+BojnfLzIE9
9D6w6SeorU26f1xtXWG1nOfPaYA0SVhyaMw7j6nWL2OuHvDlEia2PWfnSlG4
wDpYcfF4/+lkw8gxOhlnsl18Sp6lDMekvNf1hj/Mney3ZXnm/nOEgAaWibOe
nPIc4QtIKB+o7P/KMHgKqHSYRVT0tcl8+b4lSKqQtmxKh8V3ylPNpPojhJdI
pwoSXSirUTHWYUA1P1XebEWiCcQQVQTkKwhs/5sGhQAIX1PCoB1Hza0BxWZj
TTekVnxqh4g4H/1CaWkOjC4378LEUi1Etjr0Lrua9fMPovhGcaweRTxbS6Zg
1mxumgai/D40xV7ldgyB9OF4p8LYURVI/HDgbr5uXSNFEWBSrPxyTgCqCvdF
Ccf+ekDsULJVLiJD2HY9VJSQdXP/X2Lf2QsnxORLjXQfYqSnYaOEUmmi+k79
LB/Cvg135iajrWdHzPHFVhuXOteH3yFBNn1Nxaxej2v0MC7sm8IYoK0WfQsq
92X/6fqG4cJgmEDDtgNb0DU2W544n/oxUjBWQLyDlEeeC1st2ls8YjR/Nhbz
xetNWCJ/FuPEcGae9v+l/Z8/LR3KddA1vctuaUneIIvK/fD8DIDL9xmAPuSt
x2fRdQCp55MBhrJIq2E/eMLvAek73Wc4MHNvj6LFhUkFC+n3AxJbo4AjD7sa
f0qxENbEe6XtmAN/B7nzJ7GELXPtTjtMLUnQPPN7zyND4aFbVpJoYnLpO9yO
inPmsXj/78hluxsISm+ieLD2G4FGM1pw+mx39XpbETNGwcxF63e5phNP9Aly
I4OAFdRIk1X1kC6rWxz95WNN2v8w7Ldo3BsRSEmUY1s1CjQHsh7ll60Hm/3/
SlAzV1m7HPOt0sDHGw4LyTgalXhqY7S94KGoi+LD7J3MDU1RBTVmTPnWpk0W
xfG63Cov0JACko6MLePYYGeRcbu66kQRQcrC0WPzxH+94D2/GS961m6XoIVI
EWaTAL1AXBzKxIdffZfYkztdckpotcY7mK3b1zMsszfnB6AdFUDFZIftNGlV
B8ZeK++CDKcMNIqJHiI6JHtNZVd42fkyP4IHZOgR/VUdkWK2T+7PAR1yqVlH
Sd5EuG9neJ2a0uLQewkQhFAGvld9DBV8AJ2j8UZyMr8MY2qxKAcEh5WsvJLF
+KDFL3TSmOIVPE66Cq/hlBDo4Bc69rECsTqNjfH+nnf9wTMeOrmLrJ6+Nnqg
NcDRBy+RkoMh9GzwX1X+9ZoZBPchWJBNRBR7KaXkjC+wkD1EgiBKi/KMkoZS
Hu3eIhXoK0ahki4Vl2hGMcqo540c6DFB247AxJo+z+9ijOvL32RnnDvaNaqV
Lly7Ebi2+e0/kwtbejtkqQcp/+iU0ctivg8VkDxlW6Ko+OZW1OhqZ0nuh4I2
PGMvs/bgGzP9mIpNx9qDxLoLJAYrBxjc3EsPmJxIEjAp710lrKnLGV9Xoj1e
pWkMO7imW4Z4auXIqKUlOFHqO72COTbMsIhqAIYIcpxEGHGinYspee/72lF8
Ll7nE10dZZENWq4sMooWTyJEQocliL8gBFCVYeGMd3jhO/cxLRRRdxAt5UP5
sETVjxJRdLDZh4AQixQbu9j3rUHKlGD2q4OAYdvUiU52xtOvYWryIvtUjTo/
j6la8P6LG+m5yfsJEHtoFqRuASE4IqAS9+QSh9FkY3Hui5rJnptqUNTIIY1W
t2ulvuSfbMajkYw5rTBun5qPxAQNSiEu2X79KIqddiX4oHajGQB8tzTsDzSu
KFPyn0Et4us3FJsUgzDBpbljsH0wDZz+Mpw0B25fVdyqXCIQwtD97uBlRadQ
fU8rlrQmAJA+0edZ7NQ4vAcljNfiJqkI3JJYTCcceOu27jBTz6enDQGWtxYO
lUtmbP0Cli+M07CoYMrvh5PKey2fbXoZhXVavfztxeCABKeKDZlWp3Wsa28A
yDYpAr7K4bvdl35Vhw+RyVUthhEwXRO9V36aIEdlf5HBqwdnm/w9MOeBRYiM
1vOLrKlhuf0vBRKF4pZqRE1SQwO1yBeHwQOXE4omX9eP65RMlQiq7BwgdF+9
YZI6WLUB0SKfwhKT833IZBJfRhQJDmNGoqW2O902JXVmy70+fiVY4ncNmEXm
unb9ySTN+y+A5vR4xfQxHWoGv0Zzo29AQe6T+zxzeWsEy05u851C9k697kdF
e36vbWfbB18nLbbCfWQFxKJK6obiMgb7ZKICTxuH47ZKliD3pvxPVfGJXQUj
KMfUiORKtPoyNGZzJzOF6t5pAi9eKOqN7slsiGEZItBYf9gNJwv2+aNtDapK
tOw/u8UvTa8OlpuFb7WkCW0lkjcq86wgmbtvCzIu6EF6E9PbyyrZG7ylGNab
r+/XphzoOeAR/ETfLeYuNaXqKNDkBle2/CB1eiUv3Lxcbw/YQ8VbwQ9g9dG9
7W90qP8QI4CxSFlpvX1k6l5bHENHigIuiU60c9OOssC26vjnAec8BLgyLlg4
ZiN2+8959HOI+uofYsxPZzqzo5CJ7RvyENfXv1H83P+CJUZFodFJ/tViCcQd
LJYgVp9vJgdBEzew2HDOlVh9rUezlHGJg4vuQ3jMhfJ80YQ4HKee4bOkC2V/
Oak+ZKB2HImBUQFn1JrqQvgW/uehGpp1rlYBmzKzCGtcp4q2hjZX6Cw8IGkb
n8uNgWx+mYqUKXzAGcb7NLIRsdoXy9FggMuIYjH43oPHZ8yvKhobD6nEX+PO
qjGbAVKnClN3/wr5gnDiRf8uaVoc7bqqzz7B1PxnI1/WBxlFClKvEJJsZ0ZG
hj0etos2/LrrsFFc+c0cvBrM0r2CMnKjwVw/tcO/4qiIXGERpc71NUoEbI8H
8MEl9cBlFNHxQbHuVQTDV4/wJLBJmOvymlY6tSDV92TeBYrOi7VAdxPxkacA
adnmfa+Bl2QJJl0DfijrFGnM6Anq+knOYj1UCxaHSnhpkuSD6+N6maQ7+DHp
TYjAhqQm1kwzq/OYxf/ZkeWeAXW9O//HAU+EpxIYMvWMFqp6d7FmeemVO9fN
jcPerx2eyEVg1ABoS6iefb7gmgPBoAJLqj9JX32z/+XhJxiKN+0uuSM/tS7x
8+9VlS8PsxU0P/cW+9e+LdPoxL0Qp2GBMSV5Bu+1gcPjtoNobHwIUscIjLSB
DZM+nLyL4UoThDgkJ98tSM3c5Yq/q3C65i0hQF+UhnKFnNsCXc9Ko5Ykuapj
M7WZm7l0k3cktSUYm9ZzbNp0OVgjVqPn5PUVG59UvtPYcufYC4eOtMAGoMgI
acsYbazd0Lu0PGjDwvUlkTD4Cqj9cAubw1xdPKIq+u36sOnUKNDbAgQOURb1
x7J6pkkVVqjVaKjppURAzvzB/0kEhpElOvs3gVIts0XJpJxHw8rpFcE/T4yn
PMVtC2wx2QSHni1I2L+na3aSUB4NmtFpiNA0FQTwvJ5wRbvWr7k+NClND0hj
N6G6af9jRHFZwg2tjR38721mHk9sFthk3TfQJD7pkGqdktX/FiWKDAYwke+n
lVC6o8RkBhhZNLEm3oDeK66jZ1txF9YXJzSTEAGJfJAE608uv2/lwMkL4jDS
54MCqjbAd28iNohiFTcGO3gGctuGAv00Mz3a4WVwuas5u4V070KYRQTGYatN
jtNV1t3CShCaVYDZry0ju6z9/T/OZrGEDraYR7kAofD08tMbCEcLP433ZQfA
PD0yQta2nGJjyFJHnsvK+LNa82oowny0j1ZK354CYkAB8vOCkJqJJW0K+/mQ
fUsZRQHp49mwYuKxjCt9z37nULuAFK2KOcT/2RnOBVbr1MloS84JDdQCtDCU
awV0cnJv4wXFtteCSQxjZdpLHMTaWUjxHiYzHm429JjzhWIxH7yOvJ7z79+J
8b4jnyuhwYz/+cfd0kLeLfnTt67MoF6pEL1I55q9kGs+kdB9KUJMmA2WAthw
Yp7rWB70taGq+49/Vi7maO+K3M9SHA82c6EnQ+TXQpVBsES106Q7Ae2TdL5G
NnQZ3F81gh/S9O0lqH51MZH4o5VHlo8bY9jGhQIkjJiMsMkslLyR1OpF7LAj
GGcGsTG2W5vSXXtaW45e37MgftalthDoIEcIN6eMzevDSUmICx6uv6liOUmv
hC9Bc2Qv6oa4PZfV0nbsTlvjIJ4Vgx++xwWktRSyVQFdH7kO0IpFnzFycniO
sGpmsrkj/W6ZNKBipTJ/YNrgSeLCc7oa2LGkLMZJurKoatFLPas19b36AGKt
kiwE5fD+9gIHB4C8WFCyPQ5kWqoR4YXHlkJ4v2rKkMPZBl3MwqUC+pi8F/DQ
tNsFoByxujMlvZVS4X81Bk0XvZCZBCDhzwAkCiVZENWXw5wpCNynEheJg3Ac
dqU+A/z/V8ITsLB/qRszNslcHnEB13zOnr2JXIiizuEvEDZhJ5Ca1jams02M
/w/1Hyq5TibiDY/MZW03WwYDCnJ+yUx7lSqMlZqJs9Q19vPPTJSUoRGoLoQR
9RqaBLdQwO3nGD9m+5PmyhMDH/PImeKS0lzvbBLd4PsiV1BUOzmZwNBeduJp
r3slChv3lLvcVbtve2lFlW8lfkdZIo0lCSRiEN0K1jOSa5xSpXbViH9j3TUy
nkHvp3CHU6d6xZmyW5q1LypjhMwr0YaOOT6HDgf1A0+jlTB0gh6ty74aoiPW
baWpPXeeISX+D0elC+ebzn8/U4fTtFR3PZXLyzrfCMJ766Y9ZqjGSwZc6zH3
uUoIfuWwk1GJkZdJLbzE29giZwh7Rn/eT0EWahiiaDQ85NIDFoedfP0YLAub
K4SY8VJYmyr3r8q55Mgb9T8QuYO772zM5YJ/jsk4D48eN77LmVQ3X/39yxob
RSARvveo+VAUjKUQUzBOMZxhOBe6jXMAsISXbsovmddbKu739N/M0P5L7g7i
vRrsypyT4zYkAOypQwz8G9a1aPN3TAfznQ7zHUIE9UmrQmYGXMPJ/6lQAhYq
MmEtYN9G7eI6uzmlHNz5tyjuxFM4C/cwWlZim0dUJ9RMVIh9+EBeyx7ggnK7
5Wr0iITCUp/FkBe+iJ/T+knW6A+LgsQxRnLMtrQpJKTYBNqAKRPkojH3fcKu
q8Jg5CsAYOR/LKD6kGr8uO1ANtZDo5KaO3gRPvS6FKGrJw7ML0/jIkuG958a
rYVcxpQsJt0noA9swCDT0ZccJ6DqrHNXdZ1aD3MuTGUiQqvEJTDkPjG4HGon
VGufh2OcpCO8yc5/GTqYTi2zf72qrFn56qIyme8RyNdF1NIC+R6g4LM7VcMc
1q1R5xqPkPUCj4CDV6MzbjNJDwFPOM0WI4RMjMPRuzykoDWx39j67+NzuDlK
i7KiPgbpivPWDRi1i6xijGEwrdCKgmaabBEdD2njOMS7PUABeVYU86Xm+wXj
sByV/eCHSQj8pt0BT/uL/gKdtx0uy6v8LsJGE/f8MYzQL7B5c9Iv0+qWoZEy
juXUhqr0TQQycEBpakRS7gfqq6smHzVYVI/Dfeqd9SA9mxoS+HPiLdVwpzLm
XeehSWrH1hUSyGEGmn4g7B5fmD/uBNNnpKewdKvVbygMXLl+2Td9cGxsy5fw
XZFEyM/QRbJNwq7NlRR5cf3Fr54kFntTs9LGO28K004+LbQugYG0uqTTsWWx
na3Lz+80h4XrQkuGL7FLMUaGWQr1gsPy2jImDBAA7q2AaESzegnPk5sU9PZ1
uoXiStmu2pUsLLdoPweHsqLrKd6mgEXiXzZjAZYDbcUvm0qo2eXL9+0uHs5+
tzNo84bCaQu+4moeFqnkPWU1C3caqnYHrxCC5nipmb/Ej/t5xFh3+PvJDAhm
sp2CAkDedJQG94I2yuP4aO/OkITtzar5Goo8daItR0ly/8EKPkoQHNyVRb3B
xyaqVPFnRrsiKvzD+6MeUaWYMQPxG/yNdxIdLW7W5QxkMhd1BtWGc7ik4MJp
OdMMVIXkkbnic2EShDvhs+D1gGPoeXo7ijeTh7JBhMHdfZYaA4iZLMoYHjOq
NXJeUjt4ezll8bR8Lt/j2AZI+mrxrGns1JXTviPqWvr7ba47xGgdn1k1KbOI
slYEopWlQ74RqynAxuxK1gp4E09hirLBjWvQUxTeCayI6ifNaV6UJYYjn+Kt
kCdiSyZPAbL410zWjqGnFVP0QLwe21jhxwbTIkbodnYX268yrvn2A/eX0+aI
ZmqI47mDEnaKwnpz44L3EkZbbVney3Cu316T7S4zlvN5/pZG/4c92kLhvrtL
R33MGez7EVCaExC6WAEELw5KMjuh0eVXmjZgGJs5fs/bGwbDXgJXu9dIo7HV
tbW28lryjw3jcREHAB6lHz+UOFmSQ0A4sC9lV3V7/qxDIEU7vUwXHR3qUdxM
Dw/JkzgtN81OdlYj6R/iJUt6olyTIx5f8PuZLNDkgCcNylN9aKJG+GgXTBn0
bM85une/FNwp7P4kxgSllNLD4Z/2ySUJTvRZSGtIabbGn4Rhe3m1UZvM+lcW
0MJNyzcfUXuNy+IZpojLY/78Zlu4rN1p3LbcErg7LnV+wb1L2kqG64Wy3W/K
3jtoyrDO+s27Szlu1E8XsuIwubVYMLPId+ur9JsKuNzPakAluj7akOSEWj6H
kE//m+S9xkutzIJo7g8VCnCFelIriN55/AxrBxu+S1+GdWPKKvdVAgcr68WL
BRjmAdOpxIv2JnoQmSC+fZilJn7U+d+3bvD5KLabRziybimjB5zFlXKA48Jn
DHR9UGjCiJlJVMdSZ804gxGSEqbn9J+RchmFREFAAHQLBbISSzEqKXzHIDGe
VQlvgIxh+wY+2I6gJUTrX2AegcbSyC4JWCoymDjM8SWn5EdgMRAJdrc4YSN/
VgwLF4fGZMzCgLJc85dqNSbIyqy00wY/kdcPWpBdMZkKVLUWV6Zjxto5cFOG
qmCMAdGXghidrjqL1QaYWUOmrAdkwnMI2q8ZvMhk2D2uXNkyz7FIHsw5cI2W
l7vuYiB18arvm4uUbHew9o0NMdwLUFTgZVwjXKvKtqUmSWJhZVZBcXF9yQV3
6GW9kqoJMnr6VKhqb2uDxjbdgmRUaAKR8Y4Ki4rWOBvTGJuXocvtrw1kJe5u
TnihShX0sQ4rcWh+NytoLgVxneqivymv52Qaqo0nJ/YjbpxVIjQuil4dqmN0
HSWE8VOG7Ip9MG/oNPMQ0Tsj2FhgO0jx/W+cEupAWV7GyH0CSH4PAjbrdLPT
qFMFpiQapyiIeBb7mKzdgF2jl8B6sTI5RIoukoWYIcKUzpj0FTengSiPN9m0
2xZMAOxqhOiqXb8moW4SyxbCa5S68yCDQ+IsQWsjaXn6/76MoECg7X5kUaX7
Q/Jf1NZOyzQ7ogxBmExBLvC5gtlXroxBKJxg6pPouzMs+ghimHfp+DC4Y+Zh
dYbBLsr9pud3Bvp/vKrmXw1LHzryFLDvQAVoQL+rZkn6snFeiIZfT9hSxy33
FhwclEpLE56/kSFg/a6votYoCkjFBNxCNLk2h/WrbWhg2vUAdlLbDkIl932o
gogao+42RLcW2qQoEWCwXtpW+hpURfgIOyAJtSgTmMavP09VHcyeZEK/qZik
m1K/CqNRLjZtZCe+CJCpc1FKXBNPcf6L69CqvF0DVTRMe/NDqsel4rdnqa0Z
roqLNJK6C3cL3ngrEDyQLLed2iDJjH6OO0eYaqp+9V6xTJ/6HZ4A/TmyaTuB
sZ1na7jqPrR+tHtTJK8S66k0OSVVIePqzOMUj+9wYFI1CnV0WCJzooyHaYnd
6WPB+dprCgL2NoZgf9vk0hLex9LnBXJBcDuUgXqPPt/vKFTVlLUrMzrUYRX2
tBScrAEoKDv1Pw5/0zdNMTTbcOFv0cijJtffpnNzXe7G3t1ew/9Yd2mI74/W
wt6gWcFcDSJYnBSFqvudNGbZIKUVbFLSfxfwhjtufgyFyrpjFmogjtwDMrd3
mnp/BSxARnT43P+FPFMrVtWH6eXstb4AKlSjMGOoYTGLXJQPBZ/UInIpwGtr
1tOlCxBcrHLBwBg/fnl1duIkI5hSx1Ebqe7rrxg10NjbwJESmTR3sh2X/P5K
Ttj2263vGZ1NqTc3nFyP3apTn7WhgNyKE5GUh0mKPQQPc9CtN216WLJK80ow
C3Y4SzN9zDRkIcvnGA87DbYsX5W5t8qWwd/6o/Cs6jbafhXIGxIdEt0LLmBR
xEkjC9vwCI9isdVte7NVlNnD8++buFlg+lUhfoLW4186GAPghpV+4UoPf2OM
86vVC0jpW6zH39OYxOjz4/AaEV0qGN30bB6VzFwT8DnzauybxjJMDwGfo1sI
tzFlNrmJmpuGae6kO21q/uu8PJle46W5J0XfJispKMhMJZ6/YKxHzplhKa3m
+UNpAPpBGS2yxzie5woMDlaTA3LyArEBEPTZKbLgfev6mRFTW6mrZhYQPx4S
m7Z4PNKvJ2ffCA5sZ/ZNCulWiRdSA2jTqSou13jI4OOQ4hb4yfQC8Zezeolb
qt2gDET6CQ94zh6ZTNB+jPvcHg89OWd50kNUy5CyYYqo1G25Hu3nHPXjPgeT
oRt0I+92iZYevJmtOJNa3NEb/UcLBREaSgEprb+4Z6u4QrW6Y/65lmO0LLQJ
u1ju42mt42MsyVWPpPFLyKMWSzDupRyOkUNT9NJ4RBUBmk/GR+gvVMN2miGJ
E0tkyF54BEYDh0oIn54UNqyOtleefcCUXnH2fSfoPAQkNgE52LalfaPQPW0K
6XiIIIQQ/tC335L1EmoxZVOIZfowkUprhx0cC9mboriWKtIrKyOctmd9QgHs
OwrykhYvYPm/FuG+bISiy9zZv0VpZdq2TEqoWLRz9DiY6QfyyrBB7ZHotx6i
CACNOybV2x/jKDiiUF+aEAA+2S/DEaJhiZNktv7BtzKRjp27xKr3iG0o7uq+
rysA+tSPRkOS2Zoyoek/37VUzaheQ9VaDbOYMnDAiQChuuJUa7V8mEEPKXP1
D6X9AnDhw8YEbILU6V60w6K5SJh+HWrtvxB2F4POPsvgqeNCTbGnJfF3oTg9
Zi7yzmWJ5MIFv3FgHYPIBhkST74n5bEbdgsDYKGzCv+POm+roTzRzKGYcAy/
sYS8ggBBcOb7b0KQVb4dgZO5EKvo4LTA7pKjK7LS83V1d2/nVtvjWLAX7Ltw
ekSrFPwfXJw//Pie21evvtyw4DniSbYwV+6U5ymELONgZLAHBHAAITrTcxTp
wCrLIwBV4HbGgMoC6rP2J0yRfkndMgfYqVbmK+6CCL2csyvHsPKIWt2WjP7z
uwMye7Z17zR4eZb6tBqs3fbALLm/+s37gwCeET1UWp9DiRzSuh8O9UGuSNha
BZzYt1s45YSevfuk25ng//1xTEKUUa3cPK0KWZguvRxr4iMEUxiX3Cpt5X1a
p/Hkh2p0clDOHak+PuPurPvv9sBVcmFYezpWxOaMK8ywJRIw6/05bJ7vTPoq
GPzqfP6mHSE9sxrn0knfOVcR1LxKUiSDULlSlvB0N+f4W8q4H3QA9ficr5SB
M+F2zrm182Bcr1Sc7nwdWLQBFdKPcSdCqf/WwJI772jZ37ItmrnQfOy/rNQK
Z8UgZnxDIbVd2mksrZACPD1OMGMnJYsu25GER2pa030PdPwXm9fbTqK4tuBU
02s5FzIBaUXKGha0u7NUfyj8y889p0SjfUjXxkIUDrBwMKmgD1rG58r5vHMZ
eiqgDOLL60Nno+Qddeyt517Fj3GLbQ4aZi55FaXl9QOQGpU/SddNd0KX0lDE
RPpdxMKrpyKNAfp+o8y+Dqm39eq5qtY/o26Bdd1q5xS0hg4gfpJXwTaxJeZq
6frY3+ed3DXBe2L2u8Y9rtr5wNVKgRdULxPcg+XPu4MAY5IAtjk1SFrjgPjk
rP5HeUPv22ZGk2JBb9X6oQNash1UjGs37ndvcudBhi69VNeFDCJXLy1HkMEd
FJehLF0hhtCYMZoc2iP7OKKR7RMfVVIgoe/SmNf/StS06V0YKgaTHOPP/8ie
wNeUOIPTh+OpZ50ZFmrx4ci46407DVaXMzbjMSHfLLWKReGU0oT5tMlsnV/b
zeEvWCci2Vblhl0OAwv3i/uQ3kYGdw/17FzVNVkw1wdmtP0jLaRfagmmGyqA
6TZwhCIO6PVr0/nT7c+5+4qpq6IQL9DXWTuK96fNNE+cXluIadk7lPz//UO0
2FURa/xbo+nzzD6/FwMYH0d1gYj0onChAy0hXheNe/c7z8w5KbTZN4E3gOI3
pgqOEcvcFcnN+108zyLSoveeoxX9uYeNv8dVKo6ATiyNRxHNBKS1pXuSEsvy
Mdb9XgwIC4H8xqVu7vLb7ABhk7bgpVQuBVC3iHniVPKWglS2sxQCK8Lq9ZnY
tD23M88w+AL5OSj+VggC5SKWxwhWdtnzu3wRdz3hsfKU1NCatJ5qBkvQj+lx
5cFndUWWdBWte/muvXsYeJZxuIPmW2rnWhUjQLHeiKF2BVNbewoC+UEgkQjQ
1ftsRx9gNS5yZYwFfN7qc55oh6EgLRoxZVBaMbZLm+Nus+uUgIIgEeDqZ/dU
JuOXA5R9JKWePWfyWAlBlE3CegFmkG+LAxESelydVqbxqjy7usXNsfNyeG5a
e84C85kI29swb/9f1nit5wsN42AZDZmCH7qRu0GWOah4I/dNYs/RRaYXwgmS
xBUqDF8FzwxcNQfO9YJFWIFwMRnjZzwvDu0rl3uBCBqiMWRLaOg14putJbxf
FKjwkkBa0TOodnPRo2DC/W7UqBT2US9FhUIjCkhFlg+GGPWznIl5vUCWf/qD
QdqksG9QCvnaSKAmpvq7AzOKDUgRnqAgul2n/T7r1/KCTrXE6FRaV6m1FNsj
0fY2mN1A6W+8JimpiG23CfIQoZoCjIUe3BzbzMmNq2j3w3OvYvKzMyyLvgK0
C6OnKtv1elAhjK0kfxWygBb4x45V3U8zYc9Vg8/AOGaeFnv1HEk+/RrTjwNf
ohr1rVtJMYhY2pUuXA1MLwqePQSdJYTwMRzyN3h1od9e5bHkl8IjerzbM3Xp
/xr0R/plNORSkzyFvTRk5e4L8FYA/Eq83Wo9n0kmrmUHBUFYYDszH2RhXtQY
oAZGqoWnn8av3lvNlS6a4wD4c+9mq5HU+DsDyK9S3wD40BX0wpzen/NRVV+m
wqLyaUQQBXSD3AbMvS6PeM59mPtU7QUYWOJYt4iQOiFTZiQ3sVNzOxbe29zx
a/yHH0anDeIeWbkxVfODiMmbkXPStwU1hOtFk+nqeOujPfP5M6QcovqBbZnv
TfVqQVp2rb6oINX2XRDay6t6+kzMr0oalLOao/eLPnKGA239dkA5aoJeEMp8
I+U/xzvlFfk/dbiZolSzXsC2pzhWKgly+oXT8yoKvYhCuXU75//fMu4pIQk4
TL++TVYz/3mOoKtp8KHlS6eXw8NgcPQmwW34D5Rn79LGOJ5zi1l+08xwi7vq
a6NMgj/r1spygfmVhNBmoZ9UvLwp4P2zg2sEazfx1XRtnjTe6F6/7w/dFPkd
lOCE4THC9uMAbcFHNls9LX/1yA3mUsNbR1nfmb2bQj+ZeqXihVheSpZpuU1x
iDlYTgOTZiTxHNcAl+ax0a3GgS4fQD1LDqCtrfgA7DwHPAV4VTznW2TdifiH
e8qeaaVkaXjlrxd4txoEGeJ4oiPIndtiuQlh/nO3qMIiKxB82n2cn7QGet+m
wTA/aKNWvkSl8w6Q/Ikk/ETqOmcGd5UuPIKpvQDj001x+0k9KwiQZJUrdVJ3
O1XtZ3ZaV9xqh0zL6R4MzRy8tWmx8u2NVsm3X6DJ5SeZEniRIBRRyDXhc9FO
SfSIr3+r5c00TcO8Cef3C6l1qhkVsPzOe9IJ3D0gPG9foxrReYXAhEMbhet8
2hCL1NCQko0yjIBNoHTKS/ElviepI897WmqHiyL16cOXuxCha3smzkNwQy6h
FdGz/PGk48imc80KFyKb+nvGXUTDULLekG8Lega0B23AnOP87kAUZlJqSV6E
v6kNU1nRkSmzD3+u+2vO1jct4738iypeLHf/3+cRYarGeaDmO9stxUYN6eEa
HhELEWPzj8K05mKzMTFD08YgbPj4FsWI4l3KDlAabjqxfEeVWq+Kb6q/4da3
OhKd3UGs7Z1ofJCiZf2qgbs1f7UihEqA34p1Ycu2A59fQG472t1NaOJhcVvy
R0vY+QGdaoRA0Uul79JV0Ze67T9VxRGo4EE6TsMtE5vuGZNIqVPCwOlJzdOo
LZn86aOrxl0RtCEJpNAWgS+Z7N6Un/y3WQKFjpiWfhBzmPT1WDA6iOUz3NXD
KKAt/8UTzOvcTpdf8rPOt3xLLvz3FO//IUGvgITwLZ7oEp3Q68QqHV094+i7
gbdSTnFXcj7apvOhtL9m1+zeYcDvc+8J1HWgDavW955XfhiDl56mIsrw3goo
ntpC8zL2NX5zWI8SCuZwnMGv5oWwmRGFhetATP6Sbr+6zci53XfweLfhlNjK
nweQxckW0FBMwDE1GgldyUvAf1eReMkTKB3phGwVYUtrTcq/fMaNHnPVphKU
JQXyztvijOgxsUj06jUW6eO3IwQe4K3upJWJlxDvakN2rm88ySQLDYtHf8HS
FPcViiLMyDAyZ2meAdjMvA7fldmEvezrPrJtmeZrxKBmBG2TNoFI40/+ALHH
xOIavVgGvgwqBKn6Wls9GYwdfOQpQwS15TMA3BkdhyfC55e79P2+mRXf3kk1
lyZ81ulADuf2V12QketS2kdheM6kmgK+bQwDvOlHF2L6aEdDLU7PU3eYmu0v
OUjYJ/kyjlPNNJtFKcFWmMgEGYVXEaQkgZOM54kNzmKbxIBla+9z2KPLJ2/o
Lct+HPUfG1bRYwYGw57s/N1iKpGHuPMRsfBlkwduT2UI8fSmBlOALXlPWkwV
LJcj07rVLK0i6u1eNt+2Y5M28IwwB5DMscsrUnXKInAfGv3pQWTaV71R/xVC
st5bAiO0TfY0WH7auKa2DdVz00nO0MQaVGi7J3c0hJ/MT6qopAYuFx62yyA8
p9VEUeRkmBfNBgTWxjhG5Rt3wNLwImPGioWGFuSKJZPHNNDE3s9cYjleYtjs
iHFKiQc1ymwoxahdUmUZEvFu0UiZqwzkKPKkZdZlSVgI0bjh+58fvNjOx7Xf
Z+kzDq0sf6Q9cfLafXP8vme+rpz1Gh13+PXzwbiA5N6DElSCSQGPL+74z90S
ZpxlujS/SYunCfxvEcoR3PWOi8aWa5eLip4e36Y8v86ziGUtlPP+vKYyQBRP
Dj7QHHXYlKYa3k2gyHYYAg54I0dYwbFB42FxW4ZRb+Nr7WyZi0lB4cH+WTFj
+pfahBq/FUKHDLfNpvvDK7CH26Ad9TAYQVvwlUb89nkMuD8l6B7H4iuqW2zr
cqVBjdmEsTIuNd067gQj5n26PkK5+E/xu3T6Amxx5BLGCPYDXAw1ed1ADGDi
XevQ2dRwBKZE7IA6WEBI3Zg/nhe1aY7YtVvA0uRZCutaVD/Ue1ee5DsdGks0
E7jb10LBwLFZvllH91s9Z4h2NR3jdHrqNw9Ky19nlSbtzq3JtTSsvnrmg642
hCOeFt1lrAjUFPVwJT/I4Z1/ejS5uqAVwim0fj9VPVoND3bFzVkaMrbb9Zii
h4PH20Dx9k9+rzU79DHLvi8HAXSqVcWUItUpAgABQXoF/1gvrszvfbNeyypc
NhoeeO9myCZms4xM+JhvzSnzqM9qTm1YiVSwRq6ASBDKONXA5NG2JjFPkEv1
ugwW7POweJfAoPkwfN9X98L0GaOQWk6hHMk2p3tyONZ9UNy0EO/wndAmzhqR
mSeH9vI17qwji2xUwqoT2g7I7oJvEgnD8abTXcA9kgrmQYlZksfh4nbIlSaU
H9Q9gsCwUUqsMpjbdhwopGYq3fqTybbtH8izO+Gmw8HT4jUwWMXkgwEhWTkw
DWzalH1DJ56kIzI3Mk/z6zjxTHlKldvCcmG5oBB1eNVM8W5h0Xef7EiCJSmu
l6CPsWajF22AY0w0IPriJNa/pb+yLozugILdM2bSIOjFmKSUHFJLAVtIN5hM
xL0/Q9TCezX4+krye+3tM6RT+yvco/j642czvqLGEjZFmnjsOhztKgYw1+lW
ssMyvk+V/inUO7f8eD3P3pyOPaT7f9M0gruPHQHts6uPaVzDADZvjNbdKkdp
rIeJRMp8gf4miD84S/44k9FHp1t/B33MebBYhGcQccEiBOOq6ahjDjjti8xu
ExWDy80pkeujcA/gP5eUTh/iIfp19kAgWSqGwU9qLA7k7NX6hDEpQVsqJYos
YO1lZ1gE2ZPAQ+RJGVpM3OiBml8aKYhtlof607NMuJtidbwVspMvnq9QIeY7
7siiy78WVPPTZT67iy27nKMIFIz79IeWis7eRTCmYlkrxomYfk+pxB+RTP+8
4HutZ83ifCUA8tdwTK7xxFKe637U+8KQf9RejkGOfiyoUDDA8o7yAaoicGaB
KPlMyKXjKjrWUm+5TTaQej5ofgAVNCr7gG6WNv8vjo0E8lheQiaT5SraXqYC
VL0BT6t4xktnn+uONw5iMp63Ielhz2Lv/hm8zsSPEv8yz3Nz0JL46Iu20Dhi
QgVRYRJtdn5oCdevtUZIRHf0tG+ZyA0aKHXURsUzwiF6vHZbFczP6Ih9RSi4
/hReagSHalY9niJiEGrVUrYnh0kx5ptdX59995a9FC1S3u83ccYV0GEfOOfq
AgA4uAOFQ/1wVGPiQkiUK6l0qfEzvgDBkOP60bxAp7Cv45e7l+KRFqG21KFE
I1E3E1R0aqIq6fsjpXmZ8bKQpxvYUPNbEg7jfkm9EjKNcXpBH2jZAWM2kngJ
XrP1clvmB4Fm9dc3HKtiK0xGuE9HKsCMOwRb/eIi3Vrb18DID4jbMHpKP0Eq
OVdQkRrqWoZ/l5bfeXzEHKbK/LQUUTBd/x/TlhCJPBRnTbfRLWSG0e0vrrgb
8c/dcxJ7X3lhnKIefFfLrpRofJ5j6+YaaTF4lLSFREI4mQP2MgfSUpoZSGvZ
O6Gj3CNMtT6N43Hu+MuyTmPGx7r4rFL7n+j/S/w6Vsx2oZgWs63bdIABiIg7
srsH8Z9WoYqALD5STauP/ucjSh9B4yv3nrJTxTneSmyELv34U1jr9k7mS8Ag
SGGT+QYkwIV0GsV08O8Ze21040GOBWVduGJpu+PlCUGDT4Ra5eCEnTx0brFH
CU4O1B1hk36yFdq40Xga/8Bbyab2VNnlWYqkUOD1Jxjrs2JJ6L9BHP02+SiW
PTcUnU1RrnDYvknap4xBUsCbmLs9es/amdMJ3iGu39jvhno/Zx8n41n8ZYBt
LKYAl04nMtAdG2mwqEZWeoS0W6EZ5nJtce9z+t0OC/65ynXB4KXEZ6AO52JV
iVIaa8DBVrmUMWGB31Kshpu8pImRL/2A5xj/r47LkXTSYLZnR9S5igusl0dh
F7YewHDlrzJY4vcvJ/iCaPUZp636vHZ89wL9n//m9vmsc4yvKsn1DMtvNLjV
TISIew/WYfAB5Mwu1/31vSXHbxYQ3gzG/Ge98LY9qj/tYgKejPu8TNM+V3DG
21c+QVIk1IaR3QPdetGspOXC+8wB2Uje8mTSvL1u+OTId7iue8dYkdrcHILp
zG+tkToxw+hQcohGHRnYhgCSQOnwsXLZwcRG/BF7ybxKx0Zl4rmLmhuqxHr0
3rKlbI78eBM9RUPlokCT14cagskwsJt9sFBX4dC+rFt+XvOXN226vt9XHhDf
R8eXEnlIwNobuXvO6M/Xxzc4s695GdEEbHsgOMnB3f22j+GeWceMqo1WEXiM
ytJCh/6R2dkbL5K4YSoX0cMuHOzeUnAq3jsnGHQ2szliRrltQ15vehuyhMkq
wx6rFyxMuu8Sl6HmcKtN4mGtdbsni3txjA29t4f5ZhS+NLl8/votxNMQH1sk
SotR2yUdXYZNDDnrdedfUuzmVb33o/dUFbtTr0NOcX5QjxqV2kAuOaL49Vsa
S7+8Q+lDfvmHWXMJtTUjJss2yUapobNW/A+5kfqG47bZgzOC7V0cVzkLruq9
UUpJqXt6+GO9djcCRQlOAzW0HiZssvTl1av9QsTbKyh4t8SHuCV3W4IFU/sq
7GjBEkWYZ/JrURtkOrSHTUUcrb6B29qL8LQGDDmpltPV7tQSsoSbNdnKTVEk
4ZKeutk8fhMXbjaApvHA8PthE+ZqwrlMlo227kq6+bwXehU/1gjSj2LD4v8R
iNf3UTtqTauzLE8yPE90ZAOzoGQP9OvZVY4PQighgNZI3AvZxuf6wRtnWEqM
Ij6gs4fHMv0JTTLlg9u6a2HpbMYkh2B6TI7zjHMwG3UOGvHHfdXrwkOSRJwa
ySa3yY8Zeeyl10mw+1QedfjWwEAw34FDLH9aaSjW+xrecLW6vTwx6clPdBnZ
PI8usgZpFu22TcboEEIJ5T3Jy7eUvzF//MZmjn7w8YBc7K9q9saDuwK8xZiC
+4zXT8uQHOJpJ07HGSa6FFPztj9bQNtTjZdMi1eHGxlj9hcz9zI9TJ62xuPk
rnLypEctfC0T6/7G2nsgSh+Vyhhn/JzAISyC9KQnd0fgeWyqTH0lDXOAO4Vm
Xt3BZTY8HhmcJ4gPCMNJ0cSvEx57JZ++riu3rgCvpq1K1/FHWXyfVvFNAiHw
q3mCab4AP9wHSuSwbePFMftMWKlfxBKlSMQTIZT40dLWPtVsm/x4Ga+b7eWD
qAMasdPqwPjgULuONOa6eENRF3rWF8A1dR9Es2mOdM+pRUIx+zlMXg2QoiGz
mwRGTUKrzxzCGJCqcwC7mm7d5RXEf7XsgKPQMtW1EwltPTwaegWtxviHpBJt
zJgAAd31s4iz87i7I/eOKhBCoId6juSRXJF33N4jxfUH/h2i2ZAEajNxkyPA
oy9Jqrc1bAKJVdQWA/hZMhgZc+b7B5h9heELtx6z/Ln3Occ4wXPd/gbJ7PMT
nIM5DA2XwJ7IZKPa+JKDI9BBI23Lk8U58Tq7i1UJmvRJHvF3AFI3GhigJIAb
kpfU+4LpZFEjrVHUlFQBuZzlkksfLLsHOmC5Ovc9NElbMMkEyDVG4hnTqql+
yfoV0x4HFt7hhhHD8AOsodWYjQzVbWlkCw+4zo6S3Dw1WOjX7W8e8Q0Yd36V
Mn2lIoYq/DAzrVsxVc2Jk3dpfgHPs41+gxKp1tARurp0QOeM1BeoA7X1bWzw
P2EJfbD0lpgkEZNl8WUmnoGaD/dCFQW0U9uYx6wFhwB/BpuV7lcHany2Vfl+
aV2bWEpOJgAjeitih+fN23lwCwaEYEamjXHRCXv+M5Dxt91hAdukpUS7NLXC
68n3l4oCg4oOAJFnQb6X35q7sNLfJHlqdwxghiWH40ZIGzKjMRhork6APSq5
dCW+XYvT6TnVTvqfcJTOyWa5diTccuZtv6N8Dpu63aLSyU2jgkwapUL8QukM
agWasBHgUxSl26+lUJPZu9fP5ZrpBjSLnb+sjc77Vm5gVkNIzV2De0rX/ZGr
MxltlfprTFDywX7pnOEFRj6U+ZE8kM7mlmXmaO/jhh6xTwSP0oGveWsSaqAC
VPbFM3M1ZeI6mArfZev4ITmBWv9AoKgO8qU2FFxusoeajyHRNHKZ4j1NSRYb
YtHUGllbz9nB5KfyYY2TxrLjFn1fwyO24ElPBNArbURif3LeEtu71BAo7IjZ
HG0VYtQzwMgBYLkMzs757+htoAf78nGxuC5xBXRLc9oZt6pa5vmRqgQ4Ivw+
vSm1C4FFMGnDeD/uH4jWoQn/pLe4LliNdDPNjiC6OHjwN+i9yicyawK0KdBs
tdDPGYkrnVjRww16YnqgiyId1mzwV1tw5Nznm9bxEHUKleoRekWY016ytAyv
Df0NXxPDar6otVFmiMnMYjAesExVv893pUY0YgJ66DQMhIOun+aZTuV2XN9x
GKYhoLSkPUGkLrnkfR5AAC1RtOsU2iwUcAijyE8E3yjQ8rhzQA6/fhIHEdke
YAg6Z8Y6NmzbFClDA5MjyTiXeVJIusx1nCwvtFj4ETtJKoIUw3YS5QerNSQj
BQh1R4rNNfbF9I1TR0dXAU8pCyVX3vlYa8b+gk+M8ascJWAT0FALiehe0NdY
4tvOHmPWKdt+uVe6tnIb3iUwCTs3iK6IK40EzYuJQSIjtSTZMqLpV/VjdFCO
vz5hbh4slvxsEO5glGL1tEzPvSXrz8kqNGh1fRWDDEEq9YMUJTWRDW8MBIsn
hJy+lo0JSyR/HXAzEoMrm31aYld4bdPzY2IO/JqRhdNykt4u7O0ZFprFAYYI
sQF1VTOhQcnqgECXh6nYsgjjYlUomtrn2r+acsPRC+vaSDnNRROf/MTvg6On
KXkv2ma/9MKG6gyVhAiVPrxYTECRtOdFX7TXV1sHlxqIvoc07iFYgphOIEWU
SvkRHFLkXfXAVCgLNC5DhJzVsTmkTPgVEcVi4d3qhr03QlUR4sHeIOF9+zSh
/dNF8TsrimHlncQJ+E5GjCnAFiyPj4wkqVRQtngqpRlRpHdGjWPHkExqp1/R
DnZKt3UhGxj2MgR7Y8kBcMwKP8NY3Qy0Q9tn3isz2K6Y6/vuMMD2KIdfwM6H
eqcUZmdIPWfJXXfYO1PPMGfbJFeE96/Gljfjo3JVnJYxU8s9eby2j/9xX3HW
cW/uP4AjSz0VUEQXD8JDsTmdclI8vmEdUj8sofXssyu1CjgzomC1W/HrY5PX
/5dbtgJpjDxXOYoo5P8kGfFWx7jVq+Vbd88P7psFnL+Rlohixq4FqWC4b9ak
UrrnAGMwi2Q6FCoywIK3gPYckszYNoEgGwTCyX96lTQN3D1WCAzMDM4K2fDR
88rdNKGYkthYa74pm8PIfozsP9NvamN9E7l6cfD1VeXVb+IhTpgTkS1NkHY0
z53D6PUvV62pzTBnUtCrZy8wV5oQURXDUbP3hmeT2nrbTCoPeSfAqo7Z6ssb
sJATYDkTW1Z79CMfkoZDYumAX6Svg4mCotxbXu8YERSBd0v1pnOs83USc0Gq
clawCHrafkwaQ7nMMdNXrhN9IoF2grYmAJbmk2Bl4dBtLiBC32M4gC9T7JqZ
Tt94BfaR/LM6iorpHemXtf9/1rjJdY3Gl1sg9OSKFa1E6w3pO145g3AYXwvi
EqR4PF5iGu5slQrr8vz+SZAJwsjuys4i+SVpnbi5THs+M3aqPboawQya7DHQ
rkqTEPXlyWfbLMGoTUYltAW1y+RQYazRwVHMHUGE2vTo2NVt2rsLLFYVVYnF
7EGxcyaxthVfUVZXD6YEynzu482euB1LhqNRtJkbSCuIdsjm7jUFijXcP70K
tG1TlIAqzlPuQ0dBNiXZwolRvMop2D2oyhOUiZkOuKDhxn8hz2m2Ss+rIv5i
1TnLlLRSO2erfjEUMATdwfOOI6WexETy/yQD2gCPui7AgVjf4PQfoKx7fEkJ
OAKUiaadhLVd6FM1sE7x/sl+0bEyNiNMh5KMh+92J+nLcy4v6ClARUFdWSqa
T4DbYr7JZYOgEA6nfxbrmfrDfWmYgKtHjkraNfBuEm3viPvMhZcJiV7mhFY2
zMWgDfVcHq9hcrrRMa3d2YzwLQ78w9ASyDQ+yXVAjCxaJVkD+mwj2LZVcBQU
/2U1x9/0ARP13+2MqHs+Qdnu2PQLYevmPCa9Q8t4QzoWT6MNLPFQQbUjWvAD
3L+IKa8pNZa7+LpTUYunxPIRJ2+/h/Tjr0xbFUlCfoYV0kZ8l8BChrn1CYYR
Ixjn3dzVed7ui8b+UZYqOwfgO2RkSrYxZQRndKfjRnTdqlJ6HYT/EV1Lm8G8
zh9xd4xiiNQx0n/K78JsCAMqkNeLLhKT16hhPkd+ly9/fMBToVx84bKIlRw2
pnkolNeQ3BfxJNuPUrjQckaS0crBEFVNXh+nseOsriUxiae5X6lp1wbDVfZr
ZjsfJF2Uz/fGn6KszQspPxCRDokUTPoSET0izvYXsIfbrM89xrbQ4ErgiXK1
AXFgkr+to1NLUk9OUQAgL5qFvXeP2trwK/tjiBQ9yqdwXD/k9EWqp99nZ9cb
FCDHRcAQzuJ5nOpDnz3Z7jofjHHqIlfGehuGU5g990GWmmSIZ9sCj8lgvwq9
uaexqivZRz2oaWBusfKGBAw/0IqosXjQXslfm/E3j6p9PQ0psK11auBhIV3N
6c8ldc/smSzvTY9m+wzbISmNRTXzccotIG/p01+06wIAxFpNzaixcwfaiy7P
XQ2jKSD+17z/K7yWmIwjMAMXVnKseY9Ii40CcgZ/B92SAoxy7RrlI0W7v6yY
wECAVAaqeG8elXKmOI9SLJlcFv3iwi68+Ao0hTG5TKA59jTkJn+LG+kbsY1O
Ljg6OVjf815aBF5RF2NQM+ORgFPJ2kbpkjYT+pvIXxqG+zsw5L6jjeBvTQP5
Dg8YyZdj01eebO+a57VHs+jlleToUIQ0iXZ5cOHnnNjxyEsFZBws0ynOij4H
nUmHeol5zwKvs9+E0Hrx0I1lj3Hl5hNTEWXqq26H0GYXAPSgbVpl55ze9n9q
+7HBGYugdYsmwQMpXntJH6HTQhqr/ckN5kc3sgsiN82WvPOBgjXEcZGg8kof
tV4ej86uCzyfzApivKLbQDb8uQC8y0/ZcJ8hShDGwgrQ6wze9pI5je+5YsSk
vwt9cZL5KHRt/XBdS2+L/G6Oh12d5F8CvXE0xRNOIZNGD+iZxI0KGmbCr+DS
QCZpyTlX97Pc2+HCg8qmzV/IbSrpJMavIGR2hYqLbG5v9PmjiguxQaQ3ZvzY
LRvUaYV0RD6enS0fEg+hZ7yF/xeSkNHRxRGrd4MV77bQuWt35DrBtClmrtSi
0w3eGERXk+XWh1i4UUh1SaBygmNqpWM0/AvofBHvxEGRjK6TKvcig3P1ylgn
3kpgAGi0NDxI+ZHBlWjcnLxyhisbwEZcHVAomLTSG7wLlVf0DY+dcPqGxDhp
kLRA98i/H3b2aGHAUKPaRZpYBJhiobpwKSnIndnL6hnLwXsA6KYSHdLDPClq
ZB+JbE7lxAAB+kdftAP8TlhyxPtMD15lLsKnxTBXeYm1G/UT2KJWW6Dzne0B
joBXnCGDYqk2tBVGIPeAZO4V37xP52PXIhLBfd4gYN/qs0jJ/mLvaS3dAXBL
6gjASSzwrWdtNCqbfHcH4KMB9WAVAaavUnuUTrhit9LBBbaicTJyI8coaaYJ
a1I9HQyFxapdZ58PbwGWthzXZ3qkoYFe72Qf9wZB9agZ5u0RjQUnRubBf1rj
HxTawOz9xIhs51p1uDjlyW5Y7g1wDOHgB3UW9iV9qkkWwB1PMQ5ruhO3vczM
VGT/QY+Kf/oVF9QtZ7TwlFCIaCfBKZC5y8cBBc6s/cEZ29SFSgTUATH3L8bo
anJRQtETHPUSAZwFoesy2qB+IS2E6/IrtCRhJqFqMR0rQslzkwkxdVG9k2+W
Utq107XaIA8t57sN1gkIzsXaJM5D0rcT0HnK7owHeLcEBymrB1nQnqaPoxoN
DDkaUORn3zQM1vpkuthXi6keVs9hEYO4hI/S8jes0fxYFwqjug1dmnPPGPa5
BnHSwVTyoadr3TG53S+EVAw5q/XOywvIzrvV+GFFy8TqJZVE5Hhdfj1PnJlT
EVMDx8Q4R/0evRFSVpC0JiKMmIev6MNg8jYRtcTW/91/18I7aevm5JIOkUF0
73gdhVY0vbvbIg27Mj0NeBjVwKLUlpAyTIQzgMySn9YOVmUWapTxl02wEM/s
GZwR1tM9loR1Vj1dLKtcxKN0z1NaiWRhWavlaD7TUYPvfP/yoTMDt8yByYKn
Ka3CBU6WHbCILM9cEhtC1j1iCCvFGRDM+2DSuYuurXcrihsGfSrVb3cUxd2F
XMp9wDT/cZKKzALylpt6VmauL6t3LRe7JW1iTcSle4ApVqEm/zDYZRoofA7M
nKBc/8HOiz11LT36TqUezYe6AUSX0MUgTxEBsRTwDaoZ/RCWwLIsqGhv+PJ9
4R+wQI+dDM/TahO+0W3IX7RcuAMYSPgyqzDNFwva7ghCMymW8c8QAZH0C+jd
n0EUTM7p1ljEgCJoQYqq0kc+Kiie8aacSPw6HzwjTga1+y9yfpA9dB0Kt7VQ
kAj+MnZKCCTFF5tkTurTPIjylDp7Y/0EpNR/sXHLSINEzBQHiuehvAb5+HXm
m76CubmTkJ1zZ+vftGx2U75/QqrXlZrJD8iJztzn0xAmGQryP/GPkvRF8cb1
tpJ1c6RLzoKoMWP+FO0eQknvxWbVLTqHpC1liHq0hWbkRtTgq4k/JPB4ivzz
yNFZ556ToMJRVVHaCVTeHP+ZpiivkCT6F2+6oM0qRMj1nSiw9HoQXX7+5Hr8
nT0tl5EDh/NU1c/W9dq67/tLeYqsY6VVpz6uCCduqCy0/D8mbVpD+kJIy889
hwSlfEVu8e9JQiwsuLLBZm0NvdS4KvqWYxjPse0wOD9JiAyFwmZWFp+81waK
EanxxCJ3LgAI6Snpq+nFNnVALcIRQzlyiw0ChkY2NdUD6Sva7Zvok8tOQiMR
bPa6An0euEVyGFLCY0csqm6mi1+44WiamROnQIonJeVQqgBse7e26kFlqmto
xeypGUOnq56FspbEH5zTO3zhwMi1mKHxXXiFBasFOvj1WVdAsZ4m27ctymNs
9rQqvYmzKa+lHs/LY76RCYvfSjofTnN2zLBQOmtdr1Rc9jMtk8OJh6eGStyt
1qVmoCaUY/SeH0jYpqPSbt6cdCWprmi1NIlcOAurs3nb/9G1XzjY3JoljYRV
okjTVC/+jIK8Xdp793xYe7sxssm3tW+Ui/8n3ESiVvX2cTImM6xLVuNiIw4H
67FWXfoIpb0LbK4auZpAVH8c3MmPpSCPjDoew896R43pm4ZrOYWt6HVSSl3q
QTRQcL9xmXLQd9jQtke5J6YM9cTRoA13omt4lMIzNIf8vqt4UGbtu3WaVEpq
3JK/gEeqsf0Z7pSx+dxsJ+p/LB4+MGiHnFDVdXrmN/Vd9cisFv5O5upTT96n
aHYPP1V3PDcvwXW/93lmTeQGcjJrv+Nu2selNhaqs79TSBaddoO7/cy+D/Ay
VR+yGZK2Omq4Rjy48hChLdoFCzvowW41sPoGl7n5r+69WLg9Hf0bRz+E1sJQ
HDf8oq9CrbVh27HerdZzah4QzDW9ZPMmZOX40F17RP13lAFKm1yYGEr+xtvy
U1YGyAwhUmkLIeliX9ohl3NMCqHfbVXoHaBUownWwt2I82YPLprwGOO/meXa
Sfk4vd311qWaJWTbTfIJmPBB01B8orGHlUbDKng7P10jf8K+Q31ROzowG7Db
3qKr3i/d4wrrM2Vs9HkqrbHiWqgsaSA5e4IF4NnAjQ0vbUw6jX17D92b1NKj
cKmQYa6GYGjwVUJ4GXIBo2dNIYvk/gX/hh7K18qyMA0J3LfISKVNYfY7mHeA
WuD6X7UaOPnBG0GXMCWtbVS6/cMgBKgeyj8pVhXFZLsx0Vm1XIu4Su5j7Bz1
XE0XGQneg6CS/l54PbVGksLPPd3HVpRqUiReNTtNH33dhZLdSm4RHvQZgAnl
VCK/IQVxtr97B1ssr6YNu3h9/6ZG+ZZyIBa5ULEagr97CJX8sxy1QEdf2htG
p2vLkTAq1AHlCf1Ii1CxIHIlNZRipgxYvhLZ/mYQ63NtYwT+Rw/RjC4PW3Nr
pJtfOzzCpcPnFTkfd2FNMB2EoWl3zw8WQS6cGhVs0qtIEWT+aIlvRAB7+vpF
A9z0P29q96v6x5SzaZzVlAd7NCzoILbnfsmMbRXqyzRGPeYuRjhJD2HAIBTQ
e6s52SkYXTkZk76E1z4ATF0ELx1RM4wFv+ywU9qYTEbL+HYX6HuQzM2x25td
6iSYZNbRH60hf8I43gBHRlh9lnLkMB9bGJzAYtoS1xVRpTd0zT0WDZXX1zds
LwhDiVpRuIEnouprEriZsjK0hlo3SZrpv/i7Hnw//hab0/fNTMg3BWd59aIY
QmEQ+4aRUCbynus1FEJCsu125D1TrjLaB2C7SHGNIoPMfQ188aSThoujP8b0
ykGKrzrj8odttKf2kKxi74/0bXMoKF0Pg75eo+1l80zVaeEQwM9gP0U7CAoS
pIQZPGSZllWMS5v3X9D1lfdn8pfkq2K/WFIwRyQlGiFqXho4zm6V74fSy19B
gyzSjW7g0x+94HAGnMXm80qbMjk8j8cJrxRa6M2EwMadoqb8WxNmkqFB68Dj
6/2NruZO9XZvsPnIsW8O3HZ+bwjODJVvwQoQy1mfFVq26+Cjx+Cmfw0a+SRJ
245dk7dccQccEQANupaVMKXTw2XTHDGxSvu5+RftjRFxVRvRnRLEhKzgbBWc
4rI+5CEdL+UXQfatMDIbTaRDkK3kBm73UmXdQTajLQAB8qooPkpCKKoY2eFQ
KyDjen1t53gOSDrwEbBWTCw+omm1IJTUP46Nx/d6X9k6+E+nF5QM/K1/jSwq
wJrTKq8ALPOQM86oXYwArjeF3BEPNhbv3ifQeZBmXBLSo2Wiu8RJzPcAhdHG
+0egi2YKCp7kzxO155CHElL5odTeJpD5tWnpOqLLVjIo08WzCL8rToy4G84O
VRYReUwR8vOdEvXpuHPwJ67jnu3kGeQIdIsD9USVhI6imkG2sZNBVsyHkx9r
w9IxioyDSB2n8c3PUnc2WtqQKB50cJy8WBok5x5bkQyhlnYtm/j7MONVDBET
3xnKdKlxN5j2UhN3wFd/2AiV14EGon+ivV+Q/PhRwzJmv0yU/gDJsQqGoiql
ANWGxjF7tKcR/8X64SE7KNK3N25u3iGEYnDf8SfQWYUZkbvjC89J3VsuMM6c
vVRBr6WnOvc7CS8wTbknT7P5V+r00vkiB8iGA8AziB4N8bOXTBBX+yG8MgrA
2yl6vQrIzZJfeaAn5yfQL1Tu5sDxWu+t1I3SsFpdTL0yy06lmGqnOnEVYIIg
FVL5OGcoaSTPWZmZZCM7NGJeyFOH03o2TsOFEfv2iXIq2cT/HqlV2L/3Uyyc
ZdmJQd9A08gV9oc42FHzm6CileplMJmV6gd+qiXS3/8CHsJakDB05D1grGXj
9iB418osRSn2uXTK2t0My29O4BxKtxY6P+4B4jTxrwbXTKE5tOPxioVR7IML
Ka6I9bsbA2m+ntPSJ90w2d/7tUD3/NkqBph7CEHa3mlJ+iM3Pt9ljmtusp1o
J8bLzwXsuknjyI+h3SYMzkXNxfxQgYE8UUaqMzU+3vORybxy7ITXrOo6W4mY
2zQAYqp42keyt41ADtbkpx8cslpJNbRh8kydF4iekB404ROEz4SbI9AX7wmf
ffmVh1kWAa7hXy4uCv49TtzXiUTUDluqOcRgrue2jzz/mQo0vU7JXTWkPujd
7eR/fdMEOjs8ulDsEHvmm9SHeE64KqVUzrsshO5/f//3zluNwpO9OcebT5CZ
usmmaX1CCRUwLMCRlellPZdHgqQTcVa2yf8+fTQYoziBwe4HZzXSjAqccTIu
YX5aaDxfXDjQAG+0RPwMBgFhC6JI6Bj9HMVpGuw5emDHaQco0Y7IYSBbYIqS
dt5+OjufimUe3oriuoVGmW3/toBe+RW1d9fPcppKcdycWE4JuFaog9LpmDu2
dIo/qc2sWPiYEIz0xX8l5UZLlEkmNp9+Y73zmh0GpAAjXtbJwyt0KdVPy+Dw
Liv2nA/VTuU1Uxr+SvS+/XMU3cb8Jm5XaCYHdARoaNOgdIVOFXbhKjv0u42R
Pp9pxgPU9g7vxEpokmTv3w19OYzJoGW7KM6UPTLYkTUu6ceiWasc+6O9f5+3
j73E+BxgFX0QKNCmC10qqID+UbXf21e6qp9U8eDOf6enoGYiulgJbqfKmnYp
jV8UWSymWRa/JI3KG1GQrfp9MEt9e6xZ7CiKQrD9PuVU4pVAvYSVflOxZjk9
k4TX5O6Q4YK3LmUws+qlfjtklt6w+bqsAbGAE5hrCKTkVRPU4K9n6TN/2lLj
lekeQNHH3pbHNMcahINch6U8q6AUdX3UJgfYwKHDu4hTPqtBBYI5Mu98S3sQ
TAhQzPYrKLclN902zsC132emvTbOx+E5GNEEeq9bzyoTmRiiTS4gIwIWZFff
4d8EfElaM/7ckYspWsLSWO8nUsjXYh+E0tCZu0Sk6CfCkx47dJxIw+VaHytC
GKu0fhZVrDV1ElXGbf7822Nk4sLVyf5CYU8nS9eE9/0BUYDzwEfjSo4feF2K
8B0qeCkdy5Ek6InYWPwH74AAXmWY5vwjrGQmemTdbHWaKo3Gh3ULPn12OXZw
PELI5+gSsazD9uJpo8RxU2xOBD9nbFOHXB4sh7BHyExE5zseeghjX7cVbAtf
cSb5qHDHdQSHOI6PE2pg4s3M95F+zmmaflW8xZwf9OudQ9V/P376NqCf4C7l
an7Lw0m33u6ggHl2nqgK7N6T7SRtCnre93PPoJ2iyHkNORq636PU7ti4nhf7
v6BrYFex4Cj7DpZ+UoYFTrxCORfiVZ2IF4TTc7Fi72cQ6CvUSDrnmg4TJZYc
2iOhtPRemK3EBoUKkkedwZRM9N4ZIXNbNrt0qE+C3gkkhmWXaAHWwjCiiXBY
b44lVlP3r7V1JIwIFJTTXUutW76n4KeFukOHfwZyIyYecTiDdm7zSL1tpPUU
fExEW9mHCs7WUF/bW2Y7Xq1IYqnIbkEQXiWZ537Vh/mkpmcXzl5lbZxsivjC
oeMqz/8sG3/xlt1vN9FfXWQ+R7yu3uEpn4EO8rz87JzMilxNzGZSx3IdGeSA
05efwCLBE3ib+GLtCQn6kvjsKNYLKQISU/Cp6puquBAhcuBJtSzWrs3K5mJa
CC5Kpiqh/YI8g7xsRy1fI05HYEgvrkYdz4mroKKbh78txF7ju3wZiW4LEzL7
SxZhDko5dBSJlXle3cArkIgwpJYHzb7YhgYlOMowU3SN74Wj8zDUM4mJPACL
CaeqyQZrJj9iX+TI/9z/Hh3YH/P0rPjSGpoMBUcmoXfUu82ZNVyuAtsPP/TV
ow+wJUN5HdT6zTICAuV6u/PuapcQgSNVE1RbxLk1oeeKDISaW6JTMMMOA/st
PrZLr1Y/TIOtX26wg5agk1EQ722dLv174w7RWq6gJTYfppSPwLnHu0CDfNGs
X39wFO6vLmvTf6Z9+Zb9RKmNw85q/6dXDPwi2bK/O+EP74xvweLfOa3V7+24
hcrnQH6FV93XNFOHOuJNi+d7Ohl9SHlgjyLAW8FSCsyntUFxul76BWuraJJ7
j84q3+mzoc3acJfIvSTpkDCLe9PyU71T+biC8s9kkKkzgTmfTDAS5D9lZrG5
UvIx35VupDW/DBNbJxxl2qD9G/KflzOcx26pDQGFjXsptBbCFZm4m1Wt8+I8
Yg6Cb2gBeBXLgYl6aib5TRTU3TqRKrSbbSd5oHzbgat+nBDDWrR6rqDS/Gdd
RgW8b8bgXcTjgpQEaQtFTnqwtHJ4Df/3QSeYpPtCvt6DVPjShGDQhsPHe4tp
W1HSqoup2z0uB7BrRdUqQiCdUY5wpFJvrQwtnen4uzMR8uBlSM3fB3CcjriQ
HzNoG541GidcPYMpLneQAPf+Wa+Y6aPTin8ErqHxgFJdwvJUrHCeVuop69lf
bhQRQyMBmiLJNN+VzzskiCFxlKR/uA5Mayb1CWPfA1NxwAtcn6s00CJGi29d
yP9Ab16zTSWtOPh+fbq3/YcBmeIAjlGyFwsiWZuertWcMPZXXZIdYPQALKs2
6l86fq3QbMiRq5es9KjRUiVX4EtsFAjAvP3lKlJ+JU5ylLuOlnLVzUpCkmd5
tj2NFD3xV4bhyxWWL679OJBws1n53ng/4rw9Va0CgaoOfWmlW5kIkiATkIfV
AeGijQvcfuDRZ/66imFmeNXE1mjI7Q7sBxg2v+q8RBaAG0TOwSGLp+Lhhdme
87zq+8M5TLz7WOu5GcU1tehcN+etWOPX26GMXjPSRRftA7KnGLXqGv/aR60j
QZ1wZWwwANL31FjXcti26k+upDDUejf7dOd11TTILaLhXT64CK0C1PkMT08G
rE1K0LcG7hmfBLjCYUxC6f7zUONdufNXJt+FXkqtasbB2rkEP3ZHXsqmAWB/
cjVAYR67jFCpACQvTmTMEbnOLj01MupNZFSaE9MuHvtpxahYAyo+p4JGR4+6
whoTa0KI/K+fcCugm8pJYSDhwU9PpATcZ7gWXN3x4a3UHVbyPsVUkk1/M2gx
74xOK9rn08PYmWHrHWGo1eWWT3+3t/prE9/P/cxTIr8j/3CNuVk4FEkWjGQP
p0pUhf2NG8Ag2ZWEevmLJZspdBmcw2LmLgg/XYFjP3BYiVNFfceJwvAhpm3k
kAJDjoHcmAlQICtZCLsZ9zfn3JuPbMQNgZFJNYdjp3cFGtFXJu0lwPcW87rg
wHj1UaTdGtagw04l9z4u3QcEEN/iLCDk9PR6ByobhkK29DJcfxngNoCXqDCo
4HlTs4rg4iAgnBaaz2GI7hAb1e5QK158Ct2P7eNETbKtTSTP4gFsB02oMvi9
hDqFUXSnx230VvNk6safVpLODBvj3b/BBhRowgQdfIULvv7UNTMc0dqR5+LN
MQJqnpoX00pwmuVkoDW3YPHBBXfTzyFsA9fs83uJlDVny9jEPlaj7CJkZo+n
/fAmYLCg3W3NYHb7kLTYKMIoPWUckFKjakbs6/bxvWGeRTdHWmmh1bCiM1CV
U29CdMVupuEegCLWxZDmccNbFCkVvWTcyaytwBccHNGesnHvarhmqnH6xIfu
MN/RxuWogLZoqT/ngByt5Gosy6gFdCLGP54i985hoUKnfOZm3ZbLmppBW7gp
M3AcUh8mabtRSUgLwkOtnSUxZqcyn91qLw1y+13pAb50LrWNeihK600JEF84
wf73csH68VJbrUOsqFmG9qjFr/6L/7Nnswd9PUMKjvJBwFqGYKqUqnzegv9L
4IOm0TRdEk+A/ZZmlp9Xg5zMBwksnyl0/z9e8tWbOLIr4mvChTsRvlXgAoZl
kYLcJ93CBduvJRWW4ryckaxnQTPYLS/qKv0MJwt8YpZZQd1xbFHMhGdscNCN
UVtuHq+XAGMYGfxnzs2EBESctnWy49pNy+i91YjMPOYbKLRq6u7/bxD/xfaL
PRzbvkYHxhvnogGXW2DfW3WwJKvbcHTiVP9uctt5VTa7JdNw5+6TBaAdLkAG
w0cFZxzfCsKaP9ZGBbBOhHa3kREg42VNyffwVKPNMQ97onJOcnr8Bfm+FC8/
uk1Z2khRUVIEzteacPqcT0U98tb7Df7mHlIfN3j23L6+5H4KoFfWLXvMyDT1
jBrrJrQw0zb9YNgnwEK+Gb8tYn9acPOWHkdbtcfsuuEfZ1I7JY/iHimS2Dmt
+oNlkwsHeXomPib1FCALW/TO3Lv6b5Gup1h+hXe0SmUMF1bwa1lnRh60Up1E
SORh+BRdnpKOLceAxFTb/AJyKxCgmZpt8J/bBzR4WS6rONn6S1YDWiFJDk9E
GcrotYLqugprCNGnjGQbMZWf1SlKgiTJGr0oDBA8hggYT933UDRc0yHEapwN
r/wcULnwjVUhGfiKgaWM1AGEy+tW1zvZC7XiRAMINZquesfCVOAiCpF0cKis
DP+LXhxVFFDE7wxOCvplhmn5FEj2VwRGGoCPD/ndUIjMKh9elS7/A308cE/l
gk3Q5w3OACvjaG80cemeuhdlViue/yggjgBrQOQC+KdlM891ICw3RRlzbinq
QgCFQFpSKiRlhHkS3wDhkU3nVdxgapHTHKFN6bFa+F/4ML7myBMwBMvkiDs0
iCZf0Sc95NoHMQkMYPxa+HTYE6+5lzoSU1JoB2sgRI9OH8mHhgAGhNKgw1zR
FC0fiB39eDsFjSnbwRpet8L2D7PltaWeMVdVoyYejxGiU9mnVp+zLYWwMXXk
oNc1z/DDHVHTAW3J9mJPqiJNzkH3rjcer32nMpMLJ85MGOCeKb1HdVEdLsgC
YnDUE5QxYR7UZg/5EvqEAD62QvdOl5zED6poNWppE4ebGP3rQFGoyp458jlk
nvXCpKIPIjPeY6pHv0MLY7lgazHcxjDwPGMs0GFdJd2YMLMm6LJsi4TYKHk+
6yg7fl19xiXcSIq8BtslqnKCqyxgIOPun4CVDQ8ryIrUVNjnPOIVBbbaVrCF
glMKWrpFe3M0CMpQbzNxWUX3XMAPkUJUvvHoidYAq4GuswuLFMrC4p6hgIrM
LQ4TQg8o0FRhTQOwuEK8wXPcSRAC/SqKHBhSSnpZkorgwYsOko5UP+SgumHw
QvoBxGXGcj597eIhxQnpdahOvq6UpXB9rD4A0jdD3mV7P1Xrugb02+ap+MZU
tngD7VS0eicB1DY+W3mfJGTyCxkpmtxuuPLxd81rmxk1fqJHbWJJ3v+Pt5ra
VdlTND9+Guo0z8TlXIfKh641mwfXiAS42eA3BdnIg+cTSPyt4HPMpzqoas82
C6PYVXxfoJeC4jAuNSKrQcMFC4ZVTJO33LDtupkVkw1SiETs+4hVqeCIO80J
orNdR64UPNmWjpHa13jQ6bT4Bargt3Ll9dmUO3yxRQiRzXWW3vlJeg5zmwA8
fA2OPzyV+oyo0rFotY4x3FcA2erxGQmq30JrGkhIQNnz1O7fplNOfvTsfOe6
RAiJw1o8+v7j85zmFEI7biSVbZK0vbZjTVkSnwledPp/Vqm9B90WYRJh3wgh
mB48B4vWlEnU7kYy91IXvF32xrcUkA2oSv/9cpbvuUDW/nRtrAoyTlUtTF+z
6PFFk6sYgA/9ki0wz3iX/7SX9ti3s2oayAp9VrfUhQbnwpAiE2gJxpEdYU9u
EPV9xO1HUfbCGVADLTcYxlHQADiFvmiJq+9LIBQjQJwNOaq8wrWGinzi3kh5
ohv8JV6/HAMwEx3oHNvT0xXy/RmDLG17Zo1xHztO3+hClP+1yVzlnf+y0rfF
yPr4X7QbZNUV+/k/S6PfknN3idveycbRGQoUpaQCqTlXjDFJJxL7YIw2cZZm
Cv42acstY1WU9nMkRhfi53H4r8kZemAQ5C3Rqh20l02Po3o7MAxT22e7ocUH
Djjo/rOlxNFXSLM/Z4B/Q8YGcc5tGpuAw2uJxxJqQlMmsckrIwJsYtIELczX
joQHqzUmqvGNWU9phut/TPS0h5xRWVrbtYoxMHnN6jd8q89uWYIGUdVaznpS
KpbJhyvEVtoceRDSA5ULBfddsFOZOLIYt5bmnTne2cvt7EQpWV9qFSUWPXVT
hY5gXD7VzPCDnUF5wcB8wOyu1YGPNyNpC4ZZbCiPzRPc1jX/A9bii7DMLzq8
9ueuB28yYQbbR9al8gze/rgiJJ2YC4aTVkxEoHyOqovydaj8R8c6F0IVBWDT
gAcJVl09hmUt/BQG4o2Wj7RhSzQOJ4pbPhfjLN0eOl9Q+dbqs/4iv87+VmvJ
fs5VPfi3kncMpCFSkw8TVlgwz7KYcAaej0HeO0zSeKTFLbeGyFG76a8xXUsu
31zGG/hIcHnbUb6/9v35qHVNRugLofrnpToykhNvfhH2Xd4aeqbg6ZMaJlA/
ED8VFQIRolQvQEb2yOKdZsvRKfHRlNQFSRSXk0e3vzWTJZ2/nUYfKyqAxdOc
Y1tXr5hhpJtKSgi2CbbVtK56YcaJvNxaRaiIrO0h33rtIIIC8Vt9hlX9xKo2
O07oSj8/0JSFs5O184NnVpsHID7GE3JpDwWdB7jqFKGIcoJUIgfAfEj3qnk5
FdgQedR+/oRsHbtiuyFlgg2dLhsKPVk2owjgLaqmuKTmZVpl3NYzIJlNsASj
tF9a1HOw8t+wSi3IPScVMzn3Y3iWWtgKSBjMbFitEy13aA3Wy686OdePso/6
3ucz22B8ACbTsRioq8X8JAeTSr3QlJnXPhVSReLwxVTqVZ5G8N9i+6ns6rl5
gBNt6dgy1f8RbssJ+G4aKp0XQDokhnCLr/F5E3bfWgdyjPxnILdhGW0AYJWT
IxDPaUXLwmrwVuDk9/Ks0YJitkpQnoH8nc/FkEyZJFNJiaHI4Pr10OZClbq4
TzWcAeffNG4yzX4Rzh16aAIBxPyN/GsvY+i/4JjNSivulq480/7dxOnXpi2A
atb+/FNxDs88CLP4RLs83FAcpJMSVaDPO4UwwZ2gUdiNY9IlABaXpN62Exuj
e6tgmUyP/6ovO2DKGUqm4qqY1pQMtAGl5cuqsIftuvAcw2+axxj03POVp4dJ
IJIr2VqR8MR9rUw4h7W5zb/sqzCHz2I68he8dhLIQ0suy+r7g80vty4jD3+R
ozpxWoSrtZgTSSyClNN5hAYio3n08i8neLfAMFDzOGmRgu32+cB3jyUjuR8u
pExbzCmYubQh7NKp+lJahxA759mLjOJ5rb46ijWl7ZC9rc+QcIzpweHYu/Y5
1Nd6qhDc4qV22rw8O6lSynd8WJ+0W8tErgEAIDnkqbfD/kn5wvYGfGfmZvaw
joUYdIgNCxM618dI5yS9wOp+ny1HO/GnZKV1vAzf8AYypXtoQNnJHcfs2mY2
GEXy3yWL0mj2Rj8rGCEzeLugtYtvR1MuRwGQg1wk8Y6cbWMecf5ifH0SfxwL
e8LGFu1NeXWedlvOaWgPKBYl2x3/Ci8QgOkWdjG3bjakCMUqoUrly5+DYaF0
M+bh/aOCGDhivlpLXMrJ365k3iYOh6SB8cf0tW5WNeWenAf3rhT3B4hhBTjY
Cfup8UDKtDcyJzdzn6j0dNZUiRwkptYYQd5Tv5EMCtVQ0y95r+ITAz3LpaE7
/vo0awHG1Ku8eRlrAUs1ffzpQtS8/V4Qs4W/EphhHd8E4FldNgJmEtcGMCHL
cYE8fXSwjoMr0Vws5mc7VTlliMYdmnfNTdUmgav/qz2F7atE6xj0atrgZOX9
ENmZ+Xjv0rKXReL5hxz7mWYhX0elzk16cYwJVxJNy1GXrrHqB8QtZqvOMciy
dmbzHWbZA6ldzJ5AFEkNTRtgyAe+QkTZswELpSj44xmxLuEYZSJMyvaQF4tA
snqWvTCU8aGFh92Ni/apWEHrdBT0ta5HJHj+yf3ZAvOr/jndQFOB/ZNzYkzs
UOii10RuNDcPyNthrdhHFcj6+xAEFromi2Di8vU1cxUQvFVeW82xKIi/p0mq
YXdOnaEynAkXUBbtoIKr7r/JCH03uHgueHcMeAUER7sgDR6OvNxEQoWbfOu9
Vs1zzjbH+RkO7/LYAC3zxjwWxCDmqAtinetf6cTxs6Lgjp0p5J70fBLVo440
+q/4LhE+cKLgh+yUrhUIAlGqR7m8yoRKEXk8vSHL1pQHTbZGlN0lecbNsVz7
dYjh0HpAhizByPpdfZn3GmqW2n8sWFlwvl4f2zzPUAJ4fjyfQN22bAbzqJrv
NC8F91Jld61xcCgHICI4XfCVp3tYr3lhvc7ylwu346RJQplJYnuOqCeU0qcS
xa1pkPWCoGxgQ5nnGtIOv0q1GKqU4M1/QpRGBWtfF9pND3JvPVhSs5mDbK1U
ndsXm1ziUadzDfi99bpjmOzo8EzT3QQ2tSyhbVNy9GG2h772dg/HSdSYIdWk
QIHvBgg5Ak2/aNwLEeLtJo0VM5ZMp/tNVTonY8N2v97UKfsnI1Z6aLJ6WhlG
Mva5+jT0cc2UO5jIP08HuTtmOwY7zeumgtHttzfUt85KUfFG6e7lO6rcTX+B
Kvog6txBCqDKTC09kPm9SLy/TK1n9G5CUaBm4xQA1A12F2ngvE1LDHLGVK84
W4qjDbbKLBs/5giXZ6Q5S9VLapoXcVuX+IWvbLn1M8Wg7QnyLn3pdpcrz9r/
IJXZWra05u8ufYh2pitloAzElhxWBtt7Z9BQZirteQXSj2DR6ev0qV0PmP0D
jFVf9MwjhOem4bnxQGdNTxvXW8cP1KfOpIjN7XrgMO45n5Jf7nrsty0NnGTC
KxeC0zYDmeBmFayCZ8MT0BrRHm/wnpbc1qHbxeHRU5cj/S3NJiU7FhicLzOd
fbz2LSUvrQ2KU9tZ/BS3j1KLi/nCGJZ3iuzpam2C8Ed4Z49TEE0EGx1fp3dS
jMN2osAE1hwyXGsM2smPkMuc+ZTuhuTaZ1VZHRONLGCPN4e0WB2D/z28n/9a
SLHAoGjExLdFyNXm9QryprzFlSWZrJW+w/XIu7xHEixC8vc7nC5IxYyhonuN
lyZt9rQcIgN1rVzKpz4ogwVprY5Vr/me7+bktGQnfYH4xYayD0O3s3tnvVWL
CTTTtf5Puwvfw35K6gMLH+YCZWirBGe+Dna3DVvTrC6/REV1PpXGVzlxOm8C
5oksT4+P9KsokYyWfIWBFm0czP82K1712qT1Fh1d8CZOn2YYSjVTY6ukYdZq
jS1BnjSqFH7G9AZzQbwkN57qKNKMD/a2gy2boACnZfDjIhGfdYSEo1HQlkcJ
R06JLJUK2uIJnEgDF5a9efSGaHEzxA1zXnqSzJuAmr7rhAT3xLdhXi83TPOI
tsqdcy5xkzAgSd81qiiRPOtC/rnUjMk9lYQlkYgjvC5p8UNYSTAaRkk2oQ6Z
Ydmlm+8zjyUyBMZIF9kQIg6zubT70NsB20rz6+7NdCi0hBYeqL4E3jW9Ijm+
OmaCBDVNDfLWY62UUHcnv1chHTD+1VrK2V3eSsdewSvtizE5oaLUgwwoBMEp
/XB/v1gRrX33BieLNDEcpy2deVK7sEyT9ydmEys27j9rsMcJRdTqni/Si9w5
isf0/PVXL4GuX3IJD98+swJrtw/KKZDHZD65FoqkraERc63Fsu6gv/p2f7Lj
LCRJqycBTJjLpyyNO9liRWNfeh5k2uQTvdX9Re6N/TnB6PQ0RLKK0rjFdvuO
5weJ0jjwhGTlojeQ9EEtNVUAsLgtXqzTdO7LerDEPIT+5pLbqVG8eidHabHP
xEws2Pi6Po46JwqUQgdYCJ3t1khk/gnKhMX7bmEnVk32X3vvI5l6UwNIBw/I
r7miU79nPkzgRWuOSF/6VN+BOh3ZbK7c8pdPJGcZT2fqncy5euX3vKTeZrml
N4oVe+W3bsM1OwB27arOqAVBVtzc9RoidDmSWkawl+z9Cj7y536AYeto8v2Y
sTItknpMMdRbjuEmG/QTlg4BBlxGXGpOb7543eAQYWCsrJAlLKQ9Zsr5zjqi
gxSWLnnUG7Qiwd3GGGTtUyiVvJKtgzIj7Ltq9OdJ3GY186cT2e/FOQiPY+GU
DXIOw7xVNi0zY15+2ZCywRsopqPPYZ+mUy7Z17SBieDh54HEXDzdPMLt1W6v
DIu5y/bUSLgXK2m6fM5Ny9zafgcyCaIU4mVj8vtosiVSyqa+fdQHwhK6J6lu
RrZejjV+F9POObWk0mH8DleCtBBj5OIqes+udKda5YJWXLXJqQoS4OgCkArT
zuXsYDhtveM6rje3J7wtDS/a4T3yv+zeyRvcjt8i5W9Nc2USZiSM/nXhOlbs
q9MgnJLbM18P1Weu9wY7EG+xdC5UcSL79UIhrQPErnC22vkOAE9O2bSm3OHk
sFbZeE0huh1av7L3wyH8ElUmXLdH3XXvyult5rv5JcFesGUL4AcR72gIMcgh
R73uAbp+d1D8zYu6ZD5r6qFewdU+1miKavik4SpMRBGnErKTjakQp/agE2WD
zcGjzBMNp9vPVdTtA4T7qst7nQa0oyocBVWc4UPxLfx81CZvN/BbAgB1K5sU
3UYBythHOy4Hzpu5i+NX+kmv+dKWm+5YiBtQl3T1ziAPYqH1+GxlHbfz5cui
O1MQ9Segu6MFbnKB3vvrxZy4TgREfXUFMZs4RlTGd3vsw45y88DK3x9Pofsy
z74SN8i9CqsFrH201z1lprFefW79C7KfOAxHR+OFLyzUgq80xcDtoh95v0h5
+gZ1jcBIdDoNFy+fDndQnw1fBQ5n2m9AVXE/7dGzLZ0G+RPHvOljbH52zaz+
dCHtk8KeYnHIvzzoINf0MOrLJPyO0QFKpPwipmlQt4HqLYkbiy/A0GcMRA7c
w+OWlHzu0cjIfLOCrOsmmaE9NnBngvXVgClvNkx3/Gl/5QWRbtIyUPTOg/sF
t1Kx/AFMov2hPeC7BSgzlwYM1r/8Ck/G8pGROTnO9ku+booucBhZR2xTmuI2
snEcO8x8E/zw/nCWC5I0svgy4yk6DBRulqhT4N5kIml2D5mz1VYYBAm8ShnY
7ir8w96qFfzbqyC7X/IpFm2Itg7B3N1ETtLP3c+m11iOBcCFxlmLXXBgIBI5
IRMMw9nUkP9NaIR2lX86Zc+AYuXD7LCC66egUTE8FekDcqMJEC4BHEu393AU
Ts7rfqnU+kILsQT4Zbj/ksE+tftGqLl6D1UkDhFf/KTgnDdu9dDEFuMEzgRN
tX+cwb89FJAADhcL1JJZIl7yf85lsm7jcSiVkVmnS5jZ3BY8i7SXWOZ6Ffks
eenDg2uo/BnKIc/+Kf23+k1ci2EHNKMR0QpWOJsC21IJHCOzwTxk8rnHIzM4
bPbylE2A2bXvU5m/NSw9ajI+gAperwAmghWI5QGm5lC7RR60K6fgdTECTkH1
JgqD/zDVKNt2GdNTTpafAV4FtDlPesmeTL582gELg6andShmglR+kdKrL5ux
skmjwlCmBe0t+o7P4VEY6NKwpDuxvDDryJSNv3YsfIGloPV1wTAjfH1ZzmvX
DZQEnKJR5XITyn4SAXr+0p9LfAUM5RVhlawonktuw0j8QoPYyKQjsYJHFLmx
7HHpWgpcUQxoTv7CnB3qRmHzhaqejijsrxmbbtEhhjiZTkVZ39mDKjiujGxV
1m9eu44YccXITVxwgkWI04ygnTirwq7RnCz9izukI0fd9xPNCuWQL8OcYjtU
L1zIRfXoK24hVT6q5IGY1RnkPNmVT2wlOSJOzPYjzUgctuPldQ0lbDvQOfi2
SKnvyHTZ8Fck7JlBSBEc01ZJeOHBlxrAANWYoZ9H+JYSOoOueAK7ZRqNo5Dy
TlN/A5Ia1TkXdiaywdGG+U3EhyeStyCUrzJRLpSBp5/4xeAzgcnVuHXL8ghr
d9nQ3FCSlhY+dt05XZpdaJGaDX07KLWw6Gj0DFoQQ8l9/gYGKKw6TeO0spim
kH+n8xY/EjlDCCLOhKR023fxhNoT4gk0u44QQSvmjyDF01QKUgLw6CwWFR1D
EmTzRXxsiqPeJkOpArY6yn6cWb+ZDsBuZzosum/br0FCMemCfmxR8Zto3fzB
RXaJoc2GbU3vUaQUpfhmQfDoZUMAD1Shru4IiZDaV3yvcsX3Fgl68pVK/I16
mklzJPWDMzFEJVaoNC+huOKYL4TEjVxhgrT0okEtH1B7Wu7hqnjsC1pB5/Sg
AqQZjUjfHrwB8HFYp1mfXBdKeuaST4ps+UkJwrt6K9JILXMVkVHx2+tHeGtA
APq9NSo+EQIp2IYLSfPVYajuMDiVilbkpZH0Oxviu+gs230zsCmKYEN06SKR
VoL6HTLmJAqH6bK7jG6jUNfnFtRH4WWq2sKhjFpz7B3+wmjpKqP24F78G/na
VlnLu5zCsSWwnfGhXv3ak1oCn7PBk2PcLtkGXv9AKqNFAxfdO82BzuD1u0+K
kunqLXvlm6O1669+9wM/4zrKNXlOMeQSFymg804SHm3B7pIJMuv/n5WuoVF7
WZr0rTIkOzPXtEX3LhrpIwtu0n2MYOkNLzH7SDZ0tFM99MLuqjdV0gXtEl24
AoINA8cShSJrQpGIWPuMoSaI0QpC5dORuvWO9srSJs1dGkjkTgkgsC/FKodV
3XRg21+Axrh9lZvl3i0N7YGQrxrQ7ZuEu0b48WVyDWgiQF9N3Ocfkew9kwzV
RV27UqpJMTQzjeZ/qH6EI/znL5r5GJWW96aPOpY4Wk1Xu+rffWWrH/MBd3B3
C4WdU7ynwJeTdhpRRGVfiKD3mYZONuPWUgKfUoirasm9v19cKA9aiCDb6bHm
Vl0D46ESgBwv5Q1AjyjzJese6r4SAkoD32bANopczcpxBiI5OPZ/PEWEC7ar
deo5cbkVDHgiGQdpDnyFZEfu2oEV1YO2DeUhM9iKaeNYvL197eeINUgfFrJt
xszIl8ebzKNd+hTgP51BnMkjbOr/p8FFWkeq5164vT1VWaft5M5OrfA40xQh
vJLrtc19vsV0VgGaeEuJad0mg1NfAF+iLaeqrVs7ZZooXwuL5Ymvs6+fz609
S44z6g4z/Rp3vDnS9pbA52ZLPhtzfTvAKS4SvMFO9eg4VrxlgABOVHTRkYBs
yikz5cnpou/PIFF4mnsHTDSDfzrTEvqiwaKTx9V3RpJujZep5x9V4CHbS1Jk
EgWVzn2Q79vuCbwwBBD8/IznsrBihtxg+RbAcnUkrHE6twfRRbVHH0D/yRMa
atL6GzXtOdwpM8h8+2BYAortDg45rtwgN2dTft0XYZjV3InU9csmNEAyVMGm
VU053YjsZFqBHqAYhnayV3HHNmTkV7uLQhENrJr3fFOUCLt82PE7BMOUPoiB
kLPj8xEa2rKMOSUu9zDB7mXhrNHnrUtVFeHzfO4Gy7hErMfqq6q7d6Kzh45h
dv/jhFiea7lYbf/NfIncZCgzysCY3bPah4NTOAwiUcHIVYNDP6XTtRZFxRAA
lzTugKPASnnm3ZP1L/0OZuKkMPxH75c8hii4dVn7Ypv4IHDcH9U7Gkp1k6gk
tAPkhfYsv1e4rwKUlrCvWNQR0awc4oM2easzfZ4dZlLG3X6mEehJWL35GQdF
h2AvqrttcC8EDtD0zvcfB9ul+UGvpAQONF8AUpd3LVy2Igz19QO2e/r70+yJ
rXjeC8BuuXkNxv/Ay0hYQQQdfeaVHq3rGSK9dlsA9SS6vWrUeCy9NXHJch1M
o3x8wjIEmOpo5OFdMhIaE2EOOKvU8EknD6fODYvqfHuoLZm3uYqGo2clOE+C
E4DRioy4A8IOJPMgxsha4/50qvw56h9xcgZuUwg+XNJNshLsp/91oL8fVdnu
YZnq1LkRh5aQhQ8Cyn+1nSftNUDzVSpCG8ouvqY+wnxr9EqTKTWXhoHZ6FnS
lohxbUUpv/xkLAQfXY/2bdiYNMBEGJ6exql479q4ZiBFz54UosQfPsPKVzx1
ePDjdsH54wz/lOc35BUu4ztA39+m67lsUsfLmV6kp49Wvw74vgF9MQdUXsDf
3wvE5sfl+0JwXCc+TqbWVGT+sUvkAFJS/co3MsXVai1PDldZ3QCzrLnpZ/Wx
uCrEfA/sv8MqOG3ml/PfNIBwg+i+NnD/JoSRX0jAZr9MSyMHIWnzHJXfFAxk
a5Lv2TlnCOAgemw9Cqq4PiwJO/VDtYXDGMPa7MECjRE52k1jqnBpTTkNYowH
dlMpNBlslxvsk5Z00WMq14Aov6aVCrbArlt1U5hP8qpAH5EMXjyrcpega9yV
tJzi3SNg16H3P3DMVq8nUXT8O3JGXxS2sVqeawieRlB52VJwYqnRuHA8JGX+
sGfwaHbBoknV1tgGEyfXy5RYmsWJFlu43E4NpEXbbErYoMCFUNXcsfQbq89X
arow/8J9ePFI2Dmomz093ZbtvgViTnkru3oi/+ZUJ2Lk+9hi+Enc78bWCl7B
wG3aYJmqfmc0vzlmkMM9i26NqSEWTUlyqsCAAF31H5ihE6g/GvVsVM4HhiVl
TuG5VzOTIayM/D2JqoTJGobrKen7bTU+qAte0jnzBEwnhEAr4HHhnwPpmnZv
9XDCqOWSbt7oXreexzdbqH5VBpUct1faX7DGxewP8YBHruAzPJBlFm8X7cGp
q8SDa64sVH5TW8FMlZRV0/joe3nF6HBLQfrbS1Ixw5djduMVRA0YPFKGhMSs
8Z2AHZ9WvZWuCqwGCLOWk1PfwHIMA2XzYfrIRG5h+6I+H5SruiWF8ZFWs3vC
FjE5tmhlOfLeiDmkbBLsAIVfPKvzxkxi8ABgU6oGvKN9PjQEdKghcaexEzOb
p/G6k/n2mwB8Dyc/oRu8SO5Q5wWQ9nu/sFtcfza+jEB9jDdWq8X96J0LPH30
xHBPZwAXLbCy5QUWhjStNmNLAqSXSfhmmsRJW2J9Aa8JO2DorwGisr5jcZme
je/GKNVhBGnUW/xQjcLKQpAcUbO49HCxKPMNWn0Mk7vY9/3oBvVcZgkPtYHx
UksAWAZcWby4sRBs95hGpebtzVLUze8i0EhMOUVS0oG2VTwSqDsO96951E73
rt7o1x5EEdikLeumyi+Lbp/A+xsSwuZ1tJQj1WgjkRmo0wNV5sWCGUmsFaFp
SpxEkuSrYXhVn9n+N34PHXn1mo3DEXr8kCtiLrwAxhkWtTGEDXeXKMkzj2WS
JYlFkIlBo1ElB8QTsUTtrpp94Ay0myPDI6L9SPydB31pQUgBumQdJ7kBlF7l
pZ0EM6mTvg10hl+R2Pk79zgg3wZ7HFToTX5yXjzwHQ9isPlFAlaOesKB6ZGM
wy465a78O1VqKoZBB7fzDU4cfDQMirfEBc6nckZp6k3dMiFaa97CaDdYe0eL
UxzN5wS3q21rSyTL5I28wpGQGGyiiHJCgDRmhUTixZZNAJAemc04XePRZJs0
0v5kE9zsMbYUoNo5L22rTHmHEkUXzpmA3Y130C4BkycNQTPzGhaNset3yC7c
qVQXY2MzhhuobKHWdPksIfrON4qRM6oWLKys3dICPQSEWMdzZozodvRdAxjC
ufh8uGwjHD7buHUIlBRoVSYQmBpjRxIvQYHRaM513hkgN4l5aRThVJx7gkkE
ZQhFWAp5xY32I+zdrCnzzrxwKTPcDHrYkjB7mqvVIRzCpprJSwoQOaw+lXvw
2JmgXigYZ/orn6NkQkTL4z+4rPbECiUK1q/XB9crHSoeVNr/10rsrS0zOrZn
2GD6nFTSoVlT+EoCK6UrIYPdLOqJzE7W5kItNd7VM92AtrWlHR6h0RV7eNRn
vDzq9gnyz2CATgKtv3JTxtHoQiyIY7bESSDwqG8RtIA6ROOqxJwkHIJDXeAD
pEjPIQEuekceue8boWGvBjMxyf+BEJZFqHveCNQKyPJzoSBk8Ud9T7dNhEfQ
D7E8Ud6MQox9ei/nXoEDd53aXAB5Vnquo7pjts8BA558oJ5peXeOC3t30TXB
+5bxYtrKIoRK76YXG20gsErX4mBve3e5ewbbqb4arlToNgTIO2Mw8CXbBxdd
8M4uuLc5TjloksHp6/dWetQZ/7x9BUaOw+AiFXf27+o9iYnMtaj3ahrAC/fO
XKn5Bd/usHOFSVhg6pQucB3LseThJCoHAT6hZO8Jon4WmWEAPnOmXyYGRgcJ
Yy37moa8NaRFOFNN1DpSHr230ywaqs1gLBjO5dK7+KwBnEeOjHEaRxAYtMwX
pNzl3rCKn56RTDvsqG4VUpCgGOZHu1Po55HJcCHkKeEpQJLxo3hBtFhgOoFC
caviUab82wkTq1qaS0mW9YpYbUzVxAaTs44vm8p9HTSR6ThQEzVMkcqbU17F
DYhJ8Vn5C59Wsg867GI2CHu44VKFPaC8ob6i6jSxCtJK7DwpNe8FzF4KIogZ
qDdib9Sp5cBlQ4kvcRmHpn64PHmPm5vD9GImcnGjL1nVbuAhxuQcLcJLA7ZJ
YKIS4EezYmRVvMmJa6pkeHnTatJ60nJO9IAX+zS4C/73tTBpI61TUZbhzNoE
l3lPYXxtBXozsk9KEZlFC7gdSd8SXJbJmmAR08DM2X+JnK9AF+syqbDDqho9
BViOewkLSuuATkwn215WqtQCvKSATCcjaQKHNjszuTp5cHtaonowqyBxhEbA
nabe2JqoSEPYZILI5t6Ur8e1rGjkcRligrin46dFzW+2FDcJN27+Zp7yEieo
eFdqNIuP4KWVhLqBYekt8GqsbjjXftOY4ppIxBIcYxXCfzs/kxVE1D2/Ydt+
qmtxbEHi5yiD353R6zn2NjbxTYRvkXGI9vGQia07RJHz4v/cvrVsw6VJ71tl
L7Bf4ivsgxezRL1kjPWztGhXGqKDbtla1XFyzuVovhg0CPgdAlaMApNoceHz
1qjInU9rBXSgqpRoxrz3EYZ09pnEtzZCpM6fxx/EooMbP58kDqev0QtiYiZ7
/KWLCJWcBcpf38mXZo+w7Oaoj1MJN7PzC6WhCfLf2UbOO2NPNQPm7CYKh8Gz
lppAJ6jO2V2tQBsvgfjlc44iKSIjIJ/GpBDrRkKHk1xGwPtmYV0X1EYEYw07
kEcXScb0SZW6RyULjz2s5pU/xjP22ZWgAmpOrX+wVHVf/4mS4Ps5Y+ptsWJ6
mPzvULofUWCA6CV1dsmozv+WH7XPtSgzqqhXlQY/pXD/GofUbc7iOnCC9PYe
la/b/Jj/6ACBJNtaoQ6NSXH5EEeVjMr2sfL0W2J+OUi6crCLxg+0/dLsWbt5
q2VPP2jGOoA3n79LIXVqD4sjErwVfR7EIIlbN22X3XgVQRBSJO7Dcf4qfKAU
PoZTCRpeGBE/KNit6GpNizjx43OMQzQQ14oVTcQEMY0KlRVPwreP9mwoOP1P
nFL1e+YoLeWS61e3OOM4Tn1PGscZcNABJPMbgs9hiBwvr7uJuyoU9oR6mb+N
+DwFaF+g0VLR3bTJW9znnLEd/i8YfMp1+RZrhlVXHWNls1WIEz7SIbnn8VjD
cisiIiY73D1BBua+j48Vr1Ku46cRKArjLwnXkLCt8XsJrZe7J8OfXaqcwo1s
k4mp3Sd1NUAoJPQtRtDicPDRQuoZeaFD0UR371jRU7VUOwpW9F+a6U9kMwvW
0o/90DK4zC8Us5sQtjU8xJEyAU2gIw3Qcl/Je3t9eHg/WrjV8lIKheLgJYzw
jKzHsnrVpKu4iTXdfVid8d7wiesBMEEdMGYiPWId/3umeVIz3Yg1KJ62DJII
8ruyHfr118eACM6GX2CTCEdaW+WYBprF8PRfooxUi+3PLRKI3R8GjW6PfeY5
b7pjOg7h+wOmKjXJkRGreCVT1LjN74+ghCIyTUS2flVZSYPVKZ1dXwet0JOJ
coxsOYUSOaA0C5gg8RyKpcaL0GnCQRwPYhUGbz/mNqLGpF3i9wvxn/LmB1xU
WS0rTbcq674W2Wp31ZPNmjRIpZvLfm08zkHxfMsN4/9lCfgeFVnVXY/hAAVm
kfYL8AFtRwbVFoV3GN7fkelSZt8VsqehHzuJWPQ5RgQmYgDZbbRfkBSUXCE4
Sh7UpYrwO0ZvwbM6wde6OdBMyI+vA1qgbG/TSxhFlKMsd6QfBwyOl+vWazIv
exl5I57+z2QYf6dip3rgCy/EQkPvS1pQLr6g12XrqR/4ZtwMfeqFUu7eYuRO
utm15wqo2PJkAuTMcjytBrqG1VlL4BjK4hoSt4cGiDGajmrCIFja3Lro0YC0
lAIG5ud9lM3SSkNnNVEfIR6DT31ISvfqWgLvw174NGVkdUs36nMQA8HXASFc
SE2NPp5Iei2hC9c4U0RZJhhlC/nw7mHBmJt9He4AYMLKpH0OfuwcbQ9oQiX3
dUy6z9vEiLddZOtisFGZV2KT40SbcVDLTHnxOE+DtvPAhftsUrcMzk6P1rIr
wVqOTHLvX3L4QYLySLKvvRvPEPW8UIytziaSo9Q/hv9HGGKy56/T9+SNc4o9
ZUGHlZz+5LMpFcJamsfYGRy/7QwqVRZes6wsGIjHlf0hbIwff+Yq21adv/dh
wLkQKfpDM74b33nBq3sRx78wVkHVlj5Nfenp14/dD62K8uYDAAQDv9ibBsrB
HT3uoHudFgzbpixFi1Ono05laGVOXWgBkaNdgVl292Ee0ojXjcLE4M8s7Xem
J+3UF7TBdu+8jMDTM7seYgCs5fvXakCKtWT3z7EUsKFb0Swy8zE4ubn0PYBX
K1RKnDgRzYgKLtGPhYtcKdLwSuDJlDJg8hQMTNLkFjmAaXstBbVDLwoims55
mfqNdO30uuPxVBGFCx8F1njd5sg7YOhL1x07poLlayfYnZ8ulv/mImaCafdI
Bxd69FmgjyYxcakNL9P+muVF6/5/HO3S7cMlbZHlSUN85ONbl7dLVzJdrWmo
3vxhp5sRj+Wy0ToekhFr6ugg6g/BLRWX6XBsfhjjisqdq53Jr61U/Mw8+LH7
Id/0HiOtKT58bZ2sGRMTRZ+ymdkYtQKYFzSfbKXlUwKjIXKzC1Do6VZx/YlG
tpaf0P4flrqL4jhrvRDHRRysUTcKMT9drNnbA6jNUzCzo4rRCkYAHpUtMtU1
Nx6lztuXFFa3PCj62TnxTUxdp2MeqpW27vDe5trG5Ot/+XVs0RGG7TFVaR/v
+QF70RS82gunOu5q+q7VEULI0bMNQ4vmNveVGWzeyYFLHYbtJ/tC144RV0TE
Q/kaQkkOL0gRoGeG981nqOv7c2ST10lLBpW/YL49hF5wjBpB7FxjVJ/wltEj
USDxf5ORcgZSYnfu2rY+bmGGz2iYxrpLidzVCAdkg7sWtmQbSbnKI4MsOVyg
MYbAyQx+RyYHS40BrslIs4S6pblJqYguJH7XiPhXkW/r/0naTjnZioObvD49
C7WJqCTFMnWVGcexhsbdGC/AGmi1LualCfT8UGaucWjhmwPglqelL62byhSZ
lals78jVxtQ/qF3iQEVIxLC2//yt0KBTAL8QPvBEK7C2mdSVN+U8IZmzHoow
ZGhE5tT0IA1CAJryCXUE3OZKk0tMxQqDyhShcDxdpRQ1YVxzvrrXfKjqzjzw
AfQlkX3feWmz+UB0dgJ3nV4dWGmXsgDq6yie661mT3RdKNrKYfk34+jaI0/r
YUB6BjO8Uj6d+8O3nHab/FXXL7DUMFB8OjEXASzQXhTYzpbaJmhWMU2jWWX6
qSW/hWYQeqET0xXVlTU3SR/kZJhxX4CGw4Dyi25LBANVxUttupsPIOnuIeSK
CgpT57rwMWF78xlDjtHk6QB/g2LDNaev2LETowW9FcnlbUUM1UzHAn/ZWCMM
qiWBmheVo2jyLrkaPbcDWLomDVvX6h8M7NlSOrMTdU7Zg3z3Wtm+smqx1Xuk
krnlRuEkTO8METGOwoRX4uuWhDIaL66MprSDDP/hbfvQU4+ig3BcGNP1KWpG
NxANtk8YBqu+5vUWyKHfLRtQzPfWmksw69TazXJskti/ASNXTuSsXWlC1N/G
fFcSyUkILcA0oP3QHO9RQZZeLe2DVGhcNFdecsSKk1RrVhgaj43SVyV2i0vs
CK+ZN6177hSqQZLruQKlXF82r0u7WMHkIOyUaNL8Ffna9ttVwepEpcRe3FgH
otZDn56V4AVRfOP2MQoyQ/axvHwJrftTEwFi5OPdM9TnouH+q/s+zD/e+d0j
WHumKzeeKNtVt7uaq3OsSBoJPj686msZnN54V34cLqdqUc8QGnKgXRJyu3Wf
E4bxASXQT4dzl6Wp6qzw/f0FyROZOlP/Y2/NGhkC001SwK3WpO+vRz0d9lD9
dBGjTm6kQB+eGW6thOZYC2gP96x+AT/A+Pnjs5uUm2ia8WU2QKNzEN3c2JNT
O4fsHv2heKyNynvjaW3d2zrkXNKhsBxZzIgPKzlPQoYQ5KcCfBUeT3DS8DHX
dSy8VSubCMEC+VSysM4VqS7CvhW+bDplPV1LOb6aEItbdfvbSDPRpKIURY1V
Ox+2X2451wvV9yOKdGcJQLaGrKEQcuoLmlE53Mj/goTmKbdX0EzAyzXsuw/k
uFe/JaHAalZQQP/r8gQ/e4rt9hgVzOKWXDzIEosmoNlGFtnNuTmzaBIVth4n
IYpPrpqSXPKM/KIbCy/Q0hx45Vw4Mlhg3ThQ867n+D/SHcGylcx7pES3nvJa
P7+qkgz1wkmdYtgvLueNp/Vke6SnpgKGn08ygY7sBQdu2NNPu1FSpH2RhTg4
zLOfU4O1fHfvdsB0vjax+VXIslMoBu7wo1HTHRZI0nZdLTwLGB83YbC4izpu
dOtlBObcnZBg7h3DfW6+wf1mKP/DgqltmTGX9fPULATu2CLZVl/3sCtZv/gM
hPbJCyTLR/HzdplRD8HB0djCeo1e3mFsam9pJgMhPrqrElWLziUTTOOwQ7Zx
qttqDzJJDZC95mN6jPflWX+rzLkSGYi+xhioVi3XFm/1m1t8A2BUv+o37r4Q
BgplWFHwqe0n4VKW9wOr2wzSvH98uItx0CxPotVIIAKNY0w5gtMJRd/A0mjS
CXjSpiiFJfrx0j2I/v/SYnStz9frhlQgPwcs3r70SB5/eYxrSLVh0ToKUHMB
3Gd7favbpEljr/7uSE/c5+2D4KUCKy1cPO9bDXCMGbYJvzLLscPjivBAUKJn
rnpoIQ4YHp86IpxMnY+1rDQCruwZjx+BhoLgjW+P9Cai/M3NFrjuuFAp7+wY
ZBBSVvfGbVPx7PxIGuVz4JJRrPK1pnzbOOIYCSQymXw55yHHpTx9A7o8HfFK
AQ88SskHFQ1byZGX3aVqikeLwmNfi+07Gut+rqZaiST8exYQBfayzNyYCm1Y
ARuLkH5RKuk0NWORhmm3XHtWTPAS0Slu7yv9Bjvyy7xmK4a6gdTO+E3+MV8K
wRO8VAIM89oxWPBCW0dXvV3w2U7aiNDcLb1SO6/UoJ+tCfgfeA27KEa3WldW
9cFkvha308xdICU1BaQv6STg3ASgjpTj4aPBmhq3ooK2XtVKFQlnOm00Ht2B
dvJhQpva9FX+kiEnD5Vnb4pZyRp0bQ2TjB8NeZyIfl7JtgDK9ZGOwuhua/Zr
2jRTQkAqXWBR/HrjIouWWnPZqY9E2v9Qe15RZLRakiIFBV20S/A0274RxtpH
5ztXEYUO3Y//f37xxdlAOzOe1CuwRiWPZD3x96v4iNQgl1h8kKKymNLrnSbl
EPzNpjhlssMq7cYoitnVgvq+W6BpLYNu5BFjWEKjSkLaDVSxQfIb+FjvKNoq
+d/pCl7RvBQLCk1atdAmbstksy+mZbqO9a7IQIyqHUQD/JWKK4J9yYjhdvBV
b00iOefGRyVurc5OPmcVXUXsYdCcIuSYJQI+/s/HoEgeLpCBdFXejFnNCtU0
pe/QluCai5ZMFYUvmBBZMgDCisiE8lmQzPUaE3hV6T5UqyYgpsS5xbY/Z/Mv
2zgIu4mJ71to1KJX6C4rpQ6p9SE9NjVaZFYi8HVb16f6GKwVpOa/aknty3iR
BPrF6t+bDzt1f0L3tuwNLA174zuT6+5x59hLTY8Sk/S7z3tiBhd9Zl07Wk96
2l7SECcZ3YoyAVU2YpPfHgWoYBV0hkSwVzYPJatCE/RHTI54WuMVN0nRIuWD
Os6dZVPuJ90rKKK4t5WWh/yYAsqDl7Jq7bDzQX1FzmZ4j199+SxOSppKVmcW
Xvi86IleHbOreU53Roaa76ntEFuZfBAsWuv3yHo3lRJaGNppIi+SsV9umtld
PYxe2IyPnOG6yFXWROar/WqDljVzXkzu57V02FsnvCUeCasbOjlG8eiG5cYb
JD3vlaPyYM8sXOzrazfd3ei1zzqOETCMd+RGubuDx51qoysYnu0MhH2sm/r7
QmnawF0/IjX4KCVuIYkVqDzWKNz8FqaSD1KxCIz76WTw8DV4vHhIEWw6Rt7O
swuYKvkqtIc24asaZ/R0kPJLePijfDEFmEmfkbEfLDZLS6IbtKFhsYl7Kd11
Uc4El8W5Ydji/41ub9dSXV9659Lyam0fCL3KSxmGLaiR90+KHr3q++z2shPO
3zyCONHuLc1cVKngd0r5EnRNZ8S+sl+YXWc3mOOHHhgNRXpL/PbNxej4SxOW
L4s+yDHuqrIv+4h5Ti8u2EvPOfjJyRJql7IqaR1hGko6SFGp+YZXb23qzpIC
6o8bGFJUyEVAz7szpKzBHDqWm3AqDLA65VYtUppgN3Jx4dkhZRwO3qG1/Ovr
C5epooKJ1S5kDZcOIGTIvHafzsXqS+Ao+aW6fdRJ81TvDaatQ+rtmOg2dGwo
ji5CHq+lZ+qoDwOQ4FFkNug7dVJ75JueiyJypP1TCpH8FmOL+TEoipR+VCnz
2LQb95c9b0E96CJ5lTUn5EBhh35ASpLTPFJm5ITMrWnNttQ4gUceCorDDJMC
89VkLCRkU1Z20aThlqaOjDqZFuSpth8pXXiZvb3BiHXxEmsGjO59ZIMl/RbE
zK1H3HOBsbs+Ng63hrC50cB1ex8qvk2uQ3IN0e9yCeD5dOUhhCyfixDsfITS
tXvDTkqFGiYcMcb4yIrBia6UDONM9hb2EoJUQhpb2FrV03/J6SmxS5cywxHx
n6BAP0wJ90YyqX19Bj+hPXKmKozR98nXoQshzkZjVtqedsm5eIyTDiVu0wmZ
7apbBaHQVdFbpJPv6E5lFocX4enqnCCYCwX8r8idbzXXBEf1ijOTEDKU2+s4
VrwWLpt+WGEyYHj81H0fRhe9fcvTH4lpcnrZf4zeb/0OiS/lBnsjkwvLicyO
luV3J98jdVUC8JFzBU3FCVPJXTr0GBIOLcw0u7lW4LPMNivYOE1DREG76kUY
VumkOoDs1Xcystt8wrgnpWZD07dxXtJIbbHwCCpaOy8cRY6c5ceAcYY43WCG
lKEt3jqo9FJcUF0ZGXgIlt431AhCqa4+AJz3GcSzSZ0p+rDXnm3zJ0HrtWrR
3AJPXKL9ig7iGMmzhTJb/Ql8OQ2oWkPt2wLeiObVqFwSDCsjJwGqTIixdVmc
B2Q67GJC+OAcH9GiYjmeiP0=

`pragma protect end_protected
