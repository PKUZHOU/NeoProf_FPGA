`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
b1GzzIEQy4/vhv17AvuhP3OYTgmMz+GS8hvcpFqi37YytT3h6Cb/skDOwK2xsyKH
+rU8gtiZL4GFoOngjEeYLxTebzOZWuTb/7ghXJuDplRAhdQaF+DgaxLub88YZA3+
GL0DQrs0vKCQiReeE73V69ZHjJgQTc8E30iGeU+1zoA=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 57744), data_block
9BGx78uBd2d/umx5Pt/rpyXTF/mZrpsP/LbB9lOJqeCmpb/OIUGcgB1QQoOo/0t5
6iCvOb6kKuRgBwnhBEWOjNiq1XTqQP/7OC4mI/J4DPWKLOdxZ3MLH38caGpdGSmV
H7zJovH1Pyxm0/WlwgOiWwXt3GS64qgXb8GFyuXiTVUl+Ydm918QsFjL8m2DnQvD
spyHWpmJCu/YZwgdEjda0RdWFwjb6FDmlC5Fgl6kY8o+Fb0mdMH/3msgocds5cj6
6n1wgrj2YIMbbtJIQY5F/xAxEWb9xTubgPh/gjBiKdwLeBzsa/2faU8skWMxWv2s
i69SspNPdJmdHWFnNSIstpNxbns9+pTh8b7Deu4XWVQivwoEdAA893pAoXQHOWZu
ltONuZeeoM5OQgx9lgu3DZKdhOq5pUj6d3R6mBM9Jes9RwtDZwJLVpsb/rAMQkL5
X77whL9SnTf2pNA8TGxs9Ac2JLxzSQ/ylO32xpCCawaUyGZt8NIDQymyXcwVdlCL
x0zIIHSn0QrJYerSZSkfUiPiiw+DMsyGYdn4hWtzB4ahNa9U84lAaT9KNRAFE37B
/Y3CTzvJINdC+P/cjKF2LwyfBQUYPjCjHxPM66ZpZEwB/JMbnwIpxfGGRhNFdTDj
IenU6k1DvA6TmCTRYnb8XjdT87/LKbV5Koy5JlNpx6rKEVwu2zdlNxzPNvyZ1KRr
SlIN2XbRLiYt8fDvm7JeAVFxjSydju6NNvcrXR78R0KMKVMF1vlYiSUMnjykjz2+
V23in/xq2gwVcwHHmlCOj72Lln9OSbXVw7bGHwoYhHLRCziEOqx20R+OLzxbJm2d
QBlEl6hUW8WpzghqFe0yEtT7nKctsm28+ra28csKLRnZTKfV24tnGzgR9GJjYffr
/AxHNwRPYhc1SBKra1rH3uE7ziYOvsZc/PtHxDt4dImU6I/IYHHe0kXntjpLHdB4
Bz2Dso7NGbpql72P0DkBOL4hHnFWrz607qKHUCNDwr6PveDQ54iLn6RWMGdX9C/z
29W7Xh5TfT00vd2IigIKhmp9KyTjNJLTuPEafS2KCrUIF4fgvwT89fNgJtCOZSh3
LrkYAE3eUzVkB7qrGxBlxbuMyEuIj/PtUkq1lkXUjjCHWHIi1Q52HScY0K5OMEOY
OZooPP7fsBPfjKsg2PXfICQEYh1ov0Cd9U347Aeg42cZ0KWV3X6kvtE6Q27At00m
75GToUE4k3w4ncgUUf5E7+nNXdDbAf5cHFP63TiLgQ6cFGGX2jtZ0hxQpfVKrNtp
aI6QiAujTcbrOunOG1wk6h3PVAamb1sI3m1Op54zpIK5qpmb9c9quW94UKrw4BqF
H7+pI8aChKH9qF4YHstRvqQB30kY+atDtpZmVMfSyjgkzKXlH2EPI6bibLbAUkhl
OVN3HHKjPraqSJwriyYRoZL92FUX0gTmySPsyLZVWxfsQyK9cq4lSwx785hXMJwS
RYhBswr2SQYZfjOmTDh3zuvTT7wQ33znufKh5n82ckCS/ji+WR/4Ad3Up6agRKaG
2v8BjNvXMkIlDd/GW9x1vOEZAT1IE/PjnsuuKDuvToPck7Ywbf1JbUYbvLZ6xtwT
Tf9AC1TT789K7iGpxkdsw4cWIekv4f2ZsZXIQgHaevfi70itA2UZoNKLo7Q6fKaH
NlDyHCR6Sv73yTypXMNPrwSf3PGXFRTqPMEcBThpMoxrhOUzuznFxftEZD5b4XTe
fiw8/zqhiSgy/SyK/YtYIga4JcOjo66PuxjMpce4VvHUoUcGkhiD8H8kXX3o+CHp
7Qyfmsxc/Dh/TyQfKMklL+E6d1M1cKb1n2oAT+73Uy/EIX8y35ZJrkpHqDPeD2h2
P5Qoy35910f5QDilWXpDxslRpkgcOTHs50pg4RodE93iTRaFMb/u6+K2Z6RwjfSj
lTd2Lv7511ax2YmvAJhItHxknL1n7ZBIH5btTk/jelLSCpJj5Og3rVYHxTevReaP
CnCT4u6DiiBnYvfbdEPv2NHNVUAtdxFMKkCI9focDo7bj8w/OzIhdSKEhGdj7FCS
Gwp2uMe8mOe/saK7oKE2h7wxFdoK6DXx7R0mBrhu3e2mfxk81WB9yV8PSUkpaAeQ
+5xf+I9OXqyWtdFMB5K9Miny+pSQlHOqr7uEs9MoJ4zoXe/eud3kXY7SKJm4w4wF
qCUGqPTzlx3/wmfKCsFMxYmmLNvbfGQiXz6x9ikY0mLJ0RPhJIRJn/G5/4lvoC6h
2vmZwG/3fI1Cyk4sYOIMdi473CV8FzV6HPJuatiI9Ao6jCtNxDg9ZCCoEVAvzaYj
bE7xKh7aa8f0135IR5mY4mpeN5X+H9jwSOihxUuNJjOzx3ZZQj0+kBt+4iXWcG/x
YaxoTzRm5ywRlldiGkcEHttv0sxUcjY7eCul3gjHP5zhrwCWVE3zHhqeI5HL4P/L
oSJDWezti8XjbBUfd9+O5sxExn2+yplu4xruqdC6I0NlPErtopZ78H6DcEUhAO5/
94rBM++c5/1FiHPUDxOckKlKuzyKKEU/BT+3URu3tW1UZ6wwhncgcNXoDDQHY26Y
1nY53hgB7e7PgfKO5HAHFdqTqfZsgJtph9GYxVdhBsuhYrMVFyAsEP+nMmP+FPTW
07iXgGekDT5Cc3IuFGXq2dXsT6ZbiTX3flWsi5U0Qeocf+z9QV0M8gX7x+rh/Xhb
POG8k8LNiLojrr5OYC1U8ls1Ujx4k89MwthOi64eURQwUmvWA9Z1aC8P8yRnPB/k
zZ15hbjxgOQTDLuuMjpBnuSqCIao7OwDD+FK23yd8yd2FwF6vT0m5iEeWEsvEAiz
rfTlp7KtFsDakrhO2VIDUt4BACspu9hFcJE1FysRlrWaqDXmdPfDrky47KfMLLsN
cZcANoLedSY/tP07FfFpOktM0RwGHts2IrxY1EpyyK4uBenqW1kqIxCYBymYFwBz
pmLkCn+grdqJrqhctFnc2iugzQgvaEbhIcoD31tcYdxyXuZlGLAgNz/kmL6Ne1Ov
nev9sA2EwNFk0QzyosSuqykxp5ZB2c2kl1VWSfQ9qygCscCoRxtln2++YwBIg03H
zzT3Uuo1on67KbMjKlh6AHN5Wte3Z77vx5QgVclsLIw6V+BTTrNdQO2g74KbJTkE
H02F+quZ4LWAjI9DvyoAo9OQ+6nyk6vfNPo/I+C9XQ8M8e/SmzQ4aiBWOMiVKP9d
9iUNFAgVFpWvwJToRNYZFDvojmSo0Z73xOuipGtAjw/vvwh9pmGxhAWsj0sjHQOO
GLxxSsKfoDGoQI0Nom+zX9zD5vhq5RkxVkj5QHp6y2ymbTlQHkfUpkZk0+o4UnCI
LOFsl2aEOV9p526iMNX8hH1UgorNm78kP5MCs5fuYenUdjCUQACGe05Fs9DnR+Bx
cpMEIYZ92i5WYtuQzQS9aRUW/sy4nGBJ+pEyiOUT9Yn764ul2YvzP9YBVjyJ+tB6
v3f5UIzSFzztL1iKyk2QSu4a96tZcIcBLjn+B7A+S8PgPG0pZtBNW/v7rjR36vbJ
2HTNtgO4EgU7Xu/Ey/ZCy6ErjBeB+TJzWGLk37nYR/a9iYoTreBDr44tLYmyzGX8
vc1vhfecmtDwOWF7Q83c3QbRdyBgvfzu4rOEbTViU4LMIb1h7kXmUSQzRuLv7qvL
DqN7eifF3CepjUcnLt7YXLDkT/hin3zyDSV5kdn3p5j7TORRH+soY0w43PsK7gyZ
s6jCqgoXfZ46ohIhnA3P5qdBfkdeII2zve2AM1Cyacv6BnivDHd4rs10qUelp8nQ
f+K9dP7R/MZprZJiVnDg/UfdIM+PZ1M6CDq9A5LITE9ns6F4yRRTD2RcqZaSHRvU
XcnemOlqfdMsR3LtxnzQ5iQ6ghs8BO0dkNN4lEnop5QIFWzgcBFTLc6UdvLx9yQw
IbPKUGgU6VfggkoCr9tbKF6zQEpbyrKC8YMlMmL3G1jnFHeRKiq3cC+SrEMKp1Nu
g/O9Mnevenn4dm2JW36LyV+dmM5Kw41791a4GF34iY83Hxu0KK0p9ncyQ80/9HbH
ap4MV14YscBPmN72Oi5GzRMUrWQktsSg5ld141k0IuADdhmk+g8j40I+oETtF75d
ltEYtuOFTtGd2uUCELFhMmKGMsPmsxO49KAvPKyEy6JazHMBQPCyS+OjHW7tMoqX
RGq6yB2yQ0sUG2pdyv9AjBhu37tho7Kigz2PHVimBWR/oLvGw+k3weZtYUEBoI+C
Jdflcxj/ZJBoREPY+dy9bhYPtfkHzXqsyDVSoq4KLoZmSywQLtOTYCNabCj6DlTC
dPw1yAuhvd/q5hELIxcfCOcq8JWazEF2Q2DV7E2fDVBGxHTSuxtgXBGWpCnUy5AD
3kWi13jRUVLkB4jJ+sCYk8taXQmtLPDK0tkK6KknljON4QcRPs88smo9VBfIuojG
OhbrCou+RK7BrTib5pZa5xx/CXMN/69DSHO8W1MOJCeloXi/Kfwq3RIvsir2z1vR
jbvjeFhbfQ/R/TUfjAxWopY7F3aaoQhnyGLACpBNkTpBjvSZsnhKWMWStn+RsT0Y
vFN+6M9tkJtPxRKYFXoHV++gdtlXMIKOlUv7DeH8Hq3NIZPxHhBbG06srFeLpJ3w
LN3wgFue6lVLVuROIrb/Rfy0gJNAcJ4AlBkmDvduI/rwYilUVdGi9kcjx6x4UhKK
DsieKMKGy60DXMafJZbAIP9gOq0FpxJnCwc8GtkwWkVVWsai4kjKDwRrwXr0iqXR
HQJnFJsm2euzbVS1ln212rB9IB/XjYNSjpqK0QImeY6qAFwyNRCNB12UqyXLNUFd
wgm0WH5kzn63u6aJECDTPYpkzxlJzDjeMPEWOigp6Oy42Ls+JCKEqbSk8Vcc90To
lvZgshFySTBZrQ6q8UrAGJ8bvC3XnK8q+iBhb2ZwZ+a51VcOkO2Kw8KQYRmbPkSD
ge9XVIte8Ytb57+yjyjIMICkCpUEEja1TjOhvtInczM/UViCDS5qTWp8OyHij1Nk
qEGHnwKiZwvJU3XDqfNu5RPs/E518adr4UBmDxQGla49yLT0sQFJcbq9WrAB4EWI
L7rFD6T7cZBDprIhv0fSeb02xGYCvftGWv+DjUKtMtVovPUWudY+m3NgdAyWS7/E
i1C08QXvrDV5SqA2IH4+M0by0rAlCTaLjn5+r6MOrefYuHJDN1NjvD+KWjnGUyeG
YC2DIO5UfgcvLc/JgNPY8zl7ESoZIb2KkfD806prtsAcuTQksd6srvgwNGCe6r2h
GumBAJdFcpkJCG4Whq/FkwchOxbQhHpL6BUyVMdiM71OazcQv8hfgAL2ZiSMVwcx
rOcSAdyBayQBvgSOSJCOq+EKzw1xVRbeDfMk//aEhCLEO2+TjSAPqihJdlBkgvvL
Pe7xlHUcII9pjrOu51+qM9K+OaaM8ZXH7itK4KAV6XWw0O1Al5RlsObWBOdVxl81
5/ljb9Q7WVLIFpBKKSRbOcBT4ucqivNKOqnH1xnfMlbC+hENBGZ6fUcdZMGMPH7l
YtP1c4DH1nxqDmzEZsJ/z4NM/A2OqFMdd5Q2LaBCWzrUL7637Qx1RCbNCPZq59G3
VEfGVvfcxLbpkgznCuqRSBVzrlZC8g1u6yQ/FMaWDq8J70reKEb9OH7j6SfphAtL
XBlxwUMXg918w40saSixpSKrl0o7b2pHb5uj4gfAjNE23l9GN40cDIgRFgw4uyN6
SK5EtvupJv2oBxQx3tuwo8enrt8BGZHykuBiHY7nBVYrmXeYtibQLNHem7G6Ek8s
OuR3M69Gx4DBU957vw7KqQj3nt7hsrDybgx93jgoD7bKRcKi0MvfpDbrS+yyIJAx
SXE9fAenexK5YUUzzrkLhI8TuuscMTbzajY2ET8X8sUT49nlROA9A2zlT25rqYQk
nmQeqIgB0VmaCzNlWCNH2KWVsXtdjCiTZjaAOejvtQ42eqqFUfG5yaN+fYMINx8Y
nwV7oF1f6+uBh0+2HpeC/ZW61rsKUeAv46SJI37+b3FS5zGcwAWbfcDjTYTBw3Rz
RFPGspT3dwKzZZnESNarTiaeFlYJhDwM/Mio6fijzSnHJd/ALinO0/1TGMk9gXsK
j5PHul8az9aomcHgI7AXZrSlfsUNkrror7JDLtQsTNQwjGT1ziH2IjPGVhdU6eY/
oU0xftth2diFDyLQeBLqZnZcuTUNtoEGYl/3tQEolDLB2Zg1rTVdLNHqClCt35df
66at7j1zPy3wM7n8Bb3o+yDT25JIIgFsRYuf6En1JEqDW5BStQYnXVu6THkfHxcC
MznZYN2uwwHX4veczK3obvfKkgcks7id0jquV9pGN2b82YNRL7EiRP0vDodeqyNF
AnVrTC0GRKNXjQ+ufV7atHRRQVrOrsN4d3gYd7rOtG0yEvQCRwWnilDxPxpVG1oW
c9QuRGInTTJDjKjJWW8xtOoTsvCMLxyZ4+9WL5uAlSfXm4VBsRHdawx7eqZ5IQSM
3Fc3oxHZi5hW4bod7xuG+TkNf3tCU46Nau14hm+URNNOHSFg7yCqT5D+w2gKVgdQ
AhRdKVXgQH9R+6YXn++CSznhiHCbQXf4oSujt2gVh5crNgM7au79F5aXj3ScvK9E
gj/it80qV1w5zy7wJ8RGYr1eA7cPQG/J2B3gyRIBpm96LtdKTvmst469XEf+ozJi
ZtO72wJQYkrALUzA7AdBlUVQO/DNrmQsU7vnfFOTH2YGwXA+8oehCNfjrNFrAlEZ
9mnG1tE0WyWM1gBDv0tjfduxr90zgQQxZRvtyOwdWcGMekC0pyIoaaQkIibKaEcn
umRi7TMrMRZztSom6lWHnGTsu8dZQegON5eNqrTOUbdbDD8uYk+7kx7KXxpvxjAB
l2TSeojQk3zgPJeczvokUChv2R6Y4qYBsfcc0bEyO/Al6WFOakg2kG8nTbFiYsDv
dUUAld5Lz7nfW+NFrEKVexwJ9pcqKLup1hK3e3eYOKusPZlrCssIk0BEVLQT8U8W
Hj4xRXpATuXZTIK9TtFgwKaejgfbMOlyjlJJesQCvoaQKf26xw5y0GdKgvtaWuYG
/TJrQDF+T/QahOoSmndZN2ZwtF3qEonXBKc+U/asBIsRXnXhVo0EhsHjQXA8swaG
LwkSs7ad26qRmBMxSJXYgjyT9Z4cMgcTXr//zK0NCatur0VCu9B70Yk1d1NNwUYK
4T26vV7/gRv4XrgiAf5zthfAJ2DqRaE8nlmb4qkjTrNliUCPBkt5mzZ1ycogb7xh
xd97pQArFifAz9MP+P+kyq+hsk2NoTe1GURohlgxMIKiJlf0+hJrZ5kHH526W5ys
6UMvS5XDlnFuTryAvFOFnKyU26t8/MYlhBKrDQ0W1f+YQnJ3uI19t+wLxGYT8JAt
AgydZeSMAJNaGfQeE5YUXZGsMsiBpafifmnfNbX8kQR7DGxhD9vyh4o8qNZf+Rli
RdnuirRcDKM6PTYzFyz1dqsLSJPWJZHK3xHhDvMIuDDWEXHt2IssElDNfTkkt300
3/7O44EziwjyvRq2Xf+zCUBSeUptGZG83wPeZK5fhOBTyiG/bN44yzGCYYht6Qqw
+nARepIpewodqOT1CWtnkBAwWqig3DThuqUULS3sqbglfBLjVUENUFVBKygThVod
nFXaL5vU68PSIanOi8lPsQO7BneSMV7NMvUVELpaIDi1aCTBuk0HyBAWNxwvtHvV
iH4+1ckcuu3S6qzQx/kFhjKgSmr+TDav6aIuDMKzgZUtSyL0nxs1JVpowYqJw+OD
QoR5RF9e7M7sVBlX3OZWPtc14riKbRcmVmucc4OLelSBbEhEVVePmne8qeu83dec
Afq3USWG2yK9/dhX01wO1K16yOO9e+hE8/n0RKhgHn6wRjx2PLOZyDpaH/IvPaog
it/rkyalHr7T5TDTMdj4yfYYgyOgFYoGb3B2xIDfUV92J50i4e5KzSEAMv1TufMh
q8/CCK1YZI+yNhhyZmaejux2y/hpvBpS5sh6rrngoe/ZnbpkcUgjKlzx2Bxj9EDV
z1/VwSL6dNCCj4DISDyrUrDBfLW1Xpd4SGLUYqal0dglIV0AM4RBebO8RcwDPd9d
U55OBFVT7V5oN5pZpKU8+m9P5w3tD0RImjpq4MRnKSl2QCzjL8q+pXD2Cq4n+K63
EkR6LrRed6W2BV1KJ5iXFNNnD4B0ahpjlvMFrbgJnHOjrlx20jpX7imwImOq4VEc
9zvaEeyJsbogVfIi4PlactsIh/wYqJhw8Qaslm25YD4aqIo1+dusUnJ7D7XzsW25
bMT2KktFYkC/G/QpaoQr7FQJYw7dm+cG31aLe9t+WBD7u83gmsiH6TKcV5lu/wcm
/wXEXYLPMmuDo2qysZvTPujzMiILN/xB0tpXHumrxrUgJ8hVe7G4grtkoGDgVtuL
YRyPeJYjHhti2hKx5A03gPCddWMRCQ61cY8NldJTme9TxK81bIOpZbL1vhcfQCyJ
HJcn+CM4ywWwF9ekbm791K32n5z1VKxbBkN1SRznVRgoYZ7C8Yw6RVI+uByYv/OO
JOhh7hiG/Wj+ZOh6X9XZ/GoT3X4WcPmv4qvgfePlkuIDyCCk8Ax6l6yjw6Y+E99T
vkeohBEPpGXLxgu4rlY4h+252iiUz2L6cyCnaApodY5j2g2R9xPQI58A7skiySDV
v5qgqb3eK0GOihVeoTU5+l3+UOqWQctd8GGl6RiVZLXtf+SYgZR6w3UtMlKSe+7k
Hazhqj/ToYmEYZ8G8IWzHuKSXkyDNDmLzrEyWUSe7KGi2DzEFvxUM8R0tUx0OIuu
ZH+MyOA1cg3+R+hdWl1mE5XQuoAUx5cS9N6vpkhwmr1NqjhMRIgU9maMnMn32SAh
YIaI8dIe/vPL9HYSHvA/F6m0xWXMnfuiX1ePhVvkiGul+JPe7a0cbVhNXWIzb0si
rGT1oz/yGDqztquUsRD4BDNjxDccJ8JLAaMqKWGTIPf+cP2lgPZKUDiWN2xfmJXr
R8CgqAjsSLSElg9R5NR47QLsfJI3IJ0OAGREtW5+yCZFVYEWrNw35wJ5fd4l088B
u26mRUha49kXpMQq3XI7v8PWR6P3tAcGW3PieZYbz+JEmg4fuiJ7do9oPc2gkv3i
8bOmZyQ/XyRaKEQWcQVy2SD8HN9OEMqo+Px02TACtf4xdJytEbvH6JBzkaRkAVXM
eZLGVoiLIwD20em38RwXheTRxseHCrgxXKgqOpwY0s4fo6fMgSvqTo5Fnf34RX0Y
TeIdypUOuPhvp6+gLcsGFv19CPPipBTpcJczmtHa/vJIYzUvCFturG2bBipZgu3n
DCA1LieD4r894Bgbli6uliRmeyEuu5itentZv1h+IYVeyltCuLMNrYsty5HwsToz
uxcsXBdWTvRno1cmY5t71KkMNChQulFdTbXYrsduo0wVr+y7g9uBl3vcLOyYRgDl
4LD3cti+UZPn9JG/1ui5WXDcAjZoSh6fgDeYhN28zKGs++uylOoZke1cc4h6hvLn
9vQ8//phy+yXUAW0/xxBlA8gphmpsN7UDmUzyIH3h3POzTbGXjiOM2I+nDAL96Y/
CkBvrYveofdxQEwwtEqWUt2Ddtb3/U/B92hlECuALerzavAEBPv9NXOdQ08TqKga
tmye1Y0DrcJY6hthDZ8CZBdb86mhvRKjeqhoEHRafIwZln4pGaS0T8STOP9y1voT
nM5XeAXZzJaNE4IpMlVFRH+/nNueMgVVqV0hmMOwm0y6ErQEhbf1ckk37PSsee2E
sa28X4/IVZ/LPZQ5Mrw1KvGZIHHdrkkHvazzcgQLgd7C02T+/kq/2g+AbOs9ITKc
mJ1A/U4NT+01Jj6TqmGSXNdqXMqz9CUt8PuyTOk1wNexXm27sIkDe6mg+OCcIFMk
9azfb8drHr4apoQJUJ9ZWyynvvKNIy/DMBequ0zTT89Yjyp0T+LnHwlJIDd8vaGX
oiHY6LnkFoaTfqC4v1dn3ZPwTfsN83q07iR0NHiuJNJCByJ/FiKQLOTi0cfv7WlH
Z4hm2TGd7Rb+NOir5XUjfASlJ2FX51YVBCI6VL3LBn4pAo38fsxsYKCwv4PO2AnD
zICGIyzSoPa+c20Hzu1otjuW2RifH5tE6vxkLMt6ONZen+mX22aiqeY0fS3rjIyK
wNoVQkie6cn/0hLJi7LTsdVQU9ozx2+IbbOVSL3eYC0EmwHAZT+TUx2Mf25Nicia
wmcO8GR/XAtCalj0HVqsDihIH7wQDdY3nYJkL6RaISf0WTZP4dsVGiaQH9Aie3aK
16DV0TKXt5i+DxPgXQFbRVdb2dJoyTnP/G8yZ5gjmFGbknZxyufLjp9tV0lhCcyt
Phd/rOQk6VIL1U8UP4a8TXCjGrJ4zLprEqQM/jwmeusgYZxfM7khHDLt2IIstGX/
fDCbW0G20FUcGw1puJTIrIh0fn6mNzoc/8CoZUtUml7G+ibfrJgHEPlUJWf72b4X
lMfZK57AYeRgT8J3FQ5zlMN4hr5WmH68zQBreH5B4Lxb1riOsOSH6wbfmooAGlDF
aFxM5TpSP3zqtQ7PM3xh3KfjatGfWDCJUOVbjE57+7hM0RjWH3sxBS9IZPGlGGFx
odFTSNb9Lp4UShra4/AEs07i/V/p734XP1lh9FIOTeY0lD0nzyaq5QlredN2zneQ
cf4lVUEewIbwHp3HTxRYKFum+WJ0Ax6reSs5dGbqRoM+gjip2aA9IuTHk0uWskew
7uJ6ijuB/dFI5CeHr4Z/TqMRkhq+cSXgCaFSEvFGUmIB4L2VpNcbcg0DOxN7PDvp
YwtWxSakTv81oGuVL8Ai2H0nh40eUPKLJnSPEG3vXJ9FgquOKMiF1Cfd0vDGsdBW
ke6xoTFCGBArwsrADbAERHqdrsN99HxtjloY6gS7e+ZCnKxahHCBqUsBahwq/4MN
JT4OadpWF6n2u1Iz9LvyAJIvd/RKREXMNbNcQrOMF4wr0loPF5pvCsP5GHKg2wzK
11PwE5hkVjcQ49QWFUP7xAeTOnhf9jJUpVJ96iw5iC4y1IfgxZvpk9HIkH5wiNKj
456FBK8prAgv895xs3w3MpqUC1DcI23V/X3dPEq7OcQ5u970JJUDo1n2C0fILbPA
DgNpqS3CJWakkbEnX5hfHI0IAEsPpd/2gFoauh/jQslU7WIFRdpIvm8yaDkDCoW9
KqOVfUtCE89lCiIT3+SdL2QZjGCuBFqoEB3CQAOZFwxV13kKxdc6vx7pMb87liyS
hL288bUYtKRp5+2WOCfEsvxPHlIBHM8cCh+GWtFHU5LF6VAuYhwDLtte7U+zBg2S
U/uw5pL3JkEFTJQUItsdmkeo+5R/MTithZRMtcapKgxWKeGDsQaBtE5CRE/QZuwE
fyU9DLgZakFf8b0xN0oYt3RbxHiC52MClEPYGBYNN/53dtJg7E/VI/tfiZZUXw1G
WC3J/ynq0Am7Rl4o3jacaaOOdEGG0hZpEvNDzQF4CgJg++JY0f56gWkcLH/eThMV
Vgce4680Xf4yQuEPR4gv5PG7p/CbBgml4vdyRa4AVMxIxi7SUZDpEuW6E+lSsYcE
iG+rIYW4qnyY60Xs94AQhjqJI7WF7znLyRmf4HMiwVe07Z8aXYGnbEbEUrYwcUuE
JjcA4xkMIpUjwMbNHApcZ4UG9pHH6dlpqKUSD6yvBTbYKz3rPrhnvFrxTbIJt+Wn
q77dCANFbtLqf+y5mIoGqpkhmorGKH73eFRaZqeS/2KlmOIvLgMBvpVrEarTvK64
++ZCCDJCou6aqr3O4bgXJKPsESR6R0mMkftzwhlPzAdjIRdWMySDE0wSYUQMzZdF
UeNN7yiXr/lf139QDPCBWiNL40/vxKuj7lcZ7bXlta5WHuu3OF1JQ7ytYpPikLXV
LZX7x4Hr02mOaXdyDCEOk6TrvIe8/BaZi0xXY96uaEDp9R84HGw4iiOJxVVOkTNG
9/GozBrsewt0uqpco3qEnhfpHV8EoDkPrGFXVar0JIQNylg6D13X15IBW/wP7URb
iUqp7R4CgKMV1rDKYG0mhkNNtkETEvQiOcP0Y9U8tho20kzNM7j27Lo1HRtCx8zr
28aQ9wUp6Sza8miagwN1AYWmCl6TluUDq5XAyvrBZVyhQd9Uc89MNHXk9xI7CnJK
QYT1iM4YK1P/0oH2PR1MXCHGEUwQ/O4Hqz4DxQ+IIe9Ps4MY9isTT+Y2+HcNZRQ9
ZxvBp8FJzlCbFxWGtE4iEuXKercQqa6npySEa0BkHtoR0+5v0BztyeFQV3b++2j+
ZJEj1tBW28bWZA9Y+4gDbCXd5Zuev4h9kZ3S404+r6o7m/yQcVe6tD2joCfNyLqN
sQ+cQhVD8XWLCAuwF5Du2hqoYaxpL+NaTOZetDK/8HkRIHhiT+wYSDZPhDslT2AJ
RVh2V/UvkyXC0WSE/IadypJljBl/125qElTevZHz/K8y8ZR8QhlId+eYTbhLShHw
JoEmhu3F4IyEQbrlrvyy3HHES5pe/dz8JcOaYZ+3Vo05DOVmPBsRbnpO6pAwLWU9
IyGwnzDqqXEqXPVJVc8j2l202irNwpILKOSYJM08EMHQqa3tJtwbD1QHhAn19Upo
Y+mm3YMYniQuC2BY93YcfKqKrUXXrkn6zev/xUGRADNcyZh/29hzXQrg7UK0KPsS
OdGJWCizKE+DdCsDH0Zh7mbW/8GsMEOku10b7ldqaB/GQZD48OrLyyPum2DNndhL
YyLznAIZRKXw7g+6q7ZQ86PqnAuE9euZ9+0OjLpUaMzfJqyo0tfEhnAnsHZE7tog
kDokHtikr1x00He0r0l0iNbn8hw6mh6/3rKVhpFdMIvqTsoRr+l5HwMeqtZIA5cw
Kvn6bJVk7mnkQVqKaZ/4/qjtYGipjCkmB/0AU0VeXWnvuJgEz0vUK3hop5UrGHF7
s/VtiGvlRS41Pb+/Z1u6dCmi6w9kPs74pI5ZFlpdsuYKVb8/T6J6qMSpiMyNtcXS
aFM5dTZWGOlvi0BetCHUjZK0Nwwpy7k3W53jJan3/vceqAzaUVph4/upAYohdm+s
s7j6fmix0SGdNsClfYsvnHk9Kqvj3s90p0LYxh3H4Yqd5ishD5zvIIrEGezqk+r7
id1Vpn22D3gpaSGWDGBlXI0UYYwEGUB6ydt9BaGVgmlMok5U2T9LEQ50UgUEQ5r8
kbogb3fdbffn4fk5cvROAuWfniMIWroqGW0DJCOc3JuXceGXxzWNQsf11pUIgFql
kcsz6EoLIkBiHdUj/ezbS29lqgm/Ll6GGrj0a2Z0g4x5X78qgbiRE7uzMMMq2pIv
ZFvmQYv6ySSUlI2XVuexkUEwfNj2upLyArMeFy86Ln05/FsT3rlvIlEbVYOlLnIz
QtcFP9o4S5SXqRcLGOADksGkYCkKCcyjIkAaIeB//DtNQXdRgygzVoWWfyHRscUF
F2EcWIh+D4qG/nrHkHLO1w107ccun3YonHdLO69+5tz222vBZ3O5LL5IpZw6N/sQ
4TrQYPhkPEFEDyPSNCl7BI0fIfR/6fKp8fNXRr46ya7tznfJ8kqOEX3hJxK1AGUv
1kmAqRKzTobP0q1ycStRnHhADJ/BAjNXjm1VU2+gHerRUgWBK+grqPWhoqDnHLbx
5Vl2EZeIVADrUZHdfLGzOJvtWMFwl6ve3GSphvXpN7v4PIsUstOIW0U1WAv99njC
qsILkn7JST89adhQrqZEWp5GZCs5OaypU8iqJpojPXqDVQsO1CmV8dnZe28fXvKB
BTA/N0TTx1UhduKJG/onm/zFZKQHi2IVznzSBl75zsbIUCA6CoMKP4M6sUffdZhr
LOw3mBCmePIjF4F40/NODTBbPT//hNw5Ed8Z3XWfUD3ZM1uSbni0Xny5OiHrnLWk
KaeTjOk61SvEt+pg9+JEzQ9YeLEnBF+ZVCAyOeO2NmNDAr8jAHjnr10eKHt6h1CS
AdG5TWKzm8q8sENZHHL8jFZFNefaQcaaVtItat8Xiyhv+8uy6jo1jDdX2glWjQmb
iRSy1jUBnfpac2FFYSH9eXWhzHJj2zMMhiVZCEjh3WuIuHQZiaFnJnBSLEn/5Wlm
jqxkvStHzvAM7vTm6S3jnoTmyvkRzF46ZjrRyB+ZM8P12dD/C/BWvoIvpegvPOIN
Zn2sTxdOiOyhquoxqSgK0ispeiOP5FbB9boyFv/RpMsH3ixkSRisXz7uVJ+RGbNB
zv5ryrloC2eNQUt0F0G2ZGyuZ2FIYHZ7MqSCfH/c+lqy1jU/o1/Akt6FEwzy8gaa
v8e3hkXmb0dN2kdsTHAFf7ROL+Op3YOvorF64QGOchzk5K1y7oa4EntSt4tNvTVu
zAahIF2acvg9yOM0IPnS9b6l5Ku8ocgpJVVn+dMIPfJCX7KBR8hIDrWdd8SzYjbP
NugdrSIdFb4xvmYx5b19jpFS+nJVrxaK704Mi/mP9k6NGo4H1P8vxyILeL/dAjul
DErBzzjyzQDHaRTJVvVNG3Y8BAMmGLDOkwNx8ZOkZciuCxHro6Jl9MZ2V56FN+0v
RFK38Rcxjw3AwVyagL47Nbfpd+NQLJS/V3YSn9rIf6wUP2yWEKbjfjAf4ZVTX3RP
ZiD+UFT4hXohJe4ztP1C+48533tcPhaUaZqh9ZtTvHwQQiK4ltTs96Bo3CMOlJrw
wTVmGzvSmz1j0qZHnPkxe+ZKX68Jv9hGKQ2LJDZApGCc6JzzhPtIEZW+WwHwbbM9
zUFcHgmWcMqDSo1fZtiTEf3+ohHgp4/BGQCm1mzoVMCFZS2KRHdTA0+QKV4ra6Jd
rJPu0T6HwTEURMxNs+g439WAZ5fmz/AkvQnaNFxHVpV2YTx+y8hhkJllT9zL7yKm
+5WHEmlTSuuUpw4/71ZFnLornaOvoQ0/MwASyPwWGiu5o74ljy2Gl+uvPn/agiSq
yep7IX0NsodZUWn87P9gM1fUI9lP9ojMX19YfFv5m/gPwie8pGB8w9xgD3DJsmvG
AiKPJA+UuX/zAwW+oTgQSlRo73gXTLt70/1UHroaptBCVoRSpLf4TT1c+JZbFd4y
h/fg120OQ39Ox1zkQRDkpecSvh7QUiUsZJ0BmFQ21scH1oq7BvPDQ5ydLpGGmfTy
yhuc6U+41eN1v45qNR6W5ZHJ1CCT/PdPvnigk0qtWvWzqWo3z3jfe879HOUAav84
5MrjBO2CVgNYdGlrArWSEQPVtq4DALuzD0P9r/O0aoHvOU7ZdQDKlFl1sfBmonUP
rGcnbIndOt5pbcDvxgITWaVt7RmDUwoA6FWtl5L+r6q/DRWd7ApJcNwAvoikAOyO
G2thbiyY+9MJz911DRHIEh1aXEIX4toH11HVB3Qx3EcGNK8MR5To0vO2FcTpLL1h
RMsmijGV7aGGTrjh2S9d8Xd/t79w0jPywGhkxowiY0tZMPG0ZUo4ofQcHhDo5cK5
O4geCHHVTpFF8QcahUS7UCUvBY1nt/b9ib+cZNISGRqjW47aYXEyPvFCoOe12LPo
qCpFwnJiiWCKwfE0DfjsYr0pi+68FMjpMHsf1jq74iq0hOgfz/F4qXe1h/0bDTnZ
Uzi0wNeWdn3qbQtjsGTfDDghJgBw7dX1yizT2yCK5EbDF3ggkj78rC+BoaLdETCV
tgu3gnv+U49UdweUPxWVYpnCJwXxaFDjKRGAMgJKVkOXmtBjaQBE589AKpgy3JDQ
80dH55tkYehhAtTQF+18u+h0NKUifvBjeF+jBEXvs0BI1woRt8siP67+cxSGNJcu
EPzTsRkskX1lqzBg7xxgS6CRFwhk+fuq2FOiEn/2Rp/mNNoz+tHz4qweVlEmgUKu
siLl2nPpU2KsVhzXiWekaa7G6JmptgoS0kw66JFbwWTR/Y1IF/fCtfq3AE3KzaaD
xuQkjU+TT2m/IleiyCwH+7pzkB1BKE/J44lU4QXWsXSSVYFbPBu+sVvPGu8VWVam
uikRK1jUR3KJHxIM9YG123m986bd9vbIM8JqMIDb43DBfHis/UK+iecbjiPmqE10
ywFVEXcPiP4tj9KGXSwdvpNYqvK5jvhwR/t0RryGbGqzO5GLLi5ASmpPpKM394sA
BCTllv0rCain7sjkmw+sketz57kH53USrvv4L9HdvLZrALAojNUMIDvOW+g+4Ues
iXidD+9vYVTnSXAj8Ze3GqaIYMhmX245+BIPrsu1IWHT3ID3K02m1MUTs63QinZT
+UjfZtGaiuSpXIx76iffH/aUvy8/OgG2CFBLOMJZcp4Q6DEZ7flsTolQOcWBPYvT
3hi92F1PaiuKiMXXTrP0pNRQdkicJuxyDvrmMPueeJtUB2eQjha4syE871DxJB+Y
2kISozeJILq2RR+95DMaRVmrUwDLaPsuZ4BCJKdg7hdD8TlqizsnD4B7PL0G4Jdw
hMPx8F/9impmtpZ39QHEUyU5ISSZ678m6vfLtxGUjXWDJlU/iECL/aFc+QexPsRd
/ZjWYQ0FoOKLg5TEoLLje0BiK9ULKomBT5ey6WaKCL0dvj2UR4aGbYoSW4nDGE4b
GoLjJHMfgFw14QnsDINx1WW4sOG10BFTJjZng+YZnacQYuS/9hzjxetgJsPEAmfG
zUHYmgHuvJYsEoUyabENl9v9ydW6lJfykZW6qsDhsPyhMONxgLtuSV2WClncCHU3
eFCkBogecwLBuOmTNdbEsy568QxPC4K4dBXDi5JNudv/Pq96DvdPXMFedrtrzWX4
8tetzUO/PHptMJU3jcwBsK+2EykJOATg0U6WrKFMIBMs6vXnUCIqcGZinjZKlW9o
YHb2ElJ4wLNZYofCXZNO0hoUyb3XIfminIE3eb/w3hZxUog8h2Dc9txfIcJ9hCDm
OgXkvPmAqFjKaxLvGZPeOHRr3A0VjqBSQSWI5HEKCfXqDOzMn+mg6QD4KdVlIlPp
aesi2OE/vsgZWCOfGk3+rIW+nasesbBlQ3o8EssbQyQp8BLg8Gm+hHCY+eOJAqaB
rvw5pxrsWFsDMCHewpUJzXFQWhQf15TFo0I+8K6+lPPa1cQqLFQIsVrit/jEtwdf
qXXSC47M7L9hs4sED4QltPWiLniq5dCSLaD41nUq1+gnavIBVIvy9MWXeGlSOy7J
seUUK4oC7fvJcHqK90S7XHFriEWAJ9F+VuxpHhieVjzw5n545pYdsoCAGKxVQnWU
nDZ9ZuFX6rMa6LrKdgF/WzC5S/ZmEhRBQD9RalqStXjegb4V3qCGc9dvcgC04Ry5
Wbuq+ftVpM+7fT61D3uxf2zEjhDTdHFA/M+KFk5xwwFAFXfVMxmxQ1wllSxHG53m
kHvIOqBdlga49m54vrE0uoMw3hPnu3butffzgSU+FRvwOZ9w6pdbECF0mNCM21wA
p+3t3UqrV4K5xf2/RKU2BcnS+bMXKOJkW8xy1m5OMr1ZLK4Xft05DBErpO/+86F+
ddvZPVUAh4zHP9ko/M9VarCEP9zEhUxI/7PeicpqJDQwztJm2kFKCBj+1xQ9CqmQ
AXxrJmZKFo0kDWw/3KDjb1EC+SFFy+nacLc6T2jv4elI61uZgnYoNhT9MBmnNBgP
1nDzLT5vSPuvbQM0iZCjo9bePTnjflpIQBMy6wJOGhS4KekobZWOPC3OPGJdDuGS
Jqfh114DekhldprFzVG+TlCGbBhEGOKtqrCv5wKsNAxeBDCArixxn4ix7ZtHUuOX
dYs+U7vQhhQSgjk61K01XA18+DSxRpMbpiPlOO5rqXTkG6OIn9TvZPFjVLAJiXpU
Tt7uX+ur+t/1MoXr6scOni3DqWCvdJh98eIvSNnQyQODjxvx7M812iTWrPbNN9xB
6PywoFnAG7GhykvS2xITDhKTg5YknQGq31B4kTKD3w+csNIZcmfjVUM15fsFTfUt
v6k09r/rHofhGUFpPSynglqery73YEM+VmrcQOK2DSjgRmLpv+a7UIeMbzD9lx6H
X3HXG87naEWv5nlZBUAiKic37TnChhnRAMZsx1RKP390reRIFbtnU4aTQjdPF3vc
+GR8EjvPibCkbZH8r4DRGToFVKhbEqOwmrgQLaHiRTz7qUCs+yxopcLB2s4LdEe1
/QTiBsFwtjH0bAf9N9XoiDfTTgLbimeKD5MOBQpW3gzRxhMeoBZwdrAw3kzX04KB
GF/0+XEnuFC76SRN+jpZdawmt8WMVmRr+W+nQVcaAcHv3cObxmPk8ICzm/U6CAK9
57hKjc1bjlCur+sCBCIEQyq7Dt6zY8DsvRA8FNDCeZdjUB0kuTwEImvl13pFuN37
z8Yid0jxDBtGEo4NfQy8LHpk9/c+XWN+WCDSYNIeC9/bBdmmw3vttMiA1g5F5aq7
H39UUeEPx4eKN1Tp8AYI6Y1QL6vNfrkHE8djONxNQAc29al0DkCM2oalKIZnkVuT
G4hSO8KLlVVBtdwsMeNrmQnP+lc2SVPjvvBlGRwvgjkgxsRyRs/wFlD2bhOT4HDw
t5fGzHDUqSaPmE7F/cIh/qX3asW00OdXRAo+7rCf20hb0zr2ZPNgRg90OtSj2VYA
tNhmL8h/ufjqz74T0pVg5Jd3FZNVqcS1u9zoN3RyQXKwJAD17HVcfNR/QUBhRvr9
ys9Jji45NQnn6p6LMyb+BpfUjXBq8i/gHnNkwj4tMUJq6H785ZKNM+v8BzdpCJQS
H8zsV4AEdJ/CyTdsVRw5WKHTP5OG/BmFsBo8VzqFM/b161L7yezsGbqwVy5MBXqO
0rXjavnQeJa70cG0fsoHTsEkElDK7eCTXae9fffLvEjZ/ys9LKr2TUJEIC3lb6hI
MLN591Jq+Dx94/cuk31cM959N1xy1c626k09O3BnEqCCGTDOI9Ojwx4j2/wksSXU
ORgb+YLxtEAoywu9j35q6jHBcZQPpZ8+7InZCplePoSZZNmTmDtsC7VdJflM7Xi8
aVxugqoc9qG5zaSIHBHAStc90gvHdLhqcB2dod/GJBqbb8E4UwM5pU6ZoERm9IXv
pkFOuJKKP563fvV448uR5mRnO68HAYtsfBTMymCf67kEGKrTaOnj81EsGcnDd3JY
uIBIrmo9GAFxYcEoFSs6ksSFmocwY4IqdNNRRLlIGsUITsGQjLjFFCym//1MlJt4
uKenhFLJsvHbH5CtsCSWfeglBFU27cOXkWyO0632FoAtcYHWo7c6MZZyC0xLlEa/
kqvoeq/EjJMAHX47erRG0sS0OuUIY6f8rK7zU04Yw6P5M9wh7NI41O9ikSFxLH3M
dFQEKo3PYR2L62B+BO2Kc+lAwpKf+cgRYqyNp7i2Ce7XwA0EyDcQjwTRyil6IcyJ
SHNnuLQGHoPzshYdbSIoEbrvAC34dLfw82xPvyNZjx5AHKXcUGafyh+u0le5dD1I
oQDLLfsdhS9xDZTLSDoRTTXoMNfRYVFrmJbTXIhnmiujG1Qdh2dx8x3CJ6F9s2i/
lGpED4FxF7fvC2r97vYC8UBe5rK7d+ZgWfhaci+SHarIorfbdKTzyFHD/W7bHCVs
woUHH780QnmtFzKsrzNolwHGU6yyk7Dm68L1YD/tqkGxfZwRnibAEyguZ0SXWcPR
trzX41jfyc2+myrt83/9qaonjv13WrIGujHIkQVLmt+xxPcceWLwysbIdUL2SuGN
kQPfLEoP9Ulom34zCELhpO/sAkhcXN+vWYM3WcGZsOlTcjj/tg5KQnwws0yGy+6c
2wn0jub4gAfnnxWlqMmRnMvb7j+bySgCNw1opuNc83qpafDvE0978WOgO4XD2Nel
7ECepIyKY8bvk1y0JL4IAjFo2QfQqGbBZ/AkVI2aB9maYYzwjcVLht1y6C28ZVSq
Qjp9NgGX0rZlQSssld/HNpQwQrLjxM1y12E+xu8hnskIPbLGlBR3OmIyWkGMmfWQ
dK1RLOgy54W27IPAJslK9g7lqVBMIZaSMitlfxKca29T0IAwzLtiITfyz6iMv6wq
PtDiSGTG9W8TfQl2JhzT2GPZDcXj8TOb+SvTFtg8Odc1A8Fv2o6tvEL047Kf5nud
U92GGeG5NtJOysvJr8qxq0FTyakR9F9nI5mN+dwIDqdvngX04nrWDVyN67Du3MqJ
N/L9baOK6oPzPRfD+kPWHBucuFgtC7XXsvBc2Kgp1s+CjnKv5S0un7QrkxEXh6lW
h34P/UcwHfvrx4fUegNwGq0s535QbsckosnX6L1hsMWsYBgp+S8vP7+aea5vbxT4
HSlLvWTlf+lQJRqka5YLNKUY29/ZuEEWBvTJ2fhZ8AEimhDZsdOnomZHr800Z84+
4y33DDMUPmwrZDYzC6SSb04Oy08U/Lmwe8IF2zRS6LyUyQCg+jCF9USlBiJMawH7
9TxakxKB4Sef6CpQoflnXhcLxSg6Nj17k+lMROfkai4bgBF8W3Tq3nVKTJBptyv5
7V25dCPJ4RnrELTXw6gu3d7KANW3LW+V6X6Mi3J/gS2Vyph8YuC//zN6ONwp68iD
lD4sH0WX8RLH7YdbDXwSUI1NIhGlh1cNZGE5p2YJ5MV618omyz1qt6L2tjfgS5QP
GSew8khwiCRvc7e022V+t0s3AmEioi9gT0zH8LF+/XUWFF6o4DqiIfD29CnUFj8g
1wV5C+6LLUCKQKU5B2VQ9g19DgMi2wT2Dfqb+u2f0nkv8g5yoHm45yc2UxVco3eQ
PMOhXhReviiM9/0Dr4cH9OTPZN4m7fXk412Ej0h8F0WOc1dOLJLgIpGnq0aMG9TD
uDI20y+lYZNhM7hrTey/PKR2OtUwyi0AxkJsmuT5Z9JaWtfeffzy8pR4Og+lcanZ
PWczhm4advgsLfBfq1ENY38DNwyqLryDzVagyOkwoN6Ih84DmmeKUDa/ijeqdSkJ
TZpjVBGwDPpBEPUfnJgyzVUxEl/QBGasdQJmJPko9m4wFK7qPypa6fIfnOsaPwDn
mEMFFGDnWEFqMIKECu7A8zFx7SCMc9u3PZNlxNoIq2haZF9ZGKDolE3wqgOz+mkQ
3WLJR/qxEbx7ZwfJFwfQ4OU+ELnDLTMBzfUf9yopy8fVYORseaC/YvZclN7HFJ2Z
47Pn8OG0ggMS1tcvCz4v0GfcJlXZ2GxVKhb8mfbkmmaq4mh4oFfo5ruB40Umy6wu
UKT4ZkTfkbxTXYxA2AY5D1QNC+rAWt6ZnrcPeHzcs9cf+l9Zter9+PZjEz6k0DCr
XRYXQbSQ9afLNZJzj8TdVXPDqx/jZ/RxXEbtArpwhCs+VHHziT0XB3TwnjxCkaFb
Hv8TWqtqqnyQFpoPm+5cEaycC8ehO3ZJO/9dUGobrM+iY7ETNbmeD7dWeqCuTD3j
8YpKj/0fnVz2q4ldLAPJHvmWvL7AMhDMeUL2VtzVbs+KFhHCEZvi8YmksWZEMQ8T
Ebr2eofbV4L9+zbtMiQH8/UwgMv+gCaFdSPCRaJG4TXB9uAhjXnSee7frdvVaMDn
YXu4Slcw5YzQIUWE+FayB2RkKPc8huStis+l4Ckhk2uzyho9hvzF6+oTYFffltus
a6RcfnooKos35MS1vROlbbdyvzmC2ZzR7F3jozwsurZ4HSuDdf6vsfGnXQ7r4ovI
Ka1/3Q6gsBwEEOGLGjcH9ElQsa6tAj92sXREXX+pgkFp/qmCIDAs0pLgweCpa3e2
D3usPsXMkg8jqoHSM+V7zfhcbCJZXZzIYtK4/jcSJOYAm7tRWEDFO+oAV3NTP0RA
twEv6nheocz3ZRPbpmnUYWVXlKJwdB3nvM01ok/+aLAhD/pCIcvdv5m91WdQoiJU
UVPQUBuY7nGumM/9mDWLfyKCDm80RIIWQzav9VqlgWOAo57KXgH6yCaKCs4cXj3m
uBVFesvN3ndlSOUD+BXxLqjXBDbePLNu24dRkxoaygrjkwhjxuSHdLMUWdaviCOb
LrdOG3fmZcp0j2kR2r5LtrMGenLc42iEzvhfLfmVN5sJW+Yamn46FwcEahepjSSr
Idy8bO1mT0Hx5Vg/UQ6c4Dl7R6CFDGkOeOY475HPy5ZXs6fzycyfydID4ivJt+Bn
hPwNmYDr6K7Gr7hB+O/dDYjQAIsEyAqiX0ILJFsAFweILbR9hVM0RaI5Iaf4zqdf
/LqSat8Zy05fNZcpNr8mOUXabfqj3r/loPYviyEBjoe/9yt4QuBMspNBz81Tsneu
2gYF8hR7uTAR4o4e/t+gvxWk677UrGLg0EyCdnL8tK0QjfCNDHJv4AcPTZfF5yKj
E8wfujcuOmu3gK1q+57VW5C0pxUW9I+aveaXyR7DG6LiXGg+tcoquR6tggs1HQrv
4jYIfflxM7zvERRHF5ilHCQYa0gw7/0/yofuNnHVNDxAh/zOD2TasOH3d4J8Zxz3
+mM5OCL57UMo2vSbtQwJlskZmfS98I86wCUcUXPp/2MDVWY16TQ/QLmNmv0W3d1e
2jTBz2PDMp7+S7q/ShDL8YAqz/Ubxy/zJwH87Q1357N8rRDeUa98ZxsTE4JmMJI4
QNRR2FJw4t2ktcenWTM/qlM2pBmNv2hBjhPghqTOmqWXmbGxD+/WfIChOZyvyTN+
iqX63HVYUhdUkFotPMOKObr4kAkPY9B2MZHr8s5GtQ2BfA2CxKL1Y0yoZmhn/RdO
0Zm6eDeD5NO5KprKMV29gGADc08G8absR3QOp9OopwR5DoJXdGAIW9FSEqu6Wx1x
IJ+XpAk0Hj0KipUUqITiwxDMA822l1+UCfpuhVFmsT6j+nIWTMUgI0iuFMllLDtC
WjRtC9au8y8PSFvQgcd70xGcYN47wgGk1al+Aw2K7j71haGK4haf9hBwfGEQ1qNT
j3innvYOXkf4H/AOa029tEdFoQvlqioYYEuDD7KWEk+w2b5NOv4qo/NfAAfnVDXE
K1iQHPuUQLTx2AaYDlq3NnZ/TFpfZf3V0sGqRrMVtD6TzyRv/1Ff8n+LeGY9UL+P
B084UuaAsaFh1+PKIjo+dvDWiAOLeqfso43nFdbE9QpipdmjFpW56iifLvTiBuuP
PtNNjhdIb0uCJ9SkNDxUkP84f4UFfDgVrxiTbmZbB2+EVp7qBUhuk6xZmvliBhow
4tLJ1oY6T8HMEzySZjJFgO2jqcOS3FvpZUfRF3Eg+cDBYiMXBoGFFLUACn+GmSmh
/cFZgUZ2jG8me1ksrDirLjRbl/MJBp3bJEMeyKS7U04Q62g+zl6L0ZuJybZN/EU3
bhT1qqfIa28QEtQc7qW4QjACjAABYg3zcu+BNSmERX0e9U3h79nisFee8qyOzbeR
YjyK3qTSDjVBBOKgGsVe+JRqcAkFkYuG5wVtvPy0q+QKkVc7tSGmtVQr7B5egm/y
6/rx7IAd4rSuCGKjJThSymhIJxOcO4H9JdQ3kQbvx2x6s6uJiML5P6eDKjKSt+Pq
DILFbEatMkRmLUUs40gU9pFmO+6w5K9u3V+ajD5RPM5UqKvFNiPjgA2Ad2dDdMYk
L5rLqzQm+le9Rvq32tKuLnXBLScDyQOF9pnyOpk2fyAkjJX2JeK/dCBf6cEBtWb0
FFNLIEceB/deSUDElTiskgqCeYPcuxYUPJOKGu0OWHOMaSyusXEM0cYo+oOx0jzA
p2iISkl7vR+7qhXe6RO4ogzmMoyryVZ5CZ059EK7dyoEWDYtek8MuljHCwxNhAdS
k6A5/4rEWV14RXl1mRi6E78YWIDtTgfbuu3iHM6JDhc3VpPRhxzZiNKnn5P7dFBv
nFFPvjXtx4TOkuUwoi23HzvlAlm9cb44eXgUdf58YpS2aoMSCr53ekf2SKqeowyb
/GiY0HlSwZD5PnqaczptBiYJUREtKKTJRcDXEB57RyYmx0YFqvm2ew+UlExA0pOX
eNTqo5vxUCJjpgEZt03tOwAmvx29159ooZWJwFZp0LHMQTZgTM7rqb2fs/UPOvaS
Yc5J58kKnXM+u644kN8NkDKjtInVHGKnDt++PD5+Fp4cGAvGRh23MobmyLMiQrSO
mxYHRQsi7osUn1oy8NFXpA6bW/xzo6KTatnZC9Xfdnn3Uob1nVofKDFWP98xDYVS
3NVlPe9AncA9wCg5lhM01aBKp75WRXpXmee+Hs4G6h4iRmKVLOvoBw/M3VYUIqPw
XNXa0bW6zWDbeVWFeuJLz9uvxrmjFlDvnYQCinFTVgQMuSceNTgyZKL242xothWf
t+wL4WAoi7JDT0qbInJ34TtAjRtlyk3XGKSSXCDCFXpFeh8M4ZEmgqRf/F1N6LdK
bOhqdBGauSidyOxBmhwPd1GMgvepuYeqQ4aNFazzHouiIN3bZEMwC/muaxwwhUPX
HQ/LVVUaAyzda2IyAPvg8SK7SVu4x7NKjbfxQHgrKICUubBRnNHC7vhbw96NHOgp
z/m1TmDNDVm0bU/7OBl+CS81VEgsWb8evT9VRpWdBpJdz+g8/lZcmAzjazgsagnE
lcjmsmNf6ri/elEz3ZubAkeOSOOygvKwqM30m9FSlKx92ef6EFkW3rrdnR8OQ3WW
ONOY1FOavHIKbhzcrEtaJ7ed91UNj8rUgmEwnbwy7fkVDQulblM5qucMOUaIk4LI
+bOGCTRRwjXFSmNit/C8V5nqG/z4XjqPtZvbeDLifiy38sSl9qNEHduoKrxfL3g5
lazHWtCqjZuzJDtxgfOxHKv8ZPavgysKIv1h/m4qAYcF+ZFWVl80xBls5kldOjsf
OASWAe+zC8BF2N87NBKGYIiA8BtGNIyCyg4/DlLS3RZc5NS2uYUk5fFaMQRy5/39
orzNN/RdimeUSw7fLtbgZo2ZAuITGGuZAxcsz+W1rtAfm3oBGZmNNDEkrjt9RiYw
oD+/eQA1o5iO77MZTaLGn+MfW8YfphTFsvyoK3TuyQdJuLTcsj29+Oaqt+xKjwHc
Fs5WI5vogSyClTffWpqodb9JX4vipWDUmz1FM4Q1/28DvPVGsQvwVAO+Kne4TIur
U/HUzUaiIja3bgVnA/YAIZc9XwAxSzBmGE7YcImmacduOTJxLzv7GssjiSpi3FlG
IYk8rsdkxJMyytA7rpdObMzOTC+n67MMOkTBYa0o3ZSuKhyCcAtNV5SuTOVFLtP5
dp+PFQ7FVCcMB8GdNq+iTU3ADMRMIjxneBqh0fHZJKP6HXTvP2X5y1XEkYARxx7T
LB48GEenC6OsWBTHpDhmxrnh58TJ/5IOtg0A/Ge4cDuzhrMikzrapMqZcvl8VR6y
mObu7rZ54pFY7SEps6FTkrvNACEtET5cmJrRwsHbCt5f0r4nUfDm054M9DnsNtYp
J6PDLSCq0k3/LCv9XoDCn5KuLuRA3K2mASbvHwwO8XJEH/t8qpGTV0pj0Y6+ofqZ
g7QfBlgXSttHye2vu+nKWXUScM+/BhUkB6L3M3aN4c7gduHz/hfDOggMiXWP1u3w
q+CCmNhSDe/vwGnTZp1zZmLIGXq7UY0WgsAQMs5pH3yVKEo6O315FgqGFm6e5uJ3
ZQrPMptVG1DaS5+oOFTWhGqO3olYkwEuxyjX4L4M8OC0pHgwmW9x/jHwSbd+0tar
2iMNeV+KzKrXwH2GhPBdDq7Brlj3naJbQoxBMLWXW074wZEMsOicmikZ4xOtdlJG
ZbFIRMoAnJ4nZ3qzKyl2RN8oHfyihBp51Nsq4k2j50J0FZkvLrl3Z6Wo0GiLuy6B
qF5XU4Z6T9C4V/FYMivzPvhUvpo6sUGgkyfFdQPVNu33wEgHEXpmL3Ocv8frlk49
7otcWaKXI3bLxu4KKjjOiKNQ2KRQBLegtNKBCeW2f6GxVCdMaMA0t1xYx/Kv2KS8
QuWoptl5SG1qlo1lXSG7FAIQr2L+/m7onvaNUIMbt/svXX0lwOoYe+esLGYuTmTU
oPUnw/Uu1Cftw3DWUgGVfEGNkKVHLMLh/tjQxcUcSvpJgZ9s5oOvvolhdRYTOCVX
QpvggNoMJ5iSWEAfHRHWTiYcoYCtFxSL16xGShFexWHlCLe53ihpns5Ijo4tHPyQ
8XapT6Jo0Lz3S25+B6dXvqIVmef6vVUgJWLzlPdkLhWdJmdbkju2dBvFhen/PsS5
epIdZ17ncHBaETqQM7+oDUHl/UXPQJATeR9BpRckd7sVQusnH9qV+h4Rm84Uja16
4AW3OviNpK1gSpjfQTqdtBKHarpEzWSL2ST5NKGqUFRBJ3HQyBLC2OIo2GvJExJH
bMu2m+mwGUnLKrLk7x22xKWGey+skxmcz4RiiVDQhW7cnWjwzY4kWxXUjYXYLAl+
pthROWGuhR09Mwocxa5UlSSrVchWmbAdW4fjbH4k0yEk9MJJr0CEG7T2gvyuqQ4+
mpqJwoOkKdUI9zXSLHlllnTeqPk6hx2gOKtLl9em7A5z3E8ZgRqSmh8GkBrNjiYa
CRyN2qEi3ptwbXvJUeKdmN9sAfKqUrCuuZDEvAEtbJiKA2imPiVAJSmYpthFv+jx
ooXTY9qQ0DPGYTPTxtxQexHmNCqnGCl558W+S2fkoThEM1i1jpWZFcmjtwJjM1ep
yhj1SixTTba0DI3D/3zceAEaxrmbmONeGQn3MidHd/PZdGgDh/+YMEMIGlGVgVjv
/os6LdaW/ABfFiZ63XndtOr5CfyJ8/0ZYucpXSXipo9nVQL9rfegoxLJVN9Xw4ku
KDybuHKNOBR10I2P1wvZxb957H9dX5jbb1snOmGIYAFAxrVzImuHUsWi1sLnczIn
pejpE5b8pfrmjGiANvpCcOOiu+DGR4qVZiN78MB3sTQjUZh2aRIdO8hCwhIWbBEZ
R33ijI7Pbcxjr3arhLWacGBS1jDgc4kG/64Bnn07gw6cLhwpBN2J/h/KE6km4CPF
/UuoAkdut65IHNeoG/BzTzk6PgTAf8qepSLX2/LdDB/wLQ+MPH1w1gDUftTyn3rZ
w6o24cnAPNJ1KQ6lFRymXD4bECocin78lXRIDWIxoIkOVanEvQos4c4erLC0qZ1F
MZmn41t3xtMVVXtGdT2yModVUh1Nm2CRS5dOF1GXo/jOPabz8HHnofUjVDLfIEwr
9Dv+DHwkk+EJDQTy+ZX9nVvPshRTMYu1kGhtdnikM8i1d4eeM2rGjlIxGWb0gCwU
GI/GAbSN568fvp6ZfCnxdkTyixXpD/ptHhA5NqqxYQdMdHBYrGJqrjvsyAVWqMuX
Z6VYZxsHp7gQog0VZTC16htZIvocyVWYdoidj+3EIpNOI6mb9ykcjn2fbsLzIzjI
AC2LotkflbZcEEj+FU8b315NKG1qVdgjxxAhpYaPThES299tH3Ov+AZGo1MDkPgU
7cIg+qoDF6RZI33cOh2piSo8B+gs+9w5yQHwnAeLE6F5pHDeyE667SBojxHiXokD
CR7NX9OEb4JNlB8ksSE2A6zC3HfxSVknxilqE3AzYV60dx4/UxdKdIOBOUYyb7oT
Oi8nzRMjAXgHw4SLR5wWk7YofkiHn8x08CYR6oZV0DXHL5ExeHtCZTpIFduFc+LG
j4XHXaTA3x1sCauST4SzVTc3E+1R2xAgm/I2boD9eoetq4EM4wq8RVu8E/uBUPLf
X0SficLIxuwuOCaAWrTrrSKTT/x3gkKAExdGiV+JS2/DBZ5057EE4niquByYBm1Z
gNevaagufSs4Yad0k7jvm2nsyuwBtKPTdqKMjybY9JYaX28scVBSea5jD6pufrtO
25XRaNYaKbCEcTmnN5wVsTnA6KXZChpX4V7bwZqFLNZuVPkU4/WBI88y/RAxGWai
/UD/Zrlm5TxuFJWo62ruDThVXWFyreOhWgbnPqVivLAZzU56Tt7NY3pz/VunboEm
nkjG84FPFuFMLzG3ebNDErMBTiLzV6+ErjzoD91dD8QXRRhDGoNUwFZrx+2ZD/BF
LlAbhLzCcJfIhb2s8I8/f+/iOx/Ko/zAQGJ7/BRibeE94Erer2/k3Om46luJ67JD
Vb7OCXo3sugPAxu8V59pKPlWXX0+R1qM28m81lKmmzEpGnNG4kf9tGVFTK2v63rm
eJ0U4RtPFJrf56HwVb2IrbGH3yr3bYGUGNXH6KW4HgFSAEgw9eqmgV/KRTTxZ78A
38SZL7xuTUETxwslNDI+UUzDtRS5VVjKyw6szWp22WW24cBrTnypMxu3f10FE3D0
0F3jkxBaOXbKnAlMKLMBZAnwg0wH1iwyeNN0yd0UlNw/omWfv/x563l8xM7Wcn1t
hOdtmbhifw21YkFb3GkAQlGl6bal4NOrz4gNbw61dODQSt1Y52rXolyFLFhfCaDL
wHo+zfWZa+m+d1WsIX5CkVgia7h/MdYlQKpDCog9offe5ne+BZUQonTrvLLF5dv2
vOressojhzIAMFGKnKBWt/YTRb8+xM1iEunbA2XnMR7mKV1GwZcQsn7NOySXrvGe
3qgPvKt7r5yAExhOCn0CM0/8U2ZECWoDpi42ByaCeaKVbfBl9jmTvN3AOpZTkPuA
H/EtpoKp7OHGnp7H4ObRrr05Pe8C5oNQscC9s6kcb+HO8+3ONmSO3QidpJTEmO2C
dnC9jawVjUfQ6pLz0nPH2IKixWEcj6N2xRMLLvg6DWck2/DvPxxODHT6z7Bsj5SY
DZeP/k6MZhOk1DyT3UHbK9Gb6n+NBsWU23wT59m6i6gDxw6Yasuc9Gh51tVMD0iz
XpHnWSOcqmz8G0ZNFwNeGFDp9xUFaLCE4h7AjoT7JdTEW0kQjR5lNF2MKQXdiWUi
qm2ILnWvODWnjsgXk1eaYpm92B66ZHf3YIGj/ITpe+hw1X9pmsAO3sfnw6zRnv5D
Z1DsMujzjWp8yhI7DbpaIPT7zLmzRQebsna9v7IFGQxcz2cCuzfdSS4pjfLWL7D1
dkA2kWh/P86I2wBn+ODSqDW8S6xGo6PWL4omut+hHxZB/O/dlIhJVYxzWY8ghtSf
GunvjP8CEjhlhM7IZ1kCDTCtAvxEjthsvnqtxmUnNRLKDFexJG2XIr7PVFvhlk/0
vMkEu4NvM5dA55ACxio7Zi8uGVd5OVVWZbdogCZhRKpYwxSjGOk8D8D+MALIxK4N
HUhDgKqih/cZS0UqkL8m7fyubzvxt9sf53/PxNlu6gmo7dh+hKGTxxhnbCSPNIgx
aIuSDB6EHu3Mv07iAmYYZ+8NeWSS3SZpKgT6162Iy4GR2fcjfNFx+8Mh9KFl6YNp
MPZC+eANenugdGkNjZaADiLNA5CW/PQ1ybve8pkoJ2HfLPhrn/7I6tAJl6PXTkit
8knmJhwQJ3XNjwatVJ4P3KuxLPTJMnvsG9UEKR5aY8XB/rbNlqg26XCsiD0uIzS3
qpxxFuQpyfIqxQcSD+4juXsaMBxlTey8THDE//izX06aPV6r/PhWVpDDU/aulEqH
1eOhWYaqCS+jySdW+QH7e1v6hfIqQniTiR9m3s0ZMwfrqHOpBRytHcdzSsu+b19z
d5/d1lRClyGIfY+7LLYnDJBtkTsIctX/I7Pkc01dqOk+iAU2YgwBdaSb1R5zNGz4
DIMX1t0z+n0G471JW7CnSJWGfkmiz9BydRxdhHh4v3V0SJAuOGY5kOCPI7TAXr3z
aVKFHc1DMx0QQp0QR1hd9WCnCiq7OEKO21MRlyLT9ROFEk11Q+TB4/dS+e0nOumE
Fuaaas6cyHdK43t+dKtcDA2L5rpMb0OkymWW6XDIehFP0eH0IHeAAfsl/SAqlSvh
guh1/8l6QOn/cf6KCQpGNE18Hb+DgBLLguY0cD/BCulBXQw1PcTl49IkmEXweGN5
K1dsireAu6aYM098/i7mLUiO1b7ns6hr039rESlDK+EPZRSgObxUYBmbQ/vJy9ri
oKL+6ms6Obc6DooJ8OHccBkWzKgpmkZSyaEgMRPgkuYGaZLaQtatnE6PvAK4saBO
+Uo4sO0KtSbOzCnZmdU7GtfZlNHkjbj1Tg/jRAy/lJBVv3KSeKjXPwe0ke6SUJp2
5wRydZEZMEnhXFxecK6/zI3rHJeqYX2J23RV8m9d/rDkaIdw5+mkaA0dBw6UtInD
dBkS9eoscfRn2gqqJvkY+bMdXg+zcTtSDmazSdsY/0iWNZp9ndX7XTlIiWtuitMr
locNoS3XUQjNrezACnFF/kCMO3kJoCR6fn8VKQ/hkt0t9CUe7lMf6ODdtR+KXFtx
3Yz+z9Oq5bWVRfwVk4XAKZuz+k6NA++UTarnSFh62+6w97VWyDmLAnBxGT2FQtDQ
x1oZijtglPHxc97TAhncnWNrPW7Z+2GajR/XkGLm4RkA4/AR/j3d7WPLszVpYaPN
3fNVxuL92cDDDmucqPHpKGQYiDZigPMVxMc7ZUJ7h9uBu0d4pXcbuBsK7uJOwfF2
d80PACjX2z4s316LB+DkxhzmRaK5FsJpQKvdDIC2ol9/fKUz6t72u0jFDLfE7wmE
lM1NH0C+I81QL5T+DzhADSt+hnhXqnsu6djeEtgmdldzRzqjB6pKR0ldLPue/JsT
rrFLT3HX9KDsaeo4p4Fk1HZvgfO0kuJQzyHLkCb05goEoa8op7GNutmPwNYa/jh0
7tc1Y0tdYsoz6MQnY4e1ANU1jTY9caCfW8GRZGl2EEnNktsQHxJjJwpkqDk4OzZl
q66OJFq9PLkbJ/BHQGmavuVSHdAssdycooio1I7wuvJY8lMGwhhAwxrEMF8G4hBj
3ILl0EdMeqgpU4D+FroQcVZE77D0JQ57094IUZpRRL2ouUj35WEnmoGeEmG2OP5/
hPTIZxeRN479IPSKwBCEI+eQytXwpAL6rbZfflEJFQv9QgCXnzO0DSLoB90ocmCB
7Hj8rTXBb8x1vF4UP0ZyUl2S5k2ZQX1sh1aXapVO6qevPNwnGEddOM8JlyFKqVBI
YfyEfxXm+0UFBejz3tZVM5H9zkRQ1uFqwfB5GLf7XIWq1Sfs623lnlT0YNlPk9CE
QDJXLcbe9tGFdxXXZeX8XdkptC1bbBKOrRTDXMgJEB33R1rhVOWzToGwQLtTcA1t
+O1qqNK2/0iWp5Rytm9/3PkZyJdoLXqKBwSNTmbYz7NXI0hU3JMQPVRKVJMm8dSX
Go+1/2mVZhtMnlnBnK3IzQZQt6Z2NhCN+his6ha+x9wihQgY5qyK47cC3s41UouM
7SNDDAnKu5i4LTOfcRylOwUx1qH/iodc0T7DUr4oQJ37Bocejjqjme1muEWoun3l
bE+WoOsOD3sVPqXz7IkvoqYlPGXJyXBtc7nHVVCiWztny/XIQfPtuOR3kJdDpNhU
Jx7I1V0fIK51aYK7wQqRcdX4zrxDWxQWFYygE/Cmgb5TryRV0ZKioAoW7Schrl9F
/g9XjsF4dw0YMsnr80oLIT9bAfJTn7VEumeyR3NwKsTwT+6Vx9Twf4FeHc1RbvgU
nzr4V20uQHHodNIFxRaYezPF66WLwCeUuqUSVdOAJ7MtMURQq3h/U0vsiOJKKkw+
aMPjJszWfeb+2KYVJvZnyvV1CV5+3GniLHLOudU0G5EM6HsX0+JqngyauFPYnOC9
ZFGabLgkxy6blRF1yb3HmpoD0Og2fmDHCR+PybuHzankPmyx6HAR6PKrgFNmZfug
mKWF7RlxJ9qcZfZksNUm+OGbh937gm8vZEnOpiWGqSljSKmFhl6wNL3MTWUUA2H0
/n3BQBHlLUnl0USo4ADaw45q4wqakPTnerjBTNxCw2/OT36yUhB5ogL9RWysEU/V
mFVOfbwRjvrfwpNOpVUvFXD55HJhpoW7VPcXzn6cX6rL8BbapY14iy+0LhJiBBY0
LFlnKN65bcSZQX5vmJ2sHj4tjrIomHvjYxgk9tj7+WCDm0yH3wlZjVEVH5ON4VkM
Enlt6K7cMmuPj9duZ8+PcDGc17zr1wBXWk83lXBBb0ymTspes5ejj0GM5UkTLJJg
uCLoeh0Wxm7eKJ8u6xFMKyHkagwKFdAS9sOwiaQIng+6WBdWE9qWZOnu8UTQK5mc
RF28WDzUtG/PZeB/NUyjT8Qlwtdjk8JRGpHtmGL7L5hyGO6YCAjvNNbNiO7RYNEo
oLQP6aO7/dt8xJXHORVML/qgzI1oQeoDc5wwEmnToK491YgO3C0VXWgIWDuE0wa9
cbCk38MNrtZQ+xXCQ2nsOJ9O7ZJe58dSbLEMF7guCGpQVDE5aeiVO+45JxXslefV
LZ+jhFDCeVXmr9gfa926FWQLlFnNbNznrXFbI6a0zi54c2uRfeSpMgmAZyUwIvC5
Wwh4xkbPodKfbeAUfIYo0T5ODhTXqG1ucv7BR8VQRelCC5wvVIB/2AaA5HFQEL/L
nSIMSqwJ7TPnrlfJQKMOKmJ4roqAOzMZqD3kpzwgK+IMPjqfZ5CZVO9CQ4tde2Uu
sO7eaMRYlxQOR+ah0tb/W1G4H5n7gPloVA8o1fzO3FnmUd3DKFjtyt4yV3uEM+eN
JntZ5uBwwAcym+HrvGSzhL4BRM2pQjW8LJowqlfo35Dz1IaydbdsTi8iHI4LFisz
kuJJ07haf1SG3QQVQgjqQTa18KdqezRCnqpah+FZHhNCWklpuGCfhS9w6OMGbUlm
vL9x2JAbe3I8072tuC9KkOXVaPadZOyJwhu86rtjWMgQa1RnmyUmA+T5HWmn/LIc
m4E4mOwjwYnmWyazPxMbjnDbguD+SmX0n8EAJ9RlJEwFCytwb2EeEv2wRxY67567
QHQRPNTmVBXTz9//xFbT9A2XniWCzh2kma4K//dS9W9gfjbLTUv3UKvrawgfTa6/
ee5wCiQW4ZHpAvUL+eL3oD4uWnWjSOPtx+p7W6fHCjF4gqIfbOTsCwcED7qKTwR8
fG5fGXXn88Y9wc3w3XHZ47lCmX09XSck63MnLSrzrhCzPT/ZbPyOHwFk903KaY8B
jUgJcKXNEfO9h6h0Z3/9u8qFZWzW5NcRoMkyDc16OeDuLHiWA46vQ+ezViweEnN2
IuZ0u9GtSRQrWmZWlQb5Vh0LDO1FWNsXztznhMbeXfzFxdO34OJQHCOfvLBOLac8
qA1ZMPpX/EJUmj+L9m2/GO8fPnQeKmUWV6HaU74t0Y4uhjN3BhPXJyZQ7MHRszHA
11iANqoza3EGP+GYEbuCSyzQjtjhSXXqzYtWWonG9myBBepycfRUZFcdgT9tQocx
3sjgU6G2dfzkhVb2JwX1JA4TDLknJfdZWjZuJf6jziq9f/WdRNzaLoK8TXghd8pU
t0ARYT1xIN2qWDP7mH1K7OxGy0QdUOp+uLs0pCMUAEkIil1tYZFGEMDGQFjaUusU
YikGL5efnDpMP7vBd5SQApqW8DwRewtbD/fdMZ/VkC5ni7+I8kJ6l1fkP2SWlp2/
Fy0qivikA74IZuT3pUIajN2Vl7hzYlli4TOvtr1ukf1BJgWTye2TWMFbWD0hxVp5
1Wmaw28RAM/qkKEzbnGZ5/hjpjBsj2KaWxjj2cGXVtaDpgtltdT2m6kh98QXuOAa
nAAPbagNWlVSC6jhHe+YzFyI3Ju4qMd/5dnjZgvfxlddh7KuI/My46tVSDt4ckKA
irMCYW0DLpetMlSfYyQlC6hDvIM8eZhhN7Ct5oWle0Bkvdax3jWYj4GDQmd4/qOd
3I8jThEaN9NIa++tVD0Pf/T03eiZA6XeDz5NNiNj4DyGnElWqOle6YUGEP9NRSwd
1AH6NhRIo1OeBTJ7GmiPoMGQ5vD9zoTrIDpIRva5h0lM5a8teb7NmErqXAc1SIyD
uHQUPSTRigCKWCzNpEf9CX2WhU4DLIMOoHdbjBpDC4c5qYv/551vWG+dXy++Re7V
2DmImh+MoG6/jBn6btOP9+6ycKSaK02TiXnjfrMQF54uoRToJMFZxQbSrHQch6BP
+AKcUUOjItYlorEO/MaP5uUpDX1dtrDze6/OtIkIAYZBFhVP+gMdoklahm5rdA2q
jU8B9ytPFH0J87Ha48STXDsNML0jfXR/Sz/fPjG+iqeyDW0ZiPeFhkvwPPmLvYqr
jpn5s9XnJXMb3ec5ARhSUdh9drxz7TWr7dVixGlgIJkR+w9g5XsJhSlX9vrFSDho
h6onhEC7GCUyELiJaHp36B+vxdC9t+q3f05/RnhfaffE4SYAoJlxEIqiHdHIKMpj
0FbdnTaweaqORQQcxC1rhs9OtfVc0JyFv1RH+QsCJ63GogDFHdlVPLn4z9Rp7Lre
23+GGnACz3MSMdE7LK9E6JJJsnItrYjBcCEzIT2W/rZsoPmxOK6hYQuyXCFR8NiD
2FTaL5NXNxFCNvv9TYKxteRi+jTD4DVn9X9to4Kt2onIdXbnAUehxvNOpx5vUT4H
wUqFTapefT1/Vix2Lo5F0fCDB0hQYOFWGGD2RFPlc38ZV8CWlYz1wpP736XzuT2K
1GvYJMyQoZ0hxSkA+TMl4PxL1LuZ0KMZ8UNogVYc6ZYVcAGElsn7wNkT+i+f2nDd
ZxiaE0PxjLh4yd1i103m7KvdVZWi13PaD75NNoKWszD3gjvXe0mPnFw23TDZqIe1
2nElVyIwcxVKvUHse9R5pWhDADaIy6pHmlYlNF/bdAwTjHzEkfjiQgkTWS+6oNSp
FFJJkbpc8B+++dd++z+FFeIcv2h5nDU4UIx14y8qedZux1tV/g/MaV6+DcxFvMq0
xgXps/MhNVKsuPX1Tc2iEWPN9fwjHmQ3AyofpIR08zww4aguFrdrCy1+KAB438/T
xx1REUZEgFl83ssWWcK7sxmdXX+JAbn8um8VKMtIECSozgkV/GjqiMwhzQu+lb4D
G7JYmZcTFl2zugKN6ZAq1FOCl4S4BB3dx/JenZiJ8GpI/4ty/Us7OUD+o/TQQIhG
xe24B7aeDLFhb7QOczj/AHdveSMWM0Tod3j1KqU+uU5gsVDNCTKWeQDWiwIRaWZj
8JdtXxJzLDpqht8b6Ynx1asVTFgTvIPgnIms/dd+ViFRNcYOgcDSDnVuk4T9aWAR
z96123xkjAfHZyjBq6zse51nCH3uV8E3wdlR6BJPVJdRrHVP/jN6Mb0Ck4JMtLCM
cpHHEMSq03jJCvl/r8F9kPyLRgrs3HROYXYX5vP8klG330UBD2iF6GfwLz4dru5F
/RYAleoTsyS4akJg3LEpdqMKI7XTdUkxj2vMSqZJXP0++jyzG+gygJVXSBnAybwu
f6yPXfpQT1btrnbNro2FgR2/k2YTYy/01dM7nZ+wsU/TVys1e7pCTds51jCWf1qI
0uFVgNcTy0Fa1PqTJDB8hD5Wv7Heq3we4J2heq4PegF1WLA6jGzk6uY83p6GK5aF
N7d07VcuCp4qWzycJ0eG1VN49pbTygygtibdY56N8fiD3G2SiergbiQGFXgFX8Sf
95Rn0vG2cKSdG1A1LXg5Nih1IDe2dObrivEuaIa51aoxrkrUD7ED8sjlELY6S9qK
yKDrqGxXLR2veYSpPnWED6a5lU3/ckWOlUlGVNhU2LgKWN6Gq2FDDn52Dn9aeV15
kKQbiFAlZPUH/KJ6E6w+k+3JR4V6WJH1/OHrzt677nzxQMB8eZIwlntBR2V6Motb
vkBOCMdmzxoWPy0u9oS0zzTSgrLQpuDpD9ck7EwGPy/vyfrSKmXsdmKtxcrziKQ5
nv6+1yEaYpG4LPy/+mPhIvh+j6ceqtRWqpgcTwVsCknBioCbNpX0//lU/Vz/ljkq
5gJxk/p+IxvWzkNH+5Vwlr8+B4M6gCM45zKWJoSa23Fp/edwfaR2Cg9UrBssps06
TtzWSuYxtWeKMEFU5unz7vzvjpErmi3JWLE3EMgH5/33W6iC67USzPkXidphKhQ9
ddCyPI06De1yTzjJ2n3xy7U9EfF1iLpCkY4iqv4mBiLV+7nsSRpb/ZmqtmHW9K5X
pe4kB5/fP3iwXtBU8GrLgcLQBx4vT0cji+HmzA30aXgpOXM2cO3XetppgCnnYof5
zy7R69En6zP1DsKJkgeqLqMm8CeIDb50Vx7/T81khZxpQaneIhOSUPchYCrbBPjU
D3I9oR+wauwbIDQ2ZfW7rp/0xNJlOrTUlu3V1jgBM1Fl1UB9ibZIP6/N2dC0DHpL
uH/jjm+bV1pxnG95rAyHnVGLyKeAMQ1P1I6TCiNXP8YmwOL4qEULaPfzQnUAZiEV
b3vSTCG9YrtN2j/FnEGiEXmCfBlJdIF5hm3LeMIChX2cGmnGRVGzfR7UR/4TAbSe
6QaAlIrdYUhH4NDlFMP1UIo5CdRZDfKf7P5qLmF8kKKeTlsqvHDY4ilacg3/LQlj
WpR/WISxiui7hMZher85ouImZ4T03M1fdBh4UowfbOJ5rYZORV0WpMs35KMVCg0z
RabaBP31EvHzbSspYmwgz1cm8i3xDpwuHEnpdDl3l9MQJ/bX3q1vQ7ZV6nZg+9Ft
28lCpusjMQ11CmFiATHeVfg14R6O4tcmc4ipa4JnCL3VtiJeLqIStkH4tEKOtVMd
1/iT8w6/rYazku9uNIUtD1mlsjlZTWwE0mhXZCjK1MT/OB0lxClGfkloalDFOu1h
IUZLwggGias7DjHpGtcPWFjDeziCkRiAHMnthOyKP6Kpops+v1dpSp4LtYCRtmq1
wSHzljQlU38E5dilXwsfC7BVrfEwjhSTxmdQ3oJAqwrt4lctgOpO40yNDcD4+c8G
N+SGx2Woi0kDyfyLjS1sQV27Fv9W1pnhu1XkbcjhQPJychukmqSf2xZ7QI5urYqt
uZgdZvOcojZk0RN79+wyqXQkGqeqD4UpHTAMBXpcl9ckKoPG/f5P2zCeNLDywdJS
rI9SbsxUpZ3yVYtCD9jUrqlTff/xroaNffzM1o4HU7cfpo5nKCvJsJrgIX5JKXAI
S/WEUPp0orj0UGg41C98sBQ7rIYlXbIpiV14npnL3NwWQKTaAHZOlFZoBDDZHssq
QV1P6zVgKd0F6IQea1tnYKYIkzMBHasPBD/kt2QB/3vy/xw4Zx7F+RwVlSgtI7GH
aJGI2JNC0bZo0lbmbqAf9Of8vgVidKuIC7WA1JrZn4vC3+2IdlaTrLroEr+wrQVc
FLgHuc7GENDPDDj7VD2P3ym+uD2BSGvKmyjOPg4uprYNFs1o0OEXvje8FpWfIQTj
1cMZXpa9yaJR8UAf0sU/Ov7CfG/WR4eEd/xPcHRmeoNFjAQ1mo+xMIizaIh4UWwp
djzDIwkq7d1G81Ghw8iyDX/PEI3d5BXPsdM8nOL4DwJayXSZNAKh2+6TVBFFJobn
Yggm7RZqLrcjL0hsJsC2zfhJLlB0eYH/l9WaEILdxIlfwctrLYEBg0x6QJibV+Vq
jp42vWSvbfJVdC2eegoqDpK9A0Owc0ydxudF5YyZM/H06qbVXtEAOyYn8TNzloxI
txLpcJfdVBcD3em07fvfnzG0aVu2wP74wuulUoS42PNHnKXQgWuX6DjSqcgJ1ede
RafbZfDvX4yy3L39ZVTkET4S1LuP5fHx0FdLU3QQ1ZtHqju3xwkRC+o4fSY9y6Tm
XK1jUwby76yuLcc0eIKeKoPtZIVwXDu8nkSug1PyxPrUVGojOZbtrO+EYwqSLG1i
iUBqbk0n2KHl/q+wiaDD8b3TTr5enwwEzDImoE75fk8eO3xKOzi/qTupE905vcFq
/I656MLsxTxoAasIY8aGFaSCymgxn3KVYvNrHqDFE/nl3NaPFuN9ZDPdDUrwBsJa
H9lY1NZ1P8QteMSp6oDQPec0eAlfCY7SZmT7JwjNXVd3F5kN1f4Un0pshV/GeGdU
wih2PwNzssdMn/DD0RyJf5FfHdfxx9EIb2dTorBp3sS/bXEuRSzVXkyvVTTXZ+RI
8NumQcy2Att+nf12uP6GgpNxUOLHJNLQYd3Fvnhr7u5G8Pa2mHtPcfgSpPySWTJ6
WRLS4paA0DGIaP39PwwJ3IiePJWN6CyJHY7bz5oxCm5BIWHr+jpKS0XBbDXA2Y6T
rfwhPIYnqL3naMNxC8HuAnyPNLccPtfsze48e1/cRERCZh5c/lZT3CBkw25lYMnL
xbudLzATMyIcucBYEgxYXUQqOIgsMAb8aEM5NCF6PgxQJd9VCpakz9VQpOLvLPlA
WsBbjTGLS1VBpEC5y5y3bto72PD2sIR1NeQQ0UUuqaxb7MLoRajD20oZsGOcY921
RUTjeHfX6R8dyoH623KswPVbYjXB4QRM9PPUiWORKSXUH0t1EIxUV0t9DHVEEaxa
x2v7PR22Gp8LDRIjSvg6HiDfxlDZ/ZkKWx43hwrUY6i521CPRmuwX0xzwV7HJo1m
b107gdWY+1gBXN8/dmVYo+DgvvTzlgvnGYWQbsEx3ayq6jJS90Y1QFXUpLHVJ3dk
FaAZZGxcZ90ZieaGZDlaPVzK/ji0Yo5/myY9bCL1bQX5kpLm366LE9pPXZEa7Lg1
AHb4u0yHEOl8qu9ZBO5Y2LryUX05vN72cwxNStzuRG/Z0D8UU6NGfdCk6ZoTnhir
8UxCyvznBDWOihAGBGmp7PGGvBqZjTWAXUt/fbXedfMtRacsjAGKLsfwueDSvq3N
07BgRUzbVglz2uJ66s1GoCbD8jy6nBH5cfrESire2LEhQrBSVK2AxSQZ2RgJov0K
yaA7X0CXqemoKcnouwrTA2JCt2rQV3flskacZd4zlhliDSIqi5fxEhLmI2Ol7t00
NRGnBpXWRCIMcZgIlhQsa7L3l7J5TvpIqe2jIyppWTm6SOQo7XAlbF+0rBqX8+bk
UpzxccrfZYcKqgIrSZdJ/0uEIbUpEpJIrdN7N59CKVZk28xt8mdo3VJtlyRyFgTW
tY7NH891dB9VkHPcc5XBJQyCETynHCvFfW6OWg+0aZtdgnICmSNwjMtokK2wCr0I
mmPyazFc5b8jcug9CKHzM6Gl+3B3YvKrZpxOSjHeXYxjAIeb65gjh6bXa3ewenOf
ux0vyIO5xyc3OzulHCoyo6PTIlAr7XN9O4tZpLdMhqG1R8JxUM7WuDAkZhXmxenO
rDxPjBbSllyt6WPfnZ2kvG/gZPIa15iQq0sqYNf38y835pypQEdx7eeXgkY6I4Xd
bmrU9HTkLsDaaQeDU6cHuftNgYiZzo3RXTTyMJKOkGkcqmLN6VkdjtUedE6hr1eP
kpNLltP3Uauva4Ojz6bnglyrJI/sHBI6moBySo4+ERHcuiyEHW1p6oRI3S4LkCt7
KVZTpt7lGExyE1cDkq03/q1d9BeUYloDxEhYLiPVVd/MKwu0p+7RFYP7U/LMGrqF
fUg47mZRoKkvWFWAuFAl2fn7YEzPcXiOAco33RqmZG4iCuY3Bff4IrTPRPB+9zuL
Y6oKAnE8g3fdlMhL+aq4CGhRa4IlHBpmUvHu/LRalyxPe3XSy/HFLmSwOz+wQr8T
p+6k9SgomlY9Da63ttUq3UBmRnyjt1DvI1m/Kya5DV11JHIvclQFD0a/0nxOH24b
Hb6uzldNNb6ZQX5Zkv5bXSWONpi9x6VQ8WOj2PJfkJsfbwwYcz7AD71GDdwV1jKe
0rDdC9heokFH2+CuPE6r/V5mi1bZPmlRZUh6ScZn+UffGqQr+5sgdvf+tKhf5Ovo
yMxVrfW4OqVJgMZr3tckwZt+U/5dixAEpKQ419gmcAYOt9u68UHq7pR+LzKFRDQl
WHcsL1bG9Xo9o2Pc8eUslUkMFFEovOIZOfblstYXiCFNY5DY9NoD8PgpV/nn/QJr
SYee0BeAdm9Ga3tfnI8G23OYiXiiHrcO/4r3nogW9MCwYTazu4ZR3LZzzZovIMkF
OTWLt2hRONhwycRt0U7wcLCy1Yn2LTw9+2f2w7dCjxYBqiWGxJk/s0nNWlc7jgM0
J/Q3Yg+4PzGJjBqp7Gw8Z8qlf+qB3MA1Cs8fjEYacjOng9ZugA9H3Iu03EIRPaDI
vi7XcMh8VjdnOK97MOm+JrWU8jGFBMragQu+zEsR7WrdXQbN1jj9VqeGTyaGAAMm
kh4XM2hBy/SlIkNCHguj73tzrQPgZMr4ffbeil+dhjbOiQ46XySXh9OeSM2oLVsp
xFEmrHRD6n8daLCaQ2uk8tb2F4u2YZwZ3sFa3K9+JibAK3nBlEUyjZrmwGKc+iFq
AR+ZUfNJXuRO1qjn9KsMV99vPYnvgtfWc+/N0KvLGDiei+/dY+1dth0ZifYtmKBi
HTEEG3MzdsY5DEdy5HNt5lvaSg7nw/wBXZwpdpyxQUyOK0io+qZFvL9+Y+aoXmz4
caNlMnG/UIsdqT7dhwoOQSVZiGUw1ILh6TSch4UUshT/eZc3uD/9ePVyAnSUOdfc
ovhutMFql/SaReBRzKwDWlun/QxHGCGb9IvckaP6Tbp64SJzYY+IbMYykxIWms/D
aq3/m0UVFyLrzTT8CDrB+T0+oTO0diQ5W3eYE+UIeqhuGYgSzPj62Up/k9ExBd2F
W+Lh3xYd/4n8j/gMZQWp9G92GC8XTK6gkeOGBImNT3yngOA6Fnq08MbQQc/uHbME
Xh+fmfyegrZ//KE8T6S4OFDjTb8E7GAaYStOySqwRwO/rUyKdBAyXJHEdHK0qEwE
rkFfg6coR+yGyb5O0+/y2iWjPxgYIQB2H4dozD6UhrFlpX7xWwUQQAQcdEQD2byA
rbbdYsZJject3NQGwc4TBV1+y7NaTpNRTnQvgFIH0wlnR1tVqeKTNExa53eo3ALT
1WCtvf6vTwBMM9GGd1zAxxDjii6T8CBtXQ6GzdSu5lGqkJFS8+8AGl0y4aWycFy0
b+F5/7P9NWxVEtm+0vtWT2qcT8ag83sq4ml8VYeDdOmm/kWbLf94voo0uo5XuLYj
FcoMwjoSWtmEM9pLWpQvdkLIsiMiWEi3akBBbH+UiQEbT1agmDHU2BgnMTDUqlE7
i3yW4cUPi6BTZ+KvHpGoanyrtfVnnA6JzPXD17RJnbOY75C/CFLLZYQNMqyZ9FWR
14cWryCShgyCIj6Bus0MqA5bpyKrL+EffZ4DVfD0Om+uGiiSvs35SUhRh784jlO1
2p4a1v8HQeXj0h+8XMpSqePALu9CID0aGRRQlLzxrnMfboIPTjsAO8Zl5jwVAIBV
co7O3K8PbXlwQl0UXYK/seTkxrcvnvshHJmOs5LJiDi7P8t03xjNChdC3hFCE24g
0CV95EJqf79RevqKUu/syvaP4k9EFX3GJHjDyDPRb6fLtA5cpZbUCM62N1q+49Y3
aEoMVyZLWUTiPps7bv/DyLzKESNE3aV+c4DhKXlFOQFOeN9rJ8haq1i2uyugJv9E
w/7pse0CiozYS1nt/xDAh+74AVJHLbr8Baz6Sf9Bm5lC96Y829IUY7RVhc4WfsuS
fYB0jlfu5e0ft40B1nAjq6xfok6UMUyCdg4Al15yZ7/p0TXk+Sj0cqkr0T4GFng8
JJr+50+t5N5uwipCVW08hj/VKD4eh8EPjUa6C8QwstBWMYyne4yQIxoZAYFujWCw
tnPvPhsZswMhKrLfzNCpYyZunyZPIChUsTDIff3bOMusRl3AS2Q9zCfipFYv+8aD
nZlCQJ/nstE3/OgYUmwkwoI7SltC/u5LGQv3ROVzZgIjb9hHcp+PrtmRujsEZCMJ
K2PgxI6u7wN+105jItRhr7aLbbVg3xOvpRHOTOL+rTUId77SOZHxZT2MW26LbALR
IkJhMCwt0UB408nJRR0tCMjzwOy4VTB2H09ToPamZnF0jmD+RbOodJj+9U83OaFu
TwbT/7J5gwZiu7ncy0DuZr6EnwvlgV1LtQknpGvMeTzME6fe6Iou6tFXA8zNaZ7s
nouBdp+SLvq4oPx93AU/0or2sClgoVGxeSfUlNAWhAC2Vu06XiQvJjlyZgA9Loyz
QmVlefpKk1UuaBvq3vbwVaF5usUjy0+yf/YbRF8bmpDJQMj6W0baYz1PQaYfQa0v
O5C86hbQ3v/1g3vJTZD+ikGUBvHOy8idiUMB7BzkBclKUXh0bx9KgIRSjsc3bVNZ
eEdDSyWbUpgvEwbFVyBLkWX8wSDc6yCXwTb95EIQ3KcVY32J5MAM0nM31Qd8fGbi
4nLBLodtdjB3JwdYfpkYB72vHkj7ubzn8fe6YEmLfkz6OuGOpQ4+sSz1zZncu2q0
9I8DIsFTvExs134C06iRxlHI4KBqK9ZFpNldlbNdJuCRKQK4aN2LxPdc5jAARAeS
ncJrFWCLzGfafiekVqvcHeJf2VXJCWE7pOGFaMJo/fMIgIMfn4uNOCtVfL2AhcjL
YaDWEio8rUzmBfWwQk+ECv6QfyOvjSYGegNacfPEt53udLTZSWg6wbTFISBisgpu
QW4xaeBwN6eJZd6Okd/7D7u2otNJ4zqSIpV5LxGjzLBXfXX9pcsVU7cS/HLMM+6e
sT5T6LgxPeanHsCIIQXj9uoSmk8C6c9dEFoBWeiDWzC4oQQHFfar1uz9QDjeZCm2
7ACjncOKQ93MmRHl1Z3Xsf/L8tqWVLaLoQCiwyENDLUppokaZPYVPwT4+6TvAw/t
YwzN1/h049ehVC6cY4NLWN+jxqX3EAbfI3plViOEmZHwt7FGM+eQGi0eqc0GP8TT
azMdlkwoXsW2KbMENu5cJGQ8u0/u1vD/nmS577hdeXWqqKoeOKgyFF1IgrD/G1uX
73rOZlJ21XVKJzzReU9mpgdFQpF9A623FnSeY/gyC+cnPiEjqUWXGqB7Li0fCE8k
3Cx6SXumUbVT8BnZaXfeyYgj4BhKVwAFhC6bl33nfB0pjBUZa1tk9CBW88NksZBB
IoHk3r50FWLBXUvRPIEh/clliNkIO7KPPTVu0vcQlXUQUBHmTYG2eDGruKzRCRST
pP8uZ6axx/fd3PeSgEruFeNrWYrQMTcFdZaxwUp8eRj24U9O3jABw/y/a05D+hg1
RIOkNvKn45OLooWfqgex0/BK1AcfehERGUyV61sq+Dz/CGPpZRMOtO/eAvfBsIkz
ZkMeEkX+rHQ7tcQiicu1cBv7yEY/dI8iPzdkv7D6q/MM3BWKp+O9zuNVDJpmZoz4
PX/LpwFeH29s9iMfvN1wS85une+OxATA9bnHPiKC1Z1u44zUlWZQ5mkA2o0to+e9
HxmGfOkiQCvBgMWVNmk2FeVnFW682skfXWiJMdOmXNDBz38ySk+RKzg4oCzYQyDs
Jnw7WD4+y5yXvAC0vzdj36u6x26uzPjmTmbJJoXJJXZYqk9fIiYUau6h5HlvPqr4
bZqwLH/U0ebr9eouCPI5QCbj+qBaPZw9Or6+z2tCaiygtFwqhLzkzikwwxQyS7L7
5K3toGEtKDrDinzton6oKHKdmzruAwQF50bmkcY9nA0JwfOWEBQP6Kcx7GNHfeff
vCoxwzehtwhP1eZqOAB3Am4s958kaUTme5vWhNVXuahBhb2the6SgV0xIKelDPxS
1CvM/veP62wAhclOHvVF/vxJRW6Gn0ay/OHhI9lncuetEL0X7b6IG0F2kY+rEAtJ
5GB5lzB2YXZ6+2PcfzZs+HJZ9OnzkyeI7d2j8S1bR3Yz6NZ5xwcOq9yVAiL5nAVr
LQpcs76slOKmnJElw9Gd2wTDEa5NzKlY8FYqSh/3FVgzDYvn5OR8eMQqUFTGphiX
oola/pyjb7o8nO54dIgJWL1wxwASY8OT8aKp2aZ8YgbngvIbQKM2rdt+4reBvRCH
nOyBcSIyFBiPtrE/SueIko+gzK9+L5W1dGuYPpfDiqvvFByRLpdkmf1ZpEAEtnQl
fG529BjJW45ozZ65wIPMk/y5h6IdiAEvFk9fGkPDl3+lTSIKyapgzRUyaXvTTeSq
q0+YVUZjcN9bH4FQX3YhVmEQnD4Tt9gaOA0OlGgt/9inFgee9WvwhSKUblGqIrO3
kAOVEql3Y6qtRCSegkG40GSkQpy6CzJHe55Ei3EEdYc0LkOFKhKiJQaLlwsc13mV
+aG9YCjrAxJukKBUw6DpRIyKfK0OX9bgW7C56xtqY+LvMS9y1PkmT2fY3V0mpzs1
iFh1pVOKVSLPlSIdp10Y/TiaBO9X9vgO5tIs+TuZBFVlf2UCJlProZK3V/6hE5x7
8HLGcYWxd4sxXOKyPOdMy3Me7uJycKeWATJR84QCIYCRsBE09dhU7t5rNxobCUcd
LbbRUMBMrWaTEUSZI43my+ITVO6q3GFkU60h4ugJBJujHsW6cXLKbOBK8I+6s7vV
WGBQN7LE0y+u+wQBIy07ymAS2UoG7jJiI8sd+ePUsgpLuWZDRGF81qs6+dOjlCDm
w3aceIw7EPLkwxji8zj/X0lQd+IjfQ0Wqs7Va6/Sn3OccNBTIlQgG/xGOGduWZ1S
q7W6II2PW4k1Lt8kTp8PkiD+rVuPyHKxSwxZRzb4vSjxYQGqACotYnVpF8NOn/Wv
cWVowXOXDS4Dz2SmMHEyjLc8tuA6vU9r4Vfx1FEtpqDZ80jG6XL97yWqEMIfKWbE
UBtZHgGYgvAih/ujcj7FMvO0SpFba+PwRY6EPsHtxIbsbpQ8ssos7DEiB2WOHP1y
A8Ky8EBRiG/38VphL4u56f2pwBoZBgxmVAH/yaqizLMvDAidH6kWqOxVqylMR1KA
wmXOo3ReltzUUvl+x+VW3tmryAM3SeqJ/QJOhsbqcOEIPpf3dR83cHg7mq55ljHH
+RUN00vcI4oXq9AMWzQpmeKliYyatKZGcqWm2mF1yMg+opCyv5Q61x/pndAlaeCc
4lDMSnfOm1dOYfoPiCDH2857pKMSNXgNlj+5JYgVLpMSVHKUkU1QJOKhOA3uBJPO
ZFkvEvcmioEEWgkxY7ycjNgdIDD5RXGW9mOIsjYuHCrQMKxfLYxRT4G3nHRBTZMI
Jlm7YpcSDasVT80B4y+kh9PHksFZmtE7blOEWvWW1t+cMZ83gw7RHq/88A6wNKqW
dIX/oCNc4qcGmfDBvjG/D66s4W5pFIwMh95mHDVdewp0GTYW6EJ6GLfzxFA6gOWk
q9ph0w3GKrlV5e+c1DHKk4FFRKBNhsLOCWvLlJ+35kVnFLXyNXUlZel8bFc0h4Zx
FxIY/T8gVVB/RBgjG+Al0FAe+1PfqRZleR30fEDqks4YtqLrW8l/AWB7667XWVkp
ULab/Dt59GADj008go13iapF5QqZdo7mgjQ6TdpS8nKSzbT0p52oDCZb3QZrNmqL
laP7nwYhmIOfGPXgSvL9t7ltoyuCLza9rHNQh1nHAWv/KXsh2VOKqkg1KQiH8WfP
5sih4NDNA1XCTj49Ycr8NzXPzmJvCifuGp1c7Y339ZsAs0SC35c4rwEgFjcu/s0Z
b3UaRQ7xHDsQqPvYgCBZdNbx/1PYnUfKr+9imbtVHyJylXn8M05JHa5KRz8Mua4y
lgTnANPQVPAqjYlvrTOi3EpoJLx7lmyhO3kynC/zlNV20Emw6tQcsvFSpL5efOoi
FiEg8+L22cPoFKflX7E6Wze19lR1UAOz/tGUkN7IjI7ke+ntIpLi9Kpr9+B2aOmY
uK/0Xwo2GgCflWiVwOlOW8Gyb7F/aV8p8hED0RH0cUQJQ6Oi6W7NFpgu0SZop2sh
m5ZmQP7ZhtuO0mHPGXySV0tac1+nv489PipsneLDWQgCkw1sNf0Kyk8lWM+tyE7d
+YgEykENbI2uxTWLpQGtIzzpXeRXvE2Azqg9KRpoWX69egMSDEVHPjV5ea9zs4+S
20Mk7C09kDlGweyKorfSkzj+9FNTaoI+zGqSuHv1CuXDSm6rbwP8l4d2os6hgRaK
8nxYKFJ1ZhmO86/R6ZRtLVF1l+dJizCwHBnFMvgN2oYZJ4Wh8Gy693SfqejMT1rm
n/6th5R4pMPe2IIMEXsd9jjCN4LrEDypiFyG5SVVugMYhAmcgqoKRlzf/AQvffuA
0UufmIw5Li7JcoZQeLqeR5l0g30RaFfBNkAZN/x75xRWRhgkf3Z1Zfr9sZ3d+gvf
ota5ZfnzZyeu9t7q5r5iY+7pIzByDL9iyyFzXhXiQLc0KhQHjtrUKcJvuMwp1Hrl
+fHOZ9IqI3Xe/Y1tqhzm7wuXuF1MiyRReH9nshPe3WoQRDpiMVfMBbRDX775N0O8
s8yAIjLzK4sgLZtXjyqincDqh3R4Iunxd7XdykhQnsGK++C6KvMKg0omkLm/aH3D
CRsOLG/eWUl3IYl3rO3mbuC0yCMxjqNJxrAr8FSNXScSqCzvbDUpOF3guWuBgHSB
WjPLVgJh/oalnBFH4pDQvN27ehDUsK0NjH47ZhojgXOKDCTqTnojTc3pEizxNWJm
maz/gP6JZ5oZpk6boaICbsxKcEtwgIBeRgUmjhB7XYJUNbJ9JJ2uhxQ3KPsfvLL9
0ardkRsexr5fSoryW59PLYwRqGAwFOmkKSPhONAq6g0tA+KetsPWIOPV+WyQK0KV
rqiqmtgmOgQvS8ojO4I8GYhyh6BAMLyZREtxPWeRtleFQkxFejznmZCz5A4yiPTy
6PnmC5LufjtzSbRk/+3I2l+tCgHB6kKk+vVik/IovM27YlEvZL6hSEDrLv2Ro6MA
hiR7UAK5zux2gSXFtvVgKXhEcsfaGursKdUYaPBQEnnFTgjQRM4cpRNzJ3poQXVj
6SU6rchbF7uelbtKLqIE9LEhCfuQpHEsWF/6C0dD/VCJo3XSC8m2qSGHee/kM6hT
8g/xGd7ItYY+6IwKRa4eb/KGHkPqi80dL9lEnM5jxt6sgKh4icE3dP703+3N4/HK
9t44tWcxjyceCeja2cQQIoJKZ/9DHOUU55ZAfCnZKUpol3E+PSbHxr/ti75zHiuC
zK5rGdTfzD9HSfv5Dc2Em52N2UsGSJNI/tPbTgP23pMfl9DkHKva1SgLSvqOAUWM
Kb6dTdzGs1VsyjjkC+9jsqVE+L/BoTsI4cttyUFdB97vo1pZcR15UC/ryriHODZo
ynxzKnSq4vcMVLjK8t1hFBrJ/T2oV+3HlThxK9qGJqQkUK0PnvTer5CXWDscAevx
CQIgRHy32Qi9MRy2zJu7Dj0LBtdJiohHq/71mIoe5ZsZoRoXEeIpjpxeeJFrnpDx
tu+bZo1baTyHrQWgahhwo1TKiwTJCjiwkhPFjnJoPCg6Y+Xg/87in2mlA/BAi5Ya
+L0Z3kjnOdvl0B81OECSKj+0CMhSMdL4M2k4mWIaFRittSQivBUCaaPaOm/9ahN9
JMUAfMPRIB7AaZbR1yVApbu9qqkMmGQExVvGgIamIRiEKWxbwlQJPJPPKQDhlktp
tzvgEaWFh1mXIXuRHeDrR2/bHJHfxjNWPtre3dvEptd/OumFm6300/sB7Ni6tuak
oTuMyF78CqoGWuwRQ79jclCqpJsTOEmo+6FcDYjRcijQW1mhWLJckfoZHjbA/0sL
uiF004uD/0vFAxejgx0QBH9XovbR2PasBZNaY6vq05JRzeIvrnQNXtRti8udbl48
1yqJexxi4K+7gICjrOCyxpe8pbj12Eher8QkEOvFVdsw3/l1i2SW7PFX73bjzpgP
67rBQQ+LpjL5F21XgIYx0cUvuo3Zp2icptue6+1pcPw1SzzfLD8nnLyWJo45jCHK
AlXOWhJYLie8FswTsMg0nlY9EInSHxslxqShA/rtcGP2dlRr6zeAyNzdPNRfpXov
qI+wuIDjd2qGc4s7+PvjLn/Z9V+dhewB5V92sHLKXeui7gtsIk5WcLDi38usrBCu
99UEZ4FC6/ki7G6pWj+sgVhgTdSok+DAbh2iM47D6/k+V58ZRvLcBM4ZIhWo0mYs
T8+UfkK37+15yKnxIXXVZ60tIMsvTCGLmQlel2FrtleAlAu9P4t4GnDmPZKIRNCs
F7XKUuVdExzHKDv5GxI1RbtXrDaqItG3i7O9EIb3Y2lmtvHCsAuINFnNO3EmybcI
DODkNnecHIKVEN8/D1LQVh/N8mhLthAcnWdGYb3Eot67VRp+iO0YIjXfokF34+Fn
tDdnSkY8qt/9sWsJZnx+pcA6O2Kzr4kZVxvPM5jmtuqDwSl58GGTqQYhVjhS/pJI
NN60l6OMaKfvcBdme2WjCgcN+WdgaINy+zl/lkdnkslXDUx8HR7GZZcIyHYzb4jW
cU4MIRwboNK20FFf/pHUN5KOzoH5r/MXyZnqQxnkcsi/Nca+KBSUkdYZ1aiRcObu
KGrS/hyTrS0v14eayNB5rcmDsxlSYESN5ga67umySRrdsUsRyQLjPG81nFeefrSJ
teAUwXqtBN+qHVteTRZYL1W4IYiE7kh+xzMZMtXJHl69kMYTxjn3XhU07f3XmtaI
z5TvVAFQcn0AoTIJsMgAYxECS/mSlmoBmOUu7AuKSpWMM9ij/i3171mdqHwwBtD2
ASR53kJc67E3IOBJ6Oedt9lWD+YAUgg6MD0boeoZ9loZ5ybTLRg2k3BYJ2F45as5
Xaqs0uQYIcjEpq3arcoQ53c2ABFtlHJFxkqjIsUsZ2hQAbC3d8HVl8Yz9jHhGBec
oNmisUiU/rs+3oZbrzryZHBHOZ2RY1idH9NPCaDC7FA3zRhAcDntgHAot6fa2Cge
Ro5TFTVbuD4tv0jq2q1QXAF2Gzq7Tr3fic615pbfMNu4md5tHv3ci/gMI8BboO+4
Y3D8nSOLmplED1M2ls2hvUyPGMxXFUiWAU+ltwD6Bj0SH4FLbAR/mNVigHgvI3OC
nyvw5j4xxc5yWcteV7GhYowkM9cIp0cnXy7V4/FSGfELc98jNtPjSXetdV2gwdeK
UZGyesAETMmR1K0L26Kc78EDPMN5XqarnQ83HilhMfRcuHRy7N/jaGr71CNaa0z4
rcqnJ4peUG3mk341iRrNBCf/tfI/ft+BCSiKUcJcZZgpZ8P/FX3ygNXZTO1dK+fL
p21AKwTXxlPKFpGnw/qspoMgMxaDNraZHJkJE9XCHbTSjRmUj5+A+l0gkSKmbzgg
OSsleYTgbOVFRdBg7WwSHQSoBPelCarfs2J1BHJ8Uzjpc/Aj1A5z0izvXJStchrG
Jt3aaQEntROoTHwpVhjWhmXh1YZl1hHXt4ISXGVHwyBQzbmxfGqhSV3lCblgRzS7
KubtqIUR4mKDoqvG78mYcltSygzmJ3OxUer1XAn88gwZY1bNN4ABWkYJNibg1BXZ
xORUCdRPT7WJ1B3ZlUg7V3nBknMjjacT2gspJSnaycemSkKv3mqwY0Z0l8rtJV69
VGQ+KPW4f7ob4chgKdJCq9psIBGYUWiEGStg5Ttj1ELFiwiFbthSlYOg/tAUgGYV
RI0IlOLPL4SVF9b8g4mXfnqBYuUfiBZXUlMqnT003tlKSXqe+P7CGSLvXu9PK7Fa
+F8r+vWrPwvgDSTgOQzrLDBLSSXauv8Qy7tPDyt0/N98zQAFK/qAagGue2ooR782
1rR7gATaXaVHBZuGz+mzfaW9tqJYe7CwNI62ZzcQB9w2Upd4vycKz2cS+jycwdJs
eHG11uHzF80P7ODF+XPUrAkE67sslZWFTIZF/xt6J7EQdWK4/CIz4xSgzFB2eYQs
NYK8npwPIZO5W1GfA2HN8pymBSe1T8sPKTVKntcdM0I1cyGGrRbHX023KwS/xc5W
pv4H9agFXVsDUS+9LWlBzhCfRF2Y7ikrScMNqH7mM5815WBsulOXRiCGc1MofyVl
ueE4OvVEuqEs/R1ua/lVVaMiZ/tgqgDhNMf0Hd7cka02EV47GajpQpiRNdVk7nfY
DdaQOqah7jpr5yT9kCwgcPmRGUkGHiVnxT8NJy6fcBMvMFb2Z/0PIQ4v/4v7LR+p
vxT5xx5bzYTioeVfeJvy1MAXaEo22DZBAu86WfYrlDz4nqeJQrmnpjoW98g+yp2C
gbb1QYhvQ6upjbTZEoEROopiOKsBiKUKC89VghUsvW9fwCN7fG+0gh1pXa4+MWnN
aUbsKbSHsZMmiaJiTeW+3MtSBXQFyMXy1I8QpcC0myT+yOAg9FiosFc6nqeaR0Vy
tkXToJPGauutp8Erl9aNaHDor9pfHoD5EwcCxQdY5HCQ3egldhjtBrdPL6ZzPE3A
9or+IMvR/qn895c6IDHTN9xePyIFyJ/Xcl/eHTT299vuTCYgXHOAd2pkr7dTpX9L
B735YJ+j++n2E9wCCbWibAOvuN4MoGx4LYkMUJ5NCmiuj2LLI91crZo5cE2IIbXl
+iKtWjzuJGhAZrpkZsvTfnCNew3iG3t1Vlfdh4OL5Q6a3GDVEq5phhrGRl0EQp92
vHg9SM5n0MSfJoeNznzP7N/7ADcpg64ipKijztnOke988IxFX6LuxRcPZ46rk7Sf
DoL2Ty7+h0Uf4AxsSWZeF8VhjcAXKAzsHgHg8k8PZuczsj9w1sUWiBfyxzdymkbJ
ZUTKkZZPkWrQJbo+ceFLZ/Fv3eygt2Vc20y12u7upXDAA65R2SIwYvxMd6+w9R7y
p1N7zpCcKl9e4hgFhska629/KqyzFuoVlRgOWKM1VQCugVaM2y9vtLaAlXAuwtZ0
YLJC2DoKNBmy+SDqdIRyGtwARTWFropTnVCHQO8LxrM39RJzgUx4YB3aowuJiduu
rVRb2OTV0Fw/24/CGGg7jEE8sWCyNwP3WVdN0iG8F9xIMEt49GyM+KPT2Kx2876v
KeySJxifnyZWjg/7UvA5Yo6MJniXdfxp1FOC1gfbH9G4UXx76UlWojejAh3UcGLo
Mp09E3wDXOzB4MQ19g5/T0mxfWbkjYpRfWbgwM5G2g6OWw83oedIA+3xC9BPot4O
pBV5RFRLI8lKFHWab0hN7gbpL+2C3dawRA5zvy44dSjUrlzm8dt/fOiAJL2HxRy3
TbRU3uhwAlGXes/LVGj/vALEMwHyr51csatxVuODwKE0DYtoWNkqWfcYG1Tt4x43
otIYUPKjk3/zv7U+ROSkbYy22ffJG5m/m4rTCoj/0Je7vc5jsQr2FC1wyGztDTAN
li28A14IYbc4EErRkYXzPRpFwMcNSCvmZ3LEdLBo3yyrWHhGpkwv3CSg9O5pxfe7
OlM0S+zGWXTe2sHW1bxdRswfLFQ95YuybYsMCjowrRgZgJlmZhpNmPUaAy3bGD0H
vkb+IxhAt/Lv3McdrOYZjy1Z+/QNGT4ngYrqX9IAx3lK7E4yMVkDaiiulbm3+Iih
TTGGAFDD6KvbWoyB5QbfcyVDkIE7DjnyIc+236r79Hx67B/RiA86PqYFfQ86P7I3
nvPhScECgXorrBSVtplDgqBlIy2xkyjyrPAHtjMl30x9dk0PTaKbKbveparSetdO
L1jiPkXKIrCMlewX8EUxSauV7BswU0zjHxh8oeb6FD4Amx3IkrZtEuHzlPlagt0c
1LhXQENnpIN9nTbAOa8KoQfesT2PbEVAagBNgTCF8L7PkTk/dQ8+C7t+u+5Mp8BP
0Y1Llb2aFLIjRQcUolHVb8lunDFGqx9DBBFZHnr+2lrcZckuTjTNsyU+qHWBGhd9
GgI6VMQlSO5k1U2oL7FBX/mQyy1GxnqizjWUJrjc4NVHe2Rv6pj5QFG7AdSiVC0s
FvpoHfEZMQkT2/yNEJO9t1NPMZsNSNII25hKVUp2neKe+hUbM9QagKvN0+c/tzTd
lW/EFe61SsEW8f1yXOyEZqcHaJOceaa711HlVJB+ZrX5/BVQh1sqbCNh+U1YlsOo
fwukSzBUhhO5Hh5ia85eBpksJqMaytXLkDIpXhi7jshlTaYK9p/oTAVygGYxs5ru
j69mNgQ7EVdEj7CsK/DtuTZeO399EP9FF5d7aa8szUfWemGbntZigyLnFgxwyi9S
OKOARQIkAHXn16nRSFSi5vozjYTwP/N9xYHw9auPC4O+wNKCFc8TzlEFL8e5scL4
YQObtic1niZFF6rxWKFv0kRO6CgWnNN87m8G1sLSU0e0LSXn5Ut3+WW25OwpjdBu
j6zVF3zd/5JQ3owXZVVW5HVLDzbkMQNkjMM/ZXxCPPp75dqF+j/zoT+QcAs2q/0V
sSJg/sTaQGBxpC+rJrpDpBrbgzBK1/eiEB4sTBjUEAsa3yFN2YUTd8KYHeVayPfE
9iW/FiC/aan0T4IH28BwTuFgP5dBIVzMzZMwz1sp0r89iIWyTJhBUnC6Y2XXLBFV
p6LBx9lyCjxrjIm8E85w3h/DjqrlhejhqvR7Pj0EIezu77XmldOyjKuOaIIEV/zY
96Y5wpQt/9antztQxlZKJsDsKypxOuJuw7Xvi34mqYpwm/wQABYrf8YB+GX5oiJz
0aJdgEvnx5TPUZvab5L3xZtVClNirDZ4+1ob7gE4/kosGl/0eKUgQyU5AIATrOhk
x2BsxODYBX0Wknz0VMZfI6hVhgQB6/yLgtH5TeTNzrZYMgWDNYStKvugPAN5ZyuR
3mUoaJdEP8fxau15ZkwwcJiFzpwoneUcAy4wYxSmT3i1H4VkEK845stl0w2vaI7X
s2pKIhulWHIx1NvFZ4nMJ53qwmnWAmUjNVh1GXQjFS1kBOqOfjEMg4ij/tyMzrsf
Fb0nnS5JU2r7e0KWklwyOkRVOX35epNM1/XMF2S4GDDqUnND2V1GneBXMc6StMw1
LCHGIjvHNGvGE2C6o0yEhAd7Vp+z5Xh94n7Rx14nbysL8GQBYUwtedHF5UEUQyoW
wI0i6n5GFuisH3x0XkVRo7j0rc1lQEAz4Uu0NGkc+OpDTicErTn9tfm/xtB+CKAE
Itt4YF4Xigx/MvHRzXov3Fihic4oHBjidAA2p8nCyvKI3uovOddy6rnfTUBc+c51
sgd5yjJWBI49UxCStph3oD9EspcvnL2u9jJ0ZO2+PbFrgqirFUUNuiXUJigETMMX
qqZc5xuS15mZ4cgxckZqdn7olvQOeTvy5VcjxLQnBXvuu3uKiG62CAp6mofqJTFZ
3YHdfparJn4jNTnv6KNdWYpUX2iReb4J+xyAK967gf0GqZVxVvKIxus2GtJwNYfA
YpgnAVrSOvWk456zEweTLSd0VGJy3M2OHyj3evO2kGUD4RxlRZZZCsgdz6/HBrS0
kVHJd0PY5WG27gyMoJUZFRhxm8YfvjPUN40wKd76GVz6O9qG7SVRMB6P+VHpMzWg
q56a67UlefiOHm7uVAIvfv0I5cbtBxON8+DqO+cVWFgJZ/lUPU4Y0tP0nHBLA4Mo
ktBlCUVUf5tuE9bkdOusH1shtX00aNxFahsQ8uMCThKjqlslsiuF56tsydqZQYPb
dnRzDFNTuGdfqyAHPDeLeY+Df2Cve+ZAa6Wa2ncfk1B8pl8KZd/M91LMJ6kaZXet
3qJNp7bgkG8WJCLboe+nNLfAFqd3ZLuw0wV9Y/Yw+xqB809QJ8pYilqaUAwOGA3V
JB/6SDcAzqrSp5WZHp2bpC4HYdOiaj1xOmv7WO2OJlGiKsSd5oVLFkpqwhYqKIhg
d/D7cmY+x/8l1fXvi93V+nDMvJ36kQJCi/PjG6FQwW66TAq4Bk3jwxXS1bsQy2WO
8jW46G043M1nJ7ZWo1imJyxXpLtI6nDCw/1ka3KSNHbmcxD+PHWusF8oHqDFfaw8
njsvax/vQx/4lqGIlvLwkj1TKVZLYyFpmSvBWxtXSjWJP/udrVGzoMNmEXZ7F7HP
gEDjQwP5NUFNuueKan8EjIw9TIyoKAkInreLx7stsDiqj6qOh0Rv6mP+0ryu9AVw
3qqJtxttWpM9MkIIsDbMCf/22NC/PXwM+hZOTbVzr7V/XM3d8cOaMXDgCN0TpX3d
FBeZJw6nO9B4HwQ5CbUE7vm4TWKp53UUQkjXAEIG9F9b/r2uQEA2Ao8zUqjiBm6I
OVxKHvhrFwzRXrXNtWm/+yeE/AaoWFDrB0u31Qk86+iUjFrvgAIJqU3FJue22S6B
x+VwSDtyAVcgazMi8L1+jHLkDFJrdQ36D1llnB/Co1ZXbrxcUZGiZE99gJGtJx7Q
IS9MHjZoQijH1ZemOD6Gr02kwBmSpDQgsXDocePU0hKgm+MyJPY1jJ2XxTPou149
XpVptL/dTolBUuFbQR9IQU96ZN+sUdmV1wSImM3mrbRnGdSlW9NyOeafPcdFVQrW
j2q3c4hphsH+V6EdU7K/JJrR+XtluxQjyxGpowOUDlutljU9ZZl8RR2P7Qt/vLBL
FeM9pc1jAq7VeAUqGZDwyV17bUqjKhaDJxayx6e8udUlcgShHONursoduljHZx7+
HoJFdvtlqhpgYi2LIDxkXK2hyOg8IrD9ILESnAR1Rv891L5k/G6UaCnKmSweAv5j
Jpbhsvt7C15HlOQyMv3oNPVbfnO96zx9IEfcZ2/0UOeQvS9McWwyy+sVgMfJUSVb
+MQdFYhP86yQRvXPnZ0b6sL3mD1e/L+7YVXTIL6g5MWMmT7eBLkslfzLYlYqWjny
w9X30JsADz35WcnmL1R4s5cpWQDHOGiEulZoOnyVsMGybkdN/tmJR4zkHF0+JTBi
Ra4VQ0imjFgi84H6qdyMGX44j7vkMP3JPsJ694cVqdpsHHrAsINbNf4Xu4gRNXyy
Jtm6k+BRCkEo4p8SIwSeFjaXGGaJX0hW6S9Hoy9UCV1uYyjRFV9C2WOCUQnTwnS5
xoTeODSSuDyYdGovd07jkCvyQGN9fBA/9Xp8S5sz9BMv+HwyM4ZTcRUoxrR1E2V8
ZX25XmxXmuDNGG2LtMqedS+nZGRofTIECFCBNGMhStkshaweMog9oEKst4RtkXpC
vi4BQyjd0Cn2k2B+zBuKatEeS9DyNG1Vm9gCiWEU492z1j+oKqFv3yWfJ8H6k6Qv
xJ69KDJhJFAh90i5h3LqtFnGW2+AQ6IP00zOidpGdTH0zUSqpfdfc962jINtWZTV
o5pJMFwhhqcEz5jjHPZGuXHjNrk4CT7UrWnB2j0Div/rkFK0+q1bgzQS8yGMBNKg
dsjnXTPSI3FvHfg4C2Q+IHfV+ySnm+Ft+qwZISlCmwqrtdKxjTBorzTyVquQUmZh
8bBq0vCtQ9nGWVwxp7VCm7EFtIbvmuPBTclNdVMDfaVtUOJTaYxUqoA/7oaAoZwU
nVJSISNfX0/nnEbtC8bzoZO+bMUoQl+GAGcpziTAvzIXTZFLJ6M/NpsDoixffnX6
pbjwIpiPoJEUEuOWAPl636QJS1EVcch0H0L+UYmBSbp2nTBX1+5f5smdaA9x0cxc
4K9qFlOZ36IUEeF87GFJKe+JPFLt5Pv1lneJ5gO4rrpW8EqVPa0SjBxMNcbrOlp0
uQ+ROSPOkSrAMRSLyb5SEYxcrl2e6IsNNTc3MYSmC1TOCEdhfdxwAlRSG1y97xa3
8dZG37/xzcEIL8lgM/eKFC4NoNKeVAuG8OAgUC0h05WArYa2xIIsHMsnXwxI+trq
HQQcxCrCIhQ6zZfeLozsVFfjJP7LNeizZ9ivRWJaHB+K17iDCiV8x/RSNJuQh7ER
xEoQZ7nQh3SgPUpKEtvATgF0kPxcQXMAIUDLkZ9huKOlvHpLw16Z84YI9tvZgeqi
5y16+9hflfaJosasikNNobZMEv6fMWEs2AvkhpYk2QcE/JCj3LR52E8v7wAbPpOE
pH9NxBNkG+k/wfe9yVOth4qo6Sa+SRXIb6PyvyaNeeHKIdjljJv41w4en3Mlhs/S
fpejJ68LSYnXOGUzW9V2wqORL37gwAYzZ/2pVRJF98Rc4Et0O3M54rV5uQezhvEu
sRmJNOf5ciCg+jkWw9WvCgFtMMPv2JfVjvUIE2xYKgVjkCcYsHN9NIejhu8KF0Eg
RevuRv4joTr5cDMk3oE47La+CKA1dcV0iyyJva0L5df+t2bPJebPeJ0C2RSi2GOZ
6s5G6m/koW80x5b8gW6SQj4DCFO+ZCO2Od1XbYwDDqc8rbxQYmjDKwZ7zEINekR/
N/2jbNerkCx4JGFXGqVBarHSX1+sL0IryyAqIJcqav8EH8AZG+rCcsqVU0jYKb0j
sBATWGZpOvAMjzbVVSQIP66e0ue2IavdsD/sEgx0+OGJG3k6ZPh6SWhTrg1qYgeh
yh1EPyv0VfhZzhmDU5zf9qd2RxXBnZzYyWZwk/xVu5KVZCxi7FHPXRH95FZtEzHC
v5IexN4sqbxi+Sn8KMblaHK5543CzuleLG3xXfrscMKyhO7Na22Sln1TVKS5mmdE
dNAmyXL73TwFFL2u3g7uOQEEDINbD6K7yFyM4UtnCmx0Anz+YvlaionVKBdl9Rjb
2luYZcwBFzk3MGFIlPmws4omSKPHwk57M76Tk05dpjuueZbyQhYzBJZqr3/w7uee
Kqw4IF7XGGoWbBqUjq1r+riRavbwzdRGsXKO+5Hm1muJ0OazRz78rKxykT2ipGAS
YAn7AO6cG50nblmIL6vzX00kifFKynWskElma7XxTXygW+XSbdM12ml6l+lZfw2S
0Km7Ri2bScIHkpHp8J1znc0/XHd1JAgA3oDQUsAXlNtE5FMdPpG20HY3whHyYnXk
81qSjoTSyPq6DLR15FvRBKe84HtwPPWzURFcp51H647GMYNs97Txoj/1dNEkD/+j
WbpfLIJY169JLppSJvqSyHIi9z+2WUDf/3z7FjLLdbrxjkHrtrB1EAXkSkLpS1Y3
I/Ax5BoUk//Os57nuN7jPdAC133WyHU7XwlgHJLL+/X4Y63o3tA2FBrUQ5OfK32C
c5Aci18bpgVGwucm5flBvy5+x10E5aJ4aR55sJHzLt9VQPC/dR+o8luWvEzvEkNO
j0UH3RXAHCy68DHi5qlPlsDp2g3x63xU3i7z3jGKP/QeiGd4mpXfPOzaHwPiQGF+
TBTDGYa01MbkOJB1/4k00uOxgOpYEimz+exlQ258oN1We6mUwJlv4hqYPI+t1feY
OAsj//sq11X7RtzwRFPKpSJquPWMeZorwQKxjnPkJv87o8Xs1AJaSIwfdDhoqHw1
wvrDf0dJFix9BXKcwomlfZmRr3VkJZSjiJ+I5jGl/pZ4WT08FFnk93wFK/xDoOcV
ZF1eRW0gSgP/NSPlVbfR2s6p6sPKgFlz+pX7kpP+vQh4LcK1QMrif/L6IlDHVvFq
4B5pRk9JNaoErjDBwuLGiHYefrpORcIoScQqbzybhZZF45lqu40814MqKA6OHSAL
G0m4v7muiBqMbMI+LR8QzjhROPKgcj82ZsFtxHnvGAJJKNjEXTgY+2bHaIwMNcxq
r28FTcjm0HTRtZthNYg03OAf02Yp3r1xjcNCk5GxDgpYuVUd6HmHmHoSDA9aOwuD
Y79RRP5hKI8Xf7WEgogNokHfNk5edVtqTc7NFQcWsjDH3g6V1AFp5j5MLH2l5VYP
4tBqWknMjrgamdIOGkoiRj99l+OgCt3jti2jswpUP2c8SVMjfhi7KVd61hT3MswV
qUeIxAjWm3lSoBSVc+yzoh++qgZa9YQ3LalvNV1s+0YDYRlK/H9y26Qf41+Dtmm/
fv1FYXZ20vpyhtSBAdp/8e1yp1kLi2hJQ+j/ixLpRdhRtEkMtXX2XXfbhQlbIqjF
3CA70G4QDQIEFt337KLhRjmey9dOb8IolIW4uciwyjqdOAz5/5nEj2IgeIA9XiFw
fNsm/9UoSF/3F2XPKDOAWtQdcN5e2IhCeuBo/Q22fCvdOXeAm4BYSqOiFtyrZr4t
qy5EuOmZ8u+KsEdvPdMhedzACwoGRnhoBISZralWBi8h/GVv8ksx+21WuQbkJfnB
0ji0487ne01wXJL4m6xkmhSGko+JiowC6EHPKorfEJaeRjDhGl9qzKNR+H6xZq5K
hGOuIJ85oB1fBpJ3zTBmFV7FNYNo8IIBlEY8wA2d9x7Aqmw9ER1gN5MsTyinG3lV
utN4V7ptiED+7HiTU2IET1gmWDZzgGBjJj2959lGk23Njo1dPa64O3Cj5FbjceeE
gdnorHUq2bdYP9XLswbMiNVNcVXchEevX8Zf8SWehUNJ3u4ES65IuUxgJIhH7946
OfwW8Rp90j77fykwvEdny2dA+fKZsiR6iDmFAzznoXktQjid1LahXUMzmnXYngOS
7zxDK7I09efrMXoZco+outQ2GT8iXxUyRzPAeXp6GGjJ1EOtFn1XJedYaKAw1d1E
VFux2DGC91bQA74AKkek65mzbMNDtTk1lsAa9Ju37meRaIl97cjHPhEEnET/RrUi
Y+akyTxbUtW/W+ilNSSZueUU2ZU9pKwuAdr6HNs/Yk/sBnQudE3j8ybJFwqGehhi
k2RIIAKs+1obAJBSBecTh/bysTvpfM/vpHG4T1V/haA1Welo4C7YNBpvU2ihG9q+
KWaiviUV4XhKU0vYuaqfvVf7A9qQc+ARU4MKO4zdRTIXVerIhwA+0ksQLjlZQNMH
FXwtXMMcMN/rpFzv6hJbxR+QEa2GWNReUcxs3TWlJQ2jAaKvL4vv9ZnDfsXp9ul1
JqqeAKQKbV/gDLbgFuw8sOq+eW5CI41ubQ25AvH8ujKodFzv/uYzWdsdfVCQKi6O
kiUPrxan6Sly1dEvfmTpDEJMj/AmcGnEiCLVg2xhi/d0aqBPzk70JsYTMdGiE5ZK
SAjdgoMyiNXLxFaNLl6sEYgv8d9gtJW2xertNh5DXUz2Zc4UbMN7PRSem1nDYmne
vwSYhbS2XZSyIA9ZFhAS/Dk/e/ZoWm73Rh0PjaikM2zQ3wxoyCcZcnjl6ONDTyfg
mgWQ4eCFDLKaG07jfLzTQ0u0pYGIo95aXU4sNUN5CFRFyKuzjT1nx46r7d2cXLoz
/0deM/jW3kuKG9/Ks9XVvZNO0AZnEC1dqpXHlg1XCXoTIK+Xdv7tl9zCKNuCjVxK
RCZsOhAs2pCpR1vcaPU0O8lIcutT/QfXL+/vl1d6fyuOKT3GmFZxK0eZrfPE6s97
ckxf/0W3O6mRGGYYA4oJEQjEeE9BKJpScOqUpMs5KSvhZA0VelV7DGBalxkTO8XT
fktNb6m85vw1doqPELBl2nE+XUiQnr7sQ7/gvIAD3KIJwWy0/8i44tclvYCwVDja
hzVDRmXgGZeA2JxqSTa+ghga/Kn2FN2FIRDf3mKsZtTJF8IdBruoFrbz5BrftsIH
TEaKy77qh0Pgr1m3XoTlzKziN0krb3lIG0N7x/J4ehEcTPmxIl8fRbS6dJzaQhuw
QucfzwduAKIsdp75yOlDjKKvhpCknX1kICQi4i3HN2MECJMuUIBVnw5wuVrmAzUO
SkkwwQcZ47iZiC+rIthwh6oP7ZTQVqy2atXKMtZ49WPhVvqNqudADp6YzjG3NmNu
UBFLl26PD//05HNdNg8d52HiQHkQaNNcTT7aduniZwqD7URFKe1M2LbP5H3HQC5A
vA6ucmAMk5AWU8bEo0poxyv4rIbs9eR9ZEE9itUNmsF/zjS9jpsxEtF1Xq1T99wu
Zo+h8Yn4mdDRhe3vjj0WBv89/RPrkXzlzymD+uZD9f/M0RhEIM1FjMN+I/O8m/1K
5/8NZuYghXxmgHy/qrb83/x4lPUmn2jIoua/XUWtnIbN5FxPE40IFRHGhiLNwo74
GpiZeGOVqn7TABOVEteuRcCazrGx6s0THsl+vnHS/O7KucLi0jzhmb6XhzzeruZh
En2vq/ZpajtkMjVFZ7/6Lurq8DgoxJDasRKMkcyBoRdL/vZPWoessZUbug1enGwJ
OwAttoVY/qLvgqc18JMyOTAmMju4oWzNbxvYHecSBMozpeMsjk9vidJB6IUES8AA
Zw/67Exmn/QXrapJjzhFlvGjSFRFtQqemPYLvtYDsYU0xPzDrVv9G/Rb2puEsq0f
D456nuqSdrCvbWP9YilZdYyk7TYYTZSeNKH/I8SUsUDC1qGO+APgyASrBzNpspk9
wMCVnNhmZ9ei1SX1n13u6WoHiqpnxkftDT83ULKZQsr1pViIWCcgeGc1CtE3IojD
PSJLY6cBve5fhEVJN+ibBy77qKiMeg+W8xfexTeOvmo01oTtnbJjA5e6/XBBUy+C
fZnAGv+XvwjisCNa5G9hJ4fvF/z5nendDM7kIuSrNFb6lu0YJt6C79aHzMljnaNk
SyzbKZ+oRmuQCsnbyau+VbCD6VNMoOatxcSKakEp3JgV6rWz7NLGBr94ibOpm15Z
dIlRzuEi8lDR4GEUXz9SxNjmxRyA3MJ7Y7f2JVkV0HE/+OkzC3H4sp1b3LeF/qap
ZE2/fP3dHM7BhqWXraDCigzchDuAlEcX2zOS9ysV5QcZLU0lM7zEYkHFpEFndbCd
zcEXSIx0nxLmGnz5zJjY+/frswoXUgvQh3Nh9DwfTKp3gSSt3/fbgwIgy8BmxT8M
nsJObyD+Jud763XRlW50vA62eRwiH/EuLUqSE3dg7xNttOZ4WXyjG6x4T7Jy00LZ
IP67JxtiWEXss8JVAxoUolBkjMe+BhlpiPq/7vZJBHFzidNePrEAfjpnCmY3pFFq
A0+lRz8sX+36DdyVIkh431O3Z/pI6wrZjaQOPaI70Prr8WW2hXvyHFmHrkQgyVZW
urTBmWasofgOKeZ/Jueh7GFZrKNjQ1uHhU4naMYta+BozcOfrsWPpZNJwS+MBV6R
n/094DA4JJ4JDLxRBTJNmn0S3fj+omDIFHJAp9D5aTrawxTkKnJa7BOm97SGpytQ
xXLww7guTPi25BmPdPKqA+UuXhgWZ7v4rHtuzDpxzcr/54t4rvtjER78JOsDeNq3
tUZzlmxMyJBX4G3dneQeUUaIXMJRts3iv/aenFnP4qD+qltJaHUSAM2saxG0hWv1
ynyGi/RCyIgk8NE4OposSSoqd06IKeNQX4brpXGrOxdzkbdUn1uAizQIO5/iwAXH
YZeSC8M9o3iUv5zEMr8JwklNwUsdr55gHoLZ3wwI5fkhsMifHTYhZ49pwLAF4PKg
gexcopeTSJoAo8TvTRdDePB7d9QxcUMLkArw4do8TItUGxoN7iaYDwaDXoSZFduO
5GJ7hwM+EfnkV3bQr51AC5EPrMDY7EsDliyjkYVkNhn3FTHSmgM0oORW5uzYHu1V
ly+pNTA5gDQJ0rIhSOA8dvfAXcA4DbT8ET7GMyPJHLiWpIcw3g3PXQOQ0vthw+ad
h+PsVLaNMwS1W0nfsAq08ZivJgLWA0MQ8lndsVb+90TkNESrhdb1AI3BVgdHZS4V
fmNGasNK2HV/tII7MH9glYiXSVYX0ruy7QVBR1Pm94Mi3PqjZMbYJWNGGiu7O4r2
iPNzbwT8YZV0IF8KGEJRuB01GgLsdwIRI9HGUObvkNzx2bmaJSQtYWnohj9325xv
AJ4oiuhtOGmgcRsgb8Ay2tG0QZ0eiKkkHdzCxMGrXb0SyLr6S4pqAnakv+RUdzOd
mGgzZnfw7neEiKVLkidX8n2RgJYcQmLViNqd8YACnwpEFZV8eEDRFB+Ixc3pes4f
cO1T5dnwOrQ9Q0KUROjNRNNZ/0BGzZVCCDmfopNXuOIRMLwxpVBJBRwBtkTkl6ZP
RkFcuq0oyatOGc8U5qNnHgJZdd7UXw+fMrObxKt7gQgxftv4Q4t/n+lwLj5XnLu8
iR0ZpG2GTfIMdcZwHdwXJ0S3miR8HobNbUBHkCHZQMqwZ6pl/TIE2F6GfByv59OJ
Pkj0J2gwPrPZMs8gy/G/GqfoluoneODQc1AA46DgC4PW18mDM0cfDLoLI3hMuV3U
g+q+KOakDO6vvrqWJsy638kWdckNZONgnWAD+Byj1xbhVlMA+qX1o/C7a6g3l8lw
SJ3QfTYCyll2o0oCoYvO8RXEmt2/M1WrZHVV5F/Eax9OuIp4tmtKGqSsaiLp6FPg
NIVw/yW7QhOs4/1TKdHz0MJaSvzeyxS6nVpe2t9I7o9zr26WJeIx2+0U6Fenu70t
cN4ydrE0cpHeYpkwUqPJQvq7otx9y5e9jAQHMu/7KvUCEn+P7OkZSMdA8tObrZN+
lcnnsXobi3mpos5ufopEgUiSg49g4DlRz21F16KvILbfKbd5OqW1Y2mEDxv4SjQ2
U66S7U/O3J9d3DWQtq9gRC4wG0D1jgcq9KDv6Y35O9K8mx315pkz7fgsge8jlv/r
sIPhgl+0Y4AsQiAoFOJoYobm5m6doc4LDVC7AzcG/y0A7byuFFXuBtSKOUNl+xvQ
YKVRnIs3OJbOgqzvNJE41+IJ9+XobtJZLo/Du1u27Fi1kAlvIDgZiQBuBmW9pDQg
RRClcB7FVGDtQZYU+XaX7qyEw3EY7lfqjHMH4P6rD5fOG5I5t3wnXGbYh7ojWVt2
85ThO+RvQsh0hnaWU2HnOG9TUrydDrdSAHhYg7FDkQ6nmWMcMO3RQlOWbNxsuw2I
0Gurhead4KIdGP40f9f1y48D1an3XWld49apzqQtn3JKN558v8xKDT+pY6lBLugg
KYyGhPG+T6R41whtX5JZNLtILU/lWK78lZwscWi+PCThv789vty7wYoIQecLFOIP
aHryvfHoBQNsA9AFlOY2zF7F7JbM2p7SwBuk2ZFmEcDHbJk0o40Kud+gZJU/zxHr
dciIRuqcGY0hotSeANQmBLklI/Fkxe7GSK/ieLJdC085J/VP3pgMfS1M0rQr2zLo
vcdeA6zceo2nBu+yjmW80mjlGMSqQI9eqzCqS01cT9ljXKtFRHENYpL9D4qECnwQ
VYQPF9ZzMZTOqgD0UPdWRSZjRQxD8Rvz1VyGhWQNDszCJV0v6RLhpBZSnPob5elA
MV0h6hYnwwsO0qdFJp0zvR3QFDNuuiNCAV8kSNSFZku7Zw1scl5858AxzqZFdnU/
9ersZQRkluuJSF9W8sh7f3YXbEueNiyNwGnZRXXjc3kP9uaRLo6LORAkRIgiKS5w
P6W6bTsD0u8fDDaxhsYHfhQNB0MDbarXj3kDlKHZXzepYuMLMz2Y4eK5gc5ZJiKS
+urp0Qo2s81IMiy9ra8xlxfjucQ8TAbzAWo5Z2JDV9LGPI+2wUXke/LuZcML41Ki
BkbVhWWJGxstAMVrGJKM3p7EJhRYzvWnok4R491KCOAQmVrPZRhnVR0mp9kESeAm
lMV7Ynqq9nSekHqEQ66azfr8gFNsv2k4fZnAudFUHQKglzZSvfqtEIWE/T2vfXbW
duW3rNOdsffEauAH1TqXvZh5YQ8VoDuUwOfpQosv2Z40lUk1QZQxjUE3hB8xcqci
Wd11tE4oH0EqXXjndaUUJKVbNJMYcfeOWmfDYFUhRwZfT9lJNxmx1/8Z4SkxFHeL
9frKZjMEUDq+vJW+ZdseHasVDdJD7IyNNENWlUHWky2lZwdzInfAPfWr9DUU8vzQ
fMmM8Dpoq/UZpaNA8Z/htMUN18N/38E0Yth7giFRA0buypZhPY3g/7Xp7QJGXENI
weCA6QIWa3hhKjSWMYnPdkzUFSPtwqm3agHWCOFpfHti5Gv2Rf86a4Twjdh+Z8Fn
Z0khfbcxkiAXbawy0PIp4ESK89oOff8o9swq/jUQiUhXKELWzvhlMKMiaYtUN69k
PH6T+YXjSsfE/m6dxjJUuMApeojiPJ4ib11F7phcYLtPpLEaSBOwdplq9wRYwv84
LNZgoQDZ8m2IubtblYEdpzddcz8G50R6eoOa1XhMklz/+qBtlQ9sL8PSeGyxOy8v
uyKtSS9mqhZNn3Dzi6W3uyTfclzARhmBWcJJYIlp56LmGmcnE/t9jpbhYqrjf9tX
ChiFvySSbhWAjK56/h6FGJ9ecA+mM2RCEnOxUPIcmAI9YxQt/m42aPytIko6JbFO
VgenuZkw6JXvCgIIi+3ff9rEtFAIhvtkb/oRIiBnOhv8kKBoAEMiUX4bBnhIKn32
UatHoARbSevHrrHiegKZvCZlxMjuxvYNrljwWmjnHijR+DBiJLZo6wLuurmGB5LG
+M9jGio9qztFziKnTTqwvfEqzE/o9m+g7sE0YvRTDiSWb62VpUKsp9pSFbKqh3vA
poP01ssRNe3eT1pRrxWlLCO7ZvvV/D/HjuGuVmK1FVZeJ+9ErWawOHWNaiccJvTL
siGjJruEb2afq3WoW1WvmYCDC6Yvt3zhFmzvlpPnzuxlnvL7lB3RJrQ0ON1MTfus
eZ6zyvn1T4BI5NHXUpgGD8CMLg6O0G4S61wZLexaHyrP4+mk48oJORCb5O2g97jV
j/6dVD2Meylv5PEzKF1xR4/JsD5YbWr2H4zhBAej4PYUVlvwbJPS8tSKqE6Oxss6
Nzr/snn8wIhnXW20CD1+fpupj9DOo/L6yKto9Ns88IWQ7vulb4UEkeKOBwfvSFw6
nukL8rIS9bi3GlCoTR2g8g0P9A4U7oa6yWIFPbrsuKGqeyLoqRfM88zP4kTZUF4Z
rCMte/jI9FJ0Muh/x59QuSwyyoSimHxKIuh94jUxJGC6ex+8RS2THIq1attZnw8j
zq+g0EtivjtCUaXxHllnkC09CJj1WKaU8DLWOEjeXLnOw0pRyDkINHHf87ZdrVuV
E9ZCZXUfymyvTWkt1dWYIgDf2rEbTHE8mgz0g9pzkCSD4IqaSI5Pm7OOn3o+9mvd
wvXEUav5ROHEOaiQIGzVl1GYvu3UzwOnhrvb3eDc2VrmvIcOkpM0F48g4oSmcLqo
/qPngmfH6oqr4RolTxw+r8tO1kJVkE6furzIUfai3sHwt3Tcv0TciAzDBOfHYip8
8JJNsCRJMNdp5c0ggJ+RY77HdAx3EegULGPHOu6tWTguEBE7NmRkPNXvxokxAPiP
CaFZOuSVn/mxoa16foTLkIjSTr+JIhdLmRwR2fqSbdOkVu4mgUu7djLU5OHZMPJ9
UXVEzoqjt7Wx4DgYVFFUuNdvwVCN3B2JH4w+A9oCUDIQ2uL3jcYfsDWLRrxJehl5
FTJUkiiPg6gGNHlhsP9awlA8QU8VgWF7d7Yhr/xsolzL+WhjE+lYNQp4m8w3QSgK
zWxdmmxlo5io8KUj0pCsSbHrEF3GIAzhlPwbmVbl3eQScTc2j2RoWYt7NqlnFoMk
4R7oROmboUwmubCVBUx+X9Gk9ybyALLZofhyIoqwGmU5eesYpu5cXKcDrXMEsLEi
TVtqJ79GYDH0BZwMnpbI/2x3BZMqsFECKBg7+RG8DiZAcYiLBWiTF+8JJsCAo1DZ
/EgIdPUFn1qtgGh04Bdoets/WoZcdNEg/xe+LgGmNEDEVVQugh6nNeTTYQCQIchr
J2txAI9O6yxZcCWiObnoMQN20M3DWRpUP5pIV4du48ElFMn0h6jjkUYPsrNRZNxo
KyRAn8+qGFtA9EKcbozH1H+asS5hrPhelWAeM7fiPpbRjb6/z8wsmNrNJiePn5WP
BnTNXMv+vG759SI4jAuYnAOpVbpg8asVpsRm3EgjsbKlR7v4BlEu8lTJfkujQrEu
D7Ver7mRJxClY9M1qtrxBWW+Rs2jGMBGPLS09WwB/06QMNboDOF6NsF2aKM8rxhS
UWeDRX+5URUW7m2jMGpkNjkWOqlV0gvSEq/jKUYrU3CGcQ+FX50R6dJEJJMhzpV9
pCEoT8YoIagGGexwhZUB1zShifEIhP3Dv3VStqPqXzlAw2KHzfr8GrV32329x6FZ
WhbjRzJN85p9z0KgBbzFYRdce9R5Or8T3FrhdEcdQ5Zzzr0IjeLJxS341J1WIb0v
ncS4RDl9YBnFiWJGg38nUBQZXjrvY5icVf6NJtwu6WC9xsa9C+0t0mjLm71JyNq7
cGJSTw5pkmorRAce9Wg1h2QRdbaNHrYToyv2BTs26+cpUQEEdPiknBwfPxMcu75v
KShSh36z3WkDTxPXKfAvpogC3jghZAH3kwqs/OOwFohXLyuCH7esQbtIvwsVYUxv
AkBPTkezulEOm85KrK3/8DDytvcdaZFmE5pmqtKzXdzMzVhJ2p9p3kZtqTazQyI2
nlfsEiaYG3qruZM3NltqeTdaUq4vWvwqqhjbjwVy8exlobQ+2Kyp9Q8jUNV34Ier
pfGYcIQqpkYJTTzVpbKgbbHe2eCSch1ZldY2jBHroa4q9+BueCuOAWLcS3uar22I
/43XhChIjpuvkiMezxlZ16dAiMz7q3Vfuzi5obLTJ5W8BdwFbgsNzlIQlgOn670A
aTHGZpdsMf8O9nV7oL15x45i34PDmOv0UAuPYzK3aiWzzCIay/SAL5tiyBosv2c1
OckGsbSm/ei00q40LJR9raqFN8fWQFWwyA79K7z7poa0oFE+/XK4PbOcGBihze64
sMkEXpA278+YFKwgxiowrGsRT7SPyo2wL2vkThqdWfwLonPO8Ol0K9eaJlw5YGJT
C9b4LKTT3Z27loaMrYMphdiml2BelnoRLfCClsI9c+fTk6lxKTLQHA7SnZFCp4TG
lrPdtX0UFls1CUTeqXMOFGz7ZVBAiYeot1Rz100g4fXGXXg/q4Zj5zN8Lp2kKeVw
vsOVg5Y+ecXr9uiSw8MPshM/IbMIUqRBMezGOXxSoml9s4AV7ISQvxyHbfWEfWI1
PeJBIV1sIIR5UHwxCDQBXQ0ueXJQXAVrjDL4txfK/fsa7tkScisoE84lCqdrGOsd
+Y3ezi7MtIYUdN3mVBpZQthm7QLemqUSIQvBOwQPvO1wGL2Ni+I2C3/yNWbfWXoE
+doWZ+nJEa/kog81P1MJVcHYx1M5GEmzX+VGL0KsvrK6RhSNbJsBpzY5lr0I5QVx
XAv2tr87qrZHuVQkkMGu3GW3/Mcqzz1H+qsWRfksbfTRtDU5ENOT1L45idSJRr8I
TebW/7s//KPqGkOShc8wrNWA9M20ULbg7eS2v/HVFNy+7l9kZfUC4zL5xQ13DV01
fbRQxVYiEI8avynKRBirJCOsXuScJbI2Nz6YITYvU2MCFleQoNTMLXUzmezUyKVV
/C0S39EH5nALhlxEhhpFuMGIlpfnil2D6UIIFk//LRLUkQIK//7UcyEp8xhJE5yp
t3toBo/kZuKQnjj46vciU2DDEx0LiqU+G/Dl1C2T3gxTQ0iiWu33HMOe3ml7d6v9
7IGzWQ7ohQkejEgdnWhEO8jfO3xuDbCTPn90oJY0amGFqyn/TlGbs4BcaJ8UvQnP
+dMwvRKB5HsIJjR8IySYfJpqO1nVUDt9zA0QRB8ufH5IjRnj5dJpv3UDwuXT/RvC
B3K7t0rkOxVf/gVVxoP7BONH8zV0ON+oODS4bRb3wQofPy0+u7ZM/HpKwb2oDjgc
kua3FV/iqdb2T1Okdtur0KL7VnCMlKJAUC5co6Pd1OLWhfnt5SWTG5tOA1ZLwxCR
oZvFR9C472O83PRrgSquKATEqn3gPyJai1JM3VRIEGjD+UzKa30dciGyzMDbar+l
r2QcjXiGHl1wbJBq2KrFc+B/VQNk3E+D0H3vPeveyH+QJEexLnHO7aEpCBhN1VVX
SCyq89eZOyaDzkxM8P9f960gSLV2N92z5KUtPaMo1lywbbzCMIDa6NAsTZIB9O9U
V7PzVdUR548UEWFDOo8dBe+RngTxyrOrBCaAM5ejKF57VF7VXJdku088wv7b/p0s
HSAk7yME4rCX3HzZ+E4ImUcN7WeK0U3uxglT8jV0wFRPLzrQZOrIREql+0B5P56p
JtFCeEc7scsSzDa4gCSQBIp4SDwUa89h6hBo506xeEvzf6F0s1chpRy/osvMSWeM
baO1mu9sjv+aib3pbLk2Y2AW64zbPImmunsECIajWvvlDebKUqSC4VaMIpxgDJtL
Nov9NTlZx4gt4s37yh1Au3IOHuASoDsisqwJQ6DOT0duKG5xlxWY4rCty0mDQr4+
zFnjwXTBDJf6ULDT0sGSWSFtNmGTgpbA2Y4RBj1j2PIYlgAl8y+AH3uAvGTJRJzP
03XlByQF9O30bGUHM97kySDNKQ/YXCH3SZR+m3NyJeDDNL5H0jFJuny/K+ehbu5L
5fXROw+Am7ajj5iea3zjFXzUW9ZyKKifFJoGKTBlc1kEc2Uai7btw9FYS6mHf2h6
J5EoW1jZ85eIgD/dOOnXOo8q1eNcVIElHiWuKE5ePF4pkKtVy8loCG8i/pWMl2+X
XD6ULh0aXh8Cx/oTxvGTEeD5Z4mBkDoCuhEmvbdIpzbIvNFn6rKysrCkay2SihMV
DwAE+UxLwD7SLrSvhuVMl9mbv1lleasCjziqbW7ybQ5TghFi27CHNFd5Bce4vI/M
zpAxwbK3mU12r1Qpuj2PFCydX99AkmrmcWbVZZ+b8Ep5V70lgm2SBDEKLuowzSNL
QsQM1z6uDEOIiB0aTo5LT/QoXElFLagw2DFzOQJJOVwoQEjL3iaOzJD+Ljc8SXTU
ZGHingTNlKMb/ljl8QQxK/SG4e5tHkU+TT5qsHv07tzXtelMZLLZKTs+OIkBXBy7
gYipOyA0loq28im5DaF0x2EyLWlZOkwiC4riDVzRDVBwFWrQJQXoYCCO1CVpfd7W
8bxdecfpIs0Ad54/bJI5oAB29R6gQDoM6kO3mSM25dfiz9aTAkn1obi6HoZsfTu9
gAnuV72k5OtHipDuNmAXjxb5XdJkGNTx1DQgCKCF56QIT8EIz5gJQS1GilHBPUKo
ux7o0fsW3U1vqY8uqHFOxIPtFve3t9tnjV80sxeuqc5DM7WEs7dzGXToHh+Kd5nI
igiGwZsHPUF6twhXBfMKrdMedai1ueVXKyBg3xGxM3zIkkU3Pg24jv7JQ8jKAXAS
LHeIsevfFf0+XXdAE9ilELiGjv1Y6CgDDOQmLvRGvsXCADal6OoLkvYIGdlYz0OV
5xtPgX3TpHVnCL2hpc/1i7mr5QLYkELADqxSEdDfyN1XC4g9PNYgniVxbicrx17E
J09HYnJbrrtZ38A9wLl87k3TTHxviLe9aaQtEFtbb66WRxx3suNoogLqiujLrZZq
rZEAPI3eosTFmNksJNaYgf9rsv2HS/dqjvx4tlxU3Ooae5TOLuuCMk0HdnLXbNV5
H68ufLbzDWaXnRLF3RFQI1IupBR0/jk1gvHlWQ9kG1qP4WP5fhtiBKdpphZJS4DT
fZMd3vKd7XJsctEycxEnCYhIeeg7wx9SVxs8bzBwf9sHzj/puhLyDSXVWQCWwyyS
eRIU0s4xBJqmvESGo0peENBF0IFn49LLrfI6fbewDYvkj89mNCcXHBqmosr/wJGz
KYeWVraC2MyfFx04a/gRkeiA2C/8NHUf/1oe8EnswYjyO+hGBqDV4D7/bb2c5p5v
t5/ZOEMrmqnuxSC5qkUjDoeb4h3rMXe7FmMAaaSVoSXbXJwbznasj0TEB3M1Pm/Q
S7ipilne2bDcgfYa89MilL3uvCAeZ6hjaZxHRuXJO66r80hbgFsynzsQO+Of8t4d
k84CEbBUwz2GqRKGDWyOsnpuQuaCDTNda7ADmkvvUY2VkuoAM5GuUS0j2YZx+9rp
sE9YHXUHxSnxHZLcNIceKasBiiAW0cwrQ65Yq8VZ6gEq39hbHGbIIpHsPse6UVRk
U5gBF8DxuYu6uR+6zQ5y4vmDXLPaYPnAOMme2VkXGzKpdq4qVKSfmZHUMNsrZixT
gNA3htrHj3OfyiqYTu8qYWKfnpZlmwWzam49+AN9v+e/HqlORsr4a9FA01DZJlHX
xznZq8JY1PM250/POl6xuCXOdFkirBp2/Se5X6/QGviHVDE5OeM4kgJ/9X6JzlSH
zz5dWBRiEdY9zpWKxPyjKb39byzPVlXFusfEzoEAPdoLrBfJTlxao9d6ye+lqqnp
uwuKCsKqFY3g49cI3dTIWC5m3IDxJxipR1dVL5meULorc89MdjM1UTK1uIn8SRod
2bRcCmBHUUMULUml1H2T8Om6t5ff8Kzs4SZ3TSXtj4dNBMicmRfwQOOtWXBhRAxG
cQ64MWZ5a5WuadLfm304Ckf+KxK0mk61aK1Ji9fKl9eGVSkHjoliUCxzZdtDE7HM
ANmuLwnhB4bYviMLu2k9BRUOYoYmAP3aeQ616BKuOI0r/m4bExA16pKAO0FOh5Jc
KHheOhiIdLWPapok8nAs36360poqkNbPEZxCQQ5Adi7O8qW/jVB3W3xj0RK6xMlH
FovBMmD1j8If9LDO4tvT8qIV77BSy54vwjqeSgspq0XXm5oUX3ItS1Sng0TrCni5
fR3+Z0EcvDxx94a8TOPKhN1f2pRmz/PRoCr5txXj5Mlgj4NQ6Caa3sd/DZ4pjXOq
uIQgIm7BjpKRGGD6D+zYYaFPEG6VGk8zwL8lX2Q/GQfXnrT9PdytwDY2L4RwFmjN
xiF1GruKlCP1z3OI+foVBWW34Eqt156ctsU5/Ijj6QHquDecqIxU6h91bLbNUeQK
36LVJAMoZHNp4FZmwkBS923Gq4hpiANzhKYvyh4yv+MxRYT442FxIlZmiB0+w9A0
DQgPAG7PXQq39/M8YrEAneyjyBTBF5w4t6tAHIH6J/sAY9pjGSOVrX+L57XNA3R/
RrsCB7tSAstt6bN+Sn/hjYkMpXJN8QmeytWD3iJmOYNI7nrFIyY4lSDJyS+r2wTd
os1woRudfVJwKapa/UuqJJpYLP8c6Ed1EhRcRBajBHo3q2mQn5hNQoPIs23G95Vc
ImRj+OdLyzFeGYC6tOS4+WmWEWsipPkJlTqCkm1ZWQ8s1QHaZat9xqXZKi9TNpLG
gPZyuEI5G2G1fzgNW9+qoAh0bffik8GvTVukqGKm8KVpdnjKlFjGto542UtGaFoy
/SavxBAzqgDPjZZfLuWEZgx3TLU8b201xgcETN1N/jqLEpYA+8l2PEptPL3J4nbQ
XgLL6GljJJ7jmwKxDGDMBM2qnSBPlKHuAN7nEeP3Nk0SmqECSBhateIzxNKAvziK
a5pdztWgQCKfY8mRBuz3DkcMrqUMXBZahXOG0JtGNt/UlxMoDDLOKQKeglGOfhLo
z0XeLuPZ4KsIFRAuWQhSjvQfd9FJcMYrCyPHtvWJjCsNZXTLLnuksa5s4RAaSP6o
Eia4QU4sSANduHWQazfsvgfn00YXJUfyKOuQOmhmMCvQDMjmh4Q4LfFtimTHfhQA
cqy/aox+IYlXGift9nnxLSOmBjAgEZ5XmqVRBBWVoq8Y9eggOHude764UJQLYqRN
3jZU/ub7qFOcYIGKLHNbIlAQjGCQD1OxGyHj8teNl9rxi6gw/aSbSpIbOci0eX3i
T+8OenaT36jJxFeX/Q/IyK6x0HpXmspZOPorhOyPut7kGhtqfBXEqfExhPyzBqVM
GjMnSmsh3ukB3woGxLImfqAdS4A7qdJ8bi4sBBoSinAJwvJoa2sWSNp5mza5+DiP
vxGFjAt4KELY0nr2tVNk342Wr/i7FvmZn09dcASuUG7AgkmF73XkIGHmfkw7G6Nw
/R8BjWyBb6IBCE0Q62uqVPXsdr8uadvrGtc0Uvr+n7/p4pAOsyps0feWVfNvow+w
UQRIBBIAmbrzzzI52cBn+9U9DGDuzlkjLKpIjBx9vgTz9W59DAtkMZpee693XqDF
ZU929kxem0BloCwBp+lJbUcWx2956I9x3Tkn3tl5Mb1p/Geaa5FSrwrfCxRK28sl
eGR3nAe15/j9oVJ4u6MyH/TX/kuh3n8y4EHNXsV6ppQ9iM1mwWWxB7JrjcSqqU3E
3jrtX7oef7N0w/8wP/eUfCOALtXtwy/38TMqGfhsfOUPbAhgPzIqOro4ZyRh3u0I
4C46tonvKP8gnyblo0aCm6ofgrDUTofZCzHQExg0hD3t5hrSDZQRJWDOr1UUE568
DmswV0w9xi1pvBwTIWZAvlKuLxkq2bSbrf9eB4BO6nDp6vSfs12nnAfhw0+dbOD1
4KFH0Is8sWUpXsUmxEkJemS3ls7Kxtx9hT8uqBzTHiJRdWZc59sy7C4sHCQ59Hfj
yLgLgv+S0teOAYxrUFVq/8qOdFNStJiM8PgFxVsVmZMd7HStpPcW7yky6GfdT84y
Yw9hl3XtCIzhqKrysNZfsZ2pAL8SHaClBV0mT8XcZufTWZJifG3dbggWQwkvAQKM
bcq/9Ian45m/l6MyNPErUN0J8I3/bl1CPf/FHTo8qtN0Eja90D0fE0utLcmC2qNP
mKwsOI8Gpi7t4vVq3OIumUQaHBdaogAI5fI2r7ZpD++PuAeDPHQIuIq+OjL6l7tz
nVafBFHFV3nWUFts3WN83LPSgOKceeLU6sC3F6ylJw2FRJNt49aPNuIXPV1acHCh
tdviJbSYl+dz0Wg2xoAUlUB3TtOY/J2bhsjPFmFK+V1aMy1aklR4JYxEk7KyHqtT
s8yOrGMIuT2+xOkwaNZ4FiU5lAQpsi2ESUvFC5d03gTiDXL1H0D0hteRcoEa5Lh5
hlT1zHYW0/rwDYbTItmSp/5oYP+vGkqTMVu5IqsVCDJMOVT9LbSQkgGfFpYKVJNa
c4yYPnssFw4vlYmIjc0D5aHFJ3zHCOofR6UqLIqLBqvOC1+SYBsBCy27IjKuhMmH
MXuxOa85cY6AgdV1x24YMY+oxY4biH9fM7RRa242x8BTFtBehGxhZoNpxAN+9ggj
i+H6+kO2LUYdzHVa3lrLXA7RsYq6yJykJj6bcNFskbJzWyZ3i/BtaDEfp9jAncPP
GTPPmxjhffb5dfmfNjgMwncv9i3UFi8CW32SPrfgeJRkfYIq0hRY3zPL9jLQ7u0P
Kn5M6CJ8zBp6iNgH4yBVDwnRxqVpDA2/Pjijm0nKNKNIKlVTIUejR7FS+/RqRL2h
qXI4zlFpV0asP27XThUnz7oJkIiSReNCyU3fMZPGgsJcZWyi+aa8Rki+Qh4yJ4wC
y49+dLPC/1nUoGpepLvUYkTuBPHfQPMJ6LvyjzsbTIuf+dELbDqZAok5SF0I5guA
+/45FL7DxLucoP6w81kcx+xuXO9CbvJVTayQYYbKAvQNyYbBFBZd+cni495YErWq
C3QNjR15tmqN+EQGCHL8i6a9/IeXeKmkRNuLeACCAmXySsNNiq1hZtROD+cMWWYo
rdig/sOuXuYr/ihhnwmNJl4i4ndpx2fc19V1I+Ghy9XQahw8zdJmxNvjM60PVmId
LhEgXIctT82BARP8lPlgV+2DTYPgteqbLEfWMEJ4kg0AoOCWqTmG75JfTkpclDhB
zGuqb3PlueLIlZdvUk14J7AELSoccpB+LLAnMLeQFxLGKZZEmsn3gWwGf/agSvcd
AUji6zARo1NXrnWQ9IxbT+RvkCEagAbfJQSiy6WVr1tJjDwQvYuyNtvpu1jMq/kY
PS4SHzm7OzZ50SppPSmCeKUQK8DVsIAMPi3EYOja+jR1B6t2r/aTYuIIzaDGi/i0
GTv2IOVk4OZ2uZAh4O3/aCGgTM6uNOqfmZ9QsNIQNHYmLJXnfLWP4Ej1E+Th+Oz4
jOaurjioEwSUhq6zegIcQNb4z2wYL2m2cefnmypAfndAnh7NKz+9KZfa3FKVriCQ
/Ga3A+cnf+GbShtyPeFsDuejh7E8ep5rzYc4CMc5jeMxws+Ka0ZESOFPf5U8NkIY
PspXtFnGDhuZFOnpobX8p6RAZTHQqe4Y9Gm89M2S5rdM4syrtzl75sDvvREpfsmA
FcFz2+NR1g3/m/A8+aRNFuJKKA0aKW9AVmLPux2H8yrs+gki7QHiD05NBDqq2uQy
SzMG05nfCP2h06fVcrMXolUdPHs9FANS7hJyfrGzJuHssL3HO6vhC4gW3gJii/Ru
J+Pv/YvdOhv75YKitVxQyhStsGnKp4jubw8P7b4EBF+4KSCeFmEyUbwDGv1cZEWS
rTsqnuli6vr9SPQEKU1JA9q1wGjek8p/3/97mSmRIpjKYn6ZCeZ5mzvbRoijahb3
RDdgjJQELUeFU9JKfirQM6SOVgSG5UpYis3S6GdOGtcgkpMLYXdA/kp5HMiFn69b
hjJ4mZm/+nKn34+Wxunm3ssujyHwCSUSDt8bGFlvbmBQCVE5syIKgKJG9v3YaWnP
ben0RJOJpToJAh2cRtNLp8lQSGsq8fskD+gI4pHK5RwMU3ev45SFGFfEfIGpeecV
/KgLJS378t4ZiWzTIF06Qw0Rqy7tPD9hcpk3MOwx6Ak6wWBiNMenyPVKZTGFRYmW
VpDMOfvN1ChTW7gyltHfYBXW14PtaEPAa5U5KZyfXvD29fDuKc17TwWS9rLy2nWO
m22/KeZDeN4AO0WXT9Fn9PUXbOypNwm3Pa6lcZZb7/eRVzIQjF2D06VOX4v4YnfX
eQQXQ86kyCdeshU8ilm4t/GlOFOHufzKv9443uGw3inkghBXZTL+qyrVXFpBxFkp
M/TYDQi+cwBWss7Y1Rmq8tvG3Ac3kbdyJlU9jH5nKP8faja72hrbiEVXzsBbgYIN
AWsij1SNC43df4dxCbTDinNWDAibCksHZ0tJjt00yFiYiTCiO9yU6uSAqPRQS5RZ
aNZuvYU4lX45h1HXUV0SlfaiRFkgJEBuGJ6h9LvJlM/uLZLNpor5YriZJZRcrGhh
06n4aUNMBgo3OwFIeVUa0e8x/siBKwIB0Vmsig1JR3CoL2vY1DZ+sWQMRL3ml1No
t6IBmcOUpT75JCh2A70joPtW7KRzDK1Vfq3Fm/GvntM+cK7kJMvkgBbplKPzO4eG
zaIKnUPXPcGBgWE/tifLn/rf0jV22wLG66mvXes2BpiuQtQ8ooMbLtVwPYhni4PX
Dasw4vBlFTrR0BDHTwQInZ67Z+2fyE8H2zSQpljosOTNqAY505pbAS/5U//iBCgu
knJuB7P9HlpncjXBGgltmP0iQepDzezO34YvwOaaKvsNG8yp7avyn7jNk4rd60ZY
UcJpfXMO9UxzPPxRqH/zP3Zrcn+gqkq7vORXIMKZBk7CjLr5mrEyMQ837UzAC3j3
IiNWMYfOL61hWUW+BhvkNH/iyo45GfGkCzwsUgOjWx4TnEhy2tFDC8S2BQnm2kfb
8flsXMsN/oQv5Am2G/sabZ0hyXXkGp3SY8TqjlxV5GISDz7+gc6GZt/sV2+caUEw
sdQCaFRHFnRQcDj7YCT3ZGR4E3PUYvYsM8r8UkEk8IsJazwEoN9YHngoS8PW+mwP
9ayjA7I4kauinaRYGUfS4wiuiqNo7AsopuB+MTtKv26JpgFEnoXLFUf3rQMCTF7k
Th56z+6uHzZxMDIXdGt+hZnD5QK96LARBqcqXoE+HBBWNo+x79oAbk7/HbA2y57+
lWBK0drd8bj5DznHm50qbzi2+w9bF4fy7LAaeqLjE5MMP5A2iF0CSB62061ETKQf
ZP6cX/Dm9DrjM98Q/TStBVlUQzspMz5hkwwTqGD9xlmYZq178ZssHJbJk1+sPOVN
Fp6FiNPFQ/O+MvrC9ITRPOO3hkJvrIQV7Co2edXqFYcU12C8xqaa/lEA+c0Cp9th
YzAq4Dc/RKSKzoLrFWFkYJbWS7cBActWLmk2X+nSLN69VY0n8FYfXGtrd1NHdImU
4cknHBijbR4yejWeC19ZSmHDXRmutswPWwacxLrYNRiwiTJLj6DDsHJCltWhUU1k
ketwK1B0r4R517XgJGUyzgwdvKfXst0N+9erz7i5OIfxNA4Hg353sLKDEaS40Zs1
2rEWR6moX+zitbXg0bdR9VDmTdACiQ43PA47Y/6sC6ABabRXHvDtGiUw5Zpjp2gh
iR7QuqSMs1eNFIzralUjVbLxQYa8lBBAMTMsKcJXXpICUJn4oMDRfOAAGM6W4sfW
Z4l7oX1pIFGuHrqlS+9TUS1lP5CKxgWRTIq7MEfu4OxibXYbM17oLEzynrXEus4H
heDWsSQ4vKmxJaqYTf2tAzolF0ZMUNej4pQhYJ580RalUa2rfyoPHLDcY29d8qdZ
rtyNXI3JjyKC15a52nIVgkmTBd1EmbIi8E1JURdNooRpy8FgK91HvtPSt+NiOl2S
Ua4FT2Qxj2kMi0e+uBtwyW4l9KU7eyPI7O6ntRS40+ljsYawq9jZbVYNI2mWUpRo
IIwWhXOXgxjhkYhi5k90aIi5Tzm1Yf1jx1pDNTNui5sbrPMLonRuEWjDvaJTq+pj
UZzhspWmxAoIuFN9bv4tOde++XFH7UB8tCktqgp2rOX4duL08Orfrw8FDLm4ym20
2VZnivBBKCcEGA5z57yqSmjFfzzDfuLgdlDNKfk42rkWP3GTF3ayf7ZvyJIckk78
CaJfIqM9IwLt0xB43V9O3awKQM5+HM4bYQPW9Ph6VjMXykqdHmEDDmLBe8ahTjdH
J3pNweIy5/p9LONNUhrThEnswbRFWj7A+SQpyT1MV3EXSazlCS9AO25HN9lst1Fc
pg+aO2rbBfQ/F/xHoFNeRilGYxBj2tukIu03FsRYxsbihXsylpIqQw3TkbnkE6BH
jqCw+cXfAhV0FH0bqCVzyQNN0zG9sOs/Gkl02V9P3BQOp6ysdTeVypAZKOre2+JW
atPYIcdrmLcO9RECgm/+AM5DSJ8ar5bQ7se5t6S9Gyhmgg7NptC90/9qz00rRKh+
OYZOCoUQVnNnsLWKZrGliaffvOYDkMBFjmeGKWwes2JTyzW4vP1zGA7GHzhPdnBb
AMMkysGKKxch5yaFQ/PsK8BvyJBJ9r2FVi1+hiA6H2Sxj0maBtQMHTbdgyW9Ut74
TH9ZtX344deZeLGQWa2QKPHAqobM+lPNEk1TFIiKSuxXIi96PZy3DU1LWyvMqzJX
ZXrVtjK98KtozVSjLeCokBF2rDYzeiEuu8Pjxof34KNDfKnKXjHYpGFs/LzSAjFE
Y5jStynaCtRaORuNYzyWD/rED4x/FltA+616Vya0Ub6uOAixGmkhG6ckhhhd2U35
iHMq+ugD5pg8LOkALrYYJlpBqnH4laqBZDaAxtPfc+yeazmqh5NBBpcAZIuDufa7
8h9Dw+BeedbIpVtgYzmzC6y7lWMYbaGnzet+Ndk7gxscWb8aJsh1cmnTmxxkyI6y
6vDwy7djLJmZD3qusnpAr6Oxi2VFH4STEeMGXsY42VBfWqBGhyYJPLuN1VMyDgaa
Q+mwcdzw1lhTdMxuZNyBPHm8dMeIlXrDtUWOFz6R4lRfSK2zuhfAXMWO6Yh2Yj1Z
cZnTn0deJOU+TVdv/r3sGorU37rehD5whbvVtmoHwPgpcMr3zfR/JEFHZe1AkIFO
e9OMT2VzMrURDNONNwlEu3OZ+IyYTsB5jSxMMj5Y7SCg4pPQHvCjbZtbu2dWemyh
YLZSt4JGB26fV4pO0QDHnq27unnBGQF3V4WylweYxvRNkHntpTkbR3kGkEu0QaeE
cD8nWmg/TpIns+9nuH87eT97iciM2Ucey2WfJk0s3mawO4BrAxBOqDcdW9Wf2t8X
x5bivcJMnWM5GeVfMYXAURi9/ByShvo1EybFKdtrQhbM5ZC7VOyU1BbLw7TcuESc
NUp3Re/Y2QLZVfzOSvms4wr5g2jLs4e6R+0ZnZIqGnei9jmJ140IwowobvOIW1ym
f+RSeUMRGIXutaOTQYE44KstjZjesgKtkQ9E/6au3ViGcw2t8K8fL05cRMAQ/Op9
AwJYspRzNxZ7DSDq+mh/QeoIUjiVutpHctwkZyG3i8Brs6TvRUvJHKEKaWw2wLJZ
qyG6PuD3A0n5kt7drBTR5LxlEl+ZX0MhpxkTvTmrUX9hU9ZS+q6KwyhpCtkJS5/F
LLQep6V72NAShOj3drWLwQJ8dCknNOLXQ8jMdOrXqmMTSJDGTEtyGOojRUxJKuNY
D6+ZfHP2wLTrt/53hM4sSB/zej5Ba2+dd2lsDdLYgsIpQmjs6Fw37ZatN/3e15qm
vPY5O7zcCYFv06PtD6nTAjWL6k1fJxFOaO12dLmHknN8Aw6ii2FpNiKMrVpb+CcL
gbh3aOz+rB5NUy+bE6i/rYVDa7B5lp7fTT4fRHzWrTlAB4FC0vdic5biGNfPbWC+
9gW6eEhWR8dwzwBmBaYqEZk0ATQ59yPBUc+oXNl7tF4YOIhZQpkIXx8rRJqmn+iZ
`pragma protect end_protected
