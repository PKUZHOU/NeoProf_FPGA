// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Oe+fkK5B02FKZsfjzg63Dbm81j7O6+tnlfEicEzKufGPoMdK2XFR7TesPOhx
GLhOSuUCH6F1smJvDID4XIvLdFgYRQYQzCtm9nmrTz9JxZ9Me6IZh+a41nJg
QbAq+CibvnfLl+TgYPXBEMYtWv7Ih/Qf3gSCcURR1/fmCzzeABeeN9hf4aGM
jgORvVqit+kV62xlJr6KCo28085R/6A7HDkg5mKVWoV3K81HB4tWmj/D6JDu
fFADc6TSzgexC3fSkfkOXvRS2DPrR5HvBdAhZkpLRsSURy0PUhc7+RTIJuND
e3kIrqUU3Ez/zg5YFc3Xs7/VE/nXlZ8PdJPgotGLAQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bb0TN+V9SMDgddPzvTymgh1e12KkSXWWdQncof181Bh77lD+vLDbf8685JDE
d/sM5NzZwgAICGNMfSfoDVxLJwuM7aYb6FD0qXCiW8mujLj6zGvorCYhdLap
pGISr5tAHGHGnImVZEkxsdUOYaa79SxOMnH6aNRyug0Wo7tf8yJJ2VHEw1Z2
pr/eDVGhZuWLSwH6nrEvgw84KzhQgwtvVuLjZAWDySuRwVN76ZZ3bAXAUvUv
hK/mUx4HSrrcFF2X22B0XPssw9PGs5aNj2vacyI3ghrt7JfmsDsKp4ORhtP8
C2PHSOwnX8mOkSasWNShnezsZE+mU/6dcRz0PYVYNA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mWMjRb6kx5pkgo+PMQRHDOJPVGQjDx+58BNI/0T58Wjmvs4n7Tfmt+zwOcDh
1dP5fy8Qh/kj6Bw8wLb794BUqko9xGf1y0UqSW2aVgY+nEX7d4CxdHVcSKbR
by1kIiHQscTi29dBj3qmeZ7QSz3rWfeVEm7iZ3YK+j6Hu0XAeTgOi+gm4xaM
ZOgHlIvo9maKH1CAJ+KdXLIX0hXxetxNQF59Tqh+VfYnjj3jAGhsgozFsW16
/XwJBxZbe7sViGgvC9chCpdaz4opFZxEgqPvEaq45csuVR4Kxf2mabPds11N
Xsjxkr3/z40iXWayx6ojMv2LAOSTONE7vGR7XsMtbw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dmGZeVwuwagGYtibjy7MYp2QPvrWWuLqDBAuH0bRpxmdpPs9p8FB6zCt2AOj
q9oMmZDIEdxUwRfoZufkSIyR65XJpOLz2KVCr1FCi9E150OY4k3HSsfYymIN
tk+ZxXA7qaSt718iS8dz9GKM5WIU3naaEK7lTg+yU0zjw8prBB0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bMgot9l1y2UUZUIyZn1J6KeDmE20smKA70diAO8jqZUPovw9Ibp+eGuymb2y
Jm+rGfgOXEVHYXn6kBeRBnCN9QdQzyA5BLnQkQBz1B9EzBbNrF51mIDXslSq
DtWpeXeT19pLstl+kmfFqxThYmU6MRK6JZCGgCeNENqwpcDtIiLk38fLVu/k
0ahJEa4e3O+wwQ0rTOWBxOQAZWzqn/an1cFB/ssQf90Iv3blVrI/d8do853R
hmUpe1t/+1jonA1757XByOs1DfA2Bob4AZc7okVg9fe2jkcMnBA36C4pA5Ka
dU8fgJ56Ru3k8sDenHrWTF/9dVScrI/kvtGj0epM3+IGiVmBDIdBI4q9PzTS
BVHFUwCwwPLl4Tp2yGUfOh5L12sr1bImK50117K7XoDOE7yTibDvFRZgwM1t
J8n/1BoyP7SWrzlUagNKqnFuvPRUu5Rvg2Jj7re2STDJpiKunFCrtgSjTffG
TzWdp4nWc1bLu99GkcO/ZsV+gOqV0JjO


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RgNMAvTwgQNgH45lft9pGPI4nKqMrlvSpWCQhj1P4Q6k1rwgrU2eud3FbDTl
z4TSJJTrxu8jwFL5PMOuMB+PYQQcJpyNj7ibkYpMKeqyIeD/K6tC02z6QY8p
/yZTY8IeZcvB1Xm+HiWmm8sImMzY9VUMnbn8vd8nk76t/TXtpjc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qn2lTfEDtp9sAhH6tLbtpTBBKZL/FNLsUC6R2BQs37GYdqP7CdOYb66Hcpuo
ZBFrkVqZdbukcu5i9t2f5s93lMsSjkb3MfE2VxF4TU+veFHh3Qw4bEfwWdko
VNqmCCPHW7JpTnYhLLNv4d8cdWfQw/vA6t4HdnS9JtI/D/ZjCJg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7872)
`pragma protect data_block
yjDqH549bGbAzjAion9sB7kF7XUiTFB+RpJLX3jjwRbEZsujbTNF6TckTy0O
WcTj0aalgPNnE/i6cw9/W+3HljIpfFItdxpybQGVsMG4dconXAa6/qfsSegq
ZY3lCJYXnI+aIFJ5lSWhpohxPJo2RbXGq4pZG2wT9TMCh6/aTT2NVvDnNxxE
LEoWCjnWcvh9HnCQmm8SyXTfkxe7j/a60HUTnYV2Jwpv+n7tuBR6oYE4DeZi
Ky70+3TH2/DlXOtDxrf+V+COHzMC6YJ5z5FmZ3w97jTDtWakBrjNrZLGcTMp
+SvA8QhvYwA9vPNukQ3udKKyBAwisT3zmIQ6JT06aZlyx5z9QV6sH2TbVKg+
EAkP5qXrLj8ciYZ3Qxm8WE1XtBlAK7Jko3p4v/+WNpavNF29yja3ZsyxRugU
dX7D47yxiaCYorqjh+Fc70NV0TlUTovrffmFTI81Dvy2aw7R9LrXFhpoCNO8
F31aaUFfN1dfWVpBDJP/cUO8e4Np6Yhi64+JXjHMjKn6oUZ9r8o3YyV+C6PD
zJqDm+14Kyd/08RwegHo5fLrGhQ9tjhh8S5L74ClXSZeMyKWBNoGxwx4au2r
lYSquxglpHi3JtjKyLRjdBtyFHqWZHoRdYjnFtaAAul71i/FZ6s0MD1DjRy5
6RYmaMWfygLSH72nWktUJpJqZ53Z7i7xtIMPZYv7J1ABAQ47AFkYk8ixP2i3
no4p2XR8Qc99qBduhG8Pxuhy0LnaOCjCp3Q8heRiUTF9CCmzOVLDVQt43BsO
zSvAl+CZOuqgFaAUmM/MmYASLvCJQ0CyeGD7V3wOLbYSK1LiC3DFDZGyYilo
yOm47WxbqsJYrMxyKfI3B0wRW2ZsXBVVIP7HcB7gZVJpXOje4KHAVRxK6rj9
kYHTsAeOLkgH4XbWs//7pgYfsLccRO/CHTuZIt54BCru14suUS2pkgJZtPPy
SsoT26VV+HLxlzSPtuUObjPRO4b8MheNyOWwu8frAkYPMcGAA9tMISU5mdpf
WfwMiqONj/TbYfA4CzQTf1DNE4alzXHrUpXveetQtAW6yzV0xUvR2nVmbf8g
ek7hxLqHOTsm+2xTcgF1sNbdYkYX5yvdw/AwDh+L/Dd0RkS85CjldhADZls/
p9EbJv5IqR3cqPErRmXWRNa+cbzhAfbtat6UZ5NoN5SPYmL8jDopuaoYIvcF
Q388fZruNKM+jbTouaVqjtSwavdA56m2BOgZrJyISq3b2o5zqw9cd1g94YtZ
9Z/13rC2d6+YIi++kfRBZnXZZf8fqUVLBdfedvmdUGljGBuhzM9JOzsjtjC/
WKG/c3dkS7/R902xkNF5GRtxV+Ihn1wL126BvP/LQ03YfBSMGbcbJY+qHcO5
ntahfVweux4yCqdXWxtpLnCpMGwiUW1bMBXAcbxtKw1nEr3VUFbJCG8aaUge
ivZDwNUh4ZS6iSnizfcjbubBq5nuKEJhu8DzUqVCyRlzARW3ybjNICWXYtbb
sOq0JTRwdtAX8ZjgqUKkesWQ+rqibXd+eWr7Xji6Lh8fkJUE4TzR/IOTFWz2
4r8PJQkeuWQvnfIFOFsda0FD9YH0bXuMsAyn6Mk3ioksCXrwzXLDExbYrrnV
R/WKpYA1Hle2HuOMuihII0q3F0C00bnR4Ono219SZr/AZJBQj9iVRdEwy0y+
5OolsR1xpLcwjrR/lOnLytpuVxcpL8LNZFMqmeSuOxlOm13jUBpZrqezVZo1
vNpKgW+d6KnTbHG+ANr4lBDZ4U2ddRH+hioIfYpCNBEoVzYUIU+mNQXqdXFL
9HoKDR/ABUK4DxHQ9xUDlS110sldU5aawP+1s/PVWxqbRK88qlaZzYrek5+9
Utt4rX4J6Dt43IHlQHLKdsMfZciH6hC2orfSrqmlJYwvfUqB77dbrNOHPy/M
Dutkl2YweOcJN4dsirCSZ3Ncgr+t2rFbEn57ZiTCX+bakE+zU81MuW9aQZuz
P2PxV57tmBQyj6rbxs5Q44bYPNiRE/Na7LshJo9pOI0jtF9z8nkZRCHitSy2
7XxjXRbzKRCcnf01BPO7xyd5gUTAdyCol8wloIG+AZe5V7MonPZCiaJxFtlc
MMIvESjbmr6p7P16q4VuCsocgy0W793sSyNcag62VvV7WzNa5dqboJU9MpUd
geWhlIj6aMRe9cLQlnBg9m10X29tvN/dcpwX/9gzbxsAyxwK6CAg1TTC5LdO
eW+bTtBPoV8O21wfAEHWM9ZqMRL2mVQRw+bx6ckiLNXf9WJxafFoDY/CFPiG
pG/+i0bUKrvytW8ZqFaopkWjJaIBa1KS82DTwnXNMdtWThVyPwAmclDoSO2z
7VMjt7XR7KNsRp/NlARIUDqk+JHQAYLIloFl7rdNE352R6FMtRa7fK5JPFuU
Afv9T/6a4vTdN1fUGIFYm68L8sx4nMkJUgousBTbHsWJuuxLKDGGgORXUHrh
kUoloCZOwFwKfQqrs/Qyamjk98WxYjxb7xIlg+0LYTqt2cwu11+HPdPKl2UX
avFQuIG3p3JrcCaORKXdLQ3JU3b5bkuXEYu82FLnP9wNVTt/hoTDR8aRYQVB
yeqF9RrxvaVn/AxACVzy5ncVNfcsazIVpZqy9DHog62NlNUOXHhywX4CEBu9
09RIYH0ilH8SGUAb3qoJQaEjb/z5dQtm63rJ212Wlqoy46kiMnZOS+HPuNyo
oiPUrOQmfVwziFPaCA7M66hohvOvvll/Fh+W8PTPwhGll2nV5FbtROGLaa1+
LSFWPcnAknQ/L3VlzscNZnTnliaRYRfBCfChPB1gWejec7oRM+n/DbxdJd4M
L9ydpOtxBo3t7Y4y/8C7ysXhBLiP58mJ4XMQ2RVJt68hEYYPTohjH4b5qXDh
WcG39bwZgod5Rhnu7iiljRQlSfhDxD5zp/iftN/FrDFIN1bsTeSTDfdOzWV+
2q7FyqaNZ1TEFT22bQEJlxPNejIJKBOo68LolPtSIbwhJ52UujEmXOJwGREy
42LM8a/lpTlxErSvfQlurxInXYjMT1V9Qs0GApeKUGUTAD63vVyWeC/bTf8P
Y9UaijT/DcvtTIG8PpoYw99hnuCwQT6XFxXpWdw31kLgDrsj3lhCvDi4rAa5
SuMe/82kDX/CKeY5uekVP1aMQ39drxsdFAZ2vKdX/c9FyUIdeaNJYOIvS+PU
TIQCt71fSvX1md7PYRlnkHxctB6M5JdWddWZv38sl6GCZ0yQeixA6Mb9c0uj
oifYUcEbgje1zJniSOYcFBCD76RITcqO+Z2hJi3XA+MCwSogbL08rLlqkva7
n1uM+scFsLEAfmU3WpFjfYh1AleSQzccmTA8Bobfxu/W7Xjy7bzRBHMpq++6
y19MDLLlV8zKiN7aBTwo5NGOQl8Lqq1b7KF57fCwev8UgPp4Wda6H45xpINL
HEILd8ss9HvQYmYmY0dZa8xAaPgC5ygUdscu+QuoePvucLrpdz3Fda8FUK1G
9/QrN1v3xgczXTv7om20L8D4Wx9CZhfBBYZmVZucP+/q27coeNFTxzmL5Kdd
G4AL6JOO/Uq4nrVtnTNLY61VP2+EgYOQbbUEc44oju1KLefgBWH177v0rIqD
VKHEdIdyqytfEjX7qCE90Q45MDvsK60Mk/5QvOMaSyLILgjB5z2XtYWCORty
dvpJsrG5TkGJQ+BQJvVTmqnd9BzJRUZh1biOU0G8xvoX1oHgkX44LrDq6xsL
8t7USrJIoRKe5ejeN7E96UOqELkKAfCFs5llL3jA6+p0PfbCX5WekrXg3NDD
rjz2LLZIpA8LXVPnc+SC9Pn7cjK+f0hy6F4NZxbw59vMYmpRyK+iupdZziea
WoD1xvEAYIXDMUa3mqgPebdCVcIuu8YL6zDbpeg30WZSOLdK0F/wIeVrmVgU
Kg4QQfgJ6V/ZvwObeVE09NidNo5ZXsIq+UuLRl6P8owXSsZnEWFYpvMEHGkT
/ATAy5+CSswahENyI+J+oDWcI8v9sKlfdP3/d0Wo7tF9aRAjA7nE83a9qWYe
bc3IJx1p/M5LyQr3jweDIqtfbV4lclMCa8lOT+qySwtmPnJEmMuhHXGx8lCk
u5j1GMms3EzfQ5li4UTsZnMtg430py8AT5W7UKBXnOHA3wAlUPuuGhWl7U29
+R+BpB2lFePmYEtAgx8ZeCmlMbrit2Zek0RC3F9uIOhNcncV+axbjYteyaFC
zR3g0TW7z9g6JKMPW6+y7LxstbGNOKytYW7GqGcbbwRi+ucCiqU0tqtdl3yd
RqJWOwOYAlTr+psuevHI9kzK4ZneE0R1vtvul1KT6zfruhHA9xS4/QIcBbsx
i72t+pcMRUpXMKxncrjaMF7PJ8LMFINYJ7OiyGL6uTHCYNTkPitWzFe4ocuG
8ON4Vxf5ytKM++hvOIGZFHdaURAXiiNaMFhfa0onHUYZcL1gj4J0npkuP1Yj
5wXP3yAiZsfXWSRNOEbcA0qRyJ8FuyU1q8ZJL6iM8LM7921elwmIN6l/hM2B
gFj9C+5N904haj2D6PHOBgWmYrYAPNeMVZ0gjWqbQteYJ0SQjQr01ro2w1+c
4+a0AKe7xVSprH+0SLicJbLWnePDxPKtwBz8GK9//1d/FrI5O3K7vvMBaQGu
Rh+wbKsbqVLut3F/h+GoBfB2ujlpfKYkVQz3iz8KxTeSZwg9hihnxVVMjGbU
cXAJDVYTB2/by00uVb/+PJ9rzO0FSApL4AtBoIelSVW6EH1saUbL/ZvSukB/
efTNblu42XnfdPklZHWkeR95sAYGMCV8c59HTJ3bz4Gmq9uK00r0CZIn6Ihz
OydsuSvTS6FaRfo/vq4AKmXm/iHxMbfxaGgDXRvCiuUnIcd+hyUXp8SdUpzy
5EqnKwNAW1cMz5on3aU06D6l79k1MamC86IYCtp3NzxdmqUIjHaZWZkjLUlh
onFQfFZepPI0jmH7OW/j3dXfjLKAwqPbCquVsaBmTaJux3y3xAThGEnNjsFs
dqj7tzP87g+D8DDyJuV86Lx+fIri2XicRHLz3LH2PIq4h3yFONOC5cCyqcH4
AV5SnYRHdWV07pxu+sOEL/9kYBa9Pz4h7nEWDkPuVMsCTt2sLoXzbzyg96Nx
CDxfNjg0ikHeWBDz1PjgjB0Wxg1YwZdm1wBFGAzfKoAz6vy5GB9dtpYpssSe
n7+5JdsdGVBtKOF5uxqHovr3iBQmr7wqbzU1mEgqmGwXt4EKH/M/lHNkRWQl
Ym5Fu/Psi0qH9LiAbr6zu0SMvxexth2NFb+pVl6V2iswswn0U/mImfAG7R/U
D1+mPbgggr8HIWiTxXjJ+BvI7I96iiZQz1wmrWH8T75SM8U1g8CEb4tc9d0V
ijQoOKfYCeMxcZ9gb47xPGwoWFN+xUBfRMsgp/4qrDwe2QTGeluJtoCuZiFo
npXqHfe7Z9kfJFu2UWIvDxnm2iv9BJ5ViimiDkHAFe/MwVqimNtOIrTb5wdJ
GFvJczo9LkPO+xAWhbG6HYwiNV9DbLprwUbzQxNzg/7vRwrKyt27vNHdzrUp
Fs/YnawhOD1H8BLh2rnfpbFtOvjlyfKbOF1hMaqPaipMmi/QC/RoZJlOgFtq
5pq46zfzHwaiPGn+bfmdt8y8qQXg5nj6Vg+LNGeJitYQE1K9coOzZcHjmwV9
CeX9puTG7OJnF4VKXjEIDTtD6k4BSNHnamYYoon6ToYNE6EQYykDTOwk3fR8
JhC8oafmzJiy2CNEcOd2tgeLR79ATLi0FRGeF94YCN77yBtDCwzoKPXxIPud
5VTbmcVA3imDg7Vd7cINbe7pUqx1NplrUAoFbxSljim/bfyl5yiI+NAXF88F
64b3B19noLDYHEZeK9BtbTVG0cpI2/Xro9GsqyKXXljkiHzcvjEjqRrHMW6D
589kLmDWV0LeCZ7BuHXCOV3sEngfn3pl5fVymcJEdLIqTtYDOfWGkQSwkd04
0iKfysQsShz1rcJ29GoKyhXGaeIUTHY9EZIok4SUdL6haev7XI7rZQWqkcuI
F3aPSMyOpwQ42OhlfxdWS2aECgMZXAat1TTHVtSYxrl3xUQ8oZmX2L6bfNq3
OeFagR6MqIgMs59QM096Hl7U7nvNGQdbIOrVW4XDew2hoTVCCxRiB8q4HZsZ
XpxV8ZhYapfBSDLjSRpFx+m+EUeyoHiOa/rA5fLdNeBCxsfIcy7woHRIbmzy
DrLUhXWxin1SZMa2vFR7QPX3p/lpCswrkF+EUisVpvQfagluz/MJXCbkW7V0
KjmOrW5q7RkAWB8WREMqJtzUD5U4tvl4KYGwKnkVX6VQFKlpXx/kLw79l7a2
urofh8fWAHqaO/ZUe4cYzgtkgUJ3S0GFq31hurOD2MeBNynwx7q+ZmYJx2Iz
QR1/0zcSoiXmCx52R8CgMmzT5K+PRTCq6BkMHyTcjWJzGZBifZn/q0c0S5GD
TAb0wRBlpyy4UoqkcFceiYDx7ua2aTb4y+sM9Cw54E2THzo1fb0hyYcRvSZ1
NhHntCsD/ykI5q3UTlnDkVoq7ZpdtStVsjYw2G92ybOiNfw6L/o6ounUwzmk
vzuyiu10EJ5DDr35Elw3SOKHTuFJPVRWPnONFi2vT7igK3Hlkrgmir1dKdZ4
SBWgiZgXqbRtYx8vOX2xmosscnFYc1+YheinzFutx8QeLfcVAW6t2dr+eZq3
SWt4BMdDWK8FyaK5bMy8veC5JOLoH0LXBjhCBOvga5xI+TZX3deVK6T65Ez/
Ko3XgRwVk9ad/SaaV1shKyB/H555Jxj3EeifYzw0tyBCCfDr9jgX7TakBsj7
Q2pTzzjbpVqoP5EE3v4n9TXmenExwssQ/86DzDy8WoPWxEvJRt5b3Oruk6v/
a5r/Z88lRHgds3pdmVP46VjiRKibS9oj82euJfBxNlJAlPw6aoqBcP7mVWr8
87ER/ohLBaLtFxAuSOmKcVwGXWKeRMNMCfQW1Me5KliG+KCA1KbToPxC/z5G
g8pFtCCy3Uoqa57Bmr9+NoQ+Tm+AcGf2FBC0TWZ78kr+BDOHcqRSHU8f0tzz
S4Jc6/whQbfhfhw/fJdllcaXkCzVw8bLBdTzx6js009zbbWfyFYpzunMazLx
5zTkvuSyMVhYB8jlO5AOx37zRaYXqHfBcts+Zo/lMXVtGxZIS9dyK7XCQ3mg
nWpb6ftAeuX1sB6aErYL2w1qlg7rrvLYmS8FGGCIxDaq4rSi3nmCrt/Ay80u
n7JX72/L9AeszbUthKKKAHqbKlnb6q7PAHwRzqhD6jEycFcOJSvLZPHE3k1m
MZrZ7orOh/25AU7K0pa8T7YFvGYjqa/cH9Jht9FOKlSu1PJ5JBPmFuPbhnbs
EsLoNJeN/1+tO5neGKZoEwfM/3R/Cwt16MGPZXTkCZoXqNxtPsjmnNb7mki2
X0rEaq58iswsDIszb/YXBXMDeEkdL50xLw8V4eJ/BvyB53mim+WatL5HFl2l
L+jST3gPZQuwnOKyKYgONeVMjvQwe7eT+klvRRkZDTEhP011UcUHZtvrFrTv
h0nW/wNzvtaHoDESXdfTv2m5ehJeLWa3OX0dMBQs/OncEdlhMiU+R74ZwNSQ
ZcgXZfNB6jo4Oloziz81Ko3EIOzZBVlQv0vTGrpGYoUAw2xqVTTDA5TH+7tu
9f4qbRsEP+akQD3F1yZQBswmMR7gR26wPjwKVI5orpc6E4wx4QKJE3+59YQb
Q06vLSksmsZ+UeE7Zn17kSkeAawY4dXFUy2okHJuSyl3sZpmcGSJNcVUitSF
68AU9KmH0jfxA/8Q2V+wRpPdt573wfQTcjwp9Dkjit3ZqnEcPvnx8A2Mhn2w
f7pKlNypNA/P5O4sgna5iDb1E/SS249q6fQqebVgx953SngJlJWjXe4lf1Oo
YDXlauvVycWFF1UujFH+0nVaJxMpQgPcJYmtxYzYFXbPOW40oljyhQeMJ4Rn
Qq0TcMEDh/HlhY5nW/n6/pRskuZ3bwt390EaEGPRIoui4RjxlwsJMgvzydxb
71O8byC79C1c6dqBb4su/6BmTJkxqJ8PaZBwt45W3LA8Y1AKSbj7REO75rAb
vICDjz1D3vuxHaLJAhDzIFvvQG7uUXbT1iOMXmAYfWN11EQ9+IWWGFEM2Ixt
iIJlrKBsuGx59pDFUZUMGY6jg11RybDrRHmggrnNspxYCbdHVtm2wsayzPAJ
TvxlG4RbHSde02QL662rNsmhBoqFmg1T7h2XT7D0A5Ma305J0oPQjXTWBvOr
sfxXA8P4aiwkaknNKg7iWaapmCmUNhndAxAD95e2N/YYo8yfhrr/yPL5uVn1
O/8vTSivLnPhzuKaUELsLlqv1FyhItZ/8VMvLk61/OY4ZGc/mDPrQReHxYNo
h13NNOerrjZvkbuiYB92+EwnifMURsQv05+t3E/vDFF1dfQ6o+Cpy535NwRf
+3h2zQ5diQSBHMiBHRDFvXEoBHrd9ZwUUwKgymsRNLtUCEsrGLJJhmY3Apjm
Y8MavPkFUELSeqNjaEH3slRAa+AnWYeW2NUpOwbvDCw7xlokA+nV4yGLnuqo
62SJQQogq6Pcx4VSzLrrxKHaYr7XtcLLKGcFlGjejKtrP74KfDKIPGqfkiLT
h6Pmpbg4uvfAyXYaTi9IW5V3fdRZONm8E9c8lpySvNGA4oERdvYQ+CKrMbb0
baRZyAlTOgWBmaAMmurNG+pe8vMJEjY1ma2hE3cCK+sbbO/1zR6yvva/PTet
DUzhIuoEiauOhndrWnmdwog3Jb/7Jm1gRrvAt/rVmaZfUYmpdJFFcisilyIM
pvUoF6DR2oQilJjQyeVdHp3tFbMql7bVeu/uVJR2hDrOn9hE/Ig95NQ76yCi
zAqZe49e1Bhwl1sm98GaIrtYMfr4CXDRkYWDguCmtZHaJcCxpdfcGtWOnqQf
tQXeYfpPMJh7x2TvUFNAFOSLTIVIlZZjJeIf6JTyZpgxhHlMxGA+DUs05W5t
ZBtl6vPmqpk+vX8f0WrtJnD/gSx5HO/CGT1ROm0KfX/Bcx1MjCYN2Ft4BV+E
g/Qjt8hajy86cxzs+/1ycBhNSrWDNCW30D2hv04dq4It6bhppN7U9oKy9/dV
nTI58ID76CkI5P2o2PmJkvbYGBhvSTzC+1VWGaCsDDGwfKVliGTT0dA8S7Bk
t19Dh295mO9NypYKNa+a9DD433JTgJm/udnT5GssGRVtp0cvF7CdkewUabaJ
cVTQ7VT5NwZBoEKCYqViaMGfJGs7zeymi0vDOE54fy/8mCWjCis+TB+syiBx
pscqIsTVrd/YKQtYCIe72Jy51XgHjh+DfGZz5dxPS7U3wdkNXTe7sHmsdUtQ
JbO8pRQGJ+CcLbB8qLeNcClnmVidsq2BuO7MTEC5WUaKsO1yGyU+XdCDx4wr
AH00F/qDyOOj4g5CkjMjZ2gsF+mTQqOB/TtxUm3GfD9yUHzuVmMmiOHjYBq6
QFzcjEj8r1V/M07S4aa8cG5USAkIhw3MEWaJXI9mVHFzPnfnGU/0GOr4113P
pPyCe/bza/agPaiWtAo4f+jcD1n0hE/5PgpnK2dVhpCSX4Cyu2Jj8AwTWW8n
OIlJ7LcjH83Wxf2xx65PUrz+NrVSFXDsDrEzuunwHYy9EWtrX9VlDdadzIGA
GiSarV94IMRSHusrykcmh93/9PFV6bxrIyMFzUXkaAaqGGabqgxF7yU4Xu5d
6Rj6wcbd1AcFHSRY5WKO0PQ99791FZKU3j1TrZJcjMFXeB7qNP0b3kSRHLwO
NtF361+dBCLu0CHaZQHCGeRQ6CLh7/E2yJHFvLQY9c2wCvXHAd5mVFYjlZ3P
b0CfzXl7kYi2ASXOHVcVr1kkUMqDbISF1IdKDCnuKDjbnngxmBx35GsoUToZ
T5jvjkraaejYFoYK4ue0KUZ5qbtSfjHYbNUVkMaHci+pnDPs1kf5WsiYYr1a
mR5WWgNnPabtcrGCy3U8hTD5Ms21L78odAM8pus5kSu5zVzjTDYG4qFdZK59
T8/2Gl33RqbjK/9AmHY3+Ydq5RLy/HZMP5Pi59AIuW9ASEB9Qwk61VdU1cHP
Dm2WBjThmEqLu5Ymy1/WCHLiVujOVDHnmDr7P4+GSzRfoVyv46KWPj4G5sx3
wp+CRnx7cLrwADHQk4RX9CjKGstiModX2Sd6ol68UqrzuAkyovnvbFe9J1w0
egZdndqEIbn4infGzT6077vSxcXkLhdddsazUbZ8awu+R9mIC/zy2O1kz62y
IYS9PfqLfl5BkBDQuxay4UG9x32okylLmhgBkwDKz8THiHicGZFHp4eyMRG3
d3rkTntqv2kZ66GH9iUW+G4cOjTfsUGeGIKNfvZMnVkwF6OYELuOWqUNruMU
9HXS3SgZb4xYF3H+tXhrjOf7crf7F9ZqcIbGmCb5t8JsxkEbKeQwDTxDzoz2
mQrUBQxns0/N+ov5EU7qGsaormBr0vmuURIktkERZCGWxRlX7SPdd9u1oqqE
sG8n2l5uNvtM7THGbkNk9SsvBi78EYNoB8ZHAvrUUoKG7SEiVN2P4npS

`pragma protect end_protected
