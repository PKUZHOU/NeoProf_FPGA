// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
dkNVHnPMlMQSMnM5lRoWTQ56Ie81BKy6sipc0AXBLDzYDbyi2KAGWlBK4epQGcXq
aiNZ6QbH9UmEEA+Di1EnToxcLunk5x0joYm5ZhoMpEAJJ4C/W0xHeSXgOMOHfqyI
gM6mIG76JEaCaBc1Ov84BSoiTVchc7TazZlFbk+rUZcmSYXH38sD7w==
//pragma protect end_key_block
//pragma protect digest_block
j/Q5hrbUbGUPIsDQf8DCV0IwmTQ=
//pragma protect end_digest_block
//pragma protect data_block
5tNqM1xEVQXG+Gz4w3qHWhIGRQ+4YNZnUGMeuxVO/GLU3BkZ4JilGQR+GDDFOW9O
UsVH0L/GTTEwlXqS3b1PquRE5lcu2HjfEdldLBNgO7zELelqUOtbJo8lRFcVK5lT
Z4VFltiz5aTq5qEooHhdldWkTLAictIvRwTfeqaxoxxUffE+KcqgyrI+rY5ZlCLt
6Vod1mzZECQMZkV9ca8bs7gxQZNQfUx1NqgWchAR9Ao3Gw+RzDMlaDD5TIabLECA
SIlkCu1YYo9bq7fif9FPXrUhvcnwaZB3LZFaPPPYdI9hP/KvSTaxCC7Vh6MQXxnE
O7Llk0yxSCEuv/sEcIoiY1/4vbHYQx1uxacaOgWmYUgoViCeRmQS+19UyTSl+4Qi
aOteKBlD/B78XM1VJfxTrkxVMA0RdIFeoM5epP4RjQL1zWPWmRUNcLibGEfsJyAf
czQaZe6zrKOxhkpGhNwxvEZfIYcfkLbzQ6PnRTPPRLtBGJg/8PcjP7Lp2ujl8npq
CvYB/x3qVBKGf1hmHp/MQQBn+ih0xDfPHOHmKBcyuGS/qo1Ea3AQYn0Yi6xCuls3
HqQAEmvn6MDjU4+tOyjWWZpiFUohcuiamRhqIfwodLhvnYbeiqg4o/xWqjq0kbiZ
21SE2jbIBag/D+jZWpo3R3vNLDLVMvsuX39y7JEZZ72yLt2JTNdN8AE2+oYgxB0w
0XaHlEhTkvkLavODW6afsEdseG0QZF1KYrTwSUHYqwLx5o2w+lOZQsR92i0kCrg8
J7qzOddjNVHQuFUjZinLnkpnvwWXcqTZCvljEJFfqlT6Dffiju96nzo4Kiig5Ats
VIjH+cMvjL+j8qP2NWkw17c9xW8kAwMF36fiXJx8NueKPXHtPSIUJHkHJTAiXgjn
wiGvss/abw42tpa/oGQQJ0AyHKEtc1uA2fNe/Fi5b2mZGeMYtoEtruDPE/EV5vSz
1xvDcSI9F+b5UeRP7+d3+XFk7+beHwCNYRxVHuOCvmHOC8Erqo+zxxH86o0QuTZq
v4WxjZA886qkolsqc2svUMmRamTDqS1mywZ+66cKmrypdAHJ47AX5NQ0L7smjyxl
aRm3qrOXyTUldPW+CnFqKN7zzkDBBSSPPIIHK/eiOWtneFGVLs9ycdBTfPahkEEq
Pwi7S8dWrtINUMLpDbppsnxN0fWdfvhh2tA+w7ZibIFOAWx0D1lOmODN/2zl5CRf
2yZWe69HvwzIBr7ASl8Mu3etde7A2dO0ntULjSh+LNP/T73GteZ4c29VxjECcsgH
NYMQdrxoRWSo4Z1fjb/N84UCkmrlfI4/L8bWgRsrs9Txr/+wH+0kMQ3E1/gG7DZh
+vbN6vNdUVyiydJlWqYKza2InlQlNL0lRiON8npB6nsUgkL5iFlsOEJOIn/B17Rm
rxDmbMLTG3jrThKZI77DBu4GDpb50DmYkVTo6IpSATb6f74wW67HL2A1TROFlCOW
TwxW4sv8+blwTKlbpshp08WFoWcv8aVCKzU+JyxG9mWco2cHM383k5JbsPldh2DO
DsJksaNJvW5VpgX0O3MQ5HCKqJzK4JHrKRLxmZgrK/W6K4M1eDFVbAy85FdOgQdU
afg1LqDjKULqDCMeWDJ5nM6wHopd7LxJ91Lz+lMSQ18KzgkLUTEoMBvL6eGt5SLI
CQEZHqu3rSJgvPvRb2xoINuXlyL0rJ/bgZnRM+ZWcipkiRoYaH44JDBGvQeKW0M+
qbLuhkwV13XWy/0UCusVoIyKDFq4dWLSFToLx77S6FSE+EvRdgQA2VMPBrB37uAf
CfYdxzoiIre0WvVqfWSNd/YNy7XvANi6kS7u2sVRhqzyvuJ2WRnZLsLrsZyUUjzU
/hc5nmn02PtnJDDkWe2CTmaxH5HlDA0Qy4OUOeG0MsRWkCE4q0jgHiXEarGPPpAZ
dkSepIRDqIMSAdSlTvR0vnHoZAkazbx7ZeBmei8n2tPyPsvEMJWNJ9zumr1D2VS/
gY54tS/jso2BvGbbX3UOydUAXpO6Wofhto8veOz/xWwc+acW5Lx7sxSWcXyKdmmW
3ZVLXwgefXlcMTcTEs9JL7YNFHGFXj+V/kWMAlvSjEuwF4yNWPJ3ClTn+GEBqm7S
HhWNV/J7NUeZaqGqRWcmlt/46PjKAw+5DZVh9vlu0c8YNzuzQMYWKFyH6YORRXSN
RNTCvZQ1b7pY6HcP8UNASPzD9B3p6W51nWOmkUZGLNhxYiHA55qGCYOE3YNp7fCo
zlmI/JSWOsFpUywJ8ct0Cs3z561LI6YsQBc0VK9gBaYXzSGE31/AsxaE+WV5QXED
3tNSttWQi3ASgaONc8McjEfW5Psr0t3udaiK9KzWMSWEpxBHcgQGH6JGRVeeHyP1
uPhQRsROYHXoEzPqrz5dyCPb65LAYusRcswB4BP1FVu0vmWmjpaDDOsFsxgmVfJO
61Pz4l1JCshp7saSUxSHADDKye8ZttO/mTTogg3ZnRye45AhqrDhKwGLr+yDHNB0
n6qHwkV+eVTYBbtlP0ddx6arR24fNNN1xHnKY4jhFYY5Q98sq8Z0Pf8ls6R0Jz1J
1SimtAKwajal0apoky/kQioIXjEJGr7nwBHe8ZagsJIvGuR5VUl4qlRGbPStd1xJ
/hI2wxFOEY6bJvg1pLHBRkBZcCXoSplCjavf4Try9viyh5UcY/xftdlxajRtAj29
VyzGITdsD5Do5m7S1FRhTpEn7o+fgIve8gjvZDmguEctGJlWjh4Ci6RIUm1XEnme
icZVaLyRsENQXZZqwVzKniey+6az11zFODnB9+Y2brCtPgurPABYiftVgm7dOg6Y
TDS6p0dH4DJGDb8BtmUy9WD1TKkPkHkzh2m8cYDKUCb2m0Gt6BBPYAME90dNtiBW
eusCEGHpifcCZdI5uXTHNjRwWfkTQE3ImaANwrY2Jwc8YDrxbPYQXvabKtTm6vQ/
m9kWKziXipARhMUFfxqKzan7KIDastYnD06vVucfsB+alSlfzrfOlysfz3tgqrHw
JuvHvMkLJyRvDPL7xMOpZL2iqNUuaT8d2gZVzNmrBxj7G1lZqzhjPBefpMnQjWB7
uRuju7GKyxaJPG0F1L0GHIr5QKzOKImBhDb+3avL8+jEdU14kzq++JD99BZeNwTr
BtJJy0gH6RetihIOqcwr1TtfBEYt8B85dwwpQWSFmF1Yg3D25AETaywomJawFPbP
gQozkC/8/A5REMBhRapTNnxtcwx8rb/jXaMMu/MG4OLGnp99NFsBdG8v5AklW0X2
Orwen+jOWhgS+V78Tmd22gB0i0hEQXGg8bWa3MrxQqdWVBh/noBrb0kOmcFuMo6n
7Z1hyDGXzGo3kYh3novsSVHgwDGCGfbM9d+rhen5IheiLmb1gqaHb0i7QEnd0+gS
yo7UsP9ZgMHOCLb+KhNxKYAWfLqt+pNRwLZCtR5mYWXK+p39CtKTxPBNBALywCZd
jTQPHTWsxJWqVuWtgt/b0SOckxRDTzF3tbXbsgDYGHbjHh4vBsurMB+qGVDpqnIW
M9YSLm3N/LnIxfxyyp5Ueo03mhEmuyUact1b4y9rzwRfNucNS7oYoLJchx47n/rJ
KKeHoKUAn1rPJWwmCrs057yuEDEIK+POq9u9rLVlRYl1m0sZ4blPVMDY7e/eJBaV
t2+AM1T50nixV6a9hkt1Z/j5EV4kOsm97q7ZHBQm+CK9+H92oS9WCFGNUTqk//2L
WTv8hLY5uqYd2RtlkiYx9PhRhRzng50kyFORkzNJKUewsVoKozGsZMydu7K8R7Rz
xJH7MW5nBJajghTopzqkqxFhY+X0gb6LvGJk6OBL5dxDuTDYxGe2oGwI5uzdXpv0
BvqCYk0o6l1W9WFG+vqY3HGabsGFCbpO82AjMbq1mpMX8FjCdJnXXFGvUbwGQSMV
OK5M3qhf1bfv965bNR/AQaATM8BwxZNWscKbBY8EZqg/Vc7pCBIwe/+wiSYRirss
0eg2TjvaSp6zb1LAYkSzAcm1gljnJB3/cfx/KJ7ZqzbQ2a6HU6Nke+W4RiUoNJy0
Mcb81HFcx/2s7eUUJGD+Y3fH6bp6DAXSdCzlQ0+fsVyaXIQ8huq4kQyBxJoRIeHN
6aCxJC/MM+uab9DS0NVRZ7MQwP50XuBQQxLTN7VONgPeStVGm5oAdBYwX9QuX7Mo
O3c2WPXDL/0WuSRogs25O21XdkinKGEhcoDvQxV78nwD5QysdZXun/q0nQkcpEH3
yxy1jhCvd+Inh4NgDMaRTkYNnltXIUSiwyjQDg81OBmHOx+UW8ST92WMoklvTrTA
R1DOe93NOpD+SYYjDfr2URuM39tF2WBfNrdZC8UsHLj5Lq8WNcA0iJGx+3UAZvSP
vc9JbqGDC9AS0Q8vGCsOI++6JEU9bGIdCK1gM5ys3e0K8CpAIsHwiSRoTFDLMPo/
bkrj3hIb6rdI9R9GqBFpf62aSnVV+PdPVoTA/bxuQseR43bCGYH9jRQyFYfmManQ
pY0+BgcV39JSsTsWR6FmijpUmNrTKHli4GvdFP1vbCdn1F+q4iWv8I/Pf7tzIFVI
0XW+tPCKks4WUpLqwNGsHylx7mbiVtOA30N+bNIElFeph32mhtLGUZEygsHX7UEF
ijS0WQEodslhlUfYtyrpPD2wbP8XGu1TKIdtbfOpKBLkO3XHy/m06B2D7vg4p4lh
OMZaSJC69pBhygFBdkAx/tRDgOnRf5h6CUSXC1tHfqigR2LtZntHj2FniyJ67hUe
Dm4FSWTyAY9QdHDmEKZZ8uZ/noB7k0LshxUU3jyJH+njkMGCGN8lv+19MYdil4aP
1lo4HylikX+J6Y/g7UNwumpd2ZwTmINc0laIIM5VTRE1+jCezlPkJ+Ym+UEpnOKP
pDSrhFZF+C9cTcf5jeBRX85C0Zuk8vdZ4xzhnY8sRbBGUVJfdB2UvfyG9Iea0xyd
wES4WuILli7qSqVZxR+7S3Mo5UhxNHOeWoMcYbfDVL0hiAGg0YEvEBOO40GQsBtJ
27Wr7fHzu57YPkVLZk11H22n/YlIrw3hS6fXXUNsLvc53yd3XxuzLiqYwFudEqMc
j1wonbmzj1OUDZ2CBQXyuclE2WsSsk5EnTxexpDnIgPKz17k4M6SIbUup7qziPGF
97vsK/emOXEWq+cRAxZbdkGd2w9bUzzkTkHMm2lkEfWjpmOHlDCOdnyPwBgnqAdF
ZuIyfE4OIU84F9j6fy1guCoT0fxS+iDDLUXLiwJiLwaQQsbzuxo3v5pBqXvuPSte
ixQgqo7OrmLOppKu0Q8K26o/mCXiJ/SLctnjVjeOYi6ipjaSN1/0nazAyZhkm+Ii
S8+o3w9vNKywiQPXZ3o8VmkuBThGJttPzps/qjHk8egF06JUeWWFBHsXbLgNFRQa
PEHLBj159Kr79s99UHxDZ2Gz78GAH6L0sEC/g5ZXF0qiKJhRdanI/vqTvGjYx8mf
4cu0IS/t4x56o0hc2MWJKsFfZU4H7lUuUU0oknHB/4Kh+qO47FiDX3vdGd6xN6EF
nOPT0QOv0m0jnixsz+ek+9fNlRYtZr4Un0bth+1e6VZ1FrB4EMSbCBTQuli1pZsl
F7jUDZ4GElxVMBlBdM+nY5FH3CDzwScXNK2PGh2Bdzg0rF/sDhKOaNLCu8uQEuMz
rWDY05s6PtXvAaxchH7hO4u1/jgQu1nLJlVm+VZprWoNRu6fKZi4Xufp2WPVwJwG
9vdKc6TnVcm0R9ULwlVfmVM7KCXvnhE39o95dVt6nRRNGOmOua9AvgsQMOHm7qAx
USphcGdEwnOFP/cMt8EKxtygNZ4UIk/7b6awuryAgFrG90kog477BouuXqebxTrg
Ynu2raEFuoGDdOqhY0UTlVBH4CNUnCVkybPB11JYQblQ3a6hQ7eVRiZsGjqCX9FC
Rj8OlkDlGFCSB53AtOxDrKGjpQ6uv0ktpplBr7HBUMSD1A3DqgTLngOMFtHrRzII
Uor7rOqD4U7zRaswnu3B63f4GosS4G6IhWkzPu5tnlxmF/bfC58xjRICL2103QMs
t8/U/gxXIhDK67wFZLLZzjjUuZzSL3+1MaRKspz8OU7lBciOh0QLkHXAxxA0jTSh
WfjXoLdvKirW7OGrqWa1dbW1nk1WywSlDQ1UMTjokwmNi2iT+WBbbe/XfmdG+D1U
IOz2QlUSh7mhPyp3DmBLOcxZ9L6kBD+GxDQ75i0Dh4UUlzaWv8B+UZVPanohtj/T
V6s6Jjr94QnBL2cVNXWQ0uJcrKjn/zf2QtLNh/NaHr1o+29eA2VAxn9/5qXX6miB
yJWvnMVDFUHgnMBi0ReX2EEI95Pak6Agd+l3ToOSR2V9RnY3g0KgE90Qq4+Rm0K3
WLCDVnKcCyVY1jQTfvmV3ztKJmLH4X7dXGp9blAUyCciUhme2D6hQZ/o+6Mk2vGd
LfbBxOHS90LmoEGuprdwbpMyArz6ACxaMp4h5gkPATliQ1/8G2IR7grHVEgHuaX1
h3k9dxNXkpf9DgJUX+ZFsuKy1UJnAx2Tkpn5Dv8htj3pbLdiJbMwasu+8iJODGZE
UeZURrPW1qSGWtTgepox0uHGu8V0SJSJhAFDxQFdESVMw2675zXw218jHaKXVAIO
GwpgLLyc5DwjWqRI3DvB9PwPb2Ic+JrwS1364gkSovknbIw0ya8KZTDaZ8onVD8p
jtx0UgtS+v28SAYuMWmkI0R59QinJnyI7S2amDtLaVuSe2V2bRwix/tU7dcf46AF
nWeJWroH1taPQWhON+sxKgNG0uFujNAg3EGQ6bltMkBmdUU/u1h5glvI92Bv/Wul
RKfbmWvfmk14N1Tv+cHGGKsS4cLPpyGIflsPeMMtaj2gRSycEOibOJZRs34dH9ZO
WQ3ElVihtHahn8Ls9XCqGfyvyPwXZ2wHZcR62BP4lS2UYh5jRbI4voy1OOF5uUfB
1Ri8wXld3LoJuKd9uvA4DGDpHuBvS3ifXBNgh9vd3Nrw82Gd8u4/wzi5aiI7yxi+
4/55To+JMggJ1OsSwEdp282n2KlvBYuIjimYWo39Dt5I7WX+wwiTWmlRstfZ8kGh
U4kQGF5bVTRXxQbqClyEXC3yAIJE7FThkdHxeAOsCXkgApUFRwuelYZR5CA4NIQZ
+1CXEqV1SqGfiZBhvPcbSf8glaMk9q7wA6r4b7ob746TqZqL1iHoGQ4o/qbUWAVK
lPtwLejdBBgS7idV3E8DVTXIeYwzFP0XQziO02gVtt7lhCIJyCyrWzUaOmysx45+
Q5yOnD6hoyGl9IJgOgs88Cy/qv2e/3lUNbHBuOHmwxfNqAay5659alrYfgAdw5Ra
ieREmfOqUAE6BzNBjv6C7Qq2pUtq7PEoMXgRZIqiasGfNLMOAkYwkbJtsT7hsLGr
HiXIpN52Q3m+4cKTino4K0tj1bDHMNXi4NQOw4vC2PzHGfEzBtBkvKMbL7S+BvGx
KjOAvtgR7cNOcFnyza5rYvQEnrIm76BAYriz/27BXkq2iFg0WscgktLV217IM+E6
mVfxJ/WOsN2+tZc7nStmdVvFBSccMk7lEHDcgakMegV6+RclTPepPBC9cTl1/gKL
953NsW2vnhjNYHWPULvShyCpIpOQ89RhCRHjkiQwQPfo/aA7RuyU1MoGOYD4rip8
CnLdDGQs5ZZUeFugTVZqVKhkj7J1qP/7E5IN97aSkzsGiMdJOdupi78A++N+ltt9
osfEc5nd3Com599rixuIlb+yTYeTq2VclHr9lIzv131FQuIQjEC5iM8CBw2kpNO1
LxnaPB6FEGEFI2dowmJASh8E0REY/xgkTjyBOHpCe6ED0dmxJpqCy0rJETWR3rOZ
fb/0dxCvuYyCFYNpWR8OkMavTdWKmw4AtssAk11sw3qFrfHdjnsAivZnoEAeA4/x
QD7TYthpsN7SpveJt/ixJFDbabscXG34rdu1OkKYqRq+9aiSI19eVKQc5YTuebYY
7/xaw1Ky4/vhyucNHapTG4byRNuPI3VdR044oyhHyzC8zhLZlBZR4JxgqAkdhhzA
NMCwU6LStAumGUfDd88Z6PLhj1G0/UY61F7EEr69+CBBW8S2MNMlUqYOWyz+awSA
Qz3ufrMsFf3Jf0noQQ0e3wz0nL6H6qFfeGMenLC9UPtMsYMibq5JM8WqbPkHl7Ga
3mtpvaTkKNqN2HkF1K6T3udIsfaecaZjBAjoHI7lhZato5pcx4hgKxdbmO3zSSrW
QyT2IvYj1D1JLAMfVyG03wVZiBl8O5EiJNLkz2M+D6m27VpYg5qeU5xoE4gLsneH
z+sw84uyp+aXCikosFO/JCuATtKnW5bn0d0/JNNL7nokOHbGO2JlsT249aE4oCt3
KRB5nbv8Q43A5YEffxYPJf+t8FRaNeYEGpIWCpp832HFAFgrPfmaw48MLU5FM7l2
uAXuXH35iixmRa/Bq2v/Nd4LHkaSSVTmH9iKHiHDMzD+iB6pS3lLKG1bLbc8TX9V
ivQDXzq4CcdCoRDpvInZJK1yROho6DHfHAzOeS8H1p1CHo9fzRWCbw+MhE1c4Pk7
RW3qn2MeeXYmUE00C/xhxxByR+Vkp+/ifgKEJFezKqaFICuCTy/jGJ7hqAZDF+5n
wgf40WVeTMiPVBgtAdXuBnxM2rL+jwGDjyD0uBPRIj5H90vHFOYgx626VYzUiZwj
S77R7jD4VFC6QI3AoqDGFZYamCq5Ig45r5vUsSg9jYtCW29+H5RO5NLHnT0YC0lB
TGV0VsYDlX+0uSiotmQ4fkvjGjbGP4feIee0krHxJuKUfAu9oHOTqlQKN3eLNU8h
7RuKF7lN60q/Q4H8mqrWvJ9ck1AZ5USJ7hSYmqtuESCCBp3kD5rjd5MY437KF/Z/
cLJwjM3b6JmrhdcHo3zBe5+e5cs04RUXfyjmaRQOQYdzc/s0XOsTW/gIQMc2yfu1
0+ZqNy/JXDPpBeSaPQwDJk41VZxwso4gaKSZnPAiatqj5fn6r/6c1mULwcJCDEhU
UcxDtsr42QYuJuYkmIijuMcyxtsV7fro7JHiqCdluStHW0msjMAVmhyieN5VTCvj
ghXN6QmB0jZu2+h3W8Fso42l5y4QLp1QNrM03tuB2hGvdX0mC/GiPJSHiDVQazCZ
WRc1CeIJm5bQ6nxV3nszkmhukVzMjkrONKcv8kXiNryfUUQGAue+fI4JbWASl+1P
JAWEqlx+xOfTkNCBsibP5LjQw2YUBC6qdk0d7o7lPN6f0rXRxLaEBgJEK4NKFJJB
0ZfUm5+UbivylvrGGx1ARHGaLcF5t/hqLuJ9uR3kyQ/wZMqX4htr9DppbqheHQUC
Ik+TEBiGVk/VPSIJUK1XW/wT7q5eNrlarTt9tiN3d2lIrIq8aPbr0wkWVIVwCtu/
X0AZjX9kybY/7oxe/tB8VyxfVsRbwge5yK2hJvNVyryIYHo02hgQfe8GAR4rQEBe
fpG1bJ54heHtvfsgxW29yRvfqZ2SJS/nHwiVZ4dbJp/mz2gS1v1Sxx/1dpPdxU0W
Axjtcj/KoZ8oxVfFIrZflQout63PWK8Ww709x0O0Roz/KzIuYsXm9Q7Y9PIrPRP4
N0xrzybHcS5PZGhlWdrxV0XdeHkHs/h83LXJzN3Goy1JYht9Z9SMehk8R2XV6TRR
tOY/SR54sJ5iV0OJIRcEVM06YTgkiVFa2F86cOHh2FmJBn8nezNSIgyzM6XTVYyF
UE12RugsRCP7rYbmiap3FvFtRZ2qlr4LAwP+na9Jzwbkovl6gZeaOIGByDyU3d4q
Ud2h/2K3CyiAe9h1h0Y/vijeFRF7NCJqzroA296+u8PMKc7Bu7I7XA8B1LG+1frs
vAq5b6CBaSUk1uf+lmdyyuKMgwIXjsCXnneL2qzVya8yE/FKHQo4QTdUwwimhs26
1hVmtMAFiLzymuAw0TGBDlSqqTFTwrz4eKjTxJsCKKiPTFbtiYN3nwqVAzGiNEw8
Rf0gGffrOqlD56pLYj38XQPUfmENQPDlOf0EQyz4EHRvxDYBYMY8U3PX8WvNoddh
xzaGzpplTI4OCIDe318Ekk7CdJy6X1rdUPHijdZgrvP0qjcnGnW76ab0PCjwEkiW
QWrxZ7DzrCUALaTcqZX14elRvG6/uxxUmXRvCBH5hNGW8Y3NGLgNsq7iir6x/oQJ
GwnCfojdBf1CtdDYIkYB+Cq80yiLQiCHlWUDRyyVp6ysA7Se1ux81+75VNEAcPSy
izUBp/ZiL6KFqRQv1Ac53hR25Cp04zulzRYId+D2ZGtUQxAJhfHp3NJITrhA/LvH
TOlJB2vu74AxynnH/G3RnuKhRWwQi4vMfZJrdvdSQut/Zr/b65slyhYqcw7bXAEo
Vh5jFfHKrECpS52H5BoHZiK52x4ZVLJIJPwX69DePj213ZRspK0Is6wryrxwLmKJ
SAYb093g3+5ghW7YCqhmNgRVW5Q/A5VwLeDEblkj98Ji0RV6QJnInS1gOFIlK5k7
mSahLb142N6tFfXrVJfz38itS5z/r/lc8EyfP+ZPJ1dHWWgnIK403eCE0cQs5vPT
38iqm9zYaXYZ0/j9JO9NiaNJ0f/iYgg8DVMejdiH7AQNmjSPvYn2keW4IfSC1WWa
7PbzS6yZbWpENZNWfJ/LK8fEkv8U4mKPpx7HfDACU9+7RazPln16hE5bxC1l8O+Z
yl8XuVKtbU61xkpKSa/f6m+IkqbW0YIiwgfq8Pmw3y0Xd19K/5DD8NZL+bQrVOOF
azUThI5xQuvfgMe5eWWL+ZhwvBruJsIdCxlV/B2RAzmoW0/Vat9lwu8akig07VRT
ZbdVgWaeoTNFBsmkB0t9j5ataVgYLNjxpLh5Zd2NfCcm/Z65FkhvQd+0bFMf2R2R
DoFd5AXqVWzXSbgcYAIicN2KBcbGxc8jLX5qEw9JxnCPuDpA4ai5nrJb+b+7a9b7
206B27vC2M/aR95wKWnKZRH0hqrIgO0un8yQTnHLm9+Yp7ELg2+9SOdyVccBeEVH
SzyoJiS4r9stwZyDxxoCUdejMlxFKW5nGtdYBcIRbqBqa5dt2+LQSSHunt8XxSTQ
5JzQylqlJ2trMRu036IQyMdkGV5Dqc5iKMlPDL6vlcSDMEkoxf5D2Pov/rg7xNfQ
kZdvryLmwinkg+G1U/ZU0B6R02QE9HXqvzKaaqxxjlXzXmTdMQQ1v3M0dkGuuXCL
LeQmFTrTnLZhF+Yp3GY7duPGXBsueeiUKraCQAqct4o/vsI/kUEtHAiOEmAdHt5Q
xK/mCw14dhRPX2U9fqEz40FlZxpX5u4YjBxdBYN3ttujyiJzsGH2KUj4+lLr7Yx6
hkWXibx3d4hein7sjW6W8SCaA7h2uEr4A2uJwFLrZs8DGa96kHMjbCmd2Xjz+bSj
yip5OdNsDAYZk7CH8SmHZh6M/whE78h4gkCKTuQNLsq2aWfe4XSS1PheuwJ4L7Oj
KdG4LRaf9N/n578fBxqGOIdxgrNzdYoQ47GdrxIEmFV5UYVrg3rguWAgksCu2P2I
HngRdDVPA8SgFScZt8k/0N8yvTI+zc0H3wQs5w6OaZPMPhEQXGbQ16PKLIPSA25X
PkyiHIwlqJp5P92A/bpCxdwamd7HMeJP2uccCDcdv3qjmGxpsgOG+aWjzj70cdYV
4ZRwfEilXrkiuEf//w+pITulXK+G+B5h2zuAt7QMeIETmp9AypwScz9tZlBfqN6X
sOQd7Jv72WVWvStbdkeM9i68Eiz1Aw9Lrwmm0F/qHUxLk+ssuz4twG3VaqjCoCX1
FaFkhTRYB6hbXrAwPb6VrwSq3ZhwNko/elMR1alfWsQGaNp7R011njNCuirdPd9F
Hn/XrWxbi//T+oiqjjm0hcpBrdRdfeBGt48CZ84eXjb+2O3+d28FHN/QRee53QwQ
PNRhDChgJrOiJ1t5XpVHsAcJbswZ+YY5OYyOM3aPPum54FoGTaK+8u09Mrm1zdqI
fQQmvZT3jyz9/C+77nIn6BN13oDA3dC5ua06GqAkZ1vzuX+YGr6vJg5TmdPYGoge
56vxgBSF+ATFvOoX9TbnUw2wqbqHLE7A6jf2mmonefspXXDoKk27V5fQyuL+hj5t
Uq/yEhUNncRD5m4REwJPtPWEuBSJHCX0RFkcW9MggkRapxmXpYdvpp+c/iG7wkNx
cvqSZVpFjyNPyEcC7z6vKlI9EUBaytopIBV0XdD/ZYkHOsmRcnX8j85nvU4BVHVs
LHwYgEM+a54rPQRccwVtODYRuBrxSZFjlgK/UCP7uxjTAt0N3uD0/ZrKzoagWV/A
iYU5I86j0pSvCnB+Yn392p8cVFk2cUbHBRDn7HXAu1mKC+vYj1Bx8k9A7ll/1knx
/xm05Qo8TxYjpO3kKag+AWXZlbIr0RucEDf58a9arCODKn/qmssquW9XyGxu4xMM
S2gDYbRVPcpQM2qO10sVQLc3x6O0dLkwpeMoNXL7TnHTJKXxAeFwWFlPzr1zyaUL
gHQLDkA6zjbJONJOeMgR9IeHpq/DJtEWD4JUNjSk9js2lGcn74S7exNWZZ5rvycE
XdJkmcUtdeYCrV4+1vCIozVcnLHdf1LQYFV15ZgcJOkliJw/0/WhPfQDYeZUBPnb
HqiuhAUg3LiB9W/pQXFnmzp56zIAS2njUfwHcjrp2lY8ActPV/Z1lcmLrl3cj8hx
fbYyrEOrpyWiEAO/52hmq30Nl27cb2cDxGgYsF5EtCe2mHdvQ4MG7Adzx7DBIan7
m/jcDlcckFTBZcT6gDqRT8b/lXyMsD4iOwWQlpPPYQrHJ4CQxDuf05XatCCrZFJx
JThwzU4qH2AenIq2DG0zkC3VCn0GaUZNB8SMdE8ij04QgJ8AGa7UU107+n2Bd5YG
yZCIT6XcdBfLwM2hSK3Ldl653KgPPovrywLdIhlY/xv9PFMfef22leK1GDHY84YN
+tII8B6aAsR3eenoxHXsoCHbZqVVgOt8go8TkilhSyNrifJGG6IWNUiwxKZxzUkh
7HHk0fpcTN/jMFYhe3dqA1r268X4W/Xn2Ck8WQixm3obe/jaNqqQbSfLIej6dZc/
V78tU8n9lvorXVdYEvFsBppOKkTk8gqk+AMFZ036102x7JImq1YDMSKVO94WFPk9
xU8TI6QM2WYk9HenaZE/JC54ynVkMtCdgw8Bl7ihAmHtwbh6oiwJ/HzAU+yJNl6b
iIdVf0DvIbNu3fL1i3j6N+oa5orOKKtGeYXaw1C0LDos0Hev45+q/G+vcNtGEBJi
tMfjl3kwad2S+dxtepO+Gs97uesikpGe9wodGK0Jjgw3AKjVyBhLwv6A5QCZ9Ax/
rbpCF3IxGPZkSq1hgMDstnLNtpG+NEfv6jlVlW/d8jHJdXxExQpwyizwczooFNWp
B5BajN365czrK1pXO/7IzC5E51XDxIHUfxipqZ/17+2uVBXQDEkKQ+go1BcahEfv
+64dDMjx+CDtAg+3iT0MiMb8H0H++FmkeQ6jXFzUG3d6jAcJptEVfLj51yW1SihI
OfH3rTa4LkvobLOSicDeYBDj7M6PPhMYIHrlLb+9AtahsRjpAFLMIeFhB1oFhwlX
8iV7ARZciHVQrnmPvilME1IHvVpu0I6eSM60TFKYV+AK8xVuiWXp+iQzzmW4TUkJ
EvsVKv9Kp/nW2P8KqZgC4gCvIyUB1XJgy0jC4/K8St96e0gJz2ZDwK6Qvk8h3u4T
6ZX9Wbg6CHqbAzy3nhNGIsat0JiA8KvvqQJm7/JrwoQt5dB2bW1y3rNTEM12Z8lQ
XcT+dl90igssjG+wnNohlgX1kJmvXdvEf2Hv7A7j15zN6Gup3BmKymBTQpMAJ+wx
A2ZAf7Fm6rpbxQjv22l+yiGIUKRmqTJvR7uwaPhPuHl9uX2SRZQW8cd/Zu7fiaZG
VFOsUOwT+djQTai12XdGHkP9eGIwhD2OgiraIsJ+I+Qo5wm03BujMwUl+mi/gb7D
t9JECJNbbJ0kRK252zFwPcS0tcB0cJAx1h1vNWhcF2QRMKNKoQxlFm1KUabYwyeM
b0Adn8N0dsyFU3ecaV+9+boq5dsr4xupCHI4vtEEWAWdn8ExaBuTGAdTgkNMz96j
L/nIIaFE8ErxRFfKCKwnmWKnadbGODghV3K8MUECtuF3kGdZPyhUgEd6ccOyVuL/
fqi9wzfdSW+qYL0TXXnIF+3IhTj6/OSBtaPuGS8iEYEP0464yaLPLeG9pSp8l4Uc
vwlrzGFUMXLaYAYClCoffgMr8EsPwGN3hoqElKzbe326a1wNa3bMktAPsKD6w411
rwRjzbVBpztjJl96QRTmOyIscuV9JElEnr7sX/Y+hOQC9kQFIzno4HtvDGUZN5wz
qjqOoT3HfvaHr2a79lTvj0bHT/W+Ek4Uzirw3nIiwkMrDzxd7BK+gSMSHqhmnD/G
Dljqb3C4GE8sjNC5sqmwH4WXdd3jv0Z+PHaSccLoditr71FDFTcXo8TY042ukrz7
DBHXpCG/8DTgiTo8Ie3iv81IGKRu1vvRLR0JfSbq9DfuMvGTUVr+5WHl0OEckX4u
3EuRcgUrxbRAfB7OfS8OzmYs5xBraleuUXYbT6Rok2P0WXiCRKQEnHsVRNWnkf6R
7MtEFbRRBuSmYzMO8WHcVaVMJDyYOVDNEwv127a9w+9I0dfye6SzUOaNu+8jhRnX
9dQC9vHwFalH4DbG8Ug7PskxFJIzGtHr8y3xYroSEYuXezDsurC1vonMq9OSzOw8
stZQpQi+RgXskQv1zBGsWjK3mwQ2zHMYb70/kH+IRa+TWqhkLrNEacZtKlYM0G0E
gKyiSHAiHs5f8UCzCXGd4VZQh3iY8hMdnr/XZYbWZxLoLmGFmnz1ZtHivVOK4CgD
mlyXaTkuLcK2/N3zt9+eWH+wTGO9ywJRT8s2iCtoIbkh3IlUvRzjbWjnmKcl30lv
2+e7givAiAL0sobNuIPFPkYLGLUTZj+XFUi1ypEWcs5GCdl5UHeL23r8AxEYNzTF
pMmDKgec4nlIoB/ob2hic8R2Cwo2R9IzKNoHyhzvxYI/HnN9Nh+8wvGvfbdmWSmZ
NIEwjXEGUJHpJyopv1fUUxVL6E21hwh8fwR5T2LoxpLJ6BV+J0Fa5E9D5ydAFlpn
myQnWl/r7P7RDDfp4ZP+1HsbjK98AJWTsbiIB3nhpv7xUVdoULakdMbhzyM7dpwi
GDzNwo3cueEDy9tePW/5LzJQY5e3LaRySgDkuT/YvwTa1W2g6qe3VwHnvvzKJSFt
IZtB02X5A1vMNlH/UaEIeAxBrgRjFy5M6gtE35zG+ihvK7+YhM9N3S5SeLEkXdGS
m8YPAnwHlDoXTNcF7n6sbGBjuILwUTF/rGbhCGVJ8pHfnr/A/+jd4vlqzGE/zfGS
0XN+RaMvkKLk6QDZxq6NBQCdn/2kJVnCUtfjWruYP5xT8H3ecOoGoJK/FS6Ff3z5
XM3iqYRoXrsWFL1RgavWojjMtKeK1p7NmQR+TOqYjkEBCh1Oxu00Xg4yaazCJymS
dJZ4Mcp3vi3zD22QsEX8rMy08N1zvG8yx3Ai/bR47sYACLyJMSGtYXkGW18RQp6/
hkO0nwWSLrXm40QQUesLX5q7Xd90BEO7lw9jx6fX5Sr9WvWHhJjE9Z+B+t4iLPgS
lcNMcWb3t8e5iy4TsPE0IRTcjS6Ikg7m+O4M8KK34XFeRGDfhcAs+uUlkD/C06HO
nZCPzSLHzG2nQQNYrsegVEeCvDWhr0iydvqjRflKKwJydWwlb/g6XsE9JaFW/wNW
OZZKcXYWwaZQJS57UK13I13W572AR3N8gJLzIeFxX9TGyIaR+Lc0KFqv7yXRhGZs
r9m9DKmvjjuoY/iSiOkexb95ztSK4B50bll4FDsjbDp3sisl2A+xnw0bLm8fSSua
Kw38q3XWhEaZxabjwFJbXftYmvOnMIhqcr9uK/KLynTfZzpQHVMG9kpD8uSkg91b
Z0tEDLhCDU/bbpnoIDUyfTFnKCt5O5CZgLoyckr2cq687++iH4Pq1ITwuvcm6Fh1
Wex2wBrI4B/MfNENG2cHcvdHbJaIczuVpwIKVcCvjL9pbDYrosvh5lpycMNPzn40
px2rJRSvrsJeYhdSYEEN+oSI7cQcp5lpOIs0CtzWLEnSWTy7fBE60ssWXxiJXLG3
kkIeC1jT5uFjFX59LP0MlMN7F63xAXJbWQ66Fw2z7/rgGrIoubLmaLF5Xwga3mWT
PfZ+DOLTqHK4NFxNzJAeG+I9fjU9zpSPoydBX6drY/u16khrv21fRMJsvDFwLFig
b1dtbbuQdG+1uiYTUysFBecMCA19JiMtf/FKMd2Q1U5L67lMIjMFbgemFi4GPo42
I5/on7OqESG4ebCTuOvPlVz/IfxAUqp1YjOAl1uQ7L/EOiKhhnwecQApmNeD7h+1
XsbBZmb9RjyVH56x4EPsM5S1ZlkVGSU9d8rs9KRNAimFEPDlwSDlYc8jWuG+5ooB
BJtG+I+JuBLfKkeWs0ZhLzDRSQLIUQIXyRfWATKq50KELr1433bjW56wQam+x9/H
J175OgEhmh3dXnUtGLbUlhuBhQMd6kA02Sw9QJxQJKA+SFPmrywajDjw8ELj8nMJ
2PF9uKmiMVXNvJrWrjjwaQ0PlQ9rnyKO1yGfIMxF/MFyP8w4f5BDtDw3BS0EoODb
V5dGrcKDmKvjDlrAhHODYTJ9kvkoQXRJbo1NQUcHyBYylM7ToeI57eTuz0kPOIrS
7OomGfavwQOIPz2geaW+/hQDjcPtEQH3FeREN2mxI98A/XGLX03v3LqGf3mfSuYq
zTyubhtp5jDTw2oa6UXyvu4xVPGQQoiUDfe6EFO7Vs4VGWF8TOFybYrbWHwQwc46
0psCpLuozI6oA+KscZT2REkH60IBOWlp8ti/zQ7iqYG6GvU8MRJBISL7PcFbQMBB
LzGQBbJ3N9Y4uChDmUYXKoCp2DO8yOoPIBOSoCBH8z6zjOQHgF56SpSPB+QOLJ5p
PeoiNo58wSn74E2Zpt2wImpZ1gow4RzjnkqaMS0cWVnfjwCVotwKTaI7DW42c1Xr
F0Fmg4LKnVohGVMC/U2H+pPzQjv25yQLcZceaBh5JakGohEEkYLty1y8wQDx9dBU
KW5di1/g74I5jh4+0nr76lv/YCrlne/txT0wcF1ZJu1XxHRCMocdkHNppA6uALtU
pR6gRv5v+zcbWBIfOSz1DYFTLjxa0YwYnChlpVSXzG57Q1NPad64Bp3+TGbno9zb
t9lXQaQcHTKmdX+mFCOvK0go6D3cbN9SDYdOx6DAa8+qkQDab9JWEnS0/54riGzF
vusEx3WYzvp/D3nVSAL6eDafjF4vUIWhJu2d/UuYK8DtX813RBReGjxcp+2Cb5pz
WBf7HDBKfnZ7wYPn9WFf9HJF3zzIb/AUo9KY0btcMHj4Ncdfj53k45qt4Qm0KJa6
lGDhPx6zkD1ivQDZc1cUDZfn0HMj6+F0nmD+KxDrGngiCOvvMkuMCuqJlSwxh5vQ
99QeaVuXwJuCQ5yPTenX6E4lCzdOpgb4DDYwb/bo4gE64oqivyT/CTqGaxUKUsJc
THEaio4vq7ch0wZgAZeX2lpIlQpnAetOwNfr/5TiVaXS3r0wyaF9p6bkn4YY8Hfx
B1BFUocsvoQasLgQt+LtiKrcm/AvxT8+4n3q31PlzMeAfl78wsa1I3f8oPKRa5kL
9hcxw6X06eFsJA/nzJcZf0eE2IuFKiY9ZnvQ6Ns+Y1Hgmvg5nMB2tO+4X/XOTPLy
bUOE3evsuMx8P8rL6NdyxTszR1lFbxksnoLRl5VBEoj0IKx2s2yhpSftnE9j1AU6
VxP2QHMPZmtygF3cbWDVasnJqEe/AdAUPYwmcD9dSOw8NScHDv8u1RqfKe9ZGL2F
re8ioYcLJ6iOmguC8sC6n7v6XXlj1CxMN58tofUfusYCHKv7tdoWF08nf5Y+1S9/
tti0wYq6lT/iL5RPX/VtN8tqmF5LIpFXt0fIZ9zAgtBWeF4+RwXCuLG7RvXaDS3V
bpx6U3mbUJulppuH8Du9mTpEGd7arZYK87fEFyT2rtzWtNOrWe4tubXSl47GvoSP
Q02Cd4YWf9ulEbyhHweY+K6aY4k8PNkMd/aNBurowk3Kj/56t+PnW1aNyvpYzRQa
3w/SY0BvAQhEolr2EJDGJcnPISS4RIsD7P/rspmdAKZ8XL9SqspbXb1ala5KXlJt
qWiy/X7Liit/sKIBJhKM0fUu3n1ZVUAHN0dNYBHsKlnVQARae8XyDd9abkp9Bur7
pezNY/goF49zymXuPrQPhfB1gU1vp2/Cm2HPncHjJ968oDGfhE8FvdtvbzyGt5Ok
2H8OIidiqqaaTJuo6XmyUkZZ2EEmwIcxNzH4oTLAnEBOVjJcKF+yV0GF/1mc0y4Z
QRvYDSKSMOGDBGKAwewXOMRxxlbSRvDN8K1GnK4Nd8b3mF4BtF/iqrcg5u6KKugp
rY6wGzv/97iG1IyZSuR9nV+9LFhY1gpw+tLGXnMXhgWN8luC6C1otrC217AnmCje
lBqDmEjbpnxO+6mU3OOBwVGx4CN8cZybCgFA4QhFfegvKBMya6mGzdXXSTb8luwf
KmUYTgPvECEMBydY92mk2yPPxlG1BOQxROo91GlBp12evPalX74rSaBUTuwZNQwb
9keqI9dygBhHNzvpP2YpZPALA69rBy1b/TxCVATqj/i4LBNxRa/bvvmT5T+jfE5I
uZj13MqYgI2ym9kcOYWKA+E1wsYF8FowYH/jK0ZC6YeS6MeaJIA9O7zPsAccrSrq
iyTlRP28vCVUteZ8J4SzHTLfm/cXbF3U1jCC35ABvXaUdBMggqC1XAP3cloEaXPk
ULjds5kKQO8xZ6vRJ+r9LcAas2z+Dkm7n/8bbDJgbeWuGYhMYM6uq9XOktK6UpXZ
Y4hefdEK45GH8ay/pbwRBNmc58ghLC+/Z6/A3SA6beId1I13Mu75XzpAUOt12Chx
XgvcZgrfx2prB5/+NofrkCT5b2dBHM3hJyK/K+AnmHHXcvWDQBr/QR9gQHDASkDY
dUw6U4CENjaCKEIQneIEggv9NFjr8xbPYKxV7hejkyOFDcY4MwIc6DGjvrFuRCbk
gksBJy3nB0nouFC3+WaOedZH4aQ0256SBWqh0NfGki2Jgi6DqhsHNmQ3mQyCKlr3
KZG0Nuf7+rX7EA4iXZ/2Hf8ccgDRKqc1yyF4xc92s71y/ViHxQJylIZbpr90AypO
5dnh8YDPKIeLy9O1EYYe+uXcuqDMH9NxuHnr5wtEO3SkytDkKpivIqh3lToTTSoE
3a4IOS9O6kO8hOWcAqDOx1+gEU5FLtcnmkCZLq2hPAcvVj54cJgMsmNNOjwjZJJF
vySGTy79tCpLS0h2NtW2wMkUTxlCzTt9RrpFy6oWm1zjo62oIlYhFR9bWNMz9DfV
H7MmNp+5v3yinpFQeYiNfQRmTJozhbZPkb+V8/g2YC6uzEplllgOY1R7F3+whpqi
fW150CILFF5h7IOfns6tjjc5MeIQVseMtttqV+ilCuevuKvH7qvtaHjdg8kJkE6b
Gm4R0ncgje1SzaWnrLFHz0VVNyaOG79eHSuejWcH8hHHTwmbvXZUPCvhA1QhqBq5
QzZRgK6VJ9qtXdBpj31zvN2y8TSnawXb2i01K1q8VFSuZ4RX9xGRiJyPcTIWfECi
NSJ+3xo0BWyi4ohya0/i8hLwGT0kI2Pih+afUZjl1gvqNvRc7RYfW/w5Ah8l86Rf
r34hvuYzhHZXcWTdd8h0G3lHYzKw3RacKlHulG86yQqgELqlK8lbKQRhM+FVhG0e
Uyu0wCEEQbApsupk2X/8ouVKbLOVFnUgpnLYLF7RuyF94fCuchHuIvFkDeEE6RQW
BgOg3gSnx32SHlfi2iaf7DrU5YTt5B4IoF1M+enRQXQLgSNIkeBapXl8ZLEAJvk8
nYHHvQhcpCff1lCekKq+uX+f0C1I50fdlfWCijkhy3DW3rT855SjYlwLD/pFOhtu
uSUMuqGfUjisIPCLYpqaMSgg434um0533KmtfSf0w+nPgSRPggkRPvJEsI7U2aqC
q7mbU5zcf3rT6v9HJP76twWpGWqtTrSooK1Gl8l7HDOUDi1CTyYI8f7nDmsDrc8W
GUpWsuACtJQe9NG2brNvDV9QemzS5yLz8TMjbYKyB0OtBF3wZaf35GSioR/Yca3W
6fkU0j0dsXyFkpk2FfbuUOGxeBE668hFThD1YGAPiPYALYFU3snoXhK+yEI+avPe
iG7V5vcrKDdSM3WZiFIxhF87NoIa07C154mbC6PfVvYxovfKYqPw89k2quNMzGnW
HIBUV+YCDpkL+XsoMAlHhxm01R5a373Hj6KP2/izGrY3R5sMxiNXlikmcxIsIQ2o
Ro/GTv9EXHq3evGqleJ8j+d0FFTHZn9JAQCfE5oWv3SsXniW+w49qN9VVyQjYgTx
jhEyl5CWdM/DDJwqWrk67+bsD+QABXS6Mv7uxA2FNkg4CgDRZbi7fS+BY22H3Rn7
QbR0vIypFTDClv80GM6M7+icUZTqaVAnHX+Ys5sAH1nHFiM9OPgfRNYnzIzJF6Hb
aT0yFzJHxwP6/feiZcA6hzdFEr5E1Dk44mTXPhYwNM6z1Z/ciu+JqqrNWW6csBnh
HWm+5CzGCXYLpDrS6/L/a2ckEghMKCulPWobuVsAxMo8ppgqQGBq6cpPgU6IYsbO
eEmy0vBn3D0Q4tOIlm5v8vr4FXG9tEjJgeySXOF+Kc9ZbTRrgPkh7BnmYkI7sIhB
b3MMRyHPqbF5N7bDw5q8OL9iv36Nd5D7ttm4sSk8BfpV7wf3qUC8/t+yeJKGIER6
G/S2fJcicF1UXLKbTE6koal7xTB9J7gMFaPIaCLFGXsT48vVLSH8xZrj5p25vuGx
TdrwIRDgeRpxKWLx6HN3BSZ8xpVS5uBKosjUaSAANzaNzHzTifbfDoY7S6WMCgVc
c7IUayYTi7c3E6xia75taMdgOGpP9HN7aAb+jKVPcBOB+SN0QlTsTZSslEGlduFi
LmpVTH5+U1NMesAw36wksmWUkjHmdTDqcqGD7ov40ICi4ja3Vg/YzGRGlHJQCo6E
WOGfh3j+fvc8WNt2VgWtaRisqQ067VwIqAQgyeIBe63OBZE9/x1BHIi4s0u4BRNY
VY5qUhHUyJAO43NyDu/fBqmGOCLBQJBVvZ3giCS/R1XsWTWyV3ncqp61VQpPOi0r
pn95X3Cly3DcJh+/tiO8nWdGyAQ0NyIzzDAAErIZScsVJvLbihS30rjwVxXae7V7
Way6VcLoTRWgyEVFFwe7NNefHfJumceHmJC+Mj1tWLgfqaBJ1Jt2kANAZBlnPRSR
exF26y3VK30AbjyJ4d7y7m3mWzRSJJXfIVNUysFtPuxMgI/86JieUPS8IWQnothZ
n7ZE4x1NjYyXzMxNS2qvmTng6eo7xcKlc2Hzp2GPe3CmdqbqsPQvVUpX5cChjBJy
RyTU0crLQU1TlfMOEL/laTqGULK30v7CAfOPGZrrYKXfejX81wcg1YJs8DK7noG8
W/+GZ/R/IPo7JkGxwkTMJoTE6/Ifa7Cm7P3wd6JvdIaEQPIHofzBgttzJc93Us9+
TLv5obKrO18SZY6fRo4mf6hdFp8W49VTFexJ9POItC81JSWP0CC1NV3UT7l7fGbG
mR5rg97hfeBSRigNRWBpHA+hEfjTsOxk8Y2ALHZScdFotIyWQSj52E8/mS/KIZAR
1w+GTL19vzOx4+c8olYBnF74hveR17SyZg9QBP6kbKCaPm+RwHZFNg6cBFRhLiLM
eH0wWvU7qm0gjiGDd2DEiYH1H+3xMpaAF4+5veF252qkfcuKOrNy1d8+okW2t44L
sZwE73UrVqzZqcSkotncJisdS3nB1skTyosPUqeymsx8noQCLbrhLo7mK+8Aij5i
DhCM0BTRVIoqOAxqQiipCRyUhivjcmAAJatrhh2d12nSUzrcqId1QjJXbSRtDaCb
+YE7wReXbHlMtnu/CxFYuQr6Ja9ru/xHLitn5IQPBsuiUL3uDVKSxteKYaMIILJm
Pb+sc0HGI67eP7CccGzUUwY4Mtc9y0vB5oDLakHERup2Z/DCt1U7c5F/7QRU+qwD
vPp7qkzU5xARSWP9O8D5Ux1gYSaPHr6ekssN02eTPVP1+hLgYp+o2fXJGn2qsFkf
4UfR7E0U4kENFL+PstnO/Phrb/kZ5KSjY/YFsSKnjz/GOs/eAg9vheVmqtE6y3S2
TOXldrjVaJF9PXXDqhVBid4akCHV6G6lMDbKox3NZofDnaWcbbIFwDX3ZQC3xjWN
mblCj7Tu6eyxaqFkGyORaOjCnffvuicfykQlh287t/+r6Vxh0K/7kxdhTVPO7dcJ
OmypjJQfHNcK7vms9UuJ1CBjPohdQ8tBkIeRkC6itN53j2IvrASB8cVStYKQdMbb
gCqiGMkIl9nzMVjTqGlsXlreZUO9kdKtW6+Giwik5SMg+ltITW++vEL/PCiR13/4
duThiVRGp/tCos85OaPVZLQeCOlC0FZjEFdbvE9Zm4NOTQxvdnVhXgBxNEoQVyzs
0SD/Suss7fAgtkBWT6DkxGNK81SoGV41yjI+92jDsCMQj26XptAvm+YFOT8JM5Nq
x7LYM/4FrAXHDk7BsH6fkLRC8I+cx8HUw3VkhQhcN4pHfKE/4kATdFYPHoYp2qbq
Zui6aXp8ETND65koedlRzfOyGZVZBzxxt5J/80PuZwMSoRo8RzBLn5A2ekUYzmG7
8RJ8GOlcswncoMVz6ZmpDJI06LiLlondx1Dg9gXsZZc0Uz1z5we1gr4brhVJXV0f
OQcKjUgqIbcT0FIZkLp+MVwgMNlxHVLGNvMCbmYNygKfxJYrSMke7XUZ4fxqSzA/
bmm6bUCjUDJ+Zh7j57cLLi5sHOtGs7PGnSDak2+8ai3TfSJWlTpNI5v0x8bdQTEO
CdfHI7ZMCR76kxdw4iRPKGcqasxVDNWxfcquG7W/AzIyMY7oQApq2P02Oy0G7kiy
3U7hUY2xfKnE9eYCis71PFgC6TAhgKrZ7bWH3wbic0nZeRsVN0yzTk5RpDExduMN
eIvAaphrFrmckLXv+b2uKmjmHZ4mfrXVwvKkFrvlB6VaOiSCgkP5ydPUhCRIa6Eq
n0/CAXgyxKruaps36YmPCPo4A3lGZ0XnxQk08QpaENsOmfKe7vQf0Cl3cOnxaUnK
KbWJ63u/8bQvyreOzjHUiNDwceAQgr9yMUowrY6LvvFIbL+p2ftFiSyNvVlcoRw2
jM4meqmmUt+aJ6wOrHkDuD/vQb5319H5wo/19sNBDlI/VKba4xbPEq3QvK+oFPsX
L5yHrCncIMFZ3XzJKp2T3LRecys3bKJl1FLZVBxr1IVv31UprUsQvv6o30dIKRqd
3vLI981OcbeLYlpANbASAfuhfLWQqwC5qWR/BgqHEW+VuDKzJRFtuubjsoUja/7K
9+ArXuDjqfmVK7FsSz/OY6nWY+uPjC5e3OrLFy+Xweju79PmJUPhWyWwClkvajoj
Pb6qBWaHpKsZImVJy+EaU1rcPHUMnRQGlXn+lD2P/H3M0nLwKA+USt1S9eVrEyf8
UHKmKpqr1Q/qK3UpIeW65EWYz63eBkEJpbhPrdHWxaV7/wkrDcmM78SaBoX9l07A
U+F3K7Z9DPezsZebKnylhpUAK2rifpJmT9kjHsswWVxgFMDMGngD+FAYWQRtG/kY
aYcqjDZQ37Y2UN4KC3dl61IgTsFRKYMnE+B3BCKAUxPY+Nsy9Gbr8hRlDvX20lFs
FvQJuv+wzezZNNofC2lYCZReJ7N5C32vkmJ4KZpSr3eUr32tf4Dk18ryNFLMs1UA
3FTg9nU+HBEIdFiIS3bYeV+iUcb5/+QBrheYmjC4Qu2gzsDK6pfom1h+uQr/gqUs
yl4REyMbaUbh8AIjtpWdd1QOiBhT5c+jawW2luhSPaB+B3b3oZSC9xFNKeK7Ogx5
Ag2lCDkL+zIN5viz2Cym86T9hW7nYMIVkL0BJkfMANwZWI3R/T355gkwTtHQGbEg
x0cCzbQWxC3DRoDyLjlccadSji7Wn7cESbUajo7k//bACaA2hRZM8kTPYreXA37J
WDgHA0OqsSuJyb0WslQaOI1VUxptlM4HUG5DQ7VPpQRM9IWsjoEyJbAct3WLgzsm
yupfhhvHAIAIS6famcb8AfOcQGoBHvswx1hQiY91Y0GO8Q27Rmp/k2QVbPgHp+ZL
m6UgB7Qq2rHfyI3rEBL8WG0mWhSLrdeSwLbZaOzfxwiP9FuhwS79Yywt+LlOdJsx
O6fapuLLaIRkz1j/E1MM5JOqli4YwQvs4QPhujt1yzkqWDsc88u/5iW/LV0ooLlA
z5YTIr1h5POPjG2reQqeniPJXMx0+S1H8UVzHmE13CbB21jx4DTzp5w6jKjwUedW
gwcI2xkzq4BfqosWnQvO4ZeRzKCMVINIsA5IfJyE2UhM+KzSUC3WcBQJ1U4zUEzK
ve+pOSP3FVBTVKrwGoxEd6AeDn8xbSzk0P/SAitror1yD6lzSi3mGez5fHTBRVX0
b+nzO1dtcAhUmRO9Ju0AbQFos6waASOFGLBQvRhEHUI/7TwbPyEiwwPyJTUP4Ahk
VPl4M7/Bob1xfZ6Pbr45RDWRsfmULX/I7FSEvMUbf6TLDiwGjx9y8O/t7plwH878
0B8HP4A9ZuV+/u0kDT///TBrMQKs65zMwlJLh08cYtG1ZVBIIZAlPkhUq1jfrQdK
dTfRcdkuts6DE88doraRehjPcb3QXkK1mwcCbO1jQ9FUefr+MrZVnk43j4ea7iSS
vTKK2IPOHcaHwaCZS9jtT+ZsTOKD33yTIXvVKbmJvASGXHKbKxr1rlh0ZMB/CZ7c
xyMDQ4Aa2VY+jPM3h9DKR698tfLrpC5Eq5Re21b+y2XNK6AHXwyuvJIGYE9X2VVE
rMV4i18/YrvnyiqWFe3JdYiWsuFEJ2G4gA/fQR7SQOfrAPYOqi3je9LwJMzlkelC
MN+r8+yprneIgsrPY1u0lkYW6Q3ivIIAdJfUWFBnA05ou5Bazsj5I986180zkHVE
biZwfItRSXwl+ehR7Gb3jhinXzgUiE3+RU8G1TuNC9ZZq34YT82kJW1jufN5vz0x
tXIDbIoJVnnGnyrH7kdNmNRO8Kb4xs/tL74xggivqmQ8Ldh6lvPqQ4tupVcjYETE
cYOriUsIPsVuhtAKvQKpkfsBklHKJ81uu0DpRhsa1jzwjcM5FE0dh4yC3xi/K+KI
M3KR8olH9eatoAGS4h3j7IXcepMwkJDS/TMvj6TL/Kc6mm0nwLNsEOh9wtaxOc3Q
u6QHKBf4yI9DSO9yOM8Aw8lWd4rq+DTsaY7GUJiT7dQ/GX5X4qtLINZt+hIDtJS6
l/InVpVP71QhJuavu/vlfwB5BprWunlj80nWy7JUwOM+2d+aRj2Ku7tMal2dxFZb
9c8qeZO6bMPQLD4qe8de1GA9GTAkQZLl7sC0FK/SgQ9hlr6vz8lVJAsrNhWnq5Re
VeLXIKC6R3PP5kVH4EXsbv2m+1IlWhFymkC8ajk7Yq+I2m8uCii7DMzvGmWxXhlv
IzA0lxGr1IZwgelPXgja6Q4ubzZfneC0AlVWBoKWsteGHnpOWyh5sBKxc5ZR+S//
KvnaQjUWju0QOPk6QCqex3kyl8kkh7rOqzSgxVKgnx28T1hZCHZfjnGKOn1+rs4I
Nu71Bpi/XQ9YaDa4IaBQJNtWJ1H8UKjBEaChVH/qQXs+JZtQN4uNhzSvhf6tXZBk
42z2Hvo29l9311lLMRf5ym5a8POgVHdSCkCwSNvXk9992eWDqSe8KnTMUYuZEZQv
58+Ae0LKAfGan2EZoR+TOdcrbENI5COm3Kwjjf7pDptOaVfz+osc51BXTfSWHq6O
8lSRkuRMzQbPv0mMfxIefVIt9K/xwOzLIwqVYkDWuzsQ+5klrMVBkiNwu6Dv3fPG
IFRfEGH4NpkzqALsslP9K4YQXLtpQn88Hj+hRz1Mbeydjc2i87bTdsw4B8XfCRie
9Tcx3tqk0YyELKruZ/khERSaAM1DREYhkXmJRbKlukKx35oBv5aQRNNGPVdPJIPv
olvvfLnfbdOYY0SHs1vKMCKU/uOP/AHNDIdwIswT1N1Klq8b6UALG4Ll+P3vTciO
CKXwnZhKnAC710rr08CuAdLp9K4mhkOu8Lipg7NX8EgXwyfJaBgFpyctqplEf9Ys
Ux5gNuC6oSczDKSBEa0zrFV8bfM8oXPDd3Y+tuhrc3KnIDtIaSWbWXyS2Xm8Ombi
mXlknRH8MVyfNqd8BhIieZBrcCtutixGSZpiqoPnn9l66pmssjxHtpS94fYE3/MJ
w1LgkK6x2eQvNkNM+y4A9aqI1dKNlKmaa9LBZICrY1EHREOxBVPoNkHDObsbBu97
xRZ1Gzi6ffCHck005WQdfT7akjSLbtLt36SXmFF5jdtfCnuNLXYg2dE+dgsxNmYR
K4reo/6qnfPZ5ObjjwBx8GH0a+4Tsa19pPuknPhJjHmEy9iFCigSZ/P1oO9T17Y+
vJUncIl4XSPaGw6q5eFU0XFzOAzpIuOPiUcMElWsZatX1Uw+dR+9M+2GK0iLc6P3
9AzlwLFGrUUL06OrP0gwUVrmsQgnZipHX79DH3k/ZRzPrPXkweR+xC3kv/A9UKIR
vMzF023tRfKSN81gzRIh9ex0ZHvfgNzpFCyNrAtah5jNDeccCo2jOyr5shBdCNie
GKJ/7Uq5h19ujQzNehT3hjMXRCCLw6uqEkHnYqJ0RJqSusmO0dbGmeZiBLCA3Ti1
5r8jvIrmX5QML1V8RBxo/v7k5/uTNAKjJRS2i6muevmFE+9Qwn6+1LqYPVMJa32F
kQ5lQQkr6dmoVe0k0ABJ+ESVWcynuUFNUItv3rteNK8YDYtlXDvD9BW1ilWbWBf1
XG2dEboU+MqIZ+oRj3r9l+VMXKtdWsvf74HgvX34dO3g2TPGnvb7wGS9JZr2wwLI
fAnBAAVkT+h77gJUQizaF4kw425/Y7gEacj0HPv4HO2i0qoEag5OlfJmSEQLT4ZL
NhD9ROpRXN06IOgt1nukED/UJxp1AsBjAEaXABQx02nxbGWSAJIAeGDWqaiJe1/E
y+DPKtmjXmzs6v8+Ykf6+5+gZUFONEI/+W1974T/YlmrMvudDaHRD/fCB6ESotvT
LPJOInwWIwiWKLHLEmIc3kOomrPXZU0S+b9Mtbs+fwJGPzZgntT1ik9x94a4IQ+T
0gFriVqSBFHJsNml1Ix/Qv3EB4d+GoPL7Rciap4spJ/ao9cqPUmHGTELeDvQU+61
VTvuKvEXwXYnDS6B1Y0JZupa4ojS0eTzurwrcDuDn0yI5uUy5fm33ngdPJZBxg37
EiFBEruVqSGwEZT+aR8nfznDM+G7/cIqMqzNaWm/61CpjU3/rYD/Avn1WIZjWfUU
8FEEbfrACQsGH2AdAEUp2E1ei3A4SHXeehJc76hvbq0zo3SZWrCs9E8yfiHeiPKj
kqBrcMfhYywrR9N3pUMtdeBmdUci7YyqjfYTybCKHPm084ixR4G93q9yKTQjd9Ft
UyAAxL/EtLnuzXUzw2H9sieDvUNRuT0/WMoHs3ayCDpMUs1SjwkYt7JaKu2T6ojF
q2qrnbrkErAjTd9pz5L6TTJz+0vSxm3UBtJ81BIVu29zI/pryzyZ0Sy+CaIC26nG
w/tA0Et/IjZJrTSNG9N5nU+Txs4Ia3WuXsSSgfDDAO+6YILWStk4Cr7CjZIKAA4j
fl9dd+VOJYeajfhDsvsCng9KRo6mYEDQKatv2DgK273YzSjlJ1BbqZZ6q3BxqxdF
y7FRSan/3tfFTK0JSFMwqwS+St6HLCiYafUsIGSU45QWQSfE3/VlXoQkJ79QJuPu
CvsSyAIV7v2w1X/G8k8CpOrYnuweuCRb5ftTdv7dk367PJPUG01TnFadsiyl8nig
e20WGQZuCfgD84MmUO33+LGOTFiwTwc6ndak+gzf63hiA3PjUWboVI7gkPM097pB
ttwirVmN/r7qrBL3XHqjyeYdrBUYAVYRE639Y8FeBXYIBjgOEcvRP6aJQ/b5HGje
TFGRWX9Wx3o+WXw26nmmRr1veOrUwjAemU4/+f2RsxB4sHLYfZv25kW0qzZCjH+Q
SH6uj9bctQ0pjc7FPcWrMsN+Cfm9kiEFODrhfg2s58jG1jhJB2k/kOydGnHcVfdy
4R77cgN8IVk9RiXjTTPNQVZAD6kxNbzq3MymeXcY0yZ637UMUsG5iWS7kDvTgH0R
k66M7T/Ra15UtUy9lO4Hwd5DYw0cGOaepbm7101BYD/qOJ/6pPf5LDokvPYG3PzE
YIiUBP758GBxEzIJaUMnJd3doWhhk8faisXWRw+Ua7CUUS7+GRBk4hDuEPX4KjhW
fGzOq8Y8NnCYGNkwrgswFFmSMi+/s9oKr6tFuUuc2EbC6DGNigzTz447pvJ0hIKJ
XjgkuAUux9b2JoGzknm3B12/ZNC//wiuux0hyNlzkuXzyhOowVfUJcjbvosKWL//
Uy6CgHt3kM36EPZ2Lzzl+ScX1EFdQQc5A9TMEmDXNCFB4E6YocO6NFBJzeLvtWvm
gqxR7GBzLVedAqWn5g+73CbpxGRtXCfMUzkjW6wJy+fKVHyKGLH4mzAuy3pQ4Gpn
SnftJJlBhxgV1L3IYAkWYVq2n1Cc5N/86CyUI17KruQ+CX9zFg1GbKKXRnLWpJ/U
M8XNw/jGaNmPIA6eOQ1CTrjzMDkF1/qeucCFOpABMNgLFEGyR1hxekpdW5dEblaL
t6hMlrapcSy6juOHgjGABXaxRzX0ieJPAGVhxJr5CNKggmjYpuGGEXvQk/+zPgj0
CKBjLHboJ+3IFL2BVgf3o8NlT55fS9cKlJXF2xpyImiNcwPuHHuZbDVD0U8z2X+d
5pXo3h0fPHy3TiQYP1/OgTo1YdoMKLRqSk4jJ5bsvXsugE1SftRKgOe5u86U2qtf
++WsLjoS3pwjszN7a0Uih4GgEsnDlFNHq0WvXm0FRO1g6oyEqt2SmGtiKoz9YGDV
iV5k0j1j+xYCi4T98gWCExNu/XwchMaE2d+1JwqQDXEU5NTZ/F2WuD3CNTmRRcIa
3KPzmB21GvCxne55Ob0xkGEcsh7h7RlzVyv/AqiutQpoxf3cfZNkC1ja09VT01gW
1PprrrBq66NvoOBDkkCLvEg81LLaaRkVpw7JIa1MrIIh+FBfDtBPGVwlXnZgg6G5
OTOtFhRtWzSCwmwUd3MqYbKh/dgvL7e1riLaLhEmY4YVHb3VvtShssJevk59h6h+
+Jy4jpNJYa0f00aGFBcE9oh4oLrJWtfxOIiax+mVmi+RDfqL5+MXjBgrTQEtteEb
hAKRAiM71qEwsiR1J83iHT2jCLOea+sQgNkRuajluzag9qNN1g2wqNqW0GUVBTsY
obCZ1remGZMDY6swZcGZFMvrpmYsdGhneGxzILJ74R3FeQ0JfpSdCpPMW2REk9R5
ZtJTRQT+pXIeJDxrFQu9y7DSs+XnAwyz+zHskFuLJC93JNXnh3TGeeEjMa5IkWZV
v6ShS82OAdQkC6mxuAggspaIAJDUhuyOrskhNVo3qFiN27UPSdHVVLkN8HgNIiw2
SyIn1trWy3Y2AOVXNpzuvOUv6Drps3suTTDFTQHKo/hqRzo8h9ZnibO0VIf54/Bp
Jc8qXt9Ap5ej8y8cr5afmJHUqdB9Rv+j/N7lP3yhsmewJhSx+D9sX9q+InZbmTFs
izq5tSoJbbcQhQnp/zCymrlqP2w0aHOnlzRLlDr/XF73JD0sNJeKq4QF1o/XczCR
yvkV5Eue5XcARGz1Vse7mA1on8rP2dZwXkoC/AjiNDE4ZbfejSSrU8nm+z1zsXRS
yWM+uknHqNALipLPEmPNVhJBKVwmnkhgOQV3o2LGFE0TiIwKriliI346fR+m8e18
2/aK9V4YZfwv9MZp4BilmS4RZJRDcdQErQHu5gtGhkzcmkbszd49KMPaXlFiKGpj
Op3pnj/1faBqVHOzQ8/GOTvgf6uOyuUq4MMqgOXYsU3nuaKcRDsJcLnwISLrjrIS
64JDdI5YVLJ7w12TPgKkCaZNVTQW9X1RnZt5ZsCBJDzNXke0Bp1LZ33n9V0+t43l
TTe3FWmKry8ALlmeFTIBApO2LXgnJelbrmp8yvRAr8sjSJYAaB/OmUvMg9oy3AMZ
4ejyHRySNoQBtmSq8erSMIFDmvr8BUKlJtn3ycy2tiLdarnW0LejLxoDOBeiC5JP
ic6BjoGpQUwuOn87mz6Wc4ubmDK+Vi32MFeJFOn6m1p+oCjUzoxYwyNzMymFv6bl
33K9oGnWexMDn2mkal4O4mFGWPqtHUR123ysra3RzICHVcvddwsDcZhzJQIHVGjA
JH5qr5MrNWscQbydQtS/80zPUVrcYfXucxZLCyVXLykZqlE9xeUo0FMYyyuGAC3K
O51TbXXHBImVIQ8csrQavZnZbvnhhpCBcAUkMhnHkuX9nOQVevrUKgabkrUUH+Rn
dIk3bjhRXLuCNgi/QZnlimufQQJe5XRgFTROHRR8PDUtOhMQNbSTMnVSuA/ZZJ/7
IFrhDlN6Ew2G75NSGc0JeEdhSGcweTtxtYzJcn2xxHFjixNug7KDFCsi5i+SPSwk
RG5WvArGQgnV3c2QDLQWK3/TwiWd4lc3BANTOa9asKc50h7yc8Jz5+diImBQOTxX
V79rxW+i+XpHigF8SH/Tc+2NMagDF5tEtP2osMAFg9gHe5GpqqwUyaSezxPGMJhu
TIb7bQq8E2zdfjqohbm4J+rKZKjwTCDq32xAVmGoOBw/dyNOAiATfOfp+UKghAh4
wQiLEbP8X0Rb9tsKlxRufihGuQ1iaXe183G1dmkd4nKSumDvXeMlnzWkd89xsDcz
omDslOM4vwTjQ+UR+WEGWcGVXa4vwVs5Ya0RED8n45pdbirW3ytNfaUX1bhNImth
AQEoOpcymG4fRjnzJW+tI6Qj2aAOjkgetLs/9TWQHN9Who0hngRxngikK68+K26n
MMxTHYuAk4xMRzaiODyFcE+53r/QFuFiKPU25fSwlPfZGPnGC8/MCR9w7cVG3Sv2
FdPpBsZkCwTjc/H3FxZPuUr7vrkdXiZalgTYNf/RrKG/RupRtt/Yg/j1QyJToC1j
/Daey3rNqCLCnBmLVY10xTmzf6MIuByh7MEdTYaA1HsyedLAAWZlUiKqselLKjbG
hPn5aH7Iv7dJyT8EvpSUklTu1tO92GMRAygFO6A9TXc5RvpvVWzPzHnJeAg6fDhG
0MtHRoW05HSeNR9G8gHlvuqdczjNvNosRMs52TEiW7Tuje0RQqM3Rjxl0hdu4lSu
DVjkt1C5y+YnaKea4KvTzsO+0ksKgCybZS84YqBvko2xdC53xN0ya0nuQp6fHP4A
BrSWbEKHxvgW4/5F244l1BtUkJcXLjmeMzJ/ZSFxV0hDP4ZlG1IW5lcWXJwRJweJ
6IqxegoQZP0uG2LpE+EXpeWGcI27tCVK6H7aLAbgxKIYeveFVF5nf7otdwTSFbvm
o6hLZmcTMZWd34DhgZ6zr8jLQk5zlbwAGnNwCa14TGaWZi5dVjyOufPO/ZnlaePS
odKKI8yJXzHcf1YMD4lHQxYXsQNKEONukD8t/QxYLUbmiI7+EZMM420Uds83Dlxf
yGa7itZ7ciRmF6+dcB4XYV+bBDb6xNr8DsuJu1VeQ3wQdwqhIauNvEXvpoebvtU4
JycRmHivCdSob95jm5pxaKm6NV97kTpbehH7vDlluPoWjqf5UWxHQEh6o7/vL4ER
gNCM3cJbZZ0DnhEKwvmtWx0t00PvWejCK2ucb3Wx6IjrW9w7XBGlZm+9KeeD6o+5
iMg5O80Qbm0cfdybgpJVZdQ1YyVGm0R1CrHndKlEZuLOLMU7ZXBHfIRFlvByZ+hX
VzVeyRw5hbU7cqZuhh+8pxGlftW7NLaEmyN4A4pStbuOz2Fu817+Z6JPtzXwi8sc
0mv/wU+j2/HM+CUrNodjM20lQKMfZk7cIhBVUkClESXeAS7VPBPPHk9VB9AjUDDH
xc4+h1c8ZssI6vPdgaMbydUA3i6bQe3HuNsaQ6I/RAi0vPwGN5I7I/f+EwstiyW9
3c4m2crOCfFj9p5Tsmof6sb/+qzGeiPNlVYLw9S0gEwVe7KJRgv0E5/y1zGTP/th
9NbmVLMjlxX0rVaCYMvuLHZR93HCbYNr8A7XNipeAefAiAFTGWJ+j+jdfmUHCOBJ
PhJUyHKIlp/vrBleRL5cHFbYEeGlitRak3LYQvn1A6pOoBzP/ByJpayI+SAy0x9I
1M0vbr4+GuIfUMTUCxePtWL3JBrfuB2j83gqLlA/ghkbcvkbHdE7WSRlX/xGm0yc
L9SndD21SJ0L9uNFomCchhO7tW09XPsQVWc7PHYMz6oDq9N+c/KARZmnNhpwg5kP
ywbwAQCLwTsUib4ptnx7npQEUuXWSSGmvoLXoi9HqjLDOtJRJv2WWkaq0bYDimci
OQ/yx0p17dIcGVo9w+WLrD2BVySQSLszItfp2Znf1uWvmnTLre2FVs+xaBswUvWv
IF31uj1fPh7+XIhKjfrfZJeoOY7EBT/9wwE/EkoujwL6HPFwaaqckBUVlyGbBXCh
pjbVJ0jnFEETG39jNjIe+HAN3CI2og5zoxCoLz+OLYuJ2bEfPNIsZsSc+DjwiszW
96G6auYbie26PjcPlTHYDWgS5U0uspPR9lD6cjwq2L3bo1ZLjCSGRzr+EWmuyve1
wrfmXkqRY69F+bYBzDX8N9iidX5Sln1K03ac5C535zhvxnbd6d1I7wihwYcrYZ5S
6liz/ebVltGTqAc5Uy2b+lgbyFuoQ2fFw+/oiAwsHbh7vnreSC93SipsDYlNNQom
E6519n9nM08pOBvVDByoHsV6M6Yzd1XmJHJikOvaZyh1yFEykU6luU+mIvURZcix
7wZ3Llec+Wynwga/gwe1EWA02+VZJU1kjkDmMxMAAp0CtSfT5nTT4Z9eNIyzJ0z+
NnrxjBeuZ43MKRrk6r3Th3L6GvPB6ASYu8P113CVCb0zlw+HIFCJVJ6ODi4gtx41
TdtC1H6zw9YPx5yVtJ0OelDIrLfL6ndyTXom70v0oSlO0+YCIw2SB3IC/wyvT3k0
2Hpy/IceXo3qFkFIQnEEwfRtyXmNK0ZuI/Ab+XgEYB6bIBNQCs0kFmz9blZAEPsk
vZJkdlGhE1UprrpZUPvH9GjfW2o85iCieHNvhZACFvF5j9/q07I2iBFy72o91jJn
1a90mLbA6l5exPOXJUe48c/xFsav2sNLRxuHpWN6rSsIZvhF4dxnGMakoA2vBHe0
8cWmTQdRjeVcJVC7NKLlN8G23wgVmvAKRmgoFCikvMx34d4EHe7sVffU0bbvOCkY
pqn38tuEII/IVZb+nMyYoolxBaYAd6iGlsnGAmzfPXl1u5aop/3y3HQBawrTuK24
MfcOdCeqOuA4XKslfrcKj+wKr9RyosCCpfxncvs8PG+zKE0wwDdSceOFgG2BtXrN
VPrIc7v3nAUC+yZMxT3b7EiIU6lS7+Yxexx9PTyvXVAqtGyEy3O9U5kw0FAqEof5
MmjfGZ0CznVwRwdr+D1HLfe86FHlMv3uqw2FnLjArS5/2IMok0vZSrjxb1YrYOfG
oCWDpoie3qsIV2+YgpOEmOu1/omjIx7kzVmIWPsJw1FuP9pLHxXC5B3BsoO6X5IL
X1hbsfEoWhObkqGoNZ/NyVqdKrWCZpb36rZEqp6S/bwtSAIKCrHhOesOHO5MHvAD
y+NYgypaYX8L0d3U+yC8JV2I5T5IFogFEz8vRVVrhryu6NTfYP0LZzdItwOlPh44
c1RGSZWmcBKwkdXHf1NE+8uPs4RyZs9BPdq5dljAyuxGsSQrf2xkLML+EV/c5Yif
A0C2dpE1hDXCW7MU7rQru1HsMmCOGRZhlk6NsBWj9O1VqMVnIeH85Xxp0LoK3IGr
TsCyJKlzTy4E9TwHGTmY6ZsF++WjDtKbaKoDZ+zNfxr2wvAhZSgmOpWfqK1Jl8bg
oc+VEieVQ+eUxzgyZBYfj2aU6LkSaEMpuppC0u5dvwr/sxjC0a2Kj1T47yljpV5z
0RwO4V7lcj6Md/5P1t7TIf4Xa3FYOCs2Lurgcn7VJJcBHGC5QtzChC+wm24QfGHa
hKjEhIuYJxu44F6LqDfMOcSJntzAvAqQYPxOc1SMQomJsRGnDH3D8jcgBrE+AlGG
oqiWf9CL4ieC2XV1j/3QmRxbZPD5iCCYrm+3/zVBSwPLnE6udYYpGspzkxrWDkAG
pxrl4lDciBN0eB2BD0Q8K4WP3Gojf+KDel989xxjaYlCJdqejvn5UoG+f43VmF1O
iHRpnzEBCxrM8H5+ve8nc/bIFAK/ptBw3Unhkh7EWqapgGfuS7QO83rG8IPXcpbj
Kw3KQ5xD+cOVOy95+Os4F9/Ndx/RjF39E4Vwka8Qr5GX2CY2EYz/NWPjr1pxKuED
/+Dld6L4Z5wWZAc9jN0LkSdJfexjNEJOLQaT8TACkOLFz2lUB3NY9SVbxz92ha4M
0YqjB7ZnPUJflgMHcyzpz/96swDRKMUB6ejrwmnzdv/VuxD8Xf9I2GmZepIuD2wp
/Hk16JGzxfTRHVZAttL1GpqQ9ZJ4+qmbLjkg5IO2mABnLJgpJiOomBG+l02NZG96
Jpfd/tCL/mEOq+vCscYLLO983GE2y780m3pzm11/C6oq7UyQC8J9CMTgN8khC8Fo
+XRQ0KarFjTAXyXLwQrcmFJycfHtNZCfwmaioDaRiQsxh6uQ3J4RSc3LV9kM6yDv
X35UxodHHD0LacvVTGmFbrGCE1oY4x73mYbzPYckCA5fC4ksxjSu69ocnSzFhXow
Gzza4llH42Yni/Md4xWQ9/H1EElhB2nmZADuJEOUgWNXRd0rCH5cCdEZ0NySZruK
4//Heb7caPyeFeFivwaBowL7o4UJjVBhwZIVeovo+bkLZUoEesED7PymwG5a+BQg
3ha+tto+1ToYmieawZvkMCajV0fX+MhpDA7nwi2zGbTfLGKIEr+xtN6EZMZ8U1W4
lKHR0gq4G3QsEIgr37DYkZ9UWQ1hzbtYBc5OF2DjQc4jXTiQPu5AGbHpvSzX1/QJ
ydk+CJbWwaXnsGQHCmbjR9H94brhh7Qaq94kX7KxrxlfgJyxD4hjOfncpT/Vcnaa
vNWuQDr9dtN+mTlZ7I72T3CkkzBKI6+N1ahFkJ4wulVJKW20uIXb4DNNxGuNSUEw
ksjhZwXqLysuLh2uaSDI5ymrmrix+cSCU2qRs/fcrD8bhbtFhxICYKb9CIi5EY+C
UK1dhds9Lpr0Pq3QKryEOo6S5dXO/tfGw/g2PRjZfddZiMeLeu/gY9wqwKTFZEs/
kTXLBTLMKYonb2ll9AIJ1dDjdxicIpljvxWUGNaGtUM/ZVRZ/3toxvpy2XXtW2hm
Xe/lu0ghxFGnoXMhdxOSl0qTaj76tM8NYfV3npXGAbOxKelfKlTWU5Puy+ubIGmK
jZQ8T0xMR30YtBv03S8vbwm1Pw5FHl7DKO3+njzurMWci1tRCv0mSoiZxWH6EvVn
D3+8x5iRVg+PQQH7X8J7vRvDcemJuhvVQdGh3rM/OmJm47+Q9SPq2zcbMHSO1X55
ssMCv0OSEFvJvDCxYhPy92v1b1vqbzFju+tNh+8gXAtXhCJ61sTLBOrJWGmmRkHh
Dm2OlszPD4V9ttMgXHCPKN8VXGvCqUpxU/VUwjdNykL1H5IEW6n8GPX30xDhKmTV
1xaYNiHTYAI0q75tYAEJxr3qRfwwfD7BVYigR7HQk6j6FPOWLUsVScFMYmWntF09
dS9DWaRMVnbZqkS5jiNJEMrANriV0k1htGuZVjlPgp1irHWf+hxxgFOwEG3qGGf1
ZiOjSneJ628enxgHIzpoW3UmYEJrglfQ2PF3vfSd71QXZk2wzOBFq6J2JPVBqTo4
HqYaRt2rCwxLqm4+KiFQQvzYAEv41E2tu7sUaWBpc/OU70MIi1nhyuxPkdaJjzSv
Mn8ijJhtKuYylLpncW4JlAN1+lru2K1r5nBAzafu//D5zTfvwE00Ehoz0zTMCVYO
x1sqAYXiHcommzT8FNW2YzzX/MQkkTGuFEIqIjKgKfUPmeCzKuHP/cEnRBdC5Uak
BdY0AEoHaWBeHguSOgr57d2jN9Jte4PVlJ5/Bxs7eB7GD2H3G+XP/qQEm6cIKkU2
s2Qd/EQDYz4G2WRpDrDpCPuX0OIqOF8ARAH3O+EimJJ3rrTvZ6bsl+WuQyunr/8+
Ub6MQwhtD5i8T6LC7FlNhLy3+vkgvDej9QewgTZVLsh2RPuf/ueg/qO/OEvQc2L6
t+qqnkDYePl5bHaio1voi8Penob8SdNNI2LsFVgr82eyEVpgrvqJJ5EcQRRAK4cF
dU9brawXyqmMkGDdYsfpo6lK0GjnBh5Wiv9ooAuDbizMFiS9b7VCmeDSKSgibF1t
IPZ7oNMsR2pit9xiZTxuzW3lFv/R+wRVaSxCu3AwiqaRpZ0TipUa9VQPHkHyrsH+
VsduWCopXfxW7gcEwOfBQZB+F30fbDMvx6bWyiEUZkWX+XO0j3DfxM9JmBPdj2Wg
+UlWS9zWA3E3aXIA1PhKLEQaJrcdElGysXbq54KraKZinkDK7XXk/Zu8DzaxBAt1
9blTvwMrUIsO6q5NLq1OgvQkIm8HiWCJgGdDZQ6Q+1o2SLFKvi9Gytk02qd3nRBf
R+hqDqnLBRNja+9Z8gG7FE7fi2WpUZMBEBH9posyS/eBDFt6O1zEO9tN+Db4soSn
FB+U5aSoaAAqHBgNSVaC+THiW6F/3EORH6l+aPE1tDlz0tfXsc7FZNnTVeHkwBP+
4SOrqC3dNSwSOzjJ11ljb/7qwwIdw1q72hxPiZ+n0H7z1CmfZb/7L8Qj/Ak6La3s
3ZcA6H73hwaHHmrYk7gfPiPLxIRDeIhgV/aq3tOBpRWCelTsQFCB4laK5RFOaeWK
bIvoYG+ZAqfItRyeElSa5qlMhhXSUc3XzGiTMkYx/NAK/TYSsH2d9LX5tP/Torl0
IhZhuifqpfUVLwmvQwMXRvO+7TRfvxN/UXYyh6Qb8WdN77DSeiv34Nc9XjowYlEU
Sz8IzEWG8oGcz0z9YYNkaZYXHDUe7c3FdIJHsR/Blug/ftJUTaTbShsHELgKHWlf
amtdgT1A7P7xcz66OF1mkMfweOSP6PgPkv1LB5x6tOBLxKYeKjJesV6mHrBKLF0/
dxXSpCKchQyjPUH1XGaBzY8RoIwjSnEz0CuxrcVyP1XlyetMYgnfWF3xk/EZX2lV
R1+EyBoHcIznGrcEcsm7Y5g1PrMlATE5aBWRZpcWPkAUuiLxfhMd974hClQtG6s6
+lHYU7tgHDRkwhoDKeS1dim/Dl86O9zwdDubt6rkUOt5HmXdy2ILsQH4GwR4AkmI
CoAWERcLE0fSuuvIfxRl4O3g1ab085AaZxYqaCigq4j7dd8XEWjcOzoeW3o73Vys
RwFRL6tLxSTappJv86D0+Z6bsFtreB22wX3jFFQUa7nuyjp1rYG4wtO14jeUkvQ0
tvoV0Mwx8Qq7tGNl8HiyLnAv0Vw2FJ9Dmx+KLlDoYLYL5hc/36KpnGtTAJUMQIL+
ASv2oWskYWEW/mUYVDygL9RI0NHfD3E49Hcmv1JmzRqLHssVx8ogRDM9+3WVIDHX
6CwR6VDOq2LkcnZdA7IA0CxMEJ4xmNpNXIJ0SDRNgVZewYbOwj1/aag3oepN4CAo
lLschirhr+xPB7dHNHmmN6cdYLurwcaUHNiVfoByO790FPzAUj/DJeSH31S7esA4
rDAOU2j9fk4JhEHjC8D4XG/OnfjzPLTqIrkDwBVPVx0vgYJS21ikIHkzwg5Kb2sm
u+kY+AMESKBpjrlVIIJhe4SwN83HCr4O17BQ7INf4QRZ8JZG/ZdeZA7tyYFlzRL0
WTH8WB31fJuSw7hbmk2Bf20Y1dD+piFy36sALn6H0iXdmrguqcqX01KVZ2fbWSak
2lsqwhw8N7tOCBsXQ5dcmxVQK6riMR8Lcz5RIhoHgK441vM10+3pdb+BIvBfrnUL
IeeiWhXpiwTSFmAVVj5kh8vxm/fDMyRfpKCvF1eBKY/YI+iyXQuFNE4F4m4e2mOg
eiedhQHHa+bECJsPVvmxIxca7EmKcykNx7gp7CD6SegBxsfEhgC+3VVt97fxAKc7
D0BFovXD5So1sG1zUNSIivBYNF8AFrvv5gPCKQ4hflo9Zo2aoUjEB3DQ961Pjgjw
lNKLfwMGhlmCvmEL5/vDe6k919KwKVkbaUezBgyKxdZnoXowiVyLXnwwoiUpTNHA
RaIPpLGs8CjJoua7wuQ9/20sAp+lMMk6Vp65kMkAtscBpyvm2C4ec3Gr5qH9B/7T
qIicFivqjFeVqAiOAExxeFbHLQ7o+wSOIEk1eud2M9PqAv7kz+g7/NLTVtBQd9pO
uymuc0yw0/KbZBGTxIQWHblOYV/xLuFazUs7JuM5fjaJ3TRm/zIJFS1fVO/1bawQ
xcDKaW/KvfZ/0DJ+21daxLcLlGQhxptxjhmZMRY+UiH5lXmfVKQb5VpreuxR7dfU
2+Vbzbi5ZRSTQKajGnyCNI//IU9u/uL/RDdpJu+rnk8ytNZFUtiXP45Qm+t8IapO
UUzRZtpzP02B1gNxqut2JnRe+kcKkO3Z1Bz2JGuqw/chhOfeiaCh/B1sVXOjvO/V
Zaz0vK4XzHtoUsuuL6+n02d7bn9HMfl4dsOV6NV7jPUi8FWs4bk/KE7B3gLv48PX
Cmi5nZwkI2fhkXZIH3UrFJ0B2RRf9S0PAqolzAOMkWNrcHZbew7p0BqgU6/EoO+U
hASYFArbGeazbIkDiXow1gApfdbQ9iOn/0Mjdni59FoWkSwuZOkr7iyLN67+KMPI
uKCjapWqpJaOWvuhJDr39oh0gvMXHGHNBD+PJ43/BrpI3Aw6WLCz74CoBcSrFhQQ
3NfF+j+g+Bpn2bHI6AyqNcz6liDl2cIVCxPyRVBP6s0zWgroArd375YQGINpUoIJ
rc7yCMkPdINU5RaJgeLBRQ75lgkfMUhUftVgluwd0zod9FgmUgmuUfKCp4+TEJXl
zstQSN/6IDwbm7yxO3It9hE+AVo4dBbwsefRmuctlit+8XCD17u/FdgB2zkxVm7n
vucVH4g9kENAsNeFjLBQxWqOm/ioG8L/1gJYHOlzuyBnFHW8uqDYL3iZii4A8shY
Ob6y8KrrVVGe99P8cla1f8IizXZa5l+zutNBH/t9gheW8V7lRbZhHXqg6uP7PJ/q
bT80YMJN+pafjQED9Zu/lGVDPGwelRep1slIDEbF0zFUk7sstUtY07pEytg9c8fK
mauA5r+iXPYdPYej5FZZKuwNUtDlTNmA9cRSjF5i23kjqjs8u3OFoIvubk3VJu+E
uHXmDWi7urMQ8AwhnKdcTtPBDXdMIbIMfFl11Q4GqmqwW/6Sp/4J4USP/jrUGw5X
SHRgXVGvPSLtQCoDHOrtVYr8+wXTSKu1Uvs6n/LsNvSttU9pOrcjLjkiWUKCgiTI
R0Uhb44Mn/a9XY88GeVlwXRS5Jz3iEjoMkeYRXmk1kHolRW+lsMCUTl7+HeDFlDX
6pk4ePOC8vosa55HUdigOi1oqrLZol77u8aHLuzAstBdhwMhIL6aijBw1y3904rT
qHOA7EBTStFRMZOP6Qy3iF0q3HOJtHWDQdN4kFg3hjhceTlO97ehLmbvRO2JdguF
bSwHBWSfwPlbg/gO3QjlCh01Gfzo2QMznTYgPtTR1ZJtRXBLEEzC5XLsBC0gK7To
X1XRJrWzoME74g8K0KynKbVNi1y+BHfJPki24m10j119ij2bK+A8ckbDfwgT/pZe
ixzMkYlKxmekquaSnZg9S4fOnt5sF6g5x/IVK43ZvS6Fq8Q6ukYwTd3+Xkzm52O/
Owc8mV2bZsgBWMTfQWmoPIqTWcMU5iJOu+U7mtePwHWWUB9SjI55zOd6XkEzeUo9
IZGh11epjO9W35wLWXmHHOx33+jBThoUZIbDBpUzAZSXAy5q43GeTHgXFOvwDjeV
hH8AqVQlJuM1/qfJSD7nxa1PK3ch/6HZ4V/egQo7f75+xzX60HFgPuoMGT0G9iNT
Kr8ErtxhO45mGq2BAP1n6qtbc4Zt5RHDCyQsueIZwJNguT9j754Nb2YwFJAAFz+e
+6QYiYAU30QL5QonzXwqJDmrKHZ1LeMpdlGqNKsl5qCOCFaPLRKATGjF9uYSWQw2
lBv4spT1ghlmnCcZrXSjQUwrrEJOchGFqZ/9/Cc2bQe5d/6QSZhxDdZoQzivXbzq
ouhPYMGXSVOnQF/FqJImNDbkf1raN9nJuBzGGl9YVCeFnI3Xkfqk5ahbPjM4KR/j
4OkPtVtn3gXomudiA8ZC4J8F2H1BtVEkY5ERKXK6a3bilbt9zyCQoX8bGz4WGgVR
tGk0CjLopFgfbLy4z1UTedEiQAYldXThE0+WoZYyrjSEMpVblme2rMfIxTzDIUFL
iSfrh6tjsocYR/bNfYrwSCGcxfxe2G8xyDfvZuqvLG09l0o1sjt/VVMkV9Y3rsOr
zWVRxPRMfGkcqcqXSQBIFrjY9LzosHDMmtV4092nZXC9RnFTYKp+5f2IT17Wd40g
8eHjgSQL5L2ypxCHNru0/bkrv3f3a65LthTmiixg/1NWVEl4XrCfGcxJT1Sm14bi
Q6vHIM/v5rWdX9rNDemOrVP/e1rmldDKRW85CUpQnJbCMcbp+CuslgXRHKbbIU9j
hGF6Razs78QjqAr5O2rFVVsxsU4yxO+D5IKxI17UKEUNbeA1Kf5nGbDIX0WYU0kX
LUy3zC726c6df2vrKHD7lK01Yprjhxe39jXsKvx8p29XUdMhXiGIdwWI1Jnadk+p
I8aeLAsE5NJtn8hqbrHzznyRi6TbuD7ZtFTvFRSo7P9jfhYILt9GKZNuLe6kheTC
rHwEj98CqXupiAYB5uNLvbFZlKX0GPfX+s02ZBez4UpPgYYz2cOtVpoJc6AYdBzp
JdMOfQBjsjINiS9mk2nWIOb51KHz/+CDotIHeaR9HlhM3sw471bfgY/uXWVmCL8F
W41HwZ4b16N4VwpJXe4bdhDpENsOIqK3BNGIwTzOhQrkGgKvUKLjPx3LF1jjo3PP
xX7OU+09K7jW5Cu//S66H3YpH6YC216TyrbVgOSuHvntxGqVHNzrA8rQ4ehQjR2o
z2d8CL+fApSAuof9BH+YKmJTnt82qei7s30VlfXXGwR7Us2xgZfdtK/8SaAvwj7+
EMsQTSKVzkIiTSDcK65VHR7NaKdOl71mmD4ykpeW3ottCrEpouWYIU800nLLKvm+
DE3q866+sj5XpmSxJkK4ysNs3onogReMAw2LxtxZictaUBTvu1NAHpAr8Hjt1zZE
o3mx/Ofln3lGqGzgUeabYJ0y6KssXbgWVvaeRIZaE1qdnK2Pk1EyKiPJnQjXCq4I
5HoRZ3b1GNOOSzBacNKXXO444grRDWhRXzaZsLvdaRAOmJ8UES1wPUamf63zaA4D
8Z3PxFNCqaJllKPPgJhd7RuPNuWU6hT/qVqO5Wcza3fYhTCwVr0FnBGnH7W/djGh
h0DCIYmgGmE1CQ61+cU5V6oe8Ba9Vak/7nsFv0tk0nVnzgdWK1gbrEX/s0wL7iBL
PQ15SHTi4S1Y/alnNcxVGWRq6lMuISKuK4NsolShbbTi3jFCMQkbwho7xhYhghI1
9knAZCsRINu+A/EhzAi2IbeL1Kemma3u5M1gzAKuZ/lTnHAPVsiDZFgGVZ6n5fWI
KVu773HZKl69iHS13cLOfdPYIELWKfVXzUB64EJ9pLe4yzS884btx002u7gWBMjR
QL9NZsOGnFDQkba2Yd3tVTgGDyYeTPapTT1tl0ZQSAVSqh7ZOmRcmOz2arJvPGjm
1ciQ5u4cHwO00opLYPJPR5m2wFMIIcXp92K69d6oahp/rML/QaBC/3wIAVcY2RFv
e1UkHvB31knoO6oADIXjwIcC8UKuoJ6Cz6511gdqIFSA3LQzwVAVrSF42LxOuri6
dOjVwqS3u7WC2kEgME/GHvk7u5qVZvA5XOrASemRwWj3VDDX781ivaSyoFfKHF73
tj9ypsx/RQrKYna8LxQg6iM9dRPBvHuRE5bo/g5KoUyuSuj7+nRaaSTzAHiBJVtJ
i4TZp3aLnsQmgNOFuh9O6Nx6Y8q1lC3Kau1X7j7fdvaRu9PiP7J1WF4Lcq0tg+/U
LHhXVt3JrSr+LR160vG83BbqKT62s/Tl6ou831gHs+2F0DSKL9NqCExitFvZVEwe
SGYWIme9MYBk19vbMSE1i4jODD+SrSUo4CWF36UdmBZo3ieALtOXUJje0YG3zyrT
m9uvJeBECxWW+3ZEUBvDRgHshaclnVf0YBYqJUt3fK0Mh94km3NL/efyRP9cHrij
Z+EwZw5OvNk5PL+Te8wr5Yh2FVkl/AdfwvLkahjhbGfbw98i7J2EuQ1YqY37QTe6
Pve0MM0QoFwe7+bICwTbx4x0nG3WFjLUBmEwice0SrpLbDs+3SEnfj44k7WW1dbd
+yX2vXg7x5GRr78CmMSrCV/9W1F1o9O5leCFF0pgikw7E3xLeGXvqu5nJTftOHzY
VZUrE4Do1gOhV/swKeb+WQm078hGj6oCyxyV4B6GXEMBP8oJWi2TKqNrlIDf6bOJ
yrNFPEB0/yuUN2kPX3fCFXjSashv71qHM3MQjymYmpbvqfW6e9f9O7zfABssWTtE
vCq5X5MbwTjdqA4lFdK1F0gW1cUKcvAQIVH3Qk39LwRtmHjFcn0O2FhF5T7PsKKr
v7rKiWIjdhE4kaO4yVvkY+K7R2qWoKUzy3OrW1zjlKF+X4Ulpb3rUf5uDP9iUm5D
hJ9lLvcOj86yOHvhk8Kzdceahqx51JVpk1TeHmbHsoCKcNAdYE+v67Enn8jPiYdy
j5sr8ejfAJdjEX5EdIMr+/bSF2zct7dfC/FZk4clWkTHB+losFRPLBzWCHdABXA4
XZvDlCzIXD0AUziGt8pih4K7ysDd21NOjbJJHldEbu4U8qikC4YOtkh09l/ZhsZe
r/x2rmVwjwQH7qhexcN9G/gZ5Ed4vUgCxTvgRyb15j2NfcGydE2DykmqQyVRDDUW
OmeFvsbFfhhVR3qrZ+XErtZ+0dhERTpCmNIkhnxAHoEr24Dp+zP2gvLKbxWzU3l7
qdOlICwqjc8rG/p+9EP4keY++yqhMXb3PX/VygZ+C9QYvwWhxwxmJKfJEyY1Faq2
ng/8capAr2zVm2vvhOQaz/RqTPyMiEye4jUgTuztQeATESnsouZu6z9ZJZ/WD7xZ
bIjVep/wPH9v/chkQVu1wymIie6Z+RYK8o5A3IAOsokm9qfX68T0roxjjdkOJYGW
uBSdh8F+prn0Sqjhx9ns6xnp/1aU/ypMvJxQnuPPkAO5BKiXgEggC7gCcNSTOqlk
tH3pKnDHIZne2Out4niiuP549w4Fc4C+1rBj1p1JrCnRacUav3+D4bPdhNLacNVR
+o962+iBj5ebCY8O+mVs7ypd1HW10PhTItP1pd9iPMHVT2M222VPWIood//EbWuS
dMRtzji/32gQRTwkggQ/q5kyXaNRgwg02L927NoymMSVUpZtKg+rvtnKkEqRhuUq
0ryUCZqtLWNygLKzEsLluhafCzyASw/pUhdlRWWOPmq54TTuy+U9bDsdqB3dvyKa
acQeXX5A38XO+IZXML3jyeKZf1VpzatIQf7zCxvWOtK90oogQwLJBo6IzZSAJr9g
4DVAwh/VeF04Qz7IA1bqyHFIO74CKx3rMMvRRpqEaHoNu3361GifXVVrNSE1CHpp
P5R6lFJTpFJKSrbXAUIK7P+HAfFTd049/4T2BqxN/ws/+Nh4jLv68euG2ZdNzyDS
V8h8YJ5pEqZETbbD0zD/x6yXgRpeYCfbTTxk5hufAPqoqyJEbQ3AGP0F0vWQjpAU
0b9+855Tcs323kpU+YbhJDHd5LDh5LdRUxWzWurATg8Mec3gz20ZQ1tffC9LwrQh
ivvQkfT8VUZSzygrR+vYpg1hJ3DB+ILK+flLg3Z8KXn6pSfak31ltXJh7yzNn+w9
Vky7L9Q9BKTbQngo4BF4EUpYwL87svatEy0olzYE0Mbz9ifGp99qSq6XqL/MtS7a
6aQsr3QrDMo1iQgr+xCRCJ/q0somhEknhqjZP1sI+T/o6aUWSWs3U/prhG9FMokh
MZ5AZMrtUM+mJDxPjYlSZlmG3gTUcjrDk4HufKDGqfMvYNx4EvP5VJHlINs0AteJ
47OZnKadYISXY8fWaeN7Y0Tmqo0WE4MaAdinE24l1npgU80+tLJAtATq1qo2s6re
uz6iEhL7Y2742VPxK8zAqCf5r39/UWAlN/OQpRQcIC+009DnBJdv2OMGza18cv37
k5e2L9fOsMNlKzy9zYpO3WaoxQQR28V6YQp5eZ8iYFt1uPEFTfnmT+ctxT18Zr7A
nL7+HuHBCRTZrOQtxJAPQKMzvb6iW+dtYfRa2Z/h7nBraIpJ1KOC0ESeG72xmA4m
bPUubsO/bD7xXfS6+AkNhFvBOqV6Xsx/6Owl8MaNK1IwtcTn4yyTyV+Ft9oa7shy
mA/HsCbMF2rXXj6hwNbapQl/Jp13miPrCpkJSVApdAdThbQuIfGJRHFLe2BD2Osf
78oxBt3669KCsmmoKucyfsNv2sO0wf68LNW/QFFBdHqDVj8rA1TOEsp6gSThvwaL
QuAXmuPdJlegtv72kZ72rDbtTO6BkJ8QFeeQ6TwzSeO2AAzRGG66QRQqYijyPOWn
FHJNUlg9k3hz8RcANiIEi0hgC1lQy9jRlN//DOvoTUhK1wAX2UurJybXggWyLcgW
j2o5HpTSVPbsr+Dajq7ZM6Kd+sI3jqAjhk4EKU5sofBWVdJF2ojMAbKw8VjiBkOm
1ExX5OOewtv/CoYJ6aq+e98EB8I+hMxGLQn8+7TYqBj2+5swgkf+jYdkUN+G3PNX
JLTJfnUZ/BiEE8JA97uQqe57QW5pFEODM2dD8QOLoG5ODFQbRielvVtNVJFjet4x
OyQH5/q1YQW1iG8m2adGO2CXof5hrsb1nnX+Eviq3CVz6vJ4rLdYJNMfF+kvsXyx
1PqaNEO3dAhI/LZfBBeTRNha7YY0bor6gVVyvR44YhV44VTqSDjG/TzQe4vUh1EZ
anVlYl2QmUQa72Kua9APf2ZJlM/LGmWoRhWbr6YjSoNvIDVPBd7jAbj0H4MKLwar
qv+7dhDj6Dv05js9LpM5qOo+LBvE6B4Z7lRbZsxIFB7wHI1Kb8F6qZjE3ImRY9sZ
wR1+WcFuzSK7mNieBG7BQYhfOllO07xrl/AT/7vC8vBoy6a14lkpNdIOrTqCe2tx
aBdKUON98CUEBtNt4rO/sAxSlaC42iJZTFnkv897r9Oq+Iz8kz6uRazDk5a7EfJQ
skCvjFJMo0uH+vX6qN9arEi84sxAoYAfPiliBgjbeyuKKmUA0SDYJqbK2J3yb/dW
M5+bOdGvp8XL30PEle8Oow2zqxAc5JoW13F9GFxOxqprpECb+/FWkuuU7ErXqKPs
BHNRj2OOeTUA9FjX6KfGIwn+860IC13Xez2lDQidLKIrwDAhrso/+F3b48EgzIeH
YErAIEegdAj/PMd5uX7zgZ2/yKKoeOdpeyI13C/AiRnE0XtO556EglYeAUEDtX96
9I0/tsRChcBA9Zd2XU0TMcuf5r58Rgn/5E5Lt4wcbIh0Jy4kmZY9tw3vw62Gt+O7
qWB+pRlcl4+HbkV7Xi0r0r+czY06fxKtGd92LeVxnI8QxJW6DNNs7LxtvkvP/49Y
zXPDipWN2OiYJLO4VFcruV/OUcieRh9e+m6rW+Ca+T7WGmwqpzSQx5QKMPVI9kHd
otg3AerZdyRyzk1bwC2iosh9PTkOt+pjrW2o+WBuzN1oxsKK2hkrKrfdaV2dtL+S
Bs5P/O8d3qDfTDznewPT655QNR2yUGh5D2kkwoQtBy0CrjJZaSKRiSefcU2XAKry
nBEYsJ8aak1TGShrTLBEp5Icz/ntTpdBcEFXGe/Pt01f3sW8GtFACsrXDXUfbZcs
TQUypuLc98iLnAGsl74JX8e6V3PK8d6gmVz6M1fj3kmgMXmA9JixX16g9/6ujnSB
CU4O1D9Z6mun0zCzY213NKsSDRQLNTLhCHJHHPl7WX5iboOOj/PWgNDP/UL/Q52W
So1NtllypjwlRJvdDIjt1+5FinZuTnTYnR8YaEG2/sDLq343zQpBiCzZHcAhBd1A
s8ZdSgLlC7bWtZR057xRQB3dG3H1P7p9oALKZrcmKpVZAe0rWZJCjpC3oo4nBt6d
iuWrHV+SF0lZr0vztFmlIGCeWo4qLzGF7vtY/A+5Zm7yA1yk0KbPJ6LmURx+NgQh
kj7w4eOF3gEhVCI5ZnL4IuVc60Ypp8j+g9b75wHmueKZ/k+fNyljJ5CuIKgQZuib
Ag0XzFTUylmGkB4b6KrTxqSnAJCqYV6qwlP5xPyOLknPOaueQJnpvXAtQLz7ux0e
MsTBjjUGyQTeBts00biLV69M8d2fhfhYQkRMa1v1SNuaZZygFxcjKo7fOY5msAeQ
dkL5qTLRBZJU9yOoKPIyJdsJ+wvbXcfjr0nErY6dWHIlD+pWuMplrkHO7cuGMKgb
gMJu7MZ7KjyupAfkXqztIeQdQ8Pk8iqcyPLg5cE8+++chqUjp9vyZitfH5bZs/jz
aFUaX5sUEoBH3LJbdFgUetCOaH1oiVaPKYvZtydmuGBwO+XVulPS7JtuYE5S+exq
yCX54WPjkN/7dGjCWrTx+7RKGVuRhkxpQmZ52lDdmq7dUMJklIiBIoXorTFpUpiU
itBCWXVVVbRkJVpgaG6DZNu+DBONG0zKcMXOr5F7I5xxOn1sFJ+7MGTibgLtcXDy
pX9e2PrC1j4K9NvDeLKLMV5Yj8TY9Q11t1mSOP1UNeIl3OcGprC1Xzuz8Oro/KAS
AgV5hKuRFE+lJUQt/HqUB8pUPsm4oI8/Lf8FsPbF+cLJZhgxusRQfGz7iLn7W29V
+11mEPk0kdIkvsvVP4C9wPJ0rf6VMRBQey1bIPIgiyvFJ2sOFxvdZUPGay7IyO9j
TJq3hG+YtX9kW4pIJXw3+y91/PzCOzo0J/YQYrgG/WDgQ8xUG2ng9HSGkwjX5stf
KG/uQPyd39eoAh/fIvdNGJ4fyYQn0VDIUCQxWMCz2h7vjrfOnIQMUtbm/brAsmun
14LNeJdxKqzk1IKktrtpy7ABeOTCQEeanlFB7a81569xXRf9KC4Jn3NmBWHIGTgt
/qhThD7Fkb0XfgN0gPHagsiuaKhuninmAE/RfyPyLGD3Ofou1uHQ0jDJmyQzpxbg
38dRRA1MsfWxHu+PeOjYu0gqv3q5SrfKFNeJqCFmHA11GiY4VI3H9PKLzx/YCLoV
g4ryzmmpCxXEBEoezu9Nrjt6vSGQUI84FYp1kRK8xRRc6tIn8IaY6k5zvOspHDJG
n1X8GAYYrCxvnsD1Tk2Z3o4iRxrPbpLHEU/+Pa3JZ+N0iXZrI91XY8M37zMQhhar
J+F5hy/tZpY5AezCwtVUwPTJE9A675XaJVkKmEZc5rFDhDeVmycA0oJJB/s2orZv
uP+qJh8Tz+2xQ1DT8xjJ8GEAwRHjLKch6tVCotBJcyDG+Jb9+yJYe1CXuvnW6Wx8
R5QDvrxdT049dWbW/tQ10ZMXBj21/OHXZvfHdeGMFkFjrzQNvjCaOrzwqbbBbqmA
47PMs+DxRFaAMwE92VoRYEqgXAfAmus3Nb8pFnXb/PThW+sXaVCIxYB9192P/0eT
5NAFudLrBYrteu6ZwGT/KnMYNH2BwdvYOB5SYgHHnFmDOuGZeMM/Rt2hJ62/9Oo9
VU5XwQhaf1jZMDaD59afhdcMCcVJRV3grLhJBNlvKwgrZl282XJXX4ReMJelckIh
DXkoyy1GHPviGyzIz+vL5PN5EF+Hg+eAW6z/w8mh5+dqXDAHcCHQ/0TIQGiMNUzt
km3oSw9t5ty/YGJ6fUbGrLHf0eBwK56iMqlFLkuzKCDpnRTG+mssljumbqCzyGHT
e2GH12a3DBeD8e5LZXzt0lTtdo3QecfAS4A/n3bSJb65w0LmNMnHqQmzpKh226PW
/4dsKdWW0i6zMbrK/Uo5VcHbJ8rDKEgkzZp9PA6SmLofiVIxG/RIFwrJbz7899to
mYHLWjU5xg64MK2FOvdR5MlWaBerh19E/24njEpRL2NTdC28zROhti78MhX/0k72
5D2fTrH9mc6zjnHOPG5gdGyw22GxZDkqgAsI7ULEFO/gUPrh654foi5vgfctpow8
jC9IlXBQHMOoFzvZqnmQys+zz6T+bdrOhND6dVVGmKK3Uri+60cUrLOf3EQiSgXR
VOs3a7t7Bj2thLefsoo9uXR/2GeRCw8OueQq1spWSqMgLw3+50ip2VvfXGN6QySa
MfVoOlwpsPMcNk3XSOAoajlVj3KJpuYMzsS/1AnUUeaLXX5st4sViVyV4b/rOqdF
8jEHCqg1JoYZ0W+tw6ooGcmaL/U+1mtZnf/Tx+BCzRpeY996cICHt0fyRpRnIooZ
DWMyVIrx+NP/2XykbRRaQtL6GtKFdYh+wp3/Pngw1YuNLfLr/NxN7TOXAHYhkVlD
2QV7NGTTJRetuQbTVJjkfh+ESDKjwpDba91X9PGW3Ryt7efSQizIuxTMWwqgBJ24
DwhKMjunZB3vLwttYRmpLqXsT5YnCu3Y2b6KNaJAyBS6uGrVeYVCFXSg1+LCE90Y
6xeHjdeOtO7MRqlUr7gFx2kz4HBN9mVxKtz0m9KLZXFky07wksAbZqAP79pb/9aa
2PMnUvYmtqrwWDOjmc1lwMNrRPQRgZAEo9jXwY/m+lf63rAkUlW3O1u5kEydcqgQ
a/6OY0eYu+G6FO53C3KlHMsdi305nReBBjp5WkGE5P7HW+DRaJqBGocAy5F2vPuD
8HzxkGcGcREVw4qvUeysSnvMPx1uyo8ebw6UPJAxBAcw64JW6MZrP2XU8UgfKtFd
FLEIzmteMoi1Sd+fAW0xEWqsXJ+XvUNhKeISQJzI5LK/tYxp5Pj0Ytk73NSY7JHo
ql62vuxiRDpvPblJOnDWcHrS+0elWfywxE4qQXsX8fewuPdO0/6RpbAqPTJ2/xYM
/qHJEzJUgQQIsRVsCsmBLbaFPn4Gmk2wYWeLMTUmEB0btCfjcRGNdt03XrTTDecM
nB1Kj06t3qDtZYzc6/a2YS/LwnqC39wTg/UIfOkSZikTB23qyO1uJbGNIZtuAoV8
96lW7YIF6fvz2W8kwli/HWdPQH7U4a6HRWuAK9mx0hoWww4APpK19mMCMAWESzMT
JLNntLh49MXYhoWiI91uY+C8mJJ2cjNGnKWSqD+B0Q2pw2yiSVWGrtUrQEMC//Pu
7mKHowdcLeIgPCnz84Twxj4M3IN24BPjfTwLyASP230pIavsNRmpm1Z1AFDCoZFP
HvL2/scvAdbstI7qUEaFN3AQvLyaqXAdfNxUefiJT8uDuITNmPRpf+135rE+3rsr
X+wbGFzXX5Dp/1xflIsghBZI5jwcs98tN67Fy8pgcWkO4ZF6Bv9rDbN7NsBtfBUK
eKSM5+LkvkaQZhaH7DIMG7wp7KIqzWuKIlLsmxS/WaTjUq5O51PziC0XzD/XRlXh
KH9tRnlJl6/LAdlyNVVBMfKbpf0vDZu6ZRslVwIzkgc5vcmxJwqroyBx9mZ+FQXb
cpV3jY5QMw4y/UxFL9cUDpIjzvLYxHtnoqdIibH0UwstbbCTF3DQdJWSSoOrff+C
1/l/T6qhLXyqWYLrRbQ4gcB8Rb+nNSjA9CRWnWVCrzu2TqdqOsat0xTA3kZowmnv
ZRMdb6wDYvd+bNoQjJnSO2rOy7kgDsIvqnhRV0o6GAK+zqTXUN1bL2WbBymYxAai
3e21Sk/nXGY4rcjg5Sr+cSJPXV6wXteuUPiG0GnPbFMYBhNJT3ajcuY+MNjYAMrq
JHOUEHs+4cOznR0Zos3DG4lxwOlerew6LCy0FuSOkFgKiIJz2IH0eS1fJm13wClo
jMfsIIyoaErZnzSj1yadty1pw9LQeU1p5TDupXceVXKEQzYohezQ88g/3bI8ohXj
dWt1MNhUp5DnVge7CbqhvpFGVLAxHnFw5+nqy4RyJL8pLk+feSPt7DxNMF4maSGb
yennzSETcY/VnSF8qpfoAeZs0Hfphaeui5K/8e8BosqsESYgB1w73CL+zbRgNhaf
2M62S8qYQX+Pksg9ipXZOwy+zaFwD8oA4SE8YoE5xP5mor+bi9fp6v2pi8S6swO9
N5Y511QWhbpHssMsxMsvm6rHDhbvWxzfzV/UkMpn7/1ocakV/+kwj4D7r11mok+J
o3+82V/3IUtaunVwHvNESnKUU0OMDTUawXDkXWGtI2u/EzosrzrXAiH02Us2PBap
RkkQq01TRYgaeLmc+phNAqSSbM2eSPh8p2YFORBKZmPpqk/gwm/NweKl/cxLYSa6
mZR5rYHt02e8V/fCxW8ooFV0NcsGr8A0Y9Tv67gWOfOtDd/RKh8qiQ5Xpx7R7I4f
1B8n6cMU8eYmJljmFnWKUW7Usl5HNHT+GrwfphPow+5rtZrqyFidPm/Mx7zfKuiH
Bh5HQL5MLk7VdVAvFrg4KoOtlxnW/OZ97Kj/y8rOw3pQPq+Cu3VS7rzrOv4rPaTu
qftVUNnSVCbbUGSBYyw/x+SEgVwrg177KuaqegjDDYF7KTu3kKmsQyjbkj7r2CrA
nDOTE+7yaNEzluhuUOntYL/EfNJeR/qWUJgYr76vFNqi+C1T+n1QEzajmamqqV51
M+jyVsnw7ZCtL+QRpsonYelk+w1BGoV+95UIQSDwi+DOr4+SRokFV+YeN4j0rihL
2fd+g8+g9H564p60GqSGzaYN7tSYRnlCDqmTzxyRLdZzZPyqL4VffusCIxrpMPDl
h6hT3WK7ipW8HbbLBSgO7tkfJMbYGiaI+oecR55Af3tiGmg9lCHUMK6K6/+XmiuU
t5lRW4MJ33i9I1mSVgijmsQ4tAqFPmeUSL0xy3H9sL36KMowNSKgqnLlGWTHWydE
JXIrjqLcKww4vRbJJpuw8szCmWvIvj2vsmRTQK9QBXe0wqIsJrsZlTi28/CszTU1
ohg+Zl7se+8awTzuvI8VFvE1oo4Cic3OZpVkOnbWq6H9Fjbnh7YXtZ8j7BCSBMaG
sfC06zQyJxxVf/oOwrIqpk00oPqVWzSkzzHNaOmZftQ4gjF7RQA41WcJKPTPH7fi
tOL/Bgkosr+3aY8rY1/2F23G0VQ2HOPdqMv+/kGUkgKexiPRJ0/F0ik8Gmox5ZKM
0tm4nsfCx79cuomE8fvtfGRsc8P9gl7xXxAeoleHr7KPrpeswwiEEbXiNSBn7wqY
Z/jpJE1n91S+x9UYZcmfjz9es78ydqNZj/LoFwdqGwXvJj4dUMZ5ckjMti6vr0mq
P0a5zbAZ7bzL7DGRhK9rK9oNh53BHyyqJZ9a2m859JEXIxyJQ9ci5DYDoLn1FEb5
oXWffzHTPJep5/Xz3Vjz9Coc9hTCnxvujE1IS5fTbArg16kEr5CS/Jnpg/DuPSK6
nccDhrwdQuRJfVj+WebqgKtS9zUBogJSMXYinlMqyA3kgpVFqCz2CU+kBNg7wAdf
TsKKwQoZvKDhi5ArqFsRpqVlV/9h+iWoHILTwCjYqEAvbWCbn4kNLSIKgBHTkq9X
/PhTuTagTTqj4cg4suMl73ti/7DIhJJSwwKOMYOpGbh8EN2nt85fteXFSPf7keTM
xqEt+p7XiF/KGqp2R7REt9BthBFV2g/s+FgixuPRJJTsKYwoQr77dNM4fT+VIcc4
EcUV021e46QOOEqj311qSTUFfNNXV2B71yLVEog08gN3oCSzNhZxE1Uvl4Y1pN1V
1GsWXZz2lRiMKyYDn3WZP76LBHutOP2EG5nYurfh3SV327o9E60B/Ewpbl6oFdm3
eZq9ZIAlYwa/zoVbqIL0cOGHFjjJiLDlEP7avu+l6d6vEjUvbdMSVCQocpa5an7+
n1Icg7npELrNZCG0wGW2esk63BKsxptJxeb/MOWmlEITU/kKTt6ekWN/hblcoVMe
buol0dPANGRjcH9gj8zZpA8Rl80gFxyposiW7wFkX1sHkMh9DJvd8vPvWwOR6ehc
SsVeBvi4rlNuHKVwigqwAQkkL8jDpRTWx+HOqDj5x9wXprFjJux2Zx8JM5YiYE1x
P4OWcB9KWYCoaHZkWsRS9SLh+7ThLzGZ9LsWly7D1HbO/d3aTW/5XEay9GQWsNUu
cRGQX7RoVNX8wRiU3fOhJqhIafxIuVoY76/AhlK1LHD65F5/5OUiWGnjl3/jZ40p
HGXCvN0oMYFSyUCjlWMu3iDYNISMy2MllyaKvnVAzl78zfWMyLLPmIDY02h3DCHs
wo4sQUeD3dbRAzOnCYg2LpZJ+51vJd9g8OF8Tgzl/aoAX7FpvPAMFDb/DpPOMCSh
FMwWvDUS21D65dRR4QID6p+HngShPhNaIkFjQBjYoo57OiVOaUv0a6WxTefZbBPW
Tb4u7gTnrUpm/HQ1U7pPUQ52qOtoM3xlQjN8JIpMHsBqBDDH+UlCECXk/zimQoW4
EnImU+I2Ko9FVr/oX3tiQdoxH1tlL/j+UlMFN8C3awIeuggkdcMnN6UXkH/b4Ugg
yiXsJDWdUzblgHuWMHp5waCYFX++ZOoYGvM46cUgAvCP1TWnbcs7qo7OZM9htGI0
1XGPQVGwbJ4nsZpOpeuP+7P9BxUrpP0+7eR6mdx7tE/exv9vyMZG1/eOyrP6TY80
g9/CovVEO3q21JdU/3LlP2QRYPRqMazsZfgrVhh8lI9y2vlIB7tU9lTofgOb9ns8
ODZ4nsTj9exxvQ8k69JaORZIV1SREmrfr7IVCIOwyOjeS5SXO5LJWRC+felIriYj
/6Pwdf+78ghl+6Q55M+4U9bzKRNDIJxX4ceRPZoulwZvMR5nJy4pId31sgG0RxYy
O9FZAaRPZyIYrLeCV5lL/0HLtt+Bh2GoY91OqkD+B6A/GKS0gncfj8Et2gQN5UNv
GFGCmDSJe7yB6t4vN+obZcQAH+bcuZattWoDY2jgM+aVD4FKSg108mt4bNeSmd/8
0WdMLdKWcf2LM4eYBosSOJ5xwj7d2xixDgCQV7ls+jWxHtoKpmTFfsZFZt644+r3
qx3CcqQSkNb1g2F6Y1Pa/j0xNKoHpgCLjUEbCKzGin9eQk0GXwm9iMRw6C2qnscu
pyIu8daXWNPdLTRkeBUSSs1S4mQVjgX+6g/x5ow/YFNJtFEXyGC7Gl1ljHbBjehP
xCal3I1G1zKxlZlZCYEVnteI5s6fAYjhB43z/fu8knZ7u4QilEfEjqgzidZeySB0
tzbk4N346UOSR1bLCN6j9Jd4KrEUtSeahP9baOXTfLnFPiSArhTyUkwH/8yWfwoB
PAxL4LtzChAaDP5MD6am1tOR1wi3vbuGwfLHRSHsEUI/fPPY3zjturFC2vV7AjrG
TVwwRDJvcrI5mM+dXrRzWD2yNE5RW6RVKWoaaryLqcCdIyLjIw49/rp4lPU7yLMT
6z/S+oHTCSq66otzGB4U28ewqB2Dx6snzlwNJ6/3wJC01KQDFGDoWTATM8LZbcJb
8FMBmOWrssD0N2qb40Y4/HmtwSsECQDXLl1HTrRqmEeaf0iAtc0Hka84hZZqXgg1
zYwaipj/FAOowlE7Qq38JUwRDdOXKUrqq8nzSVeyW8kk+DkTyx0S2cwAaHocgToc
F2wEEOO7/PXDcGG5H2Sy9msexO2jflPm+cxo+nmGWuqUlO6Z3KDwYyE01G7+IdNW
tT3jSl3KxDlcrqcJspmAG5f4iMESeMU9ohFQtjzKbkf0524/HvOJ+/Rg8RnPxcne
zDHFJXV5s8dYJ0OkqaCt9CpL+AqyIzTJYz5u6OVGhIv1VKD78te7xtpLrxheP8yB
5HwCY54HqrltMBSy9iwJXf5DJrahfOxF6BhTn9jvBdkz6eR6tNqdYJlVM4oLp7HE
jHcsrurb9Ya/6J4qOTivg/6kJhAMaMa5QkAbHVd+PZD+haVbgSpDxdx4c6iu4DZI
CqISyyWFWxXzaGaFAZ/XmdCRWyOhwVdZnjNclGbK2OtAD1vQoDcdqV9Opminxj/d
JBoMTJpdE/zw0tsXOSsHX/emZCs4gs0R5m/tj6C50NkWX8TNkm0t/FiefCbSqiom
4ROjrUhxkXX3foFfkLd4GgLTWvnW4U3nEgXGtdzL5jMMfA9at+9Hx6UpcZbuJrNX
n32JfMFEYYaCKsNXNZcHaVMlglcC2mYPftnqfEsWRYzYyGmZcEwo+O5DEGWNshVB
eZaNkzvYP+kUehEG+1wUxBbBxXnrtxENl2WkZi4f+n4QkAtxdpETt7PHbrg76Azc
bIm7GcuTjcCM3S1d9zvRwJwgAT6y1fB68jlmTUcvg2UoHxLqtD3MOggyIx/dqLH2
ihPm47Uh0lQzXzGShdLBzpVRYSlTpBxCPyVz9UbALQAd81Ms01Ehnjzcc6oI4Bz9
nYrmuLm/bB8f8pa212koaCSSbmTG5/uLAlcsTVKgYELZfSV6qmD6i6G/HDav6dOl
D5Q+zNaYgCGJotewAaVVvXFBAt/6RcrQLSa+uv3r37hiEMgmJNGvSdHSt5pomuqQ
09nHl/FaJFyZtrET2lwqAImY1QUJpyxLl49uFWZESUtLrc02AQViFWBbsaQ4KcG8
vDPx1vuK6F4ZCG64aiC/JIhuY9K4fcebAsz0r1u0Vx0yO7lnTOGtN7LZ0MkPa1pe
XAyOxWy6JoaGAk/PakSPy8QOwGieGXC6GFuF2TpkbHdRUuvyXdIqevbLubBZmEyn
dqW9TxjaiP3ipvI8/Zw1iGPXKsajcbL68GkeNSKZL/kexiVtPFTKRff874+hJZDm
0mSIZSxg7iUhVtEQ7mqlUVdFhJ+HRbIfimJK+39gE4liYe3KWHRgStfzgW9AH4y3
Xgkjx0xnE7LXaQHc1GCbWPV2f+mWuklJBT1pceR/gA2KAFvyKFv97UFvWlaHXZsZ
lbinisVRkxenpq2mINhsV6g/wVPMF7GDFsH9/AvI/TEvSTWg6vkD2CUjSNAOI7RF
Y+OXzqIKA2HyU+MPi8fK9kPJjX+mgnbOGzb/Ai4bDC8q0E7kC1NWP6nelBL9ezt9
iA6ipTuIHKLMkSYouTW56bxu6TmEWZBgccp31aQGXkJaCDYL+RphSbRwDV43xkye
mahI+mdiwilDFEWeqEKGgy47xkBBZ6Kjm+NtZdF6nNXksy3J6xARLQB/SRcq4oUj
Au7ECW7H31FW6S0+83d+rRk7an/0oO5dg+B1lOYWUfwjV77lWu9APsPcdhTqfhaZ
r9z8tcjl7S3TpGUpwGTnXqoEDMW2kesLMTp7df8rD6C52z5xZBfsA72qyE5jQI24
KexsjNfWa2yyRBxja2G6Rn1vulYKVMSDEvIW28z9InHAz5nkzepTEW2CyI3cL4+m
kYwHH26qfoAYQw0xbWc11e0dpnrvd8IudkBDPaLUz55UdGMxs7nDIWw4PPuGLqTw
0ubqSQxklLz9uypQOD4Ab8+2E63U5vzGuJvtdjc9KkbnZ/cpTSPTtUYAjihIlMXo
Oh6PkaqpHn5ymtOLT58D3xYyg9ikWrSfqq4bdCJZZgQUCUMaMVNo4TvsQ7Z0qigA
1O44z5/jOkDpkjjoJSV8ziRxisuurCWf/J4ON+3MIjcBXNFmHSB5072e+ei6Bw0j
slJqpcxYX4XA5VqvroU+gPkcp92tQLaD6iSK5PISkCUKtt6lEr8/xIaTIhY4ObsI
AcPdWhKZ9XAcg3SiallV4odlmdINw+n/rvSIAhJpKMbDwze8wVFeerR/ig2MgvAy
Xbgupwp61LV2bT0wTZAoi97jY9TKfzZvk4gHXsanEQrPyRH4idUY8uypp0GJA12o
M93JoTkBCtAwwCdPeFxXf5ukU/ah0o8J2sFzmTHkMOH7HQUqo32SKGJuFyYxjd2k
QDmVVFutfx4GlcGF/9zi1Y1dhkC8euUFJ1aEeF9uUVI2qT9ScaHxHEAZVwBIfRxT
GYAAqH+s9sWYtWmD/ImX2jy37KK7f8A8kCc7d7mKV3S5z5s5w200toPLbWXJhZdR
S+fvOQQjAQ8vgUtKluvD1qD9fjpSgT7AKGW6l4NNh4emh1jaKlY5yFHWJYiek8iW
3VuA2oHPQJNUzmqRlW9EFGEKrDevdjoC9JkPRCwc8HJXAl7L8JPjesoJQIcZjKZo
J5ULWmPKyczKmg93Mq4I0nxPyLa6dQPxAyvAOhzoq1qHQK/yGDRrRM2kT2DlF09W
3uH0jHeAW0fSYmDwDRa4WEaZExoUkF4BojwaPuCt+q0urlkO01b3NVUSsi6Y0A26
uemJ6gv3T7B31t+XfkBYiqWqZoZXpIHyWGV5XdyhkpugqYla0OXrAu5EFDuSKVTT
tmVUh6PMOXqRw/w1KOqOv88uO+JWtiyCHzT8yaFV2KSVrSezc3clbqiTuqtegHYs
LEseHma0sEmZjnFsobV1uGzQPPdq0Cav6ur6d1D3oCY61eLuyOWAbsLOivsSGkjR
BWfARtafwCQ1Bwp3dxjbZCm+kXv75z54B7hhuFvZQus1EPWYv4632iLMR2CIadx/
beIXKzvQpv4BQaPMV6zc/iKWw0nA5sk7Mn9OSYh7LvOQ+sdJIAtiqNZCA1W+RXo6
Q0fzMF1KlTgchAUaPyZizyv9BFCTlt8vT45OO035H6r2HG7hVYwxLpo0JCiM6xK2
z5O0gKblGu05WepPqU7VM92nzUyIwNutDUzeo+PHJu9Hl6MBZO/h4N8vzx+a8L6D
UKmfu+lFngIsK/4Tx4ZxrHrpnReeRScZXJE3VHbqcO2anlkJcOVDCvBdg0FkxEde
5/+/664e1QWx+KItgoLHiQ4GkoU3GEr5cn6VTfdax+VDY0GDubSOeSumsSWGIoIN
FNqVCHROPodj+5QhmhHBGNCQP+aB5ovI6cLCBVm5uYFUZg+CdENd1kF2PMMM+3Qm
NkoV3xB5R57aTXOsHu8t6Zy9c9Ljwv7pliWLuhFgkY74uMtH4Lj8+vYwQpg4vef7
F5vcg90ODCdoKLmzKI2dGhsZosm3L6/nHer/mTDdMavVAg4vDSwZTT6v8yZ7zH9P
5Rx1DcLh43sgCO7nzpdMGmcnfg2lm4El79nxgHcMjH+R6V7VxkvUqvonRlBgPzcj
NvmoCF6TINpY79qVNN1T0EXpDrR9L5s1QmfpP9IDY4p7zKidKeeYbY8hXHthNCdD
ojvICf3PTEK/OMiC+Y+6DVHNidS52g3GUdO+5zkrzhwMqG6TmXSOK1l0NxUNw+aN
CShIo73DH4Jr92bCX0Tcu9dH4AEiTMNcf4XEQXGnawKqbWsxZIB+tx8Sqymg/g72
2JwBarZDtv6fKEowm7c+QQ7TwCs1MgQC+sD2cwRb2FYQUO6chTrhBrhqNV+abiZ+
YRe3Ewx+nQz+/qJdYrnOE1eRNrCjIUpO8YhbGTYSuxcyqqXpfl2aL2BAKIYbXxJC
kgMgsXrBFO4HCsuqtZeanYixTg9UDLYCCoApD2n5Dd0+wga3BPkWhRQpdIZC6rXQ
vNIVq8dNiOuxxRaJX3bR0HpsmPYhZiE39u5aiEl1ixyIV2CTLoL10dMJEpPBY8WO
OY7SyBbKD+RmUOaT1KMDBDVrYt6Xll+nr7ZbBY8bqS72Ys4KQB8cYSBAtVquqIsy
8G3AEJ5iT7AMNyAULxCRQcYFO+QZsuL05/HiA83Tv+TAPF6ToX1zdamCO53CQfCD
0EJ9xv/P6ikUZmsnIGizrWKnw5J1X7LYinvu7VX2hJMHB8NyPGzH6YloAlcIomFM
YYc1GUMJbGPsgbK+6MG5+EWtKjxkhLIxFMew4dhN38bNvUz4hlX7CN6h4IMttLJk
ItmNRWPw3jNTQPZo3CZIRU0EKSUsdoTrxyBTSrlNr3AHH9+vJ2ToJP/2EQV1vfte
S3GiDhTbU3D5FwTKB5wx/S59JqrmFZiUsQatJhtosEfp665F5zKMQ7hsazu2y/HK
GN1/3HnLeHUkRg4Pj6vVAKx+IGl72+AyHXZW94sqZU990FGV3Q7OAwcod/RtH39C
Mcl2pXvW/DYmrBK8Oj+WUEYA0+yx+dtHwKuJLBWoVmsKpGf6UqsNqQDuhZPWXSHj
7u65q2I6kOG+gSvDw8ZnFUJiJZ6ekMhvl4AXQPh0m4JjlYhDgzJtJMpNHV7R3uf9
mJt7X5+zTcQIQv7hnK1U2Lh0jMcUOBe5V2xMjdHffsllpSn6YlZcQQ8QmLVdP8jY
QmX4ISt4XLUexHrRTaYcQJJGOBZ3Epro75f8Ln7oysHn55unXnRJJ4h36NrN7QzL
mk6EHdn75WeoxtHrCgvRlZOoabmCj8e/KANu1qe85rMBCXSO3KLnTTZkSFmlqzCl
iGLeJXtsOj8sfcCwsn4Z/Na4EqxTKXTVMtxx4qZp7BZ0N+XsMP0X6rZ4nXUM9VEy
9eTj2f+4JnzGR3OHe9mFKy+Z6SPThthzoeMch9sQdQhUF8rSFLfJ65HvME7AYD6w
zP6KID9A4EeOmObnXyiXVsBZYEKl6KZDluEbnOxIb916uO7xTlBiZGjh+BmuefVr
q/GyxizWnOauGdMAY5mho4GpSVLmqfKDKcric/+CoNUGgeBBBixMUag90QamxrVR
6iokJ9eIywG8mZpKYY/JZuIQxe+4oXrbVX/nm06J/U4k1w4Uxx06aXNZngzSe53Z
9Z44OnH7J1+uKFAgKydToIzrX1x2JXAf7f8qznQq/edqs2SlA3eub4gVzbAsbnwQ
Kb3KrIYhTW/2YpAh6gKLcpCJjkNdBiHU4DgefigfNmFznTjAOjxXyodmFPdjWhve
nHiBvHQia/2zaVFBUQ/+e6Ojv7nAskt+4C7Nvqaa5U5yLHuIxEOCUub5jds8v8SD
zmuHSDlM6MgF+7kNx84A2RmFCBRjbDLZZeb3jdMIzZd0ilRn2kdhFM/vBvJw7kfG
kfT91HRRGfpzsYvNwVBitW09lDyxkc6SX0o/qhvQFls5re6frQYQs/Tc2DV25aFH
a7ADIJPfktT58ZHJkmZZ6WtOe4K/BiLnhrl3JoOIi6iDG+ESMm5oqTbD1N9SIiaN
V08n3Z9Z+A9hgsns9RfnHgOoRePJW/oLIUifbvFEt2Sd4Cl5YoNu3CCghfcbknDh
VGEij2W0EPnM1wrz24h6fgI1SupxQxY0K3L6ghtvrzn1Mc0o1L1ihI/wmqyTyCHm
Xn38lDXZviStH13M6SvMfWRvUdGW0F65xyi3a+AsJui0hhaEyr0wBMqa4Z5uw/pK
le2y2uWokz0TedSuRGl6DS6LOleiiP6OvP6xIVdup2qBOIXg6k71QTs+Y1BP+ZZ/
zKeZbapzZcshjwC06sJrSPu0MCk6gpPrbMbDmtmYh4Cwhkfk2i0W2RybrVnALzdk
l9F3cn2MZ1U85r0hvJUPQ5UDMzYAjqbClTnSibFtoOkq6yRwN38lW3dkcsw2dftp
WLzDbBevCOne+8gJwpYxv5pNNLBDQzTsLusb1oYOVFd5BlkQoMqkyeex/+BlOEtI
DZCP+kzrvaXo4pgYn7Rk9+Zaue6rkmSZlQtH2rp3+i8i+utl3Pu3UKDQHQjg95cE
HWfq9HyVkBX1g6eic58Pfbysht8eNIrxtlDqCxLM/OO36Af2MLrC6158jGNyA/7B
GAWSIWFIPKJHKrGq+jTFi8l02K5URHYTYpHdBbWVY1rVnAvhZ3XWfzCTEF/S0KZr
NeelSn5H+BYm13AAnjcinMT+Y2xXKaXlUtVYtFePGIoq8Vn/5qTO/79qx56rQctp
UVuKWP2X/MXlBqXDkpAQNsGgDrO5uKSg+zznbobjSTbWy6rHeEAa9wb84SYAnaYk
XdkHok5QscYSkDaldY+G3U/WsIvWY/lMXFPQY2ti2B79K2DllISKjGoPka2dr9xh
caBhcJDOi2ES5PgYXWnNDe69ciR4waOv7DvPG41c8WBAIC9VYL5cDFGo0CUhf5RA
VJgKKHEXAhZ8QJ4tw7jmvVKV1DdupErpLoShdt3je/e9FKHMmzsEme19hXRKotjS
sQ7esPsQy1CEdroPDo+DBM+KNH0wBWSC8Jjo1MZcdvkNE4pxpEpKJ2BegUJRahmy
BmvjYui0f21pEWYOmxcqCnXaJ/OG3IWP+VJwqQY6qCEmQ5vXcRKnbL3pcg7/T9Rg
8FfbLHB3upn2+m6xvkqCZaGcittoBc/12Os+dtAcImwzl2pou+x4w143/BKLSAMs
HiZpbMWqELq1lXENO95hYBh1B70eVlaxxfjjBy0o9Rl0YssF0BIs591WUR3L0GXg
EegERdlU7+XcoVv9CV9AEFJZ1UhpIIWkJHsNWDeYSPjwjp51Lmzc/eV0/0m0Bf0P
NPkUbhnEPM7hNXOrcBNM+oUwwk0rPoGb6JXZmtWh9ojctLWWBJyyBAC2Spjm81D5
PDvMlQQtJy4bbuKwZAIdg59t/N0DdqgUXSIx7NKrgCOLJRTnjDB9rzTIVdrwliEk
EHVxe0g2+UjTI8tSJxxJsQi3LpBePcgJx7/eoRw5/5yh1+qgWiaiv/uSHNW4AlT4
JnMw+3RWpcHoCs6O1ceKolbvAYJi5/uji0DVp5Lnu2dlWmf68McT7hVH8M57xOie
tP0wPDasPswokDJBeBe5Ite6n6ctmHXE28FJ3RbOAa06rm9mmQb5T6kwIYlcWJ2V
Pq2X6HAT1LEgK/3q8Y2L25bK1i+WCCcKLEYXFgr4PWi8s5e2hL3M/SQot0y7V/hU
7AjAE1lNo8XVhNdFkU/mpwMFPehlVf4Am0U4q+tMWPtOuP+RIkMK7bscNSpP03Ee
f5O31NXS4rqY9eP5TkH5cAJKVSy2JEpawVA3BaA6XPiKlsug/wesdf20j9foxXHF
SfoTNxuF3FYeh+BYnehBEl91unU+XdkIN8l58k2wVzR8UwWUdOTjadL62iuiiIap
qS8ValDz/fnvbONE3/BH48UJ+Eu+iFFSKOOCcLz3jf1vjlw2NLNhTyBIX8qYUTzq
87a8AQiukpaLkp/niwSgAzH2c1e8e0Tbubri0DEEsWz649lRX8SB3wYla8lAoYfY
FNR5ckyKa8oHFgNlkrmCFcD6FZoBlQjTOVc/ha6WilhaWkVQVJvFuSWeSr04inw4
ahrbjpOcpK0mK6rP/WMAbAemk+j6CL/A8Z/SkE0PDvtSbuWpB+M9zxvjlU0KCJMU
r2l8FFS3BgR8SSXXpvj/Pzh1QaiK6kYIkmvcDsGrb2nS3OvKvLvN4Ie4NiFQpuDl
i55dKjzdgPuRV4nOHv9YBmyxLnFTP0lg76CklcqI+l2oZl0AOWb5CiYLlzV5RxYL
lDYAp10iabPTMeBoFKLFtVLYu6EETRh0bxgoRbTouHjCSXhtK4iyzT+1v8VHYLIs
VIMgW4zuXtMy4MYu+DTUxKSEF5H3rS7JytfxijOY1LTlbLPQGpcBXgX+3QCukJw0
4AT5ZepiXQ1/Pha+PC0B9m+rpKs7Oyfa+Thqdq0xwO7ukut+8JFsVXnNwrrOmEMj
IVTy1TVxRiHY5Z0lIINzQUTUYFx+yEBWCguRKIMcqIUgN26Ci+GhpOPsJF/0lHSk
4rx2VtWfUpd/teLfoxX0/pbZIVgMdCdHmqXrVz0TwIn2Mx/cfUs8asxy8CLKvAwV
0CKn/1emXdlEN801VETiCpDA2TtxXnnHNmPColN78EN8xrXUH5XmPEj+Lqy1rm/B
cWEaeZ5FqAia8tDUsp11iNF7kYcPxdeszR7K0n1Kf2606aNkv3sjMvCc/qfnLkRF
Ci3nRkP4Q1/KIBS5CvsNyTQx5zjFZWVplz4MnBK3prfZSOzzEVcrNnW7dsDQtl9X
VCI7suL+Kk95EmWwLCd5uev2fu7ac6aysME6WGfV0/Y6akP2sxuU8Pqir8/T/2kS
upz09pLjXUIGk66nYBCiol1tOVzJUBRfnZNzdW5xBxs1RpP53PAdY4YErC9aGEhY
rAglnqKaI8CT0dELb6/H8/ZDGRYp4oUGI7Mb9ZWX59b5tEz1sxI6g1qTCSbMgRRM
6bJbBf4Mdy4SiedaIO6UIbfDnbednhzhJ4GjaHgaxbCd2xmVdH7/UqsqNtcoa9qH
2XoNqHK8LsNe2nqtPEyqi62J1RJGwHkE3VXSUBGnVoBtbw+1LaGWT0efOD6whYj6
XPpcwjXShl4fP4qxgRvrFiz0Bf0izXnUt6VfeH0ht8w3fE+8498hnOqcOxl4bjYk
9/AkCLDlYT+LVCETqeq+flAbQw8mUJl9o/Qm0AZyO2DNv0M3Sy2KUOaAFaSVkopj
9xPwQjz05oy10vE70G/PV+Pj4yJSJMDduyGEeI4QVR6TFx48jzU2+3atWI+sWD68
SRLm27uye44EdDIEci6ZDSv8x79cGj+hzeBgeG9osFE7L16BhmuEAskIDNVpV/lZ
OH+BNoDGLBPrWke84dcdtsn3WoPAM5IKrgBkD+t/eQ8heEjYlQJxKIpNDhtnPAHL
Pv6o0zOd1xHDceGiy3PQCX4rEpDimSHjLdnvgPYHc4ST/97wKNeWt8t2re4CyddE
VbN6Isu8+215JEhQww9bes4IDfX4yZNQEq6bKTxCnqsikbiXAMllhlsMIiZaDI7L
1EtzHo2Ceth9nxiGfeWUOX3QRb8K9ak6juj/nuavaG7QuZqp3uCrVHcl14XbpxPa
cRLIu2QMyfuElzbCc1nf/oMh5ep0iBaaQlWKmza7hiYGj4DaeWd89xWHQK3K/796
PA7LRqcnl4hHXTEHnHhPb417mhuytZUt0Mv0GvXHmTCb0qq1kpK+PCihitYFWfiL
gWWU4LoUEsPfxeVedmt3aURZQeEyx3RWvCeVLbQTGA/eDiAVFWDJwq5DaiEOuPXU
1kO80s12gwuSVFFZRMXFE8l5r0hMs5ebTfmACRbGQt6SK6p/sSlHMBB+b/TDs96D
wlsHmq2HHiLNM9c1eu20uQQrG5k+a+6sUPkbn7fjBDdAUtbUoJBOF5yokWhwUt23
hRU8IOu5b16INj+uRfkg/X3l2oRY0u9Axz9gfe9jWksW0wuA9CZbcSak/lO+M0IV
+F4dErLH/lWtktk77/AtvJx6qNeUUItC1KhAuvKF8qTzrni+Bdx567xoVO+Kj2UN
t+qsubOnDLmoClQp7wpglI6j/e06TkfyF3fMl4io4UL0S2NPx2aFUF77rBJ78zW4
OKbI+nQRZv6ioBMGRYNLFcLbeJ2g3U2yUCAt58Mr2nrap+LLTPaNQwPv/H91WnwT
R56vNHahRsBnB8h6Lt81/QfnZQ2Ibi/wb3V7+hHvvjETiXlmV3uKlcGTHoNhSTHB
CNTvz9nz6ZN+usR5N2XZ5tgxO/ATpJL+YKMFXdM+NHNp8ABF5HdoRiZS/rVABuWb
wteM3FmwCWcBqVcbVkB7aGYCqZIVHh6RJ93e1qDbpoAs2XXeQIEhww8J/7sDJ3Jd
5m3Mn5+MRhdXCY9AedIGPpTFIl4ejfwdHfTtk40F1YuMYJO6tXPQOEjioMs1nutX
GMwltYHJOgXuCD+pNEFXBv7GMK5qdxdjfJkcTfYKvC3Eg9Hl0FIpVtX9QzdEkU5v
RFhUhCGD/YNgO+IzFSXuPeO+2tHoNzhb4wSHyeSJXOPVh6EaZy0pXalWkwJ0n/sM
2Fj9OI7dT2e6eZIPCuZ7fgr98OiJSbw8FckGz5brITCYIGil9S0DWw03rf82lfXl
EQJRPKa3QbSwSrWuyX6p6B28KgrP0l5AI42jQIW4ZjuFYYIm5dZQVIWMVMcIM3S4
GQ+6vauR4mh4joVQU0x8bdInSZb93tF58QNPSykUxF8CNVoBouztZm7HmcCu6LbW
OEJKvbTFq6awqIKU/LPg5UJpTSRAcojUJ9y5laUIsJgzs+CUhGx6e+Cv8enHG6uE
pkIH7ZS8RTewlGqGVEHfj87E4FyF3DsXsk34sMZJhNOUrnU6xRtD6WglD2GnBGLH
cfcY9IHcS0yWy843NdhSeYcECgwn4CBAfcj+h7THD+9oBbeceq2cEQaQAE/UdK8F
8E8VX6JGnOGYYs4oIOni5AEoq7NveeMAawjuAJk98/VNkfplkOVoVH+PYKdDJDVw
mXDvD82tIprobVkiDFMmytlxgUHgl15rq/1DjEuMC6V7POiTVbI+KuWr0B5XXDXi
ZhiW+NZoYcpUEEA/Iul1sFHWm0ivbRZukLpZKJMuKmFev0Kn+OrC7l4p7ySoCqtm
/iR1UeXGIIrDwqmyRZFg1kbblXyTsGgt1BUpgEj2afMslT7NYy038aWhiDTtXoUo
LXMsAt5n0Uo//nAzOMV1dcmQrU8F7O9G/u+oqVfO5q45XpkPZjaA3Y/iko9SK/Wh
2OCf1AFMacvGATsNL6I0dz4Q/Csf+Hl/KGagYHmWwXSC2tShoLQbnBsTIVAd3A5N
Uw5ec9MYTiDhn9hlleWqpUSxonaC5Kqarz8F/A28RavuoxWRdAM1TpevCRTyaHNa
ckiwJzw7+vhRR5H4R0A+e0AwJqAomsEcyghNpNdJgu5uVLL7FZUz6ba6lqt9o8Wk
tsBZu3NBbwrEixNbioQ9pYcn6o99r2hjpSTKAAjrNJSnhQ6QNOfVVWUkzV43h5xG
IkQDqCZwMTi5bMdxH2D4HJCMvMX1F0yA4xmFkl7Kl9Z+dDXoN1nex5Z3W6f1IXJ0
Pc0m1gNY5lpQB2TNErSK4RNlrQ/HOw9LAAw7XL2ZzqPfhICoo8WCd7Ai+sbWdXhX
qbimfjp2rigYn41A7UX8qv9bUmpWS2qYtUPoz2aEa7fMsYppLd5Z6mIip1SCYNHY
sCofNn6S8F3lteWdMsUQYeK6ebfdqAo38nqOkzudr/SgyCx3KvwZdoczq7MQi4WA
F67oL4ZSUJy+DXOl6kQmZcJDkx7XXUAPwiy+ucs7FABm1Zv9iWxbwOH9liYrn3v0
0LgP6qO7wCNPCirgnOfCM4ppln4ftkDJATwp673BfHN0Qvt8emLZIlryZGyMmzAo
nCDfPX+GhpGt1cIQtnpmIZKPZ+D2aw4DivJhi5UZiau7hGAmldGdS1ssCN98zq3O
lYNADMfX2AbECPGjjv5JCVaxaBjUbqyc9Bvo89lRKzatIqcjXG5cad18aQgT51XW
l5k6vS00fduSSUwhCUuUAdWrVGb57/89QN7KTHkZVg0EqckG1dpc1ygTlTds69Ki
kGBmWpeaJxYrOyskIwaxYeX3XnI/Ou+rDu7cCDfT8bfbm4eZrDmmKabNE+rVDRqd
VNRyFRYdF/7Pgw0eVqdjsXIAI4sPQWYvqt3qH8Y0SjIKpr9fcv8zFRRUcs6+yjxM
BblxhzkQT5aMhnBgwWSlJ+AHoFHVZGhHWu3JWLD7WOttkicAqwzAjPWtXMwpTYqd
KX0atANcoAJoCMCsIwjbu3n2x9lMcqpoBZ8BtbTETDQn2PQdXFozly0ixeUJ/0iL
gGFKBABWrKmyRvPITD6gwyna3yJHgUpfeHy4TE8SmRJWOINagGs4oYlq9vcev4zS
DlyK04rwABDlPX/b9EjlJGRRb91Msm4Kvzon6e6HNeoSel38ySmPIw117gW3JKi0
JLvqM8Re0jJc31NR4SK9ZuvDtDObQDoV7XhEBOBjJr9KYEGo+0O17neN0Eo0uVhv
Y+W4zMSGeeMHGS7jBqyvCYwxtFELiiSozx9bWIbNrntMUPnJt1BK30fUOSO2qu0r
s0IystUFUuNFipjZKcLXWvyfNK3/4fiwjIUt0F6YjD5yfFTY/wS50Nng4GxMEz8s
EJTum9/Bx3fE6HxzMFCfLftTUXfQxmEQ8rBar1dZKVDrs84iyf/tYmWDHWrIAqNf
lXlMGduThurvo0xZsSMccpIsfsZrayw7oJiffEccNIHE8ZsUewIAhIFoeUufmjel
gdMe4wMtMMyoDl0KtRtDMumKwTC0ir7G5xFN404yqKeymb6l+tD9vVI3q52CGKjq
QD+f7RXxWjvEvF000SbCUdc0o1cV1J21SaIP/ZQS6PZQwSt0pTMBOLK2dLvblm9L
1yEnz2jFYioXRjbkREZiqdxf/69PV55StHzlVsyRlvbrFoLXgUwGdqrP0DmDo4rk
wHihiJMcdgG3IQvh3p+Q2EzMyjHrQrUO8m88T+Eer8etBBXVSBLPqaZEKKgDowsa
7Q1lXrSob/WhbfKQAs8E+Uo3l+fgf4/NyFTHxfsovsJsm5sp7KY9UK1Hma7iq1M3
MQgnl7APthv0eAGWON9vPFc83yJki1HyiF4DQ+UV8grrI1KyTRgxG2bFvVf0M9fn
15rQe2uCWBA3v3S1qhWe16j6NyLApvbFXlfDXaCWVQfPdc3Y9fJEzShou+9D3ap5
fpsPAcFPV6XKpn1rDYEAK689g26vQC5w8uncnp4mkShZ8jdpTxHSFc2ts0eeichC
A9bG1obrVREix6j+J/hli2seRuVnhSFWrZOD4TgKFtuLIKgz96GgG2JWoekq9HhP
1e/IAqW6vpbFfohvw3RkHC26O4LRx1NNWNlxDt/REczJc7KrdLFMK02MkjylOJRZ
BL7OGGZgGegjHHBnVkpFJ/pdetGTvz8nfL8Xl5KVjFVJi0lC+OesByhLIZNcl4Ul
vmrJWm9++8gcBCSqGBkGJ3FYo3Ezy+Nh2WO4p77Bi1TZPgg6X5jfhGaGqNMr52nR
SsPbPAXny8SCQffhxKN0RcbQ06UB2XHAG0s74HLu7bfpFb3ozzaLEH2PdprQD/VG
3i7+7kXXNcQsPjZfZQzyBsEu86h0jFWn8RKeiZkD+52GEa1BSsWuy735y+alF2G4
g39tfcRRHEFBMsjwUYtpsrnRKm3CM6vG2XSKlYnAY3yPi2y69wI2Futo9A+tsWA1
33zTZbdMRJCUC4JhOdp/NPbKKYffoWeVd+LKd/rbh9Qk4xM7oaa61yiqfyNspg6T
f4BjFDk8b+vMLdt7ndHqNr/bwveUHblz4FtGLKX8R9fixBiROBnDtaEaSkkQGd9c
CCNaSzrxX2ByPgLwCsHXlvtje7aVr6qDlKVgPayXaUrrfXdS5+Ft50O4OjM456eZ
rCpWC00JAgUcPt0jAJA2AOaIjuaxVypIScctUCkcPdCxzySlMw1QxGdOpMQGJPqw
y6kkNC9ixGfra89QsFwVVh4xjQ2es1+nXBpEG4wD7MJHiT6qNM74HS0ImNAlNslT
CRpkwz1fPaC+ZkuKG8yigLyti9XhfuA1t5bNSa5pH3dUkdNGfDLlSO6eRnNtNCnw
t0Jj3GOgnrfcgyc48lZmvp9nGlUK5xzgluSg+BvmGHjSnq2c5dFTLzdc0RoCChR0
Xh+U2BCfZN3R1xyHRJO0yDLhtUS4Orp049H8S+3D7wxR8Vj880t4riXFj4PVMjWF

//pragma protect end_data_block
//pragma protect digest_block
lZhEsQqRAY8rQlC3QM+KpTPi+qU=
//pragma protect end_digest_block
//pragma protect end_protected
