// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Hp8PYrTVRQxPq73JE+K1BRpmsztY6uwLI0OakbDFccTfYS/n4i41xYfsI/+a
qe266YUQ+Ic3A8TxfvriqsrYhT/19gpr3TOvBl5ceubXAg0aAvHsbSF6Yk7O
yuT4N8SjBnn8jBqQ5EGQHApiXfaYNbJ3Pqh+LoltSow4bVligI1RfyMzLPc+
6hUQBxLu5+2rmHzSO5YVUCEDNG+DZsEHofknCc77eNrhaJ9HSTTkpwpvts4F
9Yj81afyCaWtJI77t8yNqkv1f4ltQ4FnU7Yca2yHWz8rn9FB9ie0E1IKhJoC
UqP0g765FYliqH7LAakqIjv5MEtv1qWQVfylncfs5w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h145JycSHbIc7lQJ90vtGBhV7nrgSgnugjsFeSrIJMisj12j2MXq/UBv6rAg
czZwxqD6AqN8E4pqPlwi86BOxAT8sDPR95RHO8RiHro+wyrxeydXL8H0KFfF
9aWLfIOkIICqhQRsL8DcCRceum8XFlZrXvLO9AGuQp7SxnL44e/SWdJpAQUG
KJL+EItwaVWc+Trx0Z8X1MCoxtPqpyxM8lhFMjFM9alX7kt+c2gsFESmWMRV
V10mpliStqmifBL4FifDMc+WfNSoonld0YIngfWs2/m4i685VGhO73O2mAym
JUzYIt1YRvJNlWyYpcl6r/6tOsRM1R5JfiFD8X8znQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XLCQc8iIxaVWxfkSJ34WzBWSuIyZLT1Krc75zQAQt7Cd4NO6c4Dq6U5ZxpTy
xnQvxbIetdwPEOssX+xoDwWJ+0LyYFWQXMLZoB55Im7oGJejJDJBp9fq4t5x
wDRiLibn1EFQyrpnzfvDi0wYdCgeIe/EOP0p4qqPBoa5DLUsutwPOw6YL1tq
WhlemhDdy37mXYgCrvt2kSxtb3s6t3qColMm/HYstmHH8cPcbeVN69UjYQPJ
qbYJl3NFiHwJaK+1I/TmFYm1hdWDwHVIsv3PrGSuGFnfMm1gbq8uuvwkHURi
NCRegjkCML52meLZUfTMELPj4k1Z/4ALKHUTkBqMtA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h+w9JRE5JEXjcbIw5+FXD0cYbH4W55pQYE53Pz7e7UdFnZYMtwIQynDqEiMu
58taIS4hakze0OLHAHmKEVTFcKBZDiSmtJapeLTG1hQtdCf+QMh89e7wIly6
Q7+v11a7qq3BGMdDVhHGKKwni/Ir8/FpcHwIcCrKOSxJTaK02NA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
dqMs/i6cpL1nJRMiMZENvU35N4eXuFQtbqdH/B/Ql4WcJfUUXdXhW4sanyQv
ivF86HdAMvhlkXvYEYIBDKGgFCU2GHyALc+lWQXJQ7TAVGaQt83KbSU0hR20
x3rRt3gEtgBDDX5CCTJvRR9w7wsE4DqQ9NVb1vZ1OZcOwLjq+AF4rOgnRxEl
jUZ9+fS97JPP3xQRdg5akB75PuLLqeT4syEHvdiok0KwzG0Ga+CQFYvAuv+O
P/dFFClK73gL8ICJzvMxsB/isG9E4C5fKXU/Rn1C+vFFmynJPeRtyXrhthBf
KdrqsanE7RG3HZ0IR651ZwF2z5irolgzh3U0xMndxA84uHmBsqpX5dswbgqA
yYxKvgKIVQC+xgyh5g2JOWeJjVWteSURMxnQDt8pno2H4VW9NRe2dlUODSw3
Ey0tNY0lPRWLovHWV5XlXlBVye6wBDXpYwvePbnyUtxBnUChnFNy7TT9N9qX
VxTzpV5okvCVr7bDoDm3jEYvuZ8SCfOc


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uBnWsO7Ynevj51PoHG2E9iAA4Am00uypMu2EAcnnGja8sG/zbLDqKRdyUVzp
8ykbBjz+7VX9kNeQi61G4nZFwa2dmveDQITOlP9J7WOZO2ZQ7VXLITm7Rq9q
XuTSZfnNfjxVtXpBJSdZKQXvy7IXRLw1qaw+xEIPaPBJEE3/SIc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Pxrkrx5FvXiIeUO3+ODiuSI5buPYttrlIHAG41eCLbGmjRPmuC5CKnWUFcf6
6HyeDKB7Es7dDp2tkLv1Z9u0yHTCZXOld/mQcb0aGno7GxInOUrk97lZrdJe
DqxQQJxy17MIIRGLzpF9Nr+PUWJ7dfcpdawRGKWEAg7/b03L+ZY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 44048)
`pragma protect data_block
0c5880eBpSnmIFkWYsRKFBETBzMlBTzg/CK9BxrLvtiUxyUxPzTjWnB7SQHG
lJ2AP1n83E/VaZghwp4kHkybcHGN3sIFu1kfOIKU+vblI7jgGsMPfcd6oEcF
NemFxB81m4qGo5IP1g6KS5TY60BpOsOyHM0T36+t09h3WjTQ5D+aDxXR5R2k
BoQ0mxF0Msibe/f/F/ETTucYN+YyWdd0/3Mk1tktjwdN8MLrn7i4nKVj7D7i
qBus8JS80/V8KUozEH3S5qEzVwN54NFCbUVB5rYmpeCqHosHPVk54ikkzcVz
lD26FGF/rDZ+ktnUWkReY9YPraU4iuhEEmi2XdLKAZmAh25ShjHMqo8N5mWH
wUHWH1WAda6NiSNCPdvGuQinZunakeup9UlyLj8es1mIeVdYNBAwOfC4I2By
cweoCiHZ7oNHK9bnKbwM+iRCByEYVDhws4GIfDSIYXvQlG+RTlD63c7c5hIB
eULHiOdJRQeLTQIBfyg0vHFExFNFPlqtwsSwUAjSI9SFHK5ACrkHFTbalrvF
D9Vqen9SXqIlU2QWsW94go9iJ1vALFQqmSC5OLmLQAl/RkzfTPmwCKnb7/07
RTULtEkJPIbrdArnvjVJ7eOqwLQoPgwWg/NdeVV0RrR3JPnUC2wdJ5AsHJwq
9cfKVqk2mNzJ770GJnZeVITTVCx4Mx8bjYpUnDAuRR0fSYIYSPShaMz7rxvd
21PC7ia5u1aV5zOtbzTixVa8/t3aAu+gytC/igZtEWW+g1GdA67vPTuIGecp
Id0Y2PcyUxMw/1czMJAanWREnRxEubGVSCEh+xnh9fP91J27H+p2/VBtdXvB
3DK+iQqxjqvE6Mo5T+zvVN9F6XYZ9Mvbj0VHRu9rqUz6nrb1g7qkAP1/uAkV
c8ef/pY4vnMvLrq7S/LMSdzPbM7K0wDkSmJ53H8EhJkvMSIIobNNWfxfHMAq
Zu6I7YnybkN85OFLIIBnW3Mjmtl2b7Pl6tKBbb5qvQjbAwAvBeyTHiWWBRq3
k9Hvfrz3lEWpULU+/pxsZb96e+67yNAAMr1PZrPGbfkbWnSC1Cp9oPhTh0Wr
eSmaXPd2MGjcKrtgaN1Y4YNhxr0qnx9zqXoySgD1sech3pzmP9adLcLk8Ua8
E4OUhK9gafzkeqfTEsK3SBWbvYvD0c/4M9xk7PGqGu8Hl8LJIGFYbWZqM92D
xfbl56udBkammxGZz6NXu+BpeOs+kzL2MKsMQntNBZ0ZcynsBmFpt6wtyM9b
8wUmnHKfrcWL0/nbf80wC2O7URjML6SQp+jnVy4CkU71ZAIUUsoFi+T0tdLV
4ndmZoF6UdkHeNRLsTEVjxVIEF+WWzieNWmEp0eugG9cHPHR+/ynGtEJsJVO
042++e9DM36OSvPiTA8/0vD0f4nAwxS/B2I9H2IDRTF8j6AsMXxzPmQxK5rF
yCEeTEJs1CR46Y63cnv48Kt/zf59oOYXU9sCjmLNnuWtxA8Ot9mwKibIXVq9
XWZK1FaSiv4+B7e+QfMC7vBXBZwaBiOQlUHsCq3gClK3/VH9zUEx2a5NkvVY
8o//WIlASf1L2VKUHYQWMhc7Hg+LcPhcxmyZUEXsKqlEqo5YqF+YLCMSYCOe
FfuEH3Ny266aso2k6czT52cGOEEAA9m46IBBdHPDRR2AQhSZkZ4iUdtlOrkD
wQZTnjAoXpllo3F9GiOZchs8A5/6rebEQG6vrH+H85xFrakXKEsZzCgY4z4x
LLxhPqtNGqa1Ch8XeN8aYfmOEtAKE3vCLL7m5UuUE6hfpH8bMLEYAJwGaFZc
14Ji+hZlT8rOTJJa+zGf54HR4RmUxNZn7z8DdML0N5roL2D+K5kbL/sI/P7m
J10XPd+wRfrbvfD1lS0AD+Wn8u4ZUO3f/ZEibUGTtxkjmr1tXq/M3tcsvyNm
/5IgCeDc177TMNgBgiZYO9aHHK6W6D2LGeqda2gI3ld+Uc+o/yvtkZTs3OlQ
WAuhHfxL/G3dfco6c37IWPHOeh5uaxMOUXFhE0FMfAbKzcg8UMvL3xK6vDU6
M7lGNP40XmnDmtTLsHdBhoFuFbbZJRexEopI7e/67DKm3efSpbfU6ODcQy1K
V6aKaDJPxVzxTsUuqmMwkEGSzUijiiPkfB/HDLLlwQlJKtj6C7rrEo5tIc9H
7U1bTvgJ7uDJXENxwXI5PP1SjEF7DkMtZXETTimfj6DCL2ajzXvcelMgtaLi
S8ST6F+ppUYfPWkJNfL65113lSBMf0hafXD8a95nsz+nmf35yvb4eshrYsCN
F/xhI4MBA7kC5VHXEOZuPP5NauHSqaoP5jDtlQsbWRZe9EHvZZD5uqqZq5jE
I55YtoDPBVqegYoNKAbUvFGN3CMXSnnuKv6UqN/gS0MBFtQ+ydLBW9Vt1I8p
3ZvoeFaaXfES83QYk2hT2zhcC2j3RpiBcPE0Mqp3U8SBS1ZWatHZ5Ep5Pk8A
5MoUBE5O2uQLs4h8s1PvMX25yYEnewQuya/zvNj3kWlrHAJpBt/IC9VNazUk
C1g+NhMv+eTvY/Zofz6SQXu/HVisjrMChxIkF8VO3FVN+F3bG3I45nJPyh+/
RO6bnoLUM7DLnsdxuMRVxKrGKcCmOvV+nQEa0K+Ym/q6rp9v5FE6iCWhilnB
wIUKUEilaUPaNMucFummpGFFOYbD7YrSbTGOjcY+NU5ND5jsZG24ZL9I6giJ
IjiGH7+8mjjmXWC8MGe15IYTpCGufGPA6O/OCJwYoVfzX/qZwd2D6Xqbb0Ib
a3GdU5dXMrnSInWejbZZr1dW+P4CXt1qF2WoBa634TVvM2+lLOtGs8T1RDgV
qz5G8uPGwBDKOoYyelNS1MfWy+1845Yl53rFCHUVYbotJ0Ow2a2WdSq9KEUi
YDMeLOOSdNjb/RXW72ZkhgTHcGVzLmw2moQdFOt5m/qK83/WDJPq6byJpxTr
LTzWDssyY/nNswFWALJOHvvBzaeNFSqFujeQmFGnrku8Zuy8Eanr6Y2tqT7T
cl4Ux5tqqCxveLSCIKCaSeFI6dJjOVsAm4VZ5QlplI0KJ5EDIaFSR99goffl
Umchw1SUnFeeguFq+pD9n/CWzkr4O1wzmq/22QyqhzSbchHfeBtIDSIoWMwO
W7puIkaZyAKNCWjmi0ZyQT/b9hwpiALggeSmOwEhvkMzlBob6STjsY+SBfcC
xMqBCQZhqq6ZPl9BGCchvUgoqpkSR4Bt2LSNE5v+hovDx0hz/trQdSsE3The
WsS1ZaURQk/ucqxzlCKfQTvYwLKv/CA9vSctsL3OIynbxNAoPNX3tmkdhxEd
eNgtaJm5rayXdiHcDuYmvFfbVqJvxValhpbDAvUiKIE2YB7ARbC6Y4mqILru
gulcWt9aV19Pd+AGaaR6hsr7LPXUwnxi4/yxMZdZVWm6Pi3h+Sn9D32zSkhC
3d1xYBbYkna57P4RkuGqJDrNcm3kh2a7HgFpIPTVwKTbFsPBQiC0yM/U09Y/
2V9PKd8euBprV1kyaVGg/uNQjqHtMZ2m5IqoTUGzrD39xzl0bMArDI7oOJvi
gsSZQpcUdEEvdbfmfla5XLva0lhBEDHzX0p5Ina9hPbjoz6dzTbg4Bi8cQZ7
XJifqF3hOjhB4VcEosxKQ5piY9HXwdkiQZMEeWCO1H21XE/P/xIldXQNcvDH
iUbPj7wLGPk+LRGInRtC7qx2Q4NQ7wOZRKEklHsk+6uVEpq/iTEZKOX+7l98
CRhyGIK7akNpJj9IFmij3PX0eGGkpc6drWmllcrH/ig15Bg0+pWgFnJWX2g2
ZGkJl2WpjDcmiHnKtLyNUuL+LvQbYBHFTFCnWBL+0kT7Kqyddpasumvf2Cal
eqvp17clUmQxKO8JYi8VVBepbOs2aSMxDix0SN/fiwb3JAayRux6JK4Dr5/3
QnMHaOglrO/ezszQ+PIznaM8vh2VlOTkMwxTPY5294ntVnUlNYCLI/7o/smU
gZLD19jkoEm/q7zlcyefzJs6KVu2JAfxPSrLWEDCpxuPWcgmCoqoP2KH0Muj
mdBiyaCEgLXF/r4LGVhJE3DZu8ZpEXSBUqoWKfnbb/BJi3CSKqiGvwT1wOqO
xwHfbzg6JzOdlOFlKYeml6jK1g5Ah2yTaE34hb9/yfaQQ6VrbsQDHg/x58MP
1FvW1uQPxSHTRwMkC+LA6cGE/pvMGJQr4En1WpGtjd8b9fglMvjTIrDQAaRD
5IKhijfezXRZsmka6jAw4B+CqW0y+mL6EK1SvTGDDBW+VSs//MU7Lxl3ixyB
1wjzK9hjmcnmG7zbx4f6iF36j/yS2WgL5i800V1VYbbFi9RK1+BUAdaEuGtr
fDTfWJGxBk6E4vPci3dlU6uoYRsKEvvXlLuZDDr9pw1YEmFa6DF4K9YrczkR
X6el7kMwjSi6yRYiK1cYQL3na8FfYEDSLGy1PR/83SwsAwlAq8A8QW0cYMgB
IqSfYcFjTRHoU6dMdynqRywYwiPvsVlEvnNYqgCHCVJOO9WMAoYIRcv5LCzd
vWBcwPogUTGJjlbcwVwwZKEZ1YSsg2JcnMi73zqP2eIQOJ8tJ2Gywi//S+2S
2O7+U7sU/yH6hn7uFWilDdga+BFoFMAJxL5dhF/6ia1VQun+gXLqB2RaE36v
/LXDTuSv3yt+3ZnEC5EcEq/NX+bo1E/tXt3O6tP+T8wjZpDrbT9A03okEFH7
QOEtMWdFYuoPPMMSN8ea/nkgV7Oqmv/wcM98sRCq2cCBBAWh0MR3iODHB71l
YeQ8x9DWLqDcxCXDcVDKnbAVLXHMbFYnVFTqZ+Yh1pdIaHIlQ90vZdGXyerM
U2KcPnu49MEnBqjJExb7WN4Y8Xs+jYYu6V+4Fh7dTpl8uY84Nj3NCbpr1qVM
siCKhN7gQ8w6dZtJmjzARyjtxjhxtosQLyl2yErxdkW3Iv6un3gyMprfS0Pt
YoQu6zj0DE3FdG/aLvnxKPhJICnFASJvdHCAtasXD1HiSVZp04bdUzge7ADX
cOkYUjsq1bWkknP/AgO/cpp5Oum5Au5zFmNmWSqx+zaoXA7d81E/Fkp3h+Ie
qJIL7+TvMboT2mIC2nDgUxdzaYP0T8Bqa1QhEkK+mMOpRZH3crAN3dzMCf9V
cguZoMW0ZZnZvl2AcUvd9fY/rk6T0yaLAv3eGbl8z4U/iP4E/O0sptMIYawp
Wk3ERV68V6NcMZYoVsRSjl7L1//mDpQkGQwyRm9QAvnEsT2udTNWRv2jOSBC
2LdaGbwffF02miefzykE+344tJFWX6YhlKZ8Lm0lWcCGJYagJf9jj64RBD+G
SzLK3RGC+ww59QJTBWHbsYDcDB0tNou0OVFOax4+NPL15p6U+L/dEQAEvHfQ
HhvXexH2i4f4KMVqVNGh3lCZpPgRZTVYuYYwwLa0RwwjR745E4ZGQDafXZ7y
KeiOG3waeW0V5r+SnJFQEzrQJB2xKEPlE3ehGc2wVb4mYHWcq/gOQwp3skgK
anrFWTw0qk15AinLlI22cA1jAFSkjttaFNk7ChvocYE2TiJef6GXCjmjxnv8
EM7lqNJPyr9c/wtlNS7oda63vqqUBzTwYgbIjZ4QYQvbTfWJLXs1+rbw3otM
7JbOthkAEbiD/WByjYHsKuqtzOIU9/Om0ZzzfjH2penOVaj1pkTJMdNzTaxZ
utemzC9hi5OHmyqMKjDJzaYL2QXmeLNnzIFMMfAhuYbJUttQTppaMo/Z3uId
myIc2zhLG94Wap/NjGDvRngd7aabb8DxtBjdJp/x/rBxfT1gGctNItrtwqP1
/k46TNSsKQH4EVCxWeE8kknpFGuJFSS4l52xTdh/7KJREW4sUAzcEZdmCFMf
BSCTH7w0m6xrIvwoyb7qDhl49vDdqhpeF9pjxoK5WLESl2sRn3CmZY2txKkw
ypZW3MTvQPtlqKpvhmGUiNqBB8MJTBPrJFETFsemdiutoUHQhGb2yW7ZhZNo
wL/XnIpRzTA0S6QvpKKDTJGxVwlsLMp0t5haTKiosbD4eRfBPLWz2K/E6YEx
gIh0iK/DLgp3hFdb1txuL3bwH0tgFddeFORppQsBZKXNiLaZJbCMzzXU+49/
tTEmBsWgTjIka9o/89WHRQfZsJewLhIIcnLt7kqtsMtyZipk8ftjsoIV1jsE
BZZKG3yrnXjbwiV+lBMsOqwyKSXIXdL+gWkHj5cV91ztHv2AFU1F1PmEW/AL
pUZ/gzZ2G/OqMFTw/c9bC9JqjpqeN1tqSDMAzWCkYava0rVnXZegbIQWaXCO
T5tHjm0JM+DgqhiP5+0v8uTnvm3py5LOzEanJ3LaKRsrHG4Z+FQjl6qHMA1s
C7Qs+UR8XRQaS2XUsWlcSdpVwGXfnNf2CIcDFU4CcDPWNoQhUONFzdrABnD3
gQpZIC+xRWmppZRMa561EtDIWhEnge73bFuCTvtMGy3giE2zBlGCLPTrOWe8
ixEe2phITcRZzSbUe+PSAJvTb6e34q//ncV/eawdy9An67x8UeFv9vflhAfh
EyViUY6shNqx2AkEo+4jXoxd0pliTfYZhiLnaicpFsAP3YoQbqBL7LsAhIUH
cvtqnjKjubNY20xvFTfon/Q/TIlFkD7nnPnL63UAqOQFtvFvFcdbYrHFx0Jl
uHphrFTYrZRA2vGSwFl2P0IGSHHSaEZN0g2Dh6e9I/EHjl9RP/7yoWVuTU5N
WM4k0JmGGKDevdVJm2sarOETDeNkq/OyO68rG1nm8LrLZ5Z767D8z+6GJNgM
Crkodk8HGjWciiV1Lpv7z57QrVO2XyazvoTpB7P9tC2CxaCMyrPUfPIzKcC7
bbpuMMdybVFLEF+yhesY0u+H17hm6WYdAt6PR5nL1X7bXn+PHvNsZlYqK3Ka
c171mMK+TGskIrHTON4ZUx723LTOmBml9QJ36T2iSrnuCN8uaVUZjHbW7dk4
luZ3rzHYPc9gTajAMncaHrXLc//NKazz86fLvKeq5M/ZGDUdHBHdB9ZJNJjN
akb9iA5MboLobSZCJDP0IzPzzLmgfXQ6pyduMM0S/0sHe9izOSgdZeq+PiiA
cqBMflfgtQC5NUC10/mWx2t4sBgJbXe5oz8W06KtRJSbf/RHjnMKs5Nx+s0F
EXgs6blTKYd4Qhc343eKWXSiRKovA4dpnx8gKAFBLnciT7CQCUf2Dxk3866h
rtCJQJZjat8lkmE4w5dpv3FtLmZ+ylST1ffDzvAOdwdaaVvzNQSNCtkT44/e
Q9MTb2s34f6suPWeQKIEc9QqPJMtpn/ha3eYmKQ5JbVbnae2SK1HjVnY+uov
2z+JBeQHsxrHomuybZapSzq69pznCZMpG15FJaVhD/QifgwxMk2vsM/aHPI0
CW0EuWOG2f+O4tX2ih6keUsQ5Wa5kwnDk9AEWEuDprgrVPzKetAmEUExbpVH
W6rJvNlD3vLty5SFHkh4zJow8/7ioljiUGaVkhp7mZ4kU6i2ifZD8oWmv9fi
Q8IJ6aL7530cm7pdqyClg2XK0ycZ9+NfjCSEcNfbE/zMci1OsrHtPjPJJmG0
CmU85gK/7AX7dvD5sqtj5u21EqUqA6z5tWmMFkRWWH6yZ1EXKn+r6RmKMHeP
1UppHcUHRWYltOu21TSlT/Ug76jcK9uTXKEBFUy6ynDB/7tl5yQ8La1E4GOG
bp5u7c5KBM6Si5jjQTBQnVNl1DJP27u1m4j7IX6+NrZwsXZe5A7MdP5l/wcI
/CIl5OIBvjD/z4hB9spq6VnBi4W3SpVCmLcsLTPcqLSn/SCkYYQgIAqi2qAl
KEyk2T6A72FTaLj7uokkpdEdGl/8bAY8yZaXR+J4o7aozu+SaM/CrFoKQLIF
kGHJEZLGNJ/6jxbgAY9sDe/vDmXqtrqRSIbXmDNqIWsijwL6HviQgbwO0un2
Fuc5QESEm6KVdnntkFJOE4QmF4YV/umzJg/SI21NoZNFUcYwzunxkmCrpt+Y
4N/hUD0BulTRs5GOOiGfwZs28M3AvvTt+lEJTP878jP0GrTcVh6sBVcaG47r
ua3L1G2b3+qxqUE7RGddsaASH4fLfzayQEq7XbBuDGTVKtqlgI7BTvor/HzB
aCgCP1BLNJ2afhOuUoA2z56S56Z9S4ayraY82Oa4B3MYuf7q2hkQBdBgmvYS
qK0hamOoLFWy1idN9RzN/PZlS15YQh524vwphAkrm+hwwjWEQrGixWL+HQMM
poHdsw1afFO4jT7j0LKwn0bwuaC+uNv207s/cIE0oX6RZY57zoFxi0XfHs2R
5cykmRlRErbq+/zafAW3VejdK4Q06rN4xCk2TmYWjbVzT3ez4tGed+jJAOHc
5j7aLZkxpYcXfDQbfObiuPsLkdr5H+k98mtOB2fMDKdds8hedCXkb9IwHacC
fyv7qesb1pyOzUJO16dOVVO0Aj+RsvRVloJe5wkpPMDpumAFii7qIm7Oo9O7
7uFrs4LcCePWMfzZooA0LlE2GBzlLZ2Z52K4CKD+s+ZXj3ioEShYmbksKhj1
1VNoGXyLHxQSXHwHRxqIgQwyHc5KeC3Xk3TAsQ+vXhgP/TO++EbZ/ADlW8ho
hbOONm9gsaHHXRgSH4qksksDmc+PAdUqsbrjUATIxclI9yu8qKng+6/QzeIh
DpBoRSWZS9J+BWb/ioMB24jbosSDp19t5RqMZ5FWY/SBDT6tGboapRBRHBS2
iYWARFceC6KT6gaSw3t/1KA4+TNRYa14//ePnodtFeKu83k4mypCodyrRCIZ
+oouMg2wvecBCpouzGaIbKjcqEhfD+qvLZ59OJGAwkstVrrFFt/J1iWZgT7g
Gd4QQxH2rf7/UrLdYcW2jdZLSrn0eNPwxfHfqjc27sHq3/1Z8lyPRi0Kf7DH
B32EVrh6t9zEqsqrWyviT3NX9qQ5Upnj5aJ/Z3N95dX1VvXyLVH0bWfL0n9I
KIhXhu9UVyPLgMcnLSr9OQV5lHeaxNBYK070n5Ih6OPcyQmJH1SVC/yH6G4t
GbOHMIn/w9d4ssI09QSwSQG7Yb3opLQOTdr6gk0l+wNXupcKPvpjK2lvW58x
haFK9hwUnZHXCziC4xFYUzVlkvxdNGBcji0UObiXTMoS3rWJgHsMkqgh3wgu
SpJ6T5LgWAzW2zSzdYj+aWW/jKuXekVqjxwGIn7T9MXhlcnJ+y+YuHgu7t8i
jK7OjGuQtGAu8NHmxQNypg9g7L1SkwrMg6aiW1wwzHJjWb0qRnVGh8jx5XB+
mcd+frSPevZb2sySoHKGAyXj+Bpg6NORxTsp+CzwtqYQkbx6G92ICRBST6YW
U6pjnPbnqFrKgonQyBwV/N5anq6IvHHRCu4DZzDgD69MubiGRkDsdrDAlkp/
gpZOiR4WDYXZQ7zlpK49oaVG6iAYaTkd63/wTdoYuS+xEt8RH9VZni6GSclv
GY59cM4q+4gBzaDCP2wwbxysYcK0dUmSqKQ9KcjAWTgF5MdGKtVoUxk+3K/b
+9YjhvoFN7P/O2KbzOCUWJqWqthKPJd88XaQL8dYuU6JqWYdMrg/W8EngWSL
J7sLGE3L2+tT21D7Nb6Su1ogy+JIHveljla6gFLNtuEN1AJVZFXvQ1hYFgWa
lVfG3M6y7ePR2GGmapSRjj9tLKW4ce1iYdpGmRYjRp3PomqcJM/vxxwoPxvV
8EVLH2Ux9yS4iX3g18E+LbXVU/pNL056vtgJLPyXvuzj53hCft4nZn5WSGn+
rq0u+9pzWYzN4N080kAi46YeWWiAQbzMrJVrKFfdfjattwgw2tENl5cGeY4/
/jDHtl5MkOgLmN21umHw1Wi8EgcjS45LTq14EUmwB6ehueMeXIFHvRwG+XSt
PACuBcD0Jcdg2KNokwDxlf8chYARHKa4P+uMIv8I30JJK291lFTSowS07ckS
tirMv/rFvkciar27oZUiAFrHQRWgpVNHzzL6kItuOu0kG79cnIFyMlz4muha
4olcdNP/lOZ9VbVF9XojUUfhdjZNZHFHpRbYpsYs2AmUGjE/vvUXkZ0MHIfh
DTNOwibiQIaUfq8jP7+8mYSv2LixYHlBbjibF1+zK3Y5pjXqck5d2hVpdfjh
kvPuKwWCzjo++1f8WT4TwZ8oj0e9CUtlRe9xhTwdqbLh1CCdHI3Qzd6udN9E
6se1oVL1aseccq8PEqsGkEIQnW/n7sh9JpAUTR2XCe0MXbEtOdzD5HLSrCDY
1nBufIE9YM1Fsy+vt92DEZDcrX8G3geFogUBuhT5yJuAhKXpBcNAe6F2x24d
Nobsk1Qo9OfO977HZTtHDRQIIQCU6HSDyzC/fOXM5licmi7RMZIgTjCk/y+y
TvLRercQI/3DQ3NTgrQtjcKL2xDY9N0QxjYF+LyRQillD/lEh7AAcdSQ0B4B
mXZquD4JoaP5ZpPtt1QSg72jsh1phWVUoiCCU9iF6VMTX2eQYpVk/wdBG6f2
X1G/4Yp4kjZNua/8BzdZCUaRHYWwQl9axAqQ7/1Iz3yqCa48SzvQfMAew1Jr
z4rgt1xnmFPhGP3HDIP7d2eXkz8e7z4WTsVSGQjQDCGdh0r7JBJ07MgVOuag
Ygpq1v7lj09jiYPL8HG05mPlpWcUdPWlcCrYV4itnDMbzusS4tBRkKB8fTCb
AUQmCtI+MLBv/Hswo8zvz0w4Tz8rW74dAcRPxDh0ATKPQB2Ug1826p6X9jwe
C6oqsq6BPKJZAsf3cf9hSCd24wbAJntPR/vCFr70pVDxLD6iDRNeRaUwl6yP
VjuaXRe3lHMZq8NlnvmHR73R8KJzpro4ArH5huqut8SwsTCuYHgfkxDvte5/
Y1BYgxgTDM1C7ajJyFrfbh+ya2txCaT5D6F+JA+iUN3K+jN6IiDD0Qr8NpLT
yM1sQ4P20IazDYHcVV+k0HSUFtWJTdQre+e7Ul54VIpXupdGXlTpidE75hVy
83QUas9E6rsOioJiHDRRYmlMBQK2iaSH7Sg87gZQBThXqixx9GToh9SUbTr/
W9BM2YS3c6YjpCYqYbwMX2FrgC/B/nE8TZvHMBmakHs9ORoDtWvCzpnzB9IG
wbsNNEL0Nxk0jAbwkkmjN5CdPxLC1u8VN33Gh5Qku2aTTkldTFBHlnQmKaOW
L3RS7DiBSvbxt7atBT4wJWVhItBCEKanaOmRJF798BGcnqM2oQWF3ixlC2rV
pzfzisHJpSEN0BgVwo09Y2Q1jxPc09SvOyd+9HRq7YpyVo9/x5mfTfJuzEM0
P4LpH8uJ/lOx2YLO66fAten7axHwUplEnDa8thmiCM/NnKyInw/gqttnoq2E
SP7n8kD2EN9ObJCamOI74HhBylk9j6aiHYJYLrmBw7FNxPN1tS5rhzdd6Ea4
bRu62uC2ag7y4lN5oacvGSddw3qqKxoyVxUyqBgPwYCuyFikNBAxhz+iYuj0
AmsgivJekTLiY0wXfiPueuyOnD6nwy72tP/9LkCMTz8iDrtXIEw+vZN+S6MN
nksSKN4AHuMr0406TXUYW98XisbWLfzsOr1p53ML9CLQi3CtOQPirsJ4/Qrv
dqkh4/0k4k+5V7KL1tLpQKKa+WFpI34dUm2uJ37GhxE/E8K8qIs40NaM+lUE
XJzjNd9NXNTj16QEhoh1HJlTRFbct+TcOTy8TyGTFKcIf7BJ+Kdgo89vV8jf
xABEsVyL/JvZTU5/o4kvSTBbfHWDyVI4ndWIDAAhDf/RrGm91GVjmTInjeoV
BTR0Oi1DSyTo3jAt55vn1ORLu8qnyunKJUorB/V2iPqEE9ypX8LNjix66flG
X1XcA34mzscZu9IvNViBMjxUxLGwX5sACN2wAZWwVA8YagkfuKcpabvRLUtu
oX/vl/g8tKs/iZeDVclvfIlnRamizxAMNSV+bGGC8yZSvr/b35wd3tx+Dv3G
cNvToKHUIvXcV5qrs9IQSf/B+zi7edeID1uJOMkpjofhN1yMTjSFgAbZoPp0
I/Zllq1apPYrYx1Tm4sD+SrEfgFaS+y10d1rGGxzrMyJPNbUzavI7hP0zCBl
wjC79YCK2GzbXDrmXUSiCgPNfu1p2Oc+bSSCxzvvfsh99UByh0nLCTcom2nX
BKrS2kR3KYV4VxRJUVfSWWqBlG/w12p4OHHX5sPdLFr23Ha2tWKKosewh9my
I0AB9dY7M27MZ5JPtShwvSHBJVMJpueZ31SqBaueYFLEjYtW8sIS7r3HdF0/
VbTkY4T+Z/YoUd9xEdXlDA2tsX5PNx/aYZ8zxVV+oYjEV9IFIjlTuAnPFgI/
EJ5iPkre9wbAJEC+QdFGZSNZtPDMbSvcCWkQllqzcSnHGa+9T+XfrjZaZrvz
4dv8EZFvFYRmyJxj39y4hmQbxmMU011yJUB+SV73O2HHzV8xUY2FU+n+CM7T
BWBuK1gZ7HFytdKOrQYN4jWv2ruGUAOACSLEtmwpNNBeqOOnVV33dy4DQXfS
IY/rWSj+7RIy3+TRAZfrgNsvuPaKOE2N+SP+dM/ojpishlD0qWoidSBqeUmy
FUSyaCG8Y3TKKaOixfr7Aj/SZOBGpeF8bXvTDXEUfUc/Z6F/5bjz6RifX4lb
qAWc0zIsGcLpLGhVt9Q8dFHZ9Zf8Lrs6tsird/WNBrGkc8PQjAJPPjwE0IDm
ySx5u/2U8sIIVC7EY7F4xnNlHURFfTwTd5s652AKeW+8d5fV6nrwiosvKg6s
MryGiQaN9ijppXO/pJhhJ8MoCXbSu+spllYrMJ+WwnESUabjOvthZmjIwD9z
fz4vhjCZu2DxCvqyYA2LOIibn99+zAAtU+23xSdcJUip3eLvABko99f4Rwez
T7PgybdVpyn/8WTSwd7atT24hkN8TX2ogC4KB63X3fGL9xxVxPdb04P3csFH
yqY7H476/ldUL5OHXyv51UK0piVZ1caztmamlvek6dFL4BHkdqSL3VOfYIZ7
+OqIUiPsRTSuZ069ANKKaxfdCXa+rJ2lI6SwlJehQwhH3T2X9BycZDSeLrO6
4nd8qy8cwklGlUHq4iBeky02K4W6he8u6vwTANS79KXO/5MSBptbfGHebS8w
Bl3w0Id7W2XCsnRRmLTBgcNeEgX7ePzqyxDmT1fO6uLsXuU1cmjTiKEVuZi1
PqEWKTFM7KC4IUU+nzQx3zjkH3dPclnr/CQfpizH6W8NnEG35dyCY5y/uwJ/
sitEIupCkZBnTkZ/YcLj5x87MBcVLprrMWfjFqWS6wrLOm+VmriBBo77/+bE
dNzPLqnJzgrAgfznfypaiPc180IxesGWcGuQlOgmjH8X0BuLwYiwntyjtACH
EUrvbEpGFCJujdw0aEyxUjyZAeRY8vQ7/NiuoSl3kHGBOd58LzDRUdsiHx9H
YJ0uDKQtR5a5lnvHfqAIMyMOfFhrFgUJm9GEjnuHAG3JyyN4rweFBL5icFtX
Y9EcYnUOr/hh5Rp0h3CkzbCx1jWGyLZxFrx113RWEFbU2ftVxhrJxWF4lOpy
ja2XLDRHtuUe0MYi3qG3TTZwemc8GrSMVMw1+DaSR9OsdvT+RQdQ7ry5/O1B
STTpHAVcva9O866OZl3q92lpEzLCG3rX67SUuAynUAG5n/5my7wqQ0i3avZm
/x/jlMwXsklw5EzHOhoC1JlKbKejoPYUnOlk58JTktOLGQi38cuBybv/VwrK
BOgyTm+SU6QTPf9mO+VIWW1hudraa2J+Qnh6LvGWOCK0nMpvc0DNxkvAun2y
Hq9U+mg5YhkQIdIM4V8hXRv7ucAR7xFg8AAro3qFpxdg5ku7P5nRW83TuR5O
j/3iOdZ+Wknvmlv16djlxiomoN4M/5AhTET/KImr81wbEAUjbpy5R3l4gYCN
oC/GGz2ZV+kUr4NXgS47D/WaFHm83fYt98exxrMOSUTtd+EtZrBuS+EHn7kh
wNlIzM/JCVxfVS6MUnsQNXWtK7bSs9dbAf0ESP7S5bx//yBh/CAe0lzwvhv+
aSvE4DaJfzy6F+5h/W+B18/HYSwIfyYCFUl/bAtzhxQY4NE3Hf9wi30nS7lo
QqHNNJCWtjhHMznYZcT0x/5vacHmmht7DH3kC1WN/Bi5WBA/HCFif/ZqCPrT
S0RdtIj9oGPV2uuawo4ENkGSMvS2aZxvtpV7RlhDLFCnUXzyvp3FIB9+oj+V
OU3EMhM4f3Vfkv6pfmneTFEOC0SzqhfP8KWVXpATYbPDltYrJX2/VfTD9UXw
C+gaqEdmPZ4gmoF7zk+Jwm9/uIKN8UZilWwG6jyHBJ6BP3fMA381IUFuPIel
d8xpV7TLm82y7i8tR7cxYB3p+IRzUexXWE9CdLZkjYBBON2MsneXobheqzyo
Hqud0lj4RxrnI5lsRszAdWYAwiMH3sp4lhQkk5V7WDxz8LCoFbnRwGcFnomF
SKM8+2NEn/aEGvk6/qHQba3KQltn9x1rRrG/ff/hTU4cRCReksCOIXR1fyoS
BqZ1Sy1R69jGHSgBJXo3JHknkuAB26A900LljRcI9LqvURWyiem9VVA38eYq
iU6l+DxlJ4Sk0SBXmQuwzTH/o636PInpNnjwVZJOCozObDsfDRxw4eleTi8H
qFrSMPw/exl7uqYzetJ3tI45gSxgQK8VDMPxm05BYJYA5Stsav9Up+0PYCJB
JbnKdyRXjRvlsrD3cZ5AolufkrbePnHn98AHsWe1+9t1Q9RHuF+Vd9hM2GeS
dyggFbxVViDzLfnefMcJmW7qdYhr9MSz5LVIjLcuU23BdolXSSmpVyxooyxg
6wR6O4bNr4dsBQfn0vOqoRr+5YSZCudpgmqFzxnmXbaKFAQ/MSMtSHYaQX0X
sEUTphkbz0JoMTXE1QOQkYQz6Aaa4KnrOvviLkIvBkStsHBV2vwhkshbnGbV
ktEbb9Y67aPHqQlJaOF0zN1LVY3pZgytDHxq1OlwiI0dEPKA39OdDFlmxvv+
3vkOwDoT85YG6I0o2LWgcye/e11KIM351Asufizln1aZGom3gcguY8rVk0mf
JXN3htriEhhREyqTmKND8MO4PpmgWommnOZAF6XBCvnk/AFw0dyj+cjVKUwI
uExlB380ORk+a8jZiOnxYxphak3O6yAurtm+bu3oVBzN5DjOAnhozgau7LgZ
rLT0aptzHSKsizCP+rR6f9vF+0Kj1H/itqQ6kZrJ8QkvWBgGaIwPBBKSrCSS
Q+Ka9tSBeYKEeEIhiIbKjQ7UF13mfp+1eOwXLug5cf4zKmokZwVrRHK16lkt
iGKrBBqzn/wLoOxMUCd/nWeq5unS2y8ltFXSWbENCMVIZT4DCMVrEWobFgcU
lyyJ1cjO8mm3oklZz+m0JLONKQ19zjeo/VBom/noYhQCvwqLrpyj6BTSYGDS
9c1DjHSHAEP4EIPiYPsT1kpScZ17uGt0XFHaYO/yW9w/FrvD6+eDfd0nnGQn
cB3sKQnP7gdjuoue+kW9XoNwqXy7Bdq6azO1ogLe0749Ca/1V/3dQIIzq1Tx
8dUyZIys4R6+x4iAyezPGO0guizl8EbhVfK8h2cDQSFfKcOB71A0pcUFqM31
kShsL99cPXdWcuI+KiYIsv+OMIxQecpC0oovJCfzk10gEfNz9hf2TBfFAVjt
IGJyqPAjpJ5EuW6SlSWDkv4JHlJh3Y/DCPeORkVudLkl/5ia/ji5kOnciNiZ
4okFpA0oZCPMu5GW0uHeCLfvlFIpiKmVG5qdqEVk7p66GgkcpZ29UUvqv9ef
+yVYoxjeG4MNnZ02LOw0h1CWJqSzKc1mWN62AOYju774MwfI6RuFvHR1sPRm
iS/tqoxR8pRKXdbsYakwppqEXLkFDP6/r8wXlqIT9LZKxMIyJTJWi+p99Io7
Y56VVXDtqL58glOPvqefPA7Ba5D20lELl2UGO7RA48LB2UCUhh7LA+WeEA5u
iFs48XF8TkuoFT0hnA63kS7x26PLwFFN9FR35kKzCSRYbnZO99nNlOc73xja
5gQi3+VHTdmat4l2CkUR0g/NegNlnt78Ofglu4a+Jr9InGHH3oOz4Jn76588
qh5qSLSeIVI3xe9r3epsE97n0UY93NhqGWFeUqfB0FuIXf7R0QYcGHz1GC13
DlZP+0i6iYe+kfGhbkFzrXYqYz9PzQvjqbJufQpTNllLXaghFR3FcfpCgFsa
CMzowLVPBIY8m4/MKtqUCAFongsVrVktgdMs8pxobEtgYMYGLN7m6h0NPwtQ
hkIHr8QWRRXpSYIwYlB7p8HZWuaEU8uFnw8XDzUIxVpwuUrmdeTkb2cSiNyt
AeTlBHzLkfqB180XnE8YTLTmI/iiDODfHjeGj/ubfsQSKwFItZTMCjqs8hpS
agbCf5hp0eTB5JvxVkdGllniYlhoVXDjDBTsHVHNyHwIcQX52L9VpFkWQfOS
hIfHc8EET0ilIJHgOqbSALSELCG2+xMCJ3lmgFepFvqt08EtDolU31bPmErx
60siy46JVr9xzGed6P9DiPGCD17xwg4wmhOfGUOhuMFvd/ZSEQq0M9BMvicc
7EjYd5qAED5TrDrlPBDOsCAnLOAvda9dlvqKf4M2jK4+J4bAGCgo1Qe2WuvR
d5C8FkBiJ9VW/y4rINsJVRf3V8UGSzi2v5DSbry42jnLUALT/LcOTLk55B/w
0agNcWmgndW36eJCnCuxmoy994Hhlz70PrXAV5VF5YcgzfyuZLXkAt6DdE5p
OIEXo3fq5P30gyMGlysC1VYRcc0gULSF4CgFDNwLZ9PXAyOyvSvrIakc679s
7EBYR6kCpAPM5lc0F0cBf0I7W95tIA3R+bukl/6Y3JdBgN8NOxIERLTxY8pU
i3YHbnWBvFn9p4Y+J6lOWhxR2llwFh3it7x8JigOBX+XNCDT23to654xdrBy
QdMlTmVRIligBk+fpU+A58gQYjkVifHVvEyY6dwZjGePnrchYzfhOEEyZi98
NlV0yFq0KIxv+ONZnDtp6xQagE9B21FPJhMe1Ic5dkLlKBt/s+KzHcteg+D1
feMoL5vXV/JyJicHOK7qpSctw/cw1Pi36eq6vJ3lByDmGxHc9egbCMgI46u1
CD3eDXG8Cd0fbzVJx3h/fwMZr8Km0J2MZfomY9kDVUb0B4ajCaDaY/XKyZ14
VWKI9YPs/RMYsxIu+cAb/AgvLoXAdGTZ9MBJ70aLNzSZ9M+AjPcl46OeBhJh
bOOt7pFpv8ukTWcIBoNZVFcAxNJ7YzvHYluy01Cuz8ExE3EGyN1IC3s6ZCrx
5tlRNg2eR7Fo7tA4nthiPffxVXZwnhcV0FTg4pruWcVTW146jgzmzR8OR6N+
9N4aZZgL+tOTtB51QLhLUEevjtJM2JuWkheIbKirFO192Krs7RYG+I1rZY/R
7rskwiKUpiei4Zfm1CGkjrLpqg+N1BxWB86R60o7hIA+8mZhN6MiMo8CSC0e
4+b/ZpbmFh30EcngsfkPQKYhPH3ZawAQe2u+QYkSvUFBS1QLFJ8+G5L1rjxk
uyl6hZ3MxWbyLkJqFs+s21+TLH2hhgJv8nxtWvBgLaxi1oAo4mNtvPDkeN5p
YdMmAsb9Nidu+A99TJAI96mcRou1nCx6hJZsj8PcWkpkte8ZvweTbrrgjgaT
RVuE0jOU1cAhdsXR2SYiZI05oS4SrplDvUrH2KlzhTZjoOTNJT23IWiiUb15
KX84Y0mmPzpFMTPAG/x4+9py5cNybnv/U9pgGg/bVWtLgMVgOyRO+I5N46+I
nNloLXv88cWmdi6At55ihw2qfNaEVLaz7cM2PDSgEz1Yi3eFFczSBMhlaq6+
LlSsy2Udgl8QnddpysSTRNEn5r03Z41tZVZ8aNsUykpYa+JWvuYMS/GOtvZ+
8EqJzL0v2OFE5Q0LC39AIiBVJyr+5tn298TAdK/ZpqKEL7U0ENg/2m6YLeyj
zxTpXS1hvgRq5qarh77SYdNHax/maqRhjJn2WgQ0y0v0IMO+Vjdh06n/h9JB
Kcq/Bvgf/LgGIDnixewAuaUUuqR5McBkD77h1dEgmo4Sdhjg3s/xpUgyJBgg
ChGScA5ggTdgc2WBitWZQXEppERs2X7twmcSotKl/vWuMP3i8ociz78WqE7y
LT30k6hjlqsIB5UTeP8fw7ovay8u+cM5i7FhOrbcqXg5BinrfdPtwKclBVph
ZpkT6qHOzaCbEiyRcW1GvXIPOVLGgIv4kymf3MEJFrIR1BojUvRWbA1f3pXZ
qc8jPm/Yj+7ysRMmlAVqLJ4zC63zVClolTV9qtwM2d0qKrok5Phq/8yG2lJu
DbrlpUdR7x8MxYyV/2TUnjXBMCLJICj/ehp/eb5h3NoesmrJpEiIcSXbw5bo
9ND1M6by5RoowiGAJrzfuUfLcLPUsiUKTXAjdQ/i6s76L+Nyn0kkS98O1EJA
jyI6w/McAOX82XUQDjRproFUfVlcvFuenVQfrKAoxEzndeYw6iSbYV43tMea
uvA7knSHnp2ij03B8fgryQtPh9gPrzALGnU9pCD3hbbkgStvxsdWxI4HiCT/
dUhgc9L2et5OJPKoLE/aCp553U5D+lkYRRHqZNKAK2wYjqos/nUESHy4v7rR
K+8/cqTuPGWVD/u7JJeus+xftI74tazE2M9rnUKGE2EQrIyVLbroIOnX1qwM
dqG7Zlo9P8cs2NI2H8Apmqq8XpnFw5+Ogv2kjiug+JtNB3LZy7G0pRidV5Cq
uZqpbElhlZM6rORd+U5RgMrIuhgtiLPeSAWtv5lZ1newP7U41iN2lTBsOayZ
lZhzKY+Ff6qbLjcBXuk2UVATgGSBbP+FZQxWHU+vMHodsAa4XOa2uemhACbI
92OlWFnL74RhPSIZkdhog5W+WengCLbhLwAh1ht/ix4TzLWiLtojJUhmcutQ
i8U7c3irdgJqTF/Xfl42VLtpfPgluWKpAU7cqLVLjPyK6E9+1Tw2lwT54YOw
8Z1xeW/FZQ7A4qMYeEAIHgtcBTwmS2AxdL+4BFLxhx3BrWTOOzaAY8inF7pZ
5Ci3tGeDS4TqaVHngsLpEQ2Al/XJM6dchr7M5NnFT2uaMmiYyvECLoDR/dt1
QXxD/TDZiLjwl6bJud7W7sGQjJ8NYJ7vDrP+CN7ZKYrfHbUw5mTKeT7EMasK
HTmKbetPRsC1FBXpOe+NjAA7bWYdVz2pKI7qcQmRmSY0d9AYj2+2BgUH1MGK
H3w96GLefQNxcRnI6ZLFjm+LfBDhX5IlG0pXfTSDtyL0rYS6xKv1UDuTVuOy
9IYYmsLHpYce8I/EV2AMnEPV4qOHQVAr8JQfe1ZA4Rr4TIcaNm2OEForgEiD
HlW1Ssz1/qMmEIPGNSl3C1fWGuimBnkwh5vZgTbPuRRo2PhacYAULZUs3GP4
hdDyArYCLfq3I6pJ31wrBzCQyMZFtzYrXjtLVRvlTjtpBFeMTKpWte3i+you
XaqBySKwR/SLjaaF5bn0vWJyHD6bklFS7sHUBGLnJRSXvE74KKTLi2BoLrux
AEIar4gfqo/tGNJX0qIIyi23ZekKSyAyAbR7wsUTIkTR2ZS4wdlTzA86j+Ri
vfVI8e3NoPnE3/67APWkU2tKq9jYW6u95fkRqbTnMG0lO4wIEC/K6gEkvrse
dMB55RlYXxSMx+dx9QPRH51WZkXyeyWxvYvTV78HFT7YkKleAhIhUEPt1kB3
5R5M6H+fjDRDNqHmplMq+acWoZYc8c+hw3h+OXr4xdw2NDqjgGaRqGRA87KG
cvfZSw+k6zo7CL6rAY3ZxblUwkmFJk+5DUaYbH6qohw04s529pJWb1yoBSc8
H9JUkION18V0hLcoBfsASFuQWMByGZEMU9ac2wFK8HbOuJ/d0sLKiYTerny1
AT+KA8z1Iuqiw1F5gZ6wNXkcbHw+75wV1y/N9D4L/dMz3T2BkbYBeCJIWxPk
537SRlUCdREe82Lpv466z4xa8dQwDOJq87r6TLa64ePi8N5EVHaX1CNmj+oY
3vrpVdjQQJM/1bpQdgqK+lWJPl6G5sM28Gnzb0Uzt4MgdPqkGpa22fhcvS/m
oTaktOue/le9p0yh8XD1AlXKdg0+ZCiZNPyrOcCM1RgYHT94A5iCLuT5cJR5
0MC2J/L58Vcy/M6qKmki/RyOuO8kYu8Cdff5jzLHpbSPTR+lwNPQpKFHRtf8
+r7G0fawDjWjYHGxYehsIjTzDlYJ1vP5JiXVrW9gNoSy0E2Mcm8qh8Paxpkd
NxrmKo2l3ktQpXaI1cNoig8mhnTkO9VV9OWcxmkETbeK9WNUthYqvEG16u3Y
ol8diJGhHK/kH2low9ygc6oeib9M+dxjRDyo2ftAu3ldq9WOsbgcPxucdwXQ
QFilDmEh8LAq9rTY1SbdrfMiR/xuUYaAwRr8ZMItkjRQDOcezDty7BbWXWnR
4xDCzceoHAUMocETIc90oTTOm5iFBcgsa36kEzQlxtXPfDMUpBaw+IgIJHJD
PBfjYGT+yg9Ha6Ky48Fm1K14+UMlSwBviKbRLzUCTghrmWZnICP9WVk5rxRD
t6Wiqqfvp40Ut5ChtiYL8qymLNRp9/ubFlhZ43gZBSxDrIjM50hIAdN98Uwd
PcuzFtNF+VfcilBCHF7tE5YvkHFmUT0KLv0BOGoh+VaazXuSGCwaVP4B/yQ7
mYnzaCHK+BmM6huk9RuIG3FU/feZEHCCUl54xhUjVITFp1sBKiIiFEQtHEnm
+MVJfmdeONc2HDpHXlduILFaB/jOY4dA0M1CWUoZXVBpn1sgdx4Wc6KLcLB9
tlr0wcRAoISbU/t9QntLWdjHajlcE66LexytZwtjyFZJIodw+j74p4GEsfoj
vCXgf2MkuuUpcSZCu7mN5mo2DkaLOi4CW3DnlDwVsFZxBzKbOKBpRJTx3s4t
+KkjyuttxxKsNmoI1bm3uOBLEvqtpx6agK6cdlfs7YLEcxOFn6p5G+vgPikf
6EbB913txOrvjNlrmfV0JW+v7gM99psThPBfd5HVBeoCq86mmr16jmi/qW4n
y7uCsTBhZOwt4d5vEsbro0XVF3oiZAs2XAwYgQmb3JnEbILBhBpUh2wytp6g
ihjcX3HtgifvDseBhqTYdo86uw2Mr7tTI1/lDe3cm9JmSYTEMenP/fzJ99Wk
/FjJpRfREHQ1wZvHL7RwWaYtxfE0m9xqaxkzGp/Ws1B+RzwMfFawpGWm+uip
ffjQ0cdFk4/s8MkVHcC949a09Kzkr9MEeZxoLmyodN6REFiBYe2M4SWxgIz1
2fhQOXnXnkfNjLxMnMxhChsivMpm65FXGASSkwJnS6/NOxUuKymRocEovRHR
Tt6MYR1jW05x5f07lO+gx3zsVYNwDJQ35i0sAC5pg6rThBRCOq4vNNLjMWGG
1PUoq1dT2MDX1WE6OGBnKXsjMeEbJgsL20sWazRGJeNdnFzjuywVzEZeF6Fj
pE0BoWbNAr5ItPM1isXMOSQ3s5Vw0Xf+cuzzyNOAUcHmQ7wko7BfjB4HgUtq
lsM2tt84QV8CtWO1AScx2nlYDLJM9fy5ajUZshLW8WCdZzLlIa0tIS3U+aNz
QMUOfrjp8gy9WmN6wiuoRfFpKzEAN3AbEAtZ6/aYGELphq4ihdbNtG+b+ya3
KrhgJ9/swq6Hn76Fk42sgpwsIdAWI7LTL2BHHRYTGkNMOxcOUo288Ax3otzZ
FoaziBLWoUezpD3MQATuob+HxglExjQQkgfcmrjpX0J4IogF5z9BIzKeycYh
bD9X+AR73qsDOzzeW1klCTkgsJj9x1CHSUJ8Qxcpn/X4JeOqbfkpXL7ELQj0
qxmjjkkpjHHM8kAgLcJXaSYQHcPp2td/xYYcZnhNdgFFZeNxRh38n5Qec8Gz
iQi7UDWsI7A4nSRJ7Q/y+g5OHK3mSZ8XNrYBCTsoUBWIMgtn+KdU191aos7Q
aNGAAtexOPOHmLaDTeGT8VWTbP3ECl/qiVMjRMPQlnmqvPu3LWj2RJB6JS2/
TU+H4wSmG1S/kGhhNMmXZuR7ehW+za/O61PEHYz7a0FOwqffPvvy0FH6dzmi
Gs/vgJavVxgTU7nK3MrJvAzjG6BUKdhH0fnpSyzVqKi0cbVtrFtZen3T8V9Y
sMUTf4q1ddZN+GMURn1qwdaP1BALeWCqrhOjYpZDUAqXFT8wtGjpoOKHenne
b6NU9Rn8+vfmqXxggpB/GXiQ80fSYBVpTfP378Ycya0D+LGKCHXH8L5rkATT
p/M3M+O6ygcV4ibAlla+/0MJHS7W60baJeijWnGbOtRld0lVlaLJZEf+I3LR
PR1UQkskm4PNh8nSFSEt1YAkATFTfecB54QfqIyvWnJchYcnYGiJBtg7g7pG
fanRfBsrBphecCuRSptmLi/WeBxRoe1OXMsrkGjGTyAxMQWX+eINP59dtWCf
4qndTC6LUURj385tVxGJM4zdBhPwPQN37cinmv1cTzUuyDjO+zx2lip2sUo7
zubBwW1Hy/HxhVMoDba+AWV934WmL8i6uxcjWy6tMPHqemIL3np8XjHWoByE
1/IbouE7aL5SdZwMQup9/WORn6RYevu8zv33q+T0Kn8wrf+S4mMl2tftquyp
MBdSSHn4XQ3jpeTMd++mkoMErEudo07poJHf58QsEeYaVguocQreFxc4gwJW
xQLODJTdgjEcXI6UKtMIsc6x2NuhJ5B8s4eDU5BX9NlRdNhn+DzqxhdcEUq8
vDuUkB9enS+XaeCcLf26/mpEoam5Hh/ujWMnRugo57E0yVN+TIBXTcxiK0BS
fW71QBE9g0L5TAAKqckJdLui6F6iwMML+LOFhBRP8p1MDwuVzIKVFYJbKD9B
xESRqD68/pjwnvC/tyOWh1ztW+VWYvI2jFeaGW1nv7QX2hmQuHC0wNpCys3e
s4nVEf5c+ke5RJN+yqQscFNMSPz6cxrVgnBB5c/MHfm0WGbLM5V0aLG33B6N
0bDI3kD/Rzs7k8svVi+DA01IFJu/xQc5gh7iI2FoUtEcKs6SrsKvjTjn4hxP
qJx3D81v7xUPI4d4TVkgwCceFoekRAmyQybNOCEc2w6fG47joBLHvtjUr1KZ
FcIbBfkIkdesX/OVp/vTZdYULvh8CEfgTlYaRwddzN8gOHDA+HDSzsP/U7l+
LzXx1Crqdx7B9qYXO0dCckTj0fPYK4Q72jhHd0UWbljY+HLj0L5vL3bW9ELR
l7ZGmH6vG/5wbfGfoE7ibeuC5Z47qapx8AlRGq7FG8oBq+1KKJBEvwcIzl29
9LLoD40MkTNbnsNds+bHIZmscwH+ODI40zwSSW21NAS3nc/PImEu3Y2im+j8
Z872QK/jiIbfwpINeam3v9xeVX9NoZ98EGPZLs6JfXoBUvsqegLTai2GjAlk
1QDRrYK/ZDnKeGg89YU3fjC2S5j9CFG8gyP+jWXLERlQw4onYH6kdW5Q1ySR
eKZR4iDZZmVhA/TMJBVfMbF6djcAdHl491KOH/WJDIf5O0d1wQogiA+RvaL6
Tef8Sl8pXt0nnLzi1L286KuH5xWUtwSx0OVqK6UGFBUoGc8sUhEiBL2SfZof
mc6LOr3DeCt31QAaWc9OEnIxOHOIQQ5zpG8Oo+evlgzKf20Zo1Z7lvxbdytL
yU/HZ4ipEfUwrSs6TSwouCjR56cf49WZbS7z5IM/SrKFqtY9I4pGgVXR1cc+
8X8W22MVeYsPYcP+sviVNzlEkLoaQPVsPyeIoFqPzFg7EfbXLN48QKK5taXX
S8DaX9NPRq193baiMz5gypPtvI1rvFKYXQaNyXuCxhMTC3iX9xJxmW7JJSVB
g8CFZlVGs1RCDSz9BwlKDd3da0KvuXW0TOhDDwcct0+hKLo+XpPd21uGIYFZ
yIRQGuZBGdbOcrkVoOTTcG4HIqx3+X2wq2j6Pa0acrGj7pFhsyZTJ7Zh54Np
IAk1xMUjXBNHHwSLb2WkootvWxgC/twiNtcOFiXOiCEQx1PTTeQNNTlgbpiW
+Ogry9/mkEw/PdI22OyFG5FUWio7XC1GSAaJfMOKIrbzsTCCbQHWhHDjHfnP
7CDf4oYqZDfM6ZhSeuvs/im4Bg1bhPRi9mBYdtwBhkifdUE38DYiiekARGKP
rqmIXmDSm4N5Bmru+MQaNy/rwTTJrA+6jNDH2oiumgREIhUuYjPxBc5T9oVE
HQoZu8IrAAIJJgzeG7ZTin8fj6urQcIL7geFfJjThedEsqezcVXK6pxmW3ej
DC9s2oY+UhDKDK81KODy7afS/BIakk+hbAvrr49qYdCrMtdcvwnsXTnmGpIG
4RoixsPnm/HzgTiuu7LVlcw64PGZRRW9rN3jbUug2tja+wdUx5QOv4Avpiwd
xkeOoy1qEfhClw8DJf6VGuv7Gcu3yqNirll74gxGzQPFrYI6EN5GzhBhDEUG
Fz3SOUiPK0N6ygiLg4qiqiSrs2ONCMoSyI2Nd6cuD6WvyVF2jczZShm+YBce
GHA2Kg0+hFGZU2ur9X0RlTVSjIlJoQBS/F3CQjpdtPcNvJQtJFfzUnNoaRrE
xdoYdYXZDid75hhS6oeTXujiv41425m4r0PIjTVNDblXo++EouHkfZRIH/GS
DbVhwzPGalLrQk4YoqxBjf081TeDV3OZb9YtijXPbyJebdut3YnA2YhSo8/P
I5KizS+cZ//E3hVIQFF9p+MGhumNTDhmHt9kEnDIteMqi0LLYr9b0vY6qicf
adW+l/LDrE9hBfrr9TPpm3XKS3NWy1MSSp/lETIgH5X8k8nQyWsIAicrV2Xn
6c/xuzdiCaGVOn4qZwhCzB4ebiDa06gpbVnllSNM2irxES7HnXeMRFEo8Do2
XIufWvOXEx4l0TsrVwJG4q2GhUyJuWs8OPqghKjDUY2tqeJTeMpZ0yphAaSv
cD5WXQ7XLvTV2fjOCLhFmwn1QH9NOgLOC5rmuYK8jxCseXcwhn28NBvrZ1Nb
krQZNKiEYmFqOkw3i3qstRtg38SbMJMbQmhDWpzy3NdMyZLN3v9mXLQjXN/c
IxSJoiSruNhFQnwLtPUbwAo8WCRgFkdy3F0sVU+2Ob5HqE2EauDliIJkDaLW
ebD20vJB+WDejxjUdpRs6Fh04Vgpz7v+4CYbUCxtZk3Nx49YG3BRH/z0PCS9
tbCTXjEyiOx70Vnr8T4kO3/+HA/jD6DdJg6S4CnoJwNcfvHJpNDVb1vYoLB3
Gn7SKEouj3oBPcHnkFXUaYRfRKU4Q/L9omT+ZD/sYbM0OILHP9R7A92g2Ysw
Qh5ul1eafitmMqNr4hwyn2L6m0RctT/+jdSgXWMeQ0tipCapSV6U2IIDXdH8
0LoUHymz/Hh1ZBBDafAP/Lixla6Zj0wj2xUFnWXaFrFTxePJV5YJ72xYQinx
q5vw4UI1dHgVuqYsIVB/IsX7GtFty1oITiBB6vQSjV+8Gg/KzrGCzfUhgKip
i9IUDvD/nxd2RIDyjbmJPcqmQ7HHg0HnKqOk9wg4DyAfU2iLE90SoIWtxjGT
qSZ/lUwC7m6YAgNozIqKCzMcQxd2ogLGzH46WbkeZtTb58hWlrLL8bl9R8Lq
4xKkzLmnoqciMgSIFaFyc8hIPDsiemOqHSB/2+ONlCDJAI83QBK4r17M9dvX
0qtq3QeuqFtzzlxKoHDpBaZi82cZ4M023Y9x2IBotC+mRbsTF482pBcjvIVd
LKUtYga6dR6hB7xDAKYH9cinf34WoI4c0tqHaotDlkCRBVZqhHXUojiE4hQI
8SMdgnIaS1ddI5xZCHcF3MOPiIGDarWFky8nA7FNvzlwd9n8uQjXuC7ce8CW
w+QLxvf+Ufig1/6/DwASBRolbcUulcDhqCj1bZK7jq57I03cfYPL+xjPwQrK
8h2D+1LUrI6IY8AitT95bb/bti24oe3h4xM6vL5hizWOTfveVdkIAe3zR82e
nxUtiNrkWRrj6vKC6Xqi59N2vHPHZxfNgSNm65oaR7TNjrJUYnDznU3xG1NP
DWMxzWGvvbINyNBl2AfIqzJkDv5+YXKZczwGSYFb1zUUZ4Ijzoz0L+Uqnjl2
UNWtTl0UbfRCSc7YN/EhnCoSx6exHT0Zok3MlWbf7e8LSCt0UmWjqeaAxmsv
h+zxGVe1R+Gfdnm9TasGZkJuLPcmQTAeOiNhMFsd5zxtnoi9QoUcOiJ7Hygj
IBwZyGFTokFYv16t0PbAkLCBtFxyF9lNVqamXHLtFKp22OmVgAuy30MThH4t
h6IMs+wUYOtjEDCUsv58zw84q10JDoW7rf/2p6Sz09vkWIDBUIodPWOWdH7t
q0JKervfUFTqPXsL9Y9IHMjtj373k5J67UGs1/VmmFu8cBWKTQ0PjhXz3n5f
qdFqbVgtdhh3FMGdsvMjClNICR5V8rHcONv2tDELtBphsUxw6BGpXWcMTHMC
iK3p7YAmn+YSS8MHdEWo16JD9EoNPNdfd1KEbaZVP13/iF9hU7nWAEJs/WOl
DxO6pIiW52wpakdRZs5fq7eXRe0zdOPUbw5whmHEkIVfxjR12R8crmdy2INr
NG5gbqr7ICGzZ3EhKz2akMiUlvzQ1VKvTUCwWndXHocMnnxXEcdz1U6kkBXR
hLP/AhAU11AvfpqtdxZQTPG5LCXMci22ODDGcudTPikB3SW0wNq8fiJbH7E3
Lm5j+t3XY6WuaKykI0Sj7yMpiLxK6IjhxgLDpgR3bOKjrtE2d2mE5+hV29fB
0T1pDoj8K1uNtBG8FKi/4ZnVEDQ6d+xnjcoCZyYCkL/AW9WKlmsZ7IWyA4/m
M6eesgmEYAOTW4dK7woODqVY0XFU9WrCp1dhkp+Bz0bPp+YN2mJ1mNpn+0s/
OxE6uZMF5PmEpraty6q00nL6+ntq78ZMuNIS/vH3/XwlYZYthmbsLHiQ5K31
C0tT1IX1BT4GLVW9dgoD80mHLRwVGI2rYAE/qwpMTD3wLt8jCx4tcYiiy9K6
1B3GoPQJr66TN6dtuwgGXDrOYe6+hAl8TVUr9nNApxbEAmSE81fIOh7X9Y3v
O/UI3NeOXJ+jipvEnqDD5gk3LjxP86bXGLePRREZoENth4wkAcRxXejsUOaM
xUjd4iB0MJhJLgeXLEhz8wo+BwzUrr0jelbhL5WAIAtYtvp8UxGb0OehqO04
nlpdn8d6poQeWGeL+Rpa77EPLdXXGYrSflz3YXvGgW950QM9Z5gPC+l5vQPH
ENJ8WNLQRk6q/C6kpn0S5KGdTX22s/ZijdmEdLiUgGCv0xth9m/4EiQhBYJ+
wcpJZLsxSge0GQ+KuZvSjyFkS+eHyd5Se8Ec9OK54MkVuy+dkhXsQYrZqJwM
VAyiz/ZKwLcn62RkHiTOVpP7YMfsgi+EJEkiMNfhDrrofNlJerk1+Mu/JIW3
DT8vqAfTto7h1nVrr+2T6ZR6UAQQtXRrnQxUfBIaTeVog4EAi9tCu61u5Lub
HRyyMAGFkbODK+mNZ+yq9uYje5qmdWA9iu5Z7NBhUx7i96poficgvZqs3p7n
RS/4+51rVkV2exDHcUbthliz8FE3cJKUMPNZC7G2INoz+8flZigjH8D8o6SQ
edzXxpcvj5OLZduwa4noI+gIue3bTQFzpbEhgaHd+XJHmd20QDnO+Hz/oKj3
BZeE2FHM9DEdjOolMKuHiDQVPUNU/XTetiq2WHTmEOTMB3t53Sa20DKS50Wu
rGiaM69r2BMpi6Wq2WqcQDemuA4DsF8X5WvGZSd+ZuKlCDtSEEWwLVURl+cX
FK8qaoavS/39NlE1F1mGZVvYLro8o+/WOgtHrJzduCs4nq77Gm3LJHuokWIp
VoFK86YqDVacvqHXUf4rL6tuuvDLuvYnPd1dlbeerl7KFLEWev0E+7mz2KqV
vibTfd4ED2QlQqrGNt1n8QcTx6ECVR/Qodi01/eF1nEstRNITlxvNFnX0nea
Nikqj6qYVr/19qHJwkB0KqmaoL9hvcLZe9PLy//WYDOaiiIXZzfc7MEElBrZ
X2tTRe3YVV1iswuM0DcTefF0tOUMzyRDA+G8GYiz11JVsBw5yy3aGsPtaXYI
D2Y2OiFFKM8uYi8UtzaT1u6cp0ZRy7rUCIfOMxCA0XLezg8P+XUD5CHMVeZF
7OADiWeKOlRqybTjPRFoBbUvoZXsLeLHvYZh0PRCtJeLCMPNd8BsXKFBdN4C
HAaOkzlMpVhfb8TWjF3F/gHUzllhamm9BGSov025KqnBw6aia/pdLeoYlEde
UhKlHFY9GddA8Ei1Sn5WmqP5p+epVemTfbDlkq9l/LEs9f7I30ZtCgrJR2A4
pa8LCEJKzzYi28K4N+k8ZvEb2WI1hLX0UjHNSZZE5Ob1XrSbMjCjm9IkYIcF
hr9OM95nHFZ/xE5MuMPPM7VxueZfIXcQ7vexiXisTqqtosjq5uWisqNjjHZ0
yTzeDIx3Fhjm+wNVR7GqmvnMD/Q9ZK6nSnaag4xb5VjFGkkhUCpiph8HM5bo
5eCVVRKb12fkKKrOF/wjBGwWompubJYQGIiRTH3XBU24ukXy8xY7zXXwMzTL
wXnVlZivuEMEaAGPSpsHrNeYMhXNSoW2yFeQd23GmDUzTTiCDZUEMzxSWAgh
/vPvRuLbmJbeghxS8yhmeMnig98lIbjVPCvrbKG4TXh5usRwm6ER7OG6nMjS
vkARZWdGGSkOyvFPqcOj5NALdgr/zAbG+LulMxHp16aAWZQoHsdY8bYwwQil
pZ125bUqTCCygadGlqVd1uliQH5XG4A8T7X/0Huh1P7zH8sM7xXjxADoKU3C
TnHtw1fDtVV43Ztat+tDjsSqmZolQYCBAsTkkKHvEKbZRdoCI8Uxz6c/PMVL
ef/KtKbEJLBoTpVL/mQqT1cNf8VPQuksi54MMlnCewvXQEMt6fzOV/K2Cv33
Pu/OSi5l+cqwHL++lVQl+4igZLgThnZkcPL6Ww/xYpWdsDNDZNexLq7siq+u
K4Msu+LLQpb23G1+VJq0ULMbL/YiJsU87aLR1oK6rZuhS1pFDDTjdBSt4Cle
XaC7BcLdKLLDaG3e0hgnFwYYWuRfb78tJQaORF5hoCZFj3O0c66qOInpZgb2
T95v9mjULDqw6e0oUcKHTGbPYyqjjCc6t95+PLZCBx3H53jnfz05ZmPLkPgV
pJLkhmebg45kKjnYhPrJicLNG8lO0Sh5u8zdppOKQ1tKjk6woBciZfDxCEGj
/qCmz1G4KB948/4CEE6lYT5t04mBj4C1GMhMp3FOUEclGtz7kvH0VqN602IL
cbn+bDfcqC8+ggPMzFrRqLc+24uvV29+ljpsJz34K1SLEO1Cdoh9ohHdV71Y
vmXLgbwCh3Ldi2Fqm2H2pV+HCCB55e1QVNRIcToynmlNEWGrZCBBvOq97YZe
cjh79k9jT4EFwBbM6lFYQL0aEB3xOgvALZa7idogm4/3ExRXY59PoJ2vZG4D
+7XLypzREXVsOM5OUNf2AWAmAqt27qgkCC7thgBLo+SoJAXVq9zNHmAkBf2p
y8QLGAB/EwpTbvMEo8rbBBfZCKFMMmm/m3fSmBZF7/bkRRQgKd6zoovZyo40
2n0RBwXJAToxtcUolBlLzqew41rUQUN1X63VrTopHG4MJTR0dwtZx57yEqwu
derJECt+++qD+vzZgIO2uCbhIvQxR21Ii0ABlzAZd6m3dqdvkwgZSKFb1yf0
YhIZyeXglPsfnQ9E3gAfmL/HmfrzFQNbmSgtFbl/UkhLUx358mwJPHALN4/6
OdS4+ebAjnv3lmLVCbGSFuyLM3VKcTaQ3IQKIP06/H0WJnJ0SIOiU2LldEFn
iFXmwckcnDZiAMUu5rOhNx4k+4z6Af/f7SqGC8YxCh9qRc35YKxD5Bj89Rse
SexKKnX8VA08vzNdoDtHDHCHJ8gozgRCFDFBdDyKHX7Oa4lUnCFLg8vYNo/b
uQ7rl94CgOisoYZiQMhBLcukrJYpsEzyd8XeTWzvg9astsHWFqHsVOFySFlm
1ChVrV7Q2YAG7xt3nrfq11Tu3YxSz78gAWI1gwFpm35iFa3GDRiPBjtp4W3o
ZswNAQdLqXmvx9GfLTKK/DyMsS/PuXTYToupvcsrSe7UEtmikd4pn/Rb6aS1
EUtKeyzqyc+lYbKhvN9EeVhhvowNdAAytEqdK30UmcYkC828sXNxMmKxhVBa
iPewT7YsrxvwsidH1BYO8EhRvRyUVnjlOf6GN//+LhriaNxKSd5D1UCJpT3J
gdzmjDUrEqJ6Oh6/Dywydh35qpZytCzyHiK0QY35Kzcidr2I7n3jDAOhjW+u
Ye4LNtUg6jaXmqh1pUt+cm0mOyUdMZ3M3Ai14GnMkMJFq31cZk0CaeEwYdPP
LXsihljgnmI5doczNZ4TlyqVNpoRY60JYEoJjaiK7PMA66WfH4Iygw9vl6U6
IAFWiTMGv1orIABcjF6ebtZVf4WSEX39W6SnvaTMKYW+lPclpkF6w5tc+YUz
0WyX9ud+qxORcVzQXbb25Gvz5oPudLTgz/kOgwN7eihs36OoIvcQNYVgO0w1
qbNqWcvPdSnZ7hmcoM7jngLHAWr6S8EG6MkTAaJGowlk3ptfhuPHtMg2F+2V
2XX430NCGX3RBiAvL0s0HiaQVPFFb9QD8nh1JyhrTzYbB7rKFI20OyhMgBzl
Iv89iuDxpiLAgCWORQeo3c22VkeO50Bz1MrunyJyZFiaW2HqOD8LRVEdvZym
Ys63V4CtZ9koLIqVQsFWVSzgOHAH6Hb4Rm9yL7/9a9ibwhagUPvFp8v3Zu5U
7Gzg5wGeD/Zbc0Y6UvUzxo1sbPi0OSjgounz6+UKgMZBMra9/oDFTlE+O3Xc
kKJnTZ8oCMIWMey9SMIU08zoX7+ri+5DiOwnR/Moar5baloQKN9C8t/5CKv1
jaOkLmBZQoEvMHmZBHxCbC9B16NgPDVMmlAJ1N4FtRTIIf0it4zewDm2q4vL
LdTFtsKNeMOtzKLv/hGcQ1c/AxdnUV8lzkOp0CTMJt/A4057fBSm0WRArjNu
KgNVC3RkjUgeXLDlaxmRJ9uyhlevvB/BECr0EAYi+fhPwwA9csR2FCXwRQxH
ZlHCHMpI7lzCzPjqOGExr4t2pnEv6WnxRXOHZi7PKJVxdQKssvfdaBoQMlxX
mGGSRmgSBIzbd9+b0F9q7ADcUtrJT9BipNho2rWvWohvy9v5ngwz4fNIqWx8
G/+H9JJTbC9hdgAsD9Ht4igu4jnHlRcWjF/waLgVaTRva2pDRSoPVuyYJtBc
P7qmxIHMQnwpJevYWRuzYbCjfXuaPZ49pTBOxJ3FAV3cxoyRKFc26qpOmONa
mNwxdtxzSvjOj6HFlJhkqNsOypYYKLmtp7ROD1pJ5MRkVOQscIw7FFB63TLE
2JEJyltr4mpg+CCZltwLwQQkfdlvygfNs0wDNoOe71LdCqBezBtH55+eqEkj
0txfMY6ZMEOi7VIC8UWBjl8awDiMyl0kzxRkzsOUNSItx2VsBCe8JmQ8IX97
Em/yzZPi78amN0CmzxRQyHqO6d/DFwha0YB0STvMuLHmiUmUkWBh2QYGK3qY
GgVXTqEYhfIHKZAguThhJMzZ0A//mr3fMPWWZa5thXySzRIewuYD7jKzgxJ8
MNy1E2VQNkoSIiuwqLA80HM1vQ8KyQRpnFWKlo40h2gqkVLm7WrvDpZm7fGJ
jjU5SLNtFZUs5cdQ2McAzDA16baU2P2oYgB9gY/4YzLOGjRdSFSzQ1Szzj6c
+idb6QyvrZfTg109F1BV3JnoILJeiXMkyFS+ugHYmszieUld7YxAtD4Yr+J4
Qmc7UGpp8yvckL6t4gRVSn5t/eyXyW0mgTzQAGAlcgXhCmx5+0LSXIsaTPuA
r7Tj7a8uCv0WlJ6cwcz3EUFe8jBhhPSw+p16ILKpAgXt1UfGm7pIhg9ldYtc
0SdxdSdL2NFOZ07kwAfp5uLEHVvvd5xBNlCVmqZPigimxO1XSmXEEo7u86kQ
HxNPyvSMRr0N4C7WEvzdhIIoOPWrUPMI4dg9pkAAcO7o4uhTWjFn+tP4Zx+s
czBo9uICfiLYgfKBVQzwEb4tgbBiBq1m/Fv8CUO3zCQH3fNYcezXgBs6eccB
TeudpdjxYZvdoSgejiFoTBM+iftPZgY7ZqqZe2igPNEdt2DqXgLmapU5QuOZ
pAlRfxMHJ02WwWqqMwQ3jKwDAE+rRi5OaDsH5QdADqN2FmR5CwrUlp0cPIty
9nlLzFDBz0QRig1AXimPZcOxrr9ds4skeL51VxRtA7UPcns8YUrIJYp4wVwW
2mLIC7J/1S+UcLoYablRsekPDHg6qOHujYeMvVV8y6oaAk28UiNX2sU/CTed
2dFsNf5dulSZXvYA5OEUOPUFaK0sIQWpTqAks/3nTNMEO1aFj/oA+cODo8hm
mk4gIGLOakXmqYPZsYgqW57nB7z/kLFf7EGrE0YMAJ6snDbBSOfkJlz42tZY
qU2fYLtUfYezC48gwAltY8XD3w+/gBAFAZRreZjfE5vX5PaR/PS5dfFQxE/+
xvq9yphVzIkrJQbcw2q3wp1rarflbP56VbyxU8rN0MToHn88sGh+/0q2AGsu
ohHoHJfyMqEv11y9JCpftsYTPShrZfEmHUt2rx4U2eA3VBe4JKKMe8uygCRo
Bn/hxyGXWuy2LZbJWHJA2wY7/Q9QvTkCLiK9W09+s1vB/lhqaIai6VmE4neT
RWGDsCNRxEe3IvhqsyOPM1SnRcLCyxLRenPyA/eT4VOrjTae1NVZ9/V7uUb2
IX1qLTL4RZjfhyklZl2m/laeeaqBD7+N+x+gVfb+oVWELvNKju9kIwVEUReL
fgkIUoGg26MSBux0/WagOKyliASvl6yseEydW+cxF6FE5b1Owxi2hqTMUeI3
YV2UHqctTp/Y0iHZ+P31sLvS9XJbul9fQrRu3xMj0gNIhqyxeKL3auli41BP
LrtVn/8lvIWgNltTDNfyC3j73bBsEmWeFkA5+3K944b/j2cpKYTDRCa8HVDz
pLuAMco6taeH2B6l0R5HYGEEV4ocQIQeX8yiv2OHAfPQ9rmLcdCKUbi1ejRv
wTMdPjqlsqmWDvi6pQb2l9n41fOCXfRVC/ap91YOYdmXuVTY/85WbzoDhecd
UdyF1pKExmj5CCxaq9EXxlhhU9WF/e2f78mRxUzWv5asEqforvdYSe/meT1F
jy7nxNbLJiHgnkf+kEHTxP2F8WQAna1Wt+q0pnz1oX571vX76iLA0YxnzqZ6
NbRteEPvxPy2bSFnEpPxo9reoXNvDB/6DZ0v3PKOBt0yYdcfrwo8RRYgRBUU
jYr4mwD5gWiXFRhoxwqSTnoKFzcKdOoNxZIipG7rsBgGC4tginPo5XFDE2gf
hj0IsUAKJs3ve5KGXkSygAD1+QV0t9Yrsq7FUhNTBI+WRrDDlp8RtgTkNc+V
r0/NGqUKwa3wOQo2hZPt2aaUS82UhW0d2xFn+vE4OxiGQjJVsDNBhITc69i7
753P6zSQHnO3V5HpYRVekC/LBh+bBpDsq5448Xydc7IqsuG2giFPhcvjZOfj
sTjDHJSJUD33vwhlishiLnkxLm2S3EjkvPARITWPSTshXuE4+lsH5RgjSkrS
4duJw4sToncJE1isHrnHM54MfjhiCSLQPc+XR8Vg78Bp23jyFqFs8g5MNfID
wF43ZHCWd499D20TLJ9luZhUevuA078ogmMlPniY/8xfj5G0IjqY++I72BZb
r1czVQlyksTk47lQpl8wxINpCml28pbqe/oyIoko5v/AsXY04LB6UEZcDS7M
hIiq8AfOQM2DjGWiiEV1NjNEFckKRODdV1jZM38ixEGGUS1ArDbKWrIjOSQ/
e6p8Az+eQeXEJ6slVYHOglFTNPAwtUSphza85YaifHXApPLB/aI/+qWFJLNZ
zDzXm4C6CryzY4NgHOwp/QWetxsmFPx8ZoJDilV9pTrK42Us2+ZNi1XGvcJP
0HK6c4IvJUKR4HK4uFQ7qULFisUtr87Br8HHFAsEMmX1pxDKZnh90y2mGVAz
3jnkLlYPDfgDPlu4qjP/YGWFXV3np3ApBdh/hYb2g9chqdbSaDvzYv+aI/9O
nIpRNR1q/GxduGc6TQELHrtMBG+wBGY3ec7k7M31eGNStetOqLryRA4ZMX16
fhz3AAbePHelYHllSTql/wRXB+QHHwPOXl3txwlkfFI9tPekFfLvNONua5uD
LSsR9EM9ANzt6DiNuX0M4W56X+LabetltQMuQhyAcc30o65VxNVBMnXp8Q9Q
vZ3onZN6/H2kv2BPfTWdZ3Ydf8MysAZ0izdu2nd7d3wJSJjboyRJhbdmcFWg
s9Q+dKz2FCoqmulF6CT2uKaHo2YGEY5UIx6Rmmf5eP+Pz62AW4Kl5NQEfJA3
6nS/DB3lzG2+vdBCX1uG/NiX5JTv7gmhSMX+WKQ/PGVBAVKZizLLvIA+r+kH
0MTP+ZXFvJGPTlPtGRcyktPEHNaJsZ88iYwZBjKWnXsZ1xvxuX4+nr+ySvCA
3DAv9j3w19fkNhUuu6lMAwoKrRh6RYlgh82L/tlln37CGcAUbrSmRI8KSNrL
sNEsSItZ73a76ESJzLQPjyIYMmGOS4O5gLJeEdAu0OtVILSVSdLmHQbcpwK7
C55XvCL2lvQpR+uVsl0tTONKrygHIN9xxT7RxzC2UyfDhPbd4CtgslwJ4sUU
F+1rr1kFKbCXHXGgCnxqArh/cS8sFLSkDRo85Ph+YPmLWEOyz8WqHSG0SPEW
uyHqrAABN2ft8+dFkPjomWMsVtVRmXjGOsxYh7T/ZAjPOTgOfe1Wck+pCYql
fHEq25z0PqtEp1WjGZuqTF5oxExV1GNKTGGBX+Lp83HsRfDSgSxe9ML0RgQL
BQ6RYOd3mc54HuPkO66YvIkbNMQnk8JbRV28+gxkfis5tmo9rgvOjLPz0Z1p
Ny0W5UiJ1F68SkNtvFTovDluWlFeln3To3OZ5hkPjpSPkg7jbZC/P64OUJrk
DqbD9ffHzs6ka9PT5C9krCN+zJYyNGUfhh8yWb9ky+MQHgYnB55Xukvp3JgY
4yRL3wkIT9dZDMz0R5toJVLGSMQV9radb4ov/PwumjLone7pcRpV2YQvPfOu
vEBRL555DJwaPkXS8JvWx/UvAaeg3iH2HTqIawjQDESFmu2uQZxVGJmxzjtP
ejHplrsWJDO7bD5HzP2YN6wfdY0KwQ6KaIIoWywy7s3Ae7BjsVBCw5H2OFhg
5oGUYiOGRQTem/oIxJz65YjeKByoj3PWpLqwuak8bDdUMX5K+MbJ74qPr882
i/Bxg58iT1SSQlsrM7Tc+YnTiO+P+qS5BBLQN2wa1r2/Q7U9kcdUfN50mJpP
5h8N69hpBGHZyT3WRNhy91UDd6rmmLdF4/IcmaA9yMz6fKtZMEYpFDSJePb4
8ZGjX1nN1I0g/JOjQ4TKInBM0L6uuvkdo7LKhyd4Jz8qjjYorWGlZxXQ9hQW
2KJUfPr4dNyoW3aHthsTv+X4rkER5O+wcX0DyLzkvE2QnRvId9vBAwW6v1u2
Swad34WrRH6PvSiUz1vn1gAeq/CT6GZYlssMRAoguqrqzxJ79w2vQe443Si0
jnrYDSI7BVki1RRgHhWvp6H3BLCzDPDRwAOony7YDLRJ6r0MlfY6iVQTPNHr
cuCeZXz7WFudme7Lp3VFXIlXQM4ZgXw5vVJ04pWqp97yLz2hFVV0XwHVH7qx
SSdH/yk1pvi/ZV9Jckc6xnaPHftQQB9TwwTsV17hFGukFDwlXXwph7uzvCs3
uje49T4TE4wMdKaQQwbqZuZD784rSYYJeMHEzAWxG34WmGJ3XxL4NoapEpze
EMHvtZQotVxWLF3kNL5zn3gzRTi/LwMjFNCwB+i/w6qeXdo+eQeOZN7sYQPv
3YwcsPuitelchn0N9sNP5o975X3nc2ksE+Mj9mIE3qJlnpbyd2lNB4D1PUJh
qr7Q8YZm70zfAD6PAyZnn94Y850H88d+NzD6Up6XyFiepF0tEhPU9sZD8YSN
MpKlbq7xRtyWQfTkmUnQeWrr/uNcppq0QfcNlSPPILQhV9I+tymY6idHdm6T
sSQnddCuL05Q0i5H+ZBbK4E7s/L2OCE/3+tkocQjJeqeYWb2eKk7Tske3XKU
7IQpSPcK1DDp5YMUdSK+m/aljb10pKzNPO05m9xi2p4OZJlIUCWgeGz4vmSm
J9wcb4tPp43GmBDGK6BHq+LMhJJsWPrb3fx6DsTMuXGHYGPHVzOTsAuT5vI3
UNiNCQvdRQzbUpslxaAmIInVP1xe5ugHEPrLAhORyAYPY0IGOu5U9tSXTR2b
UY1Lf6uDZ5ZrUM+0mMq5K0miMV2jfjihF2/IbIdF+DeXs0dWYxQC/4xXXD3R
O2IuIFrBpxm5//8Hbr7O33upwiQ//b8Qrd6B+gKIRtodxaRTymiT7n52Xi4R
YfmLK7JZPw3jyACFFwDLYtnQhiZSdXfnRWjPE9qExtoelZNOcvO8DqWn9MYo
DfcGSlIV/X+T93LzXVFkY9cZhA84ZosxcjSnniYNocIMRvwahYJiUTP2uvJn
kvSed1bnWQbcPavLpeR/KdpAjaqfWpluVlDSduRIeaJIQvDCOm00YvfwPED2
XiPe+n9LOvqFI6jSogA1TBWPv0wuyZM25ApMXmvnq5li0gpki7yDw1MjNDZ9
LPE4UnVTegl1WaTEza+v2ZiD9+/QEZ/3wVYXFOefforRIknIDjUJ1FmuRxzm
5iLQUKkPHVGdLxUuw7e5xzwQH48zQgYfScsEMWb1mzPSRySvEYzrjsFEtxDe
Fbz0VJOdIJ/SsChc9LpCkbclTu/h2Uyc5VWUz+3J7zHcU3hKZA4TZgGF4BQP
Un6NhqmZ0ffoC/xNCYd2arLu/2KZpR4vBrkWr0lZlNeWAxdwyOQ/hlhvLGTg
ikbRaFOkcHjg9ghjIM9YdHBFWvz92YTZGZu4wj6B6qmaR7sHTgE2poQDV3dZ
JTdF6aj+8by8rVpVZ7x301ZKY3kmOE0iUXnb7E2MgIJNct0SHCAhCOEPSO3Q
8y7iKq8Z7S/TNRv5RjcSDNseJbtbrgN5UiTnvMCpaS/eeh9pLNIuAPmJiDRM
rYbGjFFT+7vw+GnfNJC6ma9RPKzdm8mKdx9811BvEqwPtmpz1Pr1wqOQALpJ
xdeIrUQdNYddTuSxoP2nf+rX21LkMA4b9W+ps/bhvJSLkq0A6g+J59nXbd1q
+rOwxyNi3ePitY24kf5msqR6btpSWb43Fsz+zE2cOuRviI6UT5BS/sybTLoy
+FUhnboJxmXvBMgXnPGyUQ7xctS7fQcLnKZpAc1629QskWVr7kn9NSBiSREe
k4EJ3FcvtQtugzJSbCXz/4jjw7PudzZwSNCsA0XAjQJlNIbU2VUoCg6vQo6M
hy/OaDokxEQKmIZQGXiAYBEOE4q8zPozxC2nvWPvKneg0Jxd6A9iClEnvNo4
N6Yv2Y/WTe+DaYK/7mqPmbtln+qqsFMQASxCowJEyshwvFjlt9rxIOufuRSD
bg0E0zuj7PcvJ6WdAH4DlVDPhG5LcEjNd5umcq8DAWzWQ1C+TXIoysvq4bnU
W2UYUG2BY5ijWlF5b4wHE44Zow2Gx4yBJgjSfxWe+vUYndxAHRrpl3HHU4JM
KTSk1DvadvQstmVJNhKVdrC+w+0CgJBpPbjy4XFMF16B0LiHjDT4k334TuC0
azNY8Cyzm7Evi5uC+vgyUDE94rh+AYUFgF9ovgoDy/BtFfiY33051eF8MTWT
6wYCF+4nHqqqAC7q6cHiz6XOIp1JACunBtaVgcuikCIfXVLroU3TuNrW4sKr
ZosnNySslK9rj2sr5WS/pvG3vSDiXJeTBGQ++HnE2vhcrqUFy2E0Q+HR70ow
yotemM8NshfGoZVSHYYFaBAf/K8FROAea/840xWiIvAyRYyTnUo8UUYRaAqx
PNGz/OWa3fJXGq94/G4h7vo+mG94cZ9r1TIhs6Zttk+chrwOsVA4iPN3y5Iz
mP2khO51IEnOBZNjWpsZ06N/eIHb6Tm16d27pQoTQDp9Awx5NFXg0s38eIbQ
RR1pLK/6pFMG8Iksc7UF+A8wTSvx1t06aurZskdjLhRCAFPpf07jQETb9wx/
RaJPyrpabzTRPucxLUSxCuNB7Ps/5gi9CSeNjgl9GYpIzN0A5U7DOoKnxAjg
LSdJlwg/AJIwF7QjKZoBnT9lG4rR86x6zJCdhIL9Db8uktkczHLW1mMD2SgE
65pxqvbzjX88ZPRrfwrfnIRlKFK8aYPO5DBaC4znhk8Vq7HT5NOBq9/XWBaN
XCnOAcFICAoIiZsMy95GeAvwHZrIA4x/nfb6VBB9vhwEzaoqY0uCZ9oJ4gFM
oeLlLKlG8C6yyeEi2KfSfhjqceql+S2ktotBAFrxTW6QeUcF+9lIyMFUk4DK
roFnzYdzybck1D/Rp1HARTl+b6fVK0h19ZLPo0PGSXciIWVnloVBxzbTpz6I
JrvfwvXVYTiHDdxYLjJ2FY/BfgNC7T1BBBW3bcPHKlpFRVPwzXMPeC/2N+7b
NF1ngXAwMzqDXAN7WW0G45ZKVdv5QMVWMVePQ8uCx9Tp5Y1PEc7augYA6vDn
JyOSJ5AUovNyd6wgsbm7zYS2U7bhr8JuByUyll6+cEBF80lBNKYpchl3xGrJ
OWY8X5IG7CLK9TSsZYhlreqD/8qK+c8BIAdv07VEuT/y+1aaOzagyt7uEJjo
5XTG+oo+F6YwKPkR7pJuqQt1nLz/uaIRqrmVKCLR05WkXWri/DwGdfaS5tO6
TuGW3FuYYJzDRQ41CrdeFwI+H4ox4vACBCd6l8mVdTRHsbrGw5lMfE3VoE1k
rWA8mILHFwZFaQVO0+xkUTkrncZZU84pjbppsXV7HDHj+3GP/KF3Bxrb7pnw
/x3B8n1g/uIw2NZuaeWxyXEjIKqCbtKhO+USSRJ/p5a14F8Gxyse4EdvH+sR
0bRSheYKlix9+3xHuf5U3Oc12fe+6YkGf0Xn+nkGljUMN3WWk0fBEqpbKdYK
PI2JRDR9OQPup9Qtn58Yjvptage9PXjHGhQTV/TXEcBo0s0MBBOzH2LBehvh
FcxAo4oW4Ne9frCK0rCOSWN5g/tmoa3KbobkFn357sB9fLO07hkwsECl+bfB
5J7vWGdy6rS7RW/YJh/OQOHQ9P8pu2/Q/EDYkcC26ecCU/UX4h0+h15hgBeY
MJIT7gbRQCisPtYn5hfvgdh2NHYQLp+Udy+uRCpTTDhrb0Ggqb1zpz4ZApUY
23uiZxSncXQuCPoiOilBCDB73K8UVA7oKtT2xdvVWlwJc0NcajAuEweA7nKx
sGYQ8il97HzWquZUrJ6MPYPT+FGOEdbdHcQ8d31yuvbUbn0Nv06LC62meDM3
RNtuYfN0Xy9Ar/nMs/27m/jAJWldFtSAShWkLjpgxXkGC0Jki8d5jlK/1XCm
+xtw866Nb3CUYFIkM1YZvRpzdqSaIOETGFZnSbM4a9h6GKzOvE6VANG/XypR
cITC8E6asquIbuExY+m3Z7VNj2VW7xAmIQovweIc6Nggs5wcDiPg/XXzWY0g
f2Ekq7IoGOouamEzsRdhBOK98U5Lzh3xoTjzZgmd4gZIknkKj1sPSUVACnR6
ocrvxSOp0903cPyBoz9cvWliE9s1+CEsCpDlViK2cJNoxyCQS0l/Je66oa2N
y4J8zF1e2Na5LQOnXl1nfstgCARQfjLa2aWIU5SuuqGXgVsiVk8p0hP/h3lG
ZkpnEN+FyvSo6NnSXX1CM24FrOWj1upnI7gziF7kYV7JB80tqiqQ3Rl6xyKK
KYmofVxGdq5kpZ/jYhY+wwj9n5jMtOeo8isdQ4GgOwBkiuyKurnfR2CUcRBG
te9k7q4XMBtBeQtpxeDOtnRxUXlEqqfE39jegdmu7mVFJ8IuoogNQ9FrSi/I
bmWWwA7l8ejOgL2T2DI1FQksk754FnjMhv1lZKJobfRdUL0Lw7qj1L3Kyt+p
9o0yCzQtD0Fi0PEAVZ+oJDorNZGK6Z4D8VCglNupet9HidqvIJ6THaatCI8p
bt6dTgmTdhuf8mWoltH0gadibHakdfSmZi8iS38Mv9rSG1Ne9JrM2W7WEO3J
WUH8jfrWLUMreUhfqlOO0xBIYCj0+9V3FbXDRJHjCOry2fZkZtfjBRg4kEjx
vFwJ1T3URozf7esZCn920Aoaflvec2U7TvtxqmF1fQ6C7qadfvw4HGpP+vxo
1OtCHLkoI7Nr4CHDoVZbYh5Azkw//mNg2sB98htCGs1JzipMpV4A9as9SU+K
zYa0j7n9FJDkS+Lhql0bdVeS5CfWTRo8X7ZYsX8e6wMXjVdpl6esfluHQLmL
EDdOH+Jdq6YSZx32Y4Z1CR24Luk/Rxfl3SFSLuepxYB0fNjMums/z1ZalCAg
5zO/cljczwPsu4lsmjR5dac6+5H6zXGP+KV0GaRR5p4/aaWSOfMHUVXTS/Yt
X0tEaoQODemIwQmMs1eSkmy/+Gk4leI7vMKochYszabWnhkW6Z8kyqbCT390
6STHEKWUWrI0N55/hTlrUQseG5k1O6ew+4aaXZZY3kbyJKYXC6Vx3Avclvpe
bwSXG8/pHAkGS8NpjpBwhbcgHzrAnDhYxJ/C9tgqPmFt7I5qJlq1uCFvAse7
xIttCbiw0+irU6WKixnTZtlwoY+IRieQNOivsWpcLwmqReaPe76Odj1qCOLC
KR4aAQag/1kxdtIiCBEFvRcPhiBBK25rkeKf8iyOtD6a3yaf2SJP3SLJQu54
n+DmTusaERg9O5Yj+J6wrwY5+Aw4weUfuBRaN2h2fCZwNpQCx/U6Soz8M8BR
gB+OovxnimESljQ3gt8A/0gUxqAwV7hmQfREU7b9Csv/PaXzLyvhs5sce/Dh
gpl9/e8xAsY8526+ZIypYUBuUmrCxB4lMCrQiwca1rPnwxk/vk7yARpaG3kq
21KpbWByt8BdXhSeZB1ERgaWfta4RysCjrG3PA5LVzjsQYqQ4PN+Vjb++QF/
NW3ade0JSTP2ZJbKluuMc/AIlbCZSw1IbqZ+LDTTe2a7OxPKRzqCPriAhZuO
33b5ATjyZaPZwspkP9t4eBOvjGufZ7OSZm23A6jZV6CSZNHrahzXaumYUM9Z
pAYFr2eccce2iV30WfEVImgImc3+bA9QIIaEEGZolSbPBFeIPi8EF5+aa+lP
U0IHaJAM9CIfjUMtgr8xbw8I0pROGLtLhMCIL5KH3NA8rGXa6s+M/WhEiYFM
vKxoEfqyRyByWLHTWcZ+QjOxfb9cFWRPgVvN6I44To/j3900f3bf0bhjr7zJ
lx01Vp1ZupvJKusE5MLDFjzF1pVDnneEUQp2vPOaSTaJf0sLKZOeUOW0h1AX
4fpA9KjfB1tHT+QHWs/dmVs4XewtWojKBtjugdJ/L/EiF9Ioju0PXYw4zPbV
/CobheBgLqcbR4sA7wvdZVwckwXYwP1F3whWCWHFfO0t2Iu3opmlcFe4EIML
hwvRUccOqWbdVgxITg9+gMubSH0uj3VVHiYyrjqooznLp3OTLWAjHop6ihsG
poHU7uVkTOqX0nUDAxJ+d1azW0yv8q2xDD8O3K4ns8eFVo0ytiyPdhYYZc6w
lrtbZglXGrQ1yzHP9nCRQ8YfbGjG7/n1V5apcEUFK2yFhBH0FFBGT9vEJYun
ILOwXWnrNX5AtD78q6UZvglA1zhg2d55n2FvQiPttSUAtThKp94nPpZnxJYB
VCYKBD/jw6mk5CdsGCg1CL4M7Hf8K8Qxxyrzg9lSXDTCVjQGJhVXRd9EQ8pF
wlD6SJc4FcaFk+TlI2SyP334FGtq07uyUYo7eBMbwS1oee2QS0T/RGiaIuet
iHddmJJjXo+PLeZPeUzmhptE2UY3M6BQB12GfhEXgETkLD0Ge5OYJHJ4ZrK7
YslZGzXERnn8/MKKOZfn1yLI9OfM06LSjaZNwhvvHqfTIebB4DudmpdSnkYx
Du+Lnl8h4P6+p72eXzFraowwtbVfbZhuSFDdnUkTFPwAc4nssDVsmRPH2FOy
fMXhprWRw8AIaMi6a5cCFV2csMbqgp4K2FHJD8OEzb/fSxN+/sgH4hHp2qle
i3UCkKGJY9jeM4XUXW9Vf+wYgGA80OubSL/mm1CF274rqp9x/bboALK9gmDj
8NwhQMYGrrnMHod8QmYHEcXok4Y64Fbu86x9O6jE/lG+H6/mdpGVjZDjeSLs
LJcMkQ8FACBoQdrVWXO8xXcxEweuyQ8HVqg012lileg/2b4hm1yrafCoAsSd
lqhJaHtPrG9bsIfM5fgRF3Er1V3kB9cyA+xaI0Vbgm7ERRO+7tlcqe7T5L8F
t5nM84bvm1mO51LIrFbFR2odZ8NZ83AGMmg2zSxjiKtZz5E6aVHoteoRzAI4
akIdgIHzuweFiQxNqGG+q7OnPASoj80SBajtMbyrmwIU8/yu6IFoFq4KlR5X
RxAkQlcBVlyCp3+k98wP1TQmkBOzaqYd+PIDmmRHE1pco6aUMq7AinjgDGqH
gAihuqi+SrJo/T+cfzP4wsuo7Q6GE2j/yYoZ+xH7z573wxMUf9SmGVj8WEZv
luYq1o4YHlgGxwf3G2doyl/mPV7QBKrpgkgFN8fZPWqHHPg3SlSHFdIQwkmJ
ELzli5lxE6MBI2a+d5M+2Hp6yLXw8ftqlaP5UduZj5PysPyaiTvhXDdoCjDG
2zgP72RbZ2poaWlwgA8jeVT/UzbyOom2LkwTzH60MijQLB1RALZUPDCQCPuU
4+mVo7n2wB8zmLxln3OgiPjnz9rBqbZUfRY8nfKKAOsJy302PN+CZZtJ7uC0
LNoHOpFrmcW204mh/AKejOdWnHJRU1Oraz5qvpv1fbUu3tKC7q0xcdJxmQQg
DZzD8lzuKZb8His4qy/4aR0LleO0V921fio3bNzNqWt7Rz2dhNcPXfAAwkuI
Q9bjXQYarL9bI+GccEbhANR8xK4KJBVXFIdc8O70JO7VUbeQmpYN7AwbmJGX
2qrNZ9Nm8DNhkES9t532ObuSMrfutStdonTHNE/5aq3KocuqkgLojBt21XYZ
av/xrDEayIZNod5DK9dKA/24PHqqouittUJxO3eQaMZD22SQx+jE4zjzAPTq
KIBDrwd34RwtWR4j7Ga82/Mwgh8V1Kpt+ebyg4zaac0tASyTkC9kBpj+sguQ
+uqPgjWLtk9J6OjBye8Ih2ZhFbIjMxvSWz2OKoH/9K6ookPI/ovFY5x/IyPv
voOwvLODvwDvAAlKfKQKpqmOqDl5yShWeFnMK9yPKE2Y9TYOgYhFWJK5DiYl
7BfcGpDNQBTuNy95L6scG+6ieZvZDYY+rbI0ZVbzZwC+fYVi6Wp+CYmCybnm
xcBfSfwCxa+9KPaO7YGrH3CIGWdgHQ6JsfNRHgx0r/a2DneH/S/1C/KAV49l
VYjGzkZzHAbneB0yPIqgWWRhW7gNyAznqvGMQU3h02e6ndIZMooXEpy7Tl/j
d2Ki9acaePryZlhYQCWeJg18miXpn/MeMs5kwhAPO51ZbNU1VjvneX95Nlr1
DitkjD43wDYlrGbmhrV+AG1HIR673q8GtzqmzjC68mXQZmd3QBc+ghMnzoEG
w1fs5pPTVcfGOyAVl8cvja6C7LluDPlEQHvt5n1LOrRifpl8xMkaxhf+9u5a
6qdoTGL5jW9xCfYI5rfD+Xw4VBqe46GXbRNj21tYIBvycMQPU9EAryrK7Sxy
RUO0Hai4WYDfvfuBMRzn/SfJrsiIPnRcUPUt1KteEhd8z8MVGPi2AaiEP2Ba
ATiJ0xIYTlnrPHt4yD8Ak+4oHRDgJS1BH6Qvi81fUk3rShNUfiC1PIePd35i
ECoWTxqDWHz4vSiSxetLfjaiKramHcfnWjDJTV0kHUQzFgq9pNEUOVxMrvK2
AKsfO3LhQ+km5cVqlv4UzkaNpvKiTX9O7XbaBMCRrb8neakATPPlTnPeyuq5
3gMD9G5PYVZFsiM8Y+M4I+ng2DlCdI6w3ae0t396EoAwHsXjqlQN0iZJn9ID
kbCwi4DUrH/5A4JVjBHGYBSVdjKP+K6q9m/ppITVlFP5LAFzMM5fRIN+51IX
N5B3qJ3eAKYGxJygyBWIBsi7fYNunR8wQ6EpreBSJ45wEckGnhgpGDgNkfxH
eS+V26j83w3E2LFSjvvf4ltc0zROkuqn5gnVlBj/1Wbp+kxdua8affX8vINW
TDC7ctuL4qap9t0XAelDKPXgrXAbkY06vkivu3hMEBr/jiqSRA6wGdhLKp2P
qYupasEmzR2A51rVhDZnnQWaiPwm4+lUT9zXexLZ7GVQk+jzp763avlR6o0J
FTyafbi+l6X67pszSJLxGL3hOfMatNt37Dz6QxYrp16+vNEjnyzxFk6t3U9p
wT19lMopv07q/XvC1rzFuQJvm9mpgDSJzYTGOzjIkY5ng783hLVUIX6m+wOo
xti9eaI5Gvo68rMWSZdrwe5uITFP9DZb//PtXEJFoZfiCiLXJGaPoELjcnQt
SthZN2hG9SdnBlYEySsG/IqSSUqqXv64uozcWOAPQ3jJmUn38gl1rBqt/4E6
/rFisFOB0JL3GvnW5mfytJC4x+dYnhlhEtwQUOUn0Wico78O9L9XJt34XBxx
Io+LMK1LFMC03SbOmCg5GYZ2R2yBsk7iyXypYx+kr8RVbLGm8kRzK5+17ziQ
DSS7uhG1jwEGwV/EHoMyhOp510s54XrfzI0wFZZCq3XeRR6+5kzzHhjvldou
K3oY9FodYgW3LmdQs3Fx5IlgprCAcwKkGpphyhtrgtww/i9VFEA1p3+ub+d2
TvgnEni/Pf7Lvjxx68Ni/cacZXdw4w+Dw2N3Nd9fppI6XkiDRA3S5FJZAa7q
mR3nT0jXQQdL8UAAjNVJGufBsTy4ZPaW81dwvL+EMvNdymM3lvx3V94yd/ba
48pJdA58P1mk+VHQMJ9H2V5y96dacWgwEnTXbSIank4dE3H/uE9z9PfNE9YJ
UQJrjFvwjK2wZ0Q5C0XbKUklbnZSI621U0zYBGLf2tEM1veXIrsRhYFK54qT
vOercE27ug57Xlq+WB/UjR3ARQ1EftIqNK+v5D8H9tf4M1n6ucQ7y4JZ4Hqa
PUilRPQJeOYgAC4HqlNijUvRqjG2IMCoM+/jOT3ImV3JukSkWOTk4BVOqNDj
fbqZiknHdQMNv7O3nLKoDenJRHmW6QJyyi/iJpB/WhSxOjRfLgZR1CB1GHnQ
vgaDx3pLRsmAp0XwsDtQhzC0d1l2+aFKA58QFgNqkD3qgJz9TDz7tcA32eAr
o68PdzLD1bIEPiwFpC8NmAD90+7y7D+tl1K3Sy0YcsSu8z5bb+RzZ5blW64H
TFxBkvvcsWRgjbyd/u5SphHGCpGsdvzysM6dhwwSVZL6p6qtvTUafKYQBgzr
xOR3tvQiEzJi7lGVrg9E4brLEdE6S1H8UtyCjfZepp2W3OmDz4JvDbKBTbmo
D0qObAPqV0lNrxLVHkgi9P60orn/xFKH4QsQS7tFadchXBLFqfHNcnx5UZh9
Lrw0zGZnwmLmqBC5Ei+23ofLnOCWcw8xD8kH9oHyOsjcujJQDBdI4FAhk7Uy
mru8p9oNaPkLUgJw7WKoYH9VHRJunetdNffVnphOJFO2Kas5CRY8ToDmE3eO
yp6N9vlAbhT9PFcPh3OyTAwgmnxqHRUXqmPLbk1lMA0C/1K+yXyJihq1LCFt
I6UWhIJj2J74Gwkk7eI2xABUfF8cCO8y+ihfJbXHCFogNq/JNpvjeMwL/TCl
072C0T7Lm+y9+GMxGPmvmBBtl4aZimWuoYoZhzMpPbaGBk0DmFhYmZPJ7/p9
wPWY2KkZYXpeDrTNROahPNE75/mmbK6zzn6UpJefOukCF+xUaRlkaEN4+t9A
K/TReCrgSGrM+3cQVGVCFCjuOs6cHzKPsy68VEW1M9atSoUdiWp3+i6OYERw
8QWTArJXbFWObXX6zN7eowvBjLY0xaF0E0/4WxjIJscaxlCWTfF+NAoMsgqt
WjUPyR8pzaDQ+LpI/RH+KdN8OOnBquqPwFls5UTeyqVWt4MvgdkdfrZkNWN3
MFDTa9Hy4hIQ5b8NScnumipI8AZH/APZHZOcvkw0s1KzhsR3C5aMZF6joT4u
qXc5hJTR3C6jKNMCpLMF4D7A1zxg5vSSOjdr52oCai8zvfciCONC5nvckSVS
Gdmih8BEQjKtedAtcwYHAYFSV8eqMqFXbTok0mW7stntFzGzuSJI8bHbRAtI
wbGM63YnY2erHYpQJVevHkFrcf8kcpINwVg6nXb4YsdnUL8XWHhkLgRH0YUV
EWdFhTlmKU5u+lQAsIJzle72VgZSvOqZckv+VoA9MDk3XS91xU8E2U83Z46N
v26kkDkDe7xUzwEAzC3g5zt7cNKZ9Qr+flDFDzQrv8pCoXDzJ1RYDl3m4Z3E
b9GDxdIrWX5yxYN8X3VwfjUf4yV+28jbHQe+znfYO4g6bY9n8/w+7sR7Hfo7
vaMf+/eInveErK8tIcrZJk7AnYz5lTUIBVHsJMeTr00TlD5wwJlylydB5x/M
7cM7acKOJUyIZruKV2mtqRYPAIvF+i4Kgpaf6gxeKY/AWX28K+ZFyUWWBFEP
B0wywayq5mm5TfZMXQbYCVVeDESfEywwxntkcmx5zTeijjGUbj6zUHbpXz9T
YiksjQ/Rq0gNRUVXH+JGKcrovSBa6XY/Tfct5cNHYNagrLoYw4+l6ktr6Ymn
xVnUO711xlwh+0d2uanHWdiNMALiJe4G9xdJAj2EtVDBKHYcFuO6demsoHdD
ENnKj8cv1BwvAFSMDJbLfipNsdArbd2qm6TqQpF49OFHDjGP2pnyCz+k/rrJ
089twkT+4fPCow6mU5jXdPAefdn+O5klaMbzsuQzHm6hfJaekelUuBx8Uk2Z
wmcRK8/ySqrhX3j1HeFzq5NTudrXW/DIEc+hIDXbzpesezRCcWdgVkw/FGj1
OWxPH4+wlL3WkeU9ZVs+E4JDgENgN9Z4a057c0a0SPC/+b5bGFLIGvaDv/7Q
qNL1/5dj6ZpQHzmEWNelZ+M2k9FO09k63+LbKMSkN0/4VXt6GwegQc9nlWbh
rA3vCTofe0EHcyUwwZW+k+O8x9JLUyJ6h9veAaNvLsg5qRWGC/3/cBedLZxs
Ym8b3CbB8BtZgPQBh/06SsnjHqtlRiRViEe4YwLasBWAMsNVNFrYNVtv2Dqr
ZA8cui5WZ9hjFQpW/IhxLFry5iWDLxfc7NTXmdBOVf0KNISDlF5jSzSUn5B2
CcES46l5hOTgZGMJGbq/XdSkbqn6aFnyRxLeXhUnPJMmWJ3pAVnQr3h93KdD
uvYUHJ8FJA0N8xSWCc8R1UoM+jCvZq/gMe1ofhs4bEXUZMwdqam2pWMwCBNH
lJ8LzsQb6dxlrmYkdbT9aZcJJDt0ssHDj7fExmQRNoJbK1b6mrZwA1U3uHtg
cInZDk2Sfs/2dqnvhseQDy3Olt3ZVZ4lmtP94pG78zR82ZVG09vYdYm/tmkh
FOCsfsTCJR6ZMUFXBbSv+XJREgwKyl0gN3IKJgakpg3qcq4RaiSkF64jkptK
ucpnWJBq3KRmcMqAYQkPDWkKgw0bfy4MeVZCcW+f8ZufIANkAuk/kMyf2Nb6
wPwjQ+j3eNF4R1fjTdPA26zm2gVQ2UrP1OQlwIum+pcv2PxqcrXSpPlijZT0
5NH6QffwZo2GGyksYUDaoC8MNaEbG++0ZLBxt3jBVy40PBXUrT2SA1WqoCdl
I2ERvwLHKWjxzKvAfjQ3TsPeDDqS2P4XU5sdIsCGMpoM759ImS6o8VoER0nB
WuclNXq5JNN5WefQIejA1bXG6oimR/23JtikooXjyQzHLfoGK11Qpe5Cu66x
yV0nnEI19reWCsgL1M6zWsvUcYgHpfzEy07iyKEstHqzc9QSxJSiorGruI3T
D1qCv33nJ/j+SbhlKfBuDv3OhwYmNu9sB85TdYYc57oCN3grWSeJ4jfflUlP
Dw90DG5RD3m28vThvgDLNcPaz9Yqnflkcfam1RFL06knE+q73ppdKg58tA/b
b/LMQLmpvaYJX80s/Xu7hvG6MLzQvJe7M90oK5U9mHfiKSQ4SmZWthsYSf7+
Xh+4/IzKx5F2KfllbwMB2VHa3oBi6iw2uMFBD5SD/6EtRhrk0+5Xba1mqg2M
Jbb/ZBuerWlpXseuvPkqhgUU5H2FlQhWWGBNZpIfcEAv65r+XUgqAjYAwhUf
9W531npiihq0J8BPl2F4tIgfOvnFZj5uLktRAgV4upaQ2ECzz8+jZaCUZpWY
dpHBQ3fmakJikArK0IjiAdb+VMPq56dYkCf50FIiOtIjP312s/HCWAzsVazJ
80lvqU7NIa7BOsXqX+iHeX90ss+wY2+Y9bvO25H+Vdo9yDztODRqhgO+mKBM
j864zeoDhWIivqo/ARpHCjBKltOrXfRukvrjUDa4H0sxRzaiKj3uGjtzU0o9
Cn4OLJvnVuEOFG3422VCKxsgE7lfoVV7yFiOUkIdaBJsG/UttyXXCLFFddv9
Z9sNpNqCp9NvhywVI5bdrDvyIbGERTcGJ9wrml/DJIXLNZnLDEcjtk84Ruab
j9UHVKrSJ1mWVHNWk24XFKQ4uKbYjA2F5o9i5UClKVSxCV/ffzH+0V0FplGY
ri+1bihUagdAY1l/6MIxbvQc+Q3lX+ts+NQ9ZTJtTiI89dj4Fkaj4KbL8M5q
XrsLYjDLvYRt3BfD0xioF26nbd+f0zzvAC4sc8s1H77BIY1wWiSb4P98OEr/
ZQNmU5L4i+Jr47Q2ocNHc48r7fxApxErSqiXnTwCbNX3rYLSspJAnuWMkXTT
MHci5FGuthtxMFYA15nETrrG6K42VUS1GVWxE7rev2T1iyyWHuHqpf7iKlbV
O0IwjfqnqdE8gp7dyQpQhc98NtIHiBgDYtYLZUm690IJovU/3h87rtRCeH/r
IOl6IpOCEcEygDK/xNdXUqA86aBrmc5I1Dm0Wq5fNHFAy0U4JT67fsex28F9
DTM4l9nf0AINKYyKNie9uwiCDjYpQ9n+yQtfiL79nD6HWY+PXHDfZax6uSq+
FftbZVjjc2xoFVw6Z+Fk2U8At/qfElvZuvDJEDGkFdzSyrV0V9gkcA4yAPgu
A6ntGIigq0hZKWJciFTiXlbMAVkkGpxhMFNxDGHyVT0mJdBQIfJVrlvdisMK
OGRatgifxh1kY10ES+mShjLd/MHrQbxCv4iXB/Usumg3lzOhb1G6gUP/YOAI
WiGsgIphM4CXcrvh7HfP620mGwQUAKXksxm71hGxVRjOK+9Kal65bSs4ck12
JJKbG/NMXEm3DFQNEKyFIBj/Qh6KzyutE1KOOwwz66NKRSOkcQclYP8n5dFq
/mob6HGHwQ8JG81eWZxX1/hs7YTpSfUmEEcJ7UbsinOXiIOgC5nYVt29zzIq
i+mzvcBGNjNEY4fMvUAmNK4dtsWyUsMj+Z9Eu4CwKA+N3PC8dqbN3dKFZ9ve
6VMumHNlk9L9E/mqwrrTv6ianfMsu7wZJgkWRFWIta6S3Kz+MxsAzUp450/I
EJMSGVK7V2vipligfi838W1PiSqpkTJLRA+ir5+nwIANXlAa5K7safxOCWYD
P61zqCVGgwHq7pMeztaqkR46Q0C7AYiM6rs9DkyWW/A4rA54nDNlmdUFoRwt
gqVWfA1DCzx5lu2OT171N2nNOBw0MX4t7m6ANabEBHMow308U8Yu8hS6U1OV
9iXRTx1qeYU8HkIWE+o5Rool4hLumqtrPv/oPtg5dQT0FfEJ7wytYmX9s50l
Nu+K7xh1GfUEHKKPSjnP+6naBohPLKOQWU9BgR7HuGJyVLgW8SCqLgnbWD97
xRLY7EDgeACnU9Xpnk8RU0NFSJZvxsdliITm4iwklExV7ztVbF8Vnqv6VYzj
QzlgxP9PshTkAoZqWTQIdgUP3WOnsrvT25vj3hdKZhrIfHtFs7RLTQofrWI7
1WOQXQeiWHjW2LMiWmQqlcUV7TOBgCPvHT4COIvZ6R9XDR9+C5RVcL5jyXfm
G3tl5Jn3eCAX6j8rc9xfTgH11SHkoiG94pNfdIGAj8XMWW4plc3bc5Rz9njP
xhb4f6vO7MqEzXtjVdIzTw5v7RogTP5sXjYNm3lbdaUHeKzW2lDVxZpHqvTN
Jj8ch66p6ev8ikRlcEA9NOspawNYy5m8QWbloA4KMKab5dScgTwgk4N8Efqs
V+thoIxMvgDauYSL4f+Qd39nxtqOfRvt12MGqRQ/9fsvwusVwt/aO2OLdR19
i7wSyHTFiNzkfFW8YfqjIMytP0WBpk5cD0br+bQ2LVFhr5tAHzpuNXzKeygS
nKz181kiPwsOJj/v+3zHdp/60rzsYxN/TD1MbVKMt/UeJp27WoGNoZbr4U8k
jWg2ZiJ0ECk8vEkBBtJwix3726rvzu86tqwdlVIUsCz/1KxNftHAQNt/zF0+
NgIg+a2I4+yc4tz9OZ4jV+IVWSt/st2ALQNuR4zXV0XWc+RCe+UUiQXWi19P
Sl5mYf6NZdR+viw5GqeJLljfT9DdaItt4Nu3NzT6Ze5g2dOWoo9PluyU3eyC
gdbEiGztnzsVSJN9wAvCL6pCSOZgB+8Z2DSILMXfF+fALO558n1gOJZcIAFz
ygdHPXPm8wCIvbkCwKhr9mebTXEW+2D6y32U0UMu9ecVTFqrj3h44UBH+I8d
roMkZfieV32gW/3Kc/U3iw/ZsKOCIScbvYCDopoMMgC22lt98SzvqPUYdZjs
JAbrbaX+nP5vB6l1YSXXvEOMg2ZjMT+7enzseC+oMtCnOa5/kxUMM23C5pco
RlL2w4ahMzyzg8AHjMdCn8sm/Cf/fqYj0IwEUtBnEVjFu8Hnb8nOWnXGKs9k
xnRxwI75fS9nzJJ0mv4/36uwYmR1W73f0OjIqgFWmHE4xGwpoGn6TyayG3kG
RE8YRlEbGFWudjrOvfLPstATFGH7k10TfDqX3WJHx6KPHF/HPzAa02AjMOIe
/CbVtXptWNe4ZX2pydfD3AAUefKOiecBQQCXKc/EfwDRJJ3TVowkwMNC4HMT
L+n8IL9DIyx843PsXngVXc1vHCWpQ1doFtyeqpUMDmtfn+K/DLxvlK3isKVQ
hgdBZhOVhgOhiQfRh4uvIKryo21ultbHBZLFeY2ViXtvOHEb6oZsGyQd8WYY
xJplycu37Yc2c2Qre6shuESqqaHX43rnlwusRSG0w/4/b5nC4sqYSkSyz/74
sb1PwGA1G0gJK7x/YOTzTpGZ5j/bR5r/SzX8YC/nEwmcT7H9s6ojeGHeSxg1
5zSlkOPRBqBur6oJGb0kQrpNQt3kDQSJvXw+1K3ile0TZAW6WXm5hXQf+9Hn
YA7GtpTNmSQyQTZNaTU7XZ5Ub3M+oYZ5+ZzNY6akvV416m2c3CUt3TOwlaF+
Wh1Byx8DpgLVCm0PnSXNiVVV7ceGQEEGil8pv6iq9plwmunLiqhpcbmoYJex
x9BEWfXi8zvZVCpYuOZ9LZ6Zsb9JpMAzEOP34hxLAG81dO/z1FdWUFGNFmxE
ZplUDo3c9DNScKJNwVo+ytXnbOY2mIkrB53k6RHBUwhUADXpDCSU9mnE6kKK
dvkHso9bI83Oy4fk60ZH0GgDHIbaKKvca7O/hM7WKkEziB1Q7XUno4QFeYV8
bRcjJHrrwZS/0lD4sSzmJyoVT1S/HsyvvJ4VJH3kW63kYkkgvzvXRZZriHUs
5FquaC3ydSPWgw0493KLNNul8x0BO+n/njslJE5zrRu1YX6bE4a7n1eI6SJ/
nxPLXCBpy6FBm6AnLKxRVXOirKTW75+hXBGAaLUnpWfjFowuLhJujcCY/CsV
VXAOipPFsMZoQIhIbxZFXRqOcwE8seWa1AYpAEOih6xdssm9L+G269LF8VsH
jPwmB6xL2a6cZWulRY6G5iGMtos4NAa4EcWq910jSv29e7eNTGgcKZ42iP4j
4RJEKTECuKz8WoF1zAisAoZSERn4Ri6K8GjJk9uy0segYNXN5aFZL2v9UNUs
T5WNs3HeFVQhIUvMRDADQR5bBBOi3qluFYRShEYStQ5cnlVj/IgqwZQbh7Qi
4BfzMzuI100eSxyxWUyoMYQYz6I76KYKQKPMvebnbWdshGatgltV0mwt/Tan
yWaZkO75Uflq7K9SVCCN6qoGZ1cMJ46F2NDEGKUdvRjNZnJciIxBchPo+llX
50tPQKsiC+cNZLYSjTLsT0xLVUoJ2vhRGd1miJIqDdGK9m8n7EHUu1NfwYfD
qzAEm5fS4zPcTZH2/70TnEj8Mz9f4vaIh9wNvgRM4SMxmgUs8kniW7hcx1nL
ZofrXnSI/5b0oLrbVymp4GokAo98rkeVhe/DN/4CM6hOrkGiVJwjhXw2n/rT
zpt+L/Vv4pN8m08AkQRzXzHKvJx+OGZmLo+OQA3DLI+Swbc44tOO1edmMK3M
tsJ35Z8KeROHp5eREH7pJd3WALxm4nZ74CEE9PFBo/SS3HcrhTHPxCdEvALn
4DwJB9vPwB7pDIU8mJEJBhSgP4rd3COPdjhrZQ9YAqMFThKNgotQgivk4QO6
XckUakdywi2qOhWo818ogIfshg1ADIgaejnmQhA1FFaA8LR9qRerfG3XOpW2
oype+ySLdQt4SQ660MlTggWZWEr4c1p3o5kqAHTbFxRwmjKdl+AkikeoPzBP
8nsZ0Kml+G6NVEuBTLjfHg9bGQSFZb/N+DZDzhtpZO5DFQ9DCxhb2LZ63Wb+
UVmgKphjXhIi0RRe5Mjd90x3GFojT+uvCcRB72X9i6IIB0cM/YC54zZRmrp3
xwRdMQB2/61zgpyG9mSluUD+XSkhAHy4T+OzZw5WItYAskGNxFz3EGg/wBce
YGJOdRnXfShudYgDkcTy8i69mVfmBJTTkYjcjW9tzyLidi+jgM8/W5wl2zXx
MVqCmlvdCwF+12fvOqdyHHnAF4lvOJmRbjZbIBqqb/ccHbGuUO8xAZtOwyJF
zTsi6ejVrT4tQDczPzMo6METOXeqCqzWEIdfX8CGdlowNx12B9iZuRd/o8rb
iI/E91olfgDjjNA0wVj1+TK906pw+oXf1zHjsNblbYb0R4M8Q7viFdgnLQo4
VKdqyxexj0KOtrmipnMgWrlodrR2RnkNIRn67ARlVg6OWq4KzcLUoptUnBY3
V58WM3DGpOjpyaGgIcfpoB2ZIh1fVu8jDy2crBtVi/k9yJ6BsIjn78kaPdF7
ERhORQuGChOWoFu8dad7rVw3kGGygDKbVu4aybHKt/34VapzmffT1r8Be6NR
jyKEtdKFg3xIgfjJZPpAwZEt1YE17R+hrTYUycVl9yWCxcIfyfdn6FCEUe++
S93UkX9x26M7AsVZUSfvHkTAOqZXMPzVjycbREgjRwjEk1Mo4AGCAckM1Xxr
uxHKBc00QS+908d5OSYi/jAHR2kraFw1qiI2jqD39soipUPWUtcT0UdXlz7E
FYD9GrmRLgvEfjkdb6WRcgiJmcscT3314fFq+8b7sgjNHLsOi3Wn1zkUbwVH
k7LOvDc4I79jwZZ8dJOXpYr0FZqf9qia31cgFu9S04JCmWyU18G2UkLdnwRb
AnyDHSCHsu3zSY8Jc/xe7NKTduaKadvNZmWBY7jjdWKALnNSCFwW1sWiWlbP
PM6x8G8RkhIj6bHVfKN6HU6WkebkvKm0wvjIS5hcvk3pTkSjBJ3Sz5QRLH2g
oR4TOd1hQ0ejPWwIWRgrCaIMRfWbv1q4feo5DgmZiGLmASZKSOoNXsJ38iFi
6ejmP4CyIcK0ouitptY8gP1vf0dH2U3oDDIWuea/onyE8uVRb2gQsWHDKjqW
FNrrb7i4iZyeSiEGrRY9rLaHqKn2HNfCV7bcOhzFw/Q7J2GD0I3msz+Q7w8P
RBZn1j3L+15z4Kv2ftxz3vvQSR2Hh2phYem943IOZ/r9tgm7D1dgaGA+fhbk
w9UFHj5mt8kHMAm8wi/KCwvBgTYtn4oPh5EHc0IN/92ug0shz0Tc9p53ltPL
ZVYKWd5WHPL0z8hAXNPehPrEKw8mWy1wPdlUEFPoIfr3X/YTMqYHow+TtoWx
nnwyTVQE92dVK/gg1F0CusUsHg8oGreCV0zbm6QFHT4gZTH2SWeC2N+EuXEl
8pkqrLRxz2kLJyNIW7c2Zbx6rVPsOtbh7/YMGZJhDPAt8PMDrRQsRfRaYG+W
5fkJe1Mgm6502vFpR7cf6gUdPE8VbUUF8YrHG4mI8GftBOm+nSzuDAcqznlJ
lQRw3vEaxvy3yoGJTJR85KhrnYhrGhOS9ErgC/Vk1jZga00Ztmy2ED5tGThy
c9eyguW9eY8u7wV+E4FSQe3UmlEFQF0omjFyBC36IOdJVrJUv9R33+iJN8CI
JKEa+euazfk0tqRjUyIxZ+f8PCXbxCP/AKJheR0sfmaiqGeaiI3hq6ABQdua
1d8cXmjhVoInp/btl8YlZ6WandgzXqTtJ6bnBMrrudgeeNCvCnaHSJ+O04xL
VO43V7TnhsbOTJKdaXg5ty6fDzorsqqQudizv8RNpmlER8CCdelCCs+s3pFo
IdCnb+tg9ahJujH0KoAxkQWG8fjaMpzU8VkwzA3ZajpHf4qPxtqlAnSa5QIC
FU6DDjuNwsUygRflFQg6GUs0lgUpfIlQfMXUoI+S4VgWCm6S3WYJCR0yXVc2
zJ+j3xEJl9Rhi+2ZrxIOdsOSJybbaVtcR9QA9OmR1wz9QBqyD83yRE646pow
s614wc/XrK4fHxOPl2nTRmDPkk9iqlubb0tvgv+pbkTTM+rnTGpnCTSbH/7S
QoIhe0Cq3wadriC2Uw0B5D4gxTzKbE9dTyCgkD1m7bKDXLlJRghlA+RyvQAv
+Ld9OJT0jE/UdsyFhOUmGfmRXcu2Mh8/0XTShXwFD/D7IJKBd4Wtzboc1Mik
O1SlFijPZil9EXYEK+zTG6Ck6o8WVEFy4zzYuV+H6DRszr6BW9LSZb2CNR67
AKDx0FSexVFaZF8OcrrOCaeyrEnAd/SD+zp4dNE4VJ1c2GiLTlAhPlw08FTo
bXNTd6PWh4VAkC2uGLrEWoAzqVsDxWHZu6EnXEZBkeWmVmIQPGGlIF6TLh8H
Ikrj8q4o/JZw2QgUqZbvwY0VQa9GzTyB7HrJB0OuZLr7rJm6Pyy3KFJedbkm
sZ4e5+YeMS7qfILfUgLTXZ6w5dxNV+3GL6xWe46XjC2YpTQtDRJOSU4XOUqo
XyQ/kLItUo8RSBX33YxDsYeypnfX/Bwx8kZus2MVYt4yyW4vYTFHFYUE5lnU
YO4pNdLwmgFJkor8G22MmWJ1j+HgSl1J5iI5vF8yp8qbPj8qB8i5/mFR+CJ8
odxyb86/SHb4lLweNaqrMceJ8weaC1/yJM7jHbOsJnR2N/ZiuK8al567B+i2
2E06CgYL1lyH8f0lcPe3TPSwSkOe+8g8s1qhejT67PqA6LTvsrjaK/WrYLvm
HQCFqo5pt4vC5rm5arQCnxQoem0b5c6fAGNZxwRm5DitXdEEjWG7PkPbyK9P
zcgUSXgQ9glOkjplYxCkflhkLHwn02NpdkVrMyyvb5xrAGUIz7VxzbHngi1O
/IpUjucNyUdczlhAL+VnmprhZHaVGwM7MO654EmeLzXFTaiy338aG4sOYyT/
N+jP84iXEBsBr4UUfeMm0hWfSWsYB0blbs7jV/ctT556DDUQoZSYypnxutf/
Biivl51oZ88voy0Lx8Gi8iMDj+TNS2/2QZCC3X3ofEwPaFTlfM3e/s14V62l
/sPNQxoxt5nuEabFw8+Y0pymrZmRN2HD6ho/a3A1K/6G2rM1ccHDICVvVbvP
V2nj9cclYScOwTjEfOQUxIvOWpCMsd8KL4IHVXxdHCBrSF+7WgE0WBbuhJfw
CW4FEO15HpZcItr8J3nzlUcRSOfJK+27y0URoo56QSKbiV4kygju9H9Q4av+
lh2akhI3CiyvpHkeSPY6duQJ5SB2/M3EVFJColxyss30qh07BMtUZRLk4A9H
0OkA4jdQrGKKpf0B4he+vNRXpJM3+WYuKj4AwrvPGkhoNNsd5S+KdHuFvUg5
cJsGPwbcF0FnaZ+S7Ba2GD18DPBXrdJegdeQO/Tk/nmIZKx5jw1dGOZwfzeo
cYJt/mpJ4RvMs/Tt9K1oiQzweBFXtQHDevQtP9rxTIuG4mi+FsdzGDqzNS+l
9r+zrChABeqOAO4TU6tl0cUVFcphv0JBxbTzcnaE1p2Hpmrs0QfreHsBMzMt
m5GYyse8d13kxiOv1RBfgwTFfslk1mlmCbL1EtPBAnBR9S17Fec+APUZcHCo
OkdZzg6lPe6NTXAkzy+tdjQBckv10gOeSSm06CVsNusjzFPKM7HZLLckqifk
yNKx+8JDEHz5vjcokqF0OhSTyW8S4MTJhlpLJTzxJWWE8GygQDneJDQsyAT4
Rkis5MHSeQEYBOqMWIhiNzg01U2yr1Eu5OKU8S45/36kMHBdw3VNYCYRkyba
cLZbIzXwrGWkFRvx/5jPzqsiV2wWv9ft9UIrGJfo8SRVBIOc/jvvxilZbAEl
D7UJsvsTjIWWObpI0lHBv4o+VyQAv/0w75ZxiYCHnC67S6vyaJPtoZNNOWIh
l6XlnKPBsOAkA6aurrFfEzkJmUJoUKo442zddd/lqZoMf3jR04ypMg8b7D7q
ZMJCJvPGiFXpFbIxU69n+rgayKpBl8y8zID8TlwTu2PcUvn1HcS2FJTD7xfy
jnwa7K88fWVmuCpsXs5cQIyvnXUFzeQY235X+mWROWduzMCowOJ1xdahuXmm
ZsT0F3xt9SMuNjRRWvBrVjRvz+GltVbjM0PypP42w0l3nlrJM8HM7UU/lGkb
rAnAsxL05OgQbyDRZy6o2qE8qzYtlwuttaNfp5ril7c/Tysi9hx+/VrZLc1S
2HcamUnOE+YwkCXWY5V4ee7S91sF6qgdbzAJ3u7MioDqu3/Ys1h/FNJZcuYI
doe/hs7WPlE1TbohmTYAn3SsJKswHIO95WwVrhIz+cbecwCrubK0UU0Y0Gi+
7U+EkzVIOl1urBMiQ+yIAskknrM4dCG2CAGlrYWkgola9bt96nib08mEx400
mxsLx30A5vXEyU0WFAc8z11IrZZkPqRRy33h9Qr6+0dZzn+mDmnYtoLvUQL2
uzpA525Nfci3mn+1ylOihLzKbY0gvYKuSmB93ZGVcqJbvcp8AaCMG1z+9w+0
1dmN1/M2hu0V9WFOuZvs78X75jDaZOuJh3CFdUduSw7J10+Va1hb2DaAgyH1
gYwvWAy4tq1UN7GxHRUueZwNnORXNcrHurBwOgNiYSALAZHDtByZXjMKAuZF
MlTT/3U7xuVO33dxSrxsTXN/PFba65G/mBK2ndzGzOy6+/DO2k/HtL52b+k6
xe+FmvmhOrBo0SgrD16IQz1Bu1ybJTiXtMJzG42ficG4Qk0f7pifsnyuMQGV
mrpA8qIrYe0YFFd5r+4dJZvBy3mvqM1fAevotKW0yQ94TXqcMeKQDwiMZPAF
9w3FhTdCYAErWOQbrVKvkG+l2DWizGN20YrAdbDDdgmzmkdJphQjtKvNQFbr
zE9cPQNI17o1e673m/YVqHA8pYLonn5pvTRFelELnqqDoY4fjDPZ6KnRpLZ9
/+1r2VrMVPSXfd33KSh6hrDbT6p4YzTY4oUKdXHZ9v2IIsKK7LvW5i+04n84
Y2EI707O8jv+tScOMZkxDYi9eWbGdhN3UtUY5NIO8izPpqnXQ3iyjnaEhhTQ
VrHrERmkC7w3RlS7rzqYpJ2uywK+YJU4mRUG0kmRs4syzpaNFXNSu/ZozXOt
+bOl5+xs/nsiBQ+wlf3aZbiyKdIEavG8GPdwI9laI6Yp5y+EoCXGYsNSJhe6
earMzG0SklW0XtBVavB52lEfk/0aegoQwDZxfqajEufu88BvN0eWj04CLx11
pUWQdkWyaZ0A9Gmi1b6HxO5yVtdwUw0A0J2msAgH4ZP3+r1QIxlhj8fHX7W2
lquozG+/pM1upsw/wXP+XXd4Uxb4rw/+SUD1TLTIgumhAJDPGvxhnOCjWhjP
sG/1F8xZWFq4yO4hXsrDSBzxZvZn9GmO4W/JJXoQhWniWkTwVUZIIw3xCCQx
OSF/LEB9ovDiFAND1fUNnTaphaj8ZviOPTQU7Kj+Er0w2PMDO8GfgcHv/Lc8
Hkjf++BNR3PP3tKZEc4xel0v9EFlT0PEA8sKgSj042W1cbcLsjdbgKNfchmL
rYlDdKNvAGAAxRYp8McKvyugVvm6MU5fLu1ojui3/aLA9lT8WjZKkJ2/bs7f
s98+DvfcjI9dzuMZWpN5U3UPZeU15yWVs6InaDUoPpMJxL3LXNS1BLIJBjUi
StVFlFp1SMe9Q6et6miCfCOt7D9VTMJlexVojvhgzzfH6sVXKGCkfuXNr9kw
cT+gyNby1QKU0Iq1Rs6RRBSXIsrErUkWDkPdoWUxQixwjdUF5tiKSiZI6nga
ZmFMe7aQ2bB+MSokDPUbp4fB/ROCpsGxoyKQBi2L7eijUXVdzJSdp/EjCqNA
xNJeRXrT6/3mAkDIrVqt2P/JWVOrSXRsUCmbQ0FKhGug14f1ZRxplmLdN3Y3
qSUAup7GFf3dcOS7rV0ZAk0LMePZ5CC7IGSs7rezquuvvAGesEybD7InEZHS
q+JQgmtVg3jvwMWeUaFFhT3HT8jlNg5r/MHuCzlKLhBtzLkm/S442jDrAhRN
W1zsUC175Zrwgsl1SyGIMsjc+7baaaOsqGjdbed4KNDzL+aUI5mxSo8UQUeI
8TonVhVm2L1iOGZCudhgzsft9h3pc8PGRS4hH9ovl6601aJl3p0IwYXJQboQ
tB6xLuLJSEXrC8heXFkMtM8yf1HMZ7B6zM2xgPNFSQJHt8wiYr0l+iAfdRIS
y6NSfuJY4/fa+2LM8tNG5TdB98rDkLB8NjQzptk0QBMiuxweReDhD0ZYjGhw
4HswnHKELUHdEgH7sbZLaRig8vvVcyJdJs9glbmtORVzKT+qmjcUzo3Y7Agb
YoDRPcRUocysXZUq4DtbsawSIGUX9otWzueN811EUXAtwDzI9kgcGwAxEcQl
KjxUhe14rH3wksXoBgJxwH6y7mOSVErzQRFmfzG7mpuVXMk/VYE=

`pragma protect end_protected
