// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
JzRPNZAngbUS3tHUwh0qM3I9GYlaxoWtCqfGhWSJhSXMCCaq+Bs1bBBVWTcZaLTB
Ln2p1rsYI4k1UefSZcR1nRLC6bN7LB1432VjsQFcFB+ocioO9HBB9mGPljWGFdQN
vx9NkeLG6tx3oq8w0HCpFswGxnpd6LmjE5uWWRjzKFOPeVrqtK6DdQ==
//pragma protect end_key_block
//pragma protect digest_block
HWyMVGIUSa/yJjnSWOqKfqXSn/A=
//pragma protect end_digest_block
//pragma protect data_block
595naomsH1M9dXCeTaFeghgu4fLdZ4flPF5CN3j+pkupVpWVhQwF+oRRP9PdqLXO
yc+Wcxz1zvk+nTkDHjW4LOvfAphRsmnOw7YMiuRGmwD/SX5G1eQsdlibjQmOUhEM
zT25m4aGROeEJT+n45sEOEGGJEq7ooYtxH9B5oQe/LLyOqUW8QgnD8Lf+SiBIUc5
fhmrPX/x2XaOrzOqJ+ESU7sMcuyse9CW/rHPWfeLlFlXEnH7E12IWcN9Rndm9/9v
5z4ZacwYxdb9vhsTQOyZht76yWcm7TZzVZB6nMxsLEKYPCchfgy0Ef4DfE70OrJy
9shbRhEdHiUK9GDJak2Skm8Y933mTOnOwc6QKvd/1WO942RjKqK4ujAY8LAl/FD2
A5gZwx9MJ0Am3moigYKm7JWpl3+5apsZCmqYBmdIbEc0Nxb2+OYjQVlYHVdnridO
+3x+kNWsCloD2K7D7i4bVV6/2kN1EpeDMVaqH2BrkUcQKIdu0wWH4LyEej068Yxw
74kFt/zThtKjQbv9afshtWit2Fc17p9Qge5Tq41kXkdvhJbXf8v6GDSKyLc84s9c
Se6IimwkRUmRVaVvGlY3w7eIqDEbLv+bxt9BzYWzkq58EMI3jFnIm4Wm9DMDFhCI
yQZuUorL2cgn6THSyTbRWZsLPckiVYx4B6xz/qO8XPIm+XZytl+7UeKOqy9wmZI4
2t854kTKQNGjguwi3kWIVSBA5Qobz4+OhXyC3+FdXWKhy76ZDqvzD/rPRcuNbKsx
x/3IGpz0YDHgHNV1BE7YZazeiiQpE5f/td9+ZRYSDM7QNHVT752M0fm1PqiuSr0L
gas9C0lq7t3UpVJ21iO8Sp3S5sNsXyvirghd13JY6NwcxZnTN7xssp5mSGUP69kN
uzA372SzzFfFkrU3xvT2II7D1+e1KSMovlwSXdDOYC+zBt/2HSvJc2KgsY/HkihO
TsoY8phpHWRwoYRyX4eyddzK8stjm00vwa+D69H1RMAE9/NbW06fAURs2pQg2eAg
jFvHaahBHlMSz9rCkWTgTZ4zE7kxnVhKziHw599vVVcxxu6TmoRIzEfJuhX7/jcn
lRYhnV4oBKP/LTy/oSg395qI3v36pwqxBVndmIXySAlFRwMqzq9yEeF6ArfQEQ4A
PuvUSL0zr599wuR2XrSsEplDLpxGbBSRxbn8MbKsbjqTLbPEn8hBSijfHXUUYgcM
G3c3qaRMVFssrh2cKyywOW9DYsaFp0vKqC83cYy/6I8WjvTrbJNf90fvLD1oNMce
lV6LK33NOk9Zsw3VvKtOlAqj42iu3g6MvZCYpLsAIhbPdujvLtWc3iOz8NUeFFe4
v/OkeTHlG3zr5TT2314Gg43ciOQ84Okwc0XJNn8jisGn5sZh8qveufNi+tEIMxq0
wdPPEMw4+1ii4zYN/nYjZCGm5f8TMGHSlFM55BHJTpnHxu6YnvPcjWkflPe0W6sY
QN0KcnLcp9kDNxCoDiTTgTrUKyDVVshahp1HjyqiwT42ytuEKe/yaxmzQpytTTh0
ZhU0wQnLC+7vk56WON1ga4sHfAW8dluSDW1P3v6YEZZDkg2zwUwUGHBOPCYdXS+P
vY8xAzuyN43CKgHgwyv9FY5iuCdQuOwFFLKqhMPFKy6bms49M5ToZLpMrCc/yLcN
JkOS2T1R8PyQU3EIZWAB4EFMnGf88Uu1fz4xBa3R+vcbuLHTyZmuPHrfmBtauDwu
OBnZWzYDKMZLxYTGi35td+vq+g2lVggmkXGQxi+Qk82Sx2ZRx8GgTIAF82f78yxQ
xpZN6KGxw+Sj2tTQS6Jh24WM2DlYm/dy5yNsVB2ly2/Sf7qbEj5XNS0Z2cUyAP78
LIHSlnUh7LYaJJhuCHiP+PgExDtz0xpMwfLfxemnMsrrX9vTyBAcY3X+5mQKIFiV
ueWcq9OcozhMxoXhuQcQYnYIri5YX+CndffdhBzoO7p0YkssudJR//QeoiEvnTkk
VDeqDd+0YtCw7vYM2I3VzKlr8JnI45q5QQj6ckUTbf+ja49pbhgL29dgprAVr7Md
WCo9trygnp1HgPL96E88HRgFqbGtkezsKWCmB1pqGaO91jTJDyMzm96bGoBPYXt/
EqnISqatTsTRh5khG7uvYPdTohT3+MJPLmpbu3qWdF5uUtm1nnwsEVtfTlM6fFGS
Su3afbILc6jwKcp5AnLMT2AyktxXP5tMCs2TU55LMjBeIf/VFeha5+fmjF19AT/K
K22re1KDbPxt8dOH8MDO06z1pgYOqMVYdacsPPUAvgmmVp3GSckv7pHGFtiDYVDh
98hHrAdhxpebaHEgxmemINVDg+n/grdk0OzQOutaQfHN1bEgZCgoqTHw97geIR1B
NGOqxqFemCnIclVaWzNTqzF/Nf4R7u4DN7aV6j+blvlmC+orOIHfatP+aPYDsg3C
K+u74eYRtZU1rKCWYc/aAcQvMPuvcobhs+jpm4lU3dgo6TFCsr1pIiC4T50esX9z
1ppnR8GUaIaCqOz5Atghn9ycDmYaI4iK90Zk8iprtX7ruwo0/kGXGRf4zH9fSkZu
7tZMtjiSOSU4y9lkOKeHEXUwfjjSAufXfNRDwzPfx3mMZtINGKk464wSJtcprgYQ
ip7MLfCmSwb6h8zx8c+e1jvaobjD2ab3YDpzptYVZO98AvVXUH1ssRCSVG3SkCAt
wIV0uG82bndqMZSLF6DO7jG63AIAAf8wNWQ9Z2USBEQt6noP+TkOJIslO8YiLtUZ
fMPwasTA3j85FM6BoBPjByFONNNFXjra9uw112VbUGyi5NpxTXTK2VpmrVr2qjce
Cz59KljwBbZoj7A1+AGmKCfV7iRCt1Flr/xgSHpOyqAm3xAyWt/5kf7ziP/yW86z
WqJUe0NYyZjkZ08YfiCC1LUWoPyJUnzAEsgxgkFm8vBnfhGKoEajWcBS7jdSN408
4P2ny7JOnNdqQB5hBvVvjBh4np+bKGvI21HA+15m4SvUcOG2r6FNfvUlsao8zztW
pWJmweUET79VhZapz/U62/pvj5Vv5iM/wOc7pQ0Jx77cAwQVTrF4HD72s4nAs7rd
zahMjmqeVUxvtWtZ0jiHmST0dZdxr/RYSIjdOVSKzST6IlQlejU6HhZbiSY6pMEZ
obh5xdvxnHb58QSVCYg4UPt9vZoRKax2UAFoQKF3h5M5mKw5lLmpTZkz9LrTmbQ2
ab0g27ceJqgwdSkdjfZXK0EfuY9EMNHZr5LGH0d3LfqJa6FZ+xny6f5EKuH25CNL
+EmtmKW05Od9bdFyrNWaikA7UH8OzIl4iaHmPwQM1d0fspOP5T2yI1yGc9qupn5i
UiLqgNFpU05GPcig2xylfPUL2m7ZeGe1tsT+A69Hi/KjLqN2xtUtvE31TRETRxMR
cyluddedUtdd3pzK3qaA3aYueCfwjvbBNofmnhssTEGFtXOre5AprbYaYeAO1TEm
3WQCXZjEsLBe8cLFC8nyTzt+hDOIudN02sPLW1GMy+1VboMLNV4XgyOeteOBu/uU
1dxEF0rDPxub8FcukxNq7FSQ9i2wj7rwGJAzrqQy7so63WsVIi+BTXLWEP49vY1K
0/OfToR+2tIKww5odrkAtQgDraJDP5tihugiuOsLHi/ESpn1+tlpWA5Odue8Iikm
ncGcz+EnyIkqathFTW8EVedXWwzQ71TvXIvgI85gAX+u9allONiSw81XHN8883d/
7JIoCvhqyq9KKtXn60PePmkJlpr6THS16Jjs3A8t7B+9rNakJXv41oZPlzaPsW+v
a07nIzRq6Myb2bnBziAG8/8KDfEr0bisi93U7pb9zt38WrdeuNQAY5z0Fm9HTyME
cJo7nWXoHiSHXaV0IyA+2zhaX/Ccqwy8gqeLZIiACWBWm8/LYRWHXkFG+EBxBATr
Wbt41KyxPaooBxnn9uhwuvsVrbd9BFzTAFbQn29wz6eCb3iCOuweu0rnq1fuUYjk
YKoQpcniXfkRzLLk2DVGBp9y9K2+kp8eW9BsWFxsmKJYRSNki8wQTCyBfnp8LM1t
MsGBzWOK+nVsMa+kMRy0cyvnNBbRsWH2Ocf6CZiEj7EHwVdbshMjZmWsbnLGCG73
GiewQR1qIOUE2NqJL7iVGutuZAzaumnn2ldmumazeZZVnOtVWuiyp0UrOqMp4MrT
OQa3cR56p48F0oHP94bLfsL8fmnfbs7C/QwNFx3HLIDjdkVMb9Ezom1A0mCzrW4t
PIrXsGgcixIrJ1GAlrYX0PGMtOOmZbAT5qhlb2lAJOqzBDV4SAR7mX9J5zB8U5oh
+XFZ1Z2wx96zWqwl+XvfBJjsVnUhJxhMH6L9vCJ7oGHdXMq+0EWYNHiqsddfa4gx
BCIGIDS0H8Q75R25uba8fCgOQwzworr8JgogkcTK/jldpj2HLoh7wRBPrXD1ZkeR
02wJpNUU8ywyIRtxKaZHQ0Wv4sCxFaG2nWpeHWSDsPH9k06C+siVMivnClndlMEu
F8gWa6ehE2qxXK2TLvMbWGoZuYLqrVvJficW3d0lrPtPj7y5CK/YHCXc71HxYjDv
pVBmTOZpe7B6tI2ht3bFdkfkI8bX030z4nTmSIEbHTI8QEmD9bbu7Dj/V7Shbdsk
fuRQsEel6Z630jsOI+l/zNhjMFM5AZAc2/o6ZaV11qHvFmrVkJJDqYri8cmvb5Bd
Rh37LC77uSpfBbRoPkAYnzRhaqzu4qck9/t4OlyGzlVwL8VCjUbIq/5AIxTxon+g
CvQfGq3+wJHQoBzcXj/QRiButqfidTEV0BlnqQrX1uXGjur1ywvU68j/5UdyapkT
x0Ytu+XPyd37kR8DBZZ8O117Xqd4uIS3f2J3zfsa7hNj6AZ1BwQTkWqb8RcjBV9K
1LdCsfU6/xC1nxHd669MRLUYCSY8hcxE0/dvudFKZ8eirlmYwq0PLUfWUygmvel/
WEh5S9ZAANiu9RW4u/bNNfDq1MAWLswg5wV8f8gJjuH5Dj4W9nHE27QqF7M7dT7z
4mYQOL698ehJRlnOeM6uK1hyTY9o8HUYbvDSyYA/E/eZBdlW6dsuBdafMfmREkAs
PsZk8wXi7YcYQskHis5e/i4nREDOXxX4QtM4VDoUJkBKGYn7C9LzAkMYLOkTiz5m
WSZYSmyK0++BxyopA8k48nJifEGMT4DoUWSGJ0w35IvKer//mqFoHA0pbEZHA/cs
tfkDtq0RVGX7A6R9MSkszc0xA/ZjCAIYAon6RLOv1AvwTOY4QG8enAA1D0rWCHDr
mMcsGaxxyrcPLdch0T9y7heKbTYCEX2QbOlRNXOZ0+6EyFrGtCFFpU+JcuZ3alrE
aWD4IgP8JLRVAb84ngvoueOaiqQzCpzSdkMjPj7ugAetWDYzOjS5fyz5yLrzvpYW
QA1f4Y/6d3bfKWsKwMJpwMh2KXm90zhUVCBdkftf1MwBGUhDZQ4+9npXkYRbrHXD
hnioACYhq5+gdSXXddu3wKgjwHQlSiJLItp98KLqhkehdjx/hLbdchVdgt0SWzzN
ShSUZjFYr8LS8rZNHTsB7BHe1ANwbvX2/hB+5sc6IDUxCEbipEfIy3YJgOBlbd3d
ABbfxH+Cd0x8Z4BLV1cntQON0ov7iH8XiOYyXNwL0f92IKa4bx6DGnLdVNSYX4Hu
ZGqsR7xeYi9+0FYywb8f32GiD6tYMMUmH+R+qiRDoxmVVQNZPx6VJsCB3BODiCnv
gTMtTqGHAl0VJHzrfS7da9ML+0f5udd8A/UYP1lmGUdgLY/h7MrcxCo0w/jlTTG3
uk+KJjyQAER/2znCycCR5yJ9RuwDFn8d4e+b6zLangoWS3Jnp7NYLawh92FBPiAf
Fes9rukI0KWV8U/GGykPl4rutNZ0pJzAN7e2IGnFjCiaZlTx8PuHNqB2WiToK5qe
0VnZ7UjRHrJNqr1Zn6HQ1LuI8uPm5iwtGXTNWcXzpcwxE/pUt3d31PSmvQPAmrRi
bBoOiGXP0edXikqfYeT42x866C37fl/xsJG6ynye326xgvss8niUXHpJhW/TVQhh
/rWn3QtCypwAdESnk1NrVwP0sA1mg2y/M3tU2wgZotqVePEPkVaeDMIutGZgG5aR
FGTR6wUQ5c5rFwqvT68OZCMoh32Z+4VdDDbnVNyeaKpsJYeIBxIJck7PHpNqxbIu
PDsTWGNmL8y5T/fCiQ3Zucmghi+QNbLFmRigvtFp/mjRkmS4FXHRVxWIrqJFXWvS
zK7chnkeec55SjGBUtzzmqHLEnrmQuOxW68ecmg2NIInoiQGLxDBrpxx60K1cp0K
Bj+RyVGVEjWsityojunyDwEDAyshaM0rAicn2XLvcvLWTojV0JTB5yJXBuhB1eaJ
m1pde80nmNtpSEKQ62nIL3c3exwlrAszoVPBmRHt18HtOsMFyPptQwe8wjoV5N6o
b10g/J+IGDYZ30AGDLkas3j0FnWeuRMKT2h8az56ru/RqLhOOb6er311ivCPGjE/
xxUS0EbFfpLImYznpjAGdju+sNESX0n1ZcxfY9Nhn2od+LtG7ZvoOuQwnIh0EkF4
sL/VRjMT3AV5ZaUyCgZ6IWPcyhBHR9tYuG5k6tS5sB3xtrJI74pHlAEvCOLui0QJ
Q/qIHEr5Nr2iBq23rOutZebxMexsU3mc2SXuMHYRsWDZg79Ety9UgVyAb/oTT5sL
FHJohuFUaqfBlhlrkrkDO23kpbEF3JuEAD+ZbxGFpZcgcvtm2IodVcrhWSXFlavS
cB2zp9bLbGf2vcxxNwH4q6Sh+IEdnBzNS6KeYCXBryWh/S/24JMf47glSg6jRLsr
0OtpMbc0/sCRFJUaqM9UORNjj0+Ggqq3UAB59Yfl6A8zT6nUFOpbXPtwOx6kKbqK
G3pQIvGPRKFP4oFT2ZhCDZHu3api0kjwF7vU89I/mv0Xuns1RWF2p6ZLtBDwZpvY
/wKFilLTiw3HQnq8oSV8uWheWZX/hMs/91iRRJ5PzYU2eEsGfuK9ZTKMpRY4Le03
0XixqNSi86+1D1SnmdYDYivsDqbi56rTAb9E6+lDD8Iou5xwcNM6/cpY30iSbcZQ
H3oBD0P+aUJWLWGEV+B41a+fwVcL2eQoAGt153QKyOWSiZbOiHxRAFnzhyWU5bvE
JM+vSvPg/1QGalNR4ozPEelq4S199vh+OjcPi4ZPN1RI8Zaw+R2SnHFPkaYmdNCO
KDlW7CRnPspEhTYnZ69HauhbIF1dJQWmt4w5qcBzQfIW1eK/6Q0qyzwO/QUCGcnf
WF4TMwtl4DwKxYLFn23nsxMcWEatDxkir3ZZxflYJkDVBUu3pmK3jDmJMjTNlpV8
+8u5vA/dT9GNxXo4BLstQ5M4gWyJN93imEYHeMPf9KhknbJ9OcUTW4AXTA2G82W7
rc4QJKZ60T7XztQyin3WSRDLOjbDARRmdjK6CrfQ9mUht+C91x7Cr+wBUukZoNbd
ra/Y9BNTjaVc+ALvZf/f6qdzctO4ef0wJCZ2Xf5K0T4DclaU7TsTbRliMgeumWkI
X6HayPpJ/BHQ2AKmkwUlyO672FiSKq6MGVmJiNQXunB7o5L4XfyhryCjp/ApQMyN
oGXRwECJECJqVfLTORI/9nEslnzMRerymieiyq6BqLsUDLpGeym1CvcKrDnl49eg
qj21+/kDkoTkwXM807vag3ipy+wgkmyKwCXhqTy66VHhjmhByoVMLZmPWMd46niL
vlUSifUdSGK7sThkuw4z+qj9o6ad4lGZnaye0nW0xrRJvQ3E4TEDyv2vXtAblTA6
JR854tv0OEXT1DyCPXNS86KKKHwAoKGBmyNfhkkwQcx9VK5x0iFWIIrQV8oO4nSO
2S1gKC51hkARN0aq+DldV+5Mp9J4/ckgpH6Tz7/y/Tz9Vy7/acPMyQur5DhXSRGl
INcHFWVeoc5ZbTBVe43z3jaSlznuwLOMjKX81uVEGRWhE8aIAIu0r/3P3zKE6RVz
DQ8PSI4Syu4iTF3ovwhCw1vBmJbM6SIY019fo/PawxSXFx6TLGpw5II22sXIlscC
zd84KBhqM0zhU/P7tVutA05D/8yCRxfV/XGc/5loDyN/10Ac7BGdPavlIc5CIm12
fmIeati5Zq3JrP4lWsAu3lBnN7sLPEOn4eBeGq520leduvcjMH+z1KUNlDD66OvY
S4PBzvlyUfgYlmhRDNvg1gwJo5JnmMcK50yPDCdBZ6u3c/lDK9RIL+rOx1LJ++CM
orHv+CCV1Js+fmlewfBNxSz9D+u78BoyPO7+IePLmesf+IRaFIpREouTnqAEOAmp
jlRo9wEqOD+WCc4/caikwALoi3xYbr0kPyj4pTxEl9r/uGw3kkUed2E51jPIxAl7
AShH1UIW9VZS2Yc0x3Moi1nOFrTV76sWyn6ZJoxMfOkdATYuHGU0jvuFbOUFEvdK
5AqGIOh0gQ7MVq5auO3ZSaO9XOwCFFKFysBHnTefAOfWiZYJ9uQ/72sfyk2uR8wU
HYmBbk+Jpi68QRQCjDZ2GWZ8A5Lspuxja5Aq5+/lXYr6O0VP2nzAFi4ArmtlbNTs
7bsyZlcaDtjdE6pttVresThlGZPSyIXMMsmoAyhMbSPomST4msyY7fDhnBYZBFEv
cC+tNckfUrHs5LCvo0A3GuJaCubP5+uZi89ZcadCNQJCqw01r2ZdXFyKuEufMc+B
XolzBmz+J+AnS6qqpq2ql6kD4oHYhGfjvPpigKznD02woQjL8qVkrL+CNj0WiBKT
P9B1mJ1kOXGFTrX4ebE26rkwxR5rRr/k9HlpI5C9uYDBceGI+ZKv0x6Pd587CqXX
fYx/tuJCSWy/gAZquFcpq6xIjSeJgKz98rAafC4yN2C/X4MFAq15k3iwYk2423cC
91G228L3JU6O0YXjsbc/29oD2d+5gphD5YS7lKX0Ip9cHfVLqATdk20FnoSFsug/
4C8HU1ZQSNlGvpyD0wEBB3OehHPBh7cIArQzdFj4Gx3ZZq/KeKTrvn0Y0UU1z38r
EHV2IxyerkAebt77ocW31oPY2tLN2o/Qjs+Gg2146B0M8WGX0JL/bbE2WwfSjXDA
XB15VITl0iT5iExxMirlnWXTKGGhMLJQqvcc64l0lmXgzrsx/cZyx1plMe9eOov2
jOKAJETw+sgrCZUvANiVPrQYILFyO5a+1QzBUD4kNkejBw0/B9jDu3JhyHby20zy
SsmsXiMUTRGKdKuu5ejTdEhS+bbm4raij8kslu0y2h28jQYXBcNYwZMglGx6T5Qn
qkey3xPucrlGJhu4/3FY74Y6Bs30y/Cf8DAYnws/bJ4FVJbdUZRKyerTCvMCkvpa
3suyLwb6qh4HNwaiicmzs3Rz9jTWY1SW69HgSf1AGvXRE2t/E/mhK5KrE03BQbU5
300mHNdmRZTNOPvxoqvO+Of/ZeGZCvbmedn8j2vfVr18gEBCfjwJqWV60mPnCYBC
ybaDgacj9Ha+htoJwOrw8Zf/e58G84TmDfTLM/dLj80W4a/nOA1R+pmhc6mfYXOD
1Ga13KBrX75xiw6NjA9wsHsYUB1xFWFhX7as32Nn7u5wTwyZzoSS4QXblUUJl9Fs
VixCEcZgPABd/OwCxYHY79BRxZUB5UCvYefSmQa/BRJ+vNcK8nP1v6Eykhl2hmaG
Kv7e0w4VJ5sNgfu1ebFWMTdxoiF6rELOuHrngO7mr4qGeYhIXjUxFysUyu0mFQCR
a7Au1gW/ISwFD9xAvX8xtIMe/q8J08DxMMzr3PszD3nHABZaJ6tAhr8NxGOF9lIz
trCa1C9V0Ogx6Rf4ZlBsfQ1RimqfKepv3nSqajb6b+QQQ0r2tWxKrZe+9RvhOSE0
jpeEm/uzjdCI5SFE0DCJjC0mOGX+b1uelp4petp3H5y63G1n/zo/AbtAg2bAODs2
LPKWTLhQFWDsUjC/L03cDj3J2rixZXfbc36A1OsN6MiVNsk3glHNQlqUBFUS/MuH
yqjey0rgMc8CoqGTCswgKL9Ot1KesGWH4nXUzaM9anIDrkAKXdoI0Dy5/AYqi4fj
j4diAIKjwIcAfmRjyA0ipvBh2ysguTAfa88VLh/ccm3X6fYlw42d1PDsg4e8K9AL
Mo3DPObNTPtC2aTXe4+XfVOJFTqfV7OdwTErVBLrB0n7jD+Nfe/tyMINoIYc3/pk
l3YiukJUcMv9qQGGDD470HJ5zn80nzYAOlxsU1PA3ZuWCvQGTRWVjBGkygFMyW9b
BLpfj0HtqIpwX3vYyf++2CFWYuH9UkxHR0ll6IGweNKyHngfJwJwgJ7hp8xCuui3
Hmc1zjbSOLIcBN2ooNWSU+qMjr27klnEyJJt93C1VBlD9HMzzAUhZDqpZp/DIYLT
vxv6+A+cCJkC6Udx0mreIsB6ZQhMjrdBkPLJ2PTxBAh+Zv86Mtqe/W6qj5mfG2mF
D52/AnnWlMqLRKuNMtuoXPF+WqhZhpzpwR0EFY+vTHxH2uvWv/sjscsV26wKkiFD
AZEYRw0JgwVBDDeE4n75apcg24HegsPH8kfV91L2bQh+AqG5R1x8tgFJbwxNKnjE
5PwondJM1y9MbwKSF42MO7rtBCK+IjW3iwch1LK6JUPoRRvX0NZE08Oy+LgnZFir
FFt2gLo58UPKYp5hitQuXe/TBCNBQV3T9JE7uedCz2mHIuTsbT2Q3yaxN3oFXYet
ORpU5qnEGh3GMCMNPviACfXuumH/kbRkLy502+Zf83U/s0Cqdj3C12WDaiKLfN/F
YljOfbjEowIgcST8TaGBiv4ZQHvRxwq54OzXN9CPPEBn3WMFQhOUEk+iNE0o3TA2
xhhPeaP3+THqHyeMzv+hQJ9gdsnJVviDNBr6whhkO4tve/oFvZATBohy4ZtoY8XU
hIBGzSlzxfPGCh4dXXTY52wiobbe3J3+zZYc6EXUbrTciEVnj96h+uIsqL/xoR/e
O+vwNNTARvJmgQFl6qajKsRMn0NIPm7pbv/hLfUKcjozcTy+yZgE3Mi1iq1pmIhF
xGfrCvNPZQ9wiFKLteBlpUUJyhCGmLUftMxQsCjTPALFOb1T9fNKXNatqJ3Dvnxx
GWHGyOs7T76lYPSmgk3lGjhEAS0dEDlUcm4sVBzKfzTAQYCujf1LFcxuY9sqU6i4
B2E71N/Y3wTVupBZEMz15J4rbG61p708zwVogCucRsCQyvGNH6EoGLyYhL4WTSk9
ueK2RCaoHvPbxknH8/HLUFV1J7YGbmdb2kumt4EwtHVNeeLUn9BuHHQo8WFWRUFX
z1l6TZIHEtCqX9ajAA1Opb+kV/LhWWc5DaqSD7nzhwuBaxQUbvZtC3lpuv6Cz8si
P2VfumRWl9taz9ax43wubb17Br3KQeWCRbSOvkeyXKWXsJdWXuxyXDf7X3orFD7P
dRBWcsvVM5aZcJXA7oEoAx0iF5Wwod8CveUNzFPqZICuXb1wRul7wpx6TKQSPXfV
G+fQBca6pBziXPbth6FdiK3nwTKX7ggDfZxVVNy1gG8VY58nGhvA7cyBAauWoA87
N2MwuriNgBtXGOpx+xNp/ppWR9JD1WaqLTsPNqLDdK5A02SfFU9NSg3udRB4pfDB
WMQnWVgwcV+c/Jl9wjJzEba1iw1RNeN7KOrlkc9qLPWPFCy2N8746ebMXFfOccHM
5JfefPL8Iejfdfn9FXU3VQ7p3B2zZikCFo1w00KyjJ8GcXjWLitQPmPb+7MLPkKb
t16ZhAD7tK+8VXYv4F931WF8c8kHaA8wBdI5bdMrYnztXg7gNH3RkZtSYKUvhmN0
0feTlVzIymMVdFfOUkBAHzm7RYA1HHyQOTVqslCIDdzPHZ+i0fot7TmCYlatgYal
c5vlp8EV9XUL4ltnqNpzk7lw728nEIKC9AdA+LlR8766DnQd4NIB4Nt8K+nkFSMs
8NmX6rgsBfd1nvlpdA8uyJ/jwfZfrb+mQ5nHf7WVuygkrxbgUzZ7JeJFGw1DcYai
zPdUGJgc17SFpd6QkkVtiXY4YvvvACOFhq8Wzhf/UCXW7FrJwRs4DiIDryL2FP0t
eP8wK0oVRwzbQ4XKo2VsthjOkOyrfZIPl0V4uyLLgSeBbND3pYeahubpMNfTPVFe
GXia5WBbnpPB90k9QFDwvBNnyEUVCGQg7HCeHllmbDMSgtP3sTXR/XqhZroK6QI9
30B5FDfkWtIL4/BVmDNtxzVIp3KJDbiJaoryPo2khExiYNSfEFcrvItdJ4YpmFkg
7xWT7/7b+Iw/7les2JWdiMzUWLA2C5KPrks4BSCFdzCVv+42jiIUryS+Bnk8EcvM
vhXTX/TqKH+zD491VtPbiDUm2+yByZ7K8HQfLRaKDMkH45TVOtwMvQF8OKcFa/se
BB2IjT86nHHhKg4mxe52iUxcucVTLb9k5tiZraNC7jy+zbqlyHiC8bt747pd5CER
p3M/88cE4GaoFGVtbVbGZdZM9jsJJR6QdXQVTVxLwBapFAvhxwnsVVFe6uS4M3a6
ZAvx+u/7ofE6+Q+sZ3Ax7s4L98STe5m3+rq0NM2Xn/Kf+71kL0KE6pa4po96FdlL
eoaKIzuynwEdXsuZm9JY3AMtHgAD6IXNjCtVdg9RzbDauwmP5rEuF4xPxPL+EL+u
xR/oTYz0UFmxQtUcmJ2fPehkHLQjMB4elKX5qGVteokE9Bajcg0evlW53lpN8Cmq
JUGAOVG+wwPy03hNkrbd+XFImOWZE83fl+B80SFPA0u2toyKeTHHPPv4BuTUZMzw
gzDtjlv5oSgG/sO2MuPZM3B5cnRcqpE8CaPenDOo8VrfaoQswWK0ImIz1vMzAHVr
/ZCO12/Klqy+Va35yTNqlXnuwE+LCUCVr2hCcjsbWDCCVLFNw7tHhQoqa1UCQRvE
criqwtJu8mQ1eIYfT3Ge1Mesi3q9BYF8V1nbAv30kNqk34T9efPiz7HYS08Xu0f1
w/LkbaccurAXprDSVPY3/X7YCVePsf0GmqvDbV3VTosbqS/VYA4ODSXvMYmzkWFO
XDVvd7Bju6eeFDDJsOipVzdPvQ4TZg0s8q/f/Kgtwlw0RqCch2r1WL5P8vE9GHA5
ccJ1MBnEE4T94k9P8oSvKGp4PLWdL4nvLxalB7RPg8mVEzFGcsPfo8tEQAVHT2Zk
yB53JAKdnMtlYfGRRO7s2th8MesCK12lwqwp2SrPTC639h/0w7z0klEnIRNnoP/V
ww8Nj4TFn+JIXhnnx+EyYnktCNbrj7OqAlWaqXAI83r6KHHLhngjRb1JX3JkxDus
rrQ0yiFLZTtwRapUxTdrHMsq3y465XOjKU9Y1DVEP0JbKdXArpsNjirF10PCBmyi
jC3755tAacPf74kkZ2c8ne8gq4OKbVQDOehJI71od/gfbKByQFWqqcpoFuKKEgII
FpiztyPD7mxIi/B5yaOgaN1k1ehtH2i7FOemfxSYZd4QBiVZXi36RNnhYjLFCS0M
iqNm1z7xFHUgXTtlPrfg1ur/wD2dHZK7LbzIUxKlzQ2gKU1fVFO0tZZLYhWBiWDC
n9lOh39Dlq+MhRgibt4RnzgiSEBPRNf8rpEfiWpjQF44EWmy88v93jY278hZCH07
K8tR/g4i4Mpihb5vSiP9GzBiz5G/2N4Kyj2urLVkVGhNuKGMI01X2JKLW1TazJPM
nKzEa+rmssvFywLX+JQWR324IN28x4zNRNyk2cVFyLwJmEWnmNuMqcuhQ7xHef4X
XtJhNmWYp1fjRls9y0yCY9TvmD3D5QUYNYWzjLdm9Qepz2rs6RVaLR5RhCTk6n+M
bMwrQcenvA0ICAKu4zQB6bC433wJ4EWspKcpUw+dgDG3pbAXwxNbsq2UkbhFtpWK
ZT8u+NYXhkTGZhBWl2YW+00zA7aTZXbbxy5gclUP9lT+/ahN/kiWJ6CnBGxzmZSY
le2grM3/yKD64uJHHj/nDWkozBabH7h0BXZFDuT/DrJ5NFcT77ikazteks9GwzvU
2x4a4jlxyDxufG5bKXyCZjpa8MpAJTJ2gLsyK2xwKdn8uUWNwyqm2GGTwiAJY9bu
/2SBLdKN0FAEx1e7gPTteoFazPq97DlGAvmbIocz3B82ec9W7W8fTcDhd1RGvRup
BHlvMuJC1gkoii8mGZlgSk7aPTGTKp4fXsm0JDAW0l8cg3UQ8tYcgWNUfkJjNA61
xztHzPX2Lin8v1oQecwuzEoybBljnZKeWxKZ4CQWl0EiLlCYGXuQopVZg03zfolB
GEZ0avbqdq/oLzaP1vtFqkEwVRks/so7kKCfXq4r/b5vtBw+PAGqTZ1OrAO8Wn3w
cyzokpyUdWrDdXrp7/9KRKZFvLR2R9yLxdQwZh7nA7aklwZZrwmGtoDdjnwMSDam
++uSU3MLrBoLqAzkwWmE4VJgLMXCkWjhcT3kki+Ig0A=
//pragma protect end_data_block
//pragma protect digest_block
07Tc7ALt8FJQd8OYvi3JYrLd74w=
//pragma protect end_digest_block
//pragma protect end_protected
