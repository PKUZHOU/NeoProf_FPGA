// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
MHSG5BeKuxgWd1LEEFlD1IHDalFIJjPcLPRZw77YxB3CpMDxRGxHrkNIK7qOFylB
YC9VhdEQdSpDiQ1aPAoHmqIFy/5ZJw4hTH+z2S+2uWPY8VGe9gl/bevdxuEWCiOJ
DGpjlVUlsocXBO8sLbG1ZDYoh8EOxUdJEh5lIHOas3A=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 18752 )
`pragma protect data_block
kAb/JoJARAOh2G2Oq6KrARCiGqS+CQYlZw4s+qeEJo13R5pgeeeTcp2VN/i5HoZj
nd2c6MeXZthmiGyomTTzydeDCYA+tHjewSLfaM7pQpnPhTppaMk80NB14bOajzB4
n86lBlBd7mBXoZAS5rZPDfRjKvT0ZzzvnmBzz4XyTCQNZyuCo8q4lBPIT9y1f5ar
EVrcmXWKIuKCCnepU0TG6cENTHD/YJN5qehJ19uMnY/JDCVWwrDWvoNY6PFJGc1e
vggcg+4N7JtS9XjnzzqKcwcLJGGLgUFsjrHC6cmQSv++usc2gt3DvOY7RttOrBeR
imMEQYJM28DXmtROc2zA+DHqEGtzYIOtnYosg0L+zfqkvufQUuzuo49fcDuf/tSA
OPNCk/CQELDLJEitSOyAWzQEbPDTFb86acxo+jf/2HktWqVt7huK411Z+PzPeQij
9QfPbxDlOy2QhtJ2poFKHTrRchhGgTq3hV9YIyKaXgYlyiyDI0c/ZjzCW3CgPXu9
DJObwv5Gu2mAw/gQfAw9pyGb1Hvu3sqPvWd+JipizsA2xEmbYc0Mnl00eljD+mVA
N2vWJtt0veRJzf7BhzXlb3RYcjKH0Y2ndkjBaHT9rJb/xz+4oxKQr1h/UYD+Gi48
EV/7QWWnahEyESZZ6ffIUqIZW0M5skTYNqXVqbRrT5TIeFTQyo7CTB2nvK7b8Jhp
BpSZbawCJkzaiyW3XpIIqmooqZU+Afj51CZTyFO2tnQclN7HNmj2B0w2PB0MQRva
/qIdnhnSOGxydPZGEJ9UhBqoJOwXvuBbruWLXVqvzQLHrlHENmohmnmRHtugcj8q
pVk7ad62PE5ICNQbclt4SustoRT+pW5wFgYV8XoWC6mhMvt8/1DUtHuOTkw6PG4z
6NB1tVgp3dxMQcpAfnvMGFtLBCMZBrIjaQqoIkfXDQW5SDVoE9HhqVLksJSMGkG6
c8k5fJIY18JG2oeExaEKuj/llyCmCz5h0jU19gjgYzbu+DAQY48Cg9swf7DIqFcr
ViG+KqRJDEjucSBih9jQmRGlneDKNwlBvbEyquTHHNc+wxCYJt/C2EKYpkaBS/wH
t4GekaMUxbGxJd0fNIxI8ifJXOqBVay3k0rKDCrC3Gn35Q33uuI0CCt6kdiucXNU
N/UJdFHN5PMuSuTprlIXjPKrLA9rC6uy7SMMHR6LO1JneeBkp/qN5icBOQq+Scvm
SGfFZ1wHb9rnfLjlWCrHLydgCXKz/s7eyiEiEj+yzaqCkwk3yeBtU7E3uFjAEBDF
l5tVBV+5HimhkpTTJ0m1x6lNdb8pIhm9KQ1luqwMDLGzGt9fmeNC7YZte5JmDiQI
L5L5h6SXe9Iikp/Rvdidds2tcNSoEDhQw1tJZjfu7miwD3CjWCA16q7xP2bPvyrc
xgZyZJcjm8f6NhyBLLCeCkuRXTgdEFv89p6k6Ctj++LpvtgkptTt4W+Nje1G0xm1
HJHLlMqHj5K7636v3SSFkDKXONAuAOFUxIjHV/pYxyeZdLj4wa9KyvWY1nOD4Sy2
W1MrNMMtPsOUH3Q+K1HiGYKEdTW9YLrEwZPnLcGyb3D5gH4xyAijgk420ObHCeGC
8VfLSIU2JzP8L6LFBpT1qWkFmYQlGXz64Fc6P7tb9/kzmAl+YxQT1Y2epjUMDfi6
XlV5+YSBsxEEI1F2VXS6FDru0kSpLBspmNtxZwnrtyY2Vq6QLzHFWePeJzXSk7o5
IlCCaw21Xwjd+jMx2VuZ3XS7gN3FwyH8xQmk1+PsQQ2FJKIkSiWeleOssq0+xUiz
QZOh7Vx6rtzq+0SRlnwR9y9CH9kB/36eaELx3G9rhRcrwYVf0Dd6ZR9cP2EMRmlP
4vPQ1tKw6PYeu9lxTz9tl8eFg0q0unaTxuRKPyfFEOS1iTe73KfOtwc/bnKvkEjv
LAjJnFx3rUVao/Rey1gF9WA7Cdxsz0Zmc1JaZWvMdx/zknr/I45InYc3wzV4SlRc
M7dSMxKJ9oUNqdhqiSKmmGbyE8xCeXxHemJCizgfF1wHBg0kUa4ryy2xMivU8Qqr
FSAXBBJGXLtBCM6ml9TPZxp+l8YSSb2Xhuq/SD8/g3sO08MuguSUXdh6/ERS0iNK
ieaQ9s8TsOkKhVzdyC8pt8SFvpZ2Ins4vos6CCJH9rcG9E6E9SNV7pa2b3L7gTEU
LtFN4rzdRfTR+0jxCOgsGqrSAJ3k+g7T5NXQYkIy1tJA1hqniO+VPS0n0ZwrFsPp
06NuqcT2UNVrb/Lkrezc6W0yR4vnhLUdgt+QjSwa+4n/IjCcj+GufGSnpyXuzfLD
m0+Ohbco2Do29Xm7vVbHxJVLcOQW2fZEBla9V8EC5clNAAOH6AvJr7WSwS0YaWek
KJexITXSkTiXM5pa8R1RAe3l64sEs9ZfVhKpC8J7FqEJZqeov4vMSBz6cDx4B6bH
/dxzw3E/VQxmaVpwmM15kTYAXneo1Ihqpzg1c0y1DdxFv5mMW7J/JJPRvDrINemR
/CCOCrWk5VXlNdsdoVJ/BddDqSrvaFkJgM/ABNzwHKkdQwDitvYQKhp8DShPTu2W
ABI3c1vHHDCSr9lG2DwvHcx0ybiKjAD9qsHmudS2zUCN0vUqlFMVDMpTK6T4RhPr
7SvWCroyWmTCSMTRILIgzg26ACz+tndI5odNfUjByAXBOj7O6lapnDyTMSKdBBBt
F2Lx1/HQQhnHI1u7T1k+2Vuw5ryLtjxJ0NCM6Qv6R1lF7wJ+zqZrQFbdvHX07bn5
uhy72Z6kaCSKG20bWF5FT1wbIfFgV13V1KJBPqJenPhEheTqyrjpLy04EeY7WL6m
IPTsIocaDUD2tGHxKoLYvZqtnD3QhNiheS6cVdJsG90JEElw32tZuwlAxcI/WfYr
PoH0mdmSic4ehE2eaRt+GWzsRo8hqwkyG6uGQ+BT4cl3OaPOMw2Iz03oD5l+WFNH
0nEDQFGLQ0+zTSSEDZOCjFGhyXrEGFNqgZ3QctvT6EFOXVPnuPj5qoFfpxRdShhp
84op/JYqY3asWNMhBLVeeBUJBv5CIwBC29Cc0GQtmXr8W85eIdvNu+4IHfX0J8fd
W5JsAW2LZRHio+wBTTA0H3FVg3WFu3wUXTAcQWe5FHIzY83v4YckJANaP/PR8Ae1
6y8vdJrCPlVWJsR8Vu54sxQkVWisaCyUweIqaVha2ZXVgii6t/iAIl9CYO2L25ac
f0sLd07PMA+Zj1ZoPdK+sSG/tuTaP6CW9zrib5c9SoYd4R6/n7kf6zdWbqYBGnRw
/wBsH9zD/2we0qQ5QItNs62t1lGKQ05sh5dEiinquKkVeL8tJ5KlPbEEyOinBIti
n9pJ/VfsTdnGH0PE3QBPWh94wwMaYGavEAIT3p2LbfXuPd/aL/YldIUhzXkXVEOb
1dYz6D4hz8fMeCjri6yzV/45Rd38XqjmegsLPGsIZePU9rh85hh4Pxn7azEurNAZ
7vw4PXSWoCNWsZEmusb/7N8YjDSdE5/p6em0KmQqHRL3Jr92q1l80VEtJXl0NQ86
21SQystLee3lp42pK3ySJllxdTkqPPXeviEbUnFmBY7b5EORWz+0cyu76KZTqCV6
YE1tJD48ihBD6rHCc/hb0QGx8Yh48Akgj+HSqmVf3vaDwXgPEO05O+qlhMYuIp9f
osUduENBDf+yc9/mTIa9ApGz0jNnspfZCmpFNrh1v2VTNi2JgPMh/BsxoQ8HtwBl
1xoVIh4K90sp5SiyxyE+ursB5tj7PMowWcOblo6jPmBEwqK1AEYbnDTrMS38vtIa
lwSZjnMO79qSzMY+QcKAy3w1gW4qa1eBFqZrBbND3nwPlKKiC4YnKK24cQsuWx8d
xYMzu/zmE5O00ZmMLDVDy4TbaYfU47ejeAfUE6GTEYo0xUUQcY1JFDjC9LyzXBDQ
tYkrX2PG8rMwFJ45nKsQmFeSCfB2kFq+vv6WhSgawgwa5p2fSF3//kuw/K71qur1
4OninuAK7gLA6fO1QxXcLodamQ/XuSqfGAxvTV4wgF928lJLZP51r0EGXGF7qF3c
6f6BMCOAZC/p18yMfj+7iDfpd1L5o4Rz8Mn5ZRPsT1MXXetsw7em+E+eRIhY3VML
BUw4Pjis7Cf8wEp5Lr8oZaDsuNc8R1DD3QQDustSwOi6KjRCSeRokEYhv2qrFJPa
8lqnP/EEkVPmzLtRsSEX/1ymK46rIb+IWxM5ZzOcsSgTKn4y0QtbgP1XZ49y1yr9
Na++YAcsBDd6+oa1Zb6x7NbsaVcIQNphJIYbjeymz/hMab3dyt9IzC/olDCyX06h
3sqqBNSEBtxbcMFBEm5MvKbYVR0ufS6/X5fYM94OR6+C85oHW3MjGPuYXZGvT2IZ
iVNtYbSx/EiZ6MbOBbf88lVooqICZKLOPf88uvMQIzt2u23Et6kM5FO86JZPv6YN
yuHnVRia9hvkASo7+IreN7Hu8sNTaDodGObg/IA9Z5KTKCYKTj0CNyhfzYA63OAy
qgPbPFaI1GQYyO2FXQeZcmqX7BOj7aNmwodOqDW83P1AGvPNOJ0yrIQgxtAp88PY
kO2mngJRQJGPcg/jd6CBeBBESuNMR+PAPgOqPFfXd62IX+yDAJ/kV56U7RhDlBV7
CzF9DkGR9BA6O+L4mxKz9XlERuYqyMolhvFhirCGeNpGdeFUMWLZIEpETyh4HBvp
1J5heJv0T9YxBHSE7apZpAHXweTO5y4IZosJAhJ6GD/gy0scUTaVDyPNVG3cWiJd
i2YNZmvfOTSej4Q5LDvoAcyR/8OnI/LAgtcMlWZZNXtGYzGILUyGNwl6B6rDD3QJ
yT6UL3m3IXUlSdaMafLx5uhi1ij5GDyH9b/CIU5VUMBhVpItWM+6zlL0dt0QMigG
m+dbiTfGzzTcKSQcSaHYA1s1b5xouL2OnDkPRKXk2DYK4vuzqvE2CYSVNIU2MZsk
k7BH1EbiopEezZOlwPjwsxJO3KC1AvYnMdnJ0CoFOZMcugVLneLfNYoqa0gQzDP8
rwBst/mkgbN8KEDomByh7cgioZeXXIK1OnZpH1FE7lFrpfOJUP8OOBGDEW/D9iss
lAYmJR1xkXXRJudS4OwwAkj1nbYHtEUJuwcNxcWhZd0nwA3WpFOXH0MmVGQOHEV5
cK5jep/9KNAerBhboGHvwoxKcj1HESi1uY1u2dh0AfhCM11HIDtULrVxbUCxFfhe
54Km1QHbSn7gfpUzBD0ara47SBwiHNzWjovJeyHrRSEfSx/WxTBUvndwRY58IhMg
9Shhnr7BJ/xFy+TfD8Wy1qCq1rAXefw7zO4vRHAUtsSRfoF8p2mpZ+TDWiw1GXkL
gvL4wcG3AhFYj5IPWR6Y4LR8RqwDD75nB2bezOEPD4Ea521b2HmqIRgWhfqFbB/C
aK0QAvZJznRclHpBH8ZD3084okfUx3wI5NYkOuaDORn+uYNLIPB6yGo4v4McTrF0
sRUGDiQ1Zx7Yh2pZXDZwAmo6+ykKYnCY17AW7iV1LWjpCZzrSHLnv/ynLOM3quBh
jn9PXGRuSyEgo6tlOeYmkTrp6KOWZ33UD7ZSGPexhn0pB3lyVdQhVdBR3FSkVSY4
wcIW8ARBXIvCFRCGx1/SiS1S1/VxcoIFr0kaT/nbTXToQVOIHZyRujxxOLpxFwgw
DgUwhzG2UdNhXkyIRoEMFuyBj4wHu7g/rtQvMLy+TKXtWcKwzh+bgsH0MD/6l84S
sxJqEeSEs99qaq0WQYC2c/tGdGle7G6cBoV1EWZJ6Xw7QhL6WAW3vuOn6GWRudyj
tdVin+29f1CdGmEjJu6fAFslK8HDoQPPfzQ4V6xpzi3uLDg4u0q/hs7k+N8dhNFe
Y9moJbLYnEyATSwfJRs6mpOtZ8Wycl207PeWTTTq74d5suv3k0cFiE0Y25oQkiRX
IhJrEQ14QFBBdXEDJ9ipZm3D1avspOqmMXJmL+/GFI+WcWEIcnL5uy++j5CxxUWY
M1xAKdkN3wHmcQOSogfXJmOSkBZ/u/9QTjTz4auzLhF2vdPakfFI74NDlsakYpIG
l4jqv7HAkQHL5eeX3tI6/CWucrmAjlg8xSrKI4tNejAgmGPyh2gNG+bZz7e8z8GB
jP1kCnoF/Zrc9P06eaM5MgqKfOwcx8cNEapjZuevO35xKn1/v4EN+umBf1j6qii2
2lDIiaCTu1RmLc/LPKrVMGUWFERd4Nnj1dVUzmhnBJqUNikBYAdMVD4veO58t8u+
4kVGi0K4OBENIDy669MqSH8IVj2IBwiaBb8xat1LBVXLZAkxPHGe/nUmwhO7D66C
3qTiS/aWJiJpSa9wLlcWmsudG21SQfnoeK9xISPVuSqmT3QFhfkz2Uxks9N+eBKW
kz3fFk3I/nGwjgduETlm+4uKcKTldrXRW+Isu4R6MxzEUI0g9QJNwri+1aDZRjcc
y7J823WJFM+zLL5AYvlwHSX9iDQwK36QhQCaDp8fUW7eoUp09iWs637H5MSMa10V
rsoUsEsVbFVrA1iyBNHa4bMOezRkH3qfaUSnKuNiyrWu43vrc/9d3VjNw8XbB5zo
xZG92G8Yxkag0mszaK25Mh3vgqxYXGvVFDpzOfszkSS+BvGAdJqoVm7D6nb0Gs5s
7SEbVQeAm8LQ5ZREwR5JafYcPN4oAXw/TmpY4PCNVXOgDtgBsKoKYwyWsOG0kaZv
mGiifTE8XgDDrAdyiLJh2rex/K7SR4YuM4VanEHKtfECyYUj9q3wBSTAi0MwtGUu
ZcN1Yi1MnBpwSWjEGf16IvisSHyydqH68bat3V5NKdiP2RLdlWNuSIpFTWFZRKDF
/HydG4ufLVJWbsxiJnzIgIkNMF3hAP89T/H8QelZjpasvyjsdz+UgCLg7nYYCRHe
6mi5suyPXbP7oF2QTMnO+mx0WIk2oWY90AjgZ8cy+e8TuGpLCQVmjAjoLy9YKD9T
0EEMMDGUe4gbtCIPy8cxj/LdhlAUafAKlEdtIPn6V7Ar9QWtTR1FaEPdqnHQ0RRm
HrvWKvS+dPqgwDJ34/iTzq0svor8RibCnjWQmx16fk7VfcrJtrrHepIxBkfzBIEH
2hozBteaN1zFteL3lEvhcpzhiFd3sy+gVA+K9b4MqQhijlFi/icPVZBbSnGRaaj3
5PocDQFsvocRv/9yB9n78PAjrSJu1u6flQ6QHOxo/rywPos0lYuC/ZYIBaShlnkm
Zcgcd6GZp3fS57fxhT05KJWgxkQInNJBwf1GphA+3YzTMoVFW9QOKmKsEMvRGXJu
KRrCIdsY6CtUhvnQ8bYVKd5loTLlBEmh2o6Kb5iE0tXnA+zZtNJerecUA0BiLN1h
Jft+gmtKRkZLBn96tiYY6l49u9upElTxcfm0+k7oT5nux2K++NXgaj8Lp1TDlbZS
c/5Ix5iOlle7j10Efihqg6piVSSXH+kXK+xBP6xdUpjoOXTuuozoLwJQrkQBJEHL
S0CCbGqejHDT81ZMwwv4n0+U7KITnYIOZVbUpzYI1Gcy8w4i66j96hPP5HB8IL7U
VGJwQaQErV3REUgNMVdONQxx0JidszYXZe7Gl5J3cCxOnK8Zy6cVKyugx+e3Nc3b
k2ep51+tkurI+g+MMPtLx329KD9mofhkXE2/7OCCHAMJtUH2zng+umIhDRLwP2tX
U1PptblMYxJDZ6VigBaz5p4oxhsx1zSNjvezSpTtJMcE4Xui4ccqfO32R4p8Mg9l
XJYHUanI/AHI/RqWEfPWTIGcopGCy7SZZPfK6XsIL6SfyHn+H4llHLB6tKpuKewS
kfY8mU5Set2NvBDGxS1QrcD3ROFHeOJtBQ0ON9pIpMjs3vhK0TGN2iS+g6ZzA03R
OMBP5OoN0oPsaKikDu5OlOXKnazrAAYzAbO0P3LLHZQ6rp3VCHKgp6aUfu5qUMDG
84j76xpYGlpQbOEg/b0fcTGQzcbh73H70E+tnOoXv1tsYZ/Uc8wYVQ/t+j8wtl1t
APyL6+dQC8PeDkPNA5oiiMJhSRyCOw0ihVbLDXamJ6dx4M/GBM5iaIzS74VYzPRP
ld4/Sp+4Rf5Zwrt2ot00uuQwtaTGdl1wk7jYF+X5yxhDaXr8Cu/bgly5XXxOkvNi
JWq5tdvSPvcsh2R3QhNDzO2jfrC3KO7d8nOnv/wBzExl6tij+7KR7tV2FckvGDoH
ypI/j7X0ZUeL2fx6E19CS9w/ZPlUK3DlOiMBrujdfiasM6cB7CvxBuYoFe3+w6ma
JejBuz9laSVouoCFwJqpdb8W7SpRLj1UvwFpbsvE7mDwgt8CVfj1NCYGBQc55P/v
5FvQYQAdug8epSTIQ/3jhu42fSQTRk8PJ3BuFkYPUJfV1HuMmH/+NooQV1x1ArK9
k9fUyGUW6xd9Zj15VcA9TK1SU88gJPdY9ux6rah9pgq0itFjBn+AAvUfuU6nJoe/
yvuzPzqxbXhKYpzXaE4QG6MzQruSt1Fys8rPqDWxfAwNGWWD3R5tgnxchRjti5cG
Fud6dSLAWfQc7LwkBzOzriJBTn6pTGYaQuUG2V6XjYkFCIoXLp8mi7UtodScbSKh
jCXmhgkIL1u5BBDuWIjKl+Ah1pwsUxhNsOyQoXeG/XaxkRBbgWQDGuuBF9ZcTzXS
+fjoNWMNWO0Nb9ifOdRYrcHKSj0DB7cEXE+CIPQnnk4SYiY8PAGBdzdp7hT7f5Ee
Tmo6jgnWfilkfWB35I70BMKzA9ZgU/PZjXOQqZyuA5QLP07fGCjA07HrcOF31ODG
rULuIM4a6OUtcltqs6jqCYzLzUR3QhjNZNRNbhmLhBYnAc0B5s1KKDuqh7Ixn/dD
AjWsyJ26TpIx0NYn6cz04cucsJcLe5t4NvzUteqhwBrWdY6bFquq9yC9dfsPg2q5
q7KRWMoEAZ2NSXaBvrCMUIcrpC+5kSXahILAFx6eYSO2gdrJPobyuoE451+fDGHn
WrRRNzECPeWdk4nO2K52vAFCDeKg64tQOHXWHOZtgeE0Au4/iciCQpQVAUnGcpY2
zOTAyHYI3k/4ehaBE1BGbmR8MEtVinLk05ILRxZtcSyKF9lqRptLjljcp94iiX5S
7x660xtXnEv4Sk6bCgC1vp3g23KaREoRDJ+q8qSXmGTM8iyG15cGvvXb6Xz1S5gU
xNBfbm1SoU2BQ1w6BJMWpei7iImj8vsbDWTK077ubd0omqxw4Ab2mG+Sr9cabqM0
mGNRT9+s/SxwAX4FALFG/34qgbgir/bNRNU4Oe9uZ8s77h8vJFD2faTzaXorVsMO
o/cg0lkl8Ay3oHJzdQcNUmnTbzLma0WGoGXwvh5Chd1rtXllVB6HFPJc2oiUfd41
FLldFJq1dBSEM0EI1BU4TVUJOSmgvAelhRYYqxQTAPODbDv28A1vW3RMf5kAzg7o
D4Luko62z2lWhX0LGStDLmOjpHJMPKcBd2+a7hGTbI6zBWe3rpz1o+pkygO+PwVD
2smZPFdoYOXllqUOrkAoj6P2JScTgDWjzSoQi6S+5ZK2OuYlAQPsBaosZGTQ8W23
dfpSu1gG3Pgeccj+vU47WVQ7HD9grv0ztfFBgx4Hm7rSrAd012cPAWq0EOgNdWY7
rJESFd1P80oiMa1GpDFEAOqHOhcMz+n3BYkM2pr0gV7+go5Fct5muLz9XR1TFBk+
Q+7oPaZioUALVOgc9x7B4rJOa88yfoU+i5PXkdXOWfXS0q+qd34D0mVPZ+jrM3P3
1YYm5jpQ3R6gS+OfR+C6Gagepa3pakNLGnbpUzfyRay7gW6S/fbOf3FnrMm783nc
GMZJo3kMBn3ExyloBn1uoW9UvJjSFP25CgxbIDoVzI61Bc+BAHcjamiZAechtwiP
ydLm2rBXdFpcJrcHqpQkYaJ5ySrX+m2lSJlq6EKkXGO6dBvjrIyVl2l8mAyLgUbE
BQqHMYYFdQI4L8VIHKwqMp88Gq1Xd5bHqygzYB8SXVgxXPVsqzcEI9Vv+1ZB6Vfy
pCdIibmpC83D9mX2+DJ80NLJDpegyBo3qj7Q1H2OO7sqaGO/7QQxVInQjiRL/mCR
KMLLa9sd2hHTGqzB5v2fjB5ZpshiSWXjKp+OaRUWTfN1rlQ642SAlfiVz60VzcfW
f1Hv4wf3v4FvJfF4+EBbZ1matzJzADlsQ/ORQLTa80SHJh9/FgwuOBsGTZaN71VG
r6DjHlqzs1aRsIdsTY1V6C4rVA6mAmrywBtLxreok8FyQEdicitVTqSJnui2208J
RMu7e3HMVwekn+Qj1rsPTWJZfoZopgtGDKyAZEa5O136oubel/7CD+KLiq3YNLrK
+S+EJ0HDXpxD6ohavEH7A5wMmZQVa9y/pmQI+X6+uPGBoaitpFA4Hp159HvUs1zB
ZMKsTWeBkzr4Abyo5qQbQgC165dmnEj2aYWcB/CIaPllOiORtW1gn/wB+judckd/
9VhYi17JxKHNku6BJ+sF+HMmrLHylj5A5Cd9/8QLChhdfIatP5mula6MX/++9fxU
coFL1mjDjf2HaPwUNEvPemBVdDwcKHH9hajJSSjam0cUDcOH3CDJdCsEvhekPwVP
J9s1bMKr4YmTZDNFxb88eePEq8YbUM/sqmQuOGKn/0VqhOuUCINHxFTm9RiILNLK
dRInn4sKxTpeluzcv5gccRFTkTHnFu1Q7Eb4BY40zG86u09f8DPcJpZWtbxlFIwW
RT2CWO/9hp0p6YJmDrCE8LDj2Q40SFkZyFnp1Xm+VCArDx9x7ceFaF0+ERazAqXo
o9VkGPptKa5LRXViTJKGxaOXpVDPJ5PMn0+I6zZOktaMfXTKdyYEz5hOSkz3QV/a
vFrxorOVTpZw3zcmDKIOPrtZi3g914Aql2HqgPi/ylDrhPI6/lNEsTwJW7cQjFN6
Y2txvfRzZjMAj/BCB6l4+/wBJjzaw1alWnIXhcFDN5IDmNMywFQau2/3KBeap7q3
v/YJv1MuWSO7lGlQP0iujKhXIzNqJXWk6BP52ZBiZOBncnLKlV6xfbuLYoTH7KsT
INUwozBKHKL8Q8aU4Y7JiFyyzaTL9rVSSiFrDGNkAEb4T+lV1mlPb5cKJX0bbwjB
nxRccrj6u7VzHgOT/s+WYdBxN1q0whv7D9dBD8MSE3CeG+6Z9q867hSUDgJLmWUh
AoYzp0bwkh7WCSdg0ay8ygGYCp67qxTUIwxK/ezAIHgdWMc48QO459hhpcGzvyW7
QIL3HVWF2WHybMZYH5xHzHqqzymk7Y/g6lzt4uMV4mTB5tjzdxOgwO3i6AqNRUNa
YgRuPwJAd3N/O3YceqfMK1OLqpcW48AxmZOG6o6WXmxqCTVLF/WcHGpeMgirQjz0
K3BIY2bSbxdKigWgrez3Ffzv+iUgjHIYqrxPQdyR2ixqaI6o9C0BGF9qbHW8IzLV
v8ZnfZmjISe3BZgJIgHe089lbM3Cdq5T93W/dQlQRBctAZUZLiRcO2OqprE75InN
/frPEHLSGWVLoWS019dRp0RtyAYtVWG4OFVuzJfJ57KyBVzyZVaN5UUaO+LyeQE1
+2xsUisfRS8S162xgv2AoOVNdHxwzAym0s+v2+InmiQhqEOd51bh9yR3HiHDq8MD
XP+fzE0ldOkX/eRLI+TnAqa3XZccYs5MHvnOFmlBNUE4MNn+pkQal0ZfNldiuto4
KSMxz7BLscMyOi0l5h3hzwIJWAazOxZQ+xWEFXb+ZFF0lx5kOfOdXyWKPvuNut5P
21KlojDOqoYy6kOmQksqI8qQRfiABTMPh5ArK0b+uYrl/pmekhw2NbwnmSC9DeS+
a3hD7aC8kjpPcNvp/l1l92QanGNV9Em2ikN3190eU1O54SZrUJ9BDYRjY/d/urDh
D08L/GyfnjYbW6apBLQfYAxdIOuDb0+ARP4P1tBpAOXMrOwhqvURDtKVq55MfWG2
Of56A/d2LEkUOckb1jn1DL7a82fqbR7xN8Xrr8MHWf0JhB5LqISXEamt3X1+vkEZ
3s5Uo9f3ixXTLQgmjJvKq66OorvJs1LiiuZIaCrcqmwXMRtCIV6/zI1J0Dfha2J3
M/nlhr28dAUUjKSomdG6i3jVljsqQweP9KPjC3xkRcqKAaf5kQB25XwcvdkCIA8t
x1W+ZY5ym/tIfnCnJfmj/lB0kCm/7W23nJxywolhto2Uz7BocSSLAHknicsdtdKU
G9mGMUVU8brHN5Dblp72PPJSDJWeu/qOU1O5nEVN6V06QpQsYdNLCIluomRiudc9
uoqulhg9g2TPziR0/7iW8vlMqX6QE/CV5Iqvnd4jAMUzcZs+ohUXzKrTi8Kz1a2H
mia4lgh6WPa7LghG2JZtBeynIQUxLlf5eAuSWOavRCj7GkWPKByBjsAeAoZ4EmTu
e5mFPbKGcV5qTHwCnS7zvMz5/onUAMB/8AFtHQ6jCgBapHcbvE1Be6wPZBNqgN6V
vzEHQjYUjqxAKJlxlMPkZEcfbPFT5bvbS/7XI0q+Ntt9X9vXr6MJToWWJCbIBeUh
jdsom5ZOCJO4YfXj6EhSa2DMfh7WCXh7kJWY3YTaHFXdw/VtjdYk0eKzZ2Jh/YJR
WZLBqMzQxPtyx32CB7uJwgbq5U7rOjfl5cJGi5HxY/E68lEyERtZoQcODYCmIvQy
sJkG8KKwFc+WKiVP6y/M04Q06SQaSJESyfGy/q7YLdqo4VcB38qakSVPnFgQEULc
Ix+x9IO3JzTJ8NfQSAaxmmj6obxkVUeFu70o5K6UHqzsd2UXOHeofGOSXiM7y/A0
Q/HoObE9KGJh7ISoaZ4G6cCm05dEuNTPY/sn3Q0OGLwp1na5n7zyBWUNXp21fyhg
gYsuJo+HUYiUA9Dt9b+vZ3voJ4q4E1PE8x1VydOy66AkpeVUBjHwRfKRuoMgOLp2
E49l05+5aay5XtqMItrMGGIucTxJi3CVqIXpKZVrXxEVmyuKyyozZvY4lpAmJZYY
LyvgF/PHQMbfubcXWi5lUpG4IxfKaUXk7Ak2DTSJDVVjEcv9HGSj0wqWgp2tn4Gm
SvAFDKUWhpysfqvHp1l3HQjo7dxQVMc00+2PsydKHleDxMWk3KhTDOhohySpblUd
zjd06Bil/u5Ykh5Yj+vXe56xc0I/uelFXbIgD/nHRoJ0weyUNqv2Xmgj/fGoLMQC
JD268BlJr+X1HvVNZV3OXYThjEn2nAF+ROiXLGbgZ6Dvbi/qMB75tn+bthol6GmG
62JHycvUfVpXWp+gUZacGusgoRXH0KjWPgtPb/cppP3UpOrR/HfXNZ+VlIq3IDZH
x6VPkspVpyznlRoGGtOxuAbm8uVfrZI32l45T9X5T+w8ZUkE/n4U7N/p2W3ynoFS
ht7kzpF7lSWhy+auPQjlknSGs/BmVRZrzyRPS2W68jAyWQvJNwpn9TVkdO9Mz7ni
cJJsJVvKvMjrVHuc9oG1I5bVKbP9mKTzAH9TqR+/ZTwjgeDynzBUpBKzInQuwFhf
BMuJ8pfpcoFvUq+hz9TnnFahhor2FBR+dbMg0SBjwSu3lLJ5RTgA7MBTwL8kx5wq
OXZ65vl/qiiConr3LRqIzEYCt2gx34ZLcl+QhK8fU+VeGbuFZUUuPI7Td+Ozmh31
1+RohF4vTLHUfhve2xP+DL+U6sR5MDJNHBmySXrtGBNsqbi1YxlExJm58RfTx1vb
n/yCG/fuGAFgGaR0y90Hb62bLKVf9iWFVqeOBqds+YgNwMKz+VEFY5IzIvYE64ij
N2NIqaYWUMWZaQcnXLt/5FOrHRFOqtYaDrnqHHcttQL7WEYJYXbf3I900pa+Ihsi
49p9H4MjqYI5mx4vnpFBmRocr4gsvZZ/5pBvgUt+36GTdD1JKiilmKu9DSFQ4ZeQ
fmtA8ZfZmCKVFvkKz6u21AXNC90dXilFgIK/cYVM4eOdGHKbu/Fpb5rJdDyeU7RT
sue6ST0YUggw+osch4VWKqXSAcG2/JH3MXKMUNTx8MmcnV66ewyFXp0JVvgcL6fi
WUMKpsAGHmjxIRZ9/iIgLr/dszhJmDE9PnJjaRa4TGJ7y/vGstw07rB5DjfsbvJF
Jkf89YY/aL0hPboBYXVT+kd4oYTt8+PCkj/li6pd5V4BPRuyQsC+nNQcDfavx1xR
37lWtSbZmKgk3T/1bBNwD8JGFoZcWomXFTlhMJS4Tj5+mfy2wm67X8Qfm2Imi5e+
xSOxr0hDyg7rumogrX8bEfNR6KrTmHGwbTnDafQ6l2D4Qa/N+gNfoP0G2Wc3zveo
2IeHp+amZNrnL4XvFvkzZzRRhajZYj8aWRTadRVnGdtbMe6ufTz2r+3tcbj7mb3b
ZuKAiNmth1MNUBFp4QxZlOwj06qt0IQWpFr+rqSoxT4lMytTod3i+Vi6FUZmZhp4
srbk8JhVKb0eycZoouwG4Mpq1TCRUYO/d/pfwZW+c1ijCF3raSxiHeLzrRh7aFz9
ysK8ilUU3X6K/yQTD7LA/u25IIOSNVp6YEFIDgx+Md9s0qPJS0Xl8vo3Cz8NMPtS
ewzgUDapUGPCMKcdvJy96ooTc66DqOhSOhkwydMSwb9IJ809vGmpSJISTfyMeh1q
VZtYJHq59bGwN5qewFPWQCN+RA1Q6LnbBhhbbNgYw6E2TZza+SfSD3o0OO/Mnlji
615d3fEMsmHHNlITqWzffRq4Ysqr/GVcZkuMBysEVRYj/cPXObXHYLtHesIQdqyo
GdIh1fF1h7tIZ+0dDRMD5gt/m+P/oMqag8t+E/MzeBhy0W47n92ZQSS5Z1PxRE11
+YNQSlKN5XcmbrhHpgW85z8xCorYDIuvHB0nR/pa9lmQf1hbgILLUbBpdFA+j3Wj
d1as2ZOH/f+6moMk9p+24xcOTu4IE5/xRSepGZvrYzXR1EmZdwMQAKtBVkAv4zTp
fEGinydX+L/b/ObJ8VPFkSc4SmLZxuyqvdqyAa2Luz9rCND3ZZjE6qV+Dqa7Sls1
s7wAR+KIWRZxicjpogtxJhMpzyurC++xeAqnWNI3f/wwOXl8t3Himujgsw7J4rD1
6xLhFH7JiP1JWosago9kaaLbEWwaeTzyufCGowhZu03+W7ZEiiLnrw3joFVzcxn+
WtZsJtnK+JvYMyIULwB8WjTNmTv0BrBZEsut1fuRGduFdYOzCcQGoBgBVkOuxdtD
ZDhbrix991F7HMo9yEvdHBtmokQfWQ7ZZerowYZhP5ounmCFb/0BcIgVCsrG7Nyv
2J5infqDNh+JrL34NyNEWILXGnRzka6de6783ifY/6Rcg0gud9ffP8ajOSXOzzmH
dVGcTCL+BvBzvOmm2e1kd4HxLgUBj0+PY3fM1j/Gk0urFtlSc5UyuVj1N3j7R1Y9
6HFGwZ+Xk94Noo1b6NhgGmkx9htgApd2LwjDufLcEpSs2+GVOGQG4LtK/qBbAlgI
ZN60DOFpM4YuPcAmzmGX8QMZHzJeb7TldtZYOOjn8pMaOhonWUigZj+ycRkh5TBT
nBk4onQXEmjni7/lUwfHHtQDPX8taVa8qXvuGtOChYH8QNOcDnAR1NbF+rjNF6fP
NZQjPUBMai2SgTI5jcx2trOP7Wt5gOH9mrbvkNY2pwyDkqHyqXMOxds0rzMh9vIs
NKI0biBrFcSONhkipa7Ni+koGYpHBTd2sY3WnOvV4zRKXexKeU401UebRQQFe7UK
PgnFVITJRXkSuX7GEIhHdAAuZAsETiVWLbqnfhD4am6URWNbJlMQlF2c/x8gqHfR
5LsBXOf2fk8jTsuJOFMO9n6rUbmMRnbwVvrFOrdBJXkuCNaP+2bsAec+wi7VDddu
3O5cOf50F7BheA3mC+j37yuGh8lSsOtgL4yfqp1g0/yU1YwZVoeOI3g12RJKSWHi
uRCZ0727qUIR0sHshlmfEL6rzlZ0rngxO6p3zWEBHsfZovZlzSvMSOcMTp9+zHK5
Et6e1rOmMzuQ3YJ1/h/1AiQgvKe8HqWL3GDD7zTMnPcybUCFJz8uuSbBPSw3o6z9
z3cldZTCEuVq+6XWflzue8GKk6w8AG9gjpccfHfCoPa3KFyS6XI4wW11C4PqCo3+
QdR1iRCVtTStX8KpSTZufb+SeQYc7kEC7OoKLdxrDIWvljZ81IfdC8aJ9jUK2X4a
8YEgb9kmYQvDEzrQTxtKWWr31i3wB2a/Ijk3gyewGxfUlZ1a6CVCuG9zUjNGHDot
matpSW+fXeudoN0uHYg1mu8MTxGf1VCDdMM59iNY/dtB71/xrSu3vPVwJ+DWEKSZ
jRQI4epV/1EcpADlF9SEkocKpOe4u5iGEF2dK4ch6vsORUvoxzyxjgicjU09NFIF
GVpUbjSGnUqR1JHa4Rj/64Q21MqM8BVot9XZPZeySH8uwMIZrTHEYjfRaYP7QCKd
5AzIikmNKWLQ5YzqAebVGa3zJDm2TYAYy4fKP2ftMLv26yGmfuC5yum/IVD5orOF
ehtA1S69QLmq/ybGvtkAyW/URKjcgJXN2A43yIpkKA9X/8mP1WpsNoDIOo8bFnDI
gXoqlSLd1mNNhAUF8eZxzY8gMSXhtOLyDewteK22uP269uH1GhR6zizMIDoNhWBe
A8LR5oVao1lzgsuG30hx7ISuMty5DiWM8yxLHXM6sH7S6vd9qVu6oxrzC4iRrzzE
h9I9Wk3VTsUDxW14BOma1aqFP4Whfbds1Wnk58hZP36/CRSTq0XYKfCOLhQw2j/z
IxTuI2uzKiSD3/Z5BybTwBmObCro8FoGeS11b1z0KwOlccJDQA9Cf9dZQ7e+IGEk
bhA58Zyt1AubHHDjPtjahJ4PCN41oPNGiRi9TRIMEe2NgrXLj/giW9GrsUtD3Cly
IxL0n6Gdz4T310YHk9Nl2f/Gf5pDe46gQq4ew4VBDcDQ8MGKeWRsA2Anety5hZkb
+eU7BaDZXNWbAaw1SoNgyICYlNAyDyNiiT68JMT0e9p/DuWGweakwb9zSBINCVs7
fNUy/YtQxA2erjys6vJ2X0MWbsr8KxqNZaxZYKvxVH5Kn5FnR2etKlzY0UpJeBua
9S3/jeVQn1haj/AYnEEh48vXLk7i4zo9XjqyrjERo3+hij8jCHK/fVsSPUuU+BJz
ozLE6/IC/svQnDu7zSaOPCD4g5t49N2zZCvrzuyFKq1oKnQHvGZL+0t4x0TPEnvH
jD+kMS6Q5fhrNeFHHH0YM9f5jdh6aqhzLDHsNfKmiDPtLElGjz2/mr765b24H04P
B36ML27MGt6LuT0me2vgIhbcw1N9961CWkbW8duSXfMdKiNT41he+Mx0IrjctBgQ
k9JUDsVYEHAulpJpAkCBv6qEtp8slOu7RFThwmCtG57yqdHLMKH0kCAbvVZxFwUa
zG1zp43P/ZV30fmnkdT5hlZtJznyMZzf3zRghw16ALTjSo8ZxHcML163oAazzSfB
8lxF/xAg4TzfQpG/994PV2GyuEEs04YG0WAnT7aDGPB+p5SAPEbDhqOOr7WFoXap
MEjZKTJ1M5mcPlxE+OWd6XlAi8PjOMUT7r3IOW55rXE/qWUETcKWHuJvCJXXoE0m
GqggXkzlSz9/KUt2GC/Ztsbcj7ty6+7sMgyePiUsJRB1JxPVIrNUV7Wjkiq6+i2f
FnLwMIii/48UtHlGyuOqjGNVAwLKGzmO3wgvUSuMTFIsszc2/1BijJcY//5Thid2
Da81hByOW18vDouvSVCIapVsLFQ688NgoKT7asLNgnWxV6ef5FbA9i2P0Vpbqvnq
erwFt/KNT9UFflm2ktlCu/BdhbOhyASx1gUvrFDvQ8mYuzcy+5I7UdEbvRiY1EQN
Hz7+DIMe9MnBYDIe4DU91IE2YOCdxf50b61jNsJzc62d3LJdHtawi3H3L+0+A8hG
pOYzTif6ISOUSsxbxSKmZjDWVf5XjmTGTcptoDks9W6sT9YCDu7lqBFK2liDFER0
N220aiN55QRG4tudqF4aJGs8Huw4Nvn/4ycmSFdhvo4S7COL4fJchT+3va1OAT41
uAtB+Yq0tvyQKTrUmTAiQ4lLJwtyq0cbSBHfz3RLbSKUlssuruH2YR9SIvg3oZGD
LFXG8ZmPRd3tcOcSprqyg13DNb8kpJw12wKlV8qyj+VZiUp/Wkugzfyb+R1RU/pm
U2CrbgbJZo5hAYvP81VznGYM9bH4DIL2nS1VWubqtIC4tofPJ+El11H9emsz1RxW
+9tJYtKxFrFe0W/CIrfOX9jQrA6JITis9BDU1SxCwxzI6E/2i/nHjDnrdXBUTJV9
vvyTjCtEDnxlRM7C3ydb0+tXIOIIREWDZVUF9yQMVglJ73MCIURVKGoVKOiMTSl8
wTs0hzEBRmafStEMy1bUuH0t256Kv+45SCbaAXpT8xjMvuYWndPhq1lumfz1LhQM
dg9BNqIVg9E1MJXBj7IfuSTsk2gA0E7ZUnMS3AIckS9oMwiMzVjvRktgXJ3g3u3T
bippDDg6mSj9vqaXZv8Dmvrq6kZLzUf67ZyTQdj41ITU/N60cfzL9XYC1COZLqZe
vUgePXoUZepI+t5Vxx4pz9Osj7PUQOT3T6AbFhyn/C8GFYXwG0x2nbxllpenloVN
Xg2Jfl3luG3rCSuzV1thlsDPq+SCIi0rLkrD1bGG0qf0CTphe8I9DkMn0CuR/ZHZ
qA5FOgdcacZlm9vyz9OPCRt1R8VPyhHcWGljsjEf3AKBnF5h69tcjg/qRZ3xqnLj
Pczg3ly7gBuiNrXR0rVxPsjxJr5qCoMGYmsD3vnIEgdeU3BOYPR/PM/CvGeGeKMe
8Ldqvuqraz7f//JqhaZCe3a7uH161ue01re3oF7OcfpkMxc/lHoZeKWY6UuZF5qv
p1veiG7Y+5fXRNSjMBsyLpj0dMGmZGK9MQQemOkyayU/j91Qku8sQbBnBfrPnU+O
nfWftYLdkh5YTNNo4Vc1H+D2y1FE0zSgn0zsCUec4wM6sWw+yuky4PeI5r4RiBER
1c4yIw1tyICoacI49X0i1i9u412zVIz6c9143CR8SclL8UZKu8yjTwxIZCkDmGyT
lbqxqFIrsvnPvGQwp7rQPNI4x+QPVLDI74NZM2JdiQrUN7f/Y1BZWJxoLMSE+piE
832i4WnTAXTF8HLoGbac8Vcb94u2FVNpyUmvPDgDxq1IrlKQkrWIYiAKDFLg4zWV
CMnHft366Ufl+Vo55RyUgBvmhDK2klm3l79WXd5VtSjfwlWCmnWf0i7VZ78JvAh2
QCFgK+7RQw6O254LadTmeXtXxsEi5NCNfMZva5o/11r+gZdjzzfBjl99tOQMsuvd
1kKBSzTmquzk9KI+0B5uKVUPInhk8E5M3D6L2A/LoVlItRx1M7+ICkF1AoZOx9+M
vwBm6IzM4d+v33jCnmMuu88lF3l8pBMLr/o03L3Lg2YirDP18sBmecWwMe5iecKg
E7lvSfDURGrNFfDOK1iG/l0My6957DDNEb+Zv9VMKl8Z3H8ZRA9LEgLgEg8T81Fi
fDIVj5q4XCsimYveUAI0G7yCWl+n4i3ilr/08pi1JwXNReSpeLDr0jGqaq9LV1mJ
JuiPtIJbwPlVY7HBcxWzUtWp59eO94elJjWgi7M6gR8rePhcX6EjTZTF9iE/DwMy
BSIrWtBewzNX2aMxqmfMf5rl0vKer8SWyk7pO+W3R8tE0jZ5/QVySNksleqlyd31
B8WpJ1DmL9sc4WJDjZW0lsJQ2Ohc/7G9vQGaQH8nyqAeKWG9NCmnGnLbGsEngJDU
OkdaPS58JGximft37EU/SNWzTa2E13g/zTKVooGKDA24RlVRCSq5NMVO2yfeJf9W
X3lpChW9VGgj/kO6dLP/pDPAjLgbfg93dp8SbZBsKfvWZfIj1VKKy588gqwDBerX
TDwBrrGeM7xSFBiOisitgtyDoMD0c+UKlVw+dVhnlhVh2ueg90Im3vvAk1g9ZbkE
zyKtl+n6Yk3pNU47lj11mPH1ng1OJaQdkLTkZNSooDi/q998l2QYbWxIsizHzUlD
KBep0+ew74YifjyUfBWq2kU7P8xzyF1flQOS7uvRf52ZIn0FxFMSIVdqa+in2r0u
ZjTWXtUqj4EzhR1w4DNbM6MmDyJ4M2JSA/gRfEXgaJ2QZasruBxLdJa2AwHcGoyT
Mlyf3OOJL1kz2A+qMoDuBIxMfK8v6dCuQbnTm7IaKtR0LUxj7TOZEPBbvAda7o5O
0Usl+lIc+FfA44BJzCV2+ph/wBGm0uWFRVp4zGuO9z4bN94BKQd0+vYU8Afyg6ya
JjH9ZwZrRZyzHd0nmHX2OVZwiEym+L1mM1ftkEpb87k8qMhks0vasynUY3wnqrZQ
PRS+WlsrLsQ7D2RO5zQihwk5wvOm5tC8pOsqOAmp8qHcJvKxh16sekoccpig1iaH
Cx5ibfykGpYXcdWGibCWU0rBhFbmEBxhj+iivnh79vDTd/tagRQXyfTSwMEs4/u8
SAL6N44/7tBBBtVhWKD9dTaiHoM621Njx9ymPkQcYmwq3Ps9yhCujpR5ir6U6+Dm
kGry3/FvZhKB1Joj0FxUPxxfT0K1ZY9oLETCpV1vsNovS7U7WpMFL9wo8T628UTt
P0QKWDeHppFgXK1Tns5xuh6Zq3HkHQccyWLc6VdJSd9dodtk9HdUrsRdFzekhlJn
jz+cMx6YDo8CCp50vJFPjQyDJo1IkqU6Kwe667H2pWa7m5VmVuV2FbQm1/n/6z8z
fWv56ciLm2hLbIeYOpR6I4xy9tbz8PYHzGZ+mmqIDvO1xttdj6Ur0iw0RRyMyCVl
/ZF2aWwKMstQpuJb3BWTdbZAa4N3zSYaSU4eeHzcvbXZKkM0pJWGuyZvWrIHyvhd
Rn3AApAdThLz33dm1o8TtF16/5brK0d9EVSUUIwJjCUXpWPO5Wyj2ckgvw9XdhRQ
Jmw8jskhzXCSWyWbltq+ABvVPZZMI6WPguj8D2tEst0WTa1HyFgL6B+SPic/btke
JbxX0AJD6yt5BQHxxl1D68oV0pIYBbiLnJ3eDeovNtotk1Yh25Q65RyPgUcnx5u7
H+rIzZ/k36DKlP1GXpqf9tBs6Qtb2n7P+DZ36V5ql59lkxauXB/TeM81v1yabby8
nsgO91AAfuAF5cRdSxSiKrHfKnhDRHIaz7rk7gi38WM3u8xGwD9Oc1kTaJ/ICJQO
92Vs/qLp9zc3ywD9oSmp1jPFYYJRlswbcqojJeTffWm9E5Rhh7rmRdFOdufvRshj
HHAV3/Tu1vPkTnDe3Vbm7CtaametyGBq5UO81Q5n7ksdYpujz7/zHUwMzgSL/kPV
mnvqZGvMjmZPPyGker0e9ww7SBe8tVwTWYvrBZX4FstEeVJhc1XPxxjpu4REm1dh
68NCkeqOGeSli0BfO43VEC2N9Wx89LFg96Ml2Q+Sq0XUnNNYxInkdLlV5fjQ2dXN
1bIAt9PrpQKdFPL/gX5mMd/pYwgYupDQmLoi34rhX8WAJGFck4+8W8H6GerUJnFi
CjKZUKQeFemuRWOxQDo6DjPM9gYtC5G7NwbT3+x9NRbo2KkaFzKLmsjhYGmgkn9D
INi6y4T1wp+rnnRv6F4ZUWedWxdgPJj3mUgSQJxAnUk3/ctlcgO6M52YzaF4E5rR
KysMz0ADoJpvRU+ABtbE1qo+fznXXrUtFs4azxUGQ+NcPRRQ5HUxhOvX4v1QRclg
rQhZwbGqF8HtX58jKo/j8BryQHhWeGkNxK1TLGpvIp6jKRXOXPV0ovMQ12EPUPrh
RIeILlGQmACr94PXb3R8pBMScif7Yuss7yKcrBbn8DAzRAeuyFV003hHyR/yeDx2
2E5T8ZGh8XvN8oRAAJBIlxLPLGjAtOXIuhSKCuYVFfwBRd3diBjrsiR55kR0i5CN
v/eMrosK+GMutk13Ki/pBKD0wgD5Bmli1/+H6/nwpMn8issm3Ao/Z6aZLzMBQBZ/
Xzlc71Nr7uyLmeHsOWRYg8K55UkB5eoQVx8UW929FaTxOasUzYmnIPwV6Kq4W4ZW
Py1l/6vpCzreevurhztQN5+ojQ72j60jdSG9XrsgmWBuiTwT90h2D/cyJ5pHGukp
juxV9redDXq690Ocb+C0nFkBLv1ahzgx8Agrqx1XHjAsNyBRWi41rLRi90aMqLcW
kQ3/tGmc5Zir0b9ckfHyS+P2vHeZ1B6BP+SWLT0tpt6yfJ11RZ8V5s4wNKGHgjbm
UfS4ojqiBj/j0lagDJSUPyxgQ0sObDYg2jsRF3QfSdQjeUefSSTcV9/nLifgc82k
bsuV28I2PIdHYyiOr9nRdOHchMNU67CKbnECFp7qHzCxHShAQfONWCxIwcq2ohBN
yvxpTA5RbB9t6SnP8fdbgANIjJJDw46Ei0ZnhRXDE7chp0rZjGu5Rd1J8WyNQqbY
X+QMjD7nN7UQYqt2daVOqw/7yy2tXUqDAICIZuwgT/hSQLeMIaqvCzxCcHCB0cLt
bOKguZxDcFuLUrev0tqMltm+9rZFiVPgcRDQEwq419WGjbfkyi5ipblaDPBcAT8y
7dxics098CqM/I2ZovhNBuCJJ+LFHXmfzMJTmD4etiCV8ODF9DghJ9w8QaDMj/jg
4DPHCbdfKDvoTOF7z2YF3hXXKMSyQGSYiuukMJQsoaeGY7j4x4sbHcmWWZicOLoY
sXEi1SYPiqB+v9w9tgyDDJHWtbmX7EwdMFAfg/B+3O0JElEKshTTo9nsou5hML8J
L1RIYc4gOQ5PceNjeScsKpl/j/fVDornL2Fow/CCbtQ3R8x+3tv9+AqUSwSTrQaW
OkR6rJIgQAPOiC4Pgpu+m5PKbw7AIy78ff35hLkDwlhBjuXuqxwMzFrWcBAyQGAd
7dmQ5eY+feEEDhd7zH57LiN3V7qA1Jf8OqDxBwTu3E5QndzzGBuToavN5QGea+HH
JZzsyYnBaA7yQ4QaqV5YJJaQWgSTcjlD38I/S2EwOlZKgItTuwJGcZrhhx0E6D0F
Fh9xc2RuKqGY+B9hi3phbdDQzVZmrPpOOG66MvpEiLVYlBmyuTgt55cXlx4hrVF2
cGPZC/+BvLDlrgUfG9PSzUrhMD8t0O8ikyqDrqcbF+k3JW3NvWfPTRD1bVIHWosb
Qqyy3yL3hKDPyReCwwyxR7nJk8tf+vlCWbbpEWU1F8hi7d7GwBSJva+qkzpQ9MoX
f5eQFJLRv+FhZNjonLYMU+/YFHlDKVqTRLU5ZV+9G/S9619aCME14x3f2zrWF4fr
4BCwf6dBECQ56sF/3yuOW408nyK50rv2HaeyX6FWp99DHMYtYZeiR/VvTAGt8M1h
bp4WSUGbQ3s4/1qVwW3TGbDiIyHQ9Z4Urb1qAaxuQDllaMMMkh9Tt++eM6ECWmBj
xXrJrgbBQwLW2fTq7R0MHmGErPbt4tAiKhFPHDoIGQhfnlnKyjPLACAyDE/oI0/f
sejVuEk4Ec/MzK4bI2DB/N6HF//PTOgnQsYXrKL6NE3o4Oyiio8rd+FSm8hHid2Q
Qr9hqF/PXyeHC9Urm9HCLBtkUXzcH4pkuJMbs3WoMOsbeUF1eKLWF7i0PAXKKAsz
qpXvVpMCPXB/65hGVs+hqE6XUX68Bs6/HLvf1Scacwy1RmXcfi6z2J3tzZx0U+iN
cV4noQQZYKNBxL/WGuUf8dRJN3du57sM9LLC4tgNwcmFwJ47e6dEXT07hIrCEaXj
BHcye8YEBcqwRJ5PTmXORoUbaZv+ixyz5b+vDUwfJhEPffvSCaRzJHto4FahztQc
TWQhtFbbsskoxaPs10MEnwTw0XM1VEdNlgL5e/LmNkCfs5/esSWQi8ppIja4rodl
MaHJKM9NztzR178Di7+e3fIHYMx4YPeArXhOpByCsr/niyS1FZmM33M6Bg2tezzL
X+AZq/bRWTcttVtVE9cOhafkkhDR147qWvWbg+KDoNpA8e9npWyBqKLIpwCaB2EU
mIE9N3yXBCHrv+3LN+thL6EegmTNtCTe+vc8o+9zpn1NtMsPy/DLDCzJ7moIC7rV
kuF6u/SlhlpqDL4FCMpVbtV+GRPO6xxiNIvPEIIET5a50AR31wU8n2zz9vCxCM3A
afV0c0wC5HSeSBdFiTuiXUqcx/jKlCcPBHkS1rT2WYB0gd9jGaq2CE5DHLVBz5SX
K4gzkE9pDnJjjXrvXQKc5dGJugOq3nKaE/MgEMghC86Kat9ZrpRZftPb72RG9e1b
9B70eDUaqiCJJHJyjB9eyyQDGjQIuby+RNG+H4oOtVeWOQEBrAnc+9XP68wzB41m
Y5+C67Btvx6PkOvm/4woJmck8NB0enWS1dPm44YC/xnhl3508wi4U+RW4TiLAsiC
s8brsKQTLbtQTYGeq6X3x7/ONz6+KMImLZJdZaiQgh+NwVr3RzUtREKui0Imgkq3
inPSy1ZRBKmpy5JDZwgmhgrt4YvE4bkDCQgpFdMKGaT+8KY9vpd8gt3PNPfNfAHd
/ksPUVu/tCki3mKfS4CdAheJQ1j8pP35skcGrQX1k2m1gG4jf1K0GSUo/AveQqPV
/RF3XsODDAeaskgDB2yFGHlF38PR2asd5Hr4yajFGvVeWIhG0VvzoCFvnX+fnknN
kof9PaAvj2LRRcuMpGIMPoALQs8Ck2BLgw7DjMnzTgvrL/g0JuU8hkyNOl9wLNUB
hZI7wXTmPcAu2KV7fnCluFlgZHUyoX+sxqJChAWgmfA7lSldIOmaOyLPITkl2DGk
Vh5xXuU8svtSUK4ceoPX2TsBCG1AiYeNxdcQf4t4h/jqcCoF7iGDlVB1p6b7WnfV
jhNJpuR/1oZbJ4MGTUmATofuvK6tpKF0ajqBhG76DRyboZrUx0aMqEhbqwBEQ9H+
Cep/8syOQNQby+PJyiTUIHYGu2IG4GW61cpDYbQO2tz83/lRzQ9sSvGIwpCsrCa4
CHNFnqIC+PncZe7YQUP0A43dQ2SkFRPnSZapG/lzMRLKNNZO1Oh9Wr7WlNp3HngT
XqjitMk4B9vFDlDufzFDEA8YwrWUDt4/tfGfiNTGWD4DqBESjxafAcqjg7ioL38a
2hdgff/UiQ6Alcm0+xUMIHkhjoL06IVKk6VdxsCYQ99Opv6EB5q5J0ryEZxqA+dZ
HO2H0jo3WqloEzk1iVupzwUIpjh4PzMTQ4xjmPgCATOrFIfpzvnGzKPdSdTqcKxh
iJC0Wh+joFrpbHv7pWTBBnvBo2dp1MK05+oiWXm+5Q8=

`pragma protect end_protected
