// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Hf5pHGpsA+YoEIzPCmWme9A2eLbXNUPZOmvdX5Asx6Pp/RBSP0Iejj9CPyYt7BMBhHxTyD0tchof
oSBes1DeUi9j6djnZgOxcgAWjGNuBQhin04VaQu2hXTsuPRmgh2zAQI3BqQxij4s6HE3mVxL68VU
aMH4CJjwwK0KTlLg7EUKkN5Nm33pOzwrZjFSUtr+B4kq6xkNEaBDtKuaOzNF9Gi+TLkecNOwLatG
LQkA8KOtWGh32UpZV5txqRT/NO+EhBhZw8I4yh0wiPNnSchOd8FQSonh+9DRbyOgDJThOXAPho25
FeVfhwmLaR2ULhFEvi/5At7ATnNrQKtP2SR1HA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 15472)
oANtDCtmJry/uablZfDNhmWx6+oT7tYhFBzIWGBzER8HTFO9I+vUiLLmd/moxLHOUiXRDgzaj0JJ
DEuRLzTi3NN6uAUxUVmoSRHK1Lal+X7AWspacafEuA45bU9tdPRfPU/t4WkzalNla4YUwSOGs1Ib
BUi+XuTdAx68/829J5KYq4XJ6zlSbMwXRLBCuoM6e9E8BG0GE2wS/Zs9ADqgkvf0HCqBRmq9d7dS
PWoQO8sz0ZQe4w16l4qFMmgOLMCwGNS9kl/dxuZMWcumMIPeuZ5e+9g1TA6IewPuf+8Jp7LG04FR
q12erzCCsVD+0X4pe9mZnopyw8axOGxi3Wa2HfywLG/xp3s6hJiBrCC7KSVl50Qd3f+wynKZjOuU
AVr/Ki3xNd+3cisYV7T77yszu9OB06xmVkWbmI8hJhJR+wBHb3BmKJvTAIeCeQlNso+pCWy7Y+A4
oTIMCBDgo5aBkO2j3xByQ+04esH6kSstgFSi6N9IB4nNDfEQWAZjDthINTTtspDKVUJml7O8/P1i
KqArddN/wk4Gz+6XGEYOFXClP/0CJ5ShwMYRudaP5phy4goLnGS3w/ya9pwIb0DviFse0pQXf+v6
xnHP4ZVDzn0sok5EG6VcKR3Y6gz+H7dH+4AZdQTkObuvzZnIsiqSeTqKq5tSG+GGDtUhGxzQ4xCN
sUmHHrCTy0o7qVAwxvKdWZwzzjTiJn3ER34dUsrf/aN0aytFAQI41eFXZdtryIxwRN6oG9yygbIr
+dvOW2wiNKzLm9lt2o7cjVb6wJ5nQxiJEzplY6W98x6izBWGLCWWtP6syT6z0SsLXj1wtNPM4ji3
VZjHOezvaRuwLtrRUOLlwoUHccgGxTTmR42+YpknoD6cnkgVu1PHnbIkXQN1fLe4WbOey3uakN1a
rk0MyC3JfHL6o/WAUwnjRoBfQv9hXtFnAIDuQA1PwDFhOYmhLPHrHTg1uV1DpYvurpZ8AG0rZWT/
uFz9kU2pInLcBictSnM2oVBKs1EBQXMBH/uad6LWele93pBPyi1ncsD/ap8VhcBOEBO5Ntcvbx+8
64LTG8O/bdtom+JGKvi31TaSO3DXVYuuaeNHAsobGeyEU0wFLDm48uGEtpX5XJAnlvGkc0OhSqMu
6z8glmpx1+UsEbmF/xYuo/CEY78C8kS0QL6ku1uTG8h++tS4ZiAQ3o2dK9XhIzn4P0dYnWY9GW27
l9iYUTD2PzFwf2Jl7q1vR+PR3lKLaWLWwPOYLK/VNG1h+DkecZALJQWcLfW1NXXOxbKvLSz5jv6x
fBJn8N+CBEjBFL5a7s3n8RbS2WFaetvhnbAIq3uUm8jYPHOOedfBgAGso8JCVXcDKCsXAMIR3Bnw
/R5rl2aCEnyQR84rGeyB8LDid8nC8T94MWdsLvN1NbQrLnewieBIRxIi5eiEPXxD4Oho0Atx/pcs
HZRUijbLlk3GwUQrTIOceQ7Claia4phLbZPFldtaaGpqRAEGjB8BAN6gkvjI241+1y0k8XuVT0Yt
bwDQF64rIYLY/tPDzcikpZkouT7zDR+jYUBCSp0h9pfQDoxvH1WOStVi09mSmyKnUiK5PPpOYtzz
E7NI99F7ZVkh2Uys/YQodUk+shSSGuBR1a9nnBinrSaMwneuuhHy2+EpzvuyZPmQ+++Mk+9ycAc7
au1d75409u+Kf0QE9cmXHVLFaTAnCAH2d4AljcW5apr2w7pj1u1h7ibaclmlKTx/p3CHZqo+Mvph
xL7FvxZSku4222+y/R1FDugGg/nnUDIvIJFaj9DTQ4YDXygjy4ui0FdsnFYECfZqt2U78L8Ti7ZY
DahZAFgMrROu31ovNyls9M+8D2J0wtvas6qLg5b2t03L0fbYb+VTNv/Qb0rwF0G5uQ/egMhUCfg1
XBy4e9Tl+3dvJNb2tSiya8BklOG86CyzB7a6t6FMIXrPsJ/H3JyfCISLpXyjlZMAQAQvRLfctBwh
fE6Fhaqf6FTHhnZ5K8WIXPZ6YZlzCwkI1wsffxMgqTLaqpW5REqjxEtzvCJo+Af5chDaP+n1PaR/
zBDdVlgkmM/am7V85/iz2nm9nMDaTbxQx/qK0wdZwffltyKUGUmOcZ3J5A9YzSJ3zwkCQueTtSoT
x3Kn1RWriWuACiqTi5W6O93ZSt1XJiprvkvyFN5yy+BcRiJyh2khVy2OF0aHpXsyb3Cl4OV8MoMg
S/NEZRs9HEZ/3L6zoLwKQGpsWyXp7pfO8mTqgmskdtyZhCrbLK+wbwvcF2ve5e8v/1sjhg105Bxu
H6KpwYbksi2Iz+6A7cPwhKVl/RiIXmGh+ACdij31KKOJdz8spJmFEcJq/JmcaVvv5tZ2Yc8ek8cp
XieZ116vNgMz7LK1SCS6PC17Z93Wg7/MG5e0+X6vr1igBNn7ze/4rgC9SvKWWcMmGWsx1v6sfyXp
DUFViFoEAgHRp2VaUJyurbXSZItR7LIY3S9d+ad3S6N3xfajp0d68PIMGjZUhXRLIrFjckQSoL1o
CvCZrm2izd6RgLAO/qBSISfEG+/o2+cFtmK31vIBN/E6pXYzTRiAhVFJVObJw2Uca1LbDv9moQ+R
KeC2t+jaMiBRMUMYQFRDyPSuxczoywF3Y7/rOFW+JrfAvCG9J5cRtIjW9vikSJAShc+YwHgJmHQP
efVWL3MMbpKyFWwCZX3SiloBfmsRFOsmC5yo+ttVB42iQ3Y1YHl304oCWR0d004YyjuDJWSDpJLW
1cNyZrJUyFn4264khxn6dwi44yBdVUYL0M3xL8iU/6O6f5xrEmJj/mUzW2zRxqXuRZEmT15cEAH4
0GWFgttiIOyZWv2Wna3O29YjJ7DaC85scYgzZZhoEDVyWr0hROAIQ7NFhHavGkgXjeCP6nSsVxqt
tPdIWB4l1sVwYyRtuGVWbdpzxFCZs6EOHPlwhBKXsOcu7QS68yLW32TXyZ5LAWiMmRMyLSoqhGvP
cA3vCjrtTeLmZsc8UT5J+P2nQPGYmGWmSxooOmoqXv88dcglHZLpSOme0eRhfmTiAYrlEnayf+vA
ZL4Sn4mljQTh9+EEvspDLXd7blMMceyrgAinY0S+UWbcPjVIeUgR1w6+vPMNHrA5Hpu8BRX0t/iz
eW2zn0n77bpSsg3NLVa9X/1kqNYEh47O5aIRFHUMFsDfc55h1kvI/njzX1nLKgTUxOK1jZ8Zap5L
J9YJLc758Mr3tFqQrmsVih85NrQ6cM0Ccxphd1x48VV9WitbHNjed1ELD1dfWcLez2pLji2UaK4I
AObuohnVoWlCy4nHIpzU/wNGnjlXxbxwn7khcscGXnG1wB6MA+zf5zV1TPyXDSjci7HFIjlJu1Fn
SqQgx3DhqDpCPwavkfyKLdXRMSTY6VrQ4CccpaKtpxvw183zjmu8jxjrRWvf8zT2SDgyMH88qPW0
+I6sW/3MZVbJQLpb3lYJlYmT2mi0ExU2Jl9MCEHP5YQLuJG4M6FptKF659AHLY7cnxF38WLhVtgS
d0IsKI8I+WcmDZrt55uTxVIEl14HBLWrpgu6f+GKwa259hwMuNz9OF6WE0oUDFyBNFXJbUierqCz
9JHn+xpaQeUPWSAwDTk4n7JPpJHF8PKlAN6zG4+9rmccJfaH+wJxsyHThCZh1ELfmY92sHDzhxWB
+jAsKDg8muClQuo0G5i97e6l0KOMq96xyTKEcp//35GIdeochzalWhy6DK5R79Ax8NuXMbI6JJuL
pRv3xl1F/z5dkNgSOo0wk26CzLFSAdfLNIOeSFc3c7gMMDqxFEt8RGFZEblhOQNMGemVIvzW7h3b
DB8cCPeRWyjsmsaC7CYDfGEv4byTotXK3pBAynEm8xHJnBGxTYf4RLEb3mdsLGjXeS8awFC5JdUT
gLsmysmtGpoHCkBzRt5euxoFjOP9p2x5Eh2BhzvBgpojIF5Dw7P96PqFfdse3j800dX6By1k0/6i
RBukwRzW7C6ZNjwcsdry0br8iid+KAvYwoPIHU/qgBuD5JBmVO166mF8NTafTQY2AtKxN8HXSPHn
gsIXzpE6VbtNktAGribA6yIemVpBGpczi+px9gHcmCpKWhxY0HpbLDidt8mV51fkHFrX3bsCV0pv
cjPlsiBpfiIwq+1bOQAe3QZ/HG1ZQkS9Vi21LOdffEG+IX1GtXHw2zLH0NWmWNonOf+awUPP1tyX
6Xjb04lVC7qWdYtOQcE2ZO+SbEvUmYiCpQWvTH/lT9oheAypPhlP6hdPkkxPHUAqht/e9kqiWSlb
8KtDFXpJLhITCHHO7aJ+qF1ieEzeF50tuX5tRtboXYVjxUIMRS7jF6ci0BGnSIAxDfgDn7kWAmom
F4dY9b7FGufnBignKrVswZObCUdMyiZ6HbD4qygrkJAkeMhro3UwLqbA8nogS/cnymM8OADWHMiq
qcE4JyjvSqMp9t3WE0HAgtGl/qRL9cQzUzOM2oUzD0qoZLjMCzonVRi/pHnp/Fbs7pe0yQt2oAH4
lTIhpj2OxAs3rY/0Elfw7R4lEuvQoTHJ/bj8drUrTngPT5Rqczd88r8FvEuGvgZCPgQ2wj3liq0B
TjXN4ED1nLu4E2015XXGc9j+xVMTatmCwhq28SnMqx5JKonFVtIkx02fMYeDMGXZOQkncOIeNW5q
ChOG8vGgOGRrAEtmf3KuaG0/OPhJpIrhjnuHV5T8s8qOwWdh1/zsOmnYtsvT71maMLz6PTOQhccP
YMoC9P1v0no9J7GGfGJM8ImZtn9kUr4Im8aKgUnM7Ful/zuY47eE+ekGy/x8B+uPKUemZFhdApE3
ctdpHB6fIR0HGT5APd/h4etdCqF9FWH9NTBrO0Wn32ugQUdJJI/9fKbho2PrElt3nDIBMPrf/HhE
z8ZhKgTEeX+op8MOV/aAm5MYDlmWsop6stcKas7OiiKdvkTkQsCTYra/K706Q92UTYxfuj/q3GuX
ulbwI8nXXpC6a8eHLF8K5cq0I5OpWOPmAVzHjdkn7S1MMUd93nPNVGz6A0vQfVc5MT9SpHsCCgbZ
zjFgSGubD6iHrlkHlNlJw9SjJUhXXXrgE5xz4md0g1PlTJ5JIkxBva3GxCNStFNR1BVY16ly+sdg
sM4vMG/MxZdRxoxABe0PI7DeVWScfaQ70DUqjU1dkO1VFyuG6sJXUZf/odWb5lwnDf/tYxNncLA4
EwulYIdrYbzCup3SL7HjJuz/UMK8Bvtt7sU2F8AfzMni32eUGytY8bGgFEE4QzyLZoY0VGpySTg5
mIjFR9nPQNBt3QkAGUCqLsPID/bRGoj3qeczNBWvekdM0w8jx+Jp5Uu6GkPnXuC1q2aikURL838P
ZArsdmJwyzhPQDGG9ai2muWEmZosrCgh6ZIsi07GxE4owRrsGsKnpdRPZ0wgAc8eEHgL81Infdm8
mlE8upbvlqC+DiKDy6t4DJDq93H8eEDLkSWBB38vhwmSsWrZ9EplrTWq4fXDaxWp2G/JOBYUvrnc
HLxDnhdv/ImB7Mh/agl2EO+sRiyUhmqSJbtPci3kqwX4zfSnFerBlV90hD9pdxpwJfSfcpvw7WfT
OCzgUd9Bah7KkvKQhtfQQuUfNMScfD5aT6BEHmApZlU3aEHedutQ0pJvrUGmSnXmlWsxk+DgdPMk
4iyGzSDfuhY83ZkQYc/w0yJa6juREdgle7mx8i0q9h1KqEi4xPHJyfJlXgcoMHdU7C82uYe7ouiF
bU62j3Fh/YO6cuANCAxZJ+xILXJiYbc5JilcbxI2ij9jaGgKWkFS0G2QLn5YqptR7mQWFfpt7hKh
OgJhyJvceRPQLw5+6/gvyuX/hIMY37APRU37EE3oEu5I7uRltHsvysCzhaKDuQH4HpO9BbPAtFOU
rk3kaG58rWOiJBsaBvNBxVpJ9rYYo0sD7UTjb6OYv+IdRJ/hykpVYYZAI7lGpMmWbL/lVK65s5oG
xO6sUmIlZqbZHSrnZhWIxeCQiS2nk1T/W2PerIqKInPYtdLgjB5sMZuPC4etNRdf2WwWibCydjV0
5iku+krZh2HBNTTuIi0LTFiIC/a07a3GgEz7PikNm3fsnVLa+CCi5WKBmgi9Al+oF5VqG0C0XYo7
NupagSPgZ2aBvjXqvJN9sVooVlI69N7LMY6pTpBCKYYFWNDnqdwxKt/TmMCmrPKilz5E+FX1RQKA
K0WQO01t938kvox8mM/ZbTe/JXXzspHg6rUoXUW/F1F66WTcUctXi9klQMaexMyJgTwM/pRCqD+s
6Wdi0UAMw04Nl0udMoNmr4B5qtWKKFVmQd89H+A/hMWj2OvfwvH9Eb1bjPRR2KsmyI09ATwmKSsA
UArvXp+SE+VJWAL1lc03kC5cmXvfbeqix6uylIqtpqlRGMazC0shDnRTe5nONzffQfwO+mxnB7MF
Iyhue9VvZlVsfcSKkZF8ER1gMQa9KQ/THwEWfLTekaqge78RpBJWqiSuWZOGTq9ab/15m++b4ZCk
xe3d3ZO08je3SnlJ0pbB/Jpd03rDJbAFmW3puKnPaLMKENejd49HsCaVjh7G0P/N9QiojsVrlQh9
VV/hpXwhoIxTTGBHxa/8H+MbFAM7SfuBr6suM7NFK7aEvuOyDQrb80CD/wRRnLCWTqAOdFCXY8an
1KxWHCIr9f1tAkN2sutg82sjqUYGiW3OS4B/iM5F8rvSUc7X+Z0QTxB5fYu8Ammy+7PTOs4Gu69J
t7KUG/+pTqWwRT0gEIcPols/ubsAlvnUyKgYs4Q2vyt+mDjLyA3EHF0PEUy5YqRhVC71NpI7bHu0
yRXIiiNTJATTtWcJcMBEmCpBg/7vv9F92Pg0CYnxC86RpQ+R/z0IwQvLWmyinqXHoJIMpX2XpUoM
o3yrr9DqiLg58uzYFjXbibRoj7T7xr30YriVN4TSNcXAM/UKa5Nc19Tn0iZHApBCGAUjDpeO/lU7
gQihRUjaWFJcMqxXLsvsud4qsmdfsO+A9vAXxCf9rcj/GUheoLET5NjqgNwGALT+x8WN0kHGZJiD
ftAtrgRRwmewVI8w0Z6g/P7RN3hhEGgO0qhzmn8A4hAN3XtUaIfkCQ06z1r7Yeh7vU3hDAz3OAd4
EiJP5dRKlBbO5iguXO0tF7TpKdOn3CwE41xgIg2/r63XFEb3MwHjmxKMVEelwQz2x+8nB9qrdIyX
Hz53LcmJ1c1DqOg2Kkf0YGljuztkY7ti2W0RnvxCgajPy0Dk8eErgsjz9Kkh0/R+Tx8lf3mNO3iF
xOcDiSwn6C7CuO79z1ojlpZyjtvYSCGMMEuNBjv2S1leZJFaxZ/9oXdQ/BQjKK2QkD8Q3M9Fhc/h
UecQEL38PLK2xurBenyuYjYkiA9os64fZVkb8fp68VdIyUh2D8YIxaz1XHIYll6cZvdDePoed2hN
1IFPpJR0krmpnGVM0hQy8yLfUTOItDcWHoKPHa/PG5EreI1TBRkfKU9CfYtsKVJIHK8CvIP7/2O7
SXIQIZ0LF1TllfwExtrWxqubz5n86U1vpq9WEscQWtOfkagUFp1OL8CR8MZdC0fwh32rRwQXksC/
uQtbtVfrp1qQNpJBRd5bMOuFGjprj4eubkcVnv4KyGyQDiKAUJGOGR7h2FsPR+4mbs/eqjuPG/Fn
xA66EccDsJo2yrSbd2xb5x8NzHUCtZ73znOS12ATq86BHS2AajnVGnyFMbUtzBZRK5OrpNusSW/W
l5WAWJEJhz91aSc8n58IG+4iGlYpfrrhXq7vJfQGgX3xTpQnmQ4bGwBG+puwa8yfFGE3AUZmJbJM
D+XhDHVi7i932fvuG4DNZ2V07TbawtAsOFrHLaPvBJxabxDZ0P8va/HEFlKi//FYG/NpE415HyNO
qbnAElKnvnJPRAKR/4EqPSB6kitx5MGH4EGz2aGyYngc1Cp68igf93aEUvS4GoBqiZT37/H2o+oy
/hFrJer8EmEqLeDkOYJwJc/EeW9jfW1QMVtYNUa8+tcNAG9P9e+qbp+cTn67xfzCjA6H4BNQqSf1
xIcbzkMwz3aQ1ka9keDs/Hie9XOmpdvbYmogbfUB418wv1/xUH6lxYXXTa5Rl4OefeYTw6nWPLpg
3UET4xvbYQCgWuoBs3gAOlBf5Zsl4Z3UDG7WgVY1t6qGC9Tvv478b5ZOhftP3VVvyDQSwvebdq3v
Echo5b7YFI6Hcl9o5fkBRaAlqU8yW4kQdeWi/QDfb81+Ot7wDeObh0M5BzYHKmxbJ3oubeqVFGk7
ewy1Ol8VltrUc3s5r/Kp4FVB5tlaX6fOGT4UbCLmW+EmfzLLhJ4jM4GVxljKOuFGC+DZBwupZ2or
gvJST0eiz32nwYyEwKhf8xZvpmrWiiFbPAAFI5K292vNld8BHccBel5V60vxZ6Cz1Pwf1+e+FG8V
OfyLLA2N+Cp9q+AL6fwtI+zffVT5FsUsA9uDRZgx+o8d/MNG4kRKPGB5DiPCg109olcFc3nT0hyn
sf5g4TvHMwXPYl4U8EdknQl6OMoLdrBuNINmX17gMvTKhqAPwZwgm5hGniowDE/z42V3A7yNoWPj
D3VX1p2KUeJIUTJkbGAkoEPIAMSJlvYUjqYDGW1QKUNPDtzEHHUx+S4i5ji/LLN2YQo8QOA2lGYO
9a2SJXt3/Smrq6SoKo72aPxX5SqNIiWZKUAUKjXAni81ZKzcWM6rosjIBTKFmnceCNNA319qQUI9
2CYCWhKB8t0ior0/NiC67rWTDByBTTlstaAo4VYC+3t8LdE1BGh24TRhRjFWcc8lPjk7GzA/SH57
I6KpBIU+s8wyX0ly0EbZDLp2VcKYItjCGzxDJR9C6Q+Fvw02skXmnjtLa5qxUdSprwlo4bvZVj2t
nKvdwupsqyiLYKG5fTgtDCvPmHptLhMlgMZU+Opj+B+s/GlGB64redPx6Q2zwJVoR3dmPx2l+eNU
NvKyajSaLI4RzYk6GYOhDLoMaS48Byh0T7TWgAw538wElLnO/7nqVt6ON8ydU3V/Q8aMNGhAB6Lx
pbK1KzRIDGBBWiqDvF5oZ/6uxdU1DbMtd3rrsjwdbWDmHK4Ys6ZcZqEofJiyt3fwZE2hRmEIFc0w
GHTrW4aPxUNjFCZWtemqtXp5sFrvhTmZG2JfNPzfITHitNbFIba799hmoKg4oKW0FXcpye/bEg0J
wlii1DgNrh8DFsUrdnzzyqDamS0Z7NKO3fAux9QS24yKA/4LGLDb9udD2bJPlQvQJHcnMYTbX16I
bwLeCGrDeVPUOU4yxYmjARD/A8L4rCH+iuj0AhKcSjiSVWouKIVkGK4fDP4mFJ8Pop52Hsh+Hvxu
+Hmsy6OwSMHsHoc6IE7WU+/ZNftIYkL/nYRL5B4gJkJedHDaUIDj2nI9I9413zHhLc8AlEYWWr2Z
MK+tbWGUpwxXN0S3g37uiF8+vAzWrJbKhcgZlCMqXjLQmRlvwK8A6d83ZNeVOXFcfzKkwFiym+NO
8xV9tJIlDKoIP+NgwvPdx8oKByVkrQAfXIH9WRVe6xJ6FZuBm+OVoRsDrZSYbaH8o3n2oY4mthx+
zz1WFbqAS4Tl1zEN91pT3JlkItuYWkXwMLOF0A9rRMYfhn5ZdiHGu8lYlcSvkK0ZTTL8EHMR77cU
R5dPSla3ClJUrc4Gk04HxohFrZu0O+bTnZVyUM0O5hC5v7vYs8nNGVkvf9xYeSDCTCjbpvzEDycD
4YPOsO9hNwUz5g26nS2N+/LkxA3Wzw5wC4QYk4JHsjIztnrVHEKr8gs9vmY3rag72iJsU3MLu/Vv
sS3/9hI42whljv5mTixdiQrZgHuU9lI7NiGGJDxKtgfyoQavCv3p2qjLeLkJ/SWpW1B+eQ1RYLWg
QuZ0maNiKgYpe7Dy9uuK90tl4zA5HyUBk9sAbJb8AyxAgqEUQnzYDwMSTpGso5YJ2L/l6/Hee/xY
RKjji3q5ARTez+D9jAcUEvxywmNkVvnfN/EwysPwUSb4j3YcVqNuWUOsjXSSNEBqxO0bXj9frao9
Q04jfM7d/dcSl6tAp6NaLgGaEFrqKTu8vSQLz1xkIFdqes2ksJ3ZS/GfU8fZq1SgRrMKL4qUo6/e
JWZpuCKtyjp2KIpU4hoKZhfbDa/TI3He1eFQA9sPlLdPQM7CMHY4iP88OSNsMJojdOQOS7DJIBxm
fIZDox8lNzrbnuUhrxUf6qXqnHmht83p+OXKxVmMMgFJTcQ8OQVE+r00180jhUBuZCIEWTj6SMRD
OUoUzQNAmKdPVrOaSICLTRdZMIo5K1UuQcDQRgcD6qzJAWg0czEqNRyEnWGOh3XDa+5dPdrcP5K4
1TiZk5X9BOHrA7quSaOnHgOrnxXPnxvyD27HBexPgCydD5+22xxCa1L5ugYSvSwms/EirHIuJ+bY
PM8LFyqwZV4R70xfDSzuKGQ4+dS2YVGQWLNizc5zdH0PKAxuqbVrwSor/mtDcT5636thZkEM0Dxm
dvygF3mICM132WfXieQ40DmUhm8y5vuWAFqKKt0ri/qSfqVbP16K6rfTVQd6EdLuTCG553e2nztm
anTND6HHfa9W4vjdz9q7tpfJFbfrLhvxHirmuYwzAZho4wkK89kDc5GD5RHruCPTLwp0V/2p+fJw
T8ag2EXwzwRPqT+QAO5AW5hpUwCgFnqx6rMLxxJ82iXdvEvWlQtaovWMLaIm3dalfE6Cc3Ge/rgy
Gpw6hDp6TZoCd4+17yA9ntdJ5nuP27hApnv9mZBTvy+puwTSE+L3IvyqDAip1jYZ1YsKr+1DM+5H
5MHUdGcbSMQDMuiWg85ABTfCAvXGSCYtMZQvc+a4Z5fkus55OEJtUaZmpFS308zTMXam5ekV0Jsc
tUQUIbftS3367Dbqmy5W20GQWJr5f3DKGID/+DNIcBxh3WdkQmvlK7srU/HFsfCjxncGzSwG8uRt
Ke2zr3eD9dK3O+zPZ7zQ7tQi5UNVQbqo2znupFYPS+Jj6mi8Es0wrRgmxoe86jIDPWT/RzfMMKve
Y3TuL3+kAV3ZOPC0cJdou7n/WSJpoQNpcbXp/6PytK6bSLpg4af6NDEYXFFgXia+opoxJWXP2EXY
qHl7wv5KmznH4N2Umttjgr7T4TJiVnQNPpRw8vxqbXQAs7gd4vDYpmUyZ2K+XQYn4K6qmnX54yZU
/lSq2BurnsgmezMp+SbbgUfFx5TRBgK1Hwkza/fnWv9eY0POOlk9MdJPjZ+6uYIqQt1PrKcH7Vkh
9D/+m0KmrU2lJcHnuyi4BCYSbGo9JybjWrfcor1jHNkCW1hZa9tYInjLBVMFvSuMzupHjTuPGbV0
LS2VH/JqYqS5ipyTfx87H8G7ZJ3ZUh6kRQlpGeY0NO3WuFFrcL6UcBEMOpm5jKv1XKBofaUiszvb
gh+YsRlQ+vxCqUXFaaqjNRxL89tZfYVJpdXt/bI507BZ5H97WjhPFZoUP9KP7iGrhlim+mz6sBK2
x/hSKHdeb0Rm4yepT5zlceOyOlOKuqAx4z4dQjNVZycBVYaP7YXOhZbf0Gx6gcklJi+SZecMp6x4
pYp5xxx8n0zaDW4ahvRwispi1uWZ4crXih7SQYheEBobqvdi4sWu9SCgXalHz3j0mbm6dDcICvgV
Kdy+lanhuFcRFTtVrClryer5dcdYLjnK9VMh+qFKaEdFSpko95+b/ZAUb/eNZ6j0neE8h9IVDj1T
I5gTSmLIvZbVRsii96bHMi3y3F4yD00S0h69Coh/oCHFsDp67gMJrKpwtw1vh2cUH9oh3N4Yk1DM
mLuFNDk3G51nfyqOQ4minUfEEeHnvp1PMeY5k7lhVLM2jlXCFwpEcIY//409Sd2nE5391KpHNCYn
CHR9kEFN29v+6r+/iS7YGGJk0P2C5nd+fu4yRrmMy8sDQo4vC018Lncf/uU6LROV/7f184BO4+TY
20/jAfX68g42S6nxF822WSQ2fhpCJuydTLg9K6icc8MxNblh9i0xJmgQT3yu+NLfiPDrjJP/IlO2
NXxlBbh95YNa7JOaBwdk1ofCgVESWSCylI9mJcaJd0M9wrbeYO7DI2eGBlC/bQLKKB3bdpZ1uIHh
s95WqzE5EUBbrwWeyYMnalOgfIFnbvxLju5vC3kKrQaQo13s8hohCdTVz9vDVGZnan/w2dJMOQ1f
579XmUBuVp9D0Oe+UNydJFV1wBSQZki5n2odYOsbgoyN6HrK6bK5I304ufdAR7S/LMaW+kADRF/o
Uw13YM5IL/HowCkPX14nHVOJVqmlUQjFDwYz0arsWtUDDY0iDYP7b53J5Isxe9Jgm16Hvcih8tZM
XBpOciDvbUEL1jYYJ8PnhtkPy8si7zQZZr1YXQExA9vYV1eKzGJXL7qppaxybmkfGR2jPYbl5Shp
t2Ces1vbSO6S/Bs3WZWF0lKizmMfGDFDeNXS2JGth8yMlFCHSrPIp5hXjoF8BoiVcBXQu82YNO/n
snR3PsFN+c5gS/ZxjDEmETAQQDIHKl9c4fwL+a7lR4fV4VfuEHwdNmKKStZCVWXXYR4v9rsycZ7h
8jaW5NrGGG28DM+llliAFimHRjO01/WHHji/w0N2SYOyNA3uDH7g2D8/egjC4UgDCgEJUCSbje3F
7IGQueqyMxWzCd4rMhagiTfh5Mcs8HLdwgikmHN2QqaDA/ekCP4OHQaEqmNUGNDQwNWt909gdNgu
7giS6MJSJXirC+9T1+DtSWPApEgJWJIYd2w3CYUjcIgg5WLFAAgMrlh83ElAGrfKGBIHOKSCKv5A
2WHxScXonjzEnO7FbvFA3wlMSJ0oqOLbF5eacHbqXvlC1Y9BxO+nmXhr+voEEJFQe8vN8/E2yKIg
PqhMDSmxth0wI6FGmX8bEqKksAjuGHhdtIGghJol6qn3OhbTpcaPz7TA4iup7EKhlBeg0mp74ksT
CwmhbIf5tTcYu2pkX/TcYA/tQrPEBDo4Xla9E6Se1O69miym7rk1p2qmAg3gbxhWXyTOBJmvxKjy
vQynmCwQWEMWlaFb83hzSEgITcgZoNal3PCUkuc2jRASL3MdoOxPzZrKn0Mqvxc3WZXbF+kw0b21
j/V1yzC8m/g4aTPyakkmsEmzWeH+ZGQgf8/ggyxFuhDpXnLTDAKxQXMfHhabxR5oaeNjtSrtR9qI
at/ejoVfFdndAz0/0QOzLn0XQffbkBfBdzOoJ6QYctCNljhrFa8W7guP3+4hh6dQVp0pSLRhIr6F
p45TKmLq/GEzExeO6ZZUDnm7k88ZVfk58uW5ON+I9nVfEbMiSbxL6B7yUqGVFZ9Bs0DC4MJtr7pb
Wh/f6jbqb4XV5g2uMghGr32PTY0SiTurgCdkrFbh/pICIdrb61aQsn/5r7o+Ndq4MmZmxoKWjfIA
GzX4aXpOukgbTueIVtc+yxChkcfO8y8E+FVo7NUK3uGY1FQF4JEQWPeTzNCFM8ZxUm99hob0zS9Z
xI16BVJLlkdNObg0SBx2+Z6WX9PqW5J5fzoXMEQ7Rzn0FuOlCjrIYpK9Dwk8SNyzjz5V4wLC1giD
e9FQjOvnDCER6adh2oG+TEmabFWkDPgA0GBaW1MFsoUgnMKr7KhMSsscNT6obi+lhHu91ylcquYt
by16s3UzU+a1cCud0nHXSNqCtj1Y0jwss19dThdxF1q79S0dBVwRuWk8V3gk35pnqZT139glWmeo
/RmrAlKDWsWtwSmOpic7HfUCWp/+3NqEqluUY8zbG3NPCOIbMY8hOKCzwxBn8Z1DJkdrFoUsqO2Z
2a8RIeXDpHef9O7jByUDwukVSy6TQ6Tfshvy2ZxSvA5//OkLTAm6/jLLF6uxncwapAlHt0NobqwM
DwxLUentzdG3/zp3A0S/f/ICMfnoX9TqXnV4u4gkPksy4YeXIWr3awvUWfDs03oQmgzSAb4HCcJg
Qf656kcVmckXdLmJJ8kHAHPfz6TGIQ57/wjt9O1CWL4ayy1shIv6wkUtDN5ThIh6hA07G6pZL2zY
BKe85oWItgHgmBB9LObDCvonOmvLB+bpcY0k4O5L3pDfTW+Hd5ybVP6uw/hKaQKlfqz+V9Xh3Qnf
+VmkPtATRX7XBK703X/10lR+4HAXs5jSPWd3eYdT5bCDVi1KzC+h2Q5mUtcVoKXZzcakw4Gq+obx
tpiuRsLt5y9jjAZGR1gWfFftaNfxqz5oWy0nNjW9lRSu/z/oRp7KxybskqFZGlC1Rmwt3QRytPyp
ORiMuDNAe+Y0hoCa/eY7nidBppfprf6nVh1M8wyOigjSn+P1Wsaaglq6Z2LYu/JfcZdVZ2+9Ykm9
nznZ9deLxtYKmPQKiMRF2JUuVUQWQZ25tF/V9SiGdGXBJ1KxN+x4ssz8T2J3zKr6/01OBVkiOaCs
KJYYF4sFD9Pxw6b2fGbi4899sz2DDs8I/3RVGx50p/3Rr21U1XZCHgJ+B5sp+cIoG/NfSl5jCMNQ
tUFZaXTS80We30uMwJ1RdKRVhk9+I0Ht+6dUkEw7TzKe0u+uuqc2NaXI0GPqrwrveayv0zhvLWTM
L8jshvDQxch5iI//Oes/7ipHd4juCdtNO/cUc47SDdFP1QZPqnMQRdpETLQLMhy8VIXhRiv6TG44
YO19v4Mn4TBD9eEvwaoDjzu5ZDIM/D9uo5aYgXaJp9VkH+I3CTLbqn2VQbSsz8Q5PfOB/MG0hV+y
nb2ZgYtTM+tjkXFt1oGPJqexT37GmaRi7amQDhMXaj2d5i+ewOR0vGv5hqEEcRI2phLxPsMyFuzn
kTIdlL3B1H4MPfiQl74vXW2ejPlomkLINg9IO2IjpwUI2mythK/ejNCW1dTHk9xlL2cpfGqsRCUF
N7ElooUUjOLTF+RLX7shVsDr5a6zqVfXDBS0yZnIG3wQKM06uxHpU1s845LxaOMe/DlyKhm3nfgy
RdzjodBF2i2JqT7itMbFMhXjA5frmuOSPo71vSNRqtSZ5wNp8pXse+NNzp+sKxbhIow90mInSQnZ
jM3e+KZRy0/k9G6eHtDd878flTh4wQfvqMoGwqjz9NyLmWA2VB8UAbYVkI2xAddtXm/8OYzIaNED
K+G3113tDeMpiAyua9TvhnU3fJbE+LEFJBtgrLp5e0ytZF8DCA4cnRzJZ3Pot5tVMvaqixFFufE6
vrxwX8uqukiJL1t67NvfjXzlxpkpNgD5qtfwo6JLrb0Nku+7/m2vNPzN1GNC/RZXo5laLCK4p0QS
7Os0o4s2Yij1OzL5Whq02uHWNvRGzX1QS/sESiMa8Nlv+NRTAwP4oTAVHhaMLbtoTdrHAyt4YmVH
pUtDswDMm1zVIdG2IOc1T46Y1Zjo+AjCdKjSw12vZD9DCqUifOBwTR8xRwbGUhn9HAxEyrbHWGRl
DN/BPcjZ0BsoGxakzi2lIlKeF/4zaaC6BF9qi5kvdQ1hgvonEYDXB8HabD1fHlVzQPFgCWP/wZIB
mnALF4wQedybsWBP+MrTUyHwGCGsL2NIxo6BeSkv0Os7Yj6m3aHreUF4KhZTbK8a04qOuhfQfX7D
T4I205eUzKGuFTejcZTx4sXnlbfwVoeLD74BvUOesXdAQ/dSRsdSED+hgPoIAfA75UBOLXD+/tm5
JC845NEk4ze/OIWyUEEwbfVhZ9t8czYeBZJ5yjDAYWi08TYNaHbjUrtk+FHI34izNH2zL2Z+Pjdj
6lZJUvJVZcUQEuPnjgf60q6KV8qN/OzHL8z+XM4rV6fakZQrzhL0k8S7TWFST2cdsQkBYLMkmLOf
P6Pv1567CyIVw7DLbzyS5B19nCHTT7iE3aACNVYM3f8xsuf+zple4gZ9H96XG+c3/zu3hHY9W3t6
trfM6bdI0MOTYnmBJWwaZlCWkZabynIQTKEXTChZ0VcSttHXbOz2Qavz3zH/36tKQ1TQhDeT689W
5hg4bfhg4pFU0IUwKpiIHNyZA+ZIdveTQdw5m1S1xm0/2m2SoV7n39vqRhx2OyEmKuJd5oc1lzxh
R2gyadxo5oN4yfVvduPG/HuiW8kSyZgt2wDo5RvhgE7++KRKDZE24dXz/jOCXB2SLqT+1PNhLrxq
3MpndZqTiAtjMhmJxqYDx6r+jnWIU0uqw2WdmuKVGbO7AfmL0Y+R0Fcdc7nxwjVkwhl9svOSl6bH
Bh77Brl8j1Zq+qZfjTk4LnYBkBtgE7W6nHywZQxTeervfLl8GpL5lWmwrmgWM2btUQVCw3vv0zbO
Y41JDCr+fWYYac4LoEGUfDen8Qww2WaZuAlN+83vHl1olLJQSgJ/bghqGBEA/puxXbBYq0orHRfg
alr2N9UeJHlK9n3ZEDeaQA/YOIAxS/dWrL0FnnixOZ6oZ6bGkUKNUoJrgjVWzxm+PVP/vM+IzKtA
7J7jIiSqmPoGJQytaXYTSV8YyalY2LEbAL1GIg1L62YIFhLYWLkejcDJgwT5EaXw/R/LaNcteqhm
bRC3pdDk55t9lYY7ybJO5N2S/znQOT4RCbZSR0apr5i7b5uF1i1cJi/JUC2w6KRPJkHpgSsWiPOo
7FDUpaPvh/33ZP8XlxmziMM+y7gEkTDXwT6tBCBHWDfe80JyOKorq30V00b4cJolx6rJfO++2Pim
PnfJvUsbixCbM8CbDd35M58RkQv8go2MrIZZcV+2jmQnk3KACtvC4VabPs4lY/wES5t0t/kUJarz
XZ9gjdYxKyMx/3os7fdYa4Wa1fifPrBO9aEqqznk5sqZyECg9yVcUAFRY2s7EsHX3sK6AVv2gqyA
VliobFdDD8Xe4XXS/rzXEG7RCHmQ/QyntZjGdLcEuZ4zy1kFqv8NMhRyOLawArC3xkFHq3oYdkhD
G3fgcsw7CZLS6B8vwB/NAOSHs3S8MJNf975XDMKJ3p4TyitQj64LA8yqteUuf9nKEfpUeBI4RUB+
NUU286KeWTdqgC1XsUkBrx86kmm/AELq105PpBeiu1gVxhSlr+FgMOBtg3XpvCEj5AukpUkM8yHj
79ByxoUptwEtoY+iZMLK0+GGOyZtJasCPbJU8bZKFcPd202KT7w5/croZCsXvXyaqFwizIVNinUC
1F1Sl+x8yJVhYrIKstXlB+J6NCXMKKY4XfUUvCEF303hyR7hxN0i9d8RR/hgFQtvU1M/8bsVCpsh
CAEpPRxFRbE9VAykuJnCa1S6MYI60l4A6ctgDDWF27fU0HAwL++GD0bMfElIx6kVfh3Mv1J3CRUA
ye8tO6oVqY9qqmS/y6EZXS2Vz2adYEixoAdHzLreSGIbSZSm0AwXNkSRIX6cIXld6ABdqk1/6lbQ
msj/48bWzwvs1muWwI9hyzQ9LNIsmnLXOv5GUXVzYrvBf6d277urx1fHU67InzBAV0GTxdcDtJkz
nSkV8LH6aertQ32WcBvyKC0ZX1i9TRkTFwQH7tXAIf40sf7lbVifaVff08T7KfDKJDIO7acC3gfL
VeI8d8KdKVXmZOlk9BuN7hYoMS/4qI5YAGk1i+6oEokdlkFtmx5W2CF42GyMQreng6kGg+3yto9B
jathQTKcB7lPiVLrQK+9FGGK5a39l6wlnU2PfsVJGQEWk+d0IyXQh3lnqYMR7jVJpcqOcuB73yVj
vYiYh38mYcUIEYNS/Ak5or9KZz2rR513GXlM6JzFdJYTpzFV9ctgiI1zVoQ9FxYlAgXiTfIUW6/h
DrQSWAfRxghxuvqMiDrsy28P5ftMFwAPPFvJD51+c+Nowma3XqkzzClJddfXTZdXKPpLg8glwy9t
KHt11oP59ODWpDr5T0JMZhwAG3NoZiOV1c2beAY05141jzrbAXch1iO75Ux8pv//+YN0SJIQ8jIv
7usvis019qfBAyTedInuPk86RrqxaZDUHt/lSx9ZZlUWjI0Q00n1YpYQ9DfYH2xOv/w5bNhBmEss
hiWh1bJywSUfz2JWpO3XFYh9pQDYeLXLLpobIukFmc6MUG9VLHUx6I3zXX9tU5wVptlKLnNTJcCM
bVDbM+MT99YxLCbSK9uz4B/aFL6PdZ7tHBTreM5ll7klpZNCuk7MBmZcKTqvjK9KDDb+Yr6tVllo
sw0UMOBCHChwsWM5F8/KZR1ujt6QDPtJRwUIwy7tftVzKpY0yWtzAVDPS09lixOk1Qu1XCaXsb5A
vyPaZSgy1xhDyQ7r1AooE1BcfDn6S3Ynf31P1JHWarbCBu2ujttZjZ5BrQtw88XQw5EVDriSBHDr
xHoTtmD5sOetZBBCmvUUkYSkJTKmKcRi+CmoLxkUBeOOth+PoIN3Mymwm8H7zTNQisEWXeYGM650
BwWcGPainNswG/15LutswZeDh/1gSC3dFLJEy7CD7D7h8WWIAWSmLFLifJLZH+qS3HXJ2nW5Er+b
/LlWoloEpU89fwcwEAtIR82NadFXOzZzqgV4jdreaYbuIrksnil4L4G8xR0y+aQ560facHgRmu0A
9cTZWcxW/dUEzCfiRP8LTgXlffH5vCxzLgwo8UeXAj858VH/az2iuOGA4oUwGCavGGPc9oxOiZkF
sYOyibNOFxJDfnk9AcsAIwR16ULq0M7y4uZKDlS0DijVyU+hPTe1wfnWNRvcwzPeY1zXQMIaIP+B
G5Niv2u0KQasmEG22Kr+JgFhV3sEB06pP0sQgTjathaYlrwBN9WxpdBW3x2MetiDCGBUNXM5VBhB
cNRfMkii83qTQQo42cO6GC0dg3YgBW8KrR2T/5GFpwHVEqJzfwlh+MdPUkJ0fZxy8GDmuQk/4b9+
T8JhOFSvVJKRD1c1xcK5k+3fglXT6T0lCp6DpszUtK9TiDA0N/WEsOiAA0VIIPCsNI3e6EWzbxCJ
Sug6VZtl0B2RsNqPpO6/uMEAPVFrnyXLmpWgUQsUUaA8vfH90M3fDtaN+8vTWljnXRjb2RZvQaw3
9AH0p/vhYSq9c1+rs6bXoGfrMVp/AiSRn8Oiuyt5zRILWsPZX+vykmSdHTyfsWgtxNaJ5oFIyCKK
hF5SGUpBZ0ZSQbAoMYLL6yVprGj8XcS4BKys/kOzfWSqGs4KuWMLYK5Ljh9kmTUo4tq+hJCuyFmn
AE11x4EES+nNYG54H/kziZ53z3c1cNuY8W382Qlt6J27yE2I8YZB1zo3QGcwfMemRNEgFVrxu5iK
lDz/MVRlW8I89VFra7rJbQAaRkx+rwPFJPxVCRpglq/7QiK5PV5IA0DOfUQM5ehnApE8O+RIpmxZ
+cSa5ht3TsfyHVrdtvY/6urF3AQRpzSQr0XTw39c8Ul4Cwp8YXTogkWFk5rpZ8cJEnNAk2uATpA7
N0lrRE16o5fjyR2DLNM6Gc/nvX//s4g8NjPI9sHq2fQ4nvroDNHIa1l4e5+zQv0pCWa66KJbmfIs
jCyICUR7dqP4Q6EBH6/r0/Ifl4MmZcOCNdgunA7VkXixE+n49f9zz5/GPrlwbsJt6P02tAP0Q2B6
7+3uWDlcbuNJMb9rZ145F9/fPy9KlhwQjGX+GqhaQE4XRUnyjQTgV3RQzrX8Uh5Wh0XjFyxd9L13
vGkHXq84G+q7F1rpiTENGrreNsEHfZ/ptTZ0A6pfnuDEsgITMHHJ/H1awwn4Onz/xxJ6rneDX9ML
dmdLF82ejnTFY1BwgcCeS17rUlOL/3dHqtjTW6G+7/JnLfnydZX7DSfjv4M38tzAFpUBaxpkhTxB
/bfVWOz0JKZz5Z4mGaeXuvco+ICNr9kZtupeLid3qsyv61ohk0tve51cl8XGMXk8R5P2vm8gw/w6
VvJxeGp+pO+8A7wA1oWP1orqZ2YhZq3xu/x22eVhzJeo0gCWE2EaIbGIK/sZL8xlKWNiwYglgKTG
o4/lWZPeDnAsEl7WfXI+yN1wpxTC+sOITmqwDLXR0TCFEIgJYeWR4+szIVPRjOi1A3rrZrklLLYi
TEBLwJJi2V4ljQdZToRPnS/1fkhvNYd4iPTRX6mp60vCV1DD3fWnoAMP2E0p68fF/XOm2jkL/bdI
b8x6xrz3d/fHyj3++gvhUC919pX99e5ZqrVHhOyImTMbY78/RcWYTqzhHkJT3GsIV0Fn5yTtbzpP
/S7gsA8VaEF7wQtvUFMfNGI4FEa5865Kctif0wnI2TNn6YTz9sunpZyqzi/AqUHa0vg8hf5u/quf
cLlxyxSErveAmbLOqda+fKGqZXb04fBIbbFG2V5ouV1ozlpaGF4ZodOqpUcLEcrfTmCPYLRa491V
nd4TFq8CfGg3laumCmdG4Il5qYvWzgshW5wkBdFSQtb8MJKQn68O+1KmUPr73SxbeY8l8cUmfuJV
wsdBRlRx/xuhQFERWLzXIl0WT5r/or6oT0ojkJVsdok15PVeaVp8buWMwwGzFziy4PWE7w3+LwOs
IpSnyi0J1EveZ4FPP4atiwSmTDS2u4Vx2Q6J2nI1X7ZenHXZw+D23Th1YzOB5MR7/Ky5PNYpe45c
MY2UelR1WT/jjROIMG1rwEX7iSGmB3mKFnS0w0erpnxd8uxWmtweaQRvay5VI+IIfInsRzzfHplT
lM4dzHT/9T6WL0ehiJepsLm4FeEp8d0UvsJCNh5SDHaH0RUbfPf0zwGTxCKjVsEOtcyAXqnfk9uF
2I3wB7cUQ2ThumCEu77BK4BfJu/CFETZMQS85Wes8+8AnnnihIfP+rVMsQo2sVNZemWe6Dnv2FwO
0lpRkUVzRgtfH8A4XDZSQYPO77t8NyXqnZX+WSAuqqwF2WIe/6z1ztUBBz3lcoEcK5cPT6vug1nq
u02vukHMm7IX0aXYeLOiHT/1s7BwzNcklw==
`pragma protect end_protected
