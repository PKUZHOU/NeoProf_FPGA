// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
EQjbuvLX2bn85HeR9Bz+UYkB2UBDEV8QtpSedt3hqeluR+S8oIDB58WUVk8vvBl+
/vVjuOrZoS0z/o+OnkD0MaczToeTD2uCZTCKCahw5Qo3IDhAWksCqZzkUi8DO/Vm
tyYR7MtlWDLtmP7n7HsYhRDZUtRa7OnRqD9cgJhvfoM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 37104 )
`pragma protect data_block
f5I3ihh2duaEnGNfrTCTx5D8TRU6UUdxlXeSF/2Mrw6K6/BDp/oPNF5dRORRq728
1DfhDOqN76bC7Qmqh5kQfjd2VTNdBJwkEiheqv5UiymNHcVvYLp/6PK240j1WEqL
htLEKOrtgHzHfEjEcYWHRXLm1r518al8cghqL9iOfpoX5agrkROAn8MQZ+eIFXJs
0NWUeyDrhSmJ4pEsyrUUnFgHh9p/nxTAeZpvFBV9Sfn01+Er0s/VPF1u+JRkaYkw
9x0V4KVzWn5boo6+XRJUaxQfORHL84oxYNSpwF0iFDxwpE0j8G5R7/rP3bMzRDTs
781POPenNSjvOZUQhgSlIWfpwh0QDqHrlqpDCsyoiSO53BHDooefA3udvaRi+w+f
UWvK3GDLvxbnYOrx+MlkL51pmujeBA+9/vjQewsy5aVEqEl5Q1qgHkWw/G1O/xjD
ue6VFL746zvFZWnb+umS7i7r/iawRVi1H1v7u20834oLdnobUMH+9+yTRmPVGxom
2bzJP+yC87Mv2FwtLuDP8X0a4zg+DCB3SKF81sdCadkO1994Yl7+tBDhWdRu5nOl
9q0k8GsJsrj/Bx9jyg8pWLhTe3XzwEz/O6WW0+eOP00GDSGyhHE82iRRLDTG58nK
DULmslOUgrriT3+1PraBL+JfjwraEe16T+dS6ve5EXIZcIi8sdCcIhjWA8jJvHB1
fBZ32C3qlTxxMZs34sxfdUV2Uk8p8UPlmAbBZwKLDE9gbJBlLF3rYiVmCZJfAGAo
mXpVlNm7OV/qliPYGdymLF0u645O0194OTYC62WUvNHypVB119NlOBp25Il+2f1a
etXwXq3rffycfyElG0kxk8Lut+GjEXsO4dmWUcgwD2b8Z/cFA1ooBYd/OW5Y9k1e
NdYfoAM49GMbzXYxIt61LAGCiu+tXtg8iJOqZEjSnvZnk1Vhkv9Vc77R6qPO1brW
F7FPaajzxrOk146bFarhoXO0ZIw33nNah+77CiT7Latnn1IXuGrJsXtV3+aIIX3D
5AKtOltdXuAJJ+C15OHaKqfcDMR1faNHK4I21s1dUPJoYGj/zRDqVNEGFqM0ZEx6
aU7bD4jk0uD4npPtfy5KBbbydQh9MX/Npr2/wSsQmvL3lWIAE9RiVF1ALlbZiQel
G3riV85zbomWwz82Qdwk4AB9uj1xdlzypQBnJXv3AeNwajFSZCdGzzATd1uRDQQp
CQGJgAq5/B2S4XXZ+sq7cwp4xqZ6sLGHwrmIfzc4g0KIR8ZsnM9hwgqZD3RlGfOH
MiTLPFJp00QFwd1tXf4enmtTMyjyDhf067OI/OCEfOPe+sRUnLMw6d52gftxmJkF
7XQs8QLNopKJaXXdroGCEyKqHkmfO0wBrqBd6Dhob4vYR1BS1CkUXqISf6D7m+IM
B5mNGJqmqWRcGAN0Wp9zsEpLLQKl9hdzRdg6Au0q+uvxb8kENwCfAun3xJIJjAP2
HyYwDUm5GqfqEljt7v1Hi4Yyun/HZG6kXcEFlts6MDK4Mni7HeXfx49ehCkf+tfd
StnoINrGs2vRqVCaEn19u0kQThGrty+KWz2uJZfGAHc+0OGbiQ6HkmUFvxGAv53x
sw6BVCy9KEm1f3Y/JuL13rmNaGSYFBqPB+1gyLKSp/ZTJRdBsyeFCjPDd/myc8vU
MFcb7H12aINgVMAYUhresqWMhcZkGJ0HNSLZBHuzrVtsPK4iOcFBjXm4wGvzweL+
NbU5JuvKZkl/xF+3mkXIqoOf7vzeI9BfGbjoVQ2LskyZYL/DXCALW8L1Lohnemh1
KehPnjnKuL/RS8sXob/bFCn79uvu1K2pPUWKs6QNVDb+n6sVHjDOeVoQ5rpH9h9G
8g4IHNC8Ggl5OgNLBzNJ3vcXALXLnKtq235CXK8kZ89EQrPI8mU6kqlgfoKO9Nr+
csjFhKOSlpi6sCbC+13QGyDxlv4m27bleKHd60cps/ZRQ2XApvZOqL+p41KlTydF
T7/mtFT234pDqZTmxI1+21kCfTsXvZ5PpvnHXLJVLkMmzfCzc8bi2vEmI3dqMb2v
z5nKtgK6DuL1sD+5fZF8YIqgT49t9eqxioUBFvCLr+qpJsu7SYiWs/nPSGerzkKb
szvM3SpAQ5Y81pjXFsh3tELK8GEdhWZAraUnSzQjV/1jAsW0f/U6P8JG80WjczC9
iXVrkRb62Oq49hLmuqnuVfVIHZb5rvSCCj2N2LsJ9p+P5YYPF6CwVaMcB2zVOTyt
9CmtGTZG6jdw+4SPUxOdoZ/SX5eWzEpXabiPzOy5O3He/ELOx2UGFTFetxOxhxMv
uzxK/Dl/HeXwTTgv1CHeY0sIRMdVT06saRq0aoeXHWlRJ/4BKLfg9gOExwMN9qC2
iuipT32LegfVuN48EazJcubpIrJOM9Xv1AfK0yi/3HysZMJP6TNTXD6++3a1RqAE
ExrptlLJTB7WkqD4paNUnYcO5X9QLsyFbQ4Ed/eH15wYFw1FkE0YUrIYWBwTlb37
ubnzKND70TrFmr+dlzfTAWByKW0A7rOGl+LOKmaR1jXm0SV+2kJU26agC2fKWTq3
RvcdiKJIKE3OVCbHM6odMw8exQpSe8HxPsqwiMafiqbfQ5s8S3lInLusgN/hMhfb
FpZF409qcK+OqeTqvjXaQ35PLCcxFQ+TJMtcJ/Yh6dhvr1sBmgbRaKfoQYTsd39w
FdMf5jXT0p73r7yL5y1E5/xTl3kcGQZa0iJ/Rr+0Zwnz71DUHj7AhrE/LlnyRCZd
HmR/1TBLiKUCwdSigwWjwM3oFpf/jhSFzoxuv5IR62o6EYImOPvH7Mo5K/HXSwAz
+7fQjperi0O4WuA286NnlIfK611Thi/sUGddma/QfQh0roKG/bVq2/ICW0k7jtgj
2XyV9wY+hbwblw6HfBvlZMhUvIaOk+bRQvfzawgGcWhQ4AUAUX90z1W9vqBcujA0
U4/JXulNlnP8jo2pQuBQC5WW5ggftzLDIrv60R5dPucWS2HTM6d4HYBm9v1UILyc
SQtvW7yejnhUV2K0zqA7olWXTZuBJ6AKVkXX6f2zSqkA4J3RrtbgcEBeKB2yoneh
zUCnAlPZbM0sxdVybZSL6HMsnwukQomcO9uSDDH+dmVEqRr2HH42dc7pw0ApyRHo
EjInPh6VBYCrVNRj5u/TaiqfawvtEywtTpvOfuqC03l62Cl8Yn9qfC9W6uqWxTqH
abHzW5QB0W2MsFmZq4aObcnL/dEwVzQLupPAhDc8CmNn7p97sIZbQLhGnuDu0frK
KDCVHsQUgp+ItPdJ5uVRzNFQ10DdxdLC+IQKK3K5Yxmm+jMZFh5XvyA3Eauzy+ii
ztCdKYQQr6I9yCdVPdvzAvjj/grUDWtoqn1NZ8btZyTk2bnDurQhCEUcwUFVNSDo
bEw+UDHRHnSmunMmi339khFI5vdNOtL1yd3YNRT35od5+GgyP4NnWmNgrZs+oIkM
KdvvDbM4ZI6n7L5Ptg7CFVOZRBBm6OfRqNfM3fYU0Gs+FYh2kt0fybuV8TCsfd3z
rUBDhpgMDBVu4jOLmU2PLAldL8Tl4L9OtdVkuJ5vWLrzDOorP7UmgAxvWfDmH9Fd
yOu4e0RNYRC186zw54bKyuzBiIAhOtrHJCw0I8m6KTR8Ve/m4MNT0fUMsFzaah6H
ualeD2k86OuiP4a56PsH6Dgt54l1tm8iARCZe5NTbhivJy09szwjtLyrns8geigM
WjlCovPaL0dCLhLKFMwr0XjpfeD400oixsM+5IcnMW6fC+6+/VTWi88Sqm+PMYTl
Vg849dpOfwbGJMp0ZDtKEjZVKuM1iv5XQSTUyYH+QU4nFTL+aBB0Ke4/xP+Pkujg
UMxIOjgoMoIMFF2nsQGgidkg4LyLfhAw1GLPPMkWtIc9u0IXNTnFFr0HR9kw6W4O
EinCnU0O3GgkvNW1CI2FM/CX3/1T9pd9xFJ4cEeztpjE8gEGpbHYsRTwSG2bX6sy
BYkKBJzMDiH2ohxGeYcKF2e9zxEvAVxbqs9rJM+ntLLTjPzW6YArBkeTdgmXlY1Z
59Cc5s41FDIqCdFx6HQtT6dSlquO4RGk+mz6AGPJGrYGNzwO2qD7++27SQjhPmru
+yb/cGe0O3FW/59xMoTBzVe7pR3MeYxI1JlDnTi2PnbcXXyNj9wHXOpnA/tblBZF
a8Qwph9eDJr66EPjCOgVnVeL23vJqxffMr5pUfLNmcCW21RmRWrw0yUp8Wfl1EC5
QBPnEeCEmgxh/LrpEGvrUo9XDNgNuoabhozdVranz//UKaGRrXx9GSbcVbP51TXW
sprKjUyp/VxnDvgBm68iylNcGE+ai3rWRYq3PgM5kz8p3oG+TXXC55tvcrRck7CW
VjWIKPyFNjcRsJh2+tj7w8CzbIg/OrdQ1xdXE8SDOD9BoOu4nKmihZXBts3b6ypa
YD5O3h1XKwlvIOneOwSpmKwXdNWrY6vD2wY7066Kc7S2kNBuXJDwCjcH6PHRqH8G
aMpXUMzgu6oo707X5tvhCWfDEQPHbjiZrXPHMf2wJfWXx+sYj/NXdvixDVGaNWWB
vgVaeEUJnhYfToA2YJSZE9WaUBmcK9h1G88F1aUQ99CzUh2QNXNNU4eoLr650KoK
i1IC+3K9LjjHj9RoKiOuqnJVfjtQb2mJgwljE6AQ77OANjKSumkoWsd6gByYhfBM
QLksiLahkLavvY14SA+JbQqVaiXAsAVaEdRMfQXueMHI9IQf/vkHjT0oh704VFwj
327tnchpnQ+nKYAdHU1bZDSkgxTHAsIo84UV+rRY9rnAmJTpUuVshK1/jxqINfko
XtzQUUrIyAZw6No+W6JZUQAD1udpXVcFuo9rZtw1ajPO2SUW7BZ+k3bEAoTQFKZq
jjFeFMuhucazpqDfGDhzzJRSvAhiTMTUI6M14sZidhLtliRcRf/F3SwE6V6Udy00
syKnbdzYbYF8GTATO8141s/H/3nUYHw389m9LPEuAsztwywUS5sptMnYM+b1nRbZ
vC6JLSe6GAyTWKhdzc9JVUk92ku7ADBbQTBt6i613b6dlkpP8YvetvSbRIOldrL9
ia0iwN4ZZdCczBCWGJYCexgW3iHFIQPStIwIjL/CVL2/FkUcphpo2pEY+nA3irNv
LZPxsHtP9raWX+5+EUmuyGpOlW39y5uI9V6LSC+mxAZmKTzNeFE8U8yzlPrBfcKo
DDMlebwR6CVOgJJfokty4Yzr5zMpia8wa+QtwAAmM1dBGc7azBSORaaKIyqZNl9Y
iUl0THnt4OKnJ3qmGvvveGkwJPzWeictsZPxLsGfLGt4yvD21WWJyGexwIM8pjdF
0H+sXsYLbR6T13IML/r63Wvs5YivShOSOFu9jnMxhMH4w5E684nOot9wbIiPQwRb
fdvzyj4ha5IVrJrMNh2Uyh0Tu2VgqCTcYCj7YzJV3hscwhkMr+mcUz10aBCFUpiI
Z2toauNhczE0vW45S+mca7WHe8FI3bci3OpXUOWSqtAAxVoG+XS66Y5o1MqbSIPw
arMgjHKgNoFPf54Vzy6udVy3bBmHj8LsQ0gAro73xyfq4bOtXL5IQHDi1hCSXrPC
ZyxjDIoR9CxFSMaqED+vEKn/qGpBXV1HGXBgnY6lhIRetPqOTarwg5/Vrqz8JMTe
nABLehjgK/fvkCqCltiJa1jShxC4itJeoTmuCCkSXbIiORlKZX7Sy+Ofnh/p6YTY
P37TgX+6AzHj9lVVe8ged8w0SjJk1wAWjWnWxfRFMUbNnfL9nelZE37bHIwcag3k
LGjvsM5MdEEuZweM/s6FhxjXeRv3dxEfnv02hQU2OgE0UuzjNBSPB7DSC6c0Llxt
5gB+BNtgw1DLN555npS2+uW72Wcp+U4mBHaCf06KDBJnRrNmglo0ui6VINGmk9zW
2ua5q3JlS4WfDAopALt9VCPy+Sif+ccyYv24Nvdts1eiSXx6bkPGZ8q1wdZBnuUr
W4YDBsUxTqKknz1Vr8x+lkZvd6GckCck0ATcOYrlMIRsVAzWp808VtKnTbaV+9JS
7y5TikOyJUaN1q6M6vW+xtggE1hHLsQY82PSF8F6+vm3EkGN8/zKtqe2bQ6M9h9T
EERAjK3ub6BeUvYb2kB/mGNQl9Fe+26k8UrN2sG4ZPv4f1GqNOIsYMaRhyIMD94G
Kh96hUPYnj672s0AB44QPe0kkKd6THjxMUHbMJqSLybsEsrUndHP+8A+MwHwnkYk
938qZAkGJLHKlet0SXXwlzqMR7WcJfaCNRw/h1m1JX9xiWcPb9dwWiBkNam19jxk
7DTU2nET199qWcf2hrcJfELAgr771CaL8tWjjMRLa+ElYFey09XB858rrnUxh/9t
s+y7BiSv4cn36+ne9XV5/L3oO5IJzgC23tOaa9ZJyX3NtIN0hK7EXHDvc9/7va78
XXEc9TxydR1NGyZc/V8df2jySgJwrFRkKmqyeEW12IHUpWNW2813lrCNAtCdqXwl
s/n7vtLYSBfFXAo9KCYmkDHOsSGgw0ZuC46rphG9N1Xey46tNllTKssG3sl37ko8
rxjxiLAcOeCjcXPgghif/Ht+kdAW6J8YV630BsEpgfLU+EXyPQ0jPBlyxBs+XjDm
0rqhdnLLH7vLbbFZrt5+jZwnLM2w8EZQb63mLYjzzyqQIoxk6z5HC90lz1Z6UP4u
54COfahw4NVyh6jKCn5T51ypjOz3ZjgihmCmtrqiyyDvJFY6UroYHVY+9W/89vVz
PASQ1hxVXkgKMFMZMkiVX+WLq4aGABTk8Mu7YTozTPfWE9cru11fUyMF8O0lI46r
PLFQlwKAWZR8mmT24zK6xWZm52IbM3YHq1mmARsrBOV8gmD4YqISxGvPhcx7AqjX
cWGO7xtZnt6+7VNS9GjMxrkZA7MGfNzYFn1it0vG2G4NPODku+jIQQiyySmavhZs
UzSft1rtBazh7vQlZ22ZDX/nba4orq7WSEJgizDyVnBw7McD5LBF+7CLMWouBMsm
9bCT2zAU1uAqXBbhE5U3wTpYYIEAONNYA4w5wMy1zLWGciQ7Iq3VI/UNITmwhqi1
h8m0bJ07IVMxpNfNqMzf9y3x3dp5vis08CX+0jNEQk/JOd+t1qV55OmtY/2fES2U
E5M2nK8QeeBJPKrkC0XLFCJZkXdv22eUjvtSyC8V/xYWi62JXhaG+OG/5ArPHQx4
hb1PXIiU24Br7kX1Wpths2KhGws15mt7pgY2I1UwhcEKgGW15jhhSLfkmOg5o1Vz
bq/GkEKGN8xtfwzMEmCjsCIXADBtC/rhI7VqLYGSJpH35CYIA9aPGD0cCXmvoC5K
EYo7Ql6nw9duA31FAomrUULSZRIQqIYdE6MSc09cL9dDhyBwQ0lF+iHhoemyTTLt
7oNq19pDgeQrVMZXaLTsI3Oc9MVwgv1PM7EcDFOF9Hdzj6HlWSg8fdv9+EJ3adZi
wgRC0UwcpJ0dSe/P+crJ4VLtU1pjOnn23MWr493Bx55h/TVhDeEYVTt7c6DLE7dB
kQX2zO1fl/zu7W0r4afMnVqXP0URz7IBjkKSnqLK/Se1RTe1IHIPouHg+cK8VCOX
6blhDyofqZBgUjK9tVY7Syhi13g68rE25MumyVAAPceXeP0JUSXMWyqiujReRP92
1sXpEIilrvbkkqwSoD6jXxHH9cdSqsYCxPnz8f3eP3NhELVOseYZKAJW5+HUuaqO
7eewkdjuIQ4Gw1VazE3kYuRHuCxhIOfo/00MopK4xQ3JViiPMXRPdSxYGbdl0878
I8ooqerTyeC0cRcnN7+Kdlhz+lODAH/HB0XI5H7qizAF6uuVwPMBluXoicfOfByy
UzGNMASwel0VUnDJvxvH93bx08GVOuMy5WeXhLKGIzOn8YazU0ZFhGekeAsxm38J
OQiDtt1PH8PDAJakoFE21xUE2xJlbXTjJSe/7i9Ej+IoNOmI+nAvL5qRZBI0o4Io
F6btlwvx1flJsezv/g8FNBfkWus69OVq4i9b1dZwANqbsoD/YnNdoO00seA9V8e8
auuf/FYF7OrP5cBz0ORwtTtYglgXEU8LUOJus3rKjyq1Rv83y7alGXgIuvlFwNKQ
ZsAN26vDplkmiJDHyO4n5J0hWAj+EtPnR5nDCE6WG/ILGkBHmjqq2r/UDdMu1FeG
aJtASNcjFNhJeB4oeP0/jbzmA9nrhJmYWmOl18t081gsC5r4BPwgPqjBiNLc0Gl1
euan1pa++cnxefmVQxJqo3+U4hayKn3pjr/j27mTeKfSylqAOqOqJT9+FV6Iyj31
x4yJOA3qZOUycd0CSYCYefsl/0+9R7j1+KNruz/pbRfmpXNJnMI/Q8X1d2Htk6Nw
kkPh/jsZhXOSnLIHcB9W8Sp1ilC0MsQNx4SoEMAjplz1eSrEY1Gy7YjnNA8f0CZk
DZXr6S2pW0UVQe8t9zrYHOguZ0RVajZIgne9i5QGBDlj8A+vA9Xr6nFD15vI+0ej
x1KT9jZ8eGiJpNi6SkFQUqs7EQnRIu8BAINbpymgNfDlmel0PTNpFp1h3bNxQsB/
j2diYeG0p8GjOuqtvxdxJa5TtESS8e4q0vIqyxKlj4bln1QAuiOM5NflgwQF37r/
6CijicZiLXM87FizoqlIziUZXSFQwhTDWNCr/hDWjtkfe9wzYxbkp3qJEWKPkJkx
J7Cw4B5wX+EWUEnmTI9LfcV9yaTZgRJ+SBVYLbt/CZTh8+5K3hONFAaXyQhNUJJu
aWTDCI4oNDVMNRLbGcumKPDzpXzDGCtnxjA6cF/wYgp9i1IcBqUbU2FHNketH9Ug
uhdtyYwgTCaJWKttMd7XwW+kFsyHuikuQxXQfAWXJut35RLhHAMZdfF2w8EYq8Dt
RSQdvsWkgHtC7UNlOkmB4LeNj+sm+gZhqBG1dvRtC5pQ8m0inkOyGJOgTgPGns2j
NZ8MKTnjlTRm5kxoPgyiI6vldkSJZeG6hX1sQ2TxOvgLjfU1AiPP4MsZ786hC4BD
kPrGAF6+3LL+lt3y54A5VImuGczxSEYy51kZCuOsIMCrU0e1nPoLUUdVwEco+Ji1
ZG5ZIfYACZhUfsGco6v7FqfDFiJjj7Ve+B0IF6Dvk6ixVtjWA3a49Yu1gepeAOFc
YT4zpRR8J4jez3L9UCWg+a5VuxTxafkeS+dLxNvvfkfauxgOfAE4kI1awmDWT/OY
zxbcJyHuogjz2IDu1cM/HGjwcY1Bc/CGfjqXXmJAqhGjgyaPjclPsuNm9zSS6CIg
t/yj5+p63hmn21FRLUxrjU58NbfRV82GjZloTbLOsZ6XPs/OVj0mrAdfr2g+wwC0
rYUIORzBPZVsx8FPXVQ5jtCdJ/tWSjzmpAIwjdbtHe3Vrl8nKktRlOM+4Hc6VlxA
CFL3ZylvJWwugILz1p2qwI+avnPtHyKr4zB5bdOj9pk+AjOSaCy7kqZqiaKYZe1c
mmn9M5D2qR9/eNTu8h1F3UIcyROYwajgnvj6OYVU/Wd/c2xMN3d46qnj4KijRFSP
ldYnSk8lpbGyg6hu6q9+/sPpQ3ZVaoUtw8Ybv184LZqmnDlhkqY5D1RqOitoAfZw
nyG+ulA89DrAKhICBmix/CkHNIrqsBSRxpyWHCFSVZf1DzhdAV1/JBklEPm+JgEk
vO/caqGB58HixQWtMp7WneeYEltT0W+cV4gi7ytsAXqIO3f4NgQ196l+QSmSz5py
VpvhpePa37eTMONEDJEclxfZxHBqepzTmUtGgAlbaTUdLpQkUfyUzC23HcmWmSlE
Z2XI8SqzJWWgSZMeekk2xc3p2dMJ4ZWsNzZmgmI/KVUSMgjATZ1A6iQVH0zV/B5g
6LPhUYtXEkGyyv19Sk3Ii2BtiEPqvnW0z/WRBW2ZLIZ0OyIC7h/q7z2DLf5rPqWL
tcwypVPcLL323dVO246mmAJR/lZb/WrnFhPWAYJZjANLNoNTEvKMQnumci8el+Oi
2qiK+RM+au2kgKIaOpDsoHCP2Z60jKEZv1cF6LO86HmTBZWIpmy+x4tsTO8wXngT
MPJxMsosSmj0mck/fErSL3uSm3UINARC+eZdBF/xewbPMUl4S7Rc/cg53+lz31Cl
uT/It+Joc07uR431uVvj8Cpz0NW8pBbYXWtUg7M+cQiAXlUihT4FLZLOSjBe3nT4
RUlbBgBfUnI0Elt3T8GGcF6M0DceWnrIhaQmbVVgMUE3lNLMwRaF2KKRQjVzyJ7l
Bgn/HFRIYf2DWQ8Rbm4xNUSflND3Z81++wy8B5auq2ZyxuzsOaj0Q3gOAWhSJIOg
RT2OBvJhVKX2I6qGEZAJqaw7+iCQnI0/9LjMAyQqMsQR/6+vncLCktV7XFudMqtB
dAvS6ebyAtxQyhvX2T8lVUw4QZHMp7TcBhHVDzpdqHOJ3EH1g40Gjii0kBktMIjq
4pV4pkySrQg+yJW1IpJUb+gb12g0/ip6wCh9gJJzBmYUdHldM4H6eUm4xgetkuD3
Q/7cMOO72bxufMQX/p+uDMXrMwIn+9w5zXDWdQrssQaU1IvB9mBZpQpE7EzdxQ9O
bhLDDwQjyPl2ntYSQ+cJvNwu0Z/ytQ/R95q7d0xSSwGyWDCuFkHU/n6ZPMRe60JD
xU6YoYzvz1QYhmZtqzfdcHNeWkLcWQnHI8neQc1bbldWr6r1dPKIuW1imsUodtBZ
F3fUJ1CiPULINe1RDG44nrEP3GOrauC9KQHBRXDWLV4f/bl7kqGevYCp/hSid8Jz
YlajC0Q5NNOT2P/icZxq8daLAgSUbWZpqiPrmRWZKjuDKtT3uAhdbypu/6Fq3t1e
SuoENF25ImWn7VhPZr10g+CJ20wAxFSjaq06c4eC8mtOBcuqjb7Aq72G+bkkUnMb
N2aQY2d0D4S4pke7fP/Lee/F3m43o4DgKfMvT03xWxE1yRfzlgY7vhbz/dg0jQDa
4jXrwkoiybfS9H4ZqRRoMtb0utqkXqld7EzWgC4cHVvL3YG0XBOUlHwRAboH5das
wAuNrPgMaZvc3T+qp0eyfdDzVZY7NJfti9J77/Jg8FAmsRqMyg53w3sZy7EJXhXL
KsQRqpmSzeG7ugxdC//oWMzvfZ+Zun01s5ffzPNcnmUHvBXk+IQfIrFoh2rxln6R
LSP7Cr46x6EUAE1FiuUiiZuZnS3aSQ3Z6B/e9oUiyq20C8VSxGb7mwS7BtPHTzUb
ewndL/s2sz0W6js7gFXxN1uQ1QRygY5Q+GNlLsCiJP63KYsBy1y44PWk6lvLi5rY
A3GMkYlmCpew0d8WUU0e8m8YCTjR13EoNeC8BheT7cK4Ryhua406iwaXVShhcS1A
/Kq4f3mMENRMdsNk9DWoc0/ZlE50GxmAtD0Sno9n3/Z1s8e2IB9aMz6mfuCOOr1R
7jNBwspuN4LZFLLhSXM6HOA3E7q+W/VHsCS6Lqtuw3GX2QsPUuP3dGt4K+sG4BIr
z3GFDfV/Wur5g7kpJOHVMniSSUOCOpSNnogf1o897CNsBo+Y83Ww0Z4qvnrcV8aE
tKN+qkkKgonFreEhKDE8GllHZ4aO/1ACAWlnt36IUo1EJKjqS9gj5K5W5dr+syYo
8VZVA0vBnjeu+uL0sIIOcUGwfJDemIRROOhDazkAnXjyxsAYK05+Ax8BRmjhq7BL
sJjxaUlhUFXzavJCFip8b7NQpNCakYWh9Ct2/aC3wBROnPV0T+GU9F1afVJxSkuI
5Shx6CfyF9Pa5RqTLaGRdcJ6SStairkdKAcF4VrNkSYXdtCnSJ6wqSsXroldbdnG
nbw8O4cLtmvdkiXHefafu1OZAMcvA7PQlDP9PlNRkh50zoJ0iC6WNm79TcrzjJyg
I4SIMBQZW6C5uVUVX0hSnmEI3Tx5YOtWvAQC283Qgc6IyWjEVMUrELvtSCRRgzV5
vE6WrPz6BMzPrTwMC6wyAdNujRgurrmKvPi6/r2tXvIl0Sufb/WEAVyBx1p/q29y
yQxDxxI5ysIgs8bE/lZI4/oqU8puNp6It2a5eDJoI2G+QLZDhR3RTW4+d2LVPmip
sA5TpMhE0IUB6pojVz31NcLlgZgtRZFZSvU9bSXXLmOskVI45KLo8EAMmHAjTw7D
84h/x5Z90LXWESlAB+aqNGJofUXMXJ8SoSAAcDaRSCBwUfj6TlpJ2TsauO1irihY
BcHRMre464fACy/H4j9JP53E4uz79TJiOaQTQ7eYpVA08y6pJIKk/GW92bNx7KHr
Pk/5+CYdWlXZs6+tgupDzc2EnMUI39tsehvG73otVC4kkxxG3tp3PH9YXHciERyb
yTFLBde6l45rDcfrInlMhrffCFv2N5KeGHIkc+mMZUirZV2xRv2XWg9KTdcUFv8w
vI+CV5BbxqooghT4Q1IK8w2T9aj7dQQToALd3ET/DixMoa1HelYIg580gKbnlU2t
8doXtxJWVfqitjQsnHGLJ2KtwWU3UCtkN37SLyONyn1V0YaVGDH9XZJCRiFeS08g
D88QKd6fjEEMbS7KvYsR8EtgYA3ACPzz0T6mttibAxU7evLfzrF1h0lRrkCHmAFs
6EY9AJsigRESlyRkME0uIdL+PNKQOk5vHitgvA3q50d17k522TTi1mtwlCgKUsdc
AgDhI+UmKUJ4LXCLsie2szVXMw9kXUELmps3G5dhuH5PbEh1vxJQiN2rTSLRGpEo
h99hgy64urBQB/BhDjKqX+XbwAp9XwmrMYu3Y3E5P20SXRf2/zmG5y41PMDsXBlw
1GV28YRX+UJWGVAtjn+NG8E626FEE7341RSisbbVGrygRD8b0YuXBIb6gJb0cr99
KH+3rkY8rH8mIWDHGM7LqsMvDz8yCmp5CPtKKVLLMc3u9OUuXgtXKW++BTYuSLV1
fFBDrjox3OQYrgPrOGDlU9sU3GctndB6A+cdW0ScXYO4/dZACbL+B4FPa5NGlxcP
2MJMHXLC446NbhFzAsARH/2+MpDJAmO5YpfNdQcKVrfviJH+nMeoB/phbLQtXPLY
ukHcqnr6kGFQNipLoIiDc7oL4W7po61nRy2w96wj6QdkfLw/Nrzad8NVbXsGGpkD
p9EVaBdmlRW+vAbUIYIVkqtUr2nIrYPsWTLHvfTmZsbLU5I+Wbb/wa+2/xX0DWc2
XWhB3oMSGbMMvBodVJHw5Ay8hhp/u/TWIDxcYgreeAOHM/6jmX07rdXB5Oc15oHT
cHKmO0UGyqlvF6wdzYZQYEZB6ZUt3MkKaMlglbpE+5a8B0bpk6oti/FMRng/DLhS
dsNIHjqlFZVm/KloUlJNaIv7v/F2FgmqIb+hbm1o5ttpNKySXUKG8nZ+t3hJcGB6
EPNKONJJ5jJynXt1ZTgfzZN6W/s6P2pcQl1Vassmmk2RqiXr9coO7F49eVJFBmtb
TBhirfAkkYcKQ0IToCZMz65OchMr60aAzNjg665h8CHBx5cNv20mA37cNHR9F3Du
XPsT24hqiUnWYC+wMS8Y3xrI+C0o/Hxkc54+JaMhhD11y15Jo9y1bIf5qmRbomoW
CnvoKW4Kwm/wNUvTYl5vbbvkepfCg5pikJkxeX3IWc8i0pKsXWnJy7O7b0Y4JTE9
Vq5aq3QOCE8mfM33pyd0yup/R1iF8RGZYaOHPupHSJr9JGeuS6N5WBS2pfIJ/JB4
LqDmOZelXC8kk44iLZpkw40urLEIX83mfxI/PwnrHLZH6Irq46YRHP/OrfcN/5wf
vjIO/S0oV3sd1YoUIPgcOo42O8r1W7YIgwDpBAtec8ikerX+xVo5X8CdGETDwMQA
FG30QkB+KkIXuLFME22GkJm+Cxtn0NPzLyKQwvy9Ni5/p3GDtq766gemOTtJ9WRv
Gs5nx90bLcNLC5aruT3m2giL/fKrMgnDl/reYqByYKM4bmX5jb90IlCUXqmM7jZC
J91Yw4Ov91Srx8uVMfOhnMZ6Dcesf48e7Fum0yJhrI9Rv8csMOCqIeCrueM/CnXR
dyIGaxzfSN3M9vNSFLtsCxSZs/rc9r4yaN87iYZzslghQ1Ad1RKouvLa34L+uLZS
uRMGH9z0XLAgBDc06EuXLQmhFS6aXapREZkLyf7XEUw4jNZeE2LVKbW0Mjc8r6/s
yg5wTGBwb8Dd9cn9lJzbmfKXyxnbJVST+G7qUdoms8ZMOzzX4nGrT6Mb111xY/04
IdceVc9KeNMud5YmdeTAFLc7t+I6o5tC7mSJsxC7z/UAChxMc03xpx6l2yAw1tB3
Voa8lYCUAO07iQtmXFZ99ZZVAiI4fj54VP0/Iw80a9G+/VreQvIEIb5McARY+Tbj
tT4U7dahjLxdf+LmBsaG7j/lhUH1m5FA6dw4QJrpYvpLQsRLvb8jOuhZHRdNLGpc
4BRe5CkQGqgIbKIlrFoZID3gf5IqTKZ0oOM8BBOwiLEkbsnNY5xGz+VR8ALDdcR3
uLGN6EUJLL3KGru4SplCSHhwvDPeRpYT9oZM2pyXZIqxvgUrnBlc0N3lTMmb84IR
sithxGSr/18XZA7aaReLvuUc/xaQpNxqBeuqs0VpxGf1Ifu7NYfCEmuVlNEBzeoz
YiJQLstyWew8GouP/0ckvsfUcB91Ye1AtKLklS4pk8rd9UYvAtSDTXH4no/k9ZH8
gTZW/6iQKCKvqk1aM0dCDrFxZGjgZSfvFdc5/VQojAYoiOW+YtXejTTv9bJrr8zX
BGyeHcPeHsYnfvcAD9B0ql6yBRa+XadBTAaqLGidyag6tanB0QtpQezr1Pjoi1ti
vLRYYigv9k5vGlaK8Kq5c1pc70aTLM3MD9TMRrZ7AbuoFGu/b8OoHnAeIqd9mBZb
l65Ww1cEBLUMFnaMYHuY+/7DTfMjZdPM2anRCKkWra9Ooyua40JzYfuSdeI0K/Pd
77bW9lxvwuxpvjcaFs59zv8RXm//oxezz46wGBIvHFRIVp0npAiqlvFZ4je60UIt
UmSECrnOt/xf7I3p/nuJuPJ5CDahiY2BhmfC1uLeuyJ/DpfNaw9FSFW0jgNi+sKn
qt9+fDiy7Cr7BnExMcJDUruXqYPSTPYYgnuCE64JUaUMxPWfEJ3W/xgO7iPG48vb
2jb60Zv1nw86q4CZiIvUhGAvVDyRP0+8Oa9J1B1aJ82jANlJEeMO81RgThQvDxkA
G4n2cxMJdcJEoWzhUZrkb+mW3QuZJVqLe3hasWvrNiEazcQL6K+ufVaQFvBIegvl
WPBU2RTs3srra8Bt6ecyApjw2kIsYDAj9hxpxBN5/V1z1zjrBgdKA8v7lArAHAOJ
dwWcw0o/3TMBBHRBP8px71GbUzrj3wUx4Ov+jqPW/zoDdw2dHU6LGyEPspiK5LSG
BAP89FSjRsPFiImdggBTopd6XN7//MDjZG/9CO/aY89UdpTwEu0wg/mZcyH9HLQz
l31OFY0vafX3Yhy5SS4Rs8RqaG1yxTUpzl0FhY1DkeAITRl1eZ61OB+j34p7NrZs
CHOzTIy9mu6k3GFQfq7jD8gfydRYx8eETe+7QkquSwWgC5n8JtioAGNiUwMQ5NV+
7HVsB4NZBc6tbs7fgLr/RGlMlnHggJnrgDeL1ugDsLsrUAceXk56E902bxg27RMB
3HU9tkzlzAvWF6F/vClCAjb89y61WASpprcdksVICgu0PhsyfDKcSudh79m4oXZ/
zgMXGpIrRBKLOrtW3pUrAEVWlABccm8sGODJHnb2PqxTi6hW3dEjk2/rYZ1EvAGW
R1J4OwJ05qKMdRVaq8BsgtjWouZBXrGItH02+fymN8Nc9A7ZYBeBKBLNQ0b/Kt0U
fDGHMfDAInksFFF/Rpo0i6HlNo5f97k0bXkEiJ1OD8nmt/N9oiSLT5xLMFOKQlZB
7EZmusUTgxZMMdvz615zaroyhM6u4aG3MXBni5knQWF/022ojQ30h8oa7AvbOQnQ
ts3vbkRWjYTDS5oTjIRaBx/ic6bSgaCJMisEvmloFBTH+t/2znhsjlO7LCtf+WHs
o8HToq21uzwyV0IsU3swlpmw18VpXab8JFUerZGNh+WeV43CUij6NJ62iBmZkXOI
jjU02mm6mdyNfjwemumjEUBihGnE3JtnNmt+G3rrE/gLRQzUFZ4SHGxh83w+d0lh
aXTaU0GoKx9y25fqojV16F3JNzttfwh/8hZopKJO5CRz03CRWIsUq16eQUsMwbeW
s/rXnR7kgBImHlV7veNP7d42OU1M56qg3Ed5G6OdPwzKUhpnERFITmGSLjB9s8rw
W+q4YG5vYoro7Tk714v7dUrIE1dkBYJuJ0dJHeJbCq66HX6tmL8EF6bBF3B9PHdP
Cme/miWb57nc5L6kJ0fn9YoWI9/S+W5+F4KQnAopt5uNM7ixu0oI0onWpUKHdPg0
7PB/CvHuyE4ZbZRL9eJ7uLpVoVRQGpK6glLBOzulr7bxJYMjHtAeJw4v3ub+CAED
VVscR7kbSgpsxUqW63XbrgesSLu6M4PWTIbBX4aN7e4yChvI44gqTGUT/wbOSqjd
DhQsWkzmatH4PJeBVe60irXCBnVSvBc/Pg8CAAG0NGtrWowVrH2yfz7I/ItGznKV
eijZLmrtdGvQn9bEuX7HitsvzmCBLJz+aAo5gDvirSnojZoG0mR2t295km/boJnu
2HdZWfAX88LrDYw25ny6SIGoz7yRf02fX1gGj06n+5idqNDeLULopgt2zHK9Mhcw
XGV1zQ47dSyhPSQfLKiXhD2tkaYCg/nz3OvylBnVGwhdcbQCJ+KMs2rhe46RAQQC
aZDbPivUcgnmMKEDkvHYDApV8SXBt8vSZiy2O+O3uz++uQcBYzehfxRbStyIY0xz
TZN+lssaGfbrPXZzncPAC7+6pQMGuV0CCCcHv0E6pF1mLll7Xb+9M+CGQJnO1L2j
hlTDBfyC+5CrOfeWxs8pEN0ueCwnb0Qrs7dWEPAy2hvJBdj5cR92J4S0bJBzONAp
Fz2UTlkvvPIJOPldz7r9M3OLenwHI/oNNb4f8HrJ8x1CwtbD/PaNlJfeJx+jFo6R
X0sch2bqUmDQsHbDeSX7yW+zj+wV5TEv9YoYFl+8amzP3VcTDnU4CzJZ33TqZEsU
MqtA4FGf1R5Lu6fKTDOjzhez1wOjU5g0471ptRbL25gRF+DiEue8ZRYjsznjyXtv
bpVTvMqiXvm+Rufe2QSHkg7IMFjyLyCEtPsm61gophQGaVlE+KKyID6X2uoVfxBs
IYrIh98c2bBeajqOYrE3yCkH+2fPKvI+wpQHV16mEdGjnkX7K7LL1bDbbfHyNUYs
oWDp4kArudQ9oVd3pDpq1Lhjwm3+W01bFsWIC8xJ/y6FyNHPD4QCd8bZfwlA0IEz
LmdxIR0vyauMTvy7Fo94iW+EEDTAXAgaR8AfcDZ5UXKTo01fekVFzrE8VghgEJXk
g4jaLBScn3NJZdpLUbjIKKoDjskPVHlRGn8Sns+kYSgDnG7lhi9B829fNV3OVYGC
4ok1bh5sXJjiVJEIrI7ViwvIvSls9sZ2t0wMmPKhJhi/66rEpHUHRhc1H0GMM35W
InZTIn1Tq2UwCpKSWveh/d25zWgjc80a6axhXD7NanD0lDiJn0JvVuAk7fYP7f7+
9KvfqOwGVwfGB/KXaoBHhWatsah6ZwqeNHbYryxJr8Ij+RdXWgA4huTGHvQzvzTP
sE9+ypfz/4JYritUJ5sHAaYkBRl5nom0S6RjQNDzvB1Wb1KeQxwYj4GLhuDqZZ4E
BzSpZNTrONfEfBGRZfs3ay5RVsb7fA4Ipixb6c4AmKgec4QQkT8eUfP9Or1UFgKS
MVWF01KkhYHtXgIJLJThshtQIN0Xiek3wFLEfwjCGexEBwLd38SUI1zOz6Uo9LMr
L/X+q7DX+wK/t9Ku521GRFFMWfwjYDLz8wxfU3+bDCTVg2+c99MEuzMicFYooA8w
IQzGDfX4C6HHbDO5K6B7qKbvLWU10Jx3nhno34lOByhRu2+HkUOxyUzO4lBYw48R
CkJIIp9YQkhQdiIzgwRXSUKmg0r+ckCGx1vXQkvBOc9TQgRHx1pIJmYVLwqrfi2f
rN+6PSkIQgZUTpWVsebDx8yK1ayvh/fDNxkcZZlEixcF5qMleuD6aBhsZSfq0loK
4fopS1JdcEmS1pl44t5BttVQ8Npc9r4BBQiyGIvQEWL3PGeRBuCT9Yl04iOLAlbh
enr+xyMi0xO9UINy5iebVv+hsWBat79qTJ3t7pcLJYgDEFTrmN2boFhHZxBe+paS
yGGd8ExwDxLHqx/YAlEKj+MbqX5Gg2tMiUDGsg2oLnl/mXmq2e6u5wjYJlbsddaK
6MLznrauRt8dSGl5ax2aqT+Qtxl/rr+kORtsgylw50I5nmyVUICh+GHvns8y022R
wCQHNGsu6yP6S1wxBvyb8B50SJixdfPDjsrZ4D45C4SFz9N8n650qHLpuK+HRvBv
jv5vMVpfn2RIiRYAhlZ0PbfWOpO5JQGsPfQwXjU2p5smiMLBLkXgXAaKQASZ+M1S
PMEX44z6tHICSzZQ/ExoJCMzpjCEKHu5aJ0zaqmnzy53tW4BVsZy6PZtYvS1OZZc
8eQnRbPppqAPqFhWjFvb/IGq5gPXyr7xHPu+kkk+xDOiMfbRrVlyYbeZT1rH3YV1
fPWGStw5oFVinKUEhrZGiZTk4nR5tpmHbdfhjz1SuAVHDJYZDP+EAt+ypGam7QnL
n5HDxdzpRpPh05q+NdtJw6Bg+aHcCoQfLyrcLi9jksdLgplOhuLQVTWYr1pX4+qm
93ngSrT0dwyLQnV2P1PzOwEAq8H8H/OJVILfKxarozsZE5ulA/eeYtJetmLZrFRB
24bq0POnl29IcPf72Jx9wFhIZB1bQPaEWZariqAfKyeWKdLIjxHr2dS+gh42FXOL
og8mvkWC5s/POrNftNjhX9K17Ce2MZelxVOl3ncH7eFlKRhVCqWNmFL7JsH+rwkz
9JFtXqDjgdTBOYhB14KxWjHp44cy+Orxs6IcOo2/OdhU0weIimhC1cO7xwiPnyEy
xRFpas+nHpMZjMZg/QyzobYAl4USFjoDrLmowgmfUOTm75KA0aXruPM4aCp81fKw
bUtCw/2TPdKq8uGPZhNqXEM9OCTfwLNz0rTv9Ad52aeSlpstubiLV8qx95AhASiP
u9do1c/rMUnovHTHHOPDACQJYQS/1Vk0qUaxCRrBjk7SEsSAEUUl0tFVgoy951WB
ej8SRGo2zrMS3e/TyYwNn56rvDC0CO88mudUnl9+6d+ggSHTdns7G3edUs/lvjCS
/LqKBxQ/aonrEAv+DRjcWg/v4EGeLuxbzl4RxAQMh/48yY/oJxPrEaaavM755g7w
sgngz1YN5zMdRIj4OLFeMNX/FLsjuDMFBDX/ADUXuS5qEV4qESAfl0jct8u80zTN
DUBBPkq4rUpVl5lUogKL3oJOtR8GRU7t4yhamfq0t4DNG7T3MrWBonjfn6vA5RZ4
rkFz3BbGiNTsAZS3Pa9h+nw98sSRp0SYcvs4VU4ViVTu98huFuo7sgcxIgKBjJaD
eFUWJGSW/jadbRdJW3vqnXEnZ53MA0ZR0IN2dO0bmmonZnsR+RBgnJZoCmDkyuKZ
U8vOrBgbNjhXKWq6Jl3Ntax1NLQSUf8yhrLuspS1nMZnkqbMPRO9BfUhlfBzBCm3
T2aQfLle3SgsXe9XYkGlZ/v18d1e1rpjFzmgv6kPC5/caE/b3CzIkBfyCl1nO0HL
ulMSkv04m5e4V1iMNYB/oLAY27jy/NCd9WL322ydCznq+6wdop8PddUIEtf5yF9j
5jREBNmpjAp9aVDdqkRHFPvLn7E0PrT0BcEuqAMAmfGz0GyVmCDt6OdxCbp8AcI7
f7DtxV0/mfJkHAjz2OV7FxVGkWUBIl3B43QQX/gvEawOUp8Rh39Zx+aI7ucPwAPY
wPi4W9k5KvfIXVTwtAdYcFS5VRoYW/bbpeo69m//f+AlMc1/Qe/uaSRe5ZwBG913
jke3YQwcitPPBArHTSNlSXI5qvvXOmASo8k/irts6eVgFbHH99sfwAp7DILfkhn0
mwFzuHLJ9UQHpAOoDzs6eKC/cU7RHwh72qbd0ie71B0a8auEMESo+dxIl3Mnj51S
I1Ag1DsYBHz47mDE2feHkNrFOWGRljX1+d9aRskXRsJFTYaXcGHQR51dUQfjjlqO
610+Zr40celGJLVnG4jxjQft/P2vmUYqiqFiSWXX7ukrAsECuqEykHcK3WYKXwvN
z8RCVVOE1rwkrRcCFObhVOimf6BEls8xFROCY0mlqpLPZdhS/P0H5h2M3HdXezaR
HsMGAg+RRhOnWEWw+caZiV/kJJ287sqbn536bIzOKbjS5J+zVXEBKR5WRQkqsZPR
BXGxMdSRjtxI4rDq5w0WRoA2i/sKfunuWn7quKLWyZy1E0zoOii5iMp2NH4kLtbo
jRb9ToNU57tMlFFoao2F3S4qQeE3tLQPvLwrzqDs5UNICc3p6AveUBpnzw3It2IL
1akZTAGzfn/VbWfig0kGekZB6kszAgICI9OEsj4+qYcavFSYuRPt2t8otUV31Ubv
G9qHHxWyEJ4niLZuLrqNdhM6Iw6948xEC5ggmlMQgAZ1lyV/OOYwuAYAwsf0wB+F
gmrU4RsI4Yt+vwIViHIXbDeU+QcyctRhYAEL2AqdaJjOMcvRdcDbWhjBJSQgGznQ
i+d+MW5//CoVkOECTv09+Ig3hE1RITuPfU8F67N+Wo/pZF2KpFwjEGceYsBdF7jH
94Qe8/Hv5FMZGBqQ8CxvcPpCAfqZLjfXPIBr5hSohxw+kaj4ct+36LcFAB5Nw5L0
ZNK2cgRLVVntGidZgqsbJ0HpgWz04/KNsE9qYxE1wkeLCz+eSc92BJllLwwYAXH2
g1J7RSXeyWHGOMAn6bXBEHmgx1+NLNeHbz7EeTGP3in7s27ttlsTL6TzqAtWLRm6
2hmQd5g96/hDs2apQmZSozX6yCWOzD4BXY9iVWLTnPtF7XSrHOB7t1ddIdTZgaLE
EqfNozywBrCteqZMopm9xih2dpPud3UXx0ceipqtTSNafC+BOLkpJAGsSZmQcfpJ
ewQCp5L0HLc+BLWzLGH1ijICqAPdgdhh3Yt9h9wGWGiKxHQzrp8bffLaJdmu+R+p
ZwL/yGM6ldeRwog8t8JvXSMZoxnllVYn67XviDnsJMN/FBy5z7C8irMWJin3JS9F
jUge0sPcCgLIj+yZWvgIyXfea6a3mBvIMFW2wO1VUFkp/NdW8xyZzsV7L3j9rec/
jZHyOEVBXzJv7trIJlg7n7daJTPwKkA748s6MaQSPRBNjsMTficB3PBv9NbaFomd
u1OMRiqhXXU+cqr2WeaFyGDOTKSn9Ch5eEo4glvWFUT3VwYBtmuv9vWqyQoERMBy
TKN79CuCiQrhhbWGI8koyNd5WKGmUAooxVL8leFaiMnlyJ6F76Bi+s0Raz2ulTjB
3Ykw3IWONrAn4K9WQRxVnEd+IZBKI7fbyQVX2kx/rXEFm7JITGcn9F1HNwhLB4Jt
hIRvpVNDT41+TmO7cPBMRyj8HMWSa9vnSnh5tPHGqV82Eszz8vTHOOsFUavNowej
aXBC9oj50qv2sQhOqsnF1HdfuUsdVR68q/rbudg+dXxDg7eg9sy0o1yjCYo34xjH
/VaCgk3CH83FdQsem/EEenBX/PyycyEsK/BdJMIn/JVUsjYSXrq0I55/yKqrRj7Z
VKuB/qduFtB1Pdzr0J605d3Hgk2U0AiErJqzorFbmTXbzztoMZrbSn8tk5X5SVO/
0Lu9xHHiBqSe+ggHcwn5qvc0uY4O2xF8+vncTq4VrvPf35Iyk8UHZzpYEN5kPVPZ
v1xbl4/zcH/7IHN1wCp9Hka4LmiTjF5lEVj3xk5alvqMLFsJoTnU9WFAKAQvli+X
LspTKBXDjmCUiWNQzGn4VSOZ/TJ5FMOQWKaqDcPmUBgIycrcu0r/NNBVGPyfWEP1
oupLY84NNb+N+5gN/pXU+jHrrbrvrE5W+YBM7PcBgKNDuo+NcO7GGUHNvmd9W/74
vETIrQZ9DWqpGsmzZNohdq1uQRHMJg/ztXAxsOKRMax1KcfW/XFSvNJviu8yG0bA
mkwxMT/PhgiCWo9OTFVv9EAwtMhoUUBKRnq/vG1VXFjro/jFmFlljMr5z9Yky2Fj
lLOFa+f4aGXhBKhrZh2dtsPIdys9Ih+DwTaE46jYgd2DrDVEtinWZd4PokUWIrY6
jIsj2aGnodPJuzgsvzcbTn1MzPJMsnAHhA4ZnmF13ihDaqZ4Dv7OCcdYRBU1Sakt
suvkjaumOa3j6HPEGVL5WhUniTRIwlasxsrE0rD8ZmpTwA7Hkcy8ioBJZCCdzpJw
S5qFj8OMnkSsoE0k8ws3gytt19+eMyBiBx6CH85fPBBMiBfKs6WSv1qbkkS7r7Ko
YnnyAAh5x6oYMcKCROFQ+29tKXSXxHVdrvwIr5zgFrWeVTifRYAPKzaRAGgzhMnz
KfzwqJIiCZYisFvoGKywIMIjqNonJ4rqUCrck8DR20UK2qai1WtM9HE6RWfSERsK
x+z74oMLmgANC+8iZUewawoVyllzBYnRPOw+1NLuJw/B1vtTUXAdgBn0IYez96pK
JMUMBNVReIrUwPccA2qXYf7BKkNZzXwtGT5MxrseBPajjYj3syiOtV8oYsinzw/Q
b2A/bWTXcwYnPaUga+Xa6ZANG+CZs7pmLeAkjwwPlxcNTubL+VJtLn6Xu3iTIPWx
dF2+D1ohviBkQ6pkRDuKjXo6tCwjzjIu7iKb7MMKQLyCW25D4Sl/keZBpHt7cCNx
DzSz6K1pwN/pJVPAksIPgatx7ZHVGEuByTH3FBOOdwM5Js2fa8NuXS0mBC1OZcKX
tKyGaojAS6Ybl19NW0hC8ZvIsmP0H6MaJ6QW+1DVCWX7L9YKw8po0y3XbVdv+5yz
aGDF/NkqJsGV4iRogDxxWUUAF3okXXQ533MK70A1ZQ7PFkCunLIYs1rJC21p5vD0
usEyCh75PklHZlVJBG46jqmUtUHMZ6Tl4S7hNlWtIrd0XPY4XPq8Ly/jSrPE1eC6
McpTJGsVvp5IfAMz+d4EuNpPorgLCkVRaL22A2zMBWMWxTk/aLQwE5FuPmLW6JMW
3XDdI+qr2tw3yhb7oHJIs64ap5ZcFW81nsa9wiWEbe4f87AY243JFwRdDoeL+Ta0
XJ7Geq3yuN5bok/W3xoGVTKzrUJTZXobtom9x3TTKjpKBvdqIXLEg50kbUcQaDPr
Y6p/UH8zMkzMphUJrqhlPwcs8oUr+DXaW4NXNGhPdKOApfXG1/Jf9e9vTo0+QQBY
l+OzqJViguimSUtJLKwOA4x+b/ITh+EkOlRHULrlNH3XCVE0Qg7MuZrh7aU0RY3z
nUmv6gFr/H2J53Ycb4pQMy0qvx3U9+49oFVpRzK6DbSNU0DTzDDgekDnx8GhUv8q
ZatzEDu/YNzfWR8KPBirnCLeHsfSSjdXUZ5vdMJjUR842528KzbacZfq6xooBJEU
Iw3s6HQZrJ2QAwP/m499N3tBdjA1MPS8H93M2Dn9koHyAvkxnQ7NA+vpgZoHG3uS
i0FU8M2O3rHi2wP9wrzQUns3NmQElzHxEzk+uJmY/D27YA9ei4+XBr4eyWPX9CTi
qySuv2ITOQnpYHubK7Sis5mwK+BT7BDTMAUp9bPD0i1/RwwaKa1n3E7i2spo6Ioo
d34ffdfS/c2lYKDYtjn8octvAFUbtgjXfPy9odC2EIHxbfqF6mIVGmFHeHFw3wV7
fJ1pfiENA5YdotaBhGlNW5DRuyHkKVswOKdN/Itads17wkni2f+fEMg+t3y33k2M
fIw9t8LNwOVAo44RfU7Q1VdITiP02Ht4/2cX56P7g8tPtWYnCKbgS3Y08fa0QmrT
D3RvHGIss9QWHqEKivifNeXnepfu+wDvVdX1WM0zReYzMvN4OCvXfMRwWRExRxPL
+A996FnaxuErA/AXtVA9TlxGk1n/eTUal0bepSYsGPTl2nDBxl9dMjZgFmkGBqDE
6amdzGKGgBeyeINdwa/K5QMtdB9JpogEYvznalsnQZDQMnxR9KB2XbWh3h6DTQjZ
m7+gFGGxDGCqGg81Z9Fd+KVNLorEC5bYTbnv7oTGXqNL9E4kcpoxzuc6V8m6Xieg
QGAVAWu4F1ejkRYNsv2dXwXVG24D8k3hZNriQQEk7Q7ddbiRgHli+37lVewPV1vC
3BSPRX8TaTcNeNY1+MQMHP0QPglG5pEwsuHvxoH2YoAwrOFziJ0kBGw85r1JAxX9
mjDj40T+rglA1J0Ap7FQxJcHxP0pnJPfiyPhLpiEzl/EtDEzq1jK9UHxTVbk+nv7
jRpu7hLo1uJCyWQYiGiynCJOLs4+s6KCTJGV7Eb118hk1TKRxaocw9xailI8mWeb
2err42fzS02jSYh06+YsGNuJjwhdM9qNXaR/CLE2NyzelVD/VCEuX2yNj5mDSeQl
/6/yENOnHHPSMoin3LP7UXq8ygVLVsH0KNwx1gsPyG7SpBEdTdsEuufI5E/BTC0w
2QAD/WO1vQWo+Wt9hSijy03L96bWMW5BT4/u93BkF2Y3r5xrOmN9R4WGDxqWlOoF
LoiQCWSkj6ZoB0IqJYlbInFqMg3mQb7QOhsHGgqttROQmmR8x1nLAzSuzq/40b3Y
d3RHGlSri75oFYlQvDL1FvSwSBzWfyy0RyVNLZrJlktJ6zB0o/zDNLZRcDGMauPD
wFghcghf7c9czNQr17UHbV1rEY5SGACtGU5G3Rs6IBagO2kmBSoBuVb03CBnQUXB
FdX8b92YkDbBUuugBEAON048GH4UJWEMR3t4adrrpUPspmwWfmxYzQzhJpMkuEkj
o9Z37xRBg6b37dKb9bb9fOhumT/hlyBT+fZa5O7J7Q9ZD98s6UGuqThWEnEl0Bfm
Tg+PeHo4yyw0bwMBRFKSI4/txP+3wdKguAuwdg9RDvTfajD6TDaJEfVF+pXjZQzJ
85KsSwuaNHcUYdI4gyXYySR09uy8oaoJpd7EYtgmYpfmU8ILG6xILV6zS44U44HT
nfrP59HV5yaxVqmlMo8dxRmY5FpOdGLzns2dJtVWZ4RKa8R1crM1kVKTGKMbo8LQ
6zprA9DZFxi3L4TPEUIkrSCX9UijeL0GIn+Z94EpWFpjUJUnzODRrrKDKrVNw2yk
WAJAEOrGHsabaF1cTMNxNrMXXIdIyTLoxsqx3rwCX9Q02Ne57tnjZEv1OPB9RwBL
Uq5pnpw4nSrkOR5vSUIVJZOy0xNvD1+f0HHENxAyKJBZI6nO36te4rV1tbSLCM4+
6tPBIfK3vf+39xX3vym/M06iHWws+bbuASWbHdE12vaxXd0Esz9lwMmrwBc45heX
MdWS0A+5B1ZblRvKO+jnlSBdrVFyS0rAaWmPH6cQg6yDFUAafDo49tBYPbwPFVIE
HJR43ASN7bju5qXY6lnaiF9gBdLnESW6Z1jv5ORB5UH/yItLeuWlT/fIkXj36lE1
TrQk/NVNJNIuZgvI3dIfT31+QWeXXgvfGGbKLcAbJeeYcO9GitAITKgVKpOoU4Cb
pdMprD43rcb39x5PUX/WlMATrtV1tNH4rcOvPlDGkHd9HljZsFDCU3nM+RnRiCtJ
+XMsL06YOeh+i2E1pNyqBSs5eDTzVXt2BeARBAjeGKKQqBARS7wg+4PWGbgJbZvV
4QAVszX9pPotdYvQz+PCbZJGo6EKaLiUeNZ0I073u1vNq+z1dyEOvk5IX0Ohe1yK
hDs0tGT73QZ4AfKjqg3WaRrgTd5ed2Kny/cTznPgEMWnC5w5iAEMsf2Wdyzfdytx
lZEry4F5XWMs2TVf06YwLXUZhsdujbyKaZeNWb9TeHatjTvkBDDSIseUJCQzGnAN
WYOIa+MboAe590fWIQlKbSz1+Bb2vM+nvAORO9TeuDRYGecQAVcZm9KQCl0Z1XUY
VKkCDIaognQwAjjTKI9SeDBdi4nKmIKbBf/H1E2BmURfUWgXzsqipN18myYZ2vBf
xJ4zE3cOFwFdL8YrroI3jm+oshp53VlL/EArr68v0aGxZg9H9rhlUJSqTMm/8j0s
mdaLH2GKzTkRH7tLOadBa064zH8NdHx5PRl2ohMK9FPx48+IJukvBvU4UF4HLDwX
eiZcDKFr2XBYUEJ+ATQCUHCVKTToRwldfFGRGhihyjTPZZb5yoJjLQ4lmF+gPxng
BzZmqIgtvtob8pGO//PTi1dpGvZnOYMG5aaETmW/hcae0XsBuUjfKREB5Thyf6nF
qPJ2LtawcVtHgPDvuiBdDjCVfGNra1cHgn1AOE95CO2pKzCrUYANV4DWKcGmeedb
FJheufSrPkRJzuFiJEhY5kSC92Nd+Lyp+8KnkRbxXUxC/3NwZDKU7XLSocwOgd49
nzNe3WbZ+xvPO9mVGHvYLX7LSRkxEV2eg7rFZ+zqVIqsiqciwaDAgdt60XmI2nnn
VyPw9YcmR6NaJR1papDCcvISk/j8I8tOWNhuMb59SeLA/pNkHbHZva3xqg0AWGlt
Cdq6/OedTRlzXphwdfwjI1sqe6BRlZUzQaGmDBtqnSqyjuMFGumigk/G6ZX+Dti8
F+OqMEiHn0E2MYZceCC6lmR3TSqy3oTyg067WKVWrzyL+b1p0vF4bVAIBBygmXW/
0LuKax91/yd1HUsYu6FXt31JHZ6HOcj0IH2jrZNp480mb7gkZBPUmyB9nDiPr7wN
kNLPXf1/RgOCUXbtB/7idLwF2CBu0uWdEcbf0puLlAd8Id3kHUmMFvCv0F/g5h8j
+Td0QmNZgVlSaE20fGWMZ+lFFw24ELwmAJkGmYRw0V0X6HSC2Mh7gu3BAeYg+m0V
mC/QxgiVv2WLY485cnDx4Eu3QqQRnnPDRqmwYwNO4Vy6/MZS6M15YwAHlRmS9VXL
T/PZYH34qmjq3n1/9C+lWxYpb/qcbdOB72DuRkO5/u5hJqIAPhTkoHAjr4lxzEI+
X0JpwsEP1/LLsbkweTTUbaG445fd9/GtDO5D5sYOJ3fMIAp+hXGBuw94/3LQpvgX
kNmLM7fMmgoNFyFZ6oparI47RPCiSPNvNgzwNcgMMpLRQ9PpuxeotCR3yKZnf2b3
a8NqY9o2sm1A+pOEDjcd/XTtjYlsFdfFYpKCFHbmR70hbOSBg5Ih/BYmmwK2Qcfj
txgydEURayk/7k8hD+VwulIE9kVJImLKU28KL5lQz82TnFASmffUGq/soBYUXNmn
khP1+OXl0D7nc7pTXJLxeaUb/rujiek6dkd/4kUC+oChYNAyvV3PCbqsQ8YNPtC5
fepz5QIxI7ib1JISw/iC5Lnh1xEs/lk6aRbXF/SIvCx+SCNtYCvvLqM2oPHle/kN
GjhakpiGLOEvTx0lifaTHT8/D9Ujrjs4nxnxKKuaQmUlAL8DO3Sh2Au/Zk30O6XJ
I3jmWnqrcydEZIEre/vW3nbDD4ToU9i4NvN3T8TugHlUaRdGfVWp4V7T+uxpUbkv
AZQvGHnl5i3Ng9LtKSrQ0bTQPM3MQIjtR/xt1uUkSCh1iuMbgNy7UJmKlHntHVYP
9xRm8ABL0HGVk8f8UV43MRwfAxZBpBt3+SMKZ3xfgeJKhjBqYQs9sQH3DoV3sXwK
36SUxiEuOp/uSXDbIW5llUdLuk4d9buoyPfG8K8o9NQV0rW1T+4P3UxObqF6Wqll
myOJvSKGR1bzE20BhNxqXf2wl8oLakj1M6LFsZ3fgQDrrv5d/RoTs0fWCGmDWO6l
qmT77nPHTvfUiZGIPrvDSVMjSr2M+PfgbYuAailsO9/V16mv6CFv1mUOrhFIyCWn
F5/H7qxSUMoMrZCdz8YjtrLRGdm2hDvfJyZxIAqQaB0GzORugyVsA9QlOviej2l4
NTHqqKfveJSzvw38rPJ7+mm4OfugAiFoM0kbcqUHwzTjYSHaSBQXk3KFrxea4DVT
+zVwtTVd4UbYR8R/j8UYpLnWBJ7uBrtffFonAD/oGFIBt6PhiY5hetx1rMyEgjae
ZTE0wRuJ9rxJxMS3K7P9vZ2h+dVaVRn0tfjdS4ahr9OZJMpGRA0e2YtWGQ5Dtn2a
FiebKOYTteirW1zjDuuBWO7lTOaTNKt3m2XtSYcFWUIjA719QNdFY0s/9aQQnkAh
nQgl0340FQn+hYW9iYdWtz+VqzgzxHML67oNaJQBGQw1mf/rShsrpgoq0FwTM3rU
MOtj6dKU2T9ksF/noeXVoWefG86g4ob7mDO35eodCJKO5+mtEYiMbg4FLCmoWR8+
Y0ew546EyS5UvnbM52U3vS/6mUMmgm9dXwdqWclSrgqYq4m58jaiYS6U37WT4lX8
SkqnCMbfvh7RjpPp9iDFKf5HYqTodUgMJL6TDO7Jzxtv62GvVE0YNER7fv/2fXyU
XkWwDqqTdNDisWjuZUCwp+jqvzU/PXd5SWwwCIRz9hcQJsJmB5FZ/ri0+wyk+ldb
VR9cnV0tVCjTUDnwFaXrGtTCDZcX8NVydmRofdW8IXqudKGx505Q6XR+Q2XEJVrN
qCK9ymPvUIw+rISDSjbDd2/J2sf5Ts+B83bqJprGPIxzGwhNXIkU+RlWQbbPkSBM
m78BQ9+SwFyg1YxPW9uSwGo/R6NnzYG0PrJzn3DalZjN48T6/yWogO2flx2tL/eR
cb+9EW8/1iRVgS8BWzqRuVXs21VBREWZBq2TuplWXmLcLqED3HX+88dtOtcHynXg
QhABuVinod9n0VbMHdnNN7O65wAeNmXPbQTq+1uXsXhtloUgkMiWO0QRZvzkQpCb
uaIbNRrCTbgY+55jnHJbCKaMJgxNnsZBC+EDU4ec4FJDY8HG1U7QdCiHmBFn+A8y
WnAfxMWJ6Kf7cJYB3HPq4fy7O7XGVYVdRV56I5CFJJbtw8OUlZoTtEYsmWvux43G
ju87V28m9meR/b8D4m1lWdaYYSzN8DVFRATJGXwLVBF2c/E3o4+dGIp/PVEIOOXo
r3s0e9aw1kwj/G3Lgq1yxmzjY4fWyuNKA7MngPceeWtZhUAI7n4XSwkBUwqHNqhv
EZ+2ZbMKkvVIE4ia7JkUvz6N+eN0KwhwsurpJp4dBJogSxrZBOwJ3ru0SjhSSRt7
A6f5kEmXwMrVx0SCeb1Y4A0zvm+s5/7HsgwDNKW1Jztn9VeTn8LFugWsP4hsVtKI
XR1dxB+QLhMh9WuS3+C7HCW4oE1+eFLBOA9kCJTo28cHD8LZfPbZoCHQqbzCrehL
RBSygx1RR8hgz99ZkMlCxXMwvVUa7NYHEVE1P2lRnFxpgkXmCyeSsoPXsUEXezxs
6jvgbj9o/jlWP9Lk159uXW0iqgY9TGmBMi3GXyYdy3ZxBCq2OQYfj4aZMEKoNySB
dK6y1C7+7NbW9wCGf/bGMIojCuFloXIBfuotsrMm9b3Ic6RV0Yqf8/M8HuWNOt27
oUSAHRNlwF+X4WeuGbBU3pQFZ8OckB6RklM4xV0ufWOoZCBsNh/jmaCPyB9pPfo/
4hUtnvyHz8NDpS8VF9OF1VyapLmnuSpdqc2mgsiNZ4bHhyPTPD4eNOEUIJKMflq0
0HGCQzOZxrAgBWjvaW93tFsIC5lTjJOctU3VSx1EjQ+/ztyrgoxKnALco2LDFU3t
cJXjvGFMgXxsA/NYjRov16nRwE+qsQplzhrDVq23HxjzdrR84SgJelSzwXDG7kih
11ptYDH8NtsnXLGTklk9dYgbrf7f1RbVum9BeCJaZK6/3eN6VCwo4NK5ZZeP7xGN
yc5oaBfAavp+JpfIHu2yJ5nLFPNz1Csz9U2gXrLlP6DXl+/q612JlEad769ne+Dh
Ouneo/fyVTXCeju1gxuVRTmYXsKET/eZngATOTuORtohmHtTHz2YZsg9uHdAgr9Y
MEXYOtNH6ImLdv0f1r/bnnn3e6YbL2gDHrJbr0oMFz2ucyJNIG/2Urn/ff2EgXtP
WPTIUkgBX4sSM1XnV05+EIIwtGaGjWpd3kbt/ElWcfcKUbnFRZO58QI0Mm4bprCM
mEbj4zC5I9Jl3KQilvh2rZyL6crCcTCq7wqsSgzfII7pppOak/yiig0JgrgyuLN8
Vxjr4IhZtPi4ZAY6uddH+UogAiF03dWBV7uunLM30BIKSAdY51HmPGErzFK2uBMG
2nNCXuqGOgfbo72TzaH7tCXGF1NzscACvPhP1rkeAcALrunGw7BoePTXXu3nUybv
il9v7ANWHM0ktVbZ4K8Ubk0VEN2OCOcFF03XZVWo7ouIyCVjaIqToZo2aAQpDUGp
6Sfg7XGpvW8fbOUByKOSMFvJpKIzFUdMy/KXlLzV7BJzj1D9RcKxkO7TEZsz5l1p
KApddYi/DU7EtmXuGP4Xt44anUBAk/qfpF9XUGqnYqpJfqoXCLqOe9IT3QGS8Phy
ZbEdObM0JRNo+dsFK+NKBkO4Yjmny/WHou1Hgc2OeEDzmc+EHaBVu/RuL/GIqLWf
3cCC9Pymvk9Mlke3T7Ac3lFgepiNeUxV/ydO+0V1l1xOL/PQMg0GbfTV9k8s7587
nKNkIOSD2ecsGgfhAJCKzVNkQhZ/wrixog6JLuFn7cZllZHqZfXXAJEUZojf2tRh
oG163UQ7Ucg/7mqXhB2gy7GShg4yJYQAvzegHNvzH+axK5A7pAFt/vnkWl1wldZ9
69HTAIe1Mo99RMxCbNDfvaNR5xLEkUNtIGBV1b+N47TOv2uATZlZ7UnFZwu5EjYm
Rrd0A7VJwMVak+mQXWWq46OfipRVtmZmj82DsGIiPUdyECCwYpUjj0s77NZxMu1b
TZyudRoJXmj79KqwkgpaQsftgf46YjhZBAx0pL/KYMH/PiE+Q6yhd8A31lDQna6g
AYXWlDdnKuAzIqqHnX6OhBCKoqwOfClmxxaLwNSJfFP2IS1jrPJC2VxSI2ZnpQCG
7CXKyRE2IeqE/qsyxfKZAPIQIXjkSy/0KkoLQAUrpM8nW81L4yorEOWBvwe85wve
EoAzl6JxP9TQYUU4exw91Kwf+89sThwFz6bl306wghemofIz6q4BQsG8HOCSTvnm
+uWrUuCSrNaM26bpQrWU5cUp3QPha0l8Gdh5PsbbhxDYFOaOY0rNIPggXTZWDhHW
ROIFOzGnt8gQZg53HJC/BqAhLpfPKMrcRC9JhN+7LThOPGLXKrF2LfZUCE/BZu0n
U+FJCvGdQGVCV4s8EIPdNYhxAJY5xsbI2EGX/kcq/5Ep5VdWKdcMNmsMO5KmAqDX
ooSz3DkTU0UzI6Ds/cy0bvTSI1uMLczEv6SQCzEow3aoyp4dyI94lsrelqukoRFK
9FYa+S0lpDNEMbHBwQhScON5Xt2JkFvu3i23gvTH+7CZDVL0TbAGMjznemFjJD20
da/MQ7aGljv17sJB9+RLC5B4cIdOYQDNf9tmeEkWXw0OEcjhnyiKcO6eqnYT21YV
lBU6PtHe4QaFwpIZg1/bQPp9YgokEYGIL9aRQd00OmAf3HOKGfWmsCV/O8M0e78W
YUN4lvEgGLeA5r//VMfpxkYFen33C+fRwCwAoVVtrdrCEe/WxPcV7GDvvE/I4TWU
n+hRdg4btNTQjT0UR18K3pbV8iZx7kkafVtB2iGO7ANfA9+P2NVlICVgp5nVtT6Q
qtUBsf5JFpUT343vsrrKnCLahfSbw501Q7iGTRzz0d3b69M86mL0mttUN/YJPhFR
+VyejeFRFUyxmsPn0vPP7zB5fCBUPRROSt/cz2RHhBirLqwFUINxfBO6tKgL6ZJW
LPhR8ElsxVVzUskpY8xRAFuk6FRN8DzYCHOwsPF2m8kpLJNUmOL1rVNLD9cvfbNX
F+1THNwoqpC8xfTcxN5L92bqDncWqhwhFjjoQIp2pyvd1fFdGrXfSMOL5hU5TAZT
oQCJ1kbGeNa5qUZ2AzNFNDn2KsfMCi716uAsHt6QLgLk5VA+kQdrlm1z95w8XRh1
gLe4S4djDM9Bk5QSY6wnTXvb/QkHC4gihSq7pRoX0NRFiSJjaIjW5WP/wOIItwhg
0QJWjBVJ8J/hHUSvFNMl/w8AeQcsGi53pyWj/fw256fVySZI1wE7HdXDwQ4Ulz15
7mwK+6XEdXeHCxwhw5D3OZTy33u6aVx6mL2Wb6tTd5JqkX/VE/kjlRPaNheqmlST
k8zHz0P6bhlamYWrqiXZMcXad372pz17cd95klBLqh53mY7Ovkj2r2oPXktPDACd
eABGI+VEMXDbCt1sBhSf1cgYBKoI846Tx26rnBG0nRdJaDASyISU466+PAPbFqbl
BJKP2zf7JhIu9eDcHSwAmjAK3lE/Q/dgEmPVx7q8we3ph9fqsQmAGpUu2VNyrQn+
ZOt/G18wiYyCOn0QaAD1LUT9VBE2wKIkfK2s1IwEfB33CWaIMRcL+GKDPeBDgKhF
tZeAAvKYoAJo3P1ZvyIVOXPATSBuu3wcJmogFJhnxf/olzZ9/j49lt4YUjIN36EC
evf+6DcGn4iR+HD82+40sJrF4DEzq2vqwMmKzZcy3jNHko+qOCdD/PlpNuqF8EBD
9BEmmKgvul0aBa3vO3mAzFRy1Itz8AnLrZuaeOsa/cEy6T41Skjs3NMe2b+T7Sly
7HwTH69hv2Q7fz4sABqULE9/bjjurHJB8VUm5vlU4zLsKZ9omOlr/G8N0+qCgKh4
KuFbPHGYjNjBj+Yps25QVz4M8aPGZoLmhjOZS01HamSP9a2vn72PiByA54OHhCZ1
0YNMBaCBqNBK3TV0qj1aP33Z3pAx2BuYgevmQH9E1Aahjcxg8OHsEL5eTdwqlmwX
Za7QiEJCqIN14fDeeKTf0cODk/S3zkAJw8F+qdSqdE2m6b5dQASpysptDDu81nqg
HR6z25SJN4dJSjzYchhhp8GddAKAPelVcT0vWnokggwZqzu4W7DYbg39Gd/f9RVh
QwWNpAUxMkxTb2i+vbQW8GBNH6p8iLK1EdF8HslaMlkrrS/8TitLjq9lBvdE0L0D
mN1Vfn+KQLk8f5yZaJBNlKHc+87yEGGIpnaCrz8G5X6Vlug+eS3vfvhS4ZJ4xOoB
dI2sT+dnkQjlorIbw0/EZNzS7HX8RY8VROcExwvul56Lri+g7uv8YP3xqecp6cXK
U0r3S6Q9Sh/RDZUDnrBn5TfvZdM5tYpOgIfrxG0pMqu/nj/E0EQW9DckRDv7aqnS
ZBKQl2vZNsNnT41I99D406JXqemONTfQgDY7jAuHePSk965LTdT56MoK/SCM1qHA
nMAmPexpX0G+ifo/9V7wh6wvwR/6L6IJiq8vP4w7mXJWGEe9vgCpEphAacf5U9Jo
Kd5ohSsB1S/234eQQgMgHfOMqF7GhM9TOvntpjwxNXhk3g3uPMdzUY1euyTbFWxK
hXoVFk32ctj3oPdsL3+cHCrNMB4TqidPMm2yJhx34dqmVpVsUFPx8LEoIUSdaucX
iO293likt1QmvWQpJiLxg4LaZzYQuyIXVvLDPchm0WOFOOHq5KUzLw7MSv7dA6ng
EX9nxZQ2c01KVcAPy4co4MdL3HQg0suOcce77usJA8rFwgFF66Xiyw1nS6EPS95c
sLOgRAd/3h4pvhQ9nce+14Q1DnsFFvfvxoM8om5kj95CHH4Abdz7D3n+ZqriKlkv
AIHm4arSSqSzZ+z18OJ8OhQCyw5Z804cmXwCiHNgDhwRmlJnR0OearVlqRTrP3dt
VodX65a3ZsKDcFk89cOgbLPTxh/T6J9wFhVIrOyP6puu0JshQAXFNhv9/C+sbdEe
qBJSV8IaDCQwvlUeKOsrmujsgIxtc/A/K2RKIUZ96ON40QdUTglh9mlUsPwjE79y
s95mcJw6rBncjzJ6qoHeponx6MiV1NTA3k63Mu6v089th5K9vJEjPrrm6F7RTdKM
aPPAvJKq6qVaDhjDTVcZvl2yg2IfrEe4940g2a/rREHZCkXsswoFp+0yiWAvhZFp
kBAAMctN3snchOUeIWOcmf77hbOLo3sUCVY3zHJF15CM198/RW7tRJZkHQdS3vnk
msR1YQm2yoxn9Mx6XKiz8TCWaw5tL0MHF6Yj8hbWRC3JUdeFGMg9XoPARAhs0LEQ
AAiLnpsdYGMXbvv11r20nH2R5ZMBteaOT1ciASM7uQmwJ5qruD1OmtUD96Mha0xK
Z9wDyIdS38Sh1OHJtE8Bg5w39ml0FR/ZylMJzD0oqhG6f9LPtp5XtQyIpiHAdQV7
SuS1O8uO/dMBMXIgSRXN/mrDpYvHBzgluopkyOc/PWcwUvloTdaCnkrn9AZwPEuo
VW/Z5PQXERQ2/8d46aIirsmgI3ZWdaEL96u4O22DHCJB5ZrMbPfs7CppflzTRv77
41XC1ugb6GRuVL0Zci9luyeDI/cWUIaucWAQfDHiiyfj7sshnaFDVAIIuofH1m3Q
zyDlq1cl1qRzB7A1+SKxQGaSKPp28qFGWE49iZRK1JTSjdrnRuYsIXKxAYUwQl17
fxJdNg5LjmMWP506EDXObdhad4/nT+PXiefvqAG9/NgDX9KDK5sNHpQZ9iH2dxK3
cxgAD4g/DQLqdJgOxKpZq5a4NFocHAqeiywbkEpqFAsTgNXoLm9Dw8aiTzAtPie+
fX8jqJ0wPG5DofIzRpYMf4rOUsSMKr0B94PXtKav7wnTeSk6VKQE9yhDCTFnFewd
076Gg4FfNbEcxbuKbU4v0Zygs1tj7WUC5uZL9TLN8pMiE8z/GihGHSdqOJGz/MMc
j+0LVuIS03gmjVzCjIYhRaFsr4sOE/HfZCLv3j80yR/olH5qrtaJXBlXYY12HB/k
dNPyz73yKQjJOzjDVFwg4ZEFq6PuG1xLUAVGov9wyauoqvHhD/juWRRAJZyouRqA
ObEtQOEuvScGzV07Rcxz2TOy11P6aEaarUTrxvj/ie98bdN8g6ieStyeuVIMYZAQ
uSTRnLq6q2SESgw4lnxnJT0Iq5mY0TYmySET4WH9aU7MWaS+qrCzpi/moIJ0AHhx
ZsmWwIElansqGinKKrBIvPooOo856S8O43hHhRZ6MzGLYgCb2hqLKSDoZHJzXk6h
yiBJtT6x8gLGg8zjdVMl4z7/YpCWfcBozDE8fZCsiPwu1dApLoriI1hn4kKpP9DG
aAsAYVZxEXFBd4l3N7P2uHV4GvjydDZ8yQMYZognpVdCvKghTsxdf+2dDrKgWNkt
fSXrS0+gHrKokLleCZV3gxwggPhh6J9IlOO5NXhdG06GWG4vESumVFqFVms03THb
PaTdn3QbPycW0IFPBkxJXzm668VE9P7vODGFrcp4lUj8etu2vBa1+hwsLbkuNEo5
qAg19GpQVorPTuKSNqUHBXDJwjtGROs1V+MmFR361pHP0CHxqKR2TXATfYnFYx1r
u+5GWcywel0eFCW4cIdS4H1Inihf6zA0OC3TyHJb32oEceGr16Ewv8hFhB38h5Ii
DbqV1m+udgG4OO3aj1wb9e+SgJYaQYqF34IWwRdQVoifEgBJdEQzE3dDVSsGhc6r
Z1h3Ud2G442UkIhTM6PdeCWzzq9pdWKALF2jLQd/NU50y4anS+Ih5hz4dpLVC7hD
e0lpvI6q3EAUU1g+8uTJqDRDwt8BJYIBLvZ1we/ydbLxhHSf55279E2m7edx5wAY
rr2x/bbmSlHEWZMVKXV21dLKgkCy62FgQHshDnG8IPr6tUlaK99STyxyeO6pqeLG
xDY5sGZaSljEXwqIDRSeInJUJPBSHj82ATejbFNFeXRb0mr/TGkuns3scQ0KbaGo
s8IZ0ru+crwd9lk2bMMHOksEVCrIj12Ucv8SBs3nTGccy4NbI/VHNqLMPN9stH+M
44WaEgaQDcATZfPT9bxPqby1higicUr/1FompXOFF5lDKVKjkxHgHnND2OqxHd2z
Qiwuq+EMMdGtFmPn2N+h788uAJYDui0r/vCjAc6xEest+Ww5D4vxEg4Geso4sGhx
6VWQ9B5PYXKhDtJVI0NpjP3evpfa5Rus7HjPDbAeKrM/s1lpJ7nrT9m8nA+yymIJ
kjf8Rg9Vw26q5GVGb5FtYYsmtb+tFJ/x5JE9DHavcVgtT3INBaFRgiMU9LZ3HR1F
UP6ZnTmNGLPbDgadm2Dkj/8Vz7fVGZksjKHNeYLP10boFUfBDSV82RUZ82H9Amk+
OSzPwplDn6+dUZG9IM3fmSpNmRCQ4e9M9uWOnHJZ2gFzgH8TrgAr3L0KmhKyFhZj
9V6Fy74oT2DMjrfFL6gVNUzvk8vcsdPrNLbWoE8hY/IxA+5r9AgwQ67+oaVP/gAW
iFmnB5VGHeOI/ne5/kl9gBuilB6wVNQS0z7y80SYn6y2ktEedz6dgHneL5yrHR0g
iIpx3sqhlTYODcD5zGnnDwZz6ZMRTMnRJUL2qX8h5iw+2n9kiuH2F2zs1Yfu/bAp
3619OIxYy6f4EVlAq2M2w7VmAgpL43tMBlEfryFXRqVjZVnuza1xBEVwBMsCD6Kw
pg7faTtl475AKRw+IF2SFPEW0ew/HANvtimDsxdGjZz8NHhY6lQsiwhXXkuozoeX
a+4PeRAdD7GjVz9FtFX4XRNjn1lTeiaM9G4BLsJLYyf4C5a0+mb7Eq6w8Wj7btQn
+CzNz2Cqc5B/ESJ2YAQtXhesr8JLwDpTOmswNAspqNPIXpByUzBCqHc/nYIbBAT5
z5Haz6/0Vuhaz/X/T+ECMoKugha9E81yeP6/I8bwQT4Hwsg1uk2HzIABvvaeHX0Q
5LYIVzm/fxs3qy34EZ+OOFUflRFkuzECSnieQ6p1m2GIYFMZ2V0Qc2B6X4qshXle
nGzMeynzhptPbspmJTE6yO9wZTpBZXgasSUF2yjcPzGMoKU9MhRFp4yDKOlkrOcT
HkVIFj/+joFZT7pAJKIKx8VLf/hniOLROd6Rtb7VpTudEsZS404Xo0/i82xTH7/D
kVohNRSS0eYenub8DltjBuvZpQLlu1FXyiqJ7MFQO8jTEzVwtPoN4UDJCTp4fhA4
jo8BOMWVE63po7/Iu8m6F2RxsmGrXvHmJq10WdWprdIcF1NKQiuHdteXDZt91cRT
q+eZL0i0aFsKljMKAtBuYZxiZEP92JuPx+zLxqm9cNiLl6AOMcOkcXDopulOj3Pk
Sdf+JlmVO1ry2EBw/4Lr/U6Ckeysx+Z5ptnJSAIwtAMD+AQtEzZWtDM3CxL9+zEs
+SJshYNXfgiye+cKLXeRu3vUfgQXO6L8AUgooGw3AAOfL0X+klIMbX0JsyWYNSHs
wa+CHFZ0Jsp6c/hqHnk8XKXfjUnoSk/VoUp9784yZueJs2cyPEP8VQVlKz9Cr4Ho
04I3k2SNiU3mdjCOViMAcfZbvwiAj2UIWvOIPRbJVSkS5nfV3fmH8K+C8r6rvi7F
u0Hy3r3+W/knTZ64X/3gL+q1Uy/kiqKFtZTDiJmqDedKHcxOeJIGiZjMgxUIFhLg
8063a4Hk9u6Ke4qHANEFGJiOid86Ji1hLn1sKkDzfL93sqraJHIT7ElVo2nrd/pD
1IWeMU6UQdwuEyFI+IBJuL/DFwvQY3vWZ9RTGJtxla20MJ4L/rNp3tWiivMqVfL3
lannBbY+aKg5V1r9QzcY/kVNH5Tzf8M8HLXfCPstesDiEpDkZH28p88NINnffeSX
MPW/oXd0TG6k3P09fkT/QAPBhRZVhANeqS1rAginiSGdNYdR8rl2dZg0fDOxFUXP
Rh3Hq1Hl6ht5yF53ltd+9C7cYsF5Y8thqbelOepzOhTiZIRfSHwAbKv3r2i55yu4
ch4IAkFpFx9LPHGJ5/floiVG9mCGFy4mnKP5jwfGP98pkG8iVWj6wr6389ja4QKA
Wf5HBAkTXsVM/59ZuhCdoXo4ui8v9yr4VBvbtxyIvA6NuEFk+Kd1vyhTwwHiXaX2
tzeL2/4IxzSoR6VxEUGz/ZfdwPYD2Xcq+LgYcfZ+R5iVuhrsKsThDz6fmpeYt7Z2
ypXA2/UvkRGO3s4IlY7InLCkuuZ+p/n7q1xcLXgWAvi7loL4GoyHQhh/rGHwYStG
jro9JrXFKkX7GUpEpwk6A/F/7NbwWVHJjzdaCVVQe3jwmRrik7krK6qmKkwsjcmp
Usy6TFEYaMDNO9FIQGOvf8orzAm+e0xUVm8YClTu+2D+7QuEk0g6CjViFgHoxs2i
v4o5tt/8VKTm/BUf2UsKoFZz8ivZDL67mNXdBUaCWXZnpDaIhIpuEiHs95Od0gYF
4dLQvp7IXG3tvWVxhjQ2pjW33CZ/qYDT2JX8ViApOuoJAo6OCbchkdqbwb0IdV12
EjL1hAKmO7TQWVoEaDFCbVcmTDOzjmGaPHP4DWLDgIw9dn44DYuFUfgj6CHlCOom
ZZ4sVnXFw9JBdTQX6VUyMRUQtI110QTBlkW4pkxyvY3BLahTEbaTXy2limsjVVEI
SNYLBon5NUQ6BZxPsawq2LoykPrwNFF3/KOfagEefrgVBvTDPib0Z+df7GAfakHg
NElSEezb5kYvqCq08P592ZQ2z0PxMgzfEdnmZ9R4nlh06mNxUov+EF4mxdFyIIMN
o0B8PovMha4ehcJNrC1jmHpdUP8CBMfnmfzlP/8cQhJPWQD1ShhITh1l4DGWLrIv
xXd4oVTqf7qOJscw4dpXZKzPFdH4pZ1QldB2n0ukfRTn9L4aFWxLLsb0h1QFJR5C
kYaQg7YIz/qQM1eTTi1g4AYhKSUY9h4b0uXX6WQCxn4Xiqf140x8ReEt/r34o9Mm
dbH4CQ/J6hkFIF8kuhhxaJzniZuVVmeLCk7IdB5KvAJp0EjnZH7aUiH4FOEAryhf
xAi2JfXeYMjwmGtqNLfCXLtQJGxVYndojxeZ8RkKZQBlhVQfjX0ck8HWJrdLOfdK
koRfNDuiEy9RYaoZ70JtfJoPRbMSDqeAdJPuDvBtmHw2g1WXnOrW+KgRK6AOtgCg
dNSpjVFwtiGh4SbxZ8wE+m2jdm7K9mo+QX3gIgOOmzevzOp+jzZ2Q2WsFzNXITvO
/1qcAiOfywSp7ZkxgRJ4GJtD6swJs+bMdQR5bwiQb8470M966uO+sW3TEzmYD8mj
OV0A/+JMd38zr5y5A4GZkXa9wBzt6Tudk6JyMI9ZyVrGeHHLIRCXCxA6miie9TzD
rVM8xnYLUxLgTcXiaaJASqe6jLnG+hcXq/Z10gfw4oMgl3g4xJtiet0MI1QN/Rw8
ZNh+eRlsNBEwvQMEoyiiqWm4gyMPXcyHMWLKr5KPdN2L/BInlY3pyyqKd1pJMF7j
YUGqON7kj2CFtNB7C2RaVfhMVrrUbY9vBUctCsWIkZqrdwVSD352GtCCZFi1vl/7
E2Hx65HRX4frHVY+vybKViPTb7FrAOrXihcLNFFDtQR+JmqZ9e/WZHRTK6pIXvzQ
3pPRloETy7lFEiHVgoqYWoApAoKssbOMVfo2M3B3qCRwg/+Dcg+wRYV3fuUv74DY
XBykWkzEm7knPoJzIz7CpyFlZXzoDagvh9vcCZ6K7BmieCYSdgMken0dzsblqzPt
MnqzWwoXAYamungjxHQKfE2GI660WqGer8ZxJs0wKKSUsKEr6zEtzwtaIQjUqNyg
NkJ7jR/9RwRqej85u/K2sTXNJI0lKC77fh01Z/6Tx+PJGiwNbTQnScMgR1Q2DUtc
7i6hhpabOwLD9eZ74RvsY/Nzq1wUldFH5TeDr35imqL9W/ar90Q4nx5rxQaLfeH5
RVF1sRO7vi++hMuGtnlyk9YUEqkHf1lUniy75lT/TT5wit96QlkoiDTn7502kHNR
7Sbc8NETy/KHAJGcbRbxlOR+EAnHcCN3pOd1wn9TBrhW0S63lV2oRvm3+NAfnaBy
XOrPcHq5Pvoal0aUzijMmtV5hg9d3DedGDOiuCQLDvnHLcv1Ynh3rwHoAHvw6RAD
XGpr4OzecEAkwJcXhZLKHmvEa45slUFUWF3fhljhYKtHKeoLVCNbnMVSTTIFguIy
VNTRLPj07roH0aqcy72ciZNmm66yPhy8s8iygsLjXKW1Hjf/c7M/aNAWtN9HrVe+
COregnMdB1w32ABUHygEaC7nwJvzcdH+6Hxs/HwBkEenC43KUhOT5gZHZ//IeFhk
cY/MLK3yGZVEFfzXFCtDtzjmMoLc/b1FFABp5negb+qtU+y9h03JKKZV+XazP0f+
4KDT6S5xUwWVuA+tsZqaV6xV9QGYlF8FrG/JuCI9t8CLkyyUnRzotbNTUV7K9NF5
zz2+VZ4AJamX09RndVIYrBIY4qu8Yv6l8ZUyqI4nnFr9zvTm+VmZGxqdhix3DFK/
G+XLG03peHi3s1+tYjwutgffP6eVCF1Owd/IjABWYPm/JO2oVsnqXwc6HMxvNFYR
9OBunIKBf/MXfKkfhFhoW9fqDCU0jgZylSBRTREBePCDff6gq8FlpQnkFKyXNTjy
SY+/cj0DkEfVv7qv0/KpVdBGZGuJUUpxcM2mnDdul0Lyw6jwEhWI8fmDD8gXyo9Y
rxgNeOT5Qry0OQCRaS17Y2DIVnOlKTQy5w3AJhmcfyQKDEXCYN+7tE/8mLEBQLPu
7awfVILEPyvW6XBRqCUmtFRAzN2aCbP6y+9gt0lF7CWxqAm1M4n3dV38HAxozOQm
7lDikFi+BG+cR4LI2sgec4SuFRIFuvQmSzIELk9LDQ4NHYgeU4GgOStCALWA6ULD
+G+Iz7qZCewv/oheTqLUv/8SPWahMn0zNO1ZZsjEz4J055Jk9+mbEJSGE+ZXOxTm
S2uH8lyogv5FiBn83lJ+UB1O+AoiNavVdcPqDoFTlCJGd3XLFnuTjFJfQ30e/5xg
kT7w5cMqgTp2ljXMi1vVg5d/aMB2F7RUDWZHAa652i9O3qyuCZHFWjs46ab7mJHY
YTRZHE+77zYygQ+1JR4nTklS6C0qOHaakYcM1v0VC5NFt0cxC+tscLzq5Ng9hLCo
4j44v4pXjfdMcYTvavh3WsmEd4F3gkh0DMAKiyvTJrBMGxCpNLjQnqs0V8FJSPt1
Gx8U5MumtJktgmMFNVaNXdJLOxvJJKj/DK1B6dxIEuwOeSQvlLluISHPQyKFn2Jh
Kvyg0gFzOeoH6gHTK8mswPZQWvsp+rLOZOydb1Jm1IV0PoPeMSSLv5usDhUP9Qfp
bmEjgl2HeOaREW6sR7TreNqHdCLx04ZxbG8bNLcCts9EFVdmS8EwGs0Xom7R5mvo
TSy0xqgczBHQuWPgJod5oGxz6edJ8QIbb7VyAkGYcpi9y10hpDJVLVKs1PXk91uk
icrSyj45oeiJArBwIIaAA2/bfl4ntquNt+UnddRqVhyI3Op/tZ/BBHB/yWt4cq78
Kd+4W/Vapq2o4LJNjJTWQqOq+QgiiyobICeoZ3/xhrAeRtcp5n8pp4D6pXvkMDjG
HNxvYgKGe5nKoRKbCUJPHTLd8EfqLVvpX49Ls4YXyklump9WTRBRKxGj+oKbfjdN
1QqxUtwkhatJvQ69MpcEuf7ceRkkQe5y61Mwlr0dJ9H6BIJPVsLuXoaJNQSVgYhP
o3xHdCe7rHKeU61t1jkdxiQczeWS/v7+6rQG8JUJh0BiaEn1sHD2AFOax0TBehCA
Ikui0i9ULet5IRQJTCm152//3pkIJiceGvhGWBY77ZLbCTxE4513V5J7Tr5pQz0L
GQSbBZDzGeC77/2yOS02pmnlE2KmCH9KRk/r2ZKMhyr70K0nYyMr9hZTD+DGS3wJ
FonNJ98l5j0RQ0wx/2EogsxFKmMDmHokUa/j3DQ3oFpQlUvxCRPU8n/dNJoe9zgj
mYbK1eBPk5FAbVMJH6HdE4y2IUvQHPrbBdtqmaw6Ogm23ieRh+lRxT2VE8QOD3SH
xXe246CUvqmKOM5jLWEXQGaXq4iWyrtOJ6IfC4MKAF+CsGcx/6IzePrKDS1/Zdhi
mvDV9j2AmtERrHdBHMgP8LCrlPOj6VIDdpfMEWlErLhHFncGBD8mfnHLhvNz28/Z
+h1IiXxH0oY6myyKcVHDWCksh7aS+9Q0xLYvjOeZEmtNiZLJSBc7oScFUOLy2Kh6
2s2SZYiwpwmx7N8jOBEJwf/T2ITzZF1TQeip0dodyURWLbyCPOfozpIiSuRe9v9D
ToJLCbfR8+WdRlu994zHuT5oMaI7yIuMqz4vDz8gvxeDyv/omma59vwYuvTltPTo
OiYBgLphdeY/fri0NENpMpuCUpKkeFjSDYrF7gYeqvP5cP6I3fA4nl+Ed2heiD8V
YvVtyAwmk9Cm1C0n+KGY1gJ7dbAzRTIgDsoSzR3QFu6nmVILPq+7sj5YLHsMhe0/
FeJ3ooDDx1Bk0uncOBCZQrrDk1Tfkv0g6mSZGnNzXbHwuB8dOGYzuorqAHPBwRa3
l429Xd7mYfLLIrula+wDbu25OiRNOKluPNpwQgzuvmWz7FY47O57/j6k3D9d3MA7
9z6N/VfjTzGl8zFHD53Fib86Zlf9x/ck8deIFKtIRqFm3ZzK/Lra/mDtVjbkT1gF
PjEHT63CDy0Bn5HKT+RYEPEHaUfVkQzNCL5bP1aun7hr5ouQmJIOHIhcJfcIUVzU
Za50/uPma5cEJM5afO1wjBoBQgEm8L4bBTWEkQsqVGKDJmbUyPxWBVLxMfaDIOrm
3tX06P7nBiAYiSuhLRG5QKs0KhEiimnTuDMUDq50Bzrsw2p2kKpsgEJnNhsUX0SF
8nnX6FRm5/X0bhhh/jYOmWETGmG7J9ov4DbXGcT2d4vj4/XVY4vRiuPiG0jgn0Xt
kALeKyurwcIm+rDjp6kH6+ikr/1mHI6i+jq1nOXyvuXhGeNYJAKAPG0CRX+QLfbH
OSa8Bf9mmTJPlZgJ2otS3QZ0euDWTDTCG6z7lmmlG+1QZGPakGnJFyeNXUsLhlHm
v+rjgPz3v5T9k2ZXYX0rkfzZanj0GchcWKnTacfK6hluoZKpMry1mt1kyaZnW6JL
NqutLZBTioeD0sRRJJNqI4WQWE5yIwkcx28Hmn+RJbixIQy1Pzz3bkMRXnGKRzHw
dh17lyyNRXXf65Db5QnG4y+69j6vXkUfiJOC7S1FV0QI7S3pJ00yC5E9CMugoxpx
UYbiG6qYtQ1pLf0wbwTIn+t00keDkq3Fm11LxnkMUP0TlxtUjX/9FEnuQdZdxoJW
+z1jkWwX5ya0i2FT4g2liJDJbhtObQZ2oSLKUTLDQtZ9XC1ca5E8ubcNUCIBCMUG
xVzhaVIXlbTBME34j4Y3+ShM5tptwBsYrLb9tD0lFB77ye/uuojPZqMdGiSjxEIa
VNgqVcHGlV18JFlvX11z7e+vmmK8ozdJY1EQzZanKfCimk1IT0BCiqPihCT66XyU
5IJcjzb1XKai+Wh+zSs6Of80dyfTacXxEWzzrMLG3Up/RnI9x3yaz6ybFySVb1KI
84FJyUOCc/+xx1ZENquIYPQNoDARr8GCABfkxjOuQNmMqKLsBoD3emJ9EH+DfZ6i
XqkuihojMDjj0E1TRGNQPB4zMkfelSRuv5IwodETgq9Py9u1o2W5vk3BF6T0eDPs
1VzxcW7WUY6IgDPc4agLnCSL5GKU8NpOCZCjz5dVUmJDdqcRKYdilkdHBblQZ9hN
gaEcyCi3B1qZ7hcJyLidEvd1xzB1lyZ5v8ufUNby1rZUrsTeVyhgUieMBYxfI+ju
+ZXNdZxMTOHOTT1Q1mKqzyUD81a5D9zqKL80OS9F8+ILOxu4EcxcCCuswWP224iu
2HsjXtzWoC3+Qw31kHbgE6e7JxhDJkrmcbnSX7Ja0LbT8pugdArXF9xLJ5t4tqbd
ftyG5TKdf/ygr1w33XaFtgOuFenq81/5nxL1zKDdHzq358V/tyFEdkkE/YsfFNN/
ows1O6HKwyfQuEx93aqzp0IqrHy1kUpV18xJkll0hQ92UKcTZ/ZaqloQQovs7uxx
eJlo1eWqaqv5LuTaXc+m7bC5GRlS8skLRka7V/+jqJODulstuPIixuIpfjDDid1d
/CONwbJ0gdnkWWRp2PljrOZczg7BI9J38vhPqsA+WfjXHGwN23la0Htv1BuBLYRv
DrLlmCEQtE4ZsnecAyM8WqR5ZplNKF/v44O7+YDW29+suaZ33UPxpe2mVKMIFYws
LQGGxRh3aWpBacCqRMRlqwriYZCzSaDVIrV0LRx1hxyzOn7wpM+ReB5y5YAkTcTY
njShy06sDD0xT7i0gOwXYkuShiBERbsfRh7o4vdgdPqA3tOxt7yMJCEcy1nGM+sF
yZBtP6Jvncgf7dexZeVfCGyJmaMKMaLzvrw6jsBOg8C6KNyTrWIk1maIgDaarFYJ
4++/y1eNwvBPQ9yTRmtHPFDC+dnmAZbR3BMr1fesdlG++UIQ+09E1XQGa6B2AY/6
jdilc3eNMZkwi/AwW8Q3/AadtOrUe7Cb6TO2KVud+FDkZAg7KNbyWtFTcpIwXXiG
7n8NE2QtjdncoUzXquR97e1ZubW2ATZukdJ5N2lFcG+7B2JMMZQ/b5NqE5kvmKei
TtPU10a10i07qAigqX+W3WLj/iNCCT3EkpQuEg2Qh1FXfWddzziUeG+yTsZErk3D
6qiP4rZERtyPbeyDqVlcyxtww/2sRzJ40f6a2yXbqryhvFyiqmO6sE9Stbc1j5Vu
ueprweyTJkmwcLQLRHWcN2O79x45pKZBTKsJgM6Fv+95cV2mvnQFh3W3C5gwAfUv
oJmcHbjSEPdWdGE9FkAsy32yaWgHAWIuPd5szC/0YzGjmYnyb88hVBZRUSUzuk5R
z8Z0TNz5/ng+yEJoMB4rsevONeQZmylJEvdacGrJ9+oJblxUIM34si0uLVcKugJh
qiL15tqd6VZMukNmJ6EKr9721xTHCATirXYgw/iv1MkxYWFE+WLseIpBzEpsNuk2
nNne6IUS0q94nW2FbI6af6i3sSS0HjFX008hYV5dFwaU98VGgthyD1spTfGvEmxj
DxjGuw/RyIacwfm8cyouzqbXnmgBqWK5mp+4OesMnkNwHNU3LMFy85G04/uaVeSX
SUbu6GGM1GkapqQeyoQjrAW4SOhUhNR8aVB8+YCRJCDw+WQgGTJe2FFimEaTuuFL
QkifHLghVyB53IoAWBBa4rQtw1cS3U02vJ0Z7Z8Huwshtzt3IoOkWt0A+Addh2bg
zPo42ivFucv/hRbthKFF+Ts+HY0gfQQzvGWhj8I3Ctzuko/HY4aRUy3yJDXZ4zKG
f3morX0Mpz6XvX9d5D2kAiiKCny1c+8uku6kIwCrDmCvDroCo9BNprdz3at5dKeX
IIQI5xWSnN3Zl07tL1O8qX21EbaYknIthOLRcItnoz8xd/mTL+qXxjho+Asa58iN
nEnkr4VrVYx1KNYxLyLBftRrxroy1o9NH8A/UEZzlymy8GtNkoIPm1cm8CvRLrO/
0aJenqxn9UeNuWcxyKEhRGvDgNt83KHugLjFTQ0W8JLxxpjM6EGaIHpcAygWrnON
bZe7jDSIjIKK6qyt1ZMxua4TIZWcbVXCzsJLyvOe92dYfwFUyFkxI+Q3EBw6h8w9
lhCU7Qo7XqrkhTJ4UKAD+xzsDkBFF3sGftrknQt9JXBZGMV7C7WWV0hxQs1Mip1h
xaj9qgwThvxbQyTZb1JQXIXkKm8ZtOEVSZZEa/MrfTws37H1za6v0CxZlc5Vo0A/
GGMdjRaEXk5JaNyoP1txSqnGwIV0t92KRa+fvF0sfUSXR5Eq/hkmXj3/1u95LmQF
5C+eF2BKKCsH6mmiGq5P9luF5lOXbOYFw1DdkNBZjPCImgsJE6h54W3j+QLpEcZJ
j8bWU++NBIKhYeazf39ZsrIHpjZhsHkKWk35frYU+HmZrI+n1ICiCT7RDXyd0t3v
F3lEoRaqOHBx7xub5U8jaqLFr8V33oZGTLL+8PqTc48aaeS3TFqrRi4XNGhDHzPn
p2yoFrpSV8Ypho57uy/AFukQGnaGtLklaJa78t7nP4SdhuYAepkBkXUVg4iJTf6D
S4G6Wmwmh0nTA5pospOFJsiWNuRKKE2wG84qIFXCKdv4465TgSebAHBRB/L72Axf
Ln0xlTNg+44OALj6jSF2Eiok4pYHpV/Wbr+kpAUnW+iN52E6FUC/xP+GALi82TGJ
/jNn1j/egKj5ZwxGoINaJ0Y55FRCI8G9RoJCAJRdz/ou/QsxYMTv6P85rRoqFkx3
Cp+n4BBpZ3mW7CQb2X5NcVzNJwWQ59AoWgrHuKlhlBRs90g6n9i+pc6w7EF3nakK
+VSE49Ck6GjbnTqHgEG+VsyjE2PFva5Nm9IdQY308qsvO4gra4Q4pS8tdLUbVwu9
2gZ39pjFlxJDERgVkQpa2qnN3ncfHNTxlajqOOTpggG6vZkpgpKtQ6XiR81InoWA
DoumbneMSYh29wyBvvKq371E71IhLe8H4Cif7eEY4/uL4iK0Nd2PRbrk6KP7OxFb
+QRgfQVL9DGADQv/80bGwJa3gQSI3p7OP9kJEtTYep+P5lPAU3uYIe5kzfYy1gVG
joaeIDIPKZHahXM8Y1gT94IYeVb31weWvrfcTaSkhKKp9CPA1AnzV3ruTGHj5Z9r
HbQqLh2BbFAf9zdruf65VuqHLwvRAB/8E65au5OAKHK0CrAAgjpEty1J/yyYSG9q
ZyYT0ef4uqlVXhAmSl3Wqx5GhUs0ZuEmD+HFkkqfZfO+JM+0B5JKqU9QGCcG4MQS
UQTQu8IXDgrT1QbhCioaqSWeqqIgjarlfsK6eaZXfD3wADzmbC4loBzflxsdfPJG
8C+Ju562QnmDakTZHOhI7ratnduwcUEWiesC/De73cq/wplKDpH9Lc+1PNhztXSV
u1tWyyuDiENeLf+Nn4/+ueZpa2rtHKYClhFagMdh2cpBpkviAEd+Fiyl56cG3M3p
FsYyhEWO2LvByQKCnhfB4KRjPS+hCu1b5PWaIOoFtBhzT+EPIhiqGY10rHnHZHpq
cmN9huFAHUUxwMIbH4bdy5fP0AWI1o7mGSlslEa8bRPMB0ntVv93pwS7L6iXcuZY
2lZ3UlBXX5nWwuPJ0849MVqt5Bg/zcL19FxArTpeB12cvS66ygWRrC9NAR1FGBQe
LWhrIpWXVpKkg8tgw/DeTund20U1Cm+cycKDFvU/c4MnpV36Kaau5QqTmH8m5RVL
5uS26vXrbzeP9GA6y7YukN6r60zxavB4539YAtpe8RUzsPZRMpWlEQX3+aoyf5VO
wIRJZLyWMF/JFAKxsu1Dax4dCcJ2f90WDpogc+s6JSftq5hZfVf+w/kT6tZfUEjs
KssOPxCZdAUEZohq2GTsHISz0rgon6/jESNm0hZNxWI0MhmZ7Z+di/u5OrKCeKi+
OwdngRKSC2wEURmxy6oRswXT6jjZISrsJURoc3LzmFvy3ZJAPIN4n6BIf3vamKtH
BNP/M4LBQThJ2Z4htARxz2O28lxF3VY3v1uY/0vs7Yth1ugcIHyVKTy71UTLH3Fe
EO7dFrGNmNCxEWJ68kVYNksxr8PvhWbcN71lRT7/VjElD/AbAJMopZJVQrLxWYEZ
GYgAs4nb/rcnf+zzqHiunKEzt1rZo562FrKMBmU18wkzyvAFMu/iS/Q2zK/OKsiZ
yGPGNSQhaomani6hmJCCdYb2N9JL5Gxr+XHVgrQzY1JpJgNCp+XR/Kd6rQQIUl7K
+kjj9bPlBRjUbLS204h56GGNYWaf9HQ4oDoWt+3lPVjf9geP4pfsMDBVDU0s1ir6
eM9wDitrEEE9sQXYe8I3fFtGUTzd/IhTOca7st5xOWqo2EAtIWxGqBssyNKpq0z0
tSbsvYWHya0/MGnn7XdnIhqwhFQ4c6w8KsQoTvNm0LxHf1x0sS/OGE9rvLxIigtw
C0YrnFwtRvQBQiaUwltEu3O6HLf1SI2/TykdvAf4dBGUSwDhz+U5++HF/GuHxcc0
tXVJkO37A8svQxxK7RyHuLvp0YYNZHBVdJQ+MAStQSmq1RADKzVMChrqRxmk5rn2
gPUmvcUImQVdYwQWuzuYgn+wcvY+bRJCineDGtNCkQQBqktvtQ/TRNIsJ32qYTIm
prY7ASPZ91tqSbTaYrxEOG0DSk8lXyZvBZoYeZA+SKcYqhVwUa7xp04uzi0bXG1C
xwdiCcHT1hMiIdmFmKKx7EIsv7O8mZeCHZih9d6HCEcBDPKZB9p2k1BbmEg4fWEJ
sYW3NLM/PsR1xEg2lMPZulWq+Ct2V3Mk2Q9iJxCkmxvFbplixbo/XbmVMLH19ETB
RVHwjqvSudrK9he7UbhZA9hkWiH684LI3L97fYkNOx8dkiLZvTtgm/kig/rEOxhF
rneTFU585+OjV/+d6DggxiVdhAgHM8oNOnHHHRyrm/pwNZlb/gxavkG68FEnIxeW
O88x9JYxth/Mc5cFVE++i7kI7elCVw18mzX5P6IO/rvoNzzqkx144mVxuVOPqpf6
kh4L3wuBVlTBgecj8fUTMpaBXbztYA/PvxlyJ24YZVTWG8+Rf3uiKuJPpoiUF0Ao
MiKt5DwQ4U+xTCxkAuO7kjdiT2uTCI+64VL88KmvtaquIDf6UxailgfPtwPMOlA1
JoYL4o/Fy9AFMt6oGuWX19Z2t//YknPapEAehZ0bWwkLXo71QDZ3CjyyzbdbYb+I
wLM91ipFKNLaSwQJBNXx5p4J3qaMWTAaBMk51/yS+aWn42eltlXzhItNuZ3QB6AK
vp2l4jwKrBvs9fpFOiOQ3pkXpE3twArmabqMpG7tjPvT2AFvYW8FJTpWEL38mouH
hjr1xNyUzYgOoAQA4PPj0E2j1K2yM0kwRoW8QEVEGGWXyCAau2jUfQGm6W/PF9zk
IqU5tfCD3z1+FyKPWSBGbJclQlclBFVA40O0iqoS9lpxYhoECHZwHyNFSbih4BrM
OiAmr88S2VWpPL6IFSvPosfi12+pPJUPokK9ePdLT7vvfheocm7fpYcXfEN6CauL
RL1HeXxFHlvKNVTrrfRxcsF3x+YCjWVSdy0zYfOG5pfDTIGthXFMyenPItncbdoK
MAkAn8//0iKz4IJURKd62UXQ/Ar7KwkHZ+Ta/P06zhbTlkFpZWaCm9EZkojoSqLz
+stTaa16syPqzOToLp8LT2XBenj/i0WdT/eH5b9Ph+zBf7sZf94WkwxK46V8G8vd
bjWKjo+W/tf683pNbOZaIDvhPRylix6ZTdXJAsF318OX5kkfnC9x3+NS0Tcv0jCW
F9Uvk8zYslpcNHfNPTiT0xn23x27YCs/oxIrKi1YZEg3WmuRdv5loaTo7cXG0Ftu
C6jGHRp8Uw4FUbvbITjIj2u0C7bweI9OzsWQDkB3JrOhEVi5WxTwTQqUyClAw89J
5QHKYnFSt1y83Lqavt2nuE/stUP3VXNF6jtAN0HNtqepPzA03w4Toq8ATHV2APbl
5agdNWatVyWoDh+OLNsxBqabqx6sTbIsKeOJvFFQRk3UsMKCxvTfqpWL/Y8keOG6
1OymVXBfhT4c493tjuB1SEs4pIQMHWNLQvFtO6ww+l6dCRSFvlBdeUez7CdVblyH
nRrWbyeD++YlrtnKnQaP5go4joMGo/wi2/FRb/uSSgxNJqbqymiwDNFQta/IW9YF
kt/QkXJG1rXGu4I4KCb7xqATEmzdaaEBaJ7//Hstph+k4VKhLzsY5DRR34Hp7vKe
b8ob5Zy5fs0AZqdN2hrQ/4A8DJ6lYKC/d4vqeJf49Q5y2dvKLDsdhJ1YcGkdvgTr
K3I2p6Eot2Ff1q0I4cmL7S4D0ZdpJwjuf5rLDn7HEuhs8TIMemvZtOkrmwv+vkys
7ytRcO1hebAICqvqspa0v+gtiL5W94DxLdlocXelh6w66unSIO231URcR3nwxK6I

`pragma protect end_protected
