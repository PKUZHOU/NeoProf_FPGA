// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
QuviYtKT5KXQQYmz8GophQVe8LHD0JFZyVa+MsJlKOJ9Bel8296r3nCVS3zk2U4T
pQ+o6BFL6Tib2lzUn5SZz6vQKPIWUqBhM+ySEWw5z5bF1XRuMxU4N2utYULL0j0T
TV4JeyYEA3V/J2J9crGtgpePCDuRu1dgob/KOwH0qyI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 3120 )
`pragma protect data_block
44eliDaH/5gdZJeVPeNnAU2DZQAyTdF1cb2kbbyW4RnXrYKbgqeeTIGCYCQbVYAj
Wh+7bz0246zvWv4DGtN04MXZqRxF/Dpy03Z2GYLTiVNVdVpYykyFxjf/A9dDqSKk
Hv0iSnfKiJqlZcPWEaeLsy9Zk/myIIG8IbojW9tms/CN6arGOUNU+KbSXTQQ7stn
3GfYpdPfe7eJwdBue3J4r49A41m2WWnEVN9BDqrCZNf/+umcKd9jg9KRIXOzo255
8kVhVik52lYNx2PT/RpiiW0uz4SXJO4FkcEmEqKffJD+8XCwKENHs3neIexZmNRo
jQH/K4Rh70dH+2xTUVj7Rib1glZhNLD+F6AT532CHO613K83oLy+a2ZzKEGd40w+
aX/iqyM1e1ddDK2Bd790P4C4ZqLyA1qq3SZrxorQ27AD59+moj8AgtIzehrak8MI
tjOoqe22NG1q7mk3Qpk9zHyejfwvnegLT4l/y5ixZ4AwnGOGhDH1UQ5PC1jFWUpM
+s8CXajK02vr4weTlxvy9mEtoa6iF+DruPK+9o1+X1kF/+0utArg835DEtwle7yU
oIp52v3qp3ib/GjwmYLfxgCgNoe3TSHTU+HTnxjiBtZwj0YqPoCPVO0COucXNf0g
EbZrxk10LhPsZHKxz7nr8c4F6/U3546vQgEtNpwdQ3XW1VBrVlpU17Wy19PK6EAf
tRrbroXSB+R7ncg9B/YpYECYI6Wn4W4y3TlZz0XGDsL6OckypzfmBatch0WGIe+j
nZHSz9n4oJd57+pZ+VKAg+ha+AjdUcSlHHkgeI8z9JxwEhbAcYxnvYB/7SeaVJXW
rRh8xSFmUB9MCbc8BwshS3PffG3K9+bvhONIzKMaixtc+FZy58ErSMKFEH6pCoWf
Rkfwee+/5V0zygb34w6YG4a22C1hfuuPGox36OqyezK9UxIjr0ezrv91DaznEE0Q
DB7GXj5pXn9CMaSOD3vKFQCWEU4aqi/ggs1aTCCDODMJ56GhflqZwnQnL0KSyAMw
nmqqaLMQeqq+4XC1Ealr24d1zTM9mbqM9+6mAYg2mQFPCRb028U3R+RhRdrOG9NE
Vh9PxsEOmFkFeWKEqAzoEH+6/fDpWLan56wVSeznK63Jd+FPwYLCykI4+ke/UWR5
3lVRsiRXSzibJfuD7r6PBIw6dhxQF0lr19MIQMqxg3qXQcXm3yI2KuN0sApHlpul
JS1wgCknNNhTTLLhTGlzt7h6cxhwkcSj4NfVPZP1qk1/YtKCoZ3e/5g7Sq5FDuCL
bY5Qoo+cr9gb8qB5IkyPuegDliYBQVTKM+fLCpeWda6/EiHcCVBAcOrE87CHV3F1
f+dhSoijX8VvEat6lmKDJzmlABu7ZP2CaXTTEAPQylcXiBzep/q76l2EA1r8IKnO
dIwPfMmDRf+pjBCNm0HMXKT37t2xsBmHfkh/gX3ran6LMhwMu3H9zUEiMQAiwUop
HQbXIewST4STULF2oXbGyKft5k4N4wAhsXIpy1RXUDQbnXhd90ku9mlWTt8Ppg15
ii7Rr/0Htc1OeiqwnDfLn9h28koIJcgNC/ndRExnrQUnR0kwaZn4CdI5rBnJYWok
VwV8EOQPDq4CbAmv+yc0V6ziFLYNIE37u0pl8D00D8cItGMqDQQvwA3jyv+JzRdw
CSKoC2ORtRmk/ox/Fceubxe7L/hIq9Kin91qe0mOTv9HtWaGjUuhH+HbNswauqda
L8m7kd5DdvLQuFRKkvRVDvG/oQc0DZhbwKHsSDmBPbq2WTErnJID9lzRLT7t4+v+
gP3il3FWmEHnbuuISY8o53WSRe//d1+U+ovuWXJVjgE8003cHMwwMNA4MAYfrZh8
H+9VfXH0xghY2SOFn86WXvWPS5d8SxqQA7Rrh/pxm+p2vdHgN4FS1+efW8LAaDpM
CctHF5akXPLTP/GnzOSViwsjlf7L5A9MPZNpttOARZs6MZcwMbqn6L28iX6fIaKG
gABhdR1uWZ7k1ckwz5r7FyGeYzEgx2jxejk9TJL5FgxAAkvgtGbdmu+GVYeo3ChT
YQOcT3YQGlka6ao/ZSsu0OOdI9I6d1iQldt5FEkr+ktM0Th1GCfGDAr2ele0rHZ+
/qBlL8XUjaVTNXwOGfrwgqi5o0LTeF3k9AF5GGrn2ZhGd44I3IPZ0F4WBgHS9dEe
aJvMfUOHByvRjdWKHwNeiXahzQZKpiuXfmRqksSMcpBMjCKCXua1MOxOStY9XNto
qMXRX48DgBaHWuVaZYdrfLxnhepjL5yjB+7NwBeAGGeCf/e/01vXtHLe/iJlW3Qn
iQeDP2KAjfs19PgECJX9RBmazXka6PEV0MZjrCCVtsBc3E/J0yjoDeGvHz6V+rV8
jeqPEJoqhKqBaGIBZad1pCt+GYbGLPXEgUDPt4YMhQZWfbKFzfKCkpEsCB09BTlh
AarPUWmOh6ec/9YwQacWM+AS63UliKtMn8mH1r7LBIfksm63Uu7rqw2JAkmNgrUA
K/h74iY4IwWBU61kDu5ynmxHKSj+rcbOtmvj6bvUZjbdHyd9IeLF92QTI7XPQRtx
+AB8rgD4oiHwzRuwYN/Dlg8SLu72RxVcnr6OS6VChjoeNXvxxCNfw+Fp23ZcsQkR
sfwsDfbRRw/hyrdtD5EuKUYkWOgLXlhQXqYuEQ5JXIzC6C2cAFH9ZNm3n9qCFQBV
xLgdZTW4GAGOKzawtnqIZNp6qwJkQqIHJcWf/whYcF//uKwKo1psiQCX12hHoCrB
XlqS6kYVMxZtrxKlaNHRPabnbCT83zRtjfOFLlAsTwjRbk6UvXEk5hwECfArcx7B
zXLeOw0TqjctZioPuDQIRP3thJ9ZFm7mpyNZwHDrhDmNn1Kxhg2Y5c5k9nJ4H3eC
SLdsIY6PoeqwVo2SJsmJ0dUD1xJOVBeuksg40SCply1YldAPB/ORBASpoSo9GmnD
YJEs5VJ5+CVTAPVyj9IMuSAAr8Maf6AZzC7W1ym4MktMRsrUatqqnluuS4Blapn/
c0CfQ1i0G9VuuPcX8403u+D/6RGHFq/YXHHuEvj/2QG0KkOTq+yBsauYUpAxfdRL
oCA2s0iYwZakKvXU6f61oaAGYAId58YlJL0fc/0ltQtSr3NYBcWOsuuLsYwGYF4F
4GxN7mg8HRPVgdDgvvAYl5BtckP8V+eRHV9Mu1EXAmqKeal/WNMYIqE2arnZckD8
0ixBoB0Lwrrf3y6E00sQN1Uy49XfVcvuFNNpkI6g/Dr0+y/6FNUqvLcJK15KdNxu
EPHLNPQSWypv4dOoOvQYqGBN38trHX7ftT+OrEi96ernrEa2f733zOZNi6mEOycY
oMKZsnwmnBc/pc7q5l0MFULA3C0J7BBMrGvJ4fMrB103IMtV1DURd/Iavs1SyfJW
teRfy9hqoaXOInD/6KMh1GqtxTcnsQWbp2w+aDoCrwOrPpQPHr/FyiluoA/dMi4v
xsXZfeKqDEo+xqX4lvhACbtva6Aoz88fmCHqbzHjHmIzWoY7/zlLoxGEJmkfU1Yd
hOKPwpSBQHoYTXkIj8o48JI4rh0dGCfENLQMKk1y2eqc3KLPpkjlid9NiyUFvgBB
iNNtTx6XznENvyQqZONoGrGyaaTp3ZZtL8Cvl03ibqXHh5tmfZ0pVf58d051sC6t
cChkMQXmKGhm+tJrhImSG7rwjt66nwuvjuxuHUkfTgHWPytdHmqMf774Zk8tq/na
oWMUfSi2NYMdpH+UX323pFD26oPOUJ7SvXZB9snhIw3zOaIOq9LMyZmFgJm0y4hC
X72rirUUa4i7+eGX0WXiMqkZqR+zlSXA/AodV6wM4JhCwswQKHZ2n5kIr3dm6/7C
3cLdH+S0mdC6Fg+GKB/W2nf6lSYf3MCjvybrf+ZL1bK8gn7YrTo0L0EtVlJtglMG
4x7jhMTdzKHURYsZngmX1TaURvROyZdFJVL2AENy0YQPQ6ZYww3tA6DBd3S5pruk
2EE/jkJbtOyJxxKbZYDDlcwPLZ2cjt9CG6aPNzWRJVW46yciLVvHLfJRGVcTJj2O
cCYXDCO3ngfkgNuT1Fiu00pihG5gY6mwyc9DlLb8KmC9Em/RHt+9E7Jb0MmCvGen
g8QUQEEgonnm4/3ojcZMIlPa9W2/vB5caQgeUHH5zd2/QDCzHlSmqHj0zVbWUwQO

`pragma protect end_protected
