`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
jHz5zcqeK3t2+Mvrad3LIVcmlsEqwlnkt6hmCbB1vFpCsesPGPw4Y/ELE4sojqhM
h07tZkPlYmFVNfi7FXjMAPthDyv/stklJfXo/3rvlLEo14m+Vh3iXIhlt+vBcFCE
BfEqc1EUJh4v3W/4TqFl/e3zNquNK4/Kjig42si6KiE=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8544), data_block
yix7mU2x6v7fV/wkDxtif0IkkVgWD0xOqdgFw1OnEc3AMW20kXiPchvrzY5gEGXQ
rXvyRlDRAJY+c7kF5+eiA4TSxz2Fzty0S+vhg/oiAUp+gbpjuvxGjqfwXYTEEaJI
9Zhyxyzea/Sfjv+P4Vl8Of0ZKfcgFxhmmlxaNtMZ0DUer/+Z588/KnHrrWRkv9ws
CoWC4UWRgTiB1TxKeXGPdyPM40rFCumR8bIC+TpnTgyiAbpiGA+PEyiZmO1sG/59
5nxzKy7914PxxHEHBfg12B1vvp1vH/3/4uYvG+aU/utKFLFoi/0hy4pzNcT28fPL
hCituILWkMoUPw59vzfrRPfX4uDHu7g+CNzPicwMHKgeSZMkeXukZCmEYT2BX8y/
8prDfOX2uNeXaEAfKHg9NZPDE4KX/5LQG5oR5wpxDRVpHHgWcUr5MmJl7WyJ8+E2
rHO7qudUGoMYJP+gTNEi5H98UtH33hN9rmWI7FWxWLLZTuPeUEXh5DqXlE5xLTm+
kKavxuMloEuqLEN1oN3D4lNB0OzzVSNwskDMaGKhsmZgxu1uNDgSKOMC96XASsRP
V+peLN66PJGfao4xM4R90BsA8L8ERKsathrDX/93Q1/X5jtxXtmlTN51+Mx01mwz
EeG+jOEunoLlYSzaCeXQ6IUne1YrNbPjJC7bpWoCF64UZp3Vbuybo2G7QfH9bcTb
z0tDj3qnDFEdA7e+aG3PI6wEJYwsD+HITeDFGMmVxn+ym089lBmVOpF9WwQ/HR2V
VW5W4U1Yf0Hf6TksRMal7QhKD5h9wZKpaiL64kp4CFLL0I05Mc9tMA30eKrph+so
yooRY0DRIVZGyRu5vHdrr5jz2Nyq2GJg3jnwfthvJmsorJWKTRsC3r5/9H9BLP7s
bCKjJaDlRbynxR1H6TjrRkCA3//iZeqeewdy/0FbZohIdMU3rypv+aZpp9B2Ptie
IOiEfpyyUx9N5kL5f6L3wkXwhB4m0eJsY3gYiNGUYu03TdqyF0J/6GSfXsZmpmfS
McAtHyVu1nOTmPXxuGji2jzzHvUxtYxzMUiRfa/7G/JhL+greEAMSB2t+NOWFDT2
w7ppBbWIajVA5Hzd0GLHBz4/lehws+f2RLqMbp4eGxwPQrNws4/LkNc6l6vOZVFL
WYOG6dD2h99WlUFOLX9yrANLBCN5p0q1qOAnUiXXZjtt47f0GclJRKFB5OxdAj2H
2m/Np5vr65DCoY7MySLMMtOW+rxUSibbxK2X3qAGEevawVPgUutf+F6UHmDj3v+Y
uHROzsZUHOu3NJd7vbhKk3gaigR9fHdrrgUj9XCMqqZRfPLmXMl/EFj/sIxB1+A/
wVWk9wCEiFwuWQGGovuNvCnQ+SOGSGHc8eAF9xF2e5b/Irg32iZ6LcF3i31Hlg3U
1a0oIRz58AlLldIangNF+e9VbEtdpVz3pxmxLkH1upoiGCYjBMBXAZSBrM6unVXQ
ptPClEcEOeEGaD+7BKqQTS368azJWAXkV4fGxqFvFf8e2QT2zuXeVUkZUI9UiiCF
7TptET/aqN0ab1o2R8ddm5UcVcm0sxdnipFcQTnxn3b5oRxSNe9umObi0coP3n9L
SruWJUmE8xmG3M52lwGClfDlb1Brxsj8Pr2oN2/jw5FHMnCmZ4lM8XfZA8+iFJHf
of3BVUV153yyVEUBGUg72h1FKJL9cc4QzEEFghOltKR2LHU2zExL1Xa4YQFVW3Ha
Fb0+w+SEACWdiWjmFBVtGNHMW4C0ANFsNDgy+d0l28sVB6ZexAJv5pLDD6wqG8ij
oNliONKnpEuw0v4KW0LnyI465tTsBythei/Jur0lqjzqWiakkiqTPOYap4jScfhM
/+BTqdlyZnneEset5bW3QvYmN6cvXAjJdeCMKM606TUMynbWBzU3sAyq3kVva1Td
8Y+uDyLbK8AZnRQNQ6/lL0uWSF6eS+JZKUUpSYmQeMU59GetpARx+hBcKN2Wb8Jl
gm2Wh5gA2qj1PouTkEdXYvllHVKQAS8mNrzvNHzbmFUJ8A1kvXkw+VugRwtr4hqg
9qhM3uMTgHrWcxXluhBoV1ZbLOM/wxTV9dRx1J2pDh8RQFFb0/kqmBwnfUpcPoqB
pLHeNd166eAKqxsjZZC49qiVBQ+kva/oEAJeaNeoB21Yv1KPTr55aHQGyLp7Ks6A
eWyyT/sTpujLhS6Q4mqa/hQVSCQBEp9MbWESskN0h+OO2hNO6OU3FeC2Ey3Gz0+Y
Q6mELna5CcNjxbTpQtRapZMsNRgE60QxeQnXY9ih77IHQlPeBuQuWp4rHYxgKbIs
lOPBHzD02ynwiCpXG29/hmMC2tBbQruWaR4xmmW7tnHTCa94WAmafhjwfVx8pLny
Vh4lumbrTNmKnhcNGkZEcBLrBMMIJIqmwufZSWRkUGy/kYVrMsavtMpHPQ40M71k
QKH9ADJ4rDPGLwddW8EXLabl0Jm30QQHln+nnDPiBjjGY76sv7H8JQ8K3/+as2Lf
AYcGYd7qASevztt41qRezfceeh1WhOhoIVHtXGxXZjf8z++vhVqi8RmDldOHOlVn
HaZrW83WzoueKGbio3z/V+Nyzu3C6T6g/KoUV7PIyzMFHpThY5DsMF/hptX5zrhO
nHTA1magm9wQUiwO7O3hIXbimpTClDVFo6D4lTSUppufnlH4Hrjr8Hcmj0Y/vGwf
CZB29vrX7bWaKlawLR1KgtoyDpHc8Me3V3xAHHp1uh8gbrrpTGikeW9ct7raR4Ll
A/cPWirT7Rg2xR8hCnV9TEke7oJ8ra7Vk7730s2yjQjsFmPxPUh71YwXAkYfWhSU
IyuutR44xDMipzUtWtzAE7ZH9DF6mhUV3iaHucjelqVPX6MdqdIxpxAKBSCmpLp7
TDu78gawm5EbIV7iC5xWIQm6h4Ct772gsdZbSF6UPduATXkgx0CZY7HX9Xcv/mo5
nZOVE80uINsG1hTmy7DSQ3BaEZy7Ol/ivujBLBH6cRJPoQhiEdluKqi5HKG83jGP
A5+sF1jRepaJa97/kD69ksoCTXDRbmfMeGFKHrE5qukV+eAsfHX44B55tCA6iOYq
dqso21fysc7NMjATSi0qV9gukNpu3rKry+p2xMURXrXBvPsq3uMTyOhDqkmlh4Wv
xEnEwqZ0NwgHkcHY3Tadgn85kteNuJ5NLXT+n2W7RBvwzxNfoTjZEm0EcVPxRgK2
VsPbgjzDhU9MYmvtxIfVhalxb2vo3kCimlLoRrngog6n80rnZpvjjajK/KjFLppc
8bxdFQacNTUR4j6ZeQsMrUNv/JQziIimL59/s4O2a/BRdbFXI/fjyyuf9TNEt+t7
OUUVm+GPocfHsoQdGX6LrxLnEipsNiPzSpeGZAB9H3fC+izQmWsKXs8p8D5RMJpv
C1EHYG6Jax6FAWFGoLiftMY9ERvn4obLTGFvdJCuX0CGOSShAc8D8FQZsv4KGX7I
m194GjWxeC8qrLPZId7SxCqAfq2PYazVK9wUAxgxclAVR45IoUnDzXn7/QAZ2jLo
wQYGCTameaiBnY5mHU6brkJgZqcVtSLuhaWg2OrALx8eqOwibdTY3mfeZAsvTiO4
sjvxIveNGCidhILx5DNZq/V0LDNFQ8t7QLYpdPNRGqrWsbs3zh9cwNMCUe4AfQrE
Ee4SqnE1mfGy5Qu9+6X4NsxRHBsWO0M/OjNxCcQ+eZAl8Rr9YRlayO1U69z3H5Ng
Fg+4woyC7ZwDhxn99Qh6/+69K8EbpU3kUc2mkmrHPc0HVz/Oe6bstLv4P/oHtBiq
w2hOqifIQEzcbjWYSwfHp8m4kDoXTE37jwJ6fHtP4D7W0EcfoHT1hhxkt2pE+xB/
NhaUXxK/+/5nawzhYlRaV2q9+ZmDo9jdy2WROBPJW4SWDnLQrlYDF4p+cQKxdV4p
dK5xwxvv+sdzhVXK++mxbsv+RJ0mZgLhMqojxvYBErh5SsJrt19GxdsG9Jo+6j+0
5TaIi2BzYFF8iNNIGk91W4wdhAJvbHGkQflfaSwaB6aOrDPInsGWQ66MEcvOW6Rk
QH4NKAOmq9wa3gJ/DcmD6rBTby2uGbD/WDVMZ1OM3Uk477t15C4m4UCoRDdUbzFb
pVrSroAD3Jw0V7vv8gsf0WMoE10Vmrde54/FwacvI04bplyNR6jdzirXl/nKNb8G
yvcBqHiGgmSl82Nt6c7CijRUCSCyqyBaDpVUU2O0ZOBHDcPu4QTK3/7pkEDBlb2+
Y0NBpflRu7T6XCXzpMp6zyA4j6bWOSxrzDj0zxzEDPnws30dDizgH7GDnntb1kKK
QHcmTh6CGiYl5hF5VYejaelLjajCOi3eFCNeEv+Rk6cdxuQ0Npabob5tSnj8iXdH
OE1j98yAYBYNr1txb7r104/XjI+GqSiTKF6leaUr00VZudUvwp548O/8HyMZ540s
9+rTFWfECpXTcJMlmMTeIWKEvrOcW25MXCZXnZ0m9EoZtkbiM07rlcwcZer8/Vpj
NoM5y4AWkOc35taoJk97LBPcoaHbf+Gvv2SrdJhEbX0HGBT6yv/Lc3ooefvt8iKo
6XuGB4jYVPv5dj80C6mCCjA38xrUVh/wJu8ZyHf6ZZLu0dzG3YgRTBy53+f32kkj
vskUn6x6uugcvP54DYATmErahzvOAuL+L2sbut5E7xkcps22Lj2ATixUPZA297UD
xmAcDVlZtTQYRsRVtarJTc97TOnV6wMLxuFkTS9hRw/iK8x6Y2PSkKh9fU2HLBBE
3NFsWJNTNvGujU/ehMqqR3jcV8KhSr0+GIRjQgd3U2bR6hW51N68Cm88NwOujTge
CYOUpJ5XWiVLBemIZ51LYCajT028673kOTbHviJSB0XTq+k1D3+PpJtbXDms2L3z
ehO8yVOtwh9/zabCnpPqWqLWDcUFQ3YcRlncBMQX3rFJb8uVpxQoLMG30uf2O+hL
qmYaNr72K1gLK/U+SBLeq+Dv5c1+ffljfjyzOzL25rVS81HoZAYro3cn43wQHEYX
tGIXv0AGE1f2dOJkg6nc15OThnysBwTN1Eqkv4ftF9RWeKAwOQH90CGTYbV/LF7X
5f/mD6hD9CkSm9C9+4HrXtu5lZ7Mf+0eKCddzF82WUYwLkWV6uXdUYMxDCOe3Bvk
iVz2TuSZ6pkkPc/DgyIfHL3v1VopnDgdj/p3qq9kMaDbknNZ7xUHoa3qnrt2AA6x
vZ+10exoTDqNZmE/B5P/ApxLm4oelcdo7YyHtRVvqfZISZ5w6FnFJ/eAhhd8Ls/1
FuJzA8vlHXCOH77vteAk+Ny3S9kGMB/hPZ3//cxvr0gkVl438VOKWJhB756BzEOj
AXQWsL1SZlEooQF2f8rmOWJVOgmO5M0MaLWikZ8LG6uWLJoCIs3gzUxqjQrB8+2t
ZP3/NZqbl0Cqx3+/Nfvdow9S0fBbYyByhLyf4shyq/IkWbqImsaO3jAKMAooGoE8
BWv8llWYnOjIpavqReIWu/FHQVLNwIRCIu2YdAjTuPieB6jQJe3iwyg5yRiFXJFa
N4heaheszuZOHGd0WfKryeoDQrfmleFFQvPknAKlFp4wuJO07xK2pOOLC3psJkf+
2LGvj5bCH/lS2vveIiJh3CoNP6i//8jBl5nja8a1yOJ8j5QL840ZnrlSMGN0D40I
0gj9BiGFDpMF3dFXIhACeL5Xqnm5TQx1jg140xUS1fP+Bd7I3EkCHtJwVWaja6Jq
9oopUy3BxdQrq70Qb+1Ug/AQQjvZdAd1bxzC7v1/4JroQ6o6ogTKH8LA0MCCHh/n
xE5+ONoXkoqVZCNtt4hSoXQXllfJdA9TtQcKE7ODmCCgU5a2k0TFkr97BlvuNh7N
G7jvdwhvKGnwggL+vVxygRzZvPsUOMtNEiXYRGoHqG0mBbB7mIBgzBDn90F9st6T
yRej0VhqDOSuPOVQtO0uht0ogim5uNoxSa6zQwTuGx4x1cuWHK2RB4R2j108od79
O5nWUnDxo3iLStrTiYp66cqQ21oWQMtp9a6kacU2NegtXdaUQQJqLJdh82HI7Aqy
6Kw3JO6FiXTNpsAEoWEtEZ1PJeZBtiwrhCuIkAoNC6ZZf2IpVC3btwlKMrZ70U9p
YO+fW0AVp/9ujsMTSRDVkIkgEASE8q7rRhnZcNDs6R/0r7YR3zaMDv6TIdVJcAN4
SKIxtHp+4IieUTkYZ/hCc2U9N3hNLe34LCcIXTOZTHiNPE+x1+UorTVg756pSAzE
yEoVfoqBWPnh7+wvqlPvMQ42bURqUiGxWfAk2gI96pL+UeZ80wwPg1X12fZnM94s
Nu3CT9YN427zrn9iQedb4+fOpCOR7Dq4iaJW149h2lwIE7Vv8ntjBRoA9P8EKrEl
6xindbw63UvQfhJMt8amPA2aCzKkHuO8lONamgWv3chXGf+oyz5FofEVIWQfsPDs
3lsa7P/zCVgC7hhla6W50UJqvAoAQwViR3Emtx0bz6NT8jYQySpQetzuTuzyzNhC
iUXyXahw7SW4ZKwV9HIBPQ4GN7aVsFQYV9U2bEUmO4/kjwmKIbF+4o3A38ov9ahQ
nr7HhkwA9d/Pk7BGHono2890cbmEIbA7M5OFfiu/EGLej4gu/upWTbgJNIddXZhD
fxyniQV7DHx6ZCKlciPZirvSO1d8wuaXL1dD1fnlFuU8058i0JmNXvlBWZqqADi8
OZr7lLzNOpN0cItl9wrHNjBSCj33vOcRmkMKYDg3MbhiV144jiXmtBpqQ3fEcCr0
eOEzLaIhNCFJvy/iX1spBFWIz14N6qnzb1VG/dqxCSZLfFKJ1PETCX8JpC/oNRQo
n/Sl7d9/c6SGZZEKao9YBNL8tFyWOoRVEwfkElYLlV7aEmN+uzRBhv8wzqhkyUhh
N3kZ2Q2n24Z8eiYfnmhaeO/yFVwUtTFAWGdahbyFyuT1Pt06xqXvvT5FnXbrGPhh
rBr5kvEjV08pYn8cAqoN+xdZNwaXjOVfMYn71GwYW0JrIgDA9L3AvPRrzvWKUHpF
U/MVj20Rvl0ewJk7rpeWPyYU7Z83P4AU6d+HJpiDEDaRrOzyDoRGh40mr2nkBF4X
Bp9qGNvk2iwRmaBhLD14HMxTtqWCwaW5w/4Naa41hKeOeiSGjEivVFhMtBa+gx7F
T8F/SvWDLbx1xLIK59d25Sco0+G4aaaiSSPDB12gS4qM+7dzSPwNx8pPmhVYkUvi
/PyU62fiC4xlFPKUzX3Xln9h4WnkgIQ3JQhyJFZqJBLTn1onDYgclQTVW1VWPP0Z
XTxpJj0Qt6zJSZNXQzD6kNewQgbrFDzezTLHFKrFvuTKvpppDQUlujZV5lKqiV9E
h5IARiNrQeXy993xcXAyB7v5WViM3dVU50dBl5x+i51qDeHM7sCwKK8ux+87FGxG
SEV+nT7TZwthLyt7WyQhXGJxzC4AkvRvKkQmAwFWeSwY0atJr2UtMol4Qeep6Xla
sHSgQ3OTD4ddy4BiphWkXW7sZmMlWOESi17rodVmssxjtgpwgrKRFsHljZTG7JLG
EgMXI2qI6hJggTv0fOsw5mr653mTojvtyCDuyc81rc2GnBbXncKlUxDGzc+4YMYi
YVwaiNQO0p3qzYoAwDQ1T2DsIWPFnCuezvcU9trvJ1n551l5Zk8QgQgGJThP67f+
vP6VFhUam3CDN9H6R6IMXORvLkvH+gVLOyK90SnEzHEAagXn1K0e4S2wZ9aO29q7
kn20OKFyVB140IXDIGwBhj+CZllk244nHorG4/RrO5qC5XwRaDUXGGO5ODM6/Ena
cuw2QgVhRiznPhqJVyFL1uIuBvcdZKmI+JEq2uM4PfzIcJS7vWWHEO+lCoCvD98i
gaViQaoAiiFu2/PggR5cX5U5S+Crg8/uMMtGvzpleoOrP1d+gClKn+4UEcSeZ5n0
nsncqYF9m1L4+XzPzjYIJ5//kZDd+urGzwH1risfoYwvsJuIqfbo4mfPnv7vul2M
UMaB+pqyRA2iuoOlQhfXZc9xkJvVOQio0SK7EREOcU0sTYzuV0pIozwCYas7RcVF
llp4H09/nAGeVjp2khLKOUtvY6dV/IIRB9MUqkxSrW315Wd6KJJcJkFmg/DxImCU
pVkEs7yeSMUfnDLhCNVObnXolVJfWqrwH3T8pZd85AQ2f3yZSTTTPyZx+wdv9L8f
GV2Zj4J5sP1uqFGN2kD0Vry2TFN+Gcc202PyE0Y43PgQc9vEhmlQBKMbK84wE3r/
mVlOBwRtWwoarvQ7IenR3VmaHaBCs/CEVJmJSzlUJ87LygaQFwbDumeykmEIsJod
X/S7nhqwVTaz2e8g28+j+UvLLxMtsK1qCZ+ZriBUlTz/OcXzf+yL2H6Kt2fkbHf7
iLk8u0935jo9V4DerHHs5wB2xalLA6bDZUDbEcWOJp3D3eff8tkdsVd+uYEY8NKH
4uZJoc9/qUfe7YqElMpIdnBxR00eBTzNwJrVf3JoE9pFtLGeNdLZDHzsIKlsDbSV
mIVVd+kM5wFfn+OOOd6hEf/+I0WhJFhNmF8uwDVqx4kJh6FRXo+b50eOPr5f9Mct
JjplIbwcJmrUhTSzKvEAM8l/hNqV71sdpfaUY0bQeNxFq243fy/2qSU4ySM17HO1
vcDQutBoKxXD83fBkWBHIM/kuy7JWXunFxPojKmxvYfxvB1h6PnVokDCtUzhaIQM
Z50zt2y2plKXon2KD1t4XluIZk6kUs3p5ew67EQyfuG4mFn7DH53j0gd6HvrK6Oj
HtfcRzIII0JYQbm1FAU4KuZTuhi8pdOdKckNr+ScaSEHtA6WOXltJWDs38B/JORn
aXZYxNt6HpJVYXTVaflFrgUBMHF8rbqXShZJ8Zvf7rINzRcidlOroeI3el0jvNDj
hEf4kTAEJHj0oEtDtz+GhIQurbqTvOqT9QQoLOsmn3q1ST90O/Hz3G+POAdPl2CT
U3XtDVvh+oXkoSOCQUkomCd8Y1jl34kiJVyoWKfKYUAjpkL1ajy5zZrx1efJpPEi
C2kDAlBYQaxd75cbpNbe7mlLFNWEDVt/sbce7lAOnxFsDuEpm41OOBJ7bD+iIhQ0
np9TyJrprZL8RjL1wAHQ8WXSwcF/s0Rb3J11huP1TsmN1Fn/1tet8HV+T08h4GSY
Sp6VCqa8ElYhvnWeNRzTV6bT+gaj5yQbKHbxsQKIj+NhYQpNiCYrY/NXIJ8eoxxl
0Hyj0P96+CEzj+TooZElHxukfVSSiSi1P8tHYVJj9J6KUD6RItQgugr0JrIGbmjK
iNDyVm/0+QEb23zoH9N5ZbW3YsDmT1UhbzHZVHMmHZI+33A5fVi2URYJyNQigkYX
v0Bv4P6MM/+DyOXQI8cctkyIgR7El8cckSN/3exB4JbQ3Qk2XvaA8rk378tstDzM
qe0sw0YPcwN4eJ/P8BEWSt/6sBhILEpcoXvReRtRigfhxc1DtWc+c4Jjn/kSw8Nm
GK0EEeCLW4man1NdQfFLyJyc+C+L8vsNXtAWWdIUpKxstMKmwx+pacX3zfTENLIv
92ZdcQrTyx/IFiZ0DWS4MP4TvqqCCh/ToPuVCBKbBMH7cIFDCnx50BS0t3oqxMmw
/ynJ8upZ6FFUSFOPqmeU3f1ouC59RDXaD9g2eV0HxhOJxxQ83pf56S5yk45gTH+q
sx7DKAgZIlekn8M4qXP2p0h2fx18NOpXPnD4AP57yRduBuKeI+kAXk0Bz4O51oFe
+YzqsU98LigB49GrbBEJBwr0nOYR2hz0qI2RhsQdpAYaxOkbedxKKl8kZ5qPSNcT
fGLKwbeLgutvWxbYcPzrKhuP17JVNIL6OmiUTLG5NIBkg664McP7mP0KlhCpqnX6
J6/UyoXdPBxRJBgOSuCvbYBxoPtRB2MvO9zdRi1nNEXmQpC1jUVZCZsUPxzyD26I
K9g6V74l5T8UPGiJXf39Hpv6ZOeOBCORTjC9doMefUh335v4N8bk70SDk/gSR0rv
wr00JQFN/FKuouEruKoOvblQoD8bXY3fiPnVjpfeYB21hFt6tc8RzoBcplh7fghx
QyRTMwdtgD5hOJuUjE64VYGfWBil4Xhhe09Rp3VPmFWr5p2yF2LUXbSgNSsNcyCh
OfaZ7iZWbT/Xe24l8Zie7/q5IAegnrsu3Ft4DR85OD6QHEkaVys1FR0sIjN+6V40
gTg17zagGHXFZpdiJZ6HBd690ctI1XgH6adNbSRPJXToMylejflgXN9C5CsFMjpn
2ws64ySpZju1tnGKrDKBiN83UdzTL3YDD7Wxu0io/z75A96U369V2+i34UUrXde+
q96KgtD8CNj3siY8a57TPkUzojcr2NPT+CnGsGZfwwrM3pk4vr6fEJ1QmyXqyy8I
SD5BttFLhnoCTlpNHQ2x2pcVgWg4JfK4bKkFw+3yxZgxYZCSSNLaKlibfN/6Xh9p
JXOAylOlL+2yMbJF/QMWrJT+z3uQ6Njvqmu1a5iKf5q9McMSjshfv3X4VcYHicSM
vTNp+zIwJwoU54Cctx2O0cx7E+4dgcYEXmguP+dWYK5URanEHOBO3lBpjq0XJezr
UHL/vUBNNWwUBd6xZGoFxqPRuNjptlPVyPqRYvzcR8l0qZwnvXsFe+Iku4BCdv68
s8o/Iz9TU2taOdjg3mq50gCByr2t4P9iPyI7pH14V4MpAcYswwaXWVyNLTwa/SGY
mE6KP0uye3MzKKgk/gWYZscwl0lK9lyuxiOVMvrUhkLCoecnUcy32GOp3jBvxnrO
b4DSibKWQbij9l1xA6LMCT9ZSbgh8NRJM2oPi16kSf0xiVnNZ3Xwky07Vei3msfl
gCj2FMd/liMn+DUA6ifnSORzr2i3OmNpYzffLRGVgQ/HaOFysi5LM5SSwaKGeC3S
PKRSVCqp5DepmIdGlNmo3YE0YFYsVexUHQP9/MyRsPKJEi+AdoElfPWzHF8fqgcJ
rqcQrNAMdqfMoS5nYi9iJ49PqBmECwtWneBC77ZyjZnw+jEDL5L9HMWH0DIaGNxl
+nmCFGKScmjT1VTOC+SpJPs9pWpqwPqA6Iz2kYuIq0wxq1a+4kEfrNqO22qSgHxj
8Aaw3HJcz/+SjL6c+5PnIpIZFsPkLEMPkA9tkKWvK9AxiFdKAMZ11seFM/CZAEME
B6/kXxzjlPpjLaBeQ4ZvR2io/87meGXsJIRzBDMBBl/sAJqdh1BTAoTmtbVF7vdH
54rwLo6A3XDmvSpZd2whcpCT082LqPt7f4xAPeP6WQVirpKiRSnholpFJ6Pn/A0j
0yH2QUJRRlS6RGRtn8oOfzJ8gN2RMj/qa+ES7qyrVEJFUsgCfvm+PCXo4GFWXi6v
N1lxY6uhjl+5vwpRUR3aEHda5Fi8nU651vUh4qfLLWO34e36iwmcVOvJqjR/9Zdn
LCzwVoJJh551SQboUI0zApvgHKQK8TX7BxMZM/ueDPxvnDfKp2IoGAruGxZw65uR
`pragma protect end_protected
