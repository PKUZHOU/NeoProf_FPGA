// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ol8sADUqPGadagFfcH8CUCNyBWDkEvdr1mVqEmdXYIevnMd1VYgwICwuf8xC
dmFkfqWXRVHSV1VR0uB342G1rHbzucwsq8YURp90H27Gni7D6X0fKtRbKH5B
2YPG+EhOBtXMCsVW9ikKIVoiHd5cZQom3Nl3lz543SL+GZfsNlINTYdNxB9Y
6rN4+DlPtFNO9OIXPFrmlNffu74xOcatkqcKpzL74sJx1P4aR9Uu2cDvwsI/
S4jXStv7p/qskAkCjLoshslT7e/bwFOoEb/eZZkOyjju4XjbW0D0IQ2I3hTo
PHRbJvNRQz0vxrQtzhlFMCRbIBHHW1PsKqmKXWgP5g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WlW294ZZX8FGwkgD6FgVoUPjGYRAp9irlFaC3kyKa32L/a4rdDc3BXl8OJk4
SBnXzHxNi0Ec14G/3nGJ+jWhuqmylyzDqULejEDzPIbzuktNWaKxmfnXm74h
qlfcdnJFNHmvoYamrsIGQiWqfmrV+Uuh1KuC8H0ytuBLmsmv3g1h6Zz/C8Y3
69tOwwLAj/CSXLOVekNKONya1U1VTZCjPxyIn0XK0+Ii7Vkf/HdcRXyRWAuY
qMvELot246g6zmk5J+U0wTcJvZsKGJKkm5LmMMiB6w5VIQj3LywuW+Vhb/wp
/9eQCZdmGjhMfgQnFKY+o8sEziwNs4OXk/w/Wa5g4Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mUl4S7F2NTsobYdkL2DFugX8ie/xiX+c4nLlHKC7YP3XAaEAeTUfwjtHMNEE
7D0I/RNljl9Zx1DdU9LQ0kArgFXjqyO6vYgXFZUwvnFUIF0Lzb2AvMd7jcHo
dkByZqdZFpKhLoVPzIBZeuVugJGH+i5U/nQ/mRPglyk2I9pKJLQDer4vyMSQ
g3XqRtL8hQZqRUDK3f6R5p1WxR3Ua/TS4F3ca+5gqmlKSPCJfH5TOvCR8gXf
keT1CRuVh+P9EJZ3h0HEiu0V4SUcBVDJZQHAfBDcG9LVK/b4rlm4OI9i9tIp
CNvUURp8HFeovDKogVFyJb/gI8qh3w57Hl9m8DCSRw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SYh4B6Q2JbpM0fzQGFCVCgfQ70x7tIGKLHY08K5hNd+NKVesbxHfw/hQr5rr
8izELCDnBMxpQieHk/PQnZk9UVZWKZJemuaiJQmQF5o8mQjd4TtY7//FnZFj
X1WpnuVRUcShlkrBZBriRIMD3ldqB+6T7UBaEiuzbbgv7VTBhZI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ULB7MOwomRJhMiQb5DAia2V2S+NaPzQhVrdJiDzCJdAbxynootBEKXvKd0+f
zjwHyCpJBaTfiBNl/6vqBTGwC2WPcrFpDxGGZQD0qOxeX7tZnNSvmKqcjL3f
6KbEL3oLGcYIZF/5OOFTYRpXqWc6/ER0KepSSDbSPeBer8YY0RgmIRAlnKWp
RRoNJAFx4SSJzVv+oR5L1OozJy0wrxC1d+nQpwefQ5CZzmYaR2RmouO8CnEH
sODCj0rEcBw7jGwfYNYIOswYw5Ycfwh7WCi3303OKPMOFpjPFSiqtzAKx8BX
xDVjub3EGKEljXQ7lGndlWEkEqMC2uIcCnYqyQBgyLAqkbxCtP6l5h+Hwe1i
vJN1IAtD2OV7Gwt4EkOgyyJ1uvNZA6G4M+mYGBAp+XQw6g2LrEAHLwwfHLpG
zWNglkEKlCSBH+KPlL/Z7eo2h+wRPldSMH230ltC9JOcctQ39gKhTxbsBrj5
WB8FoEcyjIb2Ts7AD5Njb9qUmGkganO7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eeDeCnh1Mne0C95R8Lgf6GoixZO2YWFckz54TTH58FcY+bcJZ18/xonduVq/
lwsJg0VhFjNsmkVc5aPEmQyETJsDstufmsgyTTM+IKpTmFV6y0hrS0vUyOrq
rKJR3RIXTU+N6zRmS+P4aninAdEmNd2vvVLV/4o49IH4xeqN2BQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VfRBBKND70L6qgZijh5oyINiBMxYhVPAu+Iz3HcVvFTTsoruBGk733tdr/7g
kTlMUJoLPoiDgprN3+DeOZH+kFTS71QLshv4KIc0nCOefm/4YFNOBrqhtw5S
Ulr2DFa0Ia99wHXJE4+xRler+DYUufv+ksCSyH12hmMhcdGKIdU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10128)
`pragma protect data_block
T1spZnYbGwD+MkUug/G+B8uSybtnPXBKMXXYxm1/7AXzRVRALlNCOiT5AH6x
0ttWJCelBX7CdgDW1BGpo/PVzXc9tH+aCSLigHmLO8O4LzyVsAwOgLB9wFRI
SoqzRywklrZuF+kkNEfpYrB8G8xCO5FZikonjPJUsJyvH0aLkhJIOn45GRt3
tGDVj/8CJPHg/ARMcfkXcddTd9XroIC9F2+nXuoRFo5kBaYMgmAS6IdvVat2
bzZoqsx8/phJr3Q8TIwcnFL0RZkbJ95ASX9mnMo4fAtZp4gJBK+d7WZ5ga+q
fMgnUqJnSMpE6kWRU/dc9V/tZ43HLh/4lr0CdpDkDHXe64yTNv9S4kfh8kgC
r18hIM1lrJ9T92sEWyj8iYEK7kJMzPwiVkEHE5L2thTzw4eEIWSbRPtbP5FV
q4H6hnMy12DN/SCrSzm5Y8ghi717Bb3yAlaq3TOKJq93hOAPGgWs55LcqL9Z
DIOUnyMf17QeaFS0TYAp+xfT+BsnMCXzwqfAacRThuSou/pr5lnkMshVMFMt
83cggLMs3d0ryfOnAvAZVA+5WpwOhkj790hyk4UMda7WGjpa8knvqJMbTL/g
uQtAz9pxgMhG1GsoVK33LoGA/+AyGiR1Nd2eoDFdqhRMvV5Qq1qkkQHg7UT7
bHPOmPrQW3rnGP5b0/7uiVuxt+W0ijsXJLn3GE8b2ezOm5GNJKN/TfZnT1fX
KLv63ds2g0c25pLzizikVLoHtesLvZufZW8fhmpQYdLJx61LBOTkWS1Jr7UU
glonlOTshNGxUs/7h5+kcJpSGIhBN1pb5qG3soDYnIyEhVxgy5rQgB8xNZa0
+g8V7qjcRclVwYF/E2sW0GygORuPVW+OmEyY4mYQSRkeLoDblpoyexRt6nTd
0wWjFEKR3JC+MLrul5eCejv1jKtrN5VgozN+gXf980gdG+wdh8p4q4q0Rhvz
GvYuEgsk+DizpltdxAFqLnRR/GwvVML8JEqoMkA3EuMf/BDwqQLxgZE0xcl4
1PLCraAahz5LgOY9BDhJoBifMoDDGjq3HV9M3oCG1g5oMo885KyGyhkvqTWi
FesH2kwdY+rSfRGkrC1WRU0VA/AXVQJaGCx7I8WorzY8lgPJPqPdTNV0YA55
/JwmJ72wTNJl8bhHlgGhfE1q1lD51RytsbjePazRxIKQIGpdHMmoMvXkTeHN
ae80ZAFGtxHpE5pREvSC2puQpzOsJwCfZDBRkJ9XvDGwjCJKZpJII03V/ZLc
OWxTY9McUbQu0L/EeuTvpLEUuzCq9kK1pdggaz7HOTWZereIbe/OP4DTiKxL
TRNjvbslwADoITtTMtp9qWunSmrQWM1t6nTqz/ztc3oWnKseh0bOVZfy61AI
NL14h9Dsd/n5bqo+DXq90azVW5c88R5i9bpC8lZBIwrnHFZE3OGV9Xe9FKNX
vwb7lI5KTC3948rS14ldIqSpnevf1TtwL271x8U9kWfjWbGkENLvtQOW2TD0
sV6usFSk+EmPOP7IH/J9k96btPk6P9FMiEUiySs8VfM9MSIw330jSJgb9812
aKpjy2jyshYyd+Hgo6nLDYgXKiRPaYkUhycGSinki/95ia2SJyC37vPpA+hQ
LqluEdZC7wW5JKILBSF3mUr+xU4xb6TGlI0m48DJJnqkbDXDItr6KnksE1A6
p2I3vx9+l48wGYSVJsb4DaSiuSHdUn+LC/2fBINu/EA+2RVp16z7I3teVCJW
PPRm0oJ6fk6IF5gmcxPg6uj37jQ8tUDpYcBgZL2zOAX8QJfTWCNa0sxZb6p5
+pJ5DhLod+e8TmNcuvxZak3YiA4ql1v6nli1s/P38M+NE6H337SpAsq/oL5d
9yUqM5QWM3/QclbBJTtz7XlMkBkdFJGkxiQ6EDKy3ZtH7GFEnc4Z2hI18/vu
XWtaPC8GF56nSrDQ3cqzFJISIK5F2S8LQ+JzN5s8S49qkK63rplX7NISt7HF
GWWvTDafqyDF5gaj3Mj9kHcXZ0rPm0GeYnXJMhcPVK+DqZBnHQ8mID8zum9R
7qBcZtIapQJmvcHQPpaUO+AcYZ79bfWzMKp6W/hFNdH9Tfw8chMsYhOT7zU+
QcGKmHoZitpMomn6OadQK+1XkjLGkODEO75qTYMALvZ7beAkk7MoUzd5t9Rv
ifNgFretUqAaBTlEC3phAaglH2WvFNlLYrZ43SZo9zM1UyyusFdMtS/W/noF
keLm0NkD1gydJKHiPuC9fSXyJ+VNHy8PRrD/QbJ0G5s2Vq3L3mNbwKXjSckv
AUMn8c1Ww+yGp6r0s9vsx8GGYu3qUqJxpiVlqvpeIxvA0Qq9qhneZ3BAd3hP
qzs7KVOsnJVIX9Lgyr2dAk5lRa35NHxv5Oa9IMvb6pzMq5TXluJ8CSMU4UMr
V3Ysvc5f8se4wz4k/hfNvLKWKjQsScWaIV5zx7c48BdxIGcXDW7c6EftmgS9
cJ82nAcoChNaZoYs3QyJy0igqqU+5MhOeyje00IPRJA9BTA76W3WtIH3PepH
C4VYhRdUqadiZvuj6Lb8dj3wytvgRz0Vh5NltxA2Rhk6CxMEuY431kb5Cgnu
csSOeFc/ENYRXxdJbEHsfsdU4jfeYuQN9rVRja8EMyOyTsVqZ5S4ZfYk1dz3
D/4VE5I6q0F70Bq2vEKJplkBv23y4TGXSKyR55d/Dguc6BCOHo+eMGQl0DMp
pFqR9TOEPhw12vE5Ezfhia9JoEZ1jSyFvvQL/1nDdP5oVOi03Tp11VAYBH0m
jyU7oA7Xi0Hg1GJKMYSbLLNK+y32OENNirohi+WEJMZMknCrn7ecGVvtRWtB
abGfPk0HhZwQUTqqHcSiEbtiHqtWjVFfoA+S/TO/X8GJxgaL6FP8wKsVahL0
TtQl45IqRw54XiRiOA7PmEsaJRENaX/Y4DAX20imBm7ImTiSzxaBRlUWTvrr
LlGPGV0hOsD60odUbQtn6gECOlF9+fhNlVHvTRZC+wbeAa7cvwKLlbejP8Yg
wh6lXdKjQeHcplT9Gq6oN+Y6LLCi5u4meu3IuXKxSRJaQvhCve6yP0SUq3Zn
mrb85VPcMPPgUz+kZe8cCygDPZuTzUnkgroduAs0pTM6x6RZ0QXabdt+av4Q
LEdlNyfEBSllHoLogMP17Hexh1FuRgNWI78lCoF2g082szNPmigAOIF0BzqW
d+V4MbBvrPUpKYoW7gJbtcP9niRpEUSuJamLfwFpa2wEks/v30ckyS574vXr
b64CoZR5InVZSxBUiVktnJ/8aMqTXFBEshZX0IZcym7AOJm8AWqBe8u9T2oE
0aZsjNIdMLrC71M88zSbt2RWWPO7TU3ck0fdoNzWAkkbMep50xx33Qh73wJZ
K18e7EoOP3r/yQPMQbKh6qwziUgpO7N+jKTGo7i8mixigFmDSxOfnUSiLwQm
f5ziGv8za7yhoravSSoKvVSSAKVF1pN7DSg+EoRetrhb9lzTl+6YjuRvDXzl
H9JtyDaCARTEaY8FxU8dTQOZxxnlKxNkJoPxJpKTnikOdx6r5wUGtUJUww8a
ygL7F3mh3b67LseG+BiXFvqvxPi/RuMNaq2LAH7sCtsZMUAzjuynPf8nWhBR
DNK/cPGi/zoyAxu5b1dv+G8QLgERJO6VgcKf/ie5lXcnRiWQ5b/yIk5HJI1c
N+OCPILbBzpvaf7cXA7ypA/XF0WDzMxO0e4ecvdCLblwHg4HoPimcU9YZ7zx
VLuX/26Tt8RQ+Yx6jN+O3TKDHZmxxMpyCrfsFuSm6+/TPM0tGFEw6fL9eGNe
u6rOuHura3VQrODZ/7HTr3Se0rqPKzN0rkoICqugl3zDrqgZaxCwgFTJScpx
TSIyR4BrTD4D8LpPkKRy4cib1s1vf8oCvWAJAJJZmzeByqJh+6s7bLlgIrzD
hGWW1xJU5XpjlW/vfJSXs4flnQNgLHIbm34z+Lhzjwb0FN1rFUcuu++7Z8YP
6UCaDBoeUhaxmTHCDNtEjnPcA8pnunCLTRp05Zj6Y5R7qHIABkT2ekBqAKnX
0qKMLby12Zp86OZdIgs/3Undaff04LK5S1kW8NpM+RzV4j/NL1lgkQpQt+SH
Q3WnJr5j8J9VmhFYP1hF5ZIjwEiTG0ygip5La4S3ctKRVaab9TFk0ztHU4jN
5lswu3BcJXyKgpkMFFmeXTqld2SB7SMEvT/tSduJUbmBkBzgM/n4T3lkwhwD
ie76WHmsijX4KHKNjQeluHStj+35ZaYgORoGtVFSLzQ+rbS0Z4foGthkxYtZ
+CsEh+3OahDM5HziY7KD/UbiHSus6vBjuyCTYeV0d1Xx5l0JaFVtgYzdnY4R
GQzRVtw1o9bIqbNeriaUuP0QH5OndIsK0o9+OfwyzlgPZc1ihLRNW1YWGAIb
QnDBAoVIdPmZWcSoGPOuzB5texb/6IAkJBECBd0CCzGGAAPmQ4BElU9gYjqn
3FUZ1pb3PFLwM4zANINO2FXHXs8q8aBjQQRQEdZXU/rWntmFZnJR9iOzb1qG
UVbR2GhXF1940HhjzuT9knGoLpCnXEN6Q9OJ5PFwJKLYy6wS5Mp/BBp48bDf
Iw5cokyCKJe9wy7hfSveQc2z33ed2i0D12pSzfxrG/Z9Qj3+3IZVuINK7yln
qZCky7VDo8p3Ckrdijx9ED6Q1XFLNMQm/XF8j3dh/LiczU+iZcZynM5/Y2Ne
u/ODqhSiMrO2u5/XgJF6H4s2VdBZkIfnf/Fb0z0onbeg1HzNN/5jD5L19nEh
ZtJ6HJagaldse5NuacfqWFksPaDr7SNLiwYEku7UQgS80bnAjlm2EMBwX2Yn
2gyjSOwF+LM0QqLDi4EGIEAbajaEYeughYV/fTKqQHHNT5PpDK+IocqX5gSg
I4zd3W9+ww9Ke4XOCZsgWSFsHGiW2xe14YiADyPHmU9VjeS126uqgibcftbV
HP5fwwyx5nz0j6hVzRPc96huYgHOu53wPEkcp7kg6IWNIhBVAcuWFMx1D6am
Rqa24Nl9cTKo62NkGOdDGrId0HAtopP2D4DhQT1fVmjXzVPX7MdqufhSXsux
cH9PAfQk9ilFDPz7xRFZlYTjpAM52VnAn4rWOI2YTqWBxgdfaf/L9ziCuST3
htJ/V5TPU/Oc3mV8yPUPVhvmheoCtmRr2+Pk+sLOWqlmJ9W5enWn/5QZ7rJO
e6i9PtOIKbT+PbIqkwDCeUf5NkTSQivhwIX1bGdk1I/L480wAEeOCByTBeaS
6P83wL4t4jEsRlOmqVXOjL1SS3wfTDzd6XhzhmXlnMBZP9e3xH2BKUYhmdHN
4ZRU4wcg4QB6G6gtwT2gs1Uth6TutWpk3H2r0KlASCSlLp2tQD6VAtnevLsW
tHFuF7cdUEQo3c5W9RHPfU77cexWQeK2GYwOHEl1uFyCJ1aDLjWbIs2tF+1s
mdYMiF/j/mc07kWcbSc3UmGMaAQofBVqPVVq1WJot0HGsjs76RBdYiEj4Mqx
WxSunty4WsXqBwvb/rxagYmGcJ66hpM7jRLGLayK661e9il5lCJFKOOqXPWM
12v4WkmzOSTUcVT+QxctLTGCOP7FAJ4QnO2v82sYfYcRE+gdfbZj3k71/H36
/C9osvX7JDt9dGxiRbkvkmkzgasNxpoyXCy75GOxSsjyHUQWda8qvhSiD5mN
OJ9sFXegAJE+VqrA7pYBAzAOxlXAK38VQNTFDKMlCWIwbu7m4l5TQYfGQyG4
CRqZLv7seqWJafrtNNnvjmXL8pkHt5bsk/gZ8w59nKx6MNDyZkdRumbLHp5t
mEpFubZoD7LYqbRtPDK4bKLfh5I6sKmODQYH7/jP7PIqj0Q0U/9jOCxUDdxO
drdp1kv70TPug8lsgl78TzMLUxzU5ny/MMIulQPOL5BkB3M+THXuP3rTXGoz
icBliumXSiARRYzSMHpMhEhuielbBF87TC4pcXwGyM2WhQE/2KavmW36LPBr
EuIkXQ+gokXsrq/7YPbMI6lIHZKH5CwHb0I1yWW7DNmPGi0v5mTd2X2cDJ5l
yTBdpksfffnOt+1VCcDgNkG0xj0rgey2rp0qo6j/fMhbJhHMa8LKMJLkZSSM
knxY9FoecP+YsKr/RoEQ5+rtNvFV/FAGxQAqUX2CBwTRbR1xVLsoMRkQLMWt
r8AmBt+LzPa8MzYdafrNn9rGco7W98iuvdWu+/+rR2MPoZY2paXS5GXKHfyL
PEMCgJwRBiei8t5OPBh8P59S54lA8spe/hSCncEKnW7oR94Dnrcftb0F/k9o
FG3gYIDAObOkO/w4dDWUtiqJeGM2Q7CJ+PVDCo3rQHBg/H2fP0IbZA37I16E
w26QeCoS7oSTDISbdOZCXUv/G9y2YLfN9XP6GAcsgElAeZkAoac9Bz8IElod
4OQn6iQKlhuBIqNVOWOKuV7qdlMcnX8Y1cNabPsUANLLxRzmNk5OfpZLRGk5
7SRkFzdfWosFPrqgqhT5vQcvLnveNV4rPcQGJOQOHwIAEYSms+ZziNiBPFfb
RcpvJr3UPHu5S82vSv5UkSdVwrt76vBrbIdom1yKaszMnW8Qv/3OQcoIQYbZ
pRH/Ml5899sQubxu1BWDGCcT7ASIweUa9XCLBkglesguHnwMx58FvdRyg3Kx
7biw598cMX3lRM5UEwOPrZ3cI/KbAHkbIpR5QszsJQ/q3sRSGvJgRtSWeE4v
YmIUwc2cMGBVVLukrVFanXsumVaOpQzd+nI69gCBZ44pdS46RE86Si+UOE7r
p94Vvz/mUvlMM6Y3DG5ey2QtQiQ/hvnxXyNZ34Nwl2ZGDsbjv5KtQFSFDl4i
n7N+pmLw9H6HqjCw0df7Em9J3BCZFw1PjeDbM0FQQ56qkX4ANrrV8LcC2Avq
yWBByqa7XK1kezm0zO+3pWw4lkpMJBwvF4qBM6HgiZi3124CEpctySbBUuYw
4Q0HwpFTOykBa0vpK6Kn8wJg/DBBIhpyEPkwAuou6E+HqNhNrdK2ce7I+YgD
+nUtwJ+HgOIUj1fUDFRauemW3bttw+fEGzroMcg55GQXUsdZ6WAc4aSbPrKu
LFrvy4i4npipwA2ZGR4EkxZCf4mHvzEltVa+QA1CnNLeHNhxvAEboDfXABFr
7/A2lye4PwU+kuiuknq68eV18SHrxCH3ausBsue4NfQl3rAh4DYFKFLk7dQZ
oMM1KsYCzHun6wPDqeGCfWNGsZY780cV39euh4uLQWPU8QhRdDwcV78ACWgD
h0jsl8jre1J0I1aE4LeW3z2go+L+LjhZirPlEKrRNF9U1y/FI3V8C7bJ4B9r
FOEZh87HErznuXC6sbFH3vn0ccxliNAHISEHoGk0n+VaayBJWRi8LCtaiaHF
lHiQ/piN9Vp4YPTKIJKiGzp4CmOzKo/BqxLPVIzcTs0wN/DfzXIHP6p3zLMh
6zoxB1d1drOvCvpjaA1S2xnadM8+Y/GuEkyvuP8JTNMTPRruttY1faD1TCN+
96bPPM/KIm5vHeNKiK1Prd0tx+eCFd+XoEUBCrgBwaMif+Lg7UD3sh/bnY9t
vtmT6OUFUGIjbq9wjaseNjXKbHy3xlLIUvMlqWgL/9mJB3W4kPTNVTtRCvRN
JsAPFu2NgCJnGZq+/hEjS4Lj4jwcuNEbC1LczfUb0wV//VCEWumopi7/td35
tOPS1hSk1nsqyxuMOAsqlloALRn2scb5sPRc3D7Wiwyc4hJ6LxfEoV/ZCh9a
DkVRK9yQ22kVrlp4voIK1GdL1bt7sD5MTx1omVNHD7kXDs1XJh1ZjUf0vH7L
dzkDqJvg8ghzX/LDgmP/kb0YA6YdXPjH8Ubs7wORBSoef/Iv2uHJqvg6JfEm
tNhW2uhQeBjIRmVZ7q3oCLCFaH2RRTg3T/iDm16WLm01mPNbaTc+TjJC21jI
rXl8jHJZfu3bUEKjgqSG4CUKEjG82nOCVMVfOUOUeCaMjosaoFvIaUZEJVOr
skDUDNDxMhLq/sN4utLbtWSWVEFVaW2g/qHJYmo9kzQkRRIYkvAUEvdAqo1n
IQvlip8lqmJmZ43/oxlR38S7VB5b+NmlonDYiGvs8EcAcvdvBuHxaPuYhQY2
W8WHa59Neps5u/TujDdcFk/8MXJ3XkFvLmIZu7ck4AoeHfYUXtmdqjFCazpy
0XJS96OunK/qVHlLZxl25GfQlKJS7HaEuOFqM+hzOHgddXQzWA9ddz7esXvr
x7S/ygkAggAVvvelS8GWViFjwd/mxFTPoq38yAddSS9pqqm0FqIL7IRJzcup
GgYHKYDnON9QLkWduTIuJ4ninBOfWIgoHkFLaX1C2pWzyu1KROoe0msU2ywS
/lU0gv9woY0M+DJ04dtTPN4AevFLMT3gOJgivLyPf2qjGiJnBBgnX+FmjJ9L
I1t7b29R2RX7wt4L0FSoqzVJCUU1LMhdhq8VM2mfn6Vl8FBcll8icxX7HSEZ
r/LKpkjktohmH13Njsae7fnTnISLaPNAfhR5HMaSXQVO9xFCjIoeB3auzw9E
kV37mFu0+mY7NflcVQ68FPa1xvRngL1+vrfuJzX446/pgSM1PQNPuhfqfn6r
Y2DSnh64iYShsPjH2+zTvfynidhGHdduvohXwp3uDj4PAXTGjN11CnTpSNeT
X7qd2z72PeEuCOXmpFXLMetYWqLho9YL4Vd2ervjR9sA8VIzB8UxVK0/tpZZ
6Cni+voj1xKswtVKVyVP5FF0sYVqSjEFgKtKmVWmFkRP+bygDWv7E/OzykOo
GXx+1kFsjyT2+7Nc8miIGYsVuU9LT34wozywdgWpOTiG0i4Msa+E+wduQ0P5
NeiA+boXzFP3VBX9278V5kV5WeLi54NFCH10Lr3yWaHkaxcXdNX6luwzfZKs
rTTlNfgv8SI1T0ws9JGJk3iJh3cmRTsB41l8eGCRO5oi+Wkuj5+F1ckSIznW
IJSMHhB5P6bEN6AG0QORSKgP+jWEidif2zIK/C0/14K9L3NOXFgUcX+osSqt
eDpXHnEhY62+Z0Xgbipe8RtEjX5bdVcL7tWtEJO2qag0akrF+NEnxUV5lPH5
6DWa4pca7i1LXa+SVdD2HZQtyiIo2YIrNMhmjcsivQ9AP9yvjRSk271v/vhD
d5bvsvXKAYFddUc32VW1ISalU7u2KNIGIBwbYQIy5KYY8/QyFMXAoGZRGuXs
QSTHC08LvzYkzQ/6wFHRtiEDhb1/BAvtX+0pMenJNFwknp5oHcI82zO5ZIGe
OuhDwC/xu+i35syLVMyV2vhbrJ186j4m/YBOgBtx3aJhSJE05Z6JUl02QLU9
qdzCGMBwNN66O7SJnDJzBT7eEU/2KNpDW9WWBhtRXMg6jaaDhfZNGgUgDFcD
uCthnlsx3bNZjpWb8CLyLKY5m2XM1mka5wyvq5bIh4hBxzfG+A0wCt2IdBHO
PPguMKeViGcwbGuu0s8UwDSWF6rg+9hBWA5aAMKm9FgrsRtmlZNKaOTKXXlQ
e5ILl5bRWWRMvMRm0vBCf2E1RI6bHWPjzJVfWiGJIa9aiM2YXE8SufAyu5RW
FI+a+gfVsd4AhEYYAwXDte/8xTexmhss64FtWYi+wTXezUdUrOX6oqQjpowy
/LX0vbtZubsDNrmtXCwUZsUo3EEimQARzxDKH8x7gRLtVjf6XsDRSemPsebM
Gue/TqqcmcY+BNC6P3bZTf3v0OgY8crAwUJTBLO62EJMNj+4J3Tupq/kg1qx
LrTp11HxOXAmhZdcjUTJ7JonhhornEfDANu4RzmZQ6srcTEF4zhiVB5uhAT+
5uiykdC8bsaKV3aGQ6bvTPX11ZpNScEnqPH+Z/DIo1x2s/qHQSkwEyyLHt53
Y4wSMLGGGevoG0S5UWxpC4mi0nP7JFn2Ks9Cb/qcy2JOjRmeyGeyj2oePG5K
2RjuUgmYnSUHVUVVDStuKzHEgoRJRDnmOJZzGL15z9qZzouI1kSR7g802b8e
mYDzBTGMnLO5eXJaojUke9iiVy42VlruOECyIxHPRkCZGkovj+VIXXgNjWsu
g1XObrVSc/G9a6Z+1013KELKo+VAf+riUo2BOsO0L1gL7TCBZKatJ+ho462S
9/nMDbUSrVAiYfTv0zT0qThvdAuSxYZ2VPEDe2iud7wtZVini++zoO7scfKE
FT21qkRl94UffqrVDFcdq23d+Gm6icpMN4+tBj8V0u2IyBZN7VaynVFBeSgo
u+4qm2HA81uZLXOHxFty0rUIS1VqrLPErmPrGt5otq7Ni4BHFKrDm1tGhTXv
YVJHaUuvZzDe3ArMxOA72ne36htb+G0+0pKkAtn9Mf/pkHn6z8xvSAkbyT69
9IJAWqAoiHNtf5mO4cbOUU+sXd4R/B7hxWGmNruKL2RuglQxDiCs8WjUxJwa
bJEPNpsgIKeKBbLHZQh1az2GCUKPNsX3LXgtZ7nBKPQaNgez41mYe+BUJgnJ
ELSsyuK5NqRuv09/ujdElweBmKf3tFIcH5QwdDmDt9Hfmxw8VgBgEEVvhiuS
XUPi+R1VKYyjhE3LwljnBsCqGovcQ5VwGveJAfTCIfqOAKxpEmH1ciJ8n2O8
YT+bEOQ9lJSRH/gGqC12dvA7R1q0iE1leij3erOjxeLS5B+1pQHjwaUmsj0F
ii1K4AFfz0wNQTaOY5pfo6tp4ED1OpSUT9PH/DhIpn2jsXDe8u/2OF678OHa
hEd9pz9VQxNhAXjWVyt3YHeFr8F8cyUMvMrspC8iDm6XFsxWTb13YgvriU5e
TEQksNP7xBeFelSfDgZKDvM0a8u5hfnQvoM92cNFgYaJB3FK0UkeVsG2yyw/
xzeP8xfehgIDyVXprV/fetFkMjkhQjieuIzAPJk32ufxDrD2eFV2Lo0QudHL
yJrRcLZwY/F8GC4Um5uz9jI0Pt2gB+YGhxIMnPCweTZk7i0MAsp3hxt8/ITO
eoZ2nLdQiy6wm2M8F9S6RLs8+U3OGnKxcTagn0S51oQ3jEWQ/00+lsTYo0AZ
4lUEkxCmaa7+oeNzJAykz9j5M6f0jP/nCJ4GPz7dVfz3ptiWjUizsvn0t343
OzA1NtvvnIpbufdDUGV3NaEKGPp6v+D+6x4Q8cPlb7t8565akDZLIcFxiyw2
n2rzbGyJEy+6CDAzjXWSVf1DeDG90FwAYNHpwJgQmr2lljUhNtKu9nPJfqvt
TnDVxTIJwWbW+XmXApQyVWunh03UqU+ALbGWXTEIzn9qH9lGbZHQYVaLRMtq
dyD+yGnFNP7eqOtChjQd3kJ1A3MKObKWbJAe16ZQ/ZLcU7GLYftuHACw9mOk
3iliV5wY8ZYDqaqoAkUHa1m2Q/DU81FiBOVY0Zqsf2Fj90P7+Zg+aIJE3Qjf
abohf8BMyaerxEyAX+dYZTg9m93r4P7I82qZHRRB1EEAcixBNoUfBFmHtr9r
1JDk7lEhQ4A3ZASGjbz9PO1cwlsQ1BMN6MOIlP0TOt8zhU6dc7PrR7/Wdavz
B0C/cqZ5RcgWMaeSKVQP+lqLoM3ZAqZQujSb4A3mHDiQo5erL8xHx3b7EQj8
L5HGsLWUTb1w4sV6qWVsqJaKgC87umFIR669cQQgYDaXPrBJIswFQFML+JX2
mXVvtSx4rNfUl0O0QSy5MNAleHKHOPzO3wEHc8ynysvAwZgEA4WnyRlLzKTc
BB90jEvN5IrsP6BhJYJlDi3Xq/ry3F3B6gVah65nhH80luq2k8he114iOhdG
vHIPiud51R8kCy3AMMZbolNgQ9cTdXW6yU6wnKhCyrhQJfPhd+wsB3yvtXCm
tLomLJwqPyr7c/L5efItmO3H3bOhIJmSDFmLx43jOmBWh6PwHXaP9+Yd/eXs
q7RAZ1Sw+YMZjmTe8m+3hyU5K/DbNN32T4+pDwWOBX+8FoqPiI6SwVyHqfbw
sqJubmYRaCz7kI33ADRPwhWqgtJIMctcmCfohoSTH497DBzmbKsWDI5V2bA1
h+B+6lqzZRsIlW5LTibiIbZ7gSwRGjJqnUAgoDEdGXj6tQyqUWXbR0msCeew
kNXRVsg3WVXphFV16F4pyPGE+tYcJlzHSsmIsa2cvpNUHlhil/LQr1WU8O81
6juNXmNbgTSBBu5//9nQmF+Zfu+1GjpzOTIIF3d4lM9Z+Y6GFiPQj6wARrkX
9kNC9sAzlkx+BcXGZImNk6/VBuhXamiaeWF0JG7Kc82lGC3PaAvvx2x7z/At
+aL9srHHiA0pvV9E9qB9S2yhxv1C+bXlo48HXfsnUaN/gGq1pnfLz0bIA7Sk
8qTwjvBguLJw3frJrv1jPHKLITH+W7VZuVmKOLX7z3oFnrw80DVdCkE1dZ9U
VWepbD/RHjtGolQcvfRckytQ1Y0CNw028sfIJAn8b/CBvQnX5mA8ietCG3c2
+F0OGSsIquYM/QEQ8Wdpaci2VsPTFcPLIvWqYol1Ole1HJAkvvo90mWrkaPr
wGLh0C7EJrI5hUrivqSp/7lALwEHWOv9AMNeFPFtmarPcZjd8M26+Htk+emW
C6G+huKutKep8zBbzMWLcaLJFLBXmn8WllLfw+9pzL9DTy9azdzTOWrfWNH0
Izm+4BQw/RanY2aFKYmgvUcpzTV2ISYQoWGj1Uvrzz10UGdgx3b6QwZovfEM
HpW3pPCpx8ksK64iIjEaPtBBczO38zcABYRfeFSLGt5I5aYmf++yq6jRFzdC
3Cp7rKW4aOoVhTAF3ofFbCGDtRGkrdllRP6PJnw+0DvdpJU6cG79VM80ssIp
3KHkhJVqrgoWQpxpwXZIFpDmmHSDcouz8X5Mioj+I3GVOP7UTP+fI4/vkG/+
r/AzlGTadArDbZA8vB0bmpOtK2qhncvJU0LIXPO/bPdorwTbUt1LPWHmY2yk
KKRkuVUaZ7ZDoPMljhA+UxvCQVzA9wFpylCix1JZtrV+DIYpPWOX6Uh5Tv8R
zLK11HLRCe5t0y3l+n+oyo4kTp2iQuF4jOyCJM+jCep9th14qfvLib10o8l9
/ZBIM8X9x38IfVdhXXtp009k3J2wYSay30btKlLrvZ8ePstZuWtDrDnBjUPT
d6RJswfR4tyajD5OM2yNvXOGsvRHkwEm0qTakW8iirKfjkrbckWUttGsTAZ4
+UGdXMQyETL8RzAU+s9X2TwxTFfrEI6heivDJekoUm8gk5xvXeo31i1ImPRJ
lDr5hOHqZC/Id1q1RjK1usHSCeWq8Bnq3VXOC0kKf8PqRnnzUbndRDidxKtt
K1iz88VJHWvn9YxmoiuAgY9za19uwhtymEIt440PSaw/ts5m12vnfP0c2LyF
Ze8Hu/I76ohSXD4ygsb9ov9zKH+FlOO9oBNfJtuD4oh7MBXkPHYQSWMjn2uO
0uE8j1uKsWOjh3ZUlI73Aq6qvVee1FzbCaLpWCLNa4WMP0IAqrjiglFbmBia
3LLdr3GOgUAu/a3SwpFpM3+ru+5yz1ek+4wsUGt5RlNOsJpnAmZMrT8UM6bI
LZ851Td5NqdtQWokjAZ3uOvppKfN8O+LBbrSrU7s6TykrDBqQrfQ1PhzMnlk
sbS5u9+obLy6DtIXrojJN6sI8QeS8LlN+3543YQ7wa3InqMH4fl0FOBHGcmj
Wjru

`pragma protect end_protected
