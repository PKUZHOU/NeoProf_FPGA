`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
pvyPvsDUFZbAqNqToWCICalK1RKdLn7Z86rTs0Kl4SxPxgQieGzVdenlqPPPZ+yJ
ttmklXR7qJMUbqZtGiqy2OoCvsg6pJ+6NvzgRPEQHJnXJGXPwePSqdkYw2Ma+c+n
mmCBQumvWsE+0v1CvxBLDdTpmzzg+PPaGW03rP9tGZk=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 37184), data_block
7ICfjw3zLT13P7APvXw815Bmxqgf5ckpsj6JWdEnMw+40FmB0MGTa62h4bCVXygV
fcjy4+kP1+lyHbrlD4L2yNYLq6OC8CcTMKDpGI8n7P3IKkTyFKPbqxbPug7bPmk1
de4hCCyWtEEaDYXibTslH5zMeiIgXcf/kGzTxbkzHoVF79Nm8o3TckzmSTabOIU8
QtREFsvLe3WgSPjG8Zszx9LBb/B2vov4UYX/c+eEP0PojUGq/Cu/CZTxlDccMbCD
ClQ7PSZPArEJaW8J5bKpkzl54LIV0emPyvnWCTWQ+6HBqzlXNwYnl4FsoUKK1PdP
NGtrcSjdZ0VF97iNzpxwQnEwhNyh0G3Ekt1uEZoEJeyD3gYxYoKUllAFqlfOpRdi
8E4XP3CJtqO5ksgZWMARmyNIjsxin75eWQAeH+eRdwyeWqbXiKEDm/2F1DMF3R7c
vqjBflNA+YjregFlWxBHHQ+lyJIj0btrMCaSaVlOlmF7Vi5aewlPdnhXLQyD3/NI
kIzdxgSpx1wWJ9M3hMbQ8uSWfmar2wrhLlkeD4KIg73fQ5slpLfd5BcQ0OcrVPKK
q1E+6vVccMV1YCWITJSBXsNlEkI8f12vF7eKuneN6fj5ci/i2qS9v94G9SSraMRj
xuBxWdZtQ0hG6ot1SSWTZLtZ3RoiCRx+idUAQFFyf3SThO3bxDF8Qx6nePe0O/o3
KwMXwlOgVTtN7TXUR80Iv7ihv8y6f37AlVLXqBTWAf2ZPm4EwNvGSl3bcekaPQiu
BjkzW1yN9vKrsBc7cBSRpfDbvtROd7UJe72seiiySEPFtZoNyRAxmB6N09W4/04I
w7CedOA9NIEqGVWTVq/LKtaNccFMr4fx5Co75NZMaF8rKIxaUZ5IlsfDuwswqfo9
w9wC3dxMV1MqeiXc+Pdaig7i3p8sQ4EvzsJB2DrZJ6tGVjd/FL3FuMThADi3+DIE
/yl0RJojQMSSjsaCuk8sgfdwZzKFvl1dS9QTjHXEFk39GwYtBFnByw2Fa3YHKkb6
7z80TH+cPbJ8Q4Brkpnh/83R/cJAOdztAxVYyGkdNoSKKJ67NAWtXI1zrhxAqIEJ
Up8dBJyTDCn4YGYR6D7MIXJb8eCKQt1f9lY8lCohtKjXIqf8anz22/GwKUj47Cy/
l0VWp+MdJXPFHZUs1diBRNRAewBr6j+Ws23dNJ1ela2+N+2W221iK8jUexd24Vqg
wv8KEMHQXJPRd5Mjr/YPPzTpuu4YD5/YJsJKFzlm1WnEIAZAaj4elRp2PgdwafGK
3znqc4L6p4+ISvV2AepzRPqkEO2805f7b3REh7JcXW9KsQE8nlDu2zhi0uBP48I0
RF3Yg0jno57RlzyrafDOZ8iamHj7rg7QFy4Y8JEER5Ds72Vvt8pdINunSL/ST7NS
w8F7y6ORM/2aq598S3nYSIGVsRHJNtNkbXo7fAyi0Wf8XKJgWM4czihLeHfGwp6Z
KG2YGCXjVueKGpzVzWR3p6bOiDSG2bHfka9BqdltDa78cPvpCO3GvXn0YPkXL/pi
a8MHayeCTziS1JkNzDb19L52ZUbvScTxpMEaqmssHC3Gu1Mqb9Ii/fwPhiTQJyUc
cThQJVg4tyBp9IgvupH7BoGQQ/Zp1+zS9FPrnBd8/NSZOJqV01Z4yOVuOoLGFNIr
+AdAU/TLSOaGK/TKVoXnMps4Wl4tnwldTP9IGOPCB3U9G7FXiEW5MDga7Mt3zxRf
7qZIV+RSgalKQVLYlGRAd7VIhgyY9fv3Bc0ZXvqG4Rm54eZXhs/8tSFC0x6km+fF
9UddVJZB9ZJ/Jj6GzmiYFC1zGJ/z7cGAnUUr4X9pmrNjablUcATShwmU1j2Bc6Qb
ggiUw4iCRyA6KVwfdZOSJbvzj1zg5/VV82vgBZGOoR4iYlzoUWQI1daQ+yLT+AE2
1yNtNPiYhPVeaPnuG741jNFcmccQnjWqKJx8cpMxYOnWJtdzgDXkyheM1FKbYOJE
k4P209q+9bYHX3bMnXmDiuYTGKoVdo09l1BFlI55kAgMEiwEHnwKFSUcmX384RTr
BSQkK5Gk32sqeVt8NwaMXYYrybeLdvFmKFNBuN9eIQZAXA1l9X/SzcL9ja/BKSWq
mFaTmmzNA6JjRTynNpWcaXNNVucS9E25ET6TYJ5EDOC7WdAsmqkpjevQLUDMmZrr
W1+nn5APLSrfcIchLvC3xPqzzmsud5ee91eX85ihXegBB4NooP8VdqZcriryaXcO
mcMtn9Rg9XUbXOI75RfBCrMhRlNlKkNiGm436TyGSfqBfIuVoGkurGj1Ae0eyIL8
Ocx6EFbN54Bw3a3mhirG5YqRd9T+bpsB1A6btxDXIWd6U6o9ktiWogJL0ZzetJq/
dIh8jOCuNJQrotp8SBO/kqIPvycrKNt2LY9K8ZdOZkNtK4yZHhAS3uazEvJV+agz
xnSBNTEIP3RjzavSjXa9k9rxEUEw8zHyI/yxhrAugAYFu2opBb8BXDaWijWPnQ2m
x0sNiW+PE5blCjAZtLWtzQ2iknJ32L7Js/hJPwep5Lj8Eqp9ynhfCJFc62x+9ow0
hBWQOXEx88/0o+sg009AM97uB2OBlnYYOqKT/Hifi59enqDBtCswkJvzV1tlchkH
ksPE94AaloOxhGkSU+hjUTeyFdvqzQf/o394OMg0ZcXCIXL2FpuJ3SJgJHU8oEvm
p5UGwxHWuk1rlz8iecQj9wEx0ltNML6W8abq4cFFlprGjnn0OP0D5UkOWJoP7JuY
ZRo0BUVHsnCKtBJeLflg+xWHH3jxdA0jQ3r9Yx2qidiasBpC/tjJztCjJg+Q8rIj
bvJe87lu6lm8NHUFtbgr7ilDhFV4HQuy2x0m9dOn4j9PdWoNss5rZamsZcrmIVjQ
fVKaaq4exVmWCkFgBmFWo2eMQP3Ok9lX+Ps3xmfwOS6OI1KwiTnBgz5EIiUSb3Ue
WB2nGC2PDgoxjfNPnOHf9o1voCW5mkOcliltK6r7yWRyTC5XHifcduEbzJLw/Aj5
ixJyyX+QB0kpO7jq2EzQJHWaEIQKtU1cVIUvdmfxWh1VQVGFIsQ1CvapV//Aw6Q9
m0BBg+79vYpwlHhpM5ZH0fJuU6xIUk6XPfjLeQdrCubSViXVcl1bBMF4B7BTizjI
kw6Yrw1RhZnK2wfQlT5CDh3lxOyNKAjW4yIyl2P/EVsE2Q+nzBqe2S8zt3mg+QT9
g6xAD5Xq82IB8IZ3Rlf8dsybH4RL2JWQqf4459ZG2BDhnaoJmtD74ZunPjyyLH5Y
4Mh4Subk+0vlgXB+tnxthaZonwfdr09rw+F/XYsFGd9UVy5TS//u+06NbIXqsZGj
MnOqezPRY9iyALzvPg8CnxAMWbDf/2mWATsntXSKVZTdDTmwQ/rWo3CKPaiab/JD
blP/TlnWTWw+7nGTSc/cGxd8qPf/2lZoM8bxpF641S0thrzIhC5ePHzrA1lt9jX6
/tNW2IcueO3oBhc6uS0O1r/MNwco47OL2vPpYZmPtI0/TUZkvIsoFqTmI4A+FP77
2Cor+4YLj1xz9xQgDQVE3h7n371XDhch2JxuduMgz2oLxOL2Dp2xhdh6OTvE0ZmE
uTytD1yHrMn+EArEyn86k3E3X0PNDYdDn2vddxa3HeevRMBUaoBiYRxhi2GYw/DA
Y5mEnIN/KaQJl/vRV/kiISEsfp50rZXEPCRv6+jXjg3nqIcSU+cGRWKQjCuxbo6Q
23arRhNdbGlT8/PwtSytEwimVVJQlTRUUmwr6y4fPDAy1jgcI2Q/6uRbm6wtWkh9
r9K7kJHAcbSFIySmaRjyPQW3EoGUcbpMRHtag89MVOzhcsqiQV3hNfBNwtxNlUxQ
M1oOkn6yKK298ZKWaHDC7J7dKDrarLXYOdm63/IPUcRs8h5+ULpN2gByOYR3ypFk
2WOIZtHsQ0pfcm+NK345bE//TfSAy/k2LfKu9J4sDKH2RlQ+9iBZ0erTUX2Gzzex
dT/h4ErVkFz3v6fTktL2C7oZJI51IVM840kHfaV1e8Kp5cIlKu6H9Ip3zTtQfjon
x0juvrudcKblfh/LfErHWJWz/1aA39tbpn9QMD2nJcPGhsAmLkGjf/EIrttx/IoU
6BP0AG4Yzyb9MDio76UQ4lAnShy+fzTzlQdkC5hUkUOKMWkznZbhBkhaHjGEFjqM
AW3cvCWU5GKWrjZ0r1/E0wkCpYabahXe5bVSMAgoMzul6Pt06ErbJl8y3Bqe7SA7
Xqw/2kjwq5L0ueyWvmQCt49wYWLTMrfbskxytEJn9B+oy41BCk9Zg7/PeXV/Bu1a
EQytaWIrukdKqnJylORnrn6dlnx43ATGFMUjqSq/5jqLhFDNTPvm6HtN6txHx20q
QaVRIZgZkRpLbjvnbYmjJvX4XYja9nve+q/zdI2BGonbuyhNiihdhH1mETCNc14i
m0K0ILzgpC6uqPSfEWNwV2aucXRTTmI7qDX5+N4t5DQqofyhcIQTxGP35Ac9248Y
Flrh4L/zh2O9AVjW4Ce4VXknOWDlO4S5/Po5PgfRjpakm0pK0s+qtMY3vC4Ze4Oc
BbcbU5WPVcPcIpq03HN/qXpulcWNnfq8uY9nIxql28sXYp/Apva4q1E5mCrlTsGl
fkhaDVZcCY2Fs9fP363WTBM9AlLxOdsuMPXcBUvdQhPpEg9Av2WyjCxtBLb1xip7
tg1lQCgDzEQTIy2UDvLuda72nxGqQwLW34k7n6fDxMsQQ1VYOHd/zY28nmXc5fUn
BVkmtvrP+iyrC+0WlLG01ifHpSSwOwkYHa6k7MErHgpr0GXH6ZpvC5+BKaJnMWRg
S1s/vCe5VFQw8g4MIZ6AhIavNE1UiyQYXH7dRsRg+wBjqNwJJabAHnI7KguWEtWh
0v+bYqzvl8FUY6pVqnc0GuWWQt7sSIot87OSGsw7FMM8U9oB+u1fJrfqqtCCoeES
AY1rhIHqjOsKMJiB3XsXMkYCkWMkC5b4Pw/lOwwfQl4+evBs9gBG0S41xtpClq2Z
hMU1+8nFY0gRI/RStHicaiIHhyj/CZk+eA2hNSENX0BWOdS4OYsHP1lkf2+LXyt4
mAW3F8PojWKOjT2QWM9hH56cb+lR+N5P/v/tFX2/sidGh+ajjSJyEr7pnN27RYy8
DFcwdvaRpxiiQBp0i5ryWPJsTADQnlzt4QvFvzcbmnhvXEMPLm+Fo5DMs5VE+5jC
q0d78NTD84gKdIIYPV3I1iWQt+GOHm+sVMNaIGWqkqbo//03NszfMng38X8ZQZlj
wJ4vrG4cEOC/2yB5YqpRgkEMUhA9lPxbHBqvH7Is6JD2AAQYFM4usjnagAJUwAqp
vY6L4vF8NylaKz5TuxH887RhPJGIZ9m+mdFjfTCFoelMm6EVsHjIxnHNXu5Se0zE
uJLGmRd5Ym0uvrx+YkABIi/Rg5Cl1JMOVAoY8awtHmhWkP9+Hy8RhkJr3col1oZu
xoIMQsnBY8dcLNSUH5D4rCMrbO4lyNw/1UpnMm+d3A87N6VWqPIxczV+//WqYqHq
DH10Bh3dIM1sOcaXE1tdKEtykuheIsqmVrAfGwD/+uYN3eAJ8Slmjio1grAcFPvx
BXrHAxwuXW+A0ovmlr9VFVzpKOZWvIVCzCkkqXkhSnWAbpc16lXFWUQmF+JKyHbz
Retp7ErWg76yOpJroVvfSslKL6fHV4mqnztnGHW+2FbivRDDxGxW78WetT5rXdzo
yf51LIm6DZ+0IVmuchSvgLBqEX2U9sFtLF8sL61F8Vrs3NM2KZZf3zih+CiyezGr
sEdgeI7MUMRYNe/5WC+srIqGCY0DqRgZDgfWkLo28d9D+9Nw9Nf33ino6BiydGiH
ECOQpgZ10ch1s9V26RKynnX9Em+Ygu93Ugjrd+LZghx5Z3V/lPst8r51BNx1oQ9U
iFvwzTIufGzh3VLir+CS1dpfCLnfY5oqqQ9RccMIdOYpQiw3MS6rwc0Lqq37+2eH
tdRAVzJ/UqFCk1Dx5Lx5uqk5JzAExZNhlo1R8X7ZnwntMiUmrqWu6ekc68i9Vk3r
FIltVBLEVhfdqh1il6aXs1VAIgb848wntaxyAy4taruDYW8KAXo1uImwDPTpee5N
58fTXXs/7SPpLl+bQwLpEuYn8X+HWaZryDB0GxfqlDcdAmbNX7y03MnwXTGPMbaf
HNENJGiFlf6D7MGKz/I/BZUs+CZsxqYudZuiuY47jOla80/SovSvil+frL/1W/9t
FpfnkQK4frvbxpWy10H1CA4vH9Q3zjtCgiaiFS4+g56sKHBF+Vht8zYPgkv5vzy1
SmsaCZEkMVQTKtwORou9Bpp3RaVtlz657Yovu2QE6FlINYy313qcg79wuELA3nUo
H7KTchBnlxuZChrXXZiH68Q3DkwlqkZEC4LeDSKOn4bT6Gk8gfeTVqFCPxeLvAmp
ciductkFMK9dUmhXXMgx+hs8G/toa7xjUThGrkSkeIgaHe/0/gpiB//ZjgCX+wc+
Ctqct220vW5lVFZxFc9fl57PR9wzadWQV6WFjQQjs05KN4quXNK5zjlB7GNroU3S
VzIri8PXgQtxNw5z9QKC5C8H/rXL8BUi0w4+lrz/k2NPvQnF0TIsJlYQoAfitMzd
MJMG9LCZ66qqSW8jpf0KGCxrDXLbFBtOUS2ETjCnUhEYT6Z8/ZFkdUEUhtDI+f5b
zG1KQx8QWmJPdUmpRYqGPxytNnpn/EtFZd7PA3D1PtruGA3fvbdjo23K6ZSacT+x
cE9cmPog3nrrOuhn4KVzy1Ju/Zg4v/4+e5uV4mz6yg/1VRfW/mfCuRvZAdueuDED
xARIjGdV6k+BiTtAd9JGc6RhPSpLcd5KDHZIzVRCaDGu5xtN/BC0ZgQOvJl5NrTu
wFfhwZvWVbvG08r8zcQ5dNOZ0TZvkR+wAOlA7PykkYnsW0mHQr7RrbbthODDGexs
loc/GeNMOyLsSB6f+/zS83HJI3RMRsjnD2incgxw1Ma8wohIQDcABLW9RZb8J0jm
foZwg8/y+viSIQB6+Y1Ot5cNyj6ro0Kh4h2Zl6hxzAJ8O3hXCfXXGSR7IbyiCUIS
fOaRJ+VBvLJnKNqGQQRfFR0+Jk35SZvtSGEzmQoan5sNfLovd41uc0sI7Rq/H9I3
IIKsIXWTLS2J5P/90VlIfpCynPI5MtueY/NnM6lOaJdOvxUMsScajXMn2FuNdr0z
puJSYZrw6YnEPzkV5s5GbOvGZ9hGCHE1/2yhJJQliFLKem407VnhDfbJI4zol6EF
qPi8vKJ1T7hN33dJ5yY+NN10VQatPcBgqe+YoMSz2dpoZdTZVedYCYymT5fZO4rg
hSqZrcPolJYcb2I4k16EPff0VXiFH9ukFKE76nXwRybeztb5KeCbxpVUzv2raze0
qz+D7OeHlZ98O0DR+hVmV4+484rtgCvG0Kzxl0LzfpACUPnc65Xokbos1HaFeAy2
nd5rdoy+XeIwoJ+rbieaVseJeUuYQPTOaYVKZ7jH30KUR+IBcfTV5gTXV1UO7imp
yA3WZPrYVTVejFEm0OPpCa6s+/yCjN3CThkG1pqMPmVVnwKTQIFBya1R5us8Iym9
na54nU26C7C++VflfkAZVPdZGbJhwYEIxDouJtrj8jR40jy0GRbt0V3jCzDecINK
X0EGTOXARMDFjyx6R8m1u/q58QQxE1Z9eAVxtTF1d73kopCiCVdk/+SdJX0Vx9He
4Su0Uqgvybd/F/EOt89g1Esex8igCc5TwyCE4A+zkUruyhDucszxLA49Qx3iPrmO
EeNUMsTk7mmIppCC5tY4PiFCdShiuAdkFjUpg0Oez/t8xo+r9OXfheZuX3J7X2xU
7maXU0Lx4CXAFmnRuvI6o9xWqVxE5GGIAHZ15d+9gqctA4NWlwCuEvTlPCGxNuxb
LLLFItNY2j8EpfQUFATbZyhO7sEbUBlMdI6JumPecVJ768SJMMDYh9PtmgvxNb5+
6wyHXAlVe8KZAU7F8nuKrdCZS5iPkLA+W+jk0coYzUWB9eNe8zfkkGKgVlq+xFKl
rggSbIt/gJvzFBfdy0buSg6d7OK5unX/y+fOl6qUxH0LOGiNKW3rVFbNN98whqBx
aimcWy/+CqoOy7eWWh1rARUoY6NuREMemefvMMT+JXMdwgPiXpmn+BHAZh5i1Psr
HDX2+HdIEicE+5cLIhWqKZhik+tiI2JrcIlEfxydItvyipWRJfoppb+9dFufTWG/
uGKoxHB/hpzBf4McUmSqnwwsKCw6mhrJVrhhGipgmEcvYFdtmfnCGlhK2twOSCrD
6Amz1+vwjFoIURjjd4+v/dGTL91nR6hELzR8jxMh1yfG+P8fHo5OO5nKOd863Qe1
w9AoqBINSMWLBUEQUKOvJ87QL0z85Ini5/n1uRYcq4N/kkILUVYftl0eal0A1rJH
9q5e5S6Hk33l0wH2LTjQceXae8k30dUeE319cmSYqBfnw2VRRKGl8TGqv7OlyrxE
eL3vsxlfvyGUGrPvxtrwgGmtrDEIBV68aE6ChdltK2gyEWP9m8GVhnT7zqDUZMBJ
U2UKP1sHo3boxuLdnupX83lUbxVz4PPh9hxfdFaXdwyo/PkMCeiW9QqRMv8ozGFk
sAMD9f2zANaKIPoKGPfeUkqlQPHN7Uot9xJb0p5J02lO93ppdERwbYPYn+VKpD9I
6Ku/nDfLA2LCX+hSl6F/9AUJFal0bNO+jd7bX5GUmK34T37GbTSTicp18UKhzTu7
7Qu61qVBWQ8fwFXnM/7Ck6Rd2LMdiXDFFoLPSZG6gVnE9fZhQNeXZkNbFlmzgZH2
2q/3RlzE/SmP9DyXQSYpmm6goe5fxdcRlYSHGntMbDkMx37tl/95bbowqOOt41ki
aLImjMSieEfmYDffI1MJs9tfbeNjxTg2bEJoyhFUCyEtWjsr96NtEC1ikW53GT3F
ZR1KoV3OEy5p/lZ2K+0MaY5cxegAYrzJcJ9Muph84kXVqAY/oWWdlnmRh/xvPeLg
4P2d8hbtK1IejbIBxZLqWPFscYVrG6t959od/dd3GWAxO6AT/BrmoJXBLtr3qmqu
4HFjXcEwI3aYkytBUVzEtAqkideb2rm0EZ16cyCOEva401oA9q2G+xNaNAMxKIvc
r7MzHggg725j5tto2ZV1J2yfGfrmIjtjHBX+a2YaF0yQkKo/pGxCWEVwdKdnMw4j
ZCee0EdWAETKqtecIQT0Pac3i5VcSWG/IVVrryEUwRhcW9/hylUR5gPL8qJleb3R
vS6axhdLXwS/x9qTKetgpsArSR4iLpUWBfHjS/M7E9703V92WrKSm8nIr2gehCHu
woiEV9M5/ts+rV2DmX6jpV/VSKERbVttmi/v0GKVLRa3mGCjbRjT17gD9hFECluW
hamTK+RakToqt+s6LNffB834VePAcgjFPdM6MnZ2R0k0kkapJhc3gugScG9YfVEl
KraBKTQ+eEn/+j4ftCA+2Dxppx0iXSYYxeFAluH9yJCNO3+y4ezBH91VBgS8l9C4
vekE+NMosMk53Ao39xuZQGsyGQde+QozLz7hnucj/yuSO+R1wze+gIM24ZS1g93q
F+0u4ZP9ZdgGp+3HuMMKbuGNAHX1fYeMKVCldkEsziFdm2pn+XEW/RqW3A9VmANW
BvTtz95xjndNOebVNYGWMcGZ0RXzZM0aZzDkFIM8LBVfZyMQpYKZKB2hsjcmgrA5
encUDbQsWa86JFwIrbhMWVA9PZNQgfeaOnyktq4S+iY6QbcDvI7HPGIfRl7eN5y3
MxxDGiIs0F+/sMTILwiHymHcI75Rb1FRBqYWj3Ni/ONUCIcwN0+yKxVuFci0uzFa
oCIIn39MhIuJRsD5ZVaEU06SSCXZuxAaXqLLZhXCSiF3KthW/L3HQrWfe3ZpriCt
ltMaUsatmIw+/aHiiR0IbC9VFUSrE+IXTnUcv6q8QrDM2ykq3nbI4idIFrx+qGUe
Nn+f++S2KpS6SpSWyxcVFgrrNlG77Q9wXUZzko/AyfBZ2ADMVyOSyixTqND4t05t
1mBhOmDuC7E739opWBDzoZ0nu/zSGdHwhPjbhCdQnqlEwRAc5SHNpFn1ZTSp+b6e
Rl4TkgS9m5VjaUJgb3PCid9/K46qVOc3/sVy3OMkAtVQoBLETQ03c2fCrzNZ04IB
B7rlLSXr4g3blWejJgDjaz432zjAZH7mi6Us1its3bxH1p7v21JTLUN/mR9cn0+I
q6EJPpHEtjNWetrwhryMu2bSvmss2zmCJzhH4286+c6IQWf2TR2AQUxqO9ikDpLg
MUlzLgK2OcjSbsnTV7FinpKEcbHR0qFB9vnPnrkWq7/n76xY2veUipqSRl6wtiAZ
KYOV3gzekCWzSp62g7wbD7jF6ylX0Hs0HtptlRjn6MV1+ii1i9JGZGhzej9VJVgU
Q5SV8K8hpn9FCwds5xccFFj6NlnY6I6L3OJNlt1O2JkgWdpgKlk7c0hWPdeD39Eu
cruA10VbkzPUqjpMD7xOptwyttX+C1nOsrE50cWXo4+9C8O9KWRNFmiZezjcoZE0
n9iIq07lZJHMlKYjVd8ah8vF1VocDI7DeLwKd1Tg8nOjLFlxJD70TOyeMVNGTvH7
WZ6qV3iV/GtzKeoP6JttfyxzdxWy7ZrAZdfRDbrObnNSKNGNysRcaCeLb8toXDfg
FoHJPSKe+flIVtSonY5QsCblahaLiAa03N8AR+f8GgoHgE68b9Qpb7uoWk4QeBha
2O7bn2eDcvrc2S7OMAI6Zye105TPyYWhoUajsx33em/J5Co425eE34J86aZJXvhy
kzEmkFn1owxgEwwl9BrmEZw9Z5KoKu0DDfv9VTff2//jwVOiuSyAT8nRBTDVh08+
MYLQY39fXgCwUThVXvvrj8lGdT9bhYcaPhO7w05+vXQTjUkKat/FOUR4U36N3Pcf
5unXBNOW+kbxLvHpFvpRI6bgOVR88NJkjlbXXfwJ6BS0vdEi/yzQGmCMuXMVJw7b
ENOFb2vGcyW9f7KQGN12GtdTch5rnIGdkEx4yJzZRfe57xHBPsGBX0oj3h7g1X7v
mS3X1K4y7dZ9tZMdQZ5BIkqF+q+YEByT0x9va6duiaSSjzrNTXasHeYDt+bzDD25
dkz8fACXCabsOTwDe/BirZ33RorE6Afn+tNXAoM8Tjr5LItkUg+ol8sJxdBJxERz
SeX5bCxzEszkKa+c57Xj9VFi6Q+gao/9IkjZd/SpT57Ps3keAUbHpl89CDsujPks
uYmMpmIP0NF8v9KpOCfvDn4SObqGPLmvj4yMjUpiIRlKgbdtYS69WU3NZ4ptIm+K
IkLH03TiUzzz3b71p/k/80eip84n9l8Z1Xm/NbLEnFbrWT7Hea3BPIdYUjCU1CGZ
y1ak/H/bk2rEMyStxOpks/vc1GheV1mKVOanVg7PtYO90LJ9FWi0XyIsLiVwYaXB
vIEK8n76kuSiW4yr710wibeuKoC0m4VeKj6CN5Srwo7dSSvYPkU6lJYnaLGLlO6U
Ca+VPWRUB1FM+w6QOnCeWjyGhgRJDn+f3ppDzwK6hhj9OHYA9DUW2W65/QG2lBoa
5lnIgIC0mAZrM+tEnVZTutIOQcHlt9CoVNi4oDREy6sJqm+exXjBUBJTTrz392J4
Rfa7OYX9rILdG1RPjusH2UIY70XwUoVW2jeH0hZ0Z03x0tuBbMlqv4ugShVHiw66
XIEbqWXn9SMztOhVCEUbHuAz+xRagi2QFThkuNKtd2wEIFr5Kk/qYgbctftm972w
WawR5WDM9v54FimXY45vO8F2qCGbBVhyb3zSYC/j023cEXP9aifcVtoJ0KWuayMW
acxDeUV0TM3AelAPA5zqrF7YQ3B8geLDlkPcjFdEzavolkj9AXULYJPRle1fezxu
7Q0Wk2h4M3esku3V82ljHjIWGpSKM7RJWuXCkscoWgUYC9UvLNGz0az1MB7k9Drb
KvuJSemnJi07FZk4F+0bQMfSYT9fyBXWEz3+XL/vyFA3212612nP98Q4rZi8dnY2
H1w1JfBtcv0uXUYaRu20noomPZxGQOyzxOKrGluLmUGp64cF7LsoY3rkOMW5nwqt
3u84NQo1GPeFAjGQJ8sNRbC8gyyL4vERLRBG0K4Xud0m0Xo5UeaD/0uvMW5oyJek
3QUsi8yAZFlNf98eGQfn+qjqe6Et4wS5mL2bdg2j5lo63nhWDm6owQfnaC5vAgZo
tBDB2dcDWxxISfzRq6lpnQo7CpwD5lgi5m1MIYQnqaokjHwxcYFNRa3a5ocsGHD0
fEwEz+494XCAGamhc+sYS+n+oftvn4CURl0ks6fiDFKNjqwRYzlI6Kf5wsyluWvV
12LR8f3dof9kltfcs+DjxyTddzrVm3NTmUHtuz060Z8jWQEeUEeTvW7YbT7ShpFj
jX8RXqxKiBlK70fL4MgEWFrO9Pm4KVN4zaL5eltSKVOfQ/y6TU+YFI1dgD4ufXed
aA7qOMK3GlOcOrhuVJM8HD6E76ymHBdtbqVHlkKAYY7hhwAfvp/bBeXO5Ri/69Xq
IwRezzO1s5NHS7dgKvt1bSLAiRGXvEvyYXaYO8mO7gwXj96UnmX8vnf3bIcL7xlG
AGLm6/I31JEB0keHckm/sAXsIo/ZEbBAHQkwoiQe4Oor0ItDQKuMTl9C6hzeGUUn
xpqPGQP3yhOAohSwgN7O7Hr5i5pzOquuGDPBMMzDwerazFDQkpr+KWGRjs4saBvq
TS22i4gsrHp02kgDJ6sQ5fgP1zYybdatH8HKKn4ZRoK6IncmdDPRAlOuEDGsjVUd
rPL0CN4peUZAsEJmv5v0lFJJNSnCHm4FLbOcSBR1VsLeB/FLAEaWlEeYXOtUyU8U
0jCTUN4EaZp0tjWLQG+eGSZO6Fp8Ygk/wbdhp5fuzoNOX4dq/dEKe7PRgD0cXNWV
GkNJLpswx2NMN9KxgKIKsCO9Gy3C7+uua4VqEnmvdOBP3qUGdhgH0z6XWbI5eZTX
u3UIgbAlYl6jAxa3jLItmWxwpfQpcqAGeTNHWrdy7XJtGbBXF0VKGhmz7eBh4wK6
WiM3fShkQHfgHHotMLxg5KiPg3HeLx6DEYVH3nMqzaPILl1gO/TWp89A470lu43m
gDuAD0mXbsDXBEOrcdkkUv2AvL8jT/xyX+DGLSJdcPL1w+R8mM4G82y2w6fZJ0hb
Olf9V2EvIILpbK9gp4ROdj61ne8OKlI3SlriVbS9o/HU6FcnmpDIdgsxuL3tXq5b
cmR3HtE42L6ARXuIbkZNeU6HkPr2soUbG2jXQVyWAYyTxRPUjfAeJFPwWeJ6eE3y
5/nQ6RkAJCMc3PNBMkBdWvSrFTczx6J5uOBwBpjK1el1Yeel/UTEraC3p4uRr/qV
rYZu6XDfd4l6WpHHLo46oOvxLRKoEDsmAxT/rDemfvO4tGWjU5kHxMKUDr1F69KJ
qDddKzU0RpLWWv4rdm2rvXXFiw4xzYDxJAxVX4H/zfhncR1o4/4ZHSkWq/SrKWr/
L/8HUpw6fJi+18DF+KREWu60x6CIM+wdJastLIgGf/AgufPhSiP0dHMsUhiqdsdy
OWuzdAIMmOcijKqnPa/sSEQ/DK3Aimyejb35x2JKySY5byg6ySlriEAR865Wu8/O
2ABaCAcc9oCllm0ZWbxMdMmgHuLwLUdj76NZvaHoH37elYp7Y/H3Oer0NOpDA5mY
Rh72p9hOiCot3mbRB0TbWUzwzPC1XIin1SbVkhMOcjxFScNC9MoS0rQuwdntQLPo
WzF1ePCSrnyOhD/1lxyeKzav7KQXh04n4WPAJqAwEpvVy6y+3siLQrrd1jbngj+e
6sNJ0jCL64x1Ljs8PwYUNNI/Jky+rUg5+kAedwVlbGEbKVZ1mHrq8TJuTCqlBlzH
RsbOkV2YugpQdPgKbl/rLbhTuHWs8utkkvZ0dsuBnd29Vazwmv1HEL+vaB7QJ7YT
NJY4XHBdcfK+1hIO/bZ/jhaWB0E2jYCMaK43YP0Qfj0bjnU4Ie9jN0i24tOgp0pF
ECkrI7y+OLd5nNaoYzwK8IdDj7P8Yin3B1VgSGiDiFJGOdCyf3FLhjvas4JSC60x
YfLcEQXc2lIeQ7YyjxoZIxtElWrteTrOgMYOJugtPT+VZ2Zmc5cqYfr3ROEZz6z8
JQ7FA+1eUi+6o4hmcrttySSoY6jpww2rghCoAVr4kMJlmbxZWihKIUMb7QCxL+cH
wVnNH6/IHPr6CDnfBDk61jHwef6Parag9IoqCGzbyOtqTcnPnbRbH30KDoZy53ua
UdbLpXrtVhPIxnKsMkLKlrPC0nRvRu3L60IxrXzDMUdwW4cTo1stkP7r8yXC3v3L
EX5Jsr1nEM5ZZJ7ZKVjD8FLxBa2CyXLr903iCyvrIpvd6P99MFk3O0utop9/HZed
xam9hZO9/iu6rk3hFsT1z5ykKsCHzLtK9GVajLbIZ3S4UEK8cfuLpTrH4VgobJ6D
UDuOWgbVgxmm1WxHT99WGAe4dVWnhpZH6qjDAME4hObdzAnrlS6YaCkxLvS6C8se
zmRE4CN8Tdylntj1EIkGcGv7Xbf5SPH1koJ3C2Ipw3C7k8uzeONqTlkyr24scHh8
5xq74jduh489OjCc8yJCvLu/RWgbkfNVxjT2QGKJCy1lbTjGNKrs7etBBATrd+K6
yg3TNVE1TW5NC9chSNkPbZPEmzGj3gy7U78hGJ8E5wLfl9EBOcMOeXsZAbApR80w
+JDQ/8wukTd7QrrDlExEz0to3peWv0Kuypqtj4DY1n4HkEogWn+Zn+zM+g9lVmQX
wXCuBkZHD+578gLWqSkNZqDxdonSHDm+6R/kqHivu7TXxZKcGBf9Zvt++7JFJhBi
tDCRGPhnPCOw9AwLRVEaVuvu5/IFkQREt34bOZo41fo72JZFjrQdJ9D8HrIEn7Lk
ku75B5WzMy7tJEpO6n3eAMKqpxBenVNYJuTgFnFbEj5kOY2hAMZMCwMnhKUUEroN
FmIllN2dxqQHzPnYRMbGIXiyoDYO9tSfA/i/7ssi89PNeQRNvfKnmAqMZSspcePL
S6VXiuI+wTKa//KB/38PWY/mcM3I+R3d8ULoiUheuqL1EmxywTp/UBoaKqU++NnE
GH0Ojnre0YhkvWjS/H75IJHPrGo7GI5CoGSDiFW9jLqrGnmBi8x+eRhM1FsPJVWe
ZnhNIijyFuUXWkW3YZWe8/RHw5tzoXbMkJpUWNE2+JknJ+OhUX0ZIXEFaHxoyYHf
bN8EX0+82/y6VayIUFzrwkAk9/SqwD3ReXY1lr0GZK0G4llxFfC9geJFDqdVw0mT
+twO95619lWmoU9Fu1FirO/GECg05Rl6mrSKjXs4zApFhEN9kzspUF9T5Zx4mpSk
T/iZHMLED525EhMDyy9J9IvNry15dV7pOvFvMSbv+GyJSO2tFAHbnmzEL45Tlq1b
OSmTfvv3xG4MwUQAGz9yIYfbapVdzDTUTyc4IDv3Atxx6xt0cqumcvA7G0bQzmO1
qrFodZlXx8EcZ4MwJaQqxyOw1bz9cGh6c0sJqg5i0vaufcfX/o9MHYWBiD7880Is
lUKVVad9MrNGAr+zPiIakOXfuu0NXzxKOGzr/6vKxrd1NHhIpGj4gCRPfJa5ClUo
Sf4DHbhPR2DEl34quf1fCvSTFlKyjvieoY35F8t6oWdhxWPLzy6muJI496vBR8iy
YIwecKDTD2gbSBxbxoe427k1J3pjqtci1npdfp4o8n9qvNIdOq1LuNHYmoARaLrN
CI4APe+l81WuuS8JyeoZHBDqFFTU+JEuHVifGF1RoMQ0okGkHcpMEtvsNSXOncGE
Y2p1drme4bdP1Jp2UBB+TFg1oNM8rshDFA9xUJazfsTAE1vc9hULfshr0aprk4mE
+0Hzy+pKE6bB+3P0g/rL3xdPhR3hPt89qQMskxDMLZY8emsH8MwRbvxEVfczqwwY
WgUh4FbQ14SlioL6QuhebGmM/8tMnHO9Mq09naAeXUJPQx09QWkhVhYa7LC/fbJq
yVbxx4MC6z2PcgU3n2Y1ezTjvO9tQnwg4ObzC3hOj8fSMH8RURZLEdNdT03wMjJY
YrIy8M6Vy3nmRH/s5oMCceafzF43ae4klzyZ/MgNLoNUUdxb4Oh24Nxa5AOsoFg9
p2RJZrY8FHu87wje9xzszYHyQGYSE+2+gV4w/bQ/7CyBgdJEj3PkzydAwU0h0z4G
JxXHFvjPNbcL2JX7WTTP40dhOUbLqgv5ea+vVaAHRnBjf9IoU0IWygVWFpufAgYX
DakazP/iq/5a0ae1aMbC+yUtpC4ltC0Wkv95ya5Vq/9GwQwiEkO0tF/8MdyJyceV
DlksujsD7T1S2RDRdQxHbGvN4Lq+Hg48TIkYnWjDBjSQAaLU9/xsZGfjVAz2G/aE
5QeHjI2nAiWmuqFkp9idNhozDHfuSFo17TdnVP1qeafVNWvadNo5tUn+KtJiqcE6
CrV1qzBhHzbK/1nORTtsOdF7gdUq9H6Sfdl2XungFjaPJP1/In1yUGBxBeNBkdH+
Y7zwLUxEUVC//GT87dPjZLtN9iBxU9WXl7SGD+t9aERSYVdIvBWFmTf/mFWe/MUc
oaWLNZV4bRvbaXNYa0oO1yz8DRfXUeuTY2BkOJaqCbSqukSX6Oxyo83o3rwPpgrz
7xASoHK0445ucSLU9ABwAIk8TnxKattEqpMgn0ddY05+JDPAPjeVNx+iqGgtKwlj
2A/Iu1VpoH43RHcuiVYva8FbUDDYG2BCyT+eCgYzs38kI2LW+ECVBDa54+I+u/Eo
yYuRE4MzI3adBVJsZzrETqbJEHzGewTmw6b8H8nnwlNlVR7iuVdwKH7XPwvJbRmu
Vh3E0gZHqQBPfC2cvuX7m9C3xlDbEaFPk0LlrnsKmKlbNFXNnRg1AIX/eQVnnLMd
K641nltAV1PQ7G/sYIMGsLcX8a/UMvmoL4gUg2Fa6D181WwihypmrGFm8bMFRZx8
IoF2l0HBufaB8Oag6zyAxgRB2BGNHN2ozSGFV1KEc1Ha+22ggX9d9emFHnHLP/hm
gO7Gt9igPi8GA0Ww1OtLdep+IgtxqG6E9BU2cJ3begUx3y68Nue9sn6R0YAszvl0
UmuV2zFoIjrVQs5CFx28BfhFxjy+4A8G66zQxJy+nflJ72p6fKfNIbgHvrrp/ifO
39sd6QrljvZe8jmAHY+Tbyt4j2w0S2osbFF6hrxQWwOySWvCYOimXoLoC9tGEYVJ
nz3aB9Yyr73SfjmJxoPMojJpaKk7uRGCAOSDuWR63w5tG2rEe4eXWzmwrF3VswKC
q7X535YbMk4WF5yW87LPuaVobBU44SVqw4MIOf2dXjNfHOxEdZP/03FnEnj5Lfow
eH+XyEfq8N2JjhuWW20JyAy6nL1Nl7UvBH4wnpcNagRkt21YQK4vrIpqzedD0UnP
IyxU8tD+THRnnrqRCJxpAF/L/16ELO2hRjoC3UUpT1s1jXov2W+ssOUF69qP72V7
r/nRLqDbrKqjBEsUvo9sLITaA2HS0t9aI4dNYYpSyowhRfyuyk8GcbEZ9Ar1v8N3
NBqk2SOkr1bBKRgxeO3Tma1+I37qE7yOsVMLeR+Lm7I2miWschcD3A73ewgUVdqA
3AYkyRRKC8WNbDP8nBTshdYGliFPsIoVhszW8yov+339SYfnTI0YqHeh/OiV0Gws
3M6oFav96zn0bPg5aemv77GXZnHKjm4WPbHy2pMbL1q2+TRz1olXDkMCXlsYrRKI
XI2/U0k79fGmd7atYARmT2p70B9mPzY+NAubXNkY8oaeIoUjGc+L79lldicmVPJ6
qyQBmX5Lb1hIcxmcWWU98dO7MU3/i1gZbj86epJ5/1ygB0zfNRyy4+X0fxXLYGIY
GGuomx8MupS68zupFVtnyxLwtM3nrSulMkLJ3RZyqT1QpG9SGXDSrBWBePA+Rc3d
rK1l+BrcsJ2+fI8ycoBRDmIFBjvy7Gs93wzlWOX3svp0mYSp4lUOBZUwjrc4BaFW
42AWkhIN4bVJSlZwdg1kEjSeA3eA4U0JArahvaB99oEUvFfzUwFY746ZinTKgpw1
9NohEHGOe+lZCz5ClvQnmm3xs4sMf5AgB/PVboBiPCLHk+jDOXo2WAjb26Gc1lrx
zeEwSqshwtTB17ne/GhenIjFPOtlqR0IJ0BS2+prKQVAQ7yzo8CoVBFVJpxdDKgN
iYfeifuUfmb3doXFc0MQVARqO8wLkFAht3I77H3vPbK5i1KpjWFIWhCKz4n5dJDf
8zMG2JFs3JvDHEdLdfeHJLe154bFCpAHgCZVhMKK1oqHJlJJbuS05hYB1dpdIDI4
/Ev8VFgIBFkIIZz5Mtkc/03MTlE/SWZaob9DIykx+fIDgnBjT15+1Zuv5jRX8WR8
w+Aj4+gb+xDlyBM4JgXO4SZOUvx11FsngqNBHkAdjL+7TdMgHTXm864dj5Ov65zN
GNXCf69geG0E/ZrgaR/uk5xMCrGhbRRblioYu2GOKkbeZ5nU5gATLuCOlYVlCj6k
ddAJMU5zx8CUwra/14kS5yBgafFDC6v7s4GsFsTH370MKz6F+yaweSw77q8moEnj
Kh/g2QyN1jqFNj4xbFlfoAqhgkt3XBSU+7EoH1EJWPGJri9GHOe8/Y7L+2jzTivl
12lbMB7jCQjiY29e5HZ3ty7Fl82Vnp9DVLabScC5smIRISWYkT+MfP1hGQBRmt07
T5E/7izeJ0Wky0+8DfVZa0JCDO2MeG7AtRDyRMjp3gGxPTJGsBNSrQDyYIdhXSpU
LR3Hb1MS9AAd2YWHZ7RsmbNCIWe50p7FaM/2pwTYR18z2Xiy7fVMGgTx1QejbO1F
0M8lmZuuJ7bpOTdSE/UrE7rVhqap9zxsHnRhex21NMcuXKuklGx89glBtMbW1mUE
FF/R2MeF/BajruI0/+Xw2fGuYAXnxJHRccjqMvDNA60i5RQh3PNLsvypTWcTjjHM
4O0K67phMtw+dbXfww/hE2kz/uzHG64948i+X6W8wjmcUzKmJ9iDOWnJ7gdfvqG8
l/gkcoAGMl5260VemvB0pFx1ecredFKiGb67a2zB/zqdZVQ1j1IwRcADpkFwkMwr
mhd4svZEfO+tv2tBUcBgOgYBY31C+B2O5t3Mz2Z3JgnhbLaPPtlf9dI2FOpL570+
82m2OKRwW74PUs/fLHCw/6n/KYNe5p05mytWC2Z5SN8KcO0Eo+nHORY5xlgLhCId
BmOBxrGKJP2VroMLa11dp06VyEJGmBNIUun89DexQlUcYM/P6+GpFkWteaHZjpNc
00F8ddRNwAjRq/VOmt6MiQFgQj3hnRctFjGGt3LkpLZZbv9+ty8/WcN7Wf+exnuA
ypxa0gvT3exDVCc1FfFoBgc1fSBGB1Ge7bxy+pVjOSh4GYFZ9+eeBfWOvpcu8zdn
jTlfoBd1kB88oCNxixZmC6tyrIa5IPP9eTpXxHRZnVsT/nKwTaEoeUIi1uDOYNDS
GPKfXDWzA1/2GC3HBjHuGcfsFqd6vyrsIJBaAAo4tv7dJt6dwi7Y1DLBlnkdqwxQ
nsePcohckjjeutQm3CHy3OM9nA6Gqfhyp6+OnCE8a6icnql63AFkVo8HWhUuGlXG
fJs1DmyyueZcC6zb6EYbaOjZu4VZ5up1cuxaW4C9haEkhz2eVk4DTcOs7HHhs8oS
pKDhUD3gbbSyYpGcpFriAXWAhlsKKUwRUuUcyg7sT82nctya7Pv80SFMok4sMgOo
VC5Qyaol4WvWUDeH3Sb0k9oJ4jd4VGinaluxBNS1kjWaDMva5ib+QGLsRQaLY1Tg
YoslUUlRMy7ZT9shSQBPU4XTlm0zGjW3zGGtiwjrvM6cknPUwGSavUgh4gpfkgSX
AoI12eNq1NamKDcf1kpKDU1rZoRTg3VBYZfqgpcnPUiLtvmP4DVj8Y95BD7urQ0Y
C+uQugb9sGel3fTuHxTCCzJcdnTC2fdeWUd8oLzOLwmatfCdgPjYFpUmUGmfiRLU
SV//D8F04qFqp3DNIQqN45aZQYIrmglGcCyAaohGDbrDjfYvikNHVs5gcduta7pJ
f3rmOHzhkkql0wkNFQ0zrmSmztFagM0dXow6f6UIRf9QHGq/k/hEg9pqcjhhgfav
d6oF3qWICdsJ3b3HjHFlc1u1KaLYGRmy++H+70GBo7qJIfsi46IzAN6PKU1aTnQX
Y5w+NG2upTQl+xU6ytWibqxTOgWlFvb0SqEcqeJYBNV+Ef2zZN6z3wrjyR8BnT+i
TEgi4VTKWnIhCYfOxAWtQU8o6jHkv/76faC0AXhr574PwBPDkNIM9r/iIRjj35pk
Nv/BelDGqkMKSHpVqE8d4DUtaAH1yReFEPORchBynBrlX8AXAankms2ec9FFWLRI
S8ry2wof9gtA7nFsXDrQfkCFgy4KgwAobn/TOehM9RbqbSG3+jG0jndouDLBdpib
rJhpnH10PpAt43ZIdR0e0Qwi0oUlsWGj1W4MyT2Gy5xdvqMkFbsiVhtJpJnUvUGx
BaqmsMLLsltweewRDS9rxLeN0UOPiLH8WKMucKbCrffVqngh8TFUeoxgvdOe4j3q
LtH/jY0KZ/H+yjw0wz/bqbsNB0pa0lAdfLhsWaP9OZ2wB2opB1VmAANmMXVooGkM
EvEvVjGeWW3X+R0tyALC33gGaE5AqIk0kLHL08jPYARV9x9kxswLD5+ZwjUPFrsB
rmz0Lb720tgR/Yp25HOSpCB4fwGVb9IoJy89+1r4fNI7bB/wqTm4LHg6Spugg8ir
8qw40Yoj4LM+RDwfdebXIHFf3fQYfkOTZtw6Do438c//XUegzMM2VzNfecpDngH0
2TzDoWCJAcUAG7Kh+cJDEB0OspP0xw8Qge9wYa+aEo+SF8j/tcZZmgIeu+sOeacy
3toxO4Is8MdovavIluunMzVeJvzUrAtq9o8Wj3OgGTCibS16vIXIihorjuRkx9LJ
b+ZO2fSw/l+gAtfDIyzhbffiCQw9KZrN3UVO7dHGkZlfQJrH8+aLfICR9VTQ5wb8
gTMQALMBTpwZSr9d6f7GnenlfVh4cbp04APECWGARVgTi6s6YtyXcPXbLOg5q5bH
ZpWQyfBSHaC0Bmv67csRkLCJ8R8aXgQ5K5zK+emuhRyKQ4W75lJMswdM4UWcX1G1
xUsNxOM1sKtr3kt+HofWwqRlKGnU86/ITLoF3PELImMtVbKjXQyG8PwrszhR2KBv
89eURSfbx92ahu7/5Mit5umL4wOQ7J9T5mkFvLQsiybmpzfdxffdW/P18YnSVj9q
JoIqEZmO7lQc31s393d5HopNo1dpL5f7QwYvJk6c4wtxxY/iGBmkornLTtqX6VmG
tofFeHeU6wpqwcFDoZsjK80Qk9aXyg05LR5z0LhP1cuYbsgWUC59bqF25P9yfGOl
xgXtOD0Y6DP+ePNdqBQ8UgOHJH3E82KpYW/ZYqW0gWUcc7VbE8y3IGivm6DC8/zF
nMOWEwt2wbehNwlFkmWx5S6T/dWMlyugbUJAj2DljoWCFg/HjDM8asQTZfOnCJ8V
R4JSd0xzgCC3CgV0RZe4wL1chEqQORn7euHDV037xbYbXXpiQzlx/X4TsJpv1nWe
mBGXlUz8jhB629PH+4fehZH8OKZj1vPfm5O5Fm92IJx2gHqpNSPbf0uhzPeWJdWa
a/3L0m/uKeryxAfT7DnofyPGWqqJK+X2Ki7sUdzhEuS8CZEQAYYji1sEsYZv5s4l
z/imZlO8Ybj4z4w6/v5otuovoAeFiGn0NSXsZ22FYxyP3VLImnsV8TY5stLk8hL1
lb3G1peyTm8BtjnaG0HVh0emYZC94DDA9FBV13iqnvfsv7NRRDDbrzM3T5hDk3tx
oHaitZnkWOaqb8pO5wUF985tcR8LpPuZvdj7Ef/EUi+iBd8/eZFgF16DiZ+jsESP
QXXZOvGc5Bpe+6+Mz/bK7bIYnTM4WaDSsq7xbxuJKC1/AEc/V81SZMF8+ytFbnaK
TO0bvATP5ED6nM9IPZ98bI/VJDtTgNRqx/tQ/h8pU+cPv0ZYQNq0J/szT4rnHwbh
RzMLqyUYyKL3X6ixntqi3wTijEPnXoLZCBhMabJTP0JuXOB0pEg2gdJqWVU+bhKR
A2Ah8heRz1qYxRGLB7U2pMOKU8S3ACtPwh/a5/qFPYvI/PQ+3vcTMHz9Cmm3PbmW
pw6EkjKC2k+O1xG4t5J1HcIBRPk9IHxCLgHZHgwg6qlQ9xVlUayBS/F3ephj1RZR
4jEBdnQvqfDJ/f2odGblrm7bbZPIyDCidHfZeALyid8BWkT8rM4R4oZtDMu5diKQ
edlfgJo3sdN/A4nehBU3CY9DCSvErRlmzuq7DLeosmC2kzcqcPr8egWNDG5PME9h
AAzaFNPgJyIiEJ3Iq3s39Kv12fwE+uwJU6NnEn1yTdK9t1vQE+/ulmAtkn9KDVT1
mQuc1gW7RegqJDiw1ebcVDD9TADb/XUE5XHuhFN5eE7EnAyQIWQ/8pgEMrLdekrs
AvQ2PiskocCw+SDa9rNRzM9Gk8yx5c8YFHEUQntRUroPqZMYA1tpOjstENZZuZIK
sofzZNjtf5tGFVnKTVa0NhIv+MrRSrBpfD7lqOaWkFTgbjOHewIsGIe2oZr4pMjs
PjPWHUhcyc2L3rLM73icmfgSrhik4IxPB4f9d0we1E7kAfXwwYBj7jd0pvuh3LSV
AEW6izSlCJdQyp+cqXO8Cd9vM3lrDlBJUMfVYUqmKXBCNHZIN5sdtgpeVQjOAP3m
HCcVZcFG9X3RfIhXo90WHBZSRr0jPV6AQ5CxmeEucb7jSxWJiXfyB+fO7kasNyvK
l1NrQ13v/d0gr7Rm6t3k06G5i2DpPGi6I6pApwbnVj0wvSOhBEw2U8EvzfNkY1ns
5XR5Ds6JCMxKRX50WRmMR0eOa4FlizJBAMuEaN1aP+diRejpJnhCcZWmKCRg1Kic
Sy1D6sOKNUxHygk9VFezzpYdr7BRlHcsfeWK/yETpTd08fUKIrNoihmcnL8UB2T0
xYomEmHwEiU7CRBP/OgzI6I8sprF9jLEqOGwRYueS00mYTBawRcibtykCFOb5i3v
GfVTiJEmky/T8VIPV2y7thtcHUmysT3bjtwzOWztI9HRXA5j4zd8SpD14euZJUP4
i3cezVnpQuJsOV0RByS84TeJIoPj1o+mwoW+gZK03k2/M7+swl1F4yjz0z6mTl1u
Wy68IC0gzKFtTO+Mx6CWgP1vxuenjQCCdfKTA3a36fi+/HN4qr//LhJsC+2eEKEP
KfkZRiCafy6v947adaijYIHq4E/+E1d0vrF55OpVEHuL0UBb2waw2VstA2wEIBOb
xsnJFWixdjjtjmwdB4mycf4B4MCTCbljd54wFCUORCQ+JsZFLuE9z/nukNgrbhA+
nRoCYF1o0v7yYKnAlnhT5dksZ6RLcyFAUvgMl5vnWO13dYqEnL0BzkqgP29lpVm+
4OVGNnkizV1wAyWeFwjs0dM6GwCSgdTv+mXGb8Fp2xeLs1vpBeQfHak+kcwlGS1q
jCMB2FRGCP9v+mOX5bqJIy9fMbKqHUnXyaKofR8eRCd47JaTyKrC5o9uQH2gACsO
rbNNFMdQ/GDXkklQ02CPZCcVzgSCq0E0wIfBvJKXBit8zlTU7hpvnJ6r+rDgCd0G
LtiykQW84RVDnv7sgjpinNCoFvUbKq6kU1iT/cvxN+LSN5+A9DMXxBfmyQ3KaM85
uFkVlntB3mv8z8gkB3ZCDpOVISmqcsku1fecrt699fmX4/G7LwsR/0whx4+klRlv
m2HRkdGarN8bQ81QcEDoDk+FutoVVcDIqNcZbeGR8wKmGFQpPhUzDxXEWlgLTRfP
L/sEwN7zz6vAqpq19G9T8SvRYUaLFD6TyhQKdktNUJJlb4T512oD7GUPcP0lz7co
xBnmd/nRx2Pk71ZT2NDjkLp5lF+M8YWxSxQumyFliXLcVbdenk66RfcTQxPa35AO
yaXT9zlcdrGD89iCy/JKGTO1+Wkab/c6zU2nkbMXdYFUS1KuE+7/ATq2f4QQ6nRu
Go1MJe9Cc0kt3CUluyeZmTEX9vCdBZL1V4ZlS4PJ+jJ15RjUQ7h5M9CCjaMNpGaK
rBSqvHK5DI1ASYIdzH0vEifLyBs7qV42zhfw70SsKI7f6YY5dzZJbw9NoE+KC0fP
jHDijIR8L5yD74FWTw43RhEMLxS8OLQ/TuIBR4pCZs0n9zA38q0CkuPf+JykXP9v
eguSuEBnQRGDVpYK4sTl/bKX1EjXRTndoIUkSpFEOgWhaHswCQYiq2U0Bqyyy7Ty
y3EJLTXF1O4BMX+hWTsuj/vY+Jwah8KbXOD7a3OtJKVyB5zbcICpRcmH4/hE7W+Y
8XvfXvCyMJeOucsTsljLaCuqMZp171xZ7OyJOBR32CL2DBkDUeRVgdSun/YEX8II
TwtpB+WwW0oFsSjQey3kCud+ANT9iuGvIHDfTC3hsnH0Cf81YfQZ7kIj9FJnxH9z
eSA9dbTyJsvGZLoqEi+ZvNLlLDRT5ZD3SC/Gwtln4SIaO6gsTfBOOO0dWJxAdWiC
KqryduoFP2YX/mP7pWu+k//ogT53dt44inUUzYjLUgRZDxNfL/yk2Si4uG2tvzff
DH+u6GA/X6apo3fFNA2Jaye/FRO5hmmLXkQJxmvxFa/g3qbpHnofM0OhkFTRFv/v
CMzY37nP3bXFKfX+2sn/9kqACP0IRkYTv0Fdt2xiBfFEX9GIcvLBIyifTH6EJonW
vwqbHZl79r6uKzD5t+69MtiNvO+hrmGkbsFQQp3/JBN1dC0yrCVSqLkGUG+rfSdx
/oWb4i39qIM2kAo1kb6i834KHtG4Voo+vXWbecy4eaDWzkDTkS3C+TLrue2FRaI3
l0GCMzknVrpcCySr48Uvzp+ztPuDlIWrSqWlLFAb/IM2JTOG4HjHww7GOWSkyj2S
HhqX4gzRrC5AbCJ5JF+U0bgAW3ojiBLv6XLJNkfsLETBtlR5hMMqASQEisW4Ejlm
+sTYJdgz6vrr3rCK2VmuDrsopo7NMN/DJZ0BB5rRF5B+bbD6o1cl7qz9lvn7PK5g
y/2Nkh3gakLBu/dMAWhOJe1axOOZgWsNMnIKq2IYdfH0wTYhrJiEqy23Bo6Ou+N+
LOLpYHvwD9+WjIFS9nttuffuZhx4PB19nQ2mqGGpCkAdPg//mSMHFzdGRcwM716q
GT0XD0XqCFxK+6DQ48H38ovQwa4gbPDI/SU6BmI/hNOoQvXCHKWjb4hfCIPMaUG8
ocgWP7ukRhjK6NXT0JhhhvYipkJLYtUmN/Zz/mQgJ8n/GrgQ8p3yLkmpYVT+zxS1
MfAveILH+4lhRZ8FeSV5XVvSDU03weRTIcI7Z07bBIHbLG58604WY6XSx3FTBWNR
NW4sN+5GXP4Ajzd30I0EQzR9G8WMe2X9Fvql++1ZRYykcsfGplxAcgAuZa5ellRL
a+RAbit7efSEX/K9TOHYPrkBxP73IYf55uVlk8G2rrLTjYvbH2HKH8aURe5meCn0
khLRONBEc4tH8NcClHmxdGseK1pCZZrCKJWjyW8vqu5jiKAMzAvvL0Maj9R8i04f
DNMbuLdzWE3bOccyxLbnvAafyYVtOuFRh1e41GYA9aBdb6QazgioYtDNi57rMZfc
oXZ7YrOpGDmgDzmdVEVrLTFZcVZtOicJzR4prUrrDyObY0dwuVpIMZLnfYdgegf7
CFGR22yIv4iJKPG2ACZqWbqKE1VhIs1M7j4CfODpht3FwVYis4GBCLNAJ/Ms/QIY
K/KjxwakGRd1eo3Uw7MuYb/4iJlzV3GIjoNhacoQvjXDe1yOgpC/bvEugQBkEGrh
9tgdCRvMw5J4einBWSbh4EmiQzt96zAimc927sgKc7jmcDKkl63elkmBKvyTNP2v
++2M8o4VQYGicVMvbv0iQr+7HK2c0Oab2wLB7myGGrObLMCNmoLaEvYySoQlRxj6
aTx5I5J68jQp77rM2MkS+nWPMC23kXpR45AV+QIx+EuYfKgFpMBg90PMkEsD4dSA
WUYsgycjLxjatZ46KMQrhjET7vz1+IhoWQXEyH1cEnAQiUg+Zu2NseM/Z8WW1RZ7
89zKbTfjuQzK7uA6xb9r79AOb+wgrmJix0CUBmcab1ikiL5jm4o4wPk7BB49Gf0m
Qfcr6BEbjI+ixP0dd8Pj7hrLCKrtQWmn3uUyeSMvjJw6emxhLAuZnl77DxgXxlDq
06ema7+0NQQPXfdb+F8MX4a4hf7WuUCsMtW6qcKfxvF5CuQVmW1V0OGbaQ9qptfH
PrLKIxy+Tylu1D0R5g1yhwt6K9hcfvRjrnV6eySOy/TzpQfGV+Rv1HtVT4iJ5YHd
QduPZ6q0P346Le2Y2Vx2nhOizz3+U/3bMZ3fUOv7VDqVEPm3KwRZU0utDWM+FiL4
7L3u840IqRUf1vMkxljJ4dL1iIukkeiVmJo26m+KP6VxbevqgF7CMbtOJg9/K4oB
G4Gqv1Cde5IuXzoDMGmWdF3hqFjqzG255t5J05FEKyDq9WkikY/qPV0XSxwrdx/s
LYpePgaGoEN3EVVBbMAhHTB3SPgOJhcz0IHARkTLoHRxlxHgshPnGa9V/eqIq8WA
lVlzAXImbSVn1bcAb74uqEUUtXKpWQ5JW5DNW8icHrYyoz02aFHFu1wnDXahtu47
ThFbMSxv9Qz6DPxAdpF4+Ym+41rjXOM2k+k5Dnh0ILeD93Upvb+mvK8HFwzrniU2
oF/KGcQdyvY2FCOOKEnUapKo+0EOERYPjuGEbczmoC9xbyr2fOvsG0DkSkdCs8ID
YhKC3VEmTecTmxa4f3CUKiC5Lw2nMhbFA3e03CvZdHcT86JUZVv1qMzSY5tddr+C
vYv5+0lPSPhkCopyXcKQQ/PRuUWhJA7XImsT7ljDntOhoIyC4Wtq2YObCqN+VRcU
JHX6hSrzwuBK0KCbXMyDByquxY3ZUurhNT870EeRhqwjYISjkqdxq6TAOLehVrey
+/pHKZlQeNXzKPnO5tHWdSAp1JO4hIre5+h6QKXCnDMrG429mCebMycsXFt8D8XN
cVCmNUKIauB9NY4BlXhf5vqrM9AQKT51V1BpGOAfwyArlQgeWutLlAzObscDhKyT
PdroxqnmOlbsPTyLtQrLZDWcZOhThv98lvY1bLf7C2v1k5AoC+Xo4QitHrz48qxt
ULsA7WJPmZjSRdViVwFzMxr8jJ2TGHqJgQ2I++RDizb8u1aGmdhs6lIqFtPeoQEm
zRuFi0+nBvc366Ymc3V6Cx1Z0YPgO6VwaTti6WuGGSeYXEu0OXqCAGhzueL1KAWf
lQFRTwiciwcfuhE+a+1Yo9WSCmZfBathfIEFWgnz4RVCmcJNRjWLGSk3htIwPG/Z
1W+7KuDJYmXboShF+uJef2wNQBxQAuOUPVWFnTbCGRj+f5vQdP4QoM3hsAeNc9Wd
y6MnbBj7ODrrmupcdrdZDnW2ewSOtbJ9S9hI8t6AW2x3FYWpLBqr+yV8hIyq8mVj
iDHX4SbhY1y4ZdVdg3Ta+KKh0Ok2TjvBTIMdPusZuZRJ+ST3MM7haGB3qSs0N+OG
jSU4E6wfUp/owg300hyrkyn0m1fyd10g/MbfGJH8AJuTn/i+vhngoGrCZj3n3+yo
vPUnAUh+XFDcKcglqqSEe3JLKsQi6ogMU6ckFq9xdaezjcDJo3jFR9WtIaxdXZuL
iaV3FktOq6lvZvhmPE23JLIUlOGB5ZxlwmQx43u6+0QUHEzDry3Fl4O8iv83FyvX
kro9Mcrry24olGgxu1ZNxQvXc5N1QqAeI5D48/+SqiwbG9JMZRdjPCRnXJTjpTQh
bVm9X86COq0oRf8/egqdacXkPW85//TbfTfCRnEWdVY6waXPhTrhCpGwC8UyCdGw
UCW8b1YwlzhSKBndbnxuW+atks80jJYadILLLcMFSoYVXfOwGiNpNloG2LpGIs6I
Apvcq1jIX//upQT9ncnKjrczC/j3myrz5Al2NbbzuS2RfNrt40eLpoTECZr8ZGW1
bCE0jQ6k2tVK2IssP3VebkDb5kx8L0+xeX0zeFuNDpTTjBqtMX/WISFb/5+24GQ1
anen6VnxBp0CYzEQqe7JCzCUkRlnJpM9L6oqpC1itAHeiwpabVaMSJx86NzJL9rs
jaQTF+bqOVnat6guR03Ld3JwzSgf+fzpHQy9rjeYIEzKY+fSlbujcIn/GgWda6GB
pRk3GGd58O6Fli3ALsHa1fRUyKTSL1q6DPIOtYhlembHrLX+Ic2AKqlowiuTYL8l
5aWvYPwb4VHWtW/tLwae2tvoFou+GvEoW1SqmiMpjHsPUWdfOCajhipfQqVcAOQ2
nlJVn5hXkejdu56oGnNbuS8WkA0WBEE38eGmlwko7jkZ/v0lsFFNNS2WwzsP/jkB
kTeQdrHyalnTjXgJ521POD9ced0PwlihOJB3hpCUx2mk/lk819KNpYBwH0gw72v2
aVCEwfIvwTh2NqCtF7BHgeAIqlNTzW1cYEjvtc9Uv0Rxwzwji/ALhhwO1nvda/sg
KqaMIvbGmdWjuF5EBL7wjIAAOPbrQ9x4EIOTOtbDeaSFlY1cSJzdIg4ixND0kPKk
AZZXZV6JcJ4yvxQVfsidTQ3W5Ghe9cYvzE1fWivDGQm2ajFI3QZxSz7KItYhQGEQ
4vYxwvliUbIQE98T8DFAOKW1mcFSlRHSyMKdkk1FmbhYKoP68GE6JkZ4kATbvg6o
r+trW0opXaKiHbw0YK2N834cE7sP+Lom8Ax0sIp5qiQBJoIDE1UTkytxDxlPe6do
g01yh/BWVLl49sULtLTfselC1HULfMeLimyH4YtZmxpNI+IxtwLcMp9QLxPTtVok
/FzLBJjBWvBIJaNe0eUjhvl2skpGRllSR+wz3IC3d+CkbHtRShRkRgIbGDk6u/11
vLVKrdIlWqoA05KHzVCcmjI/A4rE7kqmyk4Wa6oXwqxwDI1Nm1505SN0m5PGWpvA
lWtZFZyyo3+pC7HRKHKDzhuuHVGtc9xc2nkRoEUuWnlZrNQGwqb+onPjfdMICMWd
RdXTOxPEuK9CRPgX2QSOrMtC8DppQGTcLUx7qh1YRWH/kfzdmV71xoMwhNqtLbQg
bzH8veL8obgYWjKFBbTcCc5oAaGH//sZEcuQlnFc0DK8ZQOlPHA08R+dVU/oMQ74
FKKC+/Vh3G19ToUNQpNiezlLb50Y1Y0gnsC2/TVV2Kqp4ir8Tabr1VR2eSLc59+K
xgt+me6E3rxLe4aN1JmNFn7mXCI42cGgObT65Jgvhv9nGFceljTTjIjMge0pF1PT
0lOOPsH9slbzRoN6/r5vze1gG5ho/xOeN6yPQIqMkEzunpttWkiPZVD1kcDXe7ln
5A587cSkyVXwiMRJM0PfoQIZaJOpW3yxsaMZEeNg7sWU/6jUt06xbHLpENzKSot9
n0Ner+DrIVM6ngE+rCVEQKwp8eI1iZ7e/Vjhz3s19IegqFupuJIbO7CIciZz8Bn5
abSw6XhRFB8FORpOv1eG2Gv0f7yJ5jojBAL1gN5ffdfo5hueGGKLZA9rkZcEnPqu
Y9jM2bji+meYeBnDlmb9Iy5fJslqLE5KK/p00Sg7Rh4BbPcWS/1NpTx10DSfiY4h
kipDSVexAG4wn4kh3wVBwL64fF+5w4l7/gS+7B/mmed3F5F/mS3Imq6mAs4cNcl5
4D52epiQfdLAN0i/20uEKkr7yfxvOCXO7Hpqpc3QW5U/kyo5MXai0cNeWkQkn2rQ
orgW4B12Dfd5yLN16BDFzBjZDVnxcC7RWsjA+9k9dg6nT66vsWTr8Q9u6KGqqRmJ
vopz3TSnLxhXy01phbroO6V2V4hLy9YmPHf/2pUKzH666FLC25jMUtIJBEa5mg2e
L4utczwFP0reCiswDn3bMa5skMKgqYmWovCqZKS1Bt9SvdHsJRjnoaFJKY+jZT3W
rkffI6cYZSxJN2ZvXDTvAEXJtrTZaWNyHLfynv01SILsePkaTgDjJ++dAVQ0ljzK
52JgwnaUzaPc9O6mE4Y0rFViqXjaPz/ryNM84dtI9D52tPhutumgfNSN59/uUchk
imN8tdfKk4Xm4R3Lm796NxChnYFoqzLloIkIjrS92U6p/iTYvrQB284EJ6U9n2hG
iCZVxJDFlj/wXhdBzXAS8oAf1ZdUVFOMG5JS7wOm074BZpbiLsX1uJHhIrgxxSL8
x6f18ebdcWCqcRV09V8nun50YmPsw6acoctJhlKIElViH+3y0ANCs+WQc9NU2XWi
Wzw2gr4laHEztRqQ5P9YYQA2ObHZeIg+/pzCEoDgdPaZa3pEJ53YAxyGCGYF7Qhi
v0qYI84OZYW61jXfJZXIejDKV1O2UGzxP9PKEjTpxFMWDLfF3d+XCaBwT/053giJ
s5Mm6qoIvHMkQO3k4xTN4kEUYTdjJqHJQq6vuV293BLQxpExyKLIVGhmcq1jLi6S
oatNe4Ml7CgmJs0xPNySyqIspfFKzlVYSY6JC8INpPaYyvXQuopDhSl6CrMzxBfs
X54HHjD1mWg499mk7N03dC0ngqYh71PX8FlmTW2OJWeXqW+vt09QcMqWBDlSaMdm
bSVqvrVogxyVBvfHAhjexHMs/WtqD3L2rKWeRAmHNreuqEq748xO5RMm0fbEBzs+
tNe6sWNOyQC9VbHfxL/bJ8QYLRMhC9TLON9hED17xz1X5qqYyyOA0UtDGsfKXPtF
/Xv1ph8HmA4uIgohSNI8eS5PulsScTBkeI/cfvYMHVZpzutaj2bNuCppFBO4actu
bbcxjqv3QoYVurTsVDHdeCKFmSnTkydeMxuzCVMidUh5/ISqTkADZ8ZVZd7EM5s8
BU8W4VtWgqPwLwP+ufDhpkYcxYZvtQPLR18MOB18ice97DEXQdqHUd+lTRg5JWsE
LWY6UFVfGfoh6B5uHhltZTb+9AUcb92PJnM1qWJFWHfmaLk6ibHAlvrC4aKcAghA
JMC851FlSYnyF33PIQwtWmnQX7I38Yq4okPrB54F9AT8yUO9deF9gyhRk8Ym5xPp
SfKejE6X2xwjLIrkPAxlWdEusM1L0zSqTEhmQW62oAOrJ8T5nzrRgWQVY3zfJSAU
31Mw1ddD8MfgUafmrbn9MpPrYxvve0TX/9C4jodM4o9+QFxMe9zjgBbMq/EYt6iR
maxYp3iRBevEgQhSPa2wTcW69fUyIrFFmr9rH1wI6Ohw5BjY0KYcrAZ2Vu0U+f7q
xArA2oUUeFZnnxU3eQYBnLFr+4vAnlPz6tM8mP1NC2u+aC91TnS3XNYzDp5yBaXV
IAK2yIIEVWfi2/nxxRkUxgU3uBo2gSxLzuTz+KdrAAU4EcEO2WJKznb1154b6HNi
tpH7jFtO+dwZpD3xqso5uyrZT18HX/c8gVHZUuvPZnWe7Yy4iREZrcrIY8w6CuYZ
0zIQ8bhnX94Yo8oTizPQg5uMsMKyItH2gM1x/K72q8t/mqtddbp5gu83YmBoS19r
raaiGffUzkoUsKPOYV3khmzFFjqlXyn2/fnxwqSD3KXawpmqhWOLT3qKIwJi1JW+
FdIb+5jwHFbAnseK21xp+7KGtVXsamXf2PL8GnFpVqW1qv+PDyC4hj0TmhQx4GRh
wNBii5DrqaIH9ii0xMsbY+FuFB8Xpu3KnLPtWt2NN71PJuLy+heyxbqq4LQBpOoD
Rl8w6j05ZPfDPixgQD1rxjPO+LmP4v7LV9DRwTt+fIpqtZk7iLpUuXbUUH34ZADF
20dfmqBQXNU4ZDV0Yh3FW+MfeDKdvbVb+TDK7Ak0z1Sa38nnNXe+5RdFihrLuRDi
OMJf1XdmoyVNQbOaXjh/GSbeQvL+oFT0H6ife/r4SAqcXhZqovwQkyxtfXag5+cM
r57c8uQs96I4JcNDY1U5MbuXNyJGdFXG9txlIEmJd5idpIW1AcrBNJiHxxPpzfPn
YjjFVIygquvTVK5wv2dWCx4Cb/Y44Ofyy8QdV0GYgBH39Uz9GX+rcimhf1hWj3FI
NtPgoCJ3LZ9LUZFX49VIL+Aoj3qyC8yr9eC6k0LHspG8heYvjZozPrr4XuSPKpkj
ehxFBozI+J8KGke+LiG3eL3pr9gBvYVgn1VzWHm5bvY8xSWnhLIEtXY9wkbXZt3X
mVPOMdxwXb8WwvcOSvux4LIuNqozbE3NdgSN1y70Dekg58bg5t8PJnzqn7W74Y3Z
aWDw64m3XyuEoaQRSprGiM/CKISjHHDYq9kfEeFqkGltyZ1wRG1WWUqQfmC0UcTd
BtUmnFfhzhY3SOxtdLpBvXrAe0h/VDCckXbFzcbRooWbEZtllroGTA2kBQE4Ro27
NUi2ydOms2wlndITiyLecgIFNdDMot4rSS73DOApi0EoO0Do06FhI4HWbSOEdyaV
QLxtgmIUvXjhVVj929JmzEsrQr63M4MITBojb2FjCT5R+2J4tbR3id0BQKC4EJgx
UMW2/46XBww365lTLK5+8WI01BrGMJVZqLvRuMmtzERD95LAzgETztNhhDqAVL9Q
Fsg1rnUaphVLEzzrs9yTkLmLF0Ny8fe/AfF4bepof3qrOYSxxv/xqOVQQqSfwSzU
EPIUloE+CTdvaGuXSSlaNnhgs0cXERp8cADTN2QlW+8Bv0i715bCG/uzRIMAZYRV
KddkuckrKzvApittLjTILPPw+ilbZJ4mXxMYANuR6OAoVRTmRqYTNFJgqRDYWGN3
8RtiFalPOSC7iqrwvmkXemAox8K/xzQJ5ndvtzDtaeS9KZaWg1spmkOA7aNPxAk4
t0V+2DF0hL4sCyxzmU7heyM2TCK//uE32JNSxeCp+lWcoB2e+oytYOiM7zZS8AfB
FjxLQ/LTx//6IzP6tx+Li5v3HhtfKQTY7D4uA6etgTa7v9bWy4zTj2f1gvttL25t
a+bcbzdBYSeO/kX/ERKW2jFRcCRKnUUK+MTEB7feufQ6eWqvTAqIu8/3Pv/VdXQg
e7XqawFE5/ylf4L2uRSaW8kYaBAtxn7qmj5oVyLAK34IfAwhIcUl6PyUh+o++vYe
xzMaeLVkDg2wMtNiDtW8jlRQl4NDxiTnnmxvh0B+h9xpPUibjkvzN/5pLYiCyZxl
H+h4x+aH3Ha617bDKmJICXl8rzU1HJgF/E2d7hzyJKZKwUmRBF62o164DdNCZVIk
hzn48BKz05Nphv3+kPYu0qMaz+5CrkMBYEqzjddJk/G+M8JDWMNjRyCBIs5TFgqf
yBpnV4E1fnGGiVlC3Fc3GeUfBM3LS/sCofGgH54TuwC5BQIwgoQmyhR3z3L2seea
Lo/2B8bpwlb9HPHHtbz5gfanJ/lhf9N+aKwnKd55p9ZsQ0kD5/UXVRMEteB0NCOu
q6CG0YZP15EJUPKg+7ytCixYN6DkI9v1uH4AGOwz8rQAujBw4a1NSJkWKw+AahPP
AuBuH1AIxTjJlPIPuKKwiRdd10bKyUibse9pzFmC9jvNvt5B1jxCxgxQQLmYOwBV
iqHECzW9psasgXahY9VS+E3w8mAqBWYLRux6wkNCvrR3SwyuBstpBNOj8zvU/wbO
hZ4BHzzF0vJZFNEasUR0C0LmsUGVij3Pt2CfZJKkjU6hsmVJJNuKFOgOLsonKkMX
VqkXbI2w7/U/DxUUrA/1Pih/Q7MRkoPzCDIDXVYXisrDVA8c2Z2JJjb52nxeParf
Y/CiiriMFAZs8xEcbRG93ywHVCaXSg9TedQroa9cUp93xu0mEteL6rOzk898acLH
s4udPrqkBSD/dt5Zt1iyJvh8BG8DZUaRWwLy1KtV1h1BRTdkeTIodOqjCRn102EB
E6kVHrXcbHjg3FS+SlM5MX9r+R+CJ4yzA2R5WrOiAmibVe4qgIHpyZOmUHrBQ1Lm
Kp/BKo2hPesxnuoUI9zNsyDUTTFJldwP1BJbWIkWmXFU1q0ZkkCqmTqbIEosW2ce
zuppV2xKZ+p+h4CQ2mKIUWAaHbf0ONxo/ju3b7R6prtAHCKM+Mt/8Z4dtkQ/ftd0
yrvyOfYd3pObUhUCE30MJUeCO2s6dgeR5GaIXGb34qzI95ATPwAv1un2hcgoJlru
8WgKk+0BBXP/+3NsfoW217JgqFGyGfCN0EXloXmgo8WzwHJuOJEp/p5TPXwZ+J7Z
guU91vt5cmwLGwIw/m3XXDXARNCDNZfnkrnUabyl+FKjUn1G/WsB/gait+38E+bf
Qf/KulnhCnz/e6TO7tTYUhY2vujzkVRvsC/iNmDH0aoCemBVl9xWnowqvG5ra/Xi
BHzX1VF0O4Aqr7/1ciwlZ5EVW8a6mA7zQ24XwrorjurQsqUUc4ymozWq1CuE+A+M
gj5l2oA2brmg1mGcqBrqaVSSK7ukvcK+wml+p26lpQMVkuPqy7lR3veHuRUq81Vr
2khQaxf/mS99v2Pn4SyiA7e0u0zeaMisZwai8FmY0gD5EhH8qp/yqmdBP6WZkzOm
NXACT5Kw/Nc3/50CnuPlt5eLRbInYe2drFXPR4UtoO1gGapqfolj5PTPse2Y3+z9
pcrNnX+J1Hj6Ulz+FKZtr31xylqH39O9HGyYqStcy4QgXP4F28et8EydgZH8Cyqs
6ttdowtixXiELwfvPK4iVd2kjBMs0aMBu2/nChIiYwNu8E4WNln0unAUfQVxGMdq
oxsIzPY1XEQfu1Qf7apuXyf+mbcf3KSloohU+rla+84IeuntN2N23YQPqexUutRC
gK+199KqSnvY4E36cWt1QjfC/yESXlVyLoA4c93PFfQK0PoqXCA+wKEoRRHLOAvs
YLFEmp74H8lE7Ed55yId3WnMEIyzrjijk5LX/xRbFW/5G0/qgLRH8D4BITMfnGvo
H0AR7HW97azc4G8q3UpbXKKagWGmodZmlThBLIpmvAc0hiNGWDp9Y2ZFRNLoToCj
AbgpLI1O1XxUqXUxstWciWz5Vci5XRyzyjsROYm8cmM6xAIaHWeMsLIUByo+7gt9
JvoVZmu5jo9gx4arhLhvLmXdFuQ3YEB8rxTOgzTlsZYIjv8sPpS99KyAAYfICFLW
bPuQ/W6SHNRmELYaKpNr6Dcw3fkHhNqJaeZ/xegibhhle9ZF0iBPWrwMriBEcodU
xDnp4C2mgyK4mxe6JSUaNpyl1sRbIg0XSPDlWA3Tfx0n1RPlocVo7iZXU6d10XfK
GdVcBajYmx4M2BHl8Lc9iqXH7RZ3yNerMWcMKyfxlvVVVydTs9LPaYX46OpUC+/Q
7uqz+GJog2s2T8Z6wuGD3glaD0UD1MCcW3bQH6pAAkn0sw483RdTb6BXs5cyD5SL
QRs+GQCOkIFSWcmaWpxz0mCTcoH11xWRbvqogyBJe4b18aDsRMNtlMYkzA7C6WZb
KuApK103Lf7ryUXlUQjDDvtXSUkhk6dVxP1RpybByW3ZiAZrmkgTYLRyY+v//gp9
TZa86Sgqyz/sNLcRrHNoW4jL4BP5OzxORPDPuanPbtZachHaOZgltoaQrlX9hrnV
lry+i7gvMjMR20TmT/VbbTRVzl2RVNQ+EM2kQbOjO11vdki7ZAIKNr8U/oOw3hJ8
6UuFQrhCryjMkObUQh9zSV26RjwKWPdcHzkyjDJuTbV2XrsHyuyUqi7xG1EdGS3t
jL5w5p/t/flZMTdIAlamT6Nsbp2g2pwBfHkHZ0mPZlowkjMKwLG/aJnoZDh79VuU
s9Dh3vUxo880pKuh4qkYG+gv+ouyh1P/c+VbmGdgSMJU3B00QZUAdH1qCEPXfrMU
VwNPsp4Twm98DRytDyYhvOzY53g83AJ3lq3meYdrka81Ir9/ShNwPioR53WFEc25
cNLWuIwyZgnGLSw7uN9kwmO6Ho40766H3kqG/zEkHVLOkO6/YM3BYo25gh8LnNqv
W2Me3xHavQQmbjBrOtnpkTf8ZV32J6RJFvpRqorBFly1qU2TvjohMvLIT9Nco4HG
ga4JVujptCHjohqR41rx45wmQq14EOVTnsnNiJWw35S6ILWhNE3GuiTRdIRbIC6S
A8dFp3MBgKkUOP1nQ6O2njaF+v0V0eaIydHYDSWBFz42A6qizTJ0qFu08bAoKrxv
oatN0DUxpRP+wFd96uERRt0rjUU4r/oX+Gz4axOtRj8VvmFSB+xGWXtVxw4Je71n
z2QWN+97VeRSBBxJky7yBsXXlroaw6KSGJCM52xeUZOMG70Sf9wzyTc2dIBoHgvD
Ob5PES0gIUVYAvQnHcSSZn+BCCaDeKFxLQo72yPZ6X3lK0rVYchZl1rRBkYumvix
4moUNMpRLHM5YGHnEHUQQT0p8XMmvPi+UrR4NCGKbJ9YaD/VszBO4aWRKtN3hFPL
w2k6zU7clScnq6PgCINjQagejI0ISgGE12jx0U/jCuqx1dq6XWoA6UHLj2ySj7do
mh8DFPAs0bwLjn6+OBKFNogmAcW3gol9HU5rHg49JeHx4ZOuzGP9Rlqso7MLKG/o
isIYtZ7C/Mj6VXtCE3BUR0g7GuqfMvH8oelvVg5UXSjfeLKSgcANzFQLN8sdOPWr
g4JUiIcnZf1vXtApDYDXJBiw688bCtE+0XeIllDhhyQ579gSfRRmyAPal+YAvjcD
6oskYgZVYtEAHL1tRXgykfRQi2Dm2jeHCr6fWq+lshwtrGHbz8AtrT2IGhMz8bCk
4LOdp3bIMTJxCNSzpJ4TvXIw7iDuI4ayIdyxaRVVbSNNCyifXmovzCKdt7KsWucR
7hXfUBMOsz0wPu5Jv+Xcb/r/an+Qa8ha2w4nmDou7OAjYKUTIVvcYsuJ1TWqUDBi
R7fyBnCRH1MnXlY3NveOfb5Pewgx6j07kR3WL0c3OlwGPA4PV/EAZkRUd8dCfNP+
HV+RLx0cv7WMOXS5Z7AFeDztaL0m6q9U97GwEF8dPYiVh9fZr+H0R6n19T4X82D8
23F3bOHmq9F14J5YWPO+1Pk8xu+fSFHyplj81hYQzPyrFem8jZhFMXlG1zFWcWKk
cGpEMFws94WasUsrm8e9CoEjv397L/dythfmJCuj6MCD+E9Pl1Est7RqZRy+MBok
qlAM8ByuuIIJ3ctNn8nRrbcv8iRXmb9rRzKnuV8vncWKvoW4m1EuEoD/0wBWGub5
GLSiVmLB90vAA+1jEMl0ugjAqrXXGoadahbvZHGO9oPJXoIEaHkkJ9tQO8LVoESM
uYnbwKfKktTJdyUhfDe7FFJeXxbIsjZsU2C7qkqzJ5JQuMJbH6mhLgOUJObTwUEy
YYdYz0wC8AgNQFw0s6XUdrAuQN9t+VsLLEl1YISJsz5SDw1qXAt9eSzrXomT+HHu
EPQEw4rLLgnqKNZUJ0hCQmmqtxXVdgIbqYOpF9FZaZd2JSSloc6q7qY7HnrF8BOj
rdcGgIGRmbigw9bSF5ZRUVEStvnINobcSr7+Pwz98zXO+vp7x1eEqMRbRwPGVAXF
Pt7QAum3N4UR782QLEKwwq7JAsVv/o9GTs9jPkOxb4GE9FD/mNfDcBE98IdhTU5U
T5oZh3MUp5Yh85/y6qdc+HQ2I4jKw/D9sjLv5/dLnv77SgZ9NThowihe+UYu4c2t
BVP0mnELll9BZ4xHk9qgYRnBt801itMhg/Fjjw1tUM5UWtmMDc7aqHlTzLHPHJhg
3Kcev/eWkOo/CUX23KRjWIOqqZggbdROwdpioNskAY/dTiLyEiMAxNHEZ8GnK2Nj
L2fHjcVSGvWAbeSwcidBxxUSG5SsdlIAbB8W3Ob8d53DCqxgzfnc7+K6xynI4CdB
h57bJLfL0OHL3VbxDZ65xptQrRtuEE1TnGGwSKMuNeABlQmvvif9W0SAl7822Sym
3zPSWp5B+gevsVYUaUcM+0QDvIsGcnh826nVjnUIcqdbzSUa+Wamv0DOIt0T5TeQ
IngxDZBpM08TbjbCSYgdDaGNaWWXYVsKqxIIH4jneK1qqH7TdRQVuxhwHU4V3caN
ReO0msYFAT3o/9iAwIMjUM/8XDKueQzI5gU2ZOiQK1QH8yIe9IWonKBZ1DgeORpY
HX2Y6cXJw4kdlOz7qYmxNWk0vrQsMmuY+2+YCM2ZBzDLRxdnJg4zYhSHo2jQFDw/
FO/hbNHRSexRHJfA6nt5hIZrMtnZ0N2h9D8HLUZ/j9e4PXC9gw8jgeqdnJ2/OEss
CIn3JYJ51IvRS8/ipOGtreUTuldyeidm9L3mHH3PDKHaPAS0eqDzVE1WCXrJ3qoz
/yEuODrgjcOQBEzH2vTaZwYgjXM8rztj54fHk+E29XZlZhFCECExNJTOY1T0CsHu
XSJ7eh4WKztn7L1uK8aPO6rvr+eVchsbm7bVkDeG98HNTyebEVLoHJXYfneNRcPk
BbsSjAyNgeS14OK4A6chEo7UUPzKN9WuY2Rp4wgbcTcRkmibuvdPkHuS0PqmPDIR
ihEZ71Fqwp3/sK9mZZ2WtKcj36lAuS3QlYkV7Mr3a9f5KIWqFs/UwYJ+rA86iMar
10Mkhe98RrXkft2k19n/SwAFrIyh1/AHMQkZTI8XcOPkHDWHQjrMuzZ9EnKwcUR/
Tzqqz72t5G0oUGkw3iLIe/WqUcE+K4ZvEZWbEQTRlFLAbTZByfzex6V9fsDrsBsx
AfBQ6iK1BqASzAvGnlKdw1xnej6kWX0UrwT0W1UU5RRWfwYB4IM1XOyrJN4s868Y
ViBki0ENf2OHQUhn+u362kaJEOnEojSNBhXwWDRvNrOYvTuKamiKxxTEctd9ud9q
IepnlgiTL2JTwTuxvqeHlMmeQGkxG3ZGz6VudVvWtvm5xC+M+wp/MznzWrRpV9g4
AV2tuQbLw2ssyTpt+dGmRPyOtEEBREyVXqIn9xEIkWsOY4HRs+pXM1pcrwIZKKsG
fZAICBpNMUCzOlZApgZBsKgSY6VgYqi/Hi52lCuckhCsB+GXxJKieCbEQzzEdY0k
YA6Y8hoS9Pe+7t5szGlxFSeY3B9DgbZ1MbNFmZZtVvTZ4SbqBm9FlehPmU9mYqBg
l3/yDNgXMTAUiEpmMJxIuy9pUn+DAD9WYnR1I14T/DmKjrljJrIDdApY6Dp4ZdDQ
F/BJN4yzSLLIY2BB05ORRF9H4aG73cbYuSoz3eUZsHPckzNQTF6AoHZbZ2eFkXQt
rhZIidLrvZP7/7QTUZ59L+RTamONNDtPWuQyS5OcFO8ErwKu1MwDFRuXLOJvA3VG
Y9uE7Q/VOoP6ZS9uQKlTka5qcMdHDt4oQaeUPD4AssYiQpiRnekbUdnUivk1hnzS
5NWrkQs/ADFfsRsln68ZARVevpKSQdOXiqkF+4pL+EbEq5BgbbqXj0+ot71S7CgG
6y1abkFspKzq9shYtBon+H32rVpIOxXq13qm7K22I6Ubr6QuUzIONA5p7t92zYAQ
0Z7xSPzmHtz7X5ZqhGFvMx+5wJPEwM5FWVY/6ZV2Ij7hlAx4axQzUoZ4C6x4zVn9
kZYlgIQq+GXJurv94xYdHqhDLdsjJHao+CumFrRmZql3UM6VX65hCRpdHUwVEx4g
Uo1ZOxN9YdsE/CxDCCSifEl4chMaNPgaUfeU6jY0oo/0f5HusSGg+gxHl28mncS3
F23NG14qISDABweF43fLGhJg/vTy6DSQWXvP7cFqCplmGcvO3LN63NyOeG9fz6ID
4+8RdoLP7QrP8Yssx3s9udz9Wi7zGO6hjwLVeFEea+mbe1ARwEPBNU+OzS4rhU7l
aZk05c+eEn6tJgcpCtH4JyHFoNaPWpB4hvPt6+XaPJzrvE0ceubSh2Iv6JB6jCEs
aqQkl/HmAT2VcXelHlUMoCyWoR5TdImHWa11uQ+4NMlvZBNyv7P8IE5Vf8nh5+BV
RD+SkL/rP7Jie5HCVbM0+D0L3BbrSsnPHnJ+CU4S0Nw7N/F8nG0qMrNgg9dIEM6Y
s/Q3Kx3wd/HfMB1abCXbrQ+joVpT8NQizzwgKB4EB3vkikrewq1HvkZ5268QMZRM
p48yb9X7yqO7jt6rkBhf2Q3Uc6YBDFKqhCsEqrQdrNPy6KTnJTs4kf/aet0YKKAB
Xl0KKhE7LU2HkbX60Mhr+HeFpSbPPfEpkfGT7v0uDHFm7e/9BeQDq8I8QfNZEVRk
G2JABSVgc0mEVjDeDHwtHbBVATNGz11HynbHApI0Ly8XPuNgsP4hYEh63Ivqv+NB
DPJTDvHv9rkhjiSopsc+8iIPA2OJlpyQ7IwBaIlQ1VHG5pkCM29qsAA2maO5qkFW
+99e6I+lZ2pQmRil+CBC4H9zJT26NOameMqZMz4zOhl1quTRvRuZXnSsCtRRIq/u
rHtPhv7f7dbJPm+lZoa4ulbCLQXJ1v0OkJKazTHU/4Htxmw9BGn7fKVCAqa46kX/
r5CxatNQFEJna5YTP4LrkxGUHolUYxqJU0ydw0PDn7L82c7Ltvjw0e0c+wCLSY8t
Mf9QaPsXtSheXYUh9KhS53pDYK70KGHAuyMQi1/u9TQH08YxtjKyLMHo1sQOE6cm
Mxiw8L0pMdLvSOsB4rDUKnsmWfaPRcdpMaS45bLfmnNSYCCN+DhPGtzCqo0RsChQ
pIOLtcdmHxDRkOZVU5jdHgZmfNqhRTWsq4d5pI+CDvTNP0rHA+wlaJZzeBHiX9gh
c27K3Y9BOi/yz3P4OM7WjVb3C9SRsChed+qExxf8YlNk38ctpnM7BdAhHj4O+S2o
yPRpjjMSTYQh45cNL219yyUmxcrunlMvaye1wzvgt0mYPVBFQ30kd/nASNlYghqr
pZjMGtJmM3I9UaBB1z+11FdqwXY9fYUEkbNNb6uKBKnqilpFp5tw3+HlZSL2LzWZ
nLb4Lx8HiTnjcX46c98m9xwlzWvm60Obx2gbuGSZwguwSgU5Wbot+lbfx36gsCvV
kBZ1nR26vS5lrsVJBoGFZf7vl5/KOo1EiilaNwsN1pWM/SuhB1ycOHpTEkZCgvP4
3rGj+48BYslxD6qlWeccGCC7Q6m+DLt8amQZhPRvesIvGgqaHSg84EvtfS8Hsbfd
ye8UA5ZZJu6FColrjxyJ8GZXd1iPTwWj4Je4ynmL/xgLjaJCoQTMafwzz0rNaKyQ
bJasIvW9RnV0p7Ymbgjk2/L/hnQOvcBrpIXzzfikxIhVqx5nw+RJx47u1yIgl43o
WGvZpn0U48DExpw5AxnrtxK2+4HbKkD4L21JdLH1t6YYYqK6dJV0dqTPvj01K2GM
HvrcU+YJeGoheeWMexRGvfrlpIHQwYjPhz+aatAtzW+k8ze8qAO5KMXYJzhB6LDo
MlOvLQLdOrU9lpv8k3JD4lHuib35kgyp1katUY9J2pbYsygMI8PU4nl4GkCUhjaM
B4dCbpFcujN32CajDrNSbpM4bQHQr2ry1Zm2qEqo9KWLXuwIQmAjFn5Wy8KtJPiA
dOOn+G2OFfpB0bh7pTKszatNYplJjf/kB6UAtzLX+NKV7YbwUO/4QYVs5ouiwJA4
XQfEwbWkh2N/LCtAkUQHWu+vB7nJBUmRSbhXTdq+R5pdp+NcoVQ/9qLobzExMK7c
i59XXowMqVdS0mxGA5O6I57OLrn3AhRDyM4AJpo+GXBd8nRA3Al/RBS5KLryoJpR
9RXOJZp709WNFyYfpwsfcGZZBx2BHsoXTbFK+nv6UyBzOE4/1+zSRi09guhcADgb
ZcFnR1S4DKWE+/Dpju/H3gk79XXKZRa7GlZIUpUyPIJAP5hTBzObnMlHVSbB8WuG
6DIsLimlN1vkt/2P+bTPJZw6aES0eFJKjykXs7AtEIgAyIbZ1e4IdEhgN2zJ8EyA
YNuv9cS4E47afKvXxF2LzIOeSC0P5vy8JIIoG5y50g4ZQ/I6EAGkzn4cxSP4F8FX
5FCdy01/VNGyy1ZVbx+TUVoopfYWZH4TKdJP4cdsGDAvMo2chhHhFbXP049VNooN
gReP2u3Sam6l6lFz8bLJ4Xbrgo8ChbKMplneGrtoe0tCE/2J80ueudVE0guj0Jv4
mHWXAEoMU/ztE/kepBvpjb82boMy/Snwqg5WO3fpQOY2nycEKVEGi5HdL05izbYP
PwaZXOoSLfmyinucUh9q+kufUC/AwLUn8GTPaG/tYz21/Gl7QXJ4d49JQqa3FyoR
AP8aRomGffg1peGiQQVkxvnTH6v7HtjdOZVBzTWrDg2FcHr7ryz0dtm/pDoSKTFP
fzojtwdfKWNQ8bMv6KyvENj2l46rbo+xAp0eE+hZFPYZPxuDKyrjgXIQwYYRz1r6
sc6XZD2CiedXbCdcbDqz6xqNxRdNAEzVr7KmhkTfVxl5iBs/DX2yNNzHa7Spo9J6
MEjgNFnAdW0Y0dvRVRhIV1x82tIDNIeRwtdWUNsHQotsHZfGUZ/j+gxAE/VcJ0fY
g6+66zytc1xUKc8+YYuUKcWmzNxNsxypDJ8ewwiE/iDLl4e/CVaDU4gDYIfjecLb
qToVjVeQjAgczyVGL5YdlNw+z/ctKFd2kvjj02zxQ5I2QfJtjWKGL6L5AfSTh18B
2kJI4HACB44jHm5B6K9kBbid2Fou1hMCTNyXOAZIyq29Jqx1xcSFTrCaSAtlN4YF
tiR8J9/jq5bYBZsRMPhT9PO0CcxqL6SIf9lw4c7/ZdoOcSmevzYOZiTIpTQSoxeh
WUrk0Zt4hcHUTY6AbD0zoODwkw+4E3GkIp782Fxg3NfLFvGAgYJpC8fOlk+KUJ20
b+XAyuspkswS/2smO6oFcS3y80PXZ4C+O6fUzMT6/x96w0r2fV+WVTJ4eoWL+jXc
u60hTWufAKmGAoFUlRP0fUe/WofjZZ/ArBddn0ASjf8usI7H2XoVkp0KBw658erQ
Z8g8g96iIPPBnq9JZQO0rlNBhfrz8IviXICVZm9oD879Z+R3Qbj5XzrULFlTvEto
35MOjTKJMv8Qpx9Hyx3SkxdKnCgkjvRUcqMMBw+hEQ38jH3y4fSHvmGQq4ins9u1
cFZfPtWB+xLI1bP7yO6OpHU38G+jqu7MX6ZGFXqPER4+GlfTflU5wrAa06fkD7MM
8R3Fkxq3igS9z+XPdzLve1ZGCfPJWTBDXlclZfS/Hilgm7JoDiOpLRNqthQzajy6
PLYBE6Ohd2AZizcBl0yz24ylohh6AsRkV1crhO4UzNeOWnl7YDZ1sn74IuSvU7xR
5nZu0Ojb3GtPumSNjyIpltFWyTTN9iqrMDYRVEd26PE9n5xuYaifQZM6OY1mHxy9
JEpFGWflteNZqdjw2polSlPdVKMLj+kYpw0/OFYzj29fY+NZB8WEpjQLrZeekNEG
e6rToiDspnmQhfMC7iFJr3CxaGjk+pPsZfnd1O9/vjI8HQYHpQ7EIbXBFXJdryiD
QYiQ8qnNxmYGMgMh3QZKTab0yZBC/wxzvH8SYfTNYRi9B9aZK/RI/5RN/u9CRuuq
sWpVNSzWOH7prjqlPcTdz1YAcgGmtK9v/350DVM9kScz+XvGXQzWQX+gdpjAHdJB
M4muK44NN8CyZshSAvSTsmTYvZSVaWjAyRMQQNXxooF0RMDPsoDxhphl4AppEyz4
Duu7J9DH5oNuNisgs+w12VUKVDg10Hi2HWqyA5wKYExBo6cHKjy23au2KxW2WHbV
rJQOeMu4pAFzXDfglmBekSXRj3CG1fx4gnSUPAylckRYd12SIlpEACRBwJ1mq+Ix
fK/HkvTq7zJcokqGzhdm7NTZY5aol85zI+MoqrFXfUkNfZtWcQRUun7tAaSkyykb
ibsJec30I9dO9OP7X9YlY/6nxHSkaP2LTekSvGjZ/lV8d/wa4XxgWy0G4TvOEYGW
dXAsbSd4DhIqxHcCnfnxD/dSocY/5NIrAt87R5JTZF3dudRE5bPyDrcOdVVsKydR
ImN4AZ2/PbH03oIon+aA48vNaZcv+kS3HYwd29PLPPPMjFonv6kvoCOQn6tIKcZj
axQQfUgm02YlAAoJHLjjZc29jKaSyVExY7tpgE6nit3I3SNd8tW9eSpnceH+bD53
rztG/H531XIQs3+TwH1MnV7W96EgH+5ffwiQF9ROHqV8gy2EzIoeFHHaFb/LoQ7o
OdTdeP8Q0qz4IL3a5OYSHnOpYlPGIcCjbdLBXCzjrY5gY3i48NJoq9AateLOO7pv
nzeCo72Dvfm7b1c/zNnErTOE+TvLJaLxOeXpLZv+m0r6wwry3pja2H60DP2BnGYe
h+WcAiF+e9nWpvCdV5FCCr4hymVJECjxZjikRP8PqgFKInF94vD2jn57wA+LvdzN
AanZw+qJ8yS3O0bUFoN2wEZDLSBLEruEsNifr6WeBrAzCQ19xxW6m/f0ilnE/p+s
JD7QP8+b2frQupkTm9pG6QsDYKFY37FDwwjTQ9pIXKf2mJjq6dYwbDAiYRaHM1g4
ynfXfhBu6FCqIy5TRc/LsmR9D18sOo/tlQbvSgHtvC1q6+ugyqw6x1+ibaNsMI2e
nfMX/Aaxcm0MIZ8GHc46dg9KYIvrB6oW2oq9yiEt/XR2j4QpzbRJTKE2XIZTpMrp
Be2NeNJRqoETXuNlporlte9oeVoCW+s5YGoIEGxQd+dLETJ1DsopDGI2WojSwRY0
JeMIG8fL0CWn8wXhrKrZjBJmT9CmN5NtOMSY+RsOEyHVFFNeGE+JZKdNAk9MkYBV
1trg9/Y4Ju3ktdXH1SAlLp7y+LiiiMcC31p4ShRGeaytEqLaVS7pTCZjVZneTvyD
I9Va/saltCnhGbgYGHaz4o0eXArJBGsai1zsk8A2taTl8XjV3+B/38TBQw0CY0NQ
9I5Hjml+G8UQyxxz6AD//1PhcSmTmqgkcmZEo7KbBOtmHLeoWSYcWj3QJukObD5z
iRUH2/uoSfZfIU8UsMjyv3Ihu9Zr8u+7w+WmXNE8J26MLxk0tMg4RWybW/u4S4Th
CFGtDGJa5E0k15Fh9Flyc1RhndQFAjjSfxmMjDtAl34KIJJUnyTVnklD2VrYOA6U
hMMhpwB2uI06E/C7zqUlUXn86pfgpJc1EU9/QGd71fkazI6GzMoJ82Rmvbh37TYc
f/FVmFroSeQx847jCQfaYDx8R2d+AmqkyKWh1Z1pX2K6EpwM9DDoFvrmK4cuEOll
thTAWJLqi8EEoMtZoFJaWSbgqYFXrWpfLoEN+tgxm8bxHu+AATv9EGfeFrh8dkMG
LkMMk8XCNqmG5VItPzWbZRFAyYoP7YddbykAFhlAwm5LnbXukfWUuj+fAjmPUgxw
caEXEnwUkHE9ZXfZ4RTE+7p9trtgzA9HURwMyyJVNj+UCZD3zpGEGwQKzW63ezF6
w48xjHZaNqJD4xvaSyIHwhzRuB7PEFUBd0QsLlDpfS7/zzb6oxfJDCkMhzwixF7k
joa0vf6adITIJj+YNiwrH9oSLtas28z14lfiWeEkgmAX26lvshyMhbWMVVKgVGEY
2gjeJAXUXlvnYV1TZ9fda8/K45c4YDHmx/+/G+xyGFUe/HMVGL+fGkggPpXlNouY
+9VuSbBPgHlOotR7klIIPknQT84wJnaNuXwPTYSGw+S/sz3tSqs559W/owC0GA0v
AnZS0NFHNZbpDJAyg6if9bilCkC/jnEf3zkD1p9+Yw9HoWLYCWtq55W1dkVOHV03
OXyytSXwK4IRbwQqZDlrT6K/cXCZCCPOC8zvC7TbeFMGZK0fbHDh3qwRqyA4JUWh
CMzMCsx4yXJ/D1G155O73iDgVZqlc5v5EWE3RXjEKIQQ1Jx1qT/p7PojbTER9xB3
IWBDMb6+c4hRw+MwDxulyoPMEAsGgZczTOyHuflKdW7W6tBhRWPnSiJbsYrmOEXb
aU8Vhcqoigo2i4VuGSLZovS0wSQrGWnkmaFt2pl4osi/rFipD/xO0I2fA6qtof+e
9q7USnwWdOHEI7h54N2LzsH1jeCz2LLeuwJILh/o33aQwInEWTkpf5ij0Tvr3Bnj
KJ2xLLsha7ULVhYaPD6c7hTr0ZxgitnfcaHqSesS1mvUx/vbdlsIibKfh7BJA15E
1ct8sEsDL8kK1HF7Re9+Oozwxk+4LCQbZcCYQHBBfO0tCfstiZzknmhoaA6ovJIR
VGq1aM29aCCNCqu5f6hasaV6+V+YYsYNmpmkh4XzPJ1BBEftedfdh35/zmVpVbiy
iFggVJMGU5q+Swr6tKOXajHUzyPXYedvW+9T/so+spTUpDV2iwXXjc7TMbLCCaac
K/teDTulka65PG8U7jjXoJtDCMoe9WnlEL4QK5stIntQLzodKXxMBSygpQtnjr0X
nbQZ9hAS4iYBJLa+mZ+kKtRdH3bRtegB6pjIHPbK0p0r+CndXAAkwr9RpIwo2fYM
BA2eZmcf0sbgG8JYrofH6ctAhtQ6e0D+HbYqAA0RpdvK/EWQZElg5EQ14JVcuW9R
31OpNqnO3021DKRKBbZNtj62bDqsFJTBd/CkCPrA4TxW63KlUNdIGNToz4lGF316
3HTzX0GIAAAPFCXsm23+nGmBfd+U0SOIEH2J2cfpEXAtRsm6CyMMTIKuUJf0Ns+K
XWnym39ENoq5QkNLUf362PnmpQSWydnR6G9NP7wNwdcuyn6Bg+t/widvzkUFc0oj
/WMezUAnbcZSYiSF8Auz9SAsje92AOduaMp81oX3iwdY7+JhnaFNvWFY0Vkfm2Eg
Emr8x6+A4J1HASI2fU0dM3IHPyiZWX2jfCIDjDaCE26j7a5J7zlb0D0lm8NO9NC7
0qLxc9UbJoP3o00UdHNEgAeyV8/CbwJJABc/HolzlIzRZyBZ2ptRVa1wWMxtkjPR
hk4VIxmqhv80zw6gKdeWugPMpmU4UMbXY4DnD1kuFQJ4Ytvy4+WSiGLPumQItuRd
BVfWVAheRTzRMqecfXRY02VpMYweaqt/GNiswgNblD9oz3tRAbpJNBtZo2wSlxG5
Ex/ZQ+yKkQHZ/kn7lDSOrKmTa8PKKAJmcWXW0NqSa+59tDk6IgCmWzkiGHsSW74a
PTKHpszEPMPXis+9DMnnbhVueT9M1gt/uQB5TOYahMLul0SE8JAa6wtiEad9Cd+W
L9O24663QjKZam/dRwDEp8mBDRjX1/kPsoJ5/rGGOKuGfw6j9HmX16m/oNWyMS4R
b/wV4sU6u7pvQjL0rBUx6766yQ5JxHGzAkXrbOjTcyuuNg8+Iu7ElS/hZxNsKawc
GTmGprUtvp414GKlm4orpJvyHNYhSCyG8PcwAAWVy1AvKBpcguda2WTP9DLOepnC
6xdvVW4CmvPdTmtLH5cchFEa9qqp24J/bGph6566SRkNiM0y7DmIHZSQHPi7QDTq
7rN0mVa/+c0dRNTuhI/UlvFyF6mc23hZVd6aE3czX5i5yrR8/PStXnmWbiKVn2kI
QuUOcWhBL7CccpQp7TJMQJNB/Foe6gpYK6G82Cx0Zg6+jS+vkCy2lyu8zW5VHnyk
Iz79N+AwGmORE2lO0kW1BCfUqaAdmYxFtvUcARWOPtkPSm6hHDWXNpVlEPU0z6W7
z10FzoERbo1mNGOJLM+AzLZntI0BOXAGevJ9w7TnnugP8+cAOs1AseTLxhGvm6cs
LFD8dKcpIo8YwXMgfShJsYUMXNY9SWNhNO+eOE8b7Z8O9cufP/9H6LG0MzJePFAP
OY4tSuqfuUFN7W51gCW1E0aecdI1zhtksiBL908/km5biTAlODwUXdsegT3vKlMy
sjxXSDt8HM0TNCJSyFaWu6BawdVI/D4WtTfbQ7ixgCU2Oy90n6kDZDbHo8vy3sLT
MADK2ZGKoW2vyoJsRVIP+YD74duvqiNytHD3hN7y0JbNq0Z4KtLAA9zm7EXe92zT
POzK/M6eOtf/kz72yeZZL/jXo1PSOs0Licz0dZq4A+6fg0mP2qYT/KhlA+T0N6R0
tOHBlIRB2uVwHmKUOSI9ZGHw7KPrh/Bh2LWKuihDors+l0oELcvfyk5pETRSe8Rr
AfVCQvjaiabkJdLyZYK1uRXVkRvnhdsiXWqNiMaur3mk1q9rSRQFbExjohkCDNcX
oEkZ08hvjK4D5tR5qudj+/WS7xXfZK1UijE5LCzDLAedSX1dFIpIUSA5rCOzK7z6
8dr3wubIZ15XYCNYyBi+ULg7QmsCEpIcz3LDB2J21AwvUvW/5IE5OAEMz1/OmGVr
CwV06Pq+ePfs/KNths1Astm1+LyYhOfKvu4JITIq+EVj7wYfIRaWBSucL3kQEqRT
mUmbN92F0t9bCABoeldrdl8YCQ7amV8vE12sH6T8ZbmVc7USf9vEKpY9ebk2KUp5
0T+R8IMM1frh0gUOWAaTWDwwY3a0g/cuqF1lKUMytxkTmZ6O9P9jyDubpOPaazJz
dYoUDTuVhUVX7ZL6IkSGumiI4yoercfjfT1R2Ug0CdPI6OkUEu1aK6YTdMZIfpBc
vl89HVCrSlAiHJxNlRCJblr6sX3mJuAHNRVBEY6ISp4aekT2N/949UeJItZhRTA0
NSLNnI8KrZ0e9w1fvyfoWrED1pTg0cjRg42EBTFoEwbLFUhFKUi/IQX3+Ccn4g8w
A0+3aajqX/m4zvOqyRIUTmNt94fHrzxgwmdqKeZVmvDHxwtSo7T5qhL3v41bGms5
PVg7q1ExdAB8jUR7OwjUtfNLre4Eg1+rOTFLHloNrZsA+MoJB6mmqF41m8BJbBkS
5j8qZYyqBS8o3p027C3rO24d6kBLujMjAoAfKYknopnvbV4hnc0KWy8L86Puegqt
kJMsevQNViZWsSyTUcgt/4XzzVJQjgk65a9lJ4MgwLIEWmwD1Erm2NQdMsyUIYhP
Bmy8RWpOQlJq3DK3n0ZOa7dbW89X+j893fABX1t0S480/y6GSKPJ/DuT4WuAKrVR
p/z8fxmaCPSDrdR45VspfDofXo5jpjvwSfogvh6rCzx5S7fruwP88WlmiL/BydGu
MPbF5gC/UkDoo8/L6URxeHFXWw+p2ovhtr7OYoQeYlk4QHc93+rNfL3HV6LftQ0B
d1jC4M2u47RMUhlnYq/gPAcEp+L045SSc2KNuBHSJuKKsXhysfAvz3q5W9mkHkWm
ayJgFcaYadAj4zX3zotO99/IkO0FHsq6smLOeYouo9LvnY9ZjBRIMgVU8mWijNd4
S5dvCOG7O9+jiSYvY9pQQHB38QVJ/4EKwzJ2g+4NRzQAS24V1qxYj02YwbSf4/0A
JYS9/3+qxe34bJCBIaxTY4E9dzeEFHTHz7xgJrA15D60HMo9SniGVuDOxxLcMleD
ajdoDgTDhsx0m/pvEmaTULTW83dEJbeFTkv+E6e+j/y5a8r8FyTMyyxGdVDhvrW9
ebBa/fOt9VXcuAPwh0HBYcOTa619MhOINLpGIcIgVidzJ6M32inIPFZFUs59sqSr
viDJv1b+g7ADyw9qK9uZK6m9pxN8S6IAnutqpudkAli8QwlQbthyOjY4NO/i0RSj
ctRhzUrnL6eUetp1685uOECFLnWU1OwYH374bP/2WJ3FCw3g3TMWthq+mIVwEbFc
6WV2isTXbgG0biwHeKVl5/ZEBu684N6N7Ee9kpaMciRybYoBgUnNN4HKQqnPmnLb
8lAxHahBRzji8NyYHF4QGrG6E9tvjURXQ94MPZxt1xmXQVxlQdliOH2qtyLBM59D
n8MFwyX/fIRFhZXzS1kmgrP/YirGgShaQVbUCKzuMxqqIhOEErYBv223wXOzKP5j
X5o1xibTIzIPZ71A2ujXtAeYe9ca/NDPwrxLlhmHSIcGF32gz5b6dogFnb/FQLtt
SczTQfz6KUD3fltQHtwsdgtCnD6N3nEwXuavcIGo4bLmjAcP9wikm1kw/XAX14Ts
pGeV03kM5/JqmfT7YUsxItDO/GQ4fUmMwuWul8S6ml4Qkk50WRJRemoSRreVmEih
pOER+aVW44DBYwR/yrv6YQ1L++JZJdu9uzj5vh+14YA=
`pragma protect end_protected
