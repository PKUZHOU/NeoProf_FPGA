// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ND5QnbobLq27ntG0z/oy2rSYThPMRgQICQpKBNvm6FearoNps6BUUvFwZTgL
1sRvqV4ZhEDogu70GP8MCab0oOAz2qi1YAjb6Ld1RR6AzOVNHAcGpn5iKs2H
byvJf/2EvJpDeLfXFd9jyGpkAQWhQQtFeueDu/IO1ijY5tOnxHLqlf+sVfSC
gVbIWUvZtO6xKKSCD81gAlPLNazLcgaAz5USKnxyA7Dm6AivK9gWGycgioOe
vGqLUWqXgvLj3c2kDcRn6mGdSrsTAsrHIEjALmbwHZ9/c5kechLQNB3XFeSA
zcDoHHdLYkSg6T1gDkVOiYo2CiwQyMUzZeRKzH1xSg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UgFTnpHUnBbyLjNTHXxxeihdUAqMgX8nWEj0Xwz0SVRgZ71X2LmM0ms9IQ9F
eRHBSKE9NHZ+UNJ7uSxwRCzTI/dUFPs082tNBaFa5qmSm2kk0paZ9evE/u4+
XL0M9fhOi3OIr0oFneuWMVzbzC0eyqGsxjWSRHHoRzJt/X0AGuPlI0tNNA3j
F7LLaXm5m1bY9J2CxZvjZ7HMWUaT32y5lWF+3wohPZmKnadHuk4QuacL2KsP
f9YUlK66Se07JAhlst8Uu66uhPvHKa7KtgDr9G36wgJOsEYbtL7C5mLNJrdp
4SeGkbbYWmzd8uzlqwFUlANM3BGSRQD12yNvlw8ajQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iaDUmppUWUebQJo2z5ADKLl7ZpcVofqbYcbpJxRZ6xam4BsG7LURwZa+X4P6
RIGOCUwg15qDfVlG3O4EQ99p3QogGWZgl1DeS5gjROkU8kNWdZ90T40RBRcm
eLkP6OxlONq75sz/GQ3ub8bSwCVl0i+d31w4ecYhZ+B79mB2+Ixo4b++UV32
KQeUK2AWBlaKLVwtlhNx64tjH2VaXZK+gPUBWZ3K1QGMt9t6QXK1l0vlxXbb
FvDgSwdpHvAxC88Rp4pQ9urqWZxfmh7hFH2yOUlVrCxRP3r/MOlNyaGdA5H1
pqTQ+yR41fZwR2imDyK7IX8DrVoVkkTQTObboqIqgQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ovA+IhEpzB3XLrHoRY6yd2a+OeZVPucu6lAof8ncTKf6xmQQpPOiiW96qWRH
GfNukj1ukfddQFsuSiDNdtC1E6BIWMk8DA5qjCuYQCCRgTfwiyTdRovzu2E8
Tnd35XYcnFelnrUy9F0bxpZsb7fMEWBGXLwKl3y03N9YL+FQr40=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
TCHDHAFYltNu+YdYr5YCnxpin/M8BcTXH2SroleNUbf22zmNxz+mXegmr/0P
cEkhOmU19PtXfbo5Exad1twIRjlrx7UKhFuExu6a3tsbMpJ7uo9MUmtCDNvr
eMZLYwAegNN0eFLcNnpPwn6x6EzRGJGD7aBnY3lj9bjgA5EOMpUeVOSCfpuP
iWGTfZEGrcLCz+VALjsTb1werBkwKHlhA/6R88SNu5xsqNwuTPqYBATVPkNK
7BcTamZrPA+aFLnbghB/nN3tjMFpOpVBzDbxubJWQEZGCEZrGH+P0Ut0tfET
SnY8oh5NRzbNWbmP/Uso0LJK8fEJYK+zp/vBxIUiU7FJvuKTyPUAJje0DeSa
TQNX7Q+UyXIZsIxgotaQ5rHve1m8yPpWsOpNjrwRKh3AcFdjfLk6aqnfMGy2
Wdzs2EMmX1KqFbACtYarvl6nr4TbQbHcuHx16f+ZFLK4a20kY5ZffUd2dYMb
8Tuvzg8dZ8iArY+F5ImESEhAWCXVVYZZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NoxUnFjKYrlnptU29gMkHzJYjxd10msnm471fDTL+VesB3JfEUPo7WUYyeMc
ANTubVQ9OJWE98QxYIYYu1ORtAd8m9cfiMRwmLcAJJ54GKfBF4g1fv6eMhDm
nDojTBeCmq9jBo0zEOY2wdsEjLeCD90/+bgmF4GFOGloGfANgpU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mfsBk677JuNlGQ0hyQ0uVRn8YAOEE+DJO4aA/pJbIu9ohXwoiM2j2/EZ+daA
OHv/cGgIT39G5yQT4lAewXFyBcQMcqLpTCXc5GEiCLKEPpVJbbTUCLIqwaum
cTJ6Lv0jQc2P2zK9lsfxcsscjRuHIiJx+nYEY+QIgVFldsC4EDw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11488)
`pragma protect data_block
6pHICU8lVbPkw+GQu4wwuXzvbUWloVZVT/GrJ7QIoHSfwM5dy2NGmPbG0Fvi
8h8qhQzax5/qFLTV7KE5hacqgKIjEorvJhkc9iskISPZvGV02V1u07KW4+xP
AjZn7ygk5PaT19v4Ib0pLo1BLprrf9zcaTANA6WamYNRMKGUoUUeGXHnSl18
rzYABuhyrsnf86EraNzgh8I6pVxnj+RoQu3pSFE92KqlChZGm0qWsY7NKlc+
b5iFtTSnGKHV1fcWZ/7+zUiwNtWhLIJXaUJWVMzKdzuchQafKsKf6sNnvHfc
APoHRXrhwIk6rh3ICLBwGo5PitZYoRmJuTEx30yHP2M0Ua51hLF1C/q/ZK4s
h8er0IvzurAhocJ+AwkvpDiOwB7psYOvpHihuYDlkQOZAjshmGmjziEjTnL3
wVSNXfLCxxNOaxqspaOtGtiEyr4XZzg45NAx+MpUzD1mopqtk9gGXJLeq5tY
qL+itbomd2QOl7etsQ81Za03IPeVos1TVkg1nVyQvXK9G55l/nxntXIJi+rQ
1mziIWp9NW1g/46E+JghLNyNIkBDBWDBCQdWpt8YR45tfGciBBVY4r2mCqXm
yUOcJHIC9plYd98JpIaW6r8eYzUOPxO2n49qf6JGqrDuYxsPaUoWZ+42eRjV
g5WBxuFcNdNJVh3CALxEFnj9fainGtgyawXMEo7Rfm/9Y1/xf1s3FTPnA4uT
t0uzwsMjeVDgiGl8XUGQAH7+UIcBUMGyOQIuu4LHbjkyVjgU8fn4C+nGeUFI
B8lJPvs8nghv9KgRSMB1nrjLXuIZIbo7lB/qdFSMvU3fs2EnnhVgDvAcJSfL
EM6wcU+/njdGOcp1c5/uoiTyzdXpwOr+ZvI8PIEsV5DJyHI6hjr/m9brsGG1
lqYeptOtaW90a2I2G5/TLrGbMSb9SWemI/si7wwQb7+Om1b68SerhCPCTMvP
1+kZ8ec3Llbq6L2FKiUZdPQoXtaELTeBlx9wxTbqfTq66pYSCzah/T7EnVec
BaPaB81gze52bnRtz2tavNSszNgp5gMskN1FQMcGANUZyxKU48pW/3VXxDC4
rEvm8O+gOVmMpuBRMQqhzFkVlwEj86bjNEKe/aGRTr+y3YfcIgdUArN9JTfj
op8Z/nd1rcB8nDclwHHvQhevdyWEUiKUmU+p6EtbOO5ScrQwetU7r/nVSyAC
a8Sbqaf8d3Uue2kKHKLTs4IEfkhZ7Exo0tgKrICXX+R9xDPJFJjCI7qFljSH
F4ulA0dmoMhdzJtNrONRi5MDgOhCsdJYZhVochbjoHwJoH2RTpQCW1cP5gxJ
4RlZsPRzdJE6ZLK2nLAeknkLJFRlaCQssvYE4CxybjgEDgfZrBos9BafKoZu
6zkjwuZov+u96mjxveBvfKqk494Y1sfZrmvsXV9R3Zp0EkSt82C0IDoMMdVT
RjBNRXFo1z5Z95bMjKwDieYjL4mcYeOQxdf0anTYHyy+YQVhRdMeuwUSE7b0
U4gsjSFNl/w4gr0kDaQgS1RFRe2lvFue75IbAIAH4z42aBxWFqtMl2f5ExWU
mckGXCTNpDvjlSHEbiR9GslY0Tf53ukS/OaAtKOmhGbUkoroJfbC6fGOd3Kk
6PTaG2gUyae5F1GXl9obJlbGe8TGa+hd3Z7otMReD10p26gEssNzG5cpmloq
FERHpXko6GhE4e1vpfN4zm7U6SemhfSxqr9A01gB1IeCyaakDQWnuapo0FqT
mzOr75JWgm5UOmjXjrA9Wwn9UhJybPBoa7l48SWUY7j2jhRCpsMyDjW/muuC
8qZajW2c+0Hk3IvniSoej2LXrjSxxGwjK+so4Yw4y4Ap7+Ze9ewoVLM+1Z+a
xWBkZIoSKSvDiNhRMF/DEBxIg67cu/GFpmK22497+AivkcI3bQjA0ucPr7z8
7/aIU9pe5GFJBN7pMcGcowJAHsKZSXr7h3YC2KzR+4JqvlQnm4IzcRGmYt/T
N36FRst8P5kkUDOwW1upI3jTEnnfZVbKdbN1LHybJ/8Uc5ENGjQK2Vpmg8D8
Y4GU/2JhhSpFuTwOZYa7TJQiECK5rgyBrQA+vMebS4EPSidF04Sf64PxmxSf
3Bc35H/sfuhewDReZXsMFeMAD+Gd2g4C5i0mccefFZYQrzJvo4NEDaAZ34+J
1ndf/p1wQW55j/VYinZ0EUcL1+GXpJRRbNLkQumKlBKdM2WwtgJfHNoEu311
VphjAGCl8GO0KolnSalqPtCWpcwaHdUTy7iskpH0mS1a5RYfKxcT4+nhhoYS
H/XaWt8XEjtlx46jXKMF6AXH3fLp7EOn+AsPBylLFnioBQ7Rgc7UAG3a9OrB
9GZLUoOrkCR3cusijNxIzPoQSZBmw+DME1Nwcj2SjPF1AMvxnWftMTy87au5
xSiTEnW3Fn9HpE/fo2q490UpdNK/uKeZZcQQWCPsYzEMaDQIQArP951ZVLDm
I5tDR4DYJjRfhWuG6fsZj9OzEhpXZnCin950qJ7JUf1MPFqW04C3ICQoeOhx
Kl9ucsa4nZUZTJmEbt42DnSB9/cv0rtzuOLHEtyO2SdforxBu8c6ai4TTIwC
pGeZEMDdfp+Z8DNKkXJnJ302b4wIu4Stro446PslozrS0ywjJJm6UHNkD4DJ
M/X+z+E2Ik8dqPpJ10u9BvI0L6uZUwuiVXEtXX0zdSRkmsoo1O86dFsKIe/m
797ql7DxSeAmVyV5O3WgdDKvgamtH3HM0JLS9nrB726ktpiAzq/0ASFbcys+
kTMMT6ZkSXxLnAKKNOvmICMsFQKqXTQEcRA4eMIopKQazcQwLdw5BLw87PJF
UTZ5iweSPDuZDwtBq13W+zg+2W9oXgJVn/R3rYDxMChEzgTZnpNMeZ7wtdqv
V/ta+JCim7ixOMdG2WZNcxvg3DqkuyKDy2+zRzW4qv/50p0i2+Cyr0pM9Jss
biA1qVZuF8ailvvEfhtkQ3iyipFQqqyxkOB0aVxlH8YbLASmBi1Z/v7iu2C1
u389+FOZnDm7FgZQ219c6hmYzgK0Xvv7gn/tuBRyERqAGyrqJudLq9TmKZ8b
vRwLH1iFu7CKqcSieOz1HeV1XvIV/1TejOVOeIvLzYt+r7EQ6QyAn4yVrMgc
gLRDE9z1MRmW0R2sg40swgiDP2Uz51wkJgwxIEfRvvVu4XYErqDe0U53+79X
ZubOVbYVZ3pR5DX6i1Ij8bE4VHBZobvPd9i0FfcxjInzyxEpNyAwFlawdsfJ
0F6lfj0luGjWEJsbfnxj+u2HTKKYhfdoyPHGBhid7tTQg6U8+ho/GuDD+tvy
6QW1ktuGa6E31k7YzsAiCobKaDC3mR6BYP5P+Bs85n795RV3evc4kryds/N7
qYp2CIkFlM5pvT0lOeBQCg+MNf+s87f5824jaYPi0gwEeTKNfhFBEV0tQEpC
xn24psgKGBA7imNitukqZQG5WntNS9429rICz9ilG/Gu9AgN3KzHT4ZGraGO
dvl/kNCpopZnKBdIAdIDpsYCWc8Be8h+DQ2qgi6Rk05BknnAc/oWj9u0AvcO
pSivftla5NtfGYnrwOEEJHn6dwCwdebCfl/mn8MlB3WEfDKznNuvuJuwSqq8
7XXd3XZeAZSQ4GwaD2dDh591PqBvcood/LH+RJxbVCIgeEYIn3U6PWtIuvP2
pkb9R+DfloZ7I1itqcpVWnjrNDRsJCIr7BjRrOG84Xs7b7ReZ8dA2djLa9+6
Y9Krf/SCkSni9hArTWnRNejyE/iODlbmEabbnBfK5gkiXNWwSTwCOFv5YHTH
tnupRL0oZIg7p+x2UP5LbweOjHBTZ0ev7vVaH2kc8CokFLez1SvyMaJtbpga
dgYyTSrOnJc2M07iEfetcr5WTNLSE57r65RnJkflte0eb1ojA2CBXWYr2XuP
B3ZFFb69z6ZLMMdQ2BD9qAQ4sRz63NZ8tPb38bkzOUfZNvW9oFQBfwB1ECZq
HrQcVNVqio7cIHPDbYnCw64ngigjQ8RRGTiLS7PjaPLV855RvNo4PYftbK4j
Y0KNq3hE1xym4n46VQAT+Sj/odZPLdzUnZPpkHOZT4gmbgLCm7WSoi/YWbVJ
3d6DRx8YIR/dAoxiN7yXwWZFgwVNUoBzHrMWp00frCiSMqVM7mQj2EWKDtCB
TljhfJmT/JNcUKgRkrGR+8yeyBKBlDvlyM9AfONcRje2MW8WIesaEh/vyo/r
r66AXHVe+Q81B+T1Lw4b8yZNN3p3MRJEkgFm85FhRPOW7CBLe0tqKi7FSXZk
N5G1drLGUGLWrXbmDZ47kZ1tgaj6LUYHPuzYGk7ofVqZVxOdLwiDUw28P76h
n5L29Y02OEEBht8A1WmaAYHi5VIEIGG1UtdvLZyRjah+NbBiwJWZzU02sbND
ETwwnWLd8lVcxQ9GpvVBNmA8GD3iVgRsiAinQwjwclg1u9ZGuNlOPwqfOWCT
FkFDhwo1Q0eY2fBrCaovPpNOSazGao1pYZWFy1Swb9hK4IsAj2H/VRD7M/s5
/OKLdlYb4I/b6w2qQBLdfN/8CwpOMBxtLUEe+TkHeDtCQDOqwzPLyd0b1Cbm
gATUi5gjsuvRr/QHC5oU7fuwSwCxJk9hUm1KWbmK2h45qxHkeV2jhLRmpn60
SMi0bl1DmnWlfwFJgx4l2Pr/0NBByOy0ryfHQb4V5ktfKtidqWeubxErbpfs
dOLcpqGXsGdoOhK/UAEWZNjz1lSloc76CtiH1gWw91Ka76aBRU0nblEhwArz
SayMP1p3eD4W/k1y0+eXTIYO2vwc6OiTo0KKfurq5mYWS1JdNEoULG4B7+0i
YuwfPqEdO9otAqm+SJDZ1NEGaxu4iohGgT2oRVmWUNBi1GNxvbcq4WCv1VEp
CuMl2xmjnxe7O9U2NRrzyj9fKeVtevUoVYEOyHkyn/cL6xs3YSQ0VtmEvevX
NRGAUbq1Z4xO+QZOR22g4zLZkC4E/KWGW94DCitGQcThXCK4m+Opi4KU9CpT
wyhs7Q8HtMn4iQceds9+ALkJYn2eXya+5vNdoxWQ//c6/SXWKfJgt0bcZmvw
J4ocBShsNWjqZ/no50GSMdJB13kA0Qh9IRx/lvncuOPfpheWdDnLVOnM2zFw
DLW9XghRfUxyuM0WIYXt8vYVp0zSc2rrgGtswWZkUo0S/QEYJYjUiZ4zNE14
UR7C957WPeo26NiEPxDewUnUN6Bxa8H3U/IjjBKETP1kWR18OSJTPxpHPaqu
8jFXU2bg1EDLwKqub861B7voAndAHo4g1aR6pn7cM8445RHHJsdRvjuGjXGB
gHIeafaimoxTEpJe/6qoAkmdtA9EoPSAOK+CQJ14CIYvWywCIoQgTAXj6ozr
H9FlZceyTZpNvyf33CIa45+Zvpn2LOEJHItcSI9tmY0V32vMZEdPL+rlaf8p
YE1R3O9LmK9PdLBijaBP9xONKBZozva+IdWRo3iHiKOhPOlJ1NvZwKtjIZ2e
2tKcRbAqrEX8FPHFDSF99tT5keicrRoncNhZmFDUiZjl53OZ3JC7fqgw0tXg
UmuxTC0X+fF+xJ18I7L80JhlZIBnTg0Uz4Co0ztfXJPOYlJZa/n/VzaWaOQb
spMxA1/RYTEr/0Eh/aOB7HEmVLZpop3ffr1rqMidS2f1ErYUsBFX8KEDx92v
vzvxAab7VbfVJSjbycXIZgl8+oQfTA8Zqwu3VbmS26CQ0pAXt+g49IN273nj
IaiHzBYCDZ4zL4RSNLNczp9JFG/zAgJAFvU48Gi7cU5mJyReGTND1cilgaVa
W+7zfPKd8xGzst+AD2I5Fifl45yx6lRuTScbISkBbfdz7kvmhQmc7ymPgINh
hG3cOON7mWu30lLbvhfaI7iHKqv41AvrUfZXi+gArVQTjVlA7DU1W3DR3vuh
wJYwhXBtgttUUHlD3Fz3+UBUI6I9cRhqMUcnuntfpd6iFXNgztW6tkaRB5PW
WzmENUMULa7o8KPTqMNpWnZcMU35KnfDeGc73VwEVxWgj6LGTo2Ws09oAIiF
vikHSPevMJxhBJu0lqs46cewYAMIy3XZzxNxr7EdvPV9i+AiSPNqJzJ/7EXC
rqUbU3rL5f478kdyzd078w23sSuB75W3xNDRZiblSRJVd7ScGsCDa1bg/IZi
ZG/H/+cYPOOXL1aCQCj1xbULYe0N7XJXIKvvZsEWSdCe7MGVymNP9JML8fYo
9eGrT37tu0hAaOj3DsHYnXjxEj4/1kTJGWHW2T5K5WhL4n1KFIrw91TIGfcT
t2MdtOuvs3s+SwSWCmZUQTwn5w/adj4OEpbj3qSx1AlxZEOe5WzRAGi+0JUe
0LdectoylKapu//zCpjBIU8RrLebLWp0L71LxC6c/6c9rZyxw04GFKQkbubm
D+2t1RaKsxmMmV3F3RaX8ezPq4MPca3GknG0mwOtM9tclJoUQrdyRbeiDHoj
NNzSj1bJosAKbT/QhR5KSB4mnKg0J4AiX+5gPrzcfN4X7UlHcsyZHKVDOQbn
bc8r7/9XQSUqck36grvmvlFUxC1XdJwAzoBQvwsGB4mNXqUUDGmlpavA9Oyb
h+5rIbV8zbnwdg5NRUAXKDZWAAWI5IctXpESi84LbCDwh3jx2f1hUtt90gHL
Dy6/V1OmAdBLHk3xFeGoqBzirBy5yZ/57+gtf+kNirWj2aFGg6aD2PNtakq/
yccycNyWNlvbAWUsyYhfk3HVymUKdQywyeA8IDUdebFMQPE9NfvU4bfzIrAk
9fGoh/0dEUZox9HXXAr7exY2pBzaSa0QpZvKpRv0nhZYhfPGW0hAxmFEdl8Z
C3Q2DLtZVj9cJjzYgq78YXZoI2zPvhiKtHucM5wS+pVNmllLyxxci/6Pm8Ed
/e8TRRd2HwPLOE/0vmpxuAJO/cFhqa//S7Px2e9jV4EywkBzxb3hK7CzdFH8
7YxiXr8TFRmUMbVBAzaZbb4L+A/a+K+CU+DP5i8HFiiww87af6dQXzCxWa3R
0KjcPO3l/hIzz8AncWdx/7VerU5HIGDWDat9h8PNbmYQOzefFZQszzhnHjLf
kkjuppXOWsIqOAGxEsfIe0Eev6O5AoRulv7CH3vDx53kd9g1mVOM9rFEpvqh
0jVOQlzCqcXNmqb+gUqviTHdKFlSMBBrI/F6AZjBDxOzGj/YfK3VgS8VQ18H
yI6Q3yEgHgQ4N8CgJuwJA7iRCmGYhvlngaK8kErG+YsOCtCGAB/TbYB2uQLa
BrxV+P/u7Q2+f66EA0/nEcqw2lXNMeqZz0q9f3lHaDEh6GxPh6ojDzJuL2qZ
6oe/SoNooEmptHdwBojCopX95mULeggssDd0gh/fdCniYEdp2PooEEczbHNm
tO5kz8qyeSEZQQLH/hicVCXdVlj+yht+/RGM2gh6neUbeH4+YIcIw3bTesSY
HEumVcUDE/SN/dmv8fuarrPZL3qWmU+zI1bT2Ku/4qt8uP5w7WJIBLbfC+jA
Uztun/ImQEPsAP8Va4O7xMX3tyfZ0SmNG8CCB52biPa18q8qrgtMfMzURC4v
8yA1gMGbTeHtA3WrkBlEw3p6S1y//6p3GP4xM63cVFAT7ORPcVgBIAJWUDuW
sJ8czZ3gwbHfYJ/YCClFav7SS2i7sz2o9jPaMsH34cM4e06TMqReNv8oX8NT
do0V5KD1pAjleOtwjmVR4eQkKV1kqzvanf35o1hdL1XvZD//tEjpBr91jJya
DsObFNvG2J45QggDLPUb4gR4kSqbFWvOOKSO/p5rwGcxx1CLLyJF12Uvjcp3
RvmCVQ2cwI2Ru7/nM2MujKtGWlw0KO3Mdrnv+jPU8Iv9Lv738R/2kOv9l8Ku
Ndd2TuXKkTny5nsg8BwNEazMEwiQK0DNCmhuXpMS4d6ipEv0gA0SO+wN2jhU
jVuCOO0rWtrGOkHUSkuQGwg7YUjubNch9Nydr+2WdA6l2CEbKCRF1I76LsSa
Y6CqfSf29yKfvx5E4hjVO201DVkPgspSYS7VCHiNyaIykQ033hcLhFH9qli/
xD0FirNkrcMw7it+F5kMwkTjkT2wjdWCr5OCiJKaXtUe+mJWUMkOOhqvQpl1
b51GJ9692DYpNjxdZzP5nRWjvUWS6zJpeDKiXx0YHCK26KfZhSeQ8r1hLQvG
yip+hYC/i+SnOtOS4RtlxLG1GlJtX0D+8J7CT1s01liym825jbAtNSIp5BWr
nNhaEc2q3UPkovVXjrmaxGbQ8xJIoQPPuu73Z6sND8gt+ib+kYFcPbB4d+Zi
KTa764suhC5pRB3aUbpuehEeW/bA+MsgsfRtjgh0v4lvMs2YBhwdxXlI03Pv
gt+qfEFjFiXp+GgcDksJgD7STHw0EUVCDwLyZmiwZ4a55TXP3QlmjA1kSkBX
N+nr5BfrBeeM5e+tbvs749SUlZcakOzxYZ3z7MCk1KL2Jua+sU4HxXX54SxE
kY6W6He3w2Z+AL5xu8fEpWYUpnM/MoA3ImshdQtxcAJfkKyBBaUiVDv/a51t
lIkyWqPAjFx+Yv02TJy8vqCBT838m1reBRSycdskp/5HBsQFawP33ieimo+S
AU9aA55dPjUhdOojX+1LbEAIqBUNB+5D+8ZTG6ggsBqq2x4yuPdeG95Vlwg9
fdi+xor5JnXENEJiK+AOmlzTFEPaYj969/1U3s8RBYlMp0BGQrnuACIhiWHQ
WbEtpAR5MRNJXMBvtGEA4ILefHIiK5RtlI3KGjOZq4giz8LmJ5tcrTQ/Gw6Q
wJn+83UzgRNmhce5FuIUUy1xr0JsrWM0EWr3mz03hOwh1kzny2s0tTJdqVl2
v61LR+ZJellckzSGn8Y1pGrijpvxjm05KcTZI+8R3vvnD/s/+59/l54MfLeq
S+p2wziFQ69L1yrrx6h0vFoQMzUj7EVcpJyOR3Su19HEaS0ja0DhUAnbtKcC
3Er31S56Oh/sYfFEnNDa+S7JMfw9kyAsS5XDR1GCPBrN0E5wz9emy8zNg1uY
ZLQ1INsVjFmkDsx+gm5g2qPFUlO+LJXI76kWju9cVHcd7McpOeQ/2t3nCdR7
08GwRH+LTSbXVVls3GyGfAbehRkEpDjyPN3IwRNRatpPDVZj5hRaWI7OU6a4
USzNo7gGJbLNV8ZGDR6oOMoXTECI+eKYsmBf9mHvoBnuezamVmS6Ty3WSaZE
vhVyfpb6oWdZA5gArT5yafJVrHBza6UqUjHhojkujjO0JP2AeKxaR6Ky9STi
LP21nAwt+Guu9LBFmQkBaRPzcDkVpU74WUev0lwXj4aXxPTnbU7v79gLXplL
Uk8Fh4dW9+cNBU77H7oizfMAhripRSOLK1kOrgh6NHdrHVrznFhlO7y22q25
W2i3SkzW98kvWMhpOrRyErZc2ayxnAJr+1FKevW2Ojn273d8SYulDCe3lwEL
5H84dO8wwQTUfWtYK+Lguv2WYoW3dfYT40LRNOGQouPLLWu4ij0tLQ2nn8EK
lSRwa2XwnKgtY+N7L/6lTVDzSEPQMmkl8s7pgJojBLKY5ZTHy559RhdY3DrT
sZFkPfEgNioYnVCFHEM3M6DIXP/S5ud4u8OUzuqsizmrtRMXi/jNfgdivoep
wJ+ydVdjjDI7/1cGOASStBbf6oNPf6G0hEyYjPz9pwzseFD2U1jRSIewb7Xq
UVD9qgNzMKrjKa7+NALFpdQuc4QanytkfL17endSS3S/5V7fvuaG9z5a6zUU
SC5q/CY9FTiY/GDGIniDjNM6nu6p+RYDn+fuMKL4cjWIFpXuZFe2oJIFdk+d
zZJd2Qiozwb19+C2I2U4MTf93FroTocJiA/vO58JMWoz6vZb6UL0gDhQmmYP
r9K4gHRzsQX4HHmojMzRosT07KrUyJH72UiN5+HsSiWnFD8O24Ke3Y7N6y7U
wIe4sjHxI1ShCwUk6D0NMeT20iYomPY934Korb068YrT+zyU68ela6KVeNxS
MDn8EdhOyASWOqcZZcZI7Lrw/ctqCoCjIx1lc0DOiq/wNBAvlvcpzGa6jYEB
Ru9Spqj7G1UCpH6s7EVufCgUiQWUxw21OwnHCZ7FQCgVSrp8k1NAmTHGY/XO
kfgHZdGL6bwzOiuxqCRRFJWGA0c/22mhBfatTXBiPBdIONu8T0iwWxjFAUfa
bFic5ZMfTA2Aacr4GwZkV7KizVvQZMDoFlG3wrev/ejnSyvyUTakC6BngudW
dVRbozomw1CjrgMxGMbJoklqTOij2nzIDGC2Nfo49Ef/EN481Q0ry+mUMvnu
/K0X0KFgz95Ld4WmC5P4YEZTGJDWM2vJ4M/420e1j/wuxvWpYXFFGg+OKevH
6CLC5+DODshA6rDMXsbphd8bqUGbGm3AOUl2bXbLCUCTGrBn8MDFbbT6f1gD
pNsi2BBi68Xy5O/qyuLsSoV8u8JFPhsKv7Ir/5cUr/VzMCP39qqIGpkXy9j8
maYR9mnXmhwFxOj+hvRH6HMaTcV7GNXiV4ucVhmKB3rRKJ2VkpHD4QC/8VBN
MxmmNlWwKwKXh9nxV7RyWsfo9p/h+7yVoz0Lcsg5oaZcumCUPArloEUAfKML
kAaZQxVHSeHRRDGTDBQVD8CkIT2wNqSS+aZ1CHsiUGxsJ2KWIY/DS73n7nLg
rAEyq36ApkpWlCHRiirtwBzyOwnY9ktOLk17rGxiS86r34T/LcfHXA9Zx+OK
N4+gmOeTV3Leg8uIqfFFFvjhpww21QHvF44SZ69/xQU9hULBYikYALv0bFkY
8qEftw2e7dM7CmWNQPWFj9Z0dhXtvoH4p0H1ihGz3FkJNU6tk7IRxptMTkR7
xmnYX3hk93z9tq49DP0Rx2+wRcYq4WMT2A0hLKh+8+7kJ47z/SY1y4kCrpjZ
a9qAhc/Tfg8gDvB6rMHWgHvRqL8Bayw9y0eo1fLur/zuJ/KPikGYYiffM3Hz
GjTdWGdkWztTcxeAM1s5PG4/pfjR7j94sUuxDSj68ieGZ/88v/w5HwIiFt9Z
lvSgBTQIk44300iTmVc1GDXesGLg/UXuyDLK4wq/kO2Ytb374Lum9Hbzdjlv
BKDa8TfauwVudLYh2m+bDjbUunGaLDaeKT4YvkmqUlNF4iKhO27Ma2QTjMdq
kMxS8zhVCPlM2nl6NQjy961N4ziqfNBMTYL9zjSdXLh3ZEc9uwqoGzjvDMBq
LgECW/RDtyVP/ZVkaAbpj8mwxBoEn8vgDNqlmHt/ACDDtXQSt627NdwEu7bL
GlcjdAwGrfcbCBE+JeynF4Zzi/DS0Q5tBLE7XjvidtSd73V/XyjLulOA69WD
u4Wp5Fmy+2B9VtTaV+MURagobh0j+Q4VcM1n3SOYu1wXB84gPJf2agCtrWYV
ymbM2+2RCMMCxiUWOlSo5VQsyFloCbniGsmydDsRm9XC/6FEOcc35ZehXx2r
rdil97ViSdhF81rcSdTziaDxlu9UXORSBIXjJGgXZE2qjgSGCXqrmzjAZnZz
uHu9rsBQZ0EYLRwm4geDfL5ydLNDvX4HsLY0Cku99A1ObSf1pSgkyS0eNsvB
VH4Vg3bCUlhGzWKzf4WXn7xvLFGh20an9g3gs3QOPomm1siTuW4y/dzoK3is
swYhek2whNcAQTLuJVdOEyO2VxyH9hizjvlYAVh2goCxqUWmLb1obCz3pqZ+
kUGQalKTZtHG/Tl0bmJgAwgJE1wTu2H2o1n+YUkdf76bUKNyJzAYL/qxS6jU
TFIz0NXGnQMdsquvedBliTpKSRVV2OIH+flqA7361i/JQv8x5ncP6UM265UX
9SkZYmMku5IN684u+dBkyVMaqAtmppRG+ogYm7XKCOE7yd8qj89DjZQ8tU1U
cJl2INXOhbxQGG+ocLm2h5wE7OVynYFT+muxZMeYC/+fvA0qSQjP2MfNVJ49
rKigRXi5B7dN6QjCvUoAp3kAtdubP5kndwb9txy/55LSZ3mT5HOwfMST7yqr
e7R+WHf6iXirCNkk/ZOlsvKV9woT5GCsI2QkDg+GaWSu85XMhDpCxaKZ1D+C
ExRECAz9iadhTHBY/HobZD+hnxIVtCv7PsXD3ipn//HdZVBjJ6/i7UyZv3a1
PO7E2+AdK+bcW4ZeLbzZkDukp+5+gw0wvdSp/BwXeZko9N3FT/034Cp6tVj+
/cBwWBa3pyJg2aJq8SvR7u8S3bcYOPE5Xjp42bNOrx0X1oSbe9Tf2/5qv75h
B1fGk/WWIUOrBqsXcQjr3DXRAkFK37Eb8NnwXM7PCG6IqSSbNipa3gL2+Oj6
lJFjZyNzVcnpK04Glpf7DlAkIhDXsT3xzAvCTjwxqX8cqdwPyt0Qp2bAGXFb
TXxuLJN4hw4ErEpoY7Xqd9ltRILJIX5mba50iGWeFIhS/+3xpSpGJL8i0ELt
+0qNZ7M8B88/3CaEJow913IjDql4LYjgiox0zcGlGqvo6O3eWv5X3VQpvKAH
zat8jbl0mJic0C9HmJya5Mxb/ckVuTzQsUQqutcazPBE0Y+GXIK7EoXTGnY5
tj09pqChSosk+CjCqul3soGXV/35D6MoJYfyqTEmIj4BwtZeFqeF3Df0/F0j
GQPAWD1lmVyK5wr5Xv5poGfxM5EMPPw7PRfcFLRoK+KZlCUMJxJVikoSQ/+h
6OALaCT8khnmhRpli0JRgHn2h37b+uyt3qAl0SUxPePisB6AQeEgwCOVqBcO
sawUdoJ/X/rlSPNFJdpgPD/7CgVZYJLXkX9WeOybTwh6bivwQJM5saNhvVst
sj5tj/RoUr5O0zE9M0LYRiNaNmIQEH9my2+97BLoJ0JWAIYKoc2MarHDOieS
odjNu+l6RrnCP64z1xXQJYFJnSQOB59lYd8NCOEzh9DqvWmLKZh0M+wvlVGn
/GvoNNxOwdYq+P0PdhYoV12rMyPc6R5eWrVHcTuOuRtqUmVhDJUt4T13l0L3
QYD/C7haYGfrh87ALRFtN/UIGWXhOfOJ7OZj/bbDganQkf4K/q1RVtQ1gCg5
gQ4rcymZPU/VvUtUCS+AqQiVyaln+5SSphEkfBal2uYtSLOwZvWEZioFFxeA
zcv9fAf4jExV8vcd3LeWkRoX6TviZeNR2/2dlUALpvK5FConxe8+NqaspGQH
1fMtvIAE4rI787n+zQr0b0z9/7v12/QmcCg8R84R28JOVQYPd/aksvZUbY0j
bA8ZjoeFLnPmXXtQd2rUl6n/IP9DTjCOT0lWcBFc4NgCOC0rtqBNS5q2TEl+
16E3AwKvTPRzBdsH46LAVhtfQPjNBgnwDXbPdEfZ2spbAO9hWhRV4lXuZf7R
0ucbX+nJ1wUl3lxYo17WIHvNhBGxnVDFxbhzy6B35wsQWVyF9fBfn9smvmFt
wAK/MCxySPUOD4oqZdMY/bdblnywbxPYj3L1otK0BKHxeYeWaJc3f7Xp+Dcx
d1iauDPUysCK1bL+rqRpDBFtV9meXGasVzN82E8kgN0ABZLZQNxgGrwxB/8q
W32ZheJafpGd2iZmtcynYoJzNz7tbqJinZ6EB1meuPO4t1mFuf/UEQwQsrJv
qVkNfpdPBrsKNiDgpcROrCSZJTT/ItLTDUz04DtPBUT0X1qJawYNeU39cxk6
EAiyowC8Rgu+2bNY+FwMgk0ritqUIRUo7t3Loqy2yZBbQHYXngqA4N4EnwdE
50fHQrN8KN2EhXJCZ4lyF1l0XwN/6bo2ZUdVbD0xeRs6yqNKihsOKfjyfw7H
+p7t/iD7EI/yVhIk8+L79ODzqB7Z6a3sDMVpKpUEoiA2UFW3c0NZlnBD2TW8
/zWH9umNDhlL71vBavdiPFMSzZEKPzgHDEQvLvIS8sjPeLGCvXUWLKjpFydv
URTl4o9DMi4D3fMm2vE+zLrH64ftYyyyQs4jEQjMUckWY79gMKaYgbsCYn/A
NUXbD/ew7+GLvHUWAbvL+RkWdTczw2RS9tYZrHLjwijI9da+zpo8GHw31hpu
9meqkOtSyJqXO7Xz9gL6MlwXO54Rhu1cJyv9jyAzMKrxNxSS4/Rxlk2iRwiR
PCZY/FHxDu9zdYSDOntaB91/MpuK1/sBRnd50t49PQT5uueWrAS3iju2tPbI
OEU375fmOMQDNHmowMQDcNF0JaoW4ajuJ2nYLH5pVlejAqXSdimohn4Rc5+7
MU86VJ80cnqKp+joVMsc7vn01tmUUdRoDRu1ZuHyBCgnuef40qJyv1kRkZjT
axAqeGfbKIMHTMV+AWvXeCkM3Z+K68rGTP/UDJDEbgX9X9//h0ALwqZ6oO+b
19MHJ7tBRSst61kQvU2adNf3Qihu/KG26pmNYbd1/CfRUb1FsGlEHpZ7OSpG
4j7jPoeY7C6iXViNL2hJJ0aDT73qGc7/R4ItkHHH7feVgHBPlgpSoF6e/O77
cZzvDfviizTT5vUK3p2lLxV9JCgqx2FuihyMOYGGEFZ0q2Vmix9BHKSRDcOM
i/CzWZBnBPX6r33Aw9/h+FvjrVNYLJuloo5VzJOeDSljjIWFuqoWiAo9aESr
9anxGJKp1osP7PFovUxDuXUseh7AG7c4ZhkFk8nDQ0Nb5ZEeVR70+GJxhRHz
etfPUsTjQ9H5MWlBoVSh7aTT8Kjxv2dHXMs2KY+HMF6A74aVi7dMPvD8lV3E
fVds+pBnFu1TwD7zLoIzhCxGkGYK48vDsBFptD5NQzi+f4lv8tkFpm5uWPCO
6M7Eg3N/z38Gy1fUzAQsbFkM4m0laZoRkZXw8Sn4AuPvTHhPvBKnKB1b12uO
+8Iv0vFP0RZ1j7WTpzBtgH3QgCF/IxSncH5z7evzePCYoli2gwoqIcZjRmkO
1qt/LeEFkO4vGuuFEsIoUdXCLYhd52QtWtaSHa8M6V68tci5eFF/mR/1dvSU
+41QC0weXeVs28cBq7szDlKRNekrTdKkFHOGwDFWsv8+BcG14BTCGJEBwrv0
EIhBCOfWPMXcih3+OUCBCqiXbcw7UsZc0QdHaRLvTiqoahJs7wemGTXMc6A4
SGN+sTbjeBOect8NtOMhgJzZQKHN1GP0Sd6hgRdif9VkKh7HW1v7bCV2Ic7n
zu+6BFgHGP+NVRTEoz9kgNiAyq3ZdSIZRPlK6Kh7qDmLG0DUrfRHEVikEP5F
mJxky94laQdcZegR4SxE5U0EJdf9rdMCuxHn2wql9h7WZaxcbSRw0P23qUMy
heRbIsD4+JK6c41Kl/TdoRhfYf4lbGpJXB4f0MtvyIub7zafI0ZZX9RN22ks
sFWpCwh//2a/9ZEu8H02L0PnBMzX6O+vJbarZPNugAk+yVrFB3qhkjnfT83w
eHVeKVPmJoSmt+eCM7gMH3evuMOF7b6WaqiEGHZ+NOD1A6ILB7s/kNprKV+T
Qs2i9azyjFabarGi9KdAO+9igYnL1XOsN01myYPQPY8p+So5Iix/OAfbS2Fw
y36YwhVspCW+EncX3w==

`pragma protect end_protected
