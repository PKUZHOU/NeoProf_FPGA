// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
vmcoBxVQx6jk6R+MAgHeiO/COL03D2psx0Zr9hC2yOtWw8gQixpXr15gjvEoIxDt
2AEH9sPY2SrxnpZCm0e8rKcmKmRyPRXjaPF+7DKsBnFP94iYN7tsMWjrco55qyzi
Me9EBlzkh+ZXLptOpUtGQ5hfshTNkStY8026GYh3gGEYrXTYv1e/Yw==
//pragma protect end_key_block
//pragma protect digest_block
vOMYXVtE5P9u1uCLzJctQuokWGQ=
//pragma protect end_digest_block
//pragma protect data_block
bMRgvFXeq3m9B/iwcHRqGxrwfYTwv7FC19H6WL6XhX+QVJOilwwCP59I0DuUy7rL
jSdgawWexl3EymA4UlKKiZo38ar68N+1fdJx28FPRT1PYqRh3bawe4MnWJoNfUHx
uWe0/zPUa1PQF6xqaHEbey4zrUGJt3w8dmI70Rg9+Zjew2LLIt1BoN2O+TRPg8LK
WiUcRRdwcXrF3FulC11N4muCk0EtJJYiaKs22JdnLS2TmgHPWMEqnK/+qUcgVwzg
2dLtS+qoCjlXC8ir4iJZvHho57qWHDQeK2Ff6JhhOmRNoSwacIzUScsQvFbpIcB4
3wQoypCB9p8WGgqjipXIOJBeS/6NijBMEL7/ZsbQAAtFE7hhmhw8OoIC7TMItfKY
Pm0IZDOfO4FIBN+zvlH6BBonuFWxuCFT7XUTD989pBd/EwkPTZ7iCplxrbAJbuXo
ecN75Bf6NhCFOgwklyOQ9nFDtJk6TvKkXHyeTA8QeasLg3TkKbhx+zbIdU6X/oQT
bOpuIubArS3IR01jiZM22kKopxjl2kEZzLEYmy1S+Prn6l2m4hLP9oLzPvXPk4ig
kwG8EbZjE5WO6SbQiARfG3786HpMXqj9MUVPOh9wYrWyAyp7M/hWNaKOo3TG2/6Q
t+0tqlERvG6CrCWZsHuQYTxHfSPmfgGnDEHbq+cujVH5lWhEaaW/Lzd3m34pIIWZ
A6x3l1s9fgy3I4WzlSEKoLGXfHz9bL8BFL1AU9Fpt1yRYcAuJCvbNLmaSu3b7eBO
/SMXfQXmrluoStqsKmnXYzNtOLxz5sM2KfTcH/v5SPGP2ry/O+KJzW1IgMvM6+NG
W7AxEaygu/eMMzWqWHD4eAKSWNRc9qz7wWm5ess++Q+Qk3xHBRWZfw5uryp7aa9N
ocokITYHQ5ESVAfEf0pSD74M1rmBvAdYf2emWRp/6VY9wvzgmQK3UBw7oTkuWwK3
NtwBOxN2sD9LV/W68AF0cLl2YngerwCAbNogI8yAlSmhsQi7L3Uu9i2k5Ty2Wqyg
9l+rkwcJCByWrD9rjlMA2fYKIfqor5Njokk+LEU/IuVfDQv4NnL8mGgOrCpofBC8
lCFWPWuwdTS4uro3Bc/pbPI4SytKv0CTt+m1F77cywlqv048BbRKqPpr5pq18Pfv
ICO576qm3PIeNzr4MI/b8HIco3ByT1Qtl4GByQJT0lokK60Eo0YqOPiFEY8ZUlZk
97w5hOmC5Zlr2MDFpQxPHLRE1LeKZrD18k0pMqaims3LO5FXs5Vn8sIwEpUcjwKy
wUrnvatyXvHDKhKM8+gbo8lrrxz5Dnl5m4yvKc/0dqGHgHNLQd2gw3geY7unQUma
f5yagP3/JgpOSbytbi44gM2BtNCKcaUjlr7zpJHrZcWSXXUBI6jNfmXOWiqLkzga
U6YsM5EVgsVoGthav2u9cUZkHLviRTxIU7mu4f4m0cm/JulRiirOb8C0ghTi7Avk
UpyId97PCdTFqXkYFTpszltT3qcTJKSIXhq4OLRjNicv3npOCU0MxDt3WDJN5xVt
YHSdHNf6cCP/fIAMU/yFpKZw3zo/2/spy7XgnlycV0dhRuMRaZJVfZmS97NXmOAQ
55ToTGDGMrl9JzRRvOvlCI6cSAbkaxwGjC1JRlhkgLgf4wqczwu9iHU+/SsaBcp/
7ztsRLlBGHCb122Ygi+G/+kbU9h9pycoahQP2rxJZ+7rJxd9r8gWMh4QrcTGAJtM
IAUYKn5gxywmKesFOS3fozRqRmZw3HgFNSAIAnOD8/+7HcZ+S7D9osbB9T51rgIf
4VEvNrQBbbJmRp8norcsmvaMfpUPwD2kfV+m2atB+MRoGgKCBpsnHkKbZ7OAvGv2
AtLqvAp5F2fBKKOR12D09S/Ya+D5vy2G3ZWVsWbFB2SsJdc6il3to5aP0YRypMPX
mp0vtn3dqf5AS2wXqQQszfBI+7DdtNaQN75qLkxIUlTkHWIJev0BXtBa33yiDg6i
jM/LsFRlhnJGhOaDaSBgoMgXRZjnIPJppPOebGHyXndc52S9yCR18K7g4pMjq9PB
GDO8BfvlkiA80oYIQYAO9lId5P2PQu5r76Kiar6yfjY1N/irGp8CKdzWxTF8Aein
uQWxOuXz+UvInZM+uoteX6Cok1dMiiezFmUzKliyxPqfdeKVRdfxMDhvNbCXfaRv
xOVDaILrEXxITc8eos9D2hZ2QFUrsRBzs0+Va/Mn/WCG3uw9j7nZ9JGPXRqHTIao
dT0G/ss38R9hixNKZP8b5cC684Z+lHKiGHRR5wnMD3cBlY/hjxWODLZfUba6L6da
oHULFPdCO8fbW+1L+cho7auhHkOE1Zmg+A9WZ7ctr2DKuM1IbnTQD3g0l9zCsle/
tzxTF2SiMXbOQ7GfJiEhPSNE58AUyxHlFqjnaday7lJZvw7Dx2M8UmWt9dJfs+q8
XcpzLno1tG1nFAetBRx9kgjX+ZCBY8CoDleGQJbrp2N2kGLdvDn49Qh6tb9eCiWK
5Df/UKbyEZc0GA4pOjnfVtJ9Ze98tUKfRSR1mKTQO8QfbUO8QZxIyP1F057KYutq
XgQ8lSQ+94vt0Kon3lflwD1fi2T+wOzkSfjM2wDcXWny0+EYQZYQGX4Ge02LG8HM
YplG5urv8cuaPjq++OcEVMGvqlA42o8hsA+aBLZx/DeI5V0of+3mT/Kh1LVsS6t8
l3VJ5lWz0e0XWzH7hnfAzeAVX18Ep5obnaSDbqXLdIMFLsOSJr7Naxtp5Nzfwa3c
EA7gZjfnFsZLbBS9bPzw8musIwICXt+HahQA03et/ssiRNpKUZYSN86wmtjXsD43
BDstyTHb02kG08YWYMqQlqUWeI8ywrCaeYaTPkRp1Ysl7AH6QhLN1fLO+VAT1vRz
VNcNn2DTNeWYNFTTPP2j9syKyeu+AXrGd6FOMOf3baDRLb2QLiqHKuTpnbWY7Z11
vdrrNiSvhapx4gZplYngnLpBdQXKB4ObbaJhlp28cmHM0LaubSMO6DQ5wc45sok+
P4dniQoU7CLxIqUiimmFgooficDrx4529JPFuIr92DeW1tJ74Tp+7k1sskmfU6J4
vfJgl2QK9sAn+YAwITE2iEezkhrxaSoI1g+INeVgPlFGHAAdyYEHEdQ5Ypx+KU7U
gXSNq/Wk5mFQh+56CpINRiMaGyQmmdfQ5d+phRdGJlG9Whff64A97UJDe/eADUGl
bf/2N7t5LCiePyKZUwUsSYOI5qh/WSRxiZYhiw2ckslDyXMlCy11qRWq+oXgXPq+
TUMlCy5bqm0pNp/ogJSDWj1a4dT+hfzjkFDP1j6I/7RmoGMdkttC8TRkZ4q4BBqz
8vNK1weqxnckYT5+bZSODRt2EqJhUzKr97ZLup/wPOq7RykDTDjZ7isJ9Erq1x83
VFr2BiG3JSQqbR1tq/XNR8Tv383XJihs56htYgmCYQPQkH8lTUTubzDcCqBspBS2
j1QxrVQD75yWwDw8FRtKa+jrJuPYPrfg3L6F2ozekS/uJ1OfwdRE6R4ULYl2H4fx
o/9Zjteb6H6n6TPmOlDH18fGChW+Iha3bCGGHPt5CMJQ68jss8EQX4JEG9lz7rD3
bbCpPgrewtArpu00YqYW6z1mNkQiLeVZ5+n16T7W/xI28JVyxSvuM8QrPT8qYPe4
bMH5Jhr3dp8v80V1pWCs7+0uF/+zMXqx33Bo36AHUmqz1CbbISgUe6Wa9Y2vXHXS
TdWr0ufd0/J+nL6DCZYP+vkwujzhMCStazpN5hsqtfsBZS0g1u6kHQAvKWGPjdev
OV9UJmiO1rAgdCh9MB9uCGggxCcEP22aVpDH6JfoFeGu2Qx7v12Ga0/FKuOibUtD
nqtV0r1uzxuR6ztfq97v1jyDpsQXXpJNJwbqVXUba+HgOYGzefpvf4q6++/XDbJ+
Fzhqcei84c1tdvel7bEwHBZhQZ82v0KL44n11Hd5aINt0uAtAxxV1zONM1Hb9EdW
NagAfrLxngZLpXqBN1s3Cim2jGeuVxb29XIceiZJszTsnq0b91r20dr9010h4uSq
IJ969QyIqmqYx1afEYgUZaUPnlnDOJSW7wKaCV79Crko3qUq0fURseFTbb7pu5mJ
DVDkAItML0Bl8msa32DJZnDvboHeC4zMLST8+S361qx1XQm3e2yZ8Bs5m+lacWAL
7mb8bRnz5JMSNtFEnJX77UHvwjsqr0PrFxSlNIwLR2IulQiDaC90RIfKLE1WEi6/
E3RAVlAOHjc3szaAl6Ox0lpcniu+mAC9huc85hliFllM0F9fA+kg8Zx2WEzZX6TN
x3fmIERGfnbPLP39x/eIS9TV86npjytaxdkxt5zpTL0H4aem0WmPqqcaL785pMwm
KN1Kqlxy0YFv3lOEkPZwyAlfWYjFC1Fxn3oh2gT+qogwYJDANrHdogQAepDQxpG9
tAZwGNIn3B9qKzrshb7c4l+0u5YxV3y4/wf5hbRFF91gYv0bDamyiIKE78mIpx4g
UXduiroagC1xCqplwsJR2p9SD179Xg0qSTxcCFqzlPESyUZ9vhnb4RjFD2JGTCrC
ihe1yp7/FHkLCNE3DsfBzYsE06AwOSXkEgBVE273FOdpYYjFin3bFL8X+sZMpbjG
Z5tPV4u98+EustJheCzx180wyLTwhpriLxBSfbv065T6UVpKDFpQ4MweHRNDdbny
kg01FUPQUfj9zgBlp/xzGM4K7SpzMNFrZo7euQnfKVnzYL/Vn/0NushbuTlQU64s
2N5+oW/aOYl3lyAiDIeRTClKijOyYuGE4diekdLvxPz1m2Vc/1DfFsFz7ILhk51n
H2PapDRv92v2Q1ZFwAni6IXnu6RLtFxhBk6LOp9l5FEkxSKJk6lLJ1oyjyqELOMR
901a4K2cT/NYmSBHLhc3vVNXEF50HrwRdrH94pzmQk+Irfsna3b14FzdzvGKa+Lt
+Qpg78yuZdKaFETtnBEEYOkIceuGeAQNmu4lfV9ADr9EGOEymawUxOjH27Ak7hC9
9fgiG6Y6C0uxvRLNhqSJIKsT0vgcmDQsu9gbwPu4r1B0mvWn3AsuD+sFaXFlX9de
PC1G8iB2tjYGXN5/rQLAeGgnTIWZsrsr4N8mMs/tmIp5l7G1lKyn42ARFGPh1ayn
IyxEuz2Ckh5b3kAQVKpEmY2bxvzygurF+4ZxYFH3FB89ak8ANywbBDLRuonkWUxW
jQEI6fXziXKgLYznXU+QbHPJ8bocdWAavrPfA1OMDtN7+ogvu3i6ig/KKU+iFozf
KqGS7u63OWEfT0N+Geng/mtBZsx2thb4gyDx5yS8z6Cb9d73CbKnAOFmvkqH3v8D
aM6CbIYJIuebKY56u3DiYEvCdcVDTXZJ/JOxP6J+f2npySd7pqgLL0XYKHk5d7v/
CIQibCPk0aAXuchU8Lvr7FZg2Kcgfcu8reTZ7kBbHD+/RKQ8/2r8P+4U9svbOMp+
20Xex1r9EYK9z/IoVE/F84+pIL8WkZUO+3ou8dlXXmEoeAz47HoKmgqxpVMjKJLK
QaqiOCG8bzjlNyXXNPYyzLcNojoR0rOwE3CKlFw1XN4J+dnUJSUPTkvYyudTGS2I

//pragma protect end_data_block
//pragma protect digest_block
Wq/oUNLCtvG4tn1qDW3r8jirHSg=
//pragma protect end_digest_block
//pragma protect end_protected
