`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
TlbrGQK6nO83+d2pLcNY+SZr6j94LNFMq+A3ddBS0LrilJzKYHsn8tJ1kCPKirTY
Jmsar6kUPlSjhnUkV77SGLo0c3oJv95yG6xR5iEXRSVadDwpEyoq+Ps5+O3FYb2t
4i60g8wNRd4t9gkI6IdNxLTZuE4Fd3GjCWfDK56kFNw=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 31024), data_block
V/Y9YKgUDzZn8gYtirPA+5LhUV0fMiJXC9J3GLnGSii+/1RpXkeEsyH7aFJodIxN
KD0t9YlpsvIWkifdjwxCeOetQaARI1ENPintt5uic0Q9jV8aFFIbQECOaSh4PcXj
rIBHPPsX85mHgn1SUdpBeUX9Tei+05NT+gqTP1U5CmZ5/iU1ADwAXGrB/Rms9jlb
5nAO0MCEtMaANsbA+nlY54mcAgcDH1jODgxRz3DXvo2b6KxYYS5yl/CMhlW7SSwY
DrHYa4FDpsDEBJgpyqsTJQkgacDPu5+5BaEimJSTfn53tuq4dy+H/cUeNqbG6s9J
4Kk+ZCZl23YX72poP0p24crN61b7anObSoVpT8iGTekDwLfsaurFDPxRFP0g3IT8
+XboWWYX9eUSuHua6Yv6fzbTuUOOaWZNfv3+XzdBuDiHYrvzQ0fnC1cXM+T14kMa
M3s4oJe035pK/SBkVdjHJljboeoXXA7aXNRM5IJtcWQqBDFA+4XTvNUL1/JLpVkT
zsGOIl7R4ZAeE/HDciP20Z49edoilDHMyasv1HM4FPmPkPdmqTYure5Q9WJigfBW
QgNOYgU0f5MkEX7IwXpfo0q7+rldtv0T+I+FKjzfWzGyIyTh4Ljg2gwvctMWZ0So
Ms8TT0d3gkuWoJ5U3nb3mZDvT7QJi2hv9pP2A+RTKaqpqeaFQZajhWQnn1p90i+P
nOrJW/nfT2g2HJDmjB1nlQdMAo7ZTsWOKsgFbW4QLIDVLFjfQE2Z51qc06O6wMYc
C/V+l1BjtmXZahs+3lZ6PZ4TXx3y4vW7avshDZRzoiCweHbEEt8wS9SqG6yb8TlL
iM0VJgNDkDfkf7NMTppvpQaQYQkq7pvxWbYL3LF/dr/HQIsdeTeRHDGE9TG3fJao
Ak9/MYtb+l+2zBtZHwFLNXjXGqTOW/PgepFHh9R5F613CPF/7BMQDTssLxzm2JCn
zBkzWUNXH7ybpX+bxYVoQCxalzDZMvu92x9eF2rWH1TmqOiww1SRI6yTs3VEAeT8
/qGtPQyzUIvd+rnnPQDUC/RQv33G2R84LXCw0WOGCCmXQz5FaCix1VZLZPAMvs0o
1FWj9XO8gyWynHoxzUWjz/FUoCJNJAlsYiqTNESax8ADJMD99Zqt5ELHg7sf4xuh
kjd3CblLNzxOuJ+pkfphVy4OwxzFa30zHblc87S3wph9zl4jdQu5OsuwQ6P8YM+d
XYrccYI7sNklOtPxFcBcJuNjzu3Eu14RE/pf0YGXoLtMuCl/CvS7S4DrGQfFsPkv
XnNv3d+dgX9yzsqQkaoWYQe5hBukbTQ4FgHwlGc7Wi0FuL2lFzgacb+AiY1ZAkBt
xMBcudJfSZte210SxxlgU9LiCE3nAQewwrSViiGTViep9zSY/bi9l6gN3R3fxwUC
XpBt8T7SKxv2VHJ1Puy52gxCGL3ga/6ruvV9y0gPzUtquAnqlYj2BBpM6zjuP1Xx
JZ8VeShXW5aUdajIHobeMO+HgvKmG3Gr4QVWBAOevynt722D3IrCR/cn6Vv3xg55
35WVMMHG2Xu6aY/tTBqWHmJStwxelTBkol63xAw9pdtH6xAcHdx4jcpd1uBlsIVz
Hh4SxuHS/qmZuQElj9w745FziVouLsFoyJ7MMcQpffqA2VEeyl8P+aOfX+TT3igl
ugMAA1CtfTiYw40fiZ8VT1XMp6LMHoj9teH0125mH+zJK7h7DVDy4fPAh2fhCnoE
KG9aTSlFWC2DWeANkWnkJqGxaThRC/lEcV/Pd5EraZV3CBf9i8SSBZed3wHLLchg
arsQ3IzM/HBSHbzimgWLK5byKRA6KbYnqzvcuVcExvO3OclRQxhpcA7WUEJx1IUW
jPxYJD8g7oXvaKyfH6USk+mSZeJzUNcCSptJDNZFjjD2pcxvc++MmexbNUPH1mR5
Ft/hnOMd0y3SBWnwM7ZV1488qnZUBL0Y4bnQEy6iiDqGSsBNr1aRFX8elHnMd2iE
KVxhQ0A3P/aFmx3Q11+4X9OVcXX3QdPUpbTs7Hqk1sRBKEQ43It2hPRmdv9HwU4t
FnrtpU1+4K32Y4AzUb6OQcCTvxI/tRsNDBBeousaPOcUdBNik93rDyLNDiqc78EU
Csx+9Ezg6tYqommcBX+B1DXz77BC/maJv9X57epKH1dGr6M/SWp818BnQI7RZzZP
bfZMSZGJK2AXSvxrFqWHRPxNvrD6uGN8F1l7ySRaQFoTRbTZY8KuG/JYv4A7bXWO
Cj16OQ8dWzBCNZBtY1svk/BBCG+6kndS9Xeceju+ihpCo2TT81mxN1pkLn/uEYAk
hGDWmDQsudZGrgiS4yDRAAPqPX/Une50mKCWBvqTmHRzFmX2XAnkSzuwDKQyqoCo
VazpNJD26WSRdHIXB4EGAK9lwI1KABe8nvbjVJWZdJhp7hVgTwanVwyZoCN1IkgZ
klds11qgP2YdUb0ac0vDlqeP7P/woyg4Kg0b7ddWJjQ6LwIWAkX29+ELUcf5lE2E
uP2dCxpkR99ka7vh0lPQzlW7JiPXOhVeNZ6uEtCOwx3u+Nrd/plaHPslv0RzBF3f
mQ1FL3e81gJvTm6kisUbeiUoVpMPqPsGINHVZ9c/d2S8n0MSQcu5fF56iYjdGkww
mLa+Vs/Cdm+/S6uGJ1vU5ALw44HNQoQCEzUnliAvH5Z4JLEnqP2eUMg6J3dLnFhU
0FVylbBVgjIGUVRACyWNd0yovL8RmTbUsAcPKm+eeOLZE6TgneR3xDYVb5sIEZFr
vSRtENq4/sAC29e4MddxFAyq0Mkb/IBoNNADPSH5IAg7uMT8SVhJTVaogVcXKuDW
KEAgXVJIXOT6pALzFiaxCrwfWOuat3/pOVLGfYfNKByVfQoiPRhDfG68M8JVRMhD
iVLv7s0Soofn//trtuQ6pGEwydFO+Ys1m7ISet/TXyG2PPkkxLaxCheRbF/rBxUZ
zhU2N0sF+azCOxfvIDxz3NLqoQKnY0CBvYl2Ju59Pnv+4iS6JwlPnI2iMxzD5qiH
to7JaKB0zGpCgxmvJj9Gc2zjkKqw7U7pL6EtIudwjGJrwQJ/Vmtal/tQBwwsjztc
MR8Sk+5LsaM+oWaoQDLsfN2YtZEEFBGyfiZggzyw5LUz3yffojmN/haYqZB44qx0
oy6TfVoZI4lJcIBp1a0lKnvPLTla4DNsgmnaB14noKA1XdfQUA9902ilBfuIuyK9
g7V1z89mO7FtK3E/quxqqb/WI9Kc4Avb7eOsGzwpmkRhD3Ta5w3VWJ/2EgUYlNS8
bK5Mj3NmNuZJK8jfNU5n5NYNLjuOHpL+Daix+TJcaW7RzAEqQVO6nu3c/6nqFnEe
WC9Q1CRUDlDvVo2VvvZdRSzZ4oEXdTon66FltnaRJrRuX0I0bSkfyk36KwaahD9K
T6yjJZCQeS/IDRBC8YTzqsCCj2LjAQDAiGk5oqG8SqG405R4sVOuCHT9riSSDqpM
gMPi8Xw8SyoR6BqHiZ/04Q1JBV8Lq445fPA/49POSmqljeJBvwkciCST2jYlOfLv
p+hyQUrYUabd6nLQSIbco/EmTe+fKAHOw0c6FSEJMLaSWQU2+I+6j7d59ttUZkbS
aijy7NOyXFX6Va9ctTtWelvFuCVr01UXv5bf1GSs6YI4CjU79U4owEkJtAJrkV5a
MfkW2vXPTifUBeeqoqL/WhMsA/by3Vz/Nad6VbR8/F3KKkebRFJ1M+gTBNczy5u+
Br988GS6HHyKf1bCddYkzA3yBl5CtMBE3nJaj8uj/RXdI4d8gyBRoKX5jh6i8EhN
JRFXdR1G5AtokGOWUw49ozVzJO7pU+m+gQi5LbP6jU3QiwPnt3wo9aRHwV5FzUPj
3ek1ulvIrxRYO4F5tJqt6W6nk06J9iLdspJujYys3u8RAu8rm/BcI+RH3Ekw2hA+
JowjGp5ubcGzQqrm1FGOaW1uOGCL8Z0PlsJEIaQU2Tb+/a8GseCt90ZJ9RapXMAc
BiwwsiuYxoMfq5V6BbQfNIjpaHBRk2aWitakU1H4hnFaDTMaFp22n9TrpDm7fXOU
XBbwSs9QVELCPZNxbqQ3PamfbWr+qcbYMwRbTbb0v+A+och/IIB3d3mseThLE7Lk
u1R7TVWP6wUSAyXi6XJjHMrYLOwh1LX/vGzM8lms3ZbQ57tVcGbhGUvTwDTmdzd1
TGT1TQSSi3QvHl0AEi7hwGfXUqF6syUjjQdQULXBgl+4jAStocljOm5axwjSgtGF
087f/yAXoL+0PQIvqm3Usp+aQmNIVD6VZWxzsp0/R+ZMn72aWG8fYdJQm4yU6FDF
ItGKYpHgPQQd+KPWN0o4qlE4wGVo40MZs2AjIb5bBJvh3A6MzSMhvuU8qKeawvsC
O12kgnYFf6zHOb3++lcCzHVsZVwNreT8HBji4UJarPSJscnB+MPLGnVs8sEYSwDE
+XdAa+zIg/RwIePR0c2WXxvufA0YCapW+1cplncJ/WsrUZAcYcNy9K48jMroWG45
kg7fkLHyqGgHXIcEB1QlqYMtGD5U1McoQZLsbcW4sV5L2my4TgC4jsRplNWNJR9L
lTo4jKMkO0gS4Ni+Bm457lARXNoQJHTbqjXZobVoeKCUbekdGRfTqCudJKHfGwAF
oL4ZFkmg3liYfl7UCNt5j/TJQwTuMAuPA6fx27rkE5N9WptdndEaF3l882nRNX87
C66FlqBD++U47Qs4IPtHOAmLsRaHVyxjkv9to1X29GAA/gCOfRZDHYAxxMMyMtxi
mI4rViBKBK0Vei1Yzi4VrOOPkkOmTR/MDtTmzvKVwPCNq6oAgDcO57lPd+pgLaPe
LIML5hqAyR2LQSgEMY/CprcI8EBthvWMCEzXRxk3uMSVhHiOAzCY5JACYvUCnoOe
Onoyn55WpvaxXtBx5Mp7CDgeLybtV4ouy40UJ5gQ/TMLlbzusAysKV6cVJYcrEkt
hfynOf4GE6QEG/5hIgv9et4MkxjuChmdUS5qymBvUqzJZtQNmYXQorzTsTBoYq/S
reBq99Suz3iZxWlQCI3iQ7iOfuxVqFXDZ9hfFOeqoz3WvqaikRxrBY4kEpggkAcC
aSFKZdeBR4dhRoQJAhAHzKoKOjNmyZB9GQlzrfAWiDkzvt/KIoNxtbnt7Vw8+hnY
Jh4Uw/e6IlDRlkpHGu1c+J2YCDsC9Wf6yzajuPEu56a9RbUgjgEo9pwdzIwCvELm
ZFRqAF/jiSj+ggckIt9WLdXMnprbOTjimtuQYeSP19vEAgnZTPTP3fJXjAK7A5Kb
XTb4+6MoFlYWdDkvlvJ7toaJ9u9/QmJID862MpbIbq0FWBjkgfk3auvoYoASl429
WJieltihpOVshAkIMNdRiaQAN1rx9+Zg9n9S9+ytNEUvx8ufh6uPTStGejZE86KJ
tOC647Bs4TArN4VGklbpqS35mj1mmuyxBM77o5pnnlBIoKJkAVOa4Jz007rIlbHE
mkwKDJ33vpwHFR/X9JUZHInat38jmmt/nvLkjHwm0SjEj7mJKFsfzMiTdW9EA4QR
RUPdcgN531ksjGTkUgydBxD38qfFa8VrfBjmI5sDmPy2OrEbzEnIAGGvLHuy1YgK
aKIBBEy8XGbZn6Eij+4p+G73ptn+ttEnu8y9fvuGHvIFVE33qesd0rnkfM8t8ptD
q8qgMHmbOmgJ6gyq3haoS+cJncax16rD10XITJRsRijZAaGruE5/zwa4kiIz36A1
mm/zmm+SP0+pfUwBNelVUqK7ZnYZe2o86AW9QR+Xp2wiGiyRpgk+AcVugUODzbOl
UW2Pw12MdMfIjDj4mQqttbNm/xZwSZDtue2sIRCOYGgB7r+HxC40jNlmBM5LVQ8r
/dawJt6/6PytDzJUNVp9axwsKMaG4qORVwwEX9hTfIvTJPK//m9pQez4exETteWH
1/ga3TWusPVyA8cRaNsGhHUELmXZ4spUejTqeSeiLZDqJvEHcx7eeKRcH1rDJ+AF
dj+FCvfNz6XGHm4SsP5TJeCk6leSvV27/kwudObmgyYVBHS7+vsSrdA27kszBSrr
sFanE/k4XN4s2vga37cJ2mzhAE/2GAbk4ASoUjGGP8E3p37qZSiH4VRAkcdB+8I3
AmV+gI/CvorWNbn0ZcP+XPgwkL8/S6Cslf6Xqjd5Dnq3iosnEoHfpmXSmzXt3gIW
O41MjqsnFred+CegYUIKRef6rSwt+Vbf68gKznKBzxHJ79QmAR04uDguHtPa/rbb
zkjltDX59tgFif0r19t2vkGTaSsi9UeztzPMtho7zod4kKAE2oCnpRmkqmbGItnP
ybZPm6740ZbWD1q2lSYXCM90ZaF1B5IUuESQ2O1HEUYK2S9Fi9QuwtDjs+9Cj+Q7
30AJ65rjuddoJbG74RKgG4UNqimkCgeSnE8ph/QygJGk4hoU8joqivqXZT0V/2Xo
d8C6rI1zcmzvrp9r9UaPmT4olt14Sp4X/WmIdKRpjdygMIyMK6l4RbLa9hiPYQUL
nJgcq109BNlkXnyH0ZghKuN8tzivXzTqjpEmIFrPqJTYDFa2uGFiLP3qfFSkEbZi
yGRmIVe42e90i1JuS3AwY8eGt4xFectUEAU9I3qVJtA6DH+B5mLlv3BAt8NFeKar
+bD5SpZT/vhv+qWynPArFxZQr4NI/OJo+k+0Lmcd+GUKnnMWO9iTzNzt5q3uiBJ5
98qShlhbHTcYVnBCFBB00h+iaozku0WhZqWLs+yi93Y30QJslrcOmcZEfPdm+b3n
whWVIoWKBvrRAocwy9gTLZSojAZt7+Bn1tbKNkU+Gp3wA0uEUYgl7gqX+GfZEVqz
OPf9s1sfE2TgVnd5eE+joooHWIy0/P1W2ZJ7XQdmFKYEZT3Vc2L9PIkdMqKupVzm
b5JJPkENWmWpXXGkLXvrgxA2kilyQBcfCMtjlJ8q3RGYZFpsQkK2wSgkpt/YHg7d
kmuaD07liaAIJ2OGaZ1iWd0rLK0bLWzDtJqiEOP/RRevksgRHcjyeQq9vhPR16I0
khczzY+dYdjiN9aeRMYVLT4VpYmIC0DtEPOOgbscVfWhQuUuQa7UTstnVPPqy6YR
55IdmuP8vzAhQQK4NxD5dzCjFmumK6hot3BdDBryOmn2BwRFPhZzq/ewdXpM33MW
q1MnjIc92Ukwc7kDMCPgbgqOisWJlWVQ7jXf/YGrA1FpulgSxeJX5+3MdzSMXVTH
0sg/E/63sMkCCmslPiVowA1yU5bkoBXXHL+PVdbHN+/8/XCGdcUejfprrYf5W2d+
c02AjJC/Sx5ORjJDb7X117QhQxA3H77MPBCDShFalGZpxm96Ayn1aME/jRWl0DnF
OCwkMozv4+nSL4Jgt5jiTwnpgoROC+0sWSXaEitOnkObHFcaQhFi7rEbeTqhKG1T
lcrzzR0AQp5UvogtxoboomZB01e9gwKYViKJUQ4Xb6nw3AFC7YBPI4/CDLs476GA
50HWFVPFhUnpLeVurFxlkGf7Mpop/xbuNj1Lfino4Y+wD3yadM4Ctv4rOlP/nP0Y
4lE2tA8N94+pyaKshRpPReiIVH6lcN/d/xZ6jGSORppAvHLH0DYRQMtbjF7gDe63
5WA2sMYDOoMyJEmt1qazm7TxXIrJG4ueMjVVItRD2E3bnXRsP5/6gX0rNlLyfxaV
BK4AsN7Aq2txs/Hoqpi93tlfLdbHeM/GslEPK6wD4+itVwDU6oP7CpLjwO4jlJMM
HRkJQR8/aklys//aXth7JOp164v0k9Mr3nFYAWeYsIz+AeCL9Wlc42fWJMvE5xgG
yNCOeVgzNA8dl0EODZxdktQmaCDkBtY8Feasg6vOniVsa2kqPaMu2L3jFCxQklEl
1sFRX7vM/ZURe76ixm4M+fPRC3EIXOpDak/peV6IXdo88J7SppyAUD6PvT+DzG4a
WurtGQlTmH6sHgwhanSFSROd2ibQUgOxG8nB/Az5/iQhCnTeBaMGVFxPIEVCh6sG
42lv2d3BluFWmkT1h6Lk1DSSnBvoG7p15HXyM2AxifJX4tNQBxUrxcUVbHD/1bq5
6odc66Sa1TrXR2S6DC7DB1v6gZSPaWBzwPwNKvWoEXB+lwcwyHXgErqx+ZKp9f0t
WBlPEbV2QDm7X4Qy5z2MZOYoA8vJOgd3yWUtXHfgcOP2n1kJuowXXuA5K1v2CH44
HEufyV+KyTeeeokyZOqpsPIIncS3X0CtHW0Y+FHjJ5gmBv48clYx6S5XIP0DUh2u
e9TBVUfpqIlkrynTJ0wwgcqWwMt6Ohd3kzKmTeWLq2vVZNR0pk7IxZUYgJ83ebZJ
th52RypPgPND2wHsBqGLFe9JLwKPyR/izV3Q67o13z6zjBbQY8dWluxK5EbWKrVN
H+I2716pkyUPCf1nysKOoz/VaESu3KDPqUHpahWU44DbSNDiQqNOLQ8G+1J96I2B
cLzB3gdd+oeU99F02+/UT0SImi3ODdgLcfnxnUs3gaw5NTy3E//XNlci8R9UJ9gU
dLq7H6OvCXDhu1dxXZZAC7IIQpYwqi0VuRf/MxDWf6FzhM0GqQLfgFoWPPqBgO62
7nydeU7ScUWg2dFIvFr0Sp6PEgOQg4ucJepBF3rp+OPM390WN8gBveoxMV4/JqZo
xpnUoVD0UzF2byp43lZjB4cchuTVBK/44Yek7aA/pmXAIpoOaltX2zMRNYOFvcpb
kKBNo+k5NVsqMkm9s/1dDzq6/wIvIJnHPO+oD5J40cLHYr/k0bnu4qIMm1Zbl8/z
XeaEhYw/AcAP0Tm3Lf0zz+eFP/YGaHSZgGfZ8rD4Hm3ZvZdOEudoo6/9XLYSI1FW
dFyOscy6g7h1e4QM3zlSyqJ447I0GT7aDtz/ZCQ8D7anhptSRi0N++IA3IFgqpIW
NTYYFk8MTtDxF5p20nSmFx0EAFV/Wy49gls996iM1uchlmyse1Hgeofl765GGgDk
C60BjGJ6y4UXur/LbacD8NcLbD+CmMesCf2+uhxxKRmdLh9lKpdE7eOS/gahxTPH
YQ+//r7ZAksDnJ6joMmUBEHax4BVSSSAj6tuicgSctZVlB5rm47pqoMB7xQ4RrVv
6G2Mu8ktjOCmXk5gSaBiFVQTIHmAQ54U/MVbyu5sDW0bI1swGPpDaDRrkdcsWlgx
dvpRaH9hvoJvLGn5+Aq0H+jirX/dW+3h4CzvvbfAihu5bOfS78d01tO3gJBssGm1
m1KwsEEAQ1NsAaDDAheJ3jwPo4zlHgXlDznlqS5Qbfu0OB0q9DkJsPO8PIdqekc8
5cqKI9yu3KrI7fepc1mdQb9jujJ18HDIWtuxzbPStWFCxiazJA4Mb+nvZq8nIxif
DSNB5ZBJ3N1/bbOrG0ixx7lcmOdFFPbWBXxKtJnaTxWs6bW5zc1qYx5+ZHyuZoSv
yKq5AFG2+447aBGSgT+AdAnyIL91DnrcIs2/IgsQT94vDgiQdiHkt0cdUWAbfg/k
xsmz6di0LeEhlqgSpREOX0Cg9BKbA9X4+6J6U8NNNjJajKyd3YJ+viEXb5VCHqru
rR3h5+Uhk3/YQprE+UijrjC7v1DC5YDiswrRgHgdC5Qp5oYRXNUcxEFUUfxoCiIJ
EdlDjcu07y4IISBRU7zax5eXN0J0EqSL+dI8jPNWb1VTjV0xadwq8GIwVqSAh/ki
cA+2MDw6nrzMI4E0O71jcfvIDZlBvAPw6XCDaaK3XN+nDwmci//+V9VyZU4irR2d
RysHkcPFc0DrKPW1s5+IZn4tJ6LUyEHDuyr53G7RX/4WgUr+SdZS3ECncB7woGvp
DXGMIUoe3cIHCubEW0+TGwn2Jm3exE63xZp1PYMqrEX0PuUNdwUL7iLhgMODIImp
ouny0CxyLXiFPZ8wB9wkkukiEWFmaiX27g5pjPEmUlYc1jvRkSouKhoQ7wWR4bwQ
qwPli8QIdots425NWzyhBs74XwHsgjiQTm7V2jmUzzHzmFM1V9mPQ3c25Ma01dGP
tXnpT1VdtSIoO7Kzr7mUiWpy3nDxuWTOrWQNjNU3YKLVAXNxtdPscpUF8tAC2Eu2
YnSlWQeJXJrAu9oZ+tOi/5mps8Ih7wqY7nAwA4o0aAm1IHZfc8PUF/M5kQGfeMn+
S8sfGYv55JSIJvNUZ4QW6AugZiRm/tKXlJQgqgfAQMYIgG6OBS1RAgE5LnT3eYCB
yt1/Pu+kcuF2nn3xKEY87cU+gbnp5DMw+ydSvaMevb82AsXomi9l6tpf1yo2XkPB
q7ag4THUwXWcQOPUOs4OL85603FTjtLBaYIV29Il/FZhFCeJmm/mD0h5hUqoJA88
kK07H1ibXHOh1pXfdyBK6yxPNHUxyQt+0h2iGDbobFgE7YmL3i2XXNVW+iXoqXPH
cVKsq4hnZQV/Ik2kTmUdD3HJ0Rm+8lUWeBFem+jjw6gIvQp5C+h0GfcpyN4Wg7DQ
ju8XbIt4sOCTJ/9dYQCZ1ONIo8PaJ0gXp8HBC6idxtv1Pkt3ncSbviw4NDkTJZqG
QFXhhKGnDZdp6AW8B+zUT55hnrZb4iX/OIF4ZN6llTw3UTT1fUbHLNK9i8jY348F
UvnTK3CUZqYQzJbF+UPSLztLustwDSTLcJBjkH6887RlwYf0VNTBLDoP+XmD+DpX
gmtTRSQDflH16CnolddJ5kdkTEBsLTyrquK7ECEYi/v60NVKIEZRzJv/A7xD7PR8
E7vUG+eIA/qC14hv5SwKwcLDGbIE4tjXg7SW2BeMdZkmb503KGGntgmuKoQUsuhw
rCDrmcjHMk/k84v82Vpy8yhgqRU+L/7qrd8Zofipvk8lmjxiJrJu4TlmjxU/SoKv
lD5wjES0JZsHHVcVaYkyDqnXIkfpqDgGE/Ax/ofkEUqhwTOQ69mWNNeMJeoJeDum
TxQZ4Qt2NeWb2/aKUKKmToc/PCChqqTbWPd+mNyaBxn0TrDaT2rrrksLW2Wje8iL
a5BiJ8FOiw+O/9RH44nsARG77dbq8qRYDz1vD21gTVXssWbleaktnz99Awz72yqS
ta6HKcAuoCRI7416mqlljhWhq8u/rA3MKnKabdSYgDxQdOxxPTJhT9nu8w5yQK0K
s8hdPRXtKB9vrGU5ZAiF1z9boulqZ56JsRqoKkJw+hbuTtOqazWHWnEpRmMq5wEm
MTupmTUD8N+G566uGWlD1S1niLFd9+/bRvX16sBa4IYuHwNKo+LIQPrFtJxQoxWD
OnC94fv8tDHQKqLOQSu0Uv/3ys9cmnXqiNd+ku7DfmfsfdgTIAJ0pmwX3mAzF6zt
vwoLppRDJwOGzHPcx+5iIf+3lbIf0iguJ2EYsq84Y/9nU2yGAC0DKHJioblbIPbQ
2MLQoEE/r93kq9DznbFkpf7YA0HqVf6/xIOcxt+eeAe8LfKaJ8bHxiR5ky3PI/A/
X0Y7RTNgjkTgA1waHLHRO+jCmecIl60V3KU90r2pptrDOUGNHH/D+yFk6cRDJjGx
URYmeEJlpOzTQx/UXNtVSCatHsTExR7nIdyb2oXODxx9JZoqIpoqQZVcYIS9bSU/
wva/kOXKAuwudmjcHwhUmz9k/gKPUuVJXkHOAI+dONwR1T8++cF2m7PipfA6SB5N
IpjN08Wr+veI40FJsKJEqqZ30NDrELqH2i2mJOu3y10yALSDkSe5WvakBwXGz4hs
xJfhncqgzmKcMLWHNNIuTC7oeOlZxVQOgiEssq8+k/GPa/8an6VoXb6Lkamm6u6X
LwPk1VAI+ihJozPGpqodVcu7tDNfCZNoudq1L0KFDVzR16ov/Z4Jb3boiIY2aSCd
CA8S0Op4k7RP66r03dTI9AfCsqs8nnMoJVtTwQ9vN9LPfZku+vt5SuLWwPk5Kn2m
/j+y82yWnBFXjYhWP13pzrPkd157gVDnR1RwQ9Rrd2hU6mhOOlKAIIEqDUBn5zqe
5t0MlcTHfr03LilVaVvBK3ZwBNbYbaZ1iuyhGCMspsk9U/OFNyCexm+uJu93+FEo
blB+QZPYtUyJRoTXp5h/6mGo0Y/NaJf1dbz5l+2ulMMfC98sqLvSv+MfRNgswhi3
lQbhU7nX67bew+8V9anGvO6hq7/WDQufUTMtvUYfDq/iPGcZMGduwoPl/csG7SvT
0ESEjHCN/hyx0/pE2BkZg+7PcwfdSAlYY1tVdwTHDS44xtWl3oxo3TpE1mOgiZxx
dDu6amGaq+Wlx1QD/0IOuLFqORnVi+EzEn8kVlvKDF5LclyTfAMcE+JQLPNlNU8y
UDRPgWUwDSjGByIiouioZKD7LBTb/xqt1S5r92Om/zaZjMzKJ6RToOQrW14VCrWZ
6EaJqBVd2ZK/FZiQ6kVPrPYeNkmh/4Pre8wWel46gcSPg5PiY0OOSapta4GVtG7/
mNET4ztuEKDi8i+tuFJuKZhiIiUFSpulzIeKSnduBNpiAQCNX1NyuNfkSW9/gyun
b8LTIh5BkiVIIVJCbBcKWryjt5xamEmofT2/dy97u4wRT4vvWN2EevctWQdnRz/P
y5faqgKEizoCKamP/HjTIl7EIuHi/9MiXXb+KWhQRYEmy5cXmxtDIROEY0u9jYbM
expkqh/sDwZzfUCpsJmweclbiHnGsHCUlHpAdINYFaVEbO5m2fdlohp98TpCZKqi
KAPNSjlo8xeJIVBdz57OHK7Alazs+4fj9gyeU6RxurmYCSdzw7tsq80oosYlyS+f
DZHLH0VY4bFGdULE5VkMnwpi/vsG1Q68+Wzv2gRk6GSPGyS0D4kZCsFRjzfkP3la
G+0KA8fw1DaAaNJBYExXZBixF8bm2KPufvP1cGLJMcbzNNb7nHBc6VhDNg606cGJ
CHDD3mD+J8ncnAzWAU8nANqSD8Ll7aalOfClEQA8e3EALy4RwX19XI5Yx8a6MRSB
/9Hkn6NA8NhGJ/jNebv63Ap5faWy5oCCA/Jt44QSjD/WoTuh8AtubBMObn1OX897
+0oEOp8e0dojS+jkUyi4kywCVAjjzj6Ma73kvQUtL84kXg1fdOrocAztinu20+fV
S3AdIZ/5OcziVb/VVOmWBiR8LX9RC6YnQZ/ZhoeFYeXq4rICKzP4LUoUBlq+kTyZ
6wqVdgQOrcUsbjSWe45gMNtP0aEPNbK3CN303ugJ5OFqMs/jPfwGexZwGNYWW8uI
R9O/VcpzoCYsui4hmu5s+biySkblu5E75cQ/jSXGNjUBiw5UGyVUlww50/PBRCXd
Pqj3q/iJTEAfZwpUpC9/BS+hXQrqTK8vLL4uVsK36kaZexRGMB0nXgKecYkdpHP9
dK9qjQpCvpw9wXBhQJEe6KVOXzkJIW0oBHF5bCPZGB9UDDo8bPRyPgMGj9JUShSI
BQ5IaMsBZtPH4KXzopIpKsa0/EwUCzduKzpKD5ogc80aYpdjEeDRMgkLo+VZW+aD
ZoIa3NWruoDl/ZIGWbJTWww+K8w3fV25om2UXITtLvDwWFhfXlOdZW7oKhZSSZqf
TzOuer28ltI1tzqm26jW8YaS1EXRg4OnAfztlY1PJ73dieG5Y0OJhsN0lWNqvrHb
LddMvHh+2GA91JxvVXT51Au5dq0Aq0669/mIqxAoTLQyr9RAH51JQESjxW/wKWwk
hWZphPxikTEP89no5JInEMMuA0FJWOjMzGkMrcU79rd921XauF9hyHu+5zIkfPfw
+zzd+GGkmxLQkjbryp+tEXZ5dwvbs1tSVtqxQuFHdK+Iwv02MK86eX3mYGN8/WQa
JRIeR3vVPSVrkOtU7X23ZuB6+OwE5R8UriSQ55qmIPwnbQn74ytydow1WIiXEdJD
wPeRB1m807FYuQH3I9VfaAvbQM/jDhzgl4exW/DU1KFJFI6io5OpnNyTgSqgO9W8
4UAZjxxVSK8t64tfOk4YNQe38gmb9GJ27FXV1MH2K1woXJKbENTP5eyKhsxMsKY4
o+etMta7/0+3QfVhFCJJBcAtlFHKHxk+F2aAGuwTOtFFYCyBKtZlouxs83PVEGc0
Z9aj1dTUj/TA1dlrn7qRFJSkNKw9zAiTuhTxFDUnQkXjxHbaompLdd2DTpXVKji5
8rUfiaID0RQwYvyOfyrf9E13JbGqAwCJEzHewTZ4Y8pxDMnlewbykrvI5g9O8Luw
SBvs04P74KsaVtKTJqgKvIbTu/UpMg+HyqOt7B8s0AXNmz3m6YvBkuASVFixVNG4
M/RDavmLOAVVHZjVQqNEgLdzQ9xv8z0YVOt3phewJSHg5B/gmHXuxX4zlBjow/1N
NscI5kDIMrPOfFNt2MciPK/kKOnBUfnij4SIbxLz5DAs4AGeAnVMYDYZXmbWyv9a
qDII0CBQvAGQzVYk52oS+7t4pyO43wJAugwNAGhXfdRrZAuzDjW3qi2cnlgOHlpD
XavtjDhU018X/j2gZ4aLdL6F4NBIpS7fHsdS4rzMVQiTmvx/sRPL6fVmwloE0eSE
XEbo9M69m4fgtvoB0FqgxREgRA6/M/lZI/rTcn8A00sSKcgLb/dldAn6QMVNliyp
JqCWQoWeWqz9ZKRBWEkr00q6lQsokpoVyHaU0rxwMKjKXScwpuRWRe5JyXa2WQgL
mT8GjbvD965oSRFCHg8H9bsfKYpGNu7EhDnQ99aEk7zaG62BVrVNFyylb0F7yxyf
v8Qwd1tLXJQLXcMIecDhAS0gDzBIdqlAu5BS3leEuKJxbtTgrT6zHslf5hOkwqC3
YJd27TGmVr1hz8n4vTywVPoAS3qSMAsnilJvoxsRne0gkr3O3uVT5yjZIzHcAmMc
kfTVq3wFNvZrERgKs9wZaLRxu2kipTyIOoSkd4Yz4J7dtxr+JwG7GpiclZXRpjUp
mbcrzkNTgCpGGjQW0IlCUI5t33j3PUKn1rtwA5D2il7SVojSDtCXrAtX4+KpA8pC
qrhUIhwCN1LGSk6gzoBY5vWBwfd3BtngApMSmqNj4eTcCDAwvN5PZa/lB59lMmy8
dW+Ca/tS8hnwgDwX4OWGN8MkLBnjP7dHFGqI3lsHSniDqH/UEs0Iwkvf60AMLlxi
lARdMfOsheW/z8VJu++mTLZJBSbygo0AdLTJfkzobFHE8IFer4BHqDSBYFQ43ggS
rUs6GTsN5O6n4GJbOPfsp+Opf+d9Rnp/6WLH3MWOXiIS2Buwr7zKr+tsodeYcyqc
8dJwUScYHoHfMzgV779Nmr9Vl691SeLRzLz9aqxv8lwxaSU2ES5TV56csdM9Iljd
ov53IZdaXA1AgLrmiVGJqmrubP8sclhzMLxeh4mAehlZqK4V3LRKCwDnRQ5KnCFe
bMyMq7C7ZwhuIoOO/Y1bD8Kcq26L3VEcxYJGwJ0i21dPYm2KYNJw3z9sjkkvHMUA
gLVXv+8YPqUpMYqkUJ+RZZowe7b2gshqFx6SJsHh/DaVAo6Z2LRxPk6SKV3MXxgj
7P0OZkmCfGgV06jFfADl0J8IWjGxSbKZR3nnIRM/HTrQy4X8xqm4qRf32do+GgGH
aOZVI8uIhxkVNa7qBKIKBQWCHhGvPvlZhwR0LRtRfHRj4NgGLbDUd1Tb+IClw40z
w2LbW6CfFa7eMCtjJqX5bPGzcRHa0arJKTyj30aBdn3RF1nUSydUN7D42TaRH9XC
aYLsCO+cdsPtXf1ZqT6FlHCXJyh33qev2Ffu1W9sMm3OMuSS82bB9fERqpT0HfpI
tKjZPEF48T4YAyR77t3xbjCz5e7n6QXt342Poeh1BxEMPlX4EskRvr42ok8x2cTd
r+2vx4/Bk3zjK4wEyZ5mGmUjxZD21s/B6Mf3RA6I3GjgTsXCVzgpPOxtkG0lwxU5
AnS3Sj9z2ZH3Q5ZeQz67pKnW2NRrqkPh/LsKIaIK6eEK+rVU0LlMtycLqrKUwmNF
0p4ze2AFpBAc6ppDfC6jFZK4N7jg4d9t8i4gGleSNJdFKL7pNZiJBcakonm3dQmj
f1VqJ6SXdMVe7w7UF2HgznlRIVmU86ArSDbcoDIvkTGTm/ikyiudGhK9dpgRES2f
bgvhPHMDK08JhgwQtCNf/rbN7hB8pPoNqjn7N83+PsvnxZImf9U8eysM5jjQAwZN
IzqJXyXwH+u9A3sfd2TLYntef5ppaJXKKfsVKPS7A4A5UmnJyiHxTXDMKbzaFYZP
5oqsfR6ZX5K+2MN4S0vTc3sFmIosUlNiRFg1DQ3PS6CnVf/1Hp/tdrrA4PWuhk8k
DBsi2k0WUwGHdLdD/Vc4Yj8Xfrcr14PotroPTgR1cyqW5BB74xlAKiexhSW2k70X
bVcIe74zInYuWQlQsfx1ODJxqasep1GwX4mqe6ONhkaQgt9DiWFAUdkxFjVwhnWq
8D89j/yj+CdhTQ7sijXGqmoxY4aTPtJX99oSTncjzqfii6vK1GjOCy79F+hUED7f
Ia0STOu9WRYfTcYSj0Yj2CIgjZgDXFXhSeO6HhY/qKaWLdFmZzI7kAY3E0Qzy9Ug
+Wpup2UhVRok9IhqctpB75saFienfD0suU8roXRhGr5uoVAIyWNbCvcjmMU1Narn
ywtov81zvEOZxX7G3P/JuF/FnfVDkM9m/WYST3RCXX6Bxlx3UhiPWWzUwjOkMVbv
DcNKHQvWUgDCDTdpKhGEh6QCYXjmW7wtq1BcTPAi0klf+m74fX0NwD5ykelrmZon
ZqEHtSwwR+aaHcmtAJR6mIYlV2JmiPOgas6ivFuzijDMu+0+tfVlvh/ULfFjnG5k
XMMZFAVZjZ0Xla2mih9HnQOC4OjqkA+eIYuB+gA1j8DbOLe+HbydIdLiBXYRcRnY
3U4eQjZYrTtklzqRK9QtpGAOlTx7JzNVrTZnpIne6iwSCHmOOhUBwV3I7Vs8AHnb
/2eXzzfLKInzRnLNKIruE+aHvTQc+tnqXvbxqPtrk5FcxIwCJgKxaY52J/GrMSX4
wLPu9qYAa9XfhW/AwwAFVwBiIi4ZvHO03cI3exkHxHWMsX92QQTwuf78XlNWWfaS
kw9FpjQN+zQphUFSN/19Hza6vJ5GBaJ0uIRkyt5oILbl7AnIVVzbcVa/HQnvHa4d
AVI5ks44mLrSkKuXOvKLBw4x6Ft1kxR91KHEhGfw/oZbUOjdkPpfl+smjTQ1HQca
XulzVyFN0ayKafEiWm+SgnW5e909uqkqePkXUouwuVD3MhvNOx2YCdvPU5gKk6vc
tgUP7PpX2QicVnQdZpDD37h2cPeycgHs02fTZ72ZgrYpcwDVxH2meJlsbHRdA4O0
QiGwM9w90PZmPLmVZay4ttVw75CXwX9JhG7CWhpwtvNWEkFG+QivYy4zkJi+Rsnj
g/0jniCDyC9yoVqPuDvdvNQqmUAy4UmpqnzTFsAhrdvAw2Of123WXFD46wQ1z8D7
RwuwKv7KuSD078xXqSvaEUC5gyQhtdKxH3ju26O4PvUtLgzn3iIUfo75yodBGzCp
UHTf7YDDKTiEtJEa28f/COscIzpa0jlnZZDKFIr4PBDaVdnKWnw5O58N+P+Ww3Ku
E4hCkh+Vo/q3n5syBHkig+6QsDhJmiuwxyw7woCLWAJUgWRvYFgbVQW4Qmes8NM4
YMtliDPLYnK4cevc8PlmvcJzu82bTc+1SG6gjmFPhjJIutJOn7uo6MnG+Vr/3FIg
A+KSIwd4oZkOHYULOmD1l7Q2eUAo7OK1RmX53yX7gLgrETFF43x+5cD5XCmvA+jp
iBiC2kR1EtSwoAi3nUbfefjc4C2v31DQRU3cSC0VtLYDBYRT1LV3StDtnZHUh8E/
ZK2XFcG8bx10lAbMTXR/oO6P4TOGyWhouzJ1zybzk6IRRtchaiFuzPgs248pFQoC
Cep02Hgk3dWA90OZZuI5B0WzQJHDwRbr1HMgw1JilIH2ju70tJFBoWMPr90kFK0C
UVeNPCa9y4pDV+Io2gyRFV3NwS9TUAKRIg7ST+zp4ztAAQPHjBEDsT6+aOL8XwNi
h28H8yJGYwM65qz3vf9i/drXZXZDLAcQiFFCr8hIFnpzUenOsCw9/7pRNPbdQtCt
ALfrqate147JkW1dCjW3XlOAQLhp0UnPNQX9R8/WYzlsb2bJvut/Wx2CnfZXFs62
7vb18HazJIxtkkBfa2IoZJ9W9kkImqZLhqDh5UvePaQeVmKpT2kbpTDYrlfsSW4Z
BgqWd521wBn2JjfRh0TcXIQBG27z3qdzf0SNCuXN4aPX6GfNi5J5zVEjntGt/R/m
bkSPf3NvxrGxYCvV0u9xRwnEa1LosDySJtvozYbgelos5EV0FRyHFU3mU/vKNgDo
XhQQALbZJtRD+hW5VhahNfwFl9O63IE1V4duPlkjMLftEGu+EZB1bNd2sk8KvTYA
o4TTAQsBaN0pB8VM/b3M2QfD/yUkj4qBq8R/LpE6CsLOPtZZ4Ml+tW8FG13cBvi1
RHRyx68M08OhvempLytlHdES6uuGTKxWFikwUNdsUtxk/Aga5rHrxRu1IhRhsn23
QZ03N4UgALUC66oyf5pPCnEr5qVLg64uRTOHifZdOe6aWkRVwdAiKJvUbSjIBqhZ
fS2DZvyyiEnomP4M4uqJdr4o+WV7hBju/UrTEGILc3ajGUJ1D3cfS8IuMxPFnRtD
VTiHdws+lXyacfwObc/1yDBbhdgdMXUPwFF6PYHbICFK5CrOrL1NVrMCyzohHgAp
zgBvIZNXTYmUmUgoc9bO6TOBaQo/XYFNA1MzJ4TmnYDTNbn3r5u5SwiZCWWZYywk
JQrrtWtcoLFnjWVU9OAofq8xF4boeXVjougYuMkj4lhNjFn97g/1A/06vaZqkNEa
8O9Xm6xvq4V5kFOC84A0XgW6V+AXfDyC6lu35dFfE81Eu6YgUB43mipDd+M/Z9K+
E0xF8xCnDsIOBz/WRpa5ZUtfBDhvjPJhY4F8gt2ZyHS4VGIbakxM2jHrOOYLy2TR
Gw76CXocGwZ6lxxR4YXeoEj+w9ZWU4Ia5QquhR5opSxHDIFBpVPgQ2ns6Lu8cRuU
lNWyBGICOnzGX32GLU3mF4sOBjC0lfStJACUI/BZ19tN1xgqNzMrSFOBXZphFjvE
rtCc350bGTGRgFqjff3dQa1fJu6E4rosZ/JwESRlnuOjCTbd/N+E6dxlB0XyWZwp
7OCoLKLOXc7ir7Q58JBe4W5LTjpDFSJR+92UsfbltCn3KsznYN3X5KhQqj1JS8mv
QnRiN/aQUdoc86KjxJOVRv13hfhGMc2RcftkuJ0UkFXtKXEBXloyDMqJWeESo/Ab
0J69SQpaOzhzlIVoGVf/VxIHt4IAn2kFY5aGTd1DDoIetuxsRAKCUA+76IlhqjdR
UOLQHQz/aPBDNvRR4pf+DTi1bdkC4T8Okgszf1M2+LMoy4zSvZq+pxXf/4IgFioe
qBF2WY4uuWlRlPXGiLJ1Zby+InJzBzwFgSOpjf2cLUrHOSqHEBOsC3YTYObQUm0V
EeeQ08tyzrGbVjznEIT2KLmAf+1+2+adg6nBlprSfNrBcW/hBFiLFcpwxxK0ZIF6
mSoKTtVwHFwEz99ywN8xSrl3Xdb2XZcY7fIikeeG+cBDKLXQcE7PCeCYDzGLDe9W
ItXJ2OUFdXG/S5E9++CnYmfMUb2RvxGOQVzNI9OHVtpHf9pKNU5yHOZ5DVINgOcp
R8cAXWeQjiBe3h0czaLTM1PlO8lf+1K8CZDks9h6H02dzNEsnqHGgVBIdmFIrZri
V+VhI6kpoL9u4GIMdHclii7KiH1uCM736d6hKRle8uKZJr7aVCZhpeV5aVqwoATJ
1vrNYihasoHEiLaujayloXdtzn8HtCUoWN2F6rolosQ/KKWltaoqPfM5zB6c7klq
kTb7rNLiceYFeWQ9YK9+ibxlpnWeOmi9n9hIJomXp525+7T85sHwozEh/mHC84AK
R/K8f1+CtO5Rrek2DyatcDBSBGaajbcjsSVXe2f3Lt4hAcatK2O+BedVTvL2/kb4
NociM37fMOcyihMFZqHVcT4pM/sChxDo0cD7C6lDRnRb3YQ1ZJxb3wM/sV20/AzC
mKiU/+QC+EYvAdmnP0r7FTOtKs5oM8yZrC5lofJ871nHVcKwQnGACQtBb479RCi1
7opQAnPeuADQqO0obx1zWuJMyNxkJ7QjPkNQIaOZCbO+xJ8wQX5J48717RM/4vyy
jryyA62pfPUDMO1QvPbAmGL6x696Jo6T1BCfNWN8AK4o7aXncbS7hJwHJ84AyFGf
20YEqJuJONd+vfJS21XS6m6GpJp4tAlUOSGLo0jO3S++LiU2v8WT1OcYUD4RJJAY
hswODkwxKOIwZRbC1rHhrtUSf6l8+w5fW+ljSMSh2DAFyajHsJRLTsnilGjF17Zb
ihHVtf+kRl6WdzbxoPlfZggpB+nFsYc0cIVG0e0T8MhGS3xAXeUB2qfR2muXJ7fB
wxeL8HJ+7zQQF6nCnjQ2VxdtYsDaK4nTpvh7spP4uM7KT/K5d8b6KftmOAUkMxHb
WUfOdRxV6NaifJ/eArbQdl1nJLbF/Lf5Ip6rTzQt+x3tsVD2vVhkYG8yaPCBVi9D
ZeQMOzt5YxvuPfk4Bq6GypMRXxMzungoKjmUTmFjqkPGqUKw/HrJp8MdjsYS4rz+
kk1en861vvh33dEakzONzUgEhY3PZDq0ip5yQqxHHyEBrBk7IOomQU5ZbYlxGOuf
0y+ZMFvt8jdzCxsXG+g2GakzzFrAoh0A9Ve20puYkB+fgqwsuBM14z3P66i3JkJN
K0wN8S4wV1OYOlatqUI7Ul6Vzbjmcy05+cAIMZR1Z5wsmwavDlagIyaFxOlmJOhS
8xYy2NrWlh+2E3jgT16BxiHntXszoxelrUzprgLSSW589Ex0Jc7Qkmw87ROhWg5r
SfvKKzSaR/CsuwEKyMRgyln/bzjWz+JogUSn1eHM2oxj7gQp5SzhfKSw+9c7rEfe
5UGjOuExvEKSodwU4LhZNpFnPcLW59DKDM6ud56MySSGSqYRAbP3dF/tEmIvNvxv
i+ydgArIMHrEEAc5gsS+wsOJWEqPHpdRaW3J67JBuAcNDDedS6n3NfsHvLy38a7W
0audob4Em7rgtENKaBMCZfCuBt2JGcSB0InJpRp9bwh8I+pP2kaw0BHnLXaRLozr
f2KvLNKIZHymSnuNoGXadGx68O9AEWQmDzI0U1QI4KsQDbZNY/y3YjZiKqm+Guid
2Kk5ZDY0muS+J8tbqeO97ErjF12RkbQsP4RUtSiYpR5g4dfSTrxl+E3bvHuaKxyD
qEfdO26AUKRMFf2OABretJvpcg086Fn+ynoa9LQ3AGuTRPAY9DamDdEuacm47UXf
0ghTA1LP810Y9pFR1vEWfKhH71wPTlxk4ndGRiq9YAKrd3L8SQhj52maiwS9TQkS
VuQu6fUxDtWq5VtkI3JmNN6Mtao9BFdJhI6/u9+rnTcmq7vZ/cAKWA9SfYOkqTdZ
0AEMFYHhSAGP5KkQBxWjVCyaDtdW7yF6s/8maqAAgdL2oRoZ0LiteTOfwPNOFHCO
/7kew5Mr/kpYDQjWEBaopt18xWgqqp9aYUthsRHzL3VJdqzKpW0ujKDzhT+GBMix
vCsEpm16DdUmDhbmISZlAz9JbkQMRFegqEWd31aoRHiBqSUaPKKKpnRSKzkbZ9Uz
zIiBnlMICrt2/TJt0V2dWA0zzPgF13dKh2bdhlh5j//S8ro66l3+o5kuPOxI4xKE
oXIX7NnZhNWBU1QXgtj5Gs8HeISinqj5O2frPQghZrWrOTPtgGK1sKD3STmQL8qW
n4o7Y8elSNO9DKeNuW4mQUHQYMUbi43A2KvVsrL8lrLQUH9Hx+8WBFrq+lACKzBY
yu3RMsKMP6VhbVMUbhhkOiAWJLXIFvMN3Ccmjxvsf5ExcZ4sehWLDuSbr+YrNR2R
kiCb79xZXyILADm1CgEY9I8coDHz0t5anjiKFIXsxncYY9elQECvbOpVwmT2Rnhn
QEU7clu0NgK9QQAiyXebm40nqtoW8vBwYKzn5bJjyX8H3vycHpdx5/Wc2Lus0Zfd
YKbYEAd8J6VGWxWkjXQoH6YIBgV13oKZKxXkKxTutnx9tZJlMcEQMP/65J92MRX3
L6EkPgcbdNLB8TfKvs3j0GP9EW0Pivp2blDpmSoh0AL+VKQL8RP70uzbCj0W2Roz
G8CsCMtpoGvtxbAL6220Ty5twlFnDHxUC1+yn8gdc+64GV34aUEWs1ziDciVdLOc
EVEI6e6RIV6nQDqajSIbgi8c4QP++CnsHyC+K0ojfhLlJCWHUEMlzq3jfSLxcR+7
MuRDDdQ/OwN+ixFYjTaI5p6AxEJ7gXAuIlUCGVevL4HSa5lcHpb0pruC/cP/HZ51
mN67p0d4otCUiUVThg9YTmAXTi9G7JJO/VPrHOxorXjYdcmsP5BAGmkzElOYmtkC
qxGDAK5Pm5eMPpH9SKaWc7NXsws4BmeVRIs6d+a+vfs85mbMZGMzS3NuN8pNTdAl
IGPJ1cUyX6ZmZzdH4UMFxNw41p29c8M5xMLNogNFnwiYc5OKPunMTuZ8Tq3z+6l1
D+MWeiQZn+N+dTiQYllqqq2rcTyEpiJmw+RTdzO81iB/t2z0L1eh+but6P4cd7YJ
cvPIUDd2bVFsH+zDWAETxmdasBvmCqHodwRT4HhujMM68JE3CxKe3J3fMmH6NoX3
DL2m6Gh4Wks4xKQbpfu2dbxCh0pVd139gk5ZwL/pEqVYwmw7hfFWPPSTlevZuiJD
FjnvMd6dQ+2SdjlE4QK4agW169FpUkyDGyVNCkx8PALFrcGJDNcyBxBbY+G5HeB3
YYE8OIav2zX43os4ii1pSySwQz6i9AO737aupEf2PF9/hnTRxpBUd8jUWPmUdIj9
Kes0ossi4i3lPr/toYVx9mHFOgBfTGneSGN/tlfoXFWDHFc1pdC1JI75RAAtjSuM
N0hYk6lT9pc63xv+brl5EOkA4FLMvpqzh52fEolhKWKUVxm28SoZuyG7IrPu3NNu
+JIxRGLndN0QnLIVN47b39qLdVwXu0+4aPqt+JfsXAJtvp0JYX18rxRLjKVQvuKh
765Q4exStK6m7Uer8hGXJopchV23vWuWjlLyZQv+ud0UA6shNmNEWlay2MJYbOJg
VlMaI/kfZ3s12NtHfU/vVkjDaRG3jTRBKUmpXMkEOOPj+vspU2olcjUKbmF55eKa
qCEqW7JHPm/egnXfSSWJLBCFmjfYpRdlamH/q0ezlBXvgt8UPtp433O3kozxZCIH
1qokuHM3ERRXXaRBuGRXXbcVzfmaUEyNLnhinGWYFmzdxKCya6V/k3FrsLo7v3fc
wMuJMiGLIxVrGY5KmW49t2cqyzOAIaa5HjzNYrFV62C+v0/XKLaNvZ+4kq4udjVN
yILF6n0QcwRezWLl6/A68O1zDwd82vd/ZJjSmUHto7w78AFaGiu5r5qkf0RUiqqY
pb6SlcpJJVBiQz8EAcbupE7RP9D1cpk2dNK9jVYU3eg7PDUVVaS4rfNARKkOzq+V
yq5NE/MgjNFzfRbGfzJsojcUvbJEo88Yhe4A/onKgb7DFvLHKrThkYstnldt2yPj
y+XbkfUynteyWpZ9pplVeWo+zsLT3MOaCiYg4t+xctl5QnOX0iLSL+d74NJQiQ/k
9n4Q5XjeOVD2z9ujQ+wrgx9BIlRWkJTonm6bYfl8SU/RPBqr+OkSk1A+XxmS0Svn
erjC7Hss6JoY4jp8d5Y78UjUxv+WwRGKJKjsydCgx9zhHhKYlAvSS9JZUIs9LK1L
0UNhjZ+dhIA3XrQ7eUQGyAh5wFHb4JtMWwclQ6gSKSnGBqCihdwVlhDdI8KqWsM+
fH+d66X1pZ9EBtzo4VWjzg1DA3w7hE8UJ1PzXvazEW3CdaSczunYNdwj30kUqbpn
v2PNNt00GDSRk+m4njvoo9XlJ7mR3Yb050sHGZBCkz4lYhTffwKjYovO/Jv4QLxh
JNxgEvxsdebX3pDZuWBnftNq+QX4FdA7SHAH058q6jWR74DNK1YV0B9yz+bGO3la
Hgm33ZSfGkEltV6JdFCjEsMC2xG56Qj4eDTor2SDhkURipW3XyXItHhm09H1RQCA
kDoBPrFYS/tXSiH0uSzbRugPMZwpqsHlN1K2kn60GucEwd8aRJ0DuyimP48LAM+J
CKDeVT21vlqvphvZtc0RxeDbA5OYHN6ajhEDxo6+yt44taOPkYJXFqLZoTAzu4V/
Yp/PSgas2WYrZfDVEgctEDzujt7bxukFBjqKjrDVbaDMpirzPrW2rpOhbTBmEdaM
RBpL2ekT6LOTrHdD9yTv0LvzMGH2kChwjxmbP/nj6UZbAzvfa4JOH8EHgJd8Ym1X
uQDDRcaKIkY0qV1iE4oVZ1TdSlwEIT4h3u5jNfAQ2+aWh8D1uscL7IYzhX5I5/8g
9Glun3XlKvEAC/p3eSJ1OKTs8l6ku5yu/v2qmROeqj7bKTFJO0uJruJ5gxED5hZR
rvuhvymDkHae7B7Jvm8ikOnrc2VyGkBcb6zbkWZD2nQxHTlu/eJGEyPmr4u1o2PF
PCQj6BwlF++AtvCD7lgdP3KDSXdEaKmOMA8jaJU3HH+KMxFitD50H84fUbuDKm1D
Zi2wECZ4wn9TmUN3R+bWkW9nzFAXGSR+FFPL4FvgwRw6WmZTyvEMjMrc+oBoH6q7
caZ1ApeA6/OCJsYBYy24wtMrvSej8AkPXZIbFgh86sE5AWTwcSjfIChTi3FvAnlQ
dhn71SYsM7ZRuZqq/o6vI1GNb33hQkDBlzZCxnDyYLmo55XN5TzAk920OL1G+7yO
9SYOOv1oSANABmZC/L1yLHtVt12M2i919tDVEtVtufk/Sp+jg/ie5/9Cvq+MCt86
Pj3kfEjG1vuyegeyynEft3aMUuHQpXNoPZuBuZS/UlrYlsn15yAnJAF8UaccerYQ
LKpTF4jR75mIZRgFCHZtR3dwuxdlMCgJYIOobotIRz/K05zLMaLND6sywQV3HaVt
J79yrcqo4pMi1l7/RJEyzEuywvvBnv99aKHz5BxRcfoTIbGOR0MzYBmcFPdeuPmE
WgSHPw4iqjR+iYZyizgRab7lcdc/bTrIexQoE+XwQyY52PTvhV0sR+EQ+Y5y3D61
vT03LdveoG+0sdBqNrOndGVr6BDknM2gn8W7Ha7TZFsjn4sfZzrdjSNu3Oiz42+p
u2shn2Bv+9r9KRzhBMCzeYeD05KUirYBssHlB/nh7h0vHmBZ7e4yS8t/foeppYvS
TqU/GbZeWKS7o0aub9mgUMD+ExaMqsaZK3rrG4qqbR6P0lv4W2cyWsCEFuin3pdB
tgYbalFU51yFCr/kAJKHa6StmwRcn409g/KmQM7xSWf6i7lcn9DeyvHaRZblz8o7
8UVSCyNSoVru8YCeEPPw6kJEorr4Y0QvWcIJXASjv8yYeknZglLXAKesSQ/j2FM9
u68G1Mh9FfMpZJotInS/QNzVYblFG1QCdXmOdyMTfUKsenpDWJm5qxHsqbX5mqzL
58G2JK2DehC5bUeyFWUMFa+VaMOBOhMu/v/uBuLfru+XXa25GiFhmzLMlTRh28Om
jHM9usynANEF6KnboGPUkU/Zv85q+VDU2tmm7X+bVkvOzHCNFsn1Aaq0NBoSIvpn
5n5O8fAwAMeE/62lLgc/nJUAhS1wF2jfaiUd5BfppF65NKxMTMczWo48TMqNWz4u
bXhc7ZyRcsEJUkkDrowi1bv5GWkIGHocDHfKgB/jhvy3lfUtElIkDBor8WxAeX37
G97l0f9YowxjFUMdV/BCbcxEDJNiO5ZnYjaSML+c9rkgnPOGEWkJ9t1CLdgP4k2A
wy2uP6GeUnfRcc/5Bc3G2FDioTxOVTNi7U9P84iyxhZoeLftX3VE9oDV38g5B1x3
QNmsw+GbsW09yB5FLj+WfHSmFrUZ6JPyjAPKG9SquuqISUEL8td5ZPGUy7CseQCZ
IpUzU/aKbUyQU0SsELjgrlTj+JXqLcZpOkXbNUaHUvFhtXgeuXu2SrHijgS7tQPq
I2wuWlZbvvY/kFzSshacYNFywecKbidoBys/Qkv+lN0EzIGQb1LDZKYFc4Eiy4Qd
5dZCBgTTujdW+fklgskT5zyQZ/bmYYHoafDaX8ecoSa+TGLKdqA5jVKoU/sZPetj
BPxIUR1Vd6pSfWqo4UUJ2rNOlCvL1vsQYdxi+RfSB7zQ1Etx3bYBwNrGpHPZbqKC
WKWzEIfUtBgPl/EVuoQmddFNSfesOQ9Gi0ckVdbdlURjqrrx7tqyYKux+7EjWb5r
U7F+Wxs+dQWd91yMAuCBG1skqxLiySczIWIRXDOi8J1pDwmR0LPkVnBYVdIE4Vi+
cqHLatY/WjBeTzgGND1Ro07eDvvK2TH6poGTCOW/j+0P6Gv6kitf4R57FhW2LyFO
NuwNYYjltbCHVGvUIJiVTM3buJ4q5W/7zSSHq3l/aglD0g+d0QIWkqFmdOXGv5Bo
r1VGgQnqUblIMRIUM7Fks3rfGxMP/U2cjQ03gNNgAeOx4slmbQvrjZk21SMx/HwD
S4F1tJilzCs+ir9arDQcyLN15VtSKYUov95TBh4NZkaBiP4KBtduAiLfdZfbkBe8
B7qBvimnGnxE+921PjtsDH30ztb9n1DkUGgz1MH8Y1eUQVQ/xA5EFA3ZGQGWwqWs
kXXWXlFSafNW6sd0WLOi+8OT2ymp+/G2qYymwa1VGzZG73Gjt4roJAy3XA43Bv/B
6psI5m5sSL5wU5iYEzOmYcPMThyMrCGVAvd5QnOLtKYo04kvisddTWl/Rfj//oO7
uEL6BbMCwrDv5XWWn5NSHumqMSUF3jzpmpAKmRyDqWoCCik50+SYk6v7agqWcxMF
F0YbscR42ecR1b4ZmuQIw46Ex0Y1iAmigk+AoHLjbyRO8td4zrbmyUqRtOTMD8oL
Gbg5B8ut56JwHi2Hct3GvgWThBEaY9h1Q32d94Z8WjbHLLeOLRA9Uwlctxx5+Zmk
MNoYdrLHNyW0+n6QyqypfrKB2Oz/3HfXFW4bjnvrsE8Bm2jxemCOqT0EGFEYLn7X
ag8b4WU/igU3lhUo3RX4Ct/zyZx/69I/5UHo6EW44NFQQvJyInZq4jXrezar8yg9
lCRFXxd03jZVHBrRx58+7rPLfnjtqW5elJzv1fdW4UWgUYfPXHaEKvsgN9A7cZjC
5CooVKV8rpNeU4kme/Qu6ca88auCCmcWGC8m8Q9NbNtHs+ZDa9eXt4lCY1QZKYZ9
RsAsnDMfpWr5hvAa4xn0GOVl0Rlcf8FyHP1FXNyR5D00CFPw4ilNpZt5XJuAWCXf
M+ofWn+0GXZiZBAxV3JRJ5zyE8qF7r+WNjrAI7yUjFRDh8tVmkhI6G+/Um/L6/RD
pJrMYbkqy3/9P/0+Zmm+QiI3NlLQvwYsrqlY8H79GqBBW/Oxe78OxMCeBk2ylFbm
01PJA5EQ6yqrhT8bmwvofeCWfE2tpEwh6HTx5ALwdsBCoHpdMrAZcHGkpAF1Lr3V
btnN57YITPvJk/Mj8vC+ytkM417stAZJnOQEsHa0oGbpn1UySt8in/+l1Xl5dFVJ
0amx6dgTtserKNNxYETv5BXq+AKXhc8W6J50YBSMRyzDreuU3QzRaSD3dbtUayR7
FbcYa6QpqBCqt1HGtcpAJl5yDrGjhaZzzMJvXq6upMoAzjkuY7M3dtm3A5Iu1pNy
oZRN0gA7VOlRyLu4IqHCGXpXopAgDHwOhdgK5i0Oe7ma5UhEHVLooVhB3t9kRrYO
KpfyHCl+HhhY/SPcf63S3SDR6fD88X2J6xloJ31bvffo6vRZk4vNQvF+RlEJOumY
3i3SJIg94d9mxMnRpWl3pTedpgxXuGLxgdTn6Vl1Xb88mywTfoRuR6RrlvvGVgFL
AiacXDr2MKZ1EDZtvhldxnvRXbJOLWk+SPSuVPbBuigKN0gMNS/VnuAC8WznWWvU
HxkBZ114meB9MFohq+/cNrNNXvpscU9H0f5dd6Bil1dw5M9BHwieuMHnMEqNKCZE
fjbpqMAWyPoaFhx8aQXJvr1Yl59ep265rcUq6njJyfdj5SuoEb1zulDUdFJYS/fM
NSrWQ54sgw+ewVS82ASyFEdIqMy/PAs+nuDZFebIkaFKlBQ12tH0XwbdmRkgNUgX
Sd4nbYTjBb26GwE2KmDxbrvZ89HEmGnyd1NfnDlJpQ3ClmrR0cGGZuWGAcpA9i6v
/WX9UrMZkNsQNaCyO7I6rFTe01Wy/9Ogll1fth25asWeUVaLjcnuNOZb8xnAPCUU
2yAHRKJaq50XhyagODfR8SdBMTxvxVz2LPYlt/ViOwhKW0QM5ljBgaJENYk4y+pt
mnq7/g7D5lY/JJs2/FZx/Vccn/iccvHiF4JPgpYMkRxlwfeFefayQJtkzBU4dz5h
QYlbPqMDlVWJa2pysH15QQtM2cGHJhQUaJq5z9qRhAKebDgSOdK4SUoMditIAbIZ
m70JDFmVQIHQ1ofQI7Ah6BAQZj+dt8TW4hq5gstzK9dor+nCZA5YInXCqClHASeT
ABBsTIh5InA4Lh4Kl56Pf8K4s+31B4QZBdLXpe+cSEXxNoRSzKv6+FUtvAxD4X/U
cExL0Qz9ShcL979FvFJ7Y6Z5UtPDwKf1CA4tQc/b4PihEIxcrcVNiWnRjrUdbXM6
kIMjkdNpAwIQX+u5WJdgehDRNtv57QHHIjohamghAk3kxd/g2LZRhgVTnAmexM5o
L7PcAxuo2Yt2fZ0ZbyCicIZoFxL60fmibTNQwWrwLa8gbJ2GyJJKoeIlrNIWNZ0B
JMMtLPweN0ALzfamcNe/Uz6eAO6XN+oSWtJl+yrtENv0AO8cWpZCOtGoKGcm+/m/
bWdkYWXiMUei8xvGBO8frW597jD7djMnSrYVyEoRvKakGp0VqDycDwEtUz80PBRE
Y2Y3VUHQkqfTxaKfCiFkHhzAWRznLr6YbIUUg2YxgaRDdzyvBbYacmMV07fPj5FZ
i08uzG394FacqF5YLRHsomAv8EiWeZYjoUnahp8TXTxzgNa9DtHP8k5Gm9n4ADM7
aVcZeaFW/cz/yYvxzZqNBzODEUWehiBNpgeRkPNwls5Q3y2hlJ+ST5aJtva3pGXm
l6jFAPjYEJVzfPPdwcj5CiQoD1Fq9WW2owFE9/xktbrvmzRgIqBiduIsvkLj5wFC
JPEXiu3hsged4zmXNTAbsMhlWT0PfYd8ter4E+IXSFZC5uG/qe3cke3P2iLLNQyb
3AHJWCEEyHZGuYNadbo83/iTMKjon/7ePv5M2OorQk2oOgbhIh86CNeHSq7kUYN8
z5/i46M426oHH/cWwan62rTmNXlC7nvnwkdQXr7iHEyoc7IfcZS6yf4QNrBOjONe
zuuAm362rmdNorC+rFHAaJpH/QzAYipC+GiTVBnvlTQdl0BLpRX3sHOzd4Sgzfm/
N1tCynktdHjjkFdSXBXaiUEmwnxlonTo1tLc9XTTwPsHw0TjOfgBASFrQ1aCrBnG
0Xq7LF2y84l3z38QovlEfdTdm0K/UWJNJ60KJ9qFjJmYyEuCa/WxAA2flaUjzZ3H
9r9snFe77RRAIUCGVjvAuR0vS6v3J8kPPcc/gEISDWnfZTciPRf/WjXrhIH/BwB/
9yVar7AIDc6Xvz+pZnT71cVvzN1UdiXnhN4uUpnhnbgSi4n2wK7BfURmXOgj99nE
TwKZ2HHRhBZu5K+J1t1ESQwMgZT3Xsb4MqZskR28LrgOydPAFCjax9d7jQs5k2e8
PbE855lqMuBgduQyj35d5Ke1y0grp5zq7EaG0EXSm5IjUrihkK4gU7D6wZ+lxn2E
xLSw5Xfzzy/M0xD6zBk0K27tFOhf1zcpEJWSUB8Si1RiQ1LEFnYK1XFssGyEiWOP
/0uHYgfGFI0i/XJqnTSBwFTtx5jG/GJd6Q8KcyCvuEJ71ym5Q3JKe5lRZYcmsv9r
4VnulrKqku/N6EFr3qE1JzZVt2yMcyOxUIcukFz5vFEPYk+O3+eY2B2iyvg+2XoF
3wjheA4XvJ0/J6wRNb8ZECmYCF6j2yODTD8NvwGEYfCYqH0AnBjXvbyVX0G7L/kl
IhP/IzqVPX30nsLqSvmDuhN2wO+2+0iRpz+eUm6NyywDDg7JxRhfqMNhJK7hK5Ng
y09dft8MMriIAXxwumhHhtRy+QVWwg14MqVVFdyUOTMV8QiJUBUXLK0cwOf+PeBM
cj8frLBds+k3aLdQd9arVfvqskt5TZlrQj5G12ul3u7X0dQxZFoHxCdau6FunPye
L3qgoQ7yA+7MENpu+x19/7DOcNGDdETUD4jZ6XAwDrCG576Wpqdve/Go9dM0d7Kx
M6Xfkrw+EnyibEdsjTw6Wx54ElfgbnyP72v8P6ufBfl4RyLDTLe1isaGIQtgBMKL
nYNPA7kUPUGc+upV3dXqeZgS+mekFr4SO5Zb58tJ+jhxtRCG1DI45f/50sKWWfbL
wosVlWHYx+a8MjayOr2ZrGmW4q+8tNckKJ6RwVvi8HOoOI8oo6MTsZOWJLmaIYVi
DMqVhr8j/uh4bxMnD9+fOVimpjt42UOOGS7sSIAbJQYPN15PeIttlCbzAgamnUCh
RLcN5mKK0WMizoYzBVKvW2Ip/NNGrOXv1G7OJMB13uDlpzWvhntS0OFC3pmeIdvZ
oEVS3N2UWOf9SdHDqs3Ge8m7j32muggMNy/jWjkGTv1wNrIADbSt4R577NSSKCwG
gcp57Q1LcPB/VcUy9SE5sg97jb3D/bWPw2iQy6KrMeB3ryuiQBIH099HleQyrX9M
muP6GuGtByIvB+RgHPKBuwcr5uJVwx+uJUnQe4ULf+OI9yKkMb274wCWre8E6SzV
Sh4507g6oiFwdyC/+4wF3g9Vq/y6g47TrRpjFDf0iZyJ3u+JXxGJg3JEOThJOl24
+3UP4/8Sg07mL2NYbxLWkWpodxKBBavNZTNGL/09ZvwgFv19vhAVtJBcg1LL3HdS
bRUzQq3gSqQtPBHoWSbCp0NdjsCNUspm9I8iTVDiCpqIcHlFOztzeZvFfw07qjAQ
muxDm6w1efpqNGUoJ8QjPW8XacYHydXTWao2Eky2A4pgEUwyQz6AKV0UOz8AsaS3
1l/RZlBTjzniB+brWweT7IS1BnBHLqc5UOOMKhk0vDCCyj5qvGpoK+WS6VAwYkyG
OF9ZToJ3qagUVdvLROcD2WTfkzJeVUGiqlq0T3INNhXi9yT48HKqUwBZvpzC3XWe
cRXwnJfoV7eSJ0PcC7Fkqls2YbhpnlbGQqzpGKX7R/yfFY+PH08dO3Pptd14V1la
OXobq4tQypzDVwSrLWhxyUpX04QhxZLQe1dgrTABs+JOaMtqPHDjf6hHyKtz0tHS
6Om3VC+aOU5GPOlcxSDeW/ME/fwC1J2sqgYkBov0KC9AsMGFLVJWhJLuKNSwDtMQ
vr2Sic6Mu7VQ9CzSoq09HXpZnciCOVA2UFcpUug+VGEdObu5gyfkIfsDtZxpgCO8
n1/2MdmmNtG6IurLYZzMEgaK7cHQvIvGnf4UHdXIOuY/ZsKXgkxpNdJK5IMpe9M2
I/MFkW4Toiwao9g6Hc0ynDW67pSh6PEAgdUCxK4W7dOyQ5EmhN3qjFNqsulqr8/w
d4KkYlXvt0xWJ2KKqkJUl+BnGu4SUU0ggt1HTv11Jn9j9hvPPSiA3OCQyk/tU5kz
6FxbvZbLxkVxZQWI2oh3RzGx+KK+VDR1l74SdVH+ZvsS7bMbdCCrPtokNBkvmv2x
xK5ECjb/nxOuewYZNTMPC2E7PKwX12V4rwvtBExGiAi7iOx0wcRIV1Fy7Jjtx8/N
3RWA69ZiuTNWddQc7S32Nb5XSPsyP3uUh34W8NO5U2kqClxoEHDGIU62jXfB0y4y
1+uJZfQiMT5TXjdvOsPfV7xYLY7zclP1vkXjdCRirqA5i/+RvumtKbOiu1f+5B+p
6MiVKuXL/tbuybZKUjCAZ2KnMA+5yFYLMu6p+/oZMU28Rovn2CHZDY4jFZfAYBFz
KNOmjhAaaRa6G2sPwbsTK1Ek4h9s+61+Mloqp/dIk7dc5mye5Whx77lnq0Jve6oU
7H80ks9FVnh+FqKOqkz0s2JLnm6vzDn3bqMS5zhIFSlgYFKwGgWhnfu5R24qZiZr
ZdlVj02Tef+KT3yn0ftPjcuqh23/TFcJP722XYnYgUxmv53BSnyT5ZEzpRIGfRfG
L1UOS3hxqj8JFzBpJTxgElxQbgdvhPNAx1wy83qfSWdLGQP5XXCqlnueElEZfRld
Qe7/eaNpijhhmSznutHDRxTjsdoQ4SBqH1vOMnG7cUUde/HCwgSQpoFtt8ftRW87
nrxi1dWfUqSF8q+2XB0Wm7HwJKGf1xsr0Cnjts6zhsGsXlsR7OIG5D7F6lEbvPpA
sQ80Bokgeu2pJ5E7ajDcq76TeJJMw5LRlXajw/WSfOS57eqzasjICn0KVj5GtQNl
uAzGj7havQE7SNwVo2TeRdhOOFI0Ig97wSB6UWLqkonIVRG1vnF2AMBV+87eEUMo
xHp11U4aj5f86GOYzpFjpT4Ir7OKzhdPpvExHFDkFS+9QHvEX3Zdv1gzSg7wWaVh
aM7C6e+W+udfcaZTgj3io5y2Hftaz4epdUXRAu2be7x5msrKBLao+GTf500ZbibR
OBghw/5CmAfM8a5aGUfVWlVIrmFsXCtv61cg1GCvOQDZd3/yZKBov5nfeUn1ricR
GnLKxhevhntehHIv/lemWYCZrul6ndRMjtVNyjnfOfAcHa3p5ehEqiT+3Udb03yD
G1CSbJGN9+FrsYI0gnx0Aenj8lWlOM1ev7h0k+EFMHCwKLgtj3Yb4riGHtXqYb3B
JmvZ2REtFuul20MQiQjuSETnBshE6qp/+ieU8DhAvoYOghZ8Vc74RQlbbUWkU2MD
TyNehBowaj1yDUvuB6AuBFqlbLtoavYGC0I/WyqcFczVhRUwf+ikzkp+8rpQV+S1
XH7Y0UgLLfalY/vwPSfEosIc+D8Iks0XAXtvtVIDZJMYWrB5dY/HMp0ons09EO0T
xyyIhtuJHaiEfHyh489aDyCVALSXasxpZe14yrG8STriKzRYohYy+w+q9P1vl65k
yVuv+toSUWQsWRNvkok3oN4NOzvL54C5TcxCZ068GoV4iv4bgEQ4cwvJGnnl5FVA
YXHOU5SRzpBoN6ZtoPAL3TWBswNn1r+gLEEnBkKpE9QCnUXPROm+lNaoEL7Ba2k5
v4qxZ0ru768eL3HBsZuMwNHYUUfENQPMK+Xp95nC9nnrzzi+JEZrIhB9nG5r5OhT
EVc1QavwlPpu6RWNiK7IxFd7917LhTRWq4GJmwVfm+Y23wF7E7/aFOVmaz4kr7BG
Zl1sMQZMyi46DbOCtjYIcsE319/qgJfOxeKH41nE3DHIcZHWb1h4auxNdYOHkmry
nARA5hI8O0lw9EljgLvSDfW2SJWZdt/VAVvJbwkTiA0aruq4hAUKjuLbRqeyfFyc
+GMQSDwfgXtAGsgmA5xqKjRONYXMFe8vt/cesrJunbpVjp/Bf+pHO7EZAEsE5BBX
xfh+FTwVYXKVkF6IQSoCzQ6sPoM+TOpPvRMTtPSMcEk5/4mCTg2ZvE7mvT+9CfF6
zSUQSiI1pOb7ceI9CXTPea0VWtih/rGDeT/aoI7EZEa43DxlUcgICWdj+I/iaOj+
8wJpzxhlqMbB11GdP5PVs02YmjGHsmCY/AkWlQhAT7qrfRNZXZ6t/yv8Vbq/c5c4
HiINik5cRo5BT3eNLMboHd6HAjXqP1T9UOkArkrB9l50KdbEMppTfp/KPn6eutcY
ulQNRd8vgzXV0QJrNc+nI3itscqVkpSSAS1rnCTmBI8+KpKmmsODVoNyfPgAunJq
u6ua23WMQGONDXKvPjCd/TuBEooZxNySYRg/+9rdgQ5LFQ2miug/5iEUbXn3qMYM
sMPH5o2bINB3tBC6v/yzQjk93dTTYMNu8IG2XzU0fSlTQ/ceyKTwIYblV/EGGTGr
tQwqiHZwNEXQO+PTEHhTEOZe9COIQx6JZ1HDGbPmnvXnB3hz6IMPOGIz+4hXPRI/
VaMKkCbC88uxYMIpj0uvj39j5oCTVkEFVWlGNacAl5AkgF6DOTDNYJO2zmPAPMY5
UcLLXU+WDeoDUy1Jy43DmwDBKz8HPFppvOaFHyK+qnjX40uc7l1yJi2Gu5WkvAPY
yq34DCDbMb/EcET4GkMa/ZVFDId0qZyA1Nis8sCd9Z65/QE/4uJDljlI5oYwtbJB
ZtCB1rXG3dKAcz9Uk4t5buernWO/fb2YVy6Ukenpz9nGCNfQNMammwz+zP2NDYOF
mKtcM99YkyaKV35rOgowt64YhTs8njvoHjk3jbw8vyYwIcVNah4YF4h30AHMVzNh
CBEkNE0YNbdyImPVOHb3Yey1w/DJbP4HTb5kayVMUWtyBbtbrbt4cRvp9Jq5xQMS
mG7C/HpEnXqWn+SBSSFB+hmRURBOJyexdZIeOqb0EY35qSPxsFztElA9BsXU28Od
EXO3rh8xw7fVvPDRue7MsQ+Zy2S0Gi5xfgoqz2POMr263HWJVHsrfKp8K2jl92wl
44lVgRO1lQilaXhSUBYr9/D3DiVno3jlOc06jygPFE36+nBFiM7f4u9jmZUxamiI
7pNxvKlWMJhybC7URflHuCdzsGhApPbzrZdegVcsyuEjCf1gsGDAVDgRRYD9qXt+
YDIJ9DfyxuEyttkMYsmyblPb/GMRYjxTOA1AGYL/lhsLbECgyxa1ci9EsVg0o77n
RMWVohfo52XE5Tiewl/1TbyE8VxtL5Apc7CjoYHkx1lbS6VdBpkjrZLRiL/NGAd4
gGV/3FYdB+1zezTbk68ojn8dXn59JGO7WlVgsWj51aKCK6ep7RAGdNCEkqEW1Pld
e2i3aNdIBiBSd4sx1s//YQ+gtFyGfv02ucS7ky2/7PeqB+tB97KcQVDdH2MIvFmT
T5CrmK4MBXQv2HHi9VMEQdixqBflQeMcHJuwWlfCzfxxSy34+qwL6GSItsM810f1
kCqPfJ4n8+DoYP7jtoihQdpXLf8AwYtdb2wOkgyHrjc0zdDDd6uzeOeig0H0/hWE
8boybgA6n4PuJgLFvN5cUnx3vno2N/2B7TwZ+KOJtmzrZ+DoeYZSKMSpqOYaozB3
EkssJO81z5C5dSgkZ6kN/2QqzwzLNvGO4cfX2yIuO2f0a7yaJp9ZpPapngI2fkbF
8bGeryAQIAND5+arbTawm1idqFrVgrzTiVvbWsi73U7PPMj4Ww6cBqzatl3d2gwf
gbFlAVqBW7IOAzn24zh2+GyzDZqy1biQuvKTdq+GeodILTlDK9lK5LZ/SmEgO/VC
23wKsMJyUl8NKdfGl4Zed9zjaEFB4vzw5EdN9jawZUTKWMmyEK/8LGFk5695QMsF
TH/TL+r/Fdxr0N/MceOo13nDJjRpIQjDOueSH/ARGVZqHTyPcZDDtFGesFHGMqq7
eUlXQ3pCbe149ZvD2p2G4BtVUqafTyYamIQydDg6uXXhwZnzkI1gdJVeEWYKj3cG
Xh5Fh5YUqP10DgNSUalHZzujADoaB5SlMti/ER0sG1r1N2ib9KpqMf8FCMngIAGi
m0Iq1uC+O8GAY5sWLUHgT+Fl4am4/pCDW8hBCi82R6jJQnx9TvUbsCvIO9Voq9Zm
KUCBkzScw1hDujN0ZzWFHanhCTL3DBV80z3ky3kiBeWHuuQnQdNqIlh+RoJiO3O7
A5gm7+0krEmvuoGueIgWeZpdnauauuykQYL/JUwcAZKoOR1l8QrUxzybBrSJRfzy
ozdHl0EhQJzCmCsfa0OgbQVnORVNxB/bZCcQKyXf/oDJuLGMAFoUPbRCR2dM1ETs
j+AygpmvmsGWJSAhdJDGk1LH7hCClHXqQwgpr6iUmccYNHkyht7COOeenQa7yPQh
LGgtKOvl1gEoxGIbqbbteqNXpxdaUesGeik5kih/MftJccFvYgN8KjbW4SaeAO7y
IvKBdUp+2cDTilvNowCMEZGR2Q0CXPYwAca8wjrbCW+znt9bILBLPk7vqZYVnlJJ
HGPjBChjQOD3lEwxvumSTIy7fqNWnvAUr09reP4B5vAeF5YYzStPST+aKIPFJS0y
c8msZ74rzC9yXPs1BrUnO3NU2Wt75/ocTXmak1IiT/+18u+mg8ggFtzdF3qtaQJv
98eSrkQoGbabGu5yimUnfl7VZPxm4Du6KxFNgVl+SQEpV43a+7IK9ag6RqhQEMyn
OCLeaZYlXbyhDeYHexSvSG7CHwYV2EUH02g9w72JlHEnLWfXifAYuZuk633bT2p5
xgjwbZ+cVYY2iQpT+b9ZTa2WPKHQWN2JoYuEIPF26mEsrKEkmZmNBjjNg+NvnQs0
rMkCnHW2dqIo6fV7RTJy6ExcabM/VR+T9IOBSchoefarQkfOyXRbv/ZbH8wOLiwq
s5SRIadwa00xhKX4viyoyAVyZYqNuYdy56GTTrnaof1S0qSQoQE1Av3P4tNWkAgz
eZTGqs0ILx9SIiqKsJyOP/zVTkqBUwx43fHlLEZ7N0oJpYIXI9Xb5GHMPyTr81xG
v+H2s2O06jtq02jOthaKPhqfvtNdWDnG6VBGlSoX17GMCyBP2N9/f+y2D1v4U8X9
tFrYM1/wyLbip8vugTT5xrFz8vhma1jXloY0Be6I7x5V3PNO/4wiaiKUbAbSBUlc
fDzEF7BtRKmKzRqHxkSyfnJ7RIBnTQyAHCe/R5OAoWnRSH6h6OgYIe6HBa/oB1me
ADy7Qf7v1ZSvxFbqvS6S+T1dbvdl27q2SFwDs7EOPPfWTiW0LCD2jBAl9y3qlA6P
CEHxDvFF+UxKX1tAgpDIMFiJ9LKVDFJ2dvBwqaAqScvu5Hh0rOH1k49xg1LpNfJJ
xSCHjSdLKJLTQ0SIW/mXUeVn07ee8v5QdsUB0yEJeeJExQqUtR3Ze/ZZz939h9vz
yrg0wh3neNKwiTjrHTb3kHDhkxaatkHXGjS15y7uX/LPr8v3lu2wY3WriBcl1J5Q
WDvsGmW0Xy//7b+iCXD2N1GT6R/FotFqvynvnT2twSlP+g2LDJWva1Yp7q2TLkkt
f7wIyV2HkfmS/IZ6Sri/L0kjQqwC74rJer9diLhhTvH19Z65eQSWQxj7542k2kzX
BKSNPT4aLNVFrByz+x3fU8/yn6nRtQtVmgRKDKN+nrWOhR9nQ3w1wMIPTcF61Pba
jsuk+lRLWl8iqbo86eqR+relyFtbRmng6lLDfipcwQFbYjPV7MPEVLVonbxoKTxo
BpQ22L0N6YPAQb1SmILCt7etgzgcZSBXUecNefXLqTsJ4cp++EeCU0bQqdafBkWI
MqGP6xQH1rRYLCkIBiRjA3ou6Zuvet5fOdR6tyGVEQzOQUcJjzAjr4ecGZMRjGUz
rZTuergRr7Qu9Cq6lqMP9bhHcN0wB1fauQeXpESNj8bX7Ca4gWHFHwtQDIO4PVbL
QQnVBubdOh6c+R9I4n76/x7/DMc5h0sokvAO9++39xfjGEWdV0Y+mPWv4ExPUDAA
pwsxrXmvZQOhPJT830iKKykXXp5aOR/xfllOG0xGtgDpxrrTgc2oVQ+7EgHxjbmP
JNtehIXMvCZ1WGFdF44OuyT7oWj7xDwW4/NF4lEAB//kGnsQ+35UbSq8y3pvf9hb
7d1Fao6tsXdTehP0+oCgs47f7uakDZFizfgojw+x2YJu8zHI5m+1oRrTFpw2y11N
xRnoF/a8EalXdFsNjltJCAXVh639Pbqgqiyy45F4/RjL3ZyqUFAseFc6/o0pFCAN
hAHARFp7W+QM1gFg0wgxk+Wx/9abHXt3YCh2Sp8/ppaT6rV8uEXYfeVKg6hB7jZB
nRbhug6fxRiZpa2t5iiDPUZvjpLDmaowVctZgosGjTUPUAlpcas79Awwu3aoTAbE
4hgtybdZ9AtSotxEXfvSjvD+EAgCDJ6hv3MM+fVFdxwrJwB2WDGemIk6SaD7R+P6
LfU8TFoiBitWHaswMm8dizpXAFdx4+k6A3XfLFQUs/74doAhwuxs/lKDFkHxZD4m
PhwQMFtIqZ8pYhJ7CnDIDhp7/7PSItbuV4rU0EcBim8mvIoJQ3zLPRghMwhgKjHn
S0AZONECytiQY2Qg4P1sRlABsEoKStGJ/SxdJbSfEVyLMW90E4/zN0r/NGYOZwiR
9xlgmBPEwK+2uqwGufjkPrJy1fvXa2/KKV8u+1Mpxgn932azcKvYLBXU6XVuWECN
e4/cVYfnYcHEJHKAdJffhwF898+mitzrBzrZHeJSzUHlQGwzt8E0JzAbo69nxQgb
R2CvkNvyPYO2FXKa8Pxaa516/QZIKjKMhzNTCVR+eQYFjPQ8gddw/qOaz46EeZ70
x/i9RNUTFh02KNOYxEeuD3opMnEJB3JjvbEZUCRJ06vQIdGzk83kZGTR5JAE8Tyg
hxRYrac3u0Ucp2T6xLTZs+U8Ug2+wgukVLUKowMyAjzyDDhfw2lpiH3sh61XxxOH
jxM1MEIvn2uxgN+5eh/kJq1Pta+5PCW+YgvYvJ00BwaKCh3vGK5WIs+a8Byr4a0i
kS+nomzlDo58Yrqwp5K57672STsc5uI/cm7eh7OPb2XqQ6y0XgxHSGdFTUJA4Und
7fWjv+rqT8pchlmRjKorGpie9SXiDFMNS0R+S0B02grLwSIP+F9rM9FNueHiV8lk
p/bGN84+ZhyjqD2dfh3eGh3o70Q/frIQGIO8dDmsF45Af9QTZOn/7PxZXhXrxwNq
iNid3+MAimBpyWEYLZBWzyu0sUlAKJgWuE0Ydc5QYRoFMykMzV+dqD3IabZbSZNk
9fgG5GhdJV+8GrYlvp2555yClmrAXadC64bd1NZRVzTBWKEUF97KonmyClKNrgjT
s9XGjUs7tX6O35BZPYgMEhpe1R3+lxau5xVTLH1dMvMLHYkIafa7bLdM903egX7z
iPMcofefr39TWl2bh55VjI3kvhH7KYLCYR2hPPShrB1UINiCjwElnSYCAbGWESBA
eaRTv4D/C5pilLRDFt8Ie5U2prdQvNvDWM95S9KYckpMMGeZkaRlfL28I/IsvMmo
ppaY4HHa/n0cLovHcRGwTJaJgTGGYrck4EeFkGTrUFvg+l6mfmxR6K8mwA+Nqt0d
XoDzPM14GjY22oEkQxkLXdt9uO+q1GfoB6UcquU/c6XHg0JgFL7IaZkCNGNYyqZC
e3xUJK+5uYKgro80WNzuzTP9K+kuXqnQOOVkcji7X4+omeItaLmiyqlpFoSfWa+j
xet1gFVTsePQ0jW+gZSpA09Wti9bWHBLFoyfu7f3czHuw/k+zm7di3Z0wb+Unyfz
Je4z71wjip7SxJQp4/3MtOkP6qPcw7yPYf0MEVCkVvM+JKmif+JVK+Rp88EsBna6
nQCyFfpYtngqC0Woe8EZEFTEZozKiR15gTD/ZG8f2owypC9lmRngtKeWCtHshzzr
lfrrrB7tcosqmW+Yp37Jltt7V2grNIKncSg2UkbkBtzP2CjDqwOuFPBs8LeOT2uD
8k+DQdWU7Ed4kRPqc20mnU562/0SYH/Ht0uUh4bjCSxmLDlvSZ/T4aNgjozFSNMX
TQhY8MOynLodcXGsakmenV6FbrDa2iv29FJptnxTOWOF8iCVI5hUnM726Fdf2pWW
LC9JtOmehHmhhNxQXHNnaEILqH6a5tuJkvq3GQSKtFq7VlX3JNR15mFGW8SwMMei
zX47n7TVHB3Igg7eeK1/ukKBVCPfA1bg06qB2iVkM9NBXFn1rGsFnZfIPSk3QPsi
gFxW6A5sUvl7bw3ZJy4WesJmVA337U7HImTFxOy/0AajrFeluDn9bZJF/q/ObEXh
IFBqN4tMxxOKwr2Tqj7OFhKadhlLeOCUWogLhlZnw6l7411iDlMjxFn70aUDw+me
FYk0+T/M0Dd1CZ7j89u4AB30gCNplK78KwTx0zo/w4GwTmDRqzuT6l3iPuJm82Jb
lOT/maRNOqjmFK1eQVmViLxLvTcS6TAFbMoq8uSvxQWHGaKrB+OIALSprbTtIDi6
IOAyatNWy27v8p1vOuSCcMN5eIHxioFOTRQ0jjB53DjBfhCjdSTDGcmptgz/2pEx
tVYBr3ds6sSYcMmS/lGV9bDO9u1U1HEavISJYoqgnSn7QJjVmCf4j34XINM7FcCB
yIrbFei6gV+z7aaaG+vKtptzM7+lk3hKR3iHdtp7/KG1F1B6AQU1nXVgJANt0ouk
/oAkJL4hDlt4dCLxizwh7aBDNlDYDrbKB81TTFKcT37EnYL7vWYc+JtsqQBxQx64
/J0kF75aoSsn3UwWWRjXIdcUU3w5jri+dTIQGE9vGuE1UWVz0xaenOcKeMpr+90V
etKwEyqX/QR367JQ+N34olMY/US6i+6r+UCa7KHLTi3jw75Y2gsiGjcEanHvSbMw
1Tcy4HLicNDtDfKIgyxBcmBaoAd6dNQzrPozWG7XFa+kFpzNf6ZjIOfebnAGWxj/
vYlI+fUz99Vo0DmFHWKMjKUiZwc2q7Cecq5MaQ82kD4CbVdtX4b9U1Aq6ZVax8QI
rhnt4IJeBjjoOr7bcxkgkuLi0j1+QoglXl3HNrK19K1kUIrqquSvaGKWuh68zS9O
BSr02Qq7rDGER+7dD+t0XSs5/sYObHCQCJLjJXOo2xINNXRWCmHIyvGNCY5vskQt
gGZYxmnpFRjF3wdpkOc0x/tKHQtYotjdjQdtpBcpQm1bgJ6s0xndxArGwkeQbKVq
UmT9gJtIKjj5L/FhX7fkCr9kMu8/z5+Jq7Ys9zGWlOBiNZGWwQc0pDojFn1X2Fwy
Z3BsrE+ajm3vhyGKMxIjLJem6S1Rwqp3wqu5XfftroNWgLkGEyQsWXk6jAYmdVZH
rc4tpfzOCSku/w9Dka2EYkHMjU1M7Hy76Pbs+cy/skrvs4x5E/K42l8s29LFKzbp
o8lgC0lTxZNgxafyD6+w6p+sK6sg0ZRdu5fMQkMbKFQpESgbMbw7XZr4R1mWk0TP
8GGeSok1TyTZoV08XxSi52HPP/6qZaZh5Oyvp9jo8YmywTSvsZWLdnMYS/ZNAXQQ
tW31TNebiZcxr/0GcDWaxmA5SelIykfRCrayIUVopb6sdKTNpgjHdRBTedTIDU5+
6c84teKbpmh1HpNGx+2Y8CppVcW8uNE8vBOUrW7xvy1h8HAHCr6hNSKVoKbjYKpE
vkF2tMl8FcSTF0AqXiX8YI5XMNLx8Bre5LJE9BbfebNkV5XAh1k8gbTh2u8+hq2i
3wqgOQOGwsyOYv11iAdNYge0Ma28D7BROicZ/+gbuditql+NuPwKEQqFHxrX75Sl
Bpoh5oDzJwiyon/L/SzJhDB4kTr46Sxj9VsjHHC8l37NjfMkJbMPgibkzv6Gu02c
SNV+c2irXU5iY02c0Y24oAQY6C/D2LWFlaCEbZpVJcpGQSmeysE9fdeVXidh0vz2
ggXBzjW9Wbp11FNdT1urU+dbCL6ldWlW4VQD+1KXZGZYla6dLsFLtpghsSnMPH4r
WgznnAhal7oGjhErLjGEGS1kFrtXKLFS5WRyT0I+bHHJp8zfRZRMzXbjQvcsp7me
ISC9gSdMK5axEBabKk2IC9r98XmJbsdIGbadXWolhKd7F5C7WCHDPzXaZP3QfRZb
gPQXBNWMzikpjYWU4bVuTg==
`pragma protect end_protected
