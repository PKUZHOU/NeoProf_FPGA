// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
AafzmXav9fsPt0XAM7XNQ6Z88tWZ9jIbeG62ZPgflilGWa0VbpxOgofa0/8gDMNb
nmD6Whvg8ccAGvsfa86zM0umviibn4bj4JB2gO95enpu/vq7pOvxywWvAxWmimrm
zY33st/IT9FBgRTrUGSgKFMtbel/rwuX42NCy/Q5T4M=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 1744 )
`pragma protect data_block
M7gg7Y0yPKYSY4RNdmMpvQaejH1HB6Q1UihaAevhYHH99wKCSmylRgUzAc/e/nMU
Auj7w7oRa4gpVH5PDhNMM4DvsecGibH7p6iCAmbl4AaptC1H9/D/VFdy+k166m+F
V2sose0egw4IA+dnQAqHiNAPixXUpVJU8JwJVldeXVFIs6+aaAsqCFIrWTiCuW3w
ft11fOTVJf+hoCxZaVeIztLxT3LflXm3chyLBKb2TjzIKB6wuY9gEQ7CxYDiABuV
smdNNHaZI+aU6DFG2L6mHkE+sJQkdfwO4uBWQLc7rF5I5pP8y7WT4+GurVT5OX9q
jKHoW35uGsyxeDNL5pNZuKq4tI2bkGLb9kzbZESS2I7rJr6i0SH3V7D04yGE7hS5
vqACdKuGptZDChmsZt9ONdZjx60YCGjXaRfnbJtBJlcNtvFEpB/xiz4HbwcgnqB1
2Edxj87vVGLby4zGR+v+JhwkNz5fv1gV/GduXO4gaJ2PB9EvndjlCcUgBrtpV932
KQ3UTkgZjYH4X9K0N4m9qKNnPgV062uQhu6/nT5BOw0dSFopfleGEFhejgZ7ESnc
9EF4s160b7/rKCZlUvNT7iN5u/bVbZzspuqE2FC1MssRZdyoGr4UTiKlx0z3v4Pd
YRZxUMDhQDI4lCQe51+c+hOAIJoq/DLmVGDhAENUf52//8mdSfio/2uFy9eyVy06
Ccqgz/mFUJ4SwO/rqH1Au4aMIPebvvk0/iFFcg4HaZpAbw2fqLOtP08lpTL5TWDo
ESK42tqHbGevBO4uHkKh6kh0tAN9GpJ5x3vanMBhG24BtIWAyVe0dHK68PcEb4Qe
KW7YtdlPC1ImyL42+Uqf5U5rxb5gUFISL5I1WzZElcFzcu19i9Xd81rH9PerN/hO
ytfA3J4IN5QMfbMTzMT6I4yqHVzt7lIk+MywgpTzNWEXa+fjm9BrVzRwixQupfuM
5pd3BGdqVLmviP0yQVwzSLajvpxZqv3eHR9zV38r1Fd3t7s9ClteZK8hhbqMLGTk
UOufgpcezQtkc+dV2gr/6N/M7c0Pbf/fqS97qrOeZRaUUyYjPZwGd0qW3OE1G3dz
feWOAmfaAvJSe+nco6Z2BGdAjVg2a+9aURgLYNcKkDBdtlRuvp28A1OiR+1VwLrn
zU2DVZQKIKuPqdxCJbYQH2qXgdBty3Jtvt2iGvzrO9fH5VML+Od4cEPYBS3K8tMw
KEtt/ZDNPRBfjlhVBI5j/e4Ka2Zg95e9v8J/tokoMc9aUBOJmYKjKV/hbhrIxMvF
TX5jIGdFEQwxANeCFFWLsB69JMQYo2BcXLADf2xa3egg7RwHtcj9VJIw//35P1iq
cvc6EC+guxCMVIGDSWatpzVY7PV6g8t0dlCJZoKnMUzqT9vLA79EA5qHNnc1Eeyg
HeI39XoFGd7JTQRT6Uou6ouO2mslTcYrbIFQ9GtP1sGTbqs9LEBlMu6qjULTJLd8
AbLNzRUpr3OPRgxN5nWAL7vGdj9ixlbK9EY/FdeMvsUMnu8DjVJVYfEcLwZlx9xC
hphR337u4z1Ujpd1hhPuhKRqIH6pV+uY3QSN6PmLAW7AXecv95x4FNA0LbCsGQqa
tezE1Rsml6ErNJSDaIBQ+d3XnIHvaUiyyRP6OzHzdaRwCSy4dCnpQ014J/+IfK0i
xkrzaazWNUscL+6hqWXr6rhJem2ik+dBhiSDgxV5p7h0UzzPQIObZgz+0xTpb4nR
0jZnBeyKmpOaCihEMoaRDgzkvsZ3YiJ4MYuqK0gbkYhuOLfe9cvylNSSc7W3MvDL
llJIwjqirkeAoLyD5QSLlMrwOwgSszCpUaCACFzcPi1F5wpeORMLauNE9ASAMadC
hvuggO+DFisfsf6Hpu0rvd6MplL0HONAAxmyUM5gfs2wyDElZYeV004myPQy6tLs
ewXghJt6rzFxj3Zz4DYldEUYjETqAbD5HBYz3/RnsrWb1CYyeygbzXQ5NhwlsURi
m8kUuJbAfN6wvnf1nEX2H8gS57V3U5t7jJ/yvROEqkURDbk+PkIqzHGEeZNLO6FX
f4gcGtiFUhusXgHvnbkN4EcQ7V4iW3eznXRgniVpqJ8nMnxEWlNMT9BdpssIzOea
M91EVJ79V393JjoPiXFo26qEcdyR0/G4Y6PNQKzUjbN65J7Vg2qVOgWPpq9x8oWI
TR/4oekNuAp01fQdPvrYWbOI9bDuKUSMBTYK9Sz7SG8VSjjKWKLi3UameHX8/KLG
c1h3IX51okCvuogH4Y3VgnbfJecGBrcWNGkTAyzGGbypHfyNyQVjMR6MJAopNUlV
oDn88SrOfQWBTPdTDt0vUg==

`pragma protect end_protected
