// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
iYpoIWROhQXtIHuTF12QT1jvYliuBVVOrXU4o+pdfl3CcQtHeP+XXujtKz8V7FUA
qa0gB2OdjvAaedblaavzXPM7SnNUfpdC2RDJTPUYh0YoV3rvBEpZSsDvoSdv68Ea
kdWOfB5q+JPBVq3oHWipmoi9YGz0pt7DW9xNCgNFs2A=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 31408 )
`pragma protect data_block
TJk7WaNtJnhr+Z32qOkGuvN8bnuy2ZFyAMp6IxVsslHdrIxLtLMo2ukU1ofDFcwW
iCBATbS5y6gtvjPegMySolThA1let8uH9/QHbjuTdZeRRp35oHF02A1FRvXmckxk
C9giZ1cvKnOlTz0cpMZ0j382NEVrNsHG/+T/pObhGqdJBs02JPmEq4hem4C6tID5
KLXtegaEbrAsn/2ArP97gC+KnxO47H1MSDE8cHAQIp3bzP1Q3aZwKfIq1l9PuP4F
kVpZzeVcemQc8TL0sTohvA//92ruGSwDLl5dI/YkdDQ/Zj6B0ozmOK5Sb/NXE/sn
/SESTSIQN5+OQkGvJkiP0G5BY1FKb+bHxitOgqEcz+gRTEVfcJBI1btYN+wAdLc9
GAH0JBZ5KGjiR2ZhOyrp8QT+mcKjZ9qAEcaoZADABYTQfSBgsFguX+F2RizYSv90
ZeDAPB8L58i2m8JnXrcjIei1JT6MNFl0XAiitQRdiErDnO7p5YcXEIBhqCYt8dkA
zgrJ+IQNYaFCHYWmsZNTZAdrRhLZGtsL7LI17C8Dz4ZeqSmbO8B0mZAVUOiXr/wo
LbDC9qQkFq2E/ZpmL5TNneiC9E6le6nrKmtxtFpBGp5dCW2/oJw+zQYdVObXx4rl
s71wwFMULcnMskoZOQ8F4jcNOIALCstrPPnDKRDTIi01e9lMjMntA6Fm1xZQR5Ia
pUBkOrRKshyumQrzvmBgEpSZwbWU64P4xI6SXmh9DpidanCbPBidH5P5ZHPpTA36
5dy1zy6lJWt09FIJc9m6wa4n0u69IgelOPnjdyMMM2TRpSbK5JqHKYEp7yyktHuT
7cv0mfjqIeZcd/AAJCX+yqVhUYocWQbU6vvxztwEZtyx3GlHwT2oS7zp/Myty1B9
5tZgeK5ad/jFle2j0Ruh1L4UzI13Hnf43yKLFlblBZ7rdXKhdExwBjuFlHBg0wCb
28gDgIAh06iuYiulAsesyw3gzKuyCbEwYzu2OVil1kZEgpebgQLnTbPPb7RtM5ej
6nrRzSwtWL6KERNn1qu9PqpdNePbZvLqHbYfQPDgYSnotGSq5uf34IzCJj2+MhRB
xSKXNvOSsRPXocW+TJaFlbc2JJEJXakEKxsm4G1WbzRYfp86EIYv7VvuCH/iXtGX
KjQ1K4GT4u2kEmI7MsZKIaJ84AxrMBV6/OrX0DVomR6Eqc7K7ntOkrYtZRXbeCyr
sMEZLfTv4OtGoidfevKQUvr+/BTojkiKhQDMu0ZlBIyw43f1/UuPwJuQ+uRVB9Xi
iaMhzQug5S2/rdp6DTyAMgC+Se+V2sqAznQmec3hzOxR6RYKcdABZSMAG+ew24dT
wTHHcMnUXvkYS/wXEIDq4pATPyT/0skPubW1lrNIJm5V70NBXLmP1H4FLIafrl9U
u9Zp06Tmo9K/q5Jgpx/lPC67lbt+SAL5iQOgCpu0ILeH7fd0buh/YuUXjwvNSUkx
+V3RnQVpDGhl+ESwjgJNNrLpzyrbRuye6PtMxMA8k6z6lSVSGracxq2Sc9VlLkbo
9s4+LXwNaNNFiCGF60hL+VcKfcyX0vLIOVCKoz6PPm13fu9F7HVVfOFqtRBP6ETw
r3ZoWDrOw/0CMOjjHAB38dspiBfKX5TK7IoqC2YYofhyYXpQH3Z94EXmPje28YcG
Tw4McBXcPvjAlhB/lYG1lcgCM5T4dDw0E3mWqc04ehIuxN5cazcUagUDSSQlu2Q6
o+XrQqP2u9rHQseom+KLhi0I2KJExe21pqtVjAZL15zou9YCXYo5956wPPudq3Ap
gcD8znApdGSwQccQFIthtcHSWlleLW5hN+VvmQH80MtvGEoeiaZMHNxhwfTMcovd
qFR8jO07s5ebK9bvebpbrqQIxkjsPXqF6lrcXc1fp6AN2+9gErjZTUQpxPEO1NoG
r6ei9rknroOJ7jo2yCaZaC5QHBh8Iwhh5NDKxvARRexwaHzSMNURWNAvBGGYEUok
O/YNc5YcoPf7nQEbvuHhXJK202N36lacBc5eGiE5lx6vAUcEnpkZrF3qv5KXQfcA
v1kJgt2voLfgokeoYmRRW4xufv/Wwvy2LIWk93oOdof6QX4IXHDve2x4mjX3Pjog
tFZmiOZ2aBVxLQFRbVEneom/zwBmy1Gvi74SXopTWj7I0T2U7P+SjDZWj4CARZrj
CHe52Ip0VJID2IdHAL3llLN/tMZMqcAbOcALMagUJeOEu3BawUzCfYpo2MTKxWS3
wCgLxWxVVTRv9U3COjTRCRxRPfWzS7bk9Z2+r4xX2TiParqgWlt2lxbljOF2zAoH
wOQoglxO47aS+r92NqMoPnT68zXXJsRh8kMJl6vQFEQT557Q4csuP023aGWb53U/
61EfoNvw5FfxbMsf0aU0bhCDYpMnkzw7f46iDza7XDxWOSmKs8ike3c64Pq+7qYZ
MjFIH1aFHvhpOGtnB+G99ta6gzUy96nXBdHoyHIOKgChk2UReSfTyMRQ1IHrP1MY
2BgxBh+7OWbsN2GLUt3j1vcFmAdqQFOzkNu5lGl+/0GhMoayZPq882T+SUihUt+/
l6876O3G6iEjGrr3VRb9MxCKyfjnxQCuwxZhfCYplYnCGDXWQvTSyJJHCDKRXCnW
TBgZPYbfI6468bJf3u7KINgFbd9qhYkwPRHfjhgyGWuc0OO6H12k0QG1kviyi5CG
93CgfG+jrFB1Z0rzWIL0JxYslhe5EuZUZOTFRq024k8eSMAcuUlUyl10eAHwPrTn
7MvAmzuoE+iyozVlzFCU3kwrmtIsWWKLB0sRNVs9e2WCBINNE7gvQn0HuRlLL0mv
ZnDL398BBU/OmaHlYol3Bozjrw5uGVTWT3I34E8vejHM9spVNnXbeBEK8RHW8h5P
3zFpKAcUnmhVyoefcSY5wwBZK7H6JWTsgiwCi/MeIh3CSTGVfqNhpcWQ+j2CTsbr
5/g54Vla0oDjMT6jilUXGL7SPte7nZ1jN5+uYtw3QFrYmUbQEy5ParbdKRRYNkQY
tpaNjVFm92WNj1MKveptmQO+2CT/EJtGAm1UgYsvDWqqsnRrVoLKh/3nvISPWXQx
1j0hLQRNo+SmlQh3N5KSljH0KyyxwuQXXcElL7xztTKa+oVAvvyU75mrUbASyR7K
BRruVoBFjTBilzqreMIWD9ZZE8IDw7Wqe5tYP6nQ8dVejDWbvpm85aTn9k6bBNjt
vr9VUJHncnuFgSlXiq/TVJ9YftUu21WpburD1ffpsGLZwy0dVkDecgqMUV5yjqsd
VUoAaP2li+RxeoWcWskcq2leeuCTBm1ZA/lrRYAT3nmX2Je+bvdy5EQgEewAZnA3
t6hxHyq/Dnm6iO2lEmQ9rujTmYBWnfJ+jnAK+55rD535ZqHE5Jy0lLf6nHEntUVd
di8YmznUm169jWWY0ES2f4qGrhMrr4z+BHtvk5vc+jOOp+vYI5v36IsAajYDAjol
E4iyYBwzRxFP2NNbESAAKxfLy4QYc6itXJzHMtSy04M17LjCEdXTOlV5tDQcZHCU
akYqS0CIBt9AFeqgv348BAy6nK/t9JATw6fg6+pWJi6etG42z0avAf+h5Ay7E9uN
FrePeSXcAQJ0VNtBOwFW94PV4XkQOsB40/3Qwz5RP4UT2aBkP1yZpnmsw1cTQRu9
WTELqJOguYp5SjyxReSFnofjeOdY3ZkF9uEqivcacV61fk9INGghmj0kMqpS1pCF
NHBRtnxI4YFBWwh1vTXfNlK+bK9hJGQJFzRUF/jjesfpbLuCz5/NM1tFu26OTaiM
Fa0LWGsRXZtjSd8nSSrjUjam3kbG+S3LPxggxjYrluP6m0hsXoIBpcltHiZirN9S
1h5iCbL96L2ITKp2za44rvgJR7NA0mtcJdG/pqlB/wiTM/VKbS2XUDgPl2ci5vV9
JBP71Hg+LqXVIAn49/MDB+6BcSBJ12pX2zT5l/XZ+J5yKnTZevJG9lyYYhPdZ+nA
35rN7UPeg8rKhOnMPRYXRlq0pc6cTmf/NM79vZj9fq7P58v7gajywVCWHb58PfrC
qpUg61PISPRUw5z0MIUZjjvfIwc8GguYleY/dNyHHvGS7SUuc/xlGZpa+A2zrsQN
jKLdUBXSTacSvGIRaLuYpy6zmZwMoDp09pTnFRADDEK/w349oBW5qDxa610skiUq
KV+BIEr3xVNGyErUFBLAqy+usIDYKxTh3y16reXuzETbZ0uKNuiwOwa4OCeIHfnt
NHyM0JI3PIyT93kT1u4ixGFE2FWCg2xqIMkfsOqIcQ2fPlj67JQQmi06cQHhPpKY
cNfsQ8e63TvZ1wF4SxrYUDF7qnUsEBATNIpnLJ/Xi3pC5WNJqxG3rhvGt8G6eiiZ
I+Sw/XbJRB5flL4+7Zj94boBeXU1kNbouYZ9VWS1f8pO/pgbgLz/PaPjmStU0dhp
cIva2ZZ8Hv5BHoecyX2lFk///p9HvG+RWeorldc/aCziDf1fmEvc0iNmXRw09nzz
upClsiTxFZht4lqa7CFiuCyTIdE2pg21GDgRto53LO/AxnQzrOKSxtDEYio644yY
eiOzuob1IuOEdp1uEFkqFyCrPE2TEpH0jrY7qa52+eE7/BVQJI1VqgaNyRE66Hos
XyRpq2zknCAyClVOZI+7mp0dbTqZiVxiurWGVjVG/ZGxNyl3z4K7nIrqGos10+F8
Lw33BqQb2ONAhuyQ/Y+ooqwMRIuKaLR+BlAbcSamX841F1BYtEXFrRWWtxXMxVXp
Y/pNX9jVDrSW2ZEBGZY0EqTg5BET/VO0+5Xr2DSCg4GcZcD66hGWgvKyNorK+1ZC
zbJargaT+4ido6/MYNz377XIUk1j7lujpO46d5MTtGCEnjcDsim0l29WaMuXnm/+
OMNBHdfBi3bc/Sialro6oDHgPk10Tvz5S222wopeiX3F1/ftlniZQZE+w+9nigkx
GiDylD8L+X+/bLDfVrCspKuO00aHW3teNOqVVZdx3P7Dng844BleGHtHlXCHi4Z8
RcEEinVYahKZOY4zbCQGFKZAdhOckUcRoyilAX7rdhH69iANMdhNqogWQDjjvTjE
tNaqQU80tO/gSAmZBk15qaXlrShBQeBCiAV/N+Gguim9I/nMbLPcQsP9pgmVdUEw
52o9Fo9QUVfPp0RIJtwC2rh79nNAHUxk/0WerZtQWWMfCX2ZeMnOWjT8t6/FzPZC
6hYi5EhHABRzx456gjfb4W0e/C30MD1pn+WCPnBZkg7bslUoy+prq+vT7+0BI2hC
ZwxNYUGBLr1F+nVbBPb5tdT0KC5l1xd17dF+5t9ADpm2V5pKO/I7O6OBzd5ZbGLY
PWDM2nWOxQ5k5MQDWO/X5darbgAEArGHPXyE+tBwaiCT/bX3e2cAwT8iVPtc+eQS
JgEzbZDHqtIY9D/eDTpMt2FEsYMIAKV40tiQH366PW2n68fRhvc90Snd46G3rU1D
90SBRfGWCeXE9hes84I3ftEHoIJmtalpC5xL88+UtO4U38kaivlXk9mR+OqI983P
KkIKkndGHVYScEd+bdhgd4/GRbfT7SR3nVxd4fpX63k17v9h/5Jx/q4twSgj1toD
frAKCx99vjbQbNzbh+jTbM2WforLqoyn6GFDZ8GWA5PXG0ZQuoyzlJxflt8baQAO
43J0WIL93SKDt2kxib1CS23q+t789/HTELjiNvtiPMKkbH+rBxwO7KOn8aCXcWHy
fcnG6pMOh5++oHxqMyHh5wHq1bN4rHGLpG86qy686u3t60qR291XzC/nt/IzsZkd
kW6FOFFTTgokzK/dXTRarCHaiBbKssAYsN+ZAbSpzyB8lgskE/Z5+lu97hwSovm9
8zFVqSJrL+crkm4E7SP5gXB1CFbxr4yj5YYsVM0FaZf7/VftSoQnb5Epfd0uI+U4
/lUpOMdFWqS1YZlTM+OM+xepT5ZpSAIaSjlTbe/WByUNoau5b4INpYQ3CWtIs9bD
S5Rj7445znfmWVWFXjBzMryNucgEmGOwHKFrdFgL7wJi1RQ+DdMovraEUME+tmF1
lyWEnTr9IohM+HasdO3A/wWnDf9oG/BjlJhWfBHYuWAjIJNdu3tyXzkqhhRPbC7x
nSFBwkEMeHrGpWUv7DUuYvJ/YqWKoeOQqL3gDEavs1B6/VG9Inen8PJUT0AFXXWI
xB7GK8TFImPgpB9zofTmL8oWnt2X0FO9bHI77Jbt+Tsz2pJvbuLRO5AjxWnoqzkf
cfBa/YxEe72sJaj5v1B1tL4Utnp0tphrr3uvEd8k7vbX8u45bNaP3Q13r5c3+wcQ
i5m7pdhA5HmFbIngDCr6Dy6+h19GGQzwE6yj5qy0zT/sGIAEk08NwWmtNIVpEf7Z
pII2TARr2xEcsctgFxp4gl64bkVCUAPJU1FzI11C7F1HVv5qfETspeG39E2pksp3
BVaLKKVmvV8IHFy7s1uShrXVlX7Nonadj9+KH2eu0h2tZ7Tk43HwQLfufp46iJy0
DWnIIeYDO8nIMhDc9/oSo2h2aJb3/1r1YB0JM56lDeoGEeq2JCil5jW6gHnytiNw
Cmgmg90kArPPtKj9CSus0K9CbSPGKIfvhqfII37VkcPW2sjALg1jX02CuoBDYrgt
7BKE2TGVN7iSkndvnVZFaSSFZznmLzd7QEcuioZ1Q1G72fBbWdcIfo3SQYS0800T
Gjr9AW+NBy+hs1x3OpbSv9/wQ/rrtXVoD7jjoNCjMYdF5paa8kb+ozUNKYpq2Wsz
O/JpkpOqEPCD58ZFF7ELvI3u5mtU/KArF5y65nO1Ih4Erl5kpXVarTIuCCHhg09v
vLgjiRqn3rWXTW+YKQN4qU19Z2fwZtDUp0JpNye0PehJxN/tZNS3iwNoDFACHEm1
Xs+1A7hpvpW67Z4Ye4AbYy7BlV0Kxsz7GG4tiH2WEqCtxeQn8MD9sUVwaDBd+A+1
KMTOH2J153JiXgA/a6mpp+swxAyCQkSlkb3lVvkratrGhSYdC5ML3OslgMIrXNSH
BIziVo5sYLfRn/lRXsxxp6XN2AIi//w7QheEWAg78uQuLxVxuY8Wr61DPIwdHpqZ
eoVeZi8hIFVuxhe506N3FQC75YPIbXqLEj3XD+zu/MOP/bLpqDzRm5Ni/GatarTm
TeTe3DlUwCIz4e4oA2OODzqYAptCUIq3XP4I0mmollpkYk4nPyLcyyZtzM9Pz9Zz
YPxuXqgwocZ8SaFhdU13k9EjXjErtXa+aphsftsz4+F2XVUZ3dkufB/BSkwH+v1d
hvxuTL2numsWCNq4gm9ib/ZrzO4IjjjLrWlhDg6Z3KB8unVA3pPlwtCTbobu1GGL
vcUdh8syeDayDB6tkdFObhR5kU+4gv/gq30cKlOqKPbPz8dP/s2pEYBZIGi1TCRW
DHwnckv8QPOQmBlncmBJGnzC4i877x/sYB4oBfOBZmT86Ecl0jWaat3IuEUNgx+3
25JAu6jYdMgdH988jvPzzrzFGdhHUek6fhaEHQC8CyXWYZkbDjI7D70oz3tnouV6
MEn921Hs1LiEdlwzPImTUBrM7mRm8OlqMeS7bqjo9GdROy1m1n6wR09JJ0HapphU
gFwxgmrEz5yPjOpubWgCc2Z+PpBKF4iucRSVom3aFESneqTNucihHktECfCTUfJr
k6dvIKpv0df8x2sMUaOGrn/97630HSe5BvN2U7xzzSgEkoYR0DhsApchqx9m/aJV
2z2O2RWdfa0YVYOCDKrMVZgT+KDdxAw1fxcKCKjOz7sQLgV5p+fwR7L0w841GLrS
U+4M2R5TmNn/if26AQVfHtIMuAQSeRKJylAeDT0d06Y03OFnXX8c3IP3MaS7iU13
b9PSYs4YKslq5/ZZzQGnZUgIR0muWHfn0uZxnjPhKsDk01rDQABKhsDSiLtb9HLn
YT4gGDxErtFGVKAvFakmLeg8g+5LQVQEUlZiF9VbgKlZzwtnIMjQgHrkgPOECAOz
upNEIqLMs5Pim0sF0SejcUN2Tb5/lb4wyW3aDrqHa+BgjOgOh8n4BiYn+voduyQX
h8r2G13bS8EF1trbPOdkaNUjWAAvca/0dR9nNzfQaO2UOVfO83rGasznUsGJJuSg
sAHMIR5SxZAzfb0fZBdvGX2OxMJMqJvKNEVcd6DlAZhdp12tq5P6JKO+EmeyNHv3
thnHuZxCq4tySUbl+avDDvy7P3WjENdiLeoKyVKG3Fy92H6SqY4SLknSWTiiLEWv
+Pgm5J/G16ibLTLHrBwPL1YTEYt9dBw+G+fvX1CJO1dvfGQ4g3BZ0jV+P/bWbOe6
pJ9YcGirA1L5ffTJ0JJO/PMRU5d14fTFizIPUMnt2iXJ6pFMHRYLWMJ5lApvtTVc
KdiJw0A5otAp5udBPesq5E5IVKQeqLwe+6gm+71/ucP55GfwcHMS8DiZBWIEJszz
Ns5Oq0zRpoIDhPw2zI8d5Vk0sGvsU7tEaICzgGUVBkGMYgoQcuKdsrEf2WjEszQG
JngjWVKUsTWUfsmq/ZKFkNrrVfgkjkhLvdZDB7HPTRLAa6czSyjfmYW3BdP9ym82
Cf+WwDlRYdjPjYvByE9bj9Z4pyYqT+TxcY1PlJBnl4NYHs32IayBrektAYlFKpu8
f0pw6U9Thn3y6mT7YWP8zw/xapmi64dBTZMMVQFTVtjKz1FUQqHtMeDJAGa1w8XA
AZ3hI1j+pKDgOsw7SBDASPZsJxiHtMKh3pxhZhvYzrmUC2c3GNv5SfSGqo+8vIZL
rZrJ7fjeZpWQPgF6HpAhv3N2T3JZiKcPMuwn56RVG6N86KRRHasa1uxYP1u6C6+3
vRy5Bd949WoQkJwbULW5IZhWDdtTP3gwKB35+rrUddrxSBrMHrpkwniVnsa3xffh
QxrBnyHk+ki7+EmQQMtSTmHqyi9VaRr2mARAVCIFr6LfWmMAOvkNVBmcWnkGyinF
coqRvv3HXzzx0cIWFJGviyy8CjnLp1EYau5wmUozVpcioEU/u7odc198IyiUulP/
7FTh9bx3wRfVqg5ZqWmu8m6H8cl/mCnoA45XOkOD2p8iNlDOL9IpDqowlCcE0/e7
7OWKBYV4nV045b+1/8Xb1e0c9tjycRFJiWLM3mebLdlQ0DIJNPURNoH0DGX1uKye
H6xFctngG5WLmTLftYAIYgjFAHbrlfgbCin7ZHLCWPHXADv6lWPT514E658VIta2
rpHc9iKhmYncj4jqCQ8MeFLsbu2CZiNdamCsFZS9AOmHEVIQV1vePMI2+7u/UDK8
QkTwKSTvqzvAy7ScZCv30gGFa+sDZ3ONJVQzsc7iRzKeT61/nsaJWfhvWgD9vnQN
Y6f3ZAAsIFw5SD1SyvqtOOdlcuFMSsueUJY7FiTYlOEXndsGr+3ZQr8hW66D/O2u
hZDSJjj834gITwB8mLjd4k1j9Ezeayf6aAP4TpK4mf7mlRcREwPfHI6tAiL/ms5F
qaTli/n9KhT/vL8fn7UOo2/r9sqUjR2QRTcszEX+OG1VGtk5Wz8SYGYHbuMyk6/n
/AiVA6DOWhoyFCPezy1+NnYUoc++6sCXnjSFuaCEwEsy3od+eRT85zn8SADPNhio
FXSr01aWBk7PoSgnwq4H6qivR7FrjNpPcstApm2yi/aODcNA0PxRr3pYUr5CD4BK
BSTYh1zhfLzenA14hoNwCWDJFKpGPc+ZuA3G5/e0xRfZ4bQIj7kJDsPVoTVjbF0Q
T7NUuhJ9Z3edcA/mIsMwFViaKTxDrEBXfpNYxed2HbYzqnycjlaCfrS6x0/N8aKl
opONWZTDSbn9TGaXDHb2vc6xqvwNEmPDg8EhdgUtoy1pRPpvgTx2Gayj4lWe9i1S
tA7T0ID+amC/QQORIPRQGt4rc1eMf3pyQ7f5Cg5vH4mfSGu8J8USuxdGJ2VBC9Vl
44SY0kPOjCtTuvyuXa/5mnUmEPM/2mk5IIdsFnSsCgW1dRosLeRH4i8ooWhtauQW
yXKaNABDWcEiRpW62gQAiihuz9N2Gae1d32QSO/NlyzpVXfUPE0SEVgyWq+3MYAi
DU546EdrmzYKvh8C6gwXGTMTqIWkYwpAC/W735bP3przwPPOqBVlw3XYzbbnvLhe
RNquAWwoas1veFPSLADjPKx+ScsyiWCE8Gb8c1MefL6RjD2MOhNokkJm4xadM54J
9VmFXLRSViwvHPIN7cfsUOj2rzxLnSiZmgs6rlMmJZPlSFH/e+9+lWcI81DDWj8u
QIjAiyugEsKZxyTOcH3ixZ2Lm4tZihqdBWIk2t1AA797SmkNavKTN7mBViPqma3m
MVyB+gkXlTKneWSxcETV5DrO4E0yacN8jA5Enj6epDPFwizXWjgJL2PBGKr4xBxI
KTq+fKlaH52Mxtk61buP585vQzHH8Y1y85VvpwATUIZY3iivxBUkAREocn6F9r6W
TbtYVhEO37haXIobsbfjec+XOhtW2GZikur3jLtChPjBob9iNaeud9yCIl1Qw6Am
0hNIOT3LjJEkGNa45GNdJxXoKZf0RF/Nx0MTd3tLa9z9iy52Y1jiC5t/73611Aid
wbR4Mvs2fl1Ys3R3tRACgQQ7kpU2Uu1txnRfd9nkkakujPFTIcY6HV2pAk2frvHe
2a0lk8NLoX322jtgB0XQZy1mZL9fL7gnwxOLj7dJvBl+NKmV2bpxhWZwAjFoeWvo
cDPwIhABQ+omaH/jY5VLeQst1i5dSYQwfu9mYLdOKGKmxD32Ua+YmF3kMNz5TKwH
SLEMn9fSclcfcslYHdVSV13P+ABLsYVEclVGujAki6kVAnirKdVlO97s3jL5qhBH
XCIypXOEQgrNyDbXTL6u5YNjP/o72FDwPN7+nzzsQS89hqAduql/SpOHNo67VaNm
yxl+wQdC16hZu0iA2UUW/6kUMphv2axLxUQy5Lnahbqz+TvP5kTzpUrzA0Z1ppm+
B6Rl64zP2KT8PTkI1RjhZrd+98BEj5tNXg0EUi3mPJya8RkS7WaSuyDImq6gJn0J
72qK6ech/C2OLBfE81eKyB5x8lWGw/skW6sZVzDR6ZOFSqQE+g5D+LFwGX4F/qSE
/DFoSE8KRN2taCzJnGb4TA9KuDx8X5KmMwRpGK6TkCw5uU8xMkS60gShZjqLoPbP
BhH0eBU+Bdhj+/6B0L7jMjfaSjsPx9A2GBVP1xP66hIlihvSpriY5uPb/w37m8Jc
nLEZ4KJqGj384CVtKwDFjtK5rNyzzV/MIZDtrJL3mxXMXGu41v6HjluFsrso7bv9
LAWT86X1EDIou5gG0wBkhwAn4OiA1F/Zv7rBxwOaGVAQAieDcKQtdqyfG897xaYi
PYWboXH1rGHZLXzwQ7wHZNmjhEi9UqHyGFB23ZQgYjApCpZ/4v0s81aQBW3+6yJA
k7AuoT9tLa5FdXKEe98uSMMemVHu8nuoNz5TxeyfxwZnLGANbAHXILwTjo/ixvN5
rMN7ZFjAxU75gR0DZHzRmHUGsCNodhQDwBf/6QGW/zC3/nvqaQ+NDFi7ItRTzyRg
OPpI3wVVYxHa5PNF9LGTgFNmBVYAc0UxFHpFkeU5ylnIzGkR/+qiA+k/gqX7AkEY
NEL9gyEbMw0bPsnYGl8ho5n/haD/VnbL3lkV4f+Puus7PoRHmBCGQA9aDg4WuZXL
bA5BPoATY2m8VlwhMWtwf9TlLqxLTpC2WLl3CMiiq2B052SDcCSdKoWA0DNOUVnz
+JjR4IsCqSt6yrTn2mn0gZAx0rGKy/N/1mqPfXQ9JL0hEdCm3yxoonw/Th4dJ9bd
fa2CKZE8H4Rxezu5FQNFDBQ1JqDDkVIvMLi83VqOg95yw3g/rurF1Dh38a57eJwz
zJHvyio6yEBl4N+PG8i3Qa/TcIS0lDV3wZsNmA7L1NGBoOSAH/N0pO3J3/81yBSc
vQ9Zf0rHPJhgDL2fGcVwNPeqoreZbEgAcsV1sgk9eWNeq6/jmLrZN6nEKDD6OVJt
FNPPo9SdeVE6ubzLW+UbSgsJvS9A+9Vaqe+NIFwLl+5XO2M9hCjOSMA4lgxBH5xK
06GyQHPM0JXiIErvM5NSQQjSGvfpcH/ugtJo45wMkluanVp+LRafejv3Kkuzh3QU
fqkvlKnlfYcF1nm0incfN7D/KPvUwLtfUSERlvEEZ8i8nNQqDU8YNe7sB9PEVRL7
7cJtlYcCEgUua57xy/3DiIxIKosvhjfd2jYApki/Rr1caabddT6bv1ieB92FELEQ
q9rzeU90XZ262LHLFJo+2cLofN1YZgZtJ2Yu4wuPSEwZ3o3xriOT8ci0diqDErEc
AeuE/WeixF4bcmoHzDLJs0EIAkMaFkRWfdxSTdlG6OXiV8sIHsat90SwkR9OMXzW
vUO/vWHIysakUTihInY5vqNzRYweIqF8N2YDaO/QzP48k3TkfYEOni5VRHeiaNC1
K1btAPmcmSV8CyCgA7WLcMa4aRUAeRGWyjZmpY0HoVGW03ADyRlJVVYVyvMH4JX8
hbJWeFzbQThJnX0C7qM1veEZo4H/8GxpNr9x5fFAebiiLGSsqbfXkkh0jlf82nhd
wB0aPCJ4X84qiZ2EoJbBz+usDILWvUa+pE9UzqGLRUrqjNKCgEbkd9pukQzowV9H
ej/bWAuBPzagMNUFiQPTRiIbMjlHECaf5559HUYhpPATv1hOQUyzzSVrzzp2ChcB
9SW+Nr2AMziQCZ3lGMK4xq4eZnx/lVq7IJiBBp0vlE+2yQ9Pob/YevNf0CMp21Qx
v/WXiVXNrD8PWvVdv0SWqvVjJ7WptgXRD9JYpq7QqM5qswkp6uvYnjwDXCngj+l5
UVCaQYVzVfFIk7av8/piivSCS6Bx6EjB+ShZwv7HhbYAl9oQvU/TBlUwwsXDV7N1
GBN8E6sIqpNJcac0q913BzCKbuxJnMTKAvH9kK3sIicfYcGaTX93Yrj0DxPdDcJM
JhfNVSvmD5XlJ3iNCpAbDKFdUU+I9gnNCU2vGgQqJMxOYlVdrFds+JAgpJwyQ0h7
5XDTXEaRz8PT2ZYVBpWt3MCqXS/7lZuaQs4s+8wMw8oc6QyskWiaqrOSg5rzMXjL
xgvEb9hsb7iSMwJ66/ZVvoFLHMyRztCp4yp1QXbTx0ESFYGBgvHTB+b2RBHcJ7/B
5K9qCd4wW+jSIO8AhwkRJ5gtEkvQRsJzcqJ/TRTr7Ex8Lfm3KUwg9HkXjCX3Lr4B
vp/PeZ0Yp2aOk6z/p25dW6aH2m6cq2MeY7F/u22zRMEteC9Tdvr0CTo76WqHZ7Og
6RKWYq54Xkgzs5vPq2m7Xykg5c2GC7IB/Fd5MtLXb0lmlYd0/27h4/ybfvjZSUQ8
aQcFz8UrY3JUJxhWkWfAhtSsGUr+2s/K35qhoODTuq6JQRDJ+x7+qfG5mSaFoAiW
pV9m3RcrAqxFTQIseUNiUYVEAHvOCczcjg9vKN6YYEi/XppErcvQPYWHYKXcmGnb
v2Bk07HkqcCcSn5fbydK6bAgB8/iwOgWD8hoDC7xTDLIojjvtqd2rv9S9wMABYXM
KfF7I+fBaG2lH3+7eJVLRbmIWgxJB37S4rGuZcE8zIvoib+fTr1JeRkSNIddZNBS
/xS7EDGWoy6rC/eXZJbklwyJKBHmThfDM5TrqU/VXmI07lZBfTHJTC027fqLF6WC
32/a/zbJM2RpOny8ixL3aqnCJmRlHi3azkfcv0w6BvAtYbQcQRnmkR9LRjyr341I
8fk/pZUXlbGqzBUXDsTVa8YuiVrrwuALvoiiIp+4T88M5In0hmOBUvZ0k7s5I810
XBz/ld0eJqoume4CyrIrjA/z2RtnJ7TNsTN9eNJKjukXrLq98qAe1GwDQHibe6I7
37AZY779N2ZdmPaMFHNYCWfVWedjelis3yZ+kkLDBYIx06sKX/svaxQ8MLcTBRRj
vvMEx3BWEmgo3gcAr0olkFhEblj9uhn0tCR+d4A3OTKYytZCgUWgYDnBQ62yboku
JLNGHJxLcVOrb3NU3r7TuACEs9kjqWWu6QK1Fb6l3H5HPi/uekRmp+YyWHkpl4HU
tcWgrdAUruHiTtvWwajEsYJQjKo0y0qYwljXzTrPiH4IWIwxT5iwbVQlT1SkP1ns
AYaxyP3sTuj1Sh2J+YDvGyyKog5C12B0mS+kvdeKmO6d+9rKHNDaQL8uXCBVKui3
wq0IVjwcYui+q//BDkq7IOeOwZzmSfrprRGlLBApMs+9TUuMPs1lFv7SnJO/bVwI
//P71/bgTle9Vk85DnUzAum+txqYU24hxOAgtsGx830hZm3WBj4hbF+6i1I7uce3
yLvgL+9KmbYTqRyQehBKH+UROMyS5SxMYus7cJmuVBhS1oknzbhStLvi78o5eAq8
MhCvvVrUavVP78FGfudL/j6isq4Ppu1+fXtPWFVkfOIwZvGIknFYdBEGtAaZJ0DI
XJMyiUpLUTB19/Q6YaAdlaL1bDNKmrpAiRaUvEJGT4DSclkgS+GB4LWo6Nqk6N+G
Igg/0gK13eO5AOza7zgARyyWS4xBi/DzgouBvJ7uJzPl49ZZt7hURHxXQu7ys4Yh
zXpGh+Flm+hQXIyonDu6MwcfZgdYWNP+eU1EoXnGFE8TyCa/SA0XYKrv1Zwu5raf
nncemYWtR3R3s5Dcznyt9qX3D9Sk/fU92iXqikrkFHLlTCbBvHObCp45sHsHkoJc
qvfba6M60Jtmv62E8fEaV3HNvf4HPpn4jKk20bL+OfXuQdpU8eZq8WMumqDUqt34
3sdQ1wEOWERivLnRJ2WeNV4bSm7dG3Lj3w1f3yPybP9NTOLkG5rtYHPbXPdSkA9M
hBasobuDFR8OCA4kYdu9yxjoICPF3/27+Y0cWtIgrWmvpSafvozMry0vxvz3Pf9K
+uoZO8xz4QvZ1xd4DzmxDI6yD3IiTlwJbe81rF7Gd3Fnt6JQC1hijhh2liqv8mfb
qlxuBzHmf7HjmkvPicYFyusEpv1lOWxYLdrO44N/rSEY2TTSTqrEkxej5olqXFRz
Su0LDkF+FcB9IvuHVKn4/X8qtzVXgX/q8WaMsLA6V8hB6IuZVg0gHW+tHrGibaCM
JzKHkW2gd8E6bWgyNO/OVCthkCVes83Pit07+QPNOtDtAP8n++SEqqwOhk7vgx7s
EpUIjYFa6w4m+sXx5TDLG1CCnFrGYDJ7KQiHp5pqbknyrWZxgUVCoPCqwl8r1stJ
1rAhVj8bnKKhz8ushC9iVG4psbvuD+ifkS83E8gdzt+zDbZw/7u9oV5xGofv39Av
dBuJmGYbOJcbwCJrKl6T0dWhTQqM1muGnlnf3i7f30elcdKFZ6kxGOOMfu4Bi9Nn
4XEuqgHXa+ovnNeQ9hudUVCOYBaCH84Eps4yFKV3JZTEIsW87CgLPufvLpZswcwY
rawrxGYA/G11uV/zqNWwrevsvjg2S8ssFhhodD8TR6t4OjfedSkewaTgSFiSW8qZ
bVmmuFANQ+BL8MIdFz/4miF7JAEVcUNsxiZuslpuTBke5jmaEHx8elOMAjB2uLEC
XPwZYzgGmmYhNActq/lzEeaLBgyEENewmfQ5eIKjyFLCc3Z5SBrDJGVc4Prq0sdB
FfpiiD3kYQ5K4WsAhRFUc7DP2RhvOlVhcDe0gLEA36s41i5SZm4ln+lpH71x7KBw
t8jZR/DPpkeVgqma0GYI1EL70wSAcZWn8U/XgDM3YWTElvEfzGdsXtR1o/rP7pBq
/phSz3OFeyGmQSC9+5chBq/SaLZ523C01qXtLltQDh0OHm5JRLiDIZy5ktgqNXM8
zHzKbmprSEHycQDy4VWHbneMipf8U9gDUCwXkzUE0Cn27a4rTsw3spxHD7fsKybX
p2ns9keL+e9No5fGzq5mo//9BkAl9/6lGse9VYV206gBuSsRZMhkvhkGe8bUZd8H
GEcux3GRMVQkDj+EP3nfuQRi8HYjQAbGanxyW27WYcn36uXzUCTP4r8d+7byH/X7
Hi+0kbtdiiTvZ7YNWsaYZBknwNOoYe2jOjBKz0Ya3eL9YzkmQg5ieVQENI2LZzk9
xxS0h3taaC/cUkfS4z/uHOaLZKlbk+hLSh8lUOqHNwCRRB5S+pWob24wmJojT/uU
1B7kYrkxNunqVk+L9BOFvs6l9yYo2jzqalJFxgGNVGQGk7lIBKFq+9RNhlKRzqkG
H82Wbt027Ct8EpUmyJ9KAgaaRZ4Iin5yFROLEMdyG9yDrIFD1KCHgQsVhdK1k88E
vOewBQbKbyGc7O3Bo12YMhdpnF+4rBhYZ0oZQmAEe1wDqb+YAEAlxkyXJ24iN4Il
3vAdHRU3GAHCBR5gO9INNQT5XvhMK4u8kudOcx83d3IzimPXe/0m9ZfalljvRrOZ
jXjZaY39leNz0kV3+XApozjCx3+OxZPkTm0oqnNpOKWs35GT7qZRJ8hfvcxXHHf/
uZxbwk08WSuFx/mR0rurb0KRWUVXfJmXzzKCPdatAXnRlOtOuk2ObsXfZ6YQUzxk
HchK1sBi+jLCqoLSjorEgNUGwnXaFWi9y6L64ZJVD6ZOEOgGXKcBeBRUTcwnYMvF
Mv1GjO5yRqAixkgUizs8nBCN6cE/7IwqFBl4hMcn6O+e4D3mqAuVpJoQ1jN9HBS3
OYNxaWKzsqykhiP0ZcmgodF+vTElqk/nJHxHOpcJgjZww0dFZ93cLUZsDpE6+LZ/
757dGAuPHFc7H16C9fkbLd/URw7THltPYgyQ7zdhjqACComEi5FhzZjA9TmVm0a7
r2eqNgjbCFmPahNQS/KsGNHdSVLCNsnpKw9GVxDvTxw7inUSWQSHeXR46hdRt4Rh
fVT4UUvKQmNV09eg/Rb+rHwCzhUsaf+n7OLmo7A9QFR1EcpsCGhDaNy8nb44mCc9
Q0bndi9Ab1+qu4OAyZlgmJ8vOGLNyNTWvLpf3DNklgfZi3F/3eAoKQR2HB2OC3Vn
2XswEJBc6Nmmg95gMfkJr/AnXX9TItSt64JTOIolyCMB525AEABzyqfDrFWYvIrQ
eSNFcNmOPoo2vds7DX/qDrwmI8uHi3phE1OwGO1qSuLte79/8SejflI6E+g4v/e4
ONTlxEtSFNhMKwi4pvS3TFfxB9wzIn7rBz3s4+6DKw86SsSF5/fHkbel6IFA6ozh
50+tLY/O3GKyVlxHQ2OEY5i9jW48qate/Sb/DC6Ubq8b+qsQpDKft4UGYC2HwTcC
jbHs5PVOQIPnZBRuJkQrL+oHxQ/W4ncb9YG+/RnDxyj7+t5DrA5RaJqluFxaGwRG
FlhFTnWvfPmdzI1QmarRhbiTwz8o5mXrWSBGKUvJZLI1J+OZf6ct4kwEFbNj0xEf
E1mt0TuD9Wms13d96jzKL4Q5fvVB0kEk9Mtew8VEOAUjjDbZcxIlihSAfhofXzg5
goqFCll6PMp6vLWvU559NjA/XBBtJKHhQpGirX1NE4m4rLZL2UPTS5+3Bp3qLcxY
5JV5W8KT9RW2TfZGqVTPvrabGtePvf7x6EKt+A8TfMkfQatqG8ZIvdyK0TTwArKa
AE/BEfJQbSyuUCx1q+k9Ng3Fd1K74scoGieG8AuAcZGY6SntrCCCpc3o05XpOSUS
J6ljVdxE7j+MShYxUbrkA6RDNfkuTiSDJB8i/iyg60vmjc45zeTDAe9aogb9Pxvk
gRWHCUDDgo+JmRugu5GtZvVzgystuZfCeEoJUdeSFBbGiT13TRGyE2RNskh68zCK
anoDt3B8cfEu8KwIbSzHAgEIvxAPVS2t/tPrvmXDlZXk/QoOW/qj1m8xKPyvIy+B
u765yGTT6D4Ca9/AWhBgBjpyeZg9Yd2NfHeCcdqn2cnTgpJccxSCBKXlaKnGY/4W
fZ81tHPwJzAURutlscdd9rTjlxEwHEjOhbN0Rg9LpnmtkI8uIfx0Z5N50IkLbwGI
rnmDoq7f/ma00QPw0/E6TA1EKLMe3uUuqGYOaGSsWfbx3lhjAwNjE9NWgfTCGaWD
2Pz63Ork/Taq+dsmKRkrRk0WMmxjxafbZ3gG0f+iCxQyM3rMegnCfxWyLCYRlRnA
y8UQ1r6b3MEWp+rIbSlcpUuWVNloE830Lz60RBV6GR2MLNBgn3TYqAbGX4KI/80v
MW5hepoew/hYxw8LIKkOtn+w8nPQIoVhycQyFnW84mPth0WomjnxBsq/MPlI2E0o
nyafP8IAzl4U80YVJ7JQ0pS3QgSZlFCnpiv3V0qfwIlUZsEo+mMblfXmyuNUDi+b
uL9TS7g31TbuC8dG7ux93ujHaVD9Q9I5PR392LvZsllM9CBQ7AV5BNIaMJOkZR7k
Gp0mceOwf626fZ1R0ifSdI9WCxpxrOwBVFbT4IItENwC3etCUQWg5/dDvUKkjUJ2
ZBaVdk3+8JqZKKPRO4O2zkijIvh0DqOABFCl42XxVdUJlssEKxiqVpn0vNvXTU2y
9TyBNu58Z3YfLdeDuRrWzbEcbrs54dMEoMdt1l2mNQ5NVP5pxm1G1OfIWHJffySp
/BtHqHQyxA+dxUD66Rg8q7FIJC0+Pj5DKntPtFv61d3nVyvAm+IQRUNp1ynnW76U
risxhC+aj+FnkhIRTYv5spzAiFOP8uz7nn5yb711TkOOpn2KBu2NBCMia4pJb/4L
YIAqK8LAH2BOZW5xKuc3lT6AcxjgNeKNOizM/wkbyiNRqfc1TqzOhFyXEXGg5KBq
M4ooM9k3X8gpVKpQ5lX+HJvltCR3reipWnrTv/ikhDYni5n9et42AllFjbJrLBR0
Kg46jsCMOPoQiWlHeMcDyE0kE+GC5erLsBTu3bH/iUFwxYbyAYXZu91Szv3E1GzG
nYJKW5umhSf06NlpxuECxLNJTnRefmdBAtVQLcPaOMTlfOxaeymQlHsTUfJftodZ
eHIVrIH7NyFZx21vra2j3VyaxjSddYkQRBk4MxJftDIIwc9OpevTvPMXUg8pr91H
4Npq/YgYiVUb51wVXy3wkm2wAD4XSjHDLSTGJghbqkqzoLvcrmzHFTZTNGsBo2Xf
mb/A/xVk0pO1CeRoKV4C4AYNsuPAXxreex0Qo//UxPS5Cg230o+TcIRRnLuNX6Uv
70owxJhI99URzpFTv3ehbhYwh4IB0jmodGLsbva5kIltmU5xUJA8Z+YCs8343PHH
PFhunia1MsQDxQAHVqkIStoWGRqkkDc/hf7xg7LXHbH98NA2p2CMNnbrFuOjDOyY
y7bukOo+l/iFF7DeFk3Ia1y5VGKqGUP6eQZL9iHJVLtkFPsGEIt4AFDO1XU9spiu
lKcBcAcKbGp6SV9l0OHKQn72yZ6ueFLVgTYwBPonfoA9kue/dL8buYISuzFV0I/U
le8S/q5jsJ0vWB2dRh+ySJ1ALBg7Kx9HRqOgxekXHVeHRLeEx+KSkv9hpid18uMg
wdMnH972lHs0jMew5rQ/RROBVqGPAOlFMaigJgGK2uKfJ3eJDwqL9xzreDlR/EoQ
YTDw7Ep3A09feL461bKkxog+JRKlTgNRDTv8JzdaykopDnk9qa8kvUkroAOlhuPp
KtmLfHZq+phfN2U7Jsap2oGByBtZrfoNuGC3q1NfKgftOgJOd5iwnj8geS4HLCaj
L5rbkWw/n2Bi2ef4tWwa98u4R29pTP6vW0wi9W1QYCgPdIi08S8Y22UpOXIwOSXx
ggw+0RGd3y8cvCn4ga7Qm3IpQWw5uzHKyqHUpKAoAr5ORQglVPwBjfaie+yFv2eI
c5pFptbEOyrulALqgXgsPS5B4dUBgcSqmarcbUy3BWqLXbT7mQGRwVNDOvYjvEhl
hluzYPILJYghEUtr5orupzZ1/HctAKHkqajxMMxNAUsJlLYnCMbk2gVzMXPo1kI7
BuevFs/uqRb7sOfGDrk0bAC069G103/3dbhPibDEDToFHE8xluNU/yiSIY+wUdQC
9pghUT6UjqX/+kRFLImXmy1tFGOmfODb+/UbfX1Sg24qwZ4pqjXGydnWpYDzDB8O
q9ve1wHQN6vtbNGyarIcHH/j+BmISp+BHpsgKTp3c6rmbQV7/XqXNrH3UgU3NqKu
BgJHTVyhcaSDk/LhL6xr5mJu9lT9RC4+3fOZDz/Z8j43ka86UoiyORisOEQO9HmX
nMmJyJ2R5PMDGqqIzZnEGKehpF4Szgkj6vzHPT1O7sfWVi7rbXfBgwG5B1fjsG+w
2WgUD4a0h/gMslMynuefLG6SIMp6V026kLlwMl0SnK0CB1jOJP/SeCRBkQSZT2hr
ytuRnZi76Sm/vZ0+n7Ny0/XELQLY3t+vCk9t/g0Ik3ntzQRRAdx5D4ICce8Ggve0
tSCy/rK5yFSP3KXOG85lmZ2visIqiyokYCtW4/po5Nm12dkFDWhOUCgZ1F9MqfPR
xBbARTSlYwg45Nx+DQoHhtqurGZSEH80Ec1vpy3bDXSslmnNlSOM0EEPTIkb/J4i
/p9Jr1p3V4IewKQRMfNhBjbAIshj/jEIyaQZR/BzEhR6WiyPhaB0t2iN+dmGlVhT
V31ihpm1LamkK3pXIL0kj2+5FtugP3Jou//4PuXbQMtBeKgwIbBsRYX0sq5TAXbS
MnmhofQ2hrQBZIWjqgPZUUJkxDtw4f3GiAPKF3lBS2rD5M8IUWxfERhF4g1wr1bG
r0UGqI6lpSsjSXv0MoqkJnXdtuaNin3QSrvLz5YEO2MRm9K8CzDDJk8Ze2ASzdoS
8KM3mX7cPArstk6D+KmNM0KZIzEVf0LrauE9Az1pL+8xjIk+Gn34lUcB2t/sXwym
ewG9JyNPG5vmx2FKK+n8whsmuQQ8jOOv6AmCKvlJDNAhhu/USMdmNheUSF3B4/vp
yYJ5JDBhSuSnHQf7oqchlu7hC4CJCTkkI3VXL92QhOeWkJUGewBrjgokp3MKi9VG
LuY0gpvvjn/PyTxf0JXT5JEx4LtqbcMNSbBJjU2ohec5GY+rjWejysfNh7+RgoPT
CC4Il+88nRzeXfGTeuQWV26Zt4P0Ai0a1ZJBk25IhDxM49f/fkpvoEKKmrL5IhU6
i59xX+D7w6sJWyU8FGxVSck8EG6QNqk0xK4BM241faYziiZnlJBEFqnGLfjyfTax
eDY0shNxi/yIXoaL4IYnF1X9/DD7nn2Rh7Fjix6ZpRJ46BiHwhOoIb522nCzTz8R
cVIL34fz2sQIvozfcxShCY6qv1XJFIIdTAkwO3zF+pJn9XuCmjGkksAV9a0B7yzw
c7xLTRsoqcz2UdnG5s9+PeDP+n6CedIgv34S3ioVK67r7RXChs3LhCArBnH348Mm
wncpNSe5PGHFGfDtF4dMbY1bPR8R1p8t0jpysZT0Y2scwaypgdAvgKbhRiPSscDC
sERoICx2ZuMc9LM8N5FTV41vbK7sousc0UfLlvkiiFgsfvWPxPcHIl4QgbTJxWwt
SiaiSbwC86AYPLQBGcwME+SMv/t0JfdClRgSOgO0VbpwyvBZPNU7f7njZIE8LsXF
k/EibcIWYgBRUbXwvKfWb9pWYU4YoJICZBvBvZmsXfNEqaB3m37R+KK99wIzzjCJ
+IMMpvAmIQ3uGx8JmdHlN24P5veEoxMD7OH4shZigElhjEt75Zr0UugoLPfxMciz
7aDvFwfb/xXlTUzfKVxZY3UPzWBdX8u56U3aIfjiB+VADaQRMz5LYrOFNmrgwfzY
689ehHtdsrWiuLlgqXrz5Ztq4y543wFY4xoZVZ6KHt9qjdyIEXOCiaJU0FtrB4rf
4iDOm/phrU0YqQELQX6uq/b1jIxqLoVQhD693UtaMtw7pPUrbB0F6iGYjcSx8pqs
0lcYy1pNsP4vrNOsyfORWnDkSuJCdcKmzibMpZvO94MYySVtZ7guj5xgVyu2vEu+
1IlrlS0VswcU9iMPXYqkvnU/9lKX/392+zz12gMLHEyJGMkMJrRws2GR17PdE2ie
2y+ZmVVNkO843y+iJ7rLNyT5CBZRrRGPBH6mGqmpOiqBaa+tkpf9KN9VpVlVTLCN
w2lgO/+5r+ZO9ptJjysasX2FDBqC6FJfX3KapXUtST+PPx6krEps3Juf5NHaSNcs
1J1NPidNx4ZydqnG5lMhbKuDxPbNjpeJFGwb20s0xOqFTQsrmlOqW78YgWRa5OhG
XGFymKclJAD2+En7r72uJjlqe/oA9+W08z04GMX/BHm4xhG7xSqQThns/Z9CVoEd
9bwvO+Uhwi7Fv+4wLGGw0UYpTVzE+SmHo5qk3oSWvawqK137oyM6PgvxD6gLbvuK
1ueOWmSs+sWvTuasZufUQtP3iWEg0iGMZFLafDi/6ZQxJozsOejaAuCE7YXvtihz
NAkldhp7XDOuWAqRqd9hiivxsd7XBcuelGhKgjr1BqQRwI781UvwG9BpxXsj7tq2
XQClUncYusibD1IGI2XbdJ6Z/a5tj3Sq49s2XvX9jjxRmqYPQfLA+yjGlTxBcMsR
o1zaaC4brsIwH2nPO6WdyyMDGP9M1DZ9bIYcPNjyAwSguQEM5Zm5rNOIkHh5iuil
tj9bGeRT/2eSzR1uPCZgRfUY80gHxg/W5o9ODk94HbOW5vVA/C5R6WxVz4Tc24cS
zFbg0cmT01AqYDJflY2D+ANg1NbACELKbJdQ6kbQTS09Nc9ezDFPLrOhfImA/AO4
PPR8MmNAEBIcEBqlt1R7litI1EHDWkN1IQV/FdTDB5mhSq2rrn1QTBBV9KRIgYyf
mxPjRbyF5zuype39LWw8BH2k83k4g/CgW70m3iPawmURvf5D0+wt2MBM+maaNS6m
ZV6eMn3Jdc3ccvyAIhVvuiXzliRaIqIoLf155TPsV8O+NjaKPEZaGDra3GGRUwwi
cIAqKba5f0FXMlICDjcoG9MHrzNQ3aQeRW59t4Lvsz8t7mAwOXTjHscAKU7se3/0
ZFapgX4Ej5xupvc56fy+osSsrWqXLfDw+FqpFhxYW1oAwo95DH3TlZ0V0x8X8jEB
1QwAAhURQZXLu6XbTcvMtgOLzRqIbKPFYERcq9eh9iMSiQcrveWTF7lelTt5ao9g
cqfXM/dP4EylWWGJqlaDEQN58DgdSmuYWgAmQWp8nuKXA1ao/I7GRyBPlH1Do1ip
Sz3CJKvWYckdFF3J2OdeXgo+KP/L/CPFWmsAwxsZIylhVaOMfPXk3eAz1VhyLeCP
pTjvGRerb/Xx/cVnBTz5e0+WS0ec/FO3N3acYZefkP72P6TUT5pFEGRYYbk7FZ4q
ZcBOAc9kOZjamgfT4LBnEyVq2U96Y0+DFtmp6zmGX3XxjazCkt503YO/lbA9jUPM
zJ0lezLLqMLpSc27MLEmKLyH7KruLh56HtBFFHSuHnAGhsZ+VsPQlaN34IJClvDn
iLjAKF7khpLQhn0AWe6MTLrp7hax/zSG++lpsoOAMdGDsTHflYWa7xl0B4Bo2MUx
1HQWnPYhREYzKhV4CR4XZcPKO8jj62i1sgEjnoVQvwVF1Y/lwmew8ck9bugzU30r
BbKM3y6UrMnPsbAUhYm3nRIlBjFLB8BZAe32PG89IlqHkzOF493kqZxWWxsSnTr5
uFGPHZXnZyJRjfRANKEyDSJvVWEM1a2dH/LqD0BW2WU+4ZwDy7LswriBaPte5Zn/
XkYrRN9oHYnH22w10xhtIryYhePuZg1a6QEbiwafwmlW/7BIv/LyJoI62R4tqOM5
vh5K4wwD6euDGTIsYGxLajIrN4pMKx/QkGm7HLJyFZmbntpYx30elG4mZKMLgq6i
NRrFk/XPf46yM0Q4Vd9org6TF/Mk5mhIzPnb6zmlkrwsn1ig/BzZ6H0IrWR3QHSN
+DiBtQUQBkDdyo/Jdud/vFKxFBKd0aricbSMVVKPBD1EYw2tCCKrcnY4M2bONaUi
1rboEclQwT4rBBgD13d9V8u/wBxkiGPeX23PyGpGm0NXZM1A+bwLLDsyQKP5lNYk
sTZr1LX61aX2PKAi4CsJicB5emWhNZRkIT1xf66aqXlQutlPGy8CVCfETGuLcm11
wvxY6AGUOFnK3bnK7/JlvuY7PMHlo1pJ6waxrJoBJOfwpwhH3voW43hSS8yHQFes
BS8AM9EnpA7Oips4dUZLOgtEn7Y0bVBLNlDKzk+h9HpC8fWf+AKh6wNF61RRviN0
QaKb31UNcwMotoXGEOnzIh/aDPoRQZ5L6Ixbk9KGf9Ek9vg4ztLc7cBar9rjOLsa
l5ITinX9yTZuGZ/jpSd7n7RWXx+oX7hFGjHEO5N+fcbOLcyjEaXocyg12t3vjAIZ
n80Zi7wTnTm6Uc1Pp863zqPcHW2YKPoEKDNS0jphaG1bmNrpS+/9iw7DjevMuEiR
6AOHfPSdnavDbkDxXLIgdesbPE2PLqUx4JFKGvwJc1yTjrRBCk+R4puUlgP3Z3Qs
f2V/tsod06R5Ai29TJ3jJ+V0A8+5uVWp7MD99T7Ipyt3+58gj+7QlQvfKSDHWzx9
yErNp/JBOrIeb9BLyp4r6rKp/WNu19ze6rQ2LvBtU1VGaZzUVz9xH5ECT5Ir0Aif
HtRxjZwBFbn5C/i8KZRiMHDLaUnPA1OCOy+/hrVvehorykZjrAnl6FYIOGRKzc2F
7pJjQAuQVUMg0N2LLm59AWMKxD0Jb6zmVeBxwns4QSrtpbE32Z1gHsHHMqHcHb3x
aiS/G7nH/3aIW1qNfTd9vcL3JPLTM/m0zNholSBidE7JIkPM4w6BwbB3/5ef0LU3
Jyd3Jm5r9qJJQGrkm0Spb7FUvW2pQyQhHeFgAzEnaDAnYtyxbg8b1QlUECD0pgKV
R0sYlSJdghYiZtuWWUazWSSgniJ9zAq/OFkqG30ZYhas0WvWn5e8kJWy2zW0Vrbi
+TOK8OT1KNKH0gcT9F03g60KBIOV/PO45XQFdWaDxyM9iInW602BNvHMkBcbPjqL
tiq6CPaQLJWxklTKm2QAQD/Kh/645kxMMGDnJMom6ORnE3/WjBDwylVN+iG4UWf1
Slyqi2yMP7H4cmNctk+41p5kZzYsrcADZbx4M+8XkMLVAaoi2ZKrPwjwpPaF+Dh8
m0hPQiYEAkiF5KhdQe7dbz1PXpFjKyAg/Ij9CiydfY46g0nwLkVgv6b1VJciSnwE
MMspGSD0kEf6m6GNJ5F7W1h57u2XK7EkTm637iyhoeI9/nZ1y1o0OhcvrD7DgGD0
sG/Abe0Bi5x7G/PuoMlZCUbC5F6l/5qNdX3oq06iJIxEEhz8KF0V+ktbUMDU8GzD
qefWvYfPu1SLLGY2AYi5jQ5JpCC/2iIA+fPgZRNyTVUrH28X+zItbnO3BEhKk0Xk
PNZGqkS3O4HmJI1x+jT1W7m3WtEXn4iZ2KcPy1QJKzQ+qqq1QXIT+peJkNc2e3E7
3wF1lD5EvItUft7TNx9AtCHyQN2pkL+Z2GIuWzTUAXHVrDcUm5CFW+BGTgoOgA5T
l58QAoaufob0ukigbvaK+haXw18Jk6ZPgbTmoGKWuUUFIWTFNv2+uD6ZFh3/6uXJ
QHhDT+wYBru66uGbiOx9fv8vmzmpgxGXpjePjugarK1BLaURK47FKKoUGzP+t29+
1fRX3Ws2vfIRD5E0JbSLMztGk01wjOiJ45nxCRmNh9k+E03Hc720+uZOOX+B6owL
CerWC/FSC7gPl1d3yi+RDBCWVRSnE7lNWjh+fLz26fjnKzrMzZnE1KPMUFFKd8Pe
EmmeDuR6L5UHyuEq7QjlY6B1vtEXGdLrQ//rDsJSTxAY6x83VA2Kbkp49vg7Ns+x
Jos5O6jheUzYuk7+K/Bj6pyQJPZCvtZczUPImDeCcxyi/lbAl9KV/ukTvUI/UmVf
MW3qPWEcKrV84EN4KCj0Mm4a0KQ5Cdu+iWK89xH2DFzJAGqWNvI1neVz6mKGz6VL
jtVxs1/bf90BweNhr7uUZVp4a3VX9oHDtX832Y6zCoS99/DZDP11ns99YSKNEMEu
L7BcBiRs07BFWs2tab+zFwlu018QRlegBJfUeTd/1kf+2ytcf+qOjOgOsywyifPH
beEn3EC68wvPJpAavCX2xfs1L4lrGNOmE1ri2N7og4dZmj+06rlcuJ8w6BXAviUG
Qnl1b0fHGtRXCr6LnXI1Ox/+yQX2kf95aOiSJBkfvygALZ+rY0rnTRCOmuGPhC81
x3LFLnZlckcxuEqca83HOKTANj0NY6/1JgLAVDgWFLw3Lc3YRpHhzSEzO2J5AljF
7mg9A5/fwo/ABS0WvWpuL2/TaOYKNjhbMtZvEnL80NXMnsbUrsSh/jhvIL6YA/gL
iPJ9vUoQOSrcN6QnFfmMIjy3sG1+2Jvrj7PF27gazt1vqvNqeQtSVK/SS5FS5O1s
ig9wikLYZjGsmfoAfQxsaPFF7L69DBJGwHdv1/6lWd7aRCC9SbMLMcUgOK0un6Ts
dZh1GJJJjUHo2vJ/Eyo/SbdJHB7fwhx0vJ1v8K69HFvSEaIA2G49GV6+1VPkSQM4
I9yHykT516V5QT/J42IgSxkl2Sk9x0T3dM86FJ0dY5INuuWjJn2HqR4BA7a3bJSc
yKaEfvhsKJNZbnf9tPdudg7vk8IzUTZeaI6reh39MMNFOOQYKywQzs9IVzhcyyql
FUijjBwB8uMd00ZOFIaggKvtVBtc5SQpfEMDUNjqAuoI4MiEPzaKkVX5BgnpHB1s
l9pznwLLnVwnLexE8rQ0gZWQ2I21AMkw2IFVRmrWPEZts24DcF705pW0jcdmS/Vj
CgmCfJSj/T0LzX4FIRhh8R1IDwvq48G5YBbsH9vjlo9E3U8c5WyIlwMxzKcP3Mpz
mcUcMGLWIikxQo5CcwLjpcWKtih4jJOlRDcMdW/drGPN7somHrhkxQV8WSVfcL0M
MSuKRXk/7Yt2/kUxtvOvQ/SeWPYO3vODMCQ0Bo2nMClVNFNgYSAk5sZbjHSgCCc/
/UAxyHaL1ITqmqcfelxqSqGimGlNknAvBx7VxvMze96NumBuDL95a4sYSzoKBzzW
vRZVk18sa/wyKkZwSVQQNaCZfon76sIvpvnb8iOsFcAcPiBJwZby8YIa5n+xNgek
laZrDsTaRd6NxZFgzCdi+4P5O/+byvLZ2YWHGr/dV/XmJ4Zc/Ak7M+bu9cCVMBwa
l0gNhX9ZHlhG9EcOswxBNp6Lv6eL+CNjbvdamia4sAU+Q53qoqErNwRWXJgyKpvT
b5V4rLVdyVFfum6wXN9Za4P2ni4kpUQcGklX7yr4mUPKmuBzB2RGMuGhDBJuYSgX
D7dN01jQuanWcQQShSHX31Mw0ncS+kw8mVL3xWvxyUqDj6OI09V6JmID7WPN3H0D
E/eXvIrph58bcB0kyBLyPvme3VpRKytNUrQsEI4bYFF1kpADIfz8oGUWzb1rBEQx
bQYLCvDuQKqvSkOQjabEAcDf4wUv4cFXT/lAcrYkCOYQU2cFquYZJGQjLQETj5Pe
zxnoVXyxCTmRvSx45sNxalyN3O4peqakIqFs/1CSJQIyzaK5C2SNzppfMwFEWpXA
/S9KiKXeEx57E3cJLQf04iSappZH/FrK0p4JTNAmI18wbSR3VbdcDqrIOTaoF5e3
e1Fjk7+WKo3nbcJmbXmGlXy4F44XvCP5/KL3uF32E7h4gG2IbCJWqWMh2egBC3Jr
OxSUeat902lUeMrUdOEucC/h0bNDnG4AEFqaLNX7kvVPMZx4bpfPmpoGE2Kmmbvo
iR4F3F+qnjTAOgDB/GYkx9FqOaPU+wL+OiGUctBIl3G6Z+XBDasCmid18XonRX3+
JHDopkZ9dAA2/OsSL7+XOF6gCf5iHIYvguRHzSgx7nTh+zuylkjWvcmdTZ1KPTyM
WyfHtpl77kRzyxMtwEDR6nb73+27ILSd2WGCdBV0i6IdoswWQey62zhdCQ2DWs1/
vT7EXXudaKg2onQOVQgYVp8hd7X4/mcI5mruCFFt3w8J8p9xgSZT8Gj18pFeQUCb
c2ET/hMKiTR6NGj66WmxMZgVVE7keUltPKuvBCsiRB6LWApEZunkqfULW0nKMhaM
RcAj5wm5GLqMq8I0J5vO2n7R7LC+KgR4YHlxply/zpQxlrMGXUDUeQECc2iM1AkP
HZ+5YmQpcln2mmqZThDE5aCXzIADq1wSTEnYyP5Lrg6zOpoM+sXcI9NcOLzqW1pX
VGYgrcrs7Se4duFnF4A285bZBAzggYmgJ4w5mmOXLXunBGxEP+w4pkcs+6UnX5to
E176PHsNccZHYY6PF73snoSlJ0t2UvO5CTG+BEbgsQpCghwWAjq8apBs50+RnYdb
nE3bL/MqX8US0+dUliEecc+JH9JIo+ZjCL68oLDqEMiOCD6yge+ewWoAk5YvSRbu
wbnRWavuSIhGi/PrAkGAVzAC0Nd3ZGw2qSBKgICet3jveT7Sq0G4F4LOklWMkWku
Q0aBPs5F931XVkY8LtPpOfeR57X+RdGOkN+j7msWdglq6SAkT/UX0zckQJF4HawC
8+7mW+E7Yhwh4SEwPUW4pQvvp7fwsWCxnpwq0bYT4MR+/FncPDT3GPBEN8LqW5Bu
Nu5R7tdXsA8QAs+UU8VowbYOPojrl/aQFKb13jSwt2jV9B4Ew98iE69oTS8XJLU4
kKQOc+wvStv3s2svfTKVUZ+Hm5H5s7sIcICxI2JFSc5AnhtW8uEFtQJ3y+Tfpu0K
Rfgay/iNgx0MmYS8/oJ0PQFB2PhBtaXBt1I0WmuON1P9tdNJrpxQgSMfxExODkcR
8Znn3QECg2TsVwGe1n8QUtB01lEzmdcgIY1egeKw18mXcQH0fR6hioRtqiWMW8hX
FXeXcuZuaqXQ3q9DIa365s9qr/6WEq5qLGuL1pKMyWQYPKcTpYj+xpG6a7lWvys7
ONtz+UhUZ4urM8Wota0TbM7cUAf9ZMta5kwYFp4fPQIuBAH6SwrsngvW84iYuq4o
VNJiTh0sG/wWURfXrnuMvFrVRI4uFgX6WJYKbGGqfvkHi2QlaDBOXdO7jhtXI7v1
SRD84o7klLuk8mxIfGe4BJ6xhE9BfW3Xsj1siWZEzdEDWKQERwdaNLm8xrlOExFy
BY2vvwGi58pEYz6xlN2pIOCXjiX7uspcYRlLNsmduM2qtKhXqVOoNYkzpB0YnXkc
cG3aIsOEnRhufofuAsScFsnc5w2muJhGMX5kmlZzV0S8KheaU2DMOqACxuHslmTe
dmoxR/eC6HkxkbWfsh4d1GBwvsa46E6U/zfnGaSv5ArQ0PreAhQ209IOJNLJChkD
lm6pNR9WVllxEXu9wMCwwKGU6+8KsswYUxcG4aMzmgTzt3hC1eD7O4lOX11K0FJM
A5wrrr6V/ZJKGE5CpaY/AbZTY7UPBOSDPYiPMahXcRe7AjKijbvvQRQJVO6C+Eti
WLy4Er3dQ8PWuYKIYz4x04AvCh8APW8x2jCoWFFcHkmiKwQRUVzduqgKAhI3mfDY
JveftB+e6J4qdZXp9jFYT//yjPR4eo5CRwbB3m02IChAGIcbDG08UGOkg3AdUYzf
EDB11xtW85ZT9UlWVd2eupd6dEDJ1PbNyrCqNTWXPsT0HU26t9gNM5qPqS8E4j1l
VJGkaKmdnowvoIR5JyMLj46u8FuNzWCzB47LcuEKoNz5ipnFbieMIxrIckQnQEYA
Hgzq2f+4X/Xf4ZWLB71/4w0b1hEhuIA1zy4uF11wKQJiVOqLqHqnuEzDngk3FNmX
x48NRmvRoorULw1ZhGcFrjfIg+z5fCj9VdHzcAac4TWknkkyQNqAw/u+uhtCgLsF
8Pn2XtrZTplBFRkA8dbEuOtYyRVVzYVVrZHre0frZFAbDdX/DAIdsnI/nugTcj1D
zBh+o9Ttjh4hPUiIRBOYKdfXVeR+0ZSGMG4chI+OGH26Vj+57eEpoSszGcKMxJxg
NAGBS97zQJLOztFZzM46J/lCQveLsk+ZwP5SClp/8dM/S4JZIIsEBF2UAhx9rxDh
+dogZvi3hfHlsNf2AUavbCrfT9LdItAzBaZulxDbxyKL1ioTnCBl6nZ3Yo7bTolx
gBlOucPeUfyptARB5TeLngae63V2+CZN3UTQw6QpHzx99qfl7gQWVUb1UVOFbqBI
N7dx7volbZL/22e7mZQteBlqnnNJ99EahWJo95svVY/6Xi0vFs2ttCOhE7VPtqoo
YMHjn/80WFbygZG0JVBExeBl4uoeQ7J7ZnvGRNjKVykf3mKdSD5qO5PaX3E8R7U6
7peqX/knYp11LsLnj2o9SfRGGKHKSVlTSKg7jJfoW1UXr5z+577ziE3PwCq4Ar/v
aZUCMBXwI7Zzi6Zgu8dtXjZoKMnm5W+ueWy+xgb4nVeVbNLq7yhp8HdxRrsJc8FB
XbxD9rdr2nrDZjezOpSVIntElEPx2o3DuPXjcQtIB7OuiiBg0tJFewiIKn1z3ZYU
xUbUq32rVlyWwbidVjlKZA1bkaj2QJqMpvXHF8EzIbEljuwalQxC1Hjpkb7BLx0e
caMDyZHg2NLsfyLZgZREfHsm18tbODW1GS/b38kuSqmRrQvVbt2kLZv1iHqh8+eX
EwUddxZB3VPNibfzgUt0FiU/oqAgVyPAUa7FfL8R0NkBPhWNsQBgchUdro5rTXuT
cGrEUVrWJIr2hwaT0d7ly+2xVei7x1gxHpwPBED3Bi6OygPFa5pjW3SZxtBT3HOS
y0vkNypaYSS/x4R070UyTVMJmI/6YQbx3bpgd4HKDRlQTPBNnMSkWY6mrgWvIgsg
aj9/n7rptgQJiQaoSWj9dbdgHuSuDCLYkNpqFYt8hHqmS3iqu3HIeqa18kRiHxG1
aaxZ3fbMlPqPh98+R9VyZqeOT+pGTBsFQo/KBhAGx4Ez5FAVm9cJgHl9kDUUpeMN
WZHG2utTa3yzc86Lh3AoA82dfPFxSrdFPjoo3n+c2n0cHMGyD/r0FnDSg/20sEaB
RXakDPBunzHLDZ/mU0P3yvM/+ZkjnPPZ30Udl0KCkP4973fl7XTT2A4RBYEnXr6o
oawR8MOA93KcXXoa7m9JkihR7TC95i71sHQVw6v5KYmXbw5+w2UgNBtjyZOlNOb+
vjQHm3Y02+Eir+jfzvyX5IqYynPNY+VMjSOK3frJvGIzY9g+dVYAT8x98EAtVL3d
kbG2Nf33Dl7p8OfAElISy5/4lME04a4qLrVwp5xhQEoNht/BLo8BzwlhnW8FrCzb
uGlSLkfLdkMpMtj70i3tUNXWSTUGGtooAhRb2QRUG5LZ7DC0OtxOdZ4UsLPwno46
yjuBKgLY6ymwJNMcyMlZrFiTfMmn5otby9tjd6+pcLh3kjAZh7586BklkzcFT+J5
+Rphh7VWX/ZC4vVD9uQJwU3vto50dW3jSCi3slcUQJm9IgYbxwhZl38yC3wGpbhH
49CiIqA+eIA6rv9PqQKJ0YwY9S04vuu+wRzoHUTKoks0S43RrSZ3LiWJ80gaFRnQ
/vLp2tn9bSAgw2ivmhuDB10sivGu/4kPqYyOCuA4nzcXedgiuC2iGa7eTJcIXUGf
vIQ2mQMnkoBFJa0S/3rpaDqDY4hIo4cVAqKb3q/VnoGENvbYsx0FeeTKBhZG+IMb
r6E2yCmXunmYWh93g4NsP2B+RnHhoDMWUN157ZFbDvARlyW3Hu0dxcZl/iW/G1Rp
zuGpOerSqouQtCy3qDdlrgpngne/jmKs1s55V63KyUbUiEoNdNs8Agx2RbK7BcCd
zlm1iYF+J5PLAWNL1hiYVjiLkteRDR4dD/i4cN42jdEXXkQbzzSGy/2ZocCZO6oy
4IgkytKusFjinvHhr1Opaq4uSC0QUyWmB0q4CNakxWFefCzuATUa0RL7sPJACTAk
Sui25d8q3sDlXme9FwUmlUIyQjbmd15/0iY1ks+RjjhmFammK40rLJtITk1nrDr4
CvZHmhN2K6k2qk6pyZlPTIRfZg7hhne9hc7iNGTqCdpoEw6ZLzX0Saxx+h7qGEgJ
qxn8KB/1ae0/y1BfN2RCfIImmZyBQwuosqyTOkp4Um00qmq0uItYw4ZJmk9uaRBT
UOzR4mOJaXoz/BkbiVh8hTexLpAYcFmdz4P0VMLhvuHTxz0ihLpgifJwYLZDIgqF
exGN49KAw1jwHt6JvSs1DoVRddjFHO426REWv/ZrMvsy41Xfj1MSvIT3ibkmiVLp
o0Lws6RQKhRG3QiDb+56MsmDKN6gixq7CySZIwsEFTYQF+O5aZ3srEy904pfkb23
bgkHhfS5+Ug2wHtknKdW8OzAcheIBcd8LiecXvQQk6MayTRgWTG/F/67GZ6wipl0
EF51uGgT0uvF1ViNTM0hiVi0MEn7WTpu+GqBCkjw0UDF3r3aq7YPbhj0BeRQjkGk
mOYeaJeQ+WyjmNt3wa9ul4o60u+oGW0KwrP7S/rzGZb9jz2RoMDH838MrL7SdfnS
9iFBJ8LrUwYUHtNHVxbj2sh6PXbNmRBsluRbDZhXInuR3IU2qscHlbvimcjp7/fR
GorXx058/rtnqOS0opEJgOAhd4bJNSA41ibIY9AnBkBJ98JkjGH9Nf2Lea4g94v+
8CpayQvahRKyRgCY3xOSowxd5kpHklikJrXR7OTHPvlWjnIfQJ9Ue2x5Whqka/0v
VBHqUZVGMl12yBRkTGc5bPWeYwDTYL02nsGfBwtXmL4moMJqq/JivG+9mk6nPnsu
ejtDEPLw9/oBxaJy447zZL/qTCTeeqRHTlrS5usK4s5/zz+gi2sXEt+c0SACjoTs
hCtPAfwXlM0QzuxrLqNC/gLugSUg965jt9GQcBI2hcQCEAcRaJLpMbsThqxG+gtq
yFa3wPpUHMduDkadyJ7stvMYqdP0hEtJS+jhb5HCE/Na1/u3k5oPGCVg65VaDLrz
IuWAxruD5NVJ3/J77bWo8/6CGMQ7YtSxb5dI3UGCwM7TcPsCzG3XKI8nySx6kGtc
A0jz+7aFxZ7b99HFdMKxprVPfG6YCBr8bdLyhvDjZKlRP43B9q7opkghA7DA3b3A
gx9M6ExfzVHl+9gkSejRX2e3XtOVsg/Rt6Ta/5/bg5xteH3aBLQPE0QLwRYJKYjf
JdIYxqEyd08prB6pJvkTPk4Dx7KyN7NpbEDWtPacUyMOnrpxgWM6rX6V+izik1QU
stOtB4at5ChOle/FJISaaKSFzyd8ONa/UPQXuVjts87uezr5jm39LLT3QWyrQrmz
euiS1p6F3QMLMgFmMWhQZ5VvWo2wR0cBQjgqP44uyYUAbegTLRuODysb+8OIxc0i
7JiuphVx/E1dAB57QIwdZUTpmDlOIfgxr/fx3NyiBOTWyHe/chZ2zGbiB2cwWdfp
7SufeUGlmA83u67I251uBL+ifsF0StqYpNZ5aIHfgGRLZ9SX628lUnBx9YmcKaH0
YhuiKJpVjE5eflEs4yWwNpL91GQhUQ/rSa70JcOzzQ4MW0KX7tr+HrjVVUtqTv9q
vQU6vsorvraB617ZWKCA1AMlQcax0H8vNQNnWYQITdyqIIit/4t1m+JZjacFfsGK
lGAgyQf8PIfN1X84pI/xl5miPeQmwbmt7cDmgfwIMBzSpV5uxPTRSAr2b8ReGHMG
8C7OqnGcWSv41YvlWJeZcbf69aGODBBWQCFBhYuO/UJFOqWisLiHAzx4RaKzzsy7
MUPzoFR1+UwV58QxtHvmxTkycVCzISqe9DHIjV4eHJ4m6zPYL94J9k7JV4aauO3U
x9JF7yhETPgQAF/hNWnWDvzJZq63v+ZIO+tg8/ix/gqF7dELRVUevOd696OTPx6u
gRo4WDY2kSMk/+89U0A7VDL9ZwfFpnzHSZ3XRoyd/x9HpQQYV5mPzv+LmqeZbto7
RKusD/C7w5KOp59I2puZDpDpGzGBy+hX3VknXsndAVyYq2RaA5oT9h8t/kuyjPEP
G5sG58LCAKP5oGuX5x9SNiF+gA+ng/nno5w6Y5+jZPR/Xv4vkXmFfkx02/5eYNH0
FYRf6A3akx4HXNlkaq5aXYT7tEjHXlsqe8vhqAgE6FbIqtkXYJi/m01JYymuETrD
FwXB/Ck4WF16v0TDStDATy1j7+iP/DV4xjgKgKXgJsFDTG6eNpWtBxJMjuAfvPa/
L3lHmSqDD6z5W35A94daKR+q4bEEKcjN9W8OLX9et899HkZO4drt7TlTg+s9KVip
/g7256av/Q+sFhKv6X7FR9VmKjTKE83JYDAE/N4H38zaTctaHV4ftO0k78lr5tc7
0870x7KRweLODxcx3W/CJAAudxMY4w+s6GOsX/P3alONXRYDPzb+e9xIw+nV+vur
bQXdZcSPyJfRETcuXSy+JwWz9LuWoh3NxwbHR/AExUc9rkr6rE2sh3l3eKmtqBui
DrQY9sj/1AsaMOZ6E1V64XL/AkOiAs7BG7fJxE1+bFH9pdUns/lSUEHwqZZo/aFG
06p2AMT5jR3YNnZFqmUN4GdZ705ycJtkSv0tDhiPNqVdZJ3UB4lvwKYNbGOw1/99
d8Z1oNvGIhypBG/HlOgx2WvKRU+PwVZLz3XjCxWTnMrF7B5b+WfdLO07E55CrMNp
ij1r0tQ+xkks6jE4GBWWSa48gdYI2+XWfE/uXC8XJ+Kb4w0ao+ULMc2AJM3hnZW8
VRjKJkoaP6NIVY8sa9eRt1xhxeeZMkAiFiMZMrhK4cQf2Mfa4Rfuv6nayrzVr5wt
c9cI1As/+FtPg4+u253NXxDiCpYFkPkFwDrz+6lkGkJe89qsPUYPvGDuMwDTK2yN
DMErtPYujOODzJXDEKZdJUuRdvyc+aZZmj4lvJg24edgTF7dXLBC0J45BA/hETF+
lzGQSPUG4rR8dLdjmASnr6kDOYipZna81YwVBkNYZbStClv8ygzPZaPusLjW8Esi
Ebf0W0OA1IwS8XlCSJyXWKdhykiDdtxkrejobxADFEGbapcg65gGvvPZr2dW1Byo
S5C3uKXAWYxDQODbYPva8OWSN7JmXAN93GZhHQs3ZclAvCOo27i69cKfftKmTthF
m4LU2TgrP9rlEgdRsT445X9zGhJWZcyzeXJffRV3DRAKCguxnQc5cmzx9jg9pnHA
C44zTCpKCTnxf347Tns24C3OB3fAUWn+qeZC/Bz5HS4sd/X8MaVDiHN723Slbcbk
/Y6ZHyID0Rqx6Z4viJfij2mG/maQRqiTUZT/U7jUM7fvmtD4QpBHmaiOeHJmtlnu
IGU3Y4XCBVbJ57w23befMzVdz7OPlcePowQN7himdgW7eX+Bu9CjRYCoYOxPlmEX
S30/n+FlW1B3DFCClxgSlwv+w7HkDu0r/bbhFjZ2Wcmfnot2teJ4zbUHLkGY8Ojt
hgTTHFq++3pAvAP3vxrWjuq9uyboJ6EYSFhzArV+gbX89dgQMSXIk1mwqxM6kUIR
mf7XtTBqMdOgcDiwCnH8Dzu0q7Lo7YVgjdAr8dMPxW0irLAqqk/Ig0SFJyw3gvF5
C+S/hly5npi2XQEqrwiwx6fx/3dURNDnGMoe7oFd+ctvxRUGIEI7l5Fp2RHl7hk1
5SkK+j/O3DxDrNToDIRjnAdExPTyrvBcmxtuSqOLDo+s42RdSMzvH6Lj6whuxQq8
dJyGkmd0ClWxu5RC/VHXYUIkB2clscOcnPXz31bVROM8iwOvINydnBSwmM93kZ8f
5hfe92R7XMBUbLWiWWu3UJuGvvWOPF1roPwyhhLW+W3/N8mg4un2i/UqYF7ggdgg
ubw7tXl9GozoJWyEQIpDrvIjX9sJF4P/X1jBLNk70F1RQXSX0ad4llFXH3L/S80o
fcP3NHtT0qquHxcTxwHY58hh7hXo5lsgn6sYV2TbIZ5PrWL6V7RHll4eYOSxI7Oy
Q5wlIDNJOhhVZUdQ7ja2NgmZyuJjg8iL383p+52/wxcMsn7Y4O9CMC5CPe99SFas
mJkAUrV//eeacFM0TjYo431QeUaGcXkR7jf8AhJotQLfzRkftWno9U4Z2ous+yy6
UZKPOUx/C2gkmr9R4t8n74xpHf49AuFV3fWcN1Zryfu9s/qFh8XTYvZSr9E5M53U
B4z6K0+1izJznOFVCuXFombLc1Z1JG4+SkTf9XIjqVdxjeDm23L24NwHRZxtgrz9
xElwq2i+JpPELFrqnBLTeWiwLN8UgBsIltixu4/lW5ZXOUp2n2GW9/EnJ6UOI4wl
3CkQNvWNLLsIEdSBLKGBMHChpC3LVkptukTYkJlWJ+Dmhqb9qAsCMe4J7RrG3P4r
8qlotTjhO87Nh1JHelLJ1m+zOiX4CND+478VThEQ8MplhSDfu6UUubN23iEzOu2R
y3t+VTUYl04FEF1Ls8REw0svKsMV5BqAxqQYk6Xd5xkpplE0G/7ij1BzKcU01LH/
4/GRuE7l7jnW3/rcPgpq5JfkCPe9mlX9X+Zu+vGdx/0zTaoLVyqIKWb9Fv6GWKK5
sSfeOBIn8fA/CUfhGWH+2u5Rtq7FB2re7QCvK7wnAtxjdSnqi2Rs5XAy7qN4tahJ
Oce38NV308WuPGpIyAS5sZBgyXfSfZ1cH8lTz+faRJoHey55VXM89NAygQ9GU9lK
iZOolfiutVbOa0YMqQWFJrj0+dQg4tWfgTaBCYckFNRqRDx2nicCfN+hP0fob8WF
dm1I3WlfE581e55K/KBRSWqzAnOhym3unlMv1K7DQS3BHEomN6GiK8njijGirPSC
s9hEEI9bhqwCr7k3NKgmD1HS0OzHug7i+0BFg98d/Csama5HpCyEWIjoyadanBGq
g9rvis3JqypvDC2JLnxjHKBxxfuKf0mjlCUyhWUFZ0/XtapuPi/DCdEXiXjt4dp3
0AJuRgjvx64kvlehfnBb573Qi8recWckpKcmqBk+7HYVTFID4auwluAx90GMhN3k
27/DGNSikoXsOLO9wGj0qnbT93CSxbhQH/KMXCIxlZ/1a2hTzAZw8MhUZIfM3gIE
iFgJXWXXI+VQB1N5iRCXxfnCiMUFvIOsl8riFdfYGmMu1XdN8fOHteAD+A/gYojb
E6sbXU/Pb27T0OV5wckt5VG1mgiXQc33xuKqzPrsk7MblWX30sGihHcP1+zRiqmF
emGDt36av3u4aBxCFMnSq1a34KakPosky6WCXU92n/Oli9KTHmt5azKj51SMV4o/
dJyaDx00CMxIlnoJr7HNuRNVDBvx3c13Qb4J8e1u6/qOpvFCGOD5bHHimBO59A+A
jM1nO3wl5/TNuvhLt4N+XHvpp88jYliUfGPWVhakjcHJr9Lw93nQh8EjZ8PHM/mW
6uYSwI1yG10Bh2aY81gXK/ggzL2yZ7dK3IshiBsThxHUjmGSpiganGwP1BANSpYL
aSDBdTRVGGHfn3M89CkdUD913H8qWp5FV2Ii4LK4xGlyafHEOkW5HSymNrs+02OG
hQ6XmPkhHP6bHFCTdBUcB+KnCbfurGWlYyxfFqS94hBDHQP2zI6baokDP5F5PTrp
IDd73QWB4MQ6+lg+kdTn8u4dQEXs/MCuJ556DyeJ94i+Zf0pc1lZFc8KSrLpavWQ
84/4/yZBdxzbTN1iEE2Kr8VScrPuyexCKf1Cmz1NTD8consyF3jf61Rg/mfI+2Y3
bLl9/gWGTdeSg11FXc9fZ5uI49NGyTdz3uGdK5S1sAWkD/9dLAfMHpr6qia/qDdy
/m1FVw/LZ1iGQ3B3yhriGiJKEXI5hCgj3FXoyeij8PuUxJXLer2Y/1yOU2h/2/Fk
VUhcPiqL395igiXptfYpoBh0775LyK7w8NpjVWIERquIX+QO0Hjkt8TS0Pe2b2sT
5uSY6cgix2+99OCYlf/1+uwVXw2aquhQJS0AdeLeOIMCVA7O41y/wvH8+c8uWT+h
rO17tgxLuIf97Q/Ryl8FekogaoTpAYv6xRplRQKysuTkLtBrbb+0SNrzFLHzhXNi
0IhkmMLslfe77dKAbj1o8uIqbrAi7uMqMIK+/ifBvtuoeqjOtDgVJBxsNixYEF5Q
2CAnsJjdw79fEszHledKubYH2MgASfKgcBuUytygnxf+/MJIT4WSUGXx9p7ZuXkf
ndw2qfRhhQjaJI8IfBV8LGb4z5NiW3WHcO4BNux/GNoq1VqtWFklJCFevF4fpiqN
A5G4Ypi2LauBQdlMFDxZhOp+Xpc4PrdFzJNt4MHATKRMQ+qBBRv7KY3O7Z/8ZVz+
XpgWXYcuORYaR1GmU+YXPHmEEH2QHqhpCV/8sioIF9/9RzrsHoPghDhnOjePA51p
5SP2HpH8AqM/UP3Jtyp2Fh7ThAxzZiXkkp2fC9K1yLpnL/8swKhe4IFccym8zt2k
wFgLlsUkUKdCzY8Mcv1j0JTYWVu0EwtXDF8xuqpIsizR/tnNfemX7C9tuZ3Slo1H
MyH/Dbj0oZeEp5iN2+aAYiUtnuuVVUydXosMhFP+ZBIDBre6yfreJrlfuOPkNU6M
EBMkf188wkFH+ph64IWwUO+yq7EDFrwCCIqZ3Cx9cxRaT+AJ0Pt8HNRwZqvMSYhS
TiPx1CUujeia1tI5hZeckX/XGwrP+apMXjM81oDJLWFjPYnZkyw8E+POnQoN69Vo
lU3xL3lPz7n7LTRAlFueBJF6lRxegx7XuOtie3okundQf6vgnfYfMj1HlUxhNJnF
MnerXb8gyHkkw9kB4NS2hAcPy84sC6l1SMRcj38HEsLvu0D+x0O3OqSNbscn6oss
S6XzspksYw5qoYXrGtQKouOBngY9uz8CqayvqiKSLlZlrj9RR6/RfwWhVk2mnUgt
HHDiZPSTlM8euJRl2V3qZS1U33jVUJEvA7LgGiEO4Nw7diQyhN9EQFzLkgazvZN8
gA9VQk93v/R5IG0HD8ZJ9xm9TCqWqeJCTGlXj5+bRKHCw4zKm4wjOSzRkLIJK85n
Z5XIIJK46IXW5x0SZgQiM89UmQ0Mw4H1gr7kdtm3COs9DFdTVBBaJvjvWH/ov0QK
SeWAIe3Bsqruz6Dr4TiKHOTU5mfcsBytz3e1/U1ruBKGGlhQ2rng2pgdrfsLUGd+
0unId24Kz9KM84GEGIkIHiSkKq7YN2QZY64bOpU/FPm4J4dXUgIAs694Zly+e4Mu
n1jFzj9cM7bArh7SGXrdeB7Qgi6q2oYS/2W+vFqTfRBtaOkoTpf3fMth4NUIccAL
s7F9gWSry4Bnae64SKrYfg1tEzfycWcBmnqaIcivYUFMFnVaASY658GpypOgBsl2
MP/QI7F+8KbLOwpVQmVDnfo4cxqkA6crKCR4ArlxBRVj7W32owQDkJkf2AthoPYP
7SSx0B5ApOCf8GPYzaYv2m/K4KGEkDs+HPqPIP0LmREwwUB5HZq/FKOS1W4UkSlF
rts6h0dRJfIhx9g5Lvo+S+ok9m5+Qj0DCuSBgSFqq2jxi0BM/vwgTeQ/QOb+9/Vj
JT/uuzr973UN8nDnUoSjGKSfR2Tb9qhRRt+3BD/NLJcCh7e7+LTsixC2R0N+nBFt
7K7YRUFDACVYyEEyOxfHqQwx4SmhzuENQv59Lw04NbYddtwvNcGTgtJ2XThVEbYY
WfI8DMKACMb7p/+IQUzYNHCOmuWPDTXKpsbzC/GNaco0ksKyuW3uUHCQmdjm0BgB
UCf7NQei6wLRhtX95nJqEw2f+tLsTL1ujgg/r7rpP0an9+jFxBocxp87kGnOkkli
vnboYe5xe9nNUqO9L3sAMW22xTblBhI9UT7EIkFi7aVBYKm3vtKs983Y/bDmvmWo
7oZQuk++jUDdbgVTZjFTyoNSLaaa3cPRs+3jDztdrjaSn1G4yaTQiCJkgVhaQNik
79PpVaQiRGPQ5l5izlB0KoYZWlxhO/Bnvryg6bQj32PIvG8EGJiAD0/1EdHUWJy5
wQyZkDBNv6SpHUY9gy8oFLp9yAb+ySjGUPiFBfPz2r86CajFgCBBgduD1DVFdVRB
E14/5U7pmmc/cmingaAsDALC9KO2vQuIRW6G8gPpUiXOc11LXd3q1WMk0ssIEB6S
8Jm26lkVSTde8SnFDZLGQy/ondQwyzfcYaqV5xrTdxPT6K/tY9QetNA3bpZZ2lEG
9KEgDBMGgvZMmXG45Ss+7DWuqE7PHlZ7QcWPZorxGFdXGAq3Sohu2Z9ETAIt5+cS
FWUzSnu4nEwTPiP7dYbTc1sog7cHjnnrjewR2p7nqKGUad30a+wJLOg2P/S8fJkg
9P/qocrzGTaMpKHavJHbAkAZ5i5CEORZlDvUshsJBUC9dguDWR1SJwMnwKrtENJZ
4lC2DNtL1ooiChPHzdXP0EoJiRcO/7yW2U1EqM7R1eEZTOqN500I2TYPaDkCO+Kg
G7MUHV8KL9+K5voPOqhOlRcfOrcoaNy/2uVB+Kb1m56EOryBKkzVWNQFqc4ByaRY
p61PM5K5WTjF/s3KHiV6wZZFSWK7kSSUMdqhDCrjHivPPRjTALW+aMLeLU4OkxJA
88J/fRXzoUhDLXtcdkoKHQrJ2sDFkDryRzYiPdSduWmyF/dWFbsxYSxTrfNPDlxX
rV4zgRF/QKipXsQNxI2rY76uRNFXw4KuDKO5YJB70zx6Uf9n8WcP5Hq1Rc59TyD5
4HmHpWpVTw9l6t4I6GPAkjOJU/kPat+Nu/cSCJhqeKY4KKPdm33xMIrz/AY0bK9G
v0FwTYtarNOFl2w+hBLlUEZvkgaztnlx4c2HZrZsg9gHNsVFl030Cm9l4q4UnyyY
I7ropLd5ZtmNBYUQ3HLdPCBnqyDhIuSu6tVyL99HdvG+pD5CPJR+qdJdmRYv9YWU
+d23M61r6IihTqHz3EaLt3qRFugf4WepNDjc/v/1Vr/MQucNCJDcdkwgCBDMFNbE
+s+Y+/u3wtwAaSSxZs7CSUaiSEtrRVq377smZFDkkpowipKM1nJoMlODz7YZ0nC1
XwZ7FnbAzWsLGgAxeREDKtSE+4sZXLj9ZQPnnbP8Ey+HncthECfOtKWAZNHJSx/t
IxQdWefZVTC81B6wwCDYnAVecxvdPiDQp4vTxBSQ8ngBIL3fzlXNjzuRl+//IsXe
K91ht00drgWuGahMG71m0+g9lpwu/GgUQ83CK8mEngsmHI3Aasp8E3PA2IrFzypW
qwJGjpE3xRO8H5C34k6jAWAa0M44XZMK4Azdkup1uZCEc/RrBYAuaAmAp/a8vDpr
bwLX5L89HSwnwaMmk3ETQ9UMWJE3ZHjbZ547zwAGjTp5sCECPyHAbsUueaOTC4tH
md+as4xoNDy/YiaUffHXF5yWfZn0jljHcG7+y6ewDOgTiGHh8dkHRKyyJQiomMm1
V6uGGAcQOqn7EDmSMC72myfxPBVZ3fWQwJms5aPwADuHpGTjddb7GFIDL5x8Q82Y
k73uRMWdD9uMwnuxGEwP5OTtfCTxT38msiuRqKCQy45oZLed6IZJ058w3Z6T7kPu
1YkfpZSTrfjclvE5o1SX6fwoM9hw5yGWLc3SV8YgoboWxY9+SRY4d4R4kfD+fbf+
5KmuoQQe6MnEhQXsEAGo2XVqstFAfBk8gQvXoL+f2ODGK5F2Qd3EmbvnmFB9ANg8
fj4fDwaACQycAwVdCLgmetphif1OvjukLMapCU5IHIORn2sMQ8PG4+JTynvibKnB
qgW9j9EO4dwH3Q6DaWEg+ncw/kGIUTk5fDbA4WANZXUVJ4TL0eQMpWAaYpXGDfqT
nyUZyjcQgX1C3gdzpmtiUlE5vQ5/rTm0IKC/Whd2+ggp5YWfjlHsVg+hghgY0SCT
SCVhEnTQwu567NSCR6nx+xf3FqpV7kVx3eeC4EcPc6Ved/zX8VNXXLEjqBn3yJd5
2OuCeCghwlKREz/6dh6t+XbKzq/U2q0sJWtoUm79bM6Sdd7Hxt2CM9f0JGS8dW/m
Tc0iiWdwwkYkKgZSR45X2aygPRIpOFMZW6PykspuophJyPjvv1dbQZY8P+CwYzt7
8J2tI6BWmMIfC97JL8avVuvQ1y/Fi+IR0ekaSCRmQoUeQHjErdI+7dB/L2GEmHfM
55MWLhe8QCumSJlM5hfzIE9hWpocfO3hM1Gae2iW1IsN0ybQid1bbQWm+W5bcKjm
iZHcVMTVFCmixqMP6dIJOYN1Z7wHpedOiWyHzM1YySdiSOIIFcUZ9XC/0+KrU43H
xeFpxpvGq353BdGKpQ51tN9aZyX0CFtAATDia5I841ZNYhMd4grz5B3IM4y5njnJ
gnBqrb4htw18672zVSaZGtqCPSKEggNuB8+oHIOSp4JW13oXE9tPJs1oPD2x9aht
U51y30XKOy4kcDNIFlhVfg==

`pragma protect end_protected
