// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Tp1nki/cCb/7LhLw9DX/VeBl11ZdJ6bz62f2lU0dDoKL8e+bA0DPPj6ShJIYuPeU
CXehnBkoRZBvYY8PqLed6Rzfi+bHBnN9Y3hMV9QebqBrEY2KxgZ4JSf0ZLYhSi8R
IKbG5MvLbsm+SFI7Hq762gD4R70hvR6k2KqtUK8ioC8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 14528 )
`pragma protect data_block
t3kq7URaQHbRZ4Z7/ytsfepqxr/FNic5MAgOHyrWWZ5c0KiQuAi8eW03dbOKvI9d
T1rm3/Hngm1EH+c0igbYc+x0moAXURPEgCvOjJDf1F+S+G/7I6k3sEjMe1N2nyRf
a5Ri2224bsEHrO9o2p7vnnaghvCO97/aIvMv/KyLRtxsDJ2aqoJ0UpqUC+mB2RaH
qf+alJTINYMJPOb+OWDVGLFMPc9hF0P/0huStfKmtuUaUy4ejdH0Bfn9CFd7gnEC
GHLy1YYpK/tKt1WiILRSQENtTdkIYfGK2ET4WOUHAnc4OEjKHu+hsV+VyxVHaTs0
tdcIqu/S2wuzuBu3WS+GdGyvUQ1OWiIIy78CeXBwGMFrwE1YzA7dPaa4mzpsjy3R
RwXjG2mzXNcttGnRfW9mFDnftbFaPQXrIj6rSPfWh0NwzZQT96HnCapGJ7/5OY4+
xJKEOnDLgpCGgv0De06PFLsytxOWy7+uFVY96XwE+UvEm6LvVG+1WKo8lPCwkmky
VYVVQeYUnIMUih4v83WPJrrKRlzKHjlQOvGjFlZsCOYL5jJCpFFcW8ZshmbrjpKV
51tC8kKhdD4OOxz+UqigtEIDRmfmwEMNR0YUzg9l/6xJtTBS30B/yx4vGfB4iA1I
y1rrKA9VjHr+SjwCIbt+3a5ys03LkSxDJvZ3lCCbQTnQP6/yI3XQmlaYy+41mzVs
6EIOOgo54tmKgMKxUWJgwLzhU3jVyyRV/CyRFgQCVLcdpRny5jd8cUfTIKp4Lkof
E8kloZyzJTNWSkni5gUVi67nvKzePARJQ9qaDbPzxfAR3+CcStYEb+EJGaEL7pBf
jVUyI0FMCOACVQ782lQs+0Q6ZE5Lttp4GDKWo9UROL9jEg5U7UKHX/CkMsJcZ3YS
6onCC3PSvX/7iDH9Gio+QPwMWCj/TP0igH6qI1kgb1C6WLMPVaC70MKPS1c5ptlQ
LzaQZd96mLXHyJ0wA4PBvjY73MOxKE0pJ09WuMW9ZuSiSEgSK+zRnNlosOXVt9BB
euiRPDUMeHy4lDMDlonKBfH+UKiQoZXOpwXuMxTAoKI1HtBhObtiZ8Pvfuam6UsE
dHr9dk7rMoR73spr5sTQsDFqrKPlhM383iyl/Ex1im40fL8LST4g0VUsvbQTiKcU
ENuTC00Pr653dzfBNEV8PJE9dSepkIVD68hAsywobLh1Oc3+6MpmPViqkdktDT2o
puyiCEYVeN88OKsKZcV00KH4FeWXkF1KSZ25Hgikr8r7QgMOLBVL1m1vp3DPhGf2
0phkPzdMKlt/S21RdJ7DIL1mu7kLXGgaCEl+7O0vDYHGqfJ9xsK0Zb3uU71kv64o
sFUV/85jOxaNnMSGApfvY5CoW7IXr8cV7Vp9CWs313MuDXqMILVtWIiidOpoqscb
rwrKbvq+Lgd+vHzJIWHGsab0ru4OQSjbV4eIIoHmnIPsO/hcP8wRuISiVSxEjyEc
n5g5jZ4Rpf/QKPVBpzj8EjlvoHi9xYPr4tEQeBN0eqy4I9/1UgLsqIDVHvn67l9a
4U1PbUVxDMUgJxGWHYqgKWc8g/bVMp3u0rEPdws0ADlz4vuXFyuslfUP/xmiCe0x
nWk9WvtCfPxP3MIoyRxxXfNbQI3w4SRuJYGt41Ocl/PW0QzDTood2UhmMkoXTiDJ
q+FxWfWz8lqXaZ/oGDhFXbGT6NEDJ5eChCMn23qiFwUNqmbJ24UcC6Gn2xCUAVEO
4FicPVHX5TUSprEk8qGFBKipDDdqVck7e10Y7W8OzwluwK9TOUxn8V0IEKCW+Mjr
4q7eW9a86xJTkbHIfnqskePMIXNfC21RJyZM3Wnd5EI8F/zfKnbyCBK7FjbE3rOv
zz0vgKEwUXxqpp5czAzqX7eswmZi7rma/koLEn888Zd04mw8/MQs+MfNJg8+et55
Vk14qZagRudriyWufkgg3RKvAwBQ6rEn2P7+GWxjlsfmumoAGAD4MfcUQVWGkED+
GGXYvZiQUt0JtqpvaTVWv7prEzJT80HzEmoQLksz9JTvulCl4xOgg1Lhn7r6y0A7
gVGXg7bqGUBDEDTH4T6SoMxSye6BXstt+vjb5RWae+YROJVFd0uiPqVXoQNePO2v
Q8sC403SGT4Ohz2CW7gsd5QCFH1AaUu1W92tG7XadYdKqMJ2heiG4MKdbeyv549V
jy+6bBF80pViJrUn7vieembtVfdnwztnbiliYNihbMq0SoNSFES9OYePUkTHPJP/
QkgebGPXm21H2M1TBBiGLm7zg1aOpRlI/RtBkKJj1iA1d7C/5TRMFFwmGnMwtDVJ
L2PyUfxGaejXONlbnjjHp6xoKKW6sZIyxZeKT4BhcwWeTMgdnAnVNNNAp2TfVdBt
1cHE/EXDJUyKqg5U0ZS2NwMTW4KQCihFInrCqy/aiKLmT/XNn4SWSXgBR3/CUJvV
mRqBz8xMkJ3Kx4veA6r9KjRR/nIu2HSBKYgGORreX6I6zQpYif2K8bv0IzoVd3ja
3UpQ+rQMrqjOSvidmI9eHGiu95z21rQ0I5cPpbVQJJYfLgHdcysz7yaryhg/zcRi
x5oIG2s6N7zHpHa9wOjL9HErAlMruIeeorvDcqkIMcey107DpHyAbATo/HbBOd3m
ZLxeHO3zYGf1cZNNtB8WFU7qS15TLEkak3W/NMWLZdiYvef9BKZOee13vzelIDRY
ejXhsNIx8lFuFSUypC9lNtS3mQXzg/BOjKrMa71b+jA84OBs9mcoMY/2auWgwbXt
8u+da732mXmowySD2XxHF8lGecCton/yNpqTvJi17oJukp7UI9SL9HvkJGl7T28O
xAH4k2+Wn08gm1yNlNskuatAF6emq84F4fPHJEu+52ToySnPG23MCb0MwcOOCRiL
cWDlZF/FgIiFrxFebHhXl/gM5rikOEkuiK+p1oJDanPxSRRRjyOv2oL+FYGmt0kb
IONFqapH2GqZnF9pRqzfNP0c+cCEVEAmaB8b8EnqaZ+vCY3NEPCO3oMMj0UABggr
EHln3CEa0HQGsGYJS2N53rka2+6cxmWjNyh5etBeQltLjbBdaHcNm25oZJbGrVvs
dees3sBjOMmXQCm/jRQlekpP6N6iGwnZFDZynIDZp7T+W3yoR53f9nj+sjzpbXNi
yLVZSIj0yUz1/nYzdivkB8n/2ERxvNNDCHoK+tTlsbTAFddw7bQU8Uf5pqeTn1xF
/DjIwYRqEKkfuFLFUAnPu2I6WBEC9xu9xuZifLQ3ldxKoYMOs8oHNBYzSJJejbov
MIOCDx+POeIqPxIRLSMueEHo/d+Loz9lai8DNOnxdld2c+6XbL4QQGAf/bq6kvEr
K303dYCOItqAMs6j2Znde0q7A8Re/26PlAxrN8xZnkZ2QuM6DT6Ka3B6qJ18FYOs
zVE1KrFT2U0GEEWrSupzklDCCmFoIzFNn9UHMWokHqDrboApDxTPsT/GyCfM7QZs
/6Eci/hgyOqGEjtVh2v3bhUJ2kV8IwvAIh/2V11zbRTZsnOX+XyNXJ5kRmWp0cI5
npFYe/IK6lPs8WrvfuiYE98NYiqNtZE4K8HhSdWnTs9pNkGBxEYHxaKmJwkgwaf7
FMgtfy5J3wL/xqnVBRj2yPyTFIr3SB10wFCi9Qtugt3SEuM14JsHkdd/M5r0fefI
VYVs9dNgRuRFhM8d62xKkK58PlYE2vMMzQU0ZHaNfFT4MXPWGW99PeKcY6LQRrGa
3Z30756L/qFloBModolSt9f0KIxZw0Al8w/HIKjZw78UgRdmjJqF2Y7x8g6elvN3
o+/Jo9PABDj+btNCvht0Z4JHJabULtGlEKPLfB1/vnR2wZw2t881wmJsuj02HF2l
KHKihtVjHCxL/IERSjtIYLEtwuxBR2BJjIHxmba/kxm50bX8KMNe8GyuuaNlqQRR
oD7CqlHA8UWjJSlAoySV0Lgkw4rCzv/9M9xVOR6PM2CCBSDpL0BPSv5xQa+WKSwa
zNngbHsJfR826mRbwr6Z7AfV5JariMk8KP/0wNtuH1HspIs4f5FEUGP4j3VJ4prT
64s2Jhk+12HxTdU5dWObz2K+KTGVyb3V8Ygt3TkOz5ao/3yFZ6D204+qZ9hwoOrA
u4vfdEhg+DgWGE5B5LNjHyQdTMMHzgwOvxJWf94VA3JDa4QYCbu1pbaTKK99HA5y
gZ5h+Y+5V51N5jBbuXQR/EblM9UB4VPvqmx6jQYxCFBiZc3l1D4ZP+NUQOdHFVva
laQyP3vyNr799tQF92L1V9HYtqYFDyOY0GX1Awb1Q4FlHllWk5GIzRsjD2aZUXSI
nzPrNA90mWjN857L7VM36naWSKx5KaqZW7+fTlbXx2m+A1iYz2LwlcmZmDFV61eB
rY+ZNGgHzdjAYvO42RQwgCpv0eeJxupV+NJbUTNBtfXpDCnoE+vIkwyh0UcC1Zdb
6pXBGFJuw4MAojdpXaw+RpOqtZv3liZD1Rp/c60QG2nj4Lk6Yi+Ca9PEUeQWTG4w
5ExLwWdx833yi1CvSeaqBv14qYpC3Md0oT0834G34i5RcQbozyIhQ28l9ryf8p4G
Ikwtz+CWf+9jYVpm9FIakhtlhnsWMoVjxn10fO3KOGiHDkn9Bm1tbuYRh7lWRGBj
jY3tmyLpz5D+xPXSH/w18uF0iwiTwv0IT+Ns5urFRGJFX8oo1ZEVPvT2XW79VRWW
fH+8Eg68aFmdwOnkLZe7zF1O2WMieEItTFfV+16cM6xILOleZLrJT+KGddqWfNoc
pOgp691UpHpiXW4iH8R7D96yyaBdIDmwegVygJhlqCjq/nLy48xZnY5tGyQqIZJh
HIyYErZgabzdZZcWe3zeQ6QsYl0mZQyl1SelKDjV5oKv1Q+sZ263Qa1ODydSXc1+
jAW66mdWURkGrBrie5bOQ9tTYKuwrTo3sL+3xYuMxevoMDbvU0tGwnmQ/61uDm7L
Kjmr5n9YsCM5HKUmeNmBgH/kw+czC8DHrGibwvyjqlu9Gx5QpDdLdxjnfOJlLk0q
5KYwKWsJyvZOtBzJCgmICjBFmvKVsBpTXKERwWtElAblsfFEHOhelXF7ixiyKaYU
IWVcjKpo5BV94CElHTMa6YbMbfYuJgWM0jIIPtHlySBFyVlJiYxWumRN6875PD+m
AdzX+/TjX40XciSzLR0xjG7FOUObrUluRPeODWRqXRkqQ8bqnNcRmvP5bpK0PD/G
J4A4gXvJ3xJ2e9IIsmVemS/KEYOFkXjD3wMEcXp+AAVRMG5K4N5cn18y4P2OxjPM
uw0N0cgHEXZPb3Gjd7cDoPklZjHMkKsicmYPpkxEebl1GVJmZPRKEkOux3iiatJA
HhYWOFlFJ+ovZy3y87ZhnlnHjRVh4+poYNew2LwF7Qcy9fQaxsDpG9OeLeJUCAmg
kSGTJuQRwqfr81pc5fDOyQDSyfRtQa9xzJ4aNn5lNjzCvu+nAUhqf3N/Q4BA0XuL
n39XlEU7Fl7rGjeJ37cJQm7Dmg6pEeQlWNPjHRqsLxf4Ko1DjUEcq0Z3ShyuqTGo
hQwPOTkmECUSHB2DKzGlQPBVwh9uZsEgUq7eeOhoVoYgMRxegaU5usYrUf0ZglHA
LXkd0c8qGq2O4usEwZvgfhW7mt5fSMjIMgi8RmVeb+ETjK6TeS28tiZO04XRKKlT
bIauLblXK2bUbdN0GuaZZhI5eXPYxkaXUNJlUC5M8CFynUJsMkNJBNXuFChVwtQt
kYJb/CpggH//V4a/XRIbOFLE1ksiWbye7YZ83RiopCAm0lpS0Toalm9xRYAmZMjp
1XHT5gYcHN2rz0IfbjoKK4aTiWLMfoOcuMirf4PT4p8EYIqGkU6reIz/m+M4b1HD
mrf3rqyS8eeYZIuhmq7HRKF5UlICI5VD/U9cE07Wl3QteeHhqC5Wc+QAQSwA3FKd
E2uthbz4QRr27hCnxYNqvT0O8ZMQ9eHnbK06m4LvVE1DL0YIinZaOIupxGrQYZmJ
fwKpTVYQ+fSG8n2mGNX8r0B8XIWKZnAtAX6jt/6ING957u1EeyVlPjTpvvhKh4r9
zbc8IYOv9sbCrevoXd66IOjjvgqF6C+otIhcusiOx8eD4ECxo9dXOd7M6QxSV/E7
23SZiQFKCKxyjoDT/ZOJnmF4Q29i6nxzjbckL+/dSjdQBBZxf7ZLenWaRSBMhhjS
bm1TgwBjPURJlpwMw+W6MlS4VZYEtmsJwDKtq+78kvY0VY8qmxbK0VUdq95ExE4V
8zwltN8EVcMyhek7ZlCs6Ovo0p0rh5Uz3WhyQhlRH8tvDmzEDNaERpVMPqLbpxin
UICJJE8hFNLbvTBXCRMixWIMaiCvtY8rb/ynhR4/HQgfzWwu9ia38GwUhpUKuekx
LRmzYsd/td9+MFQWM50aHXMrhDx0W/QAw1yzTAa1nwwaN+UkRdGAtAOEOJjVXqx3
o15Iqmpfel6fpTG2GA3aIZFAM2x5dg7d0Rwfn/uN0EbVA8d4hVkfOtb7hmFK2Sn+
p3tTC9B5KHYeXXWeP1Dm700HBbejenvl876uaJxPecnZSIafXCwyQTB9lvnFjm/C
o1imaU+AQLlCiRFqVmtFUmB0ApuaMRYXlgqY/5wXmLdXbKGy+KYUmB6VOH96waqN
rIj2Gxr8AxH1cw56ELw3lmTefl1HeyzBpz19f4aypuZ1YXWuI7OkhXSN+0+qhfT3
MMzaQY32QtIoXxQkshh2paBFcGAhNEehZs1h1ajManNYCDYu9Ym42/sD9UhRyAmt
J4Wm9f6+taW5eY9lTCMrCbLsRBFoR8pXmhx8x3oh1Xl5Fv72WM2/Akqm7sFq/11j
uzrpgv+EHJyPhv7xcrVVexDUfw1DSkM2N8RnpZ7vBxSnZsP9aULGqpIcb03GnZ70
qIDOdkSozwlj6GXNKJeD0edCRXvxiQfizbXjjlRwqEwtkYVCxeWfg79cNfnW0Cy0
zB/FOYFE5c6pdzA4ASMBwtauvkBCZNlj+n0VEYZNVzbEV+E6gvW3VmVA+KY533SV
CI2wZz/8t8GH3u38mb5oq1lS7N4q+QUCkMC8myvMYYXur75fklsTCYwZpofnqK/I
gAuShvYaZa7SysUYaPqR2ylWe/3HKIqzvFz/Qhb1RXBxQLKKwF9cd88rOECESedp
4x27w1oFVM6JoOk5ptWhGPxjJUkJxLn+I3SsTHd0G/tk1Fx+qFMqD18ZSDozhLIz
cOrzdqOm8hxpPEua/TmZxbygIq+5J5FrxGpslj0w4A6EK4YP9cMe9Dchulc8xBiv
GstRwBFlEWjHPUFde2NNj8pBBxao/Yjr70lagYeeVw8qKmnezboHvE35SktknIUH
kf7dYt2oIAFs2EhWc1Pxsm2ZWcOpDX2cAOmKuXkgmiIVnuo31KEijzz8fvv1fANV
jP6IiME3TjTDvU5q8cwsou1754W81qoq3K7TePPgd1BRAk187/14+dQVZXjnz88V
GB8iBCatJNH64xXq4OZl4YttazNpk6JkJqdnu785jfdszge9GeaLGGaiKQhHUNwV
LNad8gRr6XPLHFOKttmiGovvV6h2HrqNkpl4esgVKyT6YfOG1VWxacar4v0tD9eX
l536VpfiAJPcfoQ1/3K9uxZwvDleRBtxS/POm3kdMYX9l+wbKANguGvZS2lA3qTn
lzfcgZMysQW0jrPp4BnAeHCrPQPB68PQyCCTnlStUqu8Ta8ImXdrZQ6vXZ+QtroK
/nPmEhR/GQALFRhqyRn99QMNYjUJE/l3J7cWfvWywR+KT//jYs8jNwmRcQ15SIKw
ywXlC9Bn0K8yBNYVJ+U4hOiBasSbsUHw5hdFYvJaGO1JFRSuVfiEkwQf16BDqmgd
88MUfOfySZp/tm2iiVHjc2VydWTaQMQd4sNsyLVEtZj+rqsaZkSMwluexDORluaF
lUki0R5pY3rIWLzUHiUXU9svPk94y89kJszgOCEBD4ELKUclCEzaixF9/UlrTd1+
d9gTZVNYykIZW+Y3a/Fu+GYo5CI5gvNHe6E5Ait/DyLoZ6goOLOIQv9X5UFwRl22
jCqI79tQ0nLF52d59zOTbz8mIvaNmCnGPmOo1e2sTT8cQHEtCCWVuuvJmGfkSCou
3aBDzr5Nqav89D9sUxrKi8rau7NxAo2DfNmGZ/vtxX2w5SxCqXRJdCw8d2coIW5U
e1hyu7sTXGdHgPWzni4x7WQOxDzaoSg5AReavhsEVH5vsbTcDNTT9Ro5LuKbxezq
QIAZhqentEHpIyQbKEnPn6sjBvZOfbQn7Nkn9HGqtZWiXfdBZpIMyZ0tJi+MjwzN
3qGWAZZxH6/QNKD93v8B9Q8L49HZkB7y13/WrKeQhyjb02z2QW1fGc7p9PW1OHck
l2M5gt55L+lginmS16dWLbsS+PvhCCf9/VM7o5Y8PdteIFf9VSWbINDxb4nYXLFa
+SFKVeTOla1xJ3d+JlpcfFjg/vZtZbNVQ3IrEJFRQ9UBz+fSzxRmYUF/HQQT6zIq
fXi8Kvru/cnqC4tlPs52YpIja3chzyhqyKfcFHhhc/ejN/AxUyNI7x0GPDXsHjXe
kGbGDrHS/i/r5ilfFTJyLlI94GyZuiMTWBfdWkm4KElDQZPp8h2w0e3cgSk/nFT0
ubs+sREcIgyt8w+8Czgwv+jTnfjraNIBVSJsxTs2cXwQD0QAo/UkQ9aVNjbPashA
9f6yr0s7fI+ltWIpVaYLL214tPutEkQP1bMRa+DqLZH6jCKgLUaVDOlAnvVwwvDU
QzZaF3HPVs5CJtfaVvPaTvPOeQ0fctgqKgo61QrYjv/ygJmKC7O/jFi94baAcI2S
ePrhAqTAA+y1FMVbAUG+m6O4CAMSTnYUYL6NxmIX6rWcPI8Zn4AypqJwQBVWNzo0
eHsP/6QyqLasezp1XZN1DwM/6gFLJhefQkixE9jmlaKXo/A9Fo40eRRkrWNhukMj
eFBESUZezdbsjHPwwon8UVjBXSD03VV/OC+LwPwuGeYlHj4nDSUw/MRCCtU4ku9Z
5Q91Rt8sJtfFuuGYMUi70y21W7cJDH0w8WpHhxqL+Pbl91HgYz43qKvia8ctdMIq
u7RR8ADod0LO/Vk3Kdeix1ve+ZMa2vJ/yCKbJpZzGnCnVDuE2Wre3AHtSRmA4y1i
eh4GzVISRZ380+8PPnI8APALLgmrIQryttXbt2hu6tewapO8WpWthUQSWdXXtC5P
SgbR/MHc1jNUVXksebs/GQVyHY1pOKASAnOaPf6iPhHoIk2pB/UCTRWchznc2Z9a
STf7btW5TTJMU0p1ieUsN01L1k15bh1WhMrACKvfycQoAr5bIuv+Kqo+hLC/14jO
VxES4YWrAHWW4ll710JodJ0dxhLbs4JDZyBBvQWMLqzkiRTnzyM59A0ZWj0uQLJY
I7r5YJAYIVuhAYjz4aCq8oi+YhYF3nin7zZxbriE2i6y4ffCXIjj4A5E6sHgshwj
8Fo0ArO+Nn2H2KPzx+8cKLK8YmyGCLzSO6cd5G9DZZScWJASEN3ZHj1ZnuuhrK1+
un0tGfgNicvP2FQxi3RqEoXVolV3TLW2/3UKuGBk7GOyO5iqxmkYX3WI83bmndn/
dXiRrS8Z9POnAFSfZpCKiV8IolbKhJ/ZKBKloWRJHXeJrGTaFZrUPpypdfszx/HE
4gdWXaxvfxUBlewoieE27R0YDQCdN3PKo/+hOWJdv8GnJF0sdSY9okYf6KlzvDVr
aYoswp8wtutGbmoEZNmeo14LIWwVCTPHoRfGMUaYPfnL1A2PaMVRwWVVbh4m8t8K
BiMqBAUu89Of6tX1bWBgZJyw60ExGhwoyzbGuosdGGzA0eP/fbgHPyQG/Mjr9bx7
KbLQewPpUnktaX4MztVMR3lqkcd5HVrAtCkcPTUvuHDD6bDKlkM02HfXcaBB0ISL
pdhfTGsaPKWnLElN+ypv+gTCxbNG98OZMjwsISm4AYzoXxQ0vZawzQ4lT14kl9Gl
jnJkMCds2JIVTzJpsGi6HLiGiEm9xUs7Y9YEmIjdfgNh8NC+k0T42OI4zrUWQ/od
GrSH6tjf8IgDrufzu/T2ED9KYH5fqhtFecQOHufayQkjVK/u6jV4+BD45jjTo4T6
9o/xMdWAAk//EHjxiFhuJJvbq+4eQENUqroUdn+yhsh6aUdV2XrmEBFhSOiXDGT3
+WeBXF6nKjbZcQwiOTICLSEoNEvrlDTUSGu51zmn+sbm+Q/SDPMsaX9AJiAfNYnf
X4UXLWkd97fNxw1zWG9T3NyLLfcosz8aMC9oWxoYN0MkGRCoZ9j4sUbjEaWhb/EV
eadmYJgiZ9FjQEso3nfEEj4sPQiGfBkdQsOHyp4FDFe63M7b2OUaP+7SqUaMqlcj
7bXli+ZEQII3rn1t7QeeMxf/+TaMS3dqn0xWl2Yq9rs0KPc2D7JiGLJW7rzUnVob
y1/EETvKwaWOkzfkm+V7FUtWyBR7uy8tjN91VL6IxV80GvHBRPiK5LD99vaimAea
U1vdhp5/9MhNAvCWVPJWRHWlT5MI34MG24gRO8iSvvI08kVTNre1krgISjVmIma2
Wg5v4MXhdcCrbiDXO0CKOMP/4COVm0Yy4l7jk6yRfgi7GJOtiHIR925jy0IXtd2J
+7RgYKOboJLBtxkIOQ6qrDDXoxXOmTtdNJDBF6Jdb+kcn/e0CYf+LKznRD+oEkm1
JpjNIADWuOUo8vW6e2fq9MAqU1JOxVLXTtv4z2m3xoPJ92fZul/IpWiiMPqd4qId
j0c8+AmdyOiP+lb5oIbCrmdstvxwgB+W7Rv8uN5Rsyl1nkZXDHlFQfS8NNvpIqja
00PByKnXPWN7tYSJpgKqPKjBg+2cRdAwo/NMjJmWkKAM6pOejjNvxp+SCwkYI1WW
mMNuDQv/zCwzeqz7i7OmUkVW76FpqWuToZLS6gM8q0SiMxkrLVr3ko3N54M39TaM
J58qFZpy+xBk0AEGBZgqepdig0wLwdQF8DtDd3UnDv1ElQWc1BR/UAfALGPSBusQ
TmLhvF3lgLnyXPDCAp4m3lK5ywoS9PX1PUoPCzr9NbqTyQWll6Q/PVdtf82jQUQZ
VoX2ZaMWSqKNcD1Mbfy57TrumGDrV950dZGhOWt9d8w1uNZ1yEirqoiLP7h0R6SB
BrUEa1QZ3v4T8on86pFy+LNZEOL1Jwu3kYypD1XT1HFnEpZpSRj1qixmGyt8+JNO
qhK08afPJTldApG22wIb0bhKZ+8KW2MsyftJAG008ud+S4atkc4tZJ/t1b9bnwJN
JOmOftM+c5OnR+YqnRA7aHth9Xyi611sGHR7pWnRPpZ3L8WLVa4hLsLqRe0l9A1D
kP3/+8phDwGFVpHoH5KVLm1gMsnDC4pgq5xmZXoMrqcyBjKOVjFU/1X3ER1NnlNq
7GDlrkzoM9acsbcqEalvbz2pBJWLYE8rWJjOwPEo5JMDgLp8R/kkQHq0TdZTefP3
1D1mi6DcFjtBzOybk8dfLkqoBHYNTu0lVRUSPrv2cTWKDUZFS3jWIC9+aRdEofkT
ZVprYPKi/VhSifaqXyKxeN8sK+8sT32KrIfd8jsuNcUvcHRhL8nfzBGbnrRCU8io
spWwArM07o9gb+VCVkert56AzBxI6Y6VVpfzzYJdO7Ha5c59a4lnHN/rjh6p92k0
W2YCL4ZMtD6u2bBLPRfwh6pDKw6fKXZglb89EKzoSY/sXGvkbwPFCdJq5qc9FA1c
Y1E7puXdeRowxOTFGddntkCI6A2zEcM3Ddj1VHuIaN9UVBowT36fOB3T6kUiwrLS
ef13EMZzIBNWdxyeUhq9dcmH0LZol8/325N1otfvwxeH3msk2omKTRGspb/eJthc
QC6ysjTHck9g1ZuNrnhUI1Z1oZQqy961UsZBuaTg/+mQpxrua2/x0Jn4kLavVLVw
pYqQ2Fn/XtngXX66y7vAOql+JuFbP3o6jq8pCwLzr/VHywZpgXvBydljGOYmhcvu
StpPWWuBWUjbqq+DOc9uD6ekDLxvRFM/yux0+tnffU2pXA+VWmg+VslRlse8AG7v
s/bwzwypCkldpnaSpGPcNJDgFh/oo4ljGDH4r4sB1qz0DgBamS1P0cG+VdPs5rZs
2U3kIgdeiZJ+EiwDUMvR9W8L4i2ejNB6Geby6xy/XhWQPnlsCklHe7waVEeZKTqU
dtkrbH+4mzoY/y3OfdR90QL3AOTBGgmELho9czPt9Y1r0MC41sOXXy9vKA56s8Im
ghEYgf032XvwqJR73Bh6c+1CveRN6baSwE6g+lgw1IZzIwjtpPTxvguieBBz6xPt
EsKq6SOfbD8K8w32Z8/YoX7HwgMfWtkjpHncZAUVIJX9GQY56KR/tlL//l1jkSQ3
BkEqbQcrwcuH1+qZiCb1w0yLxOvd7kUGNKeJA4I55m/6K98sRXIjejssSPfyjXVj
yHdTdfbM3IqhdAwq+UAqGnefZwBV7v0PFcW2J4X8JN3LkA8VYX9Zh59TolcWQdHa
95NhyFMgvjefphoRa0l/LZYClF7xZWHV18CMLdyWhi80EeyWtP6gqOcvGoWQ1EFf
Lv+ffGfZLDdw14hI64yueI6qtgK15BQh65Vk1Jdl9lDNDgDu0Umj0g6T7Fr5ZNKm
GnnMStnyf7dd2li6DMBomT1OYIYvYrDGCf6I9XZrSbwiWQlrEXE6pVabE9j8fiBA
DbFBreJoc4vg0z6rEK4fZDkdQGPo4RLkNeNt0mUdSKBbtdRt8lZZhNhdlMSbm+Om
dsTeg8iEIUiJzXPluLttj9yw/2CJ7BJ0Pm1WGnoOoLROmgJsuLm8fDl65qgeT0cn
N/XlZtn5O82ukZWHLrGV5+0kaVxBVX2MqaJweOp2L6PBQD0w0KotqUN7tVevPRX0
xA9ihnYwmXdanM9uMt0dZNzJoPPlbBIV9vA+DhIQ15VtX93TcvefgRNlayBx2DSe
3PST6FJzJF3ltSJ5iwA8DdrdU3nHgS5cLSdJK89BNmbbmsIUQ1Yt3BKrR7GK8rM5
V5UawLMhi1K+ant0Xapz8xu4ENHkmoWE/JhLVamPGoP66MFremsWlJMU5Z9Id4k9
SSqZptwQu3NaM3LfoFGfW4KHZ+H78JWr1MwzVQ8N4bjroSuXHtmReFhhe6jDRIfW
deA346MCfyDf7s3vn8icVEP86nZ3Gt10Jx5psk8LI/k3KOFc1agmAVDcwaHOuwYy
3mdKb6BYFOE28MHc3IXEBF2tGxOS+tmKWI2NBpEczGS7BEuwJJQWSoTl0e2TKQTQ
OEi2j4tbu11Ald6me4jfRR7G54/A2HoJS36YnyWa90UktrGIfqYG9R0f1ibmAEg/
MQa9ndmj/kFo7LbRnUE9FGdXKn3WdqH/hLFIQB5xnOogB+caFM3/IxC9490CGN2U
Jnj5+nOFCkarEW9kV4FrRSAoP1Lgw0a56ojgkBMSKMSKiQnqTUaaNQuwl5qO29Yx
rbB6GHukXbIquwe53nR+3K/BKY3G8yKWl+ABNTtnQnZo2DDf6SbO+vcQiRetJohE
a5Rtj+GjjGdCzTCZj9kWi0cnuPmGRKOMTvh07afkX2OtFxQiart3U39+XqeUPgw/
ofbP8YqwB4IBIaOpgBjN2cGS/GCFOgrfQjtBhn0KSeZhRRIhfIlDVlvNLygjwnGn
N+fdz0Wzq+vmCZHmAAFkL7KQow/5qtnmd47HzOHLPAYJd8kQxaLCYJyHpcyi6muZ
/VBmWND4KA5az+PvHXfBKhGf/20ibvJ1hnbRN4PBtTn/b1OkEoYjOrPyeovz/1Li
xzBLSmVl8S9wJ0IxPCEmKtAYEIEGpmgcIGjRXyOhONsjhUlT7NPaJ73/rkEEvY0y
zXLyzs5XpfyVIZIa8WOb7AJhrVCaLdi/wYZMZXvcshfRNHAVgyNyO93HvXWtspJy
w/7VEH3GLbyCUpL7BFNPm9yKuOGqoIxvli3QwJfJydzWXFah1hVik2ytKZqVJuuf
QlBl5D+RMBluk8mX32xJfhKzJNfxN9bHCXZ/w0kL8/yo6xd8bPJF/LBC6i+d4Kvk
0OPTtCrQCveoIUGnaMkNLNaaXu7FcIH1PFH3ZdLp0IoGm5g/hAN56oPa6MSZ1u67
sDViTVzP2Luyrm7vtA5VIC5sVtX9GrOc1ledeFKv8sZ/HqIxJq7pkIDu7+2B1lfi
JQ+HT21vagxovhFfYwuRVZoJT3OUbkedx7YtCvCR9GoKW2IYJKGlKPE8XOhnvWIQ
lmVhLpV0/HSsyCSM4ZraP0W9B1HKr1Q4iasyrXaFgG83PonIS1aaO6B3YAjvBX/p
4JfXP3qNCULHoz2TQt3A7DbMJJNofxsirh1OlOrLRjj3T2ZQp61P+XGEne8RBJdV
xtcSyyjyLuVwLtcuZt7hMkiD5lS8quX2nZn4psYw0gP7dVOpLNKSnlbfsZQSlkkA
P+ETa2jtORoaMF2LwT//wlcEo1qwIBZnWKfxus+CqkHgoIDJNflNCzgrdWEaRR3T
B356vQ+ErZ7PW5awoKrzCkFRJQpKl0kcsF8nP/WoFsp8Dpa0rgKFAilRKiGvaoP1
VhJtL/zFEEelHa4eF5EJSnAqOYcH/jACLplhgCcgYy0YEj2RynLCSY2xWwmbm5Wn
hH4rQxLS5cd7Se3d0HOEmMZlf2kwHduNvtM7xj+pHRgd+CgZ/BIqC6PrNKKQlpPg
ED62BxDOBwPHbXyoN4+uOQDss+Yhg0KI8IDSKxXkJMxAuITgb0Fd+YeIEv25Xubr
Xz1r1hWzH74fD+ZMJfHpV497kjgaCxPMPz7x8iAM09ITmHLuDwj8++QUyM5nE0Op
hCWiREEp0Zehs16XLWR+FL5ZFJ5LUvBIlzg9sRcLwe7Hol86/T9piqun05lXmuwP
uQ8IB2lmHZQjsfLAQAy+PVbNH9SW0GQxUOUvNs+OyY7tTMmqkuC9wrIuhAiAfdJL
4OgSzLESKXS8U03CTPlKZJYuMsI419ovvm+QpqIn4Yt3rlSxq+wWwvzHag8A8F4L
86WXYXum6UFplYtf7uFec1NdIDrer8ys/8yKrGwJbYMlh3x1rVL4xNRPq8+72Ydf
kVvLwnLFb0SZ4LZ+E9kxUynDdGynGfUXDPFzRDkPB3pNhGVID/jtq/vTJkHA4eyH
rJwdNYu2HIAxniuEwMx6hgWnMMC6PaYTt/4iM2wDUxiBA7yub0DctdACvJs95hEl
9d9jieBc0onfnyzhBLPj5zELUgityQVu0YKFrMsVg0HAAqaZjomY9O/SK/9T75a1
ek41xj637NelKwMFhDBZHBTB+Ltltb+rnPHxHhH1/ELW3xTF8VeKIxZUBMOSWPCV
3i5I4ehxXmbKH2vR/esEMIyV+AgV7bB67H7lPxMCh2O84CtG22TF8j3snSPsKwGn
X5WBj/jFKNBUbjMomrQrwRFb0wD8BlELLYwFiOsAX0+QDllZIME80PVi24LF6dVn
PoUzs31eas0MpReLYjLx4ulHXbEVEoronfP36bT7A3FzqoJyaaNa2WmW7tu41tL3
XiV7zY7bqpmdyZVuXL+KMlyNDVtz5AzZdy/N8lhtv8G7lhPvQSpbyqUyipJ38G4X
JlkcIDDFXM4e13g/8Ofu7l74G5GIjB44sIOqkmCu/qHvw0SxAM1pQH2qu3dnI46Q
+d42EZ5PVXQ0o5wPOGcKIba8pvBly+Wlh28Xhs/SgULDiKE1H10dV7EsKgHvuXyi
5eNFBz86SO4hvyKdo4auQ/XJ/QPdYfdYx2gDs/hYlerdyyneGt3zr2qCPOOy42gi
XoEtC+7nA6fMdxcRVNc2XEaXEKf1EYyvs0dDUQc+L0hQQMK7ZxshTWNvpAzEpqD6
LvsurgmnTK04PLX3cmLZbjS6FF6Iv7sEAWLDH/YYBBAFm+J2KWGfbLfTcn9/Vufl
JDjfeySnohvtW6nDLex2EH7jHbxLuZ0mqizEvmt2Oy0ZHDURw592j88QJEamWRRa
9f44g1cvVHVBAFA3nwP181m8WY5QTw5DUiWM5rmRnad9ymzdsKdAbnb47YzrXwKe
6cWYGwhqAM+xrWf8DHAjrpr27Pm7rlrmn3uqA6Hh/uwLqMjcEFpgL9q/3+kvOaUO
a7gAJ+yiz/aUSSC4hy4TjPNevCDfR9gEnY/kEpPT7I6Gg5RVlZart7JG15Ci1W5a
DKe+XOZprnH9H/cd5gTneSjaxk+1AU27GBCm//jgBuJSxfm4AMFWsQnRXcv2shGc
XUTaWk9PscwQX2ygCPaTNh0tikUHAtnX7AtmpiWSjTstgZb5RurSZKzZvrDRsYXa
Jt3vU0wdBWxe9ETePMWrX8jmvjAd9Ffd+/EwWWRGO5cU0iipnlFuRySYeD6+SKI8
i0eD463rC5xQBTPjrFVAhBp8mz4gFBMibvZKec0hC6pWG0QsWwCUIMkO2wE762k3
7bJVCZUIgjQ0icdahZrUqw1w5H2SVV+zo/T2jshvHZ0F6/u2KP5iPhb2Bv8ej2sv
Oxjyn0xpFMxCNAhjRbEoEDk1Wi0trZ27s0Kq+DMoS1mzozXFuY4bs8kDCSoG0Bm2
dC1tsSKtLJh74+tklEIj/yBfJSgcx5eTHl4IVZguUc0MgdTuuyOcU3uygFq5HnVv
fUkh9wNOtGJtiAcaTgkoEmpO2pSDDOxxllTEovfcnPyY+jYie7Idp2cP+O4OyepU
CELIOzS4seU4OBx8sT/WY/LCfbSmsAIzMq+E9Qdg47SmoXUvT+DDy4XJHhV9Vug7
tILVai3e45wtV7xxzrEnLNHO31KlnIOYPv/IkgX5OIU9fiI3zr6qbxqZGyWa1FL7
P9EMHGyE6M8Etd6Iamr4rQrCH8WNd8cc9R9M2CX3OGrSV+TD/KA5x3FJ2HIK6Plb
bhGMFkLaB8rb34AUX21AOM7RjMdHJYlZhm/O+PW5EATg4kUcl5MwgV0cHt8LEEnl
uzumR/ykpgLts3A9XMyBbnpdbBk7uD04xdtROxhPrPSF2TqXr4lORFDiKVgzbvNx
gXe48ZimtoymRVOpX0ZiKkBO49mU+NXjNHxi3mnWjyTF0JoGaMaviDpdXcTaM6HZ
Hqxuy6yrZur/XxZxWH72AcAOM1CGpAwikORk6tIyV1ysHpCHw+vrSeYDQpW+yXHR
3U22bF3xGh65RS/yYZDSsMf8Dot2WTZGpMR16/PwMAc1UOjGjPuBbMYiz4DCg8a/
awCPAaFUm/pORC3xznxBmuO/KXY08I8Hs/IVYsT/Flp2xlq3X9gkI9qV2saBDg8T
Um3Ba1tTKRkt9zqYFavivCwrCvAcnaNa/gaJmBkwGKwlmN+sNvXgR0cPtVd+UnUO
8q/3Z2X5JXqbY3zdpfBiVqvfKuLxw68xOe9Y5FuUKFnV3RYdF7BfBtJIfc4i1FIO
0ZzFBPVljVrB9jcvazFai6dqkuKPa1TTLrqUhTpFlqS0ax3ACu7H88x/uGQgT4h2
zPf92DMUc/lK8qvN43Xxxe5FJS1C6j9cgXhaVb34pwyw7PmKWVErzaavjrI+aaDG
r6g7fBjtkLPOwNwNFJ0pcLEua5Bk6ar+WMju4krqqxRYttGSZsp8r0O4rugjwfiM
dNEXXd3Qhq4tMcH9nSaTPd9K6JvELraxvhMM7bZmC1RMNnSJJXan7OlLh4vj4xUf
jkmU5xZ72Ks5kVBh5DFDil3JvEtq+aZeQJzMYVVhuCbn70CWCenOrZ0rRmAFQRsB
Rhv43T8DqKr85Ztqd6stBnlRxycUXOeBfWLohL71AY7p/0mD/fXG6GWz8LjzFmO+
72Xqt1cR5o87Cu3FmI9pvXXLv44RzA2vxADu63L+7zfU9N+97dUiF/BtMxcb86Ly
/xxthm6eiXzyzAiZLBUC81xxvjU3c4W9AHataS6VMFMzN5Oc/XkCR9o+zi7c5ZCW
PogTMjWfo+Q4ObMdcxyP801HitS9NAOrLtxMedgTFIbNAhiG9lk/6ALarAA3Yvv8
FcLPNueC1tnykLuzvqs0bQBL7n6jMfNraCrd1lovsHguxVE50axXqobHjyZH4PYf
sycCdrD97kSSBLh7UIYZaBbXl6r7OOnuHeAXT+t8v1J8jxWfhWYexfIIIjdwaB5P
OT9todsBe4ULif5ZojfYaBEjZrxyoaw9OxzprcnDEAWLdvLBpE4kiEE0nwlbp97Y
TorJpBm6JekH8E6FDthUwFlKz+qt5N3B8oryeHZHZCAPVA0H6TQ/PwLZVOH49gFO
yei5z5hnjt4XrDgmxClnSp1C0uwiBPuJtwqMQNwyXlanip0wbB/obn/14Wkh/d7V
jyFBktU8ZMmp12YBH9gcq6UNBpTCkvm5RxW8rnssot9TKofWpknRKafCb8aaLmpJ
bFKXQ42ZepP14aehMhrTnAtXBYuMPTwhPcQpvlyi6V7DR/15qIEIqNJI5UpZ/QDW
Ik96yShH3kEcyQjh0JbTVeZ+8lSlFEFiOaK86hNXydViFIRYW7xGd5fEHWnR0ckQ
2dsBDEef5f00QwUk21JVy0euZUUIdAMLaNaeX9AqkQ2S8spcIRyuTvXMbxjsXAPF
WbAPpAJtU8nhR5EzHmagyeaTrla9hPTubA/OuA9qLD9XIqpXPqa5Vfxma0A/MYXT
Y4kK4kDYBc0n0hMIbUyWSovs7OBoblqqaZMhUW8pEBHj4k98tJ+VFt266zsGDTBy
KQGqcBrGJfTbo4tzPliy1SHUTllEAEQHIJ3j0MOF3qqpiP7SIeSs/KCk9B2GhnGX
OiLGnAImxdWu/AX7vrMotnC5uDiyE3q0kOQTLRHVBXsCuPZDoLn6Mlxty/7fLnYz
UnFcCsJ7jNMUdz3JR/y7g7GMnw/sJIzZse950wP+5KCkbxw9EiLkhdFpWSwEYCUV
hDMi2JYa9OzcAIgAss7l+QwxjjxAuoH6ClKx1OcVXLR+3P/4zb5klYRSa9rO9g+3
KsoHguXrjyWW6Q6/x1PJrN0IzGZ8KlpIWWDgstytMnqR9M4lQ/PVsKPORFg8rebC
/CfMclFyi2Fiq3JPVCmspbgNk0gGQFDBsTLggSK2ekK6hvjrIf7LAWSCi6IqBOKB
muIQ89XCdCrbqlYY6yCDV4BbCshcZTUl7UcQBDMoVOH4amsAWCGtg5xg9/mPQSCP
OJUkkjfDlxdjvVYc6LcV54qu6T3SvERPSCyQMwpq/GYKMQBGw2CwsPpkCrVmWS1G
4qKOKkbyb4FABBqR9L3N272E/IA3memTQAWk3Mvz1UzaUDEmyAgj006bmIsC7yDx
Qo3La3b6ee53cZjqC3FnItFxhFNpMvOHq1BPqkzROhVtYQ1aNLGC5e7BIHOCALtx
0D6d3PQ9xMHeH/AgxTYlStVm+/Q2y8IXBSUZoSxqjLGr/wd2f/IhjJOhjdvNCrhZ
NH4wtvJYexxRaRwu7jUCNC0/9oob7XvVn3lt3PkNJT/luUdBM16GSJ4ZZAyaVghW
E1NZBdh9KZ00s4UrbNLOjlhOcyX4uparj1rXk/nSA8s=

`pragma protect end_protected
