// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
0ZRrouiDVdfcI1CasOyXoPPrCvQDQKwNnqauvN/v3OrV4QQFfCMxAfw9O++jiCfY
2/CGJQqRB0Dfj9GL/yNT2dEFN9HH+z7t1IIejt+WVeavHZ6cztIqAHA0SwWh+LvB
OSGb9+x0nzXrHP297eVFMHCzb9uSKUCPRH/nupUyDtI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 59792 )
`pragma protect data_block
4m2cMIWIU5AjCzd94cswc7g6TL/lpe6eS0I3kgSbQHCuM4nCgWwv+dvhZDOhtTAE
vTDTBypwbR5RJLXuFc0TyetREoWIFkD2WfAt56QGr55Z5pc0uU6MMfTXklsI4lge
/DBytO+LaQGDwca0Fg0mbqF0aHzYuvWkV4/14AQ91LEibSCmvXsOO5GYfaWuEzf8
rTn3CC4eRoGx6auNym74EjTCQ1xtrTCEYdOW/D7JAWKbbLKxXHIQkdpVWtNsQNWu
yniMKMo3rkNA14PfBCZWMNsG1XCAp7QgchGFcyMyVQ+CcNX7dde65tztyEXU0nih
xOLYVTl8WoHftObW1RFSuuouerRa80YuyHBkylH7PTbJP3cOO7GA3IoYGVWhXS16
vKU4eJ17hS8HE2FldX1y5a2Y3Rzoe+a/WA2kcSz+yj/sv628Ou909MwFm74zwdrR
aGwYZ+7y8QCiinkf95QPmEkyHy9c3LB3Vi9PQJLMdz3tCNS/ut5BEeQYUxDl9npl
92gI/5OwZW8pO9eP+XMl3TtBGcEj9c/OEAcqtMODwKNK0tCmf0f2dmld6T+VIOrx
FGwKKgL6xPySYPhIr/2TuUI0NEUZqPicrgrCuJFD5v4u0W+QbjzuzWGApmlLd3q1
e44tt1ZPe0gIA2sz4fEqfBU4xi+Iki7YbfbZimn1XtQ1YlV5QiSqGEz2yK1di9mO
q+MjGI3pOU4FSoA5HUPkpOHauqNkEQU3P8ZkHTw4Oi+QDiIxKebDyZDv3enEn+uE
wDB3Dv8LvU3zRIEYfkHvyLtsrTS2qJ1Xfo13QFn1ckGyXIIpN55nwIPs19SK8nQq
pWGVwDBXhWQvdgdvc1d4Au9Z8/fozvlbhwbCAklmZO+Fd8rhjTWNZ5bNnRQBKnia
8ehac1E1cmOpYc5kvyBkNbqbETPqgB7jsTTd4duBp0Qx2J1rt6P3blgl3Q2aQOt4
nnbvHLfjeYw2j7D71bVrCbacHEzSHRR5Nik7pij+lLSfkUCuhxZo9QCHcLKwYJAa
Bbi0CB0RSGCjqbLV326bXdN8ZFhm2AoF+D8NbwQI2ZHFgX7aLw+ESH3tatCj14nt
4mJT8M5ynvDE7IeB8tzjRVhCPK3eUJt85zGrXJYfQQutFZsLrfbEb9WMaWQHI6hU
MptDB8DdN4CsOOP4Ic0R07HGpSkEW64hVeV/rNLv5TONkuHm9+8PHEZPBinSgIoi
Uf9LnsKgZtj9LSK3WPrKIqOl8OBQPJWCXywfpHWICpeeZNff8CU2E4nFDswRpmB/
aoEiL1YpcuocfnOhZxHik5OIRmd4qHITBCYHk2awlv1C4R0ODRq7PaRuvB3sDkG7
rZJIe3Izp/z7b8EQZpb9ZwOjDjs7ww6leilPtt7mmV3QDzkzd/cq+ADQbFjUDMl0
uwpoF0m0r/zh4dDwkhmDngCLXqt4s6Hii3UpNtlcg3kba/+rU3DH8CZX1AsYnYJf
JNSaH8VFc7gVsn0MSDLU0gky6Yukety9jAiI4HGqu5oyhqZ6ArlU418sA80r+iPJ
KGsDYpUrNpyVEh/GSX5ioNgHqnrMpG8Io4ZIAsePRe0TW5m6nwdbtFw5+95BPUEX
PaaZF5b8ru6+jqINw8CEr9jVqYmIW4RG/4lf67WjgxxvxJU95iq26Tj6wLFrr/YY
ySr0sWxgGWwqrxaOjaIIODehJYJBuP/55kK37Ukk3RmcHnUKwcQweSJldyvADV63
Jg3iRj6JNZNi+0zzgFIwOKfcd5H43FIEfNiyTe8aMJ2H97O4FdLdvTCXDwqq0+7i
BO5XlXVDJCAghkKyVIPFcCX1cRnBIkD9uW15NPeDmpdjbsqT1lV6hJQXbklyoJ4X
Qx8pez5YSsQmwf+tlT58Pt52sn5oJIHu/wZ9qfWS95liRqH7kLkz2Z2CwJu4UWPt
0q0XTHsnX/OrxfXSk1vlzCOfuhPzxPNCNL2SAT6clgg4lcwTBbclR27xQ/DBs+I6
6kG1tnOmxFqNmMIr0LCo5nWuO/ZVq75ouXWZOGKGJ67d54EC5y5Gc5uX4T1exk0/
0Fg/sfwmay7hTHK84Ulmyr+MXKsgUik+3ELof/u4/+INx7PPKogjQscMCA8FgO9C
fvL1XbTeIBi0P0R4gOcUR31zn/45uoZdii8wbsc0XGWM1D2BU9pvtLkY9roRUiS6
SCH6tsZlXRLj4jRzxCT39h15gYQCF66nq3luIJ5MRDyQaWR4EI/jJUDMxN7b+Nmm
Kh3tsMIJ9+ZBYooCgx6DVm8P+QYROEA4ZAOXoOyAGNTFDMHMlEOuYynZxd0qUv2N
Wo286IziCqM2+Ko8tRUvUy1VdCaw4WQCy2hUK0tvEmWka0MKd1ipppuG08unxz4r
ZWBPe9kUzbWk/xTdmbghidTcFFlYR4i+VwLi3weyhh+4olxXkecsiF+asnm3aO5R
q900zDMRc+7euFIB5e5qpUBjNrLVyoI9bmUe5Yr9fMdg4yD9r6eR/YjLSVwVdU97
wpOh2I1rEeuL3gSCo6Tm5XsthzOW92kpBfr87QMQWnJoihRCVxnEa3K6r7XeoOYd
LNORQ6FVNkeqf/Nx/XUVssxz4DpHew7ft68I+ybZYxMnxS10s4CBQmLgmEdw2R6D
PgjSIsoL1hDHDP3/kExiyQ+WAzo0hR6mXCZQJNSgJ+D4Mf+oOHMhBbdn4u+Qzb19
Ka7h8bNcCDEUanHw3LSTV7o6bIRkZv/sGtQIP34PErapUBpGw+gmBOJxJXUJB41y
uALQFFJk6rtIJdGpjHdtZzP3nAu0Euc/n2HapjAz0Q6IckSJOcM8eo7Mrm7djdZK
eRJhn62GkTmXEv4jWXzif/0jTHQ4sf3hvYGstKIFHr6oiuAL+h1j9csFGPLVsOtT
y7SAxNme+0BHi/MofvlRk3aXurZO5244r5WZebl6vrmZz/p6j3tmSE5EkPUP8f8N
SgNiOeFD74E45JTc1skNZjohWV6jxPtCTDs4idYY3yeK5T6PjVEvNLsJTt/txEj0
TF+5WhXSdoLUQdTiLeyu+Ajk4L1Ekn7GVJMxddDk97voX3yrHqmPegHA66l8TqXx
Nwn7Ug6fHvK8EGrpAcjVXng9RwekVbq3xcuryeBH2YouKJETPEGQvYOfW/dbYXdg
KZ4B0tjr0YGTsk8IkY9FHPghJJmUGpG9nLKQ2rHImjkPRJ6rWj8wvYA44VNPyyUa
TE6ah7xUZ6tktHdyU1DGNrRGrawVrItC8RLrBEDpQhK81v6C+mi/Klqcg+7mYvMP
9RHyrX0sNXEMiM9To/qHLYCkkrfZrbUUGjLCL7ms/R5F6Nr3wP+uspCl3QIPvMz/
mBeBpS/UIejgFGKgafFBqVWiPBkb3RvkY2BBpvqGSbynfg1RvmQnjhjKr7Midljl
dRt/eW5JckMbcfSwl/NRIVByF1Ar0OCyzt6OzyzCB70XO1fChI2Eb2gqOFSW4xwS
YQIkhOyI0OpG7BLz+b7zKJ58Zk1ABu0S3k+Ga/caBenTTOokFEK7cy4ZordSRqfe
KNnzVPSHDTHe3vbWOLH8iRlUO/xtWtuiftAQcRU+isBQEDW7zph2kojRic27s2rw
Pf3qR6g42HICQx4AhVyPxGJhBoI3GlZqEAFxnUfpYpB9xO1RobcYR52ezQ2cSsul
j1zdxYfF4x5d/CDGKMrdSks85y2R9Il7rHi2Iv/Yzt0vsNlkuLdNgVw+HtbEV/+Q
fdOzQbh0xFNJPL/xZDNUfC8MLl+knXC+L+tltpbalHsvto30Ibwa3a14xmx/2MF4
aNn0AwbJ6m/GeoD4hyDkbk9mKn7ncTXyw8SxFnjjFqcDEIhtEoPS7IIACGeBk5IR
oKpDzozs2u8oM0xS2UjjJbu6jPUd7ZPfcDtptJTYpyahJtngYty4xXclgh2xQEqA
i3i7hWlWd6tLufR2GtjN3qW6CyIOhoKbQ4pBPLF/xZsQ94UtqZCsPhD54DCaxeMa
RbOK+6UXkoSRDClKOH5e6XzhGnqYpNbPYG01tSY57iD0jqdVIP2jPzJRvaXKYOIc
sUAEHhZz26Vrfp3mI6YrEcc4OwKhdT1D5dcw8BXH6SBRqDTILU/Kwzb5eaqagndN
bmrjSHNUtmWN1wCrsrGgC1wCA3Wki5joAAnv/JinKhUvG0I6wfYzOvSmgmBW7byx
NUsWFlRVf1DK67aSMzwpMvQ3OAWIQprgcY8SpUbMwwuhlPxtPclxXXxgnRNnIj1g
1O5rFp2+gFcon0fLui3e0KklM61xAANyC3TNxNrBlrcBAGZXQo/PI9/h6W+Rik0p
XMFAVtFm38WKGpk4dL3VlfqpX1JoCLStZZQRU+/6ZPjUIFfQSQv+Gy46r8PmBljU
u4ZCex7/PaHs0/jWtK2/3qarEBEnNzaq1U8pdNGDQeKS/z7+xmbkor1EI6UYtU50
NZnycaK0mVK5/szxb6/fGMztpRSxHWL0Au3mAyMVU0S721hSWSuEqA0uibv5SXcE
ZAeyWlgCMVmZthJG0BbWIhrRx5GiZt4Wl5HoPcFHevQE/odiNri4CLQeNzX5wBin
fq45xUCLWpg52gVE0IsGVspDcxQEGunr2B8l7z+UQaJfN/AZ9eiAqyr4LEpLMBCK
K/j036o7T389I9/FW9gbDj+hF4pZ36ybHszScVki35jYUqklNFGNa120LGd+MTgv
bVILjdjDcsadeD2X9ZA9BW60qJCODqO5P8uOO0eQI0iqZkNg3fejoQgzanXfXHrI
8sTldGo4X6Hcd+gXY6Sl124+ZfLSUA9j/Wvlf2/cfxnivwPrFXgm1FB2xmte5qh8
qS4E4BCviIHDTEVMAjeWAe1TyrqWlm9vYgPDAJE18n46ESME+AUzkldPhTX2iztY
Z4ki0y0U04GUXkWoAv+GBmYtCG/43jZDwdOqQjn//vP8d6JNMeZIaA6/fthaKDK2
p3M0Ip71EbFxELDDNw8BaaLpbhOk9I1sGLAhUJ5qNhJ+QaDBe07bBu4C6Lwhjk+x
VT6OIRVsJcGPuwmU/lILLcWlRgzXjhM2Y4pcpEAw8oAJ7+IjsetBRnS8ta9hTyvG
GcvSKsCLAg8M0AFW9gBNs3QXLD2Q+lTmeyYOcbL8VtArHLg3cjmFTPoKmDeKFQHk
9zNLd2VgcE9ZzqzuroFt1wL7UcRkbhXy3X4ckkJ8DqfeBZmJ8PePH/yQk5lZLYDg
twqQlazi6NcdHSzkcM7A1lG5O4oTeVZdkdu5ExVkRqHsDacGmpu0/kuHOtu4fVDz
su1q7UkPrpb5ulOjSO0iuLuMN9Kdjdi/M2Z3X0/kbT0aPQ2mSGVVzSVK150fPB6o
7vyYXJvsaC0QPpxAR08mXsEzBln15dMZwxGHyKRnxfYe2KNX2qd8uAIxUNZmaHN8
DcWbNKv6RbBtwRpz1SdqSpPMNRzaM52nJ2sqUEZP7S9B/hkSJJ7pJzi+Kd4pIpfp
JRSIpv+s6J16FhxuqYOTVsN2ZZl1Sk8AyUhq59bMzjrLfQn+fLawmOEll6XrPOF8
1T2of3+h7wHlwVFrb6rnNqKfVYrLEttnUu97gZVU+nceUvGcg/gBnJcSYKAkqcBb
vcHLJWgFrK/WPB6FTZQMri8XcT+yaYvD6o/SHmkj7r840zPzm4FjVmmitXLj+eNT
/dZSYNxk2EH1ei13yrGWlaMeV+AETs1zcKVWvxtgBPtBxfk+BZkZWWvaQEMeN30t
GphFzPF7Q6Jx8yZUAVIDTKVfbHDEUU6QB6vSHz73IksAv5wxsTvRKACuN31j/dnH
zka/00hUUNe4WkSZnopnusYUdnj99TJtgAxlsZMfTAxIYmngbY6lcfY++IZfD2MH
Hcq+1n088Wu3EOGWiUTsGGWyuLo9i1qy7/nOzs7yhDQCCOMpeOJ3Kn2I9eVqFHeW
qVQhL95ulvA9JgwZO+NSnx6MnlV8xTzxn+KRrv9UsR2BZ16Sg3v6glyUN8XU1if4
PWnM/FAhyD79X2uFW9kqYHjagDDfrE5vUx3N/vMoBIxUPW5QbCPNvX7+N8EvPVNd
OOMcRCGqDTvj8fNOMCvS0o7MqLF1ftSYELQfmUUFexqdDCAKXxQYz+ySWDUKthJY
rWKUUdJPZj3KsNN9Wy6aBM8SEpRYxslWGDMYiZiMaqzVP6ylynsIy4eYXbMDAIJi
vMoZRrbeMknQvxHt2Syu0nkhQ5sTDwKtedB3GDq/RUX5oB3FAGktljhO2oDIckEK
tf3zl+Ld17oXTIPUvg2eVRNFOYCF1/zl8ox/MvpfXNIG+7/fGLkq+0HE3pkr67E/
ETtNt7EH9aYovtnEUpyz64iTi4Xjvtp2FMDgD4Z7dvEH/xCOjpCD0U93xSDzM7Qd
fXhDIt/aud27BJ3oEDymYPiL0NxOhaJqRvQVDPw/2DpLO6jQ43+LXbBaLWPyIpbK
ZhTRnT0U/DcPSpWRA1d7i5t3M+F5YQqrbuvkjj3rBSzAf+j8733LfOXfmu0g+9wg
yPbH1tgIw6Rv6qzuBXterkgWqZKV5yNZ9j8HbIQliVMy8j9ZnHzlTqllrt+zF731
LYmyw/1RDzDKVRKAsP2NN88LSaBHZjTzDz/jCp6jA9JQRkqWCctjK0EjptHEwzBx
zjWHHsvbEI4sRQoJbEhBoR/t1WiPdghnKUrwlniaINV45FjlUBVK+VgVAYG3DvHk
rs3yIohI1kNqNZ7FbASMEG9qB9fCaIR+qUVryKLPlj+gm9jP6/5yiAPzm5sCxLV2
XwjIazG1v8Vefh9aUW9TY13aajCaxOzg/RffdVtIVua/G0dDHe5nzXtiUudk+6f/
Zjn0Sc78ytgs7WrdJp7gHqvM/GJGsQiR7fKwKFmI3uMeNc4HtIt1Z2VaobMdgnMX
Z2P9DbODyPACPDW8Y42WFwHJr127p7Jl4W8iwpIa31AfTxfQSpTqhFewS//Fqwvu
t7Q3Jy9cz5EKIK08cKilIqvpmynBTUkOYziiNaruGrkHUdMJ+FHqRFYfHLa06F2X
wT22LxMHoEUluWYI8xdNfHb6jadxsJzUI55tzCF6VdvJJaIWWBtmbnwuIELSOl/K
RZXOwfH31eOnEmIbc9AIBpp9zzOBeL0ebVPMwJ++GkGJ3ltJcR3fi58kvPGlqbus
EImQ9xydhcbXGgLq4JsnQoj2jWTbVW+afIYk76wDSjObZrUooTllo0v3dMSOANu9
J1ZEm0YK7dhI/KDGozZCs3wl69Ygd7kb0iTJ/mO3unkftuZIqWjxwEJNg+7UH1bt
fiwTgFYBoMICnzZXIHQToMkbeurpMLOfjDCW/I6xrssP9GT6imIelYF8wshRrtkT
gCKvPVFfyq17RrWX5rEJ37b0FRQOQgJ/EF0srTfMOGOGpkAJ4J4W1HX97KQ2yLiV
rrcgabxOeFlyKFKGxbouBGzfn3L2zo543rmrc6YAkewRFVI8h4fD/JEMw65y6v/T
8HwtcfDenEmZin8BeVIPQQKL95nB65Ei/1WjfnB8fiaeIkT2y0sEOkFHGohZOvSI
X1vI2i1J9boBGudWZJqo4g8z6+7HcaMZ13S0CYVzhfMzEgnMzb9x8okf5ml3Vohr
RWbk9xxOnhavtdZxGnHwZ7EhVQja5YWVtNi1K5J2aD5wAMqAeVQyIRazr3z8TaFX
4XtkPsPP/aA8m4pdYysK8Ot1/WPz2d5/TKXZD0DJNOUp39X6myF4av6YHBYlN8tR
d4ZcuxnitQnztqjD9c15yrzS+mWnTb893+SkxXWi/YThpx+DyBnrKM1O1SivX6lO
jx2rIKSTJmf8TfR1lLcjAHv+lHueBVcL9vfjUAYj2QMM78MOQhySbY1HYpWEwscu
FIa4UkZjjiZP4I4be1KUwkbGLE97hfWhwRvbtjvCwuMj/HS/kyV5X6Q/p35vN+zr
qQcZ0X3NPeW2yMyQ2sfY4ico6wf5T+bxCPB1hG4s85J0Ub49oh57gwKec0AjK8eJ
IlQrEXy744x/Cp4B9RCnCMq8UHw3dbU55FQl5nebLkerHsFEWIHaRhAqPu6CP0MU
Y8NSO0N45SJrnTf5NYFQTWV6zFzD/W+bLUiDtnXKTLspq6YHRrUgo5VsPO/sQFgF
E0AofaqLdIEH0dQFV/5wA4ZX5fa73Q9spLLtNPJHzcf+PaG808w3T1IpgnNbmyh5
hBSdKPBtreCjKnnbaB+9cK3hC6cvCXwQwZ98IP314ZmBwHCfqg/nm5aQSGETeSqb
HeUSDt/aT7K9sdUYNH+Q/7+86Sxpo/LQKKFsYZkf4TGqVpBGOYclC+t/kpRSSIkc
sh5kzzh0rFJ2535V/hMdz03Y1nkah+aK9EwFjVIIO81CEXpYX0wppaKxQ0WPrAR0
8qPIaq6J8OzrlK3vmqjQL5t9PNcyEM1bcgj/EWpt0LJWWcsb1EzLDg+qCbA7lPUK
1xXTfd5ANi956a5Gf/5Y6QBuioPunz3td/4uHSGVxszO+jHXUc3MbJgS5GklFlEV
sZaUOADULrePNZO5fLFbHBxdEtkGJhciG1j2WRT3bvELodbbThik4ATX3OyJ/xR9
GbJcDn9p720OUQl6QWIGgiKcfBhF8oERyuCxbWthTBaCGDQPTzp9J+l25RjF3vdp
3jpkVES2+AkC5VrongqMIPDTxn7QsfVcEijX0Sc/PI481BcfBVg9wEZIg9KKX9Fq
wf5B5QFSRJOI/Rpqj71gJK/aSPDpEyZT4HYW9CHP2LCtxQVlkqCvz1qjSHwwkJsq
U0jwZH1znEcqgeD9P/XuY+lE0fzl3Yo8fJHCZ3AMYeujEA6qJv5NQEF+M/mVyofb
tpWs8bCWOCWK2NN3xovJoyHcoI1X/70FJkO+hv+YE3r1nUo8ww4bp/lkFU8bEnHJ
F9FK7LOPqJ4LMcjxtv9or0fxSMj4YD0uz21Tp9UlRP1R2Mh08K9lmzl+Z2/HMyng
SRrC2ahu0wY58CEJvD4+mvT7pxAN/8RM3E9yA4iV0qwynyHYjRg/9Yjyhr5Qw4ou
XcwCJdnEXEmCfkSBq2wApWaDtXP39R/tGk8Dh82w675Z6BZv7RMdpg/mnZgCiC+v
itNQBVZPMH4fNW2Wt8FqjZdOqVBH8yi3q51KMKGkBgDiv0sLq5Pr82v/tJCOjK/r
17Fkk00l3dBbNI9z8Oxkis35s9GzGrp/JjrnWM3DJmKsZUeimPYRRigiYMt3ipLU
sR9m6L0dAhNoatNLnI9jEZr1fxtDoQwyHseg9d13QpWugobiy9thLfdlfhQMgmof
4JWmrrF2oSAg+XYFMs8pI5v8K9aETRcQ9p3ZxmHjBOpbswtcfIND/C2oZVmSXPUn
rU23rXNKx2fN1SZZCWrpqYb3DkS2T1NREY1wJuMM0OyFJ4BAlS6UNK/eMqogR6kL
9NuFVlFjHYuXIXLuGxacttbN7dm4hQvza0y6vUu6lIILE3DWaHdNUIAUbGu5fpsj
BrmQZkAUDmSCAVYDRCh3SvqRz4Dn8UMMJcaZip3Luf2U1II30X/9v/aQe0+6W/g/
8mQ2r/QZeS39t1/FSTN+ZcNsJNK8HBsew6ZoGdqAEVn7iiMWbq/1IZkY+ahM6EMt
L4LdrZxpSDPKMNkFEnLkh6XzIqdlyBdUvvquXL9dtNZZmLF+kutAgJQ9e10w30bc
1472ZvngWmHkTp6g2Drh3VMITSbDDrM+lnh0/wAAZlIcCl3WYa+WULSGdIxWnyU1
Gj9Z7mf0InjJrlNJ+/1hdUkoybZW60G/M1HoSh2/10w0XCdoAIlMJb9yZ32DHGbi
plcN658ZevgVfaEhhA9Hvu2MmBWnd1725u5lqz5cBHKs6b5g6nxgaekunFQcE5ii
qILNRuEGVk0PvcpQp82Seq4q5Xe3hDcv2pZsHcnwMSefCrSi+c9WrxtMhvW9SJNW
n/7WBALcXE89wX/6O9MKtn7TzD58TtBgV424Db1UmfrHgM60pjg633KWVn8Fg/TZ
6hCYEoTvHRwxtXwqw8WX+XQ68esVM3rwoNKWILxD6TibpeApTBGduXBNixbY43yI
1bp/+UQGEqF+YmyU6Vaw+yIW2i5COejq3B23rcnWbDAyKKxm4MdmfM5T+rhPe7+A
NGvbiL9Z7CjZHYokV9Gw0L4g/IcNo24wbrO2xaR2LOsS4BI45twQPtwdcIFfiB/5
VdC7kYlYq82uiis/Q1/nvvjuIvmJ9q+MABsEHbsEqw/mw2uNxmhsVXp554CIj2Nr
KEqllRRRjRO9o6Kedyp2ynCEM74BK023TINLigQ8Y8A+rbmewbD8SWj7i+Cd7E3w
XUIUPgh1B39y/vcc5UVOtGIuMCqTWZQu1G9CO/BXoFEgePHUmpHelvXkHgI21dPt
6D2iXZuxL/HJmoWwYnYdr3PpU/x90TzS6Vr+s6OsjahLr/JeJT2X10Wly1+fxS/k
ifDDnqeHfwmBWPX967/GM+qt694nlB4Sw4ySO3lcXxGji9+RllMqHzLyuNqNAovE
+rhfWrwYE6BnDE96pHLKuLmj3cus/L1/Y5OLz144mPTxzBZcASc+6bIIGRDIBM3+
yHvJniwbPqD+kP3gRXlyjOQC9nMVOztK6x1bz+sfKBi9+3IFBHFSk1ps3SCa8Ff2
i6MXkRFgn7fRrKgxf+dNy9C+IYf3EPgyKFPvprnve66o2PCUNFtX1AfNB7i8yPkz
aZ60x4VS58Kut7LVIUFKbxQVoTCpMzlOmHmHQHCODuh0VY98ZM1ZyC22Z0aRzezc
Znfj8oquSZJyjQJBhiZfW/UjVK+5fNCVO1SVNtFPydPmQbzWdT3nUgM8dEvsi+4o
CN8OWCdFdMr+p5yl1budIRCPvm4lme3bguTifMKamCs5ftSCrIVdbKdtny0Awd1T
+bihfG1jISHW21WjQhpSZDZeJqwu3VlTubnmFvQrd9i5Zu+0cj1UjLJWFxLf66Oq
zL9yhgspyaB+sxEVp/cvkeWoBZPNrORsLcTovJLuyMXkh7B9zRujMZBaT/UrfLOv
St4k80xUkCfamv73PmRluaDfbGUntO0utPqem0qW5yXj0vM90apgGii4aUpvnOMs
JPKMnmYyPe1MFG05hWXvFiGYlj3qB46eU4iZqWvk4XqogVamMa1WyBPe6JXLd37d
NNpf8Ma9ckL56ntsSP0qt+Fg4z5sxIL3NfYtYW8MHyxGYN4vcFGDk9sCxE2o6Ie+
8tlLYIdUYdB4TrYZTrLjYovUoFFq0Qf7HIUMbjX7IX7oj0HTTNU4XASNUWqu9++U
qJapKhOzO3w+unGCC7jOYi1eJAiKf6yg0N5ZoexdTPwI3IEKHRLfBnmQ7dEJTib6
FrC60WqD1nIK3Fa9MLG27cf7G+xuMORx203THLyZ+bS9rQfNPdjdKH5/swWuH/UF
WKEf49YJDH3G8zAddiZQtlXXP+2G9vRE2MRBWkahUvoH1zhfYz7vKvPqFR9T19Tj
tZze8Gk85IJn1lfrQ+kokdmNIPPKPDzywmcV3kSBHfH3L5shBO1uwa6EzVRedSuu
qmKmBMPTnBDdZisVVULRUSvch1HXD/yHSjReOU2FaFMBwhbUcECvJiXsrWAT1sRY
R/GVurxQuqDeqmEeVQxy6n/7SwvRzfFXc+oosT1Pla3/XGwFPIb+iSV2CtWmcN8M
kfjDuVVR6qtz4dYJNz7A4r9+HXcQLvSX9W6vR4SPFPKGFP6MhLYHdUxjhlVrPQS0
3x5sOr1e90K1covjrdbFowsal9UHVCD8v+RuR6069l4a6MXfNT5mqGgnEzU8/42t
zgAPPkn/FXlA1nsn55WKu30WD5gXPZDfRLvr4lJZfY2Oj3MXyy/M/KjOhyKuOXiC
Ux43V6gO5VCMFHDp1/U0VJABfBWDiXhsvyac7a0vVDoXXu92s+Yf9pdNQUNEwblx
oz23s4cg0Yk2X1UMc6HuNJ17IF2dwb1F7yvFKvV6fGM1LweveLS6p0LxB7zUSir8
w62CAfYpLIgJ5a5hJezdaaHKz+rMjpOl1gWbOzTz/vfpLrG+GtC2YMOvkhTdCFyP
SrExSmZ5O/BJzahV/mlWL3Bhpc306UUZ3m9d7gm4+cELLpYWfCj+22Oo+tjYVjBa
CIvpjq+5Zyr39qqbst4A+XvDuAax6RLGBrMqor57oX/Q8qZyhlfFhJ8C9cwiJcJ6
zD32j+NQDR/m7HienxQ3Vp8j4R81gcUZsKK83RVhk/XvDII3xhQ4MmUfSnt14W9N
nysJmvyhrh4JukUZUOrcpk006unj/zVPj/EatRD3YLf/TUOT85wB+cXnRwZBH0HT
ZSGos+caj0pjiLFyQPeMR09X37zXLycvwkFvpcUGUzcDK+1MW6anQ+TDW4zRWTaI
v0GX+2NypN1GsG1GHaTrfHvWlDnR1mkrw+FEbmMDZQGnTueE+F90pGcp3mNqH5CL
Fac9NLf7oO+OFDoRj5Iqer3DO8NaDGFyEe3aC4JFIdpBzW+uO2eg+7DoUXGJahwU
X/iYbw336mmEilWSV6tVChH8hBqgUg8reBCzwURo4qQxauVVoh53G0K3+hNnYIPj
ednaazUURKn3/u3p8vA3g1xe24sHn4eGRGEnOvw3fycfDo/fxX3gLfl3hOS7WslM
37ymRGm3sfg/HVvd6OwAByf+7Ee3VZoHAQbIHTs8Ot9j5+41a4K56+ZU3QJCBM8C
HiNuUPHaO2JqlLQDNOIeyKCaMUS9/Gqp4ijOfMSXbfdKc7UExHFtv3lmwZ3xO4e1
3mcInCYtZLaR7eTZ068HUWQidfdzlflBX0/21wpYQG4n6MlEJ2RHw81n6r/bg38t
8RRrk3sYZfDRufVWrlneTMt6XTFfJCh5YHXEYskKY2TXBjpOHUegDZkQFAdNYEq2
H+pvDX3wQFtNkqqIhHzoQmnJsS+dbUWXqxI96r4r1tPIbuwp5BIda5unl0Zubr0I
OQY3YSwaFwa+Imy1ALs+QuqpGfyqidQxI4QLDIUy1z0x4g+pFyP//N7H4UI/Rsl8
JWyA3tly7mECAOdaIn0Rbro4kcrq2rjyx1qUoLVUd0KWWERp+YuDbscDOyOjdVuX
0dC8Ue5QNdoER6nYNSr0bdeY1bqcmTD7dNylSHJGnXIVPI6zzRO8UWPmwGEF48yR
7qU3lY+DKcnynnihAa4eCm2oruYGyQF9a0s4LSA9qOFF253s6DcX+N0BYmYG2qNo
g84gDvjzkQAUTda4rAB3PDu3RDxYRytGZzv0fuq03SBeSYe/VlH/oP3w99lf8/lE
2bWzml5s3ja5gZYkGWuy2HTFFO5bIDtPHpZS2J/9Wv2QIcPyQiGbPpR7KJPoqvwd
MhkcvDUh/XjWB2vM/vr2E2g5qbvbqduYvEddIjYsZPxNmzdIFDY1Ng/8+67yQ7NS
xexcPjEhDF+5f/JWE+h0pdR7n4HCuJeEc7LJIgMqGFIjrOLrQ1LaAOi6DJPJI0qL
5Dlqowjbt2pfU7cvDAgMt/4Ykw78rDViJu8eGl2wdgVkpqdOjPLWVjdwRJ+1HpDY
9jkBxqZRW6L7Hxu1l5sFpHi7OXVjP4LpIfSw25bDli6v5S/SJQlmtH6ddua9pdjM
lFAMRiHx47sKsjJNfdMz7oe5eE77/Mt4vq6WHPwVBSiloi0iOHzPyt/gTm6K5ZrG
EUyQotJme9W5/rMqyo7ZbM+L98IxZdP4I3y5+0MNmp0tmA7cOv0RflYSL2NCpDBa
tUTTihIdZxqlLU0CU7mc4LywQMR6MbBWDRkn6+3V0sENWpudW6x6h6uNUPtH0aPv
XSHSfALP65oY8iRWLlB/5NDKHEOPKQrQDV/IY3fsum5h9KsR+WSmAMrx/junsT+0
2OPccsE7kcMctz5X/LwBZtxbJulDSkoHA74wgm+9UkgcQshvpJMzkppMJuNYDR3B
DrJxHZKIcQQuEQDsuK9tNeMrRT2z5o4l3RA1Fk93Tsq53r5+b/y2TGBWEwvvHode
eHvUn1q2TH0MZ8YUB84onP9+xemAFxrVOn13cbhePu1HQfG5w6k8RKKx3KlRPx50
ZCMgc56hgV08ly+VcQZYsT0UKvr5QNdCIrmfW3ktM5rFw8SVngHn4cuaGaYdl4VO
7txTWzwoIyoFXtWBMW6vjXJbMyljiSMLT4vIt03ZXf0yCi9Ef+aA8+4p/jqYGRK+
aopT04uvvPBkwmMB4fOIsbwlZIuecYReojyqtbOu1UioBnuFHrry0SVXqdHSBlhb
2N3GKHa6p1vbwpTJh410QdlJAU7Iu3uV7+DJMPl19gB+m7ZW7DIolXbUwDdKgRfN
BSqDuaRQN/McOYQ98+QaVcZwPKOUrDRdIrBa277fEZ7eTarstrleAp3gmvirdOFE
BmNQ9IpYmaDT2UELyUhqE+22X60Wc9LLdOg5xhWytXzbmLOjgB/7BlAIdVBT4bRi
J/y6vQpQwj2JV0q5osWmkKlYg3BvOes55ErzG7omM76D9INZN74/yO49I4UjcUR8
jh1L6cjAiSqBpnW/zqtwIu8DGAWfmaxRv+0edrjjDfEfLNw95cJrkNjGAU74fiic
5tJhy84mcIJpEWWoLswv5CieWAdPcbODtwQULzCBwmpipr97Yp0vSamdgFAKFvjW
f1/4BW8W8CzA9EOf+VE8FuKmHuoPJ2qKT/ta7UbbHqznTuyn8/U7xz5ph3CoLTH+
1q4vv+OPqUcs2HQPdNK4ZbBAdSJJ4KWedVteixZdMS+UXCEe1b/HiC/cRApWFvek
40HcydHjBxJq6ZZnQo6H2QwWo/sRqN/cQWFC1vLBR0faPT1a5fsOpb/iE5bfWFJi
Dlmc+hOu49UbbAYbLVlIoFHne4lhGnCoiA+PES/tOotnkIt/6er195BREGwm4Rh8
smU4+aX4+b5bXS1p2/jlhB9q/jGEjSaff08z+fJXaCuT6DmvLklfsBAwd6xJYnIh
pFS2xitNH44/ayvlN+Z6Q8xR9mjinwbjkoCP6+aO+iIeig5X5bbUUz5q2U8F+T5e
lpPAXRHA++R3PKplRcGuyxTqT1oMhy8ZN6tSfvO3kLQ0BmtbPqm7mqUaqzMf4aC1
ThZ1F0B1i6X4C8WeZLz5i9mkZX3CJh0qNoeR/8HDTNsXALxZVcEi9nzcN6fqvN5W
p2drkpk6C9UJ3ObmAOjNfuRL1DLs4Y0ZgE+0sEHeMUSWobJPAB30D+dIwTghJpnD
JaRRwI4N8UJBoUSQq6dodt7cNnRKuJJbgx5vD3RuhALYNf0mQqJd5z7eXwMiIAbA
GWlUpFB8AFailJWC3BD4qiaMblzC802B1OF0jGPuPiYqOMl9NybQvjGn9e5lYjdS
KLA/0o2GqslAspe06TQ69SyU9PTrS96gD14Prc8KE6FayDEo6/pl4ShZjctbGCSe
rvBpV/48MtptwqLlQK2hIwGg6ZOsPfhyKjHizh/fOfZGWTAYgydjYm3yIXCH/j1i
Qjqp+zIc3GVMcgbUaXvvfLLNSE6CTWxiqP+COn8Yf8a4WWklGTuL30nOLx5GmdIC
mYiO53M/m/3E01kijXSTi9HTITD0h+C2GpXhaZe3slMY28hDyfqnCH2sXlGOv80L
KLxSQV5L4oGqnHOkurjL+DARvTTQaiKV8Y2DhO5RxRPFO3nf/XdSaAFwupASC+/i
Xw5o8+JXdE+d8BAcB6Kky/HpFDMNgTTtIaARECFGoF6JDrjvfO/yCOwfkLApXZND
BRHdn8yj4AF9zP9Bkq2QHBbheiy6Wp2LDeQWZIz8vMenzcfp5orjUUCC1zNLMPo5
NblI/v3InCLhVv032N48frrxP1y6Z6JSGjkXw8127IL/78Nsg/BCqkg91pL8nNh1
IMp8I4z11oz0+ut9K1SPRY/KIzP9hLT2QLuaDoHAVNr0yM3EWl03+daYk0mlUcji
bHgJC1tK9PutTON++YJ5gQOz1iolI9FAjiolpmNqNZlZEAG6PsBvw6JW+uQlLyXS
2q3FipXymAdW3j8eX3+roH0tD+huywx8uxKpu5jqOgYanjhqFeGOPoCuS5Qg6hCm
wj0r6u/ZRcA/dWlRJDuTJjGR+4meC9eYgNVTsjhUOzs7WX4cugUuox1pP1tDe/Bj
VRF2GvPWlbVj13tkn0WCrHVhuiyHfM2TPY/XMgajnZRiwkLZ9bYucdDP0FLpOoBL
PzldqQUCqxZ3u3VyC9usSs21poJqZECvjhJhDRk/nCsuUnJYBQUw0h6hSfFTjXx5
SoSsZsEjZlPWS6wRHUAokCUUIoJCaPObx6NichNaslFv8EyyR5NtN5lH8E8mOZxw
1KUpwTJYUxKHRxzYW338M7V/6BhCEZFGUdBqozF/MLTl/LeC7/5pkxfL3piEtagB
JI0OQ3z3FOHmK75DR5fGwedyxsctBskynS3QbqI18V2oZ8ho31pST/Pf/uqYVhqN
TyATLW6JN6zU2fecIEtmmh/22QZSU4EKVLQ7G2GVK99GLuohgt85NLijD2bu7dVy
suikd8F4fA6ZTYVlln4/OlSt+QKqzLL1KT6bi/V0pasO7UmjKWy7YzVVxD0sqgQ4
IOXLnLkeAq1vV21KpDE1C/omQIDxCffOMiwiRRnpcf2k1L6v+fgOMCZLLevT8E+2
LJQOSYtAHXPUMJpCS8gX7VbWJ8SIDOkuRwO4TmtUjkClrP/a6WSnhAll+4nq1P5j
tPMRAEHNr0jZl2UmW4xrahgZMhIuMA6m0NnViE6PowsbmEdbkwLtQB3l6fkbtRhV
s3iItt1m5usNWMxcwOXemJtM6obde4vvq90UIvYuJ4cEEv/ja+YCUAAb591CgGEB
5g3Eh40+CHxZR+m8GDWSS41uEfv2BEGIz5dizNWHm5FGRFQ3eOHtp2HNuvbxAdJY
tvVrtkMOqDrEx5IGLGqcOiTfE0dV7TtkTwLSNZjUvillEY9mCg9l7Ql7jKIlv+WH
N9kz7RQB4vExFhJABoNXQhedj8agrABe4A1kjLzI80/89NDlysjZCTtxZj7AM2Vq
sSsT/C1rQra1nb3SSAfQYXUyixE316g/rxt9tsn+excQcB+Am9HohgE/5GFpU/Co
c3naQe1Lsbn+KXvIDP35PmdXYuE62VB30NPpiHXYBqYSMUC7iyMOIGhvSwwPoM2S
e2US1gnnCRaBGdTn7PtZhM/8Sb5shT2jo/Cp4EsSurujAPHUFMBiQRtkyUB/d6ni
IO1mP2J6w9nYFoQ3qN5WLAPAQoS6FlfYxBhiyYeh2hc0q/wfXR5vK+IvTRYMWnWt
IpsCngWH808MX/noadfK/6k8FJYCat0ZTz6Yd4h6ZXRYopZ+u9Lrj1+xU9N8SNVj
/1n1JINa5cawBoe6up4l4aF8SBm+/09khIFhmu6jyqBLUYIhz4ODRvOo6Ld+1rWG
YZJOL5a86XWGK4ai5Pa0egzwxr8BcwWU7CyTqc8AG505AsuSJV5Bw3E1qvO+KGkV
bwK0apwrf7oixuEpiedI/MfgG5uIcFZ7xpQ8LaKR5StNnmlLGxpkndr1lKd4BRln
VgpNGdZliR9Tl5GCMkVHloAioewSTiRP8cUvnbXcRltikfjv2Ap4KZ3VkwX0Qgrc
t415nlfKVMROYEGw1HgfoF/pYRH8YBgkZkoP+UneM9mp2ScJ9CzwnhidJRR+Fplt
doKutAuAggNWFPelgM+euspY4UkCmEIEhMvjWwqSmBwbGhGuz4dDdMz43TVqvLKX
ei+17XedFblc78zPXc9ER+cdvTJMYGmycl3znsM12fsllIr5qku0yVkgpdBpvQ7n
0I3f0UFh9P6Dq4EhTaQYJ9cRSbfVeH4t/kT1RgwIcvlNgFCkywGUU+8y/JRgmrM9
l+oQYvIq+zOQbJGodKzvPZ9uB98giwLaN9xmRAlSSW9Reo2AnGNhR0x11D+raLLH
yq77hwTZZ1VkexCrwhKPOGor4o0XVzRvVHe4PmDckIXKXyR0wDwYnQvLQHDrSUUg
JSF/Tw+Pwe0c10hWAdVspukFJBhq8u/9or/W/bcuph88O46vUbtNXtl20GgmAxhi
z2gUFjevLjD8qcFec/J9+2izNvbOOYqO+tSJhpEMsfaBeC9QzAPGDfuK0R4hyewb
1yst2b7usjkUpQ/sUqu43rs5QygHI1CTCTJriqNSFNSXeU1h96B1bH5+TR55K+3i
0jVaA5b3dFVEE4UnLR2bGleo1s3IBKyxwUrp+KYg0y9Lfki5LFelwPFYH+q/pRE8
uGxD0t7EgfhctW6ogwyGUdI3EVqfkrGdbGBSIJbOsUCO778vp+qD8VdqNiGsctY+
w6DADQL7M8Uzfj46d/ULLbKtSiof0+b7waz/RsiPJpSq3QsuUPV9IloaMhdd6/PR
lBmpsHq/CVl4NfvBbt/0IX9KjH3ZxOUicoOE+LiJp/xIdQ7xBpIecbBUdva3LTVN
vhsreUuG7HVWXdjHrvsOyAZk/n/TBjBeDtgOmNxaEm+8IVdSkBEvloeZV/hvs2jY
1O0FpOsZ3nmo2Iew8snhg57mKV3qTRtlk3BYR/o5jKUd8EisH5/A1LlkJWmMa4pe
6JjVYKGChNL2rBqIEq87bmtI3yIKMXt6z4+ghbe9W7HOvUMkpOPN7CEvEvOXfUeI
leDcis3NQte7Mh1boVYzzhIgGzS2is/gzsZhCdUsJVNrtevzd5D3IBFdiBFjymR+
RoK+LlBDMlXBObUfVMmUnah39gJNLq1gzszIO9lnIvUj0+aNYs9v/049mVHiJxNc
Lspwh/mA1DoDEzFzU3VQWVP4msQJgkLU85pmapiUKpVkR6AhbIy5Bo33JzMye/3/
a5qO5/bch72wa+9OM2K+XynXAETkxbSd9qccrKQsVLxuyNArUS6twx+0PoEFMU6Q
OFMsZX3FPSZlwhcB5RVKd13z7pdcGHDltAssLJKf9pSqFoq9GhdSTcb9/hAeynjC
8l6WtWtp+X5oOO2l41OQ0rSVL6EcLuyM17FRYcYYYlmhlf0PuL2Qia6NfRla7V1t
oi3iUHTrwXzqYAO3mhlhkHYmFqDoPolIu5qOBEWRG+IJ3edpvcFqDgQ0CJDCE9zs
oJvcdGzjq9ihM5l9Kdi/QKRankOaOmHDWOoqkaml3JsoPKsmA4neaNSH+BxnhhuM
ch5arecAHRh7DQyybbfFVb1uLI2V0aZz4AVrOTGcPObhEPP+a10ZDSgxt2jKrAL6
UK344SHR2b37IvkOtBSu0E4jm9uin19mI4weBjfUGYkFrl0ZJCOHui24wWjey4ZE
ZpzYi/TXhYZIwd1kxOSap7Ru671O4WAMtgYHF4B5uTWMnaaAI85d/1XUOhZ+WrMG
JP4UhuO9Xp7/qdZx3TmE6mDYUm42PoPB2hENWVSx2l8yvN5Sq+wsku33e7S33lpN
dTWKGYjNgkIXTCl7GxRDrkDv+PjDNFzVs0/JimsFf7MTrz6TztlNmLPAS+saTF0i
nRivcXwlGivCe/6yMDp8G6zf0oRYzu5u+qp7+euec3s3V6t6xs1nGBX0v+ScJqaT
QAkeLwXcilvytNy+FTMCTVsH+jDW1DtqBmGpWKzU6pD6rLRPcV5+CKsY4AlUXgKj
jbUm4y9ByfXafIaB1Jli3o/4qkiMF8Vncv/MkTHAyOqri9Y3iSwEqQzffFlQP7A6
2Ft8brSsE8r8B86NjK8SbMufP3VMh8PRlLwk5YupPbcU2ulN05s50wgwPg+LPwIP
dEkA9W0qoewJrKyAd6axsvkcQUCWvgAGHzvR6uhrBSNg4GXqHTnUNospRNtX7F2u
uH9sOZT7st8pCQmuv6dAHzHvcjbk41A+CCummbExpSWA13ioMYpN1H26st0XHgML
X72z8NNE9jGNWpkVu+lKTe4l1G6NFPo1oaoT3LY4skEeXWCqgwXRpUEgMceaHiCI
X0F29NQhqPHckVJieD04SlRV4LherRoTMkeX4GdmPK2++BZqFQ1lzo9vNooaGhP0
GqlAlDlxHhyTZMTUd04FcGidNuo9TdEnxztcNblYQhO3Q52orWT0j7J/lyqWqiCv
UMVdMyArZUTa9PSM9+rws2s4mX9dikz5maI90PKrkPHtUpQO11pP/VA6F8/nO+u6
jS6kBpUr1GCDbx/JTJJICkUO4l/3b4WxuaDnVP+vf/5ihEUOln7tA2cQx0zhMTpj
1tIbuhDvyy+W0jxTD7ooRr4D1+fyGynUoPqYGk4pSLgWZoASgKdj10Rc1V/p3UDn
+4MIAkMugeZy70xvIGxzwyYrdhJd5C75yPqDbs8OmWneXB52n//3bekDOU28clEn
ksFzsE/vdJIi0uV9Ooi558mzzfnpSKvuvxoF3yu6OJSYn0OZia8dT9tspk9sqbkt
MH4xpBUqCg85hWbNFf4xvpY3Mf8Yx50slIwT+zMr4FSuZ/AGG3/d7PSAczjwZ52r
MlfzQiHEHPZknR/SAZ5OGCnBvtrvc57PMUQJOCMeyEmVbzCltebvBxNt534kHThz
l7qckiEAeHEsEqP77NDCSUI73kwkMgqComn+NuPcV14tM3FB0G+r0RzLDu1CsxKm
Cc+c2hOxXH0NgJnOBpkOvU+TvylSdF1yNVpNFdF8FNXD9FEKwhgxKfxI2XV4pxn9
tFMcZY3fgXCnYFa+WurOcgtBbIMhPIrXXg23snY6nq+hPKVF2KOQZS556buoYhGz
jDGH/P9OHjzUoSiDnrP8K/uyVXkOSzcJTObRVmGK1cwpZouK90r8z/fNAfmbVoSS
hgYob46X8/0x8tFK7+3QyKbVWv71WcZA7KEEqiFniBEtVix594yjrsn6HSWfhAMh
lQ4N3pWMZ+jq3am+GKsQ9OVI9UXFr1daWNlebm/yqExuvlC5aQrL7RD59Kcc4yMQ
Ky6J9NC9t6wQslJn9fbkdwLfpYo/5sQA4bKtla4F9nBqzWn2zcNqLKKzzPuvpCxR
0Az/6G6Ifg0q6g5rGSOtuXwBYSgQG+5DF+oQBO+favwsodVF/U8XVHnAKbtEHWMl
OUr3rk+OvrW2kyPo1lo0IIMYehmDi2l0MXQf3Ox4bu9Nkl6gTTZT/2Nwb3QoPExp
7s6CXIAP+HNaTH0+l9zRxHMDcJHMHkaZ7NEDCtKBsRsOVj56ZSHOIf/9bGUX9lmh
ctg4DjdiAexelJIzWW5eAGhT2IS9rBZ44SpOffC8gkD0ikZ8NZx9nFwDrxuf3OjF
lWXNngCof5zkonBs0BVrjjToh1GKGGFpY0qIujAyq2NWT+QNZ9b72PbOPX/gkwTq
IleC/zaq283Qr5WN68YIac27LtDrvufWmf5CKg74bkiXZ4pQXQPbw+CDTbjlYRnC
Ovu/hmvxhjYYOaFrM5rZJZQfOQWyzsxnJb1nJu+BzOwjRGqVWri1xpSvxTrCTW5/
eu0XcWZdb/cogPB/5vI68XtJlJqHfXr1T7SB2tup9QAj2v4zA3rxbRAFV570azw5
uoFR/HCczFIkPaxBihOtHPL5MYPa2vG/hPZf6FfvkoC6ajQxkjPLoCNHcIfxaB+m
+c/M30NadGSdPaO6QO1Lt9ye2Rqxu/5xDJto4bxs4tiYZvXBBFIYVm5ieCKNPSdX
gWTNtboARm74A0MAA1a2/7EhnZSlnYRN3UNqQhaABX3zaxZvv6Kj+l2Pb8WZSmJV
NpQRcnAFSb0wAKIh9aEJfExQzj7Vp6Va9PnkE7AHDMy+391lS9Y2aj9Wy6MDH7Pw
7ALb2GBHviNKi7xNO503faDYZ8sfCN39qNXC8NHOG6PIEpDaiWPs28FGjhiVMmBs
VMie5V0euQzSHmghLDVD1d7uUK3p2D/E5yf1qpISLoY33y3mkbVohvdYBPaIsc0y
OEHfClrtJx/H+ZhXNqZQBOJy4I9SUv61+c9eYvuHKR8+J3QmwXqTf9LNDTIICrnj
A+yAVrLgxuf3EjiS9V1JLC2bGMfkHA+tUWxC91127sl2Ib9/TNko6Eeateq8YutP
JCYnJJKA4dkZQY8pO519m4HxQ2g/oZlO/kLku7HhX56FsSM5SHi3bnQgATKP0a6L
qu1vrKNbgnAorpXWIi73OlugaMOeGUYbjtqRfj5DoMvKujP+t8syJ9FgsXxEQx0K
ZI8V9bByZLt3VicYNPn1eZpk0jyU3xEBW208Qn6SVhP68IfMYiIRZIfsTR+NHWz3
bGTRa+83+pakDawuNgzfP1Fo8e6GMlx3QrionubupQSdfNQPzr03DhgLngx9BP7F
+waEmepnV6oTBB4Jwkngj+4KTAEWvzwVHo67lllzALgeu8qjDoCQ+D+FnHGaBK2j
vENELUbzmB70yNr8Sa0ykG9f3I2RFDIHTq0I7n13uQ/2AUe1lyQcnfPWPE6UUs8y
z1295xwPxMmb2TH6Z3JB1jPITQi/3krwSy3bHLIxQmX2O1RO9b01I6JxxBR9fvym
0aGkaCowmL+69oHDisbg9BCoJmOMtsOIoaFW90TodW8dQn/507c6vapbrXzA3m/4
jJlLotldAFpm9sfweSV7zkO+um/Rgs3/KR8Iu6+tP6TuDaT43WK5+25QXe4pmkPl
9aczafX2KRCdz2nOrOzo/rPMNSZN7FpAJ1b5WTmcNBjI0zfsKY5ohp7XefuvYmfQ
5t0hWmvcM7GnTcSWmA23T4DpcIEpu76G17fgc5vJM8bl0gnIy1TzrSlAsubGDFza
nF3lcKJxkgOrNhwGCLKV5O3MSl+f0FMFCK6Iy4rXxpckgXsiYH2jnXH+nlHhNjFn
YFwI/GHKIMYGSr0RH1rtxr3xOAvnI7ARBcfrEMNsfCkIyaKO93f+ZPZGHLxG7YdL
uWzqrKLMQBYeOhcDfGiZyAh9XpNmSuPjbH0alp8spY2zMc+1qYfTvtL+nX0uUiRC
wyUpQfNvxaXctUJMYggyX8Rm9BBdQJ9aLzCATnEgyhAS3T7KonpdlXluGWA3ks/Y
2n/QIIM7bwWDfkZVQU1jVWCUQA/gZM1htKOI2wa2ZCi3oRS8eEWVZLloE8MGfjJ+
OXG/POFOBJM7NjnD4T1QmqQj7r+uSDlK4Le0dxa8nYxsMjlG8szXugyGW5ap3/8+
y3iAoiRd9402tdFvIbmWEr3Js+VdHJboAK2529Q0jfHbZGLuPavDj3wRYLyCLjVj
UBTSYfTb2ywpemmaRU6t5038gGwMrN4/0wTQ7JrojCr2SwmFBJM0H1p1pPsRqHBl
02yuhgWVmBGgnelgjwF3GIZVfM94aX6IMM9A0KtR2xCycnl5Vv42shi8UwdQawUo
OijU7eKTBU3v+7gPsqq3ch/WS40oSncfCLISaUKKBZPMB2JEQT9MtQtCNLnp5xn9
ArTc63O7bQhRv/EpCCy230W5/y2oViPGU6Z//9A+Rt/GDWGPMzKJ7IgR05nf+Ctg
FMhUdKjGIK2xbIgQlyj46fDI/hir8Ix/PKzA8GQ+IxFVUMSMK+OFiyhrWvlUPl5l
/HfDxR7vwEis1VKI7AKkKN2wgz+6MfsBy3Wb3s7j4kvr+GK0aWevldMRKtAti9gw
Ch+T6b5lMRQ/+3ZNsmPTsqqh8yH6BtmVCSuNWhnWB8aYIW6fB2puWZauo6+ol5KP
8YtVKYHpXPCLACRMvON83jEGNAmShQNBL5Xmq+RBUlc3iURlRkQQY/h1kA+ANSKQ
Tw8YVRPzcwPgA3FjrfqebH3zTzTxb2sXroJsZJCwNXczJSG7wc6RKvzfvrpN5Szs
gjVs41nu2DPPTv5fm69Fy09mbR8JkZ0khE5HhtMApMffwH4g7wPHWXGb6D0yQBwS
PltElFkQykW+sNB98ZhN0xnHyMRbDBT58x7Xq7e2BJJXjHmfLF15/jgL68Uwd2Tl
C9ovmrUyn5gS9JvLrLHoHOoJNze85jQ/j4UvXX5qDPNRbx2SO3xt6i8baP3KFvN0
Su7dx4GtdO/SqSIPQQ4Bv6PuJY9kbOGGruv1J16Kcnog9jDUZDtIW6EcJynVXLLr
IZFC+VhqJsvjZRRmDvYP4kaLmVD1/cEH2XI0d2hz/j8Wr87OHTeHmFChwW1NTRAu
YA27cmgBblyqqmWWoPjjxqCDa/xuj+7teJxLZt3Hz6Hb148EeunLJe8PYBlopelJ
tv4I/U6Zc315O/yWdpTKWOU7ZLxT9liS/5/jgHEdP1834NQferCglsVKmykSgwtg
RK37PXaLvS/lc0j3J+aG8IIujHg3rIE1ZDWUhjkx9XmY4Ohu71Ip2qtKZjJ/eG6v
hYjYArrcNDAWVsJe1hlMfLdpgxuwO8cim7BcbPyWV15SRsM/18ey5E2ZMfTWtbGc
XKzGzq6BZ7KaZ3q80cP7mmjaxpi3Z7Mwn1kdjZhQkyQaZ9sb29BQpHaRq+bxYGQj
ftlzyIJOvL+CpyhXWIM87t13dRsO9Y2kZBAv8MQJpDCPlxRVOqD1QuBvE7C3yBxM
ppxVzwxwripxf2ZcT8RMdmcDBKv/rUag6XjHHjeis7uSwAJSVRDxDuP5Siu2Y/G0
j7ryxNkE6q2UzIhiO+ZWISsobKi1a2COKC9DSOrRtq1ndWQMHs0h6kdfltv6qpYe
0glAYLblmBETmV9gxjMfJR7sr+PCdhKd/ECn+Al/CIUQD35NU0iInbMFmVVxrsxm
Z2v23Pq7tfhMIAJoCraBC5YA9IRxmjs6zlPLwmy1KZOB3hmstfYCJka7jZ+TYkdr
lxqlaUfL/RCDVbpTyBrrjWo2df73fp1lKgq6ojG3+B1QKgyx2MY7rcEEr3oE4Jha
/y897MfLplIZDh1rqY7D9IGyKEXkz+jrBuBzZnOy0bPXhAVlmeDWq3A8rCRYHUM+
aq9jgxq3agJMO8Yj1F0iLmmYB9rD0nCZiJrqiu9AABZCahk7PgGqAFJeM5Elt+pP
D4/8Cvd2zwlBw/p/BblkqNGLmMxPrnfq6pCFhXMkgd+1nuyi3fch+qeuBC/biht1
IN+G5OivNIkCmOI76AtcZAUl/Y5Pg5KAp0LArv57RXZsyCsahOvD2QXAwL5LmQN9
3JjtOZMnPGwgpL6dV4VIbZ0yRmxC5m51XmeRymt2APdPInLVguZfDaLgpgx3ZFtF
j/uAwgF02x3gKPVWtIiSuMaG1OGBXZZiVi+uotPN4kMExy5IrNCXVBT8LBjyDktC
UHRkmBTHatGTVnuxMJqwudzijdFP7GhIp8W9J7Wfh8RXlRTdy7h0Ukiy22x93PsZ
JTjItGnc0G9EOkBfVZFSvf6rGZ6EwpGbt2seHAvGUlDzJ48Bdcrhe6Hs0rz8sCBL
uWt8JGhca259deUYQRJWx0Aoi3olBEIKLhlL38edeIUvD5O1/TZ0Inj7dw5oRvrs
jVB65dRUT7GoQJ1Su58ahST5NRClS+AVrPbJlhKo/v2EDcahdxyvmoyz4k8le1oD
25ymwrCCAp6JJ/nZQKJJI4PERmPaewanZllJ3EAf3INEU41bfzkJcyKlHDSctX8R
qi/mj9QsOefSP8smrI2Z+HVipSwDD1y5DfxIuhWeNBzrPJR/GV2b5/76qp5D7+A8
UrYHbJ94w0yTqRlcHaLFicEx2pZ/x+8BChC/rzBxNZvcetoi2vRO/TA3khx/nAFe
oEnrTlRnYPsNc+xd8vHAKnVPiJ2m5JjzfQ/zRubFG2HRCLXkCK7V3RbVfmMaB0SP
FPxUxacVMIbBWuuqf66cG54wbUBpZsvfwmiOGYty5gqU2+GJvA6Qn0DnODLrSMsj
bW4YE92UvrVs/4LwDOmqre7bFK4AkjSy6ZoyDYbfLiF0DtCrNIPtruSSug234yAp
2w/A83SsiltaUG3MaLgHIEuFoYIorgXbW7eNFxkt7Aq8qAgmSKZah18rjGtGIEnk
hszBj12wMDk/AbKk4zI43GGp8PnJatCQCwcpLFaOFOuuw59yQ8P5b1SbXtSicGK1
mjaBf8y11tlItdIm3wLUmaCPBvxWGNp9MG9DJp5XM4wnQHWNZbirU+Y2TFvG3Jrt
l/jfhGJa7fUUEeMRxNx4mblXNanL+ndLFC+d1bag3Nwf1Z0ieNEgMkcGgxH6kaVx
wVaRh9soS1gcsq+xmAr6N9IQ80OwFPKUdVCwQ3t6P2XsPsVbR0zj+E3EOaGsyF5v
unhTcmYc2iEuyfl5YONZCNBTIoib71emKQnFzL358rFhncws7mVuXe+9IYSwhfdI
Y0Btv+Qku3RdH5yTkqy+yP4hyMEwSJmGozYDBOw3Vs5QhUn1Ykfu+14ye1GFDz2q
5zgGYdiJ1VG4p4gZ3QwKtVbP6nbLYO12I2YIxgCBuzOf8ExyQlMv1XWKVRMko7CO
pHXESu3PurIvs+CJs6aClvN06KbJbXOIaqXRkoEiTjd/JyJA+kpRtUUdTGjjOKGV
Fj6cDbN6wYNwmHLtOunuAhZ0EqOxYOwBXuw+uspgS9WjuJmTwiNm7xZeFvwvHZXV
ecpKlDcC9hg9YYYao5RPGs3c0sUbr0yHABKTMohb4LGZzikCnP5hfmoLaGr9HEwB
sewcIOSDcJnyYuFl2AOFXsg5ygmIJWU0Wm5iOeQpyFCCbftMFcjb6jk1HuOr4zOV
WmFN9ddFtrYS1nSKVh4vpMqodMMYxqiJ/f4BFE9YOdL4CrH45sGeJQA9ePemLKWO
xTr7EB6RyfEu6dVKuAu/5NzhUzLX4xdp7oodUuluroRKjkVSg818dQb1bNjAbG52
X/AEBkARVCjjt6nBbiFq/BBeqjcwUz48omyrbWhI+6KPcdRwM/L0WikEr3fF2dH1
GFPPxfjL+qOuRA9DE0YHq9dm5O5IuwM/0y8cJ7VXRAv0Yebbx7UDqXbl0wlPdeWl
E4G9qN6ct6oSx821OLbQocK2bsqACULbDAFSCXi/+1rK6PzHY0xtRvzOuEqmQ1fQ
uETa+L+0XLeasc+E5oSF9Ieq3RmpN8k/+iGgeghZrmjaFmLHepf9EdFXJOiY5WsI
Bn6tv+6TpQqAXxafR/X/SY2hZKKXWsOEXTR/7E0dOLlBzNkk6/4MBL3sQrBLCliV
Nwqufiu6cq8SdUv45T4u+fu54Pf4/lqRit7XR9qNY0+Nw7iHj+9Os42z99a/3HNx
rB817gPpKLRDhyr4nMVDCkp7uW0GFV1GeLA2EMDA/1MTDjxi7cWRLian4OkuUzdM
rrwU+2JNGuYjCxrpF9bRid+f7cPaz43gsN11qdMMREzcAnJVgINhmrmptimI4JRO
ZAUrHHoigh98AnlkpC9btVhuMFMuM9neRNq8XlpUBAkyDlkmH2qWHl6Js/epbPOk
5fbszLd4DkFc4PS+XVnRqFrzuT4DvajOn9XhVpLXi/vu2hqZFJQtyHA3CYZ9YVF/
IpJ7CWuPQM/HyhHZqo6GvhRK+78O8Wg1SSSKSkg072V4sN22LJzt+/TJU0kE2SQG
oy9RoHNvFXRb2dBsMJV5G3R7hzU0DWQ7mKiGqPU9obY8vbm1+j2nS8rGcW1IHrPT
OgGNvT/MnSl1+LoO1QSdeRz9+smC1dlnDf8D2E1JI09aAD+yUH93Jb+hNh/Qqs64
NrbHCmOwPzP2yTjG/WXHQL3wHCs8wzgFBJRjWO1amctbZRs2SZQRjUqA7iZ6LHRP
SsBZIjEKHGoFobKpnPyKDUr3eNtynAjTFPBbS/9WvvxWuP9uUQzZgUXaqksrJHZV
tub0yKLe9vEWjOPGSe5t8uYbF51H9B9+QCjbMpvUuqyhD3mdOMd9S3pUL+JprmGB
B/kPXXVJLg/gqd6ZBwmxsQ7BTklPySV4VC3OaEntG2qgdbHEZRBgR6fd45F4rr0s
6WvmOYqyd3fFCx4Y3GBjAgQGt1clysVHfcoen7rjaAjQFW6McAtwPVVrg06oc7hf
E5Vmh6ICk6/3jQ1Wuf9McWM59s7EsNQ6dU26bsa+JNAy70vQ+BOcAUmSO+7p8wZ2
zxXDra2QFWZawL2eMiHXHtDDSfCAtO+tw3ZJCZC2VdoQhzElz1rwEp3qEIrNu4vV
ZNYJhbjUhYHyvNQlDyPClg5PsuG45apNIOt65n0Fg6W1lnWtsvKFWnCkRIrOL0dm
LkMwG4+WQ64ra6e3i+iBBxJgeu8LiVO3o6pn4ZYaxqBQUXg+8D14dOclm1J4QkT0
LnKd9LqicrVy3+9GRRILZS3DYM+PsH9FWFfYIQnX4oSQ6aCC/BgFVm8AGjuif/lp
61HOy7P0/RwYDee+AkQHMUeggbJ6GLdXfhM/uyfWjd5zKDips2CwuOqB31itK2v0
IwHSIjJFyeEiXlZqdojjLfbId1RUsnusZtaoWik/BMOnVh+vlt8iq1yhG3Vc1Toq
mnWAG/isvbjUGy0x73P0ZruwU37tPcMSvGD1kwAVZ1+UquzxUYnss/gRjoMM1/9r
g2KQScclT4zTdtUeF9DRdrRqfTSbDj2rWp0GvYtJqcduBPHsYX7nd5tNcV7s0xSc
WIDxEUYdHUPFYvILNNXhCfryVx6psZ4XwrY9qR3bxTaSee2h91R2gE4082sBSSgo
N+h/SyvaiQsNC35VANuoJAgNzfBvZQJm4YacDN27X9vhftukXZ84DGbeQZV8s7QS
EFWS2aKlFYBadEYyxPRcTLwv4NCs29F5nLlVmt9JWKDlKfg4Ux/XXPrxPEt60iHF
4hsXMXagpWekNIf8HGB3DJYAS8qo9Xepp/79UuJeJthnbuL2HKoTTf6ep59ndAoy
4kUuarrPtcMIQEpd4E/6X9JLLT0iaGSY1SrbElCYb/UvuhUsTbrHj2S4qQpw2RQ1
9lYLO5f/Qo79D0SD3bW6TJZIUodyOC9hvm9mQ0SbRX2CnnAapffdpFOnOjVdFir2
EF1DS1nSefuVAtiU3vXG9+l/ylp1H5mC1omRJxtYF9uqDIuV9N2IgNUWISNlCujR
exW6q4CNnI651fchPPKHraLOfsXRsDtpSGaoscx8qLjfIvRmaF0Knil50xs/R4FG
PjRx/no0d+XTL8mnl2A5qzzxa26b+ljkHPpdT8fWb/Hly7aX2bLeu/CMQBkb7nlb
Y3EZ1IdgWQPYVW0hmxas5qPN5oYIG6RX7HlX25Zq1AvxH5p3+iwGYzE7wJOQQmXG
5+u8rFXdw7s1S4aJQUWoF3FLWG8DaWn3fd554lEwdFZMoAfI1dBJv89CKQmc/eh4
wybj+rvDG8yXYA47+0w3PICvFHfqLjcKzGZi/VjTfBJCl2X/KipwkMAuJv4mKT9G
U86dHKEsaZxuGGTjNehBeQN9YB8VZ/oVRx5ep7Fq1+zMEQe8yqJd4/TUIfqiD0yS
XGz/d6kaslPNe/KE7QbMbWb0VxG/W1LlIXEM73idSR1CiG1HiJFLm255vVQTY/ll
MT3zhntW1dADD08iGPFTYaGb++qhlbgjK5EwUJlsr9KeBaXPiCJvoZiDXUy/2i+I
/oYLcHVt0LG0DoPKw5JyF6cZz9Z4CoIFqE2226T5FlMQdi4JmkfWcYBEfAuHseB8
UIF2tJHuZVNcZ6uSiTepDFfDPo6dYV3CpSl+fPa+3MzR+QV4cDz686eOELx5TEcE
wOj+QAU8fiqvTmZoGXHpVZyK31UqZvc+QGzAiCE91dbSjKaL4H9Dv1I1UUGJiulj
E+ErgJ5L/sjqKSv6V4D3EUolj/lq3DSVziOKGJcqLT04Ti3RHNEJ5uxDm8cL94+X
8sb+qHS5L5D7xLgYX64IH0ZHG+SB/J1ePxUH4cZZg7aVF7iUqUVcORp5+O0Mwq0R
hQWQxiZEriXT8l8AeWeA6wyXBEIcFm0JZ8HynoAGYZKMbIcICSCG1cBBWqLvS+6L
YOftqhAuuGztyNM9UdtdRfH+nIjyek+UFLjboY1EbwVTmQQ3pVNTD0WIUE9wQTb8
flhSFmkxbmdeeDdP/ycIkrhd/v2DkvcBT1o46qIxBzWpYfTFSAP1NHy0zz/K4o5V
tIuHsj3yEAR3fRrvDgeHjgujCucWf/HApu9F3cV9o1szHU86x9lm5tmLojPT9rDw
wyENLwuH9Nbj/t/5oU0EFrwKmw57R9aEWJksKUHSLodG//bnhmtpeDlZqZY/lMLv
7/1RMNT532mHx5472Ejy4YgqxwylrEcUby/Rxo18CqV2R641qHJvaGytIp+h948/
HPc4TjmU4UMslF+cXOlH7+M+cGWZ2I8S9S3EyXYP7igVJvrjc0xEe43hbkW/2EZg
CFfNghszy2lhloPm8IZn1cD/w1G/pELNdoJIhOHs5yPvc2LvMPCbJXBKe7InberT
1kMKb4JVYoZuJeJuWqytHZViZMOOvoo2yr8FMQ7t6JFPDDuFFXmlryJvlDsA3lZG
juE79ekRIJk/77k6GYKyGG+nOnQy4LlmJZxvwsoTAL3VZhGuRbuwMBG/qoVOHJYo
LGI+vfu8lBrn3Vi1qKtvW2BXumkrIy3MUMMEqlMaiQfocqh8MJjh08gtn/iy7jCT
xK+1XkjzltZgfhJDDIiCKdE/H94QL5SaulSdT74a+ewxUZZ+/dKMgAgyrEUc9eqz
YtjGexnePjgsToq6cHbxwiMrEaiiTE0NkL4OSOoqAU8GMpVDWXY/PdtWlPNiRgyH
V1tpo+H6KtH1kDBzXHq6kGWG7OSR00U8TNaKTKVCCI5Bddeu5uMbyKSbL2Fy8RXF
oGzREfKZfHKmPV66a6NIrQZA88I1k3Avj3bq2Fur9/PJOAfzXRllEhCicGatDBMw
3+A3a+VfOjnjCmdGMyMR1vAfWZWwVitliEZYfrTZ+0fC2B6FpeBSN9vjT+tHUMKR
yWLqT/dPECOSlN5X1Uyq5lBetgCE8OR3hzVA594UIi6G5+kF4g4A9QWERnG6cWF/
wsJx+U5JTIJtE2FtIts3CyaLm0GWrR9oaRB6QHbvIMLsfzIj+g+AQhj8CXAjDrCe
Bs3WCMso0rhi5sATWTkR8MzQCWJ/IMvl0N68SkTbtmNAU/S6+3AM02A+dAlG+gwd
csPlu0xZ8ld97Qrq3lgCSDYspAPixUpSS6jK6HBKzSqVTVJY6QqFAvFAgN79xOrA
REAz7IxwTFGtfvLnyh2eRbLLJL/aO+NuRKNtk+Ij583/EGZrfjGvfzyA3ZHOyj+9
3YnvktuPfKOgbMQJXhL30G5gqoAnRhE7Jgw3CyIunf+78nb2zSv9pjmVRBKHGnMm
9lr9v4TvVTGbntnFaXVqgB6n8uI6hmNwSm6Yqct8sSNGDafNBJJo5K7uRBTKLX/j
bWJfB70D7u/2KogvL4uZlIq3+8LeCyW31NAcI9Y50svDiALbmTsXQanIKW4Mip62
6UX/01t/XHCzzkkCVJ64QccIcfJW2D7hFx933/Cs8BFzxgyjmPO9ShZNkPPcEtc3
2psMXJfADCBaO3vn7tlkVCHsBnRv5vRUizT4x7mnyTHHLWYy/25zfFt+8uTuLMd+
3YK2YZ8n+1OHBNDyAaDeChdUUsXoPBUoHcyGSlMGB+hIgA+2QiTM56b1W+UsMy8h
OJifjGSwlpa41E3ZEROBpqyOqzTEky8PNzGxtaNjk2DX1QUTw6dnLBuP4VJOQLKA
DgDjktMvQJFkS1s3OZyVtkdFRkfCQNbs9BBF8QSJ1LvOESWEGysfgtkBZmLbwGVB
FpAHEam34+pGguBG9fzTudMgt7F0vmay8z8Nn+DJr+40NWn918RJIdfE8m6P8FvN
6CMQYJYYNmatuzBSPpDJtOotydwAlKxc1SORbSrshMf1AWSCm4FTqiQkeZ3KUZdF
KrCoZyY6Gv9lwPrabb0sHSvg9iDTW5LZizCqsHN4rtY9GelxWrcVUSMqZtzKRJJr
Ax5a9L9IdwdebzVjJ5S45BkZcLcss8lS2FaDn74My2X5QaeXTKgtwLl+mcCIJ2N0
MtJNeAJXv6yAc6Bbgj7Igl9SNGI1Sdr/s789gAJlH99SpfSmMEwWoinXJRwTQflT
Y7tQQQsYuXov1GwhOzRSM7ll0bpIuKJzjlIDg5l1Wf+cDUvI6TuXdj841dshMyss
Y8RQGOkeaHCd6+Cb/YBYMZtOlj27aBlc12NDl+eov16XnPeqzWnPztyaIKrraj0H
+q8SqER8bIVhIlbvK7djlRjOlTh18rfZEWpKoi6vqQMmtzRwEqd6ZJSGZSHP89G8
+1Cs0Wq3cSujPxXkefOI8i+6RCgu0dGL1oCcvhLm8ekr9mARHrMK5Xo5tx8iiGhQ
MUklVBuiwHW69xtAbQUXQpm+83L1/vj6HmZnZ81B8qF62upMNCo3qp681vIsHVyf
jwuIEZblSwtnhieD76enuIDdSdb+lei93jD+86Ky+k1LB6yubwLWT/cVZWA0T/W8
uJOLZXnCfh5r8e7jftrQMtGkHC+hv+ro1aMU2esB/sV68k2OvT/EiOESlb+RrEoj
v6DduC0Wxx664wwVmpp/osJpBhCPpxMNUxQZccrfaNm8Sn4JV5ZU1dWMjQT3BQyo
y3UqBV4ip3u8dPUUDaB91kAXBNpTv9LKO1F6uIQTIrPDtWgpe3qX5XC/DLUrCU18
fgxT4ybTB+F4g+lgSvC6Ezh0iom/ukv0RhhJ8mUBixYEDXnMWYSyd0sKcnwzVARt
ykUZWqcPCKrHsHEiD0UNMvxXjq/Q80LKJxIkA5T7p8k33s/wTLO39m5pFk6lwCqt
YioskeNb366zmQup4zmVRq2tvCZK9efKOPxSHSZtmMGi15vyTf9+oxjd/HJ+zotl
1NBNnxftd/52kQFSHCgNOhRLdCN6FwDoR/p11Hms0M+E40+5Rizqj16/XLb3wmsj
XTKN8To/bA8lOqZMd7lc/Ajlx9Meg6+N5IVu7tP+j/zIcAMu1fpXQb7k45J5MPyz
4BPPLaqTdqrit/LQaNMSFD5cngE37HpddG5bp9A6oJAOpq2UWnGcPkJ30YCYuFKG
6gZGJPPF9GWgYq2bMjSFpMvha42Gm5WQvhVvmTF4Y0X7mzdqOAaicnRWdeLZ223o
Xko2ymxrIrkJUmhV/Y6fIj0r4/G91qn5QVx5Lp1KpVlPirLA+fig65Gr7oyF745Q
qiLnI+8TqYd280ldgBOSBCRzoOYPxUNlAI30yK/jBRdfMjQIf6WU7y69yHck7OSj
qv55whTPSbl5jTlcQAzdkjBaYEJ57w76Caza+8EuCD9nZ/XgbDwNrNqH/0b7g+D1
7V0RfeZzksVeO/VRhH7rZcEtZpJq1hDhLs3vS5XBErKQIC2176DUr95lgL98NOZR
ZlOpnQAmWH36MRCzMsyIrBbNRurWwiGmRHoOu5oFFfzq+IjJKENkwUWCo+q1M1DX
oOwTdXlmn+q4LfSn9aIOd2V8lO5lnILpTEkdE3HWWgG44jFvySv+a+2RnOcaIgl4
dVOxQi29I237673AldN73RFZwAuj/DyHx9nPVvCUAJj0d/pqdNGxjNrOpYM8/ckK
I5K2Ilm0svxCh3Toh9Ox6LdnkehWyer8bDqXgWTHgnA24jAZkqzna5vP2jYL0PEe
qeuiuQy7nxwfXo3zxFwAO21nanaPmoi9ZCcA2vhN6AlDR8o6cCAJm2AIBhHu+DEy
OnYyavlLwPWue/S8VPaRVuqyy3KWL3Vj814BaKEp3XtXXO4eta+oAhpguOa6lXOz
odQs5CYkiyK/afsh6IQSu3UsXAhbfs6MPMnj3aqcsX9CJgt8dFHAUjAMHHZu+U1S
+vCaa4lnRiEFDZYpAEbeMvQG3Y3lYwXlcCW72UOX7wuaJySF1MVO27TyjI2D7+su
25kLrGAqQBLQRcPoVCsGLV+CC9trMhpd0PLbsd2T99J5vEL+mp+XX6ZkOpEhHfN+
x/rN4vouhGGHkRr3H++snDryuW98KY5ABRzn5FsOndEyoeYsDFhzH9um9U7QgpfK
9n6yNtRW9eiiUFY0qWrClk/ZRMbplEBitCsantJZMky5xYUhZ+5YDv1Y0BH8qINv
r96GWSKOMNEcgmV3f2lL9uqB8CQhErkUPPOTZm1b24zZqlTnbref9MTXnY95WPPs
Zjza4waaP0YNx0qq8eSYxhVHZ36zuaMS6BCK6B3nrXnSgTNZrwHk1lo9BiILeo42
4tGMrdiQ18p5q+j/YS1U+CpmeJsv+uqHet0v4vsAaAxsq4ZjXeSM4n5aluW/u+vN
5mm9oxMf7W6tS8/h7tGp+05Rz18rcpxlnMeZF4MuDcSedK67PnfQRj0EhTUwoPbd
jkB8LkDHYYJvMX4wWlRMb3hVZgepqmXggI2ayRJVJ7NDLy1ZyKAtQ5X+uQMeo4sJ
x1UU8vleHZfNfEvrZR4ZFybnzNNqiUFaOxcUamSd2BsZPINy6PTMKPXKgPf8pijK
4WH7evo3M+41XjyfBbbT3KStrHMYjQNBlKfa4DSdpSGrSPdLvIO9u9gRdbdKLDwq
TdkYb3Aqxww1k3OwCKsaNryuCkEkvgmf37c8ShCTyRPl8/AuM1ohVMCDvG94Jmic
hxnQPmrzL1M24ATdCjcjSU7jGNeyt4RXM2T7gpDJGafdv/ZKwa00/KSQYbnUqp8r
cysVjeG5QbwTMHcYqhvI3oS9Rk04kq9lOpHSFNRXFh8+cvRG4G8GnELexNMYuSly
NrGCkkSmqWTsRqNrb0NAzIPZ2dCc2maSrl7qcCh9tBRMlBoHhtfNiMtmF21MXmkA
4ksldCWcwZlU4ur0rII+0tkKCbTSc38FhmZ0B029U8Id8nP+CtTksbUcjQqtLHtb
BmBg9px5F7hSv0fvzVt9+OhluNeiazsTN+d2gGpGcWXM7CUFL1+J29fa183ljjN+
gENR4g+p3/XLJ7QSvc6bhcHWx/ZNh6oRc9jAdPN01W0Ckr2ZjgD90QYeN5jzTKKI
cNrTfhLNngoL7TcstZMUhpGvG5LG+3/AwD/2e/z5kjJuIRZLlX1zUSYLlYvTWxEc
CW/2TQZIQ6EQ41dTs5n3d3k1JbWoS/g7NuZZ4rU7T9i+aVVhshCgZgtlnkq0VEVc
iN4bEDogdiMS39JIftsJd0evCGpm0bbVN8NLKN7xplphjMVB6k17cPCU4UADbZ4Q
5KHMuM01J8QVS3wWAXIu1vncZl5ujPp+v9vwVHp6w/KcVLi40JcDt92oyYzNoR0w
jdgqhTlBAkYYLqJCkoPaGsCfWQDCVTZBnNIxKA1Et1Y3eWLvztWczh/I+iEZbxyR
elOG84YovgX3BYxqhqMb66TCtYZL9VCzEYfrZRCEtBRdFjHcRrx96us3Toj9o8Mw
JxRbUYGJq9Jdiz0Yz0677pgweIJbwE3Ap8QlcZYgHyNG48Jr08vdwZQc3wwMH0rT
MHaTTfF+4HT72d0tXJpN29MBQgPbhxQIlnP2vpYiKET0Btlvykvy6od0W7S3n+89
ei7uXTZcPDixVycdYVgShaya1m2F8iOLR5gro04Vzt9A0o1ICuGDCHJKAu7P89RS
4HQ/mJ/xUdc3DQeBIqQGNQ+AAgG9NPk9anxJ9O4NSRpYKl0KbNNZsfIjzfhX4ITG
pncneGBkaGCp1xIAM+IUP5JO6DXqS2eyn0H0Vr4lQooKjK8KGGHykUeBWkAsbCk1
/s5zs4w7A0WzxUCCU7cxhUOxq38YSIcJwoqGjb91av5uozAk4NPrzDx3CoEQYvHw
I5H4iRzHGKnuHuzdQ9Ogb+83/u7KQMwwWMQoTQm4MG09z1kSIyBbM0qAVT0mn29n
QQCT1bAGRE4gbcn8J+GfgqocDqKLm+YMJznCV/kcBD1URueul1gFJ+JTzfZ4aCB7
Tn/9A+MOB21DkXyF6h4Ev/912MY/e0ZJ8XIsDqfIT8ehiDcqe/IHbCV1WSl+E+mh
JSwQkbZyZYP1tJZz6V8GI8h7n+o6nQfDbk1jamzutWI4O1Vr8M9OhNzLDuY/jwCL
uJwZzjASyNQ9fRkvQ5XGpXXL4gZNq5aDnPP6cCWYwFPuAAEMS+ZpozbOFMSF8oxg
WUd/9Z3qo2MnuH7UzVB9SC6Z/NN4qjNopUCUaEZ4+NpLVEcF7erRgtw3RhVo8EZN
fX7YuIpoSAfsuAHdi94iTySo528MYC8wArPoFT78JeN0jkAelu7cHmWTdsvs+SNb
ZAPqQ282hXluKzBTjnO1A3n+JtyGzh5FPpilEfyQ6zgTYk6rw6jgnnyDU2Rzslnj
Ri9ghU5EoCKERboNesMwUeVu3QM0w3KF46QP1QL2CGYOn9hlSGUuhonP3JfxDjWo
PDjLIUS5yaR3IeEO5P/igbhO+LXybe0DB7pGT2gaKzNuZLTnAPviu0RkN6oY7aOX
atJa6Znd1/sOA6LtVXdHGgUOLqEux62uUaWmMvtUbzBeG0Vsh1c86WX/aBuDuouy
lr5p9Kn7teia3M8almkwRiCIrvNLEDUI6h300RAdkUtoVAAMN/rnmW/3PCBcBSB8
zgon/RQmkhrTiyUX4w+rx0d4SZIl+aIhlheKlg302YJ13kycTixcH6/JngehXlKW
0mnHVuFzZgPpCFXBeUQygkhgCfpHcBmhW/nBnJhE9jt0HmrVyCv2aZua5xhlFJ9Z
rtj6ihdZAcyX0rXkAgt9z0zJBclhWyjCqTRA67uG2RMjCiiOVoFM/susOakBlIiZ
nOrHuzb7mplXop7DlTiB1u0X1JNZrCkoiJaMWuyIInwLu4x7Qkg+acw7c5A2mb0F
tiwsAwDS1sCtSuZYXtWvI5AaR7w8TJuosTZdCxQgNhmweqA/ztzGJfA0QSWGebY0
8G2dhRxTozd3PVZbDmexnreNhse1LNgpe+RlvvgAWnSusUgn7IF0RpwvPOPwq43U
p6hrml3SH6Rec0wdCU801fr/T5KNFu408ce5VcLpoPKMebdGGJ/2ebFdRPFPlEDt
/Saz6QIGPG71IGH2tauji+K0RV4jtjhU+eXADiud3/bbfZ835sevx3z5BkdpuuQt
+sDDURR05WkPU7QqzvtsfjwZU65dYy+82ii5G/dr252jahGg206n9JdjtkXPP+SN
wEpowp0ecYgKM0zW8Ob8dHpN9jyAXrvC7aG9v5Qxi+dRXunb1UyjxODeyebzeTln
q42LeJQ1uUisIbe0I5walpFfpiNEircBqln/1kJ8eR3yIRKLp3fgTsLBeuSPp825
5rzWMwv4fPJVuM2CgVm3qZUDZcof1lNKp2PTZ/Df4AqatEcVh5Dx3ZCN599tIppy
Sx5ucVUrHBjrAHGvc31+RuCseHNlHkPhOnNiidm22HSxhcXBgOSaB0djIncOnvlM
HWJDl+vmq5m1SOL+r0wFwlRgIHSbUA4Deysxp88yoY1rhhNHnUPr2znkpGk2+ugb
sxbecm+n7ywnTjLcy+K7n3c8szQt+75Nu7NROWKrP27qNdocsBZRI/TGVHIlKolW
lKR8mEPwYyg8jy0paaLw9jyY/45R+bpTV4hSYjULUryBZ8t2EsO6fMGy+WK7FIOL
lviPd1G4H3OD9On9k3xkc0nPrqtpOluoCuL+H2W+wdyCj80wwGfprbQov6kSNLiP
eZZgVoNjjaF4oGNxgiOuHgL1ohrgsraXltbGnjd7yX/56zAADuozBja2O7rSLtOV
uMqvmk0gBCDYQ9ichNRJde09egJ6pX+ArsCjYYjW7BU7hrTkcEsgpE4HyR8w24Ca
Y9uCHSepbmWJkOCxALtnMmZrUG5WLOMac+nZqXW6f6Sw7MB5slVP9IXFyKVVip3c
wUonmiWTmY28/H2ZbFfFxUxYDE3wJpFhFEwXA6r+rpjxZ+AupxHzagcCSn2pKEhw
p2Fi1feGemAvgfzrf5gYjckEuNVkOCX7TXNDyUHK3c763U388ArUZU16fOPxkPA1
17d9VLoRwqKm4QXgxEBBHfQoJQXB/hO64kJ3ENAChqw63u2orioPYKbfaxbyZDaI
gvnYUgaPazBlGCEqH2vMkq5vwHzkzrBNInzSeGQImNY2HZlFp2ItpmhqfyNT1er3
j5QrdA8YZQ8J96+NI93JEi75zb6lmxoEzAAQs1ki4mCXwqlMT48istQVHVuDcF6j
dnDl6boJgokrS+TbB44R1J0FbXWnVhBwnaxH3D+utY58tqp2cEGT1C24NVzEfIrU
DPzIz5R6pct39Moodx/j89L/RkQ8VfI1Tn8eC+x2+pZN4nL81iPgwOeL82Tk6juW
cqY9id5X0ynw858l99uFOLmNcre3QG5j6FzISVQLJVIxP8y6Z6thF8LNe17zkTPd
J4/qd7o7J55FMvHxsjH/S6g9AmyLUUr1udbdCpISSWwnixos20QEbv+9Xb5U6klY
fPqcpQOvNU+i0CDvbUIa3LncrLPWZdk7ZcqcmOYRdr/q/qP9oDNp4bUemyexivMg
ddeadb4Iy+J411tyYY+n6sFzoCLg0Drxqb1lwc8UI65CAsnwifdbsCBf8Vqnkf4G
HoXALAPz0jihntalgCbXQSVKqXm0F/ZXYfN/FWhEhccw4EJ00/oYB8XsJH5KmrTU
6rfTrLnU1tOML0N1FOmnyeU0k4yOPf8ki8APDDMYKhdWSL4lXPHQUcZxUKSJmKf7
meXxgP5w+cqtubyxzqEIr4OUuwDBCV8OZ4nOZL2p/hAGf4aH+i6jh2iBRphoW4N8
lqff0ZWfY70H+uqR3WrfaSH4pCg7g5xhOG/xdpWrilUX24co9aWjdkvLQQcucHVw
nw74yvRvcu0+Jk0rJyGgJ0ABUxJIiBfkI5+EH/LpCSvdES52RqpbMKWO/Yv58lQk
7ggK+1y2oZJJ6vYhCbIgjasodN65CGQlrSzKA/Zidxvgnv+rpsCksuZSbDOKmo+n
06aAIbx9xrvCrt45ry2OimQWPXWCfMCqkRn/H7aX/y68RJUApIxybU8MezGrf0xi
1bE3oXRJOm+xI1dOdNVIr1Lyj4woiR4rOK/oC+Bb5o7BsZQkegZ8sfvvSRZz+PoZ
k76QLXQyInWCAGIl8lBedffc5I6u2ptUEGQWwR3ODVVqdZUTtvEFC8oJyr25n/Mc
0Y88aTdZw3eoQbF832KcXbnsrM0F/npH0KYaMjlq31cCx8XdoFXDYX/it9LVVFQd
sO2BOF4Q26/UtpH62KCK0oXHWc0Ng53s0eFc7VLN2dIaEuXdJzM9A9p+0ns5akQQ
obBeT0yxFlG5C8i+GdJCA2WNn9Lk3rMY5NS7RcwRUgBYH0TJYFovAPNKwoQ2bgvt
WkiAofnGz6XcQglDx30CUunwzehphd+QXYTaOx72cq1eK15i9ulzryDChsjLJL7X
Y2ySFbBgNhwisjeG2+cyTzrBcHsxnlvTaK77vZO03VA1yFfF0qHPeMZmktOdlY29
+wD+hbWWrd0wp31jqdlBQ8bnWT+cI7GDTMAWr013qKZiYySpfNmtfnWjUSmnpBXl
YVKNRkbY0kSlq8NSvkFZ+dcAULmiwjRyUu/xH7tUPcb4f9LuR22Ml7fv1fOY3dN0
eGVCNT0W+yCM+9MtN8urwHLYDO5bcs+y1pDFYAgRhVggLnAqoUbM7a0CCMFZr6P6
OniPwAtte7wJX4kEZ+6cyGR7gMICilV/rllUdiIbbtKg/3YaBeKw/XCKJi1lZCXT
sf/SLHQygEvZuTv4nNwoQ7UxerECUwSUNiArUPk53O+CE1tFACbNAASbjaAAJSJ+
2gjeMDNuqImo8vj1MxKLmfXGUV+PO86qFVhNClAZqu/WzbbEVeakt5bUlNpvZMXT
3b/Ze3aWJJmDCN3tD/lRf16FwIU26OR/tCKtWAj5CFyyKbzzEuWzYm7jSjuJUp6D
bDzXOpL7vf62lEei6cgJ9OhJvMKq7HjkdMg1tTqK2bcyeSKy6B5VmJ4NA58L+k/6
23ZQXOXO154CiczywrxB18cveirubzwve9M9s93DiUxHExpLv7dQJZjoYhcS1Ge4
ZdcNA5o8DUxxoUDRRAIrruKAzELn4ST1KOI4CYRz/pMX0W+OHVD80KPABoY0GLVI
+ueI/ZoQ+lwZT9eOy5EYmkh8UNS8mRE8FzEi0d9fZo+gdNHZEw+yKLZ5rJbajept
veSOhF8RewKhIrzBYqIeglCFDOsSR8CZKkrq5AeBVvH9FNHTY2/tbhoUafHjmkPn
FzLpR/k9SdRpvajze60Zu0RG5uF5i7qU+4LoGKAiq//n4GwlyTnGcawKg70w3Bbg
qG4bzqOjwvqnB7IP1V46z3OW6J4+WieC32vCiHIsIKOzJiHuujWjP137ong2NmUZ
8m/T4g+GFNQNbfiaryjLLNZtCTzoI28Dtup0XE6fyiIE2Gukj/3TkBeT6/BEhWrj
2BhPYxlM+R0ZyCO3uir21AYKoCS79emEfHfJBlppqZcuEyrCFSbC2Dbb73/jsFQG
YmYof/nbp4o65CoSe0GbtS5p/OM0ADwb0C7NWXn1MOC/ddeAC9pdtJHVxN5ed5cI
qggV9gTONHBFpf1CUH4Pr3ACDhxLcXfeoES18OBlkMIPNIh21EnyOi4n0CQnab7t
rtOIy7n7JFtShpILhsThBFbRZ0gkbXZMiCDe20XnLOTxtmCjjWfnGa5y4qe+VZ1y
LYcyp0tNjAJF9Kwya+wgxosPrfTPMwEql+mFuxTTaqBir97vlItyfbEhr9uqbQ/I
vYChSFOquG96mGi7iozwyFR5C+bU9eNoy5O1863953FptVgZCzGQJ7WLTNT9cJ7y
twh/pkGSbBZs3FZ2WcU8ComnwqsisT6vgY4yjc9VeVhUkIwwRCVP0TP1oxIJ1ZJG
KIY+ZM9zgpyha06YiUPFkSK+ZNIAbQj9NQcp4gsdPtpaKTdkyZ7+nOwik4j/1Jbv
1hVC/R+aiXMDlCyQ4VUFgL+ZqYSqo3VmF0jmqxsRVZdpr2PZqUK3BopYeFpTgber
0zgqsn9Wcg2nnNVlVfBjhkvZJ37eRwteR0SLn0jgU6YVpIb7SXy8z5N4JQyBkVAx
yqqCJ0ZbRlSNw4wMv4krkQpzbsKqIk5XXcTmcHHTh6z3T4ZhiO+2lwgH9au2LRoB
6174aH1Un423y90xOYEtob2b8QYHmj7qIb5SuarLSelfdHUI4/5chR/RUagnhSAo
pRTLRQ/jx3q76+cYP71lkfY3erGwmQW7XODtSiYPe1XaSOm+NvMcnr/OYt54Ka4M
DtpNKFpCOMU1Q6jOGhuEvUK7pJuAY72Gk/Sc36cIbvQHi5jwQp0cBjeV7s2FB2Ns
LfkfoknBmjrZDH9ayFfEtf6U5JgDjudaS8sorefc9OTVUZfHQJsmQ5TXoHDg11oK
xNuvcfwE/HawDS1sibaqDSs7iL3iLYndeKNJaf1frMofr9wcPd3oHd8SMZkzqxTa
NLXU3r5KenJQvbQ9u3BpEKTSJ6JfyHI/FrGNgd5or52o7K/Bj/uxxQsOWXjLbE3v
s3ic7rwUgxBn32EChJjwFOdPHNPtDT+upMza0CT6DF0iypz+7UTYJsKQJZaBaA8r
+BCwDUF66T23Oksx2Nx2KIZcTLuBCo+fxKO67t2goDPgAlO5c2sH1rT//AaGQyCE
jhYRNptKTay/OI7tM5r1zijjqO2c3ZDlpEFi2+LRysDkQDr4Ttn0Q7iALAS44kjs
7c3Yf1tTI1xrxGTJlUhpNyzTZMw3+aYwKn3ffuUusGrWhZ3OWEbtlhGQfYABHZ36
m7+ff4j+l7Vg/IexenmCT1dJLS74SW/sK7fNAbeNRGjtfp2RY7pCikX6j83j8Hqm
tfCiHcEXos4g0Y43gUC+DlRuW3uw5Hygkzg2VPeOxnTubkx/fCix99qXuYjnjGcV
OH+cE9qmp1foetkYgh2RIGnflbrNlA4sSel7/gQuuR9I0KNac3JgWXLJd4S6MGm6
pIMcPtjFZdM3eYols/yaPNfrV7+ze4RBhgKFV+DUDIegt5GR+rIk3oqZEPTW0PFh
ZdKWM69Ji6YgP9BvIF3U8R5o1cKYKfbsOH4ai3mYdrJCexMIJH4Noq4w69sWEKS0
dVUBBrHjzhtYX6kBdtwef3bvi+0c6Bvp8B279zbSIodL0GuncchF49qILfKJgR/2
8Wr+NnjK0FzzqNOpv/qWbJfI6PCBsSYitQiy45afNlLOWc6RaO47UFP6irsooBrU
nzsKvhP1Jba2+cREzu4hgaqby52sRkmFGhpcpSq4mlVAUtCjC8f75fNAT0JpIFp3
JdcrCawLCKGyuIZi+wEfbnXcb6W1TYD4V1Xur1dpNsv0hjcKg+qVvgrSBY3As6OM
FIFtxnhDCcH4ZCiHT5hlU3yr9IA5MeNt0yKKGRApKIHAH5PtQF6ftzoEjjKXt0al
t8Qw29rzFOlxwmJzNHmLxjnoOHhq58VF3MpqJqDVTurAkyLhIoOMlyvxwk4Wbqbb
fvRbFQZwZoYqDFojghmcsvxaV5w/CZjdgBMWwkn7bpD/kk0x5B9VU82ID0ReXOwP
UjoYQo6bL44cG5oUeT93FBJzT50z+5myxnGcgEUZI2cSL3qbjgc+ahgZ8rH6fhjR
hc05Fba0f6cToud9XOCjWcEGDwoW8O5goW4vCpC5E6ZvlxeHf3gyPbubD4JRx2Pa
nZdUc5YDvdqS+65H75lv+sEpA5MhJqM22LYAykw9uv3zc3r4dbErIvlbp1/GZ12y
LMTFkFawrZlTZwvRacnNm+F4TlR2+k4vSYzw29QuujYIt455h2yIu6Kk4GUXwlZ/
VphDaV8C7VUeIEDetI9Ub7FntBgPyl+kAiiTIGWQMQdO6yOas56nHL0pa2gm4Tdm
AodEydiLVCKkTAE5Xxtpzhdbg8MqByHLO3r2AwMozIzoSKmkMk6fintGGDRyYpMH
pPjnnLWhZOJMGBWhygRDk7L8ngCNfHIMxebWLFBMZgTc/aYDU2x2GN2fBiIGuslE
JrEsjRpEVz2m3iTGiP6ywVeNOehwsQ865pz/Lz3FC0u69woibJa3/aJZUGpYXZkE
JsKq6Dvr0CKBVPOBUegg8GtkCbvG4byt3e4qa9EjdWaYcORKEzuiR+0Jm+avtiOM
7R5gmSh9KXdO5Ts82me4KY5m1w+ZTaEPmUXacQ0Y7KiFh6Sr0btWHHwrhclumNiw
qPWXP81ACNSd1wQoyDqfP5c6qUV+8oZJOuevZH2sEV/12e08TClNlGC4sIRgqrPf
TOokQSVxrJOBQFmDFrUbSGegnHWaEH67QD166ZtIaXeFCvkzpMQnR/LGfA+fFcuZ
C5IpMvXSH2XD1ZWICWl6udvS/ODmBL1JGDoRBywmakSnoq9OKSjk+GoyEYanZaDA
hgUR8gpfRsX8jVbrXtle2XiA8INW7zcPwFjivjm8J3/h4QLediC43JwhvGkX/J/S
c57q64vEz3Cvqkd6kOKQ09va3TkdnXT+d15Hq6BxVI6Tr2EK4Yc7k8s7UZvX6qFy
685f5rf/VJTv+KXcE7EN2Rspf4EV/vrReLoIhCe+ISajEnfJhesurDe28KxJzA7u
qXGXtO2ou3Mp/66NfGUMlrbERVqGUpb0r1eD8tUd3TO40XPNoXa31tA1esEMyokM
vn9qncg2JqDAU6ONesFTsIJvJ0zWguumqwuA4xEnMnRxQyBC865pIZ71YB6yX2x8
X0qEdx0kt0QiXXe0jFVJTT2DvhzCblWOi6aqRqJpUQR3ZBP26TRZuj2EHL6m8hke
WuFS5ll8rY0Acvsbx3Tl7QB40aCtPo1dKYtVXLgBBoYV1RFMMvNLYMf9oKjUvQXT
eB/cpDTFjy2n7HjG4U53Urtp7QS+bOaOH9gJR4S+bRgx9S0nvcyx6wbDcZa5c6k3
GW4k6ndEt7HxmAcOHSsn5z86Zxu0lV28WGFOM+2FZRGJ5WM79Nybs8kKXn90XIxx
4Fjq35E3afBN8j7IcPJ71xihUxq+RqxvhCe0yAVGlIxR2NrS+IexVlo4e5mHgjT+
hmvfXuhMonqkihDdKzKj+POrqXj+kB+x0Ba8hd7Jc1x3+qSX60ddLGBGAu8t1AXT
UuSrh9tbkWJ+gOn4hOTN+lGDFluALQICrqYGIcvxjSrB9fRVX3czAzfaDsu0Vf7R
MQRDmeHGbkl+SRsLvtuDLReabGMycmP5ReVc4Z53S0IKnPVRVBkhXBA7Fxw5WuLk
Nf++b9j9s8IwtaAv1QzjgWt1x+Wt1qe4Pt2db86qrdDymcNvbJHMioiy4qOYWDB8
Qm7alLiVb6iTbvRv4W4A7wax7Oq/gonb+yHaCKBBAJXfvCu+ziSosQ69gsZYcIJc
B9XMm1Wm9+Vjww1CXwxK4+vUVLaM01jD/ybuG0kVNTjxICWCDu14l61r0rb4Algu
eKz054ffTWLmbyXUmNZwj6MhV66uIVhiq7tq+JS609RICBYqmRqv2oTrq7KNrbaR
c5ORvbBYbZ7D9RnkkERO+wy9R8Vwakmot4VjRA7uqbIMFYfw5dAw+aElY8M7/ASf
nvvsRBPpqP7ahe8HuhGhRNWrdCVCtx+nn8X86WzPO0BAlDj5MQ6xdklcbRxnOmKE
8lpT9a6GvgdWe6/hfhyTKKTqHWw2sBmccDRMtWzyD/Cy1j9zgyIsZHrcCCsuEFU0
ElfZqJ5KQRgOA5yrqwryKiBCxMdh/b/hySLdKezmukXn+wRGTu7udXlvxmPrO6zo
ziZ2JCD+YNZcd5UlbtY7TYs5L8P2I5QMjaPOq+KaxAzRJ9O3otXf/ebL6wqaZHIs
B+cLBBazJADlJZrKwldneUkOntR7mv8x8SzJUrh07wFjrtaYURQSbk/yTmRaq/oB
MJl2SYHF+jG1AyLV75dgEThX7imRv6CWHJG9hbOgAG8PEpqHYVlUenSQW1ZcVJol
HRV8qTJffCQiMgprqImgRXBeh7PqotUJCP6jTRaYChGnDOolvErG8aydGL6nAWNh
TazJsbI0kC8Zon07kYIIBBrbFFWAqU9Izmpaj5aX2z9B1PdoVnBy9B+VKbwkKKaI
olnPTdO2AQbZyr3/Ka1moQAxt69PlkrRXc6YlfoVuTUXlvRb5xVHd2Nun0xuotaB
1X9rNG+wlUUIl2tOkF1sFI6iSt0WhXyr4wv6fGAAObq+TbI0t4BIOiTD5LRRA5u/
gRmpngAA4HNdMpYyXyQX2oFiiq2XKquKHWYhacVF7GbOVuqw/nGdslqn1P1Yym+t
4ofHq0z6YxuEVfP8wBriHy/UbUnKnKCZQHn9kp8on0VKo+d5+2lRxhnnvq8mx2MS
1gB2Q0WKWTCxHrWgsRXgQrOR6HzcsKW58qYwsXhiP1XwW/VtWkhdrFsRmulW/AB+
Imf3BTiuQplzIh7tbirHBb+YE3FwYXa28kzjB5MTfwhmUmMJ/K4tM8SO8ofVPclS
dyQVn7QlDiF36SBXPqFmJRcnXJ/tdYdG0O7dcnSDhxTuHJ94L5rlPI+/80GIuZWC
KDLISz1y/UavFDmrnzz254TytdfUJXv6kMwjseRBKFa6JaB5IEGX+PBfFeTDWhK0
vX86ewYa9N8IyULFAGOG4Yf1hFC32B+StjUdhKbfdyZHqWYEyxs4R+upRKZCWa4p
84UcVtF37QMn4XGS8sam/n4B4CCyA8a8Ma+FUwaE6MqbLPyyQqHFWm03o/aqghpc
IJlrrBC0ryEYcujC7YH3/DWJFjYSBdJpJ7PJfjHpU2dDIRByXnd4YS0179XNOghy
0ytdpMgzOEFK3ic1ZKBncihqRBXsgQ3mjHlKYhFqntTfe1C6Zt/qNTsUM0EYDZ5T
EAlImzAREdMccZeB8ijztUyXEO3vGB0Ja/9T3Y9kTV7npF38wJKa76IF/BGa1Z2y
/h7zbrEpwfFkEEJzBEXT46agK9eBZeXrRN/HHkC9YVirg7YamJU0TdcQ6Nk6wEj4
EaT73kWpvma7jTkwpqCngKVzUnznWWQarGNpe/Bvp+XXWo+ggqQ9HSlUPTwYGQe8
qmBtZPbnsl1UaY2gI3nqIry3eAWIaRdZ8IlT2Wbt7hf9JEo+duwJ48XwzdUtOqds
4uBE87pTLexCuadkz4kkYfO4cV3OnDJEaxCtNoEkv2UnguAbdqn+ci9GUJgZOu+m
5Yp6VC55DriGBUuYz2ShOz0X3m0KKaRInkOPeJs6kGL86R33JOp808fRhcWyagkL
/2E4y0DLY2fAwII3LVDIU69yEPFyw0l/9I3Zi+pIKMQtFvrS1L+THOe38grv+vuL
dMB+N24tbleTI8oLT7QeijyscPSqP0G/+tSWzfd9mUrGKNQ4FZptNB/PFkw+bb9K
5h0JVo3FEn/sBLBuW5/bmS7Ihg3DXv4T5+nfD7SH2X5hpY6nDdRQ1D38UFY7h7Y7
/DnIMSPBUNRoZoiiXSNN4pgQisFRQALgIpbzI7DcOJHhTIXd1G8GZL+98c9QTQVn
002mHkhudm9k9R95Ka0LeUJotgqppp3N6rQxVaZWM4tAusMo2znmvSAcUdg4oDKu
obNy8DjVcuPCB4MepZPfr5cEEKs6BXRfKTxIvN8y9BREW57l5P+zx5HdNvcB0MOl
FMixp94tgQ9HFPGL6SdyX+YwSD9umzF0uopyCm7Od9+oyBDB0IQ8zTjq8p/rqaDU
g8HJiw2aQSLVcNoubyj/leWBFv2bYo2n5IBy4lgFLxR+cGV48qzS4tVGocTXJJ/i
wUDNXl7LCJlUzCi0BjczEq1+T1xR/TRgmwIBh3U4Npml3+j9rk/ZAniF3fhLvFiT
QqlXy792OJmlUCy71DsBIDMRPoKQULtfnp3v5D3x1SkGrBNrEkAK9L9cg50BLhfA
kdIJbhKaDaU88Usvfg+9UWuXjIffB1G3hc41lqnTKgCx1WvBdjgmo6UZ4CSeeDe2
fxGWxfF1hDuApDu+x+kC9a7yanj0bVZMacYtR8Y2QsDEXZMhr96KtO2Un85hF0au
NbPvA+Jhisf8a6oDKMYBxpWRN7I2UB/sZrMdRY6CvdP9MAk4wkz/dfIwZMqLWK8n
cJhAi9jZy+WWEfnW0I5Tp2PQiptJsXsz2esuzBAajaW5hzjACUmdSsRgFlSvncEU
JjGEkt6HdhOmaXAp+4rHbU2is1X4jguOWnyWh4IwgQIr97x76vbHml02bF2FLUo+
y2KDkVQYGBC4YUFeI+KAc7lwhSl25+RJVrH8ZI+wR17+t52QT6cnr8gdiUVG5XsU
/Cn/gcvXHrw9+6yTdyr6jjZ5GJcW0FY25A6G6z4t6pn6vVMgbEjkjeGxCnoPXZv7
krwHfvkM5AWJ7VniZM1x8N5UokWaws6fgv1CxZ5Y/d2ytGvtmBW57TOYImvm6UP5
oQeSsKZBem82Q1LIt07OeQRMM1Wa86UAoJs6DwruGvzGWVuI5IIk+s7Pfj8JnF9P
8c3RchU+XDumARaoLvaB7LTjSV/hXi9vkFvpV93tcsYm/VNe/Skd7wxN7bOXxqU9
rpOFYE1DaZY618nM5HSvAMMybN3ayMaTi8YTSP7OqLeg4i9Gnk0qjQhKBkLP2rkk
BWRuoZiwNMsl/IqguiXSeZPiginftOCqgTJSvIdi7jntDbxu0HZ4EwNPYA2glWRV
m9DoHnSOHc+7ihqPbbVpowdIGmO+znLsbWtGqhVesDz33R7cAgysDbej4spI/Yzt
F9WdBv71TJDm106K4X5H7QTkuO7UOV+V0VKdoXajQJwdf8UhCPSgUtzUcydsZcEI
/HyFM1ZOUxqGJp/5xWHkXblQLNUzDevQRnpE6n3WksL1hAJ3n2G8yn1VKs+SHKBf
hZGG96KGOzldXHVEUwUFOAtQNZiv8IsTaV7SO19YO2Ji+9hYYJmsp0BlCjqMSb++
0pWc4O4UunAPfR+cjfsznJpPrUBXNZiZ2yDfBbD2zT6ElOUrPX77Tb/XicavCxw5
24Gc1yKKLhdGtKbIWgR3as2Dorvg83Scbi+axaoTIgln/+4t71/EA/w03aXc4/24
L5Mhk/Di8KifRQ0DUZkXWOxNTp0LMPI2HpID6fbNyqK/a//MOc9QgYurDtTQxccD
1Q3SU0fQfSJQs24YEhhQwAxoVrsFpr3+dgT/o58Cw1rApXGxjBagc7XYiWmanJb/
wLrtIdp/+yADBaz63lr+PuJCSbFQRJ7wKlnAVMrqCQR1oefUOXYnk3EEEMTmzArL
EHlsDJcczt6pz0Gusd6g5gopyyWX8L27jZ8LgiGWTyDzwuLfBBQ2waoAK9c4sfMt
95lh18hzEv7wZh01v3UqO6DHKC0CJutmUuYk7GmkVCwLNq+MKlnoNfUb/QZdJEsb
0Zuo4boAG9U86xRUnuhi+Y7OgTUCTGCd7f9Dpc1r5bzRCDaOXqZr154RjqtNdkn3
BK33ZMRgGpviuxJLo6JiUW55f9ybXBZQnYKjQehrKULcKybOLO4khZ3JdEyeYM3c
gY4VwzlSTLJ/9c4PUlq9zaSuB92voi/UjtxPTL7CFL/EVyekBmji3TOjgtw4fXjw
berGSkqS9+SJKbiTpUNN3k1T24Ixp40Cc3oLIXpUBed89H/M47XrKnbeXrh/0E+c
mcRaSirGDZ1t4hoCFrPPtCTfm/MOaeaBPVbY1Zpnfd46uMMlWqtnFmMFs/98RX/t
/s9il1O6qbtTLrk+tZCQLjHDZ0LdXAapsjff0U6271i4z8lQdMxYp2gG3i2yVUpD
B3YfMpiWLXGHxkoOV3m2+JY3wNTiRxQZv4auBv1QnQL3BYdYnQp19mQxbq8lB7Op
eTvWWKudFe+gJGcF2V6pRTscBYJHSmUSN0Cguo2ai188P9nPwywhDaZrc1g0D1U/
m/Kdtbmp7Jnf6vFnC7CXZWBs9+oavwpVjwH0QoyEDBGvm3eUEAU9ZNvoCiokChWN
ktZVtyYkW9FZVmvuGvli9MNS5Sxv8numvWzxsoamkVffwM0FINAMjNQ9AuYM38O9
JnOTKCI8ZZ9J9egyzy7yMGEOyUrMxFJowGFXa9kY8TwjZLkWXcbAh0lhwjjhjxyE
ckv62D7VMewg89Xex2pCBo6s6R8pEtDV6hpiTvy6lDxjBCgBgfEbXi7M05trX6Qp
gUFpI33Q3jdU8LlO4MXc2vKZIBk3f3aTmsPMZG0VNqmTGhn6Yfzd9oCXPW+Wk1Z2
XhKXavkXweJTicrJwOEZvFZQg+5IZfauh8dqcZzzAhFcbaFpIJF0uZurP7QzxP43
bnv7Tu8a+o1mJuTAx5YBHrGkOGk9m750aOTuUWZLiFurPy23r6qO441DH8flhmKn
zgUKmG31Po+cBgvle2yruLUoMZb9OTDCloW0ckYE9SkR2Rl56zAdcbIIq4eZQnTs
cqKasc6SSDWXPSfYZnqlvlB3vljhSQMMWTDvx9XH5gv5fqqGZZOSCrOMeRft+bgS
o5tpmB8Oq+gObzmwtF+F0BnTBtBtJk+mXvqAcfdyJOhyKy/r1awMNqLwSALDNimh
Q1q8c0clnlwW4Pl7xSCyJ6SgwcyDOuG5RcpwIT+tANjAy/uxA39MWvcPzxMZwzyc
8eMoguYHg2U1u1yMjRqRMfFto8RKXOkMBTFaFHhErxwYdZdmZgj3WMSrXZnM6RVr
+6zV8oPsCw9gXIclf+sbERT1j2nIQRxF2Dznvd4fEYTtY7zQrTrx/UTpiY+XbXKv
iJQ7Y+ocoALJx/AXJL2KOeRChTbUEZUdcfghYnHISZ3f95Lijiw9XxoTpJa/cLIi
rTPDU9nNplkWJLc46r/5WSAotiAVH5d6Lt926cuitBB1ceCmzTMuRMWVnhvl0ems
QNf5hmbPfWbJzmVXoJAtCt3iMp8wprBYEKn8ZIypDmnXJnM9wVZeLlvKaPmKs2Zz
Q4ocUQMmJ6XbYab7tbvRHcTu1C6L/dRhGGJW3gHoDI9vhgcno8mWvvxCaDD/e6Kw
IS+7Fy9rexCVLMezWNoKHuDNs+y9Zk31sPywDXjroU/nxzeHpJm8fP3GPnDl3E0P
cUnuVxibf5CffM1AtPtDoastcoqWaRkCELnuYpqIX2vJYHu23dAIQIaWr4Awp0je
m/lp9KBSRqji7ocuf5qVQlGwkMiERg0HPy0+W+vJwZQ7iZP+C773nrXDYDMVMp2e
S+mHBOA1PYg+l6ZDdaMhrJlg2Tclg2V2NEGcUt84NoXIiWqjXsAgRpHxaLe6zRmU
2kjI6w9GoE7LxzXR5PCm+AYZqqeOz9MfYJoEjRDsXEwIhKN81sFv31y0IMMy2JgG
kds1jqzDHMQ7VYnH201yVmhq6gDI4k1Hj75T+dg5wfrrchPX/J9VeZxX1FJdyfBI
QCWkE0o0+S0Fsa+NRqG8+V/ZaCy764KNIX21E1CE2jGQc2MtLPsYP1MIrc0q4ZJl
W9T+us6SDStktWqCzYPEMKBjjFmDn6BBy5xDJ8x3jurjMpt1a7PG6vqJ3/NBZQ/e
59U0AjrUHHOFlyO7tWs3eWURT8ZYwpgQPrq9y/wv/bpT3/8mvGIxPyjTRQESyiPa
pA6oDevfYBE8IhGqdNlBBAfeREq2FfH2j0KCAR7D14i/rIPa7R1AVIo/zjWJiVQr
T9nE7pIUsIIlfV6HJaqMQU3rewiTl4yAN7FRPsVrOKdcQntFUNrwm3QDoS4yAKIU
543ztc3u/gdhnL51IwYi2N2srK0rLzPPgLpz9ta/J+H6dbrHyfjzaL5so068+vwx
ZkYpRWvpuANfrFrg8yxSrNkvJZ8YVYevAc7Y9MIe/DT+arKoOYUhcdKSdxOL3MT/
iVG8rNZ1J4lQjZ5fIrIEGGxDa5Rh4O2J4SXxDj70RCbUIPSN8ppNXvEOWNExaV2p
IciMn/P8INn5TMSt/Lt9JVtx/xNTFY8UrPkmMWSnQ2kR0mRwgws8/TMUcQO8eOaW
+v+dEmT+IWC/2+ZxJPFX2gLvGnSw7a+Z42cY7JxnhwIef4rcx0qXINWVTB1+vUzI
sDkoRkhmwEfjwAD131PxVoabM/xsduU0DnY5ndfy79HOFIPPLn53Rf1kMdk41h4U
Lp3ugKdNalgg5eGH7mLR5NLrDUR0hH66eX3XsurgOLc8DM8W0f8+K4cZp+U25CLD
p0gIlnRqfVBimGamWuRZsGXxlRS3C+Y0CnGRmjwqlGCfbhWpN0/meenWbw0hLPWO
1ND/sEIxAsRCdhkZMO1UwJaWLMRMET3MHiUEKN1wRxv/m0en7B6l9s3wWUpboAK4
Yy5tbWpcp8wQrGf+4yrc+cN6IfMjgJ7hV2ZkTzXgdEmlZb6atECLetxph7ddIqJg
VkplPfxhSd1Nc2lQu1UPKAKsQMqnaQAruAgXFmhaTMk1IGAea2XqH3XAIf7wfn5j
0YrKqZDmPGHyo7Bite0O9zLrbEJxAv44R+E5R0R4E374AKz8vKs2HfzaFO/4qtUn
lRQHk/W//+gzf/8qTFIH8MRlR4ht2jd46qK/Sl0rBnGi9osucbr0JOpaKINtNczi
fid84miobdpEDaSSs5p/7ZteT4dynxZBqFxVHX3SU1vKTsEzXlDSqQ/PAQqmLHOv
e0EjTLp+Lj36l/AXAbVpYe+M0KG6/rWmNKGtLIIDcYaR8HuWNr+ETjMFYnEbaEj9
OXvq0q6Vj/3TXT+6f9ViiSAXZTrGPaqPeSwgGfLshfiEkg9DXxfAJSrrIWKpUvAo
3V0752Y8HyAABNE6zBxuhrhbatjaRD3upeBrzn/DjD+6bxIl+TArZM5UxPrtYjzO
f1cBXTimzrm/avaO0grOpocKKWpKQr/9z26fHrKe8qoU/zz45kxbWP1pu7E/HNwm
36nWhgDf3oumTiwU/D7TAObmHyiXCrYUaEHphlD6xF5ICoFb0exV5b+qNu6h0+4c
oHNUGmJjVtmd9M5cqW96Frt/wNBXhWlEwEfSeZJV6REX41HvAGbBzQvm3uGKM+Tl
iRcFcYqHmGP1Sb5ls+JdwwTqua6srBSC5eappSDnAlwc7ibflYomrG0H49ncrx1n
r56NFoR4IjQQzZCDHjsIF8fbuaDl9buqHKNhVttB6qVvTT1HjERXWKmsLUJC305G
CG5aToe9PjfHxB5qWNJy5kqqPii4ZlMQ3gF3lJtkR6gun6/QEzDrAUZCcCyGSwOW
hpJFyKH/gW6zpkWJ9+biZUa5qi8iEt3ReFnkchvixmoq5Lx3p9OTzYL5PMJL/1+L
9IkZH4aHsb7qCEIa3kDUr8gy46sg1+wVp4KGTvmNPNBTnYJY9S7YMCYcKlt/SQ5H
706qBX9UYRavvADuiUWiJrBK8VeVpwseLjIWQ4PhQZnyNDoRHz7dngiA1manba1H
7WdfRKWTBy4f+nPPCRWdag6d989K6GuQYnZjxPEyZJae3FTW0T5gxTWP3Mdclx19
m6AZdafvkbVuJhMGAlDkPBllLEVoVSSDtrhKsa+gZhN1DQU/KUD14L+6K8XKzKEa
6foQt3Rl/7r7/Hgc9/0ey8V7qQ7szUW0kH7qsIpwHbWPUg9Kx34olmQemTKCEulg
1ju1riqbwPyuAKNtW+hLB9ODnF2GiUPxQ+5/x8HI+1hLH3s1bkFmOg4rJReNw1nk
TjgLH5SKfPzzY46HI1Xb2FXlYLWYd1cLP28CWPTkcOnL3XE+AJu50HC/SL/TgSYC
cKXcY3sL0Hp11yIsEv1lUvIoyAg0epnvgnbvrjqQQ3L7lEblMAUlzkZvP8uDelzR
Xz+iArUr8VY8kCM12rBDPFBnTk6ktvy+SSNZjVmdGtGeAjfznBIaIVEnHTRltky9
TooYY2YqnPOFuzFieICZXL4ykc/M7iI+UwBO3JRTRmLVLXngH/lZwRtpVfri1cAE
SSDhlXPD4GK9nHLmMdKIZD6cU1kuHSxjUpy03+jmmPHzIAKyAhEftc+/QiSScxhw
1l4mlvqmvNBgz/bsjy4Qv7h40BBgkiN9+SJaFs3ZPtSi97hwk7qRVUo2voP4BFgm
bQW3dPczqTmzbW1HCxCKk9mj7ne6faaGt8e/sO6AttFV5040xIh+DnM4Grd1yzyG
T/2GtD3hZuA+Depgh+RiLxSZ7Hp7qJaRazzCauf3fHNfMx09NuE+8aFtVICkISvy
QePMtgZq6Op8xQmCNmYXttvZjCrPMIjFGvkvH0syPvEK+tZx5Ug6HjqW2CYyY8rb
aoyuXkj3p4vyIPhIgl5TQL7KQrhw5eq6b3Ze2ULpvEg2fM+RarKQsk7K+sDii1jQ
g4UscddconCDSDBYQeNk9edDhTWf34T6op4V0ddtysESpi3JhyJx2siL/zVwcuJh
imkQ7N2TrS8m4xWFukEYmrbZAheNEP4ukBOBtDKNOp3G1Nij3wzC8zIoGPm1rfxl
p/eNtOyShvqqmuuvUFBlHBwuNdzIIQh5xOWb1FeTnFrmNFMrfIbbyNY/7jrxhhN9
wZ/htORjT6jntZqilD5K6dqP6ORGFqOh0tVbfIkkq0iElKgeRRpNAcjSujf6sOPg
XndQe+eO58EJ3SoqFubvM3Rsp6/DnztA/PfI3IuUfKyy2Z0zhdlnZ0dv7X3jvBQg
nMGi1kOCuRDsb13EyFFFZ0A59N5cbQF7AcczRsgVrkMCzm1aX0Th2sTTPEg1JvBy
+fKtnKz16vr/CyWtJOwLBeArai80zWIPodKUOAT/miTaj+PDzGTucI0icrAuVi/N
gBqbsufDPQEhyrx4dApgv5BvduZNbRH80WpT7uXZpEqG03gakAClVut76UavIKIw
QR4jzpydWoHmdJTZpYavxeMcVQpMS06z7kqJaqWWpne4NmtKp4U30wvhE/Un866P
1d+ow4a0mRiwsUviW8FyM++DFa1q3JxQmwVUy+jKS2JUwUL0WGX6jkORQ+FSupRn
9crSH7hXYQfHy+NeS4dFhtUEc4BgSPviu0Uown9u8DIWHn9tRHAkIqTBLUJatLbK
aB6YX41ssmSZWw0xec3ceeDEzzC933IlUyap9/Y26/1t1BpbiZjdlKN/5fpPYh/s
bMKXccadBmmFjDJZx0/scyfaSMnaCcDNAn3Dr2n5rD07Hnbb2Yo/CdvQy4bx/XpX
lBPhGSyEurHUxRLXdVda2EFceyhpXh2N3GiJLSJ07xcmziyMIU3JTwVETQjamn1T
hkJD0nvOsaGFXjkLjDx0jzBo96gVHDw0Vf1ZSxgp9RbHqI57BZHcD++y0/g7wLKt
XL5ZFWZ9ycxLlsxvwTNzaQnNJlj+Ar3ALyfjWghweF2BuNjHah4q1+BsyxkC3t6A
zwVtA8pIxdjRVVIPVrNTnb7MkxIkIMV7IQKflk3hf24S67BGUIpKXNL8h4ZeSzt8
5d5uWIrfhbMnfqbyd6Q5PNeRbGg8ENTBl703VW98PMC7ph/2Z/YeG1FWBEhl+wBd
T8dwN95pduHOJ4gedOaqpZ033RBtN5/kAeWfx0sm3GmPxxscIqApUdScfBhXXXlZ
+X6HJUyl8R/xn1YQmKOYG9K2lYGtbCYAxZnxs7FTrnnANKs5NjK0gktR7IHvAej5
hzwcmFvX4Hfict5Tc2Jvm7POcWTdKs/sJ0/7bWWD67WeZouEqPPCpl7PSOZ+UVM1
B18hYR4oaCt3dwU8nqtjEG5D1pUWk4OQbMVBQf3PQW1iJKQSKP0wcrdA/HtOc0yV
GjGgSV3HUkgb+QraMoHUrItk1kaao3ozub93JqSh7dAIHUOQBeNB82erNds24+pO
id5gQOQOB0yV2Qqz90vCg0aHaqp52aEQb+d1SuhMuVi/3zKJR9BHL7COXA0w/Z+Q
WQwNQEWT0DVdV//YsNFZfA146eqMXDSpN07K89l/+ks5KglIi6KSjHB1Ke9HAAP6
ytKYEzRtdCRWjib/O9Oe+NttCl7ZFG2Tp2toXKY9y9E2T8B9fxJyFN99wfGQ/CCy
Oq5a2ssYHExNkAsU/GqoHFx0QFJmV6fTFOs2Rj7ksOLOWjjA+kfrNeAXyO07u6T3
LIoFFS2e3Us9938AH3tODDF7K4EfH8oJjJQpBdWKEcO7jz2o1hyoyOI54KZ+Rpfe
Do1/4JqyJ0Fge96I3LVgHjBXyPnAfSseHkXDZ9sha7Mk8ogcldChewJKvmCjFE0n
LfV+ECY634o76VmXk9/V1T8XuKh0g4cqCzCU8/7cD0drEOK0RcfW39MAe1iNagkU
H+lWs3dtBLneazefTeG8TZ1tKobiNXgZdGf5e+4/rREm78zxrMhKWV7Qv/2FChEq
BuUMCGkOo5GLY3XMDEW/X5ve5yluTS4dBgRuWlEBMTtLXBZ4De7gr6jSfLWWcTc9
ZiNE8IdjHPB2JzEaWKPhMay4fgb8xMPBptJlZny1n+l/e1fQhlu/OjpVSrAWEzH3
4TQ0b/xyiMLHlQd+HenLn18pt1xFYonZnGJpGjUdCw9AWI/G/LprUl0tZG/mTh3N
5vVhy7pVLNjRkSaCiE9WjfzbvLSqfZmltMbbbJcZEDMUkq6RZXQHj3ZRlBRgoDMc
UcrC10IIKhTMIsXA63zsNxXPZ0HKM4rpVb2fhEHHFVkYMzS8GZesuaItk5FI3m4I
8WIY8q7MxYYYIfzf558QCZTWxiAQscbOncqXpOjBwfNfff1oUB95L20sKt1UK4Cl
wSKjrDqxSvsmfgKNIiUhZH/A2sXn+XN9U/HAooJS78GrtzajhX9u7+he0KIsuDDs
hcTYbklEiYOzRRsY/bDMHuBmi6rCKYB4F8MWGDMtH+n6qObR1DY9KSpvtXfelF5K
c6Msc3aBPTeyluaJoMh1jr97eEsEfMfm84Zr50z4OFFajSDQl+YAWqynNWQS4S+d
y5IjyS5m257qZhCB1Q/RddykQCbqogQuYIxm4WoAFkWTdWhEHBWWtCZLrN803S9F
zCFKYbShoIolqHu9e7KBkt6zzq0AjioQaT2vgxdslgRG+FTftOuWvG36p2sy/sud
0mz8kaLiX4qx1s5guhU+ZI8fpnNKc6ZlHiDFPlB2B2qNmHWMPjQmBxW/rmWP8PoC
mIBAEC1uYVCFKQ2PT5+FjKo7NWaXoOC7wlfGVAAdrJx+QHz0zibKbAQ5qdwZ0FA0
q90LuUDlgu8IAwDF26MqkqbONoHcwR6q7NAivsljQbUcuNfXmJbd2P6Ex9N+Oefm
M+Kn6OK5IiQ6xKQo4RX5dOobd6nTOZywD7q7IbTAQWWtv3R/GqC7cIJq5srNQdES
VtXR/6NW3sMYwOWZbdYaYx6ZbSyPzJ/3YGf3JtqW5UKLyrb9wQWeq8rcl1mbN7Rz
3wO4z4WGQEZNNUFbFsBUUovSnhRiKlU0qXp98g32NTYjxeHSZWuSTV/iA6e3uk6H
dUnNsT6tZCJVQ+3uYG83JABUfXzSf0clfVG3+NCTZNUXn7SGfl5I+uLR27djIrYN
drsHiZ40nmgymjOh3FGdg1bijGiIq6VSU7mxFRjQnUmZ01v9vAcuSE9VTCV7wCXk
r0R79Icht7InLeX+URlKaNshNcEOoccT7D8AsAtF6h5TPqsSUlPlg8H6oESdj7z5
KzsevPWeQOqyEyUAg7pbKrjZc47d72vP2FaONsFkArAoe8SLvIDZOuT2BlIhlcnu
8WcagiccQgvOviAHhCWnB3/7+lOtvQpH217sQ/0eNmz6v0WcbLG+RCayMlMavJN4
pyV5RjPexA3NybNtcQqcRv+WKDq3NW1Aw5FQt64QrF65ovRMFdoxr2//emOA4yrH
3gbu/jkeNI2h9VX021yZA5am5xODLcy9kQ6tYvIk4lg0UF1KgUD32yIA1Nc48pot
WYvXuXj0t0D+RJw6hpEjRGTYgs8j0WVkwOtLvj3fjDDJC/eFEBRTsWz8LXp3Mv8t
ReDfj792COhqRzduyllNBXp7FhzJn208xlA6PuF59J4xdsivO6R3E390Uyz5hiAS
xSpkQ51bgSC+7vOc2m8im5H/5XjFO8DGAVpRUCCxnj6GSp3fQotMQG2xt2XqHVbI
bphxJuMPydbmRTxsQdXlNj6AR8CjpSXaYO1RVbaw0wnhJ1lrvR9IM1U+T2d9+TB/
KJI3EUR29lM587Lg5jYRl4SC53faY4kw6xoagJbHnIL03a0udunquFooz6fzo7cw
dVPFvysCRDhdyVSnLJqIzYmDzISlvmRscHtIQEDL8mM8yNZC8TNKjt45/EUvmRgQ
NOrhu36NDWGRiTHqy1TbhV3PU3eJmkCStDr8BFyLh3vAigMnz5ybCWhXXpQ+Kdrg
GQVCclDYuwhON+lxTXdMKyec1iIHiRfnZTRg5ENbCD3/UI7xzMMjj17y4W9/ZhJx
jy90BJRhaRJ0C7Cx35VgsG/iWx/nMqnOXIYWIWV2vXv/TME/8qEZtqt5e4fdE5B/
E/vn12BUUMPyDUUjw5ANTHG6vWI3miIae6lyYPmuNYmqmebQW1BhX2MPGjr1HxHR
YAlVy6K/N1jU2RF4f0Dvow8k9js6ZW/EE6PQb/qrT9f1/yuCETRCysKJVjbkADa+
f6WRPh0ZyJY+2u/pSExmsvwNQyRifjEm0RlGltQoz48A6/k209gBQnYpDxAcfyed
lRMTPCLRUmuvcynUiJ/is2p0+4RdmkDva8dmXdnZYHHFYIVwNHNz/3rVLnocYnAO
Bb/8/wMv/RDusjc24Rk6g1CyE3woVVEFyH21gYuPmj/9sSi9rWwTR3SCPdPZPShS
yyxZPoo9cRXnEijAwISzOGAN1zSvBtodNEUhASyF90AwPfWLbmrcskNSHKiwEGnq
RwicPeoTpUuZrSENnB71m7Ojiy4BI+tByMX37RMXMFIT0fCY1+4qt7p6kdaxr9us
hK9n7+Mfab59EcLqxCApoZE3wDSSygCQSLng11wWsN8bQ4Gf6L8DtSiXEqxG+Ylf
rhedewNScKzr40s35WnsX9EXEOQk9hWQ4CFadBgBcO5GwFadl6hNKvDID8zSCnLl
sNKr8u/TfoHZiJl38sHaH8CGNCWLlbpOzeWVZ7z9gTs+o2sbYBCY5ArP6s6pMmUh
C7sGfh6ja2wgu83mkxiYGU0PponP9rENAU+GLNWciupTMy3Qf/xnoTyDFzmq8vkI
8KvNXHQQtyu5XdBmwlNLUsqNO8w9rRRpOyDXjylpH6FWyafM363IOmOlqS3+Jgqy
Y59K7pCMCcbsHn42Tw5c9bN9qe+QCNCSyf8ifJ0GnXJb5aIYHvhN/tis6Mkbig+I
7LKuU1djyrRNc7dBLnalH94cVxu9nV9hvgCYUo4mJ4nPqssyb/xm+O1RMD68mMUU
8vekQ+YBl18g1PvTNNlSxeNVDzx6gzQQJYMGolCYfvlizShTCka/N3oAcvhfv+Ku
Tc5gf6lQr62jVgZbHTUqtbr1yVm4axoNdWBCuyEZve/Ck/Qoyew0nP3IFnsLEp5p
dZ61WU1UQBsMfFOptAF1Ln0pTz9mU56RrIh8qGp0ZGFM3+z5cyFJ6bMeJq2LqH3X
GeyVsRTp0FOlaSTLDIFr9FzVC4DwZTeYYkvTyp+7HdXUudZYO4TInHWvsn2vQFZk
IlTtiTTxTJJmjE092dHV2yDLKcUGk3pAb04IVtEvDOKRogWEW+hLvkL5rHdW0cLr
oX/3LwGZNA2vUUndrcvYwrHCYt0lFvX03nPL8Th8iayyEyKL+nww1MFa3N3lY+5T
d6HYso+ASOCvoSQC2ZRZXXkzrQiCPi7UzYW8ItuxA915t+glbQyg+qVHE0FB0OX+
faTEPOfD0GeTIYHUNrhCL1knAiJXus8E3/XNWs2Y/LMfKkgWZvSNlELiJXxnNigP
Nxxir+9F7X8WvnZSHBI3pcLfzxE/MoPX6ZoPqh2FwlHqDS0SlH/eERqVZ+tlVSng
bQLiuuw00rRS5RtLKXvoXxbFLeYTi5V/ajaheI2qLUn/la0yrpPmRjtnIID8m1Rg
mjuDBqpC+erW8vtLIfK6ADr2uZH4F+NaW2LBpjfZ4Qsr9HDWk3/kQ7MeErJcLnOB
wGnF8zOBqZkkAn+CldgeZkfcPBZsHscSQ3+oBNH0i3KHAf+Y3NF+noSy81xPN2Ty
tE6+H/biabcoR5VPJAkUEoU4DKnqdpLMrKNK8vL6shv2Y90WPDROVWRo8Tt5Ssct
2Pj6mCR9r2+9ins1Os8NeWP9xaDgC3+69O4GU3aVMbJWDb+V13Z2JuQLfi5BE2QD
Cbe/2CzhaMJ0Ph/NTuBFid2p0EyPeTbatagR2/mGmXvnNzg48kq56kNR3j/76IVe
fdt7J5CEfSn5aRKo3KS3aXbKPOD+LMW9U1QJLZgYNcmZnwEo1lxIL7rK61Kn44RJ
FG1VxyXBw7bMoEJLMx7Se1KHuEklg7SlmCjlUrZX4E5NkhHTvvmz+z8MBmHW7QJg
nJmxmhoHVnJni5R1QNV6EuvkiKsOErKaL02wFPt2cu/2gbjJtGJEzNn+2YWmmLKp
b0R8HzVVjpDAilDqKLutIIp/7JWBu7PwhZNPeF+F0cttLQ4WGkCEa0sSx/sxDdbO
ybGhDGpWZgQL5UfMCS63zoFwGzuGwYdspMJDhEX50ePsbq73HYsUulIzQHDwaFmQ
ry3X4lin7bACZIXFHKOAIY0QYwteAC4g0jKtMA3zkR+KGN/tgzxdnZG0ozmkCQAl
NanV0q3MA8UylE+g8EjIgRP/HtF2DrCS0nuuKX1GQppFuK3JgqpxvWsCoSJG9P8U
0kGKpdWzYTz0TKh2GfPG1c61LaKRrrDXUSN/P4fZfUBqrAHajGyKBcWOKH6CYler
GdjRLfTSX11TU7BXSF9kSKIqjdA5RZwX9HVY9uzPyGGV1pp65i0QbP7dfkMFUUDQ
wpSddEcoKrbI7F0ZQMZK2GsQ657Kt4YUkemtJdTSOUfmxM/StWqDDQFgjzVgQzTr
wry2BRDtJESiC8/Ofe2GiSja/zkUVIhRcjExCe4E61GGpDaMV5KKGZ9t9C3atA7D
xUKut121ZESKBjJovtwlYlVBUdxactbOP2ritKxeVH3QGow+Oa14T/34SrniTc34
/KSkhPW0ZuwkQPfmUt89Vkm7+XPLeRaujDYli0Km3zQoAsmesvvQyAOayOcgAcrX
UklKV8vywlEb12govHfOENyfzQP5csxCwzGSDAJ155a3CfXT4Xy0WDZsy6It4KlZ
40jSYgkuEqU3XTr1PRlADW0SH8rcSNkS6tYPMIsgaWcL0ZztV/VT/51AR15ol+Do
6+HigE1RKlNZDAqC7vVNZnvmV18838ftCg/cOPveiwn79xG/i/lhMQiZV0D1aMKl
1thV1L52bmgcBmiuOWF37LwxUHx8FobMLbHSxGrjgbW2ZNVXZGaoxnseCWF178CQ
SLHBMowIKbpSr6xDUcEAlxKDtqZPGOluSBcO5XwpV5zLYccDqy5WdUdWbm/GvkNk
Z87yx1kDbyTotJ1Gx+0Bm4NIAdRvM+31JBKJBOq2ZJHrGXGTlxn1iJ4nE4/s68PZ
v8zmBX7uxfLrDX5tzJGfmvqFHs4+ywJs4Opc2Kth6odDPNRYHmLyTMTUyWXZKI2y
/DtPWbtoSr7J6s1Xx/kGAjJv3AwjxATjr1RqLjq4Gj9PqOncnnO1vCiDznhDCS+G
BS9CLY03SdSDH6sB2mUM3iofb3HegF9Tsy5HqvmkBjiOQqWDJ3WLEHen6M80WbPT
bvohs4WE+e1Hu/k+v5eVZQNZSG9C5g3uCmgYNeTy0YT8CPuczqQWOW4bQCRXFrNF
koKpWO6QsQD1tUyqoKGzGe/EczsRsL93ICnebshJZmPdcYusts7ONRVjdU1yHN9R
IqLnGiU5y7xC9a8Y9j7wiCbh9cBCLoaFNWbhjWzT2xJloVkALf1iC3akloDuUOBK
OlOspugkxVukPEV8KnfcP/0VZsp8+teZIz3W0J/Tb0Y0UBQNGbvIv5Y0mQhg8qhh
4ED+PDFs1cApE63+zboar0TwMmlyN8L0Lk0g2qdIuJ4Bvh94ajWiZlQ9UhkUKt7V
DnXz2pyAsKKyzD4KLNrtDSo352+TP/zy6Ilsj5weZ2B7LE3wICN+tVws5oBoOtlT
D5riLLwjbnyO8wmEvRicCMiChjLlntRqoYQhpywgL7JUGf4qX1S9W8X/aPIAgc0H
efDOQApHeuii97xOzrFG+9rk1FjsNod1as4Ys1CfDjktE543hN0zdlp6az6fhSU1
nP6hgVwO6HIzni5g8pBnk6PVmo8556J7TWAKxh0EZd+DtmuBknfC3yp9reQNmgNc
JeyNQRDshdgHXqbNJWZg6oNjGZUvH1KNCwHhM12QpdP+ucram4B5wupH2p+WldVw
iRwII9ZC3DwLRyrSghtTFswYIdUnhbj43Fkgeee6xIwEZNN+2VNjQWLmX7GzaaLj
zgpCOQjfyBazkwAZeKq/9bq02XiHpn0VTou7iEVpzxuziW00cieT5k7ZVlDKTKWu
8I40M0mDqBSG5gjdkt3y1hngLK9/Pgi2RdE3gjT0AAZYpgeY9azrUKT0bBcMqoRY
yZUpvLCrvMf3P7qJhWnaeUQACrWY40kwl5JKY0SvOBVdi74V6CoN2Wz0z0kK+e8j
kC8NK3paoaL39Kf0RWapL63gfieEX+3FwPrWherqoys4sRb+NX8cR9v03O5LWMcG
PhQpQ8lXlUdtqPqzTrrSyp5UX7fasD7h1mu7Cy+cd195JC4yARTdz0Z0szlg0YW+
pWEScI7ouHFKEkVtAPZSAe9gDd2LrLEbuX1h5wTWYooqUjiXOIE4rLt7ypS8g0kv
0BHpAlCrZWeRazlSbk1VrEnmWGIDo24Wtbg5hmzqO6NoqP8CpDR0oQwi1ISZSnaM
fdQhr1sGOtR8ipS/jnnYP0V+hl+T4y8gYae7A3X3jDl3+DxOEQ7iO70fKpXidOaC
S5wGWP1h0yf6SB/DDSOlHM0YF+B61BzJcUUbVoCq6QHahqgYhffF/jiV8c6MvP9F
5ED8m7kXSuUqJFZlmaR1awNPDjwbigHmqO3kuOgr/eIGeRgV0BpHVLMdgwIgqwmS
UXBgH0D5FmUV3I8dyccJOx53XPKdM2m6ZlRm8y2bVvI5f0d5FgihyuwnctdW2Pc4
mbBcfZOAGOUnuO+lNeDmlYLHswr0aExHo9IwTePg2rfl3udHCqKHCgeRfR4dg3tN
CdydYBVazZ7Bi5qnzh384H/6zeQv1rPwJ+dPnvmU/hFrdW2i1Wr4cxCISv6gc6E8
ZIY/hkC1IHA/h23CjkWESqgR2j4VSzVXn7qDrL78n7dv9fUFgUDF325lKaiJScD0
z2tN+G8DKQASG86vlfGhA80bOqVajH6euezvdjfrHj/HV24cSa1EVeRtjZxd8oJA
tjzZOXyDQp8vFX0UaEXu1W8xt86Zu/wzFSjZLMQcemm6xXqEPMLGv2oa63VSpOzq
JDximDLKWjj+i5ryLQ4AdJaSZrgwSSBlgs00IJtPOrbgwedFf+xnXq+iceprheyx
HabWxnYdbAkq7oHM7w+eUjkGBeChxDwNcpiy+3ffU2qBe281PKlNcmQQyW4OyJpH
hXbucZdxigeaNbe/0XMPgRIjZWhqYyrY3RObXHBN00Ia2ZYwq0ybcmL1Rr+P/TN+
AkVZ2UGUyVjffyEHPIgeWTLyvVzNsla3aUYIhu3abGwWNT/iMmd3DF0uGlzIqvDQ
tP1fipaz/b7cQrdxVlEWUNZoNUw8YFYjdrYr2H+tDe7LReDX0Xmw7o+/uaktvLLn
PBNfkEReIsC+VFzWp4HSn2Bi+sHdUng0kvRqQhdAr9CFobVDn2ZYvoErOhkIm6EM
O/sxuEZg7e+HCtK62k55kgBJ5HiddnPha3w067ahyIyAtiKhzDiiyWU6qw+9Ko4u
PsX74dZFeoP09RUfJzx1w+6CUUNKTxK3OAv7393d7cxh4BM+vSzxSTVdeN8uYUHc
cqVP5vPFZM5xRSbVPF7iJXXRw+QUCBNTieyr3Lddw8L932hOf3IMrRgJAZyFTYNw
0u623/sOVPZDvTy2R5/o2wGLHkQkjnEuVokQ7M1j+n44wlFvu8nwXonZfzWeIKcR
hkD9sY144ZkJ0CmS8L8HDlZq90BYlZe/3U7pE4djf6z0Mke7qheOlznHiC2bFxR5
oNvAcfeY9HPjQwxHbZyh1UFuHdVmWNcz47HoGCrl0BzNoMt3nS+RgYbEXAvdA6aO
aMKTquoGDuEvlyEBrBeN3iUjciIdvkzIoiHag1iY56WelBIQa/hIGjqMMf1pjhDg
3FeY1RJTphxWQDpi0Nx0+2vS1M/D/JFo5bP79GbRpSkYGQJShPjokSUXVSBg12A8
HhReIcgSF5PV1Z3HXZGVoiZTZ5C4Y2hgI2l/yonfmXXnEePopD6uEwsEYwWFPW6R
VMQxVIWjJf8gqRO4Y3e9o3gSPaXLkMH39CYQeoIKLeR2jTOtfm4XiK5fYMo4i/IB
sdthi1CtB6miMyaA2kwkP5aXyY2BEflDvZZ9Y1hH28Re7ckTPRdBGVDIQTwiGsJC
v5KYch4ZFCHq8xjQ/vs8zKcTDtocfHdVscGa3QafcelEXnwsG5Yf5ELEHDh0jvBx
YAFCsp1N3CA1xih2tyZ2FK0G6rSYPT3+EXrlY8K6C4XiB/xb7YI+5p/2GoCzD3zQ
+3sJI5jT+majGjY1eyfvXe1GuOZUUcCZF9AahAuN12IUZi7jH8J+3657CHyaW3Qc
ZW2QzBH2FEr9kBhFTHV+2k4ZGT70EZfo3quOfBliprVkFWtyU/6L9fx9RIn8Ieo9
V4DVsHThS14UXzy0E5Ct9fVN4IRh4VA1Roe51EDgg1XRj89gJbIVAIWEXcAuWZBP
G0Q/xfHOXiPXEVfRg/kSSPEkepjovt65HLk5gylwZsWZJ6ubx1bhMRTrBcnWmUH0
em8p3SW8c/Kiv0BdMc6DdnWhc6OEHDTqT//3iOZ0Hpw6Igw/ViaYc1VDV+99DWQe
8UzavMvCYhR16GcnXVkG89sumvt101tBKE7VZMD+semSGSq0+bniZkqJE1kamZzu
wNyqlndpj40SvMxocSOqOt33g/O+5ad9gD32JFskXzYgczZDEYqIxEDWlgQagc7D
MOMNahi41Rm93YHY3KR1MFzv1GWYLupr+v2H73izlK2S1YIi7AyaycpQMY54jZsp
VU+tCJCAxUTwON9ir/xGgX2Imj8njsXeygEqBL/TwEN3WMCrxBqEYigo5LXeqzfG
Fri5QiDS3HcrdUEFF6H5kBtP2wIpii3Sq7CSNkpPQZrUNDSQ1CDIB8gwIxW1kqDv
AlaNVlEmMp7j1oAbs1V6cl8SSLlLqA7ZaREn+STRVaniDoJmgQvtWkpRiOJe1HE7
mf3/82UUBLXupbF95iBDKL3j3i5zpdH2f1MlcBVLYpc0H93x/kguu7+25v5v5hKk
ruo65g51bH5TQrlG6Fb8AtENqzr4dwq2Skx4j8f2rLGBveuhhUb5hioqdWc7Syf9
1F44F6lCnIVpOAe3QqAlbut5eE9zrmhwbQuJR28wnKKrkeozSg9BvlQyrMU5/oAw
e1lQZmajle7/74dUKgHolXAHoSyzfgnfZhwduad5rX1aosrUs4XFmQr7qceVYFAm
ujlYsXeO48pOZi56AB2bE8eb4elYAoXQu7I9+sJIejIL/AHs9nzfZLpob1X4iU19
c3z2hnlmbYkxq23RQKEsKUQkgMWrArCD243ZxGIW3aLwQldv42FpTzf/sOkbPNw+
c1dNZmFKxdDcBUV2FE0fCikuM3JVLygG7BX/5bUFbo7AvD61vBJJUQJl0WXeCSeV
sfd+h2S91W+1ZYR05JaJ1KLWxMjlL3fzI3y7W0exkLxyb9VbVEeGp5cIl5AysNl7
vbUQJyxuN50RsxcZGE9S7EEWwKTF1ZLfXhPRk59gdAnjNEapakEHw2ASixl+JoKu
RJRHtBk2o9yr9mpWVqe6nVK6TKsoFlydMYYVVuLNzepceTR3WLeN+uTyLEZvSttN
9MdoXE+aDCc2ERtL1pob9ZvzXhj6n6dKiug4Td3b58s2J65z7av/4AIfszrDTEZG
t6CDHZGmOLVNRKpNDpZv262leKz6ESifO3FIo0DWghjSwB4m5TTuEI1NuzOQqTXF
crAm381j1+UcibpAYtlVPLWdQCqNsnx7pSzjthqDp/ZfWGhB3ZkyThbtaXcXHlh+
8lQRyZJIBPEsvAKlpoU1Z1hn/2dmQ4F7sJmXTtIjBHjQbR7JLImFmOzFDT/7XMCR
P8E5EbCH8T/qxtPjFEgvEMbI2Hx6D4rLmH4hfbSY+Eb+QNDPRJDszC1SPm8wBDY2
5281dhXCRQuTn8ey4+Sayunn6JpFITK9BdB0A5p6PCtizza0lxoRNvRHwyFRf04p
j4ujA2LlEPrinTGV3fbtceCC5gdVWzXMx84fm34amvrEgnFPl/WYMEIBuYPqran/
o6Vtlvx+OZRRJqgHRhuWj/DUaOBo1nCDLFnGPEKBsojRpyIUQwPks1CsPVOvtxET
g62rIwSl0htrBog4YDgdyn5WA3qo1MOD50QS50UFqvtF0F/00pItZCbXsR3sOpQC
uFh3A5pbsyYnHpCP7/IX/tVRDvxdqFuHeAUaEF8nh0syY+onqMDatJfXeFFNBrSb
Iz+45/OxwzY1Pu4AIWWJAHYbVIT1WHT4A13PPbfYoThBEwW3vhoQsg/MTf7IfU6k
jdVMB/ffOdE7RjYQWEWYTDF+bMEyyhZ4aVXCxkxDsQa6z/+6vsLtQYGTkGUgeXGw
UBCiOa+CVwp415vz4VPyDrEF2ItXayS2NsgJZfCBjmqjHEjMFnlf9POoJzdM5iwo
0ymQgUivMudhZDuUQIGQzjKb5hTTzfI3pzjHYH18FB9QcSMZ7ZyQAE+gBO3Xs5BD
PhxQcQV5/FdDRupEmbnRtulcv9ol773569PhHYwN14770deZkPjSzzgHh/osegde
2P9yYgoxLOr335/C6KOAUoYr4bezSzKRHafWfXvpDIIxLKFY1Nnn4e3rfJQ3Y46I
oL4OxXQp5DsLkKed0msvjIjAUJRs31B1w8L+BuB/VwJoVT502r+MN3Ggjh07JFBF
FnD4iSSdDR9WwBKZKB6cEyxT6GI7nQk30H0w9T8jtpFxyu4Coo7zFooiXnIF+uP+
tOXZYV78bkqbAof7O0Cof7v4jDREXxp8WrUOm7fQbzo//P4TjMVmwfAokvPf/04m
X6HRCp6noIdudp7LSKjLsBuHNwSc2QDca+hpJrndA4lsouKbgX1hWsLStocdO9Wb
LY1OpJJDA+sGBv7rUW0RlnBba3C1fSxV7act52m/q7YY1j94hf+4ZmcDkiCsqpEy
dpMOfne3Gsm3KDXBLJfKdmnfgA8h8Go1sW54utW7kxmroPXlV8JIlsrqM3CWB87N
TgzHHBgE+kmi3dVQWjcqysS318kdztOZf7iesU0YzHNko2i1YIwH68HFO2US5jCZ
6CSMRNdH+niquPyEX55gHGu9CkAfa4mopV2ILrlMcTxiWufjDUY71A+FGXM3lz2L
qNOEVe0vUVqQTYzd2/FHB3acz+jopd0m3XL+KPxk1X+hPHVVkdTPpigwLlr3UoDG
t9WUJawJRAlg5nmgFyFJfUCxTKFhJ5ddFUGYR81FEvC7iJ72SgsDFxjvToXMa2CS
0eaIXFR8KTdouWaNEbiHgF2lOFvKicJIEDfKHQjuLztb2SKUAHCzEHvMcZGm+ZEv
XhIBBYZq10GsWUEQ6kiAqS6+ESLoLtvZzK+cVlLMWTCudXQq3De+kb2WRG2BSgFT
QmdcPbT9+519LVIWrkDeOBvlVj/qjtapBV9GACJb1dg2h2ON2sab7VRcbxDK+LHL
ttUlnampqbIO2b8KlkbBNTMjwykonW2GoYnbt/oOgahn/1z0lmVrplyf2KQAcMCt
eip0JLmj/O7IGMxIiSIGt7gfjvZzKtFJFdGrOW3FfrgVXxkcOB4hxIRNuUmOW9S0
tp2YvdMliKyZR26IBoSi1Q2KF3aOYqVxbsv/GuFmGMzOaTRKLV0drY8+5L4TJRxk
psTE0OnIhfabSIWpNDs0rLtG28IiW6K478eoF3E/8za21dEEqXn2buG/BDxyH+/0
wAiwa9TvJ0HgzTuCGjVq3/KJ7LPQRWHUSgdNjIW3MsagRPH3ep9yZax6cxrMOZhV
K77lIwqJBew01h8ppzfZqOQV185UGLYC5gCAw9zM+WV7Do3rt2quKkZJvtsX2mu2
WeIGMZp66H61fiexyRqXxQ8wFjM/xBa3snUMUbP5DqOKIhdYCcOTYafsQzsC7heT
IskTFvmyscDHupsciU8bgVTJKH5s4SLPrPkk7sl64k9qpU7x7/U/UyLjm3hzLLqp
DyMUuyUlKc6+RrgOmuc6pAFbdp095YqM9IRnJnzm0TQgppFpDz4PxyCMvU2AiGur
AjDCSdxWNWkcfCNVO4a1T9bsiysfvsyvU5WtwiJTtrl4VzkuPIYFshwG9+ANEJPe
NQvdhmCwhYWtW3pGXYSc35VzHVrAwCx78gdPmWU+ErP2ZreIj7vy1vVBGIOpeXHP
M+qhRk9gGbzK/WgFU5eyN6mTz/XnyduQTYmHlhNqnzASkQcxCzScAneNpQCueg+s
U6Rf22Dap8CjfKsPv38p2Bx1MccqmKOu22AFELqsDaCib27V9vJFN5WzVjr6kK3k
BTlZF5tH08goRIYV3JhxZNAl6mQK2FZ8TSE1meSl/cxDzPryFs8x5Q0iMMsBgYfb
KMe4YRwK1wKllksW1GEjeYK1zMpBrY5lu7ZL1Fh4V+OWiixetBfW/AEzTMUeADeV
8HWy4q9tDHsZx/xTLZQjvYaNZEMAbyC6yuEm0TE+EFptMvb4xoH1AJ7sFG/N6Myp
wIjIuKwdWkDDLUhsBR0Oj/1vNjEau9upncvu2HiVzrWJPGwclo2pum9EpkuoDhQN
1WInSIKtldFh4fGy4l/P82EE8KdSjAsRN71BrreX2uLT+fxCt6/WUP0o4V03wFMp
NQriKVxGuTtEA60YG/KxUcKGRo6KXFsgK381D+jKp24sOIxXdPatkyq+BDFDhg2H
f0Mu3Y87NJVrkZTypJ3VStnx8VqWJRJ70mvf79bulW4h8T1US46u4o/z9tESIT0P
iPg1FivikNQ47on+5sLb7x1OBrAt7GnbxM5WHY/G8y8ixKXLva8OgjwgbNrTYFIW
tIRsyQSx3IMv/y4FLnplEoIF9mZYNrLb+RLG8Douq3b+khbLoYDpeoFU9h8KPuT1
41I1RqS3cm1grtWAJ9/koQYvRtkmBqYXBw1s+MDlht1gLuNIta/r/QRwnsz3R//k
HKSs6bJG9Z9mIHy4eZ9nWVN7av/y1psnaxOrQJzfnkgd2aGr/BlJks13QTCdQUU2
vCjnO0ifnrB9J5UX/h+NXbF5w12RifNzGT+7tlPVYDbmQEP6RpSjLTUpzbJLy/Qc
jqBZPe21Dt90nP9K4ZkAL4X0I95C6ppUB1LhSMCz1/9jdPkZs4KDhnFf+Uia95PU
4CBzeTk/5dl9NQl2LKPi0IEz/TT/+IARRhyvQ7391+Shz4+hOeVQCjU5CRBl2NMm
fYQT3Wthm2MO8A3y1oViQMTJaKioIjCO/rxFuNsc7BoSFAQ769ttb+glNXldRKYx
Tvxd5W/wAWexgS0ZFjSerWebE5goz4foqrX1aF6T26GWRyN1hasZDOXNY3VhRBUh
dXgjwacCGpOYtkkRT8nWRbYaHQekF2yoMNYme7+RTxSCsp7EAK6ZuzGFS+bpDhie
gXlXyBqfv0W86FxiRPprV7qoyHWEsh+8ayDxHQftKUlKFNs/avDd7nnuI8PxyHn7
pAUx97CdtqfzYGdvnOj/FP797Ax+6JGLR8UIMP+/+Jkw69sIfd2s6SFJl+UKuAtX
2YJWTCbYCVxGkUDJ+TVbTQCpeztNOYe5+nNQQzvVkCoA0Ay3kLnWS86iGoG0GTDH
Zb7nV0ccPlbkEmfUckPa3/nnXg29+MeW9iC7MEYyJDWC+buE2ds+1NLaPKCcq31O
7sXsHgRHdEVbIfB/gxJOnkc4lDBL1ZdrHOWRsStKIYxmkB60kWLNVKt64TPTWUp+
+xnnhL9Y5a4IZqHgWPG0kPbnrCWtXwdzD2uqqOvzoWao1fH0hzdZ4kJgWDIdkKpv
09+0W7TuN0vsqDQxnbDS0rAjJN+9B5a1fp9teB29Eaib0TnexCESgmvZzHf3+71/
gPwgRwzIlSQpITAfDODUW7hI2WkZA+hjzo189w5YSBA5qkie7IU++RpeWqFRLp3Q
CEtTtrQXnADIkM5xtxLyoZj5sTtaQpaiNDoKKz5Xsygzv5idlkrVxDNOb/imigcJ
gWYcfwhzoRzA1wlw9AeidtV1CkhWvBdwt0Kw4xIStyG8rPt5YgAn0rYsy1aO5Zdx
lq6rWA5W+9IMbdJvgAqBrm9T6F3npxzQvYj+2c2T4WbafvzI68slTX9WW8eps0Xx
kCMvUS5bLp8NQBHy0SMUsaSUtmQOypQYqs6+13yezCwY1qLapIfe8JIV7YQACNBr
uBpYhI43mdf2ydtLmsknpm0ov1pmaUhxMznY/6uKr/Zj484cAzK0jIwWEbmxrDYv
PiwBwr1yR6y6BIUxPcd4c+OZr4CEqyzHDVY7kUoRLg6ayR4cu77LZWQOSnuBhsqu
ojovs/z1jsagEn+kPfQ9aPGB0LZivg8Uu6zECLV7yIOUpjEZTnAFYcEd80QKXBxm
SXxoQfsEIgl0vcWt0OpN6nCPCXbsnJZrFwXnk9NnoakijdVDjG02NRO4iyHbrX2H
9NoDo0J3SHDb1SJGVuNH4nqEzTIS+QMsF7dbsp6noPoQsmJgysqWBKmGQp+N0iCz
qFE9He+UbevPOw72AjBpxxQY8Ir4KjGknXpZRMSCMU1BuLv5XWlnEsyO/pi0hOvo
TDgNbUrvbEhKbBXHwJkktJ1ZbYIJMruudVb5ShlKO5JOxNa26BIyxLg64kI9D3/a
LSSMHqbezJvQWl0tbeeU7ofw2o+mA4g/rnVwoUxIdxVLKrgyf2zkubwOSANrKt9b
2ElfaaLSdxe/m0N172BN+/5ETAhrVUpfnKgygj9f1Brbvs5GNq68suM50FzNoSz+
D38xrVoOntmp/Uea7jeD+0B8+fTg/NPEb1rhAz4SjbwElJyerbBK+xCqgVMd9j2g
s5eSlUtKwxyiYU57eBuNTekEYDefkQt5Ns9a7PpF8VdSg/OdaUw0JJkch7Y55MsV
Eelz8MO62lSEy3rkJwhx/tFDMIWU66rOwSTuNPK0SKx1XJ4EcUtUUwLGOPM16ZUY
Ap7/WRk8uZNRxGahtjuQ+DTs5dCVXVo0mKufZ8lune9ZnHQy6ZLnrHPsDdAkfStG
UakIUv+KutaP/kuV7dl7I7IvOXxnkVygTPvPUPZx5oBsOoK2nBDrOQyLQalMRP1j
uqFYBFnLgIXfbapNHc4ifnQuc9zU/x8IgmNCYaYpxagjEGYd3Blx3zYC65glBRN4
og5PWUvtS/A1WL3cYaF2oQOU9MvlWJTqWBDHLX/4AwQaAXOo0FavHD+zv+RTAJd6
meZeNlCmdmkZqBXSaLrU+F1smM4nkSWfk9zBaeKt15MS4hmUQalbracaB4F7Vr+v
X0VMsEJF3fiIvdG3F9mNHM9E2TpBbYnkXpQx0aJ1b1RAVT9nWJipKaCxc+dVybMc
XPO6A0wsxfErl5McBV6f8hXATSPUhd6kVitvuqnVfQQBoXnMCnPoeeO2drXSpmk5
CPwh6f8zrPMd+eGVYCfUGlmKTRgX5Ziu6hpp7WthOPIVYGc7LguM3xvw8jPYT52m
6sYl1Wh4mPEyOi+YjEjYiZCHlJg2cV7d3ahlZaOyy8lShFSFODOhjXpopx8d7CEf
dCm7C/jfsRTG38EYhlfbgXy1brV6wi/MNtv8tIeepliIF7XztOG/7LYIdhjoDL+R
s+YBel2pA9yEX4cHRaLQZwJm8EI8b+E8k+38LP9UJWkqFmZlU7FpyM7/JLtdcw8U
Vha28pgrI32KqVtOwY8eF8LkxEoYfQsVjuWW8f+DNYsuz+NInIYGLhdz3EtcRSW0
hCrJjatea95kYGMoQPDxtABm71wi7X5WmosD6KKJu/5/4LSAn1YXufqf9bsRne19
pe5JKLPHAT1vWtKbxRo8Ulups3TLk6ba625bWD6caw76nG8eEHmJW1F9jriL/GrJ
qzHZ96Ib+X+SAi8CrzfwG14T6cmN3TI8Vu4rlwfQhAebbIydkKXYnH9qBU4sKG8Q
rVh6XtoLB2arKAVgrVKkHn2vFxRQRsby+3cexcGZLKesyR41aauEQ7R9hFWAV5Ld
73ZQ96iKZxU47VBv542URd9QBJsCy+c/oATz9FkZt7+dLQYCt2eF3Lw7tNtKF5ow
SpEJsO0xit827xHNSITbohgIXoKAP3hkhKqJF7oyi6J6Tj1AiMXCbXKwv72CLwGx
3XERdT4UolBE6TzpWUg/4AbpGEZs9T8K+3B6kj4d+/kIPfSmmP6e971q/vMP6Bq2
raP4x0CliI06XMardUWJdjQCz+fawlj3zdTaLcC+o0bGzcR1aCIZEMZwVc12Njbz
7qAt2lL6fr6sQ6vsfjx4T8dg7vM0VZrHBCFaFyU/kW1+TNTuAR7gqoWxguJYBYjI
wIYifHoF/qrX5ZDc4TuHSIaz4diMjQj9jpeRAeWsqfpAS7FvzzqulYv8JfhqsEri
MSs3AoFifCeL87JyLPAIYp6mS2ulW8+PY+V4Tz4u0tg5S9klvE48bQUuvMFDulFG
UBxud3c/yIUF2ayYVNRTya6jnfqztFzf0c18KlLYza/BzUsOz5BIQq+JsP5ggfuX
22IjkZwAsR0X4ox0Z4yF/0+hMSstHE6h3A7FfaC8tiVIN62lP7DAgh9RQWipUNEe
lXTL5aYBwh6VN88Rn89pKm8XW2ol5fpCB2UzgZA+w6dYZLkFwZOqau7Z3PbUuG8z
F6g4kITh2peXnebZhIH/FkMdF8PJh8AtdCTrraoSRVQHJ3tBYBIPuJF3jmU5hfv7
TQerXjlOWHOWYDcRDdojtXDYMvvF7zS1kQVZ/QWuMqRQmhajaWtre4e1hzJwCo6K
I45Pxx/u+zkZ4Wzb2Hq25RCHctnhGd+SEWrCu89OC4cQBEj9nXbid8S+GbUerSry
uLs6ynGyeHWAy5mDNrVnEHAewBtRXtYMMchfjYhj1VdWEHifvXcicH8+nJHtrTnJ
WsliM+o/L5L5ZtF7D4MI6WKuGuuBeLZ/5HaQk4cnissWMxZeY8H0BE30yE1xp7CV
EPMg0UAhLoIN+DFtP6yrL/2r1wLP8CdiNemE3pNLyuCuNmAjQi9lQmwaTEL5HpZr
fVr///EFlodRU53OMl55GbQQVQlCV/TknrroRzSskX/ri4cJW2IZL96wXEBkZQeK
l0Dzs9dHm5Fl8eAW+bRw5caKzrCLX0hvdq/xT/S2bQqAjIQgWLc8m/rIapwjFdLs
+GezpQ8gAbgCdtrk7E9UXOGsZt5RcY/d0VYBCTsc4TAafg6HGKsbKb6oLugIis/x
iiViHGGzcMwG4//klQsvVWpCY+FLKtYMwNymNp9sE/59XbQchqSf0fHPwSCFnrW1
COuM1BdWxic/3qwvtN2kj07XEDfJS2gE3AWoPI9028NjILz00xHU79LEdYFAFu+Q
taMbj0GYuA5CZDdtXNKILFW2C6Panp39rWIb6To8BPcQm3pIdLfWAojxKoh1ZU+g
D0dsLXvZKrDqrgRNOqB+ThjzqUOYiYFAiTN8ra9e0y0M2Y3EJDxNBMm4tmAy7lNm
jsKNojaq192Zt7yo4jPNWK/1MYLz2TzLlmKTBtV9cW2UDTJ1sGYK1eoBDXV2QGek
JLym8MCsCD625bSaMFJBjZ1pnVEjWZibeybWBoY9u/p+0QFLJsahkLsM24kl7w/C
iub1SSR1ObQL/OTHu6dDlb5kDOA0/bjT/epcxqlcVx8XIS0/9wu3mvN7epOf8HQR
z06YPJrwQahyXkSA2gRt4NzQgGb77wrG8mrqEG4ZXm0SrgOzx4K2ESd4hgxF6qvM
mZcGGj5TtYyA8u3iA2hOCy4UdoZYhcalrcIUDWzHXHGfyAPSrxCjwIokFmV7wK/q
s6FXnbzgWyXWb+8uD9FcJZhQkoVn311uGY6ErKDXeB6gDP2HTABqxztUmi6hZdP+
tUet7hJbcjyRgD6pi2OShuVQa3p8k07UpARs5uRZIyh1Jny4FEeR210Y1d+j1IJB
Nlv1n7Bf5AVFITk7IGwHomkveSOJL9S8MEaP+JTViey3xLMkr6ltVFsX3Zvit2SH
flGJVmDlqMuZub6pmpw3U7/rJyN3P+DxTwjRJM2/bqhyoXvYLDkOhPqf0nDmnyQO
bY3rfoI21kT1p6dSAK8ZbA2ZyT3Cd49EVHIFTRK7DyZAnVWaMOI6mXU76ylEMnhd
vC90HU/XbVtzxEP+f6YJ+THokX0ey1sk5mCoEGy49xIII2vL7NzTW+IXwOy5ul1f
FeDXOo8ADW9i64VNJ61Yxv12lhTJTcgYZkeW/53aWnx/2eSS8D1E+1xRLMWT3Wna
PIJ/hzZO9C25HtHFQqfXUFSOgK70oIJJBMe0Tu3NEeDYDXNKCuwkuZIPfc8gtbWN
Onu7sxsuuQe2NdzDV1yimcduQZhGEZViq4laiYvGtlCYz3y60AEIz5v0NRiyFU73
4hkoYjLUVEYxfyK+6qy72I7o8cQbmIXKPtmefafoM4zgxVdbrjFw8zEl8TJeG9sF
LTosFb6YDNgGz7peSOrxBKr8GPYx/0eCHlh3cFiNSIPFOg/NWr1BZMWpQWSwWrmO
tO6zS0ctLtRH2rvM2mPOZb9uLPuaJvFL9DHIcEOE4HN7/fFZ5FSEde13NdNHEsOg
zpCGcl3r+SmaKwpOv7eVv0bukoevHWBnvz6luJ4r4Is5MCEDhs+Ll3Q+Qj2Bi8o6
mApmxWuRtp0rJIY++UtgS9K2vkH7CwdMwkiYOqBi/omSfB7YgI8tXIkOkg3+pe6J
tZXW4p0fxsontziQMYipprHXxYZhQj/dqRPHAqwujGKc9CT2Y5CtKpDWC+0jSxq1
sAXkaVzKywaLyBMvr+jTB/ztQig9ZJzyl+SxJY/tf/oG27QzSo2flDKawFj4iuyz
+y44GecX6ydeTfWoFTGdRHZ2kU3mBbYW6hxNcVMWNio7Qeh6zg/kicqBaWTSqyXa
xwi3gB3X2nrCN1oyMyjrRnZivULSQWMNAVQdPIjMKlCn6DnRQJVSGF5RDlCVCJqW
J5FL0CsLJgHipVM6eaNVoMQzl5yEnNg2Z3I0fHsClRzDA/jG5a4EwoKlfD6prr0a
NVY+fvxCPVzcEQ8wugbVdbEtUIBACOPcc7+bUkrsKDJaWmM7HFNdBD/UaakJQXdF
ROvvYI8TpSXLlK4g+QNX/cOMY47CepLhfStEKbWmvyF1T2ZB6D7JQwISllqpZoRR
kk94G+PcD/Fqmu6Os9TtzL9YazsFoLsbywSErP9bzZ283L3ocBU6T+FanwQmSgmS
GFFXRDyJbeIjV4k0aswgaYJ2v6T95yWp9qazXTPNq6tleMqFZrQs7MyHFKLUiDiL
/VkDn7fPpjp+5jDbGS5EhZntf9gQIou3A1hH39H1KtF35u2gDcnMJarRhuyrFHNN
Hrd/Niv4NSiq9hBtCP3jYqZP1B+03+heFPdYrqKhG67aBUJnNgWU5mcLqVTvY5HE
kw/eybQTjzPJIWoiNts1hD7U4QRzucQdZmxRW1HkPHh8k4N7WSS1eS3LDFQse0vc
aDpqBnbcsMLzsbH/nKqTAkBhNLuqjdCCRUoYYv6JSPZusvDly+xNCi7lfDzerLkv
aCJr9JbWwx8YXLw75gGikPpJKjg14ayAkv9rAix6NSIorWEiE64XXZb6GRUg4TF4
ubqltaa+rkVquusaJlpN1dF8DYEMBy2zQvYx/y4gO/bdXDXiqKD/VcWRJvJMSFln
s6PEnhGrs6WUXVLHb9GzL59v8brAWzDqxC4RX6/WynBZpjAhqGg19conMTZPOAqZ
GcXitEyOa6pqWA0wFmqLQ/P4mcsRnXybOI4izoc1SJ94E+/xKev86hTjjmbVkD57
O+3Znr1gyDOsDgPkCTrlujdwKU/mfylbu/CqGOPjjMMXalmIwS+xqjIYhaNbSjFZ
5QNWIrRrByYAJo5A7eITdbaYJerX12VzEZTVgm4J+sRky/PjJ/RTt//tJS2DW6JK
83nr0aIqJ1vqNnOD5qboNmqtIgMEPAP86ZYdQ8lmj9bw/oj9IMW9OFp1OVWwaN3y
udz31/dIu5LK6vquEmXI6PhJH9IJiJPZUdnGGPgVrGQuI8jt25rBbJMR4EG9m2Kr
HVv6pExwoEqh3FKcgSFQhzQgnBaPdKk3E0ToPlkrVo4SiDyWixRsqUGal3cN77+G
xCLeA8iYiI4BWbiFp7PktDRpUXcGWfQ1AnzVfOGSgfkhOQYKQWGsvEaCi6LrWSfn
8U1UZ2mQDWW/UeoG/+QMaIcf/8SgLqxH84FqsAubvKCtj1sD6Kp5JaJ8biDgZixU
rgDfxCYjGnnDSWYtH9LElcGQWJsAA/IGBmJ35fAEYigDSPuEUaxcsPuRNgzMnk/j
GyyM8MAmd0L+sGOfyz6gO/aVZceSTRG82BFDUj10TGBR28JTX0v79SI3AEBfi0QA
4LL5oSAEFHaGAWpzkuSkwXmcNnB4zY6XFoCRROSw7skl3iAidShn7eEsplO8mYUq
u30HUnMOrlGbmiNzrxOCgP1fh5FUOyAOxKhlIvrS+3u8iNl8SWsQwJNe92UXqrey
sPvFwVnXCXvvW9SHNAXJbWlZ53iHC+JCpyaDiZc7XxLPnP81+CmCqcJ+BDPo7dsB
lw68yOc6jSELYbHqw+9u6aaWYh/wmwBSFJoZpfdLi9rWXz4W09XknyWR/VJtX7PF
zTB3Ww4/V6c4i0QRpt+y3letmvbm/DgBuVHAC8YRPoxPxh3KWdFsZZN+wM032ASc
iC5F0um2vwZfr5hoAE7TgKHKf+1V8+t6nHxIg/u0X6R5p9JATv86smLLhz3oXpRP
n1DkuzAHVnxnA8iSYes3xC82Wi8rfpf1XG1FdIUcyEDiBYUNBeaAlmudhp1ryg35
GF8c+HS+b0g8gjPZ3JNRMapNed+9D3D66PCKKGIxp/SlSRFK/4oAD/mOXKFYCE7+
mEEvyAs2NpxB+82qORPxnJCyUxhvzycTUb2PR84/fODEZnDt89ZsjhgKKwzbtHfx
aYdAcVJP84rn6v3HWeO2abVIvvZEoynk0eEMX48ZrU8W6I68Hvfc0gDmopX2pqEy
Zr3vsyKQDulrp3hMD7ODxUbF1gfTdqPhYNgGjVAf4R1o/8C2h6YyEgNi6nU2EcEV
ZISOjGwZxEf8oVrzrlyTGMEijAWJcXQ8eqgbPSDmJ8SEF0vbzfbMBl5fbBdMWlbG
xu7x6C0T6fZNxtu84mP7/uJd9yIULTssXDEmZR5M0nR/V0StqjWqVZofmc5fBisp
K9Hk1AqEWeMPxwMSDA5HDsSRWz0R7l/yEmvI5xyOSXxgHIiTzFOwh+eQqDjjJhpV
dyvEgTpcgUWkknXSxZxtUeaiChltHIN4YLnwTzdMLJ4vQPNgpbNWZovORloeHbOl
AVRHIbbuHL9iPvuQeInj6AoWkx4DC0eQktNrWsv0nnpevtAl7z+KvEoHo7D9BESr
lmA8EGGNOhl4NEQX+DQ6Qx1SV1e1kvy09w/rVtczHT98Dp7Be6VKceFEnxN4UwxX
BxRmYodRp1ogNak3ZFzV9iKxxBrBmhTjbsv5JqvaC2vwLCEzKh93QxdQ4p0uR02D
ZAxFK1CjtHtXGWldnDqRm1cavxv5Lv5nzeetmUnqQir/YbGPqkPpPltfN89Ej0yB
NcXtfkaErAqNO+wO/2iNIOhwy85SzdpGtHi03Lc+gECA8RaqC9aYa/Iy3SDPQIAZ
2ctJ2JkIEzzY9SWeF1KylGrwJg5hyKSDCr6EJ9jZty/R5A2FeqQ/WARP7dHXQicT
IKFIvBBMQqXKJAjCYDzuxX02+GDc0EsKY4B4SsvLPNBQFaZ7hOipZ2aRm3VO2PKo
EEA6WuMmXSKXPAfVMrleoVKttTsguAS0pCGIZAkirDHz+qznSG//zZQTkOeNOaPf
5hX78mWuLDqQkQfUxMeCd2P6VbscvoU1MPXLlbDZk8uGMrUHXFsKiHk8xgIo3m3u
6o/j5n55XT1B6+m1cbZNBbRaLfuF4P166VVHWKnvVoUyfBhn6CYn0R9U4aEHn1ih
e0cha8GKM+9ZLCpfYhap0zchmKEjeXaELQQB8Wo/KH4CJCxD9EbXbfrI7SsNPmPk
4VDT/Bq6DJIRw8iNKsBGsRZJWLIw6DgKlY5sWPFqijELobq5Wy7u1qfsqmnSdT74
nZtWPcx3AqdAkcUMvfcpMTdjyiyCUadmoB7eTMXWxsFpxCXohE9NNRoo/cYdcaGa
sN2BOE468HZy30YtFmgz92OmELyx0OluCL+WtvEyropzTRGtm5G/RD+1yXx2QNqJ
+z61H6zRwvrgdk9fxgdqD6BJ6jYGzVEXgucJrVDAklNw/w4IJPb/7mZ6YKdnLrgg
9/c6cegNmnZraLyteG0oxWZxslLooN+HKNazlPRQK8HCOl+bMiWwPAh4le8CZoZK
1/gqWR2+xzvdPjZhZXYR76iMI0SyT0zBaxZnp1r1scjELinyj7EBOW8WmkE8Y23V
xaa/TabRbBSeSttzHzADU+WAx7o7dofIfyHlYmk5FuAXJxvDNyo8Fv179k3l7Ocq
T7K112WSFEFBTzTQu5cap3kQkwsBoG6EwaTSlpA8swXorgqbXbP7bwRWnSh/y1uO
MZA6lLTi3dfJOQTZyh5Fb4NlJgJK1m2hRB/4XC/ZH8NIXFHQmXWfkJxMkgPqdYus
GXQ0gjOmNpupt5kA5edo+btYZzm9X8LioMvc0S9OaJ0ptYsaStACMErPPoKOrY+J
0WkHDvoZK/DVAiMr81wd6rzKkexgShGcABeD2TPeNcRisSNs5F15OCqXQT/+2v0V
QSwxyIt6vk1SbzpL3nExqWY+C9Ykjlk06WZd1Gv2V3D+iDzOULjvDPsGfhbnn2UD
k/16kmn6KqDJKdC/lB3aYNrnFnvIffB0QnBfgDBGF+9ojuaYGR9tLidMR1BKLrID
6mDRooLsrMQxW2iqVZrTlOMSjDnEH8TVQLUOrDb0efj6A2gMrgShedNJSRBc6vbG
23mkwQu1910mP4mqgjW9R4xQCdJs88oONsfDjpxfyefjcKqTPGSYnvIk9y2yYxHB
Oa7ttw6B8vAvU+WBcVhwAzj6DMdDQt0k0T7fV4d70MDCf/oYanGGbQBFH9od0ywT
J+IZf9qRk64LzByfqH04iALmosBTYoQ1Ehv7sF3Vs6x+n47MvZMztNMbOM+VxLma
LMrq5BHTcyqOybDj18Aci2dqCZT9UOXA/hvQdbpGjVKKORns4ljQejjDZRQ3X/fC
hvRLYzZ99YXW8I9V0m+lGJ7uTx7J//R/7oP3t8Pm3s+oPR3of0fGLqxSlsHVU8zn
nsY2N+jTk2FNWhA3DxxZhGu1CnLGkoy6qe/+nJTY7O4L6iUSXyeNMvarh/EsaZoJ
40wZEmK0SM2My8+yaiZ4iVFYKsCFBdpCBp1gnCj+A1Uy01omvWyD7rMJ1bsmbxZJ
dCUXLDD/9ngmh63QE3M6mqnRCfRZYRnR24UGU+UdSlgqarcJBaXy+HjJOxhijgk6
XgOAIQ/6G0JT8aHnqY+gJp7OTT/FkvGaLmAIiKXVQI36qwiWlqVehzXFmhEdZU3H
IxlRV4xKSN47zZAGMj/9noka8XJTTO8qUPsmv6YqxDDDzlSElTZwhsdl1BYPD5GZ
7VtqcOrlp3qf4uf4uw05P4Zhvx8CKqCAowyl71kh0/AquGdkKrU1y/00AETKcbSF
GfX2BcJM4mJSUKGGOGWIV0tGdRO7+5iCPUXDyqbGQ28USPPM0wQNMZjMdDQ6hnwX
1LQTyEtI4ahhYsi/lB3W20XphdapAbRaOK2c6p+vva522an1SV8JCJg2lkH7pN1k
XNoECqNTJZsPrxvLwO7Mn4cLvKqGfw4Elfehpm6a7f3W/FBlOTFGclNHp3VMLbZx
tKS2MRICrmQJnlikH3onMOpMH32wiJ5iSZogDtfymsryw2YEEig/QW5z2mPLGoxY
+veEGWh2A9AW8sJe+Vf5XD5cH7OGylqZlof2dIf5rrbhDVZOGudxzhTrBHf5LwML
R0lDSORKGVU9KV91Lwl/KpMTzOJQ+JNfzIgUSxGCzZm4Fs/UNT97HLnuqkExLkB3
im5U9jG7yzu8Tv5Y8rmjx8zz6C1UHe4w2pf/jX1ie+Y7+lNSZjPoIS4GBTtpqMLv
ZO07O+am8CbwTA78CckG27H3XR10tISQ74FZFOqU2UyPleqtdy4bAfgSpORpyhj+
5KzfhzsILFb+RhMtItueu3HnM040VytC5En4qpDeN8Irpxyq3VjnQ1/FW2/qjN25
E12FPi/Vc8L/7+uY1V/9tWcUHzx/1fYANxdlCyAEczV0q81xFigWprA00sLNSc/x
ZKX2wuQSsQD33YVq3yskcR33RscCZrXzaC9PCU9pgo9OCZirhZUVGGAcL0dR1Zhq
JUHHFGft8vAPnZjBhcZ7uyV0aMp0YKj3m5fg0c+qUVzLbh8lAKuZ3QTzh6p6VEUd
WW5X39MQj2RmTFZra0WhqIY5v+uFuJCDeuO4npHdDHhc7B939BjpL8dxDwW0+j3/
Y7OmxzTtf4gyC5O/TJlbY9sxBF8MB2uggxdBh7iZQsK5/7uR0xFr3nHo+4TM8djY
4Am33aocU8LiuYEY2g69kFpBFsk5Hf7byvhATnRFrnFex/4TMEMNz8yuQW89ygqy
yruqOdgamHhT0Kp8nfqzhF2e8wJpc/lQXm5cNXoZrgOFn8msYEKO9EietL46WnzA
UWxGunjXHGPjAAx3gW7mDoZFcL1yua83NeCz2Rl9YNzx2P1RhTaGw8fAvxEWX5nK
8TPce4BNdzxDTx/0BkKtifWa2o92YAsc/p1yeF4A7KcX4pB+hpn7LRTfo3Mj3xJp
18irVovHcFuG2eEkgqVnwrd00vN069d2SZELnyRognn4j/MYRdqt+g4sl1XV2KCF
cuJHxD5/VNEyKUi3Avj2bVWm5V3m9AKFxRdmyBg4x1YJ+/9X2cXydhOaTsAedqHL
6siN+3cbPeQgbDNDHqMnDroHVXJyp36B2q9Nh9w+ECBX959HxEv0DpCM8/N32qv1
xtS5JdacQyoXAvqwDfWFW2PIpu4bRs6VjJo5YKIqnerUfCe07xKZB76x9Hpd4F7V
UhjkS8IvEqIef/4H7Lni+BVMwaSQti/Hwcj5D7tkt9M=

`pragma protect end_protected
