// altecc_dec_latency1.v

// Generated using ACDS version 22.3 104

`timescale 1 ps / 1 ps
module altecc_dec_latency1 (
		input  wire [71:0] data,          //          data.data
		output wire [63:0] q,             //             q.q
		output wire        err_corrected, // err_corrected.err_corrected
		output wire        err_detected,  //  err_detected.err_detected
		output wire        err_fatal,     //     err_fatal.err_fatal
		output wire        syn_e,         //         syn_e.syn_e
		input  wire        clock          //         clock.clock
	);

	altecc_dec_latency1_altecc_1910_lizxuqi altecc_0 (
		.data          (data),          //   input,  width = 72,          data.data
		.q             (q),             //  output,  width = 64,             q.q
		.err_corrected (err_corrected), //  output,   width = 1, err_corrected.err_corrected
		.err_detected  (err_detected),  //  output,   width = 1,  err_detected.err_detected
		.err_fatal     (err_fatal),     //  output,   width = 1,     err_fatal.err_fatal
		.syn_e         (syn_e),         //  output,   width = 1,         syn_e.syn_e
		.clock         (clock)          //   input,   width = 1,         clock.clock
	);

endmodule
