// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
w/Yrjwx1J2BrlvAqrUDEpA2v6rkNKpK6TnOXQPlboIhKPrHKGckD8LfTGGO+
SNI4RqjbM2APNT785GuSOgCxLLnFvLLxOroDAlDxLxtjkRq8VrzpXLDjWMKD
7/7Gjm03xI37yh+q+4B9MyQRv2xfQfQUmNRbupDX8x//57VEhEuCBtcKQBho
XKujsoHdf75FHAsz1GnyQQmmXvvMgKo4yLfJiip8sJUQ4OoQNTGHCVCVBOGN
DO80oinNPf1jRcXw64mW6vjx4Hrxlj//nbhFEzY70n+rWeYEWK8t5KA6YHCa
x43VMTr8TzlDduXnZRBiXtmrsQzgEZlKj3pQC2Sefg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Za9f9cbYMwU+4h55BM7Vlzh8a51k2m1vUmLhilvsi6H3jJbFAfEqakgQcV/s
g00trWUjc/P0TUkOz7Tuml8gcnB0tUp7H92AGZsXClBBFkGDon/HnARF8BTu
Wz5s6yAFkQDryVK5asaKbItyg5RAJ2raP/PRQb5kQEAu3gdsa1L+EitsRvZ5
peIXtsr+6wVahxMZGwjpavqaPEy43tG4neVEUEhmlvslOwv6DfZ8g6z4YSii
Na7W1RuPzBHbjWRSbnKgRXeRwKWPBsybHUxL+D9DTWPOekBPq+4eRr7KeZQC
Ek5CeVTGOqSuRmdak/7TK4UY3QeaxNhRUDsUDP3VrA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oKs59XGe4WurTlw/EYurGYtovVmPysiQZzziGmWjxPF4p/LiTvdzyH2N9TDa
HzRJKgs5REJGEfwqQdXcoilm0RjfzXvGGLJ5rfclhPXhDZ8P18nf3B/0poDN
CoqvpAJEHr6tNec1a10MwvS+avVEQaYHPZflPXX7NoxI9LNDelM+Jb7N59XS
DdPTxy/m5UZc3jdA1+h86OlaXcZRQ0JRE95Mud8PthHn8C+xmbtqizIpsn4J
nfLevMRQyyeQBR+VlkY1l2uuLf1dgrmY5EU48497QGaq4Lxg2uz5tY1MfjgJ
KqLIPl5CKAsBDM0CdP8AqKMFJs8AL8M2bmpT5eYtcA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
DeAKXJE2DxtyF7/aVeukg2OsfaL9SOqedJctWnNloc1EcYvJmOx4qNivoRj3
IE4aqPrglf1AeXEij4bllkHTvZZouk7wo451WZ/1b3jsYPPUhP9LFFeSbC7F
WnotO9cZzzyxl6DMB8k7uRB/8i4Bm5O4ix63tZT018Mj7BpnoaQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oFolaF17NZPovTbAbA0aWxrcSxoWkUIGRTQnw9j+EUW7SeoopN6iCjoO0Ebh
9AHpNgmA1W729y4HpXutHurhRm1RltLqVD2RxdF4eH5yCd8VVPfJSB9gslPl
CkNQGr7Mf0LzAkG1Ytz6hskXV1Zo8q9x466ACrtCQOvdz/jSZrImBtyyc718
xwqZJ8h2L3Rag906y1vgpyfoCFYHjJ6uxbFIHB7hckLTPzKM4v7i2w2VZOZ5
zF/5D7JD8xYatXP5JmNLuTEl5842H/tzeXCvRhBqzflNr92DjtXuwYQpXl9y
FDYt0qJzw8zLynnLBp5lQFyDV7QmkpTeg4kTlWg102DgT0czX2fLpJ2zYIBm
sPpp1N7qqL+bd/ymBhPmcSLlDs8YsMN5pdJc2HfZvJYY/F8C8RVMrKDD5B2U
4mJMSA/As6Tnpq0enh5uHLOvIeHe/nnEMDtY1j5O7CM38W5C/sjO2a2fs3ls
z4cl+KeQeNvjzRNbxCZkrcd0xl3oWbRF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cvJSnpJc3Sc3Y618uVT4KZKhfY+v2r4VzEYm87qbDaKcnhoPqAxSff1rwgsI
tAxXmDJNpvYsY1q2ujFIuTCnsLu1y1eMpfpOl40G7v+UqWWbx+vMeJ6HyW6c
BK0USE3o6VO4oD8z9mutD6vl+7mzGXMNOdGde1C7ZGGEvE0dV+U=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jgqU1KAlbcVCrR4/ct6v+D5ZRf2qzb8ROM5l43L2lbiVwmBjeKNEqXkPwHGE
M4x03Xn/JR1LuRlr2y10eEDIY8ce8TEhTWCsMEN05EKNy/L3/iROQaQ90kL9
KFZAD54NJ+y/r4aPuLh+nQHJ22nuYpyE8mMR+fnnUCqS8KnB8MA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 3344)
`pragma protect data_block
cW0uG05IEe5RHl4cuO23KjxrKOq7xmqrx+wUF/5EewIfryLmZMpDilgd4unI
PO6NmxxObFoi6FNyfzeCSN81L4pmPf1mKcQ80gveeBNNBoOzBjpRs+oJW8xh
SwQlHSGuUMtLO5LcVUMF5Cc/Pjm74NRk+rP9Q5vE2PhqcNtTN/yvktnfObx9
Npmj2fhwi7H/Hs2gAtB56s/v3tuJuhwY6lqVvnOXuQClmXW8zZxTubhKv/cX
7ZFp/Mwlg69dX+QXW/Eze93ozw94cqLkblAwulZQOq9oKZ0FZPuwibBFNQV1
pj1Eyt4SQWoQ5IEPMFPtLvTFwIgPgOa75fmxlquY+g6QWRXSoHc/I291DbLw
KGLeUQAJfaroC2zdGiu3CJxgZkLUTUnXtjkItChvFUOaxQ9TGvw++OJP0Gq0
sMJlafTZxQkEzJOY3qy1q400sgMweqiApfkrIcms8BeTdpsMLXjv1NCG8bmZ
1XRnVPn003/o8p7W4+E48PD65qNluaq7a1xT4ix8d8ZS9dkXqpPRN1Mlt5Ub
49E4Zv5oTfBq+W8fd4Zun8JCgz8/p/9TQBJVaSD58YB7ASx+cjh+ElfttaS3
p8HYG4hOw5436XA0gkwj9fZTxGw948xnWwffYXei5d7JVxkx7r5knijwPsZ0
E3wFddjvU6tgaGkjpLIDGS8HS8SiCyuzRqvigFURount6+cdRDaRKvu9Vj8d
Kw049jZi9NsEZCMIdvioSh1xaBlae+a75/uCDszdoJMs5l2aPVEfeiNhXLJW
WO0uIZ0SHYlZf9TNpaZr6yQflgHfksRuROfxGLelXLVW+dyPqOgPyZp0CQXA
iRke8bRMqhjqR9jourdTDJMYl8ITzgidV8fiihZ8loYDNr79Cx5hQQ0f6Gp1
Rt4ewqSEIOAQIWGy9aYBRfyl4uTzFRp4hKf7STBfT54/k+GYC+khMH8XxufK
XLXcBwazl64F8cGOkvyitZ1hOI4s7iFozhfMOb3fSKFDuLG1VCavJwsTr+dK
VWfcFzeMRYca/rRcb42SphReaTny3crMyrZ66Vd+m8YghmfxanrUD9NU+1Rg
L2wJrapkMeC8aIWsr5OUMZfov8PXuQfFso5trM+IOrFcgoA6NXKHizEwZ7Ys
r0gtdJIBCncEBr4V7HPMQGNaqHb+juf2rVoOY6JYq6isjJ8e3yT6blFTBPJN
4dn3K7uzQzyfEPJHD1S7h3AxCv6XyZWbLNgTHqZTMysrQqK9dmicTdnmUqH+
z0LkN06heXnZaCBBQA4BxongiRRfcTrj0D96XVwvKTrL1shSBZ/v+0baZwiY
gurDM2Aw1Xydkw3Ht4e0/voFLv+nOYQjy155sUyJQMiRmJ14j0zSONEjPp9t
vuxp+wXGbGJzA553JokJT61iKhGTQZe8JXyJL6Gb57OZVC2H7W1CHMOH915v
tjzDQX0A1188kJ1dVbECAK6WxtS8qQW8wf4gbADY7S88eDHqtI8l9dOb0499
xgiXQPrwb+M1nZYwH8yGdxcCC+ttj045nf8SM2o4qk4gVgQGlfm8/S2Eo/gS
n6rkGWZ7IEKZib7F7F/AVvCuJ/8CDVP2oIzI96ngr8GOOPMVHjawCJxbj+h4
cbZQ2imToPIKMp+yA8/BcK2hIG+gEBBjTy6qgcm8u1BPO76uInaY4/5uS4qp
HveW/vvY1fvu1plgn3LfIZl0oTs3rdDEg7d9EkLrLI5lGlVV8vgKQboQMSH3
ED3ZQHTSOLV+sgDRzTm/DeNQQ0oo9xwcINE9XlU7mk+RZwquAi5vNT4IqZaz
EhMzSGbxT5LyOi6P4dvNQ4dWpVgwKjKh4gKZIf5Wo2Zf1YT2QAtBKcKnp/gp
13MlW6GqbprVLokUyS/5nufl76naLO2I2MUTZba84HEZRqWjQjhoybJWo1to
tMl6zQDtQyq4TOjXGXPsVVg0ATHeE0bYfgOBAIQ7NmPL5Hv+Sjo0YWHqxd+D
pRRvfC4SvK0db26H0wbLxw0ErcuG/c58vQVTNMG3keqMGsxFQCUf0+BqDqWQ
xqXRyw8pvMtMhMDUdAa2yF0ypHrS59qVZGK32AC4yAPAUGzpagWDFU7ngVWo
6/QXE4Y8aE6PG3eWBWYgQkBphgtwvTQSR/jKYHEhAShTf2sqIvYVrfRWGV/i
wqTWqbNP6+Mlp85wfBYLaXDH3sK/n/6Ya5yopONf8Ygb3vRWqnwMYDj/pCYk
1AY+2rXOEcySx0n29zuemVMleIrifn1oiFemqXGIGwydjiDOaHmWmVbgZEmP
9hOSB8VanXUdfVJKcTYFzwi4IgEgeMndZhSmiFjNLpdy96Uwwy9cmnW9UrM0
jX2Pbxq+KiIIP/nSA1DnwxVfEzfJHYhJlp5VLAlSH8V+U60rwm7cFoAT1WM3
MwEqx8sd9dcT1epoNLi7tr2W4W/o+FTVMpwnx5fn4FhfziP1YlZg8vjoEIbH
p9/Irwwf42kruXdTLy9g0ozduIt5b12dmkLePJ4c6gqhCYIwn9ELw1lOyrLv
kdgkHProFgl7wse19XwM1mA89XLCaoVt6hDvHPtjEZ1/4ZBGx9ov0OHG88zC
hrWolHynZGi5yoDjdfPL9SSzNp1XbsOYOPjThp2CynDo/cv6WU7HuS4htgLs
giRCWmmK7blUeCe6OWBeaBEFZybF3xKwS+91z3Jfyr/22pi5rrocLTDiyt2u
1Kh+zl1lAaeKc+IvCzqgJAqvwJNdUjbpzsmYdwtQX30e04hn89qlUHat5v2A
uqO5NF+0AAVVsRDF5qsWiEt67p1KfmMGYGJDGVxoC+F4n5Z6lhwzP5Ngbk83
RtH08Ve7e3V/zLFFanVq3QPsCQUUfIQ44rxr9sZIQWdLfizUbcpqjcFKnm6T
Y4k92hH51yJfWZ2LXGw9jmjqQMgPurQSfkEuPewVY98LG3RYYiQvV8MryPaP
E+VPNionsedxuyzOIfbiX17sgWxTt00RLlD5l8lAbrzggNgRH89re3ppKHE2
UGqOIgrdpv+HqboHbnSNvneAAPzkOpmkWqSAWfS1K1pQsPNW3wAICmMbpc+t
rO1wwyicwhiqnnrB7RLTWEuC1ABGGDzdUYx/GL4IQ6cuUfoiyPvTn8+1k8TV
EF7TvjGaGJJplxNbAxtYSl1hWJ4xqNCrqlmLthh11btAYom0vPTmQNksLCmR
ALXx/i1OizU0kiMnRXPQmj1wThdpGuhSO1xbNU9aysF7BtaMnl7Wwsv+ow55
AMewc/M64sHeBxM1IgkJxJNDp9QvhA/uk7ogA9dBOEH4l2Bq3jA3wPa5o6d9
lKk+tJbG7OBDYV6Jiy+XPFRcQlEnUNUfYLdB0WBGDYZsHoTHEN5WGUgRiDij
SmEYHWXl5bFd3O1uIn3GholRLZ5KH5I+aRctrRS20TfyvGaZ8MWzgVvAkSNm
KVjZqvhVSxMNUinnnbEK/W7HMjoZScA76mcTPv6iQX52JcpuCnhNeVbOG2Q9
Jb4h7Ypkmml6KYdOUoohBGONjHeCf2fuc07Te6qY65HfOtXovlzi1vXFBquy
DGQP6o2K5AiAktDDWc4u7L5AnquFpRKfWB29Y3ku9yChRIv5u1UCMAnVpf6o
d5taxEmW23559B1aXYkqWfnaiT2ECTeTs0gHDy3Wyq8kJ9sWeVNoTPwID/VA
J8hmcY7eIMGtXv9F+9mG9yQLIyWQZOSdlliaFdX4I+IijS3lLLsxgKWV5EIV
WowqQe94UXGBClW6BzGv0btp4zTrhSEUPoh9e+VRAovfHxr1q6FeH3FvLix7
Rj45IUvm/nSxux/kuwYt/bHDBCoU6YzhfSd14rSD1u3D6SXEOo28UYEpGB86
iEKbIcPk+K7C+uCfgceSxgMQMNEGnaspDQzFMjYe4Ag06MtMu65dlzMfnSLJ
Dvt2BnVac1HBdZ6yLiB2iTphTShL9jiOCnVXWAod89bU47sD+nvnYjg3n1h0
XMTBXzbheRHYwMsazfTfqfbw1ji/jA/1Yq7ens/tbHFqL4QocE7xjRHAJs47
Ce7CPZ7r86tkTLUrLnI7xia62sGZXLz+vxPeIJpS2+QEZ4iYv9CDXbosQ/i+
xdyLgQNs/9DDVtEr/z1NNoSCvXAo/IVUFPjcQKQlVytK4natSUSXX6Vpt3T7
H9xW6Lv5Tgu5HmkI++f6u+Z2eohLP9cbAkK6T8U4s8rX2WjGB9/jEvjdkTiW
Ca+gsrDEOG27IekfkR4pxFGPDBkXG/FlMs6S2CkDlID2+G5B6hO05fbij+Fd
aBEbobdoVn+6ROoGsePO2graW23Aa9LVeaE7yY6JScvr9Sxzlyh0m5OqScTR
mk53HHWqcP6jgtd9aGcLgWC0EkTQ8N2sWmAj/9AswyHeNMsYx89n7BSYWpNR
peC7ivYXWUFs7adeGwrAm2iuE60C6I1x7ATWHrZOg+6O953ZxsLcGjGSg2I3
AjGFHmnehs8yZJ26SL4=

`pragma protect end_protected
