// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ej+bb73hkyHMMWBArFKZbuIZjo9RZ4UYJvZCS+S0W+oyqpHQvwrTxA4fo/AuyUpEPMFevCkkbLDE
+xLheyUNigtmiyPZQDSpmynBoEiTXjcJ5RF3L4o+4pSSdhX21QIoQ2MZCn2zquxfGhV8yZ4LaYvK
3WAE/9YruIQ+Su7v50dMoZklk91H3j0JEBawY2kaivniLOSyn49AyF/GrKsAGzmFlZkwPmWK88vb
if06krr04d4MEbJG5ycrRQkzaR2TybzinoKsUtWlVfzURnsxw5K+wM4wNT5fB1r52ub6K3oyZttj
rxaAEU90xrPCS5Afdz9qhklf69F2RD9DjSCNvg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6688)
RChzUsUVDH4R3cCy2aDqRnCPywvS+FCAh4fTQd+UjwpgesZQvYkTuKS4AQ4Epk25iKE14ElxlYr0
bkaYRz/0ZJtfqNpy1pv2u4586Fh5BvraQXyh0CaVet3Ew+/3RBziNmjPrP0Y5rnO6xwaqGoPmLME
fXVTTu5s3Y9q1UTpmmXFErsy/aDz2TuiiyvyMfKX2Fx0Adf5kUFq5aciNlVjcnx/5l+/mzFqmBov
Fu7j7BLqhUcjGBM7d5b3GXg/9z8BPV6rji/a2ZIFLZyGzrOEvMa7ypPVn+b5KiSGNNFPDmAwbORF
Mkyo/F/kXyjcOA4UYWDuBVvT2Tiup9PsLGqA35k0QtSEqoKfldOC0i8oOEm/wcnJkRDoW1wqBnju
0n93oJ6t6JPg05ysKaq+m1M2Kc+eJ5uWFsE/xjs5e+D3mIhpCZX326xMvILEQqkSaVSQSgttyCfn
FbLY8ohO9gYNXtK5taRNSnS3iCvcIE0fWkuieQNRMHZu0D78d+GV86BDOweUkpW8AYXG62uvlaNH
hpmAYsj6HOJ5k0VyqYtBBuKRuTLbptdj8OZvw+EVnDJ4WEOZhgj2YBHurS1tSGpzCHH+JwvMd00l
9/OpetOQOvWYPdGKu7iMX9G33Q6+dNh9KRrDkD884+nevDEx7DnV4XjqLHeuPus9+Vuk1FMqmFFy
ASyJYnd2RbMKbldpp2op0KdllxwTnG9w6+TWbymDiA5olKMKtgW1Rx+SAk7n5fC8lN/Jc9MpmJnf
rkr7anv3LKkRcYap4Sr95sjg3Ot9vrELV/hLfZ40WFLgpO1uj2Ig3AIk02N29cQSI8qun/iSLLi0
ujV9rzcDYEMm8DU6HL/Y5rIKzg8NPcgbmD5CxzFvQkH9y49Wnogmsv0uCQ88U1AcBFxsTrPn/efA
tnDu1ceGtA5NTELQwDJMJKKNa2XbbihWBt1WsRa8zp558RN/JxM4xB6JZ5zMibOhPmgvxDGqg9w3
XVecXdzdnBdGcdMohXLivGFJL1imBn8abhjkeFyYrBPMUyxLHoJrfColJ8Me/+BG0cIx8JmdPnJT
zF5yj2dhX3CcuK+Ymy7uaeODTfR7MaqLt5+yPcx3Jjvps5CbgowaNbwq9L1GA/xta6b8lbNrESNl
Y7rgRyxO+JSwMEkZ+vipDVi3Fn0Ar+30VEfk0Wgu6zyjgh9EGn5C53r7QRbtzIgAvjxRhENeWpEt
7eQdLyUxVhuue/wwZIjVT4+zaDk6LmIe9e/6mXHkvXymV0WInAyHH1DVRGLHWA/LfHBDdT4RNAQB
0rVKY+XGKFgxYrAIEBMyv3qoaYFq30jVoBiFJdMiP0L4xonWBSk7+GrpOmgbA4I87r5qVlHQAWHU
v85se/IMK8NZReoeYqobnH5YCTT82Z3+4qZkNIkwLw9obpodvs5EEfCB9R7biLc09xWZnhIYSb7V
oOaak8TCjSNZVGiN3V+05Fq1WG575JKdw6jTfjR4P51ZX6cN/3gq/+Tzvzzch93BzQWxeXpRvj8z
EMLggZQQ9Rx8fPZ4sq1h+L+YejvcF5R/8X2b80LVbNjOjRj8sZvgncRrdPh78EhiQ0P3NkGoSlKg
8fIus1rgrFeRae6BOslnfU9ObARZbFYXY9QZHH6zGfpCqxIu2iyfFC8/z+nONbFt0G5bx3jZ10Jk
poxvnKeBm8ofrYEz1o9rkJOuc6Bsj8qvA2h17E7CwSRHAeYCkLuuHOW7JWCQOgWehLx3AXEfeRRB
jYbo6f7m3T0/rc1RsHIiMz9EOJqHr8rFybo/5Mncjcmc8BloVswaetEZ891qa927qeNYPXawtwsd
zFpsUvdkDe9mCAswZRQQMkuZtMQCkDxccqqDlYC/vzxz0ZdpmTRlutLkPn9jt9RBDbX29xPj//A7
Y8/Fq0ph6rYFRsAHyTXxxvr7Po+gS6YI/kU/8fSYhYYBd9VBsKhfjCGQeBtahZPIh0FLs9lbqva9
2gc6GMYLaejmZl1BKX69Lmgvj4D0tQto3wGwawWFsaefJCAer/MFL+lGDEv7RKvfaic44eOqzIg0
Nrl6vuxzWECIcCMIJivKhGgxnlJf1E/sln0LhH1DCMoJ2zqSP9mhu0gsi3c1qyHOuz6/zLNoIq8G
1m8qsG+grU6/B5KtGJENgBZcDFhOcCl6odyI0fjmkx/uE9Bx0OprzNtiC/g+znJCZ1hMZiVR3VAT
m+zwSPwEC8UyEjPyFfdI+6e4JHch4ckKHPJBBjMqgopQn9Fg26dVVQa1huzTlRpEq9lAChDt4syY
46pNP6aPctlQ9gcAYG9g1mlvzWof0tws5hm+TwFabWSEv62sQKiFF+wfqONho85JXrteXE4o1LSk
0+y2dpcK766mjw3t4U+CK4/0M8Qj03dtW23QJoe7mpecWsX2+L1vfsdxsXCD9HZI3ixMw8HwZZt5
bF7H/tqbA5z+/pMqhmXfR9U3MVoxc736HixhuUsZXcBzaN3VlkrTnazH07zHLDYUpth9zQv1zhXS
dTDGZ7L2OECgM4eVaLPX2pD5MlGCa5C+NMBf4D+GCr9vOvb+TDv2kQSqoFVV9FIek5Wl3cKT/ne+
PzRxGav1d2RMuHUQd556NwsGjjde/SsOITDADu2Lc4LJ2xHyjtZYRbih8zTbregCpU2YJR3vhSob
YCOSUp4kt28OUxbk/GNp8doeLb11j4a2U7o01E2YGO7i3Mf9G5kbThAtXEb/3isUwrkQvFs4VlS3
Hm4QlF7DaBX9r7dfr5J7hn7O+JoqONV1oBtdG8+ha+j8xGKBkx81303FVRIT1TOtNu3+qtZt1wdH
oRDbzAstcbi62xCxpWD8zeLPQpLuIz+lMcGnkuSNqVC7vu0RAztAxKNDziTMnWx3JZCb3UNThu8l
g0zegLmNx8IraLyxfZB8ytV4bLX0Q4bYV33Q/+OnfY64pkpHtYYRVS2bnPcQFvWgbg+lxiYgWXpD
ZGZfLQqYbtItZwuUF1eJxAEdwxyxP3uKzyCVmTnrPRrc4hT8AF9LewFO6e1dBaYjr/Dfgo114y7o
1yiV8RWxOHcjtzzRfDlep/KCxEeXrSzovkLpuot8PrBD9hZM8kTtSOL+4QS3SDKpCBJAXcB1BtbI
22J/VcwQ2f00jD8EreFtq/ciYSvXgWDM+9KDGA65Vk+u3NZFpvoWlRB0iOVM56WJBDNyIbJpWiuM
5cyW+x4fjFg8MWa3Ot9PTq1ARZftIgsqav9HoPCcRhGWgTr7WnKJhD2OV3wxo+1H2oLLCbku3grW
+kr8g8FS+JGM0Fe6rTaPz11vW0aoQFyM/589JxtnN4PjzqZQMwDJWhjGBHPyFMX7jA5T0EM0a2QN
Lc7j40BbH9igHbkiuhKypW+uX1zNC+EncPRFemGlwkPbGMsUgMKLFUFYFx3+Zey5m0IOfwPosvps
AqLpEdToz4y2+zdtFWxFxkZrEZ7F9r/CiLdkC4kkd4C1MEOSooN9ZHtyAnPXdh5JLZYBDreYZEMd
Zb53pDHCDJQuZdb2vWGWJV/Legn5SSiMpopq6gwsquJcw3auSGTPyxZqcr3S2MlIe9CF0KK4BxWD
kN4CvtdRGSKdl9/zrdVfR6RXdNJ/U6MTX6se5VyG6ySrlYoWIK62gSU+rWdMmnLGL6T4FxV4a0eu
o08YhU2JX92Kf0SLiavuDWU6ePXd9N3gY/MkBEcHvXFii0GAx8cQxbugpjv/yiw1o/JJfWXkjmAF
HZ0cxLj32w/h7v8ltDBRC1h2tWCCjuvLcuvVXfmlFO0J0b7U+q7h0jZQpXA6Y5RDCduE8bBK0RiN
5dZ9lSpOfzCDRolIHydO3tzyoqMdym5SHoaBV5y2rVZFdv9k6fy3okA3ciOT6XPp7gLCgH6p2rBy
51wCP8pkarQ5AtHTPMHYcSlqOr7cCZan+qvoIJEBqvBspbNHQ8lShDWgVvaSfzuoGXiKra2q+1et
vrNw9sGkE1tyWqsl2v8FtE753SSM8dOg5ae8UxlRKeidhtH71WuBgkcOfJzjmjIeFFU2q1BG61eF
GTitsfb4Ptd2jfDFyPdNILfM7JrGtZgP87a4e0TIBXjMwllp1mDw98Fj3w/yU1NCDY2mdXzNKxZ7
nOi5yVnTrB2D6j7qcMQmvCVWoR33eHTirCUIgfHjZWx3r/4DHO/FwoyCJ5pZljYWqs7aI9/oNyvS
6A0iEFvqR9ccI8lsc3Hp3dU1BRhPl+G2U79oHdLPStVBRMKvkenzLbAU9F1YwOOjbKMQLuGq/3X1
IWC9OM/1ld0a76vmlioGn7JfEozzqiXB11mx38YVNDpAGj/k2Bks1H2JmjyJnICtVrr/aOwcVSTU
d7LqaIXiXiFl/GLsbz1xKIzjMhqUnuarxgMID4AJwqvpd7BeftDnooNw2LeOEAgKitZSZThefhOS
C2pjRcGC9AF6luVUdkzQfQpgHfEDKspr6WI6UfyC8wLIrYqk4WonkD/48J/OLbL3M2FDU7HLj+a2
d95Vsz5nr5JmMnhZl94aL58q+4PZXqYr1tHuq4U8T4UChSb7E1lCuNmSITdN9DC7dBqrzMeY6lCg
9sQYicPepWtD9vnpG9Un44c85bv1Vbmy12KSBZP46FxA/WilC3Qr25jp1PEtxL1BSBF+Z3qFRVgo
Y9OaFyM8NZ3k8NDAfl8/Wtv97SqQjH6crzz1AxS8r6/lJ64bVWzmLLnj+yGARicdoVurEawIeulh
syF3KE5u6et+bEFFU5Q9i1f8Bypo8vn6G91gpFOqVqjo1xufkBsR7XplbRC1huCV2bMcp39zhGNA
yMJIHvEA17+ilS6vvpp5+krYmh7pT6xyOLJrRuOqql1IxMyYl98x6r7kpVEHCVijkphnLBSShVYo
/ocB1IcyjW8paGGabFoiwTxjFSTfClmkzw9ZHf/K6qadPoVpMpbk/xiPCecBmswekdqBoO6+locl
o3/IerKiMUld+TV8VPlkLbKU0+XVnUpNJbfx1z0593rvxw+ID+iJJspAlxqldzy42NBX3aMYpWDq
u57+gk/S23jHY7CFlrB/r7iIpcgsO4p+tgAn4nZp0cs/5PPfDrbF+9t1X+PivFZtWbVOEMhySNiy
kxHkWFEYnP6LuJenavcw1uXthe2tqKQDmnE9WFIQTogQuOdx2Jneza0kfN69Tgw3K55LhnZVNgMt
LI/iqc2oe8kkA2YyWz9dBx1oWXnZ1RibxHQzN99m1EriFXfzsAEWcjI7BGeKm71FLYdeIvoSu7+q
rT09G58Bp44/4IN6RQMO/uWcUONYePVF+iIU1zFP/lTRE9ie4iJ5p8JKdzNfjAnBTGr5qkVZ+0M/
ZkDdfzK93w6EI8EkF1jYZkBhMS5fcdYH0IlJZeZyvQCrx/RzZZmX239RHulnpGcAj1vo9EfRwoNg
TwjxX5jC6gf9QBu5nmfJs8zwFSU7hk2qTkHe8uGBkkg2lXIx1bS9qAE1zF0MzQwWuoo1moh18Odh
QWIbCtsSkaUrpYdahaLDLns6m37WkVHS5tCVMsxnUaEJMX6kOFFv8vQCXqVCNEtCuJkV+3eRuw80
NoI/zAqBUhRyt4gWBNLftIHWv+LD9jdxargUbXDwZ6JsFTLWhXZpe/uMMSvqhCVKRI3z/efpym3v
IttEAHeJ3nSpzGdjRMh0H8GnQsw+lzf1KIu4KROsylbTbyUKQ66GA4OqGMVC/HQApayhCuYa56PF
Tj7oRLGSls+esJi6djduaVfOk8aZ72oMdD16KvKxo2uiepyX2QXeegcT1vHVtnxpB/3bG5w/ky6m
FuoNSCX9aaQPMELcQ1s1kPB3szGTiuE6Jon0ZVotF7wnDFpQBNbDOuK6yMZ3C1WJThDYwJ+dKNWt
t6A9UK64U2KiryOCNRhsseiWGWeGiDMgtCGIiIWvdJi4tzCPursdtzPZ84JLB4urry8+M5JeS037
5OcoeKM0wMk0rwI8udJTqm99yNfoOL93+5/fx2qL1kuqfG5kAEq1Zl59zq+cSdc5kisoHhm9sD6r
+PjkX7lmpGDLvBo+5WMbOgbQdgBbXWVwglF0vTdoqT4zr68He/qxAaSPfN/mhNBaNYEDEK9/K76k
fQpyt+9ukceDBs0wEw/atTPMvYSQUeIYx3mK5SHVDA3lUdr/nA/WVZwV8lsRqMlGgwXbpW9JwbCq
7jfsRr8h4OBhTfEvNdwjM6MICYjBNjqURcaqXsiYT2HQoA8FKWb1yZBpa10VW9FzFF/pm0KfUH0+
pSTHWmdRAULjqEc5dHX8ILvMPvuY+9GITHXxWRnNSYpQD6kVTlTMwW4KjERO0qAgLX7ago/a5cGr
i9Bpaoo3brAD5+r4RuNZgQExoCSfR3NRXufCyjUHXt3nChaAqee+DWrhjLyyzC6xqJQqczs15sSE
gBi4AdVWFYk8QvcxuufmaekkfvggTcmiWmLhkqI2HOoeZtoTlIAKAhiBxT1JEefveR6+Hcnlkx23
bQ4kL2ZD/lSep4qh2XT+bSne/Aa9XPEyOmMUtg9brBHogAZIsmb2rMFRi48RTEEftx7Gg9XAqjjr
9otiwNSySHntgie6fOWO0DL84gO2YaDe36mEqROPEsXN09wz/eGRoGnGSTiMX8hzD5tUcqdTOsg1
HidsDUiSrg0TfqCArpwHciAaRoOfJOPrMOlzT8ATf8lrGSmtQiBLztXVZ+pVYA6fAy10IVnGIaeS
bvykBVH3Rsn/yKL7SPzeEoWjyHXmZeDg8QseVwTpoWgok94JbG71PrtUql0EX8qx2uP2i01UlzCu
Icb4MVtEbhEuOeUfPW21FlfWlo3oWTy4Wpu8nf9z9bfmHyKI+9k98AD6M6wj/OsWfQIXyAaStpwo
TpfGZZj+LWWaZxK0KwabWFzXJDUt8sfago5clPuOZ4yvBm2HtPFRKDcqQPG0ut1qvCBfoba3TxkE
KqVB2q2BhdTIsN/hqoP1epoJkniGjFSDV2vi/5IXsQ+Uo7dXXwb6YLa+7feS6P0PCUtQe3REbEQs
CIL9S/AX8zFIWFBDg49wPcYk6YwdHbMzmK0gca56osBFexlav19VeqlJLfYnkCJTkecQbAI9bxRX
ey//7UXoJE/kPP+Dko/aHAbwFyLoQWJ5lQhG2A5mOHUEN9pWJ/4HtOn0Uc6XzFAR46zfvoLxDna+
q3n6hz9o2WiR8dYDa/08lp0idIdVUa8qN457PGM1LmozZX2PE9AagGaO6tdRS/7SdTtIQI2tWXhc
1njKCWYJnqbZ3FguWtUTdR3GRNMHYdDw7OEWVIViiWj3gt0p8dLOguhWvkSmTNzWSzeGqlwpqIiK
h4qPykIN4TzRuduAzw3PVfwjHNfHTL2BIQbDQLIj0okecSHh6lyOg7cdmN8WigaWMIXzssCxCWoF
P6UNO8c+NIQrVLq5RmPE2zQVyt72DCe+lq6G32SuH9qsdU7lxr3/kuvNxAeszx9FYH0SXCSou4eW
zS6PKqAYBD9G+8lLm3xTSXnVgbM9OR5R45BDAE6h065iaySXkxTSAY7dqqwCxRecz+VjTkgGK4Sy
N6QPJlZ2wm0IFi+oR0gHthdOyPSQeyHTEa20frnOJbFPft/YUTXy6I1L1yFaQd/J2nutOPJU5R5h
L5zJRADbzJWWGLPDUDJzRj+lCGiBtrB/iQfEZl0FNj3WbT6BgWvWe8sOl1nPrrEOFbhsE54+Ri91
XzlIWwlc0yotrCFDH6YwleTG98+mAoy6Ii3Vv/9SAIFciaFL5vfysKAGJuXBcB/N0lHSOFoi5nuA
aODiGw2RmygzDMOD+aNXGBR0Ur287N9Cf/sJuepTr9vWix1zU6swl7+dGJZxzB6RhbciWpqyb4LE
zM0ic5CUw6B9dC4x6CnfIDOiQqRNnazF4qBCdlxNN+zmnrNe7DhgihillwL0Na/G3I6BOt+euQMc
Q8794gBDI49hj4KIAMgoTD5/ufM1obWKnI+Ncq37eXM7Ns9vELy/8upEslDupob0Pf/OuuBokVw6
HRo/p9V8IAMP8xVQfT2PwbMemGJNiRng6z8/vTIPbkRu+KzLYSytwS64FZwcmKu6pyAj6ecsWSdY
YKNFMKgdVZB9MUn2W9axH04f6aS3bVWzJxdrZtIOFPrQ34sQOMeSM7+QaBFEFKYMO9Wgeb9G9D09
LdMyaxTkO0uENBi6gLZkmC7LdZJmjodYcdw57kj6kq44kdTJ74uBLJfRkEABlUjc/UuTIYH5lnKt
elxBoW+nY+adsbXOXcESSL6L8uKt+uwV7RtM7kSJooZZYgrkiq7euV4MpeBAmwOCLpCJ35CsiM7q
wQ3hj1cPwv2TYYCRSUKAq3FtskAHYSYIjOdJdmQcB8jvN6g2vFjsqrzbmj1mZPzCyJl4BdylD6Dw
mX66zSr8h7Y2tOiaIRqYVkIgxah4D29ABHh84/SJJAwDTUxMxTXmBwsmNh/Xnn+zb3LOiVBEcea3
kx6wHwGd5wRNqsLV3ezp+hBqxTKmPRF3fAszxepEfFuWq8HMrfj4NE6Veu/x+X2+a6ftImnn2+OP
3C0fWa4r2bc+75sWLZt8r0vpfNGdtFTe7MuFCWiVbf0Hnki8y5OVBBgM9yjzjBN67/d4Fi/EiKEh
HKawJFDRT5gYGyUj6f9xqFsqM7t5UhcSiZDiNPHkc5TrZ9tKTwJAA8CHWH+gntPV2FI7eSZqS5P+
R5zRMSfedl7UDSFIvkSmmSmOpIgPwcWzVG8KjyufEQHfJW25KIn4gUpK8unBw7tpK36BaP9Q6pp2
D+JsA6DFxIf8gRX3cOXJs02Vp7DH3zcB8SB8q2kM1UlzsrJVcb82BwpYcpgseMc0LWnj0rki+Uks
lWIaBEO02TDj1KtZgsfp7U51vn8dVQn5uE5OkRnutUiKR20AGcVqisxGiMSjYXUPjeCse5QE1yf4
Qr9CMkLwXzYrIiqr/YawInHYoQ==
`pragma protect end_protected
