`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
KMIPh6eGRfFaepdlslCv4o/OWnFZscB1qrux7IPWasArkHfkye5oSNxOvGEtgR8q
AVi6VEeif6P90md8qj9VU5YBOIsSTOu+0ELMxYDMIFevSVIBXp8kAXXw7hK0yg/c
oSFGBxfmIjIt8FSR1HX/cArIZRUp5TR0zrEiracwc4E=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8576), data_block
ET8XYxYnRvZa3lUeJGcx4tEtI75zyJgQ6l+aAQjm1veiNWIh40qfh+NG+ICeCYhW
S0GZky9E8i4FJuMqDaq3pE80oFdS5VGbeOL37++v3VBotlYL/8roY26aVXHxSw+Q
vAOw1QdnbXxXui+JRD2A+WbNFGGvlitSToco8h3RPVg4pOHslUF5BGbWiHtBy0qr
Fd02KPBcQDL8xxfSY2oiDBwi6kHQsPx4q7W829T0k1MvmP8BHVgvAFY5yurW5EU0
gUGtxxKDcwh1Xu2mAMTFMbtZ1UZe+OR5Hr/6/7fU0t8Jqgx0cw99yXvLCRZtvJMo
oY6aVi0Z2GKRHhL66LOiaQzp9b/Bq2uEz8ACCVX0d49FitT8K8Ct9z0rQekaobnu
MIPBNVDpnSL7JHa7LrjsCLmJ1hm0/MQ61KhcdR4lsZpk4ux2TOuDx/00hG10uDTc
DE6Kp1L/VMvjP6IuDv1jzfv6Fqo5uLJ9ySlkyp/pyVhfX+gb1hsR6/IWZXWWUe5N
H7Vb1TYnAZ3QFSP6GTR/PHKu4mZtlJ3jA9Pw01vUh09emRh7B2VpWdkBnrXv7NDI
tPB67kuQEddgPTtbjeAGKssapjhSnb3GrbFt7tNKY/c+v2ke22EZkk2LjQyg+2J7
RIVueFtapzi5ONxw7Fxu0R1232XayN7xogG6jl05at2KyabzYnuBrg91ycBdH8kD
lUT6gQcJjULveL+wDDRLmVBs4LmmhfzdvOJcHM+ziigQgbNpSiv0BRkPs0f8U8P2
OvuA7pAv9By1C2gpjBhV+v0x+ihEUXTJx8Jepg7aD09S7/+FeS7kmwirzGXX0k3u
3arsgyjpiSL61A0I8Toy2vkXOQiNO1Qp5wbOgyLhOat0FniDB+quMEEOj+86vDF1
R9PVokCmw0EAle6RIp4vuAWcQ4gQHEMihYsSGAqj4C2gMmKpaMLMvd/HiChKfBiH
NafYLOgtwXdznVLI3Od8CTRjQPV3d8QwAvpUFlsZkhGJqHK2w832y1HNeLYxKcML
UuLCA90RKQgpZS+bEeot8r1gBrotRo9naUHOa+lDZmVnWnae9nEZwberVVMFDqHu
4nbzauisI0yf9prB7C4dNIkyW6JbrpHy1SxQp7hTQSKMZ00YV6ChipXdVEvCtTag
83+dRxQWz5rwQZ9aClK0WgCM8SY1p0Jqq46FAWsR0XnaP0XyZv+LkzG+/vhwXfJU
D2zrNzhSKsb2fIQ8OpvTzFsgzGUQil2rboCDVVITbGUpkRYefFjoXzIMhX0K51xT
hHc8iAfOUYyMTP309yFDayytKQtD0N1uu+o0uOhL+QMKdfz7xGW0fyCQxezK2Bsm
uwit5RFkZ/ErrfWTBON4Z1vnYjPDQ8/9S9/pw6aLCXfcqMl0Ty++1in7WG0l6g3R
1Ke+f8BUIOV0kW57Hz64IAMK0LgOhmxyRISQxnB4MBkU2K7yv4vJpCuazdX38CDj
Q6ecTkdS6Kv8tWlLb9VDazZUfJYgPOoqB3MkKwVSQBUN7S/stlPdzz+pwakeT9xN
5Z36SuPjOGEhcrW3nMR7OdwfkNpKs+FEL8CEx4Oj0s7Nt49HftzrW/s4RG29o4XD
Tr9jcl5nCBvcirBX5TLg7v6d9aaPp0RVWZokoDD322CTEsoAQk3kK8sBCrXB/VDt
UzVK6/JKmjdAYcQHzZjft2RF7Kohw2e3ozqR5pA9kzi8462cJ7W43JK51VkBMsol
/15dlSk+JTQ5+RXUYPJHi9CklMOxCkTBFllpprwXWKTQ/orwWptVJZAnoyzxo9Lq
n+smkPA2r9aWR1mv0qh7P1IiHSmARm++lXI8P1q4It5F3O1jyyCW/OPKmxPiNp3Y
qmhZiDuq7ujNpWBR6DLG1qVz/URRX7vaUvkSSurvJqkG/o7CPWc4U18Na8vyE4HS
B7yNuWHTNGdVapRT52tXEJmzEu2CsLu4EY+b1SdWDSYvS3T0nXPhGQjnSf//5Ofc
NU3U4brLqEMbvCrza0HT6iGJtwPwr4Mc751LxOLeEjP9perRpm8xba0VrgvRBRKS
OWWaKtNrcu9CO2GAXMRd5YiRrLf25I3pHsj+3D8PTOTsidEgZk6WteGGavcEt0wI
6RI/IWrAgpZq/rWw8HtDlk5Jx3KQeR0LAcq1SfMHSsebRktE9GL+CJz0d8oC2i7o
sBzMycbI4w7K5ZDSp6/9giHKso4s0QXXgIfN651o0xRJSEVeMAF3gvQ/veLDMe8a
j7AHZ6pq11P3zKPTU/rDSiZW+lftBEVhEtb4QkV4DQg2Yae9kPzeTl41kDlrs0+f
N9Nvph5NoYbzBcfJ472Ote+UY3x0MNIiFK/AA/hQnZ3Dw31iFj0+lbI8eBhe01Ob
TjcnwqEMftbIPstNnMVEoXg2idXEvHjyKsbDbm1mrMrxQfFfvzs5PpXTS4zaYEvq
VYoZek7cgkEfP5GIEW5bJ/O36V5P4MqVu+2VAmWcvZkmswzzbQA+1D/IYzzXGGd3
8Xs1jkRhSObXL7TfJx4j58yFWTPT53TbRBD2Sxc+hRxkZtgkMnpoJFoLVRmVerac
68OGrE/ttFH/vw6qqYFN1u+e6Ge2GOffCwdU4VGQu0Oyy6S5nfw71WuDgr0UE7WP
ZlF5fjk+KnBn5fdmjHz3KVY46CDM4sYC7vNXpTalVmex5o34iCdNvbrLkM6O1Cq4
vkqfKvDEzUeCUr77dHVS2wP4JcAz6pEtJGR0YMOIKfjyjVbrDyvnH1Qy70iSD0s1
w5czc9KChmIOWV5x6KNubtpi1rfjEGw80hD0B4YbHD+BDH3VV9vyMtjE+IVUmrFB
WSWh4yD2JtX5J7KTKd9L0bcv3Wq8tkJsoGbckOOQ3BeuD9sWhpk5bF0MD7r3xX5j
IeVp537ivQK5WAi3azcMveUFw+BRqi3TyBnxrDBeKEsJWnRSBFMTJ36iV6WvNHiJ
zesaLvw1rHspkivD3CdQhHiUWM78QlWONLqHgwv/WbWqNqXWQQKdJEVhsc20PtEV
Argh+0AmNw3AX2RwPzo5llVL42CpLUt3HvAOx33V3xWILApvOiVzaMEYcqVuRf0y
RSQ6jR/fQaeqDbVmPCL6EjPNnlr7Hx0H9wFmIzO2nPIQPxoRvUkIaGTo3sN86AxR
89GhQ3m10tfcKlUVSIma+FVe+a0d2SsA7naUu/zQecnKljI2VNdTXbZAgBAIjlB+
ttG17xNmxrV7Fh7RKIq7MCrBP6qdRZu1CDtOqmTfrnh9QwUURai1F1If9sVaWIVM
wu03+sK+yzjbLZVtdedUT9pcuXK/3iqqeUFHbCjATXTIADkOPKDEp8rAoavonW74
jHTbEHma8cPDE9jOvDleKJpTvvWCt0xORvTOecdkN5kXyHY6xXLQ2afcf4WrMSEU
YFIEydyYTAtvC1K38HTiuGMLuaaWBTKm9n88EVrGy7XJD9Hm1yR8ntBiMhHSNykK
dIwWsrQM0nMj2byBfuvioMtqYl6drnmXUbXAeHHdVn6Kkt8osa3CDVQL6n6GXXyY
LoyQE/XGFNp7Lkp0g+1vV+/FNJK0aajSsYQOJEMw4cg1qw3QvUIwwnV/sVNCOo84
6QTZe9LJ+4eyNj3sS2MoXpZQZdulke3Y9uvEDR6rcJp9rXVQrnyUaAQc+dFel+aa
m1E0yn9SKaa4P68nDukY1aP3aS/E95tTk10craQWHt78ihz8GyBzTmBhiRExsBvT
R4cXfA/kvRZO9S424f6NVWGTsMLC+zTjWUnjYMLeymXXLcNrnZMOmnFSirXOpOuo
wF7n6CYFgCbo8Zq6FbFkVkvDTGUGLBWuO8KQwr5ALYh3G+4phAfkI9yvKOieHTZ9
9m2WebRIy/bX1I8MGHj1iMKvTRZ4AG1EbZGiODE+yn9JoPVg4rPEyTYM9yowbNqY
4JPxGZF/p+NZF5fNyuDkx0fmRXOILUHM4+H6BxRfMP/GhdZhcbZrmopRaoGX964t
qoiHVoeEbfaMZtbWJY7Ix3C2yLtVd4VTvb+k46MYpmkSTGGeM7NcmbiummUwFbUC
9Lm80t4tgfHuZB0VxNhVdT7uC8Sj/+d1hY5k2nB9TSbCsT5trqqTltNWkACy2x95
e8c8ySLIEFnVHRHJjY/h/IPavnOWqF5mVk7sMleNEXlmwCCDNIBoQgl1xc+iatqj
+40YUJTsRC4KhzsCrnOWqbeAhngwuQvbmDSIw33/GAnp9Ym0SJoDxvxq2FEjmQoC
QatfSPqg7XYkfiPfvXFv+lP755UieFvAaYGW2pInCjMpB/4NuzZtLFBe2iFhIckS
hHuIFAXzM+5PzqrtrvUorRQjxGRvx9B/KP/c/GtV725Bn9k/9jyAE5Sc46mqLuFv
At3AQVppH5hvekQKWTk2hfKsufztAiDXyMqSPivZH2dJVrkWv447DpUc3o4z/zG6
PIAGUBX3pl8JnxqWZGS0UkDSP0gAla4Q8ltFWY4rqvSIKJX+AL/cpvarEZY/8Yjq
44ZZngUtGwufPQoc7N9pN+6mTH1sAp2PKS9Y9E1NRbPq+oBSF5aaFzf2dSp6IOHu
juD4un0tzqVQKrgtGYq6o8DNk2jumbJkGIUasKTE2uNe3yPHKwIVDEhMEwqeFxXh
W1YtGeM97WlVmKSCjIx48leS4/Uk25rJ/rN7WGQvM/fPcp32e6P5CplXLoPIQSTj
EQv63ksQ7d1JrVYDYUkd0mIljG74ZBrC/ZbF0Uj1IYWSSVtn9XsMC+DTCXDI//u0
Vnj4ldWhBvEZQWqF2VeGVvWAxa8vIWtGJFii5egF3HQfH8mipGenPYV9ebnRnGai
nLJA9NePcGU+v3Rvz8aJmvZmKnX/0lOx1Qhg1ncCrbduh2DNOjMt/+kGAYXejn8V
LNj4z2wvOyaJxTVe+gW1m4hH9lNFJAwQXWYcaPs6RSvo/e73kbqSEF5p8YvVnhHR
IIhlD9ADz2Rqc3eXgjypQN/jopVWMXSLhdHN0vC+GkIoVksMPzD93JY99Ibe+Lfh
7jh21pGIf+amSk+MfrC4PZXOkXOdjynuYL1bCVKD5GjVqRh9SeDDvZOrQzErf/hV
mkyRyynEQuSGCgkG3v3zj+xg6jkF16cjyTGNCyItrZfjRV3dS8PXrAqQqr4eihfy
W7HETS618xKaZEAgFVyaJiekzyc48GpLoLW4FctDWnjVZUhBbq08Kaa6AnQ+rZUd
UCp/4N0X5O8aOqFaUk92On5l6CtPZ0sqqN1mtIlBchyX9qVEoS0r9vjFqX4bklO3
eu0dkoc5M4ji6WekOgrO9ttc3Zj4FiQZJFVk5X/dc9N+7JmGfJFx5JGMNAVL5zM8
NC4LPxAnPabQXo7JqY6Ct0skLFRp6ds+2gg8xdA7gv8pRIz/lYMI5wIVH9UyUv45
oEDICPksNHUkoTxfNGqAUXpsbLcMNsaeAH+RsIxBowoWdDW7iwZtk9a0O2oTeAAL
qZzxMO2/7/IsrJs2E7/VATzAXOirGMXO9ZHw/VbW4gtG1jI4sxRAYCB2YkURaOCC
xY8a4AcRndE/QpjVtE1k/TlG4YB6JEVglEB3v+P/hlM6PWIiu43qby4ztBmV8YRn
VZ/SeTAIVDIZjUYUarknNht3FxUDlupHSM0FrLb9n4kL0hOdMZ0+A+jITpkEvKO4
8PTjyq0sRWTNZz0JygOYx0R9JtZP3t9fp3XoSPQXCV/QBqpBi8db0Fuhwov2ev58
WryYE672QbV7LALGu3B9/nKWKsj3NaqIrBX146xkrZArRI/OWGahZIcOKHDTyS+k
lHHaajqIdDDHmb0VcAp+5R580p5Mf/bu8aTuwdOMAOrRkCXqPsrDQo8MrxMx5hpJ
dTFRiT4QxfrTMNWEYJSt6Lld3Ql+YAjks4yB7Qk6ZPzeKDqUYxs7OvtoGXt1fxR8
7dYPzd2SiGdBsr7ygoAZsAEMXBtO6joVjLa5yvNAvxB0uq5n7kQFqDpfxsKI6td/
RcPCm9qZTMEQawMYbAovGvM7O+99Ete50ZppNX1tbWRW/3PUotExZ7ZqQtU+1adM
IrpRVsA026kW0G5uYig6jPBXkWM62C81QMLmW4ZuKF3iM3GrzovxQtR+Sn3R+bhU
7wYPJ6jCjDVuC87rguWskK9b9JJqgj58ylFwlP6gOttdkQBqOSv8hcnmjjmB+gHn
6/D89fCELSrrs1VzLgdi2TGzG2bUFyuR5ivdbTaSZGbAIKcWHv4OmJcsvri7ta7D
EpxXyA/taaLnfe68/VPPy4jdjgCbYTPX/81b6QtRE85YShNntqp+hN7FxL3pJOi0
DgPJmJh+f1SplMtP1Nt28tm3XFUe7FkFvt/05SIty1/2P+wP52LkQIugmuy+kxHF
kSHZ1Lz1NcHzkKlOyVO+GwwuOV+/Qzhcf28flsHSvBxVhkr6/VePxpFuS252ahlL
WV76j75LDMedr3GSBtfBFbhMLTflxJzwk1dojPMRCvRdqA+csDRfOPw/Zlmh7NFn
E5K4PQf9XDvg+wGyhqB8/s8foz9aNTDDq8+dm/XPEc8WItuA9ItkEJB6Dqq4/8d9
F/1ZT/A9W3DcpdmyIBGwGzJ3nUSoWWWOZjFQAgOTEfwSrJ/QXIl0WCm3uWNcQ0aP
slNY8qz9oLtMQETNFUtUSBAbqanphjGezgV5kfHV2uWg6Oeiw0Who4a6NGW08OzY
iZxqlRHuYqhn5zQpQk00JoTwvHxZbB2qOKNPlKsS4s3L8NXNnweL+fM9uJq8tPLe
nfbltj3Fq/GEE79NzFvC3at8pdbeYXFVwWgcHCIACA9ITWGNBW6eDqKcoAJazYdS
2as1ADk/RbIAlVLOGf6UOfPifaafmvYuxvpHma7U1RLDWG64ydSDl+EuD7X18qW8
o03lh/6ttVw6GHo7LF+gVwNXP2o1Jda4f/WLFCSvOKwMAzxshyWiukuKNoFu1wPD
tNGstFGrNCXHXipj3dpw1pvCQH4JASUllZZZ5uUzwQ6yuFlnmt9TaxLGIIf9TWP5
elxxtCdK3b59iZ2eWrjqFYKxRsZEISNVoRCoxqE9IgsDMK7BK+h2rWG9nOUs7Dr0
4/8JfZQNGdTDrXsJ+ZiuLdvV+NkRQVePaMtJxOkbAd8ed9Oeq+BsncakLJ/36S3p
4/sA8oz8SUMEmUjxhPqmm5WHOVh8iGL9c60w67B757bpuGRxn6R1RX/hMTplzD6F
Tn9W+QYa/PLF6arZpuL1BUeMRkGKQcYN14P2JkCbG0f+PviomAV4fQpK0hEMV7tb
4gMOO1x+S8/05XpLisffZjRIsa2SWU+KX65oVi0vOgC+Q/Ax0B+Ujr4QFn9Nob1g
J7uNFZ5Q9cGv9EYrDV6Br9pc12HKmzJyuR5z+Fbn0HZi9MNDUJRdhCx4y+Hd0CzP
/x2poMAc8PKLMRMxbYgWXgvZWWRJP9cFELQLsOhFg7SSCLRbkAZxuzg2MbK/+vYx
lb1rhRVLl+w6oCi4OBGGJ61S2Yl3o9Vycs1NpSgKhb0v/oqA1K25SpjpytGPAOLe
UHmhSpEUHtcbZrsdscRjqQz8L9VnX7aVU71uHtAA4fZV3oTzyaQZ8pXWfystePNj
eWiDjOvOkd/89vo0av3PpFSTc16++hmxJY5kwjuG5XWSEnUnKs9AiuvNqzPGM50q
HMsNWmnbl2Y6xpM4bJuzMsZ1IO5ph0tGIg80+Ax42xAf3ihgAdp3bQ0QX+hsx/tg
5Fl7/YtLXPnP9zYDY1YLAub800HMz/IPDJTnSY8dgqfNXasdxyol5PW1eaqB/aKL
n981LXHVUx9G6RZGrKgnM7X7AWvx4F/KPvRMDhtj1D3MzS29RF8LbQbqvVeX9CrD
5hLhvyYafnuh3tOH1BmvkFjnXtNhnA8/1aoJ3C2j3fXqD5/XNeXJrryAXoMxj3xr
/Un3KRFxv1Su8/h8fyggCzHW/xaltEpGU4Z0MRXuoBvL97SXI+iTp5FItLm4B32m
VNIEzmsN2E2AX4JdGI8QaX67ZAaUGyYFx2cgiOdS+MPCOCcdwSXYvX9cbdn0yQbM
l08Na3x2RhnKwk2QToShYxDfP9rCA/nB1jr9Romf5RS6Fqq4DqUdoIb3ONjdo//V
YANLU3Cl0oyrUJs4Gm8mruPwt2q4zSjj43HFz38LbwM0AK/HNhevUNh6nghrtu9J
rCCldxADHVZcqPTxMGcvXCDl5f7OvNLcRdj84TVscVaYHCdIm+4R2AdMq8xAOg8+
yKkDaNmCcjbo633sBgvk99pYuqcHw3TjlXmc2/p6ZT5r/I9w/fEuL0a/OEiBOlMz
1AfqfwxOmi/K8Cb7sOMNEUxWF0IUAVE9JX5EQpE92aR24S/Smvu2gI+mwq1eVmKJ
oWgbAf9eBzKuhgIwDyrpWafBRIomqQDjKEISsOKKvVU6JZocDM7pBIzM1D6Bj6wN
7HxmqBZ6qTg6qahBB3Tp/RXzuYydrwnqm1lI2e7mvo7cMPm0TJwTkuGi64cHG3bp
R0E6tvVWScxLAxPFUOoGIekNR1pW6dSHq0gYnx/mtTwCKwr0MJdfmr3rOioZg7cG
zOmNtHbpptL38zS5JD6UNjTiJi7bgm/Qw64Xtx65XHJudTonquDgVK0KbSDLWSWg
L2kSdaEmAaVuXEcGjczGHjXxK4OztpwbIU8z73e8+SVylgyQwkQrhVJx3DZ4pI5f
dE9lQpN5gSCBOapLICGzyBsIzpRK0ax2qFPv7W5ntOP8BV94/54QBt1ksNxVJhfA
2On4w713I9w+KC0xfop6SfB8PMbd+y2n9Y/IqVtu40YIakGUIFx4bkk+u8FDpNa6
hWEFEjflJbHfoONgdeHlXL6+nH+Q6/BK8GypAkBYiVTzfzmyR/dEntZxamuobh8T
vt6CmkGFoZ467cgsg5zjKrldaKC33DtY9wFDwxiV0bh9vVt9pVGaGKw6SH7Oo0V+
o3sdtmSWgs26J478qjUVzpjVZP9MERRR3xCqy7FHRfrx7JSshUr89EKVKvWKCvsk
aAkDvzBMwblS5JTAhslVtJAUP0YivKdTNif2jhWql0OYLEPA1ZpbRupwscYGljWn
71d9qfpKcFcSki+kVEWkwfdR+Bt/waL8XAl55LZCwcN3OalV79IKVsw9VINTdMlf
2j4p41YEW1CdbdnQsyNfRpC7CTuqaQpgGUVpARa12UKx5quYKz2xho32re2AkKIB
tl6s4NqSvurHlxZkbN8ISdg7JZ1rN+5ODT55wK8LLcgDVri+XYWzmqEFT2yOC3aj
zqtetRfQSnJPgzUEh8J1JLjQppQnlvK1Xt1quT0UbsJAI7E6M3lD3JiV3p9ZoLbt
iDx3aMU6gUXkMrOtmbnPEjecqDUS3S2RxUyfCcSKL4pkEpueR05tTfj0Uj7didm2
rigYqZ/HWDuEjP+4QKG3AyxahfM8zjdnb9TO7IWvY6Q3zt70ZV6Zx3gJNq669Ve3
4FIeVpULWkp4LuwOPvPhKp/LNLa+GcEdvKfyEbcaUsb3ALkVuecHx6r19XvtnJ+n
TvQZOm1LQeHk+zCBkO0aiGnmw4gaG4A8KnDIMOgmXHCbdDqMzhXa/JM9RfoZU4Ee
jNOC6bT/pig2496thtYXokwQdsHeZLcmTNP14ygQTFSIoyshGT1AQzbsUEx8tURY
vAeQasPFh+XgCaLT7hYlJaUbxUB4hkc77sO3kbjbMbWOQPBCDoJoEVma21AfmRAB
kYoAZ9P9Cro8SuddLn0THNMQVw6mRndAYMBYMG+NI6tm3MZh2ixKfCLNZEEw7bQ9
udB0PIzj4Mep3TlS64NOHUhtYcunGxaELRuFgKJ1Bk6XV+YieCu91Daa1ytDiSRW
2fCqBG9hoiQVIG2SzWgZe5q69pHxcm3/OVsw0wvbdEM14WDDxyLRegRo8nKNMYb+
IaN5zPJpGGffv44ZiBGbJGXNZe04yhATwHm5oy7kRmQ/lP2KoDxFCYzmFXaEpdMu
yQ1r15uIhf749/HBjc1BpVfQuBhQegABkj6awr1ZZLNe4sWsiEk2VAUDOup7FdvK
SSTjdiL3PXmGUPE2YtLHMhib6Eqj2dvzRURsr4CczKxy/91jyZuLSXfoXTkrIeyI
J4W1R2SPuuecBkhjJGL5G69hGgNyByAjsirWw2DEQMdomT7XSuVqhsMovRwvDdZL
w3FPx6H+IU1dviRNfjxslh8zj5NooIAI5/4ZUTWCLaEqbLMyQ5xaxA4wIa6TdA5C
fFmnYpi+KgZDC0gaz4ijS7sx+JuCTL3IyQGw/ogd3LTvJxGC0BTDsJEmy416849g
GBVELBDfvq4d6X1OBn6D+AVVtm+MgRtO6s4rbaYdtDIf7LDhh4lFlfqZBa54dobq
9VJ7bZh+LKzzurSeaNp+GtkJ+HZ8qOhkFNxF2yImGBDlHtUpNezju1nYBeqQeU5Q
FZCq+I8p1KE1pMSiNKg1aJHV2GERYBZL01RDw5+4V9nb+td6BPsUzg7s5Y6EIEra
jxWnhcGFxIzC6cKrefhy5Nhjuq04Q3hrNRb8dYwxEx+XKnAxrcgRL9u4zT5HrLkt
9yqqN3BCsHOqHHXfjPjXBA4W4QbWWj6BOU7qGywVvuiMaGNKRCqCmIrJmwPKt46r
JfAU4NARqO59Ui37KAqP6Is6+rKkoVQID55VvxBbw04nfvXEQAQVgh03PMeX1O25
Tcvl4BWgHIERi6+NFOSlfLxjSYOI3mSNcN/nIi+yEQyHrXrE4mWA3hdAs2xxn9qw
DAljDkM+3vq/Opf7UeJxPIAsN6K+Cr1ZpE5V4F192Vu5cX0R/TlIeKoRPk1x79o2
fDSE39n6NrntEVQmRu26+BpLC9Ie7lmii9SXXBv4ghTC7rlAmOfRTPIb4lXKqhD9
WGajqf6ke0Sh4JGX3ZrGgDVI/r8uccWOW1XhYr8ETQCo2DxeJTzwrxcfHU6uw35V
o0/iGAZL3bZpZy4D1CSdms7ZQWl4mE/rCAjLlPEhnkJNEHN3u1pk+Vg3cCI3x/aB
EGH+sPu5zy+V5SNX/LaGvkfxVVR50IqUacg6Gevoabf1ACwq1W612clwlr7WIRkj
sXJB60mcmqvR3dvAN6AoHszirSpd8IfaJ6HU0EDbcbdKUoy5wndt69t5RUKE1gve
S2SHuEqtaADAwa0LuK2PB6P8HNfHYzmeVFxIm91VVPT0NCrOeT2+K2p5WVPWHeiM
taTpE4rQEJbq+iYLtULEQKbdkX/+wKmRSf4aQ5jfrmeuXdCyiuV9yYpzw8+kNNf4
Eo3KpIdMNONaZ0gezwleY+VeIWWNHhoZd148alfIBaWFB3GNHdjbcQERm/dxaV/M
CHql/n4iFmqc6BvlTId+bf+eIK6x3Y11q8C40CXlab50LjDsESHySjxOdRT2++Fl
r95HB3UB1s+iWnfD6GnJDDKjobhpMWEWVyVC6Is/uJkuSfZBL8lwmP40IYhSDtLf
dGIZAbpGehA1lZlAa5dPWxBDQRd06dYlpu6neMYDY94=
`pragma protect end_protected
