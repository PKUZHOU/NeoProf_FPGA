// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Odf8ZHvyB1q+pnUff5Ei9ijVd+6hRkQUzTVoUNkOzliD74fctKfBtzO0/3VReTLh
wKvd7b1WiYb5dBR2B5kv81YeT/jxMDgujv6MiZnGNNvDEv31UFLQRrpIMHiF5+aM
YNHzuPY5+OCXKGYF68BF9XMuHgSiIIiDJ9VM5r7MfoWfxABO85NB7g==
//pragma protect end_key_block
//pragma protect digest_block
N3mbFF4Dl32qqyfVOW8XQwTYgVY=
//pragma protect end_digest_block
//pragma protect data_block
4yUME+fVvXBbrbVJ83yD+36MMlMLXJsCFmgUur3ToWZsfQhrwcy2RdcUnpXs0T5l
K3oukG49Bgzv4DXlr5BLE1gNxJylTUXI/wspVewzSwBo5lEaj+wpzsuQAicCJZFZ
gA+qxbIdF1cGX39wc16ZKeYpd1mQFx3tTHu7GBKOf64INFv5lqrwI8COsMhpRZg8
DbaljO9hh3UhCpBN+8ITksjGqmVt9DVJVIaOpsczMQ95EcjFq2Vln8XDg55+sYIQ
IHqOp7cYJ4UnRY75fWb68wzAbFrLhQvhOsoxY1EXP7VvFBzoUTDZzMoFjN5Dbyvg
tQBOqjS1LLlzl6iuPhLv1UVkHPqLCwmNMKHPBn5baicyUa9sLGyDVq+i6kOQMGDP
l1keEW+P4s9ko4eMGBr6x27lQPohX8b+b/O5F1FhVmEOdEZQGyXhb8FJYOrZyqhw
gWeWT+WpsP7sWOaKmyEgPO3Kclc6lN1s9yHbLK5uq+6EGcB3JpLUtIZQg1XU4i9h
j03ItBKq7+bFdzrcp3syVh+cCGuc9dgN9b3s8xoNyV5IgbMXj3m8y4/p46X/fIkU
arsNJsaBy+A7vH+xpu4tivh9q1j5vWlV2JUQKG/3wsw9NdMo9Vt9kUQv4vKBWROl
pN7qUsQ9oVSIPmWcls6smnXO/N6CFxu9EZtxul4+HEVlQMQK0kRK5ntJiZaUQkns
wSU5zsLnTH5yiyn4yc3+LU9wG4ZKisVUXQQsYO6xrDiYCMOOiYaAfna47nxyY2ta
2DvG0+xhPwm+Go/kqqKJkEzWpWfQ/8tp7mfeP9prT/RVn7/6GuUoeB+u9yapw1hF
0VrCL/1TOC9PiuJsFZaCiHFf/sl/Z0MRnBP+RKnXVzWliuu7XJ1Y7E7mll1LAckF
qckS6+W52lnPq4vf6AfXaeVXS2rQQ4TBcZegFL2zx1WoTPjyifnAES9UFT0Pqkjv
kwJDcaEHnVaZc8QBju6A2SQBfheEzLD50wKbqsS/xLmKG/PStUM5ir/o4nDkPz70
R3Sv4Pr3FDspyHcVwUMyLGkKHML4pYpBnEBnptnTZWExrC5mzC4R8Z8AAKCC28l2
C8yYdp0CtJWpXseB4G1vQeyi9uoUOpyH0fBQRd6g33RGSTJm7RMLItPRCF8lWnWq
rV/tLonaZjrzveBdtaD3LEngWZThGQAYJMg4bJN4thbxvAHfZkxUsm6LxkyWwHJj
+g77OglQfKEDIb7ufIHq4GZY4eiwDRlbjAGc9nrOW76piahNIWJtdzBSM8JWKnUO
BdF7Sp8t+u4wcHZL5dfuK2JCsC4Kw6ODgSU/pma1YRU3jedd15oVr1+pyDc/GQZf
ZQqNIPjnEQA5WrNj/VZbKvAkFNDCRGsoCvwDPgjl/u4OMzHOvlKmXEIiIiYbmsOn
hcKpCzqNAE2yspkvQU8BOD9dHSwnAAZTJIZ6PgUTEpVRYMzebPGkXJz8Ip4Nk62n
fXmixzZ17utkVR0cXjklEtF5DE8Kctmixy1wEsJUWmRGTvyte0PA0L71snzWyX0N
lsJalh5aKhgaloxnU0lw+U1V0v4FR6B4XNd96me2XUC3dgZWE9JRwmb4oBecJlwz
Vbq6g5DFY9QjgVhGQ5WaqDT+cUsCohKizTbqwhG2kxKtF4gnLgccC1AcYllPFZrA
BXlMBh8LImsvXMgFbj0cXueqfqhuaQqtkg9iovq/afni71f/FWixF6L4WtQMpPmZ
On9WxUSOSc2saRAuEfCeVNpjdtx7UYafeuL2vGX/PaqQ/q78/tLfSIZ+lNdOtJL4
WypIS5dFQTOv9Lfru7k7aIuH/XysEuyceQhBDd6vtO1t1i/EK6sdBQ6eNgvqlNLc
9ZpHjin94+H0QDeRI8aPwKxWU3UYRT8qDtyrYNpNYAGjL1YqjiqYlyds+PatAGtL
CX7C5naCJIz/saH0f9sKTt9/fEOzxsouX6/X1X4bo3LmIX37aA5aKZNGjM9ygZb0
ryKLVHKz50zAirHSHABctqpXNd8ryhKmS1KSQrjFdrRX1DtepJMvJnEufROTpnT/
xqMFGQ/8YR8ilntvtcuvyuvsTDz11xLV9UEti1xh1uIvQQ3MhNxIrnhL3lRug0ns
YitJdutEOpBPtc8FBP0vyt2P6FQmpJYhlioXmCVcAMIugTdzEUIPNXgEwWwtPFQi
fDJ1LLrZSaN4kDRNsDl2nK6WmHsPtSrkerp2/94rJRwd+MtfSZIuidvLk7Kwabp6
F2BpaXYv0Mhexk/CevIXHovhNv51FQLANyw+0+WzKYPa4a6XxyyJJjcDDLGyOZTy
IRekOtgNi0Ir6VmZWcYwgZJ2LYAprTpGaBp7S0nuAicMLHDRC+P8UTdENVWb6Hgl
7BR3RwxNSblot+1Jn952+z+6nCT4xi6oafFRslmJRfjKowSl4bcPMrMlLYjZxLv7
0Iu6AK2yU/hzmRHbHOKmzifcpeRBilTK7ao5JRzn3B0aL/95Hg3qAKgkojSWSsxy
GcaoQ+H2IJ6EJLXChbnHBZ8t3Oxg4lRtHHwqG/dft1w1MRLaQc7zpV/V6Frh6Wcz
pJ8xwS1qZHdKOobxshkL1xeWpXpOU6KSGZcuVk8bS9+XQXmfD1kF+9lj8jn5jWvw
ttifcug72gd6PdSr4I+VqF6qx9qdKuFWIJvav/9zrA4xvxGR1+ZFXiqfo02hdLpW
2sNaZQrfBXPCnHTjgpkYpUR3wcgZ7UogrQTrx+u9PqywU/IWcl+8WhFeMjp+ZpFh
ZvzBFivQH1o+biOhqcz6KGJGw6bKQvmd/A0YLXlxzCsXt3Jy7fbMeCtWBZWDD/jy
LCZpjVVgeqpF+hXajj1PkmRR3m+CG0U5QU3aehYNNhcXXT0N0maw5GJ3VI7lPSKA
3KpdteO2pwy7PKLP865FbInV8HKiWa9YTrKDEbJT7/Gu5ZBhpA6CxnD8h1P5ccCo
QRMNLZeYQScDorizHZBN0j489Adc4QLa+nYESMTXPC+BAYAwgKGJxOcBlqhc+i1t
mFabacU5S1uetUC+IfHsmetuxmj+pPH36OMUo8FkuBgkUQDlDzYTTwTkJxfGwU4n
vGH2UKja4SNJhSoSeRSSnDkjZQ+JWgrOZ2FS7W9jRQvQleTvkREHPyK4QRfSll8S
CFkwbmZ0CVwAZc2tPJ/Jhx/3Bw7YXdO+AQ2xy+t03BiR4eXqq1NfeA4HzcqdsFnM
UpHKBk8xP6GG5WpIRw/8nbt6/Nqk8D0v/mTLIGVkJdGJZLLw6Sy47HFRGfxfHto8
/X8fJmRWDyREudiwW9PJfMi9nnm5Mlp0uNFlVGJBr3xlEn47ElCfldOn3btYw2HJ
rufSiEETP5bZn1E/gmB+1OKWNQ574d029AZClzP4KT/GiWncJR06VrCThhcOQRd0
fDensjA3KvYgQCgbGEo1n1Nh9J+AzzY6ZDqmeOdujaHESiVbTljWlQy2mRrrMtq/
7xNFOgYzs6rsM1ipkTDxMNcITn+j2stFa0EyHr34pCgR7BUsDe7sCl7kIleQTsZy
dA/xZ3pSZzkNRUhufXsHnUNUMcHvXxdG4YHqsBnKoqZQdSVqJ4/kNv2gMPwYL1lv
DkFAkgoaRhfrc6dLdoAUlJdJXsg9cEKysraJDUcBwoF7vxLEB7IutU442o8IHdPb
seqfiem7ToAu3TAGyTPjd7BKBp8UcdHy/Xv0gKbfrixUQyxb8iZxAcOGcDxsMrmw
ne2wKoA5epTBxOLrT7+duyK+3kiWdgZ4Y3/tN1/mqEIspwIUkOqldEZA29tyT/p3
tep+Omc/ugmLwOLtaeXgfO1cahjLVeMcPjTP3aMYvlXB8bV3ThXmqCjmzP2eau56
2aibcpCupu2NMoIrHSK6p28Pgi89S/SLNkNNHklPh3Bb498i0sEufC9xUahZLCpp
vHMOY4zbnt/tp6XDLjGLr9if+vCv3tn19LtrAbc9cMxwB9mFdaOPRUiEFvVPpMsc
/RJkLZcKcbvsLnxTQTF4P95L8rk66V7HvP/3Y8bB3sZZD2MFE66VVwpFvxrVlCsK
RizKjNHL+VLrSu6c93AOOm4Qa6y6eqOwXvws79kDvyfRihYakirGMWVKCF6dpxIc
HWtAm8H3RpoMTpXTNEPYqKomxXOQwz4DBks13mR9xKjOCzkqFCCBEAMTRiOhpPlP
FI38iSfLF5FroG/41k8190voTNOwmHer2kf0BjrM/4s4Io8SpH6HODpyziIDCZIR
3iJMchgKfWiPiN9hW79VbStoXrjVN2sdINhOqG6Q2OT4HdSbUqvGVVcKggYpaA1Z
oJv89lo9Jf5ImDX3DPNLlLdOQKOouQy/kUrcwIUqtrIhKLC8mdXZV0DMHnqJLQbT
aG0jRUwy80+W0wyRjU3cpl7Wqk4nRAWDevdXhQTmAOzPTNcwDKdooCrXiB42qSEo
eY5gib44fM/IdWSVMCyp9wiFc5F805Xa1ApVe/QOkJXZKSv0AWh+3LI7AaxXu5lY
jg4BZ6TsKIR81taA7hQP2ZkHeEJ2AfwWNOrErJlMgEqIXl6Bo5/IrNEmv1bM9c4/
1f/2qz80lSZ1lR9kGSCS4sVQ+S6OdR7ywD4j0uMl1Bj16CYN58p+9HA6l3rPE525
1UNnU2x5zs+ZDivkEQIeKZHUt73jXRAuNF251L3wJxpXLd8L2UtFC14hHuMJ5Lhi
1ICSeF9MCjvzkUOoZYudAEWbT2u6A+bIwqGjmYDnb/9eOjUwdjNViyHTXuMYDE1e
E6XUx3HYYXXzvdqSo/+k+tP+GShfB6Wo6IHr0+fVRGKg2lOxo4rMi4qdHXgJje4U
E1jrcPc1ZnNzCwr3t3sUyFZeBwUFK3FJZnEkVT9TSho38kO0XVvl5ZJ7wUoxf/KE
ah9F8KM6grpFYBVrnek7l33nz4It1VsEkr71hQsQ+O/AbWpnhQyWfVKZQJLzhLTf
zFVPm7uUb5uT+8qlRVvKf0mVfvcYr1ILkOqYteEpB9z77lvwGRz+ENODVD/+N1RA
X5FCxg/EPWkIu44ufAzS+qvnsJbzuin/A7xDyGiP566yNpG86I2LuvSfLu+D0a5Q
lyJhfbs3rmTd9WxqphxfdF74icARjftq8+2GUNFg+48LG0gkQfolEZKdyAwAJynV
zu6C0hZmPCTKm/rE7yuY0IexSccSWDAQ0I+etzAjHlXZogqep9kr/uBTZkPlP3uo
WgmX4z7ZLxmNr3BfVXtbMtkoLeZ3BFNP+KCJ/Mkzc+ERc7qpOmQBoxaU7OWX8aXd
9Y/44SeDd9ruCHou5wMlCFOVUjtD/Hn0u4PVmkYtdlm4VmSWmBaxCjyGDEdTd8sE
1HK9oVZWWghiNvJxKCo6HSiuFgWjtSH8rq2qqVxWxky+j/itOzlYDc4oaypx0bQd
ZjAqI01ROvEtd/RzFJMkz845BRdzLe/iEXxWyVdciPrpW+AtuXvkuusZQCe+u0Q6
beHT01LxXhXYC2qyAvXK+SEJ5dFOPOQilZJGuLHBx4hC9/zupSY51RM72NZPNoZw
a26h8qMJgGrfss18isaoRfaWZAb0XoJRf4Io5LskWr/tf5VvGG/2cAtZtuf3WYoP
prlyt2EgQW2jWDEM3s01aGfdBUWMVEDRE+sY6TNmIdJOweKJvkF6iIQOMOtFbXTn
CPk55Ooi4I4nS7FXEOqWx6+gM7XJBI3e4SXZ4+0yhZrxbxG9CWAyYt0255gtmfFw
gU2N9RKNYu9LV0vpC3kr39vbN88n6dn0lC8NWgALzKtEZ4Tw2d1bNzqk+6OmvC9b
l4VsH7xLbRQLH1i0CGWA2rf0EgXfTzLOOjADsAZs5Dw8NJof2Am7/DC3LHAch6m8
5dpm4tXrT7tVvL8iqpnKQq4Ttt/u4wi3oZJPsifGfsJwYfiLm+gUcez4uf7Q1jMd
VKeLGct5Gqr6Ev/1eJ1Vo1jMnUUFUoRDxpkXV68pPNqRVi1y+ZKTBDkpT9nSBInn
hB/1wlNh7V5RdfD3G8Xa4JZmh60X8/J7qJFYUJae6euf//Yb4Dks3umXrij2IJ+i
j1ssk1U9tN1zy8DNlIm2idzqkiVNBAofNJ0+0CXs7pNyLeNjHlpCJBJzMqjlMcXY
YskJFG6lGF3K4vl4F3OqWbdQF36SHAyYveyBcFHb+BES1KjdYlzM50UULx6zrCc2
Xa7jJCIQd6rJ2LLVc97aPYPEi02WI87026vYGulbnoIxXJYaU0h7inx0tWL41QSs
UKiufc0CopBnxrMGB5V4iNAHRKdfO9iLByggUjKImg7mMa4xcLEMFJ80Ik4phUHd
VUhYJcGSxGExtoXLFTfHGmh1ey+v3dHubRDdoJ8JFKMbanN8Uxl+VFybr61OHB/m
TJ06BMgkB7CCWgrzVJKqVDqM9xSnhhPFwlh8JBlDrq4DcVvLVF0qTvt+nlUv5N3e
iZVmlHtdRNZ2uce6xq1Z7PuxZtU0vY7rGuE4hpVO04wNCM/En5gY9utJuX11IH+O
ejLu3zLXBgmjSv5ZkmK89JAz+ujkAZnl1vJYjfVsFpO7ZdlfiPXaxtM1bjBGfLTE
stAfmAxK9IruRkt9+wOSo+fj052PxkplTevl5bZDcBIgEXfA84lMxMN56oeGDVOY
NeIXIMbRA9JxYptU28Gy60q4DfN7qvYLu5Wjz8lc7b9lRGkSsnf3VeFN8RxNgOeM
YlEFH0cuC2KYAXrke8gv1iRCS2UyvWkO3adbfTbFvojyY8Cmw0FfeoEmgb3RygHL
A8eETPWPjU5gzW9BZK6iB1eDA+z75bQw8DdsCwq1at9yiBnqgRKtww9QLlCrSwJT
PjH/LMogvdopB33fqdYWhK+MgtE8E3mVysniv+xYj2ZQ7szXREv9N7EUZErKMLMe
5XUdfFayJtk65CF4EFoSX7odMAC5GVSHv3B7oshA3F64Nw92nUErVIJ9/vUTFeaH
EBN0yQRdpBJVA+/Ybe6qer+gHaf3/tyxzrsacNQ5Gd7J19zWnzOLGK/rln7I8Ir1
oLmwt3IR8mst1GZr3l93UAEmas+4MGhNA3DiBlgpEU/4HLo0MGVF7rFw9nk3Me3j
D3wkeng/ZKOY/VZfWjIJIMj/SStvXTwJaiYs6JMgdfXpcO1ZYKgRHgRMxg0Ouigt
jwiSGA2lUkX2in/hKUZxSDOI2TONHEzQzItKqPxT48o8hbIQe5oSZl8nl1aFaG6o
s9g5DjNYqVkUSwhRHHym9w7R251HpDCIu2ccKA7P29XQxcUL2o/wXW2UAV5E8Vba
z67IQxq3fX7zK8gtuWAWmYwcrtodBqZAJGDmICOFPCITYntbqSoOJhXUqrdUH4R7
PwlxIc0oCVNxFufbpac/eCXRz7fGUGSbyL43hWCwlpkjV5sDDesysO9so4OAk+5N
4YAsZ00/35IyxOMrKGPcRzNzTB37vBM8IT5FBuf1LJ2Las8tManFQZekrLVJCxLx
0hjJabFg67bTjlUXbvvonIYOYo96OHr5uHOMyn5yoe1XwvYBVHJtmSGyKSxcW0Sn
VYJF1eJspthohL2S0/9P4b3cfF2NjGMsZ9dniaVjVQf+TuXnP11mCLpWwR54Zri8
pXE2Anq90/YN4QAAdqYfYlkMHjj18RZnNrtyIfqOSqI4F2YEh5OGnjDhCs0aCz2i
tf9u4RgrQs1THK6kUybaUzPuQxp/ASOD483MdoPxwhjjN4+sH5FiXDfhzm2/adRg
vYl1eWLISWdmk3SZ7bpB8aaLYXLUA8TctZMcgHy7646DminyAsjuaz+BdWsZ/qnf
oVjF358XIMnuO+PdEgd6Y/Rs/ITK8a3ZAMXHpLon1+RPIiXW54D58W4HJkjBtzVq
c/RYjfSrXNOVdWf4Gg/9346UaI/dXZOmFbXUO1gdyfYmwgmJvqmHTBtsZfrDUOhp
SdGiYJ84ZxvNOAlFSEzJLH7sbfFqO3qTD3Kalzj1S2DZuryI37F2rbcL3BTd7pir
81w3gAfGVk6LEqkMTezAEbJFNm9417mce8dCtagjoPnsXWiv/IfC29qx0CcU0WJ9
PoVcG/BoGOHtjamS3wkFZptgPLLes52hhYW1QbhjAjTBKkDlUdvYxCbrem6ujovh
OdpT2EdLosec7McSh++RVNzPj8QtytKqGDjqUoAhqvdYpYlxAeOTjnyIWPU0HAbG
bvLH04FoUMmiz7hIHuccG897TUmr/gA+42Au+YI8JQmGMkm/aM2oyVT/nug10qVK
g7cgNoJmuHqby14WFEVEB9vR29zpNAtY3U9VEOqlGqfUForfiREFyCrwDsft0rbp
mzzocjrP1ywqvYJaGM2oBKOgJQvKGUtDE/7gqxlgpvLLQqa6Kdas8N/3vLMBFsFi
AGouWS2MfUPu6A8VN0D5XdqEkhrPUYteGDmh3m9lkZNSprA2qZlhYg2gxM+bWQGs
M5kGBQNCIC55hRwt0tcAVTSE3B49t4Jfcxx5v7vMPUAZLGD8EphcFKEi5q2FDUwI
ezQdpPEi3P9+vwKuk46FotYmb5JvxJAup9xHXNOYc061cu7FlaetQ+7QJyhAm1hB
U1PpXDOkI9B1tf3OVE7HNciDkicEId8sx+gH/BWoiK+TP3F4sM1Ca/LCoHFm7ETA
aAlM0w3UIwMbZKE8NnQBVmpxdDN685UdG6iYgT5xWAXdgbI3TooY61JvsXqQjCfz
OZoooRCX5pz9Wc1ABJgR6T5yPIS+QH916hipe9vbDoI5/MfNzymvp4TnnrwbM+oB
DlEFYPVRo+k8pD51G4Kq8pULJO9ZEMcWXifksYnzxBNfoocMnLcg45A6o5w4CdtB
UH++0/fAtDx89SW/GfW6YHxgr/5lQ3k15ZFp9QqfDSWgEM2hZUEpRz13jSANrjhV
rWFLTCEzvL/fHZ/R5jg6Bn61prgSuyUwklf/GPyOgGrf17OhMRb9VsmDtmg1vqYP
TQOKhyB4wsUutkzKhSl+pHAkPm0bgcYLX5kbnvDWzjQ2AdKAmzKCp0OTysWWeYFf
q6wF6LkJrsCt7ASp1Xd/sj0A2jVLA+BmFqYu+CEhAMq3uGnnV6O20hq0/Ztfp/NK
v17fTPTk4oYDdZLa6GfDtS8BF/EtKIJU1T1lK++80Y6oiSamKPIBTzpBrnic+9VA
idulb4cgmz8/ow0yAbkSvZsggFzTyKjRMt1jMRm/ZoLBn0VVCa0vGiJgpu9/WFgn
CmO+FbjS/VcZY7MwRbgwYmgHK8QNILuyq2I/JSg5Fb52f1WxjRzS6MIurGzKMZrT
nyOboqdkarvWh4N4rwYVYExHYPtJxM1Z5rLuaMHdJ6miXjsP1itmLgwe/QRVLSii
k1DpwOAK4rCj5vgF7+kD8xxG/BW3YP+8s4FB29QQxPQFll2pe5jCkVPIfohgcIlC
Xf0HynrHXRth40LEnz19Ac8Zs3CuyuQiywmrfiY27sIVyEwZTXObl+CDn3ojy/0L
w0gY0Hvaw9ecR1iNvtH7OtPzeBDSXhAW4Vxks0RJiiZWHDYmYhhUKWuQrBLPmDmD
fBafoSWpA9kx1E/KqBmT+Y0sjDXMsND4WjxwYSGDjrhtnbqHcHpg6p3BFC4SbC8f
i8wfQZ4w1S54wRXz2ZbUduWBmAsSschhfdhVbI4+Eu4mEau1EFXGXLpk1KbNn+j6
Wog8ywuPEHq3Ekojum5j1LrDmm+n3QQWQVoJaWXa60MNO7OSo3WDidyIuqasQEI6
y0pwVIqieUNP/Rj1hinhzwJogkxqgyLvJPwGDPuLQtA1+S+I+xBULnAvEFyhsWWL
JZ9vHUeBzsyCSjhPbpASbq47p3P29fDrrGvgPsVoaw5YbRASdU5y5MheVQY7V8N6
yZH1I6546QtwTmEabKam3qYaVH6nzJdsLCLbipIwxEWiFfboa0ZT7ZHcLHit02Xi
Z9IJz779yZN65fUDC/hpAxiGdHk2ePTdHI5Gck2nRyhQEpD1lOpHVu8dAP/wy6kv
8ASyjJ31i0ZEbOriOJKjgt8ZViLEb92cXQ+xJ77SNiXbXBFAjR6TO3Mrx4VTMc0+
8o2ze9vNzs5yj3MrtfBqk4OqJGcJq8xVh2x7WIohMT/e2K8in8A9RwiDzosI+JQm
Y28nLarxVgbbI9oJyFUR9TeHYqUAcRjzhf9LeKMQSpqTtTDiGzb/KRempE2EqVuQ
hK0h3+sl9/4iJtSain8AEPNziwlHOpmHUQgNNNwxZ+io64xpmizTtkJca0vSFUsE
15CVpRWTZavOVOmAwBTjsTi+gf6a9gyvIkvUSiquUpabwrmom+QH1JrrOpdY21HH
ILPexmtPkFeokjxbWMuIfesN4AMIRC8gCS1fuA4VMpIM092xpQRbHmvnqk9NmMpj
tTSy7HFQ4VKyez4hcznklcBhQy0ZO1aEJfS1ucV3ZQpPlYcfBYil/kxeRgfOUO9m
7Xx+M2Nr7VfSm/z/bdsVFSqk7JZMgcDCyD3JMiGhVl/Bvf+r+lTkI+jeP0AbgqYQ
CxiGaYpwOxagm498qw7HFG+CBknewiP0kFdhlLc+WyHk1/aexEBSMXAG4vL4eefe
RNKeZoTkYEekMvOYxMJj0bDBL+gcKdMVT00uLDV3+U8oZE7QMxWrUfhltrxCrxBs
GA+/I6YPAmtL7IdMyog5qY4xWPYE1QjefuxkLGIXRvT5dVNpnDWBU0X6NFCsbSPz
ujEYnN2mzCW6KvvfeBC4F3L0+FRaAOGqzC9FUN6SBHUjEjI/x/zhChIgnY/y/Vra
D9CCOvDTQJnx6K7n4uvqiA54s6ZDDXdut7RRzPvhM5fCHBsNx8Wq9m/JD9TN9XzL
FSqCM6mkQ8rxAHo//hlt2GlWXHHDP8iDyh1/wTx2ZlyQW7Mjp9El0nPOwpTSFp/I
D0wYaW6BnoqtLbcDDQVQ/gdXK14EL9tFChlZWrVZf/2UVflrn2okB2hjaHlVlhLJ
aNeqM3N7mlkf5WMozM6nwhLrHgjUxjk7CpO8efSPipYqaJyBFywqfjHvAdxaKFpa
BalB7mUrSdXQlOMZQ1DZ2cjhMuxGyORX/Ca/C4aA0d7luI+L04wjgSGCiwws81x1
CJVsycD2DkUPYp7BQ3oAXTjGrefRyjv5wrHrhMFteInUUsWzEz4bwh2jhgeEWzvn
P+BN1vp4cO6KIXBaSLXsFKAuzu4cdLsxdqL6ZHELs9nLKq2zb/g55bKfopAm/nV6
6SmcCsZlnuNJs15HAxudIsPWdqeY1m6Pb6Rir7KqXBZ+Rn2nVToiYOZGi1i1F/qg
rZeUhkOvhtld6//RytWZJzfZ0ufjgrZyFVC1z8rzzIcVmXxclaFESg7SK18fB9d0
fZAA57w3l9vsHT8fkPfoXZaLpIvFMU9eXxyavTBGjRXDySRENNts3DNFDMu/g4cP
f+hY28Z6KkoekyfSibqfM8LaI6oNhjBy+hP3SvROf7TN0DVG1pj+6FrQJA/hgnHd
gdr0LEiOged2cOODz9dKhC5u8avJfMsTq4+mNyW8mI4BwIae00FZ+htNTdj4gDHV
phdLigMJRlX15dLmCVEV3I46P2sdjBj/O+8zTcs8upeF0mZ49vWLjyliDJ2tAV/j
YTRIfpklI15ZZj5jyUvwiMza4k5dkDHZp+3kIkLEk3DKFAGZTAYUb9nk24tT2jYv
kPQYuoEv08pq2oVmxdaFk11Y1T4zzIAq9w7HNcZGZrvTcyFMJ5RIEd345kQMTOeG
bOrhKpOyw5wJfs2rH1x6aXt1QrpqtLMEldz3ZGtxOyHVV2+Bwyg1thdRhU7S80DO
2yge2XP2FmAo+LyfeGfH4TYB6XhPuq/PDZemAfgiHcsxGhjUBk6X0t6vcOszrXCd
ZReTCtkz/yddJjPK5yhvhDWRcqIpOPqF4UNIt37GzyJ1Hxu5d7BZedsdoK5z/34/
eRCu6kzW0C+sqG6x6l+TNLiU6rtrU98WZT4sEGBa1iP04gg4VfHNyHL0So01bKtN
hs8D0v0dJdO28mx7MjohLcOOCq7Hn7H3ZRb30XnVFNGDJQvQsl6lI8pU0pEWosc9
Y+g5ZfUlzqMtWWxlxz+VLn+WVUwwh+QqyqVqZv8s7UGzhEbYXDeGXCkiliz5+dKi
UBYi8uOu8lLEewWewkLWwUfo0qmjmeFgsDkzp4HSuHotoY8wln7FTrk69i9uCzOK
WaNGRDfzmMwO39bjsIjnQYxAh5MRLU9OK1AdWxEESko/9/ziUpTF5pXBRPWJd/S7
EY1pM7mA62GJQ0hB5KKQx1Qm7lgcCYIT/JaDguD3fOQrYU79ND3ZbeBGKCWSf08U
J4R91Q6ijKc4xZLODVb21PN6HutwZG5nbmC+LKsD/0uyKY1IVe1Vxx3FwRfRjHt7
/uAM8q5LYTL+Ps8sZWQMRZuC0c0/YMp0QB3vg/iFaFf0+R4hnvdFq81x/0YB0qH7
Ixb7tTQ0PUzZyjd/aTPw4yearuAA0Vcl3qnCdRyO9MGrbcSFiiNHjTgM6Fi+eH/W
KpBI46tWuPsLPCoutvsxdozBMR3jbVIQRMhAv+7xZFHHvgTjqdb/zXfpJaNk2H7y
kp9u/N5ttANMdze2SmRkpm2xGCKWhwCJtoete8ve8e4gqHP9Xmr7G1VFfjTkBJdH
Nkqc4hIkwkWHYzKl+aBBuaq1Iks0EfQJeAHCCbLrI3Ld9/oevgP9AL0/jNdrhLif
QlB3lJzLM8E5AxLh5/2mZa7TBUQhq39AT21pb7WctWpRsiZDoBJCLCaYUqruBGRb
1wEtEgmdSdeJQB93/xWp6UK7uT+FFN425f2u15HO6Z+TIVI6w10J6PrOposaVR5n
IuibP/5fon28biUpXtxxEnFKFY/uyqH5/10ox5O5V6vtaAhHe8mDV+Pus93Jb4kJ
M12bck+sevvsTcpw53L2KC2ROujCZS7LpRMBOv8lnQNvZavIINvYm2sat4Z4TQeN
V1xZAQ6pFh3Denu2ncxbfnx4EK9DZsZm9BtS4zj5iye1lnyW38Z1yZM2RUC5QVbE
8E/jcpXVfu6age4IGphmFw5k/cqiERSozrb5oyXnIoMX7Bjcn1DN/6FPAnqCYAxP
vl6a197K3g7muIp4DhGO8/kukVsw3iXzrREDDwdq+pJMj6cuJB+npnVv9I/44mYf
d0vzsRhw6CDl+Ar/5VaRGPJZcyG4PxeBxP4ERWV95CZIgPSGQGM+8nUYZP21cYhA
pPmcByy2ccoYUPeKGEjIg1KU3C8jTwD8lKmTV73fOrhxggEfL5+fP2hRhwzC6IR5
1XFa6Ttj3cLxrep6WbY0u3Qy0tqJavGMXxNo1MRVgbbadhjifUrOQh2xFLboNLyF
jUdP+EEp199wtIyPezcNWAlO7Dcn280Q3CP/RAJEktDrY+PIMIZ0zwmDdD/JYni2
ba82olNc1TPUhJptpkkPbbXGOL/en7KOJyRRE1mGS9vbGKjOaw5y0KFO8QzluweS
Um1tcnnJA2CfBg7WCoYRmN9Q0hipG8LLmpSbiqVfWRaKKeKi8Z8pqBE1Oz3fleBu
3uPp5HQ0nMWEpUtHoglrw+FhxBxUmsCE2qGyf6auk9PtiMLlZdgzR1psG9BrIm3E
6pNgd9a77PDDRuprdFC4+nqwN/kCqmL+NCvX5YTrSfwgGe8N41OIEOteaWgrH/lc
krcwyZLVgshgw7K4+GPypY9BdV0lIPXkEqYLxhPOXasPjlTGrtSFW1fFcKAXFDDL
zJf8wpL5k3k1fMl7dsB9Yi7p3fLyLhXnmTk+OEatW0A2A/ugy6IeYbG1niM1GLQV
ByTqVGMYFaFaEbIWE5cAJptGXV+sLoWlwfV3QxKRHqwzfDunCImAVW0rE6gvY4Rt
NWv3UCLXYYSPzrywVjQ+6zjrdxiKDzQkV4sxqsTR1Fxj3PoXNEhEqXrVOCKHgNCl
kp7nHSQthjr2UOtGwN0fZLSvpkh8IaOToDPm6DV8xhsqO51t5MqkAR5ChEMpNRBR
tI0tjaTjBiqu7dqkQr4zo1efcZSNEKYCCqCiwsZrd+ghAklLdO9+jNjzjIvHhpS+
vLUgme884bt59o00TwwgNaBdPgov57Inl2kSqqTNAHEoC6Qp2Cigc1Bc49SRjjgK
lt0jUTgBye3UaiySagqJPnBsHKQ6Vr/yRpwsKxjDPQXS/lRtC5gkrNnQK/S1s4oh
jMkOWmAGyLnGWeHMw/zyYrNfR39OdiKwx7TVov7/nVmQpEsqqu5I9mTmujWyMwkm
RmGsdkOdVDWSrHrtmcuWRGp1BlBh6I1GNLxI6BMdL3jALpqlaKXvOCs85i9zOp17
S+/ba1uToz35IBhrwMDLTvEnzpPQsbpvRv4ooG06RUeIhkwtn+RFZZF3ZggCXn4G
bJufUChPtpjI2zWzzhyxCD9/HVmqRo5lpyqbb/Giba7qzYlz9ORIGLY+c6YQ7iIq
+pvzWkg6r+g1/j7yii+mOX5hvBaA8FWQhCALqX48Snh1f/f02defRfAur/ptghak
ZUd/mUw5P18NJLhJRQ2f//9u+eO8YinlKrkd3vvc+gERJtC3eaWtCbpePavsM80Q
d/bhUzklBLv5jv1l2werBRW4Q4qL2UbWv1dhfc3LTc0mJaE8ZivnSyOhr9FPzVid
eK8rgKFFcOih0IIhDPN3QVxhgoXKq6rkDAsMwyoMVU8xFZ7YCD6QTcD8nwG/d9Al
68qOBF/XuGr5UlYaMCDTfknJFtqqhfg73T6HDdqD7KhvNbKJsfxjHvziU4Aw9p6h
JY1Nyp0NEZvNgFFnmAotDt/q3mB3mbpZ6PxiKD7/QMWlA+UdT4A1hGJ1lVAFG6mM
sT+fU3hWYtunF3FjuGI7/96LJWdwngY7SPeEV9+IOaUJtibqWFxQ0R4U7uIdDzsO
86azuRPWK0I8zEsaMjjS5Y4g7dvNhcJl/xFGR0TIlfIAl63rvnddp4sUJfi3gh4y
C4wSC7W7P7/U98+za9wN1Or8bIBwfHg+nieXjryIWkwBl+Ommt9weqsm51LQEEjo
p0e81K7imw+dZj7Fgh03D+N+7KClqIF1z65l8yg77HrpMSxU1VHLrg5ohjTmtOan
B8Pe3HRep05V/d/XcBYf1t30ufbEmpsfmRTy+/yzIXAClPXl1dmOxct2PokVTyUf
0zJ4zdyC6xlOADpSrYn0axVy8APQTANk16q7on/wzYmYl7Zewo9SIseiHh68RJi0
xACzw49FDpHhT87uR68bbgSFxYQb/Bwz95Nw9fa34Hpi/eC5ETfZ7kFPAKQCE2Lb
zTs9WBZNXUGTno/5p75SaM+JEe9ZGJcmCT7GiYoa1BZE9AR0+SILWEOx/etLa1a0
BLvJeP8ozCJmB15fEuwj+v/LWF6Ngzruy3/HGEX6FLENkeUBpIjdeZP2jMqwvMr7
X7MVnaUqLEI+SjXQ4PWoEv8uHPyJYgL6IcAwnYvaAbV9ALsWrEcs1TOwS0/l+wB6
+GVDGwZzpEfbdwyxw2AAiHHk74xKbJ9J74fUtLRNL1+tTuR/g87kzcHJDnaOOH5q
HuaOiMYuBnE+Rq59cE4cJA70KPmT9Gc3fjMWR2VSzhgZhIC2FhTRKmtzj704IdYM
RNZ9O9REeSHpFK36kbPeavMMgHM3GusJabhMh+T6z6QXuwLWwK8Cr3m9iKs0Efa+
C2FIxPPfmbQHKUkPnq+crtn9MZSh6vD2lNZ/SIxq2jZt41DPSpo6f2ZZf4s9odm4
337c4pjmXoo0dM7G95CEcfAbz+hutqPEvDptJnrSVGqymCYQ0dAUiV2EQTEKapBu
HH7jMXNi66Tf6aWzao3pF7P5qz4U/Gdi3AQyw5424rMrgmppXaJpW/pQRhkg5tR1
t8+Xies6AKaacZs4GIkXaDJf20UPwyVj2UqWSySmZUxNU0OxSrXxoHJTTfK9yu0r
vD9qBrDZ6/Xcncovk+IhfiQlj7cilMhuz2sBZaxQ8TnGQDxcP3zI3bcEjPiD0YyG
i0FQr32pYKFTt3cHaajeK4tZTdD+lp/PFkSUrTrDdI6IjaaE1cBQnrLz5f1D3Ki5
+iPgw/g55y8exJcfBgHLuDoQkDekZESiqDLQeP1a7fZ0Kiva6OuGlQwfj3j/f0Sq
xuJjM9bEajUEcyA3Z2BRQwSjh5a4R591bTiQo4ddBG7lmVyyXqRHXazhL6F49rWV
kCHjuSwQk7v15veRQ1dDLtpntviipFRhgR+8jjET7BArtJ0bbjv44wuZgjaTsUPA
YW2WcrE5tR300JANOLJcwDY2f77YhUj6psB5/BbdI8FHK5o+yoUmyKYG3h7RKSCV
IEjj2s/VKT5bCcWQ1c+cX+zycv9rYZ8CfUhXfuUsSio1CwhnE8qNFQtq1sR8eiZo
jq8il1btHd46Yogwdkh41kxO3nbu5kc8g3i54TMh6rr7dJYmPyvN2HwJ4iumNJ4V
Mn/YDliu0Q/BlDcnqff1pTgUTidzJ8qAx61z/eKW15yqVU66Lx3b4OpQ9HJHE+Ml
Gi80w6ahWLR6JBPPEztc/feBN0OBK8YNZrzGRXVgKyJhik53Ihnpb0HcucgAjJkR
tOBNcNwdIzd1p1qjIkCGMfeMU16eLJxD6mUs39FNh4wFXv/JaYjvyYrX0J76JxHK
E1NGGHgmhYji4xqOBUs6hl8T8PgOWV+YH3iXO2rcN/+SkZBxvMcy+XiNd5eiDRIX
UgFfplfj4XuljvSdRkrbBCgnQbU8m9N/vC3oC+RCIKSnpt3GBNENjY5l57HOEykH
KK4lmF3naHoxPnZS3P9QcEn2kDwV7aeytKgyC7zFNkeskSH8jdpW61Z4lg9u45VS
Nac1Jj7mzQyV4AzkJEy4kTKTWX61RWPdbC5Yw5oeL4noX68XoDFAgx4Pckd/+8cH
Rwg6nHerB8wAsCjMUJZSUDD8UJb8VlCslOOxn/dV118zbzs54yr/parm0ILDeINr
zDHLARWHIBQDG4YW//R0CkX5pAyoPUg6A82oa3O04ZNBgZNjrgMKSCs98x5QaYwz
gvyJdDq1Vmr+nfMwdeaSXHYeEemk8y9NxUt0iV27QuFgZUK9oCLNgaZ3sLLRj7SH
rZE1be8cjSiC/x6BczI84dEyApawfWpvE83nxYJn0w9a0tBiTY0sTMGN2qGyD9jp
4qAMcaSeGZR3zsklsXY2zdgrJrfxBIIbA/wdU4f2y4JjNSQa5oLORu4hyOnPg0G2
HVzZ4WRcT+DT76k+u8yw3TH2/izUuFYxgvqpSy5TJRhgGbc0M/yydvircdp7h/Ey
foDC/FvG52hojDbpR2TZvonYhA+89FsAE7poCz60q4yVrnFP9UqsW8GcnIC1z2B5
KKYlH/mj/M1FJr5AxnIo19KFNCFtuJVPfhuvOSXNVH7u/VoKtsrxfWE2YwFCoWrd
6dZWexJWTe6GdmcsN1/8LOVOFcthFRHrOhmdC6pBECwIjuyke8lZGI6E530NF0tU
zProvdpfpN4R8bK56Df6amdlyv5awQVGTtMPCXhJS/FhkJ5X+YrRumKqY0HFNlu5
tQpCMDaz8OpuSmvFBcA7U1+GYEAAFayYzwl+c9gl9Mg8ZTu/p/DorgwfOq5b+sVi
YYycXZicdIrM5xy9gthrJD3ENPku5J/fWbVqROMX/cWNV3A99V/DsMeFV2i6kwOj
puIhSn05LNyUlNQoCw4IaCMaqMUKbxeTVWSSXZrAZmq5DxjSJHcNixyVzqglIH1r
qsFQzW1OZ7SqsK/pmGWxKFTMr6Q8fLfEbBIagMqz55/RtnclWyxECtw3tM9mM5kD
slCQpxFvgLrRxsMFSREnsRJIe1jgZjz3NNiJ2a9Re1PB0Kt/TxFpbzsqZyOPt0b2
mRjhcZvUg+OcPMRsj7kPcF2vZbnF0MF01qxSBEforJPOBbg/PI4S4DxC8Uci7Kmr
xOaoD/NAFDpjZJ6xC7NwfPCdMEJ9vWvQcv7Lly4u9KljfbEoejoCRfmUa0oJufiN
Lg1pyLd6u7NBkXRlKFLlequwryPg2G7ECxykgwbHPfUdSDqM0USWfcKZYd+FZPiF
WPe/0OHS+Pkc3bf3GP5gjkdBl4a82OCtNTtC6nLyyKKVrltsfpQQCxfC9D+5n/iR
97CZQrHykfDwPwqh0//okJjOmT6LgFJb7+NrwP5qHf9PlRfgt/TvMmc+D6a5bwnK
E/dgEEFIfcqh+l3+R+YETc4TS/+f5XRhBxyASWf5m8kao46S1sTUbuMOvQ/9Kd7m
Z+rtH84U7Uf4JvoyD8WnGACj38jVZlM8nYzqSij8wMghflIJ8WuAIgzRCp8CxBk6
u+AiaiEp1OToCY8F798voyDW0K7oRJtHT7FM4MeRnyHhQ9GhlXGhEmgtp6UABCN2
m8ELJAVDL4OdtEvVjM/C5Oi942+w+a2d1Om9B9oAnhhI6IkMjPvCDYQs2HLZvHsB
sCQeWjgp5XLtcZSuDjUlR5kc1MDRpN49O0uwMFBWjln/kZ8qshgm04oU1HM7b/K9
zhgW7Fad5qw+wAga1us0vbFKKEOa3OpQs9Lw9S5pKbsUnWSSBFR4nnTz8482eN+b
S+rpxtGY/Mcylc6Nv3obvdMNKrQAtGpBa12lNZecJOe3GcgqUQF8sDVP1DxiptJ/
eSHLrC3S3fIk/kV2voH4T0RVCPbl8plOY4kJvuwrH+3w2aZ6MsKoP0KOF8/8XUMg
XoGVT/Mxx2NCbRPzzwamz4ddyf4iqtAAnqspTdrPBE7pljrOWfYZZR/YPhhTl870
mC17aJTQjaJXshBweIIeFz/FmCP7eF1TNOURJqJLSPRy/w9ylfA/KgGreTW8VJHj
JWHeFKgYOMvBq9A9lQX7qxosL+XzS6eR2xFnaSLRwjLRiZooVFY+RWme20cqp+KU
QKrHpJ+ihOACKAfEB/Zaj2FZiqWq2Nkow+cJVCGja6HalJFQL1fyMUVl1TsKXX2Z
ihxqf5EW8bp5j6Em1q5rRM/EBLGUG64Wo4GE8jyV2NdphGO6DHW9IFweYWfQt5yX
5+lEocxTJq6KJ5PXasPDGZs2fHveuzDowTDPfQRkjfFvKv7Semhht7T5XeJ0VKbG
1WFFCPz909eY9oEo92u+IhBcf5r4KaTqtSKmZ1fgjSRFTXPSyAZMEWKv3PT2hf0z
9vsVXYNPaNfVRf/Z79XpC3xocK+vCfznI7PoiBkdVo37jfHe7oG/gcTnI9qeW9QQ
cWbCKE4Ik9uAlAG+EHWt/F3dcrP3VGli+7qPVvCSU5fWaNCNlWc0L2BUsexFRl8L
QKlpOOrcViNjYQQZMnTk3o88bL3dGpp9IM9v+atOy7Hjs6s3DrixVANZsiHwMDtK
QXZB4P2VqrD2ZpvNFpIX+CKyFHm65krym0aJMrBzXy9yqPmfx4QjHnGwF2lfBK/o
OsHhlejKov+NIKiOAZ+igIWrKkvkLWk7MFTegllEU+v/lF1mEIc0fyLIswzyhEoh
pExEnTuPxeFnRzGxO5CSQDPZGCw+sXJCbhcy+CheML7sqpxK4cPMi6zqQ4XfGeFS
KcP4zQTydc6WPdwKFmza9hUu/VbWL5zopxEqKMMwiawmtVFJi/yJKLWGUbdNwtXz
rhd7fHTU1/BLub4ksWt46YgvvCnbJhEgJKgd5BGQGPuxZbJBYTJJMydDWI6VJ8cM
GxcHlaOQ3h4HE6NKn20B9TrnJjpD/CcPbhaeLA0/KHjdiD8OK1C4FOBcj2NrVHRO
M1yZOnVZBCseg20Xgl8PGUTV07m5QZpUSrpQgINQo/gUOjLI7knkTkb8NMtpLUtL
YERJCyPxfKkehla+bsKxyKdLQ4QV+JHy4r3QKNZUYcicPwKYOy9chMd+lk2azKWs
HyMHh8scIZKDz3vFknjh7rqMqWWs2FPfSvRCIAnnexNVbouUnxFXtnW0sQPbm/l0
eXZVkqd92hoXXnX8kM/D1wwacrFBb3fqrapau34UVHb4HtmzUBsstEoHgCUIJ9Ni
4ERoaNMEeC69keATer8G+4+LHRudPEJggl4o03O1XM/uxU6WBptgOXlWoyPWMWcR
qavK/chwN2nVOYxWzQzlSG8CiSy3AJQY/O8kwdwYwwNLW8nXWFBcsxr0vieD+GId
tOesAlypKKPxVnEO1xQctrdBS+1uYrRYNaNtApYh1rOgVybQFT84vqyv0ivUqQjW
e56DtI3rxzC3pRWMqOS0FJ8Sqsqm0lzBAMe6PjvdIAXrxnz0Gkt9KWZzlHOGWUlo
oots36CUgmgaz4yqQo4rKqGa2XLGML0CiTWjGj5szCfTU3QhQDgo+dMj1bV71msp
6EjY4CKypSpwzf59Ag4YEM2I1Z/a2kn9ESbjMFeKrZSczhGtkYJIzEz6+SPlhvdm
zDJ6BNb5vBw8leWBP9WZehm/Fi/55+bnOrC2sqgpOH/V+tu0bJOsvPgSOZ1fJ6mx
/gBImVIZE1phXrgp40MYuHy1y0W1Vbj9ByzsznjnVwbuyuCHEt7jqYTDg5aAn4hk
yR4OEA4ca+OAJ3jt8MNQ4h1/lktRyK/tss8GgQx/Rd0Xwg1xq8JPziQxWPMyt1bG
pwMsrUfj1pnUkr9YrXQ5an0D4XN24XKRdbkdMHiF5yJE8+UXtmj/Jm9rnI8o0Q0z
GU9cEqhpEVpDmHxPu4TVrhHV6BUkfYZx5G290q+QJLk1gGQT4Fwmr64BhGkHMNGl
zOOBs9jaWR83fLmYFDuNaumb5tn7/Ws+Bo1Wu/zLiM9WreBfJoOVztXhj9v4U8wz
77WqjhqO8dPsQRELbDLGi57W0g5suijnvlXqVj3H6N+LPr6Hhr6nZQb+EioFJr3e
8vcoja+ZpGpwzXUZYcEcEYkQv3rDlJoooRi42nz9VKRMhU1gomEwoqssVP1YhEON
vFAnbaTS3fnErnkfAotMr3m9Aku8FFb+q4l/Cl/ChlMr1qDMjGE6t1ixLbbFC/ml
kAX09rtd2IiQtYMREqcNXfyQWfd8jr1qNbGIj5kqozBVo3jQ04tvotFUWD6EoD29
+jS3nhATgK9IHgR94QoP/6KNAMcO3inD+igJ1oy89sjqtSE3+DQTAgw/F2+3yA24
FulMWcttmTtUyMLInUCxC2irlFHOPDQ3LeGVXpZ6l17lp+nPGshKLOG2ig9xJaNh
SocRE48NDlvOAJxeTQX8LZnusLJRRbEpMS8v7zX7aT8wcwF0/DKhEiuS196139LK
/9PdLXIkkU+7YuTLSidXNJCRH3d85nvdi+UcrWuwIygAMeQY8Ie9I+FR3eArDaZU
RUICYNJWb1UbIC91qJipSoQ3G35pIR4PYHmB7+c/xoyCh+V11ADalPU8q7RMNm3j
PSjip1+WkZQ63W7rXX/HbrtmqeINmxeHyKjlNrG2/r1H37+s+xQSCvZFpmdJNZ1h
dqGbK7Yyfu4DzoZj4M8zPuZIhDNAOKf1IXzomP9jr1Suc7c0DrMAuhjCzf5U0bWE
gdZcsKhaLfDApf/upT1KlsKXWV5mILcxaCmDTbgmmmZ3Wb0Wnt5grzELxo+xWZ5h
3B6HdJmqHA6BLxl4JlZpwx+kJCj2QJRhIvoBfMiisTzWoIhxCcry8Ug8KWM4wQvq
XBq04T+bLaNJq0YGbL0PzmQoZIbLLVc8HXZwSVfPF6U0kH6EeGN/xzFyV/ck0eHh
HrM+YOd8qd7oKCtJsNjulx+yRe4+UO1cULWOiDO4bhu5K1GQMfMxhx866sI5C/tF
ad4f2zzzr0SDe2762M50Rumtye/rk6Gl6zZ/9xi69E+39z9idXFmrEDKgIvM0SDs
FrPBssrwMrjZywcrPLNReBu0oS0kJluQk5UgJ75Ok8UEZaBp6pXsYRKB1ApIU0w7
tGRiPMkwGU1Bm4Hfr7ngREQXCnc1ZyUtiP6B+iUN0gksn8GVAfCWPxheyfUVh8Bo
O9st2/XZCVsBkPmLQARdzNDvn19dOthb3h0bD+yKARLqejDv32KSny9nEk5l3Zu4
Vm3adLZ0sl410j6R3U6b7MizFaupy0ev29T9lQ7TytBAtJIi24Vb6YGT66/TkCmY
z9KGvQw9ebN61V/jTK0cJQUregNzOARRSC8lriCrvR5rMkVzBZUvqOvJM9nfYACn
7soF9y2uy6SR8NhXTORPt/JGb82EmsAriI6PDT6DxjsLaCTiTUq+ZCAEdjllIU+3
BQDWYrKeqwyNnKBUDqBHClLeL0sO26UDu4kRrlNXzHUpWNdNy7I21UHQhM7eCKXD
MTszaQRk/yeqSmn5USxfHR5ERVQhRrvFA168SR5tP0lkVPqB66B33/pW5GI2voaf
WJw8+t50q14sO68kb/jQeFtbuLD0/du/56pXW2K4j0CAw82M9OOzTruIfeHfXMgH
Ho0HsX6zBOwerO7qkUjWvpWppUn3SULToW87evJjxci6QeZ+DwO9HOwrTHS5nqd4
2L8FFk3REiguRLa2jPWHwUnSPboZPMk7xJ37fCcLFgVCKPMqToxZFhjohMC+4GDL
8WXxXuMUMgonY1OPtaLmIMrggoMCRzFHAEr75wGG+XqzD5aMVQPoxrZAgh/BGryr
CBhfBm8XtKknPMDKnWFJwWsynBFOtwuFIy0aUm2yTLR2wWelSb1ZXSFWsWZqzkHi
6v4eaGWuRc2JChqftVP0w4wPbRc+kF94/M33t/YFExSmecu7nP7W0Lw5cBG9pSIK
ZppyRV+es4TuoUketxh9EEekMNR+SsqzhA3r4f+8GuF7b6o2Xq0HdNPkJYyesr+X
h+miuDgtng9NSH1TB00Un6lpw49fqNsqjYe4hHou2OCks/VOYuG/5lyfg62B2ejX
ZckLly7cJseF/gftzv4vdmTz7k6FZxvY3v++AhWqdZm5FF9S8+PupHi1rBMkPVR9
dH9xdutRp8U4Q8jZQkRDLGWPc5XxJfy/WCHdN45hBW6FzRVsLSLxDBwf5nMnH1a3
mLshDcHG6Jv/DDx57uie0OZ2gE/2DZ0Uc9Cd1+LAT1pTiPiWCLuCdbpMHhjQhbhO
tK8SL2gvpdqyAWZoIpdK0LdstIFx53YwkwP78IYqV4LE6XXs9+t9l+NuQ+G7sX7t
H1e60v4Qpj8rQAwFOO/ZFwvKC/X3aNpIugPAkNvvmdH3f4Id4y5rINeC5bF6yBvi
bx1U1cI+UXLOcPQd6RU+vj56NF/caHYYNv/tUOosdrZMQPJ0KiuMeYqtudllfCI5
yI92M9RkZT7yg81Hjt+alc+yPoxE8y+7InZNnPBDj/jVy39uZE4pJ/KfS4VMnu6F
sAzv/Ah/xxuM22AxqIBSdBbcD4IB7B+80t5JOIVULn1Oczx8IJ5gbydoF0yyHToR
fgOcDFYlRATaOP6cbKrkUY5EltDShSey4gMoK0kGhGdTjf++vpEwydMP9ixXeEqA
+00FvagMtZfIZV+Dr5cPMvCRvzXYnpMcOi+j37E0lIEIdfRHBSRy634XfsKUQpLY
65EUqAEzfIanXfPh3+nMxyOWK7ocH3meN65/bJpg/peB3sS19LnXAkFcLa13QjWb
Io/6GTFUEQvKfLSn2ZdqgcZMkQA0p4lMqnsmZr/Lw2FLNmMI5mEbG71kWFeClPDd
gYmDfPDs7DjdRsCx1hAZKQLO+qwUv6B8JWtFLNO5IM9fZtgmmB60lkOtHTVvE9Uv
UCSHqHd7qdQf9NbBj6raLTuGjKzMPi1bfJfYZ2FIaikCUpJeJ10FYjp6hroBu0uq
Zb4vadMfM+lsnU6LT+Rdt5YgNCrAz11WgW7GfSFzSkHmUp8mGGzUoDHRJrQ7u+HO
elqxEPhFw+oCati3O/mXcZRTY3mwOk027rN52s9h/xCcqA6RkaqqDavnBRUvHA2d
SjMNYlU8jPdFtBTyD4YIkG0IgRNI/a+c8G3Y/kYSZ2eR8M1oDQA1wYlPffPJ+kro
3vulp5Bc0x/SOKASZG2fHpsdDm12Sb7Y9x9mjujnpzDrEG7E5e4p3cbmGiBCcWo7
zayBLtCnfBmr+sD5ZXHwfpjp0bS+5rDer9H/TB3qUfVNCjxOBt+3bOGZEjVX6rK0
WwA1acujXy2Kqgbf79vYpSNs3uXNeIaCw+xp87fovXkxQLP3s+VmCdEOUETX+ere
CA8BtMkod9DdS0Fmn3sQwdR8gN3vV34DhwjyfzxLFe8aiz/eKZUlz5+h95fnCIpq
JsT3DNVQdk4HJw8XraiHzaKxm8eN93JxoueArKzQoALkPBQ1WP5wRcRAiexyOpwW
kJ/YoxyyTbrPF9YdvQDh+z7tw49EkOlcTfapZJUkrH9dGrASF8+fLwEgZhEjKO5j
cegAxWcnY+iJbQ57jIBfcILS2J2vUE7D3PMAn9zauaZpqe3n03gzvhCWV6vAPX8C
EKez2Qm1Oux+/9gsil93mAR28KVkhij5GB6rIRAtw00GRTVK6h9AeV9pdHmICI0u
b3uLAEhbI1jMfB6y55rPQqy8GRUik7L9CzQ2YvvkT373UDsZ5lMy4Li6G4Y5sNan
kOxzmWqCWQ9CN7RWvwGulZDGQis6wyArEurtMJsErv8Hk2cMFZKt3gAQzvV9Lrls
VewRHx+/xy+ELlU/GOvbOk7k/Xb0mLCzTogCUkcYdOSHnL9sgFcGnC7kK9kaU4dv
97PDxOKj3DzaASCRgCJSuORz869qhdSMyUJTqIIsj5aXwwF1s1IpfhGmO5LV19v0
sxqT1whXCWoHENY8xdmhkPuk9mvRSvm8/O7GrdiutdlJxLPhrBDlVSED1llHZd1Y
7N97nlC2T/63XT3gMwdw+GeBld0KAinUK8u0KyqFz8PMjkzOcFzplShI8S2Iw+qS
OOIPOsJAv9Zed1zT+P1srD0Q3Hs5Dn6Iyaa2T1Wwd5Yi1lX53EWJIwf183s5cigk
dZWWZNYQnhybwSCb24n8fLHS+HNmuae+H9AAD8+v8b90hzj+0LF/uFt9A5EzWKQi
rIWlzZYO36TyAS4NtoAiVnFbHMoga1Aa4ssy6SlpDJ0CL7FWS4UsWbm+Av3sXTMS
WF4II8jfnKh3IcJyY0uTzbEg6ZfmXIDpcwvA91upz8BjUMxDDQhVgaa8lsvu/W5+
biZ0yc5TfrNLgzWlo4vGp6FagSIIXatJHsMU9/EGsVfwjTaB+v2Gjvqt/mKZq2Ef
ndjj+iUX6LtW7WMU/apCSfZkFCUFkCQzFKpjnqOazULIXhTpUNBCFWLXCaT+Egnv
nzWZH+2SfDHSTmZRNEnQ2v/bI+ClJ5zl/37WQNuXQr9oJNRC0+++AwpJc+OSadNC
JE9Za5P1+GJ/fDtxoAZ0Q/UEOn7Co2rQVXQsmA5B5C/DcepYX9LPwO8eEONDH3x+
Ys0lkxoIvY4iBw8ZyMFDOXmNFWAt1LH8xHzjiP/z0mC7leXxLUQqMTj0NSlXaWq0
NuSRGRHyyAPl0mR+o/gB2nBo5TbM5difsnr50RA/CK0Ivy1ptFylWScbI2KZaV45
QmORkWSZ/+IDgRLyTLB3OgPKb6uN/RIVHoo0M3yCA3vlALeJIEp3eNrPTYQyUsnB
kGXTZEdUeJ7M8iDx0LmkGUWIWnke7cWlb4YRnv4iPddw6jDcD22/UZuInArRrlc5
aD4w6IffYB0p1sSSiTWofPEH2v0J01g1R5uV5AHTilehoD6pZDaV9Gpkkw66dO0S
oyGyIWsjgfkvKxsdFeS0283tRyw+vkLmD2c+a65mCpKXNZtl/9dVrh0WjLkprY9G
vSAZHUnNKDVS0VywbUni5iSZIQNQO+ye0UWL27mgDqh51ir9VU84sF5JSeUU8JJt
5L12FSSs6qGLGPKmRHsdI6lWEsICuno81kSYfQWVab06t39929wojwrp2l+UqPNO
T/zEIhmAZnkzeVAgEuq69jd0RG7mZupGgnd2W+40RE0tX/HAvu9S4pUvZ7nznqeB
QHAsuSs4NWZQi98XH/uGCNc/oBZShQDFSXFurx0nqinRTJz660yduMmbz2cMJX+R
PdY5VkiOr792qklz5X77z2s650mrMw6rQTnT8ZyewAk3sU/F5ih0lBGzBo76sTLx
OMZwju308wuHCj9Ew604XkYwOx7esLxxBfeZD0Jif7s2NNN0GRN1377KgmjYvSpx
kDqt/4yUldr8xSsnnty/WZnTLiJ59WEL64lgbL/3YcsMXEEWYguJEziqMSrsDkV6
hvSQDK/zM5jYzYNDZqco3OUiB0YnF8koD5vnNE6ND7sq5Ms4Gue1BXnQRlaticbx
sxZyWDF5kLGiPHaHUXGTOa5bBYjMcQA0QeEDXg+KSwka4oF++A+0biCGY9oyAPQ4
vrBSRNIsDEIUnQzoUN1Wvr7pxmwQckwBDxAFpBWbTmLZePDUn0snYsZJ+I9Studm
D/0kvNoqJ+o7O2KPbTqlkzbOAsEXJJtZBHOuleyCfRf009PVxkYrDk1x0mI4dCag
ijT83ykQlE1q46QmEkPaXUkWlELuHBiRYza7aVSBYgKQNWxE9FX3jMogQ3rsd7qR
ykZH9kx7472YD6NH9BU15W43dwo4w0GqO98CVxY/qDjCT3fCik3QfCBr3R0woYKq
Kavbt/4csX8GDG90h+UhhDiJT5InymMiUc2G2HxneZai7xUBwLl1hMUKpeTpcC8x
PoOLJYL/apRw92nTYfaHt5M6/wByLWOTyiZkM7khh43A6uLg5Z6XeNGKYekSycUx
Ryb5LMI1jGrV4Dod6NgMCEl/jeOis0dptepM/js1F0EAQQnug2A4JxgqWToYSoAm
iNE70KUX8tSW4a207abvivGEI4KXBJemcQs/mPlvxrnMAkjQa0AhfttWkqOQoVkH
k+9s1jAVmOUHdxT+prwy6MKV5mSYv0vmXy1N45xqQ0bPNbDdOrTIEBVWN6oBRCV5
KpuDkzL2kGQp5grDn940non4xtQQ1ZBw0RZ+kJmQSHV6mMhKwgzExUQ57E2Gmfzn
SJ3wXWqVp6cY8C2nUWzAinDkdLIYMRik0NiJ4WBfEJWO3PvCiyn+cAows0/rRjKr
h9C0pS5wC0sBE2cku3FUAemeSCLKufaxozoTCxEA/57g6DiWYneRqVb+1nz6Ms8J
6N/iBAvNYQ7RiFVy9ASrwFl2OP833y+kywEUxTnJTmVj88u2cpO6yLyWaKC8i+wB
WmDrStzHIBUDQQo7NQLvC7TABhRyRcAweGHPV6ufnkC0VjzG0vD5EKCrpy05SXrs
sWWJCn+c+S8nsLdWMSh4TrgXI/u5V/oc1VdMFzHUmz6xO8Gy8taDec5VQVAE7s/2
v3w9nM5hRL/a/SBGsWqSK/9JG8t+ubdNVoN/v/6EArZuyylgaBaSNjG6ToFEB8PG
saKRxDnjr15XCmHNzlK9ItWqeWdLtXFZqPCpuBX73aNG/cgTZ0HUdpmDqmd2iYnr
jzQTwqcU+fefAnric+A8QeHAQP5QSncImGyDkFlnYh0HLmuBhHGfSRl/cv2gFP3y
P7YX57qcAToyz6F4sZ1kJe3GCgxvueZZ9sRMnrn0DHQqM70/eJ9uyDwJyPpx5LqZ
UpPrxwTNqaTYmdsShjOoejg7xqhSOMYAOtIL3E1milVflFU0rC1JvJ3PHLYdl8qI
H9VfatHF1maDUhshUIvMInsVfZ7L+0B89Ec1MceDixWxqIzxQGLQi7TCxh5pq6Tu
dwEgImZW2iGCk9A3EaJqRVbBXXj/JQ5ODNizD4Jje9hr8IFfctvh3v/33A4ToLud
Ob31wRktEjvBj6NUjMxC8mtAllXLaWXXJlhqCvMdZgzTIXG1yI0sZi0ZgtzGAhGt
ngfm5E09nrjDtwZgDW8kNy7Tb142prswr91f5a1cMYdf8Oj2w/M6zm5mwL/ztNy1
RJFUa3S8PRqWFxbkiJlSwXAd2GyrXySUwtUOIXS1cWsfDuC41m1KvGLXqlmQEh/w
NcKGx0lXcFUmxuPQhWHlZqUDVG+k9A2IqGmS/Sz7a47MY+zPFwQaZRsCrVcJFa/N
rDEDYdbEmtLH7qBnrPSJvz64ACdwX242tiYfTM8W7bXIf0OfjN8oWz3OxdwKYWsz
YRN6F2+OwrURIJPoHTcloCcAfSCpZuskI17DbvT1yHf1nwTqDg3odK5U/ASN2xVG
yvN2vfBHKj9Ml5Zw04KfoQjzikRKWwfHngO26HhGGfvbdSU/lFI3LLUD0W18AYX4
KzDC5vrXmG6rikU3YUQiETCPDZ5vZylx+5klMKM/zlfpQqeszpBuGVOSUbFfYbtk
hYdd8D00ET4m+lE8fVJamW9LNjnTK3hFSWtAYEXFTSAeSmRgGXf6aAm8170sD6M+
UP2+P5IUInja5NRSFHtDavplvkG30p5sYC6ot/5iiT0coPUZkGbVDIzC8zjcoQzU
2XistbZZ4iRpeDLMss6yE5DbBkm/N162Xvucjjltp0mqOYvmx6eDMFAOJbHunxY3
ACal38eekwdo1LlVvK5mOvCpf7uXc6nu1EbFvT48fm/3bxbgAfrJf1FSIPFhHZ4Y
PqyfvruXr5HHgx29zfmMEu85y1gEmOYQGiZopFSkLnMn/NIeuuPJ6CS9oY2onTIY
KKwzZy0FeVr37KI7fhApOO9shRVPceE8Sa4wwtTAj32Fx3aGQkTa2NuDjlNXHwjT
bUzIBsq6CyuQSQ8Wi8ZpgnOOTt0aJkh3qYMywPgSjIEHP/LpRtemgtcZM01tKbw2
fFix8u/fqLJoai3qP6yLywYFBp/7TmKeKSDaL8cLcysxvMCn3nnGXjeIskXxSJwm
FWwfpcHYy/+Rj0Hi8fARkCaAs2cNoA4t0V/QLD1zyyPV7jaqJ6ObXEDkG/PCiuIg
A7e4isdCyoZe9C6KmqUKGcGVZPurzEeba3vfykYCsxFRO1tqolpWJeu/qDbpHjIf
tkcj9AtGSTZw71GoI+mZV0HeWwdeHqBiXr2ZMmchCfOU/bVP+YS574d2vQdt+cWj
qAyOvrOoaygOLPZJL0R/KpJgtZ2gfQbbPhYiPA3U+/pnjb0oCNNkKmn36J6yZptd
24LP6/cU+en6NZfa8won5NPaqum96vSQC/Q58CSnkM88NGTaubp89cSi0kIKLl8h
+571q2TWEIdVnreALdum47x1OyABnDLjnR2H+94hVww3h7f1ph0pOYUkXT/3v5Uu
nsQLFWoJFM5yNVXe0ed4ki6iO87Kw8dTOR5mZZJ7gUEUg84h2EzcJvsWs46DyvBB
SPx8JGALrTpiDrorg64JmgEOhgLXo6+en9uRHn3JGD2mCcOHPEOqY05GLKzAYm08
cPEhGJBjCQ7EwbRdMXeuCkD/XGdIdR7AW4rgRnoz4YrrWSpRebL1Sp5lURvEcEe+
7fclmDNqdL7Vu48ee8HEGJeivTz9mx1E19IdU2yzwc5KyrGVFnH7d1L9xUmdhtH6
q7Zpq9mFyPe77wHId75WcDqpXVcI4NlP9b1wcZeBem9HP9YRPIpFmk1Lk10r5NW4
1yknCi4cg8lRIMsuNp5cp4udJEiffkTL3B4oRf12VQ8fHpUqdv906/1WkeecuTG3
1bz9MwflZAq7w1cLZDOgsWgiHrD/m/8qPhvNIqDr2WnTQzXJP/mcgenYPW6/7X0c
4dH3wqH01StScn3gkurF5nzRT19x4KyLUhKyZpbkuFSlgSSMJ2u+tlsjpQugTiew
b3r5bDfjTUwaSuenBI90lPU9h45MHDcKoKZy7HdmCBul2pXkGs/463PwiauLKjAW
cAxucblmPqRNnHIsH+O8SmURKtGZEN3YgS+NkveDmIM1x+QJH1eAkm2EKxI0EbdF
uLOxCAmjPHupPHCkTfuLUkFegqaR3ajTuy4Pko26HVG/KZ9Tsgl83dvfYrfYoaQS
yRz1c0fXjwNHZH27JxIUxXc9zg3zFVgZ2lysTND2nCzKpeDKHDdejvB9dW9OP8AJ
aMVPP9627J85MjCjElb55hpQ4ZbwG5k7pNNNCTY/jnQyp2GQLZgxgechQdQyHJF4
jK/iXWmikPNWDMfekbZ9YJ0Cncgq6LWi/m19WDeNCmdDhXOA6uW+mEbOwJG6mcX+
+Rv3SHExIyjRWpjTHv9O406fk8oj9GJSLY/KuOFNbqCCkpSDdixbb8bNAt+beMrD
qx5fAtUIVePOEEc1nccRE7Zf2mBEuChjdK2f/idzmMtLk8UUXVOZfzchlWXYzrnr
cc+GAXwsqhnHq+TC21awlx33HtTNHo6xZEo0PqK4o2qaJgntwdSZj+g6xtz4lEYT
dq76fsVJZUD2Na8uBuV48bHoCpQXzgpm7jAZOrfFGW1MCAIm148voHe420PuKj4h
QN009U6q/Dl6g1+p6cFBfzRNb9H8W9o0shH0XXD/rlG/gntc/UXGVWKg5pvNE6Hn
fn5jG6gnZwJ83Y1/9y4yY3UPxW3YwJZpeTBguYY5m05NAbISb/v+J525/yrUzT38
VKDwbDU5i3A0awhwI1vmHGCFcdr+GwUZrU/XiKFPLsZff4hhcl7BIQcIz/TIbQz9
h2i4jW1pglB7DI5SeHBVTejLVhVYVvbxwA3WGW8UtBErSwypMlOrLIvXu50UJ0fW
+51mKeldmRDLAzgbIGIP8nlc5a04Nh3czTAmM/D4FuTa8aH4D+3FdkSpe4AoCa/2
teNNVYscbTTxtgxgyDppCJngC92kxyD38gvyKManUOM/n+i2LTNuag9Q6Vfk+MWT
TIYh55XCKw80jyaVWcAvDeDDXLIgChtYTcgLsiyzHjkotZiQZuTV7ZX9K1w/MYW+
sv2UP5cLO9AEKvhRuoZIHf7KHzL0Ch+0e4NCSEiZQshF8ZjxPLPbdkUrbpVuIxo4
tqz3nfOaOeszDYl3pLGvBWz7a+dBWAGEOQx3SZJUqDvdCT3xq2ssQihJK6qKNWn9
erYI/0Rp43N+rVA4MPuAQ7qsgOHyfAnYry9H/WJJfRBfAis7jwtBgxbmM+rs+vnc
/SYEMYUkYbzXPWUe7lu48cXaEH8Bm14Vh7YulHbnef6Xhq75CDXNJRf2He+cdSgk
K5GEuuTN45OKHjG0w2LhjX+pEoOS+vav8W+5YCpLOOMNjx8Vl06Oyrj/p73lp2+t
3XPH8Xr8uMxKpxBXuYPKPBKZAnmdrmhDLF87+GuoP+fR/bhvSjUc1oMPooScRC43
NXev5+FRoWD/hefZ807xRjGDbZJyseun/39Fqko37PHe0s/tZvkLUQXXCe2Hdc/a
SgVPYvfRj0eBNoKXTEDyEEb+Siz8eQ8iQ6EpJHKDWfGP5MVCHGw/9bsRlRVm58qw
7kCraTBJWvVKGarwNPxpG4naN9KGhpBrqSf+O6cHqxpXzcD9kZTv7So5x0qstsgJ
4wGXszwLRjm1PJ7PQbQGPtZtlY+MRMynjZhO5wJSdUvQkXxCA9lQqv06EiZJtsAd
9bxlacqCWTiU2Ho5rBhnwOKAcLzb5dw2dIEmeVLgTNZdQhrgZBTjD3QbByKbyDQs
NtKSECUXu7bQtJlG09EDnpm6F1c2/Sy5UptxqkJ6Zx4zP3jIgm2x+chg2HYLtjzv
rsXYsZpStKknnfxF8aeVoewEuoZqK15WQDixO/ofBUoyGhhitSlajJ5fzE89tvGz
ucluVO4/Pdv/WpIVK61PWToHBjaRWVqx/pXcjxUnxEl7YlpLRZgsTYBlDN2wodNJ
ZC0n75aIwSziaP8/WmOdZDKDByl2kKdFmVqzkkY7gbI086PxIexxWA2oQwLLTelr
9gZfdQNEoMZiKwXny+oDo5veyNbstZ1lhXle+2P7kaq37km6oYaAhJrG/JqvZSnx
JhB9ikHzYTDJA8vE9w+RUatGhiZsAUCx519yc8boXBfA95Y4/nvnRSY+jguRHVSK
53QOT9oJeTsXaMOYPDeeIYMf5BOnmwafZ3vjE2ndqvcf8uaMSpZ1GOZCdAFOU9vt
G9iYcIUBbf7yqKxYR4v2Pmrr3RPuIuH3U5li2ezl/nVPvpIEdlZzYYOBLrddKY6I
HmyPcQhuVrpFn4jdVMsvFwRoFd9IKo0jlHetEe9VjgCralkQ/Ce+tZQ9M+Hd/kyy
T7xED9uTUlvld/k42qcmThq0snKHBHF1Mfz2xOfZxUS9R7KdWPGj4QpkkcMwvvYx
NKpEb9iPYfD9Bqa3lF3Jxq+62GwQwQ+lCGd9EsxnloizoA8OaOihbuYg+XhtbhWh
3d68hfhqV0MNh3i+wf0KF6MFkdHQHfQ/PaB3F/QaJ8mTVSBETASWe5t8OloSDfzu
jFClNKt+b5tY7Sv1B4DuAFPYAA8pnptVSYehApt+FYNhqTiuSXK/iuZubdMdDfrD
WLcV3kDIR/00pl4/Ow+Eu3tA8qU5CkkRQw+1R0qQZWX4bPKbAyF8r+6RCidHnAGw
mGZNcs9YvRThBrWegiPK+Tx8iwEpcMMdiFc3zu7DJcDZ7OzuYLen7FvbevkhwAB6
1b+aLaothR6U/rIqtGOBF/YOlO72x1w1227e/qmezFIHcOWmzgHPOPFcqwyIDY4P
YxmH5EYds38dkq7+PWdF/uFwrvtqY3wnmpHuary99OrQzBYXzZHueI8dyfhvlNVi
Orns6XFFkgBXYjypfwzPNTyg601ZBIif13f4Y2S6CM4SxjVMbd0oisCtc1JaW3Ri
HZreUkgm4T/MzKzMS0yW9kySQiIEmpHMgDSVVihrpojHhfZ42DFS7Ne7Ggm8VIkH
wwX6AISvPPoSLmT9H08NGVbacXnVXmpVJBm+VYDEkAx4Z8t8L8h2SByv2LZPJjvo
Pxo2GDIm8B7yWSVpho8OkQ034uwmxHZrOZ0fH2eOK3nH5Femt0AXNblAi1FnS53R
qXrKMoTiGihGRBrBM6TnEwu9kGXPYouVwfJD+2PV23AxwFkHTB8+O231Cyo02egU
gqvusC3uTMHjffddy0AJBy+8uwOWc16Lj2cS5Eo3eELQvsaZox5wSmxwyVDm1prM
F6Tt2Apz3tROQHkTJY4CTrqqxhNhJIG9DD5nRPexhpB7/RokpPWBK1USJ/gOW7EZ
Wc/J4cdI+lYl2WOox6BGIf560LYEOjjUnkJQFCh+lm2GwNqvEBFrsg9S4gfPE83/
7EUA7rKcaeU/b3vWv9xWNf2TrVk8x8FXlPXUQI6CUSXqwSoQG2cMo6HX+yErAKPm
3GhTg2F1ZFfx2duUU3gqDrGLLzCLvzWm/sCdZbmlYbS+6NbNS5mhiMCp9sI/QEbu
e39zDl/6EeYilE2v0tNnytns7Xdf3P6yGdnHmXowZpG5R1F3KstZVsSVMXZ3ljbe
Y81MpKzHqET32+Qml/8ftUDf9gbhAXFA1BMl7yne8gF6e/8T6AZX/hwD8IQJc9li
rpbzCJPwdvep0WxcT1SqOUBTuVGekISkW4uNbm1mX3TnZnfhiCmy53sknizmqKTz
3rJQr0mAOgKNEwcGmf7I51QSRSkbx+4ZH7WjXV6KnG3ThrkY09Zy8D3eQQZIGEgF
xz6X8AC13KHbTfkVEhFc3K269JfRKj7YK8KgENK95WzIoG8FWM9lbOjUDLpJMPxH
+UGGMcozcV5mwePbJfaXxvP6cec/fMApDnTrsN4A8YYVKgRGs7T179kq3cruSpsu
YvRccUXjVzg3grN6HmyqltQMDHK/hFHOySsC32sg4N3wkG5JIZTvm6ipgJ8id7u/
H6P5Ej6wPWF7jri5Bh3RCbgNe+GVxVw3pX+Hu0rpA5kVxGPs3vaSDfUM24f4RzR1
Emae66+8iK9ekTp/6zIiNnaki7oxi9uR9VEvIB0wKHslG3RWu3Hv0wseXBGBsSjP
BxbRjYTZucpKf5J/l7VYAzZKVuiilKiOeCBHmKWJBVr2SqkgG/j9pQZ8bkTOZ+Gd
jiPS0SnEvwJ6VAVTibphopZSlfEOdhvxVq8ROpQ9Ga2MDFXtDnZxffnWrtoL50s9
NigtxH3MRNyQGZQjB4/CJskv6k0X+ITnfj50zKNgT4Hkjyvr+aKRP8e+MjMCQwbS
6H8BSxdCjmCW1C33UtZuuuZXFbDLhFOhiZhkee+BveGK0JFyeycGivCYFYQZZzL0
3bu6droQJ+J9+BY8os7W7n+j4SEg+RwQiXA38LVbTHqs5jJ2dgrgROgbSK++YPeN
fpgNLbY0RoCmzvQOFP+XsJokOaIGgoeA5CqGw0MZsXKg8rr7pWPj7BD34nLsQSHz
waC+GGXggKFTrjCsAfh2yqrZY3GfOgusGi91BT7TRGA9yx0xW5poxk8VwE+xcBaP
uj9fOYOjsQOE7jSS9YZbv+PV7QjhQo5GeX/KelMba5h0oDqv5qsj3qEbMNbD8Dko
WUWrJ/6GVG7wrN9AuC8Yv2pV2hp3BLQlI3C2086/HUBLc4MNTGoTUlLM/5usKQ3w
M5ly9pa7hXJiXpLU59E75nMEq/WWCB8AMO9vHLgXdXSQUWFuovDpisify1doMUK4
+KvZcGWNueP2w5+6P/BFuRlMdJog3CqxsHXNsalgIwkrPiLegUaAn5Ae+Ys2rOJJ
OnEMP/PYpQUH+mNyqo9utp0ooBQhfM6RiTM6hCYkkbIsmLS3Ds11VDaMI99Z3Nkj
/opj6eQEcN1xUWC0DvCX1GZyhCiosDFfS5vCqScB3HobfX9OQPkRIP6xGavrQrBm
n6Rh3s1jaHgqUZKk0sihGv10KJ9xl313dYbdPnxa5lALrgzVAyV80Lws5QWXWXx3
S+qZEXnstjr7sz8bKZPb2KOAkw1RKLKp7qZ0dDpbs0AHwIBwKI3C/EutdQK7fU4J
yVj+HSpK5znhOzviC3crFc3A22qfX183mCgrZ/UrWtkrJVVXDYqVR1cfNTT4BLHE
Nlxl2J6OqlM/J/0S0U0vwuNl5nUqE77xBQrtBe/pEUCshx2P3GQBcsrgsSJSv8TP
Z6nJbn1+eVsOHHNe9dO565MuSbJApYJf8tk19ugA5Kuhkay3osAUnOjkF+ijYTJI
kkYo70xgbj47NTpByA/WHrWNvE+iBYdM0ht+RfMZGqubZQ1B+lm/7JHa5lwhIri3
VjZ4iwg0liBGRpESF5ky4OuguJH5RDiSbCe/HVlryquy5Lsx/JFcyJxGPhaogmXA
4jYj2yx0wNHUlK5NftU74CW2pgY5WPeP0tHZ3TfEukeUgYbvWEODeAXLM6MTkKFo
M/T9N5/KKx+oZNc2yjR0JeeXKcf3cFwTtSraUAyarYMNDOFejC7SXIrmLqZMsRlV
OD4dbwwd/BqiwlQ7cXuGnBrIF4sTWBsEGx8U/samYH+L0OuvltDVhLvEDbADpLrO
43EE18zzCPqUj+Hb/h3cq/jfSbWRjAp/Px6tq6BBZxl1mf81VXxhTlaAV97ZHD2x
YX9LJKChPEGYNn+m09v/UEWPkmZj5WxVDDs1Mn+sqKKJU0Fr2BGditiMC5UA4tHv
DQD1vD64zuIYD+P5XL7NQMFsk6SvYlPWcofWNv8S86b9enGEhyYoiaDdGTyj5uZg
v2BCs6tv/Kukb0VRPSRPPwM4vmCPmuXxba0fUCH7sIoRXO+giSoW3Bl+VPVWnr2B
dPuJhQSTtLiPqw8gvQJv8uZhocit3vvktxSTWfyM6Dvv5b53VOJ28R1zxlt5MFjG
7dQEtE4b1SZWlbIi/Eg5YVGUf784GV9UguYDZGGdVN4Ba/SbxXMeHZkk71Z076zn
GP4CAwUrBvhkudO07c9WAnaiuRtNpVY2O7lsPMH4J9T4emXSTLtsqNg6/GX0eec5
ll0LdGXBCwOt1CDB9GSc/fAe0xy7goZ3fVWdENaRu7ZhPewZD+Pv9JOv8QEvD4Sh
w5c6AMAx+fbF5tjT5VfWooROfPJZP4WoYu6YnNK/rhqd3vWr0RUC7SXV1w082wlP
bQHefpqSIj9SBaejcTch5SG8GJLES/HVW2+/fHh6Jr7/nDFHOE6Cnubu73boiL4E

//pragma protect end_data_block
//pragma protect digest_block
hT1QKZoYW1YtC0/qCvCszR0FrXA=
//pragma protect end_digest_block
//pragma protect end_protected
