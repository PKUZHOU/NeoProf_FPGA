// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WRMywm1pC6a79ARd37FIYnjPHUD06qFu+xCyZ1o9fJMPV53+cd+seWFPow5y
Yj7aRA6GDhH+YJSSywOLhBAOqmRPzTG9jKHxUuZVQIJC98HPHOfPgblYbJd+
8scSh37iP3Hbf3ecYLfOYoPu8VDPmG/ALmqdGrEZEvZXzleEEpKqDHPOIecB
nMJ+LH3XGsm5e5piaHV7rt81QZ3Xo7duNgHbi0Wq0DVjjGg4RCIALcKfmZaZ
9JfzQI6Tz6fdoWgcI/VxpaQINCyKYWuA+HJRVjgA6DkQUaQPfIKFisIqsSIy
5WWkdp2H7aynDL5NQChfhBmcXx8D5KhX+3OEU4g6vA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n2FuUcNYZFH7OzGu/YOH7uRe5z8isvZZPFP3AOmJk2rEaHsE/YWH3bsB67lX
3jlNiKi+Yas/KYOcXfT6Uc3qsW1dbfDQkWkC0yBgIRPS8BJpB/u9VODuz5x9
V0AKpQInCDFu60KumJ1ZjsqnyYm/Nlh9bpphaKkK06XGNR9iNgXf1tj9ct3f
JYVNjvQq7P51/FuUX7mSZBGdRrOGHUVxiDc8L85GXimug0tmRWI8JbKrB14w
wmcXJRQ/iXv2VHLmgCV74Yz9mJ78YOjG/F65T3/7slyS51YU4ETrYEemxE4L
MeK38Sq86rOc6r+CQ5fwUywnNYz9JzQIQ5e7sTpIjg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ETBeUPJ1iLBd8FJK1ULQEm/ro7jRtcdwF48lC8ckiHHPiEYeo1FaMB9zGtJq
k+axCxDPd5SGpIe76gc9+C9juuNh744eiADOdAgczoH7Wd3zSbqbDPb4xMV+
tv814LQLHVaE52UVRL1Owc2aSjKU+jOySSczTTLMLI+msoA59WJOTHsEkifX
aB7aZclD5BQRFjYmsTi/qL/+zYRuiRucnhT2hsjR775KOoZxP4AUF0BWCtCE
79PT9OjrzLwMF4PClk8jXYlhACaPrZBu04Of2IjnIemv8ZzZFWxGV0jPCDMn
kJsnjG/LFn6yEmxV2uaLKkDJ3r37sXcBLXemJ6YRtw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bjA9HqtX+wCbKkBN4OlqUQekVkOIdk/RYvhZ5GSzr2RdQaTKOvjfay4fGNFF
C47Xji1hBN4YRCC9Pf02oN6UCFgQX1+hGMUdn4ivaZ+sLJqCN3EPkMMQPDnD
v67yq966K1Hm1hHN1ekZo/kXklazHvF7WAGbw05aoeNOsp/c1y8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LaSMwIikvRy2MzwvSsd1jSCe4VASrzyhYbDQl4d9v73BU/v7lXOwWNcJqlBU
GrX9mSVYI32CCORq+0M/j3qW/bIQTlqjnd6b8/RjJiAt525aX/FtHmXRT5Nm
EtUocSllJNpa2NxR36GR3YAGvaS0LYUU1ZHNMDdogUIHx6clI18jbKz5R/Oh
AuMRSovXbPOBhJ4X4PczXzWyVz+SrYc9fwpMdgdnhpc8i87/rT/k86c3HWgZ
w7rAcr43wjtqwB7u9CrMuAKWclSiKseUHgP5gfIf7tNYndQd6ZnasVuarmir
62rhYwM7MFWX0OPMkmKLSZMKrsU7kVo1W5Lff9xWeWgjvYQd/Gj47+yqmTZh
ZkxwT2iIo+RH2H90bWY0LTZ/+4QnHu0oINUryPcvdAks7u03CRegxrCdOPwK
PxEvrrvHMBUa751Fv4x/xiMjQnaqqKY0uWoclFIJUyPXT6gmNx49dPGnb0tX
MTtwEmoo9SeDt7CGQmnsEf+XKTi9TubP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
TjMBRvlGFIcU7QXeYnf+miE+pq53eO3N+UT45RL7fMcUPwA8Z6TqhpD1KKCs
CpNw9GYn1ta8yhdfhINhVZ8FvwJEUZN5Dp7/xZ11dIZ/DqqvoGZ/TfsbrK+n
zzUr60xpSqpD8SbZrf+BSr/OloDQUO0NQF8reS6C0HVNXyOqFRA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tzdLnGzwtxwgPRwa26yhSDfx0OrIQIYoc/6nPM9HXurhIRlydxCdcrVVLZ6h
XwsYbSPM2m2KsDtdEaWMMPqa2YsAARhiG9yeJshhjqdDjihUw/4cS0zPjZeH
O4CWqFdR9C9yKlLke0jfCchX6ktK65IJeMzEFFIhFcZ1yur/jHc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10608)
`pragma protect data_block
tQ/fTuu/zYLTCW1tUHGyB+t1GHq1FmnpXSzBCq1rxCPvnLriXpGgHp5Mrvl/
z3zX9/T/m651n55jqm5LwX9prqdz9qDYl6XUs33kkUiPVfqSys7qZpgSg0/D
thry+7VswcJ1yI5u3fnru1V554Q+oihqlIv576zFwb1RF108jR7Nk49AcMtS
2xF9+r4T06lP55/3oDT6MBwWveqcOkGYAQ+sYGHIvoobtqjM1kiMzldlxluP
lF3Ws4LZRpSqtUdvHtW9dPscmg0WhBnO5QqYfjh6dfWuLPVgznH+MxYo7Tqj
7RFglxSgqOoUq2T8qGUKD2+HQL4VZI8hepMfqLazjax3KgvJQZZw84ZFB+vj
hoTIFANI7WRsvqSymFyGUgSGeZ2AGYsfDUXSs4ex+HAkU9RLMMPzom8wucyj
AlKZIqU1yyt5AR3uVxKtKX0dC91mlMwpoWrPdXh46zjvEK2Ivm8FFaR9wFjD
qh4X4SAoNd5LNYaFarJJ93Ak21Br1Vqq4NSVYLm7Cy7XBrl4KxamMCAdWuMN
GTtichfIerbCwcseEYve5YmUgPc0NZPjjE1rqOfMh88ZUy6PXZA7mVMFZ9ne
NUa0DZWeBOTcI8HPs72D+roz6bu6ZhhP0h9TkWuRu7YOYt+Axyj5KwH2bPI0
3QGxZ6dtz9zITXG+RxrCZrt1+YK0Bnnd5N4imY2GqZJ/l1mbckmn46YRB2HG
At4BYWE9UDc14eyVu9a0VEKy0dN1BDMMLHRlOrknlmqsCGUfeJcAtkwu4tCH
B4ZL98TfCNuCuJN32rOquXG5hdquYoN7PxEh/UwO+FNcRVhKr9UZrZTKFoZ3
HPaFNiZmpm0Vpv1r4VVJQwXUCZ6F1jKalM3t6fD9zEBmHccdyK8HWiAEvMTj
D4GFnC0t7ZfBAbhT2nApoqmFWJALV0p4QDcg8diKijRySpC/BlTNv91RCU6y
6aPSlvd2+R7QE6YDYXBJOVaD72oy81tJH52ck+DiM6uHqCPpnD5L6svmy06U
wnV4lnWakpxw0ayVMvoTI7GjN6bil/nrSKW9TGRcncBS8Sfh3aOKATy17NZL
8Kz2YAPQWlHC1kGgqWCF6fBVUGvFNsw3ufNgDkG3tMIndK3EI2BX9bFZPzSz
zgz9GzYG3DCshmdao8DHThPkbY9dB7nKDvoXCu9PA3eH27Er6PYtFh7SlUMg
ZfzSD43GGgSoKjkDR/2KREC7BfsBXhucqgzXP2pxzLo/hYOq1U9hS7jHMnID
X/ix7x0xMI/DvhNLyqDeVoemIL2ysMB8NmZ32+8MdT6ZeeQovdjJ+m7zGm8D
b9kvg7/Q+NLlYS6REoPhRL2ry4SET4PqVmBNeAnpZhbe1dkEV3Bk2Z+GY1Xz
vR9nGXSu/qgkNlaAsmxP14lH/W0IzzikiAXv45eEb+lwIcmZ9t2QAKw72OMe
9FoFHJkyhnjl3BA8+eJSYswX0ynlUWGgiKScR2EssPY/u3WZQjz33gK25kAc
MRWD2KXKSsuShikGCP8zKvxcVISVEAdsbXRXfJKhz7R5a2GxAH4UQWI3jIqM
nKL407ZcNurVo5CGI96Q1LsEGUNn6Q/hXKo/eBSh1OMJbcxhKemEvDlL8Kvu
ssNNLjLa1iLXKcN1ALzjphwF0eNY5B8lfDZCU+tAd47xAQSLiqF4U12RkiPu
KT3WtWf880y7NYRE/XsXO042ICtQnY1gNBW5EL74G/b8wt6fW+VNm1L/Soey
T2/govpl5ExSrPsuQV7GJt3PkfuDCR5PWUA8e2IkdlKelN27wgXQCs/XELby
KSjFOi1cnW+Cw72MRk33jqzVXuBN0us4KHQGwqZ/8zp0k7tXPOtiLSf0hzBP
ZWpPLtv1GqVqGxYP7ih7TPRul0jAV+QZfXT25yy4hV8CRr/JZi1e+Wyo5caO
f3NHeP/CsmjzEWBjCIKsFanneCdnjjyOyHblDA9cH3lm1cvEB4aguek/IKTW
+HELqKY+00S0GPKkT2bRAMMYT8HglVO0ZbL2OFi8+H2NTKhww6Kd3T3Jyuqj
OY13N1G170+9P0cFp+SCVz6QiD+FWw+gvqYxU8FoZZePkA9H24YqIaBHV84c
n3yMT/UkH5w6I8GE6bh53yMetSj38sudRnzAmxYw64kLc7HY1BzskEaiFOEl
9LMNBWbwDnHaMvPWaEunXz2AtX3HijEA2txHfK8bHQRea0IQkhgsGYtAvbk1
FeuO7xGeR36F6otTqwVEioi6aPCXnhAD7yxnwTctDYw6R78ccIvlSkDkFFhw
MkLbx5bVcOFGYSkAFlMziCOa42uzuOwkaK9NNWuNSiAOV7XY1rw4rc2L6EBd
6dg2SYBGPnK1ZVB7JFXQHqB8SfAU3q7a574Gy/YnA6bkvmLVPB6GIcfd8yww
dZtqtWri639U2A4hPeCnI0CXX/Ae/+BT4uIqaBR2EPvbs2GSgNo4ueuvO+Vp
O0V/r9OyDALCorDJJ+5Z2uDZyiu6DhdRORw6SYDogpgUyiXNYy74eKEjeVY5
CcKwS/WP+qlj+ZiNmefoT+iKoI1l48aOcwqKfTyKBU5CyJzOgp3Moy7noyq1
AxjMtn+G3Ot8IWcNwEclKiu5R4K5y1378ADo0n/I9N885uE6vypWVg2tjW4L
E9XvmEsrkbiNls2TUppf7YeCVrynwmmD0Ml54NF2cT9s3p7e7DP9pvmN6tKf
d77GQfDgUBigGuu8YAces4YFC+K91UQKYa0a8OY74X6RBEIUEV4EzOqKAC//
WwcLrhm2/c3GmsJiUDI/Kp3F/z9zruwm3fIjwfS/JJSadFeX5sUB32qUulCe
OliJH6CkAAfHfSeFjPwoWUQjThxCUwf/V39BLiG9L1c/CbspVq8CnbHBkiOx
MTh5wlXPdg+bLaSIfl4n+jK9OfBhyLxvD6sb0u/LsmngH1LGzbS21vWocUuZ
FuYk54HH95KlqtUABeQny8fa/UmaLb7WYaoERKDzmrpXDCcnLgM/0M40I5t9
/shhbXxLTZMYQnK3B5QqAddK1/T8gLfavIfzcyONl5EtgF9jrfyagXKzB+f0
foLXRwfGpYXZJogLM5NcH1QWsYOF37NsZRv87n3xiAmuXfC1bpMREnwuOHcp
QPmkFp7XCUb8A8pFMTkyt7EfzdXENt/dLct1kC+/lWaVDeQJ+jD+QC2SBP1D
80tOSDqbs7la1/eP2YPpYui5e5kw6twJPh2arydie8Ga64I9hhC1kT5fj4lg
Io34Cj9hRZ0XjUWtaxKR2HWA1iDouCYv6kf3TJMkVECJZTep/uRAzsJjanIW
+JMIyYH6ByNwIHBImZQFg6Aolm7dkK3kNmHyZN4OEA10hy2U2x2aWyS+RSQ7
4YnBF2GAWpuolICDxIMZEx69WowBTx3T6Co47Q0vQZcB3oGArIT2MKyW4erT
kk/zuz+dncU2R1mv9CO8XcL4RgsUXrv7m72+BcGXA7c0ZFdd4ekyHCc4TZDl
Jhcld2tGGUbV+QMorApbjuIrx8a7Suk/ZE21aCteRXuAQ0byi5HGwV78XyUm
yfeT56OKAydUdeqc2tL6m846B26UHM02uFCMws/YW1aqrTUJicjkerrmj5Nx
kx3diJIkRKA1kX3sncf9sdE2X1BHcqwRt/ZviPnRakhzD1n4rrHueK+ILTz6
H2Tk4R1ar1/ILf/VEVEGNlCEScU0JtkHadZgC8AOl8ivpJpREHC61uivXwxV
jNNLvn0iKLuSQd4YP0ImpqyBdakexVDNt4r9YFNXua/7gVRJz2CG9WW9Tp1M
9tUFo8sBq5+bsxtsXFFKzAYbBLFVmw6su5do3gRft8OFUHAIPM5JPYrLCxaD
+q/5S8yP4kvqWxEYagzMftpvyV6KBofHxBwhdEVPL7XrItKgIh5v1/eDuI0R
SnC5Vw+guGFNSqNsVxvKkFe9DoQWQnFL/ZdPqxGmnZLbcYTaAtvsZzz+UXta
pc1erFF+A+2wwws+OUrRl+4cZfQKjudYu6njRH/7VgOND4MjnhiIFKhjPIIx
jOrxN6bYctJDkBpauaM8B5UdupobQlgMoyFEXH2oLob13QA9eBbFgMc42Nc2
jo9Z2ZHfwzZ6FfcN9JEz1ti6o6x+d3CwrTGxLbshWpaoUPtoDTtV4m36CpgG
a96ghbC4BOvj1ysfI3pfo2dKHwIn2L7hFWs+Tbprra+tSBYr3eZgz5G8J80h
ZkC2Uk39KmMnEcag0ZGETsHPv7l5QnLlgphYE1F7a5B/cHqBMFqxM3xl37eq
uHnWFfIAeyK8PxoYHOphg7qAroKkFzNq3qGNN97md/shst3jlw2T+Oik2E/K
0BMLV/iLMuJNFnzvZgTDzPYjdwjsLKOz+UAU9xrTu69x7BtC2TOR4FqtklL+
Kzh0NoWuKsHjquxtZVcyDELEbqCe09TvRDRAvUxEMhAtpDqeJPsX9jXsyeUr
tt7Yv2nx6n9FYAs27EbNYy6/e/g3juHdFF3VOp11hD32vlcwu6vMUBlxQBgr
IKQlOyEA81Lv0UAUKbTDjmLr6qPkTTpvCUZDm446gzlnxwi/3I2gSgz5q2aF
ww6Q9P6KhT8JNqNaBKMjqDOfOgKOFD5VfZtLfkH54ySOi19v7v7K83TRXiMe
wfhgISBgDbLahpW1LUKXOVFowMSHzF7DHr199rJNEsKvtS0Cmjs+wA5RnKlJ
5sbhUGybFvv18njRLGp8GMbWbl/5ZSj2CUlCB05h+hcKqkM523reLcnLx4km
3Fb5vuIayNdWTfVTv/gtgc4SIGbmuszNbRiidxZUA3NEVV2VDijJGODY0DAr
iXHpYq4e4igVEtiLpt3UonHzeDzoyt2AZe7367StpY9Pm4ouB9WdZMy7IlXF
tUdOJBmPag7AfMQN8IkkACtYw5f531wrbrVgn+aMMKVNZl4/9snrw20sUUlP
rB/Mso3CcsOBEfNGTvNr8LWer7q1UZBagYPvfZT3kHQRKfssNSGUZTg2KLDz
dZAv3tLFVNaE4NcNMx2r+ByHbf93TcAMBalQ9kQJ5ENBJptL9uNWUGO+ZR9H
/uW33RUluYCRu49a6fiwHib4H7OhNA7OQyv0zSAb0ZWPt7pxlPfadvR3e++j
mCNlycYIjduvpuGTjma6vMis2lFcanJYn2SShSnCg27YeYRBeCfS7G0qPtWQ
ag97Zy4fOYtzU1B4qUS9+mlDbMqjAfSKiPMZPB0aojfOcS0DVsOHJNUwE+Rd
ugDYYnyqIM1tt4v72ADQ94K5zv9OilQa45nXwQArxCYaD5UIH9KYOIOR+9yE
XqH7A/bp9EvYsHSjkIizv+MlWGuR8gwb3rWm5sOgVNRqVBsau2Z++9449neX
0+fs4xESym7zJ3NB5VTb/U+5CjS7W12UxNKnTc0dkyrkFoY7vdZaERgzlHYf
9eYqRmd1fKkTBvxDAEBS+6ETZVYZ1OoZ2AEjE14SpEoNvgqtl8avm14mtO5T
6ePQPBQliK8WrW5BQn623WLEDpbbS+kvatVDQkql3XEpW4cvB05+UCeExZxg
P6YQGcUAhYcp7Nrr99T1FwhiF/IupSS68Ue/E/MWTtmDMkkqrH5BL94zdWs7
Lsx62CgPe61yDUiuq5Bd786fsMVWFj21Iy2pnMpUd3hLnoBgYZKaItYRek+w
ARFoK4pEtIilkSHIl9GIUqHwNCReWg8Prk4c2UKoXYbIJBE/vKDcBJWmXmPX
mmrbLZGtF8mnMSQdofdFQaFutX+OBEu05iS7hs2cq3j6LvRuHu8oX0NbebXd
yp/RulzAf1+kDeKI8kJzT+KmXaWHl1SdrZQNIjtMmFAplcwBmvIn6qP1d+sR
YU5RNI8O+pxvTzqL4Qsbpw6xfmTvSCYVoA5IAO1bgYvb1eFLah7pu9sEtpRQ
BGgdjFJZN5xxP8Xt3sEu0rE+Yt9ElTZpfIAawHUPwZ1OzRtAnk3ID403xd0T
OazR9HV1UD4Gxqpl1IUFxrj0aIvyn25/qd+kJwmHtN7DQjCAnnrV10a6onI4
TFpZWcD5HGILElVqjWOKsTtvRG4ShFs86kpscdBoD+eG3FX8yQqAwxxyKL2Y
Ol2mqMhmAZb5Y2zLl3EPMlVzrkP0VvX+WkoniC50w9BZ2YCoVWXT4JxdY49a
XG3UBKYlbLxKsdM3grLMtGwBsbu+87ZbpDbpAIo7cRSQ6BpF8BjW4DtAxJe6
Nup6jbIVg8kTXkcGPnP9J+KvAXlv6YLDurgGHyTaR7R1QeTjaARBY0Acpame
5Q8OiYyzXh6QQrRT8xHOCmCFs2E31y321Q8wEDa6IvI727yZLlksPxVet9YE
2PWfmBkSbZhXf7nm+g3SaQPLzO9XHzUjVzi9O2gshnxsDzlyNI+lXU4mtUYF
novSdqbvWUXMvPsccCqFRI2S/Ujy98GKOvJtrVrK79ZzYyPizFWrRMpfPxaL
wyEPscgNVezJWCrCE7tQ3Qr4W0VM4BY9JbG1P67ftdpBV/ZJgjuPjbYdu0Cy
9vfzoO2iMdw2n+83XQOPtARIMJBauZT2xZ4kvKUs93DlcRY2r179RUhR6Kxd
5oy8GqqAprIwOhowcS5OT5WBkbhilXS+YY1g866a/3ilYGoR/cy0+vmrDaFN
TnJHqWaCxVnMtXHP+jsvKFgdiHLtMytsB9XNGQm4JRRzsKmsx6FzdEsFUZy5
w9HUkGAP7Qz3DZ9CL6TcLyP7S0MFZxKzM4kR1uIswNzsnDexIkx8O5LguKf3
7EgnVeZ+VWEqu70g9Yu7L1BlniRPHZ7PahVtG2b6Iu9bsCsG5fbZbvtofA2Y
0hLJser3C/r/lOeZwkeBr2nYkb5dEgoqjWOO+4gBCt2zFigr5g1tAHv05/Qr
0KAlka7fNNvtTxPK4p4I2qnOlVTlauikATa+aXRjNceVidXpqn5mOUAooqM6
UploWwQK5jo0Xccx4+qvsLKz2JxlY4jHS1dvg930srKjYFk5ASxLcQ9PUx6m
9iTWA1gnlOUW01sKie80ucauca4E4ID3NjuAf5Rh469+tQg3fWR4pqZfXyYB
bn0iH1UiO7WGfXMRho1T7pXtf35qKA2qV3cdTq0htgsuMb7OTPf6t7avwaFk
VCpOvAvc7uuVPb+5gpOQg2Um5Ox+Gjg3vUxrtw0erL2Xyuy+dMBaQwY3iV0T
5NqBoOajISD1EAPjHsPc360/uuLaS9oWBpKdZUciJo/E83awsHYs1tbDDDzV
yytKGNV75TOOOOjRuPXbfp8UwcTDhsJ5V3yiVH5pwM8yPNuAv3RMzCykxYip
B8OD8Xw9U4YIlMNT0qjduXCk6wEXBhUP8FQvx1hscNEotR/cW+DV4HnfAjUO
I1nKwVb7qvQrc5Win/e1NgE/pCRv2ni65SUYlUsWsapN4kB42gWVmARs0716
DGORWSkkwMdhZIxrf8m9cGNYypUug/5/Di92Gufo2a+jAOoLG8WM73b3M0d4
tkmncBfPidTLJR861czBTyoQHQdbWN4+4eDHHq6RJeD0qwMIm0lscklgDBWr
1FdF9Lw5BD89P0VGIcLRaWumu9JAq7gI3gA8/fMNIzOAgU61dRKo2TdBpxvZ
Ch8FvxAtTab7BGjNi24p0C/QwJlGZQXkKfsDg0VbM0IZDW38haJDMu1RpIXs
P5MCCs/hKKchPJ8IwOcyYy2S82N3kDT9+JOxlCv1XqoZuHu0ArhcUH0kWmuN
ToYT6HOl/jZJusXHOmTrtynlnY7nYuR7+8laVxfGx8C6WDhXfduVB139aVRP
JY1j1OHm4nJ5k0tm7XQ8jstj0xZDCMIatnCFNl9zO8o+VTyG0ELcfyJsdoyU
jhLBTf0qJ3pRkG1o40TynWzrYmP9WmkBa8CWZ74g7D/QvKupqkockmQGbIA+
yka/MxR8C3/m9su3mhDHapXMlfx7J6g1KLQK74XEhWqo84N67rQ2+y0jCsOA
Sgr3hi3sSJkxoktVJa0APbeCGi50xhlPyb6gaC3UmkktrAd0lZ+VEneu69G+
i+287zT5Y4GVgdMeEOD3bZn8YT2ov6BndW9KAKBFEf0h9XroVdGO3Qxgh5qX
3P0Sz+urs/GhdPN9Zfj1k8FIrjI//wvm75WfyKMTeFh3odyWFyR0RVKuY5Jy
twdYgZwUimmzGN7I5I3JnZalr1U3F6r25q9w5R3S47c7eMzOGL7nM7VJM1nG
gB+zEsavGKLe4e3I1vz9VjyjOQmNIjYyQvJTnrCpoh1F1VHEH0h04MXvPjoM
ZzBmwabNWkgwX54YSfs6EEjFxJyrMDWiBuzc6xLD7nO6ktDFeafWopj03+AE
MjLM2rdSNTKITwFwZyGtJq8c5EVic1EhsHZReh1P4CGIJ+JXDMSMdBWd6QOn
HFu5+WwgXfLGehHtOjignMqjoLwdNQRHUCclXvrL6yxXAOft+jgxbcaQeNLQ
r4w2mrMPtpKbZhQqU1qyaxVSGbGDpxCbp7cJzC67j8uVmXBDdHmqiQp7JYUP
zRkZwx9fa3X6varYAkxHGPQ8UEBjNW3Crh34Y6bKaL6meySnIk3GJFpfDv+W
2ZRJfFdzO1v1OMwForJuShEVT63rfYz3NpsPJIWC+q9JDsYxY+/2M5e1QBZN
H7G2wwf2ePk+Ie97CMCeLhMPUHfj4maA8sw45bU2jyMGwFYJq+SzKo9a9W7A
VH/wIEvHeXgDf3duC/j+lo82oM8WMdL6UTWxTqW+Pb0FoKrFxIk27AcdEDAH
Ufr//6aKRZa44NJvzv++BX0/HGG9VzeF8ylaku/mTh2nK1pkvy8ZxvuvuC2b
gSLK17N1N31/fM7ipmHlupDcABAN8eqQ/nL+ryCYcMFfirI/IwkAHinCfmJi
38nkCMuRKnyZ3hSbAFWppWOQjjjtks+yF3OtpgVpypL7N10Q9OMlXFGzy+vp
hK8J2QCiqlOdomnQY48/LtrciHiesJMq9zIlE+lkGfAd8qFBoLAkw1/TQolS
rqaKKDt5vp8gkGC7olvJYnu4G3m0Bnllg8x6ujIMNGL8I7n9TRIAqhwtUQpE
lhcIgihKI9FuS7iMHOJT1FoSYWnZUS84Q5gn4oTFTuAOT/4b2gueTNWCYJlb
ijjgiZMFydXIfBjHJArVsOz8ekhWE4DWuoc89Qg3vZU3IOzDONcOHo2/7LzP
Iz8q9o3GciQGiv6x61bM3jmg1UtoxGVufPXqESckroeV2mNBIl+jBYflR1QK
nbOXu6kqeQvnDlXjAkmgSHH5oDI4UC4f69TRQ3tHIPTNpT19gbj+ThRUHgzN
xcJ0jgnhmwWYtn45g/8j6NwCiE0h7kB9gnnMWUBtipmI2pSqMLLIIriVxujJ
0+cAU7triHBcb3vSGce7INBNI8Rrhi3Fk9q/U1y0s+RVsGzaL/XTSSyBqfw2
dgRutO5G1jldHyT4pnOx7r+hlKGAntCxSr3aSQt2RQqei8PlGAPWxEK6nIZq
3Od954bZWTj2RhUSPr+cdc123qYr0wPGrEIq6itUmB1ZQTTP2JIU45SQFp63
al7d6xSwvO3VNBbJckCpuXCnkNDNH8jzJ94jEDpKQm/ogJlXK7SnRzfakqYU
zQM/ThpLn3fmeYnazCrgAProHoE0w7X/Te+tZjEZr3j0FywF3If2eY/DONGt
A877xnKUmsyVA3iXYR/7RFGCKoL1QvNq6d/TD7Oam2rXBrpdotbNFMDuJPEG
ST0ApuhhVUtx6ObFD1c98RGgUmRy9vgGX7PRSJ6Tk4NpZiUATDth7ZHltXmt
zsVo93+0ZBI44vqLmJYpqkvtrJ29stubTfBCDWIJyPFr9uoh6t42svRskV6l
SBlcgSbG5ackkdtGn0d9uHN3aOS/06dCQkgHhjbtECIFEWbVDkS3+RiToNvJ
O15zt1845tZWs9BDHVHrQqBkqsgi0k9aarrBmmR94guxZiSTq9q3/lRUugtx
c092kRzW5c3qsU/CTHIHuDZ7yqIDJXLx2+a2x5yahyv3/KCEqJ2PGXNIIB86
uFpaMDTGtT9p9AgMH0E4dfIKYChzSJvdNL8E0TOYQ7JKRWo5QvZcqaoX3FoK
+PVooqy5Vu5nhGaEtDzQXqgHRyrepQPEyOCrklaksjbj8eBfWEiJpZSSYbKI
epjmtJO6+4ePnAmGhtAaaL5yGqCGaQrLfwyjOpm9/JYXbZ/NNlS8MG5giXTz
WGzoi5yK2tHplIJxQqmcPXG0/VnwIui+WzGmBPMweIkea/t4qlc7XI24qiPt
ux7o+zWVRVV7vbJk7HFK4Zh3myprJE4WFlb3yLB5qaJybjUfY4UTAibwojsw
3WUhHSSLAxAlE8esVUYtbLwaOYRviRWXEJY2B8l/oArviDPUZtyIpbMuS8fl
G2olsq+Mci7rYQha6kYWgSSkfkiuR5PLu8O/isakZvKkCS7cEQWWaB+UTT3k
0h8JbOLDy+UcgNdCxHvX1flzev/+w5MkkZngfIfu4OxeAeomC2d4kChtegwd
EK4QUnbuIhhhW1DvRKyAxYlk0arRM4KRvOpjtYYHTwAbzBuJj99iWrjUmcQQ
GKrvjvKIxfaIHQwz12+Kd+QuJF9VgvXm2Q2oqwuA04F7PNfZ56zASHVCjG3y
sqrL7bKpVX0ZC8QQFAsBUNUM/GVhZgpHRfCdGVNxa8/K9M8eJaTp50O4Or3u
FU/rVgEZ/Iu7f0ZnNATDEkhAqMGg9o+WkN5pI63CadbSrb67GK+KbKOFGWf3
nixvqg7tB+U+YgQgGnS16p0wFU0Jt8rrduzY8wENqCU8ECCVnXkIa+JZqmK3
deRjHTal2I4gRxr9Y7ZQ/TWC8iTYlzJQvzzs/tLksav4JudwEuUJkYjgBd8/
GnmCGkIfA/rfm41JnK6xu/B6aKe9jpR9ZqXPUZy20WuAM2iZYj3Jpen+zRVS
c7QrEBFb0IgyjSuyQSrfMnSZ9Q6OoInY9J4aJu6FPIchbCezPRzotxk0vDQO
uBcMDkT7Ye29DA9KJwC+oEPCvXKvPFVuxqa6zpJ2sk5+/UjO90bgQjftd6Uy
VLVQL6i1zHQU1UHyZlUBEye35zhiA0ytm+McMyOTl8+rM4WNOBdrSE3jnDBX
be2wHQk/L4oNG1DKrIwTnQOsASzIPvFOtNz4pjzIgZG+FPbniBbqBche0qQW
kVoj475UVkeHJva9bFLr/PtXEMDsq2dx1u9m+N0PkzD3ll9JfLrUoNKF1Gz5
n953SiHPmF03mUXnl63qyJM2HaIuLGgUUTfhgiPnkTb4PSikfI3Exm5hd8Qc
jWjUbwWLc1LWVh8BUaTou6xIhfALgg4KNVOwA0YUwOXRAzE5HOmmUQqc3uLX
ots2Ivr2qqhcYLwlDkHLHHeM7sMO2yZtiLBA6zMHS0gdWznCLNqmdAxeDuOb
5m3uh5C7MqpeL/hg/x4PTZD2WUFuTLFAXIa3xRjbZB9+QlFUDoxzHX3HIeXa
1Htlx7o6gJVt+7rgxvDnRZra1OrLWhPsSlbSrNIUYXVkfgVnFkZ5Atc0Y9T5
bmS1ymZjWaWXuD1eEhcTE4eX6L9zhE/4tvJXDOOm798oOqGsPFP77nl6IjZd
Fvum8hLLhM56o73xTg5zWsIfN8KqZpp+zVLd1S4A1MD0QVd8fSexSWzHGeTP
r3OTdrUXfcMkDUpEsFvDCHF8AYj71VbjWVvAMRSixiLBVX1WcJQulYv/mp0d
U8vDfxj4MgLycvJzydj5XuAEIuBLEbSJJX1+8T0ltd8ki+71bq50UPctSsBe
nOKQXC0UXabKHiZFGSvWS1nhmFnpcntVti6klNPi5SUJbhCD2c7ko9xIzQT6
FqJ48UsAH9M9969PF89yQtSAFzRaov8Nn+gCfwmVcXYcVNauz1WuUU8Ugs1M
ZI1wt0LyFy1pRoM3PaNudP8ZseEmGfv047Ju70871NCLgsgojL99Vey7iATN
Ofk51R+3w+vO15z8d/iUqxG2+y9vrR1azU/kBbwokGct7I9NsJyV29C4xpm6
nCiqHNajJS5/I9Rh8uBZcHXuqyAWF/2DxRzH6XLKxXkl5CNpd40REgpjGHbN
76wqNUDPkRjsmE1gBhWXE2T57SRgGD0TwHxA3uQdCm0T87SNGPS+U/IWYHGl
N3+tqX7N7kD5cMz3QqM0THdVUjWgO57p5/wzN4ai2vHk74oz9b6phRafuv0Y
RKYH7PT7o9IaRKBlIpfY9KTsNw5PsZNoMkK74oVydAdXT6JXLP32diAzD78P
vZ0rWjDsSI26BFW0RdClscvwo01rFbhUcHv51rGYsaG0zCROzwDa/wabx7Gg
yUxrzxPaRrumlttMjR0di0Ro0DvgYL8BTUGUHqInQxq5AMb5nq7cDn5jTg/X
UJZTip/mrq1/AeRWxO3VEui3Hdmd1Uc8WBTbKvTPB6x2iKQvWlWR5ViCba+J
P1zrmp0MhR4K0yxh2Ths+twVgSp6u0yQyYvt1ndnf3206DT9UIHmJ3dvWof1
8aQaE7nJJYGtjLYfbkjuRIlB4jTHhmgu7umUNM/0CbM/FP0/MC5exKwI7HGJ
WNyR+mBlvIkzsUlNzU6ClFl9ymCA17KujLAMOmhgaazrxBP0Z1fNDB6gIZfG
2wbqu/8cGNOVSEODhcBusTAzj3CDqnnzQAL70b1c+Kp3gDDM9xUag+Y3Tn/N
tSXhrFe94hC6KyT0b7C3AfwH1wzWU4Qnz7a/2rrqRwrQJxPKMPGQS8MJJ4zg
MMXD7K6h6VRXTfKhpuvTLW9rTFy+x5HBkbzk6Jk3cMHc/ZPYyLUf9YXVCR9+
BTcNO8sEIHEr/T4aWhvs9ABrq+COCpBk/MgC8FJgMGj7ZF+JVFHSDf31No71
GQW7elYPNTSgY44r66xlB1D/VUnwCsREVgOgHDe61Dt9NLRFr6IriyAB8G2h
DKLwrrGAwB1SdsZE6AachcCPGfGdMrYbG6idUIddRUcU0aZsDe7BtWTU+bCq
iC1ytqqaltE3ctEERfcrXel06T8SeWUx4jnCO2wM2+lz89FRrZUDzWR1xvHO
ACdzf2GrCvLSEZ9jo0HFsAau+cHb2JfBM9xEVyW/MkAnbiBjclxP/azrZY59
HTevs+qsSyc3tXkuDMKuGaNuMWxcrj6WPanO3TbyJAHP+fEuamiEXH44gwL/
VZILSKMWhfWTtCz7/UdMZLBjnP03IVAnf2d3saDEvp7pngIIYS4eakQ8aHMx
jg1JD6uXvN6wYScMfX+yyeN9gK2hlzuny0++9tFq8T5O4H7sbn6NrMG+HNbM
Im/dIc0wNK0tNqJVUW2bysQCvchAIwSPKXsZmGhwqrvj9Sf8dTT3bFGHw7MZ
XH4ced5e4ixiOrmaCgAJSJw52jBCL8c08QbEy+qHr4hv+JvZrsM45Rp2iaar
8pddvmW9Dyxx1bEsobfkAOPYHp7n8PcZvEbts6zTNIpqQeHBCq+3ITxQGQFa
Qgyf21f/zxq79MScRZn1FtXtBAE/7HkyH9MuXx277q/+30jJWJS7sxuHy/BA
YuOU6Ul7yNkb20RMwo3FXitJHSf9ChIWkumgoEnR+qDqF9HOvD/nPj++knt9
blP4tWkLinVlTTDvb5BibBea1JnLdG1dhQCxa4CqlZAw30EQDaNISLIsIpZQ
vWBCqYU7IsWJCBNO3hBmPLJrans6ybJxLfat1g5Y/wA+ioq2xdmkkhl1cQAT
r0P+3x0bISH5O69WWVMSIn/T3/ZDynJU65zyiCpQ8rS52wL8nYBZHtkGZN33
kzVY9Vk6NReqnZmNwd/kQRsMCdNz8mVdPMF+1lHENYpdmaCgFy6rdhyv8rsO
/kHVc+y1WNZjn+eFfhCCNar9PeiwoWduIeOKV0RPFCw9FOrmESklAVLbnfux
B/BdO17eqS93sfaKYJMotaYyx+1dWvGkXu4GPprwdm7VWb0pB9j4ak4iDTBc
5ifvRkGG2hNF8e36mvOVHxABeghvNmTo7kjMwWf3LQYv3PLQPmD2SPNjDbMM
rJWT3s9PuCbPnSoVmvIahl261AYr+uq+j0LjZgcPSHdLGVq1+6XwLUQ0Lyqj
tnOgDHyenzgTip5Y55favatd2TYJKi3jTKCHvPfDIjnAtcrhJRAtzNNO2E0M
DX9jSoNXXJ6+hT89x2VPuz6yuRxwLk0HIBf9rQmPPaXLzeTyd41Knt+8JfgS
J5XgNioDv/ljy4xUE129xQiWxVl1HaDfJNKQCFqIqmRY

`pragma protect end_protected
