// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bp44cLKQhNRxwVOwmCqBdG4aX0OBSRoZ0wS7PlDNwwD4KxcuEp8z5M/U19cf
Wnd16vZhJql70zlSfuC+tNA14Mi0WxT9IZ4z8jeWoDh1NPjDC0c5g/4Slv2V
/MXKl6y+TWPx2Kg+LzPsSlhkaVd/ab32FfjQQTuGUOebD6R8A14RAUWBIKCh
kcSuviUhgNniQrxWy8u0QVthvpJDx1cbddFRonn+EqPfQl8qSt+3uYhQlCme
QoolOd2Ly4nKUOzRm3eoAb8jFTV9z1YFKc3D1HsbbUQ5lJUSq6MP+NB3wvZD
xZdmTm4hy/42aUxJna1RNisu0xeYvtnqMCPGrT0Z5g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kKbraJOFLXCH27EU3xnzjAW6R2zxbT+/avVUqwUcEfv2cW7ADVPf4X/01G+Y
fEmUyXp0NZYRnXXSe6g6sDjF9BnGN77wcLfhDbkNNquS2ZfnvCmyjYRk/IjN
QUWQKVdBHQ5fqVBXnooDJL4R8bsaZDXCWjlUB2Ok6qnx5A9DIYzD/UhgeW0G
d1GXCzfhMZCSKbBqV/mWki/SCx4q5mYWu6NizsSddoA3YpL99ZiQ8xG+9qTu
pZdUDI0Eqg3VOC9R0eR+QjNEienN33GNKtpUFYvDtPY02jAs671l4CSUdb/U
GJa7JadqI3T9xvPM6SGFs23YdmksTpykvID+y7T/Vw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kE/+3zMbZGWKqZ9ZOeAy4+b5M0z04RKj5O3urhVIdXudXByX6umEkkp9Q95i
jGTqspsIWDYAvr4v9wWKIvbyMxC3y3LRoC7KyhvbCbec5GVhK3HFB/9j/xcm
Bz4Cc8G2rN4dtiJyyzfH4agZuFHYcs/kzQMEA57xFrgxkDcWtjD8ysJg+U5I
uQEqoXH6lXuzh+JhUvtjLucvXEeWA05hmx3DbK0gRKsifo9wy1/TcC/zaWlT
EtVUN99CWoZ9TIRiRU87MVbmjztwxbdNFoSrt5C1DC1+AFBNgob/vpKYVwMo
2zuVklV3kZzWX0b2pio0W3/vA8g6gEg1o8GhHULOZQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HbN+du+O7Jb98tCm1fzYCE/7lpCWk5dwlFrsy8/KpBhMsRca+OjzL0pctbcI
5OzerBWsBwSOTyGt86aCOZqt2ICMaHD7elVA6b3EMbc7bIaT4jDVXORvEf0z
kD2UPoF4EF5oyx1mQFd+06qggj54aXWp1GV9g5ZomqDjXvtuAco=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
udcgnz1bQMEOLHzH7u9G+6gSa37MU/IFZXsyTSyNTvOpTjA8zmW4m678u4BE
N/l6TRhANjwN83YamiuwZ9+NGkgyCSBsZYXjnyNior2oWuvAjKrgMbfXi98p
qv0Q2f6iC41D15xs7W++8Hxs+WWMEcRGXjy2HSo4vAT07gadj5+aff+T7OAS
AWfGFfabtssBQz7lM04srLhRpPy966bVgLpQTL9DsBPeIZCZADF2w8SdnCcy
kGCGBZHtkZ0JFIJZFvjDTt6g3AHz1GnGQMvX05ihFFnSXf1XW8Erj59IM15x
90c0S8br9LaJ2VU/Y7eGlsgAZvwtYwlUYOG1rSTDY7+OsKjW/vvqeikEpH10
S001ZK15sYw0zzU5SjxkzWfJX22oISjR6BQvBBcgxZuHE+p92PGMeFPN4YvT
rzkG6jevZv2Msj3PA3R4BOG47DwJf0JBYZqP+LNnCLGpU2D4jW96JmBcAYH7
3z20psdN66mG9iAj+9csoTliEOmdEk5Z


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eWxrZwY9rNSKjuC+WDwL8lgNIZX2fz7wxEYYQoU5mkEShhTzRI0yVg2AAdIp
75p3GYJoJHxggjbg8Iquw2H99Lr+BdMQs6p+1TTaOgy6KOM37l86tknqX3cu
AO716N6bzLympX5CAno+RNGfGVu5h5SzFVOkQVVXRPsD9hVaIuY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fDr26u03nSsAhQFTwKhq/0ZSa4fq574J330lGo2wHyLBdGQ1MLlQcYkI+D1T
hFkSXJ/DJvNMzlwdmdtBuDi+3K3Haf/5Kj5wY7XRsh8bmNRqdfUvXFgsTGEv
/SaZ52LF9gQrfWsli9NOPLpLKnJj3fS9SAwSwkShz+FLKk37Alc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 924576)
`pragma protect data_block
PE80Z/1CBbzi5RXoqww/7matkMJ9Ly9NzvBevtaV3JcEnjKF2NCWzm+Q5V+S
VN64FGNZKcDJviC+5SYT8NXDPxkHhlTMzc/2o3xpUerAFuIC9DWbSfuB+MQ3
Lzud+n4c2gAhqKlqOvtIVcdL1N6lFiq2NCF1v3Uy37jqBImP3IcQOBZrf7PQ
CqioeYzDb4P5mJNJfRQ2wfzJCnM/LYqEOHhRgjo2V4fdgMt9w7QMVeLOM2fb
qugTXBCtKuUS1E9s7C7jCLThZW69xo7zxEgZoRzdOlaKluFeV+0tDhiB9cyQ
Jq/YaWU6P7HJczlrw7MLUM8LC1Cg4aHIWOCoTo683Rq1fjrf0DizK8omnLTs
/45you5IYZRXDBGblrTPyOQYnJMZagrl4ceqjYPUxLBGj+UCncbpiQzjgZmn
OqYBq0gcpkLtQ0z11E4l2PN24IfUP6MkUJGiOez4aLS88jTJWsMBywI/jvTc
+tPMOhJRfEq/k4/A1UK0FCTDaF1bgLNmmu1biz0rqvTfoEE/zggWE0V29e3s
MWDF1T1etuYrwHMkhQ/dSwUF88x4ASGpfsJM6Ps+bWvK7lxu4zlWkJYjQ2Jt
IaJYVQhW4dqbZhp5oQM32C9kzOlP1CYMP05+5KPhxDDozG4BkZSKCxpSSBP4
5K2g3KZqdnbdlMb5pgkDj1qt0zWJMsBbQAZB+Z3iq7QtPaTxvRont3dk/6tW
ICAW/IIVDV4X2QGeyG1Hl2tJ5VCmCYVSbkOjfHctJti1OLieAoj7fkeaqeuc
CKEToZEX9D36FUaYFGcztjNs0J0MjZzc+56gFB0PVJhWSC5FTFk8x8FYVQ1c
ANROIMYAVois+kIBvoYdd+Nri6+IicWRnY86iRjWxoJdRd+h6vjMgz+vJ65l
2k6hpVDl7l74hBKX+0A5wX0CFEhsKRiROQ4krZgT6sDQbAb9mLhorffEEAlZ
SK/btfuI58ssrg5rguDzeLreAn9HeebgHP626YC7jogpbGYNNHaqTsMZhoFl
J3zQXgUD33+mZWaBBj1sbRGqX5FxxYE/VH4AT3B/cvPo9NhuIoR6stGpV2J8
/v2bbWl/xqrt4RW4qg9rvoSq6lTaNRC5DOfS6Y/VFsb+ZerLarYEvy+vAVlg
fg0rU0NqOAuMClShrqmH8kALsSww+aNt/O/OXrMmXo7lGBpiazhOXqP6cpAa
B42ft6RR1XlNGDlS8fH1rRzSRWvnvGrclhNcaryw1klYUcDi/ALMLwfYVp8m
lvk375BaDiFQi61uhAX6CeCwgJfNDqBjsd+czPMP9v1BseYTyeJnmAVI3P2c
HZs5QDC3U8lL2Tm2xECRWFWALlcsTHgLSnGbaIFK4mOOLRLYfZhRs9HgRdy1
1hCNm4cnn9MJucn7EHwpPL4p0UcJ7fxHRloTGjHlVNs1mmabMMhx4KPlwIs4
e6LsggzoAhYH9j6Vtv28ssFg7aOUv/MZIELDtgo4lzKzDWuLEk1UygsP0AUx
ltTwEsoLy1oNZK0UUCPZuyIMNA3P0Iqkf4GPUtc5baVFbXO5U0MmFOZNQEdB
UTDY7ubxVOclZmeHS+ef0IzrH6KBu194ltjcbaKPhRF5bAU9TBFQb6DmFQ2h
7QhNfPfDG0VJFIrna7R8rC7+v+GHP6elyGIW+SaD5Fj4uVSSo9Z/lJJwpQqe
7A5uqx8KbU9gziwVCimm769ZkhpaF6XfiaQy5KE/QsxYeP8xaqiNH8HOUnpJ
qtVS23ICFxdgEXdpqEpdhUNeW6tG0IFY0JaaKfIL8gc07rWzE3zlgsZW9vxO
6H+679GfasWnh+eia5Eim0e6qL//ZHmypVCv7w81/PBFCOq4vhOBcZJenPJ3
mLJ5a/0BSb7EJ8Aj7ETwnJqno8P9dElt8GGLsGXtshEZyOgfm/88ktufZTwo
aDT8oTZISYNXEGVn+fYsoix9mTS2xoOWjmRacdwdfZA9v+amG/juV7JRMMZp
uQauXWXdkw8Vq+eOd90r4znU0W1xXx1VHKGiApAB5iTmG0cgQxuI8s5wCFb1
oOCVGMXU4ZEtxx369SIrjM8CJx5UvYqC9iUPnivqy0XV3/X93Bpm0/Fqk084
nrRF8Pt6rbl0dN+fStcf9m7KfBfYHYthTBby//63KbURlyWihLE+f/43UJir
ZgSdYwT957SEs+y13LEcFZAO/24l3mRzRI+LGOLOZSxtWRSHo9x6HozBWcfM
rnm/+korLcjDXaJOYtGPEheyW9zIIRbx+83DTPNOSYjYzco4SBnNqKS6mYYH
RZ0iPqpthv16olO0IK8ooYyqhb9jdZI9wpuKUwIfcmQDFGLFbRcFroWt2wam
SYOAT5GQi2cSqLiNQw76QHS8xTQ2KGPAmjPBqrTgh4SRxIQLJ74D0RXRooM9
+w6T6yM9Hb2EAZx6cg21LaPeUOSoBi0/wXBNGy34m0FI1AhO/UmkqhS36aZV
panQW8q2EFowbYyZrewUvEQciIdoYgwa0VVdHVPzJ9KSViFUqcQ5KUHQ215g
H5ZSxsBLaWNY12prvfDIHFMsuOAk9c6dlm4PMBoCR9FRHM0pOdTYpMHkFpgO
8447d1SPZeY3StIj61mg16AqCvyTPANttt/ZjGbQpvGqKl1DmYxCRUdI/bb+
VEeZZcQTBBenZRYWJY+boeO92E9N8pDVzI6xUe45ovnUFytUzP220oyn3usr
y2m800OGHgjhuZU/T62v/w4SRnuEUr6LzXg18wZYoZolvGpeW9T8JRcCBDlc
CTNUQeYuDV0fG9SoB2jGfB9HgMzPjshnxFAynja1xx6Jtqey1vrjL/HHhfGU
zzX9kCLDU/yNCJ6ZK/f3yCkI2UYzXc1yCTtME8qAITahNJivD5KFMpqqR8/6
y0qwRRap0Y6tOGaO4GUtRry79lEWHyVNJCQZIjrnKPx79/E7Qgyl3W6r74ic
CAalzA9je3D3kQ6MqNim0bNpvAK/zw9gzEAvkoptOKcUdvoPeviPO1ULOVkE
nrIVRPKEMf001WVdJP9d3Rzyxa3msYt4wkQ6mfAzgNfhcnnFEPUQku37kcRJ
sZu2x5hbjz6jzPzLK4CbeWIlhEjI1SbxFIJkqRozi7xjwu7QyCSpyQWqI3IV
tHXsgGTVuP9MZT7wDFnW8dhHPy0+YGEqFOeBOj4xUALsMkogO76JGh+9F90G
1fDjTksSrYz2hvgDCcoAwTwTMzaCagWAPmFJXitrNsr7dHVyIvBSqMU3rrlO
TbiHXw33IzWNAKQw5MIRdpQ2f7LisnaMjtamWcZwzD7V36VaOeqNZuVXC78K
FqhlJrpBKWotmQ4O3v7h7UOZFMOKDhRThY10kqyUafH8zx+//4FTxS6MgTup
3DPBrVEG/8q22BNJXud4NoAPbBVqpTsD3y+eCKn6RbL96WJHsx0FDu38shpM
f2WAA9Fe0dlS9w9Qs6euVbJ43Si68SMVQCoigNliw4b6TfhRw1XADzuokHek
7+I5FuRHPCng6uzf68EXJswrV178Fwsj0toYH2E9f28oG8KX758ecJ/fNScw
hFLVLuZyUBG2RFj41H4oTDAFYnFvXPyIxbZD/cIgBs3aWqE5u2RG4oMDSGMv
oShD/vvdkuyEEqugjU8k95RxC4Z458B/3or2ecHO5Vsl/yG5gH57NuOlH0m8
Zq0P98y9agX8XcWqYvWCfxd2AHQKo+YJuLJKLP4oQkJMCUew5k7VLOdbgu02
PTXZAnE8RQh/eWFviYGwOO7474G87q2WIK32VQr2JRJb77rXU9O7xcFRKsws
ZZaoQwDSNHEXURye7AbOMgCq/9CDuRF+tJoaroeve+DIUHjJMcBe6fvy2Hys
Uyj8wV3aD6iKYOwX5t1Lb9r6T8Gw4O2VKnLKHJi2NdQWZc8xBuq1hLfM2mws
CyFGcrlYgotciRdMfnCzH7tl8rzQqlSCQx8atzX2GrXs88bvwUSGswkkigDs
O5oWoDEBDSeVO07FMcG2RUanq+miqgfEtWSeOu/3FGBXACxcnp7c9Rfq3PRv
MGI1wQQX2z1pBDMRRzcuLeLISLUx9ZYH8MpkV67gxgxcL8QerZHlORy9GChR
cNePwMkrbXfNm67WVdzX5UdQ/N3Ps60WUvvtfzsmgaDf/YMSFQxsel06aLpD
1xXLLwNtBO51Ccvfzj1WIZOOZtL9zyWJ4kqU0meTZfqaVPUlnnjkbgcDYVrM
BMKOBuEdWrfAfscEsCdI/RWIxOK799+/x7KjF9P6qdGW1HFnQW0Kt9COLdr3
tHqtfDVPoLW+KHwrchzNa0UbDGQC/BEtxwxb/ieesYc785Xzj6XFVYdscmtQ
jiD/q5ZZaPwJf7FzY3wWV6eSGsFlSsTx94B7VDfKJfgAK+60BGTTc7xSZ7WM
BKFlUiNjyx8wLs8d9l6mJ8DBJ/i+/Tr/M6fYLkRMHgTVHGKkwyCM4KdqQjF0
iejHzZsYiUZRpJuwmAmOmno2WVUGAGH0Q5b5HFIVVEMhAQivC9g18ZLuIXM0
oD6HUesTzZL/uE4VpOn8+hhQrbt/mMvDJhILzXitN1J02Wbkq+gyHDSUKD0j
+UVD4RmTjlF+RC1N/w/rZRoi4J1qIVJ3MAnZpeGnPlHfbhGxEUsp8EPDWpTV
2+/aQtNHCI0ine18IbguPigYnMIy13eLwnV77NRLeEtQzD+pd/4z/4C7FgDX
CsjFJ1dwDI45Y3mgwnjWE4eWY2IGeLrtJ5UvK+46ntOIIVhDUtZzH8r8Fknj
0DG8zS6BTy/ZrXjWuH30+LJH/jeEuDpUjmeioaawRUX2rK8lookdGbFz5itQ
v1KNBE0RHuXZFMm3Nb0/G9uatsvtdzu64hccmo5+rVPegBtF1j3cMYGyd0D2
W+GRRxvTFvEwCJRBScdbSFA4mAUFhtRmS5K23FJeYjrSrjRDgyC92ZqEgy7E
X/Vf9HUS6OVN5QLBz1WKvbNuFlNgCz8uUuYV3HSs+gtDxtjUK5wM055o2+zi
jHmp+RXtEYOnrgwD1Jh1FASOVFFwjxpG9WV+1evCiSdMVoXW1wQiLKSDvgyO
xJlk4S7PO3q7TlBrOMFfpyN7DmPeW8++q7bZF/v/5jY5kNNDc82F7l10nSeJ
Ihx8DQkMWXSGX1Tmy+knSBEa23mYjbQozO7ZdstLEdXU1v/gyF63ezcN6Plx
u7jpqWtthHQmvKuEHpZnhPoedOOvTY3S9VM1ssaFDAmJt7Qzra4uN6oYxDtA
0BCXm4XZo97X4EoOn5sknJV0PtquABuV3Sz54B+av9kd57KiwWZQYPON6DjT
ZeO3BhIklnSBpz4HqwmFu7EfEO8cc2D6RMNe75E9Kecc86xOKaqzhTzrMVpR
b0gcdxR38UC1Pm4GmRcE+rTaE1HNRRNe8DfKc+uN2L4xd3wqlZ5zZT9aaeTw
YUuMOgvmMYxS8egkUOPfBOjvj0byITzNdlV7b5SDc2ZdG25zXLaGvQ9EwaP+
LLsrHVobST2xEMiJbKZZy8b0JglniXlV/Rh8OeHdb6K380vsKKhylPGb3Z0a
0m5ZXtOn5pLcKrlyoiyMGmLQNBneJsPqqly2QJOU1KamNnnNHeAg0wEAv8P/
PvOlcV8j6xatB9xVimBhHAj8PXyWw2Brxz7Ewr4nIHQAtlm1LBdzSoOdlj3h
u0/qXazRe5l+VeFqqEKouxYHD8xgES2iqco8izn2Pxnjgm9uRh3uVcMViEof
kPy4KSHl7SSQLQQdgHDl3cDbqODIfjx7WGgo/MnAFGqUimQaSwnF2XC1JEB/
mK862z7tjqOttU08lICzUpsOM1Nyungf3QSbOKOAWZ2oFfnQhk4nD7kWpYUP
9lIVh5TWRl1WnIkTOE2MWGMjGqK2CSJh80odJTZDF1ZkZa82rTuuIUUj0XfI
DVZHCo/IwgqCSdRZ/LS3WkZ/b15cyp1KLFUFLQjkjMBfhAABVl/TYMKSSz9a
Q9qwUe3Mof1P2ZYnq0QT1G1y8ID6lRdjVpx6gl4hMmOBLaekJKlRh5jwmGRh
87wxLaLqjMuRtt+e/t/wylBKSp4UGEh9mQWu1wnTh3CRiXhMo4gPmCjlEb7b
nbEXXYXD84pnd3/DrncnnsBUOueSQPjfDtkQK2rRQ02QbJ7quavYaEV5d09c
BOqB7CzF7KmGfbmXXSf4cR/Dq4BtvVwVlr5bd3T5bpZ2XlZ9njLpkWF+3R7g
gGu816OPEGmcSnKdsBneo73VjUFxS+dXqCKck5KWhvgkZ3WWSnNN0Zc3Lfci
9XlzdZVmuc05VS2X1qSFPk+HSTq+0z93polu6q+ZpLIrJVBtcK3sFowXy1wN
tDUmPOmmjPywMP4rI+JyTujh3gEaQ3vR9Hdrt4gSU6LO3xzhl1gv0/JPGnMV
zEcM0b9tvuz4LHnD59/t8biOnfpNYWQKPAtkKNyICR25NiJ8wxkZow1Wwylv
ExTKzCTyoJh8cm/bFAJIlDMe/w6OTcFzsJyPqJfeuASTlWsVCrQ7BSQ92epr
Zfjda0iHlPJeM6tjSQcZ/hkVso7hjVNzYC8HLdOBKUw2AoxtdKY3K9D/INcl
XElP4goDx60P5gjV80QGEagw8kCkGTcS2NoUIOrxVTPKNpJGuMAU2rE77UMH
w/nk35adPJbJQFIfQZSTGNao9SUAF6uOLNXW/frDVKfEYkZ6EMhI8kOLZXO8
0kST1etuZ3mV/1CfbzxKT/tYEvmGbO8V12WnF+7tSF8aFM7JVkWXH4q6RmeX
2IxY/LLja67CnYNJZm/FE6fpZgyonXAnK4HiNe5OcYTznwFV9Cz+aXlMSn8A
uNnCZ4TeDMyuZ1lg/EVhxl7COvQKDi52EVBXHd+voZ4JF+z1yeHBcj7iOZzg
1WmRyQns9Th5QvW5IzfPl724nwJnL5jXaAmQru+4CBJJsFE0lCnuAfwWxw2c
/hfMFsQc+x84iWt2m6xRlD7XKFkEFcDyftsYntiaoyd/nbT6QkfwbrxR+E/E
lLj++OzfiHWr83CQPEKqwNRm4nlQUxNCxt9V5NLKNPhjLQ3cxTIR5fmSEsrv
kKdYc+yVE9epvjtQPDo0o54XqudHyx+bqLs27kMakMnQL4xfU8j4li7LzOvQ
cvz3iPoLeyjrM5FGPKUMCK8purNii4BUTEzuQi5+raRmr8N1ilgIIx0rO4NF
bL7DCjuNxQISz7xhtDbU/npKIykQ9PckTIhjiSDzK7zWPeX7FvxqFdAqQ6UC
IA7V/qazp6wJgYlk60nccA4emWbzlnnUgGTJLKSOChCr8h96Q73WKT6Sqobp
zZITVONyBkIAmJebn8ggnEMOuhH+LKwyTKm1lIZCVyYg6U/EYvlve9plfbnP
Pa9T36RZ0pTPxxpeSsPglWGi80DNsGyJ+/F9i40G97xPqcO76xn8RqaHT1OJ
VYMW5HFszfCk52sbipMlnCIf/J0/PKnnPHy3OCfCAnUpN4VXROH+LHV531W7
MGTSgATyra8iCcKpHsM0HAWF+kjGn4nqljjqhvEYb71vJH8HmqcIPJWa64ll
LQ6ANCy3KDeyZpgTmSyF6A2lcF6pAfeXHztNqWvvqmshmEIsmaEmr4rnOMac
ra1KNsH33qkOcOJI6crgkae8WM+WYdZzWPdaixn1hKLK3FU2gqIIJBjKzF17
/XqGlk32HrABHiPo2FpV7CDSAi58hUTxrWqQ0OyZo2vDhSfR9R4X/ksHzCLd
LWC+bAH/qDJWEXRQQ5siOrUYTJbMgsbOMOzB2UXUEanKYFivDJ3dYDyqDl9n
hLYZgAwdWw3oSJILHGoB4XrcJJMOGCyC3bJkW/eDt5PVbAZd5Paf8FzBEo3E
4loTur+Abu1ldE5L3k/DInZ+i+JcJNw0PGm9cJENHMDd1ekRkxFqePpEJ/VE
EUc/+c+k+/k0eUrMkn8mWDIlSkcG7QnRPOypuAP1hShZnFXICwy/3RRiig3Z
meMFDgvpb+hzLFNVIHj7z8oLPiBXyWoiKXr5UPmzFMVIuo7N1guZJExJolto
CXEU1C2wHQQDPlkPfcsYsnYNmPW7aGVYedw5QcB6UJKwry6ZG+AGpF1LzDwp
up3HTdR8EwprDzR47uGT9TLjyNEqD462VcZvq1O+bCXTkertgCNDy1exkt+F
D2rVUwZcyNGiHN6s/ZVXmts3ghNu/P8YmycTnrsrCaGICM0JH1m1FUEueljO
rSobjlSxUsm0WfZPIZUiSeMAJvOAX5ozLqrBPZ8xUocBkKKP30rcoICSd3yM
tXNAwzMt31vktvDFxbCAgVPm2fLM0zlPP+IiScwQaLcramAhxpEdEdekp+cY
lUmWWb3ZDAJKOwaQ4yVOLNAn9Pv/WlVHIjcKgGLkuA8iznWl+N7gKkqyecYn
IZeTJeLYTwZlFubXG1k5VXj219wHWWx5SYt2TxlGWAEVwrrm6h9cMGkFEHri
+KqVTzFFuGTZhBHRdJueFKH021a7a1wW2XMBnGHTQJU9iESeRJMpARhnd7r0
c2Fvucf5LNqpNRHxS6rebjzV7WI0nLX8t8de3gs7UH//MAtPKmpHRKZNlyjt
Tbfo4EmKpkbQgGgaaruvAMDfEw0CM4nd3GY9nodZfv4zbij5K6DUA9sF0yl5
v9R2h4iYlp9pgxlaU+N7BvTikf1JAlCoZQQHnPIuhLNzarw7vsRCpRPZJ4OA
2kNv0vUn9jJJNgrXQ8YSag5mxKmwaRjcHRNebR85962MIJ4+1f3lrywZIJB8
LKzAk0WBsCGZbKvVvMqERfV+lntD9G6o+TlGRqPgeLos73ufDSFdLzubYA6q
eYLrFYdZD7zKmxbUdxJXTNTfy/efiS/DZn0P/nIl2b/XCIe6t0qJrYzFIFqs
Dz02+YFJlmNLuy3nYlem5p+ANp9Tj71cax0yBJic/+0Sbt59aSmMo03UARcl
qkdmp/yeoR+Rmdy+vpgRCYKtrHGzbR+/yCqIq6Iekcz2s+JexIEOUcw64aCJ
YFOUNXJ8G7zbXC6cT6kgOwu5DuOYabpgX93RJBZWJ+2gPX/QuZd9vm89QN14
gF6ENfN/MIovCUZls3CtTj83xQJiR5SvjKJkgNIXugsXkT8f+0dhI6uc3nJy
czYNvmGOqUl0NNgk7e6pkoNmVxTHfBwHl68oKQUK3SVnAMK/BUgXd4/HIfRv
+sW53VZVyhKQqJIwUKdVxViNxy2jzBFcICZf44Dg1gUlV9lpjDWXsnFJJx/F
YQyIDua/DRdp48oR79Djvdd6qM3pPdRi2EUDXW0aafa4d4joDvMMAQUTHT3x
XrXvj9J9ZECcJyVlWSrEoVy6/HHTXUuUGKvQFoT6tkeJjcXBevTYVJp6tT9t
shXcirIOxiB9PNj/CLwifEu+vhW1X1s+uwV1ZcbV4n0Jsej3XyuWQZ9+iCJI
TGlFzwP/5JDlIo+CEZvua+EsZzvxg192Vku5CgvFI/I3dhmIlhc3qTGE1m1G
bKuul1S+Lkedz/mWnm4ZgyIUM7aXQ/lIavtY+buVDd1DQHFUPDqVQ8cYz6uk
ToqRWIb9bMXZQGuZ9jIOmmD/3RoqRhYuK1082EW356OnJTXYdI4CIszwPO4a
YgfLJoXmlOUgSfBlz3KpD+pw5QNk1FzN/apyQwV53vuVxZNGypAM2RNNHq0r
E/iiKR7RgkMh3pRwZwAB/SeYve3Y0Ht7kqzQ2OIRYWJR+7XPumZJLolJcTPL
Z3NwU5CDtUFu8JAwOXibZPtEbXaQpSlIIgfLmcNYoU5kRSI7xszZFZPd0qcW
s51QCQZu9+8S8lL7DANPMyeUEVXqmiCgBvbbp4K6vXxYXPfERRoXJMm06pD/
hFpJaKNwNgoLv5cGDXxZ6+oC6Hh24QexOUxkKtX+TBAv0nTV32WKWpbBMm9M
AYeThb0xVG1G7pSyPF5198mimGuvq0CQ6u9iAM5CnMwJe1K4wJESBFE3GoiD
DwVstOgTGQ0vhcCkRK2sfolEiDSECEkbNtkWBwKkRt2tkSXXAyTrMns9OB5F
eZ5pSBgcjYVwG7lczquQAdTuVvwg1Qt/qLUYR2Ohg82EAbiqyTiGxzvtMY7X
bTgl/Uyqr8eeq/NDcL+yok1axJeH297/bTXaXl6dZt6MU1hoEZSCLSi0JP8q
btG8EHsLGV9/PX1mMGqGgWIC46bpTNW5/jdeC0tbe5CAUMP+3eImahBo2lKj
R3/qDM24ie+7D1WaPKlF3JLF/T1JKi5sGyLGSgpS2GmNAlDHeOx+c3apF+Iz
EtxvwsU3AE/0UQLoE5Ukdnbg0t+PRpMKKoBbF10rVqkJFohuNheLw0cj5iNr
qv8BegbhFrSTDbViiE4ANor6TSS2d1kaSzuBuZNeGU72UmV3n6+xXV/b48ub
Q9JC8ONrof96s7RgCon2U0UwnLgemA02DvmOEaeLAiIkyzS6eTaJynSbe52o
UsjGczz5BcbVEFgBRMUlx4X7Wp7/yNzW5i7vX3E9qmsDujPICWBC1C5nsTpj
dSrzyIAetrBuhobBgWeKDzUMIvA0S6AmAz99uUTTYQBYAjePnoGW3Wxni24N
gn0xPiKkf48OxjbjTEvx+z4zB1iCBovVxnNKjuvWnbpwtJtLdAosuWrsX2VA
7nEG8L+suMWGF/Z8QpWrE3ihj7HfVE0zhRbTfE+E2XfMmD9MuqRLJoEEXcSe
6sTxRFkN0J4xTaWCezxfXsSS/fmsLDm+K9mN+eurjUudwvGHL3IIMti7kSot
dkODOhNu+YPvmGsV/rILOXtR4EwFNKTKSsDT/IHGoErJu9ltc+8LHQyVmdRZ
Wkb0I/KZ8LkIg1AdJgkuVdGfDNw6arWO6YHApOWh9m/B3ydVxBRywoOE/71Y
47Fc3MtKk82AahNCyroJBRIShzRznsniY3cNnvym4fXbKYx4IlnUfFMra+EZ
tyEkr3Hqn84JK+FsW8A+PralOmMfiFqBTmMCRZdzuNHFtAApZjz6EkR7pZfg
U9I6lPaerkREuJVPe6i6rQO/uC0O39UbXMuPbzKM+ZsinL86Sa1hEUtRGu3F
k/4GCV17vgG6ba+ne5+pOCk77K/li6C9kKcLA7KlWuXXKcd4gsJK2KNwX3/1
X1yL8IEG21FEDPLPvw7BdMmwfVlJdYo6DDpgmr9nwGvXX4anhr346f1QHAVJ
UWZEya0vWpxWsZ+p0ix7a40geUTnMUq45rFdNLVn1mDnfwW2jacypbHR6Btw
EdLiLarCLdDPMfwZK+mDb+1AGIbAtoyc1GnXlyv4dRXuHdScMUotajthXF2Y
d1iiAlcHY+29clqElZ+8m0V6zmhn3/affIYIUG+nixsV/1kBSAYdNbtif7my
JEC/uGqdwgzXubYCWAdtQ7zW/RRosK6oxymwLpMJvf02MipS5M/xKFjAOYqB
HA465FqpMabkPQsQtGgPGrjDGN6xkY9JRGB8eEvJGbBrm1oKFJ+X/oUb0HOl
U7cA4pTiy5I1XRqFF2PRPY0QpEuYjjsvvT3c/jfkBgc+8t0R7pUHN1ER7Zbs
D8/5N0RY9wlaF6+xH+U0M0cBl3owwMb3c3w+79OOKQmavl1FDvlii7dkGlBK
MRA/ILDIfdNuv5S9MD5SnNtg/SFLrDo3RPiUlPBQ9FesN6SsjcWlLAcNQZzn
wEyQbeH8G+ZMt0t2Rbx3od5VEaYzFwM8ywatV+3Q4mAo4lrV5zqHp9r2k5sB
2HcIFqpQCIVbuT+kzv1rQYDByCnHnI1pmUx7kQPgwQLJXDKscUgpDjxofK3s
w+/kswfRsN/gML1wiy1HkM8ClP3LooJMfPUOSHcR5xa6yyB9brTW1zApMHV1
gtcXGLkfDyFtmOOilwYb+JCyY4ioWe9jEbuM7kEnjLMoLhGlDYm4ecXJon7v
e23JXoUgdIJy+kHYlOdDvDkVQi10MlBxHeY7qIOr/VBE+KprO/3VtJMDLxw3
8THd4EN+B4pmE2GZxhV8oqt3w0WvQ6dnaQVWjnAp5ScBY7zwLC8fuMNm8V5E
qVfOOa3s6LBByl6PVJ+yvfRW/Yod6oS+sIAFVbdUqAFW4b8xXmuPnen5Gkuk
4OW3ekSyPHHk9SREfp1rojtyV2dHWWYmtMdqQ7fE3x57R5/BTazG70XpTYZN
tw5dtN3eQYHa06lvO7zw28swvJ6eyfpOxx8p35SuYRYT/84yXi7l0kAPlYF0
0tXXJk7QGx+nRsOlt7uWUFeHwQYieMZKS7eDNC2WieKCEcOy+34XqIgG1wah
BpsluOy/iOz7as+FnV8ajclXKCVdo1GCCvjoMRjO9Dt5BihqNstv+x8lGxzK
jr6E82oae7NpVXHixFkTwQSdIbvHOL9H5W3NI+tMej/UE0hI9yndwS/UolvB
g/I4xzY9MGYGCDVQZbOWEXHcgk8X3HbpzU6RMQnJnhH5+/ioUxcAKhsSrx2I
+BzYmqESubxk8SCHuoQI9wY+mYM5/hf1hJSzA0hLW5QUbF91Mx8RQcgd88oi
5q1BCgMSwfpLDqcCuwQgH3tOTVFNLlUh98rRzXKSSPp82Iym3M9BFjAG/mwc
1xzAzvyCRt9BcNtgdUjPP0RY+Nqwc38L4nniuzULWALoWlEJeFPPe13SZdhP
d807J1qfcV3zjg8NJWEsf2tNksjkJWisJNkkoosWuodeVKxrYVWHHmXp8ZIg
LB240RHruRI5DFiL/n9rZarMP5XGq+dHaFx8vVC/u6hdvSYh+COf4f2eHLxT
eH10lxnAVMo9i2EjeuWwdUK4EJ24iSXTGLaBknoK5clxzWrhAGIgqpTcJ9Kg
e99Dsj64/DsSXnO066PirnnuKdZm+n2aohrEHCYNri3VkDSoChGgrLZprWGR
RqTPf1wcTWzn0vHdfCaeVmImHdYY4y8IkZ/FWllgHmjVCq0ULtLAgJA8BLQt
J65wxZL+JmRX5IWa+n+JLbODFVuijCPNPWYr+ohyFNv4gqPmpzP4ILogqTam
TEx5WVWSpIw3FgiMJ5BPCvPBjB2tN4q7xE/kKZ6cPIiRP5p99PVY9ekZts/9
sBEoVbM/5hxRtH8StSdARiHjFJpW7l9Aqn2ICoguYVBdvFbGwpS/4flRLimi
NgXPHEZ0HDhARSd72kzkV/09JRxt6lWu+TRMkIJx5I+IcKQrsi2wL9QMFvrR
P0U0D/8jKz8BIAGxKtFvqTpfqAOvC/YxY6rYKkfGlPI3t33ef5Pb4WJmgi2Z
uXutHEQg/1L+RUGuZVqmW3oW/zr9bApr64ydOiZl1BzLTvYtGIhVzI4I6znH
rLx/ia58FG2X/9Nc8T4F4C32eQZqiDsUIeFwvKI3or6RbE9y19tKIOPG2g97
2QapoG7mMPacRtODAbzSnq8zB5dPHH84Ai5Lr4+D04vS/t/fq5dmsTOE8R6s
YvnS35iV+Iik+pGwnuD4/Vq1V7lG2ogaj00NhvU/AFk248OhW/o5nDUqa9fH
E6ekeDcaRXBYtCyngCWAfdFA3bTf0PdB6ti7JdWuy3+myfH8Jk2qV/4izQSE
5LgQDoamM1J3AziY4pmfUGNTk67XcLOPTxpux+X+So8q8+Bc2KSCLypxyte8
jxTsLuyY8hgmcsi5idmjU08qX8rNEnJnCotUUPBCPtB4k0fLU6pvWprZqDhr
pnRjWQW00L2LTMnb3MmsIsTphx6/91SwV7YXXiGeYcwB5DYak0YaMObafW/i
dzm/zgFEaZ0LEMqMC8RlLp6RFcvP4ULZqZC01hrKdAm79JsHT0HGf47mw6Jq
zMZIE9RFxHiw+sLRxJwkIAsXyUNxLUzyvdnnLVMwYXE6c534Jr0LT9o76Hyq
7E6iN+Q8ZuHTbENF7AvruvZfc/UJ+aS2ouVwpRVp+/Cta7RxHk4aYar2c00h
0uzB5qo7Mgq7h8YT7eFJP+gL59VOrGyKCH5/1I/9+mMHRoqN5PddZ850jfgu
DdDNtj9q9WMsU6wsrafCcxdBpUCHIa3Or/+u4sVbHOJ6anbCbcEvol4o/8Y2
8jn023dZomYLXWLNZm0l3Q2Dq1/Yi+xAy/l5D52PV0Q3GOrOpUodDI1Ep5Va
tUfhqg/m5wAYIffdMCkAviw9nfg3fWon7F7TI5lP7g/ebLn7QwU3Ofn5Vp0e
OJmYLYp2dGimdeobfbiLHSM+UBgpqGOluPO05euHF9bZ10XSpnPnC48DBTVO
9jnvhXvNBh59fjPbhZwD4NXd/L35pMoQhK9v1DMi5ucUGvRHw4Gv0ecKxEKd
tQEyecXD9LgIT2mX8bNmiRMa2WEuHL8zxNhNXwgwis1k79qUrc77DXFZssts
p7KaVEwkOkN0RHQjbh+g13Q/x0q1Ry4hijlkytvEo/M/QmbSISfbdI23Qxp4
vQuwRIRHmg1eYFRSIK7UsItTCWlS8ryWvU3IUQbmVZiIa5YORhi6v4AAwqVY
5MtqfAbE5qBuBUq3MaFV/WTaFxNRbbmUIiMp7Q00TXFRxEPhUw3WVb+JSM+m
LNv2BW7dYWhr244tKKs4YuXYTu061gSpCvJGGtJssLwpBt6thu9GqXIeft7i
YdpxRqVT9shyxK/Prs7OIM7PY1p3Yo41UpvLJHpYXwFLvtDuIM8a5+oXysRF
ifbDjfnCx9MUhG7PNA8rRZdR1o159vhWTYnCmWETm2+AfBf2oClm5sRjfWZ4
AwSW2ObNO7xUFv53nJB9AybDeDSV/0Hwtc2fckEI5H3PI/WdinrsnNKyK6O9
/AxDKHPo4j74k5dioMVI0pm7w6Js1OJOVZ5gDQdXP3pdr6COVQX2bPBmLG7b
Qp8mPaGXeHA2+bUve30BcqCFLUBYZoI0d6rJNzWly6+8Mad7xiFSj6VHW2P+
a1lqtDx+mxRpuweQP1XOkMr1fhoFMaFVix3s8P9m+q3cu+KKgl6EvT8RqJv6
HdAV+dVtsNHspS3EybK4ZirU8e8s3MIKUNfOPgeCHOhpHYyVZrwKuVahUmfH
/PRtG2FLMh5GKdONtXEPE2JVZpVhlGdnvn6fEjvelcOCCnKslmdF+t8FtgNm
PR/gji2JC1tIgBrCsPEfDUvPI93FEQZTvjzmvtbBfoHJYAG6VnwvIBX8IxOK
l3A+2F79zfvtscjAsCTtBMopNw0D9TPsfumxZjNHgXtoQSeZr3luPI8JtUYE
282bpZAAxRDnvndxDdYx3BvD/4/7DxmwVzI6xamszbQ3u2dLAZlaOL70urIg
JxC3hUE869oYkDYYxqa+eAvTbdFX7lTI28S1Z3NGi6tbxH7b0NeUfPxWHzTa
zExhVfWpoY1fp47R9aOR6b17jW6zDXrHIp0523vR/H1WiDOL9kylxpF6d1QC
QsexLoCIFjXCHXqW4sIs4OBnmOF+yc+PbETta3hhr1LcKCLnbUayCKz3dR07
KRseY6NhbGCQiXoB0TNaPSgEakWz2lK/I/x1JOGkjGbWfuAtjrDlIq32oIn0
Z1ZKj86yqkQtblFYgqFChrunTaarCU0GWO3iKKE/l5T1fc55LBiYDJgANIR3
hkPGzf9j34qUEJP7guoXMjparGXqhCEkBJjgCn8g1EU5RPBY1ArDABs065Uw
SPKcB0QzVooxCZWkHSuK+k4Vl+jTvEtxq68SchyufeqSsVZDNvFvQZO7rooM
5+x/OrufaKP9ypj2Pdb26GvtFcMvLcYfKJPCq8NzuKNUlGki2rIfe780JYlJ
AWZdWFP2OEXuLtXX40i5jVLn4NjMqTV7p/DV48QXKnBST/XF/i3f7kQWbx5I
kPnPzrbY6oM4zN4QjNGl7D1YXs5dNcq+IXbCDp+kIcp/CBtLMRs/tbuHWGlE
TWOOHpq4MHLUn0RScGzF+A29yIPMvayxf7qlMRGcRtKf5wMeMCtQ1gxDxEx8
HmJ2RhN2o8w+ltVmVr6ANg/DwYx9VMf0aTBZpvwwA9VfczXFz6ljmjwT/4vZ
Xl74Epr7DZtC1YjG7pWdLZFEDUMIwAZ5yhmm3NjuUASjoH3i91UHgtQik/dv
KKiK/uEHMVEsv3jR3jjkWXsCs0C+g0fYtuF8e02puKQCEDVnwx7pU+B3En/7
fqDs7CgPWgWBUZNVrFa4401bG0jU+pPEA8tmE/JSlCv2Ym0Kq2iY5J7oOsI7
o8lxGaTftdzCmwgdorgyWEZEkxIPXrHNbDcYeVp0ct9TLRXHh6rMyXPQy/V3
N6P/uL8ai5LxcsM7Eg2/Z05/w00Egzy5VEUsW1oF9ZDE4T6ToBVU7Y7Q8bPm
5owZHMDrlYh/bgaenNS8bVA86svh5OCe5fvvO7efugSwjk7WqvUybD3jhU7W
vyfvQD0RkW4hz6onopu591KFwYo1FJfnyAGSUsoRImTvnm+ZevQq6MgoUg/g
GJ0AM6/9lOC4EfKKNkFJS5K2xqUkpQ53RLqZlzxeHUa+6KQrkkAIkz7VddS5
sfYVJ/JRsDAx89q1Mi5hk3FRS8W6zKk+1u44rmDOc5hHx/4dtqxxiSloxZYZ
m11MxCHWEbOAoWJR2PR3/oP1agd0lfAIAU7XJmKgey0RZme15cHw53G01ok9
9Hwtfyyyhznbsv4c1VuTIymSuKAl7JzlqTrMumCY1elLtjGQegZgApja8OUo
S/cCLceJWW7S/mtJKfoR8Ly/rvCFpmB3/8UnaRyk1ttTI8wUObOyZjddroCZ
O2tpmWgr1SJjQPgiN/vHUnH64CvQZHc0Nt5GNw13nxNanuiHsShMNitu96DQ
z4fOKuvideQsoAWYpL1z/u/U9rGw2Y37J9KTnVtVLf65Kr8MjMXL2hMECWu+
RDSnrwfxiu2BPkm383scCeRFk7cypfB8bvRPyrch6iGEDFsWBl4Na0MwzaLb
kPaTE2cY1x70s1SvpUP8hPxO64saI3mQxDIiEW9fmBKkQW+MpYLUqyUtnyUQ
eDnerSSy8YW8ma8TAKliXF+1Vt4cZiIBF7Dw/RGl0QgDhSP/eMHL6QrP2XuE
zqc9XC5f3Ye0U6621TQmnKt1h9gzvh8abw00umEXhKwFqBZ46ELx/uG4S9iP
xjoWLFpcbAiysyZko8Qcd3VNvc5udXvd+MTxNpMN8svt1m8wmvGGcoTcMrtM
Lg1LvWxRvakL7CiaJgE8qZL8U4Gd2zpiAPFs6xGsvGon/Ep5/PfMR+JTp+Am
r4/kDno7Bg8/C1YuQ82FhDNujU0bC75Ef7Ks5hMtJKYWrV1oprkPrNfAzXsr
M0LfMBRZSuHbkA/A0RLu4rh60kqzFsIG2rMefb8+/H+yTN7zlZzbpdJZ2ohG
67z6VvlW0DE8UTPYixJWzl36frEHsLJIh+t1cUQD0f2Yny2pJFnfJLdRPkGf
g7cLoNipWFyzYMBCMLHa6/GKPHkljfHe+2wbDI4KrMMjNLf99XUpg2b03Cl6
qvov08gf2v9eFAZL4pYmlOnR4zJGwa8rjfnqTH/goLocPwMKl4/qPQvsbnu6
vXzh3MgiL2JZdfpKygqn+mNNb4efooRuzWjsPDG7ls0t74Y4uyOG6C/53bXO
O8g3Lk3WhXWEtePakQcT+zmWeYRE9q87HIZBzMR1zuKm/oL8R4An96lKURmj
LQooyP0OGwWlgYGfjIPNN3N6KEYTzy4Svk4sH6l1cwp9trAH7C5VVddptGR4
STx8xNkcbUqY4nk0FB+xL+vd8QyuIDbgTpnAOXAZngPc1HvrJgYYrJfUc230
6cY68nrdiQypG1zlG0Mb0/3CRw82VTXrit3YZGsVG91okofX29Cl3STnYSIv
4VYemOWZkidYIpImlyHsINMWBB5AEzUp2NTf09LN1XXY897GUXBC+QZlGNjj
/LmMlTFdVVfSgv3FS87QQIy8XTYUOcwy8l3wTkzyllMyEktAQFM51OUYDNKa
wfVFOaeLPuYZimUDG0l/HJQcctIMRPYZWs54PcSVDI4MwdF7ZniQcGsdz8kf
GogZEpgVSvFixmJYIz9hf8egIZf9489ryb0cU2mR2Jd2RBpqm+ST4uscNzBx
sPigfLs0FVR0ieQp6dLOm5Dr1R0O7SI8t7cnHgiUCpZl/5dopPMBcyg+XdRr
QolU9XvWtk9xonDhzqMPZ5EPPhoUZKayj1YW419AuuhmYgvH3envcA1r9Ps1
6QG9pb6ydiGvwXq95MvCd5I8+McQpYnKgcnAbalrjYirXFX/l+VJ6yAD8oF4
wzNnxiqvBKcN0yEovK489iiSshgVUkv6QaffgHzTgQollS+kFQ3GWTDc4bzN
HyGihdzXFxK89yCl+Jk+MSQZC+7+EkO/rkE7BnfeJ8mUu9XguV/iFK4W8+0I
Fkob0IIeQjoBf2HPIv11mz8p9ip+9mZiriKQqL44l8z5MyaHt238erda0uNT
nxVU93eag0nYoiYL9/iPyXfacfjq78Jttgo+DgX0Et0M7CoQ9ixUUFu/L1cG
D16rXfINcoYxwoJd8hGTBjmYDOplZ7ITaCWqXjatdlicl0EQriCslTAel3G4
+0m459pfjN9cY6TelPPDgJPrl+w4Db9KQFgLij6+VTOAu19OS5LTh6xXHjVp
KLgV1+KuuFt33ConKBCVfhMS8v7obx2PVCGgvgVL/6WQouAkrC99+X7V5sev
WDsWNYNELWo5s7o9CkL22vRyuf40njFve7QofO0084VOq9Tpv5IqP7l3NKFn
X4o+n8yCtmyYOSk9V16a4QbWB1NSy5cwvDy3UjfYSKAgvdwEPoDaKCVOgoYz
kRwi6TTKbmpM5vEJgD8VXKWca7silp/KtXwqxKaNh77l7Ww0/LGTYY/z0BoE
k/cUKr1m17v4jyuYsYnGstfjrmTeXzV0PObTJ3mwnThirx8aySGKYzYRh6lh
xAa6xXYEHtVOzdbVlgnnRJX4cUpUWrHMDbGuXg8JvZFGCR6FnvaHCafM7Rp/
FRvpruqW8xrModtvdVKQwrGYcr4NrgaDRkzBKbGel133KcoMHftAHycdol1Q
TEQfySuHI+FQbzMTZNafRzSSWvOx691Pht3kC3M1LLOdzkEphAzby11LhAUD
Yh/OR8zCems8JzUedrKqnLTBW67wb01pUud1t605kjDshAJ9wDxORjdeFy7F
4RzOB1gyYeGR1WOhe3dkbVqXjzo5vGJjfbRz2eWne6e/VSMTculge43kfEVa
LbB0YCDxWX238BR6Qoh4OpZY8MOHSi6m3Bzwub3ij3naokO8Oi7tH5Gl5S63
SHaXVceTuS3Bw+jdevOv1Y4vgwllL0F9q5gKw+rU00AYyGLN19FeE3mR2J65
qE/xR8SqJqu7RhKLpVrS9RZUbRe9gBFRaLPSBnMOPJJh4voiCamI3HUfOEMP
Xf2dCRihgl1pybgmVSCsJjmYFOgOhnkNC5hjDoajLg/het6dm381zew3mtNh
yXzBM9H50BGPXByxRR1YdAa/zLbk/fSICLIz4OPH26Pvx2TK4Aj4p/MGpl8E
wl9R31ytUYgvQzKXdqeLa+DbXmXIhyaMnOadUfq7i8ejk4Pv7D/Vh7fQltOP
EbdkK1D+iejYfWcrk6VrTaYtnFMhZET1KKh/9qDxZSR+Jncx5ZMz+HfwEf1e
rXfS21ll66trsoqv1uxjooZYwjJJw3Ul3zz8ex69rqaaJ8F9Anbnm/FGUMl+
q1+9CoTuSPh44prabUXsxzZzOVQgpgwETIEYoYLylZKRlV+5/XQR+xsNSQzV
bPi1TA/eLEv/CAS8lpgVnHLk8I/7cVBIPyEtlBLMHsqqPz+4Xi0cd/VakUwc
TG/z4c0G+DCeSTpk4jyjw30MX01/OjYb0RRRfw+Cy7imcKilxkd44TZQqK9G
NtXDP4eQM8l5pTe0EGn/G1gCMJgU50qrcYm90QgDFZYDp44ZKPfkHkvgQ9s4
cKDt1c8Gbswdt7WnO1j68dW607uBvbNj9k1SE88OdzQgsWeGVA8wkX5vD4Jr
sWREFmQztGF8UAiYEu6cSJQszvjy61b2DvaetF+M9DRhn+kvn4dU7Xhe2UBb
/cRalwf2h9ZbcxrYTHXCzJnFZC093u8R6pXaBHfPYUUIfR0SXiazcFoix5+F
jTzpziDMDNJ58dEqTkvQIKroHIatqbkPThLqJVLC+6C7d+Ih8s+2dtB/OvwQ
4DgaJpV6cXBeC9e7AvQZKEHzAjHnoZMtqlZ0bMVnUb9VFJ5vdRmW08hzGqOz
4cJtf/Ax+X/Mb/3SFvfk04ZLwOeEv24N98Kk9/+a5ZrCPE1AczvdoSc9GDGy
EFH9HFMV892B0KtBEMht2nNxerPRx/kzTZQ7tIcBObKMSCJJwDLvjciUZlSe
kPOExCCWNkQYNjFSMup7fAjADWL4YCSRiGmDOE3BlW048/U4R53AjbQfTHBJ
WjXVvPjiNPebvUiRzy7cCqkUOBnWrUujVyzX4lBYKIbPcV3cd6dcDUt1ZnBY
/BwB05Mvb4YB1b2AOnOSbocz4ZN78zhfDzN5xOpwBPx4XXtQbChUTPnqqswz
3VSCjDfd9NUAm/FtPsLId+F6MVOGSGK4Ne7GPm2XDOu4eRZllYfaNyPnS4YO
8W7QGYSHSdad3ZhP80rNVYF3IvrMcQzMg8eud7CWP8n3vEeogufNYtjLC1R4
GKUwCokNN8z5hdJJLnEKfsNHMLUxu9i2bHBCUw0aY4LWXHNkx282Tnmd4JgY
UQ9Vg/WFC9s4Fbu71qysswd+u4LeaSin0Cq0rLq38sWX/Fuja+M+ELIsrjw3
WvgX3UY0Qh9PXBytyx8myFFZx4UUJu4Sqo7Pj6y2aeJWWPdfrUt/b7iSLvn2
8aYbt7ih19bOagHsFiGuWIPeUhekfjhz6GEj9oKH0vbzlFgmzIPnc4AfBeU2
GgZL56gJr+KQ6HVU9sEsw301C0VINxLCKO6NErGz0EelX2ponTHz0z6+TrRS
HYk7dQGR3SOOfeYgAi18GIdhivrfnXUh5V/VoXp/HFBgHDesB2+gX7jZPWks
3D3sKBLjBAUTk90M5/6msb6h34kofob6W/YiP/o7nhtBQ5RO3WFyiNK0ENcy
BnWxTidhAe9eCKce+adl4IS3BRxUqg4JaUCKjP24WwFk5FVbRDpDnc/1RhD8
lRxHbnRp9FFX/RlEgbeNPmPix6PQVYmvrx+IWD+coV3e6SiF+AulpOPWzJrO
fxYpyyHhZPNvDiAzYvcslR0+tVnpZ6zA6UkMkZ0vFcQm7G9oFu/66we9AY3e
Xib562RDStZt01vEiQFWMr0dcQszr4K29t/iazHEs4Bam1rBN/FRFimmCdQ5
zzhpAe5NEbbjRVbTwluw/t26UlmbVi+PG9sDbwlard0VxMrsi5L9j7cSiqDm
OzJndK8R42fRynuZNfC535XpljJ5W6DCQHK0j8sEQgFeTdptbZe8XX+wd7sk
GO0EhMv+QqBCvuK+qPLh1F/AvPa+GPcRgXBqdvULAMKkvQhbSrAXEjM22QbK
y4PbFWrxEoE2phPxjXEtEsUNX+tJ+SUB2ZSuY5L1ksdyhRQqdW+Z8GnnLRQS
Hw+4WqkvAr+ci9JDOrX+5kYwEBnUaezroDIATF5CXQwCVfFCf4x/zZA1tBuS
h0/GLem/nx5J52wp8BibMdA3vBMiJasbT/qol24N8xy13ZzMnPTK+Am6LtxF
6jqGdHYEVM9sIBe4qoX+mXF2csmwfo9vLTCTR8lu+p9JmaFsNwDLrGQKBfLO
6pK0ZNqVsbTYwHc1jo3psA6cQ6ZTwxL0ioIU2/vyVnY/mkMBKu4j+r0Ys0Hw
fCMKlVSTDdDlmTskQyB0vF+7/Ai+u2cpvYMAuaZVjukgRYQ1VoLnCMmCAds/
2bDiOG+yewNgzKcb5S9HqOQ7IeV00cJdcpQWklvq+g1lBWelC6roucIOl0op
FZSAG8DtADhA2whCs0yrINkh9IQQ8NQnPuhfRz3tKB4052y/JF/xGDNydN79
PxT7sFxCEHTdEpEDq0GQmnZTlTL+JGTPn+z4MejUlWXoWWzNh+dR8wNLuFKW
J/3sS5xkKXs9zFAjqA2/QL1/8i+o3ywa0Tm6H7qHdCc5qSh/ccOKUu0Xkjqi
eNQblObrSBZ09mOYnk5HHnkESBSuqGQjOpFXcSkBSsLZjYIFp44gP+a+pQQk
2HY1e888R5Zzg8Jb3spLZUdlYXZefuQp2rKkxrg78sLdI66pXjcR2pu7lA2r
nZHRq5eusqu/GiWtlwAdqfkjBil9320gWIJaoJ7m33UhhkRF8SIW2TwETYsS
1AntxZRP4Z46Gcp286JZ9c1HX0Yqk6yhbimGAP1PaT0Rlo25YFsu6qtZ9HOA
noBxtl1gB3XSU0kEuqo3VcE47GG58uCP5X26cyRE+MZKDJKRaGYgGC1K7v3M
gR6bj2bJcnwkCUjXSgwtPCB8W5z88NRlNk8bqUdShd8e4vsEmqOHRwlpdPEe
hYy+pRC1I5+fAdtwWD2lY2dGQJeh4mXRZCzfG+a55tZ52nlo2/wV44XfGzFK
i7W1iezLIaxiFOL6lsBzupCpq32mbmO7sD4gMu6h1xoJNMEy82DlKv0oHJNz
LDRuvM7F20qyWJO7ZgOOqyezQszZ6W62Axu+U5du1ICGhFgzx24Ns9q0GtE/
34Z5To6EGJYMT07pAwJ+pJCmmLY0dpeJ2I0An2WAQG3h8EBTdbgp31BJF4Oo
CJ4WeqUGyPZVFLZAssc8wOqkahXTDPbg0h6n1ZP9edsVVPA2MsIkSIJjo/cR
MfrJGTxo/i8YzNU0zU4xR7FiQ6yIGy/8LXnZZW7NOT5iZydNLPGq8MOZk+SP
pO0YBBtf+eMc/a2FEmM0lOl6VLVJbuOjOHbUIz1VJ/PTQb/jVzl+dn2iDG3f
JTbBB/bKHKERz0I1xkCDBZLt4t+GDUql/l/E7w8SXJrYQ+t2/gSpngtyLsKd
cRE0seBTS5ww2HtHm1QC4Zaw61QyPthHMShL9mM3ek5dJOXCNVeC4L0Yp2tn
+IkvdaJ7TCyv9ZdAqEDBHIKzhaHF1U99IZS12w0QD00v2YCsy9hjZRBfRfzw
QjECaokh1lxqzZfS5HsgzJzLOL7lSIkzI0Euj7hATB3JNrIbISkfnxU56Z76
JEfSh2raKCiTMvOaYquz4bGV1gKS35C/grXwcSs57wf+5UDQieG9ctCAVLlE
pH3l1j9W6X5Pr3hMBZ0j9Do3hy1yen3OYPxcInw9AWBM3QMWAR4oc7iIq+jZ
Lf/84HNJa2wUTuXFkW1sHykY7LesQn73WjykFN0FmhQWFyZ5uZsppge89EnZ
8mFEnfRtm+NvGeEjywyPhgUGSuatTxAic+vp8o0cDOyI3uxRU7p/q0jZzS8f
lU1r6wPoZc/SYuyXdSXB37RbamveqEFujnTvuIFVR/mSLgKuWPWqv9zvysop
dgG0uk7hiWyQjNw9bFy/Fz81mt1UekAIWIEHpKKuYgvdschjoLUSbOtwQulE
9g1yYNEuVfkPC5veU52xYRoYx8eJUKwl3TquF1zQzH00majgYp751nmmaBmY
uQq2aS3z7KqwMT78ovbA9ZD6f5bBqat853W6DxIw1pxmudIBTpSUC27UjtZu
EMCfmCBB0I0EPD8QQdANRMxzyi3WiYn5alJvHmwv0a1ALYjdF2LHocWEmmwA
xFILyn7lxCQW4JFsDP2KREEbQxNA+2kvzz4sn6s1FMkoABB2SZcRC1nCikYN
1eiYgkooMRI5RogdbaeSoHbm7J67NvU9gzAAumOMY8wsU0BtE6wMimpbS1YN
7mjbT3wqMg9LniV/+7C2I1GWPRpTAiayzFW35eFYUJHsRZdBqKOPM0S8rz2W
yAB9C1FB9RNt71KCap/ukxi1qlcHUzZ4G5F2ZBT53mjC+0oYClVteTtuKeF9
wis9xbqfj/T4x7Ro+GfAfoMwqi0Cl0Cmt9ShfJfSlotk2LH+08AzaYzp18xQ
M8axOXeahQt360kbNl3AOVu2z4PkMztIPib2FY9mTE260NtBcYKTlxxzX0Zw
/IinOciGW1HB6nQQhhOULJ6fjUAcC6N3JR/TQv/LQifn5Khf9FhSP1RrJebX
0KYNHwLVbwrdUT6HywZ7sj8kkWd7yL0GvLMZqDUZHYlXesA1H06zBs9K1tjX
broEn0QRofUjol6o4OaR8d4/I+1zfwEQvz4vpKEwc9E7Eqr3ddru5B30ZOkg
nqllXh64cuP3cKEL7YUJ4JwAsrxGp71TKVn6elTtHlNI9nUoLsBDg6cpbxrV
4ltzbJ30eo193cpLV11wrVtI7qwus7f+6AFhSzhJjqwdBWIE7N2wkFBSpAVc
kXA7OCQ5YFa9YjpzS7idcJXlYH/wxldCGEH2yeQLUK3E5Amc4vEEw8YOwb+V
D+ro7Xy2Jiu6Oe+AaKjxpvyhn2AkUHqi7l4Cs/0nvGL/cnL7QYRLEcqNl0jq
veko7CBsa/i7G+kOvoSYxUhurgZoNk3YF0z0bpRqsP//fZTYNA5/76AXEYSP
bV1mx31SKatlJVE7M+XG4cVomvlyMoJqRJxnX32NurcCrlVnOKIUNZuljlhf
2bXZbUM8Nrg3Br1jOgte8ucD5FnaxD+WDHClCEIxORIfcI5v+b+QiBjSczSf
w63QogH0e0LHpSjlx7yT7nhQEHS0BqDHdZI/Ni6whpLdBEBmGXREzFBwEHJE
bCjYiXNhAFlgJjCIbHbJWgiHeO824yfgo5wFOlRqa4EZ8eHK3ygveEJIOz6Y
C0ZfkYqg3rmzyfCcZMAVFjNjXpzDDFjLNPcq71dJvLwokgPqeZJq5ZPdbHX+
Hpo5QKAVOVPvDQw8b5Bq7Qvow1ye9QqK1C9i4/xFpDUhqy23+q8PdUVNEKIv
CfymYu/Fit8epZoVf8gyoejoYfhlQhdmb5wrXtOxEZjcSvVN+zAp8CkWyGS1
YsKv2FhAhPVZZEyAE/559tkl0tmprmOGUrCWXlGZiaNIXQfz+eK/fYOD1Hhp
U3Ett0NcH2vz02gFC6+1mlwIzzZ+m2fjaYdHJ06rfeJzocf89C9d/TKbVnfW
WSOv4/FDqQ5klyKOJFSpvPQf7lF3AVxTOrNe/xZ/rE1Uub3QGDCtWtRxK0yI
ayxE5pP9Db7j3vw983u0L7bQtK4jkRXEeEzS/F7W0L1twClpE88qwfFVgmCB
oq+XzeF1x/VO1LHdYO8LGyP7yhzJ2D3ZfmjYEJBHUu1xXx0GeFzUNdZ+2aRO
c/sxT7CHcgPvZWt9oMegkLgYoMLsG711y4tTBhjFV8Kmhxl9wdfaocxmnFuH
1BF7hAlObDGITXblV7fU33a//3OgVzKcz5aQdOjhbMqk8SyiFO+1TXdUAKWd
BveKwNiESQWeGwal0VZyvlutYHRhqiYXYiucbh4oLvzPBJ66mk5Z5ivhQbLU
FJeqh/44hlEh6I56AlJLUZzkrnhoC3iNBmaOAkM5HIXhBVxbTKDfPEOWqCMX
GIHDr8nbWj5TE47NjsUycUyjHEKLLWPLM5CbriTv4LgH2XcbQZfKlhwKL3Ro
Lv2Fc0+OXgqX2SA06hJoqvcubwspydlczGMiOlIpth6OCa4mOYo3rFI1PYMD
xgm0aAa7gS/H0ffRIbmqN0XB+EVRR2rxT076mWndJi22rx35Ej7FN3Hg6xwY
7Izz7SMNDiFOOi1PNgtA1UyJQWwC1t8wtkpg5q6OxPDmx52acCuPMzeoV1Cy
OJ7BlZkczEZEWgTgPFaxHXhqq1nyDoooSUCb7vCDjWPzgZuNSaBbol5ntB8C
E7wBGpwcg4UvBZB86ovfGhi+ucNSyF8yFJaqjS0zsJI+niwd40IzL7KGnLP8
kTqtZ4dfgdA44GaSQNXQ92IPGJOYrXgdqqraCAbV8l2WXTJu2SmfW92Ppzi1
Gq5KZp3nZtkJMilkmi1s4XA5OVVFBd+jGRXaqOUKYb1Lkh+f3oFbLt9MGOza
4Z3M2Zsa35rbuOBmCUlP8dDQZBwOWp3dKNeUY6BTYvs2Z+j7eptgdm++YcMR
e3peoLRhahBzLZ5p87foHo8vr8lQ9vLgselwd88e3v55LZJ2UZCRPQIROzb1
t9OtWSlYFMp2L2nYuY9FyaSAjvjfoR09Z4P5qsvFtB2ZY0PH0Ri/AitthTgb
m47v6lBUbnR30owhtvK3z8yzrfUPAFCtND9eZlQkRZAFhZwbQaY6pjpM6kiF
j+6HMbQ+8qgIhDEIA6SWgUJlWatd4rSP5lFdSxyHl2RaASazC9kQorTyP+NC
XA/1Kk+VLpqu36mM78m2y2Sr+xBqtvoVybejc4dQ1BxnZay8O7mU4/00Zzcc
GE72vCHwohsn6gqt1izeLkMfmITUUrhJOv/5dOVz3pHa85lHEYE7HSf1yrzT
k+U6cIuXJMK/JwOCr1fZ/zqGucJmX+QJlEQCdc3UIgHqRn15dwina3s/+nFL
Q5B6agxF4Qa3YswvsQiLb3g/TXQF9P9YI74AUoHHTf7BNd17ifaLlswgpTWr
CfWG9EuDYvZPfbTPLDy4B39muGQfK0Tt5e3NH1eTROef2OFZU1QR2QHTpzM1
DVa63BzTZqu+HgozP58pfLwlUw4EIEKRkUPaXz5VhHLt8I1Bzx1K2cv8h6vZ
LeKAfG89RFLzfP8gyqsVqU3Mvca2zj6hAOzJC4dZR5lLmdsTPzby9aDP8KUJ
CZVqnzCwSzxKVecnco0CE1YRyX2AOHi+77gOm+wcJefYCgNEt0umlpnIgXZa
oThSFO0sTELY7yRKvGzO++LYNfIc2hgZp08fdc99dA3KplKPDrIz2QOXi83+
CBwv4JwlwgeYSiZXgN685A7YtzGwYdXdTiI1vOfnJqbnrb2bSQOfVEW1nswM
jk944zVR4RUwiSjH8o/dKFkfadrG+fwjyWr6lPHDzqbkMP1w2P/9GV6RCuG0
Bi0/H9vTl9zqsDtfODZWVU8/WdWOJ22Lj954E61dF59u8bl+x9nDiSOAoWE/
D099zarHbZfP4VXTZPYuaePheZ1OJQNaEBfeWNLmOBpEC2U0IsqY+dqLzrCO
fQvd1WvflGSkQ77RZ70fdls+FF+sLdoDWlaDVuEOJ9GDBbJv+5+T4Sg5iBFe
fLjvLfQkGboVhut5GCtF+cQfhuFuaJ0iIVzXM+NIn+/Qm1RCYO2lB/zYCCzZ
EzF/oNturmJj52BmzWPyu1AmQHU2Nsw8h/hisb7PBVrxdK16/puUCnhWQ2uw
XYuOjK1666ztltvvpRXLx1eMeM1TISDL3T+E497DmszIgSX1Xj/XKB+ECVT/
mHUVGLuqHKLCVaMzyQqOOerpVBqyllORYju26y95Ju4qjGgRJJtz6gJ09Ub6
yT6qdN5cekn7FvU9kbDcNTe3nU/ndZzSJiuiM7BmgEBZFr2yXgFUjA2kT9tC
nmo1MErpFmdPQAUZZQNKPIRikgzlmtb2gHS+MT4LC2UsMEUsjMn9NV9Shu5p
rRW8TQ3vFyCzh6oWT28x1X31dhR/Q1//JQKaL7Xws8dNKE9YvoP0SU4xkp3h
+79v0jUJKbqYKJgVcZ4Kj/BzRS7gPqbrUv7ZRNcDczd3BdGFJe1eYBw0F/wy
qNrO9UeFBjuxBkedTimQDw2o2pZIHLMrFNhgu6CmNpUx2lGdq4W+qgzRJUmJ
VLtgYfzUwRYbLTeuh7x7TJZeivx204h0TucHvikMaBwaVTxzrfjJBMQP+JJT
fcZ04ax1xR4XT8FYvkjqx7ZEbWcB0puixAj1SkDQLpiBiPUyH95XoXrNv/wF
usLYR+F2PRZeVJZUnMLb00mkE3LbHZ43M+0/FT7tf2ewUdCxR3ZqAr5BgUrf
3YmBZKC0z2FVc1eSiS3t6i1dD//8OSldPj/vGjgoNKPMzPmoqyDzMQQDK1Kw
zcxBMLzu+QQdRn/VhYodz0FcVkNEC1jHcl8Pz8yYSZE1FdBC2nQjTrVRXGsw
sBtzYCKe4JoHGrer/4xewOMv//9vLl1TChYe1gvOhgWL9dix7Y7zgFYQkcFj
80vBOnNf333SwN7gZvmXVIzffM7Vfztzb/VVZ6D1nJ6YdV9EoiKK/ajYhLyJ
lZOPQRd2D36WbLQfkHTC/uEoEt+w4Hlm0i+k+8ELjv+PHTSl/ATRSVlja92d
OGn3WFj7vGzuLEOjWuOMZSI+krzy+ZcoVl17frXs4e7sygugjVDu0lzxp/pU
2CUHH8+RUF8/dpABrOhSgGj3zLHVarJ7qhts2fLLZDvFnL3o0ByATb44thC3
/xRuWQo/Pq5VKsoPl/sVxO/zgDHw5i02yDN0tu5QS2Lk8E981zJ3ooyYt69n
UAaJ6SY5ivLajAYJs20oBYZlrAOzrF/P0pvXUJf8DQhMY2cPjPN6HxAPYBMg
YtKQkvd9IfG/qh7WJNCuWxllIKmmCb+uy1szAlCY4xsZP8DW2zrSUmy1uel5
qCGpv0dPP7/yLhVTazRfIWUmuF8leu989v2gdvgT8xW2VNp3sKqlFuJlGr0N
i7EC5RDMiTIEySutdiETNbZ4IQexHsptzODo8uGPwGw7gZZS/xDn84pEs6rt
pyTyN5em9ZFU4hG8EXQpT9TeeDiS+QKMIrP//sMbrFKnQ9Q6VOK3CIotttd3
nV23e5Zj3wfrv3f6Ow4ZLBuUgONU5KVurlFoInyZ3yLB6K5xTrWtpxoDf2us
OGvSjOF5vyiwNi05jV94OMyTn4LvpIrBXD88DSBaZoIrh+Lgm2wvwDX9AlcK
zC/EFCkCSkY8THhc86WgX+Vf8GhggDbrbEzaH5TisfyRH5XD7kqQhGp81vx+
9SpbqWbKV2kSre2G1IAFgVS1i7VB+xOuRnnyz1uINyETMub73zNGWkG3D+sK
se5wnXXkqDF+tJ/Qpf/GJDLya9sIrXOaXbaeRkbklNg+coKyR9K/swFt5u5v
ITD3Et5AYhmf5crz1PT5M0/id60vMJdOu6YfnD2CS2PPoji53YqeUSOvW/N1
TQBQ6vDdPPZyszpaZEDSUO3bR/+r2i4oN8KGk72HZpTqTQVxGwdZCIOCGQBE
V57u/Ncp+7rx4YPAsDe7ll31VpjjQoW57ZfH7xpu1d+LZ9am0sGbjsi87mgJ
CeWAkwQoqP66fifNV7f/PuqiXE2EyKKvdkMuaOf64Dm/0IimUO9FD8B0aaet
ZUQs+LIc3uM6i9U4xoETgQuebe1CkMdQVo1uR5xAku+EuEtoqSo7unlYfiSy
bGewzED+lH8Ty2tO31i3NC9JezAVfN247gltbm6mKdouDwuYGNArVZs6roMz
6CkU1OHXkIdCvboSBgon/jVDtiXlC8g2h3Bew2Xqx8jn+vpmpY7WayE2/gOY
2B1iNu7APu5Shy1OEEdsVKXmfJtH1MpUFKqgOq4oqhipe4JWn+Bjhd5qZOjf
Ch9lPsIN6m6dri2+jF6TxC5BKqYHkBGHv/2E5gvs6qIAQxvDRVuniL482e6O
3KOTGFyCsTE38Olv2bWj5lf0FOpRYP1te8x+mqUklvPpKo2wYYuTNzN2Ply6
jat5bDpcEb/VYzGzfgsnJDQ4iaGomz0n7QkH/VoI6RhNCQ26LHLUF+rKna0e
d1pGc7mkBFOaNvOORksaqsSFoWhtelmT+67rg11cD+e3jAbZyZYSu62x9CtI
BTwBQf1t7jwOY+yTLfJoK1/UzNUyANn7p3PlP9LIzsDGDm6jfDEiTU+/TPRW
qUKFxPTDGVDRce6hn8T1fsRqIMkSqAs51OxcPuG/X9sn5nYwiwlppa4+PcjF
yq8bg3I9s31YjMp1PHNduY4b7iJrhMSGGwaMst93lckF/QxqsxPMb+3fGEbX
rkONuFwhdvwxB6k3mhOFKomuQYerYLyHBiiyi75+jqS7f2pFwn8XngC0WvLT
np9/OQmcseVYzszchY/l+9kJX141+7sU9NOGtpWoHLPhbzXKoL5YrfubXFUa
q7mJ5SLcN176/F1w5QLx119rk9K3ht7MxRDXb1FwXj5123Uj4bXFiYLxGrPl
CAUBTp6T1qYagSt0+baqdAc1l414nrOWjk/tiC2PpbYquEQL9zLUkBBEC0m+
eksxckMCRJmasP1/6pYI3ArrFAuNE3Q1QRWSFc6Ap+b0FmLbQO5EMYitd2LT
6NIQOYvbv8Jcum+YvXZ4qHiBX4c0dGE6Rtgt1QEf0h5FalAw/1StasvIuUGp
73oRejkFTAIdlx0dpefyVN7N2NbcY2tL0ceoIb3bAkfwX0zqMn7rBMDl2Cjv
Jg0C3ffZLM14r4GM1nO2jvOPgh9TaYDki4EpvS/JvJanHOUfSrXlNOVhvuc0
9njSXgat95xbKVmWW1eGwhN7HQ85KhhCx48aDiRlMwOh/NXYHphewQUmHn/5
pbTRJV5YaPTGgomOu0foGAAbaFt58fwcyH5eGG1FUebtLgH8l5m5+59kUL28
8dPGjhOOcYgTIBm6BO39hCRiM2WsQdesjNyH2I8zWM2YFrk0CWz9wbWoUFGi
WTd5FJjOVFe9Dkj6EF32vg2oEEcEy0V/Hwa2Tktq5ZZLub6o6Jy8sZn0ilY8
FyEzFd423lkY2Z9FmEBNbqIhhusWCZ/C+sCltt769XZW7xXP8dISEDQGCNTh
ddbhTBTqRPB1aJgV1W8qTUl/vyncNlh4SCXlpAUhCs/VODx8eucJ4LY0xNxn
cBZSwXjK8ZzTXufxhYwq5LRt+rFgA35UJtzU+Y3p0/vzyd/NytxSA2QDzVYp
9yJPs20SUxt3ptpo1BQB//Y6TkUCFNjpyMFW4PqcznCtOiPHa9y/Kyt0brRv
vX8jnn3mRt1YVCxnW7PojAikOdUNuqLiYQ+chajnlGVy4AZE/24v0wO1R0Gi
q6ax5AkB44hYBuHYWr10g/iM6BKpqpppi07R6q7sYn1dTNqae5YxJDffEwSu
iEg3plcK43TyqzUoPtpN1mvreX/SAVt3j0x7S4kMmP4gLR5JZsCDzdGo49qx
lOmwiRBC9BRC4+vxhQtjuRzJnecQFAxa4nx5W32D+RZmNfVDR0+RPNGwcylM
Kfo/7EIPipPZBT0RIu/1/IycHhp7jmwTZNX7V3CejGOAWBSvw6fq9e4K/LPr
WfEGgxP/mhOeI3opikf1uy2LjB6/7fw0o768KtPfw+pmSpcMPKtcSkmSmPTv
jEhqpWvFCIsE79QIPxgxLgVriy7Vb6BwMPA7ozSA7NsMB89qbtdlVI4zHihy
pZ4Dn3q13tIoB4wLvY4NyEEGIfHp5a6BhPQaU/SB0Sn+AwnhIDoDRrkEaP8g
k/J0i+FX6A+HFUkcKjyperC4kgAqKJ4r8jySFw41W0raZR9u2K8OBlBZZOd3
U3vCvoTLfczcGoJOuw8bbJ3AMrB4Yl1xPZYWdcEhnkjMRQBV5xl+nHC7PMwV
yD4b6+lx9HxXnCw7+XBvezw3i/7nUrJ/5IEn4T5MyRGTRLsl4276Gjnha06t
i2DT0iuUIgf4NPwdBr+uuM5e1MHJaE2CefPLMT9H++uSmaMxPUdqmhvRsfcy
rgAgwgI4RRFj5K+d9yBIF1BPZS/9/P77bYjuUGvV1e9CI7sIiR+Y8EF2bniV
pfhZV58sdh5puPcG+Xu6JYv7+I3B/68utvThP852LZHFh3kuah/0h+dkJR58
pRJgv2QeoUmSZkUpxG7OhfEmlfTQ54sRsKzPTnKsbqfMakPKm+Iqn/+E2N0m
xXEZT5umOxsWheUMJkIGr8j7ENRcz7d67tf0BObHRL+FJN8wLXO+dPINte0t
3uVEbSfWN+SQjghH9yWf/mj+4GXVB3P9Pmq9AwpWUWC2a6sCU071RNP4vfU5
V7XFP7F9pSFiN2KaMlD+RKLdIlLftQeZhwRLH3IhXR6aXEqe3LfGGz9yBexA
ddIj+nT/ParM59OS2fEYkePT2qxcSyxPUnz+cUg7yvRAErHkMhhVQZbpblSA
QFC+nQzzfUmkcHyVZiARSpJmXgihgDCIRWsBwhXnuMT08g4dD712bsn1/xQi
NlNhXHnVRQHW33qp9Sx0ONGb8wEA0qqTwdgpOLr/IqauimUN9Frs394VL3P9
QDtTqLkBfcVwmShS0PSlDeotzhTfbXvQNZgQytkV66I+0MACr2qMzNxjXcHt
tX6MUgYKhvAxXGzPXY71fb3U9H+brqM4RccEG9Fae+HAuK/JIGwSjn+8jaY9
kicVExQXCRiWrMGgSWgQvuFgyHrcec1/VZctg8JbQWCOU7lFjYtH+uwPk0CD
tkdPxyowC0ADY2rYLUJDRye4y+1tbMjTRHhm4HQSKSkcdxU4KUnViB8U5aMD
F/HdxYU6CPR1UOnh4omnlXyZN1vYSaK0ki28+mtJnpG/sOiZiVCG8iswxwg6
WYkWhjWdKVKCcTRLcxug3ESeMAdGY0w1TuD5P5EE+zG5kCgQLS6NfBMtuAn6
QLlpQYcbqNELagaytq/zGLozMAXQk5+YZuxl3AEUJ5Q+JCbsCLP4xgNbRpzX
n8DQsTWYz17/NyogMYJeLvDhY98GOD95l0nzBErhMSzIoR14l8hTnw5qPizr
Hee/PznedNd18ZCOsDk1xiuBGbONZAfTulpNazw11L2UdOcCV9RQzCVduk1i
l7GBmgiGuiK9HsfhVUP+2cUbraqadc8DEbXl3uB5QHm5rb7Tg8LXJ3hnhIY6
ce77l6H5/ZXnJE0eGP49S3AwkRHemceqnT2cWti30J6zJQCjg4bfMzP0ZiDu
Tl61rzrnsrDG7WdIshH0TWk0kUQMLl6NA3nIrBOyMq8FHObLyH/37mwlE2V9
P2ziw3tra1oXt1K7m9cgF4CBYoKfQb0zyNZU+WDYiUuOhoFwWxMxexHIijeW
055rxW3m613pGkP3H2PckF40OQ7c1FtiJy16vdlTWOBZmcjPuwZ7k620UCaG
x3DDNGsu9EWj7RW7JEITfR0WlOw4aGON0RFsXoa7RlOMsJCz8cl+WC+7fS2u
deySP1rU6Nprc9j54ncZbVAF+4nnn4MXSYmd45SMM5JzZEoIXydic0KJktIN
KoyiyjY1R/7QvxLripdGbWor/KvW1IMcyvgsTjcFi0RmJrTusP5yEbR3bx/J
75ekzzIcWoELynvEaS2RMG5ywnlBT7Vx6pmrYC9615E8qVvgYl7ojIZlAmma
q50LmKRw/XOTBWP9vBLG2Oiq+CExyfSsBiQ1bd5vLob7WhoibwVVpjtDKKMR
AwseDiAtRLR8E1UGzqxMB4LmA9LesIx+NPlQqFNN6UY92H7YRo0ncbNWwUQv
Vsqtq2vhPdMGAtYWAzX9d2SmFUWR2BTuV+qRN+zOFzvOSuc6KOb7f0dGUPDZ
UBuW9ZW0ijLDgZ1AqrNPlncT6+zTmh0ICSBZuP4cr99G4Vkr6FsS0R4Hq23m
s8fdg6j0NWKx0reqARFCrYll/Bnz+VAr4y2hx30afQaR8gMfjL5RMLKJXtSY
daUvNclr9uUvt9VCSeKoWy0+Eb+42vXLp/25E7CFHiiXUz1iX8ONHXnrg2Vk
taou31rgCqRma3+liBQFTRmQUadaxRic7j5K3KAiLd8FyPFNdbyLQFVeoHd/
TLng7NIljITaJ2dDnE2PQ2d7Gx1/Gk5bvDZ6RvaZnF+d5iMTjKYUa3VLR7Ck
bnW2Fce2YadRQ3rlkzdhLB+QESqUWQX4IpSCR+XTk4xuz9+JnqhTZkuJvAFD
7ych8UDes1VPxP8BdhnoG8siw5qf5MuMvNT21KKqnB3hPupQfzgGAYwsMu0p
mSZIG0XBHkDd59loLemiN54pm6DixNNbfHNmU0PyjhAEDqJzxVwL0JNB8Tti
7wTiFimKqlr8K5thT7LhOTMMdPytUnNf6V5EL/iym4TqIWqAECwJVYyuHKAJ
JuWF/SH+2C6dvisAUTlw/dAVkGUJ7a15y14axLgApJBtgkXSxqWcw0w5E3Y7
cJZh/fbGoXHs89eZ9YvmHjvxi6EBeEFv+jKkh8INlWpdkY3+6CLEdYAqs9Dy
y6K0dunhQ3DbUvrMffEpIvo22L/YMZfQil+pTG6NEtWULxrzfqb0JU+9L+iE
WrAz/bhDHHXzZHhS9qYzJd+1usNyh9DQr2P2mZHd378/blpvl8aJkwQrxMHU
3+D1CSqU20UBL5He7Jd2As8S6WEX441Itfe1lVm2sG6rBKux1kZ40uRdJl9o
KfkbSylVjW2PXS1dB5uW7SZrYLFO2eTKFsQNiBicOJbP+81c0AlNfLWGsAgm
c7bvao8PuOsI+NiFDSmdqkfZrXE93HnyCH7VyrHJWwylfH+6TvA99jqfvCrl
ui4Akm2AAHO0ECXEpFEqpZyzaDhvh5x3xrS0pykPiIw3ZXAbFStZ8rT0yj1y
41oEDDDKCcO4nuSGT2Z4YwiBqzssobgY464mZCEPr/UWuzeb9t51B1C/QhRx
HA5Vhsy3hk5NnX0mTIk/7vCflAkKa5BnYFu5FHGuZmkhu778O/1mllhcFVjm
FnQhsd1Eqs4kTtUQlE2aZ6BkfC/c7PjQMaI40gvM6+LQYxlFljRowCjJXVsz
a5Y8rLte/ttC0YYQipXrKdaxw5lCzPFE/+AQKEQpaahS/TbWTz3aHnIwLT76
p+95wOgZ7SYNwkzHalnuRQI2p8G2y29ZUqi+FeQUXDGr+dcRRjvF3bNSl1oh
GAfEExS/pg/pa4EFJ7/kPF/IPaSz+FZBNV1ZJuR/7NMDb4ZAozHHh2roAo+S
DrLEyZ/ANjNFSmvYDjT7oOOtwRS+YdUHO/A/W938t9SDepOlYMr/dMTn6UlE
jZJD5R8OQCAyVx/8J94MpV8InGYwlrOMW/KLS9Sa7gwtKpcV5cCisdJaN1Xm
zkmmr3u/6u+r2fd/Q6+r0Q/seFhY+r2FzHmh5emTUSYXl4X3VOf+ut5feBlX
SUHbEaEmWvEqKZbhjyKcJGJvQVonsybVEztRBqMkTkunLtgQp5jnDvt3crFX
C4OHQANIHLJz7J3+R9MI+Q5w7e6bJgnzlR+eEAUfBr545iNGmR/jMXuFH9ya
tuln5oHZ841nI4eYuycHtJwfP/G8O1vZ1s/AZDEHtdGv2OR0cC+J88osxjMN
/rTgOkLdOMmcZCBqCHY0ALP+XP4td6SU1OJU3rEvQdjiOA8wP2H5DDH5VqT0
FOFKH0uwEKQbk8BOPB38c8z2O4VTNmxKVAFifStNFBg/mgYRWsNBe2toQJlM
THU/Y5nR6bqj9YiupTdr3elbqOD/2Clmvc2vAqSuVt0p6DuamHrJ3BT/kqXA
gABUlayLYfwrXisOjf+xEXFKPUG51W7H0sfrt1njruGGOW6YToPmUjHdyA90
wONEu9ewC12s7oRfUGHtqVfNT94AnDBAX2/CltbgoEXCyHE4sNbFadHQGNc8
JNnFp27QtG2trLuM1IrqV/JxPYm+bEv7GLImWzhTBYeM0qjLdDgGN0Cqaxo2
KU1B+gwDV5ZQmof0+Ycik6Ek0MOTVJiwS29e+vLgSq2WmEcfWVdB+6bAg4zg
RfIkD55A3P2bYdLoIXi78n5ocqb+SwmhB2JP+lb4ydme0RNIrQCOnBnNJ2Nb
UQUjwR8v2XIEOpJX0tKwChQYK9ucV+iwdgnq8UT1BKIePNgqScKti/3FPKVV
BE3dWfhy8qDPOHT6E0G5sPNOs/QnmqnBRu1tHMeaGo/ZYc3QPeXkANlxAS8Q
BUzIwVQjNwJ1c9wQfx0tBOA4lkQLBtyPZAk00ec0bVdf56BS0pOJJwKFWr4H
7DBr3+wfkipM4yghTDP1QQmb+apcKmVh9FheMJgOKZ9g18Wqt3T3wWkxAJhd
Mr17Lns/XyO7QQ0xpWrUv2xgQIBUMJamlf+tQZRjXcmymVkd8wjmD1V0J7ii
hBPbVDTnf1Dvz9anDby7pCnK85FoJYQ0sVPd/lZLpohagwXApJZBZ9/aKKJN
6GGBkLmbnJcAY2ZQECSJCtGnM0weA38AaNA2v2IBqoI5kbuk2OpTuHxu7BXm
N8Ods2xjDuMjfWptK39PVWCXPdl9I4lwuGCyANxfFftFxwrKS6X8Us45kCoP
6FEIUpZ7dgdPnxXfEFOwtJ5AOS8MesLR/2zy+HTuZnXq77dzqnkNes3cCRtL
65Ncl6XI0ASCPjzri4pb6iK3/6xfTscthM55FIuMaJZV7fzxY5LHte4ne+TO
MENod81oBDV9bgUUu5cT3NhD59WYTTvfE1ztP4Yyl/G1IrIJN5dpMNG+Ffii
RniqUnGIhZiv5zN99yhNf8Q51wLqkBB5rwJCRYav6rzL1KmybYyo9THmyqT9
G+rZwp6HLhd9qLzlZ5ad+u4s0zWetPd2hZSKSo8bwGCYGqbp32rkppG6T8ie
t1BhkzFj3IfZ1QEIeqtwEqB4Lwj8B8xAvvEW240OXh5J2tAqUq1LmmpvT3fx
bNSLcyeyfn3Fcx28xVskFK5L63bo4vuTjYYjX8ziVhAiG5Zuzzpod56X7+pe
5YLDJSauyXVdJvgMZ0qFGU8SsQDVa7Vc3gcaNfocAecngy5oUY8nlXK3UEsg
ZzDzXV9fUU1ma9qQdXVJ6b4CUhnYY/LrOy8kFKg3GQfRdwjIPlxjjhIr/wZ2
TDm21YxhyVAwPhWjZgEvJL3CPG2b9aotBNhEO7oe36PF4mt2QWzXXZPfGw91
/YAzXztkKrhJPcayxEfgOpUtOgZhaDS03nEtJKx4CVsh8leewPpCmBEZsCnT
u4TyX1t1ixYngw54Br6r/yNBljqUlqGj2+oeSv+NYp+wpEUUTUMzNAvOPapg
gVyScbRcBNZafsKX2aqAlAj/gXKIhXHPxur60l9hwXjGIewKP2EN+ZKvLC1w
mbVYHLQRMTm/jvGfJEp+N3/vULPz5ox20T6in4xzjOQsIa+j1J06uQEnWHHJ
HgaaCBXEbhf2Tmv0THig0QQ7iuyVj+y1REGrTKX4Y5N5QdeSs+h2bZxBcgEa
Dc5XM2ZH0XdndDsMB40ahyikSz8/cjjYBbE3dUwxCt1riuBO/DBnIojuYDYx
xbkK6BjqF44T03Xm/yX6wsWlwYIYlnFO9J3Utbj8Ia49a287e44KKd4R+c8m
/7gRFcgAWECAndhac/MumnUWL/a2iFDcNfFqvgVU+ejm5KbnxPT9Nq4afhxy
dxQ9llPw4oAvp5Uegfp2jT9Uqc3pZnEvPD4SRDWHC2vJ/BxavvjAe/n2StPe
hGfAqwO7x1vr1iOa1Bh/6RaaarMZRd0Sofnd/Fa25fDYExy0mpP16KXdAU+K
YqLOfljkRF72SCGxE+ZPlo+4qBknf2V+vE3WqPZ/iFV1GXBNakjRcW1shUyr
w7jAC84YBQQMYmS6p0YfR1+uGYfUg1kEYOPoiqgWBdPojQDwra2jqmiRVXcr
IOz7k+U6WvCkLCWLMkS7voVxQZTxkibBKjLKoMj5ll2dQ0jtGkA+hK4X5Svq
UHKGO6WgafPhzNzEJu7TcO7B6RBazm4Q7VE4pwr1+mmibO7+M4BTYYl+1pCQ
SCATIrDY7AtXoGqfMxHe+/lSbVPJOD0nco67lrSwIojT8eGriCvVDV6Yvc+n
ZxDLTwSzUSIJRhQuQxrggsG1fov8bq6K7kqwlM5DP0460+ikdvBArQucnN1m
SW1U4tQZgEANTkoBL0kk6PSUSqPeuF3rNk2P2XBgCVlygYA3nfa+MgcPL2uC
q690t9X/vqDrr+YjYkXtCUgUnANY9BdtwyRYPGlQTAqe+zy8gUGNaS99rM+9
nOW8II5a2pqbeCO9YkORDRoKoS2eJEk9cXfY5/6qvAvq0kDj/U4hB+V423f+
RZnujObo1/4wLfG7/IeQR1Oi/hnUN01Q/YI2P24GU6HUqjtyKbi5ckUTZKsB
D2+y3jXrF2EexvuWNmIHtYUoZHUoQOdTmI6xVnnOwQpYAXJpwjE6mdJiWitO
bxh53Z2HSPA0jGMoC3QAFjJqOYFu7CBCr/qLf+kO1RCfJFuBEsUpvkl2ykyG
cF/R4t00qIkM3yTLtbcyVUM+hDtbFY42FzHRSqgOQHvfOv6timrDRF6203uS
5UaErqpJ1tMHdPMY4yGX38bqi+tc7/P3+OAqq87UmIrQfzttYnBujgh9GQMc
9Vo1STZ4fDBU6O3hcEXh/8/SJ5/kYhvK9ea3WIM2XGv8fNNYoKPDUtfg23p3
nx+YtulbJ60aAcLGTB5oISW1A1KYVxZ2ud39o8rqThAl33MBEXNP+pzkQqTf
boJBKH8FIkUhBnm2yI35baRPGgEq4APbBMdHHTJZoTuHnVqVh5jemjxDbQaF
nJHwrNZoKs5xax0z1Qnn+HNHfb4NRqjL18jaG/0pU1tb0L/stIFFMjTYCU4N
BK9jQMQkN44ZeZm03lAcvh9zFir1DJ8y8wUzA74S22XIuXR2PVkNPlmHdede
ljk4SX0AlMylOjUTUvg9ywqywHeSzWTEO4Lnsw7hgjxjqIKaPqp6j8Kxkuwk
m5qsOnHPolP1Mj1rdZ6l3qZz80LsxDajAnEzknKdsd1G527RsaAnIC5bf0Ut
4ffIqyAoEqSBgcbwIcEF97zWoSxWG5ZMfYkcE/0qJg+92hjDHX639upRwUpI
Gr6B3HY2Ib5M0cOZ2FDBLkN4yBkksvrHGLGgbOyLA4y8NPUMybuiQIk+5mmZ
DdxsYZqBMxUatHj6XGtk/084k7LkHCWfegRyFJB0sbEUEVNo2lXoLz6tJVWU
rTI6w1TVj11ws0Z6/Yq1HC70QLZGnz5UfbQu7W2hi05d59ehWtLyYxROzxsv
RVZ0BtK4OQSEqhaA23/DI+L3fXbZIanxDFZcVg5xS1JjxpIU4Dsha8BXFksp
gC7iCEh7lm9XOMurycVKkle/W85njbruPuu6W2ci7cX1cVX9TVb5XAQQf2rv
uR9gnvc4GmY0WvobeEWr2l5el6N+/xjvdhczswXqt8CGrjl7oXmjjIAZAvPa
U3By7KEHKgcTnLMGpwNDQa2Ea+uNakNxDqQ0Pg5Kp6g8fz1csC+zjrVECk85
F/TYh1txgUXzf2tDTnnH6ReL+kmgBmi7eZyRnd+o/S3n/rNd1bzKHaZEx6W9
SAUSPmrl7eyhZf7SJwYLBNrDCPbEIlsXUOWdz8bhr34Bp3lslTfpTmntE1WC
ZUvTgP/79fiMiahxE+VcxaplR2XK+Hm/2t3uPvgg6ID9hD/ko20/7c3/0/F9
I5akP1bpVvn1QQ+LPc3dVdaw29KKbLO4Glxe0sfbq3aGc8cnW8zqkJP4jHq0
zCZROPhfG/2rB5vSIYZVtpZxzbI/zR2HMWeLCdPZQGXwjbuJ+gr6ICpCqfaP
0j04+8QY8C5trE0zssm5m4I6dguFA66KLrK8HId5gjQNgGGw6qopaPtgFNhV
0Kb8kZuqWVcGolhZqUse0pS9Ja26ijbFtiuCwbcl0/5WoXKRoocwLlJAlKws
p06n/Zcbcp1zD+UPgQ05UVllES7h6mzKWvJ/O2om23xDwXkt60id59IKtLic
OPVqNHcxMsUrubI8YPUcVBmuFBppnBOEXFxaSpAq97sISJHOsVygx3j5ffPc
HWsLYNhA2eEJ6MgBtuyRYJtqI++D6r5bZsOGHcwKHm3NgTyCiEP6XkPR3yf9
mIWhk39QnAx2tb2LgyiDTBFoUBHwBpL/bHOPD7yBXGdJ9oj0bPICqA+zj8uF
A19u41OBrBRVmpRnLO51HY9GOdbd2Bks21mXmWmqYFmu7sEGQip3rINg93sT
KY8hXhcpjzaYXaagL4C5ZJM9IEroDKgQtS+OX0z6lZ3vli5JOAlNcqzaiguU
0rJwMFbpB4UvoWIsm+gtOBRDlhLCBNgzHH+sZ3l9gSoVdyVXlrLB5NPmdiG7
iJvegsxFOHtB6jKyYVSEFnHd2Z00ZjtSWr6NjAw44SINEJlW/9WQvE05yZwt
pLBgBOptaBCRWAtxh0wUHwJyLPH62qa3T2mCuo0fFBwexV2fCjHT19oRTaCS
aWpkRBBqoW7ImgYlLXXkCJqe/hFIfLQvPPA1lACCdFuSzuHi8pDMRVy/vrpn
51V7w+KhypnHILn5ZQmvhFUYMScPWntILl0cWFGT70nuxqt61hsV/GTpLCQD
V9mLH/BgmCfc3/7Mb3mJYS8FYzY84qpi9yIwb9ukbQQgZAEvDN3+9LxMKg0Z
2AdV0WFNahW1AkO3JFq2DTCcmQxl9v1k6Mfx0lZOr5QvEs212SstwHMZhraE
mNweSjRNNPfse8nfVnOYqvI30engImrgcEkXGn96jseFQVmsxnICmEM2Ey1l
0W9T/6HlYCY87QmvhW82cP9/wVZl8ZpOCtNQNtbpQeD9/S487pxEBDTO1+kU
pdJdMD2G49oV59WXFdThth5p2X6EnuQRBf8qDDbX8RnBx3IVsJitIGfuGkxZ
/3cTzkexoEYlCg1fTP+UqvYoK4Dd8/8NykEyfg4ugFuUgBl74E1PRrKN57hI
0BjV8SsKGzWAK2Yq+9uishhM1cpL8p8ShESIGFwhqf9xw9BbsTxhOv6WaKpq
46Tkjy7S26cW9qG8Zu2jXJ1Gm7FPP0MssUQHqJ4Whlos1/Quaokr7BneXG/Y
norpIoG4WqxRgekw1KaYIPOb0aqeLUyS1QgpmRsvz86VpQ5DToA1TwP42B6N
LcHGGCpBEfWQu3yk4FYtEBNKlLrIibDPTwRixFMqM8NbWJLGaKa5RkmWL5IV
9NfaPqRxkRwjdlm7dQi4+HTHl25ks704Z70xbYfVwblSXLYVMpGiAEpWo3uU
BddhwISi7bw+kJusYgqVWiWn76hQqYXaMYTv5l8Nl067RPYKIdXR320G7MMS
RPpY46oAbGgI6Xlcncg1Ih0Xt/+G6+7Tw+UcpKy19akXpJ6Al5k3rdrQE6bT
O3oBSJqublRa3LU0vW/lyWvfecfQdQ4fHybmw5NQnp90GjNZGwiCDOupyF1k
05+/d+Nxj3Tuz5ipm8AONhgENJ/mIFEJufDpsG6qvVPV5RSats75eSJzNroe
hzhMiSmNCHKB9JEs5yjm5wbikThD4VUsEvKbTHfvJl3Nr1oX+WCJhOD1we5N
vBAYCngo3bmOI6STOBmkkoMDUXXaR5r6UTQf40TYh5iVKDd6JcNJD+ZfwLvL
CcstjztdyqMzzrUTXXYR+44fC3BYg6PYzcDAuKYDtuOFyEoDLrMQHe6CEGz6
GNO2r9fuNgoXu8qeZ9d7L0qEz+RV2BTSLiv6i3ZL8FhmJyLyI76/Zu/+22c3
kG4HrrGupVqIh87af1KqqjxYh8V1j6DoqYRb0ao7grNBEWKG15FaP5I8ZEAl
L3LO67jhhO1OFCDx0uLSabBzJ5Rp+1/WBo3wtsmonC++luI0hk5D0TAs3LZv
x9Sgbh16+5z/d7UPxe33yTgulwjsCPyU9+/2HogST31vAZ+Et2nAFW5v3nel
xTqGvlw16/x6xuSLI1Sfe++yt7V8ByeGrvHO5c2sK4kYnBJAtmb/ZvYehjex
NH5rJ9qOaVGntJWiwceStGVQcxOkhR6HE/vSKpdzLooeSqOm/nGx2K5tj0iG
yNNcleeMpzXOQAjFWxOVLb/ehsnaVhX9OnJ8RDJM1H9qmartG49clZIPYicX
pbdBWut+zJ00er7u7sItHs+UOVJc9gLmdoml6XEi9+esSfx12QbKkr2MmTEM
e3NdSTIne8mOQ1oQuU2N4UHIG8uKfKHHkx8lmBlB8QD1cRXiFElY5ryPzmx6
zDnRnqgzdqoGtjYnCaJsG5SumWg+NqN5sTAvdLq/yjwJc9tYvPH8AJQ4F8NZ
T0PKF0lOjOryncq5k+GwCYiGWZqC9BxsnwfxYsDySOMaY96C/WZbYqTjTcQz
8/v61VR63yM2e78iV6u/eWQLpgXZ62aFvbCOrbtKqbA7WsxWxlcBloBxd42f
/kYQUW0CbSawA1ZfGfnHL6ELOXD9ji3v8ujjRGUuYV5cUqrJIOE/rC74Vp9u
Ss0vK1XJnTjJVYPnkNzEbvUtnJBCTjThhkPzjqyjg3gcZtSxo8yYck0Mb4Ab
2K4lZ/wPfwaRNSBHHHklL0OSM1wC6pAWZ8x1qr5LINrdE7Iy0OaHGPZv/PFA
46+HJUkAADqFrmku9wQnRC3PE0EiRhB77UYfOvR4Zjpw4HSSrD+RxEJkjRiG
FKbObfZWhoJEqL7VKGjezOdBjTnNIfTzTv8TWOGb/lRvNoeL9RAaeIyiPaML
ggTQadupsjQcA3tiLxAj5jSqn2Ko9IIcSnpIg9tU7/rX0MI88J//83BfUiwe
ax/hStkrBJgQqxb6fPHhH4T5XLPIR5EsX1IIdiA+5LshfM/hwixzeSpVzhKn
SarvZogVlNwR2BMo3K9RDzpo2Gxx/juhca4N8Em1E1TiVACN//My3saLugGE
VQtknaAVGpgy5dW0B7IGRCLuviPSU6XwTcl7LmxZtYLt/+A4ur4YmJMoViGJ
Oq4t80NuPWG3/81OALQFptGigwQ4emiK9RuAjg62+K0diboKdoAOGqn1UzP6
c9WuwQwDb1+NX0av8gRub/vZve5jnVamF86PLGorSelm/qdvM0vkmeHBevt2
DUyC7Iu6JuOezoMMkw4PhZrapLRAfUb5Uq4ESj+TOn7szzLBieZk4d2eJhrE
jNv17lhnTd+Gy6mkZbiZgpmBOf53jy2JeCSDBw1D1MnkevXO2ZTiUta41UlM
9QzW2Smtxo1k0dy7kNvMoAWoY1DXMszuby5T6FLCyfQT8oO2frNi9ZlEw8l+
ksLybLQSQSz8tS71e/KzA2Cl8iuvEA5cMkOoEsVwPoeHCqbb1QuvH60Lcoe3
2Gma1VLDTM5q9083fPqGKY9hK4pDXaRuNBPV1y+1VPZg3OdPvFsnEscqEPoV
HEA0ADNP6imFptg0ssGlFKVy1yPA20djdHzhP4MtK9fNbc2kngOiYwHhMNd0
3NwRUofmGjXySdQ1P9r4pm2QJG7Bu/IKvKfax9j0DkDJR59NkxeThptar4Dy
gjVAfPJrUO6eBGhfp/P8ZqxCDAUbJcHLby7ClGqlnOiC0lOm9wqxw7YVx79C
GHryz7uQzxz0Ug6PkZcRAtpNuExpX9LhXCAcM6MdZ5LuTKKfP0btKipQruZ2
8zWmmKVEPBVQEta0nKFVVgrl1zqCiZ18WRnjiTVRK5WHnFX67Mh1HJU0GAqd
ly+v0tYa9RKiOTP0DbG05+eGPQ/j/wLNpqER9ojIp0uru+GgPXJOTNN4yCBy
tcI0YMt/BbF7lahcoffP1wqdPW32f2hyWYs5gXSQcj5CU/8GTw7gLQhI0zf3
Di48T0w9nravKrpffbjrsb0WBTTuyhjQsCaJLPBeU6kLm9R7OwutBkFmfI7R
sWLVuuoOUzS/Lr8P1mGmg1LIgEYgSTC9l2HkDTdUrz/niTI9+jAeReg5+ddb
x0AKIFhIg4DsWI5t+ciDwT7VDszjbb6waA3+hhpLYDaksVhZnhuagbWXviqp
PqPcvP5qHEGqmSgRYgqMiXiwm0aaLQDCLXZZyYFEYQEq3j/EeZpngQWh9ylz
5VybE1bfxlIY2hwJUtYQqqwMrqR3VI5ZrYK5M+YN5HbZOsHq0euKM/1KqLpT
jKlvN1Jkml1TR+cJMuq+06gDQvPnedASYhPc3u0ru6bydphHJcWxoFDy15pc
H8tsVawhfhtZY64fMUtUDqfXmGG3Tlwrrvu7qKnbkslQ2o7KW9787CkHWYoN
saq3eV4Syj/dA845438lAY9/k4iNb50MAVbbh0ryofP2uefmEB/jGZHng56P
c9H5QlwxtpVYpZxKi+e/9+TnXq+LMaGkgbS59s/wyjimcrk+dXFyrVFuEgAA
DOJabebIHuSORnbSzZuWxO8mTaBWYDUuhc+X9nCEf3oT7yPDb0NWv+8e/Yza
9Lg0YNKN2TXJDQ+R6gQSJrP+geo2wsx+JMqmQCCowf0LLdTWS7VC7OVYglM7
0Nv9cBjFPs58nGdDGuegFQienGnYtRuS0eH5wBP8SYJTOSCsPP/0OhT3i6ta
7ZiK8kikMqmokjBEJsL+u4dDLPip5aqPjI8AKg/WIf+h/YbzhSdNR8x/4Nqp
i6HWTLExY8WT2JUwF9sU+GRlbAg1rXyAgW78I1x4QI8+ALdZhnq9DZpZ/hMA
LQYFpGCN+Y/E0NRw3i/DfAs2gAdwfgZHJkeULcK5ab2MNfKRc6+CCoEAsla/
uHDA5L2rJP7xx8YsIbSuh4Q5MGfUmh+irbyLU5DIKO6c/DkcIeULs6QgyfWA
/m4k5Ify8lkClh444bkPiRfpFigotkOgPyqwdVAUkx2Oo8BMbIoLoPxnvxDY
/ruXaO4y5o0hdoDyJV+N03YfEosUw1yOuI0slc1hV90EwuLIeHHiSatv8eL7
ajCa+68rEZIjHG3LcyFwRLd3btGH+0LALBJjkVCiSNY5DpnZWg/iXnOPY/zj
6T1jx/DNQV5zb0+dNI4xzQ5G8m2bTAD17x/ivP0sm749QrB0m664Esqje5EY
JMBsABiYelj1KsJPndZ9sLqvu2IclAUAgObChUR6P36Lz0LAIoE3kOC2cHWP
duKYMe53LjFfQBo3urXwnGeF7ThCnvl84Pv0V8p02yr3SrZTXkp18RK+Sthm
QdiEuC3h0hc4pd44Q8er0SgememZ6AgOIsbwkRvjguh37ihHZljBzJnJWD+f
EKZoyCmWZwJWhYJ4Bm+82Cdw3p+bCPJG6WEFTv6rI/u0zfWZT3l+tBqK4y+r
FM1OqVkaFR2OZZrjjbNOixA3BdRZ5FJyJOWvCR+iTbBbcXH8OTGffWD+JUic
R9VCqU1V9ahC8QCLVJ0as/JXrWqJmSYCT+GkDPFWHRpA5t5gfmgoJHK8FdyJ
dijOzAb0pK32GJNDwz0Tc2MMYYzQV9hTMHJPlH5QCiYZrVFgcADBT1tf8gvM
r9WL3i/1CZcR1SBkx1QPGBJAQjjXwvAm3ULa9dXHL8oWZVOe8Uun5kDoqlw+
2gcbuo4QrkrSDzMiODDF6adxDIWeoO+iZ86FI8c/V47wQr1oR/y2HNp82HaU
heEhGXOJpcBBC/d6bo3Rq93y4uhtPYOMuuDS0ePZPCsba+yvJwEZI/0Xj+sM
gt/EHWR8Va10j66xs7JUCu5StDy+wxjRSCc5+JzjWRctSk+g1ILVvzhLbEJa
FVeJigUE1w1R3VhnZfh29cvVMZecENQ751mBsmh8dr5WEXuLbdZ5y+LSut0e
/6+iloAyzP6uPNmuwa7wUWPFIDHa9QVx6iU9yA90XQ7sU/8FTOp3DosFjndA
PLxjK3zz9rq3zw1MXTImNxIspdMMS8A+8BDujZTcYT/lJMaxjFCUwMABlxbw
SgmOGHlccS6DN/NwNfyEXZ/SI2uJoxamXBxLKzneOLaMvYRsdlw3RLSc1dHW
OgryeE7cmGPvUf3/xicWNi9ZmCvkmxERPqJgp2vGkl8bqCew5n6Q6ost34VZ
/vDjNYyyyh4vjED45+EJGF31/aIfXQkg3cJj+3tkFIctlZJX6bNLtKQVTRdm
WQE8+67UA7OwGQHtrqcuOAHnZNS3avlsWoUA0cIQvIwWSQzvPEwRBYbKs0Mt
mo6JkC1r8+TDKUWhUg3umzMv2YfqPAioICVHUptsle72AsJlGQW3Ju2AmxIo
vp0OwqMEjoh+p7m5652hPpYWUF+HtvqMjOAezY2zKHUkmfAhSo5Vv2zcwDqQ
5ChDTbFG3JrdPm5pBvsZCYtbEEwp14jzcJlYtTpPXXPS9S2K5ufx8qez7k/n
vv0gu565xbfzqStx2o1WtobA4FCpW4Q/EWIfa46DoDSwE0uI2DwcB5V+wfPl
Zzj9iub6ZVW4m/6K5weOtZtX4WwlQvGznPtiVWl+XQzNGjMBMLwrep7JHNsP
M1+5VQfOVxUmrGp936YIm3rXnE+8T7u0o8zEjh/K6DjYJdoG7rx+XiGU4uE2
cWOn5tvqwhuJA99zdyqomzQFiDFroPUK5TQi31c+i7cGzNfwZeaHN5sFW9c5
E8Q8zrigKx4ntYXr0jcrIIOu2hiTkLKgPxuMt/NXRtoGyRRYOWLAtxFzEZEz
06WecBM0T9ZLhhUPnOQSXGW0T++SWqbW2gsDwag5+d+UhD9ABilnhr6xNT3K
x/AnM8/mk2ZagedLn3GBN19J9q1L2x2FlCGkPon8PvDqK673QbRTo3/hr0h6
raO85bwccwL5w+aBMzLMIGpDz4O2IJb293pt1YSO88GjaOxKBs/tmLSuWMjf
vGdDkUaa8Fb7sInmJF4UB+IMeZbEGQkjc0VagCE2aVYZoBInyH1BVWgkVKpO
NfeRwoAGsb2Mett97FdTtixcP3WdyrkwwAWiMYUO4/Py+mSahYKUVyf1wGmH
jXRJadIv9sp6y1niIF8gHtLpsRY23Sk/Mdp6odiol6YruPk4fU2j29LDX4/Q
N1A73w9gOaemjEK+mFg2W8cx7h3bMatvMKByc2fkmto7+NGOIS8OTTUw3Twi
pCUNdIInHhewXYnNU4xS6FlcR3d25uksYLrUgNCdm3+x9igFi31R06dvEN78
OIGafNPp9G7qby7STdTXfMhVkiuZa1xp85rZzp2SzSlk+WYm95ELe48FhjXs
AM4IG5xhmlJaJzVcWdH4BKpNqkzOk4DcvZ9PraohNd2Gj5jU1V+xCOqtFGjR
M5dvZ0VFeIeM9rsad47FFzfV+v/lKnQdy7O0xIeFfket8RokJPyPwsqUaOY9
aKH57zq9d8TxyIfau2k57vJx+PhxJCSFYXbo34ACO8KkbV3usZEEpaZAbXf4
yWmgsDmJP0wkkWdEacClZd8CE2L3AHR6wfhvLkJDheuy9MfBTBLyuk6SZJeg
83Fz9OX23hU+qeiwFzqPw0S26tr+B3mKvfYMY3yDjgOgFscq3f/jT68UNQj+
U0QoFny6t21hxu4tO+2l5uZLiv7GCuVrHzU45WWqjusFedAlWnX3nKu5oX1v
jQpXiif2hTAQLBtG2KNsWIqKg1IbE08TBwE7YpoxUrji+fQCeCRUMladdgWq
tLqBnjnnr0Fi6L8skh6WYaviwoJR6puw9Oq4qxEBz7EmCokSX3ObCigNJFjD
ssydTUiV5bRbqPirVLusXMu0N6BVdHTD/xXyhFrCofD/JhPsyxNvnXepn+R8
FmRTQo3h1upAJcV1e8xGT2a41iRAPhAozSFPP/y2Zhmg9d24VjuY1zJxjOcq
N2iW8sL8MvWzUKLfyT/Pp4htqta/tXu3WXhmwg8qhMxYWXZ0U44bv7iMJW0u
Mg3l7KWBjxsxTdBD6vo+3ORZCZK82Cbd/gB1q27ogPi+VXcCE4Dxf/0oI5KI
H3O36ZQgjDsOxfFmMSBpgslwvjmz59+21ukr/mzGLRNUgaAtFuy7bC/5cNTH
qGMLlvK/lTbFlHd+NX6pLyxb3AbnkpKBlnqdaNsuY+PSKjyz3tgxqIwhuRwr
JG2Rdw/jzGf5om7440lQYcyKbRrux8YygInwJVDrLyIn8eG8OUh+iMqXi1ew
PlfrS4qTIMQJqBC2cj99jdyG8GxGvjX/r+m6YAojkFE3YftcsJrt+hQPp5q3
CXxor7aOXfWwEBzA5X65SPEeMHb18mOHPZHodc5txuVIN5HrDqXTBb59fpG7
j1gFIYLuwDAxokuszVPeX4c0CQGrZo7Kohbc40qcFcn0/etjxPfO7/MU8lNi
BAnUeZb6QqfYcy4iaq2Nfjp+1tvPGSgV4vpEj18Mdil9bnzNNCor/fPjEGBg
b3ptc41moo6AU1Lrx8a8e1F+Pu2P3oeikDXMRJbDPz5l2JoChbTfs8jVqTNo
l7+p8Z7oH56R6FFkEd1vYmNxpJvRDUILT4Zp1tvAfOf39UthxvlVOjsre2ID
9fGSozwYikYIb/ul5gd1C9b9nsSjnLkhnpMDyZ9tFmnsxDdVmSzNgi6coVaz
ww4waFbxtZgVXHMxmDXOS8LLMC9nAFwSeDGadSnCBJGSfCIrJU4XHmNY93mH
BPnJ/uLmnZXwfSjyeG3W3AS5lFDkuXy3O7EMqZopDz8xJWT8IV7Z1y+WP/9M
zTZL1G64Vp97R1Sfn2U8LzPT74hYKBFxLSBPCDpZc+pZ+ktZ4AYAS1yj2R7I
oqWQ2lx+fEA+IU82vYy0K1eDxmfNhLxMOVgTjnsfMRo//DZnITzUtY/ZnR5a
bsCw5X9LJ2tLcgmK2IdKhfMKLTAHwEl9kgWBZ6A4dhgpORPguTlYSVOhSF6S
BltzxbfOjogkCi2BmnTdsLwUvemb2B7fu8Jxq6DjwmLHqTKvK/kbNzst8emL
0E69S+cfrNzlxLyE3aDS/8alXAc326cDeBQ9S10RNbxQW0VnnEsvV4N71YtI
qUZGjV39acjeXp4r7H0H7hbOU9KvX6l2XhNDBGDDmjOANbq13fu2jzTG8bVK
q6N6aqmdD3pKWLr+a/ymbCB2Y/2p+QYMsq5vGc58RGk7SopuS0ObwLm+GLtL
aZmoRrii9udt8jl61zwjODLi5BmIT5QMKdm3GUpFkNcOpdPnk7UqiohHN01I
Pq2h0dQp/bi3ASZyB0m2vIuVg/QrhpLbUvW6NKRj/EVfD9CZTKzw36gRttVE
moZzsKLvjtjxiHhrA9mJkyhEDhyuvH1JwjPtLvfst0XQi4GWZZWz3J5OfTnD
rty6q2Nux/YEnlPqvw9ErHIN9Aq1a5+NejB/0RKmy6/Mp68p6NSoeLwI5JON
9nZk7QjFcIqrXP9i1y0jggo+2ZU8wD2rAaLeWCLOfRA2GjV5wMTDPe5xkPhV
S+bETDlH91AaymddKqZ83Uj34tOXjLSf99/3pytCblmKyJk/UN98POPk8V4B
vIHiF4a4ZYg/ZVtWRwYfZU2OMyoZuPlPHzYxtecHKiJg1Xk6DG4mofHuNS0C
c5nd5Tn8HJwQfam81mFcRkaQiuOGvBJVlcojca1JkREnP5SawjQ3r7Q/WHwt
jGPeqj0yLAIm8KdOFVsdsLVHiWkAmgDvWh/6V/r27gI28OxwrXuPeJM8wURx
MCp+BPcZ19i4XtMyO9NmnDKVmialHBRTQMao53YoPBn3QuAd9yLZQSq0OwDF
vbzZb3qAuMITeztuWpJaNYBFCKQ595h7RDahaDn1zBU7aZo+koeCYftW+woZ
F3EfoPhdEx8WpnsViDB8nev7pDty91Q7YIUKfHqDfOEI7lu+KVgw/gcEIdHG
sILVNbmDqOTciWkLs0brp5gI4QD/KbadKGOvtqeAjvrL546gPE/4L5Mr5LU4
i880dbWT/mKYCiR/8QQti+wgDBVlzZdZqJJm9hqbcBHCeB8IRGvD75Gn5/Zh
rJmj7TqN4ec6XnmP+HLU2QKClpIXhufLFm/+NV2CZX68zbQGz5Z/f15ABPE7
Uus+Xnir89tQVJBcnUNVWQFf9zF/zp2K9BwjNzaTdz9QcAzAThW0Nn38Dc6p
7+YrTl/hCEfJTJ4ZwtlF3k/yAjvDgofGOE9kl3QMclkv675UlGvq4hPZk6al
Dqwb7YKociJClvdqzcbZbBtWAgMhXp1HQVtT/+ARXxZgNIYFLNFEqSqAxcxL
PsLGFmNQrnmF4WnesualB5HKmDCS8J9HUdbz6Hebz5yn7fFWHDj19XiIzB0Q
K7hzNwSROc0byACMmldsrCNMjv5pgChRQ0ziOGCjgqiy0LynZHU3nj8UOkSm
FlVoxIf15UeATLORqB0qMkYYOxmfsAb1szDGYvu+EhprJVAkkh1lMgrs/sGB
k/HTcps/rfmopuhgdNdzMqgdUlco70kLTV+vtK4S6zpN+hBoTiX2g6QiR+0V
kAuXbQr1cYj7MZZXMZaPkQHQxi1MzNy+6buv8EmBtLZLv7z25EjdKKRBEDxM
bnkdIhn3u6DcrzqeYAiLLj4XE+jQav3zOUv97nnYUHztv/LMK6De6fWbRKqz
7Heg40UZFJ9V2ug74aNRHHmiwM0SFU/9DTIfDjdEl5Tj+v6uPpH8kPH4/PZY
xlOlhByY+QIDWLuhmsczXRQWEd9S33X+uHZh0obvDgLaLkppv+MyX8g+NNyJ
baQeZtJ+qbG11OkvalMtPsL2358eCrwZYeiGGiQZOizL701Dg/eV1/ZE+pUh
TMfRQdfPnKfoaH3m4ZzDWeMR0Lzwb9J/v83VOXWdYOKOpnXj9QX2P9xHNuz+
PssYUZ7D1FO2LVvsMNxpg0NAkxBx+bB46jLofnrpDdiwFQls0HnR9xFXvBkr
uuE4on3pDGXUzABMrpaZwajiGTs2R+toC06lqgEpt9mr3avGJP7fvkAekT8W
EPt7OJyljsQZW7LfTpytvqgoC39F3mb/A3BNfYJKfiKwu4fBM2rDaD9mV1rC
MYUBTiewl6DC/8gXNW0gQWwgVCXlyKiahlRc/ovnEt5xd3WjXowWY/qO/22v
hvCM2TWwv1HhM37teZRsSi9AVYd9GtYwV2PITO6DSF2EEOE7vEdEqkojq6i7
QKPRyOc/5zFqpnCvFx1pp9MSW4kds/VQqXBDdyJ2tAIEf2T06FYlYbio42+S
IhAnPczGtMaR+guE7vZy2kY8lFQ+Gq1xLZordR8Ajm+lI8ShGtik5/ZHHvFw
ObD/Dp24P5qzroJUuHMpEyn0il8r1tjVjDAw6v8IInMlruZuJn8La9sIBojl
R+LP3Z/DCPEygHig6kA+oHMTieVP4OYGO854XyOgJwRPGrE0W0ARcWlFarsU
OJVOCRGAuSyTB2q9A4GKClW2jbkHOjvJ6Dp8f5FkIFucrsz1brwA/e/kWxty
PVhkpGUYoMMcdThVB/Ct5V3uNATMs15WRxS08v61AArGdBtidVlR564zVF16
Zf5J01SyMIDEzrhZ/q6dNzVTxtj/A/Ggl6jCcr1fCZFQcIxGs9RacuqniqzY
k+lyNt8OsabmFvJOctqepKes0xa5Fs1BK4AdpABF+59KszhdxT9IthmCvRgH
MUBHuP3wfIOlPD8UhVzR0hc6NADvamWraCJTyfHqzygloadySPH38421s0/E
ptGNXAr13aS2mMCIAN6bEtpljEPQ7lr/jeE65DFR46twMLap60TOx2gEmqWX
ZWOhBX/YpE/r3pIkZHui+xM2014zpsw1lDE+E8uYS+ETdnNCNYPAWO1ZMS1F
oxVy9njuRL/nJTfKcGFMCvhejr0lsYWaCophVlEMqXdaWoXN+yf1BdEfDtS+
NYRWjGxohS4v0K07lNnB+d8h1aLRmIevs29BlLLWGYB8Vu48VPszeE5Y1wX1
q22TKkKwF3USiZF8JV4LmSKdE//Oz5piBrWGlpR8+bjtvkS9sUxyJYSxNfw6
JJM6feiSqQOvRyRBWfPhLYFtdag7UOut/P012CsK3oS98p56K9O2H+dg+LvQ
fuBXyl0c6lrdgqX2uB/sZPKni8YB2gh3vaT0uD63r+9gjpnHixfyXuLCMi4h
XfKPLFirJMXwjsMQLgYPv589kpKohXTk1dlikcbRUcAgst+LOWL2Gkt6byKW
WyETsbDouNjMd/kN587OjtEWpKqjXRDVfxXYk1hnW7sY0pOTAEVK6fQKcAJW
sb15Eb82Ow/BA4ioDuS39rwxwPc8XFEZS9YcMPhDO9Zte5DRLHqJMpNlKdDq
BXttiPMjWxqt3kTJ9qjY/AQnEYDUXGwsLmpfUDJDdNITHLPRlIUuuJJhp7RE
3oucODLKttXJXhSUsnGugvMxQxbMRiZwDrlnm9hWJPeIgeRKOrg1Z+rfC7dh
maXZ0JmyuNIVoho3mOmcAO/x8JC8NH1FRTgJOa4enOqv8HkGjTrKZ/cy3Ozb
9S2mssPGtkAvYU5J2iPpKuBzVoPgi/Mv7EqY5dt9IByjzBLglTOyZoQipqmh
Qpuir8XHlGRgfv75UE5CY2AHfsvo9YR23+4UlEPol66wezImCvxRRS/N62+S
rFSOQ2Xzetu1FbaSmxHKyBDKMA07uE8NUCQi0hmFAGx1bFG5PAxccFLYkKV4
nJ/lMmaLbGRwMqgzJ38kTPFzGw/LwxsHYQT5qFoBi/wO+tzBosf/NMq4ZACM
cDhPgq3T+tYTtMcL9lzmRQa2kXmspEzBM4srm32bcS7eu2M8FdjR9RZj6TWe
w0G7nI8eF94iDW+afJ0fJxxbITcPz/h1EvQIU6ylIYu9yy+tU2ELgAJYREGF
S4NrVmqEpmQCeg3RZlOr6jfWdGEC7d3EL2B0WEDY9U1nS8AbPipwrm4yVy5U
Tcxl+CVF/v/8IsmLDz25avBNr4Ja4vFpnCxCULcE+9Lr+zfk82w5p9cCWLDY
H1fh3hrXYRgMTXadIsibonZ1npuhJLnUektVV1t1kjnPN02mVm570kXjBktb
/L19FaYzhcvqmb9ZjX09Mxw1AwDvQH2Nfw0b8Qd4gP2E/B4w2jYUfOuaPTgS
qTPWm7Obq7+4LDtOcm8zd7r8zfAQ4zBOKtPGBzaGTzHEoUCMd31crwZ2HhGD
PGdfRqxb9J3pinmHqlLcQWJlcyELD6cfUbKgOVONtf89I9+xDSZ4/0J0xhS1
xVywaVfvl1fSQlIP/wuS9Qi3kbDktjHkiVkU0NsGgRDMxwLqKRwf9Tu2xQBD
qyeUztw80Ayula3DJyRrGGPR0V52vBshxNfQ00LdtJLq8e0/Ftq17vfLT63j
xp3QpQoM2Be9EaN8+T8vwaVkhsigPamSCaIs/EF2MUOqEWZECpj/Qw2SKn4F
4L500Re4qQ0IkLkYyA8vTmJHHBuxZVIzIoap7Dy8nGCC31ojIBaTg7Fz6HXP
ceqKqigPLqwzLFC1EY17Wr86am9nkfea2xWxQ00BVOIPJLm25+muHN0Krn8A
MHGug38C3BcVtJ82E9rScdcOBrjw1n0cQMboOySZjYRLcsX1cZkbUJV8iV59
2XxXuX2z5mMm0bXwOOqKFAP5/eNOFYo1a3S/rXChbLEP6flyE0mQqphS9F7+
b1JHmBLL+CaT7E6ShQ7TqA9uL3JZnhxG7gIxkvG+LylvKOMGomcmDhNk0SBv
x+56QriwbRohfcZInwO2X0MGrbAFTnmvDcOnmEDW5fziFTvwAKUO+J1zQzfi
FhKXlLA/8yrLrfh9Vm6K9ytZ5yWr0dnvVw90hurqPMCa2LgmgvlayH/6KDBN
hKoHyh43ho8yIv9vv22BoFjTRVGJodR0y2iNahgRcfPh4C7MAxmXFP7Gbub/
jFLLM0/2FA7HKiedehm/t65tWyLT9F2Ybl0NSjlpz56rJ5flxGs3DdgwtjSm
m7TmNh2jp18irsYomUmNNeIo8PB5UfejK/qcyC8z4Vv5Y+9OcJgWxbeP+72e
/tvzesaA2lrIOQjycv1rcg9r6Q86btgs+0yegKmsTT1mmy80lTYJXAEaIoTW
FODuIf+YaIi7/9cmXGeKa9w60LApos9r5WAfp5qhHzbk1hkWgAC/IXd1b53y
yAxsVcsTSlPpegeBpc/uPqC/MWafVNeyAmqvRMoH83aG5VG7ddJVZhT6MyuG
vBBDXmhq/XgShMQ05XZGn3EhDyxUHP85bqq/HGl7mKpUB8rrxdHMcV0vLjOO
Mn2izu93+nGXJWss4VPRzztwI39Kfl9+JMj2Q5lKVKQb7B/mosSuJcSNqpwm
Vi26wHnP2Kdl/xmyilMI6VFsPT6PALtuoi+6LjsYOm08WQ26TGOdWSuLoCW/
s3yN890p4aEfjOK+I+AMQm3rHROKNOH9ubXG1rOgpqHDohQ3cBhfZecnIFin
qcWHevlYy+pstNZmhZvHWCCRsMuWfbS6a56uBCpssOsHqKnH3yeHpliIUu1a
BR+gf8QTeFSwVgf68l5PJ6iGOBsc//g15PVW4PGMR7rYSLDvDmz16Whmd+Yk
5084WCjjUpNYiF3NjC88fAXY34X/QACMrB7I0OBa3zgDNFC6fVX68G7Moy5e
/9Zxq3UWWWvBEU250OGrX63pXNS5W3h9lG1/FHlpEqzxdO9Jt9AgNDyqB1Ct
6k5SCMNZOg85snIdpROYR3JVehiEq7qSd2tSvjOOggh03wBiNFYbF1H1+aCk
fVJCcsonh2LlL8ED7ri/G5MMMcIIiXMI981cKzG0gLdgjfGeoF1bcIhY7Orw
wwsSs/n1LW8agfso5JqsniaYVRZJO8Fe5N9EX6iCrGUyVqiGUGZL+gf2Tt/A
UfRIETUoqJ2FZ1s/eVH8N7NnxQYJWMWA2ga+IvNUfvvraVKAWRaQA5rrN7ej
wm/roGzYiolh7wI7xc7tj0kIoQXZP2bKXs85HI6O6jCDr5rSxMjeaYCBaqsM
Ih54Oxk9lwnmOoJnI8N+5HFX9b0BJjLmkdfEbuSqX+srkKhIzD0hYCIE7/B0
3zZ7rHZSlrrV9DfO8NIzlrj/LPxNlV50chpCeykI4J70zTkmdWXnxO/b9s7E
aBHg/2yscjubsa/AbQQtVtQgxVwsnUvkKIn2m5eEI06Lb6MlkDbSmTKCZw/z
BwOMPXoVbbegNKdk5Hs+rN5po/MKyXKAFzN0v4q5QJSaTaUm+lSKxUlr5x0o
pqOVTyFl/Ja8xxGU4E3QHSSmKerHWmN5Dzhcgl0Wrsr/luT+TJJHC6FTfwIE
nAlj47PAyVawZa4NIV/4ltFIYKfiHtVTNnnM8ZKX2Nr9aOXN2QFIAqpi7uLK
Ej8YVVHR05oJrca3yvbBnnXc6D2/XXnTTRuUdWyK5G6zV5zdGTPjA15Hp3ye
2le0MJe/c2X4Qvxc1nAB15lb9d1NrsVChrrCwfne1NL+nM37Lty4AGlviQWW
klr3q3BrtVnKMovR8ElgZ4Xl+xbLz9G3/3sH3VpWQtGzCli1IUHUKO9qbvRU
aSLZB5IRtDyB+5nw0k5jHWG4IEi7topbwGmHp2GprM/MZZZlR95fsLaEBDmK
YckporbyUjwegQjd75URfmNrQjYZHCRCbETRUvC9DLTmCv4utjoosuHUHkpT
eJ0LTkdfsm7aDFaYb6ORtajreVZprEzyTFRAGI6TxVpBgBddlsHV1Ez5cDkC
cGJRP1glFrMnMkewOfNUkrw6smWH8tXgmnjM+pu+l/py7pJ8rUD0QmthAsbA
Do7fQTNqVqCwmbVjhdJnyonha1I3C4nmwrzp6jnoHEpKo1rnNvuyWAK5xrSx
EeyfL5wM6fl+aFACtYqEaU3jzbIqmRYkl3MaYqvgWtsfhFc3HC/+cq9KRid8
U5ceQeyiGmYKupTMarfLalgxZDT67eeftnf80+kInrlUSh2hJi9LzYyvzUK3
4NuUEgfwCK4J7rSNZQP8kp1vJ+CGq8lbIZ/VNtBrSFDdotRK9G098nS4BnVr
StMRfMkf7M3Bt+2wC9cU6qC7ZUey/0AuA7BDGmoolktiaujadKE1+spzrrNW
nXU4MRyISU5XgJNSWhH0nMv+j4EJx7CmfJfRlSHMh4Awq6ur6fh1xvsxaVzG
+ZohksluOigkd+4slkclxflOuSorGEjOGU5qPPFL7EgXdyrNTsFLJnarObNu
+HEascFi6U1ngLe1/EQ+puEx/JZx1kUFYkc6HSaw4u10bwjpGmGMzlAlVq6m
vwG7B4CXR1UqD5wMfjh8+xzrBhTPF3ihG9tToychEHmSiruu6CZ0ecBKjcQb
6cvT4LA2Bpmmmp1JCNSVIedvouGAEOIx4nv/eLggGclB1xoIoYZaiEmOQhCn
XSmZvDoRaf1ii07Zo0TzXcJxFqTk7IgG/8inF+Fmcwqb9rhCNrp92kQZLeC+
hOD4PNmnK5SrngCf3maBgbzeo8pmcFGVoAwQFzcNVawpZSFBvUFKlXiWQrhu
9VC8NA4CFOGg9XAt8qjk5SzhbDmOQH+pBwCPGOk3HJySBJ+UWy2mT/+TYwYY
I80wsOTJjYQxFOd7vCVrBt/84jpE6x5PZNhu62fM6ucRS5FCKiEFA3wRjmCE
v6/VmkEYTE+I5E/skwNTDL6LIkstToEwQChBV0U/3VsV/FM9Fz+p9c/Bvzkt
r9q1IBkZhxtrXrEvOtn9Obj/eeGXusUc2sI4ot7pRsgg7idGLC0bWJ1ca8Zl
Y0+QjQcijkRUQ2VLBv4kCif5f81ZR0RPDTrYvLWyltPeiXm2ZH0EM9aFaf4E
nx7KMUIM5AJHfGsOmcEk6k1eo0JNpmqFuHOdj6WlNLl4adWU8PABWqdBtNFm
wBRt2veD4Lbs0w3jO2bYWux/AUGF6hKE1DJTyKEj/XDT3WBTgZk9hdlbh8W0
1B8arzX3KwV9mlct6FkPhVs9vIcO4nACACCZ7qudirwquTCVZ5vCKCmYseaS
hQiLNwqIKMou3TgfXENly82WeFVOyQAW10Us+4T+2Rn6olzaN3Vh58tl9DeU
Gx7NSQWnQR7P+34ZL0jjJJxkVMLvLH8HofGzTDNRB8FiNK3Otat7ScGZaWnw
jQBASOHCpXJT1WdHaLpGMrjjAlz1g/YJd8tmn55E4DL6mhdThiZGHFayMuxL
kPqNipQT1s+ohTz/WhFCA8uLBLPUfMAmS3+c2eGArgSR3jNUPlzUIEZ8msjn
k+MTzU5ZWItWUR8L1D4tfib0/V+U3l/scb18QTnveWPczRlhVYSRHFqtVew9
173VSdfjq2c0gSSDbXZ69+qmIJOfcYX5etwN5QyVc9zSR3o4CbSMuKps+JRR
l56hwg1NoLuhft0if7FWMMcSgQf6zZdpj3gNRYldMgAShcYnU61lPz066cPu
E/B+BQ251T7NLn7jRHHxd4vLNrCfZD6WRq1Rf+ohZ294e3K3xHqgrlNplXmo
8elS/sISsVZSOFZEaIuUUMDvCV9qDu93TwxdCjo07oL2Z7b9053UYrrAPHGQ
YkD6gslOoqPvufwmrXZck3vPUUeSbgf6L7Z1LMzLnuLZgrTwrZ48nEHvd3B9
z+KMZ3WPp7t/Is+Z1Py6IBmlgw+hRigqYNreqEWVw7PaE+TcVj75MR9LImVv
HIMKCb89/KiHRFjD/y+41yBV5dGoUXgI74Cdac1ZWObbuHKm7d81xwGSxzzd
xHny4wDy1i8IWjh12zgbEfIDmXC1A/vp8MZbbNCCRl3orktkjuXnhQivCNmj
OWr4yE4G53wRlMflNAHWLHNOiHRBeYtTlNGWmuOJa3oD7xEkx8+gap4ABms2
WUaAe1+Y+b+gtVH8Lsn8fST971z/AOwAWwX0MKPSEqD4dvq21+WTf1ecXGeX
b/PhHMsVmag258QAjxiPHdWjWCtM4i0QZNfzK+SUlmVlOm+8b1MjcyrfWdHk
Z8XDa8A/O8n2E9NwpH1IE0AaihnYDxG8l6rCm7QMC67HCayQddfSfftg3+w3
klTciYeqbT42Cv5sRt78DULuZuK2gMsnIkX4n+WLiHe5+3aH4lMBPf1AyQmD
7jvLYDjbZQcYClONkQsbzsfbvDsaAvGbTju+HkcAz49e9caUqrs0Ru8PcosV
o1827vh7cK7bFs4gbWeKTIY47aalOgj9sHyeysqAffoyvWkgO5b0t1fHfKsN
a6RxQC/A2BLcwnb3CQ7B47rOKGkrrUaWq/kXf6RKpGWxXRPIw1s0TV6JXtPK
vIvnV2kDdTaRI9hY1Ckr5YIIp1atz8cdctEaWtiGckTQYlSDy+Epe4NATvk0
FAtfKWNDZPuRWxVaVJmXmXU5ie9vwcgkdZ4JRxDMwJeQ0QIOLfub3GaqD4t2
NIU03yeufI0azBS1Z1788dkMKFkTiHYMsda0+zKfgtC1OAof0dmZOHlwbIOu
jx9zwrrH6CesZQTEjVkAS7fgvnEPx+XmDYCoAP9d7NVwkPfXDi5y3M+QkaGN
LudsnYKb+Wkdb+KQ0o8CF2IK4Br6JMWgZO4KKZb8RzlSY+azRBovIPKb/12q
V6yzo6OkKtIAvDthqE6ZzgY4RWXBxAA4XwxIzj4U4NzPVU3RhxEpZS4IDbBW
ygkhJEh5oNd56JnBURVU3vpNVnfUnnGF713w/TzBHV+kdTUniNjoR2KNzKs2
eIYxTIyktIU5RfJ+8aFrSVSLO/aTGBunap9lw2wSRS6CjeBtLquu4CS7PdkZ
wppwD16e/Ixf7nAJe8jh7IEI7vpZQjpuRAqqyx8b3kBo3x8OroCgWyaU5Jyv
7fah16furj0FRLI0i9n52ivmM7aJA7yuTk+ABvhb4bnq4q35sbgNW5dPqjrw
KOYGVoKiKlha4ftfnSQEBYBxugDJnfSYzt1gQ6ANzaQz4aELn035OyyQ7wpg
ZbE4j1JE0lWRfjnF4j4+NI3PTrUXvGShuu/HUfwjKXnDDT8WC0FKDSAiz6IY
91YnFQq846gyyv3xxLUTHVJ+kUWSqXvLoxxtj3OIIEYMgjBhF/7cqL5JAN5D
6Toi36l0wPNWbKyqNfGHv4wERAsGRVDJDwx5Z+KXtpAvXSMrRLRBJgfSFN59
zNJO04OfxwyU/MlnqEe3H4dy3q5xNaOZsFVMa3L2P3aGPKU4H74oomrAFLhX
2cOrd5c+vW5XmnkKTnKQvykR3iF35vQT3L8NrbNyOP2ELzYLxaOoge1rRt4L
7FyDHDKZMpwf2twxiihyIbnfmPgpwI0Rz/llAX6o8qtBV1Y+u4V/YKBWZZTj
6YeROpjaxGW/IO+FyyZro/r/clEYYKiHq37tHcqaEJto6fot7Zs2w9pGdCW+
UmbP9fMT2edovwzZym+1kJGwGeWsoxHN1WcOgIZw+ilTsw2BsPegzUbG/cbX
02hFQIoASwKp1Z2+MqayFXzPuVh9zEuGNCpdyo2fZ0OwkSb76xbI2HmdfI6+
XJe3c2FpdPBahVwaqdhWMzzssT9OMbuT3i7XyymtqqxiNK6AdG8lh90AEViT
LJI7sR+OQ4A8oV8puYJP+qprzSLMcgX7tkm93N++kLOXaeb46cjGQNMdpNkb
hifChBDPebkvS3iLmK784xPZJLoqtBU7pW6qzjuM5D/daDp44vs2r/PV0Xak
kR0V04JUKHGLyo76VtQh6R4rEDSkVwI9LHqXUSTt6kHHR9uU2hxJ2eTwuvwP
HXSjZbLHZMfD4g+qf0r30H7nMxVOpcUPlRyGMNLix/o6+VcbrbgbuMu0OtqL
zPZsdtgoJH8TcpUsqh092W2crp9lJ9OjqvD7jwRP8BMxnUO+tJKtpnON5D6y
Nj8tZ+oGDS45Jnh4LAppPqumpiUnX5xpNNGN5rat5AoFNcn3GZ3jAD0J6YDa
htKW3X6wQoO9uz+GxYUHonCn4scKXB8qI4TGfE5HiO0cbf/b5H0LGFASkAgx
cT9AtSIHJKNawinYzVqbBBmRTEm2Vt1FEJ6cvlSLZIylFqpBRzIaVKlxaCrM
Ee1jrVvQ8bON2Ktic1Ej+x6xKc3ebdqyoZnYAmRP8SzbMr0ujsRJ22srb4Yr
0camwAPPOw42uGeSHbaZPrHR1CsuS1coNOXZqDsiGx5wtXnVetDp0LdgS+BU
Y5KGsitsGq/LpF447LQDv9/OnLBU8NeKtQriAVzgpmY1Ew768ScxJnKaqRli
r7LAThy8EQNsx/uIJydNDruSCPSzDu7QkZfP1BWQRS2OAG1r9v5jb3FSIe0f
BJbWwKMHgGfjcWt+S9436Tj2C81K9DU9LvGXob4rYVcZHeDV4E3iPwcp8WUr
3JdML1BAWTJlCz9awI/BkY2yPvqHmaYO3+sfQpn07nbILX6cWEpnYNksUT3M
VD8J1aRk4kS65qlhyJWgE1Bv/aEFF+tse9r2Nxsg0lnj3nMnCzGBCwk0BM/B
ZOT5wIhpjakzGGXKx0OV/Y8IiPuU3pNRhdYQgr3O6W0hqxHNxiFoXrR7fbDj
QcIVpCyDHucDyJp0tclrzuDMC+j40ip1//U6OJ5QwudgF3cj/MckQCwgLW+9
FZsQBrW1dPN59e9XzVDyJFZlwS8cDhpyakbqeUNa73Q0yFjkZca9Jw8xH1SC
Xasz86nu+IK79Q/urIHvWqM+tQ9xPO1f5Y7JAjIcS8MrdW1/6Z1LCqWtUHgo
FcD/MHEhAqiVU157sJVDRF3EnOjPuqF6J10iBWM5xwQFmxiVnYkFvyLzhQIU
V04+xcNW1fruQb9DVHTlg12N6nm5s6+7Red1+jk0tq5VZKnCE9FwLuohZbO0
sc8Yljjn0s2T1kU3CnUyiI97GlFD43S8wI8LqmyT/ymgDDxUBRC4rOoXTAB2
ZVknRs0TBNDz8ktifPkaxLKSLB39AKmBMujLWawCPiX45Ayi/24h8iIInyM9
3Uwsk+IafuptElctDhUgwUS0RTqcuJWnVAM8iQHHOojTxlTDw/aFgnZbaWRK
QBhIH2NDzMAatBOrMG/P0IBR4RlqWVBjB84Gc0DEMmhLdfCTVAgQgbvdsPA3
PfBn4dN/qxKnhKluI0sPW6To+ogm+VKypGbTnN07sFqPBlJbElP1E66Hrosx
i5u4deVl5iEJ+9NcKuql1tkLy06U9SkVXikglaaFryr/jff5XvRBBIS27YTK
188ne2TvXbCF5diiH8IO43giyv6lkxJAkSLfJWv8z6c1UUzRlVxqmzlAIoLY
r8IjyqJSqncMPAmCUoUAfSaeTDUKWW/5+YzHjLB+gAxQlfR2ksBk9/UsTvpg
5JSyLVcPk8KFnNA3DWYJaku+Rdn1juyMP+Qns+uxUyIEgxcQpOdG0lh8TdJf
ljJ+c+ywfIdS/jXOcTzBkZmYqI64/MZ8aV/EJVtDK8vJYldqUZzAT4YvHMWj
DzxVimCqkFlDCUtnhyrhrrBCKRThFCM/QdUxVbgmOkqSzWr0A3J8J7G5rmKV
Us9ZVaDMFlJ1TeDxDtY+OTPD0UoM76057EPMBbLLBnLsa55Wa76hnPKpN1jo
SSnivvVmMwz5WRx4bxYxHTNiFw9VtxWFxV/nfgRSlT1NvM0OqNTwaq+uB12c
jf8pQ+9aoM0+hL29cljrgRrYFfWpSSk07j1gu6S2y6U1SIiMxcK21JI/J5ho
i7psx7ZUWiKsmlK5xplAxb5+K3Dk2gHEzF0t6YwMroto+M15rv5YQocWIt89
ZHnSJolItUemnzIbExsQbEGCLuKNfdhhC9Abjh+i2hWPtg8riwA0WPixWa+P
d5lkI3+BSk5ii/rUYEN13ai0F53Zn0Bxa5HB8H7LJW8M3d6CHoj+knOD/Wvs
fvSHdkGBPOjWHt6/v12Ov32pQcllPoFvAwVV3HApzixufI4wNR/EtIazjhio
ihbzN4mtWR7KVSFnPBdagm+b2K5SZQ1R4Ujp+2h12pNJ91hmv50dyrXJ4xlG
KyaNB5nYSG+23nFkWK5XWKcWx9xVFErqWQhMya7ACV1/DGcuc28rKSRde0BI
lt3iT2tcm0/qXRzMQEpVXz4PSfwLn+Zti69tYYefz2rUQxnD/EkMu0DV5s26
u40K56LouOzj5gNoODbId0pkX8VVaEmxJ/KNAc3NqzhYECedHdHaTFdyN0cq
qrx6oUQG+mDG+l3ko65dYPu0dk2K2b1PM+XvKVGPzAksEGM7YoW9FxFRubQp
A5TB3qCbl1dxYnWNbUebgAC3JUa2/x9FSlsQ0IVgYoiv4hk8PpCUkyRMrfyV
tn1zM9uzAojG4n1unA0Vn28fNtPoOVVH6RZQ70/j1BUFdLTtg8Zf2BfMdOY4
M0sqgKCIvw5Eang158pRurE4JczrK9q0zX0K34aSQR1JIY1qrCAjXQFwSf/d
hwirOZUbndgMxEQEGHOlZxyHot0NkZEwWu/LBoAp4Lc4IOISWGvXgQk2xYUw
gI7fG8LluA1CkkWHJ6MNTLqWj+ttMHHSDDQTOmKelTasKXdEJhiQEdKq4MuR
BLdr6w+jac+D+YWcwMvkx9bK3q7okUpzLLu0dV7jm+ObuGKuCdr+kOmMdPDL
9adiMqXvuWbeAc69jRPfFiIrVBZDFAW+CjUeg9et/KC28ypXIxfZVLIOmhJ0
DDFI0zJ9unqD2w/ji11FuQYg5zJCd18o5ZslDYywbPBAZhnfy0DGa6Qotqyc
t7WIeToVK4VmaWh4W+6MeqiDMoTrzooXCKvw9A5yhxUStyg+DFie4fyuO9Tr
NLCBteCtOpCWQ8LLtVjdsMlFY87NgSaaHqBI5iHhw8IX6Q1iWLsN8ZVG+uyl
KwyNJGoC4T9c45y3aa7xqNnLnGcuZat9yOsAK9+gmqU6o5LwwfE86xH6HvbE
4cZI8raKaO4SDsFE+93ARzk9iPO+Zy7czYb1QDrsHNjjsS2UFPOxv1HqTSWz
9swhpNDkZMo3C6uMwSMJScU4wwo2U9sDgy3W82LO4qyoKLA/fArCew6NdL8I
bEityiHyCHUTMLXYYos1/eQvDUVeBi9fvXlreYeH/1pSQTSXWpyjKIYXzBiE
8LsKtSllk+FJ7f1oWaPasXzcnevSwwGg8oH7WAArVVh3/HCOzoLGghpcuX0+
Jvz7npgMMjxYdDatD/t0oFidUqbqv4KkedyreUtnSMwhhPhB1AuYxRISaYN2
kDoMpJlYHeXOXvocSjky1kAlggg5sGUgTqisnG7P5ThfcdhozcVs3v9t4l6J
Or1Ceq7fWVUuhRNm8J3wRLy2jh3jNAHjaPnp79AwjulgEMfE88wQYknTV/3u
Hcs8Lc2lkvL1YvXsePw/949IJ/Q+xVTRCZh1T4fzM+iUzc3fHrF3bkV+G9vO
yxhVVwr7El6TvnMPF43jSYcVXJQv+PBDTONs1EmsGONRi6/3L6hU6fXH3ZYC
vkRw7ipsKmVYtOxxqMDYiwWfjeGqJimRxfxxd1jOwwTbrcIAkse8nJ0iJ8Pj
Qbln/16ZfMV7dyiHEZP9dil6vbX9XVZGPxwnxSL+UD5y0RldelJrR9XrTnt+
msWY4wuH/tLFfzimZIoA+G+r1ZFOo//5j/WVdJ/VtniMKfD9fYdIZsEJmgYF
vghQkSmqzSMGcEPBnA2srI0aC1kyUDombf+C6BjHOS/x4TnDi0STiQvwqD8G
dK3zw7/EU7hlRqg1sZk19N2qQC/Ofj7Q7GCCBEdpN+xVxkN4MpvuApWWomFJ
CA/0gSt0CqJqSdzbJMMOqmb+pODBJA9hyK3HHjaqiURkK8F4SpqrQh5FrQVl
a9p6um+03xTQxqT8XyfN7pgFzp2RsRrNihR8BoZqybEXUVCPkM1fnpkteCxC
JszDHIJpsg7vHjIe0YnYYhi0GyqTDb/h/iXlB9SnAXndJMBhSNyv/+e9pdVp
0cMuELM34PG90ZVoifV7Ev47fDUCNtY+3mCUou7FQVyTp3iFrSFyOLtsfrma
JGcsVn0MUiNSk3X9aMq5wUbxIGD0Zl7J7hl7OQ9VC3uZB/sgAeLZnVKTd2RH
1K31zH4Bhb63vAWqR5Bv8QqZEcQM7F3faeGg0mdFglKDHZf1xGLry4MojAoC
0HJZavZkfyp8I9PrQGOfKJ6FOXRNFmTsNC2FZoFwmOB8YpDRYlgGvzFSEVGg
ZfOxFKPs7qqBq4+EZTCXsHSFwKOOqZeXoqAhQH368KcyZrwafiImweWg2Dvv
DzrtcIDYLdRyeULc3DbwX3zmWooubbTiLUKXgKqeMmzNZ/c+qwJ6/A/820wb
UiR/Utwv9sPloNUimsqUzluCrPkEqfcs93SZB/MhDzJC4w2HrvnY+ws2dOZo
/QFeSd+hKgDzjeVh/IibDAYaGw0HPbQiYSVrIRaTXdgLL9QOigaNBhlV4Kxu
XII9btUvcr42ji9F7SkNLlDyx7BQbTGINVwVbEoGHEB0FX+aHQgK07+q2gJf
xAOG6GpLJDfrmimZMXnhs36HWF9q/1gaLNffSTQmaXH8c2g5R7pPNc2rjGhv
5ydG7gpiLp8t5CxDBdms9ERGu+yveCBng/TU1KPbzDMhxhRCXDNRw2WdYI5K
XDMAhN+FNp3vVWGISFzHthGkVg9p4Z2GiYBQj0l47YkpYOT8CbdyTfsxosgy
6ydnBRxX4zQVLIkIgKrNzpzvleBPtRxO36w6tMi58ort75rS116qJwKONsWf
8zQRcBG0hAVPre25OMlgcR/Q75n0ARP27tYUp/Uv+HJutMAfsGdjONoa+dGA
tSgcSYDVbeYndwXFH3iCWR9aKlI1i4JZCboSYInRTxFW9g8h1AZaCjbJS5t3
q64suYiQ+C/TPN7u+R+5BFaRDdmM8MOSPjZv4SyFUA7dj+iftVfOdCmnWmZz
H04sZMP4/Y+5v1BSLlw6KC1tuq7E3zpROFO1CNqOtnC+VDjs9ABfr5ithVJQ
GaqXMQWE84emy6Jc27XjLj9VQd+4X58n1vPYwH5E6dXg6kGkh9/8yKXTmSW6
DI5XneDutudvrKeQWgE1AluBlkVjudy6cb3K5WcCpW9P8OTpyB2u4MHtctqP
Qgm8Vi6vXqfsGI9i6cuY9Q7191YZGllzHRA+gNXLX9eLevj2LOFuyortdOe9
AuClpy9FjsVNII3okR7xqZ0QnuGw0gK47Ns/lP5nsc/aKYxb+aM8cWaL3RFK
BZLORhd3cNzmE0Uq42X9nFm4EyrdFdMOo0gX6dkFe5V2/tIy0ahTRez0uPj6
7OybcLCpmgUROjbCd97kwGCjT1wBXmV5cpRCUB2RPjPDgCjkm0h/O3WGg4Pf
xMGchx6BMM10Rj9k/tJLnnijeT6F2P7gneh3QL6wQbHP8PTJs+RpJoHqr97a
ZJ/nCQmrUdI9FsmejHIZQOZfRhYAR95RGCKJo7cjZj3XJIGWPoOlqRkdHyf4
1Jb4cTkbd9M3c7LfAJT3kORygsLymClLQFFoplKXlQHibreWmZbqQsv10oxq
iVhzC5p83yGYR4anK/ANWfZyGgPvEOh1iVmFa0uYg4lsN1q0OQRvL/Z1M0CT
vZ3k901G5DEBomplnHDu9MNCxjJs09nlLHRjb/LSAu8m+SbI0uARnvke0LZR
Ira/pJvPVDbLVYHPmZwJ0AGvfjItWXvGkcEiSEWGw4nd2xHvxxS6xHuZW7zU
eFqLyLtZF34RSmWSA6iNIIhV6w9H+o1e4QuDHloKzd39WeK6Q2HFcDQsqOTu
5xl6zn2u7eOmzOsktegEuTfv5TICohHpRGbZpRx8bryz6SSnEOI3zNI1FxdC
88RnBcvBOmGqH9wh8PKRMmcBhGRvJ/FpE3sckMkJ9tRD9WcE4j2wlHfias1X
OPv+RGmRPaEB9yFWJ6CHb0I/NNlDIqHACr4JbO9qM/NrRSewFhMPKkhzusBn
5nVGp6IFoV055nqXoItYXIetCeHrikhSpvEII1M2+JyZySuwag6NuQtUTOWX
ydEw7TC94qDB1WMg9ZoGn8PICpRtNtT8njczB+8NAxxo39PAD91fhYfmca3R
rnTxH9ypsSOhtWl/tW4M6ZlljF2KfgEoJfovQS+wEkFGObaD2tsbCTad3oc+
9r/rKCZsA+uIXqSs4ZW4LwF9u4YWkuifbokn4yrp6L+Yq2B6vn3vxrATcqAa
jjryKSadaWB/YL1Ute6mAX8OL29ye0UkFye+6YWI6SNukZ/TKnfoadYAh+nH
aRiRy15LY+Nx1R6Hn6uZSI1lGbGb9ELDStv1jDYJ+0rTPY5STccSD099YpQY
JGLaFuQfW/0DcGohEnWmW2yKUCxLXQRVAX3KCSzmDi1u7+PsvRyAr2sl7CBU
bIzDKzx/8DCf4W+U3Ii1/NMoGMFDI/IQ2XBouxI4sFLJ2QGGncYr6Rh04/91
a+0mrNoQuWMba3MuYQD4Jsfw0oPa6sYRlCOZUi//3mIIcqAfbz2nZ98tOBec
c8fs1bKTt4Iql6MFY9G1RR4HgPmL7wJi0wZzwOJbVZR2ahi9069teFQwR7sH
eEUHh4h96tDiH7nJ01NnQrBuy0bjuPHgsXwbZcPpSezEasfu8/5MD4eoQ7Vq
lUxgKwwi5bMQ1paSZbpFITb6U77O2e+XMyXOj6PcfxjCua4N9gy5YlGITIlw
3Mna7zjXiTahR3ulvEto/TuM1yZSqFUAAvFzniw4JWoCMpKhg0xJ9KB+WIjr
oZI5xzzWqX7jg2drOTNnFuG/li0M1s+UCH0e2lA8lPs0qbG22N1Ku3fxi1Jb
BvAS7L0aVAqdNcYrtXPyIQN2gVZboTlfcPJ3oQcX/RJzkl3JYutIevBzEjCY
J8KwSvJFJwQMGdvcZJD1qSzrwC19RnfKv/C20V1p9Z+0JDMZklHtI8XIgnhr
x177X7sG2JIP+Odfihw1/6PNU2dNs4Gj6nwV8MjXmCAOCJ0zsk7T3YkkcXSZ
ato5zwInU/yAs/M1OaJ9IZmXUrsc89iuY2nGFOzeFytY1AmrIJeS7D29fM6i
GV4G9svnQRtApXmWAP0yIIoEY0WS9PpANIkrdY8LefnWdDGAd6IVuCeRZqcE
1jHuwatOYSBH4OgD8WCUH8UuHN6WgLxQOopGYzDbDOfg+kFP3Nwu3hR2rOre
lTA+tNje+ewhd+F0mKyGqlAC8SvRkEnAzIzO4cY4oDy/ySRZ/byB8C1J/GpO
48A1fXH3GmBRk4yXnE3uQhwCytupbwpVZZYpZ5HdNKNd4wQ0Cjmk3NljEG0I
xLVivrQ5uMtB+VbFzXJ/lnXswpjsVtLCiLF29UTooj6lXN4qkHWE5yXnNIH6
G82tHYJBmXx5e+uMzb4+ZWW+Xp3yHolGd+WVbROwQpaiLQgPoFj5kAVjGM1a
l/PePhJFmXJe588Id/FLC2shYJFlzjN4bBx8koSkWhOP45kx0XQnWesvYGYL
cHNmVSj8Q5KpYq6nSsfqkJR0c0hP3zv8tKI72sibh+LXoQZ7hZ6mj9iA3yM/
7uJ5a+SXULiQOHLQ0VbEufkAOigv7dD06Dzppxk3fOhxwffUrMTrSVzwczQc
hsyEtpQlfN/Px6C2kCkaJlSCvXN0ZCHvGVJbdjrGGljV/Ks/KF1X30HjIX/U
2qhiNc6USVBwqJQvm9Ir9tCuYGpd+jnL6pxB3zBtZ0j4YxIMesGu+2uxA169
g1yKkRp9Fhu1KS6qIxZZR3vgjRZ9fDSqD6lcCphuUvdav9DpvjXITwnnN1se
gAw963sAD2enpnJbFBd1+CywTLIVENWHnHI4hbIz7hcG0lnZnfPnPwV+5V6l
lOR0K130J2lbBSyZoXjuR0oy/mKcxGg6CXyJcTZRIHPqfSAQ3utkTIjFK9nR
uCWx9YmUn6aVJwbGEHApFtVBzlWDvuNRXrcIC7/LpLVq2RAVrZEEP+HlzMtb
gmUIVMShLdv+iPQsoRKxUIEcdW4YnnHKJL1pkG/dQDB1wo/p359ozDWUE2BA
+b5Okdgj3LNsyLqVnatI7zXqaAy6vUTGQTsQS3LlGOxNvS31kp0COyry5ZNL
24Z/lodUsWf46dlm3a4o3+/1H9XRjaB3BfRQN+gNdjyr5d2Fd5FXCpalmqBx
9GEkuY6Jv9Gj7Hao6Fr1Lg6n470xO70D1khQbqRtc81s7/pt02ywgAaPN3FH
NNUpK/g/AxtUZyHO/sddixycwq3mInD6t+ATEO6eHuEOD9RWeY8R1tcMyNVN
GOOnJQh5DuYoQulMzEtThBhnYhY6/aOqjoGtqM/OKG3uAtQHYkpNzAT3hcQ4
OoDASHtikt+ZDAw9ZnpI1fB955Ci5Jw+1+2apl1KfRbd/eIlA1X/0fjltWxO
jVQCWzlsgffWL3Um8MAiGNCLQx4q3W9nJIVzMJyLqQkoqVedSBLZrdfOKfQa
y1dQC4TW9WsUVivQ/i0p+wihmwK+4IW6mKz/hnY8VbEFk6kS92JggRp64vbq
c77m0N5qK3Hbdfhorqy1Cvf960XwRdfU5pQwRXZ72EwvBGUemUCldRS4TpqW
ZUzuUWxi7Eoz6XSXwpwZYGpxmuP6nvA7ml4lAt1MR8gOuGyEMRhc8wzFPHsC
j5m0yamHRFuby+g905leWHaWIpKka79o0s2xhShxbXw7fUakhE6NpmXS4iKf
MHPZTcaH8jsh1t5ym72KOu97O1U9QxT40q4eGhRjiKUVf41oZ5Ge0scUXz1Y
3ld7J9wNemManoCdNjXfTrt+JPqe9NqxoNRaNK752GAsUNTO05VJl0Wf1eEt
wQMB9niszU5kaJgzVKLJF84y8r0B321ljby/DD6dCHtDXCMVorPPIovD62Tu
U06mntr0JQY+oYYs6OpRYiuXvOJk5hk+xPoDXx3d6qMLZItK4y9CNw/jsdgO
sLLJyw1kf6brF5eGaI0/fkxKw6obuKYubmN62M62kEt1HoIv7dRkLmCL+UF0
znRCZIh42W5vDc5kmMnSOKPw4M35M5vS3k2PrZbix2VD18DzpTE6/YUaLDb8
JVx7LBqNPVLGJiTg6QEL6+DaWRB4s6uYO3owyUNHxmv6MKVMB6fUS6VjN3Sb
UArUtQS6FJPB3f1no3+fGWTxHTMNNqj/1h5OPsWlOSIX/hUTzXQQxJiNT43t
JL4jwl6H2X/Nklnm0MFIhjPdLUVWIGncQHv5yz2xm/jE7zWLkKEUTfOsSKvw
N4w3ODZfhg0wQPGhzXea/0GNidw/2F7BP4uiAvJQWofoGq4lB4/X+42UaetG
LbViuI0Rtcn23PBrNLvOapvrKhBuuIqL+CLE73I1F6LyJcxL+iAvqDz/aXkB
7EeaqZVG/bXPFVIB/2tTOJT+4ZYP4oC6+b7yu0fUD6H1Grcviqu3c4DT4qZV
rWmbVDGCcsBF3nh1T53t7akQ0SrUjg+Gsq8UuRAmEeZIR4rtDSUP6s/wnPWC
TYctpJn8TiOSxvEcQLbQaRT4Do97DvwjACmjO9yDpLJ43pJfRhfdEI4yOKP+
KmxGaHNWy3jqTYTJ2snUOuVDLW0Kp9nHgNGwaK4SwZJF8U/gJQDD/FQRSQpp
2LiB2sxzcyFrp1DKDsVNkMEf1CXwY0+7mK5GRVgMYpaMTIX3/S6ivJnXp9eX
VDOF3kfNwqP0HI4e6ZyjQdPoYmafb6j9snQ0O6nVIeXxyiJMUzaAKzbm5lg8
ZjOKvdqzeVJ48xqVME80BC+VnfJSly+d6N1Mfxmg+bcqnN7vkytgU5Qty1sf
LwzCkG0yoqvneH4xi4EVUhp71k9HSG/YrERkzejYU76j87PjPBrFzsqcR32i
eU5eGAQSgiKEVn+83WSj5pfYymo6i5rmt73Bzf27K5lZC2XiLZbEWynjDrKx
RjaKicv60OeZE6lXe8x0ljPITGl5Qsqi3qwmCEzQFSjgnFd+NRXTsCQ0ujzV
freqP3qsxJ27xRBuoeo6TH7y55DJHfeeAN22x8lqNH8zVHGiuMwWQ6Q1yTes
ASBmB4x6np5teWWPs/NOc6gOQQLPuNzme+/YmXvsYZIABlJ6ZzcVPZxgIUiO
k0LTokUC84GK2cA37AtNa7xH54lQ4sQiDWqaI17xfeAj7QubqwFbSeLCv5rp
eK7HOG+J8mvRuiB4MAH2Iyj076pH/Tuaf38JyrtsuJc8y5ci2UuwiujaXNw3
zeJ5+WQ47590yqZQE234jh4+K1Q7J5YbC0rKeFOl1zvaSEpHQNtWt4uDC253
ue5KXT+FC73O/fwZM+G9Wh1LYRaVTip/eyjcCvIY6nrpz+R2RVOEQ9MOIUig
O1GoebMuySM96LhMJi0doBvXY4QAC2K/a31AAH09PMg5h7shwrQFnuwVFpx/
JMhHx+SM6xOWGe4Ka+r/39rECmShDywh5c6vrud1atQE2CfpXMDSrYvS2csE
z8pCkWeZHbm0bij17ABKLrogILSlOebiPVVkEU4pDUKJWkov2J7jMu1F11s4
riCBIoRVrSHid5+6AtV9fusKqitE/6CzW42K1MLmceXaD5pzr7yQHbVogqRP
vRY7SkSpiDvW85xivdMLAnPBEPO3kxWl68iF4eb6c8KjXW35RwmDJgUi+pMk
+X2Cr62gTbbjCfZdxmiHE3FpyamCuPtqmpzfPFbt54kVSi6VKPqBKmogZMl2
Fkr5T1kVXOVDJ18xz6kSJw+wnfN94aA9Xbez6ODGkKC1xOxKY8a9CXmuLdkr
iKX0NYHmibWKUNT04JDmHX24s63DvOywAt8BK9sR+zXw+Z6KLau+3E6LDwF0
sNu2zoQsMbbbD20rj4WGQnwCO+IVyd/qy/A2jqhltsRbMXBFWEJynM/J7uiE
1TfDawyoyU0snpKiY+0qZuXlW+otOiWN9OGQhaeiPpgjUqJ+PEwP2rMTWToP
WAG5i1si3jSv7dn5F4MlpVXbS0Wg5mmUCbXfgpY3eEuiqmi+/svT0pDXyHqo
BCa352jiX2JKpSDA11UKVh1+mB4Acl3bJmY8jxHeWvpNJUF2AZfX+yzgAWqh
NBBiXpKzdgY4OpszONjjLOmPurx7dNo3OX7/7Ko7xEaQVikOZhC5yRpU+jHv
OrTC5XSbZakEuHnqb/kP+v5I+L/KJmhD7zXow5yzbfBoB1+MZqK/4540Zn+z
xcSI/EpruubhMQmPVOVcJmzyRz1YassPQKTi6+p04dKM+mTAPmvb+F26lOHB
8cO4q2os8lq1vx2wC/zfsbLhKCSu8Ke0kaW52ZaT+iQ/I7JMf6Hvwxc4CGI5
USaV7l/gv3jMmzNuPO8PEgKqjCcrb7QGj2BIMXzEK1GRvUymEjFIDsZBAtYT
gt+21cRjbVnaZSQD8k3OgBJRlWmbP77t6Fu66bjrXpa6AhXzyCDSGasPcToe
8fvFen+2QxX5vdovpHnYh+jqEXwcRvA7mPAXsbZzAmuB5gCS/zn0LkyhDsFa
5/4hskS+Rszhm263EVD2On0tsiWAxbaJrWG8LFx0p8VtrB2bCxUOduSd1JI8
tQBd5KH1RLY3hhyKYrrY/OBv+57TxlgTMx8b8Y4DitJFdx/4p02NQRjEnQNe
JmiRP442hhBttnJo1jrT8PVK3di2pQkZsQSbCiUnN6ihTqWreXyqBv/y0J7c
nbxhv4VTjkMAy02CVjP6R17KIO4mNOVIhJA7HRhU0NuAcAy2yzvWg8zZ9osO
cvCZzdXH8SC/pCphNmw432yk7y00PHPM5YDspoSkjIQu524dmGdSkk8QsLTB
4c2vaIA1NlRQx3XrNmR1lP7IWOf3A400LZ7jvFNUk5GqmEnG1scan0cxjpdI
oW2kZRousPgFb4JvO4PttxFCQwPHTn0vHNMRju0LSzWgkoiZkXRyNde4HeFU
GDjmwVhfEiwmbwO9CTLtDZXPsB7Vk9/RDlt10p5ugBRdupWbIUj1JyM1Rdej
zSgA3GAk55LlI7ZQjep/NfbBWcsONmS33An4ha7avzkunv12QkUDrrNWw8hB
Gf1+qh/71dv1ktrhxsoVpLesMePbr3AROS2A8KZh6W+10S87RjkCz4fEuZEx
odLMxCQIOrG4IG2vgcqRwQLp1tVdxPETdIuDAbTaCooHVJMr7IcRt2YvNfoS
Y3yCDSNpSapEdS0bsVvsS2KEIW77j/N24/F1fE1SSAe2CwQ+kc1W5hjSlM4u
v2jJXGcMLiRpoTTigW5dr53yMSAEKMJgGbwSQn8qcWiFK4qgLdqhi6vRoJIN
EHsUDSk3y6ZTc+FoIgH2A6FNicA/CmMc2iKE5YBVfl/RZ/YhD/fEll/KJlM8
2Cm/C937qm26L04ln4I6ytxr/nD9WZI46c93bWhuM62y4GZYpsUqnNtOOOR/
7rBPmDKPc3W8j1gHc69XSgdlYT/TcezS7TajSEmvoGiKDC2qlEqCqAvwaYbI
EE2Ds8p0bbLYXejHKERqHeBjsIeGvfVs9cZ7cInWneAJDi7Q5tfYkSjyOCY5
arOIC3WSU+yZUcFMDwkZ5CPekz4htMZc3ZV7ejr0gJovONQuzJVCjs5DgzD2
3pEn0uYn2auBYCI8wfcQ+BWbu1lSnnX0LfTaMyvqoquveuHtsiIFl6hVW2MU
UdOkI6Y9V86L5GCgNgAa1C2TOv06hXJmlAtQqvx3smrN5Ec7jZRnb0NGrXWT
6rQfiLKVxXQSagxv4ab3E6PS26ibEUgKJxlZUXEfhfciI4vx3jS9IbgTlDJc
cYzjgtvnhDTpiUTlRAy6bEM0c3r1tXqyXvdq32lunNUkd09ludkWgKqJjRlD
RE+TqxiocGLjgtqa7F3Lt9ub00Jiw5WdxnTX03tG158OIuN6Y+5DJrE2Jdwr
N6E9eK/k2cktncKUYSAGqscEYBk8tTCdrC6SQ+MlbhlXJPTQ2HbS2hiGUHZ8
Rocb0KXaTEDo/21r1vZ+D4boVxUuxwCsheGm0aNQroeKuTud4QH2JViFBZtI
7R8TEV3D9L7VB3ySxXCo1CsRfgCb9+DbmM2V3R6O2grn7mkXozE75bryYCzl
1B1KGcqUfPsDqlZJEw9y7asAvrT5gMXyh4aybGZWlLe6yy2Ae0IRxH1UCyqK
gPld2BJu0//JjoZ3Pv/3scZ0B5SPOQ3NOexkhjJitnRQDygkQLm1BudAlG8G
sX3XyR0LL0RW+Z0pxB7r/lcyOhYvjvg2I4tnXM6n8q/TXqwVeQThlH3nCmKC
Kp7odW5RlOlK2D3rYgJIBoP3pmBR44nuJU6gejuNnCERI/hOQs/37943VdYP
eNvcclHK9X16Jl66CNziRLRfFgNBFqkY7d40M2kQ0F1WXTJBKi9SEJmFulYB
ZI3ttqraHVLBo3d9tf6iv7sxoZfJOeCUVchkCQEbgLfuePJpykVlirLfkSB2
P+jW320TOvbNnO4I+/BaRVoWuSbndPzkc80q+H413oP8CMvq5EDmJoyfsBlu
/wlDvYtGAYvqppTxSO4b2euVXt0PAczbLnzS63qFHV5anBj9SO+WncN4WmvL
sKRJHfPfn+/bDiyphiLA4m1Qi/6HA0bULcwJkOY1rA4hzhOcgJY+eKhquFXM
V3PiG1355vessRxciWoZWlJ5BcrN3xaCZScRvSnxZ01iB53pOOIhYH16PAI+
uCEbHBCayHTf8AkDmrtedPeEuKRqCU3J2XFe6NV2veTm7eFFVlcGtCLwnQiN
Mm9xdj8U14/J+T8XsTs2me3JVUnzP1j8HGbh5PHiFAfpUmm9mcU0DZcdI2tr
WGsLSbq0e3EIP+oxy2FiE2UBSqSeekLEK85fDL/OyrtU+W0I8NpBWzV02ZsY
SpVERxMoxDnUr2oT1I5BLYIP9Pw7PIcMseaUddEBTSsLwPvd6++g3xOsgMMM
MG1oP3XphxYXCrEwSDXahXNvN1ZoMNYENC5BViGPbH7Vj7IYHaza8shwr6a6
kqK6dIWhRQbU0IbKW52hXqZQ/Ua+Esq7kMl9B2ea2QyN7c55mOeCqnYVQhi9
uywJEqOiv946kvVW9Sn1pUyW16oLkt/iKfzyA+0IYAv0P1up1r1v7lpAiq27
7bRJlaC3tzyDgIzLICnUUcCPUhoD+LSoO5Xl6wQwkQTWD2Vf+feTd2toEsX2
sFr0e+NxN+9Od/Vj8W0elrhadwLnig59wXAhrcyISBH6K94N3BVAY6k04dHh
hF/PCVkhmb+AHRMMrArI7QML3XsHuGRGDBG4YvuYe55Taa8R0J59KfHkouW/
VjdnBxvz4px9e093bxaEWnzDyKZN3iybmKakSoNlnkool6NvLViyJ8RcCctX
HdUaZAET8tK26XF/XZNdROGKuqOodGn/YXwDw2QxDm4Oq+DPA6xAMADIQyT2
PeFQ53DiE7kCVF4flfqVDNmwXQtDj6ZmwZY14PKz5F6HZORSVF8/u50+Wai9
CADqjaDQLztOzY50XnIBWOPPVv5J2GDeu163jn+wkNHhDg8Cu/NemXCmXiGK
3N3WZfFmged/mbxz3vB+N60WQbgzMtqOI/b5v3fIP39WyoWDjbqs5/dIhD5x
ZWIUxfTv6fakNv7zoFLxVZV0i9ShuSKfTx7646yYnDCgGibdpiO0VlAyHMZy
EMHegFS0tGzqZwAsLE3uXzyd+Rj/3J/4/4//EZx+xUl0jAQMDz0Wbg8xnqeg
8Dl2nidMNO/iOVjDLefVYjxDDzrqBGj2ezR3m87jLa156PfgOCiuv/nm+9Sx
N+Xc4FCtNBDS2FrjGGoxvyjwtaD9C5gOVWKE45Hiaj1SKYHZdx0RDLc/rfps
ZYIxMWFKZHwqoVAZfbnJc1f5qrKaUwAp+9+lQTumHZlVWlohaZH0dE9K9vs2
P4DCYalG0CvkwLJMAbdEX2z3OU1OWh36QHFPHDMWWSB9uMtLyr4hTuJK7R1R
XxhjM7CNDjmP2zysQKJpx7N2yZn8YYpTJFLMidpiORUhA+VR7ej4m3qiT5TW
vVNpgH51os8DBpogHleK+1AF7Y2oyRvaHCQ6QckXflatzZYah68TM8mwpXox
GtmY6Kp4GYXFEj3myrXC49d9fxI7jZ9XH8sflLjhpaleQ9tla475r/Kkxwhr
Zg3bzuvOMtIizI1HG1JDo2IM9Tvb4zYZOLDRlrNh6N/hxdaz9a5JSiyuFzUV
kAp1KU9mEFyfAm+TDMXAYey/2JQ4k3GMYpcGUpJvgZg3SXu0rrmuetR0ZYnK
u/4GGotFDh2/Wr/2ci/MjXFVJY+A8q9D5m6/lkCfYYpxMATmCT+YRx5LNiSB
hVOgqjeQNkpUMzYg/P1FFTNKxdTc/9EhnCjva55zA0AqKhGeqox23lRWZfKd
w0IyPA1VdYgrQ0rTAGEizbkoPWwmdjciAO0+AAjKBMg3YwLR1B3XfBLhWIL/
lCdxPpQDslpJmTIlbdwrk/Bf/VtPxzdxRQVHiajz+FNW5iPVAMM92DY5hIQL
0YbhQWzpJSc7tx/qiwN3hji88V+YSCQEWdulK8quPqpnmkZ+EnsHEbcv690y
AxuNUS4cqjas7ReY8ihOB6PNaQnbYeheBiAzRk7OA0Busp2+0TRrpt/x9sxg
4vhickdXl9BnPJ9yuMWt18km+hJfpUBrviVTnFQj/gJ3kdvlhd2JSDxTuUUI
9U2zZ37Qv1pYg4a/CsABfzrsHnHvkg02Wlb1bO+L7gb3oNvcCKhQ0PCbesgE
hRv+mkOOc20YOM2dw6L7HqZ3h0h2lUUQ6fzVkYMl7ayP/LPThrV8YXF+Cfy2
DFOtVSJ78LYt5pITk7eAs/ns8XhMOOAkd61mP26AlYZ/X/ynvxmvrP5vV2j+
OnLBppIqrF9aNfqZmtfLOwI4Tph64+KQgQJIihNrmflJEJJ6CCQs7SYe5apF
pTFwDbzhazoS856Ki/+MmWhctjBWFRiO2oK2EKNXoSyadwYt5xnlB6ASD7iT
KsatuAR9UsD+JBcTdAhNxdPXrCuihk5ckjdSXpNuSegnrteO9/XydxNOUsgP
KSJSM1tI2HqrJn1fzOATQ0pcXM8w0fhhO3kZo6EAN69joK+PwY8mZRwOHgML
WWbnXS/BPgx5ZHLYdqWpiULT3RQTjS6RnCoItIEiLmAT7OlYdDoRqj6FCYff
blrIuy2NX1GcrwUPbRt9y2ZHzJZSqEDh+wqJFkTi69ueVlFlPz37tjwIZJfd
eItRjBv2i4G3R87TILj9W9F32T6eBW5GX1OKYPxhrqOf55tmzZpGJrv58F3P
M/r8WpcsyftF4u8IewR+k23qU17cXCOtudbvg2Z/HzHgI8MI/XS6bUAfd44k
/kxHMhBK+DXi78vmHay4WHtfhzW+pRKGw5Kx1lJlHiRSnKXOXnLVbAwKf/EE
iVvyvWZWDe/N/j2rc6f0DltemJOhbBZ3vkevc3bulkpW+mXaCk5ypscRHo7g
b8tJbT1SMKNm6scDlEEY/wwI8LhHBI4o2chVH9YK6FdAZJptmlEpChAZZyIf
UrWFqWxee9xd6WR7vH4DfPIX14nydTw3C9Oqrz/iA1e0IrSGeFfADBugT6Tv
bvLBvFlyfWCM12R3BDkrM9VBARgHG3gJcSp16TlD8P81puAFW/xzQJnK4HKh
ClH798voo4qc41IKzfDDTwhnvtf5yxZkUulBC+IgVCXvlF29nzWeS0qZfJ4u
Lr6qpnbxuu9p2alM/eOiT6Y/7O2Hb6kkJmrNP6LSWz8zI1pip8BSbXfQbB0b
pZ67hHA7CMvNRujVDHd1JE/t5eKB1S44Dp/fQ9SElumgmnl2DImwW9nUdtHN
QCPFZCUXOxGO87Zj8zIZS0DJhmj1KG8LR8pHrFDTZZNKrUBacncOgYNFAnPl
JZ511WYG+Ywby5S12rTQuYQpxff7Ct1gZheciVoXqRF6PynHB1SJI29XF8Yd
rEz9rjILHT6myFkHS3IWQPK1qLTFZ78X0q2n7ZirzZCFEo82vtUI7JTIZkkX
Jq2zpzyc5z1K7ry6/6QsgiauxMM98/QvfykZ6rS2fit0mY+PxClodWZakvHg
fj4N7ER2YQJNKXV7TOKmMQjcqdEzB3RCEZ5fwjvxblQPnM0eQAqsaHLsgFYw
IuLmBSFVCGH9hh8hapOamqg7dlLO5rCjNFea806yFEehwUJLLYTvzi2L6SfX
1K0co7Iz2DDeByV5F27SeiSeY5LdTMYx5phn0A2dCM2QiIJY1xetFfuEpF6x
+FC1r3mlMONYAZdULArvBSoQo2Mjpv7vP6/uYcBgJxdm1ThwxTzegKq/WMsG
3oH3q97u83WqxFygMgc2ce8CUvsNnhlXdrTnlE0HlOnVXexHjkhOKxqNZc+L
6wW3XE8lEUXqq5QZY2hzvr5jvYPgSk0c97xwqNpz7zYh+FQY/9+TSk3dRxrK
pKhF70Nk4qxK8K2w64osZlwUmWFHJfFGs6SOGpgyn0Moa+2/k6h2Q481mGlV
4lZig92n/+7YHHNWmVEl/PZk80Mt6Z4DM+Lf71ZIMeL1h1qmGxirWlgld648
QiK2ZGqsLePJ6lEb8fMUWrT4wP1JuvZgajAFly0o9joV+TgB69U8Z8HER8VJ
LurfjIOQLQVLWGw6fY4cR12y5c2bMnOqn+IrWCm9aKt454McSEHOHfSP/fY4
E7WLwAYvF0sN48qTUr5jptYvhJWUrhQfw1IfJtoMI+M+PJI0vtxZaoRm/B1R
hJ5aOjt+geWrRrkDqRsOb/zMuln/RaV4VepADIVQgdeOjOO55iw2aR3lWNLf
dwfuNgbWiDN42jHXW4gLFbF5V2VJ39Wo5NeUkGAw3mC8xnuGWBRdamM0P1KA
8Y5Yfyu+KviGd80rIoZ1jrnSE8o1IEW1cyIK8zyQgHfnuovF+Dop8ThNGDIz
vn/Tdd3GMQmVszFK1mVhkLbsGcgU67tod1dMDPrK5dE0IQzvLAPUeSLkWmaP
CXCIdvaDug8FjxDhevlzdAzVTYJAZh5rLQntsy28k/KAhPH6deFodj2opIOd
Q0bb46zUKswRvNCQ60ibLludKi0UkD4EuTyvZNeNM8ejD/tez5foGAWlZaPl
jQo75w++bw/XsA58U3S8Vy59D3r6Pw6Mw38zp1VCh/0+NT+LTSbvv55hmU2U
3BRAP+bfTc7Ef32hyMz5hZX/j+j6tjrVFSWgbasBxKtw8rmSKeLyKXsydxuP
qCjOhdG/kQFfbkt+fc+uyRhKGyutDUP+Aq4VOUww6forx5bC7hLuvSnrGFXA
lMM37+vn8hmzQTKR+a3zm+2ABSKjoYWGYjFJryAhBAf+6IL1VpMX2GRNRsSO
Nb4O+xoeVmrJeI8OahljJpwP/cZANYOnozv35IkMzeAeD84nYgPR6jPfbjI6
QINfNgTY7C0W9HgikT+OBRzzS/pWJ6vLIp9SiekHi+PTKNrcjh6pWUaJtuYB
8jgTBN71uLD+T5Sft/RNeor73FjjweDflQYZw0cYuJ5xbNkJe1zV3GFv+Rn9
xGYhMnz4sc7kbfOxtp3tyH6R9YTrHJ4Xk7prWXWlSozamVjKQRKLVFsG/ts/
Rd/WlV9Oy97ArbwQwxQoXWNSXLGSDZcJVHODACVgkiMKxfNGFZD+Us4KE3Zp
j/7FiukLwRP3Im0ZEYLENK+8KuiI6ErpkEfMgURBD6CRKEPtKhuD7M6FuN43
16fWNP7N8iT72o23VVGedpE8awjO2T6SqBXxIRNdamaoMPQtLDPqx1sV25Np
1HOYZpyunQ05xEIqJ06FjNVrum5ZZX+vTRTB4oUUi24Dzg5CWErUNMw9QZB2
MW1tZze8n1Mvl3+4mI0fbASU6qAK0wIRJ01jPZzORmDVWSgcTRIaGQpzxN4J
rRa5KmEQhJosToPPJlcgGieIG712SLzpSkkKl9o2YopWsxVVA4gdkdr4zdO6
vDk5k1gQi1ZMZDTi67nR+m9aCh/o5RfJBEXT+oXNceY1wwlbVBwFS/lmzLZK
K5qEyQFkGdK3t60ZHG2V66kVXYTAUQEFRnBNzLKJ7idwFWOVDP3U9/v4K0Mg
AYqzmYPrN9r+jVk8NcepAqAyhvkanNYKY9Bpy/KmBDSM1KPMBZfOLpenVO85
yjI2rau0oNEEayOziYDuKSfYhOLgkKc692J7mbYEsnnwWtX6J0vJrVlcCc7z
LtyY1eNdH/Ksx+wRJUI0BGiu71S1x27O7tkLiUmh3oR/3P1Oz+4Pjd0b7qzl
Q7w9XZ7WA8f6FGZIKM8ebrQXqEwhDX6eEMkQJzgLJPao1+Vp6O4TzdKrA8BI
TxMSyxuE/X742ZcRZ1KmaT9MQS8+X46/orND51UfFn4LCEw0ovxznxVeXCNp
xHK7pEn4FC1SkHFdmgkuASoWOBJIw9r9EOrjRZWbxF3it5z2lDPU86je4JKC
zfm+Oyk8M5y/kTPyf/X40n+XH3cahv/W7j7lbomugfG7x6eegbf7ZZ9ovZe7
lFfx87KM8i45MGcd9fT0gw1pv5RWQbD+PHHcdlmKFo2/aoVgTdsPNLw6enRH
xyTyuQoXPoVs0Ub2PoLg+Mq9KHiEkq8cdbsJgxgyusA29E4XPeRNIrptav48
9tL/f7vPHa4LfU/jrRa8W44PWsyCh9+WZg/nau85iLm7Hz8w8Mdw7g6R/QgG
L8V0JtA3OEWsyC0ZNgKTnlvALOWDLbrXYZZ0CsjvjyBy5IckodznwXqFcZuc
hrSoyqWGdt4x3gyzrncuU+mXTC9IRlwfQyMWiOGW6BqrFvzjym60xHdOqVTi
YXgZKBb+fKAnjiHXzM4Rf6ldPkV3ewz+Brpgn3iOwWZ/pgo64R1hVGo7xEQW
EYkxWPZgygsvbMbWgpIGADzEBmIDGTTrqzvkgINuh7m+MlPmGK1wQhCi0MEy
5k3BSbfzfT3zl5Cm5AW92aSWnoA4TmGbjLO51qTG7uianQjWcUAKmdewrB2R
8YF95i0I3jjQcbDtnn6lG0tuezGewnGzeoJ30nld1QCMq24feLa1fZsIErIx
Ek6QMB2c09BJDp53MoOB3O+gEc8Wnu7Kg5e8/5srBIRpEp+4hh74IHqrZpEh
kSoJLRfjPCi6Y79Ao6w2ZPCHh5Qzu2p7qP9mOlY3D1UXrCmLVFuhwH5rt8r0
cpf8EOYtL0U6D0tNQLvZOtzVrx28tBxkB3F24JtbQbS3TjECdCGgxLZCXxbU
bJmL72pJ4UzeEIvHwdeB8/uWqKgLhVJPjKr+5YcZaYDzRYIF4fkpxPeqvdf6
TAdHV4QPkK/relua4l36344fGL6rGDSCeN2+KVRGvFkvhxGXL0A9nATc6w50
rGh2g6WT64NnMpIkSeRPz809zn6gtzV73ujcxHYDRBtsE5Yu3UnzGf5Ps8HA
KnDgUHQfqvVL7l8Ze8/V0lyA1HG/Am0Mgc48BA37CmJ2IxI97jn9jjsCuxLe
1yY1fgv/Td/5vAcnHcjb4Kx9AaDVGbzTg35E+cWLvNvtm1VIVjMbRMPTeSTy
LxjjnoAu5x17Z7lIx7ZsgPLPTLjVMqy+788TIn8RWaxdGuD174EX8lfp+Cdh
mgxiYOWXxNmV2yTxvtf9V6F4/tSAjT4O5JvTqDNUQU60BVrt0EGnkEPwF5R3
y0WOU6achUWoxJVuBXfBUihINknDGxtWPnfqQWtwC0uGX0zd+KjwRLEqPEbo
KBn0Uxm7W3+MfZCiyH0PZbVK2j8aGG6823yKY+iaw3AyVfLGIJ8r1apvBAz4
mucJl1TGeAZqNBs0MdOKdzmkBeos7JSiqIPXXU74aSSQAWKdM3qqB5j3A43A
HjQk9+uBu7f5/1ffVRspMlj0qBSSpTUXsKanZx4oKwZYVopnHkqWs1o0eZvS
oa5K6LpRX3PdxHg4VG/ZSIlSa6JDyOQtXDphUOl/Baq3l9NUEgMWOca0P3Tn
AQWX/S2ReKYPhcp3g54R0h83OV+WyOiS0d5aYxYCkMSrrQpSBP11Hgq8QZcp
JtCYjyi4jHnfKyPDCSjybUT0KdXi7Hju+64GDM9B2Oh9/MZCJc8fGflvdy5L
6/JRNCyaym7P12PIEFfESatPlswNGGmZvb0yj4+g+jDu+c2zAM5X074ZkX8I
mtn3zeRg0X+VWJT9WxufOHX8Kom8VMujH1xlpVjgiVgpO6x9ZF+riL+bCH9n
/dl8nB0mzBCFRtqoORPKb54IVGoQOiz1WdQl08dphZGhgVV2n8JpQPiYgCT3
bZGLI1q3FAOfypkMA/xq0x+wRlmUKLkZtJc9yxk6C8H8tfAoMDFvSgUnnwWa
UYlPcFuiZouOTKaKBOvTwDKO7ChDOuSpYR6ZWO+kAVLkHxI/YgFiowKwR4gh
WHZBZpZIWV+O+0gJZEh425Zx2XtfGWEAyC3f4cy+kri9X3sjeepKU5X1QOw1
Bz0RnGlLPOs5saby6UkGFBTAXY9SUTMd/Uam/Dea+czvqHh3yWwkqgU3ReQx
a5FMgyfI0EkrkAuXCqiTD0l96ySu1VgxyGJz5BPS3eeZPy1ftGQlA5ZUakec
H/3gQE0qOm0CidJSLKxvadbU4pDRQyfD80vDV6dIK45B6TA4f6d2bsx7sbSd
LmrUx7GVgCe7cgpPdqwpz8K9HVJ4xQOc0EbNAi784diaUUlsj6mT6I08YY8y
BD7tvs51M2msOQT0T9ffZ4JwsHYoTanGaOdGT3b4+Vl3/qF9iv0l/CHrCzj+
WRe4QGrJnyIp1vvWWUMGOEec1456QozBsJhQri6Eheg0XICeCBblbdRkhtbv
cpoqiLY8kPe+7S+6AAsEcZ7vTsGhuGzhPudx+rLMJsDGi8zxz0Dq/83BJu0f
uhQ94u8frc5z7lmWnFqFpwutv/xE3tKni9Y4sc+6HXC6jBfq8FvmBF1pAPoh
dlnLYERKY5g+WU6sCpwoan6dcQoTDsBeVWOm+SAFNFh8ka+OubpmOtRJijMn
xRk1lVbC8tYi4m8Uuj3LW1YiVBUOyO9UyO+GkFQ84Cwd6o0D7DqDDe/+7d3v
0x8ijdJGbRsk9NkVdpyEqExtENMudmI6/7WrOMyKeLdQLZ1T7NMT+4wmTb5E
kZfI8Mo4JIPNH67YMyHRSlTE68znH9XKkkTxHF2aAbXN6IOSCj+tOSmTz7e/
PiCntaPYt0BJgWP978m0UdFBSGTVd3mU7ohUGMj7FLIoTL+bvisv6AVOK2EX
hEzSPVSjfMTAj7jl8G4qNf5vMH2YEiDK7ShmLBnq5+jDIZTpyYkH9ZUvHsfB
2s1dqE13iosuZGU8ZeqzFo3hAEHWQPtZEW8Bz7HnutSMT1a7eNs2CRqB0r+m
W4L3tZkTM5fgvqA8fqRGcxBtyMomRvsTHGaXfB/7CKpZt1019gv/Px6tgp4j
U8JjdstXhtYzZlsUYCwOVlzI8HjqSdngrthLBPwZ+Vh63ZZHSHuayxmBejdD
F+HCB394JRYCLrZBhnoNgXtpfBzth0z+21jaGGY8XWm02wQYSy8u3eKZ1GBR
J5VNfY/NIgwEcAuYtQDsbO5swEVXA6t835PbKUPZlaSOeqTFn9udWYJx4mHk
Hxu/vDQALr0NN5vs43pRzO1lJgCMR/ZrkGqUWohSihmWut+F36zcHHNzTgkP
t7Tkz9jvM3RQG4Azy1hAS6jkLHfnOGIG/Y/RDNC/1xxWx/6R+7gfbhWtWCTY
xDMfp/iDXEIY0Jas6vK436/lQAjRBBRAuSHIUanTtcTGE1ugx2u5jJU5z94t
y8dirnjGTeAxNQMyibJiG5sP/laYDFxufvs/yfGMyT5BqdbII8sEcoTPlVaV
r97xHxdrVShHbRq6jEcHLa/cLypJSSvEuvrLiI91OHJqSyp1I1j/3jkfs0AO
PViXGVzET5WbSwbxVEGHYF7Q1rOna1Wp6U3PkJJ+Se/PBI4ajcDLivy7kHep
0o/fAt+SRr30FiVsiOvh+hvoLjUL70jDzOLOuPaO3STxlLlxQ0AMF4TTw2xX
OQy6WoZZEppjHRMYrN3DXKAuzmfUwUREuzB0So6/OeqhcpnDXTvSGNB9r9Sc
qYQTzNUgdMGwqPndGHPSZwaJKfmsLOviW12ZVkitQ/UgGpp5a2usr921pvHD
A65Bh3xLKalE/oDkOugCq4PI/f9VLD27CvWvS9WT0/fvSJl1FJjVUhJB7eUe
NIekTXjQxHS5xuR3LkFwo52cvsKbgPUG0vNtdcIcEap9FQTv6pWeOnqgWTsK
KUSzG/lz/z8UjrUmzlnB01s3cMMq8FtsxOiIWxPD7kSsFtR3VqZy1QyluZ97
rvMTIkSzCwvgqOoM/ivImaqpqGXLhmRHiyKBy4SB4go0/rv3DN2pQyd36FHl
tpRBlwAQy/lLQgQDhvOzLb+Kb6lipldK7WujkK3Z4fHncqr5ft4Nj1Rl3R/4
LeTBzJKGTC69xo6TS5sxzawfHIn0V8bvAyDbkycLOW2YFEYDqQTc60Ft4cxj
lrqSc5TFfVIlXVa4goB3hLzMmCJ1HkKQo1YxyJXVkTeA9xfCs2ESP6/OO5eZ
eZaC/tdu+f2d144T/B60uepWKtybjm/UQxy3W5nEyWnjcc2ZaHWxeWD0Xl7C
6yQgd0l6xHOTQIwav03hzBkgzvlQqU1pR8Q64zGd0eBTtEsmq7sZelB+dxc9
KWjGGc4nXHlY/QpmLK7qzk8C+uhVLj0yFIqj6w7yfxtdU6szu7ab2fluV1rw
OTYf/tIr+PQlqPIVKSiH7xM8VHLwFY2e1nUpbuokpjh2LrkSRgPxwYdmhLZ9
p6E5cB1NEdEuhKHDzIqlWiktRCFMNOWUq8NpMiS0+2aLJAck864vdlYcC5KY
FgYt4+HYvsZ7fKHCqyN4IilRkriP7MkfalVk9x3Xf1i9DNRBeIUPH2JfSo38
KDlVHMmo4KP7d5HR9P7ZZP4lwM9ULYMyBuXYrFgVt+x4ntU7EmdK/lFKHJ0u
PPt5jSDTzUtqpJ+HDpPLWgAf2d15XcEdFF6m8JGab2m0MtgaLRhD8EXcgiB4
7RG1BqxtPUwjWVxsNL8DvGsDhmTWu4HMStmk5aNCGOYB8dfNPL5mDhG6hQvz
g7BVw7uzOMj8HxhSveQ/ekDglrrUbvU1iyTTWNajyumZHecceVoblYkSHiiG
YjxvXyOatwonkAe18x/y6leSDfgmx11VaS3QZlG2b6EMx5vPBC8uyBdedHW/
H7SjwRgpD4xGvDjD1mWDjsS8ktGT8VwpeF4ucTXlOjRsoP776i2AKVye/HhE
vrnqBoOIWJAMgdfFqNn4jYGvIsZaKcf5zam1hyb8DLdYPE5NVtx6yZbgkcXn
VuvNlG351a5hJTL2zGgqnYJ97Z+EGcvfnr5GqCbm5l6/idwvQAHZ7+9BQTMe
9wUoN8YJidavOeA2PlNnL6Wmbr+pJ0hv8ZBITRIqvnzl9EYkJ6PdTQVwc39/
OvOS9jCjn/GiCDNyRAxQ9EA8wjnWz6CMp7UsZx1aj7aY4kCUcd2jLEmCsyLv
apJfb6MJ+o2o+uX3lTvxusWscUnaqrmpbEosw+2DUNmVaAeUK6rSsIfo4Dn7
CSRvsI3XedwETDGEQUfDT8gMABC3x4Xsk8eOI+iE5wSSqa3tspi7iCKwNZlO
0HWfCcin/qWyoQbSLhq8YYw/yJ8rHYddEgTYbiFKsDpQM+c54Sm+RMZb6qPD
80S/PVp+hdMk+w0Iv4IRRevvkIiNmy0Sj7bdTXAs9YeTekJqVDFGJ/6oTiiu
wnroa9ybhWmnSw5U35FQu7Cdqf1nvBZh0CRN0hwEipmo8Z8Y1a0ar5+QLjxK
1DbEJEaJ5rgB/i6nEJOHm5c1MYcgentHikajM1v1INclu6AN+vl4Eb9iQGrd
PAZE3qOQ6xMrFpDGZyp4YvFpFUiaGJnzZmcoOyrdXg5u0E7G+vBvq7vTY83f
+zTiPj45/7gs8Q1QtOv5XCZsUgVFnmYJIM893GkUXx3kCBGDmHp+rMswcG9d
hJn1CSYhWSSAu3vlsLGNcS0LJuGd1okGXoo15GRZLyVcK9vX3ucH604a1toE
6/EIX0qXyohpXcjOaOP7d289DJEXitWGhofarOIsJRbDeWX4rLMULFMYUT9T
rbcsaYwLEgKk3pwzV5h8baTrssIZ7kyYytWb4HgNkqQ9KpO7aVihdEtsRF25
l11o6Al4enkyUqopMMxWj9zob2OHmcHsfqVMJWM/7dbtpF76DWeOXI1GWHJb
77y0/8x53pLy9gHkPmio7/uOqsQoVFLE+zLkPET84z0dm6gWKr6dq2eVUr3S
8k86jEtw7LWbXg31oaI/2OPeVmk/u5rXLMMA35ysUShUD+40HZClnhwH1ZCn
PwXOBEyiw4YH848HpT7AXwvoXBT1OyVJEK1JdEaZTBPDWb2rlMV3fx6Udp/P
SIYFq47RjU2SLCH17xkSnqCsLmvndK0zZTSpK5jR4ET2LjU7uQcr105NgWNI
Dfk77clOvs3jj1NheA2/VbgEdCb8hPfi7UwWqzVu51e3IzQjgQMSsSOCHW9O
voerK08BdjKV6RShLMpiprmoTHiiv5bMecRIoM3QMSEU0z3L1X3qRuOKa6wR
vdcWTLgMvhAMyPob9Pe4yFrKdCumdolVNiBtsPYOO1D94iGIXJFI9sWsspqp
Gp+3yo1jne8GQXxVPJX5RtlHj2C25sw5+NvAHgGB7g8MYf88qrleocSBox7N
Q+Hy+C/+02C4DYWt3oAWaCp7SfEYhrXmwav0XiGFi+2MBypKf/TCSJqbFd6C
TMZQqMPyqZU7otTiyXwcztxwbA+NTmlp9ddiyJR5Ql/faO2y8HukcFsuuhbv
4n4PyvZhnaFJ5hEKUqb4OhNWnjRGyTrlIGkefgxETnPA+ADWfB51gxl+v8NC
aWcs/VFBR7YqWid9Uk2/DrEh1DZoH6/fNaJezYN5iwfUpHy7Z2ycAB68M5YY
KvePPP1ZSyOmiT41T48xmrGEFEwuaYqBTtUofgDCV+7bxDfGX2ImgFotz3Rt
EXFc8JKjIEmnwFhiGspxkbiKc7+8omYi5KMVkc88VZ+LuUxy3pfL5L4FLzDH
NYUFtghugeY4yleQGSSebteq5tN+wVlM1t1vdAHa6DwNZ58hMyWtwc73AWtH
aS4HkhYf2/IU7GHEQ6V4/sW27i9ioeYhw7lZryjYsfGO8zqAlko13ftfQbdY
aqWwJGGskPPJR6QSM8qi6sMdSuK6uKybAkAjX1DNoS/0WwNon0YHk/uyWC7l
PRotNJyFxGyfqVH/BkppigkOT7HWhop1Es1E/bc4j6DVA3rjFnJZgBGFt7Pe
z3X/vW1sX31IwjQSPjXzSu0ABXhY8IyT2j0FM7ukU8HhZfmwRsu2bPXBhCEi
y1tjHKepDp8K46mBOnugUcShxzGiwImk4TmoGp5WrHd9YLHBkm93twHZn3Mo
yqiJUKmZwW55TT3cqiQqT1i5Ya2gHeIjOYA+uMpHwVOcEaj3TT5VORRYlYxZ
IhMv3hPC21kqP2YxnfnCEclGrowzEp+wypGp7XP5aEtxBca4lu7V0zudBUlE
AGme21Lf5Xg5qCQT0TeAPh7WfiURaUqq8J/B/787H42zjdwqSXMsLbmToO1K
3wD3pM7BHLmFkfNI6b1bxTkO1HUwj0jPWL6EUZAzo1kcOrZTMfX4lgChEWzm
04Wuc4tdOU0eu4Cy6PM3nCnM9+riij64wII9uYPG+o6SF4FtTba8YQtf2p96
Ddi4wGJ/1u22dNtuqU0CRfLtKL6ED9XgCcS7n5k8vWRWDWZ0Wp4GKfV+WvNL
6DBWCRhdeYUmJRIF8MjfFmH9+sSBcR7Q04KGfCvGbssyCOtTeAhmssZlR+gx
E7E1zFkDqtDmiPzUetCzyxuE2gSoPuzdYQ5EFNtRkFGKrtRWvStjMW3tAeeC
tzwux2CR90VSWFlyDFMyKsTCz9XnGJJELRfQ8N01nuVeGeXQB1lA4mj9QmMC
3qxD37YpbO2qZ2Dk/OmKkjJP2I27x0PtEVsf/oVE6YFVVj3GvQJCzCydin7O
njcp7XtcJzc/LunlESzil1+p5lO9n9iQZ1LvUI9Mv39JBSQFzPOE5WGcpWUW
BKZptr6oRq21Pbcp0feXQ8dWnlvW1/GctyAHYfQ4AQz9WbCqcvtjAeYHUABR
gt6cNF/BpraSpARt74g/87A6Ee4MlPQWAqP/9+zfhLuDwd4nMz/o4N448twk
cCDPv4Wd99u+52EPyFfQLxbOA+lA0HgmYVD1SfOX5CEmDqbQg6pElrF80V5Q
PY3wrdqrJbxjpO++ur+BNLcEwGyGfLL2GHdVv7kSS35mw7ibDB+WUwCPn7TM
BJDDWhLY6u5jW0GEGXUGWYwRBrqr6twnOFG3NLwgCei8dsaG5nQHMjbv9n/k
E0c/Xkna9iEZSMiAjysO/iMgGaJsdiojvso8oYJwqrovLwxk4A0BJgdoWJni
meN33ZPVqZCVyABhb0H3W5PsCGnHzGOXrsN029Xt0VmyRgkCQC8+z3752c+W
azyafC+TtJD4kDLAhbyYh8jh+Y4L+JTdQ3BAtU5l5MXaJoNDXrK/I679+2n8
bFfxYuqCTJbz4C1dxJ7KLyHeIievoKctaVPsjXF5m/zKCmJJHG0UNOOdtqDT
bJ4da9aYnpASm6aBZ1YHoon1XhIM4R7cZUKWEUOYJBFhEAyMcl2L+AklKYth
d8tAqj5xyd1YtUaGv4eT2nwgK/nVIhO3Wj/h/epgbiQTnN4phpy/YVJZP7C2
yBunTjJsZDTtZ8vTzzfiFkJRG78RgSLXR/FMmkE7lqmknWo1bp3ATlXVHEeS
jRM3e6rbMss7+rYHKMF2LVNPRnpavmr9fsDoLnKA9a4v2GcyAsDJaykr86ZS
yc8FaTkfbELOU5vWu/TYPNtAHvy/VdWgOgayQC7vf7IF9Qi5PFvMDnBVSskq
LXtqXyuxJNn3m+9EhFJRo0o8HCLDEvvB3vc2z6sbmDTggLxeTjWkd4AHsPIL
a1Ggam+9N/xHu/6XJ4gsOeL942Zb+k6evRa/6s3hAl2lNhwBfc246eTQWZpP
ZVxz7GQUcHxtUYiCLDIZKfEln25ghDZTXOn22I2aJmzCO9PJpQHY4CSudGvg
VDyaUBn24ZTNj5aIbDcaWlYwsx17Uwoxk+BvguElNbJzFrdE4q8F0w0ZLbRF
hKLWD3qDIEmSUaVxlrpwQOspROE0a5Dj/5jVrmRJYpkntQseZKWAhai8Uaj5
KRAs7nKrdfuGOBTG9ArcLohSpGcpZXpFOVh2E8mLLEs8doIxDKJIKFv9JnG4
MGZLbCxgTwHAux48r7+QfXq1CpVzAUVUw4ru01HJMD92I2PVFK1JMTbZ0X5U
UWh7gPqie206VqaFoO+fbzNkyNw7NEgFN4f/A8Yi4SdzT+oQZ+QnEQJnlSt/
MHvIM1Sib0vaoSmuSP3xZ+NTXtM1FV0objLFJRifi7ABZJkSHqMwudZpZYTJ
YGvWzIoqW9stf/4AfwKtQ9dez0vf4nigdH3oyZf0AxmAbQnci+amuadWzgFx
VWPT/dho9fOzDUjmx9JDXvoQaK1B9XZwXtMYe89QlM1QGirRQtPLqU4xA/L5
vxiz4aBNJtaw7pJ2xjWOh9jjFZzSurYw4A1usouzBr+ZspNUMzHiXnlwdtFm
RBLa5MDnxI1fhwHnG8UkmgbbUSAA1Jef/C6ioAbis9RlmOzc9hl0jUUFHSK6
X+6fXGTUI1iDRoemOMy15E5IHrQW3DkwDtLZGhBCpGneh2BPa2OoCdfgCk4l
W/1JZyTd3pWS2p1ekfnMu+/kLTNJ6d+0tfj1H2sG7wbOr6VEhQoXOE6CXRzm
gzQ3yACV/uslqn4+OgfPpi1JjRzS5RRHNOP9N/m5A/r9G373jCXcEsUPGnEn
CQRpcVPGUfJE+88bu2YUHzvlhv5InZF/bliG2EWzlvjMwwCXkGHDHy65MG3R
mQUeqtfojlWYGOWq413JHHBkeP6XxVvOy2TpnBmUrXEj9aV1/l1VemWVsYj8
YgTtdQjJ5JdolySAwPhJPFQ5OOvafi38bWY2ASMyFTjdONozWyFEQkG51yDn
UVI7lMdfrKuykM3dczD4jxyE/hG5EOKpSPP1LWSgjKC+J82/xbj9cmjK5zT7
91EBIlUXu+ZQAA+SHo8dHFYkBzASDaHhR0V69uHuiKVTICv6DjAGwtOLaAeL
sqwu15xFtyDmEj7xZc1yatMoVlTGKfFhgLzXh0fFyZnHo7jJf6fVxiVgSXsa
KOCj/URftoZajyIG63aqXFBgS2EtSNhlkvJVNVlfHgToCgD6WDmRcK765aiI
BKtLgYopGnbN5z4/HiQbCGwcTfDqtuFJntf7tbZDxxNJr2TXw86/MKxmaHXB
ZYnV4AKxe3wddJeYlXdEUYa3nALaqab+JQgtgh69KBS1ndouAlDppxrYx7Ae
YHej9h632xWnE4IUFoP0csnXT+SifCOOlSUtuekakgT7393aNAT3jbZUqNUz
FvZ/7MiIsJ3lgmE5Ram/5KOYs7eE3Mi/sByocbwC2fUlNb+qlIhWZ1WYNsTa
DDB2e8PmWGwjdN8M8VE1Qvc1e8eUvkjNATavDZnXlputdtnypPpNzgC+/ria
Us80f/ZQJdTbDejV2GNwuJaAg2aiNi1zliTLI3Jio68RgU2XITEnFeWi29qr
Hl1Yp1I2k8gc7sUJZk61XhDzglIEkeb0KDX21Qa9sZmMw96vkRCTT0QDYeZt
D1D0GbO44tLQY7KEM3v1IPzCTFEB9kLg0EnCxQ5zTHHZVzYL8z/TgwedpXUV
AEw4KJ2+91se/N7CsRArTgTPm/lqpW0SzphodICw1gtXXCZl+Nzk6eSrhq18
uuwPga0HNKPiUO80Vq9VmcroV6+e0EH3xC1fD7p2y1uyeoEsmKHKCQonFK67
HRuuWcA4yq5Zw4YSWrDmlpTW82usPCEy9FP7uZ1G1wniyEJ6r79F1XrLjZHa
juq78J74DPd3AyXpkAC6flLtR1IfuvDYrghZo9EeUgjh2Oxg0zn20uUMhGtM
JrIsuxWIBYofHaxlNa3MFX3U52vd3SKKz6ei/kis5JBsJAmVwd5yL5Lr1IOx
AGZTcVdPevGdtibXDPty8Q/nxW+ZAiiT0tKQtEkDNSfOsfpDAApbD1CYpRn7
I9uB7CcFGcSEtciVGbeG9D3/q2dpgncCVQQxsX4+3hCtIKDEzUK8yMlhKk4/
FcLnKyLW+ABHia6rShYwMt6oY7n4dLFv+aAL0g7i0ML5vxU84foYAC+EZtTW
4YBO0BiDFseHjOdB77BFxFIB2smM0vyHNcB+lxlv+XwI+RZh0IZRxnM6d/Zf
rJewTvU1dnlgR30qg9SwDXwwOvRMCfcqlXMlQQGff7GcnWBWPegxDqWdMZ+5
hrf0BYc724aGqI/3O92SV9K5WH4wHcTHh1Rd+1YFjkiruY6PduPipYsWkQ/O
gcs4MeI64c8nJkTQccZPB3HFAMskyNYzVh7o0fCG1kOGV3PwJzmrq9QGPK/+
iZp8pct+EJcMCycvTJgbadWpnsEsM5+7Oztv3rpAnv9Yimufg7q6dZ67AZm2
WZt1HnMOf1joMDyaCXubRZaPMtgXDQp7N9pNt4UlALxkVjQTXa4SueM8NNfQ
p551xBq5uQt2USO283l4oHIznlHxWWAXQud5YBfEZSA2y4i9KVqid9p7yOtd
Lg9GCQvI2+sAVzdMqDz/RqWeoQaqr7yKaJq5fLIKk/BoK5fFAFX0vhk6VT1P
0CKi6tJNo5MUdvhr1dhl/7n3uHGqHaXHEqLRToGjwtiA7g7JJvl+nQmf72fY
2EEjKV31wyiJ7jtoSvC2tK2dqnnQej12UB+wVginRWp0zH5b7NdK4lPjIcSm
GLjsNofOBSz9+N65KG8wHLbyBEihhhWBiE6pvVSboA4QVFNCDOATztP+C9Bd
XehCb1LevVnePsYLPIVrRzMsepTJcw3UspW1pffMhyXcpghUnR3lDVMQSrcf
1An/q5+aY+McF0xGIhH68VgBoe7EtnhiHk+N0cfq0hI3YyC2NVQanbjtievz
S9zVuyFVkMIkR9EQwnrA26B13Pl0SZ4uE4qQkHX4whccybQbT2RlTXuGcPJc
/LFCSWTLFAAtz5lZsCQBirGi+Gzrxfmf9hasIaHHfLGNWO+RjVDPsfa4R1+l
l89Rugi1AIDWIfUUjFFYuYa446KdxfK4ZTZ0JUyLdbxrXWS7YNmAip2MhKyZ
Pp/tsRKDMP5MBIvAU/U/cJS/Mq/CgJtzl5qNjZcVXq7jBV07AUaVxQxFMxZ+
0bfwt2leCPpvH+nCT5zRWmY5N8Nyxi5kn+5P6SSJiTUKsgVKW4vQowCSwBby
RmK+wnnnvPQ/oTsHm+BmQybAj+XUOy7Mmd5PB0yMs51CE+AXyQAMtjnZZQcN
45N7CGGGga/c+hUnPwUqv8o5j7TRcD7P2iy5rW+VM7tpzHumKxgRRISnUa8S
UhiTBP/2KvnGx/9uQKETAS8KMr2WWFNMCBOg6A7yr2x2o7W5AcuYI4TS4aZY
ekIwlrneVIbeN5YVO9SyrbGrMKX3XrI86/60iEy9NpAjTcnhLtrPw5YUpyT9
w71Z2dA7L17belgqZPeNw3cW7T49VMlFCUMyWtzfU5Lc7RN9Ws1qy8dK5/9/
VRwDEwWzRNKt4BXckKn1mhjPHiEp+s8czlP8JT3ef2BAyF9V4BhUnnA5UmAh
jXUPI6M3p6fy99vta9usNxHM7TZ+DtcHiDMC2bWoq3RGnDD+jqL6/Cflqdxd
6UyWR60J0g5iJZUOfpZ06ji/sYjFsK0xglDK1LZK+mK+5cvKxx9ItaHlnjKR
iZytueee+pnRSyFHZLdh2CAIxeEL7Iv+30Rti5j/WEs/evre234inp7RFYLZ
2gbtUw00iQ/KPGc/6lWFCPsrJml/OIUp/sfZhqJ81gmo6r5i0Agzuyl76hhI
U6QxQFym6Mk1ROkvcyzKv/LjSItXPj8+gS6w15JxZtEZ39WLc/5WcYxJfqG0
El6fMEUtlZL5zLBuIk5HaY7Ky8LkMyTg2G1kVPWfpNmfx1GIlWXI5fA7b011
ISwSaoCdzuHrADqgZxKD1z0RtX8I2i/WahjnD5rKGrhRcfKH4a2F7X6LYksU
jZ9aqF1cfwaVbc8iTLw4o8pHrRFC1KJPubdFSA89HY7g2QU1hfik/DpI08cK
TMIze/6FdYkUiKcOL2YHKkX03hvVcj48I5VBxpcmfEM+ccrT/PE35W++bYpn
kx8Zrh2wgyi+Rp2RUBfz4gW/tz7B7Zlvdg227jhZORAI0eKZ3hyoiy7XIevs
5tCZhgcvy9Uw62l+rhTHO7HbZd6G4d3qczch5QKKZ+IdxoiiAX13jA72hQb7
sTV9LSD5CzTdnZQiCVxTQhvN6BKBobzf19dCNmGY0N9dEvat6ULqYcOTSxms
S2RKFUai6oyn8P+4M+jbJIZ3l9DtAZLDNsfWS9MK57FEikn05rPg94SkeTfa
rAHTOK3qvu17M+ywqFjocaMWIXULRYY4msAsQMJivAL/T5K00FQWk/8QOeei
uq4DALDXC9uP6rtbT3CDSUjTCvYkCbWRs7nDAr4pSePttS0kVVwcsVkxIP6H
zItRR64H4VK9Tas7s57VCas1rCB6M0tKoI49StxGRSlXqBesTPF3CAN5qrPq
j2Po49TA07+yepibdaf74Ln96ya+hD9e++sbN+G+Pf+kwGFHmDpxqSzp5TZm
v769h3YS5qp6H97vPBNUUAwG0SPRzGKmpIvIMtDLQyEqYqUPR8KC0ZzBSKeu
ovGKSZ1tBdYwq87d4mLN7l7krXfKjn4gfgca+uYqm5YI7vZvfpfeN0bbBM+H
ImOvKnBxTZ0gc1w1E4T1BP9X4R7C51T1nk9IBuyN5hL/+s9a7fEtG7AVI2Jx
56L+eyU4zsYtkRprtq/+oNiH3j5NEhog3UWWkVIQO0dJsSRFxNqsFXtq6lGI
dhhWrNxXPeWsl59KuHZdZk7ZhmD8KBKibnGE3dgxcIs6QKbF35UXhdKPU+iy
GYDSUdzYMYV7Ta7u1C+HJJ9DAAqtgbqq7oJ3stb2qgzx8Lr1WnDq/IC1zrvG
6I9VvnqGIGzDEf88cVEyUwYsA55LSkMhjym/qNRlKtOczAorjrFl8cgGaOwW
JE4/LUtheSfhEXqOQNIfo7q41TrGzw93CPm2vEl5UVI9/ajnc67e0FbMzZZu
F/ILS2hB/jzBuuUCdRy+P1vUnCECQSGY3TOsRXhkTWqlOnDnNw+8pJ3NBUxV
5Lf9bT7HtMlymLvJJdb46zDOjM79wyZHRX6bDt4K7t7WPSKsMn2NQDwUiqAv
ERMYLU8K0+W+sH8+ZhFzhbPlGtLsJ+83nbdbGTO/1m+taqVEzuM/jwhv3egQ
NLwPak6myjsi8BFrG+RM+N47XUwNk42HBG5Sy4OHIfxF27kvtgdufN2Y4nre
hk5fHGiK4WBFJ1UfEE23OqMFG1Iz1HJzpK6QvQROgaJaljPlTEQ4u8rEFpZJ
fc7PhntiGs1sW+I/uI32IV2cAG7/yFbZnHM9HpNEY+/9EByaC4fqdhev75iy
sSKlB7wRM7Je1Lic3vFVgqWuanuvAQglg3xQztnix+ZIvCfokwNFHOgpMsBT
pW6dVmbsdIIY+Di4QoB9tMkZs4IdoOEc3Z6f6Rw19wEulSkTHLM3HorwjQVW
rGM4zH8w364O3KSsRsHzl6TaABxAifeICX/rZLkcbSwRvg+AkG1N8CGO7QiN
WQ2uMkCNRST/3FccLWznsdAxIJ1buVkb1MKR48Z1WuKnBikNWnKEIAzdbqNP
IJPZsZr2fueX6gMlmVKbWwQ8ZzGNR5jRof/PkbQuPYvEqC3Y3510isCEw/5h
3zccZ3RKk0jww9qtCJNqFtCAPLLmH9hHBQC15wIvd0UpycjgAr3JGzwM8I6f
gSQhmlvrVMB5hCTpwjCx9oE6Rnv4Ltl2ockZ5BpkTmH+CBp4brTUl75Vhfzl
8iqshAqt9CfNDHDnu6xW5qqaGEXbkYRPCBUftrB9NZvqcJf8zmOSRIH02G80
a9px7Jaxn0uiushEH4IWcCKJbC+yD0PM85s96iKhag7AUBhGCiembZzKumZi
8DwrRoTQU/h2HPPWUH+IuRwz+/T16ycZ1KPi4EtBmSDBeGSvoKFXrR6unnH2
1PP2iRzcWbQMNz3RTOgM4RNeKsbF8nmK2OCMv/175Byi8TdyrAh9OFhFyol/
aVqqUcOcnPfWITksMjxLKcVI7I0r7x7L4HHp7nWPPEvtFNDrwruIb+TiDce4
flWiyH6ThcFP573TxOJW+XqJxo3lAJB5XBefpJ0VzE1cL1TFlLp97EVC9H5/
M/r93Vpn0FvtbHXMN44C18aGWWunCePavOA8JCiQMvrAV/ER6sgLvfF2jDat
pH/F8qY5CVqVy4jNFz6hyzHrbME9q5XwwLarbvD3vvGRgDSV+p3sIpJDVVlX
Yg1RM4NOuSeUPkIQP/ijJWgo4CpyJ589BXGDE+rhx3dsHyZXHK26OJsESnt7
JGzanhUrjEJmirjgEg+Z4ZXs2sMtR17cBIFXz4KXVfDUEbRXrTwlLAatNPf8
6DxgPNGEN2+/42pcQE1f7EHuhopq4AqZGqXRJSfK2mEUjvGIwmOxZLf879Q4
pjcdiLkJkvpRHvceaZFIkxlRRo3oZoTu+z95wzmutuu2pdeBl3/6oTOfOHZw
LTeALgyYou1aVGKNepqd+taTL8UZUO39HipXI6m1zidpXtmRwV8jvexbcPvj
2utPPmYKfzMB5Sa8RpinmHpU4dpw5hu0ZTEBGE05fzuNsS0ax4Kkz7vyKkWs
x+Nfynls1+6sivrOpdfgfdaEFPpPcS6sxCkSCRRs4YcsZb7MkGBY2ELIZLE1
2PtE9X5kdZ/M8ms6wS/oeK8/p5Mz/YTl2YWh5RE1FH9Ee1bp/zgM6JbdyeT0
HC5xe8hrllkoPQJO6WF5JhNIwsMopZEsVX7WxSac+WdX4tTePTxFc7lJb8Q2
qgdWbsz6V6iRbVwbrtFCtro9RXtxOHavfvsZZkpOQr1IJzeNm/F0mjJMgXo5
HtLaszyMSc4Mexw8PhrVGfRXVcZDx/1RHLHFx5Ck6GTi6etJWiNNbJ2UnTlV
5maYcEJyvxy25b9VOYpzYJCCCTxSORpXLzRU4QSz1EfdTq/tF/YNEbBizQFE
qKDMelxUZ8icqB+kbaP9RPBlCQ5jjtfVXwJcIWyMnUhJx59pIlvw+4+h9pbz
9W7aOlAHQvlGBRGHgg44W2MnsXtLKuJvTEPh6eM7hRS33BJgYNUbhJUM38dn
B/flaYucIGe6NeTjHtdtM6sfVOYHqQ1SiqfkWo1QoyNF0vUFCxG0t6IQZPwp
uFHMymFl5EVJrA2lnAtfbIs4mDh/k1xzIitNPW/oQ6nJv8OvtGYauXW1MTHY
RzelHD3NakOYopq1sgGac2rB0qdJAuUMhf9y2FzYFGhRxmFzn79+VfLTZAIl
qi7xMTIYtO8L1C8OV+RX770ByDLqDS27hfWR47KztFwSLw7QfD+gxh45V70L
fIkPL9tNz8DtGhOj2hMLZ6X4VzAvT8GfXL+Cpk9UWUNZ+Z51D1lnyj1Cl9+A
zysgROvggkJuzETNgSnawyKE+gkPSR/aMKt8h2ubxpZm4ERSoYfySb4l5NER
kZsFpreMSO1mluGz+hyBj+ZhM/aCo2Hem8gVfBWxb5Fwn18n+ce2wBUb/+Xt
Oj4GSC4KTc2fS3ZkPfZRUo7otxourc1VjB84WKwE7q2svrDUcIOaNmsU71ef
QaOCB6mCeKXHnI1tABvJOhrPHnDRAfVhBD+VuENvZHXbHDpUnCOR6F3Q6Upl
uBFXrmM5gQJbJDa/JoEgubwG9MV6pg3ZrtYXcU7gkpwO4N/8cGRavys5lT2x
CWfH4vFIB2KCiMWNch/wfb7b5U1s1ac/UPb3/bFoDILywnvMk+hgwdSG0hmL
E05i8e8vJxecnDslCZupDePhU2yNOwigxYTk87xHHfB+1so9b+mGtN5RXm+y
JE73FCwDnYqny569iPqY3S+GurgW8VXsmD6Wzo0Lt6Su93LDlRlPMhUd/TN/
3Z9Eq10bU7dHzXvhdOsttCpcBzxJWXh9xE/NJXdId2YHBV2iezd2Kvb1oxgt
mIjj20ZRfvhsYh430X9L3q/N2sz0r7m5fzOFysbd3xUawgu/mXIYsRCGNjSf
qUrjGKRvtpCchyFz3v9P7CLfvFpCWgZHDBuaY00Ell5dmfvYi+IuCch1p7jf
Ee/nM9B2RXP0w5VgCOUN4a7MwrTxEH2kD+5D43zKkY+rqTvZdw+BhLNH6MHa
Y+r76BEW2SIdeZYesHSxDDVNnW0lShNtaD30skiFTM5uy9hux9mmPpFdo+Nj
X+RdXs+WX37QdVxkpMzXkfNEcxRDZnUseGk2nSHu1l9QcK7kiID2RN2SDWJa
kjUdz2hz1HJdKFwHg9+GovE5SILIlK237EriuAvhGpnjGySAMlvHOkuJL7kf
TB0Q9msA2A546NLpcwdR7MjRKlmf0csRyG2SfxcW8daWV3Qd73UdK1DmKypN
2AIMILSIB6Y/ZkP41Vq/9YOTbUai9UKVFygBtRW52+GgdP/59C/3Jixy3O5X
31aI+ptUnT6ffxVtsySmyjblhVOvHkaQspKf/I+8ZpGu9LYaVDPvwEPSZpe3
v9b2TEtmyi0e8WClKWMGGFyEWQt8ymzMQwBi/HdJfEhY+IS/W/jTdgyo5CuI
ghlCtajH4ufqzkg4SiQT+p7EkD9yyZzjgOSHOCU1MFBZQyS4pV3jZCbO7Htn
WULu2DxZ9i0l7S+4ZcTUaP0Qq2KoPzZE0LRrcmmmqzwq8ruWM/pN0MLKYwdK
rS8PQiQvOWhrW+Yz0st3E0tkKBgvFVg+PdgvGRzFJs08w/mdhRca1/pgYpA+
5jzQa3v/GTh/XyYbbAiDwtJOaKNhxvczblSu+UEvvZOr/JfvE0eZgKO22cde
i74px8AqNB0PS/WgZx6VvRru+E9Hu5DuqZlOSWze4QQJvWYa1T72+fYnHyZB
AFRkEg8fbZ69x7nXTpeWZy8HQlMpjjCn8aEwShmcp4NlvNYF+8hSBxC5uXHZ
wAmOavQc3Sl6oSSHtAw+yapMtZL5erdwU6RdKToSJ12zqjW2kA26J30dBetL
2RwxXTxbVZsuwd5k85qOIWIg9lVI+uXweaOviYWq1IAAXaD0H6T19qNhkkxs
RkOR0PM7AV9a0AhBjZ/9kKkuryxIFiqnJCTlH2sUrmxk9WzVIb4z2OGj04EC
BgsrHgArqnMdkkYjWaC7BEFENuIKRaLnTyaxDHMxbUqQwhB249UKyvedck9t
HVmYD928ppq6n9/sOuz9yRhei4BIUlqbjBs8ggaDRB8ARtk24HwToyJKLJx+
NFnZ6Tjx7WmST0jQ/CcfVwWcFZU/Beo5bggp1ko6MOFHJAwP+cNugOmHHcIu
u7oEEdckkyT6MYVr8wLcFtzU70dg0B4ONF8EZbd7E6jVxqz7gKCCwNIE06nb
NP+40JPwf2PA/5cZ/lCKvC+LIQFX2jYt6kG/SApn5C8sj+ZULanRcSv9YFh2
SeBFDsGUVt0QHh86AXeqxxkc75nAaFJ0jgNgK9JfbQbWSsmk4OMr7SVf3H/d
JqLwCKhKUXZaP2nces1OTtStcUbKXJKe9f4aTxUcgbo++pHq+mSDrcjp4mtz
biMCcJoH2/lpJfH1aElilpVHIggQyf8ZQlNJmKvmfo7fuN6HAtOvASxBofZY
mJkjRnLIDWRyV3iFNbfDifO9i8Jqssm12oFXWXOmLhwMo2UwWBcGwqQMB5Z4
GI7tXhUEqEgP2M8X+2DhmBufU2IJXbyrQTRxAaxCKnNlGp2PWXluGiFupDst
ZMtMj8fFYaxY4SWpn7w0bTSBwRf4vcrEtBfgJHk4Dco84YkKrIlUN6tgjdqu
mMVbu3ZpX3TImDcDjpFZA+nwzbALwbrv5kFaf2YWCpLcHTIqE90oMVqLjJ1Y
8Swb3f4w09BSrYtKqZmWFeFD7y3sNnQpwpD3bEJN4ytD3QPMGxWcvlR+AKdd
IcuPI53pSTjDeWW+qS09AXZYVbnPV2Bfp7U5+/XeGuq2Nh2St5DkU6/UHUEV
Xh8IkYnHPLMxjVhxHyveFLEhbSG9lDl9xYpxB16UikE7DTvh2QKccZrdfK5u
YdhbxcumCvdug4kXK0NJNNWhQUVpNo9EsqOt9i31aW4j7XbG0TpSJQ9Ot5Qu
2DOcFxvDVmszNVVdVxsEovE99LCQHEGVkf2a8Mj2g+JirzdmUCcksciSrCs4
fs4FZd0on6dbMDa2kzHZkbGZceDitGrVY1YEHYewa2lSXY9TmCS1BZt44Z6H
pKIuN1gawci67ExB7EDUkaKdzlOutwHR+SFf1+WNonNBF+7j6uiOwcvKIiRT
RVvttLHdmeOuSPgLcvJYLbqjWKFt6dP//hLYCQTzRFGwjXruD3jepzcdaPeF
ysBVjzaelF7D+RE3sE9iTRJevRjw0lwmjnRTqknQLRg0UAqtIXMca32cBMXf
44jDERYPMPsjTa68UVT1yXWOAadi0g2KRREuklRBl6kzo94r+Hxbr4X05b5g
Anz1PDtIJeiRuKSSi7Mr9WLDwcQFjo0s4u5FwooMsehdPqN02ozrqBj/CsS0
xjVwmrjXYyDdd1m45jhBzDSRl9BFIUUd6RORVyKqcdqCU8aCu4XGtQkXNFrP
iewKlElt76Z8KLFc7+CKzpGyleqyYOqTzkFpPT2sBrJlB1h1KzyJNAVlq5Fd
oGHBqkRP61bAXL2a0vr545gNAlXW9MCKb7cYJli2IFqxoMfGhA7uzzdA6kYg
9eYgDr6DCoxpBJVuNzfVCbsj0i7YbpobFAQRP/v7Ve7GAtxtqrUycj+gtg25
EobEhX70CLlbWevCHaevLtSXta13c25mcTRRp2azA5WFIJZwGMMoXp6w5IEj
VDjugqfN1o/22+ux4HnRUgTueiZmBb5IILp25rL4KIE8YaQ6+PH1FLiTfqzA
WLEYqeUKrlsR4XTmnCzFbkkXo1CSZj6ynqUi5iLNPuqFO669lbLCnnyZCn/z
eh3YVPNSO5tSgm4z14ZpXjxYX/YgJ//RD28kCjK+mMwmfGUCwxx2oPrZaPsr
OZEXw9a+ZYgj4H5pYzDbwJk/YX2ulMCrul8pgGWPXQY727GyNzBh2uhbaliv
D04fbWMez2WdCOMFmSdotimoytgmkiuz0HwcvmLBSOsXUuG8/D0SmPEX2RHF
eSplDmWPLdg+15aBHdMkfx54nP190Ukjmq8gSnu2BhLnHy0iwK1eU1DI9RdO
Cytv+vZDCDHbIRfVaOy+UXBKVFspWCJM6ddWyxj02hXRYkMPOfVQt0r3aTxl
vsOLOG7HytJCn7wjZNqQWP8yuj0JhBD7FqRo0FJGQNPapnJxRGjSCCEzr11t
Q96Hx+xPXOo5i0cTQwodCml9WtFfJHqTEf4wOpBZI72Z4+15A9Ua4HhzRIc6
xw8jrUPwwP802/9DMUBv+7rZTErw2CAWxtfdOobzLueL0VQaY/t+DbWPDp+y
0Tp+xl16pFYgzR9IBELm9V6CGcVfC8+QsZCoBnYb6t3R3M/GWnHuUWLmRLWw
qVfANdR+ExFCewcbJEcSYOl0cvUpbkrHQMHNwSNVNH4LP5SXi9axtDDUaVdq
9eTUd/fjniNxasMF/0aeNjQ3OOVRWD6VCpxXTE03LYKV61U8kIJU0c928EWY
HA5zDsR/9S675PjJc0lFHrKcvhVdEHX/zgGmi+1+aJWISwl7PK92hhE0SBoN
yS+yJiAXth90OyclC2bP1R4q+63RejZ3O/4z0mJOQTg5zMTQRraHzqKK5NbH
d7R80Xn/ZAufPmiJtgM6xyAUUkiKjRM8lnEgBhKj6t/mW21p34/WUpP5WT40
fYEqAjJbbm+CBNRSxUKc/APMRwngHcpU2AesTTTYpCFDdziY0395bw60gJUA
wn8DpVOc0V/aPoQptzJZhbMBnQndsRvswgDebdX3mF1jxmeG97Ez/gGEzSbG
dExjcXrR5K05n0XqQDjyffW6+CSP+fcaaJR+ZoQcB1DYJlKR3XYKI+DCL1Bx
lLEc1t6E9NXq84jSyInEXAIvN0vDwrisXkg451MUeZ580Q9F3tcnJEQyM8Xt
JZlPt2PYSPvmKjFlpLbCU1ku1URSTYfue7uIIO3UXxo53G76+mM51YlbGa6r
ge20YavwS/Q6HcHsu35393mls0zT4pI4Lns4uO55sUv9cvVjQkJd1a59bh4l
6GgLDEwVut8wPDW7qfSYViwBQ/3WuaV3fYCl7jwMTISmTPpjSHkd+xBWpsa6
8mIzt+D0IWZ4OYn7OO//ZWQtTovzG00UVyEzBcmWYiX0og4Ghgyj0jvu0R3C
6bv4GpEBdraBUukKM9NFTvBuiU+s1nzlwy2dIjtn/B+bR5sPNJxZaFxsD7d0
ya7kZfDj3hGw7sTB/7m1rgRO5Rg4Q8JRzG9PMKDGD2Y8A4Xa78pxG1HYLjhE
aALYXQHU9tM7QvxAYbwQPB2eO5n+hC/XU92CZuu5/vHJCLx3CgPOEas8VXRt
bQ0ajk64nUDSCCG2TOTuLSHLDRrOEpE3cJx6kxOdX3GPMErmC1/5Ywsoy/av
cvKX7QOaPoFEF9zPyOSi5qWjuuiSB3GuzQg7s9ADt1zCrulIa9eMcL2nA7XC
RzqaH5KQ3s1UMjjmJ9HkeDXjn0vjjIi5rS+EvoGhWjBPMgZM22bgM8YE0cpE
nzfYOx7iZiTRoPoRSbIHh0IzXEfGRXv6hsGqOMwQOr27rTWR0ZHVSVoqTmlS
FA1YayoVBdNDPhPHRU3mK+g2nd0BVkbJE8VSdG7/GOre89NcRmaAXOMgRmtM
fOsiIMBRWs3iGob5O/jvpTgQ1A+mj1O4bncFZd3Vmay1/Dbea3fVeU4/FdZf
Bwl0NKl/fDSCiOkvB8DLh5ufPH8AIhuL3BG8cOnMGU4iuBDRugSYy081rhJp
o5XZ9lCoof4eDX4gAU/CUzwyT4qShHddkhfNTc1j0bqpW5zgXsAzihwtD6ZW
odcf05QZytJv8BUVTRT2D0uupW+hEWm09gAi7RAj2vewQ+YMHS1l7eKI+GYx
Wht7sL2tc7Dj0OxA9UsHHA0v9l0aI0SHnN3cI+z57b6SvVhonbOCTHNK4DBM
EHC0ebVMtSdzqSYjKlQAXUeEuIWyfBxSigHYE/xsBACtG9d7cIWIrCIbLKEQ
8R2Z5j1R/UaPxiq4r43PwfrLh6xGy4CU5CQttTnLF+JztzuxRTxj0Df++A30
x3Ji9IrSCtJ7RuyBO06J7zTo/2/zPQj3d762nibbmBFVIrRoVWgYJWb7HVgr
25DpvjFMzLWjzF5JFaPZBO2BOJu5xas4sSvwgJZjko9SCsT/1g2fjKHxdJQv
Kuj/gXIa/rj182gHvrMYzmReuzWKBd1d3roi9gQyOkisj54Jba9QYEcAFHyg
ei1T5Vg0MMsv6gxqajSzKYM/tpJqKpjTl1kiaUcMBenEXUGYhGcZJG6VlG7+
8Jyd3oMJdfLZM3ViONQqaD7nu0r9VRFrzMOZW74l2goHUk3Pf66ZrLOQfVFK
Nq1bKs/IJnwY32lgeo0W5Ul4xLOzemHzP/EA/L7dsPr/0SeQmVXgN7UbcdvN
XSu11LD2PLgA7Y5EqxjSL4E6RI86Bcj/Y3lxHm6TQ0zyemgdOXUBCTNGaB7V
ne4uZyL3UZgPw5+Nnp76tlrTkJe2Eb90j0YUZjP1xvo/JTdwz3CWfZmSwHEb
SGry6qhLvKDw8sjfioql8QOdIIpaEZKvKjyOUzpPvCyp1jJLThcQ+GQQ60ed
NxF20qsidBqp+VcOXxrjHZ4rjN4SI84I+wCnb8Q15YLu8oSrxdwHo3o5qyK+
zP4HZiFu3+gO7Q+vkwDQMVbpWWpHRA48uY8L4bPWmX9ODt0wBfwslWO/4aPE
592okE3RBruBEwbKIffOdJX98MKVIQ/QGv5h4zXywvrwd6DctFbtW7tOT950
VEKu/MQvhugoULACHUDOq+S/TPoVIZLZvMqRTVPxOgeLDo8uIlVL7Ue28cLw
kAd1MR2ZNFmr4wdPLVIYMycspzsdACDDikMFV1WiJ3AWO5NDVo5KzNUjtzDC
7py0KAYJWrYB6afKSIdueZQPXgnvFI+R3q1DGna+ASrGZ3wymMo76AF0TRO2
qeG6DySLYtigSvTVlRUm1FSWLDupo4WKqszwtyeBz2ms14noRwv4pd57SvJ7
1CQ//a1Hgg1yiTFTlR9fhFIVvfx6CRiTgdMaj0M7ldDB+7CtbLHU4vSbnsQH
+fmhTwlQSyxbTRHlxpi7jRlm3EG4v+I4eIJXf/fcNtG5osuEyrUv2511s4mv
EuYINwEg9cGY+K0VU2ffPvK1gUnSvy344YWgirGV01jSIioDaV4htxqwtov7
0ja31TIpVanzvAy+kGW8KxLpaU3VKGq6cc/SyTFJD1DBm799gSX6ZJfF2Yyc
Z57UfgVW0JejReFJd0UHgfv+XECde1YMIUDAkN4j1kyC2ERB0qIXEe8gg+ml
x2AGP2FlBnA5Uzfxz/ffgAlGR7sQSi3UNhLj4VXnoNcBKYhuZSvRy+45590v
caEiTa36jeoJPs7DLXsRiIne+aTszEAW4v0+E17IHKAXpDIAnpBV3TbNYgc4
cIjGaQf/5kpH4o+uCsjNx0N5fqM0nLaGmxl2EVxLS0yns8SQpLji7dtxxgt6
tvJf3FIcoZBMAI+rVRDyBhwypccNMv8UOodqW0FL4drrfLCVMhN7EU9y2cYF
5bvvRSoEYKUqaOWsXt2zNvmFgATQ3iCSUYuN5ug5RLgpUVZmXeJc4tzhw86F
VNzd6vwhDgVe/sSQOx4exlyBXZuaqym0wu55lVBFg5FSuE5jpM9yUbw8VApj
6ZD59EVQMPk2naGeK7+W6YVlr+MmE7sXhZyQbQzS2AqJHy2+R3MAfHBxOWiL
VB1HqvVn1Il4eqjLPR0KSHXROljjgzMmRM3eTrOr/zYREgXn7FqYx+BaPhAS
y7wlHBLPZR4YIRoR0mzmO/HRUDW0e9sQVaWTzryU9DBuJMrgNK1PFehjOGXB
FuNXb8M1OyKYtgIq0oAvdme1QMcsuX4WPl8rI3nl82DnKZL/PRXJi+pMM+pX
OgOf9ZuE+niRSpZ9vSgUKMEQI/Cf/uuEhnrKr5dojAfMZLqkFcCJq2gegMSc
lvYpNStrW5rbsxoJ40mpiC5jd871/DI9MUrejhhfaEir1m8tpuJediT6q4wI
tcEE+wuIlmogcGX5NR6q+zHj9AOXzXmV4wgyCKT9EBamnZAWJw4WcnNIQ89w
h4P6kygwQAIvsm2xdIWQFJmEOqqQjI8aYZBlyghWVz1QxKO9WI8+VIHIpe8p
SfpRCyEVahwVUFCazRuykIlj4eLVY4edq5pwInCIx8vfQYGxYslHT/U62KqG
KC/sAusBkKNjdXYDx4mimq5e5zdW2PQyKWX55SQyxGen131Rla7vS4tNh8YH
Zih+uFs/7SlF01CbCgQ11d88H01ajdA5WRpXQp4PqW8g8QWTfgDfnu+4987g
foM3BQ/geWls+CC1djKdLJkiPhiU6Zyh+zb1P1yPl6vULJTnd5P1PkVnRctb
tMRQ4sztisBg1TdlzIp7XSRyWJFKA/bESMefOBgWqGOZZAYFwM2rDikGqxuX
gNW1gGG0oOefpWI8zOccaFekr0xZD98AGoncj4Dq6Ri7M9MXga6HAd9iuf6b
iH8BcYPqq7LTopyAliBOj3EWzsbAliT+U6iYUb0jOsjcF/KYKhBVEXuguBM0
CRIdxLNYW6S4k2hOjBmZqRhowI5sFcj3wH26+tB1VTKaStY7fHV+YYUsaHQN
b2ZZFmq8WLfYNW1U/xruUNvg6XaM5H2jyBX3jj2BXP5aNURToD3Mc8SvgQCs
kCPpa0yQ07t1UzpC1rsNOHk5TJOsy715xPqvhIFtQkB0d+sTySsXKyXUaMId
nAVH/OuwGgrIkCWkF7m47dwQWqoDiEQFMM7ITOYG0QrbvfI+wuMsHFqZyl7T
UjzwCwUyhcuM2leaRR90GQYZm/eZ3kP9yQf327JDiEOQR8T2xFEcaK98d+8M
eT8LRuUy3IixVWvlzCP+bQ8wROxUqZEz8rQ6LKMnVnSqmwrH8I3H+sTydgke
nE9L4pfchNs/8wAx0qhYEWAo+G2hbAke9D9dt+sHM4AY+yVYiYAtCER2jWmb
vX7a8tMraPeaDqpss4aCriDSIP6rzPeHtf4rbqNluontsrqnldnErsAj8+bF
CKYv05Dnrer2NT5KnM5q9Cg4AhchrlolUNJq6yTTZfvXsXntRTEC9anosnsv
jH8E5/80rBNUGu9jG8VJy07CxKhqhS+e6WWVqR0H0vvvEfgDh4M+rJ26rkDJ
47VVBrTShgwYk5V060TO0ibZ8UkK9YDg9Z8lSp97adGt8N7/Z0zsABImg7f2
xMayz4ySYLy+TDUOIMtarcMcswtR/z0Wlw7R//dD79tHyXN/JkjcNRP5zuyo
6DdgEJQVV5mSX9tKgxQDfNjYEP6GiyBdxE5qiE5znIcSPP98dIB3yFYMPjuZ
SAwnlf3DSRcJiaXDhChe6RKHB/ST5dk/bFtfXXqJsSVkm+FFXSvoCJvh/odf
4tkqiZtdi5/ZGlDHiLqsCVfXHx7jlcmSii6jxz3LxGrqpMobQiBAXZ/ULPca
SW9+/aDVr2PuWdGWd2Its/eB6gA4jepYvStQDOVYi9VTL4niDj5xHBEGVjBo
3nrqieaZBieU7BjCPH55RU7ZOUxeZPwa8sM7yky7zaAfZC60QBE/5S8D30HF
Zx3QzIYuOBY9y5ODFkWXzrnwixPF2JNykrHRgHjoPuwfAcQuL9kP2H4JgWHZ
p2nruMUPsBYF+jkTcI6ZURAwt8D7BeeTO88Ukh6sfuEtQZOHuOhGMzesYfmP
Gy4Kxh3Cj01wxbMnacsJRZKM37KsSLn63PXTRZ+uP6J888Em8wOKT89MpRKV
9g/szRcRDY9PWGxPYA2ULJtutvNUkJzM8g+F1Qw84P8sK3WzBNPBg2dk6RNW
2wbgKFaU40PNSlATy/AXebbETBgNoDt/MNQ8fr+NdE/mijF3KhUaTZtDMPGR
R8aw8ONMifhtijZpaklSOqDPq3MbKlqn7F2Ox14dsI+eEtv1D9WjakqjnYP7
38dxR69j9vyawqKGDHqnQO6mTcxSYdxFLp4pMrNdaf8/P0kRg4oGw6pv6IDc
yQjQ3fKDJ8bRoHCV5WjEV5xp6CeGtzCC3b4ZxrW8uOhd7o1pmL0PlhR8TL2B
RHyxipPvcsMfBNXFc5PYaRidUFD6+O6X8dpBATwiBMx3pLBmdkeFY/TARCQ2
dYTh0Us50gWpPMPkrAstb87CgZ1049bS396StipQnUpI4I2yIFLeM8Zj7VZP
P2Nyk0GJdZEMrRKOdyEXuITXE61uYSDFViFVv9Grr3mWjO/TAe0dRnOOhwoH
FAyoYUjJgnrKD3j7nkiVLaFlvLR3gGAKrzAqQd2U8photx2ucF/iriVgqNwQ
iUFKLSRcC9OlIwkqXAp6NYCUiKytL3mSJ7u5X2SBhUQFIzkNePZ5MnQqTyAH
khZczG8+Y2JSReuibioauIzyEpy8dK+IDrRTO31oiZ/bpG5rBt+fwUoqvj5D
9VY9fvIDOeHdaNnlmYOpLEihzG9Du18KLyuRNxeb+JODisIRvx76Dw93s1Nk
tK4ckOhKEtcW4D7SQFJcxB/BiJgCPH9SomkvshU0v2VtRp1nF/MBe1kxdtvr
J1GHT9C4RUfDtVBbUAwcyCbT2S+5Kg+WQgB+m+VrjzKUnyE594OxminrjWKy
9HHyx/DopGn7P78ya2LRJ4+eQT+L/133mlUutxw3OZYZ0mr8ah0EDKB4FwP/
cFGyeHpnsisUCq0Q6IJn+OVTtmwaKeQKXQdMs8CFRdknnhpCh76GRpYUMZXh
RIzqDhd/mjGz6NpiqoEbwmzGJAB+3lphQEbRZwisShGUL4VV9XrP2c0/5f4j
CBC5T0VCuIhnnLBGiv7N08n8SK7j55rvuaelUcPxXj96h7ahI2EXbRV6ywDS
whASLjegWC6XuX3U3R5ePpF43ceAuyLm0VaBL7744Hmn8MqwwnwBNQw0w3kz
nKDimtmQphBMnqmE7SvHjr8LGhqg3Qwuw4cXczRoEKIBBqtQa6/fgie9JzHB
K2ptb198KyUsfvOBMAm7T9SGmm3DfaR8Sya/Emy9vQITN9XZwHipnx9OKEhA
XzwGzQsxk3cundY/Px78wKOi+N0OncKkA0cEUu1dRpJcjThWeNd6dglv/WAr
+qm5hEciZAwxnpidwkNePT04VtA+oH02T8zZ63lRRrun1fLX+zcr7BrZhMLA
dmfcwO3+COOpmSqB/WPqZOHyFpgaYSgfVn5SNkaEQhbx0vNz8HJ7CvfIRpAH
fikLemt8IKoY+Dtz7kQm4cxfYqFe2g+syT4WVEdCQKZ+6RKZTnjC/TT4H+VC
YsbBFzXB4Hsu/gn9DO7tYk7y9Nu9tVDtmkROBc9H0l1yzGxa7zCa3mfnfKYd
TV/LxD8IL8ABjanc6UbF5i/wkoPG4Q7uTSt2zpoFUIiz9nNOC0TMqhEriTgb
liONfLVAGvXjlmqVqB3aYO0+F0iO8PeGGRYh7Mo8zySxGAcLs7F6dSl4azrG
WzJc3o9pWwIb6qZoGuPoO1YeFq6RvqGFtajnxNarMoFzwFeNCvCEBZvYY3Za
wUWzfzb9JBS4cNJ/8uru+SWAT05AqMfarfrX3dYFggjWIq889bUCLDunP7RT
g49oLnjTkmqM7FFtOsDvDa2KOGCQN+OW6u1XF6Rn6jZCAmx2zsT4s8ByCbTZ
zZWsrla+bRNL/sVtnaaH314KEaw9Lc4+1FpaQxdrmvsK2wvePhYOYn/rjPBT
+IsuczGybcPn8joLr1Z4C76uwRQ3aGwwnmPTQImRiIUzTUnHEI5q1aOq2VJN
f2qtf5/TmipyHw7QbktcQft64jHzFY19VWm1UZ9onXZUH27VC0BXh+B1zhSz
MAeFogb/uDEzutKgAJXk0ZvXRcanvjIWmbKy4/3i+6l+Yxgk3S03WOgjW2Oy
fT1135IPt5xKSptznZPQfvAh4MA9GihvBGcaPYdFTX52Rseq0DDwp4IDd6SQ
LQtJaFsZu8WuJ1urCoRDKE8ej8lsB7y/0CCRgRzlXBy/ql7qJOx303b1VR16
WF2Z9IL8kqxBineH/HhMukQH8TK7DRS6vDecNx9NQiDZfhIk6+wR0ZJ9YYgX
dIUCOevi6PA4Q91vUIIQMeszGZAKtziPmW1exrU8l8N5mtFbTpDHZIUBhfdV
RXxfkxIycUIdy43aDaXsyspB5fsfNRWfmXU2if+SC0sV4T2aV5rspN1bEL4s
3JMl0ALRqgOfSubsAvv7PnumEM+kC9ITZzx7B3u/VaCbmDyWFud0kFQAVRcL
iZRFTVfxORcVHkbTGwLDpGGOwYmCctAZY+qRjFpR+ibxgJCUvef2/6kzAxNG
K2hHKwYD5tokPWGaDQ7JQH+jOOc+3t4eiLOZ5QYTrTW3kunRte1ZrPfZsEcG
mIH60vw7wfn7XVC6ypeIskHMXMElkS3SR+/Jr+DbxtHwPPXDaO5aCAr7f4U4
xlm1oNVYBx8USFaly07o1s1k4BAvXBAUBNC9gxJpS5hvLYnm/7Y9rleAWAwF
hMpDhnDok8v2J09ULWnmh9SXH5IWT0Uodd8V1GlxLyCa9vxLIlaWfZjeNHRR
/TTokxQGmgwKHGYZJMneQ6d3eHEw0NU/NNz6MMXy1ITnAQj6Dra+nXfcGW/W
LnXuRIQuXTwLtIvnkftkIpYmIB5nrheZUogS580ekluE1yMeoMJ7hosrLjW4
vwrC0iVK57//o/3fJqjULNbztaqdXXgWAW26ODvzZ2nh0JRG5484u9NBXAG8
mhNIFumRRGhesv87P6vpVEicUAI8W2TS/3b8NlSf6/l+TM/uo+25Pqyw+PWj
2coEWsBYbZ1+RocAX+3GbcS6I0lSvWpGERkTtnSuusCAp4lAFfCZv3PJjcD9
qu2ekPPAG3s392Hgoqwwbahxhp8wYyai0W0YBgtLVSRVc2QT4sLHRmThEem/
Zyhr0BUbxPFVNeRt+EPK2lrQcVlutGFe/qm1G+6W2hWoM556Rscu/6cYcNTN
MgSfSvhFchzzXUaVIdH9DINvq97V4z2kgl3IqVlUjASPD73iYaKbBGf4werH
A1RSTqtvajXPFgaF9OiPcWzvj52cEot2yvyV3fGMz7kxEUc+36v5DMQ0nwar
gQHeA5+nPH6z3Ly+9fDyU59E6HvT+dFCU9nuZq5BQgSFLpOFe9te7howov7R
Jvk8SFuV8V9xZRWU44ii5Mx2rgZ1aU4MK35VQ8xiZ2FQHTTaJjS27gN1Molq
4C/1KT1Zfz8ejSqV7J8twZi9IOBQbvwHwukWmOJY7ODZwSajNI0ks+pWuyhv
JOoa7hODzl1E14Ifb94MkcH+6+dKlDgMDkY5wMhR8W9iGB0yk52BjZ3Gr68+
izn/P6j/wMfGyN7PYQRRcK0QgfGESBHPTSCdHe3wNlPRpMhnsv7HcAwtEHOK
1iw34sm9a64Z+EWi2kGzE24WdTbylq/UCuhIWAZgL++4nkPzlqtQdbsauyK8
RSaMZjTte4s5zVV77HQdpRFrQeQdS/F4A0ReYBkKM0iO0ZN82myxp5Fjqjp0
e344VW1NMJJKn+k3T9xdV37AOeG2HYwTBfmp6uohSR3a9keY20hXAMjDy+Jr
KCZ2OgMvB+Gdtu6a7RXT3MxqqGVLprFVF3bwUFRLiQn2UJGCUYbX3dE/4Qq1
PEXE9arLNyc9Sfi16RRrahPLJmbADzZ2O6gR9iCq5ckO7YjL4fgBU7hH8rcQ
Qqj/ugWpjtev0ZJiPgiO1N66to38RbbUMibEZdqbH8N40TKIRpoG4adAGx3b
5YZ3Zf22PxaAt5JM12MEkzM2W+9X6tGIhBB/Fd8Z6VIhRrNDkmwSX8rNYbRH
yp1uRkGygsf4ParYeecvKSSnnLetCnbEhoy44RYbchrDi15jswHofV8ZZZm/
vwMaJQwzfgSrIcsvGfb45v95LUdrYbUv7wJ44zuWFAhcLV46aZ1vZetEdbmY
aNKgdkgxX+r/Ur0Gt//6Voc6jUf9z1FaSE2j/t0b1c6GGN6ocvmDwpSZSpDI
xPSGx4gU5/GRtxdto7kZFtlMacRz9aESTwwhrfvA5crI7t7KPXf40ZXtPeq+
NuoN/NpXs1FvDzvT4Eany7iu4GHjL0SMhh7p2KE2MsLXAq4exuSeH26TD/ZY
buMEazcMHecraPLvQyQzpanbOA3+HDE1NIxs76R/YUCQ6XVFW9Vc6sGb8JKR
uIkIDtjqExwEN9wfEjJxPDOAGBxU7OYg+FOJpTcp7bTLzu9s5GK5y+bxv7LD
q6WLjDr5/avz2rfUJp5qLFug0Sw3Hn2TInWNEx9WFmdUPOwjYoUpIZw7H6sp
4U5xH2Zs5RercybNp1tVeibcMihfv8Mcu0Zt5RRlZqKSj80iVQWagRe2vytR
XP+aN+HfVC13TQf+XEClztaHXQrYxchIr57a8FR5R99jqm3yRvivdFOyNMzS
wSq3VH5JA4b91jxH3tns2PzXdoVanymeN61j50dISlVt28zo/Mdn/jH9v+5N
u7PAQPeLZO5PVsbSKueLoKkB2UKpF+n0zz6Gw2nfDsA7RUNCpwEDhbBcyL6g
Fc2La7CNLnqMew58Lo8R7iKhivfrhlaCrPb4cI0yBYEUMkNu1vzCPg538kxj
xyXViSKNk883knKKruEfRt6Ew1+kEQMYHxRMqYDy6I+JPA1rt4lOkZKKF1gb
muV3vFo9iWPxYr/mUfKBrL34q7sLj8EqDi/RlPovh3k/wxSsv+IGbpBkdsp9
3WBCzZ3JOuDK/bL81ci6xajyHTrPbnZqNSbSQ1uMfkCrZEgIeMm6nsizhA7D
kaXhAi4WohipdhNP+I8unkdJ9+IU2WHB9qUJ3sXxo8AvZhK5aHsf2f9tvZ4/
ZJRDbP5z8vFJqrmYHzBE51XkD94Dkle2bUOG9UuDjJY0jG7/vQtmlpWKlYlU
GBhgxcE4/Nw7TNLKCh4pf3eqgqgvYKM/4nBMDl5wLJW1R33WKuXev+MaK5B9
zcV27Zg2RteMVoxi3o8Ud3WR4jt0VyuCXIgj2KXv0lEyRLLLetj+nDwRuir6
R9D3vS2unO8JutIWqWnV2/5cTxxGryHVRJfcRR+aM848UiXtcpdZOUTter+b
jJflzhZiMDjD17W1/VkqG0NFdFpL9QT5no48w4gHTeYGCU+wZdGdfGfpCkVZ
1bcaE77Nml4i1pkOK9totHB72l44hlwPJLNIqeGT+0PVYpuoKLEaC6r54BwB
U1yEYjRFi3uj5OvEF3FD7siCPDiA3ATF5DuE9IlMXOIRZuNvMx950qgovmnI
NeUZQ6D1NuQAWUnFwXC1yKE80ZTBHbP/HksMDjdwUn8n0ppsQT6Lzt3nEt4V
3kzlEV3YZ0eKaSMcZOXcAkJ8l5zBEbApD+9G527PX9nXkRdIcdPyzM51heUA
dMUciZEEPDjb5pqEPqC5PFZ1F9S4/QlgWLQ1vZ64+uc10iVDbu+yGBSL+Ibr
LbQwlkFpDcBdytaFDiI3bK9pkrF1ZqF9Od10sIMBvxYqNH7zOXqeno3EmV9f
BXPcRASFBhiCW0mtQ9AS5dO79zVX6kdDtRbW3hU0v4CV6yU2YMdvZ9dQRo35
+JQ/WwbtfcofGQmo6PVw80n/+9R3DjRoyCLl8AXY1piU2BJNujSMrKazRSom
hqVFii8OOvgzGsRcmCNbW2L7oJMElMnGDRWg523BSbdbf8bzOmy1O9cSy3Y6
ktfyHkpNHlG+9TqrSmK+i8p5vJkLERW0rG693YCYecMWE5vueQ436FDCRw2+
GlpKG3QujKRSMnsmj97+CY4ZdJEUzWX5jE3p6BY9iH9ftmL/7sZPKQ42oHvy
QA1VVmabBMNn0vdGwRM69yPu+gOvUFH1O5K/459nezj2NE2t792BTaLwDMf1
kqqsrwYeVIcvEB7Nz4LcoiLP5bpar0R3eGtNzPfrXiUEQ7TGOUMlkIZRXY50
Q3QzaQcCI6Mpz+tqlj6efOwBdb8CZvZkQ8oeypHa4mjzIME+6lhCnwktaJkz
MmlI76AuRe1eI8KKXJEaeZMfI/nIGVoUUYMdc1Fnh3AEmkz7eEmO0xhtYHQF
s5YEAlu2zxpAAavSdYwRuled4n41SIrdMpNJ7No3gMj/Bs53j2VBSdInwAAl
Dm8kOOdSzuxV4GlJbNa+3tlPlblkYwvGnuh7MPoivSxDD5teb9ZFt873efSX
hMRQkFMQ+SAXRWKjATNtRIcHyd7B/bpw5b5oJ80QJyauVZqZTANfFkoNw+G7
r+CzqZfCvTSug3hmuNaIBDkqN74rcslYst7QLbz2Q3rLCd3Y6aQ8ofhrVowE
L+RVD/AG7b1hIkFLirxYpRwh+hKsq0zJtSFmwWa6hu5cYFTVpFvLCp62QidA
1N3rZFaEkp9vGtUucXkMdEJcyXKEvbJkb129rfwkyIH+s7VUR/DiieWrxVsC
q8HZsjPk47/ts0W4JWJpcaUGE7Hxtq9Xp7owp7rQxOm6F6WxexE6QCjk7cES
PeqB33VCKiETcJU/25e0iWBWGF7PcsiStui2jKpqRWV3yhaz2HU6WHrfT6Fn
tHMNk4CK2oqmZwDjmLbcjZWRBDq1yQPAUh3N3JgVthK8sWmWV5rEfQ4KRPuq
HujkBMajFx8dw+7tMmehr4MY5EZdP4fsWymMd0bIoItk6vqL14XbtjxcIgG9
086t090K8cOMClh2rhLC0dOO3qV52ICfR72KLFPe6cO1zpffwzADTpnfGQ+N
HgiAJU4UX2KgX2JCBlwvPe6N+n3NAGr/4msN91c7gnwHE2M9B3q4zTqN762b
YKk2e2/bci2OJ25sP6tig89oICDWQuxuEckMy3CLPj019Rwnbamk2J8IaNxc
QI4uc6MaKyAtLl/cVLquXCpGzljYBf/1l1+9ipCyzUCm0O+w34/cCVzbDhUX
K2o9VCQYKt/CBYeAY7LmYlEMof9sn5gukkm8HjcZH6QrCFPpZtizFIHIFKFF
hsd5Inp0iJhtnW8McH2C6Bdw/YNOzFBcpiTxck540jjgdAPbgw2PmgyuzRa4
TY8C0q60hOMslutu8tHd1jw9R65gozcrc+ccWOFHd5YW+uGimMrLPnR6f5ZN
r/v+NFH0WJfaorA3NEyVL4mAVerJgsoHRzSCB9FGdatI0f70h7zDvn0KW0+k
6YduHHKbAWqXlPGyxq7dkbip5jHAL+7BeQRBUCubsNLQi2ye0t2DHnWv/Jk+
MDYD/0seCuqL4w/Bxmut2O7ypuzLSNBbUBMjuYOqCbrwa/e0Fgxzw1xzsY8B
WHqe31h9BDIO0iwKcaVC4nRKFjVj70myApPzl34CZWfB9QlFHGb/1/dcp24V
a1kSSIK7XBxSLK5DkbhKer40IWPJHO2dUQXAtdRiBhartRhDRrK4kHYLCPEa
DiT3TRyv/ewoRqAD3ho0QP/zJuMjXluVdAPfZ0/5LVGjuAKwi8KW6BRJ6s+T
YdR4fO4bzTKihxpi8+n1c1eyuWgkUk4Sf1PoGgffR5NHROkB/rsinb0A2spM
3eiSk7uwpMPmNIefO5JuHQ8S53HILrni94oKnzVUAwZW6YxpuJY2t5FzE0Ju
7F0NNmF7MS7IzrqbU12SkqdAmj6C0awyhHPXa1yPVkcR/GFmOVGO/drPAJpU
6/jYkecAAM8+8g/IFbGbIYLrj/nSM78dapJkRK9G4rW9V1DhIZLHoLXYO2Xj
7usW2S8VDj/viPMg60Hi7g3DAEyvzI6CjG0rOCBOckr3WR8zXyMIhJacGDCE
di+Zz7niig1Yx2jJ1nBC/HGLpaIKQHTBR/U/GgnPmmJvp13f8+iYWSAfK21f
i1ElGF2Q0bcMlZm65lEV5ZRvrPCq/CcubfP0aWtCjkkY2NfIq7lnV0rUqgRt
XP28VsONSC7hpuOuFtYvMFpqiAJdpX18Rq4E+dwnfXU08/iXwxdmmVfhImiq
mzfYFq9svo8+SSjwsasfTGknzqVc80VkkY3Zi8aAs4BSGQVnCmLIJRZDBqGO
+H9GKCJSdaQah44KukA/WtbF5tZnh77aglGKc+o2Nt4jwz721/V7VeIn2TVA
dgrQnIpcBdTuMt283GoPU2Ohrc3G7Rk0yWEW9oU2UgfivjPWiJj5zarZVX3K
k2+5+TCVWWu+cqaoO25MT36D0x8CgQn3HSlVDgiKekhj4vuqCSpTHLdBG1zt
k6efrEiXCWXoJ0aNHsti9aS1OQHo+HFY9WQYQh9s7n+UMKrQ29NDCrTGJFlP
qnZFRADacHjvS/Df1gt/cbPW0MsVrW2uHEGQrY/AYi6KBUeqEvfimOQJmmcp
WDjebAl27ilts21K9qgT1YpnOdmhFXYv+ueRCzn7GAIT8g7SXXQx5qDyJBFV
5P5CuHzBqge06fnT+7PIRjETLO5VmxFNhB5FB+1M6L4sdpc7mimEkmxUDbLf
RdiFTpd8LhHpKeeP+cw79tbNv2tfcyQpG9v9bG4wJbHjEC+kEG8EavIiQaCH
BFmdnwpvickRu935uFMhoVMRc41qUDh7q+/IcLDb+ZfssQ3JnAjeAx+z2jc2
5Sz+RZw1+dmHu6HSveTZb8aYbxEPnQ9UG25iJlBjrZHkze2ldnd29fpO4pkb
dxvTQ8zlO5TIxxGpAwnRlQDzP1g3CS5DFt87Woi31fVKPcJYjjKhj2kNXxQa
7M2PrCpxs1VcjfvaNb5qlfCjQsxgH1+aREBSQbO8HlfFFpiT3Eqq/qj3d7To
i1S/JkI549eIH24oZUFL3aH8PpV82ym1Oarr5suBrwoGX5vPJ/gvrykem5Os
fBorPPaKCVPwQeQqKmAwHijPdpQMPwDGHsCH3D1MT64o9fHlihm/Ll/v/78z
hocbXG0/xF+zVpQzxpfEkdIcNfZ1x2+un4LaSZ3U8cljRSRl6UVkPXL9Szlu
sareLsRXXIWxHh99QmynZQd5W87zNYa3wKJ3K3e8NPnJ5iGzKznI5DPCpNod
+6cwxeIBCXmVceNukS0iVhzBBvOMe89vo1z6SQwPrrK0FzXCutkwxsfRVxQJ
j9zHFyNlOEDuCaMNpLPMF2IIPjMH97hjuAFpQKC7W+RY1FVNKipOBmvZ0vlT
Orar8ji4exZe3UkMBK/jwLptki46oXyxg19BjVVDGhrRM/+IlPSfeisxwPpr
xPH6L8VWdcO5AkWfyVFgdX2Ec4hR+4CQ0R0hpMdS8lBbVZclqvn57aGk03GX
pqXi1e8HpVeym61HIdK56prvMXG7LM/DFtf9bmafscTyIo7Q0mSnGnvbxtdn
OC1/UYCiBCTXOFLWeeZms3b1DdagK/mRqIi2u4rzNu3CnlrKk34wnd0Ggkfd
MRuriyrBc/vm+lMC5o/mDhRY887+WAU3RBxzBOZrNZs4yNLp2QsDhYCP+M2q
ZI/EsBiqmw738+YedtlQ4PTimTuRZd5kkHEf7fjzPEZqMDWCiE81WquT2BY6
eeZPbuGzrayKOsAqIY+AhF2qYkFM/+pYbDAaGVDjPinuct4qTXFhpnAmqvoM
WkeXIGZtGlJl+cURTevbvrLu6T0HscK6EEFeRBO2OxsUj1axrEg9aFFn8M1a
xzexNwPYbh8qgWb+qpJDnaaCQ0mCtINDlgTuuV81qh92iZ1HZePd4Wp+TsXT
WyjTUFnlvMo1ZFdTJcx5jzp2ALp4jPUsvgkwI6lO68PTDcoeV+Az5gaLOYA2
iSxE92NeEzceSsm+p6VoA9A6XJvw+o+YRrx1iVyxcdtOX6nPQCkHZLS8xDwq
nVdtDczaHN/gspq5xJUmBHPNRma6JbGpDoL/AgsdRvD9rYRM5c5U7stvHJdf
l7jRVo6FnM/2xgUyNX3rbuIU1DTYs45uUcrApGyI+dH+ofnX2AOAx5bmCHto
fTL+Y+W3rctknNwA47cxBgh/w7fdsmXcR9mWwCAlfoxa6GN9p4Oj8S030DLv
B1N7B460gVP2rjMfwcDFUUJI8K1Aeb4wJQizqf0ciLKbEgiyshaUUnZ/CQCN
CVafF3MK4ughZM9IV5k1wq5a83nJ9yQumuVnYll1KRZFHJFRRk+50j3yWKYl
NmDLeQG2tJvpwR7gb0QCFNANDDlMUzcjURwnoNSmUbe6LVsG4Dcm45jfCLo4
60wzD+qnBFJT4vwAQW8LLjTMMqzGPMyEhnfpVIESOAs+tWN7wDiLBpTi/Juw
0llAQNbjRK78gJONBKh5NCcRRg+Jw6AhN7lKMoD12raoTmq3Ek/V+q3icVJL
zYqJtFNVBIQDK2MrQNU/kSu1QqTm2PWXefM3F/HTHCKhaXzYioX571vTerzg
u/ywdyJUs4tDcNrEud5ddJLrVn/gI2utg/phDhb9GUPK0OxQFtE1oO5d/9in
dw9gtjW81DWr7B10DIQ0uetlmUvqOoloXn8WidW5hmsc51O6S5G6takPneTF
zt2OPOiR8SEofxEeRzJJHsGVRjFEQZ87GD85WzNTLtqFROaIzVOg8sKne3Ko
+NhzwOqE6hLxialj+tTN5WAtKx5tDMAY1u9/YafeWoYaTEt5PJHwLaZLzYvj
V0ZaHec376/aCnTBG9PVf9w2xF7h5k/nr65B410/fMdKxIXhgd31EpLG7Qj7
5iZVmKlCioUbrkOEKupcJGZtV9zeYN23Q/sGnjYXiFFOujrAXHF6itlVtbF4
Jo2pvqUZEi6TWg3ViNbywQJNvVUfxj4t9+CsWHe/Obpj5Cm3NXyvX0ggOIdg
gkONusu3hGQ3ikKG2IEugT5/ou0CvA41+R5gEVqOA0m0f/v6Re2KY9CwtocC
EYsOq2/EiVawiVQc8fquBqe790NYA84o5AX9TPDaz/fxjJkVrkidn0qZv9OK
N/s1BuGRgrMjgamoCpYis2Y+aFcdm13ZBzOLEHqfGUTwHExuPXP9StYiCL5Z
GFKAHnTGBWI5W2ypJK0eHRF0UDJkLTzfI4kqmOsov/XyjjnrwWJlBQYiF9Nm
m+KzQ/L645PsB0YqcyXfQXqWL9eXN0owlZqlmDvZluBx+5lYNaKnlJ9Jz5J4
HEO59+y4Bl06P+EZDLQAC4om/3ffHedsFYJKSNvTE3Ka3P7pE7W3EM71xlzS
fm/GC4hPgyj+kEWoTNkmQfS78tpB4B5zmzQlp38tUSVs8m/Oamqd9kGfEU7/
foYttj1W3F0es/czQviohqUYvg1otTMlCEWCrsvsT1m9GcWFZupl8RdtS1yz
4ztgRQRoAWb3dtQb3Kxulqux4wUHm1gI/LIt+hPrhdT1ZMzmRI1/wow/VA8c
47Ybo2C12W2geqFPZc5caiebttHJk/fRiZPlOv6dOwOwufNLefTM3FFAL9qs
LyOkFb8GKvSr+1vupK31eRHdTTRss/G1kRdvAXQISf+ybohdEC9DB/GkBIJw
G/aftyRxsqy5WPaJCyA03iaqDB5mgyuy9SKwcwg6WFc+sGV3ramrA7sVO4sl
fNTk9MQZ6+1iEyRCdKjHD2Vjt5VPVKdJVQ5XqQ3wwiYJUxm9WyI2VjXPCDj2
6lPMgiscfU3SxaPHnqxEikLqE8pGDqTvWAm2aSvS09t2Q2XIKMvGBcxKkXWD
PDJqv/c9JkjwMD815lUVbsGLrc9g0YSBMNRZZ5En95jPUPMBSBamkS3Qpmhk
BKemBXtDQDKtJw5XQyIG4H4keeT/ocrZ34SIUlZMRGrUIeNkFSxtq/AWUpkj
umgiNXnwINmiYLuf1GJfQYDqo6+XyDNPD8yzdxdcrnPOIDAcooHIJPVPFf1z
XFT8T2ITeO0ZbsZRPWkaOWJlRPoDcZST9DA6VUGxFxD2NZwC5c/qAS3CDJ/c
PXvV1cNDfM04AN8OSRjA+5HcZW7/m87rjH/Mf/a0EMf/o9P9dVcTtxNYOo0f
3FxTXjI1RFAQc4Aayvn+tr8R2pkT7egvXrF+5xMuRB1HbavzBwLhCwTZSWkx
Le5ww31yLxohEII0DoDafK9bEZj4QF26+sNviVBQ17NjuSZzM0Cvmb2BhiV5
pnhzPnbcZF3PojZ1e23zn+YNvdLJWCpLtNUD7vbHL0lXV6d1+ErYPzRH5wyr
4HJNklwk1sFKfRoh8QYQcP65eD7rYRdLntI8ROfdZ6QA9tkyu8cTDu9/9DKB
cqgZrWLGUrt/5SdTRphtlKyBQxHCG0/G7QCMw23rxzniL5NQ1p6jrmkumeXQ
N+QC6CAD+wJ7uWsbvvWHRHShUST8K5DjCTmEXZRmeURMtqA0k1LrYhhg3iso
cmSwUY1nRSzLLkzCKBUxZcF1ON50tSKmKWpFHDvw2ZYJzaK+u84soI5VHBVZ
kcef30Dz1ZnIX8CZfgna8W+iKcTjk02cUcxQG03eklzR0iVepikT9Ahsg4/B
2aJTAVEuGoRowVTz00yR64JHRDRyJB8Kvu8niAk+yZ8wE5cLhqnlnFFTRBos
Yde61d/LmhBC+XdOmb2d6jeQqw8BS0imrpzVcuvEJvv1c6/FYhn3epwOOM9h
tLJxJRL8AOeqcGcpmaxEm+Kj1q+sDQ96u8kXN64+gs2eRavtBaAIoSez8nPn
CXLgJNn1+BbPkt/GHwWM72vnW/gT+jIvaiwXQZfRfXcmGtDvQzlOGsUcWmXx
7sIOnsiMm7xJGKzDWlsHpaZYjE45kNePtNNRh2d8jhlPTF056LxkIfmZdnEH
uzbqVl7TLZ6bAa43fHq9P8eC5dQlHQC7QpvUpHyHyT3apfktByQ/OqgPja9K
Ti5ao1wGfOyGbkZWXeTzB+UcTMbxCdCqtllep80qFcIqHg4Iu/qIIudTcdu2
y/FjqU8ouX8Ya3ChifgNBN5Dxd+KnZX/ir4lq3IFre0HcVHZq8JeHPEQMcQ7
zmPNULVzMc7vcB1i4qdK1yUgMO+S68KmTzKm4kbbEWMHVeupIVLgZe9nDhd8
fGgm2C08Re0JZgr/WI9gdOqpuCQyv2URPqJSgZRT781igqkI4C1uPOcPc+P2
Ed13VzNhxUZmMgBYfqXHz4EZmf38F5Et9hqQABqjqaEEhJDH0vEYwzlaeoSX
LdzJW6WM8oiLx0OfqarhzrsnIKy3CnEjtAM4OwX3E/1yCqAYQ5DqIAVRkgib
acwckxMSo77qz2955/7CnsvxaGhKrETMahQxHRkgwg/IO61p9eEePVxj17gf
s9oj8CRmBxLqloO1Ctr14VH/LtTl+6gxPcsaGSW80+Wjhl4uXjz6xDGrFl4I
E7g7ZCJSXoQ7dJd8Nq7cKhL0fOlHXwDOcZoXHiOCjOBk3LFmv8UiKNXEgCZU
HCR4qSdgxfzL7SfdXw+5gtezPIB1MfhaxbC9dYLoZIiZD3A3Z+RiZmJ2WAou
4g9HZ0aZzW0HGYkN7JSU1FvvVqQ0UJvbW8U6m13V49VZVr3qKMHTMnx94T+N
i3F5YonV9rx2kqCVNAzrhTzzaM7wLp1gqnSTuJM+DTZEs0bYDH5V4icbZTm+
7a4FkZ4zrK7VvMKs/W0jG0/VHB0n6ymJJH8NmdaGqIIKOA9pPO5/hwHQD21r
7Y/ruDzrGIdpaZQerT25murFw6MQkI3YKTSDtqjB/0Tj6jsciZXa7x6t7cFV
8Wu2SE8gu8cAr1L8wGugr7oRSdlKlUXnTQ15LPyalqVB//gcOOBhm5Xfii+8
u/1kPgwg7+6DYWYKNzk4jKRhaPEdQqHZHL6rHDSnztwc4ttV9yMcqkiXrENe
qcFpT654y/Wz/F3sB3PgoiakEdKCvjKHijyFxQWHbH2MOAHmgZ+HOIhenbLI
E6XB2dgCR0TJqQJyXOQdvQd3LvuvYLY1MA04I1UxH3ms9o1Bih9vHBkRZYzS
sZTMFF1MUXB8nwEixMlKbjHhXCZf2CVV95GZIUbk5zMSjV9tlDa3ZUwvgJOA
2SvBggUsjTsZPvh2mRG13zRxSev0IVcq1G4NPa+kBZ8QtDK9xSSFF+SetlOc
DdG82hCwn8crQtHFmam5bo1C7Ltx/ZD3fCyk4NB+7SyD2K/u2iKodsQ5fs1L
UcjcLNV6s1LGzGIqsVjgwcqk+RXrkHeZMKkkdC5nlR7Swe1swAjAS+JhksDN
vN2h0WZm/NmEoHRGC98JUj/cwU+TO+Ek4IOHQbwGxJ9Ls3YLy8JWztZJZ60E
TTb9UcIdK/FXaYmNHsl22dUs+8l6by0Avv7uwpzf95DIMPbvCV7IOMrkSy7M
ns5iEMdoerJGaeLGQ5f17E4W0umpEONrz/JtZFWbC2vC4UaqaaSQ3ed8Dju+
N8b2o2ud9PSQTax41mldLjVCQysNZu86hUVqgkhzvQ7fQ96VN/2er4UuOVCM
pj45b4WG2NGAakh7DYqFqkSUkcUTOOqeSarbOn0FdddQufIXs7whcgoNbov1
uXu0CZgHbpdF0zV0dyKsopwukNViTUcTwg6KS+db/U5A459nNlyxC+LzReAj
5z+UnQIN9vCDlxGACooaw2KFz8Cqn2uXtnIAlCcPszTLj88Hh5EemiBC05qe
GeK0wC28PXBobp32DEMCj1PEYHHAWD5pkLdvPG1KtdBYAUqdRZfBoMFxe9OG
K/ixF815YW6oVYalroh5In+3O3Wf+uVgnYsJLJxQ+11nNBWCl9quivDypQd1
+9sGwEQstULn48Aj9S2BgK6OlLrwzHtnqliFU9lDBkn1+UsaTk8RNBQEJW/7
ns7vbZ9D2sQqjdPsj2Dgs/o3Pd+heaLcfZVergjNn/rRFqTBevMn5KV1s/Pe
yTaY1xW/T/MiG9/QnSirNs/bRH5fIHtTQ4ivstEjfOjT1P856ihzAIFRGF2j
nE/C686Q3Hre8j9AOVSZq/TvmnT4mU1qGT1Qv28fjWwC+iEInDAI1lLmlHer
zXHB8VDIwvQW2WhVJZpOQodlvq7qbf4aw6DbJtfftYM5lIo1aQDrkcVRNu+d
bYXqAu/rv1azyuYKqwneqQmWg9+d+buO5BUjG/f6bqPWAEdS8hXi1B3dnCbW
cDyxnj8AlJCV0A3EsPPJb8WGGANCQCVQxnJmxiKFv7IUzS4i/HYnRF8KTb/R
vg72qQZZN7LKItumJ9bn1RcY/qXJPgwdiW8n6mYae6r7BkDB84HMFLVeGlNm
lLDWpzmZF1e4+j/YO6g5EeL0zySI2BG9fumK0YNBpGUq8OP74CWhEpIxRHUY
cICJM/Nl1yLBEC7LAmGeXNgXXNbfluC3xkcySxRzuvFtRmAIqmMgI/WoMDKH
XiWV+KNAasldaC5P5m8aYMdrVjJX0qhaYyMsy7Snz3s89cBZFaQZn2Qlnwjq
McfePuy1RawX/MiTxantCVQ6IbpJzLZKXPsZqKn0u8RS3NAPtOQMeKBLHM1x
NS+rbZ182AQUtfYp5khg4WV5HOU6mAirNYxZfGPylponjVSL128tfoDjTJ4X
4NbG2oiplm8b7OjvyUoOkwfOIl6GgMshJGdr7wgWHZ+dFticCvZxVaMV6vF0
+I/oQg3mkmE5f8HvCeUsk7iEKuM/JTgCWAoizfNluUkwySiW6F2VQYUVSO84
Rz0aBeOjv3RVzvYcYz5wlnUiUtQV2pk8JC36JeUoFHypdEHSueR7X3377K0k
OxaFUep0BFcOKebJHZ/VBePN0Flq3HSfcjxU8kX30P2Qw1J6ml74pDy2UdKf
Bca4lz4tn9MAe/KSg/BrmnIP5yDWx96G4A9c5LJ/QdpGwUb77Mo5ZLGbXitq
k8CpUQhZhlLcPQtBdMLFBplXBP87aKntWLmHXKViXWH6VI3HiScVcCLTeuxs
vHFHpaaxDifWQ9PwageQU+LwrECP32od4txN5PFotYDzi8qiMeKrLKblLh08
m00o4zTM2BbKR9jYD1yf+0h253unU52B1TP/WoVZ0LJCwlAx74MaHv7P8hiL
h/zaPlalT22LC/+HcrSuwN8Mg1tgBDJgscxZ28x1pyiDprS/FtFLF9ocG8Zm
cm41MLz9sBtJjFnQXPMEQSej8kVFixT+NtR3KjKh447vZ97uKAoxcnnYNwHU
QUYOjjPnbeKKDEdiSCZrflOKHEWlU0QKKtEK6k3/aotGwtj1DnfDZPiiflLl
dc4dw86Wx4hVvthwecttGou9DVUXtUXZIke3Ong0VJ2uaFIUsWY2tY2MHyp9
FwvRBtu5RlNEqszzXwnTkaSkVUcCV3mKxhbsnMPeOUNsuoVyCSr8nKP7K3G+
HBY+bzvdSaKTf8z+bfVvPWMoEJjNrtfDlVEvoyQA3ncSBu0k+d2D2xOwBunF
9WjZoT6h8y3Y4Xgv8AyBMgNl0BwjNn0GE4/63ZQD9lpeXh8voIOEZLPtEXAS
bUgWE3XDIhwdp3dOflDdLFVhsOW0lLNAqRhyeb6r4+S2OLt7YIDUZIP2Nnjx
7wgbXDLFlnb0g4/Ghl4ESeh9P/aOVy8WEMxEhLnHFFb7iIRNou3yzLde7cUa
IL4nU4zfH92nNgYW/hc04GFssFU5qUOoNHQph4DTMqkX8XoZTgTaL7y6+XsB
umbIPegYV4CKPY9dlu1IZRd/rkXxLakwLlswYG2p0yY9HThL/tzjmHOO8ARx
b6T9f/uIIa+6et4X60yQoxF4KSMvfaGnDnU2pek2xfj4YhLkPpuAnAcRB+OX
q49qb5UpUt9bsaaq1bfhHXI1s9zAp/1KA0/8zl3bq5Rj1osEgWwQCEwS0Eaf
ZofZ6rIhHjjh4vI5IW7DkUBH7NtFIIsrA7WxqPSfkGulMGvD5U0c2yYIbnRJ
GfMo7zbCx3m5Jtbb60lIXr1X5zq9G9peTw6N8WX4nVRQI90qhlzj5L4A7nrm
GQCRkirK0Ne2eOc51O7aLl6SdN4HPLCsBLH8BFfTG8oImF7a0OEck75vrcaI
Qw1sJXPOdRFziNOg0G4pveIlx5WKXwXi8d62qNFWZ9dF+BZdulvXm3ss6He+
VW+kI7UxVWLstW/ONiprSks045IxGhS8YALmI13cSnHehSlAJyYW++J3MLMu
GqyPwcKXE/7qVp6oy1nhJ9jaLy+fdkqwyCaFOe31hdqangigcMNfv4qJtjzl
5/S/J8R7cATM0iuaFPD43sNKZwfYh5eSmJ33w0ilg19OHB3dxRcnl7sZu+LU
HX2pV91hDkdb9ALURgXjKoT9qZ6JjrnRLRCRmKwLV3Y3djtTK9CGzhO7LA21
3cvIprhi/3/MDnSaXvkKuudm/AvRbH+LgTR8cTfY4IQtAokMrsCyjFGqAW/B
Ny5DQQ51wN8cszc/UJogMlz6CIepJn6liOn6E4eYTskxBsUs1TviP4DrOhR4
Wie6mZMB9jJtZ39GZbgvXqbdQG8/PoIvmYTVCf3d8jELA8GJfVPWoNyxLjfB
JZinSJpB8M99lWBCF7tM/paeFkDRiGV1m/SV4BSD5tE2dj+B8e4SbDH1vA+D
6NvM5qiCaizfwJ+h0elrWy001/zKUh6usGcInDvxg6pdK32eJvX6xwxTH3HY
MSZdJy8lR0FpyZk0HJiFo5qXB3u0ykRGueGH6lXTOQBDjolQWZkYT/2JQRa2
HvIedSzWyq3raLyCFxzbIHZI/O2BOwVyX3b9mZ1xANMZophOva39yu7K92aM
BDJPaVD0IbKzfvO3SbBJirVkvvcoNWa2VXnQJKyltslat/7TFkz+arZyqJvK
+L/MSfTKtQGL6xpo6cgcLKQ1SuzezkTNPGPrHpxzMY4MF9PDvcLcnkSrhq1W
6PoYWtPwD/lVVuC/3wccVVh++hAf98G3+MCUZpoVS6vwLhqRd8wWtiKis2lc
rMb6raZPxZqSv9P2Spi2bZh60Uzvk1kTU/l5UYj1ly9He3uliVyowJtCvXAC
Yn/k+DoOCcwLWgAib+yVLSNss9uGXGKH9sK+lvcQcE2T3vCfJuthWdawEFyT
5JMTRagRnsK31bmpMp/LGA61Yvq46hv3VQRN4sP2FspjpcxV+vZ4RDl794Z3
WmCAyK37YLMHCHedcagBAedTb2iBL6Peber/bj8kbwIBUVFGObEkNmk2ASt8
GOqBFJZbz3z0oxLfe+lyUTSJJMvm5rv0dK7TXtJFcRge49l5NDgUcWvRw+6+
kIiRFqxO92p4XyNEkswCOCvWYpxaGsl1dv6U9XewsSgDOe0LsqPqHcnGKFbh
VfmBNeDQkRpWa7tjws8j4k4j8eD7J9XzSo1YT1pMFUEr+lfQESs1DwMWtzBp
Lw/7YFcAuZ/p/Rsz1fJyS0TXAjwrACDDQ7pfOL6yD0wFZsG2hbdtdMYclEek
0OUpo7WwIpnqDbV+tgbT6TBGb9L4y7NvIwhaVOtkMvH4G0iT3B45afMkgajq
L7hlE7e3+g/Eg0GjRxKVECDH6s48GAnhzu4gTH+L4+smiXhhE0nRrTKpuZ3R
W2BFSbrRGPWJVP1GMEJLlSqcXH8AuMuLpWcOOU4m++GQmbbmY1iA29eTEAgH
zdOBetZeEscfWHnDMxRHWvRCm4SbSGEXuLRO/XRf1jNnaDSJ8no83wtxtO+y
/NBrg31rJcU3Y2l6kQCz8v2/canw2/BwBI3MW1ceMpzJzfTJZscfIJVNoZht
Wr1olu/DmW0mctwzJQBr5aKyH5kRtb+ShEKLsJebCi1/j10svGtlwh6EaWMV
wYKxsZKdsIGPV3AYN64Dz988Jjc6FQFp1/khBIZRCNOk9i0kN571s9wUqH3y
1dw3z3xlTUj9i9LU45N9h5KzZqNOYf3I6mBmEpAhtcxkQ/zVqTyQF+otw8sN
70IcCwHTwl4WwwIHDZbsoRfEWEo/CrdcaaX4EFYk53kFeeYy4gXc/UjhINpY
FnlhQM7S9rR4YF62A+pJJtfDjq9xZLyAQZl3Chco0o3gzvadwq04uR93++oR
RXUuYepn8b3c140CgWsBEgeDLpuoDpFBbzO9D90UCDSnGvvOlTOs5X9j3W+x
Irja3xKdX7IQic7pI2XRVHfidWD57avcNGIK9+gNE6ThFLrt2ST8N8vOR3u3
C+Sy1QsfsosREBNCnRzer2QI5i5/bLJ8jrmnbC6gJxSsna3OcO7u+TvF9ios
gRupO70depziEk81IS+wxAfrk5OcD+5tWTxesqmrv8CtVlofVctLisYg7rJ8
VENdukhiUILuct33be2rOHIvUtcE0g+T3EoTZOy/q0z5ur9QjmNAvBjjus6N
5AvPMSXzN4DE6ZBwTL6DzY/qb7N2LkgVG6hRTdXqLLDh5P9DnzAZOVCeoi/r
0wG5w/NHk/OYA3cqamUA/CCPGLuINhBmn4T4bLoWRtM9L1wGIhdWwufOqy5H
ntKgH+fGJWQ0wfdsXNiOk7Y5WSKMwJEnTRYYT26pwEPbsyFyWbChEP9tomPm
leyCB8PjXek9OvQBj8wzVaJZll3SgTCEiGInWkwxmVNgp7GpJfIqujzDqjjv
Ztg5Xx3RVApfAjMFF28hG5w7binCv1OPvBuVM8XcPjLthYnEWtJbRTfc+JXI
2R/00LfeteDnRd2xAQr5nvMoH0//KUw0IgI6zMU8rz+uzNh/0K8B+z+jDG4V
mbPwbWxB0P6tjNYngm1l2OSk7wVzOSibcVBd3cViWCCLJ8cqYrpMeL2EZD73
qTriyCw2xsoSgLvaH9veNLSzjgOJt4dVMBe4LRcH7NT+vm7sqewH2BRPV4Af
xoNMduFic6Tfg69JtAqlEhZTg3n4rAX21zaaSPiCdz4Mkn6nhZ0Rb8Z4Ng1D
2d+EMtjoo9zJnO/cJrd9imHqpLMIvAbwGaS3EmBAEDvpjlif3N25QhZo0Fv1
SJlwPTDqkc7Jg5iCVBm7EnT4tVXb0J8jj2Kqj8h6FNyhGquLHo+Aqbie9qic
Kkr3XwkrVn2ORcB18IuQ3EZ4lBg532A4WUsknLzRHKCbxqn0kh9rh2nCdv4w
JRdCazSzdhIrkyPsutrRf5/O5MQix4UZl5Aw6EvJVC0aQLUDoVXSctlHBUKj
REa5tCWJtGbNce9tBLHp6x8b748ewZuz1s64xHmttAyqjRQa71ggOsBXSqiq
K+5BxJBpRDN5l8f5W7DNQxgKxFe643X8FcMVKiw9wilOxyZOyo5F68p2m0PI
CYNfd7LFymflraw5/4NJwhLQvDPSgC80c1JUDfR4UMakAgijyU22+3ncc9w5
7S2BfffgsGFJ+S0InmSpoWeaJsh5ck8qyt+3Bxal7NQf/GycZ40TZemy0lju
1QVt9hRpbT9/poBVceTndDLcNcDkUZIctxkGVenTp7x1XOzcw/YfS8E080bb
IizQoVN1teErcPNe4pIbryk+QsMMgFJdsiRHzbevUzWnype52251her9jyFR
9fYNcMNTRzPSZIRN/TCtNZb4tlt3/2q2Tl1luLeKTq9xHPPBBHyggdpFhAFR
i1wCjXJYE4wz/WxR26a44lLqW7Emq1rPmCkJZ6sSMjPsUD/uwAc2nInyrhe9
7lW3A9T1CaGtDDMb/p80eqcrjmRUVMj9fvhjh9j+tYVSknC1/dE8fK90LmFX
SwKXEe3FIbf5/l60KvGstGA9bUwlKYJA25+awJgHoGG5jnWedfT8DYJf/oya
kwBjdFak9524ZflqN9P8ZQMJGBB5s+3npPCsEC3xosEXOXoAKWEprO0AxAvo
Wtxbpzqk0hjbWxTQ2r3LLkGnxQvonbd8dL5MWm38yBv4fUA+woqomEw8t2d3
qoGorM15FKFTBDo/8xOMs0VrdD5hAfvNVIsFyjpjrpy8SStafcwcg/52nPtV
Sc7FBOqKgdj4r4JdrjK+eUslNG4wlg5wOkJN1Q5ezWFzz8zXigkYjd1/UlVT
EDgEWkdLkbHTLXuohtJ91vtgYrSSY6Gc6oEbePfX5q4eTTP8y8EgyxCZ2DgE
mcA191JlMBEn0J7I5Vts5wd6bNnwTqGkDlvAHoQGq0CvMysfuvIPaoSjB+nx
5yGCNn3TXTxLyFkjXU+mtLOAfmcQHWa495BUF+Vhzcu3ZTwm3msntQp7Wvkx
jzLFfNOF2J0FAfbrbZQ78Pq05+vT/y8z6jAyCpMw/VIaGEILoKk+79x5s9AX
K4EoKFKRujU3tJn+dNyUgXPKROkO3lwJ1yzY+tcTx2MZcWWRqPEpfg9Tv4bM
NqVcOxHqzLfNZJVmSppY91nElZ+VvJrM2EZhnHK8GR9JISIV6KlJECaDcwo9
988/8ACusuycM03h7yfCRtBxDpIzaN90Vq6mDLsNIsZ+pNHoa4sEpY0e+E7I
3p387HG2lkx+EOdjnRP+eAkepqpvIK+jHAps1BP973cQTysNwMmWI3jtdGvT
lB2Az/AB96uWJAh1HfDUs4pFYJsSc1+SOw3b/L1C0zks9UA3t9fQEDIJf1tD
Gjh5YN/3jkbCpQvLEBsFEd7n5t4vGjcvzZrJ0xkfYrnyxUKTKL7F4UzjK4Vq
J+kFOCcCyiOQmXhu+KGAwy/7FvEB7V/L69mCUDmG4uBZsvAbNm75pbZg3fU/
4Yn/7CJy22ocBrlq2aTi9ZlbHfrrQ/hByocUwLcQmezz5IWZgQU0CC5Uquot
YYnSLmsgrCHp6k56fg5ZANjKTNEGxlIJUl1m9ZFFlX1ZqvWcGeEGFVEyB2YO
Os7H+gYx/MBkvc/Wky8tIQtxvC8DmwhQGwf9WCBPaCiSCc4o5uBC5feXNCfH
bfai/cjL8Sd8pS1EgpVAdm6r5LpdLWPc//zBQKxQIESIjbKupx8RSDNKS0Nn
e7e5y2JcBiEkSfhGJchuNOLV4g/EF3xW83sl5u8Zojz0pKXn6GRvn3jQ3AfF
DncbTDJZ8oGV8nWeNqFRCAQYpL43fY/Lnxvdrfn/z/F5SPnXBaRAdOMbC5vv
3mSfQCZYD1ryIacoB/vZM8CbpgC1K0UtVWI71RFWuaxJ4biLZ3YSSbW0uLyX
FSGuBlj+5c5eldeMdv/BAUIQoIyVtpFPI3D6/XemLvf4PpqhrTh0pWb3Yjz5
FdZQHMqQvVmUEVzyDHFiU/0PhnKIQf3eBSGavXXwPf1guCUbHH6bl6PwW8TZ
IEOuM5CTgg2Q+93qUVykkjeTT6VBBM+cViQDqm6WSeCyW6Ex3ikQS3KAO8Lv
qbIvNlhg2ZKj0pjE66cv5CW6sFM0FpP1u/Gog02U+Q3wqpMBi+Y1/Krlubrz
7TWKdS2eBhw7ZYrks8pwDxPnI60+6NtI3+b7tgGkBJ2MqMt01CYvCfO5o/1t
kkrp9Fbxvr+QUgKhJaHFRGXz4SfEuD359QdDOKqu+un2dkY9xri9Wjhwv9Fh
OVy0KuEZvtJSKw53Fegqj8hGTLUV1V843r1ZV3S74aXyhyh2mvyzRTuUcj/K
mtegM1J9TELJWnwDZbY3Zu/ajQQBWQY+tXIEKZ1n+trAOE3X+OFZNc8Xi7b8
0c8NFDUps13JH0Fm2dimjHpd/mQCgKju6+I2i9dIZeHYlu9MgE/ahsPnWIS2
DBM4WDjT4Ih+f9tzMfFbCrbqgPjPziIaHAA3NSGW+lq2KgXc+IEs1YMv+HEH
PxJZhwhSAsU9kOsjJnVxq1qfpNlKIYtrGQj0QZQan6WuosgGR9zADCS3tmcc
zXSTlWlT4JuXwl1Ls+DqqQ+2wX93E3YFlsnq0/e3yQ/6uM4fRAi97fmVmKjX
ipi69LZ0xdS5E8FqjK3p0pXbZJwr0+B8ou9YOLg0014NxDQtWQz2n/QCSQvf
Vy5kmGmv+c3w0kFHTfULiQQZu+wahxD1Kb1TvTWvtwYpcxa6p7gABMrBU0Vn
c2hA3sLlmk+5rRwhFVU/t3tTsLixJkw2C7BOtawKp4GPZm3hvQtVMy9SCRZ4
g9Y8qUXoO9fwlsTzkiePrnUlCXY/ZA7HBcZB+II1OhWMkVJs4vGN11nge2Mk
cxZZxkOROpG2QKAbXfAx2viGQa1JC0YDHJqRTV5lO0QqPnfJiBYCgn7fkXx/
osC3cLNjhUT1icheeyu+4V45PZJUzbNR5M/ewsyvbr9auIx8fuF0PBmiTJbJ
v1ejz4JIOijyBaI5K/WnsF5G6k8Il1tQCeFH+OAT46yOFMoASonmv0PrVeOI
YyZRezmSXvo1GlG6G54Gd5uZAT2EZkuWxi/un88of1u27kVenhnjHGlSJxzr
RduiwwfFytwFtlnihWTGhlyxzxqcXRnzowyyHGgkvhzAblxxEI0LXwc96FcS
XT0fr4cxaoZ0Pzzu/0D22zOFr8H7fwySuAcNAail8SgqMJKTpuSflQssHwVC
r7JKCKW7D1VllBAz1wPB8y5tE2F+XOyJH07XV4KNdbceX2DdOnRmeZODesPn
TKO6u05ys6GL/3lfuZvtUuw+7sFc7CMCpr+rW2bUl8qHP6O6TLi6ZkwbK8Cx
LBGAyPnqXBfcQPd6ikviOKgTYIrVzqMmBszwiXVuM/ylIvcbc5eKE/iml7UA
Ii3CC6PqnMLtzW3pkjw1qHc0urfLqv3gAz9Q4sa54alPRjmPDiblE83keldf
oK+j/4NWsvBF9B6mEHJSvIpF1ucK/CG2x8stW3WmTMlMNHkKUUtyGIkUGKuE
c1nQnw/mdjX460o7YL2/HLA5Di/XNNi0Hx6dxA7GPqdmqaa9mT9uSf9Tk4Kr
r+uppPLAJ/5HfDhIxCsNezS6wbU0LqK4SpDBp4mf64S+6jlYM4p+BF6WW/Id
7SRd0vMHlScFB/FF2KnYpArW5BBLX+ZG6cpovBswABENWoniilxfuwwHG0oZ
k3zImPCGsJIVrCtfO5BtgVzdGH019VRaXYcyq6aVsXhNZhAizry7Ww6ENkdc
SWhZ3MrLc+6PezYdAABTCrWWSx5TbyntfKE4qFDC+rHi1u9DJ4Iu7XrLG0pF
Ts+745sG6Kc0M1fnRgeBo3zHalUM84A1576oXiawHHWopBAxxvyt2PCI7jYl
3XvoUun53WJtQA/z36IzlTKlnqNq2vYA4dJaBPXztCX1D0sBjp95p63HW0Pf
LrLMBEZQ7u1pct17KqwyuN5fopOG10P9T78Av+HQgFR6Dhvotr2Cd69t2aM5
RDj5CBgOQX3ryqyqIe//169GnVkaDIlr68xXrI9Ky719f9MKurQD9qEuaaDt
Bbsh6Yhf01ycWqJDenPLR/kw/rh1XErbRO7at2s21HBVHO7vPaKkbs/jLjgo
i/z4oVwFHcHyDHe6JGJj8HJkW5HO35MV8+dp8wK0IHso94hX0pe1Z5QMYiCn
7x5wpMN3zqMxtov6lcxsn6oQ8qacgCCJlUnrTN/g/W+UpjdJGEUvBp3ch0Oa
E/R70kr/KCB0En3L2ZVDDxxnP1G4Qs5dvstU7ByGS45PzYwCq/K7MlNTq3OU
9nhrt9B60VIKVPahr0mWyNE0oT83AO4Ol8Bd9lZ9t5B/scGC7mdP6TRjeELO
WeudUcf4lB6JvfqKIIEwtN8I4bzQpL6KrWqx4y4RRPSaa6prJPGVVDSfDX1p
wVG77XTmrF+Dii7lXftaT1ISmcbuJ6b//Guz2b4ikH3YS8bZt9s0er4cWb7D
kXYKqoW4bRz483+u0UgvngjDEojLKMv1TNhvRjlXWSOsQ3xOahtDR8gpBKuF
6yCLIEOFkCUdETVcGMNTTo0UDr36nIdEi9Dok0VT+GCPXfJQOuhyR6PpWC30
MaIYW5/fmLZI0yRBKYn8fPZWdIhj9RZENZp299AKluTc3qM9f9RR/6Skve9h
dniRRRP6he2ljscWyijFEDTbHM0YfTrSHpVzyXDjB68VnmvQQsPOumZWA9Gv
dMNyzAHFY6jYkOOMJXABnmdA0SXFhgp4zsv50SkmLmkuveFsZ8mADdcYFkmn
u+HjqL6OR3eKj2FBuyRxZUYoTdgkOrU0TR3aBwNEgSp2WnPZuUGqF5MYTiV1
uL6kLmo+MiiE2fYt2mp4vqgkCfk+9QJ29LE/AmoIMUyT7oY+bCbP55cn5qBj
HpRrKcQqqAGMCDprhtiZhtUCMDc5ce4gPV4uyNoVTVhtFod5UuzsSBk00hvj
GHHsuV2xLhf3OpaiaZejRK8SH+L1bkhBhvTLFxOFQdYCQlS09ZgHvAZAqbkx
4eHfQNoaaFR5i1XFm7+faoWCFFeAbZFqO9yXQELd14+M/FjiceXrGSe2786l
Gp0uyPQqtMRYBDOB7s7ysRD8pcOrnTIyY9UFJH6zJLj9EQYMr+WwhmXwk6rV
Xz8sW0ZMkuwbY26NoUu6E6f0DK7yJTONedEcr8qdG1/8PAujOzuHeQux0Frk
2eXuP+FFlEPJX3P/5m/AjJIaT3itrNz9I/7wZbDMBKIm6oiKeZ6fgNpFkoeX
1N/FZwSQu9hMpde6BcqHM1AyfqrQ7oXnjQu0rgBBkJeVwYO+Wyd2ZAETE1zt
r6IkWFE/NA2ZjOlwh34OPyTjG0rhqb6MnQ1bXRyLnReWC39zS2ICzO+5LhQp
xS/S6UGlI+2ysf8Kl4HAOY21y9+R24tG2Re4LwSqmCXlt9MvjmYo80/6qJ/y
/rUqc8Lz4PGwGLvLrozSovMEvdk7/j5Ng0MJITgHL3VXiTjorNs3W2FjjsWl
kUjla8hjwtQVjlyHkVOvz3byJNgJLVKrW8soHyYFSo1NkIaoBINVE9IeVbSC
/vg4+qIUzULRNqFCTKqoV/QFGi7TagoZowK5WATKUa1WGNJViF4APExSwiGj
3us/ldP0F+w6pqjEk6dUW1H8nPIMAZxbRaS+g/0QA2pMxn0AXsjam+DqYNjB
8NsVvmXCL2J6pzFCp3F3TA6y/lDzs5rlfOmwem1FVqb4h3DZePS1zDPnwKu6
nTjR27XbUk19NhxuhDumntWEtF1McbJNEqPcZrH2/eHKy8tDEh7jgG2irTli
iSoAasG31h7ivgkDk98N2La4XR9XSUVZ0UmRXP6g0Ex2kao/fPIIBrFKEtbf
hxhThosOEkLpteN6bDQl5oNLOk8ywWjwMG7SDstEiLrXDANqUUdVCLqqKpYK
/GnIThn/0bqIpySevUQBmpo+znHvPMlmsX4lGHiWjyA2U77MfYWi9IVhzAgl
M/RkFhKs9xSnqQRWIBj0ut1D/jizT02A4mctqM2Fm8FzpWo+U7N/ltRHxMtq
tQABsfkb01Kx7DS9PX5kcRGMWbCexU57SqvNZR2jtb2ipd1EN8Je8dvaOQro
oAa9Ot1b31W8mb565evgU+C/EJOV5BXq/be5aSOhBu8b1HFpEgYuAVgFpXTW
rl1hKdakt0W7S/QZ92ECfyU8bpnEYa1OxLKxDrqKF0ytGwL2xWWQOs6Uapxj
Ws1G30SFqhRtTW3o45MVI9WdFv0tu417q/SDS/4aQkAz5SiHlnIAytcoTk7z
VRAG8x82+01kyEVgy4wDnVtz2jgnx5QBZwkzjmkoL2+rGsEMJBMmUC19s97r
oO3GE58QHNKbnOvUchlgH+B4BIx9RO5nmrM4sgD9I+OJW5CDy05jQE4+Ec5K
1Qj9mu/mtalgFyo9vEfSVWBWPbKPo3FqM0ea5mKuOIktSCb1ZusIA4mg/SXy
D90IIrog3ucrzj+VUkwoHwrcLo5Jg5Wa+iP7MUEhNlsVd06MOMIY37s1Aovm
BjsoxQZmSmWq/8ybPmUqmJgCXsEwlySGeTLR1rwCzBYzRH8Pld4M8OwvYf/Q
qe5+TrSaVo5n1vhyRTIZB64RCrffIjrjHibtI0sHz8nuV9DT5/T8yo1Xe8NT
X32Yr/RBRZQReBCQ+B8gEiEJRxj50Fa5sIQr/wvbsQTwNeT5cu0wwIHuG96t
zp3HJooMq5H+2RjB/q0UYlaxkGoNle7fBmKzLppo4dVu89cZaYDWa46pSBl2
uwdAgbhiCriSs4OLswyFuACtrwfKgLFG7wRi3A9RXilXey95l5cmJidAeQNw
iVHufpTr6dfr/YTpRV+c8triDvQk2BUxrG2Q9IZW7j5Knrw2dUNsAJnEIrDn
+1zxj3iTE1A7oRg1Ps593k8oFYKjAGGGDbEzn32BmuhH7f5Ge4mm19HLtegL
yGpEkZqiBRJtP+5FIrG/fIO3jp3/dR/eNOrNTL+5fG1R0OkDllEG2P+Z3F6G
Hv/NW7DZ8cv7zE93XGFTiGmncCDW1khisJZIHRKTMmUGP6HSoB3qye0cXQ6B
QPPuN7NNMEIC92v0DnZcCuamgslViSNDdeO4mXZ9vifwgQhIk6X46TUtujpI
WY52rad/1d7jv0PRLiHiRUIHdWY+BbfsZYPbUMQya6PacQLPe1qHNjPdzWH5
K2DqdvbpJq3j1dreWXMVe/7is5yFMuztB9Rco+AePG7Cg9w0EedI8CpJ2v13
+3RLRuYr5IzbMAiK3wDf2WJk/yC0WijvX7nz5PsveEykC9SGFeUlzfyto5lc
I45S/QWVfbYUpLvORKE2ttN1BlqiNB+UD3AxFAV4ddXP9llWORVCVrc2ScEG
P9FqZ7fKot8i+UZJtlpVFlfRoT1+NHYCEWSMpkYrx7MeIL/9S/1LPr/A3tyx
WfuMLF9070nsAyZSm0XABXhoBTrwpxbmGeKezm84wPe252R+MzcDkreBZR4B
yurUu0XcC3W2IlQ93XwGz1cbCHnhOwpIA6qNWeJqY8f5aet3j9yqiFEXNcY6
+dJje+89vS6duKxHl9q0QnMgHg9ARO0YWEja/Jfc+4l1ZW92r2LkrBRgqpZM
YcPuB1p/fFIYb2CsA5rwEeZ1ToWd0eI1cPVGfI7QVFqtlh8fifxlNwib4270
4ViaSmHYbGZsrUfgg6a1zZtntavLfnMU9pkh6iWLFvTRFz23/1u8SpHY64lm
Rcz+OOHgbxaKAfHjXvd7nTMvEWO9mkDkaHNYMcFOklk4JTd3vMke7+WbzPhw
n73n0fgBPBEj0sJK4wqcmWUqFpq6Go4bwbQo5tugMO1m7frgbcttOvTtPKbm
a0tyIX6l0SbZ9IQYg7W1ksx1tyL+hZw8225SX+eDEywCYJSDPKdiU86yWqHY
ZNhJ8kd8mpVLxUdBiGABonRzT0ZkN9YDcqVivPY4gajEe/Y0+jXv1ZqgehIj
Xp5vBdeZORQPKny+NZBmg9Z0fcxQm0hKdjF6NQ/1jfZSxZHPBdDafFHr2Ius
j1zuUJaeU1gyZQLRntakezsu8NGk+FTWIyoVZxpa4J+cQyssa0pxl+40aQhq
wKFEJltiIPzP2jmyrz9/U/jN4MBnk9QFgkEsnjWzJpBG+wJtWvcOB/nwD+ip
ix9Q07VZx3LGq4Xga780H5ln9MzpM3MXLJvrdIN2CfNwHYhSBS8DkSQA7rDO
1cthjj11AGzlbx24QIQg/b8k3vfudmaOJpkt1Tjhv20o+WzcM9y92CPbCix8
HIVqE1TpV+9ddRMsqVLOa7q1Nib0CNeVsZicDgItuEZlcL7MExq3dgcysylY
r0JszuebKH1syy2eM3hIudkyRS6kwTTMwZSwMrKkvbO6AIEFxPRJWzFBENQC
VTCbdCbcMLomtqm14vuECbm2XnaINWT5gK1bssrI4iAvHe6xXotFTxmHcJrv
eFiqLdYDcd9+rpGb59vzKjaEJrFhrDa0/fnoRg6m71uPqaBM3qcEkDS68E0s
JpMKU5krn3K3mUirK1GzhnvBep22VxaFN+KSSeW7FDfNJwYer9EgLp2Z9cw6
NzINLCBDD6OeNsmDDhMpEYkYGmdqXfrLNNF+wSv0eYnof9iW5WJXxzQYdQ4/
Sg287lxdJXhuny7GvrMcOyPeUz/sYJkcPolNB0HZ58F81hqrAYyX4wAWYlNj
RqNvW2ApvonxhoPTQFtQiC7lvtqBTvSNxQ/TEtECPb464iIf8hcAy56WLQxK
mw+ozk7Wy0qoymL7ZwxJidnGLQXqVrdyo4IbcpewgD+nBV+sZJNX7CvFCbHk
q3gy3RL9mvuK7+QjMe3+mU6Ejkx8iqAb40ffgQBHsC1X8JEFdyWN5BujWhgH
Jjx2VmmH7hkhKroAgAvLF/MvSG5RAuWF9MYr7zR6YjtLQ1sT6lO8Ga0wt6L2
azjDKWXUrMJe2YY6I/x7KNUwHCiw4xuW7T5HkxC+QMH0IU8gxTnC3eXfRAD8
0N0IZelhaFnhUhjmwhPVOOBQdOskYRutgVE/81P3eaqK9EMxRdTs6DPg6dc3
0XlH0Y04JMIFhbZ5XyKECU4yEuZmnual47nQ4bzmCpAB8891FcyZ9TJtgkd4
UL4GELaBxr/im+YyDh554pmH0IVorQBDsTiAefXIjlN4AGfMJLX8FIfCsF+/
TsiU4OYIyQv1994p9E8OdrBDBULKId26qXgI+30sMDdg1cASyeio1KYi4/st
Byx17rtdLBn2VYKHY/FQJAfDF7NXx4/69MnyWSOLHh6HfwHZp+q4MRobAb4u
RT6WB5M/6n79KYlN8H8S0+QkqMXUxzJYFV7AvSoWmePHibTI3I8MDYSwc7Lv
apN965G5o2OejIDu28EpQZFdxLRwuMhDLc0t7UGzX8ugakPp/FBEf2tTMeqD
MrxMQYr/JD9axIQQwhAO08PNsb1aRU8i2GktAyZ+syRNnWBDClTnamurXexG
Gqo48Y5OAWhNmzT6mTLeXhpRcFE+ynjH7cl4nt+f17I59N1m+9Woieu2oDjd
/RJusKuks5yQII01bHyrRfxyqgSLhJQt0i/8EMeoczw44bAyCF8hKTqaO5FU
i2umJc/7OIsodSeKU1SofmP+3ANHoHfGgteww+4DlrxgcNKf7md03vZz8sFt
Yq7wBMeovVVgRrYKp+nKCFYEtmQ6deIY/ZUYjPjvpQjoackndSbVYw1DvOq6
lyrEvMpQEdDzoZqDoVLG+Ff1QK4dOj+tPRAbPUQziMcBvLCWUgvY20HVNmHE
a4bb74i3cRbu/oH4jNiHQZ6EEaPewHAdTVK86H0Y4e3a72qLZ+kbL+n9s9s3
fovQ66YcR0lBU8PnPloOuMc5CSgRwr3XwwSrLiZ8IUUyxhWMAnIZEhMkYOrR
mW0Cu2GVjrIH24Ly6SHkb3zYHntLo58WIpjOpWNNUPAn4fI0MmJ6S+MyBamc
uKwWX0Zlbhb7Z2ItKDnMpf9ixO6w/LvXQAifIaqzRDj9aJXTXgwVdA6fT1KO
nZQUvay3n0yfHLF9wpdrewQ0iS8RLF7o9kuGPGW1M1oxBrKeOF0Lg8ImBajy
je8BvFb44PtbS+/Ly6DTBJMwRMZJf1P8b+bR3zkkhVjU7l7tMdjgpjxt3SV5
v7vVarFpBnmhYWu0Xm6Q+UtA/OQtL79zTl/zHWdV/lJusvwFBsfl9/5+ulxQ
hJSOjnFc/DvPRvMrTw4bQopA85gRwG1M70ioHz6qfU1ajdJjjDC3/J76CDTY
ShMI1eg8IAjhoOpbZmLdi6JRKlNYayBga/4a5t64QPvPp3N8P8Tr7Jun7bbe
on3UXhJEbeVwRlKNK8coOtRAyqYmtiF5HCpsKHthepOLCOxGoYZtXT6uM/t6
b0DgqKsSMW/V1Tf/DEbZgWEhit1STXG2jLYCt+a2WZolsyTsmRObMgl8DUBU
LG1OjyfVLUqMzbbw38PjjaAu3msb8xlkE7wJKR8m8hYzzL1V3TnEQKov4HrM
C21yIy0Ufh6Unb9XQAOD6cH6elTlcmK9kooeD4QhdW4g69+UB81Ic1Kzlkxh
qhtL+Tf/pPhNH/JG9nhejixoT0xwsRB18j9MxPAHsFJkKX5auk+T23dh2S1k
azvC1saOe0pAbquTeZ7TNf3GdVX4yKiUBIlyhgvJKJV/NzRy0TzKjViGQn5m
88QKdgO7nNOyRcsPyDIqVUyFnI9oDnZp8QEa4YB/RlM/apSMNnoz7Iv5jJTK
N1t0t+xgA8Rh4fRdP0j/bpzQDe0tKcxRKXdTv0ogUWjGsqwHzxVFZ6Hu3cxM
74co43QJ2ehfZ8GRgyxHHcOrnEyzNeUK5j82Dmo03G1FeMNTaZp3I/x3Ey3a
4bFYQvRaLrJwLispLM+HysZSs/lTZoovnsujTOvl/fE5f0alHp//Uq9JraBd
L3CJrjIaso/b2PzT9MSh1cKSYBBDLt6t2qtUVc7SaGpy48kg3rgMsPezpgbN
ZJNeozJQNs8VSy/gKkld7o7IxfZzfwqwfAxbHS3do7gEHmBC9ErM21OU9ZhQ
x72/sxlp2WV6gOCxb+/YrOeBPpfcJAEdjffC/0brq9exl4yfdUPKb5Nur02V
YXbIDUpK9kiberbsg2si3twdCnZl1GpM1KkcWH5KqE+QyyGjBFcjaYzvH1Ql
Kxf+rz44KRasrTNFN07nYMKh+yphz8C9fkcvzjVW8e3rSGXzme1dw0FAfgMl
/JOT3tkLOp911uS7jV1XoHATrayR2CP5OFfdP7C9aAspnDgbmRjLOFKHKVk5
wR9LmyhLUs9aF2o0sLg89tTz/vxxe/17E8kApALgKJLTar9O77RhYlGtzDrB
xD9tqFpuyKh/6uLPGpI7YOf6FF6QnCVPpejYPnG5jbpQbtervdrIiD5s0rps
Y4RxDSwDC211HsFkwG6vpheaTkuvLH56hKD0YQtghSqf8MF+rLUKotU9z+Qp
fpl/aQ3eVgVgy9eXjgWRDoiL0mQ3aJ58nX3iEtL0D0oTUcBb779V2juZERn1
zeTmHOvpv5PmYdAtnEhAyZ5ZbashNHYt5VwUFwixlh9cW3WOlcWbNCYTLqWD
TeqmSo65JEIyv+X5yQWDa4+ZyJGqsV32KSlVwWluvAX/eUikV8NRIIbEgoiz
n3lZP/MEXC3apdkq8/ZS2pjPrv6hjhmzeCRJCPBZxKkYetPlSf7+lNQm6QjR
L47LrJj01OIIxchj2iagtwxyXNXG7ceRZDKHz3ywLw4PntWS0elEoQlozjUc
pLK8Kr82HMmKHHhH9b36PHEoGGEzKIvxxmJakLG//ZmLyoI4XwTGhK5ifGjm
qK4S4cqhKXtbNG98GPJChklEvi/Q9LD9L9m3MfVag1QX44Qu+PQ7sV3lR6Tk
/jnF0/MCd5Tk3HttPf2ChLmn/w4YNAutNE6rJSlOJBtWIrKng8+u+neGnB4Q
4C/be4D+iPfgp2Bdidg6VsxbXndHOy0t8fI/wK7mUFxq5lSo+ZJFdDa7WDUG
3v+E4gpQYkTIPf9+rEIgLFbnwK5rfU7OQwF55LS5fAV+1n6NuJbnRaJUBuq0
OpCF6hbS65AzDd5SzyW66HPDNL0M9IkKRThBW90S9Q2xHDsZOboS2t9pEqjr
aX5fgehTJAHB8RnFM4HWYcHMqySklIdpVoloBbGoWoXPslz0uy5HAxCvn9jK
7ZGYC+FZlSD/jCno/eY4BIabMxAW9ZC9K6pYltmRSvDOMZL7TrRIay/QN604
VqZyXnXtNWl5MvOub6AsQxgNxJexK9bgyxK930maeK/N2b2aEebT1o5RqmAA
ROy1JVdW+L1xFoAe7yrzdygG/KFBarNCAVAnnEbyo9JMGD0/zcAOv+7GASrI
7P39oNkB15U75XOh7NlIRgJR9lxZc/qDmZIDK7W5THqBnVxN2bNwgZbmw8X3
Kw5T0KzPgXms+V3IH0t+74X+xXcemqw4qceINHuPk00uEr81w3SCzPQWIhdc
fCe+FP9bIkmJVEx6DLPzcE3G/IKRATJQyFlv2yK/oPxwxWCahlU9Zez5/F0M
fZe8accDnprTfzlj94OhcIsSdhTJV4An/LzJwUblNaq+6zbUCW5qbU250tKY
gHGoX/2gQbCW//sx5HnfXZo5A8tex2WbqQn0TE9XpFHOqpwR0KfgUInVjRsm
ipuXM1hGy7NK2h1LY4qcun30cYyXqzCW0a0YCJTM1R8XCW9sloIQalCRGv6T
uBX9hMcBT7AKiquI8a7eEXwnrej6LXv4gyL54mZOxObSM7J6v/F2ETQEE1P9
DyE6SwcrjomaxpX7l2vPMzBR6pu5SaWhQwL+pgESNUCD46PwymYWgTFfZmDt
uieAdLNY3zucW0UT7eYymtnarXwdft7oUf27TCLvOcBKiL4qDgn3cgPwwjs3
TL0IdCty7RkJ81qjlI4b0eVVO1L9l6Ko4p0oiqfvrNvOSVHMbDVWJWxcolgF
DPl9sytczaDqrCz6yoLmN5pD417p2gCR3BfjwDDyL2zn6qdUrDzP8w/bMeMy
gMrF/U76MDlMB/diatSb4S8CwRtCQpr3ek5NlPtCknd3ykG0+xBDh7VKcgeZ
h9xMaz7hVJcpSksfltDeksiK2EYT/7eUHe6Hk4qGzcWVm3q4b/PCRkQKgFYA
L9bLgz8WbFsWoQlVcBQ3ao3XQkG43NYAlCQGfPVOjCGd9Lf8pZmSgKyIEnn7
ABOd4zwV5DutElIdS8TMQMjhuBDaOfHIQL0k9jGu6KT6LeP3ShFfCLgxrsPh
uRDd++VVj75GA8oMhPqUuhcLw0sJjzV0/BnaDk29BNpSSf+lUsltD/zLQBTs
Q3koDyrErWLspgEjQFmm8TgAk1Ojy0mzJUUJOuLGzwGRV73+v4ytZHhphznr
4SrShtuaXB4sJdKgMVnPg7iPhD9d3B5ETOlUMe8QsZ92s89iLWfnZ79eLxaL
v09hfWlGawNZ/Qy3WMTEM+iOR42UiKRp1zHHWLwkhj9iWO78dWufT8xqqmTy
dG6skTStqJH/4vkwsRyweipUF0DlAcVutOlpCDHH987wEaTUopOBPTcGvwZ/
xFHucTAA3nVFT/RkV1/kznAfdmalRJRl1JKY4AZiS+iYoOmzEUT7L7liSyXg
4vJiQ/2fnJU75JZ/DLgHaB+a0D2GndlZ8sr0kPcR9PRpMd9aKgI4P2QfEjiO
PS4zyN539ZZ60DlwnU5n/xju4l79y8Szx62sAVKUXJQ0Cx8pB2+ofScuadWk
rD0C/5Yf04vAJxFQ1c90NNGWeAWxbBpqbdRnIkGkks/xD7s+h43kJa5sK4RU
xkqw5vlLIs+R3YE+RlQ9PN7DYmvk+/pRQ0vofY127FpgR/XtIamRwZC7lMbO
C+rdNb1IrQJgtU+Mll1ySHS/s0Yd3nawSxag3ldMyl1sNZBK4Juid1HgleIt
Ev2RVJlmpqh5HCYmZCouO/3RjdKODthRMl36c6t8g76MjmsCv2JJx4Qcck/m
HjMqtdFcMRD5uprt0bhXF3ob3PEoststWgViGEhnR2pAF7Dpe+tvA2Jr0rKW
BJDGb57v5A5j+4NHVI7wPIWlXNGLkuL24qCQfqhipMKZ2obkE9i9FUcZkyYD
S6ghsCc23efJxxZ+aeab/FPL9tVeolOfUE6lUCJDCJKPJlAd/X8uz1C1Fl9h
TgRmNLLef+lCiCrDOI5M35ki34HVyJZCn6EF7MSwDoz2jOuQ+RlbHQ4lzAon
SHtHij1LEFtD/p77OempfFmomiNm9rbjZnYrr7O6XxPcxKrS+t8IPB1hpivg
I7kTOcxX6X7PZnBuAfpW3cAr7dPl9SVC5NEHUxJLGODxqqcGBpYDFv5tEVxW
idR0nJmnJyyisVv8JWF5dOERKJfjQ3BX7IpkiTXAe1xTPFGTZZqMI/SV4ppD
9t/Ds5P3vopISOBlmcFD2DZAaS1gMp0NH+QqqbB4Cpe/IG9q/EuKrALHv6zM
wakZLOpiGlqFjLrzib2l/ReXn54Fc9yWvPUCxIDnmrtFDTyr0weaXYyW6BCZ
Ec4MJWjFYzJZwZGbbMi0+MkWT0FKoMvfTKeaYdkT/uYoRp2XnnaM7wAr2XpE
2kszMm3MsZUz51eo7gc2OE8PG7tWZxnCvtZvLWSvbI/EiCtypWspAPsZ8Owb
KC7wQC9wsNzlbLOaSvJxRKVLFpy3IvwoMPgEO6YzEmOSlOV2cs+oMN4Tf1kY
QbT3Sla8x5D1Za10e0D9sPG72C9JQR2AXke45j/tAEW7QWsT1AVNkwkpIWiK
7J9DBHI8rTnhS9KTOS+03FwJrg4BtsxBsnSd0e+dQFSsEf2MB1hHiudFjENH
dTPsBn4sVKP+7qmFjtdxEWh4VCtWUVuqUeQv+wRdn+WgJyMcK98oZYgKhlH3
LOwONDBbE4sbpYrnJrZbyI/Y9XdxATmegRgSjGPMKJBgG4eX4pUOaIpkz9E5
XvNttVCRmL97NDvSiIrYmSIy4yuiJKVNr/QuyPeWv4c+9tUSgk6nyYTjv8Tb
FUGDZuexJ8oTnEF8w1Wkr7KN/gDuCsSxxcvf6Td+m05fJN2YfuQ3SXCJfFlz
k83hrNw2fzXuWuuGxf8DC5w9yY0Ts8D2j4dOKLr1td+ovLOC1b5hp1x2fruk
SdoiLaQjoKzAu4kmL1wy1xL/3eEejuNwbwD1zeegGRk9wApe0l9LZgAXo69m
C3464503Yv00T8zRxYJlbgnW/FiLky7KqojJIJRRNweIdB6oXQHRnP0WbuZV
pQsOCBKWBQGWdDtY6TQuHLspp04mMTQNoeW+5Sxht5EAHbZcF/r74J8qqpQu
rzlG/DcvNWG5nqOe9hI2atQDVnyuiy+cpQjcSs5sOavRBLpB2JHE7/daBA4k
4EaLcAH5eey5dIxemq3ZiXyPv47vu+I8Doi2mQuhq+t18D2Bex0j+GyLlYUo
NCpyQsrvhyDUxX3GwtbUjqWAkJhef57+uX3oqg1+Al5Qi394Ip40arkyswjp
uMO64+jnniwNvTnQui9ngzHk1OxdyNS9gdX+luxmUBDGHLrzClpNdw6v0MNs
gQlU2bpyy/mfq1LK0UW4SqgpSVz/73aKA7xVitz/yowlsbbmNeJq4oK2rCSY
xt++iuCkkTGgeJg7Aro42WXXckCvmJtB5wOrmifZfri8allboOBYrnWqLUv4
OgITuZo03xCS0cFFcAQdqNYKisXmeDjhU5AabSef/8mOS0o0D7qs/SoOouP7
oKCnLxjq2daXCdWB6BJUNhxf+j21WA9qs1tlUSDVJnsdcIwhoQRV5yPDwVyL
rH1Fqfr8j8PQZ86VATKwCM/QoIlZ5uqWODTKsiUbP49NjlREuioeJhoDyxuX
srS5s8yhJ1wYhybZneUfAvMdsdp8m9jJXia/kKRLgAtUnFeemBhHj5pBFuSs
IUP/WkyhrdyzUSFWrnZ4ddvw6ct3qmwuFWKgwo1Epc4Wdeb3GCzPffTa8idq
08FChyiu59bwxxER2PqETsNmfaJDB/oALuIjXKsGv12zClv59ZukqTZNQtX3
XJLnnqFdELgJpk9SIUj1pdOzA5++t1aYhMkElBiMm7KiXTNQHoZSFtgoBMXm
AL/tjQS/FJUf7IA17iLCnWrtYNghDCwx0wjsObOPTtd7zWcCgR2Sq1XzgSpK
B0PTwavMfcZW5za+UCwtSO8qKivgd1orPHGVRDas9fGUw/hfh7hxIG4OF0bf
5MRVKotJr8E2/+B+f6ktNJZP/2NaTTw5f3/rQMvD1SUNlQpwdCvHBRs81ilp
UCQ5aeVB13Zxs7k+g1Myi+MJFrRUGUsCCQGq/fuDAtF1UX2lb5bzS8LNNVsd
9i+bYcj7Voy3JMtTQhC76B/r/3++T/Oizu6X4oLgZLvnf5gqTTV9/fC22361
LKnOT3MnhBsvPPr5pV3gPDeOSjq9VaLumY2jXZynh+Qe5MxsqjIsPJLYreqW
/MLJjJnDgjul/aHWkpXS8iE8FkCZOuToIQCHnAIl27XzcCQs+Da18fEiyG0j
zsrkLXD/P9lOdje7xKZl1w8PvShup+jK3AdpTmboGMkeckzQp8TncViuztt+
K2Cl+RKfigjBcFp4BU7nZrFZl2cVQ7BRWOI9izLajUUe6irFaFDbmcEeyQ0B
JHjMUERu4hLg4l0LDw1bgbPiwRpoeIqPitcn84rmjRIb4HU8+IvYr+yrOR3n
up/2yJQ/dAZQ82vLVA5nlggQ0hvM9mtvhKLrWPr5CszAV+urkSQNzuVJNSxj
bLicNNEd2Hj9C0acciUP+v7dmS1pIUeAjYtSaxKIjb/G9AggZ05PYeVuAbyN
8eJyY3YtKsqAKwkIGP/zVT6b0B7NE+ejJGeg3NPJGk807fWzAmNPXOCDfQ7Z
7oSVtFjrVkwtzAHjYYWt3cMbT9mwRbVP6f0GH5v9AfdSMTgyqbNLhKfTi7o4
76dxBKXZo/vP2uRyIHQgqj4Z9HqVEcXhCqnkCFzbnFZy84Bq2nh7fRl2Yk4x
IwLtQ4XCRC9anfnzklgACRMHOSHeU2qtq9kMlZg7PRdMkWS1GQeAvqOBYImY
auxkCL4e+jlyiGPR1+rILmG8MgwmYmhK3lvPyWPvZIxrG2Jr9ZIwEzTaNb/3
5n4y5kT3rZZvLt04JTGmD9xIJi//ju0S7bL57ame4cUzSd4E/GDaNdWlThlc
1Lhd9F647XFSeSqanYC9rqYzsDwLQ12c9kXkI9LpypqcrD+6abMp8pCr0oiI
cbBe8HMp+xdPL39lFPZdbOwXQyZFdyK6+gXgZencVb8KlDgr2jEHrWirkYTO
kuOvY2++fBkaFAbyYJKY6EKTbbyzrQgEzk9LBh5xu4lMnkgqTULkctMPrQfW
bQjI9y1oq5SN2O8dYBCvAH9V2Z2yejUlxgctUyreGQViD6kDQtCZ6zM1kmBh
eOx6nYUC+RB8k+irsWDvRFvIWxMYDXrY0VAPtZg+r8tyTykxEVoJ2E38Us3q
ZyJwWg6mKfbKX2bk5LT87eGNnyibFqFpqKRv8ZKdQHBprfY67QfRqjxw67oW
ueD6qtNAsxMnEjwYpe9rMwYsEcMPuMBF6KJOlEGywwf4Th59qGFbQ5S0qGHi
K/N/h7JSriK+urbYfGD+Oi1GB2NbqcDnz+hrJRQCV+VlHgcjorCAnjUzDuP2
ANoP4Qw/6nVGvJkI4Dn8FrrtOxZFLoNMFcP4/dX0RM/UwGlpawNLq+HOePU8
cgoszQzcXHtCzDflzACwGMtawm61j2FL8XnRhKEaoDNrlDKmRA7HQY+aCFP4
zUg7VMj+OpoCaCNuknNbCCYAnZl07QUd5vhuLNjmv7e/9UxLbl4aOKBtJTed
Joht7RS5KxDBRVntlL5Mi4jWuOdBr2ZX6ZY/otht9n0lJI2dyWP6iJC7SrKV
70ts02xd5cQAJC44yxlipYiZ2SpOjZ9KDElSaPcyfpfnmoLyNt6WqJ5288yG
HPIRi1MHmCXj2U1IIM4y6d/CBUtswwbvZUT5Cr1vrnkC9FWmOsG2PSauayuu
IfB5XAOBrDh0bx7sBWmJyetHGIEkCCHCO6qZI4lN8LV3gWU2NFh2a+PX/RiS
4Y/bleaIYVq6QpxY6T3Yv14I63i0q93FhETp0YdAtVU5Nce2+fqCz5A7Pkno
WsYJcdea3uxnGNhNhkfBgFqxbXFNzr5hBUiJDCI3A03PRsiItteUIUuLpccw
h5IAIEmJSI98CbjHGWishyR/hAylH6/antzJBpQDeE7xS2MTolzH7ZhsfkK7
Dc+x/Qih740yjA8OgWcoZIbmQOFe89rPnqShQApxbOTRHk8zOyTU5vQ2ikud
HLdxq/ZiZRw8gnlkmehV6x0ab4Bk+ed5ELjFge82NeHHQfncGVpQ8lTTfLCu
o8ol8mnW8Q5lpl7DDk4P0hTzXl1ZK2ln/5gScC8/DMnIKxB1V4MB6hBTbLkR
6qkypK8znZ1LzNYQrzcqkXEn5OllMdG8COGPY9FYcePvD9HrqRDigPfiC9lX
bQMueJiBoVNq7TttSnXmh7QF0uWVSgptcI3jA0OyBiilPtV7pxTAi3+xIslS
3OMGRGihcaLhmRVfFTEixeQHZMAEVAx8QgTu4khyRluzLba7nfYqnGDjZfpK
WGs37Yxz6EKVTeg+MkOZndkvPLPisyT+yH3Y6Kgu7uMWW4vRzFOOEHBsZQ4x
MTctDtZjJ5YXXXeFMT8EnlDCnF4OjhJkngepMtSWBDCD7WEIzylg/1IPJFMI
qF9x6uGg4dkDYK8ma60nHGhjsWEmxENX7Q7FH3gUEe+vMD2ijpm2GhJ/vA0U
uJq57xhKDAi2/xhrTi+aU2t5/nAlN8nC6Vn9Zb78Z6Oe05gqEUpHI1aM0u4v
Vp4iSWbyo6Yi+3FK8ER+0jskolruiuKyR/3zVFhzMjXcGm6o85xa/a3Ka/vp
Uox0BNMZd8toBbbUU8TYIxFjwfmoYfpvvWe6n23LSZXzAcd7zxai3dNlKUcW
Mdf/dTLtqx5dyZf/aABcWZEyOJhLWLFrSBN48ocvsKUVHqRkBDMCpySVTMt1
4svceCcqhFLuTKd5I3DjfLMoAtmiHJC6uVswmFkhLooMQ5gRCrACMsKlCx22
f3oAp/04s0TWpUPfZmbTFHMnSmQn7DKWkHqgCxPnouR34nolxAUwlBOtlHpC
BWxHQ0LWkrx0eLYfXSu9UzKRgDLrmTAoW78nG9GT+oIQlVrNfLEZ/KgV1o0u
H41HJ2M8z2Ny08XYG/lOMRk20e5KYZkpgBOVdh+j68KOqAAgfwsc19F/w2+D
jIQlnfrkfU7oj64Vmn3sXbc0LupbEAUwN5wkfgZ1khFuKukqPDDW8SYPBcJ1
wG1vwptYznVdQOaEy3LgXHDQyilDOZtRZJDpA2tUJD3IzE2k+vIxRy4mib1y
w9uHOMZ9CXllvt9d8LOlShZOmFmVq9Drn0TCfCBzYsnRhJFJ0ASBSM21ya0m
IkG2FeYUcEW88ePi8JHDAecbmf3JHfPSi5eUA9795hsCVebCwrfEVjX6sv28
dxx7HtneDIR/25EWmDyTPtmhGax7iR0I/DB/cFk9M4t2IOo6Xv6zPXvGXSQs
7ClZctHAt6DE/qjei/wfQ8j06yNPqCdL1lLbZcMbWzuiWV/G500EPtMoE8GM
bTk19F43/AYOv1ga8CLa0i1OAWJVh/5Jic0mJ+RZPYgeOrCx6KyJiuMkI+/4
Iwe7R5dSKYEnMgObvt+EFykU7uHkaTkBnEbYCjM0Xz7ns+LiEt62pksyDnas
qZle/q57KU5eZYJkdR7D9rBwjQRpIz8Q2UaqslcgSyMmTlAQtWAiKc5Z/Z7E
5K4JoqwiBXTxt22Bjj+mltXleZjTP/qQSxW0ltY3E6l+OEEOGU619NFi0Rx5
3INoMzl4WYOcWwNedS4zUyjdg6bqkLoLmULoxJZxHSYk5m91UCLB6ucqwn8X
QgIvt+P9vlDStdQ+sn6UpDYfZcFGXkE78s8JXrArQkyuNzjjm0CjczMMKfO0
SAA8V61e/QeE9sBMiFR3pgcB2tRjrwVduN9yb1YrOIEE94pEFne4kvh8YU8R
Gh6ckW2lgOcagUzO5kBM5mEfpQE/LJpN6g/Levy9zqBPAt0BCecXW493yrgQ
PQXyVB7HUYN/wU5zaiYYe34dZxdi3yckEJda3O2iGkiBssbw4+lUViFt1mX2
E7LynHpfjjDiSwuJY9tNTrlsInJgcsKLarnQiYupfBPqRLHVcFC9JLHO1eXz
45IJ0c+SpgeYnrFo8DXKASbDItLKF0ttV7hyzsiW4cAyqq3+YFhot1GK5vG1
wU4LYVJPWi+CapSL/HhqHLcNBiIzANX2EDTSSfA40rfgVMWlfi7E9ps7v7YY
lvWCHkiKH+5YZbTl30b/FhkXplKh6uXko8xDK7Eud3SUcorhXFm1uEpFJlns
Q0JRNhK2kXd4AhOOsk3RVvu0GVf7nbJy2Vpbls/N4dU3orWB35/Zmch5gAy7
SYhtoIjMWSnwS5KcTN2pA9bVc5KhdUUz4jhSxAsjksv9/pqerqyX7DcB6NnX
Eq3ic+z8O45liJlQPhPkWbh/lQEOo1OhSXWtQBYzPBETXoO2wTT+RIaFnC8y
c79jFMiF2qcrlt7EyafWoHvQ8MCl7W6vi8wXPbRjnGX2tYU82iLLov2NE9dI
b0NYBD210ez7ZtCZfBNJ7vDXvakFiqOYQDiYLa8X4BOF+MtH/Qrg1+zhLUM3
uljlCEd9Q+mzUMA72KO/werVIKHgAojWSsv5vMWNrVguG8JqboANCVkxVtzG
2F9XZHfwJCJErBcQNBGder3pPAwDm3VjaG8ym05Y7wYAsmUVQPTZGNDgkNsH
s4kRim8qYew4OZHSku4aYY6gJ8NsB9pYvqs6clge7xOmN5CY+nZMS5q5E2Ai
mZ1wA/w3Tn1ALo+e/vhoctL391DYnfVKBJFP6sfs9XzN8W3cYy73m8/gFmlV
9rtTRPdjUSyz82/EpzGOvCGTJOv8S60MGBCMiH+PTR657EBjFYZwOZgwWrwd
Fyzi3ncg3ZV1HjENgHd19zxYSZkKZME+1oLMUrxr1FrbsACaEPO8wjVnMGnR
iHyMhZloEz5IV9JeUGIPQqdUFlKcSbhk/4dvRAjGCcLLDiwRhUq1y4duibk3
tHI/ePBLlpzp8fMbuJkbZh/z9X3ACqTF2cLLSpJFZdQimTo6wlMOzCKOBHr3
WUbCiIYEneny/YKFuiISmiMYc8TwreJxDbKld7J/SN7yao9WlieIXlp7qkGG
+sb94Rjf/4EaS6yu/BjMYrxCr4lkOi3AlURWHchqwtrHuUWQpklM3UTS7gaA
XRaofhWYqjl8KInTlW8yJybhQhIFKjHZXo/OY+vDLZSRHNBQZ78rHBEqc6g8
my7Ry0S+F20U9Twy7WO3lrdgtiyUgYVeazHTbKCF9shoHFSdN8Lskuzt5nMw
6tbJ+o2I1Gy4NEmR6fe7IkfT2X3RMEY7P7br9kxgDs4y+0slLDJFbPquFfJh
9QwW4N7Yl+li7QMKp+E85nZCfqy8UjJ4m+SOG0H4wVJguLGTLXVXG2aBHH8X
Fin7oDb7zyyKB269sJqoGJLv8t2kqUnzSMYLGAe6NuOAf055cZdsOWwQte6p
QXay3YGLS6aw7YiGuDteeSnw0mBaUyFencV1XQV2JTdG9aZshfvS3w95VS0e
DATys76PHnVXV+sFDD1lZXevIySDRsom0Ho2LpqtNrS69VhyB6+POzsYQhvG
RxJOC48z6e5CrvdlrKbb9LdKpFIPM+E+/uhy0+WaAfvQ6DymnSBmTDj8Tewn
KDYEg4B1KkxplDObt8uhaTUAmsCNSJFD/Vk8UCOlJvnuWAYxuS68YAgKzdCS
o+qLEGBJ6GazRD25APWGesLri1yPj7uBxkaSoHOia6k9aIUwYh4IRaGIHMIp
3mVlfDhkBw6BNsp3A1AE7GO4XSDp8DagF+wiqGznki9+mcwQtpIXWKfUCUyq
h84xdvOHNRH1olqJwypP80x/KjLWf8dlCJBnqQDPTTHzSTLxMyaUEB7h8Rgm
XvBCBO2AY1gUxl5CMpiccrA2IxGM8NlaSGy8/p1iy7LeFx3HlRuOIsSPd66R
4ZfP4wDfAb1ygnolmZ1DXAIDIvt1Jj3Ej1P4aJ2krUHU7RKvD/GwqDy9gP0k
DHh6mt8rMv0EqWhAHXq3ZArbXGbQXWifpGLNDqAWCI52PHfdQiGg7q3RDs3X
pHWCp/ABt8nUkMTdY+ufKcgg5/EcpSGtEHLv69pgMpa5v6qC4sl11Voftl7j
EXwKkqDF0q/hZ/UFeQy1U+os7cWLfZiAa5BpFxVCgy4N5ROcMOL/QJ4umqSq
LF4nnSHTvhm5Ws0a+nwgCJFvYDSRTTusYog7Of9xljTwV//h6Pcibv9B5tkQ
6I7rUAUoxyt+IxVnTn/U1TVz4mAeL63lZrSZJksrG7BHB2vVphAbkF5t0Dgy
4GezOQ/3dwLPjLD1Y8M7MpgyFGzrEvOb9H0jUAoKpxG7OlyK5H513QOwQYzf
1DF+8pvlKew8H8a39sGMrGVKdAJ4R3aMqTgBbm0PKeMuuEBl/KgZoipGxdrM
u5Db8amntw16XkT1R9OodZJFDAiS76ympieW/6YEi5A8AfSeM69I3osB/oL8
qstBKF5XKqsDtpO6tXp7xKhcUKczSu5Rsio5br0LuAYRRFLDnuNHeut3/EWq
EG1fs3NEJrskgRtcs4H2J8bYgL7xu89TTtxnPVuqqLsRWHEKc467Drfaiuc7
eDkqP8bjk6F3PgOmvnErFGdW93kS1s1qGN3XyuXRn5ZMHK1MPvdNCgUmf3s9
GMrTk+RjfOl5XyKkzWQgz2Z6aN7iiBAN7cPuyeABm9o1yJNSVzfh60pyzfjY
B9PaZAS125GmwJf1gd0uvkag8E0LoKJGm7UvfP28L+K75I9Ob+WRCzu+I5IS
k2RD3rb2X5U7O/BXFspqUGpHNLAItcQ3V6SeF99vbKV1yDWxKNtxZYSjBYIu
8OR1CeYuI+CZ8EKehK6qoq9bD2TLzzjSP+Avgq0c2DmJg6YA7kW/6Rfm6vby
HWBO1/2ScDoA35PAuxmyaBoX1dPBzAvre45ytcFNi2aMGzGbLTFdMX+t7sOi
Jh9Qw30wbGPlMtN7f+etxD60MVMBomRODv+EoAZcph3hlG6WCQIZP0EAL9Sc
TDt+x/4KtpfAYkrbufGVMkR/RzocNMVQIJ9K8/wdyfLSoafiIb2yyehM1bUf
2hH5lz70eYWJoFIGIymEaVMec8PPpwQC2CJe7+HF89vIqbiBpMXerrO1+ZP4
VNyolMXVL744YTAhLoTJZcCMFEy7dxrsVlZYHiwg4FbEj1SW0t2/RLa3PKuT
ZNsyTr1m3qMc0yFA3/3dNv2VNF5nAIblh01kBOYg74j3ANSgHcaFKsTSsHyx
FlFDDbjvhVo1V0ZnmXXG4GXTlNMxSlA/55FshPQU2d6TU7rNkhLpXaLsQ8xz
li+Qely+O5kCVr7MaUlwd8X0mD6eoO6pbUVJ5kUBGjl2XcWoBzhPoPPE0oUV
BMFOF+9HjSr7uD5MAs8D/qOIwLyaZ4uhX0uGTQFriw9Cf2uT6JDB/2tJoI0y
jYfFcrsiZVGh1hlqobPTT667RP3N8ErG8bx/pou//W8O+DGwdpYHwWnBYt/o
vf5DtBNfpAe6KMVq+OZusqx2otCtOLKPGIcbSNx/Vr8o2ovCfzE4anE13Ll+
FPu1AiusjmHlmX/9ILcFL10htRxkZLAsQDQ0+41zi/tycvgBd4a7TqQFjdfo
+ZJAnHhsesIyhc1YF7lyTq+D7WBhzIGmAFN7FFoD1trVqxUhsrAuWvEgKEy6
eax8w5XDm84UZbOd9ZhBHCUd3iwQ4dCyha0df2m5xdy1J5ba4YBffyscVDjU
6eVV1GFdgDW6tVinUG/t1QisKtL5wH7PxDZWVfVcjrtDnU29yy1Ni0NT4QQl
m8Pvrcw/AHj4zI6TpvrA1pDe9LayvDrj98BRq0YZlHIAJtCpRcit5Ajh/UjF
/9TFNGbuC+0goukMamIs2p7AT99l3CFp2JfGpt9ProJ4mNkXBiDxa+8LepTX
F9W9QtSABvSFzEDWEZyiqUJrBbcxcqL9AFtQZ3afSusG7gN2T8v70UqT6SBO
K88+WMBtzgc1k1U3A4JzJQ9KHmbj7RASSGpoAIZ+pMSq5yA89EsM83x4eIJt
SiAL529UoYVb4U8KFvxvnPHbjVR4iuFrmKb35ExMuS/0UQmxSBgyR+s61BHH
qTLq9pEoJ7FNyGjq1MnyWIxcOWcQT3p1OYwESyi7W6GLE49M8MRk+EucPflq
M998KW4ed87L0TOnKiJgnJ20hd/BhOSHhs+vBE4sMN5urN7Dq1Ezvbprjd5A
KZevQRRgxRmqK+nk5Mol5/VqzW+oo98wbGXjxIp/KL3sFpP2I06N283Gcubd
wPEnlD/RWoRKmTU3MfbypYhjD7+0f/44CbSj83TD/n9f8CUGr9xYhemiVN+1
L0RyTSQ1kqz71jT9gqR1/cn0qdZkek6ImmWZv5GHAnC2/xvIAaghp46jPAdE
B3fo761RZ8Vxx46F27nBEdsyUIF9AZd4qDm5IwcimO1QI3LnECHwKqMEcn+4
k5yR2wc8+qmcCSLdUeMFVtPqXXa7VKntSkdeeYGWk7d/VbQ65DifICW47Ubr
5u8xF+uq6qaxdR69JnnmPK42mUb30hnSbTQTCuCv9MaknFX2ayERJchgtflC
D6WujqNpKbArIL8ynxvKtk5C+Dw2qXk5UKridE+xPB5i65dvbqBaFqDgli1u
VmDmFbXnjhJ/92QkzQt5V3SagOF/yUe2km9aaSIujNS1T7pdK3+jxMFaZV2q
shmF93TZuDRk3B8M4/42UPGpaCPNLQ8wt3GJULlQh/6lYguL5M8/lopLtEDa
Pl7khO29SEMmV5yt5eQoNKmwD4iXlOlmg2D79IfUKdGlYwvH+WUj0AECeJFs
9zZKKqS2cYHgzgquOdxy1QoqWiaEDEdAa9H0bl8g5rO1HqEsUikIHwKwWxBV
oscHlM5a+SkXr4dKdtlJU1+7d/OCkZ6Ro/Sh2uaNmrg2LhnuuLOStVqRTRz4
oRD/RhkPTL4eLORqVaKMr/NBHllW3+9Uf0IZkneGmdmh1o0GXpWIhTlmpn7N
qEGp1K818ZPlAH4VOnO2Wl4fcUeOoYkHK7uTwhA7ZIRttsDGI0B4NEFp6Oks
pu7Sxz0KLIObgT4liLeeWKs4hJVTq6LPEBnejJXSsztav2HTon+WEmZD4vrx
X3PLl9ZNP2PGJKBxL3l7x/8ONl2cWHYKU3YtN0XQQhlQPEzHhGQ0hEsQZO4A
vdIAsiP6trfmhPgdS23odhXI/mSmfxv9koBET0m2BPHAZARHwCxF+1Va+iH3
QN1tGvCIHC2rNU2+dtKyVQzmhfli2fUazuTlcMsqyxJPqfoZi+fVsaJVHYHR
7d7C9PYgA2wIrglM2HqU16zRE9SWu8ihogSuZaEwlCBd5ADmbQtoPjydIED8
lMBNloC/slpWwcELPmdO+SN4E7e7cZDWnlgrajihOCO3X24zGy9r1H9Ipstw
cEqkrMnEmleM4Wbzj9URB5T/TOjc/icBY8Bpomm//CnieYdrEc3NmFZPLP4v
qGuTBEasvvB2eIFpb5D6shR8hwxW1Qaf7GRDZ2AW2vx8+lezARsfiHOuF6Xu
Ix+XClF7KJw/ot6OuaZbL6DFBWSp4sAFdBHzuiTnRtIJyKaGrfzYsd/nzBcN
zzDU+BTq4n7rWOuZxBtjCXD77wNo11ha01kE7evbm2dM0yWX3L1AERYzirKl
KMX6oQDKqa2h9tdNnWCtVXM6rIPR8ShIW5B7o2cKYjhUmbVCARYsy7Ojs3WX
Zelv8ExtB36ZziS+iw4ouyhkCm/I9YD6PjdbnPre0fZaTg8wADEM0egqgfXz
UPeA9CVFDoDMSRhkw4cOZWvBZUwpNNbYCe0wpQ2+L2j8x5MAwVITr0SaPo/P
qYX7mbC7HW2adLE2YoWg0TeKDhNZiv5UiIxZxA9wx/a6ycYfwnGfxPWm8qEj
uqzfifKUgKp8CdTubd8xHmqZ3bAHUmZT+P1vhVo2cqaUJ2H6JgeHh9Fr2zzp
ejEfbM3Ypeekt8DrNH4tmqJ363qrPjHw5b6npyM2qpmaNk/SOaRU4Wg9ZvTh
uo2kVI0h9h8ST2eW9nVKEdWOSRLFosulYTO8HRY9FrMcMu/DC5ceimy1DWg6
8dwv0C7hXi4j7hLV/o1Deny5KVur3FX7mPp/Hcx2GoNGJicuXTkWs/ypaYTZ
mpjGJA8TB2sIPl7DK9FLHgkULvtcgw5qi3o2ARte0nliWBMNkqk3Ba8MlB7M
z4cwUjFq39USEUI4hXMNLkXUi4UOQ5MT0jYMZhTKMqiZ0sjfe7+/7R1ol7fF
oDSyJdLvLfL71STue7LkM+NlkPzzzkIEPdYS/7IBuWI0n/2vrT5CiElPlhQf
4X4lO+5ZDN4yTiXspGHj+AM2zWBaERFa+VuCWrFtc7gqTAXFViR4dLiUwVe5
zqxJGSOUa8XeFDGXMck2uK6cABO/fsBzeq205rwvjeuF5yVCAmL51zq0y84Q
xL5owMVheqLXA1NMAktTWoU0zwqUsYgzZcPAnwtySUAG7B3/NFS8w7SRHZda
Q0s765zZHCvvQTOGflfddNEIyzaVmuTYFnCCwLlvbJZ6EKaFBY9PFFdIcw9T
qzy2Cc5cIkneisi5Thrm8OqSh07/cw7/Y7jRPJE7MAgEKAPtJBwkC9Zc8on/
NAKwBIZXnbAdLVv0rN/3h0RzexEYV6RBzaOPwnfVmrEKwmIfFLKCTQAmnd38
AoGykt1LUzbGMZVPGLZcu+5RxtVz3rWNMh/8HNngs1fhDyXN2M4qfkNargbt
IwZ/swG2d73nSqqAganDkc/uT+UeLhY8Ncsn2lctzhKyMJz2NVCThx3qyuFn
SlGhiqDSVIEnqlsGXs7dG2hEwzPnqUG/iqUHWCBeRZUKPjeb+e5E59ldkCne
/43eEM4kGKMzjt4eM2hmSUViH37MZr96yZxmznuDmeM1VZsG5rYQtaK0hyTy
aMdNE528xfYV5btaLIU/Opcztq1ouN7ovAxtWttQsMp9qXV2aOx3unFLY1Fi
XH2cuNyNArDQhbfXStZNt/qj2Tdl5WnPmo7hWzfRU2J77RTAWqfM6LoQvzG8
rcTdRH5ugwiAT6JUcJShFMxYEBm2rrx4ecJyXyESy8P4n0bU6+SyZxvgokSj
88wmH5w7Suwkp8qTl0PzOQN0Kud8EKS8wgifB4mb+CVCugZ2rZ7cikPOxfNc
jFE8VTMiM1sKTyPZ2qA8tKnF8JFjr7Z+J8sbysnfh+XJnEmDFGwPDbUrkM8F
Rk4MoKi/k/DlHN7jvqwWSiaKK0RA2zqYNNGDQGomSfD95iw5zKpHRJL+lGIp
CLKRb6oOR2O8Z/GgDmME2ZoAMTqWxki4RqL3gzpiDEdev4UX7dAlFl6qn6Y0
ii63aQxSih3Bns76V4dlaPSHV96rjtmRLlSdA7BqKITS3sDDIpbx7N3c4IGo
SWWRj+1xnKfm/1fBGteafoU5j9tu3b9hMxph7QIdbK2/nqaHdwMgERaXJnE2
7VoGm+inHDgMOstq0DpGw4Iv3/D/h8d+IFS3eXsxC1qAhpnMe1/+yf7wuEkY
mjBejRXRSNeJ9IJKISbN53styovEi2zsl2wQnj5/uL+kXZeQuw9/i6xoBAUD
gbP6+JAItRiTRCY7FAiPbUKLpGuh8WGs5H33VxHOHH7aCCmUSk4jw5OXHfnq
OPPuQ8p+wtZXZP0tSZgGuJ5lU/hwWpCEhzsynVMjQ5PdShgUfzvmKeKtc5q7
vQInQZkYdy9g/u/utDkrRnyPMMBdHtARC1kTw2h9qoKJ0Sf6p2PAM1ACyuHm
eg+NRdPfRKpXiLv8jiKG+sCdFF4DgPoJenwmWf+RpitWSvEDtW7S4+p52dJp
JzJy7lfVsvoBtoxi666t132jSghvoJb0k4NuUNHTuxN8VS1ov6wYmosp55rk
gd8tpP2wjgTCzHXNh/lgx0R7i6m4WtsPToRWswdy7oJ/tvO4cmzqKY7pUUrX
HYQfjuM4xWhAgn5cXIQeoLSrOqdSGHMT5tlkqsESjj9dJDPYRM9O9eIIv+7T
OCrkBPhTE/YHmefH4ZuGlWanfKOr1/OPGRp+0dX7iwlgszK69esyBB7++qD/
B7eC6n6v7Kb36dSWXCKMNb7OFmA7gLmzj9/XC0I0Ne3h+SNkxbMm1ASUfWvP
EizOsXsTU0HQV6tNQktGTiHvW+oqDeAc0pY/BnstcaAZepbqJyIu/k6yEnx/
5Q5eBHIIiXM5kRYsy94uH/RBkYqYbuT21uXpr2si2lxc+4LwDo0CRqUG4Mv7
BbLBWh2vT2zes3qe1+vHN3tqL9P3iRh2MFQ/OoAZOXEDtJnFO+xzJb+7IgE1
zdv66u0UOvVtqF/lcsNHABM3VYcZ1mf41crBElWHi7j7LhpoE1X7I0rcxu0W
9r+c1xk7eapjW2YrjIdACQ6SCGcmzAudzG9rGWnrO1+C+DvS/EwGU6tPuxDC
/qyeQa1yFSFg2O4go8rTgKKkBJESJRa/g/IJVX7WNHIO0dq7s/u7IBGjVAEM
44na4lYf8z4YGLrT5mrKRyxEesSo9qfqZAYLqw3JGjI0GRj6M3OjrF82hls7
gSyCsWMP8ywodRhmMRwry7H3Dk6lXnvsm68ujn+zYhbvSqisnoLnHIhalHfx
nMyPC1BDsuZlyymc1nF4v+8Zr2vd0cE3m7neU7qaGVJ23zEj0LZDNmWheOYC
F9ALtCwkG0pR7tCgirfaryTdK6lzWbgY0Z4tjxCU1tHT0BHQhnOpWErb9A03
LI5dRsUZaps2Zi3IJ2snIbwLw3XXfyHCaUU4wCiGI3PUkVUvLj+bGSnkSgNj
tkLYhcEMbJrg3gny4zUIqMw6bMNuN6/JZ8GQPPU2EFebHS9oHDCxY31IKEzK
aoADK+kSEUkrn/7h2ATRt1gvJRxuZnOntQ+2hnrIY0yTgBFXh1W+5uD6+Bff
EnJajrbTuonHmK3xFqHQbRMYidbtdaXBhFPFIM2Hq3kt+kwl64E8DcaYJJIq
ft1pgUeQuh0mcSqv1E5Lw8mkaxd6snfFN7Sla1iN8ISiD2FL6PpsCrnrOYEK
+A5FBzKFRBMdgcPZkBs1i82+djtTlKMnNaf29uJdsRKR9R8VHVhhnEgiJkL6
BB+Q76dg3PpougcOew/4rO9P6OO5rVIHrGX1RnQe5hdkhiK89H3riGJ47FuE
MkWwFd9Sqmk/0RXi7aK/aZuNTkI420oJcL/J3iiJFQY0ItGh+PuPFt8K52Kh
BjvCqnaHafFj/oy9j5WTf9iJXDe3yM+pc3vPFaVGwTc66qBkyrbRm0GKTETe
cWAvCS6tqSvCMZD4jSIQpeYol6PnDe9lSLKGu3gUpQJ6DziYgQ/h3OBqORnc
W1mS02w5KvhiPLmTStdYHaN3Iw4wreEz1pHH8EfnMc3TF9mIsAuz2xzDqUAv
kurj3c1CcucwwKz1udTY0Nd+gTsVNp3l12hfLIANR+2I0iFBi9gKLes3WZgB
wtn5T5y38d6a9TDdpKIB12FkDDR0fSAZKKm9vHD/rY1AK7qMgn43LKCqnQ8t
JH5q9Xv43NwJrKcZk8cTXBxBeoWmOfx6qgV3AXrwOdl2JC+wLHfON95eEQ0V
eGD+PFvplUpfOT9U1utjbSCHN69DipUxZ3YRGXHJwd+tIKN4dB5pWQxpBr8Q
Ng2t8vR2mSAtgeJZm3yLSMf2j2k8u3OcYls47W0Z5ceJPLibuYVThnu+4KXT
vtgwHs7Q8B9O1/zl4ZLoAbiNJUW/CizeVfAinNX/V6q5X016qSSyRWyzfO11
LPRDfuHOaOQRGlDB3aY/jeDWQd+J5lnePoBdUh+ySu+cbu5rrok2DR2x++yz
40QlVqX9tYxLf7Hhd3PTghWzEDeQ2ZIYqdxiGz8u7zVFliVhhifQpZuEtpIf
1yCVNAWqbRyFB4Uqg9vQttKv/hHhRg020rTMg+2BS4/JZTEf34k8fAeporNO
gC+Ozns4YzD0ITvfzfKpczLtE5EIDZh4NW9aENojXWN3at38pjag3xzISWw7
4TyF3XDwby7+5tVTBAPW9CZQSsRM7+c+7tjRoIF9TH7RmD/21MKWx13N683m
FNgwdU8gH3RRLDasiY9iRnQm+KqLuBgFKvBXdHos+n/Y9kJHCfmm9L5I0mHb
kxHPECTAhyW1ePiaLdf+eRufwb2nV+qgMYXdsM1Fun2GRSJCpvmZ9LwDxSbS
eHIQZALfGWWPF0l41czG+V6i/IrVjj8hx+5IjacPOfXNljMt9ReDiddYKvKN
hcLU6UakX7MHjmHbk8Qo9ML4nxyw+TVkZ0kI0/L7Gkl47V+KWjy1eTpP8mwx
HTS6eFD5HURDeJAoXeHHxZuk+rNDpNucFflnuWTRaLto4y/7x138g/a4YPbi
USxFzpIQ8qdQNEz1/EIYmaukehrR9g2VkKR12dTliIF2k9oXjaC5ax3rdDwl
oUUmtkp05wifr2u3B7RtU0UDY6VuONs+2qNYXhJjSlY3zxG4vHhKrkZamfTk
MiT7dvTWdcQK7uqO0/NLrpVq5YOQ2MS8HwAM9igQf18Q5AoDFhqZNNJUzXYL
xaCbN8orOY2sKLHk/HI+xkWED/Wif9wlUCNX9g9CPj65d2oz20jutotkd12v
8BbRxySXwvoXHHW/Imb2ubp3qkp5kAgieFdPblPm8cD1afivNY0VX6PpZ/NE
q28KwqTybUR42YKJhsMtI74IJ2zVd0byGavl946Y31KaUxIm3FmdJ++gsPNj
mbs37fkiOa27LT4rNevgXoUHIxK4sguebpQkyCCQc6Fk/gJI/7ZkxNLEYkOY
2+QdhXEoM0U9+gABDgCEFWVEUBLUciBeB2Tf2/Qb6Zlftlx43ZAXaChdZKSC
JyWmkDXNyWhse6GEN75H9Yw3LvEs791+R6D3g9tt+zdi5om4miFU5mCQANXq
RSTSBZ8gooej0MpCyE5a4lz1TL6W/ckJ7u/ledoyZ3zXV2/aGLfMhKKNaGeu
2yXVyGnTCl3HFJEOOpGJrbvDuHF1WEcyfLMjGfgY/JO/s3wDUP2uAHJcPKp0
lg5P4GmzZZ9/r4iCYPrFdmBTANxJAyiTyAwwa0/CBa532uT83UJn9n6kkqff
boUZtPUFmPDi5+hYb7vyb1UYd5PZdV2fRihWiwnm0O6VxKrtMG1d3eBcVGAP
p++5EX89NmBLiG7pnAGYflCBXYeyLVxVsJjK6HlWgbkOGrM0MnAT1zOeMNuZ
clnivA2dig3/nZJ8udVfyv89JnReAjqt9af99CPN16z1XyqilI3xSiXz/pzX
ScdEgDJ+OFtSIFXrrHZt07jh35zYn90Gsdq2vwJk2xHAy2d0s5yQsB4x2i4f
VtiB3nIbkJFMOnmoCWwSb+e9vz4+3oUk3jcF8TNL+W6sL6qPbZ6ODHpUVTSb
lFWJMnkEp5uzwhY4s4NYruHL3qA0qUvG2ZxHtr3XeNSQfO+u/UmMAfXHbj4z
Tvt6S5HXtdiuJMG5sCxy0VFbahLr2v+HyC1bkmEWMAc7lsy7OrNnP14IRrL4
JLE64Kf/QINyyC1ADqnsQU31kvKmHZvUAkY7Fg9QZCgw+3jKOKndIyvsO+N4
X6ES0mI/6C6SrQ43N2qxDTZTQ2PSnp0TIUCKPYq7Ret8hOUCxMBrSn6/2zT0
PzQalHHwrz7bbfd9HLJHpt9WUu5R7OWaCUEHGB9QFqqiHYd+qM3KczvQJfbX
+3z7AtQv9MT4ZTWCe9kKTo2IU5oeT8kK0du3SsRQA1KaVhk8jW41rVgCobbz
eukPQ7TnCOlwS8eTS6tUa0KsCib0sirHoYWpfpYi+qJ0oJYayNNsrNktB9z0
FrTrLjNDcT8BLFFB9e3qCT246Ns5map4rtmL7D6fo0+9kTe0iPBQ58wt41+V
eWXX1nzyMXueXvtkUC9jDxMdqyFhZuNy8VI1eTjpVLw/u+kuc8V/arSsDvcH
NKlZ/L45JxeV+dMIExjIkzTYhyI8/DENUVdNYKN/01QZcb1v9TitfBLecf1/
xTlNX78bIYc5T0BwYgS5AzJbSqQ9uXINNF1qxxHc2jDDaTTTTsjGgSb2K+SY
KDSpCFqA9Mq/iQb4F5W9SccEaII/DVPL5UPIwZHiapvAvjpVIAtWgoPM3k3w
KM3GRhDPUlx9niWBH5pl2mN0kJ0OhmkV0idFC0KpL2bkgxrqRDfh9GWTemo5
gXdXuJyskeG0I8xES4RUbvFyqraAVS54TAuciC0LlSJ+/9znRrCdcdku9b0M
Fvc8+FZnxH5XbRDBYTU+GnVjgTZDd/0ATQaIRBqr7ufv40CR22lFIF95Y1iA
EKkj+5Z0BwFKnR7DBxzqB6bMWJzWkhy7mAl/Gmj8nuCpAA1uk+mwVxYsWNlz
QUl3ZzhuzwV8d5Gy76PnFIGMEufqvwTdOdHn9fj65rJqz6jr+QN0BMind6HX
W7dbqFDuJrFKCgWmQcs1cgp+MrqB5DyIIvx4enzixatf/J0MzRNAT5LjIync
wYCtu1O4Rb0Q4xNZTZtRFpN5jBeK3NW8/ujj5a83Wyt21gLSV5gSibaj6WWZ
n9irrY509a5D+0YcvkANd5O00/7jN+MZh3mGDLL/9oc7Z9A5xkQ5YIjcr6u9
8tGjYPRhTZ1zlE1h/appxv/IK3+KwuktZN1S3NNoxnDhxvdwyR+TuIMQ9Uye
CvI3McMoLcrujSLjexK+ysZh2V9FfdEh3fxVqKQ2EEOxrrTrM1+vek8s7zHO
iS3gAjhljpqOW9Mz/1nwfo7+kz9GVKVwqmAGTN3NzLj2DK3gXKsdydYYMvzY
hiG37v8iIWRrewEMV4X9KK6R6OqkDn7sTU1cYE0rHoyFnutHyFruDg17uJ+k
W9/ZiN4AEq4QchDPGj5Ae5FSodMRSffVEmN2uR9GRr4eHw47Rq8lwhVHh6I5
6vbqJZnUWFfWmj8SmmszQu0CKUm0o7XXbCE39ANDpZHOAK74IoLifZKiVrLZ
RNwH8JwYXKNPWrx1y8ODHiLQPX4mWxipgc3pjFl7mWcr4k4tUMufcKF7x7kh
1wunw8Kib/qbc5Ct9Yr1sSNXEmVxsxGSbZ7tjftqHS8YKX6TLLu8C/8Yzt6E
lXp/K4xNoWPmrUXr83dJL4o7RBn5HuyZzvyCBYleb2YQdy1ePNhGMs0nbJuq
RrrQqBAwU7TQ2oTL6WPTWb6HiBm3kaGuycCtGs+E90v54miLxeCifmDLoYd4
rBpHfW0BDUCeTb/EON9lnDI3qaYag8oL9WGn1pnopd0FN2YusIvEq+UvlhmZ
P8iDFmiM5ELeJHxB2LSGd8TGB4cvU17G8bZCWXEfvJOrG8l0joBGnEbF4sUj
8YqwFSf6jJbmVbqEwW1NIOVhM/Ex1oijjNKsFGTJIAllmSkCpW0ILeHB/mAW
NTA1XgbciDLXw5kxVVHMusThhlTVkjt9Cdyi49CMY58RlfCKJPNQJka+nWOB
yuITeMsSD03lnAtBuDac4T6Fj9dFg3vKq0TgifRF8DNVLNw1PGD3LO8pVK52
8mN60phBgEwLfu757gsvUMNahIwvtDFd7NgkqiYrAhlICZUt7a6MxVT0EUCu
ytVObDYavvx2PZBPZYdjwAftIqSiai49n6e1gn1cM0ASolg/mTvZvht8fe5q
QeYA8sQbjq3mVe3DpxHleeykOZimwKsxb2xZ1cHofFrOhmlyd8Lwmj+2Cq0Y
jan1Cgqu5SI3D/OndpUUcKdh20WopXU+tV9xW+Xq14eniASRM+1Qqiw3PdGi
Rrn3bW3lOBm0Ufa5BlLqNH1SAZRzRp+U7VGyGv7G/eC1/nBSOG5jbPnhMitY
OwmLMAGBuypeyrcaJFYu590vmrn9I/ZyxUmYIkD3eMsqUeWbrYp0svNKFd+e
Et9cRHnhJYH9n9zcPhvM5tmus3AWoA9bue7OCEAwUgi+zlASyLEVKi/tjKMo
y/weKTLaDSuR4K6y1eRZhVbwleZ+uCxVe24APpZGZDSG/JNpgjgB/pD2y2PT
+x/4hF0iQ73Jh4oNIROief4GMe9JShejra5W3x4049pBM2FzvbHNbYDyaehV
Y0udkEZu/AamJIxg0FCwFzP+nx2A023MNmSLlTCql5AFzrFgjAbbhJe97aqj
ExwY2LEZ/mlQCJ23u39CGSJxlzUjZK65f787wQqd2My/SQ8agWOPgtFh8ZuQ
2Luper3I/nDz6mhwmvL6fetAf998E+j8jsZV/f0wXEHENHQRIZqrMc62O6A1
CsdReHv+3HFvF/80RB9enJgKSwmrvlSgsDPZtIIuA1uZpxDFQkzV46NKFPdC
Pdn508l6Tei2sOg6IeC5NajJb1FABWexaXqvw6+K2MqKtQHDWHpWzuRxJzCF
gEevkj9wBBp4MBkFx6p5cOGJasYNRmACZ6UqxY7tpb3HYDd3rXSgkROtZtD7
Ovqn8D+AlsXqpz2sCSSxu4/V9Y15300E4pu23xE/Gi+RAj4Cyv6+80r29lSX
CR9uao5jnOzzN6YjkoGZgPzzzbkjUnYWK3SLb2IvneeFCISX+47lxRUXCGpY
7tbiLSWbrj9h5GEbPGSSVMkXDbWu0nPBO+xn7L49xdsxPbmE1tPbMB1Z6xap
swnwOMkutB6m7BbpxMPZULeAYx5z2r+PNBAFwjk31ny9elujE1ianaju0JQE
b0cwYHqA8HP8a+D07evrKoz3thVx23Fvo2Ca2p05Ns4/6OC8jZbMhhwo+CO6
Gc64pa99OzHipDcZSDIjdN/89vsjSSFCORsbL2qT/Fn9sBnvqTbFRGpka/Xc
iNFO3d4OkvpgVl9VRkMh59b2RfoQrwusumwfcwE65K84kWNXb2Bj6lm0CPkY
dZ/IGgOdf9eGiostSuu0ubm6y95knIOieksyVAt+yJ1gL4lggSvKdiNMA7Mc
zY4AK3SYtbyqX5ZyRncnC1mZyZobMgmcLa3EIo/2lnByrT4Or73OpKy4Q3hn
vahtVeBfN22ITBm8/ZLQC6ITQW1Z/887UwXzvylA1wyoQFjyzR4/AE8jN/uT
wyeXmG3N4iB/FNaBWmtnUGXBGMj34Ny+VOZu7lgdpI1DUF7rOqFOOYZYbOjl
ZuqTIQYqmHqFlBs/5cEsenx0EJPU3bNg2TQS+oX/GOTnqPxF0dQr4PjWKFTd
zgw3lEUSeoe2n9dmmQuWyk81SUy58deBPw0tvS8pCaSfNMmjrf9EBjZ737j/
1LI/vTVVBQ5aD0Bk+ilX/KmoxqWzbtIhrwuMFJO4CrBQ/RsW/LeUDn/PE0eG
5O2BfuEfu+XAOctnXSmYtsi/Ri1HbxMwCAkIFNw8axiDX6D1qFPh963iUXUD
HCg8zC/xQ2G1HnJMWcGDe3S44mFJvvHFmch/FaNKLP6/kM5IPfXQuTCKZmvM
/ELcsXcBIvEe0NlAPifuXbZXePWi4fDQ3YUZYAhuH50bkrCLEWDrBq+oMhH2
c6CZZ933WXZXG42V1u8Sus/rSJqP6aN+C9//l6/1n6/WmDI7DyFePDrccNwu
bs/cVfs2LrBs8hKOwmoH7IlByOt7z9WmEr7tTNqOLLzAae1zC8LLQCh/+dNG
PRCKt3ejVEx28PLtpkhfATSynFhNj1MaeD19LCfXbf9NiqTm/6oHqMdU1wNP
vv199KHWz9U+XK50i8SWcvdHPIDw77uXQNNLMfUaRo3YiC93ebbnlLlcLErn
5e1Re5/SQsIdkNu8qQgeMHghRbm7RqLmGyOrRHc7gtmGLgpFUT7QgJvMhdrX
Nvex5eyP/i6d+8ZzbPgMN5pWDU5Tb/txyMUIyWTRD+jmtjJodKXIoZt1w6fw
9knPAAmKP34D0Qj4J4qnDOiwj+txULKwopZ0cUbdkyL/dWbObKIqucXmwzVw
saez72O7nU9px9SWowiASSu2KDeOL/WsfFb9JSiIc3JXODAezVWq+yapVzvr
ouPQHSuACEH72kP4+/tWJTYRQOCMkFy7yx0bhwGmuYCMfiZsuzU22dAZIkvc
BiwTr0oi0zWjeWJRuRaMC1DT3Ipy5aiYbtX0U1oPJXcLV33Gkxej0+A9kJwM
TsSfEEE4RwVOf5MwzddX2+UQUSaSabticw6L5XeWok3wx56vg1Nih+X52exK
S/sFh7l/jNSRwayFEogllbwmr3mfPdRVclXHpp7lBgxQINLvQosElFA/C75v
HuT8GNgfeHidhnFZjhgxyDVEAKxmh5gcn3jHvKg6PvuyEHftM0Kl1pBz2YhT
RrHxQJMvXiNcJ+noBzOH47qST7bLVcQcTu2jMutw8B3tFzuM4wZ+3XobndRH
xD4ZVOb2RH6NOC5aL6kxGZDdIwRXu4W2wrUwxr7II4x4o0O8Ro+66GaH8wiF
Yyra9w8z3hu9pIQ8bTpD/cofhYnEKf5yqdHbCGBZy32Hgk0EzQhP6VFT32JP
AbmvPFs6BRfw1+qZWJU3A6OLwh4dCOVOCDrG9Fuu9gao7ueB4+97l+r7m/aO
HNhywPn6gJZh++OD3fN0XZIuqSbEj7zRWNWRtXcWhsOsQoAS9X8cqT3ASSwf
Su0wkbSi2365hou4bs8hhkzr+TZaJM3l4RdHRxD46RFza2NSFn+6UP8YnMVw
1ZNHVOr9ti7cYbaQlvI/9S7MOYmHQkzphwaEthmCxNVu8NRUnxE0MiMYFBOd
nOMlHL/Urh6QIJmqaGmJKK+TflNIiwXNt60CCrUlQdjNzEuVKzhTLfRrbUMi
7FcYiV1U95sX5UmLDaXuHjxAh1J9q92eoddED+b/1is4RbRH3hy5IibRR8fQ
JEHG2g8lyjZ6yk6kt60+fOO4KgdPt4VGGPR5/B5YgkmiQ8emEikXGiv2CiAt
uX8S/lqPpgJqfdrlmn7PFnoEQPccrtQqdaY+hN+EpYE0v5NMoseudpPmca+V
ImWz6vuNt9rmsTLKnUNvDIzzE2pHbLZyvR4QRp0pRPEcUaXDl9/emoONT77X
k9amq1VGnRYtk/oT80Ojm3ZMnILR/ulCNtK06o4Rr9F0KglB7yBP/ypP8ZGk
ea7IftCScbTbSjdlPvaMrHY16jKiIHWvhZVBWO4T2ohbgn2XL+C+EuUJWvy+
F0Mg4M5esiPi0So3W5wXh/5Lxwgf6yE8gVrAt6hc9W2NTbePlbiyEFBs75Am
mxuCPtY2XondeHSWQYcW2g01jf5mHqlxtB54kavFca2AoaBB/Xop+TwL9dzW
PGVVZzW8KS9Kue59iapGikivX3hg64KxA3Zhe91nFQnDbknNMwkmr4uR4awh
qndfyigbvJ5xusb4BcC5sR07m5+FpWRcGvc3gx0eDf1Z3ujaDB8XKU9UNKfE
S3qGcG46Kyj7pgBkQ1BVig7Wgm/zYcRdI+1ej9HNbf1jxRkhiW2aNj+lf/Z+
sSns1hWgRKape9Qw0lJqOmEc0KtiAJmwzNF274Z15K4bZEo7m9voJ7MJTfvi
Gbrf73gTJ3gd9LBgVfNAsxknNbIB5sVoWrDAGsWlQun6eC+y1iRL+OlMSUTy
ZgIR7lUNse0bsqEW9BOrMsqKPDEYFPO9thpAQSO+Xbj22aho+lx3PPsWd+ls
QgmB57KMXucgJODwQQT1I3XiCYHIac16rp/YBn45EsqJ9knXeEb9V09aJjFs
GZq1+8r5baoChdZ+wTJx3Rarv6PquWx6HuVztEQnJRwDTwgeDwVY5Q3nz8IB
wQTyM2bKUsPGY8nZ3KOznxRtHNZPK5o4c2F0wiohD0N+yVk0x9YefXYcRIq8
KlEvW8mllI0s+dho3WtnxVDH2WKLcSr6+LBdB9VyVFeGU8/Cv/m1GG1po3+V
/U0a9i52YTL/Acwi8rpGC7nO4rW/KhZ3/urnGm9PnXEDY7hKUroWw9fOlKEv
0ssXFATZSdMFyE9baO2nE66JDcMZZnXvMQxBD2LFpY/DUTBiB1Kpqwd7LcPN
xGidBSUr6HCkZ5sbd0XveDjGSnIx+IOwtmmTAH+xC6irEyO8FJy0SQrHQLqO
UqIqM4Lt1bOlHS/WkiNINvGIeEeirLWVnkQ6MHnCiYe3I7371YQ4DWiOjehK
worHPUWt3s55QI5QLlZfHVAl+vH35Dw1jw7ABiKBERT7GbTGnXn6GjQJKbvP
maqjNtQ8jrPlmOhANEQD2eT+yWGMg7DBpIye3SIauFRbeZWsBu0ZdYCofPsU
mf6/BoGzM2OAlxGGzmLm0YTHbHjGkgDhY7j7vzniJLMD31zoJRG/GAiND5Xb
qnpjCf8JA9kib57N5qx6kZKBp4NGyDxKavbkNwUnvC4B8G2HHSu9yHqpTy1Y
WGy887gEk7RyvsUiFH4/5S6mY8Mvjx0M7mMLjxf2lpA5Ov3/ZMGDogg0ARJW
P26ytTO7JqmkYe1ohg0xqVGaUpzSI3Nk+FW/NjIgg6dPJQ45DU/otJjA2vRV
L9TnHqU/jWuIYgPvFlrG+uxD75Ck5hFMxbY2D9ZJi+nkeqyjEYAC0gzXdaOx
DZtQV18WMRkAusjOLfeKIYwm1b1RjfOkTk3eKrqSNMUbrDXuVCdKhvn0WdwI
LzetWYSZ5hveXgEpbFe37mzq+Wd7bWewBnnHP/e3e307G+u+Nm94HHcIdqbj
4jNjLF5uYIkcal0z5AXPkH+egG9+94v/bGfNz0ivbV3YrbNYWUp+kBs0duW1
1v4PZFT8u/smMC/cLauk1y2wvk2/SHELb2A2TuJVXu6a0tnE1jJLS1RN4sdi
VMbD3LrpiobuoT5S35YhbKzV+hAa4dp3BfhO+vdV2HtknkZaflLdwMFRv1/B
Dj8nYG5uYM5GUmeCpI5Vo2BRCVNFZku8b/x4+QBJYQ243p3EpuOS7MvPWFAx
ZlDmzT60TCr6iTg0nK5uDOCPXGPnS9GnTtTSlqveblrli+1HrafgVW6RB+AY
Fi6Ir7arAk+Zd3EDN4mkfKykhFO8iNO/sUbFgz7uJKRY/SW9A+TXNSiUCNNA
H1JhRnaz1teOYm4rcaijfwFfC1S1muc7RTQr5sZd4OUGGG67X+5H7sMMmPlQ
cK8Ge7J90i5uhiK1ZnitZaTMLXFcFX+O0f25uIRVa1uZMF87JH+U7L3Z97uo
hqyE3lbfCiEmFu7qkZWGW2z18fKRR4XOa96TlSIrbjiAd2q/IWkIKpNxfLe1
vOaGz+orU/J70vZPiYRQiB+0zy410V78fPaNaG4Hd12ZwQz1dHY1SAN1tJmt
0ssPWggywuI8updOtb2ozx3PXxdze54XVAOErGK4SbFJcaP3Q7OyPp7BZdH1
um2/bpFxP23atO0FvPi6nlMNr/bm57Fvr1/Tdu9Mdws8z1LZ1E/ZRA6wh9Yy
JTmdyvLmKh/zgLsrz2ipAWJRDILZ7ddEH7Gxt91p4WUzaJpY5p/qJpPeXOqs
FxbP42g2tGxRygdzoKyjBxXPfgIle1QT/jDl/n9EmSBoTcUJsIWQTZRvI6MM
mdgICgi4kQwB0huB3fcexzDwA4K8LSKa8VXqnpMzPEzZqTqTChyffrehIcOV
MOG/8GlNss6V3WtJE03R+9JarvofAlW6FOO4IiK2AYjnR0o6VtMfkxL0LZlQ
LiK6s06rOCxIBvLMrzV1rwG+QChZeViG0xtjdB+2bq6DxT9zc2YsCwEPKvE1
bq9A0VHfofVvfL5WWWH9kC70wA0xnsMpZuUhL0ti9ay6t+bo9qukdmBd9882
DpbOPEOHD80h/5K6Rg8ve9d9WDjMhxf5qK/T598FHU0XOBTYJoUhZK74nOWa
aKwnbSgOqau6/zC0tJ9bvZUM8+o+kKNEwcWfd/OtxfTtszXpH+H9RpiRSHjH
IVwdzsKvA1yQ5V9NWWqKUYmZk0kGTtHdPFhfY1btKHwPk9a1tfAx5w9m8c0N
rq6Fn/p/WAAuCEhPl9O3lRrEFRTt7LhucYKGGadj5cyKdLz726sP0YEBSNsg
v1uITx95SnLyE99FzNEnlGl2RoXmb+0hrHm4SWZAj0cK0P0v0kW8IghKYfu9
ezfvG8JhnDK8Ci8UUJKgfQml6L/vzk0lB4+XrL8a1HPzZjkxyaEPVa/AdmXi
936ityzk58r8DX0orejGIzXpWu4mkDB+wdXfQLEadN6q1bWuaieHFZ3DS87I
gMjBa+iQhQSf631eCfohveQSOnlGdI5DpCntBmaE/47D6ZwcxiCfO1UcMtxe
fMUCK9xnTyoAlCM8jg053G45D8KeiXEqRLcudW0WNfyZg0MuqhvxkKYKkRpi
M/4osExAe0w3sp0s2pVVc+J28bP5DI/GECosRdhfSGF+Tco+AYKPfOoib9fB
MMfhdsDSs/1rVl1duUP92RWoHz2HhM7P7Ar1QsPjU9fgiTMszjjUmrkpsa21
8EkgIrgFAFYbFKgJugznaDb6E6Rn/yQRmDhYTeZ3l8S6F9STXVK5Dj8LN5sA
4KiiiF0qVQWhFjChWagcNFwwB59RCIm/gHfr1t1DlLtOdolJK6l1ektJo7TI
M5R578I+LNs3c1K9TdRg0QM8lVE8d1q3Enj1O/pWd46Xq0nAypmM+K1n6TGf
ZnZOeXy3Bhd+slIcYUAzZmH+FXdfuJrVI7mjt7gtYjvK9DiGjRa/J9WbyOHC
1cLm0t4XwTTbrBQss3p7PdHxmvcJv4rSw2jV1O4gtg1hl8+5RRIn77oxhgEX
aiByKJuS6Iog9KSmsOPUMFml6T9BPee6LK82Txy/4OSx0jxo1WvllAXjmwBQ
PKfbyKTWa7hGn2ZXETeUfTwbnv2aFrBuXkPETnP+P/1w9eapJrkN3WbQAijt
Csi/4pNvmcTi15xHpD6jsmUw54XwB3t9cgKgiu32vGn9+zuODQgZW9SB5AJh
A8x1Vn2XaVxdCMYuSR28H4T9UHnad56Qt8Qe/Qtqs8e3d4w0UsM011BxO/m0
Bm64QK3/78Wy7w1D7+PIZgpAguYu2iR/+9eDptWsP1DOJq5n2UJQB0bcqGJn
gS8AIu0svvOvoMouXvq3EOtOhopAvKXUD+3tBaDbtHqj/z36x8vT4d/tLL2Q
9qJ5aP8+EwcqMibxMZs7w7tgGmXv2BJ8Kwcl7qsqCAyfpqX+48NgczinCOLK
x1Y6blY42Gx9bW/k4xWjXDBD11S2E9bMs0/KIzzKwgBJIbh8WboDybrWNMTm
QXLLAO8vCGeOO3W0cjBfUxok3lOOkclEqk7AyPHvmSZNGpyXDTcNbLsRYdMG
y1Lhw4NAgH2Oo38FxeQeIPSHSEQg8bHfELUzBNq2fjJ2sjgH6u2TDhGwkxgH
k0qX1DVf6UCsPLpz2cFzvlqqwoeF67dvuLYqm4UD9/0AL23kyQI9xlp2NjBu
F8Dy98vX3UAAQTuOmx9taD3Aac4e8qxbPbrF6jXDtjdRoLLf34iUbM9vmcr7
SvEupHSklYFKvMyMrhVzcuan7ahR/eaPtLxQrOsffyOerFIICEuo/hE3HOJX
oim7MxFVizuIKLWQmfBk97mF5nrMVJnZJa7bhEQBTFf3KJCoSR/tihuXi6Mk
ig5ah4yfJ9kyszFfH1VDa1GqOBfey4CbDBXSBwyKjMTq0kvLmgi/91qmE2GS
pTWo84QJZlO7pdCx81S9AVTsOmu+9chKcRRLHLBlZIT1ByRKX31QGnfR99jx
8LmRw8693hfZwpMDcnCd/l1ggm1LuBvDIn5nErEuncTPseXkrnkjEREtjwia
JE4NxHOkXerjBbJiXUSXL6+mBuLgHZYdmVH1Nt94HNSRgPQZ51mFhrt0aSLz
Y0B25dSOVcjEJfsqE+CNkc0qdpmxKMbOz6x+ExRFmQjsQmR4LcdKUfmX/yzN
ZiY9Wy/4PLhjjtYBmn/+n12+qH6yq4wNhM80IFurCnmYAhaMUNWcugc8Cf1E
9EBkijfFTaZRVlMrwqK0xopeir03ijD9k0gohUpdKKJOoqXeeLRXrh6wxyA4
+juYb88gyJK3d0vv0hHy3T8WuBjBMk/XsZv5BsCIoyk2DbozqDbkfNOjl+Ax
uEwrlZ+rzKpxtJimkSx8jh9ftTdWeVOfmiacugEcMOkn7nP9aUlMb3Uk+M6m
InRkJBQAOMKnNVeDG6uhkPma/BLxBkkUYhbupd73mNI/tYfspcBxWDQP/y/y
ASkDeuTcdm1feIHyghMcmLTugB8evB2k8Vb3YTp/JJTxZqOSRwz/xZ/l5Wna
FU88c97uFudPxhi4Z6VG5JusDxbxqe9lRQfQ5cotirpiaehp05/NrH1SjWwl
WiO+zJo3NJv5Bj0MYycPqd9ZELVXOmgizdaHAE25hyI1oLR+zo1Q0LjsuB7C
u62nmQ+lm6EYdU9ldgk8uVR5X/7PpmlpNuyBGoPYgIKvpPPgpHcdK8qR0P+g
BDB1w/X9KGy6m1ZU0Td0Ccw5dBCaemcWPGj5Ay/8T+ZURISZWIqD/3YUZWEk
MiNqNriRaRtC/d0npEPCQOkR1mGBp9VYUh3nBRRPcQpb5bS96sskUxKRRPT4
k+bHDHSR6iJyJzHXBmG5C/cG7RoT2CikFJ3Ly4IcNm0AueRbufD4c/f8CeQB
b95ZqnJNAsdRUHOHPo3nt9LKKdkgfo2vBx/oeAUOAy0OpNrK7lzlEjnGEsDn
lYoJ6SsK2CB8ePzf3wRcECXGTFcUTN9fiQ8RqBrjx+ebT3vQK+Ok1RCN8HfB
4G8dtInVILVu5uyPqlVXp3rb4fwnIvmBNPpIaGja2/BMAJH7PzJbDlU6HILw
NMRuZNCGs1xG0QzVPBBGy7RyNUc9DlhaUe21HYd1SgF+uj5qz2XyTJ3D7AUn
Txd3kElUpu2GghB/bUaM92losOa0D/cu1MtLO8a9MZmlmh2eqoH/7zTA4ZfE
7ATFDoSOild9EtmNnEkgmZEYOPTvWhwG968eZzunIlvxEIFIpLya9ScSytk3
xunVOxIameEFVrdD0pHrfhjMdf2u8YTlkhxbyOxX6yCOY4v8oQ56xW8Pk4Yu
9Jqb5AwjImmeRD8T2SuwO/G8LNKDxvMxP4dEc+jKzW2Tp6CNnMuELfGQ88/a
BAYyeAov9rNbzJA5OAUMsELvTC0qOh311+wjPKBoPluwDucL7o2kcqfeUaNS
BldXjEf1neggvAI/aZakXRR8EAZFuYxohAXaVyq6sx6Wk1WXlzh3eV7EJbiw
ngg5sRgcF+fZ+wwn65gEDo1EgPOWRtN164Q1DjmdJZhX7NH9zr5NgeFtNKNu
9LSkjKmV3fGyU0FjNu2RD8iQXAOUQyfOP7xpE1FHzQlfGD8+53WnROv9bDBh
48woiRppBrtrOu3GfRjzJFY/q31qx2A74OYcbFMfS9CwrAcND1WN7bPHE2Ko
0FEHs+EzivhC6Wr3v/awmMX9u6WYSOH6m4quFR26VtPl+kP/vj3+Bb222p9O
LOWOwhpWa3D4R5Ch1LUoO5d3+PNzEsGMBPLgoo3qh85hzYKD6Xrw4d0MXLiR
9n78lc80d84hX1xGLaWPAGkyJ7/v/3aCmC7L8MBnCtQNw6S37NKGxTe+JWVs
kGWGI/8pnZvQCxT9/ttNF/0YM7AwLGvA+yW9TgESQlyjP3SUJPzOegT3jxBR
pPn4ekPYNj1/UIFHvNz72avtnW3YvCa+L+Lnp3hFqv8IrwZUok2msNRH13b+
rk/BbMRnnNJo15A4TI8z3TWfJtdtCLcptqP/auDm1qEHBNxpY4w+j42EdCs6
qmzRftzWbXXnLv70UArd5pdbiUQQXhrVoPAIGb8Q1hxqx7cw/Z7bjl8F12JT
RIoVP44bFPfwq/e7/7zEOhNa7a+HwwAyyZLuWifkNEFjb3Wkm+okx7DkwgAc
5bw002ksZ8uiLDi+D3quZyjyAwKMSpyrf6cmq9CYcBvJPdhjXyRAyO4SJSAb
NA08eGm2f9Rnmlaza/7f6Asim35LsB892Rtpw7wiECo2thtVEps0Xu65rwLr
pq52LlsdNgEox6PTlUAgKFMPROytb9617m1NzzE0Xu9xJk1x6tNwrdAyPXIz
wrOTnmvT+DULpEuVEqEFCtoYSUpKVs5BF4Q65T61ZKOmnn4cT/ItVmb1E/Mw
U//7BsILX2jWi0mfFhTWUdibIr1QAQj0c7VrmsBamaYxuivc857tWv3DBn1G
rPxumGlZnJPbUG+zpR9HQkg7Akk9VFlj5DxjYV1l87GdlgeSNRFGkUK/SRHZ
W+nMADP5vM33RNxRYTaRjBGgILsVlekr66ioRCrO+8yFbE1Z5tn05s0W1/e4
XyNYJ2MSUgZoKEY5XpDCe+tRDnxsalSQoTfL2VBn/0YX2WAoK+PBXx2+s5/P
MZE0vSJ3WMJ/OlhehBmHUi5NGyUYExZIj0Pt+40NTYK7ZH5XXY8Ui42uu2UE
HI7YouEq4do0oP6G5tJqnDDyhAHAQFZnhLZ8A0v7wRwEr+i7mc0xih7zMt4j
cr1HWacLvbxDzY2dxGyRHYGSEzyL3MeZhsdn4hHloOqX82poEe0jWCQJpBln
4N1GVZnNy0zQ8UNrWPa642DuuU+n9G1R2ERCCzHQWSVSLkUSg7ZkGY2g696C
Xo0hRcZhQi03suSoywz/acDKcGf9RRcid2IQchEW6PwZ+E0oOxvTtbPJW/GV
oguNjR0bJAn53l0YcM1OMRBO5WFpapCyeT3jmTvKl+LHRA4Hd0uZQ7KoptN7
Pg+nJgdxn0EFYDjjHdqNOJz4qArAsMd3BDwF5Pf8V0w28kcgx2Wbt2dDm1yi
LsEc55L/hc7RLl8ftMpm+3kI/FmoPZuNjGkJbZgELOONubWH/k5yNI1CopYl
XGn9NKy7DlqNsy2AzE9a82VMSZn3wqNZdyje+/TnEqNQBa0qxcuMIsM3ChZ6
StjEBMqW5N1C1DCUOgHioZF3UDi6wqIQwa+3dnv9h/q94m0vh2wgb5TYn0Qw
dkN4Oc21Mh1/5dk80Nto/n+wKLNud5hybhprrPgIc5GVmwrK0QQ2NHnW4BRy
HmDwe1pIf8JjfJwNIESDExHbgm56ql3ghBZkZR9Bc5aGJmXvhsylAPzbe4PS
qqiHnfyjEyFXU/TMh8LqfzGaFggNHWXbMjnnUTvPQ9gvAa4VY0R397m8CCWS
TYhz9Ae7scHg/TjrtKcKV7VpX4cxhir/azVCEfkGcRjBHNOQnJHwf4QG6xYW
CcRwwZqBV39LRZt8SHyJGeImdXKD6WOh1GYDoVAWHEvBy5y2qcPJwIeBOg98
GtZOK8ENzkzgQEA8Q8AqQTw4/QGPjAeO4cpjTUX2U5urevN4A9Fj/EGfEoGm
C8IGbE9xtBHY6Sg75b5NofSN9BCskpnaNwEgkWmkxOuQYmxmZGwM3OxxRRhg
k2075xNqmLpeKusTyCEVkfL2WrEcikXIi8uuUZTLAiXXLlZ8IFvPlMrhNO3m
+B4BQZK7MuU41Ur1SXM8qly/i45/fEz+Ge9E/uaxe0aVShftlYatqKtLoQb/
jLKIs0y52XcX54T9bOSEhkNAdmPC1UoUvC5v+kFKV2/htQgIuTZS6v0e7c9m
scO7qHYZ4RjYWjdcRpfrHdBdJ4Y6P8l3KVmfJUNrcsioQ2cyWvAJHU9nIpVZ
s9Wj37Ahg+GYCQFNcUWQc3sv8I4cQva75QM3bsVD+kOCimL9cz5gJhe5/xim
NMekGN0otw4hf4cqoxtsZqoA8NhlfaI31OH7LQBWxOH9NSWsniWVvqJvvaP5
yBARLiVfWhAxWIAnLvMGIqnyhOmxpiagyEXFWhuEPFSOxB6VOvMqKeUxFFVb
qO33yHoISPn95zfL8dYfKOJkK9pH+7N86vdP/852NXrMc7elJGIJFq+quuTG
dNVcRQ4GDBaB4E1e9x6cznSQOeeEvb+8CoUeCMXiBwItit145eFoZ10sVgGa
gb17bFv4ga9KDYwG/dyZ1jg1oRc12lrWZk050DmojnbDZvmG4g82bamYIS93
OB0UWAEIaqUOso+HguUwC8w2286QGuLxdFVjM9avfLefrgIjSxO65e+/m/xQ
mLojGSWmbkW5M8IWMH+MA0KIuI2Gt5AbcfGIONsZwnlz4NBXeAPSBPmyVdki
MfWRekBmDcSPT/D/rPx5SK/eB4/7LTpD7MxfMqLqh0NI7k6OhMXGKAuLbqc2
m+ASemDpbEljiYSBxVAPKzx2IbWaZPTRfFqO3jeFGKv1ooXFLJJeXuqwMFVQ
SAfzDCRf+BUzMcezjJqEMzGc3qcq5UiE3lU9FXNYieZ8ZXJWgfthspQmAz4b
Vq9mfimpJ41ENbyGuIKsGYtCcENRDcEXNxrtwVFQDcQmHKenI23nD6SA03SD
qJEPgna+8XjNVYE9alVr7kK+h6SQSIr5sV9UXkZkvFF0Ulnim9nX9p+a185X
yhZemAgEOBCucXpAzjloQaKzaKbSDqhsDYOCtZLHDAzO3xilKRaGYQxxP/tT
rCQ6baNUpfTt7mfV2Xmjde6S2H4B2TXZBu+aB57Q9E6DGur3dKTOge3FlOUs
vUe+Ez3H9Zhu9D/QflZZEk+Zl5NIGjWAk/Pfnbv92WKvPlEolvT6QuHPuPI/
fObu/3eEbpXChuaLpXKZ50fxhkTHbk8GJDozApv4Ojg9qqKJHuvpiM7Q0Pe7
KkPoYOZRg5nr1Dv+dH0u9oDLXEDX6iyxvGaElRaKRDXu+yYJaKmjjxf76JB5
JpMBe/7spiZJL6abZILWlOf2Z1weYtsDvK2Hffi/OKb4RdSV4j4qn8L5CbVh
1VflCjoy8pIWtjhE9sBieFDMmghfI56Y5Serk02kDLlUeJG2JJnaT9sAlkSz
xf+RUUrEF7h6pGksiA2ua4qCHfq2eFNkbMPHlnbQUzvzEoB6AXHg3ilVB6PZ
4XJofw+uXLVaRguZ3JfPG0bUUloqa9Mf9ON0cJibkyo6fP5sFHgr3lF696h1
PmgWqMCwjP7B8C4dDHDVeE+/j1S/JBXJ4rY4Z6Gjp8ahoeX8UrUftN3BjWeF
tIVXRbokqC7IlYYF7KhlMKTNNlyNukYJ8+cHQJ2VugmOEiZvL3zf/ZMhq2sc
ldyRnRgrQrJr577mB9twj4NwAKLP36RPwkM85MnxV3CQX2sB736ChkZj6UGb
SoxbMng2dPBNL0tQ1tO9D35/R1egGi8+W9NmD2hDRKEHiNDRILEg05Kmlw/m
xXqxT8QpYdsxV993yK/jumxFrXV778RQ9E72j4fK4tKzkjGI7+uOzoKdVB63
DbsQ0TM7flZWePSLWlUkl2SsRP4pk1BVVjPRwBen5wBiYHDsEUFGgvzHCjfE
0BPGmVR7PBCzSqCLvwl4orUJPUOKlSmTQgF25LVxbeXa8mHg+OKo5cXu34M+
r+6irVJ+oCB1Qb+glL94rFAW09At5i2K/oZwmNZte3vWeEMqroTAGvQdA6Vh
pBnWcG5QRwxiMRP3vuW2GxJZiCZAX7F1QXF4S162ijB6P0/uhvkIjrW1fTpw
0sF4z//dD9ur713XJI1+wc0Ds9RmI4n5qaFm83urVx1z8dBMEo0+WHx29K/6
LqST+3MjeZX4pjPMIUGK+Mr6JDAudvA4yv0Gr3c5j93x5CcSxoMEjUFRfq34
Tg7L30MNk5Odp9zhLjO6/JZAAgSd/arV9fcLhrTdlbaoftOjpUvzTd7JoGdW
j7e2z0XBhJegFtBB2LjQ3d7CL2/tM9uqkwmG17J26B7PILWcUr8fK+0c9SHh
hFuhrlbGpBjSy6oIPbFSPzJGWFcC/G/bPfCpWDnz+C0wMknlt7rp6NEw1hs9
UI5GdwTd/szNZlkz5PgkPBRCAP40z2DAps0+Wg5MomU+fX9Q6BZnWyTTZsSD
n/U0EDjtTUrhiA1qTaq5StBiVYI4sjEkwKFlPLnx63OVw4YX0GDjwURx4bRa
gsieWIY/4W0cQdwX0hGGGO6idPjZWPbZLXKehhOjkqhp9LqCzGkSDVrW/KYk
W1vSnbifqmhr4jKHg2PMQUyu8WicMflWcLfhB+aRCYtSfXbUMQ77hx3kvk10
rg1Ucrmh5XrYyl5qIZoLLwCgWofMVPortxxKDdVYhklawIwmCCP5H5eo/JbW
C742UeFVqMalA9SkKl6Y2dLd3wMaJGJAOUqiHNk1Fn8qQgF2wW5xesZCUWIz
SqrgCJA35I2TjffFnPqfejzRb7/RpBl20wWxoaczdmcSwOG5nUETUezdpdEn
NGImH3TCEvVTSJ1w46URBiQ5Zz0+z88OVfC364ZMshpFtMDNPzv2oiAW1Ip2
a7E9CBaazwBcwpowNXvn2DGDIbX/6B2EYFrqkBEZtSNdrwzwETH7ziTtUVM5
QHgHsqHUM6GlcyLq/eGiI5I1quQvIaelkaRmdzQXMDrULwrON2Vex5qD/P5Y
hCd9R5NDxKuTzQmC53NThok1SWXci/o9qFcZIyXG81MNAZ6EpOEezVAAKYsn
8EbT57cWqWlKR1hheAa5ZB8A6XYDZum1BakNv0wVJUfXOSZ7Lw1dSmrXH2Ik
tsXLjAJStdNpcV0eNexrhqANlRaPtOZ27uuJ6wjwGNdtpAWBuEkFQP1Jg5/o
NdWw+ofd14yerUk0/PVvPTBu0Yx9As4uSSeRWm0Uq4AV+Z5iZWpahZBBebqQ
XafQgmraeNAeKr/UEv7m1qLEY2u3k9xfs/Gd04nNXRXG4ATIEwMPaIKGRZbs
nC2bujmmNcMhl1YnFMl2N8CB7old5RtlZtqVY77k3saGAUU1xpsKTyX5z7PF
359EYW+Kyp4zWoAoKEox3319fwSbP1gsx9VJIFDzyYxCkmKlSXjQd+LEvgnt
AeFiaJNIK0bQFWzyNPfaZZMftjDVCDLlIVBXAEKo2OsEmlAzby3kTMT/7QfL
gz+JHH/GgLjnoKizXfXqVHqHn5rR+DTupJhRpowHNjZbt6l+OZenlnbTptWN
F/Jlhla+B4bDyMYuf9p5qJ0HqWFbFEj3ooryEAubTs96SCFGgi8s2kKOWM+R
vrvBoOWU5+7J3fudsOE9lqxxWILeJfCZki0T7apnS+ZVlH+AL2/HWxVTF3Gk
FVn1NlRdSk4+QVp+5yOpjc0FrzVlRmNzs2wjydC6jezdEGaD+Fq0qkd3+ebi
pKghajDKubm8DnHSeJO6EmbPulpfLJyLbh1bh4vj9SO4htuR50SptmF9M9V7
enru8d4h4Bo780RVzL7GL/kmKRD2JDHmUs2126ce4QOou6y06a30cyW065H6
V2t8AHfsIvVQvDU9xD3F4DrnwAURcF00BI39ahkYzH4dwqrs1gbGmBrNdAbp
hRTmO3EO3ixkHMusF9wUPecbZA7JJ+OpQKhK3wn5OUqJ2WO+BDBUO6pRUPao
UeNiX2FjXN8uHm0AbWOgRuFggxzyfaVeDFJjj6YeiXdzAARQInH4wP+X7Qnk
whV/drPW3lvjUYAMW04Ejsq1aEN7DqVXgGvsqlR/mbZkzPM+mKcjnemmh90i
0HSwWXWu71Dgq+WbBauBhQ/ITrWL407Fd/ZMH6TrwhQjmsD7ZRInUzj8OGhe
PV7t5CCFOXg7caV+QpIEdjO1XVG1JDLi5ria3Q3ddVB0A7Ruh792qPajupuq
wAZuYmb6tQ5YNYaMfjuTBfBKFVW7fXjRNrhPjkTyu+9mOOKQWVe69VrvQCA+
XHueBB9biAEY+va4kUpBcDv5lNnliqUVMNwd1wxYvW9afteVgTNnaqhgFxGC
c47IRKLRTzq3/v5TXVOGN+bHq/9MXsMAXCQn9jLvSFcLU04HzACCUqA+vHJK
qqz4uk4MCQGJVK/Yus0rwfIA4Ob6YjJdSZRCIeODdaSr+HuWD4aHkxV5b5q3
YE3DiUbWzMrgo2yWtMdQ6ZHa+SaUyEZP+B2H/gMy2zdsOxF4knxkt6Ot5GLU
vTjr6xiZX1SqCiOhxzEE7Zu05xgZdiLNZcRu2zI1V30LVR32v2MrPs6313xV
OplmtkACfzDcCkNbfFFQtkl3IfRtvQlBycNgjDb0Gd/TU2L6PAzuau5Ng1bR
Yl5XXCeWbNw8yd7ews0Kdl19zgMok8Ew81aPSsjnRWQdYcugQ6PVMKCG9LWi
oJWK57hsXlCQqkuxi1ZYis5X4VyddXwmsScFFlL6QpCdHJBQTpHVpVkKXFAA
5PgNZaNOm/z754csBZeIrtf0vC/D9DX4C6AeCclpiWLqWB7+1WPGFF6CVMbY
Kb4aALWuvblBlVhhBF1aWljnPgBjgQ5OKkpiGBbDRJPMT6ZAZtSRM1FEFb2e
Xfq4MrEGeMyMrdbfpVeALf8N5f7DU4XnqcU7O/4XrPkqeTJ1/Q7I1BWHzgfQ
0H2LIILf+RQKPxeAULTUfXnk0NkfwYca9SZdBEoNH/5exK4HraUM1Gp5qvs0
+qaA2jF+UGdIhkYxaPRySK/JMi99LMMCRUCgN8jLQPYZWIjfbAK72PD5gz+G
k5XQjAJ9B9JpyThMvNutrVWtHrzoETfZ3I2y5Bm7DGhvgXpmUJwZfcQb1MWe
hQsapPhQAgS1/2TsZ8CveZG5w84RIubVQnjY7OHBP1jPCOaD6S5KfHnSoJ/0
+wYcke/sDSItw8frq0atiDe9EyZDEPHkLpFn2Htqb5/fj+dd3A96FZbmjAnQ
93PiMQXDwrXM3tyaUq7rIw5gta4AYFTEz2mvea5u+vQqdJ1s635/AGieuoiS
rnep2XaVVyOLD4xdS4BTH8qvzwTEmJ9plqKDlP1O7tDAgOoy2mRAWVUanHpW
lZrakaJhEsSj7ugvtFqESnFAc9u3vLCXOSM0BsNOSVuh3hxf6NE5nQ+jWkHd
m9bVMvFTAnrR6Nb0gJz15SFq7RnlKIqK/SNNsGl+ehgi7G1kNU+Q7lSnfF1C
vRNILboc/N7MsemVQGMmq7aw3+Qt+7u9/ubkqUSceDJN/USWnTsZeL9Qy1V1
fTmBUoZPytEsiXzK+yoo6W9vwNPfXq//Ay6st+ia4r0SKpvHRNhE38BNWxtr
EwNeKCpvPN/eB6GHJzaKNK7MY6nln2Y4eHNtqdJGenPy3bDMYOSfj1GBfUqL
kwy60l8t7RjHtcDCXNyEkIqDCNT/DNy0m4NT/XHiCnHD/N5hoRudFcsVkCZc
Ff7R1JvG7jG3/IGZQaaqfuL1p/drLvAK0r95ccbLMyYoVvyzlUVMhyB9vpUZ
yjrsjJsobnDWJH/4i77df9qXMSneVBJQhLlzBvSf6w8PAAQ/DKAz99YikJZ5
NlRyduZ9r0/r58PlyORm6f6aDByRwo72/4i4HbpQmZu025nkdQvTxm7x8o4p
PPDCddHdrW78JV2uYoLKjkZkfEEdcSQj52SYIxcbSu023REu3RIKTys1dDm1
pqaU01vi0AxSPAVGyAalwLVDFHrvohbxF7CVidu6yp2xx9MxJkE/qkHUJYIX
p9izTvCEfjt+t3NUzj5EsqIcsCIJCPmrc0UtWansSaGXfCR6nbcAKU093vSY
y4uBibEB9ZbneJFelFjBa8j8YSv81aIzw7BPbC/rh/H/pKqQmx4f2mB5gttW
McCbvQPHX4Pv1is6UQt7fJvf2yF0JH/x71W1Z0Hk4Fsqmi8TD6lX5p4OvXhd
d6o8GbPasH9bK7lqGNwJfjj3uTFxpyqrvRMmPWNvWfiujL2zH4lxqMSKGjYa
/J1lpeW5X04hkOJ+G6++LEPigG1BguoZxXsM2T7ZdDBjlIRIq6zbu8BQdas0
M+qm20CohNd9MDnXob/68dsjvc50vneEgDoAU5pgCtRrqztvKtdUlwdFAH58
mHR+GvjqokajUKtku6/bz74Y+Wst2Kt3oVOxiWJtV+ymm/j6GZjMZ3z3HHsF
cik0MSLozEhCjZgq9110qmP8VGGfOT17EWefXO1TjcYgYjYxfq6rry62l6qe
8PlAxFYKOnqLK3RpAAZXIH5/KTfuSdnAZ6MQ9t7o8DAJ6JqlSGFSL7IXfFCu
JAvDwZwNP96UYdFf8ublCT5SMIraqRJsQUrtyAZo8VFW1H0lrIKa43oZewzB
uD76guodu/U5hFVJAN+HPlz3eeanwBj6spjQIYd4cogUEMoqStMG22yckUqR
YOX3HJ2nZuzPvgjV15kGHpVHv21T7eTILsyOLYDfQr5iL/PbqCz5ri0/Qf8t
ij/iIR2dYUADCKERiugJgPjBIxr3SjBsfJaRYKROeRrQFH/Pk4AxrvuRNOJH
2BxA8awZLPgKyk6uGq5jaiDdoyg62iHNnzzbX2/NYcD0qS5KvePLo4yDXJVt
goM/SwRQvaT93jrihqt8bqY2VyqlpoKcULnT7I1r+GYs+DMvudGv/GO/K7Ab
pFtHvhZrhIydHI9/XRlAlF/NxM6i62wuVoATOLrTNFWeKOzFGP2heM6MapgM
z9ANnYcqCzbaug11joaHHKCZnGD7DPET8kHtw/2lAzI4zEg4O+dZtI0ywnKw
1p4m+/ltIT0CmU19x7yhAa8POqHXe/xPAu47pZtnuRToa0n+P4WUUfEV6muk
lMh+fv0G7SH8WPDhTSs8QI/NqLTQuIdyYzqHUeuIZJ/LnrMHjVf6oqDYkgZb
REAXPSriURKFw2VCS6PCkDWlCETaj/taQeYtiJoA5KA+aQzAPppnW5fe1Oup
uYjFELQJQ6IdJfoSSo47Kyh1u8sRJxh/0/7keIfjhy1ixXJb3N06vM8s0RHH
A5HFgrAUnsZG85d7faM/d+ud+21Dhm7dZOTXq9uCt3e18xw64gIAcc4lc1Ia
qP40kOynrqaPSdcg101de+fHzEInLxbqSg6Y83lAus/qU9JLJAU4b9RcK0Gq
C/YfAHd4X50koQBm5xhVD5HyWE1OgvfAGR+REHV7UsZjNtPVr5Dbuw2LUJEk
fUDw89ReJ90sLl2OOyLefi41yju395bT304RVLBk+ebu73/nX5PJHkq8i9IW
b4h5bE+RM4vsKB8A5hz7KYoYn9t52hQZjfFUB8GGeaB0et6ZfKEWyWonFnc5
8kDj6Ciq5l87LZRNgXRGn9QeIfXuMFI+y2zzDgVIUyCbtCfufDWCbFLmn77b
Y2kuDflU/urkiOs+fuZr5f2/FMojvA120bt+AyKjVGwonhLvM743TgBmQV3I
VGVp/g/mwdUAdNXo1zT7ckoqQ7WHQp1ngHsiuQlfJhCx1p6M+umcQka5pwU/
BXnR7gWHitU43ws9dRvliLDQNyhIMShoacSJVkz3dXQL67Ir73+cYO6adw0N
5YXmsTpqOOTdqULpLnSnc+iiWD97rNjIjlFB1qyBE95i2q9kOnEvBWQ+bzwb
3q1Xq/Qnd8sMH56xtihS+4RtD3KXeR5jbYkiW/0oAH2J7SWyIvsb5n9E4Xeu
WTbK8eU0reV8ti6qEE96eqEHIWoPIZM6i93ea3IWKy7gM4BK6uzNnWCuyQrp
rJtAM+1/17F6j1x4CPGevYa+18mLLtcWdkQCv1nxctLpBx7b/j1SbrUvIuoa
77ITmweJwm5aZCqe2y+w3COn48fvy2UGPI0K3ohMJ31IDXsS7a4prSzw2gdj
xHpyaE2nkFeiNxCh56iFdmx2FQreMqRfI/jFGv9NblRzPUuJRzfpRf6FN8Zd
SYENPNAfKgojkHnUwuoeLmXLQK9jLIbuTScfaLpZjmD5MDfmKWVcVhFndL3R
B1kM2lC0SEmasAHJPUxF7mgTKPGrLc2Lj7gR+aIOqsJyCkENt9aHPFLqrIRn
i1zBm7S3VJUeCH34r1QwgAYSXtVQlBb9gFO7i2i5N1EnMH66wXRBD18hbcBv
O/qkON8p7sJrdI2qG+dxuvC21/Yor/QQqrDJ4M4cSBIpwnTbp3pjZmuime+K
EuqozCgzbf+LXTRc+6GSS0XlYJ9OSGGpVNPAT6IueYCJVhshlpSWAVFMhWAv
QV/Rqmf/5FlJbbzK0o/fdsAACxPKuRyNNh/b38xuczEvVFdxd2l0D+zElbmj
qnbZtDqYCbkWw34jwvmBBD4Vh72uBF7CXjur549y7bNnQnd14R1ESn7byo/i
F/CzaIEIRCDfGRINSVPfZoqvcFpDOhgjOhro6mNl8+GRAKbgEJgNYZzuttBj
N761X2NRZIazt96rpGC2kJzypxTKNmVFjkLCE1pkxo42DELxSfV/wJQWpgqU
CUyPTyuX7NS87bqNYPR5dYxmENFO7bIE0OujTqN0ELR7V8AxasUHjF3Z8Kq/
AKBIerl71YhqxA1uU/ZA/ul856Y7d7EXmM9EfU1yZS0mKNPSY1pYCI7zgKGq
shvWbqvnZc11XIR8QKKdBZAAqIAOmgu1E9F9CxPv9yute4YX2N/SNsIJbCD1
HzUtzqBhAdom+SwMpji3xYdpmUEXvRcE6IpkkhyRjANX9oGKa5DogExxXi8/
65sOWrMNoxq2srf7H/PycR9CzkjKOeYX3EEdhPJ2o8+oHLp1zJHF2ZIuSE9S
SOaCwyty2OFTM8CVbal+WDiizz7+d49xveUuFCYgKDzQYIL89uFC7Nl3errT
Dr+D44jVmnAch1z0o1ygJBI5vrN1UAZlu/Vct+m86QDkJFtC9r0SvECa+IFp
kl7xmatwDg/hPY9wT6F6b/TK5ymzwTuNripsle7s88IInTeKeAfbmd+4Xr7Y
hme4oWQC8QFmd5HZCkd+8iS8gW2vVfYDcOO6EUa6LMdCQxln+ye2uuJDocnr
yq8sXd1BzSKn0iu61TIeB7aBmCGV1foXc3Hy5Ks94xP9z3vnWD6DGGJAGUoG
IbsLt9ePpA+uQ3QpFgU6GLnDheA5oNnM2qqDOWo5dcPprxh2rcD44CzPDLfL
+YTFS54DUBgNaWQqtIgiHk3ge/n5zY3Lsj6FtplZxFByLezeZjKzOUvlI5wA
eqpd075EtOoHuCh0d2d+Tldai4QVBtwg86mjo7cGlppkw+/QJg3x5Jnj7GiC
HLjhRiSWh0nphV+oOBC1Q65/yxrwfVVdljfd8dE34IwIBGzRMbNuoMxV2Bt3
qIdd++BEI/tkhKACK9aNKB5ARUqI295f5zRgDxoRV9h/vx992q0Qm9+057uS
z6y5bsZaKyszHCGWcM3ibKCG4Y75wR0839s71Hbl3yF2RUmNMe+SI++RNYYV
qRAoHzGieEmc3fw0hqjAdIgioZscCc176mQ5LOaF1lYtRduTIkwVAXzrr2Wy
aqL4u5dwJR0mm2Pr36jYKh/LJsrKBv2sAhZWnOOCN89imafS/ULs5od60Y7v
psmwihUpZEN0wLhIz2CARHpmD7xFz9YkaG4fCCwWoY2GobYCqt0htDHjqazB
4jvJB7LjjdCfSLqm/JfLwfEeN3ZBoTXxNc4s+m8pxX1zyzBg5maH5c/nppvn
lpRXby1d7yL5+y9otW+dem5nXfNW/u2WrJSHuwOuY5VcG4A5zEhpbk8r91kW
nGFpeSd84iIzp7SdOBbgYn8MtUtw+/hdkkutJG6PN2Susb8DYm3m3bWKroqP
HUvrNCjfMd1HO3T3NkwUmcVsfX8hRUHG9//fdO3EVziVIOdzoKGBLuQ8GbwQ
2rsIwow4jig/UE1Y+gdcRgbnlLGMOGOtIQ3hrmyf5EiM+jjEQLUUYlgx0pk0
zkaVLGHehNypL2o/TIr5kMSyjextbrInH2uw4qDUTLu/qQPvhSNtd3w9tMGM
e6RDgSSmbVWNS7IOKQa2deWhlsMvOv763YhtpFsvr1CzCC1izYKXoAI79KrU
CcLj0HDOZulLGK8Jk+WbTcaI306ZI0Od1xSZDR5ySZqn6eK9UxtnOiL3BgdU
MNKrx1sRSSHW7BklS+6PILzXQj3hYdqqPQ7tvIwOn3S/4mtPed0fb+TtmNQ8
6ZugpDuqWj5ZLp/SE1lLTJWtza9JBmglXHKDBU8aDri5zvU1cRJbiT3DmA+s
xvUd8Kv0g+ADR7r61Oqo9nAhzJ1MzWqd3UtIcs1I8ZTBmxUa85cUsLppPR7d
2J3RNUL219boPPYNrNknBHDl5lF9RBOR4E3MRr6vPzTvLVBpdEQI5Rl7ebzr
jhWOUCnqLiWUeV0Siqn94Zi+REhxWuND630pwoegTOh9pviz6dDTKnXY3AAf
CVYZmMAmzYG0XJN3FZ6kD3ys0gGKmy1OoHWZceeXKQUP1CvFOvk9hLU1mjVO
nYZtbMWCOxavNI3pp5IuaGemc5AbY8+GVoWvxRNO6cVJn+3LBxcoC8Yt4yom
rtV9Yhc4QQ+H+hF4OBxyofFgGvSWaeWyC+oQ3AqVQJtddkzcseZmGBYljgaT
VU6MvsklE6dscCu7mnwL843v9ORRAjCP2YWKGuy+QyaXGsLNUfHEWB0mvDlL
fks0FmBPjCArrb3UjwRY8V8QLbqY8i7LDulL8NdBPfRyOk1d9vWNB8LQQzm5
8Zporxf17XAWGssD0Ci4+9D26OeHjMVX24c/9+VpanzZgbaUX6MWtyuBhGdW
fvSy2yVmtXQ8BeZKsb5pipkZee8lsWUnbxmKQYKzgiONIpCiEkau/6ReOCt9
b83ByhYHRLIeWjR1GbYY9V2XrN3629GuFLf15x+sFTLoVXQ3NKM4jNpj2bnJ
gMwuZOzeh1iH7WvS0eSLvyEGVzc+sDniUN3UCc1Hcvr2WL9YJpoVv51gbAWt
gPn+uvts6A0Q3JDJyezfoHVAkoe7rt3IcLrO0mVw7h8J1PC6yYONSkiKNH3V
iN03Oxok2RzKixxqt0+Mk/9xV4O2Y/CyqZZ9ApRuuE+D2HpRu5qwDi1/9to5
jHWbg31T8AJdTlJmb/57oCmoO4aOCiO+p6ruDxMfYmIZ8wq67CCirqpyBODu
roBTJZw+EQ0QeMnxi3L6jgKZElRVupTrS+tJdM7dCqtRtpzsihSAv70W5gw8
jVDtzPKJ+WWPeJjiribBG9QMAx9juLth+UeI+r4MrXBRyoKVF590S9FKcz6t
lJiFVu+dNeuZFsGNUu1Y062hIiHHFIt/8gAn0CysYIBPKWEVP4vUwmDFE/VY
1lO7TkFFp0j+Oh6qx93D/4KwXYzu/t32v3lcumZmsGtwzP8TVPrwdzkR6OUb
rzlfE86GY2LUgdKzE0+Te4Rblqm1hOnGRHpzY/gQYttO/F9ub82MEc6f2Dkm
5SqI0cUwUN1r0yUDdv1GHJOa1eNgjHJC8Pog84ni9mf6HekKVjIm1EqcuDOW
dOtOlqOOycslHCUcAPzoxW686A5ZpPJaVNmNbOpofZB1cnVoTq8E58cs1WnH
xAUx4PiNfmomb7a3P49YMuSXzu+ShO+5BIihntmQKau7D+wH1X+TFs4Qu9Md
7VnwNSgM/VaHp/Qixq9ykCgKjATz876w3dLcdtNLsn5o+JjgPPtywiYAa7/K
7QKbE61h43sbhBVzXCJLjhtTXCy1bOpMMFCK3MibczknD+pKEQyL626GMLLQ
jFbH8IMCm8g5VKtIJaZk8W8UdrGTTUfdG76M8gu31MPDQmyyNp64IM7AZP0O
rZs2U8gtZy3Z2ydZPPzJjiyxae1IguMZVmePjgPonHysa3X7f/nckiaf7x4t
+1xxW3DwnFcM5TLnA7X9ld50T/rxHPNT1/0aukFMSdeCC9cerZebXPETIwkT
lc5GETHuCH0nPWAAGPB4SD0sRFoS6lQBfc81ilhcoNXcDyO3bzVXsX4O8EbD
ftPGpzJRqHgh1H7GPggVZLCB2Jl8nsK5Nmf4a+PU68vvrPihOOtLy0G0UjbX
uBNXq9ZWP2wKijYsRbKg6A+cOvnPFpzGPHPG/VuNsls4BI1QAFjDxpAEf4Nh
zj9xMacmbuYWzLic3dI2ITDLtmn+usSyezWQ7PRWWMER3/31M63ADruAOEgX
9BXLZ1dn2cau6kxi8LLE7YWH2OVC8/CGKFMQHOApk6G7yg/9kxfuQ7VMqcgr
CjWQdIPxAIr8DOhiBuCNmr+Y+oLrfIo84whVv43nemXfLB5g5BpXh1JEA/sk
8Pdu5qXHN2P8Z4gpL/aciWlkuU9kS4D1T4VqhqFNOs4utVFz8fR8uovSnCQX
xE0g960N03GZCqWOr/qNMZ6TRwY0ADk+4h0FgCw7kgVJ1/sX946PiZ/yeKFm
CUiIANawSrVLyfxJQH91iPkwh3odZPy/EqxrPY4cbuVrFDkFUPtpfMF7kofM
EFkOAU2XAucZZmaH5wrHtPaLZw94Axk2tW204d/LPCYtE2SJ/V53D7aApFrx
0F4Irbi/U6qtidUWA6okjUMh8icuxGgElaIK5oLpELLggeOEPoQ/mk+bpkiy
hV+Jp2VeILU0s3RPRw4VPTT4d7Jal3zEbsy5G4v6ibyTTrJ85+dLuneWxN/p
3ElUecepXJAM179XTlmFgQPxNb6Eolo0xj1KiqG1RuKazarDRtn2Dalh8L+y
x0ULpohvQW7ixJAcb5dcYOkTMCEyelDnWWANiOdAZcHGeNsMIR1NLVf3rhDV
x9f4KZK76hkJL/P1zQzv6siAoyvPYTUSJiG0AcLq2spCG8eZWZt4je3gKMKi
to8/gOnlIo0WbBD+9MbAu51ues+sIMk5IgHkFFoT8unWZeB7hB3wpMIWPakv
tU2oRNVT0bj9SLFX/sCTT1ZCB1wV5ZfGgonnLONv/O5EizoyKu5AUGTgAabq
YzxFvR+x5DNBWOeiCbcBExCmnjbeyBeqlPN8vAUvpIDOBUNQCNDrjQ3NYTc0
Qpds+QZ6vH2xI8goZDQlwYQm7sjwxNTNWeSmYTrMtjELQjiSR5H4kjjUA4MM
s8g/GL9F/dxqwtfpDN7LweQF+FkilAlAPMB93w6IUiDyapmMJZ6W3hTc4SJT
mvnn2gjD9lloNmTHkvYRbPsTRoxJ3e+57gWd/srm6iyWLIOS0zMug8SS6svh
bUOp1VdIek8n7lzvGprofVr/rDuIpun4ah4TNNtcGm8/Uhmi3XPKPeaxrhM6
6/xs2/RZo/lFmIJ27EuRqKDb6IBhIl1TVolpH5i+k0jC2C0ONEkXoEHBVSLf
53lnWhwtVWXVJPEPt+a+oyK1To6s8raqG8DFwDbY3se/QOrHQpxuBftoaq7A
uMTvR3n3o5tb+12X5BO9tTk99zJnmMZ3K+OQ3eSaMcdCyBwcIjAxYv2UwBXP
+4+ksdEuEe9hXltRIu6Pg838wjzdrBP1QIDrQhbFKCXh9v8CS8IrMYVZ9XlT
xssJKvgSrh3waj92H3LBfsK2o8wMa/gj7/bt0jcGjEV0bVG/5J/n9gQpHx1a
OHhNbj/9N16YkuAOVNWrhvJYa1R3CmohN5VaDeIDIFCRkAdp+p7eHBAK8KOE
1Mx7e+lN5Qxwf/hRzHK0bMRMGmDB0qYcLpiA8+Do5dRgFHnj6mawbCqIYz7F
s8UxDHwVXDf455U/A8lz510mly5d2Z/6vXFCPw61D57gXG+3wQtxoRgTw/a4
abdCpYiS+Ze1RoJ+p3Gvbuos5RIAjRy5tdTQABxye2WazF1qM9Hequww/hsG
BzWpXXVo5GgENLQKYhCTn7N7pXgy3pt28t1qcVYjhtd4itURVtOfnwF1D85j
V1kzdZg2hyx5Bq3IHXARKhlRDDo6dSVy29XWwgvEMoF2/O7ih7CNhEIknVSS
v67wuEOG/cwcSNiHnF+zJjcg19VDxbL1NCzTelO6yzkdRJYt1lBC3XDVmfLJ
GcD+4ZBSRBHh3JM3nqVQ0AphpEgL1Jrf7UQ8pOVx27PetKChXHqbiQR9iqQX
PuWtBpzt+hozhnCqRSa+VgDCwgx5gM4nEAubrfCYChF+Iqyr051iuzLz1d7n
oHb2NRs9Mp94bzuccic6aFEDPley95/oIPo52OCn1S8Xztsb4Nqzu4gZfId3
KXRvpkJcKpGU0HrcJjymlRs8uyJK+QCkVfZOhrrEVn9CrN5yGM9h1lquuEtt
0XofBaWr9iRWAV2IxJCM9m6T0qFns93zjc6iZMsY1bX0IqZONGM7eoslHPyP
vWj+vvVOTibxMWZhPsc3B5wWBAq1a+n7XBOln/TmougHwPnLySNwkkCajkK1
bOc+YsC2EY8OPhPPjohaEAYv3pOpi7h3pMAPHnVov9sybw1ZWYNl3WiYdOp8
/7aYhVl9pMh99JHxiFZxy3KbgnleoASWrYJrqQmgSWCRZ8HKipN2nKOEMeR0
D1xWzcWCuXyDePFJPJhYcNeeo39dtG+D9Ly/8q8xS5uIe6gqokN1i2IvlypR
TT7nnQMnXgQTavySQ0t18ExBQAuob9XPri8SQsECwEOHTLVnlL24kCNSUmQA
c73Vh/6cacK1OYb/lyhOsyiQtNVyAhcGp2urPKAjvKGU7d/muLNiA0ox2tD9
btbOLohuNVi722HP/BRFxIaHwnOcdgv7hI8cDI7MZWQup7SQQbS9X9b+HfQu
ja44TK8/LYzhplhvvMb/vMbAmcIVi/tvGk03NYvhxxy+DZnKJPMffmT74uBX
SiSGfHNwEiYXw7S5pvWmRgbXu0PXNLPGpnTFy5reaP3K5TW6jLcLzEuD0D5f
YvJt4NWR6PqidbkbRdJ1DOaIo1XVthEYO/S10L+cyU9AvKilOdaOwvvZzNF6
tPB/ObJvNGplkqiNMXYrYj/PlC9/ubGQha+inW7ugLzE8y8DYJFR/pZFvo0C
PKIMsVniiAd+jd0pt8Y+nxfPdLXuDN3rucuuMJd9NrXitwnYvDhka7iG9wNk
rp8K8yy5KSz+k7OBa2AJW/VTZ8ytZ6sGc9Cae0mxxOX7Rx1YwY6gl/7gjJL0
9o4BapWCz2LokCn2n4KKbRzEp9BS5PGo999dRBu3+HjlaurXIkwHO6g6Is6y
nXL8q9jSpR4qCCWwTGp7iRET9aRXJHV9mMXBxvdO/oVbURlRDEs1JhggUZYY
ScjjCYAEaSpv6hTqaomGQ1xNZhM3+pzTZOftT/Ty+6C066igiBAC8ryxeUXR
V+sk7r8lQYvA2hTjR49OEdWyVnPH2SyD8gqYqlEI04QB222llngjaOn6Pq/R
D85i0AKNtmzeAALJfsSe/8suouqWmt8MzF3m1w8G6KVwHQ5kJPBurtR9WFSF
5snoFbRK3YXPLBb9xRMIIC3pKPm2dC8+GqBfxbOESqRVaKlm+D4ugGn8rjDN
H8MYIq6ce/lMeAixTkow2M4BF5tUf6oeq/gz4Ex2Gzyu/K76+bj8hjcyl9nt
EFHkpF7/5Dl6C009/VLHJnVEEMWkuRPoz0byBX1jZPQPfBhRBtfAvoNQpzs4
OnQ/NpozhX/VsYtG2PdttVvfEmd4rNl+eUNMMxfUg+wL5nCkFMA8eSSZYkNe
/Xd1Tghnrpua2ynLmPLCwuNnTkDXkdgLo92Mf3AjDtPmZFcHM1OQvM1Sqkhq
k5lfbuLmy5MEhtAm5miBj55Xhe1AXLkN99zB3y+di9IIxetFbq8dMPj7Aell
Hh6F0Wexx2adaLdTdp1o3aBp6Mlf5fEVqvM4oN4gskzAukvM3eHK+TRuiI9R
Bzv5QnvBW5OKTh44/Be03RQlhvYv15LBoyiwfF+eDNOVE79K2E8dLdbS1IZ2
K8wFDYc/4vx82x2q1HCSVKM3eNt5bw6dMSrSIoc2kPyiQI+NTNBF1EYeG8Ie
Oj3B/arWVh5r0IiI9mJ9rJILf5szI0/jQa8fY3GL6Jj+QohNBfO6lFfHRFCh
bBiQgvf9gwR+6kM9SjyKJ+ixgrp8sw0BSW939OSk+RxYw0NfX5YyIMuEB4Ss
k59ppPJvnPh4RTUlxiN/n7Hp4vrv9m/CIifdlsS2PxPADQ+EI2UU+I4Hthc6
/L4GsljqCA/4f1/GTEy70cuvHxtQPtb9sXbx9bwJ9Z6D9YBLiyd9/nYFXKHk
eSiNHk85kpt8AE6jR4fA07fD3dLgJKcWRg/FAEFxZ6Hd8U8oZjFzwuLCxZAh
Mw11TpdUI3DFmuAmF1MDrxIqUjPcB3eqPAux4vO9vfPgP4t2TyxfcDbfMWJP
SrJeKRUUBM3Vh3ahhdNSBH+/o54qPdjx+UN9MdebwKg2fmqOrw9MjWwLRLis
M5AiXeZTSo48sKFTE5QdiYocAoLDYG+Rnozi+2qlSdOxIychVgu7NXRZeGiV
FG2XVuSky7nDwAryLd7kgEFbw8A0wU2ETWc1fBgCTvTrxH3sJLAWz04TiWub
g6bCndtjDdFrSW5KAOJIktmj7XZML7hsvrA656mRcBo4pojuIo47xoSB43kX
7K3HgRukst6h2xZeDbRl5kEhT6ArkVGdPubxoeghDt6tcxjavvTXs2ItnEbR
iXqYWuVoMFW8NlUtuM7bDWW5BAkcQ7UBuTzL3QF0vM7cOhUpB/loqIjX1Ypb
8D+/vl/Ay3Tn5ZQyk8CsTcg5wdLWZ4H6GxfU/Tpv6I8TIU3O4YgmCQo6sEqt
57HdauJsrpj31wvrBqQnKr+p4pSTpZZHKpVV+7c6bQuzelrdrVqbG4S/T+lT
nCsHgYFodqRKhVifgXn63nbjZP0jUNONIbgA5Ku7hNIUBb4RRygKCJ/6bezb
C7AZFTu62ap4M/EGSHBoIludotpCxxaOOcGJQI6oBOgP8hIr31HWmZ+SdHix
xmjuaWN+VF9oUAPj9zVqWLuMjIsO7oJmgReIYKbMvBhXwKoVSHT63sZIR31e
ZUOyQz7UlZcHClVJYLt1a1dhn3k6Vsbsio4zSl8Fv63Jw6o78LbVYLe8PFv7
dfbi/QV6qHv3xOU2gT4tedlY0os6II1Q59vvKBhmE5LnXQa4Fmd95ATHnGqu
Sly2eIsobUqGqXT+V8BenkoQB37rzrahtHuJK1GXFYmMtLUQwx20Fkgf/lXw
oyCiRdnnn+458d87poxRcIQwwUceM3IFzmrSvDMMD2QQcSfnG6uPHVLerWOm
OsDj19bdseDLv7QnrG3tgIdLK3Mh/RvrS++le3i0rlZWmG5pd6UZLLa2u7ba
Rnsec5ZQcwxPhCpm2pUB6Tje02c9lfL8/SmHlrasyC2uchXv73HptJUhACbH
+lKp5jBOtzJowOR4m7lsxzfDREeXV/jYBNV9NQNqok6wABrbSZqfMby/SMLH
Ph15t2in+5JDdBeCLmFnQ6ItvBUGLh+y5AWnoskiZTSxqY+N9jcbuQpHRLPm
S1DMJbpusZR74fnIAdM4plFOCaBy5XVj6H8yyqYMYuXY1WIYQHXmSGDYXnSM
XGuIDFXc5D5MXzzQLikHseUhoTfI3B8EBFO4Jg/or8A55W4tUIMth+rtgKBB
APgCnYn0zpeTbr5XSiqXDaqY+9+Bu0Ks8nQMEK950sEBYCSvrNnn3YMCfsGI
v3XfPPCEGO0czQrM3x42DhMXZ6BkG4wvxq/hEM//AShjZu6f2l8UMsmqVpii
J/aSxKwibxFzMeQ28bfU8EwrCPM3YriRWjBLTG1bcr62oAaJBlT/6z6gxozE
gQE4lt9cJSPwHyAePindEyuqVOvr4njSelJ1dWGKnTNseV53sjHOnBsRmu86
3+meUAJnvcDwQIZnc6m8a61RSKWvm/JVF+gpauJ7nWnpg/N12RXEyLpvosKC
SE0XEpJ0G9tQahNN/9ALp5KYThl/QHv9BngXHkfRttYt3DqIiNYDvToOZO0u
WTspzzQBz9ycBCu4tE4gD61eBZJ5Ic6rE+ayfZbHU1h1hLombtagKk/jwp1d
3iOfEeTfDbxV278XZvJa3/uyzSnmkfFcZ38UBHbJLczJpO/bhFmVi5AzdP2L
oI4Ge7lPONMceW/BSMJeRvkV3bjprNqDI+jvXQH7SKdpvBm5HHKJrpFX0j1L
wEqycFZP+jE+rsdHGe9SZoeo0K3BOIeFTKreSk78nKYgu1IdfcbtjtMxC6yH
aKkAPtrseM5zLkYDRGJ1RRnkcXUWGR8IvG7NAjTxS3nHh7f1gtBhEh3LBWJi
QUk5fsAowqWZoIw5V1/nEqoGN3UpPFizXMpKUdA2wcLSTSOuy5s66OxqnU7Z
bOQrVfb/klcP3kmUlYBEeDkoXXMoNIf5qFHrgWt1eIRuudJSRUDJRpZBiQUM
jv4AY4s91RMLjPv41tTTwOkVYXkeVV6Swv8eyfVaUq2/0Gll8FCbHf6UBlnd
rltC1N/WjTwdpQmkPHCDO6S9Gj1pYR0wG4dcGaE8bNmfjWy138cVRdCmHmQP
R8NsDkM392sehEiZmKFAyKGLsQWJ96MQfMANaqvKJEF7B/Eh9V0Q0NXuuiVp
iTZ1DfaRD7bJmF4cJ7smZZTtpkPfWJw5KfWljCA/3Ol3rNefIZMUnpYhFivh
LA+GGbbYjVfhKOYeSrVuIwWFiGT8TmDu5mxklWrjDCTIU3uo/H0tjEtMM49A
fdFEZRcWDqCaTXKG63m9SM4vP6SqqZ8z1SFL26IRyX/Olkh6NorFJ0axysaK
0KCjDgwqXgs+BrZSCB6Xr929uxwGVFoidQKjQgVUGxpqdkRwafn3oYCiQQyr
seWVzVC4HZ3bkNbVdNtcKGPxEw1gkZnGLG7I6zs2QKhuNwRqqHG/vWI4mrZQ
AgUksPfvgxL9/3lj29dWpxb5yJgi/w+KpwJao0Lw2Kex0qwbPg4omHEeUf4p
9dKnutgh/L4cshl1F2rhVATCcTdD5GtRavPYWoJ+/JLDeuEce7KIrsNH8RHF
Yds2Wz15NV8oL50MjQtWcvQHBS40dPlEVyWge17XOOH+oyUYU/dPHGmfhBRY
P+t2E5dBy54gEKxncqw/E96tMDl6SqDb8IU427HFl32AzptD2PeFaIv2qY6d
zn4K9keHzSRlO4PGMiTgGjmiaFYrZCM+wyyQBFcApYJn05QpizREqadxMP5m
D1nQqjaYnhDo9ELQdhGY+N8EoZQKVzcA46QPtoj+VsFeJbP/lh5fKbCzL89r
+/56nk8sTMzppqyK+ZTizcP2M0zGARDxd7y3Rv41GbAx/0zTTHn9FXNwgr/n
HMIT4mTC1MYn1rV7fmhA1E4A+jqltmzl9HwprBBd3cfxNdIaFsR44Fw4iV74
y8ulZTsz8Kx0O5YbGwroTyLMTznExqL/BbOTguXYqX2UOaBPBfSoGiHNGY0q
4dAFL8uoYl9Hs9beMGzzY1+UPdhixINu58a2M4thj09/wetsrh7dONaCjkmv
RxpAp/2dUJcBDu9m8zycz5C35YzqF2G1uX2dqYz7nR7kTo9xzofQEt1z7bnf
i2Kr6woqwwTTjYgus3OeBv4g8NMsFMwDa6dHdUP6g1uosrR6tfsxMxa5QZcH
j4fX9y+200n5eUynCWSu7c78T6FPMh6YKhZK+kxA4/vbiBBToTUgRS57tJgy
5BGRn6hcBDELBfsy4V6wlUN0Hy5gGMnTHYIHKGj3vBZ3tnGvf4gqA8nPEAJ5
giJCx+stGXuhw+IyP2Z5nvuzdcxiBTLERXiCXOfWOm5QuMEcTuVo8mocEtm5
xMXLj7o3BgR+qmADrT1dUVSR3/LBnzOzOkZHS4DmmwysfwR87+im7oeHolea
PUu7SOFJ+abWsXslgO1VkVojDDUzUGJG63t9gZaoqLvlxNxs6932ST4PzvHo
ICY50yDun4uTdnH1ynqD23Rf7AfmIWibwuz7Zw5EzNmpD4Irc5/1DkZl6s39
8FkkbJgfy6M3U7Fe2+S+56eQ70pNUinqzzeomdaYOxsJBngkWju2VNlMpWLa
xOn3YOntHRZyQNrbsEZ8XToR01oJ5xovAUBFs0PJuDs9YNax9Od3qSt90Caf
Pb25cMB53SDiTyKftm3o7kkGa3bwktDKf6r95OumrCnp5bAX6T568d/odLxM
6XNsdQOp1IoLElw7RjtRRzMNlFvXN2PycsjQXWeU0fAB/S02UwfAO/VHjzyb
q0jZu/g7WCeTJT3YkQcCLrfp9K9LnjYFAe0SQe71ah8hopZMWrNYSVepE3D6
P6fR6kgahWs0mJbF17gQHjSNsyKbbM6rHIph3eWoS2tbmJ+8iXvs3nvPhq9V
ZdREILNANyB7as6oQq3mMT4N3gseR0qC7TLGJWjzA1Y0ZGPE0VpXh2w3XhLt
ygHHEKbfFDxYjG2CiRlt7YRL+c89BLB/cLmi98pGBlKNhV1Zn++if8oiiGFc
tZbdhhKLdAI9fJL6+FDrIlqYzbBApwhwYDVS4VpgxxgY2AzInpCTAakGDMMB
osXWo65fSESQ3FBm+TQSpE39ElOtAi3xGVd3E9KB5iVqOMQ43CAx/LEZY0jf
6ZbUV5sBZXga+cljX6OiGRajKsx916uxU3+jBPdQOCrMbQN6CSRsDdmA3woJ
yT5PIa46Oi6MzwBFjzCVQY4GSXtXExq6IJuBHtI5TW8d2KHZ0tB8MI3GJVMt
vJ2rviROvA1or/hde4xEXG8bduh7xj0nRVMmSQDCTCt33cfH/E1Zbd5DkQkL
t0STPDDmsH0joDiVUD1zCsz5rutZlRaSGckElc7p1R9+YmYtBbsn02mlbgPN
DWR91U9KHTGwFu/5bdM0Tfls9nVlKGmT+XPmCiJ9zhwAykO7ATWwKMxlFPnh
468T9PU7RbYde7eqZT80CLXRE++xIUCtn2koEgSY7lSNB8Z/z0APZWKqxOeH
MJJSp3FNToebJnCWvp1mFwOdYESwfBXMrRRH+h0nuvd6zNKbs5SwrmEqPDu6
C4nDXdPU915A/XuMr3D/ALprWXo18+uAGLTPDPk7LwQzkqTmwXn+nmAPx0ff
H+f39ZnL/F2hn9wxObeSVotANvYvA/U8Q1xJMr3H82OBixhf0sWjr14905NB
2enKRVflMknibKq3xrcLwJVxjWTTQlJx739c5JiddB4KPyi/0hQKgLPo0kaK
EUiO66GrKiuNHz9O8NIP82hM6pEH5slGyK/ip+GauKDMmNsi1cYi2vw0a+NA
LPlTYfloNJ2uQp1uPEgvcbZKicO1YNR18syswZ6hjShCDKTkbhuwsMx+fgsY
9SXyB6n5ZwycWaPM02jU23hxphi98uQJjsDVTFbp8qjinTA1DwGGB0gsx+qk
X16MErNTkJenaOELIuh8ynOv4XojKkqCkydIs7IP1F4+gwwRM+/LAOqq/mCl
/XDUN4A2zdLNFGaKfB0awFttPsKTeV6yUmFKLLfUupa1y2nFDK1cQNs96R5h
6fUxepnWAxygeuyjyHBSbJzhEwMECOlNrsdu4EC18eurtw3Ho8Kc33WRHm5x
LIHTDlACZXwZ3w11kWalXDbfJ69nnx7GAeG2ATplGc9Ek/HjAkSxH9reHpsc
wewdi09lha74AVXCOJP6UgwFdMyjeRzCISBTrbe1YttPKZd1sUqsmcmco/Sb
UHa0Lo5IJtWxYdGjIYtubnGRx8f8v4jzfPYSFN0V1pbrnzV+Cl4DJBc8+Rhc
Pf1y3tXm9veDIZ2Q39Zj2zTjKSFje0u6UtdTmodP58yzHvELn1B92lHX2zZs
MaK1RiID/4t3K16GSx0geSZwkmu1bRNw78rTdEsblrilrPQYFG+CJXB2gwLA
WloQd2Pmf6PaVATBKVU3N89OQ19ehDWvDTcgc36Cd8Lf8vM7qqtVGgMH+XE1
G0dNHhJN3WKWL/l+VBigIlRh9HbImA/xGmYYQgq3fsCZj5uj8a1Vb0ZQZCh/
6w8l5QDKt6wL4r7Y1XtQrbKaz7G6AY4vMfX0pcooPAZGPajosy0nlGcg91UC
XoFqKZwTT4LNbNGUyElKbpECxRj5lfUndDPk5b/L849I1thAoL25z38yqAQ9
ggzapSbSaEYRZAB+rI29xNly2jrB3O/Mg0+w5NNwPSjrKw6E69LIZqO7WNKn
zYFjLkSnyRj8QXMXRRiTckOSKu+1H+12Etw2p3O8R1ZM77cODvGWmtufTL61
yGnU+xxT7M6TOQShFbhFHGIzobqIQv0skScQnjDHF9VumX0d+UOnRivKzvcw
6XKWppwJgqqIoZeYlZazgIKCSUEU7dwgnANDkGXDnwsMXXGxSWayageEeqrl
xzI07Fb74+ktpo733yl+hTuckW+biQKlJb2XYAJDUcjh4a9qV3Tnl2ePO173
68k0Mk41W7B1cxeVnuXNWbnmdjLjb21aa6olWDJa/F2mgBXUv1fnpturhkNz
44IL/U5vRQ8BMwj1c/IbLYcVHAGGSPM1+zfYA+ehd8Rcy3aviLCvH1G5jSdx
Fr21/oFlHVMCwVg9p4udU+FIh/v8JnqmBWudkFYtQrc3BoWzFE1xFokQrrfs
UMhcJtk9b/iuq7gONrOpu4gY7Kqm6ruxfXWAiKCX96tCTp5/+C2/NIRWtJS2
ps9/3+RROf9wjBpbrBnBqUbxUZhbYlbd0reorano7WW1zcopKXbqBUEgqulE
00PXNwjDrajKr2Yzh742YEtuOVyOC6Zhtc9niOE003Up9Nux6cfhenVqT35a
yXO5HtiydFj6u0mFJin4KtXbomo74WltL0nJIlXWsTt/TbFWEQPmSAYY3RFV
3t8vx87ugtZ3sRI6Fma92EKLB5+xAzJJp+LlZRd4HOTAkDGJWOcJ5Yiv7P3g
OnaGvnQkII6Y0p+hNjobt+h5OsXSBYaUdBfdB55JkmSksKGa3jjj6qSmtkdN
hlSq/nbduH1DsTVyO795IPGb2DtLJssENL12NByCujo0vMpx+bNQxA6tK69q
RYYqV7lFYwTt7vzDQEwseqxdZcbuC5R31VPxFGx5U/K9YlKauBtuwhJTQ8q6
i7WrHeoa+1mEFwG8pHrQ5l0jdIRShxa3qEmLWBx19OWQBTapk4W4EAZ2KkJp
cxOE5fMFEv862klletd48K+MJ2F2q1R/rk7SK9n/LMxbOHrPycwQIBSXAL4G
Sj2+8yoiPe7DHxJjBbY+niUQ7vLPAOZD4e8ceSKvJ0wGkoql5J0Lp7Z6M4P5
ucwSipfmWqhfVX5weOx27SyPZrzU37ZjbPKAjZOH6aetulmahBEkrAhLlMAp
la/DhiFAgnXwwEq+9zejMNShS2uRuYTp6k14HGC1Gy1Xkx8cgWfnscRK3t2p
6NxQmPaYZ8jSiRdJh1WI7o+2lX24Bwwz6fyA8oS3K6hOwfQ3J+ieb25px9QO
d2eotdfhphchpscycWJHeAgZ+PAT2xF/SmMxat5h0jpWFKA7eFuAFJ421L/L
1rp6YWaHm8kl0Rm4nZMXfMLbGdGkR+l3L0X0lrIg8MVBiQvUpzpUOJjo84J1
2zz+WTH1Yg4zleuO0ee6z1p9SVCuf24Ev6ybR0x88nHcT7UI/hKyrIRRowR2
Iyp70JBSJxOrwKsx/0zRm2oGGU+b8TNFoVp0FYzSYCg7yx9hEAQ87HpTkAb5
C5iLX+59YdOixAax7r5FzIXNqzCl060OEC5J4a8MWlD2GZCSROkeJOt/7J2U
r0NcNR/oaNqztegHnVXCUbtpir/hKegY4plgsLpshHaVv/Mr7WV8eBqtuJXm
clva6tO7TX6Sh5nZSMFAb0hBlZfASY2NDvEiQz5HFyTJYTzNciPHE9ouRC2f
0Hb6v/UxhT+GzeUTBjF7JJlzfwWJxHxgBzKk8mtAYZcmaPTjU6eCdujyqFds
xxEdOuoAwqoy3bCoxqJUI3tQ40xWiQcepKhjakBqPi7tis0aJo7uZamM4Ifn
mXKD0QANZc/jqKdgiHoU1R1K3qR7TBeEUllvQ2agYT83zm3b1iSruN80ejtA
w9m0I2IaNTYjWJE7NVYNDmTENoixfLImaUlAhB0JbKtntp5kjC6c7SQVoGtS
60RFoC2N6MCCw4Re/xBOnANCRn/KwYNPnHptM1VWboILMLtncAMTugMibjY2
/9H4Co1Ert6EpsZ7pIOhGLFGJNtAtH8hIzQ1ViR5fhhNVWuPsEI43fMjKmf3
o7OIgTX6Pv30Fn5O9nVWbfx0tz5djfSi02ZoqA7n8O05mqEGaT+C4EtFqfut
lmeKqOVRIbKz+2ESvdPPiho5fLbEGpnfv84d8nBaEpA79Bu6pUPMuyUh8Ez4
0EeYVFi2kjbhiaypuf9sG7IXSLEhHB/R+5cyBFhgAF29U5AO9LToB52VZ6A1
G3/GQyhvgCLMmupstah/gQD7vKLVlscZ0Tf3tvymp+XmcrZQcAs/j4WFkKMG
IPI+Vy5o1ypL6n8gM3jTw9QHL75/3bmNfkZWgBEdD/JhbF7UxhFI2Wi5a9zu
d6gG6sU7zDesYO0qB6Ggq8pMan38JVfUHCDbO/ONF6kTCvS9P7K69pi8hP71
y0b41QjWF8P0FQfzR3GxZ5hvcdKsNvKM7z7Xcs68YsU+EAWDLx0XmPmjRG92
mi0DXVsTdmEjxIzxrntt6wMRd0Ea8S8i7RgHURVzr7plMvqtoW3Sdl2zipEW
r84tQgIu6H8PsGSai9NGoUeo/YNWfj8CS1Isz+5Ac1JaSBr33nU+vVp7G2KZ
W/DlRWLzlmnEn8n7r6oo3k8HSjS6Qfz05iFTaDk6iS/cHxvZgg9t1jsvtweO
buFv1PvBSkBJlNSfsMKhYiVFJsIXAuyosH5GNpReRvvsa3Tl5SIIJo21zYiL
xNrJ6iGxtuSF/+XysCxLAySEHRkUGzi5sOZFfmPH04q4nw/CA4TVnCOV3fvo
E1fYCqfi7SoXJXvcc90MONQhc+Jhnug1XUToeE5cyVNdYdiW92o/Z1e9pUWn
ldFYYtoJAbTLBlESg0TTFtpzHtrTE7aanj8Zho8fH7UbBUQ6FH83XBXcay0y
e5NY7PZNRH9KbCTtnScaMCz2CDSkF4tm0DMdFmWhAA/iERCtaOyrA1A1zt1P
VVjx+MxpxCXcYuMMBXmDaGUAwXfmMsnKmR6asG4XQlnbJoU5fmqrx9tvgDKI
6ISMAwQZPUtEkFuq9t9SnOM2/xwP8uoR2PDHoVtJ/LLCMOkIxwj9CV9EQh0f
WYMBGBU7hBysuMHAksXkrlqbSgP6k8m31LTF89CO7T/zN/waLamjD8uMvsX+
VXtbIN7pU8lxLnbvZWyojrRO1P84mVkLUvPXWnlHluDVutvDM/K+hTsLMfco
RbyrKOKO3vLQ4Vkqh6/G/caHEmHdyVEnQT3X8HUGNVEV/WvhZiMUs2B4vjyy
wqYnSbIQhKuNZI299FOQ/IxqNSjoqiJ49ejb1KBgA0xfgdp+GiMsXgFzoaJa
3Iw3iMJ6gmBLPMM6taHbVVLTJV7ocRBCTlY7hXUrAXUckjGWokZEYsgM5nsU
AujVd/9Tvfli7bEvPDFPvTrL5xCL7ovfAlWbOA4VrmKrjxY/UIblHjr4nx81
2crgQ6qE0xNGjM6aTftVt15AORMZta6QW005kgpyxjp0Nmq0GRNVYFt6g7tf
lLGqcPxqw0XkcrLCjoXwsSH2hdq146p47isM5+8PT5UBjaAUuSbsG5K8K/tE
bUoacejR8Vy1YY+wgugKnQDnsJTRps1tVkcq2i+YP1sY7xMxMx27L1efsvs/
K262Z7aFeDz5NyUFX+IK5/Nb9hRlACqIKz/rFFytWpGnCylpgUBl3JSj41ff
197ryhBrcb7K0nAtWClquTlHqMDoyBbU5hdQqz8ZrvumOaw54PqwLwSQZGqU
QgHf5UdivEI6qzL4VUHB6X3frb5OLrYxzeMdT699klAvciTQTlkGnKeYAdAr
qumSuf/OOAZj1/9xu0juoq0R4hkIcCxeJy2AamW224w8gxx2Kzu2UJw1U0v4
7YHHN2v7ODQ0/rLGxTyTn9d5/jlnkxGjBnCQGektWBa98TuOBAmQcuDAe3RZ
vDy1gxbesAawNOrYvfw0YWjTylSb/wk/ZHixikIC9LP+mhvbEuyHbRNJv8do
RUyokm/aXH1fYXP1geFuG0xRYjHL/lk2f05p38g2QwhoY7hgizsA7k8QCFpp
aAFma8DzUySo2N/plrfGBQvVwYDY0gybjW7MMrZy3CgG2rDnlBeI0Xwv3V2p
ma8asSBeFSrNdUsYQ9IudQ1O5K6FZwr4bj08/vZ3+naVE/AMuw5bIUIAZWAb
K2nw32Z3CU/rwha3CgFBkveFM1xJqISVgWFVkHnypaecuYzgoP19awXR1swC
ofrXjCUz7GSjWJbC5BNiABw0TfwtyuKMm1NRbhNjOT83dYKBDhiZviGOGecD
dEVBZMNNnw5ZzTIaLU8Ldwje6cwO6BT5lm+sQ/5bSoTb/lTFgbElKJVUhAk9
hIKc7c8zfgytq7nO9P7bhJ9OD1D6K2hin/iTIT2/7b+rc3aaoHOC/MBgrgER
MomWuHlbL//dG2ANBuS3vcBFf5qa9R2KCgB0sXZQZUsWt/8he4O/R9HfjLkM
btkIYYQdeSADfCPxUF30t/bXn1k7L7xKHCWCoIax9ytGNunqKr9SZ7FRNZ91
AOPFHWydauCBmYG8PPKftQd5HLJvlDdPEfvmVtWNoHKG2mD9EsYzW8dMLbDt
cyTwRaEsD9O2Z9Znkq7tfkMsWm7T8oiw0T+5lDdgNjhA8CDTNZR4UsT6f1kl
dUzi9Eo89fiVJGXQuVLDqgzgMphskvV3mZHUqVROJRL6Kv6tgOL/Uo5TIa2H
2WLK3Xys6z/3Vb1ev8Me4poMwZh1rmjmE5/mUuEnEfg9ybEiNEB3yrmXWq9u
PRCWFL0rq6XK5GVJPGtjNPB+lVmsODymxbR8WHuB+ptoJsKxfJDNxF9Z6i3i
zyHd8pfRaJOB2FTTbVDxCtaRMm89wOjSBdvul0jCd3qp/407830Eoc1hXjPg
1UYg8Qt5nhMaQHEHJWJ26tDgh3w/8UkMJJpM8EE73ZAiZyBVn1+GRo8YHxv8
zjjv//SFCTpj9rtlV54GMOAe9VvQq5pivlObnCz1JxkhiT2OThALlEsD/cfV
d0UzochzffBKaJrr2AYJ3MzJdXmoLPpiwFbtEklCIZaYtZCDakDhJb1Foit9
OHRn9g15dqNYMDedtmPTLrS6Ae8GQhbuGbazDrVChmrMGdTFwkQT1mr6e7Qp
XSt9F90Ie9ST8hFBRmwM8LKOj8D4j7nHOFJ1RLiDqJN4LpwkksWCcE90FMb/
OlrW03oKvaM2l8UeowxoDnAwEobocNYPDT0Uu5Tf4v2DZrFe9QHfCKcQjVd9
IPLtrmHH4adg8jBzJb9eIBQ2XR40IVN8K9il2mrdIbe7FOzUaY8iA5aF5g0I
F3N1dEQIKJiqE1f4gA243iucaFSwogjyVP0u2MYljeNBAtX4fPfRWqw/13MG
39v2Xy2PibQ8hLl0YvMhEaV0MNOD8IeGQMD9uLY9Xa0Em+NrH0F2kbtUuuaQ
TqcrXncqbWFpqF9k6ZsdEqdr/Uny/QPaR+TUwDwnX03JItUVK/mZpt3UDorX
XIXkqep9EPTOu9sPzp27ObbpGHelXkSGfOg8VwLfysOQErdrya3Km9aQPG0H
4fnsjm2/JqiSinQwCg2kCUzZel/YpLwGcztXhw44y3HjBLxRYWvxEljNuQ/M
Eh9s8xWHo6KCXiW/0TtKwtmEst78Q9kmvB1uTBc9L5V8EYOv9d1To0D392Yn
bCWwzv5GsF5voO/q2xxRM+vxYXoNsxP5qLyiK4RE+6p+anhoYpK+HXixn084
iRjdtPgitXjKuBdm0a2AhchpYp4Jd+adMD6l9HYrSzlBQznD9jLyroFFdYpC
rzfX/nYjFcT5omC9/VIlKU6plykl359lChbV3bVum2zGgoXaSyBM5mX2/TVn
Goa9wVTHOTkrQBneXe0Wb3TqFg7/eoxLQ8DFdebUX84zVDPVak/V9Uze7XUr
XBJEv05T5Xto2KkP1pDRpc3Seb//T7xEfYAJHCaD6OwGECcPNoyaRAfUbNoS
dKsbl9GeS6HFpWYyyba0RzaY0RMNktwpv5QIAOz10CGYmBYFgZeCBIWTkEIP
SzQpUxEX6kCLjMCIMWB4T+AoVgW2p7IlHmdM6t6c3bYHdxPCLjK9jGQhqDKz
aDaa3/RI6R5lL4LRXTXiYZnHTKNwOTuNHl08URLKTWfKZ2MeBGTquFJ0H3EK
lcRZWZYnopN+T6w8M5GKM1GmXoA8CNYLKPoO9t9RAcA7SZZaaW4uLqxymFLu
eOTPlLuMwFAJRHrVNOdeEixVGpnyCYvq1FCNJPr0s1rVwRhv5w3RywhwJ+dP
omtHFyys6b14lfwGcLZqoog9C/Ei1PSfhVBIF0I87wCofa6LLpNGvx6vxMaO
K0GNEpmO1vJm3wqF62bRBkyrggmZEOUm3PEj02Wyots+70K/S6YzJqdUlkOQ
LGY4zXJDUkZpM9Sa0ZrdaiSOpFW2Kt3AtNYrtQmiY9Jyr11L4Hhe8JqXtmNk
uDa0hL3e5nv3bC2a4duYWNdDuB7q4bs/4tFpO3FDLkDYBLBg0Q4YVFIcJQlZ
kbO/WmofuoVgmSq7zMftz1RTwOcyYkKgKHMVe/Xa5C5x373gxLlYcN3pjhxV
KrVpsfHl2Ef4T9wPEFxn7S7nkVnSba6CbGfRlhOiVZbvIw7bDZY3lrf1/ShK
JBKs2pwkUeywC9KNiFOzkmYZYC7dTtob4c3ckggBFKXBK2X5VPZx6N/Uw0Vg
WXLL8iaRA3JNkVBtXEZkt62vj3h0jZ5Eoj5m17xxnGbzH+BDrKh1npsfYqaV
aRp+KYWKi+EHtd+LsGil7efPzITT8F3IsFFcYn4tTCwutZbVFFbNSwju0X/X
zbfEoPCok7/LXlBrjR2U/8CVjgkFB4OrXf/c+jUkzq1qwEDm4kZJ73jcMVZP
7WO/7h4WTE/A23DMGPj1xb/2ZFWLwU+xefbFgOkp5lqDwEnLWW7UFyc1X89J
h1r+SQI7347JVpUwr4CeXyBuY81dExmz8CO1cDmnRvNGh8bdm+Ztx3eUQYUn
kM7nl2mia4US+2z5ZFjxLgdhMJQ+COV6fZgvraTY2bc7hT5Wjj7QoACEknMy
yyfPrgykiYPAiWIgnqt+op9uM6kADL+TPYPYiWRxLBCrJfcHmKGo0qmiUCAK
joBfJ66rpKmmSvh66QMvO9miUm3k/Z+/wj1Rf3iIeFsXOwMHrFA7PfIobHm4
jjZeRVHSmkNUT/QTgjgVq+x2RGOXmI6UrHJy8O8JdDrPKv1WeBpi7UcK4K69
I9pPsgYDCpZS2iFJ/6RLHYH4SEWD+yuRzM24Dg3BnkZpLig09JDwKDsGxAyY
ioE74HRObFni3H/jCk7nYPBxiLaFNehsU6s5XD7MpfE8UwuIn12drDKLYNKE
f7TNzVDgO9kcLro64oiExJxYlwO31ER4YOVIL176pBlX/p6TsaXLVKtw6FY+
yRmJDF9CEo7WSMkh6Nsd071VHS+hU0HkFzIKd66KsB58+A5kgrwNw48UefVL
3boFRLq5cvjahcNb2A6+cnMiW2ReK9CCbnb4SD5JUsmCHjoNbyXAq+LROLV+
8WQ4TWCZuXm2bqNh0oddLmF6n3K7L3h+K8mS3x1Iuia6PQo0EFu07olYMh4R
k5eXYeBeKr9JKBy2U2JpQvvTvUthOS2GI7H5uSS/mjH5GiemY/Jj/GMjQlzg
dEjeXsan5Hj43y4Oh0t95IVpaMHhqTnEdNqSk/4KrYEcjk7rEueSvi6hdHkM
mAg+/hSPifBp/wzdxU46+WNbC3thaXQlJwjBgs+h3355OtSFUzzyVg+FeLOw
tLrLYypQkxn+nAs0VuiKz18hw9iyeeYd80vgWgkoxT9WI5Hs+6YkNCS9zQfq
RDgXHK7WSfiQiEa34SqC8HHVWK2BIymYWea8olFBRec3/HbezKYtW5qiRqoJ
vzgzUedSve5e1srJXA+Y4ZhXfzjxFOA+Lx6RkN9rn0QBhVbap5cXzWmKrVRX
VbbJG5pNUqp2cBK8EGRPWOlRLUmqsQIAQOix8+a2+2An6CTqxb6lLVzoW0d7
q2L55Ylbur/M0vx48jHxXydllyfPzTqkQC/fCMZF8CgsW8T7F0bcreiEofsO
R/EgeFaPqQWDQhyXBtxrPIILLBWCI4S1O2Cq4xUnE3iSwIfeVTY0pndKkcHx
4XugyHlqMyCliM8h9xOvVcVFW5C4sazXB8CDfwwgcALWEG3lD9hF8kGQBqlP
HnOke1A1qfVA6iFCgf9R4H+Qa8xRbGKXYzQg7gW0nMTqnRaVsWYwmjrgBvnz
gC8AbsDd7C+WW3ME5JcecrGVaz63B3zp9bg6sJuQPKg4t1RuvIMWCWWYgCOY
kNSoWkFuT7uwHC0xBMKNDAFSI47fBpO1pKredx3rnsBpdemIBfU8QPjE9hRn
y4Q4ZmuEKkq69GX8Q4zuyuZtIVX440vH9UFJWwx9GeN/TPT/7Rvb6vGHuqUW
uHNu02sSqKsIfGGsofGwYkrK5jGvG7ujD6WgVnX1PuPOnnGj4YzlHZdSCdtj
cUAHAbHxmEP6ww8YcDjJGgshXPfjW4i8so/tqf/+22+JqMyqmHfS6CsSKUJE
VasKzEw4jmbKPuiZ/v69Vp1C6nA7+X/BNV7RtwAeoTiN2k82GpPgZakIeEjH
C50TdypqNworYBf8WfJD5QrSxP/xGfDSVM3jS7Rt8NomOnAPuUsscgIoCpPy
5BdL2MQBN6D7YqXAUqDKwYpkGCcrYfYPHAl1UADpOyY5KBdW5pdA7I/7O3n5
a35O851izoZaH/31oFBhoBBTkwvSVRdlEhy9aVeA1WOMGGErfLLi6twgthL0
nA3t80XTziZ/VZRlsyOOUvF8XBryJRf0Fi13Nr6AOZpVzG7OOd0yQ8ds5lKy
Ox0QIyppwdp8Iy4bq3uZfkeDMfdQKZR1RuCmeinYhVH/hFye7CsfkifEtFUB
1M0QBntJr/ExGrFyfMw7i0/DsZqMlMipJvZDQ2UpbP1nYGHziLGcPiVZmL/H
kb/aI4owIeu2+2mSC2LUg/7xi/nnefSoFBwRBQ4UjA8kQ+nQCvwPan7OC6AP
gaiCV/KbY0CwpRU9CD7Nn6hdh7rCYgfm66etDX5oZ4dmSJcZLetgB/9zUOXq
w60fiauHOD8rRJkW0W5ujd4pt2kMbE8xMvgNvUr6fsFVCONyD41+45QjI83W
HtuNP/C7ULV5L7lsyl78y5cqT3uuTDhdtbIJzFjD+BC2FoIx9kNC01la8JZo
jHGaar7hCnLZOmjMGpF4beh2lV1HvCWSExYjKSy4BIP2WB77VBIHTzpnfn5x
26CHhTUtAhKf7C1yxwOG6RmKvEjw3kN/wbbhKTNLA1tt1uEuOxYNvaX7Q8KB
XfNGTHVXOJLCWNYfySy1H+eCNK62vyOyOHlilzcpq3eEXAQOrKzxxw9CzCPs
j22ZHSOsNl8cjzaMTor9NfGrLwt68BG2VoUa54bJFBXgqn/6sSvdV5he+frW
Cxp16uSAxxjX+cMVUx358TIanok2NV1D/swx8EeNdmjlcmSy0YsPYsss0oTL
47OpCFRDKkuZdzn6vORQDxAsO5UpoemcLm/meI/WI5ZhXc7eD0BV9BeW34Oy
JFOi2E1Jhdquymg8KE1w7//H76O1bHw20sviO6z7L6NgWhSbfjpaUIfNhKmm
M/+D6dTNd4wcuuNyQRtZqVXFfR433P48HihBdpS5llJenu8SoZIAw/HzEn8C
7mZfmDnL7g/tQ0F/q5Dbx4zFwj0ZWBO1+D6ar7859SF+Y2mu55EytoOlqpfk
s6pmwLT4OPj/D9IXVOJjkMEeJgCX0e8XVcnIVTpCC2q6MRwoz3KaNtM/ND1p
U9cfbCCSdAdAqkfzW8VtZ0S2zS6WPila4i1MbzE+HN+q5JpB3uk+OSk2kgCh
kkESGA1dX5N7LWuL7mSYVKcj0n3Q/R9mA2GhqNH6NoYXcJ6KMMUMDeC51zJg
AVlcfsOFKVIoc64ahnIOzgG9J74idQLElrDMlwFmMXE3tGZwZkLDvU86sNlP
W6SF8IDcfibFj4+9EpQUkkYobJd4Vd0565hpL7f3tilsf4FuFtFXiOfzuPS5
jerqg5PfOKnD5Lve59rCubTfYjtMEFBOKnM9kFNJE+umV3wxd0r+1p3GIidb
dy7SvGzm3ZdTvrbxOMoRgYNzSjan1oI1yJVNN2/Mixasn1VE6hUdXrQEyTNm
lHP95cbmxpoTRFl32YuRm4uSm7GEFzMBJdMQFW9rxmGXL2GQYOFV5UI1XLP1
RHLHeK4jb/ag+UU82fZ6sBFNH6ascEmebjpKSWiMR34ioWviqyta0TO0t4OI
YsHOtHJSgHb0lau+PLPGF9E6N944tD+bDZK+huwe+E6vtCeluUz44iBoXmFo
FojIxf071faY+8ar5BqNhplCPGfr/9XPra2wO4xnfXvMpQaLP7hVnLsgx7B4
yIuxEHCeImHO54B+UEjRvrASi1N4a2gITAS2C6yzAD7LZdNw9T33SonIfdnO
Lgx3zVBFw5ItG/KaRRCFKeL68hQX98jfo3wlzz1F685ywRGQX8sHDuFNDc7W
VMt258pJdbqAHQSvEL1aLhoHbNFeUVTw6ZnXvdq9Yn2CPd87RAsKlIy0rs+e
oY4OIndX4hBcd+PYXRa68Fu9uV/D4jvs5Hsb1UNPebLtxZA5kCA0AzStsQIY
wXAMBV6y6hmOkrgI7+HYXULxlc9WYuCbo6XBUTBUKRRBfOitnIRERJAFgDFp
gmrXoLHJVdtS6on/NDfo2BmKXh4l0Ger1MXgmASDZowzCeXLuIygB9jrLJAm
QSM/TpV5NoPZkK1Ea7mL8Y+IFJ40auQEgFHPWIMvOx1qytb/Rdl/cV0XIZwa
d3tiIpJGihCGMBZRMyVSU2aRS9p9HxajTwCGDznSQovz5Jwnu4/HtYEUCbI3
aPDFCofR0trSv2NnDcrbztesqckLrJPz16Laef9DoEYHvC90G6NmpY1GJvoG
x+T8p5ruMt5nUgzAHbTh/D+hUaQ+CnpadXgoHP4x0O7cVXni90lqbPiXp17z
dCLpko9X1j4hE4ifN1bKfW+kbGN7dDN8X3ilyuee3E6lPw/LKphs28PnqIpr
OWTUV0VHFxpxxKOP/Wtqzn/EA94n74FT7tNFT+cjSAJ12D+Hd9fit4CFRoFM
qqtM/pRRLrfXNdUC3rS/Ahndxx4GosRRcGvzYWtodafv7bXGXElgXeZo2mKb
gByBGtTTxOLHq4bUyka8xNne6aZyc5DrnuW+K2jiXPlGmm95SmAmLURAwGZ3
FjOMkejr1pFZpNmfGtwGIueot2uqkr0iRCO8qRO41VVvZzQcoE5YQtfRlrQA
htdJeuyTODmsSCwfJ9V/c/d79D+ifmu0gosWFBIGrQvXpU0wJJo5pRPtsCXx
omGN48SY6PEzERdJoNP+AaMgHVlYjEbv34v5frFFqYiXDj9nrB/C5pjTH/Zj
/5ZKnhbeZNBBHJrMvPeGLeSDM3u4cyoZ/0kEubPLD1RQJEY0c8PjMAAWZKIe
aKnlxbAp0zuK86mCu9BckTlhBvgiG43OUjWNUyQx4cc5PGW6D70bSfWufmwM
PzzpS43mdiMC2iVHN0X7wVLraUsW7xvTyhW8bZulAWNzvjKnQzHDa0pAylhT
WNL7TnkyE1l1FBrnNSPuVBwekkRAOz3v18HP9AbFXMv6Kv3EQHNmlIrIB8xd
nUAOvU3AJ0VNSi0g7a6WrJHiinSBZsEbopVhfNXwHYk1FbmRzOjq2nxsM6BH
6jmTmRAe5wPKOmEu8PD338v+T4XzBaRWZku7dkuasNPXt9TOv6geQBHlml5K
cEMWayrtWVpOkMP6tJheyFgepIWrvDJJMMMFaPtYGs6FKEVT3OyUrq+YlUIY
X59fQebOWaHCGxqQPtbPan8quiFxoT98OsMSgKL/RHLhigqkkpmNFX83Lu8b
CqirmDrK0UfV7J3kTYbPhUvgx9UJWeYtCVzk9JYwxfaVsnOUgBTO7vU3eOu7
8lBnsrGaUGjkxayJw1SjUpkMf75zq6yvQXW17BCXXpJzzmdNao6rqByOcIud
YFmh9vvubMlUKBGPG+KGcWbc8wSYXag12bwKNKXRORnYqrSDsVCvQ2Mki/0r
QWDuFVjj6JvUSjdyUo54WRw7U0zi5IAotU3Xq2KWKI03xYGgVA5IIh0tDXl5
FcXkjDDZx+61ij9QKAVOFE4FxeuRper4grXvANnPTFyTOslxfHRQ2SOrn6UG
IlcUW9RZj8qwzkueHmGY9JjK512ec/fwNURr/Fq5OjT6LovytLzJOGyjDQqa
y5V8xTcQMeqQe3Kz1gQC3Ve1Z+AmQ8OMYw97zO5L+28GoJ7aqVpxmxCWM3Ba
4AAuQCRM7Xwbub/mjSHoZ3yRx0SR5s6eTPUF7E7ZPnD1prNM1Jax7MTDNyyn
zJ1GSkiEeU+xVSfygUs31kg9KL3lvSk5z9q0ESaNXZRR9JSqJwUPH3yCKw1A
oPP2v52uzFYVYMrrg0nmkYxO53slpF0dLQ0TrcUAsDdTDzQTrFopfr5yHrJo
syLtG+zYfFuCA8klbcQzFc9iOqrdUtwlu1wl/flByc/PKbH3P31La33RatWs
64KQuD9z+7q4JtzQKMW88Dhdw+gesxKfcckyZtpfgdaOvbfVZO0Ti7ky/rsu
5t9B4jLgnqtD2NCkLtAoRld1BhKMKKwA7PSCpNScJaGsKJGHoTD9rhS+f3ws
5rotC8UvSRLGKuI1PqN0Tr3mCgNIS05LCHDO9W1ifcz0eCidZsF/VrguYpTS
4Tc2Wa6mmX1MizdKvQ0sPhFl7eXjCCkb1/CT0Pyb1GfANmDWh9GgQS+ypQCB
41N9vDLaxm3eHDspwX4oeZzWktttpszU5QO8MWa24FtW6LxUci9BGG0mMRs0
PSbHDQ4gn4mVUPeucNugmCv8dWhw77Sjgm3LT4bkWnirLUCRC3niWegwaJ6C
JFbzJLA8zKt9bKUnyx3Bob65wJL5VEbfmOnBFThw6YedleOJk2yqqku3CpS7
lnPTaRVodpoYisc0uwIOFeXwGTXhYrzBLjchNoPIIXFG22Q8XVG2mM+vhQYi
FStuT1njIBPJGMMzjg0TAoIGQV+SV1mLOhd+ZDr+1WDFj4ikPnGPo7curFOM
S54B9yvw2S9JnjOqThqVwvEcsmtfJ9UMR8EsH7uuLPN8Od4sKXMVP02JcvNH
qVI2jW//wZhs6dYq2Sn0z21MtZ4xaLwUmuLPG1NW9QbypPcXiC0CKPVCYUQL
XEsl7PiPyCHQDZVbA9JSCyUIu70Pa1VjHWXZnG9ZhRxwf6cSp9VqJNzJvK1X
rhdyZNgaWOO3wYXSWApYSk0sPuRDBqGpqT8aDEBUpf8vYe0eWC6+4zei38Ok
cbFUsoOBYDaYGNOx7sUE1THPWM8vLuyYFOrfmW9rvpv7+HKW+3TegQHtdR+k
hdgD6z5mTEvG5AHLHkpR2eRuk55fAFz8LfrILpLc+7CY42pnMjNb98DiKlJY
QXDNlf59UdL1nWsKH5tEJ/KYimDScOf26pJc86cbl65eJIB8OFtBhjtnVo1E
BMTTUux0+Pygwzeo86iovlDTVLYAvd1qfNl8VCepgRzjwxZBHk5Rqq8VxeX4
dFvJ7XCv1TYbPzKu2no2wqD3LomDfYPyV7RJOlJSd/PLFUrgJ3eRVGhmud8v
YPxeoZMgiB95bKRoErCHJ3A4gJxUSacNgzaVaj5EAGS9xA6LaA5oWSTGTjcl
NpEYAEyASMoRHrTrY32Xah/Uh1LoxlHdsJC/2YzqCG5NWiwAZ/vldDkT1IKw
eZw+TihTe6+oYKm7LymbGBgsRE49wMg/fjVnyae6rIEIJmISbadyrL0+H4NT
idORYOP0k6zx7aF499mcnbFVdnuzEhtYgEWxZelzwS+P6AgpL1+RfxuYpSzM
Ms0OedMv/6A10SN6Fh02mo7cbqgUct22Veh3OjkSRoGzVHB30I5uBq3RJstl
3W9tvsPS84ICUdChYBHn6ahnhQ7YlHrmpgqxKBHEoGWjuwrj8nPLHH2xV/gL
3OwPV2uSfnSuMTW8WH8djAE4pVaBMw1C/HMjANrFLroVIT+4IyVmxtL2Yw3B
o2sToEmefV/bBK2s6VPRWpPoNRlA26Fn+m42e+gkGUPaN4gTAd3BclW88hoE
+JgLtoXbPCrdl6V3FnGtQETT2jBDjpxAxvHDp+0dNZTmheUSy7joMEFywlRS
MEz2s3BUyEIv7uzwmg8k0jGbjqZJ6hxzVSCrgUQ8HFyFL1ZgGCWnUnr3j5N0
jPrVmaMRH+WE+hwiHB0A4xXEr35zH6/F+xDB+VLEwqQ1hIMjJA0xrzok4fde
Jjc3zHpT4yuaTsSlVG3iLAjLpG8lxAK50l0Cyw8khPj2zHeVW2O3dJn7YlEu
VvEvock8FX0rKazyqRdbgYFmPfZ1y1p4FSzwCKhOh+7GiRldjbDvPR5VFOnY
qTH2wA5a+QJnd2uNunn1tDaVG94zTcVsmBShosjsHva2sJM82rwdKmwPLODj
/PLmv/Ifmu9jfLtC0XfIcWedzuLob6c0ARWlFYKnHUjF0DhyJFZjOWXKnmre
JWl7YIbBvPYTxxGPFbYhBAFnzySQUmTgnQuhidZ9QHMSYZEjgR41i2d4dsJf
5w3hpgp0hTHwcbAI5r0DLgo86Ox1ZPYlI2SaM7LIcH4Gi0YCL8om8IvIdf1Y
v5h7qjGWbqBxD8bxxvvMY/tDDn9qP+owQCLa+WJpKfOQWGu+lrjK/SpINFa9
bjv7JE3coVYRoPNuWeNDPA+KsFZODELdziJ2TgZFd2aNvOaoU1zXfJje2L2N
BOgMZb1wu3BB7vVP53aWu9Up+oCB6D+1cwgH9NVtNTxfCWYboB4nDIbDb4XE
f7UQ1Pvnn7RKybolpiLatJDjJbmBDjOEM+qgixicxvyGKE5sSU67eKcLflgo
nK/1AMuLIPAix+taQwO1qJE2FKvDfUZdKBbSiQpJB3leAZ/ADFxwfK8h4dT2
hi+R5fjs87x2F0UmAFcVnXe+FaXm41Lh7CO5aRbkH5iGvMhXCWCFEgcK3FUv
Jkv1A8J1+kop0/NfL03Z4hPT2boP2GxutCQDf/3C4DmI0WnrO9y14zqSc19b
0SATYt8pL0rmmGKxadUbzcNGwQdL8LA5j+xjrQW6noJpsJuoUIrY83kAJ6nr
01gUIpb+FhC9uzQGGQmHNfAWE7i14asmkeNNqPmCoZfyUnFAa8VN6nPXow2M
zhz0GiTQ5ChvV6qZJ6fJrXnS5H42zoWDg/S4z6nsswnM3b5cg2HxYK6qqh77
yRRnu8Wfp28aZyHUDd+kPkXMLmF6r/Su80Q8MgrE7ary0MWIEEDjZ06iQ9ZQ
3NuXwAWkCd5MLsR0Eh23lROWc+v2wOoY2d67y7sc1/cDbNDXJo3S/8CGjxjV
2B33FM33yHzkbBVjSw7JX0a4M9TDtdRRKw39wTS287NL//mACc04c7fTvCl0
nHLVYLUuHGWa2kXRYUNGxqo3Pviv8x4t6PPHZGn/yXINiAMDCypX3/MMEFGV
WkOn9S8jW1D0Z91aEEvNB3qT8LIoeEc0Nc34lXMs2PzH9sdlzMRarxXXozfQ
5pdyYOoBmXmpBqV2fb798crb0tEWjFt9EGGOm67wb1hJFR3gS1SJkiXLcpcd
RvFzdKeioOieNcRoX4RTp+y8+/Wo/ynmnbbupVYZ4yQEbju9fVmkKJs9vAei
RjK2t/DqXpr1eqoJGofDOFeHiDl1T03wUttGo4UYj/ZKJmr5akXCh/qaC8Ks
A1Ra1tttk9cze9Srqwr+CeOXCPXMSKUbS38JiFxrGjUeh55qwvrkOaPgTXSk
ygynUf1Nt1yYvu1cfnAcGEuDRqEoDCcRGDyMpXqW4zB19P03D2Ql8aTPWKdz
pG0n1Ss/zn1k1XfLfr1yUOM0bjLsFeBPWRvHUWdSMXhueW852e5wyieEQ4OG
Jlu8/ouJRBwHHpV1SS4BP0PDddTaIZyHEGmWpO8fz+LBvdxyrS19axQ1gyzD
DrJCew1FhAlTaJE27d2fh0TxEZZT0X6sgoKKtiWVIGt9j5JbaUyvSeT+/1Ad
IHe0B+l6wn2oRWrXt+iJZLIlOypJDQ6g+DxXmgLPOPzH7mCXVQI+BiHXaiVy
99CcohdYN6QCgBaQ84ngyhhWBS9RFc0xyUoHOZTG31h+pW99kuokBBbDJFXb
6O0d/zSJY8nVfTdyloJ4k4L9ISMuxYVHZZPymi4sf0Vl1w5r0g3af5vC+CaO
VdINGoX7IckaRe/8cXiWLiQEPcuAU2iG77CmkqaDsxXHkClEHudRa5iCrMDG
OCsfFjqDc+nXmyEZrHhOQLCVjwArxjikBeEqzFf0aH2kQnsuwjrVQmCyyn5L
E+Ujk7Mdnnh87bPx53S5FFZKO/AaxIveJjBGCf2sUgpJu00HHp+1d4d9JJoK
FQTcdGXwTiHXBFOvlNhYBMHgfX8LgeZTjQa93ZNAol6iQdve2F3u23giKSa3
ZEM2sztsblKrv8LDhVLLWzplkKwb7VaV6j58jIpkHMQ9VhxBlAK/DDjdczrt
ywtevJXRhlLwxndBo0+jBDhgdGBQAllhRpGKil7mKqanyrDVgPijNHU5I8QT
ud1+x3Q6CICZa7T1/mExnZrfGyOQRhtRvUCJaXdze43q4PIVCsz9yZO6HMVv
Ot4qYEf7r0ApphOSR4362gUqd0t2Xf6m0W4Zs8sdA5eQcGHycy3YWVQFIR+G
Q5Jm8qLn10QrzhDkzB1EoXbSZRjc8854F1fLaQdlTfZTiq5uBc5hHLYp2Mgr
KPvtR5DBhF2nkel/Urnx2CsWvJ9Hz8nBRmDtStD/0rftuyjGtt3Hk2kw3h7d
im46w0lmwW7DiMn8uzdstqucFkQb3m9lfP83UVpxDbDkif1Kz2E9SK15Fq9h
QpMlvN6HCvKB9rUpfh7l3WmR7OCIJsTQsg/EPrUIDT1wCXzHvHkxAhuIKbKX
gMdRbDPXR2JiLTm1MOn8oyZgIQOfMPAZXywmwyrhmtvX5Zcy9b/IzDJkHLmT
+LMU5jJB/1rLD1bkhbUAUpbMhgH7hO2zxmQ1up3BM3xWjyt5ITGv65tf8j7v
nGyUH8cq8oBf6MPtN6yP+8Mg/BXMvK5d8kY4dQe+teQOmjSfaFSDxpOfm5fS
DT6QWglsdolax72Q0FTXR18V7Pr8LAEESxGfQTZz3iXTbhmo4jRjiuvYRwww
d8J+ruzTqGocHZIM785FaKzIBzMcKfGzH+PWELCnxKgqMPX3KqJHx6j1iHS/
UOHXrbkQX5fhRFXE7JwExhYw5R6vxOw/QxHht4h1GuzNaR+uIOcy5edg9SE2
cwZWrTpA6F0RMOswxIS6em+aXsfmMwHKXt0h5GCCeFweIUw02S4ow/XMjcUs
mTiG1CWNuIv+MSGBSkIZ73+b+oQq/XnKAxKqAH0CK1B3Uy4n9VCm99947qTg
vSSCuuIt2hIma/kTXTp08gBxmKRUUsr/7VnWQnRnxe4dwufCJGrnEQOMeTq9
cRbMDs9cJltBAw9MAlEn4eJwkTwp/qj7PFYyGVVnZhMYY0qzeuPXeGc3awgi
Poam7QTQs9olml1D1IjipWYK/90GelfjWHq5iDvxTj8afZmFx7X5ouogFoAk
sBEDH6gaQd9mv9iwS6QRDkxdvgu3tCV5bLbyu/+TV2mEjcFP7bDmDYKBj8NE
+veb+lM6JtE78fwhSyxbLKhSgKwIy2jbJ5f9wBGjgIE7EhZy6bGXPOsBjmg0
qKl2/35s0MmgZK6DNpRigKxrEKLvzkS63+g8Zltc0pLUPnItLbikSs8L3EeT
feqB1HIiJNWsWplQNxGW2IMkYFM44ECFYAaJiys4wPpkPU+UNqPGa4DVMJZ8
K25H8WJLoJFdXAmU4CMrWc/RxkUjtA/FipxWqQHSM8plfD1qoNH+Qd/CUTHf
um1wJ2/HwYssixwYd7x2cqWCQbAb7ZasH0OcA3suXzwS1wHJgUOnLJz3iQHk
r5heeGADKpUufSV6BkAlhBjI96bcoGI2oGYYx5EDd9fqKdnHVG9KecFMZfQq
ymG5c/JSB8lcANj8671gsFLgw1HK884IBu5WKJ2WuCTSXZqsx0BsojBQ2f+7
ZZntumMenTSj2jGey+5rAq17tBAvARzyByFuNgL6gPbehMwF9M32j7tvymI0
FQWGPO40+GVOYwSX2zoDGrxxAe5+WESGGG0/aNYaj5Toq/1Lh4NpF12lvpDt
BnRZywXu3y51z4wcYHtViLEM4RP6/45Q83tVAVWltRunplsc+6/ET9gu5qt4
x60ern90FHxlHklxf9kBMhomy4OyIsb5pzoLMhUiLcL5hUXGG4aI3+/RL0YE
Sh1foVnv56FjNWsZzyVSfq0j82/+vDCziMO9qPQ3YFB5NqHIEC5vdwZOZwg8
aGfB57RfKLdF2+fb05KSl9QyFS56bf56cFZLcYZ9XW4108sWcImWXAcbWR4d
IPUweJnO/RJQXvNNwZIuP3XC6NgK0VtJ9MSwByAyAH0dpFrvP66nGVSoOnbd
l6GbJA9/WwSzeSa8s/3ZSE7V+HAqv1yM1eQbu+X1hKebAt7pisVmARSfGKEp
8eLyDEa/hLCGmxDjs5eIw9trxhTa9SKxNOx9o0KV49Bzi0GDH55J+DYPyu73
t6aMv3B+Ntq90GSeV15YwRClp964i3dVf5s4Bovyhj7eHUnFPqPxkDOFxgTS
A+ZBWP2OKKKcCGRf5yXRobYJEBIX1dsamggYcbwc3+J0bfFkoDwyj+1UjZWJ
WyM4oJc7myBOvcs0DpzwnwURAvvzBsH1jEJgnKorU2ToB6Q3s+I/fWc0lrp0
SMHTqGIGmUAfcMQv+W6Cmik/sL9rN6G+wNGMonqkXJGEwmxaP6b5fZXvPjP0
9D5LU02fedQJolMVoaoOhezE5qvk6XK06rx7alC/GWWhIUUqS0GMO8AhzBcj
rrwqCqmntgUiHH/ZYlu4ZojH+cu8l3a+fuDSBHhMCdmtJiXVEOFKH2H0ma8l
sA+7T8VWmhklVBux0noPvXYnjRC2cJ6tgUDF6R+zygnZjoGxga2z83ZFUVTf
XckslAGond+IXJUb+rbuSzygSKnzvDZRBIUsIr6w9u3fyQtxEPsZiBtg95fm
hp8M+WazZaEsK5XBoWI2JBKIxXkNXoo+QfZKnKgj2bEnH0HW1uPeiY3S24Zo
/jgbUHWwKqsLbvAZfNfpXjDQr212MTEfcoRCcJxe2jkL5JNGzroI2bEo/7j/
fBlfC+wi1XHiA0ydhKRfgvlHW9wA9uLEgmCbiEKkNPrSU/rEvBpt7fLSUr63
Q6y5p+0tHGTG6yz1ed3wJyBy442lrhTMVhq5qec5GV/cmV8c3lv8tvvtm/FI
/tqAWYcEiMxSrAinm1yH0veMYg5XtzyeWteQdD7nUwiHLpuJr2TyBNnz+GsH
T/DzPns0fPtNNK0rWUWWh7O5vwDYm+zKw8H64mBub6HacS4nMNi09vtZLear
+WZIr+jMcnujgjKPO4CwBFbUr+1eK919/4Q7SBlHRsCypqlyCiF/wDZQjooA
IrBL78h9csqMop+a1DJRYiT4lxa4QUIUS5sgdhW7onr8rNhdRZ8pB/7kfsAI
ovs7AYZ0/AZbrUfeDaSccwSXwtqpcpWh3IkPaBMDX9aUCWF6m8qCkJwBGmYP
HGUADr2p8fQMl8TjgkCxXjHRjXWAMGvMCa+ppMZyLugNGRrWEbzkJcEy6MwD
IROAsgsKshBsNZ/7t///TZIDYLeQgtakT/BXdpeJyMgaZd7Y3nqZZf0/aHJS
qr8Ua0+weMkm0p2eH6oiV2okVd81txx0ujM9LrTD/Da74gR/BVcRSiyVnqLz
p46sgcTGM+zfi2vsf3yBzXb/TsanwqgZiu7uhKmbLSE7vWqrvM/dlgfmf148
voVtHYQTWBUlYN1EkoIK8CJ3WTJumANqBVjtGyVLhrrHROsY9/6taSQgT3MN
Wxac7dH5v0slcJD65FJ8n0mvPYYr+NRbb45pTnmNmu39zIpTslvyNUWmtB3Y
VOKQwO/TkqLJTgoJPMCCHvpEnMLusXiWy7LpEsq6RqYN/Tf3XYFjprYK2Lmb
ds3xs6sbAZf2h3ec8gAVst7rziTAVSfekwUVZm4EIrDUMhzak8hLgPh+DDcJ
p8HWZDdiShSPnq+3nWTr03edAY12/GU723800dA6cG6THcrtC4SAunns09Ri
UGlr6szG/qgyduftcJkvqP0ohGKlAGnWt0PA+tfazeeOggMaJ1OUo13Ew+2d
iU8Psim8yQIW46HI28WTYcjm79bEXd3NaOSctmSjVRFM11+PN2aLwlHs0dfQ
k8FFoFzDknIDr56cIQB+reBr7M5HFwKMJ9DURhRBrl1bmfDGm8CtX6HXSIuE
L6b95AeiKYbyj5pSRQvJCVYJYa7VLhxCgLeKd0p0GoGr0RrCzPQ9Mt5mkDNA
vtqiO6htlkN9iGp1btXpyEfhLUltWqrr0DfhhNJn4fP7G1O59X2qDlg9dkxF
ec84Z/cPv3PDXLFPa2euzvVWXyM9uusYJWwg0BA/OnIQ3vuuHG8fCw8CMEcX
Wi12FNPul2iWF/kpiWUECEJvzaiGlAJM/HYOg3LRcwbACawox8O3Er6Z9Rov
gdcygBeH5zwfONWHxqU0BWQhkfgYJX5qDLf0hskB7vEvmep4BghWWUr24yID
iLCclPWW8oDLxZ2QssWT5h5aciRDDhjPi6voEQ4eN8G+P9WuRgf9HDKx7n5i
0yZIEnHpSWI6S9YCOzIWyv8NFxSQzyyuW1KH5X5ZRGJwsZHp45mElfsDJt3b
ip/xk0tRK2+Fg5Z0LJYm4axfYlXJG0we+tQlpDtAZctFku9JSzgkJ170WZsu
cZ5OrUqikgFKLboZi2V1tjka6WSbeEEwKA+x5J64l+3Fxpywx1uBMRaZfwwK
heQIaYeyQ2o1CrUIa28kDJCNXpBxLnZwI9oAXXTNAYlSRxAvGHLn6GgATKKn
qXyxFG9EukxuSmu1VTuGGV1TUcM48jtcKtCdtaNboMJT3IMG8UfFJDE28Z7F
5Y8H+N4ybsa51NL+pqbAD0/78ts5lyJw8YiAwiyCrxWknTC+FimySgtCk64W
YDnjk3tp3Y4sNVUIIubqZWIptiKrkbLK/eSMR3CiIFwF4Of9J/7q/FbWEsRV
7hZZcPzRofyWeawcHs64pmMkjUJhB09/v9AtFsIjB1H0h61oIGAL2zoCr8pS
mXhd8osPo3rf0cdvRgA0KEct6hRIoE92Tebx0cVW7vh4wGYye1H7U1Bytb17
fS4ZrgZiwY+hxTaDG1jNwEmh/dokEQeA5oXehzbOzRorrvL2ZikX7JuSHNT0
/c/8x8mKxrbY5OHyenUf3NlZnNVXqaDuyGraZuBtBoF7JDpTRt+Ru1rRV1nb
47D2AQ6NgYBzuXQzCfghJl32ab75JTTdE9s7HCFYQ2iYw0RvR1Q3tBvbiqX/
ocW5c5bZYRv3WPNePB/v+nrNXubmQvNO0Yg1+A3SwptZ8BtpnSbRCxi3h689
+04y20WukMHfl8kk+Hp+GYg4353KXorL/Ql/5M0JcD+ysUZAlTAsBAF8I6vB
0lZZub2PIJ6fjj1qu/n9x0t96xchSQJPhrVhWqQfB3gAGqw3wSvKxTcwxI6z
2Z70MmDb25SpLgsme94w+Y4GlaKPwfVjtqv61Ql5ftX2LgS0gaAetuxN866P
On71I27VEGBs5MM5LJ9747HC8/lgy+gXbTioMZcuJfnJUjVS5vE1OojadFn1
M9hOSn39rKvnbmGs5toZURp/LRTI7w6b/Y/SFJ+MPnLOtF5EL8I0aCC7H4ot
UkQxg/TDxnptO9V7fwK1WsOUzTEWhE73jk3OiknxyrNsXPlqELUWuHYXTbIm
7KOcPt3JSHHSVBV5aPWSFXKikRPrfWHof+L6xayUr53Ye99oSlTJ6+BI9Aag
eWOHhcWUbdnK7cCgttj0AOBucPup7JdDNhIG976A87GcHWB7HpYi6opOqCMx
jc5VlQvPh43oEUQI+KBXe2oSdkf58fs0dFiExz+zc7VUSmCrI1m51OWL4ELB
PiJsWybOtdjnuovbE5LPZDgRmPjga+MwnxQSzVSchq5vurB/1RwDsdVXdDUI
FsCr1fRiuMSWntMsQLIuwg7wSj8oilWrFxLisGj2CHCsXKbKcLt2o7bRbCAA
i96JNvPdLTxbbGoSoM9CW/a4/nhBtwKt5m/Y5CVmGD1A3LU30eD813kPE7bm
SYISE5PoWXVAzcEgQW/2+gXieTd9OwjW5hjmAn+nUmrz5mq566om3L1OgUye
jdsvWknI6PhN8SNvg63p/2JiY62mUMZY/tFiP2ntl4LMO9VR1fVCLbuQj7hI
2xBHzETKB+/ndU7Jp1hX4anvTKptA6O3fDXYArqQJxtI2pizS+lKnN6K7yuF
gJHGIPC+291T8DCounkMEop5JuV9YBjApU8gu9IaMS1htwUOa4KnguwZAL8d
7evyJh0rracdAu6lzoM7yttvstYxtWgsJbIJTmD5dzDOJpOBIwQsrPRrBT6r
vr+LYSy1ifubCbtOOJxi6ge9T1pv6IJjgE6pJyKATFLyOZ6pLPDPgWxuX/Vl
ZlFgF2jqwg+55gOb7rBIC/v4OO08RQUOEGiWJJqWgi3nBouOW6tkJFZuqazm
RGsoDDUIxriJSIniHyAgqJZkrc+NFuNVThc/Pb+VDwa58MDnaa7jObPTXaN7
1fOlVCmJrJDVz8zBxkK+JJBLkggfNtsuEurFJcs4xrEusGjLAGGhldtZ+eE7
YBzIDg22VkkhyvnGYUifLgWz8Szelm2MrmInSJZCybcHtFKDkvnwCNOb6LPl
hXOggEiQLrNx3znSMmGwaeaEjL48m5Aed77WCt1md30jbpaOCyDiCLMikOrL
Aei9nvi4wRESs777DzcK7LBh8ArMTuAXdvCOW5/4wOP5JBZLiS47SZF0l4+s
x/Jj+1cepiKOU0UDAQCASH4J5HRB2xM8of0AsK6H0/u/uKWhbNW1cvA6z3ds
7KEhsYB9JqGH9Q1kAY/9WBCE2gloSYMi+TbISY8BJ05cxGmyAc6vQ+ur5YYS
Y30Q5bwKYw8KbLZ1PGrKj08Og4wRQHa0pbUfApzvEQzVqZs4PQujnWI4HYtU
5VP4DK8mX29Rv3MpyNSlMjbAsZoB8OycUqKwHenJYjzlJ3xEKl1ZGVgPQdaQ
znRjLvmeHd5xEwCowNqKHwvoFNYexe8u5cw8UjnnhDN8+Rno8GJvysKayAyX
znGyxURHOwHSXoGonvE6peSpfsAD+INPzvi52toRhME9FY/FoQi9VtZXpu+9
Yr/Boe7oXNaa3NKIEmLCULcn8zpFqKbPVirw4fDx9GDeNnVUU3aYeofvh/VV
cNrMVleNRr8I12NlMugFlampvw8k5jput2Tpsg5V/2lYkur8ZVdx3kjxbmSD
gaL870ReGecodOkgVU5bgRpPK4u0r+fwWg+PPkID2XEGIT9hRwQDQGLQCsyB
A6kJEBQD3Tl72vC9qvKSZyzelqCVjV/NV+chmlX0KFuG6aP34jas9rLR986Y
EBmcHLLlf0K+PECBVXLeUE9GhECh6OvfA+yM0Znyfsfgms4abBUSKCz7Aa3I
ZI/LKd0o5fL3m41Kkdmb0zs5Rm3L6TzqrP8hIGFS93HVbvtxu3kcrm651KEU
ojgjLpsV/iwjxLMmxSlybjKDIXxguD9Qd1St2eGfLM+sOcpiVpWMHgNxIzFa
j5oH8t2sGfcg/Ad68Dml8aMnPKinnEmjzUHVD6lGEJhnZAkgGA6QItzgvRRs
7efJYAmRzl69D0KgZ1Kez5R3O3l6mRa4LLOctAfNg4uBA7Q8SxpaGYxnxtAJ
oRmjqvKSgy1cjcAUAI8f8Ye0a9PCdxUrKMP/bH51miaPeLJtYisNC6HhriJS
zw1eVAzKTSS7ZuzPc+5XQCneY58pglhcb1D8WvH9ymm+5SqK2vFXJOZz8qEM
feHQPl5DV31tVzGdsoVVH94Nl6c0O6uxl46K/xcPCsX/M/TTjFenaDF5/9ME
7uB6ZRrAvWaZTEUXmHzWw86nYQQK1d/qeHLV3kgCshOS14W4uRIBaOX0NFlf
A9x2SzUYGHHobkR9KP4u8eC9HGl2jM7iSA+JhYjLzdStg6h+DmMCFMNFqjS3
E8anm/oH3pIQMujkloRkvJhcNe/qypKMQEgwbqEtoKMQvqoJnIbmJPSsOrHQ
q65PAN1STrQZwb9cbJ7i9R5SSv/pLauO/O0PMV7y36n7pf3e8q/3goYkyH9l
wWiQYaHdabUyeRY93cs4r+MQTohneaGHJkP5jab0zLxDVXN89cyroBYW6bCu
zIwWRfeCw43+rjfeu8sP2oMeL80xUgtLkCT/uU4RLxmj3IRhcuKnUTcbJAWb
IMviyNWffjnpUaj//RugkxT8vDX8g+I8W8Tclt4qEiQFZ1c7eahG7psBpWSc
VqKSw6XztdMAtM1dar092DjPYFtJRkkby3jrUxRYa6zNWxu1myzMPy1SfUE9
WfxKBgBSKNj2na4wDMTEPe+leOA969J+iJc99SvDZvh9YOzG2CKWqIyqziaq
+dIzFSiowK0mGf6XWzlXpNWykD/hW++FSgm1Jj1d4AZ1whGSP0n3gwhvW2MD
0A9gjsvkA/afdqsie9DWcqfL3Re7PWmLYZFlxsANmEkWECp9ykQCEOGxduZH
Ad2aPpfSu9M8vJKTvjIYMmkaO6CmU7O72K7j/absMrp/xeJMhyjviVmcW/D9
a+53zwFO3IYp1M5tUPLSdXuOalWtkmXRtbBIr9YGxMcVDjpQDJ9EhpdBnhYo
Q0bhFl2pMhG+oTrgcphfSMyOYQwF6kQMiGLPkn+nxDOzHTDIdtLvSyECo9mj
WFrqBQd71zCCV+vI3KW1hNBhb3ZWDlNdO7aVr2RRFV3i1JLwjz6V3XDqvmn6
PjauvUMmzcyt94YqQMzcFJ5ERMJjfbTfTGiur9r/2TfkwYsrpSGalddOiMQP
zViVShLjAC/KNWCdQwcHHrrtS9SeTX5VW+g+IO0Nn50d8M6FBXAiopTRWVrP
pI+H28T5riWJfNTxPZjEsWCfpo12T/ok/nQPjgvZYpzJdTkN4lbaiB/dSZNU
rkgd+ewYpT5UO6apO9PJOcNdjewlO3X4VSswV2FkBjaRQrwMmLXH3CLeT9H0
4oAr0r+wKMsNGdZ7EBe718EskJeZTksbGVcYgX/xsYAZjFO9aDCWBSZ75VCW
Wn5nc5zZlQ5u78jBudY8voweCGebLfx33kS9vNXGN5fniSpkhCZqn4tdwfSo
TlfODj2DI77QNaTzetMU9PVu9PRctGXSSb5L1L4XC5XQ8H/5qJSk5C2fjYgS
5e+fETpqgRZZFwclgZlB5bNQqEySgg612LVodYceqUAUH9ZNEezsPU41YyP6
yyIQdMwVnJ8CCufOv7f7OyGcYhcPEbNjYH4WAZZM1UHqJjmsV3zGdSKGs0mI
ENCOmzyk4o6CPKbw4/MtjQ1hLYL0U4g44Mi1+7MreVV3Q0oD4by56MhwT2F3
Clc1eHgLKitmLbbJMhNGe3+c46H6YHb7yjWqkpndQ9MT/EBPaZtaghgRl0ao
URBRoqg7CEr+go0fO2qfApwRLQnmhjXrPUoqvsnX2aCTJ34RA1mXDm1RAx0G
wqy3dIEtyzGST1t0vB6F4J1TPhdYgUBBLYBISIn+GGQgh4m42E4IxuCAWVx8
SOC9uLuUbfwpwZoHo9uK8PdlFYSZvpuQVr1t/agai2fvv0ETLfpuwZesHOan
J+fm+3rV6ShH/5u+rONt+XvK4ShdtreBQUzNu/WjfH05qWF0ffcX+ThwKonj
ukAlIe+iPRIiHBjNHDPq2sl2JF+U4+rWqAVvTEvBstSAM0Qv+Trn4H14psJz
qeDuca2EClgB4tjgdWhXi/Okvpbm4GfgD5H0XSvsEXOGAS0UPH6VV6ELwDJk
8Wm1SuxkwXTvXMshIQ9Drk4hhvNQOMpw1AmUhHxiqirV7OZU51hh/GwvhDre
9kkTIbSh1uwpx44Ww33Sw//XxCBmIoCOx/+Eh841A0Jp7z1Dwh20+Z0Nhmkm
vWs1zJ5o4HHfbgb/9eibvFoE5LVXPH0uEHsN7npI0nFxSu+vf85xPX3P7BVZ
60tBWUcRtkU+/pOWDFDOJrO7Ixf9DnQ5U4qP4a+p3CJrfyBPjd5YIL0/TiKl
5n+UVsWC1c4PL+7n9ALhUtAJ0r8yGHHIgtGHEzVJRB7uPsEsr9ATri3alcb6
2g1llFf2JCFZgZVjoNHeSyMbo2H5pSg9G+IU7irJL1WS+8lULVJ+CLxHQdQu
R/0jDuiElZBqDUfkntL8vk1v0eqkpcVe8vpOTn1WpUAglfgt+02dXh0OX+It
9E+UrToikTonuGKibVrKJOaMblhPn6LiNZXayqotwLqIgeubWh1eH/PhiUnV
qPVzIwBR04dqAFsH4RKBwbqJ3YefFqFJygvYC/B2M4/EAoGjqCtSNm0NTpiB
soPWtGG7ycbL7Dts+q+zuvQsikD0mmItE/hfzUz/WtL3P1jjkIW1/FCURTm/
9wDqt1DffAzO21QuU/OPev9bWJx0cM3VjpxodgKWaOsKbOCHTDs+8ghBvys+
qSxK9D8VW3lwUiud63RQ5FVs70KizCDeAPzVJMTxYomFS++lmJaKOv6unD/h
oAK8pceQkLW107Jt6dTD5Znf83X5rjNZptDV1wFRDGECJnBE7JIuFxeyrIia
MECbYYMzFWlLKG4la3yWFtJl8op4Z071avhqFWPe0xDheO+OPsbHZ8Edkgqw
Xv15RV+mlg/Ki6xVjEyQSPECMZUoPh8dC3Ry+2X0U+FXNhd7z/w3hU9qi1mS
Gy6Xr/8EQreoq5o50gPN7csNOwkhw2mZl3YiSdSOlRud30M1kzPXn/XsaGR4
NGi8doMGTz+/PfJy1/JSmn59egUrrijbodOJ4NVfW9tRjLRjTMsfnGMXmvfZ
HNRKii4+W6IaEeJmd42jLierDfp052hj4r824Ngn6HiUkUachaLvBf/kCEVm
hzc6vZkBqLkiRwnsFtp+fG3Sw7UDA3dqZH6doJwy0Z7POm4gt9LELchMg7OW
ive4jGzkTCRQTZKyRQulEVj9sS9uewEN/FtUlQfXcgzd1AfmF+lyJwRMSTiK
D96wanD45dESyqJqlIZ9juaI8hnuc65v3mICR8GLFzincurYjbs0T+13s9/3
Ww7AvrUkTMtqK1g0a3H3t8gI6StLsk3ZJ5aVZYZB6F2WeSBGCK7VPXm50epT
MWtPi6o+Fiw7ovE1pdV4K8p66dWMEuBaznaWNPddopUyWSfVT8mlJN6JUEt1
FrZjBNGS+3Kf6cxVrf4BA5Z72Wj+w+DPieawjtfJC6LobcMZn/tomadmsn5j
ftkLHOxKAq3tPs0Or2q2AwZaAEiZv+7ECTUz1PIEEUy5kzoBZTwtE5k1c+gg
rGlD1O0h+wp9wn4iF99nhxqvlqvplSQ7Bfkqjey3Bj/NRgTz0LnYPyVtrehu
AfkMC/OFD8+giPeu7jmBK9uV8sVOve7xnqsvjjOTfayyVpe0pEZaZrGcaVMY
stRw7j0IhSA1c4nMpLBZsWN2tAMVTzlFyEJsZXxlySpU7C5YVd0zKP9I9ON7
zjttTTW7h/RqWRlkS9i/qth5HbMcQW20sW0TRsvK1v7IVM69cjgdPR28TYjM
0UaJlaYMxrzJ1XY6/Ro748TCpx8PR9YJqR182+aY827nuxJK3v8FAKx9EiHo
FXlaE2DJjvC3YZgt+os4WzAjzvcyadyZKIFELMSVTxLWFzy0hMI0s18CXr0g
8DhOMqScvverdPa+JGKrX9estvPg4uuuj18/4PRzCv5kl3/DnJAi7OK3Sr+6
66CDZ2YYlyEdUbnil+o1n9ngJdrWFKUq1EU0YxHXLgIPTvYNrKT+CbSdnXSy
KT0wk1ywkGrwCciWNP3zdnGFej/X2ZZTykMs0vpU8Z2RwzdXeU7LIuTTakSk
r7ArZm+rXagH3snkVQfbkKS7gecxA4zAZFIzt9PZtT4kdQOnycRxgyNgUIIo
sjMSdBkYsE1eQkVVxyEgAFWjumUg9eYV4H1ZQUqVxNqi6Uh1JkRffPeZVNpT
eJJGKmlLpMlXI+JrEqLGOrNDGM5OiMcXdXBt//HV6+5VCaE5UNxUVOyTO/HJ
tQT1hPv7U7o7QUR5GpE29RFGNly45sFfcmFu7P13EHSHnB1U96Ny6oAUPlc3
YXWYAdxrr50y0Bw2gqIKCGjYu6OFNvm7HHj4zscA7cIiKhowRTMgL95wBLc6
USXeUf3C/GZvQorEt2HzxjOxmUMpbBMaE8vofR8yVB+pVCyXZOyWhD1MI9JT
VL6HzBQ+zom8ObwZNo8hHWXGs90KK9IZBp9TDizUveOttxrzQnHqCxJxHrUe
U8dk735iWVhkBepW2Ji7y1/J3asJQkq8EBVxnUVWQY96j5S5BNyiBpLeSfou
mpCucUJe/1UVPu0BDHTQc+zr+gaBpp3fPZFPPFtntT9WF5HW/gMKIBI84OcI
fpjCAT+yDds/4XI+6TTY9t/tAs/WnAg6mYm+HhAeefCYwNJpYq9LajvJojgJ
W9lU4GE9oeDcOuGUXJdpmZ38xCQICoqRLpvcv2N+1MZzaCUV0zy0BVH5/V+X
DGDqvJanlE6m/LR1KwCEyHCu9zUzRoYv7iJm25NvUrsFA8fmU50VT0CYE5M0
cWojwlltGHH6s/gY3bDcMTrmeW7aamwPkwwWMQxD+/8xqEi2+Ha4sxy+s8z+
7rSoNKszTtKsU6lxmsiEJ35iAMEUUREk6CKuDUsEKK5ET6qB0FAxlBS9/lln
zeYnjV2Idganet6SYNGRHTZxn1cxaD9LahpnvimwuBGPveg0vUbe2wveUYjL
ckAUzy4EfvmGhwHY9vdjCgl6wzynOGjN/rVlzQ7MgM+rNeWm8iNYyJeEMCXb
2fHhmsBxBNN+CY15kFiU11nsXGVTIVKomz3+zMlMtyMYZY/efGomuMd1Boky
12ARs4siH4ktErAlNRaTO6jMp1LhwChcI/ekkFJ81GmyORgyKfZAIYmMKEOt
KM+PY7nERLvEYT7xF6mueyJaur1YooYfhwuXiHSjZE8NXM19syHkpFjY0pJb
8DLEkw+ldOJ2slUBjLZqguX4iO8s2PXTO9tseAuYfCefzIP51RUVI5r/7d9V
ZEKxMFXqdBoiono/hAL/SV0NHhMQfNLA3ChhZvqEnnG3k3EYeEOrT4bVJheS
9DW0V2H72sSyP9oRNnnsMug6TF8TQ89nQYcr5O+VU/rp8L1rIH9ZH+Yusw2t
Ijpni9FGxC4vhMFAhSJw63wQVxtF7oaMr5iIbIsslhZJdaUFdaUtGPdgqBQ0
eREHZQSfW7GtIhe4NSL3o/WSHV+Po952HwbLTS5+6eibMCNvr7D7MVNgvADh
lUd5B2sta5oMQ/63dBiGAzh7ZStoeIj+06bDWRLFsGLuOu/ICJNXiYY893PN
7+yD/oVNPbvLqqGptrAssY/ZWYntzoRJZCqUvKzJFwQz6lRqwOkSegy1PlYF
yiwNL3Bt2IRbeE6VAW+aHcr2qMElvKvJ9Znm9ayZi7vR3ufdtI3jqFRj71YU
kYr9VMt4AyPsyxklYxJ4haMjcGylPSEppfBzE3zvXh7XfY9k1xv+w6g0sXT4
WyMg7fvgiZ6JkAgfT9tHuGCa6eNftWArIutGT/aLm49z8LJ/vuzBip6c4/Ul
GDWMsB8SNh8YukzrCITGnCCiFIw4f9LrBS3FUtK0lotPsk/tjjgf9OHdpAfl
2u2PbN68og7/ham7to7zDcOOK8a56VVKmam0tXWgQJM9RpQ24GUjSu2agoNq
IsDLABGpvDOGAxb/sw2Irlh8VH3QeGw1GA3hpV+F5GwNcIdvD3f8vx86tIrN
I6UEaVoLwvR3JUYV+FXb3qlaf2pPIr7Sg4lMcIb8Yun3L/KncA+FSkpY4gol
8cBz8AZnmCjcZbZt/zaU/mX76nCrTnGOlo93rw8ASdCi597GOmnYHc8Otr2y
DsBvgOLLW25mpgZlHjLtWLSrWhvVI7ZlK2xO4XOOIPhjC/9HaKT+7OCv488K
iRnUqDn1+578thA4V7DksrJWR4KLcl1zVQVXEF/k1es+3kBxEItTxyRXxMB0
Ocnm/v1UAjKss2HWZYuOnS+0AiBIpAy+ewUwTjElv4IiXM9aGbd3aM3xITsa
E/0aO7RQxAkuvU1SPgueix+m0xFkTh/WiFQps7cHPLhpizys3hYe7LHe29m6
goDxbFMuS4CaPjV1d/9HcsrnGo5UutlJ5TxwNTi1nn/0YnLB5Js6kcM29C3H
j1O+ovvrpIrnuOYQlIPrn9Wa9VdIVdrxkG00y5YIfecA186+eyHtI+CI/XxH
HXini1qVDVg8nVUYqwPA4h/O5QuPNM5cE1vFaK0anoBT+UTTKfmZUQaUkf86
3Xbl7ODFYEAmwKtLKpMX85LLpBubMlKPSo93X2ELn1eLL9jnW85iQ5jPtIyV
0TFxhWXSMYGOV9D1uzMuswMdP/zPk68DBbg3jlMYg5vqnqMiBArl0ExX0QQM
Y+GQG3IxJf6zagct7c+t+5UDCAFFUqsZdRgZFXQ4hRWrW2eCjRJj3VNfs1BW
54DyzN7mnjc86jdGLbKj15y03zGZcgiG66/b7Iu9FiEk5bHVBEUGPiZYSXsW
60FIbannfdQ4+28rsHdXHfh7XdpC5ButBk/onQfGj2ntlvLwloo5LWSC9fuQ
q/i6LiwNcQ0zpmUdaJkU2t5z/qGgl22x6mkvAi1KCVcKUFUzTndCreaNGjYO
Cy5D2PKGLxOJSebNoHdOoKn3DMJdPJcGXr6UGAZ3LFO3PFTxD4vIje4sBbdM
rQsLba3EtulEAOO4emxDDzcZ7enRKEOdnK4zs2tTnWSVQ/yMmGLGAY+CwFzm
zk+Rr1+zer2zE73yeX0VJO5vFF7k9S5hOEG5dB6pZ6Yw4dSvZUCIiANTIoc8
QQkx+9cmTeoqW3mgsNFTIbmhbxDI6xf/yvtfhHryromUi8erazo+N4b+mT3i
12nSS+Hm8kZXDzibi9ZnWd6dgZXdKsWxyn+v+iZGxEQZ+45oCrilZAME0RFr
093SQnq1CGxOrC241vg9Z/FFcVhg3RHAUxpcf4YMGD00hdgZkCb416dG1QH1
JSUp0+08GoQl0CBR9bQuvZj4tGryNuoQPQGDJJx3Xm2xCA/oiZbddl3V2KiL
iuG3q9bi6ILhdN641vkPk1OWrTGm9hWqO27wgJok9IKmzbVxN5VCDRvHso9U
OWlDPjI/iI0qq/Om3XCrxyhgQ9VIKASwaRrpqeq1PzSAL1N4QUXaCRvuvx7h
CmrTnkYAHbuemylhcfJRfDVQRHFHcvI2jnohvZe9Fq5kRwgWIAScjeZYUFMN
907uyomAX196YYZ7YkDwHsuogVcHenifVT4JJsjVxskge0z6zba4xe/F2zTq
ppHVh2nlhLRUUuPaGKFi0qHu5f6s1uIfiXEwlAeQiUSOTwh2BaMMCseuyu29
zl7t0xhwaZs2VGQyLNQ+qbA4Ipd1ccJSb8q19aVlw4l1nXhyqNI3NnmHs2lG
jvEAnR++OPahvSwpUlcBoVQOsvR2PXqFigWZFw+zUVgUsao306kXSYqufjPH
z8LOyGbpH25I3kYADeybuhMumRR7kZdTusAbvFaXjMlyrhdrVmrs30wQ9B+9
Wj5XsFKpOYDPRyJokJiOrVcgO9EVae45y+2l7hv3m7ZZIXtleObOyDDf6IPE
eanDcjZgPFjOhp6x0CkyyVJBpWQa88ecTFG/5d00n+8xRflV31gkxRE1tRl5
ZrZhHOxo8upC+5pyQzCEJoayThURhS8gKz/dvYFfwQNFJQbUytMLuKtEAKaV
CF000tBZG7QuSFaeZRKMcrh/+M7gqJFCSceEuPnSkj9W0eCf9uEf0HFaG8Yt
LH9JxgGEE6zdpdmCBDWmtlWJCgz1OdBJM+aQpmGyHlBcVZxLziVeMllU01gZ
Qi/N2LSLf+ovfOYMQQ7xVlp1XkgWal2KN96jE4xI8KHThYjmq5xlOO5s8x6a
pKKttxfQIxQnHA2bP38dwWpgh0Kyla70MzstokB/GAwwU82+eKCt88uvHe7w
P2kZpYqGyMYrpKdXOzchThN0AysViHttU6EfQuIiuH2cNeYhjmOPA2AiuVH8
t129Ok6/aLrXbZbZkmS2M6gRieIj9TX7TLlfgyDMCPN9rnbWwZp4qhXg2GDc
TMRmehQuIwITLvUpB+AUASBIaHxDqNPfzfC1O59Ig2jVoKcZv8RP8QSUFJbo
AdHtwlPqNECUF2KlTSJdUDUFduQCdd9Oxc447h7jE7XBPuEkOF+KO8Vsn5zU
jaRa7nyWlUkBooIjzkGTzVy7Z2NII/PE6qH4J7KiMOoR+PV2nhu9dy6n2Epz
FHNK31/3zVW8g+tiDOUIvAz3eXIXnSeNvg9sdgDifAj6KLIcTMHevLvXjhT3
McCvCd0gttfruXYhxdEalyOxGajhN3+Gfe/OTnuMgtb3YYS7qhT0NiqZcSnX
Q5tShlWabHNoUCWm7154/umFcfYYsIiXFGRTFalcIcnWCyjsT4hsdcYDypTi
Q/KS0UdpPqdKRMAbZSlxdaX8waAchU/PVGrhn8a3wtsUBS817kYz0ptzqyXn
DPO7qdVGVUnm+j2Z2U8c9ZKTLUvCNBVrIVmIkQ6FjueIe66sjn7jkpu0PWRM
XuBzp0oFcsbQoAyy5i4S+BTNRJVoxeIvrFqccfhsNe/pt+iNMbqTpPNTOit1
Dkb5uixXomAKRefHZ9KnSOXqkYgq8JJr2XBaQHpmbiI+6TX8ln7pGgSpPcGe
Map7KFwZGPKDWsUQ8QUAnffzjpTO7jIJO88RcARnyzj7q0qvcizPkk2bvU7Z
N8OwdtdK1JoAyiwsBntw74fUHTqz8YiedguUqq0f8unOHnupEnplh7Gg5O0H
OukH2ZPmGZA9fDWSaBdMMB/uwllwQx3OSsJG/6h9k0Y7QAyfBrSplVZEWoXm
sgCinRC2f/IvRpdQQ0dChPEA/XKeKVyL9SVj+aTMi1w0ljSd9xIokg2hut6i
9ISFHoFTDzcPgylCdM7uCE5noAKABmtb0GcKYP/5kj538HkA0mXJiL/DS+k1
XeYFKEWrCStMW2sc4+bK9ABTeWC00XyP4yg/Gsxhr5F2lqFUbYy7nxwfr9Ar
+/+lyF70uUddlYHr1v2u4eU2SZZZemzkeOQy0j+U1IoBeoMDDqbwamoNk8fg
Rt2XcM3owV87zlp7sXd2xRXFvGV8LTHZiHAvAOwsG62AKw/sZFv5VtXMGvoW
xqcth7abGuwQf//fjd5WEv1oR4vcU4ClQqt4iXxHdaIcCEcOn8XVSP8ijg82
wsXJ60HdCmHZNVhFx3oRRYcufPU47lurnRgg8jv4IvtGM3bwwoW7jLboBz9v
nFSKQlNQP41AF4bXKlzvu/fO72Z/+zb4mQwwo+/XAKsx2gE4Vs5/TqV8GDqN
bASxJzh44+Jn6jkAOyz18nBmKX60eTa4/kZ9LGoQWExjTu4ys4mceOLsGFxr
1Xr5ioOYDvOBdPvgdRWMKX43MzzJLbsYiitgr3aHdKgKU3cqbH/VkLylAxiD
ArJ4jQ5AoR/nsNF0MSqV8aDMCTRgtLXAWmuapPf233PCFgApDt+ZlWh9+idZ
0KcmvriJ9wZqVi/Kk9hIhj9eNW4s9LX0gOZXDItbvpo1S5F2zAF+mBvornPM
MQDe80vb2Kdsl7j89W200BSEQsGWdd9wMWReJ+UyuvIHyT+6Vd3pTVlz3lZO
9VxFPCEuSbO0wvFqKQKBMPBsio6+D59jUeP06VC7yHiEdBha7p0o13YtNb2a
Fap0DTWxZy8TXKqtaLdFjRQHwZzr/0uC1CdBRqjLqWK6vpi5ZsPtGTCVlJdQ
BXUErEmW96Jl1Wh6lsV8j9xxwoOLxkr9kLaVViKq5/3xDfIRKDOC45FZtJfk
vZJTEO0tWMxf3HTjUQlX8kkt61QUsEs1pgBzX+nltEeUepPa2b5hbB4ToElK
tiSczkIbPUtxN8yJylaoN6zYbEfSaZCgwb+I1EZb4cJBXzNn8ugDFPi+vmpN
NhS/VmxXQS7xqtqgsmWh566eO7lYtJun2wRTt4RgmqhtQarYJ9JgbHL46IwV
VqurRgfkCKCaqtSof/DsMqDjHOlvq66q2rd1exRn+Vow8UTlShLI+UGMbzjE
MkGbCmXLuzDTpf6I2gEg6YfQqYm6GPTpzYD17pQxr8TbhTiOVy0hZJ2Hb/nQ
QJKgYLriNhCd+QD8NhX7D0Q5nwf1l5/6i0/Qg7TRy89wr1oj4vejE+juiUta
+2IYq23PywrMCZMZBs3xZmmZRFibWlLsNvA74/EOu7bfSUSeCvDpDQyoalt/
dF7dh0yfKC/FMHv95/uA5ONClv3YmwhzIlrl3wrUrNu+lDEsdWY5aNBgKu/o
+fMX5p8K8FhPI4aLxqv5irO25KH3bcZi+EVpOHcAFz7+ycAAcMVZcOwBartk
PH7ePnd32kegqK56aCVuwVdBKWZWQs4oEMVXtSehPl7RUQNQ/uVEKKUpcbJU
TG9H7hIFbdwnjRsODE2nLCiIi0M28wvcdtj4S10D+NKxeWI7pf5cgRcofu8a
/zTav2u+ovUHQy5jOCa5KDHi1LB3cSqMHuuwAAvnwy//RfrCL1or9lP+biJ6
xXeyOA0zkJrD1Uw24EZX7fJJNFEzlAg1iWeqURRMhavFytCz09upTM7FxaEf
Wx30QMvAQwbumzpXYGLRN7r3IgIROtiTNr5o1AWl0UstD73f1UznpE3y/U3K
D7XximPHYUBjLsSSdSAPjSz/Cjtgh6kJHv8ZszhDB9n93W+cC3mQZap09jRL
j1K1rSgjwQurcQVPVtYA9hAoInNjg1gCa+2SLsjU5lVWDm1AVw6JnC2k3e/k
M/giCK48nZ5OsotdrzaU7A55+mShVtwBh28DjD9Kc8RRQeaHr16B48snYVoH
wBHi7UgkpCgHK8Cgu/iJW1+38uzzIPGmGo7ewc/qN3SNwK2d4MDC9PvpXzif
G2hAEL9Q/NbZg40uoCdpnMhUn6T1qMRLa+lwNgQOu11uDdPaeu/4wPYVQnVR
s+I1dm8KWdA3L5F1wDOHSY4T3a8AjxsC3y8ghZdzfQQs2cXfVSQG5FFYkmYE
1NsiiY7EdveRhih6z1XZE7zsHRGuMT9QTLG4VJosTx0x4W6gHj2t7w9znI4Y
9ddMSolG45Ux/puhcwMlx9bUoqU1sAOrQBKoqLCmSYvTA6Iid/b1FBK8VW7u
WTdIO5B5hUWhnVgve7qES0Yp87gXfBipMg7zGA6arxRGYqM25y8RqEtAOZPL
9R46Ak/KwihJb1vouGWg+ybR2CHD0VzG9/SoP1S6yh/v8jXztlTCOLS/npRj
1g/uxmktUrvrdeKet9OHiT4IRtk5DnMl0OETUVtm/4ur09aMf80GeuCf1k2J
Hkd1tSZZyIJ5xJFUS7Z/WvYc6th8TWQq06o8HHg5Kiqj+f/xSdOs9KxGWY3z
M+YATOz+D9hm1RS5pVWzjb79Rpfpj8A6rNEb+f+nZYFRDD1S0P/cj1sFvJSg
l/kMCxBG0i1LVGCayAC0Hs+yJFNyIdZ1FOK3Rl6kJhJh4ORyynSfegj2LiZz
T9mfZvXpS7Q05q9qXM4fKnrk//+9Ntz7iVLp495+Sp+GvDQ02dFRhuv+D18L
sJ0mrW/7o+8AKAJ7FtuhsJpFlY+/ApMNPkFz3SuOrz6lyuW0LfdZ+HhT11bj
mgiP6wK7pBrlrlKUiZUPBvKOITXyLK85zBCu5j+k8eF1pWYw0yQSZ3PHKgV7
6Ol8mV77NfqeJoZHoQmfdsIXfic8PQ4YEc4pN/X/tqN9LrPzfq9gwunVarHj
Qj305qSWZ/m4f3GyMVGaGtuRBw7YEAEd1+k3h30janNcvIkGhVUUqim1llLo
nwc/CHOIU0Y/Lacy1o7P/sAF+DX1+vZBt0MWlkQMdLZzA755kUivuC/Awvay
LUXxOhyctptCVbA4ZiOv1zD+aNoVSu81cnjbzhzw0zvv1JmKTdIW83cJl3Yw
/M/oHG8iaCPyH1UvCNm3i9H5zXBsyGYXSITVEmYSIvMo6Hq1FxgHIJd4sFnb
PPaE4qN0zy5ExofE7rgGOX2ML3y8/eFBhAS17s0Re3jlU4QxH2EH7gARwuXs
fwJmRPaVwpdTEnHK4r1Mqgu6LeNbql3u+4/PplFXza6Pu/cV4uBthF/WlOjg
7lzCuyoqmOHaU31hhC9c8Zn84bn3wg7beAonZJE/hDI1cVKNojYTaiT/IdOB
vcf4Irs+B1/UBYNKLhcae9p2E/gxwb1nwHoba5CFtAxLjUM1F/vM+OshMC7U
JCHie+lq5Hjgo7u6gWpvoacOYC2w2D/4CoPcQfEkmRsuolsJmqTW+CVg1anY
Mq1tquSBzM5s5TwSJQ1JrwRH6okKwdZC4rGj2KZ3pNGxGoyVwBCVbrlSfsoV
gEUdnOTqsvrf1yV1mYIN1OC7IZZVpzOqtQxFUUwrc8NdXWpQXCkCad6d7+rm
HP8sdagYKPaApf2TLqPKjbPq/zj6WeMXYKbrYGwmiDY1SNga1jHMvRoPLRll
mJJ+iBSN74yUZVXk+QStjHeD/2Hwz4JTCappBtBg0v+AKrWTXUNaeOAbqHXl
1sXrVUbPzCksgTPsYhV5IvknVLWu1FVhYrLEvHlV5Kq2UiD94fJIMfW4Uozm
dFPSkbc6GUAdSO4OhdbD7Ap5aq7AxpjG+WSU+fFcVUz3ijdwCkHsrQYauQVc
HJeBrJlsMY+bXT8fpFFrh7mwEgVkpaVQoPc5DlZ31tNT8Bx7Gl3rhVG5dWU2
qlkmEXaN5BCgZFN07kU29mGCoUU9VKhrQ5ArepgdG2gExRkGPipDWDpww08d
qnO+gXTwbxdrPaQQzJ+MMOJk+Q5UZzdh1+1JJwM1qwBJFVL0egsPYeWOzAF4
J3DFnaEbt6tn7jR/Rm+GN8dPxidscC0tjLYIgQHgRqddU0vqx+HyTn8/UDip
ctWaj7GuxcPI5JcoEybQ2tdhYXJpcWq/LSImx6Nl7F6F3JQYO4eS9oh80di0
RPSwuLxTwBHUp/Ha1Qp4/OxzaLctt0ZTwJLwdQTTg+no6aqWQqDLsFhcfA1I
o2rkwxnzNtuHhC+1+InawKvcd6jNkUnVwb/i4D5UQE4D79hx1+TbAXRGlgyB
cdew2MXKslMpzetH/m1WX3EWlF3+ZoxnOwswn+JpHiUMWYagHVl9P2YJ6Yev
Lmze6IcJVXWmAc2lWsLRrQrxfoEjGJhXX9wRHLENVoKvL8gRIILAAgjqcS9D
jVCRXI4gqo/lVwbUC3q32dHhN35gugNzZ75qBkxXBjEWCaLzo9VYrP8XnXxH
zxjUD1qGWZo6c3GhNeRdADOt2YNxiudlGuKFON5Rzi4q/QvwFPFoBvPxi+/g
AoPqU05B6siUvqM/87vAUlPumNvzdFsYGsh4xp38XDMm3AM/3/SLArdJZ3Ev
5rvReIa7f8Ht7SMayRAi3jmS28EhU6tN2NVP32Dzv/ZQBYCN3MIZ11eoipn3
Ltquu1VRcGyJfI7bCFL1/Jb4o3gcC9ykUrXFTyY2Y/MoIJoLUOI/IsXEpbb0
gNUQFmIkDNvYzbX4ZQ5rNxkcHmH3HCEuLiPMqVotlM1QuIdPrQiRRn1Ejcrn
plOnkiGW+oBsEohmY3MehgpiK1knCsHaeUZFwuJP2wJG718dQPmJvseyDKN2
guSKc8QZpgdBiEjs8DcUE91jqDSoz/1vQY1tkIurPo8zJ7cgG/1zKFXnZVXG
rurqlpt5pLBucsKM9k0cUyMxRgS3YY4hh1peBwcOPG+v4v2CQbSZADpcSLjb
YXmv9yDDwKNZ8AwDExcOcDXvctHGzC/iqoVjj/jP6eKSWZNelalFnZ85VY/b
4jq2BCTWxpiNuTlADCbLC4+6J92BSMz9pbNdKeglIgtfqmZWrwxR5Eh9ufWp
7vxVCZHmFgIUk25b6LnjI3waT/4/zNkdiNvh/dsSscZEMLz25NtW/nkmR3fv
CnyS8cqjNdA/G90WXOskbF9QaTuQMxgUEOICUiEcdk74r9mybSovPr2TxpJJ
mWOYkgvm4ng7xCQo19IMmu91a2qmvPjE2icc+uctAfV4fBO7HuBKPSt592KS
86PqsL/AMZfOx7GcnwGjXaDTxGFf1mUfoHx8v2FDHbJkgAkfUcNzfhR9I/Sb
z6td3ywYPGh8yFNJtg+6rTrcGjyAwAGGNKN/z/HuiixVMRI10SgHZCWK0RM1
E2HvQkdwogRGBbRN53i5QnLY9yEh7FKP5wnwh60IBVA3nLfQBK5Frn9UKUUp
VLUCuPnwz3/5f/I/rXtfBSiLQdeIx0CwzgWQVLrnMExu0/0mwKhIzO0Paxr5
t3Y3lypfZdrWrNn+A2jOrkrpjm27J6HFAMEZcGMfoImH1JON/N6QCQF74/n3
NImNISlgVvnmK9BNjWB6TXWBEDIYcMYKfXJme4iDkntidb4W6l2uodgRw6D1
K7MkT7Wg2jY2eYjg18Z9Ls3ipjIfuXBoqxOEvlwCZL8vccOFT/LLEziFzTsk
3tumBogi32jf6nZvl83+5UQVNwRGRO1zDtQID8rlVI54GLHrF+9kQsRL4qQQ
iyE9on8oemiLVQsZFCMGc/dfQZoEPETJ9p0ZUG+WKLYezkiBsTGDYBW+Reob
S7TvqIQwTyJvxFXT67Lu5p12/EH8AD2Ah78e2TfF9Gdn6cm80MXn8O8ZVHs6
bsXRvStPs4JK3cxAf0tYJNpT9OUv2oR7bpA9/JtSLDwyLqOOJO81M8NePlb2
3BYNAyjCP5JnYDwvdZStSGjBdvUI8iasQzeeDWMigmlJNEDKPerAp3u3TfOU
kcEox4sp/wPrKyrRUQDMkf601MWRA4hscuI131/5NoVE0sfZUtr4U0amYt+8
ddnXhJAkFlLEoEmo3nS7RqxpUuG+EbYn0jhLBbirGWLsdfi/YF7LKGBW0vai
ZRW3tf6ci8SjX6kXPGL0hHpEhtPn2LWmCREyqyNRbB0yZHRYmmWegOtg2c/N
9Rosfj/Qcn5sexx/sAfZod+FPusRxqYG2EnHJvhDTn7CFJtTPp2N2eV2pyDW
5bpDku9bcRdiFqgFXYsHMF9ndyQtC/UzcSTUvjIdbg3lhtdZvr7UkyOpA8gi
MWg65gC5BRK2x5lFpIPGQjXFJomSl6px3OLJQ/vRnKK/tr96uXGD4s/yONAh
Q/vhSFdHixVxYVszMwaLs28VoUK3xIbdV5u4DeuQ7d6lwDo9agPZlSh3KSph
/h7WWUnNgZqCoD+p4QvP+2d8uamzU9AODSscPfPI1/27Z++b8wOc30Yxxa0u
O/8ZF0b1pFWKHyZUM4xiNiIuBICF3Ni/xLGr5DGZumXUqr6WWm1IIU3n9+Jo
KsdUvrsXxjO6pAIFeEvEBMx7d4KqF/dHZeiASKTa7kO1DXqYgw4Q4GCnsnWk
jRDF+yVbNi+ZeuT+8iX16fyg/69jxpkj8+/TPyA6Ux/h6cq6h9P8M1x3svyV
MTb2iG9YudGQtChH3HFWzItVPdBqQf3rpXElJNpyPrXV8KwwxNPj54QS9zi+
/lKNtJsrw4rUFuUcY5iLYbq9CsQxeV47Yo/zeoccHUHicTreYqXOutSHZuJ+
8lvtvPF2ZTrf7xaMyEdJLGzW6qTgkNBkujva+ERrcrCoAI2jmY2z9Jvh+oTq
DSQdJ1H9m0OoBcFDwJAwxZxzrqV/f4syGotsFYZAWUSF1E5DCuCSIGYpXTe2
3K8aLhkDPCpQyhpyob+wQj4JykRkPmIk/FW88hKGvdhXG3UW5QuVpseCJOuS
IfukdzXycmg3Lddua39aIDPGTswr7KAX/Gxe0cCQrHdu55E7U6TLgcS+ySWv
fY7HMpnMO3AwYG95cXdijLal6u4A1K/4OfcyU+p6UTUdoyxdPvANZH97D1Il
+8eTPyVG/gAOJxZ4KoFM+1gHbxZ+Qu4IVIm671/ZVdhIwKMFb6R2HJwI8LJv
SDWeBElZNaiwmi92VcH98hqzB49m1pFj0XUPxLCqvr4VagrjuX2Ki7EnDjzW
vI3Dtu24rANkupijggbCjA/SVVog0dZt4jyKqrmK8t3QyVZUCTArgO4ZfWSO
Q5MjzgI769FerZz6mbLzMxifaIy0ou9p2bS1eGkrokQApd2YftXdmZkwmJ+p
VlOS+sz7PeGukEMIqupm/Q6x+TGfgmhKUR6aR1gpaFLtoc8n/fWgN2OPorfU
TNbkVNmNIdjDEC6Cdmc7xbrbUeRXgUTO9yNjFOyOKn1tWyVtTHGcSXUCPVn1
2Fqgsm+anjmUFHWmZSkBN2cXDjGjBJR0Pr6+8+eMo+Ui7JkyMMztJPzLY5r8
i70HzX1fncshRtGzcQaJpo3TlqYkkxktSBRNMavO0kKgq+DZeSVxYvsXBytT
BdqJBolR0tfw54UDiHXH+hMt4X+iF88b7xJqk/NR96g1bften7ulMM/uppSh
1DbnV6wd6+vaOP19vZOg8yHLerALuy1wS5oJR+zLHuFpj6aI6Ica11hwfl+Q
xVzNPf6msm8RiI2Il6vPBI4vt3lPZOnjeQFtA1ZuOXBtlnoJXHDq7yabtvOW
UKL3hI4G9d/gr8aYxBqyHs/akHeGCaVxrN0ZKe5SnCAQ30oaYZ3kA2gOceLY
e6b9LQ3to19a1h5Niha23SGefT5V8xeDJtftA5VPIaFujK9R8kLYo6lsW3yO
7K8JYbGChLts9qSKgYLAa75hGBKaohNizyFpzr2aACwMmUPBhTCojkUeI14R
eNnZSaM6Ofm6iFuqFNmQHXXig2CkIcgYc5kGOxOhWwD6FPWesC4so80OniWx
AN9u3DOwwLEKS5it7JOLcjQuevQnWKDo9BAzst7aIC8hv7aSCw9QmM3DVo4Z
YF+Eaf824SgDZPAMQLOqOWqZgsdcY9EL/ShT3AOUjetRPzQEk2GOX70uRkmr
wr7CTGYZ2Or1OjweT45gndIPAc9MSQL4/C5YoNBogkz3DqGpAtK6+5KQqExJ
Q+IP0UWjc1nmblrAJhGwdcTK1VVDtLoOVyZaLi8kJx5z35YEjHBtAuaosqVR
MzezoYvpS9ONM13hXrJIqMwBlpeYugcn3ROr2rFIVz2NpGZ7OvC+WQgTvFmx
PvysYk+1Lqu+5AxMiwaBN9FwsLPFQeJMb/lNIe6z4XvhrtsQoXtnx6o7C7lZ
iX48TJKwCZLVHnUAgJziJs4sghwy1kvwYL8Q+TUu9NGmYbQ2G0LUOa+i07ne
ltDum/ab7M6hqpWxDGY6qvYFq+mGACGQzxU2fsDszbTVa9yBqKs6wcO+9lcF
wwYyflT+jIkyP4+05hrtfJDXGzgmkSbBavSKb7w1FcM2RzVchtivKWzWzvpT
i0AC+4m+me268XNQ9uPYooHByfXIXqX8ESi+brxaxEqvE13zimp/amSKI2c7
EEb/aMWaEundK1IaSK5CjGndANLSOzEEGcsO8hHSIspo3TZnhcnGlvMbR/LI
j0HVw9MD/6lFfHBSE40TuPAxq/DtdSaGSQN4Q6vWNZPCuHiBQaQIt+E1wJEt
jYCuoq+HZahM8CzUKllaX5nx6W/Bi6mZ0j+AoYY3qMiIIfs+crw2a3Hy2NMj
o23oGXAYbBPqaStIed9s37ARunl93sjJ+eICAQ/hu6wC93bG6ANY5IGOH6Dr
0StR43ew2TXD/T1eylY1za81GuFiUBqIi43NThpfOCIwNqt/F4MBsYgWBfsT
qFOIo2X6vYHY61YKzWS3iUWqLH0ZNbAvc3+QRSL88Bo1FjFPscmdrkbf25OJ
M9/LDne58qzK7fi4HS5Hcd1aN3nvpbqn6pUw2eqqp8F3a7YuUqbmfemd61Is
jHVzLGOhLLBalRp1xcUnn57+TBSxLcjW8WGDUcvEZVDRhfuFJQeo7tKvQnvE
4mxc3OktQWEA95RDt5lhD4I6GpgKk4sNkw9Lcjm9+QyKrnQF+i5RprCbjTro
apCCi2/34wWV8il7EygTbW+gAfJfEJ4SVQKcPPWJAKqtcI1+F9VOUArY4OnT
Cx8X3MKD6AzX2FSXYiNQflBd7CbkIPW26wXVgdQ149yVwX7TNoLye5TsZP1P
v4liguFLPM6/2zkqdA057Lf4PanSyRr2cEvL2+OQ039dIaHmJxRB6HUhkbdx
AOIqjCcu9aY0V4CzTfY/Y71Z5EUinzrBkgfxCMlA+OohdQHQ4ei0CxT1RT8I
O0QfjGGAfVQv5X9LFNbLVvk6RbkjXbeQhOQEDDQeh1/tFqyzSog94PFJxh7h
gZqIsddOzc+oWe8Diz1j7JOso3a6tu2yx2woQU+SOKFByhtUwTshVvEG3UCp
6tOl0dY9Dt+ap8rl3AUfiMpg5IYivTzFdVwvDs1lr5cO5Sg9vWIbsVhbLyM6
rfwZF+l9j/ptpfSqzXjYbeFFBBkPhWxQe3dIzfnxob/KEg0YFweTCbXh8tPu
4xwGXnrvy6hwyslIgJoSMrMIaBorqf2+ur+CmlbvlIQOBgBimrEl/0ZKhEO9
F2266MOGLtwafc3WeUvD+0tsbml4TFI7VG66HLhtMnuu4F9xcskW0T6CDCKy
SVbBi4+5HydVGcKG/2K7u08q0ZnjB07baK31mKo/RXRI11RZBsPCQlE8Ug1M
ydEdPEYYhrr2SQsp0mxhNE6zV8kA8YpBBQkSc1ciAaWpSc/4uRq0tQBk9xmD
IQ3tllt53KHQpuIdg9zwusHY6aohIIe5mjoc41RbJRMtfD7bwgpcYfmvAv3g
EYvgXKqzdt3WUZbOBXBhTyIS7KbHGrIoBLFzHM35M33mbFV4Ig2YBqlvcYNc
rf6laZcCh/c8+NGqNFMwDCmd4rlVaH52fHOsttpKa8qluP0XCIhCec0EK8fp
K7HIJg9Pgzxj6rzDJhC2WstRnPaDkAU9mcjLldAu7IArwzGpOzKfNcrCnDa+
Vfzakm9cX+5E0OE7ZT8mp4ByJYgRPePx93awqC85KXWPYbYYHwqp11ZwO3MG
Sark67kpWcUMJinynQxWfcUBSoW/tYTbz1zFVZXigSY6Vl+pK7USqdVAdWkK
pyZtTDcyEozmxWKyo8CHsYQdb0HjLBxOuqepoWabX+bIx739VE2iX60ZKkpT
0QJGbHcmnA0w00jXP/rBfdCdx+P5oUGxk5g3/oTaYc/742UH0g7RkJS5Zg0j
+FD54el555+eGrQCDxuUieICWmU1lvF/gT7+GTkLElAekOF5aZMC/kp/xsfP
TGK7Q+6C7mdGZ0vIKQoIiQ2LaCKEoRw9b6exE0FNHrhLlAabaJhSkSHFrL2H
Yjb8q4JOwTwbKM+kdL8XiMZfGOECIM+mzOpCCsPE6BRrzbco3QrX7ZtimjG9
R7420ZKnkbF21k3lH46P0IyFJzIwighvq5TaI+/WxVyQBy+m2rn9xeo/dCop
CE7B62xKneUQfOXQ1KBjB3LbLXttFtobHDg5G3ttcISSxZEx01opKj3NbhtZ
gNrin8Ys8uWW9qKkwcbeinufKRCRDtq/rpOgnEnTiZAbQ8LYSG/WoKRUlb5V
S4xXkjX1rGlirFSWvCzWI7WI2MGO1l9MnTKdtHuicdkQcUJKX9nh/hEHWjPF
slH+TKdFK0IHV1PoNS2jOVB95eSnzMznrJsMiThH6SfWKPmUN0b0/Y5lH2i/
ItAhet+7DkUYWUAzSnq3AOb7T5Ksjo+kSxVbts63QxSq9uu/ukXuKwatYrZx
P7YnTdf/O7Cce+zviKug105Xhw8mbHqWQGFIm03tc/X9C6bIKiZ3qyl7wx9w
jan6WuO8Pl33jAR59uYl7bh3uS0iKUIGwAwQviXaVzz1enQ2LG92snwFAgyv
vYFd0NS3dv6GqaVO6BamVTKqk+OYIOSV7DgX+5uxl5dMDjJT4DznaFoOLeNP
IRGjyqvjohZkN1gtxn3zbNrANf0EtSkDpiDV/dgMf0zgD8tRyFz7jYDCK791
lCJ73vffhOJ21IlUnyB60oqPKVxOcsa58KQpboIZk6Ps0jTQnFpPHRQ8+CtT
fO6IRzazS+W1LBG7tRdgbMULfl/sGt0qN+CIJi4bM/JW8+uqSHEQKpvtw7mI
SbB3cPfi2qEKClOa5a3R9NsPC44y4cjdU6YUI/7wqajzG4C1WXjkRoac1YVd
J/74S/7+KCqhv5rGxFYK6krM22dc5Pf5/zqaYxysJUtoXVThcPxIxq3TtHy3
JxNb0s8ZjQoQYhLNnRcxn0TNbJ/u1ygKY/w4MZsTQbqoe8AjZxuXWFdq99Ce
TvIMEwnYvmcbmv4OvOMXDZ7Y6RwRG03nSG4W+7S2MYBCr9MyQLL4QjRimVvC
PouaavH4f/o/5JGlFO+nq43FDIQ/lu4o5xDxglmaStTEXaq+ATJ1F+EZ2YEe
Srm7tXbgNjJ0YjrJJNgskY4kLnBGqOizekbc5hdZBaBRhXkt+l2jqOdKF7bn
w5C3DnjgScfgazfHn1Gj9P/EQyfdMNVxZ16hADIW6mJ+HiZQJIEYmDYmR56L
up2A51jO0AITJs6DTeqPEReyGA9jXvTSF0Fn6VGl1m03USgOa9p1DqTaDXvO
Ed9ZcWZyKAxjAqQFm7VNnxVP6HzXPVYuww9DAtglrlVzSZ1jml+cmHjpxPVE
qZ+fbZBkufBhCUg4wtMyzmZJ18NoZmFnjRXCJKAS9zpXXFEV5E2GOxWDUwwH
yCmnH9fkUDQufKkMqpZ1AxUW0TNbW4glXSWPQJuhr1X2+5lwaZapyxAvN6xE
Mdsw64ffbv7wTBl5v3TSn6bIzNY2c872f8e1KanidkbolhgFfrsdfIWM4hNs
+drlgKEQK5UGvihuxN10Y2cIW1vy6ZVieYRUs/uv8FA7UX8qPa2F/aIf1v9r
jGOh0A1w/tfyfkm2EWxeS3bL5X1w7ZCNmeoTIf1mTx9nJ84ctUwCFkIK5sCL
6jcBW7aMbz/itmtTtkTmdeGmcojV4GZlBbXjJ/WYQDzcG3IW1JXzzCNreJ5t
RVjxWwcje4td/qbqCPgIEWFIZd6dzUn/Vgir8XSyVLvJjEIxxVniGhCkJucv
13hS7yufCyGOMlm5etAY8MKBgUs2jvlx8mFPuUoAtRgnAxPEF5+MkZirLNE2
vDiWhJmAHXV9L81+XkduRq3A+3uqeVxXosBqIKwChWARtVpnFqTNN9+njcqk
eej9k+NgCqWwhuSVr9q7eDJdpmmNL401/4Myqyfx2HIMH7HDX4h8F/uB+4Wj
DSXyWfeENlwPKl4VWQt//mK0vn1u7KIcbu6kcgFtYGgKnlWSdoqiRcCGyndF
gOw/nu43/QsWt3YeEKXeCbQtOraKY8HVMbDo3AAciHm5BALXMOn7p+Z8rKXk
DNkHMv9MrNrXbXE0I3Lw5rl/9k70qSv2KiC75XDvgjQ4LYcchKj35g9DeMkr
u3/zL42xzVIqZu/jpEMsGwzqFukW0SUvDkSYOXfq5tXwTZqK8817gfQj2rd3
ucnlYKBXYSC8f64mcwLiFQ+b2OH5eShsaYSYBhKL7003N9ce06lwMIY9NafE
o0Y2FgWf40DMIb/fxLtcGS7ZXKPfeCJPHa4OOJqnj3nWLbzmFyU1AK4xYGvY
39tZkLN8mvOnsz7aLj15pldlrjSZ9fkd8AEUtpeiJIzyWyP7S3Cpe09zbM/D
DWGbz1YyEX0k//TqDD7TRT5w1ziTfcvvnQkGDDk/tdVyTYkf1BV0NWAPRUyN
iSLPYdpt/4C1w01ICLYCFntdHj4LD0VTWvyZ39ODVZ+MsI0Ivi66gLyu3KKK
wbzseHSoK+B3fkCmtwG5PBGWtdDrOF4D5wCZ+Yxq7nu7X0dmH18lmDPxUBsO
M0kF24B4EC3L8plBDQHaEhFLdBv+uupos9P+4SHHXeSnEBophyCao+bQAST3
+NhXWd3ddQtT/ldhqz9RDLUU/VCk0s3kHXV+7dvcGYbjDjuKTIE1CaVfUi/k
FbXemOk/UU6V4bv5mvC9fX9pkp2ZGfKnoq0RhRuyq0ew2v/HobvmWQPWv/33
Pns5puIaYgf9VSh6RfcZMDOfN1F42PHXiYvpEmNZzrD41X7XBcyQv0Bw8cI7
9Pyc8yoYRzAtftrBTBzPfBrPbmh9hSDeUcfFkttO8TilUVZIsmYxVyrAIu6A
/x+SMKkI7OroHGhtLP5XlY124ZmsphZh6YIxMkYtTkPOJOe/xvtOH0oQ8EYY
kWTZsSxFCF2tUgU/WewnVJVYlzMcwezUY2pw59DpDjK1wMnIhbjYyCjLTVac
JAaaXL9D3YwTZDRborIvtadJokX4sPkrJ8nOPQIJmwRQoYOMk0SYmefleaqu
hqT8TvJVQRdkWHleqHWDbzi4H4GoiGDwdjUCvSBDlmue14jQhJ3qxElKyKMm
umDSrMA6N72xcvecXSdQQKIx5LNJqqZe2ITSyAdLaBAae7bD29Io0U3cgP3y
s3B2wY0/jBtrnd3RrGFZG+fvDFbO2v4oRd5GJj9wEWzffBB/Pk2paKYfRCYV
bB9V1rmya4HrQEYVx+QJttDsA3wO4cf1F8CXre7lQpiGUb0myV9sLu0u0vUQ
BJXO9mhUXs1+WhS/+mvSocG0tZLvd1iPSc7yyISM2yyWQHHJCvywVqhpyu4Y
3vhDNd2ga7PS/ZIqTBEX4FB6Ix8A1C8Wjl0jzCUd9sbDDu+9Dvu/smiAa5B3
mehyMiV86aiYsMWzPTk/pH8RKH45ts6ycTeXmg96eI2jFx1lllBDWVZXy1k5
30MZzsDJDrHPqYYcD9p9Hu/9deTvqcCyOfXExnfUEIRy0bIHXtrvChRtx0G/
A/hIjMUuSs/EY7ZeB8akOciHFKR0UeBwQcFRAyNr2ux2VKkJ48fc7PgDtz4C
l+CJFtCE2dxI6A1WoY8Z0hM0v1Pg4yNCu5eYPYfIzG8qovK9GfHzzPuvv1/m
5otPtmMDex5pxFfdvprciIC2eMfdWjb3od53VNK8LdmPqfrCOCbM2tvDzpIF
0k9B3EJxs22JasGrX3PgmdEVoovEYc+FQzDeQgluCIFp7RNz012Vff4MKE1F
wZVzOB42QYlM6jblzHQGiqXYVML6YEb5mfmXcDxwQKkHbCPn8nZMLT7mb9AZ
YHkbZWwZQ3rntKgBtQ/ldc18wQMMfcAizyToJ8S3kBWrRjj2J91Yz05DB7Pt
kFVCZhB5u9Dgz7ceuTAwJPDImDpA7Hx4/Sv/nADOUIam79yZE6A+eWwxV4qz
/A2CfYk1whxCfXfSAfC7FyGvAHi64OYtnc3Sv1C3+Lbuc9hhZk9fwrDwyiem
PQZu68kRLVSqtr9D56ZDESaq01srrIVGwhSGBWCLp/CVS4NWhnAHqXIle6Hv
F0CssvEtHKkmEWYDw06K0N6u0agq+SNFAEtnzNUR/dIE2NXV7iciOOGomesc
XGqgPtIYHz/6F2oU0lVnD56aVu8+4bOmT09a3LnHXtdAp0yquhuKhExaOFbJ
I8F/fQXvlSO3MOKqAQ2prEEcuqgv88ifYwlvWGUgCu/1uVzK8/sS3/bxOd9E
1qlYlsxpRPejk15kVtRgncpxNUZxI9og/F9Xp+I0ICu70LO3iZ73Zq3ULxmM
OBsdc+YXc8suPyK8Ary94ODXqgAOAROxGhAGwGiQMqYos54UPWYgQFoRGWAT
4R9zsxCvTN5Elsyu4hlK3lL3VuVh07ueyE6sp3A50Snx+UaHWxmeO+fzLRFh
vljNpqNDXaYR6g0+OaZ2Ku/x6eQ+3KbqtmTrzRfq8kXhMEemxu5CjL2YU8WR
o0kLbVDQ5+GtnnECw4bNSmYdCExMBeWSLPrx+PmKUo5wUM6YZ9mlAxEfxNr1
hff5YVVguYvQcs63qA+jb1ujHMBMR15cOhu1yKv93G3wdYtpiyr9cGMPZev2
3l2tWVn8Y2Zru25alZzGZH/aV0GqT8/mGw2Wrf1waclH13kupS+PMBPY4iwF
slxydQL4dN2Mj4IexgdCVkASMnJd6+JIs0Ad7hqbOwMYB10dPGN6zTEgqeRY
yzJw+WsrRc419MS+y+RpeicXQ+lDTe7IcmqBmgquv8KGkltwjB5vSCAFHA53
OUrYiTE9HwVoQcdeUiGnmAPh/vPyRAzBd/r7UawJVJ91TYOyuSdUy3gtl2iV
8VGjwZpMjF1sWoeo6EUy42eeOyUwzTcIVcx8Jw1afRACn7BENTiIGi+BLYPF
LBaFc3XSyEpk/Qrc2jmK9tAcQwWX0d6Xwxhn2C4UcNSPrcFa4OTE9+GA/vgk
2wMxtg2EVTt1m3OCLWC3awOu/TtM0T+1D62RwpQiBMH4x7Zv+f7r+Y0PHJ0F
4ojvQlbnI18GP/ZVfsv3VZ1uysRi5bTevokjqznompwuPAqb4xRoZnUc8aQ0
PDHUvkdY9OgrMUpYWlJuVSvGTPtimiIBD3n/f2EneyKfQyguyErtT9F719NX
oc5da1iiuwfT/+zZrjFubWcqci0ArmRQ6+R4uH3kXitQOl/VMwpSa+WHaGCt
qeg+TYsfnKWToQCPu9qc3DMEphJ5yUDYHcWGLfiqm5InUFrIW0i2XNB9L0SU
2oo2R1SHu2dgzDaRNPRyzQJQACUblJEagmEbQM/UF1qhJpKN894yi47fgasm
USD/Hhfk0QTfqR2l39rX6nbrCy7I7lDEl7pCB35Jo0nIl+nsed7QDhtrFDdq
G5LxosfJSSUQlauhpv0SnDa4y016hDWUXby+t1IkmGxPqeqU7VtqJ0mEHZv8
Gc/N2F/WggeXTfDThXDdWwk4EBhDuvIoKoGQ6S6HR5iUIDOQWhpSOEqmvM90
c4uLT+2ZYuxREscs0+5UAQH0Obu9YXoX0WvhS2XriRqF+RXyLb/dn3suNi5T
SmtIJapga1cUOgfKVQQJZ3qaVsES8V2fzYLyzfAk4L9ZGZbY3tvk/aeKlCd5
OcpIQnyju/8XMJNEY0k0SEjSiqB7e6/YGiUCZXnzo8wUD5Ktp4UCj/5+o3vh
QnYs9iQsfS9pZrlZZOCmjf2jEAeUfERu/LGQqJm9Gj9Pehf8lripDi72oKEu
KUjE1/pUt4KIW7RuG0CPZHc5naVnKUzayFFr0WT9cE5nDxHPouwADQDx9DXa
xEhw3+AoJNAHnSb+gJV+VQSvT+wdn1fW2VAzBRYUu6RJ9gOCSlXBrrr1itDb
2WpNbJ7XMq38y6M5Q1tmHaRyoohqlAVv9RW7NeTgzF1n6/vOPHWeZOMhcJN/
j/4DzY4wAsJxihszy+zMYf5uYDMygPbt39AM0LaEAiJB/rAanaSKszwZCpuF
jBqO8/cCIAM+WIl24ELcRWWpQ9kNgkhvIMPO8DgtIg38MxZ+VmSart8pfZUG
aKJK8aOYUG3Dwl5SKlWsGQNJBh+HnWZUEbJ0sTvuPM+pBN84jqkuIYcvRWA6
Ye5FL9usz4Y6bFKWdkjMrz3McsTJmWClgYiUw6BttRU0bUrfZfGZ8ITP/jBe
cVyMpy4yH55az+5RpM7Agkq/tBpG3uL99b/KNwXrAYeY0CoJLQ0yoG7akmPh
1B3UiGMTchyd4rB1NYGpX054ccjvnV3JkkpS22qERU9CqwcVo4TPk4Wxl1G6
B7izWABHeUNL84qSxcEeBeB6ZRs9he5Wk1G8zh2Z5ti1DRPx8mTqSH/P8G1o
sM2UnApdsZSK8vgruV5ZNLY+H/joNiNT7KEwd1+DYEtL7lzg8+OlWk+3oAjN
o7pHBb4tsGGxWlXAfz7IMqh2lgODNQhSK2xL+cvB09QpWuG3jd0rpiZ6CN71
SgN9wb9rfOV2vnODBE32/jEH7NspxjLjeicAr3W4cgiARcJwPe67aK2sLHC1
hVpx6q9Hyz/9tu8gJSUBO6L6i+wi+mnDtFah4VTbw5WotDcwjZhZTv/MmIa/
pctAlBe5UdMCdFLmbORFVcuOBbGoIIlRSOFnL+v8P0j5tORcq+bkSqsQHScz
r7zgU0sQOEBsJ1mzmtJtDZOYlq44wrX1FTHzLcwicRiOiyXUreZ3WfOuC9kq
cmg4OZKQECS3gh0Zw4cummH9hbSpMyCsEv+HZzsjhtGlPkZDZXoFKOLk918/
cY2sB8gLQ7GVNkQo3jzOrrnbK5Iiqe5bYIXn+8+Jr+lCHxwv/OlbDUuefwGJ
o/F/FQ1tFCoEL04LQcyVoyVbDrMN3icyKAZ4iYoJg3xnWvC5oTwzs/FBPq0l
GJoBjlTjDkkPPfnna+JDuIaFvsyd3BoG5RXk1osKtt19A7CHk0AzmbWH0JD/
Q1uzOD9oHt/pxNfLOklWshcWS0O4nVZyNBJ9xXOE9o0eQxDXsn6JEauCH5bq
Lma6SsL4Yu3d+uktDSB8hXvzS8qlpm66kPCS0aBng/8alVZnp4Yc6IvmjJK0
YQaRjxoOdv4yvf9Q4LEEaNHhoCZW8WHy8dwS5nFBPr4VKS10fxKFsZKKzu5M
RlvDIsTc7tyHf9+YOTZ9v7ztBGuRueV8DIPtgitv+iB5xTCyacj+EY0ZKab2
XjqVV8BCGCz2zWqwk9hpmkbhuPIkXHeYPYPQMPE6mfSzg8B3Dpap/MPmyLCx
zeNtQ95o7HQ7tX2/gkXvyHMX5LOpaDOJdLAaP6okAlI2R2WxKrDmeE0vebMw
JanBAcBeOoypTgxFI94ndg7ax+/tQnE5IZS1SJ5myZgZPc+V3YIAMBy2qmpM
5vfDjSDexlfYriG+kcDFYs/6ztRLCsqcgiOIGEjyMhqfQam9/5Rx6KKy8G2g
sAPiLzokSeyzWdFTll+i7SkZVHFVA6sdCyvSzad3t7A79foU7pUIzWk2CLqt
E/fO8Ase5oUPoIj4o/hQHy9ZHuUvmwa90NrF4enEQTiusiocUVZYji/Wu7rp
97kUpapTMEOH8KPFrvOPsVTXWCWuCYQdHxQkY9O/dXLrtYPNsf7+fqGj8kIX
UyPNF7WjTa7BpF4xdRfpSfJOJftab4+YxtUIp91eTNv4zdKxUgYWqZKZxzPc
7282svTAycR+RsXlWntF1Ms6TXLi338rsg8rE5AGMS8CD2vrsWrBx10J2EBi
uMA/I8ntiCd9osrRELqUpb1TCCIV+zo02XnENaqPIuPxqlL5q3hvWPcL1uOM
4QPNgKRT/O6F1nYcbM+Z9CqYZj0URIP9dsMM6bOkNA6pF3Bv8cu5oQ8ZlpEP
QvbcUmO9Q4YwQUbQb1TxWtwIvCJK65BWtyJUPiYXgvKIXbmZqb/k+Ag5wswn
K9v9MMMs1IA2NYc+ZPUtwSFaYns3U8nOfUG/oC87BzB0Nfx63watjdaoaqoW
4S3eoUlPSZS+vg+vDcOr/HCclSmvG69GHX5ID/wWk/DdoMDHT5xgftIcc9xM
tp/R6TlyGSmSKwFnQqSdL7VdgKJKCGPgn/uR5hp/WwQmpxbl46+wBzLbK/Lq
8AyAwFcoryGXnu2FA3DvNDknBeLVuPybUFQZ8U4w3BgJmHW795vgt1R4ubCK
cc3i3FIzz16azLg7lIFKep27YMAxilgTkGwm+ornlM7LRbIzMbzoF2gzG/un
t60/Pvuo4f55c5QFcsfchR26baKamglW5I2rAGsTgJ1lq4qVBBrvvTIMQNyA
TnR6xSDgTmjDYCtT9aEBZjP8hwcNj5ZlF8fpGc0WOLvf2mmcY3OjmdiEMflf
BkjpAXYaA9cLQeKy3VyvgmArGNmEZZXUb1VYKImhDWjwbfQCwfBfSl4RZBkl
1Q0/E12Kuoej3+nodZShTSnqCbCAqin6wFi4+d4NX/o2KVYVMyP8V/esu5bd
JjmXBBxApMptfLWHKUIpnoic72PuYibhA4hEKClqLsYCKQjGELeMwE/gl91G
VFL+tMFefzkied6khQ7hfwQUfsfpfFmmf0/f0OoV1YQviEJENYhjhWRSwY2E
xHpPbveEqb0EzWnC4AzihFnbrOKl+Y4oBinch8K+bL/VIJxs/BlXbbA1fHec
fC+zMv4FeZV1gz4MdjZ2ZIQWYCu1T5+izKNGch+FsKKv/J32/qV+lb5Riurs
vOinH/cbFReeKop58fe+3LLUVXQe15iw6r4c625U4gdXOHOtB0iXYZJHZYmK
wCpf5b8p5VY9OZ+Vwx4HKI0ajf6vlTDc7pTLhBffTqwAGzQZ4MihAsynX8eh
q7IKonmHxWfnsseiMwznsChkfORBstJ6YbUKHM0JyyrfuTaYAcPbo1i8OIlM
REvWRxijJwx/cNjWvnzIb7F+XtXzdBSRDdZfm/F1wAt8wXW36RxlRS/xjqfx
YPFxphnkC3hksoqmwyLDwWUXFLcB7cpiSPBrm91gVzTpaK/XshrIAOyBK80F
0ye0/dM2/u9N25I6pf6W18nF4xZ6p8qGplipytxB3CrbNmD6NBwLPnPSBbuH
NpYYvE5XJuJF2Qt8wCQ/1TRS89BEf7iAnVxjkTI6dAm2O4jDYsbCjaCLbX2C
7CgFl4J4cmS1tuo4ZNfHuAvDv1kRntlVnj4TjtVYcOoo4qm5eWOBTYaow2i4
b7I7vx2RoaiDt8YnCJUipyTwujZPEwgeEQziXbf2UvjZzyoQxEZYhjC2kKyh
YFNGNYI/7U2mEDntm+INS8dltlGmPBwHXlXQrrHUzve2hZTSk0WiPnVJera0
oXZpD3/aX7vHT6l0Y+FJP270MzR64DLZLxSgu3jsD/gvRsFWtFPYxenHaPLh
S78qtGOcVDRA+G45m9xcCuheTm7U1m+1IAnqINl7wfvFgKb3DyAlTZo8w2Sx
QhhBPkh2bZ13rRJe9kMhUKmh6kyVVtlMHtafUHaC0k6KC3YDqka2Y7tRjRHg
Mk6hiobAcTNdUScjiZK3HR92DspwleR7OZLgAx49gV3h+Dfl1u0uQN+dqjhZ
WXeu6PWZnFYiuqDMIo9LHfJSafDtEwxkSIiUE5qj3FGGmiVtjxhI2Kc4mdCN
Lezjy0ruRFMRX+81PpSIfCQHAmJZ85+rVFfSb/QS8NzjcV4yP/UaLzkEizdr
a//AMlgCE1x1d3HdSSl0nrW2XwHTPUaN6jealpTIobMiuf+zzjTncKjG1Ewq
Pd6K3882zQq1aFnub462+62GekbhRhQeAfuXPwRmzx8PGPE/eTZgdFGIfBU1
YlqtVEsUJW7WmWOf+i90HME6CGpObiy4OYrIV/+BYqzOiWeH0bpS6TUQxKLJ
Nc+UZsNREofoSRE4tW0oQ7fpQ6bmhO0GdKkNVMiHnw9zA60vXYLal7EJVEij
0OSqF95+a7GdqSFZhVUVZhmJNVMmUl4jmnKG3SgSx7jIi0VTzFJ/77EmhhPC
lt5BBUGrt8s3PLO9PMqPnMgV3KLTos3ACzGrFE8duKG54m3i9k9O4slE2yuz
1+z8xxfncbbpRywttGCrCzYt3U333VYwhprR4iWM+p1lTf4NQjTA7bHTQa8l
TVdDwHwb7TDZ4qB6NCtZXr6eKbwtXHM/L4QzMTKUnIatAcTuOBIuhNlojT21
V0pxstY7KZ5Ijm2ZMIAq+MilcdtwYLTog6AzJllpzEME4yAFdBGE235/xmPQ
CehwB/NKULBOX2E/Iia9THb35wr6EQaHJkfbABcru/UVcdmhQLlFV2fmjXYt
tXYXR28VLzATyoW8fKqNOEk8Ujhpxah5gPdK8ikc27WVugEPqcmnebg8SKFU
Q/yH/OYMFK24SqFsvU0z0Bzehb9bHpU0GT1kUt9tqrsd6DeuKuP+6DoaGc8K
77sv3ScIwY104qXtmjZd/t/zLTgXwdvQbWRzjHt/Ycr/gmU3rspYkR7ziQen
LlUVyUAeQDpWP9lQlWdm9xr0MIPr1XGp4+SERMBu8hFLLmKM/17nbgFzO1JL
Cyf8yTpFr8i0vy9bF4UK3fgQ0mkf8o+fzjtDCZgyc56ewnYZWFfiUVMaxCcF
J8K4Ut+G48+7MOkqh0JzOrmuUCmpHcEpYmmsYaWrQ030ODZA6QU3ajyzmdqh
dgGNpLg0+EIGheDq72+CBnPJ1VOQMDbQ+QcHlmEJuIfBXV1lrvWTZOROEi1U
upRYTNQm6jTcZMcVMIq7kROq+4sKOoHhnv4laA+8rmprqc3nE3q5t0v6yl19
JU8rOthpKEmG+Qyeix4bdWucqgZklqrsBHv3Ccpf8jdwDt003CD/Pm+r9xx1
HJJx8pjW59aW6vMje4vdr7pMZ96/kWYkyYXNQrxcrKSvHBO1lJsjpgwQs64n
Og73ouGm0ZZf99YJbA/rvNaDSq5wsJa/zjF8AtUWcli2RetCFychHlpCLMac
rn7K4mwEw6urDkV0NCJLyN2G0w7XMjkNz0EIBwl7uUWCFesftrJmfbu5WkxR
LKBvJ2nsc9Qz2B03k+YnT9Yqtt/8RgeBV/ocam60XbXYfcnvgsvH0LPS/7gL
cDfZXn/rBSfDDQnMLBed7lWRv1F8t0ka2//lziDtzI1Q0D/LXikE0ccPcJPp
0Rl2gemTNMUh2zvPXCmBUTROKwIIxj05tnV631EHc4u36vpIK+ad58Jz+NgL
hdXIdUXVfPnwmkksGtQk49KxDFaz1/klB7TcA2Mep8XrCOLjIdNwfcsBdNRs
CcEHUwF/dpZY8oS0lk+Xplqw1e1dKFkRDb42HKR7lVLAyqWMbW2KpYmy+0sL
34N5dmVN++KntlXfN4l5YidlU3arflvCurrh8CVfsUX/SQ9gvDrgXY+i2kfo
mi78U2MsLRmcK9DyMHkFIarO7gb9hT96OLXrGY3fjvg41Qp3ZZsx08ArsiPZ
H6hyR08Re3Z9UorUHrKKFzWWJxHSKJ/35VUCYevf96ELGNVrODrvDzQUg8PI
yuhTfe0YjWT9E7W3HemA0KbPxsxQgu+5zTOSfaU/MP8wGiAICGux9HYKkVkk
QQz8O/up3FqCpV+CpeOLJmruJd4WzA6nZSfxxk24GDNPPYRHa6TF5GuXoWhG
gw4hh1xK/aNCjw8ByCeWTx9WJF0CrIksqIBVWX3s2m85uIipdcV9gOJm0oIk
9XsH78bS9k7xUY9+UVF+Vz2OprWVJU3dkdxY3lyBywPt736w40ttGbSTdytP
JDOsEFTQQhQhgnnsPzSKkaQhUrUR8avx0nAo1HOG5XyG0iJgIvBIptv7P5x5
5z4FN2DQG9V5v8nGoYWMUBtMsJkuOv2c9ntJLzgn/2pPYVGEt4DE4SLB0B72
GWACYy9FAzX3XWPbZwEe8d/U8izOo/cl8E5NkOOONV2DeogVLNnHwPuxEDmO
vk0XDavnPRUef4u5QWkTEO+2OmNNHg56Vsb3KAhGTxnVCbd1rrl/NUTq+myT
yhUxVe19VLkxwOl+LChFlsfYCDruIpKGVAB9vlxglsBpdfmHzUOZt3+dzh/S
mGQbZeJif/DbFSAeBQ5TsTnlnSsIeI+ouCOSh7HqinBVcofBA45NjXRAD++U
HmMC3ewL8sCT/dPcLOw0hxT/pHT+PATJUX6ZI7GSZr0z3B6E+UYezed1ZMfM
VK/7d4oe5qbbATHPtJYZ/yehUZOsPHyoo1dsoIUWtvqXHJ5YPkuTO/Qnyejz
nR18XakmLAkwYcdi6d/YtPle5iKAUqFXgEAVZrOtFYSf4S7l5K4JWTfX0Q6k
a6EsIFAz7CdvRh8KXdrRAo3SZmtqcrNBDYQ0hFRtg5LabftiysLFcn5SBC+4
JHXJnThMTM7RI10N7NZ+FJUUerWVHaTyFVkreuq352agMUHZ9ujgfE8u1v3M
UFwbPoA5Uzr51tzhv81P+rZgr17bDSHc7BuUxq/5UbMjDhdtvnpmqQsT6w6H
ljNzVHBwFE7zzGh7D2HkY1AJbiCX7oAZqJ06DPnbBD0SQC08Ah9Tcy2J3kZo
faNVHIOzWukjp8dQpEX/T60iN7CHYX5xd9sQsBR9jynX27pT6sd87fXOx4Tb
0Doh+D8ZQEpOdERl54nTRb0urGYF7m9IoQBu2WlwFqCXYsaFXNVTE/+wIXlW
kVJxfgxmezMaybhkb7OuwKikQqYZf22wQ6XSw/q83Jr9E4NZMhea64BhpyNh
H6Wo+WynHtQ/J2G5VHCQKNoPcuyHDFJUZtjyTmYemCD7q4f4C5TBsAkHDorH
iXLQtKyHuEvVEzCZMfZfNrzXL2mwLF4CmBDH7p1iJIMLVoEMp7AyqF+7PXh9
PzSMES/rsY8BadNKdrn6ahY9qCxKUe7H2LV1soTMNslq6p+9xjUk99joGmht
NcDgT3f3QjjsB6zC0w68g0k7b1FC+9cozu31ul5H5Krdv5WezxWV15sLwCET
N4H9BrGz3xA1dMBzQkgFkYjk6nE8bhNAQoGGfw7AYPSyazdiGPWZSh1/60di
MsKQW2C9qKBAhAf4hyLTMoEBZegYM/xEyHEQz1Ow9BaeaAg+eN+xRnFip5o8
R7YMMIQNahJTI9+Xdf/xolOrgqCiXV4+EgXJyp8Kd1FLVzhTYc1atz+iyyx3
LRRr7JDU1K0ffbpEtMnMAeTiBabZSNUBJoJXufuo3Gs0n6G1q3Rq2QiMxHE7
00X2jgj5iJR+2mnZK2pDK/ObxjvJIJexLJT1gmUsYNWzTJZb1m7vMxViv3RI
Len6xXQtYhzRVYedqAHZzU++Mwv6HeABMRRQAohSK+FeOwlv17RMaJA+InG5
LOBOhNMMx05indQR+qMwj8XhawUSzmTtFq24IkJ2L46dqRdoqO9/zg+4Fczl
qz4izJK1FB8AXhM3Q+6QhtjKh9vEAf5zW3pZ22HcRN6cdXd5REtqVGJH364/
LCm6Rc1xa4HJ/D/WStHT62b5dj5g1cN/LyA+PXGiRFrcl04AO3G6sWP90Fzj
oQsFp3WfgIdNGP16OQ9U33EUceKZHokxO18KpkcSSA6Z9K5OaSpvDhFfRau4
QD6aSAfMsC9Gn+fGzqGy3fIQTPz/+EXULlXnrIXrMdcqnuN0UhF5Sf5rmJ1H
zw+CDuekTbd1OXxsyYXpJLWRbUaI53U3SYanSsDcKrZhhLkC5S6cSNG5O89V
cjXojdYGVdfR8rwKqnCQ02hP2Vv6IayuTyoKK6PYK8gtOpHEm/42mN5TIVPB
1qGGV20yj8Flk8tOddXwsm9dBmeeMk7BuXw7nfE0YiYxMq08DjN34bO7DJGJ
OGkFoooUflhbRLL+BVxHkXHQ+sEAVXHk1fe/CyzBh92jm5H4XtpTpeINYiKV
5fPS9kW0oSxS+WT92tP3gbrxmn+71rJNrXK3smAofq8bRttg6uHKPmteODyV
WcEv97y6w9UfofvEcvnmLZ3/AGVKMTO+yxEv3ErulrEYjaDaKx/o51496ysC
FnooUgyZfpxL8J1W1j+mc11O7pxOWrMcoRjtuMSTrpEQkWhYMfn73S7jbwTj
NESlHDK6odzqlaQSqq30hQq9Hwq/pos9gZ1k/l4tEUkfQyMQ0veLuIyQbcIi
q6agTkrOnT9zRt5qjXyzKASy8psSnloJmMTvcD4V/xlqflglhjvDP2CrOBXc
J/fFApkRWq/uzQthssWLs+Idm/0sRIR58u8kbxCXDZmfMhcrMQ2FnjTYjjZt
8gavJuLPfNA2hiR3UrL+sXSSAP1ioYRYdRT1Wgvz1jOQaeAFuW5SVxGT0uyH
uPoK9U61KM09lwQuK9fTwWTkKk0aRV+bnkAQHjot3rRwYPaHlnQlN36vGbPK
1iObsOpTp0JyShxJZ6MSBkWUN0buESyt5BMFwrbd1wd194yLE5Mto23O3u9c
ktkJoOocixEaX0PXjZSRvmEsCy5piIn+/2l+OMy+2ZQzc08mVaF3pkowNm3T
WIg+xPE0xZArwG/ei+RkmAW1LwPaOzripeZdifQ9e9hABGSe369QKPdmaa6A
3m/Q+v5f4EhP3nDwW5ol1zCutxIsdFRAbvU54dVtRhPOVRbkRQCbP3EUXYhd
DVDnWRzeMTd+wWdodr2T0VxHZDSEEnpv8HTXVIBdRaheex3xrOBjfKazNiDo
wawMrWwt51N+f6TG2ThHs6+Fe+ePh3IBOfi3Vd0bE/AQXI2f0IGbVhZM/ZLv
36uimDBCWptOD5/LxidnnUqOK8ehUK9p77DTgi16QQq8+T3rVGUwWapcWJBk
fEGFJ23CwPkt/gybvrbmgtuaIcTVDpHP3Wft/pcHEJSSQpUyoDGiM+w2yjGL
MN3tSn/ZIKYVisDyt8aLZDiMPsO5RSpMaFCK/b5bJPTuZ+oXkM5sq1Hpy8/1
3W+If2yoXXrekpI+nZa6irC4Rl939wFdCbB1rXvpFTmocSydcgWxoqmtrSsD
+UxuDtQKY7bjriKGCmreCQxfLE+4RPkKTz8FmAC2pVaII8XOtl3yVikfzThu
ncmoR+gLtyAHeHMIurUGFeYInovs11xLBt2oIdicTXLHWWsLKF6aKczDODN1
t6hKeIt8v6alV6MNsttsz1NRvFhZuEriFSW4LiQDchRC9g6Ozk9UDk5g42iS
EYoGo7fgfsKO0CCej68MVLh0c+GOzobnDH35QKesVPX9YMfE5CpDEyBCGmJG
/BS3u5lf3pJR2JRwYu7w+jDJssamC5qrVHxfsXIJa4kgwGYKnpvi0acisQnq
km0+XePNJRvnBoe/xdkoxT9PT74qtzK4KsoACLhS8vj9v0wQIWhs4kjw4f1C
AO4A/Ny/hs+8jL5jlR1hZPXmcaEWttFqnMwVoWufaAfy054a42ChfWOhD9jj
Eao7eZfAVbCUKQ3H6gHSRgkDttwW1/e5vH9VblpTW4YYAD62nOYlQgcETu26
otjHb9fG8LoIdJm1KRAof0vWB1qevV+JgXdqnKGHICuYTQmkbNE+zzJu8+Ta
L1y44gCpGuvSyLJT9zj0oqukT07+GyTt832MWgVdQrJvv5LHKQmBgaVlpiII
u2H/UnsXYDTEr3g42c745wgXBNzePK2igIvVHUd99l1jp570OJfkOchW4UU3
IwxhBeuEdTqNCJqNUrEyeCNmyeAJd8fRhWJzE+Vof8/CJf8qxMpy2HRK5spX
fK9BGXHLtDjy1fnhSWvYKWyP88IS40ZAIBCePfZFX8bR/23CWtDop5RBMkO+
gWDlcbx6mQ0YaD5CF4KoInuuaFGGw/H1iMH5Ivht2dGxp1egvkVFbcHjMxBU
QU/NlUAoamusiFWjm0Oj+T84Y0JSyRVXjaRQPrCMdbuTWLjDb8YJAb8khVWu
OJbDTyJBR4FyxrB/EFJ8T1YLV1cLhb0EUC/QfsWDN2JiQgkqp7gcJEh9UTAZ
ltQwE7Zgmy8heF/k7AqzXgykTFzDI5kJY5ZQtcM6weMkTGtqNpz7UL9oFbcz
iqNzNeLO1lsYgFnOiCYuaK7cf0/9KBek8bBmNeYlp317Od+6hwJQIux/FqAJ
tIkT23YmnQZoIkVEK2iVgowFaZEvZPI5dfn5LGvjWrVosifMMISKQRSG7NlZ
dhAnnO9+xGT9pbDsBVIoiK7zVpoJs+EUrK88cxS9su3X/+HJdWKVV1mA/XpA
Tbm/dfWKu62LgFNt7s1BZWRKohu4K1PHOEi4rqQqAwwEs+VryvcaI38QzQAT
dKf9oBarEiBNxd0sVRAyzCiiokVe4qNJTrfQBQEYxA4UiBhLzduge0eH9Ig6
+1lCqBfdebQrdH1DisBv7774iXe5w0eL1jL8g/GuOza60hHfTt0kUNF8k/IK
aNem9EYGChsCLpL967fs63jAtfRTpO1jO9By/YrDIBAoYc3unN6+71C7h1Gd
LoFnMEie+tjT+vKfvVZsxLVzXigRMmiA71L6qtSutad3LyVMhW1lZArKRvsG
7bPlGR7BvYGNeDVyLBiBk1+kLsj6vVMkikI0c6C6GZA21FF0yaTwQvUFSnk5
0nfkpasqPty7D6Cg6dp+RAU7bO+nExtyVXyM/pZvo3mVvRnCYvIpSSqwm9th
5GQT+ZcWDlqDWdWhWpf8/SCMsBVELmtU1fEmx6WY5KvEqaDaKyhhNXj5g1mb
bCwxRHmnOSDOw1BtOA6CmdG+WSF6G2yOSMUr5iDXQRzJBrBTzkK3V6nUF2jE
GJdmlpkQnFA1+T7PwFuOxrea9m7hW/zH+0VtJxPdMnxOtawqMSFmu/En/657
Ign75Sq/EWcgBr2xKV1sFIC7cF0weWoy+pDG5+aSAH/+hyJrM1n/aSusX/J1
HHPOvmo3jZfqJ0wCirAFdF6l5enTB+Ye6DFyU18r7CHUyNqVjhGOqoJ8X2cb
R0uymDNPj0BFtmAHoTfnJU5A70q8IA9IC+0CmbCIrm+2tQNnonTGjifrgMvO
qBYL5/RGVBAqSYZyPXEbz0LMLv7qkLIWLVC9WADVYkOfqSc3ehaNAVsNRYi1
s8SpBQDViCPH8d1B+QHOO17cBm7WhaN9ToDQh2PPMP9aTf5tpY8S0D17MZTq
xb4k0XyiLAU5nzYxpsPC2/1OlQl2E7VPr+9mY0WRCXfX/Q0gHk1bOd33IQhX
1ITpzqEn76E1OzOyx+mN3bG6UQRlbo+SOwgGmMMxEMWZAzm2edTuvDVh0gtt
3VDnAS496o0Ygww9jOm09oEWtXGJYiVc8K692k+I7OrL/CVLIiZAlZoCs7AC
vSaP5iGdgxG0CDIiL17ZTzePpeufHr4f7K9QwbSTagmMBpgaUmEOlEjP1se0
7xA8tlwTdUqlbfMKSdBL368fsac1J4O8pKip/Pl8ukZcsm2psfake0LMHi97
2b8yIorMz8g+bdVVeMcFG/3A2mUfT+cNCPKMNpmL6PNgeuOlaYkg6kc5poDh
bBm3qpZgOtMSJxFFwq9wpoy7M38+cRqt7lP3KHqlsqCCbraHBXfvFDbh7l/F
cj6TI6hlCFer1U/rgDCR+v/ntHzRHYTIAxRIgD5lzGSsXpbYOzYUABvf2VJY
Sczr/nN5YxAXvtdIznRJC+/1BgsF5LxsNkf5+wcHoLcfzMXieoliQfWu0oi8
B6paoxKnODTo36oytcexnIXDM6FFHoRsNr4POKgX7rkbVez2mQz2SifHxc3g
AVCYyLkSwBIZCcZ2wWUn7aSYxvlCTakY/9M0ZTqcxrTp2MzB8sx1NVXttunu
hp5OJcR2rCA/glqTP+cS9FQjwwlCuWgNdtxdnGisdmnH5miLpxs8LffYMDuX
rg5eZ7PkQMOfGRhfuW+UuD0Y1l2wxJJtlF8Bqs91/6J2r5HqMZz38O9eK/Jo
Bd91vMjESNn/iOqKsOOlaW+zJz2HvvrXFTIBsrTIw0GZKknIvU1hMSgo+rp4
d4qDcSlbv+18Ae6FnRoneUpR18ugf/x+fRYL3Lowu208kPP4ooMl4Wv34T4v
R8qRayQgn6nUrpAzCQ+tJiw0ru6kIIX2hr1fIoWvon9lGWFuzBGee9tz4BFt
9+lbXiE/8FKyQx9OgvoV22CYnQ3kJtzEl2HBKB84vofllUhVFrW7c4r0p7/1
Bp2fpcVDUh6vJIwDrb3d5PCEVcfRNVgwZ/mHeqYFXJEKgehVvcYNa/vkIE46
PGuT9X7Qk9Uu/9NRWTqM3IbLJk/YK9tCCbaKU7qvi4ighN5QS8frt0mAN3zX
0FKQnWNlzrtKGi48+1cMXTwJE6KYwyZVBjU9Wck/o2Wmo1OSW5vFP1jx3U5Z
1KGdQ62JhW0QcouKIp3cVpkqolUdr5V3gMUy8sIwkoRMS+5oAQqKILtUamPT
k8Di0lzIOAtHsb3MpKyw1slWC081x8Llu3CP7b5Zxz+D/7k6OTXHoNJczzrY
IGiE4ReA1ayOk71iDOjM78YDwFl0fFqUi+BvSm5jmoH4cEQlbPW7d961pc6y
k5809pbzBzAPR1kN6SYaUMn5VVXx+AQzkdCZ9WoHkxsclGySu8L9dO974Av1
ZKhRUrym/JkApA7zNf1aLUB0ulKGu2XlNVPCmtGk6o2KVMXZomLNiKxRqTzo
vhhl7aO+8fcFis1r2jIBxvSlwp8RCIPSavOBDhwf0M6bQzX202mbMV1VffRI
JKReqiTsJZVR93K4EYKt9DicQzOfyLMggYXjloqZIPfeoHA9mI3qfcgUunsg
I1p/TWSjEZp+it1djXLaMOsTK7S9VZfvWbubNdIOmcqRMkc/dkvtBIWTcou6
SFe7RFXqs16+AXOHNDVfrupuKogX5CcypTR1ee/oOiJZMoPaZoigSFoTYobF
sHIT+5yVNkxB8v+ey0spXfHydRC/gEtg9ruX2UqZnItgntOoDHrg+wnT95c6
ejFyv3U36YGcbrlSq4vsGCoULqRRrABaNKawKb+JLzmGWgYmZSVmvEe8VOYE
wQ6Vbu+W3C3T2TOpIQPEy15d/9+XBYWTy8RmSjGzVMzC/z4DY+U8Qj5fvsiO
DywtOhoJOskNk+puNI1PQ9gNjbRbLFcF5SVjsKoIPnLFxNq+oPoYAdcmLcFt
EtO9WNfBhyPD1NLBIqqOriyvtLwAIjSdnHW3KAL7OL0O7CR7DrLL1S/Uqn+p
6tS6u4Aqk1p1rIxl3yPxwLdda+kLTTwrUMMIwL4YNebVoZus0PXqGlDWeNoR
MY8IC20XA/N7hkiFDVFCesHBZz2UPlJIR4aOpsoyjPLiSfFaW+vj1/tVivDN
N9FPctPJITFLMRMd2MjOf/3KNLINEJOxalnshDtl98i1ISFVIjNt+T3nNfM3
fjOPogNVkNE9OyUGr2Wp5BFn9z0bT54viLk9E65JzrtNrTG3tCmJL1TlA6tq
7xxWpJneJbXkDuSe6iLb6jT7LJ+vVHG58bcbWKiRJUZP0eJboxngiK787vl5
YpIcdJVaUq4VaGg8zPceTcYB6QGS0wAuqROgO/irJayo1jekmo2q2fifMVe+
Z/v49MaMdDx+Khth5KdhMpgAV7LftH4jzV+xOMxjDf1OqCHa7Gt7Qt0NEDdq
HRJg8YfJ9RWIUaYUiefQkqO65bFLTnr6CPWyS6xv/c6O9fdxhqHXsilJSmMs
XVaXuDAysbQZKlW3KaZuVYZGkRyfJy7y13+C1bHL7rahWspvyJCUDwhqdMzm
E5RbL8eJFtLptIU2cqD0mbWR3z4H7NQVK/s3KvHzn9ASCLx4znqe2R3n5i3L
+697rU8rMAqOzh5WEdVM1AOx8stGWmbvA47HdqOLRTuXtZsALlb0iAK33dpz
SYJurkO9y+Dp+4x50uPLgVimL8SRXcETr7N/ItS/u7v6N5SVtfgvQSqK39N5
SdBD+jBj4BgUWKhOa6YHdZcazJZwK+pBgBGKVDO+OI+5USaznLKfkXFqCTPe
uFVAfBD6JXHBC5OFrOkowvGclMd1hdZwfOef9EccTKVOz2olkSVz8XX0BKSK
U3pVT9UaYWoo7gusGKtecgm08hcPaBAc+cxH4PwI9KHVg8IDeRjGuWa0iTLD
qNr1FsLo+ti7kZKENFozRBvC6lMGRD+9q+sE9uJv7gMlgP6JEU2O4Q3b8uOS
WqogXh0TwY8o06Kckv+YhyEDZ2qQjkSj0Ffl6HMRXTqrJxQZAh1Ez+ax69bt
iKtK0NfDdpYM9TQ5x1y85vHDDLYSSPjDVkYvZpn+lTViHSiFgbUeud/xlXit
1nGXBVsK+3dy5IcE9DgwnEAE0cC5kOGI1XtruofDgcRahpWX6NIaNbcrlI8Z
WPvOtphT7iv5Ca3NYZUZ8ryh7t6szxlGChcGOH+GeJdW8IQaRuGDBI1SsgbV
Zi5jKdxyyZgZ40yfVJHgJYPLzm6hCH2ZNuEDYDnUoAnXM9v94X5t2d/mKiWe
/3qme84tvVl7KBEOrjj5cYltSmgjiJ3e+ViIvnrihfcGnSFgTh6uSetLcS7/
EdGip4VN2etDDJz6VrR17piKreW/E3SvQYHuqzBL9DMpLjCTZAn68ZZarwTW
dYuYQVR2+oU0Azb+OxaeAi/OSgjszE2g1X1VsAq/5jm9n/WlyzQw/j4Tbf35
fJKkYittzGMfF1c/ZYtldmZ3fQg2YJ0Gnu5BbWoYeeODUTZEwCcZHqthYhK5
M0FVNuoL22DloXljbCFuxcVmRhIrVnIJ9FGb18CNUtxHuFObmCnj0p8JNLSE
SfSARvTYGoWnWR5Stf3BQghavx5I56XkHxz82F2ImsP9tBSwi8+Zp5hDxVqo
+RjnIQTgozjL89lfmzbfBULERyX83o4GPKHPnXsOOBmMCZyP9vewxnsEI4hj
A40BwEQ/olYAQHmHkIH/biwfTtC0zThMjJXf0/dlz1KmylZXrmcbYjqSiGMb
wVedfNkkpfJIh3n5OcKocWdvTCs3PITqV/ya9QS/NZqBGhsUGPhz/rXw2tx+
/ihSZWZBcllIVXagZG5MxpQEHAbmaD3EbM+an4TaAsIXqB0zrrqwp8cG+4JB
abHiPoB0Ne9moIEjy/Awu8Ik1AAbLGGDV1TRe5CWoroHfUTLB67PrGHx9Pph
sUCnrisjnkJ3BB+C0s2mae3gVnqn6UmRkxEWEQaFmbTF3G8Oh6LdE+hB87YZ
4KovS1imYRUOklZAcUrzGL1AXTYpF0Dvi+p/Pw51sQ4VosJckc0iToKup99z
otFijQnkuy1MT4QZf7+wh735rzcxJnUZ10WNRj2R5byLfAsdeTFMomBL7fTZ
zj8jq5EQi+Gi003iUPIlYEYnxAReHkXPi02pqe4b4xEPy1wDv6nNQF96tND6
cINLZ5hmYONdxYcg/mBuTHo5W4mVm4w43QAtzXYFsHhjWf502vxvs+ARiTfU
3xwlS7/hf+pSVvm0M3CO6WcD/E0Z/51B41C9ohnUMdTpVPyXmrRNJvb4tf1J
/LHvGjRvfWzuDuu+Sb1r6uzY77Y7XRSEcV18WyniOunJM783bBU8zB5FiNLW
4G5RsYJbq7Uoox0y5MKo5C7Hjidke2C2O5KzzWhRH/fGLBhXTC3VDHsyodJE
06a9TMEh5nmx5JpaMcEvc3ZEw1tEO5eVNprJSaTto2j/eVsaqFukc/4v4urM
FXXbC7sHIIUbJaOCjXF8mT21eIwKUke/fGk0Z0CSt1BiFHoyDbhevsRthA51
sA19pGivS7B6Nt1zSnwu/jRbtqB3iw7IqZ3GuuMWKXQYLD3q9wiNMBvech9q
MkPdeJ4nt0ra/OrxdHNvGy2C8hTmnrBitLwwzumOjfRH55t9+k4EHjXqcyj3
8lga7G6/GNqh8owdR9/2h/9WLlP2Yc4Z+z+KiexmmhOxnToDRFXR+ZdPGhjF
aXoSacQiKsytEKWNHnvux2VsH8/8K78XGJI4CLg+HwThfgQWBof44UWUQxAs
N84eVDTqaAKuNhqalVF6oy7zUVxznTvZlV3SMEIvmiNCmyTrxpAxRTf4aYqf
gKa6ulQl40ezcXg1enk6XgziABLQeeLS63sAzGox5/kTYpmyDevOXYSYncXf
zfe77duZVmLJJt/wRO/S0zfAFL0U6HlRHcW5tGHGu3qiHbxrXhIPoD/ciHFM
U5Brw7U40k8Soeu5NJvAYF2RS9vH2c6rX1GkAKx01+TpTjWNCmmOavkfg6eW
mN7hjtzt1ga47MzC3uJILFbqWI6TyW/l7GpBYWTccgT18YkutTlKkXIMG014
bNEQ5sqi0uHLbq+Z5mzA3kR9garrALYmCzSqgyXA3Iitj4Elac4aPFU/VW/Y
4Dp1uJx/wKObKmqc05cZnyaBC4L4eypsTeLpNdugHYxYMOeJ2BPrVTMK2hsN
sly4ECGCM8ZvU5ED4RXkRocCQuvztY/OPFYLZFidru5vtLj2tuPIcyKFTT2S
BLqimZRwVIqyMosM8k6gsua5VqjjVPIwnZQ8baPr2ddWxTs0ri5U0K/XG6UT
4dsEBUA6wAJuVRXFPxJ2ZJn7SGvsPZns/rQl46mlxLOA40Xudys2AKL1tH59
xhk3DxC/FXaNq0Opls6zW5ZkqMu2g+BDfdJe8fb/1FANEZ/r7D1jZ4hfsj/u
1TUUPQYi6c8OPvZ2f+WO2DD+Fhf7VuwPHYLTOb3WTDZMviU+1MuLpwFKnFhr
AcWZWlGOD0J55h1VQeVdqVXB+dBejOPIbh6j4H3uMNYwYsoub/buqhSWYSgF
Se8PWcR1N7zaPp6CxIzl5gVRckqlowcZ1aqDzgGXLTCY88v7ewlNLdLYsQ4z
WG8+LqVzg5SiKDZQQSa/5+EBeFLVLjTfqn1ZfZ1dY2h5xaqV/cbUkcY8C6Qy
tfC2i8KiWnFWpiILftYb4pnaTI1H6VjTC0xs6S/QhVz5hzdP1ziSQKEkEvx0
wWxAfpnaQ9UjRoSgo1emcVxUKxX4SiGSkzklslk9TjSVOzVrpEyH/F15F2nk
RKjtsk8hiMELn3YEmiXcf2kNiyDw9TlZq9qrDYGwRkkRi9ax/4hilti/CZKL
etKgr5rh2SJ08dpqqXbD+sqypCCkT7uGuuEPNDIOIX5y0lJg/a7cy+98k9J1
iMhvBBtUou03YVbS6OFtYBH69JTacT9LM7SSbscvlwYqMGRUp0dzl7o/NcEs
hzPMIS0CDFapvyojiK9IWcQh/sXjRdcwden0Ajr1agJY28hgE7ifrg0gixza
cRFIiuh/q2HsU4RHflWaMQkU49PtUIxFE5mIbs5n2jvg5tymLLb4Ucj6trhe
06n0/o8d8nlR3TWLwLofkypCnewYvl0THxCE/67g/NQENcZiKaJiKKj1MQI7
3y3Acpk+gs/fRBJYOiJBRZxnXVvxQIPIvH81JeYdhcEtNdx7z3cCq4sCdbNX
V1xNZn06YMHfPR5tayRG5OPgatjBKrnHZ+u7soeQ9FdfOPHinLE3pwA9oWkt
bL9+Lbm/h26hB4MBQKBHwGtNvSn6NLmeuOJRP0uTkFjK16qpGwp07yrtDhyU
iwlSza4SzzLzyhTo2fAGCuKGgrVZF8frBp0A+c4Ypx0a9YIeJQ7G3h+xu9mP
VcphdOg7vAb3EhdmWLdte+myP2BWVoUq7cPJI6OI5oPoWP+wtGUxmKeHwJu+
QTfgy3dRGHTTNfD6MNWYg93jq9yuQuZO9+PuPSq7wuYrVXGXMkpWgcVb8C8q
blu6VFtM9iv9Jyff2YZYAPRnEIYTokZu1LoijbKnp1YTVqtI8Jyw7cqcerbc
f5vjp7chPDxBzsN211xZ8lqEcydMGzcuS1s+zv7FhOEof+UinQ8JKzJLY16S
MtKo0S+o9xKIBzNRLnnkurZi+rbf0BOZPdGN9DOWa2xqOJ2z/Pl30+hGETid
F7MxwfjHtuML8XpEdxc2uVJ5ud7LsyXjGfYPkyMLmfyIVC3/zMnK2U8tzmmj
ugpSK+18Iy53OBK2ZL6ApwEo36F8hE5AmlTvO3EHVXaV7/86zur+vj//fOj2
8g3IhCJH/NTwzNy6BBQ3FDlZI2yRWFRl1sEqwKh4aqTr0NfOlRGZcqgC3Luj
F/MBZPEm3i2l6YvQOWsRHpjvWEVgTvdJQDz9MrRhgp2oDscfoCEmNLx7efK5
3Ru+kZqPx0C7x8e0EaWFPP1PTOHxYgbgbMIQnVkJW3Jc8+0f77CeaK8b8d5C
EX3aOSvPSgSMryqpcr712DEXm4MB+8LT65Oy4/v1X4vebEYGiCFRLvq+PUGO
l5BjJDRcPUoI4Am8xIuU2E8QGIEHa0eZoE/rwez9DSWX+FWPq2YV+a05dX4f
H54uqWg6SptU/Xy1h8Of2r908sGXjsk7Qqm3X34eSS9ngqhnP+DjkTLoP0Se
Bw9QXE0ticwyQw4zYBsi/uyjlnxmX4lfcHTgXGuk3MJsSplXcXHGQKkchLJA
G4RdHKQ7LOSOZgyst3weEXL06+oGe/bQjWeQa41sgzgz+WxrRJwMEO5JJKwO
4qfk0HoKT/TETsIlILSE9dqsr7spKr+XISe++ORD59edW26B/Ki4hscR/gvS
Ig4jXFqgtpcuV1E4uQjZzB15A/O0C5+wJI/cUCruPvhpUc5JTQ+H2kHQzIul
BU2PoBnuheupC7vsFSMHO30ZISDBF/MRKKRPgPP2iAi/kie2Ou4gc5RuO0uV
alZ96T+Y6cpgIlSU9vON14tgKbOqdGMklmeckV0hPTrsudEcrF5WQWuoxywi
5F+FimWdhBzqIe4j/h2gooCHFhCzFnR2ySYXBwvbL93xQ4eODPkAtivizx8k
leBTuzzzIPBJR1SozIwqJlxr9vvq0yWySLzh8YdseBS3571Ez8F/n3opWFhY
Zhb5qmk/rNSApT5500QBABhI+PHkQd7V28b4laZIb+9T5m8NUQRwEEFdBsZf
p/DtFf/jnt1E7cgXK/vL/AoIcrsYp8I4nGzEh2tZglrZnGGA1Rjxs3l2dVat
U/QfnMbGwCnVGht6oMjZyjySAnUlx2au9xW3KbpmI0882xK/yTurQm9BHy9Q
JqkM5uGEtIsGQSUVPIert8F4mGSkx9mQW74LIZ+Ftq+nfbfDyvs/QB4pG968
WG3q9OJmHj5PpB6+8+4ftAK4KGClf0rl2FANf7KQksgTRM+xshArhgFskcCI
b/qOdBWE6QZV02r9F+E78eeim7pw09zbQiKXtpWSapEDm7DZKDOpmM4peiJt
9cb1mKBejB77LRlZBcxrVA3ZYtgSbbE8iOk8PSPnpRu/4gw7CKasEt2Wl+pQ
3u+SlRjwqBoID/ENY2R3hZiFso1imZQWdNMSptrh36IRwsd3z1FUkjG/FfzF
M+N7aZbJUTXKolXKBZn2x62YX5RQbG3e9PJLoXRTbK0m82/TyBkWzRoqXnkn
YpdL6eYUQ3n6O1+T97JzYB2QTo1FYLlxSi7KKCmhc6vYRB+EqDKpekNLaJGi
7u5ukwIm2utXSuJpou5qSbiOlLn36jCjnZZ7UR9ZIg8g2liefRfoex8ZS16u
QJI9PN3MDn1vWZ/mtxbKad/Xcu2YEJqjCYdwHimEh9pGk2uV9g6rESeJQed0
3eiYPQ7qU/mP1F6Egn6KzVWkVzFJs3zFhCe+D2egB0MKkrx7gXYEcI/cdtjO
yQgyEG47Ep60VFBxFRygU/jMNF+cFf76mCNYwxOoGO69sVL447CTIJcHfpH6
zABZ+NiIHYPiAN/nilReU8cSfmaswm7ky5NdTcNwBlgE6LbLhYpniMrBWRpO
LsuQ164nWhJXCfMl9vaSEaZ9sf0WMxHJLr7ubjjKUsJLiCWt6LvJlqddB7sB
+oxXlBbjuxn2vw2fkqRWp0Y6cpWHtTClMR0LgdRTEgdJ/BEoqVcCQJbvf02J
UBrzUUrWG029P7LOBt27M6SAhLSxvVwXc7TlqxNnFtUuQqr5/zQ4VXZBr4qO
NCIOa3fqdm/19WqMyoWQbahhpiLZOiCn4YgfadE6kGdSWNkcz3q76OZhkY+b
C2T7gjZh3lO4JH7J1TwFjexu2t4pv2WUFGxpfO1EQGWObGRfRj4DUWLanEXh
kByvGE58aN3wIizuGVNYumMBEg104HLG3Rmktqa3FMOgZ180da+WqjvWn9Zl
Dnz4HoyAc6quzO0gJAUldrC1hnu0QO9rSRB5V5q2AKsqV/5lHPeWBoAZSskZ
FqBD8llsjvq52DZ72WhfMprO38yEZjesQgEw2VKcNg5iNYK79Ky3qW6oPRUq
9Qyw6IqAqP9FuAbBXNsjnx13oyJd9MYqFGV761/mpbBLsZ61BY+RlMoA5Cg/
Am4EeKp+RHdd0C+jbtVlhhndchv5VuN6Nr2HnEjR2O+XdaOabc8+nUh2zTVo
4SXw4HHgqGmzQQe8XXY2kjcA6Jity/bjlJcii/qnuTw62QuDqNlEsG5ZWm5I
LyYoBz22prHV7dE1IasB0OOzI5NircgWwyE8BDNICMZA0EWiQU+lXd0IMihp
SGXkSDf7X4DU4VmY5YQL7iWtHFxqbW3Vjm9edYtCNwoFxpvI7x1+uo3YDAm0
Vso8LGsQ1FUZXLCLvvNXnJA/iUnNDZpmJkVFaTikQ5lIvA8DiZMHq2w+K300
PwXJF8h+JL0Ng+/qMDlptC32hCn8IAB6074Sp3/jZqqCjFtRd80wwFtbXOeh
tCBXu2kqOHEys+X6VJVOFKgqePb5h8O7Jr4rJZYfIoy+cThU6MbXJuQrWOSc
Wp/GX7MDXt5CwZj+XzsA1eTAn7AHWBATKuMYXc83AHee1ju9MVFpt/AVckyA
uc2sGMr22rY4FXBkhUYO4trEvUKq/CF3+roIXGSo/CH7O/rqfG8M1scI5XeO
sFwyDLBENvz88+TKAakzsJ7oTMIx7LUu1w61GXbiES960bbf0Av5Tj++HBGX
7zpwipQbneX6trsLG83SVGrd8MZCMbH5SWvxXRV9np4J81r43tIBh8KA5FQM
5TH8uomwo3llR0gX1D+JJZLCSUsL9DQW2/kkmOPbebo3gAXtir7jijLOPf1c
XZOD7ZWHwP4e3Yb0PVKUPXRE9BVZJDjRRGcdJzuK+lnx3voZ64q6CARQjUz+
N4Ug7+4f0T806Pc4ivWrtSgJ6+Y2DpxnywHyA+yCou6tIbL5KYv/GOYyIGQc
AF6ttjSPPaQjRsUVU6+9jf3hJ6sOludiOBxrMf+FzZpw+9QG2IZeE0s62El4
6Wr9+FddhhqJIQyjdi7s4+hoxxjWbAo0l5jgSxDfeqxyR/q7G2GMPdLqPWUJ
s7RPHjZ5EXvb+yxB6GS1Xo0yEbAN429fBbXM3pbbKP4PQj75Yb/2t7R8Yeko
aR7HA5/sqscNg4X2QTEa56whd0frJ9AqHsLBt9y8gbiJWnmPrWIdv7SdCZRb
XoLLpgB8LlXLeYh5lRdwZJ1BbI4W/TquQRfHNrSDQC+bCKlQYeTZ9m6VzzcI
LE7CN9zsvgSgrx4+TzyXCoG+lvvtTOrjV39+0aFJpcn8G4+ZEg4liw2/sMGV
tmJAuC7W969qn29vp0578fdkLKohI4bL5MtQrXmHpE8pMUm/5fJftMbkn2yP
VvTU0zGitfUq1ImsDbbqnCNAjeZl6tmuDj81H7f4MAX+g4U6eEoQg64Myfk6
r6Nmhdeg/R29muOncl4uzf9FjNeF8WnAgIALmq0Th8el3vez9Nh9nOY4uEcL
DCGvtyAziVFA3d4s/FXfcPjgP3NzUpEOSP2ym0/OdcEisUik26BiZtBNM7Uf
3vno0ntT397z7+dAvalWc70PqjIHKM52riVn8GjpEfRanDtldJzVIEC10eC4
zwVG4yeHv0tuzQb5+cGALUeUI1NrrD4EHNvuzXuMJ/FDi6qNlO7Rbi2L5eNb
PQnfZ5faRKv+K5A4t4B+GzO9kk/yiSkuLCSpLZgjqTj96wt+m7trdXCuznjJ
PfWyp2QfKZeJ7L48Ec/IHd86OL5DKkdN4iWSll8wLrpxpUs1PBWlluDhKUen
4mh4sEb3Tv5TaayZsBE93qzpn3iTLf0Yzgp6unxy//Yt11TRfnFV6DMaPPem
SjfWMRHjqUa06BR3nDoZYlbjF/JvXzi8bOlZnUyMivUN9ktZ0/+qyNgP61Jx
3yv23wrxgVajeITnvEyIGy/9jaRf58iPNPTHcIxMIvuSvfQFf6PN1/s+L5W3
Dpm8tO16NYzKjgn3UgKDD8psJM6hs40DbWrynRY8galLOU/QWfixVHOteFKP
fMCbSTSTJwxJnWPimfTwvEL+8q2irt5PuUY3Ij5SrNRRrebTHmnElP2CIYgQ
bT2pmF6OFXysTCu5mPUEEQh769rHtcgzDLBgZrT5B7B/DmCh4c1DZZbYu6Zx
FBuyszVRqk2ncacBD4dUPJtpizLDZHf9gcWCNw1HZRqTHPq9AXFwkg0OIKb5
fnLum9OkC26GiEOvli3ZGlAsjmYwaZEYuwJMT7Xs7+yCUCZCO7la793gNK8U
Or02HVDHvspPRuAy0Js1+Iu2JcvlxNP3njXYYkd8TpthzVij5sj2tNlLSmgN
L9t7fiC1s8njq/oKtportWpacmAF+dNgvgXj8plfkevRbHfkckl/mJI8oQVJ
B8Iu3oPWWu7TBSv8q3hxrS8dmVWDWdhs2/NBGG0/dGLZN6P2ynYxDXbUh1Rm
Zh/NWt4AMygh+otqIgq1zht8JRi8YNTVoRleHOGNYzap76oSbO3TqpudaetI
zh+zqSiBR5hGumwRiK2JbSQoeLcFXddjdpB+Am+UAJEu6USAVnrHgXi8NxJ/
cJGor5XtWD0S0547HvqVRJdzG2dsm7F0GxtPttlclv4rSwtJCPAiI1JUtfNL
YYmxg+GBQDEpWJdZWQZzVOFmBVRTKZjQSFKm2PqYHoJewv2fO9dQ4iA+jsGV
rvMmjqbl9U/udL46TMESce889FWad696dAUZwcs58PZ/FuWcLgnRVO2UB9Vd
dCEH9nyEeuGS9LVuDISXoSRopH1d7gQE1QJOMfOZJr/I5utxrHocBCOsDF4g
2Z3U76qrwbQbFwNihIm411h1A5uD6BvywK9PCD46g9QFZ2yDa5hSXrjkOvtA
dzDR1EcmDcSxJViRfhZtaIaSr+/qGQ6TPowdOE1qvLHeW4mg/W0pCCalIJ3I
dUV8PRo6RSpZ1QxqvC99Li5TUjzAbaRc3CeJU0UP1bG0XuCoAeuXM4jU6HDm
An8d0TVGDSXYznJgyOjK+TwEVQAnp26Jvl3Au2NGzBT/+ZuTUjCiqJ/3rE2h
cpLuVOAOITzT7bhLQJ0qieA6WpWKM661Qj9ZnjXZgbMOTvsxRZubwpZjpt9m
qs7uMyNhs+n6IjBlepTQO1Y6IPxAaRTo9V91bfsyfjdXAUCju8UXE8t3Yd4b
pJCSM7EZG+myR5sX8UnoxVz3lWlwNFLgsq84a4XI19q28iKUuAUI5zYElK05
eKyTECjmCR8Ovq/TOTmC/6cf9Ksf5u3mQ3ZutpUMIQM4fJim3279AkNAo32s
DkMYOaCUYzvxAVs0cxhXcQb44KPYRmoWZ68yTg5v/jF6m4IrF7LA7UwQyZil
NwaN49AGGfgnjO9n5lap6IcA3eU4T7vd52Maz1bs43K1WEwyyVk4GJYrFM3T
uVjjLVpfI37q3HJxRmtCtoMnsebcwLDz7RNdLgOLaW7z8B6skVQ8cwTQg3om
y8rV6YHtFbmcyXby0U2Bv6PEXWHVK4LWL8jdZ/PxDDrx6KqKt9nFEwiRwXj7
/Md+x5sqfyHzMLD6sC2V3taaDBi9Ktkfr5ggYgdvF5L3hR57yGRhfvlT41+k
tYxX3hKv0hv0kPnqB653ORaSswTPiRRP4eOzOsr/xkQGtDd5aI0RujWRP5BK
i4xVx27q62/pC8JWReKMgvJmtZLbPi2lJgaalodPpomEtSRcyyo0tC8KcHQ3
hUaoBpuvPUxs+s8AWUkYvC2uTtRXB1lP2wrB5c1Id3lT1av/6xMy8y2slzbG
zj716QwicMXoEJBH4a4LEo8O9sFufEktvPoEsinhOFSxyIj/l/4fDfTq0ax7
mV/rvJ4Vj91C04hx10z1OmKjZZrlwSVsM6S8RKtsG5+p+rRXD2IvVU3Pdyiv
P2TnBEGpwnRf7J5A4V+7lpE5vqvQjcbXOw8ub9vE9J8dNZ+tAKZXr9DO1Dmj
kRtDxjqqP/4dXKRpCAlu5IfBTTXK6gi49/cZ3LV6h0DgcnuHb1otOI+5hR5D
yfEV7Vne29Aj5NFsN6Q5jrXPJOwLzN/rYMMUzzzuvq4Et5Rd5eVo/Xt0Lck5
HQVJDplCB4eLLlsTR/5h7XqMEibbeZcWo3BwfhqA39XW72W/TEw7F7yEKD3t
5nC8Dshf+XkkMRkDDEIr+BeMleRyiuilWGSyehX3Hqu/VrsISQ0zyTz8yaUS
e/Up3zQye+q/qChUuuk+yd6alps0+Zv0oscfsckrdL15sWQWEF5Fre0awvS2
XMWVN7fdi1Q0hhjsTkVzes7JVNGmsgWVOCpTnYdpQpKQJwlDvMYfTVJz9Gm5
IPHMpB86x4Q+Y7CgznGeKmB9VnZ/pJnoHy7JH7TTISo13XcJUFZgyaS4h9Fr
ZgGBZqX/J3irX1RkGYDt94MoPIrjiYddNbnvFWxBPwGjB8rR1177a7HITTFf
paRgLzqYVoEYFU50GtvoaCQbGYdNb1thLIclf2kKSwV+xVs739r6CPhWPhUW
8UNNxLzGeWwgFE7salY0g0qtlzCw1Ojp77GdVcM1J5OlsYXRPzSNz+PXEHd5
2G1hs49bWPH8/4tbPNsHuDVLFMdCOdIONcoI4ESZ55K4DcpDzAwyrUYhlSCd
1zYrKOJ+FK0OChLww3XfnNtULr/ur9bcNozxucLZ14w+/na+JIT1+VO5uPMS
olIybFP6nOO/IeJ5X7lf5UfUR+r6pwBGFFuH2Bz1NrwjvbULkDsLNiVtrNRN
OCMDxEPntzPQzaoJ9b08szuAZFTWIXO0G0z0Hj9p1ryQavkYHBBtXzNArB0r
xKTgeeGN9XfYigN3USEoEoHd60+RUamrOlrexJ8+No0HLaLuRALC0ofVKY54
7qr27ks74kCMHhD6UU/yOwr76eUqEmNg6c5vESgpnMJjfX/vJEg/MSZfZ7G+
G7ltCs/yrIM1YZIKZHI/1aAWO+fp23VmJ2DIqry9JAUkqEYK0UTEsMtY4tB9
LYP4tg4Ts3zE89PycGOIjW0KU/TmKu6Wd0fbV1CRm+9l6jeLWdUgsK7+s45K
teupP66Cr6ZvFKjEC2WGJHHf9dNuoeTtyHd3BUKg7zbb7u4SQadhi3uW4fYI
J7u+BPZbecyREF9arIamPCYRI7DzvfYv+WUrJguQ/C24jsKaQdpVsDRkG2JH
1D2GFbkQmmfSNkZZnxP7CcjGqoixfHqcWxJRn3wC/kkNBcLHmtf90Klt8nSf
kPIhGmiTyYGrPUOgvEg+zI656SHCbdADoTBcMi62DB2YYcOdeePfCX2qlxlV
Vtgul+W9ZZBPs3vMF2kMkAKwlQkZp1jFxnwY91dCtttRv71OEU7bQH/jCR/C
hgnbRFVU7AnT5IKZOQ2SGdtGfBnT18chITMjlkZ/GxCx3sWk5M5Wbt4AqOK6
4PhSCl2G+XxEE6XrbGS0A3Ze2w61wS3ePjsPyHFcuwmwVriMgAtmZmIxNHFZ
5ViS3Q0o9w/BZTvH0K3V9LegNBBOq675DWcB7SnTe5OLofMYBoAk4b/Ht/4z
IFFUmHCx+Fuo198TK8olXpG+i3BL7rCFeqbByLHw9TNRHUYyQGMK1N8DzFKE
RmssmA8aVYH3+o5sFsevz/lPiyci/76Ov3Y8Ezx4PwT0qhpXUwR9ZnP4C0u+
j8kXxqYXKdPBdLosmBF6yPCUoD41ibp6Y43NSGjQ04Hzd6tXfARGWcIFZ5sR
Gm0BblhdzEZMbVXBT+iWUo9gN0HfylXdfNgRCo9lL8Z/pEVrWKqjmLVqFA69
YO5bfDtFRyhqFXyzQ87jhZseJje8U1QVxbNT4rLqBwuJfWvNJMiH7wKvE7TB
hG42nUeEmg2eDcuKI2VWahudQ6/ETC6jheDofxx5IYxcYImaT5JXvs/8DAo/
NPY6w6Y7SmaFc4D785VO6GBY2kC8/uc60ECi24CfKdbAOc1E7AeNUcTepAho
JuKvEDEWYU00+AZSo69fZAX/y4kjwA9/OsmjaZqzRhVOuIvppodpE30qNigM
+6ZT14WMWV3BP5+LIN37axyOEKfp3TN680dQCOG6balxz4LROVoMN3KtGQhh
4gw0LARJb7IaPYhTvXhql36FBysuc8dsqpZtK6uYPUKF/m4jAXPR+Zsi+01d
hvyXBcWLQqUcmXJL7K5shbbtYrJjb1vauyychsV4v5X/EIO1SBhfuRmkO0sR
1w0bQiXxp6CmcT2yn8MCu18OHiZ/B3cT1A+5ocX0gYdrwrVjdFCq3CsUuTKC
6CL2vNbJWcbcZVQAJ5UoGSqq5zmzyYiGlalnARDFtBfyxRV6WnlsmYpzZRev
b8rBF3c8nFLPDcshjSoaLWc4+vHz0eznjr6HUzfmdN6HoJyslPByeVsA8nMn
tfM8fgpH8KDTP72AHcZf8x+eX2Yos24hPFHePjGgEUrG9HMUXn9byUUkXlsX
w4dzHPeYKvj/fyFmda1J8Ti/r5+jzGT6KNm1GctQn3p1fFoyLrx3887eD2vy
bjO+ex9RYaSgJD81pO94cBPxz21Ik0CIaGEzuWe5PxaF03+7+sB5+hhH8w6J
/WL/0srzR99bk6hqgwbky0Z36IzKgbS/hs1w00JkX3nmPOOi9YhD6wVvF3xA
vQ5a5PfGTa5764EAMHwk+oCXc7N4q6/S6qA+/vH4XaJeBkck24VKkI1F+N5L
fRufNwV6d2qQ80ahxkt1skhH1jhy4lWNnqHIMenEfva5I9bOVEs7kqnyHteM
Vgf/EQhowHm/S6KEeW61XjGYnktN3jvT/sUqjFyFtewGdC84ndmnca3W2VZr
ros+HqwrsgWiRhkj7ejbvhb6R+L6BBqqo0RjpNuIh146WT9RydbGGqX8AGrl
3NTGOYxWXB7UGN2Of5tXNHvNrJEoJAGiarq7Sv7/firmKmfntVjobBJuwGTL
Ndx0uczj9Ms+hMfsYCZSrozABH3B/acs3ZzLTvw5ThJHaVIoa+l5UNWHuWLQ
vahAMaCNjk5KNQ3YEfvausvrruQ5x8Ix7tivc1Sov7QSwqRzq9wOvGjPjkVM
fxWB7RO9M4di+l7ZAAsZAXDVkwV7qIPQpcMdgYhprmydglnoWUAdQiYmixJM
JKDAGp3rhK6SABXqU6ROwk4NNISaibRJI5nB+ZO3agvf4TV991j1UUeG+RYe
frT50j60Hiapycdbutlqixe6dh8MbRTdpruW78HgJzEF16a7JZ8nAB9tRJ7+
GfDWTrIrODXuXIbpIxU+EqV7k/GJdx3roQt8O+ATQbEBmU95PLNAvPjohAPa
hy40N1UVkUGnL5EuroGJK1lz9qFWPoG6w6tMvyHLz3bGuPzsIQ8JgK6MVvfX
UlTd9FjsJns7+2ICsXYHr921fscIYezekS4h+p9/e0ofeKCpbpuTuj7l5ZjH
qO74npPs+h4xT7HU34ejv2Hxqr/mdnhgBeCOM/JCThfAoYV3iwJ1ZhxZfqN+
SneZ+dJBMvL5IhkunVlIY+os2NzrLSxIwzrmoHxqRLcuJAEQ0Q6o6aoLm7/C
SGORdzlrQMs0kBrEqcd2k7xBn7I550ppbh71OVbCF1mKFJNvpVRNGbl3ebCE
EekZBOnP/VTZF+94V93aXQPN+HF5IsieZJtb3p5DABEl7yjFq8BXBiiVtq/z
pVzY619KiE9dQFcAJ6dLEi3MlJseLBdvrK1tXosIVIaNYgQM3e27a3eeeCQJ
B7hl6BFoo1FlIQShIHortx0uOtrVk8qklKMXnW7IVE9qlicQqhJk8V2/UUn5
9pgHQY41m4UPiXLlweF46iSoDwxikelH40Uy4pgbC0XJl5oeWhboIdK/4VfA
NX6RH57RAKnkHLV5it2UOL2f1p06NOeYh0uLJKg+J/SHksFL5Qox86dD/Glr
slgTOL89XgWgVJ99zo5PFTTJ3i9kq1Yop9hoauHK4Cx4gryGPbQZXaMdZNHq
3eJSbps5mkA5Xiog2MitIRv/hE6hJUoF9IOvH/Bt68hUXFrefUgs3rUzGNFy
LdIfrKt8sWG8Obd4Q9EdD6pXaz1+35mzPbG9GN0MpTLwJCYu5LatLdkV1nqp
3z+rXtj0JrHeY2upNH/xzk+A/PUbDt4iRVrXceV0Z8jW+yxYJL0du19zBU3w
CRkOeB5Ztfn2m56TalhsI5KQ5P/bspHaTAMDtlSrIktob3HtXbUgLhyU75nj
raccbYLrNQ3oXaJ2uLjmh5+V/Ce4Lwi6MOIZPka/Ci5BT8TMpjYqa+Em2wGR
lMMAtYLYLrivczStq15U6St1I/mNTgXOPO0GeTuTpwMBtesgpuaThiY/ONvD
SxjyLFuAWj6C7WpDI+iwQQVq1JUbvMXdB3+j3vwM7CNVuAkM3x4wFsX8Nkrm
UYfPUKIlnPEuQglEuz9Z/ZB4KXr+GtaSI8hR1/XLINL/x47aeuLwgAFzwZQz
tynniZ9ZWHzMcOLwne7/NYl7w6veJmeB+bU5mkslm4C5Z3yuaW4oX42T5JjY
sKpBExD+MvbALf/SlvW8qgg3B94lt+8oFdCTJXO3VzF27Qz/ynNlAAk5IvIE
+YHpfZ30Oqs4+a8iy4pd0HWOVqkd1ASXguJPnIVeWYzmwDqGb31R3/2zuASj
NMLGuFWQTfuKhypOz218ZxFgiKDCN0QaSud/RSjcJyDW6ZdGkVRz30sXj4i0
gCKV6QgW/IIWlSe5ajjc8Ou86wVa1huARlfjc6LljziYAbVJFP7iv/k/wstf
CXULYZ+ZXFoX/JFQHdRQ6bgqmoD0oqfB9Aqn4dPLqWkUgFRlys3KhAQfycKl
GasXHAcPtR5nTo5TMnuvgTCqnxEvkAxYZC7r6pxJLOsZNYdDKediazzruvxS
5PQ+Cks3QH43YwWU7NUVusnIg0Ls3UmalxzSVnulnj2LADtKH+E1OM5HFgVz
k3zvHHzFjXbMphi5b+ipqz+w9hmw+li7FNxtDisuTGvg/GBVC2obXuwHMj4L
IQFQLyqllk5dzhNSXGej7Yt+L7W/XeHjd522lF82N2sl8B7toy/rBGAz1VhW
qlW34fXe31whE0aIEXvXtj3ZyTKFcXJp1hR2MSNdIDj1LNWCLL0pWakmKAY5
S4IxAmWDNfeSsMRVrj7s2P+MAv7nnsSC8pZBGXNDfY74n8pjKsKOnzAimJM2
v6c/CKRQJk3HfkPI6kg162Gu5GLK5G0Os2utknsU/dMB8RLolqVkyNK6Ls5N
HoUdEbOfcAjdpRSpy31z0JIPS6hb9BoQUXOROOsJQIj80RZ0srM+spVZHtnt
eNJ3Jj02ufnzU5za0eB6voyu9aTyHW8yUVpLrL0urWv4JJUIOS4TLNLPj+tO
+jNNHWXHTxiCMv/G2PutmqQzyb7tVGBXW10shNL17u6P20omajqHRMvr/vMV
4yOIlsOdiAepnBpDAsC5TzKsc161fzSQR5OITZ+8N9+6knmSK3qejB9H62Mz
FmCIuWErJdqupPW9bKwSWxGqaXcA3xKYQW7EaEUCVcDrFa2NBG0KEoqESp80
XgIShdQRvHSzc09GCsvHWJHWkSgG14vciv3MaBrVvXS7x/14SpwTBAVoGApy
eixLxZVk++QEB66QGwNvwjL65GNvmvqSwx5oGW9KqYMuCvOL2Ml1YkAWE2mA
v7YzHAeeBQO6bs6yHSMY+pNQihMNKMZF5/JnpezD2m9sd6QUk1n0xEcH/hRx
g7r9Hlg7Ap+SL/X+d/mq6OE4QlMg3VbUu+EnOYqkDkGxELv1rO25igQSTrhY
26rl/1ZMQmBIbvw57bUiBt4wzszROtd+1xFyKdtvu8PUXEi2NUTYRYh3PIV8
FgrRX3mbNzD9M+j3/w1lO+AqUMEAPnwPn9WyY3tGAyaLLv+uWYUzKIo2yc/8
GIgF7SU0hfeyclwFrXcspnb9zx6ehVXYzCMxsv0eTCmv+ho4vdlO3Xk2qDL/
tI7w0kw0uG4QTqaP6DIAru/3eGwA/S9xxH9LRZxnPpZJZ8PK31MDWbbxz+7R
v8xZodh47yKlTU600zj6n55JhNK5wMPu/JIblv7S4DLk9EQxGrSGV82/9X2T
GaWSEJlt9g0jabY0etC+HgxO3w4hRjPeSGtpm+W90VrQLC7Js9fKVshmpzEz
7RZPf9K9VQl2wQAdTaEqN8Nx5zUNEQUghXzmQFS51wQLmY0Jw5Aykd+eQikR
OpvM8XeHsLyViAyVdOP86RMlxXq9FRrOjAbvtBqg+gi3OTm4kxanhbUbOrYS
H19Hp03N+hbhRuNDmhdta/RZd2kN2b4ge3f+ombOS6elP/TJHK1T2gJSFV5M
8raCf4Ay74wO6bUEXQE9EiUAmnObMIQgYTpus11iGpQVc+RQMjqyUoWDBn2S
YSyjipjiqzBXfaD398FC6abc/RFfrwx9nxnoJstC9uya2MfhGrkV6upF8oTB
4BuWHJlsc3f4QeCRU/pyCW0z4z6KAYdFg0/F7z5BGWYJHi7LEh2GDo4WRBUk
lX1tUcIRqlxpSg6/OLyGmlAIsnKkWAN7twsEncA/YiNImqk/C56ObJvgz4KZ
+90DP4phDMcN5vBZPEVvPe96gOVjWYZMJBQtdvqorCdfUnzDhQPZvRc5FOLU
Ha2H4dOTGBUOKnKZUJW7DBn9dxaGOwbk4iW9ncyTM7ZJ2KohsP+YkT47bxqw
/9KgVpq3lOGMJM7ywQwIXbAZO/sJVd/2FpMcz+ykQrnDjEX1p2AZnWLO5lxl
/owLJvc1FmEUdP8lsk2ZK504K0h57Pdkx5DZAzxpSduAlj7J/HzttYinJMTo
R922ZKl+IEL93S55Sn1C0ZwBt4NVFoxpk/+LeUQT21JB8V5D6Ledmu2rkjpG
9Cwho+CiPxUYk/AqFliUH/TD71X4eq4b355+oXYUHKnYd9GEAwntOCaHGb8A
ETUMKmHqJY8tt32CBXqxyUAQO3nV6MfhZ1PkT50rludmWbsh8L2FQi+WXZOW
TOWHzWRFwK3Y+ncrSS4Okr/JWiXriU2Y1WgNoBUk+wEFRGaNB7uKyAZGEvKk
q4rOgBQA/77PVkhKVSoF3ZUOEfostEllS9IjLBw8m6ix+3f2R93IcQqUbDbF
m98J0CVKt0MzesqSpM9OxaeZ5KWeEp2+7rwCDYhyaHmZ+DT3nRcRk8AJI1k+
kI5aGFOWjzqyuAauJfb23KOj6qh8lOK6Nm2yqC5xjeJcfIbKROduKQwgORtO
fF0+P8hWCv+/8y/mFODHVJukU+eAt0B7QT2IIAjSRjgAifNV7EvqIBa2WaJ2
13eqdm6eiIq8iL/U7z+U9O0tifjg2PZHX7g219bk5LlHWWAN6MO7AwjVf4xE
RlEr0Nk/NjU6NeshyJqqPuI63hVDuS44/0ZFNFJ9imQ8eCkU0hcEWgUsESKE
AdD/A/ggc9gTm9DBmu5NKs3h3Jr4O1RdPZozTnM4aSKaT9Imfat4rs6HDLIl
tCTyLOPwVSetSjM8fg3UDUMQVinVkDbDg/6n+Qu+ldty7PfD6h8eJWcOLoLU
D6d5o42Q74lOLAch3ALIZT0hcJG03koJQHdrpyKwKYB0XvzF5poT/z508GyY
09mAbzfBpgJv+7MnXa5yCiTgNNkxwnwWo+f+24+uepmYxY7X63KJTAD88I2b
ShRtJvF2+rGWFuqDx+AxEexn/fZLHXYugOL7c/57w88mgppjrokt7EAaKJeL
I1e5akQvnhQza0sP8nBqc5YiRGyuMORJIQlqu7LAUmn/4wZHhVaYeuEWD6jf
syj/3cOEgM0APMjZuneV1KIgzZUZD9hGFz8LGlWBuEBWagYfxHdCN2WNI/7L
iiElVpzM565/s8hsjAzpq9T6XukJGahfMstBc67RyIIVwuB5ft8B5txi6G5w
F3ZKpnTrAJatMdIsIISJ7Lkp8QIkWthD6ByGfr4pthHfVxc/CNmcnFiORO8a
LoxVOa1onS+NRVu4QZN2c38uMczo0ZC/uYTo2E7HnRSmIrGKteXFOdQCxrXl
e3pKee6OVz3n9YBLRV/lySIWXOnQCt4hHEWp3/hHTC//mAzOn2Bq2GFRY71o
gqtmsmlvdEKeABIzHmSwxsi4gUzIUl9NDxcjyIzGZnfAwVHmzeyNfty7BVZR
8ekwAhLR8iVvAuObPBz5ElX0aj06QeMuRWIbUUqCmCDiDv4YbAyi6Gi6RNJa
NIO56FmkpOlHIhBzAqsAaTkLRTPvSoB4Uk+F1TCRmdlEZcZufswewk/hkWAb
3zIz++hlyIB3V3O/fbLdX+hlqftq3qAcsr5jUd5j6F6EH99vs77xA4/F8eOR
8/5aHW59jBsq1cvebQFaHP0muLwgDZoCZtHj/XhUqLWhGh1UYUim5rEEFOXI
AFg65sYaFP0Qg4N/4tLOZvM6PJ6mqduGVp8B+JjSJkTQehArgDrDMlxaI/2o
0DwV450DDotYAMWE24fzvu1QE1pRqrxZsh9+xXak9XnfB9CVGvpw999BlcD5
74KmAO0BN3yExXXUosHFV7JZaEkC+Sfxi4q5aodAgsHQSGYjf3BSuk+ZEzkp
ixWNgGSLe908/oEICQFjf7D4qXTDXPEK4MRa+Ag7+2wUsJKJ4/IqtH7eo/8N
f9dEFmLeXVtLQGMfV1cBUnoXbm6dO61ehR1AukWCpb1lrnxuqLr6/cFHtGMq
yOcEVsAhZgabXgEBEw7KzxpHBL7UEM/yZpnJvUwpJ93j31OUqW1fV6jcVYmX
+7iyq1a1whye0sEptjCkA1/m0mqcLJPG1wY9AKuOTyPJOKf/Gzy/ZjXux30i
lz8PjZzGXatEtlMGv/uTAugozeJ1OwlspS56mFCjn1m5lLnzJZSY8xoqnQ7W
TAwTgo8eTayG2DvoeLGZolPQwrf7vbRXHnUsdEfK9as3HVF/Thvsz71fjrdc
jt5EMeWUnkyc/fi81HrARbUxm2Z4fNMvRkT7QwpzJoUfaK1IKpBi7edlbPTO
qmWC0lFDOKHXDfwmF7p9mthCUnPYimEiIS7U+D0mrWq7HMQpWwCQCC9qOAJ3
Zvf3pPmFYqI3vgRdzKTlduPQvq+BmuER6uFJeZImCJj4NZ8EJMlW8YngphLq
Aa15lq0H/aFHVKTCeNurQaTOaQwF/kLsg9ZNA1v7qhRQVlFgQYFPNNiwlcu5
8Njw9VczDdcNzvnwBTxbXohrjp32Ud9mT4JoqRQVnC2y6yekDBXWpfn5O/Es
mQHjAHz0UdyKcCAWd8OEKESzEl1EoB7VQncxMaw7yilVJb1qyZGtKgfMhKuX
VzRjkB1dY8si/Gf9I2xl/zIAhl6tl+WH4NLLOsRjB9qEwLt3E8ywg7WpYOmv
GVzaxhUcdox0JpWjhUJfWW1TJHZuSqCR3NdbaIFa5mJSNVVdBC6nrXAEp2R/
9bJQNoESYLfZu9zYcnCZ/0ws704yHcVPNLVXPILzzteiX2n7PR2GwoDinAr9
wdgw/2uFmx52CRO6Z5iJNy0Ffzre/L9zX2EUnF5ZE6+ZGWIqKtJ4M3GE7yCo
cKGyzN3eIz096Ea1Fs5GWQnOUV4X/SvKbVn+Y/9S0boDU3c1MuKekDanEnxK
OTv1onz/ZJox8RNN7iP5ceoMjb6aq5lxt8mRHDQMsSHBAdfTbfZeToALJNW+
UEHcNctSpAmjhxotwghVVpH9yBOI1uT7iTFMK0QHtlvW/ts2dA8wO7JWru1n
v0HYrua3tw7i4eT4hIRvR+4+X6S87GpeQfKqZlkfCKBgSUY/abhFWc14DoV2
zuNMSjqHhsjim6hWI2b1+ZXWD7etxGPsFunKqUEa4/8muWr7ugNUFTsSLpLm
Y4KFdbaRWXMMxZNTTwRh+zg5QZwGpRhgLclS79hZnDmInvc2OBG2Ly0U/eJ4
8M9mixGYE2cLWAV02JZ21daUUWxDZD3Q04vqPQzecGg9qCC9tFIip4mgeIu9
Cd+sOZN+LTNsEutN6SG/An7UVEdPANlqwfeyoOQjK4yWYjKnwFpxVZJSfl6L
6BJ8pqA4+5fHp3tuJ7ZwgxNQ82mLommeAC4TWftijlX3AZyf7M3wdRDqE4qY
PQjEqv8361WXl7xcooRlf6tX6PfXkXcjmE511Ps3yDI2B3O+BXqpOFQGhyME
boTZ3Nb1E1HmUEimAXROBZH90JN+Zb6YZ8wDjloHjtTtBD2fEcbfAj2XqLrR
UXBJirlQ8G3PCYmNIEy7p/OIOFlgSGtP6G7z5Pf58lXJ/qJJORlJrmFZoge5
yaht6cHdMK0OABel03pGf8Bcp+ARIqCnkLoanSRLnHhwVYkVruPOFb6XDght
TkhpwxnS5p9dEhvH51Go0wYKk2sJ6Z40uBh3PrVNqz/oZ1i3KiIIobnfEawl
n9TT5lK5Stj+RcdGgxk30c+BoYx6Z4s2A4GrdeCFriijxMepvD2zMKuS5Iez
mxf5eDWVFfL7vEJvDwncRfNB7Y19oihPy2C86iJkgX57rj2z1BHVUzWv0Sc2
BGjv8qRjzng7juR5tSuhxSgeZYq7eM0nDJr1I97+z5x86Cbgk2QOijs5Yj4B
QVbAa27RAB4pbMP5I13XitOmV01vwvAgjzRirhXlFJBanWUi8RtjHbDO3+Qf
Bm8tKZVinmZXUIvIh6hcnVwbVv6UERUH6LTn9v7IrIS/pErSfdgSqdNRlP/n
x+ulQAQwYVSZf8X9WZpb+2LoHYCYuaqOHCIg99VHqfYYAT5awayl+mz/bjLJ
hgNyCNlpgNwtagKJ0zeZHfUqECjvZNKi5XuN9K4ECcZoUTaVNvGWBggiUYoI
np+pQVoSq+eo6J/+g8IIfwVEN1ZSDffmLxr8yCUWhYiaWvESVcdnpDAZm7l0
b89PcpcSngyA70UF5IaaJ78OeVy7tFBCLC7V1vypupxT7BclNtOSO1XkPq2+
yw/woGBRml4F7EgLSI90vqcRfIT/jj18excnuu95eqdiPF35LcVY4bKs2UId
xZ1+PTIgGjDqcrHjpvANJSprWrCJDXzghkmA7LqRsm6vkIHBJi6C/s+2YuWq
YI9IsyYwO8r4VA5CUuqfohsFfJSIe5l40CsGKTNdi0TKvnm1trVrCbFkOt7T
h/IcMXTrcfUPKIUNkbFrZjt5z+KNN+fXAuMT85OJ52z7/NJ/Lr83goUIZ//o
RWbaQnH7upNnI5J+SRqo/3FhcMWQucpTUaLdZ0USXS2JWHUB6Uj6TzGDwIdl
+qvubHNlhHtq8OCaPhH+sKGqiTTwTFHSmAEk+pVLD8e0NscdzutSHmtAKc6v
MhN6ivQch5VN7F37l/lWorqVzRghqmoxOSmJScAEcCGEpRQNHW7Mgxf6ljEg
tRjq1ZiFgGnJqrz6SORhVGOxdpk+/59bc6XTRp2i/tH4qQrlnHQU/41gbabz
MsDxZmkfKHXIAl03+GBgihTH9bBsKu1XvNMJat7AnU4ZuuQ0CF9V7l+TtzYu
LHnhs6fD2PVovvVD39maElSLeGnSpg1qFZH7Rf+9f8pZJoSMGlZT/DUy63iY
3nmDS41emBV2rE881bJlNT0CyjLPzDxsdNwyDoXOu9CqIIi9Aq0sWvdOTQ+v
dTAcly6Gu9MOVid8Qg2iwKMvXdPaQIW9uxA+W95exXmWSCdClRiYX6DuL6Ox
CTN3GiS2/n6MxJBzX2wdi9jQEElzK//c9YVTsYCsDR9L5L3czjQiNZbYn9Sh
sLIt3auE3d2QZG3/T7zBxItKbcQEdskHu7vcEdnZuBPoXs7zgGURLCN+fsL0
4H6/PtvNkMHHMzt1Bzqk/e19ZNga9LoSuGNQZCg3rRYWLihzS60mbNaPh2y+
bwwkd3XxtDk/Gzcnl9ooaDKcZ8o+RQOi25+FvitWSSVZyfcGPMVSUcPjg90t
sLIukXNxhJeeIVBW5dalCKDhE0wom0sFZaoO2zb95Uhc3Dle7nDn0r6aWg5S
cLXYLDBZDR8w+e2Z9RdJR3uHoqBPUfGkzk4fBbRBK2UPaGpuYjoC12pIs9vU
TA1ZqZJsqQ2ZD/c97WQFKA/SaOvZGkmDTAlgVfcDZLC0J7sDiXiNHJpRLXeV
PWeoyP4MruZwMANA1colT0qrq/ua2Z4bX8pubcxdby89mBio24U/zXNJmVRt
xZZi2gG9zTWjlJgk5kc8uezxQKPTh0xnECWvQSdRwLftQ87+xfgqvRVfW+S6
I4AabMdEjDgmeGn2jDEYzqx5sovWL/+3IBp8fz5QZLk3UAqIXXMY9qA95uUG
4x7+SSyP+TezpLzVVwciu1Dyx5FOBDR+nfMEPEHQG7pyDPQwiQ1KvTgFvZAx
c2wwu7snF3pjkKx5XLLw9qt48kEqbV7ImsMhRgL91lctYxXgY/zvac73DOHc
rCL1ioTsE+q3bWORylZn+2cQG3mb9Na8rk5OBHSCnfyHX9y0L8X2KR49ibzC
fFmu0gnbCw/AkpMbAbvGIcYTTMnd5gPaHiCf0cto+LXrw/ko/X0cxyLcwzFo
lCfxFTNdtsIu2Qwm/2IosBDZTZqWm3GD/cLARRPAY3z+Fv4CREv7FpteLrLF
Dat0bv5TcPma57Rhtg/OjE/rz6I09TdjcNzoW1eQ1H+HnXHzkInvIbWbcbbN
/Aw9fuN9nPPQ1VLyq8umslzBuj126cQYk/mkmSywkIOK48+ntr4TR1BaFy6G
uf6bnD3ZoWbwv/EzhWog8SzRdTWZqVizoNGHnXd2bpWXkajBLiUcoUfs8gb3
ZOOTpFLBzu+EvSiA6Ci/lHUIypGokpONkqvw8uNjVC1y8fFDJr0K58zuz1v3
LlPF6FD99xn5m+CmPAWn58V4ppCiZg8RTOamvLopOpv0SZOlTZZ1/uog+inS
DAXM6n7Cl8MSUaXp+cWsdOUIC714VYzZOmgj6P4R/gEwgV7BLr+KVDadf2Dc
lzYT6TVYWgVNd9xneiRc40/hXlsD7qsG4hgFud244Q6hd1Pz4YvlOmC3zO5+
3Zw2v3yBhKlz4jzMD54Qupor1ybDl6Yk9lWJppOTO3p2+AB2DWKfzYl5CbCB
KxIs5k5xhhkSCIb6DZ1PrcQYEP+ENzg7Us6SrMPeKx+ZABbDXjdg8kVp0YXz
7mZJ+3b/Ne0wP0hmCajbMJr4CfgJsWbJjm4NGDePmsnlwETOXgrBXdqOZw9z
SeWF1Wiwg+AmWpIXCerYbftkShs7ok4GFqCOPqMbxNoZCEeDAyD3YPLcDQx/
HZy1kghjDQ1+C9XGoRZeDAncbb+CEoUUzP4w0qwum6KKs8z8oim4H+vKO4hB
GnCbkXDWaipoI1NtYQfkjPWYqduYdw+Cvh8bMSw7pEqFtklAEoBAsW4z6KRf
nC1/9UHgFQ8t5OdGuW/5/918pR82T+MPz+dj2H0moV9D43Ne8a6M5vko8oXu
kw3YixJEDtKJj8hWuGpekGtyqFUqsFuivDFCZUzFR7wooC9sW/JcgwYJdzrN
vwgMQkOIvbQGsDvFLLtJAZfdUFe0AMo9FVaB1uRhFcPBemKOScawLvxz1Grx
WiPZIGc9KeVoXumyCuU9W/2SyDGl5gDmf0bCSLR2qN37vHW7sAvkFBq6czT8
czj9isk3pUUI8EMrn5pq+OurdT15vqUJYcNElrNlbMBo1/Qj92tRyGv7J8Rn
9r4njPosbJ4WwxuXviaU1rFaF1Yl7JOhsk9pIFer+4rvKUFS3rDmePAhdaEa
ocEjnh7qSnt7YRDp1m9yxzVowcIaBHLPdb7cVgX+OxWsBDY7wV1dUAWtt25U
t7v0CpS5lPQXS48LX6paGHgpk3k5OZx4NyLvwOWnF5L7/QjgvBPvMcKJ9oUU
T1TFOaZSFE/qASUmqQCh8VXsV9q4BXR9xciwhlfdGU7iXcnacdDcfnugQeeH
Zi+SI8EDvWbTomTltIlWozHz5OwurbLRPOBrQDIvacf3VDHohv+Er9c7zhsP
dIshc9AKSNnQHreIejsbl86xFkEyOqDlBtiZBpTyBmBEWzcJsVpfrDnTFfHj
brOWsIslE80DHEXzcuVyEa6VFIZrarM0g5ZSEHQqQs+of6EVU+VxuJ3TcD8R
wN2bb1z7qm3pMD9tz9sdHNvFJNyH/Nd3pS+zZ5NXmfYyvMlAEWqUatqg427X
/arACEnvCc5nWQzdrlSlLcIo7SYdzAIBKXilXGz5BWbAfK5rkYgigIVkDd7B
EFKtgmASHeQP+n3Ro2FzKfu2L8lN1OrgSa0nYxJxlljgFfwq6X6FlmiN3s2L
xTWAZNjykjDxtYprKqNNnwJhu5pdspEWLByVIWSg2MJ/zfppOG4I41lgcbmD
rsrwe8KXOBjaElEd/I1AUXhNiqI5hmPY+bNDf2kryXrrJfN4SFhFHe2by0ft
fc3hSnGXYTsL6YFhQPKzroHmPBaB/2Hkwib5TCUBKzVAovLArxBMRtDswyog
4Lu3wAt0c29bTt3teVW1gXWR4fdjhCGgPirl7/OcxvwD3orM6z+Le8TR/6Wk
r10vv85A50HIy7bhG+gtk8A4e0vwQJUZ7+DGwGaz1VQYkSHuoIPSmHVJYws0
wJwjVuwxNO30LovAgAIY6ayU5lDnXk/cr1iigcLpV9yvuZpom3IFCZbxq1MY
VIWjyzg3QseMlWV4yRmqBNF/DZrahamFoLjNdAVid8dLx2QqzYp0+7mNy9yv
F1+X0fp1EHgzjn9YrlQmBLJkG/mYSo+wIqjWWZ6Ibm66un/0UNkl77jsVPHC
gNyUC26Mok7e4vIBEhFLJwrcQJ/SdoyPmot+my4McNzNSlgCmdMYCenhTOd0
hJABfDBtbP9xO3S6UWUpe9f2REQi6aAoQNHOkrzgLdcUcmdvYhS/bK9DiF/3
DshTiuM+VBotQvLOW/BFbpI5MthBOa7kTiV4Rmtkfmdre/ZDnXRTKpuJmAMF
at+pHMSM2o6UqVUa2gCnfSFWAW2JpnG82NGWS3FNWh+iWomr3apjoYpMw3+Q
7aAR9lI9L7gmrM23E8pTbnVy6i/uhRSo1yXMPdUbw+dqvLkzex5f5odcjJZO
/NQVRHdOgfb+z1/P//huUFTZQGa9a9fKKVioSN60lg1Mb6wO2wYpxXU5uoeK
t1CsLwDm3yEsHY4D+ycYaJ3yC9Yd/X14f23cpfuyQr06KVztccGzvxCm+1DI
msWa0ofSCI+gzDOFltzZAPCqcm1KEx2dmWuT9y62/s6S5DMF+e0wjz8ieqqz
BrhllgnqNK5Dkc2MrnYt7jGUiKtW/Dr0uHJc/HurYAmu8iLxDuxLlgNwZ8OD
D1ZlbmNcx0OTQmokyuGQM7aAIyjQ/qeJKYWoSW4XEK30s5tb1Mlh7imKW8pY
gvxDAWqVkyStJDGAx3klYcPf4N6VJMJS9iY9g7HQNGopLOtogkxQPim9W3lZ
Ofc+L11aJs6VBTyefjswoXcbPgm0tvX2DB+0S+FnpMlVpq04nfanuZVwMni/
RwNYVd2cfjNgS1PiPdfl6svgGso2C5P7Dtl3h8MjYLJx3tE4tYr+pMJrEIdl
rc1gKtvQr7YsV+Kx8LW8gCFpF6lTwflPGWyP3RI7QdOtCYtZ5csI+XuMNm2X
pH84BK/9wi+lxTTLft3oGG81Uwx/0VNYH1MeouGKcnKkRyf3CB90XRS0JUQY
65P1dckYiXUwLGyOWLPiwG1HNEfN3LMVG6LaHTL+ULTCIyYwWkkOmkiEJvGY
Dn9cbDXW8A7ugM/9Gh0xW9NZ6ScCbgn9jyX8+6DwUdDxlOhLlqHRfAhSnDh2
dFIIbwf72z/lffY9eYTXB0+PBB1v36+gAaRxTM2gszGBaJDlQ5Yd09bsASeb
uF43R/zjQEZUN21QGK3b4PhLaVAcbwzNdtnQGqmJs1W9QvABoGe77/kNDlw0
dhxhBu1q0s9PjxLexQ9r0TP3iZQi6ScmDCmwdcHLeVHcMywtqIPVVJ5e56Cu
VxFlHQG9+PIPpzfbZRQrSiVLe0wX8Lz7x7Fx0ydaUlUWePbUoCYgBgHlOKvj
fRzyxzYzrh0QGt0pGpt+zGuBgJFNQVdrMWoFPgXVDuAp6qox16JgRjbEeCCB
zbbqXvZN57t98LBz3mk2g+6APRhCgK6GJQ5sJMp03MIBFU6juxQWIy2zqe/c
bu2HY24clIaeFjt/DCY4IMStgcfODKAKk8oNKKEf9n5hIs40FjLUD4mvKv7E
mD/iDXt8LDmC3/Eou8nZna0/LrnarcpgtLzEM70V4cZc0mvPxDwoO9hYrJPC
ea+MgVMKrd185pyAd/FvYWBSpXwi9nLUSJNuo2bPMknTShIESG121mvBkGp/
FPX2t+rF2gXXtpBmvwS9bKLpmuFTMc56gFOzVe1cZPfz33CVYITE6Bx9PuLg
dKuY0c8K+4dIwjJ3TRCtKt8cGHJGRKNUOmTYk1tshPe3Zg8iRY+TLaXnOVme
klj0nyeoYCU4HHMEvGFEJM6f6ot1Pg1QcWxCIfgfvP4dBWhLKKe1i6HaJZYR
O2DsjZqb5Eann9JSyoSTSktxw9dQBjZatIqW6VmaSj7U/hupU+pDHSggkTDc
rzy8gP7FhpBI5Gr0xg8fv39xuOr1yQo8n5JaFqiUO+V0PenW87DPoV/JuxwP
wPcuDSA7Qz50z6zsQGENawBuxNT8n81dK0ejEwr8gdqFZkZAV3srlaf4bZIT
Kt1AWRiJu8q79MfJAcGgdirok7YGhidi0hwm9+yHESIxzhBHW7GHD4fbyUWR
7z6+0AhQiIbJT1GlMl4b8yusRE6A5p0eNPxLL/PsoQ6xQ9/JIz+8QHgeOUul
+L8BuvunYDS4qFvGCeHEqdFJ4aSQmNsINsf17I3fsxDoh8w0WJqqaiE/H2Qv
Zyci3BmG7mQ1cCk0wR06mLica43YP/gl09hBw8IKYth0T7rGgz+FaYCWsOl0
kdm9LGyEjhXVsql+IRhRBzkQT5/OOA4VdRSFrLvokjteeGI+49l+kaIFSP8s
vwxRsysnxH5/kYoqZRxxEhTtBShQKBhe9Hq1tlUaRuLppYNTiNQZwJQu9y0W
yD2PxeFX3m9EhbehKWshuHl/wybcxWvUwkKG1EXmtsULk23T5XkfvbNvnJgu
JO73Cnv0+g9lYsBE7ncOEgr1GD5kJrZyr/6P5aaSOO+KmLcWUCuwcEVdCiZ+
hojNcHC0I5XzwZBr2n1EcoI6+P7yBNAPqg2JZZAHrMjTtunHvdEBeMih4ZA/
zE1ZrkMt56bmwmjzD7yzkgkSjtDZhA+NrrnT5Pc/fFoPYw6M9WJ5iYBP/sRF
DX0NUxfKI+pFw714soUQMc3/p22h3IWUA5wADXQf5uXrZpNmmcGrc/Bfhr4U
0bXAfL34kEa8buWp/ABpXViiYi6hPxezghs2knBE/i5MLtDmMxcU89uDdX3e
snbWHfcGi6WVYGPh1GyutpkVdQcKTpR5TmqY3xEg24jMVPmfPbIxr8o+Mm2S
f9QXVxKpnrpsAEXzAnYlSccYqXIinI+4rS+eJtulp8ewiYkRUPypsDwE4N/c
YOYO2Ny1gSJKaX7jefQxpfL8Lng8HfED6aK4nDru2rV6IBUcTWNtC0H8SGqC
5+caCsR8sDbRrnOtlBbqV1ul7Lc1pMsVE/3/Q5TNb5/p2tYFKYdZoyqRr0b3
pTwwpn3BEOFvIpPJLrQ4Crwy4Lkujjze8MVsqPR49eKogcqLzhAA7NgIwEap
EJlWZnFU6qNWXI9KVx6MmNXCe8DlT4L4M4OHgoMLfNYs0EzgUAwi22bapAwZ
98tW3yQYH7kKpGi5BtLT8h1iktrAFGS7rJX7kkEzZUyRGD3SK6i0KsR1TNQ5
h2TH4faKRjTkbRaeF/Sp4FO9RKErHzDuOY9utN1zmp358a3gNer2o6sYzIXi
gZpbFtYatFjI1XyeZFhIVfJlWkf3Ff4jBQtcwT+Fl1K/ttKMiiTH9Ok6OOLb
tBFOPCQ6uvkjhbhfzkxIKY8xNu7RUs681zBrS0qiM8SbBylClYXMNebT4FVN
P1Z0EDz+pg0ZDKILjgy5Rv3dsH5uirORy0DIDasNvFCx5YkRyhqU8uyv+mYa
7CXUGg3pDvcFgZR6QIhLBJNNOYN5Q5nEs1U8aCQNUOE2Mt0VMFovwwA29QBn
2iGo0MQ+iiI7eJbC9tEhsyuOemAco0MNi+c/l9Y8fBH1F54LbQAg35XKT8ZC
Ju5E8xDaMBCIRaKU18C8o08P+Fa/a1HpGBstmXEKA+lF/WgFtmgV4+ag1ZMk
pkkjVTku3IS2nks36zogqaz0zTn6z10R9Lttcfx6lTJ+vFvwhxXpUFWJD6j3
Fp4Lk0O13qOd93A4W8CsNpisxih4VX5nIK5Gwf3a7Ak/ql5QZhvtI2RguEuP
ff6NlfwxWWV/WSjrkbIMrH7lxwjHQ8vKWbA4j6Fk8trMSNiGk8+xeGCSI6S7
OJ+cfIiaYVNYZrrOMYccZPz7FXIVzy4RKDiBWn+EzrarRZkkQwi7CdzfLgpm
+jfQWE5M8QcsqbEYBxGRw6oEhZn/RskmeGgbr7Ac164SAKWHtzjVt6fo6hxT
SMyYqAPSolvH2cMwesxIrWauda+WdcKSa11bs1WjhQ11uD6uMdes6eVCFalS
GrZwZJo2ebr48QGK/6iyYj+bIVVCnfjFXWUP8xVtwwBP67Hx4ThB7YOe22QA
garqHPeRbCqGFqgWXGbBAsKc+vsV/r2sTODiCAUBPHGkXc9kFCIXbc3bfGIr
l4bzyTKmKSIPEGL3fd1MTFPJ3UOWu2By+oWyueoJmeKeyGcjeqG4ugU5Xlyc
Q6RmfIHnStRvW09sb2kNxWPvnmsXc8O+SZznUpI+wF/UKk5aDKHXk7bkdCbh
lnoEjj8yt1kVhqKum5jm75vBR5H/FJ284vmnYIoJdTBjQtVxnHRcr+tmM6M4
JbFY3jbZBfpRbwgk40gGqr04sZ5ge/Xo6P4ACjPhrRyRZWAlvoUuJG78NEtx
P9ueHIoJCi9OtkJTYGutnVm+lbiNMaWbBiCrOg+xR7flrggkNMVgMwgav2Dd
dfQUMUW6SlVJpNgnrFyIYKIh+8L2X/rZmAb5GR+l+EiClnvieJJqJSnIe2B/
0Fzu6Mn248aXFYSnMxJn9MryMOTcaWzQzNwldLRTi09hD2VbpfSQU3/g1CDe
4rkH2ba2zN49p2B0JlE+7kgoupWJhGVsfaAAOR24ET5MqC7IDa+AKBWCWMy4
t0vKTPhlB4Jk10LV//KXkSa6VYhN8lY8x1Aw1Dji0rZaA2KmjdTJvwaERf35
u5PFFVnJUNx2cgU04pqFOIPR6UflrlsmCFZMH0NQCff5hu5ekTi4cmfqmMga
6vs58YRE9dCnwMOCuwFgPdn97Oi7gFp2tIMlMP0C+QjDxno03NgTRkH3ss+t
myfEwuTAZwEBJMsMiskfDhOhDguuirLwjh0+X3Hxze2ZNOM3iPU9DT0mRhkP
f2LQMT8DLmJh5HIjIN/I2f/ac16aaO4l5DarA7gXWGtqMTNjdW3zWtLK7Srl
pSr/4Q5xQdl4o/GGbg30ADf1c1DKq3f19yWPiFMqqmAOFaxKtt1J4iUKGtJv
Ewxrff7+FTVBCrvwZxDyBW9SXAIJidwGZfZFsqCbQK4dqulmv8SiQFaLl93h
+xUEViIGT6IG62s6YX8Sf5JMtOFjIVg7EkFDkNdLB/dsST3QbdWKGAvQr82P
ijqyOd+2EuJg5vbtv6oi6jTB6fqAZAAMA7yysfcpb6iJxytlzOlyQaOcCa/S
yscVETH6KReEE6a1KbUyAdOhtwTo/MzBazFWLNoDsVI+swlzZlyVXIfY/Pj9
YN6qyfjS8iHnEd997JUYguwHbup61wfAk65aMNCGH9Unn4IduBOGkQ0zoftA
Ai/jFEtiT/Xi441EKSAMUbn0FNZd4miP8gkSKMhVXpN3GJKNvYiW+9R4GAUZ
HvwowHgjgBY8PyPiXkYuVlj90I19b4PETJDguj4WxBsAwQrSFbuEJZp2aNmI
LI32TNfYgAgMBk707T3UnZqG4umdMotPeu9Fe1/8c06MSuV7BGFcw483J5tN
+pcCwOsaBM7DHPnlLzgmZul26EkRgTlF1xplWENyUxypqh1bRhY63m7YcdA0
ultZ4NlRb1AoICv39lEfp3zVpmwn3jwQ+wtdVk7aKiQ69wfn9m8FOYrR5yq9
A79JVeA1KlzvypsKzZmPsvP9Jyda4kVgC0GKikVLhZ0Iq5MuM0fl/yzc3Fd8
fsYTOXjkvNdNbgMqSi92kRCISzCw88IbeZnHT/3Rl7QY4IIP53p74BmAL2M5
Ke0amCCDmWWSQscYUakTUmOQWBs2Kd3TOIUkwNI+jSvyK3FetiOYOx5TN/GG
gjDRp5OOR1i1G/I0lc4N5RWKZJkCnaSIfV1gMxdkmJkl5xsNGIyV/lri/Yiv
Z50oNL5b3TxJFOWKAuj5gdyZtfCGoewFHwM+dRSQ+qY245s9mY33BjL7YwbI
g+ybxQ3RlOec8MWNdfiQz32AAZbDsInuzDqQNPl6E9gfKvZJeISxU+zsO7TP
63my8Ev2cYf94fZ18HVMNxDFxTSEVdSguiaSP0anaTB5/x27lRQz44BJe2gM
4zIeZSCrPMUxtkn5cYkdYUvhXD9Xpgi357Qd5SlzYc3gUDag3R/Uoi+zI67T
ooPy0oBtJqc+LUH9Sjl/pctZQulGjkXYdqaa0yECxDd1CSTvk/T9LYiy+a4H
j5JgOwb366MWZbhty2+1s9uTJyJzmVTfOiUcyguED3mcpYUP6FRQSUDoL3UV
OFroPUL/OnZ/8ItMrjtz+SNmvijEt7im2RYD+rasTIaKa5YInmwx2DQqdeEI
+MBIPtc5TfWx6s5Ih+uo8iKFJwAY+6oyrkUBF7ViAP97eL2TsY5JYvIyFtrv
5j0ku/jLag5tTh4jB+p03VJ2RLcEDcoFrH5SyKVuFgR3BmGqk/lO4VX91We3
ovQu0nRwqmbf6aigsPbZGzawQt37afVCM/q2k3h6VjdhwjStjx5rIGkKWlFQ
eR9bI9tsOq0y0y4MkzJ28SW2dQSHWtpss8jubjvwEAJvkYuQ+KHPUdYa1BJx
M1pM5apXtAvsquox1u7I6OzGOSqyyuVOTwk/NL8F0Vb40W6uuiK1H2ifGFMn
Wxc5tlIlSbaXZoKF9AhZ+R+hg6e7vmua3y3R7sBdF8ODwoi+vOYYovSUNeHJ
gD5QVC+LxvaWmLaBve2i/WjPjcP5g8SrmnrfKmWxXcUac0cN1PPNwKU0yYUx
WWzS4Ll8LBgfVjcWjfZMXICpnCxqbp08Ib47FUNikiGDzgSBxjhhdCrrXtEp
vKQzAHVR+R+z0D4N2D7IaMlFbDcLzr2b1HpxziYFiembqKEYSoXxn726CgFO
f3a60EbRLb3IpjbvqWEBbxbXveAf2MqSAPL0ro1JjxCfk8ieLREiYd/XUSq2
PqxMZISveiLVzQvVgIYCjJI/3y115Ul9vNu1OFtcOgKoPAQExly4Jnc7Nzu7
3aG6voOUsdee8baabuywo0yGnI5gpPU2SJGJaGhR8TytwOSfIq95GX/0VNf8
0n/QNF+BMUsi5UczjfTbTVgJWLbyF4F3wkGDf676eRJZ3uUBmjdbc6Aa+2JR
RpLQUlAftsEDd64HA72DIelQB9UB9mz5Anv43zpOGQq3cNlWuYayhNsawS2i
jPTKcTR8gGZpG2xOkas5WzMUorrXryqrViCMaK/TWl0RUfUUijR+aFeFlAi4
eOL+pxnyb3Y1WoIA28fnkLGI4+mCqF4FJs3FCw/Xh9BL1AaIiVycVjH2z7+u
SA7zZKZpoIKWXH/oYQtnf9pT5Uipxdwk/6d5pPR9KzgI/OvjR+d+07ShNGfq
hgFeJemPFPQSXZ9Ht83Z2ICcSubidpUzP6gq5gj5p3tfc6NVt0lEK5eFAxTq
XEEcwj8M9B8D8KP0UoEC6GzAxCMWdrNbGIn9Qx4wc8oHDEJizVsUw6HA9oT/
77EHdl6aaWJiorUE2T5pk7bgZ/a5cEtdDBUFedDvcIwbWxHQMsPMr67QcDDe
x5fgkJG2MmnV4NFS3RBEqtE9fuDXK1kqnp3jPYf7zcTHwkBm1bf3YHXM+2va
2BTocmliFWYFD6HjtSUDkff8vcEpS/M837lE3tjqAoDBGTPc1klu0sfdaWF8
A54/cf4/Pp/seQ8pf0RIkFxiGhZYDucjLBLrXY8YkfqkIbGyGDolqO502C2J
TrfAUIB52VP4IDPq/GxKoTVgBOORRyOYWZVeHpU0vfFs4uOAHkCfut67LMZU
2qFHERxwg09RtR/Tf21GCUqrzNPDhSVwJ82ASw3ceUy7839GcA3A+KsucIFo
fOcwxk0U7HzCTZvH4XN5P6dQ+8F/YI1BFZdR2J19EltHkMa1Vk3nZpdAP6sh
J86owobndi0lmDVQ08ku953Znf6wmBVhx1kKlEABL0xsYQmzRSUkuB0JWFuG
ZVLfhfyHAwPBo8bEJI0C0+IfdnBF0DFtyoxHSlK49bCuGyGIHTFvox0DYVsI
9l+rDMrrm1LJUR8EvRH/ycQnPvfgXYGbMvZDzhr7egQzy/dIifX7UvkDKSkB
VxtZqJWmQcOuyymlUd9tumwYQaIkJJuvoswIAE7s3q5aoZQaU760qlERK4Tx
GYHQwRGYYYPUwci85ACFllmBwXk4e06z/0CQ7kqiTKJzapH4krXSUNBMs4DF
BdWUvsqMCeaVw++wvUT+FnVKFtEUNSv4rXRqFhkDonqRLRcVUEe4k1wfPfn7
6wIv8oTY3CF9f57CRo4hq+WoW+8ovb1d0X16q8IP10aeSluigXeM4Rlrle2X
VG8RRICLeLcXwVUt1xfuRI9OSE1WoSxXr+wQAEQh7Rc6JTvjb/P1AOOeGufx
rG9wJvPcdiq55Jnn9+2NYygKbKpyOnz4gsMwkiXZrua6yFUUkQFhCPrBaE5L
xTglHUBPRRwqza605VjCcGZuYmqDgmcDIGTSqmrmPcM/RouZfzU/sXUTAqNY
YK1orzEFQGDwD1HUlkc3DCskmOvml4NEJEqCP72fgAgsDLjQ7RW/WqcFsT5u
v9WtgNY+yLwJbP5Lw8CwHS3Bl8qZ7uYxE2LzcMw4NSiz/+3E1co0wN3ejqoc
ZPUBwvO0bIHieLqfcwL4FF0n8TMPU13EL0cc5nQPaP8ew0iKqhtltfnCt+ZK
5OPi1Pje6YnlvCkHb47xUC6KHyKMFhEDbCaTJP0KwcNN4ZwjB8wShO6UUqJZ
RIZ6UhY/fvGLA9v8Fxu7UVKlGcjKZpbNJluXpzT4ynm6xyBXMuEh9rI+PUzT
6crwA03zHSJaRBS9xhETbrsE+yhYMjw1GxgIiyxA8g+i99l0HB/QM+ABigO9
HlYB5GDtO/+3UNVBoInc/Gv0/CsYlP8D0JjFmW1HPSMbF+KDOseuOAaY4X9z
sNwPXMNlNhz9Q6nYLpRzONmPkP8Y3Xa/q8zg6pn3IO+jIScMuJj4LDalgn/x
5eGdbjsfKxJxKST+P3fdkbhjxyHTUjfirrE/1jFxLR690VySqMw3sG3doC5q
9mBEHVmlxns3TOw/AYI6cepOzu3PFKx/8jEjNJAhapGJRnFZdrKbhF4rAuAT
6ZH8VNURZ1wQW+ykbcG+g+rXc/F8RNlhZ2fjxSYRa36y9Ok+759NZE8qVjCj
AcK+oqjEWnceimqNAk+OVt5cjIYWo1q07GoRizrvVZrHrq9Ljrk4I0QccuKp
2mEJEKpKasKwBmG5LiFJUCF1WZgCs+t5JrnJR+yApUBmwZk1ASliaj4qNXiQ
FxtEIDw7JiVN801CmTvCBWxcMUGSxEBXc2tmMhsv5uzxzf/pweMEKGVbeOvV
OgmTqc13F8/blRJSYK7k5661Yj9FgE8wGowd5xWPv7CLXKYC61hiklv9Pe9r
3mPWPVEoFjnTdfGTqcckAZifcGks/K5eBy92Hsm9FXCtD9ERfi2xdWxm7v3c
qFkbqYOSjSkm/qLAhI/Tns3TV7YLjUTaWLpv0GoNXVXD8V3up28aSZVmILI+
plgnIc2nyAu/j4YKdR2973n836ZuSkv2H+fVhGz+aMjSUkCYYe/JEH1em0Vj
GyZR9iG62S+KzCSO/HB4pTmbY35hT/wOLmxXP+TPYHFiF7Joyv5xcwjNCZ5/
FFuTGrXSpMm6sAjiBYj/8WfuxM5q9qndvd8y58ebAMBitdx2WlUJ0/azZHhd
/LVFaexjIBxvB57Myf60J8Vc4QWrHrTHYwrfQifrRTExSqCH6g34P+Iignak
vHaYKvbRC7nHnDnvs9/1eQtZdXTh5q0nhn24e153q6Q7F7BfA99OT8/Hl2pd
rdRmT6OeHewmyAUN7KYbUKLRVLVcj4Pi/vsLMIQE3b3OdxaGPQhpwLow3+nx
l40oBV1RqqZjDNh6RCeUYeahQ5iuMPoe1F4SUqqPIbHiTv8TdPE1xmJoUbOd
ERe/p3Ny0NjHplr6Z7YwbmDVbymF2seCASqOmXA6JgQLTfhfamxCXAyBwh/y
QgAOkchAMKrMLxGWCCtsVX36/qdwvvfgfpTVnocwrc4vhiRLgRowmBYWrQ/5
6O7ddQQWecSwNlfd+pTebKnQwH5Iv//Ej+e0+eM31re6JGE48XOGlX9oDRfz
J5pPunAmjJrqdk4Tb1DXHKh5TlBdXhPPYbKhL3sV+9xuHvLbNE9j1x+DUHul
0c/JeB7ax28sDFi3Hn/ksR+JTgkkxlNWyCKne+tYyrwRjIEloHify+z/6wu1
Ez8W54fFUF+6DP+YpFRUZQ0IxArCQh8CLsrZb/nplg4dNh3n3Sd0TmDUxylO
KvMKi4Sl36a1YOmRLegZiLH275CI69Izfln7kmcpOhIuFSPCUSpdACBV4T+v
UjC0+Hw2/ShCcYdJsdBJqnjLEuxnCmbNqMpHvqRS5eksSL0/00sk/BJYUZI0
qf70JlO9JvAW7i3rrKl+mInLexcBUhj8YJdvy8GFbkMsuuH6QqUnK+sCWDOX
AKp8NPkqEmi8jdARfVZBv5ETpI2mKvSOnAIoDf/s/KypZtMu/5pGK2CKfwiY
XkhWF4U9KH/h29sBeq43d98n4VRIdzypDVMpU+j+8EQE/KIEbOW5p6f++yqn
SPOluD6mcW82Z9RRkVaU4mQOpwzeKzQ5ghE28QmvqoyLVohfu1fPWEsPL8nv
kp7RhW1507m4QkS5qWJoSZ2KaNdS9JbaI5cKDsCIiKtTdftYERfrUkqRER4f
KEx4wi8p0tKhH4/mDGCnTN61SidwH/kH2gJ+4jp2+OHAYshsDP7CaryduIRQ
ukezS8k2yLcWRF9njS51/mjlPjygh4K5w7kgGm50AtnoRNekyM/ISbizaQa7
QtvTkkKN5UhobFRjB5QNFXZ2xNrmjBJhX4P0ZxHcnrC8f1QI4dsbkfKcfL2s
5OIUh9v6RQMjEYAArgbbX8Cabqn/en/1Y4ZJ59pqxQEXhw/3vp3yLotc/aZ+
H+jMSdMhmeV5KpPCn9vWOP+SMaM5eTepDo8XlOiGIZ4kIGIX8J2pB8yZNXQa
zq8YkzazcKw7SI8uStfrVzNlecy5kWVB83gLXHDeMSDnMMNYAz//28kXI1jt
/vM9WwHqlEJ/lDsvASBgcc85CXcRDofoNNPGmJ1SPktEpah3oYOR9OdMDkXD
KfRRmC5EH31jEX8ssO+OWMISgYHC2+w605BAzzBroaoaviUeDJtcUiSjSVcc
bYXHK5VYepjJ3+Z0UpS+1tY/0fOgJAyBfQmfB9sQAGMKLW29eEHeMRBx44Wd
YRCvvh2m5D9RAlQkve0ko3QwvKmzX0nt5zr8XwOOfgUUX7L53sj97MNnzx8s
aeTZxXRbOtWF/CyGKSEaNaiDgKtjHa3zX8qqBe7IQUAGUzdyOUA6Yflcv/rE
hnWoMPwNth+kYeggAEOmDUqzQpQbvDyzLV2BIwBzgkrCFCG4SW0k23nrxD9Q
yvzhJJ6cerueNV3KuaJeStF/rL34neErEOIy68bk+sBk8rLvMGKV83mrmy8n
Vr0sO27crpsHUhqmeC7CxzA4KV0W6VkcT9fDayrmpXqhjcF3x7p+SaAjne1D
PFg0jtGOUKExjv95RRow3REeBtjj6l/c7j5vVH9FS9A5qJkzye/ck5KetNEm
JtBynZcXe6y9wsZCZZ0qY+uVf3Pyi0SrSDTqXJWd1VHHbaKXwumdm1C55deQ
o7N02bAS8X44/wwnZm5Xpw/a5/FOgOM1WVg1F9YuPYTw6I0Kh34pYh2+gDd9
tf0R134Bi6nigCfyJRAmM3osz7shM6IAkZ4+4191Uh9Z9MW495FHrvvzepYT
oMziAWhzC9EbBe7YnVs1E0urqG17n/iMNWZT94gBZQMaKMul7nWuUmqD6l9F
AsZQkpbDImQxZMjSrnFN2jgJHJ3c+GI+c4KsMspiIqJSU2tlEOVETgwFZrsI
yjhQZwA+NYqtu08xwKM+RDyXuuNBPP4YqvhIueijcDI1C2Dl1bT78/IVAR/U
Y4GwnWU4DwwD7SjlARtb86TXUXBDJHSncAdUVhZgNbRzAiJNOFU3sMehAdcB
NNH1/AhlD0483XmHmBVaCsKUjBqQ2ANrFxxP0YpXyTFdCgskW02oVWdDOLLd
kwlzs/9x6KoxIU8wz3BquqlmAeS+dyMudUu2ZrLhB0jsYVfWwx7ZM8aKNV+T
NishG89MEQLVZSj5q5q7YHykUMI8oQuUnzIrPE3bbxfOg9CBFyg9dA0Mtn1n
VGL40/MMnksIoqcZdBJj1kBnV7h90A+kJMwZVWEoRCXcJc3Bs582H4o6k+oG
b5rUYUhUANif7H7Q3X9kMIPchhEK9SVq1XQ17KDMnnPjNDpAPEKCfWbJAWyh
3GjxvGpMQ3y/c8kzfyC5MBgqD22LriTUHhqMrHYYSFHSDMFubx8oKr/L/HrE
pnarRZbSldxfmD6zRDsFhna2afWwwiV6dgVQCwKBi6pESAymcRR4dS1jtqj0
ViYyKmPUTIVXYEiyCRVOTNNaRXohhMtYcZPg15NgFe/MBLKdkd6YyDRhBrMm
rG3Ooj6JjVvF0RAQIDDSDy+DagHQdqw8nz6sJzkrAGTi4u07RZXDOAY6WCvt
F+mmHIt8FNeM5PyIPXdyZbqp+h/2ZyOw72/pJ8z/2aHm6uK1L9CAtmTnPhdZ
QtEd/kGGJAOlB1dnneQl3Fc1L1ZEiAavEJN+R/6fCJpuNv4x0mIWZGl9mNjs
pmwzH3qp2VeZH1jnf5dphyMmV2MR002jkmLc0PnMrOa86V77sRZ/ItjIDAgZ
yRyPsSBKSgn6Bai+bnH+FRq73oSmf4NQ/0Qr7iy9kZrF6GJ5AG2rJTXCBnuY
Fr4d9zjpg01MDeACB5Jitdkx9NUUiYk21ghkBkS44lRQLou5X9AbbcnjT4ra
YVXrTLP1ST88BsdyQCaW7IipI5Dgl3511U2QYOaiolOZws9AYzEPFLXmqM6I
PciWVUHO2JXfaMS76kEBIS/sF+A1fWhtr7IJ2DWzR4Ke+8pxoNWjTa0x40wZ
nVAEXoztOjLDYb/Cr1GcU8QR4iFBRt25l86PmknQ6uBR62Dslkyx++T7e7tx
ID1XB6Oh0YxnhiM8QRtUJqAEzoQyH1wiwpRdpCQtjVmFUYrDDhZYdLIg9MII
5o7x2MceGZZER1z7KS/jh+zVSyoo4q9XDFSX06lBOSuMNYwXNq+eoV4EdE6x
ksEJYTpkMLlWeUWG+Py+A4W/2shPVKz9/BxOpOJgoVpR68eI8xMl5Sz/qZE4
FbBwZDGBZGVeeayKy2kuU4VNKs0NslTGtohNsPTBjLdLL74v9Rbt0sw+panS
qfpwkh/AtoiOJ0ijHo/lU2Ty7j48TBYrgPmi8HxzsO0VYLLGQD1i9mj404Ui
Y7Lt7LRv+BwwtpX1BdAR4Qpehp0XfM5hJmsJ87ul+HU8bM20Lg2MuMMggFqL
2nPrBT/CITmhilGqRi7DbRuTPqt6GzY+bf5KlrSthKLs62wh0UrUqWLZZtFV
COtfcVnveLvY2ctHqO7j4v6PxvtMVM2jhT50CsX2+8JmWZKp1AOyNwx1Ef1q
hSSIuluXb/9Fq6a1wD+YxXo4LfyISePmK5LRrib/8UYwpwxoWOVVrif8wkZr
h1kQPLDtWl4ZDOZPsstLO5Oa2/iu29xJA2RZ7Bb+qidhIbI1JWiYI16ZTEK2
yC/MKywTF/kLkjUDgKdwPcU86iydwwbIl43ayf5Xm2zgNADFF1vFAY4KcmY8
gq85dz1E6SSThZNZQDhZ69Knf2tkDESj2jT4JTYCFhya19MwkbCD13Aw5bCx
/RCmBDtFgNG/jxgWutHGFRZz1ejtwi+OG/CGNvx8foqH5kuYyI9Y5wE8HYI9
Gp0QdtEqPt2Yz9oDmNJm9C/hQXt6rfu1n7BfnRyHx0ObKl1jatsfEmJGmAB7
z+W4gCGz0YMs7HpzUo9nLLqO4pnQMioS2oRfF5sIqL+Yp6aFA3lBVZmpAJFt
qrdKWwYXdB07qIdiKWTKpXd4oyFPhCZZZWOjkCYFw98wYbu3amJ/jF+pL4Mr
0UhTg2xxCIYFUI2c7xjsU+SoGb7jNQIay49CRlufzi4bwWsaILO/TsZol1TR
fY+3LKppggiS3BP3wLFpvohkqi2/pLBlQgJwWIen45w9iEXMJ/0PncLyvM6u
pm37brlkC+UGu/zaKMlAojHyb+07TKoZqTNwcDWuVdq+zSlptEnUIFGcRl/p
jmtD4y1/Evk2L0A0Ltp+hqV9ECNgN0BxA1evO+0zOLpStsu9G7xmsrBHAZVA
eearuu+pU2rUEqFZ1XCif0dt4IbPE2Dw7fSiKxcegBXFqotV1TKTTf5rHgVe
bAP+ePRLnjXtOAEIzx9Q8iG/dW1XX/bM2OvUYW7dWWsnPIXFwszgj1kj0y/g
KgpmXPyittT2ls6FruxXq9CT5AGWFC/8uzhoXptgRn+nG85Ky5KNJPqew48Q
wIHJ3PQxG2KwU/0m5gSVnERa3BCHZkqEag2ETYwi1GAieHADCoXezxWFJiNm
i2VXkDkuewjKBGj0PWVqvn2G2SuIrxzHZwRMYQjee+vVA5tCK1AnoONPfuyp
7uYMehaUS5exg1OF4NebJeKa71d/OsWQlidOWSDGM1bg5DM1IDL7/fZON+AD
XjVcbZYj+YRp//KXECv21jPt77Gb4SIuezdA9rq/P6bJUWQo581b5qw1DVE0
2zCGxtIKQf10NZIZIqUHsjCy69WzHhJm6+M/YpgtGWeSB7H4Yshm0hl/hwny
Lk7TbfgHSfOSARC+PQslhxb5GOvAMxW77LzxchXELaqKzl0cqdFrX8hyroFS
stAsNa+M3HmUkk77KVVrUIFGG86OnuQQ9qRK0h7LS3dCuNlYiNbJMSVW69Wd
SgNe8XQ63D2DVy/x+yog0Dkj2rxz4hXgwFNnRgolKEZJQPP6SU1ldVxPulg6
frbXJ0QFYzxwBDAHZqc/De0v6wV23aqNnyBoKNeuVW/FikHL7ELZ8QiQl0x4
WacQIEIPl7de6XtSVKxLfnIhDIHkFV2WiGn6xKbaUxIL5geVwi3EBhS/cgtk
DJLTHf7tAaVZUS8+smNsg3qzRst+NblsbGPGCUIf7ZF4eLy7+RQWQC5TJTsT
JQI81mtd7GUzgyEU6H+VmRYp8T9/b/y9lP/kBp3kQ56vV7ie6fpfFQn8Qzsh
CvexUBPNh2vYPcpR7/ySlPmd+Vv1eFcSKRKdG7s/Ik7v87+074xibRatweuv
9DatrC3ocSkKjAkKm0RNIRvLthM/uVpApA1p9odIQnnmVP5kX5HUm0cZoMlD
MUq3NLRf9t3k/FyEjVlk9UoD21VGVSB14z90XJdV/h1xNOV5pB+JlO5Y2JFy
ADVSxCm5FIG+mkgo0b2r0XwIFRuVXM4LpG0dG0FufH56OgYgJejIkxTSZzkW
vNcYOBl3DupOIOaIrjSPMoJodxYoMbS25ETcIwjg7NOttUYpiC5ivTvWO7/o
ZVB/gdcVUP9v49jcys3Ja0HB7YbpHrCgXB3BlSOtiCdfUaDe5M1IVXxCf5p/
/n5Zi65MeExAduoQntImLmcj9yu93+gTF7LQgrhAh3Q5RuIzlCNevufbbnqX
rpoxNozNhfTy0MJwDuy5sex1GwYNirDDXuMi0a1snjN0qt9bFnrvL9fOYcgd
ZC8lXN8aIWxyqWZSjAv+IaKeol4oTrajgfvYfKJdUvZYo1JlRPWOyBRSd5Yc
cwc23rpglyVc3WIp+gYd/asKCRyBXH7GiD9YlF5sSpwMvNALCGEir59mQntS
J9y2gQt1MMu1oh7xSWteg5Z7cPx46IOKc6gB6Tf26f8g89MBpqa1Vv4Rq7oH
SSez0Obi0pMWFFmHsyBI6MniSDE3kwjKyRACPAdUUXbmrppRoCGGNZ4dfzOt
zOCGo/Z3ydPRksg1SmWk82BRHEooOERzEGaJnrWzr6xFqpTHczX6TdPKy9dK
s6Hbz3RDtSayFiX6Wl+aDAl5jBUd3bQcVCcMacNxiraFTnItMHvmjMFfv9VB
Dhhpu2oFB5NLAtei7au3D8cNtI2tQOwCjEz+YrEn9tiNjwW+dJKsKbWbHJbT
oxcQAlJsVBbMQwVhmrmcfq8ZBew6fzkmM/t0eDzGk/rb8YO25+hY08dUoQo3
Bg0H/7O2RLt6aL7fYtNt0j3afDJTj1cSQx7i0U6eV/32eQIFMoEqcGQryC3m
ul2kLjRMfN7Yjic3yf1R7FzwXKDpS30R5iT3VO+1Y2GcoxnxVQFbbDr/irOd
bkZ5lVP0ykwV5nlO/MzbKTSrzqo7DJGtsvIt7tfCWXyLIFqSyV0Y5HoHM5Ce
VQqE/WUSkt4choMpI5AdLAxkhSFLvvqTMx5Pnb5ypJAcpogAsEn9kyMTgG2o
gba0mtj+Jd01fleW1G38Jt3FsvNM7xzZQHKm3OqEMbg7QeiSZB6lLpbleuFS
ZUbLymnHaUEiZDiL86vZE8gOzB1zonsN1PRQqqpGqE0d5ps/wNsWFcW4/JHM
g8yilcKiyYtLcb1m0ylBmsWsw6iCK/B5JBcmkjLhlqreV94819YOxQVOhe+3
bJS9Shm/R53HvF8lIbaDsJoP1HIFRUn8S6hK1CWrhvYknc1maGtqvuyFAwGG
O3ncEpSJoE4rC9PMptp+kBUIoBm2OkShL/6VVJVfJOd3LuIYvwMPHiGVL2vd
CrdH9DQu+Bg+30/ZyeC2eCh2sZgjVQzldWSaENWiysv8jZfjyQe5kpPFEY9T
dhQavbrVCxdSFehNti2AW6mSqy8QIVdfATKZn0RnUOr7T0sADbiPH3TOVp15
4VZMIzJRmJKngSonpkTfSESQP07sy/2DondSvPeyfPAkpHqNy+I2qe7hwoN+
6eiv/cSzQARAbjQeF2EUtB74x/LN80fljByRAxcw26gu4MpL0G/Mplj9ND8z
sbEbyetQIzgfml1Hy3TA/ktAOV9Da0hIunvkHIpj4nPDSDiPKPnOh3XR1o3K
eYHjWQ6mLq9Rp86T0AQd+VZBqRYotbh7aKTPHEm4rbyIr+PqAk5GzxDpX5LN
iUdRbInf4rJly1VYEHV9/vElPngTzbRyDqM0fB2c6KKKiIW9RdeBSffnHH4q
utNBtc9ioL8zSQ/RwC8LLNJ7zkMAfqZmQg/lsujw9rJndpjRGWE664vhxtjW
NC4JjdYSuNfysxwZYidCnCJZvlcwa4JM2LaWwlGjxA/8biWxFVbMjVa053In
nprYnNxyRclTx0EWN9Zxdc6Q7CD5QBagLK5+1TU20/qM8X0nW5D5A7rupGQh
LBWDwP0L8r4Qc2r2ael2Bt3KEzSv1fnhgG73mvKo0kpJ2nZVs6wH4tMkJ5ij
NN8qLHb6y3BmWYDQBhbOTeWurIkes6ZkHObGNLLoH3pdJQh+p6VeHKoYLpEW
nudE1PIl5hSYmLkfxtVLENAqo3jSKfvXF5+PvS6DjvipKe/57yChQLGNARor
sgC59Irzv4in4dPL6e5WXo7iD+SjS5ioWTzIdE75Ayjw9TQPNXwosEHZy8xZ
AYCkZ2N7C/dUQv37fe1I0GVIBaMVUiZbOw4yJ00i7I6FlxC0a+WJ83hbcKwN
IiysZ4LKqschZokOMnbVjSy052fc56FQCeB/59LY/LpAlJZyfcqV3vZuLaUn
cquJJveTP7ePbReO9gGtCr3nXsq29Hgbw9DSMJAY3Nb+6B52Ij8/BWlls8ot
ODLsn5Nfha+GTm1mFhcKEwkzw9HS87VC5iGOfz1cUAE9nM/rxqsr60tATYzT
/U8VcJe2+f/1yhigkxizlgXojm6u9II/97liIJQBUXRcyXhnxM5o8nZJG8Ie
amMFnDY7+mof7Hr6wtilYb0eL8kLdCy2+hflC8aUg9O7/L9nwnmvbE5ROM5s
ot60sO3DtskrNoBbd+Zv+CwoMBzoXZT4wtSaHy6PshGsjG6NnXioyqBZxjHy
Gl9LpogogWNKWJlM7I4pS9Vpam23dEPT9RwmMYGBNEA1is3qQFCMmxRgHveA
GaMQM5cDbhN4af2uKdoJjnXIRJyfySeSusKQ0fI3mOLDrcUfK3+XV6DZVHPt
+Y551vt8cwEuhs60Q7XnX9wToFG6e6dOAbzwAJdWFVrHMJoQTlvFplmKhxwv
WTTWSyXfVZUBvyDfjYTEljx4vrdU/hJLd9xpLQLY0T9bNMKxcYESbRm3FIRL
0QK5LYsvpjDPTDTWJsbpnugdWtrr7n+VRXS3E0vhyXL4yJbd31nJ64tXakSI
qT6FNujcKyLgocLtsfru9niEdGG3cGz14RDRNO3NaWameY6fwKFnqZkpcxkq
3A+9guaW3aF3SgY0W9Mr8t6Yp1EWVNZzU44PrL1jPU6JOPHdKif5GRuVayEF
n6bsXJxBOM+5YQ9HsadB6d4tyzItBk9Sdcnnknrs9efXOP6knUd4agMxzoX/
AKGzDqDJ23HcGr4z78+vUXDtw4Syr+yP6b4CGmuLbzdlRjtxEMOIbHbHKCpk
Wp2VDh3/M5ulKe0kZasgw9vgLwlD2BUPx76OVt3QbTuA2V0iI4r+jJQ4eaXj
S6w+dXAEGOgbAR9eQAUlm7yurTbznNK9E57SD/aiZ6+4chCOC9Bx9+6/mYI4
rLId+6iVy9SYPqZYruAEgbXuixPFuNQozk6mRbwOdSlynefXYWVvaT1y/3GW
g/8hyNow4Y4atr8oIFyUodGVcD+nyzviMdF+cdTBnAcd7xf7m5BIKx104SI3
mJMYxb1DS0OIX44RnL770RQqMvlBvqUiN6YO8HyoVkh5nD2bUdVtWySTXS1F
BCQVmCDtrzNnvN9p9+LzLEXf/M1D8q84Ej+ylmZAW84/2tnTnL3MSTi8TPbO
+ZYSunUPqriYoGATOsXMDncHNTIKKCAySaXiAdtsY/enwoXzM+Y7+bgKsMPg
zjil3ByhyaqLHqDs0CAM8eRbvSQzXAD2oAAIfFDVbDhbb+tCXR9Q4y+aw52V
MPJ24SuoQwPI0o9l68Cll01PyKKFZJkKiRN1Vm5XlGrG8E2LLnxQzAd9344u
FcG08fEDX9ifpK25sriognJXoqPP7OjlTFqlgBRF6BY1Mv0qzMkZSCnLx8MY
gOmEdHyjwLWCyp4n4Z655x5uyJf4mNNbEOG6ZePsx8Qdbt+QhzMXrOf34ywq
iYoyvB5WQ4oCBwsZhPuLCxTL2mNA9V9wOCWL2LnzoS7zABlV0y7p0Xe6we0x
Rt5AN8iAX/9xagfG87RyVSresnNC6r9NcGZrnkqofXpzrEoP5MuOB8bBDimx
cg+hUdoX0Y31mutpK6vknpTBsl8WwAN6BWWik73p7tjRBrGsbGDbcAiISuol
idTVyi/2LJ2hBaXdFVsSeh3Zxhms4CrUCqSw08E5vI+X5BOeOdy0BVQmorks
L1Khn3XPzTbMeJNoBsqNtthwBgOoGMS+q4vdNWdy2+VQg2RAIbrvjlHsOwbo
OPBTkJFdwv4HwF8eCuZhPn4C3JO+DtN+MB/eHs0uhEiRdmXgOZuz9nSmsvFS
NlD5VvMuhLZ1xYE/kMxeJfrClLpt9jLj7K2Nyvk7FS7rwxAXqwMit0qfIFfZ
lpqZgGrF2UolskoBmJKuv8e8g2w4R4DiRXPL/x8YkLvgik1GBert82Z5JwI5
pJ6tGAEyMeAWeSuGEb4JCAhUMDTiGNKPPzDulupPTb+UWTbiP7pQnjeXKPMu
tLjlrWd9Mdk1f97FcGL1Cw94zomIp94Ldnv+9z6tWtrpkiK1l82d3mrEIkV3
QFnBpfGrwQP1Zdp/bQRyGGrq/6CeiY3PSnjPH3cHSOpeUWD/Eg+5HSj/0zRR
43Al4MpOimQyR9u0hujo6xxlwgX9n6jBteszXuKqI74nNkCrzOKbhVJEAPQE
uMFNoN4Iyhfl7jCK5Y4y4MICG3FaiRfOl7VQ+oTKZFV3VJ0wfn6Gfwf8QiXa
LSUaVVSOY9SxMcTJMVBA5EcAQBIJ2ceQ9nq3A2+z5qKhV0bVgSZ+67a9hEJA
iGuiHHdxKhi+Kr0u10E4g7m/NwuD+7IIfaxEcdpzSB0Eqvt+4EjcCqPo4PiK
RxcoAa5uBfLmMZn8E7cKNY4FtzFUtUypOaQOS3vW3K0NKhhdfEyfsYG0YXzF
Y+NhggfjK2YCvE9+SDEJlMc8BjJVw3prFJGGQUzQ8i40vkQgGJbPt4KeBwAH
xjZ+4VgIV/C8nDJ0zgylnpaIkYfn2lbEqBu/8JfIpdrZrHDZA3EAwK7KUEUD
wp7/h8Sye09yFxk/DZl/l8fOfCFK+UA0xzQS9hynC5D1O82p3VsR9NAB3ami
DUie6Z3mUst0kLPt/WACqfCiukRKYvqR41LACDT/A8Gok/mrf+GqV5LTjnxM
+2DLJUlyJPNeqLg4dHnRQIsGYjGvuczWbHZoBo/wUq/nNg/fzuDs42EUrG5d
Ab0QR8wChWA1rh2p1DnSNpyllEFbE4vlZJ/rDbgfMHN2vBOVAAWoW0F4BjqB
yNMtue63R+ie5/kXVBNbH9wY4Rpg+BrUKhAkKGZsnEqBrIm2683cLn4gfcvE
gqIBrP7TUVoFyrtjGvupSwD4IqOV/a7F7fWhqqf67RjD0gugciQYo2TwSBG3
aFttDd/XuFzT0D+OTjhHyQw3qq0UrZfaEuEF0hfiaqNxnj72ruooRGQ/RUOS
IHx9b/YrC/SSx52LU9RlzR3HwwvS4xRqdNHmwgEQ3pkZp7Uh0U+Bt0Sli0pC
wphq4nUcOUb9bseAkYYyK+/6FfoJQJvjXa8So6IWARoiawheOPhldDkcwPT+
vcm7b9l9ViDjloAKRtqc2VwWnnmAP4585lIr9G+4aPnlkkBEkpTWHdB1yq9F
0x84yPdiXie9ZKOLaqRZ4Gxw7HiJxARnuQlZrqZ1K6aJTxCksXhTmgsHpH8y
SKG4L9oUX1HZ7aCxkqyzVuqsrqjPKp8M/z/7qu/d+bGrqrGal/ncKcM1lWoe
u/AX5SPkUshl+DHQbYXEib6PPzPfOiiwkhZj4hjtlUiDX/GIJHM+5bwe6Z4K
aPCsZzdcsRA1bRuEtiEuy6muCrNYWRGdHRwZFSD3H0Uh4jPuz8CpU1cuIT14
TpK/BMqPicNhYKOLHZFggML+CcfcQG+NMo3W6Wx7NhPSoT/Mh0tBA/7BK7mS
WUdjx6/qpDIEKweKIgrcE4jPTFvomijiL9yxyOxIefi1NLF5wJEb2AOZVbaA
U+fLnMl+FY93Vlt8tEd4qrEx/37mXnT6xpY0lfwBLSBUV58LYOq+vdjkwcg5
f/uDR+Wf9uOlLMXqBUE/gTz9Dgf4L/nK0YF4uPP3bb1xBW9ijFUmpBUpS7M/
3TneZ3kNNS29k6Ivw0q80SV8lV72yZPlcIZaChol06BxBfk+1E6Jo1J+G21l
5DEEPBZHutUTqWHDCBbLKZMqVYq9hrvFIoV7e60SghkvfRuH79rzX/elYUS2
voc11q7NB+lTmjLS2AZVoF93m1wbbLiW+vFn76L/OWiehkvlOp9UDA5vHp9T
aRwlFaTTm+ygY4cnzjAk5B+NntsdhKUD90MPNKf6//9Y2okvurGKfBU/Em94
4GJe7AO9x2RmUonqSm5kiQTCVdOxY9Bsh+TKOyCyjvFD9VwLpWZidZcc0p45
q+F195n5azb/Rw0VKjI7G3kadUtcD1LFE9zlOjE2PVGw8DVIA6WRh36Hk3iw
aKxg3cMg08yTn9+dq5IpmlhDHPRXAZF4qxq5fS5KmuvOVtiwz4+Z6hHX8mN3
KBgkvscxahnmrDSvoamt0PYqQZFEg7ewbk2rmdS5BWVAGJYe6Du2x7YArN94
aYmRQComM332FYDYzZt7QchAdMSIIPtwjcj8DcNf29E+3TO7HDQCwS/6bN36
ETDOAKKX0AmOInbgyLbppZLIAfAtLrm1LYbKDXvus2s+rBfoGFcy27QTy94m
RXwqKkrKa6RdTLO5Fdgf95w2EgiOwYZ7gw/l60dh8QAVVFXYN0xjYfOPOOm1
hpIh73xYnjcv4saUhK2i92g23yt0nlEtDzjLSY8WkdyHziQtGEcojPiNmuLl
pDUoY3nfetZSyEUe5XVPCbyQFlrqeLHcIKPR/NQD9artOvuocaQnmtXLGg0c
QBN+Gz+2G9bxK0Whq7bcID0heAm5hAG1+Re9i5PSEJQUDtS2qrQeKvjuDtTH
BRCg8FkhU3UhQFwibMy9TivtVep7FO6gcYTrJa4vLqYZlzDhchthUrECduO3
lmGj1qr6QQu7fAF28TlEVc646M8Q8DAz+i7Nh20I7Tus7NbrDB0be1JxMPDZ
BQdvd+UZvv9MAIj/5RwG//524orNF+sKQKaN7i5q3IGhDy3t8Yc9x2Q0ySfP
kTUpeuCZsP/9ul3wAfuG66iBxSDWzhyLZcYgu160yczRIF1krmFdy14yCeP7
r5F3A8GDs356ZZPc1C8EeHomLV8+rr8xmJ/C6LbYxpQQOekN/qU86TN+ae30
snH+145KCFEC9MVLjf32X0FMhFgM1JFPTw13OVdG3Jo37oEO4lgVhhoF06hL
Ahh/AEukbveYIZ1s4AeZnh0tNGPqfjFGNLCvwtg5wIyGG5oLZW3sv5+I7jJq
W8+lem7NMTOXtHmiTR2HvnQCmwYZ2jFHqGp1WSxtHPEgZqlIRMoSeScSe+UZ
DXaiwiVpsk3TUTPvZ59kYl1t8+8WL4PotRDrLzu/Ve7cRGzjPd/CpjK/kN1k
NJRL8op4UB/IHhp+fDjhOjyN/nxB4Do4UmLlkW82TahcWgMVv4u9nBRjrUAJ
i5NjbeUGdGrH2xYXfNEa0R4FMirzsa2nSmWKG7J/5dopPTod6PbDxHiJLCIw
Ic1pbmMy+UJcyj2WpONKWLmZQ+J2pVTKtmeUptknH4S2DV4iw231jMrPsocl
pPuyx4LuZbq7tLnxyQk1a34f70z5Vdi+HfSF7O2NHGVUIzAGZzPLcdiN9OCc
OKvL4k1g2udHFRD5H2oEAvFyIuXOAjGT3IhWdUEZHBHLOwttnu0+5wC7IcVV
a7Sh8C6hjAwzRJ+DaGT7i/H2KkyH2rh4HE/N3kLXS2Volmp3mXvABkL//j8k
siHBBX1WkmzVNyTYNfCBAFHbMsAap108Yb1nKqKR0tyP/aAImb2Zv7KHWowU
MzMSAWjsO5vd6UE0vDAWdWTQSbXLyG0fU+VK+CSRzSqvetmzdGHjbw92UeMl
DRfiLg2OGqnRwmx5RxRdTV2DL/0hRHOVaublMJNbbAP7YjXKtofBZqPaFpr9
9dbHxWpsmsSIitKfTFmEBv/EQ2zc8wWYEVARddlOe1iUeEix7015OFdU2rtw
OawZkPeG81RUWL5Eg8Asfen0axEnBnquM2tMyEj/sfK6UuiGDyB2psZ0P5P5
RDgN/AptUqJ3PkTVbUr7BvRA7h8uVtwND/aZcnVt3+uqi0enzGaTEempLU5X
Nit5OQpVSEF0BDz43ohiMFmLr1i5VVy6IQ9eXp/CsQFuEv7etTevYFKL+BB5
CWJ8wiUcN7ASuguCvcJ53eLZmpxXcwcbBJ7P5vzZqgl9egez/45wkCqmUuxD
bK7/mUj8qHFwm12m4IkdaXusKt1RitDxIK07Awbhvz95+9gysK1W3Q8w+RC9
7RoGJTvLEEizG1mHT0sFASrIs1qzVTucisQwy3RXCNIxyb21ZrLsJo//SMFn
3cIejircTSaiIN92DOcUP71H1nW4J7tdjlEnh51SmEtA96O9pUMNmbo++X2c
ZJuEAapGDtvYG5M7nI1WsmfULYe6awGKjPF7qE6C2JDSTKLMMhv8m48v053c
DyDdQV4E05iEm+486BLCXqx2HLF2jqtPC77b3WEbq4L1v6Jo9bGROjMJIKZZ
2BCV0/Jyeldji1tKkB5Ub4ic2hM13GHwt8DzEnYeLKjmcWtIZ2OsV5aMonoi
8AfUNufmp5ugiEEf4XZOreF/2PwvuCJRSDiSOA+msbQOwbtzQl8MApKfQWMb
Tt4G7HI5T1IeNFjfS0CoZVsqaAEI3TO9pgsbAHWCnpP1qm6EtX2523Ahj4C8
jRriJVq5XVMgiSmVlBuvFJOOp3CprNwRPmvbuV6NjB7M63ur94k1c6YXneLR
UkfYz4+TzwJ/NV7ZtiIlcqyxiGgk2cQKCYkEdDUgDw+h6PXAhhdYAfPPQsHx
doNb062KLTNDUfXcSdppXOA++h84aaxLa1XAqmaxab98kGtq0ybrqBYaaIq5
QR03pGKKzGUp74vt5R1iEXvksmnRtg8o+0Z09iq2hyf775xkAnolz5m9F9BR
h63FhavZPf4qc0tIyhkkt2co8spnO1UOs5TPADfHf3n/0F8AYiWeKy3RJ/r/
/WnuSJqDsTfJUZUgAbtfiRsWnRFHHiTtbqkC5TX9wYKNf1Jr7s60Bi+n8Tm6
SKn4yfC33ZsPAPqPTsuilrRvbuM+tSZK2yUZr/PxW2x6bVY2qzf1MAcQdbfk
c0/0lm12cwh9UPc0T5lxnoxJzvp/T7E8iSyEkt3G7TlO2IMcu14Ua++1cftL
d8ht0FyQ2mU0oPdUbDOv8XHMzwTucpgQ+cMRd7/NxvsFjgEyA0JSFyhztduo
O/K9S7/kyfQ0t8dhq8bGIrD2aq4e8CeZBEiJldYoKgwtOdQ+hUXm4i752mrP
S4dO7oYeU/VKpaKSFT9oz8qDedEdLS4EvrtqxZyVnWcxCvLQZIHmAk4YJ9bG
N+NdL9lWJcLQxSmuVZcbeyws6F+3wr7I9grGGjWL3DadxdWTobt6OFLySRHm
pq37M8/KbiWetnJjVAy2iuTRwy6/3wzKjGG3/dtvXsIPy7zoMZB/1Lqw4Bb4
nNZXVfhYk4fssIqnybra1acd5w+e+3M7HimxFcDn6iuWoRw7WxaWbW9VrLL2
VIgOJabAgwL2px4wbzSBKUZ2W2lSXk4J7PciTfPzinCQ5noKZrv7sVUO/tUz
g4LomKL0cYCSz4MI71bpnGSc+jtL+EWCnujEUzk1V1hYqcAkx+xG/rm97CjT
W2oI28OCGw1oONUtwwO8kdfOofI4jYbd/cDqOK5aaU0Hzt4VEedVwgkFbd8Q
kDZkS8Rovh+INV3t1NrfYo+fyrvdie8H+RDZylEDUEuk0ifmHMcQKQ/6emkP
nryeB+G7o+1Y/+11q/FM/oUO16qifUD6ZlBMgrLFo2jlwYlkFoVr2kdO1SFh
HVk+SkUdtDySUg+QnHKQJi4jdUKEPochQu8Hdrkv7w9SqXwS2PSpZ8ocOYW0
cjFuU6+8KTPalPEQCUkI6gTwRHucABjCvPrWJUFTBf3/4lcaYYNwRihNoJ73
VncSIHqOzG7VGKHlL3A7XkiKxesNOwTRAP0lJi6XSjNRk8iAWeS/lz0oISKo
bT/Mhe5EFnFlObTak7jxzVBG3nXEomEM0j/2ITQ0kHiLRM0CPNLEfb5mxO2F
ylBfkDkkiN7bD0eTOz9ZU73U9JKy/1BpOPkcSOrqFlcXnTfw3bAKGc05LJ+3
n1cbkyz4+p3ozZJ/gCGrVJHv/NHZFkiNPS9S8aDRKUjNjHm6xU1rEqkkVe6l
kQZWG0H8T28QchiBWFEs5DuxCoIaz5amhN/S8gN5tkMTP1BkniG4VMag7eSi
yR51hfHbobDKYP9InbKvOg2XwNj+HByKhTTH7kGEg55iiFDDvoGUPlg1ocVc
ck29QmAF+p0RFhzb84OXJYVJCo08XctMnPw+SVaC0BntnC1vY1AUJnT8e30D
bNm4L2BXsxt5gfKgeYkMOONIy8OprgJaqbwgYbR2lcOvnC+WMS8WfE9sFRd9
EVJtX1/OSMPwIYP3O7Mmw0dgRlh6qgbOP4eZr64f+s1UiWecbT2lQ6fddSoe
6JaAXaDtbV55QUC4eEVWVnN7QCcwO7XuYYPtyYhcrtMu9hnj8rvsVOjXHADn
LTdnfRJ/lVv2PG6FIQRnlQIwsYG0p/OLi9trKU10IBrbXWLFg6xRpIKnA2aL
77hFoQkpvk8x3zd0vjVq2JMTyPR0/lwcu/bpYRr8Nq9GStgyiKSRh55ZG/0R
W3pXTAZOqDiZsIjB/mcNIYH8MAJ4F/866107NnOHQ3FeqLfr7bn/dt+9dltQ
LjpgDCoGYYnFepL8Bg7OGRxnm5oO2miqzeUZQtLVCk35s0YedP849mJjXhzr
BySGeiEqFmJj03sJgfXW9ogGhtVb7iFNNIHzZVy3qTx4k2+kEae0tnjlaxhI
pYEe0nxDi2T6ymlXYhHRIT2p1vIONZRTnAm7Sy+jOHB9zutLK5FP3HHHOskc
kvRTyAnRiXWgHlGWW2kHcHl/MCDLqKPEzdQ3sZoOgbsBEuz+T1eVn6agVl7W
yLkob5mm7mTVEet4unZDqC4N6xKf4WlNdQFGx2OlLD9Q991D/l/Z37G90Hol
dXQffFnxOwwa6RqNOOMTq1SticfllC4Bp0UywLK4kKciG18UydqNjGXlUePm
nIUG7NnF5wEcwL0SEmNKeLa+mQz7xw5WWj6P05/+IgTsBqN3LIbEa/jlNXtN
PgRdjcOBnHb7v3+R+KfcudcvgN81J8wbD90yytKh0hHvI9JBTVB1D9TpCvq5
R+0M8EuO/cJ/VjWfRlilm90JPhp2iNENcyFz2nyPKZ6IIFFRZXeTbNr8UDke
Wn8TxY3M6sEP6SvihLbVWM7X4MCeqcPXQWjubQtHLs9MzrgplHfI3h8Xc7Tb
9IzR4vgSLGDSA4VvpDe+NXtMk+uApcU6E5NhQk93G8j/EyulZ7eUuN6KrD6Q
AMs42qvglhkoRC4QzYmp/Yzu9ddgsMFCAjc+NrIRRC+FNdxT5HakbgZgOxX4
cTI1LOUatw0bn78h1jPhZCU+flG/fusesOBsKApROvIHgwQDCkmaiGwii23S
x/j3voalOl5hj5mR5BwJfN/b7kIMzkclqG8nMYwAWCKMJWqh7Edi5Bbw+yT4
dYc8j3XwtI6u9qPpvh6xE09x0kNPW7Wy30ICAieM58IL3nNaXAIe/ERrIfZz
riNhufJB/wwkz1eyVEVAqLE2/i/BQSpVEnHoRApzX14xMiDtNJzAPrQ+hSol
mj4to9ndyWsimr1RuEk+CQnjXnYavmqZ8o9nWYY56H+UcwBrpX86iR1cwx4A
aBQ7TmVFhHioSSbU19qzo2m8QYa6cb6U3krM5054tPvlR3GkMtPIeWTrW7gg
DAs+5JbB+pShiH6tK6fFXvghG8DLJnaMBG+QUOxvvtRdNBYqq6/i+j8gtMgy
io+DHfmc8YZyNG5cOsWS06XIVyvR/NRbcO7kQ/EAOhOusymdEo4Y8zY87+Rv
JYRqDMEO4b1sPITxpMbUdUgU4bfqIC3Vjyjsfg7+CKvbViGntqCoBuKM7feh
khrhtFY5+aULUeeqXTkw/Jwdh85vRpe/r3d3fUVSlAyNSQ+xaBf4x5SY3CdE
t+zM7L4+9UYNKTS6muCLeYLk6HW4pc/+gDaVyDAz+qjidBpXw3iCh6p7jjcy
tC9MncygXcKVBJexzAUJv2l2ZND6LG/i5wsWqJncO2L/0j727z4Q3WWHzFgB
Bn2V1m/ScLOv0X41ec+8F6ZHVI3GIyUczB98SaUSitWQkMFHQzGyPIFTJRbg
1rRt6wOgCS8qCr6os8BXdUQdtNmVgldu/d8htOlp8xc3oGlepCHsgkwDWlSU
mvr8CyidRenoM/xkU/aN0iKXGrwZUXxamSChyYCEk2jQioF7oHWMnS5ph24b
laZucB0jkIQUeY3ynLSCBdKprh/qKY+6VQuvi5ezCG8VElxeyCi4/1/P5Bz0
/b3ZJ2XSvsjeDG4XGHLygX0gAoXNVfHJxv5sfcGXVrDitu83XDdob2QH6WC0
j8PSk8yLJ+r2qgRuPsAyzN+hPhHEO3iFG/OxohZRP2WjraE5R0AVBsCRvnF/
D+h3miJV8wrldjYjowc0E2ZCUKZh+TtMNQXi7FUBqq0VMlGF/rQx/08Yb9ey
pq7kGlhI2lF24w10g5E7g3Q2P0/TM/yNiiCaRQnD6BPZgIevQ6hibAXZFDSP
mZQRImSSel+h/X0hcQhpxxK7nbeV9+/q+DwxJOvOyZnobj7vm1AfgviOMs8f
VFZsuJFql0kh008LCArZRlB7n66uw3Vkom5w0V2r06/OHp6v9oTVSHeSC3k2
Z4R8unUlFfODC3S+KlxAkZmI9zEwP5qnL63NI4pbgARPE3Bsmil+Fr6Vog96
qQYBvolT2uAnONSDGSYkgM/iQYfIy7UzmkJB1XkFQHDXRKbYrLbOFhqIFgRQ
SjMQiXW1whaJr9/Ti0KElgaCFCC3Qva7HakIyzAENfODlBEFXOu3uor0hgvl
kmVU+FZfkmvrJuOw7JkJHGZe7fRpE46Ik6LL34908RmiffN090fpmF638WyS
a+3TYnKJelVx1h3tWtduS3C9/tMCtRxZvZzMp5TCW45qOB2hHmV0ou1fWFSA
ku5EwwFMoV84FwOKs2bv8xOTYhIG8hYONze3R/qH/tV0tOHvZclNbOzkXhQG
8VwMqLbGndH6Xv4W4tUSYupwctN9mputJdNc/egqHlPKYdjBdgT5dh0nKrmX
JPUNElgCu5YKMFVqDietbYi5gCvwYRrz8nlXGMQ5tBPMFlW2/vq1HGxBbmZo
Jl/LABDZcBqwSa8ZGavb8Sl6eU2tIfqf5ED5o9j3+Ug5RX5rD9wZeDPhAdgh
whnt+wKShUJ2SpdCpOHP9f2xWIxCKSXZvUwRfl6D+B/TKpCdPTddI0MH4H0a
6wjIUHSJ9VN4rQhOHC5ZpO96js/G6/7zmYhSZy8jrCPpVslYH3UzJITkH7VC
/xKzuQsd6Ufw0uzTaboxxxM3NUqaHUQwv0CgriC6aVBrWJJs4C8kLcBa+nUX
wMvh1LAt48mP8ZZnjOkJumUAoIgWwtWgrP5n73C4OiUuevJaVV8Y3PJe/cIY
MNtGowtoC5kgbb4Ceink9TPFDXeoapHm1tsnmRYNo3k1Mv7YmFNUt1q9Rf/h
A4G09/DjHY+jntrMq0T5aRZ1GaTB9UabXeKw3nvT4Sff4SXKsP8aX8PCSOWY
2vlWpftkA99GPRvThr3x/Y8d6xdqu3YIy7SGwt3EJYg3HnSxFymuzQzQF9wf
DXKol99BRPuY5RyA9mQlzIkk9+WXg79E0Q/7pnSM+WAZvR73MKbp8kVay1J5
UK8B0ioQe4XAE/69vuWRXrfdQGW/yd3M96BPHViwI8lMrIAZ8AkDj9herQQq
NrG1qRBuVNOao1Cnmu9/VxW3fjDvfXQY6Itdydl+VqmqKo0z+yOlJ8I2eTBi
0moQXSkWNQpV4pUzgbIyUQZ4rJg1Oq2ppLYx/O91bGxLxVB4Tmf6i0Wn/YDG
MvqlAM8UWWVU3U8k+rEUVZFwxAzrGAxXhjXW5xeOGvxjzUrHGGgpiDJSvD2F
w00XbpvFe/2ZslilVzSCGAPmYOCqWm3HBMf12JyHvUMX+SvJruriEmFXXqaa
hZHI2Q0tYn2AYpTQoJRpXJ4BhUERd6s/yRM04Kp7oIInrIRhhu2FQAJCCMOf
nrykEevSULjiIpahmzwls0Rco8kGuOZd1B3PInAbYoo2Usthz6rHzMuzE6xM
hQs4TcY9vNjMtUaboEQDHxPgSyNc0LzPr+O1VkXT6utFStzzx8FGkxiEFIr0
DNQktnxlzz8fDibkMndbF+zXGnK7PpO6x7cOw8XdtP+xIcYB/sSOsTG7jCoM
t6mCjlSPbMRTfvxSSDudsdcMnVa87s2qtO53oEAye5W1ASMv3DazYKu4A9oh
VI9qrTf30EvZKAy5SCDIFwMgYPhUr88c2uSvAv9l65+aAfnykFEop8B+wKap
+oKiyw++vJLzLNfr58mk4woD0Jl2jhzAlpzkuVGLrNTjdJmWf13b42iIUS6O
Yhz5Iw8STxHvw7IJQeOh3tAVGEEoq+hntgkLAouPUVAnpIwdzRTqc1kp59cx
l9d7OcnCqI96uFNhs7XOkoxZeLrNe46TohwrZcu5ZiexDVyWObzQqad765kX
igoITwzQhJunOaTXh+jkK+/lv90Mm1Pl5+WCccL6i4SY2AZlZ0C2V1mdmOTQ
JFUAxCwC5RX+IgsQYR7yY3LRxbETrrU9OAhUOoHLASRjnR2VWfT0mbUYl4Di
1Xifm1ihjWfyRcR40WzL3xJdMcX/XrZeLEDXvMIIYueu/5l0RM8kEeqcUoIU
L/yd++uNbrHWJHHBiaK0SUkNkQpIlnOjk7YHVIApQwrsq9tKRC+Drc4m9fkV
pfAWpvfKdFi5/8EQNx5TDzmYzZozkqIf5I3z45t5Gxh9J2PFSWpOEgbb/BcV
7MGLX8DSJFn7YGysvhIBC8Jiye9k3Fc9e5rEJOCyZ+QBolx8U5hoGTV8MplB
V+kfL/CGOhdYgXc3mLiWMUwNh6KjYnK+AuMy79YDpPk+Z0XsTm/kCVeSujpx
NUZKg7h9rkQQBOG0broT9fBQG9jOu+js2Qd6LVTWmL1g1cZWNaAlUrqXMbvs
0iJbupvQPbTzirIUN7nULr9LJPnE2xjWjRiAxxKfqJIDI4bCw1Rbdy7Cw5+0
XdHdb2slRJMDjyn4DYIBhEHbm8TlmO3V67jsrthvstdvjgSCF4TKjmqvfWCZ
mNoE/BkzY1IQwOuULPRenxVrjHJJWDrS7jzJGdRHoi+8cv0VHfgzxM+h+0pF
ddfnyxngnBt2ubDdkVBMxVoZkrRDb6z7XyVzIvRHeRbBULBsXruTPWyOMi4l
9hWV/UthaW2gz8Nh7oEPVCK31RGBt55eoiMkZX4Zozi5IR7a/Pn2/5CdZ1dw
2lL1gk5wEQyzkusZd9VYOgmggQCVpiN+f8+Q4bUjg4quCmjLXF/9oa+Zg/t9
EYrx1aWxnglfXKSwk9YjIzk/HNHNUj18wljYiypQoqgrfkgGcCujYVHE30My
o7Rn3uczt684UetzLt+UOCC8RmIyjdAzhA+jbmoC0LdeogaayajoskHcISPU
vBNFKrnQ5w9PDQvIUvI08Pmy/6jPFHXVKGEN4UwkFfTz9NbynK9Qy4uW0Yo0
RR9FyfEzPPasCNd6BWT3ZJ4E2HCuNiwNoCZzWLsysUNV/WQ0sepo7nZVfFfT
q2O7J29KMkGqVCglgvK569duqyCAeRa5jh2RyEV6uIsXI7FCYuQu5LahE3VT
JWlGUNGEPbA7tNXkiHMVbyCbhmb+LlZKfPWvnGySFAW86yE7XSnKbMG2p/mm
G6Dqwp6X/BdVERynG8y7mIE2gHlQ3tQsTHFeoaW2DbQ5wNsIO7FAdQItPGH7
oDwiLElSdfNKRrvLvRsago+CGj+uMEkBLBtasjgtIFaH1q9bqUhNOb6WDuQG
AKMJGioPRwn1QzZJTZFn1+TlI0qU07tVpFig2NEpFP5ArRPnTaEM9CAO+yXi
n2zv3cmKf8SkHXFtsS4SbbU5rK/H66bnTrozX8vEXhH2dQWrtdVQ0rKEmdR/
CaZMZFR/zqrNmpUKGXw7JXLPRu0Nj99qysK3sFeS3mYUIhQFFOoGr6/psohU
AqeZDhHD8qwFHAYxaEnWlJOL65pZz38JkRHhvPXsvOsLijA4DO0u04QPBRAp
h3219RJWle0fwJbindYE20q27heRjZFm+gZOgi8O8jJmcBPwQ2jAE6m3TUBy
mjpEwWdaQUIYtIir+3UrjjzdWDK8PzmnnI2JO8iImY8tF4A2nG+DZp77dmrH
I3XT/bJq9o4nqYxS4KmGWOWOSBBDNchSFFdfsAVML8UvXzno44tHmNcH2N4Y
d2Yuz2rmC0iZdWAWb7Iwqszqh68QJkf6C0m/HoeOIO98OU9noTeYYBvlG0Z7
ntBuhe38hUTnO4U6ddaS6Gk93Kp+qd+D/HjutZgWOC15C9qzSNs5vB3crEpG
klrrWqMBhypbXzzfnqicvvAmwXD6rhWg1QiZhgW+2UkUvCNV7fnjkqedfYsI
Vl0d9v1HEKeCgB5tNAgSMu/fn8TyUPTMoSIbZvC7xW2ZfiFkmDjJJ25zLgEA
T5lnmbJK2gvOZuBHMaXoNI23Tny7zHUYAcvZoHa/0P+mFQp83ru46aO1iBXF
2+KdBCYMfEmz2afi9kf8ZqAD+Fs2x6fEhu40UqcrKt9v8glLTxhWEG90NIAd
jcsAISownHHQ6hdEnCnVC/Sr7wYif95lIKlLLEI5w5NhlWfP9DTZwiDAvggl
HzNfWssmcGrD72pafbUwUoLpFf75wXFtIwmeOiBEmDfh615Pyf7HOMCQCCb5
l0c3KTdK5AZJCCkvRPBP+mj27+RvvWpAPRKLPFxf0borL7T+44S5lQ83dYz1
19WfnX0GmO1NMGzgERZV1Sg+SxYQaBorgXQV1x6m0K8R1cuk5NMXK8isOWK0
q3b4ukS4IdmEmrLBS4oozjKc1YLtJl1qHdgHdKZYvqwC0GkD+skifSd3UAzX
x7fGZD7fjMHFv8sS/F5TyvK073CCwGoRkGNA9dZ/1Fna+J4bLljKGdTU2zuL
ioWNahmmunwh1WK9doBgCqlC7YK6h8v1FSX/giXPTv3I3tY4Fc72gDlXIdf0
JzXKoAjHpMHTGXcpwyAcyVZ1Or3p1biRC6NbVhJ5BhvE35iKzigYUUVXJHOr
IoEKuWj8wvEKMz+tqwAfyS+Z65uOE4+uo/rHsnNofwriQKC434JHmGPK4BYu
OGr/8y5G8+YIebkXhfNsJOY21OwfKQseSNvRxk1MdMUTQZ9buQqEo5WGqI5s
2COm5SS0J2k6qgvcfPV2TOOQUWE/YM4lJx8R6gy29NT6+pa+/O8u1VOqk0Ml
9mk45EvXsbCRetVK7xvwkXzUFYLeIyM0j3iNZXFppLNuo0QUWY64qlPzcwr9
zFIFurB3djvMc4leGykzF/oS8cw3vmg06n3PlFpoanBj8mf8CB18rLgZP8OK
f9YAaY5u3xU6JRFkpDFXXRzXBXf+OQp5D/A2r9CV6J/7UqDPPKxtSY5veShJ
aiJ4MoBa9VvFh36JmEolFwIY8PLR5QaAIpjKeUP7GD21J36l9PHm42IL1XBF
HglQPeSasvuLP3ko3rqLKYY87vf+v3KaYQzil4mok6N0+LP4qRqFRSQbnGhb
Ucan/cjr6mGLn/5bURy9vp+x3J+fyRvJ4MnIWxwqwUMLqO0i3VvFJ8tbrimb
pyhljgd+pLKyhT2PtQHmIg1lSrgYp0VFrJXPI3TzOBSRbB8FiLIpgvvT5l5C
cXnpao0/YTiEHeJgRIZlLP8/lIY8UOvIrYwwJgoJOMXur8Gqylj4FS+Kluxx
U7jI76hT/5UF3jYATzhAx7o0Qm+wWEdml4CYav5pFs9X84Twt7/h4Qfz5Frh
xohS8W75Mr/6E6uwqeIT7+konvykjtWvaYBeXH07PuIXBi5QidKC8QwQ8b2t
Pm3lJ6ubaNTIxYEYVJdA3IC2DtcUbfc5P2IhKJUEh9/F36wXLSlNnJvPvN3X
zorw/ffB/jevNb3z5uWOu23X9wr3K8+GONuKCWHSc6NbEsJKzFXT+LQgOrOX
PubcvI0wMlrVubbgXDajzeHbPZyPFxmy9emtQVNg0qrArhAjcZYAPP3SStdr
dqgCSzSdk665neGQflzX8ikfRh7+EGYbxF5IOOP8W5mVWSoPJI2uDhfkRmb4
FU0XZSjxdfLXFxxpWsMJFEBjmI7kz6RH+11PLw3yu1pcpB3vHDuhJlO47aF2
oBTDwAP8Ws0XfhI+BCd1610BETcU/lJVoJoE13ixWiyVtH9ZUY3E3ZPHr3bI
PZU5G+YNTWyHKgBqMlR1MAwcxyFZcIH8keyO2MXDQkBpaeSM45WvE+YA/a96
AzXUb2Qy5kVjQCHcfHaSznNHKN2gf/ZaovFANfmnv8Rkw5KBH5pzE/+n3xQU
zv55pKQNMKFHT/C5XosSveZHOHUco9lFWDdtBK0E7ljA2i0nhg8zCf+FigRl
JPJEjY7rR1vvDrtFM7ZRDPlW5QiUPLH7GvN/fcxUGhnC6KkBS55M2nHGhm+q
s6O80vpRa9eB+jPnukcHGkXQd8NW+MPh/86O/JRfDxgfxBbsNSoyZKdmp4JG
8il26mh0YlIWJEQsI/vi+YBnwtSpAFl+LdNOQ+Z2amklfvE3eYTmT6NEFK5u
5g4X76clr2DbaHuRzexX8JpcdX6pU/l+FziW07rM9nPP1rfwkYlSuZwCF1lt
qWnCnn3OmrKCZ7FhPUsY8F2MQyNhHSWM97zOmDUWny0RrBqve7arK3nnQF/4
hO7k14odt+Gdakpg6BdBApDiy98eMdbHGkg0D3UxtQZpTN5etyM+oy3XhZKm
43EuUCbzLcdFznsg3MvDkjhFznwOrzYtXjrnxF/zGfWEcSL7nUIOtMhlCLXK
cJjdcgxdiYbuqulbfSS4tSpah4Xwj2dST9t0abBgE+7S72PnPEIcGxl5OUiC
IrlJ1e7MOo8FVBc2Vs7bk6CMRmhqSsRA0hQKk7EIPxb6YE3mH8tMBsOSeMtu
I06ZElEarqYUVOsyLbPx0L7LIU99vK8A90j9e4dzdiNC3K/gxb8HEcA9mB3w
ky1tr2XbpicysHalBIqvNxGUI59YVMWYgqLVsEDhPr0qmuuiR70p9/OL7iiH
HToi8lFxiXzA+gbyjSBazP6wEtKNw49aqKQfb0jFn086oeo2+LZ3ShVRIOb7
so0g4kTfBGvttH8QimuaNFl/034W0LdcSikwZN2PTU0Pm7yZH8LR94T/yb6A
ewMMnljUUohpen7dXrOl97Sd52l94J/X5i2gSttsiFPSkjgPweeGpZSF7gTp
1KwuUwvN9Atb4wpvcT6cr96VNXTekfBxUSaEHOgvyvXoMSQxeKryl1qMvY8x
TBNWnBp9bU5h3aWCFYl0uYJcEDLH+9nO14iImAg9owNcNiavXuh3s1VYeCvq
OnoY0hHTJWtWoNdvIXcod06FQ0V2431QIsLuidxByh3mX6EzfpGLFyRYdIPQ
+ohdwrC/FfzcOYYtMGiZDPOOuwnIEnpVY6gJx45gZgcmcyp4YFs19jUlFTki
/C63EeXXqg89pSC2znMzXrwmkoSStFJxqknPQ8uF8yWl68QuIetQeLsAUc2X
taRkqQVShHkB/X7ouiLOl30EJeyJ9joQrj4GpGdVPru/2d74m85ES1xfZ2Br
JNohd+xFrEBUYUZzG1FMUz6rpOCU9YuEE98D8LHvnKpS9ClXvFWepwpevlVI
9PEZoMkGJz6qgsU8irwHKm+2mGasWTfkiaExWAfAuK3rNpf0ocwSkrJe4iaA
i4IPTiG/nWgU//yLXSt2Hd0KEKuwAtGtUCDjP3USe7OW7gmDYx+gmIldGOI5
4X8S5Bt7/4Pwh+70Js7cLBj7A7s8goLmXo+/bOsznZ51qi/vEZG/18gCeqRO
gRtdgt9YwEKT7SHVQydwoBdzC+1p7xuMV0gjzzUliGvdYWiKDrwBruWEa0Q+
9WVmpeReUdlol2pTPvGef2XhppyxaoU6OvFhxiDuPFnGlFlRuuWSGENyFplr
sXP2u8fAmHIlb7Tz0uZeVv9NGnrDd2Zhy4TZWAufzbMtHJrKCf2KOTzmbk8S
/i4D8lWrbOvgpBYtrnMUFe1hmNrjES79aIcBdGYPyzkmPnLO4g2O75oRW9by
Xo2ejdRhPo2jxKCCH8fSLiep5vuLLY0wJUOJoFzrvr02qp2RV28mIn8GbUlG
mIgwAiPfmxCFa7O6HzS8ztKcWOTDKZOxkmK3ogLuSHm72++3aXR8nd6YXYMy
Zaj2vTSex630jOknlJxvEsN5O9d6d0jRF+tIXFIyD+KvkpQHOeEIzsqpL5uu
O9GBqdGCkZjP6AJx46WZnu94BsDyhDIzsSrZtziQpYcnpzrK6TGiJqCXsqJJ
1K/2dK0BFzAIkxsVS5+1ENrKLUpe1kUFldwFijXOzh820ekTRqj67FVK8LFR
5bupWbrR+6hmQW7vyFjxMZJN4CLrTh//YpAJae/gsXT6vYhnGesaYO95nCAa
3ssjzTDDvWdIZf8qLa0j5C11kZZqIyIoAleWr+c0p0cCOnxT9LEMLE9KwvPB
Rp1QXyBql+osDYxXVtiff4B4JyYCKiP2xrYnbwVBG6XyskgIi1LoD6cDoszO
oxhgRczljpYAytPXR7Hda/cUEFRHIVjHTUm2uC0iKwgpVkyRsnjvlZJoCVlQ
ayQaK12ZQWEusA4APVasD9IB4BfANeZFhSYF68oIyn+e7nuk8MtKxCxiclvW
T67ex00AOVS/peq+QHZqjPHL8QhYnFIxzMQLSVCAnGcru614JAPQA7QbZ7DO
HAjSFrTTfFq64RXztKDZ8jpQvG9hDLlST57ixVnsgKvYiWdNtmFq0jrnmQdi
NJR9eWgyEpP31EGq1F958Y7v7tRjKjuXHx4OOjvTcWUQkegIxGRfuVTlD7B5
v8TOKCnnEE+7N1OGq9bPD2+SstVgIsVEhbV0M60S/8B/g4zG5+WUZdOoOKbT
H7+WCHMYIqoLtxExxv4zGIwRUH3KqHtFRFDvuoqGHBkg0enASxcN7aBu7Gxr
8gkEhVfKRC/y7tWYJyt956KT06A5c++QlYBxuxn1xOxI20WAWncpyp/v8Smu
LUutqysWjPVxI8phiREoi5qp8ZPM7PFMQsMUU1OzQnKwULXXtyZoEH3FoUQ9
gnpfl6G5HXuQELlNdxtlc1rRJAvUjdTink2Ov4PjidXtBKDcCtE2N0Qa91Fb
oHYW5h+4pfMzjo6Smjlgh1W6keZ5aWv2RHGi7YFgc9sk+M60C2GKa/0sBbMy
rQfx/v8dqic34yxDfjlRVtGhVnWJorkE1lnB9bG5kiqn1azu5SndVoYG9dvb
/M/RxD6t9X/qEX4/e/eiGhmRfxcgDiaWSjUJvHqAz3S5KMsmRkB0AOQFM/51
RPIRK7jxLjYxU8nu0CgXTj1JiJRi03pof/sIfbi3NJmQTcVo/melEDq9XdUu
dlCgyBoO/72CRrlHxIWbzXzexavB6lVWll7zuagcU6wInJ+1HK7zEPqz6cyH
X5P5KHDeQJoSj5NAHQIq6e8sIfLVIhLiK37ZCo7i8IB1UBCDSXjw3IStOegX
g/odl/GBiVFQL96yHv6CGlCilhFuDDtsghKEaMYe6MpjDq/ZFZCSIfn1JIir
MZk2Ow/nNR68qMjh4grbIAKD2CbpC2TvqlLw9jBk6+qjo9I5nhKtJNuLRQqt
md0MYtf1QSyxFNybHAvJp8oC9y8KJayfcyG0VkpqwGKZWIyzPHChHAUhUD62
v3Yn74C5ZfrrHVviSAzgJTwgj8nJpqInCnI5jpoInY0pOlgKDcZhXsIxYF+1
eSYwa9tnH4nLHkHXLxkUdAUZamEYQh8/sZXLkCyUdbXfrtKL0apB2gfjGQwG
HPA0wi2/DrBynEsWrlY8FOTY5tGfxd+iWQBv6BxWBLMNfDo7X4Rh+VBnfwSe
H9hUdIH/irzOgQ54+nJq4wVwBzkZD0TwxPIUkRskDy1Mz1FSL5d3TFMU3CfU
nzaCwnF9vyg4VJyETSFaYkzNEqojz2UOktvkzS5S+V5jDIgZI2oindBc/SzH
/jqO98uja9S/gf26xO2H0PK1dowX5rGZyuWhDBbGHQuSJynsVKhNdZi6dveI
uYDFBtcVPEYvTugOnFNM/v+EzW+VtDzWBfjIRptONC6K7GtMNdK8Nselwtu8
5SuW7RCK2dk13kAFBsyHB+qrub4u0EcnZD+M6tZusLXIF/sfhX0x+jDa9nYb
V6hm8cn5NZ6UefjKHjlqCSfYsiIjFxdtvj0Z4DEt99NKU+wFqBJvdfCPiFqg
zcOLFIPKTwDClVVld3xkMFRoFvnlPIrmbE2PnKjV0QzkzD0uINf9DeF9b/2m
Hl4piiQwpA66wc6p4rM+/zvxL31zCPvhsU1vdlEHETPdhneFdzP8Xs/kLVO6
TI9KdoCPuRLuvslO70laLYkjXnBGUPIkcgfg9a5nvvlFQbJPpc0123xbxzga
mL1jFIfQ02x30nS+BbVLvvj6Nao/2Tf/vT8nsf3+XUxPm8nlHweThk0AhpbL
pfszsSEhOSRL0dJTvsEz8VvCXvqzq2HEw++Rj1ls+RbaKxkmp6NyKuboZKyj
zWJEtNqL8J4YFm2KJKNrztnuwwXcdN+KUIIJhZOG9fPpQXpzotMNYKpcEy5U
WnhpnFQeaFvlE4QVR+DNejSuJLxTJ3uPELdzsv0RTcUlnCWEMHmTkHN19YG/
gEtKoRDb1L0EhZIyCAxtDEYGXG61rCOAH+HPWCb4Xgjb/VPLtjwSIhngkAmg
qYVurJWvjB2cdWIeqpylSUWaSeeWcENoQqyhpC2EbTM85pfnxsTOyPVyguwW
Ja3/thV9K8h3nY0fF0+pAdeInoP/d98jtmVQA89Id4QuidDYYg2rW9TScjBP
2ljVnGw/6sTjPlhdlykbbSyYRJavbUp5HSpGMEJnbuPiF0KJzzC6q3XyqFit
u3IP5O5idHQeRtu3/xg4Tch17DQffyzyFaYYW3qI9mgY8vGRuEEptHMUfOjj
o8ZD+8PKZsum9kk4rBc6R9n74HXPdbspTjyAJoNRqsZzYhX0k2HnYeRYUOiO
yWLhui32P/kta6wIJ3vUvGNrVJoQkUkPlRQGaGcOYgJ0cPNzLZccn2+3DB+D
bxK+qUMfDlhTIM9l5vfVy61FItsS3anDGcBWLyNEryfH6vuwsw1hiEtMEbG5
9q66BQqmEt/sEy4beCIcyS/y5uZBxLkPCitwPIGUh0l7tipLzO5dZyCYWlKk
QSavCaPe/SH9jhIDTwyIgXGe8Xnx3uJWxMenTG5I+Ttlj3eSfmzkmlSM9lZo
N+cO3kHBvGIBinYEXtAq46d2PLVr5FeC+vNJV1gVgRmNGejv29+efJIxO7Gp
Ky8ANfp6jUl6Pt7Z5YEw6bSqWIXZMr0NrgBHBBYKfdE0/dcupy8XtR8UA5Tt
26hTXGW5a3IgYANDA6f4ZpqlfcoyeoUZDk4sA83YE5QAzzOX0Vdj2efx1Ugq
/GWwzOUBRZWLMmG/NOCbXqaa+RoSMBcLa7dsbb2dJj1XFigcx0aZk/iRqO/+
ps+XTzqKCwc0Kr3FXkpr28iy/oTqbWOMCOh0n/KxgaD/JRgqYlsC+ul0DZd3
g1ubWIOw30KQhA5wsdnyv4nQs9LrPAzlg5bBfgqhUYFNdCGtrIeW/M3Ciaw5
aAI99vo5vwtrNk7RWAR1qsmsIAKEVuBDnckcjbVLWRoBtfYbGeKu7eH6d30F
L+QJ4P29gzE8DVK2dRDjo9ATpQhobp/uv36nvLxyVmzrD/lN3MzV5x/dWg/C
/z3i81uws8HL1NQ61wci2XLUcDXCusKXNXLQzeKWHL7fsAvJc17P+Ekhkn37
rsFeKzgSgecrrcIqvkvooKM3OHlHjP3x4yLjSOxfg7aSGtrofiYIinqjIJA/
BsTLxUjsIYg2R+j0xRTyTjGNKx9MHac5YLC1fY6eIXWsVut0DVt7Z1lMkluC
c8zt9DL8hA/rsnkeNGojvhz+L+SyOTlF6GSR+TTPWywKL0xfOzAfklXAaGgu
VIf414kHxKK7X4Q/jTpar90pXlncn4CYn0InN+HO+SHGMnJMpfBB9g7JoP/C
JxuaaqcGg/LFz0w1glKQViTuypvJjg8y6UPXX0aL9urwwzHM01EF2kka8iwe
hcM8UmrYN1Vj2hKPcw/RH7UrGniy3urcZaMY2M338HOUhFgOYdk+UvAbJnPJ
IK8xnUhagEX2dwFLCdYEu1SKw6OKOF8kkQAV3P2XoAXuNZjMgk18KUWQF7ik
7bg0NIwvhWsf91VU4szl8egRmOk/il3FxotPreZBixSG9NU2RqW5I0IpGDg9
AXq0nUirQF7mT58NdOM5LHoxYtM+XadAkvlv/H+pKl/RscQKo6YgDchEWxMP
SAKAzRJ7MQDv2jVkbvDy/8zL5UjKTLxVctUhj7yh9isC8QPk7TRAp2CD4/bn
rq7HNU6lGjoSRrwSWw8WlYIzbNUHisDNKPiaYCwqeQllf+DSbX8I+7v3q6+b
RD0G0XRuRL6QMNScyXlYVfs5YUJ0+gnfOLmn0UFh9SMqauw4v+2YnX02J9Vr
RZvmbkJaeskpMl0Is0exeAy9mdsrPcgiOUjSnIs83oD0/sAW6lZxivRsPOxo
87J/HmE1CxPt8nNrwM+AEWANBJOEt3g3n8zu1gAclKWRklVEypVeqH6RyKOK
2oIFBzVB9r2U3cAPDbnvoujsUZc1JI+7feh8UGueXDCBXMIUKU/uZjmYYyee
lODoAkXXNlAV3XD4QxHHMXUX63icOfK+rMVVf4MXAvoZjt55/ePm2ZWy/Wju
XjrFdLkqcWIAeH0Uel1osg6+4zJyze4SPb8LyH3EXkcJooi/6ErQLPntTkGR
6iSMPfvAiRtdXJT1sZQ3nV2UOUM/NWE+7rZf5i+BtPMprziTMKLMzZgpyUco
d6M0NPFcfaFoz3vYjvuB+FLXWD8dFxKoXMweBcloaa5SqO75l3ftSMvDvvc4
MG8W+4HS6aaKNU9Koxu6F3LeV/o6EjbO+KOquXedWkv2jX1wdPZn6Yp1NmHK
RZxUamr2fp3zyJxe+UdNNihWtjm9QjQRBygksFIn3ssTWf3/rzXEsqNoF+xr
8uyEzNgwl3poI7D3OGobJwEOZgAH8dsD3OZTqhfjGxBLZySDu+Qz2nR/MJ8t
bxVHxCnC/ATCU7AH2VKvRMkdlrEdFc7sCrdLwWtfkfT3M2oAyGmO2UP4cDLb
+wUvuS32eKqflq3SiC61SqEWewXd55OJQY6Vrx0He8vqfamgAO+gG7d6iXvp
TDKWqgmkSpybmk7XlPJ3cH4UHmmFhGxs1Rrj2C0XTLAavHTU532e23mHpAbI
V4I3IISLP6lNKifOMKBVrKxtWFEICIPVSqXDMSNs2sCozQWhBtKa6r8mOFob
tpjU+cjiuYYXWlTLk4G55q4VL8Xo/8vGCqt1/JoTc8/Cq+HO73XsCcbtTn+N
OsdHxVixdk6MWT9tbWDHtUYWucrVH/9ddSksQor1DicwU3O0Fw+9Y5zmFpMM
XUD7KRmRm8gjQvt31YjEXqxhAfkIYQH1Z7k3NBGyefPkX6vk72LnB5F0qio2
Wqjv5Z8Z0EWlwXAyqDfCNdZ9wgRNFIfygG9ajKu1FaBDvEpH+ZXXYL6pTM/6
5UZ21ewCNAmy96RdiX3UMQ9bgQzAjshtMiURwNvVML9hTfH933vZsyUQFWqs
ef5RLFVzcakBdSIhhc9MOz7LOZOo20F9KDJoWbKw5YHo4yJTPmlmr66QrDoQ
XeQm2JIMx53/xM2EjIz7tltj6A6Nn39+SrQs4K82p+i6oYWiLsF+wL3MZAhR
9/+VeHguEynaceb74wOcc4uMjP615KrC0+0AsNgSHi1uePObsOX5gV5uO6a9
Vn1rJstU8ByowDM9g22ArG84KWo7BkIWn1I+9KZywWrYeplqvejQ6pIfRs4Q
ik8h53uJYatILYd1Y4WR7d5K1uq20ZOmNbL+I3qIhqNW/IcUCb41QwR6tqJN
ut3BDEOv3WXQ/z+nmlX+lchb/h0iQYVnCLkpyxm88RrMR30Ad6DQv/g2Ws1i
Pvr4mqQl0yySjDnbBlNIMFcvHNX/iGm5MupMW8YTCRm5jboW2NEjDcT913V7
rmcJMvtHepnfVJW4kW0jZDK9W49PBtM5rYL+JENg8uRj14Y/cuMSAc9V8ckf
Ud2pjwMiALd9Epu+pueipOEahzaMXTwuaTM36lq2sg7yzL61SfD3VOb8SRpN
FSkUfcY9PU3O4NkwZkYdqyIah2EKLkAHXiN6wO8k1adH+vVV2iJwrJrgOAiK
AwSE62c+X8Km95ab1lZ8S3LzZyAnyk/yFxlEqKEQd1Hm82EX14rrqkcbzQx6
dYOFRhQJcMvePJd/zf4Z2MK2mxr4+JXFcw/UlWsPtCQCEUkH/nueBqzX5H3u
CKGjN+1JQjdsBOh8vDb2deofsY44r5nqClhzMgVQqXtswsga8mbjJo2JIWBM
l43DdKTqdXP9I+bz0dg22RaZqyNB//QGA6DHffL3o2ybHAjnfiWCeLLD94xW
0g+XT19kEMgjiAiov5tE1DJ1xrGTd6YFKCBD2BLt8QNe80G4SNWhUOASvVEm
hiRkaucvU0nTM+AYt3/D4OtZ7hUM/PY3f9F7RbzNKjgFD943s8rJNv2TC2CM
RC9Y0YChEbyhLct/ZlnVR+KKQYtCz2n0AodX0hqTZYLdAGjnS+pYVvWz5STw
syQxW+Jr+mpyw7abw+Om7m+IJDc2WFJynjoxrDm1pan3yI9uhnfHXNOMG2Ln
J9HLsk7fXm5sUi2JJIgybHnOIp7dd6V9O5VlvRDIqnH8bYvsz7eFGCBAxybF
ChmewKulb0t4iwXsMptuuEe4sDLMD2AiZYFBbKH+8xbYx1aW8QIiC9bGgN7b
9ANG/bmpwgSgu2FU9DdRJYvRNzv/TppW26RAbvZLxo2ErO1jIBrlUVG+a5ZK
CLFTvitd7mEPOlzMWcTiKJwU5l9P1f6GiAIlpyC2WyZu5KNvCrhhmVs2Rydd
p+Ya50jiLUd+JNODlWw/vYAupDxxIKRXEBYyi/OwSzfYW8eipT2MMjE6AanL
s0YcXbpUC1PhS45UiLGcwMBqw+PH8fjIyDGK1WymOX8CND3CZVndWvLWaVAX
/cCUKXnBW/YnI1Rxgs8T3QhCfu5CEAcPlXAEAtWJx1hoX1gTBeReh+UDZG5M
jfg7Kkyk1Uaqme9lfzfSTFCx66E8NFz2AM0wUbuxoOe8oI7FQPsEF5k1dQtm
aLMOScBaE2/xgqxy1os2c+TM9qi/4z0oV4TxtgShWq+XMPAzma9uZoEcKTni
kNVTNQ1cQbgzNyczCEGM1HEMbxfc4pSnFfi/Po7bMMPjXuL0F7j0rYa6M3mF
xtAzW7qf4ta3KJbzvteyjk35cZmwpTTg+NhY7vUXHZmH08TCYT+csW+rSxQQ
NhK07KX4KL1nXuwTPtjj/r/hqjXbSXJUg5GL2HV3IcPyLCDoAGFrAEA2NKvm
sPEuBBamAotNTs3Qe0ao/gzkMUJS3dxhTBRQOqx2nwqi2WoyRO3KhKMcEUXj
5tt2OMtv7BDQ4ES8gKiQOHroeMjTxD5hx8Ldril/+Cy47FS9o6reuYhVNlUi
hTV5+zpMJmrfySYLxQbMXkEUyTc+CCfY4nUcfD7ivrZGrN9kVk+xOdt/vmHT
a78d4eKFhDFBL4hsnjoW7lWPII8qPP/g3dIKdfz0yxsJyK1CpLLD0G7plMLG
guKOHttQxuo94evgZdcTfniBoci8MdH/t3WJLaCGmHBG3ymtsK1cXcJnZ4lF
3GHkf+BON4ngJ1/7TpD/jHVjsmH44riitu8hx/GMoZTmNVGGOmRvfTdH7mhL
Dtct1vmeLrtEu0zko8mgTnOOKDC9i028ZFL274E7eQZdjBn+zaYD5kRKUiut
PbecPiasLRXBru9/mw1PCeSelZ1O4Hva9YLjNdPxLh9FFH0K/LSxDpKPyTW3
20Hy7O79FZ2iVX5VCo1W6/DRY+ll3GKGKfkv5rBmAFGYm3z3oBKTrh3oVs9T
Xvg+vtjS5zudV+MbXmtlHge2kUV9wsSw79+wr0sLGYG9mUjBm8fpzcAMxQDb
vEJ5bs7zZxKQKhuXiGSLvefAV6Bo3MfMZ/wiAPEemCR8kBfbmAjloV5rjDuA
WFMO/OG+2kM9bqyKx7xRMMDyRB6KxAd7lczvfxsplIWByL68jaJCSdJH7H20
URepruXg0BeI/rXkgWA6awQGyKbS9PJ3v8PykyW9hV0z4v3+xSm1nVbZcEKT
uknmmWE9eKAVdtJgzSCJ0eVBC0tOL2zuyGAUMpj9YjIl69XCzSvMIG3UYUA0
+TKdR7K+NBu7+klrajaOTLy07cy1czddNyL3N9qBBfdl864iZkDu/2xX+t1k
nhp6KY3CFH8MtA4ni1Vk3D3FNp4UEnv2dsFWa+jHW8qFalYeQ6Uw4oUT+E3p
ZoBWHsebI5TqHZq8+5ljeORwOQtAV4BjG3nCzZ6dzbUCf0nrXATjo0cysARE
Ekvx+dWb8YzK/NhGXBa+zoKdY/CfhXQEMxtuncj3fvMCB9Ax8j2s3ZyalFsv
PaOjsIV6LcIhMhWyeHVDE3femgEegM/jsvalLsBI4pjzRRpRIUgeF5pgvBss
QkAajS4HtMB8YAL8m0qNZvGtu3Fd0T2Oo+ZTRuMO/JUFU8DMQjj1cw5yfy3D
SOXhMoVPqWDx4U7zjva/Po/Dq0iCdTHWFjn255DzH9zbCsMr+yhBZELCW5eJ
PgmxGtOoKCb54fQ8lYENj9lzq6ZoI33NQQUarvxlEis4R/YMoonCC3IjFpU3
BoNZNOVThapwy1p5Y3mbcJK2Rh+OGFJfg0EwQn3I2KBo3pp3uXJOIs0ywGK6
rCdv+e6hxIIbzP4qq05ebUOn9E3fGtLqTp+Qmn0tPe7ZoGOGwrBK0JxdRVv/
07b+qSqBjws/ErcoM7zqs1vUbZEQQeIRIfSV6Mt/g5bAuv/YH2Oqv2hi06f7
+CzPBmMETPHz3+coXQegYBRbzEMyh4tkOo5VHYxKl/Vb+lQ4B+ZYzEkj8jo0
OWoMiQRbxKxpRVo/Gwi6bupXyXNSS+SspqMlf+l2+He7onVKo9upGIMZQlOL
dmPJple9Hu4muJKPSJDzPV57oVMwMC7SLDzFMimqPuzkEd55F3z8ngwUuJk1
S4ryH+sx30H/mF1YrKZcBNamqecnfdzDtRKkgxoVCkqxvF18D3L/4vFIo7Qq
l/IGUnHamomkwlCXeNTY/HOru4M3C6HAwfNFz2pcCf8pkTzc+WLLrHFK9VCF
t4Hg6mIZhcFDQCkN3//Rk0Uk1szAtsIaRGUhAWm3Ax/aJ7Fs33OwsqTUVK9K
JxlxWosJzlUzluy3loJAFYojudAO9/WfbedseYS+9hXjJGz0BJOzn9eyufmz
BVj7rXbst5Hzd3lhn+jUM+h/ZRh3NjUKbJZXeB0pf2ja98hOTC+ebnAe/7iA
dRGxFKvIheReyZIojlr1lpBuaYqkngw0KZt8s4sQiywz3eubwKDgdjRgsApN
rvDahRGjDpiAXIfKFU3nNBoHYyVwenzhXDsy+mulYq3q7bHyPEhfAhIWQoL5
a/mU1lp/M2O12pkYFYs5jj1J1t8LLRw3JBJwQlvE8RVL0jlm+vsl5ZLW/Ek+
ZBrgkdFXmCmjR+g2LP6zH4Zs9lG5STVfgyeaaYLx12Ela6g16FBSieiTFCqB
J/r88LbZFWI1b1KJWYOg7qukQdPUdKdIoFyr0vrY40FXYOGVuwQz0KEPU3c1
Fgs+QxmGZ1jdRw2DflIn+JnZIbuBkwqC049TUNBvebm3NoqXCQqaRqQ4Ej2l
R4voux9JGy6Vu+gTGR2BwXQCRbHa9fA1SzIAE+fbbA+ZYI9FuEh3eJtb1UKK
mtkzfMkxgWXfjJ8pQw/VMrfvzGOaxwq3f81B/u6s2y5HXcVzAe4BJX/Ny71Y
mTdF/jVmAgPs43agbMVWnM/6caZY52KR9Q/5+smrCp+HjINqGfNgAPPOOoSw
ogsn/wKl3FmVEtUXDRF93PiyRq56ApM+r0OLnlMmz+Ee2o/ofd7Uka+uL45Y
HwA/2pUcNzFI1hHqgcXXdHdIbN68iMKBEp8TXJsF8vgacrPc/HNwNRsOfmpM
UUmWoIjJHavMsRJqF8kZYB0bPFfUBt0Vrnici5/ehlj9EcQDGYCyoFnZak01
ZOgSeskgvIjr3+JKLhLCnX7nhai+/CvgLbO6DvgX3eeIlcbjZVxUcWmJa8Ng
wVT0WfcAntkRwdOx85sRdCsW1zH31EYRn7gLp9i/3kVOayse9fjL1I6D4/om
bQVztJTGSreDxtzgK9b59DFENu0pbVgMZAPPbmiHR+RBkc7PZHLhX0vvtMfX
5bzJU1Uz57xrqzRPYAmaNkGVAQwO1EWcp9gFuNWcNty5ALFZapNY4GzJhMcw
5b0TWBf7PRoLEGNCBIJD6mk+6dlf7fNYGM1mGOfxi4jyAOI5bSOJ2syoE9+4
qCnBg3dQ/Q8kF7w5i5pvwTNwSEWqHSJ8gscEZqEmEg76SsRDUxNE+Grbq24o
SjAnRXtZR9bbod8lU8YVDltUFKSPvWYoeM++UO1x1NMb5+GGZTugwO6XZ2Ng
7iakone8HY/O5SbIWGLJjN7UCHYzWwdw8BYUwRi6Vb8omp91n+tpzuSMx4RY
UhjGwge9nPyFi6Gux3tr9In9xwN21N/i3rSdrAd4dhLQv4okOyyiIaFU3wRM
zJJuysDozYhnrK71lAvojdH3cyj89PQy++G2T1wDTtnmBeR3Ap1fSrX4w8Iw
XxyekOkAlnyBZvMHmAn/2K2aOkqynsh9RVpzX7Kr161K1Ht1FThPEzay3OpJ
QQExR18LOlGagsRkQITwHdniJ8ssKFw4nHHKzgTaTAIKItLTyu9ZUjdU8K3s
v/ZppkQy1b9fLrOkUYa2LgDTnGQ2vGbpOVhpV9jP3BpoiX2lOrZpWLtZci7W
ZpsZJ9HT3/AGRMJf/52L/fUsu3yCaSE8k/pH1w5cBYGUiVkj1xPeJirhLzpE
sB+BFfd4B5f/sw1JFuIztm37RB7SV/PLiHxYZgHxOizAc1Uam86MMNYBXAIp
9XQqESore3Fs0FzJ3rC4AdhC8n0WRcbl6vA5c/Q9jaLbrjDyHr3BJvg4O+eP
f1YWteauqhT4BaNWFzxJ3sw7GXzeu/W1vpb6d/FVuyvUss4F949BdvgOWWcX
CZwzenRMsN//92TNB0nIt62c4llyX5kb0uTqXAD+YmFsn/Cs8i4Ibp/lf/1e
Y8mABtiwuhVoW0uLyj8w7mHConTkpWzA9d7INNnrxlRe4KpDSM9DsFaBCQ6e
3VASSpQqsrZNdOdxckgqZUyXkqWP51G5UhE5/5BpseFd//YyFEFnGy2HzmLS
BFebe8bEqwcZAtTEuw34lPJqVDy8uktIbEAmm+EfS0AsJYRq3I1p+26cXwLH
dYmCGtdJNi8UGT7mUKze0DaJ7BpXtBuPb/WciQF10dB2dj3uaoC0HQNxiyQ1
o2zgbi2vFpfu5ZfBiJcoARv8gYujsv1BudRouPIqi3EWjKkLzJGk+PS2jB46
/0ZOmrML4ybQuOElHol0iQqxaMYvHvb8my/ea/P6Ng6Che2gcxFLFJr9Trn8
8BzrQ2Cy3x8AT/oXOc8yxS8dBkJfEgtP2/n20M8QlOQ5N3sF0cF8lS666Jqh
p6sILAqHlvUm2RNLIKlHORW+g/f+H01n/XjVugc9Zpv1YZY9A6iXRjvjRJ+z
U3dLLPPHUB0zJDvjum8SYBpkboSTbds2+eLJTP6CkaBGsGoWLounV+ZnI2NH
NdzyR2eIL81V1hpeQ3s/iauf2aEBYp8XyCmMFaYv6Hwfa3EoljXKeAtLJpAc
c5Q88yFK8pts/wn83wsQMe2LMkDpar1AZD+GCNgtk2RZTs8XI41mJ6XYMulL
JSJkxYypxIWKI6eM9wrNe8NijXUrus72da/yMC0aCBIaQ4Vb0MPaSSpBXY7u
z6pDGqHXd4EkxXuZzVKh+3Xp7uKoqo5qlaL2tDSzm8/BqoEpE8pXj3ReXz6Q
tDYKsWeUAsY8kPm+eqvL4ahY5xRO4FVHKMjD7YoBdq/JItC0LBgXUqbLpygO
UrmUxHRXrJ0Ubv3WsXQE66tT4eIgXI1DwfaEt8w7NeA0c2Px4fJ00NKcBm7B
xhjvlJMnpJQXxxGJam2PwfQ+tv7+eO0KfJHgVhaZuWSFl51Uaip545ueFosY
9iX3IjQs/QGfp0+PO70kZNSAomxdFAXKr3ilNxRDn65BYagGMt1yW46nwP/8
3aiPlrau1BfaUf/YFkWFk2wLAJf9By7u1yFxV+/UzpYUEYpq8/owelztPuVf
dyeXI8PgP9n1LYP+7thFjPJLVQLNEMTZHjvcwXt7uGUKbxjsnzQcHvtZUdxV
S8DAhp0MXG0ovuXXieEGEEnNTi204J9fzE5MwY+X9Du/r3IonIc+bP3Px1No
3hUBp8Q3LL2rWvcvopDCktHxuGDC15OYW+9cgTEjbitMVIIi1Uq4tONwRGGp
oRZvPNK2EJbqmfVgD78t6Bzq6tqBglRYzNF3d6WjwUFPQzgUQ3bmcrn4UPyS
FG7QDGD3X1kSvrm88qsJQ4KhXbeo1B6d7GZUzoocuvT1YOA45k2cXIHBzBUb
sCQHCtqiNpcQbDsVZ6uNZfxUIGSdmJfgmc/CbwjCppT+mTpv9O8A2scDuIpz
zneg2v9Mz8RLBDUuCC6i455kYz4H7hJ7p0Yv0S2GPMDr9h45O6PC7tz9dkEj
KbPqZSr6teSr4InqRYsANTD54bgCaGMOQoljUjQDp/tkoVrxvhXKQDYFTDsf
dWo5JhqS6BC4CEYjDA5TFGe5O0X9TRSMWv8EC6rSqCXWwdLg0Y0/qo1Y/3nS
eD26k09RcsNJohHXYLbT8mMJ5yymWd1IVvMUZ3YbTWP/QQ5xKHJyjr5MYz0b
u6/sdmCR381IioO8SW+dAIjWpQUcY5TXGsLJvRrUVlAM88ikHXpO69uNR/yS
fZNmwmct2HKht+ai/BiU50kGNKPal3+KJAThYWFNswtL+GXq4isHvW5oUCSX
ViC2lgxJZIwSWXww5z639kkkRNg7vO0+SiBxP5nQB/YJE/6QEAIMtOyYW2Lv
33+p1f4v7iiw21KQAUdeb16N1W4bwb+HGUswQsMu42CaOFKvzVTiejzmQda3
1O1l5Ws/Wg382Z16ZH9Y3NSN7l0UNYTQcFyrDM1S+xrrKyaqxZF9mf6/Bf5+
ErWRPXuyes7+ZznYmsesSN/hv4+x8oK24JgGqd7k6kCUK/GBEwrZV91308dY
ADdU+Wxp37GvAr6nwIQ5CK9vi7ZBGev31UaiF7/BV/5zwnRn2Y1JTULq4a1/
MtUeegGV7T17tYCST9K5TKtVskPnqho8v9fSxTQPxT35ZrurklgYfgucVs0A
rYa8sgpQnPkHir7c0hFNu88/12trVSq3WkCnlw1fo+Skt0Zg3gmiN0pykpHe
U0EBTkJk9FBOYwhsXaGhacOigxAq2lMdhmKULapXGSi7SW3IrNdjTJdsAmlp
CMiFpGhd9wcFOR/BEQZMMi4b2rM1w0IsTt8VVeZf+IQzyuP9tVa8KRV715rP
3cMLVWecli7U8xxUzPsPJFNaeOfNs+R98CMFyftuTboGt2YzlXJQnegU8h+z
m1cTj6HT4AkicGYZtR///JWZtdF0+LmlVSUI4r5md8H/yXtIRHKizhR1UAaq
As5tNpUMg3Ij4+4saIDMY8psu8HwkHHPrBHxZUP2WQL3ezRQpIpQ4pgU4qXI
/anfZPUtD6JzAThn9labnXizzLU/FDoJArifGx4hJiigtaxzyMIEqn1Fd5VR
XicRvCnl4QqnNM2dBavepauKp9Jc213EWcttnJQDVSt2nRg8/bFtzCzzQGj7
YLVVaSN2P93tHOAWUtXe9kL0hsw6/txJq/6NPkZpVxA5JyHA203Ozuve9C4G
RhZ8yvrBydBJBDyqcgItESCeOcXFKlcCV/MmOKhIYyDvQWSsdKkn7vC/vgf/
9ZzcryzVmI3u1JNarJmWL5NDj1w48nVZf3G4UKLfkbMPFM8Sy8JFdphbgRmA
jEuWdK7efDYXOcMn5bNQjiy9D6smq+aybjyhWhP4vemG67t9Vt/eagwDnIZp
Hk2za9kL0CR6+GjcXw7hoIg9UvEvJfVDy+yo/r9gQ9/gKxR/Cc9GnPxk5NoE
nydc2B4qixLrN6MMSYvdYx33iyf9lT+ahkbhGPcb3Rz5bMQgmJxijQ3BBlLf
J2EsAeKk4KcD6pzMoW/yp6tIMnjr3ZTZXG6uiBPzfIF6Lnr4wgdKRsO8h03M
4klQ/UAAzvuGN0VOIwHycuuVX6Q1pnHOZRqmZjH9tpEvYY+BVQ0sjaxVR2FJ
yfSh5D3vnBN+vxOWMVfypnc/2Y8WZQqVolxEsT8leMfJlKQpXfKsvSwERFHc
pObSkki0QUZpuXSQMTlxX/a7ZslVZGrzOk2KJxdATuNZsTnJ4PY9V+DFXitf
ziqnL5ytBZcR08gXVMkIfoI8FmwEzydt/kR3mkv1Viyt5UOeEsfl3dbN6Z5o
R+QCwst7CQCOXC9JYksi3ev0Hddy9YddrBlnWcKUIMZDPvir6L7Jo3+L5Ast
uDvOfvksfU0Wa5RJoSyC8JZqranNa400PI7qqzgI4yxJKqUCBKoJG15elBmx
WSCAIpMLMq11U4MTS7+AuFrKHsh9tgy3uZ9KIjiw1/BllwMSlxpqpJgZFh+7
oaetJHwBn7mc3aiGmPo84exFeC595zt0AApaei8tamDA36gsfPWYbfHK7J3e
eCzXtnurzcjdfC1rsIXgKEdOAqxg8rvJWnz8BajZjKmi1MlDUwgilEMB55Se
bIbKsz9vhNOW7nsjiWf8VKDWnQIjW2KQnSYy6jUTPDewv+Y00bNvDZQRGcO5
0i49ehMCylS8Mwk7IDiNQyml4ar+2Btn3coNHl0c0bSE1GeCwgKuvcFmdLgu
asDsaCWBDrsGKIbWQWfG3e99Rin648P6FqcAqN5JShG4TlnohKxM6ewrUGI4
dZpAGjmjxVX9ZqiZt7nDZmpo2nySHZb6aQLxTEj/FAvRfjoVaeYkvHFKW6OY
JFWTWk/FoVqYfrbJj9xKU05Y4FpfyBEXoYNrkesKMnWyeGMw6n5fCeyAme3m
IP1yGYK1iK8nDtWY9uUSrlhL0l527MosUN97psVvOamEVLmN9NZ2cpYRoq7Z
WWbW5kTYeFRmX4kORNIBCDBMR946nk/8DAhH78eBu3+YHlOdJw4aasQDeIpI
jLD+ankYQJ470GAwV7nBbPFtTxsYWLbhHjVvl9wx6pAc2DuNi+VtFD2rXbD9
BelW5gxeiGlTXmuLUfDX1tTqY9sBf89wL3fJJhwzm/oEYJbf3H1yjWj9jJbo
U1bp9CgUDQDyirw9J3DpU17SY372dnWh8CetlGSkeTGjUCB30wt2CY4Pk7Ux
3/VGs6g+cONNrJlLILLLor5dinGT2aT6ftFccnB3jJmZaeCCc4VGPI+jYicq
/VRYmVEmrb+krjpevmnSbNcvgyVoEarCnQfpphhwUieSomL3KzLj77Gwvyh6
I5nb2iYCGFNgsoSs+hZrF5ctCl5pOnuUenu1dXlMZBJ0RKi4CXTsGSFJZ4Cw
IzbPVj/xXITnFhxV2+Tp/r6+0vaITLPvQf3B/Qj0ZZ9nOICfgZ6w+2R2uI51
NDou9ZP6bkOVVumI2V9Lbbp9+HJ720BaElBq69NdAK7oNiFiSHdIFokoYeRd
+LSoydaUk85V8N2Cff9cWBimkHUVLsqU869WkbYCedTYqBTWpwqbkdMEuF68
D5JDBRKN7WtZ5tUu8mbwujhDbQl6E5/dJ6hH1l/oqGzvdkMxK8eZT7hWbn0C
x7SxMi7LK5p9uYyfrp09BeGb1yKrolMEj5YJ6ZtfQu/CiOJyPqEwaAesyQdv
Z9hL2jDPXF/vJ3jPIQvlLG0D+y7ou3WcnQ8xCwpiU0kKzi6DuAy9jLWYPQ/P
/3oTkeaYaG2dINiRaFgjt/icQFE0s5nHgcUx6HFIXy1ICivUIDarGk1vHGyW
C7newOmvPuV1an9WmgHTGyxuaka6UtR1tv9dKD3Q2YeaIHvGuljJLz0rYJkp
7QgPhY1sZRH9GGunU3GNEjabg5tMjrfOXp58v0pdEjtGsrwfBuuRjpUz4dg9
xlIx2fI3X687vcABiSxGQxKmwj1XiZ0Luwu+bO2voDtGIpKKpSagxw4HQHTJ
puoJbXhcfpDpE7N9uqOV0oSjUqxd0mJi8VyDUa4lYhV/Cl3C8VWd93H+RJKD
+R4OjwM5XuJYW36s/Z9zA109VkkkvgWOvg3bKBKF06NWwlkfw3gitNHzwA1O
FidUdcpTPGCcxcpF7I7jyGE9FwVwkp5N3J6EHeoOgX2ZP61OmvrTtcYrh4gy
4YnYoFrH47NGMqF6D6QOCaPIDXEhIKUq3ZRGzx9cbiD5nwMZZTFrKdJz47S8
r1cf4w5fu+YNKydY0YcuMb5034uYq4vNUJJkfgnKMDCx2Zt53lYqRV0wQbob
JJTDNC+Znq1Jr28isQVTXs+0LY8bcFRpmgW603XRaxZ2MifA9p8EglyishfI
3p/cMhJnlvGhcLAi6+A2Tq0M9mb86fKmDO+EJLKgYjhCuuiOR6MRBIrWghgh
b5mSlUTWehSq/5OrDDgXuEvDSvo8v61bKy9iUfx2urWcvFY/uwvvkCuW+YUn
AQw0Ucwb9O0kw87Q9Y9MfXK3oan2zv36RgRPYL6RdDgLzx4ZHaRN2ekllAy5
h2cbqIWsPve2cJO1AMs1uY5Xgp8AeFr3IZIzF46SMwx4bKVUx2ui5GcZbAWM
Plal8oHRbPZS0+DoW+g55IUEy7KD+pUdQt0Htl6CRqYi5bXbXElNBfQYcJnV
oF+Zf/XTGp8kndIBvjY7BeEE68mZyo/eNJrZRuu6/5h4LB9eESFSC2yR7Paf
sFgPHdNMe/bA4rTsL1bRe5x/A6kM2LDIWvKOWT7lReG4wzBvPQuVG0YQ5dek
mVoVPhUpFnVBlnNEqrxhQYIm8coMmgI5IHhzcDmvd3IOE4DvJUvGEJiFcdHf
bwtLAj3JGRw4A2yrzDzrUwZt964zmaEu+CUOX3xh62ueDIIMcre6M4fkJobq
L5BXxd000Q3fhE1PHQpbn1O4zYeETFrCu5wY/aktvR7CidxOuO3Ny1PeFaSD
RntbhyDKzgpa/OiXrJ/qaMV2gbhoFmtkpTnWx4trqQ4kgLyfBZDGG6UQwpn3
WM9FopswbB/DqHol4jF/nvi7aAgs4lZ63/+ann1OK9Sam6x5yLcGM4b99jnY
M3f90HW6Q+o2Usu7BPAoqcJ+ah7ATpEdVayIzOe9TXLGxfdva8LvANwKtaYy
9o8Lng8Hq3qBzOSChIgPC7gq+lefmsfWPUJr9RFehf4AMIqLJiLTfFQo3A4c
NFPj2aR6i+oioU2MBZYJ5+cowFjGyfsWMcPpNAB4+gBRiRSaI+9JHXBS51y/
iAkLr3uRVTNjJQsQ4e6hDOsQsQGwsYxc13eJJZZF1ZREeaqUkfUSN827y5KS
yTtG55nfpu/T2DnCV5l2ctN6FPdKClYxiNBrfwjIm+arufX5qm5IN6UI3pzD
/LCV6Ya9G595DHXcnVDqWvKJ0S4OSMNPU5/S1+bVBlE52Hs1yQJa2Bkw7GDx
Hgy7B4Ormu2f3RKqB1H9Xz2CAwQYRYttgkkBu8OUeL6EGGocvIat9jHTtbDr
wVaHaIb3/udFz1h7TT+1aY4r6UfFU+97WSn7YGtkASa6CBGi6JvbkSv75lop
Ta/2OK7e4iSCUz2xkytIohXxuHp+/QpgRpE3Ra9YmH1g2j4ayhoNW5oqEiNF
PitoWsZhy57/NUnIzyO7V0ThNAWNdrV71P+s31RNmeNJ1JQ8wcgcn2cWnlia
S6IAjk8/z4/FHXTlKRzuy1XYjKzWtd3Lv6cYif82z6sdQXmG5EbEOQhjU4JS
vnhkN76yjwBzuFterVBj+Imf5u+Udcl6RUHXeZ4RmIzQY7PFARvaQNlLvVdl
V6msW2uZNlDQnC9gwWz7g97F/q5CorgnrcvqEXVMf6Z9V42jJDHjthHTnBS6
5oj3TpqxwGovmkUk5oi1BcaP9B2OMURgiDYoySbC18mCh4v6K99PUE0VXfqv
ACLlkhrXiQmVF55LognRZo31NbZy7Y8OMGU8m8DZeQyv0Fs8UeRQKJtfTldk
ptvXE5+75F27SQEb8dxRCeYvJ6e96AG0iyfP5YbeUvNsZ/o0LOP7vOo4v25S
W8bCiDSFsauJjgsrQ1iaqb/mC9YoyNnTtMiDJMQr6KURlwXayt/+o7g4CkRr
02H++iXFuYwilOHw6mOlZm0JzFvYisIzsCQabuPwbpNyzmV7idgo1s1jWIhM
Dk4Xs+h0pl46rhOD4Id2zLGyedGHIz/RtaUyOROWB+ekQ6fNaEzl/13LTUAi
xABrXaDE9cVwHYbAkWEt+XBFknGp2Bs3uniHJdbpgkaIw2+eseGsvyhIAr3b
oZtulIhpfcIAnc5u/ZxJEZj58i+reK09G0s4SzLjQNOS8KOPqB/7JKUm7Ctk
oERdSPO3ZdFmjP0XQrgIh7RlyWx8KgmSCl1n8XMIRr2QbBjYltFOErjC/OMK
LKNxjzehJjy3OpgQu0rPpM/rHw1Q6TFW31dZlUuVX0rqo2fj91jsYMs6FmXo
EJ9WGw7JfchgvWkGN0aJwgzfav1c5lHeMmFwasD9e1UwgL56VqCJpoAI1l9L
tQfiGTijTVHP9OrsyCDnZVQKdveVJHUYoK9HRVpxmeqQZccScijwxAIXEaZ0
7jl9nU3ELtzM1XLPm9Zksyx44pOV61ovmeFwDUwRZVQZ5zK0b4ImUqainKZC
uUyU4rUYFgTfPAQEiZ8hbp99jaoiSt1H6ZgLVkPp9Xz5ooACiSchX3Vt6e7M
SiN9MUnG4LTtx6fei4y+AVV07dJFPKIWGE2zjdrodi8a3JIJwPE3beQ3yIOi
9Jkj4QPEqktVnwZQRdYJwa9mVfgIpVznLoM/Qykt578LrcGbx7mGoFrbk7dX
RONMSO3NEGoIE62N8QgMKQO14g6Xw8s2YsE7NhY91CfnL6AFt9cbi3RQTzEx
Hr7Z8qS++FN6MLeKm5//FQQZA8exoYO0+fnkh014WVEH6J/K0+MF+pQaQgxw
2BFs89dJrXaeJJTeRe+tJVeJ94MnaVBpciGqF3QCs1uIebv4B0/ooiPqQC0O
TXEHZTk8VWb2hYoJ4DpB8dVwindQNC9Kqh9+oIgo23lQsa7dY5h6D+Eg/dd4
2Mz5Yyr9SHy6mme5j+pwCx6TqHK2cYwZ7Hy4tFNw/CYZbJ07YLSeIJnvb0ZJ
hUCElKLb1L1goOTPaW47BRbbk57nJ8bNZnl3eHaHcm7bWEWJ09ZWLTrek7j9
lgiDyNDotafN7KFeYkpokwMNfQwO+JAgk34PlevXCW2h9xbbX7ho/o3NNBj8
1oXbMSGGsPHr2vrWgCjf4yR6tCRGW5il4bOy/ribgUVm3krVUOqf2x/cw3UK
pRN6mx4TuSLldaDW6yIaY2cp8Pi7PmOaZ6wOay7NQw9RKbrDG6eZcqani1Kb
TzpMhOxLlY5K6HkJ3/wvVCDC8ULZEaDlEi6XiYVs6jeMp+la/hLGbfZ7uf6R
mUu9TABZH9CxF2UOY9AEfVKM8jH3soYD6ph2HdD4B2+En/2S0VcU5QHh+Mal
KoXC6bqL9HFpDbZoDosh4g8iZqzukVfY0IWVUSQk29oQ2nffeBRBD91WdODc
yJsDC4umpo7KICUgICr19A65jwwaMGHWyg3LIHUhhnZsxg7t3O0GqMoMCeNl
7iPnusY/1kCzyWWGUZQlmctMmkqZlc8Is0xdn7nxdMLmLiDQPfgX+2QQQAML
ASzhy0RkDM5DG2bpdJ83XOY6ZnZAxhQO3sD1ejwI114V2503cHadv+ku5bD+
43fuijHuwu42hMJnhykp1X033PnCGC6+qDFHg97uudlp6+BT0jtJrP/XeIfc
eOYq86l71g58LdB/Vi4gmrXghwqVSQB84S2XFzoBy6UHb/yFQSoaiue0eJ+l
Qowk+cOyzpVVnxI1JnvJz/ZZD1P2JmLgkeWzdMqrKSjVxlibTEYn6kQxgGLz
+gr0/CC88KtwHU9Oji1M5xA1odAYC/3oxFxrJTgMkVym6z1B6ZGYuQYlRkgg
vEOVcy0J4oqS3WOEtDswNj2rS+Um0dsUdHIcmItsFCpcofFvTKTJVu/3OMgD
iiPYKsYJXtgQmSJ90bVF+xxjW0A79Ix35SUznJ+4RlKzsVrtBRr2AHW99Axo
ycVAkxiY9tk8+/eVWi67rNeQCAj22XFi9D5IX5lkZWd25xBjM3ULSZo61mNJ
BjeP+NMrhBPwoGuayLRfOSJ9Ej1XxzIi9SOYO+V25Ugt/qkFvjzWe7/4NKX9
emq/pVj8gddDfWcO5CTpePKdMXUae7g3RLO+otnbjkKNAYVJQOFUIaC1/Kxu
zUIZsojf2YTFGtpn0IKkv+JJmwEUsE0++70gEDf46nlXG4KwqQDI1RwXf169
ML1xddtEMWezkufnzmWvrSa2OU+qiw16mTe0r5vYbnsVvuT8yjP9IQdn5oNa
XKnXwQXE/xG05lSIYK6qulMFNc5+u8kbgGKc9Eh8z9dqk7bhEgKwep2n+R6a
BGEwKbumqLUos27tijA9urmsOHmvtrnMr1pHuUeK0819uD6iI441eNzYj3fZ
eQRMkSfzBQWzYpJNA3sLqVVtfNgFyxRTVvU0VmVEu2Pd1ES3NuEuYDSKr+vP
KSoigcqVuhC8dtVh9CdR0v919sN6CwXuUAOJAuVCaKFuR6yc4Pm7LZdwjMcu
1piIAtZXULYsZ84D8oQwHoEQxu3kzjKI/zYRio39jnfNJvjDD3Dgx35pvtue
mVnkcnFRxLSH0Ts3mY2kfHEjxaivOX+bgKRMzF1uguiFpRf+G2zy5ht+bvFW
DT4inmpvoGScHxykH3WO/5Wv9bEAnkKNpgYaU0AJ5f22gvg00ifOQrrboZFa
kreIFYp1MDXtYAX2eCkk3wzgDOqbY9xMaAGdoXEWSxuLb3dz1DfqBrjcnumf
CCIFG7729wuxcH7seYf1oZTO5XHqBOqzpjSHZEiX6kP38fv73J94yDLNKquI
e6xGgQaVZ4lBZ8DNKoihQZZ5fjGZ8H6VpnN4R7WAFt09ez6mvxvGuTqjdjJF
WCMrEPYhIv3clqE8IWKxj9C4Hx6d9N99CWe5hQk9DYhodDXGP+48o1Uj/ndI
6bXcuNX2LQTeK8gkgIrci9AUGhhWXPd9kcsnpQTwu6R0kBvu2hSSYhh8ywee
QT309iWwuN3BtXNVV8secxUOyAdBbFnQuf/3p4pFmkR2cj0+fab4ejSPFvyG
iHGOq1TeGmGoA8yF76IJazuZwLTp8kgCejGftvN94hUKU/Xs8aWhcn1A/3Gc
J2fcbuCrTqea00lewHlzJZtJPgBop6VDj38oudOgl3xnRqSvXKjMQcwmuM0R
AG0jyL9Qv2wW6QcZCQnv07eQNbaflPTtLgVYeBkcsRNxykBjfTVekVmLAn6N
7Vb+O8PmlbcL3iJaN97bAjdv6GhlErxUOtetgXfBkxELWZwUHcwt67OE29fO
JhOmUZqyUlrFeX4UGmuG9iJR+ZPVpWFarByQmFyLKGQH1LTiRZjYxEeatMt/
6TeLjVMbSoXrJRiIkulJw/1DYNBwLMIDlQlpG8+YIft1GLq7hBwqRI0PuYuP
0XNgG8eO5a0YubZByNlp9U+x6W5ALdSWKsBHO7IviwqKyj7gD/IawUgf+t0v
zqRY2/w12JjZuyz8c3cAt7QNexljEBedI38dObN1Z81ikBkEsajhgcUQTZXK
ILLS82+5JYbd2MZMR92pE79KCEs761bcerogfDgFTeuVN9iDl7JAtk7D7cq+
/meWSvvs2aQXjfMDL61zye5lQHU/cjlCqsjBTIPHUKUP/PqWtg8LsqWCMiC4
M7V8z+a/zwxcQWepvt4xqQ3V2EUrmr9yBow3WxB2RpIKmRMZLbBsWE4BnPbH
4jSpVLSH9YYehoylOLjKCqlzNRvJBIcFDy7uMa2giPn7gWkf3dn4O20mNliI
hAxl3dtDKK2Nf855gZCfCxXEyqEH1Qda6mmxeNVOhl3AXIORoHD5uSxHuQRz
tPSQQReJ1He9uP8UYf2oCVZ8fph2BNzcd/OhfLg0GYlZtT55ED3QfpC2ZyFq
fzY13k1d8a5NhxjidWuLjyHSJV62ajnnN5qx+hLw3vqqEM+Z8jXzoJW10tmm
1T7yH6xpJ7s9eaQA32reqQbOA/htQgrlnzwN1x+0GZ8964cYFFIKmMJMyYmG
OSfOqepFQUkBWfcmD/QlB16Q20ETyBXobkRp7evj0qwM6nWaQMgXd3xqMpVh
h6DRt94yllcq1BxX0MocCpuA96LhhK9VHiSrmjtnktmuV5ATeLeE4MPk2JV6
k4kot8gWgmudUjeZNlOtYTgXxcmGi2sJd17yUB/h67K/ZrQhDaIFXIfuTV+4
YUrJJldWenOojZ5GmxgkRrLscl9u+aN5Y129RRTvd9eTMxCoyHC6ts/Lj7nZ
Q7VhwftR8btutkLlzFWC2swy1+PQpKwKWvD79YcGX23BICrjmuS8IjO5Xf2p
ls1ryETJCz+J/L5TKv6M9LmUhTPrkT6JMG29qp9zqeyH8WCANJa8ECLRRqgH
yz6hTCzGmIwt2cGx12TRBM0vTJ0WmFV52LEStkSrfzYJj1evJP0PwMQOQOPZ
HnqzJf4aRrsH487Xt6ZJds6ggWBAjT4nR/ot11eGDEM1C0wbGIuTuuUb2wlk
Yvx2lfZWm7iIPAlarlNN8KsqF1rLRuRLycvPF+LOi4RJRKwzyx9tD+Sc63m2
HEw0yGkLu34DAKzmKJVZlscL7FPBq6OLYoguJ8ME/rfqRM3nrA35nQ+Wl/A1
cbSXIUEYgnJ3eXVo2Fd1rI9QwfQGV74M1fG0p8czQbpJb60cbKR/y1Cvli2A
lqUTOvRM8pwa1y6s+OGV1B4CQgeeoufhcH/cOkmp7G5AmEV/Jw2Aej2GIyUb
nN9hR0Qk5BqfCP1BRzCALJotZiAeZ1zOVTrQj3kK8NbL/xbG/wLSvBmxnbQG
2LF5omsCf6eMD08VApf5yaOymJSMjPmqwSjsnGKgq2qkGTOQqbcwB6rvCA+w
7ZP457s5ENOVoeEZRUcVZWpJL88Cp7Iyw0ryoPHQJnzXdAXz4XVmI3GcF9yG
2NWeh65XCsVhhU3fcMaPQAqEnGBTT11c1HUf12aPyv5vCtlCgFCAEWVr4Seh
fg4GtOyIL/8VpQx4R9AZ+c7WCPHjISJ5eylPvEUqzK4Oye69JABk55QpXZ3f
qubPze3Sa2Fbc725QkgyjxuK0jPX9ge2IhH23tMSbWwyR4FH5OIUe4ByAmfR
Bo4qN6BdA1hi0X/FhrQ0Lslj/cGqXuZUEqaWpeP/VD1Z5DRM7u3QhaXCFT9O
L80mklNEHr12ilzQtj2tXJccaKfZ5DsAtdWavp+bdvMz7geoNn92Pc3aGEqJ
S3yX3mRcfBolXx7wroSZb5RLBWTmsDVxXp9JE3rOOHkJ4JghHOsrVYrdJgKd
wHChwDU6sTJTnrdFXOVmDfisw0uVVvprf/GlH0UkUv9TX17l2spWYTQTL42K
GcZSssRX8zd74e5ezM1B5IgvPQysl2DakfTr35xf331odoIGQkstJu9luzOD
ie3vYPrlD3VUhlyDG0uXBvgIBT0Cea/ookBLgraC5tSrbVcWmSvujgAAKqu6
Sy7/tmHkzOg5aO0AaEe+WdeMUDeG88n81aJluAd0wpLxh7dOc6Opoj0x0D8D
xS+gDAuagFAyLeZzjIyMi8wsC1n0HRpQMLuDZGkIz9S5I7dFJV2Xk3vgGiSF
+7rZJczWTj0xZ6baP+6R+KWZMpsdQfTo+2lTSY/nZsn+bFOkByEn+/I+gzqN
Q6inlSkPswTK+Qn2q3aVtktW4H+4Bzl007pgsmiTXBNkppuIl8AGZ6FtoQSK
qmiJerVVuQ0x0OBW1Q7LbTrvau2iZGLfAW57OQgHQlTn1/z74Yb1xXJs66Ds
x4op7N3ZNmmr4SCnJetMW/9iAsVjxnrcZ4ELHx6tCo3BGCgjBL2EiMBzjTeQ
MrjbScxuAmecVKoAUmLZ1616sTNnDBJ0D7o8dkqkRJIICm5KhpbaXl9KgbEH
H4V0ClPNQOfSvWZCk1LrzSlJhyNhfDUgFnIOEuJlUls6+MMhVzeHj/kQqpAC
oZjGOal8KG1Hj8l7eZ4NglDyxQkxYwfq9jZuNrxmOpoB6+ZiCthlUKjLKmZs
UOXboE4dvzt17IUa+SahsTEslb+JX8nqyDTn9D9usvSzOhoHkYbA4QKthBPm
P/AmWiWXJ+i8SGlZP2ItGeYzc7t/ddT7QU+g/QozkRl2KK5lDHth6hWYPeiv
qgrgFyxssH+r0lIFPhAIKC1YSeONBEEV9YB9I+ILhTlTrIUkYBlT5t5T6GFd
flOZcs2TjI5FDB6tGQqLqNomPtwCAXKsFkdF/wYK6GLFUeBwaqtlX9UPDKmS
GFaZJPRJnH1rhgawjWHOa8kgUbvD3MTGbYIH1K2nA1flhCbvh78vShor0wAH
aDq1careSuLivgcDh0lbSNJEe9iv5bH/1Z1lapUzLpoNrmj4jq8qa5DI2N9Z
5rEcTPsZ5jnWTApjSOmbDPF0zKdCJN2htIP+dsgBV0U2PPZEVEm1n3DUTcC7
HZqgdeodF0SbM4Peb35REuhLkDIs/ZwX2ofsjAvcuGc5FntnyBR0752f+g18
pCmTvNNnJhJwemiK3/4hCfIdz4JiWM119RlfqfkzZufUcOmfXA6b2R6iGmTU
ykaZ4CRlYM6lf0ka2bhyLK4WfrLMrVWnN8gsMypEo80s9OE8e0kWw3ghFUCl
hV3Y0bklg2ildckR7zqVFfydiU4jF2W6avFQs7jb7ozkYXameG8JoHpv5Gzs
ro1pJmIA5dTYcquhmPdGTNrX3xOe0qV+rCTYQOWXs0Eh48/8gXsSchS8oAG+
1M5IVooaP4gqTgXvY20LphrKkdou2wWI1PmJVRyzAXNxXILDQR5kZuaULh1K
TcbqlWVy6Q1yJ0+oAcTXfFHwisoehc9srkHbi/195Jk/TEyLE7OiPlvHvW9L
4TlNcZidcYAPky+CcF5cBnFTtd7eSFw8902tdWoNh6oZu0VDp75X64RNZVPR
kdf6FFiMCcCYs/U1vRrPKYR/EFAdMc7CIKyeKNmAkc6MziI7+QEcp0bareHA
GfFnDF0VTaycJWm9KNnt9gqZDpg2aBe+W4oM7ElHX5xLxdjZM0/3k1yg8Iyg
yOPvtmRtny/4AJ9okcK8NGhaHGiAE42JLHyvSapNzOKheeqcPeqFx5Hl1kf1
MkNmrqzlugAk6MytFKw3eeDypuepgXJ90deN7HQ3uua4zdYmL9nYwm3HGpuS
qgGTXUQp4TbY16b7wAdLexEKRQTnp+jn0XZP7UwXN3Uv8nIWHlLsJJ5KqTbu
98klajFiwHyfUiXwV8CPZi1yfLe8m+W5cD0Yt288sO9mJMlWK9TTCQwHqz1a
lVQhScBD6XL4JNK+inZHRdW2vAhML6VLmm7g6Hrsfj2PJ0xLpR9fODRP1ciF
DK1mrh5rVATPS71PBfVCMZQIUAk2SX4UcSdK5fkf9QPd8ljJYYGqjyqvo0Vz
LjT7rVsAVdHWMxNuCgHycAryiQyyHxpPX3obSjaerUzIRRqvEjNUGN/LvBfV
0uetGN/RS5ZPWkT9SmV1inEuNHgvebhVrfJWUhAStay+dhrT7heiY1CoePPH
tW2LrNVCX9UIKUbWCJB/vfF/QcijtNSZtp4urs6CXC5xxblas3oe8IJUoZrf
AYjYMIgP0AQOk03afH4E3q6ceoAqY+X/JDk0iR3upjEASnzPv+XJmzWWGPqi
AcU7+RT67tBUAA4piTTiyCWpmRaz2NjWk4xH4fU1j4YGs07JOn6yJgzs5ByV
Jyk7wV9NRBiDzKZoPCGwcuix7KJbdOkCy1DFfkKBWD0GYnoYeeMG45oarVYS
Rkurp2BN5fjNVKRTqOFWQYN9e8cdCv4fWZAoLGf6mlUkqSupEOKT2C9TSDKC
esN9ZAI8mJtYMN5CMBwHdFYNFNhIhhjk8wzDXsoP6Wl8BlqNaa01fQvml/iU
tYmZzGrYYIhto4rAeKOb7gxWGAseCOv7k6IvX7ips5tkkcXsfrvgrrMCdk2C
NMjU5i1T+X80ARG0uNbQivPW9OpBMw3env2eiRYqejYXFOePZCzZ+L0y0F6Y
vhUAVoOkAAPjLHveHe5x9AC8xiwLNHAg78kusjNoRivZ5FtPDiJP+4wzpA84
bJg7Zvbum3ep4UuZ4XrQMNPzpfr6EnElNqAXfLA+frPEz1py43Q5+D6wtIEf
aSV8T6rwbW0AEbRVIVC0CDJf/MSj01hChe7YlXpaRRxuU25rcIYnJ5Eazw5M
xyvoHSbBOFEJXZMxEpRAs4sgnbQJaxTL/5syCeFXunP6nLGWDRqF96ZYJ8Y6
xCYWxdiIr91KGnwCFS8W4STxTRXLKK5fJWqf/HBCFnbLksQ9YqVCruQ67J09
+CVXE0Y4s5DtywQPjZzMCwzZm8oJNQ0TfLxRdkILJgUuIQpwbkIAGrHfibWL
r4LYbmrujOSLh70UNg0OZJTmxhP5X6Cm/jVGcWHxIr8Es/S4iCTWZbyTNsuS
JUjifHrssvUWtJsZ5+ei0xTcn0sOOWAONtSEmkBzhGGlM3rDpKBD+F01U+ao
EORrOqt7qi0R5YTnQ/34yXtEatTMDgyYLIDJGG1eCFlh6KXKKattcYGXs5/l
2YEIY5sOQT5oNsLi7jlRALxktu0WHpsmXTb15xiTlmMTnjv+QcH97lfBBCUh
fnk6KM4mF6GtMzgzmN9wAUzClZ9nGIFjDLmNLSgbqqpse90K1kpGF1Wp4YEH
X1h6FsUmCnZ7Rf+qmHAix3DOr2z8Qy0c6p3jTrUY20c2o0bHe26FNqpHH2uP
/X48TAf5dRShGe/A8UvuMm2x7owfHeY7z11NaQ3GlvFI5x3o/pjTa9R7Lj2D
SjcW/iQXuXow1g3k516PQ0HOEn5lg7nbxi39km5OP7A+6gypErGzIjFZva0C
TME/X2rK0JDHsnNi4hQEa6Yq0/h3h/ZSeARUkFxuBxR62IC1oWguCoKiCftA
RM2jzlHD5+wnOq0UgPqdglj8zhkxtvCB+nQp5kLbpCTSu0+Wfs9y4tH8OWzE
Al3gfXZCKXfI+KKqIA9JD7jAr/uv8BfN4GTEbyUqoDCDCCc1NgNGI6ncNawM
JtlDXONW003U7iE3aQ3DGnTJ7igMZsWIEZD2XIoN13p3cxSVwSF0uxUFAKPU
qss7SZ0mfp2NLCBiJDty+mVJ1z0/aivmy0sbW50uIPzsu6sBseuNXldJzzot
ozYPjUyqU0ZkZQ3D4eB83dpp3lLjAPn1cTLFAJQqRdKVMSPnser8WYtmHwhl
vDY/tP8mmFFtk9Xje3P7IyluoLOdNgG3KGMhJ6eew7X+gSs4h6ZcjS6e+Vpr
DIaSLNWkutWEZgQUZnY+0JKEbQeUnTBeuhX1zfHSElm04QGSf185ptPgGT11
KJQB65PuG2Nc2bW7/UhuyL+LrPpES/z7SYqG60CCm5U5uBP2f25dxfDGI2SB
htTX67pBcqAvAemFTe2qPhP9eyAiZ8PnrK+QqeIItTa/ljcW+r6W+/Yl6cXM
8YWVx8MthQACjTNNurnKmkm9NHwNQ62I7Qv/coKOhyFKVcszKDKaBnFtevYT
yzVC2q8tWV60XuUrIEgkYCiziWoMGy6lrlz/ziYhsmqwjmYkGUwKTO82yA38
dbW6gh1FSA2IlHLH6guX20rRf1lyivUxEZYx+8BQk2YrF4ULNJ9wqsUE3O8m
BFl9zCvzXOh90mlXTJ2eG1jY7gtUzg+QwAvXK9G/RTcbheFJYv4CxkkPiHbN
2AKaWK2V4opjaDEuWgp2I3+zO78Dy/K5Vipw+9dSXWmDb2Rn/7OiP8DrVwXH
rEUzHLPVXTFr1qx/wq5xifMp+RrgAYUBP2X5nNT0ngG9MZlZs42VeyAkzVK9
sxG9uMhtPHACtQafkWmA/WFp0v+HYLjJl1qGfOBlOCMLr2ro23KC56kWK9bz
z6d/a/Yq81Hu454QrZiVt4UtiRa+xnofSS2QFKiJ5wHD3w6vaNj4DPN/ihFe
4LDTgAoSZhhMHLERnVwj9CWpVfOayzssQpj3O/KB670xrIIr2LOY3ElrieKg
kxUMnE36TWncnmJS1u6PZnzGWgB+kFI1mdtrCNSxddsCChjPy7laEkWXeq0F
StJ5pQC6fxRXSDqKL8hS4rLGywdCjcDN0SgAMiENIoRca6CHRnMuJtZbaLHJ
Z93ZolwjT+ZgMRf5Vsyeu0bBO3YUqTW8OJNAmx5YCKA7aCP7uGQtBPUCt/V6
kSBsPs1tKWxxnh9arHlNoCgsZPvordq8IvAqr+M6rZ0bBFA+Wh1+y4KRJ6/9
7gz7VZsXhIzhhDestghA74MAf2RYV+b4EovEGONcn3aiIIITVeX+VSdcbegL
NZ6bmhgOs3zQFGoN4S9tmMbocMmXOgkj4UwC7H8FQIT+uWg+n65886jNvI28
gGTr+dtiZ1v9/6PVNi4NebBmwA8SFyW3sph90VYeWNHe64y8dk3LJ62rkr2Y
pC2McGQFcEt1MQn4JYLFKj74WfEeFX+39VNzEAoVx5weG4p8QzOmhJr0gL8y
MqDYyfZ+//y1FQ3hstV/DLauMCWWtaJNrB/CuxhUNn16TkWkai+41M80LkWz
4JNV8x3NPU7IyRot+NQQj3dYPRqo/W81m7pozVATYLMm7bioamc+s5RLVesZ
DCZc2X0Mh5c0hNEybevj1AA/fl1u/qtXAL6VgpAXXcdtr8IBB4/5Cy+wz81G
ONAiPkE8x4tP3P1JbNdCH1QyLIXkaClAa9DYULShEmEQse3hvbGzbmqO3/eH
0uS/ItKco8Iup1RtfIa6x0C+5UhLYUvex/5aBFjGFhRjBgnWzyzAJmJkS9BU
49Q+lOvqmp9P31o1+C4jL/f7FBC3UYwOmeKrSMDKCxcvyCzZY6+Z0clU1zxU
f1H9CWvxiXEkPk68VQPXWCK4msoChn5dRkOHAbkYV13Z9+Ke7ngNChhx867v
HdqK0EDepmccJ9BHUrwIXq8c7OolNiZ1lZHgEjitd4TnT0j2RZymUT0n3RbQ
Wb/R5Ia4cytSlONPQOA3Pukar8sP8IwNU9E4B7jOh+MfKj5wiNh7HggHfV+M
323sMyz7XPWxOUXnxy5V1f/V7keqq1ENRkPUQAmQSCUHdUOqOTb+bpjoxWej
adbMoTLM2Jzh+rCEJO8yMoVITaE1bPBIEDsbaVoMbNit949c30GU3IXHJNL8
4Y1KK4cLIt9uDdQtdohzSiJHOcO17sNLQAiBvd6Cn9IQnWKSe+Uo0tYwBzyC
KvfqPmPDH77Bj66aU4fDlJ13qlbtjiqojl9qOZWmkefPmNjfXNqhxrO6CduS
VlxLnbnfenc+Xj+r1iLjNEG8j4C8wfAkUo7+7SGlY8Oy7VVIOc3iAOPl++Bt
DH7pPjJ0Jsivk6QP8am7iP+4grgwP2JtY+GIMG0oOkc3UX9BKq932SXRDZTb
sanUk3UcMLk/9js1FqxNUCoaQuPs4WkRuEn9gLYahLvdfGkxHD3S0xz5EjAm
Lg6NKVa7QuzYp29GGEHn8jGDsmJBJy6IB0WCwFFDv0DbdAY9guGT+5oLypjC
5gJewVHUU8SigsgIRud7XIbbFz9kCQvyNE3HjPnzSMnVELllOffdR5DzmLgS
1ktLhqajITgegIiIZNIluSYMxK2UwXZGpC92X7mNMi/o8CiotEZ0q96UgRMN
V42zBHvZ5/78T/vxE21KLvHrpuP5VrTlCJ/QjEuIp1irRDa0DwzOozEXTOKS
/v1s5EH8ZUIx3dELjgwT8ex6E31VAYsnsR1Ly4VAmbjVF7doL8LSZV+G28cY
vRXtiVdFwVghYGki1q5FBaFj2jtHIm/aOpCmes2aRtXbhYdZTBJkLhZfENdx
yoPFMeqIJI13X2cDHNCqiXBhyZMWbm4PK35FPcdDKcDQ+TCauEHzmu4WZB+6
+x9NRuenPHF0JGP/8I9jybZU5jxFOa4bjRz13sJ7ZbxZhKiohj/nQby/CqwU
7YNcq6iUaCCumnVX8IJEhbjlLVzrO2lOe4ShNB3OZAXbDW+vL/kICpA4X1zm
j6xhiuWUrv9RxYXu1DSEXRexj0HsVxi3d0r6w5yMASmeKTF+HpmsTEfQXm37
M/dCDjUGjgoA/h7JtMO/Wba34HjgFZT5RgaOuG6nngidaRvLVu+w0Lb2Dyvx
ibu0T0j9aFg+Y9MKj7CMAoRRSU2nAj9/qUM24dIz6jfsgQkdaeZOUoWYkQow
kGkaF812B9uRV//kkj51Bz3nwWL4luidPqAgbwTrxA1AO7Fr+vOyeL1lEGE1
CqwoaO8pzfL0dGHZKnu++q67H1sg+8VLuaSYPYiqiQAzW5LLHJtGuzuRf7pZ
jjWS1YzgXK4VJdWhwbpmRyUienyMl5pK3Gb/JJ4i4rtrrDPUNZrrHhYVPV+J
gFa2xO0yqjys47+8XWL8Xgggj2Xn+0NNoSeCwivprle+Ilrm0SAe1VenzWAR
Xj9eBa7Cm72nrecU/ZPt4W8bXmHDwWDKEPQZ/Q/0ERO1bGGL01jJ3rkv3e0K
W1UwBjf9Ct1mHcP5IvG5RjlMyHqfJXmBaMESYooGPlQg4C/U4fbPR8D71lgG
OH6MopYQErE7UjuoNgnk2EnoHsg1LkuoWSkqhV9gZHdxhoFMjDW5FzhAM6Tj
8l49XKc39iY8sxNyk49o/NYgkFIyPRSbaT0S7wq9ebtU4BPUWHdZxFa4Grg7
JmqO58toKxn+FnY2QIkN77+HWAivc3iB5ZbcF07Q5eCiL3JRRXqxzGtyqUBE
0o8ugqoOPw0/uoYI0COv6j2HuZruRVR3stNb+UwD7i71WEKagUk0j2ymivBJ
sMhZbhXtq36cZt7x1TCV4NW3pF417d+7KrtfosmI1XmZTrxd+s/R/6qviK7o
YKTC3J2vye0tfGoyHYRmc936yIAz3a0jP2jKvwDZW6iexF1080o4HtQsQbjl
3Uj8LIqWCRJbHYcZGMsvCf66nRL65QejrAyqHrI2pLA+e4ck7McvS/iM3pcp
s3j38H8ctf3uswBGRhK3rRIoZvrKFwC/elivIKoxXd0e/H9NuJQN5Gg/j+9M
FycBA8eEO/v39DYJqOw6w+Te/E+B03RxquCBFZkUGdaQ6YLHtgQobjctyime
2EQE9GpK5DXOJVPSSZCNy8PDSBI7ySZQWdzTvX5BIv/6HcRNTHRtbKyIawoj
cKQC6MbVs1vhkL5ZhPic8RJFQhq+nuS4q/4UfHMB7829GBU71lVrpEtpzpSM
s5wTBpU5S/Jc3JfwAfBMVtbFAtPJw/wtG6Il+1XocER/Vw3j9T4QiCteqAeb
w+Z++QAa07GA0mvpAS2rwTYg+rMRe/FPoP0vMOQL+KqELAtepWeEMzxH/86s
Wbg4RVz/AxSsLvilcCieu+tBZgI7jKSepQLANEouIWxnJrokMIOa5BrRyHfP
jzSvIB6BFrlIkDKwLVXolUPYEZ4CytDT3DiUqUoISfhxeoBJTyjU+j4iCLPI
nSIlG1yIWtJsstryXw/1S1q8EEjoUHmm8oq6aOsewsgCl73KVAmItEl3XRBL
cOnESjkBmD6hJGqhJ4W9AehX+03Mo7BTCGzKAqQWxRrtQNVE4/d4IUSpDsHQ
hg34EIke7uvwYpyeejZxbkwNuWuKEFMLVR6W/4HpWjOpCr+hVnGb5JSmqIqt
24eGgcmyx6LPWnbcaDjfsmEZX4lZSM+HJD7yNRxY+a43c5jawAZcBsAfFbRo
I8BoebMifM/oD3RoU5/GG31DxuThEIkAX8KQLnziotk4LJIPCR6ERimW3HYW
peD940m+zXXABUa8QBBrsWCip39jF9QkQ96gRRA4WPGqtFcu2xdhuRo75eiu
47Axn+mbeCsv5+hUFeI7dtPwN6QsWV3cU5j6iyi9yHr+VN7OdLp02DYcW3Qj
aaBl4JltwBLevpWURQiWOvOzziSR5Qr7zaYpBDEj+xqq8D/lPO3BYInwaX67
M7ubUPwZKEQaF1X+iGmhFm/+JVPN/8iAfZ4OAGTHh5BCV0ueTU+hQ85ZFbjM
eF4lxZboufVr5IRM4mJdrVavGTtFiBkhQZyxxGaf5+34Jk/DNDZU7s/tOmE0
yBqDm53VNCb5+Ip7UAW1vyNlM+nA8loh8jkvlKcDrcFFQwVuCcLt2o8WzQ3c
b4vWGPnT9mD8YKlmWYWh6rDjdU1GDex4dSRBwdavU8QOn7EguP2WmD0c6QdP
11R+6Os5NkM03piIWpXMSZwSfPLJIMUe3nQl7XCo7vQ6cbld4WQOxysVNwEY
kal8eiHYcaBKe37hGgeD+x9PFmWiOB2/swQzwGNug+jyFyDiUSwFqDRwICEX
Pz+5SCZcGoiWfYjeavGITve2qC0jD7E4a84AkJXS8+DMHiv6X6VAyIIRaEOx
sYe2YXxbsgbJUr7Xsd3BrXMkuPLfg2H3vVGP3nNUwX4WQpL1m5ypx2+CHV+M
j9YCTY+P5w/88U283576EN+Pmni/kn+GtJEdjZPz/5ssW/X268XOM75JGePT
glT2Py+JWiAWQvhAxwhEFfRqluNpM7+Qx+BiLrmMg6IehiJ1jZM4K9pfVmlF
gSTGgBGlBHvZDCSUkufXLW2O/oUoEyoZWdLFtYXxntrL9PXQQlkcN4gw2abn
EuWPhUoBpCr/cPM9OItfEJrNaChV3JBERl84vYgzfb3KrG4/iCOxFaGxcnL3
Ff6QpIgMV9zaO5ZPGDL6FTbIDseYKxZ7JUWr2C62lCtMclsyP80lMMSsnvc6
ujmoudD7RXNht9W6h/pi2091qmPII3/I8CHiiroaavfoDmxTypZa8PE3Byes
DPvJxR6Ma09PiGezfPF7C4wdQr0LYLZTE3EHDUfIpni7NBFx86HRujBVVvzI
J7Y1frF/O7eDWFrQw/0/xtdn62O40TyvhvRRB6JBS0ZZupI3n+O4cNVcPu5f
6QWveK6Tic18qfjfx+MSkrBqne2qGGzzB/f+drERdRqSoxcKpbArjufZQUzo
ju9vs9qLrgLR33TUUn1g1tiMuKu8LCgQR7MGSazSRyXQZuv6qb1pT22kMrjO
O+5IVYMTuQ3/w0NS2X/6sOACEIfwkrCMTjtokNVzVv+ILr4rmXziC1W8T5lo
YXpYojvLny9njvXJzCsivlK4dN7INIar5M+QjMTlIq8GCsRDW/aeZRXPD98X
6jxMhy/jyFr5B4b0WFPKFe8ewUk1Ufw17F+xFPpH98m21FgWHfdGdEk6eRMB
NMp/8pMpHeohPlr27r+i8b8tU8z6j2NAsKMrfw1hkEV9x7ibpW+WnK/ESeCo
6SG/1FARg9ebzW7EovAKeh9I006ou55HMOdnaDWN105rnko/AWnk7rhaodRF
x35+0rJyVLQVPmxMuCwDMlrEJN2nhCMbbgpPhanhT7rsZc+Qew38fjpFM85v
86nRpxjIu9T54c9quBGEwCiVxcch2n2fmxURwXtfrVS4h+wuoBZJTx47yvy4
/GzRNL/96nDdKmkCou4TsH64GMW1w1iLsJROAgJ5V9mf8Fl1ufa5LN7+KqtC
RxBZOeT4qF9TkTJl3BMz/IEqUJphdklOA2LgfzyPgv59P+RrOR3ZkHpHpz8i
Ywq5t6APuStf2KtGgw1oeu/RdQKc6LZV+//RF8FjlHVI9zjXmuH8UkSwWzQQ
+529dFmFycGCgevO3LlqgO4BMUOFnUjOcq6IaAddrVfrMhqLMlESGeCT88YP
5ekqHgM7iVU1Ujn82TipyV3lsw0PWbOrk5U8f7TJ4kp178Zf5oMob3BaTR5e
Z2+t2aQ0EWn5kxzLgwihiMgJJOl1oTOUUncTMH8fZMAqAzI75t7+ULdCKcgj
sjLlefDTmKmoCa2VPc5mpbnsLJG8IqeaxOGAWplIb4rQ6oDVmIDx2Q5EDIJz
HvMXbu5n3zGxD+ybhG067gkO/sVp0UfdhqZ3rZJw/Z/NOob2GbgWYdOv0HgW
IqUQrNI5sK0vRUsthkgvdt0CLEHbPrZVCD+HCmQ8wQU5BXi7Vu5Fwvu5wjmS
zceMZ+VxpWapPizxsLlFqxYuVvfggwe42fC47Qkdbuu+K7WSIyWIvJuFQC7M
J/JQ2Ehy325sKobCJmPkTRBywxld/pkszCJOeE+0HvavF5RBmz3EKKHYhOtW
hQ4jaQxsvBySV+z7xkYqKSWImp9o5D/pGlFf61DoLV9LlfvfA8PMdhzu7Xki
DI4w0vh0j7QBWF9vVBb9QNNUgwRow+KtuD04LEyj6GzCU0TNKNHfmp+PfyOl
vS2TnWugSfKSixxc+U7RdlWlAVSofRahF5iFteRpwbwpStGnEv++rDYiy+cU
J1jrlvfzWGknjxmLv2DqiTnTfOXH5V0sQB4I8bvKXWRG/WdaNB95cogLjRBl
LPMGZOOV79s0e4oxwEAd1DxKsfERXUq1eXHUrQBzxdF3XUnbQtAThDyUM2xy
O4CEV9TLKo2gWuMe738cpzGzAQhTOKf+dbuFGapl7xP9yzXEvQgxmyGNI7FK
AkiOmRQiOeqNnkh2WMypdQcXfWGkGuHY16YdqPSx3Ywp4FEIGqkeAKiTw9QA
lGTxXCS47sNbBAqjbqVzh38vmtwibxbj0aCA82K0gE4vLBmZ6FVrWEL/Ylhn
Aryb0ERm03xBh1eDGXMwv+RwlLYTeRmwHyFUmnyz43O9v2U8TWqoZJ46BWoc
U/sO94vX800iZxWxKqrzwwcL2cfVGMa1UF7ohhHnNmmWMk3Usino+xO1uGPB
HcBQN4C/oAN9W6rAS0LwvE6aJ1wPo/ygnMJZ29ibRgtshgpVOw2FwtrpVtvn
frDPgzuFG+xamx8Ilx8HnmxW+SWKwM6X/MpIs7P1LjQpIctr4JtnvyjC63HT
tVxrzppSAMAq0b/X4gjnWnTxrY1NZxs2Kci4s4brwYjqnWwQGXkvD/oo7IqW
iAVeV4aCCTxzAmm/Q0SZhYtPQhlkOcFVEGG/OJI9anRebgHnWr4wbsEyreG/
sTmoU5YHK55k0Ty+rn/Kn+XpieuhP0wt4dDMUdo8RiaoCb3nuK90hQcRu/2D
T7ITPFtl83EgutKi4Eu1W++R6Qe6nVRxk21tGjHjPQ0d5j9mHSFVM68Iyg1z
5SDRQ3URBnDxy3nAMxU5oJIUFzsAGXuZR9v2M9p5RNnpbNEruQ7nX/C9tBFx
LXCAS8adQoVvRLVHYkKTpiDnixSJVgBpj2/uQ/x+1YJe4T+gv89k2Dg0piuh
2uRR05cDyAXJNsWSSQoEax5Rvoan/4gBYMFEXPYnZN9GCDHXfKqGYuHASSRy
f3Hw0LWdYXaAqy0DFhaz8MzQGLMjVB6EbZRytONraTMPULrpkaLet4swjMMN
tz6Y1yuwUD7U5ZBcpnhoasGTOR6mB0QgocoDIbW9LVEy4Ybqtjy8beN/2XpR
UU9V25zGC+UIiJyWUjsnRArrzBGiYJ5SAjJvBkx9gbdhEIb59ZfPe6EQbNBg
5F7twmjcxiOAPPpHn5vQd6aCYaKz/aHdhRDTJD2Y1qyALUtyO7jA9KByrNxu
OQ1LOYQ5ShHEPaicDGjbg00BjcVxn2OAt6x1SRNlU9gCtcS/ky2A8BMEZIHK
c1kdwlHmC0Z45zcGX4hrIuSXoeJK2GCrrFO6Kt9WxIxOkgBUeIhx02hbIPIq
KnrNns5XjqttWmSNxCiGZ8q+z6Cz6DbQjlhrWODONNW34j5OQnQDLEbqrJFz
6fJvOdtds54W9slLqZgcIN6EPEJielh4M+2dA/0ihx1ianlk8zt8g2bcbP32
EOS2sN2zj8+yV+gx5t3ZKReEVvuI7AtKzVgYzYoEcuYNx6QGgchnavK8GJPz
nqeYUuSomKjHB/Uvmq94T0vVrf69P8PJAUnFJ1J3YJPMAqD/pFhPNNUMrfU3
IgyBDUQCryPHKgtPQY1P1dYeFQQSMvvrIQg2JmNult5j3Fe7ao7J3zq67kK6
8enkRXk5l9w6qe/mI67J4fZoeDqcA6lBrqxMv+cdaNvBZKUX2xVF42A9tofO
YaA8yFU3B2opKsTh3rpnrZw0fxUIJaucrgHCRp8LTlbsNluxXb7v+lOtUsR9
dALnkDybyCJ41JMXUxmiAFwtjlJM6OpVj13/tEldICQ+/RUTv1yToqzk/wyq
GGzaEybdsqNABdPuZAKjKW7UjYSEga1nkl9IQTfdzwMSSGxTualMwagZPurz
YJWy52CTuidceLbjsGrdsBX/6iOfj3/qlFY6QAhHoJ2ZEn01JuYIm/uhf1cY
8OkAumZ9F596yitaBGzxPyALVNUEi7boc1ztrqyiq4E8OEU38FikxR3dOupq
KQ4fIjX4FlXYVSuWrJsIw+FKupzJdqTjEAUoHzpY88lXv/rGCGqcR8mej3jO
EC3K4Sq2RNGlgy7VBY6f6clSLncZ6ovi64Rc5L7xwos6A9fymcrUn4o1oMe9
TH5Sp3Xm5Zj8ouRuif+j/1xitg1A5e9BuHO3SCk2FcmjP8llskDOkHNcuXgD
s4U7veErJCdlcY/ovI+nKuddQpxMWT2w0h+/GX4Yp9ufZ+gNUmSGnHRZPk80
9X2iguEeTS7sRBf4BBI2vidI+qxkSMCz1z/fvNIIUCDzIm4Gcsf2Za01SIXv
+PxH+lw0OqT7qYBCNIpS4zXwInYtth1SVuVJL8zDYf9wioe51bbpCP67owb5
fENQW/ZlbBdal/Qqphyom8OLtdKjpZeu1Vm5RPysHbh8gj3H/70u97iUSGM7
B2CjWB/vHQzGWbaJoNu0fnqj29reB0XMtlf5AoEDVFL4uvq2O3T4AEI8pHeb
BGo93tpO3i+RzaX1vB07M39k0RqPr5/m396nwBTBUnIQVkmAI7zfDUY0cE5w
+BsnEc4gd81aTYmRx9mcYtYE4v932wjNDQb1+FWm1rjOmkVZUj7VgfkGWsCQ
D/2/QpQczte0Qb5yc4bGZ80VlP8TEtJCybgtPjtMCYFn6NPkM2x9ZDkeoEDs
azZE2ECo1PJDfh2BNbqpz7YyRLCWa43YchcgB7mx8BGHliC6JnEf6rKwoc7s
3MBe/IElJCIuE7K3xQE2DReptz4gc2g9kBh3SmeyR2aRdBdWguTV2RIa9omE
aPVKkYy2AP5TBQDCXR76kKV0pr8k++90rgfxdvY419aSmzvX/YUtt0IR7ggc
imsZJ3yGq4pvVOFIajygP/GyWMnPRbU8LoPJNVIbBcGpPAxOv9mobaTWBAgq
0XcKbt8rR/yK7/rqDTPtCR6OnwB+QI/Moi3VndxGep3oZ4DfhFIOIesWWUbj
Zzkb4BEyGE/jjp7h/Va5LpEuKlWHia6cw0FdBUhYD65o3uVZAMzQ6co5xuy2
fLAExMBWlfLTHuBVmIVp4zUuvjllt+nTT1IaXQokvlJBVmIY9NLDFj4Qa+Fc
hqH/ug0K0QJklmS9tWtcwHA4F3aWQGsV3HoJYwqPJp10hiCXOxlPlIsh3jGz
Zse4KrsnFS1Gyg78eTT2xoAnyHkTSfY8gGA02bMv6zdBJ35yU8qQ5c9dTHEr
QOtO3Ss4WXf8DEXT+4ttqdmriN0Y8rccKoHivMR8oc2Q/cRDcjcaLjD8fB/h
Ea4LuvxM4gBEX0pj14M4zRd8+ttbW396cewyVFH2wAjGch+cgokSu7ZwGsKa
2uIdaAqIyYoRMMQ/uhbB2xwO/aQA6is2Ofkt9Fz1jvo6qUXxDUReudQbl7gl
eaEfPquYDw/0M1yyIb4zfSz6ZcxnhalfKPlOZJDYrrkyE4/L7+oQevuv4Pob
zBXp932WlNPtvzPyeH8HbamOwn0ye1yLKGIkAz0M5I/7hTa1Iockx9LaxYgN
fN4rrGkqHJvlT4Dp7skcSwyV/CVyV4LAQ/s7O5TBvBwFZbl5A8OAMQPAIYj4
CQAXkMJ+hG8Dfzcn/Nbq7Bqrf0bqSnQ7eBsfhzEYZ+yYW5kfirwfz+JN+10+
xfQpj2VXYGo+jb5t5oo977I+InO3/wjfjrHwR5tU3jUT2TNpaa7KOdVwoknh
zLStCxyMl96iUYX9rXljfSaB2foa/7UmFNcAC872jGRijm+hM8ryXk3anqEl
jiukYLoW9J08xdHd8lYIwTDwd3D7mb8wiC3cc8MEc1ln1us7AdGJ8Mk+VS8o
qQpW59a7utvnnOXS3FB3b77aKsYE8Hk0b/56mdsv47K5KdbULg/C12cd46m+
I4nS/TqmA9CtUC4CXvPWKMA8mAenOjIa8xo60GxnuqTC6TOonzMCt4K8xKMp
v7Al9Ch0w3cYmz7KnWHLuvZDgSk7bqx+8+LPr46iKTnRkq662cBV42rMt1cB
XT9ZA/O1Tnk3MMlgRgd9H9Kk91lWoB2Hr0MmgM772YcgqPPPn5mr2p1KR29t
zMgwmrlVd6h3FghvjZ9HneWtRoj+2MoL7y+jiWf8q4ryAi5bTMRZpyBtiVxz
16iArtHCNMV7ZxKTgArZyC8AP9+s+FQFcu/YV4hVmn3L7YQAx7bHFAHT55OZ
maywrboi286uE+aD8oT75nzXNqMn/33WdCV6Kq706PWTtbJn4SzA+nav88Va
lDWnHYgUHbo7ZfGiKcy1i+oGUBc1jVyov3ivxe68fyvgEVHGTAsDCmt4gSGR
0cipzfWHtCefE2ZXQLqeZ31MNfTHZgeYvFstGPOHiWYgALHWuPiTxjRgwPwV
eFL6SKaERyaW64WQFTyk048jgWiF5W7HLuccYmbnXt+1cmRy4VxSEoPSeibF
dH+k/x+BOj5gQrDpNfWTkFJGPsq9uTvxZPCDPlGXoEvTaf0lQsDVmkjj8dvJ
PR/TfzDSaZWptWoIKCQef6UByZJitjLj6UMsEJ0L/aWg3bBeVWp1dpTXyfjr
D9ngLcQqrcme0BkKldfcAbPwyNlvERASzty5LrMqSNA0m7Ybap/oMZm0LRcX
rbS6WsP4pdMS7+QUaXXYMBvsLPjiQHExOgmGokn1kaVhAZrtkqO/90kwAHXr
B1XLmdpVuE0NrbCYSfH/VQtl1QLpQmx6b63gtQ96101TKpl4jHjCcdSJyKlL
ge2Io5I82BwPiZs25K2f7OL9BBPBlfuGGgmF0sYLYlMM4c0n33aVCPUnzq1a
NfFBoc56vEE8AfdvyJlCX/q7VO+239XXrCdYlb0wWr8oeyIptCTJdQlHjizy
3PP/X/07NEUt5JVb12Co85Mup4gyNgXRoHBuCkQpSEV/0aNgr0AaujVfJL+i
RWUeJqDSTSxLZ27RjsQqxBhmQGSFcD7xfYQXr1XHl9iJNrrXq/ko+C2lB5QZ
SzkFRP9+HzDxsfnwTIX5TZ6tSlreGYlvIHgSkq2qnuQHA5n7M/6p+zRGiI7E
sAxpA34BnYR1zaZ/HbpgaZ7+GAyYoiiKOjhG3cpfREw8ZI2NNkyrsIem+W6Q
ZXoRWIfmAiWVRgI3bp2hXlSGU0ZRbEJBNoiy4zWRahYkdnGEwR9bNCDY+ffH
jfPgdOivksvIOV3icm1OOwS/s+BU2lamIm2rkWSo4ZwampItl1sKwBtSSqJB
sT09axf2foyZdAfvdxGzdB/sUpDU0VeY7ToAy9w77OXmV4VenQ6kxI9iedHu
S5EZJ1ekk01TOuwRoLDSbAaoVDOQWqhoVb+yKq2FdHl0h55dEMY/0ZuBxeMT
kRv+ZkgrkZtRugszQk9D5nqCjf/a+foC7YDleqKMLGhE+0Zagz03XxxVOgcF
0jUjswlEclG2iUz7TAgy8olK9FVX1+7QAzTz9D7o2lZ5b36ISKRrVwuEp4Bj
2jTqI5B7EoqkBddu2C8weQOeFBbEQHqWFnchpMh1l3YmcjVkK3lsgD0TpCWp
enTOH+cgZOlzXdAPeoFUFmjOXXOTnsdtcgcBp/CGpF7bmYvDrkcs3wQTNYt0
orIlBlt1WAtYGOh/ezHv0ZHbiosawzZ/UrJMczeLvZgB0BhWEEek1/R3PDon
18Z6l3803iICYQBfwiRPbwvGU/o+F36/eSQgusxglkSSD9LEcEo/WSHubUUO
DlZMjKY/N2BGnZawCAG8Gn4xNVPakY1WCY6yGX/0AExf4s1w9gywT/UCRWfg
bHebRkoLjMyNkvtIk1XN+POzRnaW2airsC4baW6m48BKhfEuAKPa6t6PY1ur
wOHJdIsmbU1+0Rv6JmexjQ5CmWYSyEH+lpvAsqQ0HUI9g2BDiG6IezMn9fDL
6arftjsIH1SEic/bareGTe6NWwdg+mqLB4m1Z/VICXXLLe3SJKhioru27vYJ
EP0d0QRHXgtyzYl2B96BPsefvFqF7/Bdlhngx7I93uYSWPReVEftTubcQJaJ
nJJW4IPDpldKKaSjPiwk/wGj+xHw4UA4IJu7VUmILhRMwwT69ps857exRyFB
mAy9ydm5vThMTNig/NSqpvwz4lw1wE0pVEFStnE7O3SUueA/5qoeke+vOeWt
LPRilC3GbU+sSSDSrn9kq/b0gDQcrMAh3aSti+FSFKKfbltotlJq08UwOROd
rTHCuHagQ1wF6dlh9a5jTtWx80ToVsOEEBzE3CoF6SVfzTw6755cCAeAZOL+
+L72Sx1HeITq/YQDx7Ibnalr0TGfmAIUTDj1szaX/uVuRduodvwXwDmmfuNe
ybMtHeR4R6PIeCKchrOmzhDXJoDSe72ynyjmLEbGgeyT8xgVQ27FqF/ugVeB
34CrC7feyyRTbnb3WoaxB5neo+l2YG2cjLsgeBGrr3WvMZdGkGZdbZAfgj3S
0arPauHEAYdWB7HtzNQojUjnrbV8Lk66m6rDxIst+FhF2+s4qTR77wGhjgxU
1m8eCVFMzSU1TRSN3mBt3Q83FjR0ZbNfj/j74IFdo3py1f8QGTCXRjQzxTig
8hKXlybQHeob+B2atTL4JYZcU0N796wDGr4hG4RIxqQXrfa+UBnlGf/ofqSY
IhoVpVp7nT++5LjQqx2QL6gn8ABw1OPCQKNr4B9D/cUvJF2Ih2ZKcZTj2dfb
bm/GCtvl1c1fmStkDY8fQOxa3ACur5XN2kFSu48j6w1whIq/tvX2mKL7sYLl
R6hJiy6qMck7KvmG8dCZ5J1nmk0t+79+JX8ePjeLbs4hA+xELd2+DgkwcFZp
xfVoJWSVGTmOxeciRz0gJ9bmwr0bBckfiV6tEmVOb+ftldJdSZPZhNKcPvuD
W2Xx0b6BA3dINfay4mE9m3iMSykicU76N7VzdUo889/XguwO3mVtrc/8j7Hw
kU8aDUIRMUnLuS4poeohCJhNEgrVCFJ9E6cy36WEUCiLbepSSARO3jgZF7wl
z4BGyf8uPVbgq8IuEORugRJ+yj1EZaw4pPM0MbhyDnCQhVFGI9nll/2Xj0/j
dKH5qGtbmk+UgdKwscNt/sfNmL0ldBlnAnJWnxItuJUY3zMVUTDuUyEISpEo
gwVzmrvU/UbfIJggcVutN3rHrFeEJx9RJvyAWBTNwfv4p2b9iX6cmBHN0Th8
4GnDbwRR5L4hv5AOQzI6tu2YoV6FWhBsiWD6sbZF1kU1rDoCImNJfZ8q4pvP
zgsc29necpy3gUFUGZYfzPrYgu6GBY1WQkQqPysSYcId16etNIL5RB8DStp/
nBeUsTc+ttlG7Di6v3Aa0OxhmMZyW3tzxecARYfugTFyXDD4NFv7kIsE1QpO
N0478+SgnCJrZady/vr9dTvBfHR/lstczbJvT8+o1uEcqZ+nfcShjU+uCcwb
m+GJmDDy864qR/qRMejU1oIJCwhtuvAIPbyiIL5Gs7nfBpyC7C+gtc0GTNzp
KmkFLKI7lC+We05uFrslTc/bA7N/FekBjukqW6ilOrNS0KYoyFiBNTuIOKGu
dSAEXSjuvG5hsDwzv7vAGxl9MABvXimq5anI+W2OrSTLP24MCD5VsnaYhNES
fO6q4tp8szaR+Iz10oeb15v0J0PhPHxyb/N4InGTfcLkEncxnwpAoqbU1ybo
s4KIYuriOn5/+wnckKn8ewdtX6Sbx0E93oGxPVtTJ8ulmMTvAL100M+97wwL
1zgxuftN7F8zErdvFus2J/E4KM4iCtEjL/apPQaZx649z9//zEsPlJpdovWZ
8evxEVjOa7abp7nR3T9E+FnIwHzCGOuPpZsbwX6+IUS3IJDHT0ouZCR6IAAv
T/0rTclBcsVWB1jxJsTckUdDyal8sQtJ5CTGLiTYcBKbDfxglR75DIOTcW20
/42gftNUXbkwFq8sXfP36++gPLB7eoikpOtD9G+8fDmnSWgvtyClBY+NvGCL
rccgFq97L8fPUFAGrfIfeNZYrBAAHtF1NU4xJ8N0rTt4u2BS0JqaPkLUxrnI
HPhtOahofP5latB9Ul8xyvdSCIp0v1iYekt+9P3+0ZdP2g6PY/x7cuOyxD8M
fJlt+wIQH7v6baw+nHTJ2XlPmEk0yR6KdaYFVtgMrv/6txxgok8iUefJ3wvh
dlwZeG2k1D3+cqUMrGjeZpDORmCzk0oxMqI6Ym6MWqppKee/MRJavC9C33g1
6ssZA5oM0zUY8ELE2X8dfeAaZ8mB3AEUqH2+8cFsl6S5Mta0G35O/zaXCMjM
2icgSVDa1CB9+V/RaMTknoxhZSJxzF6QnmFSjcQpupmlJ6RAMDZJ9xV8VfHD
UeGkzygEG9I6E4QXbh2Q0u7HhJ0N7Wwp/hZwMADgSz9+mkuG/IU4QJcIHPc1
UzNvb8m3k3arKHEqmKTvm2QhdzMpqgZY3ttc6PjYYix11peEKvD/pVpYxFzI
9J0yvP9CF9RqQXDTJNnMWod/H7vAG/ukIY5w/NJCod26/59/QSLC8M7nJKto
5dgsO9jqro5fGkXpw1LRVVCyhYZxv1jyvJ2IGxDeAKGIvJz3BPtmvZaAs2RH
Du0Zg/NJs5tPScKyu/JC7HgKvd+FjWwnFEAIdLTyxrtDGn3xre7nVgdGUVsh
Wjx2cWa8OFR9hyIkecYM7USiK0d2cM6ucK2yagoclEL/NFi5uiWTlnfa5+OG
uPFQOX4WAm7wX1gGJ44a/bYYWzUkz0MSfOfMjOIHtl3opcO0x6DTGs1DzvIM
5tL1R43CT2GZKTd9rtHOH0A6e9TDaBPxU+u/mgwo20tx8M1DBnARwICacGx2
S+Edx0cBS3yACDH5nx31jM1c8jjm4XMBmlaZKG9suJXpAgJWy3bTIpxUNg7P
sbwckpuZE81uzv7GrH81IhLcUMnIrGzv3OUFJWVfuCxQoSWF4IqDwc/znVkO
q8zs8GDM+iyw2v5scY1BX2kiVGQsrHPRGGD174q0vqnVXtHnkU9SgRUTQ4Pk
ms6kGYhIZUpLXeU/UUeWNa/2FhiaLvnYTPqHiUz1u5xR5Ot0v3RSIPx9u+6I
6ntg/9WQ6pJj3GmNxQezqL71HasayVgOCUwXHG5crytmL5a7kWRdVStGCgrQ
gLV5D3GAbZrOsxxrObtJVQAhrhlMI+AlHhbPIlPtWkU8JXHFuwm1vBQkxlUp
joUC0Ke7JOSVwktiX2NoBR4EbPL8e8bqlModzcFzEr7Dl3ZxMaIokuJL4GGg
hk9CQXegrqZ49aDB5wytbPzqJVFf12QUeA8Y5KFaMovafUk4MGPht0Wf1BTi
7NE4RcqrzQfAvd9BnmV8VXkPR3mX5faWsa+x+c2nATNSVt7j34G0sGStVOmy
jjNhM7xX0QRLRjcmF079FMCgaBRsKZFGACmKG22ZSq67TDIKR76GjNKTDvA3
W6oNvoD1HHuS9zYsBsk+rp2KyJvlv/pCbzMbZOUHojQ3/xI7JmjIPoO0pD8B
Bql9AKz5sMF8VzRAPsRdIgatw4B+7wdsW2X8YmfWpY29CUEE2hHMfuD+TtGH
1VwW4Shuxw/khjD4JAZqA3Cn5PzSZQA6Dikq2dV6Egqe+qysHjjmkeYP0Kqb
xxyF5iQ4OAkzVFg+FE16b5Pl4hXiXwixwiLHIezsa70ykQRIYrIrkcF5O9Z4
QLHuSihfKTPTxjGbnc9ygS2U/jgXOX1bWV39CtTvl43KP/SxxxadQ56pBaEy
5/9rvsQVHIcXcFlFAiJcbAD/9A5EuLQGKWFchqKh0RIRviqdF2j3L6U3Nl72
MLR7sA7clVuUwtr8lamIj/zBmuhLD5rfjwzzfnpxZlYnRro2BJwNRfCRIApZ
KFJO40f/YRhBUA5i3FENwBQKXcFyr+7nVM11+FcetJZHRq/x7JTGg7bk2RrC
rRJf27G3FlmUju9c4gNO9bZDpDbVBR9dyIXVdw8NqVGqMz3Qp85LbxsVfMMJ
aJPabDEVNrDxDquseVM0h4NnOr0LllbbPpSupAhq+bmSZ7KvlL0rYlSPBKel
rg1JXh0vYSXGtfIx8LpwIz1PqSCPETQ5phLIia7LNvlFnywMPWEGyYcccXam
JL6XAjdFpUqOGCVzh2vPGEBS4dwsReq4scJw4+zd3qrtvsAsXK+P2RkWTwcY
lB95lDDKP/V/yeWKzEM6QOp73L6HXhvIlPFXb3CD21bCGIVGW3U7+8ihUH9j
a6M2NfK+9WsPvPYrRPjD+GmR60VYT/QbA1br0QaWB4u/fR0dSE+fXefGJwGq
NabTi9OB5qxWug8uWo3a5oqIrtvkenS8BH8zpWKdAIquc7xVFMSFSp/pLOTD
eH+aZWaInIQs++jXbdHCNMG8n8/3jnSOjP7QJZAqzKXA/rwIIXS2Fv6kC8v6
mLBXS78GnSrvPMoQVys5+Moxz3RHXFghok9t2YU8aysZe0xEX0l1rJEhm8gR
LWyhdVQoWSN2DNxR0U23QcoPQXbmmlBXnoAx8YwKztWRGo24ozXLdOj31rvZ
PZsj3MD4VgiDXbylWsCF2GFG35961hbwyOhinzmhwfF7wRjA5R6cZKb0aZGb
GJpN5ReNhjaL66I3OgMEM/NbVRVEIIEYyId3hEpwhuu/EELS4XISOIRJv3yJ
CjjQLiJJW6dO2+NosEOq+zDyhS/HHhRMEXrIobYsC/OHpMm7Y74L6h2VZ9fB
SaaE7BSB0QQtcnjHEFh6gnN94oVkTs4cd0PBJ3c6xaqw163mvW1oJbL7SeUg
jQeMmd5PS/+MU3+RHmGa6+Yk5RiWne9PoGo0VHOkxGDkHTsdMXUyxSMqaE1N
ND2QothA7+8VI1tDOyLCcSFr87nfAaMf44ClryRXrQ2ZceCqqqq7Urbg8iO+
XYWUltGiczQ8+MR2N/mhzLCqgDHjlm3PdPBNWEvkHgzoVgLae8bI0g/3G39b
3zR8RZYeesdtd9tsASBWtU0LU79yHo1mHTUA5qnslp7nCLEZ8Frert1YsNSa
rgi1EPGydz2sSeOLIeyDNbCuSKoLcVjqXenOWMDE11/C7uZNCfNkAx8P0Uo0
/7r67XW/n4N/CGo2Arpyx1koelpxM/Xrez2y/8zSQZcuOhhihmPfzj/7bLFh
XEF22fzhSI7/sRdNY2HorXFVh/7iJFft4rdM+TjqR/AkwgsI4gwowLcWW8Zk
CtoN4G3pzn+8rzBeeR4q8ec5S6hLyTsy7yL+4/XQ/vYC1sNKVd9/PbzU+rnf
hx6MattoezBzwYsqY5sUDzI65SKL/b3TL1ikbZZe+GVtCycEb+XxPA3TN+3Q
jNNDYpaImUFSVbnS+N9CWIiSGlv9McG6DhJSly1FHuY3BY6CrJ5MHgGVT3QW
Zd/HMGnk4fgod23p+CtZUzSco7A8Elq97/wxF1xMnSsWugPIqQ1Bmk61JQAx
JaUJ0h/ewpd52IfKOBP1MDcRFMJJi9WDp9dIJrqVvtnFepL5MX6tJUgUFQDI
Rc7Dvl6vwLJcdl/96jGQnLQTKxGOaWdPGOO7jOovSMiKb9CATxLFOb4ZMNHd
9rpbHdAtW03E2HsFvGO0MYnDq57elNVDJimy0rmaFH8z8ly0/6Cx2ZFbpJIZ
uuExAACaq94+/360xbMMCHkZw5pC0L/gMS5kTP+9gza9e1n+EzDTaOWpD3b3
u2czOo3kuY987gfV7taC4cWpzmHlKP3r8pAw7W6IuV+fjFqYeTtgQPdnRuAU
4/1qWWoFKfW4pxaA/baFC056vNFhOCAoKX35Sj8Bb0sdYWgjitTmTWQc2aQh
K1iYdOZsgxaAmE4GZB4mZBt/5G3ih9MYDv9p88smYcNirZ/hFBKiAAERYEiq
y0boKPBshCx/4i1A47XJA61IhutXDB3YjqkjM4G0+IuLXDqVEtzCw1CkuwQE
lRh3DVZdMUUKTPacNHdlGjCctBfRDHJ+5x5avurgzX7M9WutT8q9c+Qo2s25
F+9cd/3JE6bVQkd8o/8DE9rHIsFiKEKqzJAVHifobJfjyVNvi7PsqqUJNW3F
sVnSdFdeRCh3XD4gVQcu89Zodctp4ry9WtNwMyoeAVcQOHxzj1hiOzrptsIF
f7yxaI5z06bRf4kuUlmQir7owmD/Dj/Lo33OoN7WHdwqgP7yzwTgfuDP6UrH
KPS2EDG0znNT7F0qxvuCGpPltvzhzBUKHNp3YT/PFeZ/G82ElwY1eJbkh40t
O0Oj5Iz9VoWf3LSHezG2VoV5yzr/pmBPGxCTPcD6nhXcZI+eXTnwuLiXJDYj
OldjWZSEdgvJCEBn7HH65qZFh633FliExsajcG9HVxp0hd5s1Ev+82oAIJ8m
+rHwo8sWNP8Kysyo89Gre6TDYL04C96T3O3ziM8BJ+X7b1TPV+psmzSAux8l
rZtlcLXYl6To4soSD5owI8/ZBPL/1wljU9JCKKl1tRzCtG4qslSkp9Jufz5y
YggE70jKuSk1UDmsR15L8RjTyjv1YK1SvUxbBstalr0tT6UZXetwuE0pWQo5
3BA8jv/cjXVxbLOO2fSNLuWxVBlRJxBdKJSXbfFTKg5VfLu49Y7MZi2LwOkH
UUBGOebpiaVsNJWgCIRLBr+uswiFmFKlTkjd3v+lPSuIDshLK4VOt8FASwxN
JiMrcYFgfoOINFDG0NqE2VH2BS7eE+OaDQg5CZSMLSPRCgYlWVTwaURUTj9J
TtqlZxRwpnLvHj7LvRTqStUw1kBm9vnfYTAj/A4PkgzIQPQyef8S+YvRFhMB
6+F5HLIQHB+7Cg+CB3mT1zODi069jMClqSEju2sdeafe/0fTD7GLw1OiDnVk
5HP9TsDS8CJrZpLKLKb9SoaU6kb+wOtZ/YVf/eHt8lGDdc77ZNTTt5/uMWeG
67fwqEWRxn15H2tAWyuThdKbW5TQ3Z3AnU/QhtJNnbGZHNHoZO8tkwZjygE4
Qu6ZDXKonnNYeqP3AqRmGJTIPAlnoWC8GybxefBxgdEg4z5b5P+P38u05IVT
AuFD97MWTaNrM0HpPRFW8AXySZHk0HxNrjAs/ojxgGXwadDnWvKDlOUs8ybw
unSCjZos+DJfwEzmA2uA7DXPAyLBO0qLogghDea5tPHI4SSAdZZaHooEXczP
UYE+DjjCjrrENc+T/D6ZmAceL1iRjk/GMzYJPHCQz66bRPffLuTUYPZB9Olk
dLsIZHrnye3DS+p5LXuYUrG18lBQhHdCTH3IsPgKgCuXVf4TR5WH3vBBTkFX
TF1U/SCzpL91g9ep5LUwtLSM8eO3849Trg2+ljqDIzkT9DgRuWbQOu9obYFG
lVKdyM9K0NxB5Ur3i1nafD5Dor6Xl4KghP+pYQCOUtvf6s351/is2t2k18yJ
AJ+colHEqMd0KXGcSpA6qM5VCC02SOz+VZWqca631Iqe7SboB1VIOvU0RPvA
3w4cOyCLNPXKfhoWisqdFfke1bpd7rugZITznVIEHY3EIbDAY3+xGdznCaWm
eNTcxByI1eIcMV+0Iz/757/9orkuJZZJ6G/MPQ+3owvgzhIys7pDmCJX/Rhj
1UZGHHuanGIrNG97ulWWClVXt4QBxzi+B7304wNebJseVpbfpI57K5lW3Lkj
NrzbRRTrugJCo2cN/QQWs9zx2Kz7O4+IC2CLyz+a4odDeUlepDdp3EkEv03p
94FiqwiwPmtmvZAF8osRIxo95NEAxTZoRbQkYiQfQKzhPrq+wfTr/+OafqZI
Q1OAubS92TKbXoVdeJzGqQh739d+h+tooicxmZBrgqJb5MPTKgN4ZUmGuuiI
+DP2Kc017y1uMn9Bgc8UeIIfTA698Yhh2oeOZGrFyE9PNwCTU8YfphJPtpgA
+psW3anr6jac6Q9J5Wij2mujD+9WD73QG2MFuofA7V0Xgfmj3Q0KE3Cm/kOw
+69EW3xmix7JYAt5Zd7EvBAY047ghXWbzsZJoobM/agcDkO80Rxd0ZNpmllO
B8eE2275tiAFwuibV3M/8l3rp1mKxrfqkQTeRMxHzayXp0qDgI6ROAYBu1IQ
skWyqvewN1B34dXJH28Ex0dPkw4aZUb/PL7YlRwEZ7UZQV3rgvrLGrwX1lr5
pLPcoDKr/ErPpiv8KwltSuwxw7t+7k+Tew6Zz69TVXWYphvAdZWNLXCc1VVy
jAoMknkUOP4PZ8ao0kG5cjALlL5/bP+IIu3JOOMnSxlWKfU7vyCX8f6ME5GM
3lOmXmKAXvtZTgnyBCx9WZIrO/KmNBE2SOBPGIMcL/iwyCo8e79wbZsyl29b
a3E8vd4CdvatSMae2n1JTU7icut0Fq2H8EAx8R58+P1UuI0WKWJgxDyIO7NS
k35w+C0YX7w5ALYUqcjWWdvlvWzEgGlbFaZffLVHiKm8jZOxGDeBDvmLcgu1
ZwZypO4oFNg0XpMQSZ69ha8x9U/rIt3RRYpeDBUVXVQ3Fo1QaEHdH47wb9rw
1kFDtpgdgMwLVKab9QjEIfh2ZPLNV3yPx710+AuRx58A4my2buoqP+r0ZBqM
4oLIVO7DrUvl4nrTfAoYsACEn16vVbp2W9ARyaijtzzZHz4bEMChVgApvDly
4js6Qz0T+Uu9Ij8C/ik2LbwluvwmTmFoadDnAybjHi+q0tpC977i0iMJ4zm4
o8ciynuF9ZduK46vFd01t+X2zN87PJvb01Q3hnIP+jM0r9mtUwI71m83yyWR
g+179qqpHWr9yL1AbJfs/dkNmxhKDch1znsNLD9mheKXNp9a4RtiuJPhUr5E
CGyKCd70Jnlo1UY0YVONa79fQjdxZ0J4TkhWNx/wZn3L+uhbpRqUJ7B5Al/e
6a+E+OgtSyywc4AA2TdFH1gNaJSzea8vkO3bAdyeuDJ9D/TwncJtBX/FFV6V
MEtsKVH5CWWODldybRBLlNgM+6WkBO4J+4w4JN8iOCO/Ir1PsvV63ZvY5Wo7
+U5Gp+AkDo1AlHbq+LJOJrOUJ22qa7TxrmEoDvjLDbaMqz2QMvpKsu2trwS1
YEMlDAQOh3o2AML4Snkw0ejVMvcEQTdYNwpjX5Xw3kXalGWbBbLhaa2lNBmP
Uta3k4YoHFoK9+c8fJDwzU9DNTEZJhSfYFZPc+qXZb5icpoM/WdguftI0T+l
4HzM1T3Qhh4UaNoP9OC+VsTnxS8DX9efpD69vq5qyWj3s3ugDgrqBqOrz0KT
nWoaSxpCAJteQyMvra8NBnjYUeHBvX0TjhOUMugU5vaKXQ6nckbDA/kg4Nlv
/GdfQaO9QpITbhoUKu7+2iJS0COZcCUPwUmvFvvjRZqDRvUJQvWByFACvkqM
G/a4w/I5I4HxJ0UCN0GSNliA3jronGu6PCMTTChrpyVcMvhWtVSRDnp54rM3
22PYSS83p8fMbQofjyFYFOIlHXbdL/BwGakfoL45BUXIq2xa1GOjPvNQKuLp
EPFya7Rvk1cqZTo0/8rUwktLtLqy1m/EPGHwLbkaYdJANZ8uVhzWhPFxiCK4
jQdg3mCx1MXsnf2W0gMKDyjnUXgy+cZm33p9iQlLXI+0IZNL9rEOIr0ZNedP
fPB8aAHrst9gWoPNXcbOhXKwi9nQ7Yc/d0xch4R3vrmkLlDL85ZC9ZVNbXdE
PNpSTf+RHnpxpkZvOB6B3ypUCCAncNDKSTWttie+iyRzlB0pTaoAHN39VZP8
Em7M53zH3YUCG1v55uvagEzN5vfmw24nOY94RLCeveWMv1wnHkvoWTqjrZ5Y
llDTu1cAfKhYehrPfAJZWe/fjvc330evt0+ct7Vk+VUBVpEBoLTPH4UKBUU1
EZEMdDKCX467Kg2+7g/0agtrdB6A1oKRMQLOhEqFKa0+Zgky+OAHoAYBD91V
Ux5K0rmoN1uvwtfJ+JyUe+U59Oz5swJuvCI0p0jucFOi3fQme+Ry5q5dGcSR
j1JGthcFxireUHvLSXBOEct4nE8iYhGj3J57c53byNhpZp7FykUAZcJv+/0X
xM0GdDid8qCrO5tRsX4E/bYeXYPoorwHfpEIRg+ItSt1jmYpovtLQyoGu82V
g+IFMuZvo0AcD76BvWRzPhe2d3wcpKpMrGysDgMYO0N2Gxpt6nyXCEXZ1pUN
1BD/vEdbHsJqVidE6w1Z1MtRhGVdUwm4PSs92T2G9V5CH1JCC8Y6ZuwBw8CI
ou/i829uUBfej4yGkXf4HL6llh0OEg/kMpLG307CblASePYGACTTq0+0hGZj
nmCfZc+J/kIBvEeqDH3Cvo0/zdzZwtnj8XQinBarq19RejFpYObLrDqmkBkk
tDKgXLNsEsYtQrlZ0oXe+gYWYa3jD7xGhqVvDu3PsD7V8lwvpnYt7EV3qnID
EqanvXS/++F0sjFptpe6HZ9fgpqMIjDYOcSYHbqfpS2rWoLKeRE5JL7A+GR6
MFjfifjoGFj45kOnP0JTRu2g1bwi3t107HZIhIWFEUQrlkLZ7gAmMhpaE9AD
gLfnLtcwU/jwrb1CoLDYIwG7q4AdqGH4tLymzbPq8e7lmJy9o+mJhLnM1XQ3
UIbgYy3CGs+qdq31EH65A9oJSa7UzWBuHh/zAZcEYM3McGwZN52Onqk7mMgI
oTYoscQywl1eNXr24afWSsuZA8kUukhLib0fo9Pz09fBEI87xrvTJLnTL96/
TiNaR9qXKhEHL5eY984WwdPVR2Z2lGp+AnhDakZmrzm+BI+2R86PPE2ik8gQ
Vi8kHpYKN/asVOJenopA+jsynjn8YTHij8FcmcySSodVjELSLkebPnsWIsI1
MsbYVQWQ7Hr7eyNAdqN1tLZcye5cpMIuFCmwVWoTma8Eg7YfQ+Vz1hXyuWfU
NCRxdNcRqRTePoH42sK9f3rGG6pqX91hGcv2HVRCCPmhVxqQIpcDsEYmiIGx
0WiJOO9wFId7VhRe0KXPTJQamtADaOIiUsdI1TMnD7J83i9fW+V8kz1zT0LG
RdArMuZGwuOvEIyrzduRsaalIP+jYAGUFEfaM71d8BVLTJeTx5yOwHK1E9oG
dtWnJ70ICj2FNqqQSDN+mYkZ1EQ96jFt9UmCxe2oBAgQGwP+G05NEs/jfgby
fafNr+Q9Cdr4agn2nNhK7j8k+DW0Ug6Y2sLC6hIiRMvBJZKh0semdlpBFqHH
nMRC5i8EG7qYFpflrM9+7vb13cDKWx3VIBr/7Wakz81axkhGBsDB5smHAOhp
kafgA2bydw2ZUi1CnLj0p3RqR7YxKkK4ofrQH1a3AdThakkd4m8YwlpTFp45
ji0/nB1VbM3ygyvQaZKGl4Sw6jql/4Z5sAXMJ9tJ6AuOSDgeVNliwAK72cUD
YdlLaNO1ceWR5jQC1nH/PHqiNoPMbtun8SRF1fFDI16UknRdANUuHbO/selT
f85VJkRhjguK9gOd56QA/IyzmzBRHazNtOkeg0KsVdPjOv3Offh5isG6OuNm
wrWKMMzy9/+02GeWvoRVT7YIBsexcHPnlwcg9YBe9zzXyFC8LljMULTw940o
ODBZ8uqZpwTEc34hGfypVZwivctL/pHlDvA1WHnXG9eq9i/GNqZk1lkPKOVk
V7xp1z3nwDVOxF3kg58XBRLj04cUy8uYXZqn1+3DGoTpo1mBNWzF11biMG+h
qRRobBdKz90mh/80uIjQyy+4uA2c9XQTvHIs0BF42b1h6i5txnxQ0hNRUycp
vo4sof9RNABHtQAWebYFpV6KONaWjluAr+/4BoU8xAMExaIW6fJjfchRpZO0
mtAGskIeYAg7LOejrgQ8YH4/vRVl4PPLf2jnCiDEuow6RFd8uELnSB94uogb
bd7FGLQGYlR73nDLBZIgE0CHHnbkYkQzynuGWb7Tzaj6sSPyTATQf0MHW5zM
CP8sg0BcmBHgngdHJK3HdK1WWjpPPzeqTWPuQhtIrXE/iHdZPeRNF96ld1iH
hP1Vb08OMaNPCmVyRakcJPsIY2Z/j2A8P2XW3ZK3TTKlHSUc/flHnFeNCZHm
vy4j/mbCROZR+ph4nKx9ZUZUMMA5HLdSILrSNNWdgeemibi5xKXNOTslFw2G
/WpAx5ufrEs/EjZ7SL+qMVYRUXHDuYrllMuEpXPDW4Y50NX93mvAt6S32Zeb
B02NAEkRw8CPPQw64mCtWvtgj+wXPUHk7QFvmvCPtyAi1FrzlbPthibL/+8Z
49/8tFHw6fHWCr3EeUMhqV5pkC8PgqJ3kLH9/XdvKxxSdKx3Wn38l8WMAxnO
zoORxD3zI0CUVRPCoMjjKxE4wbUSmKNbfS8RRcrxB8Yh756hkslHQY49GeLo
Z6hlfeOaF5P4YDJ5Akpi17KxdowHtjufiR/9wqNKGtjNQS8AMQ7tp0SCDr3J
lzxrf/0tILX50ixVCcnI7G4elfR2EvETtVCmO9TEzeKwVGx0WAQmCMU4D4Yx
TS0ozSEAx2TPCsaXBgY+8SrnN37PesCuB27crZP7gGL2HwfX5rnL5Z76KXFR
tdo3JfMMtbosS0ymBYjTur0hO4zaU4vwzf7CvhPDyaygfN/SjKC3quKqGgBg
oO23HtiYzCjG+7DWgLK/ubaB6MJNpAyDfb7aMg5LO/14XRQUrPlXmar2HHkT
yh2qvNbDgyRMEXX7DNQ63hhfawQcOo6RfDW7RlvIYcuC6BGNWeSxRCSZIOfQ
ISDVG6BcBkmhJc7GHQ79Y71TwujepDn9fids688fSB5bcV7bJdeWSvMFhN/X
MYV67SbXdgaB7e29D+++NkbJ0euCdWP0y/8xV3APen2PteXOsq863JL0dxXj
n7+sRLUaIJ4dIzEmQgvgEFIImG2U6I70jeaGONWNF7iCMna+tuzJkKgTi+4n
5TFfgaDlXTJEUyxO+Yr6VHyc9OeyqPdOoTs5WCot6idmT+WTCY0ZJ5oAqsrX
r9jW6ECPmdhmWuHqgNzGL3aGTs982bY6FXMriUFodAwrlsglrE7zabMvRWCG
I7wHy8oFTQLFSd49zmW4W/3zLSityaPMqq5xsZoJkS2rii/eAnnapiRwhmDM
ByCBDEW13Lw3k9HJ0nfr+C1VOjcInn5ZgIt3PjPF/omv1mOiXJ8U3s0s4KAi
pkuTLxOoeypgVgM2XeXWYekv5s6ONfjS11p5dIMHdJqH0dxM85dLqgbxGipg
9SJoZiDaYm09lcfiKEEfme3jvsvbQsq7SOXpYloB1rA/PeLMRhg+qHceFqbZ
fjXJyFK8BSu8IRKfWu9h/mjJ8cv3AzYbhfVhwotTmd0RaQwDJkVABtk3LMOg
JJTQ4qcqBvXkwboynhepDY4pB636+85kiZ8ktaFkO9BbTrPRNq93GVcRcMoU
trpmZDznHpCjOPZ5F6tWbogFN/maNWcxleOD7f004/Ev/FfhkPVmABaYqwYg
JH3rSb0KrdICc354ma9ZRDtPA+lK6LLn9pK1hurZWC2YeoXGQVICbozaEYaN
YiI50J22Z8dL0WSIq7S68/ROokmUOLsR+eDsVFPe8d/pBFLyRT7/UkWGifYc
Fslte1MhDh6ZEYplqFj8gKDE+Jhoqu24SfSwX+6j8BQ0zv2QevBoIuQUWZUo
nAhIpeLxhnAuUKchwYFLUr5UCQYv5UOavlq8I9oXf3ZRkUXGgbZGqZdxcNiA
5Ozdc7H8+szNxCMsDNQqoPTXVA2oXm80mGvMNThhJwdH0MvS7dv5XaFBUAKc
YMVmLr3Qd/nbVePCYdh1Rz9fEd6aBpsr/mEv+/3mDJfUkwashcM79XknHxXB
mXCLQMk/3zD+mG09BNKvUCPor6LumCt9G2OAN55nZlpjKIIkFfX1hdfV8Q87
n9uwA/M5MgzG3/kUoU/XW4JhpRur9SXBcxO9Bac/8H6ScUzVLFKMbS1lrY4M
o4ti4iwqT/KRn4XIK67oXCU0YxDIw13PFO2ThPWHals5QjK3IwxBRR0vHJXG
i04NqicEzxZ+LKzkirauAM9eN8eed5P2eU+L15OoRmYW+4PynRwjFS35IfAH
PXWjw7UwRE8euSQ+nTH9gV/5uv4hmkTlMuW5+zTf60s0r9Bsm1cuV/Q8/ncd
UVkxwFdrcij1N3JIa2fJnhtFsXVp8D3rZ46ObWv+BNNsBDNdIH6HxxmJ5Vq4
19I0kxK+0Xlsqgm00C8SLAsdd/PnG4PsZBCcHsDCdzPX7P47F9VcAxU19lc3
R/ejf/G7ZOtOZ8uObH/0IxoX76pf1GQaO1gRMuYz1dcZlDlXs2LxAy5erH3+
WPat07jbRJtRrXR2d6f/Au3QMUMCUIxMq2CkWdjbeYuhSL04Q26oAFCVPciY
tAQDot9Kh0XXVGE3x7j0vIDjQjJTnS2anVNeaBUswiHr2APNTN6tJmR++oLU
tZtNf20KViYDpjR9/UB/rQkV+spP5vRB0JlxkqLxzPkTzcVbaF/mZlQgAOFv
rS9QkDS69Kao7JLZJmzXYZzZPonEbj0gJh1AuAv3dCmotIn5pz/3YNmMyBQC
BGadsNjIDVkKXcY8PATTqPkqFMlpiIsR7oov6C1sFAGeMcLgBpwTGt1yv5GX
KQKNDxOHLD2K4K8o09OaIqBiXWg3sOsQCO8zng/7VGI5ZveoxiYCMSyMjUVH
yQBKOK7Hzvn1QmHbgtq3MF89jCw/bVLMsN8H5MmuBS+7aGOl3KwRz9vaLGFm
yDJqHSEKwuIVtqjxSDcPh7V+Wv3S0Bj7Q3TTCc2Lx7oKOqmAzG8hCYtreRRw
LQeRoiU6br5N8oO2wSNeaaYPwBNRl8924754NtmEejG9yVGPuLWulaMdqcEO
USBuT91oxAQ3EUF47NJXOH4x4eYhxdMz8qStTNTfk2Tc8Pc83Xoiks4WKHtA
yEpSr0OBG7OALlCj8fcRGmtZHFFoj1Yo9P7QT4ppS9ldSuhnm9rjD8V8pdae
sT6vejC09fxY3GQdu+LxJ0vIX/IXe6BdYSgLjqUibrSpD/HxprwddyMC9oSP
yxvB3dX3ugbFDOIUTAWyv7sy3FRcBfgp2RyqjHMxn2pPaxPgVbvp4oYU8hVi
s+LrQ1xbj1vtAn/FGGFPoYFh1J9Woc0e/1AJYTeYpN1PcHnVb+maDQhiuKtl
iKiX7a7pJjskcFPpyhRqUNZgx5+1PZrR8C1uqH7B2nEMjBGRVfzrLvC19hlt
dXfNq+nTdBVwDPtbw2rsI4UkiYPmW3d/NUE7wO/tyehxloYbjf0TAA7+B9m3
fTNWVSHl34CY60mHSjXUyVYXabfj9k3V+WIcMiX3tTSiqOIZvXm7OE5Ig+oG
g0N/AysQUJT1+3WsWOmStwyJsUx81RBi/ciygVqdq0HyCH6ID7XL886XjDBX
g2giDPuQ+1MqiqMii9qsEcvrCyvRWI/aQjBms0jhIvsUlQ/AcBQWvv2I4o0j
tBbDgjzQqu3c94sdIgR5YOJdcHbGno3FbZ5i0dO7iJsM8tHtpdCNdzCR45W1
ug1VBhTU43MUSzXa9vrCUqv9/91f2zc+JCsCafasNLX3OPY71So0xmxlz0gz
aKu+fIfUw1+8Pz4MkrU/uz20/TvV1pQVqpef6jAu79UJ6UgogMy4RprJO4Vw
DEZ+k8th0ecvq6zOtqyW0iGUXIXfW2kFKhnvr0nAI2kGcXY36U5K1BohoI0i
/7HiF7yoHB554E73rTv3oqs0xz4aEb0kJp5xYOeQLJi9sI4TmmDNHD4hMcA5
Ys3KeLvfV+K/hlkp92b60zGf6kSbz34L1kf8fz/M1suhCleRx0/9SVigfG99
2aeI+15VHWamh3TZzPboQJylIR4Tvow8Zd5B1UW3zXHqBbSpRmjlZB/xOf3/
W8Xtzd716LD0udnRve0Y0M1oTzYTNuhqUKKCVj5UFmUpLwBJKV5JMBozUEMv
zgMFzEAotqnzNFwgWmOwa2Vroi8+BDfHT7qK5tY/VGlXmh6lsKta/xoAvlsi
4KGnfqeqQt0P/vg1U5XiB7uxVoVwm8GLSMUtGLo9snnq8VU0Z+3yVr7gyjge
ajuzRsTyYpylFMT6XO3hTJE8cj1/zjbLb68FjPsnbcIGExd0c1swEG1B8hCz
Cigd+zXL+08sNK6HKFSUm4PUnEv/8ao8kzm13db11IaY70W+/8+xCF4TctSL
JU0HDsdWKS863pvD2BKK/amMVdzQC3qetwuxeMOxXlFxhzXiVyFBnHUddtXt
SbSpqZnBFRSOxMJLGVr8O5SreijSXHtaMfEwhsjLsOdv9t5rvRlbrV0+yEej
YHO2nHu35vZIGe4FcHsIuAGc1hLRfhPXpXgW7gJ2ITi2eXuVIiG1yh1DVJal
//DgE/5zpWuGJiyBvZDi5RUS6wruNYkUS3zzRi0kqcc0HMiG7aX3Zi4w24no
GxQSY6QVsUxF86D22+8uLIOpkbqcIavK8EHeU9n26N28RglO7EvnumElmKBF
k0cdpfhnexHBj/ypF6gWnTcabn2xOeGwbPl0gGV34T8BzuXGp/hFWUr0v8gc
2NRCWUSt/zI4gCzjTOzTd9PqhhqcjrU6lHmhEp0egeE4dIkJ9iNJQDS3pAC3
bq1wTs0SrEnJzz7QbV6JDMvO+2jNDdRdDDFGKqE15df3QFNh0LA1Yo0ObJLK
O8X+6hsP1rYDJ3KY6QmCKprzrTd5YWWEEAPATyMEViv5NqelynTnI0Qzy5+o
n8VvqMj7DogLUegkzB5GkWst6Gn8WtV+9Js8Fa2OH7Vcz/lJ0Q2Ndh0m9Xwt
w5l6L9GBSGGC7tH+qdoG7MkNzu5/9wdBmNMV+VCP59mrjU+7qznWlqROro46
pqTGtPyTme7dSE/wvX19mWnKnyAOVk8XYI59dWq3r1P+0uc651XmW1MMgLKO
guBcduoclLUm6vQmnD2I+HU7wcGSJvNmrsjxDGT6hySwdZzBG9zLvj3Fetjz
/F4tJxkh6tp3w3h9dxR/t4fMwC0itUFL/HnZvRH0UjB9yHbaaybD3rLtMnsA
DbXbP8OxLiSj/fNwElZx56QHaPnHPdz9C054GCzqorAipfSUoFA3QzMPnjp7
TWJQPeZjUSTZVuUSHb42A4Sa37YMetbRn2/59CS1OB7w97AyOp48MQRv7kzf
Sj0cZujomo95CW/CQwJoRVR94UU9FM2vPKd029Q+P+bENNvYDUEUAKA8nK51
/XJAQvMidNT6lK/mw2pdyXMfEha3z1CLXOp7iJFPg4rrD59rO1medPn1olgw
9Xj/UZvYmnJ/JObBw1rxX90bBte2TAPzsbuoVffCGcKgNxRGPdIrz2oysJHT
EcKSDSV4iyrKqn3WhjhELMws4DKMeQB5yV2WigyNU4SHriehCqMEAdThCpSg
ySgXx6gc/6BH5Ox/zCtaOK/yBbJhla7lcCn4b1b5o4fQxgCcGHFr6MsVfTtR
YxBlXLhJZ8Dn63oFgteAlHrrJbzKjmRWqiThZ+lf1F8pL2bEAUgLZJraY+dd
vc3NtQnngLVDCJwdvJX7nF4XEaNvj26WVok/T3ib3Xvc5+TGdPlcJ5cRLv45
tSqSfWVMehwCOFdRmYX/ATiL6xzMqk4MtX4P5oEXGWb/Y237hno7Wb7kAH+j
w86LRuVv3WHq7l0HYu8gaCjKeTUC+pJ/ELaVrG4xfEVEwZ4o4iqDQWHhcmWc
7ttV9RrzlbUQocr3hdc78UVEXNrDnijZ4CVMzwlZExccylcc4hRbQC27w7OK
GhWDrM3vxp0hwVaGqYRkFuig20AvkBuAwIJJGW4rhU2XBwxkOlKPzTThwMVD
YwKoQllVI50/6zaHj3vPNCpj2gsWpia9vhb0bzCwAVb814NF6AlU9jnXLVDS
3Hgq3FHJO8+rNZzwNI9ciQWE/t6FAB5BZvaDGbYKzWehLtxMrrmc6l4066OT
O2Y7/0iwX1AKyc+YdrTwh/EC23jLjz9l0DKh4gUSs9kJUZYKHREicVCk8p4f
e+Exh8lSWhKpIxxqterWJy2jR0TbRpl/s7gg56uSpHycush96wobfrIqB0+v
zrZwMNohdfo7Y/pj73I3BhuMhdqAJkDP6Vcgbz+ChresaxD4QrpbfmPLo1Mx
uKpr/z+OjwdK22Lev8AoqFnUPd1Sp/LH6FBMWHE2VFmq0vTxQPFAHlZjjrQr
UivMHG2yx+Yzbwk6GXxYD612HplLhr2bAkeIBofa/Ps8me5i0WGqIPJUUpEs
ix477iF2+ysGtRJOkez9/0Xk4j75egDCZCGlEH+D5ZgK8Chwh4Sj9yy1hEz5
P11L82pec5FET1atUvgSNNpaalxi9lSuHO9hPWHnPPlfzbRIpjfuSiVsvYyP
j6fnZA4f2jLfLDOhcvpL9RnPXCdvimpuSpKhR0hXHRIzC0gayAdZ5Vvec1Lj
LfRis6KQeqeJboN1ekizXn1ZEad+Y5SbT2YWIS5mC3LAjtzBdd62Joc3dSRc
jPQtQ3o71ZuXyzJj/cpzvME3JBVq9PLPrDNDX3A+loEL44MaZkT2+l3pNdS3
CLF4hyV10z0uOsvohfbHMvbpfnAo/P6asI4Iq2bvYXM0YFp9lyzMk01t1A1M
zX/kI8NazUyKel/C6++gmSryYUnoI/BgSngaujwcs9G3bo1FRw0RJWz8IS5/
7CbXIAclK3QB8rrOjPUv8dENbxGGVGBPfAgK35Pgd3TwQWWNtGA4sL/Uhnps
2CsSap+WcuDQlK+METKvtyOqd1gYyLiKtM72BqlTgVe47hm+GdD2mxQu4K3T
EGXuV9KOFZcwpBLiLYIk3tIvoXWzXWK2Iz1SAlmFf+CGFWQ/Ocq2Y7zUzW2d
XX6oCltjqi8BHeeJODUDfK2sgKUxz0Hx8FStK3OTNcMHy27vSffBc1DVxZ5q
FQI1gu5cq5d9Gx2fY2+c++CQqDk807OLNP7NtR7VLyRCRxZutrETZTCilcDl
xCHxQZKnXTVg6/z0OtCXc1jxJp5GcnnGm45+iWxUSzLc5dCpHFgastQzA4W2
m0Q6C+kDMwVS1PZUWHuj2ZMmbfXvMoywLmRBtd/i+1TMyszy1NIm2N+T71rF
21xFdjxI6kXj5vs7Yy9Mwcak0Tsma3wDXJbN0m0Ecwr36XuHUdptHaoCotKG
YSqh1jgDXkJrvzirEKj0R6Fien7HGelNUfAWj0FRSfKVH2AKzF8qaIuIuWgx
NmDBbOm3DkFISh74r1qV/rIqgo3Q+nN+6h8+o+Q+xN0I8n/1Tq2foq0d2pGl
MabsOGDf+N0B4RgXEHferAUYrl5ps4AsTfa6Xannel9M7qsZa0tE9VF1BcIz
/YuZNBx7fmSGeR5/DKBknoqw51FLcPPm56jF8Lggm0oqDQNJYDI9E9eMBrw4
uA/qEcJXR9jbHhqUAWqUSal4NHXOWO5f2gLF+qJSLAJBpaGAWQaNQtPZLqOR
/YNP/V6KDQH4j6+VxfEaIe6o5Fa7Pp9yLLDRHZGEQMwmuHaDUgyQCDtBStg6
tx3C1iCvWZJaumExcA05wtuGH5te7EEqf1tnEqHhUYQDzuWhBGzxoNqa0Yp9
6C3ALwlI+rs5f+AxX6QCv8wTlW1Lsqsw4u2eAUdqV/74p3foOQkNMzQpc9fp
wl4uZbPTO+mrhPSWPpBsMA5eFzrQMtOc9VmkZNeHZexrnkvyeZSq0iUdgsqd
bSCgHb4TB2ts0vPb5BxaXwJomnea/OgRD9pqGgep1X4ktzyzhpwIqMp5b9fw
2uIlPAXbEM09BZ8J/jMeOwtu/YVpA3iDZwfLkc228KxjTNHKGP6LuZ7Y8Y2e
djznD7h7Jlp/yQI/MKXuhHTG4JOsMz7+VKChuzWQtsAx2Wum7TOfQ0Yg3T9R
wNpNXkBnFi1wSHsSJmaezrCGHf79EhlMn5mNfY4M066EKxnaUR3ik57pKq5w
3/pRKs1fGyUXz1mU9VUd/4yANnZls1FzRu81ZOwEXnVS8X+tYEtcCi79TSlU
XbxtQSn3ew8lH3VYziN2T6RmEPi/edgBtyg7Y+vO3rVjswKygnUvUoyo4kQY
R3odPh/L6wT6mZ6vJSOt38ckOOFZQCUXqBqNbsdA761aWBGIDUx0L3dqcFLz
npR9dGpWTMaQsQo4C6ZNKgwohYMHJJM0TE8VDMnyrGPLOgxH9AUBimA3pwM6
ku9QUH6eqgCWc9fFM061oH+Ne8lbRa61oADeLOSSXJnzSWCDRheSI6fYY8nt
O528z4lAQgNxDJCsCBIjKiM3/Jdn7UQaJ3igBf6guHNHtw77ZCmtUndvPt4c
H28IMvf5JCBN814qvNs4B3BmyzD74W4/ZwDp4uxnNZY1FU3m5YuNuZwTJx+U
1FSbzllVwImimMm/u/7PQP6ZWVYV06J5hKIXmP0IAIkrWDn3nEJ+csOTpBzj
IH31REbCayn1zCvhu9AvYI+47kQB0i8H4PIJqzMMZqDwShPsck0A+B1b7O1Z
thZEYeFEwnOPphtg2vMwHUKBzolI902PUBUWr4lFsPjlG+ajCbyUeOs2vD57
nYcQkCETo7xMPchZ4WQr2cHiYanBC4nQYHou7eQW9ywRawPFej2ansm2uXpO
uIPQnH69D/uou55AX3uCwKZQv/SpJ0J1HHiniWDerQqWOrIe0GcuJ0UlAvrb
69qxD9eyXGXkQyu98Z7AzUvRVZ/UICqWCDVPT4A/KcpU76WfjNiLrMmhAXT0
sXBKhKT6L/Plu45sEa4FAGaGvz1IF691amV8oqeuSVSU6nDZClfoTeQoMVvz
L7gq7t9KnRv+tG+d/eJ+NRyGJoR7MoXRpXBb4fYluqsVwDN5+FGR4eRdEJZO
NP+drqsec1VyZ+utCVE25C+FeuWvWoKLm3F5w5MVHiGx+CGlHkoI8Nq0YS16
kevr9/l8hfuGR/tfhF9lI28cYYmrl8X4r+L8suYh4OmPy0yvi32dhgw60Eu0
7olAfZsEngSifNuMf2fMfanKgZo+PxFphb142aFaQV1BhbfEkXGIN0uIcSH2
go2o2uUqq52DOGbH+bbGMmQJiQORqS68POLE8XE/jTLYYl+CavORUrGtEaWF
ZBotzwwpcnH+XoILWqEEbMkNpFwom5gcb/iTCPM1mXUdmqZtSWvqw/rBkgPm
KW6fDAiRIFjACI2XN2drNBc7T+XhsTvfx6KW0caXM0WZbLj12FV4SwhEohJP
FxrG4348J3TX514EYzaSkPHwvzit3rnjEPmYif9FX07+z4Z6RZqJ4axwsqJP
rrSZr5MVGct67mhh6fMBH+pnn5nY32NrapnJBGVpu+pRr/9xTLqqrAkacMzT
j3T0Lb+kxIAT/DTtHMcVvsBtcsCH0du5/k3BDN8ah/WLrlTkR5bsGmPOQPtT
FRrDm/itpTsYd5xSQOkyJsGbmvYsAJ98VOR9lxMCrF6EQ4/dQfA1gi4OpN2J
KFYeQeJZPMUQwlOK9zoMXJjsrXhAmSSvBLzrWKwMGh/6hd+J3E8AK97ZJzmA
u1RPkmY8+V5CFJMBlk96K0PyNJqrMSVge8NrPuJbAMv0HU5v2MAywOvemydt
MXUf06TqrX3+qsiy9VZrngk+G4VXfgfWfpnLkn/jWTX6cB7bjr8CxqJ7IpkT
uaOAF6xSCKSwodGF9Gu3zxgU38a5xq7ArtjisacRiRnGRamRM2ta4q4vOrxS
77I/5oSthJGQy/k1ZCmyKxxoW+91yjmMtoHRoWjPk0V8p+ftCSict1bTa+iK
jpWuSdJyJSGRb+YkXgrD3h62pndtZazaNobb404+jRd0KoWEoVpkZNJf948F
o/xR++iy6W2MGwujFKtmESjmFSY9tkN5U+qoWtmz51F0fk0OXGBAfT6p9ST9
kCaqxldnXLN9OIq/N+i0wqFRV5nSSG9K/Le/y7aB6OtVv42PvXjgYEd+yv+l
7BlOYYju/9ET4b8Uc6YyfNIxvdmRRuzBJ3TSHBXMs0qZcFMIBLEDbiT24I4K
f76A5Y57zrPnBew/Udo0GRZafqeZP1WfMqCMoNfTjl68/SPCzNy6a6ktbZXN
jUmZW3vhUueGmBVIcMienjD/aIF3j9exSUt4VQDW16hhgCWNr9SgOb3Q1pwb
tnWBpk80prnwsL46cg1f9o3AQnjVYEVkc+ryxjLo4LcW7r2i9SLRUsdxd1Jl
dmYfY0and7Zoeb43iYIiQnK216Oq1qFm/5eunzM/usm+bu2tjY6AvLBocJPB
QeWboJ8Q5WY5BOmR1Gcld3uBlKdovbGZfdbk582iVTXUWRJAHgWUKPeQxZh2
EcCCSLXj0vTOv4EakGLlirEItRnWDn52pCTXA+HGpQimvT5qrhR0voN4Mjj9
nhfJ+fev0GiZxeSU9Aj/DMPbq8//xC4ic6bT9cY+nNhhk4NB/qRiH6rUE3PB
2YhQUraB6Km7jJpfxm+DnHSQkM7B9/BIT+9F6hiylApHpgqdXr2a6em5CTYM
4hA0hkPOyy9PrFt/bLK0t/Du5t5E53AlZqMEvqPVtFlfGFoFrnhmR9/r9Op1
gJqAmqFkpA7m0oFkjYrUQVyzYf961KDbZEJ3oP5QjjKm1+yt8vSfx3Uekr40
jxXXdHRleceWsjDdR5otkfH6ToN7OdEqOiXKupthV/lZCthiV+Ym1/78UXID
Yfanpxvx3wFzdJExErp2d4p0vBYv1dGvNoYsK7StJtImzD1cIS2KNTrua/wn
lsFYfQ7HnfyG0cbZ+z+1W0ARg0monDgzb1PwHjBhHQ56G1uKHhF/aITrR/wi
lT/d9QlAmyJH3fqT0FpXxOTnWyS8an2/8794FQxAHXsfR73v+MqttyrvmOkg
UPIlcU0ceD5z+siEY4bQYPC3FzEQ6Rfi3WeEXccTfDToD4ZqbQt6sxDaKnRh
ISFPCyMzEJhQ4OzJ4j4FgwCi7j24pDZ3qBbrQRlQw4g2MDhSJA2HegSW8wtL
I3vOLDO4W3Qtf/TdfjoqoZ3mlyHe5COO/JdIVFeowriq9EzUbbAwNQy78qE8
wpBtJlvvFpYMvB0HbsunWAvk8fdnYVQGZmhJri4UsBRTIrKD6AFgVN79Y1rT
gSwoqBprYJBXzCddWbTzxqNcZ/2PVFqxGHvmK7OOG4Cy8ulRqG2QyDIe4GSm
FOYpIy/DYAtfXdYdlgjOSq1Pa4vR1fdY0dX0AHBJeamAsRdQMri8UmHxj6WR
KW4KM3kwwaVjxWYGY2erhwyh7aO4qWU8BE521l4LANVZ1HwVyR9CgRMghWnK
ayq2U19NcLnEU4sSv7YYE0qRKfAMapaP2mKThrmPqOCVHRcc7RfZagiMdvvX
YwULgmbmnTe4YI2faDPd71KDTWA1W/l/GoTIJI9H6TGJRtVONkpgKkcrUioS
FWzgXW9o5nkxTGNdxQ/1uAllEd2b6vPAa3+EoG159wCqCx2hevHMRsHLTrVY
5CnpA2FQhAMuJQzQ7+U9oBzqgqevfagPO82QP9VkbnBumUW9yTy/gpctEk7+
f7R48UAo2eCJqdYIstoqUpclvTY3v6TtQM0zk7f3HkvTkHsG6ZcP1JcWNwmh
6HbNw1UCu+XNuF7Fpl5k9l4akeymsvPCrrqtXY6k07OYI1Z7JJE0Un4T/J9w
dnhvbuZh//P2QW7W7DypE/3xayZA/bcXgWidvL52glXykGrnRo88z8ZRa/Iz
Y9qSz1bszNKltfpATJGOynvx4XLYGdozcOG+nT9bVUsrBNLdih+gN4OqlRsp
0oMK4QvIg/1rw5ZOsa3E50+AOYxzR1+/VIPOnF0R71eoGj0+iulNdXpTVvC4
t34WeCT3yuHMy9v7A3Kyd1+PlzyH/GNJzk3dL+2fB8esERDyj/x0w6HiRBZo
+WG8A4kXJrcNxrCygVEctJdPO3ZBppjysecXyPcOq6BU3EFGARg046iA879r
nE7Ot+S6pJBUdwBZAuwfp3rkMJuj50TtAXVw5qaIfttGkcvv6TzPrpj1+j8C
6JCthdrDIF/Vqi/XLGSQjG6uxEx5uZ2bsfV9tzM6fwRixBh7H/1SCZjCJhWT
T2IBret2mCvmR64+Lxklt8d19Z5cVBREnJdsTlcBkvsVEVNSxiMiwk5MNw3U
Bui6wAqPkXqt0JSbBr9nNUtotcqBFWm2rReN8bSCccs/TIV46Nqzzi8Ql6k0
omri5Iv64e73s3q6+QvjGM3GUamihFf2/r/tnCnlbiDhkG0jcuIPJKrhDua3
laUk0CHOIdkK56hAx6cJK87Tv1ixk5sgxic4/GPe5TToWPb8PBlIOe4Xr5RQ
TsQQd2xJgdlMFKCWzZUUp00HRoCZtZ/rPpF+LlWk3tyjQbMx/Fz6DCBbzn2F
BqTEVGkqUR0fd3cdRCZdipXuzeADeyZHTCY78oXLaUB7OgIsGduIGeRj7eyr
PZAwbeUdCx5UaWtb0JtYgJpOCxwnyNYyWlEUiJobKd4ZkhTZXrKzSPoSv6J5
Jn/Cd71bntsGS52Eb8MQvzjZZySgpFM0dsV7Z+H8uN+14f+34BhJf1R3Dgui
dJyKl6NKR+QHCtdzrPAFQaQivdq3FaaKZX2bXRlqddLAIpXlq07KrVF9CZj5
PC+zUpqv13gXHmkB7J5xwZjfFX15JKb3P/02u19VkyKL6ygnPpaTOGBAkNMx
jlle1uBaI1umTEg5maLRBLb2Hy+cWwa6cyNLTBUvssqK13CJf/+LnRbxbPes
fw/M0b2df5Wp8GFngFit4g7etN/iCbwL3k3IH8oo6NkGC8Zs21ddw1r86kMR
3KSNxpEJsUeV7AOAp91AaDhi7hqz5uTY4kNymRrtbTwGYRnCyoLJtMuTe81e
n0rxdJliPStdLbNiecvq7+zn0Wk8Zhy+ntdPLhJ/ncm5gFMmMnRp6uetAoSM
HkjAbrrCeLtSQAgG09t5Anlf4z6+Yu+GbRjoHKgMhjJ82Hg1jCE3W4xIhzTR
M7qW9hUXfOkVm8AQXQxE1laKSuEu306/UrD3YzuvML1D1MTERwy/A07UlodA
rSqkWHdJam6Oo7VZEmjx2eEoN3P9GpFnHmgluEWHbopImreweomTramSQTtt
etdxNpFL49pTDs7obuKB9vi8Tes9OZXSmwsjwYCrU223BCGmt3fqg0MGD0uF
9LeGmqvpoWIZI7JyIfHvSxmXQco4YbGGq/x/NYt0m/KCNOzCQK1S98fgwmTP
wzsOQRKgCd6z5QdZBw3/RP6ZTovRsfSOY/QrsdtPKw85ALexBZWaxnxCWLSc
7ozvfbYubziawNCzV4JbwI3dLl1mhZRk0QBBMw6f7kIQ1URgAhXZm95xQWV+
k8BU2in+KeR9hLgCe3/HWtbVIIuTLCnN89OMQpMY0cj+tobkp6kFgbC5hbLK
XWVM/CAN9Taj1w1DpZyjfk2zkUo4rGkFq1HEhshziOUxhdv/C741gpEESmX1
zSpm/Ky7xG21WPaMvzj7J1YcQA+fvWCfMxcLdNcpVGilaa/DX/YIM/E1Rkgn
SJ7p4bchloe7YD1TunJwwT66hpQqmoExwDvxg7i2kYUp1OmcHpFhvlm8H4dy
Qwmn2GIleYDXQZPwYPyDZliwDkjQj75g/LZI6doorGYJrEWiRY2zKkHHfhOY
0whABrz784Z0Ymlw3GTnv9sNG00XEPsF4h3I64yIoC8XYvRGO4pZ9igu4A76
ujkX2K1IGzaDxb3FNFeUMtcznGbzb5HSz3rA5zDutdVI6Xfjng0EA4MhjHmZ
njEGtDeDwW+zsIFCwjW35dNF/AJMOM63pWYBGnNqExcdplzsIlbvTodtYT8P
ptCyOqeNo4xb4vgRm8ltUF3gDXlfHmVeHOo7efHAKeOoxfD9iOFxcUBQEHDv
T0PRMLihKkOHcud7EhC+kaTbOxCkOKTJSttKqcAFRYSjF5DvARyWe8pHwmvI
wJy1YTXZvGry1C98kw5aAnBTK/Vluew9okeu/NfXzXkfAo421XU2BiM/+/Zd
nzC0jjS+vWkVQMqznqFjLFsrX2b0NpptFmo7DRk7Iyv8K2H2LtjSSU5KBLJS
I0wylqQOpqr11iji35D1LYPAh6AgDEExyGQt7goRtbOGETuzVfCIrfPMRmxM
iv81mNO3e6iUIqB6XqcB+QJUG62p4kpsB+wRsf7qGBqn/EOrAtmSyoDvpNhF
MkjMSDpQ5iCftoxhGqfP/ZvZClu47x9tzMsZrMQHieArdFoi1sQbplRxSpGk
74Jv4nWAacIgLvPOji/k928ut3gdZ3LgHkBRV9kCqiUEMGQJKfmje8r0VZem
kvBApZtUapMPPxK9fNgxWVQ+WmkUzKexiRyN50xsDntIAFAaF/e9zacbDATI
vaU7Y8bKN7RmKwwW8XSB+8sucEcbhixqsSHJCqg9svXTlGwYonEifE4EZqr1
bUxl6y5XVGqU8coS9xVVu/YreumE8+ZKP6+EANnN1WwXfBU2Y2drz0mYUXOx
ZrfYZNo80Ij84gaEvcw+DMa7g/X8pDspQxOzL6TecmDf+MWg7CcJIzFkkp6r
Nm9j5Db+RSWEloHoIonu/0v3GqEAhWLnf3CEDV6QgCGhspKrObOM3TaPxQLg
leqhwsWVf2zuh/VutbMN4f+gFaFyLd9s9wPLgF/LnnJ6TZsTTSb08bTDZfKo
etk0iOOnrTOpkg4RPnFP3RZSPk72AhKPmXEywb53fiOEa25ei+Z8lkP86QGW
mOVmixj65ECqQXCM1M3zT2+XI3lMtRvUxtw31vUD66XQkDALZKF+UUOjYV95
YD1ZxTARmtRNu/XKU3nucflgu5EZEiexkHo8YSjoHHY2oHKe3MVg/1IgKi+q
qdNN7Fak+YCtFOZ9mV+MOzhJAMZDIRS8INUcwrffobWfBe/rfL4SNMu3ZE0c
CPkf6ALz+U3YgUIt78VdV7G25f00eOohWnnJT6irwtVyimNcJK8wloe99zZb
ExfUbUJtgqmbrBbUe916ivj49pa/8PsKH9st8lcUhZbNBJAbbr5hAfVDAgT2
KeRIYxxwK3gxqeXpUqT7fRIr/rXaervRIdfDkU2xp71opTdEUPn0N78KkdYE
HIf/ze3Mgnyq0ZjSb6cBAv2bSgwVR+IMw/DfXy/1Aa+CQeua4mHALNp0L+/E
nsjdi6Pe1EEd5mAYpegm0Pkzv/0pWG11dGGudgLvY16aV7yg6JG7qlxm5fCn
B6G6nDmZvFO7RyFlrQt2MapeUp3R5SuA2xfH/JFVen7fQ2knrJ1YWqD8UxwS
Dn9sPMucuZFFlRlPi0umuCMJougwfA25AaU0uvE3xXtbxStNCC1jIJ85P8JE
4enl2cIZxW3gwy/VgocJWdK+srZGi7uW3Ow6nMzhvvyrpp1Rqz7QG1OjbZnE
GvQ+74OOgPk2KyO/NhSmmlTq592vspcHkfR96uIo0OJCjv2inFmN2AGIXYZr
4YaEypKGC6sN8MeGh0r2aVJJBtE5TCq1JLk4dtRmqLl9fyNRcDphg/nM/XSe
h5XpMkiPwgrU6cczmBPVE8DfJSDYDovydvOerjp1acGp30PwKjxhMkVORqfg
mhsC90ql0k87H01r6t9XmlcdTiLf33q9JtTIAkp9LAxyYPmRfmAIKN88lqQN
+FU39yIfSa0Tk2HHoju5zIOf/NGwAoRjeSRd8CmXJHESV0yl++ZluwyP62NM
kZ8HmE71TQ34zvvWH4FpjUMYk5Ktr2JSl6gJzGFl5jhCCQ3+w+gybcYRyfhi
lzJ24LlIqF7U9ggnjWqs2gt61RE0ac1GJ3ln9gyx2RppEEzfE7qrB2uS3wQH
v2NyrDyoSh4en9YzfrnxM1VFPHMLJpk5Ore+1YDpBxO5S/+C17CEDZumQUiB
bNcYxtO8A6yLXmW1bb+9M6GfPWv1ApXQC38Oun+XSbt6QvQkc7Dj/aNOBMzZ
Z96crrIIFhZil2E7sQJZYp4KO4aCOKJfVjFkebfBfQg2SfIH4ttkSGzIFZi8
Vz4rP3oPiFxcvD3/dwMwoAazNqLuvjCaVLxci3KmqO6QwVYYptjk23y1z6WN
H6DWoSbS9U1Jyt7TmkHzKOs1/h7kIMEKkuFlwxZDeuSbgppIzlVt2z7InhVd
WVMWU+9g94wb1VpVtLjaO/szSbmxa+kQ0ZpYTACpU536l7XUv0Ym0O5/yBHH
oYihUwl9T52UpE7FpKKRD2FtarkmY0h1OGzE1HceV19eNYxe9liYulEccPxf
agO2rhlzpcskdv9iq/V8fY/qEeLw/S92WkVuQyZavnKMD4UaVIb7MKE5sYKE
J1K6xDqxpHXxldwGaK6c757jOuIQ5mWys90EycHNEmU9Ltu+7zTZS+2dsDkp
2Z7lKkgxjgAIFTCNUDKum373w6NZtQSAUrHQsTOx1lXFst+ur8wlFRIZv8RJ
4bsaM+63H8WL82l1sDpKiL9ORgfM3iB0bUKwOPMP7mR0LZ9o2FApOz5Pldfr
0H2N8ln/jEr1VgqhKiuFskh4NgMwKXQSxXoX9flkNbPeqZvGsjmdUmioj3lZ
I6XhGk3zK4Jikgx+4ylH+HWJ8VlpIzkteZf2B0j/vdgDNXbf/v3VK866cD9e
Xfb9AEJVNRHQSMiqfqPtx3LsZcz0ox842r2sqnzEsGnVwFe+qepllXtZekIB
T542hbnD6giYFj7icp+0h2FfG8kx4nHalGBkztzoe+guXvi2aa/dpYY2mxoX
06PR1AJysZ94cdc16Nk0iS7zdexWGtQwB14iqJcvwYiRAmB/w5L7Vj5A0Tzg
zW6xom4QanQTGn9HwxiCm8Mzzg/V6zJXBR57HBSwEqbaZiHHzoJXOhgqm4nh
9c/5Kq5h4FJWygExnQyQYB7jRA78Bt33ulfSFksv5nZt3cCqUjASJhM9jrhy
yOo3TMaV9GJnD+qpP6XTVKVmhETGh6h/8AkzqaSsOU04laIFY1a0KFiCdf2O
sABMF0yOuTJWAlOsxsY/lqfLsWaMUxD9RwAQfE23O2iD9FJmFRYkL79Z/4VR
2n10vSr9u/DKVibaC+OFMcWFq2tZRXdE5thkloIoa/c6zrypqn7HEx67bT4A
GOkXl+GvxdrOXPJhdsLmDPT409+NQtx0Ac6q0SmdhKUU/grmJbU8ml017te6
DkRQsa//FEaze7PSBAaux7iiVFCsQQrH37ccPJl4HF8OE/PyDEHcER8wpB/5
VPvRtKhKepezcT730FFBKMQgEVmpLl9dpsuWOwFDLO4iF4TUa4QZsjyTc51b
xXHe6Qv6PIveQkXvMryBEBoDdub3Mfq8BSUGTn/h5Cpx3ty1u16waAYuLWTq
Bm0vkBDVXjueuYzBrDXJRyGQ6A1x/CElcLIJsJuhd2Rr8MNNQ7x+2cqlmjRj
J31DxyFOTNv8QBVttzTSi3kAFyNELsQvy9kufOcnVic4FF4f4s8KxDCKLqzF
0JNnf1cq9VHoViroUv68/D0QLwrSZ7+aYdZrd+bAK8eR+d9rIZyM/oeoQnfp
m+BGJ9z4se54vp4YZAPdVOrY9vm7NpZnHfaI7WBHR/kycpIHu5PesIHCJAMU
Tn5Rr9osZRy64yd5iWW/ausd5c8OezzbhJbKkjzYXtEGJ6lFSvkzmbI+qj8o
yN1vzapMPFNlRhdqGmQ7BziTU6/W9JDYFokhmxEAIlg2mSqBqvbNqpFl1CCp
GYFzGAq9r8ITSmPzuH8X8YO7IukyNkC3CSq/waX8i3Bj0kVpkljdugo3Ctja
7/rWUJjVo2d6MTZN5aA/4fsb273U55q67vXOj2c9a5gR2GjB1zRmvvyj3Xt0
5SH/KOVtSadw6VLZfFGVNYymLLYGeMyAiTQ6npoxm51QPmHdNUbIpdW2MPY6
zBGfQetAPDeUGw/Bzud92GDxbP0bnyB310xAMrxDe5FJNK4K3wzJfTAXS72N
dbNm3bCkEmibN0zGdKNrd1QISkbW/8qoFArnAjK1lfOuGsDcxm54FGLRpPDs
Jg4P9j84+wLOgcAuzn/57DUn+RsNh8IA7rojeJR8IewbO3Oq1BoQ5s+XQ1sB
8S+VIXreYHf0f776jaR3K8AOHnRKeB0OxyeMTSq+et8ETOVg3UM1dFoOsTrw
0arBM0KbY5VTYQOKjxfOXXSpP7Fk6rYiRp7S1qxIYU1U5w82ECnT5PnKzpQI
Tt0YIHl3EGQXs628X0dvoSU2QyCjEasGmcWzs46uUrMB4h/s8Ff3tGEHZmTo
u2sfWTP0cm6vC6p9297NT9GZcTmoGv6KZkwSDynOH0k7rLRzi7mg+MMcDSu9
Arn6RpAvcMRDlj45fX/ANl6kaO1RN0kzed+UpzRJaPXA1n8bKcfCI7oghqe4
WDnYC+kvNTLgBI3IjlpuK42dHN78Cf469SqAlYCbCxnX1gYDkQPqMf6NhYUl
qvT5wsaORL4MuLKvSmTTwj+lScY24q8xvZeKs8r9wNgSXcJyZHDEuoRCB8DV
oIVkjKBXhjiXZFBoGdWtZMefzzL0d61WilerPgSchs8NHmbRMmDu2TcMl2Fn
WbBLPnHkJ2Vgx4Bm9TL8Mb/HErRLdEMeWaBLo83enck2sNmRuGRdQoLMj6IJ
pCSxGnM7N21eM/BXMSqBLUcABL0tletMViZXLMPmPYBw+CPiB09J+9JpPdop
1msNm9FK6tBWp/1c6rmVUQzDLDW1LwXqQukfR/6k6Lflo3N+e8IYDkVgCOAO
7PGKEhGzRVO/KCz7axwjycjvei6HS2oIC7Y0OqJM5PEaFerVYqrfqeYhcSvu
qtocwgNg9K+h2WtiUUyYj0OQEe4YQkawEM4U+MpUClUUun8gJ4yoog+wjAOk
IVkDz3OcrSm42jdlT7sDT2XCCzXZg7lFOSMfeHDoHtwkYmEvwf1pPGfgLG0X
yy8FZcPLvtDyEpc345cNsQZ5afxWnAKRdbFhLgphc/VPbK9RoqlTWhSnEuzT
u3D/C600PA88Xf6SvxlwNLmzUtrGwzrkRKEDB8JUtQ5fViZHRDfTi0ATzx0s
GmcvzGLKnq8BhRqJjgfCJboPWWGjddtTFp1WbqawKE/v3pxA0VvsXblNhJFR
7iI/x1PaqJKSSYrC9RZqiYJu1WrlNlD5PTPaAvaM6JEWfJMCrrcFZalyoEze
ZkXg4a4RYh89z3A6sRl+QsRBlE6zUrXpz7qD4o3kCQH9eNbH8RBMftQ1IB1t
uEjD/G4rMatEL3LBQwAo6u62hw0U1i2ZAbVGZs5cBe5cyqiyaka1MMolMfSA
Ip4wrRfWK4CwpWieSNaL2fNvixXysIGbABfkishKa836mel/wCS9xkttufqU
nwbo0IO3RffBq5b8AhSFVefE7Sig5BakebhAOIJOJjPMg+ERuXByI8J9qFTK
pUyuLoKALv4ATSjSYrYKPpZ60W1aYzvnmrvBU660hMWLxjdzOYBlbK2tLOhl
UGLKEZGFgsrQfIT6LbwpSknARnoDnclbm5RkosuqK661r3CLIt9mTT5O6Por
+HYaJwVjSIYl2lvpg1AXzHrMEL9xlGqkO9pVxYWmagmephr3YYyMIfO2rv/P
Vzh0Ru7JFR7jaIsJFw3YDCn3OF+cjcfBM5pQTcWuGleLhnHSBY38V4FV5IzP
TMZwayiazGROxDxVQ3MWEe1j5QHH2tKOQ/TcgA/o81Er0vY6OWAnxy2pO8mt
dzCB80fPz5nXELvZ/5bxlhtWNEmvdW8lvqYwyK+8fL6q1bvWYhzjfMtIT/WX
qNBZuJlO97dUtLEp+E3G8hVzMjF0YNYbxMleIjRbCzxMDB0+ONBbH8lvem7F
qHC4y1z3uFthOEPEtc9UJtzxUez3UL2WNjexd1+XJWyxP2zD3vJwGDO2o6DV
eqvuTRy8VDSHaQkv055/e/TV1Kwkg5iTBxu3JmS2HYYyUXnGcw+hw1kmEnms
vSk7342T9nAtbP/iIMZ+4UjgBmTNsAhl/wX7Y3Xjx7WylMH/qp+1IwP7Zmpw
iLotMTarBuu0bQGM3sXq06neKLapAB0gYB1nBtRAhSJTcO+35EGAZdzBpOBp
1PkOGrDNPdHo2zWk8H1uRnlO1LBqkq6VrZuX+wKFAh2spQkgwK8NloZOvk+9
8XJul9GBSdJPdJF2Bdv1nQB4PJsYphmzdBN68LXKqrlHGlX4dy1C5lUZbeBw
Mf8oMBEvOVDqAn4WBISgoZ8e28Eyh/lvIQ74Gn+FbQiDm5dUH94QLp7ewaDn
CIroVtnnkVB9xQdDX4YL30BGNnD8mOOV/KeK73EYvTd+Zh54PqvfBCwXymwF
3kjAjicrMLOs+XjQ4Cehoxwg6xFNoTVdE/AfTNWsgohRkok+f8L38z457g7d
uRnQo/10nDjp11q8nfjSxt8uefmIVHUzjafMpF9K+R3ZuWp4Z7wcGw7h/aIe
DC+m0JqjYgMJgDXZLP9hR49F5HxsUPapyXPgqooaJh+T2QgXfBAMxJmXUlNE
3nAppzYp9K//eRcSm7U42jf+M9LPD+/t2evUCGWQrcTsK6jdy9EY1MLjcqlD
ifB+RkzesaL3WU+VuelMQl3BOwvKpcNreZEvka9LqFcnOfX6MfqHPpVuS/1d
jbDm+i2krxNN/gtRfSz+BrF39jW7nAj/3qY9VjwhHA0JzhpkSUmC56XQzwzd
KYdMb7sGNI9RzVwGxhDYG8Tl31YfkgOHkc41f2wfR2r/JJA9d3zdRJBfqJB3
DUTmpwljF3O3nH30aYF429gugYna0r3+DsXBaSrQ0Pl1316o4kBS7YGQGFzh
x90oYPHL+mXDlnyFTr36wfJPFunXdM7nw5KNq9566okPVyXiKi44Ww0i1xNO
6V0KY+ZBCSYmsMYXLQ650g1twp03YRCB3GQy14SA373R8eE2qfb0+ciUqpt9
h+dHt9ergs2lthZg3id7TNacBOUyjRK9MeYpqXdKt4Hb4DfmajBsccewsh9l
qu6JhCdxaY0ElRKEk87TOYduhRGuA82/YAqY4edyQrG585OJli9rDi5PraJ1
bsgh3ASeQ0zhrIZjLd/HR8e3GNxDABW+Ib5nrazMZskCU6AZAX2TPTFVgjx8
shj+xG4xsb/jXh4hWPmozozVzRcMqleT2JQtH3PA3NIWr2bhZCy5nqFNCinl
eBc8+CAX+OdjYz8ypiVb7Xc5wiFrh+XUCNsW/HFpbq/vF/VBkJRG8VaMVZYd
+gQxQBLTq+COqqV1jijR4om1QhkIsgX4NXeBin3ZTQC1rcO/nH6pEELodesf
ZE5c3odIovNHvVkwjnPR+ISEh3EU28Gvnntz/EEUoFw99ryOX4K+zF125eD1
bT7YsxUEH5hYytcHdxHUvDYHkSjnMuWaBWiQrYqWkHhJ4CIn0C8v2oj4j+SF
bqmbKxxOV+qen7BtMn4vzUnbCE8Vob1G2K1NxOrHd90jeZZhaLEYahU1ha7/
yrpfX96Z48OblA6xONhqib94O8o3SIQCXrdZw0oTrHo1xbpk5xYhAOAwlXe2
VDCF9WQlx0XDTQUnp0L8d/Ci7zyC1nqRrFtO7HPmrzECHyJ3hjn5DsaTNJFr
ZNKKjI2lBnDepKwpH65iu3lPJbDtqYsCLC5jpqXRvff2d8zjdpp4xsKhTM/T
RPssOs1G3D/md6ooF2/Dba3HV9nGmSbHpZtpiNXT76JrIZSqxYay3q/GbE22
8GKujn3J1pQZxWLYW2LXVUTgjDe/SjVh83APl/Dx+hMyZOQehiUYHVGG7fAG
/EnfxMQ5OATRYiItTkr8fvB+8VbW7E/WHXQSSDo5KsyN5orhST7qWInJwdlD
q13LeLy5bO3wlQdgjDq8A2sI/UAp5VYD17yfs9YOPEGn/9fAuYA93vH1OTgZ
27UMJca0ma05l5DTLLQZYQSodo5+mNbiTo60WfSZLX58crJmsRx8Gjc4oHFd
QLAU7v6kB5bKBFYFH1cadnoUXxAHjG+TB+mdsBLw+Wb3xIkoNKjMhlbLcMZX
6FqUBL9IYt0AglgGgzbS/X7ZehKNap7ausVgHXIgZgSgaKlwtRcgqo7uX/04
ugqJ1VjbzmQ2qPRXvjXDwFKGifT8WAaRsv4u+z74pT9Wuh9P/8cVl50EFAif
XAftFKY9tlgYsmUy2SX7oXR5gFWR0DsRC/8rnKJpgCIyInGaxWPDxkpzwvBh
P0rRoFUWfQsz6E/JL9/J/zMUw4Za9pQAMYAs4A1dk7nHTuQRdXlNp/2uqwVE
MIkuEGS/t30UvPdJo+uLYbMgscRv7PA8hdQWq4YfPFf5hb7s2FlBGAaFXbZG
tYtlP096LJCt49JBLzs5FkuW1rxD0fM+MaOi1qdPIdu3VsQ9MaeBQIJ7OAwH
N5r0e2GKZfs7YODTf0+U4unKP5z+NO0L52i3E/2n3B/PutGLg7fIE/Lnq5PZ
8fGgCCukkU5d79K+3w5wDuyjcRVD7LuKMvT0BkZLklWiUplU/gQfO/j533nP
3H7qg+i2yq9YgNHAWpcqKEwVhkFpVnSBvb7ooU7P2HDNXtNyqAFRFFMn/G5/
04F37NoveronlZTNm+xw4ldZXW2sdPUt6dAlqTxlPTwIZpDZ3jfApmGdCrqb
WnQyJ2MhvQFgc1YlUkXD9kM0K7e4IBBFuLADG9pTVmZYm3zrw8mDJbZbZdbp
yjOIEdsIAoI6bQZpSogdKG814gCRes+SDRW3FoGjMrhnY9yXI9ZWrbTZl788
pgUU+OdvrlHBL94oRPt11FzLUzRV91lehOCugkhCDYcdI6IHapJJtXM+RMEn
GtlFEu9+G6wkdRWiS2ftZ2C7vbrXj91+WB3/5k0DSOaGWI7plQToU/SvHDZh
tkcPiX1GWKjLHOMOQmV6WWdiTp2yICLG/MlWuw0hqPUMu1rtGYLwbDvEywZC
RXZGT95PPNemXfU1vJV6YJRL7JjU0yNN4M1lO1a2N0QgNI7k21/lh/dohK5X
nw5CK3HWrKsuexQKxXiSbUEkVZQoi5zV/VJV/FdaXEeIg8DYi9r9/oaqdCvm
hku5r+CcmqGVxhPe2N4v+fO1ra+Psj+cUguPDblNhxo3adOeOZyQaP6ddAcw
ijo03km/bDmILE20Mv0JFmCM2D8ub/G5RxNy/PGwJH4fNPQK2FwfMxghwWK1
E/eckfGLOAYNCyWb63Vfmuid9oGqqlVYRqhpPOGATq8+xIb1Dw9HqlTEdA5c
JUylYAxl7CZpU2nqfEHKmMzB/w67f7sch46VmDofooxjjueSXn7Fseu0r9ln
KwNl/5hlLTWBvP/qBI7PVgjgGjQkbXQqwCuBTItc1yGMYeT5OSr/U6WHoURb
GWusiocx89oyqKjXDl3+ri9/zht2sc0hDXQftpxp+ifcXTtkFJO1TKXDm+4H
3jEIA6YMz58/aAwWzeHAAlXyAwL1eEdT0h8S1bUUoEOPe3AIBEWaqSZARta2
EOZXz7maX467HVHNFE3xU2NER9G34TQk/nNl36Cxf4+9oZAKB753F6pHAO+/
ggfuZx54nIE0Q+T2HxYwfNCnUcdDkBAAQEPcXsV7UwYjRTIk1Q+mQYQsIbv8
gC8kbfrv32lSjgdvP23FkzdS+bXuc7cww0eMiWvVlCtGkFJ9bZfrW96TVgE7
8c4RKHmdXf0XbUdEu8eWXfbWkqGUis9y0O5Aa27qEpWL6N6Nzi6SGh+pJtNg
SYXd5xEt9LQIk0xzZZD5s/lmtS4lYjcf+zNtmtObEr9k0pUr1y/ZbpsLQoco
ztBgqhbrMvroxLLDR9EhXRDslVml94fGzILahamXGlG2Rfk8KPEgcFfBn9dz
Cth4ZJJs+RaFSPHGF8ZRoGsZUiZMp+AnQMOeHSfQjpzeiYunPueOJkSvo0kD
9uw3rW0nbh8dtHqQigaKZIp0Qe+2dju3PpL2npKeC/6GJI9UQrbrTBEYLgeR
FxKqZs4dsmLMtdq/7npD4DnzwDsiR3bEW+55R3y+tl4AijVp8dHtmDDufgJf
WmPqnvz9X0Wev3FkcMGGM3k1xWbclr/ETYnLaikVLNkwJsKPqhNZuaosxM/z
arsoseIwHC205Rv6nqhc5E0smPrmpdHC1+ltFfgvWiqNT1FgyYvTZr675gqT
zOfDH0exob7KALmHOk9lcrzZEOcz7Ja9N1bTxEMgHYLWc2LTwqS9yZm/+oX/
MYUrseA5bdpifP5voYey4hllhnVwhdaodcoHD4bXRZ+6ljjJ65zGbDF60b+J
KAeQUSVV+6yA0GCMM9PxxPWj4ZlFxnzqRdTBdNgABlyNzacOE5p8FqYB6wgD
JnHnVAFNn1HCJfxI9r4xn8NJoY4jhprfXHsBCfjP6eonrJ3qNpSSecpS8FOp
NMR6xMFxZonATmUQ4eaHT6LgIXzmsvOGB2q707m0ATVYVIWaFA80z2yw9kXU
9lgxVipDT9CjPOM/rLFLOK7hWyMwbWXwHqu1oCgPtHcCTUszb66ksq9WKPal
N1ZSj90+xONNfBYYVhwx/kLzxX28cx6SyTFmxIxkqdEwPJNGFnlaYyIvHhH1
ck7bchXjqZ2TPgjQJJn3gApsF0yNSX3lKHqwBF9JC5qqrvzM+39JIcCSlfqN
pZj0IH9xqNWxRqw981IAFJICHNwq0lukFDsXz5hA2vfDWQTyPuqCQIUWKPRO
maahqC2NJrCwTbJqyjGJqFoQYemJpscP3mgRtZjzzsxhfdITly5eVWcY8cOy
DM4EhSceXm6i3c/3cFGhiTnuxdqk4zzVlA5ohEfFURLETErEPc2955c5i/YQ
VD5Xb9mePsOEaxHn2P3YHifct2AsKB+tqExEzb5V5Dwb7Rl9ECbSXsFxqDux
1KFuhDPyZGLhmM5dmwUWyzYLSAxbuXl3icMnaKQKl8epCcMhd9YTA/2twcsn
WiDzkqen56vRRlmRmZhH/0/HhXgem+nmx8xNrnuMxJnbVWSCcTT63tX04DCH
MaGCiF8Cs/18jUgBDEMzmMpHMW7UatmyXKiTZ4vSWhnO+dRJiTNe7BV8/HAo
6XgxM8gbSWDO5eMIfFy3/DEZrSXE3RLjMuGi4LhveNYkTQqJLo7m+z77mJe7
WxlT8nFVfS6xgEO/IPFCURaMS9Bih1T6Ohwm2pbOaySzgFB4kznRmlPswARG
slbhfbemLhcy9jkcZcRUD7AdxMvVxVAy+FQZKxbJzCnRajUNCf0rjk6ftRxa
OhcsdvENVmgsIJNkawyr94JfWrGehiUQNHaqF7T5UMWxtfW0x+WkclA0KmI+
sm9VhbdR87ursgPp4wb8F+TRSX1Dzn6hgFexk7kmDaFkNffJBaJSSCET3rFO
q2lx/aN/HWLYswDNd3qi9D+m5f1iK2EDcRMuYwOgxtR2Eft9hqL/4vdYmGsA
LZxCrFooMLteICwy0k7TY4651BJTldH3lIQMv26wTKTLfh7q+iRqC4C0jltx
LiwSVg3PQoOnpEH5VhT9p4M/WZrlMUJVE7YbOvBY4JZV/JqszaPt4NKADpn9
pMuGvn+UyW/xybZFhtAy+ucQJYvs0h+0owVrPbKGAbbJWuj8k5ahIjdvkW1H
vwiPOMtlE474rbL9j/gdnhIoGEKqrMlFDBa6ewOB8IMvpb1vPkc7H0eJx60x
QUWP9zDkioJ/Fj4ZkvmHNxc9lJW86t1qRJ60Tb7UvB1Y/Wz7y5/GS8wmnFgU
67aKxmKUrnCtIpP7ktLMTmaBDmCArOZF22038DB+KaJfce15KsshY9txH4EI
3wWOwVec2w+G5VqX0ju+P/MhdFWp9Pc60VsfATx2qRaObwoa8nsv9qtvVGJp
4ngL+PJojSl7hE2jEY6I9yuDiiRPDn0aaro5zQ4Vpmtv8ePOVxcs3Q5oWbl5
r5R+iVRx6/RkVLjQBthWnZFsCCeNpCN7bWIVANFS1xx52TWWZFnaxPrBrcbu
fcPFLnsO8c7Yii4BuDcd4TfA8O+dHrDTFSuyhmfXMiJ9kGOtW2NCybvdCctV
fDJrhv/cv2TZpz2jho8UlTQQDOdbEFoTnkyV9DIIdrZw+eJI4PTPFzijnuEe
5/vuAIw88SD6LLqLUS1hjW02waQ7JgmaRtJSnzN/OOx7uHyiIXOmaJDY0E7Q
olQ1txiZvNs4ooGs8OMgvqDPbG7TA3r+bF9PwUVHoCIPZ/rXvz680ReHl/I4
17pklLVOJtyZobs+VMysURwXSg2SWnDY6NU6uk/AshSpL+1oicGHUXhX+8Yr
JwrSruYE15EQEZR2loRnU5Qj3afjkmV+yryP3UajQqABAUMb03UYIwDnofLf
L8ohZBrMQtelozTSpjAPPNEcsN1Csmkf0+7Cw6eKTDJegPfxOXQFD+IGBpv1
OaXNA/dbzs9PRZdZrn/DNSjW6KpMojcqPXccjmMQkyswUfmWtLGn/h900AKQ
CWK4Fd5GAHk6q9vJDhZwQxBQuKxISFvCUsSWvIEDURupDdUo4xRlAJ/q8kY4
YVepz+RtehKiSDsZqXHTXJ/3wLCfmA6J/X9ZlXZ928aSGHyswhOsgiNbYrcJ
Pop16wGTL3vVdnEvoy9HI7tlggNg/n3s/u9TrgBPozjL/exVNlm56djtAT22
6mjlO3gUS5Ukj4fGAV5HdA81kN17pVuLiZpdYq3+uICNCAWs+D+ftA1wv3ln
uA6QR4VCU1NZB1S0/kdwpoCpo/vWgXfuUjpvs6LmP0dIuMvdlC+ESWDAd8wg
CsuKKqQ/WwbIMQpq5pKaot9zscXcQbB6XHpwm5qqD0dzQW7thGxVuHRP5IGn
sRliTmomXZeTtXXUpSyWApr/IjGFQ+SsftBakvKDhRpwRNUVV2sWiKwW5cWo
hbWpv3RRnYyfXFx8LEEa7NKQvh+7T5AFCwvWQFtGhbZlEZXkA812FT7mFYIR
2jnBuJCglkaF9nu2SVDEwhnuKviLBqrWmGFSXdalIxKXRHHAyqLSMM4uPoTO
gBmgIRIvConoYiQ+DS0S3MPJaQ7vfempOoP7cUKLZoFufDLrgd9klHYl3Puk
zQq7nthvZM189oad3FYQgkAvwX4D+ybmXdVtxsFQ3rS2YaNT54BmbYKNeRu+
4QRo93wZiZHJybs8Clgwc1nQRQL6gAH3ZN1262HY5LTKm1OnSPn0KXLQiKRc
5fD6TQYx9X8Y9LrjAJy/4OdXgy2NGVljxk+gYxcIzRA58cCqT1XhLx+fBTm1
bn+yVf6doluuPL7mcWapj+jYrZP+NTtGvu5RdHZyv7E0lSnmpdjZMsSdCaG/
j5o1EhlTxfv3PNWKuSf1De0rGAEvAhwfmYdxxAyB0IeVRLu0LIE5hSVbIKPX
ncqRgTPi4WsrS/sKQ/J5K32LfslcB+x6m6Yjqc50KqmaqR/ne/rpPBOWE4vf
LpscYsXijuTFRT62OgjW0M6e3Vwhefnlo2xK+D92wvQJun/MD+yqh2E5xYIW
mRmnYzJNBXnBDEw/MklnyCpz4dRrHlJw4x1EKaSpjYLcjzl7q4x5kV9BNMnX
CI7kUmdXOfWLGnHwceZtkMxmgCFcAfY5HswZ8K6MCeUwvotHf4C2e8To1l/W
vUYdE5QlV1tuLE6mSpvdZI7Vyx4c65d3r+uqUBmLI2DO6PmHKhInYIcm9Jrj
zTpcrdGMlXqODUNgGgbAKrn98pkdND4gjNtY7uEU4Pc1+F3n8k4vNdPf2g0R
4xkIeYLoYgPPBLuxPzX/U83B4ne8+WIMzfvFGLq1hsN5oaikPu064PSIKyEc
CnCfPnIEjVq6JyNMsS+hAqlt/7WD1iPu3gpRiSDT6TqUebSo0sh/nOeLopEC
WMerEENgl3diFfKbMhdxxZRKKo7UfTV/kTpPPjv84ducUUd3fEDyF5XOePUB
AHIIm/HlxQdrT83HRuaAW/5AWJqpRGZ5e4ePTnQpbfOK1/mf7gR+0Dm6z5Vh
SpRN9tUm/VRbWjqrh8q5VyJoj5ynYTy6Vhk7My6Vreu/abf/TO7R/uqPCDAn
XoXw36uZS4YppB5pg+LpaZoxQ+hqegj/YuoXRyh9MYPNo5j7QfMbXzLh/QB9
CxDzZtucS4fdmjLk23Q8tW+SmONsuihWnV1seWPzTwG5I3DaSsJN+no2nX9Q
7su5nLiYmL8XK+uJpYp3WWz16udhW2/eXEIIreRyZhDXYsfR7zLHWo3FM5cn
x6SUuy6vCmZ/Oe4gs/VJgSH/5eFggqAncy47oRfw3ghnJewS2iW3Ok8j2WuT
zmOTW/osY7lAjxT+cqVHoegXiwvMHwfoZ+svSdt5upgjGiZfvg7b9jQS+VAy
S44xnKEVO7xyGSQlbouN9+lGahcWghW2fnsV2DlzH3inoiCeLVtez7i0NglC
v51M2U/uwoRIzshw70Dl8CUpuH6Yp7r181UemJVTMJXp0cb7zYpzMulcx05A
jVhBXBj90xFla7OiWClmu77I5nUKuy1h0CUkeLrNEUw+9JK/vDqWeCFf2pGU
woGBXEbGBN2J3rC0SkIOXpxUzf+PMGvtUFbHHRP0rjhcB9IA62IjxWz/++Oh
ggnheI9k3CjaYVUmntc+vKh9W8wHkjgQeUznf/DCMTZ1QiaZwYvipvOf50uM
wjkGe5S2B/AwywxRtSYDGbDA72k7AquhwTAUHfNOQourWoHZW8mDw5B4ruEq
0k0MrvKWjLSP20hiBiVRlqhaFwHesXcO2DHtZyNrTtrUpDXdxZrh2gXi3+7H
qLnuIOAJoFYvyO/Nw4UTm7Ls8OIItCcLdV041TjYQDK5mYmK8MOE0wOhsPTp
PBgw9oqV9aTfTysn0aFOTstWbxUDJaJfy2TJSJfj509rpjSnEfsDNEYLndRX
7TbVqq9U0+VVF1cgM7umRyFXGwYJzv8hjY53zakgKeH3+W/hbOiwJ1uz4HVb
kCWS/fOe6hdfZCDSe66vscWpWu0rS3o4fxsBhOKuEoQ38rfuZIhpze+utKn6
8G9iRJSd3okutVaFDIJiyFgxh79d9fmTqOgQBXzKGM4g2PGBUw0W9qrmNUsI
NSkOXmHTz+5chTLhhcWfpxw/TTwEg42OynEKP2wi58SKG9wkNIAHhnOpATjq
S67Ddm2CcRtqSTPoBhC4DHnwhQljeqd9joCtzgsLoVM7go6oI8ppw7iOxE9h
+ZLlnkc3orAprwkSn0coHvmKhMAm5QdWaCTkhU1288IQK9ju5CxdEqBGHrM9
tSarvmQ5BIZ0AlvkTihOsPzdfp9CLZhC+kisNLGZfDZGM42KfEXLVDvMec3e
TNCkNIABCIjwOr6CXYXhadIXWK9bEdhEjpN66he/RHsQCrrLW1BrKzX+5eu5
EgYIttqkBG23SypcW6oRpB23kymGDDI5qbQ6epxBBgL067PkWpP8knL/qfPI
f8P4Y6hy+nJrNvMzjp9bFtoCtUSsG/VXnCajROwZxHvEvwj6sjtJRAZUsYjs
Q9GdQE/8F0Iednu6KxDqPh8VkOeF9XC4S7wYpI+1qcQd63AL94tg+msM711/
kAnoMSx+GnwYKoTvXcgz8joYQ0ZBXVNW+yN4T5bEJyJ/rgOUjb1jH4QGYR9n
umUjs9+plrfWO06gchoJvQJ9cotUz7ERuJ83IrtBFCu/S3UVX9RoAYcdMhEd
efr7dqER52eywSol3UkEeiHNTzlUDt9hw5u95MXC6i6WtCYy2xNvojYWv83F
+nBX1J8RvWTYQEZ2Q7dT3lkoPRxbNiDB2SccGSRrfOWVaUAFYN23tCmglUwV
+uNV1GS6mrCmoDD2ZnVpgMK0lu3ljlGuDpNfzAklAVd7XFyuiemXOc5zCKQc
6cwqe9t8CznNsjlNBl6lNE4vxFjRU9fZM1lQ+BlXdBLd4RzKzVCY4SL4oJQ9
KN65CeouhH2K1nXXh39ZMTvGNfeRocsQ19Ovikj/pF7NkK71UyONxytqRk3w
IChfEiR4qxRs2rLiiM31vhcxY0tWnx3LKk/m3kvGOCEmYL/R+WPA/wlTEePz
Sms7FUGZAFmxYEAdd+ycgJUjax77vs/bROaU3lHiNICObT3uUeVpRoo8g4Ea
KnJFhsOpZrvgHDFSXA7vtAw74Q1FEsx0T46GOulwEooBvZfQJj92OQNQfr3b
/xPXmczBniOf9Fb/ae/gj6sBrujuKTv8I3i0DDYpfje8bxQ3iq70Es3n4BU7
xh+PPlx8NVGg1To7L1QNpEEbmMndgMA05zJrI3EQeiRPcL2dSES9WEFBEV02
XbYKl9stk8PPro7Ct8zooHrLhMvPkzTVDg+4ZDKmcnt0EWgajRr1AqBS/V92
QhK0U3WVFlFzfaUmLBn746KqvmU1zsfZ64f19b83OQ6Kcc5dU1hB5Ki7xJtk
VjqIP+AJ/gEMaFs1At4gVxlAz1qRfqipUcfVlF5/XWwpWVvUwdUtEfcqKx2d
1xyLzAUzMnaPMLbaChc1pi5bt4Mppa927JrMZtcwt1tGtjjMJoRCiMoQFSLo
1ZFxn7lj+b1rNKBibU2tEKDBuEex3ZoZk2WGQg6j0Hd6l9nshT2FeZEHn2mS
of1jCbhDZwxuzF5kMZsz4LDVLw4T4ujj1QGE4gm+5SFeHhIg9owJQMuicHYa
0kWHOwFNpM1Jfph83a1Pl7GCgHuchWo62h6K7mEdix3WWiVoKOXkuYd4Dh+h
qj+IBZ5tg6cQvY6HWiQ/uMbfGe/M1gxJeAHuNJBkPgIOy5RqAL5DDYWla53B
vkWKEoJEV9LvBBRYDqWc3HF6/x733lu/2o86S/ZX1XisjAJWX0D7IGQ+NBb0
idD0FRfydmUf1q9olGVu/IviiikRk7sqdoOWemIJir4hbzRyXcAHFUrF7fTr
VQ1lk+ugzl3fl+lQ9WmAFVC0sw5gMel4rUAYmTCvJG1qrClLzb9u4bSafHzi
up4UtiU0wBexx4M93Uzbqou0dNcG9iCH1M+K4af2iW/lqfebAMMfnwjaxbqX
JEbEybdAx+epDFcpsHeyg/QkOTaV89qoyWrlmyEBxBZsB2S7zUexe8gHnNzJ
0GjKqkW35jFkYjyPtSLPb9OT9CltJN9tDkhmDbH2NZmQF0uZFRKXcSf/h5rP
/uS7Nn/IFC57O17/QqCJIapmcOBdW6q/Bo4cMBtpn0XulCvlDWMRXuUgAGCd
MoiDIZIZHnxJbRWoxcPOoYjv1P5dFzIALjzDf54pAAToRFq8w66uZuTIol6v
cDZQ1pMCDix61CrONFznBtQBU/H4Y1cbdKsnqi32jHQNaL11k3U+tkf0V81O
6icqDR0ykm1iH8JXt7DJDvHCmyNL4mV4dEvXFD37etzEdQWd+vnHLeq2IO6I
N2nIME5VA08WCOvsPVo8FgrrLOn0R7u/1UOvxckX3M7OGn+nXWq5DGvOgBNs
pDhrU18/lOhuYCMlHsUb7cGJkbAv364c3uSqBBSOlrGbp06lHXmcixOJ0d/t
FD6sOje3ayNU95Nnn8BcW+m+7th3ObQD+Y2kppCqnycWCXYslWjpihnvq620
NScCF7AsLyZbEoAe3fHDa01RjkYOkXYuYx0TA4TCDxMXNEnoJuZreT8goGCv
aTJdRp6jeztqzYFEN+4sJeqIF738S5k+ySmxkeebbKCY7oRQuwILGLBy3Q8r
E8lMHRTAiKzPkQLNm9nf0eubKLjZNaHCNfJoABCKJmPlhiEParj9Ihn3oxmx
tL0CcrBmHnYyAWPiPFd5HZMPc5V6GkNB6GSHRqBbwMAgQHCzSLSrShfB2MXD
dlTNbxyfnOdmdJppa40n038BiBhjUGxcuJ0RqlhEnfRuAFUDFQ8E80kOSPfb
p/1ioWVCCe0Tf9k1B5wggiT3zYErTtDspMAhHqGdho4enKqXTu/LkIWnLh5c
XoeJMQtkAbodepvsPqQgQePEj6SwAdo3RjMcp4X20WwvO0lzjU6iOv2IqqZw
TrAXq3iNVhsd1j9ioIJcd0C0cO/SpG7zr+idT6rpNlAa61ONPzNPBB04q4mZ
pxs/8AVP4UOeVlXmYU2ww9fj5VRy7T08R6ZqQoQGKuv+Z0Z9pXD1ZgWXQdZW
TWSIEcSo3FJzixqRXyfuO6II1qN3Ia/bqBj1Y4qYlFGLboR7N8nM7OO/MjDq
KRSaGE5mrSqM9BBdIaud/UbpdytSbnx/VaDmEFsc/LBtBdgl7jccvWRPFeQx
oXrhs1GaXpNyXLZzZIyQBCDQjVA5Anixh2sdCNt4FOmTt2k+3H6o9IrI9n30
qkXt4rX5RYydl204iCkp033a/VndOnq+/RakVXbnec8+770935VR6AGBFfoI
ZdLNMNwlp0x5v40hvGZBkUTvCFMp1mP+VW3TmU7P6zSWNtI7NKG3juvYkMGy
8ug5+bZWTtAUHeIgREcJvEY8oi0kxcgMFhXhWyw304KJc3vrqAxsOwpdFWaD
rtOM/gDZ47eJcM36f/A3nZDPOjXt8FkcZH+9BYGe0OK5aJmcJQEJbu4L5cuc
TVAqUM8Kjyg9ufilidkjDsiT5bE9M27RtZYnUrKF1qStK7QeOqjS4k6zjm4y
eZxZIY+DmJO/oOAgb6cJhb5H3OAbtmAKnoTlqE5EIxURRFk//ck34ynsjshy
tb5rvgJ/bknRFG8W6Pd4x/XkFwSQuOVdbRy8cWC3x5eLUC6gtFTfngpR348C
3UmuC/KZ8IO3lHb08ySYKR5D6bzQsSXOo1dI4VBJUcXIYr3WULPKrUx4XxO5
WvqMvu+qAJZjgwenqCDI3p4twJdd3xTXy+iXqAV39O0xAHSDj+hqIe1Y5KeU
5H3UvnhtR0azufOQ3VwVBQslyKDodwOt6kEtvj1GtaBpe34duYpFde8CRI4V
LTU0iaPGW4A4H0WzWx42RJ8QoKp9ESfnGyYs2mFsNrHBdC9csIliTfIiFxyb
D76xYUxhhIWvK3dLHeznUae2QVniwhAnmxQkTosm4HpPpQvzpxJKfmKfv3q8
rMoxbNA2eWnL70efxUZHyytwo+4AGV+YnGFSdhEKvfnRcjEkoLmr6OX3hhg4
o/nA2GHvw8rXyBlF6rvBckf2bcaChCF+mUkDlXCiLp8IMJ4SGxXwntD5F70x
JTQx9yU2QXa/wb6WtxnjeXcaRMS5s2dOdI48eegWYlC4lNWUy9xTrZ6ZGHex
Uk7vU8YBkyTQmMEyLG5OPBVGgaHlewsbaA4rqDWXKTdXJKt3+4xaKmx+Ljj8
97yOeyqI4yzlrzlU3PPfs8bVWMq4PYQdixwGgd6YlpkuYHvvD11RHbjjZ8Lc
VKKyleCdNbFsiL4WHgBwGimcEl2VH1TFOYhxznhcK1AjvG9/a2Shogbs/abG
0MtZ9EQZhMazSnFGPxOo8/ETTTLPLoRUPMBL2uRbUD6gFB3DmouNeWZDrwto
8LyFY4tYJ2au7q3LSNW+GLBSas9T6u8pPrJk88oAOxpa90C1gYBzujjJ3XV1
jQz74MUWiGm4f5WRBM4PPwFBm5s3yA9M/D0TEaUoaCkBhqkKuDT3bXt9/6Mc
wDaYNjqPvOOUdgOGMwE0ivkjibdfaX0TEWFGIB/337A/SO9jghwwCX5mggyQ
QNHCkVY3jUWY13F7JDOkH/SK9BvETYwbm5ZC12tTZJ0hETkkgDsmdl5CsJLl
Uk004HLuoC8UKhG/nNWKWABv9zRujksLbS9tb7i1j+wQHS2CCbfDwiUbiDcz
1p7HYaqYBs+YQfwCLeQJzvdvt9WSu89PzVZatdRuxs+OOcewjGWNdxBPpMdW
DIWo1K84znCaIGAAgFYSbJUvoEPhFNHEaDjXg0pVhpgEHnx6S6+KHzk3tnzj
6BLa4UIc8HLuMq09BV/aV8nNXtaX77fgBEnG1d4/2WZYjtOHwtu5PaUlQHtZ
FK6uDDN21FIx2CGSOVu9PJxYsnLkkJTVQo0mchB6m/jRn/t4gLjnc9knR9wX
F9+A4PvSRr3y2aIW8/LhWG12zcJxsnsVxuE10fIsHN4juT3JGk4eyC+++PlL
5JUazu8qhsFfsNLLELXoLHwpoUz8wWp9qW6KOOAfYCNAB6O1SpqSMjOj2oHX
DpH+k0lpE4qXzdRxMtqFUVDLEND3DDkv2+nPdwNeLSR/k9ALZr3eDwPp3Scx
RlLygXeh/N/0AIgoGaXI/Gka/Qg5nA9uK8Zm9yQhXFcnU1zi7ZinsMJUvBCm
beBivCxVhVHxHJzgEHMv/JADFIoqn8Sw5DLd4Iwed10/QPzqJ40tOaL/2yR2
cY5KxFx+OQNZapS0+29QRloCsOn88xdfjFCuf6M6ToK1tlxgI+I90KcWweXK
3ab0YUbGQYUD4I05GvEFvddoRCBX5PylRlKY1Kp8O+BRE7PNcvToljhW+R0k
1fl4ZPWA4R6JtqVdRohxATxncVoeOeN1nGm2n3oGFHdL5xgw0P15BW6KWQdr
SxsEWxBD4R5Pbh5OjhDAmn11stlpbwrLasAgpnTlB6cOiGtW29bqdcbkEJty
q1d2xKlR156idRNuO9VuZ+6xf/nHJ5Ots67FFhitZN9qsilx9J6qog2Eg+if
f2izh5orsgBqsCF9+O/PdF+LWH4jA2w59Fww6xryIG+PAw5+PYwOPtHJ+A1V
64wcd0AuRW6qMDFphMJg/y74v/0L8yWPjKlqD5MICNHEIOjQzj8UcBH138XQ
6Nas8oGjnof/eeNN4Lz0jtYKwnzhmznkGUAUbLwB3k2yCJyxt8+gO+VsVxVW
0HQfWNdRDu7rR3L8V2C/k2PgZvdRSyyVSkFx+rPA+y6hPG60ndIJlfE2U+8S
nH3z+uINbz7Z3dhxhzFpQ+X6USdeYRQ124InRd86Bpd+qZjaNeVCRCwaDsy4
49xtoCLnC/Egj5ndESGVHc3eGMfa4YYQHenwn7modnM5qvKE2K7bnXPR1PkW
o9bx+Rs7OLhwHOq5kCEMjE0lRXCMq/rGto+6/dklEiWx/eXaeb+2YjZczEzn
mjmLmavzQnXJRls9FR9//DXIhcK0QuHx4Pz++fGcVXrONu1T6ygixUA7Cxfl
A5JxPPnLg1T3MiuXk2uue8g7AkgIbbWra6Pb/0ktlLXcPiVxAjAtiBVidfS0
zBBH4yp36zXr2hfgqOZ1mNmiAmfqbFhPoPrPSPsg8+Ey/ALH9ekn6yWH0EoJ
qkNZ7crqVB6ND3GzkBulufLpxS8BwYG8xXlMz6roBv/37PALVh5UF3OdWSU2
ter6c1geYxiZ3DmlFbSUOv/yeE5BzAKP9ImDy7kvF7GXFgvLH/i5kGD37f9t
G9r1fuG/HkqFiaTc4EwJ4ntJY7HyGMHso/qt7BPmBpSW5KnIbe/huelCUH4f
MMk8NndjebECzRDZrHZyEbODnbZTQTOpGKNvElKpsb8ztp1HjyvEKeQ4rIKo
/z31Yp40v5ofQRpeLPkZggMoRhK00yqF4kLuf0jOgXx8suX6AJe7+WUUmmwv
Z4LKqyce4XmBxRvhudfCOZePys2p9iI7aIioT8mUem/gu0ugzPvPfc2wTgBJ
shnNvShKSvUev5xOQrhnehYYrvW/CPiHstQiP6m/Bk14oMGy7b/S+JW3FVi+
NticsWj3xoaz9D1QMfsCUmFN0xwbpCrQFRW5HfJtOEmLuxSCwDfy6megctb5
YsSb8D0VejOKzMF15EPN9n1YulNs7KlsftbJPaAF8F7TIMEF1+LmHUgZcKlP
ombELsotrnQChLtGzcq1/yhPbGB9k8i9BMSmq/v1jWcKe4VEqeQdt41jiLtR
VlcgeYwPzxuxaKFoH+yBwrnp0kJ5dTuA9/r/7yeRStPmuHaHmqMMiQSyc6re
Og3kSpa6eewmV4XdBGywA7bo+r2QRaB28Wtmuw+YpCIzrJZtYdrud+VpI1K7
4q33oClS+fjn38hCsAS4HFQULOL1OBgm/W5MaV63/5aS/PrXxaZbp/BLWrdN
XMRUO1L1cCAoXVS9LLX7GdpD1NbCalXw9JGBdEh8UACow42L6IIMRps083Gv
pdElF+25d9GTPCCyypd9E5308jg72pfDWCMQqLlWC+3ZtZO1CEmhGJqJqzIt
2VPHeLYWoDJKWjQCSUntJR//1L6hetEyTxRpj3ElCZGSTeb1Q18TeT7VjfBO
KIwnBDT10smad2pxCUhX5y3TnZqPhgjQ/x05m87lMJilZP67q8jFtqh7vciX
K7Jw/lkjdoo9WKFns8W3Mi5NcsCyzCdfKcR2K8N7eUzOs0TIEE42bbt8eklk
otq0l+pbLwcx8qGkKjIjFzyIV/9Wn0Sj2ywBYD9aL7+jy1O4A4Fz1Sfqr/YS
z2M1CQWegKJc9ORtcrJTZnpDdYqbGkn4F8AuFZejsVwiV0d9lmxa5hdoMS9U
42LqzzpJcXVUAN2hWSTkswPpDtpZcCRWycP/QHqhzSicofZZfZ6HSHYUd/ny
Vmh1S3OOf1YX6cpo7p7UeCnMoaz5dhv7W3KYWkFBkP8l84I469Ny5PgS+XYs
fGUHUJ4iC1YBQk0SlbhTZ4BDMBgkoFn0ACV31/zyNXU0lcYZKPf4XgIaG+Hl
wXVHPT/jFEMFqRfgWIlU2ojeYfE5bbGbpSWASgbzTz0VJh7lc0FSlvJKRzoS
HYbAbl+tJmlDkq7BOZQc3l/b3hsrCXh3NH6ZD9lVxVDF982v71PH73qaR1aM
iiu5R3I6P/OxUFGGeZEplvCE/rvTENO9wN9tT6X4+mgxMWWYeTfehbKDEmB5
cyU7ZkssUSwE2RrwD8eVwxa7vMzg4QfCfpsdfb8wEdHcfm3L0FAZ07KP5mgl
oXAQRP/TOIAx9JS0ZgetvR750zfYBCD9TZdKFPYbAsujXHKNYHQIHueKE8ve
Sdl8UP8QZOfysL0HLt5vNhNfWZtUSGjEaJGJyBnKoQP/JtNr829DXv8r9rtA
39OQsUNS5CqgI6HWYa5+7snItFO9S3gqH6HtnIvUlCcMhHn7FDzlD38allav
XNomiPtbdaAuGZAnta8vE++fOPBKiflU4jtmieakkPKaCpQZZhNlJq72gzLa
Mc/iwcUirhWlkee2qjrChxE/Rweed20YbNpEkGZ6Z/29tPWOcyhO3DMQ+WQv
vrknjNL6PJF8K2odL3KIy1lKCr0pwZiHn6GoEjDHiwDer1M1TGbjsUBl6LyN
3MwpY8svUrmQD/3vLPWmaEhF2VvHtpjuhhn38EmylRD6YurKeUuc/0oCIt8E
5LbjWWCPnOOuoKWaMMqGY1VrrXkwk2LNIBBCPgGsmS9eel4kl/rONH0EAnQ7
t0/ZkPxsZ+H96KLzlEZCEeDOF8/eMBO+Llmc0fw/wFTQbe5TypnwNbprlSVQ
uW3daQrVXK/DdUA2e6+j1V9QCb1wvuUCs3fV9wV1Kw1BZVWIXiTCgypKpqfV
60LqszM/lnnDu1qfPOHDyeXDFmigaNPzaoxL1zr9a6/MGJSc+Ju6deyDsIn5
fyIUeVwtM+ZPIBhdCD+CMso+gHOQ10Y5wJNfxY2U0mnaZvnTerf59UUEO/E7
qMaawo9FlH0ZmN0S70YkDimY4wwdOyKbgwJIFVxB+Y6KtRl1RBRClO+PxJ8I
uuIBFVxKFn73L1sA8oHfo8UMKdovWdNbI0b/5CKSMzoKT+ecgD+Z/p3/wR9B
CE6DOE/rEIjocT94Cs/1SUIV4JzXIHu6P0FeoXJl46fyvmgM5mN8UKgL2++Q
zcyY+edRe/+a65lcLBibhS78Q0rT7eumoK2BBrFYs/x7jx5cpiD6z3xDcilY
WHP9Kyuit3p6xHjfm4QFOJHAg+zajpfXBe6O7ablRYXvvU0UlBhJ7qilGUVX
m08sDQU319FQWDq33fBWwAvzXOw7s/20yLoGWXUPOWOnY0vA1CL4TCaYOr4V
8m4lQBOLFFwujzDpXF6KBxG3BIcgmigPkBgI0jz8aImmOkzFx4VaxC36ehsT
Sgb48PMEvwnykN9UoU4jy2mgKnhQPTpsQtXmkIb7MwypSc+9WMCSefPozLTI
9x3TK23efPwm4kR9GovjdNwgAmKpf7uOlP33KWUbQXRWcrR8cC2Gc8wRA3yA
n00MKO2iwOzqEbI1iIOM/k9jRQW5Ie+n8i6TrI2GYEoKRg30jYcgTGB04sk3
9stlavFFaGs7m1FIPNqYQ8E/3TvJX3ciCXRGNakh4a3DoKSEru2nQL5UhmfA
zAspiYe+a/RkD5H0OavQ/lPc79M7eO8sfYl0d3UbSYtHZpkC2Hb129XvHRMC
oxTg9rgR3i+taCcLVbLyH2z7yRX0lNpVMe26nHkLybheQpP/PshHLSL5zizj
rqoSuEgU86UalPKCd0zuHT0NBkMSBgfT3vNvhapMIHvTtwSW41UTXTxUPLxP
4tbzZF9AyZEYmSmwnwEITxPnQWkFHe/AtdLvg1xf+Cgl8PgJmCrzAb46W50F
pIdCticWo1vh1DlpQsHhpGxiPrHUODBqkqkNLEfpBu6MP7bCVR+eQ2Q/ZW+0
ApvqnYjhDJe0tTC6rmMQgNBQUsncvRt9LQyk0obay/mBqSQ9MfaZFL0a95ZJ
hZu9C3AnaMAPLhIeSflOxN+VQrfacaAcumHnWGQR3z1bS1kSin/Y+e8Cevvu
3KZLs2hbyMlc5IouBjImbZx7NOEzyHWORHDkF05lUwD6dz0dsvPTme3rtJgS
m2a7V1AYvHlebkHNWmQ0utrk4/QAgrJn4R1r9uVihEqQsJ8Z4CD2k58Yp3Rf
RE4X0qIP2JaX31GBY1mdHvWIc88BLF0xSZ9nXcSeHLAnNrpqqqxwv8L6WUVf
w0SGPGDQ073qPbd+et9bGKgltAB6v4dxvK2FoMQbl8H/0z0t5ypoOg8grQHg
dYfX8/3LdMojAnChue9XISOESytsctSskUe8WsEzVTeDegtFP5872Xctfjrc
U9PYCoVzx+7NYMQNC1aHpPxTliCt6IebUeWti3DGHYNTa1sBFnfZHsx3Z89c
HIdk2qFW8RafE/MPDea/DtHIYGv1cmWp1H4atjNT6cUcEvwFUAAL+b1dn/Hy
Hfwb39PUHiIy+eEjCHG0IbDM/tCHFE9F2Jfl3NOkeilIyhp7580Kci6cGWVo
VxzntpXzeN4zWBeiIzld47G5X4bEVPKQPNQxW8mraRFTSArMSubcSKYquZ+F
6ws8rfBNRCF6ez+OsdE+jyStzD7jzfzOuwKxyQzraGKyn7RJgWKRNbRKcPtC
kYuEJQRy72+lf++lDLPesRihMNvBUaV2HTFm2wzxuOd0sRkuyk/e8LrU3Ynn
ZxDGlEptnSHEiRHRRIdNUgzXdjETLliAqj1H4yAyV4tAVIa3dz4lGKP/uyi4
nnCuPszrMXcw1sXIHN9eZry18/7Qg/E87bQH9TL51JGrdhiNVB81+SRGlHIa
F+MuU6BMqT6rAczTEguMyx2Ay4caDAs7Ec/JKhs2oR0iY6BRG8vjvW8Nx+SC
hQJbqz5AJZvNXqONuVLdvnBVY4SJvWhdu8hFG6EZ6SKfhQJ+N0nOmJGJBYhZ
ikdUepxbNkKPjH3KvjzvZrZtDZuHXdwrW39lvEOqiHTtwf8BILGeolzymeyU
6drjlLAcF6K7Vr+3Pldep/UtFDOlgLREbrUThnmQjO4JRUCB5zq6G1OyxUvK
K+aSkxSNVL7ML7PstyZRf3cUbBrbZl4Zsxm33rzEx5OjAmvEM5Z4pCUzpqmV
lqMF0LAei6McsBGhtdlefOKUn3vg+RzRIgg7e1pB4qDGJE2rHZ1hHXMkc3Fr
/Xgly4eSLwqTRLLSy50LNTM1EX2WDej8av6Scklq2hicuFL4vdpjeckb5yZI
+43bKpsdhSWFGYJuiwWzYNwH7VCCScBHf+7vOa9sz42qYhX+Rsmy7Q/eHF3g
CFkOjzzHGxrAP5ysQYI6AXgI+w4pNKv1nANY+W9Mb/C+0q/pSk+bptdluVq+
z6duQMMpGf6b968thYgjEzXKu379oClX9NfnS+ubci5tCdMjhUx9DzlzQ9OG
ojM3GHZDEB/8VwpsOWxxCNYxcs4TrybkQYGQNF+f06DHVLq8li8zoS3vEsRk
OImIfM6lwR8Y+gZn17s/wwt9VJTV4aj74NNnSfteOmjIvQ/vstGqPjuuAdA6
OOqNOi+XCqNhyF/1CR8w/u/EHrAAfoLk31J9B+70Oz7HuVWB7QQcHpeADgMV
VazmwVOY0kHJe9GhJxmcft2PdpxlAqopQ9wOUc87dkdvhe6g/mxvtYL+vzyu
nvQOzS5JHEUEoGcVuQ1dMI7CAywzwsEWZEd0LwsiwvOImJDFOa+JBxAUqUOb
n/jzEWhg0T0XVSkVX6Ic9mHSFyA/1bBWUrrKHJhQswIZakLHB4ziLNKtn29H
Q8HrfgmR7E3gg4EK1yCLOJT0Ut8r1y11bIwSwaml8ySpANlnORAuOmnway/z
tlvQDegUDWgPIO9Qt9e4tBhObFH2x4Qp5BsKaRPJxcCXq+Ch7iyMj/YlU/JW
YFrFX/HE9FULJ1YZFOUXuPIav4VGYQiq2oIHHwI21bU0JeRYve4+M5S3l0hZ
TkkEZC8nIbwL/V/dbaF6EvoU1keaGMfe3Ee534AJMmsOtdwGoa9EAmksCMrd
cAp+dFF+f70jpCF6VW6KSRcprvG4klFk6NXrDf1/gOgMTI1OHhoWMHC6zTar
uF9GE0CYdLkY77G0kan70pqQnnuZ7Yrd/vBxRRKrFaEZz6fuaNtCEVUsLNrx
yfbH8FAs5jv4H4EbyP551rOrqMKAobTAICvt+Q4wqpcpub28J90GRF/X8XaT
c0Z9+w6odhc6WP5/yuS0oz/Vba3dU9XXyDglizPJxU74BH5ywo0p+P/MGny6
d9eCjdoyAOHOfUZtad7uTXbwKanZKLAMcwms/80d1c/VDXbPzhcT+G7f8oUz
ZptQMQYODCzGaLRGztkcrkmB5sL0HgrjX/o2UTJyFndRA2i/mgJfON6h3U6W
oNR3vxqbUiZYGL/LOjydLBNwlVOGmCBoWOpCarKL0D4dk4pXcYW7sVTAIesi
C+aPWQKPe10d+9FnW07zYrTZnzOvkl6OUr8pWoN/X8/u9OVPKnjRzZAoIqvP
3Pnx6kxQUHu/NBEiucmbMoTj4ozt84kUe9xF4GJBHxEco7Pf0fk/XkN46YAa
Qk9ei3UP12CTdiVop3NCWLDbxxIsTToDDcTmua0SfiTlpWdiyu/+wd6I/C8N
/G16eW59T9Va+8s2LlvPOnUVsMBWmuwHwcTqYH9H9hZa/U7V8w+Fib/XsASJ
A9gv9RyS2sIa5RTrCczHGeTe1MmnZmMh+AtCcTa5Qqj9tUHznuwTNXDiUUkw
eBSoEbZqDJ/4r6E94KXRujUjmbamACfXIbSNushU90NPnLGhmpGXx7alpEHv
FOPg1rTCGo+ecM+rQfXIpAyYeIvWDtJ2nkeMRTH5xRoFPk+xJT1hEcmtumby
mP1RynbisL4KDYcjbSUH1R87LmEk3qWi9NIX6+tyD4s1UM9WuZOZhx5nsnUE
QMCUjWemEiqnQJ0WJS0wvO1nUPyCUKfIwqQI8UR+T78SPMQcD8Dl0CcUXi/F
ZML37DHJ7+rOkvg3fo/sMM3ieQs3BtQ10cmqRVUoO/Y6KzyDyc2De6SmgASs
Qzj3NOat6ewndeAbTaMnQS9Jb1V5mE5yUfmJ5Wpt23L7baO4YcmjEeo/H+2x
d7CuMXecJnY8cDshDpanW19wv+PkjRmhwxE9o9j+FpvR9fZDs4SLjWEwf80l
yWiHaYvf1n8SxlC6UsorNu8kexQ5O0mE39YQceXous6FS2lnibZZX/liV662
++quDNv16z4DPw2PtQALSypFiMAlrH/XFTNF4lSyo8YVt5/o9b3dxaYcQSBY
t4zhZ9cidKwFtuK6VdazM5oPfROsBaBxm4mtjqbSnmbCKruBLvw2SWK9CKAJ
Sug8n3RxWEspi2pWk7YnXzWqzmExRYLqIMGv3KYGOiCA5li/yDJjp+wS6QiT
BlaoPizgf8ve1lSmeX1fpzoCRIQkeFH23Xn1qyYkC4PqyOYe8LpOsK7HpDd6
5XXZ4imZg3mZ5rwQHKoa9LnWtF2Xf7P+KFX9ENFM0wv3AQChDFnAds562Eig
BWhSf3oETz8DHYhrMp/rGA4tQnZ5s59MuBrdo2jnsk1DNktaoJwm6t56Yg/o
TqX4FqkiaqXvpbPAWgBpF4CvIMSV5vmgSWCB3Lo1YkR1LCMJHci8tmwiIaCz
JgdEPIo5XLS9A/LHVQqej450GMt+CEQQVwOdjoOpls/GyvC877tBYAyLD4tn
rc6kXJAhqck9hDKtD6dTIFjQf8YZSb9gu5vogVS67sqfbpAIDIkyCzckCFx5
taS/xOF57dm7eeDrzgr3isDWXHkZMq0POhu7kGYbafhVrMiswdvM3UVrBP3B
S3nHE0NPjhaqzBE9nHLPZAHomcYn4PmN/zVyh6L591J5PEs42dW95nURpIJl
qH2qexkCGbQZgnzw4jNsKXgbRyhq9OMxrvjazUaoFqFiJp+oBu3+42gj2ZOr
6DU+e7iboWlKebPRkl0lVSFU5+Nc2SmL5FBMhwxWkjHQVHYbwUB32bpxkM9u
eGi4LmC3pkmh+hT9FlVCe/o1dAzBYAJ8ysidrD2Yc04/sRV1UcvbWyPTTFiP
wqf0BYhvB1JNwhQEzJUVswXkFQqqXYS3eMymzK/dM29SpvYT7lGzORvUe0kY
GQLH1K7mgegPG1ExU55anZnYFY9pwMr3Rhd00B2yEkZG2ae/9uUUcpmptXOo
FMGq+UCmzs+kPNvdtk71CPZu91rbFnDs/d8dXuS9juAghrlaO9eZ3EwwCW5/
6H7Qo2U3WFp8yL8AdcKEh5I7Mw3WyMesMUcNC3pFMZCYx80akXHaqs9Tk3ti
HvYHf1emmYfq45XNG17/PCG3ddKJYQGtJ3d+NTgubxSXe8+ykNpFGnMmBLM+
1BXZuY/Zh343xCU0EOXDt1qkelPiqsHenlpY3Y8z6Os6HJ0WI4cqXskeUEjf
jnJDuV+61IeAsZsjxPsoP0HrSmpX/68YJv+qQjwMcTK2iQKoAV7RFuNfcR1c
+Z9qDN9YxPeDfJ2aSjdquBx6FRFqKvYsXlbPJZvoCn4YMZJcjRH6LZ8tJZdx
UPwuQkE6HQDoThPVq9NpD0KhphNMM3f/IL0yq4A7FQ5iEVNlkLO5M9BVpEyF
piHHlYxpHBuH0v8Y+gaBSls+tcJm1FN/YXCbOCPm2NajxgUuSFK3oZ6GRxhA
DyTnKqE9tBH1N28165pa7lNaZctVvCKxMoTUCybk1D+S+lnFuMoEQOmt8JCe
jjzCOQCUwmfrSR638XUcptcwkVPXpN0HHf6UOSSx6qRDIjrtsvnQbhhy9SGQ
TfTpwgVMggMHfQRBEqpfnq281aNmDi8ZGyLV1OolQSDlmcLmK9WZOURmwy6A
4IFX+vVCLZrO2JcLiI1LutIGAWHjJ/J3UbOrl0ai2Kg4KwybVXMTeAxlkGX9
RQKmAeHmbaM3/VKO0ZiAl3sVKS7g0vhq7+m9W/jozVGgvojnsjg7HVmaqFcL
E9au+71ba/XXcMKZj03MmQpIBwbrNx1CLOuzmRXbQJuqFivcdzPC9A9VpCvX
J3Y7iK8+1V41gDz546F5h3jXKKKeMRx8Yb9akXk5mXLgTRluE3k2MJt6b3IK
v/fr7L3Lnl3+C6MjAp7q14tq03GJnGy/zS6ormy1qAFWoeWNEIMbUBlaA/8g
oIPIQnRKYjgJMLGR8jXLGMs69B6XyS2PJYAfRuC95NkakvtFZHMngAwkKrDR
MOsJQF1u+9qexCzxUNs3lNEd6MyfCRby2N9wXwcE4DJ2bWXDxGWxO8joQERf
OZG4ObTZBk+hwxh97URK6DEHocHY5eIySde69Rt7e1wTkrW4VCc8TyCpl+Bk
1++Uo2Ay32IY2qOtteS1v0qHmpJcJN5dbIJqLrsQ7xZcZY1uSCDNltBOGEI9
vLm1WtLbb5/yhSYTfVCJRy5SuD33ejPck1zXrN1JgKQS37PnCon0IqL580Wa
S/BSpSbiOp1NxYAr0e1MZbdO/mQnCB1XnMfqbZ5J/kPGfY+tA8CwvGar3OS4
96LcY93kly3GVJKfK7L1XhzrR/Vo8a3BtPbKe8XmndSwuIHgDfD3d7gGUWUV
TtCX1YW8ZbMkNFV+UVe6GlUSPUq0myJw82p9SJEGKRyXKQlgOfI5jZ/d34DE
2UbYMZAmen3aSY4yvGbUdl3Gc1PPKuz0otOKTbS/AowKc89oF0afuCRlG6dQ
NlJDgXe7rpp1P5J+KugFGntHqRg+uViKMFRlnPswGAy6Ax+8Ybs6+OejMfj0
Tx0SSlFFBkd+gNkIkXlQLozzXL8RDVOb8IWH/eShldPp2lg8rw2+uv6qeyf9
0gE3JZaswv9pakn1izHmxVeSh2Skg9FYx3MgSSgMIlSGkjTQy4Mi5+PPFIZ5
57dA32O/Z5AhJHF9qSSjn/RwxeRkGHRQ5tZMfrz0NcFm/6SESR2OaFAh6ZKV
fZq1kVh5XNGRU/uvrCHonyhp6LfgtSsExXFX5CB+AiCkapPQxbgjGv194D3B
eekzhkT7GNWxG22OYu8MVJYZnXcYNhf+xZaaVJhJHiAey5K+QLXD1RY7zNGq
dSnv3jUhP+vTlz2RLvqoWI0thoIzOM9ycdyq0pxoUkGAPujyHWOemn+f/Azy
mSZs6TybTIdyBMNI/H7ynRoQAotYJen0fBdU4VTLAB+l8E5gbVwCCeTuRvw+
hfs/98iv0WB5iKjPflhDO1OmN5IIB64vx1n4GVQ23mJLvPPZi1rDc4Cnjd/F
KHi9qCfLlwrt+26fzLcmRjrQycxNZxhUlLExH9ZAqvnXPpV16jaIA2iQpv5x
DXqNutoOQu9ahm8zAjlVDxUad5exxDAaEAv47TkYtyB4dIWTx8q9+Nn7iAXg
CguuU0NgTYPkhnRRJY8S37k0ddFFULS6ol5TM97UKwbMPf8Zcyp2eQ0Rg/em
6iD/bLkN2aoHw55at1DKfvEIp71vRe/1/LtbUqhIdBvuZVTsDFxKAU0nkEsn
PqGRLuW65+VELoXXKHiA4pye7IUXdhRlvHqlBrujVGzJO3xvjHRUBlSCpdHo
FXZmGIyXl6MClxfx2++PIL0YGJV1xVkhHkuN9ynAK9b0hRfxbz+ndxTdoalQ
pTDdB5KAeOFkNJdlxzZ/WCsDsFFGtSgtWuvemY8Tbj9MYhW+8gyrl/d3g9gU
LMqB9GmHCnEobTvlMrJdJg6+CnAvSA21/SATuLXywWrsCjtJzwNNNWGcS0LC
ygFhQc97JK/L0hOF0ahmW+LM7cSlN5fcndlkJwBFZFW5eR1LUVw0OKMx0wVK
EVSGpda6WMJ/y1EmMmwF69heb/xAOT8+BPOFF29uBwGtApoZmNynWkxlnK+3
n3Y3Ha0MjROHHbAP2dwW8VoqNg21dkx+mAorE8Jj/0YQswK6eExalWNGCEls
INgy1ph6i/ylUTTrcO7JTEHKYDYQpAWy8EsIz5+JU81xrT9h7eH74BK0dbPb
Q5tx0L+zPeLRC0zGeqbfwD5cDAPa+9Pl1pIM7lSr2G3/ZjE6EhCtiqKmyd2V
NTJqTw7+K9jY2xmhC8beL2zAshaJv/sFPUVf1vzoJEYaxl6Fcotf5l4+WDH/
dmv+vJJ9ETt3v+octsjggtc6d2ChDI3KzRDBPMOKQoETlm9mZU/d7MATIqUa
nYZabxzKuBzcfURoqbQLU14f0MWFVq+GEGUMbqN18fu0G2+w/Yk5W/GlpRiN
89pONLyLUrULpSjZkTjj4/Shh1u+fRFhfHVNY6tmQPfQF4CCpGl1vVQfHCSS
R+S0qGq//x5k3m1t3/wPwMDqGmFwiVe+mo2F5Mp4Pmj+oZWs3uloq6z4Ra+E
0QX0Mk4v697X0D6elO4T1v3dyqoAq1uzVYTbta6RtvQF45RKuAzgavlUScF8
IgLGfs8VSRzp8wy+9VeTlLh77UaqTkbxFra3PUnLGI1ek0GIBz3IoQ4bPXIr
bn29DZzzrzGbVmKeUwg8m+S9+cuRWufQk/Uqy8d4+P2xTkNYxm3iGlGBiiFI
cNtimekQyHchn4LSYNiJuzHXwh18lmlX7bin49t/yVIuUiGkavOegCLTqs77
XXIOHrxegRS7WpDjIK6XSO4rozYf170pySiRTf5O8hoI0ZYb74hMjhI8IGKD
lQeRh8cXFzBfeKSj957iaysv5BDxWIuKVP72BW15lE9HFer3krSspRiocmOm
9iwnbfRHTmxU2Tfn83BnUpVsGNNqvn0S2XvaklXd5J55p52eVy1pmnUgC5CP
2P6b/HXp5amFI5/4aJD0xhBoiRmpqF8wG2hQcG8UXeUO8AHukE61GIB6O4bc
SPZP+l5tlboBooGuvuKIIWlPgeKr334xousY98LGb5M5yJ1PEz3bwzzoclwr
xD9to74NK6A1t0TuK4/N6WvUshlRomsLi2np/OLlecv+61WhgLphODV3EO1q
XaIQAd5PFh5Pb0QwR9XImKxO3/tw4JP8icz62ETa2ftdDEXqWgi64CTrjDml
St4anicd/5J4dxcyNwYvey3dtx9kpG52kWfZLX3BK2lIot2gtlyAnRp5SPPh
SafklP3asSahbzsR/+pN/4nvVWG/7ah80h94OCZyEoDl4pvpP/JZ4nYM5sn2
lYHqdDyGa3Y03+pqskvN+Tt7h3OdAV7oabdRExX6B4J4NnihblWV/RJUskg9
YpY5K9Aemj2pV0Q7FG/Lpowj49tQ/RDPyQOi7gR7mqIxruRqnYDLo7uMdkwF
s90mzB9Hvfk60dVzy7VKXCZjQwitQ7ExffibdTPCnVQ+SVai61X36f8X6/NP
4XBGvrD2KBVCLxJ820CBO5ptwLpTPNxhEIECyaV++QbqRSiNsDqDaPO8edyx
P/k1HDauP2pb3/7XbcKHoHFmgV/PSzLhPi0Vqn9kYcEGguBw51wpU+xfMglC
bM+ScZJre4TWateHQshrc3uRIuGChNwTnMBTnKCul/AZxXENKx23LSBQS7pr
E5bwhDvAYxJEoScAhDg2F1lVbTU/wVuOCEcn96dfZ1T8tm6snR0tY99Nfcmk
AfBqH8hNwZcc6ytr4s11+nE6GdG1nVnGmd/JubL7xBVcNCiXqogGIkUEoXHb
Hm1ZYsrwOEFmIysJsRtxc6ImRKxL/uLYKdqO5tNMmNaYsVmiAwVdF1KKA3eN
B+n4qwcnTacDkKlnF/T+cuAANHPIz52anoCJmvXGNLrirdnLn1ZCkvG/SLQ1
HIw5bKLk9y8MGGXAP7SMeKCw/0ax22U6wiLuIC6+cY1DPbB33qdJzZ7kiB3E
TOHJjLx2SUex0pK23KIZGlMDlkJkUK2J+uF51QkExuiqGOUJfr054Tz+zboe
wg1/VOSZWZ7/qBWYCjeHty33TMGOlNEMVC4J0paPuA6EzDHfxa0sceIhq2MA
ecSbGbRECbWXcLP7oCIkqOw8ALPmyVSUb9fN9xiFxylnPq3HOlymXHEm5znS
31p91nqtibc9ww0wxLIUoriIlEiPiMyMJmv052FjZDuPWIlbRxOgndCgumo6
JNTqCU6qBZoPpmaOOqopj5fxvF60FS7e3yJeVsIGKaOPMZglhWmB2T9BF1si
cuyT5i3bbqp42JRw6OQpgUVmqm5gd1yJjL7bWHn9SErDy0NNxKCyMqrQ6dk/
I+Re27ocYWOeyelX+HROVHZI8bYsWd84gjntWcv1Dqn63EAV5Q24JV//MKrm
Mxy5anvZqj+f1qM0JBn36giZsfW+sPow5KTrtvWQcs1b4RjaX6qzJyqcMELc
nUGWLLEuxtgAxxCDdkP59RMYtwIzOcNk5b20KUQ9zR7hLDfEhO6F75YezqXz
wKPaEOfn3sQ5JD0gDtK2Xh0bxUY+cExYUUC7mzG9cn9S5xvx3EDXFvyf3kNF
ZXlPXT1W/JtulL0qv+e6V/hI06a3ArcDxy744FwDlVvV4RaFuoZh0rc653Pw
qX4ecOe8SYfsNPmBVF5AGslsgOpBwCnpRry+CmFLcj7cjMpRa9ppVD47bjz3
uxhVf1AnRnE+WPbhKB9yAOYhJizjCmUwhlyvr3Fl58HP+tGIP7X+0m9+KmvN
FcVEqUmTtfYckplpmCQjE3dZjT5Vs3yb3cN3xQnOXQMoLoFAw6DuTRyX7UH4
SidtaChWpM20Bx3Wg1onHucoH0M+rnIx7QbCq9bEIPXW5n0lgxJYH5G8cGxj
wVJcGa66SYvmiik1FAx/Sp+r5wCmCw/vnPkaFhDI6yNiYzSXnsCQBLbk8Hm5
p8HoXwBomHUDQ5bE4HMcdslboLuBOqIHoSL9hfkamElL7fsSHQZ4x/KfFqJc
MY9t2QWaAbfi8MHaoaWkAOlWzUrAuv/mdxmWkO5xaE9mvEaw/p+VivPOx2Ko
aczBiRfRytz0x1ig+GKswyp9g/cxTYwtZu/W2yGXTKPLRdnSoBiHS8TIXR3O
iR3BgPSu4XdDPIU+f/gDwafqCy9I9k3rWsR0Npo+1yPK4A5hFvOObU/DQ/qX
ONwrXwYdeYdPPbiueoecHFcK0xBydmPUj97IDCvbAuZiaK051wV3Or5GxIqd
Bl92ZNMzX2lwke/QldecwxTBfFBN3jfx8ZoxQuLVL55nCKJFhwA/6c4Rc6zf
6tcrJGsMNMnr2bKHT8utSo1+KzooL27nKo7J8zCEptiw97ga20FXElBaNHiG
gV4jjy/Takp5+uFpNUNyul8sFwSeZE1OOuqfNa8mQ9xFaruW4oTuWU9QukFA
ea4koc2p7fJy4RmyMLMm/KK2AFPUvefhb07eVMgMXKSYI2RlKqSbAmhmIGIa
AHfBxFwxH3++N2UNzlfjLQssLjD8+IruAJLWAY5dziULFRaccwcHibNBkQQ8
66Bk/Ejo89CgChpQGNqb9YMEWHuYcG/QFrDIi+9zkgoT+/RReq/6GIMkrqNr
YT6WFM7EiM0EasD69q7srI/MWv2ke1BDlciQ5J3CU1O5nDKpJ+wOQq8GVcne
cdbcFg0L9zZhmIax4V8ZPLNGCQ8ICyCGo3RSsLbdAvevzNeynVLCCLtazhqN
OfrglJEP1zHS/XeLglsNIon+Kp3gN14TP0e4Vyh0yq3PX97Ria0vNbMDIpQy
Z3kS67Q5/wJCgGZ7j4lDl3uzjTKRHcdjfNBZYs7S74mo+wVyry7VgfR4gfN1
SoRqCsUnMCyhJUR85H9udf/SU2qLNbhMiQ2DZeC9R5b9yR5UGojMZ/xYGFlg
CQ26XAe5/b330j6LIz5ZsAHtK43bg39A48Vodyxp8J3OiFBryYLVGvWOyb+T
y+wz3mdXEuATMgI7pyQlom0Y1s9OgmJrGGpytiZWRGQwNvdhWxa5VATcYhge
ddPK6kYhdds+Yte15l4bs9tC03Xz82r/GV417+l2w9uuhn+uErz24kRM2SgA
ANlf3UJiBR8535do3M3HTmeziBaC1NH8ymmMrdl15BGM++C7jVJMUEX5cgIV
iNZXqIEreUczx+rDfIXoW/Oa9yxSvm4Odta/g44hhKPGO9FYHAaS++DtvyRc
pAE1hOmWu/FFEMe4wibLX2DZPA+AMSOBKzW1ZvcpVbw5dwXoj/NEe131Yfq/
lcF0+94qVAbs5uGoDw1UIQSeo0QM+voFZImV/Ch9RRyyH1J0nksGOaRjTktI
Cju0SwxAV77PAinkLTfP/lcJ8bdS2+wfulR12+Rv9Zg7tK9pSsmkWbAWE8N/
kGRMsxaF3yTLLQrmX1s/fS4fkTUrqoGx3WJPH+S4yjPlfxO1ABZvFtjTf0rk
KeoV+7V9HfX20ObH5FVKdDr7DKqFdtJ3mUQzzoBd2iK+KRv6GVfjiMJK/y+L
cGSkOq1wXB3F07fcHtztP2TOayzk7DgUzA/fw6ZmK8HCtXL18d5laZNvjBVq
+jbJp8jLSKdWc9JGH3Ac+nKjPE2BQo21dlXmgU8jlS6IoXwg0gikO+TBYdqd
eTC6YS10nPVzfK3oiuzEbwIcoZln30TD0JvUehTOqgDXY+oe2lRwwkBbaiau
UIx6UQWjS15p21Kk57K7/EUnw61V48emCTUP8ZM9UTWbu3BgfgWanthbzhgS
wdHFEqUxahATqzePvsHIQt7gTgDm6EhSE3IaYHcDSoo8tDi/tVur+We0byBb
ciHW4utrpyWrICTnzBP/RLU3BbwdqDpo+KFV18S5tSErdXUrCyFat2PiPQeW
MyPBTHeGXCQ7YZ8MloxkJyYEmk+lUYwYJ27Q2xgXbAt1zBQknhXyjh/dDQPP
DNbE5dJSnl1r84iyt8431fZhyTHl4S4PhVPeN/Y9Leu/DHlr3DCe3usZs009
/61G49b/3TFTTfEwg+HQTzFAa/eRFWTOSvndh67Kv7dNrwSYipNp3IxNKo07
Cy3tL17agdICHcN1lCmx9lX9G6qaK9WrJbPfVCydpousg38J6X3ZB0VhygEV
wNeH8RgcIsZ+oqdFxDcU/KH21Yy4NBvCTqu4k+AC6MJESqQ/eA3ZAtjYP28x
BbpSuWgZcp29vAQF2B7Wkl2or8te4vXZOsT+Ol4xZQxwIE8F3foZWEVfJ4Ee
XapI5KJKw+lwJAGSsza/TMc2GVAKx3Q7NygXyXVQ73SKS1Xo91m0PcccQPZX
moKfjDprr+T0cFiltpIuoHDf3iqJ2rNak0JPx+ySZaPCA0hj7VMvv5QbHDb1
JyC73TM9WE+TYtej2/A49FjryhoMka39dnRT/xyEcRBBpXHLeltQipUzB5J4
bONAJfBfV5y2pg3momNePS2fFcqGT95+5xDIziR0DRErq1IQQ48bPtn2ru/Y
m7lEyWhXDt9cCnxS9whutqZaDFSDfsiBNZcWI13dLiez0j3JejH1D2dGa6EG
+52FcXGdUZPWXKc0fwvCIk0r5rnBT5dcLL74qsrutKsEIxctdJsfdy5A7u7U
oOTa3zN9YKJkH8MBAlzdEQXpTFHZeR5ghqATgQUcYvKxldh91RTq3+yPa+OQ
SP3x+H7+nKhLH1gJPb2LIF212f7Hl1GN2/PFudnDMU7HoAipY2r01w51bIeJ
7HwOimfvhYYQCSrTiQ57Tf9WtIZqqqnxH+fjg4zbdSMjaeYZfRcPev7K8Enp
5OF8yZbt34bnWyU5FM/37xozwgNnVvWFe1/Rr0+X80nMeDC3BVT5zySuJ5so
f4Cx9D3zuNXcRCgW6K+Q3VN6j6ha90onCl3q1Ha+NUKMkXlLv9FFREhKI3J9
Bb/7QEF/HYiF748pBgx9xUHufe5GWxCmjd1hb6puiNAT8SZv67vKrFRY5tXw
TIozwa/ZzbfQoeYYEJo5SHj6iH6reBQzXi6k3BJEC/wrm1s0nrq0+B2/69eh
PYRDXPKQI5aV+IDsjjNIoYZlhxLO1x0vy0R+jD0mGCVdtmlDfnsa8kfX846g
waDNI3fF+xh0W+OfbFXl7sxilBzt933u+b+BXlFIS7QXrhrqULDTXYBwHP6z
e2iIwbo0MSTs4Zyw2/z3vaYCLio9xGYsyyLZLliFhnKGo9ar97xr+auHVOby
55UUY/XAfqkE19Ks3xK/cQ75SQxZQlel28HkI55meHdWp8CKccqga73jwvs0
7hcHzzhXxthWUbX67Ql8C6ZLOlirP/8fY4yA1j/1owuGcdMyamfG8gT8cS9M
gR4GUmraRTdrRzhJGb9qt/imR+8K13J3wAHiiRqmMfIwrsrmt6oVhQYzenUr
K7v/cv9mysu20Do08I4GPsHPgyPs1FCauHcRMIfhPSoH+RW0MzLw+y5zDQ55
IXJCNskpv3RjWmZtqnZuUYdRuCk0Ans3EMThDp9BdA5SalBlBzX9jSh9lLOd
T1uX6/fUQBbOAJjs6lTBX1/EO8mj/q4PwikoTwAe7V/osDzXfLVsZZk6X4Ni
ihFPXXZeRTAdPRz1wBIqfhhXWnniiI0zOeJXhLhh/UJQwPqDwMJb21AXNgxm
tzS9DJFKLKC9EyR0cO70mhmlSZgmnk6/EoiJQxnETK9BGl4g9Q+Qr/lsreLB
XIFOsr3GknyEsi/h7bnUJhThiXOMKNHbrDpCgbQonFm718+pA+27t+GHc9+s
pja1NcHQVw3lh05QVNX/ucrDa87QeiRiG+W471gdqrSKS7IDAhnEN5/NVF2P
j8feDA7Kl0rBJLDWJGAmfltuR2d+o7zrpzHsqg+G/UY/H2p8XUKQOatL2mpN
/z3SUnxLm1Frfl72knX0fTdsroASJsWZnRi5OBPnL8rq6lbyGADhNUIvO8Kz
mibemigNi5A3kGd42STf9S6K8i+u1rlWnYRH+R0DAWSccv/lVzsDky7R/gTB
tn4rh3rxp8HevZM9ny73Va3zrNr+IWFUr1trvBXqCOCejJhxQ4dY07mgl+Pq
gIDGtbC0wigGJhvhADwuplt8zmaAL2x6eQXVW6+29iCSuVx8mOVb9rw+TohL
M2sqKaIr9zYLkXrcMqsMIb3doEFSDNiydYLCoHAAg14RetVIP9KQKPODYG1M
uLkOtzYf6gURrp517/cJoo/zO5tzLz9Kt+Iqs1GdZ89qEXUwHIGa7ADBaDZJ
tFbaRX7aYsGbyOJrVQFUcGe4V59bE1TX1MdAKGsKOgOhMRgtdRdbqBdqwiuW
11yy0O6igXxkVGz6Nb7lpVctgWyY472zTZ4pqhtR5EEyJWIMbc7hJkhK7Iz6
jVTCTnRtCyVlif+zK37THy22fj/M/ahzMK+CrVK3Vh41UpSXGiNLCh6Eei/1
/UXPHpZBdVc7h8cqX3TF/vAXCAiS1dJkbEvbouaoKs9a2tl0oFexCyllQK7y
w7DrOSZY5lmlQmLgADVoS9rAHBwT0/DEVc0A5DAfPRTe5iwyh2uml9vs3fR7
fAAwfoZitwCcda/Gp/ZRmskaHU5xnr30u/+fObCGa1qgDMaKhZZ8bEtV7tLM
mgSNY6eKnZArDGqjJUMIlAPkEKLkxSfyRoevkCjge8AoudigsNhbAKgA4QF8
rdMAmtqpWitFD2ONqdZtRWeshMqZFhjacgZETHEP8Yx4+I7m4sl5FhwUQaMB
BamFlWorBCyTX4VqaPfgKcLsaPLcUg91zopr225T0Uf8vOjo8XgYMMxNt8SO
RA0g3dZCmxL2NxTL6DSM4SNp0/SxlEaWsHPa2PsCgdtJdiIUiUHKJSbmyTkN
LVLnR85Ayqjbw0bpt1cyBpDq5ZB3U8BlvXrp49dAZZglIumz8ztDUxNWdAtV
Lc6wIrCoDdeS9VixzQNqZdljKIhs2La2OnlUTXE8lha+N1JFWVIpBUBG+pM5
SGhElQOJWKY4RNuJVVPZRLRPB576Yt2qxCHXiIllkOsqfB5DbEp4Ohi0rHMY
JkJGyg4m9Vs9PFwpj+STueMKestlSPkq9Gq1vd6tkk1Cu5GWGigqX2QL4yWc
O+uIcfmHhOY5GUX9QYxGivWVzeU4fKhiqWc6wQCoivl1WbHiqHviLiFlwuqo
f3/31FHyRNzXFQd8CWnFDL4nsVSwTjVj6WyWjUsXe8LnwOtIhIxjlkfBQ5jZ
VeCtLZliT7ASNpmNhS25WWJIKj30Tl0H3aCNsLH/Xd3dyE6aIA28CkNUmFVG
S7hUwMsSmpf3Zj2vPPlH61H7vN8XwZ8qGaI4UiKJLWwZBiy0lQ3JTuCJhrpT
sayvaOHVdonGOUt7af681QD7WktbyJOAu0raXxMdpPGl6I4lieH1vmePDOt9
nrRVEs1JNeU1QTak4yXQmHRSOgMfZOVMnlCyjr0tj9RDo47yilNpWBnLWbwc
K1F6ViXRwUPD4IvBD/FVz6meZwScclYYkXdnF+o5prA8UL8rRtEYqw+eAQNG
h209Wn30OWYp5RywJSFREyE1zrWhC7Jp6tLUaeACbYxEM8XrBCiNRUgCX5Kw
S+Y2kgun0UBVzIJW15URpUGThwV4lWadIaQyq7o99hM2inkmGFu4gU0mBTM7
PrO6su9FEfPWuW1PIktEyn1DU8hwcJRkDD9ERcGax01DJvdGf+3QYVFaIai3
pJ/dlVodwm6nrMOH2LpTanvxlXCfyhdpz0Ee6B7hxBZ/pKyZEl9r/ogX9kWM
gYeG1eirLJXyhj8KvewW1xQLh4jShSb3pZ4uyGkDcUmqylo2gdthqxEO5Uh5
N3dN0WQiARlXyZzoZxP0UNd0tLKGxTYOIEGmMS/Rzi68EnnA/Lsw0AAx1igh
0PQN8EP7rgi6IxMUXjGqZtni9tP4QpORN5oKHvt76MOYfymsYhvJRIrdzKe9
TVFPh05+nonwVYENh8vfplvkIeFxqn+oVg1Rw4dCasdi0qgZGag6G3ka2DFG
kdfNDaBvxOnkoMrQHB2k1kA9/JBvvMrGYoywRwfSn37MzEU6cHocqX+SMyB8
+Ob1o/iL+3We1f+apc8g8K5vIhQjoxlOV88R8yaa11tot6fwTu2Xhd4/pFAq
BS/6YbVmRX8GBKtQJB9D3UfvhBxn4v/6vHe5tWpjLPruuhHdz8gNaxfrIigm
vAdA46bz9TnGDdOOllzMKk089sqACqEVMWxwMKe8z2NsBhqsEZz0HMwEgPGy
lBEVk+5Q7BxOMvm+dgzp8UFVh3JBO3ZzpHEtzcOIPbRxzOoMgYOLld8g59uX
3dhEr5M8vvTBav2SBZKYIltr0xJonjYkHS/w+UWf30KzaEjUXmmbWB3AnQVi
HN0eqHyLJkew+cxMbgZMBy/iuGmomGP8731jZIAuALS7uVmXQmk7Lscbh+kU
0N73JjF21bW28M1sck5AWABUwq87J5nEm8vBKmoi4dpFWQ7/5DNlML7XBF67
iRexO4O5Zgj1n9bv4N1qFRsbAYQ216/sCkI5fwPpLVY+rtO72mzqo9W3mPUb
7dTs/wf4lnXBtGI8UoMx83PrkM3mWGbyCkhqcRtGno93/7vtKs6iuwxLKdTr
VGGFm0La5QyIi4dGxIZsKx5Fjmtww8pAUmhGFAvjWl5lLN3Tce3p2S/wQwoM
kReDrigNP/prAEQ12lG8YQjTAEXXWY2R+tJEH4nHAzM6/Q2G4XHUwiIefPOK
l/bb7TJFiEPNitrlFVhdIUdkZTXi61DqZbgxojGRAouhreRn0nREAach2NRB
G9lQpqzkJmuHtdMKPTz+HX6foyNFrvQkohwhlih3G7vbZ6p03QYkG2bvJHxE
CxQRBoVgSus1V6SeWnbKA4Bx52g29sRhx67Qt00yzn6z1TzkjvOqBeY6Dsf/
OpQtCNfq9mjtdEjGxN0nVEyro/KhMmO7dz2/XUNtNqkp1hl/kmpBb0jO/TyN
iNCh0etiKiYgv28rfUQYGwT1zhtONzQxdQc+pnoQxDQp9UuJzPOVXZK+dWdz
VjAtkXx8QxukP7u7GdeB9RW6VtCWVm/5tfEGnS79T9mmLWPJmEduoau8CWnp
dfTVCNtOOULSaUHdpt9xzFoMEkMV+vYLARPXYDGSIWCQHO91l1g1KPylSKuO
Vttpg99q5zYkwSgj3Mtl41gp68Wj6M2AZ5Gkxvm1MhPpkAMtHTUJxSsv0qBQ
0nfbx2kugWgPGGQKTLCk13bzHcbBW4NEQsKjeYXZhfqeZG+QELn9le43XSai
RqeP1hQ14AGFY73mLjCc73wTwM9Cl7uiwlkYcBmhOE+Xrh+2YLzQNQgzflMa
s16etIaXNVwdZNWvRG1XsIiAppfBIS0mMm/p68MrZ699MbrS8wLzyrhdf1Pq
eUsxqEv24eZyf1DVwhsMKwXJiJ6IpopTws3xqTfSBXVgdlhDneidNvDBKxQL
iLq02gNGoyeIRHKf4Rc3vxTT5XPNTFy+pfdG69upfvpmFH9AhQm1xzzVUwi1
d1r1RPpHYFStOkhzVxj9cgGiaJOIi/Pswirpx2KGEbO27LgN7UwRwZGUA50y
eTQdx7LRyCl6KhwDxoXKIqC+447Vlamr5dHQsFifdXtXHCNArsUEe+JOufh8
9U8ztPJYH+NsVsxCyjEpVly5I9YBgDyXD+d/37BWDsx80hHnAzGv7uJiAuqT
4anReYbAyuhEuWWNjRDK8nijPGlgY+HL5sp9QvEaHIuG8ZfIFisaq9TbYSau
7RpDKtDwBQP1XPFYDhuh1IcNHtOebU0Cem2okNnmbVuDH6gtDZnbqlSwCVJV
ck6vXz/lr+MFV1rs2Cb9Kpgo4xp9f7sdH61+5JT0OPuFNmKmz2JfeooYmoz4
P0w13vnMfRrjvpX443wOY9kMplsO6YQOCqsMZS1BKo+yc98zbnwPc4yvTVex
IGN7bZVJC8kOpST5UetJyw3QAGCQbbD6pzs0WGkRduss2InXmWQ+1aqzHfAN
FLjOWLZ/BXHP0kexIPkR0qXb/Zd/EfLMgcjmJA7s9JKNIDIrR/IgXvpKNlaC
xyKqL9jyUdz/HtXOM0JeuIoKs0viBuofCYMrzuBN+m+HED/iWnV3fleHQ95u
348KXpnSjv9y91J/Z/416q2kvfLyWX8rqr4hSJV1hDcyZINeQ+yR4LpdGqzh
QCcuZ5RJM9eAZcDSCISDn4EXstnEWmD86UlenkavcMxgofuihAXFA7WhReIL
AmuzTNT+FP5n+Thoo4CdI5yfT5NoXFZw9vCm1Lt/imo9PSVPcBspDPwGQmYb
WRhoOAtG6UAyRgA7JyBvdvmFb0jG71Ob0i/CBbZHQEtO1NLZ/C+6YR4ncF/2
n6KsbuSWaNoSCJMeGJeFk4lgWEY+SIZIFyp2s2xjiI0oOK1SfrsA2UUPj4oI
rQ3nCplFQo5RISu4LAK40PL6iQSsbsITByk43HITy65UGNIRTmAgPf57s/fk
Uq8ChJweuPpNL+k03vViI4JDKEO6HuFmymAqFky0aAfGDpipcq5JOj4HujaN
gbY5PUe6z/6ap12xHm/6913BT1uu+ICf3YhuyKJi0xKYIkIzT1sGgvmAs6BU
LU/EISJFojq7IEZnzvAz/IVN85Nrh6JWXoDzTaOtNK3TTG8S+t3cgMlwM+n/
2aRo3clNNn7SLtpFCZ+no1HRTY636QzXnqOk2AB6ooJSemN6AkcghuEFjECQ
n3QhtRkgJydEN7gvgdHRV1eHlcjNEgXTIGL8w/Kl+oaov5qp/okLqJrgLyo7
Zn50M5Db5DvR1nQmnp3ZxLriDcpYS3swrc/bYuWp+xy/fEiDQ5fH+wOslQm0
R+LlIyFZ2qnnseq0gEdv0QEPNqBXdeb8f4sCrd7/L129Q4Zp8AW2yzTKo9Rv
bQlLIRg3ETGWLiBPe2JMVnzkrNdIGLuzxmyGhc5dSQOmsIIn6IYrlZq6UEqa
X3X6vpO0KHmRg7BTR9YI8hgOH3aOiLqAfItkLYZ91VSbz/8nyPplNP4gE8F7
1S9Yobv6UR3TCiJ8t+bacaa+02CEGzJKo7LhT/ikUlS8wauOlTmbIRkyqyuT
OzdB+229XQkIk27A4CfZbZ3gWegyFcsWLcRrHBBwRbsL97vOJUHIF4NUVAJj
Q0/55vMF/p7ZWK3WQXutBtIm1lr96NIhHYHM2XOdGJyx/0PUh6zgtqmz9l2B
gbiCCaFmTEIZCYu/xkR3n9p7tjj22uYKtNmfEOc+g/2tZPCW3/rO569zdGwK
G/qpbGRM2CBYAbGno5O+LeCSjAeAFF/cwQaZIJmVYBgpbLA+KSP254j0amas
M3V30a+M7cJJeiLeEs3umNygZAoZ3L1i2xcXdJEI7XvtaQt+LxhT/rUbGuz6
AWg4O4AhZa5pbF8EINE1czv3T+TH5C2CBOzB2+Dv9EdyOQdk1kJVE9asizHg
MB2CmtPC+OEiQVXlawRglH0GGkaeZVkJG6SaI9NLAyx9goESEKrL3xP+BKki
SmntOHYCSPklEdC+Lc6lPQ1ml4NC1X+lE3pM+X23e+Xq2o6M+lkXs3wU4ndO
S3VKn1I3dEIdQ1E6YqSaEztBZDHSqnv0++dAImOmOG3YFzQbfgQ3Yf8JxJDC
PyK47rsJK9kpZlYM4kA/JL+FrUHkwGS4v3ggKdL4c+cKUKxrNc+ATPkZlhX+
pRmJMFebJXiCUudvZVRhM03EspKxNAzfbUYXPmhgpSYy9DvVR+nkAu6WKbM+
k+ZXE3H2zisSD5LSvl4DPJez1SpvQfUTpLXSZZdo5Z9/03W9mqgcNdzD9P6u
HAJ76pPPmkvuufYd4WcGRowEjn51vOA9H5EzryhE3YLRRTa8j5et2jr5MjVb
YT1sNXwAplD4wgZGbrTl6emVK65z0oXBDNv0MAlRyDLaSRF/XA8uaz6tO0dE
Kc/ZHRzZXYJW5v0XwHaI3n5M2bttE7LxLUDZ6PYfE0Mh0Mbbm9BMLMUM7HHu
1Um/FVZ+uyqMEvBvkGG3NotqQRM4YpJx8/USoy3nwSKG5ZhkHdqSllbaqdWW
MAXDThoetXAHuZSrCtekAgDFjqJs9soosDO7pR9lVg31gE9ZkOo6ANLSg2yZ
SrOwQIWFQSzJsz4wM6p5b7h0h1bSnk9qHSl66q5Ox9NgFDvI0dj9WU5x1kwl
z3fewTjc7pusDJOUQaakjzYZto2eKfjOurAjQNkwRsHTiQK1wYFWKnqezOMQ
5xNDjTDsqT2pogtTDcC3TAa03y4GBBYZlC8XvQFVHqv5q+tOFxvx6NtJvJFG
CJVJWXP2F4MgFxN7rUzZHRbC+TPA9a41N2+vfuzJSySs5qZwZAMgesLiTfNm
NqEFyIS3q+EmU649Q5mP65twnE0QBZD/idHtlTlupft9BIGLKogwrZ49reU7
++20a/U0riJy69U4+hGvBD5vtfQ+j/MJGS6f2EVdoJvvQVAcErD6XpmghYui
yB4NVIfY09D0+eS7oC/qJh0pXL6CWhnzqiXRE2okGuOFsHKy/9GHoQdL4h7m
kqgb6CKGO7UQg+zqmBcGfAliYCyFJbKiPKuxij5WKCKp80rju/eClDr5lDUT
YjBzgvDmDq8LG/C0nUO6E80/PW/OPXDZs+ssvKsyAG7ch3kfDfpwkEBjHyMu
0MHPrEhrZ570wvA38msnKisRc2Q/o4RGo0o+06A7GpxAcykPFqUGjbMtNUok
mKsEbdMC7GiWi3djTEoqrEtORVLw/JzTCpWpbRO3/2ocQHdzbOA/f0YaVF3y
vHiH8XwF1XNjs+9PMh7+mxD/I2I0UAesrtZ6RXJnSyPU0fPiV5vdpXWh6ZNn
bDIUQ1N/j6MlS2JgqTqvgzoQ6t3MPPQt++V1pAXE/DXe+lxbG2QrtkfDq+s4
ulNLair314dMf5zvDkkJRzVQAtsxWBJi7fiVwCvsEBPdD79cxRTFLJhJPytR
bb2dRmi0Ut72QbkLU5AnierwQEYKWwn1ouZ5nlyVzAYHbYjUPmVEmZLFYso2
5ltFcD+8W8niKqyWwdBU2EZuyZN2m6LKSaLIksN1ZEGK7nSXwy+aZGQU131F
eUTWWEmj6XPkq7wigUb8yebjTZPLPIScoUnTxPXEnSXFCmySIyWRn6s45DvX
qG5zsieEbVCq5vmUlLMhUjRBHHr5RfM5Z9tqgf/CxHQL5J/EPY9PvhvHgCtT
Z3YJSTPzEE8FTMtpbKyTN6yqOur2Dq1sNIVFzZuT9HlxNa3RVLNtxLmcXPTC
UCR0Bic5zziWf8Zzl/Dw2sO5QsCG5Yp4U2ENBXenIKHEPEWIeWzT34GuOLqt
R8OIwWZ7zBj5Pgtx02eK6wZ8pmV0/J/X6IFGLFr979RvmnbXw4yX+QICPDhZ
4qxxeQHHtcGe519XbTJ6pUJwSA+gMRYCcVVaQ9UGWJKM8L5PEvdFbK27aMDI
ehNE5U7LC0JlQX2dvQHTaQyOPwg2FDS16KC3TY0dbst7+nnX8lxAnm8bEn/a
ATpxeV4bEWFIw+DNNZTgBp2RNJ9vCHy+hTBEh3nXuf/RS0pbHVp9THu/Toos
Ef/UBw49CbPzsUqK49hLNftd9ycA2+hMiw6GalpY8HMhc919dwUlgImVRrGi
ouWcBFRG2RC7uefcb1IYd04fCP/8tHjscBwBlMSfRYVaq4Kd5w1NQjvHvTQx
mn4r/6MO3Q9f6IlsqXpoc4DjJaU4l1YmoCRGJhlIXnOw5F3iEAMXWl9wF14r
M30ckCkK/nYlR3lpnbvey69zuuJd81ycdaSezWLEe4AdQ9ynx4MoLBXcjmpV
lUngX0kw3bJB6a9ZejOYXoNQYzvmZIU3HZzVGMJJTYVqST5riFHQAfMO4J5t
mVT41YFjDMqZtYenLudXxcJp6ZF13IZfeuN8fZO37lehz7aU4jEs/N+I+5lZ
EAahgsWgVmRFfc2zy1/Pf0jeYr0DRSSLYqOKwb+iaVLddQeST/p+THkSscKo
IYTov3Kh+b74x8C7DLLYAc9s8t1tl3bgHsWub2R4UMk0Jdo2ksvo5gxV1IDd
Vp8v5kDEiAC9FYd4ULkME6PcEJRoftdXCHZuu0SALlNvbN0b8LWlvrj7YAcY
aKI8/cLojiXIIjRM1/GKuJxCEFiMD3Lzci/+qSh8Ctqycv5Fj6Hn3DafmJB0
nHh14EzRcZ4/nUQLnpyqrbRKKtu+GegpAuw23BcypAjim7aG8ZPeQy3vh9O5
qrR3TT1pYS0CbWUokqSywZ3Q1f8ZFf3gj54+9H/Fu1+2dtfUHB7/Wg8okNnq
eZ/DBRkD5FJjzeUJe6D1m5LBqDX0ZJRw2d+CpAXL+c6VrlKSuMBBI6SikDd4
QIxm/fcHLErQ8AMn7/kx6KFSXru0Zowj2A6YSIDG7dwltmBoVHNuCosn/zml
PTfH7topkWjUNgQXy3ak1AtYBfdvqSojG8tTa9SYg/eGV18xF9RdCq8PYnLi
lMx6gPrFH3Iif3kjq/cKhkzHxRyMx0c5apgTjPWu3CsODzrQiDLV25kmnDi3
uFha8dh8xteLvBjgxulHTL4ckqAUI45Q2CrgMprH4VHHpcBd6xZL+Ucqnv52
InjzZAbpWMJjokjlHlh20rInjN1Phsja04JmOk9jqj3DICY4Cwai3X4a/7+b
IhFiqafiKYAvvgIm0pIh/7NL7553PkJaSyQNDAluf+VeGTfh2WDdvoM6jylu
3zr8xAFwnyKKuwr/IEB69xjml4rM9RxdwbbEr3D868pMVqotuYEvgnR2Q155
woroas1Ntbt03JmuHRJsV16igw+AZssNGfY0rYtyj15nYk5WvCEI9e66819U
oonlcGrAwFOMHhZjnzsg8HE7Pu8CbvrQV4JoJcuHgup2c+vt6iG9zf8seXtb
WSrTluRMBWPm7HAr45ze34fStIRcZJ+AcrNV9HjU09Dd8Cr0r/m8TzluXWiz
R0/jnxIVxftVLgFD8pgI6wkoBcU6E5OYVD9ZiA/gDMA8SqCz4YSo4EBaGHiq
1Iihjwi00ST8sqynTSCuOcH/GCuWVqWRlpfQjLyfrKQTIKc/p0d+BFZYBxNe
qS7R0NXuw/T34SR38RAfxKDdrboIxZvhUCVHwu1+lOxeu2sgSlJ6Cd/Ys4Bd
Qr2Q4uqF9f9NaiVzlztVIVtyzXM4DZXPEVb/KJoKH/mcs5PiN4RjxtwhAOK7
dJkGfb6ZScThuVHsjCIN6FaOEzZ9lmrZt/H+ppCKUh8oxJ7CaqZyU+iWkpfO
eBXNq6IVILEGWsBBewyrv5ppTMMKjOtGryHjdwafbnQIyV8t9Xzb7LTsXfLk
qN2/OVgE0Ywkl4DR0jR4CI7SE+e64G/CBKvgNN659LLZ0iW9LVL8t9b3/Kif
wCBDEcqBwhoiCj4d0UNPr+FHJsVynqt6nKt/uRuXhUQ8YinVvmxLG83RdRcu
a4DjRB8G6mTNwyFOUAZ6+FOgrqKyv0tTiCOgNA9N6mne8DAqXvYRiXWqeKUH
yOd03zAlEEG4QIRxk5Teqzl9iVY6oT0KHqsoFJ+uFtw+l7kuezF1WNB/Y0GB
qWBPwNYRmBzRZ7hn6LMLtk4iDNjpm91GHCQ2g7eamFk4TFUO8C6hEyNw80My
uBn3DRTayQUOBCMlj58V2li1vHS4vYq48W0B/73LcPE4vvcWHFJHw5YsIW1g
PMmRoS1bT8DLOSITBS9foF1W3WnI5ImSO3LRgcyZyJHMD7pAxXcCM22c2trK
gaAS3uek3MmTJdM1Xvm2nXMptCQzmuzBIXy7ZTAy9kc7ybL0jwCdDVwS4Fns
2cukkdKTYsYJipfT0sfbwifh9ZZbLZO9jKQShfRb/lFanqplQ8AJyyja5BtK
xKw2kYPsHol5hfGYaKFdf9CyTfuLuSwVNurzvHOJ1pUeFLluXud9s2zR/1WU
GTVGd69+/uC5zPSNUZr75fh7SU7025Dg7ZKrsJQ8k6elZ7heOWOGBNzvr6vl
M7MZzGegP0P9CXeWsSeKtmcjU0fhO2y0EfBeF2RjvP8E4kD9b8Hhs05eh9hK
nWXA6jkdXoDv7uarXoXuT6XlEMuP6ZWXlKsk4euEldKBCoGFlci65AMMImns
qbBwRksWLiRScabm1xoGtknJN9XIrvjwCp1tt7eVTQ3Ma3+apsMqp2+tjMPZ
LKbVdxNYLy0BucxcgP3VVz+HuA9jSzLy1tKPzkJLwWBlV+v9k9wlx7dzo46C
kvt3oqs23My0d+zuw0q14xRlxYCuv6AI7JYgKx05RU8ufql9Ffk/G/YaDN8u
kKvpO50hFMuiKOX+jQ/mxuJCgSEySRi0a9Fqg59hrJOvDiQGoW5RziMiTQxN
hjVBQ0b4u76knkGSdcbBPRqlZcxb/1tbGEDchcNJwXsqHkmPD3jb+AihqMph
GnBfE7RJfiyZJ/XDh0bvIHohat/gvRUdrrJmXEFB6qqtQ0TOJWa0lzwCMACr
zjNsVcNZalfjyVUf7uQzKJrGFItEw5Ej3XjNq3B7di7eXETeKaWI/dNhT9cn
4zKCy9XwgqJTaDT/Hfua1LJ2yaQIim3MBViEdcbEXSaLCXfTcOIQcO6rB7qA
nkLUFgWD8ZOnGd+NIDNqN6FuChfkpea4Zwc1i+612XHb0xea1cmFR5lldq9e
0bjmnCQa5tj+TKudS9/Qy//s/vodw9g+89bRQ0BCZjzMfz5ZrxCXoR4Q+9ZI
rwLraqD8JsvF61VZX1gMn8rMLNl4hMJCcCArrcOXYB5GPKDnZCDuJfjH/SlQ
/gpXZHFt1VSd02yy+qVyBSXl5VL/Z1OMEnr4ATm9a7gxr5fBPu6fEfonGuIT
FpogakMa7wpApS9GgdlDmhnR5XSOE0CO5VDlQDgN1pICkCaYPsKo142X9MFF
lXjy8yyJDMjTkh9MGodqqhjwdZ7sq4U44d2Nk6MLmSwQbQXqm1G42eXDfEC1
ZtQycCP0oToTOh991MM2/bdsevmRy4tH4SL9v60CJGPilH433hKhObUexwB1
UDfkK0UfBxPBnsHVMuY9TjrFj899oB1VbUo3lrYq5ClOi+btF+51FZd2SmV1
Xzn1U13dmf5tbVhfj5MudahSKOZCcLzXG9kgDSO4w6rKXYbXcVpVBLPm+Pb4
ZTeyuvvBQKvWnie69K6b+Mc3iI3sTJP/v/b+OhO75w8QGTLBHXmkwrDfgXJr
3LFlf1FI0NeOlxsCykAhwUEXNn8OkIiJzY8GT06UVLaC1xuaMz9NEyQYN56S
YXWgHRJwVlM63PNG6wxVnK1sZkDQfmAUMsbWGLP9CwRvM3Adrnfj+qsP6kNY
cbslreSOvZ+dovn5wkowvGQSkr8KofcSyZWuoBl8qSrYHpimcmEP9b7nhf1N
z9pIrxSGidAGpxtO73/UJIaBv+82QaNO5dAe/Vlk8H9loti/p47YRS1Mo2X/
EY7tGzQWG4/6gzW4WdQvF9vVBDktOaEhioHsz8iOxqBxwteTh7p9u8DVKAIj
IqcQoYHJPN1DtppDt5ZDXG+81JAu/fe/TXvC1neKIg7sYgRHlSXDZTXx30Jq
QrMu16nyQFYbf+d6o1NVzhvE/55Ko4hiEeCnvcy/vfgln7/QzFELYxosKfxj
SjU6UHfQt3+Acz6xbi9QXjz45/Y+9ZzF+f1jG/cow0CMianEZAHD9bdQJEK6
Lug9CyX6hmYLHKHNhJJp+MJXJ4VE9wl2ovIUIKPJ2r0bB4AFZJ2bDrvZ5TGP
4yABHj44D3LU5hhJuAarNjFCd30pDS/ECBTPWZQDECb4sYd2H7OwNwP7Bfco
rohVsjAY/uGOZ7WLQX7BzGIKXVMcvQ7SIhmtkeIN9fEj4kysG8mOSVsBpn3n
O8l2KPK6VowDhDPqZa/4whW2sDsN4danGZyj5Hr7m2ALxBHhueszhvPMHuWK
bYrC2AzzSumcJwytu0++OG1+lzNcEj6Kw/2r98LU56AEH04J2Oz3zo2oVXRK
Rqh8kQmU1aUySHxVWMThMDLEGkAZlRmU8cZWt7oIdD9G+o7aFSNXws7L/Cx2
ymhQh4URVIzjXmSOQNtPh3xUhD7cCWf3Iz04OMnTBKqPQSn/aWeAJLYJ1Qrm
+7lH70K4/V60hkf+Jsf+VG51wfvc0S704gYSFri7AY8WEpYetrN3aGeKElK6
d2B4SdTD0Grw4w31DL+a47+33uAosOXuTrCzpLuv29GpO8U7y+u0GAdzw+5u
okhSROuG8LFRPAKNgjYliv7BIaPixoaVVAlFC9/n7VW4PmCtSIFpRW46rhGl
SHUl9m3SpBpETG9GbSCwc7bAPfP0mGAGMDaeA15f4bu8svcbvzaBTxn8y493
RxaDV3sRT2aw/qsFJHzl1WKKu426y/hC5o6RhTdKUQbmZGDgfs3UG+Xj3oM5
++Ge0SVX6vqTZ19LoUbHisbpyKoWUzHQiVnQAFJqAqy3/z1+OUf1Is+zZOAm
jmEihkiUCP1bYcZTbe+CaQEg7SFAHDTtYeygGTLmrSRIRp3y07jDR+15oAdq
yM85LhMqnscMjQVm8Tg1jd1/9wYdzPoSkBPAwSh2nswoIDj3exLCwMZWxDhf
dJGMPlh9JUYzLn/rTbZtuOyNmCOTNXuTUI8jLbpnHosX8Udh96SOC127nE1W
2IgReIc3G1kCaywTlWEfVnhcc9IYaCHf5/TdsKfkOWmnqUMpMYef6FErGC0E
RdMtMJBMzl+Ix+cdR1mbcMaUb3P8XVLpAkegWZgokoPot0Hzt90Izrs2lPxR
FyLClKocDib2T6C/d8J1wMMdTtfqg1ZiSsOZezWsfWaNUjmsitbkguOhzu9w
pMGVdLAEQVH2xGmTm0PNsKvUZaZDV3eBHOxmx3uYSyJG2XwYMI3Oy2GxhiMf
xJNWJVvbmqlYbF8gN/XfzNfbVoa/PNFXjwijGvcxs+qJOFmgqghySHLelRXu
jjru6Dsg2OszjDllc+6NMOF/PxTSrfvxfJjbumZs7n5ADHgwVpahB+ISheNb
EAkdePy9jtQWNUdtUMmLDC3dRnceGoi+YFcPbeCpwCT7YVhCV5RvhdSafblm
NintuJ7oyJbO3MWS6Zs1htr3fUNyRZHTAT3QvnkMJxWAnMjY9P9tTwPMPyH6
QpfWMbqPWSnF7Xcl9sPIkjPimdf9uWiHvUQTzXGANWH+gSd2lE1zaS8vWtb4
nFXqkV9ml/ESPH5JBz33cgvvBxt3BFPX+DAAXdTLFqnbX+xPew6UlyjtgiVM
Eg0Qp7FhanUl2vYGfW/SQMZp4LGYeOBWSN0x23XknEmOPNamdb9fNcZNtkMK
y6HxAW+cmxCSchhg7pAFcE0RqOHPeXEG0o5H2Ys8XGR+y8GNLQ9jv9GlGwlY
kzLK3jP61P67ChNl6MTH72hcTRfzyZWzN0BIUy2MGaFY9s+fjP+M8wlt7YMS
ZX6FscG0AS1bpkA9wzRCGZ8tQ9+WKaMVsqou0iug02EIAnX/Wg/MXfzrtn7p
E02fSRAmI4WeDDIburGvpD8oSp4hWjcTeoJEzVLLsD1wqxXsAiWvml/bx1y1
vq6winY9J4Ks6eYrCMv41PtK0T1i70ydwrGJ7a7uo1t+jo0TZgOhK7ohm90M
Pa8s3a5khOrxrOxITcluiSp9MzwJH1k4awdyV/6nNZ5Wc1slLSSrr1dHBCHN
FrNh5Y7n/4r8XHl1mh6wGPhe+nuv/MNBA73IHTPQARyOuwx9NUQ9Gan08ub7
RugpfYgCvhUu2OFIbnWVs0Nuva8Kh+cFeP3IOIPrwbsJahvbc9pJUVGewm08
eO56WWXp11LQrzn+U3zEgDLIn08qFgccd5CflS6UtAyf1XZ10r/GTK893lmc
2j0d0pj+Uwp+9IHlMVyNG5j6LOkt7j/CMU/bCLYHdtrh8mSJ0aNIuBCFCt1F
lgZBnJqYkYnRdlYFlibD/oICRnDnVuMWbptFyDPXh7FhrUwWUyk1egMRcZUX
WVxlen3pKPEjl7zKftWzcm/IJcCf7dFQ60QwvQrCq6d/EJBTRh8VZMrk4poV
ziqXBE50pkhIvUVovZTQWgrCqL1eYkVne+S7wguZeOeOS8X5rFPYo/Ohnz92
vjMpfrjqjirf5XKdBixF31UyL+Ui4juorI3M11+bJL3cX8MGihoox2xQWc62
mrSPghjljtIiuw38zdZS7PLmdMu+qj/R5Krj+y7CiTtbuzY/q/msEINpQ6jn
PfEx19LrOb0a3jIyGTbzcBQi1dgtuLYjD2R+IXn3cLUObHYqOiU7h4UmdX5K
BvkqL1jLe2Kn/p6fYlXQzV0KcD7QskEH9KmPellhuLA4bj9LlWQTzWg/5Tpl
GRdsiuWh5hjuGAamJHgaolCLjzhwXTtlqX46QG0AntZHbzZqegbfROzm9lN4
67MHktbHGkO9x9yab3xDOn/GH6rHqlHa37CSdA4FQ+ft4kHLey4GSXBH/WRh
tgMXhKf/1XRgESv8Bq0Fnj3LW3GHY/CCk3FvUjtDrSbFODJ8ytpGu/woSMeB
5kOm18WHLwcrkMb4B6MChO8WgyUipC0GXFSqkSFqOKNy2XvvP9/+AHpfgD2Q
QrZ/Majv5eNZs4dRxIJB3yu5mR8od9UHuiZvcExT0qAmvhtLYEztCesCmsdl
N4ybRxagAUimOABOXjl16mX907QjFkZ76QCqw38wKkwFjaZYKUg0hPKszU+S
2zCEU9QRPEHwKxetlXjWYRWZfAfr1DahOhl3npczKdeDAyME8f6Dfk2A/hYQ
1iUQ2P1UL+iHoKwdItMSM0yhJ9WSz0g9tieBuS/d08QzPXfSKEUEnRxSZ1Rg
4dP34eXrXGOVOuTeO2LK+i2lOiGEpJUhIbTRKNQoNRt3R6F48dD/0RociIod
+Mp+m36jtcHjHyV2cHOBX55I4r1+dPyP6+D5VT7VM4gtxfOrd24k9UqWu9PQ
2hh+UmUm2aHT+KuWlph5JKUO4kV2k/u26TTnIXvALM5kU/NQtO2xErCnWNWG
P9vsN7hiFKk5j6LnA+pIlMAh4KaZ9lwonzl6VFo54Pxa4yUtWQ524Wft1T0S
FWA0Bjejk4bH94S9IxrTvNXcLwjyV/2ExOdPw1+93kzbjExQmkX78BgMdx4s
mPkqIHHu8lrUnosiiksn83xSXjtdQaQaIGjk9cAo8uoDiIcZyXwpb8+ntfvO
l9X+k4/RCAKVYEyiwvYzNExlYz+Q4e/XS1Q0NfkkoUJXLDGldiZ606fv/Ajc
POhgQnH6oi3ZJndzk1xX8HbXHscpc/RZQ/o4b4f5DqQBYss9e1JB/6tbkVlT
1bDuzGd+UgAOVp8tZquPdjt14k+srznsFxLAPJcz/ME66Y98vpfIJGTaseb9
AMvh7v/Naki79sSbY7ijUbk4kYi25AwR9Q99yZLs8XNXOWwHf4hg0X1k9SRp
woU//58A2a4S5JKIc5wtaegxMYPToRA6jd00G4iFmRFjuZqyOGYipfaZsliK
4sRj+hrZF26cTjES4INmMOm3RhjbeEF4uSvyA6kYNri1/1FynDrRk00MszPm
I4fSM4bY7wM1Ps2C0ykoo4iFqkmF/lJ8z/znTMnbvE2VP6d6A/oPyxkN8JTd
NpaQtPfpQOP8Medwfo8otZl86bPgT63V9ME/L5DvAyx06+MUndVJXJedJIsg
fJwQHWSWHFL9yWVR+vr1nwYeM08nFWtfE52SoeHBZD67mqM6vmLk8ZsuPpmI
hy8v6XnfiXnKqyUaBzbww8+E+KHWeRDKLbg4g4D5kMzRs9RTGN6SrLRULTCW
uXc+ZuPK2ddOUAGvw/j7WGba3AEURfTWu7ttZsV3lRkiDJo9joLlvwI4uzy5
LFV+cy4w3lkmBonJKj2ME0f2UU1XQbu7DngykPebo0l5YhQl7wOS9MhX63eE
rZRpu47tx+24HcH4vVBNOEgbvuVcTu7Oj1QWDpUPEO/NKidrcNH8IB6ba0Rr
+0FPOiR9Z3RZVGLr41vJd13ZdQzB1/DRRDGR/65EFvPxA7f32yQesx6IBO+y
9s3W71vjp25X7mUro2b4hwm6jxpV87oePrd1H9Rp2n4YrAEFjWTq4T81AU2S
V7qjAP7hgx6tYFwbRjr7fCGOYQ6aZv+Ux20LrWOItnfKLxCH9LsYLgQZCo3I
fbV9QR7l5hfnPFFl2N4XAPXWtKKul+XCjMaBrSfkVMMP6vrYHIADtDM8gzO+
HWrwrIL/G0ETEj0PbaS6ILaYKphZKsRBdaOYFFGuDZ+LAKMRRodtTq7Rd9ao
87e+RzQKTWiei62y7hMhhvQZgew+2OD1oSiBAzo5S7yqWKM/tDhnIQm+xQUT
IDNZpD1+jo0pL1afawjuPpygEQruvJcnuk+/29/eo2+KJ7EKUBLUgEw7+vz2
O9iwLTW5GbQmWmYmq8oDqZH3nImdF5PnEYb4K7OGFNbP9uF9Jo6OXU5WkXu7
1DbmyYeKH8E/FvptRHz0tUOEC3McHhWhXnereYvQwBuPoftAoGf8H9L4Xz+v
7vFZ6cVuhfSaYOf+XrJep9FGiB1gGtjtnkPboh1NAI0zd9bwFtFS+u/lu3LO
G0Zk6cu4pDQF85CVqEGiGyBtYFiXJQ45+kS/X1WTgk5l7VuW34m4sz1zd8/W
N2+zHiK4Wo84uE0R6p6BpB03jJOi6Lao/hOz7q9pPE0jtPACXEcxgs8kucqL
nl1d7aYZOpMvMKIFwiqS7fTlwftKZiLP9+f7KRUMBUAZhi9QlsIFEfNCDTeu
fjJs6wuSmBLxOfgF6A2oqXI9bSzznvr1TmYF9U3h6YhEPh6HQW6WvlNoZk/7
hVsBADCEFrO0vEhKlcx6rv9gIO4B/fVN2AxlotpBcmv3TocuP1MYYq2wGxHz
Q63tyvWPPp7rcViUVp/K8qVAHmMZh5e3Rz8W+BhVnuwZb4L8fj7V+GFWnD/t
6xCGTjhgy+tUmSSwF7hJ5AwDNEhF6Fpmx4VeadApVZ/EEOXqeGYJlXLo5SZA
bHCIxZd5zVMJckyk4ExQzv/PXAw9c4ilYx2VCGDB5alkWW/tHGK2lB1OHH4T
FUbfqdkkvvkMetiTY+ICOntbYn0Jh8B+okO0NqStsC4JkY/tLVxXiQAK5OzT
gYJXdOO0zkpXR3Qe6I4HTh88d9pVEZd+o3y8t0tyzOF7gIvRb7x17TO6dwwu
4aRZjNGMnBQxuvF8480rsorJmlzkjiSjq0WMf686JtKNpINe78GJJdKL1XSL
wMxxGdMP3avnknnIB3QltIjuAuvFNDSEBEZ+WAcv4mDdInqADH6fD7jNPYeO
Fol3fhOhNAl16gJTZFeBm2NJlx+SuMLmohH5sCeFe31BaQeKC9ImU0sEzMka
s77LJXvxdfF0RTUJUgl0Sl0FDwGaIm+Ut6Yr13rA4hD529CSMDelFUmKEDXq
5hGfojwWht+3Oopyah6g1RkwuEs0ysn5srp4IIU5mcM20xyZH2uKAi8Iqxzd
imuoMfgA36XcQaDiyvvd+NiF0YFOdoCX4BMs5CIAKXwQa7+jaP5kIR++u8ra
kZPiQs8L73TvkuPNEG0GOj67/ZLvpxeuuSs/g9l6U2+/f4JfTp2t1yWdUuBs
UW8oUyjDCY0SSMX2fqnyjJXaWx1/rulFWYTo/kssxfCInoXGIO/BZVjsa0C/
Wyn4TxSUTEB7F3WTY5XO3k57LzMyQ/RvOXhDQluQnP4UVoRAYGXJ1GIAiqE7
7/LDr3UhvsYr1j1kxEJpAOMOt6WukLv/82YzAGX43v1Hos088rBZQ3RvoFoi
KKIRQScloruu0wxJ1gOVrryWQOcTixS9SOrIu66p3RiVT+5HoBAm739zJ0pd
DF4+0n/ZxFWfqDE/pSXp8+zvLGI4DF57nH0hGXDmgUMXIuIzZlyDFsBwMAD8
cCUS836vqIxGup1VEZgUTNDC4GM40MPVaMT1e3T8wQwrSigm6nqG+bxAIdyg
uGVMSWZ0LML1jRqpsFSi4hbmMYHz2lBhrCucdr7bHRljqCIvTMWzvmanaK1u
zKvwEmFkj7Vrvaamt5Y3vCsPR0KpmpjR46ytkbS57cLuYXDov+izx42e5nT+
vnWTOUeGVUEl+J1nhn4ejgao+6Ml3Mc6NbkOZwpmRCzxGbh3+ryH82ts3P4G
HSA/tgBfk5WCCoYuRtC5JBpIdgUtFDOhxDXYvPjSXlDasBAosWywjUhqOniS
ss8pmbolnbVoNmQY6cXMioOzFkySOdfufF/yj68dhkdq5/wMH/Ll3Z/wMLOu
drQMrMtx8lDxdk2i0abvwpKOssImWoBwciT3Ye1lOGPOyuLOk6b9E4Ccn2gu
CwpicLbjDg2Dx0UCmDmtpnxfRJErZzMwfJ9ZzvLp55K8+eZhGtYDkTHps69B
Nq68Ip89uk9210o09GKBPtGRUItBSnd5ZHLwSgTuXSakksEQNDTMAQLTHnwJ
s6Na2dGXtIME5I2Oyh2GWDApMEwwxh/liwZac4i+jYKYFqYEu+eBaXMZKGTl
nr+y/2V5u618VPpX77R9ip6NdaGMUCR/qULylA2tWGVyd9UyN1DruoVxd2F5
DNNNa5Pqpl7RjDQDLWDMoKKZ8sc5FU1PsEWNxJB47O0uMbxQqcw5VZveYCqX
6CkjvmCSbNclpksGhB8Z4gGP6ozJl06yhWR2kBWHb5OthsWQQE91/9Oz9kdq
1i0JcRkiDxy59DLgrt2pqXA/bgo/xh0CfSmnq4OTzF5GVEhccrbSViWV2K+i
qu8KY134HeKoGMqWVHK577UOommXNL45+Egk6C7a426UYGl7wYv6FqVrJyaG
BMqaE5MgWocKdHx9tur67/AWBiSZoIVSpK2WDgC6onUG639z/q4AREBFQ61a
eu+lrmH5YJY4xW3rEywdQ/EcSN9qrpwsHd+wPQivnKzH+wJ2qR4bWlEUu5Hh
6JXZvhHHW9dk91CY/TwgfnggntVMqVTIYUwyv81qeCR/b2tkGu2wrFwUVqr3
Bd7V9ZWZwoasD6TVVkJr+LvZkaSwZzmD0qe9Zp4KE0qV0+BLTdi5tgixfFsH
19Xb2CyV2hHcAZRKD8RFXUkXnYJuEbv1d2w+G24VE85vvV5fShgY0UqLMhi7
2RMCOZC7uF3+vtpKrrDMTuDqxXwlEBc5gsj3xupw0yM8b9fk1tAHS0Oe0dzE
K/najrg+g+5uNTVuCXW1LB1tZPBoSd4XdmN4D4Yznu4JhnF4tiyaIJeB5Nbg
oHb5IOzYvq2aA11VC4SZ8U0AxE14cElK5idB9Wrhc+6ZH2cE+jHbOSHNzhn1
3KO1z4e2wwJxjTLgyZoEFHPmb8RvjO3N+YHdS36ct8BzOKf4eL79zDM6tikX
J8F5WGg+8OdvKJDA+nYRvjvlLTHVfwbUhYWpBKnu6wWBNHMQ8YUg+/XEPUjj
eqCRfmjA9DCstMf5+dFHTZdha5o58603fJbr6aDHgo9N+iWGG7KkNobS7ed+
1K3NlupyCscRg2CgVtn37F9z7pp5l07EPEZndDydAxCSqT7h3bYwWpgtzIT7
elMeAPcMmZRFKuTVVUcKC/MIshpWsbqMKyUwEWX/XJ3OTPNtPeRxw4Hpz/iF
611bY00pldVlGabfGajjsqY7JAu2P+IHQwmuiTNfMIvMPYk2kZLL93ozDZjW
ijFL/7XLgeVlmkv+mtXpItUiPKTMO7x76q9m67YVPcV3kVaZzYZDjiwL9G5a
S13SnF0kGWYU3o0pWX3sstFA8CAMD+6jPa8HT1Ro2v7axHMNjyGogF7V2YXZ
ybkcDhBRkvHVFzL86TMw0QpHDQ4MGCSILh8Z5JmsSHWYSOZx6d2yopUA8tej
BNsBMZGodCGcStdpbg5j1s94ZHLLWBjlsg1Kv2kRM4Y6PkJlA91rv9du8edV
pRxaJDR9LYkYiJA9oWqnJf2OP2EFxmJIHQkuYOQkFggNoK4sjAn36IKXzj+X
di3JZeVygp14bwz6yRdTkqjO3/CxGbYIzgw9g/+QtRP9krg8VAzF8395nXrc
4fseEMlTN3wQZmGikRddRMBdX07JOw7lhSb4/3IjieS3tAyd90DCVReflChQ
j6hf07CSmfqsVDolyQNRnVxoSg+16rfPdgmj33L9iJuJiDREkQQSQqRynbyY
92FE7NViqWRQLZsXu7JvFCHwS6MZGp2fYElbpEDg0HKJh4C7qdw/uhXLaI6U
UZADXWcqC4vubBHUIN9JcnYjZS+ZHloh6yxOf0hDwGumb9GX4EkclISZ+5+L
tqXC1eURbbB8WNgnToZfjHg2rAlgD2aVjc38+p8kYtnS/DkrVKYgp2z0bQk/
cTwgv1YLqhnNP/V7exh9Be0z5JyW9NHOi8HDs7reVUjpIQ8TYTAixnqu/CMt
82oSdcMj+1BHxgnUlxpUXL0KlzTL1mB9NHaeFnUg67Wty3PDE0dAzvIgDXe7
MZ5LxKAGkDgrRYde0I1V6ieP76pF8hzTI/clHvlnLpzBiPpcwQvQZep1lGYM
zb1ljuU3t5/6+BJBLR3uUjavRaM4wU1S5tWWdmhJXeHIfhChQIw1Qw7TGcXN
JFy8EKKgHjBBZemuKxSGrJsnTy0yPhVEt1EWh++IHnSL03OFJhjhVktLDogo
atfDPc+4VF8LN6IaS3SOXjTscIKV8dEjMrzQzqGjoHnMjWRh+4SjqI355S3t
M0cs3W9TFJa91T/2Zw5zICe8QPH6LRdVvX0zkRp5QXwIX6nyi03VrZfAI3R2
n0Uzx6PFynBryujiFw/QeF1qTTM86wLynGHDID/mVzBmqy+DrdSZdxbhHvMr
YNNpsPTuxbyB/rdwwpJqeKzjsLKcHEuu3ym11xt0E4LwixJOdiM8iYjN5aue
QYH/mEtd3B3h1aLP618LFEXSCz38Fe6GDxPYYBXVijLdgh0w08nlzL9vHSuw
XwWKo9s2yKXKflEffs/qHYXM2iqGtDE07WCorb6BnDt2mkdq7aA4FiQ3xr9/
5nXNrW3tracC36SSSBtK3CTAvklYy/+MnAri7DDtXnccA/CAknvTLAacEtPL
weLGLuERNwoe2I8PVmMLk/Od3IZ9tIXDlMA74m1QYki43Qcda6XTR9Awj27+
Xq/yDKfyBlr0EzegQoTZMcknvTWcu49/V+iNVCoObUZoFDEEj0+TRPAMeEKj
Scgr3/dqJRW45zQ8S8BCYVJeoVO8T+jAFSNH/k9XoUBvBA3pEhfWQ9JA6ERy
qG8QHElho3dbAKUu4YVw1YF0KzYC2LtnPiSyDGEQQn0Q6QnEM2pRi+zfpoEr
ppmAPOCDPmfTe26ApGe65s136MUDDsH0GvYlSBrrC7vL9r2bBRwC3l9b0oHg
Jboatn8xcgBPhA20pmrHvsmmacBp0CQoJyur0tx7/Y0RwCxFclbds/EhEj76
yM5ILw1wuAxlseRNrJ7gR1KaRaWmsyMruMJSpKn8hxJoaQXl0OGGPcgBT17e
+sKJ9Q/3mSvHkW+nm8SF6Jeu8cLdcYbXLNRaGGlDLgZbVxOlumA+P1F6PBRC
idzM+n6qeWDIapqQydypfXwjGlA+sJF1jijdAd8sOk5DMG+Srbx3CG9VwwKc
i5OLYLqPjLd8RYP/j76YiIX60p4U7uGNCwFGOrOUlWY/h94Jiu+A4ZK8Mppp
HT2373b3adfB1ohdATFMAGDkf72TjfjzxIZ2Zpmvxd7B24cBC9CE61WMftd9
UNn4yAAEJzDM+Vy9wonOGLEV5OzMauimci2wxkJH7AY0yPND+ttb0HsBX7VO
bXk2uDInYdjyoZla1LoZFJco8tXJaaSZGo9CzTdvKtdB47lABsLRYzOJ5S//
mGidzjKIVIvVrkoYmn6xN3KL5eprbyFiWIYaNkgh102DWrS+U3PPR8l5qQfY
B7+8IaNcCA/7IpKNDx/A6Iww6nI8raAO3MGiNyHLoAVUkUECSRVfYaqh5P65
+xaRI2MGkAwZyO4KTrBl8jremxX4W78d7SENf+EE973f0ampVwmOWPaer26q
IxM7RojFqZDma9XOLaFHmaKfTgcmfXBV/TJZeCQ3f21+PonP3CDl16xxrsV5
KSkVh191A7j6T1xlwwdbnyyLGTnT6PuoyT/dMJY0Gf37TEIWZQb+Zyyljhem
7xkzvTpJWR5PuYHgdb5u4ligx2y8L/NEYuzAsz6C5iVabXa8YJ2y88mN0RYL
gp3O9Yt4d9vKABWWQnYotlrv1BKM2ZEEvDLbonzyP8LFqYn8/RhfRsDEhpfU
gNwG2L8xiErhXwU2vtMOBZfBvS0cMT8pH+GpH/9zJXvqSJaKlX1dkDHkdVJt
b9LAT17JJT/FhD0fwEbcgMY47FqkslHlAaO6HzhhCXUn5Tc0AF7KCc6wyfQn
Ura+FcIZT2k0nI3vmBUa/KH3JyPErHFjHTd2CO+eRHfmeQOP66FlY+9eNQig
NFon3gg3FeD4Vn9iwpkkbD/+SSeH9VAU0XBBCKigPHvD1xfZI1ElHzo5udj2
mMOnnKJK9ggnnQGsjOW2R24qOLpG7dZ3uhKmHK2tlrRDZk3M7blJdrhdO2Jx
4ud7psZWc1xyvkBgnW2dZjKbLKNOfNbTV9JxpYlwD3j6CG446CWvzRKnDNdD
+K0V+dTt8FbxTsgv2H2t6vuoJzz4Y3lX8VjQlJLUyohHXZRE+OgGd7wIMtI7
IvUyEEB5SzvcvCywWpnRl8gKpUXMzv4RtrGwC4qalIOuouvW+H9vtMqO131v
aNy87rsUYN/8XNm1BFeUqltLJdbtLrIBP90jZQqZEt1qyHEB0NyebBQnAIRo
+TbyYo9wa3E12/HRyZDoW0NISw+JlntOpGv9vGro8f9ufhPuwmkIgwqH6Yr1
Z8iWpFxAL8gnR4yO4W5gviRw0vvaZihnomGBYtO7PQobGVMqtxTmvNTrJShG
DHDWblQ+i1v7flcvM2z0QN0aoaruUiRjn5QvUx8lcHohtXntvemIhU6CePpj
YAy87Q0Uw7O1QgOrvzUofaLtgLHmpdJQFstPLOgt1xTJRY99N3YPQoat6bwM
UB4mZwAw1+Mlk9ObD0/DqSFebOXT8JzCGHKX5CS3cz0ADIlVuRg+mkcGcwyE
tcPHpcMkSALiK1To0WOpWXFyoNTTuNk6cUK8ntHE/q4XBAq+tNkBj5tHrRiO
vnR6I0Xr8do/0nmPEYFffHXFmXD/MLS5WXCsHtRzuEGbS100C4I/Nde8Km3B
3YGp/ZT3lNvQ34wfNexf5MXaXo6jg6ASseVKDtzyaNP8rRrCr5BfOZH9DZaj
9e/s5S3AT2k405AeHNbaA9LcBoTIl4AU9eIIT+FW4FPea3YE59fnoVi93DjL
4lfZr2v+t3bjneNQdtjhFkfMylPbjq1T9tdU3DWAW+O74Oe2BOCGrqHreD1P
2tfZ8DPE8ZxJn+s397gd/kMVsybUIRObp0j0x8m0ClCEBN5W1/XULo5vPvK+
HMBDKPT0CAdXIZk+HWfvrxF8GcUos9ZKdX11kq66AcsWNygR8T57xWXB4Xjz
yEQMmGoyoeOOLHKLVF5eKQ7LVv4vKPe6Dpk4NDCrIMn1lOsg+hmNMwSB2KBw
K2sjiZu0+jIvPyjuPpyqa7ZPomRhQRimWxzVGJXO5+7rN4FI6QNXIwdEFkfU
sjOK+7TqWueSUitHcXBlPWfVshQNhcahOb3Lgom5fbr2Rrey27+XLwpvT8qK
yFK5Ztomnf5owy/3/NigY22ygJAf9p7KhKx3t3jJQSevHnsK44O26JHn3Yka
zArh9BOQGgzu7cMgs37MDgtI0ciW98sATPCDDfTdMTHc4oXUyWFPpMLk4uYQ
YgqD08qtm+IoRz2LXlf58O9Wa/fRkUFoZ4864drVOK9dGZ8w9/p0h0FxQS9e
pDYEwIA1r9QG8R2jAefIi2VfPIwB61QM66kJvnezwJ4ou82yHoeIxc1Eiowc
IkHbHSaaIwJ9h87L9gV1l+DXVi9NFRYdgiV+YQ+cFXGy/RkV0v026N3iw11S
kTqhJCOrUTvg0HKU23opDk81f83GWKSBmuL/fxrs33d+oH8DDU6qu/MldgEx
4STbZ7aKTnwTLQ2WR/HJ88Y7KDFs75Dm3EstNr8f+fp7Esm1yYlzwr7l+3N7
lxR7sxILK/g5DqjHr/w69UcxIbLa3ozQbHk02HokhhKKFqOklrdKfWaMOZjj
AUkNBt2jpcX5BeEnBFQvxS0nvkWKRbHM9T6xt+TxscUpT/XKT1WFmn4Lj2uY
5QSB03gm3Gqt/QNW6GvU5nBCF8h+hWXfIjOMAEIfMxHcrRZChY7KXwwGxYEP
bFZ64fgCLs9gUYPHyP5c9z8eZ0BRfVfFx31VOeGBq5RqHOV4AnRlkAF4/KqL
HmNLV+jZwVBdlKUM/kFSuMF6y7RCX9up7hcl9TGlK5CMGEfOvGkVOc9iPLFd
iSMnrGS+AtAFEekfigUyB49y7smQ1dzsWX6SkF4vh44JducLbxTyrvFbOJSt
ElEki1QHMwNCwqeKmln3QEHDbaZJldBvXQVPfGWfM0IBLxjxs2qdMgbDn4jx
iwF+cs+3aqWQPMzc8NQeYYViYwzvNYJrQp0CsLCpt4XGbh5asDLBSVRDm7eg
94IXIrWoE5bBI73/veTnXWCwMB0qsBMnvefjSitEkL80ybRTOi89GpwYbB23
kmHvqRdZC8dk6cyw8lNoaGc1YvLDTLkCI8C/DjbzxAzljigY55a0J+Qy/BkJ
025+eylw3BsujMZk3Wf5NwTIIWvCFdRfgvmXImTSqoMEcq5+GLKt+1FoySB0
YB5xglQV8kJm82XD6pC82JLJXf2BybM6NXNAYJU5AIqIn+K7Dur/Gve6m/YD
ZG1MrGNh38pDuKYQ7Ox58rITAGrft1ivERqh3pIk9de0nWKVJnPDunYeY28S
4NHuDqvzvOUMRoQovHK7wPf4cyu/ecnngCP7EctvxvC/KSndFKvAa/Q16FjK
L73Dae/za91+Rwc2eGjnuNlKcBZvAu9bG3rbn1QXe2wHLPAtTzuqi6hoiRde
bV3a1O47VwULN3i6rI1XpbN2Bt1DUGWghYdey0N3YavAUMxw8RuY2PTYUqck
sQKWh2+RGQvso8Aen+xB7GTEOfM70B1NX544sjBny9c104kRjrrcBkSaW1q1
RyUyLSpnAqWouh6GEKPS/3qgtab1nUc+fKlaBa94/9z+p0aYDLJbNILWtTon
4QTamQrd/pYaqgmo9bh4zIb6y4ZSLADf/XdZ8VAt3BkQMYeMkeG7cIIXwIEE
C7820+PEQjqUWF415NRLGWATcPRIiW5hWUOAXFqtwPoysl8JpmZLlRPtuVhQ
JQlfAp4NZj+9RM1JDw82uM2cvis/Et2fcbwOaWLHaXRtHt2lPej6MyFKLeNG
Vk58pqyHivC8402l0c3nJ9gMUVQPrQvawj+yXvUB7OC2kjfjkCy0TwseFj9G
KZNapiBTxFgyAVCwUyNzLLwca+VDkg48S+GlLR8Uqp3jdYrhAr6XzHLICKUJ
j3Km3jID2Vr5znsugN5P1fTxChEuacKP3J+H+EQhZ6t3sB9f71IjdnLaEyhg
zDQ9E9R08EiSiafuT4UxPSgdY8MQTMaY1HZE+YQ+GFAuJl/y6UFZk4c5iKkM
GrV9juNOat7ivlyDx9Y45vC79hFFA50S1uNDTeHGeIY2GDjDVgC8zKtey6pb
nPMpr8PX0lP8pAhbSCL4o4i0kZv/jJhCrkkqTAVuDfOv0x9vIfQFCFhzZows
AlbRC1sgxJWfBL879rs+9RD5jB/p4NpJqQ0RoDQUrLjlMu1C6RH57xOp9D/x
Wi3EKoolUn5NEnGs02mQjyA7XQ+s8PUtZ9HdlkGOsMiTj8lA1zOQRMXyA/ZU
ZEquZSPdNAN6jxmlHTv1vEtuisLTthmaiwEegNgxl/84+BPp9Wtobz/p9r3P
7Unz3EUHFHV85BHI3tq7Ol3S1fuXGVcTSlybVtjB9JGw38eWDINPEYVNMwwS
kckbDoJXQcyQz7laqZoA3yrWhqv7e0MQLhBzJzTZGg9hBSLjE/xR1m3oi1bb
aa3W7XmE5DUFM0NpfBpmflogdK5KFrsMJqM3FZEYPtd42UGx1NP/snloBaf+
UOUP2bWj7AvmgTcJR3UMgNHb9KLMGw3Fr2A4buTFCSB5TKBTJx8zXHYobrfz
DnLP71UHaZHqO73hVqlZgiIEVqsBIMH0KZLXbFvqKZuOU9fYVW134GRd4bSS
VBcD4YWq9uw8n8BJ2hJdb+p3n6LlCbTUAidvczEIusqug8V29STOwAzYwk6f
jVoHbMWvForPwYwqJz8gc7kQr7yaXRHXWoEq6xm4CLK6YuVtYlFrB/rxUPcm
lK9nOMQMbu5JHcpPZ9bAph4hR1fZMZxZQa9Ot+T+6hubTPzbww9qGtZl5Kbg
+Zdwr75OHOnMC4bvRkv69tVQEC+wYihxYngt21KDLTXIVeGQkBJGbLrtPqow
zrrrW3ZpeRsyhTwEi71+tDkc0KikrK3QLHKKCwhf+se+01KlggpIrIYvnleI
c6xv2bOCRsF7NYcjKLq7UqdpQSF3sGyz9PiX8sqEXWTRk1/hL8psVFm8u9OS
WCMqOsm/QYQpVz957aLUUGDZzVUMezhnaQhZR8h/EeVNbDW87INgJraMUPwW
mCyyxheBlhiGdI9ipZIGndVlZ4jZzRgSc7nSyrl1Kp5fQBI4O6Ip2SltpZpW
MblTd6Y0c/07nz3LMRS60+Rp/gCakcOHDl4VHDxq43cs8yA4jyAbaDXeIno8
1/gqRYNZO1WHnTa+mBdgrhi3o5ZNR63FbRY7RaUXzLTtiIi/oSzDQD264Ro7
qhNyiikB91JpyQ/mGC+UDhCES/JET+DCrw/O1xHDLuthpLX1MWnTYhgNp6yf
00PBGXnGt2bGn0S/RQnCLtroQD2eByF8cCj2iyLQ/uksd00e/e/CS8XolT8r
F6vyjMloTOgR+HgZrYbeEkjdaGpCnp9cKIRzM46qzBQ6T2GxT45qrbyOrmhX
tDWojePGkxdqj/WSpXj/0m6Swm7JQCd0RhGhb3ObUo20fzwEXnmk1Hp8ZznP
KkLsPFXXIOOragECIoCavC4XvFcDNXZhcIyn6Ef0AbBS+td8i2FFtM6WCsvB
zEgjR780l8sLWHgk85odRH3rxbz2Ij5DOA9Gky1MT9YFX2irc53lGD+mPHLm
ndiKrASkaK7TPQmxd5pO883LvRYojf1oVyCjooql0Xc0/nmjC18HQQeaQFIJ
zL474RJVgdu0caSLvHZeIKJlTwEECLRRMK1ZWYYckcoiQxP5O7lviGhedPeC
JduF29qAfqbvfpZl5ARZAbgwylQsEuFu5dcVA3ORhoZKWsZLmCfIbyOXpP0d
reKWOP4SlGpMkjL3aJiPcg2yrSp9B5gYEGrxGgcRd179LwwdrGQGurd7Msaw
8oRBgEjZ3SsadYcQD8NghVjCZ7ZNLSBlK8IlPK2dGfQ7fPRfyCY3oz+OkcyU
0MyvwuQo729PVJ/1gb8ZlTw2VO1xrc1PmbngB4/YZ/xLI1HTeqrw5eEPb/dP
K8de8KnljOtMTR34xWGtfjobBwPOQHMGYPH8RVjmkqcv1WMkqmAOiZ/TuFhy
x+H4NfBEWEgVmX5gdpZrfnvAO9tjfYp6wqOEm4YWTEIhyrQszMWFjzQ7be+K
l22BVyD7bH4yxW4DVbCRjLhkSC0Dad6t5ItpHoMfXaHTJwS+vz0ymGaG450L
UqUHYdDXno4U2rAgbFv/wNMmc0ndFgsHtqPbyME3vBfKci5fvsD0fxPZLnEt
M1TnWj4XiGj3FwSdOn2+4FXdokNtlpSsQ6ungwpn2N7t+6PFj6oZ86WAaqpp
0FQjUu80U17hZDTqSkOD1pohKsWgBlMMbbf8UmKmwn5chqmMmubsxmR1SWQY
p6TqMl7GGd55CjVaSG3EhYOeCC5rVfDm2yJc2VqqwYdZbaaMrUDlTBqpQe6C
fzM4ZZB/UdSD6kKfXzsLxtBUIcS1JrsCCW1ScLNMTnl34oP0YcfWW3OLzr+/
O13jZ5hyS2B0TgAoTL+FUJzfswic1yvnM57AQZyrMmM1g72q95UMGXxk5Qm6
QasdQHrDOzElpw0raGs6SgiaTSWzsamU3uUqLPS+NiWpz7PE1t7Jr1fl/nNi
iVXlRY0QJR9P4dPNN9MzsONScKTMxnjbBqPf49HP4s+2/DWSj0o0nMzH3oqY
fCorpghhS+NFJtVuhT+P10pMTRL36Qe46QpkS3KIaSa8iSPwass/lTlkE8AL
2M+1yrEygFT1F9LVtbwI/21A5dSZXHWenrLEfLmw1iw15VSlUk5xjEzFcDhT
hBdOApLTY4Zx9MYlXB9yop2f5orSRmItcWwYrkPVmmYUNWr3LWjQbyxZpuLZ
LhXxKujcjh3KUX2P5L20J48qrNmCj4PR3E8Q/463HVwbpxQLwzfED2SLy317
A9RfzdGEcAGSFLhl8lhlK59bDABj2Vjlg2kqkh729uZj/pi8bv0zNO0Kr3Jx
jt0x4RAiGz0AFuiJ2C/nj0KCyZTUIVJ7dkD9KwiBshWLXINrrb4t5ChihwtP
ZOGS+o/WzdUyzYykWhihUIyUTPyQzB/O3K4owXHbTPwbVIx1lxY1qj5upZSW
VPWiOwhG9nP0Bf30jN5QW+PssiY0S0q2QkwpcYLOb/KqAgAidTWi+KpgQG8R
u1AQxSrOHu4hLmVRPwv/pAazYSAVh5KbmOkdYaNVCo/hSZGZJaBIBTs9wtFL
Q/LuXlrvk3IIxCyzcnsA2jKuH1LN/T9bFARzLTppJIk6kgSshkQ76D0MgN84
SJO1/VlnwGkyPx8NycMFQyf4QsY/hM3/M4E94M38YwtUcFUke24D/BNqBtKx
EfsusLeBgr4PIk09UlCfmlVqs68l3RkOdCcebZk6dcpHH1U44IYN/PUAkXj3
a5PPrhuMkAB4Sq2S7ayUQ15AstzKdsZBeU/x5ZX/rq+QxwEams3hA96RosKa
Yx6H9cxwfByDdqZ4E2m8RozBrc4hTEYsXKgY2Z0H7/7kXfT3kSvFbVbOpVGS
RMQT/0QltVw+3ZQX+n1tdI56DqV3r7GqzsM4vzmyUMkXJrw0gyPT5rXLV5Z1
4eJFga3NPfYSuqbjNNUb4atm8clMBwTlElSZfg4oKEirfM2Mf0fid6/2ht9Z
cILQ4KQ+qAGUVSqp7hOcWgg5T1gpQF7uLVmKHKmnz+7STvwpe/a+CjISs00w
GWJPj4L14dFSSDw68yIV9FOTmgSRP3O+ljKSGQHUo83ELssq7lMzTmlQiIDT
CiZtAtpy8nvG57CfWvM6rUjXHMXn6314PF/Oj2YZPHfWidYrkIA/zrfvSmAI
3iTFWUdUOJU3mqY75CgHvL1P2yKFjoj/tkJFHneOtEK2v6CZMEvKnqy3jlCv
2rCRN/cq9sjHFA/nNx6pk0tty8Pp7WUx6JHdvHfwBfzze/phHUPnwn0grGAR
Cc92bxmno2LVDpjyTBL2efsoUBCkeoy5BV22W2l/BDZo0GeXCiCKNeu6j+n3
jOn9NrmGG6+DGjjxsR8iLGP9MAgOYY4Goj9w7CHCLYARBAoJD2GyvVWMcn7u
156zRdi8+Ho2YqSRVrUBtmS/tK0IICo/B7tB1lQqEQQ4AjCBXfc55c1qnzr+
EV0jjDpfrCtA+mzsMaDMcDoL/HvDt9AoftDfLW7CTjHCVHSeYBPQzFFaNAcv
8QdSMaLBnoq+MYi0OPeaJBZIaIfl1y0EL6RjQnYo0FoSmd5IxOOrAww5rfuD
MKczfB2eEt+4vQcmSWLIEP9jETQ+FsfYS8y739sopIzQeWc1dTSAdM4gWRYx
zQB7RH6WdER0+TwX0ukpdUS4NnSWMxPyAZzONPAmBP26eiO0Ke5sCkX93duY
ad0u8YZqjSyy9T3Os41UgpMreiZT3iqoT9G0BbH+k/uDx57IESdzW/qk6Fdr
5Gxh3b7FEpmuJUnWMOfmfYpyvAi9JWJLAO8BfKfJNl4MJheAeRqJQHKVJVKA
Rd/WxR4vqIFc8pOD9o5+wuSGHPnABCYZRZH0YUbD1GYcei/Odo7blufMModG
YuIo7Orh3x7tekFvW73gOlozE4AQxgpJi6Y7i2Tmh0OWpTV9fej/HnuWEFnD
cdqhdjDKZvFfJPsJsrrjPE0NV8eb0mDnasBjkjPX9zAENVATVKk9I7DN87lr
wwxLz0hM3ND5ycUvBZa9+tquCQhpSFWP2rf0x82TWp3cnDx+QVm2Tflh7Mf1
1NAoJNGHXKX93UCfdZfnneT/vu8Jn684A1LSvZnvKte5VzGZfOgKL4lacq1f
3Tv995wXhhFVfN1zzaT5ufBVy2JbCr8AMnsecse1nRXa05hU2VytfvbHk9Y5
sd0eru8jNEQIHdDpjADxGVV5336KRw3nBOPfxDCGZivY0J23r3TaP2eqGHhN
q8sje9OOv6724uyWjRuy3yoaeQ02tEGWdy2wm83RfkZY1UwY1p4AS5GVen/G
HYLy5F/GuYjGiVzvOjlnqvwy2u1hn7kNteqA34ajdBscWvxWI00thCh9V37q
MmzLhNuOMZ3VydxONlaN7y9G7Mahq03mQwQRiMOC1ctRY/bwzXVfq0/9+vuK
XGQNB3atgtDh18WrLwbwK82ziB+yC2Z8wIiOb694ikPEXr5iLokcGVI7tlfJ
qNRyTbzgpVpz+3MnH6HsbUpRBUbHfI+A/zLtrBJ20ja/L19QvnA32BkhgzAb
Wlvlic1NnLkQE3EUtvx9ANJPEegkbvF6Bdjx7C4KhF2WgzeIfk5ev4s8rW6I
YFOVE5Sac2cLQOggdh9/Pp+DDpdqkvSVbO1LHoyG2e7vZ9XilivAre9no6eB
qDpWif5FUdOziDm+Qw70zRskqfX6d8wT774YJqGOav43YzHL9BUX+7G6ukDC
r1ZdxfT1Ro2WK8/qQo7GWynEBS0EiOTeRPNDOBkm/ECF9AEcdCh2+kDBHTm7
JCTdTKkinclu3H+vuvsqUsKZ/sPpXxOGyuw2jj2dwTrf+UVJwQxVMO3eamTV
npGQ/3OlumOt1xoHVObhLMmclqVBLfwVWllXmVUESeO0qbIDTehCw1LnD1XN
pyUGYgXLwvLUkWos+tokKHItVh4WhDG/T9wdlq3RR8wk2f5SgfllyfdHX/Lw
6kfwOZPKwdKmPBDNy4nvVhZdn0PvO4XDbYRMynLg+DUqR4E+d3jwb8Rnaa0K
Un/3Nm66C8p2I5PYLyENPoudmMuIRksDJ+C6TLq1ZpQjsw16l7aoYWWk8GBX
e7P/J4MBBKifdF0VwvMk+M4pQrsXbm7boVtA8artiKR2pip4+07iNqdzadiD
ereyTlv+OpUI9LMz1W3XnVeGZW3h3x/IliwYtTAjh1HexrRacMeTvdgZenKQ
xidDPFzRDkSlVUZJCYM09Za4Ze2RNrv1n7Vz99wwF20gqu/d73tOGt0r/sF3
wVma+/vWNSnp59dDk8DXyybYXxhyFXnxWcsMUOzb63ns3yCuw4VIuJ1XhGQm
xzwturs7j4Pi/RrhwFgDnmHXqKNZqKhZYTI8C4swtqFi4vqEMfMlJRwP9Qs0
H1ljLKblphw9LtSframNZTOlYrgblQ6na1VjzazjbHQ0Ie07fZAJfOATbapO
IRe0J1WWd8VB1C4L0GlT0LMvwdk5hSsVIxAr9eHC14RqC+0vZxcypIOnQ/BK
2sNf7g516qRGUjdHC4PaIRhHktk1tD2pm5jU22xiZ8zpJNZ5mPMapJ1lBhQ3
G+LIzxubkvk4N9QY660OHU3P4om2LyWa3D8XfdRwtTjNI3mv/YEIK/HwSJfi
3iiPmGo1K8NnNE+2rCIfbbgsJWKoDf3hUWXMATxEyFo2J5DEqwlIcGdNshFx
k1oenBG9x0+ht8lnJtJ5ADcRLOaaX2oAYzcTXXKOZz51jshlPdPHJj2JQDw0
OBi3J/iuxZUIeqWAeHM8hsFYw3IbzCwh5+E8zIaFwSYccAnuO6aNM1ZDPolp
y7zIZ2lizEgDph+OPVg6eSvGlHuo3YMcmf/fsCQIbulrmLEpovWD5aokDewK
yyt27H1PrKBbGBI+FsaczRucUZ+Z/kNQee8VDegfDOxWynUN3awwzzq7ka7d
Cs3Q3ouL8Id7Bj1FkGUfpKa+GdvFX6QNKdqEd3E9H2TmYFi++lU+mvmR1C0j
8VTbZ9NwXpGBrlvRE7NYGR3P6WnvVhyLBmHeYnZ0BM0o15gRts41Bn1YmLsH
+QDPmwsK3UTRbhBxkXfeQAn1VbFD7VO84SDi544sOA4yIojbxDy1kUXTHO21
79hMgWHnto6d8RcQuW8tSuJtKqse643X8LcSrFHboVRkkl8oSiDEhp4kNTu3
N41t3TQXBkX3F/I6vl9NIE1KyIZ1BLpkX04b3jwemdK57yCpbu/gnXmqcrQf
KPmaK7/5qGYCQNdEQIUMEMjazIqdKDzyQOM+RMUHsldTLpMdw/i5AjkzROrC
y1YyeOtjzujSl8sxgugzaNQhWHm02RXUcL+dwmeLIbTV4r8OJvMcaASF3Hmj
craq/qpTGshFrsATJWGulR3sz9j3ZlxXCPQs0gp7/nJx7L39mKU83xGoLY1/
S2FXCDyXbGQjLXofS3qk+0O8JsKU2VrpRgMdSj2fXX6r2M0+H56jx0PzYtzr
hTySFY+3/QwuUHwb/IRAMb09i78oUe2mKTf7raccm+DMYGQ1SZyFMZY4BzbM
0kHZEMcrBfxa/nqatwbv3+mFUkoX+K7Vau9kE71Jexat5rBTMmxf5U4S1GaD
RcUz3l5zRbyrhghzIFVsu/JTeAqXmtEdo1w+suhQRroX+eKm4lhuBMTZJvIK
nWmOREPk52on8Qt6zcfs4ATvmaLmOYSxg/vre2exuZMyZHU4oOsS1ZXgagud
6b2cJRodjoxlLonWwsbEytgv/dXbeDpKr0UFQFUfyZQLQD5pC7xX7gCGK04N
jZ8PQK0EKjWrcAqma18DHJMHyswpiaZDuNx9EmIeCHBIYsqReN+OVKHlpTuE
yLFeBogxvJSU621sKpTpwDEBJS76NbYDBkAaN/UgGt7pDzQSf+Wbd1Vr91Oj
e7xzQRbsgPwyVDiXVJz+VDdyq8LidkGGKKos+MG5lDidl1iHY9vEm1986uJ2
ei2J/vi11HDdC429nhhelyoBNTchFMViibm9hyp/0UQSodgRWoPRcZo5Ktbg
1mrJiLAaIYCrhWQfVbcGtqt4nkLNjsvG434A3yvDIQ7NUmwMsza3eHN+zP4C
4KYtqlUxwOScNff6NcMpwD2hJHrab9wsay/5PSWVW4LHhjhJ/61OVKlKiBPW
gfpSV2Sv19sN5mogXBkIls81W4FwZexS04KR82OK/nfJoNFlogqQjx25tpfM
03yTAYUOTAziA3suOMJpxQ2DedZRTVxAEc7YCAAjbP0gvLQqpD4WB6uXX6F+
086+djQepsTlYbXyo3jJPtP2oCwBiSyMrE0+Ei/yzt3ua8SacFkKSWbU8aFd
i++meOJUfTHFuKxac68gnThiOneM1SN/dWIAk/A5EGvFIYI3e8626DKz6XoO
R6Aj04p8mQqwfOnjPA0tKoLL1tIXUAhmSpaJ2LwaasaZlVHGDW9KJ//UFcdP
LsEakcJ0nCNFi4sVHc7Cw1RPXRKhc6h61xdcO+pgxGFjweW0vACdZRPbORH1
Nv7Rd0RPRAOsNjgBKzxrt0B4CD+PoKSzlH92xtCmP0pejYJq7FuGdMcyfLw0
F9lTSkDFvz9qbdNCNYWmljvQj+/W5407UNylxEyVAT2i9gik7bZNfFyzY6YF
/68bOb69H0Zqh5hfHZolswO0/mqahI8UCSlzrWAZUtQGLEkumjyleNkP9tiA
VKWtescyG52zEAoBA25hkv4WffqKBY0ScP+dMqC92znJGG0aZ2qct+pI4oRd
Z1a8M4itGYzjRm3HZ8WlDhkG40hOEElLscS7gZmimMLHCtOAFNOLCokL45r5
CIvl4lABpOTMAEgb5Ze/Hii4Kr7ztLoNAfPjmx8NIYFqBfGRaoRFIBSMvzCj
Z6HUkdjrj03u+IcB7dQC3CdK9iJxrEZuSH/mMgmL9bSaEiryUZurVZlOzOKn
ouec0lYZjgJHYHDTzmoRIn+f/kHCmT6F6ICr83NtFJdL7Bybpw3cvgO8JlCN
6myG+DQ5rneRDGzHEdsmZ6mKrmw/BZ5mdVApyS8ySIWveXbSx5fLAqpKOX5H
lz40ebblhxf8wuVdfp5TabZYzTFb/qxnHW/Hfur4pe3i7ZURZEb/9oqwlCuV
R9QJr7Dff5TlNaEdaScjGag1XCgsLNCIZFX7gXVJOpgP22UZ+KWPRJlzImlz
0r8wbZNPhP0zy6UbcVOREmGhsWWoLX5DvMJHBNIE0IEZmLsVV7OBprvPfIrP
FzcWyJXq3Q5voGHwfUn8cU/9hPMhCw24RcouwTtTAtLfi5dJpeCdRX0xBOb/
laxtishEqVlr7MXexScy+Pwpig0fU6kcLbiyBum4bgT93i2RefpCLDePY1eC
nYSqeKWdGbTF8DtwpWHSNGC+0wxy5cl+fXlopmksEgoqOGb41aVsHZMgE795
AzGU1zCsFpx7LlBrar8XywMzR1wxFTDDuUUDdTgXqqjlhepEOsGhW18xa3lG
Pe8qmoJHV/FtJUEyJ54T1HSHnVT95HKllEdhlX2g8/Ectxn9UAxp//Q5rrzI
jZodijaOD+2OOd7SdnraTt71a0oJUQpoo/LiooetrIujVZ6pykhmgLjuW7si
+e1KQ/1boQec1d3riLkFtKM6CeEijYGGJDH3/IRrHzkAPLtZxQjecn6Q8LA/
Qh3+Y4f1EEt0VX9TDG+VJlZeoKafQ3NMG9rPwjU+hVKL02sMVxmpdD9yv2xu
dC1HEhSBiiZUFdNPjRmIu1v3QKGsGtF0/038KoiKWslH+WK28k0JMNCrf029
z64+tK1/Fk7pDqbMuPH5vSGKAEr/SKExfJdPbP+uZlOW+GsCe1t+xUebcQJj
WQYBLZTUnEhogdeksAzfEEXNRPNagIpav2Zs1F3Yx7ofUSxCGqw2CL0gXnY9
dqvKolmPcCRbOFsMUZGhokbX6o5u2oayJKHJwmIIuSueWqq8OJLpo4aRzcEH
qSN+ADi9u+dDIVKWyqH8aCmdroBUw1O7nrj2kI4TX30WWW0CGonPX2vVVtuv
LJw5Zyxdl3IwZqQIDDTqOz2TtfmN+cz/FYEg3nHyXnU1PQBAuXmCuT4HMMQd
0j/y/HSdWsCIsxZqLRrk/cnjzO58qxYwhi+7LmJJLjTJ+KiOoYQZSoC58vJE
XIkAaBsjoicX+jeE6Xw43swif1ssRAAUZ8mgLQ7ejuABrpDefPfNA6GVyNKy
ZBsPUAnSS8bzxscznP7P3y91I+n/s2jZ2p12dXUGflT0xzpfFno3RhJd5hM2
JWi7sHCX1vJWX8IMiMKxqCShAosp+ac7nFtJcCoT/MV5KlvOFCX2zRYGkxoF
goQwPOloINLHvsjg5p67oOLWwoVCLFiBwAMgFujHwf6QJedme/pmieBkcP4V
d2o8HCWV7WLm/kjlLQ/Jlqwfz8asjF4rLKrY0bCO9ijtE5S+zR7JEyfHmE95
JL61JrI+3Vxzs3UKpJFBvTAQ8qYIfGiW8Ku22Yr2kdeom6AFd9AKYVoRTAQi
eAgzX4BGhiwc6IWTZPeZjw7ZLfIO8+q3hKDpK/0lH2GCo++aFVLatuU9JoB/
rwaK5DsXhtHPqtjlvuSFRq984CWEVqLuEDtL58/O9OA3X/A+Nb7rRd+dqah/
/L47pfpAgk97oNanRxsY/BXahBvYAzGgi0kvv6ngrcYb9nEb0y5qJoae9MAJ
YCuFBcRHNWfAdk9W4MmuTSGwwPkCcry1yLqBExDbArIbMJMlT7Ge8MGJLbXy
O/mFt6sRTngW4vMgu9Ix1KZqZN0gFZ6BaGLPtDFtdXfv7sn4Agv3MweL3O+Z
zaPIWbbM3mbNGjOYeqstIPfyzgqOMTqLFjuVHw1oih+TlQSLM0zJNZqsGo3A
6D/I3lITLrpKld5OmrB2etoJ294g06R5eRlaCyHnamPw/lBsEv4lmGDVKM/b
+fKkAbJ4xODy8hjrUeztkF7YvhwcTIpxBx8nwpl1A5cAaX5gJIsnkAdwA4uR
2gZ2iNEWp2d2zQF8JYnJcrPvVZWmQJNlhBS3N/KT6q8/TgRGL+/8WyCDosWh
zkeA3hg5L63Rfc5V53fd2pAW3h39NnmbRpW2TUAqQh9TsInI0kHvLwv2LQ7f
yvRs2QNgV6/qeOo6LZTf/nEmukfuQdT56AVmHnsyha3FkzBVy/bYGtNizUXs
adkazoU+nr3g8Sdj+bXngzZFT9Kxw6TXgQ2UQ5w/TKXMai3hv8mreZIeAell
RGNQUvOdTg7tPVx+TGUkDxb2fRMGizBYdtr8t/fkeY6T0iGUTFwUg4FvASsH
preYW39754vdJOcIv9kQYTfMZm1I37h6k8oAdIaARhISZN3vMg56yZg1WBjj
ZytHlR6zFvwTWFx4zEACmBB+8bxy68XXfJQhMFiRimaSUHf0IdGyUpYFZOO/
VzB5N6nmRSO2ChnYu+mqYvJkBTiiDpj87KNr9qYcaYctc6VA1cDSEN3ofMtM
Pt2gQr31VJWom2I7CcLjva4LBSXmzjFX8bqWN8tngaPqMnwC78og3p4TE5EM
1enQiPKEM6KehZjsN51CuXqxxY/LpadticjZyfhEPonm/kJJo46geWVSsA1G
YH2T90eKsTb2A3LNRQIk0WywfqFZxZ/tMc5S146mItERgp7z7XXLjlNoozem
LIHRWA0Od6qofcl3oi9E21HEZNsVh/266TvGeLJMYXEzI6wwXOB5/xjV8Qzd
8Smv+BpGdwC+u5SZC/T87VXbVNdw7p5h420r2b//g6RRf8taJJKtDB1IAa+g
WYIhpTSLbNwjoy7cnqCoS0uT3eSOai2TafVilwvnbUbzh9ESVqmUrRGZRx/M
PGGhdmaAt3K8oUGZ4NiEiv0jbJXiETl4FaMAh5c15hKuOvZd2MnlQBurm+oN
iQhsH2U4Ju0tuvACmGOIxRbdwHUSlzJhpwWgJsxh/g9CqSDEY8NsDHJ+Emcf
1G2X2aW3CMh1hCktinrtm3Pod55TDv5ROu+VGsf2R9XisRMZTJjzwI/jT3Pt
WhTw6ERtJRS1KYnOhnuD30C1wtpDIG0UVatOW4Gc0s1hC00tQ7C8TxDLvlyR
ojDl2YzHrzKkEGjptbfOTkdfkb+qtqV8H384/8WXztPNOOwjldLsiC6jEb5u
3iVbE2lHRn47oOOniJYr0emtn9XV/9lasebObCcGY64udiV2l4d2vwxHqS4e
mtTawkKohzHcIBfRZsklU5QK/uSFFvLaxbOfn/d4k7wZ9hmGXWlg+lDeKMEQ
TG3OfO62AJJAQOBs4W3rswTSsIM5Zjnp3Spr2aM9PCzkqq2FU/hIhhREm6V4
AfpFfZWX3lAHjmRMU8w3tBaqY0QL02wbOTMB5qmshU4zfGLOr8j5kkFYmbik
N3kWglPXLNIPZr4dFJ7yCD7y4gigLi8T1ViTnl5N8SxspIunZKP/ZQ8HrIMI
ozFYRYo+l4wRnbBCjVin0DZrwApY9S9FKSCSzgAs9juY+TJAnuNpmLonxRTD
kEUiWPULCcxirg5SmIzGgTCHNViTXpgCcRhLJTaaAmPdZxQz47xZRn1wU6p0
QbMf2HH3VX8W2MEgjS6ngn+ZXNFswOPYUvIV4lOadDbYE6evQJhRJpXdM6Pe
NaxxNQxqhawY6MLv7PrLsk7HpLGoRa7J/8NcFprvHcLwJos+JvyVf4dmFXMK
qBTLfGChI/VyGm32lqeaDt3qnSXmij//NfZym8D5woBKfBMxrtDLHizngW6j
ddXajKVEr9bjGvo9dmVRvjedwAXQRXQY27ZMlZUXDmYuv3sUpnKuTt2IPAa7
cF/wmcVuAFiSxFQVXEFw6LEyT/05kb1NkZsakuv1gAcegtarjlCCt/XOlVLO
70jI6VgfBA7uyVxv/gD/3ipDAurC2qDAYbr/9K2FcgOb5VxJDC+oTf+bl1AZ
7DauT0oUCIYctpX7rfhk/4lwZ1Cjykb1QIViCgEadaxPkTdYdipWPkA6y1h5
NFOy4KWJw6H24RZ/pVsYTH/ajg4j4OH5OkL5vVBCFdk5yVGWJ4Sgx1ZJPDD2
DqHQ8Kb83m270mOx2AGbEQ5VYzqS4umMoKTTiy2shxekFhIcaNrmOFvOghmP
DNjdulD6/gjyhMt0VjS6LPZncw2Fo2ehNLgBHDevkc2yJjS7dqMB9NB+FeVG
u1YhzXCB/f3jnVBfBvmenle+xrYLIMQCCk+Z10Q6DhcANEsxMm7BoJPOYFj7
hFzPFzvPRdVEEWccH0U5/M3yod2qc/JA44wQ0PrUEp/qjQqTKq1yZ+23vcbl
Us6RQ+K+b/Px3zxLfHNp7GTT6Y/TkU21aw+HZjdIoO5cwmSTcf7MML6KbJOP
aL3H5sTOMHo7SS/Uz2QWDQFS2XAAqRUhgQmSFN7v2t9wLOg+PLii1bTAk3l+
9oSazAV1lYsdPbrr+Chtr8cPtB6I0/KooMC2nlrG0uEgUKjmr6JwHgeKtWYI
lhq0ESU1i++5PabQVzOMtCO84W8Lf9rL4cH0RxyOYJ8qTiAHvMe9QIxFkwh9
vr2peKpFDNNMYSPzCixIDn5duTX0WQ924roHIo2rVVnvkeoc8IEuecWjta1t
XFJolZ0fMM/wqFBWDq4qEOLqwbKQv1Zw6DcQmy6ryopxBEoZWcJbq86NuO4P
lPGTSnu13FW4Z4lA+yc/buVFURC/5uk7bKUjWRJTOTO6ihnlSmDnoOBRc36B
YEqLq9ooR5Z/VqgzfBtCa/PLEWK15j6br/p4BOLsUXgjf8Bl10R9zhKsZxKa
3pSzkVKrjITiuarfBfY2OCcskNwvkWArlmbwnsARIVsUXFwQv2bwe79WjArM
MYh47HdhhmYeNzFVTn8+wGV29Jxo+WpTc4DYwIzGeFECOluGynb24p/cdoad
8enu8F3zZ6EthSc/xV8zDSsnUsS1UOCxCDUQhNL8Mdj3KqP9/2KEs7aoK5Zy
VajfjO1vIqjqC5DgELrTjICkiFqPRc21t6vqH2ZXk4JCxBTVZVZEtBEtybOr
FfhDAMbxNnF+aglvVy8PYnBzZXVLnvUjzUti+Mp1oaZfvuBfT0V/Yz2zJD/Y
4git98YSJ5kGsJSVPYM9n5snhroluxaplk9cMPgiJh4cTYUNqv+mkNWmof4A
CmuabRzaysv4OnbjWtY4aLHhmk4pRh1sNDunashkKxmr+rfRqVgV4iZE6Gjy
hxrBa4bkMIHw3nBSxIyF3KaHX2+HzWgmN3J2q39Mzcg7+3duXmJhwiT3B3I8
Wx54OJEGHHLwVbkpGL1by8lNAUmNX+BM8R0UBeOgdONjY1N8DJykJLTfgEAY
U55BV0gXKBbT8S3hQLYS0J946UCoaWKD7wVFjyB/ksiXGwIXgA6/TrluONVW
25lt5EibQML0DR7YcI8QObyPjC2/WQI96X+geA+lCyihrWb+vfLp4psMjOhk
XZk3FRc/gmDF2GYuTAJ+qviZUpFuo+PAnwGO4Ak9iyWaAG/mc24vfjE8tg4y
vU+4jZE+dYddbWTwF4fdu7cCDviqK3jj/o6rJq8VMQa2riAKSGXB5kM1kS8q
Vt2TM7580j1znrjWKX0IeW46LzDeWL1kXbZDYaLzFO5ty37tRmShbAA2AnD6
WiDgj4xhZ8Ul3QewSbd+Mu92cxgimOoipm1AIcOhToRtZNPP808ZXxjPO3DK
QrMkxv5HuCEuDrbAdllTsMu4sHZ5dgVboNwXfjXnBILp2933AekX8ws9+FQ8
WHR8BAx2vELwAONsfE6MBtqyLQR4Dag58K9jPCQHaeIsbMUsofXr5Slo4xKw
U7V6BcnhEZTP+DjkutosXOPdXf7OxUVaEBc4dUrx0lShvIJUOYIrn+L6GyHW
h13gjVfF5OV+nNREoeVaqWVzMNVIlv27HUFukOEq4jDZ6oWMz6ckAott+0ku
X4wSU+A07tqV5rO4HAug/+OsQ/ocO9BUF8uAmEUgwW8O9U+iMvgA1T6HyQgM
MD4PlTq1sKbaFW4HZjdYdaWltyvbrBbg1YZTNgtWjILNjFix5QiiFzRFyzCT
E1OQ3O7/TWYjmhn/7snUpUJ7UaY6i0ye6yRwRdSEwsMvYsB4TKzit+vX2n4i
YzgRig9VckuaXOcCUKH7oqZd8JKe85cIkGoHK6r1zzmZC9K+eaLRQaaldWHO
VgOWFxgQWPkv5uaWgUq7LPkfzzyuJB01ytIynFHo8uX409OVY5GvW/KfP3Ep
LvQmFUFa6ZNJ9kUEhDtox/gKlnSNGOpWEkq6tljp70Va9/bFV13v2pwFzRen
ALX3B5gDha8CWAr9ytt/dpf8Y8oYj62XgB9psbkWzyfKz7bGaQZ8sScteY4y
78QX9pBvbq/KBaMK2sm2FLLPUlKGZpnCnaryT50KwAm4X/7FAsey0+YIVsK/
ksPU+uEg9oeUy+5XWwTOCGwzaPCsbCnv/rIQN+1g9QVcwOWLpzQxQ7rX68Ti
GcKaxvCSjW6/STlXRVbgc/wz+LbsZXi/1AS/wzo0mt/B0qBhnQo0lDhI3t+O
hPWP7Mmki85INOAr2lXqqZUGR4GeagzUZhUTEqSUiflSvVf2gpXHCb9b8RqL
wI1Zf2SBGf1FwvXv0P+UjnSsWkft6QN/s40Q60R7zHrrekhRMVVGHGBpMuzG
K06D9SW4UoK+d+qlofxYj6lm2i3igtNZlFB1uPuSOFyAGeg+itLNNsA+Jfvo
C6tf752ZVBX/l2Vqpam2wqhGeCJqynqyfD+sStfHJU5isJvc30Th9NDf5gBp
PwF76kgOPTwMWUiJe/CQqr8va8dxbxhv/LbZN5JFHbUyC/g+Fm0MSZY+md7q
0Bi5aKKe8dWxVDjOvuZwAWx9HhQERgsc408zc7PhfI+kBrbPdv8o9GDhEIvQ
utx9ouejrDhiLA91jCavN08RcLaIMAXEqlF8zR+4Y70gMlxM4JZFiq5IDHt/
Tupg5I1xPlxIKLla0H6ywhCDC0rI8GdpYd40gPOpKhiL174SVabYG0WEodsm
3WXLqofBphHxVYM1NDNW727vWX5ifD+Nerx9Qebv7ZQxd0Y2W/KSPoZskGAf
mgbp7IGrhC3nEaOkPSKSPPBOMVO07nuO+EXQu3Ud2eGdwwB+CS/qRrMezTXp
ppdyJmMf9jMJEZg0DAavsAldIaDaTTeTtCL+YgHBM0g6z+MxCO3X5v/ZP+sP
nGu8RJXzZ4TdK9DXD+C/4XVj2bKsWL/w90ix0dv3mcVziEmT+rIlJozCHKuP
srt76t4oIm4YUWXlA6p9f5RG1veosFE3BiT1xkps+tH11t09AVLDTHVn9hDg
7N0sibiODXPa7ZHv74ZNNkrNf+aiS+ib3F07EtDaQdNEtoug9SbMoWJlS7LH
caekFEBdOYePN/8WEha71YXNos3lhuGAXjLdvThgwkzBvd7+OEDPkdMmmaqP
y7csEOblemRiiUGzJ17eSEaXwSCWDvwlHyvbn514FfmANPd3Bbh8v9Cyrl/b
l2GYb7uVErCSZtcT88dAsI8xeUkQy/h0+J5GppzrfpqCiFJD4kjxkJRZ+99c
lLL2ZdY7eVXEE975deC5+O5ICu/ViqmLywRHLoM6ig69QYu5YtOKetv769uK
5mvlsFQDUtpAzGlV31syKwOQvXycKiHIVOT8kv2ntcW+diGJk3c17WgblWqa
RHKrfeAFYYd1jN2kUqW+SIWJ5vxZN5cSKf/0SSTyALjNvbJLAb2DLDznswAM
36cFLYGYPR6wORpGoCeYm1LkJf28dE4+6sdhPinJWfUGUWtkoJqid4te6bNK
dEETDljL/6AJyyk5ihIVKZ7yW1Nf0dOvsxVh1bTWdCj8aJcuTvh10lwPspCN
Q18609h/XIysrwBA9wH47TEz21tYqDAyC49bj31rqNJ6aGzKj++69AeTw8P2
BYsFtwOyhO6AHgcFVkai2r8xOIEE+ztjAS5cGMAZ6knfBO5lblkQFLXFq9IQ
P4X3rI12CLl/XcHEPLeNct765RUMMa3LHTPxNE27q6lNlH51SZzD3J9qQg7x
iBHnN3PdfGtbMubLZyEmYgV1HuoRn72jTWCOru1d48pqR+uQnqqpgITme5+k
EZmVrA/WSUVtx0dAYOpCPYMs+kNhklT66zV8DM5HCHsfuieJ+toiNrO/2EF7
J1NWA1co3bDsO4n1q4/5+IVpvbwZNaIz4q19xqxqk0rwA2212TuWQzHZld2i
56p4NUXUXOE7H/KGN1wL1GDmARmr9GQMy2tp/1PAyD++2Mv0DeMpYCGgdfDu
pCnjBR3kIO6hmFbKsb9q34RqBdsx+i/clvsUGTAkZSnzl3wDyA8FQ4yM1j/D
l51ScrjGm2sRlP7N+ooo5wy9pITHAWBFKNjfGUhx6oLeqEG9r2959cD59ylH
ghwJ+2+d14RFIo8p5onHqXU5frEISBtmAQYqfZL9YGdkkDfUK4h/s4wg7Jw+
3Ec5BhDtCMvkinH4l42KptHCCxyPmRwziNL+Wk5Kb8s8RJnpaWZdBS5rzRjr
58Ndu6QJ793hIbszRlmM6C6PKvds7rJTIK3TGZ5qV8mDsXZAL7g8JZtyedIp
/0tWjkSmD5qUL49N/FL+xeWxs/hR/uBQWGo5Xt2pCF3uZ5em5reltULS7+Hs
coOiJVodmRuZxUrZaEk02XOdj1uFl3mc2GNdM8GiSF2lEWJW9mBOD+KA/VX6
nbwMiKBukR6rC6NOnH7QQHiFw+iXw+LT5S7Q7VFubDcU7UaxCe0r7+dILS3G
JLoolwdWaKdkjNgG2MftbhfUziO3rB98OR4uAcsPOlmS0mel5Vi4zbBioMic
D81+fhn0BpX8rTPtMmTyq/8aKVnL6puOp/2QBi5xcadYnwZuniyC11MOEZh/
JpmZnielbi9ceWS5xWKP0pYuLXn9BEesoSKpOC5eWvbRclNWJch/u+wKsm1U
2m89ErsEMcluGINHH6VSbZ/n4uuaPxmrJJAcj0HCBvqgnZYvb9febms/kbDQ
M/kYJZNShRkdkwBfc5JqCrTkyFD9Fedi9Nq0gw3f7PE7h90O5j4FEzMA7ejU
AZZ82k9zUXNFnHDQQIEqjEDkV5dFoTJO7yT0cJMHIn4CgOzTcfu/T9Mm3/yY
4PNuXsh0mFx7EB9wvHBlZlThcxtftnXwLxFpK4nU602NG+zf5bHckxdaHhqH
o/8FrKjT4gjwn47PsSOoNxCfmYP+g8GySglB8cJXvqlwLqcpgbM2tEzu2Inr
7ogH6jjUQ6cD5tytcesTIYgAZCFFrh9irxMRX0w6JT8c/B/IEJ9sTiBDWqq+
0fAbZgZw+2H0llePoMrwnp0rJjws8wjGsYGwELD9AwEBUeXAtWUq/exI0Lt7
rB3K24gO415aACy9keCoru0JViHrDP3Cc8JveGox80Sbc5veNAEcH7FLAPhA
+Qu0hNqRNq6o5VnZ16aGAlZUiE7GYjTW52qyL8s4PXoxhj2LnQFDPIk/nIEw
01OlZB2KA1hj/mK9u7Q3BT41jek2vaCAtIyLeBbBsHkKOzoarVNBYQoxo44v
fnX8OzBS3yY/SokMOa4AxaQutGEBlaFjJzamit6LWIRl+j+NFYLpqgGkESNJ
JZ3tkWIK0tiHJYn1s4+oepng6hxsaE5RcVwaIeMBiWEF7ShKRcbbFF/RVAy0
e9Sxl0PV1SVzvrA0XB7t4tSbOUb5dk9y97AlFKe2FsJMdLIVeIkcjWz9Du/+
K1jQab9YQGYOVkViEi5hlgbIPgL/Rv6VcJe/okKBOyTFggeCNlIdJ/gQ0LgR
xGsmpBc94cRRZTPem13YKpNYT4j6j/e8FOMF5xss3N2JmMeXQAsWqlQrc8y8
oNLsM05Wyeh5r+yGv327OeQJqCkMxfW5FNUUs+JnGY4mM+q34SDK3itR622E
k6NaroZKz8rLFmiyr8i63qdgpR1IZdtDwudPZb7qW4cfxMNhFLVMIU4r8BEW
AaoQZ2OqMYeitUd8C5fEI2ASa+hzHR5i8HLMfPyzf6DzncPOnuUrZUhixaIH
EJuD/GHzpo/brnKrBXl6M/sMpz3i3A+bkJmKx/LPdBex3BNZZBOI7Q9o6Bz0
09/XQH98G9xiQ56YtvGC6/Rky7mfe0M6HcOK6uZKB6CBH8NxF+yxJ10F66fj
RFI8IVAAdG62rlb5QTBUv5f0saSMp3qt6Pi6zeyF6jlMEl46Bs051qpF9J+M
anIIUDHvf7nrsbYKJoPWPpz3HrGS2BCJN8hhMcW34r4B9Gw0wgW6m9cXDlUC
K5qFoEk6FyPcL/gwvdFrEs/cjZaKJR57/CxqtbAjteoYPTsCK5OO6dbWB7jx
nk4KK4ylpJ15QMHGuzqyaVQxXZzHZrDf5JOSC7f1YMJOc4bb9YtCMn7T7VZf
6/ZaMT51BvjaH8watO9kVkqnkUB4ByXBdxn3Me0/rLDt8DHKUFmsWRKUh5xf
wj3v8J2FbPJya8TRWlDxjXHbALXID72R1l4xgl5QHQDMk6Jv5Ivk2SE7kfJo
aQ6y4idl4Z7e96O+QDvxEM1mwXSTe+2gkIBqgMnxHhMjGfcRhZN7Piw5tXU9
ejWBneMH7wdlLJs42ea6+Gk4nCDWhOjmAMFbJKUkQOA/Ns5deiWGXjgvTnah
gBjL4efWaUknHMCCXTeuiZNxZHmVXE49vA7hMAwqN9j5CCfT5woMrl7gok1W
7shoDc7yEgXsN1FpnHZAvI/aZL4KaEdSpas1FERkwgTveFmoWG0XLk2TOAr+
EN+ruFuYGfPeL60ND2RCYR4v10yX/Sc/aq8aKppe7YH0m/QcNUZCYjSCJQ9K
10qLU1S1FegSz3Zf8D48+pUxzebMo0ojk3svSIc0NQsGSjAByoaxVUTjvrHk
k8X74VuIRyGeFBVaz5dDRuqkppZlQELs081BP1e2vOZn+19NBX26FkOQiw0V
9BQT9ji8SyTQYMqFOgwT4bDF0D4POGQRNuttaNCZtZ63/LVkxXFZw1Cbg/3O
4W1CbruPLnfovryr+xLhKvqC0IrKo/4RcavRd2TE5ckIBGL4mv+XfAI/43zk
5JTHoxIOU+V9LK1w7payhiiWQYoCalyDz4issrDl1K6Cdxs0vlKlhCAJx7EY
t1TZdKdbfoQWSRxZtfCLuFVM4I9UEABXLucmYZ8+Fm5oYM5YsIYos+VgqjMB
eqBOnTzzfsTScTlLsYAWRG1CUFuas0HBqqtjijZCrQkDIgy9TSD6ZKNWSCvU
Z8Ueu6nmx3+Dp8CDCQHbpmdzrjpYDzSA4nct9P8oZ36Ky4lLaxjzXkLvjHEn
0ZDSkPuAXjT/K6AYWlsPWu5WNHJ+8HNm0UmzDhDcB8Nq/4z5o0LvD2D4Hek0
zS6zzO5zkwgrsh0Sf93ljcccJN9pz2ZgGoKEnRlbX59BPot8vug+yiLOz5tC
YBjrpzHkltp+NJ2KE+I4Xj43sczyZx4B0nURSUOlX2WTJl+DD0GPvSgMazVf
T7VdMgz9j9hE+pqRkRrP8zNISY8g2J+aUGUBH1n8Tcn7UddMw2wf2NgmONb1
0O+hfYodvShRkroXJayR0HazIHtOzI0gkxpV0C1NpbTCu7N/VHLOe2vCvGjG
xolkTmmoFr/HpZGjzjp70bi4Lcw0CP9CgZiKgz1Wc9hWN7TgeBNAWy2/mJOa
xnoQPv5fE8jk5IfcvDQJfPNs85Wag0runC2XHAxacp8pWDJWJ8OPiYifCHw+
O03ggYg7gusz0oLfVpgBzvhf9rzMHNHre9ilk/GWntZA5e3uPOKIPzrS61u5
9jtwtk8mdeOptWdZhu4/sXE/z/zE0yq6/UwOk/xvpwSnOxRW3YfHJWHm6vZN
v8ShyagB8qQEXJ3xE88Rt+XnXNr2gc7UyXBk+ecu49cpgRqINuzBqw+a1gFs
TVsXLFc0hUAhK2dnKRFYISeHS9z19zsq+hS0SvnQ12gi2khJDGr8Y8jU0PXl
IUJZJKViknWs3DlI+wvEHIsv4L7Z4fgFb1zdK6r6FmFsH4cE4h0kXbF4i+cw
aOQ0N0nLTMFV2Qw/LEhuX0uckh9CwXGBa4bydFlRQdpDUYmEaoPCTeRQV4Ho
zPxwVbo0Y58Iu6c64Mlg73iNj+2E9KlpVvh0Zw721JW0jqLcNFgab7aUiDol
LktEz8kYaRMxnZZYy2qLgX9jcq0ij9njDYAxsPEorDyi38GQ4DiokKz1qD3t
/bKgvPvV3hm75szSSpks11Qg4cSKN5klHU1Ku+6XItD+ktG3T6hglWchzklK
7Y4ar21MK1PRdUYGGyjCSLgdnXaHmhpgdpOQH0SuEVxySxtmjut+4fPEe/V/
nav1iJ5q+jhBCkBd0vt8xQoDXDJqUTHHNffPjm1Hb3USqIwErUbFHcY6ofEE
4G/YwRS4m/Tf5RYuak8xYo0YPjQkRBrjEpHtjooeFdB53ePJo8cS4IDmOR4y
dPO8uBTZ6y3dTpzBB6wkUlx2MPMPakj4xKemEuH4DB38wQjfaoXQKBWUuzFy
NfZqKmiA2RYT16MpRyhpwMf1r5e8MHnzlzKrqM950CGcC4zcuQLEfdKArMOD
aCY8kMJwIrlomjRVA6/+/xtV5VkdCFtyO6l18qoB8dXTONiyS9GLWl9/d5Jj
KPrbzhNV8i9w/8D290YrlnXM4kwm2J5383HrLZLFh/I5Q8WyBV7/J8/gFvDw
pv8268WlSipnidIb4cTtWADXm1NysQHfz9eE4eyKc1oJHOFkp562iC6RHKxG
jElngz07tNH8MVGfDmcaCL7ta+RUFBXMbovDyjucobNU/SeOM5Ps6fRhzdeN
fkYCL6+K/S/hAJXwyVRZPAVbUBvUXxeHXYLOourmaaMN+GvyT/izo9EFgI3Z
WdobhyWjlx5ELliOZoi4sBE48AJRAhzVNb7x4Z2LvVnJUTZrBwiw9MLXak0g
2vMmJNI6QaXDBj+tGTYrGFs8+P4fyUHuTXHHuDEAl8VUzsgvNcMYC8OAD4F6
BY+H8n8pEvW0DIXfuSHZP3Tusj9eUwtRzXbWqh0nKdtzv/rhrK0p56ASSLuw
0UYPIS2QJsxHw3ijaQXv0pTjaWBsiGpCElW+NBLKcrqazYnzAbqBJA2vCH5B
AcS/+8gr4E77szkCyzVC8nNAztq6ks5pAIezHz21+UWYdveMJPIwNIWqfZPJ
XDi/tOJ/ASkJkF7sVdimqGgo+gh65Raxb+f/WgPBs/j5A33VZ4d5zhJM46bV
sRhouNsmoaEOqz+Mz1Kk+uPz+liaCRRgXYxMcd97SMXtWxvVO4YyrxFq3VLS
kaiex+5LUOohHne9AhexQeHmiGgDBBOtd+5neRxzkbu0J+qmuHvPNlA/aR1U
oM2AnQrCi+f1GP1GER0H4f+oL99I1o8srNA3KQPutsmxjB6T1acln50+0uVo
A9bh6UnKOusFxs439MW0uHndpU1dfq64HmN2NbLWOFAMtbs4FWT1PjDwfwu2
Tjc7qayG4KbPtLvdNNWhBqkLUNJk2ipLa3AFa5OCCXuZAub/7mkRmj6MLl2Y
ZtiklJbowi/xHTx2jHR5ol9wPupMYT+TuWEIxhGe9qIht7qaVs3m1s5ZSE/k
HW7Kp2J2Xjnkrs10zX8yIODNOnXOW0XSXlThetEoPKDAlf5qNGcucB78bUZ0
pre+faEn7tNVE12gtv5QP/DVcXLPjLf4G5hiOzqUWGTffeC55MMnC9XQS3wE
8k03+lVMIod7Cvp6xhpej9xXPsyNTOot64QkoBOUl1Y6CxJSyS8YyMxCw8cD
PT0HcFkqyAQU97aX3bhAf2hoYO0PRgD/WaKbaSJHxGFIA1no7QfZYiY3MgNm
q7I9llE/hphSI0EIPwz/0XiTlvCd7SLLwa8rKWrkg7ro4yesI+vbAKu0z+Uj
bOY61L13C+IYXUYVqXOkTk7FUFNhs5hLIBHEAWTgOVkayye+JOBGuv4rE1G6
kYXEWQWgb2mZ2tmHgbVSTx062FCG/AKeI+07k8VuP2ZjxfkMrXlse3WNJUa5
nEXWb5/Re4/ZPfVSOaQDCwXIH/wMhNPitmRMLjY/0hUUrc1J+L8TExghWizq
RHh3+0FD5Wd+XmTLyIFmCZNX1ip7/e08wX63HvVKuxGGT0o6gm1hCGAeuUNu
ZQOAVRBDhoxfYY34lNGInBvckoJmJ1GJbW/dIH1ptbvztR2iJ7MCHye9XT4A
QrlrBkrF4Nh8fkk3nDHL8ll55X053aZ2fOI4DmdsIeaKVAu92UWEaw68ZnJb
SW9+4oQmGpfx/yfCTNMQCvvWky8qYW7FPWIpyNQVfD9AVqdjbE0fIyjdge1/
Sz5Dw388zY+jcKES92sUPD22pnBJjttaC0SjSzA0qImZJVP00/yUN1iYvuo0
EIEWMKKkp8uXduSOtc4L3VgmrJ6lgS9vc8fKQwvMfpJkLH82JL6bhvYWhqss
NKjQws2qIClGp6Jkt1ENd89FQJ8EVsfQzfOz1mFCActPPi6ZhoICTT7LyRnu
7jGVi4Onplk6gFeJlLVjdjXLqbtEZxG0VPSOQJWeUBu4LIQHJbFbz9v5saI4
01q2oaSV51ALYU6HpgOVmhboHakAzwwwKlu2/5HKuDAXJ4C3YqHOrJGzvKf/
CHii/wLcIoSghkt0JGnFXzl+y62VbNhn9Yujh5Q74QuQ6IM+xMvvBqIfLTdn
XbTstvvzejtIjBtoq6jIxwmZjIvBI+f+BNcOAKYpaKgAjmQ8Gwuj8pjywq6y
tNLuJLZ6tYZNDg0XVEBEpysNeX5x+dKVt91obtQmn92Lagf2iHznrY3yR5/B
+CeZCbuB1B+l+lVdiC4yR+U4wmN0m4hQlaoCH33EWzC72jxVw5Woed5+uu8+
PT0M1fL5cip0a9H1b3Tdahz8wA/IzY8+8nHyNjoi/HKCYNDFY3Wi0nG83F5M
6f+VFgH8uMi81wGJm68gIbkfKrJzi5TjzcbJCy4wx+uav8CuDDrv7UQiugj4
BX+w00SL+Zkn0Cd7vFaxQXH+gwn4krzMa6+K1KzcRgf14M6qEfRPb9ZX8Wxa
yuHCVTClJzX5YFpcNEl45LOsduPcde4ldm9agzgzFvMjQLu9RdAaMTWjf86C
4QaIHCybZDGeU6y4I2zLWukivvUHbxYskHRYEd4dMEPzq8RyRS3RD1H7xM69
f51HtvLTtV6gbpuDju4/+XHPy5l/Nn4RCPl1RTLFVHXonsC7mNBeL4H3wRcy
7kP9WHHhTqesg4vfRG49VbWIDoup8iGxdnJo30QGv8jRM/CW8TAEzAQrpgDm
jQJ2yp7B7eLv0mbrvWLWZ+LzRissfav6YF6vMe1uTCXTi43pHvYGsLYvPZ1n
B8nbPZiMVQ4snOMH06oOe4ualncDSo9OaV+HWIOZ2ciOnz8bdBA+ZeG1S3HY
VSmt8cfOo/CoBQDMUDYFWLFyswVljL6vnRNxXBofwELVZOyIQ6K62eUbCOXB
47O+IZ+an6E/tG4gNenJ/QdWAdVu3KB/4FKS8C7f1msHICssDd6WhIYiSqUF
h3BQlhk//v1/HwRokaIV06eiuuxcgRs6EiL5HaqdzkKqM4cDThAFFWLRdcPv
4bKefpH+xnqtyr+av2QGiVZtVWBg2YPExaAGy8Q951jcAtIrg2FboyAc79Y7
HwCVmUzRB76/2OEYTPq3VOyiDhIj+8uZRGr6VAPJ7X1gejRn3COrSGqU+GMU
au9PEEFKXd2i81df8JJtvI5hzvOul0oKfJmrSdy5jyhaTi7Eq4B7PK2Lbprs
2o+dUHTQ8M5CCuM1kcHE5LqTUGTjEtjUyQl8UiB8zcXYYkalrTUCpFRSwqKR
kgNjVYMdICplw31/08hKr51+hMwQ1ULZZLiEOpk1m9Ulueo9dEhA7Zd8vI+h
KGb8UbZBY/IwBrIu06nZgk4TpTNz4Chha84tEMnPyH5Q0tJe3Qaeg6lPpBzM
eXpbnkpDRxMN+z9QacFgKObCCHnNTuHIAQbILP+8tGaU8IT+XIID8KBhu68l
OxoL+apVovj7toF4dqSsw0Kay98iXbbfKDXiIlnVabHWL5utnOuzRKulaZ8G
v9XNtzT+1gxvf4Js9JfE1TOD7jFz7fKn8n2FXbz3sBniIfHOPm4DbCwXsmTo
591vkhfbSZ5u9V6r+FCSMTLCRkrM4VjCaL0wxb+47cfy4/jb514CtBK5oe2F
rm5aAgiGYGZn1kkgaifOnmyixS5tqd5TqaToPKsnqjCOBBiRtfFvMD8C3sNS
kYnNxrCWLzvrdWe5D3dP4bO1Nuw1y3sGfoBMFVPsnfgdbv17FdfMHswU4HsV
HfYibM6K0TyhId+8wdIyRIGJyNVqgLHUw0ViiF/U3UQq1t31zyPty350iXsz
LFd1+i1I9jPaUa2oHRkdcW/f/dpok6M1VQY/WR3MTeiJ5xmPUuvk9EIAMKRK
L26z8CVRMgCYWO2zBEhnW9Qfe1v1VrlkTTrbIJovOPOAo7r/OTjaW5aGaxxN
5IZofGiUp+IqcGE6dcK7k5wyuwr+ldCupaw54kW630AUX3h4RRqvs7zfrd+4
m3CC6C+cozKXfpIp4aIvx6s6OGl3GF0TIYe5f3NMURZqAeSKOhWwSZKbeyTb
VDRwYM69yKdH+wGQY0+i8a0xE987fOqrcZMMakNFDLUqBE06V3gtIMUlp4FQ
L9SzeVr9CmvjErcijbuAFRsh0Cf4F8UP4ViGizEYJheVCywmIer5GrNGaCUg
wzKetcc/JH2nHxDoxzpEXSN9hG/dcWqJROGk4jNC/J/29DIDsJxdpvPpk9am
fNwz7MR1XAnS7nnaWcZpo6IrHWPeSxTN5rostEwH4gmoNmoo1d/aLYvZTGIj
nctZFs0uR5UBGipm1Ql+6OvMF1w6OXqY6sqrCsnG+iGnYNOQMH/ph17TfAgL
wNpTncZuOyplmmwRiLD7k7DVefthHv+F/B1myY+55flGlL++UiEyEzh3D4xK
qa6RGeceXxmwdjhrgTiKOVJPyNM5FtaIvwtezbhHH8Uq8HpjFudBpDGMeI1y
08qx/QY1MrKSW4Own4VslyIZ83nTsuf2g9pYL4yeiC/q43ps8TgGAJ6xJvkG
9yPnSXE4iYxwj8BoCHSBvi0zhddK/1X4Ih9H2OJKXMy19Dyq6QqFcy3Uix/y
DKGChUFaD0F8VnZEsj9b90jA8NQBKD4FoWkHLkse7CcSs2MrAcNNr4PVRW6p
ZpnvRmimTmmmlrY6W03BKc4qt86w0uZf5XVN+TEuoddFCY8Xr69FZzU5UIb0
874X4xBo/BonaTDfLSkL8LS+S6NHLOele1Y4fhfDrizkKw+XAIGDDilX4jR1
uEHzJhIx60rbJEm0iNSkowoRRL6d2QC+ty26bG3sDYboA+aJgRlaWaXklkoy
RiiY+uFs+nqefe2e1RXLszhyBPof1wiIQp6xlKEyPgTnd9qLk41eQwZ83k85
JHEc0OpZk1smN7h7X6k+PoTim96NXxWgHnXtlrYvfyCriTe+S6XLSycj/ppJ
CBTCXV4jJXQrAJX7KGUFAxIDxcaN2O9sRY+x7lJk8RGC0Z/P1utot/L65JAH
3q8LLOQMdPfhY+ahxSkuZcASw+CcxMjbZ1SGutt+ISNFvpBt1Wup5zGXn09z
bBOheCxXrJ+FWeg/pwOc4rNF95i1Z7ESQX2SlCH8GUn+popET6Jeq4BV9nkX
6AGm0F1FXlWI8cddCK2ufpMJNOywolcSOBynTinl95XcerCMEbQltL2XnjX3
TaUPG5HbfT/f00DOyPqJ15JEJ3FCMJbVt3b9jQnbXC/X06x/4oL4I6ZlCxOA
pT/NsnNHHPC7xQzRN2YeRwZE4uh2Q80V592BC/V9Q6/2tonWwg1Hp/RlBy2k
SfLx1ij3zsCD9sHWK/D0Js2NcaUQHc5BI6yWnk/sUXg09UprqT30uMqVxdpg
7akgGScDhQ+JiOEFxUcbsi44N6WaNBx2ySuivN6WQpTjitfuqSSGQUR3XiF1
+HVxlHCrSJWhEX9N1HEhLqNLSCN4E5QsQbXVBxZw7vvMxyMzSsSeYbP3QgsC
IlTjn3zvBfMOITsrtPaJOR7KRL9mOyMGxBpIBxM5RgGaY2aeWV7BZquwkGp9
wo7VFXULwhJGyYjv8SrhD5gk2aAFy2AE2xzfyDGrA/IzO1MuvJAk1dylYhfE
T2hVfO0FFIkUQu5gYO4im4JnRqxz0VxbW1MEFUT4ySuA2FqUlxiJnVSMiiB5
TitJp6oNVxFC1fMcN5wHaSe1tPvNSCU7ufgldsurIhcIrP8m3jBUTqnXQ5YE
fYQSjW4bX8yH/StDbKjviK/y4SSwjQZYTw3IuaP5hYE6sZ49tRzk0R/lGeF6
ps409D9M/ejOXj1FztE7bBcFRumjvSHxtZP0hS7Vc7IpAMcWxogmcqhWEIJw
X7jSvecNBwF8fSBzz/b+LtbYnMy/btqvQroEyUbd//RgP0UPhq/hFkphmR7N
EWxvxOYziBmnOeUpjhyhALvw8PyqE0R+6KeaHfGxwcW9YxOxfM94aMXo73T3
bIf6+0mobzFM+6LA3qTPymXTFl29TzatUEc7J4ivT9iaqElraBimcwZa+m05
8/r/5k3DkFIRWfpR0lApcFSjh0k3ebwr6tQ93auCmj90fkL0f2wHNRzgjrx1
EyF92UmvT0OQP+j6NPBQytqGSfC/r/jNrA3z0VE5I0MaHvH8EkbA/0HC+rhE
Q1zMIrESj/mVfsliLt5iQhdouA/rKkI9aH86451Z88Zrm/EnpoAKewqZ7sF+
i8wAK9K+FWevFnLes4GI/Qvc3hBynM8QmgAKwoesITFuNpm/TAAD2d3zLnL1
9fwMGQsY34UAzL9DY9hU3WIMgknqMbs+hcinNTgR1Ama1efD00W/AJfc8ZND
ZrHbtcEGSsV/7EF87v5OST8fHvqPegRytljyKHmuSQFxR+p8WGdDXtSlO8FD
13yEaK+Rf1XYUcoMeSN5i7OIAw17wRbrIdYnYtsTjjXmv+/cTHfuknS+uDIQ
h0SM2q9oymM1TRkLxJ5GMLwV8ro+/USHE6w8cyUZj1IATDdrefDV8IV/UHO2
KgbktAiil3en8W5s+cLN4uH5+/Hv1tdkzBf2gW1/sH9RZw6WKG8jZUGUTOpE
HOsXjUygBk7BNgtLg1iJGwZxcvWjSFFw3c0uMm2R+sQAWRqpJN8+aNZMkHK+
7v/fTgdIoozMg0bCJtyxt1gpMFjRvQBwccqFy3NqrGXVz1wLnWgofQeTN52l
OdHrCYZ1Ug5ezQAxjMULjO0vlhr35HSBL3QRXKhO5csDz5NIZ4EwPBPDJAXD
bdTJlaaYALCMWRFHDIJUySA8iAjXDTz3hfSvxr6ex0gaH19vfcQR9lOtLyUh
vLjzUknbcilK+viGtJdi8RHA/f+57oLCEaiEIRhYrH2Ejh4GUkSvuxB0g8MR
Ld0a+xS3jh4eLxgSM1I/ufHNCQ3zxA68Q6bJhfI6xNLdqie+h+2XajQaAMSP
Pg2UCKHOOhhgrT3vU6ZpyLBEmNCE/2wZOZ5ppcGoKWgaMpH78X+h2L+aFdZc
zrfYwDAiSGRbsSBZ6asslsY6gDY2pkifN7c4w9ySjZEt43OD/XSYm1j8Xsvt
YHHaL8fcvy+gYNv787RnUYoPhAiVT1mx03yAmN01t46teehckglVW/3PdbJu
wmpb1PXeiMUi/OSWcSnXXAc7DdM7az7O+aeHlLPB3EITZtyzWQZXziwcdKRu
l1jjfRSmAlWk0Z3hQoiYoLto5bbqt9aPnBu4fDiUBxbehE3UEVhfy4FKka/H
7lhg7obfmElxXqyYSgquMkcNTDC4ZBhUhwUfIL0r8ZZmSM99OihU7P5frFw5
hqgyQUzIOM20mvUtNQa9WzpwZRsgd1T9PHMtNOLUGh0lVvP0fncO3Xo400Kb
GEtxRMXkJhApSQV/ovIqxS8T1GLxsQkN2yAU86BGsCYz4SwGnbDcE5OB0WJP
ldGsf9IeSmN+tg0beFDEj+qsEkPj/eOVozm/jjCXah5H5eHh6gs1IIJqCzPw
jBMowhYJcz7aQ0U/VNqgFmMdDan+p6VDJYaOqYn2RarTLuibWhDkDDLnAg1h
1pybk8b2R6c8lk9ZOOnAqH6Edsxfc/HlirNqFGEKMk6L8tkrRSRidcCi0rQ/
SETi57MqFjttypH0y7kYNujPh22RivadCG7uc71S7vH3GmYkBUqdy3XXrQnS
vgSc9/r/OUvYNTOmIjRj/C3uRhkJLf12ri9I1cE2sQj71N3f3DTYGrHZXHGH
+5JYMONKj7WpZHgdFpnBIKzL0h/rwbW+Qni1pRuKe0hUPZPBHGHRe8Nw55ry
laGfbZziXKAUTu6wBwaa5bpee5zfezEqy3fqk7JgINeNE8hhS718zV1rGZGE
YoIPcFoJy7Oi6piGuQtR7kQt0zK1HUXmWAlwvbiYKljtxkCUPboUVdSnvcFY
MBKXXlIlr6VJV9B9SNkMNuzdjQ7h9Xyzl6O8EnE6Z6oNa9MV4DbBgEUfvCNC
53IUx2pCGgVtqMbXeA8VKNg28wDEAcZLeI8/gKOrM4+ggnP4XNzpL7ku7fnB
xfu+iZhuvCOasStZj9e+uXokV3E2N7DtQ99HBtqCsHiiRkJGOn5ZFkthyIT1
H9uTb2VO0RQd1FiZiF4e0P40EaiXrM2D/QDSAU5mV1V1FUOY5qdqK06TC35/
3OFdEm3b1esWqMbMKWWUHsVZjNxWiCw7N1UuJZW1IisIbWnH/jIU/LwhhI7Y
7CrHimyJy/ogFEwrn9KQi0yHgIFhqfEShZzn1GrI/plufJZN8S5nLU07dznP
uu/1tABijzCv9FJT9/hpFjHBST7kM+cvsFAol6p9itXcfCulb8xwh/z9qLfU
ADos2D2lHOFlQyxwSJlvtNhgO/58y88kPYApzXlWJ1oPq8S4Cumfb7WaVgl8
NgpL4qD6HheIW8Xd6SP/f2NCN6eoTY83/Q7+ucMCUyq9Oz3bHpZZ19KwDKbi
p1zKEj65KIiIY5JyknEcCRWLRILLcisBvOfLt9/4GAlzYiP4mVI158D4y79F
KI8i4Hzo7Z/JVlBeX3xMU585orNlDC61uK6PiGG4AcMnUVhX+gzVkqntlWo/
B6NnYopyPSx4Xs5JRhwxYsuOOtqEJbaR+gWUA/W8fFALgokjN80qUCrhGaUl
Mpb4soZ6pc+i/+8Z67I3nACqikMYKEd8rZPp46Fo6ucyykvqRfOIW26CpFV5
LP3IGSd1TR0ZbQ2gYWEVRZsK6xPfqWyfXqITcrO1OH6GkGSBh4fSZMZ3253y
AVEmk1+kEQ5lO2syJLjSz6GhmQpSAskEIft33JMOs9lnXl6H6ClC5jhIjVpi
nkAUGVvvT5fq3kwi/Tkk0ak9nxOGQZIzuWoc8Ds0REkT+chQkdwC6lKAUSiB
NKTw67PrgKEmrsX6BGcBoP4FL1ftEKnAFjPEwM/+DRQIOwPRUknyzuC3i2x9
x4cQiBL4JGFOYO8xGMfhPbDB3MxmPuWmpZ9kO27/StnMSTW0wae+Xgaf4hNe
b8Me/J1XwY/Yei6rIx7Z5iEtpbTIDIYHw1S7MN1D7LXVT85UdXpKe6SCbNGa
0rD+eVcrR/Vc19FeAYV5bqfWXxfRqNCMByJ+5zPWzo0t08UaoZOijwIwmdTk
cibbX0MmK4rnEyXVEJVU2YPKl122jgsCKNaqmtpNtcczXHs42Kn9hoKbQ1y1
Fq+jt0Np9lmkzILowocZim6zQfgAhOiz19B4bH9H9+obKyTOCEL5k411c9In
GJrT7s4NcPNUJm1JX6mT80KDRuRDCZAx6cun89tAKuzVMA8fhcuEvZW3V2Uz
EOuwkPe0/xraRd0fKpr3FzIcv0x6NAeWWfauuWQ7oqr9CeB9PwlKM/BqW2w6
lefysjDhfGjQg+rLZuB0jdx76Q8bloR+WRhVaJ9NMJQ79iWlcyyXim13VoR0
Mc5c8pIzm9oqJdGmdpFbaoR9CdCTJZV/chKlHjEL1shXAwKQmmxGPOG1rq06
PXnva3Ytiq1/SvicKrmi7kPRtIPD1BxMFz8k9B20dJSl0g0H1r4/8iHT+1Da
/QuXi7R2uJNnfdWSv5REYQST2OjDo67zyfX0HnzUOPdvah0ctZk+Ki0AIWx9
PQiXZGn42ym4WFCaz4zX70txDKOvjp9hSafj4BVz5pDPtJcI+heDW4A675+O
CGbHV+jKPN4rN1o/2XM5d+Xlcfq+WVXbsrt55aRuWeTA+5Zga+TLnupkS73S
baT7Q3LKEhJBfr74VdRIoyuPg6xJ3dwFDXhSLMLn8qLZ7L8q0AW+2s61vkHf
ucvQnfKDz+ufPaNLXux+zywqcSiA04b2GznQdWRiy4C0+o4TO1HxeyoO7nQx
vc3SshRgEm0mRwA80O9tUJe6uDPpV4YEgjPFvcMI6Y2eEWWTH2qdvSkmG0p9
jwtUJuQ1NUos6+x6YHcImdV05n8GKPqlxzasoBVPuHC6A6D/kOr7qcP7u1GZ
9X5XwMfIx9TRvVXPoyDxgEqzF3sjQmm1JQO0YMGyE42aSNfNJTA4XuAVcLMx
NMBU6+fj83Y+G2EYLfS2nbWmDsLdoeCyRFW4ufZe3/BknZ1ru4dncqbBGXqh
YCb59Vm4CjNti5k03M+VwCy/OXYOptimctBgBfKTRCGUJo4PDtRcaQnzHI+X
QAZj2madwyjgrEKp5ck50Use6YFtZJKRctnCWiGSqzGwQIpohPQezH7EYl7h
mvgAXPBk1qrbM6/hWdEqLOZyVwgxl2VMPlCBXJfGBOKs/yPiLzCIPJsfMb9M
S0aRa3m5mVvJtw58HfEoqbw7UtMWIWJx/F64Y5plYwlk2bYboDl7/domEeIb
SLff/Qf223zFkoey/c0bLWnY67dko2ei21GsAL8BPWHqQ+iXR/7cbftg03DK
tamlv+NKE3NSr6drJdYjcp4dOYOejBUzICUrXZ3zT/z/Jm47WzZfe/J43Sey
pW2TSs62OYWOmF8AZfhjta+DzrH3bD9aiX3cpO6TiCPBz2RDrfKpO7nW4CMH
ZiD9OHE0rT17fhq4T7TlKYTFAbzlWAg/96c9/JHyvgdTr4CqsMWS2tlRdAsU
9Ri78OCRNO2NLjslAswNcJZtzbZFhJn1LN1OVsdl0KwQUwg06uEdqmY/hmFL
EJA/iuZgV5LoFA9j8MAmdBKbAkebhJVvkGk1J+2EAbXZfXb5OB5oq40cCOcb
dJsA4bWUvsT30VXmcxhaevXW2cSeYBGsmtwlnSvFCFW6Q4w8khYcjLLDYoy+
tfdiBT0qmzRn95IcA89EXXKNGYjNUCCGSSgAsp5u74sFFTLADa6U2/25vDzB
+ZswAoJYCaHJPd/FvDfkorCc5b33wKQNs9o7ztUG0C2HwduyETeITQyI2R4Q
WTsFV9Gk3quxRA2+ER6i1tgqdc+d6SsnVGtKW1E+wymW2oOwpN6God7yHWXF
FeNrcZWxfkXxzGO6G+fmsmafK+Od28UelwcHrYJn1vHUG6lIMCY8M6yqKbw6
DdiG+Xv8k/54KYCyrKbB083MEwn/AZMrKYQeU5FyeMh+Sk3w3ciwAq5nLKbj
QovszFV0eUR5wwU2KyhLkQz+dgdT6Ccvp0OdTqGp1KfNBoGw8yNK6WG0jMl4
5RuwIJ9+7LHaPzr/lDVfAFQYAVZQ820rFnFx/GAKea8Fz4komJbBx6jvpHPz
9EVVQxDUwKSjFyMkXyMCc6q122ltHby+et87b1/NPqALSTowBMMXOMZ4A2tU
HEeMHxzTX1m2QDoodwZCqq7ACXw+1GYQuKuOg7yr8m/8Hi9qqnTS15BXHQCy
kgaJOHtwh4F5hCnlgEcquH2fqKldEIEfPv2GNm3Ig0QggZQTZ/CEpzJQii7n
Jux1HMb/pOED4lN9UQLfNRtEW/zoL3j6SrrdUxP8YrsOY+PkSH2A7H1yxMY6
RqFq7F/uEg0vOqJf7tX6awwTTOxjVFrN4iNaA12goNPpbPfze2wxV3WngisR
eyBG31CqoZTigdoQ9VTBa2nBJb5AEO4S2ieQPNL1mm7r1w1Rsvalb38KS3bL
SrONGkG1TYO7i5ccdKpn75VKU6qNmZnAonWo9C3cFr3uiZA9t/7zG9EVDd3s
vdFj/9sib+HPQWI0A3riqncIRxWIuwBQe+aS3Egnx+lbKxgq+C4uudvflyAl
CeRRZS7UOk8tgZnmguKmzfJyr4EKk5ViG062oWWdiSF0TGa6ldcAB/l05Wm9
dDPlHy9c7C9iwsL1sEUphJhYntmlNHfUfSvIp7doyrYIbOHGB/hjDBqzVhLW
DsntXr0Vf1JQH+VMpDHYmwfcy7SdltG3nyDvGeS5VJpZiYGz3msaCC6fIyQ7
qFACU/oLopYT2G5jd2GQbgoatauNHQPjPL3ragHx0GdKdXzZx1/3t/MPQ0nr
uH1Sc0osrrjMFunZLrbAg/mrGhd4EuGiDoY5JUwozK00OWKLnfMgR9VNbk9t
Q2NMUEa+LnQPJgR9Grq8DDr0cXmLrF6KEcwRuCgBiwPYkHnRClqXKe+5Ai/B
vUbu2DJrV/jYwnIodoM+0HupUwUPcusuZXhyTDibgNelDVM9O9exbf+MUWO9
pbuoHjZ6FRsagnYzD1pEVRmIXjbyWg8wqOj9OBI4oo3Sj8iSrWsucJlrHkcc
9F9elsu3tHgRy6+uOb239CCOjCTvmPb/JGjh4+Kh7okVlgh0Ds39ntiYbOmC
nh+EGnbmV5tFgszMbFCIi8Tbu0klfacXyG1IpXXvcmPRTh8sLyRurgbF5+XD
DpL+3GZjzQkRlp22b8QxrlL8itJh0/aUB1VcRBOZSn6KqDWaCCGk0Zutkk2J
3rXR5Eb9Tffh0gxZcVNQM4uSLz6oWcRF2rrZCvj5J7wFz7ucT+XqluqHN8fN
J7lIFY+Ugb136sgRsseQ0tTLCKHcTfNl/ER9xj52APMgYzxDucdtSUIoycmT
/5qUQLwbXwMJh09cFsIl1302UhTJ6+p0rtk7uUSPbx2A9cvMFMu7ZDka7Mdq
AkJY7aBIqOGYumgJyco++btryiKGm+QMqNIgl9RXr8zu+JkijSutCgB254qN
VTJT90TeJgAxz2Shp8QWMG3N+o/7FUxTF6veKWBoYpMTNpbFzmCMBdkjKeKl
CzbTrQ1Kzc+XoPtsJnaBN9PCy/Azj0hEv82PAaadmZkHyAlbH1e+RPC8F8xk
h5kpYcV8reOuxxpxrGVBLvIdmtUsHkFgsKJ/+q/duBbnlue5Z63kJ2tgh9jD
Pdak5BuqyPzzcoLSE9bbtHgS99J3euodxzXyxBWyhEMhAJTCM3V+XDGi8LTz
6lyEMEFXNDrVZ22kJFgreIfj80GSCv3Ae9zg4lrmQmBL4N+ZQI0VdsfJAV8e
swrEzjySJy3172JLQmyGlf4SX9tRBU+nfYGOZhvOXORgmpcDcr+xiZdTmRUD
qt73gzhqtElUY+XJzzuOOZYGA3SwwtSUnR5m3Zz1buSB+r5GtEX06ihrFaGB
XKyUjQPgx5+MSn8wYC4XzFg1xZV8KLeKsdpgJyyuuhV3unD5wzXMPodtZVk/
qLflg204joZ7y5NwE58vbuKbQp5D8IdC4psyVkQCoENv8qCpv0odkZw6RsPx
VqABefSWfKwwEq9QQn/rb8m9GiBiB40TIvj7sWOIIpvOTTx9MEc5Hm6g3rXv
rPwkQO5+UjZeMct9LaykX2an/lI8XzI+oQ/9kLvAcFDHhH4ZWZM1sSt97Lf0
jZnNGPvAZiKeuN+gS8K0yjt3HvrnYqA/EvodCYZG8ZcqPapXODaRqICSS66K
KgqFvol8H8O6MygRntZVWUVxSOWuOm1G8TWCl6Tll+MIdYZ95fXVHqibXmXs
lm4GpIzjjUXRozy9GJUkzxfKVqhOtG+dWeEEXKZXoXUbxLMP4Q7XlP0fT0DX
tuXcHTLv4eOGskARZfMTtgN9o1NrLyanILz47LFj7tsUw2FcikddTzIygeVi
LxQo0RsEIZ5LiM6uzBC4mS5hP6/CElesrV1/Bbq41FrshXkpreXcnYLFXh7C
k/VAnj8xceSzzCuQptfoi9XpPlIW+cuxjQljOETmsF8dKwC/Bqxg3Y5MSxp4
L5qxyx69qT5HkpSwT4Cx1JNPVwk+Cl2olYzHsHRxVmKZI/fpxcgcy1oGkrvO
unYbRk1z9cEBXT1sB8G5pY77YuOORf7htx1CV/Cy0RMPYHIEoEW23WeI4/to
WSPWnZoql2kttnHQX9gCDRIDYXx+iAyTmJhMYZflCvYj3Fg/Vcdc15Lgkms8
bLww5emvr32gDRYeS79xt8UctEH59m4kOpykfl++7wqpS8xvsNuvAMp4LpUy
I2PnVHLQEsgwTO2JrMMGC88LpaKcNApB5k03iYjQ8HRXnE1T+/4cfBYjV2Eg
eKn5T7Lxtxb/DdTcQmqIsYELZ/DGbXpfloJJL02ObYKL9ZKgCgus8Trl6nRE
R6Kqwb2OMgKSTz7surWKbU4vjm01MG7R5aj+jmQxOpmLmG9QcGnvM2xghHnv
GlqhX2O4tPnmSSpyJisFkgihZpcYZcc4iwMT18OuoemNqZiJLjmsr+tqAsd+
HJoibP4o3EuFMsaL7AmujqQtwFldEwnfl3W762TIZbmueO4P7BJaf6BzafOt
AdnaltUDFzyZZ9EMxAjoCQqMJ6uKoPtZyE6ahUd2Y37kbvrTG6Ix9J9xzov/
hhRjJAdCIeo7QbGVs6jEkaY3M71HFUcj/Ov3V0sNGZZPVCGqk8933iviS4i/
rOXO2Tcx1DqAz6kIWzdf3Z1Aw9FAwNKFDjK3oxplbmrX44GtiTc7q7XsrMY8
e3uqaBory4KrbUiQizjqZO+7SqOggG100gdfb9S2u4QtAI7qFfJd8lz9Cz5X
SplC2mLWYArSCBUmBD5/jeIw7L+ExFNR+xtzknLWO3Vx5g2b2CZEJQwWGWir
QuFx3SYj+t7KFf/KcSEuC0MpjAkJA/iSl1FpGdXMxzGvlgQ2gQRITw+BeGDB
4ddJFiP+aK6WWL9QX9rTd9/hOTFSFhLQ2j8T2aQ75K2msDtECQo7RnBA1ldj
b6L+/q+TJygMJRVVV9nCqlXlQN3TtsG7LDu+XWgx/jSRsk5cjNxFl7/bAN0A
q7eSbajhpptrZbb1hMi4FnkoFABou+SpQlh8PODlxmTNoqsJvsgGkm3hfsJ8
LXzdMc/YpjqFztlRdCsKxOo53n9kHFqScyUsnzX0BNcffNcTlXXLRPip5CZc
crgZC6llnCSXKBKSFBKqgrwady9aoOxyaASuAKXz80VglXhrDbw7fNUW5sE/
X52IJdN8edddMGVoFglVVd/iHNCiia7u4o/WSbIYKx7wZoNN+uS7y0HGHrs5
C9y5Sl+8tFHfgokKbnVcI3w8K3uKUBoS0g9R0KRtNH8S5pI/juGc9InOMrmM
btNAdEV5h5ShtHaEND4Nl+S3KGj1it7pfOX1S9yNtjmKM98iJ6X64slaC8Sg
MuhCrtu7VJ0NIBnsOOpsLO+jPqmva9nY0InF7Vpmv/ftGabW4BpMUYMpsQwD
/as7vNf23LkY92KSyCgd4IP3dQYqPgMSq5KzxVRg6wbilm1xqTWK/88cOMLY
gEeVsTw68cf/lvQ7eIu3g2PjxiPtxGdhGz4X8g59fNnJ3rrigM2Jf/lmBffM
ZDlIh2EGFTBpYnWpBq5nenvLhCsMDLERDilbuzyG+qXefhsbBxeu8sSThkpi
uaAaXuYS5c6ZSVGsuwYBMEKIqfGEt5OqjmkczVsAdjrida19iPqd1i3OcFqu
PwYOHLiQVg32FPbNHAt7AjoTVx+zsO8MFCvnMhUJI4vVNhvNDV1GEmlSkHNc
Dk9fIkZMZqB0LB7Shn91pU8Rri8HA4kwgPXlWMUX1XEIGyKGgBVBBzwCdt1O
V+kgyWOqY3MuC1Wff6AUNhuc/cqdbeeScJGccXe7WV4Jwv6/vkJUaRGYR3Sd
UpzDI8iZmoZhJ4/eeKbwI/BT5U1B1Nz+Zo23YC9g3+RADPLE/zSGw8Xg/MtD
/o2H/Q3/8W6gZFBsq+0WL7R5SG06udlJcztN1N5vos035lTWx3bj0BnAvHSe
bWMEJraXUhZq1pfvSqZ+23i87AqoRF7bXfv6oeWzYS7M5TEpKoxQZG/EzLQ1
h8O4UEYyzr6a89XrwmiyjHwtRce0qmiBR77/TT75pZSnWlGIzYAUHzJDhdBL
RZdeFfMDL3ajNLfoUU7vHTnPYA0CPK78nI0GgxP1WtKfgF3rN7ppOQp1eJwq
4lvRGNCL43JE0yait3wkJxzcqSEzu/GN4zmoG8h5LTZ6mhs+Bx8HsbBATqlX
hWjXqb9pfln/u4VpKiF8jUEHVpqkt05CTma796cYeXjVODpPmxZmBocuwQC4
xvt5gfMFeokj1KqOmTA24+CJxF/+dOxY18bUDILmlXwjYZN/5p7g5fot5B6y
k/dTdttzFVDabOCsGv05VrZJJ2EYWFFUn8TLilOOLZ+R9H4nsVeleksTlcVA
TTEHnhnc1WnNvKd04U2GtLIqaYtNp9yR0nR7TVA25yWIya5X0VSArVmdsJe0
3+TTO2gqzvl/NTpxuY+EdnQo5JSw6jZtOENqdKI+6L2jvL1rSp57smsJooiq
DIOdkLCkngbvSdUhJ8hlLHJshRCY9U1i5s7a5ExI9B3DpFrpE2X6k2GYkQWf
ZFUA5El9w8M9rJXuqLMXFfp4Vrudy9sSuxV6kUCYUNGTky8EKuITni9yEnCX
wNyAa9lJdAp6uJqrMvHNNUkVmzVlQflIEZAIQxt/8w3x53XuSl7PjLz1EHfH
9dnPIh+9aNHUwz3EKLHlslljKl7Wp2E5oNn8eJk68kAoReaO6dPTmSGxfsMu
AEabctHV3eE/3babHleouJZcgTlf0w6nJh9J5N+Q3WYlOVY87QRaM4jqYQ00
2/u+/j3jRjfCC8TIDqk2mL6ueBmKAQ1HPYP9Vyk1jYOggsQw/+lBFlnrWXZB
j87ussbXTi0Y7fxxIWbzSdeh+Yaeabn3mLRR+bnIOz/8YsurwFbxAlEFbb4/
7VdyLgSx+xuRoMS9RrnuoVk8o4VRGNISVVL6H+WdQwsn6KtvckGdLRap/cjb
7mTCf1YmdZjH5XPXqZpMP321aRqiw/F2O4MDKa/PVz1q+4OpQhM+2nqLumdC
G87Zhizc8sDR6kJFy+L6r9mnlSbx4xm5NpV2n/sAG4UbmKJDdhjA1hGDzzg/
KZiX2OBvGITAaUc/0xbCrglp85fh/Y+1anODavBjvw848PxXbFCMzHakcj5+
oP/U+5Ew7f6E58fYOpeDWHJ8eIxUue+yvH4vucB3XBPGwOrBzJHxMfnIwPZ9
YTTUAbjy1mZRVWqN9cOWrMXBrMw0zPC7N0asHiAEvH0XVfTjbsVyu60bt11n
hBUAhmP80gwuW78kuiid7uGUB9Dc/yTH5pPxstgokuvMl6tE+g9GXWrihe5q
yMbzUvxQJR6TtwSHimWoV0Aep6w2KIJfqH3P1UdemVyGTFXH8w7ebWjYsl5M
pGSsNn5PJqMgI1+Ut6aFfFYxf3fLm2yT6X3JYNmPNkYJvj7I8isZKyGe4f4W
lUtVr1euKGkZ8VxCKIFnkzYBUDcE8Yh+w8aUbs1vq7gy1loTkGvUN338eX/I
E3INFHRnHBxpk+BcVVXCDe71iTJpoTe3Hy01jsSwTgZYS3LNM/rUBPOBcHDc
UIEHst1HQt03DNhTodqseV0LCmsB5XmI/MS8yfVTP+FuOTWl6TtHtdnU4LWs
Dp1BfxznpS59lVSlpwa5gy3fZ3UPGpijGmLi2amV53xiBS7Mj1mlk+gwXW/+
UpMjuPurEIfOGXpMI+o5tDX7wQt11CX7hxX4SGtGJFxFM0mQ5mZ+B9cwuDf2
rzXW6BA8+QjG3qIoU7F4/c2Q+PJzxREk46k1NiNcYGjM50EDsfbhsj/tZMTU
UGvKUsrQycthz7hkc81agFNwNDQreDULDpp/XaY74/35af2W2LQrW19ZDfCO
WjszJJ/HwFu35V3huU5joX6PWH4uVwEgTLRjz7aupVFIjnvzDfCF0wCPCy5/
xPprh8G1I0JMCCtzAV6vGIh2TqtjaGPtZ7wDPNxfXVmL9TWzM+/mDoJ3SZBW
z7J+n1rKZJqc6mvpkLDevkxC1y8kmEFBh3wHj1ER94nYr1o5Cpzu0NWhVB4b
SHU8hECuzdnKy+eiZ6t/bWOXGKL7jOv4L5l+ivUhbe0H05jYNcttXQjOjijz
mJyA+j2QGc4sYxUNSzVBi4QajYx08puGQU0Nxo30AC5W7xqSiZmtDJ2gORUY
x94aN+lFF5jwqcMkNyqE25HGboXmXL4DDx3YReEq72L6eCOb4nWC9ywxU5VN
pIfAIlrIqJ9UxgRpB2wG/bwDuAz7LIjgG48ALkfbgsmkd2fZocxdM13F0HkU
PlOW8LfTibPwIqlyYgetWMBekGPA8340RdzwW72pDOUm1yL70QCF9ZFr9Sou
LLNhpNnd1sufNqB4VLZQfZNKCvId0LJjzH/gLIipAXZQ2wjmr/JlMP8GaE+I
YsxScZPaBzCJAqaBZ5iLA6NP08dy+kNWQ7MABmAtCTlPHLY2DHU3LxdiO7Ap
KVh/UTRouWBiRvZgo8WQL6LJqc3YutmaBFc+gTuEIpJmtsf4Bl1S3+oPbrrn
61wFk9ba+YmCvccosdD+nQYBxZ1taZeAHGCVz4ksbt8Powzd6crW+0rKIdtd
HgYO1wChOvNFEuIDo83j3T/BmGcPxl7N6XEseOowuk72lATn+Jm7cMQs9H6D
ly1gHOVY+L/GINIjctoocJKUT8lqemRsk7kfgOWH/tkS+BJ1+o5uASiXnqUf
SY75m/P4FMqnDJpBWPjJawKWrmP3+UxZrsWxKJhiYYOWd7ZndMcc3faT7qbg
1OStypocdeqNIttDH2PHGSbvWr+hv2VEOp0BZnuUTaaTBz480arVo04WGAhe
HF+c1eiVtwQ0o+wNLC63wuSlEVDCPELN1qe0dciHM0+YgA9+3SvqR3TEiQPW
Fn261UvKAq3pmdOjajh50SptmWCX0Cb9orKNxsL01p2kEOjCNOJAUrxsc9LY
ODjPweaguh45WmAqMqz7SSpB21t63V2fT4gTeuiN9V+poheFUg7WnULReMKX
lGlCJRHgW/1H/4YqZvTQ6+wnzfi6DACODlDDHEtVqvinqyz/JkU4TJ24s4AD
L6hahI3mhn6/RgVQrOsmw9zAynqmmLY+hxzu9M+KBlh2S00EDbJSRViEL0WJ
gJYj6CMG39YOeNwIWHIU7mOFV+E4ixKSpoXQNqSTa7M/GHh5rL9SUcUTBsFz
Kes6D5U32oh2hPI793LUEciHf4Ru0ybnJWjzPU5raWRy0+Z5K8IjKn7CACdg
gctZUblNAOeAVUSwZ4aJHSH4iJzr9ERPif13KmCJ/7rwsG1uMGQJvv51gp07
9uNfewNv6QIfFjkFTZQrB10zGUB3nlYEm9ORdWKxtoVQywGouUkCMJS5h8ku
vk2tOMJCyuMHPEPU/Xmb8y/LPUZWUklSXQESCvvSU7ef8KfeUrpPaQLOORfj
iTSL1lkHqZ17pJMa4ZAgjY4+WhD0QE1docEgGpwOOgDcHveKjYPs6r93IbQv
6y2uudC2ko/oD9UcVYaN4torDJ3tvkGNYnHNP7jP1yeViyXhaZzGNCZ1Ux5X
v/AUUHW5wYJ9IIIX4pf0aSSE/U5VPDjj0GLL9OHbvzW9/yqvKdRAaIp/NUBX
IyDOF72sNyN6dNJ/2FcgEBV72uDm4J9fqZebwvjP/nNfOmI42bS4onYvqA2I
j/aWsVEKKPfBgvKxS1SpE805Skr7h/E6vVfC8Mp+VUMJsrfJ8GhL8EPAibPj
JYueYhXFdK0Lfz5gPm88wUKKVaYXNfuwtrmnvCKQq0XPgMZt0PUpSZluAD1t
mZYvIVmy3sNXxI3RH5BdGbDPAMbTL/38srBM6uldGA9SBQXjnSbKzIGCzPxW
IPkIFF7XSl1FV6FKqce+YCEQNWgQAOCCz9UDARStvYQfZPPmWq4EdPbYU7Tr
vN7JM7uokHMKtUj1Ynrl2i1JHX1821JTfcclfSh8gwiIRuEELj4HSQbm21/U
TuNw9nK6cHDRi2sGoK87TELnJGvuipR482Szy6pcdpvvAkFr5Pre1RQFQr0f
jjZ191X4KNBXU1b9qtsepNDEE2dY2O4PVhSKm24Gr0ovM+QSnAtBAHurnScO
BWJiTUIslZDJo1mANpH13TgHEcgpNxAYJcRTmNlMhK6QrjbFGFDqe561peUs
TWGAhnRi2HXtolobRAC+Qy20pd5k3kmNoWJXvwPOqkjwc+X34hCufQ7Nxkmf
/j2Pe5YC4rExW1ufPVZYNZwlC4js0bZ0j84Qf8fBg8lB4+zbbiNhsNZQH9ME
cEFMQK1Ax+N7J1H0jDi1PyyqoSc4fEyq4eKkAtzp1Y+MROKlzpc0BtFCAWpB
fa5XVbi0GsXBYAsVYum29S6eeEo0PBoeWgiGXQliuTXFe41k+Ryz7graPeVk
hS5y5HUZK1eat+Q7Tsj8Rly/jDVQlGQEvKTklkPdXo7E7Lb7Ozvuj9WmLo73
uI74HrVv7XNHBmN2YGgJlCRZc54fbShf03azZipxB3lZjnq3RTbv/GEhwuj3
6Vsp46GljsHtQznFKZ/Kfd9Ub2Emu8zF6HqC3pl2bK0KJjuXgQI5wBVXxmYt
3EDtca9wu5NZpzbsjAgGeISgbCMMIkOHmBJFYMTVLQBLq8uChv3I8ZKRjsZz
xKJbgp6JVwdyt9nBMrQbXJGYL7iZyQfSUPGkAjDqlUIOvdwE16FVfnLnnOWt
V7DSNRZGdq7ytfv5V9yZZAQmbyxLe/ExfF2FFMVZHRFQfV1NL61C4qzrDiJ2
yH7QRQSAzi78dXdY/8Pm/pum14qH3eLhnFYFVY+u9o4uNrotcHdvMJIpYeHO
eoaukJl2JECvE4bLhzsfrU0b7jC9G6eKIqjrWU18XhTPZcCfeFn7fBYi/JJc
URnB1M8tPbyCAHGpwvb2FSnhrTIKEDHSYP3RilCZ8+cdnExNJpIfsBKl5xxE
k6NTsHzodz6d4jSy1dZUOi9kkz9IdVD8RjaYxErE+EwvhHf6bJdjNwYB0cJ5
6YQJeojNiImWzV3SPu+LmhgsSrRV/b1NMuSYoww5sFZbEGIn4P2qCgk/mDL6
d1myyCgH4TdbzQwWkfhJMr5O0R/0PcFVXBQ0D75a6CYr26ZoncCgBsV4+HT1
fD7R2nXo/q8aFdVYwbLLl51Cudv5/Q8YYAlxIeoWoTeWmkmEY6tW+n9f3R5s
fVh0uteqD/RKEiWXp2/NYYt5xYnHnSm2QcUDxRd2LJ9jyXlxOLpV2ZruECN/
+ucZE4+VOWYoqllcoYNcpuMDUmzPotU3UB3xO8Kt5vncX0g1iKVw7appqbIU
tUGYW3n+OLTEU9cn6/72qC5oXHg8WWr/wLwk5PmuLhEu0aaCqcVpN4QQS5lK
jmmlrVQ0kh2V8j5g6sIre4zUOgflPgEBsihNmkklx1SRulQbMpzwkqYwLEUp
Eis5EmJ5tqGbtGLDpAtHCF7aWDkJ8AsA76x+oZHYzPj7fW0TKeeYzCIycYEC
fdQXwTsPVMbIIf9LOIbErY/PI8JUMlVEfQX2FDk8+GR6btouRr/RQCuzbuJX
xqlDQ732BnANcoiq+qF9znpuh3FqSEa36mcDfOTDmYRiMedmT/MlWwampTX6
6OgHQuXYA+CSyL4yOQlNU3KUfmsrhXQcu/vvl5zycQ+m9Xg7DJ2RoQgxoICf
uZ8S6zZ48G2Kz2goknqQGNBPhITqbEqxYthsc/+Yldz2Me9RDyjAXGQkQ9xr
27cTGBHJupPv4a4hEeFv0uYEbom1pPlFXTiEe3Nzkkmr7SDc+RLV3LiqiKCS
0/qq15HFVeN9J3OFfbSIv4PD6VMZI+rpRZb+smhYL/qGm+N+Tm2l2TzFM1u9
/XLQJx4JzdKrPA614JvFLfkqAfA+du60nPj4tdyFuLG/y20GSkLQ0nOQnUCE
lpvy0f2CZxDbFpD75l4sR9T9lZbjIDEs6U/30PVXFssukWl5oTJnNMBYOU0g
xRIURiO/Zdkc3Hl2UlT0MPL2EufiwCj8r4geIELVvPj5ekrSLwC8gWEpuzP/
lWTSdTz/8bYW55K9f0BKwNmQemInXDcR/MDA+y6ca6O2N4RkFUit+7WPfGGc
d68hvyw168sP2yeLi4UgCPvSY5IeuQstHci55wJ1Gox7WIcecOBgOswRJm4m
Ag+IynynfKCaHaS2VSF8qxcr/qCW766uVIwLVxiJd9Jyp+QH8aPv+2Vh1p9e
E6s/FtkNJi7UAnvPaUm2Wiy2NHG3Wwu4e+GgtrRFwRAbBpd3QkMXat6CtR+O
/A1K0MwohOjVReKI5ineV9szFCtluE08r18/W3W+Vv9w2YlwokzEov0UfPDl
iXcwOZRMFmS6AeM/bygKSdbvMDyUb+FJu1XQXBHGpEQX4+T/qPBjEDXc/uxb
/jH73AEJ1H63FtdaABrhqpnN5hgRxgj6STwSFO4q8KRNMLLLBJB/I0DSTqMd
6hiv8Oos3HvSQh8xCZU5MWst6G/UgbIdvYjXpFNhlGx/lHEkbULXqbiuU+U1
vbchGp/UFPXO6qvzjz5qB7WUFXln2KjstPYt1gbjLh/HT+KHVAaMJB8qIqJE
OFzhwK+rpi52uEooHCttR8SQtEMrxGZGRjIWw0Q8Hbulvhgr6qN0OTHRQ3Td
mCYW2jsg9pzjqES7zBP2EIU/YO9FASezqwsEyuVExRGmseOR7FDWqFuSoFyz
Ilmp7phZZZqnlbOa7JK7QGKCgI2TQKb7VqGeIvvLD9bidrcbgCr29WMIaXaK
kRNh0p1xgEp7OzJWkebqhTgy0tD/h+aaQ0OLfi6c/DRgchbAAMK9Y667rrQo
HbHaiKPDyAszGPA2OJ/9/YcV4y4akdWH3Rjt5MVhn/eC+GevklmqKhrkKrXW
gDUlwjLcG5FsdCMTmbbtDrvBBOafUZEBCbE1z38Tr7qJs6Vzfgaz5C5kkyPq
aJJBt6IDCdAQU9dwhbxa4vFMHDFQhuMWwX1tcQSsG7xs10fGCT80mi3eDrlD
yQ9aEw8mkKE5N/uEZTfBmYx4+53DWgpvTuXgpNzCZx2KKkalA328SP6DgLjt
KsCfm08IVJkLG1rIDX8CAJG7GoP2Gg6pTTeaCGpaLPYnLSdBeiVkSjs1RMPg
2LTr9F0WbjHcV1r2+9SZSWk7t6U4PNWonOAISKlGtSZBinGasU4XCrqip7c0
x1022ENBpoggeAe70gxsjqBUYgcyph/p1ZdZHsvijH3RefJOpzf4QqmsrQ9Y
jRtlEDeAxNBLQjuf8ccK0PiryAqEet2QW2sg5eGN7qRI/xIPJtAqr0uMIc7J
H+nVVRSAIVaLzUOOeY8etjVJsVfJLS/j43Ihw8cIoK+JIKP7IehqF8yZj25z
jWz9PRYdoSPJAZzS5XMR5rhTrUXkqSDpJ1Dmqs+uSxJBrf74L0Q6fEMEsHm6
VspnqHPBMjJCInWbdWhd7w1Pswl6Kh/3kFhi7hyUj+zSXeYTcDI8LrgfbW4d
F1ludhADd7WGTND7B1EQGzk7rG6EsgYti6cOd+qH6a05F6l7YsYm48JGKfvA
h6wJpVWd94wleIZLWZB38uF/K7X5D6kYWJg7K+ib19Dkt9riPSthqV8NjS/Q
io1jfFc3/T+Irc+iVLGcnHoyyWO3EALJSeUhYcQFimoNklQF/jQyAgej6RZa
xn3NTJeuLOOG6WvYK7KDo/u39bbfF/qUfyAnm+fJbdMJwIwlR8BmjwpaJ8ow
ux3+t161y3fbna7SZiBvUmHUkO1x8+/A1A1KDeMmayXxLbC5RNyrqyO0/SnO
Jyu2KZJdMfqsXyX/lgJMg8PMTkghiTtLB8CFqx4EgxanaMhzh2goSE1xZRXv
eCWVhvJA9xPJTwixygmXOXBOBGu/ki6QXzISKGVBQLrtqy1kBCRLHrxxHgsc
AEH/6GgLOmeoWyQGarEZsf4fmbWdZmLZAUQIm5/3euUFay2cgf6pCfPW+ehW
dFTzP68bxYgUmxRNV+rMERI+SpUIOgI8S1TZgERoSj6BXGl49pC7szRfJ/q4
0slZWV7xX22xlTzZaCZ0dSyd4pHrDbLbRRLlIQQru0p4ULwc2gPXiaRfIjMB
oqRiwPKK5yirfQCpk6fAOdlWBcj53dTKnJP0AFv/QesN3IXfDUIUyV76NEup
y7v5HsWxvV+bHXywhRr6SI8p7PAl4S6U24hHFZUsAvviuD1BvtDUEY2xj1rD
GHc/ir3Ay433As8W+fW/XpO82B2GRVbn/M7FLRtORQhY9UO959p+Ps/I8xLa
M5ls+6x7QLflCDMuEnVGArvf5nHHuwbq9/cCemiC01rpS97auei8ethHgbzr
y5bagtjSPwUjivIVM3RnsIg0GAhmq1Vg33CE6q1YhiyYzfTkvYbJ1gNjWKFG
ufTMnXTSJWuQH8ektEYFAoH3I86t6Y83g70Zdui5chH8vrFa35vzTxwu+yCi
UpwN8x45ayLZAg1Tbvr8sSWy9+p8Mj5e8scXJPbkSSnsdgAeTR42tK/mXKRy
8VfTrpniW1r/JJGRwRfwRM/V2N7PhQph9RnOkq7iYMPrVb5dpwAO++Sxroy4
iNzbqruRpXOSz+X3apCQUH4WlAtSu9MH6xCfxoRV0GNu0BBU90UixyrJxYJ1
bNl4Ui5BDcEtzLqIgDOOigu/q+pekZKC3r+rgepuph6Y1sHv1/JrRRH2/W3a
TTKd3E0GkVkqbrSsqQa6F687mnJ2hJxHZ3IgczELZiOV30iJLNy+VeX+3V72
A8lYWOfgUt5bpXmDbC1MdSda75h3MS4m1kk25XjeryGNEJqGxon+FAaTQcYv
SCJq954dHDMAu/j/v80vbxMx5KYYpPJNwUmhPchkBNglH/RKhsM8CAirYors
FeCAM9ZAV0F1LPk4sF7uP2REOymg7CtG8uuaKguw/muQZV87TARIlv4dGXOi
GN/NvbqIzmrtof0p895oHeMktA22WWOqN/iBtmfRODNey6Pmj4hNZfpMu2cm
kbuQ9Wwwz3k0aCh192Z/P2ILjucwUH+9NyPzQOtsKEDD0Y3ydHbEdQ++WvFl
L+AqnpnqVDfV9YQfIM4PnFmbLOEK0N/BDmjDevkY2t94mX+Mfi4pvEk4sMg6
6euKo/sTeXZdLeMZLEK+dYMnV1L6+zGFBIXaJlo3JSK5pfHzBR+JW8qTCYdb
6pKUq6xdTce8e9FvV0IrSaVjL0B+s8dH3Dadwa1F6ZIF7CuU/W+DUB8NjF6g
CBuxcKO1Tuy9jFtpVQwj+x18oLb4BBMk69nO95PDQ6blY77cW800gYVjdk92
YojXbVCB74H7MQT8jvFBGWji2sNm3H067AFiuQrEraT4dVe289MIedohRO3W
mmnkqAz5G8E8MFJS8gK0dj57SihbH5JsZuoOD60JNicaD535jlz0bKJvQsWQ
0pzB+jFMEBAzvllBexDh38pnCNXrSE/hmEm4To1/z4iM36K28ASUUy6nJp6L
FGOfUCHwTFFlf+D3xWB+lz6jzydgbmP2dFDg2lZL5lnTg08lgYqB/4/rb2ER
y0qB7DoTgYtO1jqQuODVMZsBpxpO2c2srG+D65azcyDmiBzwos7N0hPOxYPm
SKFCqTfPjszi3YBktwttEM+Zf9h6G6N/4e5QjsnssgjUmbJqHioV1WiakgqF
RySb65PC/jdYT7LbeQKvozSpx9sgN/UcxQMPW5oza2rV3QVH90DydZ7CcQd9
KzuEcxToBljVsnsqDhQUyXMqGGEU3JCW7AjWwS+pBzOqYFNyQAQyduJevtem
mkidnNRdq/G06olidhlftI+6mtjFDA6fMQMNFAto6hg6PBu8nEO5UO3t82Ve
1bMJkQxnPYpNl9jR7duHS9mTgyz7W0BsEVBU/nGsOHGCWoDqhJxxnJcEOUcY
cXH57uDPzgD+zJlM6mHCTwV9vWcxY6b+0Ru1zMlbehMziOH1tddLIbILYYkG
ltDkfgmSrlNURUJOSHgR8/w4A+6VWfUrmfMXNc+PUcuIbAeZombKULLJhR2w
lu6S3+9uqQNfTA6RYyjhUpp/g+T3t9gYx8jr/26EbroJGCexHSkdLYpmgJMj
lSDUbS4rKLdsISnOAxLea265T6h2Bbx7dTsVZEKj6CCZz3SS8LfCRyl2sGz0
VYAiudmXYzSCzpxmcwqgzhNH17C67jOqpvDXcAWpKCPKk1VIPJwampn2lTb3
0K9ZbaRK6A8w9Q2E64YJFSzaIPT8Y2eD8wWVnGpvDPJlMHwSH4d+EjmzYd1A
FlqVXyCXFCOnvA/n2h9VeYr0QNmZZw24rQGjcWpBZ7wjQ3uCFl6veZNhmxIn
qul74XevNUUQNTm6Gb8atSNqgYRUX5PABtOk/W3NPL44L1gf0+QxKc9ze7mY
0NbKYiQr3VSu0dfsjv+0WLJhSpRcJ73RkEyk/6scUR427/TPShR0hhiUM7bC
X6vJB09dG65v074SEz7/qeEeo/Arsznhdi1GzOKg7ebXc1kHPNVKvJdwDafe
e6D8ve2gAmo1zv70tatE0DOIzvnE8zjDDBRbl7e+TI4iuSo41NePKE6xiCzQ
JlAWXK9SMxZWi7IfgCMLwED/qRbtF1UnhljxK4/3EZXVCuLuXWZJFJ7n43Ss
4Edq85HU1w+zTYRqW1MQR1/7vEHgmtT1RkDPCayRVZ1ARIDbvhJZRWAxGEU3
VCkxhM1pxUvtGQ7Y6FuPcfJ19G46TfkTLDaDJqa/9s2QfDuSgf+HIGM8FNhK
qvrc/XWOSzDMlaSOHljTqQSuxO0lzsi8gNBpsBqGoV+z2VlEgGQx7B+O9wM0
y73finnBUW8SVUY50e7fRDXTIht6T/P1wJQuJfRbdMEnEH4RLPdxpbnkUN7X
Jcj7whQFSCM93Y8PdmC/Z3UrN+lS7sM8oCL2XoI5NWtFvEXqds6OAAlqkfUM
QfjMbkTpgseUiZTmbe9TO1jhzob4To7zr0mMmhOuP4tdgAYadjeNmTAZ4pD3
FBpyYkcibFDn9atjVWb0fmPAK7tezQtAcvIyQl6JwXk2DmunMv1LKaMvGBiP
xgZzmVlkb4TbEOUdZwzBG/dRk9yMs/duAYexHv8wVvkxAUyZ9nIhUbEZFOSb
rOmj9+EX/CbB07pK+BFRNWBvuQayPjJxylVxMMQ/2FA9bJeuinHo7Etmzh8W
kba08XuQBlFWli40tt4mKrGkwe3t2ZNBx6Ustmu+StdwW+GxJQI1A3kGq0SI
Deo+ju0qJ8VumT6UdMVHbvh0kvuivO2cJUJSmQD8B42xVDFJv9at+AcLuGto
jW+J8iZ8bMdglaza+qdLDXC5XmxoDfXzZxxDkaMiXzG3pJkRzEbyOoHnCPqE
OfbJ1hPKnb0sVh1j0G5RAeW+23pMoYoJ+CM30cm9PStAe1TpWHG6qKhJD7NV
3CcbxtF0cS/uAIbR0ItmvR78stfKnPzdVX0lxd/duR3Exk7nvdO6OKGUZ1z4
5kfkWSxaYEkT+Ji8piOW2EUgn1+XhlaImqiUGUEatZRX8DfJKzc8F7sxwyhB
IORjuRrtOtColZWrLlQS257gpnB3ZTe4gnChTWBiqH2IsalWCI2bxj4fkIkl
+0/kRZfZb3sQtx5xP1l/9E7vlqPbwuxUKbD3KCX8SERZM5Wabrv7RxmMzevu
ypgxwxEpJnw1F2mGv53g/adhSOYmt/i44c7LC6/nBptSmUCr+nkQ//FdvdLN
YwXbYMzSJzSQEjletGGKECM2VrEISY7VyHv7Ttalz0pKZVsXHY6BxeQUuWXX
2t3wicxwuBJSvSh7JeD5rVo/f68xMi+RvOTYsEmY6UEpmAaPkUvi7PiGwjCU
EiT52O8NM4E+mesljcXpSiJL6mOWCIohMXP8xm0s2vvP7EIb9WXPwNUNFzFx
3aOoMVQ1VDB4oQbHFx6Dh3ol5TrRY9x4H/df2264hMb5HCtyEZrY6nT/0FlF
1vFo31yyh7bjq5agV9IFn8BdxogEMHiW95tK/iWfaqepfnL/OdNdB306seAr
NHTxxlr9cXlP2OE1f4JDaMw6qIppixjSfcYbSx+AIFl/h7G8u8pfD1X0VgiR
qKjM9oIeX8DLh2N6cI9kJvMWUvfKuHW9dH5zGeBldk3068BaVr9GvfNtDffu
/dsXVrdDlX+pRB+RgRucC/QB+/CNeF83cgU7dWjo6OWBGdp3iR6IGYiMDYcH
sST63mwQ8UNbyqjLcGaz3k+lFHbvmOoKv8rzv9l0AFmoIVxN58frKTarqijE
STJOseepro8xrsur2ILZFPXWMOecuu1EK5tCSNdxu/CJc7UaYjmvJteNdNpk
Ar1/fkkPEUFmDaJtbbWxDPhwqWm6QJZjAfd7yN2rjBLaImcZ4+8rdf+7LUez
arpUoR5yDcQdiONjoPgVt3yjf7q6L7eEiHBl4L5nEAfrumx/+zXJT13l8Zqi
wRdunvr7JyaxsMnDiGl+XeQapcPGYsOBZlWLH4vrADZpEDad+qCFp8hapbG3
NLvtRuqJVYqUEimrnooIhnqQslWlOztfBQp8JInDI5Xd+i/fBnWfPXxfJevI
LNWmxWrJf/N2hzWavOKPPY6nMEFZ3cPVLHa5V3YBRHS5EJJ5vmrXpz4GVIZ+
R9ad2/YjhaukkpbLtVoYOXPLDCc3Wdd2RQqQoVfwphTu6+Q9+9vFGlswQ+/u
eM2iIS79aNyJ1HlqZ/KSOgIB53l2g492NM8wSkB0pjxZVI/pUbdPABzdB1SH
Z3QZSRzV28hRTPTfiF/TL6nWMlHU4g2/mzz6e+rnqIjfzI+6Q+P49nX3sFiZ
DCTTsOguwt0dU/CLTtvmyHZpRZDyxwYZD2s1jAgQ19cQ9GMHJ91ypnVKJwBi
xpzG12qE6ZkAT33pjpeqQYaEEdUf7v2tx5gYbYiUB54/NnX+/5Xj6aPAuFub
/+pjJhGIFHsjtx9HgxqxcFwL2hsCWjbN/x4x7hbvBOYl+mFMJSlBMng3HUMe
SuLSnicIaJgevcH+BbNCkZEcDgclJaNYd8odFhu9aEA0XWh2tSZS7sD3xaff
gfOtHVS8ejl1SqJJyL6vPdbesVyTJjylAh0O6IWsz3aMxoVEmc3iOBQJBKR7
2FeCWagg8UDnovaxWNFmSXjUeVVV2zdyDa3xyxmRe5PBDHjg2pOPzYcKNhfc
azPHaQUcYbK7Nzh0kF4zBvhPiA946r0VB+BDGaMEQQuUi4nub+20hUUiAlwE
uwwUMhzwp6wxTAeExY21YbbN/l7y1/IdDvjmdUs47ogDvBQjcGJ441Qv2msN
hLEnmWUSohr5+9GVTyCNgS1KXvOt+a2OjP1JWjirmsFI2SH1gRiVU73YZHOC
Dx6gqpcJzI6J1ikxk+EbRIOpXZRD8gam4b6i9kBGH1EH0Td566EdUCe2nDwd
5VULI+8tQGXhYAX2TCFwkwWyJxKtk+iyOhVbevjxMDaFIvadUCcs5/TwGdqI
WCzXmgKA2T9lMB51P3+7+pXpGbVPpDBDWdfRzjkKkQHSs9m4Xg3JcEWGsNc9
Zl9SU8v+GuLBeumi4uf48DnuAyhTmWRuvt71wo8SZ6q2swFbM1jqTBJmA0Cx
FMWlfN3VxaY2+4Uj6uGJnLiAKFVkoQdfMZsygbNJ4lvZtq+d6FQle98wPqab
lrgyxhABqZjrseDIiatksufr6P3TXD5eHJ0sQUr3iuRFlFoLkJwEtB5gLlqZ
XrOpNy94kY2Fyj4+niT93PmjoGJJJurZWtxTh/81c1fMfAYDLi5lNRGUt3U7
kXnib5+3kfloqYQUdj3p8jGC78aVr/zWuROrrCZJe6X8wwZ9lxNNv4oElRFw
ON2nvsH8QNtKyJq1f3iyXu8wWnfAHDsHbMkLhJOn/TiygRJJzvaEEVtDBg4b
guN3vvqvG+mdz/N9OKBlZdANPkASyh3V9/48UFnX6bnm/+6rnVY70wo+xEMK
2q/DSXyJ9vsLONwlrRnh8ogm/z5x1pfD3GsQCUMvwbrmez9Tj6mvycT/ukMx
or2PwewFe+J4a1jjKfCN6Z833i24+/S+9aRFY+pA0qve3ZOfQ5+ivYXbNd98
h3ReUY+2dAP/P0caz+wHLu3EjqXRFnBH9qDjrrnxuXOFzKJ0EQzzR3K3OnTO
LJOPTMRVPm2GIu3/TXHP/8igd/NaaMp7RlH/nyOdIZacMrMX14gm4jdrj6It
uaIA/f5q10+JlDH6OWfRgdILHjORQ8uG1YDeQYYRIUxPb8T/txQkIHELsziA
+4Fe8vRxWkoHdBCF1aunmimRVZ+g4OBTf8HjXEYGfb6u2WmnvvPTa+dJjLu7
ZegXJ6F7DH8CliTkbQsCJ269d6h3u3UC97blHGa1MjObAucKTBBsjWHafM1t
cZVzgwjV+Lt60c/RKHAdH01B6Z2wGqSM4pBK0QAvDMtwBU48/JyrE6mPK/zN
rOEZTsrzJg6JBpYuWo6VIHJsQ0xlcgV60osSASI7olKdR7IATpcwseS/5uuD
IrmBazWKb/+uvMh+PyW2dD/0gmDkb1LqZPkFL5xeJu7f2Q4/EE/8BmNG8Xz2
TPHNjU1t0Aa/OAdZPi2u7gom0/RN1IMVoKnIdTa9aaJvDasTiFQJI0DZQRBw
FGw7EgnoQF8CTSjb1Q8872w+JPJLtKOPb+SSH/1Xz1YtsBGFKiKftzHG6n2b
DQARpbDPEQCuWY1iV1roYcQ8SniLofw8kpgeSHLuvAmY6dCKfguI5DaVyWYT
QcANykhf5baCIcUKpdic/Ni3chh/o9q4Sgh5pXdQ8pJCRJr/Kr3peuRwOajQ
v3Gvr8E75gnzekjg1p+Vudj00pNz5gRtCIVzNiVz8HgWbkHGEOKMhFmRzozw
uYBPDscO3h+inpte+XLJTJwRlbGW3QmmHbD9PLv3x6pKi95o2vV2kSw9uXrL
wpVrzdgPPyv5riBcObk5Ix772O+rvUfXjfJ+LJOOZRJxM1e9gAayp/xMn42z
/HF6ICPjbEtDnxdN5QWqr5VDnUsYttUhN9YXcqXKj1gdXnV2lqxVjOkTBwPr
dJeGCt6Y0BCyNlHZTKyKFVKbebm++bilQN7EnLcpAcw+zgv9SqMCEN2r4hn/
umVYPQel/x44XiQeYIkMNR2iwQoDHDxQAalSgpxHmBnG0KTEIvOxssN2Aay+
RXp/r967VgVa8oZxKmgr4Sel1KJfZPKlDNpb9/zLn89lgQgfXvMJfTtSQXSI
40JUCO+lz3nTsO8m27BdGtfTqigbljYZm7xOY7a7Vol7hnomyi+FAcEFNj8A
92jm8YF2ng7wALEdm8/KQ+1LxzcF8uR6NqpjPuPA22/0QV9rUbqZQnY04Svp
9kFtBcUJqC4n423Jp6a0AuIe/dCVxjACNgf1FST6H/IysJLROyDvbGq1vYrw
GeqveEl1Q/uPGGfjQeW/TIfIQABjrQktyMWhhIafTKneNT5EWwChycEv7n68
T9xZ/gJpUbQqZ5/zpV+F+fXAtydLL0Fktrr47NIq1xaiJ8Q0KrcZpDlTEkRQ
1aZ/XY+FUD97hOqHUNbtHOeH3rydnO1+UgV8Jgo8wzAHWINQXYg0REZy4PS9
CPSDDPizrwdVIeUv9RO6eqlk7xxLpxd04eXNvcpboriOCkRfz0WYcm9E/S0f
UOToajQIIVEzK4AYjTbC+XfvdTSIwhs4tClMaRg8Kv9QtgHhUpexhnKbcyMV
8ac4n7zB/DF+/DfA+zysevkFotzmbiQlnp/oXdMyx9lHPy5tmyrgnNs5g8up
08vt9N3tiTahWbGe/d32cXD9XbpxqQoFdk6jgNn4qmwg+MPRjTipSQBEigjt
CFgMlhwVDLSO3w/v4b+Wgbf24zYT3uHRDAnJY7HqAFeSFpSLg2UzTRtD9OLR
8z8wr5XEYWlvEK2ymFNQwbsEQDU0xdCYtejx3pDdKA0Gnb/dH55HeruYWLrG
+McmRLY2qcRFfTL/QdLL5xJn84zvFDg8SXiAHHRc1nqCS+Qh1+OxmlR2R2GX
me4swS/Ze1IZRWQ4RZl7ERcUf8eaO5RRmGqnXW4BcshyqqP2hFfan+OU8qCg
ccgRcEmshqILyUYa9o4R51bpcRfWYtYDlbFOKoknvFumxg8xeUyu9KzEqjAj
9bMlrJ96aB6sNZxsy1L+mLR2fL/EOAaKPOmlyqbcaIYAD5i3YIjaN8RuUqMT
jBFoXXLfsjNGi+RfoYUgwEd5NOVQXYCqS3oBHLeTJiWGl9Yz1mO0p4bszQpa
AopSajsvDABDB+Yd2WldHkVQ1I6A7lpE/7mhJcFwL9ETMSCBsvdFKWJ46CHy
AXgy8EJik6Xu4eclczWh9sO13AXT5HHA/sE7ZlHGJLit2mh1Pj8+QdUXgax6
XqRcoZ1woYpm0pBaLHpOL3p5gUQu6BhQWljXNcIUeOU6GWRx5OoJJBcQdXQF
elhGxqw5iBZmL9Lp/Wxps28nmKD2SJSk7jf5aLFd+22/Pdy7QmCYpLMaPCJq
SWBxaWRGV8lR+FFq1PPoajMHO61qnzcOSIj4qUBQJmzFRXWgvbru0d2WkXpn
WmsevWtGMWqX8xIjjKGZv8IWHd2OrUqRPkAGYdICjEObJ8P62mIBZeCLH7AM
c2kgIIA5zyDof3brNmcbX5u9vpZBANZrG2iS3FkXqK8RWga9gfxNqW/6a7mt
sD7kLJh4awfTg1a5DXJ5cty0su8302p2xAKrMdsDkEfC/PIGV4GDyyoazqCF
SKXRUMNtMUi0QFFAEmwURUKH/pfKsdeIEl845CKIPg8YudAM1s5blDE53L6R
CA3qVmd+lu9MBpI66/zZdY5i8BORvCeFXMBqb9WSvZ+tk+rc2iAbeFeXgl4v
4oARwi7ycZzrRogTnQc7zB9sSVzfyBr8YheGPejdy3hi5BUPpm1qYaj1YvFv
ddU3+9xlHgg5hn1ctMDWakQ9QDjdLBf9cVMREfGRDw0RAZtT9iHUXMeo5K48
lweIXngPabL8/tovNRuV5xEkHAFlaYozk5oDFkVJepB5Ysm3Tg82rK49qASY
oc+gZbg8rGAmvC2HTMRFkPiOYZ33jG/fgaSalKgLhURZ5MkivRVQPpLqQ1BO
OAXBBYjwjg8LFGK/ecFS5XYBmErvYFozhCbYfrTP6Ula3Ycdcxw4htMGleRT
LzD6oJfLp9OEglaFxRWCWo9JwnrYvCnAXGte3v4ZKD8rvQTGF46oxg3Lmk09
S7bYj856xI7+HNUKFUGssiaDjB/0yFd4QUWcmIk2kzzHHM27Hy/Y53CcXAu1
3sOxcZnOe1bdvt63T61d1UB5LzeuAVdgGis2LhcTMgg4pTkWIkQJ/zaYsFrj
0PA3LY7/5FYpfnyW2aEtnaheo2+tVMnV9GNiHLQrO4WPpmc5R6PVbL+NL24L
HvcbnKlNpDblO2zS5pCVUL0smLvoQrGKK4c3q8uX8JUsIQR1d6jFNtaBStE4
BUSzjgMENFPE3bntjwIasQ4iHoQP/w1CJP2YPaPzXTBRS04g22I04/nrGGAC
RpicZCDCszoa7hjJsJZVrrsJqvVtDlLHIgz+eMiMVKcjENstgZccBtWocpG+
m5OfyXPYX62E77ixGhixEdjOOPx1UEz3ftoz9RIn7ZqgMlKSB2DH3Lqln5o8
e4yI1RbwGzYGzRNnHd+HUGroZgOaCKQoZfY25AOkE085THCHqe/XoG2T833A
ntva2891Bqh2xa1sq+y0bRtaU2Lh7X1VjKXmXJAjI8rtOScYc9+r0yGaZEBY
vcGX/cjt7ifwRxQECErm2P8030wG/O+vlVsX3C9UEzq83boKeq2VhuhwZ0dQ
vdXjlKBJWMVnz2oWtAGx9/HcwCq9gAq8VAw+AhKrW81KCbOqfjHzaMb0xgEy
ZojwzAB9PJM3cAQVOFAQ397gJYSY07L+VmipiqOSlnQvrD4e7UVexKOPpLmm
i4OEgR/HJ4e/oPAtXm7pjLdciM9aVfBrqJeB0YgLspTBiTKRzToiScqehTYN
j6wiFmARcsTVTzPA6OLZ4ZqFVm/vrY5pmkqynKy465ntRnV0CTekf2EBzEKp
uSylGTrspYaV0/Sy/2/J0vT7IquHfNeMI/uSJ4lUHGrOGNtTAJuMSQoN+5DB
p4AWLpREWRW6j+0cWZoRAJrIaidDTck+4RJk/Y1Sxkj5OyyNU3wc0zOyI52j
56sJe7pW9R8Ta/1bvts3WbM83wQDM0SgcezXTtm7Kfn63QpnVYgMnws2eqi7
nO46NZ9uweEgmozsBOvYIn1sXO/Apr5Zc2TeEaxao3LVv5Q+QynWfSBjPrVI
5UoceGuwpyHaRM1rJogY1a8J5JxmS7xcRMTJnoL6aupID50GuaECGC+SG3TL
3L/lMXlUvgqUrwf9tR7EJceuhDtgaVg7oYhQTjC3n+EY4yLMXTa7ZY27b6Gg
835A7OfcgZod2f3SuDRoX1ASoCtZvfcKVmhLURVpj6Z3vKiNDBfB5NxHXmPY
7FmaqGr644v44Yz8qQ0FMJR3pOwI7+bvyTX1MvocbHkJBBOHgmN0d7DywK0T
28ScWl6ymPOYWU8rLuqm6jBpQ9yjneaIvNjqP1E6tMJ4SWtgqMJ1EeUjP+JI
T2HL2UyfYPwyGFotVHQmme0iAH9oXjotgWZ48rifJ+gCc7r+/mEsR8hmJEaT
0taJIvkSDivVWWonwh+9I5SqYZZwCk+TLhH3hNE+swnN3un9JPm6oqBff6il
qgAwspaJPnjOlZWwEKgW8gFkx9k1xWI3NOrVwV1SRZSzM7+raXcTPWAzDll/
brVuWnY8RRAMYcFhizVvHsu1UIxcmS/rjIYlLwtqXZ39A7nL9H04irAcxI/N
W4F2+w113BCX+bMUmdvtN+TY/mDHGo5Vxv9inG7OWlbPcbYEqmJ1KR9bwDnu
xEL+vk81Gdf6V+/xSaLkbY/A+O0r6R4Su9WKu0PpHUBdmlp7seId1ISAl2IN
T7aj4/l0xOEPoN456x3xHQ4PrkUY0ShvE2xuWvO8uTvoH+rgRepvyEcHmMTh
6wd3Kx8+2t/m3LfPRJC9CoR7h8Uy2ADHtPmacWeX1hQEjDNT5rYzq1NbWdod
B6Sm8dKYjQANo+J4AX0G2ABzPLECLIYj/U5uHbdvqg4h6Ax2yF+gfjr+wHLI
T8iRGKl3jsHWLxydQntkVe5k9KpoUOQdoBiJlAjMjo1i0GqMl3FPTQimS5r8
7EAWcxZ3Z/8XTpd5Xn27ThA/ktBnFT+YP6B7qDUzqxRVeZWggl8/X5sHaxvy
EsWJauXW4MjQ3eNaQ2neMd2yUGn545A+e7lO5sBrCBO5dpXbs7li2LvL//C7
lETFvQCeh3id5opnnH2XPlClJA8u8Z/I747OKxXgQYCSSklWDPd7LqEFz6ze
PWp8ypf8Q/pKvZ8XaS8694pMCjJGQxbfuACzjgKr7kNcFH8vV1J/mofmr1jm
8iUWegj+Jw2jLbyFlLQ7CVKFY6e7vM5ReFt1P+1hHifJFe+ZDOm0u1UlajuB
ZoNaDjJ7g8tcx2e10l/275jobAbvfs/sjvSOO+XXupptDn1GvpvNO851SAaz
T+GuskTIgE60RGf2Vb+aiI0ABFbisJtzFce6a9mzLgUqzn7t3l83TV9rOkZz
HNeJaxvwH/mTXRYX4hEkb2DOSB74zNtF+QKjnr3sxqCa9C3rIzVYb+GoqEki
7/IpBa8poGsTBm1aLTd0glytn1o+KISPnh/XT00tez414gapcLgZyOev4dAs
JQdUSuFr4BdrmHoW5N9Qf6GQlTp7Qal18Jmj9ZOUmwjwxFk14/aKXJvxx5vZ
1BdooGoFUZP6RBLq6dMjatVZ9PWfBqHZUf/wNFNzRE3GjswzRCaW2AiLAx7r
fVkn1UisHJmuUVeecKk4jkCo2P0DlfGr+sptIHqs7sdeUl+kOVHIMmrkj43C
kfUIbh2XvZjVIFRoOu40CsSJs9569zXRtehfb4TifFYO0dB7n9vdioI33Uv1
ZTueAgGefWs2Si/SO9x681C1+RDLCQhWpX8rc+k7Dfu9c8U413KS12jGIiDB
gYPkdZ5sgsbYrp1NjIcyUebgYb/CToA5JjUdvqb/Xe8xcb/FS7SL38tamngs
Ul6DiWKalngpqUAMiXxEd6oeK1db+cJgf68aD4gxJzEoeIk5ukapMwW4O7CK
5aG9GKWu5bnysp7BZHmc+piuajSn4wBrm7Qrkv3DR8B9IFnU5Ws8xSneTyMU
3Li/HXB9qCdNfWncq+43NoXhaTnHVRdchXW1STjJ0f2wb7I8ajqVhoBk12Tt
N7p0mCPXGkQQVq8GsXuX30Wo21LItIC+TWBIZaPCJBPbeoRFeVtaW2fiWwDD
Kiqxly0jZdohYdHLkTWarxj26wEgqp1oy/iXxTpiaPf63HCPOsU8gRNAFZjx
eqG2A9j6xlWBKOsLIBYxhBIHfiy0utCiL8Y7V/wcqeQQDoGVk34oQjqyjuNv
HTe1nvJaaBysO4bfLNzPPuUQgw1yLrt/5cEX4Xvn/bTd1+tJcYDgeMewla9C
7GsAhrJfvgoihX1595feLMfprD2JFMWdZDG0RCJxgCu734HmkgIxaKtQZXuN
wY2SSEjpQ+x8KdSz1iAdRvNXFs0xUwedsUzM+bjCi3XEc0hkkfEntRVFBLeR
wcWwCxLT05OUz975mcISNr8fUgaeaNpm/XJuGKgirCbs7lecWOtKQpfo/mJb
F8X74nHf9SndOPpboBJE1oCwugieHGxXbORYkM3zO283ZzAeGjjcUN0Zjcts
LF4v5omiBPoXLWzAz9oVFK5djdY9OvWRVuqPUTJp0SnfeTrr3RpxsMb8ak3X
BHbj15L0Ftr+S1VKb3XnpoGi5xJHBg+EpESVQljxHqKpdZCb3v4E4LGA4CzB
io9/dHlaY3VDBCNJXV746V5i9eCO25RMhYf1n9IEf9p36rzQLmjUob7ayAeq
EthUEgNWQhEQHstBhQj2Fjo5EfLIeR64Eq8GBCEpfHACBqO7BO2HQKHEf4r6
vOg/oCJXSTD4L7sF4sbKCYpsARMJjTFZrYHDSenuwOeGi/zgE8eWbor7dok8
NwSML1MeDnYWv/qOGYUXr6wxjW8wpFDLsYRTleryq5b+/3kfXjQg1KPCysY1
gwfwPMC/qTKoZBviQzz8NJEuDLe1n4FAcaRnHWyHUon+Myv7sHt13aheZlEv
CfZuQ0wkSpd4lITzy4CNnpV5nvHF0JPefz9GwF221h7rLLkitCOBtZFMel8/
d2VuOkaS8Jw6CGFNaQEA0SFydFnfh/I6T2Ewh5FBV+b+DCIvjmQhPzTN0lry
4MNbWyb4CHV16YbaYgTftT5eEiqGTFRrBPK8g4IfZKVO3gR1iIkJacDlItZd
QKPvMNQSV1tmVL5x+ynvvXjklkw5Nf8e+JQr0kWnNthSbv8WhEqKoZ22BBeH
d0GNyFFsM4Ofqhl/tdB19BOoB7qIbAsporVs4CJMAq93WmUkv0uuN7/TLJVP
3wcgNcpSncJN5WVsrG9ukoecNxA+jRGNHQOM2vB6FfUKTaZbcCvr6QSfCzLv
j9yL7TslWke26eeFCWQnzm2vGtv2xDL84gEBsdBXufk5qtgRwUdcLZ1dBxeo
BD4c7pXYS95fGX+T3sYKFX6jWUQgo2RjZeBw8Fo2Nnltp8O2Cd55NzAnClXS
V6IA2lUj3b5XR1uVg9KtFZ6X+TRxa83ffkM3gfNpe/zc6xBIx8Ihon63kJux
5apkuO9O+nbjTOl454zfCHJ3JUc/F7ojzdHxinQQ+q7rhHqoYto5TRSMJLcj
5FvaZAjYyd2JxDcdGF/GiZyxpGytz22oRC8o7UoS0MdmUMn2ld2/52L2vhwC
aMeXG8sQ146Gj/JWrB51f8oB1kyvef0dzS1pFIOpC7mz6JObTtXZbu1T0nhc
X1V5mZLLI4y5cPnW6ZHyavMC5xCzGzWrEQRk7JMeSU+FDE9NPx9N9bj58+KN
YhY+sbKMFJQRKsndeLRBVYamUwzL9+TWad5Xw7p99hUyQRby1ba/M+OrNEvh
p7AikEkPZEmi8g/gUCyj6fN9agRms9oGqxB2HvnuUNlLfwxU4e214H0vKFyh
7uA3ZLfVghP5umOk7V/4DauvnDPm+R2T1YR6Mjq21bJIpRt5gR/2Kt74Fodz
29UPwnU5CkSjMLP4X7Z+L0akZ7+AMsJjd09LQ0bpoBSslnjcgLn/vVZ8et23
So93FEynyFolKOM8iLYZGRHLGlGG4nrwuRFC6jCAdY7L1LgffVtkH3zL97co
EEdGpaSTOjV+BzQN3iY5+pX/kB9130G/tGNmttF7VPGB9s1KvoZG5A4fEdt9
Yp7UNbcD9uCuNH56vU1OMR+VC0dc89sexZdIEaDN2PzMCTctTYSSbgiJ+1Mk
0lXp5T1l0l784A42IEARCpspLzAg3jDkkqIzRNCe2oYRuptxcL3Vnjt6i0bd
TEBScGicdxnlbTHS0pPrNeKPgSofh8Url13qPBpGxMBq7c0avsuHCWSdW2Gm
lgs5NgX0WtTTEb/sn3lCoHi4EyZuFx13Xv+vJafm+fVhde/j0wVJPCDCoG6C
nl+ddwNS/OgDRqSEOaBM5f6+7CLEiB8IxUAWCJkMtbZAaOG7CjExQTPsO39x
168sRga7pYYy8cOZ8a3hThdyf30s9fyzg8dWGM21JJkNVP1XvreTYaNia6b7
UHtL+WtpgXL9eT5il1pwC6HZAXAoOW7fRiqiYhDPf9w0K5bdS+vSXpPWFq44
lb4e6609u2Ee/Pryvl4egnKjG6gnWZp1GV8k8Y1gmJTyvUxZkEKiCtsg8VEz
OpMh86IDXUdGIG1TsTzu1goSO/RN3ADS3lFzgCWD3HSVwyTsAtwg/NsuGZML
ReU82XoftACi6snkckJ/4fmF3Ih3AYbkAuYD/d/pVOsPQR7xbbArUBDbDyGb
UQlBio3UCJJd3CHOykY7NRWjM0EHsqHaq6YGCTGnCfpwUqapyv7tqqX+oSZa
9REGKWZKTc4N1TNYIGcmk+t/Nr3o26tjSm8CRNEWFCpYvYKZM+vPhcwOg09d
4p1fx6LkdvY1hxYlljCRZSv1KUnwwyzfFEO+7MjtEtSYlILpBPzvdqo8Mq9V
g9qE9O79trLck5nfTHfr0oPAY62+4V3bkcTAPTJZ/JEKaTqyzOVNZINbIxEZ
rme5I6T6xDcUcllIB4hUeUvOQ2FArh2B9HcZOq45LZhCGT+2AgBNMfPANcKA
EftutvSoCKiwbzo0LZe8AfP9ZFZv3pRrdzFbF8apkPw7a64CIwaG6JxUs5RV
cGM/EFOyIPA+N7y4/D7CMOWZcKPz4z6TxLNm2ZKbNOJgQJCP8NoBgo3KhmUq
66IU+BuXp0iBrg5+jyGviD0K2nLp6qvaw2ZmI773FXWFQLtzDd5fX3WjyyLg
lUhUZg6xcukllLZQRvsxFeSHEyhnqlOMbAwunmx5oqz1IYKbGC4ZnKfR7I/y
L70AH7b5rsivd5Az5lh1uyF/f2ISeEyQEhaUHcPQGSaTpDKvIeR2X2LZNmuE
r7nGlyutMhp2xz0IM50yzhBk3niUoHTPGZvh0kF84rR8neaGzb7SIE8cmoR3
vjM7MSqbxse7jDEgGjG7i8MSA8vLVrWBn6gtiWIoSOMjf+JQSfGBHUEPuaxK
HwAHAhPob5pmLiINEh3dCsFAmpVGfrIWtaQz5b5WMcDIkRYE8Hu+qj/SAXBi
EkV4f1x5WWmeFhlO4vKAyzjmHiokCmWJ0UKckYdQX3EAlKCLtM7hMBUts3sZ
x2OD6JhpzkQ1DpNbZgvVyrpX9IXmFtSbHxhlL7cwQbiucijmU6JNTNyxcOJh
gAD8Mb+Zfx4Jhc9Q1R/5qBdSaNU9o4IJlwNW1hUaN3gSbOQXh7EyNvwY0rkt
xIG7FI3iAumKPzT7BfXrQQgYIbZD86OO7tCDTy+VTTdAejoy0S8nMnN1z6yf
lUl45sGJ4K00dICWpBz8J2YfOx7l1QwyBtfknionAp12cx3pSMmy2uDKlb8Q
5G4cvosYB5uuDVbzS+kVFKWSoWHzFp79eJApVaupbXIybQJ2Oh6eZ7/FKxVF
dIY5G4QXGjtsnPXcttSsEw704tbeNJTI8K57o8VndNNknVqBsqkgushbUhag
2dKT70rM92nO3SdzeHWebq3+cXheofnEL0Os8467txnwI6JvYLS8ntK+iOfY
SQEgMi+xTSHjZ12uLjfS8uEXwkrbgi8KXsfBvhrYCJOJA0M/XP9lKOMlFtBf
Iutu1gqWntZwiIpEKK877zRBs+R1uN6/Gikh6Gzcp/yGrMeJpLAL8BuaDL6P
6fj8pQxJHjY/NnH1/FfJ8aRTIrmXk9QORR7xzB9lSOvQu2bkL/n8rWXU/WA0
F1uDa9lRce/8Dq47aY5mpkJ1LC8bTMk7zF9cMm9pAqMquqh5xhrI/vQph943
m66gd/dNZmZ2YdWlUCfduLTSSAlZSVb5ZW7ggOWCpQs3rjW+MS4mr5a27pVD
MNL1qDh/DxmjSRbZ4Yr7DPGqSM8t3PpbiFqPh7kgQhMjb6erKjw0MdN64Goj
zn7rGw59esHpm39+qnAQmKV1L+pfsaQiG43PeitEXL4OqNHji3yzHGkXxJmT
MwRhgPHssFckTKCH+cmu/dA0jIEdMDTYonVw5SGBiTZU2C9YsicWe5eqfyOk
l7NKjhKPDrtW9NExz8QqyeZk5siEfN8FyRZcgmOiJHu9qOb9o19QOMXpsMTZ
DpXPN1kWqa/e2CIwvoSWL3P/0/byFr136G44a2egPMF4N1YFv+Wan0qmuJSq
Lrp2YApPmS8/3CSLSSBXlETyGZGR0+tYkE4rmNU+r6ULcStEO0F/4i+FndB4
u99Jw1HxP4RBvjyvo5YENLHGS07YO28xduaxwQPrGOApf4SlBTdHNp/KwdgB
LtdZmbd+a5ODg1/slMywaTGZW9Vl5IkU7zNHUxpTCdokOh6rzna+d0ZEZ/R8
uTcsWhj2pkI9EatMw+J6SCEP6YXc1pv7plYwYQYN4dZ5xhOkYGNbI1wDmiKY
UdKtzwuUx58Kh20mF477haS7vG6TEuByF1o4NAjoFo+YvUlsWqWTnr+ulLlh
dy1sdxZC7ozqxUYSEJde592yNaE18tM9Y86wB+lHPZsnfjPA1eMS+G3dM1T2
Osjk54Pp0m0RhAhhFAkueFE7IElaM0T9XIwLMqesos9L0lAlfz4RwH/NxWVp
hnLvihWTIoUvyDIS9KMBp2XAbuS9uTTRvmXBkNLVAWOJU5t1TdmlMZ44ckkX
Fu2MUgknuqTM2x2C+xjygFZTFf5aIGkWF8ImxeqlCjaxvKb2XktUGarmb/F2
zHdEV12t8ObcJ34BCNcyfCeN4a06HscHI+ySVlsy4d/KF9IJTea7ZybieDkL
5fsUpCyXQ8snsRcfYHvwHTiZ8Xo5tD44pxFNJhzsPW9xMfsX/cMcC3/qmTCz
rzla2v1GegZGR8iP6lQ+4upJK5bSleiMgrcM967cypUifAxSA2rdYgJ281QK
WM7f9uA6bQ/mzL6RqFE2yZ94OR2uLvRnQ8bFgGPsJz4FXsNi0bVZ6afEjlUk
td/7+jItHDVfbWDXUD70Som788Bv6V466dpiSOyqdjCEgIDdJU2R9xnLuvbZ
NejM069NE1MMALRmtYO27c4X88cuvIS+aUhedfxwMFRrmpQbVAaPdmtuiXNF
od5Tmx256X1qha2UfTFy9EJ8rOQkywPBIBZD1MkS8In/H64rV9aOQ9IMC+gd
aLvdSL6IYh42X1PwWAmpQu+ADst0s8uky1yioKM56iWnEKV1rH5EYxhJe5hS
wWzuY6KUl26D/WQhgXfragUmQwCuI37SZX3bjGGIYk9ucOlbMqI8BHHiaGq2
Vtp85sRninFGD7LOsMRZMbvpZpefFJEvKR5xmU1G0A87Cnc4zzA56ijV5YLj
ZzaYNQtagtcmCtqUr4czHuM2DzAN9zsTm/VyLOaiGqgvT6QL+qD2vLGYBVfG
T1DjIYfwxWtVOPgBI5/ItIfuQGrL7pjaJhkOAnj8fpfwNGhjMnOcT9R8fDRl
dhXqlpFH74qvyyaFPrR5Dib5jN5H1eIX/PJddBl5dKKLr+L/yryYPKiHgy80
l1n2hpTOXAxv+jwg4Zwuf3dM4zQdHXgBz3tDGY2pxZ2gbG5wmsrCDI9GLjp1
KTNTfSq/PnRMOgGZrV1Cj88Sd0CZ5zK4bignyqSSECpMflKn8iQZiFU4loS7
PW9UMqnupuNTAwaQUDFjikvLFD/0DF+GPlDVL6Cr2vBLvVEcOvLBapFV+ea4
BOSvgFDvbAR5/jKyOaWJcLo58YgYbgUb6AmWEIX+E+cqxZuEWaF9DOaWbUh4
lkOv5zB4RAci5FaLpexgBw5SoOIxuHoJflQShQdAd/kXSCfGWHfDJAgNG62n
31C6ZfR04I9fktzlF+Wh8kXuBtgrRzxKGVqpPZwl5bxKHehqVsRlQzPgCmux
TYl30Cjp/KgQ6NO9gV+s4HfQIcL5lD//PXw8/IhdhjJaVNi//MpkN0YMvd3T
wj1UNFc1yDSFDuo6jQGQ+k/RFuGHbGfghKaT5BR76pF1VANQ4C+uoNaWAF0x
R36UVwqp8o0O1CoMhuwVAFyr6VbIwyOn/JeZbk5/zZhmYJbhNDUD5Fif/En1
JUv6SHxv4bqA/QcROTp8mT7KeTnas/PqK1UrxU4WxcMSmYZ8CR/mqcyKs2sy
q5+UXqbvmwC6bV1c7aNUp6QsTUPV9EuKhoaxlUxJboB8pq8wl5R0BXLzgWUz
CuCaufYle1TCRo6quTdcLKFMzIW6ubX1Cz8K/t1qDfFOmp7MRK/6RGqu+aO8
JMld/K9CUqLPMABaUcjfZh5JU/yIWQsSDgW/RHASOSbzdX+fld1xgT54PX6O
c4siYHC8TojRj+wHFbCXeiv2UORVTuUplvYSBAb0OBCvDN+xSJgR1zR9Oo/G
VvcoskeFbqMMchlq3BHXkELGzhdYs8oezpzhqkMustewmab9iugSFJIXYuks
H8i5fPYXi81YNQILCjt/SoCt4pM6uvfF5h8e1oru+BrK8d3oSOMoRuucvd36
5m5W3sKOOodUKg9iFDWPk4fNgSP7zay91izwA5lYBDYc2+9QKWDB1eqPOv7M
F7iVdoHoFGmmSS887T6NfLEqBbWv9rb4CBXTuClklH5dE+0MNmBCbsJivL94
J1/tQDYlObGPxYLlqz3gzOtw5GN4GI4GYjEnpe8mIiTpAzCtLHuTfQnjirqm
l/0rwgMi5XzoYJ8CI/cq/pvgMO93bF9WjMUHckjhtOzeIkVXvl3UNDK7Jnxm
MdF1PDG3ojAMJjwATTkyrzMTxU/b9vkX206x8YpuiiWPeosWlhI0M9XkVTW9
vhyuD1ei6KIHHiN6OgeZ/CptxPBLThYp0wN3aUu4MU9bwHaMG0X4vb5qJq1T
fqz3cCV2CGLA6Xe3qXSZSAK/yALXwSMd1lgAiPyhvM4uTGsLQ7EDzXJ0B9eC
kZm4IaXkcOKCdD1fZOlWCGasVEhf3Lztfxm/3+726EzW9qN3wI6/g2ka4+Y/
IeeM0kQY4Wzx7ROFeKfq70AQIDATbdTxsLTDeD++zZkQkbM7RQtvWaJ3Cebw
vf4NQ4kuCbspBY9IVjGO5v6op1d53cvLvQMLldAZMMNNqvwJi0iStLUIacBQ
TXOvO/cTkIOWWwAzhhoMvml5xkMQE3z1917BXTAhDJb7702TkRLVMWN3fu1T
lmz/0Mi0czB5upqoADHVM8l6Sc9DDuVWAhydA50it1KqcsAGYzaJtpFyvWrd
fHMHzjMi3beLNyAQa4pArDx+G+pswH3ZTkRvFqJeASY6gPSMyCPMyxV4kOWe
KSmyM+i7Tr6IYRN6B31YzzWTKi+NlLl3wIVU+GATdeMzLBty0qn0FPbycOPX
JwnQ0TyJ+yR04aHEceKX5LDYp/nHq9tvcAKdXoD3GMS2UNKjwIWFpjIvvS5L
CC7eOAxtsbXxZuaNSa9L89Msqa+YQaEjz4wDB9//VbranQ4cXwlE3iK1XYLW
PRTE9/ob0y9O5z79SLe58w02oUIyMfg6//Kq2+xaU3vRomWOWaWeFiUIA1dG
ODra2Qk7w8/0awOMnSOwadCxBDM4aoczz3pHhe9UwbBfykLVK6o+2nrVlFTP
XHljSKFxBlh1YpZxMJcUx3lz1u8a9bxQXZMqxsVcBBzBmPytIUHKWJq6CU54
okNs9PhgfzK3MREBMdjB+oX1Aayp+Sj6t4Z5U8sS/WUyp4uqS5xF+LLantws
vX79R5Vv0Ska4FnzFgqPVxYjtidyxhhDD2ex1tvyPpmu6dqhUWrdqliN6Ll2
CLwp5v9lYl5ELdFeY1PDhoZc1zNt92lbm8ZTeZryBFkAH3assuytydsc1HAZ
nbCDkVnxZ6leCu82luZaOIkib7gmb9LSOqFQ9C6wZzBLQhT1cBlhHT60zJcE
IzwyPnxhUHdk2jOQZWpWyVsTxUSYUDxiEt//Z1+GdiGG+btBto0/J+4Ny9nb
uyPrOnuL/z1AOdQ275R2IVNpDQ8qdL4n7HUDFbq1L5QcBeCm8vLn878FWXAE
4LBGqkGjS3wQz33xulMM1SyJY3q4nRsTSKD4kYCO3yzVXKKf7Kf0a6ZtY6G8
8pQB54WuK5djMFzhfxB4QYg7QI4UbXmCANPOknNWHpaMNM/hXenI5iEJuZMZ
Iztv2Vb3J7qo1wQBZKtCUzrQ1jf7ZYX9YSkzK2fGvfQ6T9uVQceblK3FjKra
q5h7r+u8TO3neabhUOzk4ktQAbZ2At9SujFEBCdNTQwZLmdsUvqp9/jiHBy9
A2chcH24jIr4SfT9d5FrWX/egu5gxsvUPdrVWyDLdnMVo/mjq0vB+AA2xD5Q
HV9lwIRNxBKfKxzExiASWtNHM7YxT8kwFZ/BRnizYTzCw6QgS3822PRTppyt
ei4BmPU+esdcWMuQXNDfQun+Ogi9vhHMxiZrzDIahf4kgLkEe8nSEtXfH0Wc
gdbu81WBg6vGyYaUQmHvqbXGpCnXUKIox6g/yQcjwfgCYmNZ3MDjHJ2I/Pjw
PuoFf8stTqIHHO//euTxACWflH/L4vwe3mIVZvlkYhbflqrh6u1FFbbTxm+i
kILTn+MTMgyaT2zNoTaNzjYX3oJo66iBEb6s40gJG63Lmhm9q+27On4BEWEl
xG7lxnFuo52DQZlR5LbR3wzpKQKJ4rghiwyFobdqDCnXvdOJ0/8vzEMvf51B
An4o6cTzWCJC9d931AyRZnFArfq35XSP8BEtOaI3ehtIH0lj5a/53XnNxqiU
aeWlmujU2re1edZE6v4Ho/RZfhmQuiKnnvaPHV1h4cHc3vcDb++oWpUQG6bC
IIffJNdyjxVj1Cjisn/VOaFfpm2A3JYqvuXGffrsgAqmAtTH/wiXMvYECGfP
bK9U2ysv01hWFf1ZEtJnhLnLZrZ3MyVu/nrU/Q7pM5no+q4uD2G4NL+Om9Qr
mj6iNGWhXulf5miwFyWXoecQ9iJy7V6v5qWcNXkSOWFhLHCwf4pk4MHOx2/x
N0VwOLNox7HouqEl/EDlL6+gS15JEZS1GOXq3E3Ys7NtJ/0+ZNigIt55NIRa
OU/q379Xm0or2pksmjeNFuuIlx3xmXDVoR4T9VKnx/ZSyErJbbMnmk4FwCrg
2YdSIgSUgLW7em3XPqbJqwvswLILZZy5fb/oAt5JEZkSwFkLsvEtsSR7KuGc
/qP58W7VzHl498q8mllrU5yYmLciVOGXskTnfuHntVEuL+w0Ebc4kp4NlMKC
reIQu+5QIxPipHhUpLJ/iexNW35ANEDDr66Kc8XinwGryOCIYtUcL78l7LB1
qFJufxVWQ2lQE3aTSUFTfyHL1i4tchulmtBKYeogiM3oFZq+udQnGAVXDCLg
pePiOUoMrpQpZBNoTcEWaXpHTV0Q/VkOmr0ujI98x8INlB4D6/WknW63vfqx
IvnBeGS5S4HxyGuP3cjI8HqmVHmtOq2GK1x0P+Yj4W2aIEgbwdteXVHV5HMT
tYxkK/4WuI4cj2NoppG9uYJ6kkXa8ZtiY9oEb/y4Ylkn5MFmxnARs+7z4RPf
xY63U+rgHXVxg+d28PA42JXq3Hhwx+sOB7gNNg/bwWOAzk3l4WXxAuizml/t
xe8n+Auf25GR7tFf8abk2+W6ysC3w9eQ6OHdjY2Mu3PBe5oprJVcpDLzPDHc
OwibVN/6X1bPEuVSV2OA23pSd1p6BEWxQu/p0aI3CsYeDvTs+hH/al2pA1Qt
CaVcRleAsZKkMahyrW+3gAu8R8Bs+iu1MjjGUb7Qtg1H3MCwIRg6zEGvldtT
SswG+Dvv279+0VwBln+HDeVTq0/C4fV2HCRF4QTs1cOGRgdiDHWFO9vXZAwc
kvwepvDLlAp7iZuWhSK2QA8WS69q3EqK77v5HvBRbckMx62mosIdEgQDYrJ3
8BUqPai4wxIh/I9vtJAZqTayCxmUkTlRutl88EnU0+++6/cczRusnSXT06zX
G8jITcjqtmNcRYLEAEczHWrF7Ynh3velpysvBPpG8Zjd5lcA+4s1AWhAxwCh
YM6NvAMBa7BEI6NCyW4F/kQSbcSLAto8hAxcs9mx8XZBhxTzSxHSsleH0Tyf
NfdJM8C52qLrDvfL9rTUAAs1g/pUUs5EsMh3W2F4RLjgdlg0Zp+LKiDvnmy7
UABrw7tigoojuBuuf7cJ4HMJ6EpK4xXkkyErPuAVdVavHdCY7yXnTXrF++0U
TbAWxoS+ilTv1eVmFlZ8KyZoRBR1xEqTdiXS70laWA6tQHFTmNihrBLvgwIj
8yW6Z2EGpnIFrutIJmaVPMpvfU900CGHVxe19CKU7t6J7pYDcTJ8Ug4hFy/K
CRVFope8vRs8n1+mu39FhNAtuMhVrYm/1HCqnfAx4OolIHz71n6jXZEIeLwr
CSmT8MQRObgpm18wijSZDwpJX4kykJviQi6xN4tPNfWe6tCBeRJQsSaGDBT3
G4dcL3ne27eztFIJMly+BdUUHiI7ooiKVrvSrXeV6hfIxsjTygXG3QsROKDp
W4DMZ1Zsk+LPqxoTKq7Ul/TZlpdzud2Fl1ak0YgvwFO4rS+IcbqtpDGCeMbT
ZnNeKk5k/QWwxNA5PSQQNszF9wrYMVMhXJPyM95iHzk2+KPcZGVidcz2+eVt
SfhYhAYfd/Nr9xpy9homgMe2Iz55zUPZJllNroF6CAg+1cWh1hxWm8woY6n/
tRL6eFX+Gl/C5n4mu/Kd5BeomCHoUo2IyJip2Yrgq02QkxX1roWzfzG4nQWO
StGxfHaU/CrBR1dPfgB63to7wtNirqPEYWQjUMJ1YZxFCFwOrKzxH6ZgD0QL
H+MbIhSwMdPaRzma+ZfyzcSdhhkdlrCAXJNyJ5tyYJ1m0UUi+8vJda+Epgnw
e2RvbqWUv5s5VewBt2KtyjfcR+QKGEpxP3VFPyNOzu+j7spQgl9r7yf1Xvgt
kZxwTNPzGlETTOMugXKHoIODu6No7uKIoVbPIgya5tqMd6qOR12+cM6J8u5f
+FEWlWUmMxD2RZjDXldReRWEoniXMlfHex6ZImsalbGL/8jp8ADiSElyAuGQ
YNFhJWh32d49dLRM+t3/fh/uN9eZHfkK/vraN86uQeg3kSm6FjLbfAcUG794
D5kyNtpclJ4IZ0TocNcdzmRFkI3mtDqr8tE9QEdOV3jkum+8HVdmGU3L/ggN
o+ZwphSC6uXeLXZE99MJWbO6Ixd2X3eD9Ec9OjCvKNeqwNvv0u+6StKQehpK
KFhMMciJkrmGv9+V/pm/DQV368SWIISspCoqiUK3cEzIEtTn4ratMZQTW0zZ
ZQUnWs+JWlNbZJHqG3h2zwn2JE12f/uM2OiF2aEZRN4RKorM2pTXJRmajAAx
6de3N9Ky/3Ffn7hBQ5LRV/A2hGlsfMi+S7LifdSauGlrfXz9JLM0kw61J+SE
BdBHh7bCirAd1vUXygk49RU4ycsArsfAGl6T8Hqe5XIcWBTkO/WP6AHFDCft
VZPYXYUnSb8Fr7jc9bld5BD5kvT7YMPytWIH7L3UJZKiRFAnwjX4m0LKxpW5
KbOFV4y6hqHZ+0hKMGkRQ5FTAkgcy5Wn+/jif/p/ltVb8YynjpKx9uZolWDl
CUCs44Z7GG++OHjTHOvOW2Aav42j9vSIdPxkH3UXHFcCU6nkpDX8ZTh0iEln
kRWauKNRKASdE7odtDUS2gMO8HuHW4oISrj1HQ33yPCTK7QlJXcfbAaDbyte
tGx680nzwCfH3RI4EhlEbLEJoyN6QQ2kMYwmmcYRP/mPIBvxUB2XMg9LK9vz
QFrbnQR7DGcLbG6HqR13LpjZ8rssP+lDkbSK4Fvrg2uE3iMhnuf5PZDT9X2l
svt5V5AG+M/ZR2cOWgEpxgSAvwS6mv9f5l8CoIR6DSPIGalDZCuoYT0Qzq3Z
0/1yCMcMdmdVJlmNk3qA5avhGhV4lHaRAvLq//56XBEqM+ktOPCZZPOrbI+j
dPKPFLMQnBFmh7UefXDSjamVGGCbf8gFzWi2JBDDaq81VXOWSCVRGaGME3r9
+erSEHaFEJ+gdc2XjU4binduDLT8qpx7O8Kg4arVPild9rLuDE886rkdTzqN
AzmGg4bIi192ikAX91gccI1UKjP68LdWCth7TnASpH2GQyGNNUPTcQTdzplU
OZoPckKBlmdKcLU/F6RJzr0IYJbInjFDet0N1pqL6nGnGd/9+/A5d1jNO/gq
hieflhFae8tNj726oS9Ul82PjrncTQ6sclQ+UfHLnWzOEEUqMzhYOAr0saai
6yol0V50pXQoO1BiB5aIN1MdFxJ0xxneJjy3lRu1Wnukjiv3ybTfN2nF26nL
cF4x8C08Plk24b/pLxx/lyXMR0kquii3PoEw2GBnrkmEVsCS23ITAiwji3zY
7TiMtbXsbrmfAH6uVHJzZm7yK8SGKr4XZCT4FDQjJZI81GrbsxaKTFx2EZYG
0IF7l98l3LzihbgRbRxcnH3XCnya+reWzU3KVhHP326HOM3DjsGkS314XyfI
rTDXlgaYBkBET39sYtaw+wUpmhvrGF3LZjp6gUk7s5cSQs7Vmrz3i6sfSJOk
OF76OFIOIcwF468Kqe+SBcWgxG3C0X9gMN205mlrSDhbMeMYr2SuzUOtorFk
eXBNi48tM+u3G8liaz8CyvVjP8JL6DZT/ZxDrQS1Z9SdowggpFc4WFcRps6n
hV404RV30nnu7wq8EPckw2QU9jXgXBJhJ51TvPFrwITuigqXi0PyYm+s/eWV
hr3M6ZEgtwLaPCQc4NL08aLLTWuJbvSEV9BfQ1ZE621XdOkDkgBNY68a7CED
noo1M7M3HccZrD5vom3r0nDw5HWughRkDJ0LO9jGwU1O84zEZT/rsA+ykFRE
9y3DVlq/FDJNEAsSy5o5A9EnfU9qqjguRKvaU9nhjAilWUhilJB1LestG/eM
lUxah/H7INAM1X6zjeW/ZyYldFrIkBoSdjg1ufXG0I6xcpIwAzk7dHRjl/z9
ERS0NpLOrImtjvJFtOdegzf+9Utd1L0ZUr7ucbdBETMrz+zla7YuplHhkRyV
UUvd9HBOP9UD8WlIU/WMi/yI/jKxymCpMpIQoBVbEAyL67C88s9Oh2l0/AOI
cotd+9XmJncyUYFbkh7W3b2VjMBM1cCjaRXMf3PsXGI5BhdievKf8s63joJ2
CmD59xR1iAsWkqme5NcNiodj/M1mjXLG8j+/6uHM9n8S1ZnCoR/UZEaS6n5g
qeTJrSsqX38aESpgajiHETd2UHUq79f0d7eMOHfu/4n67upHOisNTJwN3VAf
X944zjL2quuqqztNK8qaqwtkOqnYcywG/0md/03iONUA1krgQTVq/hdRhr9v
g/pe7VgZx5ASJqYVa5aJqkNXKcpEr2lkyGB6b771D8ZgAsOxT8Fm+sAc4V+c
1AgnQoxF2+pq2WXY0g0dBWXlgvrexx8xUShRw1AGo8h2x3k2ql1KrQLq+ShQ
jgydrvZIiMdoI3Cs3w/AtHd50tXOQ2+gjEbgJGIrHGK7Kd7MOES9Exhlgoa0
27Tob3p/xt0qTruYdNIII7UpEsHel/6njzs6xrx414Y/H2+LQFIrEFE+5lXf
8VirWUahQMo0ZgruXoZExF2ZalOZyXA7JQH3NdEPBBfoUmIW3tDD8MA2SGcu
cKDZQN6BB7apqsU4e2no6lWuR0Si8cVuHV7CVeCuC2zgVh/TnlzkKSqHbPAm
PaqJSqIw9viDin+jY016mDN2ru65+b1465EYD9ajsfgf1oDV/O6x2pfAqSoi
6ITTPCfB/ZlZBK/gVsUeR0TriHrZzMBrrPIKPVF/0uMcavjskqkNtVAxwxjv
dPT6EcnOU0ehcTmfCuKkRbAMrUxj89xbPeYiQ5kV/RrkG9V7/g9ErehA3V2t
EH50nunSPQsGXiIJldu+OZM2i6kKTU022nJD+jHory6H+dQrOHGupO/Q8/9D
fXulY8YNxuETV91BYh0i6641MX973hHFL2ptWdenuO76NX315bA+NqVxuRsZ
Mbw2QEQ29PY84Y2yJl+DQLNeAPznXZriTYY3J22GHxsED2wsNlASmP5MeRid
BBLOHhQ9UuDYpKNMS0iPFmXWFlPYab+2GO8O2sqCRjswAMcqn3q8jCvSvuoS
Zrmsr3OW2XTTRWYDL97ubmGGnfnxVI70Ey/gyMUwgXo2NEdPRMUj4BK08oFM
eku8x4NKxLe5Wat7n4brHjKim7CW0Lf6Cas2QsDIv0y7y9h8xfXk6CJ4SB/V
wSuJH64FKOK2oAvoQYFEUe7ysYt37T4HEFOQ5bpoy45Ggnf8J69ZLd0nUVRY
G0/5GixCmq8rx8BQoh9TgVBrBAeU8oOF7eEgbc9pl9Hpl9OpVaKrJS5SsE8V
dcVENtUB1mZ7MOBspPRPEVSPMDjAzIFNZ5Pbs278VkaiVNb4f9POohdNhIrQ
z1ZIONELQhRiVnN6bJ71vQGenHgj6iIgipJEItU4Hvl4kwv9pkpZLgtMNFAz
6r2o4RqDEwra+44ieJfc/Uba6cI/ZNw5GVEjueszqlQboIAHFBcHvqFhD0cW
Kv9PogRhBIV6wyBuZkJ1QR3koQb5hhCI04AX2JBciyfO08BlV1lRuPzF5pPk
x2mby5KPn11usFUW1f7nKWjY5p4gjpbCouvmdlUegekuTbwmBeMj85UzrnHd
P3GiYeOXo2TK85HwdqhVci2ohmsPh70QCanAdKUbcqmVuep+GaFIahjbj6wQ
SXLR+X5Dz22HrzyNwXhJO27VGSjZebGuieV+g1FNI5gRAgzUk3omCxXOA6RC
Gsmz0dHDwGSy3VGpPnb5YWe/vAY/xJkIE+1qpjVZO6ZmMBaqiYj+vEmkfdEZ
dFfI+04eDGyWei7k3A4uZslJ1sNzcb0oHdGXOT1JCy4JlUHrcXUkK8TuqRXs
o+l0L/bCFYsFvY7fRepwtYvXXe1o41lIkRmQIxgKONIG+5E+2MFmFxO5ptaE
FAP3+hYa6x+1QzkaFA/xgUkyOwmYFlcqKKf5kUpy6xawEIy3R7msedlMACvm
sJ3NarjlrNEq3wRlCyYQDXuP851Kb3RRp3daHCFN885W7EywVfKTU2Mr7Ary
x0Z0vJvYuyIJCJdEe+MkHkvew4w9uSPyFfXeLATVQ1gqHiQT8CCuQfifvIjK
C12xFXlFKNZb0AlxZn7IBYjieiot6eT4Hgmp51OHHnXsMEvBHmzVi74cq8H6
ChpajiaVRdpaZ+wqEmjhvjPC1/jWqYKcJLQ3AmZskrNHTzxE2HUMYayRJlpD
5gwQQ/Ne9fjO3qON2isi54sWqZDob1Ltgb0DYB/6v6AP9Kko4ain8LTPCuOU
pKMGScIpID/KXibZiUbQXpsz01x0ZS4YCL//0ffFZLOXNK5U7+HU19x7BTwD
wEDR5ZGlB3XSY9IwxdgKT2rRI09KhpW3ay2jAKyJFmOwt6svyypZF8rnOdgT
TRl3Z0dZjQ5yvOU+is37ee/OkaVl6JwsgitX8kluC1nV12MPIL6E/UoZZtL4
Ntwt6IwAqlyOb+c0rcZodRNzE86Z7UNvePpxtFjW8YmPwEWhJt3Edfihy2Mn
c9jewJH/lJleMBhDwCEWXIj9NVeNk9l6ejBLj4K0WKMAvs9+5iEQrQbpXoyj
vOQQqFyOj0oF412TaQKVFLNGRwofyTG5ptLH+DgLvHU+Iyrl0eCjTdhTcIRs
TDI0cFZAoqBsBB76ZAz6MfmzW8MoUiOflTBYEAkB2WJ2+4i0KtSXFz5z7CGS
duMFYCd4tbGQmtM7v+uTYfKbIYzIA8VbWvlWdk+wj4/4I5wp+R4kN+GUKaMR
TWl6JV3EukH6UfQvwU4f8jg7b7hP8zy+tOegM1jQ2njA927giojkNrKf/jcm
yJgrQlk+BWshzhzznBkXA8wMiqKjUutSs0Hc2ZJpeGZtHGIkn/D20t6Vw7Zk
9ie+ERctiKGJG0uaGnY597ObLbLRaHY3t+AGbpE3wk+Mh/n2prnFmA0kwe5e
XcU0dr8tEtF4THZyqQ0e7baBLrn9+i6Ld/Tw6kd72TgsitFSqJogFOP/F9sf
mm1qbkpP9ijh6pCR/CSvsyATiCmWNpLPhWj7NUgitRIDYFwkdbZXxGi92Nh1
U9UITVbsbfe8hIx9AMkZFbPPKp1FSaUAsFsQda1A0ikvw6iCvxZcox1GdTFP
/bXdqOdN3HIy5nUL/TE24UVkuI3SPrfDSvXPHc3DVorqLGqd0WAvqk4Ywirx
kykDgGo9K+FcbzK7iW1/zPoiHmjQmUJT7hISsowVpMnWKwWf+a8j04rP+b+e
hwfH6zGdUPqhi3NNOkxUS05mkCSBbjvh9LtJSFKnm7rbnYVggrhSQ7z7HhT5
l+pYGBIUiPWfQFHaCoGMqcAOx9AC4ofADxKjD/3wveqM0t5lRL/N5IT0dlHX
QERpWWYs852mR/ARYa0NUaDtbiCjGmHpx/wWlmQa6J4hzgc/tQx4wNTK474u
/1VLSRQ5RL6TLAeR4yQPIgn71/eQEP1imDl/RFLykQfErMMrEXZvVRtq9GbN
yyuOZk8Q0UkcZ+YX/6PziGBTtXJRESuyN6KnPLgX7xyY+yjUrCgaoaomTq7V
0o2UTtOxfJfi9ckloRP6F8339FxqKDEVtOVMsNanPyMByS3TsbBXdHvFQnwW
WU3eJ2EJWY1OluL5goUj5POUQ7iCED7KecAazsDP5m/kPYugz7+CQIJA9UP7
piVECSnq2dzZ6QPAz+tkRxVCH9zgrXw1E3Qj1V6iUhAmD5Qxw99j4hD8TVPd
fZ+MEJ9NQcQmYZJceDUEQAa12FFpUd/6D74SJa3PlzKIFjCtuM2buhKsS6dY
E6jqzWLLT13nMEHCnvK9PX6SzeTJU/+MbscTxObR+6+6U2fCopHCGuEeXxmj
bI5LRI6Jg3Eaq431Nye3qRsb0aNyyZCysnzdrvfc2Oq91nhCLCBHPXYpcwoO
3RNNjts3V7Yojqbs9+wj6la8Kaq1Edg8OAZE/E4GpZDfMzcRhGIgl+goRwlh
7HKHgJGJM+U4EaMyJ8GXuJ4H05N40EmSmneoXAMqTkSXbljPqC8+2CLoxQWz
isAeHRUkNFDuWYml7vduN14bx2Kn9tEFJEZ0s3Uw6xRWFuXo2/ks9PoiYwD2
SSx5DQ7eWmw1e4hHf33+tXKY3odbUmmeOCrBuaQoIv7fZTOd+3FUYpSRBWFH
1oJw7sVvK73IiQKY+YuOLyjGieFJMI8aU6HIy+Vugz+zV31eUnJZFbnSTr+2
yvVGfaBWLohpRoCihBtH9AXVKwS9X1Lq3lhFgWnCyFXa5I6RF0KzK/ri3cUW
roC0GAf1/TPkzuQo7qIqXWdRzJNKe2JLIGPuDSMsOS5FLHsvYzI6MaEGGDcW
lwaF0HFJ3xHfSJ7v6fWsyUCf9RAGK+d2uM+qVqtzsdKnW4qtXnPupZIjz+XS
4CulQpHUCOei7G+dNQOwXp27XjH6pVtb9Ml80WWM7j8iGMWH7IB7HbJjRlDD
22/fr9CTwcvTePzHpc4EaJV7Ia448PIqnEEAy3QAgFGq1w6UBZPZol/QKGsj
Eph+6zFTQpVahjSSpEavwdr7fZt4Z0DyTXGEHE3aeS+hCaMTwHQMk4LmATyJ
kYo1c/S5sp14A7YMtBVZdwIUj5GSC2Me+Eyu8Czm0w+PeMTzT5j3/DOJfgM8
NL5TDzwy9JrW/N9qiOR/UVgdAOe6S7oyQWXXG0I0WyXZgFOtbakTnOoMQklI
eHgZtAZVbleDMXlV7lo3q99FoIt23p1/wZX72861sK3fUJbNuWQi04XSySLv
XaTW10tIESqzxeVXsbtXZ7bxDULqonSapXYeDeLU+8Afuysc8gTmD47gdb9U
Xu2Vj12ioi0TVtSn6bjVxDkm64ZBlIj2CObCIztfhF2QWL4P3fUz7gc8AID5
Z/Qf2L7WNgT0Fy8QrVc46S+R6sAxOq50NB5bZTaWSIK3ccs2Mzi+WrtP9ucO
RJTdX+o2PaW5DabvFSjMH7Pq4zsUoVenr6hfBo//RS37T7vz6vkiXgvzozRM
AiUNgcFsPQb6u8bb4oEShDeVTWB8+5GzmK+GZJaAoQa8fq/nzpSn86agZ6u0
2jSg/h6MORlk9oKpJOiJFpBc7biChdv1rscA1p7zNYF7B36qhKhh3hlAtx95
0llkIr8sX+4SUTymWJC1fnn9hKxqpUWJ3r9v/kFwMBxxKh1QD5cbzh4wQlri
cATMy5+aUxL8L5M5Vv0+4tOl7wgexL+2vUpVlXp8bRDcq8Lk/iyUJwzQhE4Q
PajKZdbkp8JwqTWwv+R+YayYE4AZpyOQAqEn975Kj1Zs2Xed0I5jQEDtA4H1
TDqv4SNOXFPHkB63NHUwPN8zQG9IxtEAEDOuxITqeWU87Rnp/BJ6Rwfzyplh
iRNTJLUNpzM0XVZ0agTYV4ZYX3G2dmjCDU23OClXDsYEuCLwwh2tSmaOJZ/y
r8bcg9j4+FlsXb4vfCFxqIgIsm98rtN5j1wkI7oWGNNmShZoRNAHDvrFWeNb
tH6AO22cVhXMy2Tfolb+7QDJZ9ckpWoffYhZuc8BNf2vIbEKKsONcXNfQjwu
zb9MBZWIT5G23iYg4B3rq74PqLEpc2wXGZrP/OeTpF4E9bLQd+CniTYAczIU
CuOEZq/IYoNOrP7FcDUOha3gvaajXm7/7N2aJVQwE0u/Dg7lX/uJCqiuyweY
cQnivVk5a67/+UtyNrLtb6Oks19xkjabsmtgZq6qZ5/DvlRHJCvcwp5Jh6IE
7EatuhV19QU5qNpJ2QVmcK0BIrrT9ctoDnZFh0I0fhUEcGWI4qUty2m8CNWa
X8mYvnfavAGbm5hBK4q4/lCeaCquynMXxToCopmOupSGmKFQK0J8LGzuVbQU
Jg8P0tGSawUVVu8q+sPEM6NIRUkl5VOwxU/MsNDifRlxF9jqtSsxo0eVoJIv
PdG6HyTdeg9O28LKh2zSpOKPeYjOaM0NsaChoDaZC1b+PMcOlAZVHFZWAbrj
pA/8Gd3VmoVuBC8eZUXOHS0EW538cjblBCOyN7migGQpvHCYUDLPOL0OYn+H
kzkSwHOMu6IKFEo8BaC43RHbjbuZ6vMkiMOSQicpM5jMEOgCj9xEzcx8437c
Oxj1Jui9Mgp1vRzRxctGqgRPdDfSdxYTJC7i77mL9bYd+rSEgaMGPG5VYFaH
mg0Qa82nVcqla3opns9bUpHVf912DlW3weRizPSwYb8gnbPFXgeeiKQLvN2j
jBQyLxWHjSVtO053gxgosmHVWZJomysrKiEkSHlMltplfS13ZJjtylp9cnc7
oDxwJrsWDsZ7Qx8F3+NCpUFdNIcox2u7bu2TFjey6xXCdkZ+f1JjGl/sTImL
KBwYzmFwLtggJJtRRQSGK2vIYCZBkTRjcCJldv9gMrwceYCdbXsvp2SupJ4C
B1hQ9INp5Eyh9syb0tt5hki0CJ6avGYXlRBJeESepdvfo6vhw3nRSIwQHWGl
CqpaTIHQOvlpgdXmbLEzoeGG6fxrZ0ZzYLTs4su9yiEOK50WITjH0AJ596Vg
4fO+bbkQY62y0X0GNNqta5G3ycuVbYXTa6E07k6Ymt9BNFeV70EMB+Wg1Af1
7SES49wRBkl9GdtG+azxhTF5eGgho2YHsFFgNPF0bk5HF7ikJBp8uGICJJZi
9zkWfOkweY0zILslOPSrVITW5+3TGJJVD4CtZlTXawAu3pfApNaSdY9cxxU9
90wJ9d24CfUTYBv2wnSGqErfK6nJPbYKlOCdVsVnicHUsnfoNnzrGHo/uLHp
bxF/zAn3zTGfcd1vYraGKR4VCGQ3PRSMJiPo03GlX1OaENaEd73p3M1Zxtwq
oFBH6zKkYEXSX1YXJu0IXaMAwjfRGgXCa49AsCNHqUAQPHYvKFGkwDBq2drw
CB2XC1EgEU46C+QD6vP6VQ/iCpri0reLdMtTVcjNguA4io8P9tE2N28+2959
/NqPOnfImN6hTp7aKnCMhGOKq82jiX2w9LVW7TKx0YTbU2hpiuq+EioTR7XT
h5tSzVO9VfgK6PZw98Q/d+D/dDoLtWI+sjvlmxMJQ0/r+ecaYl1PMMladw5i
nQKyvZeDHuKZ4azLqRUDrWuAYEQhJ7gahf2lg01yJ8vBAX3TpVuvKb/9A1ri
6OtczdbiS/vYzRDirbx2aBDbE058HbzG97Bng5Nd+eLYuRfBIyT7kV4maH9u
rjOSWPgziYzJYYJksBHeIM59JemgyfTqkPzA2/2KUF/iqa5Zn38xhMta/XRF
uDEIuc1ZUT2QkCpY4Wh+sHqugRDIKCCiXVTK4rCGhhxSypS6cBVhoO3aOSN6
ktwZiU3+NcIYCon0oRVwh848tbKpwIEI1pCN3Ar5JZsq6T+RBvg6nuCOgqX1
+UoRU4Yqlh2A/eslQnHEzb3aBJWIc/8tS3dOOKB+fpunAYaFYjIJ+S+fj2bq
daRESxk5myIJV4YtIEWt2o/NkeNffqFP2IpmvO0k1bQT8+hP5bI+8iCoBzGf
rydpk/bJRwPZBU+2hYxldsoIxELLvXvFEAGLQL3chsVfDpK+dGVSYRVOvfMU
PQg7+dkAm9fdH5MR67dZdU+pnx4RgFwhLTY1uEdmHF+pXTqUjT/VmtXEyrIB
Zf25lUtwpcSu4NsQL51rqb8uaWXkjGqS3zKdewXoI8SK0NsfE7NvbmTh6mXt
8ZQDbdX5VfpsbqKgTSv1aIvjT0taSUbqYIVdNmK+zYvn5uEfVSjaXUDO6Ep/
Cr2vBtZbu9XZuWFMeC63hLTdJbINWh3ihiauW8QSruuMvsUGvP3BDkDORx/i
QJqcJXeBotKSvbpdhijRj2dYW0t0T0e/9OkBPjsI9ySctbWZI+FxTQ3YLZAb
Uu6cE/38OM70Hm0UL9Hz8rnNsXPGCQ+lbZQ/x/yv2tTz+1lJQiIsaIBca36q
csfk+ukrwo+7nEF2xqS120hSLmp4IIFB/4lG0/Ckd8QoKXw+G8X0UATsf1wu
YY4WUclNVMb+0WXiH4vuDTQ6bNfSmJz26DXpFerEhqIDhe1vyDZ1R9/yIqip
FYQLdSON4xj0Y4ovivCuk/oo8FvNE/SCEO9NK2aHTtIzjXwKnew4DZeU9mt1
JVw91EjxTkXu3aN7uGxz25lujJgThweU824TLMfL4skcwGyfJoz6mAEWicDG
SDiac0VznDbW386JkmIzdeZ2d7vco4//B59Akx7ZC0AA3jM01KmDbza7CJ/l
diW9s1gSMEAYW0kUOAimwNiBmf6ZmU3HzSjSHXb5RihJpyRdBL4LVCFrQ0QK
VZFH69nTIPVAXRzqlfBkgLNBBoVGST3K3ILbFrZLLThu9FggUzfAXojK5Vkz
r/zDO8sE/Qg9/N+jSaZQBphr56quL5Uj0Q8DV5yuobAXKq/fxPfroN9zq6UY
7DekPI0rvgvKE95uU7bZNYXwXdeHEcCYOuHpylXnC2ENcK9IsAngyS/XjFeZ
q0/HAM8n917sWpjVivnvit59ht3sxCltOAtWpEuiP/G39bxPhSBgy8MUeofO
GMlqbZ5iUgm9Em4tTbQTV5oirkNXlb44YiK2eYJ1dGQAc8Nhkwd3vZRH9jAj
X9Kd46TAIAz59/OS9dE+EI5s1zdgJqLJcmvJF4/3jgc6Y+tLmagIduZdjW9s
auWgudhkxTlH4QjB3O/7nluJxPpK+GKViQ3Tu6FJ9MZUu2DD6G0Dp2ofOtNm
sTdx+vCEAr7xAn7yTiJvJRr5ZlxN44M6aY2MtPl+IfPMgyvVqB5bNlGytbNY
dVdSbVHari0a4aE4upcqK5EXz7WM0urqT5LZQBhCLRGI+1RgZV1QD/ja7PtG
ENrD9xlIa0K4j8uOpLJO/W2jlCTy1bBIXaSNAhPYkuobp8mLwKUDVezrhMP4
m3xSd1Z5OrjLCVVxgJGASqMla8QFKgd246jZE9B2+9uDrmvaAprOtsIblZ67
dGwXL/KssYaGEhx4pX9IdoIp51qvK4PTfanyqfkEqEA9H1FUutXfqqiVXTm/
doCJZhdrN8WDi+8y9Qn0Rh2CtdSiXtWFHn/AX8yHWjUi43GhmnBq/xeI3E0Y
7R+5I1ohq2rmGc7qz12TOrgfijbS0BcMVj3+vELdvjz/aSg7p3PVZ4hfntXK
PXxZKb+HaNLmgqR93UK790JxM+r2gDwr98Izuf4Mf4fPqVv83YjTCdXGhdwY
y5/sx/OpOyJSqCNTBPaypWX0Q1pManrxIavWQGP7qFvzbDSI6/nf8a7rwRve
ebmr/9mR1ISqVPlC2fZckhcyc+VVPu9TBmB5+Vn18Nt5gLG+mc4ApW4TvDGF
/CWNx1DS9sA8qLul2F5koebKMaTQH0WGpLGgZE6z5U7L8eccHSpFuDUPtU6+
h3583F/bpJw3lgGYhoTJLigA2+iQIITRkuyuGSqKheJpLHI8T4mm8QSDULv0
wvIgU4u7MAcPle2YYc8Y27Vo+JPXBY4Fn5DqRqxt2Xr9Av32lFc1QVpaxJsY
neaJirvhTyXLOfQTj7Pf5L6IR/LDgWUdzx0n9enEG5pK7mEFQbZRePYip3gX
Q5grVsz2qUHW7gZz9PIxRj30LXLk4ebykr0Gjmm5qbYz2Ngfgdyp+TZCEawd
DCddEkR/Suj7YG2bydKim3fI9tb8H8/JoQ6cU+WWKEg67UBV98EHBTtdfH7b
xYT3iOC7nrpihQr03pp46xrhNHdw2mDOo6v/CFQEuElvm6Iusf9r3Oq4hvnL
/ZAy6nf49cBSBTwwUAT5VVNnIjlCqXvtMQ+wz82IVZBZRW4rVaiqxJ/giPJk
ODT4zwA+FRiRKkOnC+NkmWRx00tsXKo9QL7VmeZ6HR4m9FgE4ChZMWPcg/cK
s3C2aKEyHD2UVXAw5TCZktB5i2KefIRvQKHLO8XyjXyMIq4p200Dp2klMR9l
tcnJ80i9OlGjikr7dzg4fC0R85931hcCxv4bhQjmYw500iLtXJ8B2p32JYn+
nW1O0Xn46B9MjaAUp7midC4rchVIEdedrfzxGIDeSjfr0Qpdemd7FIDO7rmE
ws2uc7YK5C0oZm+ey7OkoEaqat2fchdHO/Hn49g4aHUntX3a348iUA2L4WDl
D6mMxJZ6iuKhI5+Y6GrTBx6EAI6FnudG2yQwP3U4Gx9Wc6DMDFvjATbHoU6D
RhghKLBFqpV3wMAkM2pBIQepePwgvMrsGKOSUx1wIl4FkDFMFXqbC7l1vOeX
Rj+wY0CpGfTLVNDin8lTg1AwunKA0lNXTPvABSsB9FXJBPZeJXckRc1d/osH
zRJUQdVkA77zRmuIj0u/P89D4EG/e0c81K0qQ4FSpuTVVhQeY/yCg/Y/sROi
6+dOpdEjjCmfsBKr6qwxnqc8yHC7o5K9fX5UOw/UnEh0SmfUDlClFzHx7jkq
8uFphZkXahO47Ny6SQy1QrYcxbiIeyc0LKsni9wUFywRek0TIUZLcRiHqG9n
dbRUgiEYHiJ5jDq9qarljt6rjP6u45tgR254mccfeSGipYg/h9OeiOZrcvv4
KLDpZlr++hrL0X5HtdInHWiwlCVdCdbmPClHghiOMNmVlVvgnnyLVTQimtzn
TXDGSP3lwz6YFlUnuklupJlf2n0sL9S3zr2EzmzJ6L6C1Dgt2wlmQoVekbbc
yuo6EM5bK28l/JD1JfLcFd1GeBN186/MBhaUYU6g1HIkUYYnVZ1LDS0o4Y5W
VLir740dM9ZPWve/qnAcOmSJ+B2Lybghq/njOhixi6XNJzZHz1IxkrCdYWBl
2ptiSV+rY+wqWswDaeAlnGOlDd4jGwj0J/+6LwiUGj/ruVFJiOEQ8gwV36wf
dcodrIgkRDKFJ6LtI61motVTomvI2BC6s5Vq0w3VvsqXUZWBK+4O83b2tBY7
nM90HVM++aqxZ3pLHAsWQwH/V+Pvk1zl00bNIJ5vHFqLvulMKKa0/ZErYF12
SZttqM2KlIFEvBJBcq35sEilNTnkb6JBnP74QNdG44Vvxz0jeYfFOYYmTHDJ
ud61OwUeeM16KvRFfbxhoJh+LRp1PIAqvycZGe7MGMZfPwXn9L/pc3n2DrdU
Jdc1W/d2d0IM969u17DeFQWMW3afBrM5sELvwBzJlW9tuaP5/GErIu/pBjtU
CUl67uFTFK1MZZH/Y+PSoJzF/TlZj6GUp8sCuB2tJQ3hEb2fCV4J/kortuV8
VZ108YYMO857ux3kdJbVwvmS5caqplBphY6XleFjL19PphJ1SCmOZAUNUCXl
OeFE7jKerqWSPKP2kN0YyFmn8OOmUcbndIuDl7wzS1Je+S92puHy8kOEuzAb
QeifvMX8Yrhe2YSNyhinfnRcuAxHIU9grSLLwWZLlRASHuJl0p7AIPusWygJ
TF5Zl4FI+Ua6V5cxpaVFBvUgyN+FSs1ZnxNuCSI0gpZaLeWlY6s1p0LpUQuc
EMva1pElmfZOtq88vGXy99Bk6Jm4lXTsxyi1nE11Gx3aUZG0Xg7RMW9Jf8s4
6DlNGgI5QXVPOucEpE/hZsR4c5FZc/CxEpwJneG2s1zRsVBBxtcv58zQ5FNG
oT1qUmVIaWvKDu2hYV1+sfNeeC37KPInCOcdrpUaIzbHATNUygk8aeKVq68o
Ka5rLGyaniKyj1l56oYCcwIOVfNVvx8+BaTSOgZfRMm5NWSyVVZJRLZK7F1B
c/js6bu5qedB6u6VeZtww4W7Kp2ifI0SKjVRbsy2qB/hore6azhmb4TgbOR1
hoYZS40oAv+DH1kd1Qx8UJTROGpneYlZ3PnFrjLqrORzMWQ1zKTn77gFwNct
V6NVLkeKa6gaNG0cPilBDhzH3Cb6GMZZbJEDCmqWpESDCwrVFYsR/QZBb2I5
0lL7Y50ojqQZlYyYw1Z93INZ30UZdUJI3unyi290U/nlXJP1baKyzPUmuZhs
SzGEYy3h+nk1a+yDsaNWpEnAMl6vHQ7DKlHlXNYzUubPGbo5bxeVl2Dn7/+X
K4JVeuPuSQslB1v3Px+XjROF/IaoW2MSi2i7FPQ4iZR2B2oxFDXg8pqCOMkx
jF8RhwvTU1Fk89idmMBX2au+o3MCRiIWSpmqX5OnfDY2b/tCJWf884m6cVIC
4HgUWm086IWfwgwSQcl0CGNU0Jc1jUK2XtjaIyAdsfK9vLENV9i1/d3SyazE
zYI9fuhLusFRynAkVVgCS6/yqDgsEKV9FYlygYieXOY2j+BkWg5EB0kXdcf1
2b+25hkIIomNDgzjKkD5G/TuMQGv2ZR0s8GDDv7WhNMKH/WSj7q154C8Smdj
aylUVo+j1XqsxD/8GBlEWbtMym+c9vKK0jwtvCyU0RaoNlhOUuQBlkYoBxRH
RSohwEqOrSOrlQ2nh66becPpqcDqeMIRGgd1Qh8jcAnhot9TNe6wAbQi2vot
e9508adZX5L3ORkK2459QzWYNpgRqXw6HFaLpHHmqedkrnGhbtxqHDyh0hJI
Nn67boEiyQIlb+bwtiVzZlMMbZxntmTcI+HAEWCxfuIX/mIqALlFWI4Lm+lx
oRzbOb0Z/O5sh1HqGl6cDBFK67vnyRwpkZrK+2zl0/OzYuDs1K1gsdjtlFOt
kvBGQHxtlufowBDf3gf5tFi+ecbdPrT3E4FHOBnE0hqUx5ytg9rnaM5zO7T/
+7TCg4oDsvbgFV3O7p7rt7YnqS2Kp4DcjZRTvWYr5mLDsxjHkqR+/GW3HCm2
azvL55ewacS47PH78ZOAV5QYFMrhkGdesRZRdhLh/Q/1atjc2Fwsx9UeG1SG
MoEXDJNqvKIx3as7o6ybZ0XPopbllzSE3lpgSTKHJvnRURWHkHd8Q/APK9ko
07n+cEnjiGLeN0PKKyMKTFjFrGGPzfpIq6W9RXpM+IKbBSQX6VCs2a3mn5oK
qzQgIE5Ab89pOX7Vo9LXwYFvs3FqDDHiHigB8eASZ8DexTT4UTe9H+OHU6YP
kDZO9BDfC1O7ehP2MNyScXEQ86fFmfaXU3W4E/a5wRioaEyUXkghRhdsKw1D
hO2k96ghCpSTKIijmrrB6Ej3SlWLvPScc+9iMQ/plWNJo7eDL4gYBZO5GbYG
6h4eBXWFX5xOZn6jD8us4fOktTno2vPTpA24Q9i8xqinrEENi9bJd9ry7YwT
ehO0PIP9m0KsBiOxSETA3CI79/yG1dI5NFYln8nmiv+l2AkDCm/Igt/5tRmS
TW1qZlRde11vCpcaVf/aCyZfgdO/ma+L5g3q6vwIPt2YBRu3Pf7uhUckjT9E
EGiWtVjIwG7o6NiVeBiv0h3Q8n10LcI8yH3bWELqyFkKw23SQnjNCHpPfW1C
gUmW0qHjpawubkJdnUsCbfHE6pdgutHRQpgesVA2db1VGW1ByDPDGa3Wv+ua
DavCxgfGg8Ol4QT35y7fsGcSNIRjT90JOoc2jWrXlOHlHWexO/tTwB+TQpjL
L8zqZzz8lvCo0mmbCr4F74yQv0MtXU/jCs2QTarfrJqb5MfyeBuWUTptKkJw
N0CeBFhfsszsw9BqDIln72ln5FLQ36pMMcW9f8sOBbcr97nHdziFSeBSIleZ
XZq7FwgtoRph1PwCm54oZ+4EkzXnasg+IC2LVP+GN52GXZfuiq2wYzO7UKM8
HXejCtVGnD6Rqo3TiUczXGL+itmXpL1X8bfNO/ffqUElZQMdUhmv/6ae4DcB
dUUANR4Temo9CsGv9v03KmskjCIDvaAbooXS1/VIscNaMl427f99jioahSwm
7AQMit1h52x7NAJ0MlreXMZ2qJBwHqZ6o5o3igQ+4LMrPU1TfHU9rXAIo6n6
ZOA4eKpbE8mUfB4mF30B4M5/hyKHpOru/stAaCFre5oODo8opDDoXneVIMOz
8lS3c1Ce66RqIMvKAMndBiZeHgJSLZlAsNsLc5C43oL77K7YorIZ9KrwvXzD
+V94HtSqyGwfg2rn53xe/8WUyiuMNEDsgZpEiLQ71ebmr+S62rSB/uYjXTBw
IXp4ck6ZfJAyCW59ZBZy1odOo3ZPKS8GW+RimDCI6NXljPVR5mQ7MBKmKwC9
Zq9BISkrS85PSTnP7b+FjmdP5FkuhvFndLaRMttxiOmaNkf4idqS8i1kG7Z4
uNl7j8pHUmFOnfyPwNZsduXYUBcwBKeZXJb3p7xu89raJ951NLWI3acOWN8c
7QgAVHEWmS1RCqq+Dp8yB3KNTbPOEYxOil6691jf4Je20KpNinRQYI6HvFUV
GeGfqR1hFpb510Fv1CvKi6q8tbpMN4E24Hxj08Qr7Q3/J5p3Lk2uZzoBiOwr
LWFYlW8sx/KafMAz4+Gt8CzqqYdWpO2agcj4ROmGZK15njrkKUamvqc6A2Hq
n8+od5PzaK6/IEXvphnhcF3WxD0RHaoDaXlwGuGS+gpVac8L42nymRSXEFQg
vfwbJELwLeaRg65ZJPwOeCHzZz52ASMHw3PoWEjsNfqQ6u5U0jl/iITtpEXL
36eoEaCVvp8qvkx+jn+sojaUlYlzzf34Y2yFrtNMFDb2tbONb0SffQLLs11L
z/4rHNtVjHiYhW77TvmhDmSZ2+J6EbjkZc+4Z2WJZ3X58NYkkdnezy+kzaV9
FafxuqQs4471nkr7aLCCD5yFi9yi4i/XpEX/mUEsybQx/zmJ+21GJMOJFGhZ
Yz9R3EEn7gM39OS09T3Ij2J9kdTisPLCMJqTZsqv8W7Hkg1x7f2g0TaZFrtX
1J5xaL+T/VxF7lyK/Wp/0vCXTQbk2mFnnEfjenBiiLshSjW54vp0g84SxsZw
p2o+jZu9rsHR+oMz8lxxcMvLJA7vgJMO88KqManO8PwyR7FosV/n+3/kI3vZ
/uZVCsEByfYFqMJZ7CEiNxRWKA0Q/v5Msmj3WK2Ka/FFJa/k3GJqm1NjXygT
VsklwlkXqICbJo+rPqUT53zJkuT40i5w6+FBbykc/4tKw5VcjapiCkcuBKrh
zlHn8NKlXhOopOX0I+Ur0z43dLUkCm8DOX4JhhDY6fe5WRWYqHmQsLSBz67P
Dm9yu95jazlyE56hVN1Ahiu2x7HRr1f8GAS7K20aCnwMXVtvZ9b0vpZ64Vwr
ITMTeHkq+z8P834H9Y+QkR9Qjbp/zLaeBJnaHZ5Gf5ASBlGhNb9Zu1DucVjH
MKOApGh6XwsJUE61FdKvOQ3OEPHLyO6fZIEAxitY+nkcv7M82sIw9DvR33Kf
pu9tAiS8wBHkW0wczjb5DK3GWE7xh09BRkOh4arSwJzdnUssc642EXz7Mi/l
6S/IY4G2sQZ6LVFZEjDkp9plnz1RjsX4R5d83mHpmFUFeyrbhBTrYxmzb8pn
U4QdNltck459x2x3gigW9c2N/sW4fROX3kCVG5NZgcML5hmLkbWf4wbiNPyD
zr9Qln/kwjG6PoDubLJCVoCoLjD4clbtMfKbjU40uNQPmrGf5d4YpUlsHoi+
uMDCNlME9gHVw0EytQOcaFJz5mCaz67n9ym9+xcoGqUDgse4lEdnC/DYk6U5
Dz9o1wxCIAbrxCS1KYUO1qgsYf9GephALnCTTQ83LjSEo/44led3yJpTxBU5
qf++OSHYbuwY7sKqbUjKGdXY1s9V3kJMCTsIYaS7E3GP/lJcOU8/XbGJgW06
sGGQKePOjlGEhEeG3elczzmcLQiPtEZqk7S6NA3FqIzpLRzhZtqhK9NCOI27
hvYb7+NDJd8RjgtOrvYurM0CmzyG9Dq46LT+TnxVEwjxI7KurwWtmDfDgjF4
f9PNgz0sDgHOb2RFpavjdzESLw+0h1XV6zwgMQOqOFACg9gEIZiC3+vtLDac
O7wHdgnKh8gdpsmTwOySLfH0DOgFuFh4+aBxjgSjdX6ldzblrVqlBYnS8ozm
YTi8faoWBK4U6VmtiUPFBv8rrmPoJwjkz5wIEk1X1VU5LQPYdAerUB9Pzob1
Akb36h2gcbm8GHHkzJLPbfGKl9DTt8kN3Z6rcBPUtCi/Zi7v4MelqrEEthUB
wFFdm6TFkm1xklk0MzBLMqu2rngN6Py1OcNiG0fu9vhZJM+7ZMidbAPJaHJL
dO4Q/HcicLd/G7PYT/4QhTtBHsS7b/eeovqA1gr9CUfve4irXXRkewRUnxZ2
WTwlQHYyyyNYtwaRJFO43/0SehSH5czFLpVQwnQRrJSIoUlGb8rQqpPOvWN9
BXqVlORElnS3FLQcWt8o/vg3b/GOp8T/6oORpbjVNf0Bmo6YjcxZAjhql3A/
VRGigfIzO3xq2nbiRLGn59XNJUoQ63XugA9VM2/Y61k8hiD8UH+eVkNnuecw
3k094JfIZyr4PC7g3HYkIc7N2K8GOsF02hrJg+ILNERO8TpRP5uA7XWHytWo
mTffYJQTTXyqPz6YzbgvUzNKL7nkRTCmslOJF5qPm6xZNO2CrPk3kVyEhKek
VAqYwIHludBE8RQ4Nt2tapYxbMklsCgHCssXJ+AZMmjMkfsP3pfmazKSkezs
XmYLfVOGPjmt/Jo5ujEmmoeFAQNQqMghgkYFZ8kdLif69uQnhZ/697PZI5T2
glx5RsW4b8Ftv9VTDPcp9SRxoG+IVUtYwLQjAmPCS4vDQ+WjnD06Vgju+FkK
RMpkBmlTVEsHe2m3KC2XsIxde9i9IKRrLA1PSw7F0x0Tbup5msM5xefnIH3N
bfghwoEOKGVQAZLGxIQ7TN0u2PDwjb/NNg75EWNNJUcpbV/lCiliVXnKOxUX
t6GcSMVDoooSnYj9oOVeRWf4cScLTOHc2bRsiJXjJ1mTFeOesSwuVzI3Ppdw
KOklzKD0ULTUvd8xhyDNqf4iJIWuGXDdGM27opwGKt0q0V75YRMvpFRWMpny
HVRwCaK37nt7w1sJN3ie4linJwt5eGxfb/Ee3LZupD9c0w6Ahk7L447UsuO9
2mzZtVFQyHheW52fwU94gKU1ntgIz9hlbTV4Pb8q/g9ElqDNGfLm2S2lrdZr
+KTr4kUNMegXfo6zzTFWiAK8tmBduhRlE/fWs2BEQAIS81RYjuQjP2+Fi3vc
ev9eYPwWXgSjqpdSTLmv5OF3EUpik4q4MK4G3U0d7BlCWl4LNrUjUKJTeuqG
Q83ZvfJpwCMfKmQ1++ZMW5Vpc7ec6u+pMnOWXgFoi1eE5xoIbBmjHaxcq0mU
4J7M9ei7wf4CvBBHQJnZtDMI+KcqVLC99R8tmDaMK/RHrcFuz1qwV05tNCGa
Sh6bTcWzs52lQ48edorkVQZaGExJrvWEj4ahQBNFWiBICLBNvZyPRfazt+p7
dxgQk1iI2pDjSCZ2hVn/Q70+GI7e7ekTjvPqkxsIUHbijm/P+dyI2VBLoPkq
5ckknZGHh1z12Wbc346yWqTsqlbalJQCqhi6Vcx29PxQbQHTdeg78dZTOslt
LtYkEg8uPtsX8HFgvX5CaQdXlNafdPnbtKP2eVlMeIhC3ykzE+Z5h/CBXmgB
b4Gi4uFfwakZiAHgbwczLNeeAHSNUK6bAJaBH/9+yCM01WUVGsPVFKrNidC4
KZNBGMd91CMueDvjU8N3TT5ShNGGP4rips6BcilUvB+chZVJ6xOiduR//hUp
vOEAbCVjlDoZtaeC6qf3T+DQpXeypmjlgqgjZBga/Drjl+7BK8qYiZru4Zzy
FJhYAHbOMuTx5Dm7qCkxOxPLLqlJ14fKnqsgMpxOkSAVdjj9M8XPvMmiBKJa
O3ODtib+kL1AtW3kV24ny8NwG3hd/ooitCDhtQgRoKwWAwzAtcw0+t3zAMLX
K+0jN1kSEko+lnDjMt82R3k0NlgC7fNfSi2VoPoaVdgi3vSRb/K07XZ8NZd8
FafuzFP6FtbZTgYxT+whRoMoTomu84wneHfIxTYfMhHD8jJShOU0OHBYGdIj
xOltMg1be+A2klL0Yvwn2Iq38nvHheqr3d8x480z33Fa8zI4ZsmO849t6lwa
XBd8HhqJqLkzQRZen3Yl+FcEKz1R1oRvrr9EszpO6RzNuJ4eXmC58LV/w/iB
5rEQZdh9JtqwqTj4tRLDOfdsA2O3wOp6A+iEQs+oUbcZ1D+oZU6IAYVrnwdT
/ToDCHvq9Gxg6krxHUnLVMlPsSbQ9aQEO+YCNdOMtw24Xn+2JffHl0tODpfZ
6LBvIPKQBt4+Qgcwi/TXQUPVp5VMcIyJcPjH0APnS+ptOd1nEUHn2N1s19af
zCb+se6SYZ0purFnWzyHiyxox5yL4OjInV5f1L1/C81w6vmCmeBL/6Aor/7v
78YUgMCKAP9If+m6SD++McKqoaBfAWZEIAhLFdgQ2fGjy6BRvooVT03qQ5V6
/915uAJt9wKnaeyGKGj6rJ93f1r18u/vDsiJZA333PFiQ/i3fEsFp5B2D8be
WKf6u//KxL/joM7AnX7IQxGuPjwB09v9VN3WyPe+68YbRrbQbfqEBYLJeeMc
vZSVA/emxzSawvXubLbIz5Ih/Ox2FiNsfHHrWnR+Dozr1yv4PWA1s00DwZHh
vvwn53HgByBZlNYW2gsCZBsX964UuiBEBDRwb5ILrr/ieRXMVfG5Mxrpms2T
xuXJFFYiR9bms43XtR8aHgyxymMUrUBOWrBqFxI7Ixz5eStTVqEeoQSpB7yu
VH4a+8woE5/MP/jzBWvHyBNVojzHWi+wQgfnqJarY2qwAIjI1js52JfDPydh
mpGN3IuThOGe06VlOWBoL5VufmD1MGpp1+OpaxK038HSiErfmuAZbgWIRkPl
x8KwaDgySp98g12sy9C9uWsWQpqwDvMX5nuvOqhplfvg1V+uE4QhPXzLAybi
8d+Pnmp9BLWah7flpDd/JSTarC/N5dfhifsF+FRcYlHPbnYlO1y2ixKrFF7x
0Y3S8sEbv1fdpBkUzVFNN/o2Fq/3Gsv/5eYh2G72Y3McWofuamHfL1jGQFwk
hn+qDTAV+P2FfoOOzPkoauGy2egZk5sV5kMx/rk0lCbt/STD0rPUP4GqnqG7
GmqBld2UG7aO60nvnibKWY4bIkFbrP4hVIeCA/tGRg/QWW80MEv59c2OTXM3
hr74x9ypSpmittIH8C2x5nxnuTStGj4DEwB6JpNhDJYUy/NHy8wb2gXCyjWZ
/qDPjIsGkuYPwLcvq0BS8JjGqJ8t51K+avRPwwrryu3FzWaaEMKkHtuL3EEt
y7555KnXphjHg8Q54koKg+pVgmMJsQFh1jjqppk6maj6Kzma+AlnWzx60AYG
y/dlc4BLoaHp9yY+K6jKn6mTuDReseUbfSob1N6a8sgUXz5ywMLY1hxJJfQc
Uc7Ze4pZyyxIAdKpxlk4kNdQ/e0+fUuax6+hauS9SJFJtt/X9xRaDFdhQmpv
Kx7kv1f/atTJFwxpVUYPIia4JqzUBn/ItEmyi+XRkS16Gf+oews7LhaGdVJW
88ooiiMYcbXp5t2RSAX+UPX6XWsvkv4YpvjExaMSciHeqPERlWO+ge7e7mBZ
SdPBegJ2q481LL1DyRrTtCZvyhtuq0uzLejQuPW9TylPH5L95qOccHpbryMp
bu4hfycMkXGjBubQmH3FmO4bCu1tzRAzK6KZ8piPb746mS/H9ofUafErisDL
ZK2AAPGH5DLJBdD8DMxkzT6lPAz12vPpwl52LcOZnhi65gb1MYQCfJd+WJuJ
xkjyqul55obsbvjqs7J5K3jq/poQomdjbvq8S4d+fuV0YzxJWQEohbk9lkLv
0BYaB1c8Rmkgps8F7Pm+JFA5sAqgvgNcw2CwqLW7zjKFhmPo31Swq3lx5CkS
oEJ/h1vhaHdoJwN+Eg3xp8lswcQd7Vrk8BFkS/lB2VChnG6s5e/wR0w/jOtT
viBMdMaPJ8HVOiosJckWcLnXeB5NpDVthhq38+7lJM2LmvVE9wkq9u2lpNIi
2Jb1M5BDLSOApmz4y6KoiaFZaSiYvK3xpClJjNmRa6quT94IhQyEXUc77gy+
lol0+51wLz6Y7kAxCgKDsDFDJIrXYWkCrbbvCaasN1YOosPXoI4bnNeSg8rW
qDjqQh2FYH7fX9GGSGG/IqQXk61vABr86PQONsvL+sJXgJCta3Sl5tzI0767
zYQPWx7mKHgzSjIslyBWfxjrUsI/MF70YZyq9XEhc3zAAETzuoXc4rwBZbKV
D4D2nsBn29Jmi6i9XZS/SRC2aC+gRAtd0tPoe79M28QmqJEXJMVG1bWjN5vg
4vJ+/iF6bW1Asdp0tFsFsdeSgGmAHBfAM3y9VlcpFxLcaj4aQUNmBNxdbNxM
VTYmi4VyMFKDe1mWc2r/H+eYHXLxmc0j5TCNqF0qlhFWxCO6a7jW3ZV9L91F
gGK3jWjUW7NmXJ4BQe2HymACWkIJUDQy2g4PBgkLUzd/qAa9wA2AvvWjaYHC
aivboJOROf1nFmNaJLl9SY6G073JLBdaruTpjJCbaWuZas4fi3LaNmBXFI9R
82GnAKDKBTF5GFROL2Iu89Kd2qT6hxlmWTWfdUXf8pwzAB9svepMLxC067vG
1rR+qfCHKpbJo6Zkq2V+0vRROiCaczLShfVGzg5jMJMXIVHTIxOBI48Ln9mJ
iPEEyYuA/uAjGPVHmkjSuy8e9PiexRBI/A8fxZAg4vm2SUgN1SAM/L2UjLwi
7WIZxAIssF4ydsHaiJWw5AU5CUNtIz9gKI+cR3gRCr5ls2svOCjZqJp5VDrQ
x9C6hP2K9B+I5i54Smao5hZUMwrqGEbv4i5bl+XJTqy2BKqOVtsEZBuxiIEv
c6Syb2aAouJmyIqI/PGiGchBZFSSggDNB5ZwTBCz26eUAtfULjIYZm00xEGW
IUabYXP3JAJZ3MNccQw4KU8KKLPOSB0KjzfXNze+Sf/hHjd2cNjpe5gOrxGn
LYJXjY79/ttZTbVMwSRyvLGsucD/D4ueEGJ7ngLimWKORZvp4z3RbW13LN5l
ZdWfyn9QXbHrVo27vUxsosjm/msP3eP3LXMOOlUoQOFM894YIR2pj0PS4nk5
3G8HXUYlarDwZn46Ru9nss4syXHXKtZ66JGsnKZcQ/XRuLhFRJ9rsYdwGHn6
S3GFnQgz2KyqoukGjfwgKMcwp8WIJ66BnnpU8YFNdQdOExPK3L6jfnEKp8SK
wJyfRKUhHXg/3o4fivrXngMXkVizGwBmv4tJiTebsgOrXNzYRv5L3zPZXwwd
ia9BODTDRf2yzxAr3HHI9rRG7jm0NUp+i7ID/+NsN6Hse0dVlT7ujO/p9Hq/
yK5HJLhGxk2o5SVtbrHIsiEXurf61+L5g4kGt46ozjBeHKgqSS9utAYrGoPz
gLOuFjGlPdTzvyvobFTN+v96z5pTQ/YkoJXqhfYoQ9bHQiqcGAcPRstf0q55
PAsoT78Ntjn1NjDhoZvhffabLwDhkKzKrDQfRO4gvQgTTZCy5RoquDwdHDdd
n6eYpFfSc7foyEWA+93ud9eEr/6Us2CF3PxmuvJaOzcpPsHuihiBqoCWG/Vf
ujMdBko17w2zyhEttyfFDwxPX51qQh+3uDb6hYQ0EYpqkRBVMJs7enQyScBd
YA+1AQKAJMkA0n5cb6zqadkgROVvvHdJnBZ/ROtnkggCAKpJNubtbYIYPKli
HBux9CtgLpHD34uEl/Neu62rDX6IeYOtzyuoLIuYmGVhbi+45lPv07TbwbXE
HS5roZ7tbXjndfoYF9Ln9u8Aco3t9m6uwyAtZvAnguK6mkWuUZ94PQCsqOM9
6cl7b22VGlvJLuVeE03Z3X3/hU9ZdeqPS4sAC9QXYrkTSvOMEZcJjDtF0A4H
S060IuyiYOUj66YgnZvg8RPfUPS73waDsOVO15NxKh9ExGUBd8STBTZEHwLD
LT1jhB7+U7EV2z35w0FW921jrxrGTMYOC3tiMRpuwk+RrTonxoJvj5kpL9Wg
TR+TjvVYsGtfYhx3Lm/nvS2wVHDXck6cos0XIInZ0L1cx2GWk0AwiJhltl+s
EHZ0YRk1co8HucXVfo1peaeS5KQ7Y+h/Okya3vGles/MrQnEGJkxpJZl1l0M
AWj6xVxtEB/W7SQ6TmSXevxV9PhkiIrB47dRcsnCoddARpPq5tndW0zDiJ3A
4ipvcoAtvThDww8wh1q0XfpqAC05gnWbfFG9F7BG9B+URAvBcOzdOCdfaICe
rRvIBNKDAkjqhO+BElhajyxU64CN9Fe5xLvFvTLX3FQw2NJckXSRc7JMh2OJ
p6dyINArUzJsc33EIb7XeCBnw6fspYt6mvQKAj7PLEhx0VAvldbWm7fStxe2
KMwCKDyJlToTFYfTfr8igOihfYjhM9tahiXkHSWIkRUovKBMuuvorBC0dfVS
b5mIKtLjd/0Ir5JfD1H5TWay5OXh4l2m3LLK9kk8waaY3di6Dg8ZX5IbVapu
eOPdynchhgAUt7ALFro5ASL9xsA4n8QY3hmw+zzdakdAk4LjSifA86jdXYGz
yn6zG+xmOS5mHc+7n8b0O1eTQH19I3GHnCp/0heCjuiUdS2b90SwZRp5+hLB
s+HmNRx7fGECAg7kritKH5deGhH3LJQLCHwX1acoZX+BlBHK1kFyISbOpOlr
BQCnrtkBEk5GnZzwP1hLeq5uVcemnXKtQlz/5TSk0HOb5XMzj66PmCe2URGK
fQBWyXqTic0lrNGiFXtR/k6pYJQonR0Iy7yV9wJgIiETbeJNKz6nVotZJcAA
+hRZEyYXCOu/z6EZ2/THHrwvDZbnuG0koLDpLJdjXgzMJKTU/Zaz7DPSSFye
IdzakksZaShxef8W59R3EsoIIzYCnhqSWkBUHe/Tvsdy1tQDH6x44+P9VWpj
CxM/+7VaqxCoBPuPLogV4k+EEpNXWIIz2BFmTfKCJfdlbwWc2x6v0gGMD00d
0CGgtROUQA1aZfnbtMMt0ajeuTROZPRZbBpqvTQ4S/iW6yUdRmGD4Ltk2Ax1
HsN6oMNMLTVfSRNUcMH6ub3TLgdUThfLvoDzTdpi/8+thO5iaxR1SPo+UQeu
29EfUy3Whn38WGZhe15Zi9BUTbo9Oij6Tozr+Q1GJNT0h1SYecgaR8gw8fiE
eYAjnImuzDefv7F/z6zOqecORz9ilr4Y9KTL1K+0iOu0ow4h8XCtpPIzsKOz
QHLJC6/4e5V1i+A4MJm5kVcdhWsrSV69EjWRkCCinLKAdV5W0Tr4DUF7Xmtw
Eef4CBc+/MNQFW/wQPnoI6Rr/ddhvXmfzEz6xuff7Xd79NMBKkD4w4pKvuMb
mTDSSpmrCMcs33Hf9kPbZI4qPHVbL7qpF97NrTO/K9HZZwktD6j96gHkgCoa
WwRBh4Xgi37bmNcEhlAIU4n7n3d5hAra4Ze8ZPaeg0FU1qj2/L06CFUfcbp8
v2rW6+zxwqkwFkPSowuNM6KqZ9r6FLsT2RrNHzpdMuE5GTZCakwjox9knS2k
R5qfuZrWVUte9y1WzTSdUkC5lVTK+qnby/TthnwlcStMEJ/aA4F9mgxeQchr
bfSERBq2BZs2Eh6LEwR6KJAHZLUbro6cu4fAE+mptZ+FvtrgeaZsH7pGlA0b
37s5pptFV8Fh1hlhV/rW4QYhjOHcWqOda6cAgrJrKvL+OFkI6S9NKNr4b3vG
HczHLHS753HCG8Zy6KqJj5YJYQxqSqAjszaViA8qtxzyfFUhLNwHkQRl7Lgk
zWX1odILhQZiCAekFiyjbdUwyyxaQWZ5Y96oEoQxbfTAep9TLrV0Kl4rZKFV
r4Cthws2EOAXaMic1aZ1BK26yK+qW25TdTEJ7p/bWfcvorVjFoYSNVTfgZvX
GiGt+yFSUwLwJqdZXuUbM4CmytmVdt1gSF9JxYxnH5Wk01Mv12+BL+3EhGUC
pt4aNgxdKY1xRqaXfNUAVEC4XNF/z52lpJTWmcwj9jqBA1WxG/kLDhaMx3Tl
M+q7MR/SKOmieav/b6g38QMYLakEOq5lvJBwgQL97TaYpKzGvv0MJvorgwBy
N/zv/gTXMI6SIT+S1rvBnbgTGaFYIBjbzrKkfbODa5noDhI5yOFerLl+u8dp
u3tPnSHF/I0FV5Hcedr6ypC/NfiFvy1sjmgnj8orkm5N9LeSH/2gBFCoJZeq
+PvUzlNa640laCXbWV/5/rFC5j1NyNv8qbJPHf8N5UEdoDqMrM7MkXM/yyoZ
EMyL6mMWCqYi5cfNFHB9aA60It6bPKHHFzlOTSE3GMAjeIrdDJdo8B0y7/rw
jR3I4z6LeLtLvi8DiDOptfhjzshE4YB0R26TbpCCF7FntFogltS60wMKGEcd
642qOvIcRihcMMO5LJChnv37cZWn7JnuR51DUkspLk8HmyqSQgL2bquWawjU
q84/RmhzOyfFLzOAU9gphV2hZwZqUOZciMEguD+F7WDRkFEQN3OXCoHjmPj7
Zo6vUXhwvgzWesrn+WHkRGpyUp7nEWmltxyPQg583jr8P72acgnenhSjURwJ
d1ZmhaRCdf5d9Yx6BlaQvT99jL86SbF95eRsWCcGMb3EsXU0wX89pEcsmQIq
v6wyjR32QzavCXsHs7lVDMcv+4I/68Ivjz6HIVAJhqe154rPfrZQVNF9tCy2
Qh9N5yppBfayBmi561PPZF1rRo1WU7iPZd62ew4WulIeENLp05CZtY2uBza4
mn38ARaCviVWHjajFRNp+S8J6NpSssK1Se7ocj3pFjwjLL3dWGONsiXkmi25
gtMZZG7ZGwpasp7DJEpfUo6LuYQx6+aIGsDnHmgAvfExO8tmnZ0dE0kISv+B
Sj2CNPjoOFfmX/kKsKHFssZbbwu6YROapjZv4gpbE+OMUOdnVpB8LQjXZuIJ
cbsqq0KuO9oaTrKxwlQhWdYT6WqK/sowb5KEJlBX45he7zGltoLYY/o7rMNk
Mef2eZisMSQoZKbB4p2AJPbIembNRg9kDRmMct4zKl6YYUV9emUi9XmMEY27
RF2fBcfXOejqlR3p9ze2nIBDDmkMZB5o6adgKgUL5l0NoFasB1V2+YWVtdE2
vhc83ek5r2P/ba+L9Xz0jaa7Jqm1vy1Fr7GfVA23eWTprqvXhhkyPCfldbDU
3YFDSTMWXget4TMl/j09Xm5QFe2KGTbPSJCjy0JPW3nLhRN1gYEoGUeruuH0
BMtyzfPry5+EgSPHv/8WNYKeN13ZhNP82oKQ4ckqkOYo9w6QD1ybjaIrC2dN
3EV77W9AhrXxev7NWmKNyaUatURKeaP3JWC8+qWr62tf0nVF8rMsob7LHlB0
wrWEaUPsmj/FBsI+B0EWz+y01Erq7dS8Qs7ya8rU8KSqfADYSvUGg4aGrTp1
svHWBhlPg4b4xRLvVxUnXHKHGNctPwfcEdodHG66qk4HoSY9NEnZHewdX7rW
bW5FvA/A2LeviO0mH92D5nqZnYYSiYDbdijaLcn3PM9Fwfzy/J6Zhw1Pac+R
cHIpll2o/YYN83GTyla4+cC0sZYINT2A+smCr5KexsdncRFWDoAOsKV+aQPf
wuI2w2pcVVBM/Vbzx2afZ+LiEX+XY8bBdTxJijqQPQ7W3JWTRjGnfJQF00+o
37f+TcvhKhJNFBQJM2GQz+boxY/wB7y88A5A8gX3HlCwaVfH6jLePpkYGKYv
VvLZU9xSuIqbHJiYRdL+Sxhb8jCltGDEiqq0XuOIh0FEdjQN2rh49F2eT9gx
3mpkxSUeushjQ7P1SCat+m8QYE6iXZHJH/frMRBUWdZbF6ZQwhIBWDCDm5fH
vqTkYO+5fg8rBM9n6ms6lqQQ6lSnnKxvKi5XOMTjnnzXh3TqihGEsQXc9KF9
ZKtv/iI3sdEGQAyuhXPTFMoQxFMPN77JsXUo4ZZX9KBnCgwu8VuX7WzdBbnl
ntezeK6xCPlszRm6hf2xX5x+hyRrBjzrUvE1PW8uWzs9Q4vHHH3GJeKU1ALp
mB6xW5WL785o3A1wdtuv6vn+YWEJBIe5i0XAZvsZCjON82iQPpBjiuHGZBVU
AAGnh0TUQY6fNotG2aORL8GeD9biLOi6HCdlS4b5+OOnoF12J8lcnJdiKyic
dzYszAUGa2qcQ/bzmYrDVx4WKCXZfTeVkooFHhU3hl8nDdkPY9WLKdzbknqg
7eKLeZKkbX5kJ66wlig6luA9eWQM0TbYWoJ5wsUHzb3XG6vOmIjbr5EIxOBm
3/Sqgidwi1FnkXFmtUN1o5CSK70Hwhg1N8NWrZto1zyZNE2SEX5qkUVF7CSN
j1hgh90sAmX/cmbOhskY7I/yu4q8d7Hw6blN8soJGGW89Mh1LbyBWJ2OVU7N
JOGuaebDeJCgwC/t3ZgyvUuV92I1ul7iV6QVKmt3YhATG8W4njHTmOJzx2ST
jLJklI0ZjgtLMTQlzwbdcUbZs7JraL4H6Mtqplh1p6Nv1NF3JTRRRugHA/hb
VsWy3Eznf2tYplfk+Xc1OvzQHOaZYWVB1FgOMQQa0zy5AGJFIHWXYYWhrddg
GlU4HSN+X3BO+hRuW0OiJeu5H5WKJ7wCjSwMAbC4MzTke71JMgAGLRFrRHtd
gNnwmDUmTu2a4IDntRy8kSEi0BsbBDT6FfVLz2VcqbPu4X3nYUX5aDdJPi7C
lp3JZB4yz+BHaVF8hiEsE/mv4hiJOqXYFaiyXJbh2apKme0pq9kTFEdOXCrF
91p91GQueSkJqNCeh4aZQ+4dhKtQ5HrFNx/wXTM0H8PH7+Dc5LiFiLyMM5Pi
WYyDwRe7q70n9rD8lJfe9EApZknwIp14fpGW+Hdi45z2YeYU78E1TwyPUgMD
NBTX8wkUuZDQu+FIIxRLIZjhqxWyqwcuXKe/w5NUp1mbQugBPuCxVyy2a3iY
TiYB0w+Kljpu2oC3ScO4N1L4lsBhNhCXrzl29D1quKHLoRZC78/VqSWTqb62
qRiC16WHqRWRUcUdhrfpoOS1p0cLhh0/WLX1i/4B5LlPl6sGl3jVo71P7KSf
FyvYllQPqZi3+YeUJGHRiav/9irqXhUBCwdgN+JGygDIHzE6pH9wNvDQkuXE
G3ANSQf/klbaCQXrq1BbLXC8FuqUMVqXAbCTcW6SxBS0zAKCotgI5P6mnK8e
mpHdiR6+INTHWMudp4ZD5RpXPYbbcqxTmb56X9RFWwq8st2nv+lwWDTjevgm
nZB+ppjUHSLkKIJFTA4kJJGytTCAb97iKgeXR+wXPvlJT7FQD6rtdR0zxxmm
Ea2KjbPIUCTHaCU2fw8S4MSscydRV7F3FsvWmoLpLsdRogLBAte2ySPbErHl
/04sv7GOVgFwaexwLiD8WMldEU75/v3lGv/+veMUC+iqzd9h6oFD7Fu5a2tj
m4pC/civ12zGwxl+xVaxzjVbT/hB9BkIpXF306qzvVc1Le1BppLSzLNt2G6u
fhFIqZGQf+OCnsNJsMDQxEjRfDUirPg5lSkq4h87gMPoJ2PpjJGLjsfFtmgA
5YDKv41S3XcWAzm40CWRLSvPXyXe7D5nKY3f/zfG9fwGqDVbQ+K/z3cF9FkM
ZvGJwHFFyO9GCBYmKub0uUSWQoDSG/p6skiHNDb38EMb5r/3wV45CdqCbZ2r
3z7/1LFKLQZMKnSjUWCu7j6PsWJEu/WdOuZoKUFT1E/v9X2lacX2lqvEcvy/
qah0TKowoZAsuwAmphb92VhsGkBblf2o5zp34TNKjL8gsHXjLtHp8uYFwRzp
L1sDt1YJXyZmo6lEG42SgzBhAJpMcnYSNirXWNic0QeM/I2g6uD7jWCqdD78
BV4MnpNaftnBjnacxCJjJsmOUdDK44FTGvi8gCEczdftgBszIy1FcvAKMqzr
oT84JPLLjXlmqm1WugzvwNbAkXyCY2gr1mfVWeQh7+XMerUuSV4MG0bBAlaw
+GC/MXUIWB2kUWSbEefdN02+0MNrJ1S8a7qnIIt6EuSwY+CXTmhNqDBsQEHS
GGoSrEhE+vTq+vvgQxI235SiChHR/ZvUjP+rHrqJGHJoLmc6MP7HjuX3T3N0
rJRIQJQqyJh59R2xDoylTUZyjqONOtj+vWdJCiQA7Tcn3RTMIIXdbqcj4sUy
XFS3IkAi5KkoHzg/S3HKXamFXdiHbodrWKRqBDrz7h7lWPpo4CoetZgCTve4
ykwzqoe1RrZdUTwcUR2f+5cIkfFVEYAcl79rXkKthPjIcuGvijj57I5MmQAr
oq2Mpy1+DU6Yh02JT0MDiZgXBzXpbw2PFTFmU1ksPt6xLo8DUowB7ny9bmMH
11eADgwPW02i6X9EZ4OWfNoI3zqUC4nVWDIkKwCArJ+r3osb9Z9VSCORBBRQ
79yOURtN0diXJYhnT5z5OmRevqi912DXWtRPdjoFz0jKrIl01cifbRhP53Jc
y7pWDQcDATX9GymHOxMkTfUuiZS7BZT7vkvJM7UCJcaqdhHcI9Ztnv9ECb9w
6rnmeA0Jg1fgAXD8HR4mVasraIGicuFVFEm2NU2vFFUMBm5zTZKL5zhzBvAB
+8ahsBdZh3xboPgLoZFfRCuajmIo+KaN9ka4JPXwGnbKxmWdAA8HFnxVDKEV
6SLgSVh0PhOgZK9iZOpVBFo1UJ9o++EKwCSf/s6ZP1BDXBHHptnl4MrHpkq1
wXTQL9BCmzG+VhlWU7q9E5UkoZQY1qXeNgaBxfsBxra8CnCzWgqdjBixO2yZ
nHyrYg7FNs3jHZ2ZHudGNqT1YQ1/V/C9+7jDjT2ziN/eKoSVTHFBOdFhr650
x0yT68fVqsXuYreyJnyKJZcButOFACRYiriaLVZPcOtX+RuaqMleF5DJPYd3
TbZhbz8mCeQeAG5z/c3AkIDNZU2AzgbT5nQISY54i0khruIrVaYZXJVR4jKP
6sCYrjBVCm0o/8gIcdg2Hu1N34v+kZbJqkuz/2AKXqWx2o/ce0mTAJKaeA0X
07nqi8S6YGQR0kSWXHoh+d4t0vqXmXt2uxTxe+FSY08fuO1iRkRLvqbTSvqn
dSFw/FiLgT8SGSTs1PMP+iRgp2MJukGmmWKKVifSRz4ZQ/6N/lk7Zt1qCOAI
ibZyzG1RHimxQkcVCkNNYTkIC6z0gXY/sMCBNp+9lC8s8cka59x3BV03kStj
+DwfDE0LMxkrsNcXdTCLEYLr9OG9co7Hp83sGHNjIauRSWEQvliIpFNhZxOd
n7GBiUXmF/Z7Vg94FnMWIfiykPmjQ4HhmTh4UJ7nHEqZh/Q4O+AW+GsielX5
djMk+aRYh3Nqblivb3a7YL7XpgodA427nzjLoyoEqAQ4D7j2Ija8q/rISm3f
UulevwafP8oyvDwxRfMqAydgmFQ6lCkonpDNEwbGW8htZ4XelQ9cwLJzG7B6
NBP3XqNsc4imisxhMTHzy9K3s5EWX0aNf0fV+TJZ8+E2xhY9NgIegErrscyp
45b6+OPg6cL+2y7Tuv6NPkvgH0yeJp69/zBV//mMqgMIqW8hfTRyP9Ls3Kfx
UWDSrdYebbdiSJleGf0L0ESUW7ZbJBdnhHJmWs0oDNYh9OVYNJ9eS+jxyzb9
j70FVmwf3yduhA3DzPKTCTVR26JIVhYhNg8Ow6nN/qTatK5yNiQIO9utOkZ7
Dsg6kgdu0g2lJ8uUL5v/3THUj24IbXf79GoJgD87PbW3p5vKlyEoN/hLT+RN
xNu6oSlMZwv6yCfx90kpsd50cvkZ84bUTU3h3DxQj8ciKbsiZwcRhwePlQqx
Vxeze48AsByWGRv8q4ixlbvR458EjiG4RVHX+lOOtOTJmhjxTBtiFk9JG+Oy
4wIWNFDsodUp2a368yYm52yabKjPEoWdiFw0+rPUk5ezkq3j/DbcU3sc5Zoi
4zwabvdpK3fosdLtImkHE0VVphfrtHAo97w6Ynqu2Txf9epUef5qvpNsTbgH
5ezDR84Ew2MseeFAcgJ4U9KZnREsHjXDZ1tAKIJXQamJv2OVSAKyu8VSdY50
D0WGVOVQRxwd+g35SbCrc2IKMjeS6OWjggHt/uAytgMBNFsoPSNp7D3G6pzR
blQnfzm96BsE1MJ84FHDistYt2FC4mYWbIRZu1w06srBNd2CKk9KelUSQqud
Nlr5TIX9TLJuEqrq0WMpjkDxf7quqUBUFNjHqURgbK/Z51PRu2suRj6TqokF
tWsH2HrjAXkr9gdhO6YIQIMda+IcoGf89YLVlydnP3ibAkQ7xFOj1tA+bo+K
r1WD2SiLsfJ/8s227Sks28EoJlkmlTlQwiMIJFmk6uQqSO1Z0umPJ1+dqMMA
m5nwSbL/EQi4TW4ihKQa43UwBTLrEsHwfHMF1O6q4/BTnN8xIv1/DXxWylCP
sFPjvitrSfuC9ArL7AJPKx+ez4ABlSlkuXBHmAHoXCqeNEnSoebn/XLHEZXR
xKpmGQkkcOCxTZMOlvFbd60hk8b7QOtztKnXIgcrgD5jAv5M23wqWQwg4d8m
7kUBxXkYySXggKwc6TziLef23Wnm0goWp8JFFq/IgRL1Cpa7SRJxu3rvOEGO
rZpW/VhwBPyY6SqaiVw1Db6je6PVcBRa902ng7oIWng0p2wMksD8TZtGsMJV
OfajeDRr9qoahv9qU07C1JW+ajyKkme45U+iKlnlvYKTXtUTGPaMg+dmFEA7
UwKIIdubYXiSrKWlP/F3YsdnfXaINjogfKGCy41haT3wLLIgegFZMRjS+YpM
DzJmTGW3yRIwETRFK5tZthnGk/DjBH6xaEliHDTKPuRYBgOdOrzZTo/iyWia
irDDwa7xrUdjqGkzIF1Uhw1r20xQcwMWfNMlTkScI0hRW1tPNlt0QL1ysPAD
TMW40Rc49j60va5V3wQqP4PWq8NAimfkLjSlW+FB/ZxKn4s0+e1fmNImcejQ
UwGGRKPhBvps/tz5S9WiDAze7ZBXI0NvY4nKeFtx7o29RsQKM4StMkBHq81X
7TEyLiLWrkX9krETWyYTibOwYbW3FDAj0aCeBFo1yaAbtJhHvz6yNO1vsnCT
K0Fuku5ni2oJmgRaCiR97CyZFRQiI+YGrEFLnUEK1h/qJkJBL1MbFjb/ZqWq
tlaV8FGVxla2zVER6Z4D4kmWzkos2C7IxFFmN6j1st7Jjc+BpuUFpexJ5yLC
bcoE2ioL17sC5whPMouwfx70A6ITbUAi5oHLNXTX75q0/x2tG3ojnYV5/uuR
CJvTc8P6ipLHrAX476yNOJgnsX++63KgDmv2XchN02E844rBoaTQzp8rBzeb
i4K9O2OgH7qkE0VV7J83ZkpkcQMzolZNr3WHKL6ydUwJnXvFyLJ2tzlBTTyq
YM9VHL8t+jmYa+83SMybDAcMxV9NXHYqGjIUbs2AdQKiRGdKspwMDasycBe/
RklGu+HAVHOpTg0FEijygZsqQ+bksvr9mQci1kLRIOMBnWgk90C+2ofO5Ot6
v56r+ZwiCo4Rj2Np7V8sDJ3Reau3hkA/NR6bqYkzSwarXqJvmga8yNdh7PD0
rCoBnNKkHQDcRo0woBbxhzoANMm5IKHfe0n+dnYIuVgJEGEbpfquqcEMM4Tx
w2OTRzduv+Y3BZnjaJa47ZMP3MWHQKn7y6XniWHVkrvHEt59N6gVbGYJSmLw
OXq1WM1b9340PiypL/pT2YyMUChNj6wfEDYah6tm2O7UrcppSM4ardT3vVdD
JHND2NkJ8ktEFLeP+r9Lob9Kg3YcUKdiVEh98Te+r7wVBIQFi0ZUyeHBzBnc
1FnTc3HAYbL2/wxsN+lmdB0wdbCWY6wdpemOf1ekx/Uk1OJWTRgreoyk6W0V
27FHgFNvfqOWF8y1DVW3OE7zYkPQ9JXP5zfpX6wYlnSNw9aAKL5HvIWJTreq
DMoNzExrMhQWGgQVFZku5tXlzNe+mSqfFXKbDrD3z5M4Y6ItAg/iZ7xevI0K
ZTU2rJHaHVLSGvpwnUdfptLUSGcQB02GicsSRkFXCoUISh28lLKSKouTDwHz
sgY9iA1JJ4ky5DdkVqpZnvPoV/mVe3ZIQ7D6OHPWm/pXO+EOMiWJBNXYFfdZ
E0qQZn8G7xbb/b3gl8nTLImOEcKwfPC4MYFCmJBnd7SRettc1je1ZhhI7a2b
i2pt/IXGUd/C8jAzeNo1XTZe41pLNEKM2Ogp6jdWzvgQkEHgBZuNhmTuRpoa
55qNcDgx4N9EybbOUxL+jJg2/ABKtkuBOXj3FeXVOxJkd89g/Rz+s81Oahc+
3kCrGh8btAzwUy5GjGmviaScvdozXbzspludZSnvC8XN/ycT9UCQ+QYtjtKg
7nMk0CaG+u6k0kCpcrWacesTe4Lm94hvrtzxZ/fjcDToQyGmXqWPU7fN1ygi
kuPbxcQBMCnEj4Lni4ElTQaksHnsALevR3gx/z1SFRoybrfHJDHeE7nYjOk8
Ztbo6HyILQtTpKjccgsKffRO57gbXQf5wFMsdkB7B/GA4VfpFdO3viaAY8yS
O4Nx0WxjAKvpMdurv5iBrMM97DLawa2CW6PGYHRMOWbFEFM1QxziuN7MOdpY
9/yA/r008d9FXUjFAlaNfDOqP7eazQeaCIs0EzNtXLrfvSt4fU1oAiFEWzRg
MC7zKav1Xa6LWkedrGxRR5U7jgSzv+lpKSCwcDMlSlUlUPZZtt6Hk5oaiJp0
XFWtp+Mt3HFUwC9UT9AY+Dk33IHPmFNzevwWj1EdVFowo4z9kAQrtwSz+Wll
NS3VPGKue9+vuxai91SDm3OmHY8K3meihHzU8yoGtaHXaNR8qKDEI91CxDsp
w40Yk/1uKGOZGpLTLZMdrs9WMWz/I7QofU861s234a3luUi86zat/8vjwngq
PkzGpDPValp7rxQX8JzuS0Fn2PNFt7dRkfH98POEcRMTd5j3tTCxdBp9qSfb
9zk2LJj32MvE+i3wAuPLlJs5OM/YpQJ1scnpNA7z05jy4peDT67Po5Svdq2X
3xyQksqN/8SGItcQDvPJauxA7oEnV4NWIVBwDNbauHhwEUnZurHv6cDqcbi0
Bc14K00zG3EvHOAb6Yv5NlIJl0P2ZqrfYXHujr2Eh095Go0WVkmsaB5WV8L5
23tlYdnxOJuQt4DZmq+WjeSY36cvuJHXjNFDqTrmzcDDZDsj+mB4oCnaygEF
DScfhDqGdhEcTZZWZcWjCkcli9qAuunVX26kz0Z9yvZm6jDnK+yMe9VKPPN9
rsxEZJp+39TyQAxUeF0mTmOrdqCifSvR446m6PxivtFo06Ko08TBey2bDc/S
8ZfitvOC6JRgExs5VduPatFYav9Wk2EyrmFTCNNuX4IemlfGepboRKNJjkIs
3YFFzSnwRPuIqrs9TPBWz7DpXmKtS//yEPTPKUvVMVVk4xP7DO5y6WbTQklK
AVpOoNKO5uJjYcCGXajsCyXpLkkOkRV2J28gie2EcPrxFuDT+xgKTFlsuHij
xoqZ0hDl8d2Un5x2jKmt/BC/vDfsuGSRTEP1Y4m6zNI/IyVuWfd4cT1JBBhi
E+qv+FweFmZHsghdA/A+v6qCdy+L26e+ad28fAslV31+30aRj9KHmrCQRnNR
5a0VPR4ESkhhaZKdyld+Nsj/voUVc7TnBif02s+MlytB/pQtkq4YyBbZjUFV
6WyYwuBhHXkOp47cJuVhP+pgab/d4oTby1D7cZa1azHg17EaFqo7QLC5YnX7
jAaV7jHpiIGZc8/togsRp8JOqDyLUC6vQ0TBVaYf318LyXbWdxBzgoSfoTb4
JrZb5TRlCFNLtB+7MpF7RB+qovNjgWZLedaLrV+ibxwB348S56shpYHuUdvY
T7lSNJkocJVG9HIFLLxGUDzBiJ/PtJi1z8GzN6Vot5+9fcZviFZn5McoPyZw
6PNtyJevUig1nFIxLsEWBNtyN7YugzWt9uDiI96cbC1Xo8JDUOE2C1IngDZD
UFwl1wMzVm/WZyppBtL7fVD8/2Q7Fc7mRXQ8IH9AMaTKkAQoBAPo0OKYwuk1
1Q75EBpXYZ0AB5lZO0PrAUe0d22Y2EKVsUFhByBbPJoBxrgKHi0+v/pt6UoN
kCMVtKm5Y6syRWi7YuxaDL/r6BGLnRt2Kkv3nSZdcv20lbtXz3NZa283Who0
SrpvqUKvYgQRLQxiaKG2p01o0bgnvPuFvIqItDxrNSiw4jYeE4KH1mSUdR69
KNcTlT4HVETYzw1IMjtsPJw9ycic2IutV9n5ysIFzF/d4uzqFK8IJU55ZUgO
b+A5dCqRje7U0vqnksl2xRdrfO+E4/fZwWp7F4JxZI8jlOYj+vW/UMN5jW+2
qTJbuyB4lr2f8WdzzwH97of2vYix68f3x0WSt2Xh0/lCCnzVoOfJ6uxethiA
G3c0XHHI0E4f7Lf+ng2RvVJLI4PAroxgrWNiL8PHeo0blWhxO631Ig/TNBzF
WgNuYY3hxUo5iH23x5KFDVm3oinuwVR/qDI6T7iX926CvMZ2UuR4v8JsSWkq
EzLh8ZQTAoEMppPL4LCUzW/pcCD/JE6rxQX4bflTruewpKlRzZnR+bT+jJ23
0suRxcq8WxNexoC5HpBE5uEehynstY8oKy6+Onk334J+f0rnSapP7aA41jwH
wkZ7LyHFIqKc1oO5lm2M2c1DrSNU8N5I2fWP7eD5cGsi9LluCsSKgT47aiAi
N0MrGs7sOGF/4no91IPxt89w1ceIhdOxpj7Qn87RUFYR7KzRazsXmflDdYO1
vcGg/9GwEBJ/Vyb0jP8IoD7Ylsr6f9ud3dzw7Cw4Z2K+saQj/5Go2wSVCzFH
DbZgJBLUqt43mfzfqsqccT1EW/LkYdY94knppL6t1wUiiL9ZC7GFHMRF8AmS
TkHmaVaJ8OTkWVX+aqGR3quB0BjI3v7XLOtjw/bchZFlLbx5WElHuyPCDGP4
2pXnHqjUQHsQC4VhvxKUAx0ywRC+UcHeW159vDAvLrAKIIER0Zwhs6hfiu/X
hct7Pya6By0j3KxMTYGyprAdzSF4P2RZi7N5rqWFcoPhenZIrJsaSeGVAZNt
pNZ6F3DnWaKPp4zCkVWNnz/qitebWyVMRj4tZnukYD8hrD26Mdhay9uqo37z
UGg0plb9O8K4i9OJxf+jhxEBDg3g2qOHPLA2wPMTVhOFJ8P0dGxb6lMPLGXp
K+jlVRBdPodZba+2aJbm/qjwgAM40Be/cpxyanZWpx9yBEQfxNwZ3rf3cCGv
aOLbqYktwi/5Qqh2nYjxloHreYuO4C/7a5518YKIhtlJ207zxV4dBbv6vwC8
fHs0NgGcONAdel73BQLTklEbwgngaW+F1uQNgF57srEVkQD6j+evrz8mIL53
86eMhtjpVM4CsSxGd1oycHH+5dzMi5dFajEFhyLOwLYOKi6TJ1zAJZVd9nvi
6sq2+GWPkaMRsP9gG2oN/ImVOHHeU8skjgvqQ3DfSItMFpRJppFZJO/ohojc
5Bk3CZg4BXg5WsvZZ9aLM6yySiCCTMTl2ruXxAPmGQEvYqEo9ZW6nieEe9wP
0ylhGHtG1RG52Eu5esVq3Lqn+4en8r8aZTLk8DeVAjOdccx/bOGQXExheG/L
IO27jhj7iYvJk5oFvC1s+Wziw1d+CTY/82Nm/FRbFL41zar/4GoeHkpWwwFc
FVqWfS26xmnIfCL9he2DnkiOH8AH8oybovwMEj8UoVNhF3DuWhS6MGmdP3so
CTMigZ+9hNhFQHuuvYZ3WqoXQVKzyiZQaV0a6Yzn6KzGwL0MMct/g0HV42zE
73o4kfdl8JkxgeSFaeabuzaT1tRMwkkq58YCUvYTBrB3+oF8Ff8h1tqpzPtc
ii06zScOqzaZ9TeUiDxkexM3cnM72enmuif+yq5w02A9djzk9TPdVmnp0G3Y
8zxoIcMdRHQBV2Fr/b3XsouSB0DDcwfhvKILyf9M1JaDwezXd4SxfO1PeO3K
RM+zhVFIiRnKc5ptQzIFIuKOQz9854h+tj4KfBwi+kYO7EwZzGDsryfUvdMG
WrlOp7SYLPzZuQ07bz8U1X6Acw9t2K5hJKm6pQVoGk0UL66vLO0+VqX+X7pV
kmKlUr2TE9zdUX7q3WN7u/3Xsdr6IrPsBn8xS6P5nLFqCjZLUcvqAYDCIfwD
D9KmQWMvCrPLLa+L502WrCA7AFAdYoaEfDukjbCCz82RT7OJ1+mtNFcSSqRc
d3YSpmbTCKx6LK4aSt9X8+fis/stXTc5CjIK+EBa7OVIccVvnjNmH5VnlTud
oe3t0VMb9HVifVcvXaFVL3krTQjlRwiNbLblCimeGiHapyMUNzISYj/CPSUv
JaA0v2CDfnVNFhEt30KZt7uh289g7Rdi14vDB39Igxn4z0F2WWMmLfAqLm8z
R2oHL240AQJSY9I+i9qdbbWOxxForkCNfTUmj/UxiiUnQSfmlytWUQTjtkQo
t8Tk7xkN/Hx1/hV2uh0s0Txx1bUhbNq9C6rt7Lssv4rqREqtU/aIi5B9TNlN
5IuAyjBnCIzGf2zObl6rueSVS+fyxemBTfsgbHtz3L+w8NeFv6UpTWhRI16v
/qnTXr15A2GoOKjfAa76GeTzT/wDt8axvf7qOXlgFhYIChbKKfwnyaYSI++7
xWR5ZIjiTVkI9WOlYgg52rPLfltIvjZ/CyNDoXrgbnoJwTpoExltVLokYfPN
NaCEeDb12y0TdsYGUBwdufW6Pzu4yT0ZDXVae5olaMeNLppOdWbIGqAE+97P
zJLoCidnr3HvG45T/Z7rvKdUBvCv4tk8l86x7otc9n3dRjEByZdkFNw842DG
twjtpDlP8FHDJm0M1sPxh7rpDJUBemp/4s28hgR1gKTQkd8DC5dMRvQZJLod
r+fhD3Gg5LHrddqb32rXt0ArEIhZCPt5PZDGB3Y1fhbk1bwBNuC6IYb0P2zT
0uqZuIh527hf+cbt8DZN3skZ12PWdvydDAnd1EjNbgYogIXT6SE1QfAXbeua
H+ks3inRErndWnZvJ7GCG697j2lOnugx6Ek7slDYwH2CdONFXo/mnUUsKLg/
hfdodLMeCt2wnwnkWsiOeUN5mdcPjL3+4f6ReRF12LHuUnlObDMpKX1Fp3AP
WTCSjuyi35KxqStq/LF0b7pSuYyS0drShJt9grVup/35xspe8M4ukd8s6nqi
qHvKxVxucaWSI+ysjvSVqiEAHTodKRT8BoN/Uj8KxoGvOHWANEWpCOEp5wNp
3zBhwFs8R2rnJy0I1KJYUiLd7uIH50dtjm0p0yGke/ptxyat35lYcGPHRJqh
Z6bhMn4EqoF2Ar8P/aaaZqOg3nyxrAVSN3GbeyQOy3rJO+y5geAXONGif8iM
JLFV41FcBTKk6nq9rkARodi14ui/LEc3be8SLhvUISOn4lb83ZaFlcQVqUdk
2hMgdCAfZxKPSI8fWpFLmT1oQFHI45Qc7gIx45W3hfp9mcsJJ3YJ1EjSWP+R
tU7PAixuyOUba/SWlaJkL0Vu3KTk/6uah2WWeY8dDlL2cB+yUKtyk2pCtoXp
2xg15+ERMyjHbQCQUewm5ynTjuxVr53TRVqvNlPggrv7vU6Hz1WXZ3fhx1Nu
9N2cLyiTlYoI66ZyFReZEJ1IINpqfE1pTR+4iSyfKQl7Caz+6uZm6fhhCpNc
Hw6n/APUiuuQSMIC+TPmi+JFencVLNTa7Y5hXeFAqziWXVA54nu1AldjcDNu
ChsU5scyxmDBEJ35varvvBt37C7L7GmCYfmMXqOjz6GkCYbj20Y4nb9+Jj9Y
oBaUbDdn+IPDTPyI+L0JT9TaGg8CDIvpmAwyiYAAJSwx4mjPOcXime6L0bXA
F5FVT6EUveqC1AapVno/JDalU69URAf84dcdGHUAGOjh3PnXUnP3vcC0sMxS
daR7kjsyBqU0k1O+HnjIv5QoR4zRZPSyBT2zWQH4AMNg/tp8qzi9jq5OAqn6
YXoVogcQDGQaKqNRh5AnPGIPwgzI1EL0P9+ZS9q+dT6+bIMsd+Maofy8j9Rk
30k/0BbJdmpZkeWbwazKjpVmFfvNv5GmFXrrCSNkQtBz21YntqNoTiaH9SzA
hpU8ODKpUeSmx7V0v10x53tZQcJSKdESRuUR59Ydhd9DxmgXmw7ttO/PODts
Th1FFVzURHqdq6HUwdbiruTEorTrsID0OoDXz/Qf+hAB2z3re4ZPf7JVageD
Uo/Ql9tjpCmYEB4p6QF+KrzP6FYfjuYbq4nti9QHzVP8V0Z14ziqsmR9DCE2
0EDqBnCZHCFTxlqNPYIe/sY+umhVOu1HVpVSyUKUAg0iOshsmRQCau1zu+j4
KvZgJd604F46/jx7cNH4+NB0O107HCHbzzJ+9QmAntqwluEm5kAzujP6JKAW
S2ntDc8QGk/kcP7FwU+HTk9FskXwWzuk80vvByioVx8eGl9B5OsdVLrO3XQs
RipQ4SB5r0ZTXO7cpzw3CpGMAf/BnZJ9pmHlcsARbETiEEBsOY0n8hqlldZY
Gxl6kQ6Zf0zTouDIZv3GHYIYrJTcpTHQlnXxI+RSvDHynn1ukRCR85+Ko+vJ
eizBYkMGUbpu6CWJYxIpHsN2L0ZQBWNiVVTb+/LaxZLCqJmvMYbUqVl7OZMN
PpUVo3F5XmGS8EdgYf180m1aLTN5EsK9OPvtnhsFOeE4tetPdO51R+iuzrub
8ZwTxv38WR0cgP/FLLARvDwNhJuCBefMyYvqQXOug/aNqEB05HZ8XM1ubf6j
6OabAMqu36lQGIEQ/+/gwtVkMRHa/nLAwoGsJcDAEU5Whes4/5zLYK6cQ9TM
3EZKJIgKlpqqvt4ZXHH954m2bZCbQKp5Wxo+Iddshp9ijrsgZMvVEktYfoUE
jAgJKiqbliCVpCaBdSy9o5fK51ct0HBdwRed8Lqhxv8xGv/dV+nx/MvZD8pE
tdR6CT3aqyhdMrOkzC/kBsfKeaCOkb14mYuiCTkl5O4iJ8uftHRQ8qkHgurJ
2HkHyVlC+b5Q9FsZNAXu/Yg4NswArVHzRWiBXP9y2W+powN/hJvIScIR5eCJ
UoMKfjv0y0NK59M8bE9aQ3OHYSjax6z1JWhQhJ27sBJCDDENEkPOaUg7sP2F
3wQLSmwp+X1lt3QoLLFvbImGfum7X/5SETyOuN9rPolzv7c9SuIamFwDtOAd
pnAfCv/7h8Knq9IpAYjCiXZPru0zXjmmFBX1MP3++T036KQkk+PpflMFykzb
TFEUiPJ1oVVXIEsIbeuASzHODbGcZOiIdsjSAy1fTPXQ15Tk8Zt8y7/8sZxI
vru6LsUtf7DVfXIhoWGMxnrVynnAUZd6drPVaMuNXNPNPBQBiwT2VqoouAR0
m4UPrr7Sxdr+G3zCYHU4ego4nZp7x2s9JJwiAg3XYQE5MbEYv3Xd9JUyNtlD
InXH3r0BRb3ZWyEFzuDtU74rYJRBq06c/6BkjK2Oyo2IunKrfcEO3t5awT+1
0lMsr9sBFwahpE0LGGxXJTNL150Juve9dIpNsG0EdqdSl6SCOQnPXBL4thf7
BOphaz85cZ4Hnt0H/+N1HrnCwiLGSDplmdM1rwydb/XELh48tHt9nYfn3P/u
MexZHFzNaLgqC+ifj4YyiLbEBSEAZY8mfwjSRiwe+q6RfF4AYZkKpNUsi2/E
PF0X+XU/OXVtGJvgPKOodwHPg4+IBBlHr/bS0KEPS0Kf31hjB8B4ovvpqn78
9/N2dLsgcM1BEovSTRd0WbPRvOjDnfLTiVE+U3AbkSnrKhOYpG2T0Kcpx15Q
1sN1JJ+jlAIPTP14vTLv0FqjFxZHv4kRiRxic4co8GXXl84k5X6d82EdWBrs
MpraEApqJErEr42fmAKmdd/NOCJeW+EYD/hPs2UKDOhES57Pv2PTk1JcLB+F
sNXOaKlJLOGjQzxTPaSMlmRlJP6R18/hHPPFNov34Bixo7Odqu9tRSANZ4/M
L3VBraPKHOvL2p690RAH8L6SITTa9xofXFbiOA9HdGzaYbaH1DtzQFs9CFgx
p4E6JjGKaPuNc9WZohGpfHRKaTx17z96iuRhr2F4oC4pOXFjMD9alJaz/2cr
gqeOS1Caeyx4TpSc9vRJEpHtI8zmHaVS22d0VrC3XZspMN/J8Fh4qworfsUj
/7176GHQ+vyHQgMtp/lpkLAa/P3pPt2/zgMP9p0f+X4VV9sW50WZ2wrkbh4p
kPfsNCkaiBO9DSEdsLTFnEtjWOtRLorQaDL2UY87TcvYSy+kbLF8DfqIYTHn
2VZTTx+xfdZJ81o2fBj9CvNtlspiRzQVcy/sCy5cx6Sp6LprqZNrcAhIu/Ky
x6prAKybVgUicPfRbuoKvficH8T4MG56MMaWkoiCQ9bw7zXjqxbc1TLYK/lK
wSxkU0936NPUC6A+t5rJ8BuIOgzOJp0B/95j9bgvjCQ/O/RNmlz8O9DnCWbJ
OlMuVcCEBMGBjuDjLFE+nXx0vgNa445+/Nmoj3QlGHhcmW/+Eqf0FrvTeoAm
DEVNMvyNvBzkUoW+6ay0PxuFw4vR8xXmITPz4nHkbOEVD/3jV9e8kdsbPNWl
k9KZJ8gZRLVyr2AmFVroLWzVC5nWf1LkKOFYRen+3dm9EV3GXffKf0TpbxBC
N5XVCHMHb2VULdNNs2Nxt/zeqEnv48Xqg4qAapI684j5KLdd3Bgp9F8ALSa4
jKHP1eVBm/HUhgoeArUMvqEZbcw4q89/Rpsc66ab0QD9Wx9zjxZPj/Y24jb+
9a7V/do2LukXO/spXLtSFCEh99j6FDANj1fkc9aJ5SQ97K4yRHM9wK1taoC1
5rIiIk0GVbJ0jzx7vVU+djt50+Gbn/liu8bIqAl1Qd7d8P+hxpEa+EBe0WNc
yR0VAz6PUprmM64ZV8IyUoxX5GqL7TGvAI5gpimtajdyTUx+uSEgE1r+YXb/
riC1QdOFf/ibRzT2clDDDxwTcKS0YNouFYuGh+3m/yCm8vKUkfQrOvegpER3
0zOkMTCC+ikbARd3vQZXyyekQ7+OnD+42LzftBvBXrT99Hb27fyws9kLL2h7
oFdSLfPgmDNW53e/G6+OLnwkpAB90XcJKlxMM4FpWEhdZWRWZzrB5DqyJHFT
CEnQ2WM+MuVkubeSgWmD23gfIY8ZU+k2FrF3qpOtWLD7MkIauqUhaeDYKZ1O
b/XKYrnpzgoijResLfZYmWQFCNTmUjavIVYI/dVlDLaAlqUYZIrqBl25Ih3G
VyZG+7KLVuU4mkUKrJlBl5jP2dVaCfZvPI0VLycwJXCvKO9Ak56SLcuEBrLc
2uQvjHy0+o9a2XpN34CBOMczdjh78FCbCfJQVDRxjqhlXCxMsDKY1JBnd+dE
1oZrJIgLVkEUOXXjF+toCgADt99FIc8dahAJUkQLanP0d6XXeVhvrgPA1d2H
7rh+g88ErLCUqI1HTrAs/ycclm7lpDkTuBZkt4ChTx7tnJMKGOpz9n9nENVM
TUh8nosbZtgaSp5Q5FNjqKHwHEbpAY1Wiu3P1OvorNNATiMVEY4pgBO59Tmc
+i6rYzUVgTDr6avus0VdkaYnFk1pyp3S0uFPagOupa5d63vXyjL7ooe4r/La
z2lv8YtnJ20ZtPzXpODQjvkNPvWno4KKxiNElp0Hxuo3wrsubmI17EmS25rm
O0KS8ZvrERHep5Ye4i8w6hoqsNqWOrx0gel/B3/qt+le96gCoX1ROM02qsB+
KDk6Kp3LJgU5mPoiOcljt/kg3xvhFTnhcV+e9D9xZJC/X9k6N4OwnP6knC45
t997E4XR3oE9fe0VE8ETq8kTM7PUNlUBWK3YnyZbLVkaDvYGVcfTnkVhZucG
VDy3VdA+RT+N21qIcl5qOirRudVJogqeUBhfOcNJXt0aXK7G1jETmlLUXfET
zI1mDqYNJjj7KctfZE/q0gXoSkAsti9qO8MfP1cZPpXogMb1183cIomDsF75
uO17IUZgPRcuK94GMntVM9Fiwb2RQd5rP4mQcX6BxatMH1Hoii1160qlXk8w
HerT8I9m6amQkrzXmPptnumJ6R8aJ/btdPJ5CmALaO2xVA8iYizt+bzDf+2H
TFr5tv9q1rEB4t2qFc70aFoUYcjNFl9a8ep1fco2q53RT+mP9puFFjXT8z7x
/sz1mTQ9GKGr8wRAS3JHWiP7HSynGoblTWlQkNZNhUWWN1OqhyMaLid4UqiB
aM+nF1wjZtTVmT4PXoyzm8RMk9Q4wNWldJ2kDOo8iN4CBICBsUdgal/+3AC+
BA3Bz5zV4WSOAyjSIjGRihJk4Yuqqpe6ZT0F9KJabtsOaM5fQrq9pNPVg+65
QNdYldBq93D9YnsPlLLWlfjnu+Z66czRM5Q//8dILeFYbwHKNvZZNRotymzd
jrwipHwwbPwHrJyd2wrF2MONZEhqL29Jwwl6583uQkj1aOx+SYACD+aRCUgR
3ixxJ6pon6yOk220FapWZ94zE+9sRj5XlKmlEJqWFXM/zeu7epKgMpENMow9
Wxj11b0yeS8U2df7/52dKtOxDJKYiUoxcMcH6UdWuGHbcrkLsGW2ZBX7ls80
+qUlIBkLAAgsTd30UpBBM7axlah64a2YvkSuVgYGiIxwCTUtdKvEQV9RObp5
N/luvV/UZug3F79M7ROJG1ut1Y0ny2kUQeEoEmeO/QyS775CA/Wbu12vUB+1
tk5jyAtx2DY1msnG907Nyhg5buyJ0udX2LUukmPf71aD/GpCEY1euoDYprdT
pJxe2+Iqsy3BhXQGJayfbh2evBW670fgRu75+AszX8Q3UIAI2Bl+5/xHFAqQ
UKg6bW9up+v9qclAdN5IuK5LHBpVEnzMXCGrdIrymvZtTuBbSMgQvGDb91Vw
ybwl2kwC9VS50vezex+s4ruGs9P5v/j6jhGybp/o8acNd0kOIu1lP6sGqNvf
/IsMIIBv9WshwkLOaiBXNRQLpUs+ESobmL1/FqXuK3JR35cFrU16rFIv2o1d
t6g3PjXspriFW1hJYYPl4GImI6weR8SlscNqoV0xj9G6kNEKtvAwNlD6Vjka
b9etyocxMhgtYVwruweTmWzoux19nJ3M01A0SOs013uScU+nO+yg/eeq1u/P
Sjzf4SLJVi3Xy6NdgT6ln9llVE2MqcJdFaSchLCxlgjR01jJpOtkwuingpgP
2LBh/2LiVKLjGXPLM0y+szSttozshQX0Py6JYmlUlTt9PrI/VbS3nkX+sN7d
aC2a+hOApIk5Vff+2S10saCoCNSZOEjaL0mq2/e7017jRKI868WV+NVQ5iWc
auHK+vv3tWt4mBWV8lw6YRRDza7/8eqJTcC1filLU/qX5pz1fNz4wXWOqLbp
Vl/iqywv1TAhT1p9vgS7td8D/Mt2x2Cehl/JhCIG4lC5lPxGACsvAnSiAT6c
ChreNZu7/PyA/5726knADhBagOoxa7QOjE8iHI28PJp1R2j+UB59GKx+TcV9
90FBjUB/h3kkWcNhyF2zGLgsCSDmHSQ3pE81XysXz7JiDqSPYH/JgpvJgGb3
v4SzKMJySelBeFvU2L8PofoTGcZAaf10JwToON8zeeW+wDxkTjAasalARc8K
bp6JFejBhTOpaNzIcoSChfdQoU+GFaPZ+WAJo+vIw6EM3Y8jqe85jrTUfC5c
VOay72+03PWZyn1i2W1IwP9N96O3kGA2I/J7suKSyMqTNRzIDQTDYjrLqu6w
r8Mh/sGiAhX3/PIqhhX1ZPFTwrzBWUdFQBfO1378vDA7k9Q0GnC37eV8yqwB
42IY+QeIL7NE1/wkb/tTzYaXFWcaMW/D2/nxPS3yTpibyUK3pcoJYIHanlzA
Av9AzFOedyeF5rlvBIAOb/q7ZV+tz9192xcuSY556MJ0mfJH0mCUlwe7Eizp
iPSIoQAnpxvBG1ue3LUQdcwoSfseXF1IG7ww5P5xdpA9O1X2OXwfsGCsGeBO
4iCFfO81TUfwtNr4iY0rR+nZ3OQc5t5vNaYZhU6qfm6F2tybo5MUORbMjSBj
t0yNecp6wUbfeiq3jYLeHS5Q5WAX/JeP0EYOekzI3W4IUQxn5yNLyvYsacz8
SUS2pvRXlFLPuovWgYidCTBPuc4/QPq91EgmJDIamaVb6O0uW9WO0k6Lkm0X
XuQnWsGt2/0mropo7I3pJH5rj6DqEPeyK1bkziCGN5hyrL7JvFkGCPoUlOcg
GHo6zPtiJo7Xb9g5DLmvnuJwjIA0Eof0IQ8KfsaL9NT9qSjYCjmMFQeu59dE
qZHb5eDCnrUbp95feqkF47ZoF1iHSY20xs36X4xWpkLof+zDf+rmcBe1RdO9
H0nQmHVf4Ks9ya8P9cwU3Z6kvfLJXcyy1AR2Jwu6NakJLcpoknbQggNPCKLv
piZvSp8T9puFNCBCk7nMO3zDA6keiqToPECyzTZ/BuMoqX+cBjxzFBxyEjDI
mXVMdKJ8q6Va0Oy9ziZhaic4XibPrtKU/LKrOK0Krt7qj2832djfm5vFjmmx
uy9sLuvckJ0caHaQJTtYbPjIh0dRqlGwt9LlMLRXjys3mPl0wxMgw5zMY7sS
GUMHJEr+238XReu3wJIoFbD6nIhbBbHXU4Ev26g0sXIqHwJKihdZv6eJuy7N
9BQOfWjD/9EGmz20u+f1mOPrYRORy9w3D/Qcso48tcnaQTTrWT3BtTu5b1f3
IGG7ZUekXl5qqO7PqHbn2VcEkWk50rL59/Gj5OVrMmXNSkbRdBA44ilau5Y/
/PxparaBS0sOM0Rnolcxl8t8P2WEgJ+wDXIRUq9R6gGCpqcsRPD8Retz4sI6
qaqoKHcgB/OpE78WNBzkmA3vzodwMUzkvc9aW1GBF1AM6yz3I3EEPKBMJTar
werKqSNloZ1oweeP7mdDUXfH7C5zNP7/8Ts0fN3LPU+oG/nCsvx028iZbykW
lYXRLkCEcgMHaRJ8zmB8aLsrc3rf9bOw4yuP2eCyGfdpGCwNyf/ceqapMA4k
fPpNgNu5rQ+IkOGaXzz5eVDtvGJztRuo8ouNMpSvNFpvBYapDUJxuZYD8GNw
T/P1afkTrERBeWGtaOmwhMyb2NXdFjICKK30xqc8/C7EeDtoG8ORw4Zrbz/1
+mq6wya3kHaB/WiShwfpKXG/X5QGxnZlbAUDh6L4Eb1tCxwroSSC2+i7tQPc
5r12f7tC4AgJZLnQCs6PLNZuh0oqyA8Uutu4ZhMSgsgalkdeoAxfyA8JfmrY
TVOIT7kn8DXST0wrkAJuUKNdjDXSzSWnpBOM596Zbv9tybnFBNDvhBXqMLmZ
CJnSKVWcwunzEg20/XHHJ53r5h04LU5UzL8MC3BRRvwmq6pJ5RNxEKFFVPCE
wEZMl2XgPBdQeZFhW+4wdoCUvB/+xGa6lG17c1QAPiLCpaiknPUjw04o+9BQ
xotbu++akdgTRz0XFwtPAlXvrv51BC3K1FyWW8MwHG1TRnTyIAzO1ey/X/8f
WQyVlA5/uGTrzLhRMj4Lgmp6QWiKC0vCq5XOGqXsJFexpwWt5sXzGzH+RX8N
bebsD/gSDDdMpq/sdZO2pMwQ3Sz/fNTuqnjzUCThaDvbI3vjMzDDiu7l1wUq
v1QDkzvmRdLRM36aR5zxgzDAFjokS00BvZJ8Tt318iBor09K0g2K+zpOrf+y
aA32eJIen5oNQ9+q/9S8UhKs366rpgMZGGZMPnUx/yJJlj+98JQVFcNDVu24
ZZJH2zCtyQcEJRxNJciCIAd2asVcmkngBU9cMexCoUfbgXpcOnVGm/m9OFKR
3x2S9Zg+Rp/Hu0zp9BdJ4Hxbe7H7LjDVb2qHDuZS62ahH1XBJseOMdSDryVM
uL35103Ai1mulW1xEuT+xAphcobhR5sGURXNjJR01/q1eGCtCIWG9kWi7wq/
WB3zSTyaCh77LJdUNge/peHqbPEY+uJ5Y+SNR7hfktIC4Jw4t7k6C5V4Xc4c
/4VztZgJeAtLp9GeAUfH7xFxULluxyH45gZz/WUKSLa12zlWTWwVxJ4t2xJm
HMOT154IaOVk0PVPDoH5lnQza6oJn1VNAK3BoajJhheD7fLrSxEi+oWbEoZl
re0HWUvkM3XPEgPwO3vzP9WxJHORif84GyNAUuzccWcYsxCQZlnSyEugH4Mq
QuPj8tw/cjGMHALNrbQXzfhO7wrZesejwOItj8R26UV+G5jXMd0xPziEby/m
3sz61dSx9wSrMYkOooA9za1W32XOKeMLz+/j4IKRAiezjo43LOvfoE1jpPVs
LFnrm1gPTeR0fGMWVApIzUQYZ/NE2BQjl6M2bFSh5T6bP/yTU2uz7wao61cP
OPtjMz8eeQGgdopzAbkU8wkF7NlBi6dFU8jzzBt9wn4KlYbJmJat82IRsCKT
sQO4W7E2PCRO9E+oa1uJWltnswAaVNR/LQtyZI3NYhaZqH4SkzncaP+bQZaD
8+dP1RhWgmfSXI9AZnSqIQyFOCnJQr0+O8YoGUl6mtcmd9lSMwTiMvb0wdxN
3EgGKiQmp5rj/it8jrlpV5aVBN8k3p0fKIEMXiOSfe7XF2gqTh7h9tgyQjBv
4y3MUr9Vwi6f0jqQlWLcJCE3Uy7FBXhF0MPPs6w1PuuWm0h9AcE3+K5UwOvz
XJlDcJFbMmeuZV6RD/rGhteys34oRyDvsWzQsDPByu3QXAjlHY4e18MaT1d5
38ZGGnKDr+7/mezHKjbXvGgbYHyisjnNldOy23XdBA90fOBN9w9GvLfbn9Yl
Wnzc4BYU+UuaZ4MwTSI4YNX/6dFCua89WfcwToxzaIOPMUlQsEmKWIXp+tAR
VOTJFvOKa5ta8+1uHFhubcMpGFiLERWrYQ5rXBCSi5c5xMDE8loWrNLkAnB8
sxxjFR3x8yA+3prZ/4kwDJ2kHtUBlGaQ8lOeKZPdfne7gRLRMm8d/xA70qa7
BXzRog6bWctHWmzWqE13zMGnzHjf/6LCM2ruGhftSohkI6zgPHw7vgFohzzR
AS5x5hvZWK+Rkq3caW/zc1mXJiHX8CuXKmjY/AENc4KHZPDPUx3odFn6RKuX
tfwLte7rfxk9tAs33FNxYYyO35qSVY4v/S0d2Mq3xPy0Jo3GPvN8gjOpXJJK
p2VkhVVN8KZa1nIrSRCHukPra7XMPiHRhTVoW72mrMxAkY4YvAtdSO3rOAkW
TlEYI+i1eSZmwGgydy8OU+Rr7UwbfH+1gXGgvyalyB5vL8tS6Gp83sb8vYrB
292wShMMicn5TE/cWMbiLkdA4OhH0S1pn9esReGclnAMoX/qNXgDwL+CQMON
a9kNnworQbIXINgzb9hNGwldgRneP8rwiLZV6K2cGevIGcMojXkPT12TTXMR
BHFk+sCK9wNmJcNTNQ36COqdG8dehI3xmEjIJmyusBEhOWFXbAxLQcCJmy+y
GBRIgP3vKQJFrjG2ZNIDj2WTrI2AlCXIBlHYF7ef9TvI1obTPYwLw+8sGqAi
VkJH/dL1VgANeWU0dO4jCw44/mdGaomCIJoSCa15zAxcKwfeDTJvXlIm7JjC
59TuIXsMXUF9wTavDzRZc0QTJrbcBUD7ccEWgshBpbUy9tOwnOhj65aCnd3C
sd8BeV7jKsLO9O+9KRPGpcCe44uNJJQpFP/6+ei6+B0R2+jgnXTQl2Jh8tIS
FFRDGx/0d83Cn3AfVFr5Ro5Q0Lg1UozVzonJXCJRZtbjowO5ACzx68MgGduF
eJSPXwm+VsGDuUbKJGN+vK32EkP1oEGKOtPlFPHT5vH+vNfAARTeSaZoF86q
Hqiw/Bn+zJ6juXI6qVye2Tt7e2HtNIuGnUkfufKycOzcDmDkzu0+N65KYnjh
oLi7nVEhTsqTXa16DLS8qPdeV0xhOVXaz7a7LF3cE/5BqwvWPWciJ8qJ5DSc
rRv8yBRoFLzrH2s5lMvlWFMZqXqMz7JCjqnQgpxa1H1vhxG+4LE9cko97d11
xaXC4rx+O7YiykhHkwnCG5WqQHOaeD7J7idMmskrjeliZYmNkhbtNESht+JW
cYTNXHKg4jXcPfkBsyNuGlR7LdLD2lCgH8aUnVV93k4nqE4Qsu2qhAZxVGIu
5EucZcVzUsQ4fCjHj5mZ+yuNiD8j8yM07RXrYyNNucFPjpHGPtnJdJ7b593Q
Un5XMWdAK2s6T18jhlm8GimfHP66g8nVS91hob8unMdn03xgtFLko9Y37Lvo
hIUHKtDnpPzqHr9lpAuIQWTLBjDvGNar0iMtLWDCHJ3zFglAfKeM650OgrVz
6u9KRpfjJa2crXJlrnIkbMvMz0jGA1qPVrRy/eDt4PVZj/RUIgTjqwysRumb
6JoJ7f41zgU5JWHp7pxdiFRjUsM2ml6emKRJz5c7RvlGT/7Pbt4RNBKXMj+K
UIgy+kqyZPw439whBBJ7hEI6eEzVoKO3XhbRL7kgCCz7l+XlVae/p52TjBQU
N77HLE9Qu2VS5hBrDQ9lPfEATTFLhbXuqdtgTz8Kj15+xNah8p+CLCElnCbd
4LRIlefwxC80wjy4C1+3zmL/78zA9EGDJQ3exe6v6LiDFweh+QN59gJxwrKN
76V0phQMsgxbYGvY4ZxGtLms+rgsqfN30zFrn2MuwW88qCc4qt9C7eX1MQtQ
9tbiuWS119kvb1Jywd9uZHydIYIwz9f4uWE8YN4rAxXV/IHibEo6pYmPoIWf
HWZlEcCC+h1+sUPJb1xUZ3iysaP3u0RrkYYUlFfeTpK0UKnttOQHJ2jvjCG+
TlGH25z6piW0ItWIk3hm2iXZPZMH7OHyyUJ7SGqMhWB9VpgJVAIKLKjXhykq
VpUdm4IwdIdwMv3LDp1bGAGJTatZ5+pHU1K7IK72Qgv85THG4r7nkyGh6kC3
6BuDgLa5PQcFkZw7bM91TN6dM2yUAssHNpv8GdQrBe8dsHJUME96kd6b2FGu
NLyryG43mrPg3fMvfGxu7thiiVpoYCFoD3CjTDbvH3sBvXu3IoaLkhDxu55k
K/zVBy0nvvhmI/LvFG3Y1RHaUJg0Gbx8MQjrp74kO+Sa2cdR0P743GCL6N7p
aujI65A4kajtys5v2+e7e8T20FbvFhjr0rDIt6TXZwqIsapuXClDAkKqCNx/
W9vVnSmy65L0w37fyzOVYlq28vTLl9wzGuoA5HBUjaFDD4YpEgJlg4YLaKIg
SrmEGTrSFWum45AxteG93WafQLY2PixrRr9rfwfe5WoxjG8KQC+sGdeBPeZ8
FCy2053bPNqNKh2HG40xwG2tt+uRRDMuhy+pBhin86jNAqD5XZThpizEZmzm
6n33pvyA1QUcTFJ8IfZfnPDYjEpMkqsO4wr5Y0zojXPAqR4TQ1z8OSCfseIp
vMSjSbOclkUXLT/6nm5fXdaJNv4ANrDtBSso4KlhlXfQw7scpZajP7G/a96U
yvLhfZxjvHpObRP4YhWfouKGcyIKGHIoYMzdzk9/Bwfm6K2yI45MASmsMt84
vuO6oiWksuST+foZRqy1IwfwHoe7ziGlfYmNco/fVssgjCE8hLbz2JiR18Gd
bnnMOVMkxht74ap+0hpFe6+kB6sQcDLEHVT0ucZ5WR3Ugp+KcdpsBgi2k4vY
MJ9edEl93e0v49IGQIXSlHJsCmeceJQaU83j4hh5HK2k5PxBKoZ8EPaGl0y8
x48KggD+hpZKbYefMeTKZQOY4E/vm2KAkQXfvwcDG8q399qU8iZDM8jnKVHr
rCX9+1iZbX7VfECZyu8E+mZwnC7POGvIWUL45aMB8nl7bsn35VtLObJSBi8/
lMvvt3KCQGfoMONIZVAo8WgbXVpeFXzH8DH4d4E/UTyWQ8nCZTO9IRlpD2fn
gUIjiChyUxHeFOMg7NbYzeSdWi22dDQ4k4/l1JJsSt7CX+gkcwMmwjR5m1Bp
iibZo7DOhqurLLNhxnpenv0aPv/gxsyQpE4gkEs7K6e2Dv2cAIvIl060MRaD
1AFd4DrOyLjEnMlLhR4l4dmDIsByAi+mcJDXnLzrJpNRoXxesBeeggXItZcS
L5F7tOGGlQqtV85r+LvVadUHMcvASPZiqgSbuepOE9stxGthEMleXqLnxOb+
+Ed5eOjR3lUZyeLcJhGxjY1V4SDHP5QBRHKqIso61ozpFCMmHaMIykE2REjr
tH4ZLuONzM25idCMexKxolIPdhs+Mib+oPiUYGoD2R9DquJNclCi6sG9zwVs
0UIVPNVxHWPrXVFPCStUbYcQsjxaFW/PxhZbhsZSODXX+mtk2pnO6i2gOxH3
NYUy9YUD+epxK4+1hqZKoQqyZ/NlAeE+PS3v6kDqxL0xo8mS3g8Z5dxsg/FM
x9qG+fBivrqEIWGMD5wy+eLQVTWvRB6vk0MYFRDPzBIDB1DjQg/4F080mY7D
vQv6oNAfUGDsu3j7hej5/5MBerJHtiEKD5YLG7Sf7C52a9tNSYddOGT/1490
3j3QfVhEboBTCQl8GK88txzagd2Bko2zwihVsJtib3lmyEFmM1t6mp4K34Fv
SeB4cTezqu6b5FnWiZavo5b4MGfTWu3NMhpF6S4t+7OqWSq0nsQ7wnM/EBrP
+342170Mjpn6k2VLLo1lLwzX3uagejKscx4nyOLyJtMD8ZTymNiOfbwIYjfB
BZFTUMg68kp+MjIwwaHjZ7xGhqidauhAm+vyKtKzku0pYqKZK8vRXsbvGPDM
KGilgm6OxuiW4yITXPWHFxAZdKSlnkU0mFVYg6s3XgRFaqDF/39+t2pde4ty
tEisLwY5c5Bab7NXyGAaail3TZSEdRUaRJpQfFgsDs8J37Q7brdY6P/oJd9q
XzmucIiiISdDBvvqxkF0hKHmnKo9nT0L0lV5Zd8m/PyVRILEuXRe9e7EOj9t
pvdCtUc7a/+G/FvMD/Dt18+K13Gc1NeLE3EMxhJGoLy6j5DalmHKg1W5vCX2
Szu5mamjZn8/GQSiNv97caXKnBInwTD2CtsuffrPVM4rTHq2AVkKauGJt887
qSjuLYXV3sOJkbdeFnWSVd/i1cmQawsnNF5c15j4EyCGMM2DzvO5etCKAxci
lgkwQ6pJH2yEIMTuoOSrgpLAwTZHRDrMePwoSdwFkMfzwgM7pWyswI8wHM/A
vsIoJ3yDESvzYYBmZb7bq0gutz4uDlkJHd61ZjZCn+S+OklPJHu5pGafUi6E
FsQk7U1wb5X3n0dSlwJ90IMFgcKkk0Zftgb+gIB2sTZYoHt1XuI9dQGYzfce
IpLk6P2u+MybsB2hHTMtJoqWhCYBr0wXu9hSO46BCDDCdHZrpCfNYhtMlPJ+
mSnYLEunMPAUoVV5HEC9Hbtvt5EUSrd/49I11ZZOb3LsLbtXAmEy7TwXUr/v
p/DIxx0vjY59K0Bdw/WLWvz+gcqV4yPVJBjQMy5yxaK3/8r7Fm7de+wWBwCR
xjiXDqQWAb0UPTMrYT8LQFjINywaU9JnCvoKI8MCHAARhh/HpUPc8bjA5nFB
egqdEIMEq7k0e8pUTpSViQJVNoXtdts9yD8g5pVMJoyB5KIpQ8hW74g5c7oc
g0amujXpKrSWGB/MQ6CRA+iMiZ+jHguvY8SNmK80CRXpTZ/5l6L962rWTKeS
TIiuB084/v9aBpfnTV8uMc+nlfLmE0itb4dKmgQfSHG9Wt0gdeR8UeeP8Z+D
PLaI4CWVAHQljoJppWWMSOOpnWJNrcx0EszlqvnZFquJM+slKOLi/kfMGIIa
8JK+A6Vb6jm/3Zg2dyz3UPOYdZ4bgFfPD1ZvAXal60FcflvbalEKykP7kx1U
v9s0/vjXzH5Tob9dIiFPgwH95uE2JXEOFgMlCQsHbs4+O1QHd7XkZ9QoMeqG
DpGa/7ippyjIfvRtQfBFEsZhQt/sCKbDEQhSxeDvvlIyPiz/qDkD85wMZ6v8
L/H+EwjBEacCWOUKsgY2yRpxUzt2itQLN+NYBs+so7nm0GunlQSgYYxiFmA4
orSc4VrhsqzKPFTF9LyFnCiZAo+Ud0IlmbZM7ZIbgU8Q28CncftVfg9ibigW
M34PY3ksAAliAvcnQlw61wfZ2wqo2O7kLEjrEtOueAshN6VuIWV6uDz0kwlS
m4gzT28yqkrE8K+2VuhF7qos3qIMSGLSJHV0uM1J7Oz+TN5kYa6f9xJMRQ3j
4fnQPYISyjqCTHrpyojxJ2+WXlXmeqU2e1xwtw9qK9nH0zzByB52vOTYay6n
o7WBqlyScJKh52Rf7+lHgyVpifx1h/PdpBsHk2xI1GcWFzzPOFGJEOJCCYXf
gNup/P+ZZ9iwZh1LxOZ4i3rGOg6mmKt80ERCl+NvboWooZoVRGchiWBL1AYI
dt3wEJr3Zt7xKRxs7CXiM46Js67QPQxygQjyO+1xNrSDw92KoBAgrKdfHj38
br91dr8tw1DIPJZvfNS6wx9K/Nh0Yn7ufRHxF7P0Pn2mQg4HWY2O49SQfH7O
t3a+kON+n8gELm4REZxbjKbf5+PMSQgdU1mlVngK0OQvl+ylCx4v8wz5sTGF
61WVRcW2z2R13QmwmlXcMjL2MJKmQBhQETpxFv7g5xu3DnGhrof5CB70E9fK
6zcc+HbN15u3reLWBWlhrZNEOiTgzS2DBbVHVTItKs8AAUGK7OLfRHmP3D3A
U2nptOdC5re9G0rKiQ9JcWFcwHhl7d+yaB6WvrACa5CZqhycf6SeTrhp52sG
QxAen+huV9De3Z+wUGjXRK+PdsyiJn1A3G93JFaMQCIYMDnPgSvkY+aPjY84
dy06A9veJ1uQsv7DoBzH7QmF383WpxZeptqLFU1MGAgqB0/OeL2igFDrTF4D
WL2R4oCeb+ti24SUMDHPaRozZf/BG0xch4/dcEluqwx2T1ErV1Bl0+ZoO9Z+
6ndGrBpqK8z+uuWc7rVJJlcS7RzPYMP4ZiNY2D3B3G76BwYaP205LXwJcxn8
9YgnwNDZZ7AB6+JxNIQ1fDSdAXQhQ2URBQhmOwd+lbck+RXhCTCnCyu6HC4b
0t4bXhETGXQ6ELduhHRoeinR1skO1TCRWNW87zEK3TN3ifyPN2i2mzFKSwr7
dBZhuREcHSF4Qi2uM4hNPGIPTAZIK4srzSjXRxMojfWc5535redKl6bPZKE6
WbhhrAKfxLksgWagNbM8hSnKsHBW8kBGmg125Q3MNN3bdFQWlPlOJNNXs0/E
jEKCQNxPoipvZBcH1wEuTPlC4O4RPTOAdaMuKP1W5ZXyegQEANj0gbgt13BP
fdmel6bKVYpzBGRIF7jYhSq7JcoNU/A9xEIZT9zdE9yjGt2izDkvjTls616X
EHjwJi2o8xP9+2B88MVXelTd9YMPnHwc2gLq5imnmTma7MneM0iqg7UF1cpD
v8Kvy3LzxSC+ji85cy2NqM5B2G4cs6CYDbOeViQQ7FCRUwgl/vgHWwEQsfEy
yGWhG/T4+ykgdFSH+OcNeqWldKpyGGasGSgGfQlDrLeuEf0jK02dNwcM9aGl
ASpTJYfKTrnII/JYGTWoVoWcn46cioe6lxlvBd6XwpdhP6ERY6S/TZGsSysY
LbB5GZxTsx7kqoBxhkvpXJbEWC2lWJeusESKMFesAiMHjn272FOJq0RCyzl+
GBhpN9x68jVWvZBWje/LjYMCBbrbRzJgGNqcIn8rr5SE99iekYthdR0TsyMp
3Kwqke6aOs70XnlVvCeJMNtNh3VJLRz6+2sB7bNlSaNCE8Cf7Yo3Nm3kwK5a
v3oWDH4PdQSs3L+/3eCSiDqCwpPGP73TLTEXT6x4ul2btZCWno4+qi8ddiaP
XGMp/fBWUJf4I17RzUshCDh/w2ZjppGM0W1CQjCH2aJdVaWahRmHk0X1sE6a
3M8XakH/omEcgknNELsVulasPl2LyhNgKDNYCZ7CLC3qmsxlVlJ8T5UB+x2I
rfPyH9If2Pm/MlZvIohXEAWT5cOeSCE92vfJRfDyyBEbRrE3osAoO7I6U0oU
JZwR76LH2Kzt+vlsRKBc2miR6uVM8xGus3/3M7/C9CbDzR/4LBYRzbS7seJ9
qsqqh1ZI92ATH/SyLDbm0d18PWc5bkauSCqYWGWBKxZhmsi2jsnc3QNI+l9J
R2+/hNhQlIp5jvOnjQ4mBSrmXiP8TwixtpdkYrjeB8xfSVcAqY7r4RGKaorN
ovAICkuUfEKwwejHkrot4NdGZ1XpnDP1+6x+UvVRKzdvXqY9iLi7APyvpEHX
KpofWtuBoJU4FK78OSCFlPmdQBbZJloTfEA/tLuylGCxexNypnTL4SPpYwg2
V8fDH0jfwm4MDUujegNmczT/py3A+A/V0AqsAEZNQ8avfFcGcBSIMGaQ2LkR
utxRiLqiRO9jm0Y/Lmt5ihYoUNGuGFyIGeSEPYAolXtrwbb/T/HeosUEiLLc
tz9SW0ycaJcRJsarQoUVF2aSuUNI1yaEow5wbF1cAkn4ywjJGgFqvGYXmyPL
7aSioSi7x0G6xa/LApAGwVHZPrgi3vUKHgfOPW/N31sT4oy0AQgtU3j2KceN
93QNALJi/N3A3k5eZcaUoOJZMmMu1uUUYHsAQwyJ6idukFQf6euMInFurGmv
Uw/yG4GlLHYtNZkepvOihZ3t9ZvnNfFJ8jSpmQHBvnPmN9rUtWKa7rD/5HRf
CPKUmgheXd8o6picqBmjvytBpx44rZyFQaihp43YXtsx8cQDczW3wWzTUL+h
9mgeTX/B922kDAxNVe5c91pGS71OsJ6ZsEGuoBt/fWDSZreeRhYj5j3gZy2o
52ucg8v4Wdm92YMnNWTHeyBxzRPfOOygBZb52swzQZcnnpyc17zEX4SV96BX
v8FX77GCgfwc2I/S5rlHfqLVSq1S5mQsyIBb5NNYaJZnJr+7N/Nc4QlPFskp
rKzwK+YY0eYQ6sRcpJTjk6zvc4S+YjIG5KlZRwKKe9xW111UMoiMFJkw1J1u
XCuKKrymYoCYfMvuZakvnecyytlyv6AAcoCZtbkP5BzmFfZwACmn4NM+jGVv
UfFDtFBOGiK1ehttzwoS8PyINFlP4Jf3+EVNu6V1hhEpA/wtJqvzXMT3FQ1G
qgLJRLyi+0eT4rbhl3bK4X9gElbEDFvYl3IP5EHUYi2dICPwQNeHLUUB8xLx
9ZjH/6J1Jg3y68wlsghUkzZzoTgqID7cLqpbtoooJi1qntI1xAJP4tIaD0jr
+bBanb7meF5j0jq2AC+p9t6YqxwaqYkJSU9hOt8Aum/C8q6ipoxO7VRoUzCX
iM/AzMZ7XJmkoh5PqQ8l5L9tdpEWVuE2nPyEcMaRSq5eJ5E1H0lafg1Otdrt
a/0wGsNSQ3PWIKO0g/fCnJrWtaxrfrjAlJzj5fSjF0ZYLzd3GYYv80wyG3+G
uNWLgylIb2YUGfHvcvvPhr4aY9MojN87ozYV0AbBpQibCt1OuL4ChKODc/Rr
heyUWV0NAb27hHMSdoZfdd3oTbRzBXzQMlTDwmRzAGh4abSGpT0Uoj1M8Rkv
tau6QiWT0nTHXYVG2cUMORBRJyNIcw/hjzf24U0+x3SXwpkLlwib+4SEdbGE
+OoZNE5gezGtNDaUq7fOHfAUITbe/SPT9XGV18fqjXNO5e7rfUxn+5trygZU
jZbF4PubHrB4AZZgHCKJVUp7EoMrdZv2n4Yqhuy3KhSjXN9SDa6rDMsh+HRP
mnikvZSKawr3aFFDOQdif9LxdkWs/xxdF3T5X3ikZHQTWp4b6pLxoP2DRrR8
axdiCUo/o2RWEKAcmZlhMpOsjxMEsdiIk0BICm8zKsg1zuEBNemPFeWFNkcK
zx1MJd26VXHF/GdPOvCRfKoMIKSklIqet1hcxqELXJLqHXUouYEOczwOoi6b
VzZDnfyTd5I/RK4u4VBp8kdB3TmFXojKG0SSd2XUPehUEh0Mt2NHeaFG7ahe
7PBHwfIaCKnvvv0gJ838AWL/WUS6anoi9Z5HTIE34GzWBAwakN7SGBQHSPw8
v8yJqNgXOB1yMwFHv/ORAkNKsUVWDPSDaBh5elnRUZmvib+X/rQu0KL3QFSU
G6Ph7A5gtiJ6+8bD01NuSmY0+mQj7i+iQX+Wd+hd2QYeVaHH9G/DvRGr81xo
Nb1WCMWq/Zee69TNGeIu+wjpiUQEzSNNr2tjgMHSVqAibJ/gHyxU8PZDI3an
IEacgBkw0/5KE5MTs1ut1CDno10v1odXYeT0BmnjKIkbrCfluCa0R4nrSJwV
syMBFbA76nrtf2zVzGZ5yX92shAdWLEpBR/EzTk7K8L/MhTqp5xpoAPXQwGE
2KY5VPU6EnfCnfrWCS4tNKsF5ljxcSH7BuY4V/Wzxhb0bBHyK3nBcMTEDyxC
E5CG0k6h4Omi4XAEcMxpT+8gi0gOECUMwfmGyNYWoIwtRIDkVBJeV4Xz4qqi
jkT76nV2URcHcqLL7l7h61VwQUSgiJ+X6lvj38JvfnIVWNozA1qjDE1o6KtH
r0oEdG4nV8stNFMX7xWM0eZ4fNAGJNGJOga+6KLig9Oc2QUy6F7QHHMZWb5j
lpLum70cZQd2IkLzEqiluHtDlH6nAhbts06WT0LAYkgaX7NMcJJ58m36i52L
n0AvZ7BZ3To36nFOAAHqoTHE0ueUVfdq8HlJoqzZAXbrxMKMuW/u8AbBaZir
XlJBbfiLtbcSNoe7QUBUiiYKC29C2s37GuK4aZAnyN8fPUyIDN773DQ+LcBM
R0mmDn4JaW/cDk8PrrdFfyY5ba0xvVW65VM8XxcOaefod6uQLtNZ9IoTo4UL
oF2PvgpFEGA3lHPZpSoE//M2u7W3omzWIVnRUPRF+xFD07DFA4xPEUhv7wC7
W3Bi0ruBLHARUfr+EY1qDyjPigm3NMaf4j9zs17rfSx813fhikFSYgF4rOhD
k+JJ03E2ETodpq6/eFr6j+ZpKXojNeRYstdRRtqugaEVYLnfJ2d1xJYDY2eU
PcsrOavQAE1548DEYjX4W/Q44GyELm1ov4D3Z/KXO4UlB+sSo5LWa1qbvfTA
UqFiSjOdlTUtROsmPFNgLU1vQ+xx1/bl4A+ovrZBDg/agBWnR8ebEv0fCsS8
3DqWMYbQ9FHc09EYfPObvV9B4COdUDFAbu9jO0NQqRpowUB8ODSJNf9pv+vt
l8tkDiPIlsAZDL0jsaxfy9KVVFVLZxe2Xw1oqCycdvNUAk9Dlmb/55VuKSuq
0i2Kw6Z+7doQ6tDmjbh4dJIlRQmSckkrfxZ0MZ+veSfDxJBPfNERpCRC9DN/
vr+pOH/sTRCPX1S1MewQUbvhcv6rsUjtiv/8tSPy/0YFQNInIcBIEXVbT5mX
dbei33gehvZpjRFDsbx6Y9WY8hYrRJaH4+7ktLVcPSnRub8XRGAvhaIkbY+v
vs8SKcQN6dPMjNs2FBdAIaf/y0NfiA4JWfAAhEEUgQODdMXFMrIyRDKwT3F/
zVMPo427q6T99AByNXPNA090KvrgQ3UjMax04xzW33WSIGAkAYGxY3pgepsI
3EqO9sWh+ZNZnB4EhcsRHjVh82W4FBcbQe4fYmuzbqFnGw5F8kmUswr/cQYG
n2ga1XERaD/Dg76PBuh9jkMASeGFXCxCfhiEj5Ftle2vllZWPiKSyvQhjs/K
uNx08JRle5lDo2ttunnA4BWf9W/oWt6JwcEGLHQUA5WS+axMzeIvm5TYrUot
4wYgo84lZFONk7zGnQ9uxMNJmktoSb+pm4r6PsxJWG9JqEAaNPy3UP+XNiEX
NqI7nPjJ1mZHpD9XoMIzB+9bczqvarMwW0jqzpvHJVcUHKk917R/MUo2vIS1
ozcWrOJNF0C85fOv9Os4/iHSx8NNOJMi2nWVs5pRxe6voh7W8CfMsZy90MuI
ISAPO96Wv86CiXGemxvJi76iyGF9+9vlBYvNvetRTue0Yq9Z1ARFzkpHjF/p
EBUdy4dFA5zWqACaI+Vd79YyJ9OL76rHbJUzeo26td29QQ+oBjvGZDcekNd6
b4n6yueTQfcuLFwP7LX80zC+nNQWf+rJ2nTCGLUSpY9KfDqWbeI+0lr6J0Mt
BLF3vVSLXElFK1GkxT0dBXf+u7Zjd6NntgR4WBz0C4T1zTd1od412p36tHgE
97AUOME9xMJkVY2+FO4i7sV4yrSP7my1vSZJx1QbK8kaDEBmHkDclhAHV7uj
crM/Rapx9jn4BRaD3rJu2qk83YQmZqYkLkuUtjfobO+Th5J/dblCWYx7tv99
lCGI9JhSg2F/T30V++V/evddIRQSKfnNGfCiDV1CHrw4IhldGQDcU/8XkZbd
9xNpG2mY5JlCF45RwyIR2uijLu+y0mjkcopkrtBpBXlm1djYI7M+RSAJl2Q0
kKXPf16BiyCXosMaKpF4UJE9HD3azrFqn8+y3nvOeqrgVUaqqBTZSBS53wSi
w4goxx7NNqM/Z8Ytd2/q5XsGGZeZIo7geSNESjV8/M0BiSqdCOZS3IkUusHh
liLJ2sl45sIcLnOIxgNrOgQ0G/X9NcjGoIcHm/mGsdwQ6IIxM5afN+aJtFgz
R2OR65PNuaiiS+ZTB2pC0Yaoh115oC3rGxShxiqP4L0WgIvDCeyQCs5b7gfg
fXjieFfUseYbFoaAuV7ZkrLX3wKKkHrybOUXjXQbbYh0SNrB6fzInZExx4Rd
VHaDz5TESHy0LiAUx0riJQTS5sKH/VLrXWOQomyCm66q6XJGhPrT9h4eG9hh
mU/sSUJdPjd8QxThtxPD3DXuWN5my3fDACf7fT5XovzdQ+mX2pmVzI0Ic7IK
mQOtkEBUYMe3gN/nHm+gabsnXuPAuD3eOpu5+tCHFDBZynkLizpuQE4dIz1T
gqnuD0+tI+loc7JTXLWLcuFx4QrJ/dIdwbwKsFgSlbwBplZgcW6ffHp9Fjaw
1Kh39pQgKfYhinZEA1vVUccT5cIJu8vI4M8Dn19b4lGBc3jxH61qlLm/hVLV
nl+xKwVBo3cIkivlsy6HoOUW3QW68s9S4bWr79LtrNl9wPTyb7ZIb1CX+sbd
Cf51OyVeKSxIRH6OhiA8joWbagNY3XD6/evYb8/okRz8ZeFdme+Jccl25yl+
a+VP341H5za4Vpm/6Y0zy+qC3UoW4XGcWZnSD4z3qjPOwHxW4w06/9C91997
cp58bBy/+yKqTe1ttyLr2wD7suQ/hkmoP+fiaSQQxDW++TT+usidzUAOqbE9
xUMP4hpVMYVlcDJJLbJDapBT1GZM1qxfeYoOXs8Og9wYVTZtqrfJh5fbDkN+
PbAJHldaQz9zEWZHHhe9FDCUFxxaeTpqctru2VOshPISTZw2G0nP1apLDroj
9mq0LAzelp129jaFf8hJZFBf224CO7SjZh7C3UpIkWdBBJEJXHIi4zM1+3D+
yUk4H9gASODX9UY3Rl95th/1BNELvotUmHjvlv/EKyJ8wVukome/ioayDq3x
oXxflhdKd7+MQkBHQrABA0kNyGInpi+xJvRowUmLnt2W5ljc5c2+budTjIvq
Ey6sMr6dY70w5HKrDC67Ow4ViVonbrOdLWL3UK7JU299R1jIaMHyBxch2pyI
AjdWZJzRNA3oMWO9MjqLpuFcSZiFnD1FGV1AvHb0RW0a8H//VG94CKOIVt/K
4LRiD8SKCWLfOzaj/Bypn65xwdP1BEforO6X0BYWVbKg524LODQANJlS73Xr
AgGHXXLQAEKOLb2ROftXDS6xBqdwvPFE8vVu0IZEluW9NopuT79OBlG7FsEd
leUPY8eAyloOinJj0REhCiqUFKzi8q1o50LlUJx+5T0oX/x+o9r5D+TivykZ
uo7m0EkEHDLACGyX9YJg/gEr6L5dq6aGqFqBBMaSK7RYjTbOoYQwuZsXGUaU
lVyDz15LPxYocr1V49/aebf0V3b3Dv9DloxqkwgonXP5kYfx2o7OGCt9zr0I
ycpaM9k9v2VunRprsnN+TkVxdooIKB4JVxqIX4bTiyu/St0RJ/zp9ZpEcq6f
1A65qvR+i/kr77HZYxYKIBBfBuTrk9diNtkSWK+Y0IfqUrIKyjMhUW60c6wu
ocGfoVUi6A5QxH9xqkrUAvUow1Z3spabTMRQls3yqnqrGqbDyQinV0ghHJsi
+/jwvi/JDFA3SUrj268lIvymUn9UoQF9DQWRifaqFagKwiI/p3sID40vxZDp
7PQpmph1mhNoIzWfj3AVkCANadq+Q8/K79pSUFR9ElOvUOj7ke0vvWZh0u+v
4/SY7ejd10gzwhU/ELS4ij3LnSIWdF/mSKGRD8tYIj4yTZmojhAtpEwSS/Ow
3iBV4HhVc2rtx7j0TWuLWoLfkv7JH7hV3dKqfg8bVSZ+X3Yu5ylOZYU4NBAr
Oy+IFP9HhZavfa3d8DoWG+Wuyy72eJgIIbbQmfAPKHbsw+5AXTvDX4Rt4y+p
JWfGg2Y10oojmd0ZsjjCESIc4N2OyN8oYUiNT/Dg5hVP97TFXIfw/4jMwS5g
rAwwPYAgkByDPlz9v+qMmo7KaXWW+ZUmYc5zfUmSlsj7C1YVh/Tdisso2CDf
hxhefxvDao+BRpx9ipyobLhl+iarpeWK9UCFw3k5ZEwSbupg1B74G6q78cRX
az3Gx3i2PbLCj8gEMN4yo4J91JTzQMcGmy7mc/u1g+dlvTDZRMOkS8j6W73V
ptbCzXA2EtuqZiSkxmi52LEdxkg00519w9URyGI9/KpBdvGzp0NoI0W4YEj3
AobmMjHBJY9rUx7y3xSB//+vNbCfZWz7UyJREYqYYB0x9btmISHYi29UYGZq
qpF/ukRT5brnou/6Kyar4LxC4jOcJwG/qgyfbZPw5Fs0XUYZPyTXQkW5vGV4
TKJAO6Gzpf28E4chxo7PvX9WXLeRKjM++b5oo7FAgkSPKgDpqaThIvK6D8g5
xc08AU+pixO7Xh3bOnevZbveND8AXJ5CgXogfFcSUkj2B1R2aE1Nq2BLqQ6/
D1NoamNaS1lN3xRQzXuamszMDZ95E6iQKlJ20go/5c2VoaUA7veDaMTbBsfY
gf0G+HXSV+Sb+Pc73R4CU9XxEGI65XiRBQuQiAfqWjLTkNkcp8QUp3dCUoKf
3J1qo/cohO96j3PT5QHrpmI8V0sCO8j0H09JLbKw0gDT1WDvkoWvX1XoMGyM
gliNqifK/aBrwKfsdbGstnc0QXSgLj7M1iepF4SHUHikOxMFqoUv4jBtpShE
XS0u8gW5DH1jfpY34CeqFJPLQ278ykNptLOSAY8XmPNOH22ZnshzNdXdcA2P
ewY5f6gtFGnQMVvQDOhp+f9S1EF8genS50iRaSnf+gcLFpXJ58+5ASEH7Psw
MDngajRp3qZkh5lv27HLQIiaBFhQFjootziZObavr8n68WEFbUIMr4kD0Eve
+iomXTSiSjCi26zoCBmhXgtq+3ULxDd+CxSDNctOP0FPxEF5VYo3j6GcQD7I
7NXIKnlN6quAcWsbGl31/9yzSwfE5VPJxNJw1U/x0xzpcHsl4EJgRjLHB3PL
FDzDnc7x0pCR2lZ/1n/E5BMgksP5um6UWcf6zxoUghFk8waDxgMRCHnrm+9c
El9bCFd2+p3xGPREGn7tqwD1Z2x46nniR78ol+v0ILxLrOp+NK/pT7v5bpd3
3YGPth53jzRbvTHnvilZy4TfsjIsvSHd4yxlhLhdNi2liCL7/YVEEbdb4417
5e5WxjEcaAm5H1u+ahV8uMUEPJNfXt10W2uoP0i9qspfYU0Y1vowoqbbhPLd
cCSKugETWWwZELI4IavTHKmeNagpNhyDx6wQ9Nln0HM3lomYszYlB0aPp6tx
wgjKdMNLkdI0NL9+/6uV6VmofBbvD/zrm2O1MTVkhEbSD0zQUI2kQZu2/xwc
iteUsR0N5f6kMZ+7JdXY+vNWFj5Ph8se9P6CGMhy8guhDuaWD6rMo0yiTR79
odTjvvzLRHqlTpMqUVID53usVdvKfPx4Q+9wLkH68iXWr0DQp75NpyYqaPPG
/Lloi43KuSKPbMxSDvGBjk5dblZaJaf8N1rZ2cbaxHHitRWeSt1/rZC22f5l
hB6vGAfQC+MqJ9y84FgmMubiFDjORBpOYp8bHBUPDoPLTGm/6xvVkMdskXfO
EdtEasds63yGDBs9k95YahcFhPhjz1Hk5zATm1LQqY80jFU6St/8VhiBoTqk
sglG1EbQe5aokMMiLyB5sNOdQAqDGhBNF5Gzll3hpr5U2WitzcDi5EILRrFz
SCwrppeHSaC5WAu2iEdMrhumWouGjOAxlcK9sytB3TSioleusAxTlRxElQ9y
H7w3pCuFSIIVLR2vgzD29VhSujDWoXh+LkYOiGabMxoJqYISQmRnjG0xsAPx
T9ZoTOjNGfsOfO5l4PFcpKP5C5kupeZNIXt5YX4IvU/li/il+TT5fbjTuKGm
rKjqlhOM5vaN/iYgk9it+2NGHPImMrS7vBALEK/u3GyITwBchzEIV/jOpgFM
LSNH4Nj2VhhOsEw/TjQMWsxcD8avD+72WvUxxRSZajdgeJ9KaUtcyWy03PTc
3bJo7f2m2nFu0UNo+WxYrORi4e9MR8zUbOrktc/E0GqV1FYVaxOMUd+5saap
ywUZRICfIq+d2xcN79duo9K0hDrA6+E4mf2sdcVUwHjQD+5MhZTSXuoIqMIt
iAX8k9PnDyTCdy72jhbE97OoKxSHK/2MiUq8MA82ZBKfmoQqE9ydwkokKjcT
z2ClcIJfrumKBJeczfkVms/JZawJI10Jd7LnWhZUSKd8jva6EW2PZ9bJA6XJ
doP4E0aOiXfWiXerrdUi6ioNDjA7L6AaMpEUIWFAdZbYAA8oQu1Ed6K0SYHS
SvY+6AENVfLvuHZQ2ifw1EBMRlGIj4QaucT8zR/+yGUCgIocPDzX1k3wS7+q
X/7TRALQIUjiFg34gFzyzhSVGn3ZHw3QzwlqyCrxdhXFVZwHoTD3mJZvYmHj
+fSiVcKtEE6WsyxoxYLeBpMKToAVnlkz4z4jrDbfKXoS6Uur+jOTLsdbOICb
hXpuCGLdHrt5f3DToRQhiw/TPm5Wz7j5xpusAczItKnL2u1h4V9Z/rDrzMta
DwlEwPw5UqTnKwtDwMfFFwVJtSYSCkQHl8GuuPTati11+TFVpN8Oxv9lT+lX
yuddCO9XPRTUsBeezlpynyiLvJWV9BiO+2LyDUyCDHzcBG6AXR4Mtkxxng+l
xOMEkVh4cUMJ5FZqSkYkXKy7Wyt0fuVaDed5UwF/6Fit/4vBQexV+tMoPSiu
zmpRdWkz2u1AiWnKP1kZTZmtoJKFVtUq8TdAnveb/9fkyPoVgMy5/MeRucIQ
ZEsaKdYaUtswfdDTP7lyWceoB/D7jsIWSyEOgq0IZn2rlGb7guyFvapjYAZE
j82T/pBVGE10sZDjULkbC+98F0/axiIn4s0deakYKww1IQCwj0hrJddRjpDH
zwUMrFRbgVedH6+W0xeZRAwvBB8lYRqhhaau2CLaK20XHc+eCm1f/10v6ASK
s+2k+y4LoiNUd7/hAQ0W6PtSB4WRpTVQxV5wJSDyZ9VPW0d5qtX9kZvowORB
zLy4TlUsmj5vtDov5qXUjaHho6IFcDJwjzVyJuUDjxZ4lI4IpwhswSVXS9Yx
Z3MFajCP34olOu3xLB6jmxrsSLEv+yX+lyvoy/F+PE52HT++ZrgwG5Ld0pzH
0+eaJ4cwwmXLAbyMjzKn5vHYTbgvB5Os1gCoVD9SyuQ9196+2PF/gEx3ThCy
hXDzmbxohho0CsgYeYS7O6v6KIhk/Ew90+vH1/4dJ5/CvnfQZlpB/Caw753o
u/49E+8EiMCiy/ZbQLjt7Rrr2ANNe2Lor+8pL0d9DXZsctTfENKWL+TGY1mg
pe17e42PfhwhXWT4MHcsVBMUQwi9Vcprva5lp6fU1ITQHyy6PntrguubcsZH
1ALft/UMr55gcjTy6gOzcF2A7QnulDyHdT5+kqsKXZAL4+d9AXd70SLyDqq5
H7rWkpglUHv6XhkSSNvWMh5ebCYc9cVYEy8pRuz0vKHQvgXNw9YV1b/O0+FZ
gfxmBF/pmany+jWYxb0reCk+y35GAH7XcsLonNXNo7SJhP2nooJqap8DWhD7
3jhKN+bRQd7pOI2YqUb8TB2Hf6h460OhwlOtVZ4Jw8kDtaDxgezndn9GKgE1
wHw4a5PxLdTeEWNHdKV9269SCH3DZwMRYdDc8wVMDkhLlxw2dGGg0Q7rP0BH
LiQDIokoQJOQtHktdQpl/4IjePdKLNIYoC4eP02D3r99kG/eU86egxE/Kor6
mJSB1MImHcQYoJq46qFAA1vy9rm3aPKOi/xfe2Cs5BGl9hOJi2lrp8Kmhzxz
FOLpXs0/haNZUTlB97P2mJo7zFQZaiDKpmVkMxzHVwdwIJEzQrWY5v6URdot
xBwRJ1Hwk6LXcUknUSa20zRlpm3JYEyd/7RKnb3VmBPz2U2NifMg4JwxuaW6
/4R/RPsROnkTrSAw5oYZxKfS1UaDMpbhmbfG6gRwX39MHhT1XqWQXeNybgVP
7VX4RpiuuCyU26dHQOCsN87PqBjlz1AGdaVYqvGpowb/c4Fug0cpmhjaxJZj
f2DNi8YH3xGNOSqfXpQz1buOofDOhG0Gc8M8aq6Z2Pr0wVmb8Av0DfmqaOYw
NbN50BjBoWVixXqonmhn/Mrw96npXKWveFcy0YHgIKBwP4RdcEh8dye2kVLK
IpL3aERalM/eFDihmvl0T7ln9ELUx4NkbA0zao+DG+a/bcNUdk+egejotXuu
c6HG5BBMkhNHsM8rqb7dIWZ7pq3OS3RRFBZpX8oiAVCKrPLuBx705E9Ufd2e
9H7ADMgmss8vDNTxofHbMOsjIO6GucgaXVrul5kA25RvuhNntfgSUOtvIgoA
EY2W5oOory+ch5mZwjF1E4v5rULR9rWOLg+eSWKgKUFp/ORhEDwIh39Tt6tS
NPgiYig2BTNSkqOeCseB9c0X0ML1jOWphUqCaXGqR0kWlH8CV8x0aSP0n2kj
98Mry1iLIJFLVsdiX3/Yk9TTD5Lp+kaXKl7f+5RhNJxvXR8PEVCs0LliCCMZ
zj8lUtFbP7jdh8UHJoNr/1Hp7Ic2c9J3kSb03bmDMi2aKXZDrCLixCyS7EIC
3d8tF/2+ZeXMDAebhR5oN9ubkRC7v9agCFzE+W651aER9E9YFBBeOlsCpc/o
/rIh4qKeK1JrifhmaQsWCeS3DRK/OSJpjPjKFbxxf3ofb96K7BPHtBX6mKzr
j2spEuyT0g+eublyX/m95qG0/QIdpAZXP5ZjphKIXnQ1OAjXEybzSEOHqudY
XPkTV/SvHLnndmwerFCgx79vEwd5LY+GoydxEk55oTzDYv1g2oNJfsbWJDKr
dgLQm2lJJv5VSuhx3+FspVOM9xzzIukVX6yqdVq1gAALUWTphdFOc1cpwgWY
ZHmm9uWdphRqqP2pQeyeW+ZD8WTmVfcd0bRTlKYLAoLY8T4arn55Ks5qN+Z4
d5S7TCt0wlJ0WAO8Rn0+bgi/cNkEA7G4E75hHqz3qSWeM4ldGr52+Q4M00oh
iS3o5a/k33YUmg3KOH0K7Pu9ZRXroxLF/Lj4MPuIIgpqg+wB7LHWVuzWMED1
kRklLFUgptkvcvRQNqszEDfhi3OW47k3GeJZs7HHmOYdH2jFTib70wt452N0
8fjQbK2g6HbzXhisOky2G+aJCJURpD2sABAWb/0Bt9lJ4zueKlTHKn/byV03
cXU4lLf9CZ0qr8W62FzVGwF5CJKQ5v0syQqQ9PbWQSvAzybLqmnRGPc52OEq
v0VBYCQqqWM3YWHBuTZVve1jhzbKAJuet9vfW4aUWg/D5K1LmQBYQ8huGXG/
SrtzOEoBV7f1l+MUDR8UFKfVXmY/GMGa1PG4YycXDsnriw4JC6gGx2F10Zu9
K5KGVieNAgdYAQcVEwGfNwx0Q1zK9Rwvuvt+6Am4sR73m6esccA0rrDmJOCl
13KoKQFwE7LZMyLiTQP7Af9p326rNLQBDwfhVrMcURx4c6+FPiFcPcL8j5I7
eFdz43UD9aXO7fwkYtxUr04JRosJkv4H0HBGZ1ozXEX5UQzx2ApJfQSkE7nq
r4RAQZsK9u5LurcZiKNGQZoY0agZAzMFFRXmK0mT7KDmsqe8lVfImO2rA3wT
IRQnwWzmjjQkENAsDyAPfUc7awlA/EeGEThEea5N8e1ozkcmww7EBi8kbFCs
xAjRO4lqdq8cxILfw3M2xUi0Vv44VHyh2/qSRoYUkZAWnVWtg3LulOnT3tT+
iYWS9KyKc81BlEcBUtLoQN5pELc+Z6kpo6W/VA+Ds95Evwg6TiB7388poNe7
NhqtiFhnBs9U791kzyy52C8IjLOUyY0Qml1MbKDuRW+/JUwe55iLHIcXoSYP
eTGzCKkqjrEKKSH54+1d9P/4r0Co6Klpr3xEDrl8gq13S4ze2m7ml1ZsODT/
7dwwTyKJINndHSrYbARSH+WJH3aZXe0AhM9EU2Yb2A99kL6wJHgkYwBAzas9
SNF+hzATGDwiedo4bZzPUCXHVrdxBzM6iCMDesRbANq4Yz8awxI5AzLdxcCi
TBXqHRSBuxvaIgFaTyf0WpCD/uso6KDe0Hk1i/OMGv9dBKPZ18EhE1LqOeJd
xWwTz9YDMxC9J7b5HpehYLRdqaU2kW3PwF3bS0Zi7GVZfqxUqXF8oKGnjL2c
P2xaS/L0J+K/UHw6e8+zUUS2EZxDzTVDhPv83op0qIyoqZ4V/mjYTBWgwzJY
TVjccZwIBB2gezHZsWX1OeLJkqicqaCkoBBMoF6fZaflo+ulG95ct1fV48YY
kanqAnaxj/GhEajQ5UtTryJ0xPnWOEhOGmdViEihCvFvyOLkpd/zVd8FUGa6
ee6ULb8hIlvvPrM3kQHNDgG2tIjdKfffNAr+E8RIyThk5g/8ES9uXVi8clXp
YVyYAcaVDi4KZ4oLxNbhFmVGKXKnaNJiKIknl75EOhfgR93xYwbFrR3ztiNV
G8Nohzsi4pf7jj/jhBNMMfqSNACYoSorC666DDq6P3LVJLYcGFKUocHT23rj
SUn3LGy9riLN+Q22nQJn0giQYoCPV1yYxsGKqbNUSJ8eEr3ofZ3KuLrDF6Pq
k4PwGEJmJYyiIu2lBJf3iLmisJuoJMrDjUeYrEJesbGftO/wt0vRS6WQ87DF
NDpPvldf1TU36CE3oMXnjpxWkui8d7aglDT2tLEmqAd6VWKT69cpkIAEJHkS
NFC1rhqkkrJjywryrCuQ06JyUNZatKOWHyTkeUCuITSj709PoqCmQY/c6GPP
WHagFC49gYGUOH8+t707LDmH+eG9WuVnBCMQ+JmUR3dELvq4OQCCSHLozr5x
IvBxjKICVU7ldr13MMFU9bpa03mTep+Ej9amgcPpjNdCxwA+RpaudnOJc8+C
TsEvwyihMlFlMCYiiOHnFhqYTSTFYZXEk45WVmwlsDlSrKliZPCw2Bqc2wMI
9Z7Aev6rFZUmLKHFxgyN5v9Q5PMQdHwwPAMaXkzLv4Wi0NgHJMs3bi/4faMm
MIpreQ+OZH52hN7xJXD43KQgu2lF+Qv1RrloiZknSV45MUi/ry3z6tPnMYX1
350E0oTVjWaILOoJWFRSYBtZhSeZPYTjERpS1+fC695AE+egz+tyjUQWXDaz
mXhpNR0fzSPXezZkCE22P901rTZLk77j/lyOWJBieGDxeVXBi50StkS+MWNi
vmdI1H863LQHm3d5tw3JP46iZtFpfMG1pcdL5vgrNuJa1Hpvfcq6ze4nHN7s
MXUKfJ9TOrEfqE+fkrpTGTbG314m9ttf8R1U7AriAHnuLZ1rcdeAx2uUMGgE
Z2k90Ig+FNXZx2i1gPwZ0ij/Mk1XxNM/unRIlL+4wc4zAn7lDlHG3Gyp1Vy0
gC8zdfzV6DBJmOm7yiFnO30Ewr2oqvSwMHonHG2u3EFkVF8lIeIzX9zgqrun
E8kfrAN4UMrDy5hLN7RI7+hPCfHkEmFMIUHMlTF4cQrbS5neLTZPFLHXkT5U
ZXSctkNnyrNG5cZEGW1C/2QIwW/FB07J0WVTjsG+CkkxtiWTVsuvWHsRdv7y
rBKVUSFlflEOVfZGGOVngKKFYeGuLnxAewxG9pBPwk9QkcjeeAGxIWwzLQc2
qMwEUZj8yFdUFQ8vx9yNVFOX9mITWWleP9Pakxt7xInQEhc+MDRezl8tDsyD
DdYFs++kAEXRFDe4gcvcfPRF98l8uL72bWzhj7DSeCAAq0b4n8ifbRQ94sT2
Ryeabhv8b3HVI9rZ0reh9Fqff/snLUjL7zsTqvwFhlTwPpZO8ORDlQwZ21FG
6TAI2cKntIA89o/mlNxOKRC7WzuzUCQdEMYM6jI6HYYHPJ4zQmY0A7H/0Pws
De2S0u1MD9inW0KO+TxAdLhCQhjrelPQotnRJE4VFpp7b0oOGClurbg1vyBr
d/jwTNReYCKucZm/sL6OT2xwyckpeI+sk9Iw0jnGWfXoufxdJ8fgKkRguKoO
4ixwUibjo05Wl3pDToSXC6keduf6Z2xli0UEqvsInVjTiSD4jEOPuFBqpRNc
Zp4UI0ENBX4WMoZmTRuwv/Uh/jLVTfGaq0MjNkaJgOZb4tIunGIBaSWq0+oB
N5R5q7kkXHBRHQ7/T2sg9H6cT4Dpw0lJ3llzhvCj/WY6BdHtbKv4Y4T8BDku
SHbb3oSTMMI/V5rI6Jc1ApoB1zrkHdWABB9vRhEaXuyj2QPtoyGHFwMa1dum
PSeZDtlta0pSiRslCBbn2jAFyjLpLCrz72JvLlD3kSZ379umdCBXponOXUjH
G/Wf955pugBQTQQiij4BtyREyjSG/09xkB7awL3ZLSUjTowo/Gz8KM4DGani
FRsTlJl5Eaip7DLUvjxeXKmzEBK3KA6gUH+ZlCp5uNRcihJm9pWvrM6XZNW5
lMBO9/ySqpuGeNSfZCnRMNQhIs8xT1hnka/8Bbd3R/f6tdfizo5EqD3ODU9q
pX4PyoHDk9EeVY0yYdJitl6+IvGsS5BqXlVQPHPHF6JSd1sBYQ7THNjWbpko
XeZJwmqVDdRjBdEvW7W/257CDfSAOOjxLb8js60g/a0EOXM3+sVARNLc1P4I
fyX8yTDELYmeas7ogHzeNW/wCrE3sPiCFQyIC8moPEZ7X5t1HMjzlO5K4X9P
pHpy+AFiBZI5etMAgFbG9348v8WAtcRJKZ6ZAo4tUrIZy+dpKjF/65XURbgM
Lre4sy9bvS0hR2SEzMn/BWV18d3wlM3myvlTglxubJTvW61owgZdmVxT7mXb
ljzkqt/fLviGfqDyf5LsCTSt7ja3ZBjxhlKA4ppIgP0VzqSQ6+8/gtFL2T0e
jY4fTaIajirON2vno7VDQpiswULBBHmECjRuaoep9MopQlZgoWWYCGKw+d5u
gqxCBKz2VvcYBxJ4+W80s+n4s89bycP9hAtEkXO2fZxmHaq1jVROXsiYIVcQ
0OV1lQnFt8t8B+CEBILz7IO3Mpy03AmNltywcC+c1nngSWfb53C5KRSVIAJJ
j5hi7crI9G/20K4J8XELDOONNMgfLas09mSkYfh4T6+NWFHtgRqw1voeG/aO
SMFj3Cc4xH9X3TVOyqudQc8m+mEV51w5hNWhbbVJPK9VZJfdTKa4CZjNqZB0
rHa2mkEN+IFJV0nWdfb5cFKjuF+5RAgQSfhiessCekSePd+MHoCu6FDTR3IG
LXtoPWUpaNs5elzbtmrXX144YCDhnX9y+HUvZ3AD5erlsSIxQR4G1ay66Psg
G4PwjUjBAVCB+LyytviI/zy1LnqY/5lI5UbHFbsQ1WqfEJSxM966vZhWQUAS
5Hb5s4Rzj6NY26cbZUAAT9qa6V+HMHJeb2oFWwV7QsYVKXsM5W748jc1SZeK
hVRENQmBigusljxt1DjonuZO/z7lDdnOAGvLMRl2q+mz1Hfetra9Yw3qSrxq
QXUUNyiptgChf37Nk8nBdbUzN41HUvuXRozsmJfYqGEqWXbRA/P5DJdqDwSK
ES+/3veto+GWLMxRJNSznKOqQv4L+zGALbIK2J0cxFVqH0U6DL3zmQH3GVtz
9Rd7mdfwa1FsJQQeSzw++quoOtQ1UkSc0J1FBWMJor5TdwysFMBOzh62zxlV
wGpX9uL5HWPrRi1fhAhxaKA2/+ODPlkHBDey2G87wCSJi/VVSYqIZD2HLbko
rFsw2Z3r+DIYZvyD/SYZpyCN59lbnSrlJyILIV4WewgQ0cQj8MrKVYEYl2WV
j8DJMcRUxLGvA32K57Un265g1+ziZ0AAoUfMUP/Dad5QnTGkz8MMl9As/ixx
WUoeYG0AbPI2gcQm8udaK6ISM5eqmX2D4F7b1T4Gw4t7rytO4Z2BYUoGtD9K
PxH7ewGZNtrHfTWedi4EDV2dIOfodex7JJ2T0XA9QkJXEAGKandOaktyaWDK
nRK+Y9kX0IAeIIgCXW5Pz4OPJJR7GkmV4c+XvBu23WPR6ZG86OMoN1R5Wmg5
cPRbKv6xCLpjdEQrkSJ5KxJiVnOcE/rYKz035gS1Rl0cNpuPrxr6Z6HI3Xs6
dGp8ToqUr44ibM9dlZJIgJg+HhMtDD8izZCQ16ZF5CdHUszdrHHAMpSwy/I9
OIZl1iaRVgtGPp6or9u/tQ3GAQM4CAo45fUialplokD4vMK80qPyLKdf5rmF
M4B0n42sb9MbHMJXEDfVbtf8kS4cf7I7KfaU0R68OdhDsRD6eTLxmuYh/U+o
OXfHn/lGbjRxMy4bhu5Uu/Cn6I4+EXolkVHJFebPZHKl5Bodxm+dmfn5zWwT
yaByEtw5GLoQACJ6q5mOlJ+QMAXKAykva1DclWtY0hEQoxU2GejF59d1CR6S
nz3C8162lMY0SvRUzrqHL99z+ipnKcxNO7tbiZn00usCqSAfyHM4GUk3GH3j
HCLV630WyceFd4DGzTsg/kfatyCQ1/HRPho8OITNYK0jBv3e5O5z0F5aAcQO
NQOLAEXfxdHbFQxb4c8sJGA7+lfs8P5BcYPT+uTed81HcQlMrMgDrrcIYVwf
UgpeqQmyGJQNtzS4pPifi0KoqUr4f0IiLmSA8f2uWFtUuuebVwuRDMsx9Bb7
AnnDp9/WgSNRQ+niBDV99C9PdJcFBfCTAcRC6uEmc+riDRzdfqj/Bcbj2FIA
SpfWGd9RHkzZAK5tjWk1bkMunzGy+tlbA/GmXUmfe8m4TFBn8E7Klo1X9m29
wf8ou8FjR0jndI1vmjTlQbSLit4rikNRjm44NMLEruG/YSwEC9v+TGqjULWz
FQaXznJuTboBymEYIaq3R7wgynkkSm2XU3/eg8SSaur3i5i8rX13p4NoXg8D
kLRRBj0VTq6vSoah41hHOAk80AYk5Qk0jeI+/8PsHu72pBVXHlqR1oG7ch+Q
ADmxGCCIC6s3ArE8eukT7DOQsU1PINuOK15tlZrTnSgt54tO4sNIhuszrH42
O/h6dcrJdeCxLptaoZfHR9aNxCdPBhSYwllJWVPH56VypoFcGMRA26dbvtqA
G5ihhkhEnNHbUmrBBtPXiOqfmUuRfHXRZTDsbdST+PrftEknUmiahIr6ztx2
//zz6Vk5DQzKCFsFfIkh238ca70WqkBvNYmEj+kQSfG3x4Pcj2t+LTLwWkKp
KDyA7lZfyIThmvwFxEv9Euji1ElSHNAJnQK3s7LTwJ0ArjjGWkVHaAwW6gHS
ZHh3l2VXBEIqCBe6xOFmDOa/oWQmPuEg9GqaHzN71+ASKFFFG09ywiuZNxdV
awYxP6DHzxfAqZNXRtW560VkD6dDqlD3+jMbb/oWBtVGDU6JBcvaKnpUC+zU
GlKnRqtoCpe716kMtlA2+o/SH4rXSIM0GQpPirRwYiKbES70HGVFfDv2blUK
6AMfSQ3CpZe0tgHrDhPNyRkUDo5XvkJB2/82KUI4SIz/veps3SPMPOG19TaB
8SfczJu/YugMouZEwfOIHUBLHd35MBo2R4J6VnT0XGU2y0SOm4PyRTnXYVT5
mWpsW0XMWqVtTxkmRCW/QJjmY7W1xyfcar4/9aiwzYS8Vr9pkpoNmDztsBD2
BF3VgVrlU7sPJWRf+8XvEiQbHrvypkOFaHADXAgmtfrYCdu8iFGh2U0LkcFo
1T9XMutQcCKgbloXv2YyfuRtCZxbo/VMMVDMTr3NDe5dgx7cf1EXd5LkN0Mx
3wuyNRd8zTFHf4Syohr0cIiG23fph2Wtwbb1gbARETbTr0f+uAHDAwNFIoSZ
/+SpgQ2YT64tfdosTL1wPduzWm7YfZf8VLWp18ijqv1rhPMEimWmQi0O85Bm
6iU2D1ZkbQYw7jCSt/VeMPEpxQ6ZQi+oMLorLFoiQN+rJsJp7L9QoFPn9LFB
zZvOM+CIEnnZVYPS84zTL7srcVO6uuhxdDQdKvto60abxvyREycKSrPjww1w
YkOGL3GgXZbNhPGwx++oSgD5jkUF4Y7DkeORHQHyVQCka6ECBrHwSXi7qOER
r+V0rbroTi9K/yM4B/UDCUsNTfphh3cfIsPpUfZWLDbJF+gYW3/lo+1m/DOL
pao84OhNeM5XwFqZw4O6mP/rQWd/VwG1m9EqVjim9rjbPtDxGzTv3gB7fGl5
u5uws0QaPlehK7gl7+OzX7Oqxvar4QoNwjvZ52pN1s6BNqOxHSOpGYfKH5MX
l8PLb5xWnkNUPXGTrWFvtoi+8xCiXHQ5kXzMNeMLxBa9STm2GBZ0V47SSJOm
lk1ZJ05YTBGksaWXXoO3VJ58RaFIWvvvAr/Wk5c7XaPevu6T7/i+lDOGol8Y
ljho/7AU9w0OKaY/Vg74RSOjhTYv1DKvePxbGW2rtvOJTIOjmyUUIS/mIcsl
UVcky801m6KX7LYz4erxhjwJMhGtp19EQEw54IKdeUKh62lS6a8NAcMGeImy
tn6Pnh8q92UgKfagptY1ymNpXldc0rgP5KMMmpF03OItdFZGAvL/LJ24eZK8
oXUm778wE2bEmpd25nOGYHD1rWHKqDq3We1awunYL0hENHqo29vJNVOKCZSe
XYa2mYvFVob4KQ8DcOPWd8UAaWtHRrUqpN9+2d+n7RaoMxcPIwlJG7ruTtAW
K05OLRks0m3YEpi51siGbjgLs9hPPn1+QJ1xbabJf84o3W6X+UjSkZ4D4QIV
/vKqzkgf6ZdtjANbde0bOsA5P3xsneiEKEpYXWHc3X9PgKWRQlujH/sy9TVV
vUkYXadt+9GMV/6+8LkXtGe9wwm/ggSBsB/k1wNsE0s7f5q/bD4jCfp08QSJ
JJ441nyIorU9m+fmRyQeT0IgBXtt6BJqQZdCHl/ZNeUxjAroTUl0eXQjXpF2
aqZVaSbeZTwUkB0RedKEzSekp4GCqsx10mJAV27FmlD75q8kp1sIVL+fusQT
vHxAKZtw/IzLoXsUWl8wdeJ3C6XyjYQzHS49PQcX7ym+AQGOt/5EDDDr4tIh
LarwdmbBFmPlR1qYote55lkCCy1WeViCeoECiewNd8H6PiPdq5jyuwZmbNeZ
7cPMVt/OP3GHm7Ai8AGHfRI92FPzW7OARS6cesHCMeGKnRHOLavhmPbwCZOA
eneVgJ2XVmUJMJEh7cK3lUsP/YurJlvthbh3IdZGo1J5TphRnyyQuUBnxngH
wyqpINdH7yYPnVyuPEa7Vh9wIz7Wsnnxq8P3EX9Ly6pt9GgvqGTHcczRoqNN
AZ7Jx1DH3KZ2EqNMCrDZqaRxMHhEmJ7aima/mvLPWzaNV82JOqnlqtgYJ28+
ZkYIP91YNVYZgFiqUtc1Nl2MqS1hbqljKF5+SR833GKurUrPczUV6BmvMkpL
H81SXTXfS4hsg/g6tBjDy38FnvY5RX9cAn3xtXCI/Ypl7sgyE4Eg8W3TVdYD
/lOra9kbjcFdai78810AXLM9XMfJ0vqeR3zv/tBoQJK7/wj+MmolUjKZxCf1
P2yiW0mC3qTOEfnOeS2F6FCafVWk4Q15YkVJje63bSvWMR0MGMUUti/qta9C
xp1cMYQzY7chnyAwB/N05MQMH8lXtVFDjCz4oZhjkldpXw5XEE1U0lh59rCH
VAyX2u0vkk35IwcbvZ0KU0tug5vLb4jCfK9QxDXkK2YGkiXaQM9yIkc/Bpbe
DeGuv/EBkyo3+WAu2RoOANH0CwJ5kTTlVe2zw3QnPQSlB4OL3TzyzfwN1Wu0
midaCLjggIToAHvfjDlzr6XXekUCEzq09NDyvXo5JzIs7ecw6V2WEHfuSE4C
gjtVeofnY/Wix8ribKi8u+ww9ItXcXW3c8f04bswpOimGx5Naskt9FBjBWTY
qCdeFHW5ok31FqtFDD5zAUkYFJ8PzvqD2HWeGq5n/GrqixfEiHcfLwTHVjE7
t97zsgzDUXrHRpDGm8UF3jIm1nP00UV/68jJdNvdNOg1NRFFIczsqmBn3uJF
wCGl25VwTxpvA66cgNvrdWO6TuN7iFTZDzV+UBxeeK3zfKXWdRR5RV8lIcPR
HCgZXUUIzMA9SIO5FdEzsfgdaVzpEEr8mb7uQZah2sUbHJmWet8QrQnIA+gP
3oG7xDJtQ5wcOVTB6A6L/xJTLJlIELgUy1VrvJb/nihkWsBLwbdZ4PXEgqXD
KBlEuXZzVitRaexkbM3+Ki2LM5/fpHMhzm5HIPaOnxlq/8IAzQlrvb71+Qin
S1AHqvKpBk0PNJ5i1WoaLkL7L5NyqBQhbkf5c+MCHqU+56+TxNx2WcFDDdmj
mauyvQyczGxGuqxIMty9Ue63zWzDOuf89ePFe4G02TSzi4E7Eks8yMtXECSO
kYJtmV3m735qVCWDiNJYE05Eu7XVmKm+USmmrQix7Mi5zu2TJhYKLqM/1mEg
WrbjHWR7qCuc9X2HYDh44gN64sA9kFHNsataOec7Xmkf4/w1kagNLn0mxuDK
Wp9C08isDYYVF1NbwiRQnzVdmIOOlKyqoiIpymkFzrdn6zshqtOvZ2nkefgM
GBaeKYc6ehAvKRXo9elVZm9KUIr3SAD/IuWtoUoeiecVq7Q9sVrtS9JrNEfe
f64Gq93hUnphTtHyKvgmhX+qGlgTLyjYiSi0f+/PvTFm+EFQXYrHRB3XITnG
2L5naQVhVavIapeZS2hA/c+PBBnBV7Qd6B/7c1+lLMdSurqU9CovAEgFYfgu
UZssNLi8Ckcio9cfC6mOv2NklVW/yI1FK460FOz8TcqJGH9UhoV2F+x8Ek4x
o174QlM9L9G5k+YxEU6Ugz3BuRpJDC09vKH1oysPM2LsQBhNhjHRXRCea3jX
p/daG698coI/6Bj5ccqaM9sA9bRRvlxUOTlr7yFHRkRgo/ij/DxDBlzP37C9
eaMb5Tr7wj3VTIU1BfnIrTPjzQMNvh/u4o6wCq4Q8k/WB0ryBFcQJMc0VgpO
mcx59DG+En7jxmZSs4fZnEZ3ytyNSPKkYCDpDeekrkKcAuLfqo1rJsItTIwR
y8UzmgLfN8vdX2guKgMSpR8vKMSKf5zTv6NhXvmxWjmSRB8mK126oSeGWUUV
fWXfNC4Nr1iExREvfoFsg1O7u9X3GFcwzWKr6hHN1atPs1/brjFBrd6ytyGG
5bOdaASRCWm4l0iQfSJXM6X4IBWY6uivwlICA8fPtHaoJM6ClvoZET9FnHDG
KhJdLJQBJuLZuZ0JhjwIG4UZPJyDS0dnEpgImEUdsVIrCK9XKJ77HR9Q6AD7
0aAl10Xvg8rWcm1woSxMmsRXcbyIOSOh6JPBDHiYzI4hS2+vux1uTHFOkFCK
zA460vTOdqcvWnkgDxiiognfkRR6hJPVeqbllm6GSqVt0NoVAcxcLAwtiztj
06Ts/bt38mUDKbPUuuO40A1Wa9W0/Ge7/cLJxR7obtqhUwUtDpK5Zij7yH1A
FtZCfPdNzr9caOu7a6C79KOOSYKXkdAj8wIboPV35qQOg3gy8pMo20i/DsA6
I/2nFmlvx5TQQh4kP0wk7pYXPKP310gTLO3Bsa2VX6TXyUL0C2O0cStqoRqh
gZ2L4Cl4evwRkqhrZacjbY5o5EaOqb3kbOx3lzyJCFCb5Pdj2KyDEkLLeaqQ
NQC/ggUEo/XELziI/SKhoEE6PRTYPpwFKCv+D6po7fj9oGa/sQ5oIkXhG5+k
gBhsjwQmAn7TrelykbzgnkhbgoEiuS1IcKspI/Ko5bvxCKXhhcZOTothaZeY
JkOhcg9Ibp0jlxiq1zMCimW0xmIL673GCF0b5QaIUk4TdswDEUCHpDytmRaq
xSBJSWOxQQj/jXWrV+DsI28860NltLyFPtpZkBuJ8xd9yy04hIHYuJpZfEL0
HrRDe9FvqMtGZHzZkUcwqKr0bsFVDB97ZdiSWCzzCnU4Z7xdu8L1PeA74bzb
5puuzp9QLji2nGrI+FXppfrkjse+6OYRYymuhV46pJXvU5KrBRrEPjq1HOX7
mJTg7slWpw9ro3BpKbOd+DNelwFZZwMPxP7E1uXhOdgOOQEZPRgjoyVgaNuj
uSG8XocAFqbZivEx7UZXDSOrS89lRX3Oq+JI4BZVdpAy9PVhkBHB6rGFzeFb
c+WBp1OP7C8s+e3JM4ASBAiYGYIO4zW6QATXFv8qStexD8bd9/zvcFsHt2lH
pBAKZguSwqPh8QDoy6XYtLBfv9C75QDVd/i+4VfUnaUfvYjt/nfk4p8VDuhz
Hq6K+TiGEBlFdWAxJTmJyEYy7EInrfb5AyV6QuF7Wj2G03/Qxg+boG6j9H0J
wtvzZlDRgF0aWifuZQP2UEDn8pEZGjnhqFD5wZSjETWkvxniqm/JsAXcv5Qo
yXaKCveUKCQubMQD9s+EiXqd0NFo7Xr1nxvacAa20QE2E+4vLnSuBtvFcCGt
rmjsIczk3W1/C3mm3J6j/YBDAFhSiCmq1g3utTrQVOti41NelNZrlf7eFTdt
26hzULAU6mIzAyDZLovdBM8ahhMPnsDOxvUBE8M1iEkzezSKOxU21fBGtIFD
XMsncp+h7LVpwzBSdyh8CddmlDAT2VAYWueuCXQEy9yy0IkmYisrBDdSqhx7
WWB+x4x/TOXUTh4EqLaw+WmnomOsitEgAkXLkWzYAAnvyZu3v55/1vwIbPhi
CwIzgwKQUAbUIo63AxIBxOT/gPAf9NNvQxoXsxQw5VYtxMlg5volRp4mymZp
///8Bpip1FsQU9c9y7WX/noCxwvZPyRgS43uXrXttS2LpqqLo9mZeX2X6mP/
rFqHwuO50PUB3qBuU9mfuxOoQhZcfu1gpBv+TKuMgpxjYhDEgBhmQ3xfmu6H
rKXD+fYPTkE/lPjs3Ocf9AGBtMeL+GsfH9n/Nz5/fLY1/HKvsiMQq/G9c0c8
yuXrFLLy8JtY5OszyGoALZqDo+TYCuOsPoIdMyhh+9bndPEFXka5vDktIoy/
KvF2X+RqRa7jtXALs79s+oW5FMM8ApaaK5TfBcdWuE+0ifITtg3bYPDLxb87
VBIJ32uem7raVr81kptUD0YK48kPigqmjEqu2pknEEjpq7Qi8Viu5bF5XVgF
QjqtJJEEpJRKWlQO5c5aNwi3UkobJXmKzBOkltZBPUXj9TdmVZQEX5MNXz2e
yq9w2MMFtSr6S6L3+G1GdJRlQdBCuy9bNsYmqV/VqnJtfeHMUpDr5qBXH2nJ
yJF7TnUC+oOGRlujpcNFZjMCi+qBg3AbylW/ZLmUAzuiPN+SOGB4YjeobD4n
NPuAVLcdOpe8dov9AmbtapHcTByl+amsNSOmanWTZdwhSR8UsUh+a4DuRzNx
QeynZKcnZlYGcUAOAKqwCs+OdGze2ChQer3j53hXFitldt5ILDv8+4VE9azt
ZBsgmokdmwY4YeNIcO/AfQzpmrHpj5Shu/QU6sIWS9QzJPfWlwtCIPzzIzFi
K0T2yfC+Yc8rGgqaM21QD90D9UHRVgH1ID0H2lRfSobRJ/bMLcXTd1oqFKTN
PKZD70g3xqw5dYM2nmV5hKDuhHiBvr1XhwxfaDVZECFsHTLwaX2IGuJzHEvW
vaW3smo8KDw6oO6W8i69Zf5agk+/aNh5elDcp6xJy74T7AZU2C1RDtk5F9N5
Gc31F7Nb2fR+z30qJ3NIUB3Og4bB1lIrs/q8YsSJAcuHF6kMnKj3iccnuvi/
9EaTrHh/gJooVhw+brJBN9zH4gfOhrF3Zf5kwPBKXvjBqtdPECfYTZdwR65w
wB+yLSZ8cMwT16bYLnnOn8SZF2R8Rr5PqSXtFkUMzxYHN+67p8L9d1bTihwJ
XL+tVUviHcKcGNZadS/Uemq2tMo2qFfiJV9lGBvn4hfqBPJCwFYwkK9QceoV
qDbCdiUdmdeQd4IxpIxef4W8SMSJUYFxOggKLVYE3hdWjf5kjo88gRYdmE3e
o+QQ0Hg5rMuKOJFm1buP8HBZipMGt7feE9R1vZNfLlqj3ZKlAVsjU/PaPzYk
ieU0PNtiM4tANAESsKgI2Ezsg7KRpJQWtVpIWR+pBAyRCwnsvh5q0L27xSkO
A97rueVwDf3R021PLiJhYreXu9UFxc2Fn6jivgceWKhlf2T70UpefkBRR86Y
w2GFE7hQsoddi/3eUttxXYU4prd4sthqYg6BZhSOg8SOTD4teRpcPwkvRQ7m
Zodfaq1d/ziX44FxTEo84u/uCJHlr0OeHJT0xSbgYJxSX6lX8YV63L4tfGd5
9brHKB40uWyFX50rf1/32PjXnJHp5be1ftwl9qhlkLUnvzZ7s6w5H0fhKPDV
IlAqmzo3LNsyefKGESio0tLouwquAW1xi8uZ3p+sRgQezOTLAPhJr7OgD+Vu
ih5gjHLkibQ+7fTmMztznKkrtwp+EVBgCNK6XXe8bKRE0I/+j+mOeB/itMen
uFVd8Dn7aYYmQ4XqsjNKlV2EnC7oUDWUykggnX9Jm7RVbdVxY0AorfYeHtF/
7qM2MCHtN81H4RtCCNBJr4mmAAc0nbk4qZNMfmuGwuI81E0IMnJy10HvRf+8
WA6C2GCjped+Hxw0/Q7WAOI7RwIGKPhRiVuUw3AMkCzV7ig2lGgKcewPjrML
+QnDmeHbfhaseYUswChkzN73MvxsZpYZnbhoWC4cevPSC+ArsL1LS7+GPT/v
406ua5TbCpBfqdWaTTDte3F8dfO1t7ZZ8mTSdinqdxhnJz3RK41jzKqRGNE5
myHLtwWlvuEUWQOJToEB6QHmSzqQQRFTtbLAqPHVMFCZ1fm+d9y41y8tQLec
IKMs1XqyJgAwHP6KINBuWfgX5XyZH06TH2+1snCw0wSj0mdfAhSdbruezCsg
Em6wNkZu9c/bNrnQ2nCoQmsVajxTye3cXSqZ4nU1IjIS9nr3ScKdTbjZtWGa
v5NmJkEUNk3XBfZJfYn7U3zHKlHZhY/bJbAagcMSH5yPrc5QJaasOGAf+dSE
yA1hOIv8RxZifF2MZEv7UUT5GRcu2IUr/10HKo5QnmskSX3i9+Qk5i2l84a/
UVHbE5nLWnx2HhzsiIKEcB2SfnhWKfse/SqbL/1Uh7/Tn4v6jxw/6Q7UVpFz
1TXvjGpD79d8o1og0nP0R0NlGziEjLHpwXduPuzdjGzmjXNsnihmfzqNzK3V
m97GRW4nR46dNFHftH7rjAKfAdzqfyYYJIvo9S6QoVO4+rkRzqMZgaUc7H2y
WjvObz/TY5GDNQA87NWUNNSTKDlwmmQxkbjx40SKXm/6Hte9BFb8FYjYDigX
LOR2/otppIiqx0DkhIBQm7QM0vZsDhxljj9nhn/QvAiyq0BQBIo6jaUBmzA+
3i+tx8EsiwbTFtND6o48Bn309U0Fry6/X8kputuZdQr/gSfy7jSUeOZXgk2B
HlhMe+XRfAwKQZjcNMJ865S1XPMZrza+QSBzP41s47Md9LehD6bpcqNo9wvh
kwXEnT93jXwEdXO7ytqGUhWxR1kwa/fcIlcvX8LXbvW7LCPGzk7+PdWf1h5M
yERd54ml9UNlHSgr/I5hoZwPAAcxWhjherQ2sSLzzxYwFAu1VDLy6NpE4j4c
MFut4/35Old8/OjE6YiOsC07+lGf05HTOZJf48lHpYhcLlJeR5JS5Jg+1644
A3Ba6t5jLySX4VX6r8H/hyxlXQDHS4s/cVpMgvFdbC1Ux1RmFKR3vGt+QniG
Qtuk32J3o1PHbi7UM/XpFBu5kpGbb3IwmQqirikp3ewWazY76CLSUahwwOfX
OkysmbJqL/E7LrPRyfSI665HTW7zOHzi1cAjCDA2/81tzsbmZWboAheM2O9S
ESzMwA6OUtK1NSmkbuo86W0KVb5RnndOiGkVpChLTuR5tDbmVb+zVZ2dqRYr
CeyGtm0lY9zBE0bRxT+XrByWtmiB9ilJqS+2GGbEVlKYrjNMHg/ccHzoDQ2l
OQGGr7J26EAH8CpKMXAXqZFlHmvAcpVtwOQB829GfinjeIBYm4RpFjn/Cw8E
TtcAkXOx21dWl+aniv9LfdbVP4kJ2AOvQqXg5a6/+Iuxu71LSg+UXmWPUOvv
8bJno4Fm1TJxNxjl0mBsWdyxLlWOwVaMsDSrko9NZfnwbCIbjLGojSBZy3aj
Eiob0lya7oMMKuWQDyz2QwC54cd14G376HLo+Vu62Z6M6EI/xiUDozy3+OJ+
xAOxvU+c0tYAU8w0qyi7Gbf8AJaOuL+QcdTAPIqZbtqbsLTPgXLGkDLxcmfx
GigwcpvCDR315466J6snfBvL8C6p50cv19BrSKitpemWqsHVjwlq+pDU9MSg
D57aQkqs13d8Z3WGegLGOcakI64iPQhNPUGwTddBpvNeoBLQPzIxsGvlkznS
tcvlr0y/Q3eZJ73WvP7j2uCeDRFhH6KZO+KMQ+D5BOOHBFuiQI5IeGn6BGaK
qQCHNutIKqPS4+xCOYkri8rH8WMpVq/cIRPDqJLlR/uDURLheXa05f9SyTUZ
AfoJP25/JDtajpYj6PBcstb7gsf3TQx/V8vebOxW+YTjkEDxFBr3xA0YqhIl
f79mXpmMZIRTBmRVrO1b7lqxc6OB5UT4c8ncRtl63sph3SUi4SM2RZik9tc8
RzgZC8xQj0tdx9MYDVDCmRz/8bvMwX8f6mL+tk8aKltvu/PKl3FzgVmm8fKR
O7G9aJh4PPistoEoQiYdUVRt0cul/VlH6tp0CM8ZEzS3YaOFf2zoXd7GjBad
lr0dCmg+SUBIeF/6O0o6DbO2+IUL4CCLb7H/zA2ndLPsOWYsA391qwsgeAxp
p1JvGvLNfohfFOQHMDlkwttoIkAKu8xOkIDNOIsDJWKWE89rBaplRaL2d5BN
aNi5eZaoEJBXMKQ8fxTzfcvWNZkILSKata3MJVS3+Q+tg5kl9ar0CfFDCkQg
u7bQP1E3ssWxwYvhIxGVWhSa4fpCGJrJIau+PIqPH44GTjEhKRjE0WZuMczT
wh8uytStOdXf8HWl8l3ueZvMVP6RJCsM8+DcJuy8dzz8D5SEPlq0zQV0dADb
2YIE/fI+HGJsufQP8YEdzCp/VseWBB+E/HOd/sZ4dNJzoXUrv3U+7wXlEZMm
KtouSnvpoAa1tbK/eZG/MQaGqeDlls327lWsPZG4SgfZyFQgnCdkCl2IHUUw
Mv0e7iSLqEDs0p2co83Zw5Mq/lGZZoAiizdyDVkf1RHzrIJwOzp6dswVJuYi
f0lJWW2tPJCtWx4r2Xjyj0n9KrOUvkNz9vNHylkJEnk7S/zgkICAvyZ1Zg6J
FM16l1EajpHjG2ljcSib3yD3xH1hx9uW7YiYhIL1apuehsMtLcpLPT7xTD+m
qEkNRbMWpv7D1/3sTCZEFJ5w1WCab4g8dqD65OqFnhFA8gHyFDA/i0AQXqiI
LR+VZHtcU8zf8shaZT32FtdDLNlDiEBw+/1Q1UiKe5Ppa+gO06k++Id3zctx
BQ4q88VwlQJCpSmV4jJkCxBnS0CB1jz4prJjDXY9Lg2+i2eVGUZZcaq28bjY
RJoKqlY1P9Gq4cwahjvzQbB1Mq4plCgLnAtP7HVRRGFFa1Kj0TNuLRoThFQF
oMTvSaP/S8OCaWPgmw/xj7/xEPtcQN0nUXJuSxbfFyIrLAordPfcmQRL39/P
DM3Gku+d8aBghLUt2Xb291TEVp46zxBIjGbEkHqj36fhGv6o4Crtfzd7YfIR
DeHnKlOxmxfVRc4ePT+wBOh7IK6m1twlk2MU+jLlgUzjIqG2mC5mJX33rCOW
ZOnB+CucqgN9vg3r+PcQHTUuKLGgbVSJuiNIZbA1dLG4p/6JHkGTnjTT8F12
06o6mnDzjGp8UfTGb4wBuB6FAVpHj4h4TjioOcvurTHWdp2J1laMysr968iX
KUR5qVnF/yvOiONJSMK2E3w/h30CB8603RPGQyl4A329eyPHRC6wOwQRQHiq
U97plJ2I5SLdhTVVGS3fg7Bu4q8lGYI/RhaLX5TneTuoNHXT/vhP4O1QtfJN
WT4PHzOELn+E3uPm/aEPPTdEZ4igfKZd9cdfiRSD1iZ3SGxB3MfrPSkKCw50
O5/s97BhyljPzsgTORSbQxtQ18UtxfkvnFvo74ThNw1VQDIbhN3Sfto4HHlF
64RXdheN16l3FJuhBPanE6YxKp62geXr54dXemHL5HwJm9D4dvOfALvcTn8A
ll53wVElmeHZONSkVQZiOrNk/vsPvt+mOVopJ+FxfqvWE4BpYHeF7lZ9XG44
8cq/3tf0kCyDH4snFqIXH2/f06Q0kAq7fAN1HlDoGNPHntErBmQbyefcSkeM
faRuMpgvwUu4mulDTy8YXLtkWxTbZVM2S3REPnsE/7mp4rCfRW9cNQNvXS91
JMqohJvhrhxmI7q1Mxas0DdtEcoF+Yxdt+83xzy2w5bXWfjCzP6K5lk7Q7cb
v9xedhgGVu1R69nrGNCOBCqZX6XurmQio6bxpxWhBM66kE6+BK/qi5TjEo6E
2D3UuM/UXwj4mUM9wcggx+qVhhc9BSD+yQW7CbUaCS97nugnnMKFapeFfK6+
k/Waw3IwaIXRkpJ3LYxJBAiiiiuZ3Zk2M2vVpbN4PF+L7CVaKslYUzP6OJRL
hV4sBd1qmVF3QanXEjSohwEJls6pDmK3qKgy+BtT10Zqn4VVYhUiCJMSL3/q
TuLrC0L5d0rJI7twofz20/xSK3dl4igWkr9N/GxvZteCO7lPZkEZWu5NMz+M
4ak7jEOSsNLfHnhMHa9KZQu/GHWVf7CQqjnYbNa3TfkP+JndVge11UGf+aCJ
agwvwNqcd6KwGiNEAUAHJsEmLo5EumAmB+AOP9Hc7gTLd9TuOZC6JB1Z34+R
rGfP3eUujlDAFTGBgzwa1pYiyT/Jn2ZMmAKw0r8Do1FFOZFm7eE4JP9UpyMU
0zDLOLsn4IQy99fhTN4Tc6x2pS4llzwRKSf+dDmgQ0YO3PzgSiCmUhtsFxQm
UdloyMDguyDAMv2YXLByyeu0fdNaeTMgNlTLHE6fb5yNQ9EpqdGunY1xC+oo
jJQY3YMmKU6YtDPhlNND3q/7fsOlC823F0LMNwnmOLpk57rxHnELLpPS6uSS
IVmP7wUC8Ls1Jja8kqgRVdFWYJiKJcotTG26Gkbr3+ywCnDPJus/YtVgZkeG
iHfCDyqfctRUNxwZIg23LLqljseI9KIq97I4Kms/DclUh0suR/eNSvku6HvW
z3gtyquDcbV4RSqyGkWkCL7wZpkDMXyzurmdcD+KDb07CjVpzXh3VyaEA195
/8vyAZxRNO6BqH4A/zy/wS1gkhlSTviZDND8yoy7d8HPRdjMO+H4d0QT7K8G
FP32gpvm1qk/bwbLJEjCyuaqGuI+rb7LVJSffjsIXBwHzxIjrN31mWjeEsMt
F9IdK8aroABj6OjIsFscFl+xqzHHusYDF/xmovcGmxMD/OrcDLmWuZuuDw34
YhcAmMmWWvmwaNp0oYknl30w+qdw12dWixfDsDkEyqxMQ5omIJcxtLkopcpC
8T0qKrvgAcekazrhT4sqX1CyEJbwRcbej/4IK8tzyT2V0X7GttP/RCVRpOpP
bR5cb6eQcEgqgGeTDs9R3kYw4xBk0LE/CUJtPm5QrLx92cx+8cmEQLg6TU1Y
38zY1XRO1me94Pb+4yHlgFz8sXZNHNIM94sk53Imjggqs87ASpYAQsG68/pU
Cc6dwmmEJ1I2GC+S9hIXs82ALJt1xOevuk07rfVjHpedAsmFcfwIPip4VLFM
5um5fxPa8M8vlB0r89rk0JMGXPr0mzTHp/wshMHxzHfbGM8abUurJaFuwZNE
jaiprEjBZtzVIE0SG8SaXNzHfJAwAiM48pFkAnnNMVBevsrRRxivwMlwP45s
r+PBUXxoXDUqC2CMx2wzSA7QttrPOYFJZrd2SqPKkvw27Ox8kRwNqk6OU94o
3V1dNqxXfa8ZcuMNYMl1rop4+UFz6lSLoTRi5XqZ/2/6xqVK5WEuKzesNYJg
740HCjQsQ/9X2tmzxeMljLzknw7yVF63NxNh5+9QGo5Vssg1LxIUILITxqtn
DDfK+ogVkZ6QYmBzJUcAh/XA3QgQ+mFpXrtc7MRbWS1sn2uSMqpjlNxm5iCe
/DgBj44CzX3lRvOe4/zOrUAOBDlhdBNSn2j0xMVjHn7NPtYYkjmO0a5dQ+f5
/KXCeM5UX1rV4W/2zDscOM+qOGdJQaakxkQM+7D9t9AAZm7sIISeI3q2vH9R
TIM1HuRNzioKjx08XW0kuCeHjYmR/3cQl/KaYC+vJZwrCX0hfkWj+yIbBJMF
Zf8erD0LpaWELa+lWrEAcsM7hCvrdQX7XCsoQE3Sa7R6uf0cCfODA68npe13
n7yWUOJA4ZUKEKuxDx/e7ePy5SEYw7keyE7VUzcHIVm0gRvKRJc2eF0xM4CY
TSr/IFxN9GpRwfE1N1FUpGCoVGSjhqszKA8WXLpPbDtyfpZUVjd5C1Wwyo/D
juzwumTOOLj1BDKb7q3lNknRTYslY+qjDox6Fo9TISLv+gSE47yxKQyZ9qZ+
Enz2lieW1+/KPWkwC/hIflYUfhqkldOYm2FnvXl16mgKLDY26mcfwDfcQGFs
3AkNrSdNuEp0VUYE4zFO7+Em8qicUyv6Oqr7I7YDH42iy0NncablTWMi70Oa
HSpmXi08uBTnRRYmqX3Sye8hP9FdmbGEeHDAGd/ASE5RKRyc01WHpktDAaas
ZaAVgDs3o0O/hrC3wPL0mkp0gES4ZxDLG/dOeI1qti1XZ2j5hmdR6379rpdc
BaFGr0a4METwsKf1A2W8wArYg7DeztWRT/WKOaBoYiYTufDvwsJ6WeYlvkcP
4C9MIRuTEOTJkc1P3bnwVVOxD2OHaKSJ9qRX8NK2Ud2Zv1UcuovSLm/mUj8X
Yh91ec03POK6sfoJ01vmoGDLdUNgMU3EBB5yOI742syM5DJi5s1p+CHgjZUV
o2MwvFgWz/x9I40dvNv76ngtMTcnbFYO1GphMm45lXw4n79FWyyOQREXxWtD
HGmdcUC/HYfY4Jmyuls5Cov5rb03NqXCWG53aIJofyN6rsn4CRPeIDkznce3
OBiZo1cEZAcsYam7fGMN0yXI+QEkdDqT3X+hW/OcwqXLxkoAyd060mNTU+oR
4Xuj4SY8ZMkLTqZR1axXWDeW15yjg7mEZE41Gy1jYJIXonrRcrPKYho3dO11
1uIrcU+LpuDHJB6hlCJuAo9yP04dw+mrR0pjqA1XjSusmDts8sw5iwj2Oxff
b/aqVER4s8gN33GJRSScltuotdvyFWXu+EISfJ2jRLeyF17sNtbiG9K56uVz
SYgULqWl9mZNVw2RHmwZ9CFWCTj3OyqHNuCjvnezph5WSLhehbJk7g9G+qBv
0CITyZskk8magGh1/tAwvuRfRIU3ZuulFKPQUVslsZVcaZHSXhR55z/C1l6t
Z1pVc9y+nNDPIwC7uXOXqbzCbdg1mu5X/RrFYqXfa/JUQUMRzlU9unouwuzO
sqFyPLjgjR2L50Iew9rqZ5oEGdpiU8Lmka9lbACciSDNJZpDLyuQcDnVtcHm
QxNLByzAIDgn2EGCUNXsaraQB5pnoc27B4rT+7PKZ74jjMKEbmG80dBYt7EE
liK6p3He4yU/eDcu9e3aaX3AvY9v8q6QZciYi38fnkrrzMLZZqaj+gPCPKcK
zopgETj9XvroMjGLFNSGQD2PUp27ldXFrZ9X3vaXAFkWDIEBZxMun2XHVwr6
XZYY/5ySM0nJ1m05eksLdiFPqoQ0uOPhkCRjYaAnO+Np22wB3Z89RkYrpHec
Q62UOSoM2Tc/+ovtHS9k5onBH8vTsU/Qa1VBDsZTkCVpuXlSmxcuD7UDDmsv
LPOSzQQ0xdzWquc0fspHizf8qNSsHuacwH+ouhycUj3zfmMrrpw6r/rV8r9r
P49XtiVK4mXW023mkewxAAXh4vGCqJp2z6tpbJ5HU7qw2jcdq3fDHcEKAQuA
fCb66RfkFlswhZSokfcuYSkMJ2SQSX53NTtwRF/DEMbRI06X/f+olYY6Ta1G
RFkcqxsYLQaULHfivQvsWmaqZRlWIm76zS/nFJpMVv3x8M46fF1ELfZO6BgZ
n3C/71JnJtlFsziQdDHOqvrEvlKriDKIy5wzvAkuhwkchJ0AMw7UhY+Zzz+o
+6OIkfuKVGgZMMB9SALr6+8r0HIRq1fXdFMxkpgZrJMlb5yY8s/wj3AKZftm
gKIXAauRtknA9gZMpIAsiSwZgVtOlfOpQ4xDLkcJAwLSyfDswe2ayq9oIs/g
q32uCrh04PpJjzfka28+Du5HoHDZQCgDODk3/uNGkWKt8EpX0CBWJ1L0lysA
RVfPrJVWy3KzKiUittbV4RKd3m73T6tZ8KU8916wg6oxAubU/YkgVtwsMwJ/
cE9k1DdVrxZpeCi27BBI7+sqr4PMkbj4tiKnEz37EJ5JzzXVAY2RHq8xkQKo
lUM67/bXKLc/yhhC6Z8Hn+lTbHMNGyk8nB6VmAWB3OAabZhBG9S+RJm5RuYl
QeP4nvHUMcFom5PSGMp0y10ZdTrZFTrfXxYlH8r8CjqTwBEcAloDMhdGcw5m
lw6z7V3MYmCTcakWwPVT4gLp/UElNLJnaBjQajoUh4sztvUhoZ3PlWcjzZzS
r9CB9ftzUUOTdid6f0Hqr6bWbos0RNeETQN0AouC0Y/B0k9j7GNNptC+W9XF
6OmSWeV6k/i3YVcvyE8R24tLhsYVeQ5Z+snrk1PgGi2J0U4ipkN1d8JzbGb+
XYnJPUSBAu4cSKi/Fejzl+ACC1O/o4KYStvPVTbs9q05KEfHrqdZt374jYxv
Rx90rOZQM7fT4oX/5LxkHN6eVMRW22ewavmJx4LUBUUvMGPyhdYiW09nee59
1jX5MUMy5nKZSdPKtve5emMgY/DoNrXV+8/4OCmJ8CvaVH+8TVSbszI1MYtX
zS07Izjo3DELvgIq6Hh5svdktKw7U9Y3fp9QOBbmbwJPqvbsdAYwaop9wLs0
U3SAzkdSwKU2W010I7S1gnVtq6EOZPRV8+ljANcYCFA6zna8r7KiBeQT8RcX
u61XTcBnupjLavK13e5XZ0y/GFxCvcLgU8NRB9XfyelrWea0VQa0DLFQn2UU
FfvUNwSjxaAVA4Uv9+7+fXIXJfnLPa2Ann+LPC63ZhVj2fju7Ut3hAbTnKCK
iJVQ9waYGdsdPmbF5XbQjns9m4pjwp16lyiQ2a+Rwyjrjnj0fhVCV2ibOi9K
jA5AKG7bo0zkuG9UiGsxHtsnM5CLk7VfnRmu6J4tQUh1C5RkH30awlfQOMaF
S9f5TuBTJF3l4LowPVL6pIZeU6qbMZpKmO/n3beR2zZstggWdg2f5WNjvy+b
4d/WeyuUVGj3QlUhgl0F9dCOh2bR3mVM17yewp5mNwPxr0Cyo4YG9ojAPHj7
k0me/uMvgD+3FmKU46c4bPlERjYVXbyy48wYyMW9vQMYANZUZlZD/l9JP4Ma
8nQmjfM3YiF0JYeLSMbqfdPB8cc0DB1LdarZbroJWfqkkvHGbplj90/3wQCY
6dLWaMQd0P3r3rsBrgtDf2kFACDHG9/AtUqQGFj8myntDq14UAkduVPncxKY
8QgY1HHgOtJJ4K0LTW197ynYp8ikjBdSnKpP5plbxse+bGKjGgNd4px2IcmX
cyrqV+5uwJ1x98A0PF93GKJ4z9p11T35BcoF7fuEjc5OMaf7wFS3E1R+a+03
+iO468D4LBSVQUVygzqittjFk9X2liTwc4F/+7+V40KQMZh2oaYd7M4+D4ru
QMVidWfj7pabF99xDUOOvCLRMJmTenUyEV/GpHY766f0hb5K/4OW9v5otAnD
Vfn0/j1Yb3oqaK9gpksqh8B5YN8KNcXyQJxOu+aZwMNb0Wcf29vusQxUlWtf
FXZ7HhHnmuC4nHuMIwpmffczw3WSfFYSKRA/OlNtp4xo+6n1gE4yoioB2Exj
JIhj95GTNkfw6EXO3vO/T/EDUf6TqI78TGNX8fki2vQ0iMxndVXWZ3HK8HSo
koi9gUmpWGq8/rGA+xYAX8vtlsIl9FhXnqMoeN2w1XdiI9KK5HSOAG4oeHhI
YhYOk1FIAe6LN1JTEiHKlffAoiXkpuubJAjyYgg/wZDot7fDCMLkVFAXxEoh
kkfjJ8d6Zx2ZgOPE43GQZKWB9TZ42tknFzOj9ttfRnncSk+t+uGvvUJcmixa
Kj2p2/kPN5U/cZIb3eNUxtFGzYSd2RCT6iyQmBOdLoDHA1l262ihu0aHrH/e
geEcIJ0JBzS6HxKD1Pj+R9olw60wVMXMCRxAxWFbhfDu6mA3gMoYBG/1QPgo
En57UeQTdDzuSOgZQjE6u6Nq5lgKYK6A9ZYJKxg1QIJWmIskvp+E4tughR0i
Bo12ywvbgCCr9Kmd8Uj7M7bRDIHYgHHxxeN7ZEkc6II2iFs0L+EpBRMWSxPK
7gjlO6RholQ/ulFU805FkaXXXBt0/HOJFAk1LS5zzGKCt3G2+Whlm6SdLCQp
NsTn4zZzjalf9EUh7PGxpm24PX+0h7xSH0Rn+73RMPGHdjfFRl7D5Y1Y4qeq
e0WTGLWUR1FThyOfspztq01Ot6LUGpHAVJSblPJva2Jt+U1W0K75cMrF19iF
QHxMLYLsSlMuGoiOt1vKH230oLA5hmL3T6CUi7TQKl2shZ4xtfw5dBc4hLbE
BRC3IPB9YRvDnhEUOnSr3hb+WJ8VCg4hvIILhJRyadHr4DMBDSoHdSAq32N5
xKEGHhLZXFpfbo40bumNOAyhiuNQruzS/YfmgKIPJ+kJInZw6iQj7d/eGNq7
w3wk33iifwjDXzCC0NW8tXoHC7yPQqeGe0m5CRkwskq2CiTeAGt2wUCG4jmu
bvsDtQwAYUK0en0uA+9HWI/6Pw69LcMC6hksVhZNLas9LiemNqyWZSTd6qoi
KToeP3JN6zmR2IGMus4QkcUpz2bpmfK6TSoQj8khbC2431YmUpvL4WCG2Zv8
JICZgS0iTnBD3ikGad+1lOhNDACkY8OhrjSmgyif9K7i7ENYW+01bAsln4gH
F9pcFmz47C4vftgyusaIH4TciOTCGF1fl+xYIksi7IGd9TFfvC1py5HCzQIR
q7j6FNmYr9MUGZSvoE/gO/js0kmEf3W69LlayaQhCVGF3jyJc3d8dZXPuVjQ
9hkBQNPJBSphV9TdxGrQvYmn3P7Xt1cSH55H1iaC3XBnoWCPtdeIUmR5sA2j
LBDCufdfuDSfzxC3w7aQwO57TwgYTTyGmE8HDH0jkj6DDcVlOf0wJprDqOBN
nOKkism4asU7KoUvIt1euAm+BacIjrDjzc3Fsfnby4QiHMcIZ0SA1p6e2qel
EGVcedrYUx475jgLCVBDanmhDCZEA9eckFyBAiLUCOHOsPm1IViExTQXavA+
h4DsvXg77I9NafBO8DQ5GYaStjk8Iv6Gz9NMB5n3z5jonzXe5t0/gcMCXO9R
H2kg34BIBXwjHeAAEAnd56X8w/9ZOuSDME1IU6OORJRXra5WZbg1dFjgqIa0
WnKMdb6ImvznjkaTDzT9N3zIsp0Z88DYQM1gO+W1SYH3MsXoL8Z42xWKa9b2
NcmuUJ13viDIMADshUkTMWd2pbplU1zD1b6EEdRSoi6Ogch+I7974OnxFAlC
lHJ2tUFbml7SQccq7fi18XqV9sVb+oc6M81BkyYAAhh9XkmsBjBZfczN7aaH
bK5f/MBnUu3PKOIrj0RQ+bnUecI2GCx4vPk/G1ESBn/XJGeNkq4fjssLy6Cq
YSyBJrBqGslzh828kbfXzCOAfftRsIeFnTGi+SUpKg0he70hdX78x/ZXLyTp
gH+XhRTddrLk8uGbhSXRYJdDOgPu329Tnirpc58/dSGtux9ZNcHhQS1JxMeO
lgnbUcOt9uGqsCHHzF2vIAOQfpYmdC9ZwdRxFdJfu8TxaV0IX+GpSyK9BgpS
3g725yZ1vrA62+pjLEyN2Ae3nRLXbRIWi4YIoVxKF4sdn6xXi0h9U3X3c83T
9QtxDDA0W30FmBfce33HjJ6YgPhGR3UtY1bijH0aS0PuPq9FBHz/BKE/8UpS
ealxJdbrlVvy6bc64aRlTGSUalLquLYY4KbG66Gyk3YD08QnuxaafA9sDD/q
rhvPLcUYtXuqMMq9ufwjJ8xZ/lJC2cLGaqBn5YiNcWcNNpt2r3+GZp0JpWn8
NrD5p/dK/ZtKKkFVbSXgl+6crvS/Pemp7h9VVMdvvKv/SXg52Npy2VAH+GsG
xRKr1YRjcBJKPUHem9OaM+Qqpt+K337n02XTNAMaPORnBFHTLLXbDY8FC6s2
u4XSfmoxfj6LGZii1ouvolBMnaSYxJxJ7VHAplFkwHrJqBrHWHdQgE418TB8
jDJVpY25z27ZGshNc5gIEmjZDpzWCNXcb/pBSBgW46/zTIr39RcWM2gsFtZz
wf4CBPAHT7dVwTTkdCTJgQkhamUQcRnnUYkddXqmUDeQ7dJWaru8YKMlrI6L
ECJ9luxDrxIUVzIpP53+xSiETVUCtC6E0ahKGyVpb26nnYmYP1LEQ0aKitWV
qEqWvJCthQFXE42NgEQjObrTAoUGa4KwJ6XAG+oD8kBkglwjc5XlORL83rJ5
tezqYiJPqDFAhEq6i6fVnJpRQsbKSuza/lbMYjk4l0ywCFzGqL0GVFCKg1rm
fDOA66JpYZTh/e7VdpG0eoZZIuze/2zXYoMoNdnF2xeJvX2Haoeo/kD7FNbO
mn8Nwqf0FAwTY1WDM6ngqZB1dQ9vitf1jOrT6HChKMFkdYbmn7cOInJjKrZd
VZOKFhdh3rvCe/KuI3XGdcKd/do5zDOwwVrFgtZI389WogYA9JFVVZtfFuM+
X3YgL6HX8j9lAQKY03hpvBH3ME4+LAb1/hBRWpXpWyKhj7D9AVhwVl541MkK
MPZFoZC9ZIsu5mrfGuMiudd/4AgAZ/h7fHIBEq+0zkeatC+TeMq8RUULLYpv
RivmYYGOsattOh4KywEBHwYU8wevO2zVhMhxgvH4DOAmB4EtJc04VguEu7q5
tZmYZu20LL7enUbyjtbiMcWdSImIEL20OUMaP/cTorwaJ5ZAj4HRVyACRYLX
O9VRNYCHh3CZS+9NA5XiSoPbZww31P69BROy0RNHrCMGpLU1N7bpdXFRxo1V
PoVvHXcdXQkqoeyoQ75gHxkLNRlwg+YnwYdFMh0zcrfJIABUX1Pa1nTKqbBW
5GEh/2TQpQlPrnEIN39DGHvayl0y9KCGBodm7SU9DfX/viYUMcQTmWkSuK6+
Hd0dtFYrcyWlGvS9WU6D1jAcq2OIiI0hn6hoGu/ecRH/XJke15j47HSn5cOf
SYOPOzPpc7D5R/DVmrUpPdXleM2CtLezyfEdzCgmATE8eiYUrR0FEey3n41E
1L2f1f8e8+5DNtmJEaPy5ldEDtxSxnR1IkGEHRPQVrws6h7J7bNCVWCWMgFd
RH7YJ1elzLHRO+apNKjJlE8WY6yBpg9zJIxzfAOgbHVwEZ4XDq607ZE3vV1J
bA0gzPiZKlw0dJ9C8G57exfn2pd5iEJe9SavU3HqQOjEyVtam7zJ3kAl3JoC
soPi+0HFokw2rBdOprg7xZixNYTirSt7+Ymig7EUZJ7pGpkmSnfpSP4Y2J8z
xr4h9RIH1I2dMURTCh/bzzz1eXw1wlTs32nAQIzMKaoh8ijU3MuVVeuHu7b1
J9VzEgIpaufIQ+SPKNziqOaYbEw9cF9bbTH2GEEm25fOH6i6C6n95K3F+q0c
KraV0UzURsq0t3r/ruHY+j1+wkCOe/nR6Z+q9hC5r0sPAF3CdzzsgWmpax6z
S/iHpv0N/oAhpPj2/Hdxr7k770QbdGVDvSspr5UVRaMszGTFmTzSXuoSNIJR
l0gpYeWN1btRm/Kq7je2pSt5wfS/m+/Q2Stu0JTFb47Z4mJSvmgb9Z43krLt
ycht29oOXoB00RimVnnUTXd5+UH//nNF2ytkPbSVvaUXh8L8anXwFtEH//Pq
/LA2lcCtFUvwYryNXSKlly0aDubur9Kk4kIwBCCw1a2cV0RYIFxWPqnGut1t
kcHLmtg9DTXHViVvBEQly5pyaFxlS4+xRtibHy0fC8sXJlzEO5Iow270jFXf
MmipyL1C+rGp8pbPRVFRGUHg/rv4m2oWMF+E/HybgEy2XvvQrWs6dIYycTpQ
gRT1GaycYVb0dA4T+1Bjz3ppVUKaXePy4PxdjH8d/Ugm7j2TxbtWKk5HegYm
XRt7kLgz34PLhZWY2JlRt1Mn5y5i9FAWqT1lrvg1qRNQO7D7tbSR5Kr1HLKY
63xirQyiN6Ib70sSQtQlF+aOdnxJ4JGCxJMGoiPqo0DHjqxBPa7ezEh5e/bj
kHyJDLuCWWLL/H2uekomvVc2vdMw4KOanwdU1axXNClPGE4eWC0DwAbRaKFq
6KQcLx2wWtVj5mQOviOoP9bC+mWN2nHJyCItqfVw8Oe2lHTAU9FDXDkRVP+y
+u97fVhR2a5J0vrZYspRQuJrd6gcvJ3uUu39lBsAN8Di43Gjk01Vwb2NAjBe
pyMZ3XrzjKJQ+aPYDlXMJk8j75dKwUpn8z7/KgwUDbEegDy2uAgM/o3bcEIJ
KCpfvJMGDdJuyj0z8TaKblINapFLi8fV27RujYO0eCj/Wa4JET+5r3srfVII
xT40956yiwg3fPr/6shY7MrRzmPkHNynFpf9vMO7eXHlqX/zrTbQmSWyT3gZ
Cr2cud2Wid6Fo8h5g/bE4UMy6CRcfqqn+4bXei0/B48OO+YbVBUKHT2KBz56
Ag/Gc7DygYcO5IjlTjcPA5QwnISPTVFFnkr3+ijJmy8YsJtmBYqfDN4Afgnv
kzDTuAuhHddNq7Blvz6DIT5Rl7gcYDaz5V1v8YAUcvWRdHNvb6/tA29AYZl9
K4olh4unqy7Hq1K2XXu2P3fD5GLqUzyKUjwL2izSKJkAxWFOq31/l2xPtK4W
GzGvLATevvxrkxKNQplQRudObQx7BrCU9Gtev0fqakqvX+DUWxk5wqMB2lz1
BIxp6L/+UlDqeFbKy7dRPo/mfmrRxAdz+3TPkB/FDOx84H091Vpe71JasnRG
pc2Sq29cxGm+St8VCiCVxWDzLmIJn9jW0AUW7h5jYcozlXUgR/z1XO7AC4FM
U+N2haYRRtqQclkV+Zu3mW5zs89bEa1LwTJNlQ2vQLvawYoKZuBGQLHoCgyf
20nUfZf1dx1W6QjNZi9E5ZRUU7zAKotPtJJaXAgj7IN0WjsrjZpZ7yzJRmmK
Zilqpv3qWkZcVas3f8raqjJPaI/QiO+SiuLho3asDLpJVpXWMKT0jmkZE1Ko
N/0BS832Ban1XZ0SjlRdz0vVwBVYsDrREyPwoTec3lycqv9Gm/7tWdjhP9xE
M6K9yZKuFriJN9rf/3Szw2EbfvAH4lq8bKev/QjSxjc2Q4pB3jJPQlyUOKPm
2qJt6QzLDLH5vKARHeW/Mz5jSo3inrKSZJ0ZMRlN8plUlQfEwtYuF4+puQju
nRqcHPYusrGECa7wpX246Af427/kgRJUHHiGzbS/byAKrmbvYmaABM5SfG2y
Tw1FnTNSf29OgJmhzkEORrPaRN6B3eUbB2H2Rvnj5upINnQcvMMJThxYjdkL
WrOkYSboZvD7zdeuNm4ceEqifpLtRTSYveBKXwaWYr9dxwndcWujMxy8PrYJ
7A5+URyLaWxUfydXOIKspVd4MYM5WDdiPJ1IFFCnp60eDYOve47UvRQ4TvBS
Y5pp1CmpAFU1Ku7SiZB+m+LzuNzDTinT5zeASSHWV2ZoWsQvNQQqV7ruU8gR
pBF03ZSmRRCsbIJQ/6BptkJxAddRSlsUN2L8VY5kjSJDKWcNTW5fApfY1E9v
3sp2V13KOGH/6h45JoNyL7y764kwoJsLmsKFwlOGUOTbQ3lT/omegwntUSF2
qrWEgcgzNzm9xL0+7/4hnkc/MyMHPQz9LL5E0XqzpykIwFF9sagF0Wi5rOgl
Qs2c1PlJaFcCtIfQQq1lRjB+ppHCEspbMV/uBKrmvVSEYrd5mBlSAiBg9SQs
w4pTs6p+qLr7RfCUg9kOdMnHZ+JgCt8e2khxnflu1T4+43VfMSw2ehi/vomb
/z+VRPohMOfImxvDf1u7BTU27Qyo2P2y0M+LFJFMgNDGf/qPkTfZzjdnJpz2
yiE+HyxE9vm2Fwn/mPT948+eyTjSrrqmnnhunlPGeFX4pAMfM0GW1tTIQK0S
JYZSylEN3Jv4YmYvMdtR9mpW0Xhw/UdtsR3UOiEkEyH0MDReLTqaKfVtzJDq
OJiBzGZkCS22JJlD0uPitaRZs980OReuu/ZhPZnvv3XAavpjJJjSX8XhTrUX
pMIDpv5erTmhTlY1AI+0lsuLArqdgSGWHHEvYLOvwefkaNWjrGR2ouy+ucIx
vqg/u4WCcABCv0jM0QCZBsfHnZY2H2aFJjdZnxdlHz08tKKU+9Oxy21KpKyd
XGN83donNFCPQLyMsA5K54VdiCO5PG7JEL6f2LM9JPUHqRyiCK+noLy4aW6b
OcvSxAy4EBFghYtNAWfhUZ3Nks+F9uwQKhSppFhpyrqW7BQtyb1K/wRTv96f
eV/mhIkCl6JWeIBIiZoWEqOlFXNSSR/BeiFFpT6Ecru0G3IFUd+WDOMixmwa
p/A/iRDzJ99m7QQZmG2YTtzKIbj1jMdExnidLTM9ikPCX3xPBpDgMBj4M0Go
ppYzYB1XIyqSkL6IAY9bzK4tSATljfURKDwB9xq59UmIXHpg40msL/9segpd
AsnnSaCeyagJlkNbjBq33t5GiRp4vgqgXVAd6ZRigfoeCUk2HZuM8A9CsUBM
GcoKBmOM5tCEWvjJA7mMRI9Tybhf19mEm3d8zWxSD5ZDmsL/H3gheRz0162q
NhSRUwVRawiD7CZopXsCxayVsBXR/sWnI2ooIxwultnVDQ7w0vsgvyXOK/DU
kJx0dJ7PST+YPEPyWZ+kUvl2Ww457QPPY7f3EG9TSVZYgWhLWKJM+oL/iOgq
bMKjtmWcAthu1M06hzEFFuoJ+2/y78FXdieM1QJmpCC14ASaP7OuJj824iIv
/5lLyITahmyjNuIophvqoG9TEQoRVmT1zKUQmjkwH1y72AmzvBpjp7+2Z/Mx
eBPjIJrluLEnDFks0jaUdJJogOBvyy2/EcUoXPfonvuKO/6wLFjQ/L3FPTqI
BjTvvodR9Hsb8w4hVh5Xy1BUUg7PPxLPDs3saqBu/Cik5UQS3PJVYsX86nO/
AaqxfmKO0tJtwTJg1bUAU52gYQneLSfnO+GaRBti3g/L587WY9LtiC05ttEY
M7UtDVjCyD7eYCPsfw4T9O5HetJYSpq7uYBKA8f5+FH0I+Pkl/Psu9RGRqXS
wl4ZtfpPNuiquFhilbGDtVA4CRi14swQiW7exRJI5CyNi/qOGX/PCLGlH8nv
gHJM1HY33is4OBQ6HqOcbfsCiWxRxOgs9ePpvccbjx2G9xl8D4BVRAvTWGfO
iE1O26XRHhsYrQMV60kruebkpgZoO5wNr0Wf+6mvhk22GJLvWjtCIZbh7pCI
niAg1W9lV04oJ3bg/WYzMD0wMfiiTEg6sBGa9U/5BaSKSzkU/1+u6sYQnH+R
FvN45N0ur6nFPzGjPa9NgYmC6EdWMZNM+dFvEnC6q4quHnhUyr2UNCaowtj+
Cyg2y5ySg6z6cpC6M6Z2l41aWh466pJ+yhzi/xPnyxB9i8S14Ig7XQIhd1BY
v50OOTYkEgP5XwciLOfbb5IewSdCbIjsd9Ii4/4zAlMUAYMQ74WHe4Xl7l7Z
5s+vd12+ECJDPQxqcwdyJeRu7qOejIe2WZHo3S1Ambj9gRjEILQS+gSJlCCF
QIFbggdkTOhEXcnqmAD0UgBFbMs6ErLWFf6aCnYQ5p6QQCEvrk5NcLUOga2h
acrKB40c2aOqRMTiLUh0A4CISG5esOZLVZ2apDNpqNA1yt+FI6FRpuH0EGoI
T4xwIMrFoxSqDdX/auarhjtYU/idiFxJE1bICGfRciwOVV/gho3FkqWq5LYP
GHB0cOMsdPLQ0OAbZYnuby/eBtTBVcMXgVwSxcLDso+iQAFZdY0Evh5M55dn
6Lf27v9U3TAj4fgv/DKznhehXtrbBdvL9n+YfEWV94UAqbTW4/JWc5iOacp3
NQzASDDFjZ/UzFFkSSEbh4r/N8o8n2etJPjFyHRqPAVPAPJP5mVuNxr54ZSE
J7qIbF0V/snAHLCfrFhHuZEFo8oCDpR776yXmKSJRpLE9aE/jAWcfDEHRDbg
1NVvOQPDNWxJP9DiVs9v/OvgQKoymJHNy24EFr2HiX7RdEgPTll6YmVDEIUe
FrrAZgHMjGk86T69ExmMOWFnDf7n3ESdsCKH/WXvHvhAW6CHR6kv80/9km0n
str81I7N33ucdte3TSz/y+TcMIFsqmACFXJm7IahvyJFUEWGaNaIoeTqNYaS
vbMYERQal4yQDntp2MpO8EcBYfJaAZiFBhncHBc+h2bzsuq6s6VGitrQDW0t
j1/0DXD+RweManwZQC+CoEcZzpjhD+rz6OZCsVdPpWnf0MP7mqMOKThhrNhd
n+g+fWOF8oCXs5PoqpySqkTWYbmfEQmwW1kwJnrWhY3XmIdtA2Kw1OiJolg3
PKUDsYcymli0hbzuGsA434yYXGd4DvPa60W6/ERfJ4klBzYs8T360Lo11rK8
o/9DrEzzQmz7xtVL++VID7T88T0JCwwVUYA2439u9bR37JAKbm30NS6d0B7X
A+8kER+jV9EkMv7Kf+M2juyDtOEndJUF7zsbgKD+FY6lrSUm29USTemAEAFP
kVhNqRG8QBd0+vg9dQLLnMmhLnD0AyttXb6gXV3DWm9tQ942s8DftQYLRHRq
ZvU9yPoSHqIWh80Hhi25gRhYZTRFIDBRsI2bHxaE7Dzbw/OYb1hzrx0sdeWy
QZMnHEpNMM49vfwVfMANmD2ZVYdlx1ajK5d6JyaLG45ddqQ7BPClWu/0ZexC
uIacJFu/984Ttrv82bOCXyXYDu/DzTFKlLoYRWyT/cQS4dkuc4oNTF9IcsNC
gH/ynm4uU4zlikRQJCL1uSLq3RetKvvvEymNsA3AEEHbLH1gxiTWi60h0YNI
tb9tycembRWIwDTDM6yrr4nVcDJH9XrNj+BF1qhw9g9/29XA4NI23UljbFv2
PuCj4GOZElf4iDepZevktrJ+wIcLr2BLPBd11C1xuIXWB0UDI1isIrxQKMtA
sFkW+otSduStiubpmVmVd+v6eMMCBZsKMI9LIjJzwcCXVkmLbfL2uZ/74/bO
BPUOovpYRMIDS8aGgZisWa3crrRWi/HTYu4CvhmAqu9pKVjxFYXvx6Y//Fbp
hhLq85XZi2PQ50wHxLw6Q2BXyGRv56Xm81LXV+XA+65U/6g7PbfhJDag39zb
td4BbYir+dUffUYhZd+uTK02a0LQSMItBn8aJsabXOzspSJpl5supuXY5Uus
ug+PdndYlQNXDorUJbJLenM5KUgvWXpo0JN7JCrOFEu7M7l0Q9INtQRl4m96
2HyomRWzjj5fAookbK/FQurPQ3afm9d5AScaMxc9S8OyNb4q4ui1aNP/eiOB
j56J8/unzTZJWcN704zKMArvun8KsxFMdodVed8qITRVgJbbGWBc+3hozscB
6SMSQApTTD/b1bSuoKWlGyVd2443EhGdxzFaJcElXxTWXU+EjT2EoK6sWfUS
yMOzCIlcJEOv3vh2ujJ+XYRsW62pJ+hUW3WkNMUlRWe5qCvjhgNfXEYfWahq
6z5GtLe5mHEhDJTazzPaM79wuxR3rT6xo+9bJUifWIPPivP1Lc1+qcGFLYW3
Eg6KnZeu65pGP1k8+iMKtxlgrY4f60MhZe3PgD3ZHJBacLLtzHI6kRtNUbpI
9oKHEDsF2c12xY6q9bUTWyT4XBAiHmnQkhFfIEdSdm89cxEk/pPNATQsDIpp
5g9FBJ3w5bdg8NwMTQjsVMCIO9NPu2WyBH+ghngaH4RgvTy90bhds8abzG+4
aYC4zpwF6XzRicYnV546TyhBWvE2IHbBb2WJNJgavIAHUEk34NOY0Yh86Fj8
GXHdGWptqTXrL9GuFCzVhdjEuv0Cu/TlRHlVVhoqMB/hIz2juD63BVaKa+ro
ZFru8XY1wXuShIp8xHcPGBW2rIpIKBUWLX68C7teZN8YqkI8l7ad75nEMMEW
lD7zCrylh4sWw/Ws7+14Gf/3spuPgVn38Xp3ebU7WbaICIHWKMM2rSfZlJ39
L61hx7OKpQuxFeGyCmbZ78j1cXwEcAA1uKKvCs4R9kSPZPfjDSDwATyxVZQF
VXUJdn9hR7HQwdKXg8ZM0Ufvd6Yi8EkKPObIb3uDs+xFhMd9Gytlw2Ih4F76
vlWyD4XFLM1MxXgwAV7IuOuzKCoiPKuunZ3KdFIAm/7qEdLo8jD3qkPb1Or3
a8jOVMhLiDl4jos5hkJDPxzb1PK/N/jTOkD1nApdXf5XFoudgySmJJQziXIH
yfwAiMEAU5f3LkPbIBRCtW/sHa3DzEz8nC1ne1OgJczD5H8PwwpMxLNt1f5s
ebWVVj3AzcK5RjjCK0Gfw7GpJnfzAekxu9GVdK/kbhnyQB53MRpLVKLU0YUe
zXM+wJRYt0mykYo45K1kJrKdlDs1Njim+SfdPjpEez/BTVAMl04Wz02uUnj7
l8wqlmxhntsh5zUNNA0Hyyfnh60jOh8c8NLXQjY6lfzWc7kzEv+tiuM3nSfg
EtKmiCbI2CZVQpS67LujxagetfG9xfXC6sjo3hXVIXsnv6wMSo9lTs7YBhVe
2JoAlUzCPZ1r3geoRmQ6bgM2v1AYH9+TDWDaa7mbsNprKXvohP67GfqF94WY
7qN+onD7Sd1sOsCg8coRCkQhwPAkxXcecO41YLJRACs3cMbt80BVvEL33waV
iJmKA61sDgZnBdSy0XwjewKaaJfBd3BTqUhqKnpRR4Xo8dTyOBIu6PGKfb1r
2AnAHyAOzmhPcch2g3tVvW+ER9qN1R07+SxvarzvSQbeBv2bfR7I7atb+J0c
pQDx34OYiTArZGP101rAmuOxUy9DA7bd/TzzsyMZ7FRm8NlxEb4KAbO9TNVI
w1cFWAr4qVxf8gAqCAvJo/Y/ZjIPrFnPxto0dIdKQao8rDfZ795W5jqrhFhH
AlEVcPC4gyVh0iRmEJBIbSYTrsJhE3m4BbKNPpg819E26DUgSaKVH9oC2BGT
sI7jVOxQoYILJH8wT2zcLbr//MTVzPiE5wMYpbI4fbpM5C6EqIsoZmvmZjDG
odbSuV5YoKfbPLxkXmDwEK5upLG+Sy0fXo26XDnGeW/DT+V71cMxa9qcRnAu
HOzUqUWwiuG6SPNO1qHg113jBf584bApQNgfl/hRDR7lG7T4m/+ugVM7708N
Tm+bA5I6DGQWJZSfhbbXD00cGd/qYzvSoo+r4d74Qlxmc1Z06FOhErYBoAhs
Vf6yhdnDv0QjsVKR75Ihcy5zrPi0BTH5I5oEPw3b1gcRIPz9+ldmOL10CZb4
iSsZu2dsiz1giGybtxetRf+DNRxU2XrSCitLqcZh9vtSLVl1Rb2GH9W1CA7X
xE0y515jCigV5aMb9xlQtgapDuw91OUhBJjm7fm94Rhz1ciHI0M05khKtgxL
E3zXAbXRsE51/QfqMjMxVzl9N2JS7G5hJkuLvhbu2gYCDJKIVQ3UXhCnfvBp
wS3pi88Tb892rLJ7+qmkz09VBbgkSGfG7WvPNhTxOR5EaJmifpq3TMShiRkC
sxYUhvo5XsuPH2SgIwcejuuzZzSoteh98kLMhFMMS++K7oxHD11ExDX3twm/
GX3dXQnHjA6n4XArN1Gjt+M5LkQ2V5wMDD4iliR1fAlIO2h9N936ehCSJv07
pn7L4mnhuzovw6IFSxyxeSA8snZ8VCcgA0QmHNv5OUOozp5sw6JETfMrn30Q
jdma9uZOS/NH/dj2/Z6/9o7CcWFr/jm2y/Jhlwn/MSy8Aw8YWGKCTlMZatt+
GNOLi/nh/GfSZr+65UQbcpifAeuoHSqvYIRO+pKMxxEy2/cgLdfVbCrAbMmx
dEBgk+LQu3GtjTXHpiF/cwOoN0JY9jNRH3gizGg56txz2arlMKTzkoCNOOQi
IVfLcpgdngaLK3p7Z6AWSSlOy4vKOulNWidTxUWdOoqB9vqQuwuDFc92wupX
mThg14ETqFfvP6Rr/g+WtHeudXAdzYySdiDw4qrlYncdWlVuZPpJlR59DwPY
WrcTLG35hDY5b0jQXULMFI+wF7S39kZREzY/wLwyDs0CMd7OKQH7l6S5Kt8/
fFruW8FTxWKogrFBWpzCGIqU59zvMAJ9SWJhy8nISJl4wSFX6WP812r6/dRi
Vt4BYsyZIR7oK1ljdKrEssZIRsuFv1S2VeQ0dpO/CLNgJk+IcswBaCzgriRx
uw8NwcZqT4fXeHpK9IKgXDj1OljOSHnHTOp6tYwmytZnQ7GWH19cz3rk1fCh
1TEiEYLrWjRprgkpfUKXmK87thdL0ugpC/wQ32tTUrhGa1IN00Vha9JXvCZK
IYKoPi8Jeptde+lZLKrqId6LcMjSb/IpRX5YJmSxsfioBS2ta53HcM8q/fY1
RNam2n2zOBou0hACA5ZS5NrdGdGpFanYZvdsbuQUEUWL0wCrDMaRZyKri6oZ
mzrtt+tPfN6JxOUoRtiAI4FCYAYLN7UpkdXokUdnnw7StVnW7Lny/rF7pCIU
w38/rIFqaE9tik6Ur7A/AQU+8y/6+DvHOFz/6AXpTG6g9y1JePLigFde3WkX
kziqlKO+rREDVcRom1lwEw+OW2DE80K5EL4nMiQDWP5oxyACxXApAgdvPvff
MP9+MCBtcs8sHP0ceyIvgFlgTucKzW11AOSnnWmIu1nUoxH+14vlZQvq8n0A
2I15e1GBCS0JULmRLWNFOW9mJTUIS73+Aorv13Jupbcc6csQfCIS8IvgrnGd
drkvgX2eTE8obkFFsGoeXcpK+uBYwNGxfY7YZD+z8OhRqz2110VuUhRHB1y5
XvtKBy2csEP/smTEBFnoTVM0zHM3wUn0YFMt7YKmszi611YCmBGRLi9roNPy
7TT+tppb4SvE40LlefI+3To80cl4+1FZZi1ergOamMD9Gw/nw8xZ1WZWn88v
0bTgY6ie58IKBLbNT0gM2ZsTuFS0m4ipXNnKOkaMear1x6V3H5exenxqucdZ
jUYbpZ4Wo78IIzLUYNdOB/s7ZeoRBfv+vyeBX+W3XgxVoC8kYiqN+llONgY4
ketu7tOPi9qn+UV5km9TlbF5M3Olv1v/v+g/mO0zHJFFoEtH5uXrRkbvXC18
TqkiCpZbAmjDPItQIhr7ORQLMv7lTlDhoxfxIqfZFwbry0h0wR8HHZzydlKq
UEfBPAj2rLULP/T3grvnRJfdL3Jg3hJAh+GIIP3+m+FduPm/fezLEXv30mNa
J0/MYT/m5G3yWSVRt5SSsjMRE1xQOpGcFJKr/WzSeJoY7nN3DQgi6MyyRcuu
jJMTJJa7KzSlT9gZr+MJLZqSJO75AkNv7+BU6EPqLhHeqrMhewxIdoaZiAw4
2lrV//btBiwScb9L1G03ApLyapSPc8ADEM/ydvQUVnfOWz7mT3QQQM2lfiQS
dWnx90NjNsBWMPAUjj2uamxFZ58WIteypGsHSawG88Dd8yw79ODRLzV/f5wp
70oXHuZ8hiEpOq7T5LgFEgI20HN7AGNXDgD4miSAeCB+X+i0Fvei1DxZQVNF
EAfh6NHVn0u53Gg+0/Nt0/oYAZYEl2p4l2hgYjGXheEHNOfHXINq/qEInFTW
9ZGzGT1jfSo1cKyvIlHfHQNB4HwRTOC5UUK1eKZiUTumBRgNhMHEkWjZkKBA
w05LjUVtsaZY4TzyEifTi+QoUbpUmIVR/Roqi62Qh5CAP8Q2tjBZKff7vSNx
5xbpOj1KkmOzouoifjZ4VbytJIGz7d9NZzGhTgobj7Q3Jif0/VsCDQTOAOxH
mFxJRch/q28974MXnQUfXyiloh8rkuyjxiKnD2ZyggRI9OIPlZWkEeXZX0EZ
fEhz7eO6s5p+/hOGlKUjOGaks7R6ZyKeCJlUT47tENqI111Zc/GTYrCubcYK
WUkRo1uBEFGHwFx5aERyT5qurNltFoHH6lPsL6kvByncBXyGDd7tX15zlqbp
HzcIPSar5gfbU43Hukv20JXNHk514JcjIqPpQ82kXFRYJ+WNc4VmJ8vXuW/c
wcP/AQBsxwi4epu76pDFxQ7H1rluSFYUNDwu2qean6p9CUN/BcofsuCtRFt7
zqtuZvYUV0tCsNPlHW7BmPlB4tN7GHkSRed1bqlibwLjs8+5cKw3BhfnV7TO
JGH35ivM8Rd783gq8wJ6uVwrz/dgUiZpBWFyYN77UAQWAwXHJEgFa/sp7Hq3
4XAnAmn8y+57gkuazeuRG/J9uGs9fgUtPnMyFNwYW2cTYMlMNQ9woIW5zNgn
L7+nhPiswZkvWKDGw9Gh8L57uxcWWJP0OCG/VokI7zpRGxia3Lw5eDIZYu0U
mbmU2Unx3X2/I25XsxBykkYLpLLM/PDUhhKHM4lq4EiikLqSO4CiTBuoLbQG
+f0NBgNFeJGlRuARQ+/itsrikFBV0CUCBcWeoZ161v9q9LBY8mt6mNbNIHdJ
tAv3MxfqlLX1RRqZHxoBN7XlppRfn+pz2d7EzSPF2kgfEkSi6TE9w53A6CjE
ovoNt/aFS2cDiyg03g5Reamv0/fGdJo4fyV2t9Q3HRJaS2TNQ79n+7lmOevw
1t2fu5nLSAevTqZZVdhm4rnmHsM5qPIq20RrlQdGwIjfZVmx2YyacSlbT6id
K7nMxBEjGSMBPwWvJjXX8Yfzjy9UrRlnBmDjCMWDnPfLky6uBv2YFumyF1jF
im3S0OnWBz1SUDVXj71aNn1Jpvsh+0Q4zs8RLpE+PWgANh7RLVngHTJWCBRS
A6x1vLVpJyMLhc6YT1LEDqb7KIdaAQP+8YsKsK0I/iYmbhJ2TFWm6ND/vO6h
/2X7SSJu+hmjgVOdELAZ99vFmCl/yify3BpLZ4klhqgTA7su+HPip3DUtioV
f2FmbGLNfE/gC4U/CORPjppn7SZ+hp+zl87Uk5+Uf+cWbOfzaoj/QBVwsL/m
qdcJ6+BYIFfudprKNno4/8Pqb1bV/fp/YhCOGQBUa6QBWHyQuTX+8IjKD9g1
NxBSafOpiFPYNH1W6krP4A9tSZXtznE6snrEHbqhmvdahegmrwhkhMZbISTB
SqbuyyM+TrLhrgNZyfGMzEXGCZbMWwIZxWvU/CDfWAS6ArQe9H/moprLsbp3
WNu2crldTo/q+g/OHvTd2iNz44cg7rfxeWFEJzKy2psJPGvBj1yY8cOp8ZoI
xrIDHNnVHPEReNsGdBnxfuIiJwYZmHk2Ll6NB/HXpfDSBjSsetJYA3U3JftH
xivGyzwkSdGaex7RBFnntaMa5wVrsNwURQUZMwZ61weqhjvqggvKU8AV5Du3
DI6Hbrq1ul9qKqejYUExv3Y+wcaafAwSa7F2+VmDQ7RPtKqeTnWejh5LPo2P
Ewi4ADqIuuSCfVSAtDVoQvdfssVDOCmDVkwqgyLkbnHGlDso5UnUPKMIjmKN
8bMVWT+IFM/uWcxtZmkC9U3/g7ogRmBXWSrMDhNcnJ7ItsHFVCWuHpnKjTYQ
J7FaleQtU8IigsTJ2mJw4JpwOAduZqVYFCZ+1U57OVY78rII0bJmItGoFlY4
YmJjjN9tmDYwaiZgwZGIL7ipaze4MHjt0JZLBdD6ygTSdkofyJEkNTCV5o/M
wOAHpNH7+LmNV+XMFSiDpPfH/ZV7mVCc6WcKGauEcH77URwkzCRh1lcc4dQz
c0ZT+7WHP1wGx7nT/V4uvAW/yF+M2nfCFVwbr50owgoTzuRS0s5KiJbto0C0
MRAFz1fYpbWPF1MlGw/G40G7gjkq2rb4Fi2+kIhevO9GtwXEY6OkoLuczHV/
c5zHMfXvRJyeO53xidVGaa/4MnbTzhpgirk+OulNO0REnF5wilUrex6zohZM
8T1rM+os41TspsE0HXyDJsdDBCwzU/MW3wLvuCmo25PndukMx658TEl7W3j5
2k6I65D7hLlFLjfDJSHiTXb3gEXsu3dA0xpHlOzazdmD1Su7PQC/6/la9pvC
jk0NSAR12A8bo0b+u/xphxXNXgtrPN9sLnzo5U8WiYzKYeD/yv2Jxn8mWEam
OiPkK3i6WThGlb/MGeHFWliUWZgYIH9nPRPTC3aLNDnOR4BtJmDQLzNbywMR
DNE/JWnanT7NS7fa0zhOvE2+CzsDXIFkUehKz4jcy+BkjkPX3k+KYoLvQBAH
TnoMJT2DpjhSMXdGxtugB33acPjF3iRju31Y4BnrTMo/z6SXvA8v3S2u50es
U3meDmB0EMybG5iIhDxnL0tttcNQQDrsGp5rdhwDf9Ph9wSZed2pNGoYQPyW
PC95jlDkeiJaeNL7IGLOsjoX/gaoVuTW7iD/AH8yxfgYZ93xXm3ic6Fb9hJ7
gizckELGI/pbTFxzn3KZ3ztjozfenKzuNgXvQsZOHMSKvOg7COku4Hb8nGph
Zxo0Jm/Whjx9eGgBwGCRVHmNOBiONmm/ERQcm6FjCKzt3dU3rlOIol8XGSpb
a0OkYoRnM7QkItMiPwtAmh1JSiSsCCbjpTDItzbrOn9SbhTxk+PdB9+Qj5LT
Mgdjwtug6UiDoLEpECDK/Df+oCZZAIBs6kac7vXbmuGwzLKaH0k7gO+r8Hqn
OnE+3NUbeuPWildCRqhcK4+hOOst+MrRys3ZEnAub2R3Icsh0EQdufTYQQwy
rESJ8S4uJsFLQLAGh0D3rjhgCWpxC0p4NT9XsnllJZzy7zxCl21mgNAS8b0M
QIByZ2N776CNDy/1lrtoHOT1q2kyp7Qbpq67mWpiQRlWs5V6evXBQg1iqTHC
9/Xo77Ku0DFocCdP6KwN9LKxxGvmGj+IcPwHNefQLjqr3OHpcgTjsa1XtbVg
piZR3GtpnoOsSnF7Za8lQXmkWq8mMM4J/+Q7KxxrG/oXd1AT/RR0uVuO3S9W
vyHiRdw0z5aZUvLCsn3iAzTVp56mbJnfErZXJcPP0+0enHjvvuRbfKMpjFBM
k1DDcOXYc0h2sGufeDaCR1EID3PBTLTYvogtRm4Dd+JK+25fg2xfLPyDLHKx
tmoW85o4E7d8SDcDo6sKsGr2ZJuX/mdkKEQM2Vu3EM/AKuN4FO+m9zS69Q7k
2QxsLqWMhMwhAJaSzxC6LeQoYan9t1gZUA4MIYHSduXln733mym5ZkXLrdjz
xb+3EZjqKmUxCAeyqRQh7+wD+Q53KN1EX4lBWbekfd8njYbwGo9lU0wtqvsq
rAZdyz8Zy9UDtVCXHgK2DYrMTnanzb99KW1xywThGvn6mq7/+gvbgk7QPKfT
5hFdzMNRi3cvVYM68T8OadGa9X5/G4//odJmO9FmKe9MdM+I71KPydeA3Kv/
MOSFJag9lctL1hyW0IoLmn4HRt5Joyc2hdLg9lPyzf01RgSxRc824doiKKFV
btv4YaRlbx5gHPAiVMUqpBWoBfEHAamk93/zy65hUFxwdez6C2L+3aQ1eUbu
5n548fuvnZCdvJbTZayE5lsgNHVJM5B9RAZf1rBeb1xhFnFyMDKf1+B6v8cc
3mxdF6bOOj4Q0mRJgV2BqaFdrJhmCElfhiA638KQJvWE9ilYEB9VRTrXAAyf
JF/BIC3ERYfRxHpFWnHBYyNh0TwCau5Hl5clSrH96/9T0gU9aZYr7DwI2Q8X
FnbK+fhRyKb+P3fAPLDpXK0CVXwg2PBBs17IBGUGBtZ5QhPmy8kw0lDtciy3
BL2VD+Hj2riVw/Ilkqz2OsEFbOMq0qea53rIB8jL0xRXR+eK+vYHB1JAdO3H
dFAm3CAPdlDPPscSD5VO0w4tCG8e4ayDBOYTejyq8C/EJgVLQc98QiYMNT3D
iJ0QaXq7s1jXwbTLfRvmOocvy2ovSWyPPwWulHdKGuFJvlkYz9vOMnOzPM8f
HvI+hq1Mhgw4GdM6la9uVblK04RnOTmhT7n+6dCaNUSTes9ow6Xmhurq5icQ
V/smtY/IQ1TaBIjlYSlTxzrzFTS9fefIzIaQ3Wbv3OnB928Vbd/uoVQm0NGj
ler1qqYRp+oGenMIlRGj0iWdDETo6BHcD9JetsFKlbNcXpdlyW7ZyRrvi0tY
3yBSY1URR+VCe7JaCciQQGe2Nm87y/AtTCfRUFQEvyZ2IxAxgnjd0FIKERRF
JUiXGnYyCJ6NIuEI2daxtKhFLNUKryl1+FMRxvKgX3DtSdZPIdmyuDCCNA78
FiAOCtYmrHzb0auas7XZwbwbp0p5WRSIC5rrHE6NnYTTCsF6sj13nEbIyJCN
b/A7KJl/zhgnUHOKRE4FGtl4LQzBRIwCGZsNVGSMOwcJbZolJxuVQofod03H
NGSHv3YHpv7B0b4atEiznlAzKP+XLgIdCLpvYGSgVeHLMh37VqwSDWslWVcF
YkIJrWt9ALzmKVZNyYY2xPggsVeAdiSQ8EksSBZ0R8FknTLaJ+DDfoBX46LZ
1iXj1Gr7Qhc0TtqCv50Ca3tVWwQ/jV7LaJfWEyL57nLVZ4kCl5oD9S0Q2ONI
3btuw8b7qGJNOuqK7aDc6/uYdiW/AitWtWdrdU8OI5iq6Q9kAZVpPAzTpEtz
H2hPx4B8VfVCQmgJat/aw3TzMm9fTVJvgujcyATsNQMBZ8wvdrEgWkvH46ja
noJFqZCAbLP51FrAZItG4b+H996kgsgAGdFX0iKgOlJMBU+6Z5FPBaE3kbuG
ec3xd/UCbHJNqg5KnxeJ8eWCBx8DvWhKMTqpxQcglflrQo3Lfm6EtoCSVuy5
pDqROAKesm4vVV4768BBxrZvPF2eW7caOpygB3Qk8Mnk0SDqvd7QCanPv0bH
5L5GauqYiAPjt3J75Sh9oMj/xDj587zMQNH+NbvCN0Z4+jOFH/P92iEOoETg
b08OpYPCfu+xOXaIltjkNgJS1i0sEoo5tMlUovEUIrZO0JJGcSWRvFPTK4a3
YnJsKrJsk5oCFIMdTtg5bWZFAqV75cYyTxNKopwMGVy85lZHd40kYtvWyLgr
zKTOPTDB7LFyCuMEAgQG1lDW8J3UcAkNgT+QBdzYY9e8d/y/7pSImgcSBfLL
6yYzihPP3zA/BA5COsXC5scpa4mOuxIjYmDdVIfAYsBKPfN/WdWLaBmGlYeY
X6qz+f/s34yWaxS8ZGe5ekp8WCTZwmaRG2lTn1qd/3yV/ksEzmmpA6Qoz7wW
dfDRs8PU87nAGBkJ+YtpSI/in7ESHsXX25aRX+91sAMLFn4ppDKZeUA53nhy
jLXxb3Wyea19EsmbZ9YquThlQZuBJD6Ng7dfa+dJ0fLxpHyHqNYZ/XibI9o7
QABbBcWXrvkqOjjQP82qzJZF20uMi4jioBYiYYF6PnF1n8jX/Se/9jCIThmy
BDsO0PWQ2OxUWhguQfA0yR5Q2w0o0orlA3u8sltGdHy8XTX96QY4U1hoP982
Bpx3zt8zVWRdvTWx3D4vQpT1skMOedC/shkxyf34ql1/T4hICp1hAfqQPBxi
DtyHjHgoX4m5kSgaeyQqhcGmzr6zADp3iCuO4Q38XBfcuLhEteH4oD5cuTsN
WodAxwJjwM6P5nq/IhQQR7wE4wMkPohJ6h6ytoPRfeOIqJuTseVSG8YnFZVY
QjQ12W993HG43hT2hU9gHwV3wgdybCz7Kb98BKsLICYH7G6AOJsGwDO2m1hC
d2F7DkcRMHbnLivTI1C2KAe5U3NmVJlpQ74a5S8sF9Yutu2sm0pbbeSpM6Eu
3Oo3XIxD87TNjEGCNl7JVcdbaA0UlOUh+ymGifkxgwp6BnJw9RiTKfGhPSqF
uZix6UVVXeyjMI9i6PFjKtIPTOybDqzx+ndnb8JjFuyhq9wGuj4wChdjicCQ
bfjFgArF8zYkOxZzLJFyB5ZPCnxhgADmAuxEKUipaQ52fnzhzKBhajgropOm
kgbqgleJaQHWiY5uHakPdsFbnblAWn5uP2H1f4DSTfLX5uwhAc/e4vnAI5qm
vISb7EEZ1Osu8UcCGybTUVeVfe3MAmS3IDxds9za1NDRNjw6Y2qXY/pmtV7X
i0jwtEGEQimr8p0iVCLQHX/GhqDVA0Zwbra02p+95Vr8lI+a3o/ti6wUmfeo
45g9Yt9JzTa0q9vQ1y/JCLFeDjWlZnO7HSZbYmq0+upH0/tC1RtzoRLTAI11
71DRb1fLJ906UsibU5p1+Do6mXipE4NbI2/kEpLNyEM0DT8MhUxz1wnoT1OM
VcWd9AcioTbMyIoE3ySAqTF6APwDCqIiIJdNWGL1ZXycogoZpyCEp3u469E/
JvJVhOpOzyPYMSAAdmFLSG74EbJWHavHoR9lNWo+cElEn3+dtbgv4Nwi6PWE
5yG/fxydERY1dK9gvMhCPCgfghnzF1gBpdGN+Nbx5eQZMQhgT5UtzGLTzAAK
I9rzKusvwxAX8EuxivfpakY89aHmvgL+02lLC/LPOVdy/HCODH+7dmBUE6ij
cqJ9rUwnafazodUzutby86Yj0Bhu5SJ3Ya5QC6ZrJOuYOPGsDsE/uOhvpW0Y
THgulaKFwl1c5w9OtSUpYccayGaY1/Cq6+jeyIkRLJs511QgnaFezOXUY9BR
uC6nEK7ZQFXmNTa8teW7u5yP8dYcZaAgdtQgpDBDSlkbENqzspchhzMuqWpd
wEuJhf0W7dD2+NwtUej2sGp/xOkN5AzeBle36KEjlvgdhPOowPMeLZiKhuC0
K1kLskqco43E535IlomKDkEdv+ixSi91/rFCFA0MC/JthOaNVyUlL+Gy5dks
Rw+b2pvzOx/ekPFw3ovxqqHXqQmt+T6y0jf2ds+YtRJD56NXdBzmLMQUN1qi
6ivTohPZcQTsLcoqwZN/qGvZxbnJwDUbabWlE6H9OyFJJsc9Rz9Adg3OIipE
wugqhzzRAN876ySZo5kqeQnZwuD/c3YQ3ffc6p8hhow1GOuGAyiNmz0V4ecl
8rhusIs32EYIpvdo+gkTj3a7ECdWkYRuqvZQ7xxLGWn0PyxKFFi2rLd40x4C
HmWqp+KitRl1ro+gh2QFFHu+NH9tAK3MlGJdP4X6Zk5nhwbYgNcivxWUV5dQ
ZLs4/6QQ0fTjGF3ZwsDvfItELwmST8aiELk2lLyMyXrK0R3mu9e2MTd0/2+H
yWDuIRs/7uKUg6Ef1rnIo0sb2TUm82YoGcFYro5ogWH3Eu/EDC61s6DukkdU
gMOoCfdk31BQKus92ynbo2WR77+hPyEEQMgxjYatalFVB142fIiXLPQFWIZb
+s7i+EgHdOf+wMt4Xvgdw/P8dq61MK7RHOLilUOcNQExPrpVytBJyeNu2K1p
+aR/BHu2er73GqhFiWYRNdOBcMfqK5AQSl7bgGeg5CvqkfzfHzV84wjztkph
kw9/KfUAD9fflVWHF0or2UuZg7TWRk5kViwmQQ39OogZHY3sYca2kFCHd6k2
a3u2e+UlIiD5SiAtZxfIhSX4nE8ZTALnL3pbCU5tc8V+X5C+vYwOEEFMKMTT
Q/vldB1EhcDOjp62imO7YNWPgAYLUXYI2SaOVh1PkbyVjmtocnlKJ67hwTbr
TDacZj4Ld8A0lTBnzOHaM2R5tkGTKw4qptFdBR9hmGWEIl9cdkyKLO2faSjb
WbkocRgjHPF/PL0wwQ/qZSh9oUGtmqLeykkNd+qavmWT9ltjSI3sFsS63wLx
yA/5NWUahhMExmZtXsFT/Ok6IzPsxfEppSGAoqx6S10PEx3Q4d1P0lij+gdI
RXG6BMJWcKRTgCktAjlbSEqb5FsASOYceEJmEDaOb0CL1tBZlSew8y+SAsrG
aYniiHxom3qiKCZLMM9Kfz5MD6uyUL7MYmveakyhN9+vNjm2kdONp6JmVyx7
uWEXjtsWtBZyXam3Sj5fthL7ifsdpO7SPAGZRum5AGrCqT0cpz6OVbjEUR0i
9pQJ3SEuN6ukIBStNled4hSy3Cw4z7HdR33fInTnNCihrmE2pwSf2rclUEYq
paxykfXVBXwFNJQUMbH80oXa4wK82mSUiuvdsOHRmvC99ncITj+8H38Kle1C
wHcocAOJEGSjiUK/caoij76cdKbLdAdVUy7tMmV6UYCPFsNQdCrCJiZvl8se
Fni6KFgHhQEIm4KZcXpZB+asHC0ANAZSyL00Wvva1egSNU444f/eVuEIlSZ4
vKKVnzLa9HWNfLLRzuVO8yQ7MkhD3j+lDteo25U5/ONGM5QqrKyIkT6PRsC3
h008z5YNwxkt4us/MKYKuS9G5iHjcJgRc2CWmGueB+nMJWBdXzAHmj/846Aw
sRLxtOhTZRogAocMttdrZd1dEgNkkvg/rLWxDIBU5f2rFnpqSRcJemklX2o3
xOt4m4wDuhFzxC0KKktHeuexa4Ey9fWyRm2602ZyKSM65oOyYtY8zy6yDARq
XqMyUywZbSRsh1AcHDN5RIiVmWoCT/ShB9A9xFMJC7sb+DPPWODwoCLQAAAq
aimvn9JAVFYrVLbj1vHOUziJeTrGNoFmLDEH1GenxpZ0uN1zw5Gd5wwckEVP
cDbbkbvYqLXLbg6uW9WPBrmg5T3h67mK704l8WXp5Fna7KvdTilk7Aw+UFzC
BQdFxwid/UC2VL7XH/sqHnevQwbbb5DikzK+3/sCdvJZGq1rwRU9ffrtJlgK
kqhThTTRKgoPiO6RbaxiDaYwQR2YQNXaeSai0BNL3ldaDNs8WOhnUJU2lGlw
LWZDJyMV06wC5DgDkJbPIetxa01CIWsjaYgq1jMGEiJvaEuAlBeecQbyukSa
M+VtbfEi7+yhD1rDy2yx738q6FZ8hLUkaWk8XEnfkEbmFRwaifTpaYDrt0Tl
XhrSyANyTtFAybvYW49Nse5WftGI73P8ebZh/WpefxzUMVQZO4Zp1WwNYaZj
PMclZSvqFkJDkokB8Q5ghupJitHrxCSLafueva3EdKIKs+uKzDyur4IquZOc
TOI7wK/cfLnJzTzHJ2K1rcPURPtJ9stdDtZF2L/t96xfquRpdEHImuyBDKyr
r6ycSJlHbm/O3T24IlPJ/285RE1gHgSy0UIlKr3+LUyfI4hNHh7Y9Bm1wimW
hrLReqVCjOa1kAIYWWEwylSzJROVMuG1hu80xnYEyXgk5M1OntZOmdjd6KRw
+qdGRqC4ZVwn0jFHHYlh/9644m4RnqXfssd+8ECLhAFG/xdeBv/yrrEVFz8V
adntI5jYMNxU3W4nafhTklPjAtwUjc5ysg/RF2uLlkOJhcBJHKpeC3ZPSf0q
N+illWtIWn1B2hGNFQbMUAatjwcV53S3WMRm+bck9ITRVmgO/zGg6m5yf/w3
N4JIHf6VTGB7LMcrZyG+JOZhZ4vdOtslEB+maqO4R3j1lEo7yUeIm1deu2K7
x7Th8iAruW+e9mlSswzFcsfMCwboqj4wWvlXzq563GHf6w5nqoy5oUtCKx+H
Mz1hEHxAQ37kXfTz/1BVpn1a9qwiqPP/47MVS+kGxpSZJeZ93/Wjcq19VYLy
Bon3RqjV58lFWeEiJxqPT0UN4YtNu+3/8OMCZIRk2Al0GUu74sO0wU7QirFJ
mxUfuPWpIa+yULB1BSNCAPPkFw6ALs3S6aZ4YCy+lYCqTNjDtyNqDQzAmEcu
tk+HzutljyJW30RrL+phU1Ijj9R3HropP6IBHbvjgAXHGd0VvWHThKaHWBx3
fuwggfy896G8f/3HQSkUDHXaGQLONGhHS3SuoMF+M9fW9C1gcyOmh3A7Dv7w
fVAErJ37VaIyyrJNMJZx10Uo7cby+GGyS085SN7dCEK0T4Ge6+M9QxX52dg0
VPuJoMwhK8C9oyMRQnJBM5ZbWO5fYwmuBnKXDY0mvCiMsZR8GwlNaTLBxLi9
q2g5EA/dMw1kTQNbLh1VqiQa53KgQT+F2w6zpk7P9K69DcPZaJhnP1/cFiTT
mAREsEWeIkMjwxDdxUv/bGkXiCzgfZZGCETrH2FOa+uNGIS2W2VVEiW0oGB/
TPvQJp0jVR+PATR3Bpp2bSpASQGDhRfUnTLbpAOrnB88jLvKHraXaftrcMRD
XuwHtCE/voQk3tWsWC8qYaiSXaWtlizlZu3asav2Q+ygLl5RWFny13moZjrV
yShOsiB6no1yI/lTHRFUATczANIBQZ8u0xRjkJIjJsje0xjLZ3566f8349nh
GGbx6jVlskBpbdRpsxe6LEsHmMI0rM4Q3XAW4OrOK/PV2cGe3ZidqQPq6+Tt
jG7/bekRwisVoLe0yfFEfiGIBa9oymoLP9DeGg5qcX3aRAspcurO4WPQBluH
t45wS+RHxg1xcdC2aiHBENEUqL9IakiSa651hEh1d+j+UAwawseG9GbSRjXa
VSPQXXB1v3v7wKcmbJIKLMzuKD0z5o3DbfTBRimReJPGOW+jQk6SMOIf6RMK
93SwyuYsblnQGmAdvZdZJZqESgPc4jcdnPyGkbco9DfXa5WHPr9oA5y0Mzhr
k6JCucttZFWS1omXN9+gYDGy/KbkRowVd5sVL9AaVpjGM+zXnUFGkzhkLWpa
ObeYq0hLUPvNMCnLIxLms23IHshT0iPar/YfsTFUxC7foqFJZmCnWZl4cgSm
0S5HeKlnZYz8jaq6d5BgpwooRgojogFGSPYpYAU/pRHH/stlTk0m7iFmAsII
V1QKSERjExPApPccOgbUnWD1FLysXo1gWIvElfZXXB3PktOlPgEyAy+i5yWB
w2ScnVgKSIs/ySvEUb0oDPuqWDYTmpHuMbA5MNp4qCt0cca8zbLfhH3wZQq+
FRTrYjdDk04D6ocQbzQVQYo0im1xpzJYAcF789UGLrJBfqX0IW15jwt2LJob
AuYcU7YX+l0vIG2BcNCnGLiumP83FOVwZhpU9Ymkred8LDDS6jO1pn2XoYij
or5WKY0YaiVRRTbOSGRW+magKD81/soC2CuEIo9MO94kcTs+HMDGqGAYzCmj
30amr8F0T2Wbs6odA3CqZ7Q9IdRyNE5+pFsCCtvkV0FCd/S9QO2keCq8dEZf
sQmFczHCAtfVG1ZEzu4hHWSkUkTAMsAYHQlk2IWvgq8GDdmY2K6MFC7r7nqO
1gl0LKfxEaZX045/QWrfiPGrSGJH7YB2vJoP5285RgtPX2A2oo9s+QakgAQm
Ja1DWAMhtCLyHMf8zYxWCxFPVpJu9QU6AKJ2Dj56AL7IiB8CTqw95Y20hRcK
yL2OBJdpeaC4N1ple9RWgenB4gKfjHfzZTep3OLoOuspMrxXKlMuemb+A4Bi
xVnmN2phMHd7P4Jl3E8PHT5xh3BgUn5vLdrIhwjPxu0S76oiknCMR0Kjb/jF
c5kuv1UDmM7hsQxXEqK2EDvMkIMmD5skvaNTTyfPnVneqgMPS0swpQh6Dmsn
cNI45ZyIJZm2627zD/HIL6qwy2N3uNzA2xKflyEPftBIJlcw7bYjFGK8y1Mh
5LnU7iYamKynmO+ZZjUVTheIYPZRITygdP39PF3/SoY1GMfWd/WdgHRcZ5lz
DL0pX+hNrs/wiZtve2WproJ00PnfbP+8hujDCM1/YWIeLlkyBgZzOCJmoPIc
BIbz1w2iLxH8jTgiX2+wJJ8myykkYXPHdsZoMbLkeRwwBVaDf8zFhAkbGn2Z
cRlJ518OvpmV3Mzi3TMhAzBdJLdPhKtvtAA8KXC8WkBiByOiaNAUmUB9uPvu
Mpdv5YnUfKlRFyVMQ6OAP2M8Ingf7MOFScT0MYmvuCkLrBDQtR76LlUNPWNA
scoNNnx4kfSRAzEk/XHazCHvcNRThRcOnML+nV7/e7yQiLajeVWI3UsYdgyc
J7evkZn3NYJxiRWCympvKx+G7eEcvUDa0X7M69fC4lYEguIFwc/QkNP/VbD4
g5g3XM1ljDXpWXp1/l2ckNO5RdpiCzsp0glM/EMf3lMGiff4RLxngjIrWG1a
ln/t6ifrIJ2scyf5sU6Gc60UfLO2udwYTBY0x20wjig3DTF5cLsROIMq+17A
melFEKrsiks3X1eRaoQ380StuQTF5hiV/nubMb6v1QZBTxe9JglDwx58Q4+y
YOX6pKuEZ+ofMaaLNMMZtcZ5jQYDwnrHOEaMJJneG0XV/zP/mQbKozNHZs/q
qlWafISRB+PrZ6nGU8/z79oF3ZDBq5jXTqMh8Z/SvBbqDIPzP9BCcOKLF7OZ
q7iTQQ0uv4CXmwwTifjoy/oY8r6hnXGsT817/s9nWAOFj7a/rH0Mt2kV5up1
cxqR8+mEuTBcQK1XRTG1qFFVpnvk4jZEIfm7efLTl3WNwkY7UZX52HCJq1WD
j4kWSJrwkR/Dx1V+1DNIqfNwA5tnBy+y4QnxxseAKSIs+oGZ82dzv/87seaA
v5B6/JCNfDyO67kwNt+bFXxgvEXB6NLQ9RhbUTaYDL3o6Hw1CTburvGuYMg3
tfdDfQgJYWOtmkTJpUn/uUdxIDXMhH7OlMQS6e6AaW+zLlYS4Lb9r9p6RFoG
c7QSaRwom5JHZNB2GTk9P4s0DkfEEkvCEVrrn6U/cbS10rPcLSmqXu7ISb+V
6+LyqhZHq7Ggw/mpxuOGYHTHf6eq1q2CVWgnnpI0FQD3zXkMJcrbTvTd0Ks6
RfeNLFX0y9JISY3NSFMiuS20YIrbBkHHc2gVW/isICPyY8uBMucIno59qxbi
NqbDbgZgACtCxiPiHMSiylUxrAwdOehSG2/5W4d6vbUHJ0cWFxcY/5ZWTRMX
rLr+LW+1s/QmUQUGSkkCViTP4Lfa9oEcIQ768MrT9EUyzac5D/QNMD/+xtXY
SkOJB8cwtB+1IyRPVgNM4YaqLuzuGeILHDMaK/0YIYxfVk1i5IN5Oltxdwwt
aWrft7hWz+2Wj+Rq1QJKAnQjYcDfrkyH49z+kYxOJDYiKMnfTpBIaJ2V2k/j
DLb8E/MlDm46PMGuB9xKnPxIkU3cHXLgcED3WzehVlN/qB2c11Oei7XfejN+
RikIF3zUZRkxO+xWPhXqkkJ0FX2DQN5AqsuMTuuRj0Q5LDGtLAwNUVUUhRE2
5/vjXDL3Hcmv4fAEXlBUQXHcV9EnRbQKvgPfvckf4qHVMEERXxDYSa88+5qI
ULIa7/QA0B1vMtYSb2e+edQutec9hmKSQcqcVFMAaphBE4QWMAKpB5W/9Vws
5SFafC4PwXiiKtSl7sRFybsbK8o5dXclBSqmUyL+otvXgCmXh10VqqZkR8Ry
37tj0/AMBJDDXo6AmGj7LhsdWB7qCrJfQ05BMy/IFT4Fd5zUj/85k5KhQHSc
tlpb6K7x+S75tBwVqSVEtidPETpBNpOJ0Z4uLlyBXn6kc4UCAEQlz/95aqpl
2GpwDcu0jVoCN0n7BdPItr1yMA2hzPV98oVYDW9P83BCRsPQA/tz52VsII6r
LPgC4jrMXxXity49vv5e4U05oGe/P5lmZu7HG23InZUR1sBvWuE/o/LRuXOU
0bpeo21Sttf1Wzt8uru3gxQnVwtdZbOjAj6OtwPYAniqbIZvntCVhLeEFzpo
DR2OM9WRdYmtMy8q6lnXTDWo8d0G7Yv7QTCMX4NVYxi9U0O+kl10gKazg96J
UQYrhLmIEaNekpJS7qZbL7juIVXWuTqSkcQDb+BEvh+TKpqCk+Ay1qZsnilS
UjhIX/i4u4Rss+29mWBzXG5wnOv+vgRHXc5FbP1z9baB55UK+2RTA0CZ6Sjz
+8dsS+ZHxB7K7quF+c5u8SVZ+4aCnqA8OAHCc2ih8Sj/cCbkg2M/Ls2hf4be
mu639ccUHlxdrbjmODdJhPR5z9Cv9WbAh+6XXP4YAggS08qUr7g26rs+nl8z
KM9du98AIIyE8huy34xFpilyXwq7oSvWVC/sD1hw/iFe6Q+O2foiDyU3PcLV
GiCodg3Yko16QbeMb0GbUEKeSikNRuDNkGZjoLKp27/34IXJhOocv7tdBxyv
E67z9zkseLH8UOnO/oPHtA4Dyb6NFbignQAgjcD1fFL0Tkz6drOwTZDxg8Dz
Iz/zKYkOjM4cxXKy+XY+DVpYJyL0iw/ePC28m6VwHCh1AUvkS3aWOPqOsDIy
z1h5HHbv/+2W/Kkw5btx6wNOZgjlo8nW7jjqxxUqCYTq0ixgHJrLZppsOgib
RYvXjKAD/hucRA2/HlxWxBriD/zJdFT5SI3GtbQadXw32ARi+hAAw0ainmPx
XwiOJV4d6pV/MTpds8TEPriTMySyHkxy0kIm3YmGaoJvnNwnX6HAeWnqcR+R
dqO22LUdDk0u4mnzFiUJUKPXjCY7uZTWQasGKC0xXlZaEiSObqQHhsB/4jlR
fohMOxorPpi3DgdHIYKqSSGJrnO6Tg5B6M5uQJfp2IGMpHh6b7TXQDambvwO
LjWc3nEfrMzHFiE+OEhHU/Fgn/jZirams2PwFlb9WaoRnJqwS/121byD2FbF
tDe0y5CvzFOT8ctMRY+4zXjCmEETo+UVj057ItEAwKgFT6cdBu1WR+zIQLL2
x0Q/bKIC4T1iIukThGNlZk8cgpErmByuOaWYXQ6RsXcdLOB5Uil8qs/fTuSm
Pt0bSnzrJrKBQVLMekQCyjM0hJ+/DJR5VnsDdVyzzNbLcLXbiJCZIO1M/qu/
54O6ILkKN6qhQvHnGfinI+qMsWVP9l4BXE+FWEsFn7PY/HGc1dwJbyxUzC8O
tjoF4a6FslA54CDal9tWzi2LXQpmdf6aRK82M2WzVyBGY7JdWDCg2h3otC3i
2QCC0JoIHECXrCLmVGtTyhnvsEuteoAl90bFAUYg8MgwXE7tkdi0MfY8DJg2
OzdcpK73N3o7JpYR+Hl5N9uspxvSB1vhG8MYw3Ha1dwSW5V7h4WDzV1J6CTV
h6MIrW0PprCDYJn7INu1pdXZmRRrHDjzanrL7EKqv3zAoYJTp00NeJUHxv1N
tlA1eCPn/n5nYM9Rr9OrvhIdfUbZM6ricelsSDmC2BDXnPYpy4Xoo1WloiWX
Zl8EAxP3lH2ezYU4GVG+NIIVA6EpAp2XiwIAjfzmMMEMlmyC41BUU7IGLrRy
TsYylyMa6fovaLrjUYis/BICRykiio/LDkBncBDcZ7+k2u2GioCYvJWmqwEV
5C6LLQYTMjs5jugZ7xCgVOI9I83wWuiF+/+LoOFba15jtiP63flJlDCHBJVE
m6gvKZx5/u0w8wXBfg9ufCYS4K3ZQwv/3hmwBle9YEL25QiK78XZoOQyMfsl
gCenpfcYcMI+psyFC2yXhcuMzqwsfjMqF4dFd1rSABQC9vSyAFQHcN3LFB95
dj3VsoJvbt6wfDCswcKwpWMYCxuhydHUhi81rUEQcUpBHekZIQSsVrRxyRJR
LB9D/eAxnWJJhGe1woB8mK3YC9yA4f4k9jzbnArvxw1DZ0ZEOJcJz+WcmDRW
HBzbTPsKvp9CBsWEODuA1YdqdN3PC6wDJCTW8b4XqxJ+XxtS9CSw/2N4do6q
cAIl/06wRtnAip+4JyYbo+/rH6WHpbJcFIhmX7Wm9r/4Es3dl8iNc+prtXNj
rbycf6gpdD6/qE9dn1qPHVcP+kR3sC9xkU79p+0c6RAFVQEQ1zCP20WdZT80
BRfpf+gUT8kf4GAGu0z+H6yeTMmWg4SsUecSAnxNGIwRBw+JoFgzcE83PIEg
ihe6VZ8iQqrE39SDa7Xp0AZhSOkAb5Ckc/UsP+BKwVkbpx/NQT9KCKm9ZUpF
mli0t5gM3uFBUWWjTosrIidASk2O8cUVY3Y2NPZIzoWX/FQEC+yb/2KZ8RJl
hvAf21WUNl3ChZjuMDDCZMJyBvNfW9SCEys1PkGawdJw1gyolceJynp6suID
JKc6d+tFLeobKMno914g9u8rjrbnE7AfSi77weQVphMszsHFgU7SbfWHZy3l
Q1MHUPn3W+651km0ZJ7R4hsbAZi/n1ohpQcHzLMNGl7GAxBntyStt4saKfkR
wozVtmaY98DI4gx3rhvxHPw4RZdw5rm6I3Wvvq1ovOduHk/u9m57BmMxlZQW
cMWBoQD4AnFdwpaNSjxcfA6vXYEc45t6vgn/HEvqkfe3HkxnnDxh05Vlo8vd
ZgZfVzgPwMYBuoGgjkYUl+YJGSaxuMwI/yEbHj8fFXifqR68s/5etdY4F00V
KXGgj9Y8tP+cKHSbmBKlzZaTSbCsqJlCzj6BAAWyV1O/YFcED1VnVp5A6F4K
GeCHSsbSBQ3cxE3FrGgkKBcmE411QvK56FiiaeFNO/7dD1WVQfVI4PSUzGNT
xGK4ubmY1VILhiRXveTNUmvmlZeWKXY23slAB0aYEIlzSTVqCS36atZ3yscS
PQ+sAQh+U6EXEsF2LFTzEp2UBCCOw964eQdl+rQBth17esW6GiNso/ZalLBl
3EyoTT4GaxEsvr5b8SHP5N4jA8FDezkg0gcgjD5hfYCFBBigRxjTepN2LGkq
UAIDNL4YTSwiIhD7vDEZDf0ACgyuZcQFE8ktiYyCgMLsDnQ1SlId7UeqVNJ3
ittDUBEK+W9wJlcItwYHRQyjrgKrdt9/1EGB9qbnqIfdwjzTj1pwLeOJZ9KO
M1yMFiYvwsnf2VRTWk2hk3mi+tPNOG/IgLVYy13fyW3KmBbnMaNAYsX6eAOH
wUunZ27LgXBoirHOGGX9Io85ACNM6Xt82Dmr8Hyl+mczzSb5TAt8K3g3Z9Jg
cdyWI+0IfVWYHeGjpt8a7j5YtQAj8Ped1GFHFxwskyvGS4i0/IF85DfkqHpZ
alAR3emh4PuwRYMgRqFkrtArJp8+gGrxzsn58QW3IfTI6m7uKnNarj2tVxBw
w2m5VT7wGxruu987ApnMVtCUJtlsO/U1WRk0uT9SioRP+hnFeHo3e6l28cqr
YH3Lv1BwqSnxfamOVjbb/M0CQgCpTWQR0F7RW/LGEiZ0SW88NfNmbgXsLQEp
bAPKWIodeeR3Kg4eBfLbDFciE8w1OG39iJLKgevv4gB4W6ugNu9VMvxdbZL5
oQ1ni1c+PelRh8ZABde1H1sWGg7VJULNUMBSGeeKPoljGyugxUOiy6IhT9Oc
eQJJJ2TSjgSJzQEZl1DC7Q5DmNTutry57OMitT0cVFfDGlvPzJfv+t3zxM6f
kefsO7Fo+PCMuMBSYi1G0KV6U6GGCJdqt3V5GcT60C41pD535+HXqhM5M/1J
8zEmhFTNe4wsp3vYhuSfc1Wg6y0ocZtJvha/J3J9irRTgWnNfHVcVL9DZp4u
UjA7RQ2BFGnFW8XqkXFOlarTMVNe2IGcmcByCYWN/5NFNvqIGT4YJ+A3Hmdt
oMtIIei15fDT/18XBtEY3Rw6eZnGVZpfV2GLJ6oomV2ENqchraYHLv231bu/
vjntNM2iSnjOFpt7lqwKVP7Js5Wb/sSeAjoUTS2aGLDvzyoPHMDjV/FRdo8p
LETjw3UwHaQYopvmG4qwf/UTOsmEOBBzjLm0kwFHXmHZ7Z/1T5LqUWJ5L0of
fYbB3nz/c99vqiYZhoQVrKpxVkGp7h14fB4af/DpWYalK4op/iYrQs4IriUi
+Xq09Q0HFsx6q+ZW7fqA/OWGt0N3ZYNsNhVcmCDtOBWAsEv3nw28XrbBigE/
2Lc9P4d2TbAyXJn5Y6jVoKALbJCKXwPw7kjRFIw8L1TL+BP20nPYXj01NwYF
nFXRpOTxVQruiPqbyNjn1kVMwGfRkX3RhqwVIACjiAkIGZ3uUfTc1Muyk/0T
KEwX0GPOUYsjVukKBoI1+y1RCsK9/OlWYLtm3ZoxhSSeDIi9ECkZ7eEv4mng
r5ugb82+BtnFqCvx162eDN7LIskJnZ0SCPlPC9ZLNUjOtPnRiUTzxr28OFro
mJD+HuKYPziX2gWkqhQ2jbEcc5ZBEavoYGO2v51ReU6W4AjbBb1BN3hdvlfX
2KiV74FoUT5Rk/M7z2cVrv0NHkKVRt9VUMHkgFb+0OofjBB3f9eieeHiXDU7
GWtki8FQ0iW9LG+YY6roBAu/yR9zYg/+0PqEmWS9U1o6oEV5M+Po9AkHQ5eF
FjfwdUPssBJR9BXAVu7rG2fpSnsGepD6WmoMe3XCu5JMuUwMKqbRsShWsCFY
Vt3KiaNJqKDGyNivjpuDmjCk5OqZ0AEj4YgbIa+RFNf4/4KcoWuoUkRAIj5O
r8AGLedKaYCOd0NFfBJrEphLL4hOOt/TWnZaAfTxn2Y2OdsTiEdrKfPsb/vs
1y1xgGLnLcvov80CLQl3bfSvYtlNBiY0FAAStO++mwahDn8GCsLnzMGOX1uQ
NHZinTYTVKZ/eipNmFOjxxqQG8BPZsl8BNmyuh9o/ovfG06B2i4bSPHxFqAM
7OTsUjkZN/Npf+jhyGLrqD2EeUFevkCqOuobFySj7i7Lvf7bwlnGwg+3Couy
gqnXIHbaPKngG7MzlOEnoH32wzEP0O8qnA8lWlXymVn5HEcjw28AKtzjljNM
U1s/QdgCo7I1fHy58pmrKFfHawGiiwBJINCcAQGEpHxKxsM8nwwgD9aG0LdK
+MVKqIw95x9LJzFDOW7tcQN6TkRRisDH8iOCMKdJsScnDrQsN2Au5ubb3zp1
R8ng9BmwGJeDd00IENa42+IQ1QZQTDVDRgjPYJgMRWEHzCe0jNE6JziLWx+I
pjty4XQ7Z9lNYQV+vcvM0luIR8KFvkFg7j/eD64Lng2YymGEg5m49Ds0GCMV
Vcy7H7YFNHwIrta3bXMmtJMddJt9/6v7PgIbeFh3UyAcGATzGN1fr1utKsTc
69tB6cU/it6QuyZ+ZNJvucw3HjC0YUHt6zwW0kM7pVRla5iBgZKnMBBvCxia
5gnMWwbdWLd+uyCtQelPNwNpDl57cv7l9BYAo8fu0lnBZCjr66d4Uo8RBAjT
IE4DLTQXCi3onymuPMddtOaiaXXbUnSdlbKjjIFVFuzYvr4v34kXJkqrUhxf
5vQDMjBJbx1eFcXke8/hm0IKMbPeK+TMh53huwSbGqL+C4wePc5htLnS0orD
VBNJuWxG/SuEm5RV1RPq6CcfTrTFmEgrtf5hEI1zhSI9hSWtwjbFMWTbSt/N
7TXZkVufkUrzeQ35x6GjxiKkrlX/zlrA0P5jIFzgsYZhUU3w0Shr6ik2Tmqr
5rpti2lNTsqe2KnSpPi5SSVy5O/txUPEzsw75wekK28S4/5dzVHzuOA+t/RE
hPo29vYOCiqso4R5j18DH7p3lAbOT93MjidzpDr/Pzu08qwJvzRRFdAqDrMD
fmz/ePNmC5npowjlNFb4m8hJQkAvmL6i9mUonrxiMk073hE7ZmuBGzrSGaS3
UWxzXRzHWKL09GPnn4CpEBP8mdDrmoWG0Jx7uSpVo88CWEJRCRI4S9n01AHm
V4zUfzbW599FtEgZcEieE4P988WjZ/bYZ8a5EaZO9byBqkKr4mFz0xsiHmgc
kP0pbgSGVCW7FumHdk9x/LCoaEwp3HjGvysD+WLOnMvpz0M8NygBEXuGCO1g
pRc8Y8rff7EkfGbwyzLREHK9+pZNJmPDzxG1Tn2ZFOoDnG72ZD02SU+FcBix
byjAbs2pVeSElxrWNAMjUboRkXB8IN0i+1WFsS1GPPsVRt/8ldZgeMolYghR
/QKATpoO2tSmsEzGWKOqBwelPiipb2qDCvOFcPfXCEKW8fOfqfyRsJ5zfuc0
b3KZwHZflXElj+1PDgyYsepF7TL1z4u5o2TMVf9VQEDNWQ1mzfuHrHLAcR/U
CcaPIoUCfDdY7W02Hwk+hHq6GKQnNcP5UFxsIakM/Cnvyb6cTiKo9/eo5MGW
nJW3as33SPbo+77Y5tooxQ2Seo/vgdi9ajlpDg4rLN/j7p72uYBXBaKYsSh0
QwQ4idnt10/fI+XYj+oJPFMJ8OLi7rRniO3z4k7+4sD42uoAKA4iAqgIDgFx
aBale2gwXwAtCBkF+eZepIo9EYXrmPHw7wF0nDgg8PHZO11kzG6Ib+V5DmTV
SutDqZSS2t42hCfUkwNsVJvM7wzGfyyEeR5CfcooENF2Zf2gaYDBYYPF3jKC
1wAwerjWF8A8JzJAKx22xQNmXz/2jXy02Zn5H87XbYrr5P7d66q1608AzFLh
S9D/PLwj0mJLAjQoLkClK829lEo3Dn9xEv/3yrW4tdOn1Cxx0DEyDb5m/Gyd
5ZcqWH+9l/p7OSbn7oug+VsvH4mV9yc3T03L4mbBkIEmUBn3gfLLJf6+XuzJ
XuqLHR+x1KvJnuCM1pWWOOszCtPVq1cje9bT0C3a8+CPokQcpxF2lzRrL/r2
2PgtN0xzH6i184Dv/R0PE38hmLl3LzSVpa/1ry9ej+UB+clV1jxvQ9dhtOaT
I1e/TxIs08L1i7j9dY/8juz/qze8PJc+sop3ONnBmfTU1nttOyCeo59lv91h
qbHiLAxzgdO6dI2f8nl5012jkgGZcDAjd7AM/DM156sP8bFqYsMXuzWNgyok
F43M+OPzostunDOh886zjiEz7J6xVYfuGMcM3r17dm2H6RhGJZW8eURKelkd
xQVjboRg+ApkrSgxdOhfDCC8TqEjQEJp0Seqzq03OaJIBfgFjbpJCuUELLtX
K5ttGTKj0Dg+kZc2gW3ei2tImVUhoxc1h9lpadSRubk/QnF8fv6HnOQUGVnR
iJiFzsusvFX7FrpTN6eWucqU2XzHRFcXRwtxNYm02UG8OSu1HhtxFglVHMUu
u+PuzB5sVk4yBTrHdVBtvLSilwJwkE20NbU0RZg+XzVN8YEJGDZuGsQ/7NKA
qpJjged1jWyGy99tBiNZbSdeKfJuqHMtAYiCgKRWaZOlCHQsHRpRdHFFipSV
imGVJ3f7ID0WZHdiP/9Tyv7BWkcSFTWc4IVT6ilncIN1i0+3INaf+fK51N8S
YX3br8p5dQ64nnjpPUM3buoYSm7d/i/PZ3IViXEWsZVBfNE3uwmkyd1svPNM
xKtw+dfZvUmkwLIjvMFBf/99LGz2ogK/U+AEeiAu1h7x8QGLmkqA+DBqO7EO
51iuXYlf0ugeph/p3PLsGnVh1VIwQfRG564MKgk6HznVRg87ShTzEwGqirKk
vQ3KQCMRgzo8tKuz5E3orhFGQRaWxHQ9oHe341FFcmqzzt/mo9j4D1YfIp9R
ghKlu0wliR12HVaWI43Ubh4EYcuyUN/nr67Jw784TqmxbJBoS03Op7CO3teq
UD0AuWo/BrmUK6lnhNu89P7955ggRy4Qz8YKSdFNGwgF03Hg9ig8wb3DU2HL
pYZGkwXULY3Q3cSOFNS1D7hKApMJCHamFMpMQjgtggXCkZ/7tBYtvN3wncus
/WnJVhBdt+o7eSoXlwdT+yImThJTp8T4CSPUckqIQovVsYGsyKSULiiMVmAF
vto88dheTWSiMTTSac3sMz4kyI9MX669BhP/gaN5qxqWpcFxGsP+gq4WoBcn
f7k/HmjzK/bKgHxAPcoNZrhaUDl6qZbxpomvrsnaHbnF8pHA1BIWmjYB02Ny
JksB7XRVb3dvtW4sjgOsAhV552BaLwfMoiV3j2/lh4nnwldCCJUfrLwl2Co6
IhrDUxDgbNg3upODhwNQfaR4b0WGQiuDpHGsbc8/GHAr3P1zxpAnVGvflNKO
odAB8UCpp/mOhspS6kNAdL10zR7j5z4txrEDhogQmKAF//I6Uvf+YbVkZnDl
wLTc0487TB32WPhlTYGpu1HoQoD0Es4W2pWmD+7m4LSReH/8RCAWJHeXP9qS
9eUtibe2ZXH4v2To7KbMuk4wmN/YWiEpXOIk1PY2SNnYsGtoOQ372doxu+x4
3sGX0r/mgDISD2iZYTD0gQ6OvWZQAnQ2Wtxv8+GDTm577639pjJ7mIPCvnoC
DAl5fwCeRHbwNtBOxQQ6WmX7ya7Vq+tiscAL+sAxznGCO0D3WrMmyGBQ4d7g
UfldsJaMmx/YqYPsIxMrjDsrsLv0gc6S/k6DCWDve21SsBYvpKFGfemvDj9B
NoMI0WY7bRuqeoGL8P4oLXwncMJ/3S9YPnL5g9CIC6HgeTWpr5PmqNqkVXCs
sVmMoQZTsORuEQCXKexKVYDCD6sB4QO42ccXdSJx4nBninjaDI+cgBNcyckJ
jIpFxrNo7sCIvFolvteC8D9fUOFI3fa0dUJrLpePHPMvrYWMmCI6CQXfo3gp
3L2rueY13uA//PkZr9SZbMqoS2ZLJ7sVfq7csKox/Wo6Lp5LIK4fCpBPSPOs
zrzv8ffhLvKWEUzsv7CAQ6ZOhwJBRKgmDR2hxFyy/RdzZbIXNPi109CgofSR
xUJn8EMc4o+vS1QMjY6wQqLkk7allr61uJh0cHBIhJ7FPSi/VROfFhlJ/xV+
/Lv3dVaP4m18qgM2wc91z2FXYDEywpAZdn6ppFSLOamsX1VR+CCTaZ8bIUbQ
DwKFVWHqvFeb395udm9HdG1EP9P/IaPs1KJ/dbOgJwuCMUyvdGNUfcM3vk2+
KUZOS25j9YVcCeCVjycXN4GUHYYHo7jMajAw4qM0AREU9zYIjxbd8nY2p3X/
cMct5nTk9EOp84fgr45vAV/G/JEgQAtstiHNooim/vLZm1YXOzMECXCiiN1M
sRDYMvKnmiXBgLx+N9c/NDTdFxbZuKaX8pFzy2voG8/k8jEB4MwFzbRVpyWg
ajx2gJv4nQBr717lrn9ho+X4PKpurqgiz/X4wf09zzGU2gJastfc+EFSK209
ovNBnXaBsLLZL2wusRpM6QOyyOHOtd3MQwe5lmQ86tWLDX9WihoT+qBA3buL
/tvOKRB5a5TNhB01pE6yvKZ0Ib9vbOnTqniWRhe5AJdmMuiR0GmkE1as/4W0
HnoD0gnzvPI7RfQEN4UFpjV5gnVpiPoDGOWRCamz7/62kwfkwaTfmFfvFSGd
HgoxyYnBbIpOfdYvGy3XGL+4ASwyJm8Kj267X7sK+By31Lj6vASPt4IpEFtr
n87hNglwTO+wGAMWwJLsUm+pjnkQZkPHSS8mSjVMMcG5Emd4HUgDO3oDhALG
rN6PP6Au7C58ygvXQ1OiasZfI3px1ds5Dv7/Lt03OUhWoPffTob/vK8vdfVl
pLDLp4hnGZ5DYxYpDOcwkEweHH5Ya+x4aWolk2oDsvRayyBbm0TtHQ2vW0sj
ikfLLveD2X5NmDJ5r13dMnEw5WXSXj5/SDYmsQGFrOxrptGbykov/HA0lnR4
Vc5LPpkF3zAIQQUhkULynK61fLONZGUlnqdF7plx40hK8/3etpfuP5q3eHDm
L/WVlCxOqaIUJTBykofW0jSVq82ysSqdJjcKL9lth8xnHZCIXQHngMLZNr9c
3XmIshl2DkYsbJt+yydklyz2gvt+n0VvIjULRM7dSjz/vHuAHkGYIfGczhk6
3v/4/Q3YTYdqUJEeIs9pVJCHgsAU1YGnQTFjgg5tZRi7Hk8zzApksL7NBwq7
yvvPnVaJNCPqsoyO2rhx5yFPdgiovm206MNE9EwHkUkWJ4rwbg1iZw2azmCw
pxNzFemf6bR2Lrr0dqqgkg6+X9lTv+3zgUW3BudpuVKs5r0ByIrVLPAQ5dfS
vFzRWvB9eLlbUhXn8vUBSCKJN7G+jGf8FURd8/YtumfzBf74EI9XwHgQ+Tzb
nOk7keR9wvT8CdYtN2hjqze5ZoMm3fzC/xOqb+FmDqgcoWkhGpkYDGfVuOYA
TfkAc0BtK77jkhovKOQlRzH3oDaamcIY+mX2AsRKKWeViNgeA5MJVQf8OHQJ
DsjpDSGFC2G6Wra7Dloo1NQZSrU/nsebk0DWbOEo5C/LpMAXv9vcl3CwQF50
fyhqeNIFDOChKmkok65ED7dI8441lFcsdZV0rh1MSNdz+MaEok48EtAZtpnH
gGEIC+B3VtoACFjF9UIjdMPFpZX1v1nErqgwhEmoF4ZPB+ET8eeeaq9hs5FR
SSuNsqXX78jPvYA0cs/5WQg0iQYXjuxkA68afpHvVT+fe25ATkSt1XgrY/2J
3DAaI2t7dCezG/TngVctJWim0D8IXWRTwxpjwTIJMdmihigY6N0hGpw0einJ
38wY80WRoC5kJkvZkWzQL4iUvicqLxSElIj58Vbf+hYxWl2gY68pwj1tRh5T
NA21em24WTMJze4Qv8qUa8OYgTRLtwnz39y1GC0FRKZ544igWyos9G9/9WqL
yPLUiMlz9vIj5ZJWs+j7tqs/v6eekTsoJQaRpYwMNJeJJpen7PnnN6G9D0rR
DImsZG92LdDQ94VejB4vOw18N0AWshgV/A3Sybr7IAapw/l4kcHv0BtK3WKe
daBZZCz+mXZ+hZuH4BNOuqWwKgg+g3YA1MiXmErNU1iff3fxLIYMaybBSHF2
laH+Pyl6KsroCDgjlm5LQLCWJP8OJN4Uq6znDDDcmT5DxLC6umeDA6GDDoti
tT5hkq5vmdoknrOwd8tsjLD0f42Z5lPXe+JTJZ9PkRv4GeZSr853iLAAXMO8
A1xFncGPzN6/owOAgQuLJCc9UviA8HQ/S+edWnZVAaofBf0XzHaU7DtHzGQa
vEqlYtIC7lK0acnTjEMEXVn+OuD+wJmcflgjUHjfoZdZ5oqqfAxjfHuWw7hy
FdUA+iWS0Tos2J9dbuf9qJKlu3PJs9PYGJrKWz0Y61p+IJPy+L7pCo1M8gcI
bPoMEN/wyh2P6q5EltREgB/uc1FNBMcXxw7tUe0NOrFKZDvs3/bfTqw4MBQR
NWh2VW4dJCr/kVg1s1wDUm6uOqH7wPGEiPHKJQQ/XHhcL6GtW1R2CDraXNi8
4ewxkFJBFBQbCv1nHjF6E2D2XE3bBnCukpjgPCqzkp1bvXQ0UbwJ2ACvjsdF
pV9JpOiwVbD932D5f2Zsf82pda2r7swkRgKh9eXSAY7VWcKJ64gNWk/mD3/A
/eeWa37PWpxmMJXhOXv833FsN4SmTNQrSCrnl+zOzrp03OLNtsq1Nw7+8DHH
+TGYOuB8zEs2OjMHIhXAaK9ZnLgAEnzLsxvn9dzBk+2jPRrs8q+ZAX5r2vPM
C0nVp3it0MdVr+y8aVJYu4dn/jeLOrElB67M5yEpAH3/WX/MWvHyS9oOoo/g
uAMZbblbNpKPUIDbESlRLEW3hZAsNKq0no9MGA56Lpdy0RGWz2bJxHaMBuN6
zm2oSMR41msrfIUPmtss+fRDyR84Oxv9oF8kGue1kZWPgwX6oqswcT9drdp6
Is6wp8fGjbbf74qHZRP1eQQlOnZpxvsQ5HxL9j4TUWZAlU7w1xOjBCmTqTXw
R1V8vML+4jAC6WFI4lYexAXRlHFI1VOXLG9j/vKsIH9y9WeTZRyY841jCFcG
TGBkgz4mUNMOIewIf9AB1Hy9jdiND7TLubnyJPpMpH7tvFpE4A2807b30POH
6smn49qcnXOQ5bdX8HYouvL+vclxi5ycgvKNbmtJX3RWrZp8tMb/Lm7I/4Fz
CDommlXMpxXX3csjVGZ1JxRPYj8I+cgNWNib4B1Sj0Uuhuv21r6NbQxC72CE
ScnnO4zsjZSbAjl7Ob39bvCuglAEhJ9QsMY530URVy8Xt3otXbdiVomTCM4h
cRG4AB/zdcdw68LGOZcuoMG0nlc8IpZ5ohfeG4XxrH8CzQx1nwJRfneZ+hjE
wt88ia6fNU/egVNhRqLOOA+RYsG+TEf1w20nFShJDlZkTR555GcAWLA83ISk
lo4TqixFjkIm3/q1avqxwbLX7vWFSoVnIZxZAiioALVutuoelG6jNKKsBZ8D
dymn8537IvrS7Yi3APKQeM9/uSlsN74aoViiCnywie6ytr7keATHtwaKcVK9
LEhy8ji/y8Rmpl+DMh0oDq1A0kN1g0Qf5o6TGDywYRo9teTdjfqeQBA3sndi
NoF+JLgl5zWZYOmv2fbUXIf/nbCJwLWBe1YKi5xGgzruVrq4JuKBlmYLBESq
FWDvbUj0RgKhr7grOE1t/487zu3VD6WP3lzb8JdiCdkKKolMZYax/ULVQF3O
hcpra7dxlgTUCEBBs2aLa/LnUYwswf1IKjLrzLujsge/kRtcZA2LwdO1dPuP
yNgpI/eo3Ri+4IOUnsj+lUobbEjM+t4eEPYZrE1hubr6WTQCDR8BPLYYk/hA
3Fh5ZYG4pgjM7katgnXfV7cRHmg3SpvVDsQ3dGrS8BVaxoMa2HQ8xbrqttMY
d3moS6QqlW6ctNolxtYMCCj7ar+qDoz5l3zeIQ8YpqNqzphfajARkHS3ujo7
+2Cq0edSBkHqZgp+//AS4PkZVloCPjKm/4T1oLlrv0l5vY67BkSrHOSdpWti
s/3FsEbRBpbbJ7P+EqiSiI+NNakWkhvAeOvBOCyQki/L6mEH0QsTK9Nacl9K
dvqhj7vR/wJ6zaP+O2zhV6PTXiGwdAIYsx2Z1mk6472LYkl+Bx+GNldgBF2L
ajgu596IE6fLJHrW6gE2fRvrOebxhPZUUmT4kdF3dfuag9Vni6FHLAiuCIp7
HTki8MkzZv0va/Uv3rJEt6dL0Gdm0W+UHd8r1fgTItZubfOAZ6kg6kA9TgJ4
uFe2YRkPENOP4pT6IWNgaQJm3Xrhb7JtQv7ui7XKljqsj1Yx7dTTCw/YEl91
mvZZkZoZAUeOelMYg9P0kMb5eSa9yroBGYgaAvT1YebnZ672EsvCiZ7tY3PT
w2xj3Q7icS2eTgeI9nwB88paTQ4ImZr5vxUVG864/YGpfYYxDIHuVWVyYw1X
ssxzewUek1H1cAaI6g3pMdiR4iRA7zADZ2Zgwc/E7+xiZWzunZzYpdzB74kg
J3OhQrDChxFzou2ScFvEVlxPV/XtaUy52Koe0FHtW6jZlttqADgzIkMiqkas
wLlyVwjFKHcI0pvJVVq/TEnphYPUXiwDAS34FkHB3FP7OikALU04S3iIf0xv
hCBKDaEPBMkfC7b3oIr0pkLX0tgtftLnmUNxKdII6a8XXbRkJfEmHVsY4jOi
mXXJb/PjRQONFn5l3jrjnFhhsqB6wvj7ucWydC9ufSUs5b+ozE4eDRi/2MLx
MMYm/TCnpYzmv54Q1brtirSK+3Hny7HFjzTx57Mg2HfeoBMfdaAferSu4EPL
ULvhFG+b3qaBoNUgw5DTPXACf3yApfcr36DMLof6mqKdjdw8e4s9vMf/qOyF
koogq0VtM9YIQQgrHBjpVCadOkRLNAjvxCG976G/aA+fhCpjBkv9sn3pkJ+a
Wz/oSuq5nAZ8ucZstmOxxHsTyegC/fa8Ter4iavBUsb0NszieUbd28Ti/ty4
xh95jmbgVLDjHvyHB8U3ZgOBcD7YPsd70LKS3sahFBB9QjHW3445nIXmi9MH
qBuOpYVL7Il1OIibfiw7nTNjcVa/Q98DEYAPCFdmUQQx/SLBTcxM2jN4X0J7
5aq3nBcIyIUByjD8R7+mM9V2xOU4XzSow2kF7mDAKlLIJ0WrDpriAhAji3RG
qoEVFNVqTwDMZ2+iHU6Vly3csH3CxQWDuHBm83p5cpqySpD83KIuxp372PXz
QgDUT1B70edDlY2yCvPFCJsIbDTGha2hzrTq3S5rNQoq7O4UXNu9W201YPqy
yic94jjmlZbY+G5fGrHAI5iMQzhe4LPxpVo4eld8+b6HF0lEm5UBwN9PA8Kr
1gIVw1e4VBPSCIYFDDLopr0zGCdNVSHpEPar7qWiQO4ocGYRWdzFAPoDkXMx
Jn+lDsCZ61w9bj9Pw8TkooeiPJ8Sq9ISdTbmmY78LyYiLczlEI5OI16rJpKj
5deKud7UN+BLSLF9820vt2AZdoe20DvF6Cuhgf4Gx3E+qmcVg9pvMhNfJn2h
5TFE/hMjLswwfPAtLH57pggtIEvLlyrLl4aBAeXug2E1w/o2mtS9PP+leZsr
lRHKmlKpk9kU8W1lXlfx5i/Q36WX2JyXjRczgO/fRqb9qkioNTEedVq3KHbY
Hwy5d6nbhQXDpV7cpRiAx3Y4rcnhES/GTEuTkt4BjXCVy4fnbd/sCVVCa0oC
0kKPXFMIMjEI3RtJ7NbYuzIgNwhP0sm4U7rHiDTPnQtftu5wLK+6RXa58sYH
DckeRgYMjtQTNeHy9cm744ynBDBrXyAadUKbjV8IuqGF0QRhGXTq+0c7khMv
aAcs95omI+VP/msfViQkY+0lLQW7AWCfYWsuotdtig8H9blWcUXKm9KIRDZV
Q3FJJkvwxjCF6zvwFL8M7Xr0FVNzXQg77KtA8MS+KFO1V925mC0Jdysf60jU
H800Hm1uMevM4VwIuGGyNHLVfA1YeNmSyBUz97mc7mII8Sg4amRCGKD5kBKW
C+FEpmtqH/nXp13EOLC/CR9ybPocNbMVOWXtBmq5qd0SD9GjCvTU6+1XobDs
EPu5f+yrbTlxRSOofMT1LX4+bqfjH2UGQuTrRQpd7wmSDy2LUMZItrMDq80t
xJcsCXv2kg5mOqbG5acp+zDHlT92GI84bUwS5p9CB2BkzHFVwz66Vol0/DO9
kYHpSvD6vEQfRHZRAYGIwQ4ClqMeBQ2WClBzRoF8o27iH6FltK7Lp8rOYJ7C
PGeg3q9EjvSSz+bKSFAiAq8rAiixQ2c1fY2pfmJFzvd5USQLmiQTPes1X47w
Sg8V+G89/ux4EG9t16VyPqUmnjH0ISrQR4Q4BEUfd6BH9y3RE45wRfzVoWbc
Pm/oLrpblfWu9RsgSYqv+lCoxOfWHnBJAa5XpNvI2++aeJ50VVewlf4smhgw
geiCJplIs+6p9NSNWmN0wDXgB6COk52x+R7LO4Sk5MEX5Mnma6uMrxQ1YkbN
2kJ88Us2clqnVrw9Jm3ZDTkbHpY2zd7xfEtIIju0cYDkkLq7pGXZ7afcsV6L
SVXhvRkI7n9NP3b+NoYns0jebt/6kkMaGXVnpVFZ4qgSO5MOP7jB6Z268YsE
GnPjAKJpP7b62rcF9RJUQiLinZuwb1hvlNvjSEw3+f+4PT+pI6G7sH8u0kWr
/tQQOjNJCFI7cZ4ynxaXGW14pSkzpK73GTwGfoDuIUtau4l3TdvgJQFnBul2
wiRRCEE/pmVZ5uBTytDBH71k17ATgW24SbF/4IMlD9J2C/onBc5gp5aC0emp
WEoUGS676z3w019bDdSzhXOYSxjoFoSwBbeVbeXS1nG9sk3dnjE4BvAl17SH
1lngV6qwmbVsOrDvWiSo51vrKV3S7/qw6SaYOiVxowXvcXZ82IPuP+iXSPOO
vQaK7yMk7NE2ZbGy1o7ZehQjdwc/GSKr6MihQiUTPkKg9srSUPBRcDcVtW8F
2Zd5M4VjKGEd8aj8N1TwllSPtklu691MtFOKrdSCjnhhZXgGUT9+w8v9rDj0
ACOFFW65aSomLHeOIFUgTOh1X+wV+bsHwkpGl0sRpNTeGAQYkVDQAAmhI9Mr
uVWR4YL+J2g69R5p8xPhANuBwm8zmfGgupS0TdmmEzYt0ymtIbS/C4toPaG6
R/e1hjobZJgJg7jMkeGGmNtY+76knHZRK+RE1J2qhe6eePF7Ee3euLvESed+
2CV3Ld59Wp4kQiEttudOiA/aa79xcW/utTyQ9DgdJ3gox+J6dgoCCsA43aC5
0gkTb9PDpS/v7K7ujHH9nhgxsaFWpRC2NZza413+/cOF+byF/3c2lBKPhNDT
36rihmmFQaGdjLh3kxPf7rZmJlasUXm7pgNdTl+87I1KUru9NaLStU1Q62cL
ESSlygAfW8URp+Q4otoDWBbBk+03FboZbGWPjUR+bqGSFgFWucWRusUxRQji
OK4JcvGJVUbBPeSsnCcEXyNm1qvomabqdZOMpx6pv/5PIZNp2Uk4bdlqAVvr
Kh7m8mcBEPSJ5yghRg1NtWcQX5w3uQlPivUFMJc96mdvW7mup2JBfH+6i+Cy
/cItQgCS+zJeu2CpMQZaDoZLY8RLir1It9tRwFz5TQCCyVcgybxBs+qitPYt
Hubg3BgBwC3N4aZOu2YajEDMMM7wOeu280G2gGpKVTUT8O8+mI69Ff9SXu3V
Qfphc5Sf2Hg/6Z9Auo2kyHzBEYrWIRRZTxmqs+LuNbbLgZKASS0q+/oMoPrC
ypQx/93ODrRKd3LH3jAdV7s2DOr50BUHZkiwB4PN6CQ3ODkSN1iHINmNGwwJ
iC01ZOq4ox+MHPOTizG652rxQS6N+Hj9Ld4BDYMSMDwpid9dBJYpepkXgLAq
inr1szgL0ZbjyFzX03MVcVJw9PrY1bqI8tOr9G4YwekuOqMSrWr6w9K9rjp+
IFMee55DfP0nSlZKBMhqYzT8hjJSGA+yikt2O1Q0B4IXwzgaaWQfZsLyaAFb
XBuaS+nbU4Hfl6nI4nLWO31kgqK8cVi+5f5TTM81auIXCpKyQj/rwy3SqAZd
O2Byv+q5ThFlODR2DzhktwM6LClestkmAOwpxxdYDf1mDj1F+NlFgCWigvUW
ezRFshhYnPondv46SMHnE9zBNS6KmJ8mrJbVhVwtXzHMBXFC+b81HrAb5Rch
8E80DY9dNQ6pD8NkbbVCYvVnFXqd9yZWioAm60wHOKQjA5HTq/KKDsK1of1b
WIgoSxvKIUu5OdLE89Ly4nbzmLfLXUoaH0usYLj673NDMkAtTC7Y2TaaRUyl
YAmBofxD3RH8YEav/lDEMO35oT8HJRoXy18zSovXv6WWRx3Pn0AfFZpI3sF/
9m9fhe5RaxaNm9sHe8JLaZuiwQNHL0vxRdaKtR1jdnpVkdQZXdRz+JSaknKZ
Nsyl8Ip0RGoXheNGe6UHKubIJteNo4qdjfcNXZJ1HPK+K5NQkjievWRkbr06
Py+OI30f3EFPZCJISznGdWmj1Y/+67FdzYyoATxQQQuvedQFzlT6Gji3u4SG
25/dLmQRxY7ajKRqoTIbFOjBKhqIHHg7LU1BOS2n7TbLACZdNvcfMVZj20Se
dsttK8NQ/eUXfDnbBHg69nwoD9sqsu/66n/M6n1DwU91XQpxwH7zSYTKHBkR
knoeScKXZaUMhiOWDsHvVqPFdmvptQoMOHVHik5cFBlF+BjzZXPlzvcuijZG
2PrUG2c9E1IkS+M1vYtK1M92APg3yBB9VAev/OYxOMdKeU83GWuASKNaF46Y
WCUyXDnGjrK+gpbYqBLKLNFND9MwPAlcEK1n1quNACdR7kMUcixYTW8cyJp9
tlP0TT+9BhTfZoE+P6GK8z8iJ6jc87TR74T7qBruxkn+PeOKoutNOm17LC1b
aO0s7Y7v9EyP+lPHCeG2zA9SLzsSQzPBaLbFfjZw2FJ+IwhNvbTS3J39Je4W
opCK4z/4o1Gf/3Hkla3jkjnTJj0LiYBScqIU85x5wFb1CXfGp27EUHG1TGK4
S4arKD1OKEKQ6/hPGUfUcFEYG2eVXBEWHqIfwC/AoZFgyufQJi4Mv+efkNfp
IbnqxhQ8Awt7fV1JvzIGk49LOh0JWgRrYHa7QRPqu9a93Hd4bPm3NCdhEI8u
6dQ079Wnwsq+uc3oysLAG5PXa/yWcsqHGmbtEri/3PyFt3NBOt8A4xL55yG6
Rw/eeK1E1RGqfkyVnbcHSJ9HsbCLc89AKeQv9yIvmQON73sRnrb0P0cSw9fZ
d9CZV8kC7os4Wl5s1055uJjrPMBbgAocjybrRHJ681l0XMb/1I67KN4okel5
JAkj9Wdn+P5O7ejGr7eQbC+q3nltCDpf0L/CXDLywldhVSlUWtgnABV8Y/23
X+aC9QOvturZrLBlaQhTqTcISjNjZc3grhNjAVcEQ6Ysv8MW2qkHDH5IMV1c
AD9K93FnAmp/k9Cy7dxjwp99xUUy95SeqQljzB6CKlOqyqGJZMhjNOxByF+8
OPlq1duxfgEFbrWBrXlmGRVySjMuWo/3U6K/4BIyUeDWYuC96sfN8UwJ2SWx
GNq555UA9ja7sKebBnykPkDQ7+xT347U4SttnBtKCLCkP6IMutZQ05GjTXsd
J52ZKjvCquaMNjWWLVYfa4FXMyOSrVtHWjC56NznODrZL25EBNftEcrb9mAY
ulLdpMY03QnBOGcNlVG7d3ZOz2RStxNDhH3US4soImKBaV8N19F+k9s4uN+o
aD66SjEK+cqghqlpUdbYhQRgHqvfg56krVUFK962UIbaijCI+OMxuGuwlFdl
9Vn2EobECoohK6Fya0crdMWknSgKtCoTyNriCSOasq2X7sLm1uHMZCoVI1Gq
h0TPKFdKMBz7yTO2pZp5R/wYIwf7O+NYGq+z0vCMye1ZqZqaL30exCYDA0Zh
Xj9KTTWs1a6yK1UcgaagsC9mBWAaJ1TV0+6NAr4ntEnyQphQYI+8SCHC5+8Z
dYeFrj2kdlu1D/zhlhoIsT7aH4HnESJMDc53B5EurAnO5n27NF1UyJabypjl
nT8utYs6rlxGW6KSNPe/QyXjJ4f9k/SHIgC6CWkIBRKjUDf+mf6wFHN1rHBr
tRhNEKwlbmM1PWWEQxV2TV+DQ4XP+etXGWwJkHxgAftXUDYDfu72aOFMwy2u
U03NUdzVjCttv87rnpp8HxZ3qc+4scNcBlx9KoUDX9YsJbk6ziC78csMYChj
qA4/vqVE3lRHMdTn/VKs35a+lyJp8/BpOrmYdClAtbBdFECs/G3Mf5uaWRDW
culqxM9Xy98Op7JAYXMjiE63zmGzhUMZ90CNgdfpUQHqwxKKqg9hsiFeIBSX
LL9Eb9yzccYKnMVY7c/uQK6lw9HeDRf5IbACicszYWojVknlmjxDmY+aaLW1
WTxAvIlV6bjyuvLnm6GlMV58ycyUNNVmrJ20QIwNGy0O2eVmfWIZXLzi8wx9
W+lPOsiqgAsRAEXZRQYjQB3gN1/m8XGVsbNK4r6UFOlK8jijdscqBhZo5ISB
koRXQ0L9Pm+MLSV74AFBnzV6oUBasZTTtvsPgwu3rCAjjZXRne0DsPfjyh6x
zufekIQ5/NCiOENw/e6kocEWX0iuLk1UbDNbukOLCkSzjKWTVIX8Uz/Q3XOh
5L2FUY7Nj9uliwYiEK/m8/iB7PdMy4kCCRGRlzB0nfDVk655RBHn9VJqjfXN
mV0y/IsyMUj01PHjC1Ur5n24ndUMKonyrdtio0vxBhKrlvUpgD3G2yID2L/n
tw/fT+vu9XvIdl5s0C6AJ76QIEke86c+w97Go1OL8jq3a9sfxDAg9kErkgrZ
nidgiA0npjmAntskhKuC4ETtFc4UIlsnhfAKIQD1j8lD724v6ds1BVBUWOl1
ozRjJSX8zI4EPr6TG40M9tLM/uzjDaUyCLQLpAo6D9nmSUH7yL91MUjozDiN
lK0vNkLXmrp3LWWsbSYogjvefUO/fkTgA4cJvM4dR1O1/JhasnUeKt/2PSwi
iBXH77nz2fzNRnW7wCVKEi0BxMmLasfPtAynFF+7CVQAr3DOCHhHwU4MbI8P
TqAP7bcRbS3NT+2eQ1EYJpbsRdj3V8X7Lt798s1HPz+2w7pIpAXbgYdSJwF6
3bN9JMvXgb/LYox06ePKyovj+FH5XZoPV4taHaJ6e+IzhZCkkC97EP7kEwnV
hwL/pj+Zt2VHvck9di6/HhFOW3ftoKbiByrCW+ywv4nZ3JKujSXknYDEEqhi
E0lKEyyKJnvHyfk47Pa7Ci6wv77xwjWgYL2txzr4jPC+Kfz6hMqhUSX5A+vD
CGf9D1OVJraHrwtLfQZFM5ngXYt+8duil8qbDPAKzbhB1EH024FtNTj82/BW
IEYUlV3DAp5fi6KHzWz234pSvhyipCQTgR4AcogkaYAuxg0ZUuuG0k9g/HPG
3pJVkEyHPmjVBMyc4VUXl3VkirhAk+ZDeMhUdlmdbHKtonBIoXaVqwgi3qee
m1RlnP1hl+vgNIRH+FkoiN7dXo1pxi1N2WZFRnMpe1KzYkI9DJmAllvOVUx/
uI2+X/F34e96BkqNwREUlicRJ6BI4SP2Xu8KAgYnYeSg8eeBRnjrc3Oz8h7i
k1Armo8mwx/yIS2Wk27nHl6JHWcpdB2JqT7A8Mvg1jdFAwz25P/CfaCVTZxT
1qp/YmhNOjcNYBuREj6E5FdZonIjoum12BmnScrRTEzubs/87hcOWsdO35rh
ZWUGgxLilzjb0ki/4BSjlf4G92DwSG77PxzYICjGg3v7MU5kPobYqNDUgpyH
7527OoAFjAek+/MeLJDrs8ROw9+yyOMOMWzarwvRy3Lpg30PzTkre/+wV1sD
4JYJ7ojBPmlLbUCkQOcb6V9izyJryPpzs89wuiZSH5ytkdARA9as3uNMpzcJ
opEH1ZyRsAWy2L4/atUEC76NCkXe+4T/GU9qK2q9+OVZ+PmSgjwUN0fq3k2K
UwB6KQv15ldWRNvLgBzzBQpk1jS0wTqLjfuyZuUoGqXZejhOPfB6LRL2T8V+
yAKolpz0iBR21wAAS4Qqqyv+EzPjw5x/0Po5h2QebO2iQxHlzZzgmlUPgyJ4
4HdBo9TPdbMwAIoS6rO46rjlGCGkBtw6xPzQkNoZW1VaQEC8mFrBlu0XxxkL
0G8MAHSRdIHrxMC+d8mZZCKXUMSpsiEcvBi/n7659WClhylWlgE4tP7MOkrw
mARez2/83FoeNtU9PgA8OSHRbWX4x76ETseFLjLDnO8wXa3nZfGKpYMuZ2+e
GtbLjAHoE/S/8DEkBjKSLyCft0z39xA7pD0JReDi/vLHINBrpvzMjUkglp/K
vXXiS96l/DjviHAtIBfdXrKk/wcNepjYaMmvyF8Dx66z/HFD7YY4eq0Fl5Ch
hSD5gPX5dN+5keeCyR26TPoFfaxQ0awzLnyvcIKTwWUQ3x7VBZ6Fp+ev3jvG
sqzIzJGQfUps6f4aL04n3jtxf6sA0iLD9JL5Bc1kroSKVpTJK9vpmHoDEBeR
gp6+6kjbiv7i/jzVZLS3V3oZwbJy9SXnxLrrUMxn1T9KItXIuQksBvPpb/VS
+5+6PpfPXI5MYC0shC6h8S2ITc/MrurCqq2qyxEQDUPwr5o5qBP2MX+wQMSj
PIkv/j3kZJMIT3JEk/z01MpkM+jWomR7YdxzxVEHFl17k1wNr/rEOxN1LRpT
WfB6y8XGGVJZJvdPbYX2sU9bldbwZKAXBpHHs0XhfysxL+VoJ9m+9Q4H+7PU
qJHIEfpH5Ibassvt/Q9BOlxAzCQgd0KoLKe04m+AqhcniuzIJTxM3ya0q1YG
s69ZI8In5CrDFqUnJcmkLaPPAhNsR8IPj6mLtJD0rNut86DYr+ObWDnt2WJu
PiLDn2/bZ+5IiS/XuWQQk+XQ049hunwfHkOae48xo571l8XKrAJ6nmYZopZ1
PqlBe0FeepUxXEpWCOpheuXXNrk+MVwTuNk/+N9e10cGZ0a/jEPSkxU3mipk
sLD593OtVH7SSew2Dxvv+TUPQSyxzQ1OjjnVdeINFJorSFbevZCVsRteyI+t
qPUMUULnNhogSowJtge9g6cI3Gm3lMschLm78REPQJiqlBZFyyUIhr8dRTqb
qtCd0mKyzzwMK4kGw9bd/ybAZdHFF77uT8P4C/nqU2ARPVIjE6e8RqZkyJp9
EyQQIQLzrP0GpOM/dfvF7T4P+ZITGDMCgbFzIzvm34Hy9CeUAjQT18XKO0AG
ifVppyuiPH0ow9J9PkWgsq5k+IACC98b+bwyISNi+EwOTX36twuxNCyG4IWS
smDS+pnd3umyqgy/Mn95TQV3G3StwTuH1wJJKa6b2EQUGHBYNL4NOreroopu
gERY+XZxMplPKrXcVy3+5L9SXzEXqag66CnqMfmJ/+kyCFffR8r0zxtDJGTz
j9tKx2qzViRWv52CJJRoUxN7AdpSjhoGyJwXIBvemgXdZJK/+ca51ZBsVBP6
wqx1vtRv5LPzfiKrs337j2cc45DMlKS3c1r9DqPBiMUiFtrYRglY1/4QPmze
dMchpz/KQU839kAilgZkuc4nu2Gz9PC8JM3qviKSY61C/ICX77i6PJt/wS/T
HI2XuqsaMdlJfWeUxzLZ2BYELB2AnTkdWwjw9fGQ7ffA8n2RHCi5G9Vr6YVI
556xrpSHnx4gWoQbPrSqoKvX+HGCx2hILsgjMGI4OoCI13ghDVzJ2jtt2cmc
g8SMcOmUG/zQDBv0kdUi831LKsjej+cfMGfYSsAbEql95T6NDTdXV1BEN78P
ADqoKgF+6Ki9G/qoU4DKng/oG9O8U+ty3EAhu+aBQGFuRUdxb2w9vQVoE25U
ya/j56nCHmxpY+hGjNfzRmxxQRmhGlHG/e5sHasJJ1PVf//qRlPHEjmiRrz6
ZhC0xXpn5xrInDNkopo8/OdyiK6zrlPFHwDUwa+2482Nn4eqDXSQqK0C3ejJ
3Gc9F4KT1EWEtbzgr8DzP165EJVCD7lH1J+6YSyaB4ENcLwcmPlQX5TieH3C
p8A8V+9135jH8aZ1D2Ic0YD6CeiY9Eb5FCHvMR80mO/AHDNvtKQhHOjiQnf4
KfW58y6asSExo52/FWoEpQ9jctyRrmzUhasxR0s3j7fyyyTiL1Hn2lEtGb7u
c0c9TPmVcmb2eRtvhypBA/Hsd8fJdS4n05Y3RgvgwKjnwguMm4ZMBgclZZ0N
jZeWFPfl5YK9ixmZgl/4OQFe5anC5HdifNIH8LPFr9EZ0jJeNqfZuQUpY6eN
tQP2VCE3fnAyE6HIPCwMlMaVucVI6nXoAMcQwAX575PhoRfDYKaue3BlJuLn
6rIY0Qp7j50ZQH7QQnJ0BzRGcdFdHYK8quzZ1A3/UF1siNyYpQDfKhiGUy+R
A9Ga0Ka4WDW36qqwnTBT3CLM/oN5dj7lE8vHyFDJrIB6fVcAuaN10Ehm2qYy
vgyIBmThKj71przIXQ+zFM1M9Qy5Q87NXOMSMfcYld80LU8VklZh0EesEx5v
YM2oJouE8wCD9IaC6FzyjPWKgXJuCl1N+9i87qbluCwkpVin/faYopsbASjW
+RPII36ziySJaDomkMCW1+pz/tYVyNKFkbGGTxzXB4A5aK3U6pb5a0RyM73R
MH4tieaKea1CtSTj9Kpyw/Lp67+8OVu9CRcaASvqsDp/L2JVBJzEYp9m+1qA
wjYKKr2gDYybOixYUlzoJZEopv1SxHfEGivDMRwIGf4bA26h/FgQF3Lx0YQU
d0dIXWVn/POu62d66VFu/IPyoJhtQBO6PDTeB51lG3gAwzeDne0b5ZtRrT3E
vC8x6EzXtHAlzQwUOwHdWbzYOqw8xS0/k0w0WwNVm1UV+A/B3+7db6D5J1SO
JB/mSJSOoKxktSPpXt6ZM93AtyaPefwJX/0ke7p2G5aoJTHL5hLIqXpi2m0M
gqyoZ4uYHgUogV7fbG16H1GybABmj5ATMcS9GMNVWp0PGs6Q7cPCrnmZWL4N
MdGXr1RU6ROaKJR0jbHL4MNo6+Ml+Elp2IgpsT7gC8+MSEKemLSMVz61bd0C
H/wJOiBmyC3XW747dSNA+U1IGwu3CrwOsRCL320grQl5FYTEculyk3qNyOB8
9PcVOpCwtrcNFWfs7nJlYXF51l0cPu2nh8cxMt37mYWAqLOE0Tel6Z4O7iWZ
JAqVDDMWOAHIbMjX0DuWFAdThMUgR8FvKnALxa4q2ApCf/5sxndaRi+nUAdg
9H9NNsV78Y7GAnm8f/P8hSly5nxvHGO0VwtUR3TsL4GFQdkvm3xiDwrpIZQg
pcXiewQauXmXk7zb5TY+Kz72u1PCbiIzjWdeYiGXVuE0V7NpSK/6IDqhPLuc
cZX3pAbseLmTatu5ZO8zdoHPDqrNtLp51dlfnhNZsdSAeCepEDYEAqfIz5d/
fQKxaFYS6/v/yWKu+CP78cAOKQ/j9E5/Mk2FzC55vIKEJhTquvtlQyWcKmEZ
WHnKIZ3AvYatb9WNRcS09J8sKPuSG1ekT89fnFJ0am0r0W8RGDiG42DlAurl
qOOzH0iIAWBpbB08gnfuCQGoLReG8UdW64GF450/RcTknMTs/iN3IkIVm5rb
3yUhGx2NuAJHhgJ4p+uz6A2bqht39of1lSbtBwj0l6iX++pBzCa6mjfOwmcC
82evSHGcniclvVfTFqF5f6wpwRovA0FqshHAFShn1vgHJQEEKK3m/rUDOJMy
L1e9IaRNlr+avwPEXPLqE6glAv2gwhD3Yy653fWFUudtLA19F2xpKEm+MiUG
XaLtmIxWT5mLLJCx5fd2pY5fG9yWvuPzh9TYiS8lULcLLsTNSY8q+SZFsZe1
TmTaHnyXfI3euojMLlnOOscJkRF+afrJxOgR04IlwoY7C4r/ii1fR95PVT9x
kvV7JC45IWUA6/7jpj1d2nIhIl3YZV7SdRVsGCeOD9Tp5X6iM8gzGz0KARgD
kjfM+9u64EsBphHjVPV5vCw6FekZp/swhtHVUIeBg75piT49pLzrQak9O20H
wVbmtHJvguZGsdOAZyuUMYJ45fRIzfOGocDSEJBD7YTSs3GIqY1/Qf/e62zY
xgSUm3DOR+8+AuLwgYEaU8Uce7pIKhgcPYE58ZKFg4lDQ9NwLepTMe/pqRID
aGX1guK5BXqHxzjrZ583vEHL3/oMG3nXCpnQgGOEyLrAvw3IWFDEC3HiVrD1
Ym4syQPr6qiv4IY2T2FViBPQ/tjfk6vgF9tElZQje/7ykWonzScfeo6qKGl6
KnY1pTuMdGOyynpOt0zZyc/4Pn1lGEwbR7Nnk/epW2PtEHsi00HRea6Ae5x9
Y+yyNOZVsM90yLxnP9JkvwXIVxJOMQBWLF5qe+jDgU0tiKGxWulu0LsETKv3
FZzjv7MhBRK89JskWEi/nyQ+UUEbNZtxWe4XhCzR6/oNgKnWWmzpqdHJmb/K
2vHdBig/qHe/96XRHRbmXAjmcuWjbkUXklPhE+OlyoQ3IkhUnLW7Wnt61xrI
ThFn+PxDx6uUnkXWZqa2kMF+JeQn4uVB6V2A+bwlG5F6KXMJJ3ZcyB5JKXXz
1V56ogHSegmtU01bUN2CtcD6NXcUnR8pILXTYohMcYD3FlYBHOuOYVDFXrV3
uas/qOj17+2EBKzsle/aCxcnWERTAEsfxTb58nkMWXuGfKFi7VU5v0RYyFnk
u9lU1jLCc+oyQOCKQLvY9Ec0b3tovp4lg5YyY8j5IFRppb4/bJesIu7oCHo8
hka+JfrPhpGEmDeF2Vy7gdDlaJvQzOyIfHpQT8k/hORbX+6tZ0Ps9DsI3EUu
/lXN2CkRSqiRAcCbRW+DsA0lPMQrASSqnU1IyrvqZodj7bajz/Vyqp8Wr5ZD
sSWyAc3+QBwrLJ7T2Mza0lyiZkNGfqXN6ZTLQO0TNFv1NaWlZvYfCd/T4zeA
Ny33H/2I2YgxK1GTV2XJa48eGrwm5l/KVBDDsH4mDUY/KSp0jBKXMHGYzXBI
zLkZLY+g5MQxXJgAl0K6GQjtddmqFKpHdgKGNyxFrRkTC3m61gu/Lz5RZDwb
uUSbZXgq1FKnXzqcYeyFs7aE3SYjcvly7h40N6sMJtNX66ujHpdHUTxGuc96
UR9AaU3o5p+jNoiTITqIOnwi8RsJxj5xb8lwto/lpimuqHM2bgHvUXgNLDNG
3Zzb3Mxa2dMcrv3KHU1oH3tJvJhFQUTP+4ULW7DakOf0fLggwMGE8OG7FaX7
jDU9T0vBkMGp+F3McYQqrZM11NNOPzGdYRZxPzs85lJuUWW2gT5gfhSEDyG0
gZZnkD4ygCriwc1Cll6wwFKbGkKwa68mmOH5Seq5FYkqSbRyyrGdBw85n099
PKLkgTw8QIb4IqpwKUepDdW+FXlGhVQZK+9c6JTOed/wKCJ06J+wmP5cI47u
DETzHwZSiMLXCOtxePJRD/4t9hqjM5igqE1JnKH4jBd0KM4XaVcRcHw6GI3d
SIG591XbKFgpnlIWG/Rcq+D75lSsTAoSwcEpO/1VZP6RB2QTFDhvwFi0+uz1
CD8x5vB2Fir7pYyUseqKKBaG1ySMFJ4QIh/9YKteEaDpoWVzhtA2kiPJ2S/X
TKKlyumZXz9OZEsDkGt/greYN/6sa3o8kIgQYTXogagDEg9ti1hOQvvP2opm
53epjb/E7cnukfXfKs1FLrfsb2NahvlgV1wDRkrg6Pt1XI8EfnE8k3U23wc0
IzNkzOh+OCM52wqqThE6aQIUzXjWKplY5SEYiVXQZrdndsdyz/qZ3zKH/Xnr
ymulqiohJUOkVTcbVBLG66lQMO6AYfxr/H3yDFU503k39NEtoQH/xQml+7iq
+INsqrgF84w0MJpHE6rmkDKK2y312bdX7WrTcdWCod1GLq6Fhr1s8vAYohSp
QkSFPSWLavL89OIoG8r/RWM9S+1v+aNfgZMO3/ChX4Ser8dFi85RM7JWuuXV
eGhuyulb7DVX8Dyo1iL4aIz0FOyJJ2iTVnE81Tv2NfQiWcyJuSgXTcLP1ciY
Ersb4Q65ELeFxxGTcV3+yU41hNZHqBDTOyfunbk3gR89lhD+bRp8mJeosn3L
QZw6KZgAqIKn333ELUAMPIk3k/k/wUrG/+ZP79v41KfdpaGvwRWsm3zzoOgd
FuYqp0l0JF4mMmaCL4HFFyQ9gF1qV2eGAkp6h79aGTHAAJYvBtr5pYxshlII
M+9iGNPCPUg6dzzDGUeDYjjQVvJ7Fn0C7p95tCFpQcyNqASmqeUk5hJcasya
XEK1sMerjGCyjxfTg9tdMqsSU+KvqYaIDvTZhlxeBXDIZB70m2KD46cNAgK/
DizGEKcrECgSqQQQJFuUreTh6fdQigps4k3HJuxXP5aTj9B5LJvP9U10Ifpr
hhR+uBMsYEZALISixw9JcX5+Z1d9EP4glEIDkFvfy4Tan6NJIwo/1aOOyVNi
4afRUgC94YA0H3F54JNzYSUTj5Pyp2rQUDrHj0qGYzeFGD+o8NH6duQGZvSi
OVHw4XRedur5+Rx7rTIt10IkDl9feFb5NU+ZaozMQaSvG0sIljAY5BK7Cb+d
vVnvxbldBQmd0g+lDCmHY5r0xMYnpyTBH1gFaqlWIfmMdAUchqhXXuDf4NSl
La+Ps4brFEONxSkoxFYydk+C/zpyVlcliQ6u0Z6N0HhTLAOQOEppGSpiYAfp
PfIs3I/SjmL3P9b7fO9K+qN9dCxduDhKZib7n660Vsdyl+dfC3bAI+tDOkG7
YE3IzZKhEF9Yef3InuOPTOqahHRrhDkGka6YRYEFl4TOwIb18gOkS3t1f6zh
ZxZTOBoSfmvwmgIGZGALlndILNZ905fGlGxeARToGuvm83sSN1U345rcX64q
QGT0d33Q4TFsQarFWkEA/+L/+eshVwqqGfamXdCnDrE6n6T7V/jHefW27WOb
SkVp7BzwfipEXvl0yuplV4lyhiidl6gMNorcZ8ZyfZhHmBv5Obp2NylVUfNr
9y6dc3RJ63MqixtP9em8pmYedUI2yJ+dGCdDczvcbfRTJfU5j734w2qfJ4Q/
gWNaEY9E3xme13psbncshDqFfwMheZzHqsfkAQKBA0ZPjq+QP/fBJvTcsn5L
6Kl1j3sK7fLdt1lS4JtsRJXie0zpytIgPXysF3w7BpJ5viaGHKFJnzt8M5Nl
QMZtJyyTQ71wLHnQ1HAM2AypPJbo7kGLgwOz3S2/kE6HczDgHzxDuRrbA30l
7D1AFGRM2TYtCGyc8kKyf0baakqkx2KySxh54hu9P4QHTejARS8u4qO0xxc6
Ny+XGrjfs8Y/S9SwYEQRQBdHjFLcZ0qcv5PUw3dXyVxhbCvR90Y4PszfoCrI
G0lnSn52h+kGAJyzowGp7Qemg0d1Gart23iSEgTDRC+p2lVlyDWE8KBmZ6gQ
aGk2SE02dR7P0EPQbzpRMBbtASkUWtfBDMmdLMsxOPEcX5pj+YOir560HROB
M0QMEJ6cYGVuXdeoIuGHTZXTEbUCSJ2tRVYu+39PO6dg8WbX/tH0AaOrIAS9
fo3P300GH09tfQbOFW8PfAxdMEyDNlnLglM/RdIbIrojRu9VmIYZ0EnzLnxC
wjOa/bjJ9ckeCvh+0hZ69SOak+5Apy3JNiGcE4L+ymvA4TtX9dZifsrIDJ7V
TvMZLbhEQOsmuxnHoLp3ogmH8lLDVLg515gLd1gbcjWSv/dnNaGXpdEBDn7l
e9TlvkKQF0y7rTb5QJEOgygnEua6kAu33T0Ay41/AuOCSrtYf2SHwtJfwaTh
bxEv7xfMCd3giNitOxXmFexobuzv5ufEEt6K1VnBQRjHkdGRRhWJIx+V02WG
vAqiyta8IRXADBngw9y9g/2b8qvGNMYv225joOfwGOpLmpo3IjGew1SjlbdX
pa0OVHDEgNtIKw3F7gnePyCwFo2DybUN6A7fVbpHdd8IEq9vjUELSAt+ZPNR
YH9RYq44KvYfgh4sJ0pBMxrpTBerQMjhkyftDEaExIxxpNJZt1N7mfmLZEek
ea66JF3mKuUcDC07belK0YZvLVQlNtWWFPv1mRKrLMGgxzz8y4x4zAHiq4mu
Nmu6YW6ZwzTwD84PKNAXWvO2iMh/vLBZ4DQ/KG8b+fwyBPddauOMYWONb8w5
MumxvzUPLZ2S7jtk4Ib+tXIxLE1b63XFPqNI/dEMBT04LDOc+WwPj6Yux4m1
PO33o0+XwNU+ZS/CNewNj5E01qCPGsZB/QiVu+kSr19UE9ZkXathNcBslblT
2qwtSHFPzz6bodnEIUtecVwLbx+Bqu9nAoj+JAuB5yeCEEZV5VBtufG+gQ8c
X7e9vQft22t5Gk2neOzq3aXomqEk05GO5rQVKRv1qdHLPu6t/HgIJHfWZ8M8
j/mrQ5fecalp//bzIQuZzNLrY/MH/7iP5peNGTdFje2CXvXevW7Pjz1YydXZ
gh+mPWvq4CrRxnSiWslJsBljCrwH6fVHep3I1rYhpElho6PCgUwgM1oYieJu
mWuKBpj4R0KrSHcBSCgNi1UOw/RdobL0egJpvePaMoRkYND+ABMK5oD0anPr
F86Rj/6xkozBAE7ZU9BgJgmLRWgONohzWuPOkRxmCvY0i1xMbz//1Ib+9PvK
HB00gF7SG5kuyKInKDGk756+O2/+HYr2YXUp/WsWaQtfslUADhpeNrKSa7Gp
yfRMpqB0emsCgyU6MtGqY1vT+FWyebIRZ4bXQ3ATkDprGbSQwg3rxEyaJ0Ev
6aOVF3byBufdrVpXEticUkiCsiZ2l101htZco9aFuzpJdqg3fwayRFafoj18
H/XkE+CCDk13yME9qal1Tcsvf0GwmtXe9MQBoznMk9JC1LKo2Izmxi2EeGw9
ljkPyrV5gNirpj7IENe4W7VCy+QVG+H9q13lHwlob7GE01I5CN/vrvuA37Q+
EyKVtKd1Y7fh/phsCcrxt6sRfQE2TbhR7kaFY5Bczy2kwaWMcTYE+cAvSdZF
K3SWkkQo4YiK85dad8O8oigodlp6wxrbG40vU4/KWRDm52dbLLaOqzi3QKfh
LX6JGK9mJHDJ+mmoBI71MOhp/WUmAHOYi7KKzC51U2L1xdm5cCDbLijuwyFL
gpcZefRD+LCLMDI4tlfNnuygjp4y+uE3Gon2Fo9ahaloJ57Q5Id3HSVP/hIi
4uu/gj657nKDbWxddAwIpOhtcNGJR4DGsxwfdXMt39dPY4e5SBB417rFMuIT
wbwmAmEw112f9GbbtGA35KErcc67JXsMmXzsq8fWz7L0BkXKU9Aaz1/NMC0B
lOYhMlhujQuhTrP9kKaux9TcLdoYiItjCQUguoR/nDVC1foFr+DR7CdeHfsB
GE8rrJYojr4aLUffNdwOCvSWYO1UYI01O/eSgMUzOJLtHjLmYdD4YDAFHMCf
Hf1Rk6L0bj+lbNDewtzuJoMmeKiPzv14SScq4L+gIBIUV686TtX7rhB8MLWB
iyYxNPWfuFh09BNHgPOXBefFB49xjdJY3ji4m//TViuNarquVpciEik7cvJW
hdBy1mMrMaS8VHLsR03FjvaLJiHT2wOZN+I3gX3fJdMzVfPCQHqLWDz3FdcF
UCD4nbVQEQaltxSM/+KBdHzn2AcsBra4cSkpEsk5OsbYgf+hD1HRbtnfE1ji
RsXbl16h7d7AJ+qTuBmdEZeTcKQaGkyfePSyiKoJJquWkwayLTmESBTZzGFI
YcFP13VfCs4Og9uYYet3AxJtZv8g9PWbNICc/2KuwiRnPVKN/uO6sqQNaLAL
HKuQfiiYwLeys6KLg5A5mCgB31QahVxH370DWW07tXkTNURy5G0peapnq7q5
nnEHS5UyJioGWXqzO4Ru8x4HRfMfxKEG62b/J1DPv4/1H+OWtRSNQuwuJnKZ
pgA0jU//G0mum7Z4Ykrk2d3bAjOVLJs4cyvfY3MLF7tdeFCS8Qxbij2rzcC4
NcEYl0fQeT0RNGSxbDqqXht0xbxUpeG64++1nADdC/5WFwv7PNGnZcj4iwfW
AoqVrROjlHTnfiOLLRwgTK1SOcIFgHMRvQy1Fpwv6gfa+LqbH4HO63G5gdoE
43f96uQjTZAEB4ILHwp0y0QBnDuUHot8rPxK5vHDOByoeuqpC2c0jKGx54jz
4JL6a0S+M6Y69+03Ht9mGYUo1mzrfbCxIEDtH2GQaVlgk1yluUy+VdDdD4WY
HRd9FsrpQbxNocMD+k6NmQpwX1ixeVpaCAH9FXHpWY9d20p1LhlnNdz77WaV
6WcV9XqPFxV3eK1DpGTCXY8LV9lC5vq257wcGyt5yAq64eJ0UdkaGx+P2XnS
Hu0cHSiY37hPC6Yh9AfdZPrB7QpJ8NOCgioJYcNAlJE7JzAuEr190QzuwX05
O8L4eOZOmC/IWsBSOZ2M45Jyr24QJRYnQAxLZnR+ifRB6RuVbFkRZTnQ9AVc
QK5ZnY+dHku6Aiw9Bxx+wQ8md/GHpbkCVzX5cww83jetPlkFgiBRZo7th6Sd
i4VNu1njZtvmjmwOU7wNJNb/72VFv9SmqyvJSKZZ3Q9ooyYQNYtDoeI5HFaJ
TCWS6idqm6uwyms2b8XFa1WF3V0d6zQitBgbnPoI5zS4yz5zE5uYuUcDBsOm
NvZbUqP+K6ezL3McfWMfPmO8ruxuX66hOF720HwvWR59dsJ+e+2LY/MgXETT
yHE7fhZV0bLWPYCb0zSWk9i3YCk9YEi5P2S0+9uQ6qhgaKlHUeqRijGK+3bT
ZF06FZI+/Sl6nrs/ruM8tdySSLbPd2KDL8uk6sKkp2zHQ2sfrc3XHQx9Bb8B
efaYWxnO+rszuD5/anoPQ24du0pj6DAZglqt2pMvLc2FIaqESjaBDgVGeeGm
SVrQvuTj/g8zp4C7Me0BEP+QMuXoWQ5/hcYiesFrqf912bhWVJQ3QtYVKRsA
C2rvTPZoDeKBUvMelhqh0XLUPN2/TIrgOWGHXSSsnFggW4RQ6Abwc+pUIipA
AhJVA86m5URIcfR8irzkkm07V4yKZWfnD/KmfedZN1BjYu502smUZqOOBwn8
/f2G13EdfAwFHe0YrgXMp/QBy+MBafCOJddF8rcmUT7yd1gIOkqcvjIG3BL8
rFsg2UnUNFpufwebE94aodAyUdk6BkNRIhL5mqA/BEghxZbxr/xMphqH51o8
DmGp5CgrkUWpRPZFCQm0uU9oiAHeiOp9f3euw7ESqNRt8zarc7AjhU+rLXFn
qjRMrABxTxcgzig7akFQZ8+t4gjzaALHaPPlfWhpYYhCH2fMUeioe7WuHhb6
n/ldBKjPmsdJU3LARw5SwHr2zBsAL7ZwnA4v08UqgOKtZxj7QB5ovCiwdjGo
3Th3dz5UwPFPp0/yWpupcUIFOZ0P3GwpJLxTJcVk8egoLcq6BCzTYZmg2U+n
bnQ5F1/GvVyfJGtNsdBLyKhfeK+vKHpmS3HCn0fhujx46XV2s+YZO4skcKA0
PPP1owwnZEBDETSv7HfzrSqCNOPKJMhX/LQTz7iCBCJzlLeh/DNsF6CE2rXa
IaEJmUE912WP9TRmwTl4SLHEwU5yqnhnYFpV5DzdNq0dnp8m9fheKxTreMRi
HdO78An1QuCMvwsxzyYgrJcRNIy3A0ROhvhwRTM8sscKqEaQmV6I01bgJiwB
Oib7LILrLx7mGF/Ve2pHBiITY8DTc5fGeSkCLnRQciRco8fyZb7ZxcsKW8T5
Hw3e4s+bbZ+K8Np9HDQU855fCtexK4MNJC4tHZLVrwIYQUeu7sk04cL1vrHZ
nZCDLzzCkgKjEIJ369HkSzqTDT1oEAzQJiFR2froiDo/UVeqzEgtoqWrLAH0
iFRbF2f5xxmhsRRxCkqcmDcG2qGVSgYgma+1PX0iHEsPySspg3XUGrmhINqd
Xb6f1hnyrygavKd5vFZ7JgXaEb1W904u8deSshh9kHaFjNA3HNi7JxmmFU9o
CBjvwKxUI+QyBTajLUcgIAlECTGAH41AnP8eWxiQfQCTp0YEiH0FmX0Fqz+o
PPOJw/DODdN2DlZoRZQ4IYFuK0nUx6uc4nfP6rELgWKcTxQCPQBHXCvFpbrP
M333GQHOv+Iu6g3AwlHLtCWALTvytYRIvSpDfaEik8epZB9YHabaOPy30Yp7
W2yQI+5pNFV+xGmvsnjTUIbUfR8AiWOaQhs19Yc8ckE+E00Ur2kgzvxudd6i
AEAn9aOYHetm4GjZ+/j2U/udxvk3J1NRJsFtezUr4WDma48HkJsNTs5EQjxo
0NonBK9ilC4wSTcwe4W6SsvzkbJqvvneNYc8EQaQCkN+nyyxyZGprhJ6tF3p
3zXS5qk4m8wZCioA5I73lY78WsA/LqrPVNV/pcalSyPKjgzHEa6txAEo5gbL
psLDc1MW7dvIqeTxSPcBT+zHdP3d8Yaj/830fzIEy8MmrY68Hy6NxZDLF8Ty
CPWlsvbYH+DAn9eJvFdeDBIcPh5RpWGW6pYMYPUDVu4QrT0hvSEmpSlrc5Ci
jjBk5NrFmz9eb/2FAQBpqPjBXTIcQl8VFrTW3yHmVmfxYKhIaFDhTlbQi732
tDToayswfe/cCxxBK+6GKsk+WNWR6V4z/bRmQ7SOzgrkc9Xfb0xU2viMrg4b
0ukC8fXdl07or8P/UbwL0+SoMDekWmfUTilcu8sZefFNV8XspWq/0cvGbb/N
DLwl3H2JItcXryamyXF2YVn0sLw9XiYDQeKO+3Pl0N9lS0DGsDCv+W4+FIXc
0/ZN0rT8ECOzCh4SnMRihiqhfxM3+ITTkL0BvcLl9P/vLEFMkSCfONiMacAk
B6K+gMaOTXzIieaYS5JXOPFzFb0smqr8HhHwmG1DPDIN264G+xLR3a/Ao5xl
OrBxTOkaDyl19QJWN/f7+855H+aTDq3DhyQR3NGexyWLRcdzM3jfW0JjyO0X
/ZKgFcmuD6d9BwddH4DCtXQYIPL5O/yPhTIq/uAL0ma6Q7p38eXYR8TbOP27
gfef5JY7uBSnnnc8Rztd8jHSHuWSlhF5XCLn+up75cwzXO43fBMGvpnRa4H7
7wFKQv67KFF3pH3CRG6LUy8cZRg2XRQUoBzyIC4/nUEPvqV/O+Jd1LPLRSHF
ZK8ZAN59RXTlLyx1JuWffkwcrhfXjM5LbJ6GlbyrJenv0XSvZkn+QW9v5JAo
H6Z63cmNIzDpFIC8aotnkFhV3bXQuAWT/WuUshbmFmY1csC8KhkScIvGFHeM
c6XQjupzbaTQlybWYqP/6uaSg/59f6F++dygAFe0nXVZJxPknlkg16akTXoe
TqVGteBO2ltNNhXNRkqaE6uUsDpuf7blDxl3GXlEN11SZtke/+Or0BzvzqwG
1wDsmYkOEwO8tmj5dK0t0PFV4GWFYfce1naepC0SY1nxwnvK2GBnI5zgzMc5
nMr3hClOlCtjJrbULqeHUKU4dY/WRyv/OiYbdK/l9CBWKLmfETd0bGLSR+WD
da8WNjJykP6BL9liL0R8fY5WwpzFw6Dh30AUIsSoXXzBiFE3HqxczMTlhHIt
HZ1cCreEMzKB+zgUUMy8M2xl3axLNWY+MhBb1ZI2OkgoRNjSK3TGxl0Mp32H
m+ZSI3ojjR0fcefJ2ZgebgussRPKarhxfMZOFogHjxxrJccsNS/fR2YaoEOV
UdUF7WLZinK7nFSJDfNETVx2Eb/aVwE7zLoWOEiILLjLdu19BRg2zD2aSFU+
Q50wkro7qmVuy9EO5PXRz9+qOnp27USRonxDPvuM9D/h34YQwR1uTRzKNtlE
hjTgZT4pgS5vrkDad37ndsxKybIhm6wYYcg2FWbtVfoOsoOSJFZR7YJyRduH
ZUMmF3J2dSpQs8rFTGcajgVaqekRpXLgk5S1dNmcjdeHBaQYuR09Z9wkJaHC
8iN+OgL6MnODXLgL9r+lJON68nVIOEse/1Mhy3LIQnp9aKWmyLqDKQ32tCeU
X3uIhgKdDMWLKlCA0cxiCYQVhO+//GOwiRgqqxqurXHcTzy365pVAAjSV0dN
Apvkj/f9SSY/qXyYVNThPQ3seUj3tq5SYstSpJNkNFj5aiQzOkoYj6CNvmiN
NGt/asD0Y36twA5bv039Ndjc9vKw03q1xbByM8Yr6eJkJeYyg+280ZQwCerc
pDrtS/XTAp4Y3oJX4uEmzDfJGkclgKsALLsbXuUkhUfd0FcXX/OhkFx20/rj
QxHFki5NI7QCWU/Gk4sv/y2RMh9MQ66nk3rYZUoST6yT4xuj2p7QVkPSb3mS
boRkKmKa76byjUK9R7ZqVJ4EOACZlb3i4pDm+pdGebEXtkAhsn5voBw9o93l
5pW3xS4TKwzNWLnbRLS04ZBNuq6TOrXe78R53vxV+CN2JXpVBM5RnpHsvDiN
oblcfThg6qzbUcosGMXwO8IksWOCHiDbEw3sGhghV8ykV+ZJ7Op1EoLr8mL8
86pJ74fTsTLD3pfZmlYQZZ2mwRVY62uqw0sOrpxD2EAVIvntQVlSaYZtiiJW
iPLjlOoFoWcOzNEfvCMVGxy+DEVGxfbC2p6Odlg1n2yOWEmZZEgcRtrVGvRG
0Srh2AK27AoSDKuDxrfqtI2NladYVG1mgpmiPqjH1qwp84nFkflV1pdGaKvv
RXnqn5FuhuSBBztihv7BWv7Aw+Z7MNaz+LV9KFR51+XnohZLp9OMVSRtN+AN
3BPAElxYZkbGVrufGJ/80JB0m2OU1cipK9CB+ijvEgNau+j0ymay4fiBR2/e
oTUrxVufpXd3Pr0IJhAC96s+HhWnINfKwPF4afzTv29rIhPobGpc3/ohSvps
mhreOQEY1DoN73X6Y7wdyA8OVqLj6lBO5xEFF5EmXPVzqjQimPfwze6G6Q9C
KLMP2M3gdpFB66jQ4O3LJBCbIB0NVZZsgV1fGwd4n57ll3BDfU96H4tFXdwy
s9A2jC9n7sq/Hd7EC7Ihkk6r2ueC3NjDz5pOrfQiXprpBZzQAFzIoi+urrpo
FtxsPKk+vXcGjtgzTr7S7kxAD2aMIaNX3FI/v9llGhgAh93Vn0houQajZpsW
13rDlVvZX01pJpZV2OgOdvSqbbbiREsoAc9XMN8OhjkeT2TBSDuFogml1LYS
TDi5Fq9FJ0GUPFrcNFg21e1h8PXhgmnPyZSffr3ty0EAFgtjJXSeFXrb2wt2
8HH8LJrVSDkYzP+VwI2XRwg01M6FDS0XUyjgZ6xMXqJiI6uiDK1RsHS3fMSO
pQc5HRPujivnTY2cMeoQrebnrin8WZOBvGVjYbK1N7erGY6PlHIRIRD86GvM
wWpEh2gX2A/WaAc3+uNxHI8jy5hCkgUEyFxTcckRTa79XhoG7VUFLQW2yn5B
ltOzyT3RabvqK53fxSbM5iykFFO2O2vg9HmxhH5oG+kbjRk87x8vMBvGnVhw
vSG5sRX15ZzxVeYS3oOKhNp0csY7GsdOV0qhgJ1dE+5rOav6NehxFnbRw/Wm
8gk6rCgXTKUPG3c8gArYlop6Ef1nuce+Kr+GxOo4ZPHO6WBbm+qz8HnUSch8
qVyDsmfb/WdiHieMMf6ktT0UHbJ7Yxeu8WMDTxW1h3GT62FlVUmVPeeJaDLL
+IRAXnUCreu+rXg6yBnEYTCUmcNwO3TsaFYhQJyWDrPxFVrubuiJlUw/me+L
vjrZ2+pU1PhASqaG9y2RmCTFioTorWaDir0aWxOp3rOYnNUEW6d7YNjFjMDZ
rNFDNSJSlvcwX0WFbHyAMKpiKZNdyCUBRs5RFPMspzckpe+kRwLkWfK9oOdA
wa3jkCopoJWEwA0/8xMFcEQ330OpcCw44m2OODVqWckDFaFehslqKtOOxyWN
le/T50qMFYbssj0kavnr9WCDKs33pGYQT3UCcYmO9IamcVnhNiNg6hTGNFze
8SrZjiWzhRCoWbeh7uSBiDCSoOmjr0izDliGWqSBT7ny53bW+6ne4wWZXSqU
vFGRmXZJo/10ITHBxb42f76Z/TFJ4PGUuNPEZA+T3unPk/QoYpidLqkn18JP
BhQestQ5eP0pFhfbueHNLRzKJnWGy0PsgqhXDbI0MxhAHNOrIISfz8VVg4On
1EP12eaGC2HIqRHeJaC0iySuRgNab6LBftxLuXpifmU3TNE5hxHrdtb2fNVt
4RQmDL2sVAl+NHBDOFtfjoJ7SZJIt6L0Fb+k+//3ph/7Ueedfh+CcGe9+AZY
2JsUpUI93DBMjw38IG4Wf9Y/9nvi9hzd7PYqxam3l1h91ZnYQCJL+E53sU8C
V+ZSpVmkY+qQISTK9PExKVI2IU31hK/ZL9DAgvXhNVzOKNttAG19nVxI6jUT
SCU9JGCBK13TmHmOLpOPnwZzO/izDEJrOZFmCw7+l+kwVE/rHMorVMOj1ZKH
IFKcVJcex5JW2dhRMnIFhIQywYwUe25hLXLz+6eNw1DXp+3zREgtodR1jj4U
MCaN8lMvt7xhVk7FzBuwQeDSOTPjOGuDbjTAv2g8uSsd/JegfY0y7YRbLFmh
X7EqPZn4xs7E9YITNy/II84M+ufu9U8Wyumr3Jlr9faGtH+QcTEUIvXUc3tx
ba5uRhg76bOcF9S0Fyg+jZm4d5UZeuLIJKJN5qQJxDevdfGL6GLHolaynJQG
COAf/ZoZWX1qWUSSNL5DAUNZIFw9ueIuzEHleSbqgrL0BKoVQmTYt2FHT6rm
hmaap4KlmSUvjidxOcK15kTVSKxU+w8iRK5A1Vc92R7JEJo004q1KfaGeEuL
MoJnHr3E6EKusw7QzAlA31dDjtJL1/LDMpfg+Zonsk7pxmx59NhALrH7L8JI
pq0c0I7TGxxOtcNl+kf9ZY46gcoMjY8PcglGkvfhzGDzmoKFfgHSNOdBGibO
/KYjLlseh8xoytg3a4lhrwDIU+gKKvfqIdD+mPwrLZmSXcaqTpJmzczE35Oz
5qdaFl1yrLnxq46KVfMmN/eoUcdnt4YQiL9F+zmwTXfXd64faH4m9gX0qkQV
Kz5sMDhrVJtcoTkzKL9cqzrUXWpmzaEsl+XW1oaYhUz1U+uMco81BtawgFI3
pH0jzawjAMSlU5j0yHTxMZc+QC7dV4hyS7fp6GuSIf0ee3F+MDduuATeeSfj
O1VvYBTmbRCGg3xDtIu84zTUH+GzYOJW2w00l+ootqjmrz4KOSOBnuljUKPQ
O5st8wJZUPQeu7WS5euyNID1npCv6d8hO9hv6mmBBeRY+S1tA0N1tMPZ+saU
lomkAO1q57h15UgUkN0n76mSEUTlVBPCRUS/fI3snf9bFD5drFqyN07vwqSB
HaeeJ2KG8wDELsP85hWaPH2P/NX3bJxTbsQoRT0B8F8TFEQ7ILdfCQqeIIl5
NeZ+fXCNDZX4TjVgtth/HeHqI6F/0CRQNteh+G6LYMLmuIvIOyodwJGT8Lem
ALC/J3IRuQeVSu7GO1iCfQMgdNp00TuDCBf1SEfMj9D8thL3KTyYYFJ69n6c
cl39/q7XE+hwo1966XUWTNprC7tJRl+k4IPG6ZpbHfSHDPnGQ9/4ZlbpKpvU
N8PrVYIa3iRPhAZtGbVdTNnxoT7HwEFXjbXM2sgDmS+fAzcf24MeiURrUszP
lx+ijekUi78vlyJHI4+pmBxG/eKEwuZOTgFVqUJe37RwTuBk/JQYTmFN1NJf
38ow4CqhoolNAeIln8qvgdmq0kJ76iFcpGn/gS21m8SGIAAzWl87IHsiztr8
8FUptPZfQQEwghZbHhCcHBHGwh9G+EsoLUsvOJ4topigMDaEWuos7grtdeKI
oQZ/gN+OlNqdGY0o0timSd5TgKaxzwQKlzwBypjiaCFa5jMW5bu8KielxHiS
g2uu9Y4K0NuZJ+TIaJjgfKFPg/q1bZ2I9xUa4pFZwVEx0FSpIZMYo1kQFacR
E7zpOavS41Kw7lKY98ARdXWQtKMG47mR18uTb4Cx4NSPv9hnZV2ozN4LwvwO
R9BwdG+5ixqBmdNwYgGOfc47rMbdHIVqVPZ2sSqziBSpSAW5jrhUsiABW9Ih
gEBrHrqAH52IrtgRm/i4KuijD1VROBtUql0yYtUMlju/IalPtukjKUd9a5MM
d9QciMQnUDQoRz+BG+u2x+DIpVJcJFcuEM7+GypYQ+D/Bbyo9g0eN2hHY50B
H0Qh9q/V62JqEcCT98P8b2dHaWD7gRxa/Y24ClNnsebETvhO9B+LXE4d8Rs9
RAFnuPwURX0L8GiqMpi42yzBdl36j58N1iCQraoiH4yWIKe1QbnFIwfrvIJL
xB9G1tEGI6oNilP9t1sbiemfPOHetJYngUoYuRK3jedqz5/i2LzXcpTt2MVG
fnHFOoJVfDFm8ybeJZgfg3NtfmECQq4iSJzD+/q19xOQYd4nt7gcsEqZ8auG
EIUSBwrd9bkfrPVPIO2yGeSPiP8xBBchd4FiJQBRioyj/rTGD9eMMO00vNvx
9m79zDEScbXMSqkO+x1g2vFCW6xf6JlYPcDMLpdCDOd/AUOGYmMBbqIv59ou
bEPDUjAznWQOu1hpeFr9JkxnUFrUF8W+dfhysD58qm07PshA3JO3m1m7bWZw
LJmCVrGR3Pi4gwdBK4Ru0F3zmqmLb1aUQszKT4l52ESMRXmB9LqAJmznXPcL
HfOgtvQvhADLZTHoX7nZUzj32yzLRYlfWidFX0NrfcQynE/LbNnkn3WS96AJ
Zlg6sSu8d6EZxsx3OvBdwiluftg8PdJxuEkm4sJPXoBcCpwJyz59AtxAuDND
9OLgZWBCk5Kk88FNjtbMlh1TS0J5XdjDRQ+sCD+Tj1vtXiPcbojZs/Auvf0E
72/9TWldFEW4tlrnF0AcR/Hwx/mRDBjp9ix9Ez5qCxqkS3ilKeGNJhTxO0W8
7Q4h8crTslnHaDVDmZJy0nmNEaKgHImWtW7WGOquAbBDCs0NKk+efnjecMaH
d6GGWp736PDq8hyIpFSJTTeu33L2gCvV09hs1ebhfrWh6SFIds6xvGmGDNfB
xPtino1tIaH2SAyLXYQceNjwMwgK9jMLlVdjXhnVM4eEdxN48VviK6y0XC3f
5UvV351wYYJJ98IMXTw66N/04iCi47Norwa65LRzdbJ5maOTYLRFcy+5eY/8
OVrlTrlV+WiPUJybKIvtKgkBSawYNepvBrcih3Mi3mSlJ/y+RUMNuS4cxZn6
J5+M0xFugKASnmchI60ZC19hUJaywH+9QP9+ip6GjtFv/9LE49os9xmA5EJE
f0Eb+3Fpav/H77UUUgp0VmgPtgKP833/wzKhCjLcpPee/0mSbiNOKJ+qwAny
MXP4z8lx06lQjBDDp0D3cJA7ehAajmKzwOpl1mI18vNaw2trbUMalyhXDds8
qfITjhzXYCG7T3xHu9rtnyNjqkxyej7BHYAPYxfDRzoajXPxmdR3ZE9ozIzM
5M7J42tmqXrs2heUOTt9jleHRGVnV8ACWSB22pCoB5iRYpLs3QM37vqQ9n6d
yrmFEjiObmODXrHrWe8PewurvmzeCIja6eatlczZw/jGBrFU+FMh0FHGqBLI
DnWMbBz0WHdurlB+ExWJCd6r6Z5vXb+Fdtl3VL/OSl+ibNF/cxHA4pILv6eN
HPtVGEsqVM7CIgbaFQTQcGnST6bcodyLDYnopNhm6Wq+p7c1uhEeZMkjVlvH
W49E7JAS9JmdZO+S85w74y4RMgBn4TcBN93zmo3GBJLJGR/ZUo9s0uKeDHd9
SW4GHbivwgpeLrpoFr3d1bN3senAPNxJhpbJDcpAR0g0ZD8IYzurBVDqfEdd
WbvVZscuA8G9aDD43PKkxl6zTFokpJop9uRtTTIMEDmnm+K72VCIj2KBgb2V
DnLv7DZJe5GRN2v/fQNwBqudUKHlU7fvfEERlKSKLg/R7atrn87nVam7INRa
bH0h/jYu1EbZXQXIWfI9m3VYwIU/aU7xMrpFBtsORvviyPejEBfg0Cvy6Izy
eUslFz9W8E/riwJ6302RCWs/i7fWN5d9Qe6HEGad0KfCjksTkKQV3NnGmU1f
TaKWic8cW9eJe65P2e64F/vCbZn38QZLjchSn5F86gKYfPIURkpI78bYUhI2
HrXvrPKx8aHkLnEmMylZUpA1yw0azHCfdtm89IkXxSDC3D6u91h9zwmZiuH6
Sq18Qfp2zKb+x3UawG6pMaxAleH474BA4ZdsbWu1p6rS0zCxEyouajA3xkGA
eUWWp1QKns3w+wv7SlUyS7vWvz8Cy9fxTLVdLaJxI3tlJhpKwED8U1lfUfR+
1Gc/DP6rq530oi4djX4VeYCZpVxb+8MWvJiTI1Y48VboaUpzvQ1dskmJu0/6
IiTBtJR7jPPJos+xiQkfLxFdk4tj3YcpKI5+zEqufjYys8W7OG32Sc6EkpEf
sMvojzP8DHK4vIa+PD0kymjfj6wyHS6WkqZZ15YhET9SE9+dgR0RVflb+kDO
WufSkp0FIQiTgsCHAQIL8Jf1WqVqji99W1mOTLnLrVvSNC034Q7J48TWUCFc
OaFOlp4XEANhTML4IYhuRUvz5THzp43rwFmWNhaydlzPwYIWcr8cxv+0rupp
YXWn7MiD59NQ4gB/mvHCC89E7wyDk8mhzyw5gx4k7oixXqARR8PiOiNu9noH
zEfwEdQ53cmTfqAnKZhY3oaVoRZwoz7AIpjlqux2u/oj72i377fx68HNuO5G
UybHEDinp8V/J7tRPN1bC1FuKmfYSQ6190QITbo7hwXZjf9N7idcY83YIq6Y
8JtSGIODlgXyrmqAUFBqUKLkAHqxteIKVbkoVN4ulcmelye/BhCaUs67isn3
QlPBfaF9elLq6LGYcgKH1F/X+iQx6sRvHKDuJ1pz1VvhqRhG/o72jvlq+QHu
3VBm5Mz2qw/ZfAfUArEQfQwLXHzmTLlsHt0+X5V37dgZ6zHGV7eYZd+KfE9m
3EF9JL8w2MSyCDoaLE68BfLyUwSHNq3GVOXQcq25fdAkzkwLyETN7cnVk96w
HQoBuFU8jpTbTbzrsAGC6kt3L5n6JvvI/CdSkTpy+juuNTXeHQULDLsWHtfA
W7ViP7+NNsFWNHhn2OHnkKz8S3AFTTMXJb25QBOWf4qjwdsvdtqU5PZE8sXC
wfam4v9Bulhya0HWvPgXaksqAqZ9ScozsfyMDFtqMbV8pz5STAqdI5dZAeNw
Og4vzRefArMrRVR74QlRkyWrqmwpmCP4xxJcDsjx/Iv/ktDLC3iIwJdYVbDd
tqdntt5pVqC9JUVMw4i/rKlEE79o+fW0W4HHaUgfmPwcda/c6sy+P/Ux4YxW
qvD/J6fOIKCqpNbKBBAtTJOgqeqHTDdQoGZqE2DKcq5xxrfpXNqPGosgT5es
ymCR3I/Mb55THXbl8D2+cMu3bBP/qT6A88r09sw89+VK+15dmE7ekX/RHbQU
tC2GK/v9jxmQIriKCpGXZHi99zvatMcyTPm79Pl184m2YM3A/aXTXJN1HX/w
vn/n4AseJPiQmy1oJJk3UItV3v52NFSaUdDBq54D/ioc7rec+O6j4j2ecE+k
toIsXXKvda2yzBjRA+aaR2ZKpbTtqyitqWIjZTSRyAf5P7HfRlg+E2qVtlvK
sLYt5BcVvowhwqPOTUigI3EY6Lb/lFJQ7W0yywSZ3EOk2ZMs+CM+te2ltN6Z
kNyILbqrakRh/C8fWxkRQYXlT62Tq0z9yyLHTn3SSeWcBVYo0g7plBuYn2By
tu+2tliKUCK/tpv198bHz3otOuE9M0c7Nm4QJotgNWAnk3qxxlCOeQQoRZZn
84qwig+4DQR7K8vnvRLf9BlQSuWe8t9hFU5bY/GM2LUklQYgxfvEo4r5h3h1
JePzsRByzTUAvuBchLabr6vuccqV/zbZePdxgm8E3/n55E70YegYwT3hMNnj
lys43cI+d7x4KE1/NvGPpe+U+s/EsTv5BGkGxmy9GHV7tO9GafDuUZKp6Ifw
1Yj2NyHlhLwBdQEpwEMnBBdGUQ5NL8KBUJqhd3xLpRLXrdfE3feRrYag2rnB
0ENhwQuy/N8BlhVsYwzSZAybq3hycVbK4z9f8LhQ4YYCFUmCGNoUpJAJ9tVe
EdoeArSemHKMybQNHDUGyOuk6DszfeDVffc/9HgF3sBfg2rtAN396G7928n2
nt7nJZ0JK1lLaopEfhuAvWnm2uFJeE8zzAu98JOrPguXcFFML44JrQFeOajd
UgJ7bjvo/F5ZkcRqJqh+lzIhqcnQkH/VOYZCrpYJJNcdU9Fxb08CjfT0o1Rv
tHR39/TWdrxx11clJlCo97E7r3+cInjlZztz4avj4zKOLD7skUzEUMfsWQki
MU6if0fSFQYGOAURq+HeeVp9SrFeDwBXBc27msmUXK6DFEpDm54uDMK21U3g
+XLmNsFlNRgkYC7lve9cb4gzlt+x73abfPmojtN0fdHNjnAEnVUmixIEcNhx
bOj265jxgiMX/3H9plFTDFNo6PAAgW9NIyi6s5BEW0scbpwSyvJ3ekIwxqdC
cwpjCqiWki/pUqCEu3+xOQgI2WOEvCBvRP1adNoUQ0XLdPKHMGm75Ou5L5ee
uATyBAZC0/lPBayctbcmVgAYkA4gW+te9j5g7EyJau/Yw6h28W/d79cbaTZF
ukRqa/P4aW14m33siXwciYBIcStDFCqR9uhK1p2vFLuhKYI+E49V2dX+vwSl
UPWNXXvS0wrAe4mbkDpVBKvMFc6E17W/NdiOuuS8mmO/CeM6iQBNSHIa59Zx
VCVpAFsDofZm+RFSwcuOPSLU0U/bgUuiOtq8jW7lm9LdjdgHk/VQrIRb/S1f
HEpaBbMlvKFs3JDVPdExemWEnB+QwnoLz/bMZSMjXdcsn5hHnFMSYQSjiwfp
4RLItRiENWVE5KLHAAZePeNljS0osoK+ihGS4m/gggCCBzjb1BJJ+a8AWhDB
O3fXihAKwrEa56Nz5z8vjuwYJkGJMhi47Tr4jWEfD2ryL/V9geG79XIYvqR1
DLENxEcJ1dD0z6Od0dLUDJZswIlBAdRFhSU3IxYMNl+uNt1Z++hiBZkJYYSi
zEEj+6NCvaawJy7p5AaqN+qfItlLtEjILB8rx9JE8chkc+m3qlVJPAy/BRop
rFSDssadoT/jNTYdNot8lMmy3gP2jcdbdHR+UaRNE3Cn2kmJNVRBe8HZl63Y
kTtyebxSuT9+hREaFdUhUcNMObRZJllEMG1HuVhqJ272LNP55uacgni8HMGa
og7TBRYZBBbH3cbdrwEE7u6kBTzPVuZ1eujDALpmoGBm+wJJ5AwHzFNO1aZj
5XYIIFJ0BdW2DVPBJDpaGM9wH6CFitWfxT0q16+rs7VbHeRjfJO5JUIbfR/T
Y47jbXdaSPStwhPVfwqNFO+pjPXwcgVgwgsUXc2zfXj1WW0NGwkBL9XaZznK
ljSXaO7aUYG86RvKRNM0QmizTnjOKFJKuRNzkESP4jLwVPLhNr7426BpjEtU
oAy5IQXWeW+loTqm7L50LXqr72JtLA8m/9wtHS1ZjZ9oScyzlk/bc31g6f7t
0zq+7q+BDw6S0pxfPgUBO9r/xYXEb/qB2TXCgdvIUYT43RquyQ97pXErIT9j
K04BzoJNOitBLZl55W7GgV2BJ+2eKDCJRn8mdb/XK/7AeRFQLwIGeuZA5GOZ
cZvrwyP8538ntqkJ3iq1xv2P2QMeOTyuvvfOiN2MIMUVFgfYuYbjAyCWRzDg
LbDMNIP/iLRPkuS7oXiJXQdDh1/Ulc0TWSs8oefPNNoGomOkVZ/SjXAcDBmB
8vaWlGtPGQd4jwGMtqi3xRhF37Jrr7srSxcPrfNn8K7cPcz9PEV0GQe6kUc5
SuqnjnLXd0IIZiJV440mpQ45zN/2EPd+NVOG89M2Hu9wqN2tUWj94PFssinV
vYbqrWpycfxENcskuYO9NmN3YJYymdnu15YqjXbnlLOGJIsoo+8TSsmTS3Jh
HknL1VQPTE5BMocX32f6EcFSGTxKbeQbSeAAftgZzDL7CoeVit4i8CEHWwc5
XZ8s9pvMqXiV+RL8iAN+7B/vOSYuY41UdHojdTmfk1ktSq93Fg8yBnHRGnyw
YCKRJSaH1a43a8N3t8FUwg0ILdooz2C3fc742gUyw8VBH52WZNV+g9G5+pST
V1PoSTlPTw7UevA4MccX73S/AFmVXS60gkcMhjg384UYFtJbCwHeKOJyQGWb
6koj5rcBt4veKUzTgNirfxBI54oW68sINrkhGfD5YZdP+Zg3hCqjNP4Hjh1L
Byamc4ghySZFJ8fFy0VtNcYfaaLyStpX2KWoPS8kA6lmltnRRE+85hmKsB7l
VisJshZXH2GUuamtXBPHrlY9O3+Sm2kl9+RTUo8bCu6/qltvi8AiETMAumuH
kWfcbGlCldz7zh+dJpXsRmWsiDMXl0BSFaSggkklRYvDv2VLPlttbsywYYqu
rRZCwqJAYTC+pVbR/Db3x3cxcXK1nJtTmX4NhEEAoUrYdGxguuySNOBn37sw
PT8rW2Pjcqbr7wCUA7rfImch6Cv2nZfMDWEIQJ4lOuBTfGNiHi/SaLQ6ecJD
Wxy17/iAv5d0/ugDUsXV7qiEi6xK1YnsgBP6DkT/CrMg37AIgZfgZKKyjnF7
ukWFA84JFi+RuJl4uLLfvDBt7oLig+79hBIAbcJKj8sA8dhz7+6oXlxyDInT
QXodV38r1npl3zx/a+8y7/bhuWsaI6EA/297P80zDVw+4aJv2RtEzvDl1NYy
QSFOfYnhZ26sKNG6qK39MyEzsRRTmGSsjqPME+lKGah92oogOwVULJVwTF37
Jn0VCe6J07Nrd6Y+ZjmYIo78G7z43HV+Jwju9Fxz042tKbKLFlZrDqK9PmAe
ZVH+wLIilghBhktAkF9b1SUtUAsyGpqvy3fsk2MeSi1yQgkFtOH2293t8cei
ZLNvk6SW5JRqoDoRFcXgqajdVKaT+R5ZaPtDPJyRz7ruLJQj0MQPSnmrKOwL
7QqvNkPYW/J7kXU0Zs4pJ1F5utdjVHlD5Myqb1m0M14y0uFZmMo7+yF4XswE
jmRoAjz1glGYz/RVgZ2pCqJL2iUb/syJzhchl5SEld5OAuvAmmf1ifTBZ6m2
fo7ZLSTntmHslM2D1oW1G3IW6YWQeu+fmzP6Cd2W6YhcWJY+HomNjYE9rORY
VipALUpZzoZMQd3m7h2TgzRJJBP2Dk+PcLbpcKVfTaIqT2kFvonhWsjeOyEu
V/HdEcLgpVBbzU/6knSnftDmn2idy5yTw96kicDhe6zVu84P+FFhD7onYjFO
7QXI16QsJyG5bgyP20/DXjOn4zipHx0sQl5VecQU6U4EPJhgK2sG5TMGl54s
4K3M/3Uq0VDqv2vAI4KaTb6XALxTQ9FHwjOZ+VhHqXbInsttndKK857dVHH3
fwdM43noXPfG1u6FLeO9GZpk39be9OExPPrM6m1EmAKWmTgjefCVOHKM47d+
FxFiuNK6/TbXrDRi8Ul/8EZXD+0eL9NRhvVXu5ObMG9aH+ABCeaRWRGXT4Ns
dMdOfsc5rRqFFfY6B54hEpnVvES+TaS5xnI2hF+akOnyN9SbLOeVWuhCpNWp
XoIMRILF5UFW9keNayd+EHL1Bbkwwcqqhm6N6GhKvDFULL7lRZrruEjwL8yA
o8mV3vdIAuzysCuO4EV6OilvG73RwmO5TWAe9GPYXXTssWbNSVaUajLFKRCy
vsYr7G081Wz4D2uyqybv0FodyrrR4gjFD5kTXWFL0jXOU7QkJHFW3/4vxvev
sHpx0ouA1CEKSD7ZPSsx89rafv5GsHUoPY5+WYiV5csIweoYGy/YwE/puO+G
jN0z3ra6q9h55HZv68Y8dXrZLsJE3cxiCA7wTi3FpMcwLD8akGCfPZxIJ9nJ
vEmLQfB7hLP22n6xcNR/26Ghhk/+Bzk0V+cXheKZDjN9+rzcDUrCHNC4TjEh
nEZGcrL9lMyJHjx8EBMyj4kveDNWCSuBec1IivzxgGBMdujUE+RGoC1FFezR
//9IAgI6I0Fw3i6Eo81IHf1SGXWTXBWhCzRXvRI4WKBCtnkDKgap0GTSSZYJ
5mJR4aXmw+41nfl4LzN65IYfrncLf7N6N5ujeUXTRCxuUj19gI3J2nKXa2LF
/LoroyLhZ0HsZCbnOUhsEPCHw/N1WMT8IS5uf18jlPSTfffEbog8zapqfT2g
26FQg8+XYUIbMbtS9EyFiWHbfzIDK9APk2/BPS4RVXAsXcSpx85vHma/Hzcj
MK0IcJEcj70zaaHUs6MNbqKuFTLDaZWvcHHxFVdp/fqy5gDdUEqWMy4H7MOv
Y/k5DoMMJCenNSmJ4pE4E7y/Cu8ce81L+AnVY1TIKh9v0qmk/7bTy6LpZdG+
LwEcpqrfr1VTS+0glvm01wAtPl50689IuKDVe9G0lO//e5BRW4D0k3C8BcNt
n5Wb9Gbum4r5yJdCM1EvIF7P68iy2NUPowgU+Qosy9zhBf3Rbhnx/1fQajE8
L5h2g/Kj/lKbRu4xg9HE/0bpl1fvQ8mOZIPRbUcTh34yfOy1kDhRXdVMR7tS
UoSODrTVlERcKisveCP3u08MIbonU3kcWOEQSMkED5fyTdGwAi1MWqSnbBBE
28nnGMh+p5NrRuQVx/9MbeDhhoaQPcPmj05Zn88HovIUxOhmV5i9DDfPNHXJ
DxvQ/Bp4x//dhZ7Szmrp+eqhmimne99LFaJ9RbxGjqp08E3iFZjZbl4P40uf
gmgqGd5HTgxutFvBp5CVGOll1SEmJy3dcT++LOZKb8Echbb5qo6RHmKnpyls
HjRWcs2Wxczisa+Hcor1cd6hu2N9Wedcu9HgpE57EaUFOE4WY72vo3a+2nSk
YIpK5KlgccR0c4JBLl+xSkDGVWoX0MK5eItFoo2/N2+D7T1NRlQ/XDtlYJYe
2l1gw2whBgq3yhgAeJKsIyseDMqGt11D1tpt5Q+i/yqcKwvibsURdA195Zly
lz0vgiPTMaQwbKKJCPQrQPiFdBfmmMvz4ldy5SddX5TIehC6LLmMxoN4A9WU
FkV0aRfJDrRs7Wbruo9WLqIc7wLz+euTV1fXOTo/+sqFeQY48o1kYpTVheTg
TWF9Fl0+lMAJex3Mbe8nZsyXTCUQ+/1gE5BRQV7+YB5/5SXZoIwulo1yqViI
FPyOEb5BuyAuUwFWlPx2I2rxUDm24Dt1Tj0sBJWPby8mOOR9TsVW/d9FfRQj
S5vSSQWmiKyBWHJugL6XT5IeAsZbwKNMDsOys3pse7biyweAUDiCpnhNg0pA
4bi46XaWpDSPkX2iU7RSzV/HZ7gA4SLFIdaYEtmtrArnGJPQ2pt3fvt/Ce4Q
efH8qKZSznF5jgp1uFN+qFh7EMuoaXTnkDABD5+c1W94Rsqhq7rKOFg/1dMa
pMONFV9o/COu4764qIi8pgo7VTshmezO8uoqVRyc4u9TdeTueAOPPuP8hBPH
Z2uPu31pqr8FbhYK7LlkHoMjuVPJZ6ikb0ipTueHaeSCvso4lXNpduLoGvbH
NsKIPcCXucnluCwijg7YBcjGUViev7plKsh+qV18xbfTOaYV/qZ0gVdd/jFT
e6VjmMqKiP60lLRhfFc/TjxrHtQL1j8SCRI2zaOhjY23ZZwLSUnIzAHJe8JB
Q2mBE120BR64hdGcPTv8NaRIE4X/vgspo5hJjn3aSlnAUlBK75ey3pdn/u+b
Yx8BI8j9qbhm9+8gc+7E9NxUZNtgyLJs1gVmKhZvAEUgtAdQUqsuA3oRXu88
XSUQR+rEMMt3tKpY/zNCjvgIKw+QWmLU95Ml5G8oWEy+McYjqmRLZG37pfC8
Hx3cjmGf6+i06Yjp6GKbFRT1yvDQo3UFxU0j/VlY1ndPbt8uLvH0RCQqdxI8
HIhNrPFyBsP0ALUG9aJCmyb2Aow1OC3nDWyKfpkYr7aRYrx1h/5TjYCEL+Zl
PkRANo6NYbn+c8CbW5SZNtWvzkrkw0OxfZpWgVvbzG9Y16w9ZLYU9zb3ddqh
DbkOfqjtzXTS8OtKcSp/uJmJNVJg3AIv9qBILkZd2qM6nHDWAJdGWtaEcmx8
Pwj5Ikzimn6QCadVF9//z47pWaZgwShRowRZtqW+hXkcqXkndqJafcWg16bu
zn2UDjkIie10VgUIIYXZ+vPLfJkURl7W2ljFQJ96ZJbryyJ/if/m0PsjLl5g
MLDMSBcAANWF6gAkYE4QwlvUTALSh5O4H1GyDh5j0wKicONAh5GrlzeW4MCw
AoqkqzgFhOi7ooCi3xeMFQiIHPuDAirBE6Y0cGfTWti786hnuaDeo/4aP+3S
V9ifaw/ELttjRHxlUsULUFWyjJlYFG5QUyndZAb7s0jQdBI0z/II/K1ek/Jb
Wvm2VA/M2d3umsIHER/qlFlyFpOq9vX1wc3nBYgvjq6W10dq7RCusp9APUl2
LYWL0uMgOpkRj6e24wwjuOp97EDARFkFUoTTfDL4iYJqx2yCQArbUalb6Ctf
V8/5+AA2JnSkT9TcQfpcHFQKrvBj5av/rmcdQbwiq1vu3cT5tFIvwmm4aCXI
t6XywcTJ+ZyhUm3Hi9NzkuoocCpp5XxigftGSPqxZ7n253aty4ZDyl06Gfip
Lrs7DHlkDkzpdUddx5PIa92BJeZNE/skz5oadqH819MV2/bKnwJ/VOjzY10H
lHeM4fbSEubhakCYjQ64g6UmWVHJn5jkcY6lo0Dw6BMOTeo8DkVvF3rjyQ1z
tIvV5dKuNHJCZ1ZvDG8uX9YHfHx5DV3qG8iUq1hqPYUCXC0S7ltnsF5xsF8T
Gotg8oVGkSN1jQzE+8adl1cBjoE+99YQ2CM11vWxdMfsXN2SEgu/dxNGZLZa
ylSbqhFFxNm6jK9hFzBeb5sLopXYN3RdSV3HRiGa7xnoApXnKSx+5eQeTdhG
MPqVgQBnbpTWLSSz8dbrhA7QdJPwOVr3jcS9OdsFWv6nWJ9t30N2eD7vjHPM
oaLoevI7k2w22zf3vHT4I6xfbOjcmKYpamANgorQr3hs7/U/kMFnufYLaodg
NqluE2fIMmG1f075yCUXj9hC7z7qIzqrpIfsl0FiLGV1mGR6mtGTedZdAG0i
P0eS6yitsAJJh2yTtPLOz/ebQVEWvEBn+Kb9dGUrTwdR5cbBbGA7DKUVcwsZ
kO0iZ9irWeb8aw5WxkhSrB7YshuIXUb2mG/44ABLMCvyWbIzCm2HeNhKyvIz
RqSp6f1raOKHgEzgxaX62TDLj/dGusFRB9FQpG5+sXVi4215xZ/hZUjjrHOL
Q3dbb1NetVbPwoJVl+UQcpOzdUx37uDRrjI10bhpnsEWDcJ5Pnkct266ckH/
hseuryPlrenNHjHAqssSy7RSTj2V8NTRd9Ybwxm52kP1LnF94kiM5JDz7U2l
fKYRxQIiQ1UTj1hzCYS0p7jh0HrifOKmXPG7F30GnWQW1yogOLIrxSkRvc4G
w6xJgIIMNibAyMJrz+qC3OFP0bJdIg/6bqtrFNwkyyn//h1RWMKuQLUh3l3L
kApLI4lp0ieTPNpCAW5QmCqFB+dL7z3OOtFuNSUfe52YUdEGsQoy7bd+pQmO
6aqKa56LUgeAcHRBj5QPvFFIahKQA0lEKZUtLgvkNmLz4mBBR1UYNAyakFDt
BqrHdHpwF608AUHweFXelKThbhYX8tyfnWh59NegXPPB6r08JC1OrcXaBgli
2MGhSOhnH4FCqRzFdSNoqh8VYt22qbkzMzHYMXfoU3RV3FZ63s0zQAFpJKVX
o2zw2nwM+AlxDB7jexE8cCIowYA0aWq0PbVakPH2LDl8+tl+E3vBQe9ldRyg
zYSCvtyICWkFEtJi02iwXTLQ0tE1oUnVpc6MBL5d7BsEdfEw2a4dJADJFIN3
aqt+Vd+Ij2aDcUH1wHEfao8iZB2H1N3fofFflpYpfedo/Ljc+qauOO5TUTj2
KzVZOUI0+koyPxaFxoEZ+T7NsGLcM5twCiZmLZpWl45ZoR11AhXYobAnQ7oL
QYElo35N5n4ER/evNJWTJ9T+vWotd1d9uSD1A6CxNiTLWMe9l7zR3GZOZFRF
IrSGdGZu9pR/r8BiJ0/asTGbxmOj3qFzgGtOHPIz6gi4NC/xBN/IuV3NmaaT
TPvLgRtkz6br13UzN31MVE9Z+0CAHF9EcKJwsl/eNtjhT6iFeIA3LyHuJ47o
Zq/K0T2wplt5qX9gj7j7pq6CA11z2redPGPobWDucFfInx1tYJXLoGv9Rr38
BYq2Tk0+r2l0WXYuhzpuiwen4g0oAwz7rxKtxDh6avsXzpxEEpA+qt7N/Xwf
jSQUECyHd8oNMhYsbElSHahO+EsXiOHFfsErc6jXQTeKk6Tldr4gwUPc9hOS
u5mGB348awVCNMFO9Bxmd2fcoqk43rzMZOfwjcfiqv+9jX6+zgb4A+9RATFu
eyWV7mPpZWQe39iCqza+REWF7InoGzy+ZmKtvFDlrcz/vu3TIm6c2xHESb6+
2mv8ZEJJQVpsO0uO77GUdLIUtbaOQvXaNOzEvyyc9lppjmILVV7EnZQFsjo6
1h4PwoH2kzMJbDyP8j5vYejKdEr07S0L+Wu+cTEaqtXKb65atsJ6pZFeSski
EVvf/eiAgYxUnpO7JVFGWZ4V48FJRCo6AXHPegQ+yE1cwTLrE6gG8Hyp/YjO
/iNDgL+FPemhKJVWCEimAtcGgWxhWuFiTcPVu4pVZNjIzNNo5R/Ia4GoTekh
hcva5AGM/6Y1TOBOEnobq9gEyTtq6qion6G8A423NjTOqO8/N3Ccpmhe66+w
nLQgbPiFNN9El/ZRoeOM6/d+ycvH9eI6pdfFnuywq7sPV6vPf9nz5ui5fX+y
HC4XFMT7rgupCP2hAPy7A2TKCmJkFcIZgN/7RKRla2s+YJjG/BwhZ2exrsQl
GbxMSbs3mQH9Z8ZVuVPBVEaolS+P60fea1nNHV8WEUm/KygqVYp95bUTgV03
uTP+6wJ0SbX7mq0nXadQICfZwGF0uATwQDUhMDSuYb5XFCcoBSxspdLVjuTI
frB5Vxq5w/8JEti4IhiRbaAaNEhlmxmQSmsme/STI3wZAj70jYd3cSwntjon
6hy8dj60WIwehIDuu5KgZXF0nvVr3zQbjyAsG8WL7+inx4AU8tDKjb56TNbl
UClQu9xL+oF34Te7qavL6QcJhKe070uQBtwSzP5U92lBb4+GwyhIB1FsqkU7
dyJJqznJNGPmo/EDZW3aFGKVFmROUjLTyPkECgVgpwN82HJKrd9E+kMtIw3s
T4VeTTlFweCRONSn/zevX2kuLN6QD+fBMw/k0zMFoac4mVJJGiXp4JBxvuKN
n2pYolcAy6RjY/NuegfMkgQS4VgEX/oUKxuBATNO84gMId2HqQDopCUwgm6Q
/+BR3w7RiKaG6MBgG+89GvEWa++ibKcvkKb2HqTRbBz9jHPscu5ry4uU20Mv
fguR3/OLRMt2Dd24Io+pylY8WGkBIg+bt7aT8laLeeK72LvmU6nJ2P+hKLgb
ZDxd7URtC+2pDTobFcrWVWr2cnwPGT07TQ8qEWRmKHmBgOMJaIFY4QCJBhrA
AU8YnyDLeM5tMe9TFCeY6/qTiZGMoG7oqFEmWwv5sJI+s/M+lT9I7cY2zcJ1
/uT8dtalsNB+df1iPINjkHbJEegGEKRb7ObAVs/dQb7uTKVX0IxWwRoHDZTe
L9FJyIklnhazqwYv51FY+5z5+gx/zZBKoQ7TmUre5fNZWlaTmW6mMabngUzZ
zlSaGwwtaDhqDasmuJ/x8btbccIG1UwkTlnx/60KdxBUpO1OQeej7bKn4Qgq
JRPhv4Gf3YtjmlO6N91as9X6WIM3whwi7nx92CCMfkrgmvWJlkoMuJ/RfNz4
mL2sPROJbU583M7CM5kThEgAOOCBeFzZegRN4FweprsNFgpqrnbA/szyVg5F
s/3DXphmXJWfdiUEua8+bYW7J0Ay195AIA0rwDUbiRArpoBuu9TbK4qzKR2z
cWHtu6L8RvqyjRU9jFo2A9hWqDCLGVipg/VM/mTLybQ3xkJBfTaZbsRqOixn
5/DW0YL987Herc3vRhVYI2dELJelWW+b63EKNzSIEHlwLjpvScjFM+OrFmPF
BEgF8gcOEHsLwRoaq+9n4OqleQfILkiPLU8U3Rpc7+J4K3/drrI+2fd+JyKS
DTQtg6ujbUMXdrTKfGcczsCbiv9QadxxT2kywBHuyArEMoVHm07Vx/0QQCiw
Cj3LTp1sBUV7qYaj4FyMPTg/AfHYrHRNAB0wZK9iknOPTJTipnORNSAc1meD
E0BvoKcY4elQ+GJDg2EAxORyu4eweMuQ3k9kYQgw3wqGAdlSey/iV3cGyYWJ
8xGZPmjy17P+wLkWajBgL/a0L5I6HbWHUKpM8n32EPE/VmfpOZ82HtqHpUyH
pk/A+nsw5fAJKnu7P+OAVeHSkMix7w6w3pvRUXLcwnsp2sPrw11sMO7c/0TJ
k/DX6vYQ+t+JGlliGi2XDSPF4QjCA08x3i6r17SnDnLKVcM4FuhyUJ6L16M6
tqwk2A1WmRL6IvScyU5kYwAuaGzzOZ/0NvyacOlpDURuWMbXUjycaZ+AaYCA
deChYRc8CouYrl+6OEXt1QPqnLFr7MHdpNI1piL3ET871koGm9vD/1QC8mKP
npoXFeXRFjF1o/oYgfmvZRTiObmH7azvebn8WbUN+BRx1dLFxesVi/AjGKp2
Saj9PSluZMn3Ez0xtSR07bvVvV8x/mLunFXqSyPYz4VFtRWj2Q+m7Ndz6IsG
8Ex8kOx/AITJj/hwGnxPQwS6d23oDXMbllfg8vU/bh5f5UjbWwKmuPGDr7Gq
b/5ka9TV2Tcjvta+CIB4+vmqQ+7rtHZpxp0OOi1tQtpKhtzbj7LuJo4yB/aW
IwwKZteOhAvz/32ZhQ7Njpk84wfuUuMEtbjmM9UHQYUF2WiW3SOxR+M58EY2
YLs7o3uday+P7y2wcbr602nU98sLstK8c3s5hxZtjIJmjJ5r5OFLQANalBdB
xcOlSWTS9gk+HlPDFU3uITA3cY3cCZ4/1SLYc5G6AbwHgtszSDBKOb2rIXMS
LUSSfDNq1cp3ae+uFCThsPef+RntW9Dk/wZVHmGH9Q62YXYL1BmvEmcNkhGB
+rQYmtcCAWuQUSbNXiVh9/uzaCEIv/Xvh9M8Mdu4JzQ8ljsEMyaS3F8sUoP9
NDVY2hbkjxtdc951lqzgU7grPPB/P+LlgAgkS14bXQEgefVnWAUdYbOWL3P8
WgTc4X/6lgu/oQoKj6VsAdT7x+17Fx864r3ghxCFWJhXia5DyBaQsYFx7Hn1
G0juXtKJ7ottFk3rV3iSEfmcDm/544V1O0ymqkfSpXcYNlOaFhOmG0Cdcxum
oGb+ROhQ6dOPGcUArAxZtutl4jKnK1vLeS8SwZs1mAUxhySyZR9tZo3O35t4
poO0jVBbnOI4oZY+keetL0xjohm1ESo/Blx8ddhlyG4DztUeuyAiZzYt5JKC
X9rCmCz0vNYyDN4DK10igWj+y8DuzskG7lnVr4Jr0SaU7OBSQ4QArkCz1AZX
YtfFIaiuz6GlVxsb/V/kXK5R1rf78EkNWYh0hc8xW2+6aPiY7jYAgtHXOE9t
24rSORXl9omwoZ8wjFrKE04uj/nUxx2G1O7zI4Smhw1T4y4xdOKfTNZXSDa0
Rvle/iNeaUtLmLjbdFLIVWfX/WNzkJLwqINdsr7fKhzSo7oHDJcZupZOgwUn
6Vhl8b2r3Zrbgi55aC+aOjZXqNEFqAuT8iE9jIwkCVSXaCol3KkBgXkH1VW2
yOdVzHME9WaALjr+kNd6HnXMan4PjhO8xa7iThT9g7D0icJry0l1SubAf4R8
+nKT4rmF6e4BZm+Kjw+RmL5oPWk7L5kfFpZZcDbjUUl2C7xKpKrX7iHE8O9o
wS3x009fYjQvGHmJrg+C2wagl1l9aPNrzsOmgoUSsyMey54T/BDQYAMJRRbJ
K+wI1PiRSSnB10ceGYHZ4bAbmyhE93KeHF0Hhfo7TpfeOmOzBA/USy3ZA0f2
V05wtbAIfLem7U5PF0lHJNqbpGFs07Wqs+Zw03HlqoPWY8e8rRSQhCjW3X8R
SvEauLgVSj246K2KUrNB/Saam5jPTlVQQI2HJppU7ATinZhOnuFY7ncqHYEG
M+a76JyxAks3FSBGHMi4ZHguep5XzIpz4Uswx31UPI4AMi+wjZLo1TXPSxig
Vy4SSN4j0aPhzqzRrJedgm8p45efIU5eeysf5oinYQUavyJPa0fHESp0b8mR
hBGjaRUJEFBCXKr6XLc6PWmwIYtEFhtBhADjD71tHfKwxWgOw07TFU6K50zZ
y/ObwNUW24iLFJDpQvGobZ6fj7VfSxdKW9wDYwdSTvGw9BMpPmreJizdaBOm
+zwBRDX7keKY5U+i5FOQMDpNlOtNKSeP79tOJqMjWS8J7YbpFVXDpZLUTA02
WqnCOKo1GwYTh4YWLDqsFj6yL+j+PIWs/KJ/4SgBQj5nUqIDkhBmwJ+W5oX2
xxkGMe8Tehx96pLqfCIAFbidVbd9wip3nwhiNrehYKaozl5rKTPHu8HZEtX5
b5jYGcJq26206BDfOtRmWFfKMmtwqBm542FZ106HtQypPwvW+Cue8tgrWuJM
75RehqAsLaDym9BBsFbKqOqOcfGHFcF5TIzgNlFJbzPN0Dv0Y7fuI/K50eua
qaorFgJuMaMJLf5PIN6rMIYagTKV+p8iQHDpf2lPOTlGuSiVuivXR/aOSMwz
NUx67/wFXtLdPySTgJWTJek0tb5F6AaI3sB2WkxRj7rGwn2PQsQ6OQQT2qzD
FizxLb4y0vbXN0kQZELp8hISsmPg5ZCo/Qzwsft/37rppUEf8KvpWGWxPvRN
CxDn/5SkKf10nZFhW1xaA/nbyKiLn+OI48YXNK28A/i9AdzqNfoH0yvf0UQM
ndIXCqzbTdALJpg84yTJPBZmOQL1fjXWdo6OhQPgn0VrClV+b89n4KgxxDeq
ybwaVrvU/jfflm1BqWOdqLwXcw2zVqI4wEazRbMJ0S0SJpSpKmR7seSERiqw
pEmN7upVXuwG0kmpLnEpJQvkGFjTF0g9qNgjSbHsIGC6UvPuItUn9qRi0StP
G+ehEWdXzKarBpP7ZI0bOyOLqaknU3v5V1Cg/In1PSkgU8NPgA5GIP2FdsSR
q9zCRkdYmCeMWm9YCQT5cia3HZNfD4o1/LzJCvwhXV0cYAfib1lkUFmFW43l
nGsaAYiLnF2Ak9c14svjdN0tJx08vKBH0Q967qgQ9C05vROcKaSVEE4tpMrM
R858HtEPKu2H9RGENUK4jXyNf4j/B/JBxaJROglsbh2jdtBXj4ka0+mEI81u
oY9J9SEqygEdV5ETtcvk7qtv0zVUtU8pbwTYO1mXIKaGbwaLvJYOgthhjDrP
saP8eL9IQqwTQSjz227LqrHSKSZy3zg4ZjeuZ4E1kCkc6OE+gyb++lH4R5Ys
OhECRZyvZ6EP7B31WjCUyQoXBv/viCi99JZJPmSObWJyvZB49Yvug84/bFMa
kU/yrleZxMJtdQjd+ovM4azsZZLz7nmUMmv+Ah+1NgJtc4YMSJeqLGNbURrW
0aOjyhoeXCQza2zaTCbM3rvb/YCx00QW4cxT2kBrTy4UuS1ei0j4uY/nAU8h
jJFxo9ZpCgwViTIezjehWpmPG/yzq1J7x4Ce3KOxV7JqZyt9/xV9hO70VXrL
UtsPz7C7UYpHRlVuPbQiZzISRdh93ElwN8JJrkCV++xazx0mbd+UfOsSwj79
bNagd77PdEnJHXO5hQdBAevrWN9KCqcYEOqo2laIe8xTz2vMc//q3v5GLl65
NTGJpsiNUV19yFB1csiIXcJwyischqISshgBty7rTqhQzl6xWvOQOrtEws+I
g8uuzyD+dl3+DIh4zGUmb8SR5zsba9WF18Jd43mhGYAK+niMkpXTee7WYCVl
ap3vUiYQyso63/b1w4o4pmbmf+DeGgoaiXpVE4PgpYKfczbQh+hQsPMpoNkd
xAvpL3uMPC3eiGd+9Q5+AOQOr2i40yGyLrMQZmjvGsZgTbvt2i44N+r4L+8c
wIvF9Mc2zjir0cONTmos3ePEFB5JengbfPEccmz/ZhlnqZ2Bh2IpeHnGG449
rYuUaNMiMP2kNRrHc/ADMUqfjuD8Jivobc4Dvg5QtFkE5v8EE+p4tc/URAoM
qqfKn0B9+9Vb7ZGXqqLQWFIv+zOimgmX8y3T1PqAfek+seo6wjQmm+VhYrZd
KvpXXjugVtjMGsGRnwsELG/h3FCOpzamfR0CrKEeCYKvHu7th9tujJIRH3+t
CPpZCL0v1LaPKhKIh8i4NQDhj7QiDqN8TK3Esjo8WRpZPcSDiLhtySwWIfB/
qSa4+trYjMkG+Q2oxJVsYejmHfO8RpUdBHS5jpdJ0mmzJub1Fdcxv2V8xEwC
nAT8+yssbFyXBgExbJMSRdd9Vq9tZfawoI5Ru0MPcYkXWi0UvBqJXwly323O
6tZaI5A+kXBb3m91eU7+S5RJoO/UX7ENMpGE8Izjde7IROR0UaCvvchoyr2y
qAs/mvAY2sm88W+ezj3zCpyLnjc7PEruFjbCVCiIhPKgbqPLnrHwsdznF0Pf
z92wzVK2/8aAP1lmVg8msvI9VK8fSAjFKQFO3iCHd6mnV8irwS+dyboZ7RO1
oMMmO1jtjzAFUX/kSL3hJZyH+bvghg83tVmd1GKyY5FcsK9Xq0boPvOoXk/D
vBoeTYlQPLTv+ani7IJ+Caw93yr7i7L38WHCnEiRBQn6iwgr1L9wvnj0XR4l
bjeyjE1mDtH7KeSIxDkYzzt/D1pZHKx6vFREAmOk/IoFBchj5QCpnTbOo06t
Q2BleqnN4c8YBVI1hOVfRviR5ea3BWftfjPzZe4ZM6Ql6yNe7EFJj9/JG1tj
/VEhnjT3E0hNwy26l/CzfqXp6kz/gdmbmf1mqlnZl09RLtalwWEelwiF4zLb
aI7holblFys6iVzmjIQLopoGspYu3Kfy01AjF2xgLAtJA5meoszHOMLogCll
42D6uZmx9a+Nhv1TUL/iSuDbrjEv6/2CIG+R9CzaEB2vJEVgv5MfTWQRawbX
Nq67PhC3reqQB9H4BNasbzAMZDoOvmrStqXooMhglkhQgOYShBWBbzla1AhH
rqkQsBBtqz69U7wmxsBEesCYBPNpv2iz8gchMi3P7h1rSaK08+F3oMPJm/EU
+NOYeUhb1vSwikm5ai2h0DkK3mHU9p2T4yHbd6Y6sz4e6wB3U1gPMswnZkKL
FBQbeK+oaDilNP8YDfLO93adf2bp0IKgvuX1NEj0o1ON5v4erc7wHTPHycNb
8nIn2AfXGi+qBtp8M7dUyoZ3mASJdLdDZ/XxhOUSANDZzgca4CGkPzAWKkBD
d+Nkkg82IbLT4AVg3gd2nnIjq1gDLK3oORWRVFkEI/EX0mbpUM9Ky1xveAPD
STsW52oBMhPqAjKnwY3GjaffYN8zsEuYkJ4SQQ1weYzqNxY8rGK6vj/PE3f5
+fGOOO4mHmgutwh3VBYSkyLOweuApUfpDylrWUp4yOi/n0wQIRDrEfUINEgq
feXa+uxyHpGnG+MbxjQvrzvK6VdQ3UXEx9QK7xmQoHIgN7QDz2esKTiE+WEd
0IAThx6BWvLCgcfpOBPZYoCFg3dTz4DWWTjO6tslQMFIV/gtgPgAyWx9fk//
eNsELp+LvqIfmx7vuVrao3gYOZ7Lz7+GHVpdldkKmqQ5l4Y5S0BnJ9hn405k
fCwj2T7GIgSQ/f4D/S3xsIirUdHMoSDNt8PfI11gEmljqUvU3taIbD3no4TJ
TR0Nq3ynmbgOrP6UqttuHRzxlZ/9DQKQWDZIK+IX8dj0iVQEVTZbS/5hFvYi
vgC8lEo6uCEheXdiuEQSLH07/5+wLro4NiETT/PeXucg1RHPBv+JbvDIqvUC
WuxISzQof9jozJobEJIDYXcVfQ9ZLd7ksNjBsMJqbvbdEyz55E4YXdKGzaUs
ryuzrPojFcyIjfkjx6Q54FiLkYGs2uU0RczgjT+MMyENKfmBfH9lRGqFr46t
9vcqm7Lrnx4ZrfzWPZEede5NQnwfI/uZWXZJBimCZD3bjbpL6N849lpGl7CQ
U2uG+RKJ80wx8cT0PvndYcRoeZ8e7PtNAk9LlwAxOfSB9mcPw/faJyAhVhSt
B2j2aIH9VmGpHhPMzxlo4zcutuL5fnH2NlVm9XTD0YoYSpt0LZXqTj50sDC8
dgBNuCA6duG+nq6aKItD8RfTatOKWpLxGgOI+ScHLSfozAxF0fi/bGrnnjTT
yWDi5kqN6kew20lFsf66kZsMRHAIwIoFdr1keDJLS4I13W3Jb6rbZQv3TpLG
Wy6JJcJyGPed6cKBYgFzh1VTE22ogvIpksXAwG29ZPvA3Q7GSbg7c5mzKKRH
+jJ4tTFQONQuPCIC7s1JsBt/VualDA42c0HjlqcoZX9ynQRYrKJcC0mqjSSc
7ZuRQ6r48vEcDfztJIBTFD8VU1b0vTSooaW2KB/H0Gefa+H3rPf5bVDmmNuI
wuOwSBFyvkVmf8c0/ZmK2qLoEeu23BV0+vkc8SHHrJZMc6x228zZt4u3Wqcl
rdlrcfSAbazeHLOLUOWbtlfBwVzhI5kX8JuwXXjJU15W/B3GwPbiGXN/leU6
vJtfgpVU80966O+DwfPjEXYZ5NjmXxc14ELw+N8H8kP5dqT4TbsOihubm10m
y6d5O59TTtZzDZxpRPLV8uppZVLCI9ey6Ime5zeZKexzMCvfEP0d/lkSSxhy
2ncDpze8rNmHMj3aKumSxB5zhy8W3UNwx28kIPuMHs9Jxd3HUtnA9w10Pecc
uCwwlvMvHGiHrpdTB+SgyqHy+cfRycrRIlyfmHi9L5NFSXpM+fzPjJziPhTF
naeEcd4l5rHLWRQPZ2D6e8ZHmRVqYcUFv+V2B45ZcfSivP1/nYGHrDWidNgr
bb8eLg2qKlmanxCyDpHnxFjEEjt7Qkv66v11uRKqsikRK2BbLZ5XqfnljL7B
YHSMEmTBeiiccTPGWlgc9si5x6QAQctvJygSiYADUOZJfnV+VSAUdXxEeknB
s6ihlBcOkXBFo7l5qQo+b1JXWTyBoS+lIPxOrvMpc6Jvo9vVWEQxnH92MnCW
XvuO2d3kWnE9TNLVQQYNHDjkHhobAoyGZOJ4qVGhnmjMtMUTDCVN0ZrltKym
cuQUb/zuvqgwa80OmBVk1BU3kJ/m32LbLu33hk8owPqCLWrH/Wsv1MLtxASJ
HL34tQUMe7bsJEvmhYkY+0U543QR/h7NSNmlzPw9w37+ZR6RK13B6Kr/0Et8
EkgJ+23qq8fRiAelilGuxYmHbBf5B+UXZcBSjL1aFJ0bswKJAxX7YMirTrc1
ZnfalPAiscnyQ0tyWkswo3Q3nCZjZNBp4mygk6Qb3DrNYvd0xILnhaS4GU7i
4x/XnPTWBeRyC2KBzYlfX6X420XZUEYt6B8bo19y58uVm4O3A+2xY8hf6yC0
+Zs602Nm7hrNjeX9fqUG4mVVL5q/O++kKlcQBeWxBmr5iQKVQVPfNzharQuu
C8tL31gs1cUcjDIO5/EHxDdeNwu7lpwq0zjovIcXlpzIa+MKlqixIsiAg2zW
xuTi9tZCZj8kVms2e4fFoUMeFtjjy8wOAl/A0xs9jeMARBnuTelLVa32fLGy
ZUPsWP6SMlI6HtxBwMVluDdI59/CN2ZcWuB0tS/zMNrXD5XI4h51t6UA0xkd
HTPmNf/gim9kMnoXtN6q3griiJZi2VW14vtsxgwDlVXzmsfa1s4GI9p+JXzF
9L4w/BFlCvrIdlwkY5KNl4LWwi6B8Ds1VGDG2fukPU/XhBFcBNq1klFLeN2g
n3t2e4BQRWAdnVts4CQaovvSHcqgHeQ6FzLcLTzf94vNtIZ+AIobLjdkCQrf
2ag80gIgA2qPW5fIvgbWT8uXDg9akV5dVgIfDkl1Z7MFnAkq776TNymPXfwY
OcX2+EcVhuiFud7X9835c/5AhXuGYKI/uu4BIWGpC5xNVLNnvGL1vMKY+QDa
+d8KKyw9NWwhcPCkFK8t6A8l2E/LZaEbnw/sqlJ/gw1hRpjg+1BVgg3ESICo
edtkgQTMcbP5y6sRShGGodmzOsiWSyh5dVm4EJqsJZsOwtqrjqTKDrAooUX4
fQhlSJ2/rfwc6hxg456lZdzaOPmRlbwjDnBBi8a41RGNYeBIJ7LLFrlr3Do8
jMURCGfwlsO5ESafFsygTA3yu1n9mkTd6fG0Ytz3fs+YKNcdQqNwQIvNcl4j
yH/qThRtZYWkvdey30P4q6aJRPxvNenZePdFteLz3OY68mO+JKgNz3WCoZbd
shN3ZJTIx7J3pxIxqjFGpyigWe8XvXmF4TAfKqdd/6de4GyqKNOgJ6s+hkEW
xN4oRb38a5rVLxQ+wFDPjndwMGDN0r3CDnH6gryf/jYY89IVQwPBPtvAEEjl
Y0zMdcb2TmTGgHFDU4XSBP6wHobEUQXUVJPhlzy8wMgvJqBlpb3XNTql4RCB
D4EbrNm8ZgBUMnXgagd9OqsqHqPx3U2Xv2hY/ArxVhZ7wmoyjFKNLKVjV9bg
OZ8rxYpkuC08FnzEABbEolXmnRVf9v+DPOB/7YR6zhC4ea9lIQWfJ/1eizq3
/E6jUYlcYX9UpWfAjojmadTmW/uHJ+jqmek/aYeomQfpJvjkUL/NxTZ4vdZi
+/iS9X4SBJPAostSBpNiMWa3qGANI3R03NceFitqVHcSPmx6bTBpvulEdWlR
ZngeRGlId2+6gTwygMuzzQe2TGJqsSh+q6R4XRvk853dmQOeCWYy1dUBSzPB
G5Tb4l7KZDLiMNLxedNEIN3EFmdKotpH0THYtzifb6ZZkSARMqs/V+9F41KX
WxgAE89GOeudornkZ3XpJXQvgC6oMpqtb4IsLN3Md9vImhukDJxpgXsw4S0e
V68ioSojaudhoB9NcfGY5E8m3oRjYA/APgeUqItywjfLjVDcz3VsJZnMVEFz
Uzrlb89dwHJzk+niL5a1jULQAdwGu40n6i1gUa92lZQ0GiwkDYWz2PJCEoY7
isp+WSVEuDCX1ODoZMKC9xxlIwk4t8n+NHzaIGxaIFcTQpLpPhosC8QJqCqh
cD/Cz+hRG37IBXWLyGZHU8loRvNxJcfI3Ub9S0nABjzIMFg7hQ9mzD/+JBna
H/mlY8eOfdObrCO7vtxXsUrDywRxXXrq/C+jst9UvRaoIDYzDWgUL076bQgT
P0uYAaRc3111EQUh2a/goL0w27GGaCNTyOtDR8/q5LAwaNvpTjLuC6/7H2cT
qrZEmTHs9ZyOwmd84p92yKFhCgIa17qnBoBweuq5yKgdnmoigh1FPAdjWNFM
+97B130CM3mT86de8M+CoGgP9/Tw+epQoGi7PWlxOf2oafooZg0c7FNfR3g3
epRi5OgnHvalPMCyYW9PR2H86r49jiGSodIufU/UQH7wHfM1W431TK3iHUuA
6Wt+Zcj+jxxH/6zkLhoHFWz7y6d8QOIEdw/b9l//9GEWIzmaJ/L8zTVmn1sK
HdtZTYgvneL0g8w81laOLawv2PD1JV89XLjYvnUKcG0UcOY/MRyGV+ngxaSo
Xyss7D3ncyf+2hQTqMgJJcpe/ooL+HAgvgHH7Bh3079dHTsNHMXRYXnWd5RK
3yYGwofV1oK6fzfpSEgbiHnJ/8dKk7cVo4Ds95zAmSnmpEeP3hDVV8M/KbO4
LbsLc1qey4pNULegkJq6B6bow1ey4FAflll3vPe/+2aZPz0EgOmyf2xWElyh
Q2dZywTWrWZJHQUey29ffVRuKlh6QM+TOHIRMcP0u7nInhrs54bqyvDqeK/4
3pFOTYDlwG8XM7MxiF7Z0lB09NSjaf1JJX9tecmxTV9Dq1iogQ21Mo0yVhdg
2+ba0rq4CUnpmBY8FlmLEdBj5sy+6CCnAphD7Gfs9pH4Yjm7Sgk2FjXdd+yV
kz44+Ztjmog59n+/hC2WqrYYvpt1hIEvFPIslDCuVPWHS0JsOjokAqrYjS1S
mBB3YwmismK/XAB0lt9kc319xUESnHQk3rwHhlqJvz4NkG1F1Dr/he7rkYE9
+uOsNoJZg9SvgGnaJlL+glEMR0JleQB+fjhfns+AkSzKP72qWPCGdm0Ffo3v
67NTCzc/ZwQCdRV2brra2mRCZBAXVhB8EfdiGgC9nxJAo2RpeeHZWJufzRlG
Y9Rq9UTn+drg3njRfHfdgrfqSF/5aH8QcaYFq9PSd4XN7X0IpgDbj25poKWi
BC0CqiEdIS42xTMTLhy13e3ivMCHPEj1Mdfx71JlTaElOeHJd+LBI5ihGcZN
4xRg0AXYIHMk7vGHDMCR4T7zu8iyMgT/xuPfdFwqit6GfA6e9EWYyLrJGWV0
FoGF5M8lKF65nbpHPWGL++FpQNvajuB6RKz18GuXTs/ebQuyHYNkuzeaeaVJ
0jIjQZA2osJ+FUNYOiW0uePokVfjamdBYO1QuOuCrkhgvAZzwdRVQqQA0Qf9
UvXm01zdgsPQeFcNhqGrBLrkIPmlc62crYdxc+c0J9v3R4hPavgO09p5jFjq
89src+NRC9czrMAYWZ/7EZU1uHcsKOhfbrGXGBcksPvJPMnF3ZOK1THkCtKl
lbZFYesdrl3eYOf3wAUwE8nDiFddimlLfSKI/fQplkmJTk4WQCO8eG3ysVQT
ii9waiONS5nH6FcFLIGfKjTdG8+xNHdu8XtL1JGHVCey+OKwhA2jNpVkCDGq
CmmKCiYKlPuRyfsVOK5P88Jh59KSZN0eJmS7rK4+VptHN0njBbNvzxrAO265
HrZugu4Op7EwnURDnBeRbGyUinq32D3paX5WiFDC/7NUxXQvJPqL7I/o12aK
krRf0Nn+E878O+wWmRiYMceOPCxb1egOkQcxnR1E8ZZAd9VYhKs/xKnCfPbE
uHfAbbqnayDxkR/LHNbEXqJZrnw/GMSfGApP+7e7Uvh6OB62Ok6P6Kb/uWUA
DQxcxW82PJxz+3td42eLdb0eFmjsdOvzgnTmuAl7LlasoCttl9l1n2PNQ+4d
QcEZ8591+FdM0JXyNJSEgSIgVPMCdhn3r3/hB4u3O6AhmZt1FR+Ws6Qmw/E5
2qJjZPo4cCMNRW3BlXiLbfD7H3lt6m2/HuXZgbv40xz/pU8njfrdY/61GOX1
koL3f0Ae6rofPgUUOk/qxnkHQzUl3TpJTwTZT2hifTmG0k/ugV+Il2wA0mDO
U0vFzxHO10vyqB2Qk+ZQtpdd59vrWR42inP4YeWW3PmZ+W1IN8+EvXWruzOi
sextCrBio+lnsqV2ZQmvAmOFi1sf7RsIj05hVNE+xlNxpycQoQ2WPpQJOFpe
ucZPwCh6oTQ+ESgwfkqkEjXJTiMnr1zQJliG6vwyPF2Rkyizfq6AXuFtXS5b
URFLO9V6yr8VyB99tydzedJswNLZipBotkFWgBaYMKw99/RVbUi8ltonGS6R
mg6weIbpTxY1NhT7s0Gy+qx1sjFXx0DVp+5Jax/5zSTcpPtJmEaP1w4ARmQD
Kld0DB+QolUdHPZ6IyiSpujm0s49ZJuvxq/LiM0WAiWdjqZsKUX6YCjoH3/s
AO9sZSheo75FdriqhNXQ+Wd8Os3CvLpI9f/sT0C1OCndDWKOXq9lYlTPmKtH
8YXJjTrCTweNXpieBa3nCE2b4OnCYCSmVQmaoSXtk/6wlBNI1uuqN3QDwzrE
eX5jaym4B2+3Tku5V6WKqUvXKt2PeUDrMQi2z+Kt6iJUj/sJSG5poujMrYt1
8Ooz0q/a+HCZ1pKoQ/+IqdKn4j0jydL8QmTRSqIwhjNZr6V6Ivbi5913fDPr
h6iS8k9UtuwQuRnCbccZpX7OjnvF9B1CYvsqGGTjLesv88mGEVARG27DFghb
TFhiiDSzTgH1FSd6aQYPBuTCW9pqoK62mGGcaRdN9Iqu6fjm9LrpbgU1KeSo
K/Si26167Pr+78pwEc7JQ7nxRJbtz4h0U4xI8FlZCRoMo7HhvXyBgR9R/43I
+JG6vG2hb2s60w3ouyujYwIeo1FBS+YISqzBy93YjcrdzGlVJcKoCKJIjYu5
dRA7+PLiqV307Uv5H1XbE6mW5foeE0sqUYxbSHSqiHj+c9GaVcLtvdww3E2g
nE6WxWm2T3h+6maSY+c2Ff40eEjtLetIQkXB5IXyrL1vIbbe8C6Bt8SpzY3l
aRwG+zxLmGCQQdU9GTJT8Em4+ctZ76LH0CMskqySQciJgJYPFGRBoyoKExEX
yt0eIQOjHHnlZz7yecoaumeqQ4lE3CyFVwx9s2OLgoSsYg989A8WfwB6pk6Q
q9jh5LyQ+4fEKdG4m3CCCyV3qdWHGyn4LW4nq0vz8Y99nNlqmLR3kG1JU5Xb
LKhWdNx/UrHhreuMLvchyRBuA9tlcB//7P41k1a/gCfMJ59KCoG2TRHT6E7r
7UacTTJqvGmnmPEcri/fIIJSiRJKC5dVOwr9GfBat31ONGLR15J1Eg/jdCwn
sSGNIqb/AtQpqOQgXzZUW0sz/mqctSJewtrOaeO2Cl8GZljFCGco3lLSHxp4
EPzmtIFFpVjl0upR9piObA/KWg8UbZldJ/V9hfjam49iVpn0QUhDsA8aKirJ
AfzdX+Xk+GXmDYo/6Vs07WFnYYCkHmgKDrc9FHp4BJRMqLnmcbKRIxzlbN14
X6rruE69jzGS2twDsZG8Jzx1rPD8xc/mjMrg+UFvfwyTZkcnRdshkmebopbZ
g+387scEeuGncaIAnz71m5LPe1Z6qCTnLxab3R3jg41iGG/TTuEZ45j4b5bZ
EtPikrmTd6CLT9NRZT/CiCsFSzA53JvSlBbu5a8qhD7XA362RVI6Kv3HpXLG
MJxm5jxxtn8jM/fNiLHgDR0ToOhAT2iulixcCUBjelyM4Ss4Gki9q3fEP23x
ZTWfmiKIEFgytVQlvfketENK5BGLZjO2+6xXZBfcy/Qm5XPpoYhoFG0mWT8U
exrqD+OV8hUi2W6Xxf4u6qwI2h8LbGiMPzaYVdCT1MWDehhQj/599byqR4jV
grFUUwLZmlid4preSi7D8TcypuOpproYTER1uhJ1bomEKmBPq4wZ9gwT54nC
NR1Ngcv3Yj7E0B+qYFAzWMgHFb0qkBFMeW3CEeppBTYmJaj7Ia7dYq3SZIY9
e8w0s7t++ZT5eP6X8XixF4hj144SafaOuw669J/sOGsph1pKWeLEKihM4T0a
zyeaFeOiP7XfRfY3no/v8dRkeghoXYdTXzDihrcdt/I9q+5tl9manE5/2uK6
AwfnQnJvXJjM4wlaNlqUduAZ8nB8PMl28JjjtYksAQYL6DxstodiTXxXidb6
8aMwFarbwWSV/kZAyeti61Pi/Yxu7YrAw3CcVDelbPzVeEfoSNgcFsdDqNJe
XVZXz2ImP501+Pu2fU/rrYmc4mVj8sm9NgDteDXcHJu4GAIKaD5Mje0g1PzE
F3xhQgLo/g40HM7KFyVlKWp8CPPSrutLnDMr6scAQt3eyzpeXPn8WA5bZTLd
/BnstpoCSlKZT+7nVwXcUn118IJ66k6ayCwlLBys6Y6G1TGPmnRGesgpUhEx
e+Xh5Gbs7KyE3WkYReaoGnF8feWRX9b7eKdUyUi6EdkoGPGE4hVwRQ8ktFKR
AmAP4lBjCwsExFUmld+PK/iRIkrnNX08eounMG8We2/0STB043kgSzYSS9Qq
nAY9j6egVTEA+Kr3trMUczArb6Vk5x3DB1MnWFRLYBljiJmARIKDs/R87Rex
u5tXFN5snlCO7wmKk6rVZl9GILD3Ist0RSpAoAqhla7ZF73oEkmxTcCg5RIp
1+fUItDUeb3SoxatdN0cj8oaCF2gpT6Zwr9z7dQJC8EGAVfpdxNGeG4dOStO
5Sd1qfE1eRrgKWpAg4GxkBQytexNkla+qto5slHeKvMvPdVTV3dUkiX27WWv
OcrtVJxZ2RAwzZ+CquNY+4zeXy0Ddx5GlFOFiV9FtFVHlLCEM19Sji2rf4K/
Q4uOv5kuloKq3VxHHrksvD3WmMQmIT91jwQ4uxmNWWn8StlE93glDBigC7bX
X3Z4I+GecaZ7B4Y/T+y24FdUrSozr2FdLpnxxPf+H9vjI6NyRn+5WRK+CDox
G/V/T2RcgG42FI78TrS/iYdNyRuj+9EI5YFAXxu4j3sgF/x9xsFOj7IDscf8
TrpDOsYJfP0fCFWl9do7sq6bGVd1XEOAZlSxcBc6sB+q+4yE3AYl7OECNsi1
Lx8oUMJPals0cwHN+FLoK4yIn8ODHSXNznA14sCxh7c1GUD2uaolbZ/JtF9s
ye5RGZ6KxqEaY7c9dHV8u4ioSyou64ZYUbz8Lk3mn47PXH2dUtdjrcPCc0Nk
24Ga2trobx75M62ak5G7C4ShVMC+xf2hAPVY1Ul6mzimzy/25mKnfXuwTxSp
BE9tfOPWfFbo52fP1qGfTxaLj28xJ6jZxTKH74P9H7osaDCLChzlu2w6+JN7
y2flG/a3f3Fnr8wIbDh/VrZQ1JfzTQPMPexTbk01O7YYEo4cpwiMuXC0pKz+
2ch0zTS11/IznrAkm06/XfyGVrIlUBwNzBODJy0kSXqlsWWCM27V286neUM0
WVYd1tFMY+wUClrLSPKIqXsVfiwD2PCiHccci24aRDksUddwBivdb7Em5bXS
fK2BVOyVElySqRMQcUJ0WFuGQM2zDvBSXl0i4XXxaUKCS2ITLz3Bs8b0uv66
HvN+KvBoG57WIBzyGawYAOYhqR9zfF3hy8glf8dS1B3wzoDOQENL5Bnm+lsV
gHaA0mFHk/rVjXgMrf9lctnVxTX72cfQw2oGPMLbthan61RCgHv3++lVROlp
OfIDIWZEdCNswdpIksODe/q35qrF4PobBV2hS1DFW9rr5tkACww09aQadmlD
75P9t09OX8mVHBIvO6Su3ozduLhINDXZ5s8aHSu+3aY4T/+pjCNBOJzU8gxH
crnotuIasN911wULbyW2j0R1MDwjt2gYp23J5DDG6smb+VotuXHzmaHDIruD
jQGVYGF0bmFkzDjz6knjMfueAzb4DLgeUkLZF+TKw5L5eS2yKYb+LEeMy7mi
LS50XF3cPQDazlXQbl107Y7g18z2bfNR47ksx6sJgZzqcJUuFSCZsGpwVvrs
uFRt0dQ4u8nQxmOxYrRcoZsHWlzht36163H2VUfsgoKLUJkMAYkp3vjTHN+K
5HVUeVYfywkDlO2vMeIALvsOj2EuEphjGQzojJxGE0J3s7OluivJ5BQqbt8j
JkorwS+iZWlCYeXCFQtxhTxx5IKMboVtK/xtUJjzXfrQQZSRJFYNWifanfuV
hnSqpqzLOZFG++Zt5Bo9mVJ8uM6jElJRjl3f+8R6cZU7ArnY+1vVl55++0hu
OnwDs3gADcJz+nIR45TZX9jk9c8g66ccDkmcr6+9BW7sbLyhraO74yYbkgCE
NHACfI/gjQ84NyItbtVywC7+pNiKkpF7mxpq/BBhY1tKsQIiG2Ak1XFGFPBY
oKIkLAZNfKJsH1Ul14BHMpgNCTHR/dD9xgp1a0eP2r0NOneN1EKbnuiGb3R4
9f7ElpYyLdsZfkum7k2AN7QneGnzsAI6eyhXpFQOGWFnmZFVe3KhP4asK7Yg
ODRxtwKSIHTD8ZkrZ2rzzdt8gMX9Q6ASKiiy23suWbAEqmyw7ivE+MhmejRP
1vYHJ0A+hlT/PhNrXqLbiRqvTDjY5f3nhdD0Ziul3OjsYEMzkkCwAMHg7x/s
APf8rOidWDdVfIT15lk2leE/R6kDGcUL5QkW7ALP2S5emuzId+xHlTZ82hCs
pon24khJA7oEOVXNTSUyOhcnHI3s854+chTslPgDV2d2fMnAgKGwQf5fgbW4
d0HAWORal3LzzRmCvkMtdeshiPyvdMU8EcOVSwuH72wja76+KcilBisNH1Yo
WyxwQ6C0Ta2st1se0EgGp335bpUcuGZI9P9rfVACJqzTC2YayZaNo6gbW3pn
ohbE2Roih9AEInSfXGGk0+fH6xiw2UhCRyynyA7PX3SgO3nbt7dIvYJ/5u0N
DCL9xEsDILYIekwMvSQEwRZVghiCTM32e1ml1/FGtFTTOi45zDnQsqes6SQb
hh4i0BTvBR8brwlfHQudf46PZQlOGrcn2m2TKVoHbCzrfkFYZRoLybKCIxDO
+/3unSwqA9tvdbOQQgFo5/gyxyzTRXthgAP57O/DlwdsyIHP1hjv9RJrzxXl
gFwEe0nCQxkR0vyt4OqUc63C9/B/itBTh7qvAYJiXwz9jYwvVQAPCL3co2YL
znSmRBaGMITCm1ADOrC+H4j3koD00cno7fbC16tk/r4d7TbU+mjpTfWwPBAj
hRjkCuu5jYrL3q58t17rJw2+zsqL/kEZ/2Sj7kkLuukPIhDtyCBJbGeBZZAp
Qmftf6qhYM9GRorDtYtDbKWOVWjASpVwMEOu0DyPSKtdoBRyR21dXI0w9iZc
UVEQdh1z+xd7hlY1CeqGPOIqHdm1UyJ/j3nG3AaFj/obVlrJ2jvzDCqvdp+p
hHPiNZnP6S30Zbzvc5ElsK+YDUOJGV5u6pDF9BcYM4wfuMwGen/MJaUAh/Nx
BQSnphyzvpdI4FAbCjuv2KSADKOgwk+A2Z5qf2VuhlkGbUDiFmpL4peTVLu2
yNVsB7H7mr3bnumO/soO8/+WMyxszu4eanIxKJrS6Zju88CrnQceLBtdJa1A
g5C0KhHhHv/R0alL6bF/wSllrJB4Wmf8veg4OSWELCwmtOnTIXaS0EnwyLqX
Ii10AytXywEKCx3d1LVrr4wTrq2Z6jWcqNoG6HjzeJ5+TEssAS4/rMfKa+dH
jBML6aUpPhcul9cpjE4vxLPsPSjn/Gu5KbYksM42yZC/xf3BIqalw5KhJ1E9
fpbppckoDP7zK3qzIdCR3rGXA/MvdojPsxFD1zOBrr2RbUIreHB4eVZgJzJW
5EF6QCAiuo/HVbLJ4MZkVBY3SSxU+SpbFpwwR+zAOlRPyUU/k3ak05dXXvVa
g9xNrzmrjH/MFu2HJqtXDn8jQI8AyeT1IFBewBWywj+ikNx4ESi85Z52kyKM
A3XZTxYp3UO4164BNNijLdIuuMTCzKLbD8Z4Pes/L7CGyIEtMuEqAtEsumCs
jOAPCB/GnCGy01lEWgGatD+MBfJWkDnTXN4RBBBSG9uh+vEPyqZSBEpNSlab
UUwIPnB7vThMnnsBQqZGQsQDRWhrf4wpR3pgI+Stpi1qOGhm9wf0Cvz5MCIB
rU3J+xbaRjTOmtpcVh5bSQ5nqfrIwEAq1CoYsMuMdUM734RsvvOF44jetle9
X6qB3ZpwA4EI/9JZDQBdw7l0gp3SChyO8/XFNXSflH6fPaOiOeoE7H9x4OCk
EBSveuGrW2F/lN0yxcVa+2aKI+R5fKSzVgRMQX1O6rV44OF/DS1ZKnr1mCFt
lcLKf0n4WFuC0FLG/HNqLU+pnYnam48WmGxwz0QIzb40eotCvO6HT85AEioa
4DciD7LHglCipAvimCYKsaZVd9vALAwMYMyND5jix3+dzWnjqg29DJdyqf8o
OyAxg+iDBHe1Db88o6V225bVUgqoltCjWzpKHaCk2/HmwQq454Sq7/I3M80F
K2sKfNQTgbPcfLKiCWfPoNr7kQ6uEtDRTbLc2WO23WjdLe0+Kdfg8fW0bhx4
YgqryATP7DJolLlz+CNdaPnze69/guONx63KAJZPUghI7iYLhnk48ixes4jZ
ZQKYbVIFCO2h6YNUIlEo0gAf58pDlKQWGRnQUwrLRzYF8s+Q8ERsT1+lJdVO
uMnEPOO8aD379RPC8rikLY/xdE+CudR1dYYoirisRhytLxuLHkLB38ZVVYzk
kuQCPVP6rFhXeg63MCM1NmvXdjeJvAcLoVdaW+kyFASEbcyh5DXP7KOz6oRt
u0hmt3IoxdGMT1+1XyAqB6zPgrmoxPZNq8HqL4AitaitFu9j/Ig/M1MMZ0K4
K+Nf+176jR3T4AE72UyJMh+saNYOnPYOF1kqfKl0M3wZvR7VCW8nkt+v+z+D
d5ml2+n4sv95b0YGZuvlpbdbY+RMg2TS7q0Tg4ifJ+z0d0vzQU/tHss6yGnm
aAcBv4HqnO6Von4GQG6UdHEVlf5TwuW0glN1oyaJS2cS5BNMCb5rLGsD0VsY
I1KJgb0CAeeP32sim1AEhzSJLqT6uqehGgXetyrIp88nGPlVlJbZYXGPz2sb
0EqMyAY5E1DW+F//T14qYWlbrewLS909GLBnLyJwl/iVgYul8x2t7sEyXTJr
wAYh40MAQb+JfFjsLYztxKhsMKlce/KZjd76PUNqfIK4j5KHiJ7jcXbNFqpa
knN9OhMoC8Ra4F7D4QbxE9+OqDM3NXKDmgNEf8RA4zdFLxYrurPOICjdZGHU
bcYYV4HFwQRwb7yTtUk1UxDbIWHRkvnO14qFPKfpqfzKMdUhJwlmYsHgMXqq
Vbwhr3sW9EGe1Y82p8wHbqjcx76wQeXgsEusi8OVv7YUkMdIxQyDkOLR2DCq
pXjnqHZy3bFprjklrf4GxZT0SjhHlh1gadivc267AiMn19YaDZs1ZV/NjAn/
cQy2dO7dj2Pf6A7nk8wvBewRgg8vfpCcCDcASGYTPerI1W6LBQyj/AcNGy/Q
Ofbgx4c/nUaLcR6NU/DuSb6iKhrUL1MisYLg1NkvH0moH94ieBWasAXs8RGp
/7vNHLnl2JSGRNE3rhJBrWValEvCy4UHQEwXCDUhePwMLpGYCdHlti+ydD3v
vYtcN5quXaWICdUTT1+uaiie9v1zbAbc1UZu0ljIDQnPBLbloJ6ludabqJIq
7F1VeeOxz+l6VUkpXPG3/2RN4OfcFJJQ3FL/ESIQvMGYlh8OIf40qazl2Et+
vGT5g9R7hM6EX75+z3WzjRMrBNYG672GhxfA8w96WdprMV2kgDtGQftonHpJ
linfJ2fdCiOd+3lBBizHV7wWOPPPUGdmdvGcrM2j13a9VyaVPZ7d+S1RSfJp
tdyRugBeepWUZxdpD7bEdzHLYnCypIzzsWiQ3Jn3JGdkkGjpU2cj6ZO2qXSW
vJPUl6lKAoDi8KKEp8/rYfC5Ag+sdhPmlHlnb5q2NOmTO6wLX7y3ak+H6SfY
uLcHljprE8OHxIzdluJRhr2t6onrQnOpHsJBfzc0YvHukJlaCrnEbCAPfyzD
A3OXSu0xE7/kJ7sQWnFVDtZYN4aMG9E25qLG7b5YcRTRk269IHkNVUlV61ry
MpXnWk/Aw0+gtRcVMxqdSSpvtnuRWo2CTdyMLdCkIDHH8E6E5YtZiDaU26Pa
t9ht6xavet1SlfQYEXjoxK40EScbSNbUxwUI3Izo/JJOY7SgXHwCUDYceiQR
HPF0nOnfT6MBUAKsFOkV3lOy4baSfKb/QxPGkSZgLyQ7HvEWDFAR4PhJnZIB
ER4nRHG8mkL3IAeH5zhG3U51c0SGmXXdBQyaNs+9kXKCNMBPNrx/L17N0sXO
PWkNL6n6l1+0DDD8vDtxAj2AnBuheClQJ8rgGCB7NQumxny/R4tmv/1rHdIp
hVlQQisyYJ365MRouXKkgSbuOq2/9JJLyCJr0yaGRS+9UfH/27v26fUYqtJJ
tCAGsvJGeCaklPTWjPpdmNxsajZ5kK2KQO51lqnuw/80gUPRtzSZ7c3ufWhS
RS/n2haq60jWUSOiuC9dMq9y9gTpJM2BjgNlWmDwRm4+EeBtnwSZdx1rhlbO
eye5d+biWJHfsC1BE6UmX8Xxy441LjN4YbAmCZzQ++uonHlmyC6Y18Ju++sh
Ks31Csm4zo//5WNYMUYN/Y3HEjEc/GYNcUVHkSkC3rLGVau9d5xsonaQkYdg
S0Kodo1S0AdZGcy1gD6y34WkMWlboXmrr/xq7C8U/yJJwhxrRxR0aCVq4V4K
nCoAP1CVIvkNL1Mdi4pTiqZlm/8/FxY1ZJmewYFiyonUJpohwGGpBG26XqbG
qv/m7QKFfig6PoqqecgZZldGXpKf+4jh/9SOuQuYnfFdYE/EsG8F76gLlCTk
VxAxUTivxjQwgoiZqzvSZ7LNoZkWJauvEA/LkYMhvj282v7aDCeGSj7+wVMW
GyQxpUNRVTd4gtV/44rzafbaLe6RUGJjJVgSPnWYoogpHOJeFZsw6IJq3efQ
s4EJ30zqjJn46pw8WGrd8DJB+EYETHABW+jiAPffAK5y091Y1dP4jxGgsaa7
1YD+zgsqBjG5ovrcx+n+z0ykv6ZISKfbPbdjJRmA7E99aA8cdEuNY6gbCGin
9QoShqIWX/lHDCNmyOgfQ2w/oFxIVW4hUaozRkRthF2AmZz/ZgApOzHrjDxk
PgY5s0NTlO5P3xEElnl5dkIO+M4KWA5EpnreKBje+nvFz4kKs7FVRuCxUda8
JUDTEuNw1Dwr9/3mUSiTL6rja0oWY1F86M2HdYmzGLDJ4/mGSxg9YVoieTsN
mLQD0OrgWpbG0C6IKTgdIpoIsz51Ri9uaJgsq3CNRncQci8yLxqTbtaI1R6l
3V97OmzCU2NbHYjc0mjV/gmbEd58sM/sDZwRJbE4WogFdMqoqElY6IE73tKA
97S5AIzH9Fbg8hkcuQEfOfNW25YJLfJm17rdHsQWCqD5R9QjVwn6hA84tKtK
om/UZQI5MPF8dfBcchRhtL4Sj7o5BTMg5TWvgbrJKQ/7f1I3fgL9y+CYijHD
Bz0oxlgYmBIAjrG/l/9gXtcjSgmAnKGIB31XhKUi5QBDh885qsPcEfxtU1SX
Gwihes/O2LZ+QfLI6qdQcnqGBIbXYSnNHY/g6UDVwAHWzDplyb90/tR1sxRQ
Vt6mW6n16pdd1H7llAHNG6WVQHpr1OXFtxRPTEGaua3FyBqOSfg/WtNYeu2i
ohN6lmpjbY3VQa5V2C8kOaqa8TunTi9DXi3UeX0YXhc8yv/2tkMq/qc7gRqf
D2UMqFTAqx5S1HN4Qyvvp1BRmsegv/8AFbpJksMlatATCQz2Dkv+ay1ig4dc
BQa06BcYCX/dAFgpCcn5BbELg2RdrITRPgNr5JOn8Ag3FAVOdJSDhlS2cMqv
lHGX0osjw9ycKB3WtXu7bwqwktKp/m2Db+MCh+sTO01n+g+a43LjDEPmP55h
H+Vj45Um9+IrrT62dnZj5+6M+t+z9eC1UK/SNiMU0zcyD5/OILKZy5HsZMlu
wB23WhmHJwoZWWwe5P4CPJmpGbQzGTPaoeObO/iuDGnT7krk6G2bt22ZMhxI
8hYVIOOz+Bp4hhxj4SHM8ubRJPA2hk8X5pUIk91cRtVVfmLzQZDeCJSZWcsb
/TClzTrOwv7RNwqMVBbtVmVVcAn4r83jSUVe74GlJyJC8LuWi3OIE5zqpS1v
YKBnEz4qrNl/qlyd4WPIFDrn6TwROO2pMFD00gWDlJw95q33Uxiq4nkfXt9f
4T781+umc6BuQASjQY2elk71Np5beHUTt6obGwXNy99LGy4ZVisV84mHQy3i
99/laP3MLA4A/DtwC/ebEVg+OGcmoo2TRX29pVgU2vTxVblznNJpGYq6fpxX
cg8Zrla3gE2lxPWYiLpNVSIKQLSM3Atc0SKExWvHh3yS9dBZLX0oWvtJRxuN
4zpY7XV498vV6NH5nBNP+kq61373aObIVP2aXsIu1NOi4+rMOY/7JYUCfKdz
Awc0GGPcmNNrBScakvPGMS15l3c/KvdMqDivt9lRT4Y+BckKDcrD5Kyx8dYu
JE1sTb8xoPsTnWwGWgIxPrGF8zTSP3bHCoBA6oqOLallfPEVZxPQ3zA6oNHZ
0rzDo4tZYZ4SCiWxq4cJ5ca/iaQHvHvYKCSX0CQp/DLGoaQSwyMytNcoFLQp
uAzrg3rq7159j8d/hTtO3dFrj+/xsc8xC/4k3q8WckWDHoVpqLFWLwVicWUQ
Vx/j2MQxSVARgER4OT1SHd2hww9ZkPLkyfcOgyG/D4Q6hWxcsRhvOnv6vb8J
BSygNQb37zaLYFYfsYLw5+ZR3Ty9xFKf1nJbBvK+WWLW+W+p9XIBFCSAVekj
b4GP1zp1NTrzLKXx+8Y/lvrvCOe6v+s0g/oVzNpIaWTZc0fXpNywnjSfNUwA
jsTndZIioZAXYewnDrJ+53TUNMLqcod844/XmmUMOBy3DMuZP95CrFoIyLmw
NY4mIESR3ZzbGWA+AryT7Dyo6mPpOwINDnjCDOYxzFNPQ0BCQjMCtZ4u7JS7
3TqybpItmgbHrQ0en2Iexu5G/XfEbalXqmfzRaOzeJGmvLYerc6GI2m/zdYs
DGrItmoGUx8hnyldlbhl9fnx2PDQXDeYS8cUyJKJkpf4YEICkt6vxPVo9bGI
ItVHXK7kyC9kj5TYN1rSviCg/5lECAPpdmqi/Del02PG5U3CYwj6A+HMtoxq
82IiI80spfKEHYzBtnf6Bt04ZkmuhvUBApByCYc1AB9jnjZO3hGPtqB+/bxt
eBFxHfYR3TF30I/9zh+gwuGA7/PlXv881nOWd7ytKqbAn/ZrYLndzd7lcgJz
zWxEU1IOChMzKYTtg5W7CnC/ah5oUcqXEQbRvuziy8HjYxzBfqlhmO/6/62R
wRBxshMTFRtFN/ld6i18VGe8PUFbXVhSMvrdddXvnpg6PqmuURHa+CzIStiT
Br+5zroHnlCfo+NX+J8cOOJ945RI6uX1lk9r761GE8dntvhSSF4hNHJbNuqT
rFC2GR9PZciTkKzY5lxyhDsccthlafEhuJdGIoH1HZ67XagO9jsRMOtcYYtr
8xOBK6fB+0j7/7od7OkkadrkgFy0y0wXLbNKlWV93ux+Hz+12sRdDStoWmsj
iPmOzrijGUQNw4XtuGR1ElK6vZZyU17obDREiTIaa4NruYSka4zBUIQVH8ec
TlkMBga8C9VdfR0jH2h9wQ97EdShTPDy4x9v2aTbrodl1T9KHS/USPgQds8j
xx7HhcC3BHN0Ff4eM6cycLuy3lRDCExEkGsOYF7kaBnMagHNN2kFUircV+j+
pADKLcX5L+4E4qSXcJQe0m1brYctrwsKEfaaKUg3Kv5hIK28z3m5dcNtSZXS
RoH9bJixDDEqnEAAnIBZZwp6W13Lyi25kMLX+nwBoV/QjOHB/qqXtHy5YdLu
vff0dOB39Pv+80n9avrqsQHdBR9VZC0GOcTcuVKp7coYA9KGvtCVwcm1iL3p
s5cY6k65PRRNuxeC3M5sGTYBXLxnma9gjDz/ZOmCuKOpfTBldRVxc8wnljvr
mnaUN6z9xkKncH67hjIAz/DhnpAS/Hh/btB36X9SiMnvn5/gmREL0ORyEydf
8nnd3UCQRABWF3X4sBCWcvvV04tV/ljfnuzzNzEslWn0XFCG4sh/4+2RT38l
i1nScnB9QSErYRecIV+qPAbrJlLCUP1vspJBp76maCE3I2cdAYdI9yEmuvOM
xmqOsU5izLGCHpNFeuWHl0U4tdI7DQn8kCMPUaUJNfzJemvuU6478SkIXPz8
dNskh3BW00ZeKfTonrCzdH+ZUsGWVvPhGilDfM6QSt7xqmS0uGYVsWIO8GI+
3Be2CUAIa1ZKP6gbUQ4s1fZrgBR0GPnPsEh6msoxSSBzUNFsWcV8t9yfyJUf
/8jF51vzZpZpbUXkyNhpuiLsdAqA/+AxKP7PxYu51VCAOoDXi2GreMi7LBBG
T+bXTTYqrgj8IEmglgtF5O/kcYgA8lJjNlDT3UTSAbt54AYaTFg4/Mk5SXJs
b4twDmvOiij9da0HPZjqiUJRSxD43ZQC8vhvUdZdzbxnuFhjsTWBBo4vUqwD
OWyXHBVD8l5F5hO7nCjaEmSAV8snQRWgB7Z7CY0sV2n4eIkj6X8NjK5EkmKC
dDH7VDMfgD6fJ7sRbMarHIAi2nJDzRqASQRVCArynThCgd2mC+ex3ubzHonx
XYe5d9ATuNXuM9p6rK4TQZ7Iv0MNYsRhcvgXo1I3QfDOFac877Jo1rJsYip+
6xu6Px87G6f5YTSqdAhyx/3VD4eS8UPOJr1L7WoKwWgxiznV8xEON3SPGAO9
o+1CY8nVp8AMK0MRQTtyu6Uf2FFAoKfefaa8MbIwE0RXtmf4NON1oKtLwUJ+
37Nnm6ig0It14iTH01evb5/iuLyRr3X4pDxRIDwpB4Cp3HilB1nFzhRa0u+v
GMHSnXOpaBFF0umrnGWvOVadG1uEhZ4tInua4ELg1JUJ9Ski5Y8JKb6WO5fD
VGA6HRltjZiSz6cqEIEziZsZPOZMEFLQ03GUecpOyR41EaV5bRcuNl9WuXdn
1h2hR4/5mq/kOOqsvcHUcix0MZY+mAyxtUEFqEIFD8lPFvCDrJTvZMHaJd9P
gd8tgkuo/uFYZoYqDoWH65ihfwXQIdU5wyMQImcVIcaw+sxu0ybYonP35MfN
EuNKSsITLjAFXLyVeQL7rM7CUZkOHkPDXiMQr5MaxzQyTN66NKBbCASBjxX9
b+5x4nq9gg/lLf9D4T15ldFbSqaAzdOkccmbJ7YZXCjV4z3XkJSaPwzA4YFx
wMyRrL1bLPTYqLD4oo81IdvaSi6GtooMs0fxAew6ruHHxfDK4c5i+iPwQIsG
/LjmL6WYW0QeoFkBjJiRnE8O/wXYExm/CCDH6sIs1yJlJaRsmoMnxSS9IRVA
ffofqsmtVawj0Qj9yny5aVFVdfCeJ6fuc24hA/UMdDqPZoxtsMEW8lKh0mEZ
urCBV5grS5WIlVjGJhfSzIf+ke0YzF3cRGMSXCX8L0rGxe88Mrl9SyVig7Vl
6TA5oiWKCE7eSXQJrhlJ0nUXCsRE5bdpU6/MZMDXYtkrK3MULb6sDGIZNf/P
JFuN39lVWOfSrbM+GBhF0RTyp/5J2ayiuizhUIe3+cyJlmYONh9gpjVTCgMm
oWbAMZFb/VoE2H/DRsDSh1ijcDHqChYZh0qTssFmjz6KR4eH23Tb3IxOjNFl
qo86dIPhFdxNJmyr7E2bPn89FE9My70S3h68Fy1/UOASED0mWAAcXA3syBsQ
yOo6+MoGqb4g0pWNoyljgqfZ9Trvwig4oe3GiAG943Z9UFRrxQpGteg7PqIr
NbGPPO80hWcL8Z7O3W3J+Gn+NJMLxTE0aDtLxIl+g+OHVHoPAKMM6jYO8Op3
0tzz6WstQ7gA1DS1HaN8+ffjlSyBs4e9CvAwppawtn3QfG3fB6PS8elvsRrw
Sf5FvkZe3wy/SaQ3ladBAED2DdeNouYwMGVB/i59qicxs2LTpnyKfozcYiVl
AxQiHLx08GBxyxoqigut6eQCEKFjtR2GUdKJ/xbsId4pizehDEIRML6Kkrtx
W9F2vDad7vGVqKN46ACIpNubJDY6aHwmQHNoKlmXGxsPm8ZBbaquUpDbkOCk
wGQQd4ulHfkb2txI7XH0PM83ZEOUHCtM5OakTlTzCgl2e4ktoELjKFNrR0W5
Afw1COC58ECG4NjQppCdE6F+0mjNTNJ3JVxjIQMzFO9VeLna6jeb7fgp2pJu
mzY6mnlZLGGmyYDdKlPXqtJDE2Qv1udGwqUCvvkogq0RysEjTB66EqZqGqUE
NFA18LCHSIV9XptSVfnYjh/EgKXuk9AYMFAqvA7crb/SxpdBS3blR4rtYxIj
Uema8Rg/wu65slC71/Y1Oh0LKs8z3NdZqx9XCBwy2SETZ1M9tV/ABRq7SEv9
7a1p7C9SxAF7FTJixgfYbz7xT2tYeqvb2T54gT/yvcEEMgmYhA3P6sOr7MFI
sod1fTY5niLL3pOiSNp/+dialfonVnyQ5vT37/IiWEV6lf7E6dvKUgTxZB+3
MkqsFs1J9TGWtcqgAd3ukrrF9X8jfN+6NoKbE2lBfyn5e7O8tVRiKV3O1eHt
ImsFGULQ9fLSbcVATME5EuXURhlJ/BO0ZUoP0Ruy2YgiCi7P48+s5/hvSCFh
IMm0lWpCSngwHWdJC0DkLGE0OYGa9JGLwsJ75oj5n2mICmmKXH1ahDd65sY5
7fXeufJdpSZWXlcV9ERdXhxXrzjcOYG+Let4oTyGuQSmWfP0uxsa+SWvNWU8
Ec+HKXKCv4FmxRDaWSwLvWDr+DGlgXvftXDsuT79HEoIbrGXHc0GXYNOIBY1
iGs1x2YpIMzSl3hd4KEIdTHqXSzsf9J1GgPMP2YX/cThMwkIQ0x/PzveksF0
jIMW+zfVfDWIiavFxVg9RomNsb5WRqE/HDgmWDR4+wYUkJTiUfWQ5Z18FlXg
1VMPrL72ompX46B85kKAsweduqgTASNZPmXO8QoWAXoAaOVQ3RHzPMr0Oyu+
ua6rZbK8ecgn9dxsP++51xQr8rbZN2R4RO4yvINkgDSe6TxXu0Nt0cKhLL3R
8+yWFd3GfZUZPTonxE3a/SNkJD0tM9eoYArHIYzK5xgr6iA9QGb6hxx+QguX
yC0hVX2Gl7uWZ8s5CT4x4DSQridVdeJ0EDsBEI3PZI56JEdEml8tFkiD23lX
LFML2TISuQw994gpjTmD410KselEnv9tEgldW1zs8iTy7dLvGpowwLVH+BAU
/FRJzQznNAcDNOGH6FmggLG2vW0iRaiBgFr0knstX5iH+ZA1KN04k5cRp/BQ
ZJJqD9SSg2NMY6IimHy7/jTJenc5XzDaG0FkPk1oNydrgUX/ioIUqlJBjrDY
DcPP24X3+cZzRvgEGonsmw/4+RvfL17OJ3P74ue8Bbd5hbhUjG/7GqaQ8Vv0
++fojIxKQv5EWlrjRWJ4Vrf/JeQr6WlzPFYrvvUx5ax+h8+L1lwweGSE9jN/
7VuCPwtvFVLZdHaAvvnxsMb7U4DnWRbgcV87AUKvjrQVu69Cjd1V2ATK0E8/
nkm3Nh/quWJHUGW1TS5s9ppL/w+7a51A1SHKI5SswHYOtVsdICuUwb6z2bTo
u6deeVH7aMtmZzIYg7rK/mlNlyFUtWyg1hpubsUyxH5YuQQR3KUiP+dmbcIk
2lFi5YJC/MbP+K0SBljzFATb+S4EtVFdWdWYzefu/lb/FBYc3WtSQ2uwzo2l
mlesHEl/cmzDNwASUJQ/0w6ouxDAO61IxLBVbSZnkLzNw7XJdgPvwWI/H31v
QmV55W4oXVu0urUYu8teQ5HqGj2qzDAGknT8d0deUPyFkE7RViXgB47uMBaB
zP1L6sWEoNw3xdrHa00bv4qotNaM3pyW6SM6v9Td3JMH4vWXB9uoSTVf3uUU
a/FYYa/YgakxCJovdnaA5syGX4/mTwz3AOKM1i5n9XMrwfpYRTZk4TO8jpMi
7PEFZBS6zNlbGPsNPXNrUVCv1h2JZilF/4QrHsI72a4bZVJZs+cgvqtEfXq6
PzcQT3vITyS4q71xLUUiI5JLRby1s3N0gEqk6pf/7/SfPSj81NJHHTwbOCFj
hKCLTziuF7QMfOYsQkhkVQLq7yh19JshTRR3ac2U6f5dV4QVyqe4ke/cNbvq
It9O9+YAa5kwEMZeDyzyqrmPVASjB41ImeFeC8v8QnlS/EYTi+c00qZYLM/P
xMSbBbbR1i82F9b6Isv33GXTB/ByR+TxjyhMmG4dSeH9IANFg+re8ZEc7XrZ
4aQjn7l7l77vaks8SKGJ6NRzHJR43XwkkVXZfUAl+x0jAkxZc7kodD22wSmO
hCaChJ7e2wGoG82R0Ntk/qZnPgqgj49B9/xtYHvo7/bU/cAkZWg1oyq1gTM1
89ltLjFy1RvuHwgRjsS+FlUs8yL62NOCl6PdxHcIOz6VbGFW/I3sC5DHVfCL
CHeIxI5+D/A7o3USXcJLr+ClpyaeF32U/CsmFtH+8DI8OPExQch7F9kbmTSh
cJSZxhtsIDR6fbjJiTdiojlN/uQsC0Te72yVfwmz/+A8XsjUv+5r8SMbH+Cq
1Y+jfwFRdM7pY3mXoyCe4Cpbwgza4k8BAqqVcRI6TgfNTcpTMZPxLVWdK2kF
i/PHC4VtxCiKa9RuGEfNyS7xg7vodv/4khmujkxqeTcLdYkHORy4txhaHZSg
DNhIyAtST23lnWExOaeBJhHxK/205iHLRSUvB2hirzeS7zW2MRU3gdhwyCe/
awqb3gcfEo8YmGl9bRfRakZ4dUwNsNGDyrB/5SEx/ouq+8nBksGikemkQ2YP
4guW8BeUWa87fH9Jq6MyPcMDN1qilDoeb2/BD4gGoyGWQTmH8Gq3H+pUm6Ew
BfxgP0NgfEQ4CmvRlekasn7TKXDzf3RzuC0dCyXpRGOW514Hmayx5t3mFjON
bzUV+QVG7iKCwjmfL5VBhKuZEwn6IyA3I0P6j5DD1HX14YzU9xwv2+h0Rk3o
FsRYoKXauXmMkK/TYuQjgjQbP3BPO/EKtrMPAyXQOZAUEZGzz6yxk4p75+fE
lZScOD22DlyKfyk/Gh156YnLj+6WERC6Jet5OZhlAmkpOyM3fSp7HqMV/A2J
XiGafRGbohOuCu0rNc9d8MHcdikvUS9KggZnVXsVxCPTIZnFeGLT5nFSJ9A4
IRVd/NL0JOQnd3kpppgmZdMMoQW8gcGzQbaMyF5Q7jyI/+sQcTsFK6mldTVE
NxQtV9tEq85gHCb3O1n9P1z1mO/amy2kjdLnNHfe1So2yrgid4A16ivF2vr0
g7he5Imz3hbT9OExvEjd2DiMTJOAezCMAX76jls0Q3IunVVE5sX/CtFX4SMZ
61wLzLvqbONqKVtiSI+5i1k2OYHuzsmFyHDaSNPKW/s3VbkYykSa6cj/N9fg
WPuZoz1N0i4mfCMI/JV36JeHtNb4fdj3JTarUWZasDILc6FSswcwi5vj0I5o
gL+e+kPic/YXkWuWO0wh85Ag1D9vfPFs66EaDJrGLem2/CysHNA13VfKdYTJ
KTXMB1MAIGkWROu8+PjGah7nznCSKPpB9GvWTaOQ0QwYnimfoGzkB0xBphGo
yhkMHFWn7wBJYTglIgOXIaFLZUpe+jGXARDKwxRF/ghwnXuL9nFyuVwIFjOf
HHItnbhtwNKVINcFtRtTmhP8TvsYjvSBpp37XtF6IFee3TXhE7G/RX8p0umR
ZdZh4rHm7j7N9+gjp3edQzNUGFbmwnExFV0YrAMJ0aOC+1me8qC4g2D5HNsC
ADZJvc+/HOoTCyfgg4NKgoneLsIyedls6WDYtHqvGWzxetzWD9RC1bA9UkNz
UPtS6+r3yBrDdtTo/qDVDNTauC+fBlYwh+i6dnCzQEjQCtUSwGUV/bDOCcOD
OV65H8ZocfBANmmPXkL2mQQAKgme7As5jn1Z8plpp1i7eC3WhjOedpDuRIm6
DR+IjBvBS+syaKYEAzcDRhVHM6/q/F7lC7cj2qmAveHP5+lDN+M11qhZQSB+
+vrjURLsg7Eg5fnphc4XY0DLCXj17+V6tacKPrudXiv224S+leu8h962tI+k
E0nFWuTkf1q9nObpkjsypUwKDbDhrPdEkRcDXrQuardmldiqCWXB0RD8kvDt
8eEC7iSK2rgUEir+KO32MdOlI8iETnt8ztxfJkkrELbFd5ifoAdIIonpjw0o
DV7+IVXnUCQ5iEX2MVtcgQYz4dbzojP1iFx35Sp96A9dHYe/tly/rQX0iegy
6Wjrt3bdngDbY1alA/o/Qpouk+t0Vcgr6rJY2fDrUNo4XSyJOPdzuP8HEpwW
AqW2xxW9lbETiPCeYGVLtzPl5HVc6M0r8UW5rw4xByJPSnIKyr+LfixUwLdJ
J1k2oKjmErJ1bkaOSvpqyUrhZ2vGiyOczNI8xYOSx49GEF7KyzTtMmqYZId+
wd6/d8KJi2gOEwOm6rlIU0GxPG/p45JkWRnuFXcKPRFQkKAVJ4BUIycxjK3S
cgTqVJWJt8tdNzPy0nbnCtvXhFS29xnjQRDLPa57R31AVcZZ2lNn8/ys3BA6
XJmhV/kiJ3x7GjvlVT+6M9S9OvRrHYQc6mKP4ya/sCup4AxMy7NNuZFPNsvF
ZNz15pQ2LqN3m8dN8B9oK8sbHV5oVciR1b8+qFSAyk2EADVqG1IczN7MtOkA
fMG6OF0PqYVUTBWbosHHXoHFM2ypZKZ88gTikhdu7ooaIQ+P9HHWkiAOCOoJ
81DiK0DGoPSl6AhxJOp47CW9i9wtQMSaB7IizIGzUf8RzbnRixpmqVLSpdpR
BJOuMyKfYCNRuorhr9UrXGiGkOhRAseHt/jsWX5TqMG3XLZlfkmf7NesdG3p
BlomJIP8tVBDryxfcms69GsEbzAKrFpCgheH0lGbIN+/rHWWJoyfCGuoozoB
LfRfGhkK8NLY0YrOhN8KDTJE0BgmkXbjrK1GTBqfdrnBQh/uuccyj21edwIw
G8PbHvRRY+vtrG6RUeoU8A1ZaC4aasKfr8KUmp09tpELYo0yDKh00om5dL+J
vRnsqemcbWbKkQW2SL957194N/Q6QuSV99oKf/ci29tKLsXb/A9QZmRMQEhp
vQiR5NhDruibJH4L2orBB+GmIXsOjNTr3dglEoOXHQ0/y4QHYHGixZUf8tKa
anBIfV++SesUux8o1b+DRMnmUl9nKJPBLmEtWHPNUrUoXh/PBjCmuWIIb+rA
CuIq4QZhTdcADvBjBBurCQl1XY/cCQhRSy+h+ICfQPLIC06hQSkyz9nvWuCi
EijTbVBbuFK/Zsr5KtZCKsQtQlJ7jlcAtk7BTZKE98mLkSW9tHj/LH9quTOQ
aANoIEJRfp9T6dsJJj4M0hnR1STUbrqHqjSCNVqWlpmWtNuHRD1STEsOg6Ld
hnKz58CgeRwN1OunlZpT57QaAtElSj99tIfoybIDxWViqTO6k1GIawu/g+Gb
HV8P7sZOgIU/nIghM+hlwXjUx8wHnWXeZ/bktWdfYCkrE2M/X8V9mk54a5Qb
cDUhJWXqTNAWgV6B+YodIPb5xs9NuoV6MSzGvkKed/r5SKWc4dz0TwsHRI7i
g0hLpqVz7eE2dFQbXJCkpLe+FkGGFPAITnsopP5uxu6Q4z8kX130nkiXdFIm
bWO6wLdMMV5uop+3BBCvFaiK0Q6JVoJTysFoQeFifjbj1+UJ3FsZMqtT2b4M
kMmPIpyZdkfaPOPWTs0KwNJPJxx0hPZEt46DU5XKkgw23ES8mF8C8JufBMHc
7ybI7qAGmPWietAHufl+U5pHXatZMsGoh1SVso+uP77YiW2wxPAqvAjtN9I2
NfXMk1B5zyjV1dlL7GVZ6rxQS/99/F5q4b6kThz43ruFPvDW2TIcZn8yAOdk
FqBukVE1LqK6D4Ftz02rGVnlhwdfDalON//2PqMZYdwpTRMvbcCjHoDl6zkd
JeYjNYkEnYWv4gtip77foCw215hpkBYwBBZVFrwBXpmpeXz3WbjJdNxTRAFQ
Y3ZkTtrhjcSDNdLAb/A1PY3kaeMzQxIMo0lQv4yO2SWkhoOVkt0JLWDn4wN+
FecYAph2F4JV0flIbOqZlIUmCVC4CtDimjTcXbF0Hzf6w0WufYfiUd0uiHS1
GzXBA6EdFeDQvvKGs/0ACUOUU3N+wwL39Xkyg8q6FY8fFRAbwbF/CfMy4Ztu
0D464KUqy5T9cyRKyOLW4BdFB1vQpZOWnu9+xyOzrx5AlnbTQAXa7MY2tykG
9U6HkcFSiKWXk4aafqGr4HGGiI+fFhxCtk/iEFcs7o3n7BcWUzm/So7UTdJX
1kXXHgKK9JORiekHxmy8ldZti3giRLia7hdCIs0WjFz7R3mtGOs8na1mTQjC
AQH5qaxQI3CYh3EZSZvJE01R6oGE8ya0zXlJ6NULaNy1bHP7VMizOyHTSOMI
byuMvFXCYmef4VSsFTD1pMsqjReWAq4PgjKZMlb+f4uXUZuBjapWbMluuqKB
6ZS5dDq3g3BLUSbLQC7pe76/ZLtCxc25SMeYXM2uSHUAL4u5VR2RA9n6invD
uE/ynSftEnv8TDYu6iRI5VZR+bF41iZyuk/MG+F7z84cf3n5tQcr+tBcavN7
MEfA5WwMITjxPhbtrCpNDK9ZAcmBUBqQmlTkd9XQOlQ1mzFMcthdWrLpWc5C
qmUH6ldeLleiD06lATszsJJS4nImfhWrGIBB7NdMhFArRtHO+5GjJfwdLjEj
Us4OQjd905V1zANcyE7928b3QM3oF/LS405bemzwku4Pm3qQhoRp7irgtxf4
THnJHVzmSQZ8i2hR5KmnFjREdLQCDAM654oOuZsgKO7509rB9M3chf/fAmIS
U9poFcxnRfD7OX+3Yqg4DUiluyvzAy5UN+S1/EGMWEto3jBSEIyVR8sj4Ewg
0LyoGX65aczD9VlVJv7hIo+9VWCi7+VbTHRk47KLjt32l9y/lD31GMeD3jIt
5NFUP/RYJtZ4gY/QJ3daX1nOF5mlM13LKdpRFONbkJtBOob5ZevkSuiC0/D6
gjoe+L62wf8CiwBsAJmUd7fnNLGky+8jWiNqd2T+JzclX9HzPYWFFsdrCKG+
hIwCppssL1B/lICQDiwKVlSL8NaaSuQs2m9Ged1bE27x37QVFLbzzMUec4LJ
wEuSk792zJ7vjquoHro0r6I57WYAzBgw0i+u6ELEQ2kVjY1lgPocgqAqsWhd
QUs0nxMDmUOk4GhUnFgyA8WaC/jy8iolx6FBQ1Pj6gpJj6FTEbInOKexsU3w
bY7/7dhaXAZ+tq/hflNyEvLg1iJJ3aummj2F0ln7/nSv0fYxZ3wfq7JosTwc
q9j/70UMTjl/gcRENr413Jczsi6x465fRYdPNpZtpybV6tbZ7V4KjwZFcViI
Buef2qr9OhKTXGXzW/9whg1k2FeCEg91fD/YWgpiWgkqZZIMkusrvg6RPVCi
gFSO/gu+ADLCqo3CYbqWqpbPuzThuijLXuyZ1yBl5aWSIbZ3YYMZe81QUvN2
CSVktGFNZpO2qFQJlyhei/HrvXlL4wX5NDtirrEj3fcz1ey5kXSE71QlYpIL
g1i7qtq4fdR3I4UB0yS2ReQgyKplKPkDJzH7sRdv2VTkWJ1g5zNh5B68wCsK
4nxkqjXIovkb4hqzaU7b9YlJ3Tp0cQSB6D0YFDcDpX1qh+jvh5xH8laFBeky
O5z6uQGqe8TmdFSG0uR9T1BoCnFRe5EYq0g7Ix6ZBQNNdLIdr9zDfaCxS1Yl
zT8ua4cMYRiIJnDNbb6PLfWYImc0aej5voAtgeof9c3zXRqG+MxGPCaDJyOw
T46sRk7oQ+eWSvqE83ojMT1FYk1PhbUB12wpSrD8Z0A2vqmr8RLdWYPy3ru6
3+PZapN6rm1uyM1UFed3MtuOEai2lbpo3dVn2/wWlVGexvWmhkE9U93TYEzc
92SpHeZBh/hTteMmKDU4HTyFA6TigFpqYP+e90FTpc4MlyibcOaHBmUGQDOm
yLtlx1i8uydDsVqIkRTczylWLjf+YpuQcGNi5qfAKofHVSG9jYqtxPKBORkd
TXi/LRjnVIXPR2JsUncvWlZE6JDgebvA+zw6XnCJMGBw1K+gPsz17BDz6e8a
m2sjyFZ5HQQblk83BJaOupGDalox3lfvpMy9KhsF7aligSA8s+RvxnbiQLz8
Dly34SEFdRRQ2wneFiiPz96zf5QaxjDZUAoe+eu6kIsy2GFwaNQg13piRNef
j7MaOJv6nrHy46/13/U0zKyz4pHWofyY30ESGhslX6Z/5DhiBUxmS3GZ/z/6
i+AFo6RV+3CW9Z85XyXUbjGV3K1Il3qrfCu+F0PQngjlzL0kRO/S8kvchOjd
TigKm0OcgCySRDgPijp/TqQYM+rdyma6ZC6U/DhaOTz9f3d8CXriGIqf8ZCE
p0oXxLmgN/lNtWCdN8AFP9mdZoGOgGFIDVhR533oX+VnUSUbYeDouOYb6bLg
AlG4D0ycXqLW0aZeJh5YoOWPfeD/hiRThOWlYj/XAZsIGbWV4pOtddJYN+BP
XZcBuT3eSodOJ6H22fnVKM6DD2n3dclOOVxtK+isTdCwJ+dhf51jYG+9Ewex
Gy+TS6UjwBrCK6aL60gicY8zA+G1ZX8y4O0D+wk429WWZ+Ww33FTRDpGBFyJ
bpK47ekoheWDsg6bR42sug9+ig4z+ZMYVOW+9XIAbCcP63bvxS2ggzwB7Wi8
2RYC6dQnujkcNIZKv098I5uiXrzzc6849Dn1zWCvZ0DOIe5rDZvdXR0nyQjo
ZOqoQvNosO/GHyjfHjvYCIpxYGE8OIibFZG+0FilAS3WUx81PGC1wrfSadw/
TQi+1Tw3b4n8J+LqOsAn1gYx+OQutkLEc8HdGTQ6uRmhuPHkakQyqj4tkvVz
IMkBpzy6teT5XYbaLNxG6T8rJRO2brFDQ7kLt4DKesakOuP8/j4snQA02Weh
tWhwktPhg45ZCV+H4/WG0KKXaWMQbpL1iWzzy0n1EwKIHVCxxiw5dIqyfjn0
antkcFG0M6A3Smfcg4c1FheSpT/q1KfGjqFDn/kWMOybaG7YT/90lowMWczN
io3ANPskreOTYVBr7QxiZ8+pZGLjq97b3SNNsroyTizE28P+Cnk8G3dooORz
F21XcwSaGyp/dCzETS0sWa1LPu3gDzcQIf49eNwHZ6KNjWYvnlLOPz2Z6b/k
vQyyRGebo/s2LHnP/MGkJu6P2NiNbtWRxv0bp26VatMi5vxw8OangWnsu7HP
sFUQ445/NSE4S+Tr246+Ss3Sr91nEuWymabai5v5rGd69KM5z92++T0wUBPM
EVkyrl3zVCOmHwjzBQ7T8OkvDXSGpR/JWIetWqA4oLxzfjR9p29AvFMSLEKz
p6Ercq+2I8IdHD4nU9X61bbiOHhNkHA1mJLFmsCryb17TLB1sh/Om/9f6IMn
Ip7h9oMpniUNGYImCKR11U8OptuI3TlXx6YvmmPV7Zs5e7wJM/l+RLUGv+W8
ZsmKDHT8UgnZ7LUx5T/ZEY95rFbAbyrp1FeLCpwuTxK3qVGqlU+qEP/8Frpw
X8E9RtXckKadkGGem1wSPcKnbvk9ssC6Iv3lV7ltBCBYmsp2mc0OWWn1Jryy
QUav40GcwsLRhvSpdYr7VWBhB9koc1ky3cp8j/56lPui5rTJAYcRmiTsZ1aw
rrd9EkQZZta55aacfFWHR1WOrKmkAmBBh3LAxptsZn6MxJxMU4nW8e1HRdB5
gfd5wsfAkqQSkzNWQ7gbAxfrj2M+1NQKQWilG0oPebUy+wff9cpHtjX7+5B3
vK3/+k8gewfes+3TWUwKvH//KCc7U+v9bLs3YWz28kUqqwAV7fKlSRJG3L9o
6XF34g/YoaImSbXN6Z/uDkart7rfr/Flq09K4fdNRKtr8r2Kg8JVY//dS44R
+diy3fGxrWnzvdXOckbeYqbUiSYdS7VBOHRGTb8i3Mm+kPKYqDlrxCN4UFfN
5hgYy8HyFIMMvaTA9rASs3pQ8LiF7EevalBuDDn1l1k7ba6PAJqGFZ3Ams/0
Y/SKQrSfrMNX4YFsywMHk9HW7bVZFDejv03CatYxV7OsP/2P7TQ/bQ3Lk81C
3lFja56jBrpx6GmjkazKOL6YNkQiVLpuojXnx9oFyiwN8xVTbWwpzEDNshyH
syeR6CGhvrSZ6a3SQM24z98K5UPlMHnv/6gq1VUxPRXkY32Sw+jnwm20Gtn8
Tnaa9e6bZypK+zHhKWO0zCuUjIXtaPdkN5V4XmgvFIl5hCxLEzLHj8Jg5jlb
OmPSzQW8f5ApHi11G0m2UCZNPFM7xa0EXJHY6nUf9lAORXRlakmH54Uro6YG
dxZf5nrFFjZRkUk7Gh1wSnogHOYSDkT+gYO3IYyN1ZQRJQGN+w117H6fhlNt
q0HABHkWl83eDTnxkMHjrLJlf1/eA8iA+v7mq3MjM4D27tQ5QJzHTCo097wd
kGjLvxFBREM18RX5MNSmEVFg1w9cfGU3nl5VSuYsC2aRopJIScX7c/A8mp6+
sEzBx790OakVP/4fERlMaqzjZXWq6rB6a7ezX9AMgjYjrImQEfrOLEhPrr3P
yWNUAe59f7wquHagJaLDYaRapq8IxoEdBZw8E5YesFOCK9SHK38Z0cGo1Bpz
FHir6e3bGp0ysQnsKIXECNsLWKyZhrwpvn0ZmUiwJhGtAqtowXf96TyT/o+a
+w1ezimtE2m6zweEl4tzwdzzFWCkZh540WMU4EK/Zgz2vKb2QLUIFJaSdDSw
Kr13209f+XUohHomKVW1wPqBgHiib/7LFYituNMAuygXSXiOwp1VfLLoKX7i
A7qmc4Ys10fbf4Pho6ZUT/WHLxyj0xUvAaN8976uyapLYqdG4ccU4R1RJyvO
XH2J3w1B24YcCFK83R3oyp1z8bklUWQ6hJhVsbxXeiKdULLRV+VRnfE57oqh
AglGjbryA3J6HBhSHsTQ1mc5LFyNEih9SziX1Zs/qUcMrC+F7iKXysVi3MoA
KsQD5OW6HKLsqJCvAdysK2PgYcaSsaysufeKh5L/06PoIHp8sb9Qo00md7mN
AO5MxgDVCTfx2ABRnAH91S0FNXUZk4i1UDPWwb+sQRWcRmi3uQxQ1ZWYecZj
uGUiI3QHdcJC3hQS6tePb0nOn+8gRNGyFEljrQNk5vOg07oS6u2708YQ12fK
Pwk/eO+jTx2BWUVggTOtaK64XIQnjTXG3i23DHAlvPtlNvbBx0zQkfUC6Ki+
aPDvQpBhmoDAiQn1JyB772S4Rew3Bkw3MAzGQemwDbqRpJ0q5GVpOUYEAbo4
oQxgG76D/49uXAzixVcrsFEst9OrlStX3+BZqphg1ghexbuKf/M+A1e9IMlg
fH1JGiowEiXt5ttGgrgOQsBIhTxFAZsRqMy5VjMytNoE5LvT5JGKXFBc7NT6
+H/NJft4Wbbiz0+XFvMpzmkop7Vj3ytsaZKMXbYgT07XA7LQuZS2uzUyL+Ik
7RrEy0ChWkM2totxMFBKHChB6YrQXsN67FoCXOCWDftRkwFkgvw19GMY5YyM
bDTLFFsdJaD6cqKNtczdOO7BbbNJA9Crn8Tcs9iIFFiZtNoa7eWXGidCSqBe
pmw+ipYHHOuOajA3k6bqMa25HHyx6wy0YCwAfn55fh2tl5n65Whrl0X2RKqP
vgrbQrglFdszBLxDtvtmD3RNBrWfisp8rdvHp4HRhsjrc6cyZuL6oVxaEFdb
RuOKvOJ1tLnPnatP+TIXL/Ba3Myqm38JC2dZV4R/JsDoJ4uoJ5ANGYJwGH+X
RKqHgUKFrmgLs6sO4wKNPFSAbS8vnDgLnIfB2OoBDf/jsrsBHIs1A5hAN3Vi
KsLWdkmtK6dro8KeltSBIGjoqyGuOp07LHPF4Sbr1eOthZwGvAZ/o5lchfIe
jZjnhQj5p5K4R4rONliThWUVSkfP8wh+vsAZQuV7YzB5V7hF42509oIx65RA
mWpD7miP6hw3n8yR+j2/8zHpZ8wVNR5/F5myC7cagnolHxdBPgkx0PzWmfyh
fsQSfPtpCSxsvIw1KjyGUF/ZJ2TNGy/eOGq+9/qhNR7AhArNjvWlV+ozJiAR
cVG+NMxoRCg4+G/m+oARJHdE3WiIqhrK0xYPVOlThODiuIiqrT9EhSy/DkeN
ld38dbtgW7WqDZaPbkwQ/hArvuMWDd/wVOl6ORyw7X2i0tNpDemwv1ZC8Iwp
CUK/ZWJnTHIozYNUlnZgfz+wWzk2ebYGVBWmEpOxIqOF1PMpPltH8JTJlotz
USdZ7FabI31nBeqn3DlfvaVss6bN/WKu7pqqTySSXz0i9QsVTHIFryAoUlYg
xrCxbaLU0aRha9jH/Qq+bGrBcT24B0ztM/Ez52szfYncjSGCBcrIOQ/wghOc
t0GEmxVkEVL+jPUlwWBCjwd7gRSh05aLCqSFVWGU3hR7EXFrljVNcatZMhKZ
71as945m9lstIe0J3ETpaCV7KeGto3TEN06F4+7ztX2fu8s7Ae/zIsRojxsS
GXFa1iTzC1tbB392I3P51z6XcYMjmLnoGJz/C4snivouB7yorOIeFNF/m+gE
bjDWuBlb2BW/SvnB/nKYcvn8kwM6mxBdy9WiPeBqqp8p5txWT3oVK3SFvq4z
DUABEDwIESTA7/x7Bcyxz3wXCoPWCnw5iPpjGMgcoUl+xNWuVwCq7TCC5qVp
2bWcORvHLStjuOi7/x2Wk7VEYJcsFFajwEROlVuirxA4JB9Hov2J6P1SgOjY
ejOfqWtnmlRdsU+4U615TWbFKFjUN1BGbx1YhaJ7uAuZPJjHr4o+rqGyyIMF
4xNIYpmGawjo2kdjX7j1nIriDM/DFVHHSQIfQJDsog+qE3/+pa+QuxEe0eHb
1Folr89XEKXYOIDUEtyuEsEq+Vn/Y1o+xj8bZyyHjv4qOBwLXCabfaajLXxR
4/fPb//Ky4AZjJUGvaLEw7bbV8Xu/CEggWzgFxC4jC2xUpS4CUjo1UCoCzCq
olszb3cxwYBeECGmbQHqcunnn/6/fDndT8DKXmTPrIuCNzqc1JZuGSkIqDpD
VI9F0I4LsgZqm+IPOs/lpiuDqBUhAGxZlf+cZp49lcJkr1wAnK8eHFMejs5o
fOXppJl16gw+XFD3o5wiYm8qT1+pKPOXNHFXiYh9KbjQRgzBVxQGbnC4yvaY
50Dllr3bIZkH+rKW+m/TbVYFdIHGKLG3rHonbV9rH2f8L4yC5UjJ52ENE7zr
3rM6hyi9GFCNcA4SX2dCc2+ETSPoPjjBaf8q7lGBrGOhX1iKy9daD2ifnNCT
Waf2dBfE6WTkq0tabnExalcQZ9rP3f6TzN8p8o37+T8KxEGj3KO4YWdjqaaN
t7vdVGoXiuRtVk9NvvfSiFJgAcjX8LUPk98wHx4lkInNkKhN4IHUSOCtFGeM
An/AGfCUNWNxIZIG6C0BSpQPL4OWTSHEAdV5JEVQ35vPqP21YC+29gb+HnLx
NQfSls7Q7YiVNdm/lTSBJwM5QRUtBfQ+XZ3FZ1eBfKtlRWNMJzJorkokYlC3
S+ebV8+nCuYqszhTJlrN21Zl6zo3slk+7KWC/uiq43dPpZCeVQEb/HU8jZMN
UDc5JSA/t9ea+XgFUfO07kgAZhU4xxBPSGHKVQwhjPH8qGiLVCFYYpM8EIAq
USxTzChITr52cA0gYKbYOKpL0CXsNWqH1JN7UfJJ+HbRTkOv8kfd1Lla3MMg
Vvo8C9L0oLBg05hwN/RI36rIR6SwNN2MClxveVlYfQvLKG3KK9K3489BiPYF
DtlQxHt2qJ4EyxIrrQ73T45wfzqTzRKEUc52C6DlwIiTohrpnoPONmQVioT0
+mLeID3QilmVmb1nPFGO4SaBQOVtz5TqztusO6dSq6f7qDe6WR1y8DXw3yo2
CU0TE0stOTibv5n5ROZw19H6SakNvyzrj+v9nDe5dQKvjMSUl1/cVS69TCMg
0xDD6v0s5/jSL83pAEcT+f37TexoYDNwfjWHZqf2mzLM46iB7YdPIPXh5c+z
/pY6nRsyP0yU7nLaCe/cg7I6OQ3fiZkuGdaZlGwm/uPxLzHY8Q8/IBXhs+h9
5yfByMiN7W/yeQIZlfW6s3ZaFfAHYgh4W9zATc/BPMqSmVOlwBV4KTh8z6lA
BmtPuneZGhoMmynAAJQOIjQMUZT07IGpp6GKA3s7Yx829AU7xzdBWbT46jfq
k4EhUOfCYzvfG1IDtp6KLR0OHTA3W+dJPZZlgSU7Y4dOQqpDWFY91on47yKj
eyVXHtKHYkwhibW87crePxw1EQJENv79kyXKg/uYhT3KU8NAt27oZrWzb+uu
QM9m0uiR1Mp5UemRrNef3v6j8xzp35gofGRGyEem9Dyy5OIR9eI0Q9RDoQ6M
wV1F3ZVdI7tyn8i0uDlTZyic7JjIIP/XaM6IN8H5KxoH7cRYuArtjI8JCF3Q
j10vSuBJl2oUIq8A+KP01KTDsiVG9j9z1Lw9haIFJ4wzctjF2aggdU1Xgw4X
/SE+hiEv4L+lXk4bH2YTEFvDP+eVR1PqcoEW+gwKw5fEEE9XT+JeV3HC0DA5
on4ZmQjmIOjanR3Q6hgqJbQizXE3gi6q1hZHDrBja3CIF/EGKeo2w9n6XajU
NJNoen2XLO0nJAQ2vtNS9Jh8e9MRF96nH6WQbtslWHkisyaOyiHe5au5dlnE
xvLSN2zZn6C10zTeLPfQ3h93s6ibmDUpqjfcrBciySALFxlgVm1b4iuW+Hpn
+wpdBKQqSSiAi1AtUloDjRK5Sky4XoCnVtww49eX6RpcFY0vu/4WcyJoZcVO
5vSfcU65RMiyy9pUw4975t6/k8eM3yZ81BNM0KIrGfplrmL9HHzsXF4BZHWy
33UVJ4kQb91RHNrrb8jmFjX+UPTkrsauXdiq2ibovA/WMCK7Pl9N/DUI+vF9
XjyaIIu/uCmsB3hs7bDaL/5pdZeRdXl5zb2R57PBHwq4mSMy7Id7Woo+kDHV
FyJwWKe+ViU5kqhT2FaaEz9hf1Zot/HOk9X1YjhZfn5gXqEGMIqLHPGvXgqF
9LiBzJaJR4OeEVVinBBSYh5I5SqoxQ2i4r148hb6GJe5B0oegGpWBJoQSPDV
WAiHVeYqk6ZKPxe+awBRpezw4AxVz5PyN84jdqi/F40j2FkCshJfoNAp/Vtc
CrfGhBaVgh2d99g+xAaVptEAGFoGiB3tPzSCZbQfZE5nOwQjErIf2JxEsZoU
3SGZdOb/o+v7Ko2PCtg9JB0NQxTNSSmEXDNOg11+IL4ZjJTY5C0hXnmi1zGN
bl3Gp1tre7bxE8bPW5qeog6vbbboPM2Juhbgt03GX/BoZmybWhD5c1K31afT
glBoMjTt3YIWLnsNTTaGKZcGaT+c6zJGYKkAjGwZsbprmAvatLKsIP2Y/8Sc
bDpqNCPQdn1HgUZhHEayWOkGrg/8T4xorRqkkwHAgaEKCNQNu5E+m4a1dGSy
NM5MbeH+wcHMEEafhdG1f+MImRTRwwSDvWTG4E4Xgb2KuAzHrP3NRIaEka+O
QnZuZzw6VO2ZomGIkupstlg+TmP43Ai8Gzov8QQj0o0LbmTD0aQ+ujpUeZsW
KdgLx6FDurRteTO8vmH8gdLJLrRTxCgWyUgMS2Ss7GadVKephZ9lEFjM/OLr
jX83c7V0QKit7N6jKcmUOjKvYOHvvS25vI05GW6ARxn4Fd1ENPzoNHeqigJ8
KJB4exqP2C0Ut9YKdDvODjE99IiWHVhYZEJ5KlvVx6loYTyYnQtiGnZyCy4+
5//DnkYyXyE10UHlSOyaYAg2Or3IhDWXwIuAnjrh7SdOjNbUgiVrgFWAMjlM
qy4hCw/+IU365Nzkx8vUaaol4Sn+AluD/m2/ke0ai/bJFsaFO5iWISJ+lPzf
QrtesUEms5l2z59v8GtdLxMhNJ0WpSiptlm0E6JC84etUFSy+rE8WPx/vtRw
2f+0kIohrhn1fbweIfppx4dGz9BeZfY8qj8e1JsuhnECXn1+v6WpnRyzkMx6
A8mY+iwPVs5kiwIBq4KKOTb51NfCZlaUGzfZ5o/oD1UYZrKYfpZc/loYPJNU
PxFOM9Cgu2wuseA9+yWzUp4+oaeUaq8eV3oOLOQ9/BHnRGLBs4C2SMiFs7k8
/x4ekVpto8jH0G6pjYmWeMz3dT39pFycyKxqmYCNWC7XTP7UZeTsswMucuco
V0OO+GpHMtF9WkSQwr7ldUhXimC+6KVcEkaafZYgtDYav6Dmx/oX/3xzReCS
LV/nJgkn5fmeVsmeCQhL5NMi6Zyi0YnacDEfsAsiRgH/IpsYHY/DnfjkACRR
6cpWuUKzFJcjVIZRPAN9kG3HnSbQfH/zWc/Vgb3seuU2Lo7oYnQIqinbz8SA
mifsTeWdDDu3SZthY5TmhPADcTzLyFwLlVs6f5oNyF+IcGq3+uY+oRRNKFzy
xoFanvh83h+LVoGg0Gs3aSf93t/LVniShd8qwUhwjtTXbsUITsTwO6LFXSbY
Lds3xzDUyyWSOCTW9RmqHqOO8sxuAzsWVB4CqHYX96ICnzoa8nx/BrpHphq3
8trZdg1D234BYZcR0r9tZxU2sJBDLnb9mhEPh3VqJpaCFAAzqJRERXbuJsFu
EVlFItJz+4JarMYAO6RERwkP5V19SDFsPtamclqJqnrXRfZm7TGBSYWWJt9B
FQwY+MA9QYBOd01TNyIexQl3muinmCc9pYDp6pchmL51Hl7yPCd2zzfjtEVF
Mx5Oc8gQ/ukYNTmQVOqWtAnTqcceaQ1m9jO0X988V/cNxiHtpGi/XmyQFBE1
6agmugQKnju3jnFFp8pb8m69FGyOLEyPoQ8TWVx7XM74Cn2ZvRLbI7O1gAaO
Hl19K4BpjiX8Ogg3YDEW0z3/e4Xy+6Dac/e5uYUTEfs6Zv7ilHLXx6loMqRR
seqWDSrcGmyfKK4DQVa/mMNPxQRAPYcc9AeHP7NVupNFrUE59T9O1YD+7+Ro
W6L/vz0NGNezzymPouoz7C0m0fXh9Dee2/adQFt18jO8OiJS/DYE0q5IPlFt
QEnAB5iPM9EvbHwcZTWn20/zNomiK7elenXjTLrOjHNmvLB3lSdyYcfZ0piv
hTPZ2v67fkZQ+lm6chdzYgThtf+e9vyWYjWqVZ1dhUR9veatk+5wsuGFqUxU
6kL4gZzLgWydP8VC+U8Mh+kYyK2WKmxhG3Q2Pi8b2xvPG3HivxJyt1oURuKq
F58ndjgYLRBRKRqDCZE0m1x1yzdbjyMXcYEJ4skLllqVTYTq1L6r0a0kTmcG
Abvk7WNX1qUe7xFj5O+zTTPpU2yUNjF9xHxk2ZCSOrhteF+Mi/OG6VyotuN8
JuVabABCuGb0XveUFtMXXOvGh/fzZzBpUfeOTE1Dm2d+uZ3rIsTODobfmWo2
J5EM4S0Ymk+08pwL/wOdV0024G5uundh6rxBoK6ET5cBvJnitiaQfYmQ+Kdr
lX1+bpd7yZq4MUtVDniQhRzNTqOy4EUjVzqIHteYM2L0YV0f6GSfoZBvL9uB
PdFQ49WPtSs4eRjc99hzIXetwUyD+W49O91chWJ49UG/LOpZfYbhCxW6uf5p
5Y8GDQrb0mvQxcIHKEuHx1hFwFZeeXarbdf4dGnVlDo5XgeXxstR229TKpro
Pvv44KIiRbARKYL9mCBCUAewbV6bmI27MexIug3WYHfhJRIxWjbK8pIMQn1l
S4FCkqGIdb55qCOLAWzDjBTmeXnmx9+Zy+2vnsF7yUurwA7h98CZsvH3DgJO
xxF9rxsPE+vSBB3YVmqOwRyNujL5BXAnxKN9KNWMtCcyuRNM1gMg/0LjIxv1
qozMXgW2euv5oHk0te4FmNwGIyaFNMvuN8igKLTzJo8aIaHficWle36WDdPl
ib40XNi1QsXPX9ksdknDcFiwZpRea5gDk4f35y3a0LAcl1dT7sFm8fRqh7Gs
bgQLselM6ombnmYM/3flfLdA4Zdi7cGPqB6olKIPieMwZVMAiVq44h4tMKCt
BNbtnwTwo7y+EGVxBZjL5qYawU62lAKQ/QWcwm2OuT7pA2ouWdkCPbMNRnSA
34Xdep/3fexTqHx8ymvR+R1L+BeI2436/nmAVcKFREHZ2Znjw4C+Nv4ijOdx
7jIxkwbLd6d3Jw2La1nWUayvkaI3MGhKxjVlhKr3G/j8DClmorxbp/uY06cF
EoYc8bL9uOtwMOtN+U6tQIItPKK1fvqhtjGILf2KGJQ/e0eY4DPls7vko8hS
Mypn5vm7RCYG8fuH4s/StE4vQaOiDUvA6kRGUSLm8B6nbxxs9IgsvY+YcYv3
d3QMQ9tESOn5mOKxGvQwzpP/THneuKb8G9zmUAflGMfjzDlu9HlfWswMYUn/
cH09I0HVbxcNDNicLG9Qz2fKwLq46fWl2cGJoFu/kzLgdj1JIHAYWHRWvOdD
N2+1yOn9ScgDFtQyysTzIsAQrvLxxzJYMq12YiOcUIrgbXNdAVGAKoxszUkV
/kJ7jWnA1Dg+k3q5h24VyRLWztw5tqYlmd6yZ9V3jGpaNyaRv31Mj4gOF/F6
3+Unyj4QTM+OQP7/bYjecb2e+g6LrJnLOref0B2t54/XDoPq3EcpQJpm1uWb
Q13oDvgFJq2FYq6C0G7Pjh9P3xBFF61R0ts3EoZbIpuphXGXUFyEwBnaBk+j
rpi/9kIXFjd8Gs0cY+UzN5vjkBvbZO6u71qmJqB5/bkkkD5CAUsGE40yL6SN
5WBOLcyeCvT5wEr0fwijdsdyvkEay60aUNFphlshJ/TQPbBR3HrXvXYNWz/D
WvAG1/CWtbrjywpPobKASgP29EejJFa/nh9YrkGwWFvJLlWfj4RwOev+fA1M
r6AiKbUy/rsu8Ep8Y+NYC1mTsd2Jh1AW6Qd+9i0cNzpjWoSFMb3tFRB4GpQF
AFwB+MTVbZaHz6PNc/ncYizRGicUhFypU4eyelY6DhOs8vY2Uts+rcPBe1yp
kPV+3BenoVrdrH6YGvcBr1BIOA6vhnGIijVKwbF4OwA2F3nLjAUGwQ756PwC
v+z3msCjLsv5eNEd7uNZVg2KWKWxjQLMUn2vLXMyUvFHTCLbS4rJFteiAAJm
lZ9jprJZIkVg+/JnQfYTdMq0hJ5/z+ok/Z82NBwdJM1NcK9a+3DfPURb0Xyz
H96zRBr8YC/QIGA7w+3WuSQqBzSYlwkK5ZtLvIfskZAZlJr8d7ZObooNRKpL
alIcmp4TaupM4kFd/X8OjobnraUuM3hUcQPSqcare8n/JAbJKZZ9axpsqtZA
9ig+Z+jbPMmGGB512d0c/hJhwAJvhfPHhEy0tnmgLvbcGH/d8SkL5goyp+Rw
uyLi99HmxEKMg9HJIlichredUhbudeTj17Km+RTWKVumz3HcbTMGrcq5R2eJ
LCkJN+qOe+Wf7zYSoukghxiyoD8ANeu5RNssOGS9xlHJ46LlvKXBDDt9WCSA
TRm+W8XbNl2Qujhr3hKMqTrdWh4utePCNEFjFyMyaquENOQ3LECTVz8faQJN
BaOGv6A/aTztSrfaT1ruPerTTMpPy6KuOoQlRBVfwRu4OXhlQoiXHwSKvxI9
dBXuj6o+KVpRz0sYcjLlgxpwGslPOYes6UQ1iJAscJj+UszBsVb9doht3SeY
uocYvBga26lnATdg4Q+AObrwQ9SiZyoqG6RednZsoA9wrhZiH2VIcK5MCVh6
qjYFdjgZPLut3VSfOeC7i1ePFQQ1W3obTId10Ull7KGLR9AJL4ibxoTM2vwS
wzKuyEb//ma4FDoj1F9ZbjH4FR/f3gCMvYQVxldDnbArkxfSxbCzv8eBz2DV
ByHaqvYYG5jSX4yknxIsIeHKB8MQOXX8X0Pp36EEXtQbPVM6AGcs6BoGcnPZ
zCaQ0z8De2S0zqN9J+HXXijJJIly+58E6OQDTU5iNvae3w7sZ1S/A9lD7Bdb
0Wxs02NT7Kg1F8gGhNwKKMCCYylZfjNUqN7tU5jYyMg1Z0Akz/pZDhKxn10d
QFs7lIGyTERbTORBTsZMqtAMCh4KtEGrak3FsAO1z78JmJ754SWf58nCJ28p
oznyg7TqGAvhOjWxeYjOxHjycqERGyjYqktAc4wM1n74hUBYJjhRvOggZeEw
fUipwOIQy0d87bwKle1/dvJnHxabmvsnK5Phdryen6sjiPDaQWbdkCBvquIs
i4xGf6mnpJfChLRHtkEBsrm/lSM9DsSto5egN2zawK2iHTchnFwm9WLzBkdM
ca/hIWnk7qRJCxwCI/vbPlKLRxUYBisarHgpRQtQC7qKTxhvx6BK2h591662
GyKRON0WYIrW00EZuiHIq+NSQgpJ0JzKhG1nUzDchkV3cGJYxyrIdOyBT+4G
yljMMsW2+FfDevbBxqu2DTKaRXbtopiLTwM6T+8zV/OeZvsOvAYpTY09IlAc
qnEcN3OTSRWEgPS6eG4Ou2zyDl6eyFTrlcrIoot5djr0tUWoCX/d8KwF5F37
NtA1oWjWKu9igWqleYrzhyuO28BBmo/HvQUuNREKBOvm0bb0wH1uhkMxWFHL
HlfwO6j4BOD5D01F2D2MBpMxSxAcnZc9wXHMc7sJ3f0efgW6373so8XndDYW
EVK3aYW5TJeguo+ZuJpIaGfAHXUSIzM4Spd+ey6IHBoCl+CfkvJ9OiX4v+qH
s7LjmE4GheKCmTXszmxXdIbuT3Bw5b/k/VCO6ry6kxYCKHu8NFonqk4zWIN6
gf0bFYi95BbcrUc6t2X3xbYDshKuzrnyceB8RVG20ualkJBuUDXN6AvImCSw
nvX1+WUaOoaAt4tMnQY3wQKZ3xhN+aObFXW/p6hRizKJmEJApX3XM1YLfAng
fHxG4cnFgjHpV2MQFCG3Tj5OAUuxB9BExDcCRhYCROKHpveYfHFUGOrcdSKD
gldcwVqe126TfE6N1R5J2W2MmD6lI5/VJRej1nVO0H3WfUpQNBJF24hVtR5o
9ds+9IgkqUx2RrLzlBO/DUp5HVeoGZ7uelZvjTZA/DsjK6xw6Pge4S6/JUko
sGnxwCO3qsR3PLTHGsrMgSVX+TwpDd6XSiKFjrRx/rZtQAwcMfCBjU50HhKE
k6m8QOy243G4ulSIDPgVg03lQke6gOg+JE7egWc1BtsiWputknLFMFDV1t0N
FzhSdQpdK2aVre1FPbTXUzaEBf2NZQCHxrCu/9EmCPQkEHuNWYiZEx4Ak04S
Fs7Hos5lIZIFKa5TFz89x+bxYKFgeOmeBJT2nwl2B+pqLFKTqW0lPVtFR3Ug
uTRoF+zh8/oz+WVQXXOWadrJWRjHFhwvIcU9+N/n5Z2+Ez1zBo4IQeQxMGuj
j+Ugt1Ju5UAIwA8cJUypPPlSe7XVDQWoT2knrS3WONS/1MKgiZquDDTgXD+w
p4E9KvAbEE7h5XinkQgUWiEjKWR+hb5v6TiSXoXwhXIsjW44uCeEPIm1rZaH
Bz36+1hlPyrZjuO/DU1zFtz7ZOf/OuzbLWIirb0A9Z/xMDs4CbFSqMr7Ec2v
9gHBcvY8MdH2Fq+G5FzyLjooG3Sltnc2AbnvJWkTltFN1JDGTGB9ek0lQgt2
rSRK7hFRhxE9omphlGr/kJzqtTMKeBsRhYc8AlJO9Bv6ucC9tYtCzI0V2NAa
AIr8GwFZlTGQFT7AREc3vcxf7org/+qFJqODJV1rabkqtLVO+TB16p9rAJyZ
W+uXlX726UXbjn3gLrb60alVI43ATaZ4R7674fxatLz6DOIc8fPXhWb6o0EN
9bkMWVCIk/NOZjlV7j1A7AHUQSEGdkMHKbxW1IMvQCQzGAko+Lrq8rd61HGo
8xFHedcuXf9tcpP9ppReVQ9u6vjU9AkvFhsOOc6jVQVj2B6fapQgFyr8sRO1
yArIF6efJJthK6BMNDZts3507vH1V8pUkX+XLamcHnl5cMfBXcxmCNefGao+
vHA/DyDG3Z04t6TxxQzazScwrMJXCRYBuuA1ZdD7PG/HW+/yZReff0xsgtRB
o7mI6dHr93Q3UlO7/+rlG0TJGMLzbyDJ9fm4UPCW5wZGS2392iRA9nloQGMb
GFZcft4Qv2O3li3H0oRgoTr0KbeZvA77PD+D/1U4leuPYQZJ59q+s8GdOy5X
/GKvDni4FNGqpKK4GdsAMOYy9Hw3vYR1h48sVstjl6bn874VUR9mxotDW488
QZAJy0q8qn82hET948WIpzcSIpeimNULdZLZ3I6ZbRorQRO4fjCjxodrs/ag
sBeMaxaarxbtsE4h+IZdmwxPjQEr+VMuAtGFpZmegT7YCG7xhUQCu6R+nfy2
WFx5JlQsUMrpoQTNdJ8wbbM3oRpexes1gNtRrUS4aUrL54JFTEsDvyUEHHgt
/R+dmGJbCXYJXuxciuhc2AOUXdnZWYFNmhWPEFh5R5uWGs2IRi5Y+B0MsCj5
BQA69uNw1BLjizv56BR+fILsGm3wMDIcaf+wIC4EZsuK7++dLjDAs+v82zTa
9tNKpfEKyKkL4DIe+tcn1/hCDFrdeTpQBACv7wNiPqAp4V2t4vdzw0BpxGXC
M7QBcyLjBwO/m1w50NTKRaNMqM3kAOv+ldVhg+wuxzPIn7dlkewNYE45ForS
4x0HQPMYnrR2HysKaJ3QCnd8YnouOH48A5+P4j9pZbbIIv4yPVPbgkKLuYeh
ECBW42ws8KxseIjM4opqVpbirU/BO51l0wY0EjM86DPNJ3+qUhNZEK9OfcXa
4K/9zrU2UecUsYM+rIy2VFB5k5s5ke6xtijEHyTcFu59C7lLVYEZVFBls0/I
tM3JVVuyOyEt63XEGkyvqA5Sy7QBosxtyqYiV2v22pRTR+mvzQ68ztwkJdgX
HtADqb4qDXdOVuNACF5ezPrxn7Icu+9IsC2BoUE/c2jHZNwrTzNyPjIK3XwH
VMZgVPLavc8M+wWtzK8ilMRbpL0ZAdNZ5EE2XPjKnNhqdeLZxQrZwW+LJjXD
7TJzSBiT+kOxIZ0Zmi1DXOXBx7FOwFsu8JFX2H7SOM6KdhuXN9LUhtuwP6sD
mqatK9BfCbomxGJAajKYXamCGGeUDKp+RzYSNxf4Y3PG5WVC8efNEqzYqWmf
hFxVja34ROxiQHxiIojur1SnB7niWcdgRAEAxJM6CfVkrM4UN4u8AslRh066
CxVN253Rn3dRDnayeqRK95egztZFfbTISTG9mUh2oOVk2cX+qGnAKGXIn/qP
L+LpkGM4FbvqIRw76G1Zo2+Jnq9hSQiVdftxreuPanm4WdU7e2VSGcFp61pR
xvEFKkXRkw8LT4WFmrAK85R5rL4h3smB3YUFcIIOr6WfwpHZy7qrBRnQpO/M
kfbnSbOsPAa4nUaCPRlwisBVrx+8ZeU3KcPW8wWOszPm1D67dX3j5mw2k1Gk
JfyJCSUPxHbihRS5TmocLjifXXvexxvehts+e2ZpWLKi3vRTrQW2lYN+BEXd
Vor89UabrClHSmmcsEJx7qsm5sbcHdX9DQGg3DX7YOHU6qbwH7H7dtoi9fyv
4/b29Pe2TvwRiWKABTAu7i40Mu8FG4a50TZ/QBGZCMnUut0oaVr8hm9ySS6T
BChxAOfo2hq4LRqi+7yyn0oGrNkX0GkWNtdAbz2J/UWNL3Fy6Vlbvbs0B3ne
KBNPquRSC9Eqd9L+fVxD/kwhpF1X7tk261hbFLb8DXTG74/o9l2xuab50AFT
gnhzwHGEj26OFuO3sJraPukwTxwxDxJss7QX/kZiZ+w4FwvUNAk/eB88hRtj
SMoevSCClOQwTONtH064dIc9UwnhqtUWIWuUOlAJzFnNrxTx1sMVum8V+GYb
wxfbDrnToj4jrStHF1/oxgSFNFM89ZUzi8Xr1nhfoBHE8x4AThcTtt/0ArTs
9PYjC7472N3B/dtT0GtCjQk3yFB8Kfp76JpZGlZpITRgD2mTOFjuKKnC5mWl
s9AMYk3wtZlgKEF3FfDbLj0IqZbt0XxQG74E3PTaL63bkAOosmeZlDD8nS3S
ZpPAQJ6ZjWdzIc3mCSbeoy6CDfoLsDlYwyq2aWMfZ2ZjxZfjkPCVNwPEah0f
xsctRdlS2sqUsnVRnSLHrX6PWOre0OUe597SWGIZaoq6eRuBikU0kgGKAcc5
UP0WpA1oLUAoPjsmTNEMGox5OTPIR//XTSd8VhEDD1bkukMccQig3ylkgGyD
px1YrOzuxgOCWvWkfKIDdfQd7Yq0fWXFYVg6Mj1O7eDagZkyF7HeT9Yav6qV
7CMpw1J/dhoAuVe7ajF4TBIJLpw9KOJ9HF0sRi6skfWKjezIAsgZTEZFqoUQ
TIME5rdxaB0CjY0WYRc6asfDdNGk/3vjJQ44gad1WnAYjXJD8tpd6h53cZfz
nDUPjZUXn5Ig1+OUwsJzQxAyH7cuiI9FRqTYkQiUgWlKA5WCogm6uFOPfVc4
yU8/OMDwzKJg4eBLqu/P6QPMPc2pe/yzsv6ck5Khvom5+8fNvjwYrqq3q7XO
oCuhdJM2QPKWFG+2eFEqpdkvF8YkRMs46JZKg6AjCctIBYp5xHbJftPPhUpr
mpQ4BjHtOXniAzI19bcvYRlV703f1v1vFwpLV+T3uTwyhv1u4bg2wkpkD8Na
0LsVk+TrzGy/FhKCvbadpkDBqfEx7Q2rXyQ1v6h5K6X3HFzJFyUEeEJY3qaO
iYqkxuVQWK5EARncaSbHvlnmUPDJ3AWx0QUvF3wEmvFr1rvGmJ8Nqou/JE/E
Xl0RQUFQ4KOcj+016ktsYSkNPKUzl43RSvL40CiUaIzg4wn6sw675Hmt1Os8
ILwuLKmLvr8pv1LBlr03SbavOjTR6/mvQl+lQoh8cNi0TlQr+7eDvrC1Wdf1
8gk+dGWCP2suv8O7UKZSqCxxsth+bOw+rj1qiTfwBH673lSSnn/Ur/uZ2vYb
kb/B8itoidyeZZ3H60/H3EQb0MPJ0RK8It5jbqa0VvmfYtsjKisH4Y8eNYn5
YIsFb3EDpfqFi/OZd4PAeSY7igHcb/OhHbzh66IDt0MiVDvYWu63qKqp0SZk
y2PPgVWRMlaO21lXujxvzmgynriGBa+auG7z3nB/TvH1WBy6wrsAl7gAITNl
BQoh7G2xvMX41Oa5VdNimimb609KvDhI+2etaRDRnZyxeS+paW4l/8wpE8M6
B0oQtowDIHByAbaD3/Ieo0csRKKBfsFM/544kK3IZ1tq2UuVbiCBPJzKlPek
hEfszdQRI7L69FkXugeSNEJKEhHSANAYqJOskUmIw5JwriAGmWGvFdLpG8wu
KY25evS0k1VjWHVXBEDNXx7KVAb1YOg/JO0X8XBWzSMetTzelAEhEnYDTU46
1ryCTqTCe0e0JcRRrwiWSGLqtIdU0pI8mi5tG0pJ7dtk93Z+dgBq3q147tZm
LW/yuCA2P2y4hNBfP6lY4H4KGFb9bG6naV8B4Gjw/C7URLD4Q+/StXd/kp8J
DUIdPjWWLJsYdsXSBi3RqeG0+ZdiC33Ox2UrdAdgfb1I1u/bz/QVpbycnF9p
SJtsx/qrPrW9qklLr1gk1R6rn8znLwTwd0mnsDi6Io95Jey2K47MlA6H+/cF
oi39hsg7NcFjOO4dw/fbY0kFOAA2fM1zWkKyWmyDpMOfcdUtE8jG0FEReUZ9
9uTABOWB32Kkp6+hIudbl4qXuCX3RCy/Is+4lEVN9zYux+4bESyTKPxEIHos
1KoX+zYZlHsYpQngSkv7GYhSMaZ3MTqGZPkpKNeGBhPLCjY7d4xqQBGbSAD4
iHV7fQNnTdJArXfGIHtAPkd747L7mSMOhhFAxvLuORdoP+tM+tPGzFHI0nbY
VkHoidx6EL1eVi8d/oI0yRwl9PR6S+8NNxtaPn4iUDWzL6wHFsPkMvofPxjJ
ayvJgRL0QEn7h41/XnvGp7akS86ELvsEmeeXrF/UYPAgRLWt+PvCxjoQzptt
6IT0nJHxrbcYMi97r32UMy/nk9/QpqDW2atNLiRetLITjUT0+Fq0z1AHFl7B
lhfxf5sDmfy8hxQyNimNdcGVv0G61cApQCZd7AKX7I8DkL560XcWwvEf1hF2
RALmrYi3g4LlkD68dvIKoRUT/hl3IfMSPsgJypU+0gcHqJGiLycuN9BjMRip
XTXfsVX81zbKud5UndojOWxltg5+/7KnyzRdTCxDRSVhud3OTD0BrD976uqE
HLXYrD+NGbg7n+Rlyei9XD5IRW98akXN+eD4d/VNRNqXu+//A+Q5eWvOBcN6
nmaZNPYFTG22vS5iS1ZDp4sn2XWmOHLl9UFoJGKZ+E4FNP4Cm0+RP8jFmVyl
oTK7T3A7WrCYfqabYr97Q6oXNjiYlc1KK7Zk0k7LyX+sJ1tSngD+0/B4W0Fu
+Odz0wGt0UlAFsb0WZ2rx3VBC9ev6b6lr83A1gTxANPElubP6AwaNhq8MOpp
alrsUU4PWucHruSHegrxO5zCWCd1ZUdhGPWCFnFgr6X1HcPUY+IU5kufVK88
oGkVssW1BpARA7loYn5k3tD6HRl1p/cIxX8FPK7QnPJqVaC8XZeKhuD6U97F
Q58DFnOj2VavJvOobexHVEHcIhJN/2boSFtBhkmoib2bLHWFW7pp06DPRnuW
e1G0k+pB0lChPmVb+p42VJRxpIttNkTqK7XmT+kbwFvNkrUXY87dBrltTTE/
TBAUx4HPPQusQD4bFxwbAh3dJWbfxpMteCD4U2b0qEyYUBtHsfQRkvf2N307
96jH2YikJ6q7SZdm7gMXzcRLZIE68kJS73O/j53vaseN2QpD6Q747vulA5Ch
sccwgYxoZIo8pebIcGtNh+RTHMsSJDE/atlaPXQuvyARiVsL+b4+YF1s59I0
KtKjkwjYccrgBBhb03lZjGtta73NVU4IIfmJzhcHuve08RXD7E3AKXLN4fVb
S+QXZYX431NkXkS96PP9lOXZpJHya60lKKPFa6tNgpSGt2p7cvDtQw1uzPIn
rGyjerY2e+HhKCzxBe+gOAkAzE/2ydbFpDHNjqdeHUVr+J5wsGJKunodgYvi
qeGv7KMo5l16YNwVaaAKv+Nn33Z/BDU+gN1rTgsKBtvcMaRTOnuEazVlD9rj
CWrLYzP2q7k7ATm9+buQ1kpGnIRXitwOD3gL9bbtvDWTMmbGLn5Xgdxp3c66
ax7Q3E0cmAhtNwH99VbXWWzfNLXVMVTNdvPocfLP33CAN80hOq0iamcqVsm6
YaBlTHEgfpyI1x+xipswcB0S+pvuLnCDxitlgDUbcJtR+nAPJ2VsYp9YkzcB
3tQtJykENAxhSMCjyFAiuwm2jxwqfPzZ5Yg3ZFQc2TKjf08xkGQ1NE2kgZR5
PvevVt5Pz4GFLLLN7VxHuNw4FTYalOFOR5KBkVnnTHeusKaC7ovTdVtmkpI/
9RFu4dH9dcNYp5Cle4Ce3NgL7ieTdLjEwL9enk749VQQKVu6CljLWieZ7FBd
/kFRzRVf+u6Bok429AHqc07Lfaxj5TR8Wt5HW7DoKhFTOiGjsfuqjLvOe3le
bW5SYV1MFn4WCC4ydVNeu2bApe3oJUG9b1Wo+ARjjHcxGL0uHO1UubBEm4S3
Yl4Dt1LTTrNr4+CUDe1uacnLZtaFOcDiGqnuQ/2l/Gw0ozQbQlBWaZVIQ4In
lvmR109AlWpzTHNR1wSzJm/Bw/vUBhFidxCVeSJsn9OeKuTofiYPvMFy7tyP
bW1cAZKmgthJKhzaA87ST595Zn5xLkpzc/V1jGrRhsWsPUhDfNVuSQs5j0gO
eS/i/NXANh7C8KkFPc7/BtSrPUWDhpLimIjpDIAbWxN5GXvRIZFrtOww2mC3
8wRbR8FVX3fWmV3Kb9Y1qP5BOUnypo2REsvpzdh8o3Rk7UkjzWbNyiftwK8d
+mER3ZbQHOgmcupOuVrSw+pSjY24fJs5WBtTpLMtFiwv3invCQb+LCystiWn
x2LQkmf82uTbDx+dqTiwVZCq/StgfW88XuENCQsqHnv92ufsEDkJMQjqHxdF
4pjhGnnsY4Fd8Aaz7i1YroQEX7nkPyqp7VOzKFfVPsbg6GvK1baBcSx6+Gwp
HZ84LQUV+vDONYTvtk6hdDqtItiZ06aGL6JY2V8e5apHg7t3GVUQvzcMsTvQ
W0uXtSbtLqRrXfbHx2kbsZrwSE7HLmwMuAdN4V1XKFat5ouRS9hX90i6ppMb
cUwq6godxByQY0BpXanOENUj2yRsOQupNK0fubJxpZWHtVeO3Nc0bR3z38MB
0sWQdRFGsBLuAnZXx8Dyk0uxmjZFUHpYQ/heS/uuaTHz0Lbl+Xxy9fpc8CUj
izJ2o2qLl5TPqfDY4J9wXFTEOAFJTBJ8XhNiFl/rAJu5xQiP6HwO98Y1L+Py
HivxRHwV8fVGg2haMyVY3Xh1y/AluvseV/M03zINjVca7sIGhYhesQr/xg39
/6TlfOsIHhD0Xd9QTFE5piWHOvXFtAAfV6Jq9OTjZkehdZmJuyHUZ0OSem5W
eDnssKxXUxTXOdJjfPbQBWPrMzv+oXnb9OUTUvfEIvVs6fZs6Vy6FyL2NvSK
TAJmkS8i/uckdsc262ysplnQxrHFmULjbpNzenwWOUUSBe3F15uO8sdnBJCF
efZvbLMx8nPSY50/Dk2LfJowTFf7ZohKotFNC86QB242OIlj8AAjhQ3ani9z
DCbB1F44rUbHNndsy9Nna4SglEZbjmxzy2U+xBqgBrCONrec5UCDNOxWnijC
/k3hPoJjTQD5CxxmA6xyPOMtTM5V9rDTuKv6qedYKxgCJjysoX4oEtCde2nV
bDoVtJvkTksqWnyvT+4cEFeJQadgLo1hbUExq5UvFm4NVvlrhi8mX2igHxMb
B5rGO0LwO3jrB9Y7nxAtDpKA/qQncn+w6vFAj94H74aUzwnrRHaolGtzjWNn
HmmqS3zgtM4KHRY46HykJqSZKC7KAc3ChwUKXNzta6cYcImtKlghlxO2UfoJ
EYaPJbccbREq5J6Km9mAgB/tXuNFEzodKiA5Zgtf48RogouXFZqD2zIMNoyA
kast0X9XTd7VRsxfZ/+hHXJNfRxaFgAmYe4aW+id36OBcQV1UUANYmjhkYem
0+6nzk2OfL4cCDRmT4/ivPJPmsMBFgOISofOFYOEILlOW/5KrE4yi5+SlRXx
x7D0TZ2hO7kB29S3sUolZvkjD4FALdcoZNSPXUCF1pCkbIQafHHtTEE4Zk51
kWhxKDTzol9RAA/37ehL37W1JIOUXEA5ntGOblWOjBTY3vqHeZvohLP/BezZ
xzGvISeSgo4lWNCKEqz6tPOYEYCC36ji3HkE2uQ09EM+QA5UYTHSK1zsUqkE
MMT3UOQXq28JgNmlKPS/ASQjm7opJ8hlNnEIK48esI8GO8vusGq2StMMO5Et
lBwfNQjU07T4mkqhY8o/x8SxiXpIqawRevFE12Z88qpXO9xj82W9BZRv53zG
PaWk7Y6sgpdeFGjsO7/ptvVwrrT6mBJ84RSoC9cAUSSHTb8CPrfNTkjdcJWS
ExYVwe/ZLcS/YlAk+AKm+cJXXR4CUnatXeJEIjy7nBjtfehDFnLuLjY3FVSy
mVOVGnLdEpH3kRWcegoSl/1oAq+P8ZE782xQduxXYb/zE9nRW5lUMhl43++w
mKyWHJfVLbaU/cTKC6dIj8KL5TcvHb3QW9TSWo/vVBZ6Qvstzsa+Z+dqjmzp
p12dDQF23ny53LjcE8X4jfg4ZNH31oI/nBWFKIIU9VA6oVRW7uRnsOvzXVce
njy/LfJ/Otuyb/tktKfRTJCwtuEEJg2EdlHtKrI1LWNvGHQy1n/G4bTiOnXc
DjPKI2rY7TiuZx8VBHmK10vQIuJe5j/4PQle+jT11UNldd97jAY8CmCWnVCn
ldO5IDAef/VuJUT9zx9ikA9ToeHHwcGmjMLqbFUWpi9SHTwcPdHVqqfdok7k
LZIbl7jKtwmtugiyW6Gdz6ojV1y+adOas93oHQVXKxO+mCXt6leNVK5xEfsr
84bXiJpHUXvqTounWJU2g0aeb9MWo/s4KCdx0K5OAta28cpXnTpY7LaKwXJd
WJXZyT9NAYmGKAeeCmTK5B/SsOZJSK6fdGuMx1xit1b650g1cwL2JFKIVHgR
svbPUSP2PQHLq3caneWLl5xH315GTPN2A8t28FzEtMKrdt7gaOG+60Lyy+/F
Dzkxi3eNwoNNsWPD84UAIqZ7/qUo6xcckE7C+PX8CuJ1jRErXKqj7nr1/7/x
x0dbasFEMk6DA++nFP4zhtZSURi89NbcgCJaBCjboIdvffQLMS7CGlHmIqe2
0x+KFUurOU+DXjdze5L/Hz4NwHqxOmmDhN5+KtitK6uEUDbzpVtp+d5stjJN
OwIOPupI7e8vYLdqR3HP129j69XHnBCc5QSV1eaNkt8tf7Eb6WgkPy9Snglv
LdCcssMns2HhaMxJJs+SSXMhPekKSpoldF3bAQ9LosWtq+jCdEn4HhaemVy4
fv7htthmp2Jo5TtJdd7l+T3X15Zrxy7sSAKgQmGW6IXsdVcxbKELh8ZMyi85
EIjjWSRuMW7R/7cSf/vnjf9ho9/fxxMjwg5DFWLsER+TkkFpF3ItyiIFgF4R
cZ3gkYXsnKg5dUvKW8frjCIq6ow5XK0p6//d5Ql5QA1+a2/8nb1ARXZ2/phd
PsalbvKps7pkfxui39P8tLVB+FuG8N6Y8iV0iCD6jGCJ+iz4Xzqpyub7i5WA
wb2lvUjzu67FVEZindEfUlFsqfGOhwh2TQGq+UrIabJs8FPidrq8wXM5VmRx
V1keRJXFiTx/ju1pFgY76SKVR4rkK5ru5oNYZsmCqZbF9IP1mMRaMAM0X2rb
D3OYGjMRwgglit5+NWvJJ98gHHPKWKipMbBLcHJTAXJoZz3mavMOxvV9mJt+
jUgN13tUYjOKRt1B85Z9ffKIgHiF+B6pR4AV/4ha5a96d9e3L0nxD7nTy3tm
rWoxhNiH3mS/z3/MpdSNWLX2q0YGhFzEDPoYwNGRTg6VsF8lFUu5AFl1pi1Q
V18AxNllZG19HtUsplrg5pihsAuPXSYmlDDHpHzBkxrRzBjSno6nNnPlwoDV
JODqY+RMhda8CWvSYrbb2Ary9n/g19vw+LMhFpNsRNIyjpDVJo8UyEDzr2c6
S52KABgk+01z97wUuNFc12oBR58yHsle695sen/AnpZsLFbf7xK16tDCB6k1
IAMjXDRrFF4AyuHlQ92Tko5gkwmJhTCjwSvKbjkCP50qQzvjy9dPVQe0c19v
Fj+n4UOaosQx4buYKlsZKMdZ6aMf3eRHxlY+ACsgD2yboql42gIRcxBePwMy
LZ1bObDdCPQgw1ruksaQmgz5KbOKCgThXz5e3zUMrWTfcLOwXmRv/4SQP+qa
zYYcPyw9GhpDJ6pT977vgIm/goUNzzDjMJRYb3MNbfIuezS3cNXtx+FFrBI4
CTiXGBpJVv2DbneyQQgcBR/QUks8JnnKlxLBUhnszJPt5RoIvuSpPutPCoeb
nN6btMnF4lF1k2R7T3w4EvxeFL+PXzA3TDJlkM70OckzK2+mazYVL5wBLXZU
djtyLNlLl/aY727XcojkO5HJ+GbCJDDkYwwgeXj0lpz8pnALxB/Nlno4lSUU
hcJ1A0qxVYbFans4MBQo7eGfq6F9iuZZX8k7dsxO1vxmriWgpEZn/rnygf5p
mCl+fvGjbx7kSYNEphkedPNxrQ0Fbfd8H9c6Ku9tloniNQZ8BI6uXroIUtiU
mNnOHWOgXyLSs88MysRxXQBlzm0yq7o+cVzah+KpPzHc0ottlouXD+4sYRR5
Zqf+LIiIUGahiofWfROOREfRRH/HDDsXEuAYIWcD85D3GeC5eJdjkSjP3ufs
W+XIpQsZBOBhCi1Ka7Iz0JpTFftvErzBTput/DpYWvGOnbCvimFkuJC5HydS
aOY/syXsZS34bBfmit3gqq+pRD56Oq5q54gQDURgOZ1+bUl9bSPrslGzs0tX
R+0YNXsdJr0PA/GTFKgASGM1aGYKfWqovSebb4GkO0hXK/BQQNfOJt1Hr4Wv
s2Xg/aGcJZvZWttpDbvXfmcrY3q5CxdW+h+oIZsJB+r2mlkCdpcdH0FEsNP5
VGBqKBthBZcpXb15c0R6e5O9FuAMZLc7rbAHMULKRH4JNfQtUxtYgQi89Nwv
/lN+qxzf03E2NLjIh3cWJqpOrbKQW72nZArWh/7vIUHsjcrzuuS8x8ILWhGo
zyZd4Hts+pKEpVRVQD3GyXa6rM8nadpWh5fQv6dC9AS1Ydo5eVNieu2XBz/e
oanteVH/Z/uvNb8cx0ZhvSQ+P7cPYnn05cWN4+P04OUpCk1lFF0fphpRvciL
RzMIJBqMPl1rAQKN9HT1gCIDpf838emJJUzVuzdQnNXTX8Chx1Psck3DQcye
LKiX2E7ZbS+K1cso+RYqasZyKEdRVHt/RClNtoeHwOZKS5awQZHS2ZNFvjAo
yTsf7VzP56AxSIGBCCtp97BnAts142La5AssR9WfzYsUCgos8n++KFqXAWjh
fwLxDoRcl/GMJMiw7rlM1MU4k9aXp0GnDrEQc+BFAbIp6St1iqQRugFhxi+b
fA3zefwUElN6nBVXgjYF2ebdrmG5LPYZO9fzi8RarhhmE7cJnozJVLlFsPT/
U6sh+WFl9WOcaJHYo9TGEhI0KTs9JW6LsyoINEqaxn2Ms7pya7eWrWFrgnbZ
ba/si6kbE8PByU3P7enXYzF0VcWhCyF7zOLPgxhcZutigRE2j2sMqJuRLRwl
0Y9jJ4M2YZzpKe5UtzMukPmMsDPK9Pi6Qyo1Asa8yoOuNeefKo7pYuXidXNP
u0PL+wE3882hExqYNmOO6+H+LGeH82hI4IzMWlLO/fA9Ak2zYHC0eO21H6vH
+xTKhz06rKoxxKNgSsSto8w6Mjd2/flKfukydWS1iKMdlUHTt0tB0tRyh3j+
Pku30Hs/flAAR5Yp9xG37gLm0eTCdtqmr04F/CWiOwve26TSV9pYYIeJSUEV
0+4xT7XneQstu4qOl05spBWKyHx+TKPlsg1bZCPjQv7IVpZiNpHdg5EMqlMf
ErGN91hTIWhTBKhu2iCwT65ZYx2eJCNJH3g2rYM4LXTcY0oVTk9WqHs6gXaK
N5RlTm4f2IU3UYVGZHdN5IqDUJRej3KZxXjYZ7LQ1le/aQLKtPxIOGSQFsZl
jr3Sh04N5BnMXiJommYnbGwWLsOjXYCNmhM0AqLGEh+otcFnewafjFUo0L7/
6Xuyedjn7QY4Q/On4l2kPoC8MqN9bKPAuX3b/9S47nMeBoFGypCvCYafgtyI
NJNMQXz01sFtR46bgq9Eh6VnehBESYIOSiDoeaBiVw3tgD142iT0xfKTxXNJ
SHSkLbIZRSlFMcVifqlbRiMFqEJ7jIRCZsdst9wQ1VxJKG3RF1IE2BjNnLiB
j/FUZP4WtSWO7Zl5pgkjBUBMreuIOWX+M/srokTW6VJsu+kvi+wnxwsqTsPA
8bCOYV6auBxcHTrpt/FomEweidOEkN0mShB0+B4lB28+G7xf6UYvwsdhwlb1
Mjj1uM26YMj3S8oGpe5lKn0O9AZBif0pkzbkOnodW6LazeVxNRLJJJMLkSnw
XmY6jeZrMDdsahzS0I3pvQPviQdPtx5PbsF1SfO0o1HsEPENWQ66C3Mq5gdt
FxZwW3sYqbY7XwHAjAFKGm96CJMandZZ1iIOVYCzoQj06n3lEx7yPqdXH1+B
dLUdnU9cCrnWKXvK6KIDb3Y49ZnBfg8llLb3oTE4LUAPWHvTxYe3ZdHWgsKh
uO9mijJHLvs3sJdg3rHzchnUllFb+jfqw001dfqHkvYp7NWjBPqtOcqzUdSx
KkRKYrnBK/SUxDi/un0w0Y9FV7FaAHnlnL0h395eAs016D4gQkm49mIr4pvY
VPrRCkFIumLsOfC0wJnTpXYp90F0GcrOsDQGjQVY51ZCibaut+HDz0Mzd/Ma
Rv+Ml4oM04M2AFyXUibNdImZkkrrMo77M7t5Hf6bmvQEfr0utP5R+dCWTVyf
sSV+zp/aQYXWX+WbRLxBZvPbnJfkDQqPMNL7WtCr+7Mt7k5uxklnIkCxFlJx
uPTb2QOugKe2QmQaj1n5ZozPouk2EkHVw7loi81PampnhflICiYnAZ3Oqbhf
VqgJbt7T0XxFbOhTQCo9riZc+YvksxISWeZuJ9tGX8JLehrelX+JyvpMU8jR
igY0BbanYUP3nHSiVsn7ma4t3xZ5CLH8E67JtUs1rrHsyfKkTlpcZ3o/w5JX
Xz/yCqcjP84dfEu/XX6W1amu+bapkJe9ARj5eiTWdbofdu0MpejqB7nBDwQJ
+j4gyaJYpTGW/7MxeLZu+fY8JxNpfVzooH3li5rKRrzT4YyGfMqw9AZabqeB
48/0BAYbNwF4zO4rWw1YQKhimgagfW4M6KuC12o++mDig8GzqsjMvj6mMXHQ
2675ai2rBB+BYzcOzTMt33b7l+VS9hcngItfYeTyoDzS9SEgOmmGYCdULHIC
EyCAld7iXnc6N68VOJHELLqcXDApi+GgmHcie42LtO03l6eHhs1fSH/V8xvj
0nVZncCgb50l6tu2lUW8l4mmPzkjHfHYZ5EZG7a8yA6weNBOQ/977Uy78o0r
NXotoqD+zTjqiGO50X4GnXbrocFArxvZQZlDQ+48gCbLtGReuXqfnVFLF1yC
r4i+h2tVxuNJ3GpIs4uqLHAc9vLpRSkGgAZYT8z15YW7yhnVkBHN+pKSWMfE
dfCs3VTvnfi4J9mQXKmbykQ2R1kciDfsf5xKxwVAF2EZ+MptzAGwK4/2dmJX
YrABYuXep7VA9O7WV9QIqKbjOJ5NWc5PyyvAp0NOZg64gDjt8MyEOIYWYXjJ
77hZkvA7AheBp8Alkh9vj/XgWEmqnIseQjVNTwDH5O0cCrhQxjogJL5AYey3
vtnRLL06a9rXZXakRaUxVq1ZtlH9ZMRqX6fm5TTZNzHI0gDH1Mf5r6Zrsbcq
xCZ10uzXf5NRhuo9Mqv0aL3g2UTl3WNq3/Q3qwPqkBg7RBip/cd1uOqBS8mc
fuYBfL8GrYRbHvfGE/Zi/l2n8cX50f4ekIqjT6/l4Z5lvsIEq1jImVTaeQY4
Yrk6oDpYpnbfSiwC5sI7+4x7iOEUN3OjnQfav6Kn5Qnblspc8FhBnRIox7Cr
QiPVtWIeXzeZeKoQ2vjyZ2BOqRPpP5fxWbqVFPpOGniYx5UFVhBTLAVHUztZ
mkF6GEFprruIwRn4qc3QkNLf50UZCjrYXnjiSXw5nEXc5ni8YYwAtuZWYY3b
4n52QXE+Dq3Zg1YvkmfE3H/ZfXuVFtn53HsWjq5aXA/G0vj8gl1cxyup9CIx
x6KWrdfUbSjaZRtpY1w7Ch9z5YF2of0Kjxm/JHqJpeVvnkooh7XbfjoI/PtW
V2dLQAygemFjmbrco/MODLDhd3i9gzpCmaqaGcPcpjooWS6rdqVGOjQA+IRU
cP6OTOuPWJVECRn3C7+IRkuIt/xBo1T7GO/ib4NS3z1EPR6vZts0EXfpC0az
gvnE57vypMdmFOqBQW5GgxjgUjDAhtS9lmvBAKCa1HRB9YPCtMLyOeOXJunA
p6wlhjnS2gayLyZ9gZ78wbWio6EFbRUFXWAsPlH97ugSO/k7oZlIo8JDzVH0
eHYE5lI5jKCEnLhh/FLd4waJqT6XXGHBHi+qZY1vHejxPgvgIMzGD1qCLXIu
1BSE622/XyoytBoR6xJgr38lCvG/9yxxiVvz0h06T/jeaCTVwPqtFUypcXnM
6hF5z3WR2sUQln+Ky6LrdQ4X7OISVskGQXxwidmm6ucXIbYarwNvNQahmlon
IhMrS28vo8za0cR+8IjlM7q2TlUOlwGC8LJrSF2dDg+aNI9J/gQa477Zz6TP
+RyaZr6nEw9UGO4NHUjjXX/kRO5MK+hvEq4fcEqIvXYb8nzP5RrfaNdFnEtN
72h9wY2EOp5VL9+q/lApaCAy4qz1QZIZO+yb/0Tma0IqVIGgPDpKsVCa7H55
Twkidjt2LW9jc1shtvevVsbN17T3gIR67pM9FW6GHA9BFNqQ09A8B4Jor8jp
8i6x2p4axWzC2KXCzSoWHQ1+VvHD0d3YtrP8bso497JOw7fW8YL2tqLABEcg
gD71nWuqS6EWa8dzYSTJkQOU1S/kMeB8UzvzrpHFckGhmNKiu8md1jbZw0hv
e3dNRkGibYRnKbBoNMQRH1OQbpEu+AZ/53JsNg0N/zIwqUj9F8SJr1zo5bln
Lnz6IoCz1f403ciG4628TCKxCh3mTDZJb6IuI6Y785wZL8Rubs9eMBkN6Q4B
3K5H4nl/kMIcnE4OAyGXVL+8az8eiwdvy3MNd49ZgQAxfxgt1LKfbStpUhQJ
1oAm/SfQjxzys7CO/uVSNDQ8/n4fs8sZCBx76UcRLLSTusRJNNRHEccqC/7n
zggWLODKWY/0h4vzHP5g2tb3+wv5ygkQ3Fbd8CrSIOMxOQ2WIR1ZWmJRuFaR
aDapyGT6sRYTpvrPBbINc5Dr8Px5rra8gATPz0AqG1Ta2r4+8dhhSbJ2bX2h
tK88snyYduZp7VpEMuSMJeOsEzkv0tGKJg0gXfmupgPo/OiU/gy+wJlprFOD
UmPs27udpQae3kV0fVEhsMfAr90Lw2x8knnOK9uBNZbBGp9V2qFWgwcj+l1R
Bto+66xbbu2z1+i7ij33mNBCf5bQ4s5Yqks+ewHQcuEMxwT4q6oK7CBi9U0r
0lMmnDncV/MbPFNLexpn+cOdNI96et3WVQFFe7bnjJ4iCmSFTS3O7DdyKylf
xINq2wDnNJ0BFif1Gwx7+J/y6/114KPBoHgBfX4pirQwU61H433R6XUtftdy
O0V7UuT3zV3zD8FeU3C7nKoBXUwbV2PGzCI2izzeTq1LT8pvrD3n9mAw5KiQ
RRlUowFrM+kiAVLBnjBqsG2X4ao6LvcLFR4Y2YNqhnTWeDAZVwC0X1wbljKT
zUTaXoQaMskKjVUU8kRLNJR43e535tdjGXfQfTk9FvzNg3OboMIhyp83QrTs
mwQKr+AxIFVD13JiP0SDzRyAMFJm9RwtpU1vSY6T93yFcsfkAFscQfxa8WvH
saG7w0IOyGBf/odwZ+DXSmCDnOiJjtIcOMR6brBZS0KpvyvOMaOCjRlORsmU
afbUoImvmM7PQGdzfTwr9IK9+YKmaN0dHGQv28OdjMthVmMkdkHWIzDnE/BC
SpTYke6/mI25Et1c6juiwrzUjGGivfQP7uk6UFfPLnkwWUsuX9OAQWm/UFMO
9YZX/jmhfL6SiFDUsU/qFd8jqXJ3k/WbkoaJJn5GX5Wy+k+HDGIixUZZ1AgF
FBdQzhyX9BSWxwrImmvAStas2sBUOgaZ3tVLNLJ98veEvvGvpSdB1sRXJMzF
TBISZw2WKqXamk1ABnVZXDIvMwvfI1CJdwQqU1Oh/KxesRAqSTyh0i5LhJgL
F8kC73YocKy7pOtuhZ9FcIuSqGMNaaexM24Uqiuw6maR/dVT1qGzL0X6TevI
v8dAjbk1zILvcWE5IDkW+f8a4MsudB/nD6DkaY1vrnNoE71WRjrls8gRMjT2
3tNPYruFuQVUILAFfBqBSbfn93cO2Oh8Pcq7kXHUZZd64uhx/1xfqcDEqoVz
DrAvR++iOsU7BulTOmxBzmZqiABL82YBltIYn2pq+46cdpWLh+9z4OQyFzyX
yEkkXwZaJWuB26KpxvekJwWhQUV6sj6TcMeWoDw8l56YhFVs/z9f8+CZX2/L
8ewP71wHGNPYEdwX7zVJaSBou28kJ4vt163M/D5hm6d30PRafDy6QzO4De7f
q4UYWPLG94nY3Bbu2P8phROFtBLZGvo3saGGfRKoI7fVawcxZWCQFIzIq73R
HriLPNfvHW10TM3Vtt9E2hkmJbbtIDclXICahEttb50yjQl1x8M0CTY+E7By
kQdX+yxKj61G7uhrwmbl6ndkpNJiFUtab9q8npO5zBhbgb8I9D9ckJUk/8BQ
+9LJqg6AkE0tfDUVRYainAOhEQWLACxS4mBDXYXDPdsyIY52ZWqsn0oDAKuZ
1udLCGbeVK28sCNWYAglcfWI6QLUeJoYtTFvJt/kVBfYl/hKgO1zO0+6rgYJ
VUtJhBSe0pKtGRw8y2L3WmafMRQL2paHErSpox5lG/nuLRAfLUEXQn18hWQy
I3hJbf2ZeM8hLKCtfRBNjZBJX/9A6moCMV3JuHxKxOE5xZ/hp05BjZilrbGn
V+r1mIf4ZEpaAcjmCliJaRsMxbMlCPJ7bjoXfBd+WsVg6oL0odMyvDa/0e0f
AJ4Ngy1fiJHv47kFL2OGqcJcSokCVmQcB0xyGY7ot3p+Xt9BlHBaNApuG9aM
Tx2/8Enb2zagq5Xn5zMX7oQ4Q5SeMolWfcrKA1ZcEeNFoyFWox0lTWWeqBMj
xcvM0a6/zK1oOFlsMurIq+rmINue/IIxA3Gw5nGIW5wQac3QweTjmz0zQHqx
ASEB/fZ1g2VxdUCWFpImHe88S10AS4JCzy39hnGCqQEikox1ZKWELii1WUTT
HZkmB9OfxDS3MM5flhExcB+mXOpt45jbCQLc0+DX12N5oEO09zgEevIZqy36
W6N8p6T4CS8iWsr3kYGTNz83+ij6I4AaRzIEsMdeJJJicL6Vc6/Dkf8CJGDU
SLBF95lILIrfpddot42y0XCFANBqzAKd5GLEsqVTVOtw4N4YVUoDLQ1WhmYE
dH7MtKW0ESS94f7PSwbtugRebQz7D/bB/KCyaDG8aNPT/j5xYnJfDY3wuV7n
EL2U79KwNVPPI1cnJX6j5IOhvWL7X+IqWqU+Rs6QpiZvNOktX5TMgJz74uW7
SSHW+rsBT2nBpz4klwPzDY1ZT0iD/4rOd98hNGuYX5uzBjUsAS7IC6eOpskL
UhpUjgTK9xp/nTB4RriyD8oesVE0fBjjSYqBY2XxVjcAkaAUVrgGQDLZsE71
JfNSCdDHMoWvrS36zOB6Zv4M3qxaxhms0rwVKbm50gOYc37waAKOy/mZJRpe
Kia89UPCeHxnksefEyLSnw+j5erbQhaw0fDfC89upcl2/54t58qACZg7WYWV
XEaWoBT/GKoM3p6nFNjOlCTEpHuzTh4BUz13ltR8gIkSF0VbQx39U4lc3cjy
aIEDSGz5uzPMI1hCPpZ4iEQ583hQLQF8yCb6BqX26k10j4OOr9M1GsqTo7ne
neGYHnclMW3oc34Fk1NhCp6+gxQKTo50gPROhOl2blva3nzAVOfT/U3QvJBq
Vldjy9SId+H4LB3kKnvpfaUhj7CM678mF96ipsSO0QvQXI4ib/7ZTxmzeJcY
N7bhvthFGminetBEWx+FI1R544GhRXTLun4zJl0pd7ha1RPvHQJ/UYbVtiUY
8vLd7n0eN2hufvwpT+Cc+dT0wS0UIK/ho0fBIBbZz8G/fkNl4D4cREZw59W/
oWgoCmx3kc2TAVkUAMip4RFmun6NM+wpbWLBt/gbdP7oGG8CG/bvVTeXghcH
TfmN04pGTRTVQmc/o1qRm3ij45K1tBvLzyz0/YdNWKGfAC29lmlcHLzsWK6m
DCRtQmPBY2JgbgANPSbg+qO2XzRbaJCB78HcZGCjWB53Jkaok80Ugt287zgY
hgYqi23W1OPCoUp6ACiKolpWEoZlkH9pPvSm+xObkb2v8rs2aP2k7AOMobCM
E9wjjpaGfjgORVRhPME9aaGJJEWVjUzu02xMCWWdarzxmCyOLQ1fpGpV9vWo
BfcpWQzQZCcNvu1d0N4Q+xnngUVnmqbJnlB2TOVLUxSJki0tKN2TnNkfLklx
T9hTyhL+B6hJNuzlxe9a2hLNw+wD5gpZvz9t/z59pTnZf0CPB8ItH8eYSGKN
uEp3bDW8cKUBTCIRXpA6KrZZK1LIEBhhTfF4prwzZTZ1ImDlTjeQgVIrp8Ks
+djmHUXf+GORlQco9CKZIYD61LIMX17YgytgFV0FTR12s1C9sy8AW196dKmi
04QA7ciiczkH+VYC2qsp7RgxQvCtnNTh6t4fNKqPzoMT9ZStLpgbmk2190Cl
lkMqpt+oVV8W/8KKRFJDSnUVJ5Zt8c1hhYN5kg2wjXAYVGVOoLFSK5MG2S4Q
SY9t2FwazgRK5AwUztpA7LsdrWxSGJZx5ed3oykBCeR8Hi9GzhWZqFx7fkXP
R5hd9jmRrrKDgxVgvhZbQVyLOq7Y/R0mk528cHSUv59yr9UlJWhlDt+Yto7K
N5Cje7AW0nG+IZpTeVF8/N+2gEQXMA5ibOkZmBq9KGWMLX4349R+5aANdDlb
yCUEjILlxnT8/rgZVQPxMxDNVrENRSHJkh5w827qwKbpKIgKZwhZqicgAIq5
9/LPfeVWRfmmQbw4xmqY2SstlqecTEHJEtVBysceYdVjaoJccFa3EBmJM9ri
W/9oZeTgPUqcxBWwkuEvLiW9MQZfiAgIrU3tZyId2h7Whr/Ky82QXcpJ1EEs
paz9/OmZg+ZoCBZLmbg82HA29XtI/YXJp4GT8h2ALZ1fQhKCor1ynvP6tLTz
bImP8Himwvgi1PdaACJrjOZgc/6xmaEa26HDWRlsI52+iCZ22vEYAYpYfyl+
ENig7lu5H+xDgz9wtbmxMaH+o+m+zcKsvjjMAla0552It3RsEuvK7h9iB/jV
UJ/IXhgvi4nP5Uvx05uT4VfZ+dQ9ze5eUYOFZ/CLQDW6WwcDN2BysOdKYYEw
ctGqs5Ktd7QsMUqNBOALzTwB4OEByTnMbriMljQD/YpLHCfpjJYAV0w+gYfJ
EFlSVjf4lJ+ySeDVy658vZ5ZWLdV5K7UfNnc9StKA9+KYE0sL2O/m7/sZ9pr
nA7JwnO+xS7iTr5gOIA28r+T3/AVc7tK0pez+fB/WuUOUxfxHZPadMr/ajui
AEoamrhbZ3KmkZLm9qYLQLV4qJ77m4Ls7E7UapSyNwekQB7GiURduXE3B7vv
czssS9szbzZ5rRGndkqm09UFG69/naDPFg2HhMtSVMAQeHeMxu8qvNkMNuwO
daZCDSsBZWAFpkLH3DCHTCuZRtUltnFME/k0sQaWrKeHSYHilwXtuPgklNf/
qLjAk78qlUjyy9qcHuJ4l4RGPU+XLgfMDJdJs/BSU4u5AefAQwmaeLw0KkIq
eJWJSmyia8UaTSFHshu8GyU+uJrMoNbDPYQrQxtpWm6FFPhNBWdFWJQmV1wf
FZgAEW8sp+guG3KejbOe+m38BP5m8Sa+PkFZAR/0cyrw5XIMInXYbTR27U4L
iRb7UD9zaGfeXU+57DVY0B9igrgdegPlhcfMeGYDO7vAAxY6Hg8bxJDsv/fZ
+SHNBg5o3XhLtHUrfaWKhi33lEUjuSRj9o+vhL/lb6qy86nt6qkVFe899z1y
VUS/+Q7uidStvHr5TuiEeKkNRXPDk0G7i4bM5kr9j2aVSg/Az/qqP5oP/PyO
48j9b8R0aBJ12ZnbUPx++IgQ8qAKqF14eHk9qOe9HRH17bi2EXcs/3uXR1M8
+vcyv6swachHXuSlyYXs5qxaNc6RmFEAgu0m4Yg0kTmR+Bsmae7aq6kn42e0
O3oFUdOYyJX8huWV4bAF8vNAqZbHUVgt6gMfBwmubPLGGBLXTpeHR9OcnhPl
dPejbY5riGy6oCwGQbDCh38jRBy+9Tve9RxGbtFHkim426+fbu3j9fh007tC
Li0VZBrM85QCStg+EOsn5sp+vM1g/OxdAdm/uIIhrWXcxcCRpiS1o4BDfhyc
Qv9KWRYO/qgt+F3cKgOW/+ZVuu4C/WzAWTaZkK5yAhiM+Wt6wjuAYdkGqH3U
Flfj5nklDblG4x303k6bJUeQp9HEAAJhaRuu83aGiMZYV7X6erSJeB9VRhnE
JTMhMuTpFsl0VhzfhiER32NXkJpYw7jIs2blLzhy/qPaaH1Sx2XSMN25N4XT
S5Iz4+cqZloU8ojboIOgkUMFrDwihP9VsUU3R7smuZIgXU4BwN5q0+vP8/w7
spDIZ58T/QUYQcDgd1KJrE/O97pAnSBjOgneL0xWBZ3PM2YKwKRnCiMTd7hx
9SvkzFFfSmt9wUVCceaccaHD0KSa21cm7++RyODutJdpU1NXBwDiBR2YP1od
qTlJ/KkMKMU40xcYeSgDgyuJOdnbuQr/+ZFw+oJ6MMTAgT2vNszA0bvTufBJ
OiGF69nugyEE490u/W7+wnOk/sO3lUCUnOR99zz/XkDeeAgN/H928A9I2Mnq
SVkolPnsESjdqcK8PEfY39jixFqS+mYByVYmI9BDqvRR89FmTjn058aguofC
/Li3sN8ll97Zg45GCcQEKL8+Lu6xEZSwdXvdlUwY1SlNEC6RXJuCfGnQEkLk
XaqZ9uSPKb8iimCZ2dSAO5yNGasWNo5ZFDjikCORIiz9rvwsIIkbt3KCRnyx
MW2d3qnjxmMOmFhQgTZad0LQyEJ/SkUqCT8WILthZ6L6h3oluJWagqSo7GK0
XhSXZO/TYIzKMOyamipf8Fh+PQEUFYwGcVU9FA01ElexzVepr4RP7UqCKtNq
7RsP/3dBJzIZ2jmCLRxxfnZnVpg8X4fVbeWeEXWHviq/fNxMgFavuX3f2iXb
X7aNHgx72WvsX+kmmZv8+Huut8ak+GCuoW6WebNV6/EVFJ85mHdm30ovURE8
+CUKXmLErFAkglwJCIfSz6iF3i5Xh09oEBvHBbCNQm030sS7sNFUdUes9s7J
iy1lHo4xbdZMrHGZl1JhrXIx1E/B9V6ZD2VvNAN0ArCpaHn5F5jt3D5bCD7W
hs7LUJWyuQmyxPJyHklmcc/PQ41Bo64CFQlwjxhY3Knkb4tO19A0J+XNWa3l
i7vT3xmWizw3R7/clP1vsY8zYjIXHfASR7jzo3PdmJqccXClAl4FEcX6s0Vm
eUZprQJcQryEZZlos+2dUP6f6v7/DNWBT8w5BClp6+WZQ6+3prPNQEPPfxqR
t6hc/lp1UvGxD0hTOP4khijFueXPR8hfjH6PZj0fLcKfCASCyr6z8635f4Yj
Sk9E90d/b3NJgoYQb9+0lFDRVIJvGWlBkfopgkHM2gGoqmj5R9gQIdCLJmFZ
kDy6R9YAvqizXzIPqWpmdnmYEHX/WOJS8krLUAW5S6xplpVOlcLZuLgQJe3+
qzajuAmlv/Ux/zfvq9Lw26GIaeUxGLJVgpSnAZQjaHsyDoKGSEFTlN7Y+sqS
EOHkGFSEe1CV+GDFvmt532YtcpuM7MhaRXTAmnmHRVKTFs2+DXpTIZd14f16
0eD68GB+9EggDYIvgF5iLBajNkFg9VCBLDsOJQe1Vg2djppX9gSf64sElJEa
4c6K8M27rNbXncFAlMeb8gdgWwH2U+A7k1tz3fIH0tziCr2mSCxn20qxwrZy
SOALZKUsiNuapHaZ8mZrJYD/YRGC+Mn01MSursrm9vZtfZVTy4q/V1mW2x2c
/kUfcoSk4tHlXAcVlIcFP9rh3syHsGN4bP46Vy0Zswk35idJTv/8hqZhWylY
MPnRhLmjt314Gm9SzeZ9cNOHJzhSflLqCf+ygq5LmAz5MoG1+GK8ES8TtQR6
iaJEdn0nicknZVnzEOZxBMvSM+DCa5pqdB80gVutU3MNF20cwTTRCiQjFgoK
Olex30CbkPf/BVlexm0yWA4okrYg4e6+lMMhA5mrMssgmR9MGC4Og0xoWbB0
rzYRCXrxH4EAQQ/3itBK32EnKx+GIvscdquZVhSFiHK3z3LwIRdyGHlSit2U
gY7m3aQFzt9ohQDCgUIwnziNRzuaEw8GOLAEevdatYXZv2s8V9TEuBVuUipA
yGf8E5aRDYFqZsI0YngHEvxDgqk3ZAMt/ovCC4Zs7goxdBSph6fEqb428zRw
CQAyv2CA3qaTXucfCmD9hw77yFqKWheHuZJnhU7vNTis2rLrkbyVnxzzMm7T
Iej0ThFWX/8dFkCRjsLa3pw/TsIklqWnoZJC8dXDhZvJUaAM1+tlrzDHIVX5
oaG/kXhv4AQLnUAUnPVoKcZHpGYh7vhwepLwtRVBtX7V0CpqealSwqx31GIh
bnROW+2uzrjpbjovGbGDzoCKpx6AMzgofIUIVDnbwlCPzq6NveE+0bnCCnlh
zYshw404Dw9Eff8UAjMkSvMdV6pS7facYeUizIaDjZnoIc7hOdI1CfzsreXS
NRF8yrHHqo8yf9AZKuYBOIhZygfTZp4ye/JHTe4FfA5cNDPJg4cvzypEIytz
hrZUf2Nu1gsuRVuVVyxZMRH6ETc2VN7C2U9mqyVHbVwQmC6vwPsHqxbpOTe2
5fKjnAHPI2dm1emDtNShFpEWPebYi9I/i/IRY09HzwL914deE8B7BFkLmiWm
2NzmdPI53vnhotYNDMn8Lp/IMCkbqgJr68VvKRxn7OsGSYIOUwO0LE/i+z2Z
qohf5A7tp6SN+I2DLYVADE87Xy4ZtlXxN+MADn1YeSuMzMAhzQxQCWGOTL3g
lheyI2Khv6KT+sHJjDi57hFiSwM3hovtWBJh3t9gRUW80S3s7jyo9VTRXWew
s1yj74m7dQPtTAaAssnUg7tTHcGb2K4OSUzpRSgUunw8lkh3FuU1rN1UXzoN
E5oWcA5Xl4+dwRUqrv3DZbSBg3fu/V/5vx4erzsl5ldtSJEIfBcxH6fX3PBd
6QLzqU4EPFNSjikBDDpdTUScDiEfp+nt8uSxUIxT6S3lBflyduaQTc3Q8bih
dZfYlEXn+1zsJ60RAzJ+L+toUIeVwzjZqREuskD0wUww0hCOGI3ryQXdk31o
WcIxPeTUaQnME7sAWhFld3Crq80r7bJJhvFxXHrSidBxjfAcxZT7JcJe5Ra6
Ffw8ojC3/+ycmyS8CAyMjksUFR2BiK+7LFKItiao/olxp9iKZhC7RxjIPPNK
HjOzweuBoHCrEtzjYd9hyHprRL0Th7zlTTXFaHyThwtUQUD9ChzZWN5ztvMx
wSlFdZdoa30HwkQBy+PUmjm0IjgbPHytwzb+wZF0JYehgtjVxvOV+xqYILee
/wnNnkDXShuDlHkGr1fYt71Wqm0W8kH0PUEDoY9xx2mZxl8imMYN0MBDOilK
4M58PLGpC1p5AyUGHW8CrhihYVUQVwp7Qf4XZa4mayndOe+L2Oaxn/4JBaDe
W4E3osMF4Kh1ECS+lnaWPNwGhNZcVymA4ScD7iDvPLKDtw1Tn8Jeu6CaA5H5
Z2xIIWJW5GrrAtWaqpa3pDmyEYDs3iQeN6GKxipmEiVlJvInp4wwIqiIS+Gt
5gETBi8ljrtiR3u6AatkkG8wl4QuQNPYHy75KrFTHphYdGpCH8nywVtavfdd
SEldkPQfcwRuzCbcF4CPeGNNC293x995TsYcUI2Ank7bAXYgYTHYkF97x5gm
vynKMIDfqHk2ID39y70S9Mm20iXHGVQp1UB2WFC1DTEVDCpRaJ/e8RrL+ws7
FxiCSVJLAz9Ii/pGSqFjgCO4pzQHgr8Iimk+O92PVBvO7sYr6jH6vXGmHBPD
H//yF8qac4Eenldkd7qQiL1Rugi6l1WNoJc3GjEMOj7pMzkak4cKa+G8urDJ
8y83jZ1SXF2EwPr2GUGWe589HBXwYavyt8IubAU4/H3+PZxky3vOtzlvP+M4
GpDju+pu7aq+FlCw65+C1pFMRYsQBM6mfQg0cVmXJNZsmxOTX2cBcsFQJmsV
NnbEjgLLN+/oQw9rK1s9kHsP6jQEqgqK88cnQgR1QDUKIXxJfM9KiHbzsG6T
eCPf0g6hmKGs+3V+zqS97UPcidRPmJ8qbmXVELZvgRhWtT2zG+0GwQkEjqK6
nvF0RrlkdRaBAYrvypwSoIKR6LeJAPkx9dpUXAQYCUDJIp4ypRLpWmWbgEZc
D2PWttSR2Tnf4ekO0zXic3W/uDbGIDOvX0bf70LZbzVw0e1ruhZo103epebb
/Jz7BQGYnrnCYf1gOXcOC0iw6tav5wXtQEXzmnFQYT2jshMgXOHnKae95qmT
dEPDALYUTKO9Iv4mJslRdVBIZlmXg173qtMvgds+8sM6NlCgYDZab1FMVPiZ
aBzllhEx6StTQ9gAssadHsHwWlSZ6pLiPCMGA3EbPXJTLkOMaoWr/eM5mCUq
HRBJLS8uHY8ZGB+e1Gho9bzjkq4qM0bnExJXslM+KAGhLm5nROUXxnc/gsdn
z7UvHOKmtz0JIqphUWmJsFJcPt88e2LksrrHcNcSJCk/sb+XgX7NvKwpgfsA
Ng+HY5Gwo5uF8z8osg0tKJ5WKANq89rzn8v0Q4sH8eq1jGglcdjLqAYgTryx
q/J83fN2ONpKhdkozEes6GMDyg6meqYOQ5w7rCKuSq6VpkLDIXZ4xtneDf5s
Faqx4APWu3dLhFj6Us2tTlYp4xpIWJ4ikU5g8AhmXx8esDxCglZ8KCUToSXy
/Bk7c2Gs9W/lDY08KxuPz1pzQb3de/iwSZ26W2l5A4/J3t7fWc525Z0jcb5F
zehSh8C5Nq/mgy4sCy3HYZDcTOEYQJCKOeQ/u3ZMh+UqkRwuYp+N4kn2lM4Q
zHXxeLfJpqQZ27I4cyGCovqBX7ccrVWTJAm3yIqAq7eIDLjMnUzHEhxZ28di
XzoVhOPg9be1g96pb1/CrMEQQh5pLgwqz7XJI7FF5UZ43MaozsJjT4v+le24
1C7WqT3rg/tAjsIl13EHhe8O9QFR5TJrc+e+lD/8TDZq7d0ZGNhGD5wmZixp
8ydh6J+wbzo6KIW+x5q4fflMjRNvnQEc6Ks4czXix3jbbjyU7/5ETvcDm9L5
Su+6xgFHYNmqg6K3AFsVoqRA4kocUUPOWLZuOnoSEHbMePwMaPwAx1Golm8j
3YBcnwuIX8USTIyEv3DqK6nzomVpM+midnvdquXHIfbvfMUvqQ81nUGUKyFH
AvH1XW3eSVvQLGecJcg5WoFJTTktQVKH6NsQohKi42FaqflB39H3fA5HR96K
e6n2In7w0PM3uLL6F8/Vu42cDcRHw7AxGzfH4FkOsrSN1GE4lRsX+GPbS3X0
vZMtf/3JOzU/ms1mkkBqb4lUYv7agaSILQIqoQZMYFB9kktOkymoOieu1mvI
i7Y4OnUPZ5KbKxuJTKYYUj9wm248R3RoVto/+D2owf5QanuCCsPfJ7gSl/v0
/XITtMigNFwVc4cdJPcmWknNSEvaYbn31hv+2examBuHRZlLj8WkO86ubNvl
UQGIBPtdNEyOia6wxEhG1P9UtQmawWXBXWuZjnGsX4hw5AA6O1ApHh37mRS7
rsNupV3vzioCmLomFGQMlRrAEk+erllIJJGcHMII4mxYAazudT8XWeKWiEo+
85WiQfOFjoNPbxhRBKlFYeOdKUQDki16yQK8f0yWIIB228TQrgU4xdxLfqPr
3YzbNd44ENqQv3sU4riG5QEM4ls+lgJy5UVJL6ZMdpuh9pjzgRVKEuNqaDiY
Gn3arEPj6DhEz5XQfJZtjrwdFJgoaAgKKBwY/TXVmV5VPynt4FrGYJ5YHoUp
Jhqf/XAYh67KrySj+9Gpu+K27KL4h+FRNfjTVt3WDwFqgbgKTERbkvs40CPr
BJr1rA2MROGiZlTb3/B2ORmZ48WIUDdZ52PC03/m3B91ROWCqwEX2QYve7S0
K2zeT8jgMpcmVFt7d2EMl+AslTKPa3k1CazjyN/WpP5xgCi4mPVpZdzyIgCv
S4KsGJlIhwUmUz1tC9/39cIfv3sWykm61oocs+eVWce/S8Z7sOFSW7BV2+yV
vzAMDKH2zd0OAffK/rla342Kfx4JIAOEKAkm3DMzR/jSJD4R32434G0eCyfW
+AKA533llxEdfxjJFjv5wF3SUUrfNK62z3ZA6lX4BVYN6RrpoO6LXgVtGTHo
TbuONBmakLVrXB+5afMNnRbQhORFDFM9UFwu8qcgfxlHdhw1w3mR1VGj1Sm0
EFS5tEEVLXZTDAM0ZxOmlT525FKq3OSGQ8sfvDq70NpKV/EO++m4BcS2DoZr
TswQlYzpUsGOcClQjpHaKTEAFg92ggss2muGOkIG17cz7jbWzZuMIyQXaRqH
+0A6lNpR41FKmWmrGUsmAg/SUPQTigeUuREwSgvvO2ialQJir8Pc0NV2cBFO
nlvy3a0gKmBnEgIRDRMgBdQqwUhncc7J0kEIvZGUEqBDdNXoZonGGqQS/S2f
cYo3+fRDLWF/jxEAPbEvm/oT0uw3h7BzJ/BvkcTsMvSvKxwG8/J98vA5WYhs
wkXswk0PthOT4RZeFLSXrc/2c31bC/8qcdaNpjf4LKj8U1RnsZk/nwmR/FA5
JBVBeI7PPA1YzgjDOzqI6HNGcUTGZCDhw/uGdfFcKLxcfB2e2PII1OX/R1SI
1l64aoaHwYPHnpYLhgqQsTZM0LkvsDpqGrlJqkk9Gp+UkNDsgG62FS9h2k6o
cd0CDnnV35u3seXLdwwzL3HW6TCIS6iVJePs4zxXceeMIwdx+kluhoxUypoU
WcFhzz+qA+ojx9QxM0BVyKKDoBph9QWcootn1TGe7vhHW1G36MWfLLtSV1Kp
RIxuPzXDmzxMpCYJ0xdwP9vtfpLy3pL9bqj65EZpI/1Z+htLC/Jdx4KJ1llf
Jm1tpSAAj+yyHvvMlsOiwzEME54DIg5PwcQpOTnV/et3pTbNnkFzBHjj8L5Q
HhzrbPbRYqAiBFn5am0CDWZGhtoPK+wD40u5hDE7lbo4pfAkoBvRyCdxE5g9
UklbThiCJl+kvhgp61gtvAEHcdpNH6xXpPKoE7SJWrqr3pDJGOCElAPnNluk
rZ/XjgcD11IEJfJmL0W7ec7z/943t6PKYiA7KUU5QJtNiZ0EuyrEzDRIPWSi
EJ9Oa8ZiFFro1MNWjeWh5BgwJwx5hP/PHeLGNL/T7/mpdVkQXJYVVrfTiUlm
0y2C71uXGUudNEGAcx5nI0HfhU3AYcPN64OylX7X2yEYeX9rYEGgX3WjquId
V8HemWg5KyQ+AVQPH4rhHz8ViK1tqZA4fsXnt1VrhWqq/fdgIaJ9htkPTSiE
NtNRNJ6Blb8EX/YBSD+2OymwC6CciR3m5n6x9jAuvgIZKs684U4hWjBvxIue
qbFfM7sA/CdfI+EUrK/jMoP/DJjb3AlORqoGNx2pp6BXuIrY1D2jlSXR52rC
suqPNF1IgU+c/XnVBXehkPbLoHgFThfQ/jRZiOcQFg8wZvGT9uOCuRqRdLHW
JxN4dPZrmEvnX/d31kKDlUiSgw898tZDpODJIbPF4p5yb3UlnG7kByiNmg7V
eeok/ZY6/hc8IOYn44RojXQV6RsYGFhG+54DbHAwvcoedMRvczHOMr4hRc21
3aF8yhBx2fxnTk/0N/EJtAB/tU9dw/vjHZF/YCDps8DDG9vjOQg0V06nRcWs
GsoA0wV2gkUsWNdW2XerIGt9C9MoxvbRB0Ar1VRrSB28IDpsKwTrlrSvfKIF
ZIc9Y2PprodX2MIvb+fLT7hUXPP+etYoQ3JBkaSxW3mMkTee5p0aeYyIqJ/P
/wQtKAuzLPJWjVK8nOwsQzVTZ6EQWQDmpXFESehJoMSMldjYmJXqHAfONqvS
fqsftqPKdlamC2mD+JcSapvR03Qwj/KvbrSlhu4NqgK6dhkeRdeE1UwAx5zr
GV807KIgMsuigSdeuFKHBGSZKL4y6u52SUrpJwLH9NovKaOwTgW2f8KE8Qwa
TLVW9lyPi4D+TDZCXrL5C//Jm7fW/yDoWD6CNIYlfQyFRlNCKvkzlM9rw73i
vOSk0cMm0feVjtJMjKBXGvKYaW/rHkF4i+BCEqtM4WYd4rWRKkMyufAAEtPF
scI+/fn+jnJdxZ38RBnY16fyRlPGKkMVMKDma3kdEb70b06vCR0AVAhQ1XVl
LpAaQFrVabfNESB2AIKd54EYb1D5BI+hTYrjgWsmn1VSxRmGKiZFrqZXOLnQ
NitPzOXPL4OBFlIUFyRABln1DYJZv8uVY6ZN/99IZkPS8nkbF749XemSBF5B
9oxM04E6UNdpSBCutlpydRy/uZyoAFBQEqPaGvcUeWJ2wGo4i7ULHdvIENPV
hAwR1SMpzCamdp8SulrehK6LqHZKE9fS3psY5j0VhNC4J+JdLCr9wXpxOPK7
WCLaGS3HtA2XgLFLHUL64mbFxcaUUVb1TLqrTNOoSx9IUlLgc+q6M/9GeaYV
yIjxsSgWBWze/jdzf15N8amXpRpvN8wBeNWw8/QgPVX+qKPbIUo/EMjCN56l
7AVg5RcPzJIFxjjy73GOFs2E4duzoYN1OIgBwma9MPCOQSnffPZgiLn+nJQC
Eoyu4azbZ0kEfMyzzYwma1eX9SdZyF9UlxQCLHdglnZEwbVV0pyMXnaY8yyQ
72Gmju0pESrpTWercjIaF8sSDrSwxqzpErmQHwEuTk/HOM1+JayliFDgxtgf
UmvYJItWWxS14ppI+UOZ9ngr5nlS0MGfyTv+RBJspNs317dc6t1bgSj7EpNo
/f5z3L7jHeV3FvjzZllM+BmDLS9JJJgR2SskbWweAu+G9cpn3bujp4rVwOZl
SGVc7IMdqEKRhPXTtzEQE0w5VZfupFDc/Fmu3XYqM5+NFWBHaBinZUw/aajW
8Kmac6MFvEM9Qe5E1UkQiXUwlwBZsKNC6cdECO20ISAfnL/+WWTa7K1M65eU
+pUqbnYyatVVPvVDHLwraOpHYSkIGBor3elTrbeQtdAESX4gSJllLDxM4whJ
D4wJNQzU7fV0lV0F3Tox31z4UWCXLVRBghGYotRM444su06TatEVbqcE1SXT
WYeIrTQeWGBeSa0nkpCn5LBKRgRyksw4GzGG+VXo7VHvkzpBRt4BcrzyFSDN
LUZCeiH415RTYncj66yFKXey2WO6/teEod+LwOHXf0i7IeRse9VOPywRDQ7L
DAJm01mkrylNcyh1U0cFO0phTIKv9bYQcqrs2S6DT1aV3uf5vXHhd7Qjcx1Q
xfE9mIHGrMTHry5hGjru/uPKOxzQxZ1KWHUOeGTwLTE13KCW1Wevh8op6cd9
Kv6Fs3QHaXKc+jQaCWlX4gzjqp1UsyXtSQM2ZMPTSm+I5aZ78AfkHcSYMuwj
IXby2msPKZN0GSdPAB6d/avHmtOhrIyHPyN8su0tf02VZTyhWbMfNnxKp94G
vH0enhhVeEDk3/kh5gRFsWipQcnSm5fQjN8CPMTDgZMmn30FjDCOBLxmRMCR
YKhhARwSEDdBtW7puxyzlc1CUA3EEubBkEsK3hwaifIrw2WvEmZffTZMZOiO
IfD4EIubfZ+d8i4kK5WGDBTnVbwElXLR+2BY3t5YP6N7mjQYV95YXe+fHZv7
yk3Z/b0M54hjWm7QCIluJED+8vYXBAIYZOqalWsrzQlde9RbqUNSC5Q0WCwK
6v4wpZG/6pKZedoDq3GWsEAuxGozGmXuYkqsSf43mJdPgsxjz+GZvtDrB/t3
45qKKaYdPuEW4BXBK8h2T0ZBibIUyO8P880TqQvELLI8XCsXP3O+R4jOtKJA
fDXcus5UlfeqtMVV9FcyzihAP0rQzfBCKP31G1nGgfnyF2Hc//pz7xC3r0Yf
9L3wtlzBsn0AF63sC7Mu6CbewMl5p84XaiqhZe0EpK8Ckf7DZ5puKVxWO6TE
6MjA/GFbZfBZ15S3zgXbcMh1/7ap/Lt0Bnd1ryuOCgso11ZNRm1/UNNYYrGw
zGY7bkiuEuVI8jxn7AgsSUDmuqvwlUH54hGt/eTMtSm+JhOUm92LpNdT4YTy
R9W4kuQvBIbdgkL5DCQbmrgJojPBzk6Ujwe1vI4KdY8siKf7Mm3IORZBBbY1
ucvyWSs1bhRmCHCunM4lFGC+KfmJWCH6KUx87KoSYpWCfMe/pPTk1AbOE4Re
7D6FrGI2+YFDSz6go8qrw1pH4BTsbYzMsHCKJDegx0TsSMtHukMzWT/E1dmo
PaQreybBQPdG6KqfCwWcBotK6Nqkw/cydp7Rm7eM6sqi0YJ4UqR7EvYOtvTf
oTvE3+zK9ZDQ9qoZKDD5rrsI+jDvxQTurNP4nqeKMG65rGfp75zEwIv7DZiZ
F9WH6pWFZamif03aZdxhcm5thIxD8iMUIBEwNY2LHtZTIukvktYM4nPJlkR5
VlM7OvWEvPkIKhZfzxIldPOPyiqC8EaOVpWQHxp/iwmMS4pvU+ORbzF9IiOV
VnQ0hIrHKO1inaS12h2km77+5WBywLNOY52c5q6/LAPvj9o4SxYV/wNjpO44
NOBze7VvMY2tQ8HZ1Ra6NHfKgHBL3k+bfLUWymBsiuMZUYkQ/qAp73KwVTvA
o0FtENkTTO3ltQE3Ytcb4MiHmQB7F3Gfz29iaXMSRCkeosHbX2bW5K1DDnzv
RqYWom0w5oUUSCyYvx7I5zqiVaNjpFKDALaZWzTZ9L2LZ5udwOlMmrrm66Jx
h87l8bZHwascbYDAEiWo2vkBAs7XGFlFllUKh/nq/Ypek/ZyXZjnZIeo1dRS
UfXn8y9fO7+MPvF8c8brI3VuPonqh1dJcGDZUoJcCBD8O1vU6x+AViOiVkKg
C9M43HO/KC78KXV730yRtYG3M4dqTJb32+z/kYyxICjrAhN0nDHFBviWwJtC
/eo1e40c+trwiGL/MfhqhhsDU6XdWycjgKw97z8ySEOAv9FNF1ODY48c+nwh
HIWpe3PSWKpDpD/jYdvysEaEDQnu9dYEc21wfLsoimb2BqrIcalifZCBp92D
l3BvzK4/P9vb9/+RQPkh10jGy7D4an2z2ITUAR0wacP3kxxxa+xIdaLYAFV3
lCMBAMpQK9g6HUVPEmI8PAy7kVEp+qYra340IlDYCw8X39AkDL7okgmOl0tU
73KWvW0w6XVitRlZp6ILtiX34+2xC3wyfmeh0iWh6PuaEzi0txdmCra526TR
MicaG9O8goiCXJS7C9zNJ77RUjiaFiOhmSUsEsLuy+1n0bO5eZ17f+eebz6r
/yvKeHEf6ZOSKPXqm6iHTx4d2FuqmyUHML9tkCjyNV+uRXA+OeiBIbvMph3P
/JNmlcEcHtSdv3cFg1KNFVY+DdO29Uf8R4Ie9Oxk2ycwQeA/rrzfQPADQPJ4
hunao1zawBSRgvrLoy7CIQlyTlTrHleA2VCH887JEXNiSClbG53WJSMICpwL
8VYt5CnwyhUDEiQ0dqXXGCEE2YWJtTa/f1+lA+axcZeqHQsb5Vs0wg1c0nKX
Y7E0HT59PhEXY9xmfxCYyLDh69QFH6DwTjsiFK7U9CeaSgNLDwqbWc5JK3NS
Sufo6FXEv/jSEU01dUgQ1bSk7sHBgXZf57kF5vrVa/r4q1DAIIUT1QJrehD2
vfR5wXvci+HtX5raPuGyrFT4dWmXL5NxX7WMyvJSFC61IzYdsdT/MVxZc4om
5R8jUbvgLw4atIe+Une7UErX/Nzp4s2HttG+H/xD4zi+qCAwz7yEu0EYKp6N
WYaohKRHCC7di8oiybjb4E4LurSiT0Sx2wXYlhVa1i+MD3K3SJNQetgMWOnP
bxfmHmijFKf+fqgCbv6qjVJb7SNXQFELcYC0TWDUmsKristD888w3bmDCNn2
s3Em1LzaWCxtNUkCkrsMcnbd1q1NTGRYnrOzazXt7y+8ZHGXo0AHP0Zb7qEj
jWp+8LsEUlw9xJSm21RDv0QT5ooNoLyMw+DVGcIK04PaUkpdD6NGPO2nW8Px
k3qbT2NMg0aTU9Zk7Q3Xm2gYMNMAuJK+UD50mV8alvIyFsY4+fiaeWGWKomT
z2brSj2mRw7nzNW/zcglqszmOfYQFXCAGVZ2UWNyvh+ysdH2mnm7SbQbXF3L
pOh0YgQc+1RYlYNMfV8JcBlYz6ao86pPbYmFjWhPEnHADFPeDrfbUdBq05rY
RqkNGWtxKaU3AJPYwSXwEXtUj2fe3TaVqe39WYi0TjgGK2iRGrkdnHPPpYho
EMmqHn5+6WzJm6IB+A/0Gw29s+VO2sAzTOre0+eFGK4F5CKqS1UhVD7pNxv7
blw2xf0f2ns3hx0ZWbitQrcLhEekm5YEglrICVThjniwwLHnTpwBJ1F6NpDn
1it5lLSUn3InTWSfYdj+sAjux2Bt4c9XMZfkdkvhZxwZR/fEsOtkz+Wtbnna
1rr4/I+BzhKVSHDOFxAuPjY1DhGOaxh64uBi40Z9O55FLsb8BOdImaiWZkP8
9KP4oueuCT7rmnJHuPVjm9SypDSkK4ahLJRj6dV7cUdjxluIqk7YzZkGnlrU
ydy7R5EOyw8cajRnz8DCE4v/ZYcQccSbKNvz0wMxuBcS4cgPCwyHnBGj1+xc
ebtcT8blaUpIPRaAu36ELNPgsvDWlxvjxE+TYKgfdptxVBrMaWkXY956C7kJ
LWCFVkUm9v+CmbdQo4kZr7LQN6iAmZdYeyMli/w5gDL4kccnoDiHXQtM8BO6
J6jnD8MY1Q4gFC2OgPToH+wAhJF+N+K8bGneYUI52DXJVVyboKesQ0TrH6cY
V9ZQT5BwthWm976g8Iy8CKvCyb9zbI8dLlh/fREHBvyuL4hYw8qmCZJLpng+
kEkWmeBH4ugP46/NYKfQROyFaJikUwcCVCb28V6sWgMKQ33r+M4pGhGIlC2u
dYR9ZbRuqIf/TuL9WKT1nHJm3BlU6hQ+Ag1Ck/LVyGnHhd443LqB9bltLvQC
l6JCa7Detrx9uAqLsE5k+3e9UWCR0lAlID4vXHgPd4igOen+Kqk4gxvb6Zjh
eNoooQZ6Ds59Y24/mPCkPJORkHEbdzzS04kdEgWaJiMRwuyueZIFNqhDqJ24
iCzL/57R0EYZk9bl8ibmn0OdnrJvJRkAgqWA9/xOltcpyQRLIeZRLpKNuzw5
sbmVlQAuiIvpHT0NvUKwqzAtY7cLpB7hTbokr5WQH3hCfSmJM6WJOow1xjwx
uU9mN6c63yu6uciNHHSoSljW5Y2EoHp9sZwqCsnHJRQyuk9IFLh48slqIES6
UlaYiA04NK6wa3fzYO2shVfBIWpSKc8dcixh85lMxFHDFcXECN8VWJVz10/z
n96tqPTduQr1Btegqd5/p3OW8aVZ16CZ8GLHMU93eoHqtVyz0Y0TdHRd9H4X
nwDrW4RCUYCkbTasgrdx57hquW27j2tcs93H29VChZC5an4BHdZhZ2NkPmvw
e0tTomUfpmB7cMEBwgpcybkDYHUH8KlSpDm6u7vjwkm8wWkGNhPKO/GsRNBy
TBSPN4ufIucr4QaOrZhhoKN4d14fsFVOg8L/jHIOzRZ7WCPvT26rE03Ci2vR
ZZPE6tdAZ31DaDECfiPbyIP+BboqdM2KCN3t0AD3H4V8F7YHiYK778Ih3uR7
1JwkDOZVbGsytlr3FrcI2j6F6J9gbI2PL33kUKDWsmRgGeKDTf0rnAzLxZrC
3qRUhB3rrX4Fh/UaYxqktFliF8YOQpVHvfESxZ4zKLWeGPPsEJ47XFYQerfg
P7L0Wgvj9D8xdps7hHJHGXOu5dk4tCieGpwMwR1V5kw13zp8g10kGxqYFJOg
M8eag7CKku+tnKMuzOqc0eq40Smx2bk+UGfcE6a877voWSuQ2zFLSlM4DrWu
pfzrr9WdqZ60LEUYIKecRCxpUZqAhO14L9/SIVMQgD1EzLMBvMPUD8Ewm1kG
D+qt5je2Jy2KNSxOrc8htzOE0W4m9EzHSw0Eg40ts3K2sVxFoUNxTzNCXvAs
PGt7XoVyj5QOTCS8y/5Nhq9ylj5Dj7tUggqIs7tMWpRkmMEKWXjEVM/PecRh
Kn3xFFF+hL8ypE1m/LTGzYjKmfizMC6mLbjncIY9tf7cpUFDKubJrHX2MNFT
ORG6kxttOPbl7Xowo0cgUjvO3jwIOEwN394gutGXMCaPKiqYw1UXUHmK+Xdr
4sq5GBoCfKqg5xQ6fXLDL1VF9twaSPiU1W7NJB53x6S27+RwtUOw7yOj5lon
SbNJ1cmkLUEc3FEQV0ar5rUGVWie6OBMl76z5loY4PyBnVTKbXu2iXODc8t8
Ta80kQ4okZgLrjLNkLByrRU39lsHy+ZFEA5MRNCo4GOVy/44KyNS5ChvWXje
7BfdBhB8dYTuhlI85sdsadewy8acKM9WrfOFn6/VYSn9X6KPyJM4Vd8kad72
3AUzBQbarQ8OkbY74XZ1GFY//hWCyYXSs8seCOr9XgcTdcJWO+omXAISq8fC
c4M+g7NW0MMv17dx/ObumX94vjTcjVFsKAU0G2B85qeRvEdgftwv7DgRoZnX
aTcjnFR+roxABQt/tNCPzNL/2fR1uyNTD1nWvVjn2rEfO5+fDAzAunNj3MLs
x75f/QS3/vFyONdFWibGeecKsL9J0MS1UrN9v25U3lZYPZBHBsFd2kEDY9Oo
GxwolhkIw9xxPsnzBbbF3IiO+al7Evsv+uSFeq5siT80auwaQvVVDSCJKPRd
iYsZxj5x3JC1G3SeL6CDBuFsJeTdCSihipR8oeXi1lcl9xzLtAWEuNMxTA20
N8TiA3pOKHryEJ9q5tUiyVtDzUZclNugaZDdr09VTYd4ZpzWH2ChpGhvymB8
O5FyEvheUPYaa3cRV0/4WcMPgBPLDVIv8Q9rAj+TpBvnGkxMIi3OgJvgWh+C
5qF+pd464ModbPiFtLfaVHO2g3XDqYWU1xbOBK8yN0jaL+wSyoSzQg+koX8J
8TUQeouH6TJPsXC6Lu4NCidJkOGeOlFRTqygibftkgUzJolkwQy5kI05Fqaz
7XrJWI4GICMEO3OV9DvrQIrjkrV+zHJPLcKo4st8fF0iYMtqBUbTuSnri1yA
KkY97JNu3HJgj+mX38qfzEi0LOj2zLVmPfk+cp8YRwZzKHyXc4XZso+fmmdG
TWCJ63otEt6gpHZ+b9xOnBgQIQ8R+rkEOFnaC663Y/Jezj2AUgxyoC5OiLhY
npwWlEEVU9LqXMvfcdJOeZMh38edLHKBrI7+YZkehWZFCpXhKCxPHxPVvoWQ
QMPqTghCmm67PplIcbnKwEihiIDHNc+CiOQ8cmbJyip2WmP80v3FBNVaOO9B
5ttlNxdR1JSt+hNZKU4dVtzoZGf1JgOHlHc7FcWsSlB8Zofx9gJjUINyOnuu
zff3wO5f2YXjUxuFA5CQIZ+DDz7PDSIjycT1mb7Sro+GjzlrtE3/FfUJKr7z
KttYHdpcSSEXRLWRAuQDxVbcJCkLWw32D9bEfpPIFcZAw5Iv0aMSWLDjDE/Z
pN054g5bEHLkWYMGkLTZTjqrECanbYdhDl5UIOa35KvYWKYUFXTdJ1XfqkJR
mvU/7K8hRWPK0ahQla22WUiqgXncQ+owqeVYob77b0USWOH+pq+n60yUI8Ez
OkLFL7KyHE3X23yIywnlw6qoITnnWDptCql7NVmRdPxfX191M1GUBvDVY4wr
uKmADdRgH/lvE0NhxAFlhmROrkq6nZ3TKZ0lfdaahed1xcp7gKKJR7LadkpO
oiKPCeNtSQqKj7uG/8Yd4dMu29hu5+2huVc39cy9aLVLNZ6fBBJJDKZah9H9
5fBjIKE0xm98LPRbjDwbJYuZMme2orE5PkSTZR//XZby0ff2bU750AhKwKl3
hxSsFRn7o7f08W72UOzdRJr35Rufr7bpcRsKROG0P9j2jRu1V/GXk2YAOFj1
NJlk8u7t84IxW3zzQv9/ZxWyExWcRM+qeTotWpOX2MJX6b2jUZEy2mqFBm6p
IuHaOe9mneCfWXW0d3c+/ZVSPvvfzaLax66U3NyLNvZbbHMdfVvSXiZDK69U
ebs1qydDi9a8AbtMnQp75Ku5i3R5xrzBouOg15eKsCiB9HBu8JDrVl8SBK3R
BkeMfwH2Y4myhe9PYRUqln1EXDkr2Pdnk1cdQ1MnH0yiO6S3UzVDVsmGB5Lx
wB6e7MQWAGTytOHnlEGvK7bVd/3l+5PgeUErRIvRRLqv73hMf92hLGGNBWBa
YHoYoZ8nRaBe/Gsun27+6A8egaMyL8or+vp0DEVnQSYjI9LsBfnYzOHDNag3
rs5bw8kugzxiv3x63pXYAjJQFalcm72ucpYjLSIkwqqeZpaC1tZ8ahBFxqBL
eSf2mFWEqhUHcySsemPZmjNg6VIqEs18+Ia7e+3q6z7v11zCyBV8ADA9IADv
+MJf8C5jqNVIcFKI0skLTKkZ2a6D/G6Ie4/pJA4sscWG1eF5YFL9srs3FoH8
RUtoF3XkbDgr4JUAr4Xpbdh03PU+lNEmQwemJ4tBvFlMDFGH22ERqjYgDaNS
dCGdkYqTVQUjpI4vDjekRrTRn+pyuyR70/AdBneOWis95qysqH5iqA6yAzeS
aRYExhc1556btPZIo2IFL3uJXmUsutNtawhPZeQzwcsHc7i5d6MAyDb10/M2
nyYd9WR14rtP7RBykQ5q5io0CTs8GiOsPpwsj2/2TqEB/OUQQz/OnpFvN7UV
f/zKD6aT+8yJVWLN/qHcifx7DIinahKJEIGy/K6XJ+ge8Q13iw4dqVhz7eQA
whx+o+kFekRTqpjE2QbhlqyMUin5hXskEIzawDmYLq54J/UV3sMpiH/wDWh/
P6etFWLtOx4LhytbtR2b9Q4c3WO+XCXGXE1rbHpt/X+JQtgfgCUZpkzghedU
8D+wC+WX1e+CXlozbuEyuMImaog3u9urg9h8QaJcQ97w4JiNIgQAPVSrO1lX
9WASGZkINBxYcpvv/qsLmp52DIAAIfQb7dcEH6vNEH6WIYJpSMGk5muBu33m
+O9/Qkv8hsx6QVlzRwlyBIpOo0FCd9VGDUbtr9ae9Qzaz3/8Fw4UZb1T02NH
Unse3nD8E1VThl2rk9x2xSGPjOjDRM6mavlXh7cCBDDHcfexWePPudsF18X1
tgg3VeIAPOBHsDzSLoTfqXgrCjHQpmTWEzRKus1DmAarH51yDEulJ08xJYCQ
6dz3+25UFG+Ms0hU1NJEeYs79LOaar8S2qmb/Fiw691G7VOH1IG8PvYpiL6n
fxJhruP4IlAGQF8tcNvJoAZK/gKwbh7MQ1rjwqe++nKRoeHXg9cvLuRouRMV
8TRCbVtnzkir+xGS+pBDlgVgFayyrARsUy9Uf58bP/AOaBbcGAe+wjmEXNKZ
8KSGqmVRCZWoUWBubFdK+1zS11LcwXEAoLc+44+3zwc2TqbHQIZ/PcXsJ4EB
qRJqad23hkXOGvS4LwGAY1Ju4QVlzvUUmenmkkb/6tHF+7vqNfUVCMycffkz
XAcxidNPy9AExpAEQP6/OcUjxETFfqU6kmTcUN3jO/KFQst578MMMHnXiiaI
MJjWtL0k6qz4rOBJLzyEX/WJx/STvo8H76u3ickjzbwiz6KqyjqCfwQfxnT7
n09Rn5mDWdVPrkGItQoc05/Fa158WEUrlGLcjFhaOVVc2GFABH047llcwH0i
fU8nOj3WY+8cgBrWHLkkB8DU9m8jbQXfHOwg9f3g95TMmXrgPnCLU6dazTL6
F8LQLgQh2yvq2aS6ki06jzUNyTlSUjmE6Iq0LVs4T8LcjaODR5fxjYsaeYP0
w3Papjc2MjQ7eGIcoYjQGOtlo99clDrVUbh36UyWqKPt7CFczbN9dq4SBtZq
cTb4oRnZj62TiQxLHQxHmi/MCGrEfaEo0LdYR/F/EM94ejjoNOQ0yg1e7IPO
14NCds27vBmvALK+sqa0jJXnn3vXuCFo6c63bcPJArDp877sCEbEz1nW9x1H
X7bsR2URcn4D1kb7a9sl+fpkayTIM72YcMRdQMZX1Q5XNRYQEp2sm65i5Y1/
p34EQGArE6Rql4NR+oNQJ/BbwXRFqcawgF3fAxvkD9l1Z+oyFxqvOm4AHXSY
okZzjEK9/1R6OXlze6+05uLaFArC3UepC9JooiwVh29ffAupn8Uc/noJIX5j
rqi2aGckM4P+59bqfIlfpdVRa1d+91J91sqCFxPgXWptA6Fi3Y5u1tPbrPPG
BGmDJcwFqzP625MxAPOwcv5+LPfEV9jf6I/YCl92sT0ymfRifwG4ZIfEp2jg
MFTWmDOaIO0FPhBt3rxQwXgdd0Kgio3kvvtLaJJiHFhY+GGmVxOJlZk5lzhz
punrFBhDw0O0UnsHYuq2fB/cgtiUENVcXW/QrXIrh5lPMOz0L+dvU2MskUrR
u2fkjOgGW9A5OvUxH5Q40dlMmQ5a+r44RtXnSJGKkZ6+zaXNHND4WI3y4wjs
yjKo9xJxvpldlXCwWV7lb8luPEnZBl6D78DNydr+GADC4R8og97n/TIibzGz
ARN2MXSgUUmMFftXf+UAlEmv6AwoKgX81lEfYiYkalTWmsG/uxCwab3As5w5
sEiTwyG+Tr2X04uTNlPdTVjA6gKA40jdEajYYW8rwWBoD1561A8IsbLAF/qP
Zvzy7PvlFGzwbbetDsAfw/3WFiQiGRROAF71eHv8YbHueMeo9oXQefXkXiYm
ENTptQLMIS2GQbMozXAzrrW2UVCckLhecganvTEgjNjmv7X/lS8T4NGBCguP
yuL0TWlImUB3WBoog/IMM0OIFSRO66RSIITN2wgKXzeZ9RVFdDNsjlOXBk0F
klJKE5LxArsO8qe074lmRetBw0OCWi/LypvhDVFwaJ0nr3s9THU58O69c6vt
eUlMoTcOon2sRCUriyRSeUhdaW8EFPbyfUEHQDMo/xgGbQ1nEUK83RA3gApc
4c81OI5Nq8vy8DlDAz2ah+dd276F+ANo4vdVYivx1NIBT5pmCF8luy40crEX
3z202aWS/CxZYa5xVmZUrd8jjNInX56/T3fFgjKQCKga7bpnfirGdHXUdFSd
7fFwBNqIaNdGDB1eS9w6HYXD2jEvcjwEkwdb58u1lsilUxWZ0+X8Nky1XiVl
RGls7F5aWVbnq0yrlC/JvnEz139zI2HAs+hMzZC/POfftkn6129/e9LIEKy7
caChnXmCv5DEfa/ueMZqOsvFlYF7Em6J+5Yl5fDEsVc6EiyZ9bRDbXG1LlSI
Fc+NQ5/RzpOy/8ZfbgviDogvywBLXThJuC3NDmxSx18v2AUcXtYGbUYecIwC
RX2ear4kDQJSCYP4WX9eAgjj3g9i3RFTUmGWncZxROPs58dhQcYpNCc74eN8
pIbwFlxA4JNs62Xvpo+Lmvba9rI5ulKW/uHd6aDtm1YwV2cVHwgD8t7FMRcF
HDYEnOntyMRndAJ7OEdNTr/0yqJKPJmBPnotD8w/I64kOrwUBII9igA2d0uW
e+MAEIED9+3Rv3wKOgosVZYtYMS4G2F8OPNdS/j0+vmlQvDUyKVY7PyHbRqi
aYPDcmH4wJW6+ODUEGRdkQNz7AZTtGhj89B18pK7D9EU+QQnhvc49PSOKjOj
jvxL8HgVd7QRaNffnx4bccSn6PPSdpirHx4O5sRXzMNU/wfiY7z67d89Yy0k
wx6MbcK2P65SX0m1LLYS3LdI1VRAj9Zk3IOqQdb0oerAvY8FndgdtT9CKxVG
ARN0FPi2TwR8hI824RxYzJk/Iarhtu6/ZP4tBdSD6iZO4ZFSDk0664jw3Hj+
jcPTNz6Uc2kisOlVimVLJGWTwCEBpXmE81nz374bgnsxCfhg5RudiuZAKjth
24s3ecFY65OImTRi6++HL0vvtVH3uk5eRkAyMmltAPucnP4gfI+Eqv/Z6hYY
lyrYFVQtn9UGHP4ZV/DqBBjyDgkz5ztns6Zqp2q8BH1vZg9qem69XnV8LqS0
zq0Wy11yr5USjzCyuUgqbsh1V/0qwU0DqASK9b3xP1QVhBcCvZrJekzLwnc7
iiuQ9xYRjdRXGjApUkQwj7YKSSsmJWX7gMp+QNZVwYloLPGcF8vF1f+9Ujzk
W1+ffdjAVlZb0k6GvYJhPY3hW//uAXXI6DXUXK8eWpEJf2SOe5lz3WbmWQ2k
bZ/h637lS7rNO1tRCd+xihwkZidUL2Hqu+FAxKjRDWWmYNQgoO50I507ocTq
huvckKr6NlJ2cP769fT7GHSRdd29PmaCU/yB4sG4Etz6wzZFYxaIKnvEqX/2
xM+2+kZIZSnCBXBjrQGDLmPBfDFWaOeKalC2wM2wNBDHFZDx8N+BnapUu8/e
brhu3wi16BmDUnSxJnd/tXO4GKPnZq/2nZxb5qNp/jOWi13/Z3dbHnfo+Ybj
xFlmafRbtf2uSP8Ra78sI3QC9KGRxJckm++aLI/XXl5BSugBBGX/23dG/0ZA
GV9TGqTEis5AO97UFDb8My5ikf8qq2Chbc2q3lFTROlNTB36miWi0T2VcN+U
lvS3+mxZ2FGHuHCqS/9KSixMJ0n3wliSvqmfrmwuaGQqZ60yWwHBLcM1T3Xb
6i3Qy/qIvio5fSrhoCJsIUvkWa5NYRiwZCghFYnVpBILDBrFWJK1mHiv0Y8C
Ja9ZJ6aArf8wY8ImeeA2efZEQJyRPhPcblYcS4ksuta8xqOMu/wee6yHvWDA
ZhI4tlq92LFzOud6qIkGa4fMJMI3vAUW2FYfDH7HxAu1sAOGZhx0WwS7GFaD
JjPXcVY5XZlft100ADTOvbrlA1E+g5FeJ82DlqsT4Y7p9phWS+h0hIPd5jR4
PJ0Ol19GMWNnV8Hnp5zyCUwEV4lfQH+x8Qtqhbjs9H1n9cHSZrD/tTg6uSCV
x2Cs7fvvkceyw7wcm6Ooopn/BeBpmRtpF8qIdWpEWOn12cVgeq6gNFoSTkaL
Sht3c2tLpKeGmq11ATrBswOIL9qZe2h6fhozceGYur2EZiPRAuAf61yPudNa
+QyLc0Fb40BDusyEwZaKUt6E+bCQJo1yr2PNArN28k3dJUekIf03LnwvN7S/
dZmxZrcyuURbMvy/lcA4cTjiXKtlvZIfin5DoaRKcAyBvRO0ms+wzUMp5/E1
UGwbMLfb0+eEnKTkJdX8yM7Wa2XbsDF62EiFDf7nC4R1F+E4CIVNB8r9zl/1
UBfwkthHg02HWAiL/6wI7ALRwE9/KZzgGa+q6nFOMkX8Hv3FiuMcrMm7my44
oTIWQiv9kw/xwjDfgC7r93lzMU0sUf0VL/nroXLu6/e7YsKzJxuJCuKjs/ZG
rfjLwv/7DOuVC2P3f5qgWl3Cn7H2WQGd0/wE7minbnRbEJJRXKvfaycP3qjn
7IS7E1DGWLFx1z2WYhJxyGklxIQnlPpzBCwqAdQ/KIMYnle/09qc2SaiAjCP
7ixtDN1Mw8k/a16Qz934DS6tc4kbUDPy7PaYQ5J1ch31MDxAAfHjGR5bYa/7
z3bv4iI4KKwXoshtnAB2dxiRKwdRKf2s3mFnKc+c0fp/RSjACWQbQSZMDxmE
4D929imY/+4ArmLiaTfht8c2H98ZntHoivEVNCNXyeFbDWuH+JMq32eDf7Tp
yBaZRDOn8eK6asxedrYJicKYvbz3BgLAk+d5SrPFqbwxx8dhRUrLiQ8hE1Hr
j5YM7rDJaUU4W+2vzbTi+vW5s7V4iaurQQ4U/+i8StEbGXqx6wRExruV0zdB
qcU9UdcwrOmeKgkd0tggpvmV3em6IECdm1EDDS5wQkqt/iiBpsPKCpnz+QYJ
13ACPOihE+8y6n1A7yfCSgoadoivr4Ap0v5WvgPRV+hBulpJ4bH9lJGlUDDh
cyOoeiqiEA+zUNhvmJINsmqKQC1OxWL/YgRacB4sOgTYNWZwNKxYz5mpmP3Y
yfnBvseF9LmVLCSo4WaSYmog0Sp1apD6V+nLTfL1cHLcINdtgqTkufpuFzXq
0aMcgxt1MwXyjoljZfAgH/Y3vqroecU+9fp9JW6L5842wmfuFwvW5KiNG+KD
vbIU7XVEmrADPFb0IpLaHLGthiCEuuQvIG54RPsqzwShSQQ11Qrpn6C3e0lZ
4LJ+rzWcLBfySSFe1l0jzg1MnNyiaF7k3AImiVQ4iv87y265pAeguU53fk57
bPCT4umuKiiaz61vh4YAjMvsWVCvjBrsxfu6HM3Td7i+YefvUNvxvRg/EwAh
4HvKMcqwFPTr4awVuygGD6/RYfOEZh0ULyvL8nA3+fdE1lToFEuT9sCCOhfP
gOPFJfuit3ve+hnTeCXX5P7a2TT0Ly70wF2FcX2L3G3dEch52LnUqE9UW373
SJ5DBHwYF+bWJOpDPArTSqw+JnB0JwuxcdzbPfgWKoAm758bHiPbKBgj+Jcq
DVhLbafN2BRHcBbZwxkm7bPQEw4oWifCi7po+6rtzleZY4UYRtESlKq+OnrG
ZwOe2bOekE/gGpcp38HQPE2ypKp7vhc+Ep7U6Ffz6vDVgBzPuIv7VV+ZrPrN
lrQYHeRySVeOJy3byBapAf5OlBn29CH0OJ1Ic1odtumq0twnGRrhcfFnUmkP
VFB4PgK3QPXZykfmPy8m6zJ6FoHPlylK0yjTSHxC1Ojt+0a1LKccsdnrDuvY
70Zys6t0MqLCXDIWNanC4LsRG8XyqjUMC81olSQvrbSrPkpQqpVYX7hAz57s
Q4nFKSwPx08GRN3Vcs8NcQL70YiwNCJU1VSNwgu67de9X6xffI3ZCXtB3Pzo
Wrg6JTqoUTJ3/NBzZFSu+v5Jk/zXrXAXk+uLCn26IOdPdtSRlU1ox3oxJ2Od
/Rw13pVvnaVAh/CXttVAVR2z+RyJL9FzvciTOJyFYFwPqjXduT5nmIgcICQV
2qKXKx5qr+nVda5mlbdunYnlX2fK1LQxpqRznV0De7Z7ksielPG6v7J4ajGq
Po94CSVf6ElSo8hZi2Z46LCmnNW1aMp/QrmwkBhsMyj5XzqlDs2MtkWE7xXk
JbgIRS3QYpprp27RjUYIKMXoszdccDB0MdIjTHIONkJ+U/tNNARjGVtJ9I8x
ec1YNMz+Dkzebsf1/Bugs7Kb2cxuylcYGubZ2zBJVqCW2fwz7yWVBf8l/P8n
ozVIf/ppeLjnK8TWAD2Es7S7FgA4xqGcsm6ECpYj48WgM0CFxLTgKxpiPHic
Nxlt3fsb/RrnP8GNYtVJd6RKTTdx2+048gOrUtjVTvEqyzXvHD4q5OVhV7ma
Unsol4VF+KH9LOQnH1ybGUu8DRf/PwPYYsdJ5p78ascLqdmBldzfEVWyi9oP
AlFydFKnvouUzyvKOAEh9UiQT4cmwMQBbjzcG+BlIapdiJEtIIUX6cMOFkNy
sLIUzZJLuHF4GveJdFWVgZYRJm6aTUJ6btfHcmvNTGLclFtv5m6qmtBQN7rx
p+OCTxozhVh11katWOBpPI024qEm/DANbd9zs5sIbDYd2VtiWT26Cf6wDD1l
QML0/L5stSFii7mJ6V15IFJ09Ii4vd9YNUxpdK5H0vRwSGe1MBeoVrxb2a3K
AiG6RS3wxEgIDpFK5BH0EFC8QEWgUQZU6tUpRSkO4Gt9CpLMlBiqkCxhmlPB
N8gl27b9bXqoYngh9oIzMvK3G03AV2Z34G++o/BoM5CpprEHIznSLlpOus9H
/vwQIsbLhkdoet1ZC0eCoc95tpamVSkKFNI8B3NgWByHNy4qswgee/UaM9ib
xkcogm98Q4bQfeb/4DRwK3FMFg+Qv9q486sPSTmRJzQLR1BdkgOzdbZtrtmJ
eNn/bfm+xRkBXzoFysW39jNmTqsFvVgT0JkeVlvhy/tqc8+ibrmkdU2VMh89
njHXmw4QUhZhwH2bEycqm13h3jXKm9iAFAHMciOXV/fX3Ql5BEoo+jOcyLuF
iUTQ7TyjPnt7FgJdH4V+6l3hChuAglT/7SdJ0qqqkusBdvfrgK1Eb/sEp1qD
kbhUFY1BRiT0QB9sOYSlOsEtWw+C38wmYyO07q4ARL1oYGZV31X1FAaaIv9O
Q+UZXbRwZWJwHuVDGXXMNnatvyI87kYfV97/UIIXp+LSr3XRgbwQB5TU4SF1
gwzSGJep/ygwQeNwTMFoImEfRDZczK/Sndv3JXXIzWZIRldH78OkryM4NWEf
dgEflLxvlBzu8oJFZNiif6icywdbil8HRpkAe9v/0ZZZK1S9YL+GfhT/LErp
Vx6dTFNJaklpRYxaI3JxAsXUuBPUM1XeGoWgIrQE7LL3QvjyAWtGzCni187T
3bRIikF5fv07zXLLHbCfdz1BtkCUUQpeI6uBJ4rY8KtNoe8OPIC5fX6kmnKQ
z5m8C1zXRTWx/oYhWhlbB3rVTx0r7WXgGsG852nISQ8/HDj04hZJMJO7GhrB
mwdKgs4KE2UAaUbWamFruUaWgGg4uf0BFoPRCle+4lZeYxoRgh/dkBbQsGYi
lNkvmnxXy8XepjWNdHD6oeEGEg+Bn5/+9I+lS04oppTIvgA5CVoIM0ie18MB
oBo/E8WnoYwSC3aksViVTjeuEhM0GlxRfgCtHqq4aQrrh0pNzzryHg/6EGI+
A5KRYrOUadtwkODW+OD0nEUbixPPvcfC+ogdhC/AwGurcS3A8eRnjVXEOANK
eEpaGHUnmrkSOG0Jnu8bWZhh0xDLXG7AWBSSBDu/xfEvEjQf62KcF1wHrCc6
QGsl5R7vVrnEY1RaNbGAE5e7qmHFZHkBmVd79kSjo8d92DxuKpu4/PzuPGKg
/ogDMRxAHAGbW852HfNCfAktyAb5Djib7hHtY1rWzK3n9s2uNpTbWypPMgGc
8munmiZn1DxfihkiA9V6KrZTGJ8C+gG+CjOPA2scsdMuMxd3i8m+G3l4Fyru
+f7a3fyeGicbut2vcShDiqz64N7u419N8qjLVmeHP9O0UMmomF5atheDrVjI
vzjeK3wcmQoulhvWjNSP/2U0hR15AcYTtSKQ/0OGtLEQ/gVww0sD/hrfX29V
PQ6FZ2lxi2ntCzfnGUAhdZwIM+TWdtAiMd/izKr6/+/E/3/5rITkg3bq+p3V
ltBT9vH2vZo+HTy2EoLXg+bsyILmRxtIS3Wzf4F2x6ekUs/ENFuc/V1HRrS3
NOM9hPOzW9kp1ClBdWc3X9i6nLvwiwnh6tze/j64NDnUGH4emXpgx8oxKtJx
R8oMiD1YVWz9WwImskIdeFJ2F8OwB6NbO4IpZV9dxlzZQFGSSCwp/Pc4yJQz
GnAvnSg8jFwnMaxeuQ9cGcHccLS3/xYML5t7Hx8vuRjRDsvMs9pd7UpEHVm4
/WJ5qKAgineJkKP/SodRnWgsN8wL4IPnaERmIAJAz9lpIZnkJ/Jq4aWgEtPA
iLH7GB3APE1XYSKm4KvtONaOK9q7f8i0M7plFCCuzmF6aBJiWPKeFgjCjEWD
gv2XpWSQH5lQEnr6nc6uium5GJxGtFOQ2VfU9rNHga8qPgadeaEruLX3VciH
FBX3HkHsODFioWnJtxdbL2bbM561Cttgn6OJqbjt2AGZa4B63+CkcrJToCG6
gA6O+HDSaM/mJwrnbtlMEAgwHO+P9zTE3MIPTN9vxrhMaTqp4spXJgV5R0zd
SFPvVfKZn85OdEwyf81qFLjhLAgNm65xzCn+mJ+QZ8OQiElQym979PooEccD
cpELjIUHE3Bx7ATQ05TSb2StMLMRWHNAMPpBn8x/Lt18Hmn9x7LtccJDKdQG
HemyuTXZOeRy7SUaQZeLB5h7Zlf52T9T2c6G0wA34rlVfMLLP9LZLgwY6X04
DLQPUE6lVFly4zRRnpqfmAL+sjfcfg3qXqoJeO2AKTZxXMRw6rnB91eBdKa4
X3NcEytymlH85S44E24Xe+IIHFOIdqjyt+P8I/ikAcQ+QbbzeF4QTuL0cSxG
hhi0jdDQBiojrhSD9Ql0FkNGosAzRaGzr3Ppv+X5pCExYqMTb84J0cPcJuxq
Y84rSZuNAJ0v78fkuCMqcE89fLvpjzOXJqeVF7wLx8wn0JwqWWafOA9R3ErK
7koYUBg4HkVgSanS30HNRP9M8ZmlNbcW9fNetbWlwaiifdJMs4+7clAjv8ub
I47Hok/vpcQFRyKKVgIeWlD0waZKymGfvsjdc1d9DPMytA3bORLGyM9SnqjE
ePY+2/TKFR1beRbjiVArmwVi8IHvbXb2N4Ezi0iASGxeq2r+40Mvx1vXO6UL
OewHlUq1zf/86xQHK0+9YDdRHyQXezj5Xz21Zpdbo1eV2AXi2IGAKj7Xz4S7
RZeA44dV0Gsr2k3pGB8ixj9hRc1hslGBlIrr6xE6s+UEbVFb2xOJMCu2pK3o
nNyNIWc2GoIuFchgt4T4bJfLEdtm+NuDpUnUHvQsMbBqUhGWKp5p8LGql8qI
IR5awM3WycaUw4wfNVvIC+svudklgBDb30J3v2Y26aAFy2dk0IF3UWplut3c
3zR44QHn9HPnI8fZDZPgBdhueI3ZsaQWLsBDW9+E3dK2TH9A8f5aWw3f2F2h
mxWZsl/1JQ+WLFk7XmC29B5PHeqwLZGODzZj9Gk2FV0CQCKmvxCDEGircObU
wS+M3nlfrHJOSaBAZ49JUmIruP+Nwym0eK8dIwAQ3KivFHZRgJo/UaAtY1VL
A5am/TCjLmCILyw06eTHbJuGQkiIPXaHi3veI+Iy1XDs3RnRz7j5G4aky0Xp
sfjj0HL5N0TPIKzyLrEF7/KOtlFRpW90D7f1z36ecblivUibLzAFmFcOpDuX
iAZrhdJZbraFrbJ5tHKE2cDSGA2BplBQNt3au01NlDOSVg3Z5Iw6wMArzJwC
J+iMvK+YJstQzGJW/v2DxSOMnQv6e5RPOsNsVeV05gx/hfSh4VK2voq3KIg7
gH8gyJ69q65DfAwHzh8xcFRlrVdi9FM/P+qq1DqDL2bjlSqNDYhzYPfY/wvP
D/VNpRfX2FM9IYBkG2r4CLjktaAuYYUhUCXZX8wFDxRMcGA7JdXP3JC8aUL5
wUTj4c/Vtu+R3tlTNA3kO5qfQvBh4U41p6xfrDiCuviMhQaP+m5Fk78OK4JZ
r7VXyFgIo+mT3/zPGkkwCfx6ZUoD5+mdbvBejWkNXhulW3Tvz3TDeIdAQ8tD
+EveLvHz5wBknQfaGQvJQMZSLL3fmDNSET6k2RjeUP9WW/W3u5kQidZWNkfy
xa5QuUn+zsOFRvM1U9g8iQr4l0YGy1+tsukdpd8jBpVV3h2FV6BYzRJXZUXi
0bTlmQg7lWZz8y/2iIEEHlQGdgrpZBP0Je4VpTim1jdi+vwb+YpownWlbT6k
b6a1VxOdnmLSDVbrAUNgNXQ9LUDX91Frf4ENWM06aPQdTrGXKew8SZI4az9z
k6QbXLSfEvtBZGBv74hIbu3rQR5gEK6KUaq7pWNKaKc/CDZiDv4av4XDpBeq
cVodyDcIE5s3cKMnRNsvGyz41aABpVk0gGwiqp4jq/dDCwP9yMQe/fpWNPrn
3K83/eJmVJc5mxLlavbC9Y9blgqtKypL7Z0HmuG07jKG85xpvJSS7AiUpfeE
yz6yjgNgMlbceSduqZGSzfzyVd4KOibvMBY3Y1I8fhEueA1H8ubKP2krFill
3n3SPtUL42XJcFOmkLlwBvqN80GxkBXxco5YTVB7AgquJyGU1QWXbAG7Pzyn
F26FW87AQSiQVMfa0rHd0JKux+uLDs5q+MC032vhfGJqLdcl0sEXPdjI1PvO
gFTxVaInazoIDWC4lLS6hO9Z34uRzIA7pCu5pOF+uV4XZED8SrWzE3YCXL65
9t8xEs6Si+zletYWalQjKO6HQwla9UL9C43HjauV6Q7ASAtQXFYiz8xYN8EH
16TQVbcxrLe/vOe/ZJiWhgWkcRBUEyRUyN5hfUo0FgzSR7eobI9S2JbYX5QP
y+5jW3KVXdqYlTgLbhgVCX1SxS9eUsamdoGnCWo+aRR8wA6wUfcxcxz5ZicV
Pf09Y6G9ld+0QIU7Z0uhhFXfhZxDKRHpy8Z+JlBLzMIQGlG0YYNdX7lyWXgO
RrXOLf+PiFEMAV+1xmH6pEElF65wJG614nmIw9TYlG9X4SELzvjNNYi7peSn
/R0fRzmWzGXAYlXf1qLm5TH//i0Yo0MIy8f4HwxX2gPad/jVUGEA8nghqVRC
xo5TcABtM9YdyeEzaeQY0nNWySqqypTP8Yb3iMvk3AZRdy9xuD02qSOGwPb1
+xTCIT4TNsO4t3Js/wKsdw3UOKNd+B9nP5LhrwvW06S0wdzFaTrfEqfZkrIQ
ApxQrP9odj7LRaJ25bDpX74ipTtT8x0vhIn07+p2gXmvwCLSflMJZxJlxQRE
ic8+9eFyrntNbck0vEmXzonFgB/4A2/Q/balSQwZ+/G6bDypSnd8RCiKdB8l
QuPpAzA4cjeZmhlhNLXo/KD2argHcvda3T/c9scsLqujDrvlGPRGqQO2Fxor
/RtBL9cFdKzyGxjYNOeBsHcqGgAwr8/WFrKxnRxiWkbPMlVXyiUgDsuCAZci
hajJIqlI6mrv81ld6K8PQVOP+yedOnuQhDQDEzSn0ezWlGE55IBvsYlWnu4T
HNRTeQpBGcVFdc2+k6F+Dzqzyx6PIX3w1lydcaqB+srVoSL5Fl1rmj44/sBj
Sroqgvh0EkNeM9+vRIsvjeiIyu8VVv0sYKdsZlPN8CrlVjEvZiCbwQNuQkoF
fuY5qls6YvrIVkYTXZnVmJqYw4rCktCtbnLLXLaTzXaw/ZOjXejcm/Xr1+du
7dR7jwdZuw5fq8jilsmbGEG+hEaWcq2JVIk9z9mz7fb76pXPdz3QMvQUS0/i
F/kRCKziTWr1a1AyiW7KLyLcHbvMoewjXguXNp00Qd2t1ZiDVNX37XjiHYkm
DytmjG/wqN/Fe9et2QK7M8k2VIe3aal+renbXnqByX+lHIO0nUPao/VdVboz
rOsaLr6Jv2lz9MN0TZ4wFVbnM1eQIyeNajTqcMpXqCzYVHd1woS+zu5rXulY
t3kfggQ3fJN6bfJjtcAgV+cOb93jVy7RpjV54chNvEYZt5quxTxvb+E3yg7K
ggX7E5OsVUC+lSIOhlZ5G74IJGbi50KiVKCehA7kQ5J3kD4ff2Z7Ld3bXB7+
qAeI5hzBFY9zhib7jPoXTUgrXJ35ttb7BhfN9nCtqnlTkenUXJQwbw7WdYEA
bcyMZs7jZUJiFWE06EFiwPFXqnoYUq+D8f3CghPo6oq+zbVon6Z+1nyJzrvU
tjLuMnZZHh9Si7dzaGgattlRjpMXZnTrAsJR3IYkFuUtGxqo/bSaq/VuJa96
pdO420+Zpislmt88waOM5gG7ZpXlGWQFBnxMdHVM8XgXzLkOs41sJ48MhZ3w
AYz3wp690Z47t07dqwCitGpRWptDBR8QsHBPEaf57fvf//4BMWMsFD8t41i0
gtSATpwqONamf69C/GfBUNqE1Kakfs6GB/z8uPR06P0o9a2VJNyV/35q1FwI
NOzgGOlEcmY1DIwHRjRCypZ5nGXzCyNnWArl+GVGtha4YK1oOCgCBasOOH7g
ymetaBvadWLnkAQjuq1K9OfHKhjyELq9wBWwLkUSP3NVOWeLvZz5wqOR5I1w
LZy8nOdLQzEKiaSgjwCsv5H4PNcF21rvkq+/B8ljYm+H/jbqXxoG9JS4PHfQ
EDEL2rNu12YkXnAYEXxYLg/9frRWdmf6HjGJQ4gMvSfPpXieoVA/m6zZEfOE
bsxybNedBBAVv4/QNVGC2qyNa5b4QR6ZyaT/l8eJ9bYBfzkOwB2f/sSH5p/Y
AgaxmDwl+y6iVKv5Byn4SuhiNWpQlhVFirk7ty6x+sMmz8ygGjddbaRJpPsa
VpjrTdPU7sEglafQPIsQ6EZj5bkpSX7T+oLFRjEM1cXSjA8/mh35FQQfIqKB
4gGV7XujZNlv62gYc/YcZLWHhaOw2s+rtx6m7slqlP0bpgQ3PT15Cis/DdA9
7Hp/i+0BnBIDdoeXBhXV8cMZXOpj16ppxyz+EX088IaqxbtBqPpkW8o1DekE
lqG0T5JL3pxiqS27sUUZ117HI1xO4sVFIILQzSBIzvMt+1/dOr1JCfbygQIq
Kt0NS3GM+MFIMLoGTVxOQClIb7ISMnZ5eW+LuZf36ReMK92hnrsbKTvUExPP
ERrWc0Q3rW0FC3WQDfMpHZnBxI/Ku4oaBpS4Rcc2B7C+YKvuUbjsGvVDD8cP
XNn2JivyuxzEurkS5k53+JEH9eoU10cX0yLxS7YCJ6LBR/12j8er2wfAqENn
rs8C5nQsJgPonKH49r/edZMJIdYhJtCUhr6JQuZ5cXkSwOCfpjKJfovVvaEq
W0DCm2XKZFyGpca9g/cCmMDkAUASZPx3Y9mwHmTOQfg66X4dxm69NbypFXfm
cBwwI1f+qH3z7OnZNno4l4TzkkD3e99JwRHnzYV9gbTN5zfyK3NJUY1C2rJs
+IxYv5T3G9+81HI8g/2Pw/6XOfMkEmzMPe4I/t9YQw/KIapgqFPbykiAdvoc
F60VNGRLzLmiT1yGFZJpQyLQwao+OwDCW14yBIbLyKP2qrO4kU808kPwLkCF
PqFyik4HH5Q/LWdVL3Exj52Lpm9BCv1OVvDxZ6odx5pDV4MO/4Wh0uhfkymb
X1JSqpgg5SCEkEDSQGejerxj8rAq9bSxQb8X5V5I+ylNDalg3srp765EwuQs
BjBBQMm4vwQTu0/2dnW4EhAwj4wweaQBsT5yoE5+RAn5uhH9fxBZcNbSXDGG
DE84wvEA/85PaGz6szeJnF8Ts5OmTScsr8KwRbeMpPHp7HcWf6dUbVlV2/gO
fmU6DcKfq+jUWiRIfgpYlR1jdMrir9e+VNU4oBMDa5UaBCDTQH50G2Oj2cKs
8FtxIF9ixgaGh4pRTNV8Gl1rZpJ+euc8R9CNK5dv3lD7qKfLKL932N4q37uk
9qbP1x/cvUH9zbibtrtM2bYKSokbCoUo7oVTf5+JWcUU3kIS174OPggiGj2f
W5QaNmBl/C7CIl01MS3ScP5qVyqgaB9rOphx1S0kKZUmgAylL2qa78Tvck0h
sVSW0eYpNLOljuN6EuOpUNy/+8LXru12geYBtj450/SwnKC7JVSekeXDE/IY
tJsLCUnQJEWCTHfALXB/ClJ89GjrfekqLur3dsnog5YKOQya1IIkfFDLQn4S
mX+3ctWUPAfP2Utk54sguv9WTBrAz6esLetFuZ45qNkoBZ7LYVAAtxyq7NS9
LqUJm4S2nT34tiPtOv/xCmb6x255sb0/S6mT8uYGjU8mN7O8asdtRSFsgXF7
GsubTxX6reKN+R463EzN02q4+8dXT2E2RPH/2eaCncdITXDeQO7O8Jzxbz6c
Ysxg/M0Ur6N0ajOk1wSwwFbSpqJ/OE08am0SzEkuysD/QJTjAs6PlhQW+OtY
uvKzAyZhu6cGFOHlc1guYdiGJU/XHX6uVYAk/R+Xhzzp+Xu27+eHwXK928W1
ubGnP2/bAMbhLLy07yVdBoAfQcyZJan1xYFFKV5/TNq3C/Nh0LEpe347IJil
dhH5M9N1fpCCQptI57CNq5N8g9CGwt3llTwU1F5U0sJlCHBGlT1psVv6jW9V
vq5EqqpPLPBtMZAVhxEI0GnIfb3atitLePOnxkbp0fhXzsFV3ifqNXxGbxfj
IVIOOQeqMD6kk2p3jkkPlE4416uQPTTug9pVXbQH2/sY4oo9VXztea1P7Cui
hye87H697guOrBTOakmzw+yKQF/kDPu9fl0Ix12fpEFv+5CwCw5EwSIpCCJ3
E+Da7uzWEc8OZqItABI973RoAqEtdBhQHSB+RrLaJ/D4LdMYKzOyUBhkhsWx
cAfmEMWRaVB8a8uF+v3kGSRiR1MHc3FBAa0cBez0GR9XBelZ3z1kSXryp2ia
W/UTvgg0jTFelG3BwfV9V2Eu4ROGX1dbV6z5QKLhUxuXMs/IkYwLYmXmgV52
VRddynSZY7XFzLCIO4VjwO2nWedbwng323k9lHVO1kKyslbuxhBU2EOtuyw/
ZUhXNWzqdzaqjTh/t7qp3YDvRR5AaPyCTwNiscOC/8IqljFCgMUY8C97pSkX
sU/guk2x8Kf3cEPoG+mjEk8mXaNlIdvIZfr+IfMbA0IF4OaovrmQM1XvosVl
VQ4/t2Fd5n08bBYugDkZc14GxgRE9TM9PkTezZSIO946Q7GBrPVfWAUVT2Wz
7DCcgGr5WbaMMn6IHKzp86bmhOD8ibwucpC3nwd1ERe+QIHJaKZr/bOIy0Bv
MTkk+ZDjHRaXU/c9LmU67OW2z6C0BQPyXbFvRIxBsOY8viEukRBuf81GwyCg
hUxGkOjdPHSb6xvqjIbodeJ4ooIc0paqtp2477mz0H5MV0b/GwjxXYPr2LWN
a00+4//wg01vl4Xll4XJWgJSlttMTHCRgcVvnS9IdPswdHYCZ8IHjb9LWuc1
Gs/jD3F0OxI90Mt7vp4xhh8CHZfdP9oCGSnUkONSmCY+YeDJOKaiqbl/DrKx
Mo2Qr5vaiWE+Mc9FiO/T5/Ig5tqTKgNi24eF/BYsw7Y4fI9k3gU0hIDQlBVc
9BF/CphFTedQ70pQH1i6esd1SDqBwE9BZbqMrVqQI1erzypKeYfxqEnMy4et
fxY62ujq7JoWConpNZH/m5rmsHlVrbhk0gf41Ai65P2P6qfNsgPrlKrEOQfj
BK7pWIIN1h4+og8sHO5hVDAOWRPbjCIdDFwr8WuUCJtfg01scM1bGVLFgNFM
H8wPva0vfkxSUm0WVrBW3X6vSvgEWxvRCxJKMZQfpGOKu3HjqEKcWC7Q799J
RIgQpmmn3miB/HALYYY/uRMfaFuZM4DZjKnFj94xONe39rwbdBufOD0qUQzt
W5j332IrTen2lzEeaoEVoLbzw+IYiPsnyy6xTntdpy3Lh2f9PKCW77gQ4w48
r1PS1vviZkwGFomWWbed1wJ9lfD75vSpp9NmgSpZ01B2yzbe0PZOh6FwwOtM
olEqxCoHJ6SjsEkI+yfjyM3ZqwXzGw4gmKbyR88lAqmMbySomu/91TQBhHNy
BH6tk2wgQPfXYwmHuvRTvm1XxUaS0WzJjTPiTa2Hf6JorpitqgarwQEaFBBQ
K5e3ktYTvzJGpeNQwhYKc3MPNQuRRDf+yWCdj4gDo1hq6PsI0jUePrLxc+oD
SsnTX+n+wbIGQT72UtHEHkkuZpWHtOvU5c9BJVVASCO83OLSUBYx9i786jMK
E4Z0V+5K3dJY8AEnNqmZEcQ7G+f/0besFwRuWXj8aTiqWrMaQ3+1Psn1qa8a
PFFxquaeH0rgYzTHO7apPjJdz67yJ4R1qqK9cPHLRby3vxQxJJ3EwR1JAm7K
BsUTnE93lf+ME0ykvEXtr93TEuvFYHWpB9PIXPmAaN3/QtLnGQDKJAyXhYEV
O9ipN/YsBBUUMjalkt55PRUWzMVlGBx06bKIdBrEgbANptw3rANnNazMYcyq
adokQ8IF7okDVtgr1um8bxjlIN8MFgaAs/WtXr5mbEtvS1TE4cugO9c4TXY3
jZKM+AqA813p75W1ili61uPoyRp8NwAgVp8wN2yn94/jDKfKFuLCdicBUsgC
qczBQqB5f3oBXnmlGrC8Ubl8BmHLwQwVrS8pob3Q2q5Wa1X0vbROYXeRBPex
Mqm0qzmGQmDi5W2BBJpaeGOLtJVGXgLrJViOmKkLbl/wgIUQnLZp2EYawNEd
KgDY/kCcDIorghKPodRv6XsM+s8ZHda1xcrY/01To9DGfCzNibW9++AUkuBK
UTDoDlm3YyB6rNw0wvs/rgbjU9c+ob7zu1Ov4dvE84YAlGZuQgC1CgzlYaUU
Q81lgkCYzZ1EDBysl3NwkTU7AxMF6HGL29FMAus1avjTfU9v0Me8ta96i+Zx
0JLIWXDU3erYjZ2PEmLGhd8eEBB4+pktriopx9q2QtEDwubZ3Qc5/aqXjQmq
fqKEB9l5g3rwrs8o95O4t3AuBwfpx9X7Q65q3DD88F45LTNeNQ7Nsoa9jQix
SvsT74sfzTrEiFqipAOd4DJjTWbUABfDgQo3u3hi/13Li67sFGXjNbjEAsVl
+FrIuDGxFBbTA2Z6VEc0hb9VfzTU/0DhRTHkcv1yP1AESp/eCUGWMtfb/Zde
U73faaT4Rnq2AJ4IApq0gFqOBspeoObKsJGEdU2csDlk/ZJxxl4pIPENKQUC
G+wXH65ANn3SGoGzmGdlg9UoI9hggh39IOwbMlRaiJb3MPX9u7oeUvpD2FvV
3T9Glz80rcBDY2FEL+IXtnXHyU5OGD4vNoikh+0jr3Z2ACIxTQIiXWMJ08ru
FLs9+Vv9sZl+kBztHtQG8151RTvgn5QUQ1yGpW/6p3NVuFBQrRDKDfi5WAP6
WQieBVydCOXirpZDUBKETRWR0M2ILvZVZ4gEHCn127mBfpZTjLtWRp/EUHXu
Kuw3H8REUC+ZLvDTVzWGSvH6QJuKdJtq1qldaoi8kki1xsGelMCYXp7Iyymj
209wYv/cBhs0FWt2o1a4seU2LNBXwe3cJ1O6Ge5GVGTqVRlurp0sxF+OfW1k
P66Pjbnqy7yAsA0ASfWmG94AHvtj8cVuOgnOPbVQAdep2SeXMN1us964yok3
cSvSaI1Nul+5yYAG7a5GEEcBhOb9DuU8rgjz9UPFOzjL7WLq0R5NWEQWW8GE
Yweo1AKlIe8AoAPT2mNM8zpwxXDoiQHa1l213qAaAG8Pd7A54Egw1F+zmdoE
GdJ1cw6pE8t6u9mNvCnwQfibXu2HdsMCzJi7LQ7mVff9D5ltwlH2lCGcVG4X
Oph2fzNZGf1GswIArexLrIr2PrgDztSP2ZpYuobzyiuPEjCEqOHEUj0mHOG8
is5Y19327oseEHkkLFTouQHhonzXnndFbYamV8HZ5wyTootzSgphFHrBnr6/
oDgTmc3W3h0JvSYHgSl5Kl5kWhiV1Pg37lTohze1HplahKj5QRAvibceJ2Xw
d5TYs5Qj6d7gCqzxmo9uZwBkrQswhM6fmTxnu665TXU2neS4s+eQXrSNsvOq
fpX4ydlyA0nCwy3e9Qc+MSXM3wtht7x10i2Yxe57SyaXKDUvHdWsNdZ/fu/b
F9rZp+x5ZKBj5Q8VNxMCL3+ZqEhsl8wbo5PxRwk7t1F7lQBW+fRuKHD2ABLg
FjpeV/avQHWHg5KeN4hHb3u4vVAVBvKn7KtnD0VquqohFa2kTLFMk5G/rBmw
cpwrd9UM5Hyo+FzQ4ExhDMiVGssixbAFWW/H/2CTclY1ahn78L9n6NuwBHjL
ICbeT8sWKSiTxetHArI5JMPXEypuanubQNXgxxuQy/az89IDwYRTw2LHA/kg
W/Jw4EKXBH/EZpC+lq9Xg60bKbMn1tSMOClcEcK+AzWxrG5j5LPjZs0kGFpk
LkVPSwIKmzeK7fVS+1RneEapUXrztNCHXvWpLbmTWe6yfaEZ+MTIlsxAjzxu
bmVQmLt4JZ9goUFTMgUdu1ONNEgSljh5KekOKOqzUntBU4LAwUI+UeHLERon
dvE4f78er3yKCm+A5ESr4j3Aw4r2EaO6GWzGHPl4Jt1Xp0eTC5SuOwhgv3Ph
XCCgVUN63ISTfvKmOw9P9/Q5yzR9nKUTHNvQrJ0102hXRcyQHPYJ+2sm5pNS
OQkRrFAfJhsYFNLKAxc92HumTRS1aNxqvKBhg8mwMNiU18Cn94xnZj3MaNCx
jaH5HAKHlQFUVNNxt4EaHDtkhQ+RUBmPcUIFvT0S/X+xCcSDpPQlsQpux4Em
MXuuz6fwgJlWrp5Dm/KxhMnzG94jsngcR4QvvL5Onlq0VPf5jHfdNrcH1uSl
PuXmkXkZpfIYxo0h5J1YYJUCNDFKmzavx6ANKLkxCJr4o/GAVxR/6TKa2477
U/Bfoc7EUjSmX8zmZ7QEIv87a9zDTKTu/bMryxW9CCX+n+l0M+Kd3UI1rN4Z
6kZrE+IDQLK1AA+dzWph2+sdiDRykx3maJ2J7rMyUALW/flvwdYAXS40dbBr
Cr03lnZCJA8VqTKX4rk/RIPwEsqZBPxX7BFw3/557ALQ1KtgbKISWP2iBJhP
KJ8j0qYSClvBdL0dhJauNRhLo+NnuRSAOIOWJxpAWsnU1rbsQ0HfxhDhtmOD
LreZzZGaGobg9LtQWcbFYjuA2iwIo/ie9Hb4SQwrr8oigt+hoj1ScfGi+Rzm
DKbldpcTcrVjgz+tITy8gv0szbrBAiafdNYZhu3v9aUOA7xyS4vyLsieDQsD
B+Y7iu2FqOt8ERWWJKDX/cTBq3BSDIeLlozsLniKJ2pWVxDzmPx4kfj+FeSF
AU/tERhKzlXD3XxarI5y6uQu8TligoIDbbRXNjyctRv4BUa7Kc0VV3dkzQ2D
eYhInXLxXZMujwyauYKFqtdMdYHP4hFrxSG0ES5ntz2m6rKhZK9aowJyQm/6
7QKBh7Ti3zSalWWmxPgU0DFMio61gZq3JSO2W0bkb9cblHY53dnxzoBLV1E1
7kqkUS3TuBxQasb/i3s6HLzWI1erdQfF/MsctBl3wE59MyGAHqbkMdxxapRF
r6OpT0R1sC9V9QT5P9ZB9xk0KKspT/cl8+xNSO9ds8nxHX8oHWGceLueNs6r
LIW+zE30NEgZdS5+4c8GV+74pB79/tEqeAuQTfjgqtJ1/tlq/zewbgwqlT6H
MBvEYWRNrlxgvnVWm93j8JNojATpZBtboZIyR+YlwrZIg49xfYLY/f2CMax+
oSeiCMkVv7dFbwG3Zg8owySK9GAHY0HccjuSl1OVggrOeaW92cVJC0+ytAHu
J9lkkvsEqNqT4FqyQ5Qg8rN1ugVC+4XyYTVcLi2/4zJeBL+4rk1mikyKMwev
KV+0MXdPc1BY9+mboENWLpuZjNRejfN5DhdW9lfmjr6pchtJqNH2KELlzfpt
hZdlI7sdSmbWn7JO7rG8mxSRgY2KbLwBfvANsmG//CTNpXuIM4lYIgkMOeRc
nsUflV/OrVJ72DiTLDAAL2S0WPO0IORGY8Rm+3cX4ntnv4iIY8Vxwoy2ruKF
fSealTJqVf6HkaBzhUptfvEwEEPIUIWtdSogtQZR4YKU6CgUhQsb6ou+dnik
3owgC6I/xJbk72m9iNhLqbmpF/qpv3Gg68p0oVYdWEe8tdI4btaFb5HEruxv
RqGuNEv4nugHeeVLWiZvFKbAkJjhUQcqXduCcg5oZiTunF7ObPFeSafpeeW1
MWeHgqVdL3jMG4IY2hAxPwr167ZR8cpWB/PaG6nf8erht0JliDHx1PxJD0EW
FZncDCc/o6UQOqNztIu+Nk5jW9zVpT7cnp3DOIVCg5zWVpuV4fze6O4a7ngK
GHmHd7yA9uE80yJ3rrQ3JBY9GDHH0CPO/jrxA5/ZeKRQdDZLBxWv6e3atV6C
3ztg53xkr7GTUiIbe4XRzEHMDVFTfPY81ScKc3rvvuyLwUZgWx7dNOBllLhb
ehKf8ee9d3MIDSi3vrSKtLLrZOOKGP77mhQJ5cejMer+BqCCVDyF7X9ArhoK
zfVy53MOuJBJwnal/rQ1DAEi1mfI32pX5RMH3Js0Y8/QvbHSRbPZzBVa6izR
Sppz/2lQc2EhwQpcWXyW9t8GWd2mG1mp2yf00rjfEOT4aYgQLuH4og9yGFCf
4SBKSSkcWd0qi+M1aRsmjFbut8aLxpN+B65zlVM7w5S35S3sJ/tykvMC9EZO
C4Tb3d3Vt/dt2aID0bSDbMVbDhnR2+UTMVcR/2P9LNZbqnsE/xxB7ZkfI9j4
JS5E/nkG5mUHvrlLRfaRkB34s/VKQ29psb7tUy0ZN/U6gBf9Jqaknr74JDkL
g6ot37KP/kT6oRek3rk0vMP5Gv/YSIfMPb4B+ByHPyJ5J0pjZjV0oWVEuTV2
1lfQLRJbg48917GzG5XPupMY2i7tODKRaCagqL/lOgR0Z9dCco1d6Q4DPRhx
/ewZV51ou00ISJkc7Qior3phz1qATgluqvn0TQaWF15mgCbTiQGW9PyKPWTp
k4kK+Mbe/ocFLASufv7CPS2ply+t94zpalbgR0eWGbeRNTP9Gp1E0iJQigbV
z0UeHlVtZq1cDaPEdl1coXihXdcpBxR2pDAx4/no3phisq3evSxZDIZRwDv+
J2uv070KgW6E+eWZlRtYvmuG0/48f7Ax7AEMQUZFqWwwCN7Zllkgx56erGuX
O9Odwr5pLKequ5Jb7+G4sNY8GSPGHD8DCemK1l5gXggLozsD+EFMhFKx8D62
mVZ3QR3SzynNRK1rHW8e1rBiWhBHINvvZ1I2EBNsHProp2cNcewoXMzPHIx+
4/RZvzOTbsdZl7eCXIz/IARcN4IsryRi6/SdbS0hWAhhr1hmzKZjCdIh4okC
V45HhmddJo45AjG0dfMc2kiEOx6lop2ZkV0Ds+gSsgv72g30VX5hqbMMfAK+
F1kbE4ZsUDT9GSr7zafAFEc4Ib3AIxjnxuBIgGaMKRSwYfzLkVVOmMxgm4kF
ygkg+zwI31n6LfgY8bkGEWl7PzBefUyZNS3yZALIiG0h1haH8KfDmKyZaAnb
h9jD65ZZiIxVJxjURbyJ5tGEf1vd2HAP4ZUlijlBAEfq0EiJdWyN3Om22oP6
5B0N6/Kc0t3UlHjKM1y+sevRxu1nhqray+Kqca/oJ5hsbchYpSw0qV5ZH48P
M1iZntaBv0GAqmjV+NiDRV3lx/BeyobEIWYaBibT+A8/juUTtjsieQ1GTA/l
HAZdE4n56LzA1q+GAUkJgCnokZjQfZVccuoq5LVANWKLNf3dy+xaZduCrNu4
M8WfKROu/C2RrhC86uV2L0jSzAyssyYRSIO8LzwO0LuhAYITTlSlqALPdfee
7q6eCAhF+4B4w0s26fgAE78jkVTphU+HRJbezSxRxA7kkJrD5HCfNP+WKcMe
Ovi85fAifihb78GkfRihqM1JWLksl//VZ9ZdRBtL4gtiJCPFsEJPvpLQQggr
XY8aObDtdE09elWN1MYs2upsbkMewoaMwWL1pNPK4FauHthSfMVUynWy1tfo
WuqIGkm5gMq9NJgKMk/qtHhO+7x/Saq//fEeHz/dRovQhky6QaQswbQ/lRWO
kbN2ek35Ikyp4yOhZ5cizgiZSYTQdRBn3xBRWy4Df/A2ASbkXsd9+LNIYB2Q
2QRDtQiA0Izb9zFuDmPBoCNOb7Dfp5DgR6/M7HWKgnZMMVG8AUMTKiqj5I6q
MbxFzDiiSeIFzD5Py7KKa/6CPuuiAF/l667c1/Lkd3oLrwf28kzeQkgXqwgU
8zydZ8605dFtD5/T7NDMUDySxG997xBmLnXgMJXhDATQDQgf3kEO/EuXMqBO
DnUy1SxpC11hi4pjJzcpupTGh5P1+lLnLZIMuDAA9ubkxLGrceEAWHhf6ngJ
LMXNJ3wOkQaUvn1rXrdW2Efru0tEoMoHqxlop2hA7CQ52CnQxHqiL3bGJzUu
yNscbVZhpI9kZO2qvN9zFr5WjJrZFz1lH6IPIw02LvMhnJ5X1SF4IdDMpoTS
DZPEugHJnRn6pPOjLzx/BOypGMGVNJybo7/1ahaVuWaC7gPh+mcYumX7WAmA
SbJl5iMvnvVZxMAX+IptjS47pPa1+6fvNEY0EAmLbxk72Gcxvo7p7EC+wCXp
/hiZ0Cdi/1SbbckbqS8pOzGstVQHg+syG+nFlJYr3pPOyfnux1PqHGwp8A/a
qeDgCzyYMOrC6+WYO9gTffqe6yORvaPgk99sx50cFEoYGiy4o9/cPlm2DPEv
J88USJ8OQSi5WzdCd0Bd32jyPem0VVfu7ATmEu+zcqmf8Q1AdckaxQ8W2aSO
feII4fTIKZlq3H+SmhPBtMu72xK3YdYhWbdmubfwVxuN63ihb8yNPTdSr3zr
z7fP/nNGxKYCmYZXPL6g5Emf0EGra49H/sMLxgJ3KeB0VBea9Z0ce7svAGHE
DRubDXjjlKnDwDW5FbZ6o67jr4RLc+QXRkwsACHWzhoxOijyz8MyV2TT6pm0
c70hjMtdwUt1I/vGzPSidJEJSci0dIZG01u/rjN6+6119WvreQmNR3T9Z0Tt
UfvJ40itLmT/1ozbAXCYn1MvRYncwk4vH61J7cCnpRPe/q9um1keuc8CSMQ5
fZm261J2qNv2s3qaODSfINHUPCf1Jj8iRm0hDJUW1SPyWmdDUbh7QO6ThZoE
mu2iWriLYBvD2+SnEs2QI4OVkxVjGKblE4SXHv2kMn+kdt94hJIlykbyrVSc
S9R094OyRTK8ISTkntwAzRB6edmzo7PpSR/jwSZdN5aFuhfphtzJFh+0r6st
V6vAyAq2oLUlKC74kuKpte5cO/8AJxVGDO6fZSsHRCPIk0mClLzlOuFh2Jnk
oIsg9C8f4PcyV59DhT7Ij4tmLWIPgKqK0Wn816SCI6+3I9iHoTnJg4PULafY
6wDDa3PmXkMsNgzCgnCuBmtkq7iyr+tUaJlXZ5fVJKkGsNyD1U4zFbXNa3gj
BPJ4Ft7bqZO+fzMF4bj7jAJrQOms7lKalIf/K8xPHwX2cYJc6Akxytrrygw1
wC5wHbprHz3XfxVXqeLi1tXaMrlSl6DiZpSrEnplLp5tdFYftveqn5T84h9I
DtjStlPt/64dPcHoxPwAl+RpPYRIy01fxaOzp41DmDUG5zhMAQLIIC27I5xD
an2PLsSnFNtdM5myrb/o1MYSTSXEE43TLRCj6wNWto/1Lf5eaCmNbKahizLv
L5rZByafamgtchdtzGCU8Ha6Ji7iqfguLZ1xymbE3tK7cYvcvY9LQb4B7x+5
oWeYxRZsyI1U0lzXDUIlDNBQBtb26Plf0QWDwaAMcma92LTTp0i5eKRiWBhq
ZU8IosHAJk1P0ZjRvW9k0/JhBaAgY9YAkUNnU+vqo9OU4BeKPiBeqqsT/HiU
6z5a1YRI23/r968VZ7aGOCJCBIF2Qqnv+wF9hxUCxHMeuwh1OVUiL/iVEvcE
0WNSBABKDE7ke4oKi95bKj4595u+0gm7m3j3xYuqQuEPrg7XTIpHakZ883xg
BMTcdRYxdUeX05uFPZxDoUv0Eld8q3tb6ykJhIV855KHQqIwJd2YBxZMfgBP
CPu0zOdfSXIlc8g60NbJSyKYM6Npv+yXHCmGiAEZMRRIm1dR3y8Tge7FwhUI
fgV3iVYa4CXPaW5/f6etcuJ1g4cj9czxM+ozJJknxos6/HX4LdrpIG1SQ+FQ
+v0nhtbSVMuvPfeapqYqsKFaA7W9gGpNKVNcxjiOcn9bpwCskBPjM1qrVIDg
tgR2NcJkO/a117CinX01fVbvX8v09hFw4RcpLZS4ZL26Z1JwKgzhPK1Tmvjr
iedx2aQ1sRrKqL8ZD96WStamMNQ0+EFvaGPQO4uj3Mh+EVVbXzPVUKILwzo3
xYkIhhGXV7VucHTI3u6TOX1nU3dfC4BCc9cE0VxAf8kSh8m2YFdFg1E7td9C
AzEY99UrowbySTGYBkbBH1NRFnouso4N79wuVJhJ1TsHCU2Tswfe4pG2y7dt
lfjoNOxcGyt7kqBjDl+eGTJ7z2UCDzqeF1PCxHEI5nW2FMGUXwA2h/wiCp3v
swmZJA24Mz7N08Zutg2HIV5NloC99H1HS/c5vbqqqkqXX2cH9iMo+Bo+YmnT
VGqW7Qp+IKivkg1SIlzfUoke2ENNyAWeMQXLZC37K3Or9KM89Vhyg3xQUG24
PTOMbXg2l5GDdmRHjwuzfx2ZbDkTn6hd4JhkdZ4CGBRIxkHKhHlqnLzVfbcj
UCHr8ELznfl1GpWlZwguCoW7bkkw4VFG/oWSVh5PgXQVQHP63rnXfqwfq/MX
4nJJopbz3CGJbM8dDtaP+yxdS8yWxCfIVRvwjeY8yNeKRxxHEeC4nNb735QY
9wMKwfYpxjj0Ty+AKxelFJt3jr2reNmMciyWRtdu6fhd1kgch+Lz99dq+utU
awcUUjAldu+qqcbEXdjoLzOQM287ANgZZ/sYyHK4E576ROA/+gkxQPdikiMe
NhDX3d8Z/TFrs3PbpBXtdA5BLCpfA6vyAit3G33Edulq3EMoDPGGLdYvtrUa
VZLBaaeGi80b7Em3r418yCglNJcOA+0yIRZiN5i0KGjsntxwGf3o+sSB1J89
TXv8dabl8YOdx9Qifa+KKuzLtPQM+P8PxFu+EkInrhmZygExwuZ2M++r0YN2
ai1KKW3PvDXlHLX01iyUSdSU2mxhFV2a088VO8kLa8xJMk0ER6DUaYkDJw4w
Lss/NM9cUPEx+HaZythrZ/1fNpsKoCapnSpKndrR36srCg4ZiCwMdP3dB5P4
Q5TWMyy08rMCqAQGizJs33muJWn75PWhHuwJ3tNsxdSRVNveAU6LvhKr1ZOd
bU48cUWVvFXRwjtYj5e3HEGsM6gz2e7lVDnvEUsgBOKMYaYU4gGD3/BkjPJ5
mxHhMpOhcGIxPZOuzE4IwwaI6upA0trcsGBD8BjAyHCncVjjS4OtaIsKorUb
2Juhw/lbHy7DuINfYYYy+LbfY4LlvNngIPPuo0qtYQYRZHO0/yME3ay3tCn+
4V3uJAsVo9iylKXbN1g9SBgcJ51ciTs/v6hn2XwL0u6AFCW3bcqMnhQ5G4fF
QJZI1HuPS6H+C1bFlBxXAvG0iIRqxbaEdMpLk/DqQXhsDBVyxKzaR3q8IaEr
1jebtNd53CsoHVPzKVugujiftscmBZYro/qaXs/08OT0lgpxL3r9J+h8WOZJ
EMdCg0kW095mezS1WrVSDFAOL4iJSGOEyL3APcsXlmQJEACfnUCYUD69bcIA
n3UoAlU8GTrcHimnOP/E14cnWoWVZvLdIg8VdZZ5X2dpLWYhuEGoALLT+TkN
Zp2xP2NZSfa2ahxgxCBy2MxD7cUSlY2gafHFpoaWb+MpiT3GxYTT/rpfOLWl
FufpRS9vGO3fGLIFFPjaG+QcVd9CE5Jk8eTTTdbvC4S8eRklLtboEle6v9tm
gzKNp0Lmdlb/m/AaVeWbUCF6o+cfno1Q2gd0Rx+zPzxgjee//h1PjYeucfbm
iLfOjF4ORNQbtP1wiOBhLl/wC7cLia68Xll4Y5jtcxNu7uyOt5sGt9f68vH2
7a4c0MWqjjcAFCMEPWe+oZlAYzGYfORb+ZPhnFKyAnj31mzcUJuljFiHxBNW
c/S/037NqmwRmhLCKPXcRI4PcBl7DsZME7wFv2And5k99nTjYMJDIMfmlEd7
ALccUim5nMcddAyV6Z+K2kChYIBG22HivrVB6AzNGfq6QxCaqidrazbMWWE/
522PRZY8TZRasHhiJz5vGuO/zEAp9nDa5m2BmNVGbQyFesD3IG5/7m6f8x33
K3ZUZD6x9lzH6xrYBJ0fx/I8OZHs78EIHNMJCyxM4j3Dc+3yaqqPqvVIlit3
NQXOCzWb6orrybplfy/k+tgy8mlaCs8VQCSADVfPCJKyXlogbZiLNB85dE49
KfDGoIDmW5W3fYo2wK/RosMvacB/87dTerJhC33j0gK4whJwf24zgr8Ms7kQ
3LZINzODGpM/sBW0eUqVe8G0dRxWFvbXJWRxevbjqo3eeWNmuA5DvYiZayZY
8Zrx8K34zxGlIFVQRDdYVDztNahFW+hlCv91qMPufgrlicfvXbcQAgh/4Ajd
FcF2h34GBMc3IzM4LIsITvxwYUcFGYf7bD4nZoiQCZ6nOrl7Z09Hz94xY1yQ
o8zswmGcteo4JQcXQ1663o2tmFtQ86o7Rz0NG6fmksfhakUG99GNirWkyaeL
8wzEFGnzxnArcVkD4/ffZ6VHxl8T4208L7J/ah6aVOcIobhelTkcmPOFrzwR
HJEUvZ7GAFvyjPfqG2pDx6540RJ2UOBxxmW7vZE8lrtHLzgBLzVSktmJWBaV
xqcM4Dn8EOwrMf1mddMPeWWTlhlIf9U8xYvDu3sZj5nG4ErMcG6LjZK8hjcF
iI+4MkQozb+IVgM8f8tPoFVhKYlARAob8qAT56/bIHnc64DZgJthGoz/QQBm
xzuAe8gBEi5uW3vlk9qctE9QrcGUbGet/Ymb1+kWm0GLDTLCA/+7lJKERrHT
yeMYSQNckpGvzciSC0t8BALS/Pp/UnQJxFYpcGHPQCGFMGKutbsLrG01ZT6F
1fd4KD2Qv/AlF9DXMAqGdw8+u4fYCUW4sA1UQNySnsNjApN7MV9nbq4VoHRO
FeUTG2AiAnLT21rEsxvmoC3Q1SlO+ipAa0vUitsHvc8d3QxEvdQPL9QfOGnz
znB0esXgtapU2MI9rDdAmHExODsKva3EvPMhSCaycfqulNVxH75OQ6PN1g4U
1+FDoySUKF1WEgW3HlWwQOxKVFyfrx13Do61bGDzxjuvqqRy7Ocl1KgPpk8Z
IxrwwwxMwZe5BS/C4MOCzzLJ/DYRuLRzciOfW2sLOGjKzfnc9piJU+DD4UxU
sAWRa8W70qfbkdSouKU6Ay0v0s8tj1nmKTSNDliMqile182yqKZ5Yz70WoEW
vyiNW33d6euNdIp5m9n015L51sxraSuUlk1yIG3DVcWPk6uqgASZkeR4aiVE
Sv2c57C9GN+BEE1K8RQ8ytUTWP69S2AhDbL6b8r6gowW3jUKuhszB3QcAPlf
HtdR7MioOTuaYb70cdFuvfV2mA6/fkneDqPpvYQLgVOOOPKOpq19bKRJf2e0
OCqmxseOv321IOSMcT+VW4C8Ntf1Avsq+cItUjWHZyLpXqMgAejWzUTOngI4
ehUbxgU6TDFVV1OSMjrGEamL+G4Y2nxY/PWLmY7aYc/dguUjWjo+sHpx0rhL
O7Jm5cUYWDsMGnBORjMEt8V/lkKuybqPVHvtiRHdN/wqAaSPChqs035mcyVO
4fenmX5tCpSTfxKXhHc/avlGYlNFYqcAVCPPmGmCcODCAZNM8RJkwMoh0Ll+
vZJO5EjtI5CvuUEk3ctt2TNuGxSXk80tPDkozCIW/aNQvushFBXex93HFVmz
TaD39xqp43eKDxJHtdNOk6s5T2nhFgf4Ko5qne8657HOWgXUhfFWgSjgLO4y
0lrPhJYyDvqEaiR3i4rnqpx736tFkzNn0oGx32C0kt4qFYZqq/H2zR+zfYHe
oxKJjMb1WiFPxylr4guTE6nWLKgNPLaIQLFNGdnFcrsBIr4TLHYd36gM0JoC
mv8Zpdejq5/CPg6LSiNNfecEltbeMxr70YDSYoDjA3cTDeXAt909jgH61+7d
r7YKutXGoy1iBl/hLkB06/Hqjd4D46kfWLvj1uwCfhTZHgL+aCm77DOrewUV
+XTngBG6eIw7HgUVTsZuKCNjLr5bEWWkNOUGLVprlb3U7JZ/O5Pe/4SZhA8T
qypJxKJV+7lTYaRrHjMYvrVgvCdFMufJvMldcE6Vnr6CsYKq1mFo3B4XrZ1k
3NQehUDMemsRYK4P7lD483i7REO2i/gYI+TSx7zqQiMnyW1iK98z9XaADsDm
OUXwFzVkQgfaUbWX3slHCiNzUiv9sOL4cTnudkmoLycHKlKOtCQt0HBHgGgk
J3LPvaZIyu5bXJfvhYq4G7FJXomJEudaeljLNAHkFTHEfuRA/TDDIIkseIBs
41HYNbKHzbdfNEO3t1UGZY4eWcnsUl0efZ+FQ5/uD5eGmmbt/XV1CRqG3nHr
FmUTo4lnKjfq1l7rHD3mOXBnYgEOy0ihf6iUtRjlnLA7yr3+Y21OiayVLXRQ
E0yAkbIhUQX/sU1BfM7SS/r0q2ozEkk3eIxgcef1ZkhvpJnz91OyQtgFNIFB
d8vg8N67xbMYeTnV97TvNgzyL8lJrw/Ur5PlI4TA3jduCRVAaUq1SoSsKMY7
1Qu9EIqq27c/diGNUO/laoDtcfe8Vt6KuFcjupyIwc6Y+l0RVrOR/NoB9sK2
3cfJDfVBRf78ujgNn75RjJVnF1oItgAOWZZRNakaRaoNbTLdOrfIgWGOvKOF
V7OLJ0Ot3Y/iQ2onL1Dm1BEAv8Sx85E11NDYo0AjmlSL3UabyTol92a8FYYJ
uueRgMkUdA6AtJ2SYqgN0zbGf+nUZ99ZkN2Ub8qA/7RETElfrb14kDq1H2y7
XHr5Zs/UbnueKwkOKCXC7wuxB40iJYKUy5dUDJe4SNOf3fsY4ofXDOz3IF0N
MG1linGvxcm8oAR3AM3Rxo1cn+9utqZa9Dg5ig8ALAp+hNp60LLBogiw5P2p
8FOL07yLBWn1fNBWr9EnJWImJcDFESJmBd5BXFVuRAZ3j6+ALHeNdRENTHuC
nTwYDkGX7Le2G6UTpIu9I4H6mwZRQ6qKTdnH3gedNJmLbla5zElOui7QDwcx
ZLq5GclgKM8r8zPTRqsVuVMVAhTPbs+sd0BUFqfFRglVgXmNozT9nmTRvA1a
e5bMwQtEyhFHpjUG+H4XH+WMB4phmtz59r6mtqLUSF2RhZ3ZssRiahs3IPed
zNq+3+ReIXiyZ3rMov6jZO27k5PpfOGIlHLOrzqAHY/GDGMHOEINkcJ/pZt1
l3/iQECA9e1EqhLPwOvoT2I22nIVrMn7ZtRuW+b/hJx1xUBoPyZd5duKbQcT
Mjy5XvIu8f3FwgEt9C+Awed19aWYPTkd2AGpbFNB54V9Sd7p45wAPC2Lictz
W0Rmy7tWhkGufkQFBUgxoAz2kNDtEFmf4eTEKEcCL13w3VJ6iRLTvv9k7a77
9qYN0U4+13fDq17V1SV7QcVt4GbSgcudsRqiRhpdEWzp3sOioMPWk/OB/AjQ
/qBRxgnVpEJcuZusPWGl/yEqxw7u60Ha0AgQYVovOgd3GcTP0vGtsAKnBJbd
ZB+G+AyrgdeEBY+T152rQlMsnNwdB8w0YimxsjgjVAZlmKNJVW5IHQ1ZAeIh
/nfJfbBHEn5zXJPmqkD13hUupVZky+9vmmGaMAivnx0aUmm56wbMW2+WpCYL
Q/b+TvLvBWxyYkoMpJ8A+WW+yI/mLWI6d9nXlx8SR2UGuL9kxDyxz+ZomHpE
IEecXSHBllcnkkk2EUG0Ot8gma2wDHFIu+hJabkju7UZ7Glytjw76QrJg+lf
eIQCpemX0pNp6eAwGfDpDHhMrxD/b5YC46Vldg555By+Y9NkVe8VNG196cZO
VNlOTuRxOyIoJmKWqqls6rDqugBgIQDY1MWnMRPUmKf34ClwCsn4fLsq7Nlg
v9R2NNq5uourSNiIZsJW0N6xDZ4PZ8WoDbkEJPYJGMFpMl1cyzWUjVz9FbPS
FAlIxkgwn/DPj8wPc9B0twn6sGCllkrHobRyZUQdwiX+ZCXTnOb3wKdtpqVl
cUWRDblAQ3ry8/Ws5SVDgMSlbgwK63mP3RxUuC52+rowT12xm4Hgbosj+KPS
+ubpCiMOylGhHw/aUht6Zjb/ewUatpWmGpfHMUsC61QUKh15w8Y3sqL63XgL
KKDIT/DehqxhbI1hi28ZhFS3WIC5hI+7racLSLYHkeZziburkKf7WinjafwT
wx/dAbsqRGmgSHCcUlAS5Z4KeXJwZCGZ9tbag5ZZkkE5zBpW9R0uD4yoyrsK
WZeBl4OPKDzeGeMfAjVfQJBcif2+zOGctzTo5FYS2gl8WCr8KKfD15DBO80U
X7If0d/Oo76wkyUHnqNiNKJSmJPP5+175lfJ12O0kGHt9kFuuNNAh7ST6XG+
KXAg4OsKHgLlS9ijq3lCOc2a4mB/Iq3TkSyJx4FVaeF8RcM2NhH7UkBH9bcm
gTJaqzRmOdHdFZ88D2NXjt0i16JJxxBl9EmfhCSMFAb7DE4FGMTm3w832yZm
q0Fv1A63XLNN8LfmQpMVscxyKfVIaAEm9nK0+T+s94HaST0+Zr3aq/nmSOrM
Ktv1j5xQy9x5GqB0U110+YVJm7M5/DEnp0nWDXje0hcC6vTqwPkPMMzY+BvN
DEa2EQHzDAy9/KMLtQFqUITJpj7gDb7cVberwbiTiK77HqHYrW+yhEOUC54g
PtlbCT1BcjyBSf1lvviQJ031c+6dh3wbNAJwlabtxLNaw99lhMNJ1PJ6o0Cn
aXN90QHfk5vam3d3acdlZ8TM5gT1VZLQdJMZ4ARfD7gn5+SBox6/POTPy30M
n11PTiOMiWfgSqPQ/u5HRj1xrHPGoEiaiaeUHhsXM38KVEJouOOGO298xPVa
JUEZvhTcGGRmen+tMISAdFH4WGVe8zo9jHbyWSyi2/DEEeIhL5ji9sh4be7v
Er7Mt6JheSYD7N8DSzXepmPDfs6xm79tsTZvdIBaYl+pXJ2pVtgsMeQ0IJf6
7ID8/js5PputHc8gmyRuYDWOrRTpXQS9WPyZBfR4gsnuG/P1iXW398e4hYn9
bGSkP2gX5h5K/lI/JZVf0pKawKjyDI9JAvFcvoz47aQzB7dlxDix40odMvlz
JwEPJ+uMKgAiEZwE2wHrkRZfYqcBQs3p2PyTJ5iNnClECGETUUQul/ovU6+w
aMAMiR1KYyvHlGXj89KPINeUXeSd87nEEjHRHLULp78YS4BHTlktuvOjlNy4
8GWidzy/uuCmxtwiz05m/v6clzA4F1aufyRZqAC8SeeoqBsh4aQC+RyY3cmt
/6j+MmKbDLPfF2FgW72HDggE3LPyvFUvT6OyEEtWb35KMwCERpZpRkEg3sGi
B42yaMrv09/f9HfFqtB/9+5gFhPWK01sl6T3HO5hqOcMtL6HztwZ0DNVhVnj
Dd/Igf5a/FupvMib0FrabDR/1pWfkuq0AgHieCGsDNx/+Bk9iBB7wZ6Vv6db
X0lMr06ubgt2VrVLoO6OMwFKiK8PgZr0qml4VY/FMuc2mesGy/ZrKjRzgd/d
ZXwdXeM7Pa2hdGr9GShXBOtIxrH73dKmzQGpMr18twg1B3MktGAsx/POJUgb
Frot53IA/jQ+yw5fkffsjryPuuwrF2jB1J4vYtvqgIub5+/7qAuzgMcAt+IJ
kmd2sqz37yR3f/S74c2QkrsRN0E96zoXtzXWZGOJps/DsIdeq68nAdulSruZ
uJA3+P0ayYZXlhLEmKPmH4FXfRUtXTRsreLow2Vr8PAqUxACfjJMPMrGmFq3
bDm5kPREaTGt7obLYaDhlCLf2HkhVRZ+nlDE4gpDL6mzUhef241IewUfEbI7
2sp5UPXnxv1Vu1ZAiNog+zQB9u3g1EFOYBbiH2IZgwy1Ws86d93NHAeWaW70
65LDWWtDjWvcmnO+ZkOLBYwmvOlk/Ux6S0ey3TeFkPL7PkOZvW7ydjr3t52M
RaGMAy4kB0HQP5Zcez855sVMdCv9VhVzBuTjqCsLPEq/Crf/w4Ugk0p235Sm
PBeJ0+HzL7L5fyDQtWYWBcQAlyCF9054/4GitLhxGgtNQpoxfphMhZZ2e2De
TUSH2GDkOpj/yAhbjoTaVP3PyGboi71fDR+tJCPUwm5o4SMWItI/EtZFhpiy
01zRw4Mtk6YGxPJpaF1z0szSudc1AoEQpI+OtdHzjwBol1muMROeeXGxGVRw
K8G0J7toOkS0xm+DxMGryaywkz27qipz+Tu1091GswM/iZSokCLg3piJ0opp
lGF2BGnKFckaRiS1t+bN9RU4jUnRdq6fB3dlmXoVRjggVo3vsLhqBPrzZYpD
jYTt/g2Wqq4THyoH/gFkjotvbIrDRBdbwH7A95wPt7xSEbjDFNDryFY3sT7v
rtMj4f4+Gbs20l8DaLfQKeMJFk40SvbzcO9VikOznqZ1n0CgkwtcBZmfGX3i
JRWweWC0AcoWsjU2wWXfGeKQk6OyM9Sucfk0jHba4yXjb3tpoxdfM514qs0r
AGKrt1enWc/wcT5lAa6gyUUCwV/8ghwl3FtvJqh3UDW/6wOj498O0wnkBGJS
8i4Up2rwyhU4qo5FUcfB1urLg7b49DqVbrd+u+SxyrCOA5Fv9SdiHCizbp1Y
L8D6J6cwEQoStaMoM63MU+xij7AxqtkKEmtFEbWBfrRXGgtbuCyX5QFb4w68
7TFUSO7VBoJsIrPyS+k+SkaWZF56FVwBJMieA2b0Z8JLsqKHcXCBqISXz2fm
1f/tYIm7LpyHmrhQ+rLX4N92k58iH70nZwrUgH+Yoab4CntrV3gcZeQ2u4eS
wyis3an8xZexPaHz4XlklvRjHP1gvH0lyNMZvNaE4tth2r+H4QpZDRwUS/Cx
myF3jPTinCbcZR8Z+wOTSHwI0k8T4utYIuLqzKQss47kHV3YjFZOTGSZtykE
aAb+PjPLoDzmycyfVo4YHkvzZTLMHFS5A3l4eqwNZz+zAIZR6tMHQ+sWl0LB
exukMy7oytEoskkvHCLm7weSRA2A0bMLnK+CLO7KaO9hIhNeBf1bId3VqtG5
bTB2n18omM5qx/mCX9oz0WKcZq6FH5gwsiI2q2Es1tCTiXw/W3O/JlhvHnkr
p2jbCzjxBXDXlwh26Yn05XI3233xYl+e90ksDh9SxSu8HqTZUWG+BruuI9Yn
AhwSlSzuuC6IxcIJ3nMakGhKpHONt11/xrAcgc1jXdufn4X1xWElBoj4sl4X
PxWP/djKW3M93J/d+o/YhL9kdtnSj7oF/xo9fUEAgF7SRc707UlbQouKH08E
uVR/B2c7CKEgYCCOR7ZtY0rJimj/naJ8wElat0oaE4XKM0aKbhId1ezk3fGG
Z4S+TY3LutTkc7pfTfJmqEhINuhCxE5hwY8/ybvDmx26rYs++U5v9pvcY5FC
xuYmBdMbDOv9/t88Wes2srpr0UcZQwrQMPtToGTHkPw7W6oxG/Yl7A0QtIKW
MuUfJO4zMD52cr7/kFXbrzJUTpaRW5bVqiZUYA/NXys+n7bFPDlKbov6q8t8
/0ncdcbBhS+odeRsDU4D+bqJtktvi5lml7NBRAWG5e6ACWlaShUMCjO2E9ks
f/3Lm2q0rv46wMu4MuzVguDyBLDXp3rvr2FDJ6A8RHRZ/uNrj8bP0x3C7Pv6
G9mbBdYiK5RndwVXzwA2DZCW1R8ybq69lu8BZY1lwFZhs+19O3Y27LSbfadI
dUrVM8VkizgSCC14ZmcRq9DnW/ogGSKwTKqtBYpgrlkFhHlT5jt5SrZt8QYC
Jr59D+WnbeNUohRCp7QMI7BQWlvkMmECg7gVITQj2oY1BHzLJwxaOyCmz+Tz
NcnW/29I+Yk0KCMngPsZ85SAl6Sgmn9GXkfarvE6b8oZTJDgB61cvTayD+q5
LfzbA4c1fLL3g57a12XG/+7o+b0ivhZnRqPCpexP3XjER6TdMJTlxjhdGfNW
P5iSqVKvClRCcWM/V2Oez4cMcezuq8K9PWb+oPC7qXMz1Wk1CEjdiFTCahIl
D3OaRm9Gq9v6Cvyrt2zqiJlHeKVzAzZTjLBlW7QtgTT8y3jDgka9j4X5oClM
2L90BWOPWsy1ywC57qcRLc96mOsFskI2nKmsVOzoZ39gSF5k7v2xpO13AD03
bk7k+zYK5zbapQfX9kFg9VST/tFyO8sFJIquguPdyHSZThpWexHA0YplOkyk
BqAWhVqkIiChB5BdAUC4u4M6lQBmk4yryOo6L371CI1kpHFVbw5LbdBRWM4x
sLw+ot6oVQPbyqIfW07j3rMekyb+VeYxb7Uc+njKaphc2IWLUgJKVP2v4N0w
fGu7l2WoomTz6kvebIHYC0PQtFdriu/eCXWcwiLZ9Q+5dLZbHkvduR3kHfM9
DYSO7EkWjctDmEMC3Hw0NzszTjKNDuaj/zdN8YXAdCsvyB8tgD2mACU9zPY+
RfAH6blTFfn6EUyzY0tkqKbJJByrxv3plc1p4w7qRXMU1YK7/2Ojc2oYIIr8
OmyD8GblwlT1deqXHtPhSCoW7P7lDYzHOUF9RiHzgBBdFZG1MtbxPBTVNOPx
iXujuE4zHzyFNS0AadCIazHQ5OigAW2W/G0YF3CKppA4j+zozt1P/iRQwz1C
hXm7sbROCHKtYSsxlEDFWCxiQPBLOV454/0mzuqF2QQtG16zWpEl04LO0mnw
Kp6ZAopuWXcG8pKCvhGykZ4VL9ANgWXz563uLjnXpbYhFEuX02FTMi6IAcQ+
rqnMwO6518myS+J6yKclCQmUoTNhhEns/xAY8HN0O/Kg+mGyA0PCWmnFCCqr
ujm0fXRCciWqjorbwrssVBzG3B3Hscv9ZCFfwdkenGYqnhIfAzCALCW7NQN1
n6XxH0w2es5PBie4nqL3iEWwTKnLwxEVEoAWFtyHL5qTItXQIdOfx3fgK7/T
cGDNABgYLSrjzmAyIusR0VQBu09Zawofhqhuji1KfaV0KGuXEDukB8XMPplh
77pGXwv/nD/qf9VFSKYIXE+cVluds3oiGD95Zzpo1wDQzU1S3Q4HLDU7Id5X
1p4+pguMEM6+i2GEIG67Ub0Lw+VKEgTEmhpQM+sJKXmMYNZXJdh+EoUFvCWz
ITMlH3OrgLcY3YO8VupdrX/o9sJQ/aYDIUcd5E4aKIZpqNESnfSuC+/W7p3I
9I9n/eWIMvbJtlIyBv8qMfRoi8/iwxDqKWBWVr7KxMBWVz3oi/Wgf3bP4mp/
/0Lp4B9QpPzKxfT/TZBZCUIuZcsugriWqf8uC4baNLdOdd5Gy0Ee9uiq6BPA
+iLvL2l3BC+fNAs3xfhvSc9gN2f1FRPab5tAWjr4vCRnnj36p867ISzqgyg/
zuIqZ2W92R/B2EV12hm7oaufgDL5q1Op+t+CBcwUjMWwH4eJlPpq0wolRQmw
XavdCFazlp5gVO+wwzXE70F/3g2ELYqUeNpIqmm3Yndw56DEB5DhpwcCyAuZ
W749NU+eJxYgTv3+oPNkgPsCyVhYoabRUUFqDql0gJp+Rxw+eHsSZsckxvt+
bjcinG2qWB0ZuPH+G9X23g3qxEAFsnjPLaFwQiYcb5i0zYpxetFTLBaN741S
RWbhreBrLEeTEmKJn8YhxWqYm6KpO7LrrupNjd/mQCHA+7gZIG9fiKTWiQvF
RwUKHCnr9y4LghtMqA0lpuBF0djrSuSDpBJOrKYBotlUKDj0XXi6txX5HUD8
ecp/qe7hLINlbPCaImd/E6gdupcy31nVqL3cdCvPwzrwzegvY3LdZCHqv6b4
pHD3UFApVjX1sjo+8fYKbriTSv/ljtNIkKjHQ7qb0OLDxGX1IPVclsqycCWw
1Gm/956oeD9t1UHH8nAY9Y9Oq0sBgve25cRsT8EuIh99cSISdrohS/WkeVSl
8bSAfSPenmfa+qyvfdTK2aWEv8MOzKV20IC7Zoiz6+8mx7YwgyA8vEZ6wG+b
3drAlYMZmv0+md6RZN2gv+plVTG2LiouE+0skJHmOx8a0aE6Gwobo+1z09U9
BTGWyCHWijx4/2TI2sL5xAkkpxgqYpG6ejfgiFdvtNOTWpVDg5KR45jvW6XK
abD63dnvPyZ9rnbhOMLixdb70yYY1mmtDD7I5FGolMz85i0L92R6a30woTxx
bl9iyoQnjvHpKh+d5xAN7PGB93thFaEwNTuLi/SFZXancktSQh77sOXCtqms
JsmQlrVtJAFYk/M1778f+Y6HGzVB6Q11hNPJZE4tt/akYCKndLdhkcUSN2YC
Mn5qcHY8z4Y7Pkbud/GOiqMonOn3wCVCTcZHgru+tvo0hF5RQmQFLB+g/N3p
oLwbA/ur2XhwAR+9HSOzLGYzUbKAmtdxbOMGnPbPHeBdNSJfLzTdGrVKE50I
rDkLh6XFrGytIlHPa/5RNxIM5/oS5Lsqzl6mC1dfnljjDqcvZBM+ufz1QKml
x+7QMKOXMHHETby9xVN2NkJpDRXcNupJVO6b+BtQXPxIi/WoyfE/iwCbZgHE
xZkXL5ZMtAdH+zNp7iQLMF8wsUvXtRHzyhDQw/7hycNw4Cu48Z6vCuVwOG1e
ZuhWSjo/M9ehnTXR7UMRdbkM5l1lZuvTOx2jxb/WBLx4QuScIz21Gisj0HmR
M/aBqD22NZovaI7fDXwJrVO8lEUIp7KW7C/A8KVmTEA8gPwV3gUrL1k72GeP
eC7EcqlL6QZadpT+BcmFEhhIJfBujQ2T3+/MZQoUIUMetqLWggwbnWA+Jqsu
g/U54vgdNXGVbuT/A3EfzrUhSQAd5PIAQ/pp9DdYf/iqlAI/w0fSJQIV3HZQ
pQR1cAzQtHYCEK3t6bvQQ+7X6PttVqE7kpe8LYfFkxangrz4XKNf/yi4Do0h
WlbUpItVB69jtEfRnVMa2K71TXtdZvtlEhsNHWfGBmLkViZ7ae+fLnaUjppr
LrmyGVUhoEJ0GNxCdgCwCu/+0gNwtrBMD5SVdEMt/o9RpKKHWaK0zov/YSxk
R/u9EqS0xds2wowoMD/TlgwrBmq5BWOHqynAAdrKBo5xA6jGDNQUdFOHMP5b
O0T5W1Oy5Q4y0jV9IrXin5M9qMJk/1UyE1o/RuqtI3tpSghg2T6h3bgJtLrU
6oHtl9IINW+wE1PkLrNucUZkQkLc+C5QVKgbLDCd3kgyHjNsCNsOHHxfwYaw
fMBJYEIWKx2tPNzVHPIbFKlWu4NkQjDiawStg7aO5VYqgGj6W4aIfwK2bRGx
otnf+wHMIorBwjdhg9bc12dORnurNJgQAuupVS3y3oGUfFgdyl1IkIVBCZll
MUq850RmU9y2NrGOqlkQAaV6m52fBcb6gVE0XPt4zGCKJsQWHY/YdTL5qZ3a
JC7VDERTqr63QNukQ0lFBKImELx10ncI4tgKg4y3cY6u0o/eGctuqPpFJVlE
1ctAeQOqiD5/52kXC+oSCdKrXto/lVHluKuifZWEggFSb4fPTHBrcs9245z7
c/j7E9U1HRVNa5XHWvbxi3HoJmtNeehdMvt89Najf+t9GiwcMVoD/oVl3IY0
tWPwW5s3LoI+qFt6ZuU4ZmVIbZ88kfz8FJ6nABi3bi18nHSZMYD8K7sb2qCm
E4bF7x0oU536T/S/8vjVHM3kSDUxF+vUUW1AGIWUlaHyBHnXLDs8XFwxNL2u
nU0zqbTQ21D6TWXIF3kCU3kLn8baXD+o0msPQgvJs+5Rlx1qo7WTT8UU/bx7
ehvX/vSUBUg2w/lOh2916H/UTquCjSWlEIKW/1TdGNrP+o3Jm1DwS60RkJJH
9QvsClptI4ZiQV2hW1l7A9yl599R1gzfE2+a+x2ZOLRXGzWr39Od9VEi4MER
h3A2OmGSFIda4mUQOS/VaAbtsVSK3KpFt4Eq6FWopwBmDQQj66Ca/2jZyIio
teIdxrD1Ys7eYv7PpdVRpbQhjHy/OErftugbKHG0xcw6OIJjyinRTR75lCUm
aX3hRzkGY+KHnH/IoPXEaygZr72Qt4MCJzM1rZQp3y/oFXO2CDzOTk8C0yJo
UpMzua8mAH15WJMyi7uzbMchaZJSY/jqIy6joMGPDL1yJ4n8aGDXigESa6i/
ieKBTvDtpiA8ogoZYcfOdbzSDfsgc1gIvdnXJuCthsNP42E8lqiZCLKY+I0F
xLq/f9fbby1RhZJbfw+omFVs6hM6Jktr7iCGZ00aHeYV8lLwTlhIEU64pYmU
0MA+X/tXdFYuAwoRZlMkLY6kWzdft4Js6UhYq8atOnSF2uNUGVAKxxDh3v82
It9ncNouGm6qQm5G/KEJioZkNDQdy0LUPEcRiBNnc1Q7zPHaDZErxgzr+cVh
tdzxUjKFStTINpb6st4hFR+P6yfCcIWmXfKwWOi6Qp4eJ/PAD9DfzGY/r9AB
KNTQiDjEXyCiA9NcCHjs1RggjltsT0/eaY9KklRL8UA8JHYrJs9ug1nsHeUo
AAQglz87FjO+DYlmXrP5G9JmWoB5dBhVfNp8DBvGy/qXTruzqEZYLriUd5wo
ADOt2hmCZIutIVJ4yBFuIqqnhFff4XTkKK9ty1SLu94hFKXxkZ25PX/417NC
3Tf76n1/qzzZt0+oldsksPmWDKybPkqynxKO8HiJwo5CmnSd5r5J8x8HpKNr
ClLxBfIbgciTqeyuMPNKGgTmzWcNRtSeS/xXfYvrwrgcqoVPCbPdg6Qkgr8B
3DmZICG7xzi0YoC4s0xx3gexJvX1cLCSdqkpEQYsVrADw3fRFAZe/v2858vL
ufOBf1bkYYWiJACYVHDRn80U4UjhuJ+GuyQ5MCqxvyK/ajBI9aQRjRzcRrkr
Ehgni9AbyEKeRjvJxAatoYbo7qAv/kL66yXigZVcFlSeMODalK7MLwsbVAVN
M7/s2ZXgghFpHNPvrj4B9cjmW3Gws8PdKf7yn+QKZwbMkA/XD0g7MpO8UHsx
fAfIz8YTO9mqIdifXZ4Dd/TVQWbcSiD5JHDGimVGJXYJBWwynfodaIFTlfoa
pww50cQsAIP7rLnSpizTTpFcdr1Gr9C1MWNPUN5T0c7EDPi8LXAZcXVzgH4A
pxmMUoOLO8H25tFr5NrVqfXO9WVx0xd3z2jBXXgMmN+goABPLKtgX6zY6Azj
xeEb6TN9dLLXZ8HbM6J0cEIQyC9tWoIVgkwOm0OcN3wEEYaVolcY7TR0PoI3
FT/AJkELJDwMjT1lClSG3sJLxFOmT3NDtcBzwRtXMyiFt8M3j0UJo0U+ZqCw
XgIr6B0C19Xh57GI0TrO/Lmnyt3NAKp7KPXwdxst1kInget73dn8umw7sCtw
kf15yNCAG21Zw8OdoAvBMFl/qdhDPM07HriGbA8j0WRmZou9DrxMbVmzZI07
RYuPQIgyObirGYfLEJLMUMdYmxZCkXUQoMVHLi3zcvL2b5ak3/B45TGbq8WQ
Y4KNhIKgawTqqj9V2XF5jgj3T7GYoM2PPrufkYxZK0qzrf/+HdeTCA6RIQSg
zL/6f8XW2n72gfF3/tNShcT1hSEVqWAFtWQEepJxjaSrwRIGXMPZpBpJhsWY
fYuBftdAnqOxxkw/HB2exRtbOsbVqi+udu18asRGZAK/nc4ByoVJiXw0Mxtk
ZEK00jfZ4/nxK+upSQ6EFgOTKUA6UFSJnsh+jFGEe6L0MlylDEq9WMgA+Dvi
WZq/4yKfiJ8Ts17MisdFJltpFbb0InQJ2STIgWaaXxhgRgg3cANrWblKrekb
gxyq71km07I86zsYoiV+8tYu1Ut13Zsvgxxc7z0Qjmx9ypTF29XFpqrKK41x
nYlkWkWLps8r8689WiQ2trqCCU8E0l9h27qAGvEp428Ob5dOt+af53N+IG+2
CpLFgreR0rFHQxVCUdaKofmuGj73QNM7qbzR5i0CWVRVvaU4iW1wWWP3bRuk
XmwPudHbzhGWo8Xdmo0e49Q0kwgxyjYD/shKKNJJIzypXjrR6BaP5FPUZQMT
HBYIGQce3i+19ksw0T6v6I8Gb398iBlspkCs1bHWN5M7j5B1OXsh/kIUNO7/
nzT2IfTKfRoUiGf74YWEJer4kEHCMw/vKhfOg6/eOJ2gZWchpe2WJcWnTFLI
Nfth1KRiYJmiFy7tATNpGkLda4PtEn936VQK3bN7P3f3J+ozQ8WL7ALz8TRJ
0LK67Qpg828kiP+ahj/VRPDxJd022hRKhjrGhAqbhPn6PP92pbm1QwJE/ZQt
ymX7FytmudYgz+wxY6OessqWGqtYk3gSmk+la4EvvxLoD0lZ4lCiqLfSDJPs
m4BdmCuj2miIYeS2PVh8fLrVpDmW072S0tH9UOwdtS/907Vi+xSV6Xpwy/xf
FB4AFvq9BndndXBfznOeVFYgDMUVJxokGDUoO+4nXD0Gu7H+7dZZ/oVG9XyB
ELROizZaeWH4mDot33GrdPwwTdevxvACHJ50SOFPtWqsmKNOcyaQG2Xie0Yk
QWj0n/sGfkFjvmz7Njh1kof2P27VrQS06+XFSUsCWqWD7oMztDpd/pycVRkA
kl4aYfzmUPfe/2JDKg5JdAMTaOLNVylqCLVF/cbLHuzGfCNOdQATEaK/CmCD
vlMy6AnluNOKD0qhmMYP67R0R2RLWit2ZsielkrX+4Pm2Aba6aLGD7vwuzaN
iCMleQC19dpziXfa8WxzuoQ9ay1DLYIrWz5mTrPufGnP1eTfhkm1H0dlB9mi
5HiWtbjLcqlG9QvwsoGWHEXZ+W7xBx5ScGYJDQNb/ul9+Xh8/21F18ealAiG
vngJtrcuMLqzB9n1cdFYYmBHDnWoXhIkAnmxmbtF9v5pUp9BPevogw272MNO
PIo0pD4a8tkEKI+WAxbLTRz4ne5Xukf+wjPi5a3YVPIfFPmpWZYLbE5xASwe
91BlJVcUfjVUsS2HWp22ecu7L9bR1lXp8psD1yaov7c/yOuX3e2YUd99slsA
X6yHP6d/y5y82jfnL07wo4rJitm3OaKtQ+TFB+vHBEd3GmjFG7GC3O4X4s/X
uFd3FPcHkdYUyrj9QUqkaQ4JWSBcrtuiJvTP82JrLN6pdBBVxyp2eGhpM9V6
z4hN8n+gWuinlLm9nxk6w/fLqCp/JdgDCi4oMnfgHtsalVASO8lZv3E52B6l
VKJYU6ylyqLX8gCjjXflEdYqh3pL0zU0Yus/NVGraXlkmzNpl4XISrg9HrLK
DbxDSq+wvDWQLsDtgHizLi18/VVW6iEFyp1xrJfziqngmOaDwaoEqyjno6Iz
SvBHMZ0u00lFIf+VWoVsQg2uore64hRUAuyaMMeND830NmJK73tCPoMDNGBw
vFY6T57fn0tQSyBIPEPNWzESA7l0AeeivaCqK3KYb/ArvbiO7I8cO7C4dIxj
vIHmVSTuXYLhDTW+WPxR5xYV8z6+vy/WshuFzQtIWqoR2AXVJt7mo6KNuC9c
H3oJyXOednbK3mEt0phv0VmobKtwT02YDA91NcLXBxPWhDX+7b8AjTHqxgDn
a+pMKOMyMgoBb+ZRMHa+YKXbiNYljZf/8P5xvS1uHvuq6fvmpbrKVsRGvwJ8
h7liVDL4M0iDJ9o88ye+Rl+ZCxQcKGb8NyF4zYIeF/XRUN+2DHr4lTHPJpnP
lKxmlXN/rgpnznzsdBAl98jV+qw868qUGJydWzA2/hqqPIWancOKcnt7c1vX
8hocRBU0c2bA1HA/QyvEBQw6Tel+6gX5usnbgSwmWKyGMJqb6E6el4sR1esy
B54/FUlS5nQUxP2g5R23LWSkG+PCuBSP99IkSZPmEJKC925DX7N9CQKaAxLj
KbSL40s6GO3UOQE9N+EpYwtRdDGIM3VjxA8gzm3qauoyJIl+Jzt9J16k39AE
lB6lVv3t8BYsa3Cj0bu7Ja699BzSj/K4UbXXsf3hpamG8L96VPJqsm6HgMIE
Z/1sRc5HEhBo5OROlMigQXDKijSUo+QmeEzY9p4U0NdtPGDOUYE+9TfMpE78
AwAC6erduLKe8QxkOvAolgCAfB/mclYhPL3miQKmRSgmTQon1TSx7n+pVZEv
mayjTvomBmbkI39dVqM+sjgd0r6r6mqqKiiEh0CQta3NwmxKCVt0IPCfo9dE
S9hwGxmgz6KqSXa5hrgn9GzOarswVUOcVsatjGj7VCq0CjbnyRE2DEtAD/fT
44tt29XiTwCXi0jVG/Gyg3UP76tUkelMj6akX73mQo0WurPgMx/dryh8jBZG
oQ++8+SeHUFRjDnUhprlW6zRk/4yLZZ4YvMKPZcsX5UgoWuUwvMn7Ouaz4ga
rQv4gV5XU+pEYEISryKFCJ4kw2uCBoUJ9LMc1csMngR3ZoaImioxczCiTS7d
jne76FABTMljD7zguZp+slWe245zuXjuEFQ4gz12p3Pr+ng5Jjj4LP/2EBgH
bNS372ppM0jk80V8vJGWQYjas5HET8RSj7q0ISpM1GFhSYAlZL2qLhpn6zFn
HU+J/5m5LG8I/a5w+c7+JbOGAnO4It9o5GAHwRUiZkq+EcYasw8l2mJxffRX
D8VCDvA3LoIMY8+IJdYCL1aUEnjg0j0Rp8qFPqYUW+fUrhNsXa2+jT1KL7mh
monnSHqNGe9gVAl9H38nsZo8KOwYhNjdjkFYDaeyKHGHtmP7FaHWTw2Md79B
cnbYLHzy0+ERRECsBT4HMmRIiHrlRdVevB7lc75pZ811nJBK4cBXTLkhO5jP
wzQacNw29tt6FPQ4PQagkKwLGTwbsm8hBEskE0IoJf1+LwrEwCV19fPV3pwR
XpQ9xJfzcXWVmgMrUQ7uCJICROozMI1Bx4mXxW5kw+7Kz2A03ak1yEszyEqf
uNPWobmYtZPoUhPKHhbPk0A24GO51bHCkFgNR98+fKDLEFV5dmKfVA5NmWux
I/Lnyu4uvD2zsal2mZfcWVNys3dMSVUDmDxDz+40CARFy7RQybOehz3kfuWz
Wi+lTj4cXdcwclaKGD9usXdL1SvCrLZo5QP0HEGj3T+7lE1SC3fub5C0/sfB
Aalsbx0SoIw03mrkWFOXT59eUqUjdMADw9JfNW47d33zd+zh8AojrhHjxhHq
X1AGH5u63d5p/PzXvJxVZLcRNWt18bdmXEXkvcvirs7spd/sIK18g6hJwCvc
fBsxqMbKWwQafpa19VUrtd88U35+bClP6nNTJYqm7InEwgUPxRgQsObrRcKd
h8+CWwRMcXBX535yUqWoNc2EKFki2O2vb0BiVTs2QtzxKddFCwD3na8u8dt9
CL9LddVrczHp3zLJFX5s6CuF+rkUhiqHp0gK1tXTYif36fLjEkHaMjOK2p4I
VcR5PK0wB4hUzaD9N03MUN0OG+qEwQyJu63a3yUXS3E0UcjGHMwp4wtkIJZy
Qx0kgTbUhUjsN6V08XsU1c2aCxOsVYcXxQKwPhH8syw+1/6L2Hx7L4bLoJv4
1zY2rudI6mmW964air7VzkU9SkRFLavb48sYqMd7Q8PJmAfS9i/DyTHMNS1v
9MHs29IIRHjorgo2RClXHMwjlwXLa46gh/sOR6OuLyHhaXk2q++fJXdqmkif
XnvZdzUcZeW0OT9Jm7DnvarrYc7CemNYfCJTgO1pq/Ca/gK2EuIdkzNPaoRg
pjd15lyR43JLfcoc51e6XoBFiYjVrr44kAhN2eVcUf26DayE6J9rHGq0rjbz
4d8H8kHizL66VhOcet/kZetFD/KHi4WAs2Cyaa2Tjatozoq8+6LJKRvOEevu
Bpy5nPOfSE547O48oP6NMQnoH5JqtcMOG2a/F4dCnHfr8YRLrsEaBrw1v1gO
+EQKH50UdTO00w3T/+xpJvuCfGtB/WmYh6YTOSLr4LWoY+40Rk3s42ofiHNx
MnWW5ws0AthcdO/AyilmgowLIZe5SYOUgnJvfxG3/OkQ+7gQmHNhgaaJySOp
5T/qzwunJLQNPDO7JCys1l3v4cOQ3Gfm93sq2wq5AKQodJugDHCpb5Pi5iSJ
jMB5av21BVBn6/POqKk5HO2A9FqJfdm7cEVl2PNynjH0u7PZl0MxXRd5uqiK
ZfodXA/z4OHpr/uNWqIwdyujOPXq41NNs4XSoudVco9oxB7v2mwpMpNGatgP
M8ZoyotKh4UTyNiWkOS8FOSjgS89HYLLjmvj1psl6/tRFDpJd3h5exbs2RMg
D+Q+GxaE8dgChaGef0vCEoTpjUdBniofzMU445AZiV8LryxaqR8pPg+ghoW0
YZh4qNIkYFj1AHKGkncb0sUoYxso4eoIzx4ETWroaHoA09LDF15vp6Fc0l54
nbuku84Xc7dAMPxpzbZ9h0uEs63qgYx/aeAVLIinqY7bsxo6Yki0uxEzhWZB
xWwF3S8IXRRxtVX8nVWJ69DC97hTTip3KLetfOzvoB1TJTVHSkpkRUugWsye
hR2rbEmzk5o3tL3C6rK2xKBImhvj+1Mq+xQITrx2yoJsb4qjz0iFlLWPrQgU
6JzzxK+noTPzSk23On94pJeq6J0vRGmaWLt7s2rA+ducOg4imDYakSZms2sX
Z5PoiyZtsPHOrLnOfBABgoLjgQGZKSpVxG3VlRXdfbzsvJ2tRj1IWD8m7ufX
usjXxUWaNfasIG3vGhf3DSaSGoQvDYeKxrYVLUuFmIIsL9LUYMUIzOBXayjg
RDO6T6GM5XvjI+GIJS14CjGCLJH7nM4lnDRFXRkWWO/xsOlCR6uR414u88Va
ncjEAQpwrr78Jbj2hnAW6oY2BCmq6MOFa35HSqNGj6kAE+uw6ubS+GCTyAVe
FsF09905+nwRob0K7UQ8+56k08xtlsge7Tu+xpslDd35y3j0gjoSMw7Yj99m
ogxba/p6GdkH/hUdH40uq/9bxWrLkRG5Vxwo0gq9DvK7B5UNx1pPaHO1xW71
k99DXau4lGRJ26PZb9wt1rRrdPUrwkRZ2BxvON6N4qVAwYSJSqvccrPAsj+s
/JfltMnipWcRoFlBjDMGNhWiTmJRI3UmCNtpBJYGuBxCa6yLsVCIkbLp0qAS
EDl56FaKOh7ngoaNUpIsHiAjwlrn6WskNWhTS/EBCyMcuEdlVPaO9a+ssK8B
/D2ZWxcwApnonBF5tE9WDqsrHFLNpCSu0RwnLQyIijrGJRhDI4pdbwlK0jbB
zLQw8WmWNp2iHXIrpZNWrbrk7e276eQVsTMcHJPR2Qc3Av9QHcz3U5BqvfGz
ArD/LKtTOViIzexwrsGbYLdrT3nHRFUw9bm4TRvac46ZECalI0MtwmgTqiIf
L/QhrSjj506wXisHjVjP/PhGTf9JrnnH/11EEet1au2DK2aijytA0CNaeW2E
7IR3GjwMpoXlGUgfdQ6IjEZA5X5Wr0XnLITUfdi2w3+kIykLTtduZQxKnY7E
90PHql+LnCQQub2R1OOK6p349NQI0BLTz/AbDgHyW5+lULKc+X3o6wyKUjWz
fcbgrCadtuR7CnjaEyZx9W6W4l/zOoy5WiyoUd+OdBCp/sVMIMPA56wh+aj8
1+tQnKkoTW9Ck/88LTCaDkdeKB5Xfagbz4hLBWd824+0IgPqY1aS6L6Lm1Wj
jkhzmWmDL02VHQ8mmDVT7bzUKBXfiOWQt0QjRyJH6As9VsJxy1h9z6Ly7QmE
ZN2aDjpXuOMlJQRKhacCtpmyDksXnARNvSsxDRiZMdQNyfsGzzRLo3YfrKDN
mQW0zxVdH462efSA2Rv54xp7JhH1VS2eS0m+Tjod1kTf9Ph6mIxXoKiaohFi
2mltECH5j2TFcNNznwzi260FO69s0UO+KpsOAg9dtgKycPReuD/O7HcYZk68
E70pyVwF5GDGhYzSTmcGRZ2uL5Lu2EaV64R62xm3LbqdDGr+bCunqJaLR4BR
caxQXe4VuED3QSMSgWLJ7FTfkos2CTwCmd/s3+v1uBwvMgoMzAPunHNZbOpq
2C36BK8bWH78wt5RA84W0MmY1wce8CStYcBtvOcVGsZ1RI1bHrMeG42wlglp
iyxFpoHDlkvxRTR3ahxvpO8wKMeBuIqdH4S39fODDA/b8ZiBEea/tzoO4YrB
sKP2jmzOK+FhQIVGPE7X2bJ9sTRLxwbKR7i7WpH8xnycu/aVHKaHBtPJK2X/
LLiCCH5pCnVyxjN4BYk1NJ5HHaOlUr6pxj2usIc2EswkkHyG9hhKQqmxqpWa
dHKyRzxRZYO4wNzaKSKa9hzf1HOLqmV3+xFVogtw8mnyjQWVGleDpU+ZZ363
dystfbTBBWVdERuFsCCRFxG3+ewrjL/ufCS662unPJHfsHihN5sgsrke/9oQ
Ho6c9rtUq8l/QL3i1vutEPGWVa68U0cIeqG6G+rOyBUM0infRVabuD7LoODT
ckqUxnp0N5o7lvVgBDl5po2la3a4zfuVwcBpKWW6IezgazROhcguw9j8mj98
H5WgNK+aCNL3kvqSGAv1IzWzo83y3xWhgI3uaO4GI2wlx1S75kXmHsfKv7+w
AHkAmf3Xc1Nd3fIpgvsqwr59avDBnAly45fdP+comscwjVIzO9FXXHwNKtyo
L9IkZZZPIzIM7Tn8fWF5vECb1AlrfmD/zfs3MmECRaqsB+mn0/OyA8pEs+0g
jw6vKBUoL7/KHVwndcw8Vdxu32FPf9q1wJn2JxtzjwXPsdih8RCB/Y4MGmqE
Dv3REmPvxdcr1xp53dk4kaR6K1ml15xjRc10t6hd6ThRoa1CHrINJCcbTRPj
yXrhBr+7yKPrQ0InXyJgJKGYI18P9rNgGQJZAZx83JkFWN8rn0tXabeFtawY
KHHMheXRs116avFzZoIQPzXvGJFv6w2KSGN6AImRFO30JzsBvHINJ2EHwZSz
/ckaK3+8ORyRTmZV4lm/5lRc9Tm4XL02TY9UqSP76UsAXSsOmsadlLp1JnFC
BeJYbd0khtC9EZ/QZU9eLUIhip6VvVmSKaRZOZLZP+ZVrHrqFIiqXs16JwJp
F4/EeZfnChycMgg5XXycbUq+bKfrlCf1GjuM3LQzPG9IeOdq/S3VNizm4/8a
no2VxxyNW06gj6vTtSeZ2HP1URkfqVemykMY/HHUKDwzQGmLnhUD+AZWjJ4s
58tUWA5fdUtVS8t1EElznjHluT8aYYjRxl92iXLGpZ5a9waTM9dLghJIUYHM
tjhopwj6VKvM4+UFpgYwDu8BSOKVHBPAW//+LMrwbLOMTsRTuMNOQLxp6Ot5
/6WXpafLmdykP57rqT2kTq1q3rysi3A0/UYTLezpjfEw+Hv4oHkICmnk1vsd
DV9jA/FTsYn7kygDig2B5yRuycAGIToI1e7RxWufg+ZUOh1U/2ApzhOEl5ij
jPp1IVw16yZsy+GPEz/a+M3dqZB0Sp5rUYUEWtJndVPk1vJLdAC4ha4XPNQr
CkAfjR9TKxu7aJ5hh+wAhJ8Mu0lAmW0z7c9yLDI0oSGPMGLVxuS7I7YJQr84
eEOt1TaPUjrPEOXLt2XD5unLe6i86a5sk7ZMNna8d+Sa7ndIQv3y6W7c+fEv
iCSMOLf+AAosmyNHnCDRsA/t6PLBOhgw6asMrbr9OlirhliT/3h6U3EE6GwN
A9fOSFSmkiMF97ZGiJuyahUNc/5yz8XCmakVpBtganngq/iV0+8S3pcMrkz0
kGGoFEBFVeCP/4B0ZkcvHl2iw+cZTMpfD/QfSDTEiFdNHs9gcuqrJXJKWNU3
soK6wkWd1r0xQspqt4LtEJE5TWh8lEaI3GL6+HLFJ+nbORCUK677wogck0S7
+NASkXnQUYdxzmuskg8IvwNy+LGZWqGJAWU22ZNRmMUyPrrhcipHyBU+MNbG
wxzScnGrFM+Rc/RSpO+C3Uv2ZxEDrw7ItdKsFefFrPW+aaFj84fWQPvW/EKv
LoShya/XFa/IWDbReO2SWABLmq3QmBkBwfoAnK9fBsW4xPL6vKyFn51xv2lA
puY6qmknmfTWIj6w6iKnZBsczcXOFJ970k2/VKWjlGc2y2JYvJc4U2rhjCrG
fQeNLupZHphSXmauOQG+3bJvrfSxybc/8bgp0pGDRb1PvqUkuXpEBCzH+0tf
ajgkADeuYSJF2toc0i1XpfyWQoMmtlt+uMPk7TXNKwwxlWn7zgYm1+MSpy4S
pdqcAItKDQYBBaIYmi1QXR6cAaJHxpMiNg9hzgVKsj9IGUzn+NnSX1XuG5uX
o5OX/v1uu6xM3Fa57jEEL3gcXCqzQqlnH1H/Z+zDvfwQjSNmhobLYbc6IyTA
CRoFjLYzONZ/hopOZ7M5PA8Xq8SqEXeh8OXRQQZd0ys2BvW/zplbOy4BaepV
ceq8tEnQsXoCPVkQthf5GgcY4sqY75t9gdNB9aoZHFY/aPAKqWgib0BVpVX5
F0cyHbMxidNzTOcQ7VKkKsNkAzp8SuV2YEt3zHCYmOAWcHm/p7OO+Xt4esMK
ywUO47BqkRDGmNlRwjlQH0LG4S00amVtdS6V7VrG4v6hlyz2x0fCBHNxMTLP
v4R/chH19KopD1RLuFHPQCevJ7tSXjjo2ZEKJp31CHnHODIwVb3HWDHGgYZL
VZqXczcYwqCsAD1hhaoHnzeWVuPFuLVDFCJVZM9k7hVSRCMF9H3SU0xaVV17
2raZdg3ncszUu3CCy/DY3H3flKQqUOl0CnzYEqJ1rSMXhwx7u2ma/ASlZIHq
+9sTBUhJMHeuIOkX5aRGKhGFSWhv9EJdtsjSpmQTfvHWK1skPwociqiKiuA+
l61s+8AvKn8jiJIuU21DnAUc5z6mKzJoPsa/8OFQ+WULPz7zuFTPPSy1QPdV
LjMGTE0jCG+VK+KmtYHCwvXCxIvU6kn3RpmISQJaumCZtKgdovouXttTnvQL
GBJP6DVml7U2crPreKbSNGMzOG+Q0BD3IVbofkDcg87LIRF/7IMIcldfZVUg
AIuqxTd5tPn9aiIhtSrJmGB0ezgL6Td9REqDGygIHFGd4Y3VZWiq/XClq1RD
NrfdvRAjgYVcxlFVBuaPUlOXuMi0MD6+hmklGMfdNYKu7ILFQLo21ATQYsT5
GSEYmvYGgUjK4VyYdWmoPqk5gbFgyzY5pP5YJUSccjFyWMXFnDaoUhlHM03P
te6M4IDHbznJvkhOsyqYZHkk0ASfRvoO0UXkxKsA3oa6FpXuqIg6Y5Wm2uWC
X1/VsEmgQepMzOXfYxurYqRgAYtTzcYLz8I3L0euj4dnGTLaRI3GsMrnNP0D
Gn4TqNFjdM/sw2plyGClVbAnL3ikUJsS639oUIYjm7txGffB/xytrkT32qCD
88GidPkgNX7DHEFt8gOyQ+61eQktEg6yBqbCANpPyEKBZ9tsNMmj2Mdfa6p2
Qdvg9MbN2vBotfuMbYUn8Ep56p8UBEZ+jZaDafLCDLTtg8pTOWPO2gDd/bNy
nlq6XP+phAQIzN6vdjY8L34HTuVpu/y5HXCacR4UMbkEykRS42lMSE8PGyBv
brVYKbe8YjkpPA83l42deV4wAfrkJpwVXohFydzqg2AA17FM+YuqU1/fn7g5
MAvu1qM8l4GHqPq9QUa/jF5SQ0kOcA/wLFt35/1fUc71bQODa7d+htiiM6s8
9ieix3vcr83OYQ+RFiduJ991rSfG7uuRFCIbDgmpejFCOMuJGnRkUqzIv8Ms
XjfvutSNVK2iUNAkOjRWEKAMVkAddMMht+sg95vOj/tFFcgIzKPz/43SD8as
QWJ5WNAwnCji8ii5FPFkCNHqhbr7zLF3/rPOlM/ame7EsNO63CiWUClSRtpe
XhmDLTbYgFyZ+b2HbIoIJoNtF/YVhuLIHSLrjSBy5WfMja1wsXL5g4QhvzwE
kNS1vQplG8Zf3+wBR7RRfCA+h5U8QSfbJ0UpPoigR+2NhOPj/rRrgSaIZ+eo
72Yep7p035IYrV7QOIYqs0pyIzl1vuB686P5NcoygoZELr18egn2z+FBBPvt
68Utf17b3kG1UOCZQBNlFGECv2vM9syD2C8GA8CCU0wj9w8gf7R13EsQcJrJ
79Wbt2jhe3betj+3mrmgrj16JMZe7Q6kUINSPfwjms92anZ8RAvQjR/nOm1E
LerACZgMfk12RVfS1dhk85CD2IV9mU3Q8XCds5U6oChKUn2hL0Qnl4xNDhDx
CgchhCxZxOBPj9tROEPius1YfDdWw+HjqO+kDFowfRbJoh8IFdJB/P/veVr6
KTl+Gltr4UxqsfggviAc0P2MkGDpkicgGGBMSpWrKa1CE4+z4xKxxRUnNSxv
je+r3vStEDLc2NCKXdEb4lBy/fo4RQ4pH7nTzOhM8oVIpqW9j4EyKqqy2iyh
gh47R9XlT2LyxGWY4oBqkhGZ1O05BgihyDwWHL3Mxyhpkcp6/ajDg2iIuDYm
lDhhKiiTnFJs0C2VGFVDbtznYH6Wk85ZAg+YcnrzsRN29dTwbpj3DiCsBWWh
qZwaSAB1VAU+rSbQkYNn9ziq+AwkI++eUqdJjhQ6In5EWIopC52li/9zQSy7
LRns7FKgE4+ha1A7ygZl5qxA5cYMQBMMIbX5oHlktdmhiRxgNAnA0tf8WbnW
8N2cMG4BmJuelHptJ33c1Qsg3JjnkTUmpSbwcz3/oubtaNqPWiTBtNxUM41Q
bR6wJYkuHAlJr2B+2i5kbO15EaVZySkrryaUi4cd8UkaumnRlXMp71rJKgUf
AIB6jr+8ZUFRt2briTYX7DAl3A19v2qSWVpHgga4bm0oHYfOkWuj7xr0GQdQ
RkDvl24ZG0TBFh2746KdHzQuDGoYS3Ow64gZTWpvOCh0cPLyCMCMfpmiGbzi
kV3qpqapoJ1+3fYMH5rpGvYSIHMyP2siF5ahTQmi1CvdHKJDn17EDg0QlPyL
K9yGbztCX+UhlDK7J3XIv0HBb7AhXzyYCl3mwQJZIp/XnZgWXsUrP8gzN8tG
uyIwonqvSznYnuTrUt3h+hi64zZKvaZXjPZ6zcVHUePGPpng+byKfH3LUKCm
fdFGY3n3AKMOD3bish+RtqsZI3y23ltsfnLZK5BQwCzbpPcRM36JBre9Jkx+
pRjZPibnvWtE93gKnmycv7EoXs45cSP3PI6fvSHonlHU6fDbqX93cKdwPaM1
Kqy4pZjhuvcXGnnuoYOFctSKNKmqNCgaCpmoMKbfle5rFHuL4F8F5IwUrDRF
dLXr2fNT7BDTab+nm00u7T3r0Jramu+zFYw6dTH/wACS1z/hAaxNC3kbWoVf
IWKm0lzA0DI4v7XMLooclpSKtoGNVS+MBR5X7W7VYjvt13ly9QTTogDlAFbr
leG2zkt1VnJ0cTQGpfejLlMFndxZpaJqRb+b/oEkKpmVaPwyOtovxEbzijG+
63X8Stl8zN8jf4qQgTYKJTM/vFmyK6letIEN2IKaGkQ6enRDF7bkqGCk6+wV
yLT5R1oOq3aR4cao4Mn/YOhrXNH+qYNz3jBZ6yoM9hltjavCKqfcXaC5DqGq
mBFU+IGXzeRdGW9g9qgArwK8bJWQ8zjn9WQsAfKBZLi2Q8IILSC607CV4vDf
HZNY2aiL5cvPoRWSjEEsDrRV0Cqu+EsxEC5jR95/yj8+nD7PfobZl3C4wkiU
py/X5PNZSpE1mK32M25x5o9JcleWsFQR2fLB8aKmyOvkqFKeG7GRrnWqb+i0
+/mm8eMtrvevgU7xdAuo8JA/qPve73jKXb1caO4/uXn35zQzBWJImN3iqZL9
A2MJUiHcyuqEIljA0RFcuqfurS43+a76QvmsQ46t1UhZJMvpagudfCGiPy+O
G7lLOQOtBq+RS/Jof2iI/HEoYeRy2XsLrPZ+xEOSlBwMKVPSmmwFGA+Vlruh
qBFXmwHzqjY1+s4/FkBeaysoAxP3GY56kUCi+RlVW50obWuT2NylwNvPmyRD
TMZmzHYwIJQUor8KzZXc4k+MTtbXeOXl8L4UQxPKYXws4KCKiVVz38YwGFsp
UsbUPjOG7/NQJAbsV3QgWA5WpUCN330DWKBToRIFfvCU0dPzoZDVPuSS6AFi
uU0a/D4Of6XTYiS+HFIWmaomrVJFPArmePjpMzpyPP8RWSiSwIo0rnnQuPr8
3jGSPjY6H8nCl6WqBkUlzA/gLEmSoMv50YRpnpXoqriwx6N+m490GFjY3dTN
M05BGnT2QO1HRe492iQkzofnMD4kz+OCkKQJjFyuOApDoyJvICl/EOiMJQ+P
hvdO8H6HifiQ9K+JOjVErGK4ruj6gSxlmDCnt+lJKItEnufVlY2OTv75eBUs
PvIIVbmOUUkLy5Zfo7fvzWyvCURDYdyZp1Z4L7eTWakOnyqNjdKJDfDcp7yw
MQBIH9UbvHx06Qk4t/2HVBS72wD4+Rh5pJHDJE9CcEbZkmNv4XkJYNVt7PvE
mf/r7CvVFvGgl3pYv7yIZc25HNjTylxj25l6E3QujDC431wACTE8ZdexUowz
Q3FVUqchKkT6OqxMtjbl9TXvMgwOaClVworCb7wZbsWUNvzjwYL10+Bs2Tdo
W1FkxBHS0GLr9XclHGkjIfJpsxOXP4yaFrdlSylJLxq+3jmZUC5k3o54LbhZ
qySDu1V4xvC+j0IOBFVta1Y1bGFs4Zneg6RXxX8fB23YKqOChgu7jCg8GJB8
5geCZ2/j/y08SnuoZTEibbtGyesMhyqGuwrnzhWKltGagLdG+zkxgzk2cZAF
96syQgRwP+6ihVCPWNNYAwrCCRXohAta1xhBobM6+cVpkg+s1o7Lln767kwQ
zwruseFaMRsnW4hcMNnbNswztKbvhvj6EhZ9IegI1t1RGeOP+ObAHxVhUvGv
tO6ktRqiBitlNGocdOy+/1iwkhY/CMzB7mnS+WvQovhMWBWNIO2NobIyv1u1
SAMOXPGGJAqXfIX2Qp89jeTkN525/txm9wjaL5hbavYEjJNIOUR2us+8sTIC
/xO6+IG4okkt0utxNUeBLDwgNC9G2/6qg/3b33+FElKebmNNBOTZJVUAnNTm
pe6sG01y56/77duISrhlFr5104Db1hdB5rOU1FFEQjhFJykj+Ctf2y9xJk9p
A1LYwwrhN7R3nBYdBsEaVMmDjXUJ8aOkMQZ1quNIc4c9eQ9i0UxyR3mbEdin
lJwDGxrQ+ArBKYOcnRtGLdBBRqUFDpYQR5L0cJF+BCv5wL6r6BBgSx/V2VOQ
6aiNCHk3PgkAh+4Qx3K5/qepd1D4ylVxGZP4cid468LlOZPkshoJNvs83dXX
knmTomh6dE/pIF79uNMT0WS5KL1evMrD0wxy2nHju/jk62bfZWYLhkuNK1jl
VtqNN91Xa7dpMh43cDZEAmDeHSBLC+Q0i2s2mBC0kcTV7U5NN0XPNMJ0sXAO
6DJrro1ctBm7x4KhC320lvIuSFmF3BDhBhw5HYbTtCFqG5EirSznw0pWKpUn
CjjXABz+zDiZcLkpzAW5HXi5NiGFztZk10MJKMNUG2KI0dHl1tyrtFxiFKx8
KzlAwJD8+fgYBeFRL+I6YAduBIncHJUiEup8S+uyO4wiSiQ6PqcZ/uXSjcCp
5iCUYDKCOkbk9BNGF+ZdAtRXG6K+TaqRtNbItwLHEx+DG6HBmeFiqnloIOU6
ecQqOswlgE6bKwggzPpR5gZjfVqJoxTRVKGmmDiXHX8GM/97n5lDc6kTJQF/
ZhrmvYV+nzOUaQeFSJb131chF6JVoPZ/+/3CRVdyxOHT7Ey03zgJLAlDCxDn
FKDYtP5VElK1vAG35bDhg90nZmdNnx1dfe1CEz3a56HAdjkBGnRJsyjSzZOU
uDHKlnbf8+v2fHaSldwLomnYfbdHWsTcuY1w+Ml65XrOwK0A7IedvaEvb6Js
FdzXLA+BQ21LOdSt57x/n6QeZgXVibm0gAgACjxNKf9CGpW84wrxyenCJH2g
ePEXOv/BBAZ78TEx2yu+iq/adYYTXQpvtklGwFMsrcbF4Z12LWwqfsWLH5Ej
fgtuo+bMub/QSQ2e9/NT276IoKX8VyRQ62ElDJbJsX5x+vX/RazUgmysPO3q
227BZ5OoIjBTTok2vheF5Z//Qh2DZvjlnq0PfQ5W4VT/rwLIkU1yFEJ1obv3
ci6iQsfZLkFQEeKi5IAD438+VTTW3VKLtuS+xi0DJCvEqs9FlS2UlH1EMsiX
CYnZZ3cArLtUJkkSLg/ZttTzHU6jnaYp4PcB513Kx2Wb9McFf/s3nXK2boiO
cJ9jJz/ar1ikwFMTOwQ8eX2I3GTtFSVJc6GTkOa+FDPJFvBMIWpVDva0mM0a
wIQ5/Mb4ryKHgfShdWAFsJBucBcb3W/9f0LduSvZ/ZwcnUPCDZnrbVuxN1xt
o3nEiqAGF5RAG9e9D8Y+qZyVdS8nDsQZitKaIVIZGvJVP72BllHfPHwy5Z3o
Bq3dZ6Vg32UbdJX4KISe1Ep1u/PZkLOAJ2oJEjptoib0xBH6Bv9vp54iC1O2
yD9WOtBlAymx8DzC1nSzYOXx8+WoGfT49pN1O45cw5T7joT8DoHiHF4QPQfr
UHUaXnXOmpQjWLB0V6YVn2C41w64tlVSdGEMels03XQRHjJ8O2YWrt7eki54
5yqH9t3KQJZonKPCDHZKrD9DtNHF1DQdYdhr7dKxZTQEwD/bJZysVZWtNiHK
/Bwr6JIoxM70Cqtz6gp3XdKXOnJtesqIk4NRpfuzCZQVXBtl4QHV77DGmd3a
yye/muR5dNnNXUwy/zJUF/8QgBQOMdXtaAWEejromF4Tmz853KHI3ZEBxBXD
0h3xuTUwLh3g5HXAXk5qid80t4ETdJNw6p5VjYlV9aap8KJZSFQS+weZsTmr
BhlygwOymo+X53/HmQX1eIxU6XbNfdN959QxhEYbP0egjV2odf4ZocgLyx0N
tbwWKVdnRjJG8EYsJujV8YNVEG/06i0Kz5BBSg0rJ4o0mp4hGlpuwlOfHQmf
AC+Lfo9mryhs+PLjN9YrRiMtEjx8DPtDj6DsxyX8PpRqq+C1k9UQZHMYdZui
3d0cwG4M4/wPVMj/2muIGg4q4uRpQlG2Tk6w9SM5TQhncek/vB7dlG2Dq9oC
zzMJCFheAG53bkRVEjcy0Qs2Y5pnsxmwvadPHTjSlx+QQxak8s7C+eBhG3Ar
3E30SuYmoGzVrHNLY+DWN9UsxdxBUWfccWhnV4Hp0CcjiXjB0yBbRGdWsE/o
XYRt8SwWJM+P+q9rRb9CsryPpEz+Yo/nx2Ot1rD97nl+DORA/yatqWC0Pj/y
slkFrFzsgrd4bjBC7IIltkgRvmPEIjsfP3tkSVWDWKPDwT7c6bKmuLe5yCxV
BQnP36JGnNK+1YvMJPqq3ax71d29kvm4BIQc8EOPVUKqOq7oQ6sc2O+VRQML
qy4RLxJt9O5bxGG/ClIkzr29zrGyAAI1rCsEP4R3DKBjA8RCKZosZ82USIJf
52A7EA86/NJPT0LoDEOEYHKfNxUe3ayDFrHUPWcDhRDBQsGonHWvjVhL8pXy
YRqRN1uBoODwVV0hl0TIGAGSus9lP9Kbz68im5qQqw1KicuD4B03d8Vms/xn
8iQLiVPGZ0JMBhltUAPyAhbyLQ0oBOpjEF+xQD3Ze5gak5fYPcCHaCLbYa4b
W/dCLg2cvEbHXBe+3oWhb4prNm9pCpDANjLC++KrcTvHxFsB+XRhlBlCi+tT
XHkfxKThkfXgyB83yBTXawWf0lySM0Hxr5p/Mpnx6jOq/u4Gj7pEZym2o8DG
CbuOy9erLy0U+v2v1LywKZGBJD/cs+07JKDA6AqJnOd4X44OJ2RhcaYtHAEc
YiJwTpBtNevmXBa3gX4zqIok6sN5vl+bJBieFpvNL7Os1okcYB6PaUtOqjkg
TlsScROkUu1WF2BooU0l5G1pyfrKhMpz5oCe6VdmZ/Hwlq5HwPTlhVdEuic9
TjLbFzkmOnbL4REfRVDFVkN0n0NC9DOVfSnGiax5+ysc0BE6AQP1FK6AJCM+
hG8re9cXn+IMg7MUsQM03DLLx5to51Zm2r96/y5p/Pgjg/EHqJR+Gb/XmjER
bZJzKiDesec/EzRW+HP0Z1uvqE3cASebyMRUcSqYzyBaUDWY54rK8QO8PcD7
P24DBF8FmHezZZYoG4yriKveSxaYAtmI3nIZ7K80tuVNTWUDfzWtI9oV2H0t
Ozo3faKsec+9aIGOHxcb1aHXlOsXx7sGeMeg2KLekZcezBamfyQNBZxZAdZu
ZHan7nWV9P5g6fVZU0d62sAixwoiKornowlAxmyO12BYiGmzxXd63ucDjID1
EwTtjgB1KqzZYLMssv76aOAdlm3tMpHviDr/KBKcIP76IBkzPN7+5o5ZmFr4
F2brNjpGElSlvHCsK4QGdJcdI8ft5OJLFXK02lzDb4x0yU4HkVNCzwPhJW2J
XlnSdpyxNzlJpstrW+PSc3p7AXIE3G0ELkBP2/Q+dohgCElRz8GPXtYoFaqt
stVNSAF4cin4JLcgjr39eIWz5X7P8hyN9B3LGrRwxifIaYxmYQD6b55Ieab+
ASIlLPPzzQy4giwLURWQ5S0DvDMubDhC+fXmYis1VRAzLljUsh1HDsNqEAws
iPBOKH8QHIudU4wEUnK2ai3MaoCqi7jZFEuS5qi1zd6QRYlDNzlt5NP2+6rv
0mHqca7X1C54xnGt0PXI7JKMW0Tx3NvVcJs/ktTQGKJqvK3/Cd7+lk6w/OnU
uuOf9IJ7SI/OTKIV3W/EXw+KrD1jBMVeJJjBR5758HqwVwUOSRs2bPjT8kIE
D7aUrRRgt3XLxP8pEFY708LguPn+/A/vCWVayJGqBMF0qVUF8PsP20qrdHK/
eaRyXRHL/J39g+YCElZn3m3OntxhFecOIZSu0TeBmVB9GUthbyvT7Sg6bhpp
sb21IQUht7vMAkjEV3+KydPPPJJNc38rdUm5lyNxP6DvbQLq8SRIpcqb/bj0
spYiUT5eBkkZPmcOeCRV6FAXt2rQQPg+9JRlRXc4BVPJvkCUKuWq9/lrDMY4
W38BG0iA28YTI9Kgi2RWwpy96K25sVxMJL+QlRwRHl2hcAU8i6IgEUdY/r5p
cVlyWH03ffWpWjHa1uOsvzXUHH9a0VW6T9/p8g7VVSeEImCUpdlUW5Kxrzb3
Lnb5CnP8kitLOOyYc8MJgB+RMtGReJSnGaT+zyUIOBCHZ7LlEvuxonA66/RM
HgZP1b7ItpFE6836zAaaNzXC8U0P2f+pRMdsjH+VGgLeM2NqCO9xQZxsQB7L
+NZ3PyDX/e+8i7MrhzPwiSKT5apSjWO9av4VhQYuA+EPUt/VsRUTrBvOK4/O
4s7qxrdMmoAh6/BoGFEXQyyYZI/E+5U3xwSly0kju1/dbJTvCnUckL/qz6SG
cOVBoRMGcFjxzTaaLs6Cl91yhRvwCAM1DMpCVI+1IIRydAODuVMtpxdLhxIY
+MkM0NQz7Td1DzJNEoYjxlUwMdHsFND7aLEfcZQBti+WQfzfkTp+d/MSwQKt
+SlRWljkJ7t7F6Ug5ZOrw/eQ/WFN4yGd5SeV8GMJ2gglrHfUAV66vCOELteL
p4RVqrd0KTdOg11/mbmHGDgHjAWDxQxH/bvtqQ+/udQLdbJWIe3wvwd0N469
QDAep2YKQv+QcXuInAvRZOHH5rfUFpOIQNIWMwQA83tmj2FHQxA7AB25SOhe
IzvHjg6yveeNAyKc0CbBInYKJQx4FCXUu4Shqjj3KYVsEYNFEvZNSnXk9Qaq
zEEezBQpb2WqJ+GJ/wtN9N7fECU3ZCqtRaMQXJmMwB0s9JD26LcKjsncxn3b
kys3O3SI34M0RBOA0V2Ghlyeyfj6ZLODQnmGG4vujlBMVNQ6BS4BZ5PGIzFp
M+lJy/K2ntsQYPF/8BAixt9y33vitjHBXe+IR69yfumL12esflwLTXuBIitz
miXDXFYrIpKa5Lx/EZQIyJHWIkvkTqLMJM/Hu6pzs/ULbyf383YI82OjM4rZ
lDCyoiayCqqSmgMxCLmwLLqPSgqbRdFTQ4YlGlCpzaF8L3thIcDoX5XGxMNE
FP0ukEU/AFjx+yHINgUEyVg00Za4AxV3QFDK+obiId7Xq9LQcbOYxaklBC+8
bua7K8A2U2kdPLLk2gPR+0S1TV7NegfiHT8pf0nyBWOnA1GrHo6/UUss9XQ6
OVgceBM/yyI4h55MdvsmnMCiPqjqS/grNM4rvx2GrrdXbC9osPqmT7vquVVv
wgt3/3YPprQD/1okKYXb4sAMXPzVCVmATDFpq4mL9gLrveRWQ1JM9stSidkp
if7YIYnsI+1ifYxwekp+4utz6GkFlTNroGvjogtUWaPqS90KPdbI8nDJbeqN
Wkv9dCwI23Cv7UN+drpb3bArmmb0zyI15cyR6Qh4lgcW7LFe8EOJLrMkaxcJ
0AOvdNlUm5eP3sBissfzDVr+/cDj1m0KyqOGiqiDodGCklR7KCyCt2Z7G7WZ
T3x+FU2IDdkDeCiEVpTyKGNYUb7kPLY38K/q46jItVcG1ivE98SxbblxZqEJ
btQeJKmPm/1BkPu54mE7f9QrEh9401tM2gBGB938/4/qKbyGUgAhWdo3PXpK
3pt6CePdkUluorMXuCTUrUlwUw4ccO+awT4vEwgGovFQTI4Dh93Ub2ZllJKl
qVMWCQbjGWvouVBCzMu+e5qsLTtm+ZrjFbGMKvBWbNMpY8OJZKuH1pJXMng+
XeQILXlMQ4ZavJ3BGEah5L1vrvaOmLDbJ0aWaNLHKmWp4ugosigbqZtY6U2E
/G0/6tsPCSUTd+dQAxsSW4W6YDiLR6zyBL9KCv9WhVc+W9qmMdneCv5FIb0/
TBpsGVbw1/Qak1PrFdU0NFrCjkL4xmztNFnpRgoVeTOze2tiAKgV3RUgML9/
oRuZxaqmygiHAKohIa9Ae3mM7nzoThQU/S4AhgAhFfVeNtAjXoJfDDAKsTs4
E3jnbRAJWpWTZGpQe9wlO8G0PPdMu1e6j3CbD7GimrU9y0GwgksczZLSrIAO
UTrrAm7NDgYDj4vDQFIDrlpFIjKmFvoAStUyGnbCnDtIzQWd+GNoE3HWRNHR
Sk5I80tIVh3Ntg6TdGsIRY4OZUoDz0nrYHZHAmcNoBolciktGhxls+NX89q4
g8XwHNS/v0MNxEORJrrY9FyR97y/AYJvuXjwQjxwKMG2KxqpJkemeM3JjQZ3
Aa3xLadKkKjTlP3c7GiIk+3jcBYD4RLScZe62yxdEV6CcplJ+dE2dkS0yF3C
yriSOn3zaaqnRZIpApVOCVKOBYSlyOgc49tdCne3ovgbfp9mZW9OXL3K1aEU
bWCwjKTrBl21YRieT4Ggz+HSgeiNE5skwUu2R8E61UiYgmof/uJMLCTc72NM
NtaGsNTlZTKERkMQLYQgAmBlYZtw2UHSv56J9vb5aaOniAF9WTrQggCQ56HT
OdLPFb9VyE6MPoXzl0UGtaxNPwsBzp6NYZyo8BIe6Jc5qmHF5tbh/GZIvRJC
bF6OqFXPhzOcKQiXQaUmiNJBikfmWWafEU51gVycEskMcnC1SDnlt4N69DIx
Ihk4EOYZRDz2rtjW+OirzWLBVtvi5sE2X9LrtbrSG4BbIY0eAmZOCaNH/SBh
DRbBa8wxkOU5MujiPPTyLQB5q7DE9Ac4d5XcXfU4X/K2Shk7ttcrgo5vq3qR
wKA7R09iNvd+nBrIzcUFCXukYuUm0SVCyeX9fqARUKwwEqSE8kpbHAQY3OM0
Gyk4dxsvqdexBAVAB/NPlwZbHLaFM1uceSrrtHYHBSu/aAQvYw+bOQy2dAvl
1yZ9USs5KeqTtS+wXkRacLJPfj4UWzkTd4ol/Lz8gLLxCDzd/7phKtPx/5Jz
Ph2NvBydlXQBuraO0n9Ia3aNMxlGDbxPcBKGB/rOG2izyxk8c0ORhHzvElOo
wKztstfvyhVvyvRnqow2GdNaf7deSCmBCB4ZwmKP+r9YvCHBTmkIXKFPvI2I
Qt/NTYTfqxgNzPj+5//QAETCZEFjBgCvgmu5UfmmEqDukqxmpm32pvwZojIT
mtW3KaIbXBnGiUscdO5WHoPO/VjCEP9u5pOEta6nGENxPsV/CZk/iD64OWkH
pbk14qVonz4a/TZ9pnaYK3jA0mPDWmv1IUFjafdSWTvAqmDQ6S1J79RSmTm7
vOKIVW5CYdQAC4/7TTPGmqOPjJNMEn3Kfe7wEgf52avaBf9/rMMGLhAp4VCn
6xgDFAAxaYM3r8r1Cc/HKMcxvAnLxd+AP8EOYx68iIpqjECpCv8qqwuv7BYQ
uuWtFlfUmDUSFckIv71YeKQ9AQjUETlECvXWBNZdXYy3XjRAtllv8zPbChhh
V+28IyICkjY38pITW3eFbnarrUh2mrNyboEAi1zb+hHE0vYN/zAGetymQmlq
N5Pbjg8kcvmLjX/j1ZpVZc9k+S4XR8eAJH7fuwY0aXP+BfTFAWXa/Zdha2hK
nBezZuSb30Lyf9z/R6qePx6GLXyKd0C5cShUWNhNg/WrvSrC0oD4kmPOgL3b
b8ZzAGCL+NSLT136M1FqygFRwKSRmMt7/+ijPv6uyYl7zglfSO8DF3+qfnkw
I1A7B7z8daR/FfT4In2d4n5KFIP6/8wxbEW3KhEydgQ5YIbxw38qBMZKZS0X
iub/6m8g7kbUIGJ7nlp9FmZipvG7Z6Ea/uOgeSiv1mjrJ2CmSUgvKvB5xaUW
WdAzE85mGmMO2bKLFZZSG7FGEEG+6Dso8n9CooRBcV2kRKyYb7wlZ77IYOwx
pDESzQSVll2JAcYWJYH46ZPX1gzpTw0utARAJhMuTh9HHJnism1NY3dLlAw5
3DRSvLuDQIn8kd0ldpo2FQ+gC+KP5I/rqQ3xn35PHODZFXUL3NyP+EW5yzDU
L5QcNnwPgaW0t75o58HdNEMCGo/SDdb3gr6a/2k1QcroE+o4yMaZs7guQvWp
g2/C6O9O7RRp9ApARHyBzHgpEyrW5NjgRGyxndH/616csQ2Wy84blDU2gubO
KoLOOYXjh+lLexvXDdE7B3zV8+entb6cgNWe+D4jr74JqNaenan1io3/S2tl
WtF3whJ4X/Ff5NOz7ZhSO9w/EAvkMbFTPByEmHri46vgOsgWnTc8G7tV/XDm
Lehi6HjGT7Ido9bFj90qy16bV2bRAnpXYdmkTsgtx7OfR5kvs2xVnEg6WxA2
HJu6XRPLQK7+NTosF8tagIkt+tjglg7+K3ZOQMlRslxnyoz6i0TmoULC8V6r
P1kw0q0p2b4UZKsuuQe+8CrCakr5vbwTX0lZrV3jMwMxklMLYvrRwE0nBoVu
ERMtzhlxzcbN1eMls0figJIY5V6bqo8BZJU2/SAsU14hTv3aRIHjV75AdZUB
iZ9HB6jfOpTu3SNkIycI9jau6g73Bv1C/1zTYqfLqXSNck2BvLtOUWRkeNz0
kwbITKHPMOgtSJYbuagxk1Yh5215ZCwH3DtEvbozQPalVH02nThJ5CNr8y6B
CC3Bmoqj60xCSoNm/xdfrzMjOJZHTgK7G54OjQRvxr3ag5bLGYHYoJxeMFb9
7JAfEcNLs1lF9frfe096MpTC9v3EUon6l6c51ePn2mzJN64IltppKK7/Iq1o
3Ywp1DbEi9IIPq7w++v6UyIJ0am+tG9RymdaoDBipMgmeuMcCCitN/brS+mV
iOxVaEUO0y15eVZE5j/fB/IZg15MAM6g9PLik1gg0VtqPlwkicB5UfmixdwY
2skFxsUVYxGDbDPdSyCnthZqWQy703DyfqJD274PRLM5HVIHTttv4BY2+ATf
O4541HmDTHHeZhdAtfwwK6KWEs2cQ3/VBOQvdj5kMNPEJQ8PSco9APas5yFA
7s2HChIJmW6O8c3h0thyDbljzQgNvueF95dqOsNU5XSGKgF0oSKKOz2nxaph
bXhkVOHZmzOCWaeGKaz2z2AK4oRoXgvWc6g2ALWqKL9f0+tpsbt6fKYaC9QG
G/w6Yiy3PX9QbNkot8a0Wa8mPIhNEHFBqWAMQY92OsQ1hgrsRYD5CYqBAzey
PJQfMYesiKyfeZ6OztwOPmVnPOCKEQsBMNynN+ABAk5QN9vT1/2sx2SH6128
5diVLfw+XLiCnyGob9bczQbDlftqwrhGddnCLz0XuP/ppvN9Y1sTXPw4FkMf
4c4n+L2Kh1JwtN79IrVRWmEeLjf1wU/06W0IEb/2gIRyKMhz6KAV0rsC0IMb
d2k6BTBF0u/y+C24fwGU08gl5OOt6RVHTA9D7ceaZgbv8wGphwRsGz09LzQ+
ci8+0lpvcOBWKEWsfj4Sm2/7JR5134730OMEdHOPUAizvZsaUQaSfUEFBxCW
NYKgdEA2Tf8X6AvFyNv3pb7pHlws0iUgN192FGd0Jr8W5IJvNPeDCqMStLDc
xZ6bAvWLYb3mmtGMl+4Q4LORn/O4PJZ7OPY/uqCKwh2OEVbqbTIHxeTtYUYp
OI/xxoT+3CgHcp32JAT8Tx8lBp1eP+rUJqYf/9DTqrpMPNLRFS/iltWFCF86
r/S9rAeFHwHQh1O1iS/LKBKobNgNKGVNYiUpM0ufkTs6lpbcoIuCx8DdFPVE
YCsEtG7y747AkCBpOoJU3B9V86Sk/Z0ZiWxksyVZ7b7kBi1P8iuE4xNORTPE
nVb9oGrwJwSnRlN35ZY4BgShlQ1tg9oTc+HhQ2SP5eBeuT7g2xzqGdz/QN30
sM3K+4OhzZ3ioCHNh0kgceeriJ4tK/QiVvGjDKNaZnTjySNZx4KIxDcbfND+
QRMrH8vURkDEkWwRyN2sR3cKp1i/7ekKKocDY4h5d6PfIxXJZoyveeRY5sV1
D54mDAcasmH24M9YZTfnAvemLRY7J8k69skBhoYiCd02x37m3CuFVR7FtSft
AGCjbchlz/AnHfPm9Avk3Kjlgw37leD1XHFBEE/FQtizwpYTIeb1gIR13gPA
P6aJzR0OgO+sgoL33YMLozMOZx6zMqWBzLPMeD4Z1miGa1edbkxMku8mmNgk
M7TJpG1glxmhLIccpwTU9noZ1ATGMm9FTggToPJ6lsA6R8Evj6wyZ0fyB/fr
34mcdFjI3S1ShFoYAxZuzcEkAjjcZQt1VLcvyYGj2HRVn2/1VO4YxI9CPY00
d98nYzv5Hop4fVtWCkjqm64BOYmDk/S26zqxqvi6XgM9uwGVjNLPH9Oy9Ydl
wtlQmGTlf0sy4B6+y7bTYR6Vr7HgS2Y91RU40GVpWzpTIKn+zoXvEWE/05Wa
J8LQIRcjGdgFtzY6sEaDE52v2UHv5xcGBZGKmYKP7aiaMkRNWc8CjBqG1iOn
bPYXJsYJv2Z8B/SRDrYoDPbYNxDRYQdh3yGzOWX7kN+LANtkix4xCqZo8tC7
BM6boOjK5HO0s/hWqAjkKvk8p7NweoK5XJ69+xGPn4oEI/AP+O1D3vjwBgXa
rH0smqzaiHUI27GYmmqRxe3Jg6/XdQFF9gnVW65em2z4Wd7ZLdnp+x/44TD6
V88tF2do/sLvHhrvmCIvH9tL9KcUSasAwRljqLb52Go+1yUZk5XzqY26//5q
YkEgRlQqaQxpGJj53T13lFWCevJD7rnSfFoO3NamZAprHmyA9hG4aql7EmTP
5+YcMyB3qNI71OQU3i5+cqs2J7J+ZFjoYaqJahibUZJfGhFyzDcL4D2rsysC
hCdLPIQbKpidz6oRoer+2eIFS3vo0X5AVufC9uzHJQ3vWnZpfyAoBiqR/f/J
jy1PGanrKbSnisT6jCd9i58P56zesxC9CLv1pMtm8p96McWemGgzvUqxEfvf
UiMC7gFmYoYnJ3eJ0EjR+NdRaC8kiEfrLISqew9CoRGHzcXf8H9xS9cWdLIa
fsr3PMnwbO1grG8XsD1x94vkwvMiIyjf01RlhltUyBZmWeW5hYeVPl/QzbFR
p/8tc+v6xPKZTEs/vt2BEkWFgP8x2ZJH0+HioB7JRm4Fxb17xsbElQKSAqx1
uaI3WFkVw9r0Xa+VJqq7/KnY40gNKMQx7p3wlLGlh5baV+ji6h5BzZyhRwQl
dR3D45DUqQm9/VrCiPDN5Sy9CBWIgg1M9YAiIGz5Z121l9dkFNLvzSBbmJyv
JC17ijUJOjl+Nhxqhhdwcuip45UX4b+aHWwqqKUvUfQPg8Ysv5+TlAD39xy5
8QHJeW0/zLomVsHCLhL7bJUFkp2z7srDvo8H9zE1XkNC5k9hZ61lKEqS0yNU
qRfAJjoSMrWMUKTl1oixR7wE4iLdZIh1u+hEL+peWz1cXZ75FMcp/oav2x+b
h+bFbITsBhA5b4XhfCxpVcgvd3WGggn3+raXcW7LurmOOc2gnXu/GXonm8QK
vEG50UGPm2ZGb2HmKPQWjiIAuB0zVB/DCJSjrEPpC3R8WRMxIkFD9iQ04AGp
8bcSDfJ71gkDRxL79LGr5j5f85g2K7bxkY/rxqKpLV9u2pqhQMxzfsJIRCig
/uJVkvNXTxTDFrR2mIHTpN2laNIrzUgnirbVZtzioYwJtc6Ye7OkDoA4ZJAK
ZYs5Dnz95Xi4R2q0/s1x3rspZE2pnKBGGnc9/CoSa0WYT041AZti/uXxwN1y
2Kt8kwvhzJLI9rv88o5rWWqB7Ifb2XmzadQELPz617Xd4f3zLvzIl5lh40DZ
lmBhJwTau4hPlVt2yX5+OB1t/QS4gwu/V4esKGLHHVgPNJlFQj4htjRsmdvk
nUtafq/N0qxrxnDAHOebj90vhjndwhUBnRy+Nelh/6N5O8UjBt4AgV6HKqd/
R1U2sUZ/QltImtB5RPiQgINd5BMzH74ZAFP0AFQpttg67pIb8p+0hbRCr+ll
sV88cM+HnQFzU1UHmqPNFR2MKm50qniAkq7+687hgCARAfsWhDDbHshMc7jx
GRrrFwDTSzW8eR3B7SGN25TL/zVDwCTn8hnlSqVpiN2wckrQVc7v1beQ660L
mwFNl2VWO+bmtSv6y9o1YqAkaJtjoqRV6OWWCt1N2tdpilbsF7SnFknZ0Eyp
s21xk2zy/mDp++PV0jbm9PrzCzcrS4hJB8xrFIziY0wONkU8XQn6aASKqHmi
eXIceFt11f+zp1R9GH9eesbA9GwlKX3P1ayi38QWsncq+Acsdi6893H+RvKY
JlYzFSzJuNWPQWTaLace7Z9liSrTQA0HSw+chvP+q5Ms0GZg+8hQXCmRogTa
BRUYRO1zKf6XBzJbv9nIZRG65jQHSU+FZ8gi4Wl1hcbqnkBquJw/WIvNsfAo
E3ezxROFV7kGGJMow9rUq/ZV03cvaJXaX5zUOTELhYeLY56QSakBZq95f8sc
lqt/su8kLvWmztrp4Cxfpbusc+iNo4rp/ckNhKI91ipqZFMdEDNOblRW9385
wVPBKEyvSIZi5C7oEX2enlO5PqqNwgFWlkQXhgW4Rm/XJAbezCOeCaqQWD/m
6h71KaAZnCRnyc2gA2wzgmsI1IZjsyadcO8DxG3Uc/TpZMv3lFdEybK9R7dC
4Bf8H7ooW/2yTUcyD1lm24TPDmQ0raV0MJvlXCMTH9QbsuAKa6G0MV1IRRKS
PejFgBdD5ft74Z+/our08qdr6oNP9S5eIk5pZzGT9BH6v9Whpp0pDXo1No6L
7G0DYuAJptJmlO2Cr6kvF/f7P1iOXqkeL7NtVZLJXne3wsxtbRJVCqcPFq10
THYn3ezteD06lJSGlDOJJ+1ooFroYntWQf2f2ms/wEMvUQyydqFu9G5a19y2
fpqFuEhBUocMlD3v8BmHP6a6tj6mgOyAhyUsYz9JhU32MEN441HeoeuM17lv
5T/VldggudtPbD1JiDOa3KbQVkCh4w5yEPctI1udUY7wx0xo9d+/8A95E8T1
Fi/sFIeOC4P9P//OKM7aQVFjHVDn0Zff8oXK5z2xck1+OZbHu71WAwXLE00n
S4xztr6kCM7g6X6TFnCUE7trAf9GEiWFM0qPzyUtfBvhjXgkh7EaAvfVZ1eU
lCEHlr/Jfdb3ibpWpfnn+jjLKk3wT4jmgyuzAnjM8tw3pbGFsr9x57sCdG68
HBF0G4522sZtVZixiPl0CHYpf4ET8GnSnjHEBhQcPs+mtXlBCTnDRbdziUY8
Tyj3K4Z4MYHZqrGzuBL5iyR2JBj0C2N3vndNgzva1x5EqMaPJhb0l1YX2j8G
vJjNyMSI5vWy+JuVDEmQhjyeYEzce8Ek/AMLia5FunbxsrtlBPmF7KdgZxXF
3VzxovoWxbKgAUvvYWtM4WeBXBZoFNTwItJSZnOz879QMZZZGrcTwTNMei87
glIWRGjV0SHEPoEq69zl2D+8N6v1VgVfcl7eFD2DbXaVt88OEF6ZNxoox9mQ
Urj9AISrDmdg7OI39I541LcpyUnBv8+6VGaHesYT6ew9XkxF2ADiRpb69XjM
1ExsG4ueR2NnAbDyWNxHo9PdqghOYR0XZt8CA+STvCmmOuwKjTQCztEwcBD8
VT+wHKNHoBF1VW68I4YmHqMApwW5dgrDWiPCB1g/MloW3LIpNF4J3bMlgck0
vbJPssMjAJ9DKXuyfnjrP/d7lFf6H+7cHrui5MBBtIyCvmgnQWm9MuXI96ie
L6f3q3LWq2uM3JRE41Fu/xOmVGzIBRuaaZ6YxjYXcjw0vAPwfPKgRiwCjUOY
iEi2yJj/sV2jnihA+OHgkWchTs407SmJnqrhddjhwYsytvrsOCUWit0IDtsj
HJvwamBxQAY+Aq7+gzwu/TYl8yG9L/hN1vpNtTUVMS4squ7W/7ZghmkxN6kX
A4ez+e7g7g43rYjoHUqtsErXXQghY2Udt7x2y+xLq6SroErkko/PmTl6i/uY
2JWVtXoa5hq8tSZbYWahX1VYhAsLYjdf/QryPogQ9GNbbPEczwbm/S4t+aDo
bANqhCMQlj0jP8fl+xNnnynsWk35n6IOxAO/Qfnz5WZ3iT5pZdmvAq023TLa
HhBwEwPvGlcLJ/464NT472kCGc5rln2d7BpH9/33e8HMZhQTP8TH2Gb+135X
ntL1opTg7PkMSqCZ/NOMhdN23BqhqLXLuquiYRpqJ5dc+Bi+cqwYYsJGagqs
5i9zPKubKHNeS9f7flxpQXxT0/9ySzp5foFnRuELK9+zV6q6b9ZtzB7+E1xF
sI6p9siOJyCKmN1DuMSsrRgemNBFpPtZ1OxuN26hJdIKXclKs7vmyOSMvbkR
U7mOEMf561ocBGXipgXglC1U+cRQ9Zjqmw5HdO8FgUsystB0FFcyUErPURUC
yEIwyS6FHZALN1uecHdRmyHfYLM4oQSdxd+lxCJXNEY1D9jRttgkPl+fKdJF
lD8Cp9ZpK5wG8EV2yS4T2i0WEFAbV4+o7lOFiiGIB2q17Eti5nhb1lQ5hrVY
YVL58+wb7Ux1Y79qfxA2HCg+MWxuekuE1akjcZRt+VrKbVEZEbuGQaZ/J5Dr
IzN+ZzM0YHzrqLZ5g9OVwIPdKAvFJ1VKARgBrEHVkyKZobjx0LktZhO5WRa9
2jE+TzWwg1gjP7n7nzEP0Z6odKsIxHD+GzTT89BeiLQSMwAFlQCx1O1wzw4L
oURkzsqtBxyBAWMjAEkRP/eyk1bcRweSPMKrogTlXn3/uGMAdTitCQc2VP7I
y+JTgDVTTQNiQJK0l/Ir96WVQBkI7ZI3NlDt+dFnmsYTQEA/gEGg2kGGu9Jf
hq3OedSQwzJzz2qCFZVspJOPQCqE2JoRehD1jqJ+VIcbxyTSGB+0ORFxhE4S
UK31Boshlfn2jdnZjbbqCurVVMA4jO3bm0xmZCfPofRzLlAj7H4/A9+fFNNB
CYccTI9D1ERgWT15MC/LyZPFw0tBIFkhyPf3eh+kbPta5n2dJsSnYKCyOO8l
JY+zxO3DVGoWjqoG4kZDsbulnWJIJA7aZjg/V1J5N/XO3l2+MwGpAr4EtV3C
cMjr1BCZw0QTX8/i6bog3VnI6/0+cMYhcVbS2P4MLWPgadU5fR/c0MUnSNug
oFkQsBcMZzbqXZg0lgvuc4+QK06+iP6xP8MFzxtZRguxcZAjGWZuCBqnfgcA
zVyz4V5eZFly5pJLi9y+q1w8VS52u6QbTYJb5gns2sbnXCcKEM7aM7xzZ4dG
H5xcRuo1iPXpL34cIAUqLZv5diXL2TxZoUEbLLVri6kpQMNGq7mw8O+DudLz
SLnnXBE00MmSupYjU/yIJdd+g0+Tj8VmKkOGwhTweOCcE8wRQota/dgUW50J
mUdxuMRksjUqEec7H1Tsu1o7FtrokkIAVCIA3A+ZKMqrxMmDG4I19R6gCFLn
d3Ml0y+ZVJ6l58EJ6txY5QewjRtf7D68hSoiGtxPvGKQOZRrUcRYDLEc74yR
Mf/qCVJmAKeh48yojQOPRVamUXy7vqMkqWsGFEGSWMJHWM7U66OGaWWmYRoF
wkJl9GMPqQfTldV4kOc2HxmsIYhuL9eVTMn3jVkO20Vq1tNqBTf+xcc2/2OV
6GOfe+Dhgy9O37rqZGn/634rdKH1cxssyH4tRyxciCUf64BKuI0in7lD7Guh
Y0bRXDrJiCVAfXWaqMAOlcYZniqrGTD1W7aMB6LiC2ZOzQp3eLP3mjhECPOF
WkxjSTNQMPcTVLft0vSLB4JizaXyNlAPDWOLtEspdSno0c4650uG5PVePbWG
+lTA6e5ukT6YsFLzVp+ZWx5OBg/cKHZtP1uxpJ4VkH2iYU0QSD2vIKaHBg5n
cNlesdigBf1l32509ilj8/9MZ7d25HqkNbxtRmCyTRpAT5YxvGyVBluTPE9Z
KAFpd9TKMsf0qnfoM1bGFb6siyxyKztVKAmDQgWDvvjxygcflw9cO9c/DtKi
amPzmRhU1oJGsEHJ+jdloUvZDVSR0q9Bg8bI80Wue6q+3pXFaFpdWpe00QOb
8eQsS3tHLuf7QFV7gW2zWqRnbOaI2EKgbWOoWYfQyrGQ4j+v4tCBOO9eAMH4
Adv53iitp3XVpI2PBkjEc3jFAlCAr5o6i3a/DW6jbJGI4KBnEmoaSMfla9jO
TX5AZLK0KV23qLbUDpUC3WE96kpGnDyWUaDM/5XPvWBPKKGiv9E77tJAYbP9
iMCIOf8VjhQGOfKJjPyWNMJ9+Tsxhg5jORA4extlc9P/9ZwONjcrIPVJSVBp
EXbuO7kM0R4ILk36GBrNf9Wf0YpZP3t8OaFnD50tRJbSuof7GwKcRk3sqb13
1KPZ0Sp3d+bfbFyczRO2CcfZTELYH7fSA0KVqXsEbBlwywOAANK46bfSZOUD
Ow/WF4YUa3Fget9gxLwSdSoJr/P7gtNVpNrV5e+VSyWsQKkw0ietHlye217c
kqwYe9eV/zyiYVxsMHXjQdFRflAucHgdErT+5Y2OW3KHmBeId+Qi/QLXQfj8
1F8Z/Sd/qO/jlHTQVpVq4zr7fIv+E8L8jGh5z01fgb02QS6P16aX/YjyN1aT
Fu+u+EPB709fTnM7qM/Glsf+m8EXS/GF210AMpIP9ZSJE6gN8wlmjiDo/+RY
DVvw2+K0K1dPDaqpGxskpJWFw6gNq1IYqylajhGjC7PrQDL9C7kQd4UOKEE9
w55/E88RQpvMBp0Jkt8TB02IceRwnNK+na0Wxl09vKsbk2NgfviB+OJ8vrDE
Ryy2wvU6bJrckRskaxLoJpC/0Rt3iSAFaMX5nz/nh4xISMFmj09rjgfN+Hh3
2u4B2XO9s9IDwsl2QtaL3gATzcp65++GhiahktD+85tDZwtkaC46wjbxGvcC
7+Qs1GOo/c/GQiZwsA7hzAw1grQTisgW7MKr/Fvk3J/7YAgNSomIFTDmHwK/
HztCYsryaR8GA1IxvMRBIyMnwHUofr7goUppKzaht2uEx3ryc3fUitRIXWXv
PybKUTx6rcJwBx7PBOSgWcn66A5z1twMRGj1+3p4JYo9BmGCsJYWkcvWoR1E
s3gbgh98T4XAFStRaFKUT0QxGUlRNcUPCee69air7TItNHStnCjiZx5ZIdHW
dR9dQtFkiQKR/8yzDCTmmrisxIIkFQ4pKjajVc62KzCquB1XS6eZtckOmzDP
r4qRzS8Z6W2pLBFjNRpb9W7+KlckpSSBWetz9Q+R+tEpYhVn3TB37ZbgxGaK
kfNyEDmQsDKtcscHYBOlVEv3GL6bBEOyH0Izs77bSHEN7zz1cxACJ3/MDOKL
zyHyZR2M9bVkEI4Ya4Ugt5nIWaTpoN0hteVBWzy9yAprGzW/I7pAIesISuds
7AJdYc61+rhgyMSpU7A5kHeiYcSAoif+ZRx1ZTITn90SYXh7MUoEeD2FtMSj
n8Y8igMuCckUFReAP4gsdXxsOnF5ytBWkmgMc8HGrM/MP7BPv4wQ2m5XVgVY
qZtYNXZbbtSBKUrYq1K93KYmLrUCZHFhEcny4mMLgIeA0uGLOkXbQ8CylQlA
T50176E4Hm/HzNqRGiLCbCjCA3JXrkbjHipJ0hGHTHTsmg2Vv7IacCYLp3fK
Fi8+Obc6IlITKPKq67MEIKKQLM6HU8V42LDHEMUGQCoQxiXemCma/YmMJ6PM
Qpja/QRtmLQRkUGNAIeJAYABLXHj4gTa9MP/bIA0mkpwisYt5ErBnEhTMqn5
po2otTl7OSaZwY/KvwbIAUsSZLr30MxpShtN00igqMuWTJ7sl/WPjYByDfj8
lRATzO+FE9BfA1ijh5/wscuiZwmwXVkjkST70zq8ES8fhnVmQKHwMgM73uBP
6MoWfWWibjVQ3024gdrQuJAejZKQP5heqMIBLXDjKGcSoihGbDen+JLEwMmg
5TVgmoYZt4UfSYOlxLSZUYviJQsldxicGzH8HVCCFn9NDvNWjvlvEse1Ggy1
5reSHMO7KD8Ec3yQue8uVYA7yyWRVmL6T4Rp0Iym3JlFY87i/rE2kcQepOL3
exX/gxN251Ky36yrWPRXA47hhKdpiUO+7QPgNFfLlNUyiUzrTUYXfKHlfD5d
GTNQaspUebc2zWXoBduZfwSM81WG+THL3GJb8r6hMhHFYM7UPSgUq2jFRFRF
vAJWcbnNIo//hWgiVxuXDbdg0qy1aW/C37NEt6T527RYetpGwyxgwu35BioP
OfMNCPofDu3UWJui7q9geZ2d5KbD4Hcep/I9/W7orsZovEB+2iNaddMF17e3
7QDDWO6BjzJEU4RRnUO17DLD/nHE5mNbK8IaopOpYA1dNsWx/6zamWc5UMu4
GXKsqP7tJ4FRWiU+sk3IYGRAfs1XxLGetUt7D9Jbi6/vLhkt0BulVZqItSrK
dizWXcygcO0Rnq1ilxCQI3wmtZhO6GdyjXzkiGElWxAukyiCoJd2PKPGJtD8
7sbHQ4cwQmzp7RjuABZePGTV7Lbzh8/Yk0P0AUnjvbD4+PyX0u6T2SwuGgs9
xBzSpi4pBUBai3ezo0YTRyGwV2ozWqWrsDIs/W6WVVF+OBAJBUimhlNhfn3/
pbegtqyI+9DfgMyw6S7nT7iE9NnE8ciXRVv9mvbAvF4wWdOaI0PvDXOFmtk7
uRT/aPCIZA9VkPyerykHsOztQyp03TGZ3D87X5zHo0p/Xrnr+z71WjJIVBht
CxIPFaxh9YDAbaXtqaOc7UWfSOO8f0Ew4NlUW6xN95tsyGAJ1+pdRjfeqrf1
Zp41qaC4xJLKl8TBdll3ed4fR3A4Cjz4TKRKtDn9eyd59TIFX/sEH0xkvxm3
5VULOc6mzoC4BCSNFYNxtOk7mIMl+OqjJrSkX4D/6wWi6gPDy3LM0PdJBpGF
iPtSM+GkoFcmm/CJJQik0mcejhnOQAPBu156VNJruUmaaW/4z5ECt6Vxwzh6
3XZ4q0f27y7969AQmJEnL3Noz+ZkP7XQqZ2QoSAHpzrKnqnwUlmctFcPvi55
2rEPLp5JlLsxsl5aK/dGKpSFsUIOJdOkRtk2eFkIH0XYKJWnqBX8ciU6TenA
O+0VkskZ463k/itORLjZ0OovBQLZgP6XP0f59XKsqaVvMNj3JzhSCG9Kf4hX
2qO42J42V53mgizJFF9TH5dU1fysUWYuFHIu+pbsnQg+twjwq/MdxxAMUUD6
zqgN/Gin1PwsSCK0SNxIQzrbZPS8WqhpSa9mJCzALhGXn6UJzJrEiJYejy/Q
8aRWXBIOJWADi22mks1UEtF2ET3XegKrWzN8N/85QKrAkiWweXhCrZyTXObP
1+lhCk/PzOmwoHt0slw6VItHeAxN0BDufYr0/tcdw1rTRTAuCtkYHD6bSeFX
nNE6NXYnFTTP26vGEjJtX4btDttRZH7Glr5DIdFJs6BBh5Cv1eVyMLjyj6+W
JyOJngsD+RfxLhvLq1xj0a4eIhfqqCaTNsRevDB2LT0Re6ZBmFFFYn6nSJSM
2gYi31xkGHJgTquYHJ2IAOkhQB0Umc+6cBOdix4AFHa+IVmYgub4AHXmk7C0
vpTADWeVFKmxtATQkujMFaBLOAT2+NlYpQooWI97qZFNCQtgkLT+SeQSOlDL
RGtnfRSqX7WjR3LLPER03SPiSk2Z22X4h/CAPjMahiGIxpaj8CPczX3PcGoK
/ZK5KlE1477/PexEQ6nCFAiynupkdSRp0mjDryHx4Gfs4P06CVQB3+XZU1Py
cXBFDM9qB0aSAax/jyJs4UD7mX7F+qOI0CHTWely6jHhFUIg1JTBCVRUFAS0
z1LATYUZCFCTm4YTE9aDxMSOQY35HLmPbIyGsm6YN+KKNbavPM6+3e+nWQSC
ZnYVP3cnxFJvqA+H4qloJeb3ftjfc4+sp65I/0rcrkEziJRt/8ouQKgp66nq
cKWrVctFLIawOzUTE2mdQv5Cl8m40zOtKS+VpEWJ0tKlWtdD0rFmW8IypD9k
C2coaad8XU7iN5Z+kvM5Rl8f+38ICS0IYxTJ2gOY5LFrv5MSeC0zJWg7IuBM
5uNMmUCO3FTjdeIVKUVGZBCwELEqR25sITwu6tYCiX2FwWQpsLlXPyYHI7Xw
JvolHW00SiGPs0j7CFBNKV/pbRpGH5SDl9JYVgmNAxW3DA0gNkmqmYTSIaUV
1U5DtIi9kDzPT+skdf9mXcd8ZuBPdkiaLbDBSQbr8Mada2DiQoI9F1pSzsqC
OYk7rk36oyJbmqzSJjumvYWPXNsIEUtjyPM6PAJfJGinS32GuJnBjDi+FTY4
FTWyX0leX4VoSUi88WEffvLSXUHoY64ZYT6F+Mq1R+0suXFLu+Nyq3yozt0V
xW+1mvn+9v3MDft3Ac0Tasv21TGjJokVinvAmm3pDix0G79yoAnUfHyuJBRT
qziULHHdC6LX5Dt+sSfMA0Zut1fKr6u5IYBTJ0OgIgnHJ5Phgatomef7HYFA
lL9UOBZiRzcAd19xDFSDVZegZuW2cqIh7f3FtkOS/NRNFflBQY+81fKWEWqq
AZ6rVzKFLRAKvmRw834GUIl/3iLAGqImuLKR5bd+ihR5Ceg1AOa3MLWc1RuP
xJSifjKVIRccNwA2frQbg1y2dSx2WomRcv/C8t5aAkrUpmsrkdJa8cu6VoSL
2DC/DgJuP3yukS+Obk+lzGGY1iJXudPK2oRB94ADWGhtvIEleYp3Aom5Oqjg
3KIq6kuqOdG0pqyTXgn3h8lNO/eKluaa2tFtXjMYeeDrXtwKLQGzgcwB7ECi
y0xfWK5zc5hhLg3Ec50qiznypeLQ2ClMkn6Lg5qzFhbsg/Pem14ePtmgj1xo
H2eZ88YsVFnDzMKSAz5XNQL7rV/7GJ+ZO1aAa26cKAfXhYmmgVTl8s5JPFes
MREr1IEmyCOjWSrpOQ6UyDEws3RrLN1NtnGmPmZVX2HIaAX7RDFNTydl/S/K
TRijeZ6j9QBHpISv/CHFy10EIa9Y/h6lIVrH9v969Htzc+1l7qOtoag1N0N/
0/0JCvn2ttNFJj19PymMVVLYzYCiBFGMwuk8JwyOqYbffQWRCAB/nnSGXIWz
7/t8wb6yf2G4Vv69VX74+XpYGuWqHM1iei0w+sWtCcb+IEZEjawUQMs+xxDP
ANC+SzoVvLuI1bart0XoGRZbWVP/2gK7WXFSAJJ/HzFtI+pdzXQp0smiDE2h
fbcgRBChOy2wkCVrsluniAY7Q8XEGAWIlqYFuhuuleJc1snP4iSzFhHQCqXU
PGBpdRGfvekSJjUdrYNSA8cL5szwuwuN7sisAK87qSQUAS2EF5yXPACbJzCa
4fGJAeVHamj/SHvUiLTchg0On2BhlI3bH0aTHhedZAFIMdq1OXFvYNEZXJ56
rh+c1FUoOD4oJDkU1SIl1DO4xw7Yve6O5MYvEhASpLzQP/N7cwSsb4In94HY
jhXroTqcoxO+AADVOJGgnvh16ppKppw95bzlIM7h8fVXT+76LtV41EaLuNRA
GSu/5HgN4HbCH8+PuVlrnNwe6o1d5426hMD8dUmZgz3zwIGLltGBZIf6li0s
Oe8EMzShzEe3GiZv4/s7LDMFnlui2L1clBCrdaljh20Ds0FfFxc/iOrjwvW2
ddNMEoENul0LqGWqpLVjolV9L/Yrum3zzt178hvzBUbmxiFGUXCJNMnSMkp3
YNT9uGMqpPlU8hOowKt95D5J8ay0xIER414mVSNIQG202TT6IVhz2gsv97F6
LXUnkOa5pjn/JdT3qQjiEJ2cPMJb3kyGyGg6cTeDsCx/tFA2+G9e9A0jp9xB
rQC6qocnQIpy8hxYKvolCsFLcwNB1ZqFwhqj0bLKmpGJWkmZsY/plGwMqjUu
N54zDI7ZhE4lQrl82RT2wxg9bgGAo+Cn082il6WuvXCanOOEha8WRa1NabEv
DeITtone6BEiQqIFKK1m1vMOWdZQkLOBCSDWtUtpbjRUO+2u6aZesBM7HPYk
AUgQ6Km3SYYYZjY/LwHKK8NfZFfiMpG88xopcBXamhBi2ANFwQT/c5UUhejM
iIoe+vtKj7Dp3SH5Sw70PJhDytV70KwvqtqAh1AGRbeoNaO4KajNdRkpcrkd
L4t9ZKCCR+V36RS8QDRMXhTzixfyxr10j9d7/GbzFWQh5CV9RfBgeqtltaDO
QP8aQ8DpeQttQkU41VYFO/CCpQwDsGe1hJQUwmKIEXOI7BJ1DcSZuBnSjw/q
ePISEy0Yakj/BKRWZFIDvf9C75CHBSJeHSND8QrMQLOhlqn6jdOmI4vnk/XZ
54ETMFAAWodGEeM8VEIXpPt77GOwUNrawlIRj62kf5nWKoZJRMbSDvxjHvvS
TWL2JByb3d0h0guZ8ZFCzAxeCi/el+U0DyfyXWvKWuOGOc3i9gWwSRN3Z2dO
SddfsDTQ46HBnp9kx54KiwIoaNbX8ohdWuRI/6QvLtjr1jv/GV4UmEp/dK79
uW4eHLGPdSnn0mnf27wF4eHS+6UtS5L5TSs26whfdBl9szq2uF4iRo29cAED
9UEuoq58WOqGDErFu8hOlIwGgnxx/rq5YFJPqiuUoq59hjGQckGlipo7e3Yz
aALAg+BTw2od9vVhT0R84OtF4EQ0vBd1ifoaEMs1FkGAphV5mAs0h2biwgKy
QUd5aVSsyQIRHdS6lHx2WRdPe83qBS9j6RY3MgYgO5rHYOk/v75ZEfpmoIsu
oDRDpRECIt5DJPv2Tc59sMzvC4U2upE2N3KpjsQxi6PvruByHNTXRufT3m33
ne6YXCVz1m7FJfsDy7MAFGguROPaPkVMsOTGBvoa92rts9tVeEehh903ojTp
CCLdB39113ah+RgSDicuuRA8qAO8ZWPksDTb4zUjb9u8MuN8dKJKxSwe5NHu
mGTHG9W6KYvjvcIexusM9w4jup8HtaQSJgvbxUoJksw95UGsahMUTYDOUOMS
+MZDjGSJxbgFazQs6kC/VpHoOLFWqpd9ODtDMSZGzNOI4rb5fGV8aOnBfyce
xYS15AYjwTGxSAi1Ik2ZDH5fRvROCn+uxn8A7F/r5iDVQSN1MdyczgF8+Rb8
uwwV7TxTb/kH6fbZerlIxCkD/6rG5zAVqdsuP+0HK0bqqWMADGyOD3anL1jt
U1gxdVTzjZ7Z4BsEmAU4LatXqw2Dg2IOlpOUaq6vy6ZkTdT+D69UGSAqMfMA
A+HrhLnyKOr/4s4/KNbH6ZAv/J6EtMYr3PZovOJtrfLr5OHVhnff4qdhZLuC
floWEGYzEWo8AZWnobPpYPmNXNQJqxDvWcvlYC8RSDlSVupIYpRoAorLc2sG
D5YRI6zrBWet2fHmTMJJR5MeC4H7rzeRDpIIMCO46PEHDKXOkCcsc/c4LaF9
2C25S5QedlfWR129d5cm9QP4Pj3ib3+TFf1pjsTDHtJLYKQWqR6qcozgInZm
xwqdLBNVpldYCeAt8N0tSvi6X9O4RFcs0yCMOd94WJn5VVJl8tnvVpZFx/o2
LPeFzM2TC2iCFUsCosYl+i1R6bN4yKHCuUbLl7KoZBIkA+nE1TZfUlgOeNVo
VCImNwn3K7RY6oVOisELq7lYJy+bT5rBznY5DbiXb6QC8GUgxSeER56x5Iqo
ZHLQO7kZ6umtpkVoZ1k9OIn1ItYcqEVpOOoWfDQymmFyqvHGHljH4xe+3Cit
MpuS47p/ZLCA7jzQ/CnOdi1dc2xI+SwsqDsbBC+TV6qypPD+faq6ilsqKwT8
gRCm5yoNB731PX2+Ao66mJ2iBoxNs85PWDUR4Ue4A3j08pDr51XBLu4l87Cr
AKkFjHx3IU/IwcO0qQe25JQ7aSFdQZRBCm5XVh765ryjFc44iGq9RxQgVSvB
tm9aCryV7nsS4Q0OMEKxMqiOBBlIL3TOjI/5an1V0X9B1oG1oaqBc5CnMdqi
crtJjfOoKARkzjJHduwX9srhy/yiZb06crLyZQmY0a5Sxijew0LizDErN0r+
iWwDzV0eSrMznaFAPHL5Oc3r8CorXaa6tRISXcacCyXzmubOuZ0kzLQaat5p
2qYsVKvb0R/Ye/i2KJvqIynl5RwKX5vItK+JwzyG1ETo8ZnP51nSbwzrS/tN
slkd/7Th3g3LFeJ9EwpVbkLMxFbQFY9ck/Ki3v/4Ald71Re69cOZ3VIs7cLS
GsPU4sccarnMEh+/B1iaAjy743SEWLhWK24WHSSnBMAeQ04eFdl0LbAQjkez
JMbS9duPja+ekjybCcS76fA2rWRSzOJjCTiGTdxMfJAPbyiBwQuaHbg1UF+k
GAhC4LWwWLkgObIVirdJaTd2vKu2EvP/qnPlNFwUzanczD1s+Mo7ktEI5WvX
SIMxmDjdvCmeOPhZWHEPUYqASnkPEBjGwKwRv8zf+q6N1qzi0TWIOmrdbCQ/
w1vL3vVhCpHN4Dl5kdAbl0B3C+LeQFlUsB1xuaaiRQYMy1tiNGjHUIgVnclS
rQbcf/EibD7zKSObPYrD5AQbm1TuplD/UW77yBdKe2zlO4ZG0zrRKxr/9zeA
GsFpcvVQWnvncUEoomQOghvmwiQ6Gqy+TNxcaKiVUddut+DfOm6cwAJNXvbO
stivshT6/025XK23LfeUm5buOuhgoYPyjgQvZLmUCtlxPVz1Et0p0rQjKqH4
2hAyIqu3Cf5Ea9mg7ZWDJsWpoodCtqdWXOsjsgUicIR/n9GXXEalUBfRoAj3
BRS86yeaAYqxzxHSykcjPXgDPvRcnY9cgsE9kbfcrO8oKx//gGJKuo0k0f/v
MBwIgdFEcmKYIVxf3MS6sBc4kGEtqLQPFAFlO3br1nBk++PpxWKfCT1QhNfO
LtoFvh8qUpocDxOsMw8lZiF9XcOcLthHd93XlkZU+l7b6ZA+nhVpuIH5S+sq
uVIZQBgkU+xIaFV5v5s3XeWVl1UnmrvDVlX2r1dxhOydtsehji0HUFkrvL0I
CuTVNVxaFO+/gsaLDobhuCWugciOcAZ9WmrLYu3QntRJiLdo1ohbFBnnW8I+
L3vmrnjPY373bt3s7hNaqrFsd00sfFbQayosQDN1RVB3o0fH7NQbNvYcIuxg
Xf4Cqo9wRppyOygsA+ajV4xI/98FPIwKMoP01X4sXrY7HyW1jmvA5UvPwkiO
xfHOIfBqr9cDamZU2hG0rpSw/pTCL2auGMT8ugc+QWmrOoQ5pEWBxOmTwL6R
RH+HqlCT//D/MXbx3dZQiQvcWLjGEfybMZ/JqzKVxNLbhoheorC7wA91iEXE
Hi/bflLIxt6W7kgK/gfIRHdNgY63iuPE8RAd6YyjwLy4bPdTmuj1J96QutsX
U/qCc9CM2/Wot4hBDpIgxyC1bRAk7EHxvEtR3rcFp+QKAYRac20t2zOz5qN3
8otfLAOXfPyMJvE6VfPaExoC8RqSoFhheY2F9KlUPjZnK73PkTGbqEDb3P+a
M72u1HWIqdv9SnRwifznO8QIF3E//8VPiM33sQhxy2JzYAHvhUxEM90csUhy
PLwbMTACeKrPft/ANBtsb3cenogjgxsM+hgDZZqqx+YwQBRZj7rBKZtJp9cF
pBpAj7riIR1EG7ueTbaLGzbqJNypPe3vhxtTZcivZeHYYT2Ss8XHX5/tpK8A
9YZ6AFD1OXGbq3AQyICLzvHXqf1LORDzEOTHeVUF+2mRt52KCVDsBwBUlhRC
lpfH6aZ9W/yJsirvqaRhmDmXrIDWhxZGAIVYpmHGOiCrVLOqPiRfWkXH+oqy
0fsrTkiui6YY1K5OLMhhDX1W0iw4CJGnJzXAp/4OFzJgdbtJ8avtohDbSk3P
/KzD/GitgwSeZHGLNPhR0d1I1iRz+vs2bGxGuiJkMEzTEmADav3K4EH97gi9
E3raLe/0ecCQTRL43lVKkGakND4eikaIQybV4tHLku8VUphB4k5zyhqA79Oi
UYW2Gdd3zo2lOmjYZ9FbFmywZPSOJZ0E8yqstBKtj7bc4LYQXi8JtSax+7i6
dq3Skn4lmSJol8Y+/Yb3rGSajaijtkJVXOhd7NxsGhaCDP+igQuA8GqqE4LB
P2XZgfYcyxEDffjfbMOKCHpLp47PmpacXbv/AKEFgg+JOZ6jvGrLbYhW76Xm
mkKKxsAqLas0HToYIeEXt2A5bWYNJwM9pQ3am0IzKvWI6twal5tcsMmrtyat
KdYZGPI9TLEmNMNfh8fx6wJ2DXZxahdvXHIFpmnEtnIo4VDUOma873axlsBE
hiWnGBUw0LD3naJNc2n8md8FaFaYCJqOOijeiB9Z+mZbiZyXxqKtrzzU/Ub7
m2rGRE/rYvkoyS1txe3RQiCz7nViFi9+B0AtnaglJM0Ri5t6sFozR8qwmoNK
BCMYWxcCzWJybkteJCu/fUWyjgaaFVN+ufGlMNXYqQbkAd5E16A0Gs2oU0re
kUJ4AMk7WsJohqMWj+MH+89P2EGUySWdX6LRRyTGT1kU7ElcJ2GwAYVMlHot
2sb6WKy/31KCWkCYtrTlVjE9eIGj7sQLsCPQ2+XEposa4/XFUXSlVBwVeRCY
lAUc7j68alxmeadiXRmpFLBDfB8tC02qMuB5aIiwEZxLZdb2dIseMlORQmpW
Oe1pJWogPmCJP7Pf6UQBnQCEBfQ+n39Uj/EbELo9Kv/RAPHQrrPLvOXa14Iz
Y55psIHwJjC1fBGC1KGVabGDpNSXY+ABg5TAjwSC5HQ70R+GY9U0sbgTCDVZ
I3rc52ohg+khyZb35nYpTqSxtzphrofxvcXKYWbk/lyvCIuNVbbvIFYdK+sA
Po/AE3cxwVJfiRSt3xThv8WZBhJ0rkPRaJlIBz7g5PaDUB9GTTAX8auMG2aB
90RBznLp6R9NTwMVnWnnjru29zKPVTTbeuHf3m7JlgcBSYS2PqQB6XWN2tni
sTyPi8Socg50eSVHSexh6fLuGb+YQ1qlj7fgiauzPlj97+FdgnBa3VxbaNEM
rHhfBYKF0pCNnP8CqziWmMQHxCdDltGiD3/5k1pyBGpa2Sxiw14bjUiNUZXd
JFGZDCefnwBHQuPwpi9INd8U0TWeFNb8n12/hjTpvUvb2GnXU4Dq1gEthX3o
BD64Q1vLF5mGRoH6maIleOsRvyMrt0oDthKalyyoQcZDpAD8fmyToi/j4buV
bN75vihxChlJmCZ8M5x6570jN5OoyiGhV0UfSxtgEmIfr65dcTOM0znIkyw1
NJbZm1Cyj3WJg+D/ptktiqNRlZpUy72AGtrLFfhqEw4f5g01QDdEsy3vrNdS
eQPvMW5IVW9s12cPeDnfkLxWnHHnbjvXaNG17JkbRBWoOG6mi2iQHgA+8yOd
qZwHKjiIsZGYiuwzYmr8Qa82tNL9L0l7Tw7iUB2jI1chpU6dHj6vCIJ7RApP
qgsJNpSM2wabOulj+96VmLEV8MWhJPMC63EG1Reu3yFefHVa5bQNGsqltIyv
vmcQ0JSb5RSPhsnQzLfI9/3l4MullclMbslRQLER86EGvFrfdzcqD434BqRN
uVw82uC+tmVqKQzxL99awiD4Lgvb869Y6dMQRurR3lQsf3PngBWP/aM/WsUT
8p6yOLCPTUOUhusJRwGqfdAB+W080oputGkR9Ilbw571pnQd47YOKuJ28l3i
WeJH7KccRH7CNaO69hS312+J19DNfIs2Dlg2EOpVlSXn+a7PXaELHPap56A8
FMyYB8SHt5U5Ctr0Y6iw3amhfUz4joa5aKOJ5UM9hCG57p5heTVm3Z+AyMyI
xl7d8OW8K6t91uTKmcmEZfWHtbm3UoEn8LVYABXpVTUUlOi6C7pf8OYylqTZ
8wszR8B8DJ/cXUkLZXDARkVqQB18oG57Bcek+o6o8EYldnzBNajxxGobQOuM
e8vja8p0wyCQ6mUWwZ2+5J9b85SmrznIsWe/d7VxojvMLLV80hdSHgs1kD/X
6H5VQqtscCx8tcme107wVT9PJ6qCwf7q/fgoXcb0UP8neU3LELA1PkkV5yg5
BiQQnn7b4Izk4OjqWKSmoxNBl5CVwMczFvzF+bQQM218n1arBtTAGAD0RYlF
DlbyXg1uS9AbPlz4I71gnjKO1F+clrlTZ0Px29jZ7kq8F+timCD1RuoP4Nnn
Pxg/XUWAxVdusvezc9fxvILlCT3W0dOPP/yP3Mducm2OQOB3gUsBgU4uQOSB
a2IqqFT+UP07j48ntuL0igs2dBBRn4EFZwyMTCz0Q5CaGeYXoleHHHnSl8vu
jHFnNxL0MsYeqojtiwFd/t8tV3cnCclsoC5bMzJn7hT9uVK5AKr/mNkZZnCM
/DjhErL67jQgFTgHKDDX6fGNWIF7PrqRrCqpITflay/zOouTns5fqNyyFMwv
GE9HCI6c8sfcSaYpcwAAdrLr3q9xQeo0zcWetVah45tVhgee2oDwdAfow/33
MRNsD4cmhP2hUDia0OQ26qQo3I/BcXIKLJ3CuLyU7QZRp4xKEDbdpP1u5gae
zudH3L0HralzjN9zD3jQBYhkEYPo7OvBNnFHe73lqnXGiUgJ1LdW6WmwxFhb
vDQQi1n8VQuM6oz3JVg1NZS7VvwFa3xkTOR/zp39hVr+BvaK+0ADvlIdUx4A
jMHYPPwxHfCDgMoJdAyAlZ5vVkDRQuBZmsf+jXqn0FNyJzkD055Uyn7XX4Zt
innPcdr/3KzhXwBlhKqrOoe/Hn0OVfqgPJwAGL51XgWj64k0BxbrOd1VsUyd
hnt+MF06T48YoeNT0HhGVDbnJKKs8db617AVlhRs/pXzgNV76RYm55DbmLUl
ul5AYUyqy1od378Sz4yEFMX1zA8MkHat12fliAb6x1iRaPHXutUFNaWF3XoE
nV6WCkLTJ4uF5CFqyI7bZo34m2ZjfO5QLZRWK7pgm/K6rTDpP7rLvYWiigF2
ckqlvBiVBSSqYoTJZ2HyJ1toJw7Hcq7Wdgjw0Cnp0FTrRlOmwwyeqolda80W
laEqnEo3wZAb9r/iPZP/eQrRtHV95AmJXafSnDiniRbI7LoyfeI89SXRRUSW
m02mQRfez3nVtDLGN0ztRzkuB039AqFULAOU0QR3JhaxA7k1kCJpMOtQ6tJJ
432RiI41kno1KTzNBKBQKQLr7rkkv/5IcwMTjZQ3uW6p898sshnbWM0I7kao
y2A7+L2+Dn6u0k2vXd47GlsVnu+/K2YWmGTszZI76qaFKr3Ts9MqfHjiTQAX
S3I2rNqphgSrrITwlsqXvhFRqw5HJcB0gYiJ1MfUcvyJafdFv5MGQxzpQ9Ba
X6RtVPx3v7qutXt6Em+fF1mFQ9fnfLDG6v3JXegZpBjdMnzrEH7txSAkgop0
1uBpEvFmLOXdgcq9OTRJpxeP6JkhEjeI7rMcUT3a6OJFlBd5oN9hkeL6A7N0
ruHD+05vlQ9LPZwgjygxALabDyH5wUPNoJUI/xdL5Optbx1zRx2rAnJvGErR
ukiem2I8ecNgN7BAzm6zs+5krcs1SnFwO0mErYrzLz3qJmoS8GYBMANgzDpW
2rQi1pOTwIlRFuQARDB2EEgVm7fgvYIs2O5MuTC4iNkM/qPeLp8RDmRx104y
wQddFLT5tm/Npq+2emGuHFppEl7wR2AJoehuIH9+lyI12lg3GSV3q82PB6In
4pI0Smp7Cu82q7vrf0gcx/ZfAmJAUwQpw3Kcx8JWnKtKl9n/sWel+2nqFs6Y
RLXyDfKgUurbNrQvZNJ7oAfFzg7BzjqB3ZmUxiCUC1VEDGyihkvfi/4LQQta
+APdPJCDmspyui2ZNwTfmobjibIsA7p/jwG2Uz8cv61qU/xSlcmsKXJonub9
QDmBaw83hde0VnMA4DbAfXzUpYkypCFj9AztasGfEf+TUSVymLeC98vID8mM
qQYCaj8S60gV9onz6WuHM6TTKewaLT1XtkbKH5j073URDNDy5d9gtKknSG1o
XHLvjEB/k7kWUpnnR2UkrCC5TBreO6rXRuXCURv3RdOzwDpCEtCYG3QW1S/n
/y3/FbV+fWgE7HXgmU0iCyoUXhiF7LMMrzdZGNtaA0HlIMhkxCvTW4LmQSTf
z6GjtrrbaOV/qvwbo7qqT4gMF3czfV5bNFQIBZKsMrvhfdwd3cz7AgP2m/0U
LJ5hv72BX6p8KQsi0zRcob8o+ATzNg8x+U9YlyhvK1V40v0NhM5AEPDXg5Q7
7qiI9+FzyCJF0neJHujHgsXSb8iyeALKe8W5+qYFiDohroZuvRhCHDlgCX0D
/eMaQ8wafVbzNFq9Ib9wp8P0ph9N8m/e0oHUjc2fkCCNLNYcz9UhWUWuFPyX
utO+B717u1SYqRxs3Sm8k7HhmbcJYGG84PHpYi4Lyx1r/wMNVfLhThvQB4/b
lKT3j4Cts3UCzbY0FfAKWBXAOyvSPMYlPNTuTbiYh45erDVAwg4qCPviml+t
G7MQ9rcPNmxpv5qOJUtGXf0KeujcTgU4SrFm+rZ5+ceiP9O+jxyNdwEog8WJ
lIxwUP7E1holvKPumz0g7btC7CCx5oJXvMxi8uUtPQbx4OZ9sOd1gr4Kaz+f
eadAHhuRKzB3ghd484mVnlNOe3kUgeDSkacAPEgpc922SY3m8THvrUNTgl+r
hfmWpH8qmYjyYSyb6c0c8zwfwBcU50hj9zw2yxqqtTxbb+DWv5dw/YDaGzT6
rGAhauz9iOQ9VqC8A+ScQL56q9RSjVjd21TLtljPYZc4ZSHT72zr1PYgm0/o
6f0sPjYaulc+2Jo81nv1WsT4cwjYwZt9CurlmiervA8QL4f4bihHIsvtfacn
OVL7iW+vmW5vM0o3zRuVfNOkc+8V0eFOB0EBvARnXIvE+2J/xygIdB3MRD3m
xgd96e2Szsx4oeSrekLURfA7sZjs0xHgo9BuUDqC5r0pMgxlbjDvnTllSB1F
717JfWSJLSe1A/znKZ76x3kP0XFl/vjFCACJykiOGOFUrfkLNtun7SMqbrae
RoZP4/c6SmlxYINPfL6nlt3SRfKNYPthCXbGhk4VbvTJFVsgTcd42gJN7DAf
2jnB1OuBrMKszgEyx3WYMplhKGSoafRwGl0iY5PMTK2E0HLTTsc9UBWX6XKk
2ltB3vQ4aDUhgVlDpPcALz9I9eHpjYS+tRLPV6IhwmfVNzRwKm6E3UZ8XZ6V
yZghuYDS3oyDME4HhUVy1xS3FjXNfdsfmU05NLcM1BWXA0Cdtp6Hm2f4Val8
/bZ3SsCegbyzKtZqIFea21JtvmHrJAZIjRyyaSOh/IsWNCzVg1R7H2+EZuO2
lr2XGOizUWNkdg8ZRvSSzWc0uDXJ8JbaXIBKQIQ6HfBGm8SS3ga31+HCVufX
Or0Bptc33AuCHyQd8S1UAJCxLfZZHmerpauW+SP2vcfIfobdRALK0Q66U1/2
CgxPWPAESKreC4VJ87v3d+Gco9VJSqpCRjrnpkT+pKsezqAxbMOXeWyrDs+2
c587ca1IqQj3BG5xxoq9+VHhwDRtiM8H7GVwFl4O0s9KrItc55ZvizOunH0B
wbhpj+i6Z+9/KxURsOpn8k8CKbyJmq+JhfCmwobYf93+03L5S9on++TNgqrE
wkPvPZniyuiJzzzJAFFqUP6Sulgz6VaSQtm76Dn6D6NtnaLyI04IGjiLME2O
ByjApXb9XNmr07Oxv1V/gXQM/tx7exEdQf2PiOtMIIdXthlBTbydkUbN5yKp
Xh9dp8Vp/GUCoVyg8nCl3Wi+D4+7UXan72cNkOXPO01Yb/nbUUO98luqNLLB
9dcMcJNQx2aGsCcNIBZt4FbO8eG+NxWgy9lSzkp+DhqIyVtw9RmCUMg6Gwa1
4It1uAQdFLs4JvbtfcjZLb1eE33gLV1g38CV7nP+b30KTs23gUky1HvTNvvB
eKdicfXnGQ3KmUW3/+0dGRIbv3WKYQ7coPSsJb3heHNRUPi60h3ccBfuSJ3S
eZLA1ZSXr1aI/NiP/DXBC6p+o3R3aTJW5Ii5SUFc8SJGibbeGfvT2L2Sf0I5
BBl/DE7VAMC5lkqNr2DPzoepA5nP4fh7900zd/gk1UQNXJwqai76PX/EIQSP
AWTYNWdcSEZCkKCDJHAyrKhEeoSqowdyUsIN3I5IOfIFO1sLyUG8AbHd+uMC
f9ZZpPhJXLyrGFR/ukyBS4jYUteH1VrdQrTX9QAOrgY/qwRJ69Pp3EpBhbrz
DXMTFsjEIuj1h3Cc8jCyztPJ71KULLkeLEKw4IMTEFUnv+bxtS1Zs6u8b/h3
6ZJ5pZSgDCB94rgrtjq7ast9Dbr9KcyZP1cicF0cmxErUFjK2BVuPkrKFgDr
nK+VZ1rpgOHcS6YmHcdGV083SN4+S4obbaudzFJcd+FqwQZBc4VhCEmb6gTI
ogP8CiramlVxMUdoNC/coBM/YmwA8ebpgmaTXNNpwRjv8HNzKQFIofh82hAx
tvKeDjzTQ8Zc++61dKG31AjAL8fvV1GtEZNOazfc5LsDF6NRJMUHyQGE1A5X
14T3nTGeQwi1r/r0fsjMAMlf33Z6aU3j+5hEkI3zDv7I6AO51z6juuHq7fpD
9rI7h84o6aDuFWdsvXoP2tcXY06GVyehSaqBnLQSF307477mFn0CzSGwLokM
Dce9TgWwSek+6CjqTCWCuAzojlc2tq47wFQ6lJeqewz2CWwMJSQGVkayCmsg
Qd/AParxniJusXqW6rxCCkZzBWExn9h07VOQybIws1s6sIYwg/bvTUBKfmaP
t28hM9e4qVH9GlRPXGBpa+QKKwWjXWxGwhjaxRmxXqh6imOYjnkoguxDnycO
lFpoTvjqvty7Zs29/5ms/xU7sNvsAMJiQ2+lN/SX/t+oVxQFNhskSma8/I8g
U/80nJvxZcrAWadC3xwP+krXlyfzo9KAo72c2Fu+fHODHDcvOVUDsTUUUFHW
eVLLM4skrg3qFTPcFMUo0GI4mzYc4C2rLIMjaeFpunb8HARUTwOktrb0/NFY
bt7CT9HXUhGqZGL1XfFFAWxBroshLk+yjLKaHtUTY18yR6nThBgSsOPvzXMW
nL04j2C4p/agtNdaC9POYKtRGUi0NyDqBdLj9ag+lNpjFGAWBSB22hNMTXIq
tOS4JeQHrdl5knGCtM4rt8taboh6/R6U19wo4n+ZfOwZ4+qoHgwlUI4aOx+9
7ufIWBxNdsa3QCt5laC1xhmFm+vYBmcEu88V54NTjS5BnEU5yvqn4rFM1WEV
/zf0J1MtgKBIEZfGjBg4rxU8AH1U505RA4o38ti+sQAnFq5sxlJvnILUitzb
0s69IkmwPPBMU78eb9Zn78tOCvdsg621hjdw35I6ksjUHcb+YbVii5OT5cwb
/zgko1FIjEN0Z/n/0FMZX6xq7fuAm//q2ZWpo7GpLwfvTrVYSPY2MEvcWIeK
m9HwKBxLV+CDY4vms3TXRNQ7RZTqTJxvFF5GcXm0pF6WFNExrbowUGxAQFhf
n7UfcpK594ENIJ0yKvOD9664VnLDmOBmp+bdJ+VNlhgSvVXEji+rWPKQVe3v
pqRMjQH86oIOcLMxj9PAeAJstAQMv2gtuJP6kMFicLJq6tkJFMfevU4WpD9U
fK401CO6XIA4nJ7tblnvqyuZKNohWWqPeNBSuDDSvyOLqLO3mRF4pU/p7Hzn
d3jFaFyTmCMJCXX21ad8ZrisKN3DsCr3Z/pn1AkST4D9Cye80JrKGPjwLy+N
VLq1S9so0z5F0uHgG7IgXqHvXWO1GLCUaKVehJLY5NNI44JOyHL1XpyNCpDN
bkV4ugbKEgh+5VLydtwQQxLtFRQI9gemaytEH7EaHNHEqMH2Axv/obRkLzh3
QJxoU5rTBxcZ6fWkFuUUJtTtzF37LPdfdXZl2AOUYnayG4Runm9WPkoRFNUd
3iS8VXOepG2889VRD08AEtjhJmWsAutAwV6hq/+pYF9fbuul4CWPyW8wNWpZ
0CjJViOKOCRhZtAZOZw1xldNWmY93jkjX1RAdAjv1FH3Yd8owzlTPkBKZFGW
JwG9yWuBhoTE9ys1L7Ax1fJ1vuVEmb13Lzv6VwW0ekIpUWY+rv+/l14v7hhq
puL71zFsSvu3M1hlG0EqpQrNnTzM7ksV5BwN1me0fs4y/JApeUlP1gj+ayYY
Xj6nRkMATmZ9PoYOG+FUV4nY1i+syplCMnVnTiMgtteHTbFZLDoEyCDDNwgW
9ZR4r1XC8h0YRJtdazpARoVb0XTYfXB+GXrdEuEDsdHZwMk49Cmpc5/FAS17
TGefTYYaWgk6zXXU1J3IXaZnfHIIxPbnw2w7QRjV4NjE2xikE/LsXKa3wyak
QqfHgM2rVvLGzwCmwssLUqjMnS3uRQi6m6RYYweK5DxAy1du/4cPiKQCYNyj
CQW98GvJUAIA9qh9BtP/sQV9w/isC2tZmLIMFng8nsFjyqYq6R1BbaiBGXwy
jIzP5OdFHoDU1OncZGW3gce+4PMBWwVBT+kWxbe+uG6PTbBN7leCY5jh/7Uh
CJSd6CLWaLG86ZEdVmVLJt+v096F306cmoP24UMMan53H7SH8jkqSs525saH
pcF1bKFJxJ8HIhnOUXGTDU/+33fuC4RN5Cqyd/TXE+3/D/3THJjFy8c8azrC
d52hVWlFcuMUUKM/YnxWuUJosHqPWoJj8lL5UnmWrhQt0uxqMyMf1TnZwZ3i
vF6mvUfQ/WguY9esE/Uv4hRVEkudd0yL9mchi7CWKglPz9khiECdfyui9DW2
9zBiyMnc1m8yQnpA3GRoITOJuCutMsR+Cw7A58UprOO1JVWS1fkM6NxBvqiF
9xuF6LqymndxMPL9IYtBAYkTLwNKRufywQvxfS1m13+u8FHoPol4eh61Zi2r
dlBQVI/yHxMNZzf2qEd8zSIU0L4E0YhJX+7T7WWKm11FiRuc3P90fsM71nxk
ayqjb+LJ9bslvpXxr6HhKT9tBZlFIK6p4g/tmG+iKxMA5pWRjS01dinl4tZo
/VE7HAMAsGJ06r46mBPD4+7S93NWeaubtHKuipKmSnSeP6Z3AL+XQ5gS4HJF
Zh1chBlkK9QDaS8vodmW2G1MFg/t5aqBiTKLp5Q8E6nmYsY+1y8MWrqZyK8b
Viu9pgX7xRdt9/7v4vK6e7HgTc79WuomtEtKBDC1oi5qYuJOvqwUR+jnqbxE
zdvE1J9cGqQ8Pbmtcn6+79atFxsnnrqAxTv9bbwxOBKvvnMh4v+Jcf3U2Hqr
a/gjBwFCjH+WXS47zBMQnhBGxieJBIkppsi5UMhg+GBlRe8E+lJVdu4oPCtI
7bOAOXrI/RVI1x7cbnsApQ5vBqmUIWR+e8yMJ1DWN3tdrlA+xJkrpjdczRpc
MhENyWy355IGBRHdAf1dFntl8yevRI/umlWn/3ebCe7SyGjj1YSty20UX8IN
SyKVTmteoSslSVPTWxYLLhZB/Xld+DfWKkbK8waz89lPDSQuIGPGid36p+mI
r+R4cthraCB3wsgrWnKNrr/FbNkytVB3Vz8E/JS9FcppDnQuUBZ5mTfHi5qh
TnWkEZFMxa2JPmc1bJtXPpsCki2IKjlC9KNDDwHTfCr9T1OhigyHpln7v/h1
RkNrfKykWu0KsNnpqfLhgdU/TOkox6qbIpJexR6q5YTdV8qEmbW5RsMkh/BN
ICy3+JBXjx0fSu+3ZDTKMLeBnVcQpYtKQt992KyKkXQiakmTFMcxwo8g2CLe
AGtXn4SXHgwNGtQilTShfHej+AvVThiuAOTZ12MzlwSHg1uaXEIRIuWPqaV5
h/ePZ333sst7ybZDUDpdrmEWhCe3s59PqasV88Hyv4luvqQIXYCd+Ytndd3y
PbbbkHMQJjqAsXCQQOBDf7eN8uTHEuxoxjPN/7dUXb6znb6QLsOtVHdY/blL
6qWpLajbKTZjQZpIDRMatgLRzTwA2C83TacPCA1+g0QoPJf890hYWyM5FY0Y
tsqtbaNcC0o7IHTy4Nfmr2U+mK4SZQq49L8Hd3qPCRbuQ0p4Fap6GC0hXO48
6FoBC8rA3fQRNsdhJNY7J480sNsZmnhoZo3nCJbkYc/4Ij5H0u6wR98ln762
Z1FaXpKE1xT3ABCHThWkYJSG03Faa/Y+r59Rta7l0PzN6UxxfzxFtpyaHDka
P1auP/S17nwELXJ4vquKStFrBVdIEpZHajDl4nE6XalXiKL/QRCeqtq+WFBT
KuJ0cb9flH2HSDiM0c0ydZB3cIX8Gkm8qGHDmudytnPXKYzgWvRsh/QeZXoI
HHpzUN1dgCKXD5nADFD0o0B0u7aVpOTdNTtpF17PCtrWACb9S67AKeL9dhqf
vNN1Ta7g1aD4L/JThpu4c28287zUrMsvxFnDE7+q5q6otqXAqFo3Bz91qISy
By5ouVMudDQTtyms7LKrxYM9YCiT98WOI1PTH9IYNmjF9cO1ByEkXyEzOfBm
/giU5pU8K6PfyWM0aNOnC3gGgEqvelZ7XIjLhobEEuGjkBT1MQ6/rox9ZaK8
MXvcjKejBpeSQTa/8F9dnVJ8PmNO02ZYtqwFICIB46FrT9aa1xYR0MHFSAs/
EQ12ItvqWUFHN1Dq+b0YAC7Ju3V8T1kLPzIh48c0RpIn/WH1l5rMhCF1Ij76
Mei0R3dgLqJauoNZDt636nAl26+LsMS9X9vYFP73c7QndPRNPKB2Pp9rmI3M
R6UqNO11etM1pPhiCpyaMLFa5Ok+nmea+BFJksX8jWWJ6izWl32PW0PSu+Eb
A/99NoyQoiddIhohfjN/zjJKAwOVW6Nw1n+imjfSSu5KaaNmPoZEvEHQzwVX
7dswUfmKxzEqDlD9YgWVXlK8bubwkVY5F6LNDxeY72INW63zMjgYafi74nOy
gEbTr96zC5mmIldUGwE/WK3iSBLtEN3Rveb/O29WBpW2o5ilCQsqOVEzbN5s
Ol2ZJfKmDG1fnBnDCyKXp604Qs1xdTJfdBQuiHK7qDheMdirnzZQlgrpf2gJ
9PvvdzcdHlOuEjG0BToL9nmmwIcV+a6KTRIGoJXdoEy3q3/3klyKqqSFhdEM
y0k9uUWbhHoYOnvTq/BFUJmxZkeN2xvsmjeciQwiksX9TN2kSYrbjPrpWAmS
oAcZEzdSqcSg4tKWsKBO5oY5OeM6KBofzmppxzmw2dNV2bVccYRtZxTJ4fzz
dBKnksHqL1WMTRMWY9nGax/UhanI+DjrqzBp2As5x9eVHgq77/bPml/aAnhk
YN/tiiW53FRFBKrgvsTcX6NPkTFu3xmosMf2Qq+dnbcI0GXfUMrlmSaMPfW/
tqHPP6syw6EiNc/usK9LDl6PnKS4gON765/Y9/SZ2DwcNDERdr412khg0q0t
fOCBlmsdrQ3AVvgQ+/kkYHaGMD7+IgQwb8eLEAx9C5o1eLbe/A8PSLZkGrDt
kuSX2/i8ae25DmkMroyFVw05k4dyx6K86TIjpwFapvJHBpJW8Emr7zS5rOnu
fXKjgHO+tAh6jzMbkATT7xYMt54ld2hdKlW39irR82ZvEQhsm8jj0OCOV8CD
0WuKHUaYL19XEQGFKjCMSU7HMxQ7ussrNPABFXlZY2MqZAfE0S9+pwwJY+ZR
eU6SWt+8CkJ3ztKaWa9wvP+JZUX05qmVx5sNXPL2DC9gFrKLZrF6w7baCrfQ
QvoYeUj9bB0HJL7704hiztmWW5O2JM4cBrvnLWKyRK/SRrI0dINSQSiRlpi9
+sj8hD0ROvhrFn/lawk3OytiO2oq/7LpEe2HLYy+ljNMif56buMcGBmH/zY7
tA61MSe5e9S7dmDoxCfZ9Rb1sPfkcEQ0cIHDgVt76dc0jsq0gcXHoKJMUNHw
FyznKRajulXUzHZdrhx3wTdr7ci14pifxVp2qjg3422219QLXxzE/P8u0fYO
tVcrP4zIw/5GCpsCZnnd5XKBFHm+8Pu98vaeU69AJpxtlyttZVpNNXgqZ0gj
ucp0ozDZo3Jt3q+CMDfD/Z1yjLlC+8I19YqaccJAiNG1CHrjQMSfA5I0QwfC
wtIRyRUpkHsm+TNjHwAyFNQZy41cifMf/TtzaLukHlEdUghGgLoSBNUVTw3w
tsfwyQfW8/MUcQnjcZm0vnpLPiRAgh3SjDUiotWcjzGLL+pbW/qxKBg0nLPQ
8qC4Krg7QoKvqfWNZwZ26/Ta61zWGX8qnnLIjtiPr6G2f9XOvahif7Mf1zPy
LsY0Kh18O2W5HIsrI1jbQm+HHu4XZvf4vIjSPIsKaWOGaa7xPr3D+ls7LLCA
Vx+X/yuSy5l4aaMcJoERF1U0fIH/kNfyCxuzVMjr09HTzotHVaQ9/hP9xrJF
fl6uAfkHJdIVulSu0VZ7uZ1CU4Ja0QapEsCjjykvGvGc2xDfH+roap6IzGIQ
uVQvBHxvncIX8gckddzJo1c9wLfIke7B7ePyD838I0ASImn4f/1d/Lt1GD04
8o3AiQpWfxUjlQIjEIMb7DUZaax2o+nd20JtpCHGHNdDcDcUDPE/4yQyZyj0
eoQtiuZIdzQyxwG/stvDl+XegWIIyo3sHpq8W9nKHHtUQXofCgCcYfJ1N8aD
oiamZrCN6ruwFnK9pqcgL5FYqxF9mfdsyHYN6IciZxApgxLOUaBaxp5ZoIdG
njk4/ww2ITGngEl7Hob5WGm6cZctU4VlkzY2or9s+NgZNKEWjXahm26/aQBo
J6mWQcqOjtotJHmbJt/PBRQ47B3jdXA20huKjRy3uewNDnTW4l1yDL2Yffan
Qj3zsN+vuwWtK3OPa/Ge5MgbcmXTUVWcupK5MTq0KJmlM3ncKwBzoeHmNNZL
3gjGMR9Uy+BFWs9H1j81i2LP3+mviMeYMfHmqKd1t6w44ZM8UPtsUZXOS8ZD
m5Zx9ZRnzXmgO1IhUAAfBy19HPWLJsMC9Idvd6dE0gKx3vOVgiOfMa/yEjgA
QQDIqANHMOFeTKM1RV0+xtzZTQpMmLCjjUNH9tDrdoncueFCn8IraVBVTj2N
dK1c1RKsreNF5W9wtrHzGyPoZrAQ3dVs1ydm9lMZ2t2gq/y9ZjrTFYpa3V5w
0f1D7dF3SIrlRND1NJ3FjVpGlAeJCZfkpv5ghUi4bEUkuGRZQKnNw1CDjeJ/
LdNmYugSPY3E18aBzqDlRMb2y3JJPby7RiqpUx1CVs4s+D2bQSLL0WJLCtPn
+DIQe/QZgCKw2B3swT+gcr9lK988t+by7qWF/Hr/KjeIo+fUs6/TqvmsFFhk
VTL/wKjWllQTaBu8PwdXSYVMWiJuloVlIX+PdXJxC8hZCgPtPcfd37iVEUEH
jSfW6/HZUTQXkZ2zEKim2VjnR8N1ToJMx44bi3JaUipRXgXoGPBth0l+827h
D8e6L3Q4QvOS2nCrlzUDJZI16YCcwOBVY85itAaxlkRoFuPzW4zN46FsMb0g
tzSMuo1agQy9F/rXrGDMKkdtTtYGZwbIfZHGZ4hDq/h8cJ5ll/6DFglS7Ikb
3SvOVgpnWdwv0Os2omPbqMqMgR2oUum4Njf4ePqJ9VCNTh6pUaXtKa/luQRS
AmoH+kE12jZZGqocJ5iVqL8Qlr7+Fk60aDZTB66zmZW8xz2OoKKjcZ2iisxL
xjWuRp2QmQqbzT+1Cir1zkLBTp2sKip1LfZ+WfHXkNiJiD4VLyEZxX3jBOmt
fzKZaGcQgeDZONMuwz7SlQtSaBZg+fxlzM/aVuKHMOt9/Ulpx2ytE1chiN5H
4u+uX9Xn9Nbl3cXFfIH5t7vXt/Z964bXrL853AU6bQIXHfwt7RInnJJEWlqZ
nFt0xq+ONtM+GP5xk5YHvxdEw2Jnog87c+AJ5K+iR7VQNlJVMWuAECUVK3qu
sUc/4t/WEpwxa5hpzUQcEOkHx9q48hQDlvRVBZMTTX72ITNyFlMgJebfg4DM
dWeLpfNFAJ4S37YDp0iKx205ueJNqP4j0npIlVzn521GP5JQqD8kqrvaIiSp
4P/WSl3MW80T0rY7kHUhPdqS/0MR+88FO1Ijbg4sqXMjGyXW09MeBG5Q4zU6
TXZ4maDfKK6h5sfmk2zonfAdmumW9sqE1ohOTpPBsmyoEpF2Blzt46G4Ykcl
EitPkAUFov5vu+HPi/24+9xh+AF13QI2KATkNSsLTefRha56n/OoFD5e3L6V
T7nL1Bvlw2I6XDus3b5ZJvBV12/v9YVoTW75ti1fLR7pAiE0PQGTAZL98ekq
4bMYjjde2pXRJ/hrSusqe3MYZYOSJoRYJR0xBmV+NZn/8QijDCsAhyLDmvPS
nXIVwz+bJou3prIEGuKDwSiOQZ76s+AujXLNrKo+cNYwmlF11cc3ub8tHova
d5vG7GCSDLR/Tv2TaBlSi6rqdH80OlE/kshaSniG/ihSU6gIZop4uNAMYVWi
YJKuU+EGXZ1TvYss7302PYrOurjKp07x/teU9ObtPOE7QoL6lRXTkoR1FuoH
MEY2IRyIGky2bOn/p1FFPzNfdSdJuqRuGDvtGJ32iAFZgwF+A+N6kEYY7EMB
UqIj+txDtwHWJ9GMcXt4v30fdb/4fcEtLbFIMJzswKope7LSPalmqSguacWc
fiy4MWEEKFm9bV8Zw6qVG77FCkx2wAe3t0NEd1kEnrYX6/qvmJIFqkNJdda2
rLEaQeib7vMmrjbcfu7Sj1j0xtIg4gvmX06Y9qQfTH8+iGM3oWjvtCSkTqUC
colh6Qkcbz7/nKF1M4Z/CgWqiQKu4ZIbC1Wghz0sRSi1HaOCOd99B81g7iEY
Fji2RmCM+rNRiihd1pA8YmEjU50wECRxio2OiYjL1o/4564c1R8bbQGEW/Uf
uPP66UsGg3L2MPV6/iNUrIZaUudmg4/gS/zDSNGRmZw+5UWZy9tVp3h+JnP/
CnpoZjNfY83gsvTcqwsnt7q8XSjns9tMn0QtTRICTUo6C3toWIsFjy+yQC5I
9FZtINUjxDPky+UN43Xgww0UN4P31XK0xZshNbs0/hsbJJdxxbg6Ceh5BhdO
z1rGB1cMBiL6dDj7agTXYhAtvt6RZnibKJGTulJ4ECJmsN2PjKnrCYYH+hix
pstcHqdyOQKBNIMeDxb33RMnM86MsAYc2g7dQfcrQRPR4ersy2lyNg45kQtX
prfJJwDwH3HzjB+cSrhVSYRgGiypnGsVUHXPqAVpzrHHV3TdwsoQLbDDbGYB
S7qeS4HDOmQPijMJhHjMC9K/zsEOLNe14j7QCjDUp4Efty3VRMhronvydg5j
A00O1m7Tl8oXTa6O9RMjloUhPEajSr1frsFepZiOlorHuKkS/rOHs8D1FA9R
VWYKjnx6YhC37GSyFn0HGCOFIGv38ajquxxd7D20shGBQ2fNgiY3IhjMMq7R
RhLjgytTTGepZLfo7GTFcOvzqzEN3Kg2Sj8q/hl54f+G4tB5LbGZxoHt9wRw
5lgTnq9hd2aB5rBdeTbM+tTlwzmMcIi9Nusy8piskGmO8JELmDGbbP9nPoEO
bOXCKqvKKuCNCDv4ENHhMszVn6gMHtBSSS2h/QAjKQg9ln43NCD38XatDgCm
yvfk03P205kxt2lfM6JvGZpFKpWxEBtM9iJcxfARQVK/0H8+/XNcUtHCNk0C
alpoHUT1Tj77+LNVSN+xS2ONtpGihHvFb3IhI+zeFyX7LT+Io9133t1LurGp
fuPKmywg89l/nnpa4kMA9eU6EryKkNKhBhUmfbcyuneZoFtT3GosBUFWuB92
l6AuY8oJ0HEhFKVosCdHIMjgvTvK/KP6GORPTUkl0ikHC5iNXxKEm+NQqIjs
+wnStWlw2roB3+SQ72bgCPp17dvrTFtBuRI1qCH4aFfY0XAlMVx477WA/HcA
D7oXaBaTe0ZNrmpSWRCjy3rjrfunf2fdzJVGvAWXTUdDNUV1cBIUTwJMFRfM
TwnuslHliGjLoEfH+LoKQzi4l3Prxgit+Dd5f7W4Dd1RrfUfnuBoqcWyEsRk
W74JqYaehb9INkcchOkD9dXDu4yMrwA6flMCuG/wwd7ucHMiXgmhGAcpJ1mv
pBqpdG/6vw+6Uy/EPAyJs5dPDX+ISsA2A34nWVlsWj0FpR54vbTj8NXQ3O60
5c+zi9yBKLejyLp8M9muTTBcLNufnCNotKjR6a0HPm841W/bMPpnwXN7pM+j
UoYwRrdau03s4djX7O/u/o6jv196f1gOENi2H7WqI1smGVRH/6qD+BpyNoME
WaHGeNsrTQy/ll7RJoA1nQcVA5pW/RaXdzoliZvrBpxZo8SjpzCTrRPsSlSO
/NF9xi1hWoMXWjPoP6z2DIVydUgjYGC9GoH3fXtL6vw+4xtCHvR9vtdFuFIw
c9ISdq0c5lVZiKSXZAdUObPy0r054gAhx3uR4V0SLyofZHc/nQhLBKS1GCao
BGknNTxk+EyO5cLfQrHf5oWfImPV4wRevH8PG/RC4xY6ShqUOa1Km3rjEQiM
vy9jasI0FVE29T1TYNoQe2N+l6Z4jbxaA7sNaTcd+ni7j8MrLilKwjK6ccWS
O4hEZJ7CJNwe22EwWOzRgk0pbjb/G28deSlCkOWHH2EXUuHRuGX+hB1VZzQi
BQR//apU4bo/oCK/Fbyj0S/3huUArD+iL/s4WQm+y5atOcaGfJPZAsBVsdit
2Ix0Df7HtIDw4m/LeJKP3ugauWg6ElnQGHHkcCCu6hQpgwKqTcR+mFO5gMiS
PciAc3uyBA2RuBi8w9gZ1LJ/kv9faA/cQ0h1ssZmgN9+2U0CCaOI/qLt/yNc
i4dbQgVaQPlyxn9X3V/AtvCQzW5LB6jnsPCtJwH630WyR7oNOVhP5P++D0N0
edmG+rmH6eueQn+xNP5zvfIz1ptbyL7xJvjpfcbXvdr3RDmVUGd6nR6b++oB
6t9Q59BR0EugAZ1sKJB+24mMJ6Ah2Gh2JQmf64idtkA+ZZ6Fqy4CIHPcvYvP
Ob57HU0tMUHnAeQ96O96WWZo+7jbG7QPuxDF5xIww4AVY7Y2rVOwqgfefbu/
1e7I+lUmP0LIsSHeLhYNTgGjBGb9pijIvow5dgJKanBREZ8y1T+cCFjJsG0U
0Z38NCviOKXBknfCl1LT2NLJNZ6t+b72UuLQpif1K8lQbIiMhH5x6omeF47y
KByMzWpQJLgWUKrdMLmJSzEpUw+y3q6sQ5WH8g4GPmjX4P5c4bXHaOgTfHGi
4Gl5hlpAPnj9q4IESA49O8gHoO4ATmh5Q8E9kIkdQ0neaKA6bshy0GfeorUx
vVjxTFA8Tc9YgYAY2heyzQ/mBuPkj4CZOyZ0YxC2elCqHBCTf50BGUIU1gHB
omCmm/EFsdze3icPgEYG75hPVTDv65wbk1IYEGxiGMrDBEsZRbBywWX04X4q
mGe9RIRfqdaiHFtCSvztYnA8+uARZBfF+xMrkrxvmCAKPclZ3nDEKwps0Iuo
3Hpv0rfFtutcw5AelJdEaN4VnScUsudnHasrbzAwM+JZcN0wy78yyvbc7UDX
SGw9VPpmWrSEX7VK/4+mqPHpB+fKLwIRuSCMRV1yZD8M4FLLuco1t+ln7a3i
HXd2Eab/KSXTn33etIStXoobI1k5eSVgv+HUPXXUruM2+Ieshn0nfsTXvVb0
VGliILd0NXavKj0uG65BChQ2Q6VOFShLz2/xdy3BbVQHUJp0wcMUprwuhihL
hV4I1H6juTk8Ou+7+4p0OHLzbDS1sCcVBH3tumSER769vZ3BrmGj6E4rKQZ6
qvMOtHztGOrH2yEUqgVI6ydn3Xm+7xwCs7ciUAtB3p+pzUFr80a9gqGarRfM
P1euFCHJywFdRhSkZ57dQVJdqqs3ZTS6uoNl2JTEwh+/1mJl+L5rjeJvWEDC
eCPZHyMBDQzkin3rjN/VMnTrN06YIExtYuQJ6IB1S0mbt71cdlBiJuhobuiw
SeffjEDg5/igei8nod14U4iI8gmk6rW5zQfMBhT6qwPkQvPllvUO3wTas5Tz
id4xBxT6UJsyi09UwBlsCAXVJ3IunhdzEEVvhp6u34Ki1ydO020Tbh3Gb/S3
hrjfw7EG+RvTKznjrT4zyEFl4q/Fc8IyAzjwPDxmO7lQIpvvot03nWD537A9
og5x9I0SPTVm4wBQhf2Tff0vObqrwPM8cr9FWosJfEFo0EyKsdA/RcKUOI0O
05ZCT5PW4f59hFwizet3RxIsl1MvYvRkt1RYKD7vudGDnOEaId11rHlyBRV4
DKdIL8j7w7Xu+LUVOnLS6pu8FJ0CLHESlbQ5izW8IeNxd/6SJ+81zISgHmLX
GWOQoy9ui58wdh4P0QMrAtuh1xX6qR6997ZUVS3FTHjG72NlDndmZHM6IEKs
/IJkvuDJeEhRV1CR4wslgA39A76dgI/Nm36BCB1uq8sKpHaiIknxFUhO+kyF
jtx4dH3TKbDqU7zzszhThMFvaYGtQlji4fUzCsQ9IAhpQ9aUrissXh7NU7B7
BRF/mS3FAFaQXFsSBe5eFBOGl1jEcthBYAyTnY5jYEX2YreGdF9BoLg0jE80
hiaF+zr+n4kspMK7MPn3iiDrbKai1+PPbNuBURJhrZ6FjxPY9YuHdxfTNo++
mmP4m68XJ/wvLmcjqM6tKjPNwqRWQqjzMFDLRrbiN54jTXhAbUaaxRbfbiMX
HZ+Qs3G5r6K2Flap4kQBRr0z4VG+n1r9wSO3zZLsFytQ38W2ci2J6b7O1K88
ZZr2XJ6+N4zmg7+Vl2UsCS0cJn6CurvcFmbgrsThPKeEwe8782H2cLuI6gcH
pL9RKYae1uPU88k0ZisvtLY7bP1+f3ERszQAig3ybzM4v3EfU73ocilErxpd
Ju0sW35L1O7aD9JcLNHvl+9bjbon2rLHVSAF9meYBoEp0Sr1E8XBzm3lM9RV
qzgYQr08UoEqKmlFd2s1C6peYkb6Z9gkm6f/EwpsZ/wUiN7PEk4xbBUF03ao
vd5MhBQCG9ZDLdJ1GMnJQ7PtRLW65i+fw3PXnLVOHIvB8oFbk4RKa9rFdQDG
x51kxKeQQa2I9EJ1OVLOHaJC/k2qDNeRy4w3ZQuTxVHGCK2uSzv5MMWd2pe/
S9fSYcc5E9O5zlj8+wLRWw75yJNAcQpnk2wR8a9hM1cF4dGvzlEWgcnThRzD
t4KnyX+Hf6yeLNsE3gajtETe10f8p8l6FThXtGx8yPAy277pjQq2s7YwHA+i
l98cYr3VU/fd37OvFOoPhP81yNnoYWNiuszvh+p6ys7dpEwlsKZGpo3vktaM
7u+8pKBpk/3QLnL+9XGF3xUDhKDiMWWYmgIrw1Fi3PPreDBRYDX/guAD+1jz
OWTXDPoQqWagNL/OWDf3rfIFLm9+AlvfF6ba16FF96cL3zsY8DdLZF0OlVxt
8Hkq1UApsPYcWVcmlNEVVZJe9VkULNElc3blkC678I7KpmXBh+uJkLKnJbhB
PNN4BmPKY5D6IOjBxBuWKlbp1fESM4tzX80WajId20vlUg6Wm/9IuKSBqT6T
/i7/Gce5f2U9PfIyI3xTbxQvLjgzwllQU1EoIaQBSgAZFX+lMkkzSLHAfkTB
dsjal5Nr/zRXZLbGvEnvbZyGqBVu6oO6+1qNrNm0zFxOBQGhkWjQZ4yZUpPt
AKl9rI+BNIYDx/mmK46zG1YGgZNEj0HTXt5wrJJ3bIIOJc63jW6lkdwOW9Y6
ebolWF1k/+Hrqce8N1n9N8WN21ZafXIPGljurTPsf6ShYwbXXVhQZ1rA3mvy
Oy3h1mnIsRjLLiqRksfqNjT8lOdF+Fm09wyUTbL1rcM0cQV/yEScVM/GB6t+
28TgH5cDkgMR3JlC4Zm3tvtXSGWEMlQPFl4x0aINP8+e3TS0ak0N+Lvcj1m3
8fUtgcuyYfGtIoMIi1wQ6/eeBiRfRRUOa8Y5u4NkLS5ifZmym9MPxM/k7c4b
yrwfolTYMQNmp/e9bwGhbDH4vyBS+kMrZw+fCkAhw8a0R8ZY/vyQcGjyOsQq
gPVDmqijbMwgfmSGNpR6x9grqOZQH2IKhFHpJdV9FJKHMQg+Zs1cbpzi6ezL
UqYOllpE6hNSen0NxGAehZUjQnwsPYiw3lfJHap04KLXoadW0MSba5BTSrEO
TdIZVC86cdgkhkvhP1eSKYrPUWTHrR/TjwGsEn6XM+mAe/DTng1+E1Y+SNK9
YPGyynR+CXUO3AagqlOUdn+V4YgncMK0w0Ji8yFloBtKAlRBe0HchrK1cegU
ABP8pfgx2/6CWp2JoLtJxQGvFbECBypHauB0x4jQXW+c2cCLNABGMAwVhs0Z
A9dKDY+o4FljLp5i/kuoOf8dbpR4aW707/9WXWl9N8KSBysx1AzbV8dFRHzh
KK8R2tPyQ+UZxid4CY30HgUyR0UcTRq5XPl65bL44uy5Gu77u1cyX/sK8Fva
64wH0kFCApbFaKr5RWUErLeCyROpKF/4Te4nF8z3x2kA6WhSsRMTT+gBHVcY
VbT5WE58tccs+HSwxkv0dl5i9Uy9FH4Y1JqP+Ynw/4+f7vyN840nCW2SghBR
CmKSV+/rZ7lFJp16s+GJB4svSLGyuasCeuxs/ReDSTP0OJky0QxbeALXtTUn
LcmoWPdG3pdqGXl1YK4nEhcU84SvvJNFXKvFygXRELg5IJhKZZJwJUleNBXv
BTCTO+TATNlNTP1D0yocSZA3EijDrbfLjfXC+1RG8Ev2IdWXizGm02oF1GsU
BXyee2oT/THh2Zyoq4OXJtfFKPfUGe4ZReXkLgnEvrQbg70W2zr8x1yV/wiN
hfz2CPhgVaHxlIjKv3ernAms0maqCuB/ZRLMR9dsPOlSHcKm171yr8T3kuV/
lG5FpeLQqctbiDUsnGYIcoTwg2V5TPIxKccbhWm4Z+Ov49EaY90DRf5qaH5R
JUysjwR6pt9Q4hoeM+z+idxI7rI5TCfkQc3qI99qeuUh6DuAOQTsPwn4L5S8
3apj+jUWoaUTGbhyWZ+YapXTSoVFKpkf+AFYyb4MCZEH0qGRiDHg46XrbyR4
KkDEN9P0FJhbRmggiUqIoOtabLbsByGXn6m94ebu7djmHaV/eS3C285xVmMc
fIdmZIKXH1ayKerxpZdPVqLEIM6gTy4KTipr4gYOP7oGEgBzxgHLJS8cOAS8
pzxskEoq/IcZJNN86wryYIdQGxEeFDeRX1PS8zIXyWMZir4nnKmVTNvNxeav
sSkyzne88+67hvpPvPv7ZRWY9pmKpEz4Tov8s1PwnezRT8uOaFiMalyuhwzS
sNlXgybcxs22K7U6UGvv2qOIwqQ25eHpT3OcZQFcpUNNUsH1PRkj24OTxTrX
cwyaiD0CZrfF6pJ/dm7PpiLuUbK/eVGULxg6Cv/9izyLig/BxwiVsMVkafoT
l7iN/al5wPEEAosC+RIPETvH3bxlHp4XRajDIP3AaipD8xwYSPbzDBfvQhyI
S31znIeuiNJoyet9LkuX+U49kMEJ4fGrfeHT+UtEmRI7ckAzSnhIL8sVaG55
RyjMOU4ZXieRSd2EqLjn3MUh6v0xoieX4gOoo50gcgurdwtfE4SQslCdAlk3
VhkIRsGkXnS87D3/p6k7baUjtVEN92uRIBcQ45KWaoAmRKJ8MtMV+iWazR4r
ykpXXl1CcmnWHZY+V0NPVYolk5Aq6Xl111namHMzl5UniTJlvoEPmtv+JMZz
KobKOm8w4whyNcIVGO9zA50q2ovx78CYHXC4X/GmwPbOuoarflN7lwmkS05l
jqNSIB5NIsnOuMXUw4cZLPvOxrXb9rFqOFCe4kpQdqXE7ePTDX+0LEep3IyH
RZb3NreBYMnxW+cpZNDsnGoTDub6zLpYUeCWmRBFPnz98fznq4SiIsVr4DyK
bMu6+EgRbTc6ekgx4fb9SfWyMy0tP7cbjgxk7EReaRDjp5XkLXO3hPcAVfSE
ktiUNcL7zKQdz3t9B8LQYMm/NdLrhuW2VFJAoPWaaU93M66bekTq+k2hcL4Z
aciScbdoOHR7fVgiYffJZUU31bR2yjW8LvNxLKSHol574AbZAZvHNV8BwhmO
QD+O+ZCNEQ4x+o8TISKSTQnALdZLFOmZo2sxLqcHhniP13n9ZVANV4UY03qh
26IroKHoiTnV+ycKqxltjBb8vk3nro6C/DXUxWITAMZyFs+mdR1Yh5obced7
rNNK19L8pLtk7QFPLyG5JxRPRUyeqeU8ANO+Tg3SxiYumqB018yA50MTrf7e
pDeqn4wzGi9gNWxwD7qKwIMlU3B05Thn9V5TZ8I2AtCPvT/Vv71pztxhfsOn
VOjRIH3uzk23eK2A4g9UfUr56QVJ6KtB8vuXDS+7zcTY+UnoInd92qSPPOXM
UJIAOic8rmsX3aKkA/T5nBzZhtv0dVxmXC5R2qUjJhS5/3rZB0+VUXs5OunF
DvLz+1gZOYNOpW3wbbhe/bSBxk8BNNzy9DCoZujFvF9q8BpDHjxlKazowXvg
FKFQGYngFrMP0H2cKwP7dQ/dacdyJeOKhKDOTV6XYi6R/S6oKt9qN0X3sJN7
hB6QQnK2qXAhZSnTYC9/PSiNlgyPsZs5kEOfu8FatMSP0aE7myMMNy/LRrjN
wnoDHQqca9PjUmbScKLRGLKibLZzN+TXze8Vs2gbvVRIxG+nLeup68CKtiiq
eq6wScRoG4BaJB5x4LBlYyWg3LPglfYIspEJyFXL/SJx/5c3Y74XemA5UTZB
DmzJ2e53ZVkw2ryC+Wcw6SOH3WqNLZO/vP/vaT6797u/B4p02CuSQaN8mA7T
mr9pipUUB42qWS5qtl1JIeEu1bxdSEekNWVX2u6a4Vvbyoa+iZQVHRJTWTrB
Bn+jb9byPEUX64lRDB7/+UjaCUW/HytzMnYR56No42zqkW52wnZU/T9dYsDT
4/+b5zHST85jLG2/MjK++hTv2oi44eVOu0oq6+IQvUlGB+/8+pJas+W1PLOI
1gW7GmPi6VGJTSAm8WRhXqp2MRxqtZCI2dEJCGoK3BHfwvk8RcjekTOoMkZj
Jp6hel4r8r6RSYCujbS3TuWGFdSFUqnOvLtZNJYe1Y49r3MencFBMC79ZeUn
q84cDJsRaOG/cNpiuxQhdpYqwaDX3TPall1TNPDXY5z4neh8gCr256ZVhQIT
O2hzbB2vo8RKxSnMkbcj1TN0emopsrrKfE1exE6DemI0xPnoPCTTVuBf6X2I
17PtC6fd1aUWF2mTWIxyQXe6LD0633L1FugNYYRO5+N96JHK+peRQZxPdQaP
+Rfwv9YPiYeVAt2MrFscfBYDAcpI58eSg4+yWIqFHKneNtteqb3VHAiUnmcC
IqFCyOdBCOt2p2YNEsgNMAfv5ib2uCmT7YdQBOF2UNVfWXPQyCza9d//UNNU
1NYUTCBYOLRT/M3uDJTnD06/N9+SLD73snLOh2AGijXEm5oBObK3GGkvfGgA
26EB/eCY3yL1zS60yp7wFYd5kjY7iWc6Xtnwj0lA0ZcBa+bTTW7/XOC+QjU+
Pwz/b6elHQDXXpDrYlpD7rM1RtO14lUOK8jKeVL7UUhieSCGNWoz3tzoCQdW
c58K3LHWQXK/MqC+K60JKCq+D89GTuEyoVRAXmwLj66lm0Y5OgpunzGBkFYd
6yxGR2fE7hBlc/TIXpnQMs6V+oWXtGFuxi+4diV/uA/5xyZ84oQWT4LfJs4a
ah7KUAIWk2PDqp6CCQT8lnMn8ML6K9rRO1sJNsEqwKtme8wTVDE3pfDp9nAm
Otj/CbezKsFLgmbbyz7nmkPmX/c41akYOmQSRM73/iKqwQNYvdYZBVUmDw+I
bJDT/wZlt0z7j1n7u+rRf558QYoSq2PVIHJGH4jKLldLu4tv9U/cghS143W2
hUHozAsLqhidLUpgdyO8iuBTYkMFxarLAfI3Y7o91fj4MlKGz8Er5nnLqxrE
yCLS/v92fwCyiDPURMVTfnztiIg+73xJ9bjTgTGFrQsa3TwEKuuNAM2ujeZV
fu7NwpshMQis+IoCh4boT43N7zgwN2yDxaELUwdC6AqnBeH+P6a9OQmsyBmV
N4uTO62KyPLA78ifKEuM4qphsOUupxkKf8iNhI26wnxBrcF+JZpQ6N6j+1I2
rpbEjTvdscOuA3rW51nhCVCZCzgr0zAK2zZqzt5eb8FgsU+lrAxYBFZvQYOI
i+cCyB5H6ud+mWvaRs8QsPb8xENHbOBDp8QVI2aAXHpl9N1rmOKCJqviHSwl
2hYNOnKlz3CF1rc9hdblYYKrwZUIgC6aGY+P4rNORTy0K/fvZDYbOOmmqrfe
hoLwah0DX6ISonYJVpU7wuCLbi+1auEkZ5/WWWJsw2dIyhc3BEqsqwNQzQL7
8sxYJ1aAT9wdbT+kWN+PLWSon3FYZc+WHURHdGDbI0RjsrDbgpKQMGWA6qKj
xvBVVNjqWZJvmooXmsxfMEw1iBW7cV1th8fquEY88paDQ8J7xHCettMeRbze
GpL0TQuYelP+azfAg05OoxtWWF2sRrzMW2GCeVDky0thjInyeBd8fwaVYoeO
Kuwy4sliwEe73AP8wW0uqZJX430g3P27ODU/cBTs2FDyypDfL8MWNvEsUTLZ
2/MxE5mm+2Q8BxJg8HggyCWx6FqcOMuU7LSd2FRyuNOKc1AFew3g6bxNOx02
dTDZuTQEJL+m8FTcPn45KLO5E3F+b+p+/iKX4Xg7Wehy2cO+WA/XY04WN0qR
n2qjCO2d1KfA+5ZxWdEnpYfk27BSpGPX+fi1XWcrASB84m9+mCJ3PM7SWUwk
6NieBrduLqLRGmfhTZB/iiS3ovGFtYhXXNoIB3gNVTPwdU6h6wFydXbuEni3
jdHlLhUEHUCQPlDK2n0K8HxwybTwSy9Clk2rnQaoDk7QGS2FrwOG8fUqvPCf
fKej2YkjQxgqOSqwM56K/QPKPDK/9JsYjn+WHKX/YfcNQRlwoV41TbNA7Plk
Zr0Eiu1d5dMfkSY9YqMl8omRmt88vyS4WCkwaZ5I1KKZo8jIyuvI0s29S3H5
KoGxpXV02RR8tGx0GNbUpwH2tKV0SiS1uJVPA++ONWF3HpdubLGY4a+nVQ1b
1dNZdvTF2z5R0w4+t9/bjQNSvWce+Vo8z698E1Hcz7kyqjcFkdmT0NdHMMN2
LarpO0G0Paio8Fbg4fjM5FGg9OQBmNnwDHHeQHZtLgAx86n+paoG45oPe0Iy
8vxI8GpO9crnDCVXScLcx1vuXBr3vpUsm6Mnutlvd/5eTMNTAQNVVJgHXwea
Zpi9uFXYQ10vk6JCpjM1caqfG1gbKyCLvxI93L6QVWq6EUSqpaew/T68LJ9a
OWizH8yea9h6ryOL5YCsPKrbdOBx4BL/OYr5IC5gsurPyXzeEYveyp744kPK
FqwK34qAR9Cm/hscNQffDWmG3ixVOHM1sCVCEqkIkDdU8ugkf3OUi25gnmH9
6a0e8oJKWysaH76FI8eWSueadxg9GXa9aOiqM5/IehbAyktiUq4JIWguJz2R
XaL5x5yKQ92bsmYLAQkKeruTELkgSSFNgHdjAF0vLUkgi6pKWG0M8BTewxAj
0gZ8O11B+X6pn9qOUAIiUb34VkCE9AWVBDf7EPCzhp2DaG3l27CuZDROid0q
50qXC+/iR4eR/fq7tX+5AO/vDbnXuw8evVGq2bspEY20tcT0YV6xYjkpm7zP
lzJfMTlzSmMLMwPBM4SmuW98jULOhtaUm30H3GlpzA5Fhf1Pk3bAs1Z2CO0M
lc1cEnI69Sy0JSlpqe+9gpMAQSbNRq2RIO7NiMdM4mRWUrBbTmA9OFL9bVn6
Sla1PRYleUCAUKWSYjfaj/0Y9WW1hC+KasNVQYRE+hCb2Fbtw74inZb5ldct
HlALwTSrp7QBqxh6lPfWAGO1qGuItDCTdvMptBWF0D5Urryf7+UfU8IVPVaY
IAY9dWdHxYra1Np7vOYUoOKUuxSzxCv35XQDslI7wzE0EDYj4SfU8ASmlRPw
vr13KfGyN4TIhrffp64FVgxwkpOauvBt+FRxWWjgasvlowr3LhIO1gqxJbGM
LkcClxGBaoRywRo/A7B3pJeUqIuJjg4o4UGbWbWqVQty21bzk0QBD8mbeU1G
rRcHtf5U89j43aFZs4YykOQwaCJ5WOZjkWLIG69MSbeR7E9SSCnbodgqBySo
31WlOfwzeeYJp5kjz2ihxdepegsgdicnXYXTGSQYAsvYE/ryFWySGlet4Yvb
8G2wYiAPEkV/ACoan7al6D+e9cIwAJPavkveF3aLSgv4yZkMEcgGI/gklstS
6TGdERBpDbJFOTtmNkWCLKluj9lhOtXaZsSEU8rslE1zuLlaGyNSD680RPD0
U3W1edBw6bVKFrxC/5TnsRJHzXIo+IJJ7pCeGTJqYNIp+ND8sJXeAdmGztMC
jNexOuXYEQEhEYtwaRXPKFbIsTJCQPjGxpVBQUSYwcfuj+CKuQAzsl6Cy5AN
jZWzfpLV8gVS1LuC1CvHRvDGJByEOTWdbweBkakuoylBzVOdUjjtlFGD7RXa
iZKIjkB/5TRf5U2Iq0FCN3D+l5c3R/FM/zkQBhK7koI3j5QaGe+LRaahZARQ
iucIzdeoJy6/LBZ+ey6RBSBwhQyp7VZDAzoWA6SB5x/yyd9xGJ5/p5a1mnxO
gOAQLy70/0YlgF9XUYXib4vsInKvxyw6H+cg6C1dobzsSlcN91KeKrb07iba
dN33zVSTJRhpdVijnvAGvbOvodM+MlfDJ9fwRm6MqFvUbAP56TCoGGUZr7wq
ftxztiwboSrPoQ6/Oo2DPCpKEHtYAIR6A1KE/1JbILrwOUg6ejrSvZKlvoI7
7BMeN3LPKpNJAOaamhARmsHnv3UY6z3oPVke3JTJFlxLOLuYzzphBr+fp2W1
lDMRWHmcD+IByWJiH5MSv7FU/buwOxkYMp573FS0AgLquBhEzp+LzJp7oqRH
Jvq+FqDooEeYQUTB8maBWqOk3TZKkuuuzaqFbECzotnQIA84cbVy8D/oJ7bj
ysGGpC3iniMBECKGSXs0Bk7U0kX4I9mOt3CjIoiH8f7fGNmOqCut3Y5Hgo8g
XMZKGgAMwKSYFLAzgx5UvklhVSufNTLeR66ETy64eMxwFlmPNcW/p/gSNPjJ
uzjfk/IArZBM8nimIs7RyPp1WLXpbnD5ufqMMcgDXmxmM9AL3mYnupuKzbWj
y+3Sj1EnEisbRW4hWXlaD+Pai1VktidUmv66WcHYY73VNuuC2Su1kzeuUl5o
iuce1x9r2xHORn66BAi/dv/nG0bAye957HvlxFPBNSW1R6Df9awkc6V8Ks/V
ITiEusDmaaWSQcD6xNjCxM4xPCVQjSr6V5pV/Erc6ZmKgrykkfdaJzAPAHq2
f8ZG9fX4/M0tqEp/h/inc3FVkUdcjddHrPtzD3+YgYF1O8fd2GMYUqAlFU3H
mpYWZAvwOgvf5xUdHK/yzt1Ggt3Y5pHrlUQlLelJ0B9NlrcKb4QZ30vtBvJb
uzRzKL/jrbYPnJhFjSnomNVxJphnVLSC/WqLW7SEI51m1hbwEo+YeQCmqIHo
n0COg7dyVBgd751cRsct/bzVmKQoOBbAo2rU1DhrH2w+LEtV4qClv8EIyeXN
cZ79Rl3qqmQw8lveWwKXa2xrnD44obyjfrgstcixIhwaW/iBmwFGyd9pbkMz
VBBGoeuF9a01Gnx+h6eO/489+A5hRI5iGK3K8y0pdlla+tY+BtQ5rw6Au3OX
bPkssy+I3GnYrZc100DcN7+hHDqeJuVhCKn+RAvNEcF3smx/UGWPYF9El8fD
iHaCLPlOAcVm49ZPQAe0VNDshGGgcqZiPXWOuKDv5vGCmaUUZ9jcLcPnl6k2
gSjXdH/WgCYbk6zyoTRZjur3BXZsUHkLMPHQhAJQ0Uc2TvrTfXrwM20EmKjL
fEFPHLYSpbaEWwBDOMFXKKNdmmlF+52BbzNmq2CCWYqjJGUvKOUu8R6UAsT5
PLdRzKBHWIkdmwNV/TAughkr0v7pYmaZWPFTtCWLaKlZDKe34exQtKTLeD7Y
A6Ji1YNBkIeO+7FRiwiad5GSBEsNacIrBHmH0vH48+Cn78QnjxDTBNPrJpY5
lSvBXxJZYx2sr1zjKt34X/gmZw2bPgT3e/ti8ps8b84IBgPw084hNuHMHc2J
NOSeqFbKiM+W2v8VZpt0tt8tJZx4o9Z7oSGVHtsukeDus0DjaLwVMXAF3HSt
SJ451CvnCQFq7bcgRHCyknht+VH6/qk/jeOy4qCPqfvLUWaX1tAHZuqQvalT
cdacFGwBK+1QPY9tzVzlYfCW6XxkN5lWY8nA8bw5pxkYqXDUbDkptRQc/J/l
H0ZxWziSQ8uVvOpIZPuRbE3Dkwa/HEPiHV9EUptfxzhu2h7PHavWsEXo96A5
IBRf9Qa/HaxiIGYzyWGNC/TK/p1lBXV0PFh8IAZIKuAWLFtbdo8lnQpRjwA8
AXrrsjT8gnncGNuUHG3xYZa5ZzIETq2N/2YOjY8QPSGpKCGV37j2gmVhny0y
SwYD9fvAdY03BMzZzl1x2szcNrcUE4Q9G5/9SNLo0mpdco4edVQ/luixGdh4
J8tqJm0q7A5IR8xuu3BdUSmikpgEjAOWQ7cLaPNTtHz8xlUTT1pNRfhtNnyl
E4oZ8W2spyUWAqfpirRMAqyRukFAkA7tk3lJg1wOA1QsCqJJAoRm0WZm8dtv
L6WeDsfV+QfNXwhVM7cRugjBz9wlZcHZgwqgEa6Z4lJB8nx4MjU+fyWVi6Jt
MUqkwDzzHKDexSnJ4/p51jPAQCtgX5va97mzHioAqdmL3B9udLKNKX2WSgYY
p3YwS9iPqizVnZt1+K53nKNxPiFg+keOz5/LbACb8DsUMgSlieq3c4wH5fOX
z4snoVVHyekxUihmttjShEIkXZ9w3lYgayYTrHmSpV86JCFEk8nHTIuT4a/5
wxOsH8rMiUGmp1DBvy3CL1hI+yf3lqLxdn8PG2dIwSDgd89elVmg+F9Impn8
5JFOw0vNtMbeXIwh90g6AB5546efYODMT0l3ojs01Jxq6FG6tH8eRR9zVggB
EmBENxqknmvNZzFhQQSmZJ/4MOtWml34iHbGkoGwH7bGXHNpg7z3qc8Q8qPI
WoYJ5lK9bOSL0xi70UF5RUYiogymniY+ndphcd/FZ7+YebCaqu8Yc/yXcOUI
AT0mv+Rg/tU56kqoMzqPg3s9UbxnQIlFNJ74vEy+w6X3iS4RKCUs2dLHI4qX
sbdXY1IzLb2nF8k5HfFHwLDaIyuu65yqVT7XHLQGVifYpQyllsAIuaP+gkni
3VFXu0fjx1oWoltR9vnTnzvJxI7MTFzZT+3WC5YIGp7Vy/MlFJ1LV7e9lR8i
zvu6fqZ3bYW/YFFRqMEUGfxNqFaMK/OqO7rVS9nyVx4dfo1/derJYy7yqUW8
g/itL7viSv6vdGZrfcOqCc94BsGZrtJm3jMbmxqz3iWFljvP3hgQLJ+vNf6q
LrzTRV+rU/KWSoiyBu1fg4q2NO9k8lAuWnjaiJIz8xXk9qK3tlaitpRtlho9
NL50YfEYWlm35dZNrXuZSS20pv9eAe9RzGa29OUHB0eM4t4pRKmGb+eD5nuR
xxQs52dGFTZm/+z35TdTgx5udX1UvZnJt6JMQJi6h29XM4LU4nqxW+3tErjK
wLoiSqmonF7W/knDX8tWaca/N1MKVo9Jw1JUUeDQ6NMrtXhrbzWfn482blh/
5pUiXoh/lFGIplYD6BIFO+5GNIfftZncRj8IwebGSEuYXiq0+Tq0vJcRUtc9
EBpO4CURgCS5GA/Z2rs1A7uAl0EOW9u6QZwNQMzOnglOK68wE5olViUsifQt
82mBoq2IS+xB0SfaxtWRZFz1knTbZg8E3THxQ0RWxaeVdL1Za67a1buJLrbt
y8DH4gywZiYqKikQuiNKlLEw0rcyAirv50TJvMr/hnQfnJu4NYSSLfHTerew
UiKZVXvsDP1fRd9GeWJYegj/dMv7YHrmX0NcnMJmRurzpzOH7NgLm2fdoYE+
so6dh5LBf/3b7BaHlqN/wHjrDyKvZ7cNRIVVVQ4OaSMSSiSl4fZ9myelpeQF
VCJia8JHodqW/aCuYaNXcS+ezZn010JSh6mXBepXjnlZZAQaqe87vMMf8Vbe
oLOEFbrJONmUvxLgx40eHqxBJ92VnH2g+oeQd3CDfpYs2IfPetgxZn0dogGc
345pNlQ14m/nm8qIPsNvbYy1abEMQhNwKaxUQy1neK8ylibxKxtcWl3mmhaV
3QKbF6J/OB+BSeyyIsZjX28dAhrNMjk655oGzsAeGM79F20/Z6mDYdwuyHw6
euWptuj29Y92gmJ2k/+KIrGXEehXawge5kmW/fkeL6viOaB4rzHCVf86ElbM
knwsBkdFQHJ9Md+iwIvHY4LQ1zj2mJmR4wr5PtUiZnuO2zEiJXuE3syZruwj
R1MuwI0tR/Ysi13wWHkpBprc8bVvJU22nW66qqUjR+1QXM2wjQln+9ITlx5V
SGetbGoA1rDQUgmB60dHeIOpt5dRrPO/CZOSc0IKm8l77euMkpYt9D0GjO/d
6qOkujilpgxR8PBCwGq8EfvOUbm6tWv5Njur6GiS4SkJVLAcD4CoPDdiI6dl
zEj1yUy8nl2c/7QdqB5RG0N4ah7C0sXQKHKRJVEFPRWcupgBtRRGPetW8xzG
awuzQp/iVUewTF6BpbqCa64dJVUSZwMi6yBPGfggPC8ji6XiV7hJqnUsbcoe
4UeWdnKAJRZh6En7WE0NMtK2yalEIwuARtYppmpcKez/Bgsaq5xo/ZTNrTOG
dv1tdwDjTOQ7kzahiD4o4dtvrBnKpE/oc9iasH1OrcFj2DeUK8dc+TSLSinL
I4u62sPxkbu7s/0VtjIU+N6xnxyUVq0sAu80TBwHbL6KnopVuOVhRDHSLcZK
MlkK9KRjtoEwRVI8CtQ55xEo3nXY5w7oY6Y39rnkYXWP6j/i7x68w20wIdJP
y90t4LqDsKRo+Gl2MKWth40SSpc8PNQAOxMuGhJk7bpNQZgTezSAFMvL1+Cv
QzMUg36ghztPR4EXJKJtWxDaW+L3vzfMB5aPfxxBc6XvLgZ25s6035Dr55L9
PYhlsbbLaVOdt6HtzO33oxkTpFt0QkQdTq524ZiGAwHuJp0CEnd4JuPQIxMV
3YqqTfb8BDtwdKMOgEbAXT3n6L0LB5wmberNFMXtskxXkSzOYrrXVU6cLpAs
C6bzNi1FM3XidME4Qik8d3aLj6iz61TNnhLhbJ8rQNkohdfTG3w+TM+iRv3m
584jl1C1iM0ysuYck2Sny4lQcFXkVJvQOyOF2s4GvEj1s6ah/whlqD80Lnls
WGYVExXnlTpuP+glG3b2RvXSj/F9Cg1aRlmgajzv1vyHzIhuEyc8R/dBV++z
MrG0NgMkFbhektNwGBYTFEFRntjF02orGUMwM+w1ENPTmNGG+Ujf/gf2lQy0
Z0VrkXBQ4G+u4aXNhbeV9hzQZq7nwVoTWZxxotXhxf+FHhFhtbzp3iFbtvGG
xvsb5keAvD3BXUuJuEwPtdWtThYB1gXHjILMe8eIqYULSVnisbpTi1rRKONe
WiSPyUq8n5aMo7Ia3wVW24NCoYWa8WZGhgQQvJPcuoVIaY/TOe9VKUHgu8ex
RRRxvL6b+ZqpKM1XBMLN67waGvArAYN4FAJwUZH658U6qEHMrkHVK5eP/bzl
2NXkagOT1ffeUTo35Hqe1DPrajxxdnr/7xRYl7E5ppha/OTeoo8ib0BABP0+
JOi6IN3TPL7JjWYJGM1Y3MIOStgpth3jY55QMQntGwFJnzxVqYbcFA22ONCC
paBPqSmSi2QumEp6qKhDLzjVTZuYaMC7vmB2O91rG5McIU94Q2zXDFhYQHTw
M+wuGkzQkEvAwn7EZPZhVZSoyJX4UNb0oBjW4bkPn1iGxgZK+3uDyyeYT5Qn
SBdkj8oYmuK4VxuwigG/DLMLN1zJbXiLFOilEf/EmtQVH+uXl4oJOD82uSiR
rY/ml+H+yoYQbmPFyf3qiMIkbf+JfpqbGFJdPIiVLfj6CTLj1ApVcfN76J3S
7ZoKafdPHPyT3pj7Ywsdr9SHkfdvctuFx5oaZzukkoK1TYdQfkFZQVwv8/he
58u7rX5iqmqkSx45pxFU+2twsIVGqSWkEQVVqfSfo3T5bpq+JWE+az/HW4EF
6aAvdxjPl3lpL1CRlwuJJqIZNeuXBMJAs/zqTmca1kQjSAhivtWPRSUn5O/f
As5uwPeNW3Tl9VsV5Zg+IhBtarHahQ5U/EHzhcNn9T7sKCdXhjrem9Q+Hz5i
Bk21fEuISwP79J87pLvCc0Kt+SenQiWLNKEZW2itwqXivDg9Rt0VCbcFqJcc
BmuHbqrVKdVXg9VQfkEgKmmAFA/Vd7BrYRqK171l/SLtSDaiBwHjb013j2vs
g4NgOM1kkvkrzh3D5PkiRUYIqBsQUDz13vO6OcdA42Gr4C0qAOFAyYoEUriC
IkfN7PwjohRoOvVil11w0NX5/Ieaiuw0bwJzDip705ArkSNH5/2C7Bqo17LK
WSmsNUsMw+iBQleQx97D2YMidpVCpUZgYrNlO9roxrqmRQVAtzWadYpDToUk
FfIbSFk9UYIrh9/nu4Ja8HHUWBYx/wCxltmhpF+/I9be0PYn/Z1/pM6sABtB
gvTBfZH4QFzXTqEnN3ktb7nEKWShQceGBHnGA8nElShnfDqpAk2W2EKuhH0m
XPGh62DsSTBD39qKQyiNaOlEU9xb+dsSfC5KSMJmMSerQjK/FJTUXZChPrsy
7LuwuBWEJ3/U0qWbpB5lMG2NLnsv3Lz9q/C1BYhWpV76ICiR/S7PudLhgDWu
FXjTbIvRsSbaVpc9TOWEjq1UvjFLlHm7nlQ4GgrjJZVEwzTYNUC5nwhhN5Ii
WKgXo6onMOuarIvLvXSR56WwlV35DUjZ8dhTQtufs8kK2eyc6PKBvrn2bfiB
35CXtRG2CA0Qdvb2FDXvhYwvIenNIkUguWTOfkZwKxHV9SRAlOt5kjTPs9IC
wxsz9hqt1vUr7aw3mJaWRC31CHGyl+tUP+Z4u9r8jpgv30DbTyKnbZhvPYRB
l1kR8if2av7hysn7ECp+KGNMyCKvePEiI1S2nXS7nVYknY4yjFHkqGGRjF9p
GQs9LYYzbaQhRZopmBKYunJGWE/rINIKoPZ7RHckOtoDVxAEB+33rAIRrXAA
+GU4Tsxap1GaSjROfGzJolyL7GUl5OfM7IinY5UxuqEbwVCpjR3cxyjG9zzz
za2XANSiAvKF79JpF6rNTa/lsHHmk+EBRuzYOBVB1Npifzv8mxoL/Ujx3ASF
wu7/NSnz1+pSHnrH6en71TO/K0fCfUgCUlQKNq1E3UfRhEQLdcwbZrucivv6
SoZH7XXHwdJ6XHRguAb74l/+oJlDHHH8ynGY7iBsPr0ltzWIy1Qu20hEVlWQ
kUvLxHDMlt15Pd7bAIZnzGfdWpvNFl6OY7el9xwMnKjBEoqKbnlZkI/WtQIy
SKPsrRKshmNuJKSjxTogHmjtSYI5DQi7hqTGRKvXp7n9BwwjRZl8COGpb0Ov
McBrNg23ojWzz9KF8fGqsxM5ip67FDoHDpMqj58G2q1FaPZyB8T/ppAlV78Q
T8MUDKT3yG11RCABIF5s8lIVRKPDLGKFKVn8WlTyEarK5nPmUOPsjmxAX/FI
KZ6xqovE9fDGES7rDgEMytXoHwCBa/Epfxp3ZbL9MmRwi7cgb2NSpRSyuImt
0a3NfbCv8HxX+Erf1FT5KdVeWz8ksBiPBPYXdyVjhF4g1UpJFxAk0mHE/KIT
E8+MUnwRHauqhlDtuCfaEyC7ppXrcqf+a+81LG0wBoXQHLrMF+FBkVNrWgl2
zmRyBeR2/rCEOmmq0CufHJD/lFPEYVAjIZILGC3afcnO3drF9MjfBXkriqBX
Jn7tyn2E78DRjPx92+lhvQfT8bg8R/fcNohAxJYgNHkI/bnhfo38Zc3moW/0
QV9IJ5EWIajokRoWIXOXIVUbvIKJkvqR2JLazpHuDjCsBTVdMwmYxZilJ/rH
CSmsKNN7TyOvzwhpZUUB+jluCT3JqM7PDEz6fgwlN48GqIeqHcVClIQfY1Vr
S3uJ0fx9pYx+WylBvHoL55cUqma261b4t3UtSiXSoo+Y9B+lTxp+quCHqwzX
mVjX2Lw39Z4t6oz0abd0Rj3SGFMJhS25LZYEHq/POcd4cXCMRcdX1WUhk9b8
u1slgRkFZuLnSxVsexXyVyVSB7zioqhn9YjQHi1KsorQ5jeZXFxRX11XTn0U
H5LWxw4Ixf2xEFHTjpZ/YVBtjeqgnVKxDIt1o9/xxhwQ+8pVadAy5LvwgMss
IAu8sn2xsb9IXooFGQKsRcciKNqU/LGE1W+aCxirseHURpJ4gGqZEjoMXE2L
9EZNl7mC3I+Ldf11AyVFuhMjyWeDLJXf91/9sACzSjcxHo8SQHwSZDVh4xhW
fFDa0jrES4e0kJ88JxuB9uJfMSyLsqncGsUX3lXybYP8ZL4D4NHfAHvK3Mny
KWT/5JMmeHsUlGH7sAUXZAZQXVZAFMwsbBLgEzpR+jEshjY6BJ3hqWMHDEOh
A8zoSi1OINNOTrLB0HdMg2VtluDq1zR0GxiVzwE0+AnBYEzHmcHYG4S6D6A2
KNqcLwwKGSQm5tr1NOVZI8AMn/NjWVfAwd5lf6rJOIA6u3AILeeaTLcGc7xg
sATbo3cWl5mQSx+Ee6Cs9qlILuEc3qVW729KntO4tciIK6E5CBvXF2DDnBOK
CXyNjnhweSCNR4INyMhiDnrz8MMLVUH9W+JHgJafD1OzbjBCeZjsVjbHgsdI
PYnF/dGRoR2XprWMdjwF9fn6HUMDGaGpZJgNZNFQhaN/wxyNkPNjloz3u5gA
4hLXGVyrIHAAxszNoLU1g3DsNSXrfip6P7tzCjl8UZdHY6YDi+lDXkbd2Yio
jmkA0YX4eRqUdH18S+xzvE0kDRfc9NqTKEJ3xIcwUh14nlgynAlj1VKga6O/
Cfr6Q4Goi63m73qUVcDPpxdQit/oNo+npCumKU8BHo3NWYNCaDUkt7fSB6ex
1ilFl+91g7D3F9Cf1dhERdyMdhGFsmpbT6mtQ57aDRzG9iDfhTwF0fvyVQrY
NnZvoiyc8ku0phlEq6JhlcjkaalIuxkbRYV+HDaVOinEiiiLjZcfH+WF5Joy
V3OwLLcYiq4FcSX36dp4zLtJd8eegRb+0wNCXdHUU0GhoW4gEcshcW776B3u
7c6hsLs8b37EnRXrreLtqvyteOX5qjw5A47H3CnEupcD6N9xAWl6tk3GxP9L
snHTz0MJo571bp1gBcG1bc0uo6zZQMBtRL0dzF5t1fRNeRngX0oMx+njD5az
H2Wn5tsMtmTcv2jhsGhDC3qFpmbZmzXCCU5eT2KxXxGAPRTRM05Ea7KXxpkn
cX9DDlarXdD+ebrtQxDdLNQWrYDByhnrganE81KtnG76a9RGngVbzJWPYenN
TH/Gf3ge+ev9BeQqP0VraZQpgPd5KtCqC9E4BPkh9j5+VvUHNS+jOmQhU2ch
OH7U/MH7SA26HmLl3dwLkPTzV5hOLS/niOLBB6LwY65kT8hOmNBzFqCmZfs8
hQzu58tnaBOs6jTq+aQKtBcV/7vfKtvdFt6qApcJW18p7BJnzPqar+DQ6/W1
m6ViCprpO9lZQ1x/1nGQYKfHRORl+dONA4Xg8ThZr0SOEGRTpluMJk6TgvJo
+0Km7/Uwt9Uwc2WDHClfJy218bzUiLVy9bs7dCqsF3MB299bA9ZoEcr+fzy7
p3oUWT8+QYCRVMUGpIOPF6C7WRL1X61srkOFyG6qDSGamYtE1rwZU6md7qiw
efq2bMHOfUcS1s7ubcL5ILAjhK55LTskYHtpXvQRkAn2J6RpIZE+qJX+cfz6
1L0/0U1XnmHCBlxZViF5o1qvMJQd6Eijss9Mv/buYOGizWdgMwmxLDVcWOvS
ldi2QczntpHP+AIi/wKOmoM8O5Ri/KDWTSdsJgaUUiPTgxCLbFkmMW9MBWrk
Y5lfKmpJpRq9Y7LCPZ0tOXzs+Ul4rqMc7P4YmQcFy27JmXs948jU3bwaavSd
R4DOADanE0x6Y5D1k0SBwt+A5qCiTWwMYABLCOdEpg94v64o50H2vEuYyYbF
9/yDAfdIn0ynzH8Vpz/mnYFfs8WkQKYgeaVlpBtQrY0WSmZ6Ckc5HNXM0/a4
ADlJl5kitK9KVF1jRtHgWHfZFILIu+JGRGzKI0M/abESBhSUWlpFCyl4v58Q
OTnNglHKTz5ht0OK87Jta0dn/ceTVBFQhwIVlDwfxgaLuu4liMN7cIvfnabj
USy2S3kGHJg18D9vBwuNFPV4FWEByIz9yJ18HSo3rAiCDK/30waMm2nlZa1X
2sTQSWsGPTa0gWGlxcthG3aXVGAd/NhYarKscYqFlZtV9h1xV+2DIN6aU2as
MSfxx+9JEUrnH3IhJaHls6I9SrMEUagvvRtYsFPuYyjtcGpZrxcYY7vHGZMw
NLLYkkOLEtL8ifCO2yD2UOYBYm0cu9ZF+a6COTBf3eTCRPo2bB8fDZkLXH5E
QywEg1STZ4THRwOH4pmWbn6YnTUt6vsR0t5Z1wNXQyAJq1rrKZzr43elsjND
DAxTqt6DXm6OAXZr4n2vUlg56a9jxFwlGSJBpBMRrgb2UvxdHV0qyjj/kpZq
i/ixSBzIv5Og14Qx4WuG71jVFbNvJuWqGD8eWborMcZ1EAGP/rxgMDBIY1pt
I17Uh0YbD0YyXfNdBwZFG6p1sAurdgPm5S3bLbYLT11rkUH6Iu95PII70dwg
bY9/Oq2ez/RgSLjUMk8XPBV7HCCkjUdSXiUJg4QC7NnUAB0btDnoVa3Esh+v
A09giUTBbm7JR84ZNnHZXKLGmfw2rqyaqGjE67o8Pi6NebyO0C1g7VVVVqUo
hfrv7UY21z2N47e3gtum3AIOObeNz8VE8XPyAh3ilEEUf4Nt9zPKZ/51u/Mm
RxZJl9llsPZPBXEggE6UjRwQJGCD7iEXtbgEgSocvv7wIUiyj+ub5EYnpuNY
8tqN0i3kOjBGOYeOIC3KvcyLwlnMzdgb7vazuc7NnsmXp5cKmeJNblSQejIt
F/FsWSalbQit6Vx8Mzd3a6PwT10DlrusjGPC8dKjc2GBD3KopgryPUaI8XQq
IGXR9xyQvG6imXCIhkdvFT7sQ5N4zHQAQ51RKXSYq58EWfmZ6tQK3VK7J50t
+fltbfBx1+gPRKNynZAopX65dJFOpBca5iA6X+K/mBBq15DS6fIXzZJxvfuN
P3xpsZajyk8UH8is1PNikcRUk2V+2IFKPR+7q+wBmTFdOY66Imqn5H93UFsI
5dI69bGYOW82AOupkKdFcIJDAJjQlL+hp/sl9Cf/LrwWkJfrr0z/Sbcneves
QoKuliGVqOocW9lsrLHoatmWnjUqVJWvXSRma/ZKNQm9p7LM4KXVmbkTSoq6
6p2Alr8IyIDGcAsmYJ2t3CYpQh2aimmPY+mkZ++mhyJe344t6GHkAJNLm8tF
/Zmd1UBnq+beGVdLxyJ05YfkDrih7r6+RmW+8sRiEOPHltYKlqIGHcjFKbD+
C1Nr3lRxDxnMib0AqICcTWNVyazySuFiKVCR2kPnvRRt5FusjgY2FR2fGINV
DM6i/xn6Fg6j0FcZq9EybwfjpZNqbvKZVv/54KmCq0QSqnOS1c3rI8eReiWs
CJaDzLpJArIE3LKFUVaXyJC5RCNkiaUSEMQn+ihNikp/ojfNgK9f66Ipe+NQ
fQZUQdRpbK+1Aj0k90ZjvzEQNaN/R8S7Yez9zIFTAE38u2rWbLzzxzJz/FCH
uC5BP5Fa7eZ4ALk4A/4A99ws6QkE4NlHuHVfkcLRb82mi6Sz3/Lu31iq2HOD
EELj/66g8qIA5v31FJsZUBCr8qyOXDrWoy4RYYnkrHftwRMq3VJiurR6h3/v
cMKNK19U+kxeQ0eBASAa9BsSKmwvTlRuuKWRvrFEZ67gnyPJza+OMbVf9XSG
FYgUOqVMftgLBDPq1BM1CYf965XXc9wdMMEaSElMA/yOOnbAeLLkMhfBz1BL
nOw6FZRCXSie5x4JZdVnv08RD8mDYfLXX7fnuVrDGKEOYg3EfDw/7hHL+aZn
e63vud4slrX5wjs2092smSWFi3O3ITBo23RV0PR1mvDdwiVw3K5Ba3RKGHR0
+9UKdrtZk27imwyN78VdklEvF7GRUTad4bNBuk+egV1uD+7eKjoXawjLk2Xv
1zZvTFAwWjU81Ar/odNDE/MJyypNe2f118ehDoxEAX7PVoaFv+wpKrHcJSvE
esUFmz5MGeoX85A3KH3Ff3oRBGnc+wrUklLQP677N7axoDJKrzq1pnYjlBMU
cfMNee9tZ8FoXZZLJDPEdC8UfDhGvYcwiumiTfgWbTulG1SONyVxP669adVJ
Drk3c3ikW1K5K8iFj016Mlu6vi9P2Ht7NV1w9aVhlI5bNZiapAHiUN0tp4w4
msodIk/Vors65PA7gbjY6KmmnvYaCVinKqpu2G4dyyU0Ps8TRMlQIB60rGzS
T2TrE2TEnv44dvuQDW7A6bsV/tCiCOMKX2eg8USwFrHZdOwATwJ1LVyoUgZ7
NL4f7QwHx9zksyMpGotMc4lnf8vHak3LyDIw/+dpjVCMGugA8PV9KumIJUkQ
mEuhks43VgM5pV9JCiZ71xrQwnFtuLEI5nCXrwmLMviRDcT60kBAiEE67ukp
s2YrlW89iCwsiItDXf/JyS+BEIFoNGPp+L9QdZpNKHyWtaXQ5ZsqprwkM+rD
JQwkG8EuEj0iy70FkkPgg28H+Xn2HzXwpz0CuY+y/0XDKIK9mWW24PE0nDsT
s1mQpFhm1BHOrbTYo8nnl33JWLFAqVYokCoUKwWuI8BfwH+R/nOW4Po4+zvq
8kPF5fw7LObYLLBkRy29o4eOZaSBUUP5yP5E5T5j4ef4cdTI2Fs7C0nOddRy
l3WRttDmieSNA4kI5Rl3R7N3NyJw3Op0Gr7zXDOfMDVhEJmQPtFESZ2xnoCj
FhVTzEaBIfi16Gj93iol7/THJJvCq87W2mLtvWsbxXWB2hhmCO4fdqamE1vd
pKezAGm1zKxPUfKqKhJI7f/fSvaMGExaf+MZp6EVKf8LjprjJk3miAJKc3em
EMryLcJE+hwfMVI9l+PqBB5g35mwgt2Dp5GvVseLMIh5gCzMvL3JyeIkPy1B
OProkH9o8zqjlj/5QYC449GrArjdsSPvaOZKNhPb3wJXHxZhjuMN40BgNtpQ
OD89HzksupS/ig8kwZ1poyIQZUy4VQss8Y9gQrNS05GP7didLPZJ2defKwyc
iRbFJPJcPdHLJp4V47EGs68gRBG0pCGP4y6fP+i4hBdWfWqr1PjiEks3oK9/
Mnmpzp2Fb4K7loAdciepkA/n4atKPt8eXu2Tr7Z+5vpEDH5i1n6jk3zDCfQ8
bScGcXRfgFyQva/gcKIUAFYSbitUQuTT0p7pVslBHvwu7iqvAG6amyITFCwd
r5Z1LxnQjLm+Jjh6+BvSZrUhZwo+bOVttuf1MNd4E9UMsJSB2sUP5iV+IRV/
x6fVrL0kmm0Oo5NCWeD6lovIzvI3SrohwHbPUcDtcKfDUuADTc5Qm6kwjeDS
nn+rwYEnisLmkOIMISLo5Y4B6BWw+HEJkwgdRk3wrqJWITP+S+40eCI3yfdg
bqDYWVwxeDv4P2mTP7D15GLppSzybVYyez2W28GwKhe6sZJlPJ6Mk0LaE3if
dPe0h0qA+u7KyKOS14aiEQrg3kDmzo29/IOreeS3BqA8gf4rwBlQp1lNPyUJ
FbUBh6+vzSK+jvdyy9P+n5q0ix++veOTJXi3igax7DaxTESZ3vjdBEU7cWgr
sryQVLxZjKGlUwLKOd93dbhM+bAtExgGd8fqZwpFOPJB5lYzTgu4pGkENpry
zcwAn8A415lOcoS18w53IizomhZJKpvgnZAMbUXSKAZh6PYJObO5IXdnLRb8
HRQx/FeCZJYqnzW7byhOVkJjfkvOAWiQUnQk04dteHmWl0LXoZXuoB1ZSsA0
bh4SYEFFDfDZ49Oafcl2zZep1p3VLhWv4saKleCfHg6yC15edzVOwTK0eOxn
aMUw2yIpjuW7syNQNzth25K90cCjfKHgagkbYu2JjpBNpBm1QG6APayHQIiy
XimmCr6/DG4Ct/tvpK8sexhTkyFYW8+Xor/MVFZE5b/M1R1EdbYg7mKYejgm
I7Dktj15plv17EpjFMpzjdGKeNnWxV1vyKmjdo0qc6ntUIEGh1yDygXpYxea
w+xQszulgzTSJl86ytoR3rEP9tzAAPEqGyp9GhHwkR+nejVYL5QTnkxmnsnu
gq0nXtO+hrq8lRU05MR5VjYJZw+CaJ0Cjo0zQSQdgw1lar2PXrISCmTj7SuK
lCOGwtMBDXVmnNcYSMQYyNCQpHVOHn4Se9wB/T56MjrWTu7Ypj9gmtmzuxRR
3gOuey1fOZgPoV0Fz4dQj6KLonvHQsrGkUi0AOP1BMAhTEc2xeS2FjaSCCLd
53o2Y0Nk6JOGPrZblL3aCOrugtXAsuxGyH1/nX/7UjsRpxVtw8s3fZsd5ajc
b8h9WBG+zO4b69H5QLvSLr9pZYEoudJhgObiArcz8bZlYmd80LY3YBapP7N1
vemTejNQvxsiwZdI3QQ5VuLcl+f9x5fKUDhtOve11DEOZonaiSRcaPf+liOm
N2LxY4OSNTYGtWHl6R/WRZyr6bvFXzrgCoX8NA7XMptdbb51AZaEK3TprCCp
papKt/L+gaSW8p52JOe3FkqYqhWZes7UV8GQmq5OMaE0lynA7A62pD4RaTuf
MxtNV5ByWuP80XkZgp7KEgMWZiQ2nQztqsAIQJLrszLNIvo2dt57AV6SFzCa
eJ/1STyAgf1+xKNAxg2VgTL+8+mHrAJ8ZXigzLuFFGEhO0URK6lrmrQIEvBy
He73Ib5yOG9oalR89a0nY/RgFMR5Pq2aL5gm0UkVe17YAhicmp6AYCsOVBNC
boN3mb2j5EFmsKyPxrFbK+Mdh/N9ftDFLR7V80J/9Ytw8Uq89IqGpBfkk5s7
L0UuaiUSDGa6i9g+4zernAs4qbXReO3s+UDN2HfF1OEJrFWPkw8zAIYgrBDW
g3z1l43gO0UqivVmlFzQlaCbmPfNJThDJyrQbyS0wmmMCM2wJHb4D2CVvfqs
4+LS4RhiEYJYNK4W3y0Px7XAVg8xh1xIAOetmmbSWuBO36FU4E10LOFgYbEy
1CQJ2wZuP6gDnmJNfufMVePLzSvIo1O2G1DEr6oLbbWDYy/3u+uxBeJgzcHR
mdafNR4e5mjpokqG70Grt6Qx+Jpr3u8kkyaEleFn8fqThdJ7e7+igiRRDq3m
oLG7DqjBklnEp7FXRAgJysiAbiNY+OAZ+5fbh2Ikhe8zql0p2arDVJIOI0L6
+TFphdz4Q0dPWna1l1pu50NOzgUBE9Ef1wFQ7YLCCklhBL1gsCFyTCFy8gzP
IleiaXxEtRomfCh9A8FIMMwR6En5kqDLGbDR3foQA6NoVPfPvaZLfhgkUV4E
ZBn1Fskib+ZMqbU8vCMbgO0II9YCl/bk914Gk3/memRAQSoUx+XqcvACjlh/
a5qFUWpgnCnxncXHyWRfpKF4zqXpTSMkqFcB6+gBRKJ3MJcW61hVa4Xw7C9n
38NG1pWxODJUuyMKYOZvvHPxfT9x+eRqvZBD2P8TETgtmYQnybKdi5v6hAtQ
8hCYtQNIcCiWpWiNDV8bzF42N2VCky6V5JOoK4A1C6TFxmuSlFDLG0iLnIQP
0pf/qesN/wkE9uvJGiajywJWRzxl0Bl1oVX/JgxnF8FKx+6wVbS+e7z0L1gR
6Hvz2j5hi9JT7kR96pws2q5H/EJnSeycKPD3HD1DFmzk1+KhLLgX5wwBAFgW
llLCauKBPl3bexTqF4Dw95QB6lWOtnlIbBpRYtVuP7r9pGIcd4SwX72vFbqF
lkJmcmP9uYPVNnj+ruhnEP07uqc5sRN3kqEDQwMsPTYDkxiea5ZareWTCGVM
nQ5EMycN6xfqPmmPMoIW94miC6MU20cZM9iVM5InqjnFBfI4jbon46+D1WIe
0qNjMu6ehTqipq9YauKH2G4xrGP4mTPGf7tNSZIzAsBGpNYlxYcf43e95rVc
PtdmptnItNDBP2tiBEbPo3iOJ6mrKNpeE0/HgLlb1ObaXQE4zgfYy/K+QBLs
msNS90y7mOdyXMHiXT2LI41ZC+bqNgz7e0PnmRg3fjdbY87SPnk4lrWLQiqq
qMb0PEZWO6gcXjZfQfUtrFqnvxb7xjkFuNlJVpEvvGIHiGJM0hXZSMpi1Q41
ECcs8s+AX+8GH1PHGx5kuRXHfQc5Dooku/PQ7PW3O0cwqvJC3GAlrLR8BT6r
kg8K4u4+ia9T4yJx7Mt9ASD3trHSf4ovXLWVlz9h9jiMTGJxERJRbsIJTECx
t7+SpzHRtofdeDSztYGaNEGdxra6bFd9SJKhW28Q8ED61wYWsx9PNCsmZx5V
GnmU3L9KxslEAYQ8oHR1IAFwr/TU0B6VnjZpgbqxpRwgTXVylVvwASRvF2u4
tyUZu6RfqBuG40BdbAh8zj7OioDrv3+eYXBtH/epnGxZgPvTxMSRcJ2lDAfc
O/KiayLVnAtGdLHv4pWylzgO0c3jS7zK0fEKt86SXb1bFb2m053qcBoHrsHv
wiEJux2LI4goe7yfZODHtOMSkTPKO2XmXStGFVbX8vj94AOWCjLAeAqem5sS
m+pPFBjN2J1v0A+4PoXxOsRwjONIlBBHteBEmaQPCYKU5U8MhOE0SSwA5nyP
vTCM6Lh/CVa5ap+vJ8cMi9bsU4XGZm/BGQYong9/Ny717qcPSvYfPzBfU6qo
EFdYBL3er9llBYidDQ4OEKOFtKSoobIXte+KBXdVW+uRBCmLwzMA0xOCpvAh
tbbDwcOC+fnApAfr7W4TOQWzULzYBOwL5lrqhyoxKDkXO1Fzffm+hS4SRxgx
mj7cvBhUM6okdeTYH+fp7HtKQsr+y2/yPRi8nCtTWHpLHSFeTuBoI8te7GS7
jUTIkIxG1dO6gW2M2b6P+K7UEE0pJOX/pEPDSeZTXBODvu3g/RwqjpJsRs9K
LxNiW62M/1sHOldlSIiRgUDyz6XBEugNoGP91MvRcZBcT6Ez/cDZpAOz5S6n
u/ydoBVbnR0qlYAzmEGLXuwqyfewAg2kU+AQd+ZA1tYPu/Z0KGcAbXHmgOo3
BH0ALMwUNDXPnlit/2lYRwSbgD/UeVpsnm25tK1qz59uMllwrat9Soja2GKS
Bef7g/xnALj5VBi4lw/BPJ860H7KFNTVwIJ4lkj6POM9+2SIC826DDRgzelA
FZBuNINu0ACMg+y5G7dkMgNLWWfGgKNQ7R0jRVQ0dKg7rPlClz66S+RT7xGc
NebYXUW0bPh3Np/MgTsGf5NttRdEmhAQpP/bOygsvXOqc6qnKILVxxcCvbtU
BfErswoh6PFiRKcpo3+MsaDdix503a3W90+KP2BwJ2SyTtyYCKyWY40HFBh0
c23l8DOzu3mi/cP2IMt06ewI/LIliZ0XD90voZvBfAQoEC2csE8niemly/c3
5p4sYIP5RrnrZleVOLjSVi2nGTtFaQpK94gXnFg1KogiLtu4TuKrnWCyNEw6
AIVd0yq5VK5cKGIkgT3er4ZYvhrc0Urfn/QKOkWMZS9AxOUqUx0US7Xc0fHz
gmm0otI+apRELm02ldv8z4SeGQEI8mR3dfCRJJhm+x/rzb2R7kgXU1YqXPUI
mH3LPBTe9x55TSY6yi17FMSoYXnpIuFVr4G4kDKThWgwGjfp8Bv5TLWOog8r
AjIlgNLp72ms+5O+Al4YzIcVHc/FAZKc6FA7BtXi5Fr0yFDFHMVWUlkPd8o0
8EaYX+3jBWZn/YxWxNrqmRhmPnmlDi34i8MYe795fP4SGIDbkPftu785qmq+
lRY0Uxavu9RGwfGdrf7KsJuryIvutLGzKbrheN2Qb2uwoepP2bE5Tjl7/J+1
8b0UpwBmphAw/jiRLiq1k4CAd6CAgxNjer2icq9Z97aUv3EAZ8ifaxHpHg+2
STvWlCO4spRblMcXt54R+WR/km8nh/4/KAT4NaU/i8Hq/CGt+fkoN+eKxnf7
2nzfowQUmFEMiqyoTSwB7Utg0bNdp+H0EOPp2nr0rerOvXT5pfy3yffHoEEC
LhVPXouc0znzEYG3fbo2MgbAAc7LANcAfGRl7zUnq4VXuJs7sbEnkb8BhqL6
NCIn2iIcHpz8atjaf5gQwoNg0kjW1OP83CPPF62tixt4qBssicvHIt6KDDO9
zjlmlSw5J81eY81Uat8ChUfiNE8B1ZsSXOXJIZVgGTcH8aj9zd7OOhT0iIBh
C3WjIFSpLNbjark3ALwvp53aT4ffPW3b/BRcoCZ/OoIzrYJOrlT38SrlrQLw
GbwMBJQPMSemI3IgYTcbTeJrn73NT7VaHbHLLkh/8/+VvbODDcfLrD1pdFRh
uyxoEhG45hUR3//q58v/n6yFHJ9kL/LVv8CJQ6psyr4nYqv00RH758uTO655
yQHMZI2xJ1+QVpThF1UQ472FZT8eYg1XopTuUmCwmahmB7RhTo0l5bwPWfxC
VBknBiYq70Eg3H8icHG/hz5aks4g/cq5CgboCq274L8ymmIS9xOYn8Wfey/Z
CKa7fQy8/Ze6ylOJGbaEO+OGSJGj1HNujWFMtpimBXRXLlJYkxy3aVQa+hAk
Psh516Sr4/zNDK13dfi+16X/a26CFxk8qp4L4Tn/FWtQaIJmWmOrxS0ifI2b
jknc8svHrP+W9d3Dl5AO0oRG2C56VWCyQiwm/obcFH5SzbJRVl5lWU1BDiNV
ZouKk7Zwwrnn7QQ8myziOfJaQCvJdo6QM4Hv4d70VjdnZ0KFryXECn94xvP4
mxcY37We9fbralzBrlJb4vkZPlKZBtKo+Wdsh0opcprde0Ga14J0BFv7F8uV
R3w7UxyOugySHfRb4A8UzkD9UAUucXXceXe3PRak8EnMay3SdV+yRKnWe1sh
8D19s4Ykl2cM1MZd0p/87Zh54SYcWelVuzXFb9t/owMuQfGc789kZmeHR/rl
Y0VlmfEV/LtA8J9/Tr/VLIdphuX8mBsczhV4e/kk+uBkpIyNPK0A0rqaJs8r
NaNb2JhfkasjRdcZxXdIi3aejUHF1z4Rhw6KfMp3vjdSoLzyYyGz98okaCzh
0SXImLrk82q9Ww8VcJTIckfF/LetkBei4noxia+Ao4wj8BHx4WCJGHi8Fz8F
VC40X3Lnhsn0prqZuQEiH0AYRSWobJpG6zHgirXWHAHDFy7J96gg9liJFoQg
kxyrzcjgGzL0GqVjW3zD6YUZCq+Dh9PM0kYYxOSHODUKB5Vbn9DtNS/2At5C
QQRpGnbT+5ofZACKJDld3HQYnvtwI3ty1xpyf3xhvUicslgyyzWIvi3CmEMj
RBR07wdZdM/PyNe6NoPHntIO4tWhMjTOApQ95WahkomyEz2ZF6OEcOoksyi6
CzBd2mWlNIfL7a6odgSQ23cQ4wUse2sbGJDO/CLR8sTmaeyAFybloZvOgKoE
6Q5aN743nTSsmwtdwsLhDFw/HrqtOhF2iJwGxoCOVgm2pDGiilwDgHyYJwoC
S391Oike6uUr0jXd+dkwo4cWdKKPRes95P0cxJgznZtl2aJPNURZHm+ZRzaf
v3m87P73r93qvK0GotkZ+z5SyweRplWtpz6Tpb1ppMRqxqrdtF5fcjFtIb0v
SJp2r3e8FRKe4pLcdpiFs7ExvykmBZbFGKquWgV4MNzMKVpbpKxvVkOpkdcA
0O7dozBYZPcTa4q4shpHuz9iR2xSHrhY5CU1dN2juzT9XrwSrhAHmsKZymLM
/Y0T6NO4KXL8hgl5fOvBifGCywuMvzEApMr0EZ1b5fwc3HWzahSVXdtD82dn
V4nnVgSfekLc5YSGEomIwJmndGLZEgJvz0ziEhcJdd3wVPlRUXE+fWZLzz5y
509brV9u+KhJe/I5/hEEdR6puiF3rLb3e4fXkWKSeJ9X34HIOPY600OL+c7Q
V9spa4f0HmAfkbHICfjH8gQdIa9KSvwG27FkrE53uRmHsePRRssHNmwRnjBP
yghIvIn6WRbehNx0+DO1x4Db8SFm51WuGJzTpzu+SDyjPSQ6CSKh2B6TkoEn
YFFGG4JZU4QIZRYGabqkdVZPN3Xi9f8RDX4QnVi/t4lcyg4SCXe/D2InXeFM
jWBkZiVM84F0V/AN2UI66DwTeELF6lnv6Obz1uJqr7V5uRMBoPCeJjjl9dI5
vybgo6pJ78NHsWmVY6jBKPLR22zmYFGwgJQP8hX6hf/FmDDg2Qcc7StmAFJj
nEP04+IvoumHXzjOAL3lDsl4zwWJ3YIMEy8/LY2wctAy/hCc3IhWXzmWdG1B
1e2wOjz1oPt/VaNZLA+dH5KZsLq01Bcrl5zzyITy59WSZps5I4LWvYMc7n4w
fJ2pyTcDvIy2ZZ2KRhFl6092HrvXYvr+f1Opm7M4mWdds6eStwqkZ9/wjORn
H/DEwKMwEqgN7naGuTl8/1mlDCfoq8rVcZ9aokjTu1hILr19FZCFF6VG1Qjw
iPNxyBvU7Xr1vfQw4aPtOi905kWqbDFRDjcjL8ANuC414w5oBjWRautPM9L0
EbbMG1VN7tHwD7VkQyMKOEX8SLknwr+rKBxkYGHsb3PPli6BRnExxsUjqeRN
RIp+r6rRRiV27GR28EO/dPjNtuRgXgoqfbE3tlkANDzZOPq14RRpBitrYCu0
DJFsx2PNR9Svh3YoPui3Px9Xkgw6GbqzcoDPijgJk7BuTSJLrooStx0uvUSV
YTfDfvNnm7ENn0mVhBaUU0uoerkr3muloG9K0UF2KWLYxrtGHCGAnUzrB/GC
bzPqnbRPdSUrxsH7Ap5W34ZEDP4kb0f/VIYGzUOVX37TQLpM5OmC7gIMUo2c
nhxk9hp3uAiNlCFgQn6opaHYLm2SeCVdN4/opttSO07zJPb7q+FQs96CninA
k8BxI1kpdfwAoG+8PwMqoaBciRMRyKLcT9PKnBIKqCvOQ4WHM371ZZrsbk8l
8kOx8/qd33+WY40iNBetwa9NP82kaTd1FHdQg+3K5M3WqXEhI47zvcvfYGCs
3YjcF8olpjvPjIlGyU5UP9DLog+2ZxoyG4749lAZw4NoMF2lCxZ6hjT6VFEL
r7tSN6c2twN3oF6o4kcOxgPPiRaou7ShNPyGLVMLkenvUmpNtyWiE2ebImxV
3qEa7iqNqnW9lOB9/bdf4Bmbz1Yc/vS273skgGElFmVQtCSBZvFyZDysFkrK
VXxGJJpsusll3WIpIQo8LHXWPTLNekIbAEVfnwqsqI9EpFCuwXdiioAFzP6S
w6fR5PmXMyHskqg+5FYPiU76yyLH2XT+JFaJhnoWASci7Xthm1GQ0tTnkPHg
M6r6iJ3GJ81OiI7v8XQKHrAzlmv76lA9M3vi0hu8erDp4MuhYeGKfQrAtqNR
l4mJUAiisXRvlAG0+HaKRrBkyZknC+tNtZJoOLuP8qRbl2D9xEOKfegGQ6UV
qqyDxXHohBFjsKm4kLEw1jYUPy9LpXvmrwOmqNaVoP2DMBBZf4rU7LXEznr4
gN6mR6uDMIb6iKnb+MrUI6WgAW0F+GaWjlqdV361bXlbiynyiT96fLzX47Ol
w5aPvp5AuPXipWHq2kT6vUCxC5fPDyLTigMGnDit9JBNUKSIMWY7LvMJw9dF
RbzDUu0HitONyZ5i38yt0ZA7Bhhh7H+TcP6VhIRxSnw2o86ZSU3+sR2TSUu7
5DBY/PYQLuvMrmUcF5v6r9+YFE0zGFnfMENcSS+YjUbtExckohRVzQpJR7WI
UpWMWKjjZOwOXSrgUR+H4eAgJjaquSoJDLw7SWqgCPYvHp91dQ0xiN+Phl9g
GClqJ1s6zcivadRU1h545Z5lzuUoJ4a5NPWVrnHAduEsXqePpbpLX8oh/K5D
BBzSThC22W0qzJjXs+mmuANfcJ1chyl/C2ij+O0NBHvSPkV/jtE2oFbSlhQ6
yMABwYxzJAN9ZebC6a0VPiEnjofPf/uPLcFJ4uhADr42CWu96Mx51DvRSf/t
wj2rcTVlWXn3xSv7xaRlUPz4KszrWz0b0BoMz25rH2KeulbSz5EYhgZL+WkR
RVdiSC+59RBE30HS5nTmlGRftBtXLpMR1puf46OLpPevG17kU8+Z9/XgW0cw
mF1XuOk5d3kY2rtBH1wjy5bQnYEj7bJnMViFmfY1nxqslnnPOLjAlb4HivgN
2oMkTxUUsXumV5rl4H1GRvw2FuGU++80HIbt7soT79g2eCmnNX4lEqe0wWop
V/dOm9Ea2/1LZkL7LhrJ2DPYiA0fi/juTPFyJzQFxf5hvLYpfwsrXXyP+LU0
QntciAxsduPVL6VsPzIOpVFhquesV/+P3smUsg9bFPhfhN+75vSL3at0fIcb
vmcJjt5z2bMV66UzmADugRoGfXmcyMzR1jSdvAa2+9xWm1TKdjBTu/uoZ5Kr
8FHPLHZOwE1iWERoEjAtpvWBQuFKscMJ4i6WyMEquPqxlVTX0Uk1pvKNJR0H
28yxyasusZvSKmZ42hGqERnJ/kjTtO3aJoAeTrrOesaegmi6MmxYIX9HFojv
ncFM091sMFsNbqtY9jdK0r6AjvGrfK0DOOve+mLQSh+DHUW2XvqwBUl8x1n9
ys5nvYVn54iZTJvpiCBaEuefETxc2HTcIi7Nnt2/jz8kU5ZY40WVskX15kcr
Y9JFTTk8FPLjZISIBjcgJjwesTAf2or9k9SENa8kSCNQfb4qwOnSa1G4UhWC
WMPlrfGEk/WmtDi3laI7hgFUn48ENIJTUWXaIS3YB6RxlfDmqis5DbuI7iwK
yhYSTiy8P2Ar6GVfnu2qeuz4bfHq/+d++WcDL8SRU7EwEXJRCB2h1V7c11S6
vtyprxQpYt/22aeguPe1iBDHI3sRJn88ry0x7+2MVs3Iucf0DsqKiTxMd1iI
SNWwFpEjKe2kl25tRNuq0uvHiZ97JY8VZvvNMZFBEqNKGjjq4m0i6LHikSRy
DCUke2rdLut9RdQnLBRLc0nLY1Bbe9NPUVIRyLo0uZbniP4IwEGBDsfnQ2wY
KTFIawDWXZWLxXIH6nydetVrNxCl99iUvSm0b8dUSkvVQ/yLhzDrepU2Ee13
ZaXREXLp7TRg3oZoLzBaqDPoJg81pzmUnFz3ly5z+BQ6xgI0x0A3/fkHgCiM
ZXeAnhlzpk6TAdB7FBH2sGa5u3FmCY6Gn6Pr/EOcgGhwvGNmqIK7p0ad37kL
qlFBphs3dYhuxstIbzYJNnWvcFLLvfM+7Iqmf8t/ePi+blvfuuSE4aaDVhFV
7psCIkJzGOrw4VklC90ANOjwuSmNb3upJpH67S0+hg2Oscn3FVol0n/Ze4xJ
Re9Zx3EO+5eqjiuCgn51ymkz+3kCKmXPqTnmyfKkPi8XOMMnY9Uo5TDK4WCQ
TeU4K41hwaiodHOOzMVSPsnXeHcC7aX5cmB3JQJ1ohnXY8cEnzH0GyC03k51
X8sFystEfweLBmxghHEyvBe8WibYeeE2eX8wRfFOkaol3S4SkvcmPPoJP91O
McC8tWTSix13SCdoC61YsbWxhkDqOaZpmqiaRJZDw/neOr1Ao1xZR/gaK0Mg
OFcF3Pb8r6dKNQu/ZwkmA28y0lrjIGDywtID7dlI1vJqKGUkziP0GEJH4zxR
yamjZaqPAyZKQa5q6kpewKeGnNY4jyFfwQJcIBiW5B648+WhtQAhC37BkizT
0hg/eHze9ziNIQXNpt5rsjqp1YSzrIy5qNqZYnr4NlYnzhKALLNF6olRcBl5
mWqpFzBYzBEGHWJvUzoELseOsTR7gO+jlG4U4zf5Sxs4UQJSxt38HOws6pOL
CfRXGRASpLvUrnGfzV4rjB3Q08V4y9dhbP5NCkByVdD5kjKlwIL07vcdooso
fWdmOV0wdk3VT/7J7pVueD7ryow0w6Z2jf3xnNA9bonpOR5FOtUV1uYJDryh
fMjMgImSSpvgbP49ak9njFUdntOV6UoJqx3l9xUnyg+c7j0uySadIOQm+vj8
w6T3FzZw7G/fUutVP15NH8yXyMC3E2HVpHc7PZYja9xJrpJSqcQlks936PfP
NFOGV3TZ1IWs/PAcrHhXc7leCBBCTM7m5mYggUmiYmx4UiLWb2c6CBpN60by
Iwu6ucyOGgJMdRjzq6zb9V3WI+hkpkOvmCWEsSWofpfXE15zSygzq3XDBJKz
yvXEKRivsSD7XT0Xk/MUvi6ZYB14JD6eZafnyuMv4qHd/3JPmW23R6XdJdXy
VSoNNi2UwGa+1s9HGswuRxxzxfLCg/EBtlh2AAwNQmMGDUiZT+a+fBRmevsk
6jbMcu26JRjPy32WgkpeWm9z4Pf9Kc32odiX53yUl9A0WZQ75dKF5ZqGJtzY
beVEx5bAdvEc5mztLWOzsK/xA6FS7PaQr4pZvjjEnKCCpHvHV2DshzTp3MJ5
1QPONmH/v+lgVXMss1VtjBTsoJDCORhIsTPQbBA4hrATlj5mHNdc/HLfC77d
1jzbrQ1jSMzEwMTKeNlS89+w4ZvedBh0IvhdWz2sge49XKN7WLjdiVPTtenT
agFuWN7PWd82Ju9RlDNf96uNyOocpH1hylTrph4wRhyYVcgM8sG37V9Ut94W
7retG7TAGK4lJEc1rSb8F/RQOOVMVp9AmFuCuf2uFMx5rMmLZ4zX+f/VkMfg
8xTXvdy0vHBJQByzN7J1wKWiXP4pFW1phRlon1crR48f2FEkDDlK6gTmW767
jWcNx1zdDJAOojhbNumqlRamC0e2ek/Yp1634HWJpRWb29ggy34tcmVeQqZx
uEj3mwi06zXCoF/dihQOX1utrgaqBsP8N2dJHutRmuqAAORJgNzjr6JvL2j2
QOUkH/0c0nUmKS90Gz8po7yk4i74C6lPp0BYqYj1Zcm9Ys+dlk4EJ5jGY3ai
H0ssDK1JRj9zc1egE/iTXndovcl9paTzYXK89lW1b5yQDO+gubnm8F2UVHk3
/0sdNuN+kGGe8rnsisF0poSYXAV1oh8BeS8aF8NOJOH1h6jKblzwHmIgTECs
PUXDv2pHOWrW0FQl+YqRKp6iD7D5gZKGHyQEmKOis/ZoxGNxsI8+/MPOBpAj
EW1pMUTOiKPPdMCnBg0PZeuyk8FQ3EVvVgXYXlxvDn5ba0g8L+/wes/Pq+Jt
DblvLhI1JLZBnsf5Q0w15KlQitg2EpvKeqzUJ8BSRo9OlKePj4gtkPkR9bhH
TETD2sV0VpBquMZGbVWoYKALqEK7rHSxLmE3Tke7vJrPTzT8Oj/+TrjCtrwU
PQd6rKFNpJ8F6Um10WEb27v/qc0H13b+nqLi3tei9CZ+Vyx7iZLzPPdXWCmU
E3P7JhGJ+Dqn3uCzj5KLnjFsdnyaiT08gjt9JSto2vsxg/YY17BkEYC8QeNk
+fICic3kr9Vwa8Z8/XXtB+ZYcbe8IB9krk2Tspjpa9QYGXsPOouAp1DGKWIw
9ropz96Zac2J1rXyFCR+3cjQut90H4bTMkP0yx+DCNlFwGD+gmiEDQSwl1J3
D1T2aYxTl1J9A/1BxH9ebEV5H5WwVMbcxYwFKEMNozbMkgAR4oXqigeq1/4F
lwTzNTem9Xl6E9VlU50fJBNMl2W4o1HJ2Vkv2m4+yB3aoGtj6Ntmn5vsbi49
S/E/QmScf/DhkMAgBYAZX1shDANE7OeiVf4LqinQyWqoiRyqYt2KS7M12BTL
a2joJY3n5wuUT/k6heH92TCsS+JkXqsZ1s7l94xvlVNjeHxj0ZYjSpoWCggT
CP8bJA6j5SAw5xTck+qrx3GLJwxRw05MyBv9xLS8K83cqDjqjiln6U/04Ii1
BMYrAF9xahMHWWc8fTH98kEKhikOKpjQTIYY8/POGoEThTU0Ya3RgNS4RMPo
aHiHYxp9373MFeL5LkZzRkRHAn3Z+05LiYNZhalaIzFGpR5Jsq8BXoW7Brsx
PbhboJam8nmbP9pjcz2eznaKLE1c53il5kgFWv9oX7epfSG0nC2B2CSQTQFY
LknauKPWJjK5G8OJwVM3B7rxccgBlorGwTnUziGOHo+MxX/rrC9uG8bDb0f6
z+Sc1WTQK6avfftzbkaFAqFzdQegzyprIfJ7T1NCQOr7qNZbZbCrI16CmZKT
dl4+KaMRaIgRBOPQifNFysRs5vty5GBi9xuLLvCPD1GrvZUzt/VNFpRJeswD
ILxE5fXDd5lLuJ+IHtoGP6mpUUuv9sTck2xodaVNW6a7gkcur/AtHXnPohPz
D81qN3UI6GYN/elusbHJZnV7EHTh6d4Iyrwbr1gTcuRR9gqavq/yNkSXlOdz
ZLcMAKN/OILXiFrs82n/LHbu8RsIZJTRVCIYeJSJL1a3v+3KCtZ6vUZURXy2
zlLuDdV/PdhvdOgHkQ6+3sZYW+Wb/2psl2+L3E4+nsm2D1RfQptsMUudIlTG
UAoLmCxrMOTcg2jaNuNmymDgSFCUPv7yDeEV6KcoNnitstMgpeHPtCCv0KxV
PJ6Fszq9OCKc7QaMh/EFWEQuMYn8gNiHhHn+iC9ug/toxiZ8uZ5comUdo9eA
xRJugEwNb24SnCuJ+a/ezfLwMXZRX5/qi3cvpXZ1Lt67iGFfON+bXtC/sj4/
gCVG6qeqDYC7t/Py1oL9qnCB8eiRNwDGfasXvs1chxpC8q0kGL3N9MN6WVQZ
el2buUPTAAE8i7vX/nxzqruNg+mDH8iVa+AxwCb3alqFTOmRGoW3/oK4Y9Yb
CaCiPbvmYOJKuwAfVogXeOyTF9xCMpRI8G2wKw4/2EIsxmII1KmxSnTVqagn
mEvwOP6tNRPqs5RpHNC+bYOiukAQO+WzcEiuZWsbhQZqYnPHK+wBVnuGHmTf
z/x/Sz1Kc2KVkI+cucDP/RPDyNJTdta6xFoiF30oMkqzuRu6FOtioAva9AGD
5ROiDuECxMNs5ZR0p0VmQHp6zAKDFdVHRvy9pae95mTAHJDMw+0/A6OOYKCj
WtBr/c8tUaBW7yDc3e0jQX9w9itIK4so3zmxDHPm9LNMUf1q5ChrI7D9vwBQ
hPer6mPqAkKTgUPE0lE5VrGRXx1Ce2muLeIyALHUtgU8q/1bWPZAHXFRhX7Z
nUwjXpD1JKIKppVRLc683sxD5/ortLCYE0qFP0fjdA5IvEhQTazcjkYoPcHV
32hxPlPWo3+8CmTwH8sBpdfzQupL+IQQBBdeOyqYAJshscRGujNQiaXGsu43
2ue8IZAbZjY4qwZtfj82FHYwJGeODzxiFXpYUCIELTv7WHGkGa68NlAnWyAP
PKkJrOaS1ALCaZgMNPzHO7VBzqh/Hnkxc6rsnxRH98LCdXy1zL2rJnbO1NCj
mydBWtnhNnUDygZhzUQ8QeeEV58xpsXZUjwizNRydSanazq2ejJvFSJRrROr
h2kdjmFdLlmFzs8S09hGiXXtgXNMAn5/pCuYE1LmeauRtcsM+TE7y2WwLsy4
plxOhIXEGkYGTkcOI4tkYFT0h7Edpfy9VBLjbyQQiYFadhTUrkOvPc3muCRt
+Ps1EjPs+TqklUxfUEv4bVTgCHQ1qy6CW/429rpTs1XN7ZfIglHvjmgnD9uX
tU7t1h/Sjqc8pdsaDRRMnCmaavuyOSrndB5sBwEoClWpYo/houJd3ZwyMuPQ
lvWXP47H9oywEKEbu5y7EEf/C9dar+m8A3TnYKJ/qSRqz40xN8NdlycO9IpO
ZpZdi16WnioxmTGvEEnxJNJjFXY5L56JTE8d0BIce4tRdOIb2FQDszZtiYpc
8ASUm9Eo+yM1mSY0YQ0h282p5uTLEXPhu9zlFqXif2phBMsvHCn72f+fe+7w
yD41vb01FxgEOSnD3JW0d0c4IXTbZwYi9qum6G9cHd3E9i8SeO5EpRJIzA68
2tT496Y5wjko3on5U9eeUUcPtMiuLYRZ9h4fr98joOcC8mNNOje07U18KG4a
LxZJjXHfizNOup3GWQe4YUhtWHr21xiLN6FMlqPAW+AXHG0uNTy8suJwV2UH
FiFllDs8D+28EeodXHznvvY8kU3znFKcLVemGqkifFOqpFh9gjUXQt+S5/5j
Reui4u7sgXa03cbUySVWPDnhyI9lTzkwHHW5KmwMke8QZ+sUEg08bGlDh49v
BiaAgg6x8L1tkdURuck6r1sOl4BQKGfWOBPk4Bk6BITNWbR5NElXXOFkpIzK
J3kYsuCH2RKz34Ttei8Of+JUViCwGpRl5D5w/6PDKCMxhxC8ajTpZS8RTYsY
F+0v0VGpqm/8kf1YFlGFgCw9s685dc0mHh2jpweNkPlMBZgpIoJZDyqehDpP
cmqv+q/x9JPEiGrWMFQqGJWs/MN2OIZCCqkLX+/lKeT0CudIaDJKXSl1/8JM
pNCjuDz70q+dhDUbxi4egEJWC2723ui4Ru+FyECntl3s5PkG/3QeX5qt6m3u
opR8n/j2I9Ihhi8FGEwDM1EGy0uuyicuitn+3dtzOlz3WpVSCZJqbNTM7C/K
rG1nfT8zWjMGcqoUyfzqEtykNdWXRGvkGbjwYtWpVMhzCNPAEQICQRfDbv3H
TKE18qHKe/2VIgTd3zmI0quR2505TLYLgy9IptDkypBVOjyFzutdQoyCGmy2
xm46Rf4zry7nos0aMoCRMsA9lQx77VRtpx0J4KwZrAnyxkHdPeR5K5PW2PUQ
B3SChBw1RhgLb3hI985zZXVzyc7iQO31Pb7OvjZkUu/mLyrggmQcQtQM6lAH
PwABK+9u3obDdoxvdnW/whvpsHH8IsKQ22SDERQKreW5Lwp8aVFNU+cR00xK
YUdKfV4xEPjRYr8SS6U8VobZDWNhnXiMwbPI2i2o4F43FeX8XlGRdg9ZAtIm
rbDITdax78J9RNx+Ku6lasvzH2R8vMNH/hKMuaufqDSV5Jza2+hkB4Ps/G1W
5xXvIa1gnTN4qaFbQVRvf89HjW2oWe8FQMPZT3pOg/PxNpC9wPmTNTesB3rr
MU8YieONylvYz7aJeOKMPiXjGcbqtmaVY163HJnNMkNFITo3L2svnFvSrY2Q
WNAOUOOndbVDOqRYrq4n2G3eTEPnKrocejLgYIVkAgBSzgd+G1uMWus0QqDN
1yyOxcpI7hnCbnqisIQl6NZFf27Gv6kDQho+qsQsKKGCeYz4sR8SwWeTDKZi
2wKJAT0YPMkdfFwhgHlyaW1omEo2YzkKZ0cGoqGhRAwmSRlBg1VpkRzOcQw5
yAU9ZphHujjXnrxdLLW8tPAMeffiHc9Yvvao6gi1jzJH/RnlbfmSQhokLKbr
+LIMzKbEipxFJGasbgL0gkM4l+FJURBtzEKtebySViOFcIrI3UAQVbG6XbFQ
lFys2Z1e/oSX9hRuBg+NZOz7Bs4Tj1Rwts0uEReHH8KGNmAvUsrQ2AuDiuzr
+hAmfQjWJ6BlIjisMiW4AoH6jA44CkScuJ4lQbg97s0DqNrwafbzywLfFKmx
hQh72uVzyQhTA5KGPs93hRl5o2ZmehxikqBK8/IECqrUKfKnDa1YBeDsrGF8
EqOOdZ1xNWSdcDYdWtFvX4sIjyXjvKdhZHFbmETOvrrMJG+zOz+zLSqbOaCp
+l1af7pgAdjDn5vufiwobuHj0u6iLmCsQldC1mqUWT5IA9YL0lTMgFJqBmuO
/Ge2fvkM5oIcgeSUAqTJzPwIb+bJShEB4Iv5i6fjZaDKkThqTj6yJxO5DaPE
RpfndMZ4mOA1p0t5jGtDwMqoctiM14iloO3UY6x/48RuNcrFCBI+RaLZC6zJ
jWOwjTS+iJoDXzGP/Nrd1kOPIaMkBSxudfs9RRL+Hp/hMueL19u5zoQynQui
0qUKJcGsP/EI4UFzncaqD/gs9w4EbaxZlpyp+VAqzRvQakeBpXfrD00dEnK/
7oT2lsnr++sqXfUIYpszm0cF5nsEKttwdXWPPHQ4gUZ4Pi2YCJayfceqBGNV
LU1TWQQgg3gZepaaGRGp0KD52pf66GJOR3sYTUvLt3BUEtR6WlzYOo9jwQI0
BfOWd7qcZKhVNhuWTeq9DB60xbZpwQFFjY2oYghK2KHplot4rXK7O2+C9z0u
YQqYGZu8LhQlSQFeNW15m0LaMdkeUlPtGMNHbhjqHYf2gbjzUwxmX/TcGQ4I
OtNzW7HKr9DjKlX8bNs6oE20Hv9YUBgmvpxg0u6xII8da37OUpO1ftiDUzlH
TO+DAV7AVOm3qBl/Kh30TVsIi2pZBGq5KEbly0AWQ5sARd0Dv6s/OvV+hB43
vJYF0JnCL+vB36exRZojwugGRGcDV4ZF4uJ9kai6pEXnOIL6lnJsMuuxpnGq
Ne464nuV1VHB9uFdg/NJ34/fH4C160hWc9WZ1f6vRuj3hnFtaDTHdAI+FkqY
ZiZ9Qvo/X8cLs+jjm4QE5gFm5cOd8v77OJKY+4tQ9XHCp3dODpoMLM3JFSaS
8ESsVtvRBSGrgbkX694rYx55RZFq33fIzk2t1Fybjl7TrtXvSeK56gYNvP50
2ovmBA1SbC2rmUPihDVaO0QJSJ8MStHMkPUwiUXEym6YW0jyhOa4pNVd3gYV
fKUs0C71y8aduj7i+bCMuuGzJr/dEgdlK246czZlqpXp2xvGgeCfwzNViAXk
qtfWeoJrz5bF1lj13KzisrrtIXGaw5oiSJtxzRSGGLEa+26ZEPtVx5EYcarp
DIvTbTghEwFPvJX50/Cac5RQA9P3zvZ6U7KW/SJ/RJvn557tUvWOmL/apuE3
CkZFqRvFJr4LXyAei5AfILSk7SdcKWJFu2gmuFxxtqmveJddmhFcil3DbptU
P629xeW8KGEK74QIaqW1KGRrsTRjr94P1V/h3XCQZCI0s5lXXKELBmwpizi0
KOC7lJ1x1dPabL4m8KVdhY7a3cZnKc2Mm5nd5M25MYZkZLUL8ahFOQLnPFQB
xm9HWkm1mk6/0tkwMHvTa6xIM4sfAt3VkFi/f6n0GZL/sK0tgABqK7K9SR0x
VyOMF70EomQiETt/2WSzQSVJzVtns52fGrmyipY+n2nLS3ahMIdwDfPS9WBv
Hknv2hTLZRnKtcO4gshgo35WVIMfxHbmms4U9B0BY77oSOW8Wh6OXqVjQjEk
nG9pLczOeRwScjYxjEswUBwHxjP8Ipu9sSYr6ESGQa9qq0Y37bSJiqZv/8SV
rt/1fcQbwzpRTtK0WJ/Wwe1mFO2uo2Sc4Fw3Tzw7fcYMer2wAAXSCy26RSky
l3BEfErQS6o+p9r53G6vcfS9YDxFXvBtewrpirZB13TcoQslMMiy60R8TzLu
dVU8W40Kcg7KUUS5a0fR0bUZZW6ydGlNAd/fsJckTUEb+lcCswFSU+46MMli
QCif7PencAduB39q/HM9FE2hxsT9yo7iZo/+8ZjwjIKfZxAnaWPJH+oTM9Dh
djak7O059nTnipenojAbkxGJXFKEH6xbtRsVHQyFSFPR+ckFH1mrBLrVb8Yt
NnvwrMKJIkO63fsjuKKCpIGzMT4OWVOkGV0AZz74aLUaPApyes98iUyGtMeu
+Pu8WAk0gel+UPQ8xcgiWYo2d/4UjRolCsmGQW1z6OkJDvNhpOFS4u0N+EQu
SJ1plgqKFkMXLR1jGWle80niCX43jbWDuwo5a5F+rviwHwmLmzKRZBSe67hJ
6LZhlimHNkQUGhjQlqDEdPdfQ41G7tH3+z1bQS26cojTj0GplDRbh38oqK3+
MnSOxWM/bGCJuD4hChb+C2XjOTVjw7yNVF0+Kt87V6CBkyyZBweFAixB5cJw
eEX9a2DEwD7/badekHM8CZ9oOfS2l0UKWU4AKuMW9JFY47k5dzQsQSZmNo2D
waBOqWvgasn6R7YrpCnUSVvAWAJ7nRaz1A/TZZ5SFlAwVGlCXo469mTtUeRM
DOrjaWvJ8kiDoATQThMx1TPn3b21dPfgwFEiwwBwlHMP//TM+O4L4pjwt+H5
M8aga/ZyvmgUdcVgol8zNiee8W+NQ0EnBosjxZQmgHJycW45yiXRircPjCsP
vD05hcodp6JQF5/1PD3wTo++uDinh9GJvdoiAflBA4gXS65jv+NVaqkcscP2
xDm6dMCHBp0yDqj/PxQs9axVB0n02kmGyrQC5rYeU/tbTWEIwrOH+dWVa55n
bw3Oy+0OYB4oITgSVc7oJ9a3vxTHdw514tA6uQirtWsUcFbSdrA49idtXu4A
2zN3ePQjCmzoKK11sNVySm87G602uH9rVjw/yr3DJ70Q5zSfzVSENweP1wba
KAQB4MLaI846rUrn91XB3X1nWuKz6U/rmsVMtVt+jyNrw3QwAsa2HbQ0Ik49
+0J6gB0huJeF52smjruur6FjVKvTdaj4DGbiOsBoLkSceD6qBu9zyC9OSMhY
BiYsF6z2IEz1Hl5+tbd7elk2wklhseytH+ym6A2F+ACKrr3nc5mm5g40QZOO
JjJR6btZFXHgO6tL7WdTmqmGbcriU/aTfBn0pJZG6wXcDtwuR4pQCzT9c59E
naHU+v8uPI1DCS0iYrcR0Bb6oZ595//ZxFdzogx0XguiV+QU81QZ9ZY9oROn
5OY25fW8gviFLJmqGB/THVFCA/DCLuolNFAPDC0QQRV28iXLcuZs2bexvOGa
Odz0nUyA2FNOne/uOAq16M6sqfzX3ytteLUrJN/Vv4/UzKLvwIQMYxAKqXKI
UIHp/FP1heCaK3vZLFw0iikyNe8AYfGj4lV3CQZBwqyR69cPkDs/vG2HPs7u
OQIYnEgPyKyQZy7FO4cwz7em58F+Y/nXXSct/nBYcIa4PuqUY4mcaZkZGMbq
phukcvFhYC96OK7waUSQtCwqzg9EbzD4O0RGLZzoXxMP6SSPvypiRxBgv5IU
NPatLHOdai3dg4wZk708bM5jrIFvX2gaMkCi4zznlFOppvyokM/I9eGyaKD7
im4GMA0D8nB7F98LbZYaIkm8R29qVkMDanUZoy4Z7th+0rrxQja/5K7tfmhK
R6kB6gb+yGvt0DkwXqwlNY2TNsIkhrI95fS8awUHovpWVZNNxxTCkoLaPg/K
Whfgor0iwo604q4Q7Qkdyl6zr1GYjaBxYwA9owWGqc/qxDxQA3+nmwhRkVBy
9y/s3BUSJVjKdjOeXobTEJnrQ7pxfThwfqF1eHLGkWckZD/eDgKO9Zu+SPqg
44eLeQTy54B1yCZUjNEdPilTUIWEBZ9DSI/4z/9yS9DHk+ijagD7cS2YiVtu
Ccg2A/HeR7/TZMlil12ZNztCtOu/20xugUIsLs/lC+8CBh1EG+Odi2GkciFN
CL+CuyM94MCbbWitIP7kgv6kClbNmHNLf6U4iW3UnWFO/bREpaMGQvWhaz9f
6U5knG0g6idgGcEtUMXMVZbFVvcsLahyot5VxhJRWu8B6aJwSURMvf5aJElg
96XyIJENNUJua5aplXDl4A1BONEXSjQ78SVrDVjocJqmA0G1jp2TJ7q8Ii/C
QxfsGAyj3shRoXOMuSUNkQepdGIUD16LQgT7RnbAKNl6Nx7pyu/YGUxKTlb5
ExtjGgP6zd1q4pcLIgzw9cUBBULEEM2pXGdHUD/xsWjTWlhG7ZeDyhwQgJ7i
jgJ+uFwkToYXkO7DHViUteLWCfQfwIeQDsYwk91dSmUtRFAfyHBc0tjhsjny
aeFLCwwxaaX/sXAkrnpJkmV+QJ1ie/MmUq7usGC8eT4OEo5XM5ZjZoaB9wie
TI2nh73ewJda46Nsafnv8ddJK2uI0ncy10IAt3ffNO10yoi4PiXvZondCeO1
NFZuLGWCAfCMOSY2PB+mNtVsgeAIxONsr2Csc/zgxooMCYP8y/dTk9c5f5tw
rYye3PksOezDo5Sodzue2xNMA4PdlNh2aU4E4JdkzOVlsDYqc4EbCQDa+ak/
IBke0F822NPCHf4vaBiliLcCiTCKsleFOy+xCW58leiXKBQQRhChrldWjjwu
o67wRtMCENg3cv8inCKp+snIWSAfpOqk1l4l/TyptwfZUv9KtsOkg1FWisNJ
IhMpb4m81cqFUZnilHmdA+b5Ngk+4scrrF2sdqRbYHwYOyXzBKWQMaHBV88q
y69L+Kjz/9S576qeXtfUmeggQMf1Sg06R9H/YDi+S+ebOpn0k0uyNDjK20ZX
gC+hC5rnnEQBRCSjYDDCNJw9GUY0fRIT3HWTHhb5t3UpYTCl4tFbEbYcUr/w
1/FyV18pxA5GbldUGK7bqigcbl6TkmNqdclNW3fCvOr+6exd2w32y8PQcqHz
4Vi5uUrRaAcOACZbBHq8tkjjzvT6BH/ggJBtYZROMLVyz2zxCUhE3cWR68Et
scx4zuCQLx6ad+cfWhYncWTzGbclsBCIYy+rjfg8HNI86cwKn7oNUn6aE2E/
pRIqwdvVBgCudgI/TF/GNQ33D6vMar214MTW74YdNl/xnOtOimD6elE0Q0W6
7gq0prT7dGglYl4Ov8YXPSmFe7Y96EPfz15go9Re64MdDQZnet1VvSR0M41o
v/yfZvp5jwp2xB2lVAtn1sM9Nz5xSfbsgXXJCiH3fLDGMuGjo3zi0Pe7U4JA
xslzNvQFoW1VPNRnli/xQ3NRHYg42vyPg//QOpJ1NtzY8gowfdtLBkO8Vk5Q
wPJ4COKvbH2Zj9R3faPBl3VCVWrOP9UjVM9XnWlQDfcbmzjD/3SBrsDqaNmS
QsCDghzT8urPnREskCFSf0vGeYyaw6tZR5xxJkQ27h3FSAij/B0rrNyVTIhi
VkPdPTvX4+9bZiGb/cHRAM1L++DbBFqS7QCnqHU3kostCqJkWE1jTRDKFzAz
QD82Vw/6bkhaIlPcCqiNGptBY+1pGWITC3ZNrsUqU3zFDUBNZmNUaVZ6DkPA
FtoRsdNzgHzmVUFpXQGMVcdnnSoMFWaP/TFwyhwyHdrfRIHLhNAuBEnnjTol
BOu8VKkzGC/u8wqVGLaw8sOTuDYetjsphuz72O7altB4f1Dl3egAQAPt7a7P
kC/yBRWKgrHb3ixKQVx84d2FmuVfZ4Fo+19vsExQjpEUHTgXSjkwDBZ2n2lC
pb/xfW8aPiDYr65XbhfuXWnw7Cf4t0Z77wGsQ38dW4szBpGqTDFzopPu1QbB
hP8R/dJ6CrnpofurCDAyy7Jd22uIm0+I56ORJNb3+6507nd03qjldP95oWOa
67fuc6uGDnkVHoVyyzjeFG1ma0nWnS19vn5JQEKo+vFg6o73UMXJHjdpRoJG
h2kdkl/wTrGl9nlJwiCW8nU15GerLOKNnNVw+38UTpJA1nkjowD9BnTJliYB
FydpRMo9rxYWLLReBP8MIIF+eZ1sxFBcntoc81uoTX9KI2icXtPTplnmwTPC
SAB6o1ugEKf2pOHQ3W1YbA1XRzZjt217Bv+t4l0m0Qk1tdCyxYCIHRlROQgg
5NDwvXwHhxSBNimmp+9eItieqEKkYP6qHdvYCWWjKRfaGzG89ErCr+kt28tS
0VAErnXIOl9wpXOY71KxOFvUeqkUn+AbS5swRX7nI9/rIqUYGUEczIsJ5MWD
+rNQlqVKHz2gRokahYWN4F44NaA/Dp0PFvb5WBbirAHtIVS3i/ME/9XN4SoD
CCwDXuwhG0TXGz0IhKXYnffJJSoqDXYzoV772e2aTmNjZZwhaIsirWZOPdVP
GS84k4THu4HfIw/oXeQ926AR+zfNiANnPurUk3e65xnc1VIEzqn6y99Eb9NA
Tj3rcMtA0cR1WhyNC7adwcK5ZPDeEaMLykNs8+3AwDt1WNl9EZaV67QD7r+T
hp9tZRO+5n1Jw0/b2M98kQGpEDw16gUXkkyl51EXxmh/aJkx0Mmz4eTPPGDb
lwPcVkfPWWRKD8Lx6o6Bov7hHlCuEnZ9A/deP0AqCcaSKg3E+WlrmDPeSA3V
gtHka0D8+fjETDQYpEzWjwMW6uzqjDUQdEwxeuake6hsUz7aG7ttu9nAxD56
pkcbFOquh823da53w1jfdudOihdtyUvJ8xLQgaXzlbEXlVL0dcLH8mtIeo+N
2kT9AkXianPsfZRqN6ijHLPB6lT1RgbPArDgVbbZ8LxOwtbgW8V8bgDKfmiO
+EZJ1Ph90UbRbd6iOFoTbIYu5gj6loDeg6eqLlTAsjYoSz0oymO01m42ilps
gXzlMgbuNBXGTMOVPpqkG5GKpwpWCghHWT2GFKjD1FuGWkyVu4rDN7TiP9gD
bTJoNPkInmIJNZcfM+wA/zd3mc33aTTQkxzVc2NCkbH7VUoWLLIDuS7MooEr
7qxKVO1dDfqDP4mzVUGWKnMmVLywb2fnIQkeiqLD7tXcIvkW506/V0FJAg9J
EZAH0OY68jvA2f9wANRiZYeOIh5j7Sf90AuAGUfW5346mWR5MpYcOZuOUPNA
PWM8UHKLgDDMOXqqe1HzYQy8QWpjeOAg0owCm1miK8FTJZj1o/t077rmrQlu
8uk+zqUvAUGSjuzNER4hFGbtIor5goHvMmosrLPhqOsHDWE/Anp1+oyKzhqa
NnMYJ3qilgp6IBPaG29ZS0TaHGBxyNnjGhG4soR+Ewvxq5OkEyMIMwy3rJQy
f+0ZTYblDt0StdOIsRC4NiytawgoDt9lOvBy13orEPxFbtBvbmP6+L9/r+GS
afsRAO4RiDHHAaApWyooSZUKaLdrH6kRI7xaZqiGIcTK4joXbmA5tf6jjqEu
sncV9b4mjfgtwLwHRKoHLONVmEjBddRkEvO1R2T7FQU5Kz7bZKI2zvsA9UF2
Dzx7Z3cWFdB4p8g+bJ87zCX2VnBXLmBXcoGmbzfzXeuT8NcPyIyu+1lYXGln
rE7iw8rgE3vpt9Hgl1qcWIZpcj5yFCHgJ/an8J1ndafnt7rdsfInJ9Lj+Cry
AghnfU/QPFv5olMgUGqP/wP41aQWeqOzAkFuvb7WbYtkOUo8/8nO2itYxnsk
a8EBGo0dUrKK7npFKGlPp4gH7U5n/bcHc9cOuyPRJA3q3XTMBze3VOv2guKh
8xZKElmquLk3jlzwy1Stp3Am5mQQ8qcli3pyW4bdYhUJhXiXEmaZrFEGjcEx
ggOjvzl1zYB9tfANlIMxMW7GJ9VYG0tUN7UCO8DjTwXkwgEBgT4oBnEG7HmI
VuXFLQWcNmB5ipJdZrZ4ZQAmYnaZvn5ZXMQN9v1X0pXgWawD/U2CbijXK3ob
UFPP+boWICGWQcqtH+SgFEX/8Gc536P9DuN+UrqecMv2L4PC2JJbuhHx0qjI
mQjbW6QvvT2P/VklTys9IR0PSn5XiYZBBlOD8zLEB1fVLCBn/T3tly2IdLRj
T7ELHijM0VB2lErTlGnb45xn9eSOKpGqtfWnolNBD2s8iVwsXLvp2LQKLO9G
xjrMRU1ZYty7gzkuVEVZP4KOUs6yiEVcdJ3E+Jgde4PlW/frBzaFu/yBDjg2
TW8/szcn3ukhzLR2YT58CYqRCg0XmbyIVk7CC9//q8dlGTbYRPFxp/kcG9wP
0Hot7UGdCiQsSAmsEdpkUEebiiqfh9cjraA8Fttcl20VfKe4svybeCPLJrHn
BfyhMe6W/dqJ2/gM5obhdl5lasbwDFeKBMz4IaetkUTM9EtwEYPgeemblpt0
v2JbfSA+zeLedPkVF9jGOFMiwpNJOsImYcOoRObtNf5Mq4XemiflK9dW0jQ9
B7MvT+AuXm8GCygo0MwnxKwlbPAZTPpn7KJZGEoygxDSyDqeyESia/1kDJ31
avElJz9ZgiMk73tnZPfAaqjiTT7Mh/SLnRYwAGp/EQuGvf1MtdtBzx4Qx4n5
fKwoCHLP3Ny4SLg4VptQoHFW01BeWV33dA/2bp+A7RZ5/vEg83mOTIbHbL6K
qTatC99egBXE6/J71Fn9zatBCsqQBTfd4vQLS2MdqbSfB2seERXjP+Kinpg2
FdeZLNo4jj9tY6vvhlvY3sJLGOOYA3veQWjlBq3x90QIbxAvUQ3OCSjSsyqt
Ei+cXgqS4RdyVWEsJ0fvC3Vth+RACn3a9grbo7IvPuQpTJW+vSucBlfOuKJo
vhz1tBTN5BznKn6fbHWL4nybCQomub5Y9iofSv7ybl+x1r/us9UZguX6zPvd
ZTmbdut7vmt2e9HTiBk2G6E2iun7ARNzQTk9a0NFK/gBzRgNdsMW3m+HawDN
odV3x+/cjrxPy5R3GvXSO5+JHgjzsYC7OBE/pO05DCzfFDVKQcAHDwMK6rB8
vEgAgAh0k5H/DgGDITT7nK1PUhPIgZpE6q7/xCZxtdfsl6F+ZNwUZ7ggCi0F
cAdjVoqwk9rR+U+5bewqu6MbEQC/Z+SXu/JV16qT8MS3q0ixbWUUNj6XnNh9
cnbBYyIg4Lp9J4tnpJH7S1/Y+okHETb9/VMO0YPPyd3gztMPgrDrvzlrXtAe
3Eo75PO65hnp2fILwXciGGvN6wtWsXKX6F8/t/wMYmVr5md3N6Gh/mD/WPn6
Er4dnG2d0/ok28oLdrQAHXvbWYNY1FtRqPoh4hup929rY+BNEJCD7doSqjEV
U6NaZfQ0KUVn+ERdvJBXnB1FWgJbEggpsFWoBLDAl/VzDAef4oAptxWwgHpV
UZirggWzOu9rzCLJIrRmvWvvzzBl6U34ixV3jYWGpjG3Wl57VOYWGLLNq8YT
24wD2VKong0zTM0khOr43kHJHME+FbZ1BIv+HXm9eVmHW2FAKpWuNPARutrM
yW32Ti9JV5nZ/kYxxegNFmwN75z04SghKr3XTYf5BbuAUIlkWTAE+3LIXZjB
4Uo2aBEWw8BzAVNF8HLgmarJndQVzZ2AgyvkHbOPJqv9VYNbdsRLepR8lJmd
ilyJ97f7hoaRQohdKOuxJb0m7W5jFwkGzqK6zxiZrEzMBYuxL1pyJlQct5jj
OtPoXqPq4U3TFnREEjdnXN7GBeT0Vy4e5NsFJMi/FvE8oXTfeEU7FYtgO0qD
mMDOGrWQOhiBNgbySkip6JStAHgCkIHlcO0mxNtBxZjYoOVRejTnVczXyQT3
H0JcwzHZAuKtXzxnGvFxL6BLop9dZp9mH2CJI+XjK/b9QtAmKDDFuSB5LJ4h
fE3fqqmOSsmq+zP1STYlxdPAHpphCAoJ9/LdEAW4GgQ1wacdwoQvE6d9NZTj
ONB3pkOkfKY5ggwhxMRzvVVwVdFyQZ2KwcuHK469PBe3h2CWIrBcz7sT24pK
vhqyiDHYvoI0rEHTtv+p2yuTyBts/8lW/8bjHjQTAldZrcLJes0etwq9wWBM
Ci1JJKDH41qCxldiwrryXNhSgDzm36aBQVC+AW9x2Ml1WLS+XRck6HhL48+T
1pZ5j+t+ROM93kVZYM297Vj6fZLDcJKWbGUCnoiV9XFt3zGoLunk/d6M7A07
2vuvgbyjbQD8/dGkgO4kE+eXOiECAEb85oF1KjuMesi08l4wf4G4sZqDj5Ar
HDxF4g3kAJ9h30JbbjSr1lnjiI3L7FXPLXfEmk+eCl/o+FLNjBn5AqdKV6XQ
bk1G6KP7HrXMzbdzpoerHUVb1HZsHAfOaD4wALbDjugtTNlAThz78MXTgHWX
w3Rtwli6PDPG3pXVKVReKBepBviO645OQGRU0FW+9hJ9xB5JquniMTjgUqpX
/zCPtNjNMNso4OyNyA3Mv1A2YDM/nbUl4P4WNGfeNFRz8+zeW7hbNyyOj/5v
em3T0j4nfOAYbAUmazwHARkClUyu4yzaIDinDHZamXOTwcdnAI/OIr/0Ve3s
yC/Sj+rM/3gNRzpa+tDEjezX3Xrub9cUDOJAooU4HjL0lN+AWMhU5OcSrUA5
NIm9vraKFZQ7Wr9I6kQR4nYqp0Ut3C4m/HsRS3J7gp37r0TclC2m/iZFfYI6
+PBCBPqGklRW90T+GMvHnDih9W78HtIARje9ppOi2Vc5qpWowHgvcfYCKkD5
5EVPH3sLl98rlaWVDRF+jAd595NcsZFV5X8jGsFjolKSDhzFx0MMVFi6iWli
YE5kNSpCvL+grBuNoXvWEtZr8nc/6fFP71KhPyJ89Qm3fS/GgjYzCOesY5Bw
F8H1qAbJ3jMwgG9G2bmPf0EoMy/JbWNeXVuFCKXueh5W9H74456K2yujUGct
M9q3b+DRPgsnWy/638Gf49wEX7vepUzA+xES026joK6vJOWnkZrz5VIuTPUQ
SKpWU/6Mz3Q6WaH4QhprvRRDDheZ2UoK/IQtwB5j6zAy63UgVz63wtTKVCqr
2PqqiuUzedAEeUQVOn0t2k1PD/ymNjYRFdo3FHtzinIJfx/E265/KtvVmwjq
0zTL5LSg1lu2hJGp4cu6z4JEfMKAZ6OurCw7NvGZ5dsk9/qmBt/uAbl3tWb5
OGtGw8sELlS6s+R5QN9hxOmiNxSHujpm/lhHKbxTV0y/suYmuY4NZB6I9kUx
/oRRZPuc3QD4p8Ufm412t6zgrXKJE+htSSV2Ik1ep//XJfZhD8v5R1DhVAfG
sOm8yP1EDlXIegxIu/yLeIDUxiZn8zWr4wlP3TXCrc/Y5kboi4aFXYd13Xhn
G2OAOu0bfcIoQXnPaa+37Usxg+11KpV5gfp2Teb2URPAYOJEj3U1AY0Vf3/o
ZYCBK1kITVrvmy1LEfipvBuMKA1o9besShHelPNdGYvC0pzNOi1SK3I0J2sp
TcDPEpG8cRWdboMLhqR4eXcGLX974hZh+JBRwlSCj+uPMG4H2mlXhgX5VvPv
n9dVlevSzm7Yzy6IzTzakq4H/gq1ckReIKRL3h5ZG42jm5/N/S6+Mzvcy52x
NC2XXQRQSM68XJf+rbrEoWD672M0PyO78CUj+o+asVGlmi2/faTVstmPFZv3
bk9nJZLbyGCYkr5yFZyhZJg1ZoAb5fRHZ0KltHTolFsPYfBH6HoFTqDJxK5b
D/u93Elee01JfdSBfIqZEmr//AdfTzDzrE5dp1mvrcCbZsR2GZh9mdcQBBay
e1UU3MGRlube0mrkGPwlzO79cDT+ExiVdCsuhS59WUulFvIlDH5fxoWGc/Bv
TvvI1Bqk7Q5/gi539UW4I8dDSwXOBYFC4KGTpcRzDwVDF5nQIPbiPkyPr5Vj
Rl+isBYXxqLSo+kl1QeCp+qgc4qvhxELplLe+xAiAKKg6Gv8iI2AKzKjyzl/
tdNbxg6anE5/znDfCp447hRc0Hx0ikMZpSQXOUsvvpofJoFB8pALu7JJRtQe
A5++lyCAvJ2G7Dtre5/i/E7fkdYvexEcv1Z+ck5VoCOtOo8ZO95FFLOtDpAv
H+S6yHyGni7QGr2JhGEAYhr6fwzebV2dBFLT7HtiqldPGYHEdXaf3r4KcDB1
1a/6HJ+Yj0MynKw6gMZNF+sJnf6Q4f4opzykouO334703mfB3mpYh3MwIoON
Jm/JlWU3yov5LpcNumFvJVWOX8QDf3oNjhEA3p58NE9R2oOuaLs+TA1wUw6+
IYC+1xfYrbTBSuejlHkHygN06SNCtV1fBQUG5fKKW89IhC54yrOkQulKiVQ0
fHXYTnmX2FoNlk9AEEKV7Llqeh/vS6RptnMNExWD23go4Slzcb7fiSJuuWqw
onLt9f0NYlMxhrj0T+O+gw8dUgN+aayKhP8EOPqQvZUppfXCe2lT+Pai6+ml
6O0sCpcCoGB3Gjogr/isI1Fgz2t8mCa2196AeEa7fM3fZPCdABR4SuUjv6ej
lRUX+xSnkXoymnSnAy8LFu2+ush1XSfjtl2ahthEUAxnliCgHsKgHkGUdBhu
gIcMPeWX5s0TPeoljWsavX4JSBBpDfnc0BN4x9Nx8EC2DeRCQwr6AnvaSHV/
4ZDWluwHFL6AD2ghxHb0v/OSQEFahOv197xSBEMXcyOkbHUxjqs9mYVJfbIT
L6rZ+pshsSpwQ/WTat6nYxRNVMcW1uYQPj0UpKMPxnRHPCHSWEQamvSkfYJa
0cseo04KE9ocTiqJ4iDzwdmp0X9O29e9F5oaYUOqgJuAVEm2brG4Jw6w3z+O
DX6VHmEujA4zC4lqYQmwIiHbfOBB5sdLP6+goVUR6Uv5kKhYEX93rGe6F3tU
w+25+LAQ053lh6M7VppTxRglYMDleF827sUcuHVLirJvUGyHGArQFBd75k6b
1jCjNSfa7UQ8i7yBY2tZdRGgW/XgIuJWjs7XTKG6Bq9H+d6kSnSbfgh9X4P4
11LycSpH6vVg7hOpGqRe33Ehytz329ZDJHsp4GUNE0r3YElUwL/VrCM2Idmw
LHhLNfyI0qzAhnGX8wFnghklTTGhzrcqAnrUr2Cpo1xtaHhB+bU7OLp1ZcFR
j3r/A5o/DlpB4oMaTePdRl8sU+Fh+KZwoJ0JuRTO8/qfDXFF5qETomR4qDPA
YiysYjuvAM+2NnGixIMGERBHB1ptTd4ORAaDBU9dStB3AxiRybtNErdOavJh
mqgAASG+Kvg9FPzai4EyAMTEzaXqGYvA27a2EsxYtEnAp3PhjOkq8ybce5rw
VpBqGgD64lFdytdBDPF7n1ootalEUyUN/2a3C6RVtiZlVRSQRKbZua6wpa+J
pEL3C68lPVkTC24HMS3QpKNgD7IPEuIgbUT4FbJ/dKwZPoPacHgHEp4dbi/E
48pvyNPSxC0/7ADjYey747ekIoRlEL3MbdPOMqR6zIG4KuumARjVZBFAbZRF
GGCNiCv/xO1j7srnMHnv/59/qxJo4w4ZQvNWxNEPeZFiSTWmxkcM8L1W33qE
Yb9MU3VwlfB0PYPzt+8cwkGkYKiGY4plfgpwj2CNrD7bXGUQL6v8BzK+a9cv
HrCx5Ycehee6EKGG2qkXqoF0873Z9KIkhj3nC1D+OgF7OJcEGkaDup7LVvcm
s4hz2GR7yMiLAd2pWvQxh/VYneR55ioDxFJosGFMZ9TgbD2Kk9P1b+m+5Q5o
GbFJu3gul36CbSYOQxm4cVprmSwCu5T4nzWrQ/+Un4hjHenphAgget7LdkCg
3bU3O4p01EZUau7rBzoxvFyEEVz1HY8E4k6sokPNJhOSY+DagfudKIcdOpce
H4fhDdPtdKNnB1AH8RJDXnOxqLw7yluLFD4A9A8Fkb9U05mEJkpoPLDQTFM9
AKRY46tsaZv0dWzvY4vbYqn7S+HcaZ/1+9lTNjrsyT7tjyUZaVjNPLe8Sn/G
dsoqeVTTN7AB+1Zd8v0mGT/800Dp9OG9a1mrjhmBhQ5thTkZy6l7Nb77SNvn
E6MwpkCLmOq4375/ijGYqWd6dBC+hztngTktGGAKpfAhCkNcWDjdt5EansM7
jY1Mac0cuKohKnRHgOMhz9/vHGwg4rbhVFHVctjVrS9MgeGETUif+GGCRf71
sgLlsi7xYT+4QAT3l3OdFfLCi15x/We0ycqB4ABbxd8eLjZjy1Vhk3yAxxPw
ql3enedCpfAjrl/b9ty8a6QKycI3+1xpahk098kcPTIo5Y2mmToFZ+99605W
8a9LjJxoiw1se4hPv61q4n2/dO2fM+6DUP1SZo7TopVeV9CuAP3ezvvgMAO2
DvqDrpOnYYSPeAlwN3+rkXjxuN9Q1KYtcYASYdGev6ajtoSTwHG9O5ZKDVUv
NmdpYGjoKzkrK3XN9NhqWTqYVI+LXVXMVWJP+6THfN8Y+xVafoad1gl7UpQH
nnoEndd3s5wkwfY1VAcyBCsuFZOmRJJcYvD5vD7axMiZn0EwnJF25mK/61Bm
s+6FBAtgsVZ+fgA5DDy3vADjE/zR+ZjyPhILXyOe9bR4l6GDJ2GethBhFQhk
uoRYduwmQRF8R9yqi5s28j+jFdzfnJYdcUK/7xUPkFoBgcR0LtJY6nXbTDpm
YjWhi0n5nVMAswWdAd2h0vAnxr+S98+9fIF2xcV20aPzT7sxWBbkbuO5R8n7
TF6GepG59pOXcQSoudKagXmHIUsFBfgwuiHh03cFX8nP/zz3UtMnVL3wFKQn
4gq7Ll0zzLQwV7B7182rR6iVPRyoadltVrBsnnN7tIpPYt2fN+9yyosQ60+8
hPvV1lhnSXbw0AF6Ixf8KKSazHEdVd4cIzpM/K0+Z4G1nUISF5mAMXbiwco+
yPsGIrnZvueepcIzKBNO9oKCiqPwx0KqcT4qHagNqfcgqie9fzswDBqVSEcU
bumLLrt+MDkqkVH2A9O3mBTVkBZS+KeTLZp8GrFfzt8yLXCZlgPIpE22Isjl
TbR4y5ZgP23+DYFD8C9865ihsMUOzdQM6JuXnHn8XMAuN3juHXAmdzh2RQl7
1MKhaf7T5mV8mxgDygs7ghxnZsrk3P+eeeAmUWqRzszzffqY5+yFLyQ9Ytxm
3SaGNKBFsN0RLhIV++jrcMy6bFZxJR9tCzB8DAJyzL+Kx4M09yGdj+4Vcdi2
mifqn4cv1sOur3A+W9VDuf2yosZ5Gxmmpj6v1Sm5ivCCgckaf7QzBmkkZdZ/
ra7BUj5YI0ATY4iNkDjTYacP5nsC8EjphjtzPqmoomIuWsb1G4TFuiBn1Z/M
wW6h+egOjCaixaNwFKuqeFo6cPtyBMKHpofKJP9RKjNpCUrk7W7VG4yUPv8z
QjkFPSFyvlBDgWBjmLRPeN92LVA8zlcDAExpGUwdAjEXuL1pbVL6b1b+OzpZ
2DapOVe/Xyv2e+kYJhDEUfhcibsdxoT67mAjIy7X9j1kuYbICaDtEJFsE/Ig
Ale9BDDxlEFo7Q0w7OZ+DdE05dT716Sjyr7VUVlX5ZfURKDEMPjRvYT7wpJ9
Mq/TM0A+8P0L8ndclVR15NGp+HUwlwjbF9AlTMpAwuUnPJ7rFwzKtxv6mJ6Q
DesS55b3zYbMuwDi/q/rz61rJ7PFirYbep1koJJ5o/0ga5gc5boLaMnxQU9/
AxaSF4TnpRgnLtTVjn4Kr8v74Sstmd1z+hCqJBWJpVpl3YHIJKa7xSc0j4w9
7LzwlOSuqe8JsBUAJT0ojw0wg2Ku9aUfRzrg/9ov+KjP2pxyaCVGUcPN0vFs
deiZXbQsalRCB8roxoFB6F0KdINbM/r7IV3k7ISCSRG/18TB0hIGbQ/6DMA6
2cDoOzPh1MZ1yeeWWUGBLcy2jGhtvlYHkltxo0XsK7N/uGLC8P6v/7UY4itc
b7JGc7h9X/4eFfOSjZ57Fevn+pJtb4xmRPaT40tvVUEW4STTTc9SOjtgpQEQ
aZ2qSdqSi0i6t+JlJzH+2g7xBNXbmUsu0yKIS5fAxteJuEPRq6t8ijgFVjR9
+QuaonHlP2mbokE/DlvtjntkWZfU4RrQIrUZJNR7yI/rie4R7Av4M8Xh7dhl
31VY5BnutCz4WJvSaROB4I/2S+9evn5h6uPHxJoDb8BDTzX+mVBNTnNSvoa9
/Hxo0gf+KmmMWQUyLJFQA1fRbR2gUZufiYg5PwyAeQTEQ+YpW1ELOhwhxBca
uZkW02z5wRuB9aAKdv0Bw6WXP3T2z4KILI9MnkhafRW0QmuEV2UlaijaWj4c
XpV7WYDr66v3JufB67CvziZynEy9tEV2gpssiDT30+pFblIvOhCLtVCyhXQW
cMAeFpoyYC1/e931VcZh8aOkRvzImvaCcljY7aE/dmcittoDpJpr/YAx8O4n
cu88UrnJ02AkB4Y6CG9sSuPktkLC/k7kg3LCElPnzHbowQgrecOLZd6ShyWF
YZbDWok9YTyMDAOKKZfcBU/asRBkpKbrdoNcvI8U6c5Yy29bdM7KCY0GJ2Dj
Owb5V4MW+z0yLw8vcyfvC6j0NZf74DVV5/MQvGdv/Xm4Tf9PSpDeUKpW5hIB
gwU22Met3ZBNHFmsZLd+1/77OX1Ch+QeJh/gS9sM4D4XtsnScrgNxU5kCbW4
hzcbAVNgIw1ORDl+/hqRgqt0CdRge0TiN5iNvq3wR1sPKz0cRndYSihGorDh
mdaTi0tnlcwDCClci1kn1Z4hMwOPJXK6JulGufk1R9Q/qLGuA7oI2wuDoUqj
gEHEbtnyIix2gfj+ks0w+HHeQRsT1AIezc7k88Wr8Ell95gkf6AmcAczIMIA
ajYGI3fqFbQzbV9uv77thqtMhKyg2Ky/yInfeqvepfeaRRgPyC+fC9MKViKN
wcqLUhXoQxuKUXemFoW6chc3wtUHmeii8KbfFE8RYjWIvdP2gaGyBNZAx+wr
r9s71xViWOaj1hOd20PtWt/anZcCVMid2JLAIGgDigUojr5fTZdodQnQFY4U
mcfQ8ngc96nCcLoSQaDXCbiqX8eN6e5L5vZMA++yaoNE0WiDottQq6HH1kl3
WrEfiokat39jkleg0WO8O3SSekOHI4h7BQ9jlF7U8vRQpEYQPdfs7b68kOtm
nr9ZxyzSrNjCYzz6qs0b1kKYKbb8frDwp22E979sMNvI+ilFLuPp/ng5nldv
gCmiJyIkUFvnYwsP9QwDPuenlOrlAuTmsQt2libUmeXOe62dy0kb87JbS+he
yoPYYWKYFidbRD3UshWQfti2PxfxLnwYXOQU6l9pD14+EKSoLPtwF7GVKkGW
k3JWkn1RiIm1YI/dEhbq75hV7lokiM6rdhHfVkcP79xuRJdWVAClHMUvRzlG
mgtBLBKKGISOOVxp3JfR6BzJTB0avBKTvbooftCbpvCwda+wgN1NAtmaL3Y6
RrlHrOhvEG35lzjsZC/xiimG4x5dJ04uZ9uYC8acbrO+hKa5hLJBQv992w2B
CvIx1wy/geavA2J7965kldtns+/v0QN0DGS+urJap13wiGx62z6pbpE1q8xY
SQVl4AXyqJCrv9nUWiZuUiXUTGwUSdCGBVuXE1VqToujfZhtCxMlad5QTUgY
ueKHHX00Klw9dVrHfFlp2uqxcB/jPVSv6Y6XbutL5PPp1tPk6Tx+vGYY9YiX
CX4lG8L6+Ls7rXKk8WkG80BlqwqK5k3lvaTxhc1ldcpZhjMGKpnnslJXRPoM
t+M+yEp+qo+Hq10x5BEqBl+QenkSJ6+qGY4JSvRk81DJG9uajRkIR0OfJJx1
l8t1Q8PIIuJVfAV3ga1hJG/7/L1S7xlntu0h7xobHVbDg73mKRqo+mFn86Zf
csGL49e2W3m6wAo5ET526k2wdbn2edyPeqBJL34K7v33kY5u57uRMdj/jJmD
BCN/VvMr7c4b5apBVOGTcv6U/YRy+Zma0rYfPrR2dkVgCN0HRl4DMtWXBYuA
EDntJD4EXBTm7TEbAbwICCi+ya1WxPzqz5A9mKdDyiAsfKDl1f1SCXvklyn+
x+OTTIVule6+HEmeMuNAkL3EprmB7WRo+n1vatuPmvOg5bRdNFKC+tVxqXT+
5/pXxPDYCLC1kPbn5NeP54AXhQlEWB3iwRnievQ+M3MIPTW+cVGw4CdDy1oP
OSxvF+8/JCgWZNfeRU4Eacs53lurEA274/zw9XUD2s2RYPGKXQfVSAjvzyqC
6j3L5MvnrrfpVcyuFe/t52Mia9N7A5Dv76E2Wmwyxk7L1QwOrOIbnOz8Rrwt
7RbMj032r3ZSi3minl7xBeJrbC6yeQvu1+eEaU9FKoTQc7gkctBBhw15yFFc
rxW6z6ojHJ+FF1HGabq7YV+DTuE66OWjXHDUCpzW2i/PnqMck2gVERFTTLAT
nH8PTQAcPB2e+W7S0SgXrUoDaYZWI2nKefa3DAFnlioMzT+KRUKOt4pECwcq
XKa40GHaMaoUzk4776LMyrutroUSz461S4zndmlyBwI39A29GxFWlyN9i3O6
y6q4HqO2J633+S4WoyYZhdsG/kpGoN1uXzYdT5VV61or51oAWHevciNKlaV4
IzfJNtzp5ClAYtL5Rimf1duTXqxeiugk/V2pdSDve89cpFCrsMi3w8ZNUyXL
uoe0ZWgV0tQ+PeEsyU+4xZoaf6+6FyGS53Jq9pBlC22Ceib5r4bmqX6aQWTc
FZlH+kBdT1UE5QewjqaYCoAtkXRoEv2nnpoUvW16nByIPhh9joqR05QqWUI2
BG0I+T+8OSwJCS40KBAU2+cedJs3h7+SgfHQ6lwWPnz4aFBZqKWXPC3hFZum
QuZC0tpfAAF+n8Pg2B+ut+Bya2hdxzegeJjgT5uwa0YK5PigwIgxzXWuaD8r
ZTdRmXQ+rxQCWLAoxw8uok/vOa0TjccNlmA4UT7nZO2Gq73i6Oziy5Bxm0i2
PFrAQhu6hOVEu4ghNjcRbhmK6PrnCzEYNyCNl6W61IPm6QUqkk2C0jcart2w
oSmCm+avdjbQu4G8W/7LKrOf+tPTvvfQzmyQ1d38F84yMD23XE5Se3qN9MGo
IEZAbaEIDnHSjuRcNSPZ5E4JWxZeb17PPlHV8Ig3NgNzyH9nmwjnmqvf4Gyt
DDJ11lciLDlHqo4K9WY5yieW/n5Qgon+tvOB822Snu2Op8Y+aXbtt35+LojK
jHygf11UXLxxxp/VOOeNeuAQcR9kjD+EQdE7zX3E0yF3yqB+6ZLWTRXYEURX
5PxrUbtuBOpikQA9hQfOHcWh2/7gXlhLEVHUhIu403PW+XZsyaUu1qdkyfQm
07nkNG0zTW1IbXJtiVipjxkv1zS0gTVkAwJ9PC7iTxAorAbreV61pbubIwZo
4owVYWtQb9zpWJvUzuXO42MzoQ+eVMckHQnRSnuRSq1/z6GgEaluKqmhY2W9
uzMgWzanG1WmqgSOdZC4iV9XOHhCu1hMjGD0eeCIDZF/CI/RvBFTMfEf5nlO
qfIa4dE1ksMvnkylaKF3b0fMIvX0sfjX6qcZLddoPe+4+eIToLOShvTwf2cn
nxRSPQW5U/ghVlWI9vAJtupbfonw3ZcUEd6R/fhaHopIN4Jit9vGmBN1d+IO
pdutbrCgvyXLPC8F68i1qp8sFlEnBtZV+4HveSb05H27Wv4JB8Lss1aICUwH
CLqfz4yw+e9715uP2LpGKGxyl1RXJsJF29dpbKqucmVIQssL9qbdyXRtxvQu
RhFzyfpmnAw2lqIMxNNBRUBnEc/VcRw3cCc2fU2s9qmiqeETW6ZNN999Jgnp
z1HNT/bKKUgKVX8vjL4TB1sJJcc0gTvUyyX+aq5K3+pRh7nqIbsh0SgZqSwz
1/xiaexgoDccUGdYKzqsqR/78vUovoFuYwiik6eOVQSLu9uCLFkcbG7iLm62
TWXPaxHzFNVADjRIXeSLmjW6MSvxBv39b5OI9CZTdGukRmTMxUST7tj45jor
hln1GeJTmv+CKOcuV0HCufoB2tySzCm8Orvtuabgm54pG+KZeoc5f3+5nuja
XU7+vyejO//KFSPgBHzj7Rw/6M6MHU+7tsQNZec8pBXqqtdip3IKXFYb3lJo
ZT/MdWhdWiWiMx7h8MyaX4AN9FXYP1Ljgmt8sY0/8W95MJyTl+qazmitKPw3
MlGKtHI4vnC9rjhHCjILNsV/xfTxT2UuCH3NoV6j2Pv/qKDxSKbMQRUHy5HA
i9HbxpMX4PBUkDyfz1soPS+s0dKCSsUr35DUYWk2lvkH8RXdL8wm2d0SC9X7
/gl5zv0CvlQg4VHXBq3vywJMtN5ij57oTgzx+JoLm3YWc3azKK4FtefBnFnE
LQSOak8BxWxWE8aKaUuxk4yGQCyJlyhfN49VgUXcrEkydGpzB9Z12eKNlEj4
wcW1yz8zxsRJS0EUioc2xZaSa5bBalJiq6ONYHypLElVlN3IBBb9/hWVCjtZ
ttKfbtacbzR9zqGrOlan5ajk6gGd/dn2NqUv5Eon7Z3creXrowGsbP8b0WiO
9W/VZzqofI3oHFmR/TmafMBR6aRMLVsizz9tD2xNJsPiIcfgpzd0igyeJseA
CzDj7vNhjHZQEZkbdTDnQZ6x6ltNDkPBq6syfKVjRY8xPpD8z8mrPsQKsKAJ
NM5tHDqC7FgxDOJD71VwDi1LB2MB3KVNdGA91XEwiRyRiGExZtPBYYwaY112
YeUZA3KJcV2p5oBQsKrEpJ+Y+H4zP2nP1Hg7u5J392etKfqA90IBJdRJeDP0
EL28b9Dws1qMEZGcVmH30JM534B11cacQC/48KYt/myD0veU8pcHh45CY82T
+ycphIWaDFzldiQXzETZ1xbrrFmKJcai5Mdqj/J9Scu8qaPRxJTq9+1YprGG
qHxRCxA+hss1hsi6Hr3cJg/sUtnsWxGRBKaodMMpWdpZgyYMRTVDo+H0nXdB
MsjfAxjxGGrwS49G94lKn2KjklH18ziinRDr0P/QORT8S6NFW6E4/SonB0Va
/X877nAwBYF7b+HQC6REYQDQh+hwtOzYmiwztXdQoFtAG9YAwXMLx/d0st8v
AbtvHGVIxp0Jt/jk37Jz+yVIrkrJrupoRDNbf69Q7mWKZu5hr5/iRJnI0RaA
NhGZnP4SZaCiGxILqRN6Q3OPZNI3+kDXUZA8+kO4x+bsP4uIvvcsKB86HQcj
+EpaT7p5dWCmcAlWAqY/Zvba+g/OyS9oNeEH3lNbzAJq2/3/vwbtAV7zEaHr
KCpTYSoMWRz8ayRNuyml/0OJ39QKWfDUlM4fP40wLWDSjzWrE1SkOiIHD/XW
XgXgno8c0JfCCLAxV3HZAhi9wI/nvTAu3rUSPdi7Jzsva+UgNgQUMrStUuJS
FE9UXT7GWqCV/CjSRKFGy1uRod0RPA4EznIeUYHjm2n+Yi576KyGS1A0ugiC
QisFV/2aLFGz75ajYHbOtb/Ko9GA0to4thE9DjCY5pi/dIhGuvyuSYkhNcyI
VaGol7iUUv1EeuyCqLl+00OY7K4dCTytUdPJaCnvJXwFgVUoGxYlrwD7t/Wv
l2RTGKvq6n9FqxQygh8SbHP09vJH/tCo2jM7JPANCQkjls4ldovu7kLaT5tf
AgZIMmCMvMt3LxVg2EVjf1Gr+fmxOIJNcSCL0ZVqk3EWzgoWHnzI/69ocTmf
nUV+qzYGqmq3ieNSccXiahmpLNfC4zHz5VICxPCE6B11Y8QEfJw+zCtdzhOS
DkDv3KzG5/g9hy+M4z66o1h74xMoC23yBUVdAs0CVH0ygJxMbgz/aC3+hNpM
aIgNhuUUwD8zy2q2esc/pGsttSAVrXG40g/j+SDoxmIL1YNtBIWBP+y582Eh
9j5FlbZi3BA31doPWrKxBmXmwIpgJ2Fl9UmZk7/ew6FcKHxJBEm7YiEYAvHI
WLa1Rq+/QXeUjo1yecYwcJsbBe694iRZNZxLUp1OqImh/qXbGfbllLgsqi/j
B4vViTIPeqBbiHNk6x3Sub4wi/HkJkcigORLKXporCUmsiMRvpxuaCeCyuci
BTEYU4GaJ3j2V64XYkRPgn4u0UuDSpL7W3yDwjUPYs8IotaAQFjSUT+pImPf
kJC3PKZ1icxe0qi4AaY2Biz7S6LWEuYc5zxgA3BM0a46S5I1rZIv61HV8+V8
iUp7X2QG9IFzoCbifBKsnr+PCldDkh+151tLDVV0YJAXHoouypHMuuPzbIML
bn6iID47YUzmfMYJvx343fRlv5NqelYx5yuq8DmHSzl2g6kBxsjsX/l08/9a
VEezoIal/Ny0FC1CqSGvGKQw137AymLRTCqIEUk8AlrFN4cwC6OhJXbPjv0w
30/d9LI6jzsu5sLKyhXzqjWlhRZUV7U7r+QNBl0TvTzfD4I7x2VZiP6EKWd1
jsc/dz58nKhlenA4h3EdUGMKqhuP7fKu+RG4DC5OmMjf2DGBMOBYGfIrjfu/
JLRVDPDNGJ7DKjzCgRdTPhn1DVZ2VJfgOqbQbI6Gt9rXB8DvHdLp5nzMhtlc
IiVN2m11VXltqqfE8u/L583PdgBYNqTy5TcSMLxn0izCAjAnG/TY5m5BrSf6
/zbcT0CpX0NeJeMckxWbLzoaBWATkjyzolx+pSqrhjk3SUfmXx6BMyZwgRLf
K+Rfm6cH3RnpMplD+ZAGERcqmJyJm9D36Y4NWHMYlO9q5cOGYEJmXdDHQ4Vr
G8qz7LEw9CTmC2O2IW504sMKdhCVqlBkAqPovhDZHPEDlxawZk4m7L+/D6I4
Lhmc1f/owo1Q2rEaFzXtR1hh/nNCfYOrSL/CsKpZU+MSJnSfIn0dczUdPkCC
aaVZO6EltnpCcbyXBvjFwVs4RMpaJBnnkIMD3ZlSrdiTSrLrAVTtXd5n76ov
wQqiBkZsSaO6v7+fDZNg7RqPkMF28kg+zlgW0csEMeV6UaGpbDWcKqDopQ6u
FEyfUtU6RrFfv9USR/ArUOHPzpw6f0WV3ggsFFBxTl0QV/Fgl43szR8Jb1Hf
Y6cszUozIaO2JvRyatWp19DCGJzk3MhpA3L2lHdD8bIsrPxqd/tciG8IAPI7
etyYLjrnVxVNBX41rtE4rSFeZPRwqMnu55LgGkrjzt/KqAoG0h/z91e1ssaF
66jQlHsMWhLYTH4uIIUx5i7FQz9YTgO6vgoEymIMhoTPipS3DNQySof6iKE3
RQyd+WgBL4Ds1g2uoLtYN84F3M94StLUAVNPLlk8C9gEt86hy2rq0HOFKSx/
wsXUaK+sGWK9Y5R8JYvQnGZFoqARC8vQdufbtuYvUmJT3eNBgtmKVTDxinmS
zoiXh2diy+TDkBv36oLyLut2WwTG/m/3JzIdqco+0MhmPRj7HdrhRBT3xvUY
BK8BGMou6/5oD0od0Bm9ReuluCK15UU6C9x8M5TvccB+1zjcO4yLA9Nx2UXx
Sw4nzHyIPZDq+vvf4Pld6Nfh2YAje2ptSBCIGdUuM+s5L5FO1b1+6AKawiHO
+I0XKr84/AweykZXnXO0B/ue3YULffvNz1uAfPobZ4tzZ7sVWNMbrBtTgIua
YrC+ko5/JEtD6NJOvBnMdXI/+omu8qCyC+m4Kg2kMceXTEliFBiHUnoom5PP
kLDOt5zd52I/wuazaSFRKfifv3dSmngBf0u7RAVzx7jjVHMsFjOIHujENIz2
PS62LBWfqJVtuT+SvPZ3b6lGSANO8HB9i/3BxaAjR1GjBYyWu4ytnpts9E2P
ALXKgVXCtdqeb8R1A7j69ECj10zpeETJGVf6UFe24hTzm+0vcBBQTIMb+HYG
Zg2tJ+Wcf65whe+dZ9ja11UIA0mZsJB+brKXZpdqs+uqTXtWd0h4TUSnO+TT
HfKFHZWrxrk/Ttg8yJqVW5YN4+OXbPKLPHgSHWnxejVd4zOhPMTj0nnZyAKJ
W27AoEmWPa3RTRV0RLmg+DpxJZmcAReCkwv+uHeSgLr2lIEqZx+uLGEtzVKs
0+HvWaHWr8KdkZiXHfGOgDUjJYw3+XZzuiCuXKwysMEwnydCbFartoI4DDs1
/Oj5gSD5lwEEkPJUlI4Ck/C2lXbpDzGxiVsKqlNCndRjGya3VMnKc81j2y3y
7OjE5rVLBB+ESODepepegnUN2ztswaIqmVnxyRMP3FCMjH3MJHIe1CZeVN4o
31j9B5RuoN+xZUIlwj9ZrLTZ1en1QVuFqmvbeKcNBHgZF1QUuXB2vBLpjYaW
Et1qgaj8S4OzGw0t04gFbWlKWXvQWJKURNPVIVdKpTLFUgO6dBa41D6PLTtt
ihPu6/K8XQDh6a0gZogc8zFNdQD/tAgxtmnO/MIdel1N0UfaFUFo44sk1thG
roxGhooJq2sTqTtNEXRDE8onFR7XG8sCsLPxznv7G7Y7zuZ0FWY9fEhhc4qk
9WNu4koAg8rMlcAOOSVLOfGTkJoSq5n10oPaEvQbsdGrrUjsoMB4w6Y+Dvel
g1Quf9ZhmyU+nQiR0LRhxQxnULCYSEBXHqlKVP939bZkNYW7IvmTF/Xb6pNd
604INyRc1RgNG7OAjBtSYfI67qmWUaORszEjHYqv8e+N/0sWTWMim01u/rig
v4LA/ZhHXza1c4Fe2WppRJbWNOFtjF5kL8Vzh4yNrXHI1FbL6f+5naLnQuF8
zrsBlLc2AnjkrqqXIRLC4vKTfD4ZPqY3H7OEViodcySJPF2QxUNFi0OeH86M
2NzSaDQZMNiwoIvZfjzDQDWxhjaqfYWydXJN1BwKriUQGFwusaxk2ROKOB5y
lT+KQyeMcp/wtQlcIf3xCmOrE6IuArgwTsBxXJs/eAj3roWKvzcqjaH0Ed55
psAoGE6nMju6TEeB2sqgBFKUEzYkwwmLBZIN3Kl5FdZsiRe+ZL5ThZyLP8Z9
ea5Jhr3EVpPGBozZ/v05k9vu2KvUL7QrtY6s0Hj4uehF3TpOT1eUDLvvWf/2
kH2hm6cmDpqcdyyIci/hpysROB2fW/KFjNuPf7IQkzejnMrJO3Pz4FJghgND
uaOfAKukGHEqOPSWzq+/QrMIGX5xTRF3HteAtgPDvsKc3YVhAYhPfywzrMjX
cvRTrwbFbpzuYppdbE0L/srlPnPMOr/mtm9HDnt+jg2D6sPCzcHZF326V93x
O3s4SBahCtDK5CkmjEiD5JfV8XEYlADTAJoMHTjnR8ed+g54UmvAZIllhg99
2OIHo8D+217Fz/hRWD5Erm59mu7zq0Y4hJKXT2tLiHsH9P6gNpANNejCs9TT
2bqSZWoF2EstMRZicVDvLXnZmS24tKYWqfo+0Ey/w4lpYlu0fCKZs4F2s63I
VxULqrvxi8CckLyGAG/aeuzjD7ytiLYHSwsMdY2ngy4JbxVEsrVeKXD2BIxT
TbD6sNisErrfRH3P8dems4hj0dK27BKW/lGHOQcyXUZItIzrA47IjHe3HDhC
ou/6ndbDwARCYXZLbhVpLHINlInQBHuxP4B0D4vI7fXqemYt1jkfSqMwYyHu
IQhK+7TJSqMCekEIX5s1fVMIQIjXaKaomyhzxDWqHj5aNG8z03VyH8iOVGX5
TOb5K0sqhAk3jIPbUtgOW2Hvvs9SNDN1qsujLA6NWovdcmcRtCZB4b0Ehtcd
RxwuB6DPrNLscrAocgJpufLh27sRC0VqnStd+es0aHV7mlfRtwscmmRmGgwp
Fz5oDboKun+YVM8FdOryLqgCsR7GymhiiY/HqzJTJwcHd7j4MJQfpj0GaDC6
qai+mCnGICY5w/aQzsdHbAfwDPNc+p4QbrnCMugeZvD0BEtCHFvBqnmMuRyQ
2Gr8jAsx94XWtjtbErM+zD5bfnmKGr6OE3hWhHBlMcOBzLXm9Jl9rUiS1KQH
DHqQwGf1NP4ETNpO6qbYxbt76LS3Sw0rEhmOkPSNclxUYUqGV8P2EvjPz3r7
uaSw6ULwzdwEtdvaLO5/pZJlv1R6ghZ8pW4wel1xEXK+UM8cjzfn1ejpVP6H
/YN0+urZNMWahfYc3MjKEpiRqMHp6W7GDwvOFUsAkWYYB3fEbIAXrG35vtkT
D6Jf1lvUSj3GCe0hX+uYXX42geQVUgurVb6eyJQO37Yg8xTHM/L5oRzkExbm
Ifi8RcCVwk7NYtz/5ac2mYY/MqPH0iUCyaPTXq+cGWvShkwhIq95FolBash9
CpqZllVjW4FwmFbdv5oZa/mQkYwyXLYRxURDKFuaN3N6lTQl6EdTA1L0GDfb
sWuUgRMQeQ7ykz4ICGrGzps3BQjurvvxg2HQ848HzlGhrm9OkVJW9oPSMfpG
u8isuwSr2hFwlIe3pEsAfTOlZZ0leuU3GLQrZloeblhaX80TbbIEC2WMEbpW
ya6BH6r6dFTIr/0SMbmlAQBFGXOmS3YkNzug/yV+TT0VNbkvyJkxeFbxTrz9
K4Qaj9ZUFIjdMcWiaU6FgbKB7NC370vM0og8AyEmhLnTSDwL18l5GKRSQNZ/
S6VX/cgI8Tc3C4jg7f0ZRkVHW4aIkvfnpZAmtWsqU6IhARE81K2Mo1gxDtyj
wqa4QuQ1hPfi6y1zdqOExl7rzh/buZlSmVLSxqTSZhOVpF7rluUt+UWihsVD
bAw1P70iSxEjDWjSpI5kY7DV5VYao/aZ6B08dv5x+3bv/O62HLM3U+tTSqp+
FU+3ll9Jw2rPc+ZK4orJ6a1RvpOhwW/3+QTppeU0KMQuH8vcVaGHztSzsR+2
QxaVoXqadGHfy+1LvYcBGUR8X4TIA3B+xfeTNin0cKD9Wi4in/4MfDCSoCyY
/AilmLCanYW+KF84lJgYdpOPQ5FMu1cL05ighIOZQP5J8or+oKJLB7lVVD1t
Fvhpr4vdPnxecmZEQUQa/aU/amgKG+uZjCQ7FqFSPN6XCS6NSQmmalgZGLm5
LofyfrEjOQdmIh0teeDQMq7hP32S4qjOgvXTYj2W1Rg/zUlDT+spwfEFtwKX
G7tLTPFmL7nvG4kfFjKffWkViv9S2nVUPGg27Zr9cIZOtxOxynCOywnlziWn
G1PGCVIgIh2qyEeoMXZInBZxTBZLzLhwAui7dD/EVP0yB74pchUWyExL/mBo
6rrFG4kBpb3z+9akKVlWydeTydL6tmYYOcKkeRBGpNG7QXoGM9LU6SwpToIQ
pUOxWP2Fn1wZ1mvjRsgTT1zmVM4eHb68gXQv3L9EV+Twc8FVFYfThdQw8wHs
zOsgSePaK9uoMnOoDbJ+UERmivRBPQ9L+5goO4Is1aK0cF6L3ph4cEUZIU/u
qbVdtX1DTHLwv2nNOF2JnvY+yh/F+SreF3tthzO42BBA0NuTEuIBB8qwcdlf
NXoLrNr/tV//DKMAVmRZwZfDZfGxvfMsQ2HdS3K37tBdDJQ965b5wI6Jgyxa
HUvF3h3UaBac1pjzoQT1w88qmzyktkwXY2RN1NNNT34cBuO77ZXLmAnV830Z
KkTIiMgNh9WAG26abWR4oKzV9fOdaTRomee/wLBvZqEX+LpKM732GGYuUHr/
gVakDQO6EpdgaamdvFWcRsLKYtq7WwUYQV9OLB7g0/4dcGaQSo2Dd0KjAT6X
xS3/OMvJ/cpOzpAyMI1F55ZurqNSSOY3FR5O2mpzNfm/bLSwK1mQbMGiLVEv
Ipw7VcM+/1NkhLUmqwsZQOHNiwU9fh5nngqGA7NzzKOdRdfMpdF9aVvCAgq+
6z1Jq1vivyghADUjRlvJ2L5dzhxWEn/NvLqKyz7FxdYf9GbIxwU+0yIvayyf
53e7hwhH1lgqXFc7IMnFEkTZmSrktCEGi/aCoxfDUauU1Z96w4Lo+37sxqkO
6u02nWkk0s/YTZwwq+btdWVSJWn7iPEms+f5pZvsXQ0luKWDEbi8L1nEdx0A
fDYPuktZ4kwOvFI4vuDAXcZm+5FFmnTZwICYniO9DfaeNrSxQfUrzxM0RAXw
lKor4Uzr8OUGDAtUjPrRsWx3Bo+GHIb/wPzlb/m72ivAZV7+HMvbQRCtlous
Wg+oWBxjEZVLbAjoH3Z11PsR4OhGvyO7Ei+ngZC5R/E5JCRrlfei+8GxpgXb
nwGc6QvgnI+foTYFlyT4uhGdYvqbU0xAuyjOBtrSoaFMkDWG82Ny3XrPpZg8
OylDwDEHZEHjnA1/VeQKX8ecRsI0+zOKIDiuMw9LMTTKqgHAmeEcTtYbnfc0
WkeS7Eb4ArEumAo8/3juLZynBQSdfiVFQPPRhrBKozhyCWx/cPhkzDOu6Wpz
DIAj5a/m1LYfuT6lCKTzwp+ycWcwWWy43iUEslndCkgmeb2YO8srj/3CPT+v
bhiiRmYTRTBe2mgoWf+RRUFUK4mWqh9OTLFN7qRDIvAcBYNXutWVZN7Pm4J8
gpklWG3r+tocf6qGEyhrjw4pRuw+hgDTm7FErjOCswCfjI0v/iYWh6s/NqQv
H6+vSTCeT5GYZYRR2eb1R44KZ3vV9j10y/H4fyeVjCT9Z5Xa9Ra/c5CPC0Zp
uDiRzLTmP7QQObFwZmIl3DPeaPXKKSU90PB16nwKSp17mlGnSH9Zb+7SKGY7
j+RFc10sP7VUgi1QOu/qhxZWaSPb/2d2va4IW+04KO16B2bCstPzfnYcHlap
JvR5540Cx8TG0rBi+Vcd9g05C3MXc+H+u470CVkTYTsfH9ME7M2qJEWacAX7
2yNTcuIuphrcnci1wnFLyGORixgKexRcVHNi+g/Gb84kkpGu6cb7UvjZRfyF
Ru9Bcg3BxzWdFvBLxL5B0/dz1+vAEj+8mQWrUzk+NsmtouwMbaHMN5Vd1xrH
FB7jBK09KzhM4DtlE6vnmjynpt6AteF4XkiGhyYQVf24/SjlMQwMq2158Nx5
BbqRTh7M3CktUbRalX5QBoGSAtQNtIiV1YKiP1zTUeN4tjD2heMQ/Jl4mLsY
WPgE8uTNEilLaL2gxbahH1xOBtWDJ5RU4PPkGCvgt+BfyQsXQICUs9w9eNe4
23N/OFH78E5gvIGzoxb6yCP7y9SQGtZO9etkLcE402mi931EoIg3/z3tOhuY
O82kzGl5QUu6MCmg/27uIKuHHHtS0dHTz927Cric/vJEE2tg/C72kE8RuOoT
YV//7IYdAjU++RNSZNz3xpZdwSJkjjgc/8iZa5aj2EeXTRMZ73kRA7JrmdPL
Y/3BKaf5SDEoolJC65YW88YtQwj98Ehobho8sLRx8LvX1rWjgxWEeY34e4Vh
2t0pZ+NFJxJjP5aC34kgBd7eeuycAxdu6sBdR17ppg7j17jPRJomegMZNwzP
MmXaMd+6r1q/rO5aOl8Es3BQ8umMgT10XWkw9MwPcD/0fxLYt2e6E0isKDtn
T6aDRbKUTbhubmNFo5fOkBZugyuiSQEQFvBdiu0JvqCne991Ox8PWVAtFZUj
DfK9EUbHCUcLWn0W9QtWBYukXqnvBhLbTMkX6Kzc0QnzAVO2yJzRoUL8BRc0
6/jb1NT+0gbtluXRqQTh+CJnJy+5G2kPJxJ7sGBnDCRnsIqR6iSGN168ik+7
g7JKigwaLfXAxPN3khsSFNITTjE31RYgb4kyN40A+qHg+UwkXcVhFL1KpsyH
LULfsrFs5PwHcgqlmAYDSxh7HqVlozyO2AZBYIhN3lK+aeTJGHS/cQfzjm8E
qMusaXDXVJEH4NNQPLPhq3j1QiAiCYcGWt0Q3v8qAT91BfSi5gWXutqzcT6/
XsPkOCVmOOI6+FS+vsfhvnOkC26QZAOd2T2yI05IwQDg7BJeQAfNA2jhteDL
VvFAN4W1G8YbXLoGofYtXNZyIeiHHM28vSmhP3FaTH4vILEwUAQqYo6HeY+7
nxsSDqiZgVKUboMc0O864NJ0CTahZWu8VunuC6dQgIz6YXsOsQkfHZF5lbMR
yeuu1cldknSxcGFQ0cC8oq84ebpo9DRUIk1kg7KGDJFqXPHE0haah9XryrGu
O1ILyi3k44t7DVD06l/M96PJ8vsJJFcCRMMxsUnMaExaLhyCwAmPHx5fK1hu
jXdeE0s8pvrVL/mJ0Ufj3fQy09XSWVrhsIPkOVXrTNv6347b9MtSwoIvOGPU
beoFWfgbilYq98IQTJMf3x96svTdtNe00qez2fv8q7NuAMdnoAwGsppxR4Sa
sHxYvRpsyP9OKAS4GMB8+r46IUmz3x7lcKmgufaC4dduM7v0XBtdbt2iRFS6
DE2qg/S14yZ6Gv4FjKCZPXPhQzVk6SR8qBvko+s3gB5KLBGv+rRoq+jh3+mk
yKZMOzOagGk1W53/9sWUqmWaiwDOPi+zkA6+E2TL1/MDsdSnQoP+yJ+lA0v2
omKaBIdEvR5oCbUaSfpLZGun8byK92QInSG6+rJMeaS7nb2PmvxBGn3qsVcB
F9dfANt0Ja6E6TRNAJlmTEmbgCull3lBM6GvzqLYi5J98PmuU4L+oOR7IL4N
dsIZtXHZYGnn9eX5qGKd/VUMtIT5NLBJmqGn7wBPkxqUVN+/Nobrz+gQEQM5
ADCsQqIuVZI7AL/qn4XTmgaarRnNJ/FlIrrnCSRO2oFSt3/PZIW654nSMBXG
msN46maV7qmwe7wXRuMgbVC12ZLdqqKV1+gqlnRGxRXJ5JnRZLqUHHud7o87
20c8m51gZ3yIV740Yi+AsBA6Q/ej37xd/yJ8zpIJkcIE85jBpmITUs93YTI2
JKOgpjopj+9fNdxsQ/NgZGDisJnaWTqQD7yhkwprL84GbXKZDHUZXU9OLm4W
hxsNjOUpt5JNRsIzt9hi78MuO/kaeTRrtP10N1JHMmUoUWBQKzs2QhT4c4mQ
xFyUNyaRmAmXJiQdpGRHpGP1pPb1BBDp+El1UfYYGXC16h6xQUiPqCIczFUl
t8ZoIT6AKrJbjiXevfkTC19kI9uNonQrT71P3hf/l+Wg1H7+4GN/3ZlCaP5M
VhLbCE0Oyh8kzCdltnhZtr17pJyx59X7UKAF6FcJ1/qLJZzaUjWpKV8ESMgw
SIDitOxjittv6G5XlyO8GMCbf+1t3yseafwkr3h/CRlwZBczzXJVnLUUNNWN
5nd8ZUXR1J8G/8xyIJ/Pevp1+7n65ocP+IodA3zcmTCtqfzSmIvc2VK4ub5m
va3fHQsYA7kWbFFLU6Kiz9AjHEVVusGye3DYqiEXVKUj3AdibL9erI9EAE6H
0kMYsfSkF+LBBRII525+sC/Q1YH4Y2hHKTZUxHAW/vf9b3SUK3XD9OOjUWYM
c1PbB/XDu+9ltWq9fa0LKfLPFXhOEZKD8uQkXEoa20L2ZlyKYqCMd6Ff3CQu
EM31x6s+Xgd34YZKJ/B0faM1RWp6Uk0JwkGRTEnv9KfVBwiKK9STA/oJVgmc
SEII7xBtnkNCgUIn5Ry6ZPUNbt2atjoO1v1lMGNpPhEhB8eGEcnvU1YX456R
DfcJo0RsVpQWYSu3Z9eQvr1plF0Z2QLv+X3loQ16kKCkQOTp1Td3mhtgXsNr
1k3jXTNiJWc+G1k4dMsFwj6tax+Wf3ajAL5WchbebEiiCgwuwkZvKJ2Qwsq8
60i9I7fTWDfSjslN/xZxS3lJfYrfvP7J6saeksNx+1bCoqXn2Q50AheQPcKS
lKghKnDxf4DeUaWtyZsETFXiscNFq8Y17wpwUmJb+2al5gC8eYYvgxC00gfT
mLYDvEcTfNUtzNuFcLbkKHhU6WDP8HYcitrtMOVL4wT8sfSUY9vn1KwSEGKD
A4egn9KBdOSk9Il8A7RIvn7Zoix6PSLdJZOEy6fcKshqLbz6S9UymeADG4hi
hOx8gxFTuHIKFIpPpArB+9Ds7mld1iaTlMA+i2NYB5b4Iwz11uLcwaSeBUSo
TP7jaoS+8QGv+/uSDSuLDCrENcG/RTuoudp09W1CZMo20vK/Ym7urzdYZQKt
w1TaEkHYEEq8DZervbaSajKxtjV9cWJlm69Ujhn9cafDzDb/1IDd7NZZYoCm
zvLemeQs1hKGhIvLwk4B8AdyiESPKuToLVpXl7aD+/flYAKtbvzCphw0PWiA
9BgS18qBJU7IlMh8QR+HwcRHt62b279Sjfeq+s6+9Erh1fW6w7CR6Yh8OshT
kobcLnfTUtkg/q6ZmHBVJsCKR4J8XAp4+BHdE67iloNNBBD5SKg0qOIAxvm6
8M4lIBSs+MIAciyqTlIt2kjOlHvVHQFEkHwcZxy+DMprp3m2ZaSj3edUWKh3
bm/xdIxVEEax58WkZ/ttGc+Xxa2j19cExIoBzRva/Jw6ARIwXPWcPg3F/vDk
/NG6eMg6fkP1gkro0yttNzN0l6jGi3rFshRY87/lKyaBels3FjVaJNPjEgAi
ODGtVIq1i9PQ0d4jHFWk3VOMNRNK0JX9+dhID2c+15czD5Y/ofibpJ5Reo5l
ljxEYVQfQ7BYJJlIrPyw1TGxXVnTS7VcUV+ZFp+QJ5NC7dHltsIY4YuYir0M
zCumyx8Q3+RA+nAFU123DXK95+f3ZbMSlqMmK9TH4WUsNKFtJ6kb90fDFrTd
5VE3bUAItglGxA7VB+XutCoy04w69wjhRmFV9Ik87YfepbiA5AKd8U9v4DS0
CMoXzVJGwXtxBhaJfwvxCg7px8b3x1ApLwcmXnyCBiH+PwNfd/TGyZaLq4B6
jKqQN6QzUULeRLgEFGjkwtFIR+YXbPdRijx+WkyWDuL1AG/hlJDK+4PvFJMd
rmD/LrLUjSx2lDPA59jUTgw7Q6NHbNZnJfhaLSzVl4EsdAmmd9eBY0fVQuWL
Tt1VOwj3brVUcLlMbGlDTt0R5ul+bysCodRNbDfybB3OU05EHJLh+fr2qX1M
duHLqmffzByTmxATP9cciMDQFBQrV/w3ORMuzHFRhfw2Y+hnt6XNlEFMwtzs
wBNpWC2Z19npFkknwCqsIvrJdoVgX2ZQpMY8A2McJHbG6y5v9xGXaeG++uJT
MVYEjK9joZAZLKtR0eVtWp3dLf0lDhEs09QoRxrqa5eZPzUuReRq1VC0jPmB
laIW92VVpCqBxpjrjk5sixrFjr1WQCHG2tILrWtuGT34QYHSDIxWaaQ2C15W
CZD16ICioGinDPno6tzQTwm/NcH8qH3YWQmsdnRxiai3aVqqqVxQQs3z2RuZ
RB/YmonitFAc+cUa+YpPBZg3wQ9RzjaGLbCSRuDGXwFpj/KMtqEaD/kDzNDc
77yx6NcfmCm8dlIYSI5ydXQLxZQONAIUDeSdfYp//6HZ6PzNZOUk7H0T3m/D
xN8uwGeLAdDJeCrwoFCU3i9M9cOSoP177Po6whLlCsg9vJnsr9c8nVZJKY0y
R5QVrXIJ/w7vyWt3CfsZBh3lrR8PfvCuN3yh/4Q//9X0WuAR4SPdpROsaWJw
e/eWLlu7kF92rFoMBCe4FkIoCHPMSjTOUoW/gY6vWZkw7YxqbQTOFeYoK+0z
e75Z7/d6/a6JTQ2futPnmjZjIRitEoaZ4x8pJVKT0+xVsOB/bjaZ/Zh1Mi6E
MF8tp+9ImAR6mcaB1tF6hpsB3QaamlEqkrQoEycrtgIrm0RP563NXREjkg8C
KDE9ujsbYjx7KXhKchyWpTRXcPfVhuyFjiiMNR5BB9vl6xmf0LXCxBCgFmXT
DauyDHMYuVmVjcdRoeAICPCz+b0zVsW34Ad6nyIS6tzFTz+T2dyPJGeWamYM
DTM06RT1f4Midv4yE+GT43a+y1XKlNtUToyeMu7kuQuZM4NFNkGru5nH53Ug
8QzJ/6M8vjJHCM1CqaqXr/4tTqws90xSKjfkdsReWhffUJ8fD3gmbE/pzhJl
vTPe+3oVpA0niEdHex54ab/y8NsYCmvZ9Ep7FGtqaFSqUOQxq/I7Im16Jk8m
HsQod1qrx8Ze7ymK3xpOdTxZoy9Hka+K1cnGB/udGtRVDgT+07EDbu5JCC8k
W65LDnTAa+kyRtKnhDRHm45+SM2vm93mnFN25jWdtXVrbSdoyiyeovcFDggD
YXdaRQXOsBdsyBL+i6Wn2rK6eKt3O5x7r7bocodd85EeCQ9Cis1GZBxRBoVk
ebY8gpQb7Sjx+j6NpOoyJ8iycU+FPykiXY33oBAytZtL3anziGwVhgmyUxVP
AS6qkhjXtMB+xb/CAqMGaerGs+HgG+zIuiYWmIyATK0TcVr6jvpXQKxn1hHH
0IKV1U2DTf2+h1L44lMaScqNie+OXJq66frOKPG//O2YTT5URP/eZPcBLzei
DHuX4KP5wVnrywEOR6ly5BPQW9vQqh3A8WezffFRdJDWDlTIF9OiCrb3Kvy8
VptCeOA8Nit87jEBs5s7gwh7Qrse55Jtpq29C/oS8NWkDoH2tktOwSu13YvW
2AkiR9dSg81GdxPKWDRWjrspIIEQ12K9RJ7EvAhZSLW3j41wD0y2S703nmFr
Y6ng68dRvy6+ZAz5FkCEVhVgym+jRLizfXjltyxzY4TTnZYPIoJT+h04GtiU
EQ9qvvtJ957s0149r47d8cp8YGb4LkjlViPc/1PnNZV9XwJrnH2wKMlvmgsV
GbvE3GQEDscADW0cF5d4yBYGu0vGfoASakx0au42Ra7kJbC42SoSQsOkoWVI
g+LyqjBCPpfptqUjHAYwi/VCyesT1ezBJpmJt9ixZmk+KRXjTkC2Q3ZfYPNQ
FVqO0AVJtXa9slISW3m7d2+hFbjm3v4G0mmujwepWFIKBHOAYYPseYyD1AG3
7lSHilsokpRAHWnT4XHpBh+sIEfzozafr7M2Vsf7Bzmic7qt9xjOBvwRh2rg
GZfG1+2XQgWJ2Sy5DkFcDuyLwmAvEqsLCVgNhT35S4sVpsZezgob1Tghj9Vj
B3wdC+ydpD4EWLS2X3DBFKGl3QMNMGugeTC6aGuc7eShJQOSPAqAw7taAssk
YtLIDkVhustG/ykh1ag3NBfhPrRfmfR5A7vuSXDTXZZZsvFeYXPcFPjxGTOp
OBjkQzS38HgTynb5FRXjq27Zz9k65BA3Zv99e+mhZtfvxU39Iq3XiaSss3sr
rv+sZXrWysWS6LycKK+bkeTai8sO/PdH8Mkup4EzaJ2jsP47fcmDX8bc0PV8
6UP8zcxZ5wUnodJQYSAnA8KpM6ugq/K+uqpWL5QLkxIPvL3V4kZMqK/2Vy26
dqc9SL3bmps2M9DExRIrFSYZAPnwOTu7u/Q/kqCsCEwxhNgqYcDoj8TOzv1B
DcANWuHCExwkQvwUmPP7eBxZQpVBuT8yg9Q1Y+Pa8arDi69Z+5HWMz3icH6I
V29BSW9TCLqg2iOovpU6aTAYDT6IarHoncBfen6kpBRNOkfHtGMFNwkbzMfY
MjZxa0nC+LYcW+EUPPp642KpgSg+rVUN4h3ehx3GbM5caBTYV0PYK25BuxCJ
akMLoeWxH9NY7G1j2QsxYMC66QSCgnUf7YRtGBkYnx3WhvAHQOkEwuOo4c+X
rjTvYf/HuJp5sxn2o8+ISd/nnRxdYSYDq9W/Mm2xPPUaqUf1bTlYOvTtX/0G
QIhVtkfWYoF5sI7d4VK0Gwe+WtfhlUV48D+x+fj8mopbQ0oV6sJ9PINgqaUq
lNr4rvUnC4ezDrU9k+AORadfqpFvEeLUQBLN9W8sVTQH9IdMVxsls/dhPTC5
Nph8eKXjenCb2dGHo8azIkoypEUCLy6rPexzuzBhCzv6iyenTmJYMmbHzvyI
jMuHGesEZA4wb++rK1AIxyu4MKjAY2ZtTDAQFkfny5VutVUBj69fGrO5KpTK
j6QKsXVF4XbeqZc+lvrHCXw5wIMQmU1z2BgfzipxZcQapfUAqzFVVI3zpDhe
FL1EHfHtXz6HqB4rI/6IxPk7aUuGqxuQno6toGLbmmtySUCWO3Nnh1/8OXxL
mIEJkwhGpj3Xd24/h5go8MNeYRhXUJNbU8zbOZ0nogQj1oGT4FvMHDBtD2IM
ZWF9ADv+D+jUoDma0TLRtpT2ivMZuTFhYMj75JQV3ELvbrPlttc0vwbK+NhV
hdNifLNgcbi9r/6IYBP0XpX6PGkDmKON7t9OMnzKygvlKAmJtNXTYnDNwzt3
5vG8jE4iX1IBzK7cCJuFd67HlvQJFuN4D8Gwga3CP+LL3SKy/w6Kaaac7BV/
zGjAs6lP/fnDoc7gxptJmDTS0PalwJCyCDDLs0U6MuTtE7yjbDPfPmasNOUi
yh1RBthKTMsUY4vhAwVup/jU1iaC8WXjhfUfhow0PTuDosZ1BB6/Ab7KpsOx
Kk/MTk5lTcdUGdaZaRuckX7BCFaH/1StVda0CrNngw+sMjo3aFHOyjlnjjg+
0y4bLYWX0eEqOIcyej6Gmbb3Lwkj9h+Ilha2WDJr1A35JI1y3CHunEGaVxs9
6sreBbLVmwKQfGysNV/+vCmbDJrGtHSt5XPBq+C7x3j4eJ52mwppKPFF3mWJ
O0umyg32nnHKPQeichpYDI25M+Z1G47nKroNLNwyQqLYaTZ1QdnHr/9txc26
hWcmbk8s+M3xB2hyTqyxzt5mC8iHqCe8DuNUCh49e0oUbRIDh8uWm5mqi2fA
//FUjDtUsMr2YlBsjY0JF9hP/KjuH2GaHh/HzXSf/Sng8ozPJ6ZvkZ+Ikmum
T3nsVGyJUGN8kqbK1/hlOPBtiB78KSBBNkSMg0JpXy3lGDlWSofPsozG4J4j
1hkemlTkOxx54zMw6QohtKXjjPbZvArXShfwdG8pRcKyZJwRozMx2ytzssBi
VP5MfZhsNXlRYtLkV1EpAXSUSNwYHHGHQoStjDcwhfTcecI2y01yM9uruLyI
+ni242CSz/d3S2LHtWBAQVzgzkqksjN8WuQtjtG2UVqF+HIeIY1p4Wc2E6V3
LQ3DI7Jv0pL8hfJe8wknKnjaT5RnUGi/yAsehqL2rOBZ+oFevJH/FASkNgOS
iQP0+TyZxcke59OSLpIsJhd5lY+tDk9lPMapSZ1NCk35VAkJzL2Mpr7E/AcV
IBNqadte43Uyt7xdWaivf+h44aPqJug7nbUvQ/DGP0J760igesqhjWHKEsSV
09bW6FIqZp4qoExFuLLsqLx8R6NXC2ulTHs3qQq4/LtK8OK3/PQDMCWak1R2
9HS8ow2BSJQJRkEj21HyX843eb+Hy5E3U37COFnrm4obfRJ/yngYKOj/jM6M
XkZneihONrH00AWjY2tLeSEMBA/bOaB7QZxtXkFYBu8BKtGUpaF+ThRLUMED
yDSpg3wugWvaGV/amoxYCjQk9uFRxyHz7IijwxUluFxk8/Z4xFN5KI5plbMW
n+oV+Ja/bDXxsfyK6IDdpWA7iNOirvIz3WCL1vMKMOkUIf1Hy+KalobJJ5IA
S9RmFQviOlxwev0gCO+KLG4AIr981C6vhWydWLuEdurPYJpoJuYEKAzmz+iZ
SjcJ9M+PPlycd+5XHy5mUMH0H6m3DXk7rQSGymSDsqWERFCRDKXWA4+iqktZ
WlYMGEEtXhToZIqTBU/0cVDsSccWGK/Ea816CswyQjgG4heijiA88Ql0gfFC
peAmFr2mJv6izwH8IC6/9IAX6hDz12DkVRAG6Tl9AygrdnVFU4/RThL+5LA5
op1MdsXs1j7s91Oe28zEkMSXml/Cno147KbBqvfxU1HylGJdAgN24XerI0GE
GEMpes+vL9bUqsNzttx1Q3d3HYXSsNDJy3KTzdBkzPDsbY1aZsWe1HTOHdkB
2PzMmmONeCPshgeIqjc10dZF5sTSRvDAQX3zYXR3QCpFqJwVNPfVuv5e9FLm
P7giRPJAIX15R/ra0o+VFKSLNUf2+K3Bhd5x9yzT3p25mZKrOCkIFnmqhPBb
HtmH4MpcyKhBk8hTXMTN5M9p3b9eltvSLhN8o6fTroUxX2Xmzh2KWVJd2U86
3unUaAiJRxAX2ilJS5G9uv1F5SoR3QfxStqpwp4lYIa/JfVWYDfr0mnFg69c
p/CqztnssvGqSJn0ddcIoNywlTxbu330n0iI86xA/fPd4KiPMU5zxUW81IoL
p/oOZgDPVdLlB7ixTT09N0C4jZmNuh3L61YMd67ZFeYhQfQY634dQQ/9mPJa
d0R63rHmn1RrBxX0vBZNlkrwP8+Ut2wTyR9K5Mwb2ltzK0Bb8O+IUpmajjE5
r9v+3fEeFB5G6YnmVsJoFhLo8pNtcMmIxpQ612+v6LVrylXxZBgq8mqCPkFS
aZW2Z/VgaXmDaxXDgKxZWFp4hQhw9RJGFjANbiYQqe5ndyvfqfLMakYI36/j
nuBQI4NccTCV8d7oTjpP0JXuLqosqep8tf1SruiPzcnoCHpGZTkxhVb8vjr/
sPG203NvdCCkS2r5xrsPBchFVc+egj2lkowqjavZQZMi22RgZ5Q6JMZWzpl4
YGLOUYeIwGr/6Gc98STCOCrRwsLbTatWGbjppCsu6LgSHnKSVfDhynh7Q+4c
Xhhjx67ulGsjXJUJ+pr1jgZMxAYSTx95g37ANOlaWBqgS4eXrT+6OiJTt4+g
Y07GLavgEoavRcO0TRtn3TrZrP/jAI6TuA8n1CpuCDadJFfEXz/L5V3TDtva
o1jRbNO6W0sTnELTiVOJpFqNm/yoGLxgmOVIhw42c0yvkQwg4Xx7i1GRAWeH
aTZnFDKEvdIt89urZyOM5c2uj9fiHrG3NcbBQWxii6MH1UR3iIkOW/u6aP+8
E1+nBIUP/+RSjjWkV+EWczBLbaw3nweCZNYlvkrOBDebWa5JJeWGZFLQqntw
EW+VRo3I5D3MY7qeTXVjpUdFwkTuYYRTaYI5OKWFmKgLL60nWUY88WUll/fQ
cE3Qajm5D+9sNT5/H/Vz5Ufz+qiQU9k6mL3ANX7aJDwf/Ual07S5Rixvdi3X
9qTgoJtNeQt+GtLg8Xv/E22lyvF/a3l//+0Fud9IdgYM6LZtrCjjagnK+0YO
irnTLLowTLy/dRXtkaiNJ/5UII+Aq7gUXwYB7eGB+PlIs/gKcyYuUhv4PDLV
bGeg1b3jh6r/wCPBIq3GXb7m7aisVFo17J7QdRWz2LaNCpWh+RAZoHEBt6v9
ud6PUjR8rBsacyGZogGGshRoewI1QNF8r3UXC4zK/MQMAFgB/Df7u0P8RHPc
UvGSzXtOKJEO6qwgE71vyeK6RluQoEOBmc4YSPTOW/6Wc19RlB07Aq6SmGYE
XngQRMJhsJtR05Vu8Jj3+Pm3B4h+n+4AqHSoCdaoeqG1lhJc9vLtP0+mS6nz
16OpXZWZt9uAyHq2k1qnWCYv7qBcV9Sj7lcIUrSa2nYj3rZuD4XdC79B4Vzj
BNzQQ6oqpMUC+1YygQurhZ1aUF8qqhH/4u80/hFYQVs/0OF6gCulcLJKQgwR
SpXbhRAzmufKy9bOpRb9PKtK/sKGy2HgDeihi7ai3v90oiqtCRrw8/JKiCkH
tqKIeWVn7nOsWuz28SL0d0wiZgh2R2F7YD3AVigMk2Yge2lSEqc1Gnuxwuv7
fdP6IDlpK5kWFmr8IOi8AxmclUHHhPeIldPNEb/USoPhMZoJibbF3GIQ1sYz
FSeZmpHZemxqtz2BmdHuPPJLXFkHbhDzabB0498EL8u2ipzBh9M4F8hoFA8r
+lqXC6SpP9C2x5cLm18otsda95xE8t5XagtLXYTvCeq8YjaZJSYzsU7CZ0to
ftNRW43ZAN+2Tu9pcY/2OMgZCtPQLH+kdJH8BmKib4n2hr7cJeQyPJZF5uD6
4roVd98XLRAY4trSxZepuVOY4W+/Wj0PKedRw95C5Xek4wQGB9rdK4Woe2WN
fZVWtuZhNAFPZG+Gbv1ghm+L8l6EcxML7jj1kzCrCsm6NlzmKVrRKeDClsvd
/kBug6Jmb3ldcYDBjf8WSQwVPT3Dx1d6PW96v/th0kCDzxh4/4MzaKGCM2vr
vgYlglsVDG69KPatqEanbQfPC8oKsmUGMVKuQsheCKcvAS2qxfd3h9d9fMbH
SoU/WxBE26YQTXscvFUOSlxH1hsMJgP6etFVrgf2g3DbMOSgAhLk7gOaGq1i
BFY8PjLyK25KQsc1qQCtvrcfxh86dzevIuhqjEzvCnGAVNzUWFYH0q/1qyfO
Ysi/boXXDQABKEDJqO/HKKlrR8rsdWqvcqhgAqxPZ4yaDQQl8rpWFVz/JhWe
55Kh1RfcNF4RiErEcozTJmVfAgVmAd4nkpM6ItiNrfTvb4P/FzsWlL14ePO6
N7KdYkTypGnRZ4guy08wa7qA9M6ZPlXzEvoMDt/re7aXHbUfXCYD3l0sfpOX
GGsMGLoctDLXLIZlHICeR+QBEGN8LtXAX0JuAJz4E2S6aHVLOTmOoek3oNKi
nuw9NtZ+BnON8L4EaR7rj4WGw5jfMWqZfDUqdaPo0srtNSgdaBGG1ca5AGw9
U15nemRQuQlLNxnoadSSFFlzXLcJZ+Zrd97Cs8MkvqSQHGE+ga9ugoQcsiP9
gO//lB0+JKrz1pplijMC8vRt98pfEU5ocymBxHa/LvcoKCeU1zOf5IgFgvgz
2z9RC3JkZxBw3L/mAioSUiEzy5sFpF2St6yQDepqFdTq4t8e8K0k/AsZn7Vb
52TSw6PzjqxwJlTVu+sHW5ntqAc1O8YA1pXlxLyDgMJSIVvNF7hBxdU5/L5P
A8JRwJc2ZecqSVVOTM4aQhdknNZck4malZlr+8JWU/R0ydy0/MqNf0P9n6mj
mncJi2QgeFMP4xkOG37sRRsDRrXzzO0DnUtt1xWh1CE9HiTZlMKCvc5b8yHk
UMsRk1Km7mqCbMqUmRIJey2LbRNxvuSZHJHovDKtHxT9/d+kakgF9I6eXOXm
QkCf94r5GmMNQasvvUiWhxn9kxjC6MDfAB+9OqoJh0i8ih4G21SARQGnYMsk
wzKWTG8gjg7uEOwb85WwpRmBUZK18aq0mMZkhGaN9SiUnk8pl7GJrSpghdb9
pE6js3t/r9EweVcdoHzPfIHGFEIyO9dOmC8bsPaUtxkdDQlQIzsHrq7I6WPg
d73BHQMl75p+AIPRN2uU8viBJZJ2uvXOW6bML8N1iD2lglra2KA/JpmSEZhl
gEb4CA2fFXX3OtCUuqVfvmM3d01U5b0HAOUmML3CKy2YK5533bRTbpVWnbRt
jjaS7Omma+eI+TRZgbO/aPCYWreYPAieZr4Gyoc6yO/HEYtaa/uDntQQypcM
Lyy/hcRZNxG+Lp1g9gqbFhXHaNtLIcC+/632FgC63Tk4+ORz3nuZut0oQKlD
hfAgZl8WC/dlwm63LmgHztQk+t8ncvKI1fxURWrbgEK+KVcxtm5gK528l7DL
Z9535KEAmkFSMxeDjwfPEJMYspzUnMZ3tciBKck9Ac3LwNJOC7wU8mLCA30I
92GgSC/aYNJcoQC3d9mKgqdCgKh/4/Qnu2bIVY8cbwLmuRHrWN2892hVQDh4
OPIk88DklqTRf1bK+fgDe/5aJehcI/CKNzuwJ8JpweyMRqbPOgJF8N+qHzm0
Y9iK+PSHuQ3yXoSLZKggujO5G3DG2A1G091Krn/voarJXUuvuYiZ0cvdQ4cJ
8vyqYns0s3sjO7wUOazhxhUOCSI2XUGRtwv29Syb3L7IetVM1zi2eFOiVN4y
uVEmek4QjUTARZEzoY9W9nzijfhpr2RTCAEqJ/znYazA2BTcCHoQmUfo3EOm
VeRM8RbaMCpk2P2OiZqEWPjWIki8mPxCGlvon0RMOnz+r3hv2TNcuF2X6xEN
gj/6fA8E+Clpvx8VtggzQtNmn//t7Ke2OUTvk0eFFJYir8qzNMMgGCHiLjZv
noeHtwwrCPqil9LN8j4Za08U12OvkAZ7kAKoCzDjC/BAGxvWm+WRVra2P5wz
0xxeYZDm20RpB7lAlA7RC6VpSQy6rjIGAtfBsReSYSPy7JK9p+dwugfENPPl
gqs9A0FxmVcwt3lLeeC+2uKAXOKfFowKXs0ztXqOBVyOMODe4jlQrqs6OY+6
V2uVPrOKibGwEgp3VJTycsPfStagELLk63XhQbQdRqBqYm3N8XUhb8M+c4By
G6jduwwu+9XuXCZqTbVr0yBzfVdr7HxMWYxgAb8WomMjJ6yakIEfocD3mmg7
9Va/n1D+Fho8fLjqsrUQUDefvfQL4NL2TFJyAHh6BzKPRpLsR52mvGIczNR+
tjAqcpgUJN32AbwFrFdUus9HNilKaihTE1t8UWJR1+Pk2xMhBYPkUqTofc62
amQT5xErfCJ6al5ELe3obh4nRpBOlUuztuPwLGBKFPpRTlFQArde1QuSqXpS
r9L+WCE9eLvlHBfL9ykYCMYMWQQHXJa0e7xOoBb+46X1s4obY9nK/hUl7xMK
PE7Wt9QVhje0CV8ZWkwmUsf+b/NzBHQvEdxq04Y3y1BmNPWSccymhWimPFWd
36Mm4NQUPqSnr7U0vcY+2D4+Nz56vIS0az5yUPleEOiXYCnjo7dN+8rNKOOt
OFicy9QiJC8909qyRaG828/qXefvR8f19Q78+paQgRZG9yoEP59ZEk8xanYF
7jFQV19Ws0iCxAcPHFoRUD7085VHe3uO7sYud7eV9EOE2irg/Ev048lBOdPp
pdCQp9xivatlcW9TNyPmhk0g4tTrdJhDqLtC07hQI3StXKYIAWmNoGZJbDk6
ixzl7SgcxIVbxT5ancVaLEmBAWKhauenGeB3JQMVGTBMsYLRxYBIL2vaVGE8
6szvCjUQWSvrquWYyTLRLag4H3Ytq+81Qmv5HpGCgkjQSk5Bist6NpCXcLwz
qTZA8QgVlEymPFl5w2S4pz6orl6o0alb57zK+YK/36POqJuUyrZkTmMLHcxI
Lt/UYC9MRwXU3aADymMxNWjnh35I9zJqp2o4VpjIurA5TaCof/Yr8XXMZeZM
O4PD4biioq4g4Mk8eR56pOb0XUbUF2B2b0gJMqIwFivqiRsbE1ZXbl+mt9UK
bEV7oc+A2kNk/X4ChwgaGu1qgU3dSKH0/nJgBAD4h6yRsdygHZlONLAxtSpN
6ljzr35ThBDMKyOqDVqViMQmUJQ8pGyKWcl+lcqEt3TRVSvxL8QuHmNknWo1
yKf+L5SbaJoci15wLvXL82VTYHT+pZaYxX5DAPP66aM2Wmu9AxR+6f7R/KZT
KTuhFMmFfjR8eDnCq5jIzgBbJLRgpnOdvRLh+fjrQuqbMI7Eze3S5/DNUrnf
0Djao5Izu3YLf6So5rrFvImN70HBY8bN84I3QDn1iQWuBzox8nItrClEgzxx
uqgQ3jL7S9boe7SiOkuhtwU7lvJ+/r34UyhYSWrKH7zTjy5IudYsXrCaW6qv
ht/D9vbM7QAR76Cb01j8FcpTec76eZnf6eAIhLQdKcYPQuyHsXbLhhDR25ca
vlcUSl9jryWl6++Oc9NLw1XDHktKJWLPZ5wOTIQ91Fg5hQt+iV0i8OpbxoJC
O1jagIXJ6OoXugmfgwf4kiPsZEHkFpsplfC5j3gNL7pQm1no1qzAwncxKZ3n
Gwn74ha+BC7s1iiP4goXZlIMmqCbRxfN4W+uZ2BaT2KB8wSpzL4jFWU2kQUc
elsD3V6ReVx7CddlMqIQ0R5nZ3YaR77A0VytsVp6r+A5lZdEVEoQJj8rWoEl
+vBxdbJjZeC2m46ueNsh3cCBd2r/2md8GmW9r+Y1PXDtcpf3kC4uqAJL3Eqz
VmroNJbazBrFDQe+Ui9ATp4OEoKBRfB7aaZm3W5rfk5YrbZaWZGo2kZ0i56d
LogOY5QUh7cbw4Zl5GcaMZUP5yYfB7zQyFXGpSLpbM0s/MxJgO3r9iy5V7GS
9PgL/kQjDEbUcWRafwIQhGwFP75ksbQu+1a7loeWgrd/84WDTJC7amx/Q7ag
lunw7GzpiuZCFeI4xrcMF2qeXhqS27ki08ZuHdNGqekAgBr2/+UPG6VNvuSK
OxZwLKcZxrXit89cFStAXwvmKg/vcg0cOTuR1qI+4QG+TP9qQygWzkyzE0Pg
sge0TIu2BnR/Jk3+5P9wSUGGBKPQlrNNSuIcBe7JIy5Gqhv+NZrHzeLVCzlA
1l42ElbSIRo9W+V6QMe6z4JMZMFonPAtb0NHozUofs77M6ZsGgvGRZBJ9DKF
P7C7Rp8x/ccSwJiPfJbSQ7RKli/ZAcEt8IY6EKIo14ODA+N+t/sQ/uZ84M6q
clyRS92MYDI9odN7QLh0ez/CaLD3dOTS/qvRoL4MtxDIfVXniTBnGIcxVPN8
mg/k4mWE/gbIyyM2szUPO8PT6suZWltUOa5So3PAM8XnnVfdfo8irs/xnNIF
+EIJEzQrDT7JzzOJrKLpkPY+hLV4JW/QNWzM86AqJZFkasA5kXvtnnS+/ej2
rrar7xjgFDnJcKTCPH9VpLpS8O0LFqxJA+C1PxOOoPjiLUSmGC5Kpz9ANI3P
gKk6sbs435WoDWrzq+1Mh1NmQgxMCCFa5yzSe5Qb0xZcjmNPJ8Za+J3s0g3z
OHTcVqsAK4ccdmbJ0DimTVwLjslCMzOLo3yP7NcoleUV5dH5Aixajg3XfdVp
GjgQaNBBPURTjZaPhkGMjn2KJl/gxn0ja4S6eAptpjLguMsRbP46y/uCFZzq
wvI+XjnPO5OzEugI7rgE2OtIH8iHgkF4aXHet33t9INdaicwAJoTGhUXQaJ9
ADkIapszIO8JbOyauDghmWdDChGYi/JvIeeFkB2Yw6hTVb4P6PZ7zC2cqG8M
GZhoOPQfcg9Fr8txLMWOtpetqDpsKH7eRENrNl8zwvszofBVeHXFro/BZt9+
T9ypPFA3kw05b/st0q0zoRt3eXPmTiHv8N0Qb64b00Ilen5Dn5MU/68TAYZA
PyN+B8mmht8mykKt4fEOmFnlN4Ptl9IyIZu2t5/gR9NAF1uWUuxb9ISPkAOK
v6t9JYHzweCNqM4+WnPpxUze7bvI/rIJ9TpJqgWyVV/oAo5vp5ypoXZC6OQv
RIAhMOz2g2SauBKBlpCCxfKYG91L/H/NsrjP3Zb6zlXuecc9lRhwVPs6o5Y3
egK+g0GBtU6d5k5OY6MvteedjU+2/afcSbGlYy+SovFjzsWvq5fBhhHGshJU
c9B7km2FK0YewGZWBVemrv7OgKzaPoYoUDkEil6PEsWK8h7IFppIAjsfyTAW
WWK6uThoUm8p0/mmuwPPqHx9i7Q74IwTVv1Lr0lltJtT4FNTI7/iCxvbTqFI
wKYsQKM5CW7TP4XCVqQFa/18/8nLwC0W7epcWOWnKlTgRO+X0AuC9Q0MFNZv
cuIsLFPMtUybRJdTgvhFjz8U3EPFuD6a3PXX6zqIbWxMCROnxTNWi0aX081y
XPTmQdqWJgMGhUYFDKBhZepIzrtdYhW1UaaxD0+NBz5nhWjJar4eWkKC972q
Mcf4AM4l2Csj44OeJ3FOIG5jmBC9pr+sPNzrHNAlXnCOciqQWAUyhiBWhEvg
XQRf3zmFfOCnUsUVH6b+zbDpO4Cdb7wWi2xZz7MNZyO1A84/5438bUM2cOmT
1fHId0pO0/Dhs5n91fDxTbATiTporKGFWSrR2EUYhcvzl3uxbKVpfxUUxIGP
3oQMPNnwOveKxZI327cRpt+SnsRurVHLJ2oB1OXzrTpGdmbF66FgHcbmKnFn
V7/s6reHbRoMoXsywlrL2NhLOuOzHVeUuAninYbT4E6NfZeM6DBu6A9MkNFc
9MiS+Yn+7TmARMoZjEKJBQjPFoe2Ke8GTHaN04R0Oq7NmVslt4W74kXLqvWx
DyOVzj3AvKXclAoG+535fcI6/LxFGdbPBLDLZZjBtHH6RYSADT1MwSNPSSkr
o5rfvBRhjfNxMvbjK2+/HvJ1UHCh8FmpD3W4kQ2qOLq1Du5gi6Y6hazs9xMq
1v8AxaSGwtSfL+ixEDvcZFqKiqEe4lda9WJlAo0JDN+kjDs+RFHJFbvYfKAP
nsWDE/N4kWbvBNj/jG2PmV3F/ebcEYPC734LxXZZZG+FdEA/zi0hl2et+2v2
IboqV/JH4+3a0mEcsWFOnDHZHkkyNNyltbF5ljxQsNmb447/ichJpS9BtvTB
xwmaOvsWH2ptzy0HfrxKIpzxCQYtLyo0h9fskqPquumu75k+wlRMYzi3GpZ1
Fo0AMVZicoIZTfhbctiFtxdKxh7Mu9fcxqDrlbM724oX/KpEkT956thT426p
/6zKlRoXewwRLsqGs7gTWxBQiKBoGEh2UKsuAjMCM5ApvlnAp8SK2DJIY4Wl
usddTV64yHsFP9X1kgHcqzjp1uU0y1G8ZZlWB0B6izfxUiWKi0VQFCwMTYnh
VbHMhRR0YvvOeLCI6FB92PGq4BTZW8EiCbwOtM5u3tAZk9P8ft7hAWq8D655
CtIrBFizrYCyu6zjQFJZhTSvcajbPbumi1y1h72PuGk+t6ID1KJKrb6SrlBD
CWjsz7j9jFTV1xopNdzpIPO+JICTgrC2HrjA+YTwtJqDNYpfja1Z+qeHbnOx
vw8bE4Bakw1Y3dIgl33BkGNKXnK6/WRSBFwh5GSNJvvnEiB2Ogh8rwWrFmHJ
HFf3rhiSLDOZYVeCh3j3bW/KusmKXDK6sJa/kdhtLZsccC8BPEn+KTAeu3tH
Ta7jEjkjJpgGqO9j1mMsZz/taipuw0JwbNivTM4M3bLk3zH0kv95GD/qCLr9
ARhnlWM+Kdb9IzUHQWmkjWVwuWqsxFxYLOsdVP184+/o2lLbditF6TTSZ1LU
zMVRxc60ERAleNNHz06VotVAQzFuT7GGlzt0e88HJRGWuKBZk9A5WGt64qiA
/D7SPotBD6YRVqXanzdmC7kDkMt+u7jrBND37qh7sO4JshhCDHXpgQfw0LlX
rkFb+M5L4Bdnvnhi/VgFzqP0O5kxkO8kjkY4Ib8rnCLpsj4kvrL9Nmdnn/Ba
lQjtIAjsoVsqgJJ2PaMUobOYvi8tpun0lSdZ7+651zYKsJ0XzBkL3U1qe6wm
zz/Ru+dwjIHcy07ZSJ/7q8QzkkCy2GP+B1oOrdD9wKctwoGM6Ko/G3iajlQX
FknhCQZz4miC08eVmcJ+nKn/E8XuMPBi6NKIjazxMTJ1LuZfuJq9szm/6IZv
edtMX2TduifnDmcVZai0rGnmw7TuwSvUU2X4UcV5z3t88kcJ/E45z56JY6Ls
fLVA0MLZ1RvkhLBviJrOIGjJ6hnJ3SvRqFDF2+fjwpwKd7Hwh95Ow6bv13sy
5tTaBq+Ld0gY83DRbPRVLAVmLDxuLiX9x9CKGZ+upOMzQ1qrzqEpfGqSBNWu
RsT2l0XdwJsrwRPYswss6oQiwL1QAldV0alqsUZmL5tGvJ2zFrZY+ns3E0IH
9sweYDsLBAwKZTsYKV0JT/Og66Vga2PyrnzST0hwrW4c+Dtw2BaLLVPB3yXv
xxMuveey6MDc2xIqKEgYVs4M1hNQUM+LIgGSIMfSgSTNYnP1UonSZcLIBhwg
tZt1WJDmpsMBfHAIyVJ82rjWkd1rqDAN8ezx4bG6KPiF8731yZ4AF8YV6tp3
S9i5b1pJb9KreknPnXt/wBl1lrNo/XE14r1qJWxMgXae1PG3k1BZ/735X3+Q
mXkIfkXNIh9hu7tYjF7x1VzcV71peaqTlOXKRo1G/CuhtrNaop5wvx7oXEwB
9n4UayDemsdTj2C/M6q29AVuR2FEyhN811CfBQufLsdv30miw1jTtBCuWD5e
kHKIyJfFDHgkCGDlHR09BCn/UfSQvyjsyqSLRczHoVzkTpFjljmPAaDDRi65
T0W2X/moqTdDGl+cUGnIgHFnExpPAKuR+YiRMDAjE4aeqB4PnBlxWcCNbSkx
gArBmLzBLsnatQ67ak/GDY6eRfJUbFiKZZ+SeGb6zlHTdPrgHT0SUBx+BGir
N3uz0MyM78J0G5xSXbzPWOtuTKTh60sr7L0+bjsr/g6dZR05Rv8RIuPh/+/B
ZyKbqMaGu4ST/QwqDtbYzYmgc/qgoquerI8MXufwU1sBUR9Afr48DIBXQCCm
jNx2tY545vuQfp9IjcHxYVaS9w2dvoZPtt4gwY0MLIaqsoS2Gls3ANuZxcDl
UQ2JIZNuqlwEY4RAyW64mwtkpDL18xi3KP+HoISyRVH5uNi8xhn4Er77CL8h
Bfxjl8afb8a/qW3tqdMaR6LAer29bKWSCWdmrNT5o0fQXDh83hdVIPR1Ul66
ldbCmMy83LvFDRRkNc117LKBbIJmj6f1dDOt98IiO6ADA386V09Ydz+zYpVu
11qBcB77/ZNEVP1vmpwy6S+kO4MbCij7aIQOIhbYYLzLFQS3FFy7N/VdSeD1
Y749j+o2I7XeFcB+vrtxaT9AYom7bOTrU2/YzTYkxDv6lOoGU863ScQpotgF
eIBsFkpU1Oric7dbiOXCH/yCcohDfh7xuVRkeA9Fn5nYrvt+9MWftdniFqdD
n9DHGbX0nrG9NnSXncAci5BqTUOmIXwAbD5x/ISZjk+uK886y0jpwskpFgNd
6QL0a60u5jgiN87aXLalWNnEolfIOAUjQqh4BNud8+hnwyeoCHsxF0lJrgrU
IGGFXdxXVWf60QLT6nj2DAauImN5OPDSoXm4tw98HFKcW1hSU1+EWqPXpKjU
8QJdxwS/Ol+ATqpcnfDzKrBE4wPIL4mPe3Zb9Cd58C1ecE5ebfE7im2P6SHi
ipCO4kG4CziKqnUN40C2qP/WamdktcZq99jsHBJYzFPAlRo7h8Y7HqZKmxu1
UBsBWiKWYnvzeo2izuDVuo/mn9fhP3x6kF6rusUYdEWYeGMeb+A2lMxAtDKP
XYiRCc8+1DMHEH3z7d8bbgQeHB7qieBrfywN3aLBlGxnZMtIjvCz6S1xljIZ
bV33wgzGiZkVXQlej7ktOUQ8/ZsMVlflsSmVR91jhQ1GSlntdqh+YlvdNhGd
zBP0dBEOVPciqmDiEmQFjknnmM/HMP6qHEf2L3V2B8n0KFOoD/XziydS4tio
yEVx1ctfYJqZpp1DHZPPb/jEh6KJPV4Q+SDv/kiwfiXWw/XXXd8gh2NfIRSQ
tGjMgCT+jppef1iAaczcB2tTxOnVizaztVYpsqek5r5uSzoZQXneaMvcm1rv
LmKUbyBrtucdqpvjOvaKm7obo4VADyBqAJI2ALrsTn6TGtimLxOLz4sDTAZY
5sSllWB8eVjtWmvBSzl+V33CIW5kqRhTGoKjC7qoOLY1ikkP68qQ/X07b1gG
zYS6qgsbH0pwO12JJGjKHjdILRIsff7d4Hnuz8/yjk6UMwGtJxg0gkLowQ91
Y4JcFuAteJfZjupm3Qf8IgCX4bOa8UY6+1ySWpDFnXo/K2DF+4gSunzRi1pl
w7+zEC+vvNH/WIT2pyCA3hb3dPlacGof+3BpSdvgmZbXgnOLRgH8Cj6a7iNY
2KURjYZabPxbJs4bZ31Fp2UBpxsr+aCw8rzbMRUTjA38bOm7NYyjs2PwGjJL
ZtMLvQ260ePuC5M6uMCHIVJjexZoJ/4oKMaZYSdToFOtS2fz3/sHOhsnECIh
/CFH5ldeImaxQZdtmXChrKqaWQ9OBDvQxnCbpDkVebsHo2cNEebkJ4xvyLDL
0XGULCN5ONWIDtYOQdJig+cYP0Tg7Rtk5sxQQMtrtqPMrQsnH+HT9iky7LNc
3OUA27rIwKdgKNCeXwtvX0nzmTM9DoxWew5/W9ESxWE3sWestTha0wZjD0C+
SRl0Yq0X0Jtb8U9tK4n1hp1imjPW/+ucmW7fQrh3t/1PjWGCkUld+iNd0tbm
3Rc32Obw89a9b/WuZPfp2s1QwVLiQ7nRKOnPwvccnBMo0/cictbyMDaBWdOf
C3m3v8z8uhdtaYohLQlLX/Th+nbhG00sd+Tj/+TXb5b4srjQUz7hB9VFH142
op5xqBaaH6Gz0/UIJTv9Z5408Dfwm/5zt1heFH07wS4xS8is/RigAVvyT8lT
q0TUMFshyaEw++wZTXgmZh4VJlss62pQrjaEG7sU3Zc79bFCwE2AbhDX5BUv
Grrvop6S6lnHsULu7x376USxs+j5gqZFN16jczrxMaXeBzR8FGOQI4mSKtmF
/pJ9bxmEGerrZh6lEaCp2YxctOi559pXJVt7RqZuBh4BKnbfPgsNmHwkl6Gd
A/E8ubIEsZUKon+7eApKs6r8xtyhniijNCurnanxvcFZ+SUTh+cyqDSAaICP
h8xs9tZS0ZbsEZg9sg3Tv7quEBH6Sgrb04zw3vxPAijWUyD3JF1XdBRAH4ga
aImgxNtGnr3V+OmBqsLBGS3CSyjuuMiSpWU7wnEWcthNbh0AluzdSmXBmOmJ
k41rQ4wHFwz7wOUGY0Nk14PKf8popv1bFYoXlYeG9qOM6AGMPZdeVvGTZ2qY
IhjP5bqcZESnmpkDDpAfoJIYSauoQM0bWq/Ug0bUAe41ZS7F+FLSOvyGHqVv
Oe8gcOhcQl98LtuXtHSLURPluIgHkBNygtBuHfQPdxEALOcVv9Z5j/6QiVtR
KBjinIkw+3/2KB8SXYuahdZVKPIY876cdwpDGyh7Cd4a5Z5oKCuvN7cMeXcw
5ynzT7vT1dxMS4cso6lD27B9Ooz+S9cS+8z434bKUo3E0lQ7RZledyN6CzC7
Wo7g9KS5zZhE+iICoZkHXikbb1XzkZIvmhsstta+hW8+1l4tJrsKDoQvVgRn
zZxOaj8iW3eO0l/1kB6yDHYDzRfqwzzW7eFGDAnDAHpZudG5TGHp9SX7oIzW
s0aHscQAgJDS8lfpPtNQSpkFt4MBv+GEK0M9Wrd9my9+JsmTR//wzMbORcwd
Fn8RsBDledNTi/4kjIKvDLznaiyky6Ov4j9ZM5sIcWklbUbRBqaZVuZXcy6t
wmRNCPs3FqMkMFI2+6VAA9d9dXovkDAlL/gPimc4JWhWjuCGjYi8WdBcLE+z
sVK/WMLsAw/xVqwXewq27sL2wO12cv5cdIItoQJNvjlMwYspYATEiuix+um0
o4sYM3KESf2CmmCTrJbTR40fwBu+syFaDGcd2kFPJBuj4LpVXz2dmWrl7v7m
NtEEeJibpqLBm064Ofe9c93ZLXtjdE2a3l/ydEoR9HKLt7lI7peEJ7tyuKXG
N+zfPrD9/m0hr+WIB2fhyKJz88k8E2k7MPFRvqnjqnp/6S78NqnhUvZZxeEw
Urc8uLddAZjlOAMCtq3Zeq8CxYQyVBxTlOI4pmD1E5oR+gvkqCpuKawl1dEv
1I7rVLcw2lLAskZ+3Zx6X+f06fx+4sbbv+eXKTATw3aQRpr4ayir8pGRElO0
WJMnKxLpVtX1NFpDqjynXsDDtxdm8J6s8lm+e62yzwg9W+JwJRCj1HFUzhRI
0Aed3cUt9GJmt28qgfgtV/e4A09gh897mOLcgl0tUz6YJfa4oLsV0fL3vOgx
qqF7Si2NZIYrgi/+qMGPJGO33Sf4XBlQ/Zky6DvFWJf283D+00FflnZ+R0l7
slOXwIgS9pLbagTn9pgjVHKE3uvXi/eKuBBLA2PlmaIlQZIDENbc8Te95VzX
DalIrtTSXf0iB0oD8K353zAP2+mQ5UNIB5a6/dPgBcxG367GiviL5iaUUytA
6MhqN4MLsTRUb7ERReIzHl2vqAxCZCUFAo5efeoIXHlXVIzGHJwJ9SmaUMB1
hNievbyNDiBjkqRJ0B8Gp8qVkwRTJkixYY2Wo7isBMj1/LJ3ZU1bN2Mc2tyE
N5SmaQLhdfiPS0WlNlZyglv1qFs1EO6dc+oVojnmH7QcLY2e5vLY3sgx7q7T
O3qXSbDV8tbzlQNT3kqdwP5wpxjOU8C4eA7k6+xCxIVfRH8ySGsDEsdlvd3X
8F/rRV5p/lpEuC3bllehmMBMXH81/Mf9p2eDvklZ+qv9pqrW3eUhDUnTR8xJ
IyeQeTw9m8O82XD0mkYYt8wpNZ6Lv3YTuJw/0kx2BIGBCZSULDNV1jArMW3Q
OwzQ9KoR2ijrxwP8oqqEs5vUM4t9TfgJtk5yKG7dS+Y14rf2YNz5dObH2yVy
Dm93Z8Roaf4zEYqY2uzO+LIGjpwh0Z88eZr+XBDiQwfpt3NtWnOROoM7iZTK
ef+8lMmkc/2HnbTbZl1mTnwEd9QMe/MUb6xd+LBHR5KMtb1ROCzo8+ckNLUi
Cj2GnaNoIu2oiIwbgtI1gm0O0LWoHeqNIv9p/8eoOmhyYn75gSDgHqR/sak9
O9jdkJl5H42tU7WT9eZ5ONod9QlVX9px18GuThylEUAXUeQHPPj9QedDWMhm
gXYvwc7HVe2Mw+Eh9IPaqun9ek75vFm9F5avuCD/75Twn7x1sd6AwMk+FlER
zkel1LBQH/7o1//dBKplDcv1UhinJKGhiG50iAzSM8yGbjm3lEJ0GMhRSCSs
sYa8mRVTEnxbH++oq7HQsJEnWHaXMajvHaPfpfyVZ4ewmyUj7M1ahrMqzOyV
HTWc4/zl1UsLOoRoTkntwG+9hxMP2ElL+CO0rbymy7mB/0/OO37sI6zUBt2x
+zKa+ziPndZXiycqMcNek3ikkIQJu4jlAyLMhGK76mJ2e2zkAmwN1wIYOry4
20QvruphcEeXCmIc9k0b1cp597JLY3GfGPWdLAMObFm/5SvVYCrds7bfewgz
dnA8vvLokIA9qTw6MzZlTnapcvvyvFMEDyxL1u3qaSXopvxwQMYhrplFhq2m
JrGZrLH6LGZ1Lp4Q5TNgCsAzEZD9/8CiAYKBYFyO8biTPeMU0EryAEMq0r6z
8P8g/eabp2rV8Be+HyAOgBNXNE40G275lKZkGqrW+r5gswdtSzoguDQu3BIn
W/gqEgSxz9y3zbL4hXiRnNb6+2nIsLx0dOWmqZHP/77w/C/Xu3ov65kGyMlx
zseriMxHnMTtz1F2erOoFu+K5BXZ1xk2M6oQKEkoVrhM5uU+IvffX6i2fK82
Co2/9vlrUNlozKzGpRTGhBVuyvuBKViiF42DAWTRAjkvZwB+YDIfECtLz9Cc
EKTwomqGpLj+a5Qgf79XITITsMh6Kh3040ZIF7VFxlSLBoZlfAo1zsURqBfk
LlOtgVdAdJf4q3hl2JJjxgHdwLNv4HPz1BZMKNegVLQVMfuCOFptYnuXx4QN
gwe1J5Q5JSX49lFzWA0QBJ71k95r7V5amsaTlu7YvJTe/a5nv95TQ+WUgXwY
eNKPLDPV3vppKzRwBdf7jBx0jwc3vmXKU0GLHBM5pXzlqppsmd2jgL6QYDAS
XxUcbdO2Gux0+470RGkC8HS7VHc+Q9H7Ebv0Fr9eVYtHnGPilbU3mtZW2SIz
OyEWrHFAABY5S7K2QwXDaoCNm9C6zPw73cNFDbR9SMtc52uKM0+kaK4v5tN+
qqDCxz9gfReOqfQ/pPXzz1p16f0zWi1eWTxXjRwGF3Z2eH+MxSciYMG0TFZ+
haVGlQUot7hdCl+USfoEfxC2NzW/fGiwD7TMgZvz1Me/8X3QVMs2Xt66KpOR
HFKZ76WdiAFwQOyim8ijObwoDEb2tN7XHd20SPht47p6CRmK3a46aixIOwK7
tzkf1RFfbcTftbea7RW+lQTZpGSRMt1n7cQQUuAbdzKijXlw/mHf0uH5AGZ3
F8PU0EiOdoCT0+AiItKS0l0l4plctxqQGHydWLK1rXOGoSQ3r6FSDVXhr8nF
/cqdvdMGjuj9gd0MNH4xibmmOXXOBj5T6G0MZgjnTVy02W+m4MxZGuLG3jmE
ucA6sovSqtRYHZxygO+Abti8+gAtAlPQexkvHGycLiSNJ5VXSaF+yjdm+K8g
AiTdnvi4LMRU5caYOQBcCcZzOWBr2zf9GL2RucOOCs+v2fmLD3SGD/I2xkwS
I1ikjcmjPzT8b+V6ePuQ094lUIkkMmvpMSAcgnQ/0BcKQ1xoxeXdxlnHb0Nl
XqKn5y5cZvmpo4j+nBovcT+Xam1aB3AY/Dzl8bT5W07O3IfEc9HKivx5nChH
APUJfzcl41moVLYyExN/PElB45SQsG/gPzZWkNU1cFB64bzA8QDr46V8mE82
pKUGVQFPjpfdG+9ItkFXRDD+EDpg3UmYvRK9C57wuO22ovph2zgBS1KbBMJR
XlFhV1NW+k759iCmFoRG52+kB72Ivm1f0RcCB4gHYHCq8i9EB2UfGm2jfXxL
3/77XeLiRcmlwwcyDaOnOonG3wdZ8Yr/Dj0pjfukSIzDDIXr1x5paBTo4xss
+iaUWY2bQZtfFaSqwh3crDCYIg615mBWASSJDn49n+x9d151hinaAmzvaKbg
j/ijO4d22TDdDnX9/IYZeiPQd+2veeO7teetYfV8gtGIpY+ETj6Yn2v+t9Ql
KGSgtgbtonJWNUhuDESwtlycGLa7OiKfF3miTU1bqYaKjplS9K9+7pthX35O
6P6O9wd50ENaqknOdJNtXN60MZNScDu1edCIKZncI7QJV6VKZXoe71iLmwei
+cor6PbEOgDyCzddYOmUhNxw4hUdaMorfkQ2SJQx6CCcFI1Gkr59s5NQXdGq
rSmwPu4/1s16nwh3zFWIn29MNRTDs0z0e1eNsbPGBFpBs/UpbcQaI6HnFCiI
+6F8h7XEXimYNs2zcWAhLOIHZFa1IYFNylDkwWXvQvKKa+JbhV28S0bFqNnc
6J7W5Q5SerG3UvX+4ppgIfK2Ct/K6nR61cYbx62W4/B5hTI2+yuD5vyypWt4
T5NRUv0jDMyDGkOpK3/9G6JVoxRyJp1mY170XKd1k3Z44At74tU34+xdqxzK
vHaP9nRXQrtBnySQMe2vQmV9lggA3WOI7CeIcD92vfNZQ8yFpXj43IxehjIH
lkYqM3XpiHLupKYYCTgmm+swM6HUwH2Fx2agYcK61Z5+bN9Bdzmyf5wpT0Z9
GlLMdG0hY/83efWdN3XE3xtL3RIZ5cWdDmV4ahJVtyHugX+XXYLHdYLsMPu9
3VFHG7apdEln3FBEa72v99GY2LSgfoVxF7CLayktHhxoj6Ua+Xs7xa3ELXjQ
dVvsff6a/4K12x8Wuzm47ptIvbMhuv/7AE7a6CTsOqXrYBeBYi69PDen8x+R
QkAv1623VlTklW/4XgCa5VJy01qRs74uIKhxE4Lqq5PObuQvsGRemjJh59Lj
BFGWH7nBRWpoCh4dWRwcjHwoyJCjyA7M0kWb4deMUykwe2uK8p4Sy6onc6S9
++yW0akq8ORrzhhvQXQ9cJabhARD4tN9ht+v4WuDgT3ujHhf84LCRSGPpDGF
qLueGgeC+MYjgVf6x3ltSLWRjezanTqvU/5ewf4ACu25L4/H4v3TR9bAeLrE
iQwmLCxQyxC3l+61M2aP4uQdXLNCX9S08lA5604xB6Vu5YZkNbhnK8+NQ8W8
JkMLFmX0MjG9eoc2I0GohJGExmx9OLuLCYYKkEdcH5/QfnbdaX5tIj7rbGhV
wtRmQzfmqeuvXY1v/AUMaWz55qnnJpnRSvHIK9Ld4+Qq3HytPFz9izw3kxxv
7lqW7MJckSchklzSoEqGh7dpRmSZSiEZzS4mTzoDr2U9/rmiF9kjEV2jarr6
HyGEDf1lQv2C8JTnYKhuRIYPZF0PjgT0/KORt2yTe9d22lnlrC5jyBrPPjVo
JKf7RMeGC7NTbP2P9fn9i3TVejluGuFVsU3xqJokblmhZLTY49PO+OSRIhsj
trCWfs09ymIhwjTqa9TCj5jevDS3+NWpNee353Pp7dlyouYzCrlepAiGpeJ0
854jYdAUBJCYdJpgBSXboM6EF8z4lOOraBDbrkCinx9Be4FHs+bI5UZNlFkc
ioClbOGai/URJeg7Qy8GbnFm1Uxc+GGC0NO/6KudvHKwqI0jffPs9277ocZZ
1btUsUa3J7DtowR2cZfHv1kYpbiuSC8qNOOdBAAqZLHtGs6GgsrIb3Nm3n93
CtMkcmq43uLiNxDDMDKQZfwCK3k3r4YXP7cOsM07d5A5GLUGkWkIzPxtDPOb
Z/efsqQkYxUUHsUPX5WUDBc1czQjY1Dym2bqB15q0JO/Oy4iLJZQRe+T8ELw
RurpWRqklNLeXYi2y4hlblbtD1BNiFCj3TwSM4Abt2g65dCPEo1f7MsolVBK
X57EkehQeUL9YELknHKZMs62iUj4dNKGJjvH+2Ec5MS7/HCe4BYbDu6IryHg
Dcz8z5a6wfbMeY0ajJGiF7hJuXddY9L4GHLxesAypYjCQeH+DGCSZc3LVaru
zUeJZqdZwNBbK2O1Hfj+W6iJcOkSqE5jKtfXmJ5/gqH4ytT7v956IhZJDJP4
UFL8RacxRWjAQg8f3J9GjfM9HemMo2qbp0Hx+rSpOHYjvj0MPJAiB5qhWkFY
xTFjFolg8Ln/h8448Fo8ZBXaXxoqRhqS2edtyulOV4h1CWZasDAnoj3gyCS0
OO4qi/GuF0tn3YVq8H9tkRDMZAVyofRhCehndsy+zFOnlQHNUH99pqF9eJ7Y
eAA0a+jbd6pKbIm5n4QQizyl9xQG3MGilhUYdSY5R82JgSyLaNE/ybgGlVm7
k2uOyocKSRtQQGSjeRZRFgcrVbGr5gdx0R4kNfSFY4nZJdGFCgiWRx5BK+i+
jtT6b5qzNJL5nkDHymi9B2Qse/H8DfzFZ5je1RWzZ+v2c20Fw6HqALBOwLgF
r3nd1WQWH9wTa/bBnaTaAbz3jTA8BJFr8SjqH3Dd1z3zKUsEkQkXHz9IZgiN
nlMcbxgW0a4TXnk6fD0bukycs4yrZRVyqJYyMFK8w1AzdPObNO3wB/0oMtwH
IBv6kodkfpNcTyJEUQf0iUn7HZFvRNN9h326u3KtaIWFLbR6K3E+H4KSENy+
6CouLRBq0OLKEqafOrmAe8q8m7TcG8URN8+sZk1XmBjmJQdjrOsHMK0GUuZ5
xbXQ7egutuDaxqmFGOHxlF50h+JPGX3AzLXBL+YeGz9aSQDYRPI8azfMz6/A
v/HmW7xdG41BGHE4mgnS/GVDDrtPl8s0sAlDqApLWOXr3DAZq/Q7eOlvsUj3
6G4Xhdw7VBCL9BOwwfXpGKnDCgqHCPB743ija2LbNoc4XQYXLZIpuU6SYXeQ
j8MzmwCUWW22KJwulwbWXfDuEk6H1N11lnxrOVYYlg4VMJAlhvnZjyBi9fpP
84Z8zacUjgPWcdRlVOKgbMh3rqfg9LI8V1gW+vXnNCGe0C7LUhusFb4TKv4w
35ShUvvJ2PMyWvFFshvNak/HIF1kbAx1LNRYqwC2FiHsM6ob+CpLhtjMz2gc
BkeOgneD2Khho67E7QAZ3GCSWAKBoL8dZFm6/0aNfkZaEkDPGFdBfAdDvzZR
6xzvCFv6AUlTLnSTL2dV9aHUnmP0ygY+e7mwqCAWVmkGTwlYu0WTVbhz8oOb
eua4mqzzfsyxLQ5rTUOt9jCaBBba6tITNilb9Q6CqwD+3ubybAJokopMTZlA
4ebRpbXn85duSNESnr8kF5QEn0oHuudKk1VKptW4LWbgFYpzuboLiUhzKZH1
7/4BCaI/TFJwo5NlMoH/T1OE0Pf48GGxmkDnji3JY+LktNDI0XK1ESb5Kn6g
dTBgq9Pk4+7ZxGGULsgpWFMFU45joFypbxZcGnVHpOT58RosVUlZZXGB2WKV
tUHcCgO63LrQhIKPOIBvGtNBpxWkRwlgt/rey+FDVyE9qQdiXJuATN00w0vt
KcpkRlnOhkx/9fD68SGY62d0ZBgfP0yjfhsAghd6bqUp4nL0z8Kg8GoRyusZ
cN1azY6b8T0OMZiAMd9le0MdK7MwgrvurPhN8jk+p0+xllnj45jqvpzee+CO
UBOvR8MyzvHpslMFUIWCeT8JchZNDiJlbDGKWHFCbUU/Ao0GkFC30mEg7zqk
kmdctNj793Vic0vZG7g4KzcCFUTdTSwoPXK1Cgvgf0F/LZ7gpbb9ntXOvpEy
Cec+PqBgI6lvLwi2AbKQnbTjI20vYgxEgyBKNibcoAI/CcKZUnzIOzPEzJTI
RBLhJHyR3RfExHDyu3ByB6LLwUt2xMx6LwsI4wuuNLdtXs+d7WSTEZT6wjyK
QKcLbpF2Y/NGvhq1KartZ89l6GqiAJ0JJ5olInHPLLhngEDXmbDzlBosz3aN
YT4BWaZo+j9gdTLOUAeJQWykryda5Q5gPqQObnN5aIYhgmqXkPNg752Nhqgx
tbHLwApfDKXOLOELxy5LWYaREvtq222twr/auNI2dZTgVZebKdC/ksS4g8wW
pbeWDIwnXIdD1LHVIkE+N02p8trkxQZwg25TtZkGx5ZnF0wANmgeVbcwhP9P
z2g8gx6DY91Y6k4BGwfrnCvSRYMTFCPGwYjm5wsZZgn0XRDE9I+S19k68PVH
7+4DAO3leOhlQSN7zo66wE9scgaAUbOq1vQJf8tP7uv0dC/7HxNGbnf5qmam
7mdqw/In5x75mPp1TVoUR493VPlPArziBnRCoN2x+4i5A9C3LDbB/j7YuiCp
mBbDDlwyEYNfoxISQ1MVekSXfmfwva0T/Ys3Y0pKcKrG+9IquyxiqU+yOSex
GHDib9VcXvgLUQxbdsASOde3JlTep9p8Ksw1G8CZ/BHTaVZ6eIbxJmElpuoM
pIlZbJpCWqhAo+WL6vesiyyUKz9jLsQ1zQLOIuGB78o8ctKA9HKY7/tHO7k6
rJ3dkCZbIvyYZRtiDJj21k7YIkSiokQgfd2TdHgWNsjGeAUtxvDCi000XG3v
nmRq0xoCbS/RN+7lYR0+UOKlsg8yVORETeup1AgQYeIpT6w1KWUcQh3JSyoB
ClJJBDn1XHvWmKUPYq6J/FMaQS/ElxkgvPM6OuleC+v1/ZLfpmC3PMbJbxRV
DpzGSC7RMUhxHlQ4ULL+awfDXWNSN8vIwSSs/OuSf90QohAhirbjfgXHzaPN
jpj0LO31muD71uhCHW07CYWMfwRwnLwUWxsVcJ2J2evnEcapWQLaFKr5Ahp7
ffDLUjC0BzVo9EJR2r2d8h7xG4YuLdO8H4K6nUPE5Ao76/8W2Ga5mpz3rWEH
FVWQZvSsyUh6FKsbWKMlB7ZC8k9IqninHBwxpAeDKRVR9JAhh/L2ftK2LxPB
ab/Ln+X4zttVoPmdA9IDFs9tUP4hpaUrYNo25dUmQ2Q/1n3O4yzJ5s2NANW9
3rOLM0R8jNfWRGQpVh3SxO7j+PCeqfKzaZWfdO0+Axl4WC2I2Uk1E9FAQr7L
HEV9xzwygCBsLbmalxDLqLVxoLRuZX2b9XP+f69VZjs4KiHq0mab618ZavY5
iH+1yfvkwZ1LKzch5sqrd3McG4rCbbEWg3KUpLRuD8hFieKgFPZfEvSz9OwI
I0Fj9/kiu6IrtyvZXjmOaQq7szsUGLNfjtSCjDZHrv6q52/hN6GUHCMkuoV7
d15h78xNSt0Hn03nOuyOaTsWfhOTEaOsl93KuOS439hvSsBO244y+KahDeue
nhMxhNQcB1XNFYDys24pFyN6vwGm7XuBluj8s66hFGxbGga1zRGjxT/OIoYb
Hzl9MUE/o77iKZ39lVw2aUFeUCU/f1z8hPhd2BsUgnwtVgvSs6/4IyenTZvZ
Y/fdIdRC+s7HV5Q7grvJlKCmdHR0m0w35Wt6ris2h3n4GBjXnrot5OFnwnns
Lvs6C+CWm0qRzCLrDNsRvDLaa/u7hZ38QjkkbySgn2q3tymFySAORJ9dp86J
HxkiWTfOlzIJncZNUhCO6qdgqDKYYK/Rk3WnEBZli10SU3q+USt1+9tqAfif
sEUufQftEJ4PwW3hXMNGpmYQmT0L+Xpn8z1cNP7SlVbNd4X9gMwBSVZCc0ak
HRZL2aymrpgOHUgwbATfj+2zLjEKdqJjIm2hW+/1EEZbvTxtgzD8sqa/FM8T
HAOzQik1rnrpD+byB53e2Uy4UI/vsCFVSrEKHunB4kE09GHnH/Xnocluk1rc
XYXblE/zquIHQ076Cya2tPU8HF52qFG1lw3ixBnEHB5XWutDfr3sitfFkKQY
JbYowYW6/0r1Z4StuYvw4oJOOJ/fubC/fGo/RVewtnT3Eby/NgCMuLC/NUUJ
afYSwB4LNS7VOJoSRKXyxj1wSUkVwcJDoqbJXH6ZvD1L5fZRQm3teR+UlCp0
l4KcLj2ibIZKB5mMzNbgzHIteeB0omeFEA5NBunhz+S9Kc33zlIccUpaE93V
QXYeJNbyfgcsBgH/dwPr6ZOYnfskGSjOt9IgWQ1UY3Bg3FetSW+7TCB0C71H
dR/SfcudkBLtM+4rQOg6UIYPu3hdZe2VmjRZI571C7Es2cJIcQMtcSCFTcJm
DeL9yoSn8m05oUAEG2bQDaKu48NPk56u0ek2HnuHSjCurHm4IYo0cdofLNtV
lRY1A8hN/ou6YTxn4IwbYWsW8YfiBEMzj5O5lwfBpBp6oaOC417uvAA3B2Ue
9UhO7J/oEXQ7J4Fh8ZANP+0MrG8m1dTcu/K+YRpJCkPcW25JZ34s7tPStcjw
NHdTiU3I23ZEYGbUXRpKVA9RSyakNykes0/Or+Y3QbRe8yQx6Hd1VX0MavRL
wUZk02BGh93tDmmSt9h3nyEWktXp0KTWmBHQElqiEBjXVaybIxHcTutzQmYX
OGTws1g4wtPEi6iVKp//1E5iD2p/nmfTJeijwBNix76gsrHXSZkSrtNjzR6Y
I965T+maMiH0HiEJLS4YlUT7QBQ4/ji/jh65OLDfuVNwWK5ntuuJYB1BVqgA
1G1VR4MHCGhJh8IzrW0DZ80ZMzpUPcUlSEgBefD6t9t6+F9sBYkIb86rp90K
tetiaZb0gz2RhIf/kPntnhd3Zc/1sb+32xiaoFhqHM1Qwpd/gD0q18qbNuQG
EKpDnCyZvqPaP5jIIXyolk9vx8Nsx1QQ7ElX3+b7adBSYoJGPmL0jzSVG/+g
XVEkaS3fTewS9ZAkqd8kFl3vOMqdUFgLmyxgS07Gu2wME/FiZvz07WR4zXkf
W/HYOSbqiClgJ7IgbmYCY0TifL2xfJe7lSfFv9bPqViMQtmkI1bWDQ4ZNNSG
CeG9aAIU3ZYrVA8I7ytUn4EPtZXfllrAFbetB+UG1aCMJvgBRC/ykMwkNxAP
7l20oENTSMm4hK0OopL+20sefChj63p8WR8sMSo6u37sM3iLAueS4OEtXElr
9t5FXpmzlksjgqbYR2IpCQ8k5x/BSTSjCpA06Vu3jyWSOz3PjBStX4VEW3gn
E0WejdHkGe6RgKqE1g8+lyFdRZ+1VGus7LWMAErv2ueuhrOhl8mvnSW1H1A5
2Ra7Qh7MWxljWotXuJM2+jU+fGt+PDBspWTWhre4JDIDbzq6nNgE/Ox5Qo0a
8jpUGht9YKUyQszujJxQcOjilmPm/H6OyLqE/77Ewa/7Td7X/jIJ1vJ5CMsf
oE6y3lTp7CqGy/pmDlSH/sDRrAmGtMnVTpzREBmVkGdnywp72q8q3nDgQrQS
EF4ZZvQShdC3vYC+aRA0IUs+QfWwm6kwOlexS/myH5ecWle/yrqrk108DBDu
swYokAPB4mWj+MegMAPliGgmGc3gCYjCl3IuMpJMFMBOdoUDeqWGNQvzJfbq
hi/KjLuVXO9Wo6+CPhqd/7QFTD2PqgyNbGxOldPdO5Flq8XECDjQmnDm/G0H
SwkKrQz920ncYbvlQMXJaU+VUtT2E5dRWNyewNsf4OCn3TJqoRdKg5L3viO4
3ptBDk+25MexyaqoKH/w1Pg46MfPBRHNc0RgidWYvqT2N9W513hb/JYc1S2D
zBsA0A1qg/TWLkoTx3Wcd2Jkkvmo0Ss2utTvN9XBbkOk7SLUYbwC+Q9NMS4G
p0A1BFRf9mwFQ1VOZn6lgKLZ8kocU+PYhAQjEgvF1AIRj55D0tC/hZvn8yTG
vvYHSW02u/p06xlTUm1qOmT3alq9k1Jla2qI9PSXOmXw1dkwzmaMQ6tebL2d
+D5jf147KA6PMm27+3d81x+ZLv64UIAJ8b719h/MTS1BOCUS6Wf6xFJ7zJ5X
DiZXGRPd9/yeB3feROiUvqmx/BYjqe2k8KDc7v4vEuyZzcGZZW7GzLD5EAzP
S757fxfpurA3qPCjNsE/DsQ4t3QCk3qqKt3XCl6sHdmY5IFxAeoNwEODv+PT
kaF1q5pBlT5xhO7ymSzcMQomjRVzH4Vimm2I7CDC5fdg6V7TA4QL8gXbiKJb
VsFd2Kp/Fh2J8Jb59eK5YFgkB4087KEx/pyEkmDU+2yGmoU0Sr7CtynNymFJ
8izhejsbajh9/AxAUH7hrMwL9upH4wz7XVMJSjhNmcFvP0Qdvw4abgfLoHAM
iDXkneStRKSPP+/zw8LBZwkAOkMZi4QaWgGN+vFZj/pGHNGaR7GbwkR8b/ng
p9IJJd2xwS3oIS6BwZO42H4JsR68W37LTteqG+7ZaXK7r+ImkLZ61+mNgiG/
lMx56JbUECKiwdSbgzqGjsN8sHeb9aW7h1W5k0OzOOBvH7la9sRlHBw6V2KW
GGlfK3V1YP+OlEeA5AA5majf/7mDr987Do2Rho+QKjf2PBoVeMcMRwxD67Se
GUvZqm2CQ8ExzdKK0uE3y8VXoWQJlsQz6Jp8XiAP/Q4L0dnZ0G1tOZMjVKve
iQHbUrcTk6uf5oj3J2w3TaXmNgRo2HUcP7/JD1nMOdxL7a1wEFBQCcCPB/+E
3uHhKO5NIIF1ZVmYQ5CHWM7Fh6Jv4gKv2DAW6TmVdfC7Hw0fpxC53/B1MWNG
0VmDjpn7R/cA/JAl5lRu/4ccKyDSV5CIMx7TNztwWM+ox83U58Y7hAdkZ8qv
nwvhqy/sISbSoRwHNKZ164SmRT7fnfdA/q1h60VoZqE3OhNNMn0T6YUyKvm/
9BJb1hMiUucscweFWUk14Knox0b/cH0/PDSy/hJv0Z8x7zbuTu56s6X85xGP
GWsyPhAvBx7tAgUy+XlkY5uHrmVHF8FudbTzQb256kZo+SvEBpOXkXcSSOjT
+QGku8E6iHraWGaQtzJ2OxFfdL8YZCqZVtoe+6Va2Fai9qnv3GCz9KjgUka0
S+R7H9G8v9jqx+lvUIjOzN+ZH4sRQhsr0pestbxuezVUOBHXXofM62sRuYdc
wP4jNceeuqgLIMu4+XwwjNtXiCP2iE4bXi0EcfO0CtZXfRYm/0IJsdX1yGPH
ylRP+ZrrCDfA1SF+nLKzyLyg1g+NWQQmzJ3GJk4aFALOXkvszar/DXTtvQUt
1EB5y9tLjxYCzD3a010AGPQoQqIrG9tZ/VvRQvXVjm6F+2hPmy0ofAr8+U9C
l4ZusTsQp9WAuL9b+Vm1vTiAE4w9QekTFmgKJJ7YnZkvqMawhJImuLG4mEEM
qgFQqagvR3HKUBuIwFPiZp+4+T0Ffnxc/3mgc9kmcj8c/pEpvabSCt6Q8V2i
bqhq0zBj/va+Wo3uWGbcwr45M5cpFWhotUgmhmjojap8HX6rEI6880AY6GjJ
PXU3ToVdQu7yXNOraj6nk9/nS4hzZMpZap5rJm5SI47oS4KOpcNASd7Se3sE
Nm68wSiwNFOZHL+npsG/BrH/Uq04euKwzqFtZnIWySzYM7x8SMpw3yOyWqoy
6lvHWEpNZqErgvVhL852J9o8W6UxNt8GS1yH+aXxp/uIhPMQ/oh+CRMoqMS0
/U3H4WeHs0PHyts5JcRxY3It3v7nc7/QE5c+WK6hqeqwSqDJD3pgV9KEEEvt
PeMsH1YMHQi7cEeV+ZQdzOEREGSCEmGkaU9bNO+g/2yorMDNyqXJvzmXOFOG
MViCbheffXBSMb4M6WeOtjlX3J4x8FsduB5C5Dh4H6ed3fdGoK0wznJrSkKk
z1PGjCJ/7VID9wDqrA6CBUqRz0cTA+I24ejxFzRzN1coJSW4zmsq6/IHvlsn
rtd9vbe9SgSmzo6WMJonJM96g8P+qkVac7o61sldOEfZyYtdIT9FiYaMfIQY
cgo7/jwNN78rlAKPsIe1QQ8kS5sNW2wFjEi6ZX4sfKtVKu9WavLBrFQfJj+l
9X0jEyBf5LzBU1H+5AtepCezTlIRMei4oDfeS5Vy+4IrszJKIoUJ0vXgX5Ij
5aG1x6ieTXv7XlRqpXiqXrRNoNIDDL21LGeyJKdy2CH3yxi1JwXiXIa1N2oS
XnVe5v8KXeNQ7VfXXR5L5kRObzPQunZyLj0U4Sr34YpRRR8lO8BZ5W/95yZ1
FYEnp2CeNmuPI0jr5PBi6gzXAIa2185nhHy9WgL132GdU3QqeAxCMnaFcE5n
7os2VFoY6lG9WzY3FxDr3NWib0t672RHEfdKJyGlq4KtUUDxJRBPu5l9soB7
sv99KEpQpD5da92C7d7ZEJOediEvFr7md3vfssZ8OgU4Rw67QDdpuQs4VrNq
47tr3CyBad2paK/wzMrADZdWp6ha5aT9M+etcZ1qsLxYkXsIlR3ccnovYTDN
k8yyUU0SxsZ8vac3dEVNN/7TLMD2kd3uRvq57566JRGUUIRO3ido+YpfXz1m
F6+vmQqhhL6bb7eXBs3JNv3ziZAKCJVBqj209+qSd4HAyjy8/4hTEU0G7Tis
lfnIq31m3qer/PE04lec3usZLbp3nVeYthx/4B/SquljYGk/xFJDttwBWO4J
sWYqqjc9I71ljakgnhnrs3gQHUr2NfrS0HIe4LKgkNXgcje773oAjHuITkhS
htUkXYdOkUlS1Bru32EmIl5hlWVKScCN2JfjvtWngmBHacQEjR45n9EaWppL
U2aOWdeTnWmyPi2LXV/xu3HRs81pf9nT0+pLKoWSWMslWC0ZLKdX9kaR3fZd
7GSM+gW5zncmTS0RMUNf5MsiiOUIMTf9VRcQj7nfvu/8Tei475MmIfDqoPiN
nKQZuiEp/qDPVaKuGKYQFhD+QM6wH6eVfZJX/Ih0HQkszl0p1fHlLfSdBjR7
oxaEiZ0AuGuF/tWPpqYqGi2viUaL6n5a9Bf8PYnetUkPX+zkPMOKyTYktmMv
6ZvJp1JFLU537PM4SVOE3jMpspxIKskogF4eQ/+E2sSNB/3w9J5IhfuB4CT3
sQ6x32dgQcxhp4eQyElpRZSCRsf1ZTk25C2yZuuKS60hEDw1IXJtrFk3icAw
/4PQkM32f3gHyg501lTPAiWTMUBrRRAgUrO056oPJ3FTKnuUT4JpFOlvE9rK
kJiUmhn0XI46yhIzrh6a39minKqflRrP7klaCJyo6YDiq0ZQYL/Nxt/87ibk
xsH3zuecad8jz5pYGnXGgGSc7FgJboXeY1ooKDp2vHCDTMJvIBi+LgzXPoz6
TOth1xENrlnP6SEIw66CR0HubIYxuDwbdXZzco5sOsLfZZbDGfTmPCva9F2F
j+FWbH3KfsvX3mb6oTFD6vagShQcieTWdqjnewnmcqa3KboVlVvm32Odclxr
7jCrq1sG3ZZihusnOENh1kuLp+imf2AgJROlto5BGooMg2+qH/Ae28JCbBb0
V5klKwAnCljaIaI6yN6s/BVr3dXUAzXv+H7f57+/a3uveMiClLWlw8sc8r8s
pngnLC3m0/kqOdolnq1+aUrfOGlAuMacdi5hnY5cGh7iHrM/b/AIWwxVTReR
/mfjRGgdXccf1K7qPBxI0et+GOBLfe3v4uNS/hbxNpxeOD8pijkB5LFE4kVB
NMHHxq5eOUbcs2dgLwZEb1oRMcA7EqiPMNqdz1ldCTTQ4IUg0fYrpL2gf3jJ
/U1M5ShReLjzjRASn+iuJNSmFIWAbCxUDZWtsiu0vdN42s+v9pnOQIzy9e4h
wTkQfVUrA6k06+dWubfkZxpkxG1Ghllzoc93jSFSR+GXDIzJhoCN0k3sdjfD
Sbetei9I8TTv5RT1yjRqvkeTTT89+uj47B5N/eY2555ts7Fje7LxvmCjSkpg
3jzC+5WYSwBI2Anmh5isFtN5IOOXaJssx4vs7vlToFhiRO5nJBPddtTLhywn
6ReS/g39ESD+FaeT+p5Vgckd4qjDU1+A+KPFfX3mc+A0vupNamq7SZv0T322
/4g9b519eD2FJ0OSb6zsVjqkrp6j21Rw7W84zXtgD4Mm88luIoi82GDPImbh
H6AXH+GkhciZQF7ysKZNhbPgKxDnVPtrYZRmKSqpLINSCXFTrpx7cZahI78e
2ORRAi1w5SAmwvYndN8kRkZ5dK0gNCuXftN/UsrkoAkqlLWXfwM06wgQVAZL
dZJXu7wxLyoDpHthOtIUpKzCUgElviisD9odrhbcXzAV12+N6V3onXxTJQYj
VOZBck+0qOBomdkupse2wezbKmKXoilZD+E9QnzaOSmm3vuoM/MWLyD1jXvn
O6guHRfZwqyDvYZoPVy6AHE99cRKN9IaV2p0HnOnogW2oVPPoDiJnQZuXBlZ
623cMF6FtziXj7h63Mm7iZQpt0U7VBuydRZZccA+5lTbCCmO326ejNf5Y2ne
yidQDjdS/y4kHoelwyBlpZbdWJZNSNKeEURlduG7/DayAK+BmJ14a+tfsHyh
hH7kj2i4wOscIeSG9WBogVWnK+45ydkaWD2z+ClKhwNB9RE4uYIynzj84bFL
S+fCfAehotohxN9L/Ll74+UU0fH2WklbIkGNLcXdYb1TAZLLHZ1fJ+DV2S9D
gy3MByAAN+mLAKiF6ZsErStTGL8GBVZQkclCRSh1v/m1lgaSTRUT8jwK+Du1
9k7sPQF0hIhTtlGc+jotvraLiwSH98mjOP1C7SeoO4aoh9q01YgxsySJaaWV
zXnLU78SgKhaQVyZf64qgHPiSTp4eA07j64KmtMEx0K0WJK+DAzilkLopxu2
O3Ilw0s3PMz0OWS+HlPb6gws9V7mkTJThBy8d98zVVTzBvlDQv54xPbeVezI
iV8UYwtIB52qu5piU0bdEB8JmB1IN1xYqTKjbFhVdJnaL5FZ2Wc+X2t8+rCS
FAj//sTERMVLsWcJqfMoYc+yAWiahcg3H/9JAEfMjpROxtd3VMHvMeCe7vBG
WAiNgLG9fLDa4vFFoA4jYN5yT0KQzDUwh1WefEfN5iv2Pe+pFQedGErMxunn
HWf5xmEQuKMSUVC5jjwQDxxjEvPG5E3iuWr2P6cNbIzUsu7j86kG/cRfUERI
5/vclOwtAyPFY28Hb9GZt5AcC3bqUbBeaxJJ/uocNjzq8Q3o9h0u00CLZU5F
fb+P/d+E+Khp/pGu0GPDTrz4zhp8XYo82w029DSTgvV4Ypo/WHfteb942MNU
zhj1yPWkBQ167XugcllIvTwTZJk9NNSocm0MffL420nXTXY4VqYvbwUNEfA2
Fw1Mo7lfIig9x62AwAuT1xvS6wxeLAsx98MKmMFbTrsuXoOMiHrvcXR1TKHo
XAbbvpFuHguWtiRPWTINUxOYNrI+LmXhPARAD/C7wPF8NxMzX7qQs/fmY9aI
AbIwWwjaSLdlJNt+Sa0bxridh7jW6BEwqMlhS9+RMzjW4SWOKIXqKfUIj6Fq
hiU39UERjxyqg3IzkGObMREdMi6K0Haq0B3gnqA6Nsny14P8B4MQrRUIGkED
mmc+kr4LWoqH/dGWAABHksWKDEV4Cejk2HWmqk/nQSP7zNKHScFO1IEVA/96
Yn6Uwzl64GCXFfgQvfchH7crdKShu4i1V1xGhP0w9koOy5HpDLK5FtVoyWsi
WkDkDP6U/lgHD0qCQsKt4JL38YpPaLowoFOuMTTzpXcX3xPsrEJikvTDsBi9
CxoHhNPrVzHXGlekso9V8PbamwJwIFLImjeowRSDPreZVMqp8OM2PjAyEsHz
vnWkH2puScQCoZ0SXD7nldx9MBlDrohGKz+Bs6KPdPHnDR8oTpJdZuy8Vysk
I+o4Fin+eHzMhxJ5ki/P4zqVuY//RQTDEyMSIOrzuH5ZLOmFCF45w/50R2fl
7zochdwQFw3tMr4NDJebFDe7NkXM9OMte5xEVvwr0ou44Hw4XEJp7pjVhe+6
b2x3372qx6T+3U7umjqWYiWskjXSey/OhArZ9kLzHlElVPipISlvIQyTEl8o
ZE09lVMDf9W7tbfKjWrDDj8wB9WfLnaBs6qbPJWqmYp8P5XueNQ367PiVeJ/
Mqlmz9w48hVb3Fxua8u7QNjX7IjxTX8WH7iSiv6Ok1toIvqgyqZsPMt4zYjQ
Vinup6Ik45SvY3S/cxU/EUcFNOwYSuPxFjpg6FI+IC2CDnhvyIcqnAT1md2j
P01dUe2eS3KnBFgS9D+e0JXF19M4eGRPhxhR7p/sn93nKzl6OAQWNoPIB44N
zdth1QDvwfvUglJjKszENiElUGn1Du6wYvDkvjR7yT8loKwdHlIrM3TwyB4S
VRd7fqN9rwvlezCemXs6sbzhzCi9H1MvHcXLL0T+ZIOm4bdwXEQxuNHnLenQ
Oh+mK3hDQEjD7keW8H4s7EC4d9ZjKBi3N6Hmb5kvtt3bgwmhtfzHPxNRq0RZ
wMk0JOAn4+Py7REdfl3URS5gtm7birdCsPz2bzcThm/21XqgtAWXsiovnqE4
mgNj5LI4ba1IkBQVkjd/YQJrg7zNXndtM+Rm1UPU6MjpQPhkchmPpitbNYzt
uHk+gCl3SMJJr7hZjJ82ssLRj5u0vjjRSiOHOAlTy76pT0L2NH+x3gmNT8d5
D2VxEpE3oP6JqkOeEy5nO9BTomO5RkbKy16ELgGPt0ab9itC9iVUTw5+cYaY
hIa1EV2Gk/Tl+SqMTBgN0qmh4tx8vHPJ2YF8cdyPJMYesdRkkcuAIGE+VQ8W
nFyb2mRbmg92AjC+WwSPv/W7iDDa6ZSM03YtkUusvqqoZ36RMZLiKLOaqn+s
qiDvNv7je9IRbyXBnyxmBGosTqLn66gNCtDuM43uhXWCyCgcz/b9cmYtkv5F
fNe4pRuBaH4PSdQg5A+90w+5XExb2LyKfTBujoYNE7ZVRnUL6UgYVs+8efdO
7rBiT024cQk+2k3NqULwEG89sGVr3O2A5c2l3fLH5f0hV6COimjq3iuzkUyH
I2Ztet/K846+gF0HnWHPaTDe9eEUrFwGFFZDQBcGkxzmYV76XBTLHAGuNKv4
Ub+b6Px2TFGlqTvK6l7/1aTTroayC9uli47LV/+pWo/42/Qo1RnMXiDVB0Xk
E+SpsT5vYYofIH6aAVKX6D9clOAUIYflTzV/9tYGyXJAKQDHYKs+/gGbeRee
3ud7TJNcX8aR7CJXHjTF8QCtTdCfwCNm0VnY+r2EDrJlwpDjPoz44q38pCOX
yEYgeQJlyPpcddBpFAoNb9Q+//tX/wj0SMIIICU5Gq9XdeWGc2mHAsVlsCoa
UHYscg34OOWZlyNbcO8DRhRMn4ze/Ko5s2g4xDh6osakxpMxQK8kfzceuhb1
L2HnB14yGppD09ppzPLjshedp4gpHVbtRzyKlmV0Id0vHJggMRB63mkQWIDA
9VLgrGerutFdHlT+50Gh6nVeDBg+48Pdp7qyYxsuX5cYvEgMk5emafLzfFaF
Izb9W1jSSysfkFxAq0bOP0i28GrS9CMV+WqAZv6ofClWCsz/IPHpqRYOAkQl
e/JGwE3XFKp+C+X8SsidMX54PEwzZlitJE8SI4ga2gho5luRDc4ch8dreoBj
6XH/7NaX7xwyn3FpLRrjSlFTdAKjszL9cwvsfIF46SqGL1CRZj4L09Q1W4Gw
WvtkGRIb+efr9+Z1tJfOCU6xjkRoknQWoVpOPgiVvL2YGr7lQHWbbssk/z96
F+yjLPduURRKYEmqI9h0Xomrzl0xqJCleBTD36p9up17Wyju2CLIRhcrE3Be
gFhiFCwtvBYtIS5vghHAXrxLAs8p2AA2wvGDE+D6A6808XaxtUK5OIN2w831
u8ypPh6zrdEwBPkrnwu54Z98uHUEiseE6r8xPL0eXjjiCRbI0E3XC4AnioJ4
ev6rQJaSpdgD9jnjbve1nXIhC0hNqO85ntYhTytdcWxYGDz/L1qrv/JgHgn5
iCU2ViLbqNvYkUZVg41CIyDSpVOCAQHx5k+20M7WYy3naUf42xcVCRwEiDvv
UL0IOqyrXxQp5EBw3HVEEEMEi9or8wUP6t0OZdHUeLI37clcNUYRhsjIAYQ9
BWIxkzyh4C+1RXiGDeSiZe97sefzsqiSn4xagafjfTul1qVGSVbdhuGTa63V
BVvwXzJATyzKnf9JIFn8FSfpDDjXY8GJ9lT1XBYtI9pSEheRxecs8nUYRxTI
wY7ZvWdVwlmQIei2MJA4aHxoku3O/RxS9FWqxjiXWodjjsmaPHsjtRy5wCRD
hQ9av11ZnniLZAGSXHUiG8w1MVYduTYiaNXQjh0qzy5IrPg9DRYSMfRaau4z
1fxn8rOqQc8TE4dN8EFFcrF+Ey64SsWLDAM1XVgrI0t4KwnPRJMBaZMlYsx8
oqpJSU4pEEk2ymBEoldovZJ4BQtO4qoWp9mPXahQhPCspqjFdNcUcuyIXwDT
Y2Q8rSdVRvN9PmN0QJwtZQwlFZ4R4QPZmJOK7CGJP0Hw1xROpcQ3/nCXLepS
J0sssRJQsooWza3slBLEE4sLVD+Q6EOjY0ehRzOCQP+IwLZ2FxFwDdvRMR5n
D+f5Ohz0aXZ5gPTN+jfFy/mgukfZ4SD8OolphrJTZ4X3w5aYxtFFeiALA23E
JfmRlGcdbERL+fOR4OkLjqoVoOvx1NU9+S0SvK0R91CTY4WCIxATRv3LSjtq
Aq5hUUiQvkvG5vx90y1fvaB6hX4u6u31NtiLQpv4DvUFRg8vmG8UVFc6zBjB
hgcHxpxB01GjY2Wcis58I7b2woEfgXT3nxdAkWwi8X5PBjzUPuu4ZFwZ2wLi
Bkn+P0NeRbg2ctjJofdESqoCOgHbb+HEoKY5JV1WTLmFIbRynDhPaf0KdZ3T
DeUECWdDSeR2AIj43leN5goT2+F13OsTIbGTbW7mtGInLCjc8XYn2rzDs4c9
RCkkQEDiREhSomdyftqNgTC+o8W59BIJZjp6kZzI3J9ipr0+uB58YDwA/xvY
dcLulXGSdqF8jfardl2nfbePAZ8yghgDAXCwBVKGLf9my0y6flnzCYzpQhHY
9JSVFqEfud69bA1Tuc/dCHjTQb0zGHrXCNK+vrPaQHpw9XgBqVBiWAvuRNH9
DLvdWeBJg9tZngZa6PVtTkpD+iyo95H5Us8vHgC7APDjyslZy9EJCNungJ0f
RlO4CtReEm1hrMwMt6Y1EC7qtXg9RfYqxjf6knF32Vz/xa6uqCImfLJY7n1W
Kgmags+Xdq5557RvJJpFSaqoRwytvhhLuGex58S+HcmUcC2/e7kUMQlH53yi
YqDTc1qfpy+2K+CaC08UgGIc6uvNjwQgCbjgaiKuGTg/3pYiQZnuG+jWkNMG
BgzXtvwVJS8szq+5Ium1w64mvHFcNz/sD/74NZeNAa/n8yn23RtOowvUh5dS
5hjDF7LgBSRwq/L+H2DnsIzoOR182pzzxJY5q2ruvRNwlBfp2EycST/l8Whm
UmlIIV0LJjlRLWK8WbUVLSTJ1unawkaL3fYukVZh6U8AK1a9E8eG6VUn4wOO
++OTSDVoWFqWZI9sxsT/kXLzGKdeuumqoOMR+tyohYdV4Hf1FqopbbGbEzVB
wK/5/tgpIcoGWe8NdM54fv42/lKerdo2VtKU9bWk2Wm8GLrtg1+FNKu7R/P2
MmEQcmSDteJBSoGtvoDUXOM5kum3QLtzKiEqsPDPzTWQwNp25xnu6RKlEcb9
ZhI1I8iW1r2kFAzRzLjxayWXXqPQnwtrOHfLsQY0mnRvMvm/IW6hVkJG3Xk9
0Jffh3fmseGwykhgHxHVskhl0lB454VNC6B37nS+IDRFvzf8Q7hPEIhkPRvN
S7C3GGKYicRnr+rA36TCHXejMeTooP8MMZfzIo/qHPysUAhlJ/1/B2VAQrag
yhIxEwJPD55kzSOD791Nat5hgB+yVb/gC/WksNslSHbwVBAMPMKnB7IL+OJT
+D1fcnlIwKv0mf3tv1EPb1yXw6YRGPTU8LmHuIFJZajpesh5ZuBGZ4tatAnL
w57QL+y6hHbxS0mZD14kxR0Knmr6Q7u1F16MSNsHETeFnPNy2qnaNqmvXbRh
NHlqucxaVV1VXB1i+6fMlnSXAtPGkquq0A7Qs70MFKKJ0o8CH/fQ8FEdeQOY
qytUG5T/0l004xROsmn2B+ugEAyVfr5NsdpzLYx0iY38R0CNdaeikjP0PuW/
kGsBYDfmy6IdkPc9xPdzBGb7uniDvKeVamQYbwBgduFpkeG6B5FIjRXb0b3P
fEvYcW/O1G8+uiHwNseUxFZYi8xzqfaBugNnAzS6qlbsmnZyUiOBVR/0lq8V
jXM6UminKQf0TTVbX4RAAm0YUDrdasQhNY1NRvjW2vHCmoNewwp2GTkluav5
xzWFPD2x30hBo3Bamh7/+tpzFt2YQebgIgugue6rMpYe67BTE3qamXLzl0vk
Y/OKysB8+QHr6Hk3pBLCh0ysY5FJw+EzGj+a4DQQh5v7hnwz0lkq0hbBfWjY
YjIZfux3X/dVkwKB0m93AGse4DcmxoK7DFXv1wY8HuZeYvX28Yp21zI8/mbR
1HTvbTLfL8SZANbqsZtXm2qr2sImMSY2r7GLAc3pkPb6i72vpZ0aYAEAtul+
vJQTINJ8p+p32+0RaUc+ryxROmpwJ0zC8N3bsq9rVxQdL4NDMwhiN1tQRvMj
qQrTVmemEAydYsaNUMbB6Y9qtoWHXww2OUfhLGsoyDbY89nKtQxIL1k//1Xg
7oTf/IFmtRP0p5q196pvIURnKHy5X39Lc2cVq0EDnstYpom/OzSIdvHDMaU+
cfStCPV6VEEogYRU8Kb06pYZ+glwihHw8qRuJU5uScXua06onWPTTopN8j9B
VQmZFANYT6ru8hnFTu59DLLfw2e3PE7eP241MpWZZlZhHUf1hvHyAWmjqcan
PdZt8pGgZaYI1O1OtqCZwE/QpitXpf7jmO00eq649IV4HhnBSXx0ot4cJvKW
i8KtshxP7cGbEE9A1/LwlCsRZcj5OEaEWTNADn7BRVF7ZY9VQGjlYBV7Q/QH
MAyo/P9+k7njnV9pWCWPgccAXLX6vDkDsrI3egc4k+VC4ULTdEJjcKKRhpjU
OqY9f4yDh2f0k5JcnyJnqnhtAbTJTmEAPdJ0kiPi+KREiK8Q+ew7gGNZfxLT
qLX5HG4kZay/UJBbN2DftfxzQ6l0vzFpFJf0q1We8nzSfI6GbSW/mXm7G2kQ
EN/k/Hadd02If3smChVP4Hol9bIvpMBRGFeDaX+c3A0qDKglvUs4DLvEcqXN
MbzwMbIzKH63wfoAtb0rXWo8INmKi3YiZDpR7xTMCWh9W7D8o3WBMCiBR09j
wuYt/WZ+nAWOTXN3QnPRQFN2qai6mTzyv/95KnoLNpkPlRtsjeXhMuzJVtag
2kJrKcAqx6RDWDoSVyd/LD4XTgUvqEsLKIkfr0cDVzHaEav4Qt7LuO84rCYZ
+Pil/7jUAHOA8MSwFjjaeUTxZM2UhmFsVtAsDe/MgC7/R/H6nmqtrtItMBsg
JnKG1ZpEMTdI2uWKPh+gyKK0CLqDD/cdsK2iBjOea+wzfd9/x4gjhL1y2wQh
+1/VJuamDZlx0if5tYGjMSrliLJwuuLTvU44pKnbf7jIQCR4GbzTs/UvZUBI
wSZyD6idCK883JvhUC84FnNHzk3dO8soT1rnHk29s2GtfXqEovMsmoOUQJP2
UQgdWJh2R8lKn3VgwBXdMNOG04tiah0WxtwbrbbVal8lJ3mKLm3l4BjKNqY8
BNUIRz6tJjMQh7kCamSXGcLll3c7j9pam6H5ok+v8fHzWZR8g5O19RNVjnlR
S90BZmI/YpRUUoh/6OUnaClYEIzf5kjumakNhDBuBciUJpoYac0hlexGm/iR
/T4tcORFHnAwn+4pz446vB7rXX8I5JwDnm64nsVhJqucs4r5307wrJTUFPeE
Hl8Zwz1wsqkGId7dCgrSZ2PuG/UObbC8rHMjOTOn4pcnZS6BHKF7GQgbww8U
NRBzQ2eC+yFv5Z72COszjk4LEufZIE8p/wf+dYyHR+yABHIAmWsCwKeIdoYI
tbOTodO8++caRvVuJPCj185o9e05DxBbO82jE3ofF4nZ05GEdHPCQoaoFFC1
FvXJj5+IdSbQuDkcXYpYK2RZ9K9CxOY624XAeRocxk+Njd2yUDZAUewG2YoC
/3bf9YesmJsq4Jg3uAhUwnTTnEc3rZ8eQsr+rrsUJHkoLwhTctavQGNTvKJr
7AsnWbUxAbSvPSy/9tVNA0oHz3WZTb5lui6aLq26E0rtYufP62jbkwwhF5B9
Irx4j8gOh2P1Xpk9jqWQ5wm8YkblQhY+DPTPHoRuwOy6dqKMW4Ok6fHF8G9S
tR3lhvKxS95H/XPS+/FzUqmNvrkd4KguopnjbHrdYysfk5kXJzS929kPT6+d
BR7UOBHM6A9wKvsOyBR3lBSU4Bwhk8r1u70pDV5sNH4wjv4IPQRNstSRadUb
qgM3uNwkiMN1/gDwf2HvkmkTkNV7Jgi8hsDcjzxcXUWCULFkb1nzLKGw3y0c
cpxrwmoBxq9dZ6QXq/qmwNovvExfoUpcljFiNqim0QiwwyaKN3trDdORCNG+
tDeEjdU1D3/0z3UOVNX2vZeEomJqLs0aut0PRm6s9WNPD6rZ860SQbUyUl+j
bH9myG1gbN/QaK/5vTA/H5zREDFFdXtq5Hqo3uDGx32TzNxVUrteXW1W6+FY
7/a/bxuy39aY7Cv11j9fLg+LDpUOh6tBT3LgdGPHZgu6jPrGmfvDHPaLpkE+
eYsZLRGpIOLANfetBUCecf3flq9/Ve/VkekVHy76iUs1vvBAlQMD476K5hcb
LytIVHb76G3tnO+H5Sjq5jDqbdgJviUfYb2X9B2uvR3q4P6XrcY52y063M0y
02OWKOEdNQn06IN8XRrY5vDwsNfSau8OQvNXF9ZXJzZnkKquOXQlBYrco4/H
4HxTkkfWPtKH5h+2TJQZkQrDfzth+H14wwYmmLSgDSdU3YS6stI76TqtbQwO
P05zz3USeyuMytXE0P18jE5Ms0NUYsiQTI2I5ZjUciPbUOxa4OINW8BsXtt6
BfT2+xD3MH9mZkcUagqdW0Jq7+PSQkgx5H9uHaTOpc9VXvm1vX4PE16X0q9o
yOwTJMmCEUZ9hJuYOYhbpgQhAoqk23HGIV9V3LQymGjmU4NWIx39Pbyoc/GK
VXDh894PXD/2OH/5omRqcCFYhMpxFGq61aekpfTFo4+8r6DyCSYkTaXMdgvL
64YJcquY1GWKqu5aL7B+3ISjptvp7gW2kfbkZ9J7w+ySXSytv0I689RC4S4N
xghd8ydzXuFADNvZ43pFKrChvwM4EUjjS4MRg12xkA6ipL4IQLQiHEFQyFkh
UqE125KocOANAVWbbQGWYKRDmU1/zIZ7eiPBMPbDj6SN4650YHEjqh7zT31c
tSufbORTPf3t5zwAtN2f7syYV1DGhkmp21DwG9LWh0lWEreSfpK5mhOzVDDW
9dZp4bXPKvRKjBCREOj/wzwPNsiKjEQyNCT74uMqM/MbPKXxS6660atvfulM
KZtZbJN9lk4Ao/fyABmFT/HjVFGKICi3of89HtU0HxEbrjJp6YLUpDwW16eL
hI84pm4OqLiToNjfWBo2pRHSe5UrouK7g5F+QZdeUzOyh6aFENRuBHuxmFlE
QrSdkRs7d9E3ENCfLnL3kEclK9o3o4TnqPVmUDkbnwgkDpc5GvK1/5zkf01D
YXwCDiM/5VFaBfo26n1aJCFwTtTEbDi5M3165VlzU4S2o0UX84PbiN0egPyO
/1vJl+dzbQmg6p+VZC2KwdUHOfLzWZYJCHzkAw3i6T0SXfogNdaUp3t8G8gl
/HV/hOG90ShNZH5CrnvLBPwASwUfooGUOi+aAkStKwuUiOZRE36wl5mGwyng
2xxTwVubzPQ7jM2Z4o4QvREWljehHuB/XsFLUQ/JWyepZKXF/E+Wb9/PiW9K
XZ36o7bPPOx9N4GzSqN7gJ+D0w+vnSXMAPTN4m9S2MXpDjq+pJLA/DK72yvU
mwWoS7tM93UiiBZSSotH3tMBkwTqSASgAZYWEVU/rY1c50NHs7QUBOA2Pzb/
qKhQ+W8UdNifh2+zXGoBJ8AWUxB19TpzUWItul4pjpan+5gpYYEdTf1CZAKe
upumNPM/o4VdCnlfL5qwD3GbH743A31RUK0pq+rOjqwmEmYCEITkmjW+est1
bM+Ve21JmwyA6P6TJ06TCoDxo9Xbh1aYjPcSq9LXlJHG6wwG+3mJoZqcvIz+
j6qdtsbPOK+3dh2453ksqFdTPQwF+gRLRl1vT40JTBO7s0MpBnpRvIWMGpzZ
SmraMSEBRlsMQA9DjjkTDfVph06D5/6X0FYAnssYKM12j4dYqXT5/9wY576U
OF+paSpWvMicYhnVBDlh1zlwFXqX00/mCpQHeG6iQ8tjFTWcoX64gO0gJ1a8
3xev+gVujOL4DR6ibacQAzzdocPOxpNG1ClMQ2ttK1oTjLUsY7J+hYZntmqU
BwNqLT3NieO8N3EXa71oka3y/w7vtoMVMZSZl3etQdZN9Y5AcrwTqGTKWwsD
ZND9ZcdWcTTXWvnZvuK3YjvC6JafICgiMDO0YQ4W6KR8jxLI/TW7wNyVccEl
lR706aHBznnVJgAvp4ilX1H5xfZ/bqBgKzm1pUjw/3h786sI8Fh37ohepJZt
n6ozSDuGaBgHnDhyuM+2nMXjt75r/A6jWNTo3OV78Lf352Jk7NlKgI3MhAF+
y2JxlNFiCR87KnfPwYH1W0WTAXhu32sE89COsVQ1POMrlju70n1qaRoP+fgJ
ppvJShqHrba14lzFjBgiQ9mAjQi165rjxn5pL0IBniG4DNJhbdM5mhYBCq9b
CBVWURpKXrYrYdkuMmHYjehia5nguw98vsiSZ3M0Aga58yxFHoqYRJvmLAoN
WvzUxIZ+bjh+oao9GNBJjHbfFShQO4t3hICM4zE5dzLKEhlEc6N0dGBQpgxv
naSzsrGeTNKJyzidHmvvBJBLCpI/1LWG101MAwvkDrxfImacc6r6T4pDMPU5
+jvSQjtpby8qQmRSNenmXbtdkLePDiK2Ue1B/ZOf1olTYauG4oWsx33GnJTy
1VeJDWJJg0PVT0JpZFLrHHqTH/U+byREVNB1sAw4By4qqc17rntZWCX2570V
z0E+AtMG3DfWn+xcHleGFh7u+Y/PcKbN5rzztyxNnWGasgI888D7MHUcEweQ
Wn28wNH1r8ISmNxfgwFOrNP+tLw8CsMZ0kjl9Dj15i4fQi0gUWRdgM5c0Zmk
qIAoBgGIZ/CUcSqEbCmC6+rPevRDbkvFhjda6uolLna4b0Iwqrvx5Dz3GN6W
m05GTBuEnnaD56wBwkf93Fr2iiIHn28VJV8qbkIEHIwqlnwn8o+n4qMhB3sx
X/gsnZgkfrzLSiuEjQdPQjhA/38bq3KLONTK47ni3U+Yd3Um/ZjytIsQ7YET
xpH7j3PI7xXPKlN5nMpdWMWSXLZC114uU8T5uCbze2vhKvIxXmrsm8WdeHCB
aY4gnCU5RC4tff1Pp/C2VmMSboV7pNauMJRBV7XzjzuBsd3NNCNG1IhKf2hU
TJYhxGvRmCEn3xYJqZ/jRz0ueiAuqXtwsAl57aIxgiOz7Nos7XEKHN0kove7
xbg9o8eNghDIY6iHEiSKpE+ALEP2zpik30ul/sAHu78EofUPRQUPX9wP6UAH
dazXj+6rQG6RFpr55VLP1SqCui9e2ugutypHtNaUX33mVgJOD9CLxKGHKBTg
H2WU3JKD+t3L2rLz8hx8jSA3Lgm/K9QTctWWa9FMmTnb6sBPg9l/hbVVNZHg
pGsUj7dvxpICurWqK8+Xyntd9SQf8RmXyrw0t5u6oWZ059fRmO2veZ8Z7y50
veTUs1YpgDG+ljuYLfPIxOHP9+nVEHAa3xSBQzfP6vhopGSnDsjyVsJhFEwC
ny6QGAobUH/KVDqCE5rX/hJ8FNN+u+R9lj7P1MHNSMbTol49IKKtvzmxaO6d
3n16CoiEwYTn2cWJGryIUrIlXjPVrV/KzLfzoYZCeJO2fi4nFWGIS2xy6yu6
9McCwIS2p5jumUIofUW41Zm9gLdTnD56cEa65STALzfxmztLZ7s9IxZi9vSX
gtADHf7f5IHqPRM4U0/+Aam+4Kt9xMgNV2em+n2icwyiSPZLqbYAztgfbaHn
J9nOu6eYbdgimoBQ/BBqHW2IAVhGNyVMYSqBbZDsnFLIsokiW4OsowH+FBg7
Ou1GmVbka0buWdL2nomYzZmec5nHKu59JnuquM3OfknNB/zj6wdI/EuY3nL7
CI6ViNdejpS2BG6YxOcNyAWPAj6ovubbTOYxLancuckEcH4pDIlMhr0MzHWC
LuqSK1CJspifuEct0xyx7eA4KAwCKBfYsuGERaWeQEYgJqpd6rRyKmh8Pc7I
hUrVAWiJKu1TjLnQ6jHeDUrrc6O/cRcTYZnDIsafVWhR1XFOBtWbv89rJga/
haxISC7iRCLiq5g+F4tFDaGEGVkrKm74iRrjapSHIk/3VjsrBraTrKi2tuAz
xpo/7mrJFq5pv8fNZPXWHFkF6w2KWg5XSXu7f2iscicD2Tl7PkdFCAEKmX/1
nBOrrGWl957EZnKLTOKBg1S1/JLjD5x+AOAqGFckHDHrv9nrbmjoX8z6OpqT
irFc2yL3EuNVkC0/vi9uIhppOF9pGSM6stiiKk75BGYpbYcjHUuUxcQ3k+y2
4o6gGgqtHHIFtVKziXI031pzyWZdoe1oEV+BPQ1aBrtfrKEQUUvE6p9HLVxF
bfh8miPDNRQlJFhNrmsQ7yOhekdmtHWxi9dFm4VJExtoHjJ3VxPQK1nKG/Fb
rjhJfdN0WzeYKeJVd92QEYg1tuQPchoyksNjYRxedoHM/O9rWvyXgxgRHbne
ud58/bbStxIA0YA8o45F3/vrwEC4UywnZ+8xQrNFvTPrS9UUNqzEndWh+OaI
YCaKWHhRoiHGSHV3EQAwLkJmMZ/bR5fgUiWq2izpup/3P5ERBi4gpEmKdfS5
0439cXi6izDybf7kNQcZd8tNULr5/1DtVybgj8msn/YQu+721+K2MtUe0R6+
NYA2RwGacDGBY+pH4m43mtebQ1wWKvGm5DHczB02gTDSrluLrQ3DerZJ9oUT
3oa20M0TUlr++iqYc/vlU8w5MW9xArntikCD3fOLTcdD1ukWcOCEZdP2cI1K
KH+Nw6Yfm1H3H479OsTZj/YG+3J/+UVhpX3xdSPX2yiyCu6/ISCMEjd9gonZ
4hQrSlGDZL8lIRQdOP+PUwTq2E1iS2l5sEGj8aNmshGd5ONk6PqcdyB/RjrT
c28Tfk2K20DnPhIYtmAwuws7XuFBZsa7760mPCRqmmLTFkeBDTcvL4AOAGCW
DcWIt0zeK+U0AIBE56ER/wQS4OcfgeA2z1uxxlnVqOthyxZur39brLvT6RyP
PkiCrzpOlv2RQYP4QoUpEO1ToUdmdjZUb1X/stYJcuJrnqQTVy/3z7Y5Y4Ws
5frPtLajB9BwDTw0AivUiAFEr7uWVXVSCJA6w46aUoUn1DaVzHjdTIbzrHL8
D0iQRYIFVLX29GWc5nffzHFjGPRRgBU60y7q8uhuKZIUdbPuO1htXe2ohQcZ
ODSMCBS98HALgaURcBpjSyxdpFKBUMeoM0Em/4pjiaezpbS2ate3bukSdm3J
DfBZU9vkuNWz37I0tXU/kXbHAiuqdI2sjogsc3jyFlJ3Nn+BqVRiWjNzYU1V
C0PXXvHIQjyUwkWAbVpfuebZ0urc8/Izh5ZGwa3rrp73IJE1HrfC9BE68e+n
HAyraSUk9j155nixM1NjfaoWq5cr5bUiZ7kH/GvbLPAaEkHpYOV+G6uUsviF
ewMiyoj9TTpDc3wigh0Cqem9U5a8iQuWXZTrJ0rW6F64q24QYCPZasw3aqfl
tTW7ss4XtCOMjfVQ3XVR+5qIMZnvN1ILUYLx4jRZ/ygGM4u3JuMXfw5XYCYx
lZKHTbL+KXpZUhCWqbej8O2w9ESpcfCppBKZO28UYwZSwXKA01zn7LNdBQGH
055ouDTZ4aGcRP2vlA01rkk8bPniXAI3/T4nGhrbBDDCDLL2NexCXLLV95oU
tH+FEV/9sx+LADiLFVSl31OvcNifCTxb7Yc6RIn8GtHgo2DP056wmb/Mg8IO
Tt4ZhUu+1XIUXYWzZJMd3nnpHmFFn8k4gUW4TdnHzj3av+0WilqeTC8BlvdA
yuXPzeO/PoMUSj3y4VbujO2XER/I3jmj0pPwgW3ls+ba0sOYueCAWoz0qoif
S9FiEjqAofFWSLu4X1X744yEE+fTPs509t2Dcq2pCm6afulnjWBUJyitOBot
KdsiaaABGsahKU4744lIhopK4dCKGKUy7BG9VuND+Ge2qst4JjXWIlb7qY29
Wc9Kg4LEzBXZ+9pOgYWvYkbFDKvgukIXtpcr+pGgjvcxrqVQMwG9qLlCDQk8
uKpfiwor802u7ahQoc03SAc409E2jCUvozKarLTyuJbCILy7olPgeGenQ2px
0/tMjeXrTmWmQl8KyxN24ABcpNX7cUkY+6gK3+MGuM4p7XyPDFWe+DE6YUB7
SAqeI2c2v6oqam61zgwhdULiG74ePNy06HH1XTi/y2lwtZf/pdNiivc6t+N+
eLSuijuT1j565KKyfKaL6VDC2/fR18M2w9DiOLGQiR2F8OUjd/Y7H/iaF33X
HSwH15Vf/D3veFVjO1aO2WoaibNtMNwE4D8fSySPNixlv5uiA9AW6jKe/+XT
SZkpnRRvtAyiwzPjVMHJkPeePeYl/MOrqIWkJ58dwbB8sLVXU/05CcOBg5CX
+UuTm3J869G2O6RsTSzMlLVj0DP65NxVAqvK2PdMtgCU/+rFJttYtAh2HYZr
aA5ZV+ohDkVVQp+8X0gHo+DJ/M8SemNdsQ71wqJWIrzo76GwuxeDBZeqRjHt
DEtKTQy5hEOu+1EZXJqZMV4vc9D1MFii5PWiLz84L6vZOGWPrKRutiKZg/KD
bGNQFG6FylK9SSKHvSpDQfLVZNIUwWb7RnKzb/w5ytYzQOWc8qevnkXhyj4y
NPnkdQ1J38cQkuSagOfVccmj3/sbvf2XEaGk62zEhUxsE8Ly7zLBh4ZX33zK
G9i15bDGopWja8TJs7KeQXKkMpa+KBD30DuerlzGcAmvWeRQJFEb7w9WdZzX
8v7Fkir2lPjInjMVzjsSFtYrE2IQsLoEK1xiQlta1DJTZu2pmBT+1FYmpnVL
YssiIBeSttPQ4lhg/ikJKI6je9D+cTgXB+yeC2kWx3rQ0GR1C7INMbPbMY+J
yoRo5e383w1Cx9UJiiB3w/1tzhH4cPpQiTOMjUkmhIyfeDssKpscXa3cq9J9
LcIBIqASKVcyWJQc1pvYZAV/hTe4YBlo82ZuFReKmdhcr7JlWjHYOIi3p6tD
pv94bN3uvUZFosX1MpC8ZdyoaFU8aTehIS0CXgZkMlBPBr5tsMiKHlUXzTL0
E3Rc3cdunCaeE3lqfXHhFtFGSyCN95xQHbTjWePjzkBExh0WnvPXxRvYR6CC
SpaOMfD/2YEUrjC6fr8xNO29xKZLabu+08ZC3NflIxIZ0c9GE5xElPRM2T3A
QSTbxHbnctsjK13JSMCl5u8b9U9vScCmM3wpTMeLH9O7YnZIvNHqgFS1hAAo
4RG8xfPu2khspF2peet65raoBGb1a6xmVLoAG4d/ULWRvOLivay329XYAMk3
rHb0cenf7Of1lUxx+zAHPwFz9c9TwbK8kgLCzWxgdpcmt3Rk6yXj9OH3W+1r
ZkwpGStJfBvaV8BcZahFKIuvYbzzMFf+rblm0RI0WOiqkV1RU28lBMGiw1PI
ombq+6neyeqEmw6rkc7ogW7bweQ7onzMUFXslGZgL1sIHbbb3c47qeRvtfs+
TVgw9Wfs7d6ASpCnNa0UVMDV9fRIg5y/2CXfg1FHy5TwieNIIFix7V+OdjHh
HkkXmUJVc8LQy79cc0ce/UFWUVl5PAok+K2NCpApbLUUQrDJq4y0drcUNsaO
o0WmaKv1RfIFDkB7yLSN16W1tmD9fjXxE0dApDgnKkvXWbf3gTG0JTvamE2B
UyUxxyKp6Es3O6hJEMJEa1htNKAZw/1Is1p71itoWsdQRFv74Mr0/cNjMmo7
1yR4Rwz+AgjXIMwFKtRCEwu52sRmE5N4+q7g9iiosaaw5hqscodxXwRzn0+o
4OLhSWA0+BjlCIIV4w0PN0v2KxilMRtEDBRlCxrz+Aq1ZhZKXCWyNTY41ld6
UOuuHQs4zp1TGP4mIsLyGWcGtDd1U486vRgVe9ec6Hk8quqG0qV4djDwFVoE
BIRAVHIP0Mm34quV35dPWa+3p+W/cZ4ESuE35lgBY3nX6O2xqfbTQASNZVBN
taYdio4qJB8D1axrZG+mv2CoeEw/zPQ5IYcgKNa9vV8Wm+dtXdSZsysT+yfI
IAUOZAkkVrU3evPmYk5Ij9lZtQK38dIvmemuwbKUcuSucHsXsOSLYaXhsLWS
f16Ww84jMA1R/FEO8f+byiWhtdiM1ri+GF7rsQFy14/oi/uaATwG/Or3RE3V
fvqnQNqg5id29AikfXVRjnkXpcuCvMC8tO1+F8v1q50YHgl9WmSZcdz6UVaU
MXcHz2vqDMmSFEwWRYMqoaxThvHxgPklhypzuQ+UBF1+5JVxEtghrW6GDGV7
tf13seRqVEOaQVEZoaNyZihX/a5WM9U/XqeCq3u+ensIeOp9D7dKG9tR7ekE
4+r08GgTg+lpauKo6BxRaWxc8OM7ZOFxsW1SNEB2jcHgYP2/RYGHFHjLFIYZ
vIuBnf4mPN0SjzlmdtLCM4xrvSetY+Q1x1r3ZkS70MbQN1uGKfSV89p+hOGD
cw52SLf3Xyc5zSlvGefw8K+pKBKf6HY3G2HiqnhS3K4pNz59A4/y0ExpF1Z7
WswslyWuouH66wcrj3Bcc00t4Z3KanIRQu22rxDGT2j1dY2MTOnT7l8rfosZ
Wx3sQgGxzfDZUN48FJvMtQLD31uWhB0A68SKwV7pNfNGtr8inBcec+wNWg05
BjdXWEF41DuQ5ukNC847OR9hfYQwXLO0QtdW8766hpkbNkE2YdMKXC7llZWe
O2yakVMQHsC0CwMlD/kGLvN7pQbX3IlOMGbYOejyrFwvouaVpGMZK+lYcz9C
pidnDJLf6EntPL6lH/ZqAw1qSjM1eyi6Ndi9WrhUX+bodURPC5RL8IsOOslu
6mBM+HuE/M0jsQ+GcTkRoAOqxwDjybkxDGM8HF/ToSghnePl7mCejmK/HnWm
VVBh/172i24LreJ5OWmCab/0oU/vTN33c0qjU8uEaiXoYi9lpQrDpmx2jTsA
OPsFND++zXRiRJFJ6Nec/Dr4FPx7VySabyQz3m+e98Gf6/g/+BXIWKFCScXb
1L7t5tY3FmbE/7tFnSKd6IPTmsqahGOgWd+zPB5hklwtuNTzegJ3giGVEBZM
+XX835PWrSOklotk5/2ke7QGz366cenqBvp9sNsMokykxD5k/ZqxpbgZFAub
Knto/xZwmAdKhWiSh+pTWmuyo6te3obshokL8o+DwTL32uWsS4+AG2xsF1u1
isntw/yDrYclzv/m9rq/sBpKLZcOhsCBtbFKWWG5anqr+lpt9CPL8LC422cw
hWD/lHjt+yXr97hEF1iPPnXk/dxJqRMBEcUO7F/JH5g1RYqmrtEL9uYOx2OX
jKYu7RqHzwyalKx8ItFOk/jD9d+jdUhfM4z5ex3emviYtg8EEUtx3grH4vRX
wRYRwkKYu/z/rMGVAxQWUbFgAw10sgoIblnF6qqeFvFt+QWUqLDfqu5ZFmDr
fsRHyzmiWNGranbLGOSw6419ttBhDvHPJUJdeNA47K5krwKcNjrubMdN2H2u
6YDjYHNENE1x3SNXgC4tUR7e1q28cjz9pNyOLeenW7PKwUCwdji1a2CmrNC+
J4qtn6DMQiBBwCvk2gpMmNn09wfWl+YFbc2HCLkHNtNL8mmy7uhcKtJasrVW
PZhqIcWqJLQlZOADGTDiMwYLH6xkRILJ5Bv1dZA/VtX+pIre1P9Rvs1wHkXX
XU8Zbh+tUOMMPAVv2juQ8naULRBdjIH90pWE4r0bJ+33vsWsPQNgV0rsIeNQ
5DyreWpHsUJkboPQ7QZzE2dcEeUHwn+C9jVusAcW1Mxu/S6h1PeeBqO7ezZ4
ZE95KvwwF2HXua12BJr5+W/jIcr8AWi/zZw31B28VOKfO3gPzXhFUyUwhBOg
bYwexHhcGr2VokvwXVplSwuWZQJTb389MzKQiO/A/8/SwqyryE+iuwD2u4mY
inW9KFFLKMtcb4w5e2IUHh+VXbHW30tsXwacw5sCcX+2PDtoY4XmmmNp6pqi
Qorby9ItWd7sKsN14aMxDyRzeuLc8ql0F+NvecpS+z5Bzz2bjYwb1q01wm5I
GgI1rBhD7Q8u1UAuyPRVxequKHetPYmCqY/0R8BEYJ6sc+Ltdlbw2imtruJO
bk7J4B7W0tL1SiK7D4XuyHkKVUYkEx2MXk8gTUprObuFkl0ULV2TUcx8p9PR
mWliBkeYDBGmIuFVOdUsWGLUsROlj+ZmDa3u0HiShInt/Z3GONcAX4s8m/Mp
VB3+2uib9cMGSKX4Liw022/rNhhZs3Bf1Kwf6MeB0JlW1snTr1xu7GHcqILm
jsH2dZ7xlaT2p2yebNuvMV9BFioOJQWNNEyBJhrA2VIjYE61Ofg34CluYwLx
9r9uoWYKktJL6PYonvvhWhVZbi1JM9mmC9OBwWnsGUkb+2+E35KetPyv8b6h
TkxcXOurLL5nSzrisDd5ryGpLeO2eKzgYg2GTGpLCS9z4qhv2VnHsNB7LFFs
ObJfobda+0oayc8BGujh/Hr74pqz2D2u4VzDcDrMxmgLqAv4xFVRC3UhfXHo
0CuTfDjH1t49ibQeKD7ciETAzfx5ZuIacQCFBxPTlMjtqJFm0x9k2voCk4Hm
6KtG8B9Cu8MdIH1kUSyAdd7XeEkz3xn+KRqukVLexdcBUAAU5D5aGQKGIBM5
yuKc81UEUaEPJ5ocE7KxN5TvvsocAzQsC6Pr2hlHn/wadU4va9IRUIdPq8lB
ag10D0cLPUCypr18A8m3iYRzdxLyTyugHrDRKbNOGocJEE7kIw0Zx1RWqoYx
/iTbx2VQX01yfuztzDrUNUaB5y7tKm0+xpm/GUJXS/ebsA4/ChxKZPJU6YW8
MjeQlmH//WuIcGvZKAP8k0oMtEoOL2jZjV6hp4LnsC15Y+8o94BEHx+dR18m
2qmEJ9p3fpz51/NU852F8S7DFr0rQa6bw895BCH9Lb14f5L3AbEgu6JQKwFC
q6VVw5AV1mt9/2l0+Gn1MJsY3nkSxjx+W4yjSnj4C7D02LrMB/uK5Rvfeh5C
scqxOmIABcEDHkYPCjc/eRJxFWxeFznf8t9vDfu7EdswedT5c/917TojfWej
2yhT4hoCD8MFKMkXdKGTBlUgRoOAoSQFlcwMYgOr8vt1Fz0In9pyCwv4d8s3
/9SL6oTl6SMucY3y3OZ39e8OQY37viIi8SUYauo9cu2R6DYb1k4bIc/xKGYQ
3O7GlPXu8LzjjgLxKrSACnt3rq3e2Hopm0Ejcr0NKfQPL3zSB/M10LsHe549
zRRjtmCWktfFbggMpGFgaW7qDnFYc9B6NnxQ84E3pL2XrmtBS7nJwiNJCM/H
IcEi47eFttbKjq3pbKVchJqWHi9dAG6flNtk65if3mEEanRILS7riYOsnC0L
i6VCm552cL2WpohIPlmDsqpulg82seHNaLrWUxpPDWK21oNl/VockTSol9D5
biWY4EWc/m2S4ea9sFOlavh8A0S2jxOjQJK4nIBuU+WaSTfOaolsObP95ukl
dULcKMeMJOLg+5rUdVdhuKf8QPd7r+5qeEYVrSfv+G3jAng9eJ7J5Jnub2jW
gTg2U6/g+Y1HHVucEAZj6E5Ue9VFgoGBp7vKg+x99HEDdjbKw8Jku9md3gyZ
jOaGKD59L7RQulSztaHdSSnWpW1dECtl3/4GiPhRAy3kIdvrE3m6IxHWz15q
RJTXnqjq9aoArCe7Cf/5cGJzbVLA4hLaX8v+kZpeU1MIpq+/7e7pAVAqWNiu
9mUpBvO0NYywBqtCvqIQS3a8yVufN30Qs9EQSIcR9ucZ3VuU57borMJb8Ftx
F95zEBD14iWBjPhNH46MhHFEHdPg5iaB5QdTDUhMh7VowAywgI972zZ/idds
IabitETajCCYkQjgnDx8ztg0/g6jtzkNtFtWfj1rJOYwqjuTf+5sstTxrrqH
u59faLvMn/0phEyYUKxl6Mkdo6j0h1hHZbH03WhvSZwFw4EdtG5CByosNThV
ZB0aLi2xesrafhCBfTUKijEwLJF6D054+4UKizRBfB1rbddfsx3yw3sId8g/
fnGuOSd2ZX4aqO2MA48J7WMgnwUvtyJij28Fr61O4UO+PBGYCdmP6ebrfy8X
E+Po8IGER6UnMebX030+E6r1Zp7j+dq4StV7JV5g2rsrfS1b5gWPE5NlMXj3
MhsBCiJ+sPx6uzMmm29/mcduHwXUIrVH8lM5i0BYDvOpmbqF2/MD1LMtt26c
HQWaCDL4u75IiNr64XEU42PoprXQvPDTXaYO3Ki6R9iXUs9aHcucFGUq0UG5
mCbbjCbK0IhmZfmaEaEeeXqXKH/jhd7PG0fc8d1kPQ/+JP6qPuksbboNsIeq
Luo+YcSfZuqq0KsBc7mZ7o41cS4sg1IZL6u9yFG4rsWiSVnIvl3xpgIYgOES
dXro7VW71xH4GqAy73C/7Xgt7dw1TfORgpmPLuCaxXvis3j1t8MWfhxcQuYF
PwgZMkOM60WDLuH3ep3ubywMd8FgrWz+dFdd0ohcqS6YLFqRt55RYGTOc4oZ
/kVKsonpItMG+WGWmscv2s8+CgJgWFgm6NNCtdpeFLhnQW09W3dbPmvFY6LP
kdYg/I5JL+Wa39qpbTO8SHMauOF69Yce7swcRHm3QV1vUJbu1eg0C8yypctB
I/PGk7C8smfr8NWEfcVJ4kNEHnVal0dzXoq6c+kjhdExCkQAX4nvhZmu+B5S
D8tlpyoFHT58Voxlrc5RmqFtRHEJi912G7arQ+c169ArOC2BFC4M+h6PCQFB
jc/9qEEVFtAOiLd2WXwrBYwM7XB3e5us5XhuO3Kx+aWCppsrV6rvXDSbQJ40
Yuju+3Dz/yD2NGwpt8A3JeBvhyiocUIolkbYhpZ/g3r3Spj7ilXWmBDM1wUR
uGVEUZnvKVa6dd/NalZW7mJaGKBYf0UG5nWrsmdjRMoutC5pW/MkDXGE+VyG
yQDwRH5U4G/An7c/iDTWeu0i8j9br0vzY1FiDkFYTTJ6bKY2fV+/YCHFxA1S
I48KnatFsN9d+PSlBW+fNXdwQoVUKts+/+MHZULfWk+wEF2BSdOqtaLxXVRU
K6WxoBcNDqCYg8AOB6I7xIhYsK97a8ZqaIWTsx28B+p7hMe38ObmDPanjE2p
w9JGqlmzuEnYYopqEIUZaoX4D1VSgkcHyCsx4xCzuclzJlkd+oSBqSawys+q
xVsA7Al2E8+EHSCRLdHErFvEK7J3TBpyhWQobDPRWaU9kV1dlj1Bp5fGVngx
pP8tEg2Bxe9Akr1beGxtQr436xmWQPBGETk27jN3I9kYskpr68MDuItLDflf
TGjy6P5t8Ggsufa1JZ8bH4VJ1uNwFzFjLhj+H9PzoeyQtswlIfXim5Ijw7IN
ymgdF1b5yd7DG3nH1lSFUKdk/tWcLpXKTjLEPp7IxPtuXOiKCx0BP4t456k/
Eblxk8hPuqmefGdjoMhi4lT8BH/T+8tgI8RJlJRACzKWV5uyZo1DQSU42QbC
pzuRZk+4Cs+ahc3/NXcDrsIp+i/i3SX4UXhuHGU0TlfqK0ka9SyoInss/77H
SCM6K17N6lJqLAKmu8FgQft3oUpr2Uu7Pvfi/eMS0jaMYSSqT+cBz6RE7vu/
sU/tmiTnHWeg+iXdWwxno5GD1CeYcV95dFPJp45WF5c1gT05ECA85YR3+qKF
JdrTEzYLnZWG0ZlOzCRbOn72YqS08HCkT4AfhdaP3/usWcBXhiW+5Bvf7Kna
6aR9Dusf3Tzkgh/dEkuu2OKq9ZgLZEhixV5S7el/aQekqG1+52ZRJ7Kuq0B/
4JIKd+ftma8tzfWD2TemLlwkiWLMga/fh/ZgWLkR/KbOp765LCi9AjUJRqm1
whFIpivBd99XP61y+nxKvir/mJUDVcYAg2w3kY92JrjoxO+Bvmtf/5xd5m+S
Ow870FO6sMAsGOqWwNopQx3cnuCx7dPcEv/WwhjG1WNadIp54piKKGTJY7rK
Kys3Tf8ScQaZnPn/aVrJNTKQb/ryLoqUhf/DNPpQtJMk8PSvJwEqh7MXorne
G7I6DT5nlH5LunJPuISToVGsPO/AtoppTIUoH25Nf8vpElJWoGEZCZatN8Cd
mUdzNyl54DJFeA44gHb1lMC+eiNmFASLJUDdknC/L/9cPFRxeswRkrRo2Cug
oqa3Dphmu2GeLrlO421S4LSE9+4081eo6w8avBBiT9f1bZ5iRzU3uw9fBBSa
U4ueXx231EesFnXjY7X37RrabWK2/7WJiJuzbB3F+aElwVsdmc7ci3XfNviB
ymaFtOJFyvhvSeGs6kCnNn21aG7QykYZUFrBI+ta3tFd7a0r7lJapSo5oCTv
dgkg+0NciVAqTy3r65JEZDSZVYDqydqn3qFlUckMCTiPNv+2B5hpVmCjib3V
N4ep6AeoDornEd/ndYsF52ciGRTQTtQFdwvKgNwAsVJAMdfoecU3wdkcXmh+
vrmlp/3pjpL7uC4Mz5F4M3I3xGH6XRMVOuBJMKvhjHO3s++oTX9Qb7rDQesv
tdpdFEUt9RIHUTOsldRKtIEvaGaZhk9lR61/Q+fbYXR2scApq4MZDkUy7qUM
+kB6M0IOOEEqKmr+WcNF07bRTV4v6ioTbq4J9FhqrhvI75L6Z8sZLE6N/s7f
E2sLeLIA4gNzJuci0V2/+FE0J/+TftRqApsu6MElwWBNO9/HJS5R3qtcgV1T
9HB4UCg2+e3SodA/pSvN3gtFRj1e8Xq6TsskFc3H2W71jWlplLtWeyQMd48a
28fcjT/pdDYLfOai+NiratR/Nx6Z6VqO3Nye3khZT70h0m5QM46cHOcuQbv2
UOkUNAsl1+Ztklnv8fVB2ocgRA6yoSV4QGv6ybYyQs5ccb1nh9f+fpr121kf
lUaFJmRl4GNGtrFe6aNK/9kBwVxsCFNdhWZ7Sh10PNpbCKZpYbf7K/16gWvz
8cfrzo+aD4DdnYZtB3uktgpAHvf4uI2Tk1+mToDNwXNrUR0XqwWabgmKl0Oz
hJiindsAxE970VJZdN6HBnKZgylvqkQBI+d9cBggsBRf57s7OiaM1CCeAl1T
udUGW/SP6sXpamWu4UXTUvRHM6egljJtJoKZMML/s7C++eJpWeqcOAJVmYlG
XeTeOA9h/FPgjhUTMrcM+RWhFCBLmmjkhf4HZ8yu12lo1MHHJBjQIMztEaL8
FPFFMbrd58Lm86dGkeRCvkseUTrIQ8gGqjtHT3n7FQlm4uaReM9wgqbBFdWT
X+d4Aoe+6bkK1FNGP2x6j5RZd7uqT3L/CZ+icL2FSzAdS+r30dQ4/GgagjKD
RcB01nSveVfJHJc2ZpFQ0Rq535n4NKjdTwPzO6HTYAlFS+NHNiCbiTK5g+AQ
zbh6S5f26vN19AaOe+JKqmZKLDgXv3E4N1ywwl3OJqHg6rUx2Ssjz/5KqDbp
c4+PTHQgR0s0j5b8q+1weqTLBEfOQUCz8MOJx+hsEXkmQKp7SlWwX4Tkcuwo
9cJG3BV7x4Sodedxj3q9cOUl4AtTGQ6/mdywd0h8ua0meyJ5dc8jtIGSsTQt
6WsqJDnqPYowFAr89Jb6bxSawppUcW6L4VoBf0Mds1KRzUpv++DnYhN48bAD
ZC0RDpjIguUOYC5/hVI3bTh+O4kZ0cQuAXGkl1EVRGH45Dn+EA5Ga1bXvt6g
dhpx5+WJz9qVDGtbEDG8QUJLPvkytUex2nB14dDWEqbesva0JisXULxndADU
1d4HpfaT54AZdBIAsb1Ia/N5AihE/VE+4nrvOk/EmyZfkQcoPRqsPm66P2iT
L9hxCtfUIW/AiOkIrocxKpOB30GTzZbWr8k1/ygG2GzDDJKwQNLZN3gT/Jrm
dhhBePe+OCtO81b9A5fKgORBEea0MN5MeV6x7zjXLKEnFj4GJPClykQySwas
c0hSicpYOELsiKd6+tnd/XF83ykJgP2zYqU3/zmXVUpNTGJjwBEtvmo1bGv0
EUmY+GxMMPkheZW6smooyCd10gto9ZNKOz9ykn+XzLug/lC72eTDNZ+KBo5O
3aMpKMYWFtMRVB0RbVKIlE+8Vwadv1NT0pR/iq5KRmkrGwSqJdCjEesZDy3Q
pYqCMzsG0/3oFqN1AFibZVZc4WInd8iVhCFxNKV13SCyL2hVSXd9omgFLzI1
X3/HrxG19/NU3lLr4ByImPncDu3bWuIWkXlA4FPE5ik5DL38n/BTbXDd8iVb
JHsajM2AZlHVh+/K+sN0SrWGXWas0qNLpeed4oq4i00mDtqu/GqAkvKxhXKv
H+PynBXcgOAozH7IiLjSoIjj0VHsbkN3064Yi9Y/rEqk24b5SIZfhuLRHgTN
8ScIiRhVostGFspeAZwGStV4L+ur1v1LjgeOD4r/U5RVYgsqrAoKWGbjIc2M
6wHGUj8Xw6T3iaRp8kJjtNxbR5pNagQlZyFcx0+u/JQW2478uIG6KDYzPEYz
ooO12lr99YTGTQhLnPxko2DU2lY2mfXUHEKbpL1piovvZoV3AhcWNVw9b1KL
KxXe5HsE8gYTUZvsI1lUK2Apeug55+Xd5uZdlBNEgXSHDsXH0uILo8aEvoG1
tUmIfFE5AFg7m9mihS6RgDpLtQBl+BZabGTIT2kF80t8b15xxOJhNssFqkkg
v9Aak9ST5MOes1t+tWYa7aeqQAuy+O1VK5j7HBFSis5x5yrL5zVn84AIV8Zj
tK9qKc1A5laWA8ti03mDBIP6Bti046LYgL2NrT+fpHcNW8pwDLSsUMM1DOCX
wWqwife5eKn3UDQ5RIt1mQyw4WJhtp8LdPGrc58gRpjrd+Uz3IplWt1TCU1b
ojTTHVJebLTcG4wIAjlumb3MbtWP8WZQAi3VfchkkEu7q8L1zvW//FUavbHM
CBDHRUndjTXaEYTuZpitF7wG4k5m5nK+AQSDgjs6peXUVcgyV74Ti1RuZ+9g
21BJ0y6qP+m+gTO7z6sGDu/CXyutKZC6r9lGTzXNL6aIUce9jbNvAFBDha89
JeEq4YSBdH7Cp3Qhf0gyHaIufwu+Ez/8kupvM4C3/2ujf6w5AJVAAzYcFsOD
5BVJ1tnHIJ2AIwotMwOW5bDrF7Q9X2+LJCjIVR3zteKNa/DqMQstvevaIxsz
nYjHCHXgWdXVCPXwhOQYA9hRFsvI4nmdsPZ2+FzV9HzbKzjTYGN/6b+mocAL
AZcOS6J5i+D8/eQKM37sMdLdQ8yi7ecNUb3Tu19BvSNJehe1jeswe8ulhiqc
48FGQn6HX5VaQGjPruaDKb/VDRr2odaMw19fc8hfrGKdpcnigNilBjKKi0YS
G2qYf8el3+gl8mgMco112iOEYLBvamN4dEEBSozESa8DVnvXas0AbHGCJ4/0
ow0eeMEKjwkN8TPbP7UlerdhSU6MzQduTVHY+O+P1iEuf3lYLGdPO6DX5kzP
YUvDCwRujLjcs7WMcN0GuqTZbIte2huVYA5XhnwgvTpr6prahRZ4KBBQ0KAe
2ZsduufWAz9xWY+cPuDVfBn/AtRJ5+aDEfEZsyT25VjUC6zzrFRvOPjQmBSE
2Wun5vjN/l+TGl7wqVvzw4g9CX4BYWmtVf365cN7irVtIuL1hzSrvGSPcxFO
9SjHlPylUgYZcvzvO3ve8mO2pzr+Kq/E4BpAojTaOa4qSU+8ToCsfY8E+veM
l5MeO64l48CwC8QHWijol9zsOPNud9m0EPtZBu+EjmDv4b+Rru7PIkjTJDT2
kp5G/Tz3/zOjieiXo82J3NtZ14d+Z0nh6aCHtRR+amqe3ypH6oqLFYA/9MVs
BJtRk0nGf4G+rcx5FhbAVLYT4IonQ5UAfTdQyvz18vncZaVmagfdgZE9UYh5
RVLX0sc59+9z7hy4ASraHTOwzSD3ujP0znSGRNpB+MmR5sp0yTO1KmyeGI2A
tIpXuFLse6D8ZXnztru6/Td6AK/pHgKE6hUCPih1sGoaciP5sFBy00EGpfMZ
FnM0k+qhCDU0DIXY1+btjI3Lom8P3MZR96nUkJfM7HKwzHWdP3id2SMi3ZYe
SjLRItIWCiDgKy1vLcGej9vmkyQIxZms6HoYi3OuF9aK8Cfjd5W1S8/x4YkT
0KR24qxbU/HULlcnmaXsX+ntSGkPCoacBnwqcbZPiedU6vFDBOJWL0m3HUH3
ECV4pFev9tmGVW6DCmJSiO77wijIsSewLCt7KjEDeqh7LItc//USB2pqD0pm
tXemTdo9pCIygHPfea5AxguKrGQyv61OZMSOD03pln7nrwHhJEN0Q1pL3gS+
rvTQv/EuJxarJX3B8WwNXEG/ApF0yJm1Fei5Op6PIAiTuqK1wp2PJWHSfowQ
7neJRq1HAZuoMnKnAH7vynvdbkt16W/uw6lbbBJdb8ei+iqgbvV4+kPclbcY
svmi1dZ2zBIVe4bOJHEUlTn3beThauVsMdkCxc3UiWD6FV4Q98egPDutsJeE
IcCxkpb5l8PKEi9oc0IGqzvt4lu7ffedyLBsPbFLrgucDV4p4155vn9gUpDY
JusGvlihMSQT5jTZjNoIjmAiK2UZFqeKpvpv2mjSfvq/oUika2MMv799haPr
ZfwF9vxEwDHeeR28tFWH0GIt7jTBvmpzTtu9+wTXwKQVe346SIMb+iJUK1Pv
pamBu6LJJTzF5z7nR4XnzA4CwaDOp17BPOhblO5LoKqItliIefu3l3mK3akh
V8HwLE7dhV627sVH6dlqFTwN4BfOWigTM2mENAX1MEBEXdw4zic9x8ZHuQ+Y
xABMLB6QyK8CkgQmx4xVC9R4nscxB76NrC5XhPWQB6mJLA7n9k4nqUFYjR/+
23078cmHYvkiKbUmxSYEDL563ZUkIGJqdJ2KU3bqLO5CgAoAQrUxnCAOq2Xf
lyMdekU3UxPkcgojZirDFC3jAKv6MfIaLf/K0mALNGpsKlrfb7c/1AiXJNZI
H/0KPZMKSjNdX3g2NND8gDGQ7IrshNy9QUSdJhgDuv8YkfpoqADCuGMo+TGb
kTde+5jVnUOGrbfF0Yv2rl/yvPTRBfkmPxGeJa+eTfOhvIfbpt0u1Chb2JSr
IC9uGTimSGAveEqpdbkl/NZpcuD0QPdfY5OBGhmo7QRpshZoFtjwXzG6M8p6
b/dcXdXZMpIcmb7MdGuznhZJ/WttCnYcw88LeKFjPGCo5V4xmPeZzuamBKwz
DrB1NpFxay46w10+5glhwAnOGp6MlmINK3SwS3UuWbfP1Cou8HflfoUcceCz
GtiIDecS99kiLHnb7y+4QP5K8TN5AsNPDdut6leaOIRwSLD2XAW+Vj76tEUd
6H6NkH3oOMgFm4iUnUgN8OvBl3l/pj5XpiCJ2TrhvwzslzX298LcsHMTK9jK
KUBZdV4LCbMv+1p0QLidM7w+Tj9fgkjsF/Eznbr0GPwEdd0X20oq+o406FAU
Kv2Ov6kwFBc8OOMlvp4G2mvzCCzdyFlGX0oTz6lyl5CwWTnz/9tbRmr5q8vT
TOQ80zrK2FjDxj+i5yjyzLCZ+ZyDVqbDIFke7EmcKdFykNP6MXVBBG3cY+GQ
OXSXA1jZYnY7QSJ4SZYLy8csxiSxUL/3m/cT4YWSnBbcUxeuDz8W/jlWHmdP
Guom0GCpT22ksNLGmqvqji+QWm17rgeSTd7fiuXs4Pl3kK1IsRPQEZR8brHe
/nYSCPWC/9sAvSoEHgMutt6Em1n70gJnEqYV0olG6jabSTtZkFuTlmAPsJDE
weQcBhqeIW/pZ692wCGR5AqZcT/ENuO8dbFRioYJcP/ckd935OnCiBnQE3ZN
l+OIjYSsXB11qQuk6WAUq2ppS/S/lKXyJc2i/x7Ofd0VpfXbG+rfNUkKq8wZ
jODDNOT3tbdbx9VXjPyzdlseQYZenq6FHt2vAxIXsU6u4stugJz7mM98OWR2
QoklCvvWnhyhHTHB+c5dP39C6afl+WmPOGcyuifIDWB+Oe47/ZHWQP6WBkUj
gxpyh51wzXwIJCm4/K83u0o7TQxxsoqsWiJcrRnlXLoIV2yYTISS95KUUgNc
GP41MNkpDlFHWTZVpv/WRpol9MZZXqSx6MBi4ZPvxpoPksPdnwxe12ZdKPvl
bHon1LD6HwB4PP1Mes/QaugXL7TgeS3MznNkL4H4tkfbbH7Ws/eGflq8pI9L
I+PcnJsd3v/iW9/kTQddxOz1aLLxV/ybsM7s7nKorzYbx5iDDY078OgGa8C8
5ZxJPxOE+Wq2vc3TSVzqnKCvqhkjtvkMP4c2Dp+ScYreXOsxCKhWuN7XxTvz
oR3GYHBNvq07FreAr1Li+Gv8nLdjoHC3qrKrK16YF9FKyBdbJOuUw+p1G917
Qi33yPrnrVc/Yablgh1u4d1US3xBkga6gi3gBgQ2TEobvolpKMq6eMseyhUj
NwR7QKdTyF8onXv4A39zY789AIGfvGpbY2H8VuYSaEhzovadexh/Q21N/GJ/
gVat7ADi6MRc6urP+vHFmeVDNC2mV9AVPHRIunpxhFhZYfJVL0iRmeRZzQ8E
2Iz7rtgxv5e31ol5h5vS2Dxpqc+FDd+ZdsIkoQ1k9K8eDRqaPYa/De7ZhNW8
aUkFG/dXFkAYitEhaOeOWjpL4qCQGczEV7nOcDVEWPPyYs3zpqN2AUfyF/VN
kvxAqAKUkGqmPJnHY7uWZ/nKTMIDv1WVudQwIimaor9oP81YYvaXMMpiZ8nt
35unH7LR/ZKUlp4XQrdha8MZxR2wRoCrmmlQeIXEdHCMOwvZba8DRn1Ir60x
iX0UFrv/aZWmNC0kQOB1z2xhZHPA1Uab/3nLz3Oj9y9+0BDaTd27ozgFCpvq
Z6D9bjY5VeVfVHkLT0wwepbZ9n3Onm2xCIBBM/8MgEDg2MD0yuZ+alvnVHD5
7jX2hE7ZaI3UjUNU0mMPSz6nVbWnRPMHu7hXUUJgAAG1YxFgiMeu80NKMuRo
l5JyB7txDILLWiUrrFKuNE4IxlBlpdW81AhgGUauMUB2CVQtw8PDXKgG71ls
EYwklL0I0A/ABbQAfdnGbgBbfyb75RhDYu29pEJrMXhjT/v6WJfujELl8nS4
Ykc+/FAzCf2mkJ98C2fZwWJLjmJ+9j24o95JqdGpGR0HWRFoMxrYfjc0Q7qs
//Q0xOuUwMKm7h2iFhNzYZm8apEEe/5ZVKvbc9Qm2qTvQDdyT0J0Oc4UCWqm
kfViNTR6cRXhBcy0U0KU0UGlaEFlHd6jttXuKpqQhW+lf/LHVGgg9ItB+ROP
NTxfGKcQaN+XAIdQpQDTMq7JI3bWE2fxbS9v84kUXF8ccboznL/Ab+FitbuD
v8ahQrQWfFtL5JazzdO0wPFVqCMeoKXoM3jUDJwaAJKddwQNodyoNIGzWrC/
pIy1k9nK2x8L7plWRVnS6/Dj+zg0TNmRNbwwP4co3NtMB4h+j8LHBjpviao0
d/G+XI2XDDeoG5tUAsbVo/2VobDfwgFFa9fgvNd01Sy3qSeIWrj82tnqNgHv
j5dDr9kCTuFHWbLPcVvkB6EV8HkHDy69PQpLZ1iEfP6334YV6fo6gU0UGlaA
DG7rswivI3LWFxrCVDStJlAGnlBWCx+7oY6xiy18rkT7/f2ewSBrHB1NFCuO
1/SqGdQKGti81G64hemenBCZVlWE8C9SQooDwVNR0vDnlEdH5xFDFti2L3/J
Yt/jil0Z0/KIt7CTi2v2NUsn5eCcZmVN/0YDz9Ce+Em4bXGu7/QtZKGU2YHz
KoJrAclcs45jP52+G5qJ2+h6+FV1+1RL9AZaHVNQWHOU8OsTf3yVRi2pibUX
MjolhCUgZropPOUjmdDdPeiu6JWowZpPsFb28sb38dQDGCKFRXTx/bscRFeM
FrlGJD6HIEmRkN6tjODjiXh3p4uS8jvnkUJ/bmts83zo3NqN92IB7cWK/8u/
rETRZ5+ZqikoVwip45/W5z7Q3mwv02cpcyIJ/pqxebTZENXy6XDH9Cq/Zaxj
fR2np8cj20E2NpmQNG7vxuv3QtOoIpbnwvmDGxFAPEPtfvjGhnSeJORWOEPu
KPAaa7PUnvLGJZP887RedcX39ZkPyRLNpYpaAY5KaLUiuhkS5wBE5Geo2e5Y
1t/zDbAhVPANv0tXkMHQFyCfOTgz1ocZ+DD0aUiVxIJCnCJ4K8jrN1UTJ3ge
3f2l6woZDO3aF7XoHsVMMTd3xpGariuX4pq+H1xK1tObscNKj2CAXtesWPkn
AUTO7bkOGcVTRDpM05m55bKolDDcSqx3jLYlERRdNrzMXWb6Da8BrcKFE1z3
D56UTCFFak33vdusDHZKXOILZcTolpQuNspBJC62HojEEjVA8BD0ISOtMV51
187K/dL/bkaix/qagenqqMSBTfAciXir5bEfAt8CVcwSIfV1d99Dvj8So75A
ZSuBrekV4BSg2IgOSVcInDDA3zATiDZfWzfw6xWldnPs0icniPMSenTpcMDX
br7Sky/gEnCo6OquaGUPRnmd/6/TG4IL1uM7+bjHCw7ZRnM4KKxunBdGnqGi
hYSSijCCliCieSbSmb/WvUIHX8YJfAq3/G3YcNfcRTa5W+7A4fBIDWiIoVDq
NpSen1uB56b5hVu8bTWLF7cQJmxzcrV3iuyG6bH39lCiGaCiJzmLlk9y6sl2
0i56kOJM6CR+rhyl8EtQIxnwE6G4O3J64ZxZW3oT5jjwAXHeanc2KI2zahgl
MEj6BxTK/rZ1urKeiZqKJ2jFJqW+p6hS734eByWijACK8foGTMG5AWURl/Vv
jiu58fs7sDOrtL7ejFDYtYoL2B5fViEcx1heDHeFqFYgeq4SFwxigbyQPUhf
ikHj9GqIWoUxQR57Fk6/TRC/PxvvcMhOT9wYIktOKm9jhPzshuWRd4acIXRR
tcXSDEpCo+avidOxQ5/Vn+2JxS327EGIbz9Qtu+b+asZNw2gj6MnYlRdyD9+
ijCxSmoiYVDBqAU6KqLVNYeIGK+PUSIY6bRutz/RUV7QFqUmJvYlpNFHNEA3
ISa+uiUhonQAqp4vW0D01cxej2m6LRWpatqGUtsedSylFG2CjK3ikxMbXwiX
8atjizVQ5CwOBUTwlWsg9RoPS2yfHWLMeqLqpxfKWbQXV/UkDQnaAmi9E4yp
cNT8ZyBtCTqm7qVkDMFj2TVjLL7Q/oVQynZGdmEUl4+FJt9Bbzoc+hIf4uPM
3mD0EYEik3IEwemDqJgaTb0FJFWkajLk5uvd4a5LussH6z+6Of8DmZgJAhWt
JjVN8zHoCyfFhRFijgCSunG5J9zJTYiwWtvhJgwTiQ5VqN0VOp9B64ajih8b
5EMIcpwIlyIkdRBSSu+2L1gVC56edsS/id5Leg3Y6FMmyv5cdLpxvn547VTK
0/fzDrtfaXmZlby8M4gRMrBGJOQWYVQAuyRvWuR3s4OkDLENirJlfKkn8MDF
EjJP1QWrPpv+YDrVEtm98L3HW4YTPWFJxcPWCJjKCn8awEhUg0UNVNm99lYq
N+SeVAkiYrGt22p4jcKQv45zaA9dkAsL2YEmcIGQO1oMtlxg6JyCp3F6pa8B
WBXlKc3f4dQCSpZoLI726qv2hp8F4oiLpSdCdkt860SFCzWxAHP7vLr5nw8m
WTA6UrswMzQwfj1vv5cAXC8qN4HGS5yAC33K7HTS3IG5uWxKAGVKkQHUzGjw
jC8WdDBrsuBnr03WtP4ROnOSbNoA/GdhowkrL+1bl3TBSjZCWYvSmHVq3zKN
AZa7h+NWwo9pS5kjhIyItMfoDNLtJn/0zMxR8gds/bAe/VANtZSrWARIYzdu
fsOu9hzhctuGOizjloKG0tDgLWeI15dsVYkgxzUI4XO1i7Wrx5vt9AUyhy3r
qVtzD0iFGNW8OkbKGSvjai3kD8ciLowEVfef3gqsiMiC2Htz0w3LvoN1p4Bx
R7JNVwFgkWi8qAZMA8mZm4FtAZ9MEFLiko1BAgDr9OzpxdCBPcCDnS3yHfnQ
bYdCyYFi79Y5PX0aocVSWNLKyVZug4VmctuGmo8wX2IhGC/PMz2wRSzzgc0n
x3P/beJzZ1p+YSrTsytuKSbH9tLQxTyIC6CL0uCw0dJj0xpOlbIrlHnDju9s
A+Y4BHYZvu1fJOzP6bn0PVqXsgFGm8ZvL+WaiCxw7BrLS5WZwRwZ8vshDVeU
+y6d/Kyqwwyu4rsTxGq/ugNmKbUP/gyPY6IdLxTpbXh3kTuAMPRVwGYd+LND
Fa87Zf//WPKs6nIGC7XsgLek2HtIjGD6hbEw9DRrHQVYZTaD2Kba9ImpCJ7A
mwQZ3NiXh7pC8iIwscltx3BulxB7MgWyQwEMn1j8r/1VDQ2qHwR/mZ2rvyVj
ITBycMkZJRAVBbgn+SyRGrAhKbpzHI4tnLwYcL3GhkFe8QUg0O3oOxGxyVZh
GAjFnntJadRZ1My9l8rj3iDG8/gaTQkLiBnwrZre2KPr+3FaZSpBJxjTrgyB
rfOljYmJlBmzxzVFvpyIfjBYh8YSr8Pr+0fY5kdu4Ae7tasgWu3ckV+5kFOn
oc1QUD5H2nPXyD+i+1ZJ/EjA+MDFw63k0BR8tAMtZ5nr1tFB5PlYOYMehZjh
YSd+Ic0BuqOb6N1ftpObqk1wPrD0U9Te21+D6ia4GnIaasMIp4iYjUYnK8ol
sbJePvKUQ/6MqJUSTdK/U2UzizRE5QHctSLyXEw7FjcMUA+wbTHysucTKP2H
Rubd9fw2BmLLr52mBjRI4sP2ShTvRuRHQqqk9ols/ZFJoa/qz9rK0F5o4Alp
WeuhToysXiR3OzM3T9S4J/2LXbyOE92voUGKmePCI8Xx/g3k7DF2XLLVB8RL
NlI7qZe1hUlfuNAM0+JUUcdH/yo+rccXiFg0FDN0w4NxmXh1Ice/s5D0ahq9
1Ir1peQGJyiL6UmdFhcuKmKfDE7W8jRnnTssTnHqF5/UBrSxI14XA5yeL2sH
KQtQUr7BHcMAgZKTNdy1T5kdpIfI5baL98qy5V5Rw1k8xwOSDTWYTxWcwOgc
eDqk165ZyRn6mDDZAAhaKNpOZgZqQai4+oNhZw17wWRE9SEO8I88jviwJj5P
FrdC9GwsGuVxpwUMxjMIpCojLX+It2r1sfDlAVZ/zFeNza+Kn9LHSegoV9Ms
d31IW5+RZ44kXHmAF62PAS249F1v4DWm1daRg8Tq3XmvvtRWRpuAIHGyrDSg
/BWL0l3WP6ym1NrMF0LeBrFe4w25R/MHEMxlXHJrhUuMSwSzbrRAPXE+IXsz
H6EdieN91DHP9Bmay4p/32XrCW7tVoZMZ5PFhFhjYuRF1Bdu+rwu2db4D6BQ
wkyF9/zdm0jtKCIU+NIDjSnktj1B6MFh+X9doGrpi4hpJaHWH65RABZHcxah
PliFjgNbCsbfpKI4mlBZV5D1lJ8r3gZ6qXOI9deNRgOngLNEQQc1ZnZKkjer
kBLhPaU292xXFv++tUlhqxSmIBeffGf00+1pXgDrWHuyq68a1Z4VMTrRD9wo
NMeGroRGaHZNtT5OrW/CZab0SNeUs8qM6NkWqgQ3SWe1pyArpAN3IiVPkVZ6
sVjbAx4ZmRBHcLNerz8/wHCzgK1NP8zXtmXM5CAFbooEU9dlo8RELy9nXY4b
+eYhBf1iJAL8dcCaC+DXkxAJGSZHUvMlN1jMOZoTRINz2Terh/29YRN9u3eq
JdNRG7M4XEfLzr5j4hm9bryLvI3Dsyr5hcbGoViW0fL8uG7ncLoJ2pPzdB4T
ivUiSY9E91SoxOmV4VXx6RpQfOSG0QiqDzQpnsUS/KWBEUzW3CEmaET4uvOi
f6hgVeWrG86j5EUBNYIEnAm/DraCdg7B6IvWxgh9OrlrLe81VQhlrB94xMTH
J4uaJuilWo+Ba7PkjCA2SIO5BSijhFLCUpetEPobXyHkQWQmWjcjTJKblJIv
87WO9R2bzloPlen6+TuOxFWQmyjcrANlayyFTmxSpLV4JxdCAZEAVKOR1R5P
t32deOi1//E6XglaCiQQaLlFKeKUUkcvIpEKilbu2HA8gM1G89bMnGQDHcPj
cxbMS7PmgzWy4eh05VwLCm1EJjEyps4fD6M6JxpANx8ZzOkVLjl95F9b7Bzu
wnJ3wvN7CRXLw/vRqRcDqYNnZ6AXddJlHuxf9tuKeETqFK2bbriS/7rKm3Ld
POkhS1BCmgs4umW3woePSYxo622xQAV0OwRuXwNkTMozyu/yUvuiB0wTWky9
/7Qgh41kyCsnVrRRTvfxYqqLE3555a8PMCguhH4tU0HggkEiA63FnfCQqj3o
1TbBjUJVDFklvSgyP6ukdii42uYlu2akGsL7aIbtgH1rPzJBvjKl3BofSfeU
bCq03yY04JEBTiZfxz/wEuNDM/NnT7t+boSdKEJdTTUlmkINbNRNrJzzNZzZ
b3n4DCE7PDQ2tRc35+K4ulYPm4i7ySdM4AQsp3qhyv/H3m2P7M1pUgyhgE4L
dllXLMog13IDFOK3+VWYtvs5NFrENH8muE/y2hUHB9FMeI+Xekh5dymXILxh
UQgdP8+/q7q04xtUYRqnM04QjdXNuKoTkH9HKekRlCmFIcXTEGHJHyw8zlfn
lj493qLQLn71o7eH6ityYy/wfquyZBEpyyRixIo0kFJBPVzUL79bqpzFZrn3
Nvk6ZSP8yV/Nyp1e6XDta7qe9A1A9wynygVO0NbUbgTSfzN8E+lZ8BYtXg1Z
YgmDlmcYcRm8IjfLIl6JCpK7a2ZBrdppI69i4cTcCwOVgd0jf2Bqw2PZH7AV
zQ/gbPw32pO6YUX95OXs3QPrWCrUP8qoxCAK6px2KWRJV9BoRaZ9nK/Pp1o0
L35cRqcEZ0FIdObV20AEzBoPWTF+Ha/tTLyqg13GT3jbDh8qovvXsyaKnGvY
4+HRuBHWckZaKzAfbpMsZKuPpv7k1jrbXLuY95e7oGcuWmZX+vXa1+BoKUhs
7Xu0VqMSbyACL0syrSzLMjBUsH4oyHbdU7dnr1YcxzrYpGcO3WzNaOzU9KxR
bbkaHfGchfVg2ixty9RXPRUZ+Iu7UgVOXdGR8iMqtBslpFKuAYA46IrS49Mg
AqteqSU7Nh/RHcYDt1MIXYYQwBzam2ZSMLkOdmxtSySJ5VIaneFc+W4hIQr9
vu1YJYdq+43IYQ7cD3/ds0CtoYTnKgH4Im2JL+NYb6EfCuPjjaHSj1lQ4NQI
+Gy5tCP+83AZhPRt3J96xJAqnE5OSKuNPkZDwWrN9p+u9n7JiFefx7I3NqYX
HkEYWrNMpf0V1+6kabMp/RvD8Vc0aZwgnk/QWVjK0wAZhLxhDYTYZ45TuVXN
9GF5aGhODnZ4SEvzsPOOreyjdMWlMHCzDgdgfuZB0pBrR+11BHKq/Zpmz+J2
Sb2i0srjS46fKWO+H+Vt0Dwzp/8uDcFV/CNKVctS1wJSfI0tV8D/Sm+BfRI/
yhcKeqUdqYIWJl0heolUY52EeIvY9DYoLGuulw0qXjZkTwLN9ymM/qsZJ1vJ
I1QA0ea1iGEV8h0E2gyGzFnngNRV6nhfNrI1SrxIsDuz7iZ2IdoANssyIEUe
InYHrhL/acT4QBMhlsPiKorkhchM4EeHapFc3m7Qi2F7Dgn5Ck5VQXv+6TP7
gZxeSdJcC3xUn7gpxufAkCbCsXSgyblKhRzylxdAyp2Y8tMChhjlSCiKQsOd
pUF3mufoiQ1c5p9j8QIvhXm9tKnqQlZKdg/fpPSQ2kswQNMrUjhtGLXwvvKC
hCrz2zdd78ycUixaL45cCOjxQ8kGqbS5dwrJR6fGy9LGMRx5g2tBHxcQMJ+R
yGKVdvgGro52hntDiGztfsRugHROTO7yHG/jkRahxS6u2+ugskgftcZeWRA6
e3sldwTAq95AV4YsxhYPrahnXN2Jjaut7beNB4Rr3b+OQBfd18TVjaCGjXTZ
tKBYPiv4UsXDQnn/seF+rSUrCHA4B7K0UcKyI2hiWeUauiAinHZpMIEjEyc7
bUTYOkJQblGeKfVMBld3Oi9LrIEQMH8IOf3g9ZoqEVJGZuVFr1U+BK8GiIGK
Xg3Kiq9lp8dRAROeYN7DutvzpthQKFbC1He1g5hTbgtDgvm0GCAPrsmPgxog
RKnN5s26dYvFLNUPTSpvESVPT/uWOEbc0jIrI4Atkpw6DXBDQ9sFG0d5zq4r
JWG4su7sgEIYqBlDd0CId8cOGxijH9dGuqDHEeipNw/O2JeZQQHYjoBnDXaU
1IUT8Cj51Rwg1OffmN6zlqUYaTPMZjUKbpvJIXiM2xETqzvV7/mfEav2dtVa
ldD2EPokp3a+W6KbZrkH7kZBvM2QdYpmiFY88YFc7Zakb2Xj6oNBl1q79c0L
OIM24KfkvGi3RaUWEQg9kqSBDhFJQ7ZcqFpFNdffuxEmy0VGWI6vc5BEwAfH
tsXh9xjjmXnoQMxUDQndDUH/16H4hPvlkc6227/2K8Lnpw+7IphcxTaM5w+l
eoEhJOQclg5AHTIfz/7jF67oe9mp4xbNOqyKL4x4shyyvn5SJdjiKa4MCRFw
Yh/yOwzy1f4pjz195PEK93gZU1/lZa3duc33ge0uWwImx2O6SRiwvYpVbsjV
0BQ5+ZN3rz3L2Rg5az2QC4LQUBlp8t6kgVTm5IncjmoesZFFKeXTgf1nCZOX
iroZjESeEFE59YWwxcmzj30wREjYybp8nF06WKJVcsS0WNkhPAXe8gRdNgNl
IhbIm79hxqch92t0gtWWM0keshNn0lo244+fOrCA2DXvjXNp6i7Svkt5sfci
xy6nbNHZsAAK738cMme+geYGnESSgFfsjaki3eZ6An7Ti39v1Z6NHyjlfxRM
ijT5kn2zILha565sqGJgKKbu1gAHan4bXdYs64n9zxohxoIqfkqIChumYDA2
Djn12lkMBDftOWnByxiSkmxRRhnNN3jisME+xeJ4AtdGuRAM4svPN3GI09c9
/eWG9e30VNr6lzzQgZfSY4K3HEpX7IdfbSdBMIW7Dr7M5XVIhiRjOWtmtV6O
+kMJgWIHtAxTljhrq0ZkWOFWyJQunmpnVR49eUadLIHFPjbaPw7NGs4w181T
2gOoMS1upsCbmBJTAfJQUPpSA0xSdOyiwMFIViTipg+7bqo0YrdCy+Hz6fZP
+6TP2sVL5Rxr4jaixHYJKqHIA7Un1sWOju0rxp5TeAchUmnO8S8VSzFkkWKP
r4oFDUilIOq/opvP0hgasTXfj0rkbsJSzaPe7MuFgmmOSGpiwOwQNjk8UfRg
KPbo+NsjEOQJUX7ODQKuAefyBFpu2s+8Q56zcTnryUl1hibuwyyPCmTqzru/
vdp+lGXHCpN3cb+GnQLbRKfjMvnWPhoKZs19RWPAP1y9HNT0upM/J69MNKtK
fAcVLBxnVNt5WSns8lnuKNdbXJnlTdxKD57/tpfNgnE606ppIkohEUNaSiiC
wOHe7Jsvvjot7GS0fwsVxIMnmce6Eginef2sa9ZwAHmpyRvjD5KxY84NDgdE
kfX2rb7RPQNWyo+lFYTjy5jEL5WMRWyH6bdANKeLoWzo0xebfGY/q7KHtwRL
dpPzDISr3EETiwXqIqjp2VZdyjtOjcPiGaB2YUI/zNUjXGsCq8/ASCHnSyWO
Egf4SWnGpmBctvqdE+rJaQSYuc7Afn3UPr0EOhFn0MGTrjV38bxwJm7YvdmF
OQL+d2c9A9ciFnp1fROdxW6+gU0A/EZTs8A0WL58jIYRUn1GDi2S/ZHxz4MY
mHJf/qgLmYgFvjDlROL4uYO4o9mMqIciiM4baBr4+0mcxx56Q1cxSnwsjwVj
vcWPdnIj7v5evDHJU+a1ktK7vdym50cIOzaxW9dKwIOxZ470QiExoUfNRXDy
dJu0f7/u9Z9CjtfLol8MbQpRc3M9MFIkEggs0IeQB6XtA7tYqvWtkpjXE8jV
qTQJvh/vPMiNRw11s74mcC61RYj4fOHqEKkssQt1U319eFnslQ6yVBzSCcM5
lIjsae07P2acLN6AwDfTTg6LYnAWk+i/gF+qS/3D3N31Kw7ojtG0Q43Hln+y
fo0SLpvUnu3Asg9Z/kZDnaEsahJ+GI9eDpysH9xorG66oC72Rw3A8cjp9u1i
ierkhYiU8rB95L8vOTgttQJ+uehK8wHADb+cUk1U19cjSzRKlGEoXEQD3M85
4abSofb5stpLxCxdzf/Dtm//TwTHSVB40xoBdZsXEtP0L74jaNIWGwe1YYSA
Qf4OPosk7bKTM1tCoRRxVsG4f9nSlj2Sh+0H70P6zNDEYLKQ6hgA8zSXU0xy
GU8YmcBcrIka+v5n1BbS/KX5389G0UBlGkGx3DSyiqTUgveFQ4gNA8iUumzn
7Z0I6s0QO/yZK9jw+QK1MHpo/M3ms+veBVKli0R6O0Gm0XAu/txeBcMYLdJA
XEtFnFeV8+nY4U8cVMx/rL/DkXX9+YlvFBAwnmysBZGrMChPSNRfgEBeiqId
/ncI5zdvYn9BGkphHpiulFEtypg8jR9QG7IEpxFyeK3jDCKWeEOYheePwvrn
6YrKSueML0xXW4peYHjqxM4LTR5r2UOF08azzdUkIIDEcsa/gEizUjNY3gCG
vAayaH+aebXmKe+Pwyx5yvUxZP2Zp920JBnb+i91/iToWENA1G1dMIOcgEEk
4dMxyvwpZiOqIdB8l61/MKRSNgBHLNxNpsivSJAKBsuatjld+RQzvZt5nKWg
cx35nF2ldhOxmHEpKWfE7UwZtGAN0jySo5j6pMSwjgmpKJ3UDCZyJztuRttE
Ks94g9XjKoSlO1TqXO1yah9XcBIFUJNmd8p5w61k8ueBrtwybfToxZeUhy58
vjmaw3x3uxwGKDzW40H77e2IzmbKDCMWGZUlXkVo6utBNISSKZf3rpVjr9gs
W7AyO+L5u3gUIm8CbgA5fuhmlmnVbIVhLODU5voe1RfeHGLZDXuIyE0dO9Un
x/epIvedbynGSIFHuFzs+fniV2FEvAT4ZxY1hjsvJ1Uf1KhD7hS0AwGdKPVC
KqfR046puavVOH5yfGLfZy6V+NslcjxQDVBxBl4jVSIK7+0lOOo+NuHWTiNP
qDZTXTH+w7bbqLNf7hwRmkd7dkKRpbD2kpR+oG0aZQNqUrlaFw8t1H2JOOVJ
bAi4W87J67yCJFXXpE6my8Tyguw2aPImj9ChlT8j2miCcbVCt5A1pV4dcewk
trlQOpqIn/Esk8RkGn7qu6Vmy32yynP18PeBcrclKjldJ1gsDUnKSWym+h94
AJUkjNzi5jEsk3jXJw0lZC3pKAS9v1J+ThyXq1KCBraeV6N2H7TnFKqt/qSv
ulwVWU9OOmcTxfY2kkvhnlGhYtC8GUTok5UVhDueJzHwAKwEtmpJA0dx/pG/
2Y0ZQsJPePXVACykTgWemMKQJcv4w/uL8SpneKL2ER/m8x9pKqf0iKQgePqS
wfidi2WNnQmND6j4ahRD1gBcH7/yX3qLI7PRwZV6oThU4aCNN5mt1QafH6yq
fIlxvgWXMX44b//BJ96jy4AEhN56V9Fjz8rUe+ai2Rmmmv0eqibk3m71ETAI
CXlbMNH7S/iiLAi0FhSUhP26jAmBA5qFkJetJPJXvQ6r6Jf/R4BrUaEDzuMx
nTOqnHDTU/YH5Exdv19Ye51MnZXh1sueT0dKijNM2SZVjb9t5gXeAxFg2T+e
YKkPsV9YYi+Np8XMbUOPSOOj6hoX7Wa3lRqoYR0sJxQDve47DbrXALVJuShJ
jg4d2TmlinqIHv0gBi6CmKvhs8rDoSeZs9YMpP0//8rt1ly85A+6qaCeR4CI
XHnCt/EhoNeZPl7zY7fraVoFs8ZrdVPQ+uLyAmYkeKM2A/gDxukSmGu4PmD5
dgBA35pdHA8NVwyMTvO3+Z7PAuYxRLtdASPAUg/n6LcM/lzqE8F80sfZEbBF
ZTjgLlvWfkGPTQNFdEQRfTIbW7p+qHDjxtER0nEra3WDvYB8Oxaonbz/5tDc
71xrQEnLp6/z0mhVjDoZZqZW0ZYoEGm6saY1mXtatSa9ImA1Fr/YuxWvg/8F
BdCLcI24IntaAlOi9N2US4Yjp0u6IjcfB0Er/eCL44K8AZUJWiFc9FdDQ4mJ
9f2ZoPNwgo3JTpzdzhRp3Wrpyt4Yvn62S4DXBaYE0kXcK1l2vRWtecsn+B/n
sJSGanziPRY/HH+LeYRukAsl/WLwrfkoWCYSnstcX/g3VMZDBvoTedI/df7o
usX0E1L67XrzfDSf23EBQdvLokVm4lWNFg0n8eHHbvJ3EchHkeoq1Sb/CD1D
zLkyIpJgJA625eIAXenjZ5EI1IHd7Z5AqogvR6FammaPjNE/br4Q5wNz9XF5
lSaFA9r0IXzcDxu14sh5dwqYHmHLgR6w9IeubtKW9Mz1YF+RjLL7KX6biVPC
kW9VGh1ZJ9ENd6yq/3cgXcDp9nGsa6rvD3+DgHTpYoUrVxSPnhQoi8ajQOY/
9/M/v/Mu9O8+lkONSDzVpbpurJTHrwwQSK4kn9gNlGz8pQP/b5ySAqMrMozb
gSadyLZb7rgoT74oIdiv715zkXQx2qunkI+ZeCEOFi76BXPgBqAJr+f5iyXL
kpq9oITh9RJsM5Zq5rDeqs6gV1e31emnPc1w6d83kwMPgq6OCuNqO2FOsdTh
9nx0thsfE05nK4hjRosxkWnP5BUMGs2FfD/wtEswAxGcVukuksPsqlR5TwHe
0syXgr30REv8G0yg50i9BzaJaOoo/GOn2Hrc1uVsrCSfFDE2WM2c7ClQd6cp
Cs1xUIg3zqWxiAkpkYRSAUFc0ChwhJTJntm9tLjpTaBB1Zspx920b5XCSlDf
vJ4kpqKCn2KejhnXGZ5LMDT3faLciJQJ18K6Zu0bdSstz9AxqPj/GbqY0B6z
56giSo6DOcjeNDspj6ktSLppBHJlqg76XHIM9/HNghe/24C9EC9eGLX5XTOf
1/09mtalnk2rQOIRGNDxVM9U4YJ+GaY4EQFN9FakeWvaOOd7crjkM69p/B4V
f4cmCOB+eNLSdTbSX7X65uVgmPFqOlLhKxnbE3wZbjjEcheGSFNAWEckPDzR
j26bVj8nqWMd8Dz+7X2EokWp/ou592hdiHuGeFKZMcAlPtbMgBnuA7vJRtib
3qTPO5XaLg/JujKjOE/nlZv/Gul0aMVwOxxBvVZ/dWHdMNm/V+r6+8n+Yzs1
cTa0b5qAEYXn3nyz5U8290u6++k50z3keMAEKidM/ssCfRdwdXkLMXnrxsem
NY6eZJl/6WS77zCkAJlVqyCzTwMt98rI1L/WvCPcOgbvT2CLmvFxUOy807bf
aOi3+Lr12PnrPnVMhcPyZMzDTTSgwkLrTj2Hptxqog8+0V/Gxda92xRy+eqp
Xbop+mXYqz5iQjfs+RK9BrwBCyZnlzG0imNBs5Qnkkkp5DVlessGKhfF+7fu
W1nGrKIZ5OKRo50dtFDPdMsbsP9QV0glqICXJh9VRUePiZS3Db0XPTWjFRWC
Dt4Ss8EDRPSjITE/BclG53XJcAvjFKb0v5UO6FCBrM8XmF05bw9erW92cIF4
V57kdAuv8xwMXinPm1fd3l5FaDGI1X7mqxsz1Ta8vnzcubzLSkC8sSkkPf7j
Zm1eL/b16896gzJ0ARVaxwEir7t+JeeXz/wn27ZkM4thXSMMvjkEQyJhztvu
nN5VEwmfG0ObKR+iw+CSvxv2i3JiCC8UjNePTN1A62vKZOZsBySRq9bS3ttm
EYynh8SAgh0JoQ/oawIJDcApM1PM6sZpmoAaSbKCbjnmMoEWSCiP4UhU+PDA
pLjPS0DxG6ffQn1hB0APEvd0rY+gaGJuIeAq06jM/eRRN1ZRMybkCKTsJPtc
X28yGi9TmqPdOEkVjygUOChxf1bTK+YOSG70WalVfH8VSd4sGaAVaoSk0MdS
CuLghzYgVqTyZH/sENQ16GjxT4Ed+J4jvJk8xFspZrmMjxFtNzg2I06Pr58M
bsPnsuBdVC1QFFyEkj0GP3DWMFwlKM6xoDHwTYT4SiVF6sCEwvQRcd0ewCYP
B+vQhg9EoyePZtLVFUQjc9QOLUqqW7++kUEpgd1FSr3QPkZht6uwDK1lCwz4
wEoLRFHP4UgjwYVW+g6rro3+bij0B3Ovaiuwuz71RQyDOOUEs8AqhMdwuYkH
WT76pWsV0CMEMy3aV4/lMtq3QDp5pwnGZykmrCr39FO23TVR5SrJnQidBUUB
ng53IYMwaChvMYtN1Eh+FN5zpMh5OOh7uP9opN7ZoFFYKhNflEgDcZdYIBvR
5CQMMrafSLK1JeB0m03bq6szJzHWQBTMwMWUTPSp+OvXlLu9F9op30OkfmJe
gdaTOHiNNhsqfVzwccFMuBZVq9w7dS+vLzLIUA5Q1Vhif+HtgyV3TUQIfbw4
bnO63TVqjUI3AL5k/pNfz87TSyy5nOFPVZnpdwC2MTQgj8+ItroH3HVc+DqP
HADrcd2CXEq6apn27KfNmMeuR6gLdyrWF9ZGp9Q1jMGN7YmVgfBf4TdU6xc8
cb0Hqc16Ysr8VqVk/ZpsmB/lY3m2gO+Y/mwkVKTTzk2GLje+hwuE0URiv8mT
6CdT6oZYuMo6hecaztAatY+E8Nh/DbEe3Scixskx0JqezL8KzqbfBYg90Tsq
r2WTZHiGS0S6ewbZWS/Ssk0EKvUOg94Kh5PTEwjD3VDEZSXWNYBjQPLRjyG+
CM02i9+I2TdFp7jL5WGde0kEgaJwcDsencmFfguYpHeuybWfyixmaTuEltik
ReE3w23uEMyOtjnLYZvgCsCgNHCX3ypkVFeNOYBCwjy1IZ5DTSaqqIOxVbx3
P1TReJyVQaGB1s0ee+T5GEpStKp1nIIUXgyMARAua4hf/mTvg4EQ7lv25A12
bSt+QWDfb3lbREms61A/jgzht2zIYxukttkpnQw0INj/WUgu8jHgVbDgZ4qw
CrnZDSkmhmScU2JkFMB/fo6ObdLLnoibnzKvin51i6UX4WutAd35OwbTfScd
4ARcW9a6WXzRtR7v2gHiWyXauqM7nBEbYUTvbUaFVzJXaByH18N6smdEMLld
PoiV7IDFzI6akzO0ULB6WEecFT6Xk1uI+3JzyJI6VjlsEez7QEqOAoSgFu/t
b5k6mNhz1S/NvTNjyD578OZD8iEnUbBAjTrdwbJV+QKEwpsNYHhqtbw1XnSJ
XFuBrCOu8SZBppXDQB1iCksFM0r1Cy9apoIT4XMyNH8q04A+b85iPi1Gj9Zr
wqBlm25trSTcEN8PUxSSt3TrSfMrrQ8rRLe5ULW/XY7nENRTm3v/JWB0H6lU
jTL6P6sfdVVhjqFKbGmYoVQW5eIdhMMNwtJxIoRCx1Uby4yXpITZOR3nR6MI
C3/zAvFhTMnubp1ha/BPiIHv8M7//vD2Mb/4QoOEa6GXKzzrKW+i2EuzyDf4
hHihRfaeAiuOEONuP0NgNXIHTe+Wm5BOaM6j3zdjtAjJmYWK87wK1MqG6NtR
sD9tRa+p4b6sZy7/AjKnVxtU64KH9S8hU5pgDC7Fv+1tFqjED/+RIsGQ5zaV
JOn/gmDPeQhLkJ4+soeyTUdV6VB0Twhl19VKVYdFon0GoZNIJ0myAEyhH6T2
yzEfyGc3TuAXYrgNVQevf5mUI1/aR27AHTcDPeHZ4qQVoSh+GXqQDUurvhWN
bH/aiJadQo8EMmfrrsNv9n+Mqc4fpp8Px9/GpghhL5iUQWYqUk+DBrbmlLGw
NbZE8vZ83OV8svRrCN85R/6leuBxwI0P2Vukv1b9wyBL9YfT4InJXLlHxh0a
ulvcBjetPZx27jXxcxak0bQsGtsUVyS9tvoP6Mr4yEy2eQx0UrecPcIbXlpD
4XSwRjPOEYawWmLiNmq4DqIE2Wb0y+Uo+D2gM749gB8oUxf0O/ps3W9UvqPJ
DAv8zvxiJ04Yg/gDxQvbDGU/unTQD7Nrh3An4ha6USbExPLE96AARx5BmCnj
scHuMVkLtf2Vb6hjPsPfTh4ePDVaaJ3+yaa5F4/WmOF9KlPMXKHI4xul6a/2
bR6qg2Ti7SRq+DQ3awck2+XCokXhuFL8pyq0n/p/mzLEOEo0MNyq65a0yLJA
whWhmdITVcToKX7LjfBY7hNJj/uDlPRQoNhvXyexIuPCauI+Ji/Ur7PbADaz
HQ/2PB50rgEKN4q7zOomWw8PUeTaTxkHEm9fD5XtAekXwTOnnFOMbVGLOta2
eXxPSkSEmzF2ntJkY+YQINTPirCrYvd3emGW0B/sjHWHZmJ3AoTCpjEqsIDO
7hYlOv/9oUxt8z/5Pu7nYGWoBhjPcgoMgRCMeC0lHY2Jl4GHa0EpU+mEsYN+
AOmfMf1MPiRq1wTjODnNgd/51bOiL4hp8O6prVFXcww51DAujD1iiSLNCPSr
Pd+kBaSGuLHHZPJ70yuhZlnrafe+yLFob7PNf4lI9H7lwstkkjJJtFcLH0kV
4FDoMzXROGa+2nPpJfgidqmuoILd2ZcImwGIFuGcLbl34BrIKHFQsUASEnKV
4f5mRA2V5JwYG6Z3m5CqO0barWdDDGnRSgwnxqeSXFwkakfKlEg79L9ScMKu
JQdd4iCRwrBG5HBXSbfOzIMsI16DVu+T83In7CkwNLq1dl9ueVCOJEWFR3/x
xhZ66N81qG3ZkpQfzFkgHpxAXjOaYopoV/DsNM6yvuRQK7LG4Jn/0XEWq3pB
4XTwqprtmtnkEiX8Sb+kEG90Mm8SyG+2CQtCmghhfZaOo196e/21sj5uzbsi
Dwf9eBTuhF4yOHFuAuomtF3fuiahFBolJHYDZ1PIBUB0m7ljfQSDLeZ5FAXX
PzVUYbs3MOAS/N2VN250UENzwkYX9ug5nkAWOIuG/Swxu7XHKExiAaa2bxPT
1yydnPMvIXzMKZJ32KoMdWPi/kechheZ7XzG05jTPqP9Tp2KEwx+e7U57YQb
gSpP8i5ahHYjU/JOKz085FINEgv7trKZCuNR5b1qtOuQ9pg1Ei9wGp7YAmie
GUernA00Rb4WSfmPUawIQj2XXtrvYgaQhf4X/SXU/A4awpnxJ1E8FWs/xsJU
8E2letaC1TU3s0Z9D+emSHQEuQGPuRwCIMOXppNIw56k7fr/n1LwtTgeNCE6
sEw1Vy3IG6fkN1NhIL+ow3g2xogsJswa6DW7n+01Pe+exb2NDkSZT8CqFCWZ
20H56g4M8zT3yNtiWIs/gAuYb9ap3OGHB8YdVWowtke/eT/OH+ma1UJa1uUD
8k6y5fwGYOvaQGrRgr/4YhutVkTWylKMYficT1GWs6tkfJMoowG9dlX/fc+C
U50fszgQ5rWK8XkKMfKDcGO8Gq6SvqijuRLs9mjF6E+VPAoJeKwubWKkt/IM
3KmaccSkZ2W24FVNw9jnZzuw7HC1ONEgZX6MsgL2kXocH+e4NbSbvNQ0pNYu
pf9pA8UNcxHIrMB8zTOVPtkVVTWiDXv8fcp2IIu5TEN0TunNSr0lks8TSXLB
7Hz15ryTdyXFlXxvCeCid6KK1Z9NV2bfu/NIvCVTI3JW8YPG4b9/r0W2Wyfm
BJ06B1aduYiljtUVYrtL9++ODeCjFHgXU019klbW90pN0QZ264nomDuWhIyS
jSBQULap8kTesBAaDD7zAOQQKDVuLulY5UF01ST/XKtPTDeF+Zkff2LTxlQ8
R+3EFxEOuUgqi7erFEZA/x7Zxz4JURD9a/81y0znxSOYORxiWwxwJqRWRwNI
K+QucHbIEwmVRJtSzDr5s67MvoWKnIBcrNEeI/6vtfWJ/dbEh1cFPHto4Jyz
lH2EtgZPlvdySPHgSk4QU1t7Rbd2yDn9KGnPzeFGcBzKOTmkznW28dtRfaqL
jf6Bl23eBZJGEXako3Jr1M3rHDO3SYwdcL7bml/g8GV7JsB3NT+suazO3226
o8EFlcm9Kji2irYRkCtmdBDNqo/Lsa9dmrhauEqYUKbSumzuJHEC2h9aAsuO
sq12s5/3EaQfm8bwKYaj3KE8yd2DERFy6l5nD9lvrPMcqHrEYA+PCtLk9oSq
exZaFYZeVhgpyvpSZkvKnZ2uV/78mr4sr3FkoPRkjW4n80KmmZD8y6LTTIoJ
N8xaJ6K+89lReUAbg+taD/+KJMKR/CSAmla3grgl0+S7xH1L0D1wkZ/agCYN
QXVgmsBdBQGnwmkr8p3kqq2X/KfZFMm5QRnYYLV56MwtLUv272vZGujX4ZjG
1hifCK23Bsg9VEP8DxAX+W0I210YRK5S7UHN98Oll/+noUBAKJJwYlXTpoWz
IhAgi6rWE1FZVDpGNq6H4BaIEj7ZE+3tK3mHP0NIQYtnGDJEoz2y2xOHks6k
qXOCuD3eQBikeYq6YPFAqGBq1ibXwAdLzBTk7RVM6bmdkrXKvn6vLyGvzF4R
tHj6SWzX8pOhnMLYzD/qu4uAMKlA5JpM43epPWMrGPTj6L97RahemuGVXCki
rnpQ+LxRb5Q7DfyHqDH5a0VoBCRYuTQXn27HuPg59h0FeDTaxavOL0OiLVuj
+4DiFJEasc0h4vnxrG3xRTw2lZCMG3UP2fybwdAFSGc8miaY+S3arjQ6L55q
em3AkPLsrQS3KpbA7jGxMJWb0yeONSaWsroWlX2MoWoefKWV3aB1v8tkGVNp
wtQ1M2+kQ3kcJ6shO4KMtX3GIs8y/QRGKBdpt5ulfDPe+ulxIdbplfDmaKmy
nHuayECoH+0eElq6fu62m0eYl8ZaPNb29ly6I+QJLt3e+vOH4MdiWVFhEdmg
qfd7U6QctBWaEoNcgyrE1tlBVyoXuZF4HL29dE8utXbk5t9DbmM1E1ra+cl+
06gioFYW8mtvMLnr+2inDxV+hwRG06ReiWSShLSI+KQUrP1F+TjTCoAiaQuS
RSyy+YxV1AvEdSFHcQheossI2E3/k46evFryKVYhbEuIRHb4UwP437A/lsdR
zGSuRp/PmIfDItG2w5lI7D+JY+t/Zx+4UEC0eBdXW/TQ5VFn40GkHR1BLdUq
xCD0jfTh987HL+7YMlP+ICrps2/8lw4iK08rnSZ4SxL8JK0hRT62PEJSh1J+
WvpGwlrDXZsn+fm1msqrNYroDKiZG4Es5y2pvTm0+07yQKxgAUR1ehk113aN
VSUSYgKKB3yPxAK40PVyMD66MOYG7Qjvw1GdgYlcfgWclU4VGHvgtqYQq+ER
46vd1ijam48hRQK890s0TXjfLnNV1pA0SvWCMJEVJA5ow9uua3S7Xk98KswS
ezZZ8uGGWvcJk1V/BjLw0JWWk6iCwmWBPPuY+SrbtE8dTH+IEr4EOsIu3iUa
8y4sC3RE3+GusXhAhrUU2TT+HDN0jP10nzzcAWUiLbI0F/ZXLQkT+GaMGC51
Frhdc83rlMiOQ+2cESl8PKVQBJrNDTHHLt2tRtLhU6sNPIJNuUrI1pKBmsgg
Sa85RR9a+C4hYMrZ/vLv7R3AeVWZccQfYuoFihr7yOcXbIlMNEaaJDT4kU0r
/rSQ5VuzdrL30x5jKzPe+7IoFTC7Pvr67mZiKsWcWQWl5+B4HemA23O0b234
HxCwCfTfNG2l44fVd8CtDk11DSoPVGQgNsQrvar2I5SKaLBchhzQqiUySc5b
w0diNNglSA0F/QarlnEJBsdrMxzN3IzifpEjSqrZJdz4KoZ4zbFXrpVEpanb
6GmXU7OuAJJhmLiYZTRq254H4+yuhM7UR6ZGIwAM/kfnNe9eA5Pml2Bkx6Z1
C2ysEbhi/mqnNml9MNsev50ODRGPDarU4QhPDNg9C/3iTbNGer4MHRIA+KP4
0aJCvXPvTEmSTwoUVKYxv8lKTPyxzgrRifqm71dAt46th4bEbJO0FbKkYs5c
TwXoxltUixilqIgT7DW7yN46x00mLVhOw0m+sn63t5U2f9c2KMDBBqdnMXsC
dMop4ZX+sovZv0ZY9v0Hsk7Hc0n7mb2+npTKwOFLbeY+nMFqWowKW/7D8rbg
TG/oSX7PIUBi57ad0UntQkbxH4UaqjrY2TS0EYRXstzfdlW99lhJN9aOKXjT
1sjaX12yMB8GQT/fVSQiEXALsxMdfs4ByrbZyr/tRukVN9WAlrb6vS7dNuM/
kd2ADaRyrivZDkuNGiW7CMfd4U0RiLk74UdGaoluPlJPjsQp6Na/XVDLVEvg
YrfFv7RH4Y4YDuS1Ajc/gn6mujPQ9YlZriIkXN9uWu7FTl914kt9W8gNtwFO
cCv0hswXzVB1JYtlLDPub3qIDFcDwwd8xzfpnlNEycaQq4ZXIO2wTisyjXak
CWYsQUBQJHwYOH+6kHCts7L+ydEr5zjgJ2CLnoy16BkCnuZaLJaXIR766549
0tkPaQ3Z+x2AxorSQTaHotaMcC2o1bhHkX5Z9187Imr842MwfEDnvoWL+q5p
kxIfh2+rl3jLBrULASaxdCW4MPBRjFrc8jz+V9YtNfQjRIoqn0kSATCco6uT
rbL/oQSpC8pjjjdk3k5c2WFxNLaW5SOUfsQ6ouGpYxs2/JzN77xv4SOuazqo
/JbqzVY+akm5exVFqulQDkGDa8O7bUvyZ6tMg2cS3F4T70hXzKSR1aFYeQPn
HSOSO7hlFHZWoH97tx3XQ2vYqMPp5UttZyN5XdTYxxqsTeEuEnfOy+GrEOxi
40yyMbVC1L67w2iqrSKoVF3uTpWCuzOf8T2U90ylaRW3cfL1gXYWcEKf7HtG
Xyc/Y4ey+zafZRvuLa2nfecSce1QF2UOWSG0l9ai0i5nA+9cJi0LzbiYKxKe
xgvAcOKKDLWnwX8plCA5z9AoUnQwq9xkKDoWHODOjOmCej91zGo4BJ2bW+8s
HeEeAgRFw10hWKMdb/uJ5wjiiGFmkIhYOxtQm7AksRhhQ/Mqy8ac+N197Tlw
aeCVeWPob5dBTST+M9qCIk7dh+UhpQ+aWChyVecfdor7gRILsgY1GaaMH7FD
+hn1S5EdOmg9zHyyeFNDBw4pXcfN7DYyZ8BjtzXIcr9MxItflntydwu+veQx
OElyo6It8Qpqqp+ZeQ85LLdO00MQl/fsME/HcxV/6KZ4DwZ5vJ0gB5s3MXbx
M4WDRgETYNsHUxPCIG3OlZDbaCeWUZf70dOaMrgJVZuRklbVK1Qzf7haVEC2
c/R28m3PqlrP8/PSVIqDfUoYVLMeTJWnvrSjdxb/Nq88MOFNZ4U0jFZu3ANu
uCt9owt34Cta48Q38UpnYH996bMMd1tbb7pHjbgRgabpQBP4aNn9A4q3M8b5
6TLbUkSg0JWQt5Abk9Lp3zUtiKQVtE/bbqIn3I5xkxs96ZCifJ85XCmgRNvF
f1kSU0I1HTRe7glNybGGt7wf5OG/2MyoSm0iJ7Q4lL8vb07BvjokTycYs9yH
frh4P4voXyReOlAWDY3mmiOZ2WemJ9IHzGy27E1ZjMJTgdOL/3iZcNsmhXhW
J0YBu3MAxodBL3ldprlkWpoertx7B82ppyHhJwi1quOEfHsgG8HzZ5O8vDBh
B/LkGaqqxXkRAPuoQXA9v/vh4uq8COJNFSG4X1OevyM8elCrsX9m6f2+mTEP
J1u6JQVZUDNhHkhLODkxPuYeQr0B61s3pGgNyFED4aCrBFv7wbcyIRvRazUj
63ppnM14rLI6JZaPoUmc8kXc/3UTy9k9i0nYQZsMqOFca4X/kKihe5d9yVlq
TG64vHg95I0bg2Qs40jf9pwpiNSpW/ICo39CZtfehwoHMB5BY3dmnti59oTK
GJF6m/BRDIlUbxOof2OK45GhFndrIRKISzoRg/WETcs5fxy7LQptQxMu+DvM
nKKNiCTF9hti75NUBKwb9ggxYzkIt+3oHlFHDW7Gs0UuM+6lOXjChp09LQI4
YsmwbwHhE7kG5SXrN7NmKsHqY3pA8HuRzrGG6n0A20aPZsA2j5fW1Iwf/4GU
Fx2R3hELoHJgIZyQ6ukCw3xNLGNWVriOFBCyVHePNqz7jeGpyxS0QVthHbKa
ROOb3V0wsxDEFngKhsKyvQw6ppUVpxoOnHbHj4OnHYS4PuA7coDaBLTGGET7
K0cHrDiP/fzHMntRonq7Je5w09V0MfdTCnSED7yluBTNM8YjkPEMAMD/rihU
+QyJAqjSX0jrnj6xdkq4Bt5nlb7weV15LukMT3C7VB7aYmWwLR2CQ1QsHNA5
UGa1TuKnUsQZoL1cPNY2mwPy8U15HCakxRT9U7REubtPk7JwH6RPXysVW/Ao
agnZJgrfS5LSDIymEaJ2+UkO/htvBJ7B2znn6CHzEnubWe98OWtcl6xYaXVI
pciDCAJJpYAcgLpJ7QDaZBMuGvoHjuYoU4mzRcR9N+igKGww4nxEKxevASaW
zx1chE6fU4P8+RHQISPjHDEs2FMU9156xCaiSWG9ApY8cM3/lZRqyicVcsej
vJ6U33efGyKHeb37izznhwDauc1q8ShD1jPA55i8IiXj3F7yTuX5x7V7UWou
TIL/p8uLSLUwvXF6QTnV+FZua5PFhcy+5AxhOQvYW2POnBoVyT9xj+6IYkZ3
byWZIeh8HajZz09gYLPYkLJtGvow6aXKRMKua91UL0tsl57jmEQ8sI9ZQD3b
Njpfd+9Z5SXngA1L64nl6Lp7/mZ7WmI49Xzr2lVRj6fX6tt1Ybw/HXc3MA2F
I3oUWXSttKrfc761aajxT8/cmAEmIxP9vh7ID2ydK730GKgvSEBaxEbcqZLZ
l3L/C7nKUmuLRkaNJ0+n8mXvOjl+PCA9nIfZZ8IBQaTtVNAnQc41AtugDbwz
eoUO1JlgzMyiykvrRjH1c+PEroWaEe/bSFGUa1GsCKqF3Q+EETsHIvlg3LUw
l1txvvycdiwuzz1cxS6i9P2/tw6nXCXRY71rnpKFg1hTuCZky+Ep6Qv3+tRg
ChHVxOQ5r2A2dI5qVmQfU+Gjl7Y48o8Hg/1TZ7AFOJzdWwiyxQCKXjUdf9Jr
t89UGvdSppOTKwZEFLQqzXMx86gmYTGdxJctFx5uFSFBOpPK0ur0+DD75csh
pmFSRMBy/Ug7gKn44axb9wpgaClg1og6NHrXySfMo49uCuKkV249osIi5GS6
KVFRpbHrgN00dQL+uJlSXS0igiECfB43krgHhTUVmDAShdbpObjKyI3smpX9
1NGEsg8y4Ny5gv2aD1XsN0C3hi0ZCpyh9L3CgauxCEEizQduVNWchz8LCYan
r0U47aJ8ZOnlHJRastcbotHCWlYv6SLgnmrCCIZMBwvttoitrZHZy+YQ3dzp
SSedVLt4h/UMFtjtD+ynJX/E1RvDnkvFMIiYkXfebz9kavAQkSYjJACv6wEq
uhvoYAHOTDUzb019H4H/P2LfJESJ6XwyM+h6d76Mk+1cuOUWOYHg81dXR2/A
MkwQ2oY09pP3EAkjmA/YvCZLv7oCztK0ezD9x57TJzJozTwkLLnIc+9EB4Yh
vQ4v/MpFShjMu4TMTIi6x2393/jJPHqtrT0i04mMuhalII2T0aSQfbX//ngh
Ks4kIy0YhYXddJ+TRJbcfGUI9MsjKnkjzR/Lu5Dz8kagPudP00Ppl8d2rK3I
oWZjNytNb7h3KR+ijzzYCIxTvmGcAOWyXFH7Q7STMiFsbB/RyoOBz3Ba7NzT
+gDWs8YQzhH6dqB0+UTc5yk8aIlTHE4z65NO+9Aq4KMt21/l8zWI/Q6mcBM4
hugNJiPQwdr10PbFmTeBBHOpQDmOaZMYbE4UvkEbOQa2XQPACUpqPXxVTc5Z
jNX7HrkXksiARb8No+20zQPka+bss4b8S++cJPOd/o1LuBsWNwawZw8QmLuU
IRWtXwrVPrk0hlY/PVlAkPX/SeJ6BnhynG9IDcEbeAcwW90JmYGbZ1DUYqMQ
963y8OMCrdeqydaQ6fOkp+IK2Ey2vA3AWBGsAWeNLzXQgddLlXfB9H7XwAJZ
EdPMC3t4SBPs0HRl7j/h9XtXYuexT3dsYQdzMCjA9uF8EZeZ8mep1GSQWpoD
yfnYhU03jxRbHgCtozE4UsifmAXCOOVKn/7sCZ/aIcau7FFWEzdlpqB2mpeh
S6kb1OyhWcB/G5BwyZgSgYZEpoqSFoPWkt/GfOSOk7ZnduZAD7ljJO82BxGB
GV5ImHcGzXdPyJ2j9izBRbirddWaR2Qcg93isHdeYC7y0wKp9kei73IxnwcN
BrppmyqibrVFCy07XkTrk5nwm8Fun+Lc02rARQkiOhggKtKvu/i9S8TzGbUV
wEn2Pg/AQmHjB57s8DRHRazXSl1w+/hBnz2HbZDFXDatm7cwlKhlQsD9DcvJ
0yYsj6Xej3oryRXLt/pwuJSa2afD8FApsd14D07PDFCj3PYYWmn3MY2UTyDX
9XemJ+UOTIuYjkwUNsAFEGyiGFFLhgHrWy2L5bNyfLIbWMGMFwjJ/Y7qu1a4
Zm8D44DNLZhGZx6eKBdTgT+Pe4HwaKvKQ9lHvpaAFNkQO1GYi4/cn3KDnQBB
fHg1xiufMsnHGogqDbZKDkY887EFtsAyBjyKzsD1pFANJxgvSlkA6DhEOBUX
A290Hf6Z40DerjaaY7Hd2bXOLpuKKFzNBpIWuNo/HY0S+68+4i8fDCSOkDxc
IXBEpvDRfJgteK1jIbkY14/kFXiYcppozE3Nz2LbscSwEdGYcMOwmJrYUGUP
L6908lnwH3n9th+3luSJikjkmS4MdGU0ZcnL+Hj27ABy/dVPDb4rqzRctnR1
941103r1fv5fsDI9cZMfYOdtq5xhIDRzC5JR+j0nRx6k/pH5nJaG3d8/6bOL
b92ymPG9yP/mSceLni6TW2nyt+lnk0YhK/H79TKD1856EmxcAUG+56JvQMkf
TgwrO+amkhNUpNxKPVIiVyJOBwZUC7ZybxGuldBouSx7/CiH7CAQGxnAZQvF
pSi3b6lb3eAONrn9eXNS6bYNY9u3ctVX8UlNRp6Dub358yMF4pFH1bm1aDQY
HDzrbgc3IwRjBFp7gpmEkAxKtIqVZfi4z/jRMS+8JAehVIT098FlyTIeRfdP
2lKPuSEN3JZzpeylzLYMifVDXu7kzHnSmyBMAJ9ooYs5bkJi/3007Y3w37So
aefQyLMxluN4uwUt8uTx5yiUVyeIiLU8BfE8PMPE3cpr6fUHDBkJkREggIAM
CkQHahasXzlWsSbVbSlXxgLZffAVdrcGzsITzm//tJ45vvSofuOKr0EJww3O
IN1f8ctedaRNX2+oX+AGs57Oth1gbBwWPt/5J68VxezzoQQYwKtbW7x+UCqm
dftcxUsnArdxcUMn3gijE1Knlnfla6Q2ZrF8cBUAEKS+M+B/CDKst7rguLOb
HbxExbzHN5p1DsYXXqFtSAW1SbhDxbi+pkDMscO1+kQgFWb8K1/CYabUc+hL
DMSNAYITDH8SApx8TVozOpqBRGQboa/wh3YBYOG0Zkqnbe3ps2Tk0cZTQqNr
tfAw7lXXV20oBV7Zc63K8MyUEr9EP9soF61M0++B7798CL7T3hn9PF0cqiVN
7G9gQBQLJsYHMMFexny5lA6PuFQ2WTNQEp029GAbWQucbDLa19mXumKm+qbo
38s9e1/hrPkpH4q6jEpBgAj/VRg0F4JM6oOHb3HBGhVqSIBWwIxuNu7sQTPZ
IrjY75QFMqqi+cM5u9F+QfXCyaOSAw/FkHovynbZEKsUU9TLVMmjCAgZRQXt
ZLtFD4+v7US3lNZsXFCpuZYjH0yHAErQabOsXyaohk8YGl2lFX4UbNtvbLDw
32nPuiBNzf4535bVIRN5PtK4FAINLEFfAylmzMYJ3cIbbXpgGr5F7V2bdUJR
TMonBIwpH3qw8nd7zjZudmLmF2swJOpQFTJhziNrOpUXB7ilcr2dsmIk3Ha6
QT7Sx3Wnw2iW0EjUeoVAl5KwjgOLG62v4N6xKZMpiqp/Ty5kNjkPTWPAstl+
zgO4MpRMuB2xRFvOMhwcHm21zhxmlk5uBmQieGrMiNjVVbKPAF7nHSQlOfCE
K8Ue0s9WY1CH3tJ7a782IXJie0QOiJdlC2mPx3dMBNULhnRYkG0ILIzmUrE3
mArdpY+GWZ8PcXqH1NrAhsCcW9iJx4qO68G9LAs0V2Ec2SehZo7XnPOIQQ/K
82kRl5Fba1oVllfQqcfBGxfQ7VddY2DyDvr0Bu6pkAVEES08KIpNgYG5aODj
ccZHAWv48bKLX99tB85TW+4eUmv9OQ0VjbgybfxTlFXdfb+0IBuod8RSuE+6
aXwCZrylcw+37rcpze6JufqKKZ5RjoidDxKSLsYn2epuQHKzywFudRhvTQXS
zvafeg6XCYhgRvHYDkTh16jHcvrkE37YMqD17llTqvRh4N1eRLtHjd/yIP3W
0CZiOTPxRSj/0aA0pJMkC8JYjBIqRjcfMEd4RYAXPY7CY3E3jW4lD8mo6xaE
D6vrWkx9K2NJr65uXtS1o2wvy2Pu8pvNBKGKVSwbftaWBpmbXWKPINw9phhz
e/nh5dxExIZ0a2PnYxq9QWglIwY4o8zWtqz9y9mIhjeSQ/oU96qnjb01iPUQ
5+ve1o8n6zpMfllC6LubI63L0ztzwX8Kyg+Mk1sX9iF/rNpHBf2QGVGhovTR
bZF633LqbK54bXbvzEKxOzR6diY5dCjvgBzCp+ZtGCdsA6tQmEqRWg3EJLAh
P709Jr7R71vVVH82RN1Hy0q8awEnCFeB/qBjGpbCiOkQOKeXOBLwQw8yMk0j
I/ZDjcMB0OqepYYxlUYbykkau+ABA+5tGTCErqouIpGdDKdHmyxKsty1DyAZ
GqlrTZe/KFVczn4dGeu+RVy8FJAMwVIl1Bg8NouZmXV6IZyl+pXj8QpBx4U9
iHs1aygtuKezS0zAFlL646eNcUMroWfUZ/mlg6ucJyMjogR2DYhAMojAhKvT
hddJQAjUzL+/FKVL+h/uHIMR1GmTn4QvMxbXt27tGZoqS//6ySqWAG3OuqNR
UcVLEo9Y6g8Mwo1r+eRVrWvWwlvdTLooFwr196dzkkqQB5bZtZfLHqYck/ve
2+L299ZARq/n0CvDIWqWmmbHBQ+s4H3pjeEYLinIBgOOlpuuyLOcJoPwJUZc
XakNd8DkXKcFndcl+7ax0I2BSyIo98l6pyF7LSKVHeRfxZWz0/c/mFG1WYQy
H4+TRe30WY/7u61HkiV96lOtOfB/F2k3VV7uK9kAJ62CJ+KukMEum7yS4PoS
u5uMmEz9cbo1c9wKtSROT7De05vZw5AM4xdXxditx1hWVcOAn3msfqd/8lTv
jLQG1StexoY+zgclnvWCP2FP4RsN+gZl2DzX6FoQyVgg/orNVOYceR/6CKkA
KKi4uPIyV74INaGNA4xnJO/et0xC6UrRsBGc7zTCutb+e/dK0jO9QSggt9+c
mdeXNPm07jLInUHQfqosMH/LUyazs/Ft7suy/V345CVH9le8LI5Eb2aVvr6l
r4rZ/srfLRFHtvj8zSP78gpgDVUQDYiK3awC/2ohmr1owyN1xPbDRFcAQ7hQ
1XNIdnCGtDMj1R+6G+b6Fyn6Wpw1tmGz2pbGiVPhnybRR/MpdqlhtyIq710l
mWt5qABfE75b5PbIhRUVdDiq5YnZEy6Zik0u5C+EHqJ9h5UB4pUmxmE8EfH8
2KWn+M0RmZU4ndbJrWKXHLLrwi6/H47NrQWMEoWuHp/kQhTsf8W5gOhNc8tx
g6RCPYDK7SmTEoGqD+J2RRvZu7gTOv9s5rAY1OmqVGkEe90WFtBu0mRGH7Xw
tkEr3UwRFwdMyJBtPin9iqpzeIflxTCr6ht+uZclAuGjvDv9GjFB+ST0NWuk
oPISqlcUpT847r1rHbIzZbCsWLl38FlJrBjpBvaSyGw1ZjqzFeHcxok/Skf3
eI/rZ35N0fTaYJN8dbv0YaOKa50vnI/55dJNcLVCsYX1QkNz7zCD2hwiHzH/
hyXoipJ5JkpZ3KAY7FS7cLJwS0QWu5LP2WU6B1JwKPy17SRPGzx7T7eZ+jpn
NrM2ZD0GhEvyLmb6Pq6kvlinr0uRVeoi4ffJR5Q21TtrKyUrnpVtk8Y2+6lF
ZtSoK69kCqWPsns4uq8aygnd+MosNYMcVvQusKUayRI8dpcFeT4pmC9R2GP3
/5ie/EaYk2D9qxv3XzULRiz3trO8rwoSb3yKE7VpYUGZ1cqGVH7eeaGK0fvE
l43GcXLzPnArVchMw4xOzBt9DHL2jrk4jlXyC6jxVcUKYGAZGp/ZD2cev+YT
iPf15gcPMOUiZIdknBpINDaRRkyV+EtsqQ9OEblUeNH27Wo2UqtYBE9Q+FO3
YQ7L/31LRpU0g4e3Nt1vpFr29MRrZFAyEu5+ZEDomXuuRxlh3FhyxPed6cHN
TOFPN9PukmSeBdXi18BLQOxfvWPJV3Kn3OiNuGR+LSP/3bsW9yrqzqCV8qqj
Rj9BvrdxDW+1R1ph/9TcVbBoQD5cb0gmxq3uB3qr56uOkfy84/9vYTY0Z+pB
fcQ84UJESuTtWCQnV7jF0J+5o6aIAKDER1cCI4Twg+Xr1ixRGsW3ZI0Ty2zW
5hWWKyjzfaWO4cGKGzE6a1UlEmnuDAPu2ipkuAuMqc46GrVjuK5n1p2/wv4h
DQkFUXOeWY0JNKURH0zghkqW2FIU/5n84jGlNm9TUhRybGyPxaisUMw1E5jH
px6Y5sVapQYoWnJGnZLFUaSbT10XcmJp2tR2JmTF2RW+IZt/JNEUIyKei/oh
ogj6aogpVD3G+lsFvLwS1+DbigJ9893P6WZecc45mdYSBFE6P5kjWFGB6Nok
EqYLsw/1lOJaMFoxdemvrPdY6xSsVXpJ/6bpSt0n0lEZOszxA7fCU7z0pgJq
anamITUWm9meWFpk2WlZxmDAVm5+6cblx+Mp8+wZ6rU+cJ7pSUoAfQzng1yj
5ItNFfrjz3tURifocqsFzz1zYSh+Zvk2MfeQ3iSvJg5RMwRvQWF6AlbU7SzK
MBOtyra2PKjPuHRBJ2e8nrkb7VE17zIzfltrv6slVm394tRjBuPBgt27//9k
3IRIqfi1FLVBr/7ZnXnJgqTHvg04FgD2YlJXJCscN1hqQQiEOqNpjpSI/vbq
oEnSV5WLMVsA+LzNoe7CHIvdmmdXSjlqNIw48ZhU2vovjY9reCAV0miBpYWs
tZKO2B96u1MJS4TU7n66H0BSq9SUGTkB7K2uNMK9+AgEVtPMRpJ8Fg4wo/df
N/qI4JUm4q2BBjUu9IsVZcSM71bowmjQ/BtoliQ7pMJPzyrTmI8/Y9W7FPVH
rzV3yszDY5pNW/YRbwwIoPIm0XHBY32f9gA06RTHcev+GzCkfrDXn4ZcP7SR
RwOlP+4Ls7iAHxetvKePxYDKYqoBgHhUrVzv+30eo9SjjqN8nfjN4bQ5d5ef
YAxt42SUyXzT9Ee04ABooV+76q7EMxGZHrb5qNoTtmWDxCWE84XkSCPa358X
mk5NJefMPhnkussa4yiNYeV791SXbJs+ve6jVrO27F3w2ljESjmrrLkj/hfb
8aamyRpME2NAdlwjrJd6Xb4dHkWUju2WDXTrPLJxue9ib8jgUh/AIeAJ27PH
2xzW9NQY+iUe02Dwbj1NBxUkkOe3iqaoXQ6dQCNF6z5uLPgxP9XRSCykYzOh
qvGASbUpdS73s3iDw3uhLCAKQjWGrcc5z33KDCA7x7l4z9irfyVNTL4U7fW5
myYbYBW7euJ602/4hFYYRJoV5Hbr0SxTjVxazq7ZpclWGtSU9aP1aQz912rz
VNoQETWAOj8TpWH5TZmGNcGX6vpcraJvI69KWkFE05J429xGTf6itRf8xlou
ozB8fTblT0xHPBUTM3MBJFfZdhChHiOuMxA1U2vyMi6nUgCyb8EFjwa6Z9AB
pmRKyAspVRVxGp2/NWN4mv+VYiTUpoaYs9LypuVFbQVgK/rjxhDRPJKgipEN
QTBzHW6AgHODewkg2RG0GW5IP7Pjhinl5sDawEPhIMKbIB6yV78SScAaf/1Y
2IrtxKc5i673iZXvgKi5L4Krgo2giMtCeJYkDl8uKTwVJfe8mO9JIPArmEuY
6wcWfONvqfQtr0PP7g0Y64njTvKdBTaNan9wdmtd9z0Wduq/ZY2rzFc6IJD2
SWLKF6IDPayZmbCaqrw8wXQZkPF/h04BltXR7LV4cC2hcpuOU/2MHSko2eyV
IdLj2TQaAuv1RdhLNVmN4tMan+EoV3qKeDIVMgFnRCNhE5Nu29lt2obpzsrU
osLwCiLCWDjsSYqVR0wg1toXKHn5V54cROjAlqBufSEUuy03mEnvaolHc92V
sS9FqhtQii/G7f/YkzVhvKn61om5qOj9jjqbsoD1KBReN9KVNDx/wd/cBztv
dJnzw+r50HtrQ4YN7pjwuk7qlAvaWCpc2WtCwRm+W4UtrHUDUCaYg2agie7v
K5eztxhqgBbyQzUt9zZOKg5s1M/0Iq/B0p44aAI4ZC55Wo8zjyVl68DWBZeC
1D5UfwrFHOOwE2A59Xaa038MInQsDEIUmB45Pl7W1DDvRR8VF+VRFZ9Dtf7u
GbnMfVgp0EuEG8XKsaT1xdaBt4R07o1rlgeIjItjLe7odluk6RzuphVWP7ud
H4ZOU9uoaQQihVqAIuoso+5dYmEcgA+hMZgX2a3hY2WhxJby83m3QcO+s82l
ABjEAo5cw4Slum1o51aoXYPGT8OC7D9hgIbWrRyGd8TZ5HShikWJVG6FblRG
0BsLqWVO6/ymfH2oQzzQYJEACVBSDCQUF7kBWgOCG6x0CxTYmKghIspOs0NK
oQPzLE3GXXtpq2IPPdtHZLCG5btrOMk5Xq2vQZ/ZpTCwimZUXjMjq9ubHfKe
pEpVOCspRMwAyoOmVgVM+ma4/FydvC2JdNz5dQNbi4pHhElt1fdWN3aFSElK
yMH2uiwUU6ufr8zQ3UUibBocEzf1/boxzolgEEfozRa6QXdzWpFiHramDkaT
uJU6Mb//XK8kyKmY1Zv6FJTHrphQtjCjmzKx2sTQB/7iFRcO5nROjuN5i5oH
atI7PQlVeW87q+bYcmBpHiSsAy1jkjwMQy4kxLWXuP7+5bsLlRqodoKfOPLF
LpCvN9H4vUXdynuUU7tziNPFQcCya1Re7WIEm1gByRAdZeFd1Y0sQiOxJghW
MSLHlaFgUODuaMnBVIEBZGpN5xDFZ5n9VCv+I1/iDJJlZDak0+H49PXdC60v
wxEn9woGDr1SeHq/UpXzoCNQhBYfJ3b2U7HouUxGXZWj9SDEMkrWP9etOkzx
s6gZNyJ/e0DCx1yVAYsWEJ1kNmcmJyz7L6/erD+KmDjnG9OJmPjH/RZm4rdh
0mQniEz5cUJslAbWYu4ItuDbzIbwU2nJRmv0wIyD9Dzqun6q98K2WA+1uE61
MWchT15PeRCWhzxFM/DKmvVzYMhKH1r4oqqQNynIClpYuwktFuaa1AC1DL1j
Y+70nR3YoIbsYwC+RngezALDGeICxTYG/n/c6aAL2esT2jN9X6NNxrkNN3Ve
TBBFeFc/T1F9rBunbq6HM/VyOVST5cD3H+vK7xNnfUdklRCyA8UcNtUCR9Aa
/7NzOWvI/lX2XIIe0WPhznaifD1J3/wX4nYxyd2X0LCAsA3gwvhQlj7hRm+e
IaDde+LViiB0psO8L5oNkrBsaR5LKvRJUY3Igys8BTwIdc53JRnLcKBMfk1R
IGU5UOIOlEeN9ztQt6awzJkLSf2E2JALmss9V6THKnvVSUEPbnsqNUXlIIro
lPgSULi7tQfc0v+AC99KdFZy1e670283Dz+y9mlABiL05iluDS9t3rRrfmud
v3JU6KCGtskKWMihQ/GWGdYLgGbINowE+H8pcOvx+5o2etgAKEkK6/pBr9Y0
2PiedoGYPutHNRpFJ5ZsIrDfhneZYaq/FPdk7dhtgAJS7Frs5auidSwGWaFX
rlxQOH8fZD/6P/t2T6MSqe8OV+Ytwwd2kzTC29EsGc+VAJVhdoZcBzQ2gBMm
4qiwNYsgRxxmefppfq/Izy83AgkMCDqTJEqf4n2H3wdN0u/om5eCBZE5GTQg
Jvqa64ENy6tzJYX4B1hxa9ZMjtQXT0dma8QUWj3aQprXWw9wVwLJis1qh1vH
9CgU7BVfRNHFTY7/qdE9niKMMAxUBqG7RRBf9NZCUphRnFvd2L1eC8kHs5Dd
u/mLa+Me1lByrgiAYPA3gFfAMSFxl3B2b7pt3E0KuHJT5oxMMp0VTsbxLQqD
um1ZtbvgEuBjBngpnxtLqgb0vSVRDLXPo1NshYAHoUNRaDCH3QXoZAAHOmfa
FUGuROsVpqoQeXgwAoYel85OdfRRBRcUTkJWcu1f/9BCz6IUjzPT6SA9p40R
KZy9ZBK0XTP8iceb6OGc7M3jPM6uAzDXYdL3WCZRsDC39y8Jyg1Nm6xPDfbj
WK3buQT+6KmGFyiDrTrW6ZucxXVTLTDITqPTaua92/A8RjAHHRMlmPiPSdwg
v+0ed4Q5mKssqmkuB/bhc+DXtMuKxYDof5MtlQ4KvQSMJD9Pw7KvRMqIV0IF
/qKNgNk9K8fUSMS2vX2ASMaB+2MDjV4piWfYAXCXGwMmUp5IUR3T4VfHLFD8
7rqkjGMHMoyogA36NFE56H6LHNqQk1dgzS8KudEYlyAWAUZX0ly+IavC3QlF
i1oSY1MxzhI27fVhLRHOd6nZyIV0PePJQspk733wG//BNOjfbSA7fVJQ/DLU
F6v7ISlGkuxU0aPvj1N8Ldq0nx3Cz6p9X/JFs2tey3ytzOCdBQV7HCNCKPMy
hldIJKGS7KlJsmSa2T3mjiZ9nylk+1kR2aZ9Gidsm+RaI9DIQgtvhFdwglqu
MOz8jBosfNM/8H2l931ecsTT9CyN5gQM2w9mek7j83CnWmR1dSMO/YjUzHka
bF62zcg8/M9TFy4t9mejmGHvOWKPsdqjZOcXBNm3FpVdMrVd8MUQqLONQ2xF
3cndRKhLp7Pv8l0w+sYHKSB2wKdAJzBiwoQ6Mpqg9ZNv5JLh0EZB11Yme0e0
ZWFVmP6CFuJ/BB3JPZf48xwxdOpITuAo6duf6vaDHFNcAEIHub9bmherahwl
Kihh3R0hAvrAalHu62HxC3Ya50YPK3BATcRcfLgJBDaT+1CVEwKp+XPLd8r7
v1QjnIfp2v5STbxgk6cvEaHsR8XIbxjk4KYkPwZ/PlPozxD4buxaReptAn5e
W5Msj+71e/14NmBisA3mINKmh0PQ9WoL+XTFLVP8hobo/yt/toE5SH7HZ4gI
L3/I/nq1GESCE0AwSCi8nyzzErypch6/FswjwDGARBHhbvDp/vNE+WsGqlzC
cBWTqqOeToqill4b36d8D0r7jS+5o59e8HGO/9ObOBs/ytUUMvsZHovCtp7R
neN4JIJqdC52GoD7nLbWxosUYe0/5fAFcoFGwWZVkxtKOfzr2Hre5TyZm7Zl
A7CEEJi/coPucGny1Sv0OcWdc3g+n9K/4KPIS5VjTXODj6T1DcxmZlep7Xzf
rX98kr2d1U+lbgN4CR9+9dhpJ4VX6ExCdr2tp6UBoZtapjZZwtB2BLDfXQNv
ZPvSbupUTK798cUgYntXGA4vyliArMUExI4fVlgqlkMOvW6JibHH2udIf4E+
Olv4CKNfRjjZfrbO0LiS1jcclJLn7Vh/akwbyL2bHTmmKZl6HKIdqtokVwyD
2/Gel+HdOE3GdqTCtDJikbii9ahA6TsM9vcM7imhml2q9kiuOA9cuZpHOExE
15tuGnZToN/kmxmT54R4SWeCdl1x3/ZTZ8BX7i58lZ2YLrlW2zr2RY7JniHY
lw4/ZMK87BSk1J5gHwyLJ+4dtP8avLlR1wUK0K9GkwTcKF1y12jnfUCqsYG0
QiTvOZ5twg0HwHTBUP5udk/77PlwY//kVlvN7rnhnLa7PYU2AM1IMbkbwo5V
YwZRApe5eY+FsOwMI+MgdhgMlAuDTHnbXCZY7rzPdamE+JgoZ+gK8FanBi/+
VG+JIvoWzGDXujyzl21c1hmGBJFU8aGsBsSQe0GxzjDBKnv/TwYMXrUXJ/GE
BoVjDUrhNgfnjxXK/avknUHciD2yTr5XdLadaaON9mDO3XX4a3G2PWiwAcp6
vNP1yGZ5Ss3jYjGvUMbBvrjVVL+idouTPjmjC4g/37lGF3rg6OnCNfos0BOf
P2a/0Kofhg0GSRNbgfooWOMahmLuIFaS83pYCeUotvZujgL8EKQ6cGxSHZqa
vWbyVJEyYOqRbVDbTuDlPUNHFKa24zI0XL/m6CGK70RYTIJqI0uk6sHYQcKh
yBD18HPEB0h13dc4uMHD8QEIADUQsNaH9dimhak67CPAN7OUUHioHN2nyrs0
LVY5imJ7hCHGWGFQmMdO3GkDBddaQFz5TG0y2oSRoGBAc47iWK2Xincu9dvn
gxIyukA9RZq07LTpIYYQoMU0oGIJpngQ74D1OBQphK+oSRfkxezGRxt9WeUK
LnHw6dgKW1Wq2lcCFfM4FnSbtDfXCKp7drXk3XkrmisntRtCd5qnCHwuceLH
dCxW4nxwIoecmoOzm6uVE+bF/iLPKpZw/8OLGmtdSo2aopeVkCHBTU7n+dRq
5pZ1BEPuOSo5SnmlOf1lodUxJ02GjW4ive7lzJUwRah/YoEjl2Od4xaky2JA
ej03yFUQYFc1UwfWBAkUaEp8/Tl/xNlZWFaBnWLKZKmyr/Hq/y6NlK2xWhdE
vuBtR7Vt5ZFTPObjAKsew1uI4Mbt8KYMDR+YIv1Tf7elB2NIkwsMo7gxtIPF
G+B83ntvYfwtQb/s+prQXj2uTL/GrVCeaciOciJKzjh9g7g7Lx962eIAVv24
PcF4624WezG3TRXe6I7sd9FaoZMrrVtCeltTGVQtkwWm7AgJSyE4MP2JJolO
0FX1FZ7veU8954BezyicinI5Luow0s6oeY68sld3lyjBwWMODDLLGiiGoqsv
iW6/aUW19vJrXmBH3L+KkWVvCdkxZ/hr1aMUX7EVAei2RXQnzm3Sha61x/4m
ggGrd4FStjP3ofrM4YdR5RWWw0Av1HpcycZyqhhsflIsD0pVhmcNOH+MQg08
/lPjoCahQFZHq4yy4gRUUFoJwqPzvgn6tFs12aBNFCdA1b/Vh7ROwYub1RWI
P9XRvEzrhY4J55iOt3U1mYuKRPBbR/b/Untrr+2QXDoyuiebt1xx971aZgE8
gqKu8kn7/s8CKibogAeWdRge3cxDraJcBzyZDRgasqmg8ja+D5GPT64VU8Qj
5T1Cvb5BE6OGBW4kbJ80gnh/o9smEYCjNeykT+aFBZScT6NAhUtLUfQek2ON
svXJhDQcvAmUypo4Lgxxvzban+x6VS9MrvmiMJ2xCQPprh7EEyepY7egWnK6
ZqakFhUQVZn092Grjqi+5hRGwzGErvWA9C/n7D16W2R3sdZWCp0T8XiZWjpE
Eewb0krT/W41/fpxfl9+4sYNqfRlnKA8wFd4WSLbKX7D2z2L+ptG74vGPhQz
eRQcv8MWmFI+zZcs6WYnMHNfztu+vC8FB72GS+wrkuCYZCu+9KZpRfMwX0Fl
60bhbnFOprXwhVor/yEJFgKUempzwrGtCriAPxtnqQLB9Y35WzehWsmrNtE0
TFWuAapMoMdz9htmD129bahdgzuR+3HTwUWJRk5tojOCvtSmd4Mh9QBZCXYW
IV2PLfqVziY2pDA0ceYBBrt3Ur5hZf5kz5S5+WURLN72Tsi8410uLApkfjQl
AX+upjYtS473EaDRpT9Hl8SPyjaZ9cYwFaC2V3MxiDqOU0u4fvcIZg6WUNJv
SMxiy0DQLrDpRxzyR3EIjZ49kELkd4SCNk3I+p7XRMHkQXni6NXEUB/Rnf68
6dK0DcK8VFDTWOWilx7z8zAB8Kk8iZkdaa4D7IRr0WtwHmocpy8zu81pRJn0
/7YAvhBh+nnFNc46LTsdRKRtlhhWsItWnPu51tJM3X7mmZ5MAaFj3pOo4HTG
lx+6mEmfmstEIZPnEl+oLGHOJHATESuiDNKOWAFtk1RTBg9oNkO+Dk9WECgJ
L47i7+uh/+QSufEQ2lY1TSVEESt5krRhLRnoMHevbjf31NHh9Tt2HJNCRPmw
AT4bytVO2myQfYWsBegh9E3ZKVjMrXETKEpHTt+b9vBgaSqvKsy8dbNf8wTr
gcgbMfruA35jq8XVEip1TM41xbt6g7N/BbKYjkC1fPtACZ8/F0EjvWxKGnbR
opgVv4QTWv0KcDjxRDhkJGxsUPKajGE1eYx9BBPtG3nrrqDGhR0gD9bkBkg4
7hsJS2yqfHqbaUmK6e0gi/qKFXpRE/otrzHPHSzLGCi2DhJIBE+NfwTTEq/a
1UEnKmam9UD9Eb3BAu/XLGnwSPvUkufC8oeSBR5uw2wXQ6+y8KnJrua+PHWo
IGo2U+7VCQLRddnaifeWuEXNo0XO4FlpL5ejYUMTT7Cr3v66hw7U7QG3y/b2
R4OUWh9msxXbT5GDFuXaIPgRjYYROCet76SXesB+yFk83CTjV7PrseAyBrGm
1faMi5mc1UW1D3ZbXDvdK3uT4qXkd+gDeK0jlEg/fC926+Z/ZgJxBHTrHoHH
UJmfWow6FnhginfCvsrDL8fVT4paMYCP2l4JeeDiyF7Cmtp/S3Ukazl3fLhJ
3kQqbDDK4HuPwfCUaxwSjrJf1U3zVfFGTu49l/V2Lg1R9mOV/CjS/qAoa7Rn
jzQNCD9tvIyRA6yV/wC4dpyAdK63JTCOzeO1JegxQgj41vMm5jNFe2JpxMKp
w4ZR2N0JHTcYO6WvJ72sFmgex+kL16L78aNVQI+07E0U1/XJ/uFNaThderNz
XvILUyLJwjkvxmykW6fgI5tO3GmLeXGqKf0u9vwTWSjsWVofvn5IEsqQDDxX
EPcVtYIZf93eBEEo5jYpd1vEi/qkG2YZrGx1Yu22kRT85OltY3SSQiFjSzuP
iP91HnX0hVJuToPmCW+LVRNth5Hp03o/JtRLvySGcr/Evc/BEZB/SsUUUNCK
ojqbljJ8RUDV9p145whgxRrsdsCARW1FQb+c5iYwM9HbIozX3FftQiDiQf9K
6yY9zo+MWixHVZCqAwYpzwlOzD2kO3pCh64ke8K6btq6Z2mG1vwwIj7ZUUV6
C1tjjRymaJ7k163L3SpVhOsOJpE62zJpxYcEeuFuutcEmXEjngygLqG/6orT
f+LryUqTsNZ7HOn2ozalkdh+53ataG4XGg5kJe6nI47F3Dk3xioTZmMJMvMC
3EnA/EMGebLSDBVY9/dIjlpIQ95ShCelKtI1ZND4V/N8rvMrF81ptvi3i6oQ
Pmqyvsz8AZu1PvxetMMfQODYGpkUkSST+wr+2v2sfeTuQnrQrpY+s6d6wCTo
9B+xKrc9O44/UPuRGdyUBs0o+FK3B51VfV8iWR2j12k4yV2H9ieRo8q2u1Q2
Cq5N7Eoq3q5lyNE0pRGGFY/xv/yYK7jiy2aWRktjgebqtKdl9hSxutzHZN+Y
1jmzKKfl853C8NWteTjv8BzkNt3cSz96ZBFcAL9LEgL6KFzkGcbSBpOeYCSS
81IkyAIq9pfdP6CKilgPMdat/xlrmCyM/b62+5G+b0u6XGj45r5WVMgvndRI
1daQSvlhRPI6EH0mq6cSj2QXeFRy0QgCMFIaR4cRpaYJakef1sefX28ylDH2
0Pb+OmeLQQfUAcY28HGGvvvlX44xhS6hONG3bKYlu60c7ZZqliHfM1IJDfbc
USpiJpecUu0A5CGmavbA/QwOnQI+98w8ne2+6FHfB/sm42tM1/tuc8VWLPvu
7WTqP4LJZt2kINCMgjZ2aWUH3gsK02akIM1P3phvYOqCWFp5WgeQyc2sYPC5
zQ1IQJ80Nzw9rx141q6olA/4D7uGR6+InsKvFTWl33UouO7iGwh8vFCMoehk
B64j+Ot24Ie0foRlpQu+cANXmt3B5/7FRiR+cZqM6mAXVl2I2pyWp5phTHJp
dpB1YNS3421DvOD3XcadpHlkdmRwvXFDEcTuZdnEnRcOnVA3Rg9/ckYMBsqh
OLmz+40nfN04IN0jbIy0tABmxg7An327nvuLokO0uuP79H6V9Xk2G/rux1rY
TK/JryI7iYmFnQngadp3VuakaUeiMEMpS+P4ganGTrX2AQjx1FXY7h7Xjq/8
WB4RELHFIPFS20UbdIgTAxS4RINti18wUeajA7Q9eClv6no35xS7/1zg3Qjx
nNPAnvnd6F6cfLLAGAfx1Ct7YpN+0eRozCzmjBqC5XBBpF+YSWctMDQsTTuR
WAwndkUuJiCVkmNpRjQP338sUjMT4eEgNew6vhG8fhOwrWtRnmz5O6uyZ9gD
bmDKuwjO7w8JL58VGn1FnOUP2tFCHryZTsUUMNASWVnhMxnre4Wqvw4njIHm
vCo4ZXX9VePAXglcZHYtrm9fHHpYWu4GBPOeiOnCtYI2x6IuqSiPjVBgRJQI
x5p9OEf9X9A+FlGu5kpUARIkwjwQdb6jSNOGBkXkscVnbrYOYqp21MWMBv0n
0pw2SReh6acWO5mwDeXPL9fLyv745rYGQnt2ltDLUYN6Mhvcrcj3flTc/BR0
6BQ/Fh5rqQIToNkJH6DzRbKqhK6Eu+Cq75/xupMnNQtEYJQ+q4wIns2/z4F9
s5/jNFi8JJBYvXpNSlY8pJoDhTl4Hi3J036VPZyWTR7KAf1RMBhTI9i6EBnl
fHHf4BBjz3JIZZXfbNzZmNacNOXLVz3FZSA9zTpm5D2xsyE7uUFnxbqf7oTX
NTrXag9u4NSGs7qmlO7di6TO/Hxo4bhZ406qYQ3yt9Qqi07+iChCQklIXEab
k6jfX1r1Ybbr9P6e9sg+RA+zX7KcqrjpbQERVY5nyZmwDvuHtnKw+5NiSr9n
KHjCZLdGvzmT2UXhvQTwWg9FPjrB9NunVoAoCwwwEsvPrTamUy+7LDsZGqlN
ok+91SzatuubBn2oz+mOip4QeBZmtilB/uzpfoYUFN48n+SsvD5ypQ1IlMvI
xc+8tv7iyuJqIpvgTNqf72y4cmZDLMYXjRjZpjdwct6Tc2pODgHzuk4jPSip
iTBY3jWWPGRkj+4NiiZqUv+GdL5WRJ2QQrv6yYS3S/Yg5qar4xA3YJ8fnled
o74mNzr/4dv/AD7IahLqfVCDdvSP5ftnDDGGJsPb+sphoUNZsn1prsszG2t7
hYP4l+i1VuLEG3srGs8S56CBPKAvxofD2kqfliSDbp8MkE+iGficQj6QCfrf
W/HBrIwD7JBm0+4S4wjHfKH0nhW3UtLgP4oV6Nw165CstNTPovaZ8PdsMirX
uiKZQcVKhbAetSUkIYbmKcKCSoJ8rF22sSGzh7l0G1szXLpjPO3FwlRiDA/A
Eq5QiwkkaEVfZDTSbHMKES3Yez/sUuYbunhJTmZ2D4T1JN3Vd/s1u/C6B9g0
qZnHF4TlaFJSHkxgTB57RV4D6q1Stlj9lMc9iT28YZ8j3ksbhzVAIsgGKTDx
/wMT+hyH53hR3oPeK8KPlDbi4WZYsEk2PntbX4Pfrn60SdO7wyjJRo0+w462
BbdHR7izI3ttI4DmC9uWegDdf3sHeK+i8J2LJIGjIF9qkLLLIle6bEYm9Vmq
kZC7HeVSvtHFLyHI4itkhvUiroD4ElUTij/ojz2Uos3w56aFiAydnQV3JsFp
nOEOHmlNS8+kyX2shrJdEox4C5NimXxIgSFKlKYJMW6LvZkkzfWyK5N6plod
6X6U9X8lfmb6gTWKMoRSj7leACvKDCxupmB7OISLM6mN071uPNKwHlDAASAS
11USTKNH5m1b+/bn+k0cgkbpcJ3WLT8ROal1GXpBKn6/9Sw2CMmzWT/XJVIT
k5EQpWVz2oOlBkCDieYg23Oy6ic9Gt/YJlDg4+buLsEcGIIeAs8S1dRLcWI3
Talyv7n0InlEtLK6fJ6cBJCsneWQIxYuF8og50B0zpFV0Buvs0TKuk1hPFjI
WIomivV7SUzhvdE316TOYVL5HEVa+DBANAC5lOJF+NkTNBPDVcZdVluPtDs7
8L43ho67ngkejhAQDbwK6ZDPmE8V9BawgdusuLgrtInoDfuZaexgVXT8T3Og
yXN6TZNjCsrdEf2E1BOkSRog1ee4itX5mSnGk8r6vnVP3WrChKsG+qEw2S/0
yiQfBdgss578Kl/H+tAWKkZBeeO43GbyG7k4HBm3+YMwIjeWGY1yb4/+jRFq
AAEUM46rBaPFNjkd1nJxiyozOB08IWStwSqAPgkPHThV1WpTvKG4doMyjc/t
/DMqGQLlCMz6buEDS4pG54Pgr4RtrA9k+rzjetSewsSa4kBEw9NiZvVxdbF1
Zk8Dy1JRzm/PmkADN9jiuDNaBKSvaUF5Js1CIFbfGijNaaPqBQg1leQRxn6F
wFqeB+Y+18Th6D1+WAp1x3KB3Usc01F3f56cKFz6nQaHvAkImvYiwDaIrzgl
Re61qHjWLVH5TAcd8p9IEOx2ELHfaxjR6fLr7gzJhWc33SfSa+MT/UIFBx6V
DWBk52KX/ZMMB6kjBesx6ewGkRBR4NCPGwfkUI2buEHSzO0A6f4ijLNjTnMz
Lto8TI/l54ejUa2SrVtN0b4EAE/1jXOFUWI0n7CNmYIs8G4Kc/yxSobutvg7
B4cGpCycLyblAo+3aDQB7ksZ499NkuywuWU1DhdPi9JeUJMMWv3/A150cF1E
iuBKIks8M8EmXmzCsh5fxxm97cJ98fXLDyMZKXZ2snPseB3EFrI7ifWVKMmQ
VKPDhoyo3Bf/A9mjl0oZSDbrS4yctWK+ysZoqBlkwlaDP0gwGXFfXqUdpzBO
yam265oJpsSeOQfiN1mjAqfYgmS48u/7cbAKXQ6KOoP4SIfxamgfx534qJuU
cRKTjsF90MwMCI/DlYF7hNWKGqu7yOf2MkQb7PNcc3ImYF4jIN/Eplr0q3gE
935hC/MD/+N0eJRU7EslrC8wtR9WHziwyJz2Bhkdfht+c3YodVsAP7itU20t
0guq2sHxMZJ65p15LkQXHuTtprlaPMormZuuvzIafAjcoZhaLO63MCIx6+LL
Sf/X9IsQlNpHtCqK18bMDPbLhGt5XXAkSYmbR8QQ+YcoOp5flmAVp2VLbX/m
KJ1U8GSrGgKQYry/Wlh0pRqiSXdmUPyFwlGyBGjT3Ux1z/ZyJTrFzNQNeMOG
z5lS19cDB6GAA7Y096TM5zBwgXWLdNtW7UPE38Nl1hWt80UDUt2BYmZ7eZDv
n8td1dBp5kKw7aBytroyovBGpJA+vdS4zJPKYewFB8MWvZ5GItWmTwCkBtos
5qLlBU/BVWbHZerB25Rr6Er3hX1d5Mh05GNEy3C9OHnXOOtznlYFV/ejPNpq
/1O/oQvHJA89vfV24iO7iiOQeTLMrYLMrI+0a2UUeaNs5eVRXymk1cQbGNO/
ZcuFsEaG6U9dqY1VJu3OPghN7wRdV4qCGe4SOyXvrVqbxwuSoloyTc0u+z2s
+hbmpPJg5EmcEb6pzxJA+rcZy4sH2XLbuDedi4+twjUNgnNdo+SgAfFcOa9f
dRJgaVKT1ACPmAjUiqRRzPz9VYaMNHc69drxcRiq69cewYHj7w3NaOERQh2v
QQQQNbRBp+BTIYI8pB663ZKzOt3vXNVLqA76kqV9P0kKR6WypEmm2Sbu+9A/
Mckoa00nadSO6uHtKc9aK8u77NwCZztpSq8exdFrExrEq1wgN5dC806khMXv
rRWQh9swzZRzekJy7O0wA+c3mecSmAb6mu7fFM9ccAS0NV03ewAzjIkkmUDm
inGyvmzHWVODsdFITqCljo0FE+ub9b/sQitoroNCu1+DuRd4994q9rZE8aNh
o+XWXydxb8jcICRrW3zPj9nk60ZDfRjTV3eFHFZhTD+QYJO8Om0YQN+NcNx9
lAPyv0DjkNF16xEsXuK5s+zE1ESTKEFzzeA6EO+1K20kavA1ttYy9ofu33+R
/fwT68rVjRxLngFfGoC8fMKXVG/+/mr5NL2kN51gE8lTK7D6YR/Ooe5muJ86
3Nq6AI6qWNfa5pOFbvLlX0ETxn8N6CesEIlXS+NTWUPfDe9f5DTNZpKk93m4
e+Ed+Ab8VkqSSU1jAJr2XjgY+hcuTXJKC1d0NR2j0IpMnYl/KYHRIQaftn/8
4KWwDqvXdGsUdGrChIQSKEMFWywUQBBznNkNnLywlJTfoIE/14GeIVD4MJO7
iQHvkLAuIBt37mjZbUG+fX0tEORdHhezhM3xifeoMUHqAMRG0ZfjgMjuQznt
pjGss7SVuD7v1rP7lBixbMJk0woyLhwgbXdlOOJrOYF/vkO0Rq8pIEdfKgF7
SoRhTjTi2m8y9WtbgDMxtwha2SVa3i3XM66ble6K5R1olYYhr+NoNGj0WKJa
LfQgSOpqwp2YDn78tTfULDh3BlwArR6zxda3kbuRFDX+eNty7h+yxfhQZqz4
Egi12WTntJTAnLE5eDpBUjSmjHqGDVXA3AbM4uwbxHYlNzxfNIX1T5ZAgdl8
7v16R8d/MROv1qe5fRoulLW69qs5UGa6/JZj7Zbe8EuAB/jPfD2a2n40n/2A
EW1QvQIkptqIOp4rmCh7nAvQQPFYt/NIIqEzQ5Cg/D+l5OC7rq5whhumrZcJ
Dq8KKDMAd+AFPY78cEXVLOu98UmQcm+NeAO8ZEeNwCLNAl5i41NDrSzEujao
9GrNdOw4UqZS271jukV8bs+09y9Z26MVLCLq1bnaJMkv6Nmq8YZ70CJtzuCM
26j7HIRK11nte+npGqVbO5zfxlXnINpQ7QXPO/IGnyrvsvgEJnf//TQ09HI7
60GF+EPK6WKJ/OUJAt5y24IEE2abxIQ25mtCtJ1+dB0A1ed+vXfmG3WdYWMd
oWPm4nDYCkp7YK1hlEaA1ZkLBtLk9a34BgReEeFimtAd00p1fpRs57zBq2o7
GCdJqPhARkBKctjhPO87ZIboGJ2VcTHQx28dCtAZXyQM2JIgXZEBv5xp1o8F
XXEse+GVbp26uM7YUColfYRC5rVP4IZYEBlNa7d+Jh1W6a+dX/9pSW7mK5os
aChP6guPSOUnKYWypFmrnV17orlfiTT/p1q5pugFk12TZtB+XT7KA7Gl+SMB
nWS8Jjgc3NHgykeWGKkHS5KTWqqBA+XodT50MDjsZdM4UR7GnrROtXmungEi
iDTvhr//3OfMMbIUATCW7c8OaEGq5RscvJH7RnUR6jl6rsKuBA0Ryk8kjwNx
U46S5r2UDHd9Dg832eaadxhtQT6873Y1BqkeTGy1ftjAKv6JnqaZCkCFIWbG
ad5d2wA3i97mYBeJ26h9L96/bDOTnDSQJLjoVR2MVpT7yWyxuZ3MewkAqo/u
QsY6xvEKDNY61YhmU2IQ/HDK4Ft9LgcKFE2bsom070lEPfrZIq2i4QgNAwVA
xmdjpSpTINL86voQjMrbhV6S2Su38w6M7JfY3v6PFy8KB+lEbedK0LJVKyBy
deXItOnnTTja/tkwGLKkIYhd8/EhhlDpr4Hry9x2Y92ixY7eg1SlJTi6flyv
wRvWeSZFqgfOllpvC9W3RNcnRWpZu/buLTYnDxMZzmbjXndPcbgCkGHe3e6v
5syPouGOTR7izVepZxE8aDNYTyzTvYPDmeOsnQvv1DI3sCkcYhmoZ4Pf74+F
LBp4TQ8g2r4mPnGgslwQ7URxtsGMHlOnUoTeOiC2BBRhvq+oDIVAfbjlLtoA
Tyi8++ZKIJ/jYj+P2SykmOVRp7l+rSfUPct48bq3DwgaGSLkXBlcmGhXgTp0
ZzOe5ARtWFC44pBW9FWm23e8ykbmdD09d1tynk2mNzSbFG5vanAs0cYriUEJ
yjfyLwdhtMoqktBuhOS3CuiwldMIDSzlLR4bPIipxiHugcJGXw0SdPqWLou9
yDlcsj0MmXCpyERISh6QcX09n4t/op9N9O4+89SV9k/EO+zbgHheFTGCd0rk
Q6iUtd1YJnY/B0Agusfk4rb5JuKBEwG693Pu0muLE18AXQdNNXF0kCktDts2
+OT2H2IzyFMQPQKXrP8akhtJTRHR4a8eH98bT3y49poKAyXrk73AcIPiSpBv
+82SuaD/oiiQ1Woo+tLgjpHffm+PgFoEEdSGhsXupRBlaApo4mR9lAei8gin
PgCd9Zl7fjGrJJP33SURCG8b1RaT7Tf3TFdcd97QbIegLvH/4dsFfTyyXGXM
vYwa1vtJiqREB6z6KxMJrTH7wq8Qh6Y0ZFTb7KZOFQtD1fQy79FGWy5WD4up
79AhdlTGWZEYHyMGnix+N3nBoreD74a99mdLJShR9mDGKDxDk4zS82Elp6L/
gOVxxi7FrKbgkptirHZwcWeBCn5nTaANALD3xIAj+HQSdYFpiSSIJFX8N0VA
PkS9GIogV0qpg7eJTBzTJ9ctD49RrPGawi6R7BbFOoBfz4EL4I9Sy7t9KX2b
5Mqwsk6WAV9THCnm6VuGRm23lx9pPiYPWuLEc5RVhmUKMiTEiNFH/es2TUkM
yjGltcu2qGpIzxliOqqEPJ3BfZ7Ey/64vmO3JcZZJQwecrp8QGXT26HzzPBl
RsbJbwYWv+HbyTeGsdX1h+jPdrUtyl6cEB7yCbPHBgr6nHj8izEq1vgT7Oxh
/ITPw16Ughb65J4Lf5KbCrbsZIn4UlOnQG0f+Hv+UL9XoNXrACvNynldZZI5
nnoYVVmhOyI/QcHhwNWRFOX4S7/v32LoJpXYx7GkREGGAo2yTImCWgIzpE4K
zkFQdixMjFfrx/WsnlnKfqiKAnn6hs9pBdBhzNc9kHdQxEgjfIgFwIgx0Pmn
SewnSHzpJI8HtIGERNFokU54TpJXqcL/1sTob7C76ILoUUHDr2AFxIQnTuKz
U/v66f8Y4+FBOeU75lzg9j5/F217R3LCk7+/KL3p+tD6WIOV963mh1rnU4eE
ujUTxQiC4z/ERfKYa+K6z7ho3/DNzvQATpCUMmEBZcpc/D/xnSuopButKX8E
q/gE3XhgJJXkf3AcEKFx84Fgv8n91Q4T6Elmj/y4OTSiOiVOKTWxguWJsR17
7UCdL0HM8zvgk1KK6Zh9yioidW7ajn4hm93niIoPh9S+3hW+dv/VpZKbN5N1
p9z+hZys23FMNC8ehIQOc8DYsXiz36MStsKn3o3wvffpWU28gC2KAOBmxykn
o26k2I2fHBQ56O4DnvqwZhuZ2iUzxLgithbRmG0gfp2Xo+17/FomgzJJEAlv
xNFtdOB8D7yaJAFp35vMYLU/zVQTVeYAPINx5OLVMFQEmTOvc40NOWFt8+fL
lVwAqYZe97siplzLcBAcKXfeV5EYQHs/fSvaMSq50hb1+afrfGO8nF73y8F6
SbKwRUh2GR1ULbWYcnevPA+fcW2mzFwMajH9+rajRtv2lijcpNdd0IcOErpP
xi9HEnWdZoHPCcs1ePls0tKd9iJ4Aq5HDiy9MkihVvDpjuXFkdW+d7jgXkj+
zK0J+4tcFH1YuMmoDLFY+5UNRZ4tsY6QC48xGCnMbYWlHOxu9KCkh4PHtZP6
gdU7Opp+J1Sb5+PYw4yh4zrBhU9XUGYmHHyyzA03f++vhlkRU02EfYd4DQAM
RFE2utRJi1QNPjPlr8SQ0OP2Spm1IBsJGBwnWd43+IhEw3vAgsx2bABw1k7S
vY2rYHGeJwAqDgOyIFlGooUCTRopTJa/KC5fbH0e85zL+gMHeDsCF/eRFQOo
ZiwnASQ6b4nNBhMBDnf9qgejiKbYonSSBdWme+jv160H3t5RyQC1BCn34YiL
sI0C3iWOALEJo3uwSojSjMRqqINPweb4TJnJWA1uW6frAg1K5lgaDP5ESEIy
3m/lmtjE3mJmwccPkUyxyxdxjQ1N/Uw1pCHwo4XnktPHlW0p3KhklhvD0abk
jX3Jm1UGoZfKvJEkaSNUds9XdNP/4C+bg62bdwlXMYwEd12NhUyz25+W38E6
ykciyqMWTDq+hj3Uw+4Ca3nnfi3otC263Ouuul5Z2awXn2CclWGf9p5PvhZs
7Un57BOXFrQnaJRgPoY9O+KHstaeJZR6Mg3on3T7YftED8+hDiBuT/rKvjfT
vR7uAKPZbgSAGB89h2BiE8XTyJVbM3EfJxVk6Cop8LXoIG3o78XpNbI3kofQ
YNrl0QsKSLmwWhJnK4uwRR17lJQ3NfC6WnOYpkMAGytYiYDnyy558mhTYYWa
kq/fnFhRGaulBP/aF71iff94DwwbKWtfspFZULCZkV7CTeoymwPn+b8gRJAR
aTIpEE7bbEvp4IdwIUMV6yo54kzKMHYZiKVlBZQboHiqsk41kna06L3oLeXE
VkMc0PsDyyeXf1jl4SiGSkI+ReNbMX/yoN37NkyqldgX5YR0f7v/nAYsV/0d
jxEIAxIZBfvNm26yjhnMfpfmLrf1BgTKe+5UFVuoEdQplGAOkytvh6Wt35/n
d36GzCdSbnuXwhRvnNg3Dk49nXPlMsBLp538i/8Dt3YEsPGpG/U+PyUYMtwT
26JAc2mnKJCvOIMruqJjyFABMfb6C/LxX3/LT5+tziLdaClQCdvoQ5WbuSlL
wJMEtbSDcs8Rt/iFFCKm4SWp9xYsTIag1LCCXB1INhd4++MAg1QhkzZvMvEF
u/+bREMFx2Brcni2w4/vLVvYXugtQh5YEZB7YnE2HAmHQHkL2hbagc1f35oj
xwpoG/2bpPX4BTnmJp1sUo+MyzHePX861h91lwGTj/5KePiwm3FVCUAfNWZw
pZzDPaobAiQM628sK5y51NHHQ3xA5xoOO79C5keycCMReFXjcq9Ux83ro8LM
5qLuvJz+zB5K5AQEJg82FVgXohFSNkyy/LnaW93Y8U9dg9SLpn26Wi4bVbI3
oOGqeY/7tKEuD6XJDy9KJJ7CAQgdjPw7EcqlPOkU8pIU0RxLnyve4mAmCDHW
F27ysly0sAIAOMI0CO7N/+nn+PdFuUC0RZm8tqHh/bVClBUHnsdGzcHOvvMV
lVNOIQIM7yIzmIjFF0dTSgn5muRUrNuCjnCDyG5TiiwnF9bxGqK+JqpC7Bry
auHZFRLhKLvHqWCt+R3/joc1o4uOeHpzCvBCKmaA9yybSgdqxxl/vUQDGEX/
xGT4iCni1Me1R4TdmncMw2Z9oGxYUdJ0re1vRUtftrENZ7xbRrpJ+c2bfCkf
jVlJHZhrkndnUvOKn/VA20LqnNCgWsauqFAuGKGWA0ci0HHbEuDHQP6+InE9
b1k3igtEmCNXyUUVkQZ0xt7QdBKgGmXsCcknu3QQpM76H1Qmgj6AlU3ONRC5
RN4Iwgt3zNwWlFIk3v2XU6wusjQyTAnfJyrryYiqwfneRdkrKfuhrBGNNNvo
jXJj3mTfj9M0IVLnWI4ABYt0We0hFk90vuF5GhD2z45MuTpKLyINcyIvJGhV
HxkDdmJlOFzO4TTD70bB1gYKy28HLqKyNkzSDx3fxU3/tgAQep0E0/uz1jYO
isNJG6pMrXdcvdMD+fR9kabbBuhQC4CqYyrKTeNBDyVP1WHbE8GbiwY+pGgc
I9WG6UByYDf79ju70/jgE4Oj7cWNFVTvd3LEt3/LkXNIv8/pZeayaUlTSETS
2b5JmwRBJL/H1otB6DS74eQpis2wJjniow/ly2/bKz1mFoI+nQ/KBSPi52jF
P0jUzKfuF4sfFHB5zAMHLSfH4RjYy2t+UVVZZNb01W/eODmHfRt1XUNk7aGW
V5fv5MyLyl7FBm7wg+slEwrJuMH0wivCZj9OjvIUpPlYDoKdkcnvnLKpPhSJ
h3dUG6mFrwkrKw2ZS2tumyTe/43GcaE5rZNzUbyZhom/IdoFQqDaGq1z6wJb
v7ZA1odcXq8syw/DOPCLwX3pUewqkqKJ0kNnHHaWlN/U9eyeLvYPSHnu1EuF
mJ8OtfnZKwhJYOPnI5Cwt3tASY010C2kUZKNNrhsl7yeQ02cY+ZRwOkFv0mg
2M8VBvq6S2nmFHhnbHa4zgr1E0SKWm/uUWfPFqCQnKd7PQ+gfoUDi1FEVLni
i8SZDinUCn5wOMNNn+myBzVIK6OUTFvG+s86h1uCFzwx15RYsxhTAUF/H9Qv
ZFiIvc8MbkYUtdv+ZGWgUYQDWhvXsylc5qiEJOcTBa12wSaSc4ncv7sgWZwz
PNu8+C5yA0Qf7ke8WOETml16ZMUuI2ZsXZjmjRGlSz4VOtGnku95dbGDGuM5
q0LAoBKAFoPOLWUjd4fG9qtU4b0vnidv85JVf9KEDRBdyIkyfs1Q5ZJsa5q3
b6CXkh83Qx3OiaLHm79K81HQsj5zKh2Go5FqzkgQkw35ZI38UfcEQh+FJx6b
Ya0fr4nHXLGnJYQaXKhXGzP8s0otiePB6Ew08EyFhljBc8838LnVXsfwLWaJ
PEM5c9u+VEp23Lc8t8wkCqgZ7WKsNk6gGA5X+AktiftZKfD9TyY6RRHE3fym
1NpXtti6dnYn/fpptURMospwR8eCfdSBba8Qv1l3h1l6N6bwuhNiigAyJqjy
+siUnaZ/Lu12xLmnbugswg8IjA0iLvCmvpT0ySxfONH/VhleF11nsYNWa0NO
1GivE8wxnQaRD8uHPhV05FFczR2HDK8YwaijjQU1x8P5arOF36Dr5Iybgjmo
glTDUZmxHYd/F+FppjHYul1HXlkqF0qBifaGssDwyaVUdmY/Yw1F5/WzxY+e
8avtNl1GU4rumKK3mkOa38oe1ZV7xWK8Jq50ACODKxj65c+7KMaOvvjcqhx2
oC6BK21sDJdFsyNuERWB5/BfdeHV5rPMgSjl/Rr9vfXRyMxTVfuOtcpnY3oo
z6qz4eDk3QZLObgCg3aXp19Iiq+gFMDL/ImCipv9atVRH2df/VYjhRLLRASk
jPxlTopbY7YDEXpEUtvAn+dKCzGKz7l2N5mAnUFdiqJrNcMwh32d1L1Fxkcp
8mHVsHmEKEc61kUOBUXr+Wl0lfsXqVEMBTu9mr9uzK2vcAcv1KG/12Op3TSC
Lhh36YASbgGDJPkiHCjBDgWx6z8pI8TF1fxue+gY05CIytEm9MT3DxylwVF+
/s43EQhWGSxnHjzzCWM1YGP1Ih+GyHwo8qMrHViJZ/8Dz8Zqr4ajbYtNklYx
2tHGSyXeRUcEsY8I9+PYuTtDowjNMtrz2B8e9JqceyXg7K2DHtQvcl9aHn6P
PEXJoaAVDmfzRlRiUl5+uzw1sR3qEPgfWQmzeq2bPUHjmH3ONZLfWcqGXfYj
UkhoiW1YQN+8IG1TpcPluwclFoQvimfQTlPW77W1u/IJll7Oeole4wGZwxAR
oESC5GhKgwKSyLBL6dslIF84Nk4gBSlD0qeoZCFYq73l/eF7Y9E3TEhsy24T
cylRSphSy35x02tOYDVapIZ1wg2mhM8xfjVaKBBRT0mp4Jj7xJnj94SzxUAe
STz6+eT57qtcphWtgBz8F/BBpapZmkH5tNpJrdf2ioKY1Z3dNfb7Ajhq2VK1
QeDslNh4wiSpfasgYP2p3uqtx76SGGPCh5a61G0mha377zhgJLsxXHau6+YB
1v4wGbrHY3LFb49hpER0l+2kPkZ8XzHTexN8E12oWD1CiU5OR3OUhE6V8bWz
mmw73Bu2U7fMK2VtAoiUTSmuAsUFiFHsPAKRo4cnfGXqP+f2p3h0GCu6t426
a5qPDlVra2UCIdUJHb48GlN8tYqW6Xfq0Qoh4j4qefYyWrQjHrnhsWduew7Q
FOfJP4crU/FLSxlBWAHt+trqBqOLsPekKURUof7m/oDnTX+yQUS3h0J7Xij6
W5vijKM80o/Hidwvi8Asd+wDgaB3+NvC/llgFHe9XEhEOGRcY5+LWzIIoSrg
RVMFbVZ6qh8Lpfx/eKDDt8qasYdhhE8ICbYzeXiv9MRCUKfVAl9WK7Vl/qtO
+NiJuZUIB156P4mDycDvIH6ic/08LcZA7yWlH6xpDChyjTLp7t2EbVoV9rZo
vcQC/39+Tm5OxPGloUD8Eie+MUknp5rwVJgIaaMNXsRskd6ZTjMXTbtB57KV
AfwrFgmAs+XspuDVT+sdOAVVFw7vXtIREGlbLbOjlrb0SFyLoViBjpVU76ea
SqHkadikhVp+5PhhUGI8jtvh9/G32CrJvqR/Mxc6tFdLA17t5AEZtPtZUetf
trpz4j8oErCQyb9uyo2Wjuk8M0/U+L+XwgjzlO7L85i3m49wwsU5qUoqDGpF
0DPz/v80PYwcALYsxSfG8v0tjx0nir2USDM4+GExw4cZPs9YxyI8ebgQKHe5
ILh1VPNq5Qg6qilqf3RpsU2FHkNX5TAwC8hruzn2USt6CtiS5MvQDkYs6m1c
B12LUDMbVUVSNn6bnlRhccUsWccnPD3L+0H4Yk4LIohyXgR6GjPu6cU79sdT
sCvrtu6a01S89Nh6lBI59U1oyB65jSkeqryGcNH9E7PYRovG1NzzF0lwm79Y
FW6P1e3Q/lnWs5VyT43mGrj+DA9u7omLAspqQ0tyibiVZoE1Yq4zaJKqRcgY
zzYUI8+zbPXHRGtoEF5Zgugi6SLFmpFqccrH02x0PD1YrbYWDk2Ueuj1LxW5
lC8ltTcFoYkeEthRJVUx44ggni39ubu7ize5UUdbbNXSJHvmFjWdZifqAmH6
A+4L7iu7fEP3A9zrsDrLUjd2UCZB7rZbEAtC8RSBbhe7VK2Lva/n++TLgHuX
3BxIn4rVZNirHGiLaH5WToI3b8PQSaqaeAnr6O0ZSgeyPadgrn9JsHpLvbhS
ZsGgXKDq4qmOKbaGQBcjpV4+WhtlB09MtlRae+KqzFvIjxzU2W9pQYQdErZM
WdZ0QBgJom1/QxpBWeyc8M+zEhNpJpUz57ZLKW+5WnvUmjH+w/KHku8Tqwyl
PDBOOlqIVS+TCivJmo3gEGLeOy4TUzfg9KDC/8Ri+XSkAy5y4GlNpNheVGuZ
HgAhkbp+2dGageHmBiSg2GBnZDSdNnJJDp6urJvFCTP3w9b0oX3NqCHXfUZR
xFhllfVarNCw5g1JxQeX8DmfNBwDRgXTI7FrBoTrhJRsDt1zg9shzKdXnUy8
vDkJYQNdo4Ax8P+ObbmKlM4Yzr6vzjm0CGZpNlXC6qGyTFSccjYawcvNuelR
07GFg5HxYwz/yjIHF8qneq0VqsRCULW8PZ4vony9SX0rUKGKrdx18ZIjpSip
0jlHqBBsnS1PQNZC1hlWFMeEKlhsT/Qtdw1SZ6O9W7P9shoAQBHV1yioKQOh
HZOih9nF2Tu+KLjLLNO7Uv++vPfVM7K8yJJ0Mcrh2gxyESBXRMjKrJFhTB/Z
Uzx/gF50CDs5kq1j2Q8xc+IWLqoCn3+qZWgcgnOCXpUPadsRRwJoIkVupCR4
dPL30DdUyvwYQvuVmsuAA72PSDv05x+ypJO1H3VzWPlD8tTyCALtmdzqFLSF
xZsVjyoUXQKa6s3K1ajuZcvGihDyag8ba4y7mcyo9UYwpyWLJ7EvpV7NoJkC
lEVeB7Uas0Y742Qb7vjTRilZfdghpPMsIuB3CyztNUtbhuv+3dTqXcGmRJZr
7zQkIeL8yz7DqWDKeQl+J9iKxMWs/ysI04p/B07ID2Cc89FU1bCth2k+luns
SIJ9Z8HNgWvBM4ayRmpNnCA4eSjQYwZ/mVxkTD8R5mglYCf5IQfoE+6wkH7I
JnIPVstfyWFVmsfzbPrWLw+HuS+WG1QxfEt9orFWmEiV4LeHQAf8107MDSUr
iR6QIf1wFKsLz+gA/sggvn7UEm88hi39v8lTnBSiiIO3ix2dRwC7l8iwwNp4
uc+hZNADpLPS21jmzxswomZA1cVNAKq4eR5w40+LvmV9bfN+0zULcKs5hVMv
96ZEYEbeHQuV9pwcv0lnQoNNEspZNngtRJmRXeTf59k/Lb/5d9qrP+q7kiX8
R5xf0ip8ByB4sQTM/Bb5BngSPdaXhlBW9mBXutdo8QTS8jh/kSRN7U1lWD3Q
D8WpjaXOApoCo3XBYBKV/V6xMunTlDVtlZtqeuBfd6QW88NGHzjC96NDjZ+g
0MFYSZ0blpYISMWhWeuP6+n81/pXvW8DlEcnW2fWko/MX70TUyiGwoGi0Uma
rViPxFJayLzF8bUg9iXumlyrKuoO1hdAUxLr63PkKzG0Xy4sal5UhjV9Ulb8
xGTZqcqiYWfsivOQHw6SLtEG7hzRHMyx1g/6alq1OUby1Z3ffJVa3XX0ATll
RYqxxSLZIWkWtge2W6zILkqtCUS3DBIiXpnJdumxL+Gk/sJPl59g8IAUN2eB
49V76J8+M72PI6CRU8sSVrux7lj7JzUuzYrhaiPT8Tw7JzxiYiSwz46/zMVz
aYd8hzgBvgQG9RRB8aRGYMHSAwzB0Iem7xoF/pyJseDXtSQV7NqjXISQnKg4
pyDhHzdVzJZ7F2VHL0/Wex+NP3kH1SuDViKLhF6Pz9a4FuQKRNjMz1b6tW4+
2NOzF7djU4boF46m+hQHy1MNOiwWX3HBzNXyBYIepCu/Z2sYaJbcyZkgqUY2
qDplTLG/xXaSmac8hfAaYhJjMcHb2hPFFQ6SKlfKHNXOEC2ro8hJp3QY4Z7R
PM2y5wtWwOp/MXeWHbtBpyyOwlxxduYRt/AQrTzKsHjh56vUdYW9CmYC5jRb
s4jLd6/HlJXk4DyihgYewSMj9To3vj6wfGvZs3kfe7b7BE8aOrYbdWeyAu65
2JMoSKbMqWA+2akM/PZY03g2WYdxw57LLLJen3akZaPLEBk+x5C5TK8XrpzV
BtuRteMAZ2dz0uN2Wenw5ZItrpZbnalQITmfQ5q/hyMEglfd6yeEOXPLtL12
RjTDRBCTvdW+NuH8eWjATnZKuFIE6ywiy5SI0/kQVab+WE3DpusKVB25wi5X
sfmOPh/xFpkrvYJNvw8xNsocneZALmwHG/Unk1T8dxvpMcNTAqEF5lJaVW3Y
MJ8XC1Cff1P/hLUZX4VPcorQ6oIQBeXORGZJgAbgtygd1eXhN6d4G2daAjWU
BDYBagiQWyeCoMLvAmb3qDh+MUVQEtNS8yEmKDGBC/qERxEuRqy84ioFDDj8
/c0WaYn1oenF8lnWT+s2zO3mmfFmAP2uDQJ+8Bb+vvz2BKpBXWfeGYFtnSu4
2fBCtdFX8+RYKCVLPoXDFQhBLLhtnIvkw6TCiTwoPAGNx0Q2LyKzM/DgZCns
P4jTYUDjexyEcxk7cL3p8RBmlmIQV5u7Pj4CmzjN5xDJPDJYuTTt4Nv4BVoS
StMeO8S0Wznzrefmo1K0+S5TwvXiBQcXMI3MofHoxwZSL9KR6WwIocRmxb98
t6L33kpVAI068dvNoznFWTyvEDzV5UM7utZJFSDN409uvbJ7pT3K7+K71yKC
YcC539145arbHPdJjzE9TRcJxtYOLZ/m2p4pZ33JzCh0KokHGbHZaRy2uIPr
rxu2K+F6FC63fBxve8cT/dOhJhn6OLdhkNJxF1d3w4+TXw8GA8I8VkiLdO8d
fvTdznAfzCcpkoe5i/6asDM+lewbCr8oFRi21Nr2+9oDQMeRH1JfiEkbIpz3
69cQrKlvJuwnu+FdKbzj8FEULn9kKP4cDziajcwD3mcZC3STEwqHoatSgJl0
c+4QdLn3U28U71lFwt1556WiLnvklHBnw1miNN7IBFgcWT1qM2F3A7kIVCKg
nIwLI1+owUy6TKgHBFzMlbZMzdlk6sySaGmgxYuVzl8Y/UZIr6aUVn2SQd9l
ozK7aMZ9/S6abYndbxAjWMZBvLKtrGCg+R3kp7cRKb4HOMK2WKCKYSG0tp1k
EGzTQhkJ/T40Sd7cTrVh52aI0tYn5d1IiHDDO51PkQHnq5Dg022V8mhbX8ty
GERYkBFbDFTx4a7FpD5QsxQnF7EqbmYuKVDGQ7dY3/2zGP2wOhNIQHNVJx00
odfhb89A430pz6jYGFDTEIXO2I7u1ngCFsEOLE6ZJBQFt0Xa3p7lt3qxEg40
DNBnYOg74LgYkeCZJyuK+ZGr7gt3+wB3JHob8o+MRUrebNEEo85GkzSIAusI
ZznBA9zIHjwrZYgETi9mPGxdecUdrCNFcYzDPwCsDCIjm5qGHNb5oNjpqYbM
PJe+QYNnOUR8ZwsP7f8MHBx+2kZrTDe1mjJ8Nq4PvZ+VsbLz+9U7Pra73z2g
3uhSdWvAo81K7x0IZ1I2MGiWeGd1V2FWctU897YXrbopwB6RBxg1Uu+eyPxs
7VLnvyNmRH3p0H8Jwbv9PDuPL5ZdOWDi9yltR7c5TH8pI9v+zSQq7Rb9ajs1
hHSL/oU6DEJfopglUQRcdpoz9K6DR1BNkqXf5hF5oSXAMlpLcFGnuZEzbxr/
kVlDsjz1kbCuzCMYIYRvnxH2+uoqMM+t0uVvBuDnhI+tu0iTzipsy7g9Tmxj
LhuWSpIe61QEjqygEJmuN/WvkFkB8v+gTS8eHMe36nw+CRbAI6CbejRO985q
yLGp936wYgGXQq3TL8apJDOy6AgoF2p1h9mReR3gXTq+5eFdi1YEqZpBVK/A
otl/+imyUONkxjkxzIpOxfLOLf4g03CUvLHs7x1CwENiz2PKyoY9qQZL1x1V
vMFTkyDDeFfjf8/JTEkSbbJbamkDXzqbqBQewxK/benhKmqO7TJ3Vpvbt1wS
GEyUuNNo8kEFo19EUTKG7E95qal3q+7PVEVSM8QZ6Cp9HcEqxcLtucMxQ7Iu
obNe2cugsmh3SAiBxLoLqWw90DBGrOr6p8fee7KmDsmVNav+zNWHlNDFsCyG
VZdimRhGeKAbV0/1m7+WRo10udYIQuB57Hrzo4PuKVv3r3y1PXVRspmwfnAE
F+NEgeO5Zk9AfETRAhW4PwhqBpCsAqw57nIRn8iM0mr4bnF9DpWJxND8FqzD
W171u3JdzB3s37HU8pvgEXx1DZ2szBvaD9hX0asJ5z0LjkGqmlPhQMYEn/y2
NIq7F6vHx7SE8l5bsmJbGMuMZ2uT86GrwX5szPH6BPItIa8oSzpOWNDJa1qP
nTavSuuOOV/SF2v5aOUTg44Y149uA3k8bo6O/QHsuRllCID/j/8uv2NB5tTk
jelAKCKtIAU7cF0liFIxNpvXd3rRIuqVG0hRjxty3lf1cOdiXh/oJmnZ32A2
KHMKZb5LcwcK9wfcvyROYFvXWRqI2Wuz2IkZBlqkSYeevY/h1a1BLeXMHkw7
7kB/Hk9siRldq6EI+Jpdh+khCC+6abkgVacRoZIfm8HQBIbjrIG9zSGllxpW
bsJi6/GgjUbiLBJhyeEUlWOOLwMG17/7VKQ2d+paM+7yz9yMiJhvuSsW199S
vRCAmcifmlZv5irZfQ3yoxQ0R3mDi9BsEug9HZff8jVurB+F1ygncEGEYOjV
x6ab5soRBZq22ZO6UTjAnSLJ1AjAnwVy7Q40qmeuFmIlQspu100yfEKyk8jY
/7wPMS5kbYkWHijsdqpyR+R4apu7uwpEVuRJ3yxPXYKiJh4ef8ZoBOcLwwpJ
2yHPP/bDVBsyOFHBOTgxTG1VH4RGCbVMrECE7TGYV2H6p/JeA87iBScvQk6W
VPomKNPnHr6UgUGEpHOSk3ubBF81j7XHk/XWcc3I7/fMd9Bj0ox19LanGUfG
06aGEJDtiL6DDWHmrUl1IrXGMeqiLV7qgjgZujxX7JNfl4014RSTAtkp4Nyc
PxFnSOzTUWeh4KMUNmIj2Jj8DZOWVaSgnnc+fQinhh/E1CquQL4yqtfh4QX1
TFxdZ5moG4vQTZ0GQ27a3GvzdqIe0c0pf/wJqR+ND2ZSVlisHkO/JnbBdY6m
eoIZG/nCU2Lof/alZEFgIriDovkNxnF1gY60DWTpZVgg7vlvEFTUYLLVhFpv
YDwZXuqYgz/oYdKiXemBaqwKcaf2O6PhzU/KuM80M0j/RnrWVWhouFa9Qvxm
eYYr1/v2+bxWVQO27vg0r5H3cV4VaQubJPnWnk8moCEZNHvoGfNsUVcsbdUV
hAm6ZRU59mouYRVtb0/ezM92oUm4GMEKBAx5T1IT47pNJMvM3qyYLZlmKJan
k04CYE920OBYutBWQoKF0SYn61v3LxktB+W8RkNq7rSGEtGz8qpUUQxho+cA
84bNieMUIVhYCXLJP0gHz5Nd/yxv7pfW2J9gpDfiBpTKlj1+DL1IGAfSCaH1
7tOPAdP+BWuCCkgElZlCB6JJ7nigorwq2uqzfUJyOetMJ6ff/nb2oLv0GBTR
/lhQ7dU1bp6AFA88+OQ5rXm/URxAo8/jMBjHlUPkysRBIQFOdBS9GcSDPDn/
Nd4gwe3ZAPbSmI4mloZPJPM0glouKHHLYbvZ8L6FMGZ0dqBxEZgqJdgWLetZ
H5x5z+MKNLFLIvvkFfU1q0CMyfkG3j1XcabaH608awujKAh8VRz5cVe1rMqV
KJSXqe3Tzdqi2z0Q1eSuN6ENn7C38Yyzhkqnaowf6CjcVMUBC+bcUUd+6iRt
NflN+Z+hOKa54jlGB37DYuTatrqLk0aYNsf1aM4OowKl6Fvb/qM0+KdFE8CE
T598kN/PgcR+Pblqf9fi0D4qKUqtJa0vQ1QO+cKOhfx2gI7q3+jLSk2h+ILF
h00QQvL70h/wEOQF9daESxdALm0YcwrPo42crj3K4pbYhca+PasS2xZ7dJE7
tIdYve6gbhFm+nQEkZIDv+SgaoeOJDlXzuRv8vSCr5CwI2moT0YZ535M+U3z
qc176wI8RkawrK9BLtb9WuawhxJFW9k/wYFN6KUL3N6jAPqNYMD9yBAcZiit
x3Rut1H6OdCi0n6ZY25wRKfeezWbTYtGBFgu5TcWjFX+wMR+1Kes+JOKd/gR
0889tz5PloCA4p6DkbI608j7Tu0YjJXzlzT7s5eaGyC3mo0eoo1PTZ3PgMix
8aAEcFNK6ou4sD4m1B5QPjqqlHro+6ahQ0XXox2DQcxxUGmwiskUhyM56Sxr
Xg60/tZZXthVlDCzcaT7pGBhGNMIUM9XkM55D0b0uB9I+CpRpRRo2XMc+WO9
HLPhg5KevyMJ/RVuk66yzBGvXDmbyQ8NtcJh3owReXuD11a8pqqGU940Zi6x
to92Wu3wlYA7uMsN3lqfmXNgYPPdP491swNINklWCv8nudNNAOQ3UZxHJkv6
5VtNQkwRt1yQ2sjXcybrP+3JjMi9zdx5C4cStaxf8hX8KXl+4JDE3ByiCfxL
o7hDQxvQWeNsDa4UOU7TYSkZ/jS8m2eim/M14s6ms6SpPhRK4mBaGO7r9HkQ
kDjfWy2iiQ6HkydU3vXMhYrLwfP8p/ZmKLRUbjhOih0ybTWi7RwG3rO3Cu+R
XxfHSWMBTb524ajxFpz8XV8+VUtZe24BMYeKZlUM9bx46rCFvofabgD5d9/u
4eGcXq2jhWsCj7uaY4vrM8EoJ2TKlpWUHWweZCGgIxRATJoL3svV1//J0NDB
ELp70U8qOmvruzWINAphHyNGh+NXtqJlQs8QsD2p/yZt+Uvhew6FNDw3cdlf
hwOm4bgqhJFsROLxuOicC2BM4u5eTxeKxOhlqRluidhs6+ftWwE5OT3OyLLf
bBcwVFicXSrQ0D6/vYgh1G4UCqtF4Ueu0wl7vkR2+zVQpsxrmwQ+BOoGFZ6b
WeddLjL0msxPWUgiSy6FmQyeZbkb6l1ywadT+nPxCHv1fF+j+a28VpAiQ63G
yVZiW7EqLKIn2/Hjm1volkSO080y5GG88JUl89PH1N8oB0MoNNykcIaDjlEX
oc4vRx22cb1I6luq0E5RdsSsKvjd+ANuoP64xfeCyYQan4tHMIaMSRcQ26OL
QvjTqB2dzvp8LZaVEsJLEMMTNlIWFEkaLTETKKLA9aCoeSXFRgm30hGqfP6T
amuEHqUsfdHKDVyvNmAyUbfLQazSUVGqZ9mNKR/2Ni60wOZPd3ECUaPN87pN
DP4eXQeU0PfnmtGX4ZPAQvAnBfaRa1psQEC3ZGxbZepmCn3yCeQidvSB1EnU
Ra/YLVatRdc+GEsJvutjwHI8ySdJFxIh4lmSbLQULckssKm0gCBFPZBI8YrZ
Jfdp8II70TSLCm3mze0fD7gG7TFwa6xSo4Pl7dH/xhHewhXY4BwHpSxQ/jnS
vBEKHIPnYGxU0QVE+zVzESiZf1ETxFhAr6QYX7pUupSu+dvDOOLgRKYY6txS
WJ/6dwhJrYqrrPXUtF6S1fnnO5VkknbrUIoStCuGgRVZ9PIP/VbL59uDi5qx
jU0BJJQuCQVnLTinSlp0Uy/HmwVZ7Dapowcjm3kn21Lv7aH1Je/AkCGBl1tY
l6FpVkRlJGic9mF60/cNNo7Fi7gCZkpJ913NuKKXTWupZFEkw5oQU/r7kLo5
x1a3oBErlqLp179Nk/fXnrKQczV3BagB/D4SHbySwZaRE3A2JEFwDtohulBa
3PSDbGQKT8O/kxMgjt42a3pQclu0VIXNqMFO4nCj3bEXrqVJk1bX1/lsUvCR
8ir2yPd8FxOcGydRoPAl4OycHO3TinmFGJdAvN+I7e3P/du00X5Oa3Jdnutx
qOGis5KTqZo/mAWOTUjIAVGY06roX/rbR6H/9rzOl6iSj6O0Zfy4Cq2ZrXxp
Ro3e0WR1g3vN8q/aM5AO4KDiqFRWVCeqCxnCdzcuWQgiAyvrT4QfreeNHHLx
J9sW2eo9LcJx7kyHv80CS4FsAo74/GtcEVX8RK11JYopt0Gi7zbpKi3IP72F
bBw4JyEDMd8M1NAAQfXqSv3D/W08ZPRPO7InwM2PDHdtWXsOLNnDKRxyJeA4
pG/HXhMpW2XGxSckfA9AqzeMolhy/eZPudm+Arebzl5vlGsKkc2G0mCHLbwW
I6RMf4ySMDx1mLZ0AMBs/fTRBFZKzfstSQR+LEPSozqb6H2J/jZY7URdUQzN
2BqaB73mwi/4delsqc9QJc9witanxZ5YXWznn0xE2ZH0Onkj96KiUDz6gOdd
+1F4V0v8lIYB3YySZuq8Jus1AtW1BP2hTjsnwrwwsP8GdTxDCrvrN6kjjjLC
YzMZWyV6GqC/w8D95ZZl0VObJIe380KddLuMB97R9axuDW2HXcA0gAMxSMmk
PP45iBsFqO8hqyhDCqgzuBmHGblBbhoUYESzTRX7aGIPHh9qea2M7y6o+tqA
QTgDRRDrShXqHijXdkJ/u9zNj/tFAAUC7g/x9NNDtkWqB4ysH8rb1ghOQUov
F8LMQZTxB4cgU86OPrLLyWD9TdlxnTVGuNmkf1jA72r9i9GwOAJLX037y0yw
XE70vecc4vRxvxBniNRpnjZ6fRO/NMWrtXVhLFBqN+tcBx5UbGCxSmEs60F0
pK6Pxj3TGCaP8qwELnXMcwhhogECN3nmsc/mJYHWF6X1UBGAfBxpqsDwRLca
dkrzcnecGTdjAWamoyyoLNTsEAdbQwN3lJ3m5A8Ec/ziWWhouDoJw2vPwKdt
jq4rj8/4h+GoCBtAGZ3sCvWFAsqAcK6wplz+GKx+wFhqHnKFntNk3ggKN8Qv
hYYXtbTKsBv6B+yCmgSwnNJCOKa28A5NZYUVLkzEsKnmdrbjJ5x0laA9kR8i
3Syl30mKKMNVKZw4jneVp2ntumo4IXoRxfDWW4X+Lpl9NZvDZVxarzW7YZIR
pkoZIvNiNGWdbGyhVsb6JCzqre3e3Jd4HbU7tOtsNsfEnGwPCF6lLPYNKPkc
T84nyjVqVicuDRzH4WTmBxE9+Y+SbpbPC5dkgss7jIsIXS8blk4xNR0Av/t4
q/x84wqYS1XYU44PNix+j288B4p624OBZrOCM22iQnzTen75V4B6bc2YxnsO
2QQGmTg7O/89lC5YSnk5V5lGVzJZyVar/+kkpPGBgDhtDI78Yf1VhvrydDQi
VyrnYhHbZjbhZlBjurGwE0+4G+1GgSAp3Gfj/OMfgq6eVOOQSwR8L1AvOjv8
+jyRylBWqqVkpFBQL7lTKP0kkHwJDXNI3mz+VlVL9jexjHi6M6ExkGGE/EcJ
CJ7NN51IzrsemjK1tRQ4ipgbyCmNQ7uL+CxoegDW3SUOA6GsHW127SMKAh5s
9Lekyuq5smb9czZ6uEf+RopimZHb28S304yW9jlZJ2n6nzDLsHbumIGb1qWh
ErMbQoqVDGiqDzbHtwEBLYFyQ49vOkpJA4/Ev0t2SZwKeDVHXAi3yJ5PteR1
+KuCeOr37FDiypaLN71m8vxrnKZvJ1PsSChdOSDfhdsXJLQGY6kttTcELIhl
XPxo0YOIr9zamWVm/11oUZ35h4p7C0rrCxpd6lAHypowgYnpHBX/hmW2MZC/
PqPCYcY0G1WB2Y+O4BnxV1Atv8KDz/tR7nf7Bmqja+Wyqzx9VyqMgLWV5PMw
IC1FWkjcOoKYI4sVBVc7DmJ2oBzLiiRAVGs0ZkzHjdFzeM864EkLNwYrTMRj
R0fSaa4zXDLYtk+hru3rHCkta9jbf860vy7gHDY7CYcgvH1IvVbt+pjruncU
nr6PRskjWpx5dH3lofLiinS64J8YEk0ngZtpMS9Qg/s+BVO8oUf6TSZyIQl2
fzUt1LHB3mn+AQdyywL8Nh73cgt+oCIizraV5Gj46JIghmXAorKcpDC0XQrI
HkdZYajabNYs+wF50LCfxy+8dgCAWHR7b15T5iNO/yQ+2OdNj2aB7/Cyb3Uz
rpC7uix0goL+nI9ExsZg9Yb/u/vpfA628SEaWRAnpR6Uc1rQNH4Pi4virB+8
UAMUdkJaFVsOENhsLTGm3iAY6xZEIa4AhUdqoTnxhu9kFnrz2eahbyyp1c/g
oskYpVsZY0e5BDON/EwMIRyjBwPvsfPQkz7XfHSQSGsXqVDQhS0EXlc1fhbL
Dpxg0utSowT+GjttI0un+ePFACJmG507iv5rmvlzto4SzCEJU593GIS+1Feu
LtodC9VDl5KwPv2ow9ON0Qz0NELe13duJcFAEhJ9eGDd0zuCmzBey05QqA1f
oRLX/xKLj743Qo5lL+PsWFAS1PhkWYc8Gx7mD1+UtVBtbUe5wYfBaT0J8p39
hWM+bYiYrys6PlbiEeoo0eW99exwJ0phZHh18QDXVKsRr6Z1fcQAExntQaO/
cIgYa5jjfv+MlFKKSbp+gesOVQahnbP97MnBWCPtMj66QMt8i3laxTpiuFRz
PUGZxWtybZ1DVJB5krxZ1/JFyLxL+s3zg5bsqC6K1MbAixasnAcW7ZuplpOd
IwRk3waLATdX7a7WkP4TQRtyAiHPckNpLfYhuEdXyHK7cbdY4QY9ngKkyGPt
K//Tplw2s5BblSHud64U8/wIr3V34WFGiyn1qDT1i3xwi/WJC+1Eo4teT4FA
dPcGQ4GhY9W2GF9wn56DRDpTBCo9zuwuIjfH41zaNlyq02ZV0JJgHj4vgFIH
9gY74ZU+LzNv3STkwD8UZF2hgnN1BZGtZ5uqy8swM8CBxaKaw93hcmGl+XJQ
es+8L4WUOBXasbegNcIwhk198n+fONDmy1sH5WH2DXE0Fgp0frSvizJvjZIu
3uyZUMJxbGDj7L8bauEDnNlpl+CAm0BJ7nuLfPce/2JDUaBLCI+8GA9R79pY
KOrsR9w2B0AqSEgOmDW6o2lUEmTC+j2m8g1x+hi/NSku7/3+8gdgxgMxRpgY
nW7rmxctGHChAFwZyf7KJrpllqeqs02Qnya5szL+PSz+hgf7ZvNJAGLtf4Xi
vudJTShYC3F/5S+ItDVE1P3xJpjc2bASrTxaHoio8ECBnpubU3PZ7Aq38rej
vqvFBHZPdZTD1Go7KdzMABNtXlS2v4Hhmn1DNZHHyHwWGZyhj1AvHh8F1ntu
mGa5TVRgQOUKmkuDOPDU84c2a3fSnra0VB8hua1Yva29kI9kJR4//xtPuH2k
IizrWs/ymugxdXbDL5btECtebw4ogPaZCs+2fcBOyd6H8l+8xVYSVRev4rWP
1Z8AzvjEgFHhbri/p/B+fLMf55dekB9ZnzjWz88K4xRdSrcTG+pP8xh4SBPl
CLZiqPsNygzoNya2plh3+cQb/af/VX0pWl2lqjoadzaSFS29+ML+EpP1CkoE
wGIGjqk+Hs07RJCunr//zSDeADaa28dpfM9yaOmR13BkNwznWqhNm4c1hxES
OJS5EOTNrOfaCTHM4R0izebFzAb7HBDya7N4aK0aWrgB9gjMuLLWFyRssoIc
9plgaK2Y0l61JFX8doDPyuuo8VRKRxRdOP+gQu/D4ea5dbMoq3bDHpb8ULw2
jJMRC5frXJYlJrxcesQtlPcx1RESCO6IrKZNdiRoQO2X8A9wplr3w75cRU2K
mNqQQtIyuX7DbNPJ6awXJrss92FW6dGicVzFHGVCTR16VPeGY7gaQgzp05ac
NaVR3ZDTC7VU1d8rQjEJb+fTNiE5rmqab2EUxIGufagCvEntpcw74pJepZVv
VbbFGQ6+0+HeT3wUIXerQYHcAz2cJfyqPDlL8k0uK32Bb9S/fdLymx991hlL
3zTvQcim8oKTKVWIe4Ftf7QtyAgE2twQjPWBl/ZZXwb3sV/y3KPcBAhW3Qlc
itm/R6mGwKlQlJLmIRn86lRDOY3MgCPB0XbcKbPm8hez1EZb8tq64qqiNCY9
ycpNXEgRLt3PzDxYZOlmQAKfYAQXB8hSr4nMqKqUTL6QLeBcEOL4OIk2mzv7
CcWmqJdAzLrUlim+WB1a4/MRNFlYo0O7iyT4OiVCNKuKMNuo1UvGpHQfqZeG
JuibPrHjhaRbLlm4L8uVr3ZjxSfwvFIA/LKGFAvHa+godxdoaPalmG3jz083
qDpbZ6YMEmzmwglsgTgqfG9SxKWhxz7CtLGLN7jOsB4D1H6Eyx124tGALdlO
2QyoAvZxkUsj8ryt0/XzGItsTSZ+mBbWOVksNdhbDgNegmEtRSTcqOe3kGAM
H2IHZYGS+d3nVHszhuRtCsj/l3FKmMCdY+se7ToNVBFhMH/2jpGrJMl69xgK
2cLly8TNtQwuayNmgmjEHqx9/5+QItcZwZaln29mX9t//M63bd0p0F9KnmfN
XBH8ovWXnpsuOHrisMbbNdn/jlktE2IZpL+yS4KMa7N7V2fb0x6zviDoFmp0
5hTQ55v+b2RY/fDhIWmTUSHG5c+NEvp4JZ2Rq2wLveObGl0bvww1tjmw+1wm
VMWZz/5Ov41nQ27Y5mP/z8vpZEbUk6b2j6+o3KV9qDhTBkqTkl4nKnqSQEP6
t7imRM1TuxyWoK58+W9jDEyyrnuVsY/dEUn5cs99g2D0PqHAnUVaM7jiZuRV
q5jFsy6d61ZxaV2TIU4DO+96UNkJqnRmVkPzN2jCNU4dpifCqBfVClKeDwnI
s2/Uq7953tDQ/oIZ0NVcExfFfhX6EGhkeBtiXt4B4OLGu2VIiVLDf35HFUt/
lgxXxTOoUxP2I3vl29fgy93WI6A+Y+xwXfgE+ZSjzjY3Qx04tq1boH2W9G1w
6/bzPalxtDeW4H25MZWlEgJ5/rZPlIFO2jk7CpeR7bYEU19jPcS5yxq3jVBu
+KAbegeLOjYIaV8S3Z7zfEKYzOpHmEp4CisB+r5yAqa/gIvdKLcxaWJw9rtF
0dSl9ZaX9rIYZ4CPV/vrWfaa8YP3O0u/RuDopgnQTlsjufvqTsYWVN5xba2m
z/+iJfIzPcHNPJKPFYC/dlTmM52krAFr3U1uILZyh/9uEb4r7tUWVbS7cd32
aqUHC5RDgRKFVQlMmK7dyb3ePrPRxRDoUtRlT11jzJGQ8qN+Z9YSpIvbYLZw
C/oDSOq/SCVsTjwTVVnWd+KIYBFp9E2dGOVTVPn+jkbJlyZPp0DsSp1FL9vC
kKNn5isPA5giJAGomhbbM4zprwMBa2hO0EDeEN68QDxO4BGbMlFyd/EubXCP
UDvL9i7f0TGEksG/drxrI6u91CZE6j935O5Pl0xLaWo3jYWOgPULYEWDMl+R
EoaTjijvth0LR6P42IYIn6T2CbdCK3QGjbxXtiQIEektTIsbHPiaVwh3cRK9
EWNTeSarE0HCwAMCUBtI4b0vhvXhwnWJQmRA05EUtUaYjxHfJbbPQ+oaoX5X
hR+2zDECebei3+Nxsvf4osZ5JtdhRaSogGf78quPJQ0P1MwHvzJO6BbGL4WG
r7hf2KNILXHLdVOksIE2VnCzEUeul5RQOnQzxYBKUjMbjRP4Hzwh/iC4QfA3
+I9DtYiYGzNWmMUf5wGg1bKGbcSCnXEeZGV+edvzmugOzRaEIZSgZYL+3zQx
He1bDE9W9IdhQbQoINi2ZMDckWmKlhXqoxv15nBOIGw1csfo8BWSqWOr0idz
IwQBbK4rbUfP1YWHMOl2UO+ifXCqUJaXUPFlrCgJwMmsKWJpvbLgMVenEjt2
sA3YeMsdwVHzW6VcTOMTu56O89uUUaeYrKuMbMJYj8Jp/Iej/7qxBRjpC9Tw
5gPdBssYJl0mlG+2Yd/p7Zj9NmApIUFBXAuHWKs3owl/xKDL7iw4Rx3SmVQB
KticzyQLClrPBKCn6fNea0pataDdAj3KHXmwac8UNbkMJiJujOQoGskfFk74
uGfWJnREUo3AvotDWzvHQcXNA/yUZ4BEw3Z8tmiGZ6g2hFX6yst3WerHPrhP
7ikDEmx97qlrT/ulacdjZ/A73yH5BPqAEc2gOBegu26FK0y+3d/te5ZHkVRN
Iim2mItvpA3moq/PRHw12xr2EfdRAdsHRy/KkEnIog/tjmm6ttgXmKTZPtsC
LvjPetVRG73oNUjHo3KSF3mYFn8kadQ4PZg024iedaEQBkVfV/OPqp8s+1PF
HVJhcVc8YB3MkPQf2mDZJTUP0bFWa8MXPhTYmwnbfzQT3Gf+1Z9anmlS5sd/
DLnJeETRYVH8DVnuOPM2ota/J4ZrCCjteZ0DgIZVnw9xRi8yQPKzqV/x8ocH
J7O5slMZXmcKra0vBDeyYPP+2S9qdfpVlpj1HdxF1RjZieCoUJaOFwTMd2rK
sL4qPM4xQdSfXyQO3vUOCilNKCb99q5csHibXr3cBige+KATPXxLzvwC4VAJ
1ENG/N+j4soJ/zu5vimFYMdSbIO7ofTeY3RKVvirwIpQVixe7k2xIEiuZA0s
JnKu7ySkLZdZRwVq7SFCcJkhnR/dCFE0bXcyS5raV+kfFfcHWBBqIfKnsT6r
Qw+0WJVzONYPhQPN8W3KXcYL9rPWncOYgIoXzz9FE6dgHiX/Qf7xxuRcdywn
r3EHJpAZHheEqItQwSyDm2Azglh9tB+JZj8r2MNVxWZggFXPwNebl5LLugQ+
jqgvvxWTHqELYSZVUfzfkU+ibper+VGv+iSgPCWa2AbtwZFu/fXZmSykSr7f
q8bGHzTKfaNmgPvh7OVC3ykjWNuYXAdsoI1dx4N7aQquot/gdW18qwKHUcJe
vkYCbgoKRerfTUyb/0uXYogfXf7UR/JlKUynFwlSr4fv57PjwEjTfvKM/UHL
lyVP8BDqB4T1kHMr7CQl2Rqi4AkFR9Y6hTittvOJ0ryfvs7U43zUasIACj3e
h3ETy2ChFy0Ey3f+e1R5diQZn2oudTxt/vCBmJJaZfJfh8ExxHOXWh4EYTMZ
/7g9ybL69SpzaFRlpANpRiJZ/Jywt8i2YHeuJ/krMAlNsRZXS7DvhbEXrpQe
IEpOfIIankaELbdTayfQkaTG8h/ExOP4O5CvpK6MLQ0Nf0yKc1Y/qMb5YwEL
oKMIOTRQbCGP5twYZ2GgxSQJqoYNiFTdVBYZKjaEtp9/GHCxkoc8pz5qRz8e
fT1vEb62TI45p3TcwmhHLPQ3IC68K55IzBe4EaZ5LFfHYRrMduLe2AfyUWcF
VWTklLibRjHLPTzBNIxNdaWMmVWTVfxEacsscxkFt8hlYQwNTZNiXYxXxaIu
a0uVgOc0/3ZMY0dwEyfY3w/0+y/mbx/Z3PqtD+NyNg6uNenqrJrXYHBuDfEx
raSgND0z4f8M/surN1QW5py6Icnd+5IcRd1PFiJHI8me4IPA0JPP1YgiGvfJ
92WGgxAlifpkTIhK3hjGr1RfkAHgejng0/G4GeKEPHQ7RRH0edhtinlTv/xD
sHboVMiS49k0vfMLXJwrcObGhanz5nCOOyfXRWl6h+TyUfSEzvX+S0KervkV
nasKm1qn3iDnmk0VXuE2jwPX/h903JsXUk5mnkCIL8roJ4NTj74KZzHU2j0T
p0qS/FBg0WTupqLQByyKjxoj3wHpnakZeFKXwKrqed4Tnrx4ruwLgdTOngKG
E+0QE++c4WKampsoefrQAQxBdVV6fVr3c7nMsi98xtQibj+k090S+tr4EVTO
PA+lyIebQ7z3zpEKmuDOTfeP5ymf/02Ue8bBj8C7y+LHgOeSBwneGAhvUdC9
vmSuFY2+oYOgOPuEIHr2XnuvA93mOim/Rzl1cnw+9yFY7f4mEhYp9ZEfGMKF
X2VsBHGQKuy+RAooql5QmsPtoleGdY6vhPv71JEuMWrCImngOTbEZ+nNohDt
loj+YX3AVJJ+e1axJa2ndqvrY4kEqXPdCJ8mmIF2oySazD7MsxVnO5wH30PO
+BJk4x3NtT6TgfFg36bd1MWzs+OvGBDbMuaW6gFvGVN/5nYkQ1XoLWQ1n7zw
9gTcoL++HSUxggWTurQBYvFLwu8u29hQ6zMEhBppdn+SiT5uBHQvqthB8Fwf
A+/NXG1/yDCAMJ/FyJol3vXgbZkXMB8E3QBU7Dzv1xq05ch6+LMKisIxmAuh
WjWs0vH21vhmG4kAaDH2xgMpSJYblfWy8G+jHv7bJmglDU+5OZy1pkgVrc9+
UKN2dSV4ra4KOGMN/MXeC2xm/Fo2ByhYuo0i4m5JnAnTCNKH4g8BwuyY4yZr
FfcjkORUznaw4DhwrN1h+8vgqwqeDD2DqKlX7c16z14SdqM0pz5tPaibSntT
v4wDRsh/rknMGXogU3dMnaQTuFzA8TPDd8OVEZEurG28lPLN9VRLoObBMHDo
hlNLN3StqI/Utm2DtjxxluhwlokFScSVnTMqM+SzS52ZDLW68X+zbfRLjdnk
N38hR19hjRtmYHuUYfn0FFGJLsdQvCPdkTTV8asMvLAODKy8y49ktFQQ6He9
UxI6J1/gM21u262JJhI5fhfrNP0z2esfYqD556L2yDtGCn5i5LCavBXJVVh5
vpoY8/Yg1tD9vrGoq8kZikYm4JiT8THlQ9lm7LKFjYTaGbIE2dTy1H0QGo0t
MXDpdE9plmOKJ2EBpNrP5jTxquM52i4n7FmO7BTDPh6/4YlCF1qAqaq1v/ID
sqSQSrnYaYXS5A+dZogWMuuPuF9PXo0BidJhtSwykeDEQKedL0CcAz9kC/FQ
ySWz6MlvQJy/knT4fGI6Nt/+Jjm81TKMjqHaWrgTSWv8sD/muq1oKdKmIUHs
mBBYaQV/JNWbN1F9ZRpAaia7LnH2TxCyW5gNhFDSi9VpbwQw1lZhHiahb+Ta
ciuHz4Zz3D3lenbYZAgwp4FwLRpsg1VsSJmjTjr/Z4iy11Y1B+cCzX7XNMGi
loNgLMFb4qM+sDabE2MuCeYtmvKU8gHD4qHREpSKerM9U9jTTRBpoZY42EIy
QOLGbNMbjaJkcNIIkF+1bcesZKxRY9m2Tnwlq94ek4Jb5k4wLySt/fINJhXv
fg9ts1NXkoWzImPTo+5OENH/UW2wqV2+8ZzTMR2tMn4547ail/DKTKxs431i
Sr2hKs8lhoPis4PjyRhbQ08YyYhKfKir3XbdTyPW0/8lPnEp4j80EZgb6riE
ipET7Wf1ky1JSDsXdtepnH/ge3ZyOgPbdqdlFeO5p409Yd4s23RVQN7TAYSY
7DH9efsIkrxORE8S0rjFYX5u9Lk3yCbcmO9+DAyAUpblBM5AwyJ6paHPvfE7
9d8H8Z9kyqbtgyIRMo5FqOgE/+xw554Sl86z5Gt/++6ysFzVCDy5oAek9Ahs
fzcA6LDxHfuqDooZd3DO6xQWCwkJbUH8jBfQFgYFYeneN6me+4tqlsJkkLzf
l3W1qCPJH1S52EPcwNHFMJGWM1fu3dy7s2GBwqvhMIKdavTgm0QGl8gVWD6i
LKOjD4jxTVmGFAwq5B7pC8D7E2PMF9RB6ZZ4+xlh3x1JDkRSiqGdsXSChMhi
I9ogR4MQjLiRIrQu9krAFNoy05dTHtd+airAe7J20tc0PCoUquKE8JWQwbgm
cj2MCl3g4qakg+Cq2cwkoOQRVVCmaTAJAAGx6lltYvnrnKCdwLVislqQl3E3
AoiC3CcWb1nhzidFmN+K+FmRUl89T2hINx2oGMGo9PoqVC8hSiR9xsGbjh8v
FPriaj5CAwKp0/FehGce7fhUC7ANMjtt3HgLdFiKAGPm8pK8vRayXBhoBS0V
M364+haDkHikDjSslnwJmnwV5/EuzzBezp23aX8jLz5GnWpNBP2N4e/LSRp9
AoFGyqH+i3jcJ8xZiv7y8oNDd0SleBt0wTJmCyq2fgFzLFB4vMsfwWmbUvUY
JX3a7hVhlnAuVgiE0np9nsFYQAS2Giz0FgawAOCV9uw2GYGl0wdhrKtA0heY
J+TJWvS20ZDzRngbjcnUx2+I4ecSkfZA5O8oK5j7EkNapFdVAAkaBy4/tGbj
uA+ngxj6IuJifuz5UHvnXedRVbAwlwoK/zUtlsQ9NiCM2dlI7HRmne/smx8K
8Vn90/BF7clbY/ZwVpkUdw5MYY6W6Ki8yAuscMLRlSl8CTvOFGZer5HFFKDS
sXVlfziihRdX+jvNaPDEGxHv4YM7lVyei28FNkPLc1B4undjDgPvb4Pmk0/N
qiRtEuIcRw2cRJpQ4iZm8AJDiG/DMcxxmsPw3of79XgFeNfQD6IkdcmBJqt+
Z8YEQw4mPZV9V6sNpCtMIO/SKGkzLVklfoNp7XMTIGEMKgIBZvfT+gGH41Db
ehlMfhy0UrLx1nQpGhi/uUSZ0rBq3owimFsU04qMNRDzueHG8pWAnKsryx14
L3/HNVt6/0e/3bMB+4XfjbVreHp5j1kmb3FF+gJDLB0xyelct/YLJBzYMxXw
olnb4aEqTQbejmJLecl4vsdiX4+1CDxREz9Of6sQ6PcTTYNSWCHhwQ0qvPez
L3PJVldp4/P9gQTqYhvkmdACi+ebgvZ2RVIzXglq3tIAkykFMtKqSpG2BwQk
wu3r8FzdUNU3NI+YzckEckzk0XN7+LR7bAWWVOeeLQmASWBTsDlrkDzuskif
mb1MjFi97ga4IPqDEGDsDXIi+kEkkSsIOHqKZ2NsjFCuUkOqJl4AH860X9YN
kIS1K6h0gPz3FoIcMHit/VBO4Q/lsnv1mPhudrfe6mTOeudkB9evY5IkIvzW
3QSJq2moJO09IUsgvirh/aOTXykDvgoenjbAP+qiDkhEYo1OsPPCpbs+RTLg
sTiS51yPVbekOitIbQBEni7SOWbWtBXyO71iYYuUdEXxe2DGRq1PJy5VGygm
S6nqw67Co5Z9+rCs1nY4omBsRvJ4n77+LSnLilVytIlk+b7MdfgVuDgphaB8
Kqc+wEDcrqjVa3Psxl95HbddH+W9prwStf/fTRW6aQUkr55y2LsVLfKlxu0E
pzH152E9SZG3PIQXST0PfNk2B8ly8O9v9Mhy5jngD6NXvVjh4yioOyehIJ9u
7G8RUtn4wEkwJLKAz47gGGGI41oeiApM+NaZz1z6XwofatO7T2L8QzF8p4vO
ITKf4dVwv0WK8FsTI02VDN1ZoQFX/zV2ycvM7PhnaLljb7Ygsym937lRFQVo
l1UXebmkhq+iPdJ49H5SQK5DbyRIgZqJomvYjmGLHqTwicG1i53V2qxwyFVi
Ia67Os6hAlrUbVTDqnIEhj2dJC9j07+jDGkkKkQWx0O80hgHcjv2D888tEml
o23qCIlJ/WcfQkLcW17f7xzGQ1syGcS0QVaE+j+SHgrm8370lJ0q72CWq2p6
P3G/TbtZ5hZYShDGDkDbkjVDWyIyBLbwGRnL2HpVuuXb+TXbwGLZN+q3l63y
wHMk2anbXSF91QwjkuJgm3ploGRdxmL8YyPenCbeh5BJ1AfZeXYeka6M4v/P
yeaHhqKNEac0ZSM8oAs5a3kG4MpSJ3U0JnocUKrNxE2HRreTc3m5lHGPrD0e
eqccQxgKBo8zOirTDSkX7eS5jsH1FyPPfF7kRs1olSdP8mIBZrKVlNCMMl8m
uBFPBdy3ZWYHF1pOfoCjiVZ+vBCrrxMrVB6NVxGO+KmyutgowbHrpz7E3AcX
bs7ClkEGp15Tm8EJ5Gmfj28P1xdBbwYkpKa4xpJ2G/xMWcxox5Xbvo3wUUud
+gmikMFZYEyqLaQQYjxbh7QOFKdPEEyyrs9r8LzFQQtDMirErTzv9DE87ptC
00p0pko4XnaxkM16OP03MCh7SYD6FeAwyiq14vnQJoQBV7p0RfBmZe3tt201
iAHo9/PFixceUbqnVQdhtAzDEj2t+LkEKDqFUctgwUf95TbxlXNEx4ReCgeN
tLGAFQ9uOXNS2cH8En6tJDpc+IIjcUxWCFxfDEmPIEK+oMKxfWvxJh1q44CL
T7RqMJHfUX8jqVYz6IoyS6FQKO2j2bddeQHCv3b9jC5upO3f3Bua9radh7V9
jmzgqA9QpPqlHd4lZ7Xlf0Kfjy1GaDMNhx9ZtUVb8f9BE5ZkmpFhjJKHfXCk
8g6oj8pl0WNqv6L7tsgitRXSFo3wa7sOl535+mj/IwGh6JZGKDknusUtyIfQ
tY1SBpSwahYHS70eyjNouu9+lahh/MPCxF+LSrhFv1R8jTv6Qb/nVreoNcEz
I9wuiHV7SNRM7I7FnUmedrYaKCPi9yG/699XybMfMdYJAqMmRK5MBsREocCu
aJJP8YerWtmbMotlNMPlo1XW4Ipuj9yxdl0JX2cvm8ZK/3ZknVM5QNcYp8qF
S2aYEL7KO0CDaQeixFlv1pjOJCixrTE9YvLQSNDh4QVBMs5d5jT6oHe8iFeP
5Ud+ABFVzl6wl+7dhn5Sr12oI4/6IV0ZWU70D6oaO8w/x4Z53UFzt3oAZhfs
hWLHDUpUzDMjACrEjozSZdzP3Wu8wLPn4NHKIU92g2y8zi8AsC3FiWu3zHux
oTW0CKtpkION2N4v98pMWic629IICFpquwWwbYhcgxwQHc2umR6drELDSfvF
tSa20SKXXlvB4mKioOlnhc0muDKjycyG7E+WSu3JuGWgedkTFdVtk8WZl8zr
j5nsc2lB0DjbFyerN4EbNfXR6SGJFStVVOr7HaLwZSKJjNzMqbdUx6pSra+D
bijZNNtSCF8IoQLuaBcsOCkpjml5ovceEMO1owCnGklZsUsGi7GqTyuxPn/Y
h9+5AVbchBItwxAb/yjpFrwLZHaILpwWRRIOXFcCuWGRS8KpxSlrKwu6v1Ac
lwWfUPyzf3wZBTLrufN9FJ0clVc6xUmtrKlceGIH6SDGnKznelVbn1Nbicro
RRiWmRvx4+irUnPyqPmlG05GEr3LtjDWC7jzoLdcpq7tXBw06PM0HQ+mrdzg
YLwGWCYg9JX5oUvPbFqLlZsj0fO33zouNdhaEmJF42yHh3TxLU0g9MVKtuOe
XaE/fWkZfuOFPLtL199um68oJz8GN/0hDTjcq6EB5cD0rK8Nr1SOwc6efAka
dHBYyb0u4E96tTNgyQAIFQnY4wIA6s85jq28E6MRJfEVci1hjvRExgv2P5bq
pbFSKiQ2kuQZk638Eq9IGNhjk0FJnRpu1fniDUH4a4GLwXj5p+W1PQ35l9N0
aJZcS4F/agW83VcKl/2XW59MskmjPen++4ACdeFLfogqYJ+HpKqmW6qtZL8I
vK59zRzQDTLXmyACqZC8nJ+FOhpFlF6Wv0CgtZngeXaeXnXUPiWKWQpzLbZX
eHlaAzbE1/PZWlRSaDakwNrG3SK5GtFd1NDyFmV+KHgJww3ML7+ixNmqhmeY
87jSRp9URtkltoB6KE803zbZU444/l7EDz38nDu7MFsVwfPaRdp4WRkjeB45
Q5wyVSB6BZIsq7zfmJ+mxy9JI71zmuLbGaCae+C9AGKdwXK9ebULeQpzNG2+
QiU9KuZGY/uQH7hd5Yuk0/i5uaShw/YzV7HNPO9pCJEDo5oDoWgvxqf7UNo5
p4FXfKrYHOveNdcbEJUYHVVEdbzjwy8aRp7qWTM+E1k7LJl91jDblzAGmxAG
yYC2TVbdLMhQjgfnB83v2NnWQ0zECCfAs+lYN61CuqoSq65Fb2so1Oid4fL4
4cbBsng3LnXsdh8HXlAdR/xz+yXZiuECp9XfoJ0DEA7EhL0K6fvepKwCe+ga
KnhApUnPrZCkWtDiL6I3Z2+Z7AvIXhr5sNGRe0rPWqlsqya9Q7tFuzx9G1xc
0NjhfACC2gA8thf8e/quEsx0MLUAl+f8YTivn+WPovlkibh4Gv24LC3rI/Js
DOZ3FLrlhY+MHLFcypdf2XS66duQLB72i0YZrBbmzAyBN/aUMbLBxshWnGh/
+KJJ1k1oqRTnXb+lEj2OJJ25lj34XZlRsMNc9QCw+losGDTSODAy2JSaFaHC
wTZCoNlaRc6v9KJGiCq/FHMxSCScZKENIExvBSxdCMfaHGEeRhLfjWxVA/mg
6SB4s5Rwki6ZVlSsKJ+00UUahFwQUbNpG5Eo8jt/MEoZA/EW71HwsfEG2Pxp
YPyzMpP6KPXbHfuwdUrUUx1XcYDvsf0f0bKIxNrFLqA+86GMH+yaVPv86C2n
tsMkdX09/YJmwWFEihpPKIh9TI8Kzjy+CZYlyVoQzNqcmKKPzDzLMH2mkLoM
jPQHibQNqD7EbTNzRLnYNWG4FZ8mgd5SP68B3pgjPA83vCPYRCdto4pNaM7b
BAOvhqaztdf/ySAbLxmadoRf0bwcKRAYzTqN9/fZJN1hACbzA0eA6YFJDf6r
lfILHyTHgPyHvklBoP738IW/3lUcF+yMXhnbxNJUnCthwTEKULWJBSm+Ltq1
XAJBePU0DJefIE+juqx0HsaH9BUmQylrkjexs2AG2etFxYZWWY+y2g/Yd279
Steb9ErotlZWuf+mynSES4DJ+Hpz6BLxYjXO+C5y6U0Gdl9ih602z5zBBcKq
24gzhavRn5MlMkXTEDLLGLP04IgqFmG+X2NI4pZvfdVMMyn1QzxMc0OHaXri
nggM5BuaImd3FRrc62w2GFV5q89/4LZZzAl/GIGOqZZjVT6Se7jW81+mV1dX
MbUL0Jyj0k0BYNxVEHTlzMh8lA0Rtdkils1fnJIx/+1MELbrC0jkCUsNTI8Q
4FGSARqe5Qa4EUAK5RbucevHFONGYNMIPm+VmV285EkYFkgAp8G7v4dxHXvA
Bf/fY6NcSy8oUS4rIvz63gKI74mM6aMHR/WnXmvMmRypP+coT5W/ZsxpXDTA
pTVzWJcHdIlmywI0GDThr4Ii52gtcV7XEmIQhYmcVBWKJpBWcPRzM+fwFe2O
InIGWrX7/Lk0KoOYQhSufc3WSOUZxhGqHjUHWI7Z6gdZGS7ktyHqlvSUPJU0
6CXJorZD4v/Z2l/KNFZU6Utq0/O8tqVouwsaltPiUepgE8YmZvYHyuu0PUZK
jnh82rxxgUKIvDnTsiYzGyguP2h2BOP4hKmbXNP2A2X1pDVNne4EUU5QFXD4
1cLLj0YF89NSqjEbs+1ojUnvUkUAe7ZUXDuTCrFJvgrN7Et/CumF4jree0Kn
7NLWgD8B54mnQOt3FTBCYp9dQNX+ee8v3gW8joBVGgl5Iafv+lZ4UknUGOOd
I9mGieXPTabGLtimH0PJoX/FsnTzd29L5ovRSEkV9sVlXmhPnx+ZdJMpSaxV
ZEeV7MwPB7M/vfsp684rJa+A9QaAo3hL1rwQR19SFLXfKHhfaGRYncvKGLWm
4SOcurl2RAz5tqHE32yFfFB6w6SmLPFDkEaZpPyWcGXyb9hOP+uuBtD7ShDj
ug558KeCdw9iXgiKOjnnV4WBp+jy+c6ti0jIcVQ6NMWM4YxguYOvQrf64ZQi
6SbnmbVuKcho6E6V0sdwGU2+TpcjO9eu0JgAJwkwG6v288XpzHXtylWF1Hwf
R1US4EvDUtaVHb1Kkp8iSzT6GWaitYdLWFBSHuAuT+H2ts4Z5dPQfaU1Ns6A
xkAiOmWlQ/C9HwUNbN9R+9L1RUy3ppESHZParXVgiu9pwzY7M1shw0gnvJZp
csWGL1yxom4CApyFTbLeNYw+qyIVHQsSKixxgOUYuniXoe5fbQubB63zTeqH
FH0zsW9FfmxqJjsjpbuwbqG/l+cUECMrPVwjYidu1tpzEEmPCBe3syfB+wbV
k8PRW1+NihP7LSc+VmUwsQMQnOLJ0qZ2URHqkv9Cg+t+I+B3+WPV2IbKWPyB
bMiM3Ii5X8DABdk6FNej2TtqefyLVGiXjr0NTtonO8clkzHfekQ9aT7LGc7x
+XLUxxH4FmE57c56CrJJ+azs90mz3jdJyzv0d9PBAfTRhbBK7QGjFdadRgp2
JO+zTJuFHI0UmfiHKWR1vtQvwbLTmO4LfDUwZuq96FtauqCS7dDWOjwhQvlG
lsxNHa/R9hkPrBV0CPLeuMHzWVJIqrODuITAVZNgZyxDKfKZtoetfhrmadXV
hv6EMPSzrJzRVyMiDgFr7vbUSXywCOP5fsbCvJ5PTNSiQRRiZGffevGOB7Z3
2Bkp0F10jCBmXsMPlZvcahQDPQN7C4VJZPmpi1p9WM2318Fkxu76FcmbFBiL
VHeeoK1x5nM1EIytwJ6R+Lj69d/alg+as3Jaqrj4fau41gBZ0TBmdjUpCIXw
3/E8w4v33IUMTR91xPMMRg6JCQ9KmxokuEWyIDlx3QzCEGg4zPGRYszaAdre
KNSaLo8oGE8TuSeNI68IXEC8uZoVObEgEb+yL2HhH/fDqSrp3wFtk1mJOKtq
/+ORHVDExG5kEscwyHm9vUYHKn1QpbnyyJjzemGtBGEDP2QQPx0UI2V/vMTp
yQiXEW+z+A836MjiuiV6AlCr74Bo1Wn0wVL9Xe3zYiFsL5C8HP59B3y3G8o8
AgAv3bYcjpkeQEjJHLEy3QjjVaeZCFJekFA/bDc/aaC/TLtvOL6tZYIpgpA1
5FZjMLDmsDHNsRH4Z+J9Frz6cnolSyKuEd6N5PZ0tJmQ+WcMnLdEDvoHBcRu
IVW3KmGGoTw/oyUrUGbVBUgAf0A7d+TBNyV+DBxQRfj19TBbeLmWe5LNmutu
62RtXlPAjihwcUp3IYa5Nt4gdWutmaSCefQPzNlEBZxyPSd1IEdbOat9cuvJ
JOfIAf4/vhFUhUkj11IYkjRBBXAsfL1DM4/nsmOQKqRyAVgFHd2gxyOP5YtT
gRVU8QXM3RJ2zo4Irj+Fd2clZ5vaSEohhtiaKAmNvbudjDLD9cWH1wWjqPBX
BDDWgZ4BtLr8428W0f4tOq/bMPgdh9SfxXaWoUVaSFqgg7g8YoHQbM5Cg0tl
LwUSUcKAWivs8BkJs8P62PK6Th2I228N67EjhQsLEJ1FZfsh++H8/sa+0Ita
WZGlaEzwBw+nbn004gEPMrgNpNpt4myigEn7NOetWi5BvAdiT7ecAD3jc08Z
9evoI33cQF8r4WXCOF+HBkTxeG9clSdRZmdA4PF7YJa13Kce9NrGlyCeETbP
ydyjS2h0Eb+K0pmHGQX58fxggU6p/mvp5nB3axL5yTD68+JaA7V5F4J96Fml
rtet1mOflrU4e9FwMhDs+payrFfm/XGh9PNA+Xqcrm8l2m0TmSqycoX1oA09
PZB5/NF8Uezo+9+fZrhUgQIFyQWJP8dh8Tm90ZGSufw8I9JAxBeTJANkSt0n
MyVGPAsT0jNTK687bLlk/I9pOW1xgUatvZq3ppCV9KnRCqU3hdzsstEthlHR
19mOdcdswN7HAKWH10W/lYd9EZetkHtXPONGo8ED75RK6QutjZXscJA1swW8
e8uVGEWrBUeGwbDAJmf7tcrcCjYzjQ2BjFM/vVIGlBmsqq+F+bZzGQ/qkhfq
JW+xG3E9Fkv9EQibTDoYWxXrYvS5ahBSXfXUjBJBkzXfywBJFZ1H9By14m+x
Mm+ns6DrqtDR65YYPleeLgO3+HKEPk1eem2BwG73/NXZ+7aCxx7ZygL6Dxrs
j0ziLRIBAJ9nJBYkRWQlihxI3fVwZGmQgpbcEJop6OhWM+2yBckNumV7W38W
dYIu56meBgv6hIrrnC9VmGAXbFq/MjRdTVEH9ePXiku7TMMHR3L9qA9P6K1Y
fq0ZNLKImUlC7PVrkeyxTk0EmZSew4CHj+L6YH4/PCfY1FY3gfZJPCxFxEA6
1GOUz1Slw4gTXpw0o8yjZWb2iicy6AmXUwiKOyVD0gtaApn8+p0F2N5qkdew
UQOuGNJWUMVyIDLjmY3GcwOn2NqDa3W44EDvmDdMu/zHxuTC2GjjcVaEQqSx
B/lwBFgQthJdkeYVofKGaHNSQfYbvMthxgiU+K+7xWifhGOfaG/WIve3W+KX
tqbXc5voi9xvZ1pM13OvLuU0cnHU9LMfCFvIXi6FCtnMZTD9O9cv7jU5IpzY
HWtP7H6f//yZqisVSsUUvtiJ/7vbzp42ue5hOVIkJErZ7I1lk2RSqHFdqdRa
Eyfo39z3BAlHL+L5o5AeksmVwI7q6Y1qZGoYfAANJoEJa8Oo0H4Rt5MRSVIU
OSsTaaH0NBMEsPt/WHbGK7iPAZ1ogvZg3aQcrlGtckYwbFpTsi/it5e7COmz
0i/c6/frJP58XU9CNoQMoVbMQH6sVbT2QERH//9988k5BkeOGrWQraL8gDYS
ZsnFm7RL4Xy4bFMhoHuXH67B/TYWYQ76CUwdTPzcXRk2Lb+vvCkMYGJOfvvU
srdfjPMUGDbuDkG5qDD5WBglc6JM2mV+KsalN6Un8WRZi99P5TbFyqre7UcZ
l4CL5DIUarUiI9EHbefOK/G54+/KHohkHQVAz7YY9QGfmhMokfAj3l/zF9B5
r1wWGG+UAoMKD0gia58yKnUjW0dLI+e5Xe08e96Q3rsz3EAR9MGO1t4lUybD
PJRPe2Q11CXehD8SGhxv31dgBzqIWiV2P0r6hhBa2Wt4XrfU/mpxDVZvmCWG
4vUICYc0koqfHfcLDdkxcfG3gDEoYWwea54+flS1c2TMi4rU5QdI5xj48fRv
teyXLyPa3ki9Ek47sbNfhY8QcgHTy+HiZpNkxGHc46JZzBRgaj/wW5ClBO+T
6fGOgGkvr2G+Y/n3LlT2hPlXTaVQcVAMReIOdgRAYaFH68dzuxukzf3bBrDz
DBr7jKmY/Ozt+nVHBIBak+BOR0SiekeMwhOeCFEgsl+nRvoUiNNw2FVCSHm1
CR8KecoCtxirZXBxuQOOiOhoJurM0AauFbBX6QmjXOayzSBweXn8I3MxuDqQ
szTtRPkp9Nsj8maGiHLN/9bC4C7Ak7rW+lAJVjDvezatOYBv4FgveLmXWpNE
gmSR6lzrgXLoyIYUceyFIZMqGq15ZO/2pUv26+8XRscth1CAzxUdNPz8z3NL
D3NUPuLGVCwGH6NAzOFPwUhQAHslve3k3jqE0EcueWvLrfWWfTs+bOLVY10K
PPjGuyBzaR0MGbhn0z19P+rVBSFqqXrXxUEm5+doplT8U+JJlqhRKFLGZFOG
IwQnRWTJ3RPnwOENh39LjXkDqho4vozOuPUcQTbREZVDum38VIfJkNkNiReH
ITsL5bsjrrlnomBGm8GzzYs2sFtAaz5Z22Ob1DVyb9x0tq2ARW2spwBOwqsa
TBnNK+bfe+5QiC16MoXIglvwu7z1RVTE+w79DEFGkfE7Efxv9pxRnLBJI6yt
V5a3IDmN0rAvc5XzxwvZfpcD4Rwl7/CKzyriu9EQQOZMhlYEcqyFqTGv7Mno
h2ljQrLj3YADB1C5T2RtwtR5AhXHMISRG1OUvzc9JhoIlLWZ254xTPQ4lLzX
+9TlIOFhGjTuAlGHeHkPFDw5vx31n+r5uXDp3qyYgOV87ELWZkK5HKyB0mOQ
2jf+foprBcPw2DwV7JSVSrJv5/0HrfTckaCZqMjCu2LqHP52VOUr3CmN8n2i
3rORTCSMHwXN246riYZpAP0NnFpiOc7kAX3Y8JJHZDt/dqMZixM4aMruusiR
FjqU+P5a4of9KzJSWAUAPGxyfmRjqnhI0zAtgV8k04IRxeTEJZnX/nzbLhB5
4Fp1XcJ7A1IRkWNFEgAf7IxUzRrfcE5j++zyLrrGDFQqzTkOGayZ48OWu+RT
U5Jk7+K3u6q/hTha9EdxwbBJiKHXvpD/lwwGG7PPTSCu1iHBfFN99E48d+Eq
m86JdNsvo1+GYaZn92eskcGQ4uy9kVJprz/SAt9tR88ZKvOggVpDhDFaJ+V5
TESrxqv1ZR88HNpIN/xW21WjDnDlQ+xwbwksvjg4JE8+hPGiFL31yzSWOuWt
9OkQTzI1NhvsWrrpKvEjCzAaIspOjzxiiBB55DGHb6m2jZm9uJziiRq612mO
1eyp2ouYOJ6d+DmA/vHEi/5V3Rp5fBL0F6jpwgp4sn2b/mog0F2vvZK44ehn
yG6i+3B8XmCzrKUhkHXmISOTwA5UF948f0o93q+hlIZU+dRLSgdtGP5Xe/pX
VKLRynmBUNs0ezby1QTB0aFHQFCP7zWjB9u+wQXyKVPXWE+c2wZ1ZE+WrO+9
H8p2wW4XJq1h+DUsrRpPxvaRQ++coa1GJ8zXywD11DQ3k06jzHZ+1lN985R+
7GbOU6sVT7J824DzcXyorz814gAVIuQgciSjj3D9CXqZNQ09mrGVgMAmzgN6
+PTlPsOr8u3p5KhaHEgXQpFys1aEYtEB0tznseXzbmMyayMEQkNAo8xc34Ks
hHwHIeuc2L3CUGotaz2XfS+GC4hvFSjvSNTkkTp/sfvWj5S+XfBUbYWM1LeG
1mPbpGuTabQoGY0VNuXAnEkV0RAFV0mzEy0n55v2o2vP/OAj6jqD7KTKlFKc
4YUrVLkCElC4zC/vfGH6PCbVG1crzMkf1i0T/HUQYpxc+GOgq+capVjVWjSW
c45/pTyxBcxjvcG26suR7KcpgXodglW1YGgFz4UPc5T0IYdLisnLCoKjaXcK
LcuKxWQv1eyJ4oNfaDJMJu834nbdQx/4HC2UIJETUIKJQAhQuVAcPsi6WxQY
LvGJP8y1KP/L6GjU2KyJSKCvSk6qpCD40DBYMNpHI7Ji9JBBS77Qnwi8I+eq
4YHKeJq5uDO/+pWTkDXlTUVtJLHghFglmadrUbMQoooPRH9RgI/HLy5hHI44
IR7dZTEZfTqjw60gnJ36ttUBfC1zxLHVGx5MpdwtgtgNK5KVH2PBMLs2XNrG
RONo+ENi+lvF5pPi97YzDX7X7Bv7VqtykI/Wafh8PdD7tLiu7rFiG7aR4kR6
WTZ/IaB530dDJtCKMdEg17QknFoMEJagcEmiVpf2aDZuX5gHfoxOd7HLfTOy
XErXdbis7yhh+mwnE+w7z+/Q4dN7hw+6kgjhB9NEiMPM4ARv3jCmFDCMwRiN
oF13NQ5v2e9S1mO0BelFI1Bjz9TTkQspKhmEhnOswmI+vRIrlM3sPdt/ngCt
UKv2E6QIjmF7EcKIu+JTdAABtEVxHUUGbcA2VCE71GRlu7AUpv0r4KzizGq8
s5m2LnUg+QKkjTr/5m+IJsAkDeB/ROEEXqPpnjUEedYBFE9FEr4p0wydVPXG
lH9KaFZ+TPADfMhc9yR0qaEUDISmthZevG+WwGLztGe1ROe2rFx1cUtHUFsN
m0RVJF+B8xEBh7h2q/0bvhiNduvq+429u8OEUuLpuSQGXwpIWEnyS5VBGb57
44FMNGtyQ9n7sw6pXNG7Q+9LJ8hkkFDNEouMTgUEA8Isouw76Wa8u8++d0MI
IQ1A7+4KD+kHz9mPrmu25W3D74ZVB/xfDlUBDSOjy35ccvRdEMqXyHh0sNrh
9zBZghvDF0kNmBMeFUy3qw2VNm//n1yVye/OCPsjiHRxbxbDJDCBoDU2UMXg
7CxM8v91sRE+aMjG+FGt01m+JZUvTcNhoFt9Vp+WEDjZ/EDolIt8SK17rSpn
aNM9qHpGD0QiM+AFKA4svimX5UAm9eGzYXAk4X8x7btIG2gzh1ZErJakh4i5
8fSQvDgmOUvD+4xfMF5flaZBElRAd/WgfJuIhR0154lyly+jl+eH9u8A55m+
RHBq7itjAZu2/+mRN+R9TAQGTAAII5NjlBxhgXGEtGsZBjBi7IqNRPXjkMnU
sHIgpwtEVd/GYq5H+IJne1QVNfYaERJrzN8bssYGTF3TDM6AmJFyzGfJgpZw
Pc2XaMGyi+QmT17koDkkCyk1cvIksgj4zGN0Pi07qLyo33w3AHxRYumt/lxG
GpfOn+jyTwzQLznix4Ewx6ITzgwieWU3sb1/ghEhPnjopnCOSARbG0At3VSp
+FDgY3453WmGsn5rhVynrCk/w+xDTYOYrfw9UseDUZrbFVlZq2OMBmK+ELfB
Xy6nvNB8d942a2MXKG0R2DKpAURB47lhb8/hxu9f0XPEILY1Ci5dLRAE0yqs
mJvn9X4XKUOjmyHQv36dwLzRBUnEqhznvXW44AaoDHaDqpTNS3drXj/iW6Q9
9CNZyEkoi0qZXENSRx3yIq919j/8UEqOA9ogPgKs74SlnrHVIh9TBXZWe01C
6o0gik5TKTVNV3IMdgPvFI8RAFe6cwMpM+HWabZFzRXKHwXlsEy70N6APxxz
uV8wfJb4yvK1L42vC7IhXCMdrDEQdocGFvHfMqZRiGHil9aiQ7nGwMOljZTq
Ilsv1F3HviBsESccmt5HTfuzsJqkThu3WERBnGJmH7AIJ7tJevP53mdk9MBT
ztE2kWKy69IGEoG9N7wscm6oWWaVanMwN6qJEKOKM28Mra5BDHyhpIjoFoCm
cW5cBnRwYH47dg+FfVpjAhVEw+DwpOvE05/T2xcVk/7OxMkssM08aCs7gDDD
rNNdE0JsJwLxcETQOPlVUtS3oZXEei7iUZajP/S2AUTBJa9W6ACEEq219907
KadOwf6bxfP1V8C82wxLDJcZivUgNucPrlQOVelVBuJWDWdOMo9pkU6/jN7j
/e2WwltRUZ8jNmxbc3sxPyd6KXu2tL88Y5WCnk0Sl/S5BJf+l5llPsaEsQww
tJtvuVPDEfAW7/VJQUW43tKTdrDw9RMUYck/S3f9P5SHKLTudN7v5S8lnRWg
m9zux7dxrP0wqa47eaSU+zKIy69Ah0iRw1J35s+q2VJUwEgWy7QvTeDkMdQp
HNopZsdEkwWElGXe48gbYCnuuT+8w2tftl8luR1uDNOJC19331QKk3bgr4Fa
nRwhSMgOlnozOwfeykCAYAuxM3aL0VCkv8jJd3L2yDRtdQePlNWMZ/EMKsp6
YpsKuj97Ng/BqzixdS44sGxnjT/qYvJ0FVv4u+7JKpaoGTXedovp56uJzH3W
PwV75erViKpqDe8V9cCfDDLFSm5XV8nUISM6bYd8hfiJsJuxI0RA2pBdEM1y
HoJEVyHfiLconGP8IgMx+OzNq6ucIMBTchC/7ZWmRUsJ1cUloInvua9tyN6+
sbJOKCjLxZldZJbmIjUECvCYXBW+A29IkXd0CjobV+8wvo6oaqYNbDfrcaol
UypBRl2AKpoFraVGnq8hSTE61sM4fA7Gz5K0GRUvpaY3MJs2S37/L9gio1Zk
7We/E4zb09TWDXZCk78OQeOz4qmd58eU6u+bXvivp4tKXKOD3rP49NZj5WoP
lrQw343KPs4bOSPig6P1GHk5xN/uininR5B9SYhP5O7P14Ool+RCpT/W89sx
Pk/mAkcxGQfce4MfS3kzxh3L+nkSA6fWAIs9kTM/5TshR/DJnQafTVlstJPU
/odmQVPriOwF7CCMz/pvqLqUoOl2SHKuOdFKn2HGr6+69P96Aq8yhaCop/8S
oSTkuY14b+zNNDWFy3SDmByLEL1fRQnLqhKGID+VVw5s0qiX17YfpygQyZCq
bfR3q5J31bA0F/doiVft4H1QPI9PFDLqJ6jmFxVA/LwTGACdKSmZqG0srPBo
P5FP2p9hM7cdiOUwlG9cD9DX7+l8eCblU48mtaXOnO5OQY7wN9LHb+d8Ru0b
4xL3I9WZ8eggpnEv2LkfqwcqoHElJEeTxNBCAo/2nE+8yfygKnV1hl6ECcoj
0ancm5Q994PKsUPBxOrAbnHuC9HTpNVYYnLQIQDgeqxbhZPGMdDH/xYv/T6Z
SaEkUzKHWZ0eCLHgCNKwFheYWxhPgV3VdYlN2fE0ai8ctof+0gKJDlKhk/90
Zru+M54fHIkqd08i06ZFX/tm3B+ftEP7eW/yUFc1CoJor2+qebEYhYaoUjRM
0yHqU77DwyPUGIALbmPJF5FPgkkyBFIMd8sAeOWQSkLqSzpIEtHVhOE2pw9C
eCzk0N7s84l9TcCmHUl32jr02vDW5xqhMNLfhMgT8R7wLrc8HLnNVOUacsVQ
X0VKDyr57OCIyT7CGYLsP4oFhvHhOvypLbAdKUFzhaHLdfrfBbpLQDRXCAm9
AHXmqSPenWuCjqzPAgUuOcs0B9WowQoD84tFuCcBrfNcjcLDv/ZIj0+9S8bA
h9i1RXRO2Tvde7d225wsU3oacMGypMWi0Ok7GjCRxpom3O3O0Lx6l+Cmdybx
+XnkiGfwb0mCUplhljM26KiX0DQeXdHfYmfY18ogpjJXaakhs9r28b+Oj9+7
hE4yxAPzRY6qbUJG+q28yarR+MfYg9bd16fqy0DcNNrBea/dERmF5WUVsT2s
89JEprOwFQsrw9n+LJuv+n3gzaB20N2tw1LqUbuu8fFzJamfeVmXe+1KsW1V
YC+A6RwUT2HWlH3ndN/qa2vL+zYVTdKbYmyMls6zStgfOm58hjYDJi5XpdyA
lvwj9IlMESMfpS8XxqLZgrupCXtjk43ZmrI7LcMed7rNyT+himEIl9WrKHNt
IwS9gGH8SvLDdPLCbk1TCxeQgwPptXeNvRr1ltY8J3bbO1my71fL8BUR5kWp
xPyDMtL+LaQEnOr7wKBTgdDKQwzQqAnxTYq6PiqKNBuPi1GAzhJf9Kwc039z
5QbXsNRGqXjB6oFmj8dKfpCEfQOIosK30s3pIyF26FhVMWMLaKrFzkAUCQ9d
OMBUdp5C3ABM1QvJD91uxfLj4qqLksQCe5M6uyyqJZZI+oKvbvTaZKlWThRG
Nz6Wb+hmz1g88gdnq2/q1FHvWetQiXE+4RzKBnah+ehmi9f7YaQszOvJBTRD
St3JfYj1GXOJGVSVMqAOZhRQvPGEh0hK8KD0s3mUAJ4Rq19Vlxfudr3HheV4
K297FTGFNqmPz8wgUdvb+eZqYEfKgBi18qEQ4xzFBoa7yWcOPq92ffuq/RYz
LX3tez5BS+vEnzvqT8CY9ZizoKwvtQKTLgnsfy6zytYejD3W37yPFg/7zZ9Y
G7sX3bMUyMFNTwCzowxch70goKGob8qIneuP5/xK2f5IwVUom4ZJ6xBOYmm9
zbocjNzkYwb3PrPT7icBYnYJ59xZsv/w/UTGfTgrRgHQgpFfuKPhNhMuCySY
b3m74jz9FhBihku+GK3DIOkSMOfSRicCZmgznn8a7Y2phdxOHmVvMRAf/f0J
8dAbREFD8reRVC8Hv9xzcJvQ+vYeeCjkco/eRsPym/8NndgI5cRNE0ZWTQkX
FhDFuMWJ9oZdNIEBUJEHKfgQCjwhiLWvHCxg89riXwIhE8+rvsXq65KyQC19
T/CFZCvCU8wz8MiYMuB0xyGaSt3cf4/x0T4d6jV9BII+/qrFkjT7PBICt/2A
W14FTVksWVNHJ3wIVUY8ADEYa2PdJw0LRXgF//T3WHtUukX1sD9Qu5Mc30et
/8cifac4fDUVPrZWLV/FF/gkEdg32xqD/uE0d2ChRglyIty2GNkhAKLHQUkW
84LaGPqrmqie2qKrkJb8daT2G7XyYOwpTS7u33QZxLfLEm/Uxv9dUP1QROfT
FiDVEV+Ys77efbDpCBRkjdzKHzI2nrP8P9Mq4EcTocvqB/NWwdjBEL/81oGP
UA8lfEKNmkq81rqqdvvupTtg9SGjNaDHd9J6yWQmufG7ClcVlLEyhPPy6g4p
45alO7DHRoIu4o+STAGBs9cMkVIBHRlFvePM470m6cxoHbFvbcdVzHyatHfX
anp5wFeLmSgmPqIhubMMXAi6mnHIipMFxo1/+xJ+XAAWw57lZt1abwm2wB4i
qqd1YJsPhnW6YsauCZP85WWJ+Y+bhoevyAlltNHHREhnJSLywupwkVp4AxU2
PMawMhgM34rX2GhKZyMpHxRLEYK1bZj8YIsfHROZ9UtRIgEaovcfPC0QA0HW
uFiY2o78koe9RXeP9ISeGxwAS2eQNbc6hpW1TszmswArYxR6IVZPLbFRyvO5
iQiUNEjCHjjVgcDQx5KJt2C60KtnUIQh+n8Q/Wi5qQQYUk4fQ5V+FiPcDa8d
PL7gCm7CZ+NIU3zKLiNy1KI+zTxV6wuBTtJv0FD00cZ2i0HMNl+VlM4YL7jW
af83/pL85rkM5qD8ZyQvNnlfpRNo/eIQft+9riMZsF+pi3PqvMXpKAZVPq74
EYE7kVSYmljqe2KtZ4zc54icbjXibV24Ulsy/qJM8tXnoHLQcgha4iyCsaig
cVF9fadfxphbgBol0n10TobsAp8xriodfozANptXkou85sSV28BU1W0moptH
4LH7GxofSOPTJKgFUblUWTra6SPv32KGQPKvFzdKp08bo06vdhqKbfJes1y2
Bbv5K5JQQsgh+65qGCJ7kokq+i23dYHqHohvOktr97fe68jkbhSXsm9WgKs9
kExnZ84Cq/Imyw9uUzx/HKMAT0uIR/Kq3Akt/FEUrSNFADXhaH69LIKJ5AAh
E4StiDi4Bo1XjyBPivK5Jy/QZRYOL5nngzkpt3gTaXdeO6q2lyqsNy1VC82h
VHh1MZin6KjEfIBQOha+JHDb6K2+mpml/vHB4eVTJuyo7N/oMXfW6WoPFh5D
h6zxskJZrRt5EBMysN/5Ty5IN5NWKT7g2LjumQdwQ2Ip1E0QWjHCDr/2rNuD
Msl0oHoqWI//IZAuyGPq4q9EEtyxF2NKjp7p32CQEOt/OAt/Vhr9ed3jcONV
9W765u9PfN5G5ZQlwXuZPha4W47jANQg76y7ynLJPuQOEnnmIrKor+b5woxY
KYrYbDzGFJ3SBOeER4ppKWO08Q13KbNJ75O1fFl/MIVb3+JhlOW1MjDnDRci
YIUe4ZGI5pmIX5jshn48Uw2YuRX4kYYD4+ryi4xaSAbdpIkPsz/reJQCc2cM
zB8GbI8iSinU0N0dI0TIPLJx8gd/tzkA/syR8gdXsfX7LE9MNOMbLLjkVqSV
Kj7n544AYtajrc98RCKoCLrREF4hiNMepma7K1v9lPRKriXvM3imqFbZ9441
ZRNtscGsQ/D9A9fx/e9qFic16hJihh9jiO4SONLKTh93UlAyajKvgLLDpIiR
Rv8tT878pECGTuyKI1dQindHiWFLxOdY4wWDWMA5tFkgXse337K7gEMgrn6J
GjCcvzSbf1E03Sjqw20gWtTRaSC7PQbfWlebVm+yMZIku3BwDbhAzi5LtV1e
k0E5oOXkxi9DnpBxVKrImimbZoopO9AS3+8sYE2Z6QSfavqHCTZNFMXVf6rK
hNFG9vcxn0i11DoYObRjXaFdgZwhHICCWrzXn/kb9wS5wUfnX8M1woQBrE8y
UV6J7GwJzcuD8xDVPi1hrg1gF7nBzdF+9qzVRfiBndi9cujNoPsr3Pf/7eRW
I/WgKX7BNErEA5mtFNdz6SRir+uPKvjxmk36Lz3LxV9wWx0iNLUtFhEPovfR
6cjJn1q1VJhQ/1G9qyN9UYVBwiwsE635JiE2zhJWi4Lm/2gjAS8IO4uqbjET
l6iwlcCGQB0mhpJNDV6xtyo44QKGRpLrh1jt3ZlEEM+PDe9haBJkl08kjQjS
ut++jzYNasg5nmSofJ3mEx4XV2H7VQZAwsmWRxz5nnyyuWNwy1aaOfmku8nH
sMRTgoSOJ7j2Oy69b7YCghHT+yRTOOJkKWoa5l2TvvPi5al1Jb/5i4h6LS14
KJDxIN/SRZ2Ze2t1grQjwZ4DJnkr/rknmIVoLQyqvIQJbcJV7QajIoIfV36a
r7MHWrCw2yYrFG94LFqwEJmlRNl51WtJK1TdaZoqcNFVg2aufpGvAiX0J/Wb
PJxTXWvEteK8BXI3OJT/oX12j8Yp2msnyuGD7nUyDXgJfide47IueU44g8zz
RKT7FrCA2F3pXNho20ZnQ6ujyKf0jjXDAN/2AT7NM0NOBr3Q54W0766EzOHL
molHuvoOenk3+ot0PTCwKWJKRadno+osGh399Q9XLAD+IAZNuSasfkVrc9So
v+uR+lZOXegavU77TnbIAppMr/+6IllF4iqcem9s412iXEyn96qDO2DgV+NK
y9BS3e9CDyJb5q/kRGUc6CP+fYyqroTW8AvE0QbrnrxE/zoaODQ/+/sUTQQE
zQXByDX5wCpTnaRYEfvQfxcC80R/yARtll6ZyCNBYQVi+BvnLzwbnGXxZWHH
a0qjfDkbHRfzC6uWXa8IZdfuUc+AoQqHtt0hJ8AlQ7PrwyZorjyqgCbfeZjd
bbaPkAg+rWErovWFma6xg5IynwdBIpaAm/mpc+aU/Yr9wvPZEqJ2HdC3iQyd
3N4toiQLr88P3i3gRUumFvqV1QBuWnH/a/dD8ZDd3yYUezaMrwC4JvPAWzqI
gjP+aVTnQb7MQ4WluxZeKXXSY6jLD6Ou+zESZVtRUl3tMx9ruKURQ+gNdqfY
buaSjiVvYpk5mV9FADVHx/XSQEqgPPpKzMYpX1mDtgmREYi3Y2RgUo29LGLC
ySi1gpV8w1EYBClWEqZ9ByKbagyvuL3CBH35CzZfQbjMhKgkHi3aWwTCBnft
9qnLFkMWK4jmzALVHCAd1cjem6yMQGVFVEArDTP8tvQxmh0TwZBL5YLF8yjd
pYpJFOC7nK+kGHOWXsXnnL0ZHTFaL0+Poq5lmmJmBycTuHxV3eq5+gsZpCg5
bc63D7oMbUWK326F7xIZNdeocCcuAONYC0WoxQ5/J1H/IzGXORRFWzSX6Eaq
HoPc+q4VoCPCddLxVwvGAZC8sEkhfGtLl7Em7U3aXkulAEbaTUFlf7mJIcq5
EL8v6af+vfPMQ8lndXRMOF190mhpT6TOR9M7eUYegVVAGONWTOSJy2mHMtS1
NdEmMA0GC0A0PBFmSvodYzE2dBDWcKInIjrVpfAaKk+3BZ9cD2IaChDO4lXN
q/Kw4szaMNom4gHfq7MJEDTWsBXYsaZ13GPUCdQ8e3r6+ot7ls/7nhNrQgXn
nk207+xW6HNZehX2HofmwHSKDWxpdCrP0C5KjoELuFAgMkdzcxT/RBBwTKFH
gcJundu4hMK0JNTphlVSfNCOCYdFdAcVLZg9zpY80UJfah/LDIHJD3UeO8gG
lbrUUnr4qFdBkZkCYw3tKiINtk2yj+LFPKCJO8JvP8Ke34rqZGxw2h2jo8Tk
DPecH62f3GtyIz/R+JSb1+QoAtBMc69wXVPGaewI5rPmymNHXiUNHEtev0Ui
vvOMsUO/Bxi+jte/ruHA3LXyfiaHvNay285YXXbvkkEyXMrU4D0sdYiBstb3
+vPzNsrpAWNZRcbGCdvEfv+4r6WotHgu8/vXBC6/JUJUHddIrHpbK2VLOF7/
9OWfh/6TURi23HB9/3rVXMP29e+1qhzeOcLjEd0t4UFYVybL5KQwyXEyKw1d
l9mjMzYCo+jaPS4i8rVc26JE7Ae/2ip4Pf2IuLYZBuyL+QHm5g6iw8Uf20Z0
jGzkoN8lDSUbby9OrxNKd8dC6yXdScTQexFq4jfftcyFDTKl3CzHvwV+0A1a
5qS7eFC/0jEYgYYeMhHabEcIkOlzFcL9lJwpD1plzptTF3HFo+GVlkR9z10q
89asjv4YcmjucxlDNoC3oJ6Bg9J1W8F/zCCCFBDgh2ZNiksK96DKmgbQRB7s
sUKJlaM5mr+kQ6817s0032lUQqkxcOylG6g5O+OUZBndhIXfgvicXcrNvZB+
t1GST3fotkLOH4DMAUus+Rb2AOArd1FMHZKKU37ZJGinBKyBl9zPh1RLgSzF
mfO0GeS5qYeUKv9EQ4iZ3TO6BUyjJr2hp/4utHh2QCMa4siPX8P2QJmefNyn
9ffM+VjUVYo5T06NdP/J7nLF4hH0wSNjQTHQI5woXhfI1OQuDyuw7iUAc+lr
dNKeHoH1SysXzRmQtXnAPpkVVa8xtH9UEHd2iY2C7gogPmiuMawRL2EXeY+p
YOKSvjSY7AvtXw+JrzikmdCY4OHJKso+AXmExi9Gbp5jnG0/r0sMv/fYPRH2
E/YVmiFOypD2Sa2YYfx0kGz9cQY+RLbWXdLXy8iQ9tNG3iJFSacLXJHA8ReC
92mdWZv6NeMdX/gN7f3DY5nyu65DXZGLcPYoNi/00sXoAP96zUe0GhoKxn2k
xuyVHQ8yAE9Ut7WOVauPBrzzxcMSfkeJis7nxFuuEO5acquO3uE/THaORPgf
fEV0vrplMMUbiTbx+STiEjRyJszoalP6cvKH1uLAtDSy4ji+uwQTfQ+9NZvj
FuMWo+EECtI4PzFL5P9q5sT2NphehmoDnfSUF1JlMiHnH89Uj66z4za8aOfC
GIKuTYKh8OPS0eyyTJQTDZfu/0HRLYu6MQbqUfGOvG+j4r6xQxlQUpcC+Kjy
D2lVrqyzccR/LsIVXqjGpmYsy6jS+IBz1k1/3dgZSHkP06HgPyls4Lv6mK+L
Bi0sXaK2Q2QDPQJkIRn2Mb5nITRTVBz+0ssFIuCpUhcH1NNTpIdqUAMqbwri
ZqyEyaQhB8V/Jtcuw3A+e8ruzDNWk1OzZa/Ryu5w2Gr1HJvX1bydkrxA/WJj
SEMI/VSDmBZeb/zD0S+VciGghO4pTmVBlffZ0XeBxSCYFv2O+0UzUgH16jMD
SW/9qLTN2PeFkb5510Xtcwy8kkQh53K0oBRB8bZrXApk5TneQ0Zx6pyuTws+
crY8AfYW2CBg2n2AyTzEIcZrv0RFCgn5/m0BrRJsxTKPRgtjW62JZxdvqU0B
KG5WwE8NIBWgFA0gjm+BJC6M/pF1fBEiafKJxa9KLRB9fJyScfOYiru0i8qs
jVyf69hZcHZYaGMLdhaklr0o84dI9jNoowOYE7QFInXFGH5pO/TCRsuil6aj
MEsZLuGYzjaz/f1TDf+DNJP44ezCqCou5pYPUbKrHvG1SOgNcJ4HKKUPJDaG
XIeEIhU1tiC354SlgF6MGE1CIlcIjei89d/DFgA2Z0BSefSxfP98lPZDUw0C
wQzx3pekVJ9SWEqa4zkmTIn3GnJbWNTCi0W96K2rkol/zd4PXGL7FOPwF/7O
5LfXNu0xmkfotqM2vA4SEX1tvipGsU5Vkw5EDXM27fL0LCKEesPzRddc5DVn
iKMlOvuhGI6NPl9s7OgnYuZW5O3vP/ORnbumNt32xhVMZsdAqdHMS8alzSUT
N/5lulOLadvTe0tT070vN+7bDYAAuLC4M3Gsw8QxqZiv7vJL7TAyPszCU0cu
Cl7subu1UsmYuBuHIz3okKwuWpci98kjUGTb0lc664T3QhCm/z4JD1jb+1wQ
N8BWHQMa/a8crmpJONGlsPrGQzFI0ywuMPNzkXfx2BuQAXFvDtPiMSMbaTLl
uM3sAeVYKmkTe78YHTZ40Tty2dOQrQT6T9/lwvO47vx+LQMyVS4jQxIHDP7t
JrSL0WXvsin6aKBg0hB6P0nxOfjZskDf9XzuUlSZL6hzYCwkG1ZS5dZhXIPq
z7SvexINHKXH6ZgdnOfKcmyarQwERENw693FPZehQE6zszWg7qzSMQ66bvLU
VBih4oTBF6joSh2Vsglt8oZD/TfUgXz8sLfgwqh9HW4cBPxqxTP5Y2V6YQDe
SEDVt2c8ETsD/NllLe7LtglntHojEkH1xkvmjJPnDgzBvSJK4lr6RrjrFYak
onnfEyvgTM8eqMgpkCFDyfWqiGjXJ3pEc0uVGtro+na7e7Xls+mfFqmEWF8U
G3+3MaUe7n7RiOf/+7SUZzpKrPHygTThqUDbLLN3+AnDbmA8du+lhb0NkYz+
mnRVbEio4OZSGdSYD/8bHoaCd556zPZNg4360lRTI6iFz0aVAeUATviG4mw5
DN7/vRQZDY476whMrMkiBk/oxI7hS8IhukCQwUHoJuRxxuDLKRzHq2pb4OdE
jqUIAIoGVXgCx/GpeZ+ehUhRqvq+P8TZFQD6SpBqxTjf3ftBgoxC1WdsqAq6
REe29EpNBVB41z8CxY+Nd8bHACHsVvn1jHifJRWn4mjwCZYRFCqrkcMHEqut
pbEcyTuQhARVnExyxJuaSLKc1wmnv3X8ZFb51CR85OLZI92T9GD+9Pbiktf+
AJiyyWv1xHFP+wAnXPAaIhJ7CK13dNQmk898DCcqLJ0gOz1qO4oG7R/yUA/D
ogCTbuwE6BmTgAVdIxh701zFJ8sD1GIt3RUw7Pk7XLe3N4fjo3snoyavGcZT
ddmgF0jns86HKVScmXdpBIBPd8TOXH9xM4rlRau9rrUZJHxXa3z7Wz0/JKaH
YHWFYxeIKO+a4zKN7tFG35UVwahnDEpw5cGuUm82XG0Y4bFYpFyX7id9XbKp
m9wUv0/pZj2UGR56QgbYB6nFAhUcWDAXzTKNpAJ22YIfN84iV+dMpBV9KX/y
BJ65+BE28wdcThb2+cWXdEgapGS/cgl8D66NmutfTUcd3VrB/tk1K7V8WZw9
75CODUeLaZYs8Ve9A3ksRu5PFmHPIYQEXjBhMtwsmS9cnHt+5wWLQ+/0tzUJ
QXRFJBSEsJwtg3vAnrI3K/m9bLQmAuvvTw0pI61pEAXsGyJqlfePaKPAoyTQ
/X0Sh6hpuitxn9+USOn7YjSYKTAFCeWD8MZGlierzEtRAXZzVxCu4ylEHUH8
l+pNe3KWHIg676yMKCE/0LadIVhjmnMIPyjSv/WPJNBsoKptEBMwOKtet8Az
wH8dAeMgwZyu4P0TiYTptSGZg+FnJS4BRUj5XmWVnvV45wgez2WI1YpGaBpp
y21U/oNNsEmIDonsY0A+Gpc33+wq1zZQrVq/Q+GnOHrHDHjcnCPlzNWgGQ4D
H2eohBQ8mV4Tjx6dXWgHYLeEoV8txCGlAMuqOx6tpru0w3E9Zr3LSWwJtGAA
zcq/27qrRLqB8lVEfGYiqG/rfFHnfYbZtti9YJ55W7XA0ZP2PuecGiQ+gTe+
I7Fs0umYI8LAm/VHsG33aip3G6mzvk75g6+96AuCJoIInDUmGCEG/zLZH8wu
PkCj0RwM0R4o+qJqkNcLX/kjZNr347c4PaWGYZ8R1EUPboABKokgG9qvSYR1
jRmMg35HnabfaxprUtpr1LKC13GnhNUtu/Jz2v0l3y3lAspvLl2gqhvv38NH
gQRt9Cs50MwKhtqVI+lV8retOralBUhH7VgikSDCYuVSCYFL156OX/Q3wMMg
ZF4fx6MWgnfUnXEzGKxTuWJcjTlm+Ctx64DAMvUjeC3uy0+o5T2FeKTDF6Hi
RlS2xHF9kSrc0iyyQ6jGKun/ZIxkZHYp2l0gNrlG6kuZO5taduSPBmAKhIF3
DTEUmMyHaQWEzauweYT/jP51DYWoxWbqoK2cExrKq/5LS5MjIpCs2Iq5NJ1H
GNYEdLL8yU54cQzz5dMJ9QkndDQle+i4mn3/y+tacHnumr0w9Of+FvDdluEg
MRIZclElj9L3hp1lV7Ynt39zI/UewDW7RvwDNjPIwyPhZohL0ZzpBEd+du55
F+7xff3ttil/n9C5hDqEDYOpqOa52//Ds+2Z0QH9Cdu9B5CpsLTtvDVEOTq2
GS2QQ/8oC3Xa82lD3LLa9N2+6DqXrInsp3qM3figS8gOXiERcgFoODt9kcO/
RZxiuRXUo0+16lONFedhIm5JIQjIEDgPdeShzEXmDNk3LNDl+dMZmIOA8kDw
kRan+SKuYMzmxQrU3ML29m5i78FCbRLQZgMrT6MWi+41d/l3o/c+u851qj3O
XijxNzZZf2LmhRjnnzbBPtLH/kyEGQCKA5qbyEbLAsX1UkDzCDoIlj2Eyzyz
6w/llQGbnOCCDSMOzcd0Bus36m1URpH8lsLTlTlLAIAOL/KUU0oK0I4wCMvR
LU4X9v3qT1IPU9Q70vw1mQmYwrr3lYKIn9QYb+PYJPq5dfSQxrIoltOeJy+J
e+DE3YoJuU85+AaKHrXW+rsNIggVA/fSyy+0wholFuwvFcGekFg0NNgutAsU
HmQ/EZxWHteMoc0u+fOGaMi+U74SAoQOpq8kX4jIM+O6vff4FxK2nRzEduDN
GBnsfZr7ReigBZ8lCmaOyazSPP73dDMIolmry333AtdF7teK1a2UdSbLPH2Y
P4UnN9NfZP3fghyWAktHF9WP5aoGKTcgRuhvNsdytHiJauE+OZjljPLkHSgk
YcrxvWE9CsXKvL5WMX8a+xY7QpheNopHigpR3lIYA1CMN4IaqVswD5DqzzjF
nrG6qkUXls7F6UioAAkkzWUT5RLSOvSlNDfQvN09LOtaIphnDLbse5Ede0AB
HCooCGsOIjLmg0u9upWK7PRKZNLqKWbvLhPiUvnBa3tJtMfmMSp1xtwx7HwV
1DBkzGN2SRRTY1OjVlKfYvMMVcF8y8v+4vnDh5NkykPTAYtuzdFtE1WV3vx/
TYrKpg1ZTNlJHpcIuHEZvvQg7pWZ7QIHeuxKfQiOqe27FJTmAwhojGZ+g/+a
6Vg5Rkvdi+Z1R6jI3bl2akUW/hOZ4tx6UqM4B/3I7zODy/EWZdAy2monIaLX
AphNd4PeYN7Z5P8uzuaTqUgAaJ+V/n860GZd3YZaRUnIH0U+uebya1rgSD/z
aFnf2ke3bVz89AF9KNJ2gi44ZYGRzYaIpch+9D0AKufOEEMjmzpra+tALY2z
2WT8ELoT+MyG/S5ZZDL9Xt59ADQueaXFHGHOpArxGnu6Xnjf0jFgdunep6y/
n2wgCI7kwT6+hvGvFQPNZ7KgcMIqU4p/PFGl1m5OpQAZ+eHbQuQz5Cfbj5F+
idMsG8qeDOZ7wAUkSgdy7LIWqOCRU75XIU//WsXTtegFMQMxYibnhfON3rw1
R2UaFWt/pwpWQiVf2231shsWlloqjLoOFr+nMm9AsYctIGE+/tGk7Wb8au4O
FoCZiWaeq7IldYkE3CLXBUSnOfLmT00kyrTH+ovDFa772c4OtWAfmvTfsn/D
Z7vZw2ymG81b3WmhOLbXhZXghfco9S38AARLTLeRrU+bDBeB2TnwKm6MLbTl
Qxvrr71aKV9DjIpUVX31EG1zbKWjo9Fj+mVCmNj2oSu+iBcb5Y6ZLvZScsgN
fZkm8LRpDt5W6jy/tTMm8rDGtIYfrZeXhRmdv7BIXuWZ73o0mmWIq8CO/I+u
dmkSk7rVwzr50fWBirGGnTHV5KNCk1MAvBZHwi0PUIugJFVoVhOZo7nnXY32
AUd20TmgyMTOkTPXfncArNtYEyIYNukoX/RInTHClkDK6RfSPsG4FK4jl9+m
IZhzBExbIyxdqBKDV+BVMHlggzQ+sEYwuagWT553i9pn+WBJTTTwPBn8fLb5
AkXkwMyQRzS0at97OPcJiMOJOWTjDoNmzc00GZZv/mP3jLYe1zhRY8309oTM
G/iVnL5JlbmRQSfkDu3rrfJAY3TI3q4YOLNlIwBQj4iQWg2sjXqVAnLe2+PG
2+JI+hZccCHpTouxoxKgpdLD79u1eatNQZbkQSPFGDOZpnI2Ql9uWQWEuIpu
BOPUzQXtSwrlL6hyz3tfXBRok4tQxCKs6Shj8QVTh8PiKQL5hdEsLWW8HwfG
zv1TwGlrJrHpXUcqz9czil3nxsEOvVlQq/jDVYyhuohk58aj+/ts1qab198T
g7U87rZICAgTbMD1ISaN5w2O9XEdGlXeNDiRUZBVFm+a6Ku2FDKpP7dB1opo
E0b2v35a1KogVuA2atEhp0ariDWPZwjjwmBCX8mqbc/WQFvbOdkX6Uj//8d2
CPXbloAp/3upxq5+EO1FwRprjFGNrBeYZYmWeLO/1pnPHwqyOSMPUYK2PFT1
oRnVxZPnI00so7PKstcXTlnxwoq8Zkn0Udpy1owYsLpFCUtUGGaLNfE6P+zl
F2waELglcJ1Y0RHdL0SH6wOJPLC6tYkxEGq5CNLn52XNkVbuTzEbJMQhY7YN
6+N47EXswkmRXAE7+HA/qu4XOm30PubGHDPMpyvngJhS3MwdJFXitufxkt0j
vv7Unwh0lKmQqDrV2ElC4Ui1aj+Vf+9gY3rWnTZIffc1MVC8j8D9k21xW9k8
OwMdCiCIOukLbJMpFhvY4lqO5rqNxJtuBErh08LewHOhtBxqawqzx/xnpvKI
hJAHHeONYvngdGYNncqSHZ7rgBeUkTnEKqhT9w+sH9J778Scq4Ev7k+WvjBg
MZCvkIoArZHD3R/e9Zy2wdQaFR6nJkSr9SO51NsXSy4I/YcvbyQAPyi0FHzz
7PctxPIYcbRTbjDLmNRs7y3/2391rfCsvHcTpSlwweR9Yc02YlFOEK+VTBoS
eu2YBjVbgI3faSzogmZwZwTcxoNIfWkwRWC7H9aFw50ogJtXHuSvYojaak3z
TZBq3OF4z+GBKnSMWFZYQ6TP2IZazL/wE1eXZBzl+Cg7EIvvJs35oH9KKd6v
SUg1JXqAe1GhcDl625Do7xFGOh9+ID4vBC+MChxh2K1hyU78Z6V9B/QFN+vl
W3kQlRPyWXR3RaPa65CD41Vwtqb7JOVRoFuL8ugAOyQaon+oLexme1fIUEJo
z2tKm+43tjHkQq+QfDSD4Db4agnoHy1ovO2mfGFy6J0kUV4q3/tZAVo2Hlfr
+q6r40T2cY1pQMvZW/JgLNMaxfTjbbnJAqHAuoTgcKvHXP5Tyciu3jGDcpzc
wV/kNGmGjJMGHeuFDidBiPpUoyz6qFE8FrQ0Gl7yhEGIynuu6QO39Ih9NNhx
yiCkZukphvXolXKIl6lad/vSO7/FgwVmxy7O0hzrFJPz3B8SRYKNZ4xOaGYq
r14dWQZmxlFaVvP/EmkhqVWPkwJPmBlNrPQmdXKLRclUScA2iILu0itfkaTc
xkD2M2PdqrGa67E93dLJE1f7vQb1Id/M5n3FRV7yfXLcuj1moJI91+gtRuxQ
HQd/tiro+ZUgTXKMVBqKIFSKwDcP+/Cyquqb7YxDfRuzw3FMuKX4mmPkTR/o
mMt7S0rO3d2osCbjnoWKwODz4sW+WeYdCwpQdRxFN9ylkj/rN13PxiMtmsno
W37u/JSoeXCyoT9etZoR8yDw76jfONxUbv37QW6Xjcm/YmIDAmT+qftdUWGQ
5tIwxYpBeygqKbIW7yZ84OOqFr7x0csdWLOGlfK2xYr8GowNJ1WU1faRpIY8
1jNP8eQ8BtosU7rUMWgNxnYfRUlEnu8mgrizZ/qSOJVPgf5+R5Jsj1Z/+yBk
DaAJZURN4XDjP4Jak5AQEGhae7ikF5wTBp0McG4GAnZ14V/ELAaRC2j6i94p
fEMQdEXxTG3pRj0chKVaxpQKBZWBmBBXlgFPjwCH8tFTsq842w7PY4gSYqtS
cAGdwSI3aPnVOuMJ/rnX7iVTEQUu4/Edu32JXdJMjdiITq2KkgR1dn0s/fg+
bhaXAGLRPu4RzrlyB8Q2cw+X9TmJ+JRppticzhK4LU34f6PdQZRm9CxWJfjx
YJxhu9jtzS00+RMiKUdZYlcLMvosQkMTmdQ/aRhutYxH/Zw3f5T2A4XMcnq+
zq43ID+Uvtl+dBaBH3++k1RLkpBMJs3RRq+IoVD1ZCGZmnFJBS02mYgmCl0v
K+FpG/sRzAmuHOSCMtFP1O5U+Y9KbugzJ3TbTcnIGJCGblOQ3Ab8My9OnNbw
HjDgntIQLdMLhx/D9YE++ejB4ggnpYobgJ1gNZh4z0hn6y6Um8FvPEsSmS0x
guvRfCLW4pmaymLsFvqJ5zptM56Qd9p4FtPq5Id5pYz6f8fXM9AyaiJ8C95O
YQRhmxRJWItNjMwzuIZBQDiwl35XtQUuqjEDYBly/KTnZ467LFaFxk5q0U0E
8ncxcZusIMlEz7ffOOdxpKJG91YjSAY32BkTun1P0OqfkQzBGnxQAPpyT9X3
YrOZSklUBputPyRJ4v77dqHRIJ5urrsAANtNDtunCWmFKYteS916nKvrJ5LL
9MBnTwQf6Mit7RPc6cXqYX75NGzZoxZlbrt0nuoKb+kRGJWl1CUu+SHerV9n
Poqd2xRg004M4PvMGCXr/BPSyT7G3J368QZH8JUmV1qtOmRrcZ6eAIPxLLWV
QqrxOrRn2ebdzBjWrPAy64KRUyaWu5EBSs05sCGwqZS7LXosbdcUCfimrygF
STepFjl6POV8WUk0Fqw7KYltvaPttuqRlb4v5YvXCWOQD7vvtibdANRUi9b2
VLuMMuF3LnUfv+QkDiVodltNt6M//Z42Kmsauy+GxQQNiWcqiooMkdvjD0GP
+AphDFVrn1kZxhqlUASHCBj00guryyR+khFFCFOt8LkbZu2Ju0VbetYKjTeC
MpucB4eMHUFdRyN+QUDCrvinLaDuvzY0EqLhXVwlzsDvs2uTT/CuPazRwfK+
HMTYYzFgHV7Z6O7U2EvQ5ZkWpkHc02TbEvLpMGebcRePmHMRYQ0SxwMS5R+r
dKJuY+EMl/iK8GYvspDOOw+fcsAd9pVQSboRt4EF4hAYROnHyg6DW1LVlpg9
/HKxyCR/MH76gPXAYhS4pY2Rc/ZGyGHOg15q1bbTvbxqUr/iZQ1JQJdOya1c
VQL5s7ruNsr/mtPhXB3/MlYxOGoJ5QnigQ+7bjtwEgWe53z8CSiTudHpVs2I
l3tax5Qh9vidLExTCJ2nYbz1i1nx5LGTZ0mpFQVSkvatJJmnAkU2lcL+ijCT
sd4eG6iOuqWjYeK2HUBEkdIVFx7aiPp8uVRPocKVB3zTJw9eXi3/egTjguG2
93VSXdz0lmyxhBVerI3GEnj37z3IfdCATDjtU4lmcTaVhxFOz4EGGs6MxRHQ
W0pINqa2G2XTaONYWZKSb4BvU5CfD5CNJLksyUS8Fw8X54xS1vyWT1e98vyG
Tx5lxWQB/BUrsBGGh7rt+LshBfW92c+Srdav+gVUc4YBLUCJ50tamcCoHj96
Qkv/8AFyGBuSLhCsTfRyERYpIVmvPxXtCh3+B2PPfMShSxvWgoUMdQvr+W01
2G2ZUZcf4afDPox93OmxCl7SkyVXQTG3yUQVcR2pXrLMXgHysb73/fx5cLpn
VgIVtJN98WNaTlPYdm4uvfduB+iqJS2+wW7oIU1RSZmxO1BudthUpQASUPro
1zhW+ByjO2UBiKDjbnc0ObixzMb/4AlOerwiAhM+4n69/yXhFVwP6bkZ1Vkg
/RNjIi5TqJ4YEm3nGFYK0D7lZGZwmtP/xRi9LRYoWHKzcuNJ/VVxWFW1lzeL
bZ8oDyjtBkS5KnAm6DATFYEdDWWBeJXtYihfylzXxevGWMfjj4zSXk25Ei2y
NJFIC5eSroDT8cVTCOqooI5e0PaFjgLMbesZjnjoHjSKsxicdGUbn+DK+bEc
v6EIm/YJvOgvBOQzuGf1QvAwIsEpPbjnvzzU3Cubxy4RYwQ9zpwkZd9yuxAD
aI79urcYQTTaNsjRkVImjTr0jzEXcNhIJiUHoVW04wxgWbHZLpl8mYg/B1st
8j/XBbvjThkFHVlC6h2ZaVe5l8j+V42p30XcuqTklesgHZhqc4ppm48h5GGo
yLOwhNW4rMsDhvRL/muVV/EfheDfaOTgsSkRqCUOfOMWk7TA0815c1r5gFfd
9SeV1STr0sYVsHyvwW83KPzqwR7N2t1m/I8S+YlZ0A1x+Du9V1XFQMgF1wSH
s0LmPw6KW/Ryc6204dyVO3/iQZC5fc+B0z54PKl7kziavreZh6hwOXubmeqi
+9aMVkqs45Mv849gkqtHt0qe14PKs+wwxigFjvvFWKXWUZOrp07lE3hXb4d3
lpbjXS7ovc91IwJiE2YwOgkA5e5VZA0xzgU24ofqOVdaedunSrsBeRlFkBMo
WETZS9/KPswBfhFYt7lnkjaCUZtlalX4EX72gb1fGyiNWp4A8GDWUDcD9ng4
zqLAjZDCIMzWVxsdpiU08WxGjFDG2nFqIYCf+pSb5KD+ikJrmm62bl5qyLR+
ctCK7E4VSiXJXSEnuBegwkTYT/Hl48B0jz8zstU0/NSbsxsOq2MEpWzwS7GS
lVgpDdSuaSmpqJT+LQrQpIgklr4tXuJ17UDN9wKuECQyNerhU2N+8NshRPLk
3HZJlXXoKbtTJkE7Vt8lKWNBmJPQ+wG/SUuugRL2ewHbvjwgFGlEprZzkfyt
LvN77yo6iYky9NK4M2m6y/0gcdAcl0XtDgIhncvpWm90j9Mc7YSgYp9/q3F4
gYn5IQbZGLkF0db7EmrZhAXSpAU/q4IXl3IKjIVIb2ElavDug6E3jSQHbIEb
Pr3zY6aj6Yd3K4eAGWzmrs3HAAyXckvfu8R9IYCWw/BpYLDZrj5DR85F56KL
xMxatVvurkiajATYqzQJAuH1yG9khN8mG+AIZbMLI6TSDH8fDF94gvnM1lSk
CkS9NsdqSKigLf41b2w2orIAD//PTecpv9eYIBUBcOY/ljM9CHVxHoMAukwc
7N2nwa9VL102wVDdK5vyTtt0c4ca/uXqBx3CB8567iiet62sz2INM2x3Vk1P
aiS2jwYM69gN1IaAyWUUWoYsQA6qs6cCWArQ+HUUuG1iHaRqN5cSnCWMK1tV
P8/BR1ybOwUu6oxen2M6QZFSVJ1UBP/05jGs623Q0fFALvqHBybMJkOEDcRz
rlif+4hd8z83JuTsm53IvQmp5DLXFM1Mz8Non7PdA92HsWqEslrvAxPoXWsC
GaZHqS3HtDuiR5E+SON4EeDI4woA/lLF3rTBsWNrsQBDbZNYolkvbIQXZZp3
wiq5YPz5/hu/LU3bSEZKaRKCwHT6uhcC9hhgBS17FvkKxyP7iarweEMZ5gpK
UzyB4SN2pOTS26Lf667ZGzCRBipHtHGfLQh2J/xQEaS+Qk4o/PeY09hKSAum
nMZCZ7oTw81UIt172SO9LNXo5IxEZUVY+d4xdJSDW6J5Kqa2zmm5selxrh05
PeeAAk7JJahOtUuN3UFxF9ZpCsJfktdiyTbiienWVP40k889HIEah9SrmlLT
RRjAMBkDd3SDw619j6U9rqbWxYrGreZ5cUgVpLH8U/IrAeLCoOg4AeLyuzY0
xo4Er1RE6Bic0zg8D/Inzv2LIpSSqZpR947+TzCcM9OAmruFyywx25R1jjwv
TtgnJaxolD5jCLXrYC7t67VTk/W7ccBgjs2lS+42e7IH5PJPhhmvpMBwDSOT
c290EEdQ/vSfZiRG8A2rdSXZHqhqknN8Gj8ddDAadccMsdEFYVqm2Qt4bN4G
yo5g86t2sLyb5LX1UC3bkJAjl1OBfc0i8eRAA34C8wRdgRcuqldHWpbo5eOe
8A8OANY6XaQaQjKSsmurklGfzcppOLsmQ0QO0R1xsWb5RB7Y1EiUDQkntkHj
Z7MGmG8AFM4C1KCHU+YU5dTjzPMM0evDEiVywuc+5+dtMMZc0J2XudAN6lY1
GYPD+l8nSoctKCIzveKtYECs1/aa8Gboj1BuX83JGzqpuTwcpP3qv1+uXO1v
pKQeUEqLTBPnNr2W/yEzW1S7wYMfuucMoWxJDBQNupS0ZsN+I06dgjM1NdHM
OkGEY9V4iOVUyCoR/PzOQXsnYPg/J6BNwG1207GIGZFQ9ESI4q4fTz8imC35
iH5yf3zwvhXXu7DRDR4kQHjSr7OC5dXuT4uF6t4fqH0p7JS/X/702ItoHgon
nKmshzuPW9eGDRsrYR46ivfQyccR6leSUUWWfzjxWhgVvYE0fYWOXRnL6Iek
rdD6bGKSrhF7TF1wvhO6ZhamNKXxVV2njoGxd8HAaXzaVBnREMm3niiTZCxt
jmTWFymhIB7Zi6RzbjfGSf6I7bg2A7+htIp735MlHLDVWTFUo9m9nPFlCKaC
g1r95HkkBqQsr2cVLm7SN7XpQT9UsipnPFT32Clf4WS79fkYiTBHnX2qa5qh
NY2vg9yCtIzoXPIwkHJbo2A/KnlJ3IjcEH0Ui9bNR//Tz9zPG53TFZzlRQSc
IEVGwDSSF0C+ODhZ88eo4Q4rWGxp8ucjiEpgmIT6CGp6pcrhKz/QFNTv+IWF
049DtwYSW73gnd0ufgnTi0HzhkVYOM+9m0Dunit+vTPpablSRlUZL3aYj3Av
2pPvsUIBg5XCJ7ivPEB+8Jwx57lXSt26Z5SPOC9hQzLXz7w7WdY9B1ArC9XF
OaynYOpvss7uHSxgCZyqDgSKfAaV71bV57Jl3PM/bzqw5eNrZL4cRwZBg0qJ
nrEo4swPlcTaZlI++vXcZuf9I9CHC2dIfs4FzjiL54L3NeAcVZNSvtcvncm7
kRo/k1w6K970ts2ZZUHdBFnXRdno8NGZf23nxdMF/UtHWrnOKNtbRQELcbzo
D9ncO+XhPEFRzAt0oC10wSIBIDDJ1hecCaV7DPiu2MdXEQfYDtL2DRznmemi
3P+xbOrY5u0srC9UBN9OFpxkJeiT86TGu0VsHfm2uyiXUBtdbtvPIOKAPQ9k
EHRTWVBNKbJk718frqZugeeIH83zYAp8+tPfr0gobWJ9W9Ofg/vHwxdfvkcd
Fvlnauta0uudQlKvm868u7o8LxDNZSGXnjrtR54cUHOKWdkOCaTVadXe1i7C
5ctOm1ES18Vs2MYIHQRA+OF048yJKc15CYY301jExpuFa3jCr0LwdUNdmFeK
7NHC9siTQpufsMwD9wzz8q5QmwkmzsENFFh8zbKPIIMvPTeoF8qvReQg7GFG
C6LPIbKo0vBveF/K1i2AQ/HJZCsOvJWL5Trz5BIBIpTIf38URDu6wbQe++Gm
ps7/a5xs5FW/+fkdNRK3CkK0UzPogdXsnnA4WpLDeh7JFjGXzVCHHmoCeBN0
bFQwGHX4gFaCp1E0renAWmhw1fF7Iswn2JBtLrQBwZgTccR0tg+eldhUv5aW
5+kFapWyz7RkQAumu5Jjqp1I/Rcf+5KP/rvhWiC5y4JbG40CIkd9tK6AEyuI
kZMLKPC2CKpyiyovGIQvPSDm+OTYmzaHJkda0fSejow5UzWltInEwNRD4ulr
ogae2yw5bCMK4tu/tZQl1vKq3WL/PXMeepobIOhg9jV4wDOJN9fohiu/bthk
PNhNx1pjdHIf938/VNaiGbolVUTX64uk8pQQriRxeGBSql3mvAlSFKmkBoQg
izThj3va6NjzAOy6WviUhPO7fEUP4R5+esU18iPJNzLiqTSrTkKMlFm690mW
7utpmjRTHHkvkhNYutyKMIc3b88MOi1MHyo3E8XXrJzZuFyk8BOVnHZ0GiEl
b5OqNY4i8+RSB9/rm3QZc3ibQo8fifno14T2b0u7u00jI+WQmmpeJgA89MJa
mzwUambTBgKIlEDwDJqDqgEIcpTHGBGNimVoUrD8kBtqA92ynTrxwXpVH3PA
N8DLR9uLFxzh72voISjN8H4/Yd51Boyh6htA5Qg5PbBldnt7FELFgXJASj45
Ca1k38pHOPtl6pEkFx5oZeLw70Y38rxfUz2BQU/JjZWZzowt+0gRNzJSfRs7
07M/nnPUj81YwuxBdDQJiaCaYbOjWHxotjI3O8DLeAVGw2rCMFS18fo4coZn
1rnzq4dARb+6e8gUyrOsVlTFTgDWZtRK3nAbB9sC5lkq4Z5a9arJxZu+warz
O8FJU4dP0sqHJKGBU4H6sc0Jsq31cpw04QrlvDujwcub8sIvHZ+EM/Le3hTj
b+6wqYNm3yN4zo8fyWgh+00+G1dfB8OhYGLiO0CQEtk6E3uRuPc8PDYFYQVg
UkmomAu5ypHZSx402ZhnzXVIH1q3jkfyBRt9AjASJKi4rFYxhO1lciahAnH9
xxvMlrklDlvGbM5pW1O0WJHByD4fKf17bH2Ip2Gu1OWhwtuNszG7m+C3IZr8
59IIFDhLCHDU9Os3flOacOjN4GnVYemjHIOaZZolnkzwLtNY3a75TJVzty/G
l1xs1B9BXvpcfU/4YfL2h9ihYmEMltRAUGPZkGQUrbJN2KCD/iICfp66bEoP
1ax00eWkMrSKHWtsUYqDew1v2Wux4CaWaRvZPdoZyGmulO9gpVLPXw7BmpzE
wx6C8k++8DvrGUnhAGJBC7yeiuGC8FTDQNR/0Rj4rLVg3YxK1KB2zTwN0e9r
TrC5OKafCLYl5bXCtTfw4C4X9BL4Sp8ZfWSdlgARqoACKUIENY6FZxggWgK0
7xBA7K29zlD9rWrJ16KW6RGWaTF6c5r84OHyYwXsqPdve+6o5O0u/yBH46Ey
P7HFlXyb1R/4bfeE9n9hXJ1hvvvb/3sVvvYKNW4xLHgJVuFFFJOu+DIzZ7SG
jeZWpT4GOpaA6iHlAbiENWKyyzyW8dCf8GcBht04CdokHVaqkC94CYoQg9zi
PGyVjyVZpCSFeLChb0/g8BR3lbxDh6jvZF5pG0Kt+8ku39zCDH/4hY6yBGal
MLju9JAxOhAFNFamh1u0Cv7zpi/XVVwFugPHz7Dz6ifDwhY3kfuHulo/Q5dC
L1lvBqOf0tjoog2ZjI7YbYhlpwQA9GwIACmAU3mowRSooleweFi16sHp/c1D
enfu134wQBhLj8N8kMIhUdgSzEON0CLQ/OAficgGi81sLd53rVxBG9y/bp9i
vZZ7+jHo5vpPOQCVt96poNWKkc/5q9s42jY+argOhUBXIK1fsAGQ1Xh18eSb
pRrYAHRSl/B1w2lz1sFZiaKMOArzgSgC/JWRtqctJZDhyYgVGUkHa2Gt22l+
3hnTLos04tGl1hIuIEr8kGB0MaJaDa96aKBJWBaNeZQy/Kl7Q01/xB4aT0W6
Fwkud6qDMFREsdwQtvIc32pLAWJZkGD1rEj9RjfktVk9nyq6IcJbS5ryM9aR
udTCmlebM4ukNKX9NJ+p6j7npfDx3XGxkpsoACNXIfxVthr+SSnPgzUQoxq1
dXtVKEKkPVt5+80oTs8ZMfOkmMggvoeh8YJOFh1HiOMOZe3xntn1j3vPZb44
x6clAM+VWwNbMSAYpx269nmt4R4jjXZDpEaLCJto3Mz8OrVMWtXAMYcwU70l
X87ZzEGcMFp6+p8v7IdUqE58/4OTrg/7BQA/dq9+sCmMIn/sDQk2OFyo/KVX
8+di4hHlHttt3CT6fyzu1Gee2rFHM6fUJpN/d/tyxZrNEDJK5HeAGWL7T/Sf
WIKBkGKyy6RA0qH7iIPkjkOwuEw8q3KDOZrtEQ0rW6sGtnccp8mTZJGukzeI
bgsiAJqBbCu0uKenaKyAsl2du7S43DfqjYAchcRGJwTMRKbCc/FsNMp7OqLv
uYXWB5ZrVdoP7ZHl4n+7P5Fg5oYWYUNJskNgQe6h1nk0HuIpOdweNJYoy7ry
fWLBZw5wuJqH/4s1wjeBj617++kWkILxsT+IYNnfyk9QExM9BcUBfmCFMMA0
War4o5fpqu1mMZ+PBVhDaYyGLOlXeXhr6MRRSlMjIjhRLTTC48DdMXLB2lj+
T9RO5bG5AZ7E51G7wbYeYre2pGSgfMtnQ9ebSrzFWi6NHA17FlRVx9Xymf5C
tvw2Y4bNfrHdsT2EphCwvppv2UsZWzgWayyptxnaeN9PIEDAshHP80+OeUh2
leakRDOfOi/BsTdOmozbQlsbydaEOuE+bNr3coWKVDB4XVk9yXFpxmWjF8JG
AgC+6p3W9RJPm2cZwzS0dDUU/StNmANsDvdqSSpMRQikqULDwpVd9YcSaXgs
4Loi8I0Zdd+fO7tqGq9IXbnwF1FrTtUMi6Lvob3E7RWQj1zL1ourPDDayUrs
k9hMhfQQCaYFaCKZbmJBFO9NUsTL5ZWrETLqkyRhV/P/KWT2HNiGLVeUmbkk
XE7INd2NRViCd0I+sDObcqbfsFXQEdaPK9bMbT2YbB8U5SVd6HeJ0ULX+okd
3xWHKqdXMH9qVtPNSd5+kqgUgsS749wXrDPOc88Zn162Er64mOlRuPbsCyST
mbEAyzaR+8lyiDnxeWJMb/XPWByIx389mXETv9awHg+2+nwtNmmjAKounTU7
4Ow4Ya/JMdULFZDJzzIqB2dQYFdacqZuXGxtVHCogZLTDtTuqLRNhOKQW/sb
t+K3ukEfKOvCoxWYlqv3NLOZOkZwb9E4oJBswjkQwrFpamms8h/DIzy7mXWZ
it2QcMhlYCI07cGr25VJgbYw7Imr7WkpDakwbu/pywH+SJ229B8+fNkpntzE
BUXu25bnaTzNiZX0ady0OGmMNJbgAFunxhUdDigpRYf0IrfG8CQES9pQnr/8
uL5ZXeJZbGkFh+UAACqv7qnNF57jcQOASdnjWjEaluFbsZr8D0AhcdZoXkaE
4WKi1qjLwBAFbqi0R0e0XbdFlvXiJ6tbZyFvGatbH/4LGlaQ+jdst35m/rig
GsDo+sAeBbRiuMeQ8LkUx58W64S2yoxai3aOxziSc3SpF5sO+Wo0YlP2kknl
mUIQjjvDIiFANwi8eGQexAJbhLnX1xBD9G8lc00fbICnBoYCgiwkEArz2nnD
Q46ql9CoorPia4pS98l3eTTAOC1sPHD6WLo0qfHt55KmX5TNcKqLhvQ/jgca
b/Nr0ZhCnn2D6LM6I23OLRBA4VL3KhKDSYBucuqaf5wT2VBTyd90uzvxnjP9
kkCv3I90v6fTjmv8SOw01R6V/rYXChYesq3BweBs8VS+AXN5oek71eou+zRw
BuftLy+Qp6G4ov7ujor5YyRBNmaDhBxTydFQGemC62f7h/EzU4z0v1pcnMaf
Isvk4X13w7ov2GUxZ1LiBLLdj/yf5/sM8FgHYr8Jjn6v1GsdtU66DWZh6l/r
DcupATd2KiyM5+yQ9Rb3BDEimE/DQQLX6WfZIuzdgaQG27cHWlvzySzGlZdZ
AAkdjLu+2Bpjqv0caTWi8sBgTcqHC66wX/j+nCy3kVK8r9ciV47UJPQ8QZv7
q+3Aoc+jUrIxgjLSn/TuB/K1wtCQPkThB2bD+Z/i3/kkw/Vws/myQUEHQdFu
EhcsxaKZLwGRY0onA/XL6YgghaX0BUsEfwwjNpP4SY61ekWK7/EeI044EWNZ
n6pYC51b+ns9nvHgR4kN0OhQt6PYjpJqFC4vo1tsoR8mYukJlYqQnQRjX/Ip
STsimLu/UeGNXw4lpFWOniqMTTzQjcy0lAL2zXKdCNypyxP3iY23qml3KTXL
GFdTaxNk04i01mgyuWGwIPrvfCuPV5Rx5fDfh2v+EqBhwojwSiT8i5QcfyU4
y1Bl262/xfCeNWbVnFRby1kbbO+q3zM9JGCyTN8VSjaGCAnAyHmH1gtj4GK/
7En/E7E/TX4Muy6OIwub5NL7O1g6+F2fD8pOk72aazg3p0kISdFylz2kmkym
Qn7C115kSnlpaI0uZcoN26V4HPEk78OSKWXX2Kg9wUYE6JhWZeWDFrWFfTeu
RxXB0rxEP0SiOTXafJ3BQpMO53MtIKX7DpBqQekUkc63YJeq3mMiLNpV+yVF
VniuhNuzpJ5nMJIL0RlU6FHXYS3JCKrNpfTcta3bUvWIbK0x1Aa4bMh9rVtG
t0YyvSlDh2r2gRBGahMXXOe5FQs7FhnsGVOy1pHUHgzQlp0l2yDZVcgMRg7f
BMHR3Wy0ZiskBKTzfrZPE7uX4FN4zHJThCiHc6jM+HYRjmepHucdevmJQVPE
X4dy8DdfHIkC40Be8DaC8mgMmH8Ex0hGWgVzhl3hedu36fTGPRhXV6/dhojs
Rtgl7cbtLe3ysJfwF7d49c53Kp59vgzGzJXozdGP66CrDnVNLgT5YGuuGjrW
ElaEbRhKzSvLLOzqS/WGUZva53uBHTX34psa9ccLT7YvA7dHD3buBj2mAMuS
ODC4b+goAOGIK6yaSCpGJcYtrV0nSg5Ah1DMjChYgTzCP9mnQPqpXnTZoOaH
pyXYTotpwM2pVhlSb95/1/yGNowPuIIUDLKmSG9RR/8QF2wCP4JdGEjRKKGn
uTsrJ4UtfQmJEW3SkfSGbOeyP7JJmPTe5ocylotDIU6bZjofvy05891rc+SV
BiIr9j7tW5DEt91Qr4NXEuVasmFwEjZ15Sp3aDKEQpGGQvMdAn7AHKXcGTxv
JOnNmlkorbKyQGXY/49cyr0eDLT91qUhdkcXY8Ut63VYTnZnXbzx7YrzXCwF
ptcOSx3l+LXniDIzKdcPS3HFSewZv4fySFYhytLYO22BYlJljnYvDld8cZqk
SyLRR8gZa8PLcC+gLQPza/LGBRZyydvX8EO2vXknMVPojgnWp+3u3bSKS3+y
8zp2SRhyFH+cbkj1lCgjMbP6ZBvs70nKWGnVsJN1ajV0yMWE814fKQQn6fAG
RRlCkdJ+kW3/nm/G65dg8/MUJI5kcPS1uJlEf4ak47GSJAerz5pLRmGAe/oR
xXKh9lnFkwExo+Vsm2F425nVqShKUlTynmuGAH3FUajqlJjJL+HZ5+UZE4FO
UV32WSzjJJytr92Ligts12C6xZrM0RaM6RiwQXqUqVsMT+NIxkFvR0UELske
1a+8qZtHQe81YVfXGgiHBQfu9HEED9VESYnxKbFIa8Fw7hCBEOYVeArop4uD
DOLnrhJPlG9gc5og151JF+u6ZZP71c3HIO3vvVpGcCLFi8iDA0myWv8Fe/2n
qdExDUiMOugEFC0RZqtCc5hYm3gzgSNr/x+6MqlCE77dKBSkIhxj+IrF/5mo
oQxtASNSi2cA17wO/mx+MQtDWAc5JGFgXw8JXurQcEc0EOwyI36SZncHPVJq
LmcFmjXWP87zXofZghKf/2Xk3LvWyw3++tjE8IKxBJFNEZdzsVNoLRvr4by6
IW7snrEjOXUzHvM6xGDDOFqv6kPAedh8xqV3jE9mxLQgl4YL6Ppvltv4iZXP
31V/Z3EiIWCtKjeJM3p7JLEUiuGqEHnPep5wQ55QtBHEWYdOvVbxOh/EWpI9
9eHnqbb2nhvSQ7jJmol1/VONKslGu7H0kFZOSF8ES9avh6w5VR1FWxNbtPXC
5MEp+91xGP9onUr/DZORltVZ7ru1y+4yZBEj/ewYmT6R/QdPUbpN453NLiD+
SipXwpDrstXRGTw90ZEP76Oz10oqfROhAAT3LGLmw1K0FgstVC3Sh7GN6CnY
TDEe6ZWAKsyY8L/VIiCTeRG6q6ujwVZneISqOX57XFUOQxUdM2Acae3upDlZ
pCMrgbAhM03PeQhthsW76I0AXZBjt0DeAb51/TEvbHD0DxbQywL7ukiSoX/P
GK8IQOxwXlLUFtQHvg1ox78qd5wytu1oP5V4ZijjzBPmQBh4r4ysr8qgxYdK
A0rNHSnyobmeXS1pEfIZT4oXfFrFITPH5Bo3DR4k1Gbe2ZLpocEeN0XheHQV
0twbqPcrUrS8SdXFjAt+GENosxcjDOOi0hfvLsZdX06RZv+Gk0AH6G0GUFHK
0AZhjqln8RjitpycB4qYP69nM7cwV0yerBPj5NAuQEh1smGOw8KOBPSVPrxW
xe5mYk99hyoqr8aJsjK+jnRcGWnEXTlqvf8nTstB+90cUuf1NQR79jAVupBB
uDqxgrZiczrWnktdpdcpXNpM1883VNAmv+UBN2qe4APzjSjhM68bnbf8OIPd
8U7IMnjg6QvhEylJ0YmHt6owQbmzu8Yabb5ePDXopJR/B1I8Nz7/gthFnwNY
nvz3mbtGd6+A5ncXCJ6O4qpum+iSPPOZa0ks9CjoGvG3eycaDyyEwBooXOHa
bB2Hm/p1duvOXN2EDourMGr4lu6iWS5XVHvxFm9O334o4t8dppacx1L0SmLn
nee6Hg+jhh11b6v5ectzojyMmI5+7ZG5b6C0pUcckC2BWdffyuRq770otXmV
jOECUjO0sAmreyFKrpu2nTRm49qqRzemI2h32dXAjoTxETo0V0tnaUURKbFn
/qiYkMW7ixaJUvCnq7BYG6hyE5kyHV0VHZWKOP0ZV6bOl1r5CGNESI5K8Obn
X10kNghvT+AdYdAHTrvss9Gs4qoLsnCpXfutHVisKmeyOZn+DFlTXenigCXW
qjBxlYXSQ81ZZuuMKT320tGUierTWW5dk5AHpDf+b8xmgaWDhf7nZ7uGfOvz
2acQUxwtU4CJpZxKsXVDyxrg+VXhTEBKR46C0FVdSt/2+9fnCReZLP6LTttY
qHcFA5yrHITh+gFaIlW4k6KByTJv4b3NJrIjbUzvEivE1nYiR199VfK/AylB
h6XOeRsud4+/e80MJPzGWkiyLl1SFl1PcUBxhGnlu+FfSSa6w0EwQ4EMp6aK
YX5vQFpB+nbrVeiNv9nePS+BWR7LdiAt20uM/kIMPf9BHsGQyvMt0n4zkuTv
tza38gJhO919BHc52yoo6NNceV5c93NQZpC/8Sqb2ECLeUbaNQWkRJfC2L46
YF7x0/8niomwcgU7hCLDv7O9gByXGHAd9lCjclUehqgLkF4ch/RBBPU3ffjK
RphOAc3eFk8w468gUxJfi7qWec8pbWlFO+dNlk3NDD+ZkblNd+ODRrfTwurV
4nexgH7ZP5TQB9X9M4xbrthWjFatopHGsQXXStS+NlSxF+2hgRBKH+aBNJqX
1uJkv4b1peJWdhYDTs0THGzuXrsCgMcxfd5NqlbPW/4L+CI2tw+NGT8AmU1S
HMTaCNWVvhIuLuhpRCbPNwin2d9Uzy2Hj1FdGRihM0cXVIIQMQ0xzunNapxc
iJCBtvK9Nuh4NWXZ7CNoEuQhNJErAoxkfTMulzwWYgW41ifJmvXaau8+lg9G
1SbRSiM+IoQd60bYZpymzzdnuUaw/9cR81IRFQjUVps+ZCHaf9UZGIRmiwI5
zPNeMbm3QH+TjHCb8+9YZZN06zvt+op2TeOvhB0E39x/Ed4yemFtb+rs1IyE
uLj48SXIuykImbe9aoYw34yNLSTwLiurrQWdhE6+swO5guA4J+fnaiYis+fl
7qMvW5kL4jRbzC/YgTtNOCI1EqZdusYbuPk4qQc6BbMp+3LkNW+d0JueWD/E
HIp1OUilES2qtc2LR6sOPvkS75aFX/u/zICIcZ/Gx3dAJQ9kZ1m9UAwVXgcd
k5VsDwFlV2JTVT/uMprr5WHjX1beJ29HLAzdmHPettQ9w6KQhfI0ACykoBEL
hj+T+yW9ExQNZMUU0GSpcK3KokYi/UgnLfeHUn9SygkKPY5f6eWE4ZM+yTSI
MwB0rJ5gvEPg6jwUyDkuIyO1q3hkpiPW+Sg4kjpsp7+lu1XBn1VhCsKJmYym
xxE7dTgwDrD6k0bArPbxZTb/r+FAtQ5asn6MB2wn2mPcK3/EEH0sq6qTr5XF
OA2E3Bb893hPrm9BRMB/fICKfRAIaoRT2SFK2ub3x1bHDtyLQk9j/k4WeAXY
eJ5GdvbwszLHVPkxs0vW45kxMbiZtfVpdNBB6oYqwgzdL5LBTUWpMbGXKtM4
rNTrtvafaDIhlAEs3PU100diFkQA6lzWhf2eUgHkTH/ijjsb35BL4ClyG64Y
oPujcaEa5THfKEl6Q0sKjK/EFbFQnIZTe3JR1nZgbCVEOe4u8ppKpHLMpyl6
7kuLtAAvG31b55xmHfWp7w83LBqPYXEJEMbXaVYXs4/rswKLH8N8pumoR6lJ
430Q+JNJ9ExDiJEfoJfGU6puDZIiD+JTjCoC1Ya1wir9GnU/5vdL8XqtiSrc
GU3gWuF8yznNgXlAWSMVqyz62d3EbOteKJUf0/y7dxFTBUhvw9TR2WiHDlCL
btzzBOGohzxNPlF2wKzK8wjV1Gd7DK8hAfCHEaLCT4gDizSgR71kKK8uK56y
LiUTf2Kp8b78j3VXdC+u0fwTSKLUnMSoKZ+p0NgUUc80JOhqpnQMyTXdfrQT
rz296WsUW+SYCSyufRXF630a8w/CzNEcogCaKEAjKdV4g80D5GhPVr31jljP
fy7vrXdsI93mU6vT0kkiqLAl8Rkb3h9akOthDt+OwUhQ7z4bTjq6pr/8PmUV
vTRLgQjz2olF9BHHA9AfpZLX49PMxNVcjOOvZnKCks5+J6SrE1Fma9fcqpXZ
7JAi+3IG2Zyodrl1rcZbw1qr6PZwkcimtlZYH9YMJS8und6a1i+6E5GOXZbN
8KiNA9pAjZpWuZqs/IP7ekFyrDB85RxvYp1MVnFT2EAMh07T6pSUIEVbRqrL
yiljO8SxP8Q75HVb1XGL9Ec9ad6PcNshTxY+MgeTO3l4vnQop1FnV3z7lKmq
Pj8NMsTNuzhIKcdu+LBt+H6ulSiGuy1D1L4fHTN8w38Pj6jzi4Qsio5QMuNX
XzNWfVDrgP6eKKn0I7Y17uk+3p89bw4xE1+6Roxp0flyQM+97ge3TW9zgOpc
KbNYr22ccS23FPioJ4GKxSS4FWUZFANBZZh8jYNzC1ksjdB7s83HDYcEIu0q
6UGPWW6u1l/Vi0T8afnlpB7m9KXBGQq+F7NETTIbq2Vij5EjI18QOPj43D6R
Q1Pwxv3rZr5QF5L9qfUqPlsG1/hwfIGh+vXkwSRB3QlMi+CGwG/2MvqWHFl0
R3Yhj7qYhm/T/RrWWz3hjqfU7n8OVfIs5sylMPEGzq9bdAY3sTwNp+ByyCP+
juuUDVts4YHBCAY2pqRQu43Yd216dxK2bKPg3seA68ihDk48q5Q7VIbIkxmY
oR2MhOMa9luCGKxxDlfaIIgs5sIhtj8yr5K2FIpZcezUljLjrLADOmZdUGCa
dfsZlGPMhszDruFSda1M9nkWRLYa6Jsh7gkVBw4h3BwtmPiOfWvT+ocNyv+D
MSlTV+UtM5AC1177Uk164bX/QZvWBEGsAC6G81eYatvlc+t7dOo0XNaCqWfD
UBaWXtjaboAnssYqtrvmZZOb7JNUlpIbT9SUqHyCCk1xmNCFteb6Oa7j3TZk
QQ+vimrgjybFAVlskUCgwpLlj7AVbjA6/sPw9MH6rA9bUGBmIzsm7zYBsehl
CVQr0GO8Rgcvh47dn+E8W8X7baZLpMl6b4J9KTN9GFbTpxKZovNawtUr02Eo
nnzpHs8QYHHQBbP8AybkypWFs1nrtFKD2oHW733P1Kf2o0EQV2/HqKTZCSRC
RPgc1UQtyu28yT50TzB3nbha+1DD6tSB3gYJds6hgb2JvrwEXsRmfSRjW/+U
sWlXm16a5Yj9Qv2a3IhiN10CMNIfgtsOmtQ8QjP6/LtGd/QQadbx3GNQkJbo
VL91IciHFavqXpPlOkyuWltmN32cSvKHE4b3oI0rK1dsfznkh8YZ9OOnbulS
/RWsBSKOZ1SIdhpZmFkZhmE+JaA+BWo//L4xlSz/EcpuIGD5oH9+8dLo/EYg
VpYBtNTS64LSQcuZjiLTZVJ4f7zldZc/fcCJOzhzVFteu1gQQzV/6e1ZuWK+
Iy51LdfdXp70RBiXGRNETndkbgB4Fl5jvgnRRii0EmT4LHhOpLcrvCIq/gNg
6KgioVeL9RFEcxsmQFu/G0NI+hM0b4jH04qSscbJQUP5KYbA74javh0saH40
igXYqVVjHL8pQWXvBbsXjC4NodPn12pIqw+srJoe7L/eecODi/R+PqajaIhu
8/keHrHA+p06aBAQx657vgjNYOHDRxoh9AYrINMKH+t+eZaaikMWB/uFcg8M
bqveLhGVn4BTZLPgVf27FxlAKefPzYWgEuje9S8Y8oY44SmcL8rDNLxanX5v
NZGbQ0yLj8K9AxvXa+/Yzj/Kt5jbNMH3hlwmwK0GtETaiAeNzC5WKo/x/+gk
ETxqd33KVGrHsZkMfyAlc3Rzq5G65SB7GI+c3I63aUE+I9aDWQJKs7XSs86N
lbO7OWZDgFccdLQK2MOtnE+g0DW8HdHF2MAA+TF4Ei6ziHFghFbp1DGs+GRj
WHV++UzHoVSjEqAEr1CLNoNLReP7JizG4K+cWE5HJ7EqLeYj9f5nMvLYLLb6
qz053XixLbJ9qlVLxuCE1QjooKOczSDIzbt1EYH5iJZg8zFl5OIAJ9gSHB6p
KuxT1/8xnmitx0iRmhkdGV96IUZkuUrMdJ4N2742iddsKpM61ZNQu4HnQozB
LpH639pJDDCojpOj7l4zpJ9qEJcI9tODgZIQchYbZ8/r28Cjcp4s6x8XwSGZ
rnDkPBhFrI+eRqzqIvxPIBtOQj8GXXta4TGGN+5SgyX9XarCPpgm0akJ9+gU
9jJL+nvflGWrzMHwVNWjT0RkR559JuRqcXmpCGo7nCPUrdmGcJek7lwzhwQ2
gPYDxFKaiN760caQh6tcqxGXLZuSdDmtvbLBkRrmsgW6TYL5MBhbOCLiwJ5+
MdYDnF42vQ+w2mPo/MGLhHwLD9ffBWiiItiGGKTYU/Htvk15CCCjlwMXkxC7
WYypUujWMDmxHFvGntHkig4PPSALnYxRmfv6MolzdHivOVtAGuFgc9goFHBG
bZH3D4ps6dmt2Pj74Cr3uD7ajgRajv2rfJ5WIY390vOlZ4eTUP/ERqEZ+8cE
i3fE4PdoJgUFSo/IlkSPsRAHOcDuvqO45gTP9JbPsxf6vcn1QlMHkbyXbsoK
BcuK1AdM05CF0XABIXYZb2sNkosjop7S9dk2f64C6BbY/U/B+YOkw5dDToN1
YzH3zVfbA2rhllXSoa1HHFQKE+ykJu7CPCCdocxUw4e0Rvuz2MsQZj10kP9u
kMXHZFa5EfQvt5bR4oAL3U2wm1CMDe6O7LQl6qpC0UkUwh4pJrdDB9EpPZu0
SjW81CJirMtR268Pl8JUxzQF2sVwSKJnb0ch7qZiEHK1x7k93sRoG5sWlHp/
3iBp3JnvQ6RWIvjaxW77SnU288Htw4laSg499WClASzR4mUegn0Qf6ohRpDu
lRfSGX39mbxz1DcceTDJwUNbx6feQKU+3uQwjVk5f//lVgBrzC6vUdNugLUN
xLn/uLHVPkklaQz+b5fnNJsFrBZDbyqerhApbdDnI77sPzS6zLzc28a1UePf
KWuH32H5nx/OxeCKeOPVuhfmZwn9Pk74dw6o4D4WJ8ZAqeEUNylcjS0D3B5J
4iK7CPljepkNBMYa7AdSI5Pm9YhaUFWvDsxA/x04jDAuuPGsIKtJcaf1VG1c
CImBe82bQobzcV/urrHVW3TVmq92/RogAR4xZNjnbFYieVgC8c886VXNxO+c
Srp07ySWoZx8mXNfCtONdPyJoDxvqNENwfrx2VnESObEPI3L89f0v2y+S8c1
3L7JDF/ybEq6wSoJx7yJ2YWfifijI0pzA93YkgrpAOgVNVPLR0Fuqu4J9MlK
u+HMp0stTz9FcFv1gMNRwn2LVcl/w8IuR2OnLeVZpntml+gRl367dd+mBn6b
fKIE2RVv1IYP4gUwiHrp/5N8UYu20VGIacqz36s9UwomwRizYhh8h25EjfYX
9viIMMH3ZflRCH6jcNZT+K1CzoRD6aMUbJ37vjPbgpVUnyE1d5p7t+UTR8k1
/FDQxB1FxlcK+BUUcBAlajtgFyKOMB4W20mJEewq4PyNWA7z0NLQAo4Ni/h4
xSfGuzp5GSatC6LW1HeC8YmlTmwF2cgNLvFvXFTbvpeyshZe9184nOf0LY8q
BdUNk6Jn29oreNifFNQdzdLIIG0HAsYf1cuzmmRXLdxlp4kam2ojV5qppPad
MNQLnjXQuVAfZxjncgHQIF/62y/HI6YxraBy+qGimQVVT1KA+MlI5lRRUjxm
E3PkQePjQI36sQ406NM4ICe9RGehYXWIL2VTf2HbjRuBJ2uCipoo6fpZlcUj
FedSF8byGWhtOFGmhzdXvOAokYuSDb9YNjNkYK4IlqPZLZfPAQRVveCmd4qO
ElzvQvoocuVoWdQN+j0FoEHb6N/J9pCjl7eyEkF6ctJeaRB8dp9B+qap28wj
TEENUb9vabRwWS3IT1GaJk1XNPtUhk6pi1bMf+Afco09izESTAf8E3lgiZWx
MjDbxvQmTZ8V9rKNZoDHxxwD3Naiqz3kmfnb4GLpw/SofJQa2lu+eN6ys1zO
Xn+EqUc3XMXwwhBclhFapQDyQ7kv14ph9Ib2ojWP6XY8u+VDxJBAx/hAcv5g
p6q6xGfFX4OX1kVB8dtSyrWz5A00PqdMpp/X69Xl2GidYCMYc8T+AERsp7AB
z/86DN+SLvoZQ+7a1C9KnJvJrcFfiRctoTsyo4g02ykIV7xIU/Vu0wxbPYx3
MItD/qyzqB1FshgaqQcrm0mMqx0Lo5kXanX3ZuENK34eXGJbRVXSQUeWxlzk
0z48KY4MfpDCRGmQr8Yo24v0vnAffXBPjaCjupWT2r4fAS9HWl1A9qCWnKJT
+ZDCtoVkgRUzOS4ynMrdWT+gNHQgUU59ohQGlvM0+l7RqZ0uSTtKt80T9K+7
Gqj1x2wbWWTvDmz7XuFn2T2E+jx0qsUF3pVBAb793qLRbxKYU//Jk0R6KCFh
PsM3XTRHFdOIC5f5X1hOBLS3aZ0a4X1H13RXBOD4Nxu6czUE0QAzVaJtnndS
0KSaXq0X89VwMsR9YTN/vmqWlvWskqZy4MrE0DCz6rDx6RCXE+qgWHxfNXD8
pFlbEWbwRToVlIpnayUmpQiVBQWFZQo2NE5DbZRbwHRHAoZeWQeuGuPrXBtC
ZkKYCowJZafHJ/ZMtVz8KItnLfpv4EIHFTYaiqNWAuyCYZniGSLLSrZ2B3xW
S3cJeoTdc4NRWdOkrFmVCz7GFQMxmklLJi3HHfc6+CU5JXNFOLzGWXrwHA99
s9QLYKVuROGDYJ1bOmzjlEfgJQWpZXB8lYv3n8GM7RVNXhel7X/8BAdQXyGk
dfaYC83A010jnbESzWNqO9lVmEtmqFPkrEHpdPTt53KAc/uR6qxuNIay1vjM
Z0F7nee2SWpWovriY/fD/XtJ7nshugqDh5qKe5Nwect1+6bKoeV44fd5m3T2
Ga0TLawvIsi8BM0WQ1GC5FxcGHpMb28x+vKT4shKby39DmXwmB//8pCCVZdz
l0i8m+j/aSzjI1MLeUMeX7ge1h/cRGLRGpgzXtOS0YBxVKmA3UdLSyAMvmhe
YOo8QJlZdoimaxj79X7dGfR3qGMHVAYiIvOHMLiLJTyEutYOVKUj8lysaj5q
GBTA8tRijbr1kf5/Aj9yy45RWbxeHNnCUTRBNzd86GvESQ4J6mawurth9vlJ
V9pvbsxEvlj2mgZUdw5D8pXpPcPTMFyyFvqHqJJGwG7s0IqoMJ/UKLftKJRz
PjxeDWVaCkebDbrNbUFcKeTgL8hBkNFy3bYNPMTgTdBjENBx9QM+Zdv2nR5u
Yd80gtO1QFI+OKVB2wDGj5ry8HwaHhCOM6rSJ+IXgJApfyz5U3ti+JZ5iPW2
U2QZ6XoEfMY+Yyls63MU3KiQx1HiiHCXCjnmrnuI4rGnRsoec1awWKrPcPyu
pv3ymPpLVBll4+SIpeldjEUZugpdpOEFjWuoDcO+5qJeQ9u5lxsstk1SsCO5
QCFybEpsCP9sXRny2qfoF1YjlelG3NKqT9YQcZ6qZh1BRrabHiwk7kbYXz7s
jP+HALZqdc7mCUSb0kM3fBQtuKXQZ9VuNWnowiR0ymeHpjDyRVlnaZPUDncy
7QumwAXmBGqITAEbOsFnbPtt/uDi6B1zu4EScbV7YT41FkKJjF5g3zpgVN97
skONxnccTQ9nm69VvUpIzUeXzi4Oz9ZwU8gENtnTRkcCqwMYjpR9kqU0AfR7
0WXi5bHOiEu0SHIEV0x8bCan2AMDoOTbfnWqBKqu0ahtGENEM+yvuzsYRhz4
fOoZU511iArzmN+TTWJZP6A0oXT3DUn2ELYSiLKdEBRPNH0Ekz26ACuDx7/x
+t4pQoMupn6WudDlWKBTNzXmydWjugQokWzFN0xDuCrpOp3NMP/PkuSIzcZB
6H8jxf8pgy2AVOTLl0mxqBrn+qNdfH7bCRtfnWLeedc3JVZJxlqHLN2JhKkD
NTecXl9U1ZCXPwtKgVafDsSsV/W7Opa5A+jI1e93G+oNSIxMhdpIXJAk1ejl
cJ7rQajJ/h/EP4JwlLPNAc5+P1+qJ5LXF0RogLeBY4B8L+ycJKhmf3fKWDla
GHHocarqxhX04YdTAUocpD0Nqs76vpkMHAP2wIPdEAiOT/VryInvgdnh+R3g
GFgCsg2v0/XpYbrArnshI716YLwWk8VrGJfS9lv2ikeetXIKiXRBimuYAMtD
mNbviTln+hdBfj6F9auiQTXKq7ztw5g0sT7Zo5BMZg85yye3LSQI7aoR8LaT
2dzXU3cKnhG6hq6e54zYTlhtROYlBDxXyh/YEc3+EpHaW3k+Ym6hP6fDH9vh
yXkt2IKv1wSpv1EOpydWYapGc8RfFGFDxgZGMxgeLK2jVMdCyfp7UrxJDnmD
dWpfAuJs+xQoIVZSyEQQoaSu2Ej52/BX3+2DaJ64fginSf0xC1cQ5IA3dxUw
Yezm7niyCBysimZ/koS6Rc1TsUxVOX6loiYCaNjb/aDcNqTMl4CoLmmlwZ8Q
PjuRBjsrpyfsx2JErmMbUpLwKDnyvV0TXbg61jykPnvY9NZiEPpT+JUFqm4n
FvJWQ6XAJwD5Bo2/E+bXB6CDbPHU3g/P3n/YV2P1JmvBjzech9/JWzhoVPLq
NHQ2arFs+HkC12ysVMG396VQGPpJYvLmzAVtE7X/GzPZ3gCkjeI9IIKQEJO2
4HslYshV2YVRS88GXcd24u+/bPC5lHo2/ZXSo88tORHbSq4Ib6hM/+GuQ+JV
WdbmWdf2TGRPg0rTwD4hPWpQV5lwvVIpO2Yk23pdsHxpE0MAdLyeymKqU9gp
zoHi3lLW/8eXY7C0cIGnbBWf4b9SXAXryD8MJm2PY+6hPSD26Ibwgg8Gft3M
QjIOfzBs7SDJi74ztAW0S9vLTmlVpl5wBGRrxOmeXz22jzJplaq9MCtagV61
hKZP9W7LaAZlwarahFr9h87oEoXRX+oAN9vHE0R6h2JoOdYxgmyCqLPUxFMs
KtjhheB9Ffo1fiRfohqlrs6ai243f8k+CVJZ+PzeOGmA64NGVNqrwPcG7RiD
uqMU/F23c6OapE70TE+qOaucjxV+OSXuiJCzOTBZepAxfr3hJf1t/KtQ2IOM
js2PT1uLsTQNJkp35Y/Qb27R4BVhhsrhus53ZgfL0wAmROKP8pz1fdaIk3EO
P/IHFIqN+mJaJYsCbknv5qSaZXtHAY40iMRv9BXfFabwJ+5CsxLyv6gwS/yZ
0vC0XyiAvu4j9cAQnQLTgsrTN5/vYt5NiIGGhu474BxFGkS/m/UcIMVr+3Sh
jXf+Qblu5OtMxjfzuVY64iLw4g2gGkSu/kxR1xk8c/lhox8faLJtfCh6cIVj
3UgOopZEdmE21RPFSRnEw4ZF/lO8u24hZrhb2efse8J7aE+YG83cFIgo7D6Q
T3ZjK199oxGBgGmE5jlBulSPu/t85O1XQHIFhOD50HAKI9DNA/YkuhMsf4NL
1SxmKOvSKO9Fum+3cz9LA6RTP/DBGiCmOPt2BRJmb46tETrNgm2ReHFSFy1F
rbc0xaPWpHWV5FifhylbH2KOqGVgHdD6P9RJntBeuxG6nAYptA5G31JvPpVQ
meAHXjVG6dmzcN/gbFlCwYQkiArheF2yW17D1kl1pyHMgSi2csu+Se4XeBPL
T4weXz9uGUAZE67yX0GDzoZzGZ1HSgOVUSJRT5kJlcz1w7s8JxGKJQ5NUV6+
JvhgLO2Kwxqn3k8jdTkewp9qulfsIr5gQPqlRLySZ9QrrpGe8xcJ5JY4cUUY
X5mRKNK/naYaY0q+IIaE3szVdOYu5pbvVla4qdkefS/2OzhYIGlgwBREeOQV
BZ7CtP6ak9KdY7bBE7KboesOtsARuiHUzfL5Oy/gZCDUuJpeMH/EizssMgeX
e549TqHsou/e6tOg/lValCbmy9aZYNt2xDGe+9HsnBFUMuUyojd/3bNy3VU3
uORhDFuaXaEagfpDX710ssts3sCoQaYKrN4HjxCtayUIHlEdTtHMthsl0JeA
p/B2XNR/37OLOkelByEsMn2eL/3BSuaThsDXzIwNS57sOCQqmUBzMHwWZQiR
iaBEZbbD4toIuaP0CoTKPyOZvSE2RcOEgooQmqAvUqDLqyaJJbPLDvSfTn/A
sO6bEDg2D8pttudHWm225sPqUJhPsi6VZz7NUxiH3bOx+XqMyh4arLWDMkU5
4nk4KhSMVqJuyJ1hs8pW9oGWIhUfqNusn2jpPYPFodTfGPg5Wpe1gBW+/jrE
gL/VdrwdCLSxH90UiS4DWM7JJGoX7eZ5FMfJW2GrL3clib36TKm5qMSHPSK/
znY//w2VsPwmBl4fQQIZpcIV06Lb8XxJKaE79kT8DiBDCnqqwfZZ/JJSaq30
xlXEa+S8f2Vgo0fHgEw+a5gMKgVv/pfoQPZopDDxN9zHQJd+JOPS0SmjHnxK
je9zlEI7DYgvg/b7UQvupD1lHhoH1DJyxyIWwtsoTFtOdtGu1FgZgMUyIudl
vt1I3gulGx4gcStHvte3vpoAWe/fGaNtcIPP3ykFdwUrKerJDbpHVR+lMl9q
jcKZ3hZLEs/fO3zxXHhXYSh1PgV+kV3Z1iJ9v9gSnDIzIi/TDvj6zjfZ5ifu
JfuQzBNlSV+TnHWcuQQm5tlsdfuWlaKslAe2yPQufsx1am02jsky2nnQ4WcN
bqr824Kg4nkchxjNkRRpNW+FGYLsMWUoVl+Rs3+SBE/5qvv6DY8Pcbl/Z5tb
TF+TbqqE+vBb64j82JQ9KfW5DDgBhZCLiAbC5ONqPPGssVpYTmgplogv7UBr
vsV9pTnF5owo7MLGOlkLsUcBLjSh2vpfeGj4zEXCLJyIvrYVVcnnENKnHOzW
1+PqvtfHz4ZusvZaVHnRPcckirir6RSW01RLyDM1437mqHKzGu/iwBkfx46t
bqJ0bhB4fgqPWntB8AJkoUnMYyjYQ06qmWcbdpFw4CtwkL9oMIQl8eGAiOc3
rA4JdVPu245JU6YmXe6r8b7RjOTR7YsP0xUnX/ZnpMdrgMojMm2B31saI7si
DjB9OI8UvZwyhg/Wb9TjWAMr514exGuRSeTOyrg62uphVjEDXyQs+uSvtXHD
UpkkOZk9i9WnxIXX4dn4uivMQgoBCz+MH+HK1dBF/3yvkZLWH+4EgdFPhId7
fwC9ThJ35tnHatIQeKF6TrZlrlBXyqZlbQ1myhtOF89I3NxWYQWfkPhQXCWb
fkVdfZk9MehHWfXfjmY+gZLQr5eQYHxEX3HHMRg1prVYH9vAN62A2/VH67g9
QgTqTtf//unDftT1UpCCXylVXYE74dhf2fqQS/08VsBYJMCYESbhtaAbqRLx
PexJUcF6BOczJVarh/GKDOVoHw76F1pZfqfAy1rKO7wcohBKylhKjjcfbrlu
sIZbJ4AZijq4/Xh2w94L43B4PjJEdYzul9sxw1b4zmt1KvLf1p1rHcwmQahy
hIBfExttbY0zqJ78M4BgKo8AvybraSuRXo0ih2yb8/acXa2yDsWX4e/FIHUs
VAc8bGfOEkrjedOLZB8lC39kyYnxrh6kQ6UnqhiMV7AY+8J3uHs8ICpHazbQ
GnWW64XJH9JrdryK9lUwdknkwxktrhuNGj13pKBGzv7DsElTOeghLIPHsZDj
Mp1D7qS6Ez6vNWk3oUvY4ZjfRXQDNR54o+w2XO/P341+nED/qN2Lv1b8+DdK
42P1CqkM53tfwrjrbSWaSPP+2J6I7e+pP3HD8mb2P6/1kR3AtyFMf0D5kWSk
kKCsr0OHRYNupRZ7uVKzZ1VxYhTOTpmHmRNwZTdPqAdRsssYbG+WN/uRJhEZ
gprIRV9osAwakdAFavFQizzzL+63HX64MDNt/k+o0v/U6HLLWfB2pvN0Zia+
sy/NAMvKTbIPzVomvrDB/iTufK72pcpeKkfZOxh8INuCmK1oshRpcgtzW304
2F7zvEgIegdl1VH31b5m8WlQzr+rrFchp6f+o0+pf86lg1HYIFQtVZ78t3uI
9roIEtGfBfIYpmwxsYKJSOD3B5Uq85wruNdrqSWla1AWAp2UYFBKFW4D/u6+
z0Sz3HohtKdr7ZCh7isCW/t0ZEhfPZqCIrVIH9/2duyAdKm4or9Q0IAsyzs4
MP9REZIp3zbGRWrEaON0pzHl2c/kRU7ErLp635WsaXc/TZOdwF4je4ll0GKD
ylZ6duTI7ESfxRhM3AxRwLfLo4S3OGrM/ztKBArdumIS0rMa2htg5O1AXXzJ
XWTPMkBVxlX66iyAahlbpe8ERinSo0z3ow9+aGBk+RdDod2V8oQZQe5gL0DN
MUogPFktYWjw6AH4WfEyFw8pB9lxmAcD40hVSDIsURKxoNdgIciCKO0MtqfZ
Q2FIMwTx6B/cbsoTILXYQOySq/jwIL6yJyWw2iYjmNx+aBEnWvfdOT+3qsjN
u8bR17hsIcweR/Xmdl0ZliIbk4RJifoh/78eVE9vInyjGPgVRt1q4NY0txYK
VBqNVhUSUCdn8QrNq/FjFziYNvzp484+ZGoPqZBImLHRLii6G8ljZ13vs8aA
14Bv1BeUnacZLdkuPD/Q9MaEyAyP5rolalWDgEWB/ClX/6YMzlJXAgw6cDP9
DZytyhEdNYxW1lvsQ76lKNsoItoEfsY9sfJJ6XuuSHtfHqmeCXHv4s2Tk1sp
WaQOAc7mmpB2EAnZvz+GBWs2a6HLs9WLt2hysXH2UOFDxaAJmo9PMjImATDL
J97I6dhBGA1+erLs+gbkVUHODnZxr6r9O7g9fx9UUgelnl2KgzYQP4UGcUnc
hRJohiCJu+tLM8wVuItbjPCFJaSm2qxjgu+o8L8B/VuKX8m9IPvtMqtPv0T0
JmX4hi2Zqt/qOb3v6su/qZWnIUnmGGNpX1hrDBIyBTONCsZdUHih85w80tVN
OCWAefcj6+l7Gh/GU9dAhfKlpu2LoXsPKjpFp/2gfMNzlL6PqNWGFPo4YL5x
/wvlC5PP/98oWrPrNw10IqnN/vnnfNrhXyJR4+MMEGOBIyqevE/1yHDQeQM7
kmV8469yMERCtegwIToQ/XFbJLaM1n/CZfS+zYPlITVCB/P7IJrp0wiuQQsY
vsEi4BCbKW+ysGdAg06ezAH3okBJVWg1LjXr64zSWC5xfJb0BEcAY4JpO9e0
ijveptTRh57OBKRy2d3BSxlZO2ZQGD/C3IIvC6moDaQlQR4TA/08JY9pa4QX
w4QSCjorURFwgQhyJVxn8cSY4Os5KcGqlgJcIbIVx9Cnx0Vcyu7jDyw8zOUG
mujP+dOv1kl9edX16LtcN6cHpeU+A0CZ6vz5XZoLSI1lcJHs4RKbOPmAmXwT
w1Hfe9zKLVf3lSXAJ8afY97gWbrMnffnUsz63tt7pshy+4Wj9t0e1DNqerOq
mqfuANsu0WPJ+xb52jQJAZPYQXwtJ9B17gicl/xN/aAqGMJl8mz5suglaQqD
E5K6FD2I8uWdnGrjyi1wrE4Gqn8vmzJO/elqtm/IuaTowcxGqDCD6GkoWW3m
doZ4DI1DCd+5aVnaREPY+hgVW0JM14vZz4AaMgAo6qqKDFCkenrhIxu/d8YO
G2Ekvr42TA4s2vZrq1agd/RFnUYoc6CM/NQAueXGPQCbHgyWJb8O2QVlOB98
vbAI6YEm9nG/BJ0yyc8NnHtPdtCrTqNvoaUNcrdzyOZVLfvyMbipToRWNMUu
Oug4LlakSneVzjtV8rnspmFvTXLxzC1+CFGApApT59uVWAd3HA+EiHxaNoWr
dKlNxYe5dS0EKxrV7z5JB/pVUsbfJ0qagl3X2qFGyLmTHlQtdciAMxQKMrAw
yYZIvq5EnsatKk8LL+QO5eJUh4tiMuEmb3ZGUHlcFd5BQSn/38NkS2lAFAow
bEKfQov3mdDqmm2LzKjOM+ees/GzJwC7Y7UlmoQpwBOY1/WsOGXAP/U25sA+
fgCToTYtnQQksfzVdA73huy9DLAGU4K5cwJ0yTPoEoizDGz9FnGKMieNcyCy
S95swIcbpkYzT3OaLzVzPqhHREy+epW0zyCNy3fNFK8GMseFR+OCOV3baJDr
XT8xxBR16CDQTYpEf8RuMZA4PzQu8R9waRYgDQQdlzM5vKX7k8GKXFagwxaA
1en0saTwyjVtRVSQQP+iHjZtqsyvEVdxSSXRhCQ+fG14njjuHSauSiGuUdOd
/xcv0K8rU9AR1CtCnGnxjZVPTT0W4qHFUSJKr47B3oR4Ld5WCJpD8/N8EXI6
DieptAwsU0OywNQZw9fGEQqlDYqDj+9SWZteuXcbwncP8196DNOVdmw0t3KZ
J6CDvbPvCW8rwtfMX7rXRGFWxZlWQyXqbo4ZdkxMBUuPz97/mImxzkHKnLmm
Q/EoVbRvtX6Qv1UXhNZH00N0HXcNfHVlax4088nYcn3Kx7Vad3xGypnDz68f
ufIyv6nFoqAMGs059RKnCZQLh3V2j8wFfQCSYN3ADfv8cuwpWYcVFVHtYVqI
7eXfwDfz7+zsod/kXDXMIgaqRWHEbwBqdRsHDVByy0aYbloPzsduulpl4K5Z
1Yfi9BWikYLSEwt/agAlEuV8DZJm1xKKNzFmfl3bvFJju7a91Ks76izx/Thf
cVPVuTcSiFWkAwJALBUT0lSMzxX4pvNptDORQoMmW+FAdJXiNca46KWz3wRk
ueh/uJfUcAvySQRH5/cqWYrasGQyj1xI0KlfsE4ft9vpXgfmnp8hp3T+t/z4
R/8DIhZReT+a/BQPimulhHjPCjZ+tVgdyXTMUOAREtu732Pdwlr1zyqS8zRF
KhE4g/Ot2ZddKilelJDxuefDjSYOgP06CdZrFAabLVQXnJKPF2K64pW1E2lF
9ll8XNqpFwWggytQ6G1R0HJZD740BP15evLJq54cjO0NfM7XvioBdsRnWoxJ
nbgg2be0kQ79yPVzvhCN6lz/EUj+anFf5tRshWssVwzUvH2zG4M22JmOTC0x
6F1TNeQr617a2WQiGd7qGbM8ccua2G4/Y1UDmgONhag4OR5hSL5h5yZdrkI6
g2cPwNupNkjjOsQpc0EijlnNK0g5E/3PK2OUDPT1T8j2RFJEIufgJssHOu4F
LQVOPb8W3nXuqA0Jt7lcdESpw5d/Ck/4o2ThNrxXqtrHy0VxAhPX6gQbN/2U
LNFmdZ16dTCWtbjIePLrDpZp1JpfNMy04pRlOvpcgTeC6KvtCRG17h07GX3+
p/NChASjvtA1Y7jqU5hxhnQmTN1XvOZPgSyZu4NwpZOoKQCJ85YTDcwSbN6y
kmSwFJEisrEy/qyfJSg2G7qNzkjyKNgfum3nim4HGwn3qUQPNGmN/Z5byx5y
ccv5iHniEBh3xFJfVv9mFs8mrkMt0/xEcHGroKyRAcKU/xI7MlY1bA3s1+jh
jgzAOQIRkrM9KRVi7pIJLtLmifD0VdkInNqP9sT+zGtesXOZvuTE7+n0B4ji
RbXVLa8dntEqYowu5V3Ycblc4a9dbdKNzCBuw3s8C8GzmxBLSLz5VLqVyIec
J7tyPGjHi6zJrcS6r8S7qYsNuDwXvoZNspqGCmf6ZwmqhKpD/26++hkuIG8X
Z/ukbT1j0Z6+LuWnmRcTdvLfDNC0PgmpL28IrzixFBO7AcyP2nHrG0FxM0rY
+13wpSEdYbcfZ/WLq1LeprhPp19NMUW1EKvdqAIpjR9UGjbVfCY/WX2iSDz0
IyJOgOZCHVbJ+Po+AUjctFRcbMgyjcAlWnHMH2QcqsdJA793xYrq0h0LvmaO
GdOHDQEYIn0OQeZHSjQmrFFMD7hpm8Smt/sO+TyJpQVV4V3XG9aLt8ykMwt1
rwPZMY3ZpxglpdFeOiYNVVmnWOMgCxWBhqcsxkSYU7INAWNRDoBTZe2OGMQw
s5N2xE+lAKYYxvSnhN3HhVu/XM7ERUwZULBoBWba0ukNt+vfTfVoxugXaSYV
f26j++obGGjzh7dF0E8kwLLjAOYq704sGRFnlkJwYdNKyRfAuoFONeePnw2X
A0e6YlYZrD72q/RfRvNqxicH3QOVPm2UKDzOTDHRoqEy8fvUCUnBwQgWOYl1
PHb+bSuqo6wLy/sB5F/N38KfLBF8MICvsP52VEOT70nz0ywBFJ5m9C+bwGhY
HOIzbQYUkH46Js2667+lBSKFbBq2cF1KZ66AWXjoZq7iKmaOdy9am2jXSbEa
J+8epfEJ0qR9iuPAS1hQH2G80PDZYId6azC/2qnJrD2tOHBTmDHKQftATedN
PtQMVmDgyucGlSQCWwHzAo4eGFjnikTK82Qvy/6HPtCiqrDw6S8AgG7Uw+OZ
VtDGIVrrhSBcBTMam/ZeSlhoNhnIkgDqTlGscDfGAUJO7OkR3Sdnnv7dfdXU
fN8qcYphPBRwfpp43NvoeP3pItEFREbHxjQgbU8aNXXZs6hhvv5W43yZZphj
Jsuf0M8HxFGbtpDonMfYXg9nCT+okBR65p2GgsTVqEOTQbgjBAOU15dF01hW
Ibbz/7ED2Nb1Lv4aRwqFX7SX3RRu9d54UKXZ9t4C8f8ILz1F2JKLM7Z5GkUm
kLO+eh8DqJCC2FhpEz5gEnKHqhBFbgH5Uv1TZWoLSBF/A0oupBoqjTULwIlw
ALQcun8/BNc9B/aVzlqzKn72Bwe/JmBCozFKzMqK/ocRwnFRx/DV7BdVromW
YUfgNbc3x40FzQ8W+POtIghiP5A2JndE11gRrTnnJ11i9ofx+U0wz3QdH4rL
Jq6fC/cu7RKhClkYkOnPK/WOsDMgwODpfde7QivfKotHAGgcg7HoWg/X+IIv
54ba6f4a0ymWJtG8FBgHuxUUz/5Hf1Z0GNqr1VoMqwNE5SftpWtFPJeA1W9/
zwNU/eVqgtBROomSwjVv9bMGeqymAGNGgBvYuULdVTT1lnvhBI8hk8KT2jZd
wFjrk3LArx21xThDS9GaHh9n0+Ygv4W+s2vxyTWy07QLGnCjUkeU8bTeoWZn
Ad16jHMgm79eV7H18aRw9SZf0r9fyWSfKXG2oY9sdCvK1nMfCmQQ8spONkoF
B/1aIf1SDrYO9bSMLzQEFdnZOwPlEAALWAuT8WpVqOLrUsRq98HlqeQWobhO
rAdCtEO84ykGSUtc8Jx78XcyRMMDljbkI0LWoC8aPk9CBoNUK2EZKI+l3QP5
1SwtG7h8wQp0o/ITNRJi4gQX1mjMjNsKg0XtApArmDSDAvVJ0Zz67EAO7o32
ETfddkcWPEw2fenbNsgJwL4qfVlOzXgTALN7OYt575/Nkt03WRo4UOgyMZd7
vecsNrUCCUp7rC/5M5UqtyQJoE01vjTDlCudXKuIyR5n7RBcf9HgFFVJeW90
FRJHVLjwHENJsfZLsoFMpf1Qp/loK8tbUwRc//BzuukaY9xcqEqU/pX1+NyX
+F+2Z+v+ocVzgBonrCA6kp1mWai5jmdTQIFhHYgbHKQGWp4PBr3Y3OXIZHIz
7v/Zjilc/SGZxWgLYxz27BjfDZUhViSINvV42YsvaXQ7ohxBqQOMbKgHUKmK
iSWI5nvmpn5YZVbWsVp2IpS9AaMoArLLGbQHcShbS1JryZ1L8ku+ltzX9BXn
dK5rAAO1lnpEb+GMapyMlvbtqkHOBRraM5JDWcnDZUBvJ41e0Q1/B7oMUj0u
z3H0o6ENYMq48jaR0OVPAA6IO75Kf+4iMq+AjSIGs6fvOf446ijnF1WtOk1g
Co1+bG+3gVcplVZ9IqPyfX+xsinitIX80VdlyOREML7p3FaUQxMQWHMcFOSW
09bNtJWDFgtFM5XCuuMrLGrUnWuuJRgqOoJN7ghXfkB0454VodBEth3t+lcF
lwb+1mtOcy3j+6EA/hrrF8seDl/Wfk/U3gyM+pC3pF5E3csTdBg8JMz6o3Wd
pStHSGV8uDcnzf4VoQnPQu1zxIubqD5TCWNAi0KWtiOWPgDI436r0X+1/YTP
BssfjTobRgN83pGdn88K/MvtIbNWM18597/xZ042VIqK9lOaxpXk10ZaqOHE
EAFfnVoMZGLoXcZp5Nw23TuAjyn7M1VIUeVSV6wSztpepiihFit+ncodvA7H
KaEmJcHQu8wrOcek8P2AVb5f2enOdotE43v0s+rB7GhX73wm4WaBTe42aNUD
cPY+/Arfd0wOyM5RH0jETSfJO2ldbwNVNCwU0UTI6ZbIpIiVus61KTO5dk4n
z+9RYjhUnHRBx8EX8Y2MOo9bEjYI2tTu8eW1qL5EbAT57eEZ8udH7GhGe+lM
U27CAuzvOYDYRUxchUjrohx2kZxe0IHC1+g271Ps1Uhjiz0AwCDosItYUl5Q
dXj4thABSyjbvR1VNnYhNMbaTVb5WW8YZ9WZAUCsCxe17ipIn4oGA9HaCnMK
O1Jxp2HMUlk9UV5bLe4TIqh3Jb1Hh0cVcdhOVznP/NaNxZBL8iWXnuZvEhmx
bBmwksWpOe+hJA0t1CeXskR0ThezQ1gnkTDIC2ma7scOyRPvXXssBCyZWLBR
2KPeupAmbB+X7eLY/rPh/OHHokDJJ/AswKM2gXbm2Us2NUTIxirSrAzIigi8
pT5TKPni+z0o5VJ1tHW+QTFduUZ60Wlncs61LSf+tRYgOyldMBE17nQjxa4v
hpeOrtfy77vSm9QynAP6WPyxXHRsz1aevSqfVjTGZ5Hi/sXsGVhLbBBHFiRK
UvtOyTLScbIv1AM8tbYCapgidh0CZ1Nr/MFDU2YyxERqd8PwhjdYhxKfewLs
y/nZ50XYeI/MkQIVAdebqrMuJTouGUAtezRaFJUJLCpg+5MysYNscQr/zQLZ
aIPOMg7fjGg5qLnkSC8pzI2BsrIq7SrNwjisZfQP6Ogkr3wX9St6O00oic0d
hpuIOclfgZgMUW8z8ShMBtk/tr8tHKJy6wQ4I8YWQcfVAIzTttVFwPldeWQE
c6rj9KaPBg8PRiNZ3Nd3xoRLJ1TAHzn3qqkOgkKgpgy9GiMyuz9Dp+3OEXKY
x4k6RaBW4G+Z9Fg31c8sJlLWQKCnfzB6fUOM4WBAitbrAYcNNkrNqDqWR0pB
swUF1pVYskLJj9CYzhFI/81ZCmFA/Ft4LJ5e3woKbqJQOPMqtRbd3af5oU/g
eys+YYWWPbE3eu+tQNwhN4cwBd5HFi50hd4BFHHgtvwtSn1NejpWfv6HpdiR
hcBYav8E1z6YqEMRgVocnoGXMnGvj/85Lbot7Q4CFkF48KvanN52fC5wb3uD
tJUUsn/1a+faREgvtwZR+xef/amABGg8COue1y2rLrpkf7LtSdygYydqHT64
CheCHiqawnh6AuGAOLojgY/raNEfQ7gKZc0SZsj4zkzzgso+2Wl2i5pt6Pyx
Y8SE/ImwKnySceJm5P3RrbaZt+0usaTfOrYQvcVmnUCBT6ZMvMd9POOM1dRI
GxITGuhDhCBAskil5K9GbssQbzmZx62fGkXrGQJzuxleb+PMGKr7lzOunjj2
bnevlGGJWC6PyEgtUVm3aLXX9SJacpSh3soVWPcE+238326pwepjcyyYGnMn
lNjlYEQqiBkGGQ1lQsinurmgmRlzEVPsACVQ+facN4xftxnp9O9TfEhvF305
nXZ8podDNc9v4Tw3OgHFifIQ8BFlhRpC4XAQv3IgRXCGReKBiRI3uDUw3MZZ
umpv+71AU64JnL3E2lpSBTqRWumXpjag6a4kY6XRet4VF7RaW+zH8JSaSABi
MyUziw/T7AHTaa3QujyIidL4mOk4/TpQcVZQ+sXCc7FFXV0TTyyspFW+WL6N
ty4NbKenhyfr+D7Z15ka3tPm+KeqE2qniyNUUinoqQ2lufszkJe5UyIYOStl
wedkXMckPG4TKjX4aI/PduquP5TtNDrGsvuDEcQyfqXus+EhZkNDuxqOV/lE
RJhjk3l2BZIb4Ss/YnEKr/E5UMsf9IWW2Kj3fs61BG71VwC3to7F/Yp5m3fQ
/tsCCRaD8dpHHP+pdLi+z05j0Eh5Jrqf/0rq8bykJb3ovncBr0Q0KcV5CSMR
+J4tWwNdSX7xSb1hO/dVn8gYaDkZ8ZcmGQ/clHTfYzboeKl3w38Gxj3OrJ/i
rkZe5Xo/wH3tTPLvVwI3tN8Su4Ob5lNRRJUOwfQAxAQ5Tn6dS8/EkVgT7oAZ
wJlONm27vkHBiucAu5bgDU4L9IDpcAxoJsG0u0gCM6BcfTfReIHhMMYNCBxW
Vz+5xYEzWtnyiehupjxMh1oYZoPn5SOGt07SwIFl/guR2xMsBmBZHsk6y2iP
kMfGBNvaXAVJHTraKqwUfJc79o+qax+CZXYg/vIVR2zbzNGTkg15lAlt7DI/
OEykVJbGctaQpXQE4Fx9t5z9Jgk1tjMTsenygx02Asu+R2wBbn3i8OJODbo2
f1AniyMAqee6uYc/08nwsDWSZUDEMT3Q2AKCY2tKk8qZwN1tJctcmRY+kCWe
p0po/sHcU24mBRRR4z48gCFYtvuhDPEOhTHh3A3BeScBgm8oZcWqqhtBJVfi
hpFFIO5fYHGTUnFcQSXdAy8pLCSomcOrXUa59fOmcO2Z62U8rNvAnOEy8mUH
LAvznxXJEiQLotm59Oev1nVpnq43bhVb6sxs0rkn3qYbc+BzdSl7n+ylloBm
nrz734PJjmCzbhUb+Sk7mHOQm3lBcMq7a5ESdm02WvEyrMz4UC7g4QovTSUy
961ldZH3WaGAsNisBbkQ87X8SI0tOWfAfnCWY/0NxOwgibHfbfiJVCJ51k2O
VJxs0XLyPS2wCS7VOs/hEguzcvXgAudtsFBNzn837QKsuQizaV+KtNJOXlKS
g15K7uj8cbMmq/b7JB2Ir073ZCofNb9EsPjpzyMRNcxmmlvfO5JrYOKkX72Y
4cGL6z1wsz/LYYTsKyV018VscLu3FC7QtwVJb7WpNDwGc8U5+IYzn98BfQxK
ptKXIdZDUI2LGroKrv1WP318SuD3HTlYR8N3+0VLONVIRkKiW9dEzjLcf4dh
EasQzQLvpHi9YEJOxjkRHItow/NxJIw6q3f/88YO0DNon4/ucRjatzUazTBg
62dkvuZ8bEem6o23WuBj4nYiJaNd2KQ0dp99uTt5gC13kyr6z8E4+++sxWKl
qLyG8lSsyoMcjeyI7t/We2+0gpc0T93UGCTzKOsNTTlFdLVHWvZdLHOGwq01
t31YanTwGphg7Mw9sMKRIXCr6vV6hL3rrRvkIOkgStOL5QlMA9bOfi1aDj30
aIX5vyspnDP3JVlGSglM1f8WHC+3te4E9nD7IT5r7lgTVyhtNKOijQHbbaH9
nZQUmarEXV9a4HFpiuT6yNR1XxRgmYzlNmUPFsqZKjoRZ/KuLRfZCxH3nFlk
CBpJOOku171dZbZCI6dCaPKAEB94iL6Dq2rI/izHAX2G0PLDzfThyeXtOhvS
4P212TQ+r53u6scgz0yQoIK3pgblEJpysV0Z2YFq/nQjQtrjR/0LSOPGD2JO
2J1Xb1+kJfAqHCsgL6F8PGXEiHYgjMTKGBzFNuRwYe7faCfAXZ9jP98jC4pe
Jd43VN1rQzCeVjmB8c6N7kwEbmow6id9xP5xpmHL6X6amXj32fthhsUi7IAs
+pyRs9JbiYpbrQrQDLLyoO4bAHlHnXV2B5AA/Rc+wPtcUNT0BvJqwJgPhPQA
m2oekeRR+6xyo6NpmqAjg6tnDbs+vsf4xkpxJNwlc37eyb3veQMGfPmDAboS
+ATA9u/oatJyLThap9eNp59ljORNewtyT9qnycF8jz3yv3NimHmhRrnuGT0e
8+5VwSSzS8bnPTmea7JgxkPF4NuM36klUnAxqM0LBKf30dKuU9mLZFLCdG7M
LxA02kipfKJstdzQwJXzMkZ+cxOFazjBnTM6WCQFtf7yUlOGu7N8VaYd2C+x
bS3dSNgbeQa0cKyrtgJ1jb+npnvL+nhSunIIW6R1vJi5eJx6RTEKGlq2GwYZ
0rNcH557kZ7FWqK/iIUpg5QqviqW3pQs3rVvRj9nmfNn/pzjNaxQ0Xbwofh/
/48SF+cyvxczEsjBf4D6rdadQxNzqQCtsT8ZcZ8PiU4vlhniDU1hDRMYmQ3l
gZvMSp0B5y6zokOB3UNEDyPYPdQHXCwfxtiPuCssTIW4r21GTFWvzmzp7EFS
3O2M6txbuvMiA75KDm34r5bwr2EIxrjKmotfaspKr4AcX0sxXvgH55D1Xlr7
f4rKvbqxtEVxF+57BSjDlcVMBCRuJLgVxLjFCGExynkzcuHvRaZPYjOJpALd
RqfJTT2ZE4dC488OXMSJi+h8B/zbGrlW1o+2axrEbPvOMaQ1Ha/+COX3N+HY
5RkL4gFvjqS8/CCZbbmf9YEEvUN5NDOdfHg4RzlnQl6imcnLJmEBW5k1MfBx
iuQ+UPQwUoqt4Zr/Ntcr2kqSCcpEA3Z8LZgIoGUDIOCvU42TuOtNDwarVJeb
M+9ZwXtswUmm/oyIGq+ta+AEEsgG5vgEBxfBjMRhCJNcbo7zwYtxoy127dDE
Ctt/flObMNP8Ja0ZnGzPduQR+7dqx8cPhGvNUL0Rh1s+I+7ixwUo10piBark
ojnefkSVm4qShqiqkLokFuDPtioDtbSVfp2uWNi91tCwrbqJPilOUv8ogSe7
k9f2nzbKcFrbhXFaA+vqjrqNT2VH2y1DmE6HH8KvtkdqynHI82R/2Jy3vW6F
YMSC/bMpfNB4puDrSxJijS9Jyu0UTQSANP/LzxZS+BE6GBMEMkzTv6+OevKN
DqJ4H1rrRD5eqrTlrZUh4bbjr6kSW4oAQf5MbZ+J7x14LPosly1I8CLHEZk2
X8fF73jRtNp2cVJCzG5VClUG6I3JzfFTGTLX3MxatQpqK0lVpuerYJEEpIjJ
XSViNxzZ+hBrOxt68S6jbf/9D5filmlkwhebZxLVoskCYPQz0MgbRsryXURJ
CeNFXr52w6olEeqsg7U68pnJprNFxBlMunAjaVl1xSUK3d4OLLbrIU88XKwa
dJmKvkCnQ/naddgMRjbJwMAdkIiDJRjJYqTRqQPkUWtq36Q83YbsLwusfr/0
WAtzGMqHji+sejCYLuumGBhmdDiBAgB17A/QS3UCdAiykz+39tcc3PZe/g7o
Kxl1uIfWYs/lS76G1M2snSXiFXSkiIYdxyC/Rf6Ol7it/pD6VOjuwZBk3TIQ
cgqq3Ca6+PY0fy2wOA8VJjtdclcFrsKmyvadYviQToqNpzDcl7qFuPeGxM8s
Z7asUsBYbjXsvJQ5H3EjEz/J7Ku8XEFXs2aHAgaphpJAHeuRI777NS1DN23O
Cgqk8xtAslE/Io8JjBsHoFl9CP4iL36jGshwZDctb6NJT5869X0ZaB/GDP3q
HJ6UGmdwAupdq4aKOyLMop7M3GLFqIOx64+Cn0H/vQdcXdDbp/b5kdArPoxj
NurJ1v1qWwh8IIHxA5ugCfrZXnTg68dXEh597nhDqpDCitVszASfsEQPIOMV
M8EzKJQyUSz+Y2kVig3ujszEkHVhKAhTrUaX2/loypk4i3b/zweuHaIRtNrp
SGgaZGAtAFvZ5Z0wD6/Y5+vfgvJqMGgBSE/w2Z/0SA3/ohjZV1vaMOpzr7yN
+TvXfnn5m1ipZLMskX4hetpT/scndBOAzD5JMc+lDpsq7f1RFr7+22aRSjhB
mKGMY1WZHTU8xOKgXM7GnriWr200k+c9ylZdNJobLLneesmpo6tCdfpZbsO/
Ybf3v8n2LNQup2jxjUwiCwyhTdE8N5+MaVWDRdAg/G9HdnH6J+LOs8HsNIwf
Ld7OgS3GQ1rtQ8EVY+qi1EQvITfdIwZwkfifStA9BBMcO+uHgk2MzNqdI9P7
BeNZ5docuRVID5Pyq0KD8DuwVCoCxahLa9iY4jtDE3QMEfWfR1e9JYKGfBY9
96A9cxHmkp6oc1EtIs4U+Hl/LV8FdRUvj8iLe1RDRJ8rvVUbvupT0AT0YZ4q
E3zR5gip+5XFIJL7Q6x49ckZux7/NIokMr4ATYFQh8C42UULBvIlWm1p4mFa
nQs1ebQj9IQxOfucC8CdGa2EmIM34U6nL8XX37z6SgQ7Plg7Ro/grr41qt9D
qV5H+TY8iruwDxZL270mck1ShBT03v//PcbXAvzDFkpw7yBiMvPRb4RpOnqM
3uwMXWdX1H+8qe2qVse9VFN9GO8h94vaGmq4HFFnyC87BN35askQNypNd2b1
rYvOgnjSEEx5Wv2pB5i6w85gde0ko3it55aCSiVgoj22Sn5QHVsv1Tnpn6Oj
HmwDgPkRWR8UgcU5KsA1UWwM4BlD3WZ98/3zYzUGizQ0HKbEce7TDkejOGT3
+bn5fwdVPj4qDC1Jdhqpmb/r1E7ueYzHXaMPrQhS9lm19loQ0y4KPTHKSwJg
DELkvhJnJUZE6WWksNs6l7okkTn+VtY5F61YHTaz/kFW5ptJ8d6qnUhdXb2u
1ONA7ht2zQd2GEY7ijdD/fslISM/G5a0OC6sCsDqnDJ+JLidPj5o52HFP67m
AliwK1oNVq9qlgg5KnmYwfw7xizVJMkMwhfdfa0hMtdOrJXiE/m9ZQe6vaSZ
HR29ux/6BD7t5fFDIxpPq6IHuPy37pHMUF5SmKRrShyQXxIpwH7sVamywP+N
Er45oVEQ4Rnfl4XY9RUehNP2BB9yMN+lrgoN+vSzOv7mjboSuq0bm7H0rIeu
7bWXQXCRoKUSSPGkZ5Lp7MXRIfsfXYYahecP3ZIyzd+I8WYWI5GFHrqi26sL
aJAHfOvmUVPRRk1OtA6kGefoe7LFO6KvVLdsljx2Ea1HQ4fhwOoHXFdJl+tP
VKBeSCp70W8AVZ53Sm2tpIykcNDQqL+4XzdHGJHIUitKZaN/4J6L6+NxU5d8
p2NngbiB6z8q4fSYFDMRaWCoivCq8ePVUoz8PLpgo9EbkZ6E27aS66CEpMLH
kxlptB5T2Fwbkruo6R39lR+whCS3AtOA0tHciFsMCHeVPXv1l/YPRrGAwcDz
guGglMVjw28+XMS3wOByso6ova+lFoPTkhinbNQIWihqaIdzHUV0u0mqS7LD
ROH3MjObGqiZ3am1HdDf87uTBXc2K8gyE1/gW/GL/K5mq7XnCwz2Zz/IYuQl
r72PzZlKyHp9eHjUvMiJwLYy6Ln6BCrPtrz2CihetjLDGiaP6dvNtioGb+Sw
eUEkwvuOPY4byFM/yRG0KwTQsdAm8lx+/YDbbPtK0VgBjxfBIHMXx56mvyrW
8QSX/gcJ/DjcfJtEX5GTCfz/Aq3P/BAWq+y2IIzB1UJ6l04eSkT3NnLOa9jN
na7UuISj/lBT1JKfRec+XLgkzqCumtWMHd7vIsPB0z70G/9WUvVwq9jl0y3d
qxMCrf8sCe0swGa6hzLzaC8RKFqHvKCD/AR3DfQ10RTXSbWguCnvj04Y6bBq
g2ifZ1GoeTPtAaAoMQ2icPfB5MQwKe3yqBpVr5013a5Vpp4naz+8+Eb2RXw7
6FCsm6ZCIrj2i/4BV40WPozI8r42/IfD55EUx08ZtjHV4NzajSkokkhsvcj5
DM6YIehXbSuJTFnsvj9SLa6qL7m173QYZgM1fdMbj8wrlDvlBeC0rBSygRG2
0GEGvG0ZjGcvQSbS9igEZe23cVMbjKtoNXFfvQb+AeJR3ItUppEE9Qmbmqg4
KHODK6kyNGSK0rZtpGnlTGo184yIld5ht2jh1a3iyvLajf1VJ+t4hfT8W7bt
0K+Gr2C5hBflrPLPadO6kGs13Mn6vr3a1HUf0lF2rI9N5Dx590qnretmhce+
3UrHXIZkjG9Y0e5rUM1xBSqS95CS0jjRTaLFas7fXVl51gyOgjDBMPS6ZhzY
k79O8KXoqk4myCTwF+2G6IdY896IJMgoavOs9p8gackYDnqP/sWDzV5N+rwE
UPDXJ0QmMOvc6kIdvCPKs3jsGv7Y+t/gTmP+BrFv8+22Iwtz0yA9kR1jljfk
hgyz0FJVvm52DlTdKUybEwzIm1X4E7kensgYQfOfZUiHcczbs+Yi3SxR+MY1
3yepMtJPjU5TYF3F5zKpS3fe6C7bMp3OYgP+kxG1Fh5NRJ289fCY3nXC2od2
TRuMTEzAVER/08Frf5jmrz1QQnNaDYRgiFrBTufMAvmKXqnLM9Zru3yHOUik
OoukC93iKB20nNM56olP7X5jnY/CEJLKJnwrPLMCt2BXw7nR43QsC+jrqH3F
+hzesfpHAdYLpNSRPJ/A/W6NN7Ld4tErQYM7R88OOLadnQfPZ/b1huTYU2DI
xGG7J6fndZ9Uy4yYwADgVBmsikYk2HMGx9O8AXuwzIV1fFg4UaxDMHSlx/Uk
/KXOH+2jqwEiRI+/kX/jZMmUpRA60rlAEe8Q4q7ng+Tcu7IaFmBtEPO12s4b
/azbmIZY+XC1/nSEY0MzSl9qEmSSrmBK0oTD3jV/A0pvpTB2YfKzP1QPimv2
SCEb0hd7dbvcYtsIuF0Lhh/omyW5UiNP43B+lZcS+/zcoiv/hIurdJpG+R/v
BeEuDj2Jf/MLNEmwrlk1s1h3PqcluSMHDn6TL9QSHU7uJwEAlDZhmidGYWsn
rWKSDQ+LvQSiuPZ1ajoGiQbS3+IwqEuVlmUeOEjbaIYghi8Mkw9Yb1cnBegD
rNrTlu15BLu4LacBE37CrcPunD/vA8qdTnjk0QhHDw6HawZbcGtAnt7F/9zf
nSxggVOWqCWBYZp8rQFMf856F2J+5Y8+WDRcLcIeN3zlb128WInWCFvJxJkr
0b+jm56bCUrTlicC6RVu9zW8naj+tO4TfY/hsQ2fX1Sv+FdlICx+vaL0Smjm
3q8K8wlZjwglDc5i5+2x0MaQBpvAw9rmEbYhPHOjFInhFslXhl9uTbwlt0yq
PJM3cQgL9WWIuuhPL/icIY3quzkTsz7P/zI/vlVyz24lJCkbvV7KkXbdGp9C
ha9byNmLOkywOxknFYWpucXUprHPOZXejITrLTQMQNgZUdq3qEPnKSxDSWHh
Bg+P+rAEVSiC/yNmolON29hjbRDE1IgJEXnI0sAiv20nuxs2l19cSlFJhnng
0+se/nyBzawanZz8gCHm1Lu5NciMQmezkjIjpVZ8S6yBDccCFfesxyWauyQ/
HMgKwFipIwdpC2rrpKn++gZefk3wGLJDl+N8qlIttsXR80q6c4EIF6y1Am9H
8KjpZIG/KKvmPIFiaTDUqCqqbaakbJXFNfxOk6umh3A9FSMKRl5pwmcs/+eq
WZAjnYH06+k7np+VtajXPDsLTnXne6Dz9VD9Q7uHaEolKWg3BKuA+9rxNDp6
rj1e9UfCypmnazYPO4oCL5JaPP8L1z9eYXgaguSAQej/Gtf7TXCq72ZWoCLh
ltZCIpVTmhTM8IgGVsK0dhTSFzrgRRtiayoo7PcVBaXZ2wHE0C67IZWEzpHN
pMHk0ijecOPVMfi80XAndKAgIyT6wv466PSq1gskdh4W587U1qBHgX0L+tDs
OjTR+SZ1rZgYDhndAai6xOCpnNeO79jMt8TFuRjvQ+grC8vUFg3WX1wF6pz2
DROqW/ex+XsolJgOEKkNExQqcwH1uiZgXkx3s0lhntZNWS1zDQcVkMjLxhGd
wD68gZz3IjhjHBLWawBviAl/sk0glsVwI+3gCQEr80yXDsSrqmAjHS2AWIrS
NLH7Yplc4yY+LgyYZP2HsA0A027x9fa32CjTENLeHq6A+XCjzgLXvO5OwG3F
1okueb5RHseU5vHQiNEzg8iXxcjwxIQhAea7bmNIomR9txVB02YIcftc8Af/
j5+QsaEA0h2u2swviS6jkvjXSyjo3WPWNXeyWNsXNyrfJR+sca/OLcAqQtUm
i+f+vhYnyYWIWQfbMxs8myGwCaYz37WGFEqrtB03yfMBVxXx6eLK/GCQ3bjC
zvB5+ovmsAwQ4Gw16Kez8xtrLEPtnA7FU7hC7GW2Irb1wPe2ldsjSas+wA7Y
QtEsNRqiYXPEfV9MZSkK7dP7EzY7X9DV89P7eYbr+zR3AV656wF3eL7WGWci
z+My0VUoV9bJvkUiCk89mHcbE4B7xw5VoIBS0E3EhRmOWvhQZrn9OJ7yxBb/
mK412N+B49ewa13m0wIEkKYMoFRDxPZXS3o6SxHeeA+dmPM3X7m+i2ze5BL7
xPXSzv5OXYaiaJAwxEMAnMg1S851Sw8376nMwCkJQa0YDrLkHZy6eBJGkg5v
fp+FBg+CPyQYLvGdv0QVFIMPbAzOYbykccam8eZFma3ZCQ8ac9MCkmPm2T1A
4YNrgFWnYtqmXn8PuqOsJ6QfS5m2hpiPwkMvPd/GIO0/GWjFHKOzDtxENfQF
+cTF69wJ4I+gyd3mHA5hz1nxt1eh+F2lCo/r/O56Ph+Zamb8trhWFy4KvV0V
cwuMqjZGkm1AXO/RbwIt3bl8mAVIVosXSvJHY8T9tI2nT5UitzkS3/n7xBo2
CbeeQ0oj1L/PmetV7jXyOvmONqaIUEqIDH6vnSz8iNsx0Q6/nh1q79NW0FK3
nZPuBzRZcIzrBYlIqb8U7ZwWmlAI0VgTDUQm8AR8Pm5L5CZvP3TxGrP0zZba
9+7zgEqKAUh26s/LrKC2WcfEz8inQjkMk47YtR99c/5GFaHggTnlaj5NOJpV
0CbgJGQ4hljnP8yBoicz8ubfttNQ4lWtgzF8uFGNlIrEqCLia7iyFlgwCeJo
q5WpWSbf6YITPUhVZhCVwdV4zU2Wkk9vw9OZLBemtNDugvu46CgaC8BY4Uis
PAUMicNVSzjoLpbkMLbnhwIFHmfHDx6vM64lS3MF7wn4NrfBG0r8OT3h13bf
FHZiY6pvCtUIGkgkTw7cP4dcqG43FewZD2wNMLqn/k9BLxYohfxJhS4gwsbt
T0hq6DJx+/a/JeZTcEKyk4GOhst0eJAMz4m+OFN5jOJGGP9j8XITwnrP1bpl
2rp0mvJ79VOa1tFs3+AZhc+xEDFQnSNbGq6yJuh7QhwI9ifW7peTq1p3SXQy
h95Jzs2Aff/dbJvbqZazTj3bkpzToWy5kw2EXoTbYeM4fh/8fjouUFsyC3E2
vzRFA0Hn9lB/p6gN9Uqxvw9xNAl6UegEnapxuZM+7E7f2Xx3pdUJucUev1CG
rojBR0LpVJv2A9F9S+voaU1RY03iMwh1wcPK47IlvzAnY1gaqPlO4MBEQQXV
XrkCCamofXS+8xXtygtPcrP15u8lZ3xNzzC/TQEmLRaDvYLKQqUcnKl35XaW
BNDP9Ba5zHrezLqGXlGsQXoQNAdWg/JPidt2rN1NAbOGsmiwRL0jEtwTaLSC
6EyVdXsZBrvdZvX90L5ULUBM94JPdJlxDB1H1Q3DevTyljfoAbNWG3cH5uLj
82UUKS6KEAjszBvwwcQVUKwcZYjsutEUqFd29+qugdcNC63oLakRnUoCWsx/
IRews3KRELJYug/m5cSjhqTbaMg3Y0vTG9qzBy/gUVgsoIzCi7mOGBkCd/L3
fH2u34+yzdCjBnZlMaXY7YzJQAH33E/zyB8z8k3ueQdCj+KRrrLphQ6IvfaC
6EbEJ0JzS2WJ567xfpeuyUztylOFncgz/KOvp55Tk1FObZ1rODQVg7oZuG4s
xHL+Kj4CSugrNbXv6cYEDJpzSOR0zY+GC4rT7WPQJz+V9NG94ES59705GugB
CsWxufv75VafzD4RbLQRTpXsHDojEgeURo3h+vj94vno2dKONnG+mhJHDkeG
Dt5uuA3QlKRsS58fj8ouK8B3KOCLwLqd0Uv4CaIwGQ30nugUrEdoTUJQDH9x
5ejweRjMcfDtBvzf5K5F+m7yB7yMVOC3W4hzU7Qo8QT1+50xgywOBfceKrRR
OAad+i68Y/Yg0Y0UcZIJmYpOatPtKKaXk5LezE8mxV9/rDTc1OepVq/T9M7l
WnSTKPEKillAZ1JncPnOnJcqV5wWhSq68Y/bXEyitH9KWFShjBBeVSPhmwLU
VJnQIjh8m4c/hSGOkJZe4Tbv5V4+kwJTdA6wQaLJ2f45gwnkcixJPUAn6uuZ
oD2nj+vudMm+DdxarvGOsGZwqUSIlRLCEq3DjnvWY2KI4/jeSmgsxscxdBGd
RDkEaeThjvYMDrAF7GlumqsC5QNdmE13vaXxMj94oGlLgN41xW6PjLBoBZPf
++QC2vo3HXEvbTEUEiXjkp+zMww8q2If9g5gFB0PSGAXMJdpK1Hd8CJplT4T
ZcmiG6ABf8wZGMVmGtcZLqJYoRe9BPSqZDJ9FejphSXsQa32Sawb1lr6z6OI
Wij91tvLuvr21CVwtfMH65+Ck6hQ3lPi2Tto+XQu+PQV3TNoq9FyvpOjZeYr
dfIEwvv4DtUXehCG9zo5VYlS64sVyM3TgOdlaygfPy7RpocLMYhWwFMdgwLP
c/e1JPStY0ONHjoauv9kGy5NBtfPY6MhahjOSDLyUeEmbCtWiFcF54+SpVsr
G3HvRAVSKbBDBZOd9PuixP2nDmX7x1wFzXJ+dDosAixJWmImLwx5v0NhyI7/
+YojhccMXsMeukbwWNrH7drpeonqmym2E6OoLpVpSVnwpSV5FAbEIELAkPyF
M2XdRWyyEs+7247Y5X1uVka3+lmC+M7fZlEl66dj3VXBD5QFg0Bo86VCP1AD
sBoKkw6YDqlWSwljJMQlc0IKwBUC2XIfrMwp5b8j9pamqImGr/EX6ukKxELq
meCljI6jiuMyCQvVu5NqlrNYUbCnwo/V49TfBO16j/nuUV0yk88Xviwo2gnM
TDOG+26hGPfxMv3eNviyFxp7wlFqxqbRRNxldkSREHWxIT9z8EeAarmFiSR1
wFSWEcK+68vIy8Y5vnepFoA9trxPR96Jle6EEyS/68owNwFEaCKjZhdo5+TL
zC4UbxraYJoDYnF51Tq78trIyf7LdRQoEbshFet2L6drdryukgkHP3Zg/iV4
7ZkJUnR3pAz8lkleJhayN/zh6jXKQBQ0lWNkbUMoj5WDcLXqCoggoDrnc/0t
flZ222hJDWyejvwxDp9tupEtELmOLIq2bLs+bie+g9kZOzQQCW+JGhVmR8Wq
15uy7vHVVH5+gZtYfVv7rArchg31Neek41k5yOvu05F7iPP7HiqyI7f0SIKI
TxTPnEnm98GpXxBFi3TpAWd5JAT+zPyifqt+lcQAGCs4B2vTfsRg85Ulj+O2
fwGq+aqyb+V5UIo7cqm5IuQba+BTfAGHIg/Ex0nsw1YgQ/9FKKp8dJ6RQT0q
jgin58DP+hGdpUZXglrNqU1nY5+abf1QAjWUzxLox/aWUkTUeiy2IBNKOu/u
94H0ua+0bHyQwebBi5/tGaIaCRTqIdTv8kALpeD1amppo+Jdjk5fnR1h04pY
xUfLnNIBOXGkeCf7EvB+3cfw1jxMDDU7cFXqP2BQHA6TWrSSUpRVShccXveQ
GPohtPZ3Vl46wGTdKrxKnjQbFi4kkI3GkHoDU36rr15VHwBPkwinnK8FMQQq
Yyu+CHRxI9h+GffXHUInSdgMTX3hw8R0+1IovBjNTT+cKeKtXXsmlfsERnKg
j0nn9PETAe6Bse+CqJ74RR4pf0M6MFd6x30zKG/vZJtkGL8E7/gMojRs3Jv+
ebPenlP5epvhOHGtBjTcqTCsVuO3tfYXKF5jS8IOutoiq2tHCjdupONIoLU1
SxATg5PJuMFxWplxcz8rV/lJxR0fHI48HRWT3fi9TT7JsUE0JSB+sIkROYnl
gkaQNM5qGBZgDGkhVvVrJMUArqMYMjBOwq9AYivEHVIdMoTpJNqTrwJWF/MY
I3KapNvxGhwBjJbE8KZA5sC3jQzf6MAM0RedUIffw9Cxj9odC85pSyITBdVP
OETG5Xz9n0Swv+Rxhgq3CUu23pe1glwVMaPBIWJ3g4Pxk0Qf8v8YsQdQalXK
0mtKLMq7JgRXQOcTa9ejgVD6ZbCIF5YWP/PGEBVoAYbwRrtWY0LI76tY8UMj
F4p2YHrVERi4XVP7x0CqEkhbhLlsMGOlMiCdoo9bYEcJkwGKu4pS4k3E7xuh
euJF8P1iWgwPOdqyxcaI+OsYnr4ycVg98yMJQjomsVxjEvZIMZc/wpfEO4BS
iqXnZK+/4X3Mjn3KvS7NSpqdqHMrp/CIpz8augOtx2tUPJLYr+BmGx2oQ3pU
VFPEsptbfZyaBe8b/5NSK2kcACgo8DwIMmXfcsh3iDKXljdwXffVVbCXDBSx
DgjHK2OzuFAeNMsu0M+EzIybm1TCsAl8EO1HSyevzrCqjMGhn/TW0d+8Sz4A
Y4BtA2dOlx93yPGSuk+kbjfoRz9zAUfOtv0KA4a1piKBQd++wUMZjuCV33fh
7DZdm7BUQhIvOiA8YplRfhUhfD0Vkv/6D1Oo5fENnWHF15CNxbnIZ/UVzVn5
5Vg+Emd2HMsmUKeuef7MZnppURjomTr0UA9f0k+6pLarOTz3XSXJIrjO3Nlh
nYCvJjh/tHZ5AEJNFlzYDgLT8TBSyWsnhRylzrGzoQgoqwjJxfxLanPObFAu
bC7nVpahSMd9kSM2a0A9j5xhOBc2nS246Zs2ywEroidIyREtczM9QFA+Vtdk
8sLV5vhJtee5K3v823XCA4gVTrHi5vQJt7iTcVd7JAJD/AHloWOK2mIJojOR
rqMT8QA4rXq+1kNPElShsKZty8CmjImvg4+b9suJGY0tjgO7Y3Ngypdpem5g
PGYBWQxH+9BDVFlXbg68GEwOp9T5Us8ZxJMjNbI42oNWATKczpYRXBOmCEgR
cv/1/oiEyneHfZUAwMUVmwKaFR1je96fBYwPw+BUvTGJAmjY9eYq+SWzzc17
5StdrGbJgJ7AGGgCRnJr0fdiMn9ipN+e7EOH9fB1YIZzu79D+xdpf6wsh0WN
wan/7ify7Dpa1KVklYh+PuX3Fcumxu2HSPGFkIlyMC3I7wZJKW0aJV0r/tZI
R+2UBamTh1vZx12FU/jMAy/7LevNzL7QwHiDpuHrd5YAu2DAdBwxeZ3wUhfV
mQ1nlD8lICHMGpjOz0CuVmMACa9KIgPJgrqk3S/9jXaWTheBiFIKbhSHza4d
HILWG5UEQOY9XVKuHKv6rzFv9oC1DK0Iz01Ja58ljySwOPrEHAuz+LNdg3B4
2RMe5Ga+pbl1aNWFY79kF1IlGSK0aq6ffRGaOC20voDsQh0ZOx3F0WzKRLZu
sw6eZgnei1p2uhaT+/JmZKcpdYp9oTQtciDQqos/Gpfg5AIt5fM6+8olEXZB
x5A3KWLecQ0VYqoGlxNsUn0a5exUcHY1DIuJSJKJIixAN2ObXX2l0q0UhwfE
beAw5YH2jGclerWQsgLXqrm34pz3vQpBmE46q/H+1Tim22qzw2CbI2Rimr7l
VQqP6Ivy5pEOuavEKIST8JhyS/ntTyoSryOyJKLMCm8+xEYNoHjYfeAt/KQ+
14s3YngQS/R/w3NEkhDEjgem+YSQzPDSinHZi1LFeqNyh0Zw2vInBCAv7U5r
VC3k8LpUa+BExVt6wTB2C2hbE0jGAjFTW7ZV7TLUZDsp1TgKJBSrmKTEqdon
aCO1RNPubgfLOeTs2jKDBi8WBIgttkH82KUnqrgVoXcXy5oylCTZxJ3IadVD
UGNqlHSOSqbmyQlW2FO9MKVPo0QxY3X3mwQ/qnkdABTsWz5HW8bCC02uvIMZ
/f/EEBk1fnOqRVI7+7TzUCImVWsqdfQ8efbFGWKT1tgARSEVaDJwTnmuhk1Y
yUIp9Q++hx7ZHVCUpoIZ2x1CQLCmQ8p6QvU4UtpTrs7IVLvcO+xcxC413rAG
IgPUaRe5AKp/HgUUA9K6VmaS4sfgycc1sX+5gp1FZhexK+Mpf+XXNUBIIkeA
Rdpd5IShdLzmmqfD6z1Iryy0Z62Q2W5CSukR6Nmdt5w4bpFplLY+1ok8vJ8y
uz89GB+OPzKOgBUmzmtO/Fd5qoXBVIMPf+Kd+Yf60lvFiodQ1RNnl4rzbMvR
u1pi/EQjhtQ+2j07NQ58nBrtqxyH49lSerLDZR9LfYjOXDUplBY9KA+01Six
TlVPxb/H4Y5cHOTNIdm0buuH1bvuLMraBG1KCGq8lrcoVH/dTxboTuX2RFbw
HXhGWcc1ipmCnv03xnRkDfQ16b9dblMq0UHcYjTeMfcU3I5BaS6/QQGT1Lva
nRp6BHYLuwkBZIlayTe7U8UE3cF40wyn3xL0c3W5bqPvUW1/MIZai+GzAhWs
zgdNJWEbsy9mekRknbYrR5dttU+O6ulaamS88aU0bQecAwihkr2akiprSGSF
0Cg07sKXtxrznxcK39GlzUu0vYOLGtWAP8L8pPbbOZspqBM5S8y5QYf9hrgk
S87RScf3v+GnfDQAkWVrwACmuyB2NExJJUbWT7qwC2Qcm8WHEhuYbhGpMP8C
Ii/2gd3xITi1hSSG5rNe3qoIydiE+8uIYtqXk1Qv/nJaUfVrTt4IVtv63a9l
gfZiEgWNFnKqMisvmRmC1EZ38bxhmxY5BFg5LHzEHMOg2kAYTBL8MliNOrHA
6fNzwp/curHz94liG9/KQeQkGcBpWZ1N2wsMKzQvJ6EISU7H9B8oOaQvnsx8
4e/658B/HmpoW7ESxWJ7bYuENO4ZrQhPZdBs1R2iqNzfR0hz8u5ctudFW7Cs
ZDID3E4l1rjcXesD2WLU7lWCLFN61OuCA2V8fYta21gcRvy8gizlQlsQfVZV
NGnCQVwBYh4E6wkuUCXwS4gBYekAEXsCW+7x7m2pU3zLXJda4cwsnBMTZUQf
fnjWZZ+0bk0hUwXI+YOrUO3iVCb+eZGX54XUe0gvMTiZKaaxOvVNcYCqFsW4
XB+qw/2WfZRDkvHm15Ek3kBiv1ajbAOpHBtM2hB1RTvboZVs5TgCLfWTeEFO
6O8T+7aWZnFFH0qzNG2zmURbD91NBe/Pchavm/J2ZeiNwvYln+vx6a3PuGzz
SNexlvJKSuVZHcs8nmL3DwLBZ+u4DqJTEwJY1oZh8H1UkyZmvtzQbwhKhbS9
QbZ40kVEeKuHCLTe10cLyb8z5UTvWuajBRSoUjv/+eloKFqle1NXs2Ge+UM3
agZTXvguEu92d0njlEu1j5a7xOi2uII+BEAQwuXzw5Ix1bwPzZ5BF15CtfLW
W+RvOgCKZo0idmERxLYP+aXEo62jvelQU0VKH1SftaFXwEcYgKVYIqN+SEwu
VYTtxgL1PeUmwQllfH9ntDGNx96jARFMPZPt5QjagRtEOD4WGbY/FV45SvR0
NGIR6ApGx1i8kvtQr4KlhSAXpznorMRyGA7fokrORCJaN4DEzu15OltTy6Sl
pJ+in05qE9vjUs22diAKJefMEblGYGvkhz3DB3D3JBxjyx+Gpnx2fYXbF3kh
peCXTO2vxNpkai02R5tB7GFnG4Z8h4Dc7cfjkcM4nY6q5XSDYaJtSQWWWZwU
hFz1Hl//HrRcZu98gO6B/6qVy2/Xgl1Uf8J8NpvKXFqlGQHxDyD7EHYS5527
0yXWsflYvw7EzMX2zkuLn5DEhAh2TH04keUsxSRGeTM+GJ6MOO6oSmjN7kju
nYycxwV4jEraiZ3htbiJ7VtXqnPmjZC0KvktgP1l/ersjFV3psFLCDR9MDK7
gG8gS/6LPNcSWJHwbgiVL4aIM7vLxnFjP/ap/0pLHX1EpP8JYa2FFq6lnmDy
DgZdzf0xTwqg0SJXSFnrXb6q+HGcf4jvUhrxGqc5+7OwsZyMCtLy9CdeU/WJ
A5klJDWq1SEVXZiA9iiCfUmm9pUDYXZfKGmFSZRZUaS16cuAsAm8wkm4he74
Xp+1Dkpa7Hyq0lLlkOn2pPlbSKw3oFxPzSXLS7SD3wUFVL9H7qMbEDZlfSDl
QIKlWhs9So3WIEXpBBWiSPtIeQYw9Ayeut1y3HiVO8ums6ao8vtzAg6tqPYJ
5khbXbYPwnKvjwmoPgSfvVlC89QVeyaJ1AmngYO2pnLNIsoVsvU0lS2LzKAH
BSO7xxCqKmxZnoVdD+fh1dlTE1Bb1eAmhTnBsPgWcwTALqjQHi4OqGwRVwiR
JCr6tWSmsOaLr6XOGLaBFpQmysLhJ+V/nkRmRNqfNyf3ExlXrEkPvAI6QJ7J
gZOK8yUmwHMo7JFSEUspkHof6nAcEVIKd1wVbJmaWHjIpydV07T/GcwGZwgY
yjYRJ8xxdlqHWPlXStHT8b96b3SxG6Cm8tdDXnzpz4F+ljtRK2vk8hUmASy2
D5KUe8b7k1QF4sum13nkoU8L5JeeqATsNhphrSI8VO9omwnV1+ppNRoAaOnH
Jk2r14BIXmVLtqILqTfWu1psT227deczbyc0+3NaFwAtTt5ikX/9YIo2czAN
BLovuGcIYa2snahjk/o+ncg3ZWexpXvqGZHjqls90BSF62hOweMxG20Rg56f
+2TLwdCZcWIE7JV0V2zuh002KcYC+BgmsTG/wn1d1B+u+zEZqYs/PvAJ90qS
kZibdfdTcDYr0Rft+u9lzUJWS7G9McJCZOvG1kX91rLKwPcotVcUIO9pfizm
Es2FH3qYyv2dQcj9gwxM7XnqctJ0YEyDbQLvfyr8nxfadjATzfr+vbiaaicb
V4GNTskxtX9fipUJGx5YdYvmMvlTtWVePeGZ9DvYH63S2mqPhbi5GcwWFC0v
WTDi1ciAWMrJLES+jzz+n4jXScyjV8aOeSsgiaZcmfbzsgy5IwKs7kr4xZH3
EOVuwvHzZr5sTLE4VrprAtXbIXOff6hig7J1iugkk/xlMqd8jhYMmaMbT8uq
0brU0lnTIpykQ8o4ARfFnsW/ekRSNfArF2TZnNjek3mwK85Ck79btrdJx20h
JiIFgyxZl1iFMZ1xcwQXs9Oy/1aXnQ4pKDQkqezT+hQO1aQf1Dk//PAcCDVJ
Vs5nEoUS1eA/S3xOiju8wdbuGN3+4t8sblYcqTYwUOrsMe8eTAo6sgf7Gf5i
c21htf9eLgxsHzoYoJ77ANyITL9AJ1f84CTQK+vZqTAfz7aSsRs099Y3G9Rs
/5jhRP0KnAkmR8fCCfFHQ1crQXrcrW3Dpyp2l3ecE04rkANSOkqlLgqCVaYk
/QoJN1LujONM/Wx2bOWJIoWCiTnSXlazpvHmElLrFFRoJxUyAjmd0ee+QL9l
Rj7UMebbWBQFV4AYT/ssfPP2fpIHel0mtFW9TwAuyLvIcp5T5cCSAOpvhdkx
uReuU9bekDhd6FVviHru7ItgQ5bq0tWidaI8pDswTsWxl4Oj6pJG3Z2xjGUB
lpbDTjeZPAlpabJmeeY3zXZygVvAMCLqvd/Qc2cdaIKxY0Ovyi2S2HcoUVtq
RiG0c6noFQHmtmBDRnU5LbB0NmthrN8d1FNUi5EMi/5r+qNGrFKwRWEyKY1y
QOq+fAJb5fHbg5mymHuDtB2fx9q3IZPGgxR3XhhufLp4SRSvGvgtboKyexiR
OXrPWH5tKCPwCQgj9f8/5uYAlOFaOHgYY/BAW2k9TBLHyzDZX0JGOqmsbxFV
dn7k2tnqdRoBhwxutIqJhK0idsKmPRkO9WWx2yVN3gHlP6zCnCUS/SgggJO3
KtMpMgq/9ZH8bKBDoDv3e55U0z5gHTjJrzryYHixzXS8ro2vVncgLiCfPS9T
q634TXEhtcPQ+hyDRI0fua4jBoWLFjS6S3BV71eZoj3IgRlPs8cQldCKiDhH
aJ300hVxKM1ZWXFWsRU9JyxkbYUpuzTXNiFN3RHDKbi0kdy5Bys7cgoejvVF
8LXjVC8P8iJon4qtFn8KAnF1ZjLxaiNLomMq9w6e0yRenXpPPqja1B32imP/
vgIjfaZT0blbED2X0SAKJhkS/9K9wQov6LTn9UYQVuPZjpjuf8Jp1IeUaIPY
DRzCsaAvp7ph0kXBHxhFL6Ef32vhqnNXvcEdOiHPTtHZcOXAJS22VjEvyHBc
jsDzmmeL6Rdf8he9kQeF0gL6483u1QPFIr9k7kLT7yXpT3B841dRMR1zbCol
Ch0oGJUL3OWhd4i7TV6IaxdNxQUjSm7gsxz0p1b0CoVf11C4Tl5mSNOKG2hQ
F3UeTQ7AoBX5nUdzySEbKsw7DOdYkqJdBJ9j8CwLgrmVZ1X9Qs487McUd9GT
aJONg0obQZaXeEfFFrhfdwgvopXCHFVCLG2qRsCAxxvKakpdrb1RrCDlptc/
mSk29PRjj/VetW3B74mdMNZ7jE+1CXJiya91TNUtnSmn5RzUGnzCy4ZAi8XE
b0gyoQKIlijENyfrKZrR0M9bjiaz8JAfdikezrmJsz9U5CY3v09qvnyDh4WK
OXkoCFXvMhFbGlBIsz66hDWD0JVPyn7rpb7I8FXH8InMVCF+SMrpXV7LClW7
vSPwPzqJRwgGgupuy48cm5AIt+dwwvXsy/OxNK8bqI3KknyUGxaA/3KFZy2D
B0sQKaE14vIUMJTebXiNkpCQgGxdGG8Bsbp2rTJ2LrFwv7uQj7glYsqOl3qJ
w0x29JozjXC52fVId3su5GgrcTrBOSiWQr6Zj/AQv0TdqGEjEzMfMfZkn4Vj
2PP7jN0QnYA84DNtX3GUixPSJFxJCBBcxQXQ42TT1VMZ3HBvHX0VbCT3Gfh2
ndTPWmyKoTtAmBdXUPVfgNvCPTSNIDnW94odAGDqFtBgtOHO4nZ0I7riVhqR
xiH+dWqC7CZBgXH6u9PZlZpu2j8DrUr4S7VTi7CmDiaM6VQycAeaB7Oqbg76
cG2r/vAbM37vxNzQ399VphXEte/u4yIDBK+CROIXMVQPwSrcNiCmNcjyb3y7
/pP+EIqSqak1MkGF+fY323sp7v81IOHJeJBMaGaqmOfc2x+P08mz+TL6E8qP
6BXx6lT+DofQXkIobTPwAjg/zTrGXGXZszFsgJlKjHay4oj/ZG8wFbua0AXC
b1RaylpK07QccJnkTsGlgxcjBWfn24TsUnabuRAbKW7HHA64Rb3iORFDvjgC
wHmWtV/jj/XLids/9LzkneQErgnql01+Bcpmxu99T8Iu1fDbA0QemFeoVHHn
5AjHW5C1FuD3SbQugj5xJQnfHVihRT/uHB3xzvUGRnPJ2BRRabXQmh/GQPAJ
Up57h7C/8K7NV7G6C5XuPDSU/iHM9uSG6qOAogaWY0Jpom+mCFjkiJEkJSyk
AX0bbXR+HLEA0vU2CnA4PGzbNG4jn5P6QGvpR3oBR7TsrwoicA/U/KDl6Jgs
8V52Dy2WejSH/bXz0/joiml0+T57N+UjFBAmR0SOEYVPOijsks+Itl/3Dbf2
PFvP3OG63t/O7xkbfxcKnuoFDs64td5jhxwX0k+7l44jcY6CZcMd1q36RNJH
UEIfmKdUaLe7gEhAC1WFpgEuLdH7Wo9yj7BfMGosV7cZjyclyNzQTP/kTdF5
YxB5PXQ7BmLwhEOPUvGzaoGBXGyQCBHZhQ3zCX1Xn9igV96YA3zH+JQn50tH
Dyq0FYdhaiOGXNGGBnTRiF5Sr5/pLjIe64lKTf2jUjprVkZNGR9VwWhjLuEB
jEx/hVdO96qvfQf54vEeu6kulosTz0PEvscmhrc72ZiY8HfjNKE1xET5U0Bl
m/T/dvjyenJWDcCLFNVhwmYMGCkIzwyOoj8rtfFnfslnHn7D+e0j0s9TkK3O
qwV+WwYrpxDhgszmsn5UGKkeY0cfBwJsJFXkQka++DrdaqyBUhjDgpuRLxJo
IoFKP17hbnpQa5ok1McudOwgv0B1yCfGe8KQ3R9VFDRXE4p7zU1Osr937Cqw
bmbbNy0EYswbE5EOij+u7Msf5v97d0x7dboCLzQWlVKm+aiWMUjhakrOyQAi
q8Tq2BhHNWeC9nYmklo3boKo6BMjRiDETja9EqtFiG6wIlpjSeteFKxb+LPg
4niA/RcOmIEzZRn5uTAqHuIIbDok3rCPoqZfVLRN8LioZhbM9Ltur20QP7PG
0l4y9k+pqp3+8scmEHGPU+q53JV9/+D6XoCZ9E3lz3CyS4Eiy+dqnV53OHgQ
LPfL447uF8l2vsSYU2URaxekQpBhNWO17tZe/nXzR7glpv71GYJmrwNseiMN
m01WxbgkD0MsfxsBPjmqRZ+Olcb9OsOMQQYTtZY85Z2oiGCiDzN6OmksWhbc
J7d5D6Ibo0RppaYBvy6ql/zi6dtw9U4XSvaqRK9jL21Tb1VCQPUs0334A6wF
e0V/XIegn0uXuGeyALFzxCbqRZVgisxWuicHYtb0sWTR6sKJ7UZUYjCmVOSX
cbpFPTOtzTlELv20OTXC1GITDAdbQqo3FxxlJnEh6nc5j0f+ttIMcGQ0g/Hn
CfQYDvOmv8BOo1keqtJ5VpoRdW1VNx7QRcQQb4jRJvom0Ll+EZQBCToafZ8x
RsG1dDR+lnGUlCjlVLhwbZXcq7/eiMDS+E+5grJwY3KjNQbPqiDuRmvSh4FI
OtOSwJs6eShedxYiYg2wr8XBW2HVGT0K3QLLWxCAq58zd3W9M1wKCdLy1wuX
Fm3zBUUvyeXdrT/2bRrnj8iOUPk1/A2fu5bs5OBPQKZSFpRwW9dsiCc0xTBe
qmUP1k7wR7Gr1Ly8Ea1JLXzGyxk5Yrru6vuSFvX2Sd53hAU7yMFxBa/qhD43
A8byVhsoWBJH6jnEwiyVq616YyhfyOsxYncg1D/vNa/jZRgnSFXPJe8HssWY
0OWf8vYQ+G9Wd3eBc+CmuY/f1eRsKcH7RGYtLCO/hx9ORf47RjA3nTE40EqA
5nSIZrVcETosB0h0Rc02ZEbH9Vl+nlst6B/Di9D2fGt4zFzD5JaCblRkaZkf
MAlqvtXHj54hN9ndK/ihSVUrotmoicP6dnzsfsv/Pza7IFEtZiRcq3V+DOIU
kezQgdYhEEF8VCot6dEhqaps4vH70kpCINBmM1O4Gi5oJQ9RvID3VA15A7bs
6I/HWHeYJexT26VQTNHaSDmNGKG+4EKE+C8j5/GguuQkv8rHnk2HAJ2MzC5Z
uw1uXnYPRZsOeBieltz9ZtC30KudtZoEkNS+RnNge/RnxZmE5xvpPAqNj/jp
5tlcf7O3w6h6XlEh/NrOqx0+BKj2fwrPo6nR+0ohiPod6yLiQHbI9ldbi3Ub
eE9a5+w84h48vPD9nIZsbwKhI57MGgyCcyjdqJ/AKcTzFHuVVs2lkAbxhtWM
w27dE8/LmDA0BVi7F7Aw2eMiXlB81MYxbEa/yM4dxUaAfv4U3LZ5Fio3R9e8
QdVDp6joeOaED2RJtR6u5D3Qdr91V5cKSxYaWKULrvfd6Q6BxmRecqm0qJ1U
kMf6weu0tirtOk6earxpE33VL4haCxIAybm54IbgN6CdtxrwK7vyyvvzn9PF
7EtjM0MbQOJZifkg3TbitDFw5wqh5UPq8rIEmw7qQpVsxoErKMunnEKLjYlA
nuqm5vqW+V17YMhgmuLn2v4n+w7Ffjs5diVHYBlZrMDMCiJY2aVgbwT8i7Cv
NL3Yo1Go7//rhzkR8eAwkxyfYVuM+9n0q29SYo9n0uotiHu5rnxuv2f0xL8o
bA8ah3zQ+9F9wGPAa5DjKBB2s2dZFr32vuEOkgWfJBMsWsAO6ZgOWLxFtIFa
MimTGQ9NYAKXAy2ZrQpn1xszw4UmTxd71bxahgta+Zc23HJJl93KhprZPAan
kTqnM1gNYlV6pVEuQZZOeonvWKixEKgon2r8ccQYH+hc2y67uoYpLoWlYwIG
icyvm+nzSfRxTlAxQH3jkuCfkzcqQw3NgmpvAgWLbEqwL9GpDlOp0egCNahw
6eaVPphsODq75ccb+gr2q78h9dyOghCqtW1fdyAGIzdWjyxLP019kybo6qc5
OatZNFG5DKsLE1/1szrVjQl00BqbxVUCqspnHR4UZlbh1pDieLkJk4f2OZ7u
1uFBc6sCoc0quiF23iV/b9A7BN33WSyWJPPF9bh1vhGZSGMxEgRbjKhx43pe
NRjZ1HvbmVWIyTeu2Y9okPOc/ZM9MckS41Nnd4iTf+Z15zhx9hinBGWq9NIL
bdvHx0nEUnGZ1vw7dDKd29iplVfM0SBEZ/Ko6Y9etcSY5mWnbcmF/h6oOyFc
/HOxH+EzMLdVdHQ5YjCyFk+WF84mcTrO2Td5hDguZtlqgWbbxIi+MAbptSMW
w4ApESRcJD0h15KkMGeHWZYiGkgpZSdPguXmcSIu1g+4JUPDosUSt5esdX//
P11iHma2ZyMHgJnlAohokNHntL3YG8veWhW2IRmUndac9/BvD69xWv4D/0gV
KJaX9fr+7DDqO3RHLzoOC/qjjOeJaQrJEIHKyB34/OSVxVYMXJLayf324wHp
+DOlJ7z+42X7oYWZmyJBsk8MbFV03oLQTo/YLcqxdFkfLmI01oHSr+ILFyCa
Wt33DMZqCRbxRLYk6OM0uFf6zsIYUwlsO2XIFppxhdAgGWnpOfMr4FyErOFm
J5Z5oZW9Y35X0PVSipB2EB0IpSqH0nFCewGkXE1keN5fSOm6BbNz5xzy43/9
qLCghMxZogGpPc1A7bZZSAQAOEyMNUQLI+WCp7qq9Nw+JoSLVnKhdpDOqc8M
4MMeBy/AJRCgcLP7ENnjJebSLoIJ5FsRbcNxN+oa4oXibE72Pu9XbfUkIsVq
c3g/dp7cjz9u4K390nkaGJt/AbSMcJbIQUs4UBcJBCYE+gtfvIkx6XdTUrBS
NqJBqy1K6oWQXRlCl1UT6bTkVlPkUWHT14RtGd5/N+ojXk2LXb9nNztg3R5g
Hq9HFnOPZpkbKuMizSgyVISdjMXYPSrtqPjetYYFUjVKTN0bt3DWbWIGtWaF
yHPi8Y9+N3O9QCu/x6HUeZfoTrf8B9O//rtw156GQmcllOPK+NwgJqyG91vo
c8pbBRfovP5rXBTl6LarCXZWnHLij9pVyerDT31F84b2FgTX/DnYIoNT63gb
BgLhARxXrafXmh48SlWs0Rccjpalw92OOwWyoFT7edbu4iZKD0M/A2TgIxVO
Uakai92Jij2Yy9UEkydA26ghzl6xmv5fLg+L0yws7aTLcyb95Erw03UDHlXH
GjrW8zVjGxodpUMFiUc5ily33+/ISXsYhmZlK/iXU1Vc4L9tNyfXEGeirTH/
M3uk1vc8EAEslx7JPgQ83zWd2ceIwZAMRCkf4ykzk++FPYJ7uXyVklnnxUZp
Va+4DaNUvPG2/Wyxlm74K8EidtVuKRXnyBrH5HyCXXxouiL/CFrS5ij6WU61
Xjry4FW6tAs47ovWtyNmheRInZa9cvn7wNMQPFiT35SRFpVap+NA5a/qomR0
OZHtkM3r4FJk7IZ3PNuyoRPXy3cvdYXMfIZaRsqspeenXMh53qXGy4ICjhQw
HlZDAU4q25q3vrAd2B6L4Edt5qV92NBG1PO5DC6rDufNY0wlD4Jt0y0rnwJf
L5YCIBoEGMygeq71KUNzjhPNrjBk3ke60qrXz1RTiATVuNu8vI8lsALexKmr
qAzmf8Q8ANAGQoQtc0UYF9Oenqu97D51cuLeygRrR3hDnpcfwweRy4WlYU0T
A+mlU1zUQe2Qc8jQzQT3CVgYDAEQtz8+2iff6Q6CiNnrvr+Dp8glcCuuuWFF
bqY6tfT422CizolvcrO86rSUzMcsz543AKHMfOMq+MaUT3P2crzYRlcZn6Pc
oO7Zrkk3p1x65YLeXJPN5NrtJt09e9S0ujg16JtlFk53kIge+n/17ZWC5RY4
sgR8dG4PDIHp+STMhVxGjZVrNVjEg4F5uFeHenWyqYFfls+4SqzEtxp+pakt
1Q5+N+EEHi98Hl+P8iLuReX6IqB5jS89AVSDFt6KXNQ1N+s1+Cmoyzn0j5TZ
jK9Tf7Xtz3a9IlZCf18o6b6BshjfK11WlBIHDrKPO1JKLsfpabBnKO1+WIKJ
X/Rt2vTY6OubKQSb5JfRqC/C+m6W8DZORR/5j/REHzEq0yUgyS1QJ+pn80cZ
YDngMG1qSWTjwDxPIbxBkpJjZpixLkioXgALaEfK9THadj4zM3al9AVy9a72
iIpQi8hAkx+M2ux1nlvmXp0P3r4M22A8WV657H+mDL1e8jFOj3zp0jbS6Exn
HXDwigMUe4HXZ2ORI3YFj1YX8yiICVCVyd0mW1TgxU+hkuOtz18eyD48TRNg
2Dvd9hQtkZVWqGz2rRxf2DSEmrnNUToKBlgN+5iwE0SAQY7yxrsvcVpXr+LB
14GHtZWtuD6dZX0QVo6HGULw2LnjDz2uF1cwRa4cLB2mnhOPeqs8zzWIRwCe
x4efa0svpE9l1RWXCzKr4ruhcoxoRMsgqBBtZTof1CesdGXcEzdbCO+vakLm
11k8M1De+ANxuehMrAi4lieHeT3JkQVkZTMrQ/iH2e+I2iZewWqlUVb5nan1
cIxC8h0nhCUnj/ls1u9QF7Kie6+bnfUIiN4iIKseokxH0IGgYdb75t5E2Ghx
viXaqiOrZRGmn3A7lkG6LSYWzyxLq3bSy//NEoYpSYOJqpDbK+6kafpKsAxf
FZ7CY/5OLI9wqjM+dEtqwfF6MF4+/3WsNKJLvs0KpQSXdW+RwrvRBLZZSJY3
tG1hZycsADigpWi6jAfYuKMRsvj88t3vdJwxFHz3TgjteIwKF/yqi9y2Le5m
G9upr6G4zub6EdtI2gdhkQWI4slq6q+8sC62K1PGhHw0zQrK68FEcAz7me8V
ssQDosidOAPY3yWdvizuPH4EXDcHlTZBKf7MYodGqthuADmVB1YZvvlIkElb
XJJkZLG9QqZ/BHBMiF9n24ZYlau2ND/J7Mouo/JYshohLYqOXygKPT6qwTwY
NH2p7bY3jMTG8WaQRFfayHNM+hHeZCSBiX+YMjCh6/kEk/6KwEfyfVHEnuE6
9WPh6L/yevOSX6eOzC1SD1XKUuBrutIKxHFcI6uzDRlD6W9/Me9DRP5m5iZX
OeZkab9HMXBQmwyfhQLfdR/p4I7tcmkzNpRaBkA0NevjhK/+wjakZlVGTCQB
cKNUWZYw5EKCSz7HJBLwFTsFyy/WvGwH6BCWCrlARzL+3V8jmGwhJnwTNPOz
9+vqyDYZlhPHX7M88/Uh5Z/aEIcHn3HMZu9shkxBODRaNYYLSw8Qha/rKy0y
fQ4ffj9iQ0vImz2bzdcbQj6vt0LUqktwWg3asf3WtJXNfPAhumMPhfXtYwOP
L5F2QU1HfcA3ODIWM+eS1Nlst+jKkZuM6GVElC32n8ldVC9zTbONA8rMXvJu
MdyJ75NPSvOaCWI3AEUfe2PNt7rKDZfcNHLf5uWifwYaIN0jxLRU8j/ePVNY
DBa3woxeXIzslChRFckcQXN9ZBH3wmzuTCoeWKKrtdESbOvZPVXiETgjWCUp
jAbbqk6NzLKDPMbG7TTFh11uLJuduM17hrVaj0eEuBmDoTTq3A+nAyg1kowh
qL2g5S+mGMf9ly61t76f/AjVcg70riM8QXeW1Ofh/uf51psFPY4O0H22YI3v
FPoGEePJM24uoBj0byKufSmXQIloQ0eHam4k6Z0GvdVuTHIVs83Wc73FCWm5
4CtoUr/hdwjdO+kPTVheebjDK4v2uY6jI3Emj6MFBLFtTTBwXh0XejFMEM/L
ss22AMX3qsoNs4Tm/i7jiSU8wPbYXlAtxu602vGkP5FtSnsJuDuiaSlpnyB0
YfxX8h0b0YUZb23DVbFyKAHUNqIY5yc/yWwHadpwEXqbqfFDi6O2nHJghZoA
HfKB+nnzrEurSp1UfDNmHj+NywFa5inBsj9+Gr6GK3coCHRXxA4pEMv/WQEm
657S2fozaKx+ssGfj4v9bSQWOQ81LQILZcP7S42DKmBhXfTa6E5VTQs6Z1my
jkCs6dnRUfe1WFCJSzooqMmIHc74QWNGTrEowa9yTKImra+QIQtVoIiildpH
3dTOrDlNrsCDNYXQMl7QRNe/FDtfYdgZ4PT+xzZ9sDrlXxIMluIZfSPPNhFh
Ij9ViV7s2Nv5VPAmTyA+4a4LeyvW3eF573Gxe052v+FsMCWYVn7GQrd0upeT
B/XASHaFxyu392r4bpGddQvP97qyGPB5EsLOHsVoVNMOPxVKY0Q+0qYnPIwk
F2QdgmRbuAVNB/HGB7/w3zspIVy+Z62tscwhvdzKQJJV5To+XUuRFTXG+D7B
JkhtKOG5wuT2AbCniYm+Sca0dfkzyqupQzLHpm8jsguMqNwzOB2mJKqp/12l
EpLmKzDQ5VC8cYWYWnOtP35mQ2L5em8iLeUnVmeEpMZI+eTEvkfJ1LDclzZV
nlRuF1E/DJmyZuaiopdFZWYl1scJPSOuQjIGNVzLzixhzgaBlLpg3sIVcqwZ
fHUs3Lwj6Y8KHFFcMv5qTXTL5JrGO/n72Z9N3jEEB/2f8uA+1FkCHfl9Ema5
S1ptFcS4Hy5uP+hi5U0raIWqyubIkaoUUMLRDGW/K5uXpgmOpqfvqNKxt6pw
CcnMuO1rdx91ZL17s6oDwjGkL7bkEajX9uZo1BExPO42nJgsU1vq5ZrVwZKg
LhjYEZAGgy2Ia/8kurJHlvWPYur9jLrD1hrcISFKK2ZqXLD7VOZj5nMNALfp
Sa9hSdMrlniODHTB3sPWkk1avuS6eJrDw+uEJVk13dRLuEEI4rjqr0MaW23i
3D0WaHyqO23H4Ib+XV/WM4KPvvsr1ExjxHYqG0tUa3jXeC32niCCYL4o1+Is
Ll2tyGnLisRRTkDCODTPtReuhl1QIBaBE175sBvigi3CdRQY3N8PVgqEEniB
pUqovjcgZFzwNgVTAOdvUwRV/94hTnJSi0goC7lGeCa2FJHTkcTnctOfkJbP
idsL6lGjFerscx/obfvtEZ402gf5d+Cc/LBTKMSBogB9qpFoWF89BgfCQjnb
li1q2BO9FN9AQL7xBP13SnBkOAYZgng8ks/O7R3X5sQb1LEutaJfsAaLs+w0
ct+3a0aIAbPSwgXCl84yIEhq4YqjPgi+TStq9Ae2SR0Nbl7eGtbabMxhFtKO
k7btuZjk1qxE7aU3zeACVvU2Xzx5OqB0bFyahN1sqlDvtUluWmuScBVe2jqz
wyoTv7vqa/LfBu/4irfdD9bJBZcpnGC03wDjhzVOzzoT0nnM9EYH6KOvZKg6
lWf/7OyEg9CzzbUCwj23LK9Bdvkl+NJbq0P6xA/o/cvKSgfvQlwQdJ3hCRvg
yQKSYAp8wCCEbaaHgeULUBgAJsvyFChHUb4wIKVLjez7yPVgI/X0pbmbSPhE
y+wKE2HJbkNHcyLIxQnAA/LdW6a1vvE9r72fXLRljVR4asAtz74Y/sLudyuB
YrIT9scfF8hgUKiRrbbbg5IcXOkGvZXkYDfIKwAecdYMyelziHzbbpmobXo1
eabT5jAy5YpSK/2GQY4IcT9Y4xBuN5bjULUwKX2rEreMeIBWzFNKLTCwuoWG
F0g6RTGu9zwoOaNj0G4rtaQQGogQFyW6FpQmx2E+7R/sXroIwYTec4GNL1KD
HxYqzpy7b0HM1RRTnW0/qBIr1QBDnbei+9Z2kO3UVuF4/XMLycI2Sz1FyevB
TIjetG3GHajjsxnFzrK7Ccqug64dQtDxtrUwyGjMO0SxaZcBD70nVfIup6sZ
//AOAOEDaWtvsX4kWOHsuQn8Xg2ApcwCLQD5OQvl7JijfPxzFL+3FTDQ3j91
TAgsJ46l91h05N0QDw9bEkcaFYCUDlfLcs+raRkUBIwsDUMJ6ymC/OpraTy2
LmJlonjr1s2IrkZnSsQAszlMfYIRZmZiA+HpX/TBuScyrM7dDIN4/Lh3Pnmg
w1aQR5rrDBnM/8hMVK5tY64pLyUfSnXuJrjEsXCqFyAVYXjEyLbteURFj/3L
D+z0MzL9S3VvD1trNbkSGEKSWnGpOfP1ltxnJW2ju0zMSRY26BQ+k1Hop1nR
5XoK01ZGGjGvecWQyWt67xP0QnbpcNgAtPA3iIj4iUS3Kw/gwhwtKzc+r2yW
bRVupE4FXUAO9UliL2l53xycwnsnCvhLbLSpjsa7xrXJ/25RQ4pZcDdkYl9p
qe2YO1aXUUdfDj7oi1LlWaZmraxpn8q2GSdVLUGQsLSLynr+2ADvVhPvx/3D
mMEDaeB7WmRpEMDKHzerd490V16wb4lzqgg3Hjj740oktCe13GbNY2dRSxmE
rh9WCb6daVBXN3u9eEftGD551zhdOveYep8a4EAJ+qdKcYL2K+W+4zDq+H1z
ZufDDuK/pHetdi0Z7+84wGNeLYCFu0pqL5jGlhBeaNgQbju8h86s44QH/kor
O+fwrsVFBttxHarotFXVDZS+2xm3pMxAkFgw28QI1VC60214QWM+4BPg5w3u
vnkC1Vgbi9fcoVEGM1XYs5iND7hvHMdyBTgjIYWBJnyAI+S4qkVfEjdnIshM
CVpF2F2t1/k087Jxi1MOkjgu/NAdCsE1YPXnDb2ByWjs5ngGPh1w8O/+fzo5
o8/S0VSt5CXXrY0cH/Q5c3qEv61HlGV9KvVw7eiXJrzR4+p0wRnAyEms8qoF
71sI4vG4XmYVjqB/ZwpgACzHhqtQkkXxhKzBuDusYfTVSpEnxOIji1MARdWx
Bm5k6AgpUydJefpaVjtQ9kAo3FILX/VG748XMUbMWArgvRqYUb7wtcqoIFSj
jLYNEVpRh7kzNRTUHpyXT+J1D4h8nhGbhAK519Fp5yfjU2ru9TsUDy87xPkB
nqzhqHKYHz46jzx6Kn1SGHZZQYQfkVpE4qkib5cSLDu57CounxBLFD0/rdD5
pqHy+cOFcOzwWXbhAcbnn+l+iLLkzhZn+wv4iPEsgJLPbLArV4IF9v8/XulD
qH0gkb0BywFNUKGrMoj3ZS0KteOILHyDJiwux+MgjgcEUDSe5mnF42XJpKul
bYg9Es30BWi9smrnBkD/ZujA+tavUJsCkCcymBgTnPVwY2H/oNgVjnfkYXYH
e00LZq4hNW1UlvJ52GYXax24rSePx7l7vutABT9x00P5UA/yo98RQfuHuHcT
D0cR34FKIrkfbMoMoB1ckFraEA5f2UDro9ml7QCetGaR0jEgXro+ZdSlSEjY
auIp/JD/IB/uOAaJ0VHHFxDjlAuq5UjPKfNv8tBCuVUsq0Jl7FmpSq8s7VTp
59nzXWI529USGwUAbAdidcns8Xj9luvPjzPDe5c0CqFmHb06atBHXKdgBfiK
w7g4q4w/41gEnaRF5IMrJAgSdYCaH8R83hZmllOXV94vbKLKwasKEW/qwoY+
2EXA1aWXlM0TIdSLpb4whnyYeWGIXsSqh5VTaCDgXyIQKCF7xVTCbGuleeYG
zLVyk1TWPSI6DQT0kppwMxWfHKaI2Sk0nwLnhU74FkA+/Kz+alrpTePeVhHj
mkGC+rhK7F8gVE/djEzTiO6ijgEt/im897LDLaj+hv43DUNVX2Mpp4WrgJjE
mkUnmdQgw38yLA8Jm9kCCNJmIo4vHd2LR8rMiEThpEZl8A2nb6cXWrAAe/dQ
Dv9MKNdt/q5cX62hFGmO9XTi6qc9/gRJFxIOS/qUpUfXbmih1kJJ70ujve8S
Yg1H0FSouREoJunqMCMuVJ/LzY6N91DHdsFldI0tnZHz2K13NJdKKPy6ne5n
MMSvEmf9oKWYeh3REwYYzSt5S6klj8sMmF675d40WHDG3MS/onl84Hc5ZRPR
6PZh969MoSVgb7WIMzgJjzltlfP4HPjrovPbnJWgXflPAcKWclQknszGlyoq
mGwKYjQQre8AbKc/jXbUpAFouVZPp7qXtuLUyDou2btzxZgdAdLSU5yxssBW
FNiw/PSQ72greXSfLg8iGy+DUNW8qsT9qrjgsb6AGCjVJd2mlwCEokEbleI6
3Im26Ml1GBTB5fBB1SsYVnK7hI7KtV3OdFO3lct6q9xV0cfj3ZsNtAvL3fOO
J/OpcIJms+tnZ6lxOHUjE82eBdOXUp+npymtIGaNFBTc9QbCE0pU8Uu/5uwc
KTFu0fkBCsO03cFyWogPV6KL6E1anGKUnxyJVV5xC1i+twJ9HmcZXNcj3Ih6
uZtoM5AeM6VzN1j1g2mfTlxmrm6ig75LCJNNj5aPggSp5XAGmP/4Dlcetv4q
appHhdT3DkR7mzRDr+AUQ0KYNLtPMJGzQ3gQ/a3VBxXpqen/Y5EmdV6Cs29a
+5UswdAboAzp2uskWCJFGVpFx4AahZ/jvikcqC3YBPTZmYbMEd6iLealjNss
07G2LbGpWb48JziJ94v4NHkWJ+WB4teUNQRKUikwLWQo0bx3WZ9mQzR4+/eX
QIzhe1t19f6BlZQT8TEIwr77GOIPu5PoxwZoOa4ynK7lw+gfHXPXYb1odfJh
yomLP8pDck/nf406MnJIIMZGQGDlQ8SOa6mTrexgHDki0q9DDb9N5pntw+C9
LX+m3OoJqUBMUzVCKsi+XaI/B5tT0RdoYG7G9SBxQ3xJTYgbaqmlSaTG/dLg
K+INwEt36nFqIbQULhq8DjtjqZYzQS7r5PkUDQypMOZ1AipOVpvko4/FbTeY
yeJr8CSfafP4ONt+YfAVLLbIE8KGuXM2Z48S23yTB59H1Z+8PFPMyrwqAvlP
4AdgSQD3fiGdy0TKcPKrd50l9e9ms2mbnzHKFF9Qys8UfqNUKyopXT+CHvUz
qHXW2QMo5zwXiKVbZwwRYz9+UTwfJazx+VpGS/8J5QkQnB7ZN6UozzPM3EBD
3kWoAK/LPElUiG9QM4fYwecSemvOUQU8SHkkOAmdYHnZCnUOVAg6fTNNpKaM
k/3rbpcRM2YVwTOKB7VjjpBe4sMyaV4SXTEhXdbH0fAmEwnAmP4UZ5xFk6+y
7ikV6+u4LkDUwuVfNWwRrVjtiKpogEPM+2Vz9W3FS7ksgBhZ8XtBx/3xUWP8
LXEku4omLoTU09///2d/ys90icDl8a2VZq9moq/0F9yVWSayoFebstUNa6Af
95SaByqHnmlASv5sHGGr51FINCs6Yfr2K7/v0l8GDoNFKCfhlcnAejO9nDWN
DePDSH1yO8v0+Nx4CWmx4S5wjDtzW96jo7PRoP4FdmAS3RXpXHQfqu6jSadA
JnD4pa7yYTVUKkYIGuBJdTM8WGNtNsgU8LMsnAEPGjsjajoB++5rjsbmlm1b
9wUC0FiWEk4x3vYeulm080bpT4q4PjAkmkpZSAE3TJm5F5aZ6yXmqldu+5o2
dmb7sghEcpGao7EkQu8j0WmpoNWJ4lrks4HcHzlWAixwnelY5kebzj6wflbg
nU8YS8BVkSykVCFRHyjwq3k5uuJ3saVasXIuj0NcrWGQGvQT9eK6I09R0ChS
i9w6MvTKlWNcqh694Q7C5NnldzhFPJF/jpSMNRRhZy5DIvuaFhk39NU8vWMq
JRhJ0DxpzdUdiKol9RGBnMgoelispsRdoZuI8a7qGUuyuul3zFVwt/NtINsQ
/R54mXTH0smcH1acztsvz0uLwGTbDzCeuW4Zb/tblGwYqjLLhIS52d4ju0gx
B0EWzU+h2mFzQIK0HAll87unh/TNn88dLX+r6QiMX/16iXoCkwHut2jtazoj
7/LK/KZEOOVYmG5iHuac9D+Gxz6M2KiblWDqUonX1ZDRXvOV8NgXrrVOSdVK
1RpP3MRQAcwnXbDpuqMB4vZpNsTosZiS5/z55P2c4gIg6t1FwbBVfj6Pl4l3
W6kUQjdsspExOYW3nupIKNJ4Bayxww695bIqKdwryK95RCS12LDp/eNa+FX2
jAm96eJrHOJaBYM7Ao0rmI3yJ3bdc7VJexPMvPlEYkFHlDr3UsaHJ8ixk6C7
tNgvFaBTh1GEM36QrNOF/RtnKK+TBNBnxyjtHnMTAVZXHQ9UBl7bAKBzzsgl
tO2ILZFgrFgsh4ny+qCJCymDZzbRcL4bs2feYDyXS8ZKYwtJMxYYHbEzAkiE
NcnDPijlbnTHIZftuTFj5E7L/RyNSy0pi9viiHe+udL6VisfMTGKpFzOzZwF
EVWdD0eVciuePcIo1zfaxPYC+EdNK49+1nWMSIV3qSUXeMv98aAC+ja+F8Ch
f3QJIFLMiRN8+FGme7keYw0MlIu4fpRO/Q6p6LEJ80ah/wpiOOdqNDXiCsI0
79MR+kYLJELsa4HkvsHXjSNiCnZRklfcAdeQ4G0zA9ZsJizeVj3ErAJGdk4l
kbZKr1kvgoUKU0LGny1ck8p079qZXvuOWdtVMwl3sBtCI5CtLPtD0UBPQxjj
h8qPl35Kq6t+t1weGCUEU8BXkwKME9LWDKpl7vGA5WiKxwmZAQqbrvlYcng1
Szlw5qOOcDhGSZc58cTxDdf4P2Hv/dBfzQYd+KQvVKLyyo5kaJDcRn8YaFXD
zqszZMfZ7+pjZUUUNoPOAfD1Rh1BDWlEiWogf/k3o0di2lpFUoDOikuqTq+/
ppOnuRRxrfMDYB4NPZFTDnrWW7e43Fej+3fVVADYMG6bS6jpzGBa84fEDA1p
lcW1GE7UXFGrby+FP+cGc51IrEindlQ66uPslWEbFtBb0W4BBpk+/c5wib6v
jEi8WUsVFcyNduzjZ6Tosp2eqSp+SoPqcPl8ATS2IZh/22r51aAT0dKIQ+a8
9dINq1g43pcU7oOkJPNAXA3Aup6lxvv9K7EUIjvwEpevV5YCt0rAy3+oUVM2
2olr4o2hHZ+3HZVSZYd6/IPJKCS3gW+s8tJutKT/1b7Bkruo0hGv4K+nJ77U
4XqFsHLdLIJEAwF1sCzbuyNCcpS6nEhkmqwjFgdKVjPkgLjl1YgM9TKhmK8r
HUIAKAjusYhsjltGnGyLrDIrpOEpPbs77NTNpZnmQ8HE3YmtzjwNuD6Rfpcv
n3xqEEzBUPlNoqWGjUBAbBCvPYY6K9pQoZUV8q8+uE8FRRJ8iF0tOqutFcGL
Eryxgi1LnnbfzIVp+Ms8lBZiflIgpw2uBH8tqJiHdI1NmKaLnOm1mgRVR8LP
xMG31H7It6pCTrkryHBci5qDZ/9cq1hHX/1hCRhX2XnFrOIKojWah6Eica6X
duGPu/hZZqG4Qkt9z06YHBKuqOam/AdjUczyokwy0FTQ/n53lAppff+OlQI6
rnj+6f5DHGU8j+HT9hQdG/HiOpDJdNd1Ex5cTj5Bei2Fh9S6qfRuMhYZehA+
y+r6OqWIzlQ+RQ80EN1Nh9J/FTbr3G47g3zXdQPISy4rxIwMg53RjtwBgdRA
XzoqI3rsELSWVNi9oqYO+TLWtyIYCroiEoFwKAqrd/RXPoQOpiWMmfWqsZUr
D1NRqNuLHKDdDWBD4zNcIbwUqsD6djkpSdwbX5t4AQC6AHWBwO5erPrv8EMO
KzRl0SWT0e37CC/HUsqB0RuVth9KnErQ0crHsd2uIgXUJv3kGZKB39LoPmzN
o4OJftd5MLyYDj4gIvJT6Khu64GcrpP31wzltSGxBtQyFgtMzBBssnM79SbU
tJnYgU0wM74RNLUKWUNzZX2nhUC0Eib2Lclxvx3YCHAZQCQM+s1AjzAq+ySG
xmKNf7oS5gINnhpGm5SSGfEO2Om54nHjdFWdPAkrW7nBeKSs364QO7nJHp2l
5gqbEMnv6uySzgyQ6dMkPLTrxBS1v3URWwrRqBhuXx3uESFfas/i/MFtxHNh
NhshX+TIa2UcKJXZkBqVgX91WHC7n4FzvZuwMbe7mwVRGb7WM/vo8yeGc17x
PrjQm/gFA+/Mu/a8RDlH4u/tVHLHKl69GF/iFh9CdE98c3kGRm8hXvgToTZ0
PttiTXPeAxdUr2QwVtEmib7ZTYdSlx1RiwxbLzH/tTCaelPypNojlBmz6c9u
uaI83K4k2XiOwmPUc/4qZDJyTw1UugUi09e9txFm5AGZIupYLmtOQyic0API
7iAAMZKbNp5R08Q++7CifYPlT9qHQSUX1zATV0+mijYSUpvyhoE5p4KE1xOD
B7lwyMiWf9neW1F3cCl0ZU+mRwL5jJWzZk/T4uKgkEny4bbPxE0fq1hvH/yR
Y5mfSxO19bppam3w/7NpTlYoT43ge/nJlTrh167HnqQx5hU46fkb2J7sl25Z
mDr1T5Pvhy/9ju1S632jNNvxvcn/eFo4nGTxcNN6yC8crYombCuxzu3zao+B
QNO7q+iA4B+CQRXuU+EuJPhalW8QREp4D9L9AvX/ZsQu5N8ENvua8Mb8vzT2
22Zhqxzr8nrUSzzIpM6owkEtSTYDXE8HF6scgYZlBNAKsxx5y97l1UPkc3RP
DvDl3t+MHx+HL8ImhS1W3u2cq90iQ3aShfzZlHqFxxUuYhLK/3IcINbRU1rQ
UFTmbTu9sBXV0rLCZ1J9wM23ZexEjOkqxUkXHG3UcMVIvugqu0vSxGJeu2lS
mfu2ji9qv6vfhKurFxG2GMqYzSmnwGwphJQUFJ2Iwn/WOiAe2JiILfW0AYp/
n9nNprBj0wxKKrfoSUqQcclOldRyJSvbBF+E6AEnI2BrDHFUhut5Hmu/Vf+3
ckJNMbs2rhJRBQuIQsUlZ1U6glq3uTCawDbExtgMXKu0Xui4U9HqrkCPROqU
s/TlCFW6dM5E7AcPOxfVAhcGzYaCFvE7oGXH766OXK326QppLW6sjptrzWZR
ST7Tw+NX3gpcvcpmdTctqghdu+qrTPW8cx9Y8D/Zmt/hMV+vTX8J1Jcix01v
myed/+QlbnCB27LH9+OxBV7KBewDLiD3L6OeVMCrLSKDsfzPc6GFN9ZDhh0k
FSU2Er8KPSd6lYB392x19L0/PF1esAy3TpyQjLvvYXrWioXJZRAs5za6GPL3
oCpGDmCgV8DO7Vw0XOlt+rINPuxH7lzcaipTJHgP/XyCIAL6XDIvtmuI0Ms7
TXQKpst4c/AAJmSX0/R0MF9G2645MlcRQKgE+96+HVieQXvSYdIY4c4gnhVf
kUlHL6gp/QEZ+c1pGh3/hrvAbbWH7A/ICtMtBkvxRLM7mWGUEPFSVg9b7lxt
dm4cYx2PpFQN8qsrVqEae/SBHJmd5kPdNuQntyY1CBfbS6+Z7JoY93o+Eiwc
BmjaX/NARgop2omw1uv804TMD+B5GIBb8Sd+krgVmnXFLIrMTEx+6vgEnBmK
Ektugfoe/nXUAcJ53VyUN4zcoynxlJPqV167beFi03oQAoSK0Akaw5gaFz+0
I3prh8NE0Hwf7twEcScq8HAkVRbATojFLBeCIS9HNfjBDeMUZ99GoCLVnLsx
hTfFTBW5hHYPBHd/SX8WwbbeN+pJ69z2QC+WKNIA+Ea+NDQOV8mGyOyFZJzX
ki1+BkQPuDwWwb/eUZgkGr4YB9Eil952DTL/Tt3B3nq7wFMdXpJnPIxfd/f6
ouTP7c982B4cye/qJErRDQf8iWURofzQoHk0XoY4GoZAGhAs6o8WWVKn+rg0
h4QEzDY6/eum2BW6zUnyQfIgsEB1MHDG1dEeYnVxNWKsYQ1/9j5HoQTmMRT8
nFwvcM6WUCY5Ytq2y3CkF67SaC5oUy+8dSTzFsZep/wn7QpvgrRWTsg1KwQB
zXPNXF4hQcN2B4wNIGgujsDU1oW5vmp7XYSSbJo6jdPn46CumQ04hi9Axkq8
xKTd6fR9tPrB5PHerxLu5RLTQ9J76+g1OtNzI+Irq6q0gy9q7MNdOJH6DFwv
p1xGCxWfDmb5OD3wtobKK6di/afU6cpiktpOJb+yLXzdJUIU1bPqGSstDOHd
hcz5fcnTaGBGSacbdXX3ygMHNa7W7fDsoO+fkv17DDBAQCMrZZEr3VlaiS0O
+Lw2xyAI/cWvxSCYwfmJPZceoVvQk3Qiiql2BefFKf8gYldhciGITDu4cIqA
voDmmS5s5tuGkKC+pcs2B0Jxf9Vh6MU0hCDFG9m7mhB8O/qhEU6j8hwKit5i
GpTQRvN/6Lo9+zBQIalAvGOzniE1nOYE7sFuZTKxl8oppw9e17Eqbw4aM7C0
wt/JCryA27q4+PfEF85oesKB0JcX++L7WvgRBrRAeSIZEZ5zfEfhxKjV1Hvs
GRb2DopRU98S38OaQefoVIsyhEpBztftfV4nFmniY22SwX22rUg2mFFKbO7w
KOPTpV3T8pt/QRDrK4eiWRpIP4mlJn9o3pJ3SgqWBaDke5Ely6+U9ZkeEiHH
RfR2wTh6dQqZsY4fJ3r/yDCEiuNvUZ+TzbzKFFMDA3+9mP9Yc5+5yimvyzBy
omrUV+P/K2yeARodEfuf7UfbfEGN334f4t7H20n1xx/F9pkV39johfqhm5nh
s9vDTqlvdKLsljF03Q/iu8PAYbesJtNR4vbYpVslNzIltltXIoevy12FBi0W
icESf1MMWBvhT/w1pOLzFy0lQ5wwzWlzRs/KmYO45gbyxvnLGz/uaNC2MHKq
EiUgYpaqMpo1obeR8qsVp3sSxgETK8YJ8pAyQDZD8AKzSusyx/mZQUCJhC6i
VdBOk20J7csar+/gdBD6FcAAI5x5UqdtwT+TYMWcrbWTHg+HV6l9zbtdo/Tf
VhR0O51tOCQhAWYgI3Q1nXxsxamp4pC6S7E+WS+bBSi4NV6J7NEMQ/7PQWO3
Oiu1cNgdkzjMstkZh8ZXdCBZILxus0V65Wop+MkfK4jDz6JldolsDcG5l9Ek
itgFAuh7B38mpd6WmN4ah9T3rXfeY0F5g88lgtg86cvRFKEgi0ozGr3nfJ5W
QEIM57GEnhjUeO9dkRBcAHFm1TPmxR3j7Mt/2STsLu6kXk/7hvjstL0MP7Ov
682hViVubd/t1K4CDooPFXFvNLvOAC5NISneRUQFiYETDNYKJsRd7/HzgsUT
eaT13Vxoupn2vD7U5MdFUlie1LDYSaoOfiRtOOUyzjJEBEvLOPaHqtxL0hN4
tFEm2wh3z0tv64WsYMZqg3ur5m2HnWK5k4aqJnYWNr2viwGs4H2C082rnZto
T4LMfkm3xNGNPUIuDLMhPXRqh+9Pl5fFGuZ6l3fH3sQVQ90B0TaQvcdwWNdO
1mmrMUaywYNffnaTKPhRGQcolDeRXeBMRyZjk2y4LjkWsMcrf5j8fTQoetRN
DRlrUfBipd+Q4sF7jAgSEhypw3oy+wdG41ecmM+Dvt6FEyWJxKCr8hGprkSM
esWbhacTwTvLPtkq4eBrRXLAGqTZZrJrwjqAI7eU5UtdIB6PX7LMpOb01PmG
0I4coX+2aKmNkKfudRkWU+Jw8o/2a9D/RHAzrwWUPQrjO2EF8pSxdGXSG9m1
lvvRVGXUDVWu8jcfgdL6dLMVwaZosGxzPO25P250v3c3Y9u1qvMGxEZIUHrH
uJjFGqXuqkguXC32kcYDTWe7ExsH+gELQdNWOYkxrCviD05qp5/hrxOAQ//g
IP7RfjC1/h1/Q5dtIAvmJ2ondiJTxZknY+ZEmyxtUSnHTE9zhp4AkpKcFrFf
LjpnNfFz07/nGHtxGcY35gVqisy9Y5DZJaQEohlXJ34ilLOwAhAdwv6VV/hQ
cKckO5fHpPqlxXCU3YBcL+htMQ0yFlBw48qWkVsMcS3i8k/3p31Pc4XGexp1
/nwStgT1X+y/z8ouGmM+Hr7mMaQqv+TLQ1V/48DOW3SDr8p8bh8uXmmExPRM
eJbowjo4gs5UNDK46ZgiwmhHdLVQ928SipgfZMTExGF1AHNdRa0PTPotamCp
vtUi1VcBaJ3bWS01meaWKDeJgTKs2xdGRfpdDtZ6f3LIXmtz04NJRL3E9c0A
sre9lmXt7/wuXZABse4p0ukYYkejtI3VHIPoWiuRugHuRyiQm9CRWDNsE2OC
HB7O+K3Ccq0C6B6+RXiqaPSNI+VV6/3wFl2I/ReH9hecQ+Sojz/UNCiO+d7Y
ZPukyaxyFKbfXPf0+NWPsmm8xMsjhrOMEfK2jzJjs1LECiR/mD5v5xX6IWa9
hi6k9cOtH0t6osMhNPlotMNVCcLBZ5KpvZCmhVkcPLB/OVvB2QzE8V2rNE8g
IgGEL/vOIn5wIqN0G76Ytah7eES+xwAB5kj+9zi8Ebz/W0+hh3EfoRYgeqNe
e9cHeHsBDZiPmbVIxNGxmu3wNFqLE/YzaR8VG0Ng6q+xtzNPG0VIwvHbz8M2
IMlMgVgI74+63Mcf3SDY304BqbpZefbZdZ2UzvmxO6LAslV2bFHnHioFsQ7Z
sfyHNPTL9wy9TWBLcT/WKT5DPY9ee3HVb/sMLh+qgi+ulSXTzxa+eiN1MWqL
S2Bw76Rjkx3ZTKyOrjHd2LOusOqamREiWSaB8hdnVsLJgcRbTf5B4vmTTfrl
FxnyKrbaeSnGmWQRBKCpyehadrr4LmHceZ7UoEMQ8Fx8q3vUjJL0JRBQ7QZd
rVKNWXvqxXZNJMbVVpnHZTLoxwTnQ+NxoQhbD60oMDjeRQz6UkI9Ydu8/gPG
VRVXDDKDri8Z6ZlrhgS2JR7dECLf6Gtqojng4qXRzfQ0LsEjVEDbktQhlkRj
ToaKf8mQ76M0c9grLMzdAx602uDHnJ2Qe870KYj8uRb7JYLYK4pveh3bMkDB
z66OXN4DsjMj8ari3mPTd8mPZJXpCdcQdIS9KK/C20WrjaY/Tq0aipe7cA1n
pRYsbLYvevMZ5pAJ2UhUutQY3xOxybNvr6Ple7i/Cl2IldVramZiQlx/178z
mqUux7hRPezgh5wA/LEYyZyPg5Ta91zJXlXLfO4M7TA7y367ZTn3GChtCpSD
78Wbne9+2NDOAEKWoQmxYeIOfvgyiJk67n0aVm5o4l5wzEkjAy4VEC+axxui
N/4R+Cq/vYLm8OjSTPWU4NSzRtIaFvgBFvo4RRHo8mMMgFdNmTYCqudt/45k
zoiq7ZG4sH/YkckzJE3ne0Y51JJWw2/CuctOuWn5X7rEMVyKTbyojioBlKPv
WJPr6XUyKE7SmHwE0VomxmrA15nLgib0aYe4lrkOwQueJncpPt8U1PyGiBxG
bhnHefIdORbfnQWLcgMT1Aaun3lsn6k+BWmcnn0HxVAjx7uKIcSWa6UdE/Ji
5BEMHLGPY1EDSV/6TC1ZxJWxorGDlcaDMyoJi0IsFNQZQVsDHYFcGsGN+O3N
1r8/nKy2HShz3ZnUZlJ8LxZxhCBaoWQgnKEWa3qGficflrL0lZOBPV/h5jEe
NKus18YXnSdZnay5VnTLKQt+5Wruie9zGfocN5Ba37P23GDABIHh7odGylVW
2MpO1afuOfoRhkYlEEfQsMQGm1mqMHhTfIJJEcLDPga4IXavQb8493fGAJl3
sJy2ZPSiZoSSIgu5+Z2zS4ik8mnuC35W40ImLtOIpszOfbBF/ToHWf7ej58k
XBti7Tq0iMPwX2L4ql2SXDl1wTIuPnaaK6nq6DI3U3eDk73xl0JG6Z+f65Ty
Uzkw3aVkIkyMuAxiG/dJEFKqOhESJEsV2NPZyaEjZ2f2tU0XBwnIqQcI9TTO
9gnz627mqFXQVMZi+SiRooRiQ55Z7ZHLxBoSTF5MI/JX1GUzToxeqh+2Mke5
OroC22dK2CS88wayrDwCvhelyQzGa6KnhEmuOKsLQBLkkzcKhX8oukBI8Ibx
/cs3Rl3repgWU8CZPL3PLU3R4t+UYrSLeZQfRTLIx1LnGvTTEag668WbaXiH
n+P9NJyCrzCBJzLq5F7B/JLwsX4DNTVMI7FBv0Bd5JoREEevJhrvO0Q3a+aK
VIrvgIBr5uzmIUHtAZpufWaLLHaNk2n9POPF8LJD956XW5ijq48nRpa6FBUU
fktHkFjy1oHhskAW707BBFeCAwtMkmc42R2724ChoE9acplE0QsIhWCwh2hy
CeV+XJlwudfaXbSilm/mu1ufMvCr2paunuCdJPYnzXdrVY31UxMkJQQDZKTN
I9QAh1KVmHh8DACVDYcc39Itp3SyZH3CAKgG7ZP8+NJbYGRgs7tEmeWoxNf1
D4/j2kJj/J881TRNmqn5Zkq19fihPDk2edRKaHSTWgYXLyOaJOY3U5rHlRN5
U6ioqymKwJ+an4CV1EI7Z4inkwkDmnbfaElsAeTouJHxv8Li/4iK6iDLzFCp
jpPKUCkbKKELHwUdG7K2AfIPaWvSV8fTiVm/LoNipj5Y7vZHAGmdbi9Xp9FK
ApBiIUsqZFIgkZt69F/DM5PrmZ9tsh0flu6HkX9omBWYjpwLG8rSvF9bjPBq
F4MXedwGmBO+WQ1H3GOrMOSbXSumOyNunFR4tnZCcBzn2cve6RTVIuGknBUa
q9QJc50TUPi1dKiQlnRWqo4ecZEdByrd9f8k5XAdNGFfbJ4x6jMndERx2501
whWeSAIHDEtWCpG8zyiePcBOzkR8L5TCAWwY3oTBdqYmyHcqOakK38gg7xdn
v+0yULR1CqGM+oj8WNHtm1BqKUgDM0jT0661WjiwaswqoXbdChFQR8huYeYE
iYxhxhBlIwTLn9epNn0zCSbp8Kz9Br0zH0OhhsZahh4IFSJ0lEHP2/7CJeVn
ZPRPdEDxG8fnKk84Tc7d6BU4gBoTeUzLtIA1Y1x9GzwYbjD01o6G0hkwng3x
rKa/e2AeKN+as8o9Ku/HHx/JN+NUOBsx17aTpuR8pYCUl8DusJPpWdSmic7g
HqCxh9eDUUeavD66Y0BpHEEAwPmlegdVxZI+b6iyaYxqZut7BaOYbOw2JyuN
vJOe2FwaL2NC/NOtzHrYmxVIqSHWF95xtfUfRfbjjP2LwNKiG1kOMLYqRHXE
f4WUqrf6VgSOnKVkCb5rUz07So8KLuwlyoSRiDiFSBuN3ZdM/sgyHnEo/Ewb
XOpyuhGyThJhVhqcCt8W9PGfnTRjGp3zxwfwSAITHzrwRfH60ufza6Yt5Y6D
SWztFE87ATw0NLkXi2K0KBKbA9TTOhG/A/Otw7B8aZxS/qFzCqj5uQ9Ke3W3
XIwEd49ulXIMb5ly3AnlzwNFXdUMk9R9P8zgH8sho7EQKaRnzdWmzgSmvfPc
/U3fKG41oXyp4Bs81hPYNiaXSK5WTVEeEVIclWT4knbTpvGbeWg6z/v4KQ3W
NJ8n9mgnzV9fNA2Ir2bFfsKgM837xKWXxyAtCkeGErnqKvDGt+HkTO9HhrMK
lEx2VFI2hZr26+r/mOkKusSSFe7c/DV4V18AM5rnWg+WN/6XXIJmROqkKxyn
RLKVRflK24jwxncwzM0v2vyUhxoyOGX5dfL7aUxjTqpsACp1BsZrE9U04B2H
ztVCcTbwIHd5bu0UzP5noQqMAsCHuqf3siYp2Agb3ZMWG7umAzkosRap1bvQ
kSHTJWZwoQZ1FV9Ae9NiMZzSMHnckMzAVZgNld15AQ6nOsFV3wf/dA0TgPc2
YNR3H0ZD0BfGGX7seSrD8V8EeZu2h+klwF/lwgC/oeHtSzg1q9CqKOEOevLJ
XDaU0ZNCvSD0/xzDn9JaQ+ZbnDcCpeNNY4AF35PSAUIGv2dxyUsXaPY8Q/uO
g37yNgLZONT3I3bc/4VejbByrkgz+YfZxLsAZCw0gGboJI18earr3uXVVhmC
Spz5a1PHckaEj2Qo11NvOnoW2LW1LK1l6XceXn2HHwQYbccmNegbK1eZIRrD
M7k5PdzwnnTrJNorZqDv1vZMR9Hbc7BS9C3l1fPWQdyUI5UVh1mtaGFDiePl
b0kBKDNfr8UdclJPc4cfrcCgPb4TlxfFMXOfISvaeVzIL+3+/FXGk7mL6GO8
DjmqKKl5YWIWHpbdJK1o1v8roFElfHSgA8YyE3BJhDMbWIC4QYwcQiLKac7P
9IaUZ2KX4MrTMuuXh2d0ym3J/dooTF3LrGB9sm1LzK3uY7thOcIlZZPFHji5
YgG/7RNF9k9B2HVwoIqmM11CLfeKvZW+J0rYOVlUCMTfvqv+fPNFkyfqMluW
mDfLppPdjOBilUQ+CO6BNUZ/D4BQ81B5yjv94odKb3io+YhiMsBVDe967E6B
NDR6sgC+LyQsZYmQpLWm5rc7qS0kwNS7T2qqdgr2BRnOKj4Sc4WxA0VZZ4Yt
sBu+5sCQc8aKKwoxP6q/shs+6CR9FqR6xWhsWWA4ikFuTauzU429GjPgc663
CQW8iV2MjhJ/FJ/rFASqCI/FZqutOgci/wAWYN+Wtj7sfIQFtFPd++zS71Dp
3feBtunSIUf/9a11fchNblYzpUlOZL4u0rmWVI1Pg/RTLozRbceZt8lZhf+D
Dhbd1P6Ax/bd2Tk+tRcVC1WCDjuLr8Vbn7mZa1sGOs0iP8K4erjDEOeOqoKH
a6lQuYxXGPM+SPdHdV2gmk1iIL0kmFXVnnRpKvtPgK0IcFlbQFizlPWoBObC
yBztRNKHUrBYMn+Ux4WBzoTHISm3RawYV21bP1stWgdrAFSuymawO26YrE1C
72P1zYmsVEuBEGHLkxPX48DBMmcZLppNfYc6vekpQuhF+3qConB4yj/jhnoH
uwz07Y6Jzh4m1/eHzAJRsCUp6rYQTQedgjBewPavOio8fgxFPHaHQlC4FIct
N7VpCI/6L6DfGse/ep2tRHWs/rrbttFA521ZwQ439DJiu3mkpH/YRpJkkW4T
1i7c2/YnaeWLBb/HIntC0PkjC1s4zQraVjZHPuPeE9+V2OcUhZ7RIApYT6gE
YTOtvRyzWlc4C/9N7oZCrw3E2yUBpPnPJZkyYtQxwJKIYqWcYSjPTR4UKt7h
FEzKb/LwqPAoWOmiAEygXzEoQWfUgwts3LTNLXUjHdGgaE7rwnSka3Y1kK+c
a2PNb3V5nMzdJ3u84m0j4oecdpGcQLaKfOAi6Paz/8OtHVW3QDBQZJSih1vT
kVwk06Gh3R6EKd0qoeniBxxCYgUASdnHZnFWF+0hDiLD0Rr3yUEC4/kEqbk5
goAH184qBv5/+njpqp/lGUpKQWB2+J7GqDsa9VsqvwQ2MFDep/yv0fueT0Ef
0Eg5RImueD6g9SCEmGI5nxTgGf9mVBQIZMwAGipay2ldAFl/ihkNVXxxYkz7
ObiKJxJsG+8d1csoa5WW6QCNlF8rm5CvsRGLJ2aat+6BI+HRmT8XERZPDBrv
oWhSRQTOTnk6EaraYZ5h56ubxjUCkwOuXPL9EFboc7ZgoQMee7JwiN3xx+i/
9wHfBlOhECzhz9LBLTULfA70vLgUUhiywTX/YhjLG66ncNobS1PTPMJGHDu5
bWKH8LYi7nz9HVOD9bQXHt23mEn/DdMekOxy+qxlmAtoBPQWSbnnVb8oGkgS
yXeIZy8AFc+cW6UP1HS37ryF4frlou+8D7O5v/WbcHhpv4pW/jgj0MguaJ7q
3utkpe27cGC3RidDgz4/gmwrjpfqiQDJjIbVC96xMm40tb9+zYWYmkZupeRu
ApkrRYPwGUg18qxG63b4Er8AqihF0iyl3rPyxJ3+3W30ggfOtZqtCyjvq5wG
rCa0hvDbETLiUedbSq+Yydo/agGwN+FaZMXBAY68CxXpFAjBCq2Y1XVAQNCx
Al63FWLXOQlaK7ZV/v7M8pwuXLxQmsjEW8+jpS2A1bKdadwnsLNZzhFqU8RW
NL4eHjgYkE+XOnj/c1k3hD/oOiokXgor+nGpppxkLIptI6OFcSGT9b8DHXdn
MVaDgZ3RF0zWxYNbMPND8EtfPSvrED+ZYx0DzexgMqrD/09LCJqnFe5w+Wxf
bX521BEcic+98ourEVfj6czaxQaneKKbTS6+yrVFR0pJVKpZAlonuoG5o285
aGe/APe0JqPj1boEHAoo4HYmN1piWwgCSwwRIzE56PnNjM6SwmiMwVZLGQnR
56ZoR7Nxg7JEyWmn6oKGNeVem0jGI/lvAu/CWBa1gCu0PHy2+Wqznx3UDEIf
909pHSlIkC3jV84gtU4NMrz29r7hPJ1XjdcTVva/XIRcySh3MBHHps3UxYjs
SYk+Leu+ng2aJRuytUUzDNC5XchgHmNyQHG1kcDhpAOhE5ULPUqGu5xG//4g
IjvwImbU8RRBW2LmrYJY801CvF5EMaM6/YxlBK/sPHEKFWAB+5ILUGDPKxs7
eSTQkzsmURQ70WV8bLv0KGIBDBtd7uDI/kgulXsWb522lcTV+L5JWh1IcwlN
M30WQjFkK02tqAikpjATVBSut7DkNjq00TEcHWy5vJmUmnmuuOiU5w5/W3Fj
k7RjFS6ynm7Dyn5QZaBnIZOJ5Jbi4Rl/rRhMiKd/790ems3CrISQk02HlQDb
+5cbMqIHDOi+NfdK0hxhAmHZ/RSSYzWtPx6ZLXOuoYASJBG8gWeRS+7+0blM
2pOgQkCQDc2T1yNeyHTXU4cCbn6vkRQ+kWB9ECmFkzDZJcOUr2Xs8gz9h9Ev
ORMQWz78olR/C3wjNbDYR3foJwvbeNRHkQdRdaBQ8sSh11gBfnOPoLN0Mox7
Hz3vVAMq0OoFwnJAha7jMjK3UumzHq5TmLwsyMVu1618ldMHhWa1WsBvnhzU
YP5tgtTz0Ndef6jNQLGIoxMsthDRvI/QBQxd+L24MrO1V1beaaK2m7ayoVFE
+n/e4ggPZGT8OzAfaCpWsrFfX/HGDhY9kvqLFJU3zcXcBc4++fC512xZUERs
9apIdT8FR/oK+lifI2jQDHtOG2S0LQAWnbPwTfdKqRU+5Xgn7wzHzP4k+o5M
UQqsJu7P1LdHo8jseAfPFIbqr48WyIoUoMW2txh1e2YTz2mAAUpkU+Ps8unE
x5L5fGCvAfrV5dCH07rapD2lmBgccwPj0P5qAjGDHoj1mK6kE5EslDQIeIGs
fteVij1xQHKarssggT9EsjBMZ32tqvfi1ubDpQM4NgJMu1xRJ+8tcfKE7Dbf
K60fW+7FS314J1ZtHxrvGSY/+7NqMpNO02o9zxhpchrEtSbg6dFRS0eOQ8Br
zfDloUsk8ZhkIPclli2rWK6eImC0JmRyRIJBCUu0Xik0bp3GP49sOTX3m8X1
5osvcrT4ZMO/+oBHdgds8cptsBTSfuUOQtj5pJuZw7uCW3MQpc2ZG+6YGcNq
nNryuuoHzIQKgdLQaPHVTSGmZi9AzA8wlxVCgo8syZYlOIzWey2tL4otskix
oWz51zef2lb88dSQdLvBSPVNdh14UNj8cKGzD5u+S4QdMVCH2Tzi4tyXYynV
hJs3gMiz4Udv7r0r38kH3zzTlZaISrhvo3E+/a3azj/f9lXq2SeZAiG1EMlr
BHrhKecmRZt0e1Hd4ClOqndabM3mTmoPDlc/9QVXeMKOIjMMWnAEV6DfO5WK
WLBAXGDlmpZ6dmlWMfw0n8VjTsg3LLFGB8s80JX9cdJVQc+SaVyMaGcuB0KA
8wtYS0jX9JGgW7tFquLa3s6TixeWiuk8O/Y35a2B6H42ZSgDIo8uX1z9kmh6
B0h1vHjimlkx7Gt39OWn3BOHpmkSE8rYCm/V9Var8W+ed1xgUO9HqXvQUDoB
aFLr8EZpIPBg6v8g2itd7SwybLrdtA0l10LDarvRlJzi8iIzOERZ3BN+HZPL
/71fQXjQE/h/5clMun0uWuC9tbKjqphGg3vuNFk6/3rHWYVI1+nrfe0MlsTV
pWwDION2Xla98CJSl+AgEkdxxP/HzB/3lSLApPHDdXEf4A/LSYC8JnI24u8W
90pR+2Ome+ErzuKAR5/XnEmowUDSWQ69v9SIOlxnWpqeFehcJWweUwibYdt9
PxSSvFpgnFUSUcDbv2S7Wq6tkf1+BqCHSbWYDiXqLuGbQc5EZAOnt1RwZVLa
gOmiRi6KS/66QgZKRxpcmflyKFlPyFwDjPI6pEdGSzGwUaiF73xHx9w4f8St
FBeEdpQEcE0dkGi40UfPTlLzOy5LeFFoZox+FCzjeFv72njjCOxm3jRAyIVL
PPxev0qGrPiKmb+amLAaHhMzh33xZZPtnYSzYm/LcBBUDgAr1+UmKz9s03TJ
HirZ//zxiLDr6dy+c2CkW1n/3NeyUvqa2KCgpGtPlgmZWG5NSDeNRSD2ooXg
B9agE1iFc5lq+YpjeGM2sYJR3mpwN49Ee7B4lJUwVb7yYOHtCbpSzw9ADXc0
iGiaf58xTVFsFpZeSA+uFhID2XU8QwFo9KjiLGBNjBZL9HFnECnutsWdXmuF
C9fqvYDEW9+3JOoZlHVtO0eLQhAWM6f8m1ZRj1znHHs+Pp/6Oj4jGdDHWQUp
yTGXHZYyBNbRbsG7xoilvZDN4LcbleX2BF4yFRy+Ha2FoHGLEAB088aQPPRP
ufpqo0+EiCff4EGfXuWy3zM0ckw2Y65kCfwLRPMWSUfessA+L4FSMj8keSOc
pwoNlASmsFo7Ad9QIhgIc5kfa3kGozqvTo0Dk6ZMrtpDY0OVvE+SSguwasZE
xc8pZ3is8/aIlewUQ4hpIFPKsGydUDPuLa6bd72ArMUx7VUav+bo3l5MDJeF
XbSvRJr6Px40fPxeTnoVuR+l+75giss91iU4tSj6AqT+q16W1x9DSMnIFn3N
s6W72pbNdpDmhnHuMubkKDOF7EjX6/iCZMPmZ/QQGje9P05RfjGEfJ/w8nhg
5tjGKghxE3tn85hhh686Upn1czknHJlFwL8hNbV9xUBXtStCN7ApSqsCRJpp
vNJiYdhGYHNt9bgKD7DT14lGqW4TBUPc/PUGD8qaXjb8ix0ghPYWwaNMK7TX
YzZEMiTBMsK0XrOmJAqo0ni/lL4VfZTaKfQk/LszTmzemZVKqaBF715d7BSV
b89ONhZ//5Duja9Ea/3jGOtAJHU7Q5q41aILPeFIKCgbXEjKSfydC8xlx+lC
7bO9UDlsgvEQwwFBJidR8LixUP3UpVnSl6OD7syOxgnu0yZuatFf5f+ipCFi
DAUVDddWObAfeQN+J5bd+JXZ9apFN7AXYbJvKDLpqiSTRmcX0Tdo9j407Ys8
vVaVhIcEhdUtN6toJ/8Gm09v1h69O7M0r0Dm3gXExbD21WBL3g/zAR4sBxDD
q82mpNgGe1mSY+g1eM+M0QdcMr3sWoxlval6ZQ0Mh1wOUvaSMu+68MN+XM7m
6jmjgVX0oEL7UmJhCODnkrGeJYYFt9Ch1sF7xWMsHCOXzERoXtKALb3Myr2Q
AP/as3J7alAZcdjk0gHU9IbppXggNfK81ANeGMJVYtJs8JAaK1txfY9xGacL
Lh3iNO9+pyqWcsPOgQpkt+8clQeBLhkhVbQwo4sr3ZEm5R8IR+yu+kaT+Vym
5vf21VNsQo85DZfIL39KnkmvoTnJ5eDQW31snJCPt62XWb7VFKk6d9xG+RxK
F4zDVrdBpSO8uiTc2FjC7fW0L6rwhXUTf0J1yaoM3vdNIwuDWXSJgadKBbC0
azVFkPwML5PaxXeMd9/kdV1jJ9R23yxCV5+U08jhWZDotYHlqwC7vYwfctB9
cwHez2K8PM/NtX0lSvrEleq196TcLPmwhkpQl63eOJiEFog58Pv5Pc63HjVw
EEmKT9V7ruouOCnyYLDWUHCKKbGhyHyjNduuUS0Iw+S1pxWY5m0xWsj3PXSg
OQ7Zw3G6xzXBS1OV1e5h72ScfBnkl4aF0+cKCfIOXlwPsgTDpzP+hJCDGzUL
C3ubAx65kQLo2yV8GEoMNVq+DM9q0qglEGCIKiX0hkt2vBMyW7bndPvWNFDg
yWgqw1sGbl9I09+kaZ7dYvW9oMHkosg+Jn+TBmxzPPNBCzbrSfV0pXz7Lkvq
HN1N2RHbhMjRBblWUlA2vtA5WmI/xkR2fOJ+6cC3A+MCs4ssNEJhtf7Kwajx
ItWISVf5Hcufwk6KT+q2RSgJrgbomiGOFM7GgKEdwOGi643ZibJC0CtDcXTc
v4bsqHpe5olz54iDgkjeNlLxO4KXU2oIB58eYSMhkUegZWLfpiuvYcstuU/p
IiRpSaFs58rkV0TFg78eX1Ne/a5HbioyOrvgY3zIY5OhmTmBa7Mfg7WT0iAb
chBNOYA3RkP5pbmkcI9N3eM7uXjyQKgKklg50NjxxfYkmEF/vnFTpf/IyU7K
k+e1qUQ8cbv3jg6XJ/BmktdqPercb22xaPOkt2RR02oexCBACaUl6SpcgRY7
hi+P6JbMqzeJFe10Rmj45DwOmbD2oElu9TU4H9QoSDi0t4/a5CKklnnxbj33
TClDFQBALgUwC/YNRuo1R5o/fq/hd5ceajvFsOvVeHVGQ2Tx6JXs/vl1SNK4
8RkQ8OwoOJ040lj4eehu4tXIK66RHGzNxDDEf6ZMSxgUdYF2IgGBcPJfLszm
0DFlW3eEj2ka2/yFIPe/iTqD3kzUoWE4PIbfqWyvwoxgmK02z4zEur94FQRO
Xsojpd1Q2uiy036TcD9YAmat9/UT7IJlw6bMdUbO3sbB6xvyuhRUwRRyTcB1
ckSPALYwXDwC75iSIsPxkZWtK+3X+wVXD39Lig+k/z6s7pQcnjX3ciD7QAg+
LBbdqKlRPv1JmiWBM4KvvxyzGwqtscE76HHA72PD2Vj5TCzoMB9tt5C6Fr/n
sfPouucinGNYiSd9RqDhVuMak/AT1HrLTtDmQvAot/J3HAqYhQzKPBufj9SJ
zc7mc6jAazai9LZ47rPHJ0OJ3r2TSirJjJtHeOzpaQAjFnn9FjfPdYu1RAbH
JnCP5BQjDo+teckG+kezJSBKm7a8VcY/I53v/5oiN5eznXfFKTMSqTzUH0V4
IrbyxOanDljI5dRsArp+S/QB5n87ud6WATfi+POJEdnasQZ590bUIIkGTpXR
H2ki58dmYhuN3Ej3ziu+eMI7KM+TxBp4HmWtdgSrhRQA1BvTEuhl/i1Zhwhs
JerLqRGERx9HJOMcKwn+gBrto24uaapZCp5lvFgUzcjg8Cz+Gx+373c046r2
IWCSVEN22RWuaT5IIa2YKReDqDwTH85Q+mOFOc68ufqXj30RL1Fg3dqjPirM
fVMlupmiCWxFscQi5ms9dEAEFxSAgcl+dteI9XrTuGA4xNI0sNNX5DelmiQ8
X1l23YfbRP72wspBXc8pxFhKO1Rk8BLAhfUal5EBvNG1p3gQnjT4v5KrUY3E
OX/jviTd5mP9ctz/ofJGvgv7q3N25x2xqVWnfBGcPl+UJuPhYkEU4wag3CvK
bBg6XJRquDvTi3773Nnh/IVl3J+2+EI6cZeng5uuHpbuZp0zT3TkO+bEmDFS
rdooNH5FIjhR4pfyL0mCbHOiPzxXZ1HB/2wYHFmUvZ/oeN6CBS1CO3is07sQ
owKaXo/mHIMP+mpyFIcE61PPRTCPkXuszF2xFZNM/B3O8QTaN21O7P6mCC9o
n//yTGRPk4ykpbIm98bidKYwpfQwFXrRmgPsVUgM1Xh6qTjCteL1ImsNQi9s
6t6YXU3Im2EDn4EeKHVG07RVCL1v7Nw8aqv1EZ7IH8J44T803GFzXEDHW9t3
K9r59xuyALe05poAbU6jmWwT1yaMPqCDeTWhM5L1ZlL2zInosr2MDYYtp/PU
oWdQ4vGAaOqPCHC9Jx+QOnTTOA0Zbyx6mSilUgiOXqDlV/W/hBgVjaNMlMRP
kwzMf5P6pfDA5UVoCff73tkBA4eyL93nYE1b9z4fkY7yijk1ArwcjgJjPW7g
P+rg1UXnh5HiU6w61xw7zhVZZaeAgslBiKtg1bo04h1MxsoPBJruXo+Inz9f
wcgdzPbn/z0Wf6DUl7NxJtvUfesuxK3b9RCOzCO4JSRgKyajwV+3u1PPNql6
gR71EvwUEsyhGGW/Ydb+NQXkZiDzGgQUKUq/NivEEykrEGKD4qw7s0wCBAEo
LoAtml7Zl1EFnlNHfDTS63QkJzqjAesCY7AeOkYzKnzfZ0hp+fHzCdoUenkg
hdtfmsPQzFyXs0a3BNvSegYbLcUYHtfp85dt1sYBFnxlFf31VrrC+aJzu06N
SlIZdycJLh2vvW9pmHsiOIpKhKRyP39HIx4+TR59iSUX8iqrG4PcvEqBylLW
9Mb+DgeCN4KxOdDhKQt5XvznAmgvxksiQKkngmBKCMbtZgpF0sOfv5vdB+a2
j6pGophBhEY37LD8a3vDU4XyPp16aP+8BY+EhuspxWE4YqMzXmrMAFHcYjRJ
XOWWQt+prpLmBL/yqdYookqheoSGZo0OJmSbW7CwV29pp1VVl2hP/Y98Tf5r
CP4q2v9hrgUpD+mNwzHZi6rL8sfYQn1Pr8gaXYKSD5PKYVlxVhaP0z3USS2w
2zLs97aP/AkG9cJWCW7Y6yTfWO7JTd/PHLJhJLtm7v51Q7IeqQC5k7/1OGZw
jhZ8VYlbGI4sI3sMBXYsa6t/YEuRton2SDz1uA4aoJYpsI89BpceUpFky7/n
WtR0QzOAt86KzDXM64x23Eeoq3dQKG6W8isvKY9OIiDUft9NN6KhHNYqjxnp
60wkd8n/fe0r53UigLFtWlY4SiDbPKhCJ9gwXNTsVRC+HcVzpsOE7SG9LP8W
hr/fpKDY2mGFM1L24qytBbepNxst1JiWx1nwIaYllkITutk740Dmp6lKKSMe
hEIvmyb0U4qOnqVk95dlbsxwDJmy8waPupmUaxUxefU4ho7Z0leDi2nwRkdy
E2lirM1/wQnlXub7DGqXptdLEputVhuXpVeQxP7hYVm9udR+JgA+llozHSM1
FRthI7/GMV05M/8r4Q7n59a2FmR7KM6nU3p1m/vetndp80gJLeTe2wyBz31e
glNbzf9VxE93glUHSp5C4FBJ6guhcYK4UN/uQA/3vakM0osifMh7dcQNG5+W
+w5lmUI0fzINt6YuMucRI8DZ0UfkrjDSNdVO+nXOATgSA0FTrIeApD30tXov
7iTufV2Ng3ocXDQKiYZXod64Ck3u/WanJWaVUA9eI3yrp0dMm+lhF0N840Rb
AFais771RbbShOGvEhzLvsNr8isxVTRyCqV01XxEcPygM/VvvKwbQaMgAt6i
zJZTh2xMkodVed23mH/ci3bAbFsE93n66NesxWyZDSP6Tr4B/scs39+IptEf
SdSFBZnqr9Q9Qp8lDP+b76V7IuUC+MxYZ5QmoCz+7mMKgFGISymS4iA8wi88
CXx1V8Abd3p8/CQ99EiVdzy9X2MIew1+0kr0iWMakq5Q3ohzTbCQ30WQfOsX
5Qcs4gNRu1SURb0AnvXUGz4bSLeCqCq46amkKeoRDwGnLyQJP+H9jnnfdJz1
u2vPm1qWaOH05FETWVzSOWKvTMAZqmT4X6i+gha9ogMu9bQfhxMM2IgKI7K4
T74BShb7qbiYyV9WUWl9LjMYpNlgHm6i23LRhaQK3dFZwXXypr9vMYIHx0Qv
YVvuMKB7f2tnZP7ZpiVyK+37oDgr2M+fP1QW4BRjfYwPe38bMCffZ4JeuALc
fM9eWSHVsZ2XUOFE42swklwgsO/pH9iW2LepRc6nl7ERhbkZv2GLibTuSxqS
Qb54u0cZ0sziWpE5Jqi+Ymvkg+V21Oh/2O55RFyBHEwSX01S/2txxuJhqjrU
t6A9kmQr04/YNQA5ge8CU6AbFQ9rP9N3EiDap7Oa3x7NkXt6TA2Ds13EA5rS
OyfkH7G+0I5KWtAE9DBHN+tgf6WQ6tGwDcYm/G50xSiI5PSOhqvZGcwProdL
X6yZTVXc6GMCt4fg38bk1g/xiz4ShLBhyZKyceboM9VCUWInqm2Qxs9ZGM4/
7rOeIytc2syMi+aUpH8rWGy9D7/cCVu4sCDoH6DjYL4nNsaMNJpiZ1HK0vTu
7Sr6ZXr3LynMbnmaxQP2FRnrvFhq9dOoMurf/Ef+nV6x2P1jh2lVepmqyk+V
Re8ItP3hVberxwvsvuI7XyDbTiFHzsZzwb0bt8bmGiht5jITkyiHPi1FFzxC
fgpnrL8pYf9OQXOaOAoGBjRG59w9dq07Imqm8GBlRWmVOsrrp2Q1AswDgIxh
xfY8vHNHWN0s9ixH17spVjQD1/wwg2Y7N3Pi1I17SQK9zYN7wm/nvQKZTmZ3
nosBnydj8KcBLt3Mmy1GF87LQzVvxXb1FWBTHfZGeDoWNU0lpahH601C/4yK
exe+qf2CC2BqHd2Y+J/eSCUUZTNuS5mQeUZgC/FFYDqPUEAGU29sCa/HCsRj
du4RSF+vLHorYWcmRiyuqehOMtFFTHG5RvbLo4yYcam3YvufYzf0Q4z6TJ1W
S3ihnp6J8fIXTsP+47c2R1n3fMqmM4VyRxPPBY94wDuydkvnRIC2RtpgzIFI
VraMyoyLlqnYZKTcUxxpZnNaOcSgteag5ESNV4Z2OnRnrOUhNGBN7i3JnORq
eMjgMy//k/eYn46V9O6M4hGlGi4sgKDl1SRAxG7GFm4raq0LZearm/OZtaWQ
WJcP0A0zRkb7LSGqpZmfzEXDlrjOG5gHkOQGSyf4wjbjByEUNqSDYgaB370l
0hm4/pNPI7CPIlGKMaLqAlqJz00o+MYyZKLoAhm3EuoV5qF0aXl6D7CaE9jf
1T3Y/KbjIDaymHuPrr0NgIItS6zauhEXkO4P6gDlBewWZnVhemjgRDIeHHq0
dveWmr9mF2MtdfFd3Q4qUyhySsgs/oN92tpCAsZZwMbgSLOcQILcaDrghbqd
kTIU1F5jEa1m7XhesVmKbcwWbAnEvno+PhXg1SI3pkfGevM2KpITTJ3DBSlJ
e6bQ/kxCWAieLnP72d/q4EqXvIP6PK4meJRkV/OwwqSWAH3fN2itysq4r7/D
QL+tAplyXcfwMy5o8cwevltVtdEk4jsUuYW5sV815wqcpMuMGAbwYyXKMQxo
eFdTafQh6vFv0i2RuVt3nTriSVYHPDOY2ZanuISo7S4pGtINEMWLwPQ0EGF+
p1UDsl2kb/mG5txc9fHeY3d3aVDaBzBST4z9K0hfpK6mRLainuggtqPCaCc8
6TbOLG1yDQSpuDAADJHu06StDmrqe7jXDDIR4VdnjdQ6lMNw8sSrVMIG8zro
3syvzHJ9UWGmV5wDty9ZbbD9+NcZARwyHzI6hR0FCCCXo1bUiq9blaGgu4EE
LOReAnS80IINETpFMgSTsxeTBWQe978kr8WjfmxltcYck41IiE8t+PLGLBvZ
NUrz1I5jVSLSW4wA0bL/7fAProA3a3cIgWWRkv7KpIlS6hUWt+uP2NAU4srb
RS8JxIFhKgSlbA25LrseEf9dXq8rcaYe1V7B6G44TUT/s3U/EQfQ909rlTVB
4IuYu+FNndDAMC66txCa19W1Hjow5xgbpUomV9FPzH11K0w1xM1xDJH1KqAI
AK/Pd2gmPiXNICNoTPuNswZry51IRVss9kFbD542/vd8KI9U1Jr9Z9GsCGm1
eqkpfqxTuXDV1r3tzYYWLg+LEDveTTrMWZ7iGp4Qsuo3tV3ku7MocDwKTTfE
XL3hAjdCmTC+UBDtsSoslPAhOwmX8ywT3QN5qb+XXey3GiGaVcGWzeyD0QNV
LvJ0xeuWL1ClRSk4lsB0is9vz22r8xy/gCdDT/yyLintP/H4Vl6VwD27KWvD
+3QQdOqQsBnb6yAeIApnfLjYioppaFDI8C72AZkS76d/npLwphzE1j1cmh8l
ARag2xHSihErB1/q5DWqQqsUYmpp3TUfqcY4IioWObmUlWGE1kHJT5v6189s
w/4Ez4N8Fu3IFdkrxRAnFf0AwDcr8FYTQfnKiVUYLffWDvEkxYDoMiLCN/ZH
SYR7uZ8hoRdyLG1eoviwv+fmv2nB1qW2rpgdKlzh5AXt4fEwK2KAFH8Z/yHi
JABnZF0EbR9KmWe4kEUMSf9qLRp1NFae6Z27BQYRD0y2irt3YuEhHhyWWxTp
PbF3x8xp30wBpV2AIrfxGy2Tu4OeEzoNGsbLvF0h3LzBJLDD9z0MnCaIYM1i
ZBZ1dFb+1g8y1F0jUGh1z+qrsq/ZV5jSYAmbGwfnQOJqclBz56XQqmuV6xek
fG6rPaiA1CZD5J0P9xtzxqFYxuJlknQSFBTKi3G0HeX5YTyBUcMN8Q1qB3qb
dd3dP1RJu379gHeAoBtM6PD3IZMdsdlLxGwUaZ29Yz3yDpyntpGCnaLzaW1/
+uCiCjfySFlJr4sTO6QEmq0P9K0CD9qgbe6iy2B23RX8MwgO8OkpuWSwDnYC
OzhKbX6hdZ/dgCg7VYnFvC/7wWzVAr6iLK4z8LC1fdwsoU7OK9pHC/Rfs3kZ
eFxZv3Lxe+FY3ryu3dRI1d4rnoeFTuaRN2y3Xx6IuxdmVmDs5B63G9kjUoIV
ZuXqtOMGg58JlU1LhW2buc8WE0n/sRFRgyQ/KvS/CQFh2uEPccvbY28DB/uX
2H+/ICNbQoOYaBQrpueIc63Yl2PmPvbfK4l5jkD4W3mB5Z+m4rQlMcG8Fsfv
RJiJQASTbGINteY8RvbhqAx5dxxjenQyt8E78J5Y4bGCVEJK5AEH7scOBj1O
QQaqFaOmQwlhmywEesjFrr2IVNpxmbE/22miZfbus+hPgvQ+K9DrCPCvMnD3
dB72t7x/N3ctTtSz3LBPKmI5yE6BIZbHNgB3F+vbqHjgJ9CwPKEeoSfxYoT5
eBtcFRt8rcXd0pC8uPKn8XyBgodSYWyx/LiEA8zt7ejnEdAgwF7sxqP+QqTh
tSQ0wi1kxrVwJLJYyDGteGNQjA0cqRMhSsN4vBagcEEEcxWdMoJob59lZNhO
9kaJFr5tWuTeTpLPHJQg0G9X+KJeK1tDj/cesm5TqFg0OqCHaz6yyKWtMxHP
lcWeUtenZJ2r2YrgP8NE8ZLyxSODh12/LHVHvq4rxbxreBnUCe495CMCo5LF
0qGp8QAD0y9FhAVR8tYoQo49ms4RNTB9JFvQXTgSo47xjkYa5WyxHvOcQPHe
FYeLbM58JXEgT2fHPKnfRrfdnwR12/fSh3JKKFSjibhoWFr7ErGeklE73yhJ
z3A628L94RGE1IqvJNJE7plpYiYg+wSemql/uR/V8oP0bHjfuVdWT7MxOdpC
rMUtoIJ6ryOl3jCDR1+hmVrmJ+4g6aC21rCW8dMoZaNkwuA3ka44xB2MPLoR
+FR5GtGKMG/BolrkaIwzo4yY6OZ98HftAj69wOGyKL1VeOnNTSmRjM0j34Eo
qVeGBEDoNB/eNY1JRqNBIvOwY2HVsTgcBZovQPlL+WLhTAgKF5iUTr79puuD
SqYOUVBqgEUqkAZfZhVv8641FI6jbSNKpQtGCt/DqG44Z5iGKms7NFfRdNFx
StC59BE+a0d/00AYjkWcaUzP5aCjuKjpIWtr2vx4S9zqJ9PIc0n3l3JhJh2d
N81DpSJq0ij8mS9ALtQAvleXi3M3aGRoLHzpqxG86+JCX3jHHkIsbXMllLzy
4Xu9zuVPDCGy0xgTz1YKEKMveRranDzsDDLe/9Gl9Il6iBNgv8REIsTFLCMP
6uRa5N7HyXAy9kFTP4sx+wF8EfEPMRxIzlxHxlv2v2ICEhKRT2d8Rp+j/LIf
a2PezFAUvTcaJU7L7cFwi4NcRLg0NUD13g1/G65Q3HPB0yOBuEDoGLHQ4pSG
HyANHvPMz/VuwBHYL/MuGp2ZlEUiK38c+zsCOsB0NZD24hWmaalVnAnWnIoT
19ZOVocb3sqBeZGtZ6fyD87lMxTwGY4MJY5M2ODWiq3JlUZmqBHBrKqG5tfC
+WhpOLcoIi35jXDZlJLXR8KTlhE8rH9gST+sI7fHFOjQ4/WCHrFtGL5RApci
Hou0A8RIhcUEMswidyNzIeTJOvRfHiCqphqSt8HxUe1WjLS2ruaAIGsJczXT
yfgMpMpLFhZMqshOdx+nUhw4VRgX2mYd4IXf8A6OdhToRVVubqScF32UVA9E
V9P1DQND1KdpXePnUwZvXJ/yiiYCnGwTHC1wiA5n2zUk+qlewGWoqtTRZcTC
sx1w6FWX0FXIbDtbU4fY3DYO4ZW8OKC5T7OOMBUqDDqB1KKH1uVctBI1539l
rMNPiczflmLXL5wMIOkAYLTq1Uq6oFu7GLY5uRCjkiAVkhqbdfHK/LW99OXr
FjuejSfA9Ser9i6/C+SUMW1PeHWtoMHi2jNDotCXoi78eu/XGOEXdwrpAjiZ
UGtoWL9t9l14KCOJql8gTecA4JnhsTTbFF32dpQkvyobdjCAVjubnIj0blcH
FQUdB8+T53RL8SlUaFBkGzZfekIGaOaE8hNqKVe1G+ai2vpFEUOaKTGpWgg3
z+XAlLiX/E0EYWh8Ej3rw0JjMSkKsKJSX1UQiUUCKjvOWOLf4r/JaIA8ojV8
knusqItVEg6RizXjiZOzYIW6Rb2ERqyxoHQmq9pyedWkHOpw54vsfd2wZv9/
ECNNL9DMXysnn6WuipwRnceniHtTA5dAgiVX5wq2FrNMTjG10AHpY7W9TH5b
/sGdiif0L2lh0/PnQuthn8vbdSn19uQtPCFfvtUIxl7YJ5xL0WOpGf5VBhxF
QOBOx0zxz/yoa+q4McSyxwoTaJomMqpyhSp+Jbh9XkOJHMK3iCQXz01NA8T7
R1k7QyZDiTn0+P34kuPpnkztHLZ3tLG3WJFYOOTMQQjiRS0HoQUxTXV6uYYO
EcLLx93Nim3zjjyyAPJSwT+B9h8kW+bN2EGgr8tlpdiLono82RJNMMH+DEPq
YnHo89iYa/HMKL/kIJXoQ0bCSHMAPwG6XXRkYO7CRvXpWoxw40Dl5gjbsg4B
lkAvH14i3NSye4oOuen/9Gf7vUxpqTfDY+8DJtssETLvF6xoRgBpB8LltmrQ
Kpb4Ej+rqUpttCfBhMV399lRWx14gY79vJjnWrNmr+jHPMNqTD01WQUWQUWn
q9kMCG+PAe9bkV+S12j8CTDsaetyGITduXfLCzW/TMn2Ud8y49SnuKHZwNg7
UjmSr9lcPh+px81ZmGpR3y0HaZKU/V/f6OF/aPiOgmWs/gQlu65qtIb5hEHr
/+tQf0hHWw5Xr80DoP9KdRUqLXPfDwqPI/ltId6t7rhBgWLgJ5nhrssOfR4K
EviSvzT+hpvq3LzrM8SLahw6YfF1MfCc7TMC1yyX2bwt1uCQTutGdVR/jbrr
vNmmB8KDEcKnzZWF78HKygLH9YhL+Sv8YfuNEoAx4Y6hAfBxkgXNS5yTl8q8
HTXfvjBIEwlARHVg6eT3fKRtJBEBVOqEALceYYxFVOOJVAzWJRde2cboUAxD
VmY4GjhmRSPilKT31mhnYqsyLeGuU34gIBF8+bzk8Iiq5wLXggnUbl83Lox9
pBSQ7SAVaDKjA8rUcAR2tuwAGmJCZVSjGR+Y2GtklJsnqfbeOnWFsWgkeZfV
0BvHzubIOKb7DzXlR6ssAPizaBncmR6RN/LhcpGyEZVhT0Rh+SVY6BefkFnc
0mokLre2smKWyuc4bvFey/B0M2q86s2sUX9VOsNg0TAHboDxHDliDxCFRLCx
CEV552RucNUgyBajUPlYpFuJWeXk+fJLyLnemZ/snL6dZFpEuB0KUD1jVEjw
RnLT8opI/I/dEeUGXySmLVuzTy5BhYEI7baLANwPmG1uOimI3sW7PWDPc5SI
lpsdlK4SDRQn6UeIFOMpzpeU+TIrDKrSiZnmnPWS8h4ndtYi3weyr00blO9s
KTlzcxspgea/CFih68xe4bTavHMftUEJt14/Oi1U5OuczRsRDwcNROOXWukL
CW/OojhVqUMS9ACHzip6E+XVrfi1lNWgrWeBFfAFLCy/b7IdPCQJ9US1OmP5
bFtY0btVyuTzZWDvgvh/plrQaBK3iWoeWHI08wf14YQ7oykluB0EmVZi9Dof
uAlz9/jE65MnyqPieE8rl2bNXWykCCFRfx1s4shXY7qQiXCyXLh+OKFo7UOb
CMqyNL93mi+oesF1Q7bCSUlZVl5vrRh6xdGEOE/OD5VfAT51CaX4322quGm0
4yRBAv8ODoBdBiuybcPLmu5SklU1bmvJ1zlMlDHKzRQHuY5pFBvy2rEiRPFi
9Z/TTePT3vELJM+0oqa9o8q/UIltF3X8sn7ClgIx/Wpkshvuh0oGTjoEhTsF
I8ksPImm1Eo5s2JJGoc9cl/CIEep6DjdRN4pdh8xwAwpjX8iY/2L6yasJ8G/
3rZrYK08tJZ3Q7RcmdBVbmL3YY4zCgv5yoahOgLhWvWCZYOmdl3bFm1yZtCR
pnNbBo8JCnlUkAaWhrh1dTbS3iujIrsVuNC5Em02AIo2laAPphtHegUYOC85
XP3i9zngEisKTUhOX5UNqSdUkKwO9kfoh++XiVoHtyCqBtXE9PhgPElE7nup
Kxnax9Ef64fCbZ1niB2D/W83SZOI88hihPWJugVESQ0LGscQBGrmLpj/W4v4
XAhDjcRuPAIyeBRXsbu4KR/g4grjK47dJug0avSCYSL+Pdsh2g+ir156/Rk/
BI9+4Mm7T0HPh7u5YixGmBG6CbAdRn2YsmdRCkUPiFVlzOxYVzM6eRcXsjLB
/8DByfXCl6/kdK5eUv18q30mvn5dFmqOJWgAfSuJ0oX6Mo2nJkboiH7qarqQ
fvVbHZ9u/Cct46dQUhS6yMMVBWJQtMshzHVUhukI7ApCXaKFj3lQbb/hWGmn
qImllqbIFqYaZ6cBUpfwA56V1I9sKD168s8fZj6XYqSU4rCzuRzhxW5i8S0Y
FvlGw9dT2q99wxPgNVrC1WGcqOR/LjDsTkMDNwSFwDqaiLsp71EBdi6NaiI2
80AysO4uoCPQfCQDI4HcsYYeHs4vSbH8QE/GKaSiSCdISJcRRZGwXpb/QbWs
LkfkEJuQu/3XEA0efPZK8NXfktA3qmbVsmTpqBJRAeJZVtIB04WBMAaR1xFk
XBLgZs3lX8+PTkdYTPHIaunvcHrkBHOi+cxt4D8prOkUau7EDUq39fYV1s6I
d00ZLHg7XTJP6aQyLyXz4jKfP9ulWIaOjb4We3Ddk01SRoMxKPAf4JvRGjf7
OmPdSV9fWWkhva2SO/F7QcoBXsJysqXaXefFmVUyq0FUej4cD5pcVmj4zGS0
f9/ORht0qigIvoe9V/Na3JVgBQ4MGVFM6RJjq6/Hy4EATdkBYbBpYWJ9Z9R8
DipCku6epbQe+oZJM1O6QSiAz4kEjBAcNotBZ92vxyzifAtkQAhRJb9PXon1
d1rQq/FHjayGp5G715A7GwnX7yBm6ZS5d6mx6IRvd8fTWtSQw/QD3yns4dM0
onswQGfn7FAF5VepDJOJv2yo1rLsNi5mxz/MI3ukGLvBCu1w6iJKXzj9fgic
u7+oOJXeGpdUGJKAeZ3hNmJEMz0jfWzREKx06YgrGLiIp1s8E2k5ROhh4Wzy
F8A/nm0Ta6VIY1XVWHyFyxmSgBANcdtx82DgiuiqF3q+dE46KDewgzNLdHJ9
Hjvpc3PBOOTRV8R1ttq0FOdtCRUn09ZEi3zzDSL7bDTAiFIg1j0NbjXqZwjP
1r0EmuH5PT6igj4X/F6mwv2FT9UsxgGPK7/KoCYPFEuTj+aR5WDef6h0nJpD
vLPayfALb6yP3B9KPrQ6l9YcPJfvx50USaqI5Kyub50E17DFfF7MZgNO5AAg
nrX4wS+5Q+Mu8VejSfX/GNop5GMLI4eWYqXktubn/o25vi4oBFowgxHXexLT
hcL5hA4bE6zG3fx+LKff9Do3CA0BJL+FGCCgm1EaD0JLdyV1EwlzceOq2Yrg
U2C3ARZAdfrIc74pFVTKKFFwTsU9PKMtYxt4l0a3ufudTFveaB7rokkr6uZx
a8quk+CeCNclS8gpSl3zDj6VLOKJQu6xZGsErckdIWG77y1/If2r5NyN1Ngr
cgoEToRye4/pnlWLMNPUZlyPxJYe6z3m0TShzlOCnud0rzaogIze2tiYc5H0
glK8ED5ZDXAgkmwS0jtoh+0K25CoWrN/JaNA9TcxGguyiwvTsfcRLwAcRi6g
HbJvdbh49slPpfR1WvDcpzoha+RVFhvkPlPvsDGpRcbVT4H6xbeOYyoKFM15
ldRbdzW6KUtN3aUGLzs/fUxD0Tpj5X+o2ptPfQivvqBXl26fi8a1EwAI/+17
NYbBYbaZzelEeltOCxI8iEQGYXj3npRVrph1PyBeAsko4w4PXNz1GFvh5qmA
v8YbnW19zBNqLJ7aufHUR+a8uQwsyOsd6mL8EBS7Dk3M6nXXy2nv7nlrGv1g
dkk4Aej1KeokI+STeitG4XAHusjSizFjyUFjsjGTpNt7zuzeZ7FvXAM2ZsMJ
PXh3TZtJ8Mm+vDpLoyP3PwwUmpQKkTOpF3S4P1F6e/w6E7zScLl0p6k2/jom
FHoSTihGwC0m1sf0+bCkVvQJ8OuaNuJA9TMpsBojap94NreP2yBuzd+nq+lU
MKLp2HLWLLmE36pG3QV39tpHfJp5s2lgdZSWPW//ePDt8vSONDZHBWLfbNOo
pn7WDgjl+uWsTD/fXkewfPjuFMuKH5GHvmoGz++g4aZV2SFF+EZHezdxJ0RM
ExknlDfyAJZ6eUNt1mHStLmmSmITMSkd/dJ+kN6zxIFyjelr5l8Xa16lIS7b
yEhlcKkgz32tnYqTb2dBr3sJWSW1MNJDEd8/uSJwfTXCqG1ay0TGPe2Z6Jrm
1iR0pK5Pcj4ZAabhlLCdm0PoKssSjZquNvP4DKz716nfiD8wl+o7AeuzNSeL
6X1Cz1YfmZWOCvfkJ8uLFuWo68ODwAGRe1gMYyd/A+aJ1KppbJT2Ym2piY9V
GP6NBKcjnUv//eq5BNqyKctXye9epwEbIYD79/ijzgRGwauKP2KejuetnVuS
r7vCuDG1IACMH1wlh+rhVAIX8YPiJLWprSbjM1TvtLZWowljq7W2q6VeiUyC
Fj/1VYL77ATBhZjtGnpMhxphdKYv6Tu2Zu2ykjdhu3UwuR4ApyBBKLFr9UlV
FSCBefXGleBDIjiwADeyvW9S7VECzKRUVkCYgWecRpXDLJ4a3Wy82Bc/aF4h
VkjEzH0b57Rb5cjLsFXct0ypodfB6Q2hEqMWgTZuvx/L/FCKDp5SGsumsyjy
DZs8Y+qGegm/bPuBWzLo4CLJf8r2r9/vdGeRyeF3K3Jq0PuKHEXZdO2iqguA
JaamBd7TXPXVDTBhNbvKSJxIIW58XKOmz5/pkXt2CH2yILy4Lj4XokvDC1T4
uaFMv7lrEwKFPuAFcuwOf22nwLiJVM9nYHo/VPjodR+DqkGQaQzcaxHOFxph
8xq1/oLWJGAJS8IJysJZR/jJtL+EWxQN15Ej/f9GV688Kgp1UOvrLPKmzlpG
2WAzpBaFeKaxXvKY1tLALMkm7Xy9EmEEvaDI7XHumsq6cbaXqITvaNHRQaNz
POf4Eqg4StHYibp+jspxYAuyfrrJe1ch60Xsw1ppejcvAXkWs/Rk0tQ7K2ua
zC6wLOOnNhzxfwk7K6LxCCneAioiuBsfqjUYUdXd2kpOhS/jJs3yX+okbxHY
WF3F0eyWvGt8iEUMEAGXttbocot+sg97U5vfU3zvbmFGvFZoIcqrI+hJ9v/W
Ff7VwxQGWbkPYjxFqDCO4D8TjW/ijHN6+jnORnvdq/PQ0uqWMXNMwk0KjhJr
gSW132RZvNz9Lv1EZP24qO7tFV+qQ+RZat7lE2HacrYO6fpbw0JDbduihaul
pLnarc1qn4794pfPdtSZfI5dm1zFBtmqyGXTNUmVfxWBAbEp0JO8dOyOzLZA
kEOnAJrOnPz5zYUzyOI5zY/YNhpKUaskQ4eVFN58HPTcpOwMiFwm8fWB/aSE
j3i0uLN3I6lNLdsU6MvIPDMWFjIzNYNanuns1H3GBZ5wCvQRhwrMKVLP0y6c
rnbKrdoLgE4I1IT90QtNWvVZ+TL4y9kfThvIg9cY1aJ93em+k/iEIn5waMIe
DbC6nf9D5iU5ETEBfzUlLftd0Ar1yB+quzYQlCJiJDRvUQSjQ2t65BGg22nK
t2RtxkzSt6ig9I9Zyj1/bWQcRFhoQ+JqiKo2u8CCAAzsepvZBG1CoVDzDsG/
yhYmFllUQhuHRMEKGPuXf3g0GsryTH3r4pU2oVLMY0PqarrXqRnZXRigIWBG
zMYZtuIoIPX94dR7IdIEUr8aze4xB9qTezqpsLC/7mA45BVj0ycVLNU5y1mH
zbU2SZ81SO7j72QDqAc1DEGFAyLhKS8ClkQTjHCtQqLMKaU2XMbt6gpSEpum
vgeByqQx+H0LQ0b4QtTXMX+KG3NTITDq/O+j5O9pKpbRlB+JjQHMW/Ndi+ju
SkbMDXASGHuhu+PUm8QGZMBxTOFcyQC7LESfgVUaHS7WWp3koA+z3wGDBvdk
o+xdna/zgzqU5Rdj/ghRm1vqmOOimcHYMDGBXwNykS+cpK0Dtgjxf5R0zZ+V
ZiQ9ryoH2GqT0mD5fCz8bi/Ga92+bTN5998oBlHqyzIZ7vFYSi62TDFzGIm1
AdsQ/ufr1D0kpnzJMJ6GkpRGxggq1YvSTFktvWWZpwKrp8rG2jX+r+7Kx2nR
sxUVeW4FtDXds/zRVkwhbX1xispJMzUYpYaQpOaYRDvhC9rsEpHvm/BtS8m0
3hzpowUPrp6lMadWg08bZIO4EoGf6agl4zC6/Od1um+tvqjwTR64BW7Rxt23
4Dyg8t0zsu3R8M/2q1usauXN04e/3fwuVyaMJOwerNJMAEzH9j/faGXBr5yo
v4IWf+8yuYiIas7HDDALcOMSOPQh4p2CMOwVVn2lxEBi6AvkLHA4SIp5tK3k
26rNJ5EW81uMISOwlthIQFZ1HdT/I60CP/XJI6iaobm5D2TsCqCI+dhb3qxg
G4jmQpUj7TWUPolecHZZhE14Ee7Ib/68a66dOZi8l4EhyB+kNl8DbF0yAWC3
llqLqL6kx4BqmYOWwlXuEUIF8WCp4l/I0NWJWWVSncq+jCIck2x4Czb22CuU
Wax3WWl+SaveKz8gdKuyxPT7RjDBa9FF8RNdG5ZHxJrLOCIT/i2/O0qj7Prz
Mdy+FBrvduLIP8B7v+Kv1uyTBEeGUrOvsgiMXPkAT58sUP8pzT2bkv1XTupB
9HrzAZO1sQvi42gP1PikYJMG4LwGzg0sgcp5Qk5BeA6kmiUveOIPalhPgYOR
0M0m/BkouV2NNDOLynnzl+dWOoGQjjhaMTrNfqS19HFI660FrZe60juPnso5
bFRwWj0iHE0F0edMHNF9jC+3U4XGB9cqoIx9Chy85CsqtqUrbymlMIdxuayq
C2o6rHljPN/7QsVEAK59jUtpB7npc1QYvTpkDHc0DprwjTA1W2XREhG3x0AX
I6gUgNqiU0XNLiwHvG8DUoB0cyM8pgV5wPIGFNw/IJopHUV8cjEOVyI8iVpI
mtv3+uOurqm1tjHd6BE5d3S8BfDbvsdbG2Hyta9diI7Rd1P7cv5sFXc7P1hk
EGz+j/4GVACQmqp4phSwDSWQeefEMIMb15xKpJovGDBz6cahEx9bUPdrQAwc
UvGNSomQ4HsVKAP4pk1tk/pgrZYV/k4kTqGL5W2YeFJ3gWBlv6HU3DyEyYTb
mAb6UYvzmPNXj3HQvmi0nsfBV/Eu7WvMkR9WbRjpoM36BQbjkJlIyDZMCKXn
MY2c0peQC+O7P2CoVoOwUlFnnuX8+T1uUrkak5j5Ms/mjmFRmsyNbvHQB2jB
PkiIwMCPqXFJwixZr83zvZTMzjz1mGKBumSiWB1vPRijC0387l6sT6HY2iHh
0kUU8218xQFyZSB6d/TganXav3IreoJrxijososoQkbPnuidWeVXaJrG3vpT
kuEkfxS4LXhrEz5V/Vk9KvcM46EnASCjKtWKAZG1Jd969tqwDQ7HVI7FCkae
wB5SwHLndaqEAe23oJYxhkn/hlEySQ2H3zfzG9pQaWnRHE3nxjd9HD3qGQUl
nX+AuOBkGEs8qq6m8gwHuOga/yXteXriEflSftIkvo0T/yDfSWZpFySA+KSZ
by7XDgHtIn+vwCwje2Vkr0b/W1TVjnJq/QYJJEcrpusktu5bbcFTFA3G6oYT
lOghdk7VfUsvuq1NWaViDh9YOIGtXzThKuG0t32nHMy5c4KsR16MSOGkbAsF
Y4FN/p2lBTVCpAcodSeVp+IVShrTNg8g6oKxgyAgTb3GSuhxZMIOELzKioeL
+LwN7dv8e2ADwh9YT3QMNSyDFcsRVr2OmjJg6u/Cp0ofczA3dVWKFAIDckdB
r9klZHFn2763yTcD0GlfM1A2IpOwGsezQRUvQTLSL0laeyNpYJBAHQk/8snX
tLKrvv2nL3nDqy5gNXscMvj6ypDPEoujVKxZW7vC/x550+2CgXFsg++A0iiq
xhKQXk9qSAiotlZyb6Ch6ux3YYN9YU6WhJsth1ZZu86dvDCqxXdzxxWauWBD
GsqhICqPIkoEY0Vm5DQMbWgZbCyKb1Xvsnd70Zvvd1+8b/XK3VURc+WL1+Rc
yjG/dkFN9fnolWntnFTrkw9pshEyt4+6b3r2KcY1NSFvkD3dXr1W/PKpUvD+
8L5WtikcPag+MNkqDESxCdKTDbMwcn6xnIiNkPFtDceaI6mICK2KNMdhKJA3
+ObqfEL99jl4X9w/ys16hih3kDx+8e9poLbnsV8yHyecfyUltz48ZsA68Cl0
kgDvldTXJd+6X5I+4VlQ703O10xXOVj061gXOt0vlHn6mk2GIKhJ5kzUGh39
fXKVbdCr3s9h+VpyWRx7hzGWq4tyiVbx6ZkzKLUkmlmdfgn9v4zGm4xlOm1T
oM8Du1gww0K83g5QGbdUS1lRnaPIFEtX2IPFytl6eGyQ/UFZ3Kr3UXFp6WQV
/TDJxRguV7n9NBxQynNS9GMY8qkfIf2Axo2t79BM1k2LIjBYW3SjmjrehZAo
FRgfDMrzzOgudMDF9itIi/eo5H1HHB0JFszXB7GumNncNxDLiZG6lptEYcML
LGa7IaexV7MKrgO4wYDdUC0OX4VES7JK2q/yIlgRmIAKW/kNiCptJu9ZEagu
nI8rN6vKpA1mJaI4fhkwW3hNgTChW2pWA/0XtOxWiu1Ls0GEp9mFuQ0g8FZG
AA5wTXbS7NtPketLALS/Nw9VORUikwP/ViBA0Orfa2RR+lzcARulpoIWSoeA
rkIa0GGKeuox9aVGNmblD4SnZKbR30P3L1yoBCpW7Rq/TTmRsH1/jmOPEACe
REvQbabfLHrg+TSe5C9r/1wu9wxeetUAdxghAcTF3p2TTj2RyCgYDhfHVwkw
c+7Mzf7m5OZiFDhmb0SZMu7S/Pezq8zm9Va59LOLE2ASzMaYeHqfw+k+LHvI
SxSl7oOBATjrq0IQaATj2ZOz1sjePTZ51U865DQxN4pSt1D8j4xJDa47M/in
kIv26IBWqQP0hG4Bp4pLCH0Uj5JgIBhMkk0HoYzt1e9g511qxLwn19XTFnvS
fNpwkgUmGmMRRy3NgAK75+6XukOQvCLYoZCaEvi5wQH7UQggpFhOi1fEuSMc
Tk5vDE+JJ6dSqSABcgVwAeW8H3g1B22Qyj6WKYeRI49gQXlxjYvH3mDCOY5A
DMwpOwpqd1fgJB/YJQdG71BXXOMRV+mfRFN4GLnDPrX/k7mJRjDOkOKIDPDF
edGc3MD/y8oTuL/JgKSe1G2AdCjuKFclNRs8J8wGHVD2AEBKwljaZ1U8ajKM
MPa8f5wNhe0n/zrtPsbml5BUx7n+O/xACk/6SAu39DTOvGCixCYRFhnNY8eo
+WrtztSPzkuTUIzQ5aVCTO1YSe/H0aetacCk8eWPsHlwiDnIpco+8SGVxdhl
1UCp02WZMa7W6bC9+O/fdNOz6o1gfqRzG6PDsKheQDpv2X9FY72U2NjqGNHA
JAPEZFJB2OHqtpAJAIXFatuRgmD7LymTzKc/5jn1eU0OXTkmYgZagHoZCiHz
Wl8uaFlMkRW3Rv8AMfPdaC4NHCEJPkfx7Yig2diV6SWsnlA1enE2gK4tSWY+
HcNtXMQ5e0EBsA+9ntbX/b2GO26K7mZQShuYVGspnNxKQBsj4TKnNf03Of37
zjc7tp+gISObD/IGt51rqo8yCUnHDZOtAekr6q8/Znf5J+tZQujvBz8r0DM/
/BC7M4FzCBCKHWOQZJ3ExsjJ8WPy4GdqwW2rspWmiPKJ+vwFnW31mSW9KtEP
enoO4vpyw6m3vjVw8E24zzu4t9Ge1GPIk22unzpRD2aQSq5FZFG8usWb4BII
u3XuqTe4SpC7/gHCt9ro9Q51YXtWq0K++rzN2soNlJATr5q0D/Q+lZlxxkxh
7NMz9ADmaPWGsOPi6OZtJmBzXF3PtERgNbtR9B2Z5zcJpfyKpJHH0v2SFMAA
WaLItDR0WhPyCPsQ83BlaVvMkdB4dX+7avW981RHje+ho0HMreGi8a4HJj2c
RXiWUeSpxuVOqI3xxxUA4mmQfUqEmeWRrtDop+32II8SVkqjmTM9PxRl0YdV
Y3tUeJ9GxNkTLuB6blqZc+HlpLiavRtVEpBmWqYUmaBsOXsQbO8IkfiuUiq5
a32vUynDKae4cFInoyHxStS3kaACm9mPHNlY+3F3/3NbOpWsWCjzMVLD3zRO
p5ILf9AbM7Tx7SHh0Y+BxbdQj6bcStrOwZt0l/NFcwdxjALtAF4q52jNqMnl
FMY/VYa4ADtkhHLkG74xH5u6AQyVm6cag8USIxG6tlYca6Xs1WRQxAVqbRAT
VEuXFQl3VLMRu3R4VYUb5pM+zq4tVzY5XbjYIoj/yF92FNOvPyTrc0qD55g8
C7E1FF93ngUNPDTken+jh2MqEsFkocrtc33TfnfiUdWASPuVw6r5DAa24UFr
5W1QV3GoGQ7qMtDxnywpDw46wPu+Dg/NWFCdmS6k5Avc9f4Fd6+CUImMyO69
/Kr5pHatsJK0Z7CyLo6o0uQbeSWMoHOZJJCruQnEErBz7Y1+Pbr5CferBROj
VlKGLppXQZ2CLLjn2od+NuzVbhrkxl+ncqEgqyAofk3sfOxfWs4wV2UldsaT
Jq4k2ueMlbpGcKMgLsJTzuO55lL9rTSA75Vs1564gUqq/DtFLrHtOO6SvsOY
skwFKtN4fc/lSThJSTkHa52J4l9WYfS3Utx8Z8S+OOF5+2Bbeg4StRQ4pQM8
h6gpFJ5i3oNWgvxC/Hq7Tp8FetOsXoCX2RQI+feAmNFjhZQ9ng1OZ748tKn3
wmkXI0QHuB+diwrZiLD3JSm3/jsuY+OV9tBNMzib1dSnuA9Ol3mNia1FqC1d
DWsFSYZ6S47yWfW6EMhhsW3gDK20ZrAI8svLR/+uQgI8C+akg+HUEvX+78nU
SfFr43XxcgIGMAH9hLgCwTnLXObRdCrQR8sEKsuLvMPnYFb77IsSLg+CWrTV
gGyWHKQg+sIHjLrVrqEYXlct0d1d5XDLqEJVSshLd5d/GmLBBIJlcSz+Xvd0
nmJT7jD6JAGsu0M2w5ZSjED0JhMw/zrQzlWHPIlqVge6Gy2QWXFki1pCAGzJ
NrLYwGxZQLjLDL62OMAXllBmFPLedYQ0xZQUd2eVtgBiJ1GqF5Ch5HPzLSzg
eDBTe9d18q0TL9ZB0LS1ifOLsHyobbcP0lo4xqndeCo6qT7nVs3rldbPM1nE
QF+VGczp6RepFOqnM1yCH7qTVQYY79OR2hXCC5qCAQ+UHaAcfUkHLH1utJ+F
Ja4uOHUE37I82oTGzReYHpf0E9Nrnv28JQB3onUJ26HpUpmN2Xgfg7B8Na+Y
/UnZyzX4So+LVMvJPcIkanHKhhQAe5JZi5nRFxQChe209r/YvHxBzLiw/Cj/
tTnnfd68bmQcGp8Txtn+oIXefz7A07Mc6ys77q/41hd2orD0FmHYGig4AWfV
U7kZSL7lwBTkaTBqTeazyM4N3GOudj+ZOQoLyzbG5LPVyuBcDu6VOoHW+9H9
jjhwiVIqF+CG0IYtZZ7YslnMN157k/8nldO9t+OOH6A1O5HzlqmDLekA5fry
6NYAuPr6fGOJNTkNjFx6E3XSfe9sKAP6+RcUM2PyVDWauheMmI3QNTG20RJa
ULMyT+72K4d9W79tp7SRFDz5lv461JW+iWkiylW+3ojFy2q2AQIsq3TCMWMr
Sb71z9ogW8Jhdgjx+4c8Gr0j2Vxxu9RMTzQ4GCXM0WxZa/lshzfFWzJSBhUl
uhm9PxsAVUaTnRsjDFo3qYGdCHCBtfyAiQ+bUnuEpG772P9Y+DuqHNGxwMy8
lii5IGkxWO98q1hJkGNvnoRMRuvBiMdAoflXrxJBaDiPMI70E8kTMwjsSDHg
mb6/IyOizo1IWvecw/i1NRtzGY2X//qAEmrWOCf/GV/tfJXuQTiwg4vzvSBF
3hy4GK9jKt9wZzHdbpjdOFAwDU4QHBPZSTulJ+K4oZMSjWzL2fCI3VBQQwBn
IZ4nSwzQeHTgGCVn8L1sw60LESP1nYBiSD9xSBv7ZSw4YjElQGeZtS/uJFy1
MLXlEtQVxwrgc1YK84ltI2TonP1WM/OlzYnQdqCcHTP0RxMFgPCUf1bNBLEe
kAdgDfVHvwYQfuXPjbJtwLuMMkf/PUyCdQrFLi6txC6hlwtorJW7KAQqt7BV
ptDzRgBnsxm9AyWBSqAUzAfAuw0BCjPrWM0Wjwdkfcir6IYyOZ5gHh2Joj5Z
mn56qSelzk/jr+tCKhIjrTCYVtrWEYqk+T7AhjdyQwL9ZR0iYV52+tK/Et2v
8dilNPJRXQl+qN7nfywBJNbwzmKsAmtnJ1O/XognuGavwFSXaPwOvvOBaxKl
eJF3i3jZJsq2gGDRxiP6FZSnO8vlSomJg8RrLDjG1pVVKaBSMvI7qXhhdY36
j6jxSr/ia2OtT/aKkzT9p2rTQ2j0B+BfhI5jQq3o8K0t+KoxJIJoRDnfDqi3
jbxRo5P6skFyeRuso4knFs3NItgCyNbbnTCyYrchfwqqi2nJLQod7XqWtVGS
d5e6WeIRpVSkjxckFF9x0YIlZrtpcMgu/7y7EpiWXBD/IRXoru9+AM/bE2g6
NwKkrIRZkHk8IhRGSg9HUUFRI0bVbSEbXHQdKZ2RYU/oIpQ2FMgz8qaoiDYP
qtG8kxYNVNAqV55BqdWBr42Rq6+B1KafKMGgdYhkE0RWcZRYimCSNAEanbHb
KPIPGjWXAk4XNP9WX8XRqv636bJ0+3KbsgVxddqZxx8Eyl8VG7rRq8RdIDUA
relf+4bEhel0gPffuc730pRInanVyfkqIWhUvO1o7QZ8/149v1ztjLHGfagJ
DAktNw/5eO5I6qkkcDRcAOaTkbinBRT6EHI5urubkBYOSckTQ7z2PbEpIsFm
D4McKsR60ADuee8bbbcTRpidQS268cRLK7pIzFBoFdJct5p7Ct9esCrv2fI+
Laiwi37lcTLr7ZpJen12ctldKbkhyJ91Qe/u6RWFTtSQHPrx6WfYR69ss6j8
SKZ8gtAk9jzphELpCcliNQCYoyH7DpIMACLkw/2h+d1LsPkmVX1c4NWQnT/s
LYO/9ybIPbeRwCoOOeR0hHoj1Wp40p3k8BBrGJ+IfPIsL4KQhP4CX9gr4tfS
nl8d9Yh37EpYs/CeAlbqqF23OMposxsw4Q9ZzXmw2OUfJDswRT4URYwhcc8x
JGirFyG70IHU/uh7V88E4qxwdvsWlNpXSM3OSRsKHZ2ArxDf/qgNVMClf8fy
06hZYjSY3Zr5qkIwp1+OcjlGF4kTsbhNa6aecshHqkG4Et2/4z/VAJccZIwU
q9ZSUh3X4epXciDiwvDJ0WRZEJ8XvCC7LqTXv2oFtdpIpwmOPJBDlSaInm7I
s55giZkQVCX/h5eOe4si3YVXetz6imBCq8Oqjth9zArWDBI+/v0A+ZQ82Bid
cqw38uyWIwiiok9od0GPfNHihVH6+7lOI9b1P0W2YqJ+NpBl0NyVikxyd8Sx
OBMuW1XWA+Ov4rXVImjckDEv4sg3y0HtQPTeQzBvbyIAATFGCktfef1rh3LK
L8koe8JTsxP/xosz/iOegzcTnP9KcEGAeQOWoplBexp05WDwjj+96ngxu/jh
hHJVdvz1JX9x2P1yA2FK8Gldht77s0xMXnEgVxoiUAvQCVvJam4/oUI05igO
dnXOHXRKOCZIZp9eRI+nw6ic590yttwnPNFco51QbGrieur46xtMGwMf0XfR
fGDRtc4qQ5wY7thxEkbJDLn2M+JVFERuUEqxlZzrBFEjksssNUyPTRtnIp1G
ORBrQ7NuhZBpLeX1sXGNIfWY01T+r/KNovy3UI/HezYq4A7Z7IEEF5dIR0DU
g9Vihzvn7J4oPAPniY3RnWGPAyFQ/Hj4IazU10AzhvfxaHtp1MERxIDSSVx9
tnAArqvNFdRXRiM8DeW/8ba6q5ioLSjFt5eoXLG8NaGB4RxwIllYXe6Vn78r
Qpj0+vllcOIj7kL3afmXNITYNC1r8MIGzIzhQK9raZO1n+2jYuG9syqadDim
oO16keVfEbbX++Gj8+n6T7MtKjaaEq+iMGt4vngpC5bqIMgey5H1mAZ+g8sx
l0Q1G/LqjXFSGNwm03k3vg9vy+XsE8577egaPUlKnISpdsyt1BGrDkjN6gNc
b9mGjTYgAgrwh+kC9CWxYuHP7SgenDYSItpeSSvhMlhtVNeA8RR4H0Uf3V7N
YSvCyCCDrjTqxTrHPpezIB9UJEp4giyG9WQ4VwRewqEDag5vFKObxiaRQ6UA
MsugWOwhVOsZMPAD8RDXKxcuu8Bb+vhPGnh1UaPTA94pHIYLHOBCLhAxorPH
oSpNzGXZFwfDw+YVcgkTfhsScHQvGLjKU0ATWwBxqj/LKwnnlevJD9SZmG4i
Rk74+gHBF/gl40HCJLDJuppdCvBm1OA3Do+rxcTet8+12wQtDJ8n5RjDDmfa
ZMDXgujZuJ8JYg4LpKqxGjdN+lIHdKdw9rVYV37RksHMteSnS0FYLQu7LiEC
KLDBY1/VeWlJ+YbH3tndq++xTWjZyS6qt/Yoj0xLN8bmTn1lC2pj2Z2UIn6o
MIGrfFRTb1ldDQmfZXdD6+4JLHpU06T9Ns1m/yevIbGy1V8TayR+GoSXb98o
tPFWOwLT6TugEC4V6/f2t88XCFrItbPbAtp2oQ0b6gnt4/e2ojDeYvNHOXnq
FlVbyxXEsk5NZo9X4VP6fotV8D4YOBbScR6E1I4JaPI71XbsNh9wI3gq/OL/
M4vkUNglct+YbB7b1zJ8l4hHVJTF8gFvOU3qc6HEqLBhf/d1cdXArcEnVAsp
fVYgGHx3vHapV4/yK/Z7kTMfXMP/hOpgJYy/jbdiCJhVmaeFPGg0Bt7HJZzh
eHcejik2dksYnuNy4HexKP5EwTyzgW8H5gE4ij++zncNXIq0oam2+nHW6t7y
57TdmtSoCVuh1gMGK9eEUvJgOpmC9qB385WzZN99xWg28qFW1ikSxeOnxvzw
RGL50PPT5m5CSBqBvHe8P3bbVhvZwItJiNLPstj7EK+rNKI/jA6oD9wR+4lR
wUy3NmmB+yN11WhNLCdzEKO+DePaGoMerwciw95NdB25RzuMGPGpDFsfy9sk
I/hlh628noupQHghEt+6vnZntNuE8vhCWte3hC6l5bKt4HNrgy54oq9qpUeM
16S3EtSDlkTwn3W4ThstbSkmpZp7o6cyhOeqf9TJwZkL5xQstJaZduhkLIRm
IC+Q4pkXN11DPvvvmBib7kqkNB6UbrHMlT7ufuoYF2XUjkAeuTOGWQKY6ZS+
HxQn4AtWhaxk0Z5Tk/LIx8cKcKhU9QhuyZfTLUXSVNfVixxLKr8rxxhH68ng
JNtKgFD7eHfLhnDaUG19EQLdn7LueMq3BScNoCW0S524eIZY1nrpOXwYKdDv
4uzBeNikZE2cUUimDRoYD9aPb5RPJWFvvEq9wLtGwdRgbQzZIHU/tbSg3uFW
axu/r8edCNKmCReCoHBuK9ed/st3MUKLnm6B47FwBsYjQreJ8m8BJMqU3lXA
TP+NdWdShegJXK5Q0tjBQ2qmUhVmMjQE/NL7AuiAn8n5n4ATqf4KAvNDgs+L
jRr//V2PUswfJElotNjqd8jVkWgCyaTl2d8UduHXbZMz/AaQ0UMFZRT14vl0
m86hTfN+RL81eOIVx6VRPuBYSSceNIkgLrqaLjLdly11PPzWmH9NCLwjPPBP
ENAuTSi72L+fHt9CyKYcfPmXVYTOwySkB2R8UviiCWFgi3KLbpqkuxs9Uc8O
1GElr86PFHs0Gke1k44c2qkiVLxvWxJCg7dhhwvpRicEtBxH5Zhpg8CQ/Q0n
RWtBx/kUfAxoQlGLjKGi+IxJG6QPm3jtkJeqt91k2HnvR/4w41jqbB7MRIun
CzzNRonntMUwf7zruOJLpNlqJcaiQt6x5KmEv2CVNTGPmVJukuXxMhlVF5St
MG4JCc+DUx5hzYSrJNaJK4+OKAJSb1C3T7sgYP7gETuXHB8XrCDijVuchb/E
1NGP2bXTeFVPQt2qnglQsDUPN1VUveM5clZ4UWnfYTXWu8EgMPYwTisVp5s6
aVk6WPlFbQtuLpWp52e8CjRM2YutGqC201cWPOHcfPi5eGQJ05E9A8Oq6JWM
dIqXaPSpKXdQa2GRQjYN8i6AZlDPbBrN0erjAN97wy6WHF8SHDs0Va3XD8rj
H6SWOMyE5fParTkInqCjUz/+hYxLWkG/WiaTIur92tE/gGyoMC6Tpm0sl6dT
wuTiP9W0xqk6X12kYarIcfE0Dk7g3JYuTNBZFp+fp6kERehvf+5xJRPmv+ul
aQ1201acBd5QRWGIuaVzaVW4Sivt4VzCGUqQIRG+IVt7ahHcM5m9RZeG4V2I
Ktm8k9wk0rWlpRiWOXgHQe5hJd5w9GDkAOGOrQXFnN+f2bPPkr5aBtn6xe0O
MLqstIEzYt32zflGIYlkKuvva9AHduREopl2h96NzzTdxYM0WlPfVXN+yvom
lAQEoU/R7k/+G/QXjlieG5k4XpHCcwKKKWuR0R8cMjoE7NgbqVl/QtaMAe9y
REyBdZvjCW48Xm4iBoZK6IfYl0D5adNMZTx9yQ8qh/KlmxdDSeJ4AAY8biqd
T2JZ3BY7j92zGLOreMM/OLnJlMgCCZRSx2P+aMsQSZp523pWK6zewzKupVOO
n79qRRBj6eCg4RVFlJItLSq50l2a9NzmJQKIs0lms8nvPFS87u6MUszde0j/
bqLAal0KUT98AwstGiXXo4Jnz6eC9eAGcPLnt6XgB7Rkl850Iz1Ysysq/1Yj
eNZcto7QQVbnGkvsHKQukPx8gG0fZf+lad/JzyzwNJcXYXEUiGOL13VRtwFl
NJHu3cdHIT8dR4o6JnMU6L4Wv6wIg3L6/XWEbmy1KT5Fn4QQxCUFuEhaIzxh
Hu5dT5RBXOPuY0OFdV5PvL4sdOmm14tmqAPd68CGVHxrGpNMmJCG+JkR26dT
u5yPQURixzGwvVhsZq4LtS6SWgxZp0TJdmDxWoB036W3N3WutVJQ6FI09ymL
LAr6iMOlrrQbEMuIn2UYy7q8iHb/LnX//7Ss+yvc5fVV0mQ8C8CCUZUcJQwa
4Hn40m1Jx/SRNevlSuUZ3FCILg1WhSf515kRX3f6/+GC0py/V54jpfJ6DcE5
JmLxSaLZoqVOuvQW6PAvSJT32n5cnzndsm2GSt7rVrfiDLQVQFItRL5cka3r
l5dLT7AzWrPeTsfMcx3ck+zzLPTZ/ampC6v3UWYJA8YuV3QxorPXuQ9r5oT8
WEuIHa9AN8mxmypO9OtBG6VPOSxCsTlK2diiUbnoMuHLPQNv4/Jj8z23eiFZ
T2zNvulk4TWUAqHwwjWmfBAAUQQ11SJfkAmU4gSH+YstVM9s3stG+n6+1Knu
AwIhDyyQwgQe2wyOl0kaDK4vJ5LPIXlVwzqi1AkIPy43wRXk9RTnRt8xjqQr
rNdLhLZwMehAd5IJVbQUaoRBgHO+duNcgyKY3rkM5mYep9U9lsEmqrbO+yBO
1XaDhCsIuY7Rxac5Ygj+eXzYPZTQHQmaczToi0J89I/H13Iwb2JYA+Uw567P
OoQVjvyMuXpIz4UTg/gKZ6hDCib/QL6OMudwAbVQP92sSVKPXsJkHFz0fwKA
tT/kQR94K1ODjTw5S0YqtaICCG9DhM3nfi9ooOePh93NtisN+iPL199xtpmG
NbmcY9wiEFmfpc1+JuQLsDUITot8O1Ckhb6zqEyrhFugYueKYS9Oc0MzlrBz
tlohzy8qpp+Q58H0A3CjU6oYpGWZ4zLyJTCkxyMBUSRo9p1W7us9L4x/8h65
PwOG2sGbFVJWvup88ts64wfPRCm0jxGLBfVPA3FG+SfRSEJ3poXjTTAzuvj1
vTCg88DZ62ySLT0DgWvRnJxO/4ePcrfn/K55cpw4lB3t6Sog59RkzjFvN7yP
sfChUeNjPlPQEAi7UtSzdD34/1SpEhvkaWIgimbTMhF7c1DVkriGr5RnXxXz
RBaKnOzpFTfUQbk67ZoiG8YTdVor5EESEYxQJH+lgeJw64SUQ5OfNV1oB1Ak
9Okw2K0NlGfLWRijvNFGIB15clNceNjniiXZmXPT2Gdyqdn70nmm/Bk7dvit
LQIdjg9v2R9YNS/vpVl3Ltstv/IC2W+516Qcup2/2RD0AW+WassmB9f1Mves
SND+KFe5747ZisBwB5MYzeN1Nio5BPQ/pO0U3bzXRzqqqWSnxutd/qo0IarK
jQKsIX/xdaQfutY9wWWtgJufJGfMfZeI+c3+BgBKxuvBx3Zn5k7rz9MwMEYw
32pEciQTC8MK+TJPDnUvoGdfyXn4rBjIpbdB8Zp6yW9ukDWCHy09m2PNp6s6
O508jXxEhxLo+1PVRxMCh11tx1Xhb1P7kVuvH7pfVGPa7RH0BNS/Ni+cVsj2
mr3PkbqRo/MH071YZ91eTLeVNfdzpoJK1+0Ir4PoxXHlpeHVNtXi6k/EZIym
1+sjBLKqNsAjPO1UFOQlHJNMi2cCOmsphqHxSvwl9OrbY89j1W5/yKvr0aR4
eR+3XUllB+WBglk8LBo0QZHo7inOCCoQkk7NQtnqu36SOa8vdlb/tFQ8ce3E
GsDj6WGJsjFvj4duPY20OvldN3u+gPzJH2VpMSepWoeioIBM0rmvdv9egZxa
GB04hAHVX7hADgejazWd1o0qu22uB0mh3xVXkSyGO5+4xj+rmR8fr67N53uF
FcmAGCxMuWHS8xGZl7dnBZr2Lf+QyNc3BoKbFEUZJG12N8QOpAdID6SQh3aS
FroZraO6XAHaCxjFR5OTtzGKzfjsqw8ypPqR4HeABRdp1JnxUUWAM+QHbVbs
zeceRLGizPkX70Vn0uP9cyU0t4gIVKWKSxoTUT03VUfgpMycqK1q4zT6ZmeO
pVf3YsRUy9stfKrC9YKqijYD4ieiIaOHGq71yUgMN778ArzwBsNSC+tH6TFo
Cjh54zBjaJR36NWMAfZSaIvqtUHWYVEwqx0KQEZFImD3hykw8PjPZC1zLFly
L8IKFcY9L4ZnDhTi929KPWZJ1cibOljcwzBQQsHPVkOarNJOJ3M4tINAEwoQ
90sCqVAmFNFFqCDlay6ZEYUzBW+c4oo+PrU8dtmL2YWreJW5HGczhZnF8rz7
vD28iuL5AfW9aJPMLBvgkuQeOaH/JbU7qiO2FV2r3qxdKyEj0EZ/DZwemD9r
Q636GqI8V8Bic4JGMtBqLgnJ8BbBUNfkdiodNqxEyD51L8dKbxbWDZXgjMfr
o6AK+xa5vCrSeMQmyZDjgzkpoJBjICMKLIEkF+BZN8lDY23O/WMIF/XxmbPE
wdJX6zGQ44qwTCQhVbQzHXkyk2HsBsy6sH6B9pih2pwP7Ju2XFv+Ar1kQ04B
31IlYaegKYDkATrTefp0tygpyJjEka5ghL4yvZn+vZqCjWRlVzgmw9n+33Ta
WMXrHph7rhWVJhxUJMn90FDf16cnR6FR/IVtrPzsCjV57+j64BwYTDtuiJ2S
Zju51XB/jqE3q+YGMTirmvSSspjvbOgFPr4GW2sAjSgwpMbCLP5Zxvc5u3Sz
gt2rE/pRaNN7Yn/E4ScB4RhjGYzxi/70MfGCMTs8tlxPBxDZZnXyaWXgE1pR
FAlzl92AWvszYO4J0JCfer9wNn0OyB6hZobwO7ds2MUGowLozgMQSjMUuQNu
qzu5L/aKcZFZbyEq/kAe/dSKIN1usxCMSrJyCGdH8F2JkSkAC/vRhUiatiY3
KmLxX54XcZ6pgx+n8JahrrS7aBNtfDL9TYPUv8GRZyXkJHsfjHkQl+ohFKKJ
X+uxtbReWzYci+PALS6JdBrkVN6EBQbErlPzWG79cvNNRgE2o0TNjFfOtnEQ
Fa4Ogx5i3Ddvj5CRUBK7eU2w5LdK6XfpSmfaeJHy+iXsxnBIUoI9Gn7B1Kyy
rrGWGtzC57xd0H086Up1yGCtLwLi4wtzg/cf5t1lZTy4NG6To7LJ8fkiAff9
vjBAtdSOdXGt3qZjqWzim0wq07/SxZNflbvlnQxdf98SnyV+n5faBQ3EkdAR
DsyoPf/jU5znYY21usJWND8BxjMnUC1Ssofgfm6kLk5sFjzRbCR0RQ3jL/UL
Y2g/ZyXwGeJqNLmzJDqB7oQiD09kX4aA2frRJz+36wT/x0GqZUzSxqrXG71K
lo8DDPHGEcH3uFTb/DX+W4Dz6/UcftCLsZA3uZvedRuqz/coaRjgQdImPVip
kgYs5IzJekJ3Cas3kyJFSu0yHa9Kxq8gQXCapXOY6rvla0H6j3jcawgEssVh
7gIJMjI6NPPtYri7FLsDzNBr3XMXrihLgRWrqJMk7VhKRaPK9ify6o4ghC26
H2MO02FahmflnHBZ4B/AyTjaxb5afj2YliLgq4VOaUY1eFJGgMZY+0x5rQlh
wdtSf3j5bJFPXDk3kpbnksLH7jE+vZi2r+mAdGBP4m1uF/uR9jkufWyicusQ
iUO9DjZwsDNzzndbKV38ASa1W7AeNqpOvUssqL6yVKQSNFQpWCSjLXBvel3W
SU+BYqMYcvhuVMRr1ENJc/Omwu3iVTh0FfIAjKnaZn1ug9tnOKWmKXBOv1UT
9kREVOK0eDDWCn847ycsmGzZl3Lp67ccyN8uBUY3QuctgE5r91pKvahq+Vh3
uwW5B5W7+3ynY8mqxrNZrzXviTSNL4AAnZ8STJBSqcL/MniZeoc31C1QAxw0
Fj7M8hDVuRrIsEGr9emAyRD6UnhmHV/8ume9XNgJkDMulqKNEB2RI2ZF1UoI
5GH4C2XAUy95Q3qOHcYMSFKYhQyA/h8I2i6+y9dUtCD+5fxOP/M8JMgpaBXy
K0PDkc0XE2jjuN9VQ99Lu6DXSIbGHacKxLy1JaEzzhqwvv5NON89qwCKTQ8J
cWo5i1hRfu4E0E1y51P9hbtugnIPhioSDAcJTKWZRXqzdJs6WQ49P+5VZ1NI
HeIJLgE8AajrHYXjPw2puS1tFrAsoTwjotDA+XGfDmYlvta1IPubFq+VWkMC
vUETjqD1RX7MHE0vZgzqUKRAH6YggG5hr1Y4CIR1DPg0NKwWzC+/iVrKWByh
iRdpBlxRPCas0nhdbDzJOnraLZpSW33nBFJKHc4wOQHsUl6MrUuVuGOb68q+
CyhtH2GyKEviyKZyeqm08fGZ8Q+BdAZmCmvVr7CrqvZrITK3Nbkig2o7ckVV
ij+Qj/atV0fYxTvktMpGHcNZIjhi2LLddRMScHjKTkeduXPeDnoL2Wao7VTP
UekXZGiKXusiLv3yGH+o04j8dKgBJFlEOWosC2w+eBTuYRUOXRLT45wCTXEG
/6iBb9aEtEvoCMWXbcNb6d7R9QpvM2dS8Yqf3rLyxGn8qJJ9av/oRdsch0AU
V8reVdK7f7YXMZSjOYobpW+Wtr7eKKe5NgZzJea7mpL5fRJ+wh3C68phCdO+
ixlUTzsWxTQxFUC6F3gS1fhCh7kQPp/QubOrC64aoK7aF8DPWwO7VXDoSa8z
Ry6JEg/XIj26B+Xd0ehi1QA9n9waKeIaGDTR2hc1h/UxXCEJ6geEDpa8gxj0
TNNaEwAuS9OnhqPKZgVyVpgd75Z7A9rCaJcWABE7WD4w3I/6BCJuhK0kzX/D
/RKqiit+gHWCn18VpUabKUuN+YhaE36srXYHJvCuaSuiVajH6/iLz44bPWj/
L51eAt06BiGzna4+s9pmBKE1yKMltFLh03IHJME/LT8R03PNHeIVU5NIAfJK
zfFjja+QU1YzklO0bw4oMbBae0ttN8mUDq6QJcnM0l4w8csiy7Yf/oKG+gSp
2Rb/xv1+d0Vq1XNiakF3NcwZHADXTeDOjAEwZ9CanJjnb4H1+yrIF9sQCsn3
RywO7kV6f8m/84/SO+HMKvg+tFgqzNb9SSPzl4tvlbFpiywpoNyefBhiFNVA
hIEU212P5kwY2F9rs5z05aNYUVI/WLKpPGpbnctIXrEiOEIfkDIl9sbwfh/x
MCQyO2f3wHRQzQ2JdgoYBD1KEFlkZVArKgAAx04GP9crn9wjOwUznbQbhjJs
jvJyWTCv3Ol0iUzlnokJuvYX20xcKIyI3RGVb+uTJ02PofAqZu0itLDvHavb
g9nFMjVBZ1+R5gGMMGDFppIfz+I/GuAuaZH5JF0kr8ASos5XMDVOhdivD6GI
DEhIyh7ryWB9vlHIXAJYckG9K9e+IABTJAsKgaI08/jh8jQEOI64SYaEUdgW
KItxE8Bn2B7bLdP21ULZZLuiZRAp9nW/pbTHBTP4uDpBhQneQkYBlFZe3SCT
emd2qELqTzsHUkuCh36VFZSGhtXBSYrJa9ZvbIJXg5jDtP6ckCkR4Jtgyyh/
nHbp84SbOO2g0Y87V8YJ/9z5o84wn/TUk1R9L9blC+6L7Tk0I2LPAMUvLLX/
JNZ5uKs9diab3k/aL7ZOXpPth44Gbze4VS35MyGL3djFyfqKl0hyvC4NhmNA
RYKs/i4hewixnRCA6Jjnan8xZjizvFr2ZeNvNseuShRbReopGAc8IbVVwxOr
V4t6OB6onMj69CO8B8wpoZeQv4yaXg0qVI5vYTNlEQzg5ncHQJnLS8y5BUEV
nuaaKPD7EfBd6VglJJAkWMVkUW93JPuHi7CxApVpjIc7oUXELETw/0KhlmSE
u54y9PTrslMi4MOuLVziRWuMw7l/4lXQ9RYO1VyckSo5sU8FNQdWbVgegEw+
LgDeQLfBbXD7LKyAhVHMfJhw2nAfIOs2pX4DUmcs/8ozTcsrJ5Y/b6FLQrvt
FU9ifOX5e13eJwDUFi+guCiFJLCx5b9NijsIzkv4mz52XOFRRqW7g8Pj7/Bp
r5vAWFnOftmzrQbMf71T55xKd+ofyC9zLNlcDlHStadYQskQPpzjwiotICf8
T/NotEjwxvsqZ2GDniqyTF4eTS8se3R9IEeYV8i99Ou/3MoWbl6L99GQ6NA6
68MSVtQUVNivTde8JcGyvgQ6yqkNmBmDVf6Rr0ghPyOgbW3McvUtBxWCRY8/
IBF0NBRV1OxUsLuNvv0MJccxYPsudAJp2i/ZPzHXtA17vcabzxhxEqnewZ85
pSX0vonm9xi/HkTybYkU6nGeuv3/Ii2bcQFPYR74bqPoN4E4d9xAWKCo6osz
5ENg0D9j2UFhMELPRKstlUpLpDxMJqO9zf8vyogTNJ7irbSCvblo9A3kDKTg
I1BNuPakQdKF8brehMPJsdx5lfzd50ZALLxbNoyzz1RELMZvbCHmEBV0mRK6
I/OGptQxFn0Ofo1da9azgf1SQuGroHmWyugHy8OmbTISBNpRb7Xm9+xjG0jC
RvewJ9piHtsGbeuYwgmqZT6QhAVgsb6ievlQSWPXHYuWxlAe1bwP+vH9kxCX
eo9kVJ8mU+LpGkTE4oz3oUuIr7wyaD1OpwPKfAQGg+uGLM2jFs8WeEBElMCv
YFAeLO6LS4treG+sno2FCnuJG6Kp/6nHRRdjMWDS61GYULt8fKMUI31PisBb
JPZTFejtlHVn4M59VjBJmvpwKr71J7YNi3zcKSz4mxkHRfQwsyeapjXGyevN
/OaDG22xCmKObOUXQv9CzFQ1JIb6xm7mDVg3MqomAsmTFeDbInZWXEYUxKh/
dD/aaNbkg7YUWQ27QmCPhNN8NXL9NKQJjsn0Xmhmnctk2qwZSDdA1huYwNjg
pDhSdPb5CL5L5i1PluHBUW+ICkIwjYrRlUXFMi1j8x8RcDYQkFYpujqW6Pdu
qUsgxiPJbesWhQSqvc1tF+XEDK+zjaYU7psZu31V9YxvacM92nhsuqthuvd1
5fHkszI5Hei2LP8Q6OhzD7uaXEdQh17HZLyCF3+xfARTqXnOJ8txIwvqf3hZ
8SmKTHBbysSrGcZ0fL+shX/0wzQMJqQTDzlT/IAlrAkkt37Dc75M68PPvBtt
zorl+KfmJymhoYITo17gsW2CFUW441PPiQJjG1ebBlCzluZq9QNMbMwPNA3j
6ZWAoY+lvfNUmw82jFE9OD7zXZeybi/IDw40+dY5Rqto7PnlEsDL9dQYe6xz
v6HZa05ZsmQSQXiqo8a6Xpm9bIpU89FiuPDP/BbbUZ/VZPF+PHEg+MHd7nLd
RyPTwKQ34Yhy5zdIaUuDbZhj8+sU16Bl4OqDBEPPWJaAhwlYc7tN/3vG93S7
+DayW1YsB/5FkBDVLP3UCokNrIYlnTi8roTF9FYMdDR6juzukDuS2UL1rx3m
EItWbG8WA0hVZ5i3G+Jh6FqYZ2m4Ab47zmB4xWZ7Y7aJKcN9FBRagjOYCxv/
6i6IGA5QrLAXQR6Ds1D4dbt+IwjZWkIVTtr1Jp4voqFDgdx/8x10KQHcjTpp
rx06ZIAQ5QQAI2tHiLIn2FfTQEOdAp72bi1s89UCPZRVXbWX4hDt9mG9dpz7
CUO+2RRSAzf6PPlecQdZFk9mfdk+U61xHP24m3/LVV3A1t8ZTZByZhyBwn1k
UDLuARshyGtOsUzyBQcJ8kStHajJ5SfNijgB6ja1LZmg8V8pmUdI2nB3hFZQ
7l9LrtEN0W/QUbscQ/j0TDglLNXUkL6sCag+4I1u1GN9aIBLoKTZpkfBeelh
g3O6mP3yJZRxuqeKUZog8Vm9VyQ9rIcOjWFUrkZEpJZUX8NzPgY/d6zbKN1C
jutFmNG5V3V+dVybls/Hb0A/KUTrI8kW5CfHp3FlndPWjG9sXh8dwieT1l1s
eZGZN+JuN5/p0gO+JGWvYjZY3F+e4aB+/tIJXtEg4YJKMBNLyhi8rVG/7XQu
+xoiq2xETKUYghJWPbtHiLGRJTd2wWF6P+S4vPckdR7HKq6tHkAH2HiM8ajd
ZK18WEgl0uv1jAUPllwLbFBnIit7MPrLA8wfpCBVJtb2sLRQ9ZG5Im5wgaLS
EUDw04fQ9fz8bvnEFJ73iCePwQUDQ60DUYcc1/0/JftznZ8dqnXUX+T3MNi9
hgUlf8tilqm6YjiN2MsyE1ry+8Wbyv6ZtVKVJ7pw9dwu2eCorEZzuq1FsAl7
p76+1B4bgQqvjhERKXhQRkBEtkEjG0qEUPPODQEr8yx+eVDnI72Zytahs+5v
K1Q1i/yteWruRu2CxBu1akajE683nHy3lZy2v/obV50Fq7PXB3DJvUmzPX50
nvJdvrjmwAG//xru8fwrqqouuZL7oGbPD5Gj/clO9cAl7k8zQes5ZuyMnVUP
v5TsgJ4a1/A/DC4OmsNxKANySYGw+XE/r4vjF88JQvQKcuomeHENVKeYM6LI
zyF0Vunfcc5FWRJnWGwrbrJy17gV3DyDur23i7LM63MCMv/ksPXi4GvXeOXs
PpGpCNjuIxOgrnfBt9pUjtGjq/Jtj6eYz0rdE+frEm5ptKXeOFuvrKCGDdaK
UkGIbDhjsQK0+0k/fwdyE01CTFaxdAxDK1xyGG3Xi7u0/F5dsTv38lKCrOYk
pLgOk66FaY7aIbcQ83UOJbWUnoxDtia86OSxuZjavprd05yUdOSz8SXrqCNw
NCD2NyJwWh/Z83zB9zbfxhgjlZ36qdZFi6nuKAwtSJN6bs7VFNmEcedScF3w
Db8vT+IjUmhGRSF1Kwxz5KfoKCuOgBnu9jpHbThEU26YXG9NEgM0XZtCVo4Q
xJcyQCkyP89eulDC3/T4Nbzjj9IDiAeUDAdDfdwpdkWeVSHRp1srNIDsOg+z
cCm76T3LCE7eBAzl5XVt4IXwFrrK/NkqV5eM2oQ0QbFcEzIa1bRj6ITeDH6y
SmtNIoFR9XSp1w+FJAmttCgpn3T4JhqP9zxSodrTbvqGQu8j9dxVPKWcqgHc
RlwWWilkb8prvA6ddGmIHcLVZ2GIMvv/xpGL1fl0tzdsbX8e6coQIjhcxgtz
0KhA+BW2Y3LnKS800sCCG7q3TGXZKEmDbFnScSXvMATyXN3YOyIhaM/9ApXo
f9ndSlOn1wnbJ8w/LO880mmG0KJFDaDXaHRlLZC5sFI852RzQNgkhKL6t5Fa
s1SEfAfGat3ffCEUse5y6ABhFyoBy/rglrh3K9SHQnBqkds3uieGjs7jptro
b9fOUn14SfW44Aba/PMVcKrEIdXHU6Ybq4oSuOF0JYWGYTfW6uVWPhLB68xs
XmPDw6oA+YbaluRhhumRh5QZ8BksXHhGnE8bR9RGQyjbr/BMv56vUrpRGSNe
hHQpHFbP8WImE48EcWy2R4Wf92iDScn8rZ5++o7Io3NF/lp3uyDciJKIalIj
iYlOdkNakbu7AMg6v2EYQ9W2QXVnWuZ21L12gFhkFxEJZ8YU/kMWBN6WiQ30
X3IqnF5Rg0h0XaU+lRqkHy8F5PSukDweCLfVsmyrwh33eMfCPzMO5PjuAMSu
GO6n4L7YsGtfa6gozb8YGvuzt/j3TAWH4YygSOw5QPER5Yk0CAM+98Xop9DV
C/lZxu/jB9/ogq814LKHNVbDdhPRzkeIp4JNnA+2cs8RdH0Ur7PWLy7qfs9m
vw4TQlMzn87hzmv/U1K+3tdYzsuNTNseL1T12TGzCA5tCvfpDP9Nr2snvQot
kn8xzjC3BM56sUfGGdLUr7dnkwDzM9X1MrsefT6tcd0FTtiFf4xUDAu/tTso
+UiFX2U/iR2lUznYqF/DeSFlEpnkbXHYnUfT2HMjpIrkVmzwOecsgUl1jPtc
gAffYmLVKi4pgCaC4NhmqADpVqRQ1cFMuhOvmucUjAfmC5YBSbLTZ8Kba39V
vAMWEAQQU1Tc3S/BDhek8M8+3QKSRw634eADkfXpjS7p2GOl5HINOnp2EAPx
VBbAIRQGZMS7XJxCUUAGyh6CPuWvV+uctv4Rg43/a/YamWxL1erxvNwCenVn
YReX3p/jWjEQTvEzoh2ZVi9pRQgePh+v/VieY5tWu2+smAgu+YPDt4Hzh53V
x4rlFhsTEX+PA8PSsc884r39Hxi6oknPO2gWTN59DNbCEO880K80nadBEhGM
qUWtg+pWdHb8sEt9o5fhJRTALariqxj3c+qNIlALHzqButL4z6tKOb+808Y5
A11JzhZEqcD6TPBDh/Olv+JaELU/GzKfNkuF6xIqm+LzP52nFb8S3U2w3grO
bAH9+EmknqZXMCRdQy6COoRyq5RFuwPruYNe83WamMQ3C9G53jb/yBPh+5T+
hzluZfBqnfspSUmdeSyrk++i0re4O7PSURu1HuXQi8InAGwQogeJzqTyesi5
WvDtA/YudmdytvbV13Fu9FIcRVXLybFd3xoO0MYj+8I0OERzmNini6eDm95d
vrB+f0s9LOnUwDGEK6h5ovAiCRCvihENiW3BjJ3h+70F+fGiJ23UCP1AugdD
d+rtql6N6kk2g3DVZXuesorQ/BPhJAAJra72t7VtVPYKrKFVzsNnjjOwgTvJ
DnVQABaFQJFyb/tBg2T9Y6JKZtVkLFPX/Z9dJdMAS3vLXmt2UTEneBg84aL9
bo+qt+eEeHbz2T/baVN2Fsd1efFXv3df9mhnMXG95+uoLnZRMTKEqmh2QNjY
xAZoSPDDaVKyYzKxSYRwBWgUfidnLBUlVOICX47qz7J2s9mJVb8p6lAt4ANu
Vhcv2M0wTFcuYHKHMxJBUwu3O4+UoK7ot1XZrzNoUnbMZgkD7DYPe5yo0ozw
NTNglyswjnIlx5EVOC1LuHtMJU3531ipckYX0wAqVrWudV+g4lZd6sZkZOEe
e5jjgtmUaaErO/s7UDni2FnPb9Xdb2e9GZMwuo7FR+hF3z519UXz0/KVRuYr
hueVySVwMC4YtrYrse1hEMZgSM+RfLxBQpUmzcS+9DsZxz/ggzxmFHexaCKd
xM2oFn1Rg+X/32mh1bzeaUoCHFgRqVajr72Ok6gLLfAC3CR6/CdvnwKrhBc/
jJoj2WoKdYi7dybhs7P7eQAOZ5kodZDmf9Mc0VNxCiJgqCUO/clGnbU9uQrH
LBAK/faKQitpAJwG+13NMdN2f46xU4Ja2kCRWvosjWPbQiofBWuj60i1Jzrk
/rAYvpd9/c8Il2W/YCySZK6c5iuDmIfBXHC/C7NSH3sCRw+T0ygIDbjdbLQo
fvrOaHwfGtO5+k2nJzUz3oYq4UOeoqoQXycSq5Be88s3FOE5km2/IB1NyeYG
PMGaYFLCPGRREx+vFvnKTZzkxU8GuH20X3uR1nIiPRqt17TU78eRqLgvmb3p
ivxEoPamAPGdWNZOf5hMEbs/Wpr/CDqmwTjg6BmIs68mk7cNuojMTPC5LhMH
VU15VI2HbhNHHQg8Gpbc8yFx8CdoyiMhmPJegd6sJ4q/07ce6b7wrCdVEM/u
QStNqnPPkhmHY2P1lcJjmDg/YGxi/S4trrfeAvHraa5a2zP8MEXya/i2dbxU
pl6HWTVxl6k8v313ocBCMpJjzq+5eB10xg0RlHd+6mLzUqpsvspNEu8hM3YB
ebZr3rf2UmVIYZVn6jmoQvWxUmLWOrrKnDM3ohIQwgbea0PC6ov1WfbCcPUQ
D00fXdQ9vOdLYm4WBOKGSEqMBC4foubq6QvpzJlg5cDnSdvZfnuaAnevdlgC
1HgsLW9QSt1XpawQaa+nWLbiS5J5c7R85F1wONeLCAf34zD2j5jkHf5Eq/4o
KFiyOXn7lQuKrKrm/MubbydKfoDPJBMYgHcDqd4HIo3tpcZkWpa97G7p6lE6
XfFDRMSX0owhs5eYYSyJC8BofeDRuTOfWyiVyUywzwpw46o62oWqxf0fgCHs
WCgOGNYSdCS9pOAmADvCWJmb4PwCfsycyMqj6UFU57JMvt4HGmUqR3uuL8w+
E9kwj2caHDd1dmZQAo8ByyIVucy1pw8tVwYZi6/rHDmPgsHB0a0X1g0gG8N7
isZrf0GXLRBXslk1NgS7UoovrXLn4xRgsUvU5+IKPfaIXOecwuAnP5oOhP1i
yPTpG99HZoy9tDwxWn9ZtkF3qbIrXvmEIqgUR+qejT/FTLPkoE3SPhOWr98X
Asz9IUWLUaoUg74AcjgCIA5rkhmmEOW1P14/T/swQlgKCf4Uv86utEBxudLx
fzFuXNrZgtYZfVAYEgrIppTKWT1d+/tT9dpoPnFRWzFSYf50grWlWq+vhrcI
gFIfRg+1rNgFWJKCYHWGyqTkZehYTIt9K4CF2niV9LzpRt8Xj4+HJnmEZ9LB
54nu3vIKRY4SvGzPdAEjhK2zs9goR8QQ2BhNkUc7e2X+lOV8DzC7vuOjXHZH
o9OxX4aupzeJedK69vVjQnIM9oe9E7Lr1P+VpjNGCabwpSJcnkG6roJu9aMG
4ydmPAJkqlZEJM2Quv9Z/306YynP/inrakYCL6lLUoh6jqINvK72XCA5ZNOM
k7fVyvM9yHXnU2hbpgFerV24ZG13PeypjBxZGm33aFZa3WXMsBC3TKc1hNvG
Oni5v+dUTHTw+PnvvZvS5hlnsjQnn/NjKRVqwoIdy4Fo2xFfv2oQpmU0oXra
ttNBlIxdOeMJhuYzQepdgwWUu6Vdn4Bg0d6xynDsi2dTsH9Cz5YpSRp3KR4w
SMEuYY7JIc8kngwlg8YpFPQiCWrtP/vPw+x57h3LIAwF84YGhylsSnf8q7zQ
fAAZaawsKiFdWF52T5YGgjYySNArI6i5lEqAwFEdND3HuF/7yFE9bh5GaxOx
othti8lQpm/khnntB71uAswlyrGp5dFNRc12lnXdSvcO9feIg/MrLHGdqMj1
ka3tf2iJ4DwMKzmrAHGaGXwjx9U6a0lEHgahvCdpZBdWxbqJotRpSOtIeUil
TSrn7NhHuSiy8LyZrhBpD0ZflzhcSpgk5K3qAYzcjUsNI0afd9+cH8GpPXNQ
0uyFrncAazzFIQzXIn+g1obIewiVCaAvuKI5gyrsiNh1B0/3Cwy8yyOzdqe6
6vUpAA/M8fhh5cdWXL8+X20iPHa+x+KD4fc/erOW1BNRmpb69R12wigpFF3i
GMDhASECpdnwkO1O84T8Q0UNsmcTnex+6LYwGyHell110SyqOfWq5steTmqK
QTbCFRQRzdvs5YUr/oLi/ZsIS/YSbpPLvteqH1dhwzbtBUYE2aH00dvpJY1/
mVcbf6jLqjPzcWrfohDR22dOe6pqe3wPJ72uAsVoN06Z1I0WknjI6PAqlTGC
uNhVFwV7fsU8gFV5cfvMlPrNaHc0CFd+Hu6KvKEie7hEPOJ58GvtbYDzXpg+
m3SUMgVAYe0DiDYp0dnMpUlrmgnpwssOdCnSHgx9Mp9CR11ehG1Lj/2XMVZg
HF3BwW1FEs9NoNSThGc8e1bIgQUCFqEvLOrpp4BcLsJKxoX4bIuu/mIUshXz
XRHJyNpt9HQKL9NOGEeFlohiid42hcvvzut8Qg+X7p4osTvh72bbt7Idmv8l
Ci2RcvJ242B6NWVSBn3DJJHXW2vJPewhhJTkxgeDAHYjNEYvE8Io5n40QULf
f4TWC9WxvUMvFv/i/RqmwDGxZJggi07u7UxTQXlf11hTuMPlplrq0Pp9YLb+
naBR2TJRdKC+2iGB8rSQawiVbceEoy4qcZylslL4cjdMqr3r8pVIO1vN/3/7
GOoD6vK0hS8f+3EJxIE1hNJPSggeslZzXTUeGNu5PhkGjc3MjNwykosGb2pM
o7OXvLyf3lvoJ+TBYy/UnlRQQdy04oroU5RgZoI0DvlAU5PsYIb5Sm8RHARe
4kwanBsJ8YV777nA9lD9e5VILkE58Y9Z7Xqf+7Kq3wF0UMJxaId8SZvv6PX7
SDdJLhBgQcLawxQlQyeRstgERCX7PPQ9DpvQy8Gmpfx35IrzwHRaHkgIe9mH
2rK3JUQ+7SXV254P7cFnAnJ5TodoZL9yLqFre4l/VGeBRxI1QKDEUyPyr8dG
KLPkRB4vsY35ii+NlieAupondrxzxA0kbCkvYcjSIxSVNLr52Ake8Fr09YaV
V1fLO2Enuq/Gz9pY89I8jnrV5vxWlXVt1oWOam1C0ZIAs1dQvXRHfH65gidE
4eOhrK5xva0U8Mq9GuektAjee21nEGUrgiYMNWHqmWZvSVjQ1SO3YXo1O8E5
Z449C0AzO3DIEaUSRySdIwhhmlQ6dYS/+8viWHAN+cykT0GDnIGBn4AgvPPh
1/RBF0VafHHS3Keb083nYbibprSUIzN2T8RqCsXMRg1+M7mmIM09iSxPdevu
LF+cKEtoNc1SBtAid14yquEXrCoKg7RYx0HOxJ+ApUwfhDJwXeDZwr9Z6Yxs
R3Iv8qfg6fknap8PD26VUaqGDaj2aoES4YmMwxKrGlI+QSH/7cjdN2Wdn4/1
R3d1uAmPp+ScxLI2zkNhY3AQKzHus1hIUTWxDz8KSgrmulnbZk5X4HczjZzc
ed9EoVngY8EPZQKcwv3DSU/ujLiJpLNbUV1ZB/4JNlOclgnxwYsbY+1cVdKj
oLVXtD8Cr1RUjwJh1kNX+V+bjxLdn8mKCgKWPq2KJeLvlq4BdMdPc7GZ/z8M
EdKWCS3G3Hrz90EsXOQapSwSDPFsDnRKnCzDSatxKIKOv54QaOgJa5kFxPZd
ywOLQli5e2h3OT/i3+AbNyIQkbjJ5bRVwSAzEpLOaL70zlOLqWAxouOKzwhP
p1vTizb4zKmjwA4RDtlPlFMamGGs7Bm+x/SCz3bEvEdc+baRg51M8rGmaaWO
JtxHuwO71pNRqRQpSoB9u/i2H+TAVyyXWYfyhsTIZVL/CpY40KmBf48nxDyv
U1Y6qXhl+2MsAi12uBCtqKlszA8BcrhyKxmTMLLsPAMfU2fvWqG2dYhLjk4f
ls+crIUsIn833g1z3pYXrepW8rNHdTsu2E2DjYqcViEiH9pLN6hQkvPX4a7O
2a9MCcHo5Nfaa1gbg2eB68c2uGmaxTv5F2GnZ/ucNjJbQJbSoVtDG006sJKD
I888D2EnX5kSwsykx6koZ/pkrAjTOpNgqp/OGO8KUaGLBVWsp5AtXrVHKHW6
MltrUUApyLV5jTfZDyr6bxHaW/HdCOj+iQ52lkF1v1ZuurQuHizYTVFswhwI
mOE1OaspI31/emTzw6kaJ9oIxuROfvoCnNXHC4Httg66HFqk0xRq6HY5lelr
Dkyw0gdIuSnTaScummv1YN9eysS34GTDBZoZnooKQy84jFA77IxqSNif0Xyj
jZgYhs8ZAka4nKZKqp19hHzxNUtJEqRk4fIj8D3VPNdRQuEi0WZiH9XYzS2s
HhTkrg0lRIMa7WTxY63hBSZRIHo2HZe6OxuX0BpWnqBhv90M5dnvNjA3YZE/
8Hl/rR+E+h77ODYWeewyPmnuEBzyLKsvovNr/8A++0jZTmMvu9CVgJx/OCoL
toXMLG71hbfA1vp1g2E8qWjQ4EAiH1q+n/Zlkm/8yN1ulqhpdINkUr9wFPjn
0gnLKGzfEOVehCztMcyJAFxn37wvQKxQH7PiMTNIMDGZFMCroVHtI8NqF5Jm
AYO3RPpmrilE+d6LxCC2XBtRdzLO8oxixpSydPqiXBREIBrgVQw+K8+xeBFo
AVCUrFvpauF0cLBN00ADUiz9x9yiSZZijE1OeUtiM3GZq6xcsPiThrUKpvyJ
NetXRRqzdYlP+ZnaJ7NFIml/paKMgYp2TD4NNNkRiPhQlC0jynRHofbPc7Ev
XcZio79PM+tYgYoy78jw8aeIMyNuoUQwIiy/MowgSv27X6/SkcCvN4X75MzJ
JLLquXkh/rLEbj8dLTTtkwCO6FxK6cjhrz42M4FIt+sigxBNzocvmsSQVQwo
DgFqmgdBwiiNePPA23aHL3bBxQ51Hd4mF0O0rw30X0dMA/d3lM1ABKz9mqS9
WMgUOwqB7TO74b4b9m1bp+hzz7alZisSsnZ0rrONlaLc6rNKF8loerWe0+AB
nQNRnOy592sO427T90Mkvvf7LuG5j0wrxliV7Rms7re2zlGwA9xH7RzpmYFO
++tZBeGbVhVjeo0tUT/pzD3nXOaAcu4l8+cJ4Q41+SGVF3/yQe76oa9y8NbK
6uznRUl2nIN4i2PHjimgQWKja0ff2vl8kSw0HYl//puo6w5s2jhMtZZYxp4B
4akP6bru5ATVDsNV816kw4lZDZMpiB1v601PttzJnGaS10xmf/hJhthYAsHN
KggdmW3GrWSeDp9IyyKNB45sDUxjJd7UoOMox3F/h6A3EUMoqaVhe6LOzu7a
OWmwU1l6hmfi5h3B3OLmF3Fc2IvWm+y0pAGJkuTyBpnDMx6SjRclfspPZTgf
NjtQ8/HBP2tKokybzwEU4CQgaTZzEn//2W5T4hAt+9w7s6sogaiGyo/JdXEm
m4bFfmqVStEacZtla+2VzvMwADPgiob27Ys9P3lrCjkkEE9/FeyhgpMk1Xje
EBErOMcv5Yv4kRYUVDp1WljD0VrN+bhtXIupX+IgpKHyu82sOIPHkSAz/6W5
59dsNdP+/e5hnSP2OsG8sXKdfIfr4Q+ntstqfoBLChey42AaZ2Yit+ywccMP
QLPjVwmMdVp16/n8nnYVkCPgVtJcrLAZYxEBKSrVerSpSTs2cRdiC2JhSxJX
RLhdqWB+9ZxlyIDMK2N9cAnxTrNRfLI0k6IjluR0A3XJZjoGMdL7A/fPrLiQ
lYPHqyeJi+DG/eqffYSUPZ0LS2faVv1upbiK7bWqct3JYIbXGIqF2F2IWn3e
+84Je1f6TnMiKpnWxGrO/ImWSGZ0fmTVIc3f2wFpAyv+xKbDqpJKvY8tg2cn
uIVOCpPyqqhX1FZxeJ8Bk94QwSXzsCtf1/Y6Fy/cNwS7tK8hNseUUIe0Ti8M
U1Je2IwBv9N8q3tdhzFtEQrEUavgroAWM5KoU40iRM46jUniVgGn64XXMvcO
UYlNFyxVE0Ydh1ZRpfPPlqQZUgGrbM5iZiMVnB72x/asP0X5bZ+uRFeedVFq
7TK+O8vxw223FZfjsKhLqMdfudwPuK6hbB/0H/3PBmjids9oGSI6X3/HhJVp
8qc/1mg/FOqYIupPtUGuX0e93IGBUXc1jOCp50yowMdbhNa00Fz+b9zBUPfY
O8BaG2Y2Ab02V0jteHul9SDuZ6XpO+8IpBxmNOWR0TRyNdzAGAjxyXtrGJ4X
9flu6vgZtTtsohd5aX8FDx27kqXpwUPMm0rDIh93jCcZuphamvYRTdZKuqbX
WG0OVXupRd8wyfPoZ/zM1cYqTnX5Zu+jHdP0WNCRAeeyj6S85RLmZtvopu/G
9XbKCWsOFM1kjPLk4R1Jsb2NWG8b1yniK/l+pEjGAAQ2mGU3rZzrQnJVoTIT
WhaBTKB0pgOh7NLgreOx0t8ka5f96Uo1og+iBp9WmBGVvCay7LmkdkpK6dGx
DYIcJRMmzKipynib45tujc9xvcl9pVZsnPiZfmJMVluyLKIr8B1Kaew4g8vo
tt0qBddERhSBMRC/Ir4mf7AmJg+K9N60hs5ubq8k/Q2ejR1bdbe0Y4Yp99jV
ukayUClS0yA7fUVzGX9joy24O7CfqWzfONtbRtSos3WzburgZYm4YxRuFV8g
X1zEE5GqLhpUOHshocURgb1d/47vKposISsyoqTSq/CtbpyymL8epxZr9xAp
5oXTtwnIoD/j4flpKcoC8Es7dOyHolMpUVoMeCdl44MmNsrgLfEw6/hgIZBZ
pXudlDe4ekkULVlIQ7ySF3vCeoD2IfQ+Mw7+UiJcHJ6LivafJns17BIMgtv3
VUeBVWicNtuL3ke7xAuViHfIy/Cf9IxAVZN/pxInwK7Hm3mf3vFshZquTmeq
UM6TysIPt+tOTJF7mz+fMXf06tW/1xHhsXTn8GDOBUEEubT41DqI441F6L5M
wB7mZbwP0WTe22PiVPDu/Hd/cn8IZqxmd4+a7n5e9StaHjUYm0M7U6Er9fBV
BEbXgrjvxbj4o+kxdDnUNyYlKjYtjubVNfQGdwL7c48sFOOzkj3arowhdEL3
UIwbfQkmvniLz7ZvbUvkMXJ3mMcvu/mfNarC0z4cb1i0EgZutUKNQALr1+Wr
ropVIiDT8/yClF5Tt8KgQEwnYnEXZsATeomxQub6+oHtVEBf16jGgiZ2jSdx
NzyNtR/pI+fylUNYWOhKpaQt6udyqIB1qfxJD3wXnPB/7Nk9sg1lhrrvHRj5
UZAJtblbp73U34RNeZVBXcUtJvU4bxe1DPoi9qfazZlaBSua2sfMfJEBgYdI
fLNHGCgT6e6BuZh9vZJ0VLayXRl3ipbwJbSxThdAaUJJr45qBLgKj8DxNlR5
qSMZqOR4fGNJpLx1eETJZ61vfnOYDhYlyf1htW9RJhTxf2euknnv8ksk/COi
06tQnQU6lCtntrP6PuiUIfwEFNjMs49xPOnqXpH1zddYRb93tIsEOOi4/ZFP
YeKcGhZJrpvEfKgm9h0ebAjl/g0/qMZLy/agDegoQ4vYmCLSI1QjAp+Bh+6l
Uz0hCGq9p4RvGXO255OgCaASmK6Jb+N6/dblkuOXL/CRzWoJFqsnHN9FL3BD
Xktyxw7xkOpEH98+A+nwBTHLU5NXWtOsGmyH6UzzVIgg8Sa+/3LXVDXDgLYi
vgd0OtNbPwdtWEwXmJs/i0bBIEK1UFY2Zi3RA4ir0mIEFNkcIJrYZrcVnZKG
bA4k2T0H1nzFpset9hYQ+71mT0WREGGFBJnH22RcLdSUIvFAttUGdK3iNExW
UAx5z/26+AzcyOV+hjptPdBFrKEyfqvGyyCoWjxg5Uqe3pp1vGlivQh7pi6c
JcVGofBFgJVp8i41vzl3F0NM2XsxxaI5B4F20xa5jDPItk50i2Qvv71E8yfk
GgbcTPRJmocdGhgdFKw4ZSwJUx1EGl/kWMjABU2L7hQSRVCIsunrVF1BH5vG
AkczPPaFB6Lq6DvB8ycJe/L0Cj7JrEb1GhE43fB//vxR20YtC8ZRUk4YcKYi
DX43hUrCIJY+c11SO86DZS6EpxSpICWdUvtk2yJpkE5njoDtWL+3RmSvShqu
Quc67UxJTHnwykxil0zrnO81lFtUIAmiefbQm6VlCzWBH0IKHoiKmrdItmsw
3rC3j7HpZf7PA2Q8y7xLcDOSgXN9B2NMmp47Y8m+eCWCpTANYkXFCmmfVv4q
tilCCFTAxlcMpGIzrNw13SeupC7hkNkE0a+uMMkD+pPyrwdAAOyNM9UfAgil
vPIhCfT0SRikJ0piCZ+EskJFyelHZ1Bw9zpbeJL9ks34m53qlIAfeBTpndo7
2UPwg3deyrXQ/zKxrTnMlgaEnfrnInbW+XZy6ihmYkVklCXcxwZ1dm03KUmf
W5WJfqS3ts39bvbDGnjFw0WhtUPLoBclMae28NVI8GFVDK6V/0JxTDAqc3oF
O25wiepYV/RVuetwuakoZf0vlI65oxxuLv0Aa6ITaPNW8W3eLL8O8U7uG5dv
4vSvwxqa7CW2at2CeKO1W2vUyAfPxx3cUZekz3sE7alolM5WApib51gI6eVa
urNUsUZFS1Zw/FF7UHkEJnrX3Rp+7PBdD/m9WgqwBeNNc3LV5vvjFBG88rt2
GQRfrqJKyST/cCz2dHwaMa+pju1KC8nTvhh3sDzT+mvTryNp2O8xU27YR16k
IqaupjqfGcvGCYNsIHG57tfOoul++aG/sFZAnQm6IfoyJ7v5mGmE0RedKtjv
I7kSEGGxo64milFsdWcljzKWvITLOlE33Wq/9njDMhnBVFZ8p4eO+byzHZVA
olZ7Ap8qHf/KxCpr2eicabN9bApIv+ei6Y1fZrD9TUbC6hJcLNJGI43TLwPG
3gOzo88o0NMnTThyOC+FwPn1+0+h1GM14kWYGrWqsKs2Tpfx3Z94NvlTEGpI
aRky84zYR+aQ+k/HlBUrqfAEQDWfoF93ZAn9gqrUgllx2lJvqPySn1wZHMSu
46QzWlp3C5d16XZgcytUo6uwKDtUDRtOLNOEFnHdlCiBrKL8Q4QzWpo+a1VA
wu5zzmViN6fAXbdGmWm0ihNx+vLD9O9Tz9vEc13Tcug5KKvkZSjIylAs4hEm
jU70NbyXR7uwVQvbRfTyKxv9i1f9AUfKRt7OR7QyohOMzf/mA7ymrQeteTw+
nnWjnWfbgUcrLu2iFpQS+8LIQbpEA2wgehdt9pNA1AfQgKfXl/jg9ooSlVCs
s7HuIsa9JX3F9u0c/tlajiAwiBrZFK+vyZgkO7uGnO/0XCLR3Ujmam0lQjuo
tEMktCOPJ7V5Ig0XVj1OX052tbT/uaf24poMienplsZcUBNjbOlrs/G3MYtl
Q+iwwjZQw10iEb+BoEB4pkuQiWFCZFDqi9bkzA004EHkoTpe3Yvut2hHXG2r
bUk31zqJp7O0e9bT5yC5mVRuCFV5JEjJEdFGwrCRZTxEm73SX/EYnua97dPd
PyOCBk4+ZcJdF016cufgaRe2PmTUbSB2UCrSKPU83nHGDimtjOt8IrKo1h4g
XHwl3RuTtRzLFECWiA0KD+2Zs2agcwCOxjIJD5VfKPI0g7dVwuXtkJAIRkGA
PxwsQu2cIFZqC6yQKNyc4OeXUmBsA3vdgE1YmyGwF2QwnSpsDZTRIptjQDhv
+2BoEWuU7LX++KWr2d8x3VLyTubBSue48ingZKMw1tbe9jTK5Yd1RXV74JKx
koxM4PcYfl+FIIiQRfF+7PBsWSjBbV+Yb9RBZwbJ6eReIDv1DhQhvYMFnZUA
7si4mIDFrCI2b3q3iNqkrgW2GmynE20Ia2f37oFOjyy8pJGVuCLPt4aV+OF5
umqMNlUbluuLizTYUwU/u6TfxbO+AB9cMcOciiCf4lubQ1pBULK2VfyvRGA+
o7yY+WIHyCXTRToWX6sAmuNw8XzT1Ty3ccaYtzhjEmQqVDD1MFVCVsAEdgI0
EFQAIinMjwjfBHrRuFA+iVdIT9nW9VtxYOuL6CFHIZlZ6q/222ulUXtkb9JP
ItTRmjiLKUHJOUzclmZPOGKm6pZon4dLHBvnRTEEsXqUYXopC4bbAJQZnuh3
Jyvc/bH9fCc+6noxssKeWmZ9AtQnVtxLay2DHGYkUvqMvc87g4SDcQkK011L
JOT25MuacSLyoYntjPM266vOA210vtq31Hzc4eQgdBXBEKuwezWwBBYlVwdd
8Hu1OqizL7JYMN/8eD0DzvfOXGWdlfZ1U0YK1eLL2JboAAIbS7HVfvKEXM6S
DukbpHrCeYSOC/JSWlcziSiXa9qJts2h/Mf4U0tjdIn//n4Npt6HpU7tO59K
GEz9NPo3mU1Ui7E65m4LMedpXYRtV25+Imdo+ftM+4CRxbcZpozxiptN4pBO
WO5y9KeoSL9xhpau1CdHTqJ7TI9K99g/scCZM8zHQj4S0Vktrm2jVCFOfZS2
HS4h+xkV7ZRY3ZxjTD7LcwtyV+zP+Gm9VO4mb/T5xE2Wpw6KxsGsm5RLwDnj
3KK86c0LKQo9kWqpZZT06UTGDXe9H5zAoNy0AcFDXniZbcAqZP2vCD/ku+A6
IKyx6ENkjLLTEsHhtC//OYlwEHJVrhl9RMKMv/Wf4FYVcD//fuaKrN/IOinZ
Bsf8BYLQoUyo2fXCIIUkovoIrRWQa/EugUsBUiqHjmxd7QhSfduinYmpFbrB
eELnNdWpIhpmZh1rgTaOYyn8rsEYJ0mx1kTtUjy2PFoxhF7yRmOVUT1jXlRm
6/NK/oWf5bcsymZbSZQ7+V58oBemltr6yLpT6+XgCoJLY6MJhCwU001FtXmq
4DIPoee9Vz5z8QktiEq0wP+Cfj+kg5boHelvq1NJks0xX4FgmCaC0mYZLGdq
i+lCGPoPRB6q9f8XCV+NhVLlHqSiLFkhcVFFTvmtJZ+Fni+AbRj/shWTLO0R
poTdUvVQon82/QPUN5Ghrr1hx/eNStinjRcUyW/U3cMgj/uOkWoFqLi3qLyb
4FoY9feQqwYzorua0YtCrHX5azyTwztXGYp4hj25Zrn8hW9Cknj7IRbnC4hw
mR912XVTMiQElZkz/lUJmB8No4ukh8AIOfHOytukdiE2rYAKCPiSRSVBu4Zm
sVQdnMAVFOxnWR6LjEw/Nr8Qs0fwE7UThN5BbP3JV89+p2TMW456p+zOofEG
wYyW0AmX34pJ7PdFwN7591sqghjsexEUK5bj29vS41V+jd8Doo1ETj24DtPn
f6IunIBg5Li3+sDprbPF2avpXuCQCfbtFVYthrUsJXN8ir+aCEskp/QZb1sU
1GVXZpA891rOKyD+h3gLzpfdjsBXGuMw+8fkLJr34jxf+XY0/48Fotz0o/gz
k/AkGBGa3RVuzvAlQ8YF0fwIURHfJ15Cgm8Nyp6p/Ji5TYWGIhxV99VfSEXe
X4y8IhXpni138Ht6cNjbLqQuBk5R8J8pEAAc+oVT6AX1xyFot/CV+Xrwap5i
FedLmzxajvVvaQfMgye82b2N89O+AgflFnj/9EZDbuFI5Bx5SD2BbV3ZjDCd
7EWWgtfZox+O/aGYc6QDvKFouIB8fCh/FU49S5BIAoWDaYdVTJDyI1cgWYJz
MI49tQ2kSro+0DU36dxPtIYDpQRznD8/42JrwmH7tl2m8Ia+VGuhtNfkkNI/
nH/slR7WZzFmsIShzre+rnFCpJ/JkSSJEMtzTy4aGLY445pveYiNNdmwgiy8
borzOFqdYwWoRS95fO2hcVsADat5AgjkaGmh8yLIUYruNFuqxrnvOa1VPALk
M9YBi7s+eI2f5XvBmmxYH0lTrcErrZAoUOPKV5+tktGKmS7KI20uua5JgiHo
BhXQfeBUaSb/UmzG6ryKiG1tunZqanRU0phpVgt6cN7+Rdli/HUeL9IFBg5/
T2RyFFL+HxYbh56c1aQlQHgcCEzkQZAityYZNitq9SCw+GA2HneC/HjeY6wY
oe6Yhx6miiQWKoKLxwUvRUy8PYnMQ+PoQrJGw0Nk7n5XMsokptPA6tkspkSm
gG2CfO6Y/ob2vH8cCsT1b+r8MVmqvypiLRAVS3nSwhZofTrwFPouWFdDdvHr
ic627tbaAwhOAcARP5JFJxTREaE415pK6gmBbd1A6SW6uEiKyrs+w6oXnpAY
cMfTLOIKVQyNuxiiWm+v4c8ZdL/o48moplxJ5hXwa8lTuYSZpshoGfqEdlHe
UMIjAMP85PwU6e/uapliZu3wjwPc/ekGGVdqVWBx5WNm8YB9t/cAU7yZrPpV
Tsz0iOSeGDCW1Pnzdq0ewbGYDNC7oh5F5wTGM8AG6lTk/QZ2gbuMRcxFogt5
Xl8Me3ZSJBNRcf90DcPqnynx8QR6xm27HfQ90OfWnSxDFleGfgN4nwXJWGhL
kR2pqdJxqPLZd8S25abra6k0W3jPD0Fv2XM+1AqbJpUh1lHyjc3TbADtn8Vt
PpIJVEamPTMX9Mt9EgJSuvMYPOF2+KaoTodpsmJWzxTYQX4rIQJlO4EAb72H
S/FSd4Qb1dlXy5pw8nWVQSZ33qMbl0BbDQkoBrABXtEYoyYjEMJAfuHlK7sC
IVsqR6mybf4sFuih0K/00B5xwnnvzjYvd8TD3ZzrOoAMRQ6cEoQG+aKnQcgC
aE84ChRM+FFCo36ZTC2seV6dTLlgW3n363/r4OWlkb0LcE+CaGigGeYBDKb+
aZFQYBbcX+KPjVc2+n2sW5apfmywjdxUPy1PPT8oJOVZEeEr+KVFGyHEkwbm
8naQzonXQoKK1m+WYbQs0TBj/wPKVBR5iYFtQJrAbTMGGXGfPiIJXhcVW3CI
q1M8Irfi+eXEprfnkB2BE0Ugs8QHl4yKlv2JAtQK+BedU6QpANA63xDobhku
o5yiOeP09YsouiduwwftTXwubYxkaayLjZH8149ks9twMCnsziq+I3UgEDts
92IaRYageQZOwGHdtgXPFguYEo54/GsceZWnSQdVq/3pMDGWExr7rYAs4paU
gcJ1YknGlE10W3qa1gk5+ZBr9yN9FLqZXbgnOrG16Ua4tYvd0uSxDEvYeP1N
xMpnDgnLux2igVJajVwEGuD3OeZhhHy0jWZ7b54d8a2OU3LcPvTCJoxMwkR3
TeqwIeryNEoJ2CMfqXb7EA9Yy7aAPzbI6rd6UbEdbRiS1jG7Yprfrffw4MHi
UG2t3XtJbJoUD5wSbcb9j5G8uTXO1Ixl9A8przh0tK2a1lf/DU1Jw/8s5Ftj
bfhk/SBwPQ4Xb/OC+is6I07/5JS1pi3OzIGVCqIDq+vMtaNo5iP3ogDUI/ol
XFmy/EozGLWKqSZDqzlPtg4bZ0jYhL1F04p3gQjxyENbGPScYNvnsd5ggvz+
WeDzMBgQtPOAewcrtyqo3LG3sqnDF3lZENeuacVxP2I15j59AtkR5fazKFLs
jHKlpNG56xkUErXlDnvG9Wp9Krcyqc9aNE6t7obDL68T3x4T7eZdIbiutR+d
doGXanWYLhz7eDH9JJTtjNeLLxjMjWu4pF5ks/hHih53JAtDnTPSlMNr6dfP
fsjKyY+D5uo9rjHpyCh/FP1/83g+B8uUZAXln5aKxbfJqqqwjan2Dy85YNNl
GEKhGh24sxCY27zR+pQBYOQNBbPZ4+LelBthT766qNHZ8Mnfjum0/q1UiVIS
nSjCBoUKa7SYjgi84K69gRvjChPYpL+vn2UsOt3CGifIQ+1ULtIqUrwGlUoO
bhO+9KucDAl9VP/1jZLMluqE38jxDLnAmePVWlsoBsZnYh5wAkwXBqJFiDi+
FG9227FufM5Z2MV8v8n7kX05YP5t5FeUIwMiyv6nDKDKRBH5dN/aMs4ESl0q
mcFmDydYUOerkBWTpdxKKney243QEgLq81PPlGHOYdDaxavqgLkGE6C2LRp6
mQU+wli5OreHI+CiEM5HqlhFrtUWeVU7ND7v2tsbKLiYkwlOZ1aTzxxxIsq5
U1E3EtLvA0abrcqsRXPFJjB4tMiqYRqqKPYLuFQB2iOerQ2CEHnFUZGKNx3t
LCno3PAdJY+f4Ld2P0Q9pWBHjGlqPQrear7lixrgOMLu61RblAttaiKmf3j7
XDTBp977SCursy76RFTVshjmG0DaMWNF+znbtLkHHxbRK94VSVyAbAjC/wtF
s4TMqCAV81JCMrU2UA0baHgtIV6yQlaJ/LWXk2LjzuOGpWua1U9AidoPfv2/
WI0S16uvPh0P+OfskbLDopsWh5mDUgHs1EYpBAZWoT74UTHfhbXAjhcTr9VC
Y09cbUFCSKum+kwtBtjFVYVgI4962ocNwILl/sTdhm2i8Oo3G4uP5no4kw/6
zuQrhuA+1GInzRmbxO+i2V03jQ1hJRsYKD+JHsWQg1UEekRVY4x+FgJ4lgyy
yB9uFsP55XP1RaUOnuCxJuAk+B579m99b3RFv3IIgky0m/vBsAB+LJBfGvTL
BNx/smrO41gjPJlVmrHtRm/jJDF9etwbtvxfEYdoOeEtjafi7IpsiD+Gn0a9
2akaarMhRKyfCJSlfwmZ6gYWjJphPlzPJ1uolHYBY3Lv5j45MImRMy2i0t6V
YPEuJIdIpWJ5e+SffaXMbzPMD4/nm3CDw4u9Otc77w/vDnKxAb/zdJXXRR89
sIjG8yt6KmAdGXZPx3Q6esqo8/9TDmDGOoNTBrBIxA2AJwdJkHoiwFZ6roSL
U6cFs90K1VVyQj5FirCrMAY1tCbOj0tsC20g8XAc9o46V/uM4o64ZN2nkzo/
anSbfFfQYBYI2d+FUGkLTcpAyB9wjjXg0NHThyBs9QuGKAgs7HvSTPEWHVgm
aXGK4l174/HLfs8qumqGLn3xzxyriV2HNfttlEfG7gdC8neWxhvEarmiESag
XCLv92Vxhx7J1ZbASO80TRsdYGPNcsE236ECapjjKVXdM3cBvh50eQhShzDV
CKC27uZIT+Didq8N/H7TBB+uTuiK7YRguMzL90YaHF46bp0PKYk1EytpURD1
Xr4EqFEegeRDq6hwJnKt+qa/B/zWeWd4rVqMK1f0qlGwZGaVhJidBLmG05Zo
Jejw+nB9HQNRJQkf8mHsmoH2PobwwygwkQdiUAWrvcgwCk26jyXYo3C3KCmn
76S6a2JfXDz2/YgdnFAAbKz4W9yUs4dyBOWofkJP2hQLOrXcE9w260SOnSYo
8KPlu9F3vVreHx6Kpn1hd/48oJR86eybpU6QsWeSUOlnlh5ZycMNTOHkePFt
QcsbqZkfdS9K2o5gneNGNF5ANAvgEAnbjPaDc/V6T5uFaHW+3ICKz46RTzlr
bPbL2RGfXlVp+wLdzTn79IUZKYbotNjSJNL/GC7iVtaBUg1ZL0FgFQS9sb4y
AjuzoxNoUOb4XRz1a/S34ShFkR+zSfspd1ybq1Ux5YoSYqU19028yFzPL7K4
VtqbQCesz9ghjpGkUf30/DDQFV0MhSU0weklxoymypVyuzc/AEKKdpZymOK8
z9PS5uulXbvp9DrF+yJxOfZb/tVsCjp/ew5oyXyT2X3zt7S3DmuhhNvML1Bf
H+ICVDjEkAF/P85C1s6mWZ0DQR4aOx4VcHe0UHo6XZQDKxuSmF01l3Gx2hZf
2Ve8bux6ChRcNqR0L/F2FXpqQK7I8ccnNjyFOTV+uAWEYOUyN40tItiZUjXU
H858N32Cw+uErYCWuA5CPeljRCxqkTxDWWGowtkrbM90uunUfxlDsrm9ZDl+
Q27DikxLoXMQ/w/chorH6P+DSLYN3LfMOhgI29nKZTHI2NvkCWbBpj7xMKiV
cpz04Cr9YbHWekWz0Tc7f2r14hYb1C9UQzEYKaPTRKVN/y8xVmM5Z9DnGIJP
oqc3BHjCLK8KrRQrqG63davqRn81hwk+S8enYcpMtcTQGdIQQhzEeIxHGu+t
rBnjKdpp7RLYxc6pofaOnGgIPW1LPUOCFXV8ERS7ENFrGyJmZVJxlcBkeSL0
E5PboZCDNXdh7GAALh+wj9Eos0MY37cj178KmTv5NfF0pt9ozR+MV8fCKLWC
oPYcuxqJMkQ6R1mLvQZrn+RC2D62+jcXvugT5bVVs+qFGP1JROwBc/O83pxg
OwWnr3aLbdssqxkjCKN9WQawp9SSPLkDqUvgLG0DZ4NiJjyXrhzuS3Q7JmoJ
pKY1S4YgJQkLK5K3wKtyPP0KvxARhPlfIG4AQqUkw+P2y1qY76o4eTdndhrS
wgW3doUfyL1vfn7S8SzO4ymcCknN4gri4nmyiqJghlLsEoTGdxVXH+KfMmP+
UD6VhDZfADbBUfb07LH5RRrHuQ3KpkS07TAw6/nk8BJ3km2XWqqQW3Zx+Chn
GGuMfpXu1Xl7ddmIWRxqnx0Cjplr9St/u+Oa+AFrUyw6G0l5vDtgD3O7XjbY
V1Isnq1fB21xBaraDKzDyzYvv2cx51BWVv6QUoMhJkgwaRv0n513sXWLZewu
7DvWD7DQ1vXUAQ2XgWXRUQkC+VcqYB5f8B9JYk2gLc2V6Hd4Lf84xMfr5S+r
w3fufG40eyYcFNZ1aDL8Pmj4sjF9BXp3NKh2L1aj5NtgfdXHbxNcX7iLzcpO
oWVMqCQ9Kmtcg1n8/pqod3lLccaGrmJTHiBp9HA096+awlbDXPZcy6ZG0/AB
Z/diPFQz48ZhOriCIAPgloeTZhaGnwXOuiTFGgM925nlDxvrJnjGSgD9cEK0
JPbVR4tJRnf8EB5ktiXOKoUL4Hj7wQbYzXj/mg9EEpTWatw+Muk5cJ985WXi
xNnSyhmh7jAzyhzOlu7S/j6V7zBvgEFhYyAhGQmxlNmYu0tqUGsnZUZfSA+O
XF21wl8JRO1jKXES5MjaSmA1+WTyKnTRuLhElm6l7a9DO5FlQIWnRIhOsjs0
GuexFk0RcmPiOu9HSncQY/HM79QeyAF4vV6tiEl9k8rIfqHeB1PLl90DEJ1o
CWDkUg8aXgdJ+4oaCqhjVLrqG1q+Z3BXLg2iddMYzV2HtlFyCGBRvV7JgWFp
OCzgGMPce5Hsf4J8SrpDINsRe69OSr41IGWfzQM/S/R8fveBPGgZkighlZYb
hPZCZiCLrLOErbpOLvGdZ4iRnBsyjs52R6eg5yjtXtDFz/posjgsXFa+dc/c
g7nWKC8kcU9W3lgoKeM0dXX74O9/vwZOESPkDTElkBYFuyvZOnnUthjQKFkd
K2BE5k/6h2i2vYZ6shCn99YW3+eHgNVxSrxlSsOkT8jCJKgfmLNauodcbeIJ
e0c8i8BOxDp7k6xXoOUfbWmVZqU5OJ/xQ9D6ihnbw0m+LlEMJpPwOqMGo5/x
jzpLIwuVYc+1IpEvPHEom9scTrFrk+I1uVjDhJL19YccnFIkxG7Ug9Jn7z9R
d/V9PNCcwpQXi5fafshAz4WuoIjZHJIvlB9XbhWP22mLIcpHTPDGJ9WUm7Qb
z75V5CyKY9PrPp1RPeESP9mU7K2r3OyByYG0ENmnGkivFVTjWqLNN5+HXycc
PovitnydUIqxf1jKVw+dqGO3wQ42WF1zWVvkdwmBUmBPitdsNE97KBPT1VUd
N5pwRbmYU9z/whYbLoA1E5g1SXOOlMiPQkWSq7etjJht6b5BnsVrAAlFEazC
aBxtMx/sPxMIIuLXsGqQXJm4SjwXzKUkzFYNyzUkKCYzk+RcbW0DEvlIL0Vx
lJjsM6T+iEIdDEN6Uql8MYDTD7doyrMuP3DccvzBaV7laS4uK13Q7H0IvYMN
OZXwZQExJR2t+OcQvLNBMqOQPgkJv9JP6eYMedi/pjbxjxfwPONXgnfkFtCI
uNTmRWOYSbcPjOl1M3Gfk/TYOVL/7ZXdIAijkWNfMifMWCS0+VhC31DEbCfb
QmDirqmXOkiiZ08U57BtFrEwHKuSxzOppDL+9AX16IXRgyn5GZWG+IRwjSIH
5atDCmvRw3mtbiuONEYarbD95DiQZAID5McDLEA4VScLtj9/q63kKtEE9r41
eTpErG/20RMq4CBND6BSB4kzRFxLZjs7s4Y7wGWZIsFiyY/wBLImFnk3dD7G
Qb6VvJVorv1T9MeTt0q4NtBfB14/9Vtms+/4V3d79bM/gj13sMAx7E2E+8oa
4E1JoV2ecodeyKjSW+KUmSlqeEMaGCrqfjS+bHWSTHS6BR5KG84Y4ozphz5m
ChJBm1zVHYl2JavV6QcaSnx5bq6u8vrMTfShbqJifGZEF2ToVsagme9vc8J9
RcIpw4AaAjKOSY2VjiguUhrfsIudqFHxj/12Th57uiUESQbAQBoXlHTLZo9H
BaeXXaeonBsCIioIEXRp7ddzUf91Yf94kfCIYRiDNao6VDFcCOe2rBsTRa1R
XF2Qi+WwG+ZD97feVmL17BHxfuWPdPDdOPHVlPmnxPwH8vPDCYMeM2lbRrHF
Qq3yxmMlMjZWf1Ox3xiBWGk4k02QOF5pFsBr688Wsxy+rpVqgtf7diZQ0J/A
Tlpocu6papJTsyWBdAM883xDwomd7hL0KbKqXFx1XM0P948R+ks4Rq8NWUcY
bubWlfbazA2iITd8SM0kr4Lf8KNLsoN/nHAO7iCHhmiDIvSdIcv45sLrbhBJ
4rYeo3mbKPXxRP3n7yY8Yzlze0XdC5x5rmJ8VpdyfYbd3gVvwt9enrh+bjtL
vOA7sFy2vnHqY/ZKoTgYnu1m4ZrVf8OeKmjkYuZuW9PvCwBWMwkNrDExkuSJ
FeBotl0oV1AR095x8dg3fRgg247wQIxuRHp61miYfFBfS/ZJUQ43MBYMR0UN
XnsRtsuUtSYulyePGMXt0dqTKbpmpGFzF+8HRQzTXXlCuhwvB3QdLec+1jho
MUy0r69sLd+SJqfZSRrAnTpmTkfatdIsNUh/ar/8oy+OHTeMSLtIUrhwvo6l
Qk0Vz7mMj+mNjCBfn2p5Uxqfk9vEcNeyBwCW+w9VagGFk+jh57COnM+5vRWM
X5VdNuQqtYkeT0C716SKRaX/tboWPRG83ybyjA/hkNKy4wL0zTx3/5Jh9zh7
kuEsu4mWOZ45QuhwGOrp4emOl3jZ+b2jg5rIV59TLvZeZxR4143EOz/aBySA
0u5T+RTaEl6RO7jgCEsrUW0DIHkPODlCJlp/x94UzlkfyTnkrl9UZtKnkfXj
lEVGJD5+66lB8HdrK17Gt7Z7iXLS/oOTTSYaGALECUUGftrCxCQu5FhMRqYF
m2A1K/WscqpB39W3QWPzOxEvf1iXPobo94ssuf4T9bnpoDaezWJg7jHpPx7q
hT7Rp39qIeZJ6oGr7DMT94+ZGESU204EIwRMb4FOWv2Ljz59Uz0jESVprbqX
dTa6OkKVpU+e/XafUeCj6IB1lLzwR7iSwQ8268SFCdzAMUXNH6AtVwO7+im4
5ew4K7C1kyqjG8U5M3Jm9q7PeHASnF4Y9A/xHzvWlzMgU8oiuMAkxb9UroD/
WT664IxTVCJ8sm6sHdgDPN/zA9CeZTTw29UXZmSQtJw6ffZuWl6dt1zgXmVo
0qraWv1VQPAccVzrCL0cC4j32ZGnmVlOxd/YYSvhAFZBUpITJNUdCrGYiH7l
XRkhutID9nXr2KkFHrACMn3tw792jEBdQcdBqpyGWZI5weOUDOsoVTqMEPR4
iHv+hLNft/bluksoFNmFNBs2tUAaEMTaVQe7tiwTtP2SUbYeIUqCtiNvdGsw
aFuUmtVTBa6mxP2EC3MvEHa6s/eiczUp+vYzwFC8W6/PqFaIjLbLw3hZIEpI
jmUU/8M9Mi037DF5THVVBM+BpY3C7ZnbQM3mz8jWwKKfmbvDK+NWFP3izj12
UCzSkviB1+yj9GqmNe9xoZgMvWO97XnQHDuIJowziIcIy85RBSvcN0WO3D/x
6h0nRA0VjD67W1UJDavS/6hqEAX8IVswYzufePQbTDe1vNAIUBsNPN24U7+K
+qwIr+BEYPcyjOm+XQBJRL4ZZFWYtwkcQAAq8WRrXUpOPxgxlpAYkcLzkgPl
MuCUnKrzK1ie0HOfZXqZQ0oLiLEn3da6eTMxqUHhQhQ7iYDKVdZZdvIk6ue7
Wbxzugv+vf1/DYuRWxFPDK+MsbmHZd3p1DPxAQLvH1YxqDq7499sPmV0qLki
HGHsZ5UWuD01TtE3H4BtdgTkVzRzQeGHUv2wOgzlxN6nmV0ifFyhdt1Od9Q6
LVTWWpa6/F7VoT9I1AHAmLB7rqS+tzZCUGQOODmSWVbdHnybJWB/LchWCh2e
UIVFw0I1riRPV2xl8XlH4dgbmpKS7J5Uzp1lY0I6+VEAIX4Cn/PLZY73IjuQ
VqTgaYinMG3qOd5CKqxg2CQbGLs0XFn8suKs4AwA6PVvSBA2f1fIS7xtRrce
ikldw8x9DJ06lDh6SNGJ+XlFzBqHgJSmzMRx4kg2XXG8SfmUsFNA1LOGwB/b
vgjbnXs5H6LXKTds0MLRW0wkWGTmvhCrNg/+/i8GiiPrLa+de2zNV6zuKp7k
IDERlVqr68qDOQ6XMSse+0+tLk5wSFVvw+1J+znCNCl6u33bJp66j+Xe367j
yjGawDJTENdCvZNLIR+bbdBaJL3xLz2aMjtLO4fgiOrkIYx/4gaRKWCGXQJA
zHrAfgZymUFEFHkgvrFVQvoym2tJMLfsTjsOKPacw1vw5zSECXxMomtMe2V+
0uze1OTT1C1hg1kcexQo+GnuCDjbg7rTWB3p6HD0cjESn5D/jOC8N7oeK+FV
QuPM98Y1YnPFYMQZAu2yZmTfmm7W6Lygz9XZ5lBaxG9OmJrpzpbaMFBKnRGp
yk/Gzg2mrNFJHMkADCxlGa7tkmsLt5peQMShpHeLXT9vEd/7po0q4XFsUMdo
FiAFVl/bJWmVzis03P7w8LH5aEuVLKnNvTVtkt3bUKB4FqVWJOHSnmmd9ov9
+MFycKdU+b0ex1wb4EOAAQ5F8RicgDshXJLFjZsrByzkrpazLI/vefycTobH
W8b1zFhU91oWQJ/xxu4oT9r/UE6G2MO29Zkr/nmPYIBDI4XgU0fOydggv/QO
5G4UP9n7ZKE6MpPa3eWohLtzuwrdBIFUhtz4u6pOAH1upXai0Ln9zu95hB1J
ssyGD+ZmVio48sP2LIEq6gLt3jRXac1RhEcPVm4AiIhPwblZAjCaRe5v1b+E
xyVmtAWPCjR4QcTaGzf/DV4/g9g7QaiIGl+52EmpmetnojxUAHWy9zRYDxSM
rF49jc8GXbwMNPcXRuOOTN7uU4NIA2qoHmiyZDWvht6TE2+yIKYIaYuPQvdM
ZYSpfKlJ4dFd9hj+0hD+jAlBbpPSARriT6rNjOhkv+Cj04r+WFiszVfKLtMF
7UiZAb79llFKSH9qfHpVeEgrp3qoJsSisLMpraDUVySwQ5X8/gg0gF0TdcYB
DSKBUJiS6B5GWcVr7Jqw7AVNNoAZ1f8Qm6REMccl9AREmo9+fUdGSErxxdax
z6p48nQpcWlx0Vy5CfTYvZ25FxfTg9gmTm9ocHY9aDKVI7Y/i/JLRSCE2xVJ
WtNJR5TMmP7q5axFlnDukwL0U00MZVSbAhxeavz7ieKMmxfXWx+lauxqb68b
wZpqr3x9sKX1LfcsI/LXQkN8hMHL/6cpdz/CSOUHQbtAsbpVF6EVBS+/Met/
jYaWic6RX8bQGqSmusBUcfC7t9dl/hk4voqKPnDxE8LyTsZKPB3TmVppzn3+
a9h7XCEMcTIefhzbtculQ/JT5AMyBj5hPZbqD0GU4gc3trt6RLtWukU7KmYB
xOeQORdMhN2nlokIPzrZ3SkrslH/D0XmtOtIvR2Di52l2iReSafPZoLgZv+R
JXvps7TF9NwD+/n6E3nNRJwFO3jU/Yzy6m9y/e7B1G2spLc8brmOh7uoUII5
lV07/esDPizNK5qy+eI9AAV9XZifFNtq0yseZVdOXzbw83oL9ubuxIHHl2XA
U2PzZWMQkMJqdAr1k9jNcMGWVxvFsIykbW1p6xW2nUci39u0UAYTYIRnkTqo
6/aaHhGAYcfViCtK0RNc97x5jad805XxHMzDNadMEvz9HzGdZfFeFfg4PXkQ
pWnUT6rOT7lZ+sViyrj0ZMIVHRZ3i3VjHum79ToAh47XaucRtiTwiBDYjO1o
661WwkMzlil/jWHHO0j/i6ezgbE24yhRG2FDdaLqKyxcYoW6vAjaSRvBX1uT
YcBTMwZU8G+VdVEyStzUrGl7zkvoXxfJAPfFUQic0zepjMbUWPz2OUtkBbwd
TjejXKzOumHoy1kb2gutMIHTGXk2S9PARsgvANzLdDrnhJ5Awl9re3UYmFuw
VEBDKM/Jfq18YWSSIhVwaRTW2/BTrcws0SNkqiOnStum0k15+u++mUeBmywN
oRkgVzZAk53RtHp6VOeEmsgPGd3JNlegZhxlWwJ3MHLutcArmXupmVqXW4+s
KuOT2ojTRq+yILFwzGgSSd0RS6eCRBRNyqRRpjeBGj/ecpvB0Yyol7Nayf1x
CplPohvQTMYYvGKpkY9GNQyvqQWabalD9011hOMcg2Sfa4R6VoKs+I6F+YyJ
T/ur/7nBi6qUz7t+qovkRXcN4+Jedh9nQLA113pQnH5DGkgN+1cfRtCAlbiG
aIUDJZt62eh8shfmscXcw7fOL+P9IkqvpYgdcEWESGg/Zmay3G5XgR7PXX9+
AnusK/M/fiF0/rQVuIiAGu5RffeMENq3QTPDwNLlF/ZbWUWwlUb4V2Pm12Uf
idGaUDFRzKXaqsoSv+JZbiUKgdfDKZzFuws5dVqBrswdlJNMHhmv0eoH8ZLL
dSIh+PrI9XoaVMtb5QZnAxGbFG9DbpdBtD3OpM495xQzsTE9qNF5AgszpZLt
dnnhd71pdvYdZOBLKhpxckXH4g1v6T6o/Ihg9MOiO7cYMjZ1WSNltUkWN+Uk
tul3tzVGPTbIM0HZC6DwRka7Ix/ZK1d0hVkNAVkHFbRaghfnZ88jl30MUWYA
kYe/S8WFaKl/9VQx7zbqt4Y8sZ0UYOyFScrgoSgxFCepL/H0RDgehluKwop+
Fbbcq3cHJp1pEg6C8AcT7ag7k8lSi/SAnHyRNYtH5jhNoJpU7dRvJc3tS+Uu
Ul56Il0gC9dvNFeFkRrWxUR8r13DqaTSKUP7Qd5UpSBIqWAf3cmqymZcnJos
z+Z7ATTNNCAQOlsnCurBORnEyZygAPF2Invhh3gMDv9gtbwwm+Azmrsqd91Y
Tk4Z0nmc5DrRW+g/NmcQR+LUMTi7+u+rBmKBtLO2BRk1dccTAV86mDdo0dox
neFAfgnmF3t5rQxeC3YXwepdoNuggmpNoq5QjSuHlHnV8qwRgFz5BRqeQ5fJ
SlieLMJw+Dd8AXaNOmcZwom/wzMmCHELZRt/q04uRwwotrk1erqQAqs7YYgs
VeWjZP/jJmv9bnl8sC73/mesT5MwAgNWFOVX6Jgo/ygvQMLfK/VqnP+LDJTC
Ep1rbIFZoa7tbFFpWQyfyTRb4Dq5bwZB+aXvtlWHrvLnVzPAmRYJOXPulZ59
yvKnc/UE/08IUeNsZ/qwoJ6+W4iOl73caIWKDUvswkSp+XuoCqARw/Qozny8
vwDcLGhvKvURTfvVsFnmneZwdIOuLhyA+w9sGjnVfTmusJbp4h8eVdtRrz5s
XXIfEcEIJdAIOD1n09RO3WyUebgcevBnkVwGc7lhCmQ2xtKcE2TBKcVBENAO
nG99Iqdv6wlhukyP9aPFgim+NfuD17QG5wRN0Upxu5M3dPrwoLbs+FhPPBcS
GozXCZJY+YVVurm6peYBF/7Szq2noyOZJn+2DnJ1fYhW7T2UQR6y5kmhk/h6
XhRF3WxCETKpp6GHW4usmhU319ZHrrO+NkGT5e/2lSP32eB5VbxI0nn9ZdZG
EnrU0Mr2rKRCCNYsf1zM1bpgSzjOgua2oLH9unLadEbt5riOnoci3Op3PPy0
NH68UlM3pyzUmPrMmK9nIR4wakVm1I+yHtfC9N3IwFk2ALjiE/R6ctDF4w6K
YtS6xzlVjXy3dmQDJvi8qXbp7AZBSCWYH7X7VhaNbOIA0xXgMmeg1Jkk3G90
lg3ATZUXXtFR4nIYNoblBtDVsMb5Nsbysgrhon0COZ16I2MlEpecWAUzMPKm
qOkFVaWTHGNl9OGew653zJi5WbmUwtu+ECZLZWarxs+48Gt1WwpgepZlKukT
RgqV7fT43JXYMowsDTUv9saeqKsU2wE2D9Gz5urWrZJOjNR3P7E2bk9Zv+l2
4BjEYAQXg9wFSD90igRt6yGWyUs+uybvtPnXdEBumMh7mI9y8YlGXiGdtUmS
UkGyV3MPXtrfIy4+d6PPXSdOxqEUImf5it4DWe8LTRJj3/7/h9dQzqlXyzo4
hMBrWeVtn2n3XWRFk1MUbds/kKbZTTZ+pPsq889qJb2qQy6r2i6rkG1Imb0w
MlInd0sHaT5OB219L6goE/16aIUnEQcGqu7ZxMItXTC5cm9I4RepmPusa6mU
mX4QrjkkTmzAFXAApDHCaJotd26bVCCzDZIwaS7lobYH45UCX31EEvDPoDn/
mQhwA10wrP48U7RqN5QGrIu+qtiBu80E78DwHor7+m5Ots9baj7qIBsDkPZb
PFo16YY3tj2SQZsp4UQ8WEcN0mA+ZLGUManOgv27lJ2aCjaANJAKRJU+v9Kk
xLrxuky40TfmDnYtb9m66sX2Ux8khtQo5VETW4rLO0n4mxnkiSz1R2YRZVqW
iEwXOIpQKImOAQLbirfkIwFzavfRkyjlTU3D904yeMKQXGc2+0aHedJNlKV7
n47q1dVU3IhJU94Lx/AusjBsuv4dsx4tR9Oj+5PG4k7zB3Cn3VQJ+4X86OcR
v5UtqaQE41JF3sSsBrFKuuAOPdn4aHBsZpV7T9u35Qg1yuCl+Mmhhftj6U6M
PcNVqn1OkJZEmTL/rBrm5cf/rOVsaX2AQHra7vkyg55/yfepTUNouhVFN1iQ
zjjMdXEeqqh0jprwG+qxLZlmrAhoSzD5DDLHA0OIbMMrbP3pzd9f1ZQDZnPy
BZN6excWwZKHnI2cQ/iHaiyECsQ4ath2rKAzwYovts3IYS3wBY6altdapX3d
zZ8vdCs7AyXBh7OWEGrlnm30v7BYYuhgoQ6pvkRcLvn0hIJfLF45zCMF5JKZ
1TvJoh/wr4gjrilHQOHGT4b5cxyG7ieLcaoj7XiCfSGzqGtznWZ7856lm9bk
MLl5kpkShy07djgdr/lnDuXckrWNxes/IKaPOaK9Hr9tUHB/u6YBUfnZygJ0
WeU+tBXnlWIww/54Bc11Q13qtpxOGN0CYKv8nIfB1+zuyJyN1wI9x5KUvHE7
rU8DnUdQ2EQEVLZladdefzbcnahi5/GZnM38lU2V2WB6ImWYyNFDYeesPCCI
D77kWO7ZSXX/+PRIwbBBomuf7v09NqrVah8a8RgtnQ11yXC5czjltEx/Rb2d
bBinKkT/lIasGp63VZubJL245wMco+f9vp5V/Ve93D3MaKBFfDCKsyO4hGbP
okrBqFZ1DUK5V5HqmLafIBODJ4H3qFjfA+NrvL31vnV2cGkIl/xdIRMeCh/0
x6RuPrti2Bnp+M4dB3nmfqY+5+XYSWyLbcw1Jl+TaErymxBueoZOCAyFByuu
VoZKqphQ6ChS6tsebbBicXfjMfSvg3YK6erxwVAxabnDI3A2sjciZqmtzyKK
7dhrvB17SkeRX5RCYzYFo6ef+ApYEmAWUsVuc6yNgc0D1Vj9m0uwjDkZ6Pn7
KzHo2SCVLsXv/0yU9xxpHvc/udXsACy+a/fFUui3LIiaYxwl8TwJv0rXj/tu
0odBbV8gbrrMUOc6Vz82gDtE0kYSxjWjMtsWsgaVh3PpdEntDmK/ZdbCa61U
c+zRhZk1Ew4FJyu/GlubJwjl8PlPbbQ1izor0bkfcNdvTzPyaJut734PaY8S
E7IcVsiznyc/IyQNtpyaxsgPUluZzKhtpGW2idE8lSUFRUH1n6cOLTaKl2jk
A2rxOYca5610XMiq+hgNUmwhsalfxHkGyz4NOrouwkEaRuxkEQhpOI7BEfkI
BZ6qfH/3qMpK95TldDdueSRvm6ikKn8KerMlyhf3kSsM7UhGo+GorRscRXAG
DzLQ6uhrHbKheZyJ2+o5oO40QTBBO0sgW72QGg8s7bk3SQOVNc+ovlPSIiD6
k0RAtvFzpNoTPs5LbFyr0ZzJJqxmj4J/nXvUumKm5oJvQK5HFdxeIi+KS8+8
9Tzd3hMjYGYJ5ffjcAUhxmuxQF82WXxuRHBGtQWqYIkH5Uf6u+ilnkSBXaro
XFOKw3cRPCZVTvKnhZ00Fdq9exfmsA23NIDJ8D7MkDxuUfFi3zV3mzVrCuxM
f2P34d6Pl70qgFBwNspa3bVLYlzXGBJwuHKvWSbkFLr6LJ+htCYo2VNQb0p6
bIwKKbY8//5oNFVySGMi90QVKUk2p+dGPcEnhww04KgLdfVEqr9+N/M24Vq5
IPzbMQBNqebOep6irzMStbfMfYLsSMYvCIhnuGFKbb2+Vs033KOsjeq0HYPf
m/bsdmpXCijSBCfBT8aZd8apZZwKbyDW6nvWHtLEJI66MM7i7vnovsvSV/Jw
7gt8uu1jpfHAcmZW0W92WejbkSVFSxyMCJTQu01HAULN48VlDJHigFD63InX
ipyxcYalwvzWTBQBVxcnI09WPtwr5WO+DPThv3RxGVzBfHy+pI3dQF8+jnYG
8K3I0G65X5S5vbWnIMhvH+FYqf6F+C/vDA727C4XQxRjyS96WbHNNzveqCPm
19H5ORb6wt0ct+2M/8C/DKfTxqMvbRqWMGMqDusxGlpfh2K+uRkxShV216fN
hDt1dBVHN8t3b2s+feVVSFq1HRE9STs8thExWBoHEb5Spu/cVkVBY5Z5nY/4
nt4CEnPTm/ecP8gVNUcClPVl8nQCL5tdomG5ERjdRGY/m2/q/ZD+4UTEg/qj
abI/OYP68tAbv8HV9GWELvgne4xjIHw8PJ0O+bMwgWDJRjAT9aGf5/XoT3/2
pTlpNxtsE5VPhLD1TDny0lZilOuNFnAXjoM+BxwSHly3XmwtuqxFwsgUwnSW
EwLmQY6lmZanX6vD8TEy6Gb569GdqpBl+Xc9B4cr0xG0zH6YJcFvW89NcvTM
euQel0GOqEJrtZDapft4JiNk8Fl0WTjUvogIM+gLwBGRoiMpnqTUF7/BdudC
PeTAg0Afie309S+ra4OU/HCkhwSzhAnYpgytCUQE2Ii9bXfJmmZ66Ro5lyCz
u+JWjNFB2Ck5Hb3a7r+WxJeRT7fA3adRk3YR4bSTtSszj9+SminkObr926B3
7Pz9vHgPzrro9hT48ULEa1TDQOnh70QW591QOK01OviUd1ibJnrEz75kVkZG
lEc9S45phHjTG5ENT9Srx/eJzo3ZUr7OjfuIeC+X3jkk5VMJ+UYOAhKAmdvE
kOsuaB5ieN+sTbf4hCHmOqNs3gNXZgbGMAStcsdv4OmJXFnXrCShJ4W5BiIR
cTWLDSPxF991FFmNuyCgDtEmBFv3X0f/rilYxiiZ4Ja0i7oyge2+F8MxZPxl
ahCUJj1P6S5w3KErhtRlyU/DsjeD5Wbu4frsOIvE6AL5ovJQ20F0LtaNH/ld
k1yDFVGLrN3E+l0ttBxbKB68LKr0QBK+LNlrgwMcwlTRoQQ0CGI5t9g1COF0
+f5oBJ3QjMvm6a3y3S8QJimJA7KJxXr2ss5fTPBi/KfOYv3eaghy0yqjX0tA
qxrwDLSw0FRSQHmSgt89nEfWClYzAhMauz5TvCJMZfiUnpudIxUZ1Ivb6rwH
pwkzYRlULpJr8Oo/irx7AF1+p0vcZ2LXN/7TMX7X4onNP/+FLWq2gMKiwcms
PavnEN8Ffw/dWU7O6CMvfOtty9PLS7JeOPc+FkE4ho6+m3Tn5EUyg6gtOLh2
r1z5WMAKJGjZLBM6Ym/qr6RukPs6LpcGNW7U5nYf5x8yZ91HBYrly9uxzdbB
UgG2ZvQFkASyoKTf9JO5t+LzEj9gEF5Gda9bWGqsjpNn1iuEUx3G18QAVEDe
FLc2dITprSWkYIkxe+TGgvuIuVoUcHKYwvB9fiqrmOsB9ldmBsiUNccAY/ru
TSC9Sg10hA9ZrNnSbU8KCNn2y7GkuQfk6mtflo7ghawqx42KvZAt77bxVu3Q
yXcNRJL0NINwhuv4SVlt+eFdylMLPHtkM+DqBWuQ+6VsekHP6NnKy2DRYwD0
dt7i8o8wwB9H/nR+IC89fX5VDZbzEzrfxbw2IQmZ/HofJ+5+1D3Uhfskig4S
ENJuqLPcGuq87eGDushGS8C0a4NZctZxT5WgOKsVaOneeEs1E9N7kwTAoo57
cs9jvq938DbtRwO5Ylf8Gi8XdX3bYPMa5kqi3hd/sVVqTNC6vX+uACDNvK7c
IA1T4/e8KMP1LRtyte8re11ypcNUfExZ3IN0gnCKDqEdDo4XKZukk1mggT/x
WnS2aFJmMGlTkLESTBWS9ebnlUyRsEwiDZ5QpKSGJ2TvaBrkixomAGhzq4bc
/6Hw8yzw3t7eOCMQC5UffCu3BqUrLdJXt6zV/pi4orYl1ZbluCLcdyM3XLwD
uBabIhLef0B9PvaC7IqmLypNrw24+nDf2UD0Onf4sk3mrghT5/tpJy4RnLPv
zzvYiYFv3ByZ6/B083JppMhGVgIB7HCdnnIb0IGJoV7Z3/pJ7Vl/ll4MrsN6
KhhrvylyaWp7dmqMyP+ibM1Wd1KYZrM3q7qcuCP3QAXAEnUeRGmbk1ZgmAZC
2JtGtTVhv4GLNg9Gr4M8FxEA+xDfIcwiVcVwcLkb1SDe9jadh4atAFCx7/Gn
bOnqzHbwcBEupk2BxScYcmoY0GDXxfpRevxfU5Xn+uT+RkEgAA23vPm7dmAY
r48MGnS4AK2J81q+kjCp302LZ7fhyCZtWvmjSEss7jUArKFKh3Z7u2V9d0Ub
57HR0Po0abCwMp1T1+Sm1YoP3ig0htMbDDQJZrDpG8DJYI6RSCc557lt1vj+
YiIvqzC84AwPn+FTc/txSRAgOv27gHy/ZpUQ5h+4o+PJIDiqbvao2mgQxXIe
lpI3QAK9Hnu3+eoVuqGF9eX08EfDysz1i+B0Vfj8Djf/IQW3dOxmnuOgrTle
aKvcUE8/fMza5pKu5qzal1x7T3yI07nq+swWcilK8VeAAr1qGADgZtB3hZdO
ZZtonIXNAdqmMGNXxcMtZ8nNV6DWbnD8FRGfNDsXWkXTJZgkBo1N3gSlCCOY
PYA6svnOIkwRsYwe6rLnn0UM7dNaYClZQbaHluZEYa0dQzzdOlnSrqzKwHo+
bNrSxFkpwIex9+Q0nxZbQNLqbI/mffV84RnncFXbbu8ZrTz6zO3ofIyofp+X
IXwteH9gmrEheuz240c8VHMyfxa2jnLq62+U50SFA9v7z863oH0eNogFW9w6
Nb08p6gIr0RhMkcG7dmUs4Naf2C9iT6s4JDbTRIBD6ry/Zy65YrsK0VaaSkk
5ITgRKzLGQ+hRLNSfamf954EMgTVNRUhJR2HGS1z+ZxugMUrnNf4c3DvTI7J
0sveDcEBmVADPC77Zinq9sXUfDZHxwl4Qd1i8mrMBhYos5R9flccBdrIVuFP
DtMuOpsWk0RTr4hMEP+n91Nxv/uMu7pJMSqbEGJeJGAbzP0IkPGz1LTTGz00
EFZk7zCb9y/84gHQHkqwAdTA1+rUcyzKUx2QeHjE9JgdsipycwggbtM9kave
p7Ds+bTqDSnTjbPbew1nkR9e0nBdBUAb5R9gKbG6wsuQEskvAGqeBOjs50EB
+OIvW1I77jm+G+TJczkuOY5rvD9Yz8DR4QatnsoZbP/UC2zagujE37NVAu3l
yiaJc/wy76z9APG/PPv761V7dMddEQRVxO47nKn003D5c0GS/y3WeXiaQlSQ
b+exBN+1nah3Ry5Iu+kZSyEO09J4JSuAYpuXOhwyF+WpNXduFh99E2zNsYw3
0QCwuDhZdwNo/uXYSs6fPQJMeZQs7fOHONXcwyxjqAjG8M5D/zhV5OTVUaV9
Rj7ERSo9PkdHamK1ngsP1XKzR7YvmezbeeCcJX5kQTbxqpzLrfb5o7Wmw6ZD
TL4P76+xit/qRWdd48ctkHBGLVvPfG9JE6gsDjV3ZWp/onYBkgfT0yGxmfPn
u3Wct6rdY7+fyyHDaLNkWjp1eb71BFJfdc0qM7RvZR7+MYKS5pDTXPFTR41+
5ih95W9UvK5Hg70VbjO4SltYK4EKHX/PLgrMDmA7zk1Gl6o66xSm+fEMiF4L
ymGhRtVHNpGSB/f2b8aBDeGa1N3T2MVZXT+9RcjkG6tdbzH+DzxEWQabVjO6
uhzcqWCeZisi14uky9sA4Uk7aSmFAaTxhwZShpNiIeXIhS3cRxA9Hl7z1A/Y
yNkoIRj82bPcD9W+1+ACaQ0oE6kRfIem5Q7n4LhVXR3u3xEH2/o/0Jdp2efR
ABs5iOPGcZSyG8pB4lXJSWUXqH4M+TgMNMoEv7Bg3cG2b+F8Cp8UsodmtP7w
+igrl7RFU/N2/MmpwLeAH/x4mOYiBu9SHfsP6UuC5GCKqn1pY4GX1om4oZsy
SpYXkzYwQSL4nD+uqU+vJwO0GjLX4CiEHKSgF4nk1iTJ5MA/b6BbCsrQFcmk
dFcuHmeG6lu+9KGb1T4leWfVxJ0k/UZCbCTA3L+w9ndeuDjqqHj8XnVxNUtS
8xPExEcYvzPXdjyfJhLNuGV0sL70BF623q+LhZIgA0JUbsosItjeGCSAznQw
hJ8CVFaIy5q7xEzDcUivm7Kht0jE7ycZFI9h0IO3ZceGaV6D9o+C67RVTN58
dM4nHszrg8njjZim0svKS9VUWX5/wM18qoOkTpitsePD6KxzHPo5T21xXm13
ekX+DFehnW31HwaE380sMj7X3gfm+ZP9ONw6X4cRoSvXHRwdtwb/8FsGd46X
U6xoDdnwtmCFBvC+m5e94MqHvK9NVz08UifBz+VjCDObsD+lBfiP7rmY8S2e
avwjy2qop3Lf3liqyZilFukNLW68lXnFa1hXFqXdOm2h80zPWAyIgLSMwaat
egpk8a+SnkFSZhq7MBSBX5fX8etUdMXhdIlqrt07sAuT2UKCDjyd1I5DJGfC
5yvYIKLlakd97sl6XiNwZSlyfwaijk/Rh9sSMWYXDZIsgKVWuAyoXeRu29WO
FqFxIbBCktYbGq4ShHoYfqNBHor6kthMKqb9BqGQ/kTZ599c3eL/cze31Ln0
OU4pAJOSNK2Utu7EFOiHXRnzOSKstAZx6BEp5slmwiczj8jFbeffN8kcm/74
0u6Bfe/kEhq6qd93oip3rq9v5BgkumqZfUfHbGYOXAYiW/K8NNdFJX9SrHcD
W8GPkL11aSPv+KS+WkPPwx/uBUw+3VBVOY4WQE7SFw9gT1QqH9kQpbpaLbel
nPjPnpSLa2vm/o96QKfaISjdr/0q75WsK8hRo6zU3NNztNYnFJJ1CO3VzGQc
3hpUANoYjqIeZru4LKayE3gKNKUJo6PFmI1ApHI2ufKjoKb9VuGyhFEsAnOa
WpvOk5SIwQDJAHCqvqZTZggUeVGLNxf7xtMnavmOaj3bGLwXZAq5fnvjcASV
xBcPQxXCPV3Schj1S5HxKRhYRCzsyQ1POXqcz3uUAzRo1vv2iysZZdc8GS6x
zz8TbeFgLxOpWl9A2xJqj3D3hHp1Mx6tOj6D8sgtIwsipuL6Jh3qwBNlqfag
8xhDLleoQ869MffwnMFlI2Or8Uyf7ljQ+b3z7jIppCLjfQMee3YOorTsDy28
MclUYFryeIBRevpLkMoIElmD3aECK6zMNkxJrHBWt+PS+icZmkd88gRqz2ji
A/EI2v7egSLGYjx9aV6c10CXInEvpwT7zNTnQ5q4G4z8/aqVeOpFCy+tana5
ac/yTbsTdVYnCrXnj1Gj1+qZoAYFsH/51np5dB0P0VShDM+zgIYdyzbaNUuE
hPPukQZWk6/OLHNWK0ZgzKfddGsk/uknbh3anJWJivymSSXc/hoERUskG2lw
kcwn6H+3snSf1fXUQHAjmrowvFN4SN4pd+a/PX6Ual+0BEMC12EwP3mUKRuK
nZBYA7vDpYEkOCCl3Z+K6F6Ws3Poa7JXByE7F4kPuDZWS5M0X0BUi9vM5rng
f+eYsXJW+aQzoYLcDWNA9GFDdz/ifFhJ9wBFba76N/YeAnoK4hqKNwMuCpfc
R0iUScAFnwg6O+Vp8CnM4UEcDZjO6u8maCsstO/l4vfHSO7oOCoNv7ifQAhI
d3UPkTPtCwa9c4oeO6m74qYV0+qnF9EK0Wg5BHnCeSMWd63KX/7YOsPf36Gl
2nju0nGbmYwJf2sNyuYhseJdfG/G8XEDeatH0vEfkqOQkf4QdOq3ZOmQNQh4
cGFTBwEsZm5jMEwmu5AHTEm16o8S9KbpWuLbYYih5H1OzmVW619jBVBdWxx2
f+ijpRDov7z2H4VpanN2RIJUAZHILJLnK8gHJ01qiG6VSfGtjB0YnBV9YZaW
ZaV8ijUk

`pragma protect end_protected
