// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
MoqZRUwM4CvG12jsFET0JNB2JfL1ShEsFpFl5x/sn2mUJNqBo5ZqrJtezwuMINzV
zvwmbCgj/JlV7fxmeg+jS2ASiVBvnC72tN11r2LXcuEvBBAZshpapk0XmhWQ1voA
k3zLkUJa6jKRcC4aCcs5fIJHMtfCsSIB/Z82FbiIr8A=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
Ao6xzglC/zdbsMbhb7dhwfYHD56liHwIleS+uBezolPkl0ksxcaR9BUXIODSKT0E
NmNPZSTE+iktDyeP99WQVck7EslVDP2825NX0sXgD9EfbTViS9CYa5bmbSX/ZAzZ
GOVK7VQlexv3FhBW3mfW8CSVgInTwgfrP017HOgsHEdZuZjq4CLuypEn5ubUqk7t
zZJMIRw/WLIA2GqjrDtUQw0QlCbYVLxIvlXTXoUqtq05T4c2/8nLEbXSRob/cJhY
MAuiTgDUxdbEdP2qYlzKzFBnM7Uh/sV3Ki6uKidd9fajPmf54sbUSJEPFz6DPSnX
YNVxCe8fvRcvuvgTJQiXPQm73/v7Ttc59QcOUA3YEstGwAk+w5kQSo9WCvR1ksbR
9v6p6UcCwCWNXje5h89CjiVemhXXV4qfXVGVR9IsZq/aJSBE59o+qJ99Vd2e0y0c
w1OPYulqZoC/ce+v6lu/BL44+ws7ofsz4nm8JmDm3g7JrQ5x3EswDIy/BmibSsma
DQzudMPCcRTskN+otXiCoQxSS5vpqRvLAaQBv97o7+cTkzTy+4HaytshqcGcnlNR
Eqx+647eTUVN5y6fk8bKk41K+shRlOMFVb5Ch4SztsE1SuzVaoPYieNMcEZhpNHg
DJGgmlVy/lU6l/eWYD1VZ0lG1EQcc76YHrpNnO2+xvYw9lzE6kG9TCFSi7Kn97hk
xKl/h/5zRClSqJzOitpcNpENDU9nzDuQmurTmCgkqFGg8ytFX9cDWycswt9CI/H2
QG6wdJt8raFBSSeHQTE9vhqYz196plbeHyTEB7ZC8HJFiw1dZ6NlP1BWfmVE9qrS
B9mTINfjvdffkYjbTcGlsUFY5r+HxM9400GcvHdep/PQOZKU0pl1udTEceC26phy
XVgIbmL/M+KSqeWxCTESQ7rWTOxNZ74jJ0+nlCL/GcN2ICZmafcni1bWvgt/Y/Xy
Bhav/cQVW8UIAMEifGSxpIhAwY8y+tHxQy9BV9XG65jNYOqTURVqJYLGc1MCdvg/
djHDEVfPzautxv29PLOOUbpmslFK07xaKNss2STuEJHT9vARkke10awVztZcBIui
LywC4NiIl02ogCkV6eD86qqvmhaQaOrWJ4F6c+uQ/c5n2MVBU7UXC6pU62jW5gQS
qDmXGRsM10SmZ/lArevbbCUaI8KF+6f7GOrMVnW/Dv4XcxDBnECfnMwCPWUfTuf4
Z+kbv+TVwRYTc/grF+bH/1ZMdb52OrfFBBxGDb60AtKlXE+S0MB2aCh8Rgvu0Mjj
h1uhOodh8D+iFKX/ridFrweXQaxpwZAceeDbfYHb6GM1D7FH/jTn1tMfX4668XfR
MY0pcMpUD2dnRCdk04zzcDz04YWJwcdUg5K+2QzjRDWwwDxkQYHXXa7xQ9J4Zspu
kmKM2YBlI2cH9Mo7MaGvfRKn1r29DE+mUG/biledCHDRM1uyCtp+43mH7m+EC+cD
5a4ACkciAVXhZUkjkhkruECHFEsPYhVCse4PlHGuFGG8N2WH5wFFNSCcxW6h+Osa
5GAZr5uVjaVvGPtntZUlFtyrUomppmQ9FQYI693ui/a+mYYFthzoh/qwcFCgsZz1
40WfO+V8dcshTBViyKQzFnfvkrPwk8RPE+F4ap2R2NfPY81hDtdP6ksePDNL62M3
De1z1J0KtyXKR16lo39DjpZwg4GrvtxetfCtxXMJ9OnLgwLNq3b+5fUiSiZSmyD4
wL7J7NIgCLCPxqU3DSEL7vcFAlA6fk/cQT9REqmeLqrHylGt2Nzo8int19GkjQlq
4KRm/SohuB6Hnb469upYtyESamFOkpbguZf5MR98OwNGiOxA9DTzPQTcw9FldyLT
8afONapYVPOIXm6YxHaVNJp6kahzEOJDg+AxGwzzQbCRsrot4FF89kakW229oUGS
evZmhAOdFDqo4HOiqoL0rt5WDHTmKTXOuwEm41q1tliGPjFqusMpyM08e3BYNweg
dkh0bLYCERx/Xxu/eWC9WxEzLkd0qibvzeN7NALOdSkOK+hZGtwgtc/yHdvSb8dH
mEFImw9A82/+i2Ft5/1AfR1ROTsg5mO+rUiD9w0lMb0GZ0G3hoLdcEzzVCP23pGR
STvAMcIEgDXMGan94fY49fF0IeZ0FxAEcdnD8xYrxSjVH55lWrewQs8hl61iGw1S
VRM5D/lGlXFYvIV7kkfELIn7z2H2l35CkyEt4EiLqdL/9kDmAsdtdwIFLRYo9jdt
1yQSfphFqacTFQtdKNA60DekeYe+Nz1KBZFd2EhU/WVoBgPojsGbJ/MshgiuiSZL
u/yGmGCAin8XekBpDsM4VYGEQ/YI9n3ntTJVMKU3ILibcGmuk0jaOoXahMKyWU2e
wzJuHuKw4PY2QAREgUc/LMFUdcRHMQinHw1RZzsxYgzWBQsA1X2/tfQvehzQLm2e
6wgzhySucmbLCG3y/BghRfj8cR6puiBlXqh2uGFdVSmr/DB3dGNyUSexrr9o3Qxq
vDF6wMa+b+Qw39L2TjNoDhT0HSZeuVxpG4JBSbOptKgdJqTy/ShwTk4PWp+b1+v3
K9+765XmK3oP/JKhLelSHLSi4a54kiQGOZ7JcI7J7ifEHmsaOSmmsUDgL7+yJa6h
MQ6SWWK1FLpQUdsk70JMZu7SRsIJ2TGT416xhLPMDnbI9ASz2HomM3uNi0DDxO2w
PPZHk+5iCg8FQ1JBc27/X5RUdnpoIovpIsCoJSNgmPUoRDtNAQPVt+a60YTEoxXA
jXtpiRG18mZ+jaP5yzLXfCDxdpU0NdN967qZ4sgR9D6r3ll6IkLQ1kI1PQTKXnfv
pV9gfu+xhL/fAdEB4EohMg7zd7b5pri6chOlbYABbUzX0qmJbO3rgpM5e6FJ/UZe
1dvVitN7phZbRSB5CZieQu/kf73p9CphN5I+JMhhZWxetG3+Sun4JpZY0dY7lqhu
6fnejpMGwT7/UUOF1qjRhHLNuMO+UC0GFOq2phdEMAwaSzAfvI4wrJMHYO8oGT93
Kzs1LbreacqotTD/yRvrMV5syx7f6oPJ5QdyJgl2s//Fmep3knFdtLssUgvclgzt
TjXXc7XcpQFun2BLIZBmwNVAccUw6hxtcy0vchHbtPaqzUGMihwyNyjthXM5rxIq
4d/cffOn6JzEZMvMya0D3gl6oB2x4zVDm0yZJh/bSQ6w8SqoKv3zj+uSkda2V54t
FrZ4w9f6vWaK/plTh3PVHtGO+sKEzM8AFEAfCxMyL4jnWu6NHDmZ6ryJUWWQQov6
IwFxkWZI2Hmocqim6pbENJFhwiz9VkuddmiFlzeUuHZdIEbBUBkWqMPK43+qA68w
C0yIeLTQgEJ6fPJyXtpIKyhWrizKUWi2MaN+6KhZXJcXW1FRa316+7DLUG9Z3VeM
6Sz3j2dY2k3MLClf9leAntBMcrxvYNCKVL3+9Ok4d0eFqwSMeBTdh0ymc8MXNn8S
00P46F+9HvAzGUThifW4c5UVQdSOpIbTEMtcXSE4+t6EhXpVVWbFNSfqeZX+LLyy
dEK2JaPMOoXre866854ghe6Mpzj4UvyQ477DWiSir7LR/0Ru0w5GdJ0gI8HQholt
1nDl7L+9ScvJyr1QnguQGrct9RF8+IANv97LVWDnp+Ev1r3Irdwx0ZxPZjU8H9UV
VQc53du06YTOa4dDc+fe2FePg44c9dJsu/jnXw3cBjcmxiHFy3SB5qmOkgzkbcjC
WgbSE1mBMQI4CZnKjCsn1AZKHwtiiSBIv85vH0famt/LMGg6y+WfZ8Mw8CUdAwrU
sO+Lz+ZCwZdfhBx9RINxLTg7m5JGRythKOo+E+vMkE1qBs7pCq1XlJuqRpCPDLI/
7Q1ZWgTL4/BqLRiVLOHoYRpIPpT37nRyk9e262jRknW17zTmkF9EJoNeKKzEEWuY
2VjCulswr9ZX3so6ffVWBk4RcBcFJguqZMMzneSWh9udnm8K4fdqzdwQak0C6DeB
DSGRfqBG5Rk4J88z7Fw6djbwvb3xakSPDb9aJr9RYkavcqW5aA0Kar4rM+YUPCr3
Zq2m5vD5f38xSnHok6IE6Cveiu+MjKirE09HwYF6qKgvvQqoHnIsFU9qtO0pcjrt
a9nIudJhpBiFYE5MFzfU/ZtsTR/KJ/McTyVtYN8tHFBkiTp04BPP8al+emOAoydb
POingRqu67qki0HBEhJTyLUrDyjc+9IUxwI0s61bossr6a/Wb4CRNYsgLoAhE0Is
AC1MNkhcVP2Lx/SD/TR7j9FJG7bMus+efOUNRQnT7ReHFKlkGoSMqS6JrhU+j/YU
S6QP8EmqFC6mb+zGnGoLmlGZfov0abBrL4E2Wb2F/IQiSC3DgoPLgql3J0ljDTsR
g66tycS39s4kxH1CafKWlzPQ5e/YF6IJlfozcteKSFrUtu/3s0BSsnaGx+0DTHVQ
URdIwj+ZMs07WePXyfzFnvnuRAB2j6cCzqTgfb6POM94PBTuPq0auh4fohQqcpFt
sqYLqwGi1nsU+E/23jwIwbSJoPkk6aiuCJhXhR5W/9haeDTw1qeHSjDawWIhhkN1
IAdXv2FH9Yrk8hJydMRiK51rjEPI8hav/dnyYUBs0RQ45S4HBTDQ8FxJWPzBplkU
4+8Y92nQE4Ztw+YIyQiC4xWFP1V9vsFbcEJEtHGlmY+Fdk0KUiOtsy7fc8fQ5VsF
NYSMwzAI86jmpK2VXDlF5UIwXyWvBm9WYz3icYhfG50PJKDZnfI+Scr/LJAfFFfS
ed7/dVgC4/PnHst+HioIF3rai4FRhy6V6I6Tr8s6D511wWmcaSefPy/DRVBj9U/O
wnM24KHwkUbGhI3HSGFMo8Ne2cAbi2cF2pMnR6sd94U+p7yNA9Hv27a4FIQe+pdv
u1PdnUj/zRDflfoSOMTpBO21InxcnwbP3hnZO59vMQ0AXud21Ccru6fxlYDS/8+m
EdjLiLSM22BtR7t3mNPYWdcWVGXG0i+VBrZmr52zmyFOjCBOQiTgVWpL7Os4Wr1D
W5FWuVsjxTJuqHq5lpPHij9X1jnnSl9rx0EMhAuuc7SV1KyaOyaJfow4zcSIgmGm
7McUG24kxi3G0v4oNV4tC3uaojimYkN7FHXkO0E0/QKReHxQIHxPGKgORmhPSuLz
nB2YKiDaFwq/L3rboZN7WKfaurmseZtA6RJign5MQHbXs1cw3eLNxtlrPWRfDIHh
ZB9z7knoLJmXU98byVddgWrs+NP1OYDRdsK9wtIJv/g4czDOX5FZazifkfsTmBQ4
2kbGwMBUMhBTH0zvrhc7j+uxBM1SvEyVupd2BLoltcMeP6kqcrNmJlSTEnkUVhIQ
Q7OeTfY2r1/6/VkCWCD8xKhFErqbQybe4IbUrvnVyjGdhpSEH/jW/S2P61eL637u
jerQ3nL3ZonwYFVzCgvAFSMB6himA9sHEJp4j4bY2LasBUGDBaPrTJko3O52YFq/
hHV/UXh583/+XPhJiFTL8Ipbdc8HE8xXcXuB0rj4RT4LyzP+VRRrPxHTLnDKFAa+
ivGo6UgXyxHYBWZx1VqWeJMuGHUXcT69SfdpiXKtxlVuoWIa4RoWDY667RUFSumF
fl7lWdD/Ema+iQVIqsAjbJejgQYc+9Vn00hu8cpEP6x7qkTR7w7hNXUB1h9YM+qN
9dytSUWBYpab9HBTpwr6X5mnsqI/BxGXs57zfZ6SiO0ICZ8z/tD6V3L+7Uej9muq
vpkJm5zqDMBexeLYT6GBXoWsi4k6NyDYGLW+b9koVboqFtPTjaf6eWyN8OKBtir2
WeGdkchLNqWnc1S8ztfl+MCu3wOoFawYCjEHfSMM6gNWz08zj8+mRHY1DzOApnf6
rFKrP6pnR3+pXVtzuzo40JJj+y0D43CCavlpvFLXNf2si/9o6RdSZ9MmKWMx+H7N
FpslZW1rpPQc3JYhTJ55MZWNgbH30j8o07km6cJ09lVxcGtnNAsf3IDovQV5WaBC
c/EaTX0bsujmb0WbKS0iBGcDpjhwPM7hf/gKy5TRli1nP8iouDYBfJxkeWhkU1Dr
6BAxcl9Bujnyx5sWEpN3nk3KknzcYVtMWO8UV0IJSJ0QT/i+JB34Aqx1ISi1Xvfl
OQlANHlb/oVLUBjppaqfxuK8ZbjOyA+qOddx0Qu2ESH7X10rsHb6tVF0wUQTB/7Q
GDTUfTFPbVKpLTTSItbVbJnWxQCnAaAv9ePhWmwgqiUZQ60WjrxIwjQLsmbcVVuH
iHexUWfqnOQg3bn+dXAmHt4al4WK0K3zS8oH36FwPj1j0UNQU82ILtWR/OfLUzSr
Zt/D3B367OcpVwHg3Lf5S+VCji+uyofuu5vwuXv+//RUSa2zWtFigJSOFqsZf69N
z3YXWOqigrhxJd3Tw5KBYx/SVnte4Jru4Lt6Im2H8Xw1q4nwmSNoXz2zyf7WUPPj
zhCI5fE2A2gOCkKiZmnJ8h+2QOxJOB2GpBh59BY5eM0VwVVn/wXrbY89IpaBMOmr
PySP87YpqCc47Rtoh7M1GN/jhjHrGLN0Dec17spyjBarNvIZUor6aZ85H88J5/nR
ozfx7f+anwuiWsgJ7wNS6NSWEE5VEaZUqAL7b4UTS1yng0FqK81MPchINz5+HUCC
idh3LxW7aJWg/+No89J78NQZvlCawhQKGiVJfHznvgEWSw54BpyY7XESPH7xziZB
E0XW/1dvuYDkQ+Q1QGuO5O2JQa6KYnjQfAhdNgEfKNlE3E6GZnSVAkPAb5Jcflk9
EiGd8PZ/xfpEO+tRW/yZG2/Wgppgpxm1FPybzi7D6moOaNhjbX9eE+ISSnuBnJQX
aThgHkgyYbBsA0JpHUUDNPiT68pwdZWh9Na3k4N2Zy4Uphn17H0GW1jFW1RBYQU9
cHkaY++wYRsLRMHvwXVUS9sHCarBwSLTL4jlbn/ei0/JtVgJkiaytxldPen/WgYV
WudnQ+KFI13ugblhQlPak7DdtHWhPXJRzOQXtaN3oIDQCHBWG8Vg3TcTV9ENJuDv
dMfmT8HNgPT3T6w5Y5gLjBrBN8QyOJA0DQelUMIHJBkgw6nu8MwhkoM24BsgcEyO
+Pc+UyThQ78LJ2miczad8PVjiZ10lyNrvcz8HxHd4TFfDN+3kb9ty87a9Ce0q/Nk
NPiRQcTrjKsQueSJcggMzdcNLFHrcSTrsGd4Rjc14c7ER57S5gB5VN4pa6nCCZ46
pV+z/wpJRciWYzbonc5btnUyU94YKZ/scldhg/VgpsWc5xKuYBQ/FmlAKNN0vSP8
Uwn53Ay+GFG775HVFshOm88qENDtfmEuM3k/psiHxeXzCkb/oQH3VzVHUH4qwyey
YBj0fV5Rb1y11OwzbZf0nKc4KnNm+bPZk1kL5bWkPf7fMUfTRcJOJ5JkkbUCVPD2
KwmWWBC2AXr0zdJJjzwTwiawpd3P50U6Ox2eSFBAvtxDQM9KI2h6ComWJoWOMhD+
weVdPO5AWEflNgnvv0l1/A8zYtLSkqVg6OaeMk8arek0Ri8o2DVlzQfzwIc9GTQJ
W53uaFyTAgfdM08TY1yRqZDSYPR6TFNeGYE3I+raTAsYCcKFiOstu1THMimMcyQS
nXzW8rQMRZBxnQIstD4H64q9hwY/aDbTT+475DIKxHx5A7w0913YkiWpIlQtkTlg
7uvXawO25W1F5E/ete7ujcF373d7pHKoFdGo+Y/Nv19Cpf5iSUJrH8cuwXBntiCc
KL/iaW4O0026V2M90xZmgauT75HSZYml3QzYE06RzUVFYw+rntKfbgqlXmi0eJvR
j7YBhOOgh6FOXUmUInfmbYT361rqhnJ/jjSEc3o4cyEA3vIqixyt1cTvEN2PSABF
dDVbmu6iZaCYvjSD209L1BkMVwLh4LBtWyr+XI1BVFZ0f6FN3jI1XKoARptznz2q
AUPErE6rYPwJ5YxXXcBOGKVBUtp/iCS7bm23DPg4AC4o2w+GVW+pRKa2B3FGFMaL
PJrbcnJdU0JxNcRET39F9n7sf7wHz9QFjYWbC22sbU89C59QrpW0pVK/MTD7d3Mf
TJzcbOcXGvdLef6qMnXbwcQNxU8KpgSpaHUlr38L/tv3GU5MH/XUjE36or+t7xFl
Ihlw4EKy2WbbBDLowAyV/Q+R5oXOnTjQ4Nc5eh5GNe1VAWXFr80IsWYvN0bKuquu
mNVWY9KfnE1hHAZmH0/NM25BdeyY0uDMZri4HNOlhGYGVjZZ4ieTWrTh+ua6ix4+
MSJ84WbVHsO8YdJngnPpBAvx4pSLWfxr969ZXdawhYIIrO/GoWg8qP/AxxbkD2TZ
3FVVwkQZPnP3N+zPOX7Frg9uS8dJMgStPGlii/K/8ZvYTZk5FyAg/fDoj43DQVvx
+VN+Dzmn20Rm1JO6OjuWO/uE+QSiw3zojiU6UybMIPmgh+25q2acNkPjbwAwnncC
xCn8XdQIBGrbvOxRt+7YaA0to9dMpy2zUNHMCZE+mjUOZY9XaCOlsdQQ2RZIQwLd
Itm/W4xbGz41RdBCTgmBA1pv72JPQ5/txG5KBtNfUDpSCsclTWAhZCiEAHBX5j6R
AvfrAj0pzbLHCuMRBJUUDROIABhhOevMfruPmU14jLyZF/7vnKiO5lOJlC8Vp/ln
eemMfpWQnPxOtl1WSssJ10LkMnE+6sx0qBzFh+NCaV4O9R2OzpJyBniNA3GrryVP
Ccqc3JhSl5Jyc0ITEcFhpv0vVHtvbueWvZovSwjKa/TwaKBg+G5YBtlhaf+xRBvX
wwiDjUFPLkyy4OHDosY7fDT+HJTiN7CM6Fddg4dDEcvqsdLrFv0XZQMXDaTY2JJt
TFJiKhe1mk3zVi1xjaQCoeV/j/rsSuir8zStxYaZLvXZu7pzIzaWehM1fV41PuRx
3qJ4DKTWM0wS+SuqmqS5QX4rCs0QvFr4kbRcUowuxJyFSLhYDvD0S8uFmmpBRRz7
OgkcEYChIYc9R9PEWV4OshgAtWLHepYaREr6bUznbKGORcz9Y19elciTVdMWk/UE
+6HVwhtQCvbu9yhcxwhkXqhKE8bDf71AvNMgb4QtH3mgmIxqZLNW6wk0VvJPnaVx
9v6NfraFx1amdYbj8VdSnUPGh7MeyVNCS/gQberO77AzbQtVak/t17vVol6p/pD5
TqzJoqJS0Lge4I18CcvpGSHWbcahI6IkxNKtx+pSO+VYp/WJ7GaeZiRPe+W9ZJ9G
hMdbNqfDrrbHRLen/vfW2nxva+vbMhhjyPT3hHWnDR0aNf+LWHzK/HrLzWu+OGSV
K6H/QZHcuLJauj9/eM5AK1ry4eyvZDfVsNGYymB+sJwSTFb/FQTUCzo7FcON1dqW
YK28QQh9NTdZOiGtazjCy+v4IKQwCitx27BTRwYmUzeJUHWBfi1eqqsxj9rBvJh8
y0gdu4JQL4/9bFQFs9gcfU182Ek9mcU5PjTB4JAdgjM9FeU8BAbpEpE6xZZapwE2
758YAwCq1iR5sZgxBHvMp70E9LKIgOoB21L21BiKk9rOv4cPMc03Sxunk6ztTQeD
i4t/XB8h8G9WH15DcLIiBOa7WUPCKb77d3Z0KYktboywTkz7rpbUEQvk9fMkJ6rM
jeHESQ0+YqED1kPrb+90AA57IB203xCXOIeUYcp3OHt8qxa2bFzfpqnLNhn0Bozi
QEU0NpayoXb105V1RRPzxvR9cRZVf+byrj50j5lSxjVaJN8YOILjprmJBkHt6nPl
gzhcHfRm3+ib8BLStfCdH7MQ/PXp+IXSBEckzmEGLYSMum/8qdjvLRu5g4MqXG3c
KjAS7nsA0P3ND0lupwHhKzwIX07ORD86QFnLf49JZVEcvfvXNbjiW/Sr5l5PcfJi
ZHlciMA5adUJmouZL/liexNYqA7+7Lld+7IR31AX0y/jNcxksy2R+GROj98IEe15
h5mCtEPSpFxD+4/f59fOy8ExUb4tUoVvutVT8On4BDuV9rSpheEgok6Z/sZKcf0y
aR/cbtNg2u8t1xbRhthnPgS9BbLUBXpfJhZ5HndvqKt4RgcVq9uSrtbAwZHW3ooX
1rWQRAKINk4renES3SWYDGTwt2bAFgxuVHwyrh7SbGToc0p1UZoUEcREj3zgTJ8R
8VMiLjsSZXxyAu+GWYUtfDRLeqWP7wCRddeQe3QT+HSYHV/ihZrVay+SwQfsn7xd
bxWeBpz6nwOqtjR04K9TBRzb4eyM/Ar/WzN2JNAyae3lfKOrv/zdfyiKDiNdqrgG
IjC/pAs9I+GgG0P3Nm8S28wM54iio8ydZnmvEdz7FXHaasvUxvJjlkjNNfLFISsT
jbbLSHcMdERYQ3GM6waF5j2tPQGageAaqpC0nJttUIzLJ6U1pTLF26ZrOZm6Siyn
w6TEgMSmFP6impqh0Akxg4EjnCEFQ3p1KPiKvEb3AXcQzuvS6n4NG6uNedCDja78
SZW218ef/hToIltsVcOkNMmBplToWZwx9YpWlVI5ZSLHtdEOwJJeW6HOdWzvBbwm
PQKt1PAuOp8L84zuw4Afb8KG9GGwj0CSTi0gajtMuIy/Sgwv5t4jp6E/Y8qxxNNi
3mwAs2tznycaB4PG18bd5OUOCvwb6deeX/HmvVd/V/lE3Jyhdl4lnWn+K3RZEuxI
vkynnKsfjMM1NAjbkFJ6B52PJICPopM0JtqHcfI4FxxJiflzeK7Lw906ijBFphjq
w5aM0sGMQs7PQ/VFuhwBVwymkiGfLKQBbXWvGVU3fLwczQAQzOrJoRhIMCQvPxGy
k6b4HoisxeWoc3sEOEsqhx/wPqbrT3QZehSMwG+Hg8ilVF5Oftc9rvikpiyowZUq
9z3CX61EZKgVJWRX25KiBMG16DUr/EvVu48/oLs/oL2qLiL5sDbkLWSd5Eeu6LLR
QIFbxDtAqTtohWHyat5KYlLaH3lUHQuKaUzv6jarqM4WstJhLeIEmHILY/gjxVek
8lu38/4F9J6FqQVEHJnju5gnuXEPTqNi2fZ36cIKlR6dsJ/Z2V2NeIzSBUNnveTm
YTHRERQkUi9s3bm4P/xpiCD4FoVcOp9/41NXhGGoVqbXo6UG2D++IWOm0KYDZEv9
f70NN1UXEGI5zzxPbRXGtJrOHxR/Zun9e5AoTXMEvMYskAQqCZoAnNYFpQYk7ma5
vXu2y5+lQCSGBC/pbW+oRMdiUoy8wOlB5b2My2fOyiRQLUs5ptehAnhkfKJG8+Ni
HTfbB5O0aepMQLQRd1tk/5FrlHb2/s5oNyR7kEiXzp8EJanTIyHSVNCkuEgROzxh
A4kkpC2GFEFSkkbfJuMnylDc+RKcu9ZPJOei2Bd4Oc4xn++rwRYp+D6XngocjSwm
GD+jPRps5L5D4JH5lW6p2iuGkRK2rd1ChuR1VG/PhypKEP+hpSvMXvohZzSPpSQz

`pragma protect end_protected
