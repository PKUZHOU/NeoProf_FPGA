// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZeOSfj3vxlaDVpaEaSFNv64mjrBHmd3RMcI1Q60HBWH8jWtmOiRTG+yn2DHP
8MF5omVtg/Ed2cr0V/btD14eRUqA+gJRSuTcanHceqp+74iLtFnOx5i0dZVz
EMEtvmx3FAWUQqzRt774yMWBrKUQV/bA0hAb1vtNbSi7lU7t4nBIBLnqcEbH
ZU4tBSBAFyjMf7OPsNekLge5ezZx9uUftu2O7rcFh6ZPMKWFqFuPlCKg+3DP
UOVal5B4fc17Ryn0HUbiVBgpA2tHY2w1MSA7530BQsby86oqFlGyqaz8gusd
oZv0KJNheZN+Ouy3hMEw/+6+b3yMTndju2zh/WGuvw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aJMEA56UAjo6KMgBZiZhuJQ6uuo77/PQo0Ylqtzp0ldGf8XPrqiiHw/1Y4rH
3ox6lDKhJ40dY1HnXtxv7tWpJcZ6bP4zEvmgawCCR+uCtsF6qcSLhknl5E+q
uzc1xKsU+mVB5hvXhn6BaL7E6anTi0Sik7+v58niC9SMG/eI1MjmsB7DWajq
iX4vzgZhY74dj/Ew8i8DPovJFzUNlSfCQs+kIU6RCLtpDv/o6ivMC3M/IebA
VMdxL9Be04ouE8EZtdNwNPgOmS8DWY7/pm3SyULcnD8bW8FQkKU6D1HrlRfJ
z2eq2Hx9xEBH/zFVa2Iq3T9+inX+wJJ3dPOO9eUV4Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J7AFMMTPqYBv00pRqUaCFbrPwi9A+c0lqBDz4XqekKUbMjchtUilrvsLxVCm
5tcwVqPt17uDsN7+GMOGrUIWLxINqzahpFqeVGUQQVtMpzWkXbsqngMswBFl
DcEgxF3A9ApT30xqHVjTB0ZOSEgMVo+wg6Ztt6n+K/OSEBHpMF8CuwvMRQWG
hdFcX4pyMJ6g2WebCggaxWb16Fv6jt+hsY3Exc79omQNIFKeP/6wNuITjMO2
vOnOAxUX0uRfjuSQAO29RBZbPRhobtqinQsT0cpHgooWKWaiMEw2XkRxFZfY
uE+neUrdagA1tenL2srPAzaehNNDlumLG3RYNfvC8A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KdVpL76eiER9wxdj8U5nphn2iJN7NvZKUvSv5kx2QDcchPnD/CspFHLniO7H
KPB/LKlUFK+JnHYZrvQ73jPqvhc92wqKy63Emow/EApU4G2ImEE2pXMiA5+u
wxjis0RzBu79VwWPy7Fbx8hRf9Hk7GpCdeLfsRP64b+Fog2LC7Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rrSaKvqJ51lqf/QCRFx6D8+pCYmcZFMQM+uRq2/S9Gfe21jhjwLNSPPjoZhs
HD155/Suzxkovl17uqeZYyC1S/8LvufYmpuHj2j4HrHhnhiwHhNt1msLENa2
xs+ODgzuFyOdql779fxO2u4WjsXmWh0++S4hgGPON78NnBe2TSkH8sAq1R3n
eVKkTi4wT2qlrFcEZcaqyI6rHAozd6R/8hpE8I8CAWoTvnaGEmYSihmStXk4
x/PjaJDSyk3/LTBLm7K/8bQrTlsAPIxpFL8n7jpc20deQJpnsnBP9FFbO6Lb
AoikoIG914jLg+ZRHjl8xtpRzS+8VB5g8io3ky73h7PJaNqIAl/sgJBb9rXQ
ImQszzvua5UYQjvQ4ODnTnrRKFqej/SFWOi6J0YkQA1KMOW18bxGD2+Gm71v
JghHqOud4ScFA9ZbSZZaw1BBjNjBW4jNUWltc5X/Y0h9NJe74rLEoRq2zJts
SklY+F2mz1EOm5fwslYLNcOdrJRECFcy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mr5Eq/1IGWJYgIQzelzOU/XYyv7soiGrMcm68otRL8NIp46t+qzZq/75OJFo
ZtXU+seO2RbkmHadQfaC3foq3tiMo8ekwp0kpLS+g7rDE0aGmmo3z6C4wF0N
V/n7SBNS5dDhTszwn24HZKW+t5KF+VlrdGdS3rBgNJC3uohY5Ks=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Df5vgEpdS2TtQ9RR9FKurepBO7Lu92uohUajMsAB9dda5/scmoy5wmQRhs8c
v1D5z0JbEPf7vmKFoHnQwgrwOvQP2pQrjNFCMyw/HJ28Lr57ZLtpajSj5KmQ
Ow5GSlJu8k/7jQBYVF6LValgXP+V8qhcWR+MuFUZrzK3BFSbac0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2112)
`pragma protect data_block
YwyfLca5LB831E2dgpNecL/NvrFmTRq9Yrq/+cfviDh5E6fcwzfpN/PC2Qc7
NJZAjuJj9Luc/Fl7L9Rsxj2yHRuf5WzZoCx9ar43QDJxGCiEa03BztfZpVYH
Ys3p4DPcr1wyG2NtNTjIGpPzKD05rPCjWw/3ggx2c1t2IKn4Si4uNBJiG1yH
N4F9O7t4scWuxaXa56pdaUM7oz6VkbtIXg5K3yo68fFvuzOu7r16Z050HQsk
AIG9OBaU0IxIwx68xHBcbIEcpljUIuBzRvTzwvlr8QAZLzjfSj1csdEXdWi0
Gg6Rg52FLE6HKzmE9qBz1bVvDqAGmDpgr01meIYns7TknJU3kilZ9N2ob78B
FZ3WwwJsrxO+/UiANXwcnaq3VpPzTp25ieQDHRgU4PubcH22n1nZ0Wv6FfX5
spmqPkeYkDBEvvTyXeDI4AC9h57H3/C+RjPdyJxEz+9vCknZfyR5MaTEtbMO
QD2rn5AVuV8US++9Ocbz7EmcIs2YdFXzezkuaPwb6SwbvbswoirV0PtrWKLV
fBwLEJ7NE0BKIpSDplOy/idG7+E22V1rcXPtm0W07etxxE3ubehk6zqPQBaY
2br6iPjBN+h+VuOQcLceSe+dZrFsZBoWoEsYarn4cgyFxIe0155WQKSYINYh
3geqOlmOg6MyjwHx8KOLnF5aU4qNID5OSradFfjLy+LsLwQmvoqhT5Su+WqW
DOtGixyzvdXDjWzq+B3RMuB1SitdrlHT0Kq6H/sNMACEC+ngXCQuW7qmuhKp
fs276/iW8NDbeXzKEgklFDnvTZaiZH2wcYyHru5Pe80DhzgLG5zzniK6OuZ3
MeL1oKvDbIowgSl7Gh+KiW9UyRUKgm+XZgqqK7SN1hubKuL2CWriZ4fpVz95
Cjaxfv607tuogsMP5XYWKwEisnroHygVnnmQfmIIVaKVckh69FNFgj274S9e
bZI3n6smb4tR0cARO0tYiOBtavj44u9JAt4uVY0Kk4qmNI3UkDX2SCtZw41v
opyBFb7vIEfKJ9WXboIev4sJEzfQ0Q4n8qDySWK2tfZK+caxFdFyWQDdVxxF
+TiWl6PRgmPjU5Z3LTGHQ4HIrQggKas/7kqQuZ6tUKbAy1m5v2GDBCnuvwOy
BnBMwBSQY5EPkOY/uYuUbQLGaFNa/c3TxKVn0EzqRfWt2UG+zd/YjQydiszw
xm5oyjqQYFODMGxqksM6SLgtWePqV/Elcr3gctFuWvJFx57RFi2GIqYZRdxK
rt5bOCUzELd1PzGjYl4nGCIMZlZ0BNPFTVdz52qgv3lZz4NXudA733seKdiX
/B+AaYRg6OH0WmyqrKb2uLVEcsz7dfXaeYkP6CkqRCwPz7iCVuyWst8SSoEE
WTnWeZlrsCOIGSQkP/necHOg7e/z/UqBpNEMb/LTpA2n1rMJGDUFBhu73OV0
1bjqI71g/U7kByE+7/3mOJj5DAWqNX44t4EvS0toGp4XuxOGF4XZJk/UiIhz
TWsX5wmU6csp+pgKB3GJxKWnIXP36v+bB9V6K9MiBDBtpaqxVRw8aa0QHROf
BGw7nl21MaS95jHRxDLOwbJ1s9wwYni/qFzbCHuzkcVocgdccRjctpKibbA4
WbGqJF73dNNDoVJj51QVy06mUjre2clGg6+WtqeXaaWXfh6uEu75WU2V3Edc
yaILmZLtAO5nz8/hg9g3sqCF3WYSFR33PYr3LRoNzpQJF+1OH3+sb/b6w2LE
NyoZjXjlFuc/BazxIAneVaYSA5Je/iOYsn02gBjpjKEp0OeoPgDPEUDK7Fzm
mCAWxJJ6ZkgJtsWRrFBlG7CmhhlSNdQ8RrF5bvCj1/fexrD5azLTi5rK5hAf
Xwh4pZbOeIdqVLRtX2Q4oWe1wtPiEpmkoF9g4WYzQ4+3y/bD2f4CgqIL2O8l
7C9Ae9khNLt369gMlF4siFHaRx1iWC1VjpNm+Nyim5CzW1vwlc+PWkn+QCof
TuLoTX+l3yuNphjziIZOif9K/J649Wew2pbKTcY4puX2WKIs6LA7ThMSEqv0
Ym0bmM0k3LXreZDr2pn0arnFbmHEu2NoAZbWvP1zweWymfqW70VV8Ak+Raxt
gOzcZMQV2nLM97fvj52tkdbP1S/owY29o/sleezuwXkSfz1D6/2Tw1yh4YD1
NVZdpIto987sC6u64LcZyrdXWNPkBSTuXTyJzYLFPp0fWztHClHcQn1mizbH
o+3csK/SEtiid9KwrLFFk1KxJiNc1ejSd8k1wkI2NKa2iwm1EGkRzPglrLAA
hwZHi8+Ur6Osy8w14xCSCIGb0R1qRQ30OLmjY2tP85WDvhaCqhqRkQBzUpBp
AkGpLBfpQHxbtPrFmE9Wdv7ShL/RWBFk/9Ap53oSZrlaX4P0M3ZqnlowLALx
RwoVyJ6AvlRRKwXjPZ5Iiu7Ka7kvqUO0ActFbwZBOjPmjgps6NO/1XuKZmoc
9Teucyb3akBVMVefnEpP0NLLNMW9zAlIeNQyVKU9Y6RBhAMBG/+1Ef0zF4y/
/60YirStmUk1lvRWe5uzUnY8Ma8FEj/3cCoWhZJE15oPdVWvH50PPHITqbVL
gZcVzc80+MiMj3+BM9mdqrdiN+aP9fqXiaZfDwS8zhAIBALjWHrBRXtDmYTe
9hLty1rSGSF0g3jooqO75uGm49fGC9O401pFj9Jq2e9VcsolfeD+fD3MS1YM
zOqDvBu5qoLkdg+X0xbxpgOdCdlfpp2SCxrO7fhiKCYr9ih7mZvAj+usDtSt
IT06kWipz6V7gXT5RLsm90QK0Dgp/JFXtD0wvUk26txaX4RH8cblW8M7

`pragma protect end_protected
