// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
foN9r76zP/uPC0WQkPeQ3WlT9liHx3fvI/kranAnWO+22uciGCOXl3KdV3O6PuB+
HvBW7tDZ+lv+IObaQIIn8Yi5FfTkCHgCPuoHM5OmeV7KBgQC6dlEHSQXuTFD+JIl
Bqak+JRSOo50qjekpnqM9zz2z5sZCtficyRD39QPYISAOC9EskoHGw==
//pragma protect end_key_block
//pragma protect digest_block
CVvUGSH2fNT1p2AUG3BAjONw11M=
//pragma protect end_digest_block
//pragma protect data_block
oDI+r00daFAdAJ+1T/iwS1Dp24ViF/kOeGa9Y7Mk7ghYp+kfAQb67y2pq6SFbJLW
NcxZ2ApGmdXkk74JgpRMctLKjJJOdEHmv66zZUaECztuU7imhzsXatXR2k46p/SA
gjY3FpW/WhlBSDnTBmS1dAqswZrr4osl6XS+DEHowUlY4/4wmc8F0i+6AejFIbkm
6EZom7l1qnmGfVDcjaiUN6or7vHhl/fwzxviYUue4nwnr1tSS6UZahmy4lXtFhLJ
Vzvwu0nEmoQ5til38dx+aFR6Zm3Pge2aT6RHZ30dyOTi7gVDW/fxSn/kLheJQtk8
BNHyOfvhgYqmGoIZ3x88POLSBTv7yqZl0CjgYKyU9erW0i1GaIUyB2koD3uVMuiS
5fce9fQ9zxGmatqKp5+Jr3XFlelhzXFdiKkw+QS647IXsxfyZrWQk5RSe09DVYSw
kRL/s7gkqGerfX/334ODaugH7JgeA/CU4ImqvJYEEGeY+mfpFJFS51eALToBL5gr
Z/5h/XAo3D5i3v5+IWu+23M9Gx1tlOVgpnhouS1w/1p8nsTv3RBN2Wp1wkhvlwAZ
jQMfDCUYcLU4DxO1DbxrDPSJ703EFjgTk6QV+WpCaUw+zC07KntBv19THGEu4ZA3
9wpI2/vVzYColRpU2VIatdRRlqF0Z5JdQWCvI0kjuhOViYYxdqB6GaPw7jlvDEHX
oCffopqJEFQcGx2qUnEuq2iKVjUXv6lAefwp8n4amd8KiIO+ZWd+DTbkN8kbzI5Z
4OucGfkmffJUu13m4zolxaYA/i8gLTyQk3yhErWGfdChAdX1TiKGioyTsmHKoeNV
9586sUvIlfZp55/Gq80MZkTPvWmnGG3fnTdEHevEu5iqJisCrN497Jm6hCEi9DLk
TrSI8rshh8dm39a7OsL1TsneEdxRm52L6JMrxh8aXKVUZPc7ABNao73D9Z3r6c/g
W2dGZPwc5CMOxc1Kq1zFg3GpgRAahzVCyyJOFiyp+yQ/epeGAnVGNO1xIRzXafDv
6DkLe9X1fDWF/Au8t4+6PuLhNvu8WyU3OdFmB/So8AyowCZspNQLmhOYkIMSp7Lj
h5rJLGXwOr8B3C0KpaJv16Bdvk5huabKAawIfgI9FZCWKktKvM6omjEjmtj4tvwK
jY/cu41T3li82/3uuMZHOs9i7hp2lVixIxP3hcakWqlC5U/TeWqwmEaGJGuHDsoY
PX7w04/lqO/mMjOGj6cpNGg2PxkuysPh/JAzZhTBGds/De+Ks0A3GO1H97xexzDq
6rP+nTTuVa3C+Qs6d6yZ6Gwf5G7T7yUnCplzXyUxk7JZ52TS7QvphX5yECnqVyCg
f/sM/8dclmzxjURlcMhYF1YbC3iUb8c/EJPlilHUUxfrl8sWIJSgF/P2gAAiC0qq
CGd+I5cDD7gL0Kh+ysXqpbd7YyJPuas8hvEpfaFhax2ZCpRSCp3zCD2nTJ4mAK7f
zxpFpYFXHrrAkYEQuSXu1K9XdyAXU45TrogbprLcBQX5XMoD5mDLD4D/bJDOzkfJ
Jus9ilcysLNzzQ/2SX9qeAWhdZnkro0stW1h6bfF4m2HbjyXqzphwicFpncjJ5Zf
owe1hh9nxUdgInoDXM0hII8CjktnOJyKTESzIK6VUM9Dei3gMWKkTooA47YN6pga
YxoggwpO8icI2E4ykCrFLKZ1z0iyMxGnBTAzNRvUUjawlP1mZKrveF5Jzf4EWKlR
M/6cKd9712h9aPgirZSAESXGG5hUNGJzVAyWtn8RGK0lzs0JBWR4JxAf38nKB4Lp
WHOizIU1j92Eztgimx3WLiZJskROH6ekF+T87bh3pSXXVQ9C0exZbOriL+u60Hmk
ti6UfX7KEtuW/mbE+hVTEE02CrW4bRPoBFVDIFxV2Op/A6yuZxFuJsGhheavynOb
zYlGYvqNqgO2Ha93zrWjsiMPrOItREuckXYWyCOeQ0Gzm93uQwuiJtZHGMMY+sYB
yBpCQ/O6aG0HAwg10cigkhelzT86oXSNsQ8SMTHHY6CuWMrK/fHy/FLBwpUKTO/N
k+P0JDaFU/DJLGt3nFlFuEPzG3T6uBpqewt3i9HRKozWruKIitdgypWDJ9zgpUSJ
Aa3XsZQBuRtGJIQIwGgnSz5hYofcY/Tc1YpOnBJcPNSeQi9eadfwV8c5IFrDBhxY
anWEEbKR+PZHvq2yHGKwAOQVEf18bVHryGOz8uOUfh35QuVCE3//pH+VhQc8qxNR
HIxlqksNL1ioEUyNwK8af+dyAYVENOHjkG1tR7+msFUBna023PqQbg1b/GQUAtEj
9B2mDEIIST18yPBGtLoSQJYWhcZvsNZOns2YqCitTQKAusjIZ/cIgqWeGpEKTKKp
LOdgCxULw13J7uS1ORUnKaG9a7PZzqqveF4rElNs18kIaCxA+zpYK+cCodTD3tSc
wHVaHlDfme07gLfzD9f6ggWmGB6SbBbE/sgBfWmwe1QZpPdbaAILXRpSGr5zzVSV
Z5ydeeS8bkK7Xr9lm6F74EO5kgEOLuqgaZXZNisuY88/6eED5Q2McDaRqoQkA2wB
f1STSPj937X5M4AusYbKxDKFg1iuiWvBqeJnBLBjMx9NwdQ3xsgFBOq3BpLF2yYL
5Sz9AVfY15gxp7FRecSGGvON8+3/UiIEXuJ0f59FjslTVERkTdHvFi+pW1qw2Nrn
FipPUwsowXITy4u2O2+azmvxEZvlAKqS/N6HZWlEktQK3pEHvcT+nzTIm/1KUOpw
xDFRa+DmyG/PKYWlGgGcXMr7fWDvlTk/KCTo9CHLrHyMJojw8VFdJmEq1YYC8xdk
j+cu7ja5PWdwKW+dIUijZSHFT2suQ5S1RX9JqVcSE297OYUGwBwwNF/pKwPyrttU
pd51l8mUuZ5nIjO8iXoVQHJ4vuiKP42dNeQ4qLhabf9roqf1MJ5no85gBcoB8Vur
DZOv0P0EMgTQQQRROUjhumxcitymJ5Cd/UkgdLFyNhGnH8JM9/7sI0aWSKnaJ9BR
6g+COQww6LtyWURcKMaPNeGT3RlV9q6RHZeFhqbBUzqbXHSBTVu8c6Sjcpk0TX4Y
fBiSzM9ED5KAnQ8wQHAemul8/IVyOEaUk9o/ODGphkmUAHgmoxQS0u46IpoBjwpl
7G2LuBext3I8PHkh4csNw9C1ouSiGvES9VCaUAwIJY+b81PZpm7dA0/sPzaphTDi
lU2FYd7UotDxH+TzsX7kEtJ3hwXIvFqrcSDeBCVBMHtNS1AR++9I7zN8WLzlhdVU
47pkyCSEzND1FVHBVAfPEkHsPGKxkLRYlRUqAtzIWWzy44bEQ4O4Q3yhzU+IoWF0
hmFtIOhlNcos56RqYqdg+MHLRwUdgLk1NswunZw94dKVf/0a/CCqWne4R3/x+Zit
0dT0ByyhtvF8xiw/BTGKOaLjV3FPhdeFPtoBHUThlr3T+c2qIkEe0nP2IQNbMWN5
mEZbJtgqmIo/oOEieuVoNqTJJ4W9g0vHFOsxerx9mzbW//czR4pXr6mWFGcAWgd/
tBxUx2lM8DOOlcz7RWHAieeusA8gLXmUN1ZLmCetXIkfRs33O/+/x9DOa6KgEkZp
feJ4ypZ+yVSt/vZhmhGmPU5ynZAPMbdwF+C5vrTYZzcKg/rVndP6QEd21lEd100h
oL0htfGuVh/H9BNoKXIasIunxF1T36n06V8WHaiisk3cgI6YhbudqrFCAR5NdT+5
Wa1FEhX/VpvqfeRhjKEw877L6sQ9I8lIDum0acw7WPLxJhrw36TN0ljNj95p6/D6
We1c7Hlo9d9lVZvEgI/v/pErnXto/clkl4z7/uKGBhM1SKl8LCmKVfl327SJ102o
9bHOsP2yJloWG7Wlmh9Iyoidx6LRzPTd8eKBjvwJ4VC/yX/aaQV9FXsv3cviXm7j
YEB+jdQO4sZ/trETW4Es7YM/YhFl3z6Tla5vkYvOoKJpXcgzdrwcAoE0/Gg+uARt
3GbPNk76saKYvRs+38KBHrzYXfELAHm7y9at8sWbLxuzbMGosR3n+Ks7jRQXmb8d
6L2CDWI8eQoWx+eGwwxrUqwDLuuPtOeQqUHZoC6PzwqbY7dditpPgSI7uQVGgZhV
2PvbAxfOiELIdHRiUbjZzeEWBoc88Hn1nzT2IXoOmeuBkjLW+dZEnGupL9dfMcmi
RSFY7cUZ825DOpdLt3KEnfP6nYIHapWtkMGiJq5+XZs7RTCwyjlGMU5COp5QP/oa
OFGR5o2Bmbkl8+zHTdDee6yWZG+AsRh2/BuUutQOUlOxEElY1ZS1Hg3W+ETnJCu8
cDGLWKvKwf7XfUJYsIuaoxZyFXbumUacuayVveJNO1oRimBF4kAKZbA0wghRtg1M
7dnGtHdizQzeBcxDor8o7Kyy6mLJfmPwagMy1DKM5IVCBRQDRDw/vK9LoeSoCrQJ
H6UbJUFu263tX6IZ0fSgewN3guqETQueumPPY2fe8f+wsluEPFgqC+h5v33EL9lJ
JY3w3DeAycl91BCPWEbDu6q+3yhsj9GJcJYlkUoGjS/6JZ6rUyflFAj0LHKjylkU
5+eSs7aeb6PTxytLIphzZvW9BOdtjaZ17OInVehuWBsbWjZQayERf3C3Gf5dHIdC
2IUaFmhyE2UQrzMopjwpnpEPR5/2N2O+8KmprP5OK6jEscrorgg4K4pSrhbxvncS
35gxaoUwoJWdJvXwVAjZB/xoi+4fiK6sCvu4Wv+w/32oiUjGnK1KnrA0jXu0zm0q
vHLvAu5rWXYlYCVhbxPk7RTIytT6nLAIH73nQrJMpYMBB8JYgbxWj0anIBSNBdCP
W4JC+XAd8N7j4E7ldeBtSqprcTR/9WADPq02Yb7I0MXHKLmqS/1tK2mrKjK8WxBV
Q/nalJXnUAu/pzmA69E7t5OwxYITYPa4cYyk1AbnZFKcBDrdsCch2EOUqwohhb3P
cMeyWYhdfJbL19JoWaMM17aujOZRB8hF4C+xmlKcG8d+fsAzDhmjIGMt7YqnaKZq
1t4a4FFKF4BschIy7GV7b57kslyrIhpWkOa02GBBPm24wXdbWg+2/LQk8emq8vyo
34LMpuvMD2jWDFqTKxFz+2MFEFXPiLZIG53Oo+bevj5Hp4ONh5q0jCZT+Y4FUr2O
LWnNGngJgyeVq4yCxOxctdlEgLmIG3veKsp9tM8x/rtPG6I3rlBGNmZuA7NWFFPy
jjkREHF8SvHAwUtwyq9FQRwctI2/t9+vGXhv+E37d2TEbhS4C8H6bAHDDhv4Tafc
HGINc6eN7Iu4hiwSZsxImpemUgLnTawuL8J4F0yAJ5SDIlslFbmId5YReMSxaD90
tRZS79uWp5lNusZTwW/Y7JU3hoQUIUKh4m4jnzj0XPCu6sb4nw0nC0ZQ/ylVBm9b
//dTIEnXFljJhDgs3/l9s/96nBx21pSoLFaieoLmmRrw7QKbcRL8VJyJSpsSvpu/
zCFpQr8Epm5xT++W5x3DEnVvLI0vlknViX3K3kt06eJf8bznNL4Waj89lZnEcE74
3d+TlB0yXClmXHoFXROWchjnhgGZDQcg/oonFRx7elc31UjJCM4LaJ80CoXV7wVz
R6+kQUqS5zLpmZB9UfxuZeIcbQvlZNuPAJiFexca/qw5R5HSzWP0BT5NmmsGlh99
mapmig64EmAj1zgfJndd33zAT4eclyXllUhkEIAKv/WSpecuoqk5tGwaLXKodwi1
U/f3KG90zt5Sp9yIV9wcWQV6+AoqVTqs2IjWHiXk+SZeeSmocJGX/i65Y3omGOyg
Tm9vlU/Pe1/ItPt9OF3WWoCU4WxaeBZSXLEpHuaMwrFL3KOoOV6BvNQDlTUMZjnj
vo/cCPXw/COZ4q9zvWDDeTeCDdov26mST48fJofPoF8aVY38DNCqRw+We5WbjkKq
niI8Kdo9A6io7BWRf1xgI8uzo6pwuHIpi7aZmkG0FJ/RAhNsorfGYXu5H65bsLAX
vkUjREgj50Vql0DgCSHJfTLQg0cxC3E1U0yCrS9F+UHszkKtjJg+6X1839Wpl3Z0
MkL1McLTeOWLJep7jLYWa278lVjZxfgjyfl9lakf6mQCNvTOyRwxJVXHFigBrY4o
flDwqLYhfbdrzDQpmNAX1f7qwd5JXlzjZmf4yalj5daPxlBnITSE9VSPtY3LpOeL
jOVcK/xZyWQ/kRbp5m0og9PDXaKTnbJCFJLaGnuGcBrPQiXulhAKpQ8c5PFFXBgz
yUP0BhZcfe84HpjthCTdCEfTOSbHOgGarOYgMvbxTThHb05EqO4P5EamihFjS8LF
kTXYm3qk9e0okN4lYtSUYQ/NUfN68CfzIL3NcU8ZKOd3U7/Grlz1pYNocK8gGXGV
mt/yiNYOqdjB1AhsxfR44R13i4MYSuGvHihitXdWtdze21UUnZUVt0z9zJlQWV5B
yiiyLb7Snb/Ve9dNA6+CupmN6YwRNDBekfh39Uta8yaJ1RgemOihqoO1wj3qTwsZ
JpjZUPYX0IerFSv9S+Vn3o0TCrAnHe+89L0vH8rmPMFLcOoc2G39ILJDhu0erAks
GONr9ceV/HzZd46poOaIyxLlwukoEMZWKXBW2TfhaY/7UJe9WmLuZqLZn8eQ6Mnj
ySIUmHqTtTWnbKYEVYOqHWaxMlVipjJrJYT2Rbw8U0HyjokL8xuGFD4YE09jTwrI
GFnOxiiyRwFLllt5SEAGcUg9agptULTpvrOc9SwO/NcDPZubNiKyF4Er60bVtokQ
mvj7eyn0jt4fZfOYIUXhwt65uYHcwHMALNCs4MqnDk2M7QXjZb13GxxM7ZDMc3OV
XbkvDc+SIfKRrZ6ndoW/EfVUEpRi7Hb4UZN9Oe/2FgOi9ne0oVhklpii6reeMuRd
/VYDmxz0UTYgqF8lWy0bTinYWPzoubLlQKwQnXI43dj5/W2qSUQLyyhiJ07YkKb0
cqkZsAcQ/jek65miyQ6kaUE3DFn4Zbve9xxSDojkhSFwA3zJ3z9B7ZoZilb3KcyV
VVUpO4awOHaEPlJSRLXZfmE0EobsQs1e52XvjqGuSUbtILeOTYvQFwhYxnXFw1A0
X8NZTQ0QbHjPcaVOL7NDQT6eoCiryL68eoqVpee8kIKDGSfvn15IsqGF5o6R7flC
zWUnb109aAqxqSv6ROKYlbLtqvBktZiHISXZEOzHKnrBgAJFOZ3CLo/yFssAZPWj
ceMmy9pxeAj6m4gSifOdb3YLMT7h54q0b8ZGqDtCErFHclKAio9F6lv6SeP9LEYg
wE1IAa24wobl+ySvcXQ8/Yy0R54nJhXTwrU+4libqTBmWXQZN/iQlmt29Q/jRjtI
gBWkNhSbV5ARZ+Iq7DfRNN6vdXz5laYy5ritcfrpp0jgEZpuTGHSthElsDVV1E6z
kjHwoCUVwNjEYDLF9ETie+14cSjEfjgjI66bDPyoduuVa8ItI7UDvat3VyMmLESV
Pofe+jma2yrup6PVrTQWz/hdyR4gAh6KMIaE3hIJM2WZ6yMDmfSUunD/nOZdEKyz
sm4+EW1UhRCg59XdwK2VBhxmNfEgkGxpq84hiDXEyuXsUCRbn4I2lyPI1bLFj+v6
gGjl13vEOMlfx5qvvfVgMndidakoE44qgrZFGK/nsGksczmr5n7Mo64MAu1qnO9Q
NpOgsVzj2cSgC2U6o6BP1pdMwfzoYX+XmcQ3S+ptYre0u3XyWKhn3GPwa/LqA7dB
2k8QKczN2C1My3LY96LmrpLGGh3ZvXRUdPhMkAfrMglYhYutGcNdzDwt2eUD5S+y
F77aO+ACpY3cw0/+kvGtktBOTJYfXiG+ERGdLa/y2pP55wlTM3f+fHKgAUd9vaOD
XUTZsOb5p2w2F9XszprWcaq8tR8wEVZpCIWfrugvuQE46MbXv/R+IEuIyh7q8bKM
Ym0q85lxfAZTy1EhwD2liw4rKr8++chZiCs5seAlaei+NOXM9nwRB2Wl9egK/vwM
SJBYLCps3ruTvGteIvuANVBJVUmN00yD7uOuRukIUwTkAG7Mmr89yZUQ7hR8o5WO
O4zh757k0MGx+nWT5/F/mlF1RXsYV5j9c3dDl/0w/4FDxNLtjZ5YTk6n6djOO1tp
uc15nnGCHOlGtUiCLKsk8XqMAegFeJyfkhihZI6xPykj3tEK2LZ1lQp6jRPGuLwe
00T7uAFykYF41eV6rg8ASmSnc+1IFKeXiUDJcqs/J2x4u6J02MhHareYJi+2vyRQ
2wo3XtEkncEXwQzhr2BJ2Nh88QeJpXqEDDRXWSAX5lyaFi+Klqk331B9iGPe1vMu
xPlWnr7HZE5byQaNevIscDmOVgUqCddCaN0uCuXkpZ5F/FQwFSOtEGPlacnTof/Q
FKLSeJjOSda9xRzcJkbK4py15+63jvGIGD9v4CbPB2ZARUC+SGBUWNXjKrtkcv/r
Gd0hEyIHx+t52BrXMHXrSSfXDvE/g9q0LUtRXMMnFVDf9u9u+shY4gtfaInyroOW
Pr42ykJkIRub9tssBi5nt8saj5ccAO3K8+5ubKMWOY8kLu6Kc7udjR2ukpLwnHo6
IPHB1jUIR0ERI+JYpXzXEMYgQ1hTj0ca1w+XA0qzBFE2SK//M7cBLDn03xphc7Wv
N9CelAWNl1bfxwt7w0PUgqwLjmwN1cP3mH6YOXC8kTKIAjqGNVuLgWlkNmDF3rwi
AQOwAdeo3dT9sAc66yrJueNlcwE77BRwZUyhs2YrAvABEW5kPWBTb9CZDWhlPBJy
knRW072hLjVrkhLd0ELbaa0dqcBWdEELJT9hiqwVrh/POqBbtdqykR3vzNmO7Mp0
2pYRvjqnBKkYsdoB7FRSkGyrBS2XNfY1HWZ8io2dxOjVGJ1X1/hyOtTehJDcPGpF
RvLULlTXZ3tpuDCuvpsVA6bgqcSQARW4YxQ+fiQxYXRO5ug/nUou6AGt9lPDuKXD
0SvnIQcF2Hp1E+SYLnfxqwCqvaU79ttSxFCQa3SDansIioBVsYsTWlXOgVjEEPHh
MS9GA1RAq9xeig5RxRGAmllybFCesQsy7oImmFwqpi0F/9TlCouD6SzXiGTXBkHN
zLJ04fXeK3cokbcwxBUintMq+w3XIglZVJgi0+gkEyUOt3k6I6rsXV0OOEXS5jV6
Qn3WFD7Ydu2hCV4hdsr19vEAwJfxgqEcCkRxVkc1Cwzuyd8gU9o7dUD4kO+AhaF/
4Ns4mLWxbXy71okMK0ZTwUMKejcJtYtiT25TvdKwUerJxExkvWdPShL71DACIaTd
GH/uDRjeQCOkXqXOmhFhSnZeXRfs0oiMrLPz3FoFPDS/MB2tkTL8V4+XIxJRrygX
BBhOtqwj1Tp5jCOiLFnQ8QInsT2awSZ4j9JoFvTiNbwRAQFJCUF7nhk4JdQNhHYS
uyHC0eE3nc+N774RgyJZY5cW4l2jQyT/7ctnGRpuF3WFbJLPPDfb5wvaWu8iJr0h
o7gwLumzRp3c4HPoWL2S0uGaEKm5qjJPut8msYK54sMGab5XC/zm2y2qobohFyTe
jTROeg+RXiJo1M6fYsqbbkiKfzlMeoQqb/eafWnWaie9n/a+3sH40o04RmO9uSgw
xzKU0bN3Ommpb3T6Iab2t8NzHgGuY0+0RISZbxGOmX+0GpxR+t4+9Y/EI4SdfcvV
bE5LfALxLWXA4HBdO5WJPq2fvl4z/YfiD6w4JSsjflE26xKgFPjOQ0J+723GY1K7
iQS1pkOBOmo3haeObgz/J4y4WRCRS/2RtrCdOOhCbV95jN6cKIkSoM85rHRPo6rL
9QERvdRiZWOKncDxEvfKjEXe8F4rS0p8mms2NR9Oa6asw6dRkNWAv69CA+yYluQI
TWFSsUjoXkdJ6KDTDi9jRbg+5bvlTNYS3a6OZ+C0q+Sh1DrgocmjklEc0hEE+brL
Y2IsJwc1BCtjG0dmiooDZeMmiEC1Zdnib+oN42F2MAVLT8cwq8e3KpXCzJftMP7I
R/Yby+Fz8E9GaRiLEg2pKGZ8swOg1eh2N5yAoWtgLjKK5Bi9vg4eW85vvvF4YL11
cQ8b5W5d5+oSGKmXdsxDMkZQCC6ALkiERYLP4L8AcRQOmJUotK4mjD2iVMtw8qXz
An2J32fDQtTkozIwzig0DC6LTyP+4sIJQic96GtHc8V78lxzjE/ljkcqXMHMS5H/
xn3sYrVYByIpmwAoplrq+tLDcTHlFL9pyjjXClUMrKTrba301ahXe7IOQNd+rmH/
G8WerkV3PmH5s/qBm4tmI2H5REKLMPgNjUK+wQubsaKQxaXjrr9iP5FAUQJCPEAd
d4rUpOC2TqJyfhplUw1N5adktEfpHC+0vr8fkkEEiDWnsVndv6/KQrqGpQsuy1hH
r2n48z+1AtIxi1/3K5bWdTjaL64aFxeHTMtWL4kMa0m0woaStLWWrRjWwiaUCCKp
3eN0c2lMQGsZ1nQ1pTriJABKMMS9riU4EFIB4MSyw0yjOpVlgi+a12xfZi8bMZ7D
DT1eDCIfHXAQRHzgry49QJqOUxj5vBuxartXcxHAEg/sPDtcceFlhxSQmh464kiC
uMZVzU86fR/yiac+qguR5fotDK9Rpy5RnsOPvw7Rauit2M5vovzBD82juYSTkf0f
2xcfzH1osV7NtwhXv0MjPZoLJ190Vc+yWMzxZhNZK5T9jbNGWc6tLsBI7Z5GwzbT
Sr3Pd47Hrq55QMBMdNAr4Mjxu7JlWOL1U6MN9vDEO5PmaK6UpUdXjtYh6YPB5srs
c/xbWjCKzfjYbP008b39JBUIlcRK6iDdr1IpQcrENjn6S6AFXKG3UbiYJLjfPDjh
D6tGY8pQ96DcUdEYHnIvV996ovLJ7oTw1A7zhz6mMkdaG43Md19LFMwFPcRPJBJ1
ApqjPlMQvPeH/P8eBufSED/fhKDq6Kw2h2OViZhbyBpCHRmiTDwTkdVCSwyiysOe
Nwa460vSOQibSzmwmpomPY6aBG9kOYNLWawGFnW60dmM86tMZ5rb4ya9BZkc3Vvq
7J2uiGMOv3Pc2trS4hb+m4STUZ4nnUqrqVTvlIPqtcr+xyNeFL6pNqboPuxuHoZb
i67iGLeZMJCReYFPQPpH34SlZbsFtIBU1IiO1kIsYiIqLjVH3jKCrhh8LopC1ke+
lDfJhAF1jk4R0TyeDoT1zYe3a1rf/UQFKKtKR2RpDdF7jgEGEY1HlRnkhTL2ByfO
cJdQdRRAvso5mWqfwLsBxRxi5VdWydrY6YHIylV7xMosNI+VtFsjrHJc7A+N5sFr
qdB+ztVNa4oLN8/ALOgcNQFp1PNZfpg3aDd+13aygjifqKvtUUUt0cm34dHpgjVz
Sz9kmhn4v2rD8SeQvQr+5QltVeBo1g/VTXB4BxMXVlVILmSxHJ0gufxUHjwExxNb
1LI19gaml+TACXVYSOFvvbGmTID+blQnEQEEobksNKNI8xIaAnsPkH3xKi6LfO+W
wM+9zwC4RY9sJN7N7U4aUYB5EL0Ix/zMApswypi3FDCVlL8VgMV3TlWsLdAoQse4
eHeUyKOBtOsaS1WM3o+3XRseM/wvdiF9Nr9cCbJ1QVAzigrR2g2TWAIL5Yaq4z3k
A4AAvIcMerllKnMZ31H5Wxw9f38B3Fq2TT1KrVJ6bxRalPbCMYUTCONu25kgXxxV
uX5jMwsj+ldGo8MhnED/sfNmLP6AWzGWIjVZ+UIMkHRSqcVeWf3mypXZ/g/lPXZq
u9bPb49yjF5oqcT/N6/T6fqgTZy8XNB0ut6Nx0bIN+xwIZumV4AAF8T63HyS0e75
AqfNTP7VTMCN1OKnxYVELzQlEZeBc9/IHMlKnD3bTEvV857+GuRcmCIq5oBtST+8
seXAJpBFTY5juPOMB2091OSnfrD1ZwURn8YhwnwURrI+mR2TO81fZa2sx18uVuoP
ghdqFbYly81MiESCCZhvvRlZjh1I68WmzezmuNsMRFqjM5rp+ji7r9rFBOipObl9
KbcjVCQbjVaNfq/clHaHJ5fMD5kPUouyrZp0eYQoe0hKkIo4K/v/7Ga9pTt/pnFm
Wdo7e33OHQ3OBVXOxvQG6UTiRZIYd1ieM8Ex3CuELqMJtMSWWO82K27qj1HGQv9t
2UEPsbnvbW/ye0KUIt6wN/NzA504FtWMAMzsOL0LV9JfE0PIKK9KKYviCa8Hxmvk
ws3b+L6IbaE3HjnDWf3/CnwlcCdMjXrbmD3j3yAciaGipzlO0g6NU+NbuNmhaamA
B2vdN68Uj0Yo+7bc6yq956spo9RUwVQyKoLy3lH+2co8s+3JgF/UtKYL17bLPj87
jtSXMnnYwEq42q+vnjPrbc2gxQ4C/SDMpvPlwOHP8h0TiQxiKDfyMvt+3YduHKFj
yS5PkrANCzi0KMY9TJXKidcxU6NNYzT1DBTRITOWnDf79Gs4PLqx7KYVhRVTkahi
tS87VQURKBnpiDsPmvlw3+/Eo4FhY5ZeoQpwp+a+otgPTP/EKFZwvry2tessLNxF
QbEY0RbLWYth0bC7SGrqHUGtG4XyI9p+vf0yRX38nSw6RXROmWgN2QGUhpCEWdIZ
0dAyJhZaFvfXiDJLnAwMcmmR60BfX33yaOqkbmt9ItY8tj1gYCJLVsKdrqz+AyW8
LtJv9+CHoqSTFT3cJ8V6JNYONypPRdQ1k74kCoHdW33RmUfKFM4WzqpKkJfBdgdX
zzuhcVUR54ludlSkC9rwDiNHKCelmLfq1kAdFhGSokZo2zKXq+i825PT684LNcCJ
QzI0hPsH6Rz1nlfMF11oYgvMKtMg04WXouq3K3pzvYol25gPIGfXwAoEvZx3D+wH
DZXvySE+3yAEWw2IRCvVOtDle0j+yLzvlJOzDatkaN1kVrZbTBTmEa9tyX2l253z
LxoZHaV14Wo3pt7WKGnO/QFWC0oxvSoh9kCHdjbvzTPd+SS49a5lYMW8OPknqnKr
g6mznKLjgC587OosQn9K2LGOx2LZRqfSFQHh51z8RHftPoFZYrsRNLtQHX9ehxOA
/PuhDDPkq/ClKz94ihcKbUu0zvpafc9EoVIv2G2V3r9dNhdqJENSeUxLBJx5i0PU
H7pLTl2jtWwfHejnV3Zh9dXc5b/kLEOdsZ+o+O/Bzhz/TBUiGuronMPch5grcX30
2ccBetZaSVYcaWYtsvBSwnh8T1okkDJ7BYeVrxdwO+O/LmcQwThO+ScT/UwXkDzH
DX4hQ76jaDevFAFI+IlgJ7etjkipwpJuv0aonQm6DB3mWeBx4qoBDg37uxZfI2hQ
avcCvaymFv3Iyj7g/a/wFacCUZUppgjWP8QhlOXhPejCWDYXCsqT351vR3aFtQQ4
TITkrcHHSKnLHo1rCka24qKDbSS+ievCEWjqlpE0ixtcrVLTOS5aVhstw6tFcp4i
5Jz9EGU2HX5O8eSqwl5vtO2yNN39JzZbyz1Pt2N6qjWauH8bm0X1cuH70b1TJunZ
VhXDZdHU6DHxXqRk/dzy30Sq1MdU86RG/HSaaMahqL8JmnjUrFE20EyXJ5OumR1c
XsSU3Jn+Og298HueR7HjKIXCOHYpjts2DBEfmllOiuiq/Up+BLTt576V99EurOXS
5eevEXDosJyfnuHBH7IPm/j/DXLB6REDjV6uY44rrjP/iV7Wd9GBNIHL9ECe8Nlu
zdSqWxefuY/MknGOQ8bh0bCgIimyTEbypo95cJk2SkF986eKsAuVRZAhf3EqG/im
uw2BEQhZyVZ++P7Wwq+FFQ4G08vSDYmCBKtoxgUU8pkruZ9M7Ib86XkQ3cNGdMVH
ysbeMZ1XU903BOKa0QBcE67ihKg/8y6gdum7LEnoHmG/PDt0Hgw14y+Wts8pLmf8
YkLaD6cJ+MmAnUaHqswCLdW8FZ4l1lN1W4BIBmE8KL5x9t0iFdBESoG53TxLCabG
Ew4dyPOp3x9E2dT5+7AT/8Ymym4X4lrQdjntneFAHZP2KFZhI1NOT272K6L/0S2d
bMOczirujlCflMkdLmtDUf/OTI00u0BnyngR7QkvWpsPK92CYLH1NXyeVLAjz2Iv
5uOhvd09P+hDxSqpe2H21l40Br7PBgtV20Mj+t3rYoS3u8JEdAIj9CBY0bA+2pb1
UHvLsHXVArxGTiY1gcFpTY9OLzmtCeMpDT2Zouq+PzXgYLyc+xdD5IenMNGwZ+ap
yHTqYdKLgwvSyQuDZpSTcEbzA8kK5e77Pj9ORYq1ncw2qqSSVlAdw2CMMY8wfzwr
2BpJ4NpeSo8tuXHSVVzHheEkomQWDqcuUVq4Egmdto1AsU+iPCVT5ONM3ZkBKIof
NgxMQakDtrMwQWFDbmTm5G3U8LeY8Q6wmBoAkWtPPB0gJJndEDzyF1lsq9a/GixO
Ml2AdVQMA7tlcje2M2FDe/v28cIl4FH5Tti6nqO5cdHQJ2hDgpn0o9XRQ4rdlEUV
YtZRMo8Wi6YElGSLIcsqylqJ1yCvcI282RFUstFYZMwuHOKS1jdKENGLQmydOq3w
uz5oDVcMgwEOspwV/PYVo+l7rjHm73T5/h/ggkjaJdYkId0BauiGZ6QI20fT6Nq6
OTzbyTfQ43vp+rDtxHaQae3je5y9oJbX8XMtvuIVR/WPQfUwSoNYY6kZMEX+GjeH
jO37GwcWQxEdZi4tilvGljKMrbMc0Beg1rGJZKYyIIywoGs6CJtNtY9GYpr2InyW
GDmUobfhGDRhsQ6OGsNgvJIH9JA4gaZ0LK/IF4m4EcH8fDP962ifFl4QLDmycWlt
6KRZjoW0gA/v/+vhI/qnIxL2G3UMzj8DmJrgApOBC3w9nE7lBsj2GKxzWk7Hd9R0
csUPiwzkCOuEQqQqeCCmIDQ4b7HpdhCjQobD5RhoJCs/XY2z5MqW4E3L5w/uhvme
N0u7pkJKeuQpj5FGOmpR50dV3cVsY4C3CNnYg8qEBb46cQZfZ/l950bHmm3IPP0P
j0qemFh0EIEAh/RcwGFA7d3CW/p7nZaIW80jwLkguL9tOTAliAxUK5B/5xQtwAhU
TBZSW0dwHd9J6i9r3M/9VawDDLYW/k6dtGtb5khe5XlrFZFGf96Tvy7bHY3SXxVb
YgnvDCu1uGYyaGowg2GAdFppjAFS71BSWLlrZ2i60ZuAKd6NTT7kl22QFONDbsap
EfklGRZP+NFLpjTnVZ2tDpBexPfPY48BaO4YK+5/Zawc1b+S3IK/BavNT4scEPmp
8gKL7N4Q7bD7lZJzokKp7RlJGl/3UKJ1b40iZFgybTA/QvSfQqCXTN2dOAE8tsJe
bHqZkaoclvkehEdOBbGPbsELGERHcFnceYY0U/QTcIZIsdcS06xNxsQAAWIBT1xF
93PrG5La6z9dHVLfKsYaSCfp2v9zofNhtQdd8KOOI4lfgvoaMkKrIhi7CXvRNoNs
jGjXn5tYSW/lKQichtCgzvjTH2ySehMm7DMBjmEZ0MnVmWN2M/JmP22wlX1KRmu8
aNMlYG7p9Ax8RyhbJV37kBM6WfcK4yuUep0WGCkYkXWOKMlRY1HScGYznoVjV6WV
mga6XYrlI9O57G9cx9jWomOUH/UmQreMNllbBW6TBdoETe8jLshpP+wm7bhOopSr
7Q6vXiZEMxbeo0a4f5jewHbXInpwAGT7ITFbvmFAVxUDZJlGiTEBTaOm6J4zrjsa
2FttPI8iTbHK1OpHz3MhvTTSQLEUYHmihqtY5euyGnD5JzlfPVxAV2gKXgtQHe6S
gumI0DmDsUsv3Y2RCSPgn/MxuD46xq6agKvrLohrP5NVV6a8jx9fmeg638Ojc7u+
KZd8I3BjojQdXjHLM484TX6XC2eZdrP9196wq4uwueh9Ddd5oiTNPNdiAlemo9si
Ubafk7kdJ38EKEkH+9q2d264b2MuNkYE4E0TTjvoQzy6KPYyWzh12rsYmnG1vnNP
te7V1c2tx4ZTSZwsgv6MbLX6xTPHmyEcde8JJxmOuZlQfb+Eq9COPmV7B6n7Lyzd
fjk2+/pNdhyfFZhhHIEigPZamL+14f61dqZ4mY3vIgsqyYLOQtNY4VX5gPudaJHh
0HR4gmXxdXSykggQFhE0lpMOvICuM0H9+fcIX5KGLYefv1KkfskCHGWpISR3XqHi
36S3Kc6HoDHcHvjS7nIXxulN7ljh2k0vz+0ZoabVO9wSSkLI6hvRs2NPkhF8IWeI
mYLDc/YGkC35GCLzzSncXuSAi++dyHqwnhJIpj3sfYJvtKlmurHJ2rkmeQJZtpw+
bPuo7w1oYjdcNdE3SVd/nBG5rSdt8VVB27JcAa2A1X6vgaQXk+EtOtY1pwcnCl8J
4iq+1P846SLWjm8U2SBTMtJWPWGEqRsC77EXVuzGUCqnjPnid7IZgTMKGMx1zrxk
5PHPPxasMcp3BrEl29w6w+HzPS7K7WjfspsS6xVqu1Naq7e9Mk29dEDCljYwN+F+
DH6o/pVZKV7mSVgQFMd0Ro5gJP4VBzg6ufUpyCvDo1DYkY+81m8QmtBPS8VlMI6Y
tmEXVU2EL+F2kOlp509vGe2IGPI5VpdvK26Gpr061yBm5YWjhuYDaFtGISW5eteS
9M8Rd27CLbw2N8fz/YSsB+7yIg3V9V8uRnsfzkeciV4pZGwkHNYBvY+cyEs7vJgO
itiv4svp37NsSD66CD5PBkhx/y2r5ryNr6fU1SIoggxJ8uzHhbVg6VMp/ZmMRv7u
1L8SDkiNte8zkJlkhg3yZJcgNpnyO88MF+IVd1QpjM8Kr4CpNzRCihTEsXm4kEyH
S7v0SnY3W9R9LhHQHS0ydf8O3eCMhMoNdo073a+Ten/KiXYkl2NCacsxlh1lhEQZ
RZS4Qyhrbig/BBX5ZwB00zXPtljbx22gWWjuXumWdpOt2DV1ElTVck6tCPAvR0XP
V7bNBJKOASSYkB63eGcqcKep7vy6X9TS10KhIpD/3Qf6Hq665dVuanUVtPQmFNkQ
I5Z3hMBum7vdL3sK6Ci1V8u0R52pQHhQEJn3SakiYhEMUCc45iRVzZtgCedXOrh3
DR9/nb+xOa5u2k8v04vue3rrm9KO2bLpchu/kwNz1YiPtQWCWmRbHfyh00IEOAsa
pdlPZWyJ8SxWUP2ILV0Sn660Vaci9t3h2s5NILu8qvKW1qT0MGkH+O3als87bzLX
oJv96F+NyJnkxGBKvhCWwIE4ZkSe2MSRzQeAMKYJVhNer9M9MaEAAqO0QlmYo+lB
Dxh3UHXd1gY5XhAZIP4NdAupIan1NkBEYOxZ60T7Z0dTrqoqJtym5o+H3HxEfLRs
dnddpslnjGxvOnYDZleE7yL+uneXyjaILrpKW/A/cbI7C26+bgKHuLScCY8N+n9a
AMIvuN0evijuhbPwieYTQfRcAYzdY418qWrccT7koYj0+O1yXoa8Doeul8UdNUMo
/5USJPG2c+PDEosMFswCtKIzovZ4DKJryRu1jJjh1tfOSl4Yn9uSzmR8r4VQ3Ial
Lz+9Nh0VkOXoF2lG5QEoFufP9mgT2mCfpNHp+6+mUGtWrRoGXtZ137B01XPjVd9l
LHwu5z2zIeH+gKyZdKEjp0VZO9rvsnJQKt3vs5LhYRCJXUUdn4Ja0P3ubgpFR7N/
n5KydGefGrS12zQsuhPncrNn8Igzqh9LTvs2ovjdRec/njV1jMq/9lICmDUBy5lg
0OaANN3ibI+nB5VIewbHztJDOsLVGcryHCqNjbou0pjuWhPLlJMOpH8LKgktpyJj
lEIhXbcF6QYZDEYiwcTJyRgdPpfzI+ybva3wzFPm3ZesU6mFZZ66i0V/upRNSlfB
/cSZEb+FGtRstV5NqYede02JA68lPC0qvjB89I5zJ4Cqx+aMSBMtwLYHUmAu9C5V
WcgxwOMI4iqu6LRIDjwzw5a66s1zxb8yp4PmsMYzmbD5HhKsZRvok62xpQ1uvV+M
lxHaDCizxJqzR1m2GWOWtglo74fYw9O0BWZ5Gfqfz/x4Hx5YbBh+WUyEgwCF8mk7
RbZhlryczdqvYLmc+45QCJ6OUx0ZkVTLYYlQbBLdngt2sUOqwW+Sa3x8lJTwFATa
a/c2IduI/KJxWvVda+wwJYu+ALwl6JkIvrIfnVQT3pAc8g+BFWmX4xsQWPYC5nsd
K8Lj5mNyw42RrjYCIQrpBLAx980kw7hkbjf0Bd8sYhgVRJneE+VE0dxysFlLxoIF
M0BARPiQlZCAKOSvzsjluDNqIkepJsO/zUHywLZYLpM0gZuAzE4vHuih1w4rRwrz
pks6YYoSylI4IURLgT7JKkSvK2aBYhTe2TgdEzMmPuiv5ys3DGp22nGVczCfarNU
wpsAqkRGpmImkFKE7rPIJxz2nAleuv+IYW7QajixbiqjBLqpvUDQiJ1QTN1Y+aAs
/CYYIwvVmrlU6pSR5YIRflTcoBn3nKpEas/dRpOZu62oO2vGCeBKHPn+eABFrGLx
prCCD3m2iYMxme/cEIqxxZbQiVJrXI3unykj0QBQPwUX3JGYeYKe+WuL1aqHOfU9
G2Qgmf+kcOy+MO3/mymCeQm0bjjeUNpK+jku5bLAGGFbIyLZyVO90CkZH90QhQg5
Z4YNVVp4tODIvwc33cn5nrH8rPpGgafgCdoad0bh8oHYpFTFhSCVd3/eOR6FGOJK
9r+q0+X8GFBowPaX9Os1tNtQKBfnFSyTWEwCkeAmZa29ce1ejZJ9nZk8yeEkUrsK
qy/ofci3acV+s+mlt6V4MqOb4Bf1bA1aqoNc7z9458hYhtK2jlNWGVLDPbkLMSLJ
YJvFeMViWGZ6WRgMDXBUrwDz9K1Gx15eHcdPqysO1DHM5lywBPKzEyi27AdUvMNt
/B2qWRYqED+3x5TaNlBBGS4MrCghFA2I0YwGhKg/ntEw8GEQguiGSN3i1/yrb4MW
SzrC7Ih242gSmMuxwJf7m4EG+hfDZq0mTjbvA1RdGma8PSpHjOXMj2vWsRN2rmO8
Tqd5U7cjjFwXPMjUtXZGf2I9TJYI4zB/KchqRFLXS0bUMw3IoFBMb+HCs5myx/6d
EN3ueo7zJx3x4RxYR3Ol4TvBkSXXoLy/z54hKO/nrsL/RGwgaGTHDZhTUBykZhpG
kiL6qDqTA9mck21xjWjiroYDLLcT4rZBWx6soAgtnhHenKegKtxPbLRMBHwmcQxZ
DQHopuv70w0hQOIyZLS8/KgobsySwKYIym36GvWUvnrnpdPyU2gvpa427mI+sCHb
ylcBOO1EYl9z+4eJddmphWVkyHUMRWPUTCgzL1O8y39QFKaLzvrvOSSPNjW1/moG
MXkW3gsRVHN4C8TF5HYUbTxLbQ0irDTGXzJkdM6kvNpar/NeHHte3x4U6kDI5+eP
T56ydsaP6ezbMKsnHeBmzthJY3cdSYOx7NTcQrllo3lxB8ceP2UEFe5rlHAdn2kk
NVemRkiVyUEs9QXCvlj4qxgN32RS5JHUKppiryKD6TbqPDk2jgr6slgl0+A5st6v
4x6Ssutkt41QJMkt72KjLksq53sbYpa02HHX6khnSd4dZeowiYP4sSWFA8mu1UIq
AxHhAb7EWmUJwoA07DkO9hK8NbN3sICdFH7ArAzwOVcZ7gZMSKaFY0nb8UjKGzy6
jkXLXm4iVwQ7N/zjeofX7EJYUSqYLc8Rw3XwXbzvx4qE+24N3GVOs7F5SqIm36MF
JCjeRd3WavcdTQ2b0aL0SxwShE95VfJhyeCM5clzje58MuQRKbwmSLDxROpNdrAk
L8Eqou9tbBRL8FErhWLFl1GrJ3U3S0Y5HE/cpJNsQr40Ch7Zgj4FaqUq4xXeY269
DqtoH7YB24OEBb50OtxTDzkOcwWt6VBwfOqZ7ojTX/+xXuHUE1NWbhHMIejZFwyG
NLEaLIM0DO+QcVW4ESBXRKkz9w+R1mX/SbjUFKTWGYLByIkHdejFJBl9X1tPI0Cu
IAmonAl2LTOT8qI9aHbZBYzrZsjL6k9ztcR3o9SXeUJgPcTPeG/4Wp+1tDg9YmGM
D4KeHR8NSnMxjJ8RRqBATGxwFeFCcTeX5yoCkOFtaUhjwJ6YwUcg9NphMyoCNAjt
R5xd+KuLP46TQ7noyVZ+zzdnIN6oDqo3EB7uSAlUYKTQXgEe4+JX+8IHCk0st9p6
L0gP4ChcrpGHJ9VCSjqjhj2xMDO3nALn79G3kaFg0sdltAFANEAKkR9UmtQHHVpm
NTV6jLugdahtNB9DwOhh3Tj3jrSZWz+TQx9YG9lMbyXD20yx2x98MiLH86CuFG25
S5AdKP4uDGBWp2meh9WLqGVwO4f4cF6SWyZDMV/F87XEbNVle/5fA3qSzJ6/YIl/
ecq122Bdcl5TF0J/y+Fgz/hx54pwJlJfS7RMNPvJ3p9qT5lRqLZKXlQkDRFEBakR
SxN/33xfpoy/SGaNGo1aI0ybIXFOejqxdSdPEi2MmL2imfL1+viADHWmmG6fQZUW
6GZ2u1g2xHex8+wukY15EluqXobgdst8USCPZcIzo5CvOR8x6FLN3qmJWAqcPwTa
1k928fb1i3I6x+HmuwhkBt0IStjr3ACMDNBZYDwN4eXlZwsBLqGIpg+KLY1J7jcz
DS1daCGc+8N0ShkJ2W7cDG2FaiaQAGRXmQqTKVUXNudfnalibEoBqj4g04irrQgI
Qn1ZnWWAmUijGn3owFri5kOnfWF9TySKWyRHNJHGQyGTGiitUglbn41F5VEUsybH
c4Wqr1CJ7YkbWx4knrcBvb+n1p4BpiJLILsc3NGJsalcCRS5hpQ8oVX54vV0XJMu
Nf9ksrUov5bN1pzwzTZIcPXUqWftGYS6QR/SlpCik0G9k22oNkjHXwyTB6ypCtig
D7A2za7o+8MrBe/PfJy/ihgpoxiruouX7pcL2Mot4f7L8jNIVwyHLEl8vYBzf3tZ
e82e0rL0Ch9AkWtyrs66Qm9O6dvjmm9C5PTGjAiVuD1b4VeOKASY+sbgKp2ew9xC
wjh2IBqZgbWx7msFfcnZ+9oHnEasUSc+/ESc4e2qNYJw8Lh2vhwywHz6VRwwNPtS
AegWet2PPd8/EGKLN1HDh/dP6j2Xn/tbWROhROSnBNHhSO+myYXMgbGZ5rXH8rL7
Krilc2MjTzDdWQa5GRvHKzqoRxipPIVIpfBBK9ciYLaCCD82RjAQljdX/KcD/Jim
/94bj3JJnbZ1Mdbi7gHw28xeoCs2LzMDNP9t1OKCj9Obx2ztHEbzQQllr7m7pBkm
8g4GwtvVIyfWYWW3/9oXfY9PL99WreT5m8WkW10FRCtk/C+qhhhOI02EDeG7DOFh
Bz9l9ZanpEldUaVVYAxz4Ttield8ysaitzT1ztF5nIFC2TyTJsnWXZa0j7BWZRGh
8O2+WoJ+0ZaUQ73NC+2doOWWPPBRxGYEgqn8U3/RvV71LE8mPnIKCmTHSTEGVuSS
CgOKTeoWJK26CWdJ77ZyPu0ErW44QiPOLzP9qpAGxk7Yjfnw3Kx16wtueRN9C2YM
Ewnl1IqUsLCjwAMZQymxb8t28/FjrIaQIV/38uNAtsgQwxz4Mn6zvGUBHa2IlVLR
UfNAdtYjdusbdma4pJvQByp4XAz/gwZ5P+BLtTz/zumW4qEU7yAkZBCjfVztw6+z
nQ1Hk4+1xZl2iIZZ7h/miEkr4mIyxcub03bB5o+ugFyOFm6sXdafe6diSDMalK36
idjzeAmI05dNHfW0kiQqGFWlqqEM9Svuo8a1QrldSfdddQ4CjJvo4O9HAQWza8HX
jA/0fLCCi0OTlWYjwtWb9+vMa/sKs5qPkIIVgNk9QuNPPoLau3iKsmFXqGukMf/N
pzxu3VtbBTDmrL+T9UMRo40fc6KbO4Z6BI5j7XnaeElaiCVZ9cDKZhcuBaRTfJkC
JnauApg0iDKe6FetdJT6VOrREN8C3n63xonbSxcHexhWhd/fG7XRrJlADTS4abZK
A0eJ93ygoFAE2532H54WsnFXHAiX4kRqJK+5+kA/LHDJ7J0usamPRb9dCARgVGwr
813VMkpVsQsc4sHzIyZjL2JaT47J9jbweqdzvvntMNnWzkZFitJxnDUn/OD+yRFm
oNu6Jse3GwDBFhfmHqe4CsBs9IivNxlMtoRcVVeQDImRjfxO+7vXxysk+O0O+ds4
TbN10bV+IuL0p87/TvBgWn7GeDOQK1bypzNdVMav/p3X94r0uomvjqtn6yAW8ccR
17xdoYWFaCNbQmKH6dATXEA4gCkuf0GBPcHKKYjtigBpODH9Wsh135ZrNkWbDAMP
fuKrE9yWP8BZzQHVt2Dy//0/QRREzSYBGekcZaIlaoX04FI4rNAN80INBtiG92U0
BO6Dyy7d+63+BfqaeKmGpD5EW7YfPbeTLgnVtzAGaNtpDmRcrA6yW2hmus9oDq9h
Lj5rLy3IX3F0d0pWnsjAbS/d0Q9hyzTA2AiErYXTF60uBgKZ8pN4sIOF1fIQZEvG
DjvKILMTMA9cg0wkoIUkQxfssFedCx8hUOaX4S0WFDKUIl7C8RMksNfGP9GDbxl5
5lt9grePuIPKyd7sJzzo5u8PNIAbpuBRz8AayFV7BvgtjQN5vkeMaqlI8/gGfNe0
Y/7kLoOplNV2ZpIHmPK45tyTYsEQCNaORNjgGjMmdOu4FRTzelPR08jSyvpKPDNY
Fsxvuj9qvMMVvS+KMRzLbm2vaLa5QiUBT9qnHodxMjOZXmHn8NUrmHS28QCLLYhM
kdhCI6h/kXrX4WUxSW0kLhIiI5EEfF/QpBWt+KZhkZyvBWYafFZ9xI1+La7VcNEQ
yP2AC+fASxpNqJmGXE/AqGe2WoM3QVE1ZShHdSI6ubKnOeH8Su4IojgIHoTBhRMe
cKetCsTHHoJ9rNNPixdAOAYsaXavh5gh9VJ4Ge2hLD/n9bcV2nElQyvIeurNiyHd
/KVcrr/mCj+koRnImpOQ7mJ8yfTiUuc4max6SkJ9X+m/ufy4bZiZDK1Dwook11JV
S/jJQbwl5QHvvlgg0cQ9yHqcPiXf98W7FGDIUwe4yQXxijFUV+1SX4QwHMWt/ltX
1tpipKCn1lBBPzWdhNGQtYSVjYcfU/l2KoOs19mvSVqq/Z3zBF9h7TAMPdlmx69O
lYjGZ0ZAMhamdg65zfwnHftQMBlArDQ1QR4ueZ2E7ayQ2LGCq610jhyeNIXwymQX
Em7Xb20Kqrb/m5JmzzGkFBVNTiPg+/Fe3R7r3da5fnQ1YUkbFRIu9mm/DUcBNqo3
I1Uy1wCcgnCOSWZ7m7q51FMKcfK24aYmzlLpveryenHPqF5rlYbU5ahNVjJ09DSc
vaQ2GqJS8ndbIp+z391VpelUfOCw7GKtinY8YZ0+Q8lDOK3ZgWe/rCUVNl21SttR
CeG8++rpDY71ZgfLxv/c4ylZ5loGmTzQndMmTeCrskinhNLba5gnh//ImUz9ffXr
TAQ6/fO1+G3EAHPCJtMSkq0K6eqCCbTwdSzM/Z6vv18bmKNmCSH0MROTQOqCLq8U
0cvjoNqp75cfrA1k4vECHavNfnNjZnz1m+g2cbPA+gCtrMcDrBJDip1Q+wx0aMB3
NgGprv5a6ScI3ZNJV5N3NWOHVeThwV6784P/Xs4cmMOb++89Mk8R0OO/xTwPIqyf
symY+6bdvPwJ+NrBijtTttxa7WaHvBTMmkOVcEX4DGzI01jR3EFIdRPGRE3ze4mF
nsbBJ/pGOV50C72Zekixb4SYp/LifzwzGfOPrAPV5DtoKv8JRlFcA6EsHDc40lTC
tzrrEnzGyUELYa82YZj6OxYeUWsG4yPvnq8RvcRHTmQigBnNdca6Uvx4lJrm9xKw
jQ+gxrLUA5eMoM8+3E0w4MgZd2MuNzSQZXR0cNuQOwG6lNLGkqf0TTojerfUXTH7
08Z7eX9sRsVlY+iYFJZoQ78duJ3dKYCYgsiYFDjfqcMg7UojZwody1GTKTMIjBB5
qJQpSr/B06B+kP8SAB2PXqYa3wP6eEVqbhVg6Rx9SpTcFG9yYLSfavdoJt2Ky1CE
e+6xrDQbY4YKp4O8NSdcu83wlFvUvtMhyYygIi4os2JOfhB/fu0oLhpENNno5DQr
Vm/9P2p4YVKZ+ETv0ss+q+L59wRJM+bLBOqtLynMUV2jf6xl++365qlT9tlUp3mx
wVSh/nuMO/vS/1Mgmg3SZIPWmIWbnMxn3egeg1AMUdW0bUXAybaS88qv6Z9zTNG5
CPdVraeTj1usL+St0eNA1sgzzRo+tnlRiCdcrvevLxsjLeqXj8SD95H2N222O/AE
o8euNAiLcYYVb5OGE/3ovIROAyyeGPI8yJLDp5BLP8Fn8Lrskbm5gODaf98QpH2b
7c6dHnPOakgAIweVitt1EVvvtDy9DDBa/eeUYqDMwQ7Q8HjsUeaNWCOcEs4hlRPd
9fkySxfFXCLS2RNdJvkyp4wyi9P5qtJDvTIJtY7usqSY7cqMzcKJb+pj7JxaJgPO
3xAPQlUG5Rezs7RHlglv9C0ZJX53hurQELi1gfKTUQI6CcXwHnJn8BHclF8ITY0a
/DW1w9LFpQRgGdBVL/Wh77bfboTnRKx1wOzzR3ypndAV8+6IsP63o1wGtfo02pAv
8j5XpeeiPr/5PbtAVNmryvC9ULp0IgzTBsxuw4DGwUGuvCWl4AJ51QpYrUe2SbFH
B1vLbi5sKn6ZVCjsxy7W0SpnjvpZPKLHGJ9xC27e9DsGOWmGLAmRxqis/hhZyjuJ
V444hNKi/WrYpuDqLjqSR2bdu+s0HVYBt9XaWEX73q1Wh0qw0fGxjLITd56k1w2P
j5dANm8I0d/p9aEq6iUbUuLSU1MI3V69+JMxgXJYeP5A9aWZAm+ucSYqTOoxTyj1
ALgl6wmW56Iz8GV7HAYcEs1W6jDDDjs6VsnW1GejlJN3ux1WiR1ZebV/wuQQ6LBW
FUwzfG/EyFJahCn3Tpoer+T8S0c+5tSOciGUdHPxBEZweMoN76jfnp+M8fQCmXhA
Z9+vi4iUjY+gkP231NYhryQMGYzv014GPM1D1gQoyJz0a8SjMv2BWzenOrQJUJEk
19//8FwAlH/xYn3zXZR7KLj0oujqogylO2kApxW/x8ZnpYbDhk46+wTXpCmU/V3y
KSZfdedxKq/sdoWL6M41Ma9HQWhKE8CmE9k50w4a4mVCe7weTRJudM4yoxjgWeUW
5+glffhhnnuz1W6glLJaoALGSoyCmr7SpOrWjlhbguUGr0skfrF636PCHvT9kN4W
kqflx1RM0LBifkj02tVpfcxcz9Y313tAu8ARkHeGGesU6SjZkqk+71Gtd23nLYhO
/UaUHYi3wzHGLLoAstPo5PvIo6aBS2O+fKNxjjuVoiLIUktqgA6LOShyHHaFddKI
HvG1IltmJWHpecMy6cTiWV/yyaHAybJ79AwjfFtA6egAZ5b5vpC+d31aRq/dtal9
SY3c+qa/L5t0MaRzzL0A0cB9XgTPZzUpKTarmWReqGb0RwrDvBMxOeMQGHsziGe0
IKLi4NbxYsQE4wAZA/w+BBK7wJMrRLexppxdHw6bZQP68ZIi2c79xd0buj3FHo1s
WTouu5QXMlY4UPpKqS7nvtOW/mSlEc6wAQLCBKkTsvoP0hVxX/69WKPAiJTr7/Wt
DK5oibJK4/yDJjDnDffU2b1kiVUAJf7nr/9YaixV6MgZcBNOtRXuSbTAIu93XP6a
Cqftc25wqzItdzEn/cxf/Zx3NWh96j+C6XIDMFqwfAGTsvChYCEQV45XNfIDa/UT
NmkTwAVKEwh3I7DcrjwJFYszkqtX5vdb3EQ7UFP14nNDWw58zjg4peEAJNzPRe4B
k0co1t7zOHk6oOAEeDgR3eaNsEOZrHKaSWO6AEEJEYFuGVf4mc8oa3Gsv408UwBC
vCkLGISBtvbBik6nRBgEuSkO1q6sNWZND8lrUEuPfx+auKPywAkUa/VYY8yxyIK5
67IhDQgAGv+FZ4YkeRZDtfD2zYDQD/dx4lk+MzUNmgaUikQDdRsLM0tgha9sjfsP
FuCWUwGWkXm9lZ9xshl9oFAFc6s4h8g5nNIuS7T1/tQJx0StPo3L784QfhdfQ7qq
fLDd3KB0I18RO3fU+1ptiIXdelxaeERu9cyduogIVtck7AdF0rQMQ1Tkv7lEFDyg
fZl533yXgGWmoTQI5UJ7dwod08hv5cwMS9aaBbiypOVHEPhOODICmmf3BAxlQSSA
Om0JitQBzo65l6va3ofIWmWW4+n/7bjxRM+0R4jXhD/qFGlIupVuiHPGz0tQQUEd
FKgDLl74WiqxCPdjvCrtjNIAQzh4ojsjYtx10rqK+DbpzNkQWomF/4YOvuzV7Iv7
XDP3yMu9Blo1XTKY4HjFpIbCVu/+oQOD/EE/XlEnxUXGeM24fqTlRblYU7/0Srts
ZZ8n7kHA0Ip/3bQvWIZQ1ifEw8GEtsjEg1z8O9air/x6m3K5NkfjkcdMQ/xsCOqE
OzL5E5bYqtpUapWQV0dr+yBGtMn5qJ5OMiW/mcOAsmttba/0Cje9OQBv9d8OX7Ch
11puRyHOnncGer/EVKE9iPLVdkOxahEMrg7lx4ibj+VFCiD66+WWL8mjqlznjQ5y
XTqxB+jCznq/4gMDPvITcWxgg+hfq6AVYM9N3GGQF0tT4XT/cwqfUQzECqg4brSg
O8x/3Gc5DOUpK4kfZ13HGp86axF6aUjPSwQgNHBilTjw2bxyx22nl6jG7/3CWJ5B
tBIzrmWmFUI83vbX7l6k/OHEiriNBeudXUu9l98Hs1vffUYIIzUtE+MGDWyW/Fsu
XOX0EdIHpRPFoZJtdcxVEJUp1NnIPOTc24m0vUOOtwyvMUXZjpi8acmm1U43JPhH
dk+cNQyKJtl1rn7bfplo0F8nLQZvxyaMmtfHpe0qG/tMxpUS1NVYYXQCBcbYObuE
cRJds9VIj5XqoGBJKqmUT4BoX/XW3W4LqcNjMcjTM//WU3HPk8HW+0e2rOxbAE6X
3ymYBqHmuSwuufBIMT2vX7i8lio1Sz+ZFrRVdNVApxclO9TZFTBr5VfSlA8rJdVa
QzJbyC2vbl/JD1FicDupGgjTLfPrZNGAHwYy2VwPf6sUbt2HZYSaTR5xfGuSz6id
fA+uPRLtJnXvp1jgg5vsmWv8K0tpLLUhUmwBK9RORSQjPXCXBcX5Dtz6dLt8I5yW
RoIa99p1XiS49ocrPRxsQbLpL/cpx2iE968iYcZODTcQkp/dIjFPPU0HBtScbvYQ
0wyp/CYep0Z4W1RH6UIOE7xhqn7a0iR2Qf5ZanaR5IIVW1j3kL1PCADNrTQL9xRm
65vAK7M0JmQL9EBLQjYW6MyDLj7AKNDvMl5xPxyi3gtpLYG6kyn5meULVQxz2BsN
yoqKZ6N2QYf/WW8hFHog/LM5lDC1hfWDxMZRDcxJ1yLmaP5zbx3100hX7ocydz04
3XIu/hxiptOIs1SPx4akB7AIMc8W1BkEkCW5NALVJKjvLvkiA5USD8eYSZYdZ9hY
sUORlTwrde/5N/rgnGquEGcqSeztu3amAFgIJ1LJvL+6JThDnCOqtYWlpTV6CqZQ
0DE36hUnrcrDXD4L017jzPpwabVUIfA9wJOH1OacmhyD+icuVR9u6IQ/BzNKCfwS
7MSFxgEeDrvEoJIlSVSgnU8CWmxkZzR2tScQyjB+53uqbDilmX+elx4X/R7p+Pj8
/1i+grQ7xYsSl/oMydKL0/8x5gUJyyYZsNlCC5LbHebWyq5lIc0RBzlRwqs+nZIq
pmJOwcVNQnGdmS2MkZ0jt8xiaywciRPCK/2LKnOPZrYhjg6+6C5jgXiIDI0eEbd9
I1rGEaj7WTj1BduN8AujfX2YIY6NxkglUjhgFC50YNOR2sFRfTz3jJ4Ru2UChA/x
EE6imjiXOMpHz/V/PhJZV0VBlaYvp+mV25f3zAQCzHPutckTyyHel4VHu2G/qcf7
mflo7aGMPCkXALodh63dT6RIvdJeWbiLEQqn2nycWyD6tUKomu5LgEhFKPbVFcOz
vkJDWjlPG7FK61xmrEwI+PjXnPIzeGGhRWnr2wZ4Lnb1FumqDT87NdRm5n4knb/T
FaKlWX9R1Mtenhkugv/xNfQybs2P1OD/o6EGH9Jftx0S8KkupkR4iBiIbDStE79N
VneTu6eiHwnlU+nZDDmnBpy5yUnQceoJLcnbNnVm5AoJ/Dq2r7Av7cLQl1Dp/Gz7
ZLLvfiDYjZ6c71GZNhln5WPc15MAHilNpWVQ0TS9pwf/0zQSC1drndDd5m8zUI+5
SETiIGINEDeaNtlbt1APOEkzV+UOGeNgFw1Jovo1MYVUSa6Wg/Ol2it03TA2E1Li
RVlSIIEBjh3TPkjDBbPQgHV/rjVQ2xqxx1sMQ6XXWwLEuIiIkZL2pKHrbwnpmbyx
u1bfoodzCAyFx/MM/0hWTssB4VG0t39hgxxgM0odyslK12fvodOYHFDh29yH1Jx0
Dk2+eFDLng+MjOvs3HDKDXxJFKdqxwPove41GIKRkf6XsLcwzRkan0U/8DQfXPUc
gwonlHD/Isw697Db+5+hUVy+pnCyq5ctwnIAqEeYszRXSAUVwExT2P7kEi+V8Xe3
0ZRLxTbI4tSoQsmQ5v3BHvbzvb7p6hObVTKtRDz7rgw2brcDtv1TU8x5pi3qkZUZ
z/rr0ggefuwyX81O5jnCnJXw9hBeXP3j7lzXyURHa/iD6Jgk93lCi5IGwSlDAU3y
nlUqu+wrjVE1MgNndikXzEeAa3SLKOZ3Xr3ZJ7UDrbEkTALAtoIR4k1Lm61sUiMR
dhxjoZ6Nd5CLgK0Q/F9u1F26jE1VTWYIZ7U2s86Fq/wur3uII5vulgyAs7GGMdLC
3ZVY+VrSCG14a8r9GEs3sfFadVsla/MneDWH5jGhn4E1cuJbvmfjQT96ZhBwhOQX
1DpDB1EnxFK8RHSf9NKIhhRQlP5SaGMYbNKsNwGt/X+g7weAk1eXsxc01k8D14HZ
ZV9ZLFN6GAHaO/VPKsQuS9HzPhSsZmMa8cEPAdpLr5Kr85ku5HJWs3CiejKTfsTf
2AyF5iQO8gOotln0nFUuYcfsCugwHYy1wi8474zxaoiNF39jAEk0UPdjo8aS4Ctm
v3pmiOE8yi1Xn0j/7ePkOFgaUPHBTdWo6do159x9qtFWQjSpU0cpftGbIzR/+E4a
77+HckqnhTbwcC5+WKcWbJa4USuFpRvYkMbKkitPiyhQ8sGbyW++hdhoQsoE8V5S
HwM00aHK1XsMZZ8S3AkFrct5Alu5WMoxpSYXiA3gGeMDgWLL7FKd5yxUd6gOm6WL
ZmF8j3DAE/J6c82JI2RmZOitgDbOl6n93ogaJChw1d0ssXuyORB6CbG7dGyNum58
RsHM067iEhJL+xoxBI6I97O/QplpynWoKgIEWpRdpLbERX8Oju/O7tjrqR1GPxfF
1Y8kh8BgjTYHVJslr5QzJTPrvCI0VT1la3Gz1acc6KSnjTG+WmaP9uG4+B0ImJNK
e8VF4CFQjsLTSvN0sv18uWnQD/mUucZBWHQWm0kP8IpviSLP/Fz7aZFH16tswg8Z
piU+erCSVY3NPBpoM5xMmJxktnRacWUfe/xDbLQTno9nPIB91EvqUd1S8xBroNww
x8aZqNMfeC6bfS1Xm4ZudEw0+0ZBB7mAnL7ucHPM60gG+Jfa9j27xNZRi3uBasKW
RcFlQntWbnTr7JhxNed/tqIAMb2x2ICEyKm4KoPcqHCPsaYSGtiVxqnCpG5GY6j4
82e15cKPd5Pkl3+VSBQZU0Ua0Xa7tF/8BKahwzQx+1RI5EalzDqsv+YSwkt5JCI4
8xxCrmFPPHhlIgvvV1Sc3GxDaCZk3p9fhXFpja+uuVExQrexwvimsxRTcTWRKCkT
6b8TpcCvHG3BWejVrAxhFo+wC8o/BqPsQFWPYDxqYVDYA85kBQNsJsOauB8TllCG
VeP9yBCg3kmoTeBKV+6sqZohsTir4hMJ0kqVUE45VRX+J/inclkvydbzoeswBRHN
ST0ah7sVt8LlKPe59G692TSwKB3GzIDvU55Wmc6dLZrxN6KkU/b4nLul8pZT24FC
sulLvxgP1yJVjt8a3QDiXEXJbHBvLV7/GKrLw7a4lvOMdqhLJMGG8DV6dIFuE/G0
cjTIxGbbNDrXmitEyK2+OtDVuDjd9ZiYJ8IxvjY6OKYf0zhlKq7JTFgByuQu8GPs
Z0HaRm/EiL0N+ICfEKXFWV3HCKj6wFlLboYUOJ3AlXwY91hurw0+3U7HKXxP5drz
ATL8QwaWGP83fTxkM+6dQ5XWtsp0I8VKGGPC6+oCtGERtFgSAa4l43XywIRvfFgf
wctJfYliluppoiewsYxcdJhLcgpa5JmUUxnG3/+0aE/De09cgx+P4UenCch7H6VQ
M1m6SA69br9pLwySr98Ki8HC+wq/fh1rauQL0oDK6dP+/Pqh8lOs9rnqbtXsCgqB
zq/R5JFAvEY9161o+vPXaYEFIulpCTIKINLZHQsmh6K3fZT/h6cMhXURRCyFCXxd
lUeB2ZwMCHqGNFGNlb5bfxEO3zWgBik+tBhk/oLXLzrDDZfUUGiWoXGT2xzgvws/
Oz0iwP0D3EP81DwNBps6sYY8iPM23G/WZo0dp+stskPpRbKEviuLZ6zm8GBp9nBf
jfSkT/odkV98CLMCpQ3FQ8OgMhWn+ENgEzdaxgubG2/AYVU8iFSkokvxv+SHFx4e
C0xe2fzhqfVf87Lxbh8uU1bNYL/JvUxMEtXNqZe6iUsXNXivps1dpBW4UbYaT5o0
3EVZAYViZ79bs+mSwjcAm6ZPH00KNbxKIQgdfi739e0xFK0RMhnCS9EMRuIWCAg0
8ehqEybt/iUFYHNiC5F7t/G+j3eMcuW8o3EBQakRR4y6sPp6IKWczgmeKfOYnXV9
nbzYIyB3r06MHjLcLuSyIMabRnUmGSJSXo46YF4SpIlVYdFrX61peBHiGaO3kvP4
e6DtnMTUNBsJenqaVzH3o/qD01fx9D6WXADKpFCAIEEF7oog+JBpjeLa69Rq0hal
p/X0aUM/9yR8FS6lIazto96sdKVY1KRagxgo/SQ56HXS0BTXFq78xHW3COPJGxgE
HoRq9oJMBU4iYIC/tQhmHpiASsDWzDuO65wbWoOaWKvXfAJwctEJsGKknH6TMEMS
7/DYcGG+M7HU8/Ny2IuYslHVt74w7JircdJzsrbHWMidtnU5/dEzk4tfP6nkMmbK
KAon/BMnUthiC9zSvbfUNU9+V0LxV0YON3IwXh8GP7t9wrjuDxrjSuJ1J9Ys7HwJ
PQE/x6nvGdTHLGmSuWPNGnheNQ3lZk1GRQyPK865ha35C5R0WAepij6/eZWr1ZDA
Q3DudcgNcTkuxisCUjasHQE3J9aazrNlKCqHDD8hzHpXaI673Pt5QLNS/V08U2a2
tmnEXmTJfeKfANtwLXJolE5CGYTIvDgTk+J+HEX5zXbE/o6m4ZeXrCJ9iEvliFmW
Vt9WqpDjV3aZEKKq+GebzOEpdwc6A1OnPBekl4rD/WBazo0tUHugQB48lzVfeYFG
zPiNArj3rVCDmkwXHu+sEPSwHpLwR7eb+Xtx1ftXe2rWJg5r6kqXAg3pDEsJIZ6t
6sCtzH7+S2PNGs2henoJNwCeto3E6YyCeNJUroZXzXTtyUJEtfzaLyfraI7mEJDu
+PtTDb+iKOML86qN75D2gbH1hQUj1ffoBjhU6evsowhQkoj8fXXk8dZAMCae7TKP
trJ3kyZl+9APEyKzFp42RLx8f/uXMzY2xynC+FbUFSbRDRrIJCrbnFtd+bMnKZAS
hcowCE9ddhIbvIieL3sbmmwIn/rCypzKjuJC15OtyMsc5wEdnM43suaXahze1f0D
70vxRGoDlHjiGxqvKV/3ycy+UQXaYyCN1IQfOavj9Q70MBmNtOSeDFrLfygb4mA4
e8oMKTyG2wMl/M2zt+1422wUCSdi4YNwqLSQB3HA9SdyuQ/GbucRB5DLk5157t0y
3m7IM0K7G8mjra3f7uUKLOgOOqNOtAP4K3RhLoJieKI3VUNg+DjfEMKQ/HvDjpGv
61Ivui+COct+SJMLMptlpQstFWoOMl31rbgfChfXeA7+pC76xLv+xcX2230zf0Wh
xZzhoHT1KoIHQ/DRW1ODsWQT/lRDmE9gM/ztErY1xVHNqdeDs/qHj840FPkjzNIx
PUWJH+tZZ7JrmEPtqpty6hJhKAPdt36Zv0X206QzdvOVustyetbPQM4J/wSpcZWu
wgSWVVL2btVIzxqlsdfASc5NKM+ArfrsNsleWUPG+9VYYEl3slbqHUh5Or+IfdI/
9Eh9bBIC4Qsw0yY4SMSjo76rPIaImfWu4g/JpcFjQXXNx4kyZ5kgfZF3Idfqk0Jo
a1CbAxYXFrGQioKfFEseHUhSRIGEmzGL6RtDkXVlzGAz73SxnxdiDE1hYJlZApms
QNrzWu3EgG+EnAGnWcJmTyLvw0JpmaEUhabqqR0NWX+F8LBqYZZVogKezj+/Ldz0
UC2DE/42xcyok/fckWJo2zC07xRkbXNGDrtoNQXZN0vIGf+aXqQszfTtwWA/UtNq
4XV9XgwDv5lwl4Ft1SGmKUjvKXFjYHrGmWYfLAeGNbuYmT0Fd1XoSrMTWEz+8fnj
lLafcVz3Cg0sQvcSyzK7OHYPEfiM7hJ6ZEFKgvFu/5aVV8Xadh/xRBmBr6k02EkG
S6bs/z92CBh7Q+Al4dk7XIID8OS9WBjc7I8miQGPVTccSg5/JQsJpOzCb8Q22zpk
wMcRoECtsSK7pMKrzG9+1pRSTYLkMSMUNWhKvZN+ljuubcjO6PXbKrvze2QE5TqI
fxmWwmXqj1lGtiH4YkgZxhWUFjsZ4+wUtDMMhLOfZISIXb2imGCHzzNAveXMfqk+
nrfjTA0RxfZYD6h7N20yUSc9Tf7hyujBa1Hpt6r+JBaC/DmOAo6/xcmVKTlKH4xZ
ORQcE+yTRsQhl9lMgQnQtFZZ7YBDci0APJD2aDmcAq0CmNUYP4nlw+Z5Qu2UGeda
WU9N9lew/UP8yt4Q5E4sfrlzHqwickPmsrUwM1IjJpydkicOhYFC3+2XY2RWtxOT
C3c0vFGxhRQM3J+N9N1nioZUWHE+bbm0RGLWT2qLHwpGBQ0rkAm0EKOkjqL/nZns
n5HeP1jJbZXfEiCJkaJGf9HTTWYA2L/bxlngC9k0AN/oAS2LCgp194xjCJ4OA+VC
JGkdKu+3Gx4aVfBWUFRxZuVRKHmDRNIYVBnx6n49ttTwiMN0ohRYmNUJHyA7ux8x
69OtPhgS21c3sRkKR4ReZYwK8fQdkxlzaBRDuGmwilL0j7wJRGCupYAskwX/93S0
gfdoorkF1vpJMMBBN7TmOMK9Glyq1ped6Z/5tLqLrgO/bW9UR4QDABmDdasIw75A
BSlil3e4XO+cG1ga5OXzgnLXrO2ixqgeGF5SyHoBO5+ThnN5x0jkF+6d9g+WAlOY
GR2OO7gJjac8bUw+SgOuWWqSFiZJVbBb+yVHAdB426nTdqHN0Kpt1v7vrss2TNvf
1KoZSUf2jJpNPCNUg8WxMhDcxYeT5jA4e35I3t8pu39efczaZ51ZvnN+BpJHz3Rj
whgtkRdRkgH0fXT1LUOQYB7IB7/gm7Mf5P/RACt4brE5qC5si/VxMl19KQ7k7kqh
FbCFtxchQP2JUJkPGy7SAeB5PVy2DGg4IsWCQVrZ1FM7nfrbVTcIqWZROqJDjGmu
dwArUyRl7EgQ4OnPOnuHO+toZ2+b8Y8By0WE9ntG+CeF4ulE8rpWotZ620bVi/Yb
2K4XoGx8AkKCpuY9T9BL5PJbDnRF3Cu3KI4qEyQZUF+PhDc0JIjB3EGB7+w7TJ5s
AiQEtXtm3nS0gSrB5TgX0kVHB4wIHGXSL3PaEjZrR6FuGdbsxWwvpctRimDtVTPg
pmHQVMCjAtblHba4VL9wRTBhxCnhPaqQsP9gc7ihWDvpG3IcdJS4QYgb13sZWBNg
bxT82yqxQkdjVCUH9AXKOv75Ehl54QEth0ivu1yg+5TdaZk9C9VbF7DM8+SfmLRN
tvtznH4LOlKGK1Q15i97W33/MCsRVP4g4YNbltx+e0axZ5PXjPvp8BSQVLTu1sd2
GpKC3x4AReeQofAiHM0Yeg/gW9izfdFAXPHpCG1kqo1kHQci+kPeb/B7sH6jtQas
HaO1usXEgUqd3inJAD015FM5D4VVc1S/1dcZIlTKMrr/pIXEDT1V3CCHFf54Y2mz
h+EMq6qz0jw3HW6KieTyXAVeCES5p6atzJW4WAQiV5n6mAsdLmI1vHqh03BjVHW6
OkNMuHprPnJWhapHJUPO82yjsmiUFYy/5xzRipS3ubL+434pgowVxngzm8eAyB3U
066EyYFKBhqGAw9Ky3ExrqeB7WPPbQQ8F2DB5GMuU/j6MK0/jL+4H0WoLMUz/PA1
etXO6eMvDTAZsh8IsNGJoD/dddwFRpxckjPOyZC1lKUTJwSeP5BT+ji4HE469vPN
G88qTxB6ixIv3oeS9kUcGU+PuR7IOBxESlDnSwPDyP51txsJMlWhEgLZXm5gcI5v
FRr9h407+RlkplHZ+ZPFjdfnIEgl4SLKQGTsYYWZbmBNWiWbxiy0GihYkeYHsWTC
PP/5tq4BEqXApuQSqk2mntip23+8qBZ+f3Mhx5HXypzn1t3PBGzol3V7I21C/Uj7
LQesfuQlJnmPzCBZypHyez0qhjtd9qd9BuExS6gksnUxAfDU5l+BXdSgAVLHvMCG
0RDqkhFxIXLACUZvrU10+DcymulM9t2WzcIb4m0wqQEDgYnEUSfUERc+79M5XJpO
1HwwqYrqX/lsqXJKL/xWlTKGY8uF4+jZEHIQRnE1O0izMEtfyOce3zJRuNYjc6ML
KOl4KKyG6qeBwmWhbWW0PCmS8beRngBLGsen26CL8JMYrp1X80UEBovU/ylB6jVW
Sf0m4G/PfHaRAM3o5Cp/hiXwgpjFTfbqZaNeE7C0y00DbvPTcePo1kwYycgPe8In
3Pk6gkgpUlctf0ZaCfgTwD+7xqgr8gYoxMTjDyBjm8aBtZ6MvVPaJgQNQRa9fBgN
KifzlyqES6Ct1QdqyW3cnZUetkXJoHrQNdv14SoYCfOtSw7tmSzW9HinjZEWbEsM
p5nI6fh8gbA+yOOvqq1R4c2LEP3UxR0I1qTU9kZ7AjEL6eV8MtKSEh2uJONvlr/o
sR3ocqC+9xNNiNJW89ih7yFJX8nvPVx+jIIlT42tqHYkRzvpyHBeXK9RoYd/3JoR
MS4S5g+lq1plnFeGNBSQyBLJKrEEBkZcWb37gae4eX4XLMfG8w7zwLU8IOnNe8ap
CUyHa80TDJRZisnq1mJcb+8zdwL6KBO96BTGSUGIDcJZBO8DCTTqUCpJzE5woarH
bACUY2t7tutXrtkm8LfpQi010Ku7btkAe7hRKB3frOZgajLI+C+ArulWg36LPGwu
otkg/ZOKzZzOyodCWDV76/MzmrO90opZ7rDCgu806JSS8d6tFN9ot1zI005qIeMs
cfN6XraFJY4zSgtJrdgD5waj1e60516RAWYInVJWHJV0+jJ+cKXpOcQ6IzuYEzs2
F4siG5i7Gn8qreqJg15uTFlkTcMArf2hdSCDWK+CWutI+2LVmZo5rJ9m4tOJanhi
dRsuJ6kXDpWokn4Cj+Nw3tqPJqpbHBX4w0vPAkj5jj5rTPygtHjj9x2MI7einy6q
1oMT5/abWxFCcAjSVlOPQFFm9YegyaGfcJubFnksFlFzI930xrajumdo5m09rbao
NGRWEmel8qBGCb15s9JF9aA72gTq0g2ajsJQ4QPGLJjo6qpjAdP5cO268N6syBcx
D0dI80+Z593oEgwbEhaM157Pr/12LgYntcEnQl97Slyx4B6eT4Ya9PTSObkmSd8O
qqvXYc8w3bWnvCHtios5rn0X/azCWX0yXSzSgvlMGMUxoSBRLBwGATPCMf3FOYPF
nCybviPCAkTxRYGyvJkc/P6SciOHAL4RxfVXCSE5L0ndGcEtqYELaS5c1kbxtMUk
e0PKOs8mHdxy0YdxeKpm+Ue3P+RiePmvM90Jvd4MY0JRN9KLbFZQ8aHlNI0il/xr
ANNA+r/fkufdELYOAKR6Oliud2xg539hZX3S73AmcWVPnXo5e3GciSE5XJEAHYno
PT093Ftw7mmRSRpj0UGHX0EWYRUQ/A+p2nlqvMqY46i/VFNiAfm9xGZk0Q8S+FYN
Yl0b6fK4kcjUR8YAO+Dl6hGVf16j3KfhF3yCuqvxQbARKqIAiDZfoSRBQ5+kd34L
W+vpbkAtfBvSNqCpTqcDBY2HtLlsubGkXitut2UIXpkRqDl3gJX7149UqN4Xf3VB
JXCyP0bneC18gvbvrrSiq0JpGUN8dqXXkkzvzNFZKHk8nqWeVoP7iEpVN8XXUWMW
3Jb+eulMrNR6bGex4NG/JgzWR92Oj1R7f2YXwsmvr4n8RfQnutl65UoSS1REZCh/
dObRl78yF4Z8/AuCJtsbiHcDvIzLhhPEvlhuCeLjgR9UcTcPb40gmgkiEazl1PN9
juHJd6q/oc8JTGC7sx41LMpITFhdJRtTTXR53LBdxFC43wogcROyQHSKiFzvUKyt
yWooA6+9hGBNQsMaF2w7O1zwxm6Mszq8JGgKCLLL7Qjm2o1DsVCyRquT08PqI8oD
OfDTzsqcyClND4kvbsGbrTM6oHhKv+V9E2UUszkWJJ2GvMK0R3trZTzihW6iprRz
0m8KwhjHGh39GEV5k74fM8CEa10wrCDBK2rKZUYh8KhtuSSgAROxMyzUOrza/csS
QdO4HFTgn0PR1fmK5gpyum4vXT6+isYVby5Wp6T5LFlN7dJ7UrAizHt4pepmyxRo
GwNuVnqBBnE9AEaFuV/g48leTrtBCf3v/dkb3Iq9dnySTCoSwdkuq/1MIxptTH+Y
xFnYr0AKM3dRxXy9eMBbE0DovpQi42tcHqJjcSL3cxxbQYgFJ0UDskgJQBjjsoNz
38Xrq3s8cRtNN5XKFwVjW1NCR5jSxtg1+C/sC8Vsz2BLwHxEC+0K9gUrOWz6dCUM
50M6+skcU/dLUwCz3Q4gWshMvmNLRGWFxx6L6G1zLvjwWoCXnTxRHCpnWwR/y9Gb
RQeAL8QIFBcwg0trTBq4daatnoJ07X+/UmNxzgjn/Yr3yDtcIrLXo0UECZlmrKEy
tl3hNhZNYK5tk9TwZu+UAc0j1VxKB/zWSxCl8yGzlDR+F1EGJ0p8GooGFkpQEFn4
4xqpuT0aZ2Zm8yookUcnZXbomnXXu4qPwYkI9wSw7jWohL7+Winl5f1+XamJ+9sO
pHk2DSZo6OcUvHDj/V3AjP4hhUOm+h/P1E+7jGMota+GE58r5DnjdDiFuDOKK8PH
xLpwbqODyoQ7UXjG40Zz84uD18aL1bbsGitlr1EfCqNGqk1HlLA5DnPtX2CZCRh4
3543KPSQ6udzw+iJ94BGMPJz09wxSDZv3myKPyw5u+oCkAOEmE8oW6sli+S2fyDn
0YoyWMPILYzzlaFXnzM1s7faTs39yjrYf6Of2Ta2r56InJRGZ9VOpWueBTc2qW1z
ao2uyOTGNVaLQqfYSdAxvkXUavLtLzfZXoMylqYKCECktbr1/hgNs3/ABjZ0CdxF
4nNtsMGJkvh9N3MZG1iSTQS5OvOlQ3azfHTgU6eDZOf1SEyo1OFg7GnHKLTtjMBF
byos8he7OW+L4mNdcf27W1XnvG765SQp62tLa5GoVbO7vILz/itXsvOLTsLJ8FE1
xBRa0nDwMx+XAKoABgE6jMX1EBAajP9nQjkhhgX4o4vG4y5EAW5b3PycCwcQ1QVA
i2tCAI3Cv3I30QGlcQVDxA1UTidpNecNib9S2rhui9lwy6yjiJv0EJRWDLwNa090
WHpw445dzsgLt0c+T6pEHKymKNLXYMUYOjsumgV2azyoKlU1c9qrKAGxrhbJhV/I
vQxoV7myAUjQpUwpC8hCqi62zjdZfqao/8H6PhsRySOus3Q96fEdrM9vYVT898L6
np5I1abxJ16KK4sdAiZV0NL+9nEqQmj+mD3gvlmmAVuJF5SQva/+NIB0mj6yOgiy
9yHRvBzgfk55zD3ZeLn+phHhZtSzmNi33HNp8OE1JrUMfAuhhO3h/76tEWg8M3sV
xoY8w4+R8LM0CWMQwY5WEClmgknOUFS/SHrcLphyDhpQ2Rwu9uD97EZJtR+60qnH
Dhbe6cE+p5cPNH3ih3LFtImqvwNmpsWjXflaepOeMX7UmGWdqlhjng0BezmUYkRZ
3ERhFW5wvBY5hURGsTmbDrD716VcH6SJT1hh+Ks1d0msWcSlhuPk9EeHLzT23tAX
AhEvjtsqLIgF6QNuUGKeaTlysZzxcZbqP+RwkX8njj+2ChocETUrzvODmUgqQuS6
WngIuzOwrH8MohQSLpgtOhyI1jrgKkCHI4PmzBFi3h8YNKy2y+1vsT/qT2KE3H/k
NU2xJT+ayaIb4gcOU1fMQPLxjKtzHMkGboYWwkkzbvo/YiSQKRb+O2k/PQMJklZG
F2CyKF/bfUCQ54Vqd/zk0LrUDBKZodw/uqsxtNAL7V+45hrUSclOnr2ZYfV07ech
bSXKg4iJ1+qADWHxe8dm72PenolBJI+mBMiBT3Zq7yxMRwQWEesb3PVSZpwp0w1+
9E9lErlmtLCpIHdZDpIqH9+M2KFbdiHfZxlZUe6dQV5SCpVcWEVDL46jNoEkv52J
y0fV2oDuyY2O8F/oeIN3Jv6xfg9xtbn2ZLvGrmIMnh97kZ67030rNEHg+QlFpsi3
6ax/T1KHrAh8VAH3ZNDeX1ueBGq/8d3ffHjOE6e8YaTH4WcJQeptmRJDcAhq4wnJ
I4vMBVXoOOunhJerNltf9lv3h+LnkzjBNZIGu+mD2yr055pBNSlHBlCjHZoy6A17
FrVT4orq4D/sCtF1gGBmLnHgcVIIgn18nKfGqlGykXKDqu2FlFO1HmTF9sabVe7T
hdNt9G39kaDssRahHQuKM4bgcoFnvp4jI1664NFihd2pjfVizmEXnnT5IcVatlPB
byvr24CJ1hEBTTBfH5O5yxmqQNGnZDlPC8YlaeDUzhc/3Lm4xHDlXzUMcjhaLom4
wNJgdmPaX1DtG+dYHv+Ls4Ykbc5UHOWZ02JkVlG+kdG45OG3fcCCM//aVqHyi4OZ
oEXDeJEww8YHaXbYSC43fmJ1+knL2p8nSmbuB5JBAukMS8wBQ5k84y/5m++DEAxE
vS0uJCMTgUOLRYKCYkKfjNjzEpW8dLW0iINgH5pKIHXojwjQyQGwRKWP8MfS6s1Y
aJvPT54uS/zUvViwgY6qDy23DUKGdiN9xzYm/o/plAayQTF3rtxeRpnkwwhAQgD0
A/d7rpwYpMuvSxr4ddBPMylkl4vAA8JY5wmo1BEJU7qBY0OnVhTZKIA5z8Qr7CqY
LKIsZ779buCEgL86m1gz8goYhDKPVtVQ8Kw55Kz1MJKE1Bkl/Fg8Z+BZwyyewYSF
ygYXb5EsMQoEEXHp0KC09qLJugKf78W12UVHThOs5FwwtM5Nb1V8N13XIHYCrkQS
8db6LB5OydqtDUrm4N0Fs2zdEbS6dBuAeDTjVIyQ0j74eBYSrxuSHGM8Jft8/oWy
d0Qg53Yd8zCJa4VxTKCquOaNh6WRKJ/clrwhg058DbYyH9fDR1EyR4lshDBQhZ/k
8CnRORT35i1MIyh9Am5JY5EE8XrM9K1rhTJi2j7s0ZlBVCvJ1GlD5Jgnfuu/wLsl
0ta9o/pJY0vJq5aWXN1GviWGw9gO1WPjfrdm6d0mZnvTj29GMi6k3thSENbumbmJ
Y03wkVYiW9WW9FPlYUfJgX6EhD90DxXhnmkpDxvyftzoIGxXSFJRpsNKBEeNQM7R
kECNWhW0lcKkASKaLGo1kVFG2Y0i/++gsMwJnnwKGkUFAB3FH8o8GO8GXXkIkOlS
Tt3lHWCB5fAdYvRuL1WaSCef6pgOu+Ea8y5r/xIjMXTneynAl6JOWpVtz/VcN2GM
wWk8NqeJG1VTQSnd++hrPbpzCULG3ndSHNK0CNFxk090Jvz728CM8cSIL6FItkoT
jdlY185wvQOC/o6XL3d9WW5enGR3DuXNHQXYqpbYS93ykuUxByvm/Zlb+W36ZA7B
rKgvw8Sz2+RsvLvjMvyQ3JKnXSWDDW50p9YspEhDEPUhLsAWF4ZMfF2W5vqWmgj9
JHZ3Ulq1mIeDVeTKM0TSa2Lr4Tf4nMEraek86rL2cmY8ZO9+KXMrfYZE4k5dD4Pr
UQJKwbO461vicJsrTMcWOwEDgvPxTzbLD2bcy5vCRIi8yDbACfjgIrdBTo3WTQlv
hnHdrSa813umfr1TEvWNszJdoD2ui/zR/bwhH0NZylcVi0oVT+IFKLTRZox3y4aT
AZ8QqkJE+/Jtm7+Q+eCy6w6javm4zWFZfWD0rbnhk6POCCaanr8PQ2J32J2gwd9D
KgntEj2lfG7izSQLPqufuBxV45ZgC+km4c/Yh7m6j4IXu7ICxHLRw7Q0d0ZdeHsk
oxpaIabO8kZ8097Gy1o4ptNGWZJMXM2V4Q49CG32Nt0DT2tAjJWPp5RQjozWERcR
XBaKvbKf6YjjULbDp1TninZesF8BMiwMuo9+AQzO2M+EVfDpWNGb66vQqmJF01RI
62b3Se1wQeS0ux+Kp+m3MtrBAPSm7XfZLfanQj8LgHr4vRoa2NI74GfdAX2aSCiR
8u+2k4IsErGXN5AuslJJwiDnVm7yj1ivNbL0UtOqV+sPOv1Q9CsDHGMd0KXyTZoi
JBpOluWWckhacmNENvwYKHiPoB0gPGGnpn97O8RcffBOqq7V5055vkqY+nMKwslZ
UDoD8AQItaU+rrUCDpoA1Zm/LnwMg3nP2WcxnGcwFAJSMMBTIm0VGOLYT8On1bqP
nKBFVOIJZbkjrABY7wVnm/Hk+1bleLSZjJCJzYsIgAgiY8eE/rXnF9U0XwIR3/8f
Mp3NViN9s/+dQD5j9z860yhNaAV+Vx+2P8dqANHhB/WQiLcOUm3HKtkg61jeNa+E
XSX/IR24zQeXZIdtqaUuuElxfJC0GtT9IBxpvRVdLsXa9rvpOVThTZ4EDCn0HBy9
1FfCZl7uf+38amj/lKEfpY9JxmOzQlNMLVGwpWhsjFCpETsqN89g0OYcW+U3MEAe
QR3kVVQWasyl14js07dFerYW9ihivaYX5KxGI7Ld4MiZoRqq5ncfyLr3AfXlEoyz
kzG4uDVEUwJfqZNn3OgqU1zpjtNzPYGuw4RXqgYrQyMS0LqzlbWC2hO6w87TA7KY
x1NmBv9Dz2u3UxjVLrk9By5HZU/U3Lg9+oB1YxrEb1jboxeHDNS7IMrnQI1q8nmW
dmlAVgYvVj+xWHyDJJS/Ko+cNSsZbosNqhowkBM9wUs+8o3S2XD/7d3RMquBUo0S
L9OJGwd1eEO7Vp8zVUh8WqTOth+GYeijOm1TuTAH/N/BVu2Q1xMB5qgutYhBqjlE
zEgkx4ZIRKl91/WlWyImCOAGhQjhTj4HSKrAK8TQ7GNTTjP5LV+9jP5JJAvLbJvp
r9RoH4XglXFsRQKz/tiq98dQ5YXkr+VWtUU5BF18KawoZsngeX3ZhpMD17D7EDnr
wIS7wYClhcRGS24rwW63tbjARiCAssY4pgInCrE+LMN7g7CJ3HcehkFbE2dR52KP
qyCMZ/PqUb9kgNydXZywDgLHc+X44foMroWck7ai6liZSUk2ZvMLmleYSlb6ofFr
bWSIPWyIovS4AMkt2Hv6HcvydaiPFL3Giy91eMdfJSD3qBC4IBQwYNw7e6c0EwA8
cdCTP4Uyz6uH/lMZs7tric3V243QLOEkc89smKcEJE+67P6zwx/snt4FLE9npIYg
dpPHiJRYmNOLfRqK0X7lIUR/V0qAeToT5JFQPZxkZL841oNiTQGVJ4WwNAxTFz2r
dz0C+NnA2omqeerkMtH8pXTA9ulnIUtFQzkqySD1pCbsUGiAyVBXWnRm0S9HYo9N
Bwfrc8sRH8bHC47FMVhM1/B0V8wnsuUcuV2Ija5ksV0CLoxQXlLBU4yVchUagutq
9ApbTO1h+5dJhdfRvtnCQpT5KFuFEMhZsYhWr68JHBoyaxWnfZmeKznP2j2yXYyb
9tXbnh+pt/vpa3gS+RthAZfriXNUHI1aAtNpcWxqT+Tqbrltons1WsoBwVnnqfcB
1YQJkiQNwCNVqRImAz20lUuE64XS0gPCl7m0bKGtuPhJ3PPAG5v5PPaWbZkGJ/uA
vGO+8B9dKzG8igCb2RIZn1djZZ4BaWcQolJGAdnVLCzE3aqYkdTzuNQH3sg4oYoO
J0h+DMxvE4i2ktRoiBlJYdKbSA2igGhfgrL/HJUfgbmUq0KDOYebACmMW8Ty5thT
Kls72gterpQb1gaOPkpA3zBsvmkIhIYf+dS3mXFmSEfk7Q6HGBCxJGdsJTc8Dw/N
qHc7dRCnVqdGHFC5xSqTx+XZrD/p6VoP0VpvvKGl/A0oWD8CjbUnswIJIt2CBD7K
gqvw+tXMLjL9CO2S+XRKAN+lj1NikhlRBqb5G23lKt+23hm/JZX2l9AaL0LIBzLG
dppkbfzLjs+qCb3fW9kmPi6bcTk72ko62DaGLXsO6l20l6flAWl8ptrWjoREPqDg
L5zNJ7nNMYxSVKDweMjNOzOG8xc7MrDJlak/XgkG/6YnCZAmhZYm4bQYppDqskoz
o8ptA+J8UT5mBZVgyGnTLeIG/eFMB2/R+r4yFRrx+GDMyusYWoncgXHXOnLo1N9H
AXhGHjJ6MDcw2lQAV0BXY9M5c5SSKyEa5O7pzi9baLmHq7aA4nrmuRVoJAtIlOdk
89/dtGkRnBPzPamuKjr7++FfMrYsSTWTLl7f15l1WnD85FkBNPv1NxNqOSHxYiuD
eaCzw+QaLxwj+NY7dBt46Qyg7Al9c7UFtTwS82ch4SWLueiqfiXVaC+MzNDRh23T
KFoXS+gTAGLmPcuour6FtodstuojZX1/PgNq6GXqYOYUpJtlHhCaTGpj8N6yNb2c
6xLRCXN7y4zQR2Kla5f6WH/N86M/ujh8BniElRvrUYbGCtfoyhU+hrwGoxOnhMgP
UnPOU4j5RsKQFhBK/IE2BBb4eDZDVRu06EtJ63UE0ZQBtlaVpeTjOjoQtOf0Uvxo
ED+WbA+i6HLovm1mdaYdaVwr3/R8KbPK4kmDZQWqXjR/sSfcgNYTW6JaIldFlXM+
+3JYvXDGIOT//NbVJY4otxWtN2WXhGmD9FVV0OvEFzHFVYn/+z/MUHjY61iN+IKs
T12WJvE9g7nAyp0S0KeMBRBCdpRJTqETSfygisYKLCv1n0xxRssCqtJ/8hLwMqc6
/NbmovF14P6TRbPLp+csuvGuNd2iTwstBR/yFzxCLUWWCViElzGuIn/iWPIT2W4S
O5SSgK3zC+LaNy6kvuA9R1/FcWTbEDi4s5UctqjaUBUYX+Dyq/mSefc7Dkm3V98L
k4nf6JT+FF71Heh1p2QWQw57vfIR0w2kFXXvCBu4b17oeoH2bk+CnP5VTjjln9LX
66LLstaQXcEJslhM2tz1b8ZbEtDCsbcoJLL8JkZ/RVww2JiNPBo4dJ5/ua0Wnmxa
XtamLxSPYu+8KArUXKQ15W/65UwDfP7qI38DCbOJgCUkBdOnqmW2rvr1U7cwj31q
IpX+Q/yhoPM8NolgNTvDXIdyrsZ496Y0CrIgllHkAvUIqIH96wXIsF6cSJq5xxUZ
fkfqZQKKC8y9vpQmSWOQC94bzTdO53WVCr3pKk/IxaKen4JuopZKgzKItZy556PF
dIaP4SPNw3kuf5FZUHMOqLSi3bbuYU8RO/7/imwYe6LRLI1kxC3RTs+laSsMnJX3
fLPZM9LTWq2TzYHe6KgYc6BvsAh2iQIxL5UKKEwYWoq8Zj9x2c+usWehlv1EpQ05
fX67/fSzijkYm9ubBKUXhpOadZL9Q5QNm9Kv7XBrqz1Ur3GmoD30IFaEUNSzRiAI
UXC3tK4mKt9/Dnj2KF+ZpnHXTh4VASOACw6I95OXq7Yyt5PsqSdzKIPMR7x9gqs0
msEZeOkm/ZXuoSxd7LETtroHRiC6kQJJX7940Zp+6MKtytJ5vPjcbm4grvQtjAyG
1q9VmhUQwbUjh+7P7wmtKxTG6v8bc5TzGbseG3LlA3s6A/d4Gd9Re0OFvvmn09I5
JYh0pY0esbJyXSRFYl9vowbGPSTKkmvfb67xYf3B7wi1Qbh1RqEOUXkU/ajexDzH
PxbEQpsT/7EVbx0OV4aSUftp6JlRkg2VSVJMfgR2zZPhiKdmZVsB7KBslyTdya2J
wdIudYw9q0EOyAA5gaxcWcKZ2J7JhrKlr/EGhtHTdFPCRKmnIox3mgB8BAeW3gz/
4guEv73MGTdaeBV513xYYlZhHDDaBji+uC16qPtG82fZo/52/RPTbYxwS1dFo87Q
phRhT4z29jVWMZTHyQviq9noAo7KhPtxgHNzm6KpZCViMQB2+R83qnHKzTVuFM0M
xHg7SQUpw9hdutJ+6X6705tUqes0jxHj1n5Nb4mDWSa/HZSqHKjP30RMy5ac9mxA
7NtaRh4Hhr/k5reTwS/hw9YKK5QF2ETENF+EnethWwLViNPnAHPgaFufgfSwkc0A
JXoEni90YWXhlHQ8NMtTr+lwRACQRdeqj+7jv7bx5+rwbDIWUjdv27dMsgvi4zeQ
Xfr8rl8esaCSn18RHQ4GBOcfzwUMreqK3lMn7Tqt5UF1WIOamFLKviIxl8VU0M8J
gQZuQlHazgTCZuS5OI2HUXffzFa9AgayTNC9+WdDU2o10spf5JH3HWvARiOM6Ux2
P2tjRf2+ryykGTuHJFcIA2a+fWI7GDt4SaZ5YnqaxBmAgv9va8+jCYW29l4nfkpx
PAjIDha4DXGrwt/pmIc17Al1Fw0jdvDhuNRId3m3Q3xzBE+R2lvY73LIabvl0LMT
glyPrDcQAUZE1FO40P8yK5oq8zJUxY3ReFVDQlxrjSH0Zrr3oKyH4dwq2vWqXjnn
VQ+9Ycj1IOMLdu+R6Z4jUm63CdyCGDXyo3+C6OTsSvZX5xjtRlTonmEwbTtI59Xa
7U1S41TsQVkigaSiWoBrdeIK4auA6Mh76xUb7PM4H2ZxnKMLdjvLtAv+sS4QX6Po
xNIkrZZKY947kr22vQbrKjytFdmsIkf6Gqs4YnjzKgtKStvojd/5BWnJUTQ05Zeg
zR7AmV+1zUcIWitEq1rWOiPwHA/0LneNjX213PS0NhUed9zNhaI1CNVk7AyNjtSO
qR0OKsSWiq0Lja/PgKRR7myZXfVRR+H0KROrnujL39zUPJn/zQONoUUuvEOCRpkb
BnpN6BXJCID5fy5oW4dl6VSebrmaU1xgZfZ3xRsGWablIuSiQJkf3zeuDhnrnDRg
VYi4FA2FxHb/BOmRBmO+1jAWo0wwDXgF2uyEwbmvxiyySQVo86Tky8RUjHeeYiAh
p8bv2PZQ8dkYLhlkZoQpeYij7HQ9GKrD2qmx4R3likBJCk6he4CfD4t6vuzQdsKx
kOJNPKuY14NuIGXSBS2ekyx9wVm6eRMZA9/zXeXpOSDuabjvi9+FOAGrWRC+6jH4
9mMyDtIFzgq/LP4GGiJWVINleAZWS9A2axOvbN8W9RQ7Wh/egdmxA/5+TFkwnJ7X
ZYCUP/zMVs22NtebaB+U3rcxbx/fFu662Wnv5nu2uLReuS8Ylrq8B8nbXzYbn64F
y5SiolOu3qDzL+Z/2p6m973+Ax7Rjv8Y6zdhghrgf6u3RkM1kTSnE9KLNKVd4IBB
d4/vRmWbOZTl5/VwsdReVzrgOiVBfGqPrAFDX3vD66GDgPgbfeX1vxodVdWSDwOT
/tpN2jWs29ipB52l94mOmebHOVbVg97BKsEpI+UzRIC+rFgE57mHqNEF8MSagp7l
LpIN5j4DYqOQkOwZ8dD553+4qiPt3tEK58hPBP8SlD5o422WJSf6SEvPN3st6mqf
zASwsueHy7SpU0gfO1eZMpQ+8h/GNqFRQn+os9kh6sbnyKr38x/W95XRtzC4Ogba
k6KtiJ5lTND2s3E9xjICM1dd0aJgfJpJWRLosUnFjZAb3mIVWCpXdII0v9/Zt0Fv
9LVM5GYOzr0gfhonRpIM+/ulN3bUerDTlX4hi1GDHvtEJ1f/Xje+6OAndVNgDMW3
KyNnzxbViwo4fVPZ39aIq2lYx2xDTSqiR2Xh6+ksViOjF2PPp0SOeqbjt+5T457j
5yxbmrKrfidUpiOE3C6O+yR1XmJRg9mD+yRQz7pH5nuPveGglLaACp1eNo+m79QT
BO/KtwdVTaXl2tb9V7dRhQBkFZ33v4B61ZIR3dWpl4b1FFy6ta9k+s4XQ5QmOuwk
8WkRrhehr+GMyDxquHzmiHRdOTmRH1WqAaqnK5DN42ZiiB2RCGT5CdwQ7HqpK2Yw
Cj6kl0RPRIHXNwdPW/yKHRHHZbh5hoYITty43EkDdhqQm/RVD2yE/5UVEjmaGZbc
zyCkvflpUMk0cXNSNIBYp8ny80ItgFnfdjdJ+Pr+QV9jHGV3Im2vMSmPjdGBC3ll
2FTIGHUtGsH68aQ30d4H3005qv/MsqgrGgXQIh16qsmd+sPhL/c4cm4bFu3LUKf5
A5UJzePLxxYgqioxTa8wHw3LReB8rkUjJn7ahHXtaOAJs5B5lxew+p+UH1ITSd/e
lF1ESlwaaEwgdCdFMDmZAmMAZgvhQWdaPVgC+PU7eojWFkG/Q1YkwkBzQsVQuhUl
FFfpRv/uONQTDYyArkKgp1uVe+yZsZ25S12212Z/ldalnqM3t2K7W5xhxXAKwd9v
/TBZfA+wnm7listNr4HExdZwFSBYcUKdzZOAmRtfUUURcw2Y3wBTWpS5NiVhGvQ3
9WGBW65G/Rk3nxCJKkDfLQay5DGOLw6yiy4lq0zYJKZ8wgXIZHUv1GqNihEY3jiE
dsODdrg8NOubrYycFY3vzFuD+EUycol8mBUBS0fMOzOprlV5P3BkN0X0sJ+/cxe7
lgSyXyGY87WzawRu1zAkJsXalo7+J9KBdqErUDMb1geoOZGm1EdV4GCajn9u1Wet
o7Pj/dom73o65B78aLVGF0dOhryMOiWFDNTnbD015UA0oQp3OUzcP35l3XMMsbrL
l2IFjwrjH9ccx46t5XQhojyd/LQS9gRggWASZ9oj41bGUjZopsj3IjjpRUwlTAII
QtIiHaSt5VDFDp/8JXCwxTeIH7owS/+ZxjTd3hI/2UVugCdEZL+tt2HglZhPdFuj
ERMB6J35eoFAfbBb73dJiq+G/qLM/w+bdYLbG/skLb4axQG/TE5bnOArkLrbSqjW
8EoJxqXp0uTZe+rsOp69RvZYNm5wUHhHxsPNofdG3rA9UD57qkdhGLpsw1hagws2
jW/pBXGhSpNJgdItYkHW8/0h+H3cOHyNSJf+2NdZrU7mvxE4XNHluoSxb28lHSpo
E/jlEEsfhGEGAHpjLsdzrqFChti1/D0M3DrwuK9/2cdaIXUoOSjAu7z/hj8fmtbJ
z+lYcSISCLmkzQZ1Ea3X0ZvDHm/u6bMw7WTdi41t7aHIsu7upVUNmwoEclwIzBze
G7s3tIS0jXL2Ks9MbfrkLAJFbG3yopeBGcOKccHso6P0jHaJWSSGMfPj/8ATkbNO
zaz50s5duPcUWqwOFPfRCw+sqfSqP6ytH3mo6DiuYtNOGHHXmFsIufI3Aoqrd70I
erqHMwK0yk5sz8l4XRZz+95j4daW1OUAd6NZi7iY7Z2irLeqLO22GmitkR0EBzm6
4rA1uzBXXxHw8F4gFVZh3rOd7buIFaRwxsXljerB4UYqVIepiXB7miyA8h3W957u
8/OyCiYrvFdD4zxWNTvxzDf6wLccceJBDR2BVYb5sJbJSrrvI6RFrxWG8lwWj3wM
raiUfrhTVnEh4pEJ9Uzz1zuAmufLZSAhV6NMnPbbR6E/VHwBhpthfTOH3UyWYxk5
k9Zgz5D4v5Kt9YbThTfGceiKJkj+sPAJNDELjiSvBUcOe0VM/PYCo/HnJ1HDSutp
FfiiGhfci59GZ3FEYZ2Amp/y3IQI227H7DkHW4fFdT343siy6LHHtcMsx6ueXdV2
sb1PDBgoPKq+PKQqjsjT1L5KGSMTh9l6ywCRQWEj2/fYGDDnjLpZClxpG3qkoDy0
XPGW2ROP+DzJEoMbTyke8BLt/NuEW3jVtv57YRAziRn2rlb3wM73lIFuObQ4UxS3
RDThaHhHcfkajQZ9EcesXSV/4JmuASsZJSZa/xikd1VOucxTmppxkD1BzbDutiI4
3jGJbQOy+FjdOyacCSN62Mq8Uiw2o+X2Oy/awRrxLqn9bwSLVhO/jtBRF8sFrnZF
nf0nXOosgohpugP5ecXr4AamAd9LejT2p7/pTvPfojJ8+b7ryhmCFfDPUuUhtAUF
lyQm4c5JZ04SsplYOo2UigojA4hJC+Jrl01WuE8H4/MRE6+82x8btkd1JAK6a613
4rKTTG9k41Nh8GVy+SNV8PanHM4dPFPFGPO52UlxTfe4OEn06Qw+tMgmOK7On1oi
MAWO10nta39UmrOvSUOMK3fWPTUOWjx3i0ieHBBJH/dc4TlffHoCEBsVJ6Bn2PH4
/IoJJi+OEEPO+cPK1R1X2195WIF5AjfOLzoK41bGbG4KMwCPi+NnYDyoe8oTVQyh
+OApH9uIdG+2XQsAVnFtb90r7vsULaD+jwxcaHPibbgA1Ly7LSJCooDQB0I6eZWb
w0oJxJaXWRCUyXXibFkovY5YwIbnR//bb1kPb8wQNTTcC8rDjD3m7KaAaNOaUzJb
cIuh9HYJyeKidAOCjDX8Wv9dvrGDHfKjjWGBTFZPsfzGhI2iVEO0fJ9kvWC1Yo1p
MDawzlYAwmZ9KUie4TcEnfCQIg/5NJJodJ2UEGwNPDwLuxnS8BqjZgfgX+i2OPot
No3UZV/26K9sd8FA9PXcFhcTrKc0xBK1H2G1ZaeSdBwR2eW/ENrUT36edcd28FoI
+GaEmszUybgWi0eNMNeWHcVDix4v5pAQ+34pfzuti6ZOGtqUYHwgNhJ2eWzD8wcf
xrEHqhLSifEyOZJEcRkQ7QEXRU1IY1Fk5OaPfpHM5BjKJwlvBo7GxjTs/3j7DN39
d0wOCd76MduE42OWbwvUuLz2q0PY00n6U1wMdNRIqLVlzN+xIWDF9Qqz9eXVZv3g
ZIHFmyqBypK8ipY+duV+f9mTjNK45NaATr1Gk13CrlioyTIsbNhRxNSSpe3FaMo4
3WwA7oyCTkz+LRRvUJjMqRNsuGxSXiOlzPcTby1DfOit6g4Jl7FsxzzZi/KFAjVV
K9Y785NOYkLbxXEd0y0KPay9T0jhvhkoZQtOhXXUIsiKlN5La+zWf5jVPCWNdN3c
FEo5unV1HH8S/j35S7uJVTs8xb66xdPQusJyVAr+5NdkIbhvM19MtGAzUTFUmSiu
sZusrEXawpTCDQNmoiNPj7cizOgq4Acxhgd5vkyG3YoguqElP8c4hU/IBEOU/mOe
CaoKT9QHfaBNuCLGXQF7QDDytT7ac5ozaBuDiXHZ455X9MZ4XfiWigLQal/uqhAj
+scBLOy4dlzEGKPgIV6GIQtxeSf0FvOJPmXPG2E7+t6yjCtsx7S+3LyTcVDeGifq
Ql9s+CKMkVFLQfVSlIJzj0wCvMQ5EFbvfS2g+2ktoXIE6yVwVNp+i501Psn7jvjj
g4PJ/+obwhuH1I22WtoEME4MdknmobBqt2PM3WNXiQhTRL1guHrVY2gv1Nmqdhj2
Nxn56H3QyaOwVvOpAiVdWBj3B5VQCj7atyzHRI7hP1AXrUy5FtgeIM88v51rM+Cz
xTRL4YdOuS5Dws9FjaxPXG0wa5q+EQzDI5MXHVCb8scLNx7hwnrVEUHbwTck/i+Z
fVBXYOuSxywBZZ4cjq+IMEqHr0fA8lkKznI5smT1scl0ag+zGotLoDjOT+kauHkw
SWAbMadIGcEfli1HHUDhW0kV3UAaY85JjhFq7zgKVwrkVmThpLi28VqQXmvx1GHu
hbmdTh1O8YQ60mNeagnWC/k3hpMVrDM7DnOIUCp7faNy+6Qmy9FmW1SGLp9JwQCs
FrvBrKPjzpV/bu4dapM0craD3l+YTr8FcwfffIUZOO/47W2kRWBdrmZ504b3fPIA
dParsL+/0PKffajpnBwzx6bMS+A9vHMKDRGcdPeiWHaTkOJLGa7PZdEI0DoZI5eT
ZU5676ZbFKJ4ItVjTkMKdc73soelkxryUd+FMA9z0MlwDfdJuWYITEAjSp+GwNWp
9t8OPhEaYvJqwBmYqQUQSe7WhedI+spWE0lbpYp+HNW8uNrBZ8hCNas4OxeNe/V9
dGgHWCC48zfB0+NchT9NZhuDH4EOXnkyqV6r6nrtSRIveUHxBDvro6+cmzHT+uHX
GYen6bXy3jYoyW9uxG25JgUKmiwdBYqt0M4URX8ZqnjpLStrS0oJSeNV26WOAKrH
Z68qE2hwLad6Y+vs9k3AFlZUZqIc60Mfs0cisGhsb37fhj047QWL/ae9+D7yXeXk
A85XSUlHmKcQv2lYenqbbFt7Ih83hRTl21cCRfgxX3h2gvsA0qC4QhfWi1MRwYQQ
w2NciGkfcsRGbvZKw6lPkWUZPPKrAu+Iiiac2YI9/w4s4o6EvvLCxPHXNuQdos0K
QmxwhgDmqP1A9eKIQe58OZyCY0H5nIqUeMQ7yuaUpteA38wBsou7YuN6mSBIyYgD
PGdz39HczuCzvGZR1hpqF+TAf+5CsQjeKILYUB6JFYWsDSTGxBpkrtbgBkyh1X0C
piDKJt5uPhlyugvtdj+BECfHqhZ2pal5psPbDRac8iPnPxevEKI7oWlK5t9jsbl3
1Dk0oz3zVexJnt1kbyVN6Pp/vKgB4D/bYfLssyKpGQZFF8P+QBSMUbPnEt7gDxJP
7LnGgnx2BUxXf/634DT0lckMqsRqvEfd+6utyByL6COJk7MB1SgVjCEjwnfr9GUo
mxh8SuNs2SviK7vsIdC9SPJsjqiRCuds8DzK3/5i5mcuLBcs4KqEKnxjIvwDTwm5
Ws4RPjUc2JVNgq5MqHs3L6qZd1h8N37OcCnYKimdFPKV7Dk0Rsc6ZoP7DgRebMrj
EIGnaVzMSufADpWtL2WCy7QIh6O0q9RgdGxi1e5uWtMovMFCCqTVMQ4aNbSxPIjG
SSraRefHz0Ji0nIzDZ72/UQk5HFOQKesLu7GG8MylSCZJXmHvMykjQEbGwiUPXci
MgNGCZhbc8X+4hFYA7phRbUy09wAiK+0+a+EN/d3SQgpDM0rTmop+ZcmqPolAU5E
Ejj76ZUCJDzRVZ8pqP3nqqx5ycYAMov1QZvVK6vu6b22F2THDrdcqqsUkwE/Oa/8
aHxqaoNzonlGiw6itFq4KU7hktrrLNYqcdvm+0g7JLybh5DBjpMbxJRvd+icucoh
Ka5rBE6OaDqpmLKd0SKSX8e0fOKf9JvagCx04YXS4pvs6sUbCgMBfOcNFtFQsprC
xvFLGWLs6dNwoOMdO7tCdTNdLMEEVPNFCSKUGSykkKi3kTvaOwx/c9gHvrdGU5X5
UFup3XGUrc3IA0ERYxsokD5KHq82Xs9fYAHWjuljdBzHUiBrgUowgbGsPZL9h9an
vC8T1mvmHwbWSsbyjwxM1OOeCEOTpghvHD7HrwRq0YPcBhZIuzM9POxsdIvyjXwc
P0ohaNfzJRgiKGSSJWoboxPdMM2hKXPOUa1C+F/8FToM71DxFNJxmsKqMI+kKuH3
65CZqJbk468YasurAyZv0DmgmYQOC9xnkoMUOaWnoj1XggqJG8qqzYF9PlseYv6Y
Zw2TqBGy1v+0UBELG4Xm5h7hzUqbzAbKlVmKYAwXemgWjeQ5hixVM/U1LsA+e6tf
EFya4Dq+vfKXwdNXkTebod/MqkeBv9807HUY+/Ujy9B/z4jdL3TBLTLpnE4uir3g
VNwh30eX39Mo9N+Bu7gYLU97rk1K1svmhC4zSty/4RcWOEnQ/suNrCJmZip/vDoN
UjOqgvSEiyzPxsZ2jG6iISUDp6sgauzO7WLSd15qVWcLO9l4WwOPmTB2QynA3hHe
UK8l7DKpf5NHmnMvPR899tc2m/9nNdxgA0ykx+JJm8v/Hnr3DwaWjzPLDEt6WmAX
IxrSjBihXS6in3hW4HMHA/cFqiTZl2b4zYzb5XWvpvtYPNBoHcrSqNjKJZrRaeLn
o9UUutySOZlt7OOgIRLuocBpf79luE/Rt6rSYH30KFMxUat4Xfsi2Y7pSW/7wgzf
DNfEKwfLXzzQo+fVQhyVh1w97VlDtHCOFVv00kzB/9Obvg+ipP4nRA32JQiW6X2Y
735BuAu5WnincaR7rVd6utcbhBti2kLfKDO1I2pslp9/J8g8X/JxECwkdACe12x8
ggqBrsHq4z0sQ3ClJKy7gs3aRl43zLQXhFEyKTV/TJnxdiQjV4vyqFEgobCLueyf
lQsWpvPJR9eURFixA32TIQpZgnz4+QfO6oJqbSey7QejAVa/e8kwju+vamteFTbr
Em1vVQtEEfq5yS68J9MB5o5cBll0kNz3NA/EupKe7OF79vXn2nw6Na9niteBWqPg
0OHx79EAyTexUvfvzo4FdIlRol/oyAfIszgxEB+ulWIxf0bRB8M5OSD3EYwZxWsL
k9MZZiXnVdeH3lYHIcI1jIxM37vcz2lWOupZJADTVD39XADepZsvHhNpn6/UD0OX
ufdR+yMRqm0TY6AP7gEthx2MsMGl8dmS6xliGjKrbIk3pl10QTFHa/OsQGHIaOuk
8HRM5dSh9J85/cLufs2SMYlTbh7vWVWtdon/N4zmVMLyf/OlY8y0iWl1JWUTGh8O
1kyZZtIsIkNV+RofNgjML3fKgcTcdN3uvKrhI0MDMvdLqUgsVkmnyral0b7YXOyT
bPT0og5qCFLHU6YJap1qvhfF88iKLaCEhRsTIolvagMj4Hm36m6GkFW2VSFuzGMf
msIQKYN93IxYrBTbnUYXMg2wJHUQG9sWb2guJYvbf5DJ0aAN6ekjDzi58S3HblCm
VqddF/UrYgrEBuvSwRrEU+kGL2/I7JZ/4wchkObL8cNEtHu0EPT1grSdUP3i7pDe
AIII7GiB3vKPWcN/2idACWFvbzc4HiMNH+qmyNkhkN1csqnAaECtDgcctwft3PjR
vFV7A0C8EMiTQudcv+C1dTZtO/wwCCxpW6kddNryOCzog9d8aUNVY2YmUNmcVKE1
gmcvJfXaT5e7wYischB78wWRligR/lcHNdz6om/njY9WgZmu7WeFP2yZ+YWNT36H
qZxeKxU7z5fSN5/cH5W1ul5o1J7nwqTvNS4eXwn69jz0HVfgcV3EtxcmYgfr0zlU
vaq5XCsQqKzgbtGBVg5qiGrVuP1uRpkui9zLBd/WLjDK5qdpQv2vZ+5qWO7K47/t
F1ayEctvu6b7lZcUTsD7oETlFXe923rMbHZ4MR03ccZ+FzX5Vhn3BKBJNmjEnosA
1Juosfq3/QUAWq5KhQ75Uz4f54im5WJdHT3l/Do6uuL3Mkt1Mxa11dbvtgkseXPQ
YggOSmhpUpurmhKfbyQN4WH+44+4MFTd4wPnjG0JbS4pAuQK7hC0/Tvgt8rt7r40
Ho/foyDqOrX3/b3KERhDjnfzK43MSHmuSsnQIWvWMoF/Vu6RSDOZQzgvmCWvVafL
/OFavHifKtbQ5/BUiwBja2K3n3EKuWAgMMRsHum/FZfjS31QjHgj6sC4DwfDiHS1
ostX0+dEH/kFM8FL6eSXW/M2pMU1+WfWAjTGbmqWKab2CCvygAt/RTchmVHdndIZ
2MwSB0/ltEhd5oYvcS7/tqjUyJJKXcX7qTRyjNQLoR19y0KOPS7n8JfRm7iNQyJb
Mf3zV7JZiqh2IIoowPYrgyXhH8j90owFaxvVQqmqIadlC01lxfjZOxjasrjTvjhy
LdTgGeOyiwcgP+X4XLN/Oe4rY7luTLSn0U1/WGa5A9HsWnR8KvVDKKRkNiiZkx3f
4HTm2NKOxxsJ19pdkHrIzurCo5NSK8gBYjqlDy6BTszv1wOSGTgMyw+qa+yz7vy4
8dLln4R5gkDVw/kigqVqBk4F0FoREO8Uv9eYk40j4TTMNoHYii9/MWtm1Fuvc2Jp
7W4uVS18+u2P6qAW8hAj8fcA+Avya2GK8J7D3/Hytj2eC5bDkXtgpQ9OxjjUyPXR
8L3njS/YathLUhs1oj5Fg1crVn4VnjwbRNzVy8Rn7pb/dLuj2XYEetMVt4lhHX5J
Ls15GWTGGQ9tuSXSzQarDJbQucmrfD3/BSNZE7sjljvLMnR1AQjaozlUG8UUhGdb
yF71ZVduPWA81n7KaBU6XdGuf0R6YDCdHHSdEdrs1+YBcHAsPT3vCKHagHWLnlHN
d13uXHYQn4I+ahWULUNV3LkMHjiS+eBrFcZ+qSvdSyKg7Fjc13BSyieZeshW2+Yl
D81AyNRCrazql9n9Du86XvpwIW9slvXUovIdf9dbXoegJDPJE1Delc8bLxo0QI0i
rTVAwPqKI8FrTlIihrMhvGakTF9oPDhVlkbwY3PtW7YVvOwQBcaQBZtTK4Zptinf
i9FDyJtMBzokLbmEcF+tC0PauB3VHMd9UQrx1KUSvlD4Rr2eXhuHr3AnzPEALRWo
eMLDwqPnRnaqqGLtJC0/Gjz/T7Oh4OD22gFeKWWd1a1ceryiGoUKT7ghBoWZDvNb
2Jf2MYaNpjM8+YDf2ZcJybv5+eEvIagvAlBiLa4234JVrr4CC7O1KGAtjbkrzzOS
0tDcJJBPpB7Eym+Ny/u4cXKcRV0Q68eQ6CEWbw6YAwflPfTBgBXB6eF5CEr0qmNs
Ra5iUj0hwXvGyA4EbrFhWO4r6K5FI4Q19GBy6dtRXPOs/aMIuc/4/0ybFuaGBo74
BUQmsg5Em59lcXgIeMBDiWgldOy6ocuNJ6GUpNIHo3h9kU6Ll00O9xL6OrM7n90C
VkOwUPt1Fzr2aW2XD+KAhoagYeZDtQs7L8sFgx6gD89R1c3OhxQVjRbbaxxZ2Z49
Ke4bg9WkU0H9KCPi1axzpymu7JhaaYuEflYm+cLjUf3/mDem0sOUyHLZ8hLsHOVA
T9RpArhdJSTJw97MdAKzhWSC0VEEooFGCupxx1J7tseGrQADl/UP+H7w88HJW786
udVIlEQJN8vze5X6jP4IToa0BI0ZLlX7xy1MLUT2E9MiAmm8Gj0EPHXcYvJdPYgG
FDzSxcYft/SsfW0RVTQzdMz0xY9mtlJa/H0VesH0uv4fJ0C0901NPhtH8zzC47vJ
VGfidNv80MTPin9zndMcBjh9fITmbvut11AhfD74Aqa8wWvsDOWUPNPZ4q5Ij5I8
Ky4FqamguDXQ65vEJ+KnQboMTqTbrla7oNCFVATRRiT4GJpninP+0vJmlFYqYc1v
H3pzq8aEFdqqYMRxTnSOk8aH4E5+VXG9x0YtOXUMcb2I0jI2w+KB3sL6pi79eNGI
N6xQwP5Zp5brlYU8o6+me0ucoHLHOQv23IivY30wsRhiDyuBfeP8zF4m5kP8Y7xL
0hBDisyzX7KZkVffiSYOn9WyUcFp6zGeZ/ZA8dXLiHPjfhubPezKVsGErpCHBIy7
X20PKe/zuFgz0zAbkYu3xs8l/2ILPSaS9wRpMvOhF+7IF2fW0hEU0X43VCfL9m3C
KCNY1MtnhtfnQNTLBk7H0R6S/waDMEOQsadb3Zdh+G0fIbp8TAzVtWBqdN8Y8BL7
Oq4lC55o0iq8YaS0xhiXwdJtEuktIvcZalUHZQCIJq3ZR2Dfad2YZbNrZYrrVnXc
jhFvEWWAhGOJyF8IgVuhtAnLpvnNzkeAsiib9NAaX/nh8JTNn+XRdnUFZ3XQLVPG
2Xh+Klg3QVLR6jC6/O/qDmA3lDGIXY6Lj3J6X+jsOdWpTsrXII6RPVdGeD8Fxqo5
pADUepvmhtJbYagDfsgKLJE8yJ29hoEBheDfjvbl4UGx+DA/eO6NgQ8X/tLXOP6F
CRnrzGJjb7Xzd54WwQ347o0bWKJXLZejO+Heh8d0HL3vKhW4YvW39Ri9aG9JFFOG
m+FH7lGWmmMnHs1nFv+rh8ah11kqg6ryLO78ZUAa0GrNV0SEhKpTWatnDeQdDazj
P4zsDv9ieIqtvAK+7EDJNOzbsOo6EHg0Y0+rpiszRUsp5lRmdo/6qlJRcLNHKmoA
T7ZW5Rhigo3gn0/iYdjdXhZlXSeKBKcTSkEKQFOsMy/mJ/ebvYSPvTYfO90LRKyc
zcfYpd9vqoG9RWzvt87Z8oRyeFPWus+6AFRhxlzW8FVcWu+Gn/R6NDv72vvIbCPo
GOGFAZ35/d+p/X2Af7FYYZ6wk9ufXufuK7GwSxvhm9M51imyCjgZhhBCEQFYq9dO
IerfaDeAfUHPBUVEtodLQ3naSPSS0nwPSvKEQ5J2Lf6jQ2LLMNygAhVNPT7v6k+q
GWXlpMoG2/XrayPepq8lQr/Bcc8wveqYPL+zCg7mW5P+Jwv0TVq3PQzcl1R5Xazx
aK8NCSE/cvjOLdZE2UaFGQFerqEwi2FFch+759KMaxon6pn2cN56t1JPyCnp6Kx8
+A4Dpr+YaTmjcmiT+ODsNie246fb9P601UHKUxTMYjHbfaWMlYuo7Ndginqnon65
R+QvyhCwpG5QiEwJLesZUs7yttAkeBOslG+gtqUtxP6VzqgrTCeqlnzsC+YMaVq4
P7JPw92GLDG018cycBJwINfjQRURk1HkluUlHK1WzSUHI0LoQwpL+JPP6ZHyOJ/d
1oBuYrS8NUjqZwPOUH//PuitBWtqj6StbWyQMTgXxT6iTKFfTJuBJ98p0l3dSEiR
8ZAGlSgzv+jdwFGmkTjX6/Tnnc4R9uKDK2woyqxYWb7V/ROxi0iDpah3+rQF3lC2
vyFDoXsEvR4fM5x1vg9MV9kryFEtaHXPQpyi22vV+6cnbvuQSy0U93FAET7AhY5P
LerHg+u9Rh0QqcZlE9bCwTRQ5i+wF8JbClxGbNiyptsFeNTD/bWR2RG0uu+UPiVA
W/G+k5MUpK7Weca6GNM2QjJGIVlv5tGL47csmVDNeELHb9stOQTznHyQdLhfGy6S
mBvy3ZLumo8KYnARgTYxya+76sGKarSgn/2IgIojq0QpBbzNtnw/Z8F7U1xt60XM
Q3FDnC07xMxb9+QjgpEI2BaogAvsGoBVmctIcmptqtPPgcn0882LlnxnTCBjMiSy
YvWJSDUELGe0ups7iyY9JEcpbZrva7/FtuwvuBVEquwUPlxLwbZ5HvnRgWLVNcPe
YgbqtB34ASvmgjslISqQhSZHbuU9yKnn5GP9ptLPCw7yW+o/qUyoLy0XbZ3uIy2M
8OnRLJlwbAaXACAy9UjaYKh/aAEqNqO2edkR6EiEKwU7OGit2kUtBC2qpR4KtIsH
8/RCOZZwKV6UYA0ZdMNkQ4KhZZ4VXOhqjAuzba7u4rI9i5FHrudJyl3/UaG7pJEw
7e5YntzqD9h93538sh+E5DY8IXfhvNEp6poSiPVTGl2NREfVvSya/m378w9qrJrD
/3HJPA1TnJlwcnbEgsXHU4mun1RayN+PBlGPym55MgNat7dzTjw+/4cTs9L384Mf
Vc6sz5z/pxftitd1PK8Lc114g2qP1ewcTnjvTLhpSuFxtknK4Wl4qPVi70RWYPH2
pc6jZPkxygTT1zo9AWv8idNjOF0XQV9xCRxhe0R0O/QIWi81w1xOYi8qEo+6o4Qw
q73hfJapWqazdxRVezk7t/dYPUulX64BNzlM2eJ+I5x2O6kUHHzOhQFdiyB2OO6a
Vld9Zv1znDKVB2obSwlvC+e9WTKChx5jFkDZYFiIWBio66h04PJ4c3aPYIppcgar
nTF0yrX6rVSlVIxixLMoLEIjO6xWyTQ3dHFgwOv+qdzPrQZBUvgn2MzOLCDITa7o
isIr5abOMnWnnd9UvppdvF9lzQ8jFb7XtMI0X1TV8pfKUEkqQ3M/6H9fGXtTTM3a
BTh0+vGCcroneedFe/CYBY0851JiRjmlkkuEZ17KHo1Yn6CopXO0QlEPneu+obwX
TDCw1JezgTaq+TrdE652f3myhJhhPvKj1DQ14fwIhgOTGFIO/T6v9P/VO+aonb1+
7ryneroCh+IV7JgFHk5yv9Ch/IW4CHluuvvxKzAqXLuci/N2ozYhBNZ8Na2GQKai
IbMXdYD0ovlMBwJuCbXy1dmtCDxqFYfIXKSbIhKdX/J+LaHy/8ImnnMUBARegxJ1
7o4hvjKNzTFwok7zJZKgk2CJAT4uLADMfoj6yZLaRx50qBZKs9RLQvzzVSffJnja
Ww190yG1OQ5qMCgkgsEh7wBnX+MLL8s4xDRHEpfNUCZKWo2nPUWkQPLIPQdf8pxW
yR7Ai2U4otmvlE/iFEwIz0smKOwgXoI6C3b3qH8HL3uCwsczt8oJ2SlTSWE8O+jk
brBiiRcS0r6xYTiubRZJL75351XgpAbK2euL9OrkS8mtHViP3dGwRL7U2gsl/mXy
sYZKfLjFQXtQykh504zrXS60VSIXGN+FA9reSS83K1KvruHusTWvZTOuGwaxPmP/
cCPoWjxK7XYGHMBuAP0NL8g40Yzpk4ZhJ3IIR7VZ+WtGX1HE/OpKWIXvC1ce3OY6
4k2S3RgnnR2UbUkuR9nuo8WYjGxmmcEPDaYH1JpILSKTt4kPOJ5B9ZSPHjqtp3Ej
uucpxaG2fqlkLDFSdXqhQCvtbbLHW7ue71z93iXFpmXJeIJiPq+rSPy0TcvdJ93J
ACnWc1c6PoT3ps+nnP9dB+C6UF94EC4IFZ5YGTu4awTbLy6CJhxrmqvYVaYNlME8
Nh5lHRSy6cSVJvSUu4OFDz1sFHn0YP5WuQ9NRG4UdrxNqnqeDRQIF2S2u5uD8Q9m
t0k1tVcx2ri+/dachZATG74Eogth0CG85cfPKsKSGT/qZI4jIwJ28y4F16CZEfwr
UZx53Zxi2x7NlYKW0x2YbiqkW8fNIsNb6uGqB7M8d1/9h6KiZklnq3NKaCsD9fRd
k5LtUA9j7rWdPeymli3tZMRnhuuo08wSlRN/52PMWZ1TqSSaRbT68oeDmYrVVs7i
FRSBdIDFdYF85zj1fGDPTR2plkr7ccUaNwyQn6eVFJnLh4xTP9mTDhzm05CIzTPO
Rx4zmjQqA2olFLNDtREIg7p/0eTqNrgIlERR9rDmFXvFjqOM9ZDQhOpXEfECiK2a
f4N08uMyaOsKI76vGLDVqwwaJ5HnlPH3VuvdMRLJpy2ZTJPxyi2nqISRcfyJ7REK
o0xu33h4Wy4wHKmMDcLvTgq3ZMoFles0MwROc5S8yRMCh6pzAiNxtj/EzVRwIEFK
wCfFLMFi/kSe1KDYFsAy66ldGPBXAOAQQjEeZ52bC33oX20l5LDK+adklvmRsiew
YlhnqgMqAv7AcBrAMmAbFFjRslMsOr2tNHXfmyzDOFElH9uBE63AhT8go66sLSAA
su/g3iYcKzZvc7Oe1QnUe2MMtJFyLV7pMXpT1MmKL0jUCBipSPzrNx3cawwAxU1h
hpXOku8MjbckTpQZVGseNYmxdXj3vR78qtzf904A/G5B1XPa5sApgvewTFfR51pM
NQLOYS3jk53DiTKAXUwXbMXYYCHMgHLU++uMjmekyOQYx611HLQ5bkoYbHELaYTJ
dSFL3/61FzukvXzR4fZntsAwuoYwM/WY0SS5tsEJv9bAiMcXVXgA3+Uc0HCTv/Zu
9Q2+K40N1iYnS+lTkHZ7wB8CowtQis0+S38qwf7RK/PnB6LyrodiAg83wR1SZhW2
GlEZ7DeUmBboNsEOy4n7F353caK8V2Jr+GJ/asRDNWNS/tRcP7M4MEUYK1inPB8t
XMUp1Kdb8yMCUNEexiCYAT6KdEi9/KZJqSS1BhQA4pfCyu9+6T1bhSHZdTjbI7g2
bNlljIpPxeGJl5NLWg14kZYpm9TBJiz5igFDpmhCt9xvQ43UKXYqonPyL0E8yf0i
ZkMjW1J0Qk5HZZ8v42CGL9TwwqoOrzfITuvRlRkJpJl9vE0TWsrTQcLYzV9yHL2n
fekBzCSF7RmRIR5c8mBA2e0bCNKoOIVc4p4hllWH3Rp6DcK9p9dl2PVWpm+8DZqh
98U6s/JrdWNTdhTXh6ufBftPA46Ax7eZFivlNzK3l1AJb1+58NbEFgoTbyba4o9a
EHm0oiCZht0UUlxQCOvRswRgKyIPRu2FVZdOhqSqt7gAOeKuxAaTL/xKs8QN+qkQ
rpIBOktqOxPXWbsn55c68T0OI9PTgm3hVt7atM4Xx28Z+pKFQih2vjIE9QaQ0ln+
dEDR8Q8zmg3MTGpEcNiwN/5J35ks02PjxCW/t32TyfYln4NYpYv5An3olXqd7lOU
aRbIUHLynisePipC5XHsoO/fFSX1fcuKwf1p3siLxn13VqjHAisWJQgeBVk5giMB
FgAMNyJ5fO5VG9pknMIdfY1OLi7Mg3/A/3xVn1G0EB00L2Ib0s9LAYCiM1PV6qoN
9Rc2/BYlVi/cDpTdVsb+0/pBkXNvfTFM4iiyLNRUUPOHrR8ue1OzxqcLVSPZisPv
q9+u0TuFFXUO3Qoa/ciizQ4oNc5TtiE/sVeIy+FCI1IpuFHcwmY3PuW+jTsSRLNE
2HhLQ838EYHl8yiOOKgx4KH2W/Ak7CGpw3z5gna4JUfVDzRkOJEBGzjDr4Hud0aK
ovn+CAuL6DKGqAYKwTF5mEzwAfQL6ibKxfvGPR7L8qTeGVB6OUsinwiv50144qD1
dcIJfozqaQq0GE/EQYKzoliuIkxy1OkZ2LhghInp1CNaj9CoWlPvVsMu6ojFsS1K
MmrprbxbZ8oftHsJjjuhUPHXZgseNPNyHixIIDNtUmiynKd3tGtCwQ92bFJWclwY
rS/X033EYlLU3SdPhu3IDFSREY6c8wQSjYiQZjfNLmZivk+5si1jlEylfYxWn4ef
ZZ1C0GyabP4Ywfdyps6sjRGmIT6/j3M/lPplit0EaZ+M2f+hSb4jQbyfRN8y+1fW
2RH9YjgODhYEPv8XCA+Icq6RbAXXMf7PG/Ph9AjIzjnQFgKaYbCN1dc/05UGWuXG
Mv3Vzh/BMXFvkthDViASxJZDWFEpv2UU3Yk++vGY0uYif1o07MmHd0eyKCejYxEO
fGDkqrXJDkKW6MqdgwMv7IaDQ2YFBr0x0ybXs8YGBsJ4y2YE1Jnk4LW9xxOi7PxW
kv7BX6YbkXxmiJ6OLFferSWGGCofwGwfiIdB9bsAwJk/97lJZ/SDah/PPSw8xowx
KUT8zcZw2KurgwJo6JhwOXnL1pgPHyUbS1ZitaE9rD9l2lkUG1BOfx6cXm/xRx7R
38QqTco4VN5edPRgi7bmbkoZkjVvqHBhdoqrJUJq0D6kELhW07Y66XrBODCdQA3Q
8dP5aqbIMl9XEyvGI+muaYbzR6VWeGK0eS9IEmS3XtP/R03s40n0DTH+vVoI0R/y
Pi05ZMq2h4sIRm7chSPkNOht+4oTnOcvw6ztVc6ckwFb4ROy4XglyQ47oNMT/e0v
/fs9J9VO33vfXZn/BE+h7hNVMLcuWn83MXk7FtdZmyfFkwgKgRB6wRqI3YS6xL3Y
X2j/xtHzlcl0Kg6Nq45dbt6VDt9Rlp8sohPH7Rv4bL0xfcGS/avXqWh3voU0p+FX
LEHGJvAM8Tgbhe8tvbZQgz0k1HCZZ/pZh5lD7PYTlGGm7eSQ5Kw6IY9c2uU4oZOR
NOg7I2lB2Oyva/y4OxZaQTY3hDWQ436Q8xVpp4MraqyMvVW3VSlwf7IWoExSjc7h
h5eFN4kUU1Mr0kdw2XQH0ayPUMjbBSRTcdn7+BqtE25Y24Ea9qJQqLjxLqxhaMJv
eoID2MAYiAnj8IcvnB1pqYuKmyWBbYHgiCMO8x+fxoYz0Tn718GhKSyknjMUCiRB
oAJWgf3C3PAHJMVOPrjkx37GOMvyoxlwmnh4sYmpCBw4lYZ1KQQW9MgLeMlmq6P2
YTy8J6JcglfmMpQckXZs+r6iGCLYti4OzKsHDTDhNaYt800M6h475PM74euZj1SK
XPfpbwsmsi2Q0Fh6j+BF12M2iBDYxrZ2s+AOs1UAqRXI7KG1HLGWP9KiTfmecTz+
D6MDIOKupTaCwR0XkRLH2ehShmB4BmsIVmvyeyFPJpnAA39SzSA0hYsdn5GUKGNN
MRivarUEiVBm+7ueqxalUflu9bGuHX0PbmNXgEWW5cnkVslzN0BWkB8YX3tN0Mta
4DebclHjZrJy1vkkrUvEAeGPdDwk5Pn+GOZqX92vc9TBLARgS1CyJbqhIYPBWqBW
nb9BS9NbTl2+Qotisq6vrbLO2V+MOJgcw4Lz7wUzSB46/FQndByfSaectOps9dJJ
qM7uDEFNG8jYmC3bCP+3S/DSGgr0HsBV6ti36vFxlJF2UZygoL1+3sRe9hRavfad
YW8REN1B4apbSu6i71pmqQO9VhCM1may5TdogHR0SsNCwkbAEB9UM9ZkTPTv7aTo
bd3UOPvu03xHzzm5vArjORZzg40alm5bjFy/VKwGay25e2+23mKRd2xIW1HFvZ0K
kLlql1g9sposZfOUeeNaT/iUb8QQO+fCrf3E0s2gup443GGwwbumaKhUIIFhqg3l
FPoEtztEAOPRII6Ei85u3h4a/CP4aLigr+UvQvZCto+iscrz0OW8Qlc3YHYis8at
YD0Y7+c1tuuq4tRyBXornJcQmaSioy6lXbkPzH3CniIq39BOL+ZMvpT8/niC5gix
i8PCV49EnK29l7zla91GmN6GRHMucSKVj7R7XoZQMiKYsJ9gp5Du5MkQyBo2Uv90
4cNb7F/qBUvoi8z+EqSLDjP8gA5WsLxhAriUX+C+f6QAEQ4wDKMJTBH2MblRFX7E
EZEVVbRCSYzKpp3G0We4QaBka24hE3SWIK81JI0zZLDJGD+ZjG0LN8R2aUxFMK0p
G/UrWhUSwQD+vmC3J3ytL+c+KZHugoBRQEl9y1uuFFhyuuXDlYVzg+N1Qd9Bk4Ow
ErDVyjY2sM4uq7C97ds2BZ6JUd3COhb/bxDCRtmbOS5Vg9+ukdQlfzssRQRLB0Sp
8znFX65kHqs5nrsOe3rriEibkOYBneTniwlEgb9CqcnNbv3bBpo7DMHCox++ylJg
VBQFbIK/fRqajVyLm6qzVMLISKP//tD8oXKQOzpo5TVS99Cm/L/LCb4bu34+mf9m
CFWh76FHwmW/l14rdalSARjonMQ+m3TheStmqHzHwB1nVo45HXbT+UFh9uy09iGU
N9ezck2YXdYkNGOn5/KtWgdc8xbNPGpeeIpKMIQ6EtffsVOxahfsjvBNOuOIWaMX
APsLHexFyTYnr1/B6qXPPcR1P24nx1uL8Ok+MbwLgOUl/p6LBp7Zy5SqiI/JqBtb
deu+saTNR9goUlAdf1Vuyvhmv6+Vzy8E9jxn3Dy18aq9zv2uKBnGVR62wtzYIMjL
XnMvT29flgvBLSvYyKKYq2EAW0O0nlL7/8fKsL+JbrKt2iPZMb2zlbpMtrb68+4v
Gu17dDE5MEWVAwtbRYwSKYADqBBxKjUsb82Y+iWem9t79zzoscpIqlc7q1owwvRC
cAiuHRzRGkwGEQJ/LWVzEn91OVwpeIzBtcHsbu0J/mQsfIutZj0+c9Uj1wjZivHY
i6GFTTr7OKgCi72b1qQHiS2KLQ3qR7CXla2dZBJDUHcMSg6RL4Gh+wpE4VnpMnFy
yDf1Ozmkteptm87anRU5SJunm6asubdkYT0RHw84dOfh5tQ82Wj90nBwOHXLRvRA
aP/qBbSk7xPzIXwrzGkKtFhjR9IYgmNZ7/b09Wu3ZVxbvdnqhmlt602lMnf9Q/lZ
xF5IZMHAtHA1l+FrVH+dldCCaLr3AUNuf577Xq/srXkrqYgkKF5DlA5q9z0L93xc
qWwTRSq52CkFcykOLPcmXqQIWNmbi69BjnG6nGLgbWj5qrfO78deeVOlR3NuLUs3
MK5ySky3V2rGtlTCSw0bZu9zNscHM6uhjQNgfFa96UK4r5fM1tNHoVw+Ts9uw7gB
8i52KUsL8wk8k+YU+gQcYm8mfBnHPaJOC+CB8nC6wd87ThZyjvsKF/7lb12Vv89h
AWkySBTnJ5kdm1+nVpZeEkR64L73QJGC7Surl5Hys43KksiEHdqaGQgpquM5lSKn
x35GIx7vp4bbf62qIyMLFBdptsrZ1w/YI+ers45v0o0qGR7ZtWHVdlfyJrOCJ0Zb
UjIVihTNpWAEwJtVHoL9NXSi2PoDQUAn3t+YT/GywZUyzmKBloTZSEuqBVTLTJRr
zMf921xAmLfvJRIyA/sNH5O1rWTNZ6g+5btpFUJmLSZF47hGsiegHo9/YheMf/Vi
1aTKQ8PB4SO/79pvY+STtyXQ7F8E0fKjT+XcB203yPWsMF2AWHU88V0AYcDq35V1
bUl/EPUEqbxRXGy84dOZ9+ZP9Ls9z25YRTmO1AWcEak8eOGqroiF46ArRBIBP47H
y95VgK0VBFmmBuTOJDiNQXSHV87gjj0/9VexggBvPUH4bk6f96oudVTPevtNFHfA
+RqW7jY7otymnteZjSRY4DKhIT+pSK3aQ8YFEz2vnK6e8emL31VoplCboFpjqIyW
VaRVKNnKGXfp9RH/ApZN9HH6gtfVOH2zJrF9R5RYxVmCl5g/ldhUhmUcNCDEHtPc
uabz79jwBWSRcSgQrRt4nWSPDs+efzXgK+jvKXiNO68oFIMcIZv2h+Ti9mPiX1LQ
g9IVu1gdiy2OYWRI+iZsfMzQMIWhG9MT1vJLrfPoXwsWPRGBX00kzu7N9ZkGmtgw
O6WYBCkaZqgreELfq4Ig0qWjt6L26Gbd+Y5ocIQww+MHMbYrUyF7DLZvc3QPsA/z
F0dC+3c4HV5vyvx2k72ld+Pzp5SHhlPmV39FrKLeq5WV/ybIZ3lGwolAl1FI6cNp
PXjlCqzE0i3ZEm0oLItHUsVKorjsc3cRUk0ZhlwQLbs0Tc23+s5rfuy4UUYKfWie
7kpNuCPIgYgrRH/bcvuCXmMpFeI8DkTltXyK4qnQdrzxt86lEItC/oevVK6Q7PjN
4u2e2+YHwgpPT/o1DVT7Lp6OYeCEeBje547pduPBFEW4gYVqBS4D3PMjsfV5Q1he
FOAIQMmM9ZSflm0Pq8gfq6vzm7ecePLMrzyBw6zTDUTMO1hB+OwOoKzTuPmXm2Wc
fBp4928VV09vxNA1/WXNN4Ym2IcV9UTKidCc9Xa6CJ6OvX8iXXQgZJeCPAqSWuFa
bCqcpuQ4nspuWWzmtremqA3TEiBymou9uPbIgHTv101M8XJtPXzUMU4XACVVNsQU
Hp+mQ8apG/n+rAwtoiX9ec1g5fQwl5GpFkZg+llpjXECxaTin2O+HDG4Ff4fwq/b
BVBu2IaL0fmby4mWlIvfH9nXWgHuVzRgE9wYXWa44+GeT5z5UUSPOa4yDnhM5cPM
btePkPq9xpVyBGfT7qZ6rxBqKKTBDqnJ3X1x4EL9CNOzzTDXD81XUQfN5R6DbM+J
VNkiuS8b9ynwBJ0icfOTelGPPWUfiFUZP7SMd42csovE2hTMBnXnVksLtwYSjaGQ
GmWyQowMSwJYsff+bFjycJgoCJOwYk5gSoAe+EYaPbTcjpPYnG/vDhHVdIXh4jnL
B3tu8Xok/TpPH1X8pN9/xeIPCQ4wq7dA4RHoR94msSr/DcYjYSY+uw6cM5X/ROv7
C10SA/W3jGklTWKkAN4pz3V9Uhkk/8FUWtJMy8fROldb/azgijNhXy7H47cWWKCq
2arFRYOmuLFiY6jfyJKbCkTYPfPkfKYHifhE3k8BVIi3hBUpzNwh2dEpvP997fbP
F0aCOgVzgtqAJOPmjwEovUbDCwocTlhZ7qsJGWe1ssuiA3xONWsFZPn3Bz/pOfVU
DmshKL49fzOVTX4+cQUmjebfXPXuY65zkY+n/Io11ZXu6oa0gXdNpknt46SLIpBt
UkpG05k/IKoslSBW869IJSvfqMhsxkHTDqHQEH+f3DQZZ67jQyuFjsp5GfsskbaV
QysAVCIIeZzXX7CYuWmkNVxFzjBh3n8gMv7cAH06UdpUmuJEMQPGwAUDzBBbvqVH
IHQd+rEtcHp9EhYrBpXZMNlg2+isbm+zHMDUxpxL4pDDP119xnikCUn5lXuh1hOa
ubYHN9/HZXXNLjavZ6mKab+FAKpAF3DQ/hjxU3T55uSFLddr8tO4h61EieDpwuLi
ZMqQp054QKepEAhVpBEHNUVgIWFXsK4RqD6xlIG1oRs1WgTBT0AjYQETs116ergz
5IR2ashJ2Bcr4AugdUA4Fz5pUjouPUFSHMfcDdyxJpMn+ocDNpSZDLo2PmF6UsPH
q8V4L7LCYStv5AcI718r4pb0JfRMss+svsor5GQZ2ZhikmxGSPoIFn8DKQiP92Id
IJlAsZ2JHf7IN/xWNbI6v4xksXvl5dihpzMvHqqJyeTwgDEaQn4iJrJ4uZuj+eI1
K8oB4YKrfpgm/kD9Wo8i13oLDi9cF20x/yYnI3Y+xWI7fL9+U72rzbj5Rb8J+kiL
dXWNy8SBsvpENKC3zsnyjzKjBpoDeeTAEpYK0ognc+B9fH6KCG7vKgj97YuiUuIw
Mtl0u2C2FN0+YFOUzl1c6oNfnZufYqMxFQSwkhn7W7M6WSjzMK8i+fZ0RK8bl1By
vVrj7GhRApE8b/z/2lXCh6oSZHZIuyd9amN+dFVEoDM7ozgYA3/Wdl3LTruOwDAF
IuYPwJMQROdjvW/MSlG26HUCY8BkeJsc0fRDVWVB2pLQ9VuCc69BjiZVZ+rgKpJf
8ZjnF9/qP7nrSDFOaMCCk2+ky3qxLV1aKRhPWqVPdU6Z72u65OanxetTzUCBn1/Q
qsQwqDU7Rpb3QyRwQa3w02DFRS0T72BwoCqZRrwdaCnV6bLWGQhAjqQxfPmB0LzA
3B00HJ5/RO7obFXw0kxO9WfIJJa4AHiBXWuj7ORO3vaAbyXBvznSrfwpG0I/sIVm
smQzfVdkSJPgaX+uLKC6Oy5XeH4tMAxkxJTGkYm9fdvxyOGsJ4saz4abAWJDdE8Z
UTqI9gQlko89v2HFtSlliuXxRA5Myi+1ZwNTLf+k3npxCGbX1B55TCEMeui4GQ9u
j7IYzePu7gtmTidAY74NzPXNcRbRNY6bcgg2gxckh5vWgr/BH1ZvB61eH7G0RUrU
Mn9zlYNkE+Fqy7Tfr82TpnClPqH41578sNDDAY7uj4rs9qdZz/Fg1vhcm4bEFhhi
4fnXrRuWTM4fh3pu1iJLEZOJ9YDRiM5HZQ1rdh27fU1kmlabqUkMNMAid05pvIR6
byGPJ7sAT1Iy0gs/QdPUWBad+35/FR3zWCLT7Qvt8M3xjVkqH8HVNWVKztSU/NDX
KXaUPr0oVrrkUw99Mrj7QgjfThhPkXd7rFaSpOgl0l5+hivHyN7rD6CKXj4QeTbG
euV2Rpl95FulpdfE4ljbFCyI1lfgKGKFOkffqrnzwFcxSALHblvaNyyV7SehH4Zv
OaDjyyWYKEhxBsnw0LP4F7jp6mBJaJEYK88Vhe4M/DcEn8p/pe5huUCAZafK6++n
dRM1ZV30BU/GB+izJWN3pQBxTE0yOgyOwBpUvV+ERzdFI7zs5/Lbbr+9RvDrQ32x
8Svwr2KtuM+Mdo22AkCI92PhrNIQuaD//MXHZ7smHkPjkSxb5VeA5m2ASToNxDeK
dyB3vh7Y3wtCbmgp6HMeqA9S8QCOs+WePdmqQ9vtEN1/k6mv2/ltW3jIAUYzRpkW
J1noHXSabnUYXsRYpVVEUkb1mgIKi9Jd4N+o1rTR+qj89e6AM1boLFEtd02V8lA8
4a3kVJgEzos7el0/sLrKi55bLoFZtBUPqnWGxkUnuDE0OjGz2hiuoDpDmq2UGJIC
AjCc5DHkrGfhN502xnyR82dYTAny7babFLT0nCeYMJIChKlbnDrhFz/xKHpDbuX+
5FU1g1aSTnkrI4Pk+vhNvsIC2vl4FLtK8QrXYsk1uQAoyP4qyRMBCOfy2SpWvRiJ
g0i4pITIFVYje77wCbv/eP26u1I/lOhkjBt21vcVK+zGD+oghykF5dNjw9XT9Yr6
yiue0y+hkQpx7DTcita9G43iEjp6CuQRRNbnDEL3jlNuQD05GA25Wvi9KnWNoLuA
N/9VZycWGAEp5t1SRBvBE1QzSIPadubRW2vzDbvCPPmi99LhjAqXApVmJnitXWRJ
cBKkqinXQhrFc2sMmx0+jxuKbXVBQXJVQ9dMKpA6Q0LzbibHKaNoqhC9Nhz0Jt7V
+MpazinnN0vUgdFGLbXM46uKjsihL4L75Ky9unUY7fBp2U2By0A8KH8EvuxCQFKd
rTtA+MSU3o00M9LtS3nyMZDfeiywwZEdpb1YINP2Mj0WCLGYANcq8Ioug80iiaj8
c7x9EarasbnpYOgLCHXNv/N/1x0QK3Sg1+p4Hg3aFLQunfAdau5nbNzyCL7vbeU6
+ACXoJsD5LVcEj48E9viiB/c1Cnhd/9L+Eb4QdNf0JiT5slugcfE9SFN3p+T8xTa
eRlhqo03652uHLvzTqRVGXXx1SzxSPIv2U7poMS8hL1alelBE6Nu4G3qv2518yR9
uxmGD3pCMSr0tpYe1FCp/FQzhdDqgijmWDwKvkbbErXT8YHh+emcxHRwNx/Yf7HG
WQ/s3i5TUf0Us5EuxU+8VnfP0N+OFhENGKzFo7NR4JZRFr2hF0gwLy8R38sMznTG
jsOPk90sT4gg2omSaqrpNKTkIpg3mPtdvy2KGmRylcz07nl7O0HMg7+17VOfnr7R
Lxj+NAvithFo5XAhUMz+c4vBM+HZCOERQzv1yR7xL7ZTysDPG1CBd8egs39PtT30
bIMmbDUxFySVw4wLbIa6RTj1mZB4oAnD8ejx2WFbtCAqoAFuPpHgFoEZBMrcAtNA
zQbgAa3/qkPryfPH/Dbn2e4gdave7cUXZiEsNWMWF8cOxMHZhPrqPVZWCYnNRd1b
SFIDFBkmF4GTOyMia0U/CKWqsd+thjYJk9355cWlLAmmf7pDKtgCix7ZGIYqtOHB
hxYpT2bBf08JD5FtCsjYNgcAuZ11IxZBVDt0b3Z8Zs1z21+7pPeO8m1u9oMyXKD7
OpxdDI1n5yu1p8zCAnJvfBehTfXRxyIbQqo2zvKqDG/Cn6rPyWR2BsR88bOuWJak
h5s+YK06jsnqkCxxpHDRia2Zf1YNslozBT656C2CRpunqyTLaIC1uULNcX87zdq/
68ETDOWy3GfQVK/00S5hO2NS+ss3GXbcyuN86tjxHuivm+wiNiVDoqyK6FN7z9hh
Ucpz7FScyJ0p8awsWzkU9ysE/6pHQf9klMdxv6NKZ6MjfX7fElGObYH8cVdU23dI
gCJ6oQSW/Gnyp6Ey003Wr9ZADJ74m8hH7CdKuvl6pPN0u2lXBY2YJfOIeQoYiPLl
UwTm+M0xmiKjF+snkt+hc/5Wqy9j8JLA5IfdBJkUV3C+9QNCRHvcEgsNAa0DW8hD
QU0iv2Ji8NABtR38OfNewLm+bUcKU/klfb3iiZ5wlMFC77QxHsOlOwuLG39YXFD/
vaH5JFExnpzwxnsiu3XGH8EKQIwwpf0s4Zw4/obJyCmj3JNbqikkDmV5iP7/oVuL
7c3rzIdedeuhRP1QRsdiUBC3P9ahvb2d284OITSWaVL8mGPvgtvov46N0opp8mU6
BD9MU2t2YSlCtXUj1+jAsrxDKiiVmh2W7Hnhx4GQTSFqvzaSSXFLeUv9aBPuPsIw
vI8hXQrcOP8pmsMOiv6KssYFN8ITRsVjYySFsQkUkY9p8+ITc3lO5bMsWCIJR7Mb
QMk0uoJ/12ZvgAS8ShdSaitdSdUpDIMQpJZtg1XsJzUbsOmX4/ziUqE0cceqESUT
6bmu84pk+qiW3HjojFRdjWy/MvWDFbVLPWjvusxOQ92QQbSeHNgAKipHWyCXeIWP
Ye8P1yo0t6VNEp+qhIR5RteBz+2tV6a1j+8Yj5VTmMfBI9DRRDZSvdAZoXhR101N
sLnaLwguikRgQG2gTzHB+yc8yJBRhidi0MS96tRmgSz1/+w+rmEbmY6TiDpCr1tV
EGROrmobj0YI9hFwhMkBwOrS6lPW0I69GCuCMFJkhLbyQJoPnnH6SeFO/TWSs7wZ
f8tAq04SpZjCGrD4HAKJh8irth5m4PzF2auKZyXkG47akxfleI4U+q9mvyptO1fE
1N0+tQpLMChcEQucnYGnJmJ6qr71UAxhuc1LDTxoShY0GfgXR05oy3VvNE6Jvfew
7fhnM3d0c+iuAV8sVCBX8t9KGSClX4REsZenL/2RUaw0WwpUMEmXYTzdKEdJRyup
+oK2nA5oKasmMPRLI1+ZUMJRnY1Vj6eMu9TnWieQjcBAGcT4mLZ7+nxZiU0j9oB/
wquNnA9d1rogd0L73x2pQgBtDhFeaBYZcDsJ9bUaf3QhkBfAJrwyUR6Jkg3KXGD7
RpzXKnIuQ4Vb+HfdaVNFsbDIgLO5tLcWqAXUjeT21TXRWqDTIFJtHacALliSt3Ab
DtzljsyscSrIhfqwBgxrnNaFq6A16+X81eczaQ9R7NE2JB57TvuDx0Am352Q46nV
eWlAdyw/FO7K3t6A80F57uj1IGxsadR3qozpphpH6fgJl4AurP4FCVpOqiavR7WP
w74vhG4NSrT0g/UHabccWE438DzjwVR65OaSnUFelQZguIGmvjQ+0DNzIZaO1YNp
FgtdnpGNOAsUq9+2q9aOYEYT/qxVcashXkpfkGNp6JAVeO0RoXQmtskWMRTDJjOq
vaogCyavzUfV/xkXM3LaY9O/IBjsZbyTOi4c6Shfgp3GFsXlfNzGhwU2Th/PD46B
3Haj3ALRd7Kf4Wj4oyt0fVYStqiG53hWnWls4zNroM1ZqeNccqQFjpTU/RFyyfSH
3uRd8uLf+uj2lxGbvm2KFL9PpUlaDs0O1hJFWmB9FDyih4XjMtCYHvY8LZxNc/n/
1EUC2WOrHi4eLQkrtT7h6H7+sb49bhV+iYz4EcBMwqwQdFtkSzaKKyVm5gRhPixX
ZCr/LvRHPcZvnbpC5VIqRb6ZAl1k2McCD/gpxDm37TBge6GBQ6MNCISVlVIY638l
ahP9/tWaN7KPiPQ3Ujngu96RbDLDprE2tV9auzdpiGtd/oxFMRTyiOrmPAXsOEKL
oPnJlZ49Fpp/MfBsJjkgTptOHCz/t/golu37WVZTGnrtLBv+M/3c3hS//IJpGYwQ
MIFq58LWWzvwUSn6kS5LYT6wfZzXC+TrgMt9gxaFrrXwRQxDehTZE3yclKjpEMwL
0rA/xPdj/ppRSmgum/iDYaUckFzguh5e5tbu4MXAQ1TajXwQ0HFagvWW5rDj/fok
euEv6XhqN11mYLbJ5PCAG7PVMEH6ZZemDO5zhhJnbxfVGSwAcuH708IKgOAQ16UW
7JQN2cZ9bSO+vgqtjdtjZFOmWiOlcB3/7A/DnPATA5Gjbrzmu1n9LkEM82AlbBoq
R+a5tvkUsqX0kMn0vFww1ipQ+VZAaIT64gHjk0VtTORGxT/Kws5joVSq+wUgl0cK
enMVCwu6H0jK2Vr/jBFus5lugWTnxFBKNsGPxOM8D9d2zrxg3hfP+8bD5iGSF5Lo
vESS/mLgz5Ce1ndSNPcRQQFLvv0/A2cPADBgNl1WCNqOgKuzn+QOQo1Mw2L31+To
KWnXficmUF3iihDUnqZ0tNqa9hKZjcunF81ENo0h6yGesoVpNQOcKs6q775TBcvm
G2Wwc7RsXIYnrVPNctJSYt8qb1AENh9i+v3jRa6TYeCLyzb1FTgQAjl3riMULItU
2caac0npmSWkWbyTs8EDjLqA5IOnLLzQ+u8LUbSpcP7uFizozE++1jI995V8IHzZ
AwwhMosFPpaelyFj8IMmoWpcIuuMF7JWdREa5I+X1SS6qF4ZCn9vDiMLx38FCZ4I
P72uPyCZxco2Ocg8b5bBJBs3d2mJ0cLjOYLj8d904KdY5cdaQNu8tMVrqhUuAnnm
U6yteS5rROhI3u4dOoS4eaanJeoLg/aSnPfmRuiuxZ+CNS6oJWfKnWrthmGR0aB2
HzCTz3mCbA+eYFjbljLw6sn7VoqVN86k9B8UcXp40AdmD0iSBgBDIJ2HfNpNclWB
PuD8VvgSJsidaHuunIHQe1DTpKUbZeuZa0wcVJPqlXUHKyvOwZrB8hZ7oddlLMDF
6mG0jiEnB0SIL0MFMA9zXzxheAIj+u+JgfPG/dLjULL12vrCRPyJ3yYB6vlwukgQ
zO99EFZy7RdHITphnEvhrVf9MP0RBl9PPy5FSHHAB4xvXP4LVaRTGO18YlWPkvWT
fW/3rprA1G7ghAW3hdup3XhJQdnfbY3+ZmPgAog4o9JgKh7Aptc1Ws2Plv/pNSy5
E/aCnfYqsgJ9FPmXdM3p9qTm8Q0qVbqLsW4ZaDyS6bEaTwDhEydxXXTMOuqY71d/
rP06oK6viepBfUvAGofNzmayTTbn81baHF2THZl7xsbOZBvxPQopNh+ZOZFSoUZh
stH4GzAJK/OmTCnCNbCHGM6rgjlluajJXtso4vdIxMEEo8sNECVZz7Rva2VDUdLD
mpziKHq1ecBMkW3g/xu1tvue/dwDlwqUu28bOZ8ZO6o/z4CLfQhABFYTq2w3aD/r
ov8zg8tN0+/BWL6l/LS5ev7eIK7z++DMyDD1IWwyK95FYa0l6HHlmUx+YlFhA8yr
5mPRSmGShmgY7iZ0tKuAIUqY1VZIdEkaJrub1MbGh87jtpvBYFnwSrpN2lmSJ76a
qbQgmPEmqbT7NcS76P9ESEMEthAipwWRnPhytLEzsKAkLEVTPECD1R93FrRQccbM
oQAUIX4Kci2lWWe7/edvZxvdfU/SGSndLSSknBYipeF3AGwZKrdrdqd4idxmcJpr
odhxzyzVdJ6FBsI3mUci6fGVc1D4XTTEOciIf0nU++KdvJkI28UCgaol841r/iu/
xpjgKu4iVq36tQTSxtlKnaqjCIKPxk82AvFFtYzJ5BDUJLi/UWb9dt2s4e8V8MU1
oC4JD/aqFykChxYPnYgOuBeiCbAt+4fgECASFJ9d1qCpQoD+XUlXJzgOJKhxT74w
WQc5stMJ+G0DIBdZlx0sGZvOjUKwxHJUHoqpyYRrrDu3dInt9OQdXhE776mEosY+
5IVleWsdAzojdKJMP6X0dEhUliVvgwkwsGH8GUrbs7myFdw+2Fs4WpdnpVLJcRwJ
WquhBhs3NO3lryfSdC8IhXzp19slVuRyAnciSEgx5UhMr6AyPrZDJ8hlCYVi5aIF
Xop5IMlCIQCBlOrymQHh/rbIZw3Si3LR5/QeRJIAlEKsDrlRMwZk3DYT1QgAXWQt
EmPnJ6teeB2tbpBekdCT6f6yT1kd01E+fBSJPl/eprFCbCyco6XKf9d2Z82/Tpq0
gE9FTqlioqPFkVRfbCzYF4gONP79BW84JuMUfAfJgbkCEKOrxfzeFY+TAMuUY951
4PGh/T9XLQRXx9TIBl/qF/emOv6m06hcgl15BNWTtKe4Z5aKJ3rs0JgtAGdLwxYf
eHiY+7CJ+e3MkKSWGsmV1sEuxK8bIXTLxv0LBLl6KHlier6aaNGs8ASZ8rMxQFsO
IjNfaa5Yyu62X8i1e7VyjthUW/CAx0B7nGM6CZG/fbcIY1Nd5knzbSQObYlxGNSc
XZG+jV7DlpfdJkwsNqFU4VUC9CcqrjozGOTYfMfOZdO4hzWLaALyiSVRHm6F3fmt
9iwtg3VrmP+G8e6UCWHogoCnaLl/eZgJkEYA7kicbDIVqKg/WJKlCrkRWJIm4f5n
kxW17ryrTjLd29Gutjqyc1pxkm/aFEc2XBlyoU/v3iHDh+N/kHCV871hceGQ6c+b
IBeG85IpF1Tpmw0gVjuBn3JPjfC9gOUki7O9NDIdW834vSW6QL2EIwiOsa8Y5TWE
1hKDr87X43MZD0zqxwinIIIhGKyzpWNDSB1uW++7gLJ41uLq52nEET2sa05ftyq7
jarLUozcpotvKmYqmyvDFm6mb/dBmmOUQuJICsbZgLYOE6SJ6t2tvrS4OQTnilRu
jIZH19CZTdgOyjuBj+NcRftaaETsjmR8GAyu2vCg4RI/ynjEvnf9M5QjPbhcSxDH
S8v62x4WhUHf4g+g/+qrFuV0dTIfhJUj14h79yYwepLKlcVZmbr9pg3bn7Qm/unu
mB9cQG12/FgcBPxHccIBfN49bq2ov+mPqSfhpGjOdWwI+j7H8bNqyx6Vr+Wx7c+o
zBYfL+Wa3vQPDghypg9L9CK7+bHRh+KajwgOQKLU3hx4TGsKOlnig9EwPQc4kCzi
lIzD6XzqpoqP1xl/WNlrVTX+caBua/z6SiibmZmUrd+xgQEblqAp2Q4OX7hhKzHE
GT2An2jclqW8RAcjBDFEcV5fUHYEiO/ZKVyGrMAZ7Dklb4Pgd4y0v2VM57cbxmth
Wl9nPD+uqNfR/fPtskWhP+q2L2RgXX2vZOWE4U0zyM+fQgl+vcSbjsRnlkJ78ub1
5KX3XXqiuPLYYqLlfA4moPVk3aYm0pN8Y6XH/coIz6kwEZ5VNQ5kYLD1rWqAb/ba
PJ71BFVo04OuXn3m1dLqXz2w5ei+0cm3xJcp3pAGYwRuiKWYGRarpbew70A0XNGF
iwTrhNYecV+dHMQf9w6BsyqcZDY5atX8R47M2IQJoXOZLepRtEMOMXhT93AFSLsf
hiZu/QXWoA28+yeqt1MLDLJJiyq7q5b/nIsQtlEXe+1HJ0y7g10+36nthAsvKxpA
4dvK+dEE9eWtAzIXuQn7onCP96NABBjDcDkQnXoS0Sddn+HavzOQYviMUL+t20ez
RauxF9l0lqi11agohVLRlVcrfnAcuWb5Wc0Qwazcoz/WvjrkDdlhZ/R5piqpZ46h
EWG5qhS5mnQm3JPj3fs3Lv0xe+1vOrIsKWcemtSDSbrZ236P8r7e6aRSi4w6EkXg
6U/fgMK58tERkGA7zvIyCV2TDIc9yD35hFO2uanBmT1Qe27WOlbx8gR15R/8Ihlv
HWKUOsbPpq4rzn/Bo3CSdF/MXQzGr8bhgCPmOTFhsmckTiZV6P2pnLHnqS0JTPvI
jJKX84hKveyTV8ulHxKT8ge4aNOq6ALzBMnEDzbqNcH7JBuoKxE7SF2A9iuD6VTC
u0mtQmyjQbCLOQPFN5Zx1gcQ4nUqb4nQwdgNDsU+Ha06WYIP1QP8aB+sn56jiJMH
OMOgas8DgkiysfL2BLrqzYkqjvqjX4c13elBa73hCLfoKGcW1aBtvWtewiN+UcHl
wiC+5zRD2yGe+j263fUcemMj+FUAOn/ZVPm0O8S7eJYrvG7z5XCYx5+c2szx2k18
tM+Dk6WsBzZKM5DHwf4uEGesHU2RlFpY7ukNf3E1LzqiMgjp7iNF/q8JWb4fkWTz
eDOuJraRukQSpe/bLObEuTRvFrULsgktzN6bAtf4Aflav5lGxo4rcADhLsmNdHQs
mF4IpsDGUEwYeopljMt3aHfCIosXwc7dQPWiOklc+uGO1jm4ZwpHKo1ak3oFPe2E
ktVM8Q4iraNXcz67xaHqhSWMpnt7/dA+gXvULc26j3rbgei6gDaCuS1WvnvMhN3f
3fPWDDlNusRNx+klRRXv1SnSLXLHzYAOWBA20UZnycqz1V0qvosR0B0RgIhm1mP+
3LuBm7IK/cCqMRS7eMdXu3WDT11pSaN1kBKp8Obyy4bPcbuNvTqHRefHM8Dvw6qb
Ep5EemMb/5gFbghbXUl/6gKo/5npoIhXXeqE+cMUbRxSmF38YzNAjNc7RthBJwCD
9scuz9m5FeT/aU63F6jHfDeYh7LcIiQ76d8X0T9hfUC5TEB9ckMFtCn1akcba5k+
+VwBVHa8P3q+qK6BtgOLET/ns1tloOpebUyDg0CPjoV+Oro4+MdygylvxQVvNRJJ
KeDJAvExx4xtbKHYPTYUlRGcIfK8QlQKuSAaPKgaRahSbiS2FHpSJm7AuSF1wcZp
scbfD78daqXaZJc00nWdDLKIx0M8sHFbe1oPFOcj4MdSUQ+2MjX2rNo/e20dVP74
FaJjrUeDv83qmybJtZjDq4uDXOD53GVig+OkOlfsC+P6JAumGw3J8Eq72GYlKC5L
0XsACSOMQUem1N6kc/RLawQElbglW4fzL8LKWfrAIEp5NKhdHPYsz//q0tRx/XVi
45gWjU16YSOcG3GpX9ZfOg0EoIxYJzO7uL0wU/PatFAx13jcEtZQOY/7cbOlO/1c
VZU8GkEytxOrNDCZl9l1Azkzad9Bnpd15hGBYmGvr9T+A8W7l+9p0VSCURddh3t/
FHxKgj55PE2tJ/BwP+9b4/+V1ONuzfxUmzuhAhdchCung+/zqswPMMb+rWEBfLDe
90qtjsJSwug03j59Hwnj7qrNPEO3neTgFI0s7HG83fPJ6HxWTG3AjpEf8vlBLTuJ
ENQKNyhtfTNH7Ksr+AoR1FBwYya90ORvZnyXd6Ecx9maefGu7yBDdTKVBBKao1M0
+2BsKWW5BRAkIdxz6kZN2ilDhTvFutQrwNsoh39a24F7I3SV8BhBDMDiHea+bGdH
rozRRFeRu6Cqgok6lRmISLucBBxHWU9u3J0sdfkj5qb1COaZJ+w4ClR22D3GUnyI
lZCUwb4PQf+YiFVdCNYoNF1FTFV2cKAXA3Cdsb8HFnGJ2cTS/SN0tMwR9KdhPlsq
Kz0zo/Jke3LiKEiztmnc6kk9G7OBxapabPakf7dLM3JS0H1FMaza3rKEjq/PFfuz
Bg9qB4hfEsXh/HMPFIC2TeGFWHVswRnqTwCv8VpwGieSyZ1aLSR/rJ+EJS0bmY8B
du5OybtuYLne4CLky2OgHkgEPMMsH4/F5/3tujqj6IYR+zeagHr+Ek/Rb4Tjl6lu
4fG/uXn0FNwsdgfFeOmTXw3FetLlpZW5TYbp8qsQ44J0tYf6hXqxpFu7rOqki1Dm
CdSrE3jt/smMBLqrFavHi0fM5sCnpd3P8ahbXKZLa1EqiMAxmZ9G27+YnQkly4g2
Ft+MDBDoKk0cg19V6bia9j/oqaoi4bQIZq0WdtEXN11QD0qJid96Z5OsnHkgJDip
esaJVgvthWL2wN3GJb7T2QKSESfTzKrHujcFSNKwRvaoQhWw2Yz/dioIKEBjOvqD
epXU7IxJLVhDi9IvbUrO3QJF/I8ibvXhAr8DWgO97XKCdS+vEoa//h1GMp5x3Fkg
IEGE2PYcn17zjYGoaDFjwPRRQE/ByVnSJpaSDbj+ewUUL8y8M0KM/UFVeERBufLn
zQdt2gH48XSg27Z3n+rFqICgRuN1VIrGlEXzmfpBYMTpKIXnjQroaG/sdD84b41j
qaBZ9wxXzyiS08iJmNpK1uckGjQDAvmKIenmMKH/ynr13XQ/0xUWrVi8JJlMi16j
IKK2ynFmVjFipyjVxnPoQfJ5fJrWko2KNSu94DUFzfteLN1r2PCoy91XjOp+GM5O
o6E4BkwolelgV+MpPNhlboKhFWWXf4WaAn0SIVYBF4wwF7zsID7FJtGSvmVsQ9GZ
jLWYncjCgOU1EQibzxxo0MTeQvUR4Y4MN8kR9N9tEdDSzM2l+EqkaBIx7TkUQFiT
2kxZVJpftlzg5ILgpFp8d7NTvQHFBNWgLJp7VIL2PCWe4mW0YE8dzvSopcZaJ9lg
TeEXg8m+mYDgzXCfe9hpqfpy5rb8UEeAKYZu8KSehUo4TJHfl2T+VgqR4xSgK3L5
ODb3pxEAQsV/dRdwohYDOEV1OIX42ONk0oQqG9YXzcpt6YwOD005+KlvWNBVzcm8
kXleM0eyEvW7JCYtBbfnGJeyZ4LAXQCJn670QiG6XaQpm7pgB5LRA5Gii2fMpKhc
N8XlU7YmM/bs/45Lj/+AM+iXX6TCLYdkGWVJqp1v6qvd2dlNE4BpnWa4b75kp4Ns
mr9lAMPL36GiepD6IEaEVVHRBlpwhaLZGk2BFIG14TF6G3N+8u7ZldD0mX9A4gvO
svXZLzDKoHwGbWFu2Hkc84wbp6bkx8IhzvAmZQ91xgvTQ2dyP2X+YrKqSk9Fq+mp
TzAzNE6Vq56WT45Pv/2hY95tg10NBW9/CqYtNdSis7olc/iJNAZnK+nHs3DG/Z4+
jndGM0MsKHqU52YKcoYH2Xw8VKW6oJGUJvd/WRfCgU7VAX6E7494/2cynO9bYshr
TGA7Bn8bWCfMX+7S5KvCuLcGjtoWacU/Ghr4E69YESJwyjpjNMt3gsLlvuRHpLm3
29Sn+Ls01CUcNjBmA1Bvsc2Q10mAPBA26PvlJMn0OOgTXlzQZsP/jiOLL3JP/On8
xiG/tk9eH1NRZvU11n7uAWSKQ1NM3uLq03bRPmiBipiRhMyW+xsIMDOju0a/xRxg
YIvJAkzsLOOaoA7E0YdZmYn1QdWwQFbP1JeokCH2akxnb4YIlIKM77Ko6yAFsLcV
5ULhc3kdr055e0jdQF4oHUwWHmkqNAOjhzMo6Bm+CwKRxfprtBiYpRR0QnY4rAU5
Ck3jOj9/4U0iaw6Fdb5EBOCbspmOsTs4r7OqUrws2EDtjI4Gp5f20eB6tV8BYn9d
bx7G5BDnSwV5I1x3Kooq3AGvw0tEUxuakoM0lXxkXEhsCTY+iJJwjkywV+/Emzn5
ugvJBgYfJ9K6bRcbYNucVm55EqDf/UTOR5ELc7eprOAuxEozvKBMVGNnmzrTcwKg
J/dMSLSB29IxZhqmoiGJFEaDPNH3EcH7/gd2IYeosGdFuc8jo5OsWXbIxya18gqK
EYr6b7IJ8R6mhHtuGBvKSEXREC0jszyKGsHusqGZC4v3pveKWvNY7ymyn1ATMiCv
oE5zE19kdFcla0JgG64dz67tsSdTcoHQTdzxdIuC6N5wC2iSDDmSDMMAkhFo7OXb
4Pf6gHnsHP0kvCdHrbRtNR8zcxFUMlhqpgixnpa5FR2+srTMwIQxB+oyhxk5LJsQ
4J0ayBYVLwWk/aDG/L7E8bYnG/VpkLnj355a0L/V5rTrdD3GMrmc4J9KQ4dRsJ3B
ieeg9hjQ13vOP5+BO7mV+kigECo+CQUQ6rWzrEhSfgdDo4OYPEVNvw6VNwAuZtbR
BxwZ8lHKm+ApqR1FvemvutgYvRIpaHF5K7wu7WuIr0QTRoCLvbsvQw08thtYQgTx
t0zTLMsWEdQa4OQcJdWFJYF/WBQs57OBjGXvNzywobL7a9DqCjOwIKbKpxGUmiEW
gLLxFIrn9zaZvj/C0sG/3jWJAWbNLJunaLsNKhC1Q40USiW8ljSArs0/1CZITAqO
PKAT5IpVbOBaPzF5szpc7Z2HOns/+vJXCMGOLaewzhGZYqT+CDwTvO8NmkpkIif0
u+w6DJAXGnFRHC+jdB+dUUg9DmvouBoUvMP6Cq1VlQ4Yb8HHQWRDbihW7nemHCtR
Ezr4rBGgQztgstzxC+RVQngMlFohqfSlRGL6aXCODCk0lo3cSGi6iMKWYEn4E88W
QHmQ65zVbCuMZSOWksP81jj+ioN5FF3G4U0u/CcSnU4Uwih8yWFM+mH7wXZoC0x6
XDH5G92iHQ5f4mRQFwzisfXssUmiMpsfvyNryHrYeOKjmR8eaTpnGQ8mSNNKCy22
LlvbcZW6RD7uAw8rkyaK3pI6eszHrlWRzDzbJ7vZltFJx9fNNJN04ARDDQzJRktO
Tl8OTogbAgQsL7e+vfkH0+IHBrFmj3xj3hnRAjjLj1BLnoFtBDxw5okssXo8A6si
V/Dl58T1gPOQpktPBIkxLd+6QNAoV6iqmRh8FNJRnVo0GToU+N4xXh5GzDCjIr+s
twJ+jcHc5fX+YLwxfK5p4ijWCov8Gw89RPs2iaLcM5pdl237OV3ygx1mNauBBBvq
N3r7VHdgzJdcaYfBcN/f9eC6TKQ0UgVBvbYMWw+dj+IseFpneZ9Vw0rWyZ5X5jym
Hz3DS/MdMHIIJmK3/t1QVBgVjezuPj0EJLHOsNaYhm3bmmME0o00spnTXlRQ8NEz
PXRwLHF1I4Wsk3yZMMVzDtFapYoQOIdXiYhHXkMi0HHTM7BBYVcV7EDNykeeT248
zA9SF+J1J0f9oI+Zk8ukwcvTSYZHOwHFiVXBAgOTzXyUN7LfZJQS02cbarXwndLr
pzGU/bs4448zGN4w9cJPTDFKQHjuqOrBb8UuuDqznecRdRrMvc3TcGfP9PjSedlr
93oeLix5zq8zBaJZXL4Kx69n1AQl7VKS64VR26MdtbW/tY7oMFKqrNxnBkOU7C8x
mQoSk40ySwXXh+nuP9z/ddXsTgL0dN56zZvWSebkFUUz7BDbjnTbq6ZhM71QI9Wi
mbuAJl7BCqXH8uj+ri5lHMoc1XCnXMP0NR6uDd/YusbAY6XMtvDrzyrzOw03C1lT
u1DiXu3AvjgaARuj4g0s33iU31IkWSYZNaFzwy1kRCBQXvMpOrIZFdxS1JGDn0/K
WHpFrkwmaGODkNeHnHVaALAea1J+96WRNiUa/GDdaMc=
//pragma protect end_data_block
//pragma protect digest_block
em3l3Zx7KG2WfhZRsw/0/mfyXcY=
//pragma protect end_digest_block
//pragma protect end_protected
