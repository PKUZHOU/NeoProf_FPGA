// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
hiGGDqk++WByAII+jbgwTPAdB1i80etgGSflOmzeWN1KOBElIyMel0AKx5arcMaB2TvdpBEOX5Bq
eTd/CsaJXXNFTp3+iKWfuS1gC1LfrYE61uA1wLMUfSiZpI3UgVIZngatMF4wR0gRXVRZ7hbT1NMx
Eojws/NOBdDBGcD7rrX9qOfaFRfp7m/9FXUOqaTo/RfSuOYHEDB+7ygs2cNpLS3FaIdxbK93UmrK
QHBx/PJZevjbhL5LOajgzTMEhWeAfva/09j+BojOvexTOCHKRczgSJrgfWX8xTNhreugDRlk/Acx
sW2yWHGhzovKpVjo22h8JAuNr6+aqVYGeFV5cQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 3952)
Vc3JNUtlnKiKTflsRv36KOpHefoaGjlhi2Ri6rd71tjx+yEWFJnnUMuSSeyAc6719+Y39Y5V0i5q
W9jiqYl6mjL4JrgFY5mtCI0rRsLN5D9MhwFvy54H6X+qGn57BFK0L3BYdPjqze9p1fFZ7DLe4BpB
rQU6EcPCrQdflblBIF1+bq16ur4wXLk7uX/JkQK236FfsrV4U5Q6C6AHo7oX5hs5x/zz5jEMZPcN
nhdTZYsQg2geUuW++u36OH7Dvtm1hS2YdUbjwmgQw8i6hUVrx4ZiB/eVguNMjy3nBe76yhlA5Sdp
Kig+KwDJ5WSoIA+d7olamn7xcpOO4kr2LssKKCfvvXre0u7Ao0ChSKD8tXJlR/rB7crd8LP9zw9Q
zw3O4stasFMVnu+bByDoauUMAeYxkkowy5DeWoll7JTridurGXC5qi9JVZ8B3Tum8XgodFqy4cji
8Vqve2QNDh245eZ2SMWnIE2+0Ug14C1aiyqddeYzReGG/V3GLKdETYGMmfzP+XYQtJx1+b2tkO6D
PKaBZuMAyvRsjqPq4pNgJzm2jsQ6gKL2UlljRoAU825EI/kqkIlK6K14ey92qf1SO4svmMQzFRI5
ypFZMaIMJqRfUvhkMtTyVTIs1sQojCiZvv4GzD77MWFt1DjAfmeLfhh6ThRZtIy6V7hhvzOg2x5D
g0i30k23bhiqhQy3aaBiumeV2byrT2FbDkwa9LedztJ8MW58reJ1kcZ3DMtI95RBFkh1nu5bt6Lc
aEG8M+nSdR8BuTLoojABCfOwMsUb+HdZn2HJGRnICENpz5n+TiCifMc6WZdXo3EbNHu+GRX1XS/c
rUhPig7iDd34lmaVY0kXYkMWvWHuuvF00K2KDa/ZapMF96crJYY3AfQSBJ+9cKWXq4ZIpijOT2U0
yxtx+WVF3htvULe4MKAmi0bjGjMIUvwhPepjss+q3w8crSxODT70cmsVjidYv+qB4xq1DpTPOY5J
CFlMQ3OByHddA7h6uT8Xbf3j8kAYZzxBLPaVvc1dR02xnirpv50zySGlnF6+fVNt22jy/7g0H79I
swo4AuR0aGdq49LmGKBFFuf5nrhPcu+nkbmo5gtIKismO6E43nYIoSXKOEqVXWADzXs5K3Jk+OoQ
czuBaHotaU9jCLzWiEP1SEib4DpXSNZoTV3orCrjSEqBBaNqbTt89Gx8GVeyR2UcCF8L1fjcqRlX
p+mqEotOtjSpTOcdBajuvs3exs60OWqI58EEiKBDG3D8NRJI0fEpqNWzp5WFoiS5f7S4w6ZAl1hq
rCD3k2Q/+AAUFSuoIhpgAQA2OPaLP5kTlxTpH009oZetOouKXak0YRh23DXbrLMWi5j0HAa6gYVW
Fr4lNNvMHrjyWZcwrH8TOL3c5VJy7Slr6aEXll/295pqu4whCkAzJIY2m5Lq1ctu1ELjhulZl8Ox
zp3WXjKMUqymZaBORoMw277k7wJoAKyNP4ArndsSJj8o1eD1Rhx8ZIYYIoWxtWGzSsNbxWtlGjZI
QKXwpv6EFBHB00VJXzCgF5n5mm7eDGd8Jb1NSN+yBEoiQkfKP+HElixPdNSD1NYzO53mjVHOKwYJ
jLZvTofl3jeEO38qHVGYrA1wD9Ee8FZ6kq2i/MFjrxgCPxeNHdtEI1BSsOjruJy0LsfHFbNJqxAV
0sJtjkTQM8kYvhANwA6nOcCsdFGC0373oUsAD/jjN8Ym1KBGqvhMRWI5kGw1nGWra0eCt7a/qMX/
a5DdK/nyHypGA28IiU3gtjHiqEjADT4wNlJDZgAnXIVUKiZp3SdSauWkLSjZsuWqHSYZlPcL4tu+
X8nqR35MbJ7LLlRlki5V+ptY0OdFPHXnx9XPFiP/r+Js7GcX5uO930bnoAjvZXe7eoCoygtc4hlJ
QwWeqDrmtHvg+VVVkSapzS1pnkW8zkBjCVT2B7Knz/P3YHjNMAi0wry5UYA59fqGQsUBFjdOA+v7
lGuYGPLSHa+szxfeekNpBQqevUJEZwxxDj/WWOXl1qtJSUicm5J9n+YtVz7tBeXIkr/TtDOmSIGX
o6iPLb2edQNoJe5worV3kjEbylKHhdKehvV8fOnpbVdh+1WUwJFUb/KIlhJJ70dFEcn1Fvz/SpCp
lvZYjYu4NyWu7Ee+QkmdRw+1i/sDvwBKUq7/dvDuxX1HZL8WVG3hHHgDJTW2M2YLV1sa0rRiLoEF
SzfiDAZUZAr/vUBxPaarqQOTsRoZtHMxJjK9YN5BFnqVp4r2769nY+UB/o4yB+a6hRnmYmhhL1rn
CWZXWM43Hmd2TZcaNMB3mjQeAO9lktzW+zfpFrPdj1ya1PHatZgwd7Y+5cDAVl/tHJ8TRqmA5+Sv
HkVkNGG3vQQr5Lb4zO/0VBuJsa1X9WXi1AD07+2aOqu6/rclShQdoOJWNV2jrF3sTmMyUtL8p0wy
2uwKNHsp4owZyDyRkTsPH5Fx5dCBTBJ5dBbVlMoeodYX7k/NEtDsY2banoCglzPKV8kDGrWk9+Qd
+zHo1ryold/sN9hTcG9/4KnLm6wreAANdT3Dts45c/3/7Mzj7RJFujtd4fc+83WjAi90X6Ms/YOp
wwO0p9Z2zOWWJsQbISVLcYnL8GjSjuv08Cdbq4JuqtfB46Nb5f3bucqoqB0jcidW+gYxGMlUSE/c
fD1AeUuPfVqiqvSCEazW83dKXSOK8ZsilmifLTh02bDma6n6ggJZWfE2NHRpwUjEboMDZtET1bvS
Wpgsyo7TPKeGkJBFjty0A4jNP0bvDKQth6kkZV+LrAJq/Kl0HETuVo0d4hqkNxUdDhv0S6LLlzDS
dRevr4CHsyaxFJS2cyrtvXY1QoSJp2NPGylayoLGuMKjaFhXxBzl8vjUP0NCTP/CtauBp2y7K3W2
Nw4Qx77WCnlAiv8NIF9CQCVwDA4Kwc6UNS9ERxAie3EAC63YnWQi/IBYNZqXMswG/RyN+hzrDSvc
72lsaj9I3kgr9A4alkAC9/YV2gHybqxAhpPULpjJ3hi5YZPQNhx6Dgf5P/znLLJuRPq8I0dRKlhA
UteCkbVOvJvr/ML5MV5PLSn/eGrnTPoIqWqbWZ0XqvTQ+AX0CAOJ/iiJje6SPCRo0eaPiZWoKTE2
APkU5tQAdQ2IUqfb/81geX5SXJQBiIt3a+HPNvwnpk1BbFwpYPz88pQTSHiY1p02SQDPZ6UPLi+v
J2eQG+D6v6f6gOVrvLjCkReoynj3VQej1clNvTX2mEOT7nepZ1xFY0DZS3gTBtJSlLZtRA79NPDw
BoaQxm1ktakpoRdSy7o6IGL+iHVxpv23uJpIIWb870Aet3ftwy8U9+6zLxBTAjfD3pQZ2/n5/V7U
ndosLPZxhfX8OS83xta+Bp4rwuf2D4QIH9VMNcOtqQby2U7iTF+AOy3VLpfVVs4rhx4xmuAmPXlD
jSygw7XdbVgGtCl4JS0kF0PjVP5uevdAxYiuJbbPmSdmK60pHmo06Ccelz8DpIMswDR/Wr8Z2qiO
DCKXQPNp8UXHQHY1QNLX+EHBBvmIRpUMAdKz4nQPfTGqwK696Uyi1vksa4LmfKObwwHAa1ekggH3
wPBXWeQXdpuPVtx8U8lXTESy6uGngF8Non0yE0R60S1L/0Gz7ZtrLJUtDxUOm1t1a2FU8mkuizZ9
GRAUznEcu50gQ8KQtrF+oO3GmUiHRnQ4hLKHXRnsEp31jqyzcTFKpaPL4JSG4c5P8PD5tiz6mGjb
KSbXx5MlvOE69gV7eVluGKqGnLlpebn0F4qP3NWqOIFIu4IIUnlSslZIW8Qr7nP0cOZ17DPlcFcP
4/w2+zcxYpmh1oKDl054VT/L+I7zCIS7BsB6lowPF/1BGxgUskGeiLaLbWwDbxvddITHvHXxB9lU
Z1c+jaQxuNyV5pl34/p25UZERKdGIWy4WEmrbQVS34zEFEXuqhPQuSiKqhKM96xfCCOaMaUU1pxK
9kQQmMva84/59rCRGjxlA97yJ924c1/bDu9P/eRHv9P9Rmne6K/fIUj01X+rXc/fIlN2IHCfjJrF
7LDobrM4jCimKYrtT4M67qppWDP89PxenNSlZNdQ/coRtp2GEnZJy/YP8EUjF+ytKos9YFffqvWF
zDu/TeohY7kSoOnKhS193M0shGHif6gHiso29ZjMZ5mE/cMeXYj4fQK59P+xzIgHhWl0bUPF40uq
VALLjDHX/zE0aa76LViD/M78+3+q4FsjAY5TN0aGR77MDd5iWBQ53RBluOCRogQB+3a48xALTY7b
VSDWEm5FyKBp7xHM3EEcTArFJc4D9p3XL/cOl9bHoTXViF8Wwvy47TaFzBKDChjtVRNblwCJ9htm
+BiTg+E5IIy9kwfYxO4tTaE4Dhc+hhhhCBnapN8T36RZee2eTJm+LoM1jccNTtB5ZISD8jCp3BpT
+0jAcLjszgZHSUUXLGbnoaq/ZSFqlBRnkfMKEmSUgknyOsAL6IuvURnvoRuwtyP/2Fd62D/wKxtV
oXaLawoZzEs9gdgcawD0bShOQzLWIkLRRZryFWJWp/GyuCVWOLs69U2c6rmTGgnTxU05ZO9d9lnZ
wrSCBAC+xq3CZDwYeBV1fjEZg6REkjPpeeQmjtNWCeukGe1xc3Kh2bEb3J/+3qa52oGEJW7pRBxs
DWJBHZBkz4i3F26KuHHJYkaqn/r0SYTtA7uMbg8Mw1/2l6ShKIRhPD7hHVTiQyLiflwjVZ60Wxp1
mVOammmjNXxbvbQzgrqZLzaAbP2qMT8YZpPMzyuLSwO2enxDDeTJARQO+fqvzWkiTGLCce1omiWJ
MrCNufQR+wW1VsQXOv4dq+UFed04a24AGQHpA0FA7ZFw5YsAQdCEvg9DIMA0uGc72cQo9ThEKNOe
aoXSlfhBK3c7YbSaRUGzHP9qB06QfRfEpTYAP//wh53Z/9gwus9tG/ZhYMDBrJ7GPjh7CBMAMQE4
9hwBpJ2cp+ohTp7Df/YkMyBQJmxWUlpisgbKgoalvMqOi95YaIemwhXDmIFUQxjZTglg1WID+nbY
EyO21tWkEXmSOYUMxUsYoX3uYLI6Fh3YRXCbcgIlEMiQZ5b0cPSdAtDr7RX9YJZ07LDCg8p6POsg
yXeiC0alNSe7fGEaLDkYLZYYNP0UVHL/hyr5aGXcMJ97ghrG7rNZ3OXIDWyn1kKLkFj123SIkdi2
+cVkhBkQTSj0owP24qxOfK8AjUu5U9BirD5kxWLfwxukGtatorz2r7SeRH8moV8HLs6kYlwiMkDP
jmh9zvlq7ZdvDkO9EctyAaSUIQ==
`pragma protect end_protected
