`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
WBkCnVFI0NtW8I4jvQGTo3Kx7TAH9ddaG1nrROdLswl825x9JAFX1l5YPKrsAggP
tUZQIycTLy83MQ9N2RDcyOnrT0xcI2mwubgHGmA1LYgkPGjloD1Svc9wHsF+YIni
qENkI1/HsfMhshfa262TZKMFHXYPs3eqlDcWYde6jUI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 25808), data_block
8QgLGjrGndvnlPshnopuEW3EzixRX2LLNCyr9ln3yvxjWO1Sl1PoMiBqjkWK5Y7g
XOfyfaG/lQc47VLrIvu3JiYBiNnnUjhHWSKIMk3lZ7ZxLd5wegoXGqxZrP6pCAGc
r4KAwGKP5yaXt0CJKLnJ6R1teHRrQs1wNjo937g5tPNSFqHbvDBPwkuYy0ioqLyy
iWi5Kvx8vGWv6kKUjJSXlbzID7SWySFbkoIC33mRNsTrbYI7/TdOMnPblIfw9IeD
MZMIMjjoVHOCCsG9mv6HxOccVfzNnQ1XZ1jwpTalxET7Y4wQXYYQw9f3Qjq36zKY
lbtZeEDCCLU1ESqhuyFQux3T92MjWc4g8nENE6n8uxDT0Vo25/LN8pjSUq2w3LV4
aIe7/+Wf/tKNOg4NybBe4Oe7tR1+vDXx6SJI9rUWtTyRPneEyMkT6TWINaAbogJo
3pUBAjapqk6f6BBdO888qkQ5+GS/rOPQjAQQRpwS77JyYIpgqiY0n/gWkib0RTUC
1yNYXwTXAN/HrbJT08m9P5cI6cUDXj6YOI2hZiilOBlMY6sHsxK++Ky5kiyF1hkj
dxA2an9QXiFLlvAb2O+8FZnBjIVVPZX/AhPwp/BzHikP4vIbBRxePVsZDKuk68Q7
tlPDypl7VgV31c8LKV3JCgAvO6heycDicb6kx155KJpFAtMHUOZUOJxyq82ooJlU
hoItYUMO201irls5oKiu56sx3STZgjzhWUY/KheMxr80k9l/Ki5mg1gQYYsl4EHe
67omEw6hVrfYdoiRrsw4rcCOsFxTdhOR/A+XByt70o/pYPlpPNsGUnUgjOD5IdYx
q3EkG033ymDvbvB5NnyGjZEOqkhOghYwpqAo8d2A1dPTaZ+zve/rNXHGLwvgrVGK
tpxiBLWOwfhvn1ldVpdEsprAJxA4+/hQLPRSxdMwt6c+RIFMXEwANjYrCHljVvuA
l6ZSs6Gxm50WqVxIbElEx/NNYzsgufp1R3dtQ79wi5JFpEYo8GRzuQCMbBNAwrvc
4+2SpINyq/GyFihfr/4dK3Yp8ERcTGKC5mWF5kXgy2RmpDuykB9oDknLpaPD286b
hYzNNOVvQ/rQO4yj5Bp7WNh+1+EC6Xvzo9sXdHbpiFjM0BqL2qSL7qhYnQBv+yAS
6mqc7O8s952lmfaRIJQcIBv89rmqBYT54LNW16d0KWh1TFBaFhpR4a9BnefdIDyp
Ky9z2OzsXrJj5g5dXg0uufMTvnRs/NjxLtLGlIDA+Gzvzgg5OISaVZ2sWoILgPn+
hBfZZsr2HXpE5i4GSszR7DvrSPT2STxglFf4vmsG9GTllWonbMoYsIgZZC4olAW5
pEBhejQLrWIj4sQdFkrT3OkQKHkUPx9Zuwx5S2I65tb7YOSAS3GnVlcmKTpjni+a
5pDHDXKLA0n6ADbnDsptUrEfVM5l+lDjGUjijpES/nvcOz7iMaQnUxic5tDlS62K
9ZEw433Jb+v5hszzenAT57RJuRDim0UHmcp2X8sQsC1ltK/f6swES0ONDsAR4kki
WuSSWkm+/p4OIwcYfSRb0VDa7MX6EPAo8gD9MwfwvobE0J54ST0mFVcFl1+ljBb9
Gu5OWciQh715Co4PAOfAi+TiU34V05H4HAqs2DwNVnHSN7jvZNhRTN0TKA+KR3IR
COnwJaiyRG4BpAnY+HTWgQICY+EotNPReYhy8MPk+MuuhoJ5pP03HsvxDNxz0QXz
3lRA4IBCZeRgT7CAY/hTa372vA3jP1GM3CYDa0/6nH07ztB0K4OaLNusBttd6cze
tL+ApCMaZOPAKqLQwlq8uNjBR6aBbzH374BIB2qChTLtQkO7egpC/qwhiFAuhwf4
uMyBKKt++A5l0uyqJqO5GOAkXT4n6FdH/Nijp0EWdll1pc2W37/KmTvt2Qg4tCs8
h3k7uZzXcZbo/ggyJOv0lLm1kmF0QgCINeTxRcX8qie1Ei6N8ZilQ++qJ0F1QOls
EdZ58VYcAHPm3ByI/DuB6OHNaiG1XSMZGAjSV0vyBZjKaKCkHCewINbOXfBAfS/O
lgTOjcTn7MnST/6zD6gkzQ7jhUtAyLZuEGRObg02Sy4KrphbEAUVsUo1Ylb1QZhM
1Yt3SU+hNMffHS4UprGIKma9HpJhg7letGVA5e/lataHvAq1Oe2FBapK3u1B866i
KZYxc/YQWYHrhK+fijv9dyOPUH1xAOAEDHVD+X2jrKMxXlzN+PGpU8Hg36egHQJ0
YBSx0DceHacmp0KTdrAXiNUJjNIKoLWoO7in8jRU0TZUBqSdbAS3GW0cYhdr0kHG
WbKlesdeilzYM9t63Lvk1l3fogoKn6VWzkc83xYne8nXIJiQ0rqx7RgdLUbG7BcZ
6GEShf3WcdkyD4iCOEoEK6eO4HRp3hUuk+3sS9NfbiG1RkUX38ETbe9rjB3UH8GO
p8HQHtiZDANniYWnJ4LWpPPf779c+oXd6RIx0tpoaOJIyVJ6RdKyS6dU2kf/jPTr
hD8f2fnCuPRvTFX4vJ+fpr1HouowBJDHEBE8lAZqQK7041Gf+7TPpyg8WtPPYR7d
wPTco9OUsIvcu0IVN7UnvkWwEK2i1sdZG+iwd0cYFbeYRxmPCsYdAhxwAlIUVhLB
nAUo761/JCV3EMPgNrQWx1R8CsvSNeOEAhQC+AEfVXX9MPLXTCqZkvHVrx1KNtqe
WRnLQO8pw6kLrqx1+4je5qJDyutHiattPhuDpg8ZNA0aCVzsFpI6YJYRlrpY+7V3
EPuA37NdYHgSzF4CE+9fBf2Vvqzf+sibYkNZtTgfR3e9rMOvovwX/EuBZQ3kYFoL
6zPVmVa7+Oo8SKzhrXkQadVMGkrGnlrYElH+ntfE7ryrPtvxqKwE4U5+4aMo6FBM
3L7ycgBuvoABgiR/3dLFdQon1wMcM0a5trEqu2fIonWQWqlTRMssReWG9PaIddND
k+OGmHycPBN6Y7Bujq8aa/hAZtfl8cjnQPn25JEvCBkQaN7c88P9kOfiTlZkl/kr
862H8nb0+HodFuYAQRMHNvQG0W8LTE8vLNiW4pn72uxEjtYhrvuAZs5BX80TDwxF
Db63zzknS9AeHi2U2lvpZtu7qXPhvJOZv5XwfawK2JzUEEto66+KodVRabz+ZP6V
UHpnUwj40dz5GOusOgrUhYp16XNCU54J9M6FQLav3p+0zdEEN/1KhNj+Z1yFfSrT
QAwE7epb4rqyXzqVyMIjLq5NGFaTW2qaf3pTa4tQRLMiIldZdD2t1XO3AhNbZifu
Qzxzgxt6KKfnf4X33m+CFADF5qFvqF3BW0rYhuqSfp05KFOh1Md04KbrTD9unc3f
bEcntSPCav2/ktM4ET28xb+IMASS5wVIeYMhcs/bBSJxCTtXpJCKTfyyMpuPpAd+
i4yvHE5qzQPo7l54TfMkJu++5qY/62eXg3CQhoIyE4HRQmtlL4LYXEGNLMFkUi0w
IVK1Ve4ibZetmupPEVG7I9YCdoBo1i3NRmPTWHi/XbsudnW4o7heY4C66wmCc/tZ
qAoOpRttjYCbGKvf4MIkCbYUiILKRnAOP8r+E4rrx4zn23IOoP7nsUOW+l/WzScW
0AwNvvBUS5UJREz3uZ979CdU+qFvlF2a4KDOAHtdla8BMYnvtMjICoUXbCrKIurl
r8DP28J/2FjD0NMTLHF6AYOg/7Pm9LWpB4IdS3Q8yG4Ytt4FVsaQ3nYJm6qkpitj
ztj2nw8KRKXTjlgUgFecP2I5VQVqtwIgcWVmOwIR0xsfBTWwrMMT3CUFnyQgJQLl
2nd0U+Tc6cFraJNfclBBD4BObHn3GY92yNioe+SLBBbQOyaenR+Dze+4DaE5TogF
QbOTxyc+2/Gv4HjG5ZCJ1phGKdiMzjjswqtq7Y9DJ+aeD6DoimUG6FI0AGI0HcII
RVl/T5ytQcBuhWH1bkvShwIvicCyurB0dbpdtwpvPkFzm0CBeYhTayUo/wHP0mDc
3NIROvtNqh2+kFPVAeHgBOIEnUVFBFvHw3TfFFwMVb2Sh1h8OmxFmCxT5qCl6Mdp
9vhiIgop8eoVUb29246Vsn+WkTPi4LI0ne6cZUgH2BfoPjXrcXbklABG9FMekJnc
Nrxa95Rj8k/KvlNOf7mUolcYPvo6z8zk8A9Mbr3lfXoO/uH4IYLs7DERol/saKWe
Q7VXNKkCWu9tD4VBHpNS+p4btbv1icgxluJ//sHmIT6TUzSEdWWcxtnFEk6EG3aT
AqoqTC6v8r8tobGAixCGbKuz+PG7xEb49+75jKanXPqjUPoup95/AQR+3s7yuc7l
xKCLwOOsonUqlYNlKliUiNrPfRWaAE7lIVe9654T96YtVZuKDH+yJR3jocUhyzd8
zhbrPULsNAQZVTMZ6rOPIuOaWkdeIOBDEv3cAO3PyGwp+MHbMlyurvA5znqHOXVS
ZKlx8Tw/hZMpbDzJv8NGEjs9+iIJqAOOUb/1cmKtjEWbZXXToH521YAvH+q3PnJR
/ABMvPQuA9fhYJ8aTe13ocfZsQWBSqv/aHz79NUeBCv1pmxKbKahHHoTHiK0IC4l
NAj10WlZXrYN0XyVi6nlA7/l7GuVidaAgW9XOd6N+SdsVDYqZNElTDRHtUryDz90
MVenAkpbWatj+H0bMLB/wPQIll4oYrBbO/8gR5yTIHCcRvQkozcuQpnoEB7ggMN/
BrekmTG/ODYSPsAgDaYxLbHoOmXqGtM6Nd2KsrNQrKpzwUpbnHhreNHVTjl4tg89
1M2XiDXrDQlGWNk6wq28tzy4hhjT4mdgIc3LWNAHfnguW4h0rsMaNnebNy6SjiKO
dFeOQtEnUX3qMtudrm9Zxhdu9v6bX6m+tZsfBiA0Uosoopqk0WdxuEhkeeXnCMu5
Ih4zPhEdtE8pJaC4UhLbou1qqkQhb6LR5RAiPZ6kLc0pzbwEAsu5pz/XlPRm2m65
M+DcjHB3FW7p/9ni/eLklAImxZ+Lj82+HoxALb5oEPrcvep1QMsySdXKLHkWgthN
lO1Yv5NgcVg5KYBSfZ5WPaDs+EFUiwyT/N1DDIQntxZI5j8XTc69orId2GdGGNf5
Fed98MhLXbVFnShXZYGVMKMhnrbOrLrR1gv7QrhP4OnAHejKkJwzw4XCVu4+JcEO
McAqpYffULFn3tTyuEGZXEuWgPhDrulgqZZYVcVwGOyiXWyvHqiBjs3//kea5HMF
qThRTkqHnfGCR+M53jIewkWKAKFZS9wg+h7YfxtnklL+i2tDiZew/I36OWsKS1LL
EHHwvlLPiY8Y/M5orfkF1BDzGSxv3pd9UMgT13t9DtU5sXYcDMfcT21VlADzqzyp
C/oF1NNuEUS8AchVo79KW4rvcQngGP1xCeuHNLbmJoA0JvPO9YfXgd0iXY6hcsmQ
rBpDHsLrgSFo3hNNH+fJt+c6wccXNMJeSgK9HKnovujbdeJ9K6rTotoWrQglTjNT
MHr9V03bGfQgPBM/saglg1E7+tzOSWW8Z/mnUUme5cd2UQexvH4IAH7KzcnlxrPk
g4zjSMRvPFDdyJwxCZwWe7X0nj/v7814kMoY5KdW+XUuCFQaBXm6BHMYvoaK1RQl
0bp5jOH2wJXYbtFXrx73yaIfUDabCLAYeOrln4cUDrUcmE4L7z9olQz6afBAB55F
0Q5MDVlPKl1U+4Z6+6Hc9IrmdzJ1Twf6cMtNvj93aaLWEtYunpcT1SKdsT7qouw+
QmarTkt6PJ0z25K8oc2a+HlgGpuWYYLPt/Xqgm1lkRD01a56QtHTQ4mIds3MWS4t
ii2jF4SiTSz6up+vprC6Cb6KM9HsrxoZnuUJpYIz0CKXtTeCl0g/VpblSw3DZGH2
+5VjqSnczIc+EjaLbjJS8HNkbT8KfUjLK70eSMJsbN+D/YbOjnIrZGYcwENeLLBw
ly6TPMslzFbZbirsJVTZ0grP0ijN+A+nbEYns0950xf2skh7iNWKF99da4IFhuwa
W6F3O2pmZtnXhO9GeBvlnVkLQq9JTFA7KjyMxWozpDPn4ft+KpaZzuySGw3/nP4G
5NGFJefau/xAEA+1oUtiMvSSX6ItF9HrcRVAmvEptetjw1FmEEgmW/q9IKjimcWG
hbwKjmgMkNF26SveFAJlurht+Scm0SIpPx2NIXkOqskVRienOBJtHISAytglvhe/
Ji+yjwVYaq/yAYqD4W4ghCnSuqLwhZa7bKP/wp/Si0bxJ2jPIhUXLJNozRpO0cKj
g6higZDjR+TpD3BfA3lVi5WQnkdV6uw8RZj4NzkXyR8dqjrkCzPg0XN7/FQX3v3z
j5apoVu2JaKFYfWrOarnUHi1XylR0ETcDICueaqFQWOaLaHw4GzN4dk8X8piqvPW
uZ1WusMjsvTwyas9bi46Y5+sfv5wzovEaw5pmR+K2lRKBGaJjbcHQ435OxVlHjOQ
BEdUhFvtNXRB+ldZzdrcmnefUnvq3fd68pRP4JIRvbYRbdmvTJwpCH6MY7XpHVup
nZOO8tXzBM9PIFSFdaW2QXpon7k0pFHjRNuuA6jz5/YI/ne+Se9Ihurjg8LMd8OK
jrbSXJVHn5n74Dv4MbUjcQkmEloy5D8MNxpA/FuFj3IxL0Ow8ZduVpSnQUxGeCU5
Vz236E0KLQS6kotOvhCJRiVbKBg4qXzVOq7LtcZo+yspLTFtmsasmd4ztmW4YTEK
tj3AMnZwaFB0/g/6DeDltr0iOxtjNr4jMKBdOD4zz+PlzWXp+BCwoJ5G9bX5tRQf
G2XOSgYR0AckI5KwKsPeOTMTBY+rt3BZNAbqOYQBI3sJlsYkqY13hOT7MCIS+4cu
14vThFGFfjPGN27HUwR7/mzXBCSgZoKpUsXAcYhobtS11PKLh6RA1ngh1l7h3il+
f8PoLnci3Q+6NAildEt5dtvrLU4xaMv0Cr6wrUJfxxC1sHG7zTNb/DcrT+DranRn
jqOnOwmFAerUQgTnxCaG9it/CPYxOMI8o3equZAp18SNJ8vFWtBHJlV+WIIYi7ns
/IehdOKNNFJGPJESMv4RcUm+PacGmSr+IrIk/cr0C5VgNGvRALPuyDTcI23h3S40
P5HSJ4b6Ig36fURpePSOqGZuRra6ljBR8p39ooTmceKj6pq+4Y6YqY/xaufrh+aA
+DedVoXaPDpJPRFz53o5nOxMHo2k8YgreMmynlNRbGHvopSexI7PWeSf3PxfNYks
l6UGQYguixYA3Po8A6KfzWVFC+wagkOtwNla9/pxqXTS6NbY4AlWYptQvBd68dyN
0W3bc02AckOU/SGWQf9T9SMgnettRvd7YGyUtc96Yz+jTKi2NTEe6sQb7hrhd9iN
jFWCLDsTGDEUnGgjjYrwFaheZCQ6YbDD1G0+5HnTnVuG8ITmJ3aDunUgIrZXlyuT
BNPHQRaye+WMQDCWQuNrJ4tJAZ+IBTvibvqqpbxrfWaWe1xsMhu/tO8li8FRo/Iw
MI/5THXYlgN/e3lgEqoYbwq6qd0rhA7nw976+ugSfyO1fKiKCKamqy9Qj/LWDD2Z
zuh+jwXh0Or4/U224I5UWRMojX1Mbt9MDflPF8EwbfTwfGmEyEJ573ARxgKYGGO4
1f4d0P+JHhUolpZoz62hrxGKxHRDU92bm2tTHPKK5IYkbx3fgArSN2gygqKBkjp6
V6qXztCF08nsXRUUX/XMBRkUmB4ZvtZXcN8d8kDaL1Bj4Pkb5K2L5BKxPBA4dO5x
0P4HxaqA2wMlJhJ8oRuRXfWnOVdLC+M/uABbZvKEHLv9nFoguNqDMoz5fWv0NI/s
14gsqmK492e2ER+5TlfLgnbXGrLmfL6ZUNklHgGpoC/smyBlq0RPNHKDhODP/blo
EiGBuibBIAHFQxZquCivm1HYut544UDFEGwyqYeZYaC3n4BqPb6607S07gyeh98+
MiCG/oluxk1FBhS13h1Vi9eGuoJA2/FQyYcw+9KCy5hrxNQ8Rr0RVipeh4A3Ntuv
y76F453ij2bSYd9z1vwiEJYNmLnKFTaEwMi31v6GczRGs5p/BRSvkehq2/otNvck
BcxSHhjHzffl7FxJtz31xtTzunkL6NOzvbIGkgcyvMVl5CZzjXGJkroiS15e/NAk
7nB20dzm8Sd12KpxSR/4NSb9KRr1c1TJvQ33o6c/57hZtsuq/GZ092lx7Lgp1WJ2
TTZ/Q+sZXUOP9+lrMswlIQr/lFdaBV5teF4OIMsuWDUgq3xFJLWDZevtNUZ5sX1m
WUq22GPA/WEmtrYEyU2GfSnk7frjWTZ97Nt/hwB2/h0E1Bf1ekD1Hkz98QDaj/Kl
iz7dQ2hqdNwbIqfapXmLaXy2SnoRiZJhxEPoH35GK4/825sitDRv+IdTKlueRobG
MFzoj7e9LcSM2/Xc0bjyYpOFBYqRzjjbJTqalI28upgdm4Tc0+Rp/tK2+sfOG3iL
RehqQzvwdNSnVDueXpSvGt8cMve0dDZJFXM7RO51Qzs7jhpiZtzXpUuDuUJ+Tvvs
BxrvsWgqBrGvQH89qKzmLuZuBCZEOHH6DtddQFeNpZhwNsqaNJ9JGMWssv/lAW2y
H77pVntdS+ftXADzJ5suuLiDbXse+cwmCRbFo/oeNKdcQVOkAn+SINGqE+/p0ds2
ubUnBvvN5cpYD4Is0sRkDmKAPOQbXrjSSEs3c0eptqbQxR7xHxFij/HoEWX+SkmG
TJR8sVbNFDLX6PDxsbzp8jPWhEW5m6pITg12N9sZ64F36OKM8dTN+kEyqfh2APmm
7htURy/WBY/B6CttV8N1jCLsTQCnmjbpCVq/cSe+U0xlF9tQzm10iRW+YBBhp+yA
VgA4WWrrEWzW2teTrxv4Vn79REOGeZHmLNaKnU1DQ0/6SLTLR0gXKPhYf4JFmfqN
q5j9XArK4ijU3o02fWdOdB8Hr9LsawIvY4V1d3M4xzzzNILDlPsbf4lgT6gL18E+
4GpjrSCOqg7Apr9hRef7EGltAlncBu85fpIOFv9cAkCWFRMxNF47A/Z+b5abY4vN
kDuz1qeAOUEnQnHmhJvrkdMBjaiAK6PFFIbDTALoGOvqL7TAENCG8gv5n8cfR8i0
HQezY0r/EFduY78PhHD4DhYtnaTjGoxRqGGo6Czi2T6JrU6eLhpYgZ3+sG28Yxgr
MhC9pgqBJ2oWLfjuPKyw2xeNRPXMP43SqES08ugDINDpBTn4hA7oMtlOsbWICXlW
TjVKdhjTrGatW9nNQZ6gLUWAotdg0XLRab1+QMjxnhEDipBKKVFyxuuxN7RVh63v
SeK7Obi/qV85AVSWePcVe0+nuuecphOLRSD84MOa9IxAgS2+Z7jkZ0CjFQqgHzYZ
xvr4HsSHy63kdRuJ/sWZFYW3P7nchFl8KUm/t5dj6b2JOozJ44pyH9s5Qt+oq/I8
sJ6E6J6w93njY/TaOu4dFqx0hE1yFcaYyoHvhw8ApG9AUKIudl0gtxmVMnPAHHCH
pivQ5rJxRsnvmP3dJyexkVE2q9RJYLSKh8GEjQsQZcigyF6CsiNk5HeDoOw0IETs
UXbGZ2C1+V02kIQBeoi8YrTKd4/1wrhE8s9SZrBvzDtbKC6MxDXnpOpS3hwErxWy
nFmi0tROzIjeETUNaJ68aNZcAI1+2AXQnbdrROqsjeUbmdNtzhS2JqhDTymS4gG9
w3col+g4VY6mW9/DuJ1bXUPNH6br78Vos8bkigFRNZFDrBF/CXZeyXdjZTAnFuEi
rwNZqXCBC/EirL6SneeIm1B8kI0mneJG0wGFiqZ2j4P19Pc1I9Bomj6buvclZRI/
bYRteT59lxTLv5yPEB7YiJZbLcuY9wjgU56r07U/2ovapbLsXxUVFhUWTfjR812F
VrUS1xpfFoEj6PT/1C8HONDh0tHDS8K0rTSc7GVeljDCYhMriN9K64/4A3QexJUp
XLj9W9gPuTkSkV3tiOKvzss9w8GPYJsbiALk3K8W/Fs3/e1MeAcgr1/akSaLvzfA
K+V7IQ64xZrdhcas9lAIRBr1gVH6LBIadJ2L9NPYwQQ8L2DmDMvs4L4ULK8vDisz
Bj0H4v+aduUszbdpYjvsVj8eGcNFztpPvRycydPL1SAn8wcdXrxPCerEi7Kol6Oz
62yTKxbMjr0Z/zxXCdpr3n+BzD/ZYggWykR65C3BmPHnuBRe0zUbnhAoTJxa9VmZ
Ay7i5LDr3VOS4wt6m0HRDpchSBfznoQRtkK76PcMJ1KLya9+jaUkSMnPE5IiZpzR
xpI2WkbO4M/oN7mSfMTSPnxMfHWd+0E27IcRUEkfXUj3tgNq2wbyWuHs2/CInNU4
VgdRKCn83yzjxZKtJNrfc5XawfX1AJERIu0KQVdHxqSIqMNL8ARYr90RkRnGxgu5
EGynyeOoQ8AESFn09dLZimmUNK8tH83ZzLV3eocvsk7LCfGSyY3b2v9txUqpeoC5
0oUcyPmDpxVrmDgmMf/Z3M/U4UocIysQmvoE80DsX22St7Gog4OdbFJhNtCFOHYy
koYmvdL9+DO0rEUj90f4GC2Im5piAQkZcLBLXZGrkybfqu0yvupOi/KFUv3VvEzd
5QpBLWiDN6AuwJdmNx4SpIAVP6H6OQSeo8GbGumXGRCuglOdyn3cbqRqPqVqDCxJ
t5MM0GRgWNJbk92W3+Q5sUC4uwQ2tHXDfKHGSWkXw7vi2smK68mcbzei1rpx2A5G
7Yex/83Co3Qa69bttM9ESjei2DfziECU3eGdP8KjBmJM9lQG1BWD9SLJcdoXXLC9
cUEn6vRVnS645kcWtC6aDIYguwE2Y6nZLrZrgtG5+Ie9zPgprM6sM6TK/Af5IOm7
jq37iMgZrg5atxi4B4w1ubBqGU8axRoikByQD0XqrOMlew4bGsUDzVeEVCKEUg7k
n85Wnd3TaB8oYz4Xn2+Lb78jdGcll+nvvyFKykS7u/4RHT69qq9wygd6CkFEW1Kp
38C2lzgsr/CKwpZ6tFgXz6jwUSKjh06DwiLD5LzPoVjGzu59J3obXTtbidi7C6dH
lTvVfSRgJ2wrNj643fhGp6NPfHedDU6YqNn95h10SFvsbKpkvLJJ0Buiwq7shmAe
rJaeID9tM6RvvWiTIylpfnEiGcVV4PgCaqH5UVnkoDp2/dhK7Sif4zPX2LZs3V37
voTxboEADaPTiJ0+aR6mWU/V+etJ/F8epQMfhXl0WS02DLNK51jAwgZnPivzFTjC
AM9Ljc+XxQxlPlHOIFW50Vyx6NRQgANqKkUdULKLxdzU20AsB01SqPNONpn32nxM
KCf9HTGV4bGfCqUuKcIBeaYTcm4+IUVOEE/Yx07p27GlPQESqdj0GjQ7Guu5oRfS
eBUtj4HKFNTTqzQ3Syvu0cVtVIsV5tWoDG0N9zC4YLBJ+yYqd1t8MzQ77Qi3Blfd
wcEsJU4Lg36Drbtv3C8nvWr4N3c4FwcnA1zVzZ6aIoScloYyHmwkxmj/NYiiWlyp
09Pblah+NFFsEY/pTX7gWjvfDa308+becORKOsxsaBqfjGccYKN7rQQJQqVDCnNF
mvYAStms7ejZEkrDb3y6p/A9OvrNXuGnJUvQlvbSB/VBHtV7Yf/qPAZROGg/KBl1
b8naSsfxT6NYJzHVBF9hHucjNNZ+W0GHN6++V3YdtbceHwp0ukhd9G6Af7aKzv6N
YzdJExsP8sGCIxhPQ7R9kkLzsJsn+zvC/CkMK5GFPRxjXHtEeGT/nv7OvznJP6e+
Ic9loh1vt49fsBvoPFhDJ7TN/n0oFApSL+iQtg+grJBRztyJMqlGYhqrCD4qkXCb
54AqYa4WRZQF7VMxuS7lSE5NIvN9Oqy5hDPd7ZAXhGpLoV5w+usMLVSJFIUQ3zmY
/HvRrACkSU+D7FhSaeHxgGO/awmNEU0KnW9pnd9TYdlNM/gZrn1PBUGRBfRUXBAc
DDsGNJ4+LOz2x+0N9YsOSNblNzVxAxAfmpuqz2XiPcQcb0gSkPqBhaO3ahuymI0f
0tXzaZ5p9ddc+LX4OQcxdVWEkwixcUiLYOUwfIZs0uW2hJvJUlaiZ7mswLAKwL3r
buM+0GS89IoluRZl51CkeQgRHoX259miAfQhEpwcoI9FpCueiveeh1eLeFyvPULN
DUyel1TfcdtgXB4Wh72G7ALbpwbpgRlM27ra8oC9HcZMmKHtJhVfEO+33bxhxgJR
GnKKRiaIwLdsBNCE2LkRVBz2QHUPqbUdO6mFJjLK5OTRsJ4ZzB64COnD+c2ZV14R
u/Gfhlka9Yg8IJEGw5x752hPxUZPtEHmV9XJvbwQm/ShkTNm1Z1rATV/m1OvmHfj
TFtvQGTCh9mzw6Cjw8Cw/5vKCN7VojYGSLdIDa2ukiHuEogw2OlopeFUjvAOhUtZ
CRyzKggnmnQLLfpTIp/vPmWQS8NB4WeNF7SgVej4rCXZRN0RtVZW8/v1iP49rJa2
hlhVM+a8A+7iHRZkUL7bBJd7nN/1eryu7HX53m97EIXsCXRo5JAvmVNbJBArou16
w0hRKQsgAF4rfZQrvxEnVLq9AW+Fp02sW4l2Zh6NnEZDfN5XPOdvX9F/+813eVLT
7gvJsITOlyA4+n+W/wvBvYt3/jHECjNjIHtJZK/4ai9UtJlwnVR6oCu0KjI3W8B0
GNLBmty6tETXM+Tf6GLlJ7lYwTlcEYCQ0du/XGKggziFl2C459h+qSVgkPxHCaks
cWywt/LmYWexUyh5fvR9Ikry1QxnheJLzXFskyNYbzSkVTinNHNCK1RGNovNChUZ
aGw8QI7k2Nik+89hwRZ0Q8L9EdrWP9AGpMNwbQmUkJmq5WH4TO5i9HGvk42+9eFG
3IDxJHHeqbKc1TQMzhe0YeNaCO4HYLghnHriVDwK64ZDsKJq0KaKDjNZii09H1FJ
Xx2pjEwPxkgq3yiYLf/sTje/RFFPF0iAfRe5Jn0m0t2r7Po6zTgV8TXZO/y8ifSB
Yusq9+DrP429uzD7mt3ARvBU3ly3NDbVUmar05MMEGXD6pVXzpDuQUVNTRsw0Wej
J02r0Mk8a5MBYcDcXwX87f7QBARhDc1WCT6WmGqvo7e9MlGXZ6OI6rgocXRVE8Ju
YKVOlt4z0oeW+pHWJQyyWsEPF+v8qWB/Mm5XfdhlizDT0ivD3bw4hv213B9ffm5A
jwGcm0rMMupAY9WCYvyPejlC/6NWbjzQjZZwGalNVqiVCPAuHZF33NHqW0e31/nJ
ufEIxFHUqrkh+7Efjul/7fbY0a1/bc/T04gv8qczHTWYX6/uY6qGTQfZn50Y3Mlk
2C54JOia1tas15HJkHBFVdV7H/1oUy8y7Byn82/sY/LaETImmRglw28Kw4crRnMY
PLk2TDSn4BPEYZUjFwz4P7W11HRnLbS1o3L7g8oFGBvc8U+BNwJKbJvxt4cQobf3
vK9zayDPAF0fbH+CN8j5w5LfIE6Nr3h2OT192cJoDFfgFZ24rJi8ajfkIcMkHnBy
A8/4BvXSq6BzMAuM16dBfvDvZI4arA60rkpR1hOMo9ctfYik1tLz4gkFG9JpDKio
KwPrx5HLK9QOHNGgfq++xr2HTVOhQDgjBhTZFlVXMCJ8lgq2QcCXLPZt9OAdp0oE
WpHy59Ye7lMqmaFiIo7n3BLYDXUYv9tNtNh4hyxDrK9JVbE+1OY9v0tIe2HqyCYO
6bPj5nZIaHcACZyDQZtOSeloZnrScfGK2nUm/NkrkqTV//0IyLViRiCc2AYh23Zm
4mfEJAtToPfStEM5HofRUHlVrGO2rFtEAcOiVfAOXNWVAmAHKKrvEH1biz97K4R4
+0vP2sSbuWxIGmwOi2yMNN4eN3dx3mi49IeF5O310+8ejatW2HDDgysSvo5/TM+0
eQdo5vmF4AhWceJKLbMJoKTm3cJ2bpf2f1dhMk6w7OA7nA2bz73DD2gj4eI3NUXK
lWnmAi3GdJ+9fGofO0r/wLweritJJkr5QQMvvW13+LwzXv8/3XQ+MeFv0Vxha101
h8zEG+X9o+4Tm2YEph6gk5GR9FIE7o41HlVeVrGwaRRuvLvrMhMjZvjK79MENKWc
vFzoiNVEQ5QNR++0priJlrUuouICUUP2gnSdKN8eu2HrFBucmxGKP4fN070nJK/g
gnSHlrT+INYQqp387Fj2Cu580TaLw6QOIzDCCF3SynihV3h2HcVd0OGzDV0zsZtz
wyKnVzZ57Tx7csZ5quQjGEVt6RVypBZHsHwF56HBshKbRdivDhJNyEyjbvlw2DyU
gxUsc7eJtAcSrA/ryEK/HgBnhjWkKOnkunZpNScSU/hU6VrRTNcC2e+nulZqNngq
TNlpkAyr84Gr75lek7N3q+4bHrk9vSkhR6wBfKzK38bmkyxAnA0/jRza+vmNrVa5
eGPAiyTQzNcTLBYguopl6kfKKZcIrMS3fKu2/qVB8i9zajsslYTUZ5mTcvaJCw67
+yRD+iZUQxtXD9+BDm8CKwVRnF8fXBRJsbQ80iYt6B6FevSWoV1HRgdGfIFYH9yW
MFxEgE66r4xwG0x5TSqNOOgkyWIDG6IyEPATw9aTdap9GkLfH2hh5AaF+dBPfiZR
Gk8MXxOaIl0fUaFUQDNcoZ0xLjY3awVishfOLpSt1XDHHbFRUSb3qzHcJE6ByqUR
XCqfkrqebtWpJz05n+pTvj2MUDQeoxfCwh86FMeR+sC80ouSqr44ly63Wdq772gq
zSOcme+oEiGhh6B1vsErHfG0hinMzSVHA/j49Wyqd+bfJ2DjbS/ZHoYBTkSnGnIQ
ZXCXGWg4uZB43IZipBLtQex4FA5qZg6E8jiis2cQJBpmiNesNwEQfgcGowIu1wev
DjaV8jfEZc9IyxveJ/2CEX7YNAA5wLXAcbGJ39i+d0dTdfcA8nPl6CF7Wmsxz/Jl
C2I7NfTUbDJMK/WcpPSU69bPBw6S6yEO3JT3dA2yqmNLvt4tZ5JwvnsZbAG+6JFE
hA3imT7yIF0YSIX5RPF+oxwbYoYq1JE0rmvQE+jl2MG2F77gQtS1TePA7FDmZk0J
cDLFSRz9LHEVU6QJsgIseyEOZotoRDyVp2pFj74EJvgyYo70mIvGscMMGNV/Or+Z
I9RQJkvy/zmrnoKHBXdZwLeWFrHzQvOSNfcLoObeW2GSnwcnm71kxSVM/5RPto+8
epHVoXP/pvpzlcEsA18HrxNNWBI+4PmX11lpi/9SDgWc2azqh5bYe/jrHDpuqu/Z
NKSGosQYXJHIJrRo++mw5OwOTBsQPh+nwRLBdQrFMGc+0NAezQUCtG0iiR93f8mc
TftGQVqvTBsASV7Evz3A7c8uWtiUbTJizR8VS5PNApC8LFprksFUyVnUMuIH+HUC
QNSVIzk15i4QzW2MhYO3giruvPNyhVBwKqSaY4Ow28uXgYZNQzBR3SCKDQ1q995f
Fli+3dKIAlzhVEARtWnR9Y2WNWLTY5VOAPGtPQMRCIIt1zx3O4xGc37qofpgbhfO
8tYyZ/NkvwJbJkdS2AY7CHcJxOoM9csLuVTuGwbMrSmEhT6x/E1vXfFnP4W0BHs0
ZKw0/KzcOcj7byeNKn0FhKhqeM9322QS4TFjdt0X3OHhRhb73gBw6JnNX5DIUUyY
CKlaVAp3ZbqWB8jLVVBH9DoqSzSTQEupVDMO0oAoYPdxeRn9OLO3w05fVdXodcv6
HtTopPQIBIfwAysE6tSJKBXU3jBiYE9tDY/yVv6P2vXYooofQP+uZlQ5efU3Mv0q
Y1SRLKv4zgXqUGdtTHVHg+RrvWMizq1hdU8smcdz2re6QcYQNocvHFAHgwXGyQxk
w2qHQ5InrdRSWjzlTx/ZEO9ty0WM7cE31uMOKCqY4GhwZPlk+k31sDKQPuK/dPJM
I6MlMtzQD5/4wwgeYLXWyO2a2sx0wsnQxwKmqJmYmksb6oWGlI6LW+dAW8MSnkz6
dmeX3iKrKGpUKOhxCyf0DGc1cUGoh9RQKuKAdDJ77/0HnlUEmIxt/X8TidlbW0YP
T3+r5ddhiQcPCfZFtqlmbwqAZo07d6BjYfszaorcj2JmZaTG1UGq17iI3ohSBn8K
546niXkH6I9gWP6LWIEC1aLu7RaNy76u2qxDbK6hSLUSgzLOulHBza3Jy15eRi61
U6DYq6yaVumD+4pYDPq5XGVvpaE/NmIThaQAl+5mOj7F/WQrrn0pLhieI2uoo4Cp
ucUryrIS1dkuCoRQxeMX6mYlI54UQFwxXvByp0k0NW7UHnnJ9x3wkZ8GEglNnjQv
TeAI53Ydd7Ryi3rZE/3k6nB+7GTHCz4+U/o5NjOJ8hjIYZ6dZdzcaaWL8DB7nVtE
zDSZ4Caqc4f5tosGv9jMfjAu8LQ3/OWPOBVexiJcYD0Hj057Ia6bdRKMWTkN7AN+
EX3lXa89TxSCHtOfxImq2gNAIQi2ZgUO1AVsv0NBLvTiHkmaemEadOl1G1ciN3y6
+Bdp+gSRHxjHTQ1d8V/ROv362tybVT8fTae/Y2E6229Wvq6cRPbA84dszduefwsC
ZjySHGN0sY+mN/lZkMCHy5Pcx6PNo/oJvUNHQpbceqW0wwAh9SaBGr1RLZURzCns
lZl17BWAq+Bdq1B0ytJXTjHS3WW2w9xncTjl9U37e/BLLijhRu4Z51jezzdI1EqL
fl+1BlnPY3sqAy3SOhB2lf6gEYiEciJypZu6PhCOg6pKA0UbZFUZitwKSseDe8Hs
McJay5wx4tWfU0WciMc2RzptV+W33k7gqRuQjTaPp7Pm+IzHPPPZ34Jt3m9S9wr0
REHrZ0eKLFijOzAti2tapcLcZ8NJB+yZYJgIpzvPU41bk47ynRC6PLqLIE178mBv
Ve/U0DMuZRnfRl40wW16ux/m4hkdlt7bjxlwhbIOjQJBRoThUZRsBucz7ZChFgjP
1Tq186cydzpolSJvygYZl+TIdKRvmCwny/nugp9suMOPgtCAYUzK0qN/XJFK7PbU
1AndE/xERewCNo2jUJ/AHixdMALLF2tfqMpKtZI5aNkRzJsQLqW2AoyPzPE1zAAF
BQauECUz8nzHBuuvQyHlU08irsZE2YuVASjKrzbEo9Phyuv1paMX0C9Ng989tPyQ
/Bbdc5QW+N1sO8XxsXIJWT+GzX+ucZ7lCHBwsyJwVUFHVpJzjLa1RugU1MDsarBe
OEh1tI2dtipdo35K9QszLq/iJDbn8jsAuLrRM9usnnqtGnUCzH/PE20CcD5ItwHX
kauwEd7O55Quqf+DM335OEsOJ53ZXjIxSGR9GvlAqGH1V7wkcFmiit7ADudm19WP
yiOOgEFBTQPPAmboDMwW6448s6vDQ/2OPGC+9+CUkiUlmAF16I0om7OcID/EEE0K
HSM2b5/Sz4HbuzQkpxrC/Tkek9alCokZtPbZi+/oNuRLgrHTt/YdP/WM46Nbgj9i
09c4U4VIBVAZ1nC9CH1F/GDxu3k863cmCT3A5IFEM7HSmY0LCRjliNXS/KZwk3WC
iNT/jW9UW+J0JNKuZqT1bXiyzSKforzcmmYuGAx8ETeFaNTrhoPaIdwBtexzxhCv
BWGvcX96dtjVzgIYQa+Wymu1nCM4/dO24mVHWOdKvFMUMm5zX2vUPy7yUCi5KFxr
OX1/IzOdQxCzJgkdcC/QINa0klmp4kga3Qsx81WJX3ZIjav6UKfjJQ1wlFl2XvCh
9WTOkGIUGdYjQRTdVLpHC7qwJAR0AGjBv/qlkaXfpr6HOiQge574MdmfZ3bv0Vv+
3lf8Me1DpQpMVOr0wr5Vs+j307OSEhjlqskTWnkGdZCnFeMKhtOFwscdnIPMYNaD
gjA/sHkHytdVc5nLx0ieVLVTZY7zL/LCRHZLAwWjp9D3oqJ4A1hflDoZkjzV3/yP
yAEhHn0zU5OvqhF36RpENMJBKysbHdbxnutr9qr47E2es6/rvBuYx2l2+ZRtYnNn
CcXHX5ARTz9GWSCdN4q7xB+7pImHOI7tiX4fPWi+7neDsXSxUn0ye6tFvv4/JA6X
UCcKgc3LAW0zwMWQX7Cfg/flsRB51iGiW1DiCF7lsvx4HkmK0KsHDSP3Tlb9r0Bf
xp5V84hAa/u8yjaXSLKWgSZ1n+jzoWI+2wkmGaqkfp+jG14ex6XOmJeaeSHtHGKJ
kpzLPWiUg88LA38GJnWkJOvtmq6gHcQlWzd9vVlWr1+22SqBZaeF/9b0tRyhTs6k
kgp7TOAwaIWe6Ap6QpMhzG87RS9EjvwVwTEAkqaMvgERRJlBQJxA+OY/wYoz68X5
O0LKZdhqVPcubxD/0EUY3Wi1yMmRoEfQ5q5xDmqAVlgQ5yS2Le9NDlAVBqfJaAJ1
986nXd4PXP8pADiRfc+6P9zkQSbFRkKcdRmR+ox1vy4TfuHtfE62xghLAnWv556f
8GRO7y7mRNzU6M4EDrv5D7OnvbXgfUmU60/LEOlVZh91a3cFAr8e7NARBHDKEYI7
L0Y6+A20Er1pGE6EfkwbXPInXCADzWkfvOF+Blovvjoh0/cjtaGvWd/3vrKgXXD9
uYqQFCaSmWOVBnWpJEEzFagWf9B0DW2ZAw9zKCzIXqwz2DsjmOAZsVmPry79L4HF
+NQu/n0W4PpIFv/HLM3povztNhQ20vG25NjscEjLPY4q8OhDmPR8QauydC6JtDa0
21uMjgaH0ZVO+IdiNrSEePt7sXJz4tB9l17/BpGIJJbQLy0vBbTc1yx5eFiCdR5Y
FOi2YPzNjkl5R4SF83dWS5qsyN338kT+TFy2OU1MyddGvvWmdZIYWXwOATj9Uae9
AKOmruXzYfqt5nsPh3x6lt/orORxWERKLE/AONg0Ei7RU0owvOaHag5OBt7On99n
Z1pQDAQDV/bnCUemSblq5JqSlU6PTx6UITDVCgWw07xNcHr7ybwlT2SAOGxSilM9
1jf0RcoYiYWIZ/Wm7IUt2VJcI0tNagP4/FACT91QTo2TT3i4jILpD36OAyEhJgIW
FZSN39VY5hYTk7Ey/GIGRFcuTDef8VsIeAoc7QU3R4piJkfWqxiElQ2i7RSdW1kS
IaImKlOXPewWdh7cJ3xwXN9wZhO7OK95E5Hs0sajrxtQWyulfV8XUT057hDh8tjV
1cOUxisDJI4pLU5l3Doljp9pQVM0bZtVXKiyPEV0RI2x3Uac816tvPy4kDNmf5uX
qr9ktzf2634jodqTnyEFnrVRC85YjFBENqJI9qsO/UsLKgvkfF8kn4FFPLyqpA+S
X90h1/lid9vajHU4UjzkmzkWQdSB1JjahB95viz8ep/ERtDjYp9kEWDtMIWxGxME
benS2vhu1iYmjBhWFOgI8p1XKei/tEwvhFNsXGjJqzKbHZG9XQke6h16hk18ZCtT
VV1ZFOE0pq3HNWx7yq4jkglFooeliH5lr76Vl9Hhhm5Y9FTaAie5VQ3d7N5G4u2b
Ognjyu23o+A10FoCD/QoxDqa5tbpGoYl6gxJBGtyC88KNrP+8UGX56q6kib1QUI8
46aEmgiraI+XdFbI21aZKWo8dD6l3JPvRiPz0stf2aP7ZgBAtaNZAqn/ThiXpI5p
1Zs5r7ExasCpDuSLdtZpQ9u+cjUus4mFWt2sjsVrf3xFeZb7fYwIh9bG2psSNBIn
zA4vu500g073QXnv/z/+1vr2QHbnr2krlh3uduJyXmWeohEIZTR3sp/HNMGI4v9v
uCgVYYQu4kA+um5TJL6/4B3lIoxIIzaVdae60ytLTOPy8PupG6nCGcWyo60fV4B4
gMGQsEToLXATTNPgOVlIsoskphCcqiaXcuhMpf5dWzVpqnzb8Y2N0AywPwi39RU9
k/3VG0pKbAgAonV+ZNJt1FSl+n3j5+5DIWhB8XWED2VZn0h+GIfhW37zPldAhdrZ
9XMLOgvLX4at0dWut3R6ypZgVWPuPqQh9neEH4R6Ms7caM5VS+hqqwQoIIwEpO/P
eWS+NIApZcX3ydKFuTUdfru5Hs36KzMJ4iVFLIpDWfeKtomdwwgVy4v9fLCtdBT1
8QvUhFnhAD2/mWAQP5OOXrQVBCBtcp7yaugHasxfOGLebsBVMOFKaHek2T6k/U7x
lZssLAOJFiUabE7SVBmLtmCeWrakmeV2tsUXv7FIRM0AtziMt7DEXzJ8BnJhRaVg
S5V24TQGkXf5bJ9YKKWt2jH0GwFPWIbPNiCq7kGxMsauOppyNMZT/A1xcSSDO32U
EtQ5Mb5X8BKD/wlVCxF9NE0aIwPA+5NK913ZNl5LG99DPRNDp3QWUjtB/etfUZNO
odKtvmatSJcncZJrVDaTYClykIcSudCUIc6cew2tL2PjmDc72YFCpLMbw2Ly4FhJ
encL0r6LJOQWYcwgJ/JdhDXgB3ye+3KV0Zpti//1Vfo/k8T7bjRAxjrWttiT0DvE
tdFScAjHgsFsJeeWhRzDFBGO4Fgds68iPTgKIO37c4kPaiUXhRz4lEi8pJmnF6Cx
x/LaPxzqfKXzFlGdPMtDaguRvErFMfbx1y7i9juLCk+5+llDMw6zK7WalVs6fVof
44s5Xz9ZKvPB9qU3aqfvSfU5S8kcSQbJbuym03g3VDVgTJxcUeXwnyQN4yLIWzUy
sudA7giMhKa2PsRRlZ8mYLMLJXOPwnHhO5SmabhdOEdjSdQcbu5UxcBfRhATW4IE
L72asv88gdhde7sx/0CdHaDABywg/FwwXooGqH3c62MM7611z5KtDk1/ClPqwk0o
5ZKKMw004LlPfjvUU5sjR3TUgSpaBMUz2hDBTBBMFjV6b434bCZAa1wCQzHMZz3B
NSS3UxYG1qv9NECGLjyIihLAArvOZ6i/8elBZTG+/Mkjvvni6il0XEKBj/4nyv4U
kosNq3lRAfDjRoPDeGZQv2HjpllRAyQ0v2KwuA4OG9wfnQnPRS17e3athlgpkjYV
/MY+B0YuPBHSS1FLBDz2UaBHo1YEzVGn114Iwih5lCUhu6P/XzM/o6jiM27sO3HV
BlM5wuBBYeqGmFAZqbswS/HT5PJEe0MLL3G0kuA8sRYfj/hltjfYIAV1nS0hz7dv
itaKoLjU8L67shkfPXZymQXIHF+dAhvsMaIeHol/pyXvcAhzo33C7SdDztLwFFsT
AhdkDKmqXp0udM9vYwnTR+wDRqAkiZEIMmjzL6azivOeU7XZoU6mpjrulluuu0aA
lUfFFgHBByS97z3JQdr6JrFzABM95WLfbDmKhGz6Vc15amos3+ao3jawf4ywvYLO
GQajCvM74qtRICeISf/POLfGMM2hI8C7AtRU1CCSTT2NMRdPnPZz2LsVVVFBD/VR
qGFYlbK4FpRGQDN86U3W19yiIAqZuEt9/8t9iu/XXkufm9qphMiMn8sLOGtp/w5X
ZiJk7uLIbPbVaFOaV8U+u2Q5Jx+OPBSiCP6/gFkFMujsMHXYyr4vMV+FrgyL+bga
7FwzFaeS4yTG+fDlZsIKqvSBaA2/q+7AIUSlM5E3JQCdvJGiYLfvkT60ujqNYF8S
UDSrPs7XoOURt15Ql9KnH6zQy1Il/dYaFILQQltzCV1n2NdZw8ndAdwx9681NEOg
uVjLSSyECgMxymVL8XpcBYQ1S8ExcU3246CcqWqolbOvR4KcIcXDRgZavXd2q1Wj
BVa3NT+0r/RvWVwPgO7Nj7f3a2dd8QEp+0wtrbaXkeKC8nZAvOh0GyqgTWjfHZXI
lGjp+a3f0g2HbYqbdvcZkO5l6R9VWuI780uOaIl4WGPAkEfilqbnVkXYaf6cEOII
042ckv7EQr2lsIMFg5ZeW/9XUKZX6VigWelzBnUA9LOyNYmZGFadmIyve08AWH7S
pMyCCfqlw+PPbnx09+dwdd7FruEdoiWCTdA1py5tKONUoGEPxnFWbPUbM1khmDnc
+u5iGu8Ze17J1POllvXyuoV/27IAcfi2p+X0wAIFcaTkQTHrvsDFP9uQQ2AbPdnX
wg3TxT2sT7vExmw7y5LDrrwegoV/NmQEhhdIUwT3adyiUiiPCIop1fU+hTvjMkty
WhirddIp604V3/LjpA6+Q7QIjBAYqdlfp5fuSBtTTlNW83ga3eWKeFdUXj+ggOgU
oykAW1BxOczCOxZLtYxrur0U9RcZcDfiyNz7i47ROV0klBzHCcngDHjB1N0t6kx0
kTkfZdJm5WN25TPzNYR6h45y5aS/5xn0guUR1drex9ODo2LptN/NGzmHvVs1GiIg
mnY69pOuHdF+ruAtHzf81iZAGD0JLqoJ5oBbvng0EI9Q6M49+c9anGJuEcysuKs3
qlOio4Mdc3V8AuWS52iR9pFq+n4HR+sik9HgdJAzSHVZ3KW2Jnwh6NfmhIKu3A7b
PeBZ+qMuC2PNlhkuu54YuCB0IWloMSiO5afHXmg2MhhnSpx7HG0kG9jJCikZWE6u
wOM2CzC/7gUk0z2XGITR0dTaYfdtCg/shzjt7R0SUD0kcueLI+wihgdBnUbnjo+l
kvR0jMHg9tGoOfTCYUgOlVh3Aq2Ht0p657a2tVyqQkTOAvim61u2Ncz6KcuMk2Sd
hMmA4pDbsMH1E0yTsZtfmf+ll32r+834oQ6PPuCboYaGApspIRBH8hhKKcILpNV/
DpmdfbklUBkLPkdNw0H0+QcESBkqphxadT7fymhBdlUgqmIdtwRs9TDlBAmhi071
rkjG8OHWTxi7rrfk8eh0EEgBeHJjxC0eulG52h/MbQjhZ1Ph2VkrPiUJaxAkzMh8
GNQoLqsfWJu21dn4609UfTV4RSHoqJS9q89aAbjzkTJ3NWjZW+YtN6S1GROrImFb
DeFw36g6bilVWzf2KFxnhDAG+uiH5lvGjZYu9H7uZ6y+kiY1vIkYVGMwrJmgcepI
0KO8mbAvL1qO3JaGLjwnpySl2JvDehYqqOmZx+RjKFivXNgN/SJdxR2FO5VdfRrl
BUYUZfrtC5ygyBrR2fJ24KwhrKGgDAsWj5V3V+RI9DbpcP1MxzOXWD8thRGWRCHT
uF6Uz4pVA/Rb11f14vS43BetX2EB40FRhTyZszj56KCP/jOWWRCU2Qz2UCb806hw
xscZZfXYTIveRomCL16ZCkbywaMRcU2JahJWcROiDMIpJfLgYwv50znv4nHnEejS
WBAv69AeGT4S1D0yHwrfNAioD15EWMeX8ATXq11DDrRZbY8Y++khP/De4RTn7mAZ
wCxumTm4NeGmTlMokUitE0gE4S9+ubuAHGric0RCvFxYIRUzzk0TC9Ps9oQseUTb
jarNOhw8+KAxh9amQvQgjtD2fIWsfpqymsk+gkNgtwUtQygDS+gy6rMGzQGbwzsI
h87+OxuzARJe+H5OqW/HLvusIJY2Q9HZZfdBeyoOaFl+DKPTHUskrDXSfVptf+PM
/rO2zyQwkYbVjjwMj56+imkRGI7Ufrhz6ApdEQguQAgshBK1vetyuZVed6aI9v32
lknGXjp1+BFqDkd7uQOJl44FRiF0j7h+WnpUeAHAON3xXnkmIFOK/PE/Zv0LFBVs
s7+CVBBgOXCWMhvqY7bQF3rp33e6YBx1Rh350pTgHXoo2u8Gb20COHWWso+TS4b+
/CUbBULwaOrUafbMOHFOfwPRsKSFLwNcY5/dxdNTVkldyYWup/5cxg/VFpIdO4tN
WE7io3zOmNi64RqohOGVh0XndigPZibfSG58+anw/ellJCPxoV6HJSTsKDx23b/O
Ml9pXml72Vh5e4Sw4YmryUKeBp6g49zPfHVacphKe+Yum0L6n39htNXzIHock4IJ
h4y+3Z0UrvEzzVairAJlZXP8X/m57Y7zS9QnOUTw5ctpPR7DWqW5LzPBlgJ85ECA
S457X5Gl8v/hn0hmzNUpmmP7CMDMBzJqJEg0fW8HAr+qCw+WeX2C418Kt3RKzFLG
SonRgmiagqRuEHa/N02cK2OjJNB75pgn/1zJwoBXgrr8b5vuk8Kz9S9ES4hy2KFI
568Wn7mFa0WfNxmImGhqypVHmY28L+UugGn2FjIpVNo+QgA5TkYKUud4qWRRGUk1
OULvbcl7sEK+ae58gPTE5zCoAeRaONZpup3kGWcnYAvRnV+JhJU1youpgc8B328+
x77q20yMa0+GPuOA7yMIftRZf4yc+atSU1icDZ0kAVpJLIIsgiRomftPvk1REein
K45uU2z00+T4bGmfP/KNz7i1V5LooT/KKa2ZY/E/enPBBYU6gpiKZAiCTM+5AwHT
drDMZZfr7VzwmfbTiUU/bAuwyJUdAJTcMuJov7SuYvbfHvRYx+g2x7oKpmxVTwLj
oQ6KIjEbxOi1aFhPzmlyCHqYpfRRPmh2guwY5b+QwHxmsNkMUlxy4Q5nVGIgvhSL
rTuqkFock/inLB6IisKNTnLt9HnSnY8z05xB1I9RmmXHvmFdoa3gM4P/Hti8u41y
IxHDWPtvdNSMHIvTf3n3y4QY0m2O7YhlWTLRuZEwEs8Nu0nejgqqLSOKu9PB3tC1
YLc/0S2b2/LwJH96+e0Z4YNoDIOcEzAp3OvXWrZtKcCWH4Kdi2BrOtvyVruX+c29
ERMBEOUS8phDOKgxljyEzyNKgmAtNZGNNKRMjRTQM/UTy82RgW1phpAZZ7cVMPDI
qdOChL7Zn8+zTbbnaccKTsZ63Ts352lR17kGXUfVRInGRGse8wwskjiQBBiLZ57/
Htsj/HJgXjQROdziQ7E1oumMmUWnPZPymc95ynbhxJk82bvSXY45VFTdzT43uV6x
48KXAPaMUS/A8u/UsRzsGrFczCkwQmaoOjMpK92H7kHn7OOuHkrXkgon5a0Iwkzy
VB2lJnmFsLBRIAwWpEivsGeBOpJ9hCX1OQrrXnOnXo5yN542S1qE6hb8o0PXg/RY
/P2+1CeoYJj8rFg5TCyq92UMgO2t+30pFco4LImyoAi0wP2O/UjDMBjdMyAm97vq
ghYOEq7EUhijYKepphq7FzXF3R4++a4umT0i3yoLAEOy0skv1MzXaIcy2UssgVQV
XS0oYWlHUJ0zLBG0qw8YmFYPHtfSsS52UjYiKKCY4brSYMZlU0rWEUrLPZEAf4TZ
N9mTcttuigYMjqE8tweYdvS1xzvMM2ng39fFgHbeqzbu6/wDdHWwH+Bt7T1cp9ZP
G0jwdH5XnN8MAJMWLrFXDV/RNERR4vH9lI5pByPXGQ9fJ9JKvj3War4HDxrATNRD
ViMMVM6FNKMR9cl7xapeaALSJvEDOqF5fuO9Uyz7N9sxjtbPFA0Ch4T3futjp1xf
ENCxc6Lya2ZiDRhYbm4A7mWbf4uwQlXpWj+KAfdPCpiscZ2s4Tj/6AlZesY+XrPK
mkTQMgCq60FBzB6n5i9fztQmK/EFO6U6cGJx738CYo5lG2lhm0XrtEQBjOf4qtN3
XMS4b34ROZ5xKnNeqJp08I+uBaojKG1glaj2F2R/v0bU4UKLmtLZbRBm3ZL5C48n
T042GZFspS1QHnuINj2msspXydPT4tNesdJnAWA+XS5TXOuxGeVmBMNIoDuP8gi+
Xgwq95gsRqOsl64eCIK/cbCTU5brAzpD2DoVOC4eBAo6f/28f7ma04VHQaJXYxQ8
QqKWH4UsMzZ/wjFhcJUbwZnWqjgieDJeBe1R5eexUVBhKOB8Lp9nOLiQS2nUWPRT
kFb8sO3FIaK2mbLcs636cBBVN8A5t59vCw0ID/S7UcvgL2fGNmlVFjDEnTMTYzIg
d0XLqv1aiS4A2gYjzZLR74QiUUUxhcoi/GOLwRnqZDkwwTAe3ORjB3T4KaL+RBSX
EFPolVjEy3zhAdHWWnY+n1m88u5Tt4PyOQ4zJAUVjsHWWimaaUwCcfsd016ja3+N
TUeUogBD//7lK/sUMWHnDbMiZFeFXVp0TTkSyL9ZsAvwynu2/y6ETgwcqc/zl5Lh
nzBg5PAUPvHhw031RLE/F/doq19xKZTEEtYLKiR7g3+Vwnk9cJsMRdl492+ENkix
NYVoKJNKXF/EWTZhrvi/aGqltb0WB6aksq+7u9BDcx7F1dkRwomFS0MIpkzattBI
R9TsnDgXoerwn/0ETU/NmYddFOAV5HRwuvAPrEd/SRNEnKQqviVFsJgqDuGPXKjc
iOBqRCClIf8WRACLLunNZE6GCaPzyh8n3atFgEkGeFZo02YIN5emuWdSgsAeVFAO
va1riYtHZNpn/ThEbPvrD3bUkBtbw5gtlL3uNgwZWOhksiwz8L3PoernD/qqdeyO
07JNfEXshHcezNgQOnM/TjoaynICERyMhz0SX1q7RzLfD2dhdjbvNsLK57yfetmo
0aPSd5F7wPeplcPj8dIBOFSwNmQleRs3Hb1rt85GffBnu+Jg/HR5r/ZsUMNntAth
vOr6XQxOHbVK+ZQpB1jCbPXJG3S/9G/6lnkgG7KStRIvIfHd4z2JjWetaEaGp27+
SPNVgqEeDhOwECURSBnMfO2m4A41ieNch9WKGM6ME9gEQBxdxVBczlU5MrHtuQEz
mUPjXlEUsy4d4Vlnt2c5yCmuAXOSv2Q/QT34DW8rM57Zd63RODTJKB4kXQ0wD9Ue
DZlUaDuw/gqC+53asRZG5aTo3v01VMKE2Nwy87i8EMIdESiOlfc6B4liphydiSSe
7gX8YkOtvtRqx4NaKSz78BR5JuIhSay3cOuJSEo01RS4nSu4oNdDTEymLL0xbpqL
WEPTf9Ap9o6AoIXrfu8rCZwj1sG8Yzu6e42J5JpijSFaW+0zwRYVH4qs/P0mN8CD
AFFFwL8m5AS8Nna/MKB1qWSzq4AQtiLuHzOV+P0HVps2nCXGnDNzqAZ9WKFB6+kx
ja28qutw/svLVjkFbTA4dMQvo2dk6ZqEuP6WFaWB+JpDwygzzPHCkAc0PZkT3w8I
CWKzCf3vR584P7IAsbFsaHXO+XV4rh0BlhNsSqB1u+LcSQo9y6FDmgwSt9RqcDTx
Ed4ipsiMXSQUzB2oVk6RmuwKHz3ihN3TikhC63begMp6nqJ5Xv6IUVsddQPy2Pwz
5IKYuY+QkKGAW2GDoZBynbYA72I6ZKwr4iZcdYqhVM2aq0H6GDH6CTLONJGgF8eG
/o1//SbFapiZ6ufw6sgMYYUhqYDgKc0bwgH1PY1hmmw7jF4O1W0yViABEFbKvdfq
hY/jPn5ILEWxePRqTnjPJ5MqsSi1mpfkD/EY0+vzjDbpYUIFNwI+FC2b8nsA5Epz
FpcIDLtxQJwQVe/Oj5VHSK63DDTZot+XHBqIEijeQD6LGdyCef4Jv4fbRQNy7DLQ
EFy526LNjI5fpz6VqW2bPjKda6krRtTKPkQ+P6EPk7W4tlB4N6S/EHCNcMeDBGKR
PUDc/Uoif8rANeyHLYtA4vw5OvT5/i81GLS2PY90XosVFl3vJ59x/x26CqsJ+NY9
RSXFUVedtptyzCTeI7CHo+TLMPt29+4mTQKdjMsPOhWmk5c5GOHgJpVadWz2gvT6
O3wsMSwSih+WsXG+APWMEeqf9wMHn/bOWJ04yecYzF08oqPD9+JQhwTQvC+AyWTU
Vj/1Bd0HTISqsZQJiMaicRTV2Ghb9OGNpaXGNvFVW4HeIznTk2Uzmf8Bq8TC9kwg
meud07K0b/1MhXuhOdmYNDR1gG1rGsUSHcGiyCuQ7ZV/R8kXudjgv0oaRasIY5jn
1zrEBRDcjoA8Uf5fFiEwfcjXzXPHrUyd4BXw1fXey07oy7YHvBqHzkG79jsIr9Z9
QaL68XrK9IwVDUxPV/8Q7YjHtt9Q+lUJNyFqtV64fY6Fq5LexZFtbAVYxgdaV2J0
A9IN06jsoN5KzUI4olw33pwXhkNMrH39leOgIZoS9zvFrWlsD/7rkTZx2ozRKRAt
Ow5iZYOEL5IgSQURKR/GKYxl3Ghaq/S9ySD7JVCwd0EFbx50ot8iy3Pq7HQWytGa
n8MDskC0Yubg1ndA1qnpLoxD12B7oWs8bLA6UWcLDyUU9P9mYQHMwH1BlkhChC+3
yJhV6bl42Lc9Y7y7UmO7GaiUaVw8UoXSSkvHAaB/c7NO9P3T2PZcvG1cltidIDR+
OBVu2geAY2hbtrE8nDoEoDH0HB0tNTBE31W8qU3Adt/CvshmG+3aABE1YydoZlc6
IZ5radGHITQntZrArgvw6Qhngrs8N6N8O2c6D+gudVdreok+1/IlToasXYZZ7XAq
Fbv+GWjWSM2wgA+ZZROB37riIXgz9j8G6fYdDzEDOJdUOvzNP5r1QXZDuyi23kmW
QnZXI6tpE0gEwm0Ufiva37DFkBq1Nxwki8yG9G49+jC/sO656j5I/s1y5cReJX/K
ZkFhg7myEXE7GLuLTCoNg7XPWz4zhV4PRlTL2atMKU5fGOnuEuchQZ8vdQODwwfU
7GVhCdWs5jmuLQva0yZH9YHqjZBFIE1JKqbFvCAf175FHSAXzrAuP36E/asN55il
FyGMFtJnNtVI4uxjS1ib8fifS7wcrcU75PaiJ+RC7LeHXyVEsq9LJUEkP6QxNq0o
h9+rOaHK7Z3E1+q6BQPLuZGyUYUq41uIEwrR4e5e0Rm0Xv/aoJ+BhFg0UaP/8+cf
mLKi3I4oW0V1/mHIDksbgC4/jhMKUJgMssxHMf0uyJqSpVq2Je5TKC9FVarexPdB
KM0DF/nVQ7sqPZfFcNmegsMTVuWOdo1b5l9VLr3e2lzBMMzz5rLAT1RCUZHzkDbt
IaHRvRVzCOLE79dLGCsVm/TIVAkZ6GPfXAQyDgsJM0vQblNkOoIQho4/wYIA/4D7
P+UZYKnjnROnUggc/V/VCHVKm6+sgQ4bhLfozGm7zlCKvUChNBPw9fjjXVpxx87O
/0qIucRorUo18/Xn/9KBXZbn4SNJ0KbCqBpO8ncIqPek/PbsxIVsHmbZZ+hVxAha
k9J8FJ9Wk2MBCz2+G4uWt3XRJYcma3Ch8OH/JkbdQdxVRqPo5CGWAUrGnxVIEv8a
bJbOiN1g8AYGigqCPxBYNnwD/vqtt9edwZgOw7+xgIEdUUZDEhGt7vGVDpldeLnR
bvrp0VvaVNWxPLOdozhvZljQKV0bT4ddRMuR7vaJs00RroFyMEhKQM3dBkw5SpXo
YsS5/el49eDSZNLVQ/bBSSLWoN3EJCAPGp0h3/kQQpCPx1FU0rljjt79r3IarR6+
0EI6SvwVRP20m45IQF3iPF4c9mDIUv56AMaf/7hdCpkIaDHCWITYwbj2MtPjzF+A
7zQMSROZ3FHjqK/YBetzdisL6yQgCMT4MfUZfa6k6nLC18tricBn3oCaO+BA7iVt
5BwbgAJG9EUbqs8/cfOlhtQ6LNBjkGp/PFNXOqBRhFZDqHqlz9kpWXhUACrqx+jQ
JyjuCV7rlgl//wKxzR5LlC04WttKKtmb/NSLR7CtpvNvVLJJheYfi3dItz2rbc2I
p92VQ7ny1ul69CLd4Kgs1/m0k3tIzApL//ncVmGT4cjFnkwsz0R8ZFe0AvXTqwGY
ECrodzEQINdcjj7ZFh1YySj0Qhqwsj0lvK7EExD1iiarxBpDjOC6IG64DOFxVTES
WTbzbauyfQo5QDpx5kgGMnIe8sIr8aKVswCwAG6oQlEdt81AVjEz7GgEKJDke0t7
kJ9kGKxN00dZM5TM2KTFNJ0+sVSH4wrOqK8/nsHa+1pK7yitDr08rhDCl8yU+5Mz
lQeyiC68PJhi6cn/qOA2K0nuSci+qLy5JgGdsdrcVuC245Z5DZ0EEM/K2qAyUbsS
RTCBxLmAqY4EnRqfLlKfG4nFNOAnLyb8b1X3K0PMDexjGajU3nKQXZC1WvDJUwcp
YzQprqQaz6iZxXkRrg4eahzqPixIU8aBYtONr1CiqY0mDHv7bxe1dcZFq+pUJ7jZ
+UcFs7MB7pdLiXvAc0yKgad7XWI8yEJDvmP4iiAspNh2ZSpC/+2QKfxsfWdWPdDc
LZOeQHdpQjPRTMwx/dr1P7U8yFQNNy4gPw+Hqucp4iI6Vm1MbLBFINvlE0bc116H
z9ZgBHfRqsOEmjYA66dcQsqXheE2yeiOUfsDqkh4gvI2FZnNl6Zxd2Jhe9zgfmfZ
+wLCuI/AWGdRX50iFZa8iefuA7qmezn04Jq++0kzcVE/xSQjJNMaEhM3NRz+NNUE
4ZPhBAKUkQhRH0zDRR2Nuaqx1oZR0bEN06jMrHuHo8Zz/9++67Qo0O5gcL6GuP3l
nepINQRsF7d3bQRQLpQQfFfD/Aa2hOZ3lh3lbHs+b0LsbzzWJChss8V9KH9F8EB9
7GoyK/tEixH1mEHbTddO4olXQR2JQPC1QEBqPJOtLNandvJS4+erD/WUKCoXUhRi
sjtqcaFsfWYw8P1E9EKqbG3MdsFOcykBM/H9csDLSpUArejcljLVWCVLi0mBvngA
yNQzUk8FOSJXjL+FIji4ePWJQSVxL6C4R8c6BpijUAv0zz+5b0Kpn6O5qo9agWy1
Oq0aUGRRordAGFr6zKqtwAWQWxBK4OcGNfeANQePRaAUa/QTGjtCiAoNFMKWZVyn
+KmaHT1LVI5HEGNsNMQViBrpN5E/FGKBiCcPKHzvn50OvDOhaSjO9SBxOndypp2q
tjj+QNk7T5/Bw99PAZFvQS4BgSYweidmaUaN7AJyyHMV4eQehZ9S/ZeyxykFhkS7
J5cqMJOuYgG3Ad/GKBWYZkwEcdf9DHyh5Dl1nECqi9RoW9WNhAdaqRGuIIRK2fhv
db4noBht4mT/Lp6+raXGSpSJg2jZYlEQHvoqFEQprBW6iXXK8Na0Zx8kZYNeyKEo
++Ldjx2fbIp3Z7nZ1Frbm3M5yvkn33QkJlU7HHE3/lV6KdnhJpLQr9rkkC54+njp
uS08Ge/Lwu9zm7cGRprxrxwwcNQXWoNTEh/2rWxm624Wkz5TMNkJRUIw5aSowhLl
u6JLdML0TFrOLO0f5b7wcazDq8M2vxloFzQlyGy7D7SpR/gfj8nHVRZZvlVpBXZr
6wcdRvZiZ8Np3IXp3zyuBAseQ24pOKmK0viM1VCtqd0KbAaJTcDn33rS7EWQdYSH
L3OJAs/ht6nP2Tx5BSYQPW4Kuc9JmpqfHX5gIKwI9MJOjE60YE8GMllfhBjUCPoM
nDKILFOPxYgKHyh3bVUAWm0kS9a/TKucRXB0RpdWHytt/yzACj9eTyG+j/YskZdz
2BWwklXzhVOqO0MZEopNP0vUA+xW7i78L5d6PKVpPccChc6ooSc/gyUnTvsUgfG3
QdQ89K/g+hQ5/DyYXVxFHAfBzPvy82PMu0+/rEZHZms2Q0SrJEUUh97vLHJIqDuG
8CvqLJHD8xDLzfJKyDuJoEGFOc4uTOJymzGWBjuaBXi+Oeo5r+gxSWAYXsNwmTb3
iTisbD1zhy0K+1NLsBGfB2LYeJntjOWqJPg28ZOmUxDmMWkA4XMBWWJs1MbH13rS
SMUiHVEZGC3twKXFPyM2KuidvP9sqbneL9ELEA7zLo1jdzewgdpxdTyOCkuL4jTJ
KPiKtHxUjag7AWmW8Uxee9+uhNkb6GT5wLtfs5MA6VErus/FgdhZdETo1JRiEN/G
u4gOVzCEorvBfWA02UzLFJ8eN9pbgotri9b3yc6EgWpzwYkJjJwIwjCW4H3/Knue
mvMf9XksHmEDpFa27/YRJfRw1tvyWrtiVm9dtR6vOjGJ6g6rkyfwHvAVYJtDnlPI
TeRyylJv9M5YgS3RMHWbCV3VwmzJAyMLlcT/wupd4fqVrO6kDw+z9IuICldq0MPq
qy4k4gew3x0wmwcphyeXtB0Nyh6ZVJBh9/T6BEq4yYQxtoBSOJ1hoEyTof8gaHsl
pIiWerZcZG7ATc+5oNmJnuhttztEbvDp367Wsmh5VBzRqDY7kQDY7aE5H1ujQByy
T7ASGYpx6CwzQNPEPpSXp+KOkIJTbCMFx3/Tpfv90uJZj0uHGgGcQZ8SoP4mpnOo
p+u9Q8dj8UtlKl8nC6n/zvFFRO4x6ZbjrQXGjXbAgcxd3l7at5l21aMRme+sNWu3
fdLoCMdAQ6WFrBlQiIwm1VZoVXR8YSa1LcX+lrXUxXe20yOW9TZCaerwtUEUXDhQ
+JrBTJAFHeDx5+BICldg5sjy2UWyglP4Ey6pqF3sOVzLKlQKfeR5HgdYVjc4G1YZ
70tzQWkpTh5tJTQA/vFTtiIdwHvO0dfQ8DN6kt204KYz7Gs6FGYzpYzV8RSWcBUX
o0URs6ZUNqKbdT+aDPQbFf4hjw6L8KgVeX6/31vUPPiUnjUHIO9iBqqZSpXQJb6l
IBVsutqMfs3BN/+3lj3hcTpIHuxmSPkY8igRMQkZQ1UEL5F3cSOG1CouX6xumv+j
d2uoWFNjOares4KcNXxc+LMbm1YNH1urhTJpFMQjdDnhKLbECgnGjStc71MqnCwW
QuFq9j1dfjIli1wmJZ5ABoO9enwXgyXt+ifr2+JHUbpekWxyd4muVNG0XC6UZTM5
1y5Rpjy2d3i757n74jVaCBgB4LQdSIDXiuo7skRnQQXRUdPbwZcSA7dfPu6effrL
aIhxhgvhTQb4rrD/KuSleqTB4mbNWYjx1bSM493pjccdinf0RtyzUngmA/b1qCMh
FZofCc7Y4b2evzPvJ5kS+gvg6FFF03/d4hZyC3+pMCm5MtFAXokn4K81dTQKgYrH
k260xYrArzHy8xi04LHj8FikO66i6Rd1wx3R6ylLXBJGN02Pr0Sxo5uLM2WODZc1
Y7uiExyE50LlJ5btoEeQohhmVfQ3J2w9XAUkVwZRR4w+wDOEeTvwzacQDm3biQxj
+hgyqj51cEbBrC4AVleShl5SGn6gI4+0uEWDNXQfSY1aA6qQR3JCVTXRCqw8/SLS
SBT8ro60XQfqOPG91E7Sh7KYIdnaAvTxVNM2rM4O7jhogz1Iqr/glV41Mko18J6Z
on6F2SHLpGt+sqiUtyvAj89zKy6RoB7sTAzu4jTB1QpOPALwYBH7LlUFFKBwfQm5
n8qx719zVUUnVa8HZvpsm8wmpc8BCYUcyWT7hjP4ZA0F72draaa00YgrAVsJYUZC
v+M842lC8WZiiWbBitVPyRSh0Ssz0+EWcoxT2OR3/AYX5+VcHh1Xpb/YjoUsxDD6
5i7FUltd8wuKJHXhdA0dnZ09GEBeTsXge+Ff9LylPr0hJlPFH0mk6GlxXES2Um2U
4sxuPOENwmh58VYRC6WH5kiJgfOAngVv/BL9ticCNskvoJ03unCWOLwkx2nWtnSt
Gs4RtXwpNTBHlyyekaT/75/cmn8H3Dym+9CJYK0jsWlu2NVUlVYzBGIh0xuwC7+6
n7voE4RldDHAPHThPUaHNueY7jUrPdbcfJuln9Wy4m+d97DICOV8SUrXSxEvVhdE
IQJZGeWZ7a6kwnvWvg/UGG+I8fwPPzMceS4mCyEeUfshdH1oLTiBjOJw4AxNdj4e
x7wmg9VdFyzP5iY5Zu1j9yH8Wx2cHXWzhHT9Y8O2vYXvSMIMv3tVX328DuMqlo1w
bWZYcAM7HcxpvjZj0055da7Tbx87GnbfdTAnSI278QmNZDvRf8OiZr01BApRpc3y
BvLB4FmFJKct4mv83UIzx/XfQVOYlG+HR6bNiflFNggIYFP1LNRhpkI6lFblu9Yo
8zX10byrKZ1jpf0+z3VmLWoh7lx0yKiQC8ez/TQV4XzLqAPy0osFoB0JAnM4t3vR
i8AdBaYXiMKAiQRwkZQHlVIytaCKm8QiPn76v+efMGPjjvXqUv7WUieau2Ajbh07
BvVGrxPaIuClgyLIkWC/MXWXNiu7ornvdd+oE0HmDrBwEIbPi7889GICyxq4Jcni
EMSDjHkMYhEZsMgjD8mxf2pFpoaY+SB9pvU6oKKB27E0q1Q4rOg+PEUt6u6hBDCm
KOaoijA6DY9ovV3hR9JlWo3Qu7EpkfiYbfPYba+WVBZHF+42oiyCdYK2R/9MOWIp
SZbLwPJm16uioip34Z/nUg9M/Q5LQSPGc2R2aobWUSiK8RpRiNpqhpgRm8ovDc8L
sIm4xnKRLJwfX0rpdcYMxrdIQutJLbwPSLLXdy23bMKx7IyzBeCezZpVqyAjOOsB
Jw4YNq4aaCUddWvqBMe6YnqeHdrmq2gBFgTTnAeQGf602bA0jDeq/0mDsSsp0Upj
0dfky1AxEEsXctC5VoVbr/bAUSNvkWLbiC5ftZwbqs7T75SJ6YTsj5pJsu00x1C4
9y1YAz5ZgMQhUwYPa7kzVTLp2NCoOX8I/vSNa5cSFONbbr+r25dw/Cp0AecK+M3f
xPf4zSAufXF+xvBeEDn7jythlg+Kfk3xWIEr1y9hKGiW99xfMnUTWBaJY+cHBIDK
vDFSgI7fdsjoF3La0cqu4jKR4/0J2hcWMxLi4xombYhqp69ZD0XSQ6DGQ3p87MvZ
CUW8+Han+b5mpK6SRb+bRGhGpkPMXj9iQqyAqkUc4v3j4gOXW+yIphHN/AD+DVq/
XByGdxaRCrIxS5GCMwlPXnBo61WRROvaLMTKSWzxvab349OjgdlBKvJvMxPl+c6/
nUTPsit1UF9IQmlsCvQbG2J52HTwjbz0As0zRzcNPhC9UAFDmoiDb0OiGUF44t1P
ZX1WGGCM2T2TJgmw1TT3/+UeUEiAR22/9M8NxNK6UwV4qyzQN5FWw0PFnwoc8aIm
FRAWIDCstoTJBgfngh619RcpE8N7hTL2k398OAe87m88Gb0Hq5zZY/6Ub+S7JFFT
txJFqq/GMn/jULrmxrOcHkEWUfTYUVW45Ox/SiFHpJA=
`pragma protect end_protected
