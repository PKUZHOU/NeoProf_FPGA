// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
oVvkNrzDv/mlAA1cJTxFFWnN3yhM2eSd4G7XVY6a5/08KdPnMKQfYcFioEIYMerp
fbc5bRCsPfqZFO5vt4rWQN7AHQIelaEl6ywazUnEGPxZo061SQUS5wxIBd3z8z2a
sbP7Su4KpE/KF7sOceFOFo/4IhzksIDOBEflyguuMQCNjAk2oBxo8Q==
//pragma protect end_key_block
//pragma protect digest_block
vblgv8iyCmnlvMy11QZy6jRhsZA=
//pragma protect end_digest_block
//pragma protect data_block
v2V7i2fFI9ZlYkgmImuVitkoN6f5+TOAB/rFpZyWgMAa31lXtY83IbC9zPa+lmmI
CjlHp4IsY3oF2yZtBmOV/TzIx4kCc8QTzBm2BYAwIS/LIfDytoosw4YJPpxwrQq3
wHDXyx83GfVzWrmblJvyIugPvwp8jYbCD3rKqbJD4oEANY6Cjcz35fHU81frelrP
ZOrYIeLLALMtoLQ1S4N+NR8rJU/vTdLS2FqhP3js6nOhZVTq1JJmlnIqj4PP5I1m
r0r3QQjN4KCuZZUJAHd+nmYeH53gp9mbl19WqsPWE6FprU1e/3YbmER++k/zBgMA
iMO9TyxLzEH5DwTTqUR7ig9rByRnEiuuf0GCJENHjF2ozR/Km69y0vOxJkAxjK6W
VERZnKERg+igg8GxG8uRqZc/I9qyGOVBAvwnMcNI69gNVAx7IL15zWv13WOoVdVA
9giv1DNd/cT3oAo6mKysD1tfpSN0TE8Ts4M66LbHxJzErfb6sO/9P5/9WCWs/6b3
X3yLeKCrqK3wozrORxmx7yHRMbfgHipbVPHu8z6Dcj57OR1y5J++Y4vNaErW3GZh
3QHtDIvTGbL1b0Xad8ZgqPAbdcOW3oohv7Zo3r51j5I9LmFpVTiOSizcssPMBNEI
uOjZuO0vh/fVxBOws5qjn35bsw6K0Kz7Et//M42FNPr/UQw6ZEX38YDy6PHFsNiN
Bf/ndeJffzi5Mg5gREnP+UGMwpA/QywjU3TZ/DBjzpYorR5GwY+HO41o0/hfKPhd
7zk4bYAsG1W1tOFi3XpSPGyr2NUTv2eVZL533qLQg7NqeKd8XYdDyOGXVS1grRMB
kp4C9I7yATxG9b5z3PrcA1WNqVxYkS36ciRH7LsbTcYxPNTxJHm8ZK/jSQFnnuK+
Kk7NUzMajx8NSD+V24yVum77WbeF9VoiX+zFAhHgbOQ89Q3O/bW47vHKM5YmvqMq
HQNJ+rhppaqVxLgna3Jbpucsvx5IeFirZAPAzsPzvjLE80ePD9Lkt+KIGCfArw6h
UD2Zf0A7afq2Qn3Ys9tPv93CkqH4xggY0l/0VYQHx/5Mn/uXu3PgQUi4k8m9yhy1
iBy6c2PS0LwBOx3DyLvQsQkaKgpi2qhYPARc+fCsxESJn4GkkQjTWpDB5ZGqUsMr
3XE/8l89CyQrBBOsg2Dbr7O17QbArfLevnApfGbilZ8rUv63qm1w9BbRRpUk/9m4
rtXTBHOqTOS6eUKO1FTTV0+q0uSUCg7oK+OcEk9GXB4b8HREHkXovHvPz49MZ+3t
LVNh489SRWubuCy2Yz39cBG/h8ue6NapE387yKBzubl6j43UI6d1uugXjYFN4nsa
9gP6jta22kMG67un0I8t4mvG4VVNI8ggokngAvClpb+/LTHr7G2JpJHDjB5y/ySu
xGHn6HeT/wwzfHtxXsi+dLSZfRO0PwtalALXtd3Fj8gJXuvN0gXoPWK85BGJ2ir9
M1azHVxTJArNb1tHRo6GIwTapyXgymg9gtC0v0Iyf3Tn3cZuvgcXhcvLH2DSmN4b
ljC5vZxFrs8hjd6OWNlmViUHr9UbdFHj7W/Eq3FepPZJ/NMRD+uBQH8XhNNpsF1P
upw5ywAXQ6eKwjEyGNqtoTDFdkzFFBkdHhkVixdZvB0qSDbdMYztlS/MeCpGnI3I
BTszvUdM0xw20IqvAEbk6kUXHw7oiShu0UZABQZ76Ob9oWBDFZBidCcLxw6lGLBY
YylJkVr1tzGiJsOJqDCXHIo/5gRwcIx+fsgj4ePW/nbZsnWbwFCzYomvg6gGCaHW
qBDqED5g9iARbG+RwP3XG/D1GQMPvnGbh/k20pTkTTLrS+vgZ+qbzjZkvjuwN7kB
ceMF7S+/eMPi4gwXoSpKdxex9mRBS0MADZLCBGOo0p1JtR117Mqz5JWfkNUMmx5C
zl3sOx0uwtHWlo6G3Uogxb6n+yiDMFzn20RSTfeZo3DjerQEcAEP/lWtSfTp2t0y
yZphaXjMMPNQaqo0O9mFxrkWCCY4QsqTqEkIkAt5Ndm49GtSTWWVnTkeQ1kxPqxE
lhXtGaoH/kmhDuuqmFgo782R1kx5VCIRAfp/MGAq3jA1Y2EOfIv+vZXEcq87XzSF
vpqx3fe/JbbPzaGWtzOo15MkKGU4WtBGAFIZAAOU/U7KZH1imCzZ3JjaMBjqNkbk
zS2B7TFTzxtQkgryPmzK8zGN8BciOLgbWWdfsFgc1HuRr55fAsJiZInu3SV5pOQP
3nj7N4/J6R/+giOl7Ri5bICBeNasjXUf7l1+yBNMJLTE0WwNV9OtfdqsQRywE0xu
ZnWNcwlpP0py+oOxZF0N1GYHxuPJe7KJ0faLORLrh+xY9xJZVuCM1cWC4R8+p29q
nlQeY2QrwKnQ4ncuLYUaldm5kgqR0a/Gf7pJGNp9NZmnpKYSU6gF79UaAYDfgWZe
jC5R/v8QYeYry4WdotVAiLybjKll5lOjUxMWqo6FfU0nEGzMHkGw+ioLEKO5VL+0
q1HI/zntrRvue0MZPBf/LeEsH5y12uIsAS+bxIVuUmNByLFPCqEm7g2PZNt65Rd5
FbcusMjQ24cycgSG4Bd5ybTqY5HpfYv4Og1qH5mn5S/EZRGnL2Q11I2BM10/ceDh
mDd2LRGBMPkgHbFagzNq3v24QBenZNszPVbMuljZO3GNf/F1JwJ7VPHqKGqeBeO9
yVnWiWXIeUHBCFmrDlE+Gjv9wOqdwuKTHYU8ZLXnE6astefuSw4t/Yvr8TGC0o/N
cFN56Im+HW0PqldpmJY0DAnll3rk38/J1j3NDpUvScpz7wcXcKwdDziIgH4qgfis
XeyMhD9XQRAvY/q0zVuzVftxNpuiI/FDa+3Zk+0ETCXOe9belZGDhbN0L0VLsmr3
KGT6+bM8ZWSGpY7bSuCObe5/ZbIQJ9kkAcD6d3/s/pQe4NBhcJm2Iug4AljpZ258
Qfpd18bNF+qLCMVX1RgU+TS1P7uqpZ0f1bXACSqW4YfVASshHNUaFumaj35zZ6k2
cMtVHvxnDeaSyvymozK7MCD0dMweTjNzTEaXKFsMLUaLznBI1g9g8PUCMX/9kiVB
bZCJG2yJKQZCkd/PbNhsiHRs4+a/nwAdaSAxZOoVDnl4gj4Sd6icBEwZH7ilP65B
48SnVpaaQ12ZmADGnCrJkObJMnz0dUoQ4QW3ut0vM8qtw92vWcroS0wGP3kPSoZi
WR4ywNLjPlaoRYosMjNPmoLeXdt4jTIHB/wxVTrxb0gkHKRv9bga3b1re9zLSBoN
KSueZlEtqujnT/YOU3neO8lmRpSt2grob1mb9PNvBfDIp4bWZop51UFUdngepWAP
QkeB8AepT+hcKU0EQ9z8uZnFQ/pZYjS7mcpT95WBkQoq0/ZnOePxXFGMXPhl25d2
4uM3Jc8tS3AfJRLhCSz4qYueVACMbUEqswJcWA/CoFooSJi6TNMflBJ8ydQ+VHHS
ZLxaQFvl791ffACG4a/6TvApt0wrLN6LjrW5pYYHkh71YO+JSm384RtXy86AUP3L
BpSlAeVr9dgqm7nrHZ+qqCPeWx039g8XWQZyoFMTC31zY7OiJfMvNKeXN1E/seeE
5KUCPUdAcAMtbumhpNmesCazegMHsU0oZoW7/3BxjlHky/qDxrwoyIfIoushOe+8
nSi7twx5ucGAchSt0XMmhVvrei7IoDG07XFxwA6OumJUiLypgcFFet6DlrsjQZ9/
KK6ln9g4aEmSOipsaA/6uam9/PASALanowyvs5UpXYho2SmEKHrDy/JJbC9VAC2s
Owuj6YJUooXU5EN3RtuXlt7CO8bHcMe2oGvwapqPx0hVy0Bd80d26oPsDViS1sB8
Ws3qgg49AYajdRLopXTJy7d/nv25V55cm81J0ZBs2iV9UqhKcFOjZhzOLW2V1pkZ
nGCW/lHgXvGEqLX5Yehv9TtjAcLW5o0UblVE8J7Ncwa8iCJ04j/qUbJdmArnMHhR
XAFl06mdL99jYJKoygMnPi89vc1AQbw5sHAe6iHNNbKvsgyy8dsGi1m3BOs+fqNm
u909nC+0Z8BXcTn1Wvh3oQgGfnNswj0ofxJO/IHtSQa94fxo7lU0iuN+E1TBjP2u
qPoOUcF9zoCsFN1+SQsRfqo/sM4JLm91MHO4B4VlVwwsZRWmy0//rmcjDxXoYlEI
nqWlYI3qCGBrrXN9eDMxXnAAxrHU9kXn5sFxDOa51o0pENfDyuoKDTTzwmx60uCB
8oyFlBnExM6odm9yVgM/E6bw1eZ9KgaHZBnigILLcKi9xB4Gs2jD8tsdDga96TSo
0pUb5x9AzT+QvI9BfmDpq/A+UgRcgSTrj+1ZrLX4tl1uGuZ92Smfw1e6DjxVL3sC
/stRJ6wjtfezidZ8Jz/HdluiTR8tJPwcJWPCon8Hz6IsrwZvqPN3yLSIYjzJ0INw
TN6OwfDzvkIMbn0W8cKCcjC6JNRohrOJ4EpaB6gUHFQKJV9QD8OdYjTatVfKXEyw
t6Ahv56u8cqZA9T7n39fHG5KjiihUg+NjMZ/Iotg3BNpDpeRc2Ze78xl80XxVng/
vA7OJHjprr9CndJ+UNwMXbglHlNwzQiN1nLbGEwNEa07/L5mNtbjtxfKKKc2SpIJ
OFuIfmH8u5k5AQX9VYsRY+AAyzIjAWHY4aL7/cS9YOpjb5Eq8wnHtG/FaZHRIKB2
668KU4sQPacL5RLtIdBDFqxUN9Ikp7fEtZHRhs+QQzOy6xK8v25pMAfE3b1/3qel
IhAgSC3xux90rsUkFOZTRFl74wBrhOJ/sNZ+eHI5DckylgNSleV+BPuR9ficcIg/
frttyDOXvKb31kMK7+UtXmqOGQ60DkPD/Rd0m1ltdiUmfyJlpOujeFBU+yoXi8Tt
EPFwPDt/ilp97w5tqoLFO/tjnJU4Qj+uU8yYCTvm50EuJAWiNiHcLNbjkEMUOWm9
YedNBn3wgZaXYswD48snIP4igVE4X6zio2rgSy/OQfUuQpmKWLrBPN23n/Qk1KJV
pc3p6fompVXisVnWNcXq+2quZotVm9TQRIlTIf54yr36rWkPSBOY7CxsuGZu4f8m
MFRVWis44lCxQmDcQklb/5RVNucu/hYNfYgn7Pj6jbT0eUpYWYEn5zk90pHvfIuV
QVpqKelaSFqy3g/rli4Vc8wHRUC7IDwkxLKmc0zT0T5Dnq+sQVH0wVzBfamy+LeT
lMnu+CnNQUseLFElV9IJna7qZhR+uO5r2cb+IlBsuVfqDLQkiBeLM/+WlbIbU1By
cruSkXetBhhToPDckw4DF+gOMgbLHFVaGq7sq1PcOOXV8St+MybMzlGvYXC7WC+R
0OrTt8rQyLw80upOVYTS0AMx/7z6Uc+BueuivLDF2orrVwfxwTcFnydpgA6CaRF1
rDJfqOkn2JYSGw+KD1NfImHJ7FgOUp+sW1Qd5wCAcZ2uXjSVk8oEJ84gDqlc93jM
euAkwVRy7yEBGh2UkBsRWUnFgzYVVjPr9jHnqxEhS29Isc+t7z5MJdkRSn7KgSj0
TcBCYOu5Zo/Rz7ySiIFO6ybXXpRyv0DaSBxhJpR5FoU6Mod/gywfa924EAyyxXvM
25P5vhiBXgfnijvgGoBVSF5+63mP47cMiLezIc9ezhWmo+SQOlVbgvsg00dKnJ1/
FCD1TcjpJUoCMLVJjyd8o5oqY3f5TOM/DBVWOoq6tE9m1pW3UyDv/uCrkfArhBM9
GzJDpfG865Msj4MDMSh7u4l7srRY9S3MUYuKSWrgoab4cZ9Wyrgu4pZQC5L7w2rs
u/QOw7PGbjvtzRVdRCjh4xVgundzH2DlZnyKTVlg6r0ieRtQSi5vdZ/2mffZPL7Q
jWhBvsy01BxVpyCBERt73nMEzdiITC7chGZJhKN+dRl0G10Ksr6Kx43LAUyLhoct
aq4gO7M/zITwHrjGjF0UMBegAOOs+SWiMGMaPT8u5aNqW8ETyZn7ZDLfrbXFsApD
F89ileULXelz9IH3LspinJszL+niJccXG+nmnE5gi1FnzrnCqYDcBZF0UhC3LdOA
Lqbfw7e9ri8uyTZwWZIO20ick7d0dxxZJIn0gVwA8A07EYRsMOr7EiduACvIADp6
M++SIsFMh3ZZguZxHJDSQjU9eioUFZBgWL4srqz78Ks3NcEESMiZuRaywJSjRLLk
wXhRJzLVmfHkeqVH4A7bSVszKXh685SS8fnyFfATw2jmmSTidp3hnt7RWxqg4QQX
9b56E3ZVVekxstB6jrhcLyiUjJ1DzbHWZ5b73dm49kxuaHX+fS9rl4wHrwmW1Tmv
i1On1RVL8x2nxExupvW0fJAfaGskHWFNcZbR4lRoGIMwtkNQ9jrcy9c+wJIFSExc
NakMustojw9CH7p08wgSUhnA6wlABmfhG3twuYXfuGsUfOKAmiJbE5L+VMCB9TSS
oOSHgZrRJLdovFS7/VJk1EFEeHvpFNWjZkEW2AoOIpaiv6kdoqRI52LMEaPu0utW
VyK1FPPehglQ2qdwea67+yWVdpx7nOdXNKg8WjCybAEbfNibE7kayeR13vdITr4R
ktShGCk2OTlu027jy4YXHFRhqRlKENxa3d/KtzsgnLRsx79B9+noklyV22cZi6be
CJcBvyPxabX0favaTG5nMLjJwJuQUPwd2UWAsxKB+z88hLJVSu5Rw1eski+7LyHT
LcR8T7zHvxdtm6YHRDUm25PC2i0Zl/x4ZcJLX88zC3EuoMHGCq4PCQ7pHsQKb+py
q4wR2MDgeysExKsCTfgih5eVEy89KizMlhypj54Mrz+oYTRf01QjmN7fxZ0tiwyd
pbu5/DfrZo9tBMjF1mVZ2Hq2vWX5ucputIIIA2eBywn7rx5D56sAh3rlT3rsL+1+
VOKvW4+GuEZhrS7F3Moh36H06WqlknpSkM7ULFsm332j5cqvjBGlRrYGjlCoBbcN
/zANRY/DpdvZf6fT2CFnnvhc6GNbuQMiJqe2Q5fR6TYkg5y2YPVQAm0QEDcap9S+
9ePoMBUntbrovB1B1zIGbKGpOrae/hh2hL2KGmA4PnNvcgr1pI/XWsvHIsciAUSj
b35B7dokBAZCkM9IA4ovampLrRjmfSTpGUqjP/gbdq5VUJwt+q4u0FTvzqojOCDO
TwcPDBSq0epuPq867WcQpxdArY+MUY+xB17iw5Z8SZaTckTOy9dxewGEt2oN36Mn
+pHBOog8HouzscSbUbjHZjnBZddPR9LmNNxFN92vvbLKCwdOUTRFuWMMylFq512n
hWrl9QS1gUDLXkf2PXgPfb+cwvbhuj0TXtYGnyY80zy8MTuUBSNDftap46wOnfRN
mMKRwO4sN68Bd2OvjpqgqeUNLox0aMEyBMFkr17Rahfo2jDeKCtjF6DuIRpGHsI3
yBVWsUQUvGL/hX8wyf16tC5/8zcCX5Y1CRdwN+71So80He9JCwcEg/jxHiN3RhFS
io/CA71FTfbDVMWOsRCzTdL/zrsWdYNH9x/kTbSj6Ib/4WY5E9Y8c4TZ6RIPHDOz
QHH3rX8jgor/fphnE1f4j7R2xY7HpGg+S1faWfT6xxer52+xbm6bORJTNKy0f/tU
aTm15oNDrK6uXly7tyzo34AyK1xX1M292cktFM+aI+ktdFYvXUTG9pubmfL0e/3P
nqWZcOMcjpIR7nDNrUNsaUcXG1iddPDlUV+0/PUboHA9vwXU3ciZItzOr8k9Rpo8
iTCaCfmeA3ltsMWG4agJNoRbERGmF4aNoDxp4aF9eFC9c+n7tXstYEQ0WR/dsSzi
SxFvIIJ2GUSuj2NjKktVz0RT89eFCd4pC81Ggpe6aX72lgBqxI9b2X/hAHyqoNEv
84/3m9Eqk4RzMXfSCmG88bb3sSobnQ2/rkciZB21MYNHAui+g1qEBiGXNOL4mKbg
lLqjJ7zQxMvnk3J77MzDEIFBVRYykZnM0njWU7hx3KPDmB5QhjKqqvKuyWzlpuV7
rB/Yiqc91MkAbKGN5y7VX9UdfY8mHkm9NhwUztZuKfUUPYsAYZrBqojjbfX0lT0d
i8v6XCL7TDdaR/dk6rGOgRu6B3dbXN6OAKEZUcyQl4JXxh7ZedjDOj28LAH13ve0
HLugZj48ezGpF8qJ+Za5vA8V0pixCg8o6c5jmXq80ovVjk1gC6wJGVt04wHCqENZ
9b6yN7YB2XwMDat/DvY/U5UBEeaxMDnO9YpKN7rAKO67y18bVGBywcDfhrTWikYq
Bl75Rs1Gak/yQWGdR2yeH6nhZJpVyRne7V/JrVUQtqmAjSWKrtyi4SxeIsNnEv1k
JiurisT+e3i4DGde/781danyJSFoHN4cDVXp4IbOegkMUXAjb/sIdUPxaZEGX3CT
59bxTqw/bibxQn5+RApNzN1sAfVIkRsw57Jt89fl9tIuvBeaVL/hz5AMC9HWJ3gX
+wZf7akzBouRw2MwVoL1fN7eQxTWlngXQbwd1LCZkoP5wgDAPkWgYGtPx/QS6Y8a
tdV5qqaMGu6ymA7iu141e6aybvHqQiLtEx4z7D0UfsmFUXxMRTfE1Uo7E4tx3U0N
txlO8Bt/pbSXt0f79rKM9WgPNNR+B+s2NdJp53JjJxgnKgGB6c4XkZOkIsU4sp3E
T8H5PNgN+H+IkKGNwi1son3kra6546+oQ7kiPSmuGx22BQsVFC8zXf3FkgU49BeE
maE36bEpu1D8X3dm/yaB/Q91/+Xg9NQe487ZcWLh9aaw/xSuFcUkx5n0e/ScKQvj
ipHizYmf97IgVadgQGyswv31heVvWS6QzC2f5dboU9Kwiyzzck50mhDZqv/LlVh8
ZPQ5aobVVLfU99sKdKQ3glbnGmx5geGryqO7mlwN50+aQ7ryk6DHLci4sUCl4tfQ
OkbqEO6IBZ7dDl6v6/3FVBzvgpkN+kxkSfIn5Pas2s+rSWf2XBvpdPTkDqD0QuNQ
+xgRXecvwQJD2RSo1ocdtCUQDgTkv2yswI2dscPPtS+5Eo38hhim1r+KKSdVOZr2
jURl1pBbV+8h4AVY7nmtNHSvuPC46a+T/ZcFIUW1wIUB0/n+hSFX8VOcGQJnV6JZ
MBQjcDaWNG7c19VG0txTAHmppREjJU2sUA649UrizydNZalSQeTU2QQpkprMOMU+
WSKFE4titoJaUDOf814YJVZBKXmovg6EH7wcp9rHCX0ZSeuHEUf5BWuVETYYuLZT
fN+0/rXfUQiwiXPHogSiPchNvuh9XoV6lOdoiKzPCsunTLXyzP0my3v3i6h7lJpH
DTg7juf5A2NoG3WgiLUb9CzF+IZsq9CnAhCkoALiMuGG5OacJpkdLouWgm3abqrk
mHkISsVFj2GczVvXhSMF3TcvPXNOGQqdwIbD3Fs5khKPbXir/N8p7L3nLZs10DGb
ZA0rn7C5FA8A7ir4cq7GWlr+mXcKe8revHVTyxM+9hPnbczEuW8GJqutM+KquAop
rwdmExGBWn6GoVBBR5LkvMWCo1irt2uZvg3Yd/G8r1iC47L+PcxDp/878ZnB0j+g
9Llc9xReifZBtI1ysdunnrFFt4PDvkeZ+bFy5n/XVFXPIjQTN/j8QuzSIp2//exp
4pjkzYTAOg+wqL28rP9u18g1zRa4k8qTMNEy20PEw7MkD6VYLjGGv4eN40Jlze1R
10wBkkN1Dmbp7EhYRuHmKm2xIKlp9Ruu/TGlG0M65Vmx/PnfhAlIfWWPfrRaEOug
85AJgmI8udajX3v4Vd21l9i2fBbUcQ6DcnaRh7Sg79E2vDldMeGNTcSDPdzHWPKO
vkyd/qhyAZHVlNxgpHf1tsdGXvGOmIB2ZmQisfzU9r7pdNMKVtR9+rtyrhJUEOyw
HgGGV30NnEl0SLvgyKZ7nMACWC4skhOSYoU775wREYulp9aQocVsLo0G3FAm7Cgi
p95zgIQZ2O4dHwGiZ/Sgef8AVC9Ufr49Xul6OuGlehzYFqPQL7DAOY78VQ2oOCMG
8a1ciQGeEDxRi9oBPk6b51jxfj7kFeyYGffd03xDpP8BrencwwXKn1VUkx6hjSu4
63C5LqEccCrQfRCRe5T8JnMuQJ+R/zkcgxi7WABEMTP4fxTWhXI7tx7grib+YIks
95qYTKiT1044TSOfonA3EY4FmenV0u28QoP97iuGEHphx0L+HYKGyFaej/7zu/cI
ZwfPtUIOxx/yMcnz0b5YEsS25q+Ibb/yAtcbQW4QD7Q=
//pragma protect end_data_block
//pragma protect digest_block
PQAs8YRLS1ZvOSaanWPuDxXkka4=
//pragma protect end_digest_block
//pragma protect end_protected
