// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b+2VcBcdLFqldyQyLRkjtBpTDfFNLzJRBRf5uEtlZu8hAMTiYI9BolkzKujr
q1+03Z6Fhp4wt54lXLxJ/2G9SQu6eqhs5GJvpe72gEbsOC6NLFdGw/eXectK
iZyrpit6pRD0s7nSfbLUVL49q9PaFHqmuv58sGUEtsQ0Bs7FKVG2bsfb9u/F
9bLuTlAgYSA6UMBh5WLkS5oZSdvBiPJLFKbZY5JuMp8GQioz5OHYOaNZtT5W
NlV3z7jRkJlqKDXr+2ZKEuNjnvAAq7BiG1EY4K11AewMYJcHYyAEhxk+OmJz
+he36+3+2WwyoCYYlBVppvtQA0PdV2oSA/NeMZeQJw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
d2cJ7L7chHIYBAAWqk+31/FZkBRs3IY1c61keYGaBw66IN4lxkRwkk5cpfjH
TUGZeSEeFx7L2Hw3pDAF/5+4dkCGVl4dM4KZn+ZYTPtNIhLJp4L6E4ulcGLA
0DLJewNb12N2e+JxqtdPyMDgjFXcdMNsfYCuQYBSXk25C38xA+hs695lwKAK
pX7f0e5gH+UJYC+3NVe6TPeoGLRwus+o3UxxsXV6zx6LmInVdSuEW+eYMRva
fKctLoRCFSn4jcUg7DiMCoOjQHBrpB4ojQlSB6+UcRS42fq5D9v1I0UxhC7k
KvGiy5+Vaej06U2isdcxUnH1m83FAvvjRh9GtkzpMQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XAziwfAcHmEF6OCChHpCR7bfLUxAvDzqXH+5rFGQqfQgCkSpnxb4Vl0BsB4f
kaCr1qYbIXZils33yyPpHWVvNuxUB0EXDWm4TwpX2pv5le5016zdHE3A9rEd
HoRbGmV2R764ywg6WJkpG2t6lM74XOhwZ/UHsPSnMWMHHLggZ6DTa+PJGiuS
cPi4qfqaekKrAJvKtE7ZxRE78X3ZFq6IYmLllvh+wXSGqARgnDmZuBQXARBn
y3Mubm+H+fiXwOr/kpZaau4bU4PUTbFSERIB+CiGB+xWg8IMW5o0x8CSiUpv
amDE1EkhoZZNviut2gXiaVhu3WcLIg4Ty0ETO1AeLw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
spHRFdVcqZaC9NeJlFgD0NPON76BlEFBUmIGiD7+1TEw6qwqTR0OqkTv98jt
I5bmAv100/NwQw99tvhomPgaWKMgupC9EuW2njRJTSV7cw8TaSnxY4S0w32r
rytrOQlMYoTr1aCIoC172x15IuohNImE2qIC5d6Qp5I5gPmzjfU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
JIHp3KXC963vPZTcbP6S4m/TLyfNM9REauuNbEn6Qfl4PsuitICqZu0CIFWW
sYmFjs4pFEYjUFe7FvYDgG1maoGBlv44/uVSydXFtboQpUnOc5dmCBuThj9f
WJkSdNIe26JO/g6FerfqaNABHJYr3tebeBMCFrGNJZnf5klubpojh2y7u49J
WsX4J3wQ7OKA/5wdXC0n91PiabFuFAY9v8qG8IbxzJrt1TucxJC/r+1AGZx9
eEyPDBtkvHAv0+GuAFYo1GjOTykcYfQT1AXQ6fBedFCQHQYkmisD5ACduNhO
i4CE59MXsOh4FpNrnNL/h7RdGjYJSVBqri59GaL2hXCqXidFWMH0d4kzXy0s
ZkDL4OlM5541bF6pHRCHQWa1ty7xM84uU7ijVU6B8d3gQJYZp79AK1BMns1w
faKppq/IBlBYfv17uG1pFMcjwpkQ1//rd6Ky7mu9jxVXVNQmBS4paXsFWKqa
tgxUAtM8MgD5cyLHZRexcuj37bJjJfQL


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cCIYOU2mOw5PyzxqhGEhldOM978AN38rMR6ClqKlaBfpMi0J8SaRw1BBeM+B
6Ef2FAPFP0OR8XD8WzUD7bO43lHT+Bdi4Zkdd2xqMzeGXnGsUre4WCvwgIP5
qd163moeeZ5su0oCYcWtTAS4xHTr79FjHvIosyq7cj5DenaaTPE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XWZbfIu2ttuRTBa1+LQO7HgHGogbSyLGiZzkosPV+m/1DpXejhiwzyX+Tjkx
pqqautOYy5/zpw+zdGiYPQ2bODQp/cdsSMFUuR4y/rdbeJsUdeKTK1MFajZX
wRQi1PpAPAV5UeK+BbPSc4zZQBNPDPBFLvRCKDX2QX6cST3HGa4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 15088)
`pragma protect data_block
3xkiarTudt5lomxEISnJuBhgePnPaIwhbqQuYD/RwjL8Sr2UFXC/EbD/DGJZ
SRwiIBmq5OFd4QSHE2NY6iwNG9HKl8WpU8OPefEefgW60QIiPhOoqNm8fzz7
JGmVhq8pVp2SdQCmA0rZZdYn8KCUQmPHLEJ2na7hf9GRH1qQU6zsz5AJkXcu
TK5vp1qdyhxpWeu1tY3dttat401JR0MhDO94/MQi/sywzrPrqBLsP0znR3+N
cZzcuyOKSVmibTO/0I3GpmNMPZVeOnc1CK2tsfNkm8h8+HX6whWUGmoT2b7l
vRVlu5Ch6E5+OaWitKX/+TfcCw2b58WT0Zdp7xaZxr7K9wS0GJOAjVKR3LHR
5XSptwBtw/d4+Joav2bLRHjIu/gEKt/avTnK+3MPS90tNIhHNOsICbfkIVfy
WFxy+wonKbdHkvHdX8Qoa0a/4UzwkFYpTi02bIHtsox/nhlB0vst64Ua+ms0
2uFt9xQ5BV7DCy2+gpRsvWd2MozFiHucvL5M3cAsgw8dnvbatIqQyTMZMgoR
SyzkeB5qu9IXkMj95zj6PiVdo8yd23WCHnIZRPb8m5PFLto1JsjVN8WkOPMT
IhB+HZu+bZSJRckueamp8Zqxlw5P/UzK7yZSOoEmTYPmhvb1Ujb3QlNOGmdU
TIJMLpEw37eWAe0R3DZUiYBBi/OVG5ggtNJa/5i+0YFuzsgDUdGd6arPj+m8
EwTePhQec6Wt08sVb9Gtgr+T9z9j/4PPl45n9n0AGDAUCotnd/z6Au8/65RG
VKYqNdCMkWS4knpTmiRw6GdQXVB3uCwxHu6qn75aA7wF3ZPze3wV8CjNso16
6qdUKJ/i2d3Kybf2aaxLPzXqwHIDHXey5cuGTalZ7ttl/gpp+wNyAd7GiBuM
DcqrjMPfDDsxu81gSXF7fpM1qsSAiAlmSIajfAsOEuBtKF9Ith3gUZoSqWgI
2C9/iU4ZCDnFzwiB3cAssZd0XS1SrH2bjMtoFPhq0MayPHB10FEWm2hCp777
NeRm/0uBzExrtp1/LF3u5PdeBR3OuwR0Syz1ljIWsY2rD9hoTGu3gUjtRMVO
YtGcc9SPHaiY0/cb5U5GIPVwwlviLTZyPzXnNeCgDt15f00VZFUlUtLG9U7x
IQZTCSIqVu2UT46wNJcJsOOX6oZUfZpDBcfkiz31DzGFjtJOcSMn8pibt0b8
pxkbLIeCs9f6hpp4x3kaCI2ae0hDsbY/dSZ9wuf5MeFfzj66mslCG/tx8hCl
oSIwKwm0syuuYfjRlPpgU0xJg5k8RRCusWI37gyyXbmcrH5c9xT9ZJTfOpS3
2DPmlBCMGLUA5nQe2O35tW4IRe1B9RpFIlCFcXNZm3f7MgOPfAfjAvLumhER
E8tTJQfk3ZV04Qc9lhuzW44wrcWkA0aNlhlH8YWsz9CicP6SnzvNn6C4X/9b
PXX07ThOy0KjXDC+begC/cxFiioxwrVk2T7flKOtcoNSwwiCuJNHegLL5oQy
Ytl7vTOUepIf9Ddnm8VExsOixwsPwUEpj156eJAnn6lOawPnrWLgSHjftaGx
n36nNjEBhUu9Ik0NP0qqk6+qBXkAG8JNz+XDQXe47kHHnyT1Wv+wC5NtR4f0
3cJy/DUKyX6YiVqOBktqijVKYtaDDi3RWwv11nBy5vewXtHdCnTFG1dOMIpB
iTExhQ7T0QiqDeaQTyWw6Cv4oB7A8rPPAsosP3Wj79OWGLbxVGI4zV56j3VK
RIbUgBq6aFzFCE7MDc9lOMKkpSEPOBwi4linapNiOaJb2ISJBNFEBemEkSHs
RTsZknHSnDxgiE0I6RYmTsvPX2CCnQxNNyyQYWdVLHNTtwMVyu/AJbOXMTT4
nPa8nOvc8DAB1wjU76I8hLmQ0vJOHLpGlVsafO6xBx1nWffZ166rXQZ3DoPr
0I4neQv3nNKYmXtrELvdQ1Ja5wnV3XBFBs9aN8nyXY4+zlDoLEN2E6ygIUbp
poK27Yfk+ddYF/NBodEFoO2ykJk96hWWQ+37r5uAT8221nXBaKXatboxJw0W
A9oRCqkWWHdQpKwSVKIJi4+OoywS5z3CzNxCsji/H/juNRvyNQpjPJyBfDgS
S+JTw46KNaq9MwsPeL1I0tM/EHbaiQHabC9zVkT6f8KY3En8cdiUOwKHqFM1
ERROEg9m3+9NKHltn815soehIZswvSWXogiMvH504rG+TwD0gURH+Q0EThxS
vm0Osg/eHa75cbXxuFMeNAH7AOu8Iq7anmROcLCKLP8zJ/Nejq0LjeKwP6U1
dvrrOmUkh4rW+E4GaxNSjI+7kPmWdITDWcHhQg8cvJjoi4hDdjKYzjg4Zn9/
4EV6cTHbjJutpyyWX3UQrT/jcB6HfdfvGKDLkmeaoYXgxZFSemCJNz3Q6eYP
gdx7oOMCNmDVircG1249oAHhiNCcV47yml1pOwzBEl8m/RZ2fPq6rgjxbThV
4peUYi7F019dLsG+NJaLoiJ1rMLzllBjxYyxw8jzOhNVckDHE2VAaBl7jiM/
J0JCL3nSPLAR98/Z3t7Hh7XQoqILy0iSdPL7j0FbNG9XaifAk34Xkm7qyCkm
5RL0xy+9JJs+Q2v6Zv0jFVUkjplAfjCsMhFU2lp3IMbq8AWASVE+yKfCwWXF
h6vnkCI30pmZppk4y7y4lqsrd0lOjZcjVQY1BIllL/U1/Paf/UQJzWP2mKCD
N0YPmkLmvlAOp4MX2uC5hNhE4sP0K6smQBA7zXQM+dYQmhpqwAC7gEhO+X2f
31oPrmMTWDoY5ToB1j5cNZR7L70QhNVDAd05qC3QX0n3Rdjawfo51skAcQdt
AQsGNf4yRmEavR1rRBHvZWIQBo8xAHZ0S5AGe8hpJe+T3cu+BtFRcoRkkFr2
eRiblUZjqcdsuTJtz0nt/9K0vAAayD15VTvgE7UTUMUhcFbFX91ZatS66P5W
CvhOcSxsBuio5XVrfb7Uk927qTkqVO3/7NrzjdmU2/sNifEHNp4vSL3nFPWH
xQwXEJs+d3FSZBTYD/ljE0QzFOdAbKNM49up5Lyud2CEBpNO9uZwoVFBCTYk
ySpxQTdj0kK9O9fVFZAmrNOhi1KinFDxk3d1xrIVoleEfg2yhCVxx+7g7uPR
DBGEtj6UAqQn42c5VREZU3V0aiDJjIECzmM9B1b6TGKykcR5d2a0Vdn1MB3C
+5Bg34qjibBLXlzjkx6ePcesHzPlgftRMhJiNYMK2j1qgJyuA4xvK8ewqLhz
rXaJO8H0jfMz6oNju3hJeylxjQKNweUu4WAOFwZAD/p1rMqA/aKe1j1gJqmi
UgZNro7e3VgR+4eoCdvSiUNkWlnKcJQTBh1BIHzrODmYPMey1c7BHGn8u97M
Nm0udAFnVUaWy30m3+1a3hkfC3pC2fe0Jb1YXzMV+sLpC0dbOgkswCczbAA5
tEJlR5E+iIKT3DdPAyVXM62B3D1Gu/6LX+DFkCNr+yd46VFioD9LL5+2eJs4
2MFx5V605NpD4HSQyVm6fn86X32lTIhHwb06fs+BOMUIWyGimqm9IUUi0Tbi
iE7FMkHIu7zZFVoi4aW3EyCaM9AHZjA9C0wm7eAbzN/xGJtTJsy4zIgqH83W
OVYmYE57Wk4GjMr29bGHQMUIz7F2LofAerzmLiKUBYmIae7kaoMcdDP+h569
t6iewuK/d0+Zzp+QVUT4AfW8fCjoMyR/rjLiJLRnbM/cFfCKudWLEb6QeU9x
NYX1s6Mo14D1D0lGuPqRpXepDclj7bYKq+44HBxr72LdB67D3HcbAZjm3Z+A
eIQ3S103la5v0wVzrzoJJomeRuVDElWjBOnKVNN9/4+Czc6yb2EIAhr7WVAR
x/98qZpEfo2rlfkFA8trcrg800RJON3j8G4nyWr1F1FTGh8ACet91fR5Sawq
bQooDyNnCzkXTIVlckLeIsFiVtX+tEi68cIvD60ylL+jeNn2Sm4VmESR+THX
JdNOqu0agu/ztdO5D1jautCJbtoINU2kv0sd45Va/NVPeaPCihxLl1la+xxF
X3S0bntLBfLnR4ulD4OIOKdCjj/G14KpbXMrE6Uauogd/G2v1CdXLQM1zATB
LtcvIhVhhsMF/ovLV0yMgx5qc1685k3HSATlsr21U7dTOQBmugNdMuwpIpl5
6vIESjI4hwZ28zsEZa+hOWM/uhjVntcD5EOFt2NP45Xa5F14H3eNRpyzWmHB
DXkSekyDXsd10CDFEbemexqKnQhvvp0X/A9MKUI+tf1fJSDOxLUCHha1RQCM
6MvYAkkD1bzuObmv4bDWQb6kEwKE0oAQNSc5xcJyz1a3A5QYHdPfe+pDuqKt
w7fejeTAx/r/FxQs4AVLaFTBkqcj7bTu+42ISUstqJIx1w5vKeUtly2AU0pf
kRmt68vu7BcKL1u7+gtE4FVRLDYzZCSBP6HV9yuyI/ijgTKVGkNcYqIKOjuE
qhOhvWLZfdFXtJa5FDRf+qBKPbtIM6/VXim2GEgTWtk0/NjSaK8eWi0cefzx
IfDwHt/6I5N/Hx0OpPi2Ek7QMSSo4zUxlY4SEb1llridaj4GhOQekb1ubSaZ
b5K+YX7Giqe2J+c+AH0QMd1JXp8WwylY0qpOAVbhtBRZ9ARljW77eKOF9BRK
crTXNJmh0lEtGGvZvQxv0/4ZwhDgon2La6clIHuHmnHncGdmbISHV899ngpq
tRlvws9YrdqJhTj8bd1fUxpDOUkECMcbk6eWFl/Xz3Eu5fNTRzPPHhLVkyJj
ZgvW5QoiyQ+LSxlm3R+imalRYmXqPrqZHS11OyVAmeo7KaysYcakt8EMKXzh
iT4ZLXIDy+PEVAsLJfWGNiLbpFIR3VHC0gLL79zSCOHIH2a7cu8HsHBZi2nW
LJXlsy2zBjYvRuIHWUzkVdqYCuvUzGb0aumliZyoGYgjyU75u2bYOGmm7qsh
DebsRKvQ0nzfTkxN8ymjq6BYvpYYPIn6BddWWbJmNmJ7gnCKyVbPowrmSKX1
ctiEC0kch/7wOvVa8Fl+lN5elvh8AgaRF1mq3NilmQJj7U1EobQad5w27HsH
Cd6aS6GEosgzt07cDcX2MDdILpE+2T0fQ9SLRseGFWZccnugmXwDvb27zkdq
/D28SP/sdISFWpJfkRsfSumLKHYxokUE+ZxZm6Bf2SC7yA8s+nU/qS8k/wZN
CKEeE2KHbd8RmvkgcwOQ+XJkqody7YsJ79LBrmMvcxk1xqwoNv1LlwXnodzh
0DtDqdoNf4EqRdQiIMFNh8Nx2FMFhSaWrfXeu8lKhCxTAkSXxKCE5o2ItpqX
+rVsA3vJ0H26LcVBnA2LdEMvoxTQQI7AbGODa+2pNpQdlolbFDAjO2G5Pbqp
bjg4ruaFq6H7bxLNY/LbtDuSwFbZLfKfEd88gP5bbO5LW3yT+egOB13DyLkT
0Ac5OEDrE0kbynAfmLua0mCzGaOAPnblbTMxBIdJNo4grksgpP6oud8lrt5D
75H+9hk1J3TzAeSzbZRUkVLck/S6eC6bqEPRnuUgjYwoFE528yqxpZyvS8D6
tCfLSm/F00aSAqyKnuEx0oJxMt5Yg/NnMK0p7vjc4QfJBl3BGm9ncYc5+71E
H2DNnNliv0jpfMPnkt5iOQBANu44fRtf32ruujXaToV0gp6J/Erib9WCsZJo
IFX0C1YN3QwS6cLT6jKQActfKepGRi1WU8ZtNmdo4/Xhoz0P0+zVYGJ7Rtg/
fJzKishQRCdeM+KNgpjs/MekCnQS4mL7m/5TTYLWDW1p3C6H1Elz77BHxHFs
v8azu+Iskhbs7b9Vt/WFXNHKEjiuFEHJWybPBQmJ9yqiKXZV9cF3ALNkJ4KN
vnb9zNtSNWLMWmQ6Sgh24C49+v2p3HQdhEctwep7ltFz5hsM7Y6FSUq5lWBn
L87+G1KQ0FJ2lgnMl7fFl8aBp/USsaxVmvLItwLXBv47g4T4RQLDO591T58p
C1Lm6DpPWTAcdKy0bZN1qcQpN7hHZhhX6cZwE0ztkXqSsxV2KBTP5aANg1y3
03xKSuKzrBV6K0+P0DWVQPmrWXWq5LnRJy0rCT/sMkJNzK4wbm/yUL2fL/Kj
Xp+vad8j+y3qGUEC8fwnRrIeF8ODugZFHPYzlWEzhFRPyLOYdeE+CqAJ6f09
tyn5gEd2XFvnryUodbD2jc9r6HoV9//YDcOzmc7WQRDv1xqS7MIiqarkhOGy
u9OBaiG+7R+C6tRkc7DfxTxkTVuhTNO51/bKA2ymYMp0lJLee618/Og7XfWT
Fest4IBjGeWkphxtHDj6EzOBEVwi5PswfAEWXoo7Qsz26xqTggy1egKXfc71
E5s7Piz9ffaQpl1wELYkWpblM0j4g2eA+Evshs70T5lGCy7O9PGik/+Rmstr
Mj/5MIHt7E4I3f5iongHkIDTOC3SzmKPpClZIuQxiIPfyN6wrFsIzpadsBCZ
f+INyiCMYiPggMScOhQvK0VSa+i8b5shi3oKOfV8dxLyla0jKMVvZrAa2Z0K
XkZx7wlnL8FVRM4xSACLmq5nkX/byfCpcXARHRrkCaF+QQ6YjF+ifw02sJs8
7ZAk0S9GPPedkdEURYYPiKwWwJGAA6xH5fREEEuEOZs+stZDS8rB1pjTaHCM
9bDbYqDm7frC83Zkn6QgiHfqdO27W36Lv9Eb4xtuegwwuUV5n2Xg9y3ynL+c
cpNtHQaNXgvC5L6o+snteDp2ffYsQR1FmQ0YyN+gP5AJwVXD5CkXB72djYm9
R7A7s7+S1gEbKf1zFlRUtQLOK9KqDYuqGubaoQfg1UEpQ73ydbbbTTFxhsPw
9WV+s6A/qgeB2+flbqG0aevC6HOcPeerCakVD9uUROhm57Kopg9e9EO3EE8/
x/wb2GpY9npWCZG5AcE+D0V4e9Mz3q9xXU4c8+wN6lAWZAytO9k2MwiQFu1Y
wiHZHYmCaBWVm3YlOoqvSBC4ZWW8VH+bdfaEEB14BoL+AuvR/h/r25x1ITJT
JSeeIEU6wxlCuUIvlDDuBPOOZN3svhr3cOQftbdrDxA3fOqiQ3PhGgoGCoVw
H+xVtDo4H3yzGufvSQ/EstzNkeRkpcTb8+JOS/PDTAa2RA3LT9mrnqmxMy8y
h6cp20DbJd4s+dUVysD722GZXbDfocW0zDxsPZKqJ5hG8518iiOMLx55LwXT
XURJJlW+ldmews5r8i1dSXUu/k14Co54nrHWvUs4iVVfbFMDiADR9LhpphV8
w9VPmHqCc+9ENygPFiPTjuYz3V8yWF1K1Sc3bPjnP4BgZJU9bhngwoih3ieM
1o5+wJ+R/P/z4akvZe2itgTFuUH9KK1C7VXMpHsQNyLbnuWf22sAMDCBZdsI
qnULiTmF672Ico3QS+cnEjGkNJUGCaOsnQRbEKUGb8ar12/i+UreT2FkP0oF
nRpNoQaoDRhtoa0g6Cxjh9QaBVUQ+AT6cImF6ionmhub62ph/Lt/V9KKaoLn
/o40tZ+RH0XrKYywBFWy9Y/PeuozTSRbqS2s7iscTRGEBdUL4TOzBjv92U4T
dFIzLO7K2yqgv+EyB97ytIhN9F9uzhn7eJTezesJmLYS89dYCHATo5qkYaMB
L65KA5spfkiWopWhh5aM6A8H4DyxaW0ZyMFvdD5GJV0QzezfcUO52zMpoS9u
Eb8PLqYFH1ryUM2knBe6HfnTwNc2rdf9xVNNly71AXa1eIyp6X3sEKsjZtXS
HRHKu+jjfjdjpIlUfsVLhULYYo68woPgExCZS0QdAFZpUQcHFAzEjN3GgpOR
FcEtUNfTDGdkDdVXsM+f5F8rwSyE+2l5/i5uJujrQjfNLJ/EqDuZ+Yf2H3Vo
6uCUFGDSkGoL1yvKCHBcut1qvQgmJyeAIlXjLVDerWDD8l4wwI72z3VLy8gU
SbJclKINoOJW71Jwn1sc378IWj8Fnvf4O1XJ3h7yWidl0FTiU/PKeCyuEyJ7
Em8EC/2jYs3bu8kUj9zXTAmx63rgHjMcE7H2txfsed7mxiaf2c6rxCXLOfLl
pUm+H7ljwy0DWKJSiaFVk4vsILHR9Gnaao2t6kz0OpPRcTp+gdoMwQJkc+28
bn675OF9ozO3EtTjUxJrmnqruJIo81BMolgx4Tkf3FZr7yoxSgG5QfGKgZwD
CGaUKswnSFK/cNDofUkV9tY/Gn7D2ocZE3jSX3q/3KJVAyN1Cw3wAxvqDL54
CF2TebouvevCCS5GnMnonef2kM0VxkiVTdDM1Rfsgcvsr7YurFqT7aqRkTck
tETRMPk8a3yxjVUsa99S9qqzJaXlygM8ae2Xir6h/uPIrwKxYP+A+cOyXezX
kY1t7mDIs8/s8qhtqn/xm55uxGXmSuVB4taqbhx4lE/N2TTRUeJ2K5wR0vHL
+ECWRhLYQohVot8lL1M8KLdrRuqscoVyjwWZXa0TXLMt7W8n4Kwilqknz0Rw
mz9k7ptfhzY6Gu5yWDJHQ8UOSdjgUIA/wcoDGjb7QzuEut34/nSDPCxdF7hK
JLPcMjIk959wriO2T2JIRiGhCEt3mxZl2FTUKEerenbmtJ5naMbTREqT6o25
YHt1P+hUjNUp/KuJFVqcgqNz90xVhGcW6w9wYeCCYgdVoaa1CORdkn6kLtbA
/T6EX1yiKp9brzwGUIfISIWQ9Cu52uA8dkSXN0SlGagyxDVk4DzUWSed5f5x
8JqNeU8EIOSiLnRnIh+3c1rjvzaMVMSRGbHOrYAPUmR7SOpeIEtPNVYXJkar
lZndvzzUqIgw3v8o9X9+/jT6+vxfDHZqeaNX0qo9IgCzyKSUBp8aW+59UMNh
rYCo4JiTKuKmuFqDDHhbMwMilihx+RoTIxnCpAUu5shxoqjnL6Vwk2UjxqTF
SLIjiMrD9iIntT1nOgJdzKgUsEEkfSjOhRXsl4EDEz0kBJoXurS36KnzJGNZ
2RVBOb7a4FTbfPE3kKAZxxT41LQyQ/7HkALm0P47Y00uJF2i2kwrj6lBM/jF
L+IqBhH7JxVId3qI0PekV72VkakFfCgNqPuQSxq+DmqP6rcYC0s5zLS8UHJI
lMAq4sZsflZJ1TtoMfRz+IX7h7XyrkvE96cZNzkTnsLqozb6aL0j6oIVncLW
2TngU/7MUqpZAwgD/t/ksKEavgsQa6ibsy0iOX9EFWcMQhZNlDBuLgmHOMvA
39wE8rQOuMNzXpiGh9LgtKTKMk+GmnxSeWoMTVAub3PI1cVd6vwc7ZhHv/RJ
Il9Z55FS4Qds+sb4ykNqXBy/+HP6BuCdLKKziqAYhdvw4PseQpKuzi8UuyDW
SSvggCn2Lqymvo0ymssKcK/+4EhTqdk3/FzO1D6WvJeHB0IRa6Ui1r9IQI2b
To7HSm5P8j2MqPQobhDmr2tGOhB4GV4UzTWWpzykBW7bo4ic/2e5O3CahuZS
yF2NhAnPmKucB64I9IlHpUYQHd990wmbVbqfbXgD4n3foSLq3X3jMg7RQ2ll
+YP4x08qQaSC8G8cBckBpsCNHNkcbWDKjGF/D7n+IwbEoKL57D37q2/IsYBM
V9cErSOmGHny/5NIT8pztxdYoV9N4LMgiefJnEJCB45tTmv0S5AnG0/ybafn
a3BMt6Mp/tpRxQQPiC//Av96tFkR5OOFduJ/oMnoebxjlp4XUDX5pz3DPZf1
xRMzXKC97//7ucHjgby93AF4oJFnawsuffd2QO6UKF+ZGMXg+lYctIR1jyFT
MXk3IXFtX9tGlBN/vQQaeAFQoN8Of88B4dfSy9SmnTYvEq1shtWrNJaucr+T
0WS4B1vRAkaljfKngPL/6BjMWBsVWGzs80l9c5kaoX4vQcCdOLu8ynFC6GQ9
N4Lada5s2skCOXU47kvuH4Lmq4kn0SU6AcUvUJ+wq4PyV+qUJ5/0dvAAbd5S
m3WpFKGH2pHKqVVmWa5DTHhIj2ds4v3LpDFlX3GJMjy/TMmbEO5ZbN6lG3B+
0RnFQAOtMznz89dbtZ0rtGCQh+o84naMlFf09LI3o+6Xekb4rm43AaarhHEx
uXD4FK5rNyzvY14cuKgYY4S7Tc+dtBJ+WV8l+jc6IdJv2Zt7i5+gGLMzyhEH
PNKYNOsw5wMt1i11JsDRa3ROrRBsp3LLNRUCaRfPwwtYPvyIA4Pfv4FllJXa
7VKHUsC6avCrER1NVIa7un0BNax83onCCcsTJRfbbp/IQcm52rOrqolwHRFa
G6E6YLhs+Ts6sNj8ZJjzIbAi7HD9LNxlARQa4K0ebisxwon5DAn79ATqY1vS
fj/MVlJNascpE/OkZ2zbDeNySgn7Z13bTuPEvzrgjFRNpVNlHzqtGXAmE29/
5fKZ7YFzBh8LpKB83+zulK8YarjTOrQD6om0TBEcizRGjLxXTF7lDecgC4gz
nNVoSUiv5M1fYaXJlYhs6UkJP67DZczEPymzQV3+DtQAZH/1Lx1fiZwx5GAU
yN3NLw75E7vLvCcoxKsXVHQRSZHwIYOyTqiKxifhRoqwwwYUZc6Z/u153Fn7
zDWnzCrguw1fEf1SA55NxWB9FMhtsHDsIOdVfDP4gFkW5jes4xoIkaPYKY/k
7blVwJnp5sZ4raCeEjzeEK4wsVJWClVjqWq95qpvQzYoPBUsAMQoUG2YMLYR
l2Ebi7hsAVViXC2JMh/lmFWGD5HvGliY5HY7dgjwkdKNzRUjYoiCZtFwRAz2
hM+SQa9WlhLN58cDksrc0NdYcuwHPCpq5j9M6vDtQUwyy1cyFHmiC+Zm2UF0
cMv3IvSE9OwQOjffQqV2eL/dXaja177WFOue6dLgFolckQMprFSEQugAEzLD
WpmSDYaSHZ0o6VfWULfLUy/f8RrX6enahMGk+OAD932jsOEtLRFLWqYEGusX
KijaPsFjTdRFIGJZO7lPC1K/jFk9QwUsomxpDd6ALEB62vgqkSTxKLPkceGW
d+ivgF13R7HdvNggJWUOzWiQ1SVBmyD7oxxXzS3mYUxrSOC4/SE8uY5d44FN
KrkIV89NPLcPBn8LtDafSee7rDD+LDaek6edpbdxnJTla+BxEKzPYiGRPs55
vXFBk0GvMtCZV/Aa0BV+7dvTqQmUG93QhBRApQyC/xwnEouEh/5tCEJcZ6Zq
J8FCaSxXxQVkNsaMG6qe/lX047yMLZENARh6MN+YtloXiR+tm1mqGX6x0kXl
C/m+E1WZ0lCNISBCgWPCYcrtuj1VDNJ164lbWuAoo9hX2FC27tPD3Jrt/O+r
DdaT0uSlJEZzZStoI/Eq92d/g+6TtjML5EXyhE5Hpk2N8EUuqwMELPvcbj/z
vDoBDkrhtG+Qe1SP/U9MFuo093Ay/k60LD6bQNmVhI7QnoVUzJetWixgpwth
QSjgnML7hPIaZ7RMqMQdpxPiYfHi007j7vBZfbJC8nrixvSLQlqEBXdWZuvJ
EouJJAauhu9xqrMwYEtXQUmNxCVddf3sTjcJNBPE5beJfU6dzhypN70tq3cR
/bO770qjqUxL/sWWiADG7Cu3QSol4dYqmYhTEodYc7sSps6o76AYcUNNcWEV
L5OMrxFUQOZdCsYnEybDg1aUIEd/EhitI/lOrNggXo0HXtPxD8vM8+0QrV+i
MrVir2Ipelrb8B+J9EbMfFRS7Xfo8Qf4mQmX+WehV2W2i6blsmXyJk5uFqw9
tyF/vaH2NldkccgcOGMaVeyyR1Vh1YtrPRY/sXNt3Cir7uJZdT5PkuYox1Gw
wWI4vXFhd7JoJeJrxlBoB/zVWDZhIgvLsXlRUx65drt2OcQZzl/oWcp617vp
WbYBJ8wilUs+X218Jx5HuX8HS+pPYB2CXJtLLG9zxstPzouneT96AmyIeuyS
wNq62f7r5j+wTGlR65ajiWWXjv81R2y20FOqlmRfpzRBZQbSjedkM26TptaZ
PdOAWbjeTW8/XEOxgTMzJIwaq3OhWAyb0d5+EWkbKhBkyQ03lShCprme9Rc3
xonfTnAAcNc+dkNRFoGDzEXrkYSoWXjUGuP2jP3xrDd9WEGc0Op8lfBedbaU
LV59nYSWLUn7l8tduoVWYgGhVQFTOUojcLKANXPzSPN6C3CZAi/FAGY3y8Gm
l3R3DGIEUfj21f+phIOOu0rTW30uvUbr+Kho5IRCCW5HcfrB7Pdz9LS0EpIM
qXecvXILzbFcnXwdwgfuaXgPko1ggSJeU8Ux0HYqpgG4EKqQR+mJGdIONkD1
8T5yFB3OHIbrYN67qZuyTfV4f3cRXBtYYGFl/SHntZ6MuLOCpB2QFj3wDLWB
fXslX5YlRjmZdbV1DMsWBFp0gCv8Gjq4lG/QDA97SDEAyV+wo2LO6VU/eaqw
21fLKjHlU7v39PYCI49aCZmZCjlzQ4Ro7TATwrhDkjBocjzZ4v3632eGar4I
b+gKBG/bZw7LCV1ue1KSzDmsq4fUq0a+P9DuBH2exGh7CeBxQ0oJ6SNFQlAT
/ojaAWNbHhAvQvcxc1TVJJztfXqj35hYgFVvViNEDJj8kv8O90XoVs99a96Y
NzpAWGfRT1gjTFnTMvR3LYpb3nDKDwL/lDchZ0/dt9w2xzsEBSMOE0pptWBy
VbX3KH+XpjLxFrDsxBrbvB01+Jzr9grBKpDr987pWe/4fFSS5ZJe+B6mMbYe
Damhr7DEI43dyfDWw+7MI6SuD+C6YFe+LRLGxU62jpcsHYM8ZwrVZjH8BFjz
BYi4oXFxEefWT8z6j4VpbLhYJ6FpkSADtYA8N7uwzT5KNEEGKOjmoFj8cf2K
xxayjnQSkMNduZjUtAxvo1kDdpG8iA4uQq4jPv16oTA44qhCdm85MBUHakSq
KfATHpx4u+O7uB7slxdeZilpW4gr34oAToICxLHmFl6qXNh9vK1UhdRzf9yT
iWYRscfZdl4yyCHpXS82NIWPFlPbdoIHzu0OMTVA5USqPvTCBQrFd+1vgjCt
DthhDSEMeDaY13e6BnfAJmHkP5MB6Vbw3KNDo/GTgMIFHn0yhtsXDFMHBEdZ
qM4hlCEJfyE7gC0iSFZrO4B20qtzvgZIQ7/0x1RYY64sXtmCytfUseQ74vfP
Y4wFDepCylaP4ilaAkzK+OyDWgqRDPfk523rWFX+wkVC4iIHreUWTJwQ32Bl
G3koa4w39ZcjUFgBnhlLKDjAXeqxC9oBXPL4z7MUPhD2qvV78WAsZ1aDsqqJ
GbKgewgcQh1CORmbFsHGm4c9/0DyB/TzbJcN1UG207I5F7r32fX0QNvfg3mR
rhE8CZw6Z0rdFNbUocMlAsEphBKGJ0IxVfGyPKSTzHWZ68NI/2xfW0FthGKP
4P3lHYvvCQgdxIsBY4I1Gancw/tlWHBfkHNNqLFLUkYW9nHri99csvMWjxfq
UQwPjqnUBGd9nIAsMNNxoakrLbt8SaShJCbaGN125FiFXObBgnkcH8irNwzG
2vufzlNuRSl86JlLiLH3dHFmbKj0fYupPQH+GSH6j/MZGpcqy7Wet9reXdaE
ejeScM8tg6SY0nVOHe+XyJgvRUR/pMss3bC9fOn82WvZgZTDT8SidXYROlt9
zq8xlq429j+izd+1fB+f9mr1dVH9iCRvL6QQLZbPprbfvK066opTdzKsvlMb
AqMjY/IwQQvZZsRwVFiSjusPDW1OZWeTxnvfSyByLA6iJK+WGnC6HyPLQuF0
VliBkTot/uGDH7t2K06EXOaxlFMHXh2Dn8oIeR+mBXYfFneXYUi3HqndoZzs
LcocXNgKSriiJ9xad2qQHy8im9FDYwYSwpLHPlqf1fkf87EChNNh23cNVnLb
CHRV5wexZgbJ2UacPzKyYSV0+thJcgcTc9YgiOqHzQTBsgsmcv5mEMrVut8/
uVf65dOeItIcgA2v+cxWLYYZvCj89sTl7CSxLpJ8FhMgO6rGjeV+gQSy1WCp
1jqssHfF+TUDavpeQ5PInYed5rWwHPTfRH00UApNWsKlsCAssKM9cuEz+YVv
U69ewI5/Su9ygNh0rS7602SpSQnIxy3Mus4SNtfQbBDGjaJ/E9P6nDyC8r2W
Fcbe2CN5bpy+bluGkb7XtQiRGTl+vM9d2kkVDPaYH+ANdeaFdE+1H6Y8frVj
gazrSdQAZFypAJh9s+KBwG29ieyCvaySDRWT5fUY97F6wsCv5Q1oAZ0hrky3
FVnX3Wxq8CW0D74siDqvTv9TH5lFGo3Fc97qZr9jWj2G9mQf7rkiZbltL3wh
581rV0IHy6L33dYPnRamBzxtG/iCVq8nm67tC0A4vEkX/5XdtLV79lKZ+ubj
N4Apsj4bCyMVTGaMhrM4tk8xUyOYcU4p0CQFkAJCJdkw1dR+r7priszZl+0M
xfQaIHtj+4UfkXtRzUAhE9UM20knGmf6063ELCU8fjIOa1aZu9Si1QYZDC1C
KcJOdPaUu/9yQGLrXBWGtukJFDhBrCmUz3berXunhk3N8jZ9Y+rL8nD2ehkD
2j2qDzU4MupIWCEbv4eG0/Xg1BqELuWdrqqBD4J8fhvcgjWoaK0Vj06A7O4O
ZNUs2gaPDBquHOX4FV41us69k4LK+pKpKrWR8fxB0JYvtjLjtAszNtOey9Op
3U1m+1bBO+RsrwqPpSktgvRGC4Sc7u7AmkgjULKiB384xry4rMZp3cAup6oz
Z3Mt5gHVWhrO7vsNUszj3Cyjti30+Fdb5v4qc1duc4DRjSjG3+IzobndE+Xo
A8HO10MUTU0Lv8kOY69g0r/g0Hdf6dZ2SEM6bQcObm73McdKNVIE+x0gIrTG
BNmvDhBjqwN3308vOvZdiM7plhSR6dhFTREdtYnhZwGHuymGnOGmpvQejoPf
nQY3lXcLKQYSPwtqB61W9zT7Gt5pN3I2esW/au0hJEM5aEknQoO1Ea0Q7+iT
X62hLsD1xlitJuEkHMBrqvWXU/XZSWml7PteLL2H9G4TuN6EC9qWFhVqRNyo
zFCzoBwbOAZUZ6kVc2CLm0mItoplZ3XATCBeaEBmf8CJETbOeLauUu+5sI3j
BInQSHLAnA6oyhqumwCmA1GVoI7scXENjZvUsv90rLVQJ78YdlMS3NDcR/Rm
va01sl5qpWx9DG/MNJFYbWkJesLQY1ti+nCKXG86jbp6oMhGBoQgqpVXdjgF
MQXJaB5gE5k0E8PEOQ38AoJX+CM0lcWWX7lPkiWIXteTUiAq18iUOzY/Me1H
V2UED0lEjKbQUVqKSVsvZx6d656cZkcO4JfN2IpQcI9EoGfvgXUMdlHBJV69
uqPDdXVJwoDexccGVqgAsk3NUB24M6X85XiYJjo52wUxpBTae2O9PlujhkuS
SDb5jTyqcJJFuYYhEYrlHTVkKOl4nJ4yXWJAk3DinfGJF8fq0+mj/2DW488M
DtG5Sn779X3jI9mAiF/dg+6Zie7W/IGa1oxNKIoVFOhuZCm4B3PsWFPtWgjS
fhHufy/EIkHvE7pOIMkaEDPM8PXdq33RzBiMdvyZHWCdb/NqpAgBIK2GXQ7O
fwlrw05d/hbmNj28h1rgNXsw7sI+rwwUMJ3tA4HoQbCUqNQUKGuGrx2AQRSf
96nqI3JeYPEJgkxGA5dpeQUMUxOdQwxD8H/m061h4pcpaBGcuLGrh6xHPv8y
9kGismtIG/yt7PfZLrdS6T3bzX1TB99TrccFAnmVQXcJf3dAd2dekWzIvwGY
eeYco1th958+vCW6YHe05ISxJvlPzV2To0MOTFmSPafC5OmU0NEOQJM+oZgP
MuCimFc1TP34aG7SKt0Ywvs+jgW4J2jchzJMsX3wGp0NIBPY/Oo2s/JWohXF
qoEh51tuNPGq+s35Lnjo/B8hwnTI3voW9rSu4D1dL+SjbBMvFA2lrIFPOdWB
W/K8X3c2P6e6IpmVbXt89eLa2ngsTUmtAE6bxy0NA0FMlnuHXkRe/aWT8HqR
NnpxeaJGj6TchJve3z8aQnMsWzynkjhT1a1VTvP32JIApBj2e5Id8iZ+kwSv
YjS2X02zgRWIHYDBgYt5Jjd6NZxUePs5dRhAJv/jUY/JjqW9H/8Eki0bXDTR
iLZ6rQUH9JgDdw6rkxKrS0JtxI9BMnhts19/xXOgFIyIrSYqwosivCfmjpLP
8J36QaXYx+g7iRN6JoW8awFEENjLG8pFoakce6+C9xegfhyPkihWulIYZRik
ULoCmCkkVL9qwpNGDjd1USE4PhKGAX51HG+smuretCX3cRP6SbrOkQW2JJg/
1aRwNGej7gbq3ZsG4R7ThDh8aHfgjWNssZ31CbVh18b1yIKiHNvbXE0lklrI
mcsoX5vxMD1u8JT7KCqFDQS/LQ4OftW6Po84vBVX6+4hqJdhdTth1arTXi1L
LMyRUcw5xDqIgJUgKM+NQKyzso0o9W8RiwqGn48goQSaERRIFBlkfe5ywz3n
y92CLtW5Vw1dyGOPY4hxZ0GRiNzQjpHH29RR9QFJuXF9r5MXDmwRIcL4olyM
0U95OAnBSjTQzyyiQJGlI5/BDtoooyQvrr35s3u9yBOl6uNM8ggo/ieQaW9I
jHv5rVZ47HsfBA+Nx84WhUmnKdxL96VX4Wo/CfJADzocvwDqYhJ1iSomfrJs
+Xp7hI4ob5wnLQTrDilX30ekPnN721+H2eaSa4YbLTp7gHcrCt4/m1aZOK4o
g076w2s6NkvyGMLcnbsYJ0N/juGf9B6OU2GbvOygBrUQ8l++4QVg7zDW8U/I
7LYjDwHbrhmrqE6SYIAJXOA70ac+rCiHQlYMS3jyTmOUeIJ/JClh/ok5XVxZ
gCx4SqfSGFtx/osi5gcrhgKa+jYOCXcgqBZo/jvoaBaDKNABK6UsIDopE9C2
LR3MSMlxUdG3gi1g4Kt9PyKdL0bpK59+mOhWsGMz44fdFsCIoKDeUzWsKa7O
exF8eSRWG1YONHBfK0jSbpO68olRFPz6uJdcliBhhuGzG0UoLzXdmMNVXPEy
SwlrmZlCwzKuZ5RyETsOn0BfsmR2669q/3A44oo1imvmwIlYNran9JNl/IW8
vck0OOXo0sZqWOmsViZm+w6xdEKbtDhh0ySBnQzB70tW15NHgbrHkmHQMqdH
7mBdLd9EdoiH8EaB7dVAW7cafy/9+ZA5y1rpFLf+WkhlLJAH32GKCOU/79gF
ZK9qMxqbSjCXWlVL3IHzniEkb++Esj1q9wdMdsaWd35X6McJQnn1JpkL52R/
bqzkEpJ+2RWdZXaXRSy+8hi6qYrzkjP7hTz5qyzU9FIYnCG4SbHSav6V8xk/
VW5mUnkZRmGei850hzDlK/1/INmWJe9w7btnBWi09qAGb6JQFlK+oVXJ0dTs
5Zw+v/W8dCVlUdm4SZ39gEy07ypMvMa/nlQWW5rHt579ju4nvgBdz40OjHhT
zeOueTSRnHJsd6KUD/xxDf4oC6fODrlBHCOzX1ZKd2ttMCi+7FrJ4feWvhkf
9CCMoCtkCxpILgspaBYnePtX1NzhJu6VYv+nucajBMEaEqQziYH+lIvU/jzp
125X8I8csmX7++0M6yeZisjzbdLNtLOGkl45a0UINCkpWT6vOhdbX3eYUGa4
L02NTWFu2XeyTcgbzf2U82zCy30SL6bN1r3OLX0atxrhRc8QxS+QKQ5yler3
Ohg/DYv4zJnskGdRsmZ1YRUkDND81mjUTL/H/Rq6gEvEbuzQQbFCgcfSKoS0
9jJIRch0fcSZbLthdXCUJ4VHLkVz1hV7gP9h0Hy8aHauOwhGv7TH12FWA5vt
0XyU1kikhrwJeIo4mw2ut/pzB+7DkGEb4mqfqLIkd2IHdlmdj9bDoME9tRpf
iLIccTYWy8Yw+EypJOugvu9+15YT8dyF3XwgmYW6xpO+or0Pics39CZtYU5b
0ReEZeaFF1IK1yEDm0IOPNxrGqJJLsyCFdFfPJ0RMUuvAoTY/j0AL9AhreNL
jl9XTRmyDxcyLiC4nd9GPpzagWZ89AlR8qFTTd5+MlTxo3hrdqeHbUQrzUZx
y6w4GSD3PSo262/I3pft1HEkDkGEtg+Ofms+F/ErVHKOF5CRNkzrWaNtFzEW
faRqA7z+tvWpx0Kgmnm1om+x07YQOHbnUDL4GUwSBjdRaKssDlq4zfcANGIl
wK8kEx3JP/xU9oVioLJMrNOjz+xFCC4Yoqzo2EFVMVUDPr8nHW37jPau/VU7
iC+shv6Ouce7H9fbAe5A79IrL2tj3wfZYy0vSBTn/AmlFi/G+tivaQL9AFfX
WbVSadCjrGenBXoD1bp566y1yxFR/Ty7TDiK26hnECvDgSjPSl1rtLiszsdS
2G1UzVWl/H+6nUNOixny8y5B/KlEQL/GAOVWI7vi+yGJaDjhiwOy1uF86fDR
AZ+PHYm1QIvGr9/l3Q2svA5XaoWCLU15OGBtNSp7cXyqZDby6TBT9VwAHyqE
AUv7xTpCls3zfHCx6vK4mX7I3GnJV4bO+qcO17HFK5QJHBntCtxjjhq87cv/
e3kpRVILHXqWrhMcz6DmAvMLs41bt8TPyRosRTVnWn0z6MUM/spw9NuEFZsS
74YSWAqCMuTVMf2P2XZSsQqj3oTqRxACrU8o1RMzWUTmL/28Yfqobcqtxpcg
sEkTho2bGVIooVVOghYVPu1BkT2Dz30dg6py/bCpv7SDNuGM4mosctjsxRcc
Rg3U0IT/UPppQTZKiDXeQX0uEaIYFVPEFunslbtHljewzRNMSISxoAn9cvhR
AbDnNuEykYqgC/6GE1CmdE5ipUsRPhFqn/dghTq5WhqkhRA+6P47fZOoIqWo
SIztR+aATW0DtkjeSH1W9Ncb/sfotl6gLxdTRDXGbfvWAGW7dYF4Sg70pNsA
2tt5Tf9K34fFhKxd6tBju5WoyO7W1IIiAbo1QwzQMP6D5B/kVZ53lannq3ZI
+HkBDnRU8uUSd7ir/Zo1EFAHo5ivVMjay4riwWz5PR4Jh0RwzIs7Oa6/UYCV
DU+aBs9ryiPKdkn/LVAXo9yuzZUUuiMAGtzNnoLzW+sKRsSrSpPZT79W/PZT
/mNqHkzeiD8AW8QPKNK3iB3eNK7pdbcMmBSrR63xD3pcQyLtoIcq0ndPHsWi
0T52J3RpFj4B7HG8vvMshjm0rYNtiYvTEMPBQRUhIrVt1BT8QHAVbGS4QnX0
Ih0BjhgH/MAoMv48bW+mI9zWANdwdB4BzmS8im1rjoxCT4lb0KIQ0JTKJBlT
+EG9MMxNrouoiAL1BoPCO8KLrQhF15X2zDLxRUl55hzE+ZJJYa1QnM8TeUr+
Ze+r2iKoC3/JLj/HxU5+v4LY1lODW1DbC1rlbY/D0Qi1OABTmJwmDJMGCHfJ
tbwIstmSvFnR0Wsk2FMQo7cbD15CZNaKOjLeyRcjLV6LXezxbiG/1cBkR6qK
8of4VfMqMg0XXjFaOCHr092db4YECqgaGlMoYMaHTTt0SBJqd0gjJc0IdTVl
FPg6MFLI79Awj4wBOO7Kjgo9Qz2rFGFjKSWhL9lWkPS34opMdJPF9gGGCtNv
aYd0CqOn0+N2k3782n7EJmLA1495/9vsgztC8bb8dZLbz/hz2QVsvQIAwySV
pcSiv1FbeZs0NW2ukiPu3eSBdVGd+CRE0mf8ux+q7Fre7huXgC2dCFdv98Rz
X6i1NpgI8VhcuuZZ1sPVEOeZafe1IFV6prf+IZbO+y/q7+pVPz2MbRcKe2TK
jRyMF3O8qtYPcyGdU57TLTBUIozKyYZoq2z1NBM/0Zs60gX3ZB08ZI73M+Gm
v77SDz/2aTi5bTJbTv4n9JRSdi9aohGp4k2t7u6axtEpCO1uNyvKwnU2ISki
P4XWAt/xpesBoyRWPgG0LTsO0hkRWsNML+znCrs1qSNBwAaX313v22BrBohd
P/OIr7EGCTQDB24SbN7QFdRkrWa5tPl6Z/mOfv8C6xVFYiPbY13gA6lDB2KP
a9qwnXE5FvLbzlO6qaBvBI3c1F3hJXt54zuKfZXXzi1chiioOn7gXREa7ztj
ZwS4f8eCRassZx3049tLH8gsLvkVCdwLAhfJxRDdDsPcAH7G0oG2sFZwb/j4
EKLSmlQq4QRrM9XoAgPuriEnnRO7kfNiI8qeG0LsVbIAkHnwgu+aA16ZUoTF
ggH8B+ShHLTnw5CUusFAyVLNFrXvot3XdhoSSc9ihSXSE+ZjtBkaEE4Tmd7F
nWib423P5+fwYmfXvIWZ/gfuDsHnxirPHfU7m087P9C9AmyWT/tPoZDZL+dL
WwjVMYQdKmSvqoO6OQw0U2daAPIt77aLbKSUPuWie4372YUf4Vbl6t2o5YEC
2hKy+32M8HyCMQ19Xg==

`pragma protect end_protected
