`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
LefbzRBIbaQ7eyc/fVs9o2yOkfmbzCtdK6ls667WUWai2H9db88LGLDrd1C6glRq
w5w+Crqk1P1ggW9TN2lgpjLZiifIP+rKa4uHBundI3Lkb6ITdb7An8NaxLxLj0K/
GA5CMk9ZUXzYqYo64/yNsIXPfOyR11SgEsukufNBLvA=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 3552), data_block
jnMlG9lRLmrE8E5z6O7d4NYuQAAwXQRwljBoZUogspHvhVya54l6FK8U1UR8Y4uT
75JOCGDX++028G9pPFPyiDz3Les9VXewo2ZZqJgQFCQ+Tj56QnaFiYII7x2HA8rB
CGkFDs2J21SMGTev0M+IfCFMPmQQoeIlyIOSQ0u4fLJ13pSGsxJQQUzBB/s1BEuK
lAW8Xh4OIGcc9NTrvVB05Q+m+BPNOan544rOCa3lA7pM6pRsd0raAvZ8jiV4r/Es
Ix3wG1JLAosZgX/H1Ke5UKvgTQZUZiJkuHeWVanaI6n/XpO/dcBMSSMjFwCKioFl
l1vNs/908EzNMxeI5C4Z8ee6B+rdCpcb0NTEyMeAV3DI9y55oWz2slf2yfDwOHPS
AoVQ6NAglxoo4uzm79IkUQqOZiWUO/NDRB0c/oh5xlfhzpZuPK98Y9FprNifzFk2
s6mNFsuWhFb2m+AqqVLWd1GtA9YpjhgDB2LuqjzPgaIWsyZZTHKLERIAR8UHdDvP
g8qr3hHSsLa+8Z7VXJmNUOV9FtoaINx9LtG+6+OuS1BKA5t9FNjqfPgLBveZ+RyI
T+/xrUpY7XCoxXUTNIw0vOySV06hj8VYc4mIEl36O/yl/9aZ3THHw6wzeu+yBd5w
blh3ZfAGOAov/C7QfzCOLXRRBM8wlNFyftrCI32XhI4Cxq4jJrz8r+LwfEtAy1Ut
bSOHeIuv9h/UffEELsmiglkzNdnqyqxtma/dzinfR8wu5ZiiWojUxL5rpOnwt53o
W28xNSRK+8Y5BFkdkQMklZr8iNInrL9Tc7ZxnFyrCSa5VhxkjzLpi6CdRPiiN/Oj
FzK/RrT8+CdBEiImf4A+2BkNUiP8sHqcG3R37ZmcYupLSRId6npGYfP0D63eANs+
VaYc/NheGBh4TNyQSLVOPX0LwDi0usMFQkH7GBZGJGMFfqURnx+XKeImylcQVvFj
+C577i0nl5D8BHNJxZVEHx62rGCxD2rvNO7PiXeELYR95lKJEadg1ruLEGXxTnoN
MW1HFlvon9yStROGWUCDXgp1NjBssjg1VUSrvyv91VOMOEfPAGXa58nMEhU5PbB5
KDkmCTrildFRmILuqt3k50V8o7piAhqqCIOn0uGEnCM/PVf5ZwlM1byxSkSRHd3H
4J2nidXk4nRXXEBFUf9yf2P7ShWc0drO4ffjyZ7WbFArG1hQH7LojZyr9WCK/Nj1
KnbRoDpjx7U9HS9Zk+ALMq7TRO0oSJJKAX2vQj2qkMkng07GYN2UUPMyCs2r6YBW
UV40SSmxRaQQ0TxafqgmXrH2ulG72Af+WfOPZd5dtRadYbzLQLyVhBDKdjaGsWG/
eI1wwoPPTrw9r/CSB68zhnfVb2u5MhaxD+Wvl/64+tsSonCTyoT/IltwmANHQvkN
3K4xrO+oWRYe63TktR4+OFuWO4vZuCBO2uZDORPezn6oWJ3jkebMVS7WmaOOAxRK
WQ2ckYyVchlhUUf8Ny4vE5IMaNR0WDOmpx4ZjzqO2Sa8mo+6LFGtVS9uYVUBsqUx
Y50LQAyv1MmK7rPt7wRDRlx4IwzAt8JDPgF9//aqDGZKqW3KLrFEQ2Xf7OXVuVxI
30RL3JhDNTXgAS54bAetr0/lu58MP6LGD1S/bhhFZ5J6PnBJmDAKOIptj8+rUrGi
4rJmtArW05GKduhzvW5CtSuwYQ3vK/GK4E4cv/bcQZFTC+k5s8z467gN61U5D/r0
mDbomMe/Q3Nmfj8Q2SHUfi2tU3rqe3eBCFajlAahXYgpKtOMQfGwNvsApicimOu9
s5f+8wSRPJDrpFOefCuKTmI6/OuEtj4C0FzNTokK+Z9oR3IH/gPqIwZCmT8AP5Ir
UYw5slc7kiNgenBLmwkP+75rhTMHMRQ3MhNgyb+UN9nzD8HENHKwNYye5LGcduAr
qbSU4c15da42LCnEYq4wEETLMmO7NBQHx8m+nZOMtgH+JabdZCvrpMa6wRJtpJaE
vgXYjb3pF7RnEpy9MyHXe6u81oVB/cXElEEsRjtguCaefM1nsbdsfjsmYqoBfjLy
mGT+diLz1sX6j4EtgwRjdFA+RiT+ieSfQFi9iqPAcl6g6TBjWkxQdRwefzEN195n
JR/yGyaSzfIkcEN2zBKY9+k96C4oTxD+fPS14df5OuJrZQ4iJPpPbWn3FaiuPrmr
71g+igI/if+iNRMFNYH8HKz3pg0r9I0jRU7FyXXWgDvsM2y1YPzdHyPQOn18lmC+
65CfguM8B3GRt/XLX84Ikt6CZAxs8h2WN1OnEW9Gyddy53yOqARpOT1rUZTK4Mnu
jnAzGdW+1jOJI/aRJQs3/bKSHz/zzXG3vbtH8djSJXpTB6KlCvI2gPn8jylEanCv
kAEVaADLiDKLJPl36M5VlMcFNDZvKvi69nmBliAbgjLZ5BeNCOWUvLvg/wh1oUkz
HywQO/xt+pvQPuFgjwwaCLXBBrYYnn/F+Er6WII/ZgocC7pfCozzVVLKoGfg2Ifg
+zys9NwB8wqt86Qenr4nQgCP9uR2P8R+Ahuciocsdl35zAqUJOsMPmst2V4uszhK
6M+BG5gucK5pTaNYwDOq0how1MAY/k8qpqDNdZjSzVm5ApPdZPQ2cRigxwJdpGLG
NV/ZU1GSv0tYH5mM4p640XsGWRoMXWtbZSfv4fXEDr0dAPCjuiO2b4wQRPKGZHW6
cAhihv2AwWy9WqVL80iXxdJilalrkHt46GLmQFoN6Afhe6qJP2kn0cNJThqKFGWB
PUXBSP94gxZv9h0sJRZPOPtecEZ0++cQXLaVavlU9iW8QSYCevJcDD81w1O0v/bn
y0f08nOrg809RDiB+hP4jGl85YpSsXkL3y/LjmCoQ/O7QVwqwllAKAcfmtSs8HcG
GfwE6FZb3fuFwmCcNlYDUb6MWm4EreC2VrysiOr8EOVbl0KDZ56bzDKbV16wUITT
C+ADGwBkf8lYjjs9Z+nnYJtJqG6kosXKqlkTWf7NKKgfF4ldWMZcO3ydl4Nyl2up
AOE1948OMRDTQ0iWAqy5P85IITxgMY2qqHFPi/QaFpCT/YXM51mhgvahlmYCb7Z1
XySmoIKQgi7sd1XFQwY6v3qAnv8zQj5voMLMtMVZcn1tDJncQFPbNUDtJyoudqxj
jk032GGrmipIEaJ+QBUKEckkKpYJ85ltOzchrl5BwG0D85ZaO53iX+WzuWNHH7h4
NtngLNkL6CJUpPhPtRKIVroUNNxeh9k/tIkpxl+qYWVwx1JhEv3+45nzmksC58P4
ZKKIlv+RQdamYxYhaVkhw2/ZqEXMuurtbv3k+RAuNgWTOjqOoHxBzIjBbZpoMwNN
qUkKQlgru/H/xYIeyXlQIOOsx2PbFTeinMSqqb26F7BqnUwLUOfKj96MYK6M8EUU
u3xbLLra3IWBh/Vp4ibaH9yehb4haAEo96f1B8w/UccrbFSjTv4dGj7LZvEIbCp3
ZvhMK2A4mrJsu+PMHGNLE0i5ahJ9sADQSgt3qV7YFGZkZrDNsf3vbOzqpNvPwOVx
bPJk3EevDP6ds0NtcTTQSqmmRrEHS28fXwJO20G2jNnmCD6/6wdmCalnSj5Q2+5l
otcpKbxX9V4G+zoPXw6C6gclTSvUvyDP3WMrclY4sgkhsBx1HtWO2Ic3iXH7ZaOe
ub4OgvKsLKrYSYl53xaYfI0Oj9eO8Uhd+AlRlkZsaukqqA5Lp64VxRarFkBFPJCr
pc4du+JbQDbzVI2p93qgp2XNmH2P5r7Bi9QK6ozLPoy5LxoI3vmLkck46W+iD5oQ
Z+KH3K6nU20r/adqF2W3CYNdGGWHVLdyx7v0H0hFP/J6rHZYULZRBcuYuzROkFvI
Zi3CKbw7NDwER+7EV36G3R+ATbzRD2kQv8wpHmJK7xq5w5UmtIrQ+Fs1WC/OWA+Y
Bb9CSj38WxMvWcWjVv2NnY5ccmBx9C/8e+V7zrMWm+XMskisKi5nngvE3L/wvGCj
aW5mbGQ+nJpqdNxG76rkjoNzgkhHkCK0zG65+8vLFgDTOfNVqTefeynSeFWdoI6N
7bpzYbuTZPuxL0V8g0eC3BWdlV3zvCS8k1PNvsh90KQNQnldky8+GA3oVIbnLdBk
L7NSLPMC/2E3pr98uV3Iu+CzthjLVnA7H/tSCxC36H7evHMHXfQ0H1mUB6m0YaoJ
qfbROmKvdPjbnQ5NrRtCd+XNN0bCZHwjSaGh0xM9i4OY/RFuy4HcNZcsD4oeFH3G
BYhZGYKFIACe+rEWEzw0vIMPtUVU0xVGRrbxRwSMLijAgbNzGLXSKPXxZkt8dnbx
I+69CBvqfulRwLdBQPaWFxX5uH/S6pasYOFBWkKRbGr2G5OrB5I9bXlf3brLWysy
V2QuOHCr9ThpN4vmlaPfv/E3smwr8P2NZyYBl/cWs7N+rvVm2O5cM9JjcnqVhBZ+
tXJfUTBsYW2TeoM8T9T8vVJ/InBcAriJrJ4iKejjpz2w1sD/SwGyteLHtIbkFja8
SXohkpPGecon0HLEtYrcxfdgxo1+pb1OcyQ2IArNF18ljU0zAOdwOIL5NYsVYTIs
s0t1LvjT3rbkm+ZePnCwGL3TPWiXDiXcH3HtNcNQo/mOg9sxjOx5p6PLA/h6aC1D
H/YwQ/JgYL0nzGbWqqLbIr9bI+a+ZkJjtrSfYMRzkxOXAs5yVdLV8VXAi0G7J8CK
EdG3h5+qkyJiE/BAL68TvGqT8q1zb9l0fpNbFN9z3kdWZT6eNsS1dml+GDTRFaRF
`pragma protect end_protected
