// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
mo7tvrVlu+MKqriZPzXk4FzLYXD/JowqA3lHEgOQ0XH30rEHWwzTjz0z9rvMpMO0
KCBT3FEuwO5aT9dR/b1wQkKjPT07NM7ecIqQ7biUiZgTPALoIE0ZbowL+RW3ykni
Ea83zc2RW+FEpYDv4awCEZ2Df2zRMZayYaehn/PLP54=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7376 )
`pragma protect data_block
3kxAsftMPSUpWSPgmqMg/CzfQuyrbBhIpI1HzjI6UdXQrhy9tjg53xZvuvj7ZYQo
f16uRzwFXJsZsMiRpKpWT7mvg57j9/bwisTjKYq91dUBasoklogjBKXN3cWUSIJ5
/XI0IvvGu8iCyzQG4yCZWoa0MnhMgkk+gs6x1bQ+8ICFSW4a63HCXnE1GVnz8jfd
mnI1BPJwl/ijUlH17Q/40JW8ZFeiesyEc2DUCVM7dp0ujvcKIBKh0hN0lR1G2PcZ
8ps1BPoUmpg07qXyEj55CPQLJNlL0Hs8yurNMIlDcZ8rtfMNZcMnTMvj9su8DZT7
eDrRQB5JCCiKH+ybcocsVNQgVeBZ4RJs7Z0gU2vOx4QtXbJn3glHpvaXf1Tg7P4S
+1NVrbAoWyF99POQaUgGoK1Tk39X8EAGrHBw9vLu2l2akeMYHueUsXzbALQbX7VB
AhyJ/0WuxRLufDziIQa5yzDIbgUwwyqXpC+hktQu+3plsxyM0OOSfT1JyRqUXKn2
4FALof+RkyYzhh70kobW+cNWbFvVZ5j8z/5hmRSDx/954Ju5HKHo2gKoy/DE20ch
RgHJqk8HjDUfdZtQm17CChbVghEnIZ23iB+UuRNe+qQEY6TkKm/YyZdGAXWO7urc
qXsfznBJ30AOniy3MtKTsHpKzn8GLlslT3XcCm2udpnpH8tbmUncStMiSpbe6prK
WDCOBxvIfIP75uWTfdblDY/VWcAh1Stu79gWCZtJGAF4K3xaqlHFF+m/QhVFuIs/
MpJfKWvsi7cf+gK47f429iXbh3FYeG0hXcwI59OPzWGIwe2wR5OeA1xm0YhPPDO1
XWbAQQrYNc07qEk9+nSLucXDY8PWyDA0R0vYXmToWkdiBHz1exCAz824ln3XTgFU
X2jwltnktNkVnUrvo4PyVeTK79/rWc7qOla1LYgBQOI5zRotw6/wMr5vX7PSK3m9
tmlrxlOldI44gCuZw+//It2v0qiBts1P8Z/o/3aEBn8/cI4D24Z2nX6v98Udggc9
+J3cYIKS6PWpiBUDiAi/d1SMKMqrS6gQMauzPwzMU2EnZmCbWSc2PKCQ341hHRvu
KDLpaQ0ogJWOsiSHEulxwJvvnbCUAE3+wEEC9Y6nQmUJDDTXm941TiEm51LQz5Yc
F52/GhF9wHruPG+ZtzDqAjpZW0wNPfZe2YzFSYDPXDPmXu/554p81gur9pl1QGBD
f6pmeZDvpAtW3Aclv9sHESm6iSDWttoRYw1U4cVk66ikxx+im3CU0pWbD6HguFqC
NfEBOw5rF10wbokX8HlFkYGAggZYe6fHBy5lrwjlFQJ7YeshyzB/V6e29EYMzK8q
w7b0e6gqvfadKqQ4hchFjcJFMhd38DK6lmwEabjl0ikR0O0mSx+5P9TAenPKnT4L
N2rN/SvOQT+gUQO3VyjyP3diZK7nzCJXV5lqZmwy1pNS+2MQeOI4FdYerHrd8R1f
nT9lGkyMAY6zs3pklJ5y25NV1k88hS3+VslS7jW+FyfEMHM5p7WJ6vyQ5gsK2+2v
foghq5hZk7IibNpkJADv+XDjHdGtMYIRlmZMFs9GGFsC0+doef3R4VsMZx2Eyf5P
F+1lL+1A2aDHqWidBjWijjJdOp2K+iaaKFycTbYE4CTOhrzzLJSfEyxN2X1Zp9J9
B6icAmGio0d9Ka29p5gP/KTdc2ceeq1kXfkEcaN+DG8L4frkDUSP99Ov9RZ4cksP
RA6eXpEZRLhPzVryG4z3fUEdJ6V9EPFAXBXyDlMP1dVslS0ST8oT7uV+MdZ/jojb
yTqjTD0Da1AF8oXwm7UbUEZF07ybnfQIIJng0H4XfFxrx+5BmVbJTN9ajI46uunU
sttH3aHnFnP5kn0gVSixNAJByvVjTSpdJT3s0+stlxVdp/9DKyiirFy4iyafLEcf
WnpP7n8qCedoihs7HkVrbusN0tCsWZpZrsN8xFGOF20MQY5V4RhG4t5K0nKASauX
OqSwfDU4WE889rIvh+jY+mFl88JZtEmUbyvK/RshuOkC1nGZQxNECNuyGfgpXSnG
SH0jdNSpLcLBnEsahV5ZqbCkH2CLPoABTzA0jc+f7nEAOh4I0f74vozK0LLxd4fN
phHzzNSgHKDGrGGJ9pP3BCB9j7mfcjq6q8dlxCqEdfQXvCbqQhKdc3F9C0Jr5nlV
SfBCBH8qMbFka+TMltH4qU9aOlxzlMQWAcudkUpoUEJbF/EujQbjjm1kzO/KLU7U
hoF56boWOEu8Vg1zGbxIfed4t4MiPBPP6Q0jbhyRErk03cdSxa5jb8FG0knC3Uah
DPAX4+VR0QqQdyt669k5W6/frbIP8eNxhfEBdafGb0G40BwPLQXe+Ds1J7/lYhTd
kNRoQvrOEK8eR1IYMhUhtLDT0/ikOjmrAMNKhi9AP0JXdTjqQERS2a9MPpdtV0Y2
udarKbwlJvrTZedaLqR9JcfRCfIIga/VCG/uYml+6r6S1vHkonXKIDSISOb31imW
ZtnbYF8rrjz1h6avjeDRas9pAxzHwpeyivz4HZjVt9SeIcbpH/rkM00sx3uAyF0u
ShIV8WdRN0UY6B5z6ucHSvRNYHYsQ/bFdRnUG+af8+LG/yd88LdBLMX++4hV0pHC
yIzJewqmXqVp0OV7RYGGaqk+JUOW9oXak4rGy6gR+Hwj0B0A+IPrcuEo6okbAIfH
WQtVcM+/Agv/nwQudkOL5YlqcQ87NppIz2Vkf+6bV729xgXLSlQA8Nsfv3/9NYOb
rvpkhSaYQkD1f7p7Sbbdl416atIlTph6X1pi5PwzzEizXr3Bfu63BcaYAIhHJeNe
z480dsyupIS3+ZgrR9C0yC1ceS+hUd26M//TOCR0c2zmraSlrG9ihm+ija1DM2/z
ElAMzFGKX1fNQt8ZcPrcoseJBXB/qsXN7G5pQC/iPrZtLGbECe+053Cb+B9EEIOD
dB/KDtvg9+S992FmYLGkjfZpNTN6mNRNZxQbz99NrL8EPURmmN3C/8W/G06nbJ5o
EmFWcWama31kFAsOYsGOGRCWyBvv+TsbrtD6ZOkECMNk/B9MBFUisJpmMnLxq0XJ
DtTZnvzCXuR1L9aIs3iSXzzQv0diBTnnc4KmmjUgRAWKrdmLQZOXEmfVZSvafNAv
kpo/pSVqyC2HczGAU7IEU0E+E35Oqi5HYsT/33RVxkYaiAUEHS3zY5c6Tg/nDuhk
xNwFicsFFzEFftfrQM9pLNv132zt+PijdNT8EGcXW0bLVFpaqcB4XaiR66jF744z
hNIKBMvbgtf789BGteRNTsH2SzvSVZmcNC3ZAL55JXGhmweaueEIXijLzQfIP5s6
QdzApqlvgWyg7QyK+TfrXOwkvoDdIfGgg/VI0kuL/ZDbrDg1/WI2Myiap9cRoUqW
W3BIaVsVJvyqrUTOr7AHiep2t52/fHggKMaCv1VuMKWjKMpOiVTHmyT6BQ5yxULc
bFnBjfG+2t0PPvhz///fe0t0R0WDdtzo/mxNsRcss2y26xPgsTcPeUSag+nG4C2l
tnGuDKckMkWNvZ+LMwZXvrwlVfRiGQ4jubpkBPgOCXRqiUxg5w3/oPYH7nQzTuGI
HwYdFB+8qFbQuPsExXkYCrWGHhIdZzDA4z74fFUXkx+JFp6x9nfS82A2H0b/d3XT
DkZrO1XvUwG7padlLtn6QC8PjT2/QXmzw2m76Jp2Oj/vPAYwizbYsKdyWPueFAkQ
VR4ZAmaWY0CrfAkzOwajfIR3Tzi5XIRuVi8CZ73xr6QVERrOurmA056JsYP4NbIP
7R9dDlqRmqfy9LfQsdQF0pm/3s/6KAf3kYGa8Wvi2zxJXEdlfuLz847q5beRDTti
0bLu+0P47hv8VuiiRnWW9PGF2MWD49LfAs8mCxGMw4TuCObS4fijuELX1a3jXdEf
Ekxiw6MDUpuJg7FJhWxVev05g512EFx2norxQ/x1B2ZdqLogwPnuDkei4sklfax1
Kkh5W2VvAHy0VzMKmhKvTf65IACNnFLooKnHrBuLUtWkT2hsN3dTRwlTFo/3+OWd
ZHg5qzFn8U56vl6fYCSRwXpyTbFpTl1CAUog8Y6M2HEWNW23tcN8c+JxuLoJaz14
TMjy6mNoJPk3P3mY3+vYgeYHQ55xgN/JuM2EqYoKn91wbSiJkRN/0jLd5+AVswsi
z3fK5brnJRlno6rhtiHNfyqum1jbts515J5t3/1Nn7YeLNOm3lrc2uoNwhTseDkg
UORRvnpYNZnGF/8kURaKxw+No5tUSfjFT6L+uShboXq8Z2tQaEaGrJNxVfqGAxVl
4lZZ4/nA8NK4FXSOi9xIG13OSIJPLEfrfOS7D0Wp/LiyComBQXH6Xs0RS7C4lvEm
ecVPjtIGSCmUWianqg7QJoubWZ76h4fVMiPObpmPk+SoyR4BfYrOW1f1QT3idQpj
HsbEevVzgvqvpow+LnN7pafGAp2eRgI2ZWmFAxee5shRaoWYka+Alx2Jtwh94F1j
bTPIClNDtCuG53/90aaDY+fzD+q9ely2v92k8r9ve42Qix6utxgXEcX3HEnsiA7E
wic4OLfQlGqH+NVxiC+9fhE/l/bhudiEY3y7HT5jCHPS1kzfA0xkXQB0Vb2qROgn
sUcWUVcYDRzvYKbwCI/uMZL74WSG0WauQV0KJJmGS0Vietk2xKsWVBMdWdpnP1nE
MGYS2tH5Vhv0HWZLaNz1nvKPtB3lr/BBxZKlzdXD2qZMr/WFZY01zSMghH5Dx0of
/U+UWlngjKuKoohIDBWPra3jl6w1E5VbL/x6yAWyK94324TlYo6Hhq2Vhw0fA8uY
DidBPYB+O2SBWTVNtFLSxAye7Eqbl2ssi9d5CyeOFgQLZ6mQTfZV3TWeZ4tuElkY
Sh95O9e5qga1y/d7RWUGlDGSMoWDmZpGHYiWac38aAMwdfXn2UT9WnVPgajQw3G6
GYsT5ukPM2WdWujH7UVskFV8m1cQmM5/gJoSRdjOST3wZP2CGCbnp/iCVL9wxQ5r
YlHvhNgZMlORnlHi60m6PzK21VCoJQqhQ1EC5STpR3kdif7uBgOWHWJbLpMllStS
ymwO1JHzXdkxn+50IJ+GF4wQ0i1aaTe5BLlyW8iPbabubb5xtdY9QXDsgOBm9+8N
XtQOXtdGo3w8cY8cVjDJIAzUlMHude3CVg0DVdnIuHlh94cqmHsyT4M46ECiWw/i
LUK2h8z8mYqGX4ALJjKftqIm/yNvT6ncGEWiyrNDKBIYKgbtp9AhUMegqVWGgZ8S
eN6onOUDEbBHRRrDJJlTIdV+WP8uJ5uhYNLqLDQ+JTh8+D8hACdmuPNI2FIAbdtV
EEuyw0bdQlUCvNKqwuXhySg6BLV4C5KljcAHcKEy+1gR+p8FuzwIK6KS5P68UWby
aPifwcWbihHlLIJ9WoYPWiZMsuD25H2vS0Kb7LgLKMLKHEyR0axEKSIcBg3Sh9KL
dcgBI4HYX7MFgepdc06RmDFQ3lUwXkGI65KO7AwxHIfaP2cBJOXAaU6ovkoLhbfp
44EfawMXA0rz/SENRs6Mj37+HSfznYQV//+qqIxp0yoli/YJvmwkSv57lELiBO+d
2z2L2n15WChvkxYcgqrTl9XBW/KfHx/rQoIS2caccMJkT6kml1fdVGjhPmkE7ZFf
phUIn6yc3ABM1ZUhzqlft3rG+wJC7WCNSi8oxIoeV5wB1CoyQGT+iyIQV8+/EIRr
lJcHTGmtGRgNtGseEzJtEmruyEbrmO+U4SwV2xC/pergF+shEEDEF8Cqf9r83595
Wj8424PUHXgV11ClvqCbQfI+CtcSJDGQ0PWEMbz6tgOQaka01nfoFJdBVDguUce8
C0x1Xv85D0awlClD7zzkWvg779UCSPnG9wMLwgwFCn5rrXKcPFp7llapO8NBvE9i
jw6/5AuILSuOzBQOcOWykyx+1yptrEVWjn9GEXea1CaKseN8xV/5oA9uUTQQ2AAS
V2XGDvWjXoyoxKrOGSoWey7sz5OECEMYKmosn6+MGkFXhzdDlUjRfp4W6oRJUk6B
hhPDDEejKqnlVSTSxggwRM3C2RzZkfEIyyngstdSJXq/0cMCCdTYGO/zkCR0Oxa8
jI1tM1YKb5KOv5hDUyU3rj+Upwx2kC8ukZc7OBB52wQuNTNeXfcDFzVmctQGgKUZ
7P5f0g3FaLcwcmkrHY5w4D4TVPUZkVAkqZwT878xH087BlPIL5Ncs4Dxfh6RzYay
I55rzJZPcodmQwL3PD7IP58jIYkvVrYsKcHCF7SSuwtYGkDGyCHIp1JA0DYlzzS4
3pvPBbYuzC9mmU4ikRbHoGOiIzvd6pwLNLbP5tzZorBaBEMtxlEAxbVrv7anQm+v
druAjJYyo8Bkf/1FbW3SS3JAiRbmDSCbU7KIE8kySfNbsJubAoyzZeWAb2uzRiky
IDhaL1Fs/hSD2TS5uIorC6gZ43fV9/xQzJwfBMGJNnkCEZ4FmzdlrmTbbhIHDb/S
dzLJChPp7vHJW6qv0V3XzM8wMbZjGXiUi7PPoiKRGfS6ZJU6H/mwGAL8qTUng66Y
kC2iUKJyR2iwYThMRRr8DW4c4sfeSKyJo1GL3uGB97W5bQ1PScqv/+xzxR+N9a3e
5B+9emvJcRoHltNzW33rbC5Jmx5Oir3BJjhPwg5G6JghCRSsjOUDd+niEOAX1SNU
BJr3BnhknzS6wWYFE56b2WzhXX/3oguYAs5zaRmvfWf/m8IZZeDGGdSWb3u/LLB4
zqhLeNwCj4P+IDwFkmd8z+H4bV8pUVc8WR4Z6MiAk5yBtQ8mSH3QMIHU6F8pduwg
vQekly1Jizz0t6boCFTAMQJ/rK9eizLJVsv8mfKrsX7scuq7UbatRoaOhKi46u7D
xCvmTndjszfUnO0yGVAKkaaSrB/IOP2tT7WQSNQhVkkPWWRiUoOJR8y/wTNNGYPx
gG8U4C+cRBt6AyP0SirFMGgazOhiKj1ZZpdSwmLOqnApdSb0DgD4+NUYpvIjvrgy
DJOFvpXEexOB1qk2cv5qINxwOLDz8VA1fM/aNVX96dFBdVkOQgU+eYwP0edMV1uE
YaWUjCr+kZrCsZGD1dA3z4+lxDQGokvNELGYUIPkoDoYQAvDz3TRN5HGDtZ8PRc8
GAE0hx/aKJZE9/nxWgMJcFaVkyDInDt1566QV3rJKqDNZoZeiyXlZjnF7rvNnm9P
qJSG01cBqIHGXcVERRn4WGRIsnOJXG4xKRpZL92gZ2RGZQkiM81eJkInMqpS9MGc
DYK7xXL1bBOj32Z1KXRtQlEhmRJbdI/ENhM4As6Ju/riqh/toGF0RfiFIP9epp2k
znbiHYWvQgNZuSP7te8Xa6riF1LI5Uf1eJi23WNMBjsWJE3G19RfmBZvpV83gyub
cTapykidXhhKciB7SZYBg+1cndGVqkP4PKRpxnd+dLKWe7SfTzVfHihdNUCT/OZw
aHJIHkZde1UHKOFyKe8aBg0L1cS/SKkLfO8FGDpx8b8bHo9wNDVCrXPwdsY+l8m+
whtKCSv9ig7sSUwEeuM4RGgOwvd+Q0BvSL22PXrksO5+O/AgTGnZ2pgOtnw4RhmA
eVuux41AafG9+49DWqPtdxh1cdvxJmCVWxY62DAX3i9cqeO02v3A7t5a2A+I4fZq
sciXirXGdRodhOMVSKFsBlEWDF/6vWTpZ5EcQL1BpzgrjGxS84y3G2m48ffims1O
Ja8axscjVbJiotScQFs+x1tQNiiuJwkDTX5Yyb0ZvdrPG/tepI4z3dak1eVt2RBX
W68PaSGhRoTyzK6GyqPC3uQOFGtRb6BcjqOkeMK8Hgs8hpx1hzjy8ju9Rv5lmFnh
9+4iLIrJPhr9eP7tqpplRgOCbJpep1eJVqyQUkTrP2sHVC9eXHGxW85DvO2K9lML
c00RA2Z4PYUTdimWH7vGfLwVlu0YAvtoeHa0OlcWKg5lKtB3MUU8IEb1Jc8aGpAn
yOWcUAab0nfp/2Y1yVz/cyvrAMRmF4+VxYHEITslVVp7XIQL+DGhgAkI6UZg3OcR
5FUBJ00z6PDApkM6rjpToLUDoTP5oK1B71M77diBCGeptRGVyOQCmE53/MtfC4WP
XF2PYhtCL5g0M1B6XpSwU6x+2rJmWjWxys/wifki53Y8OgdK10YlGg+caJj1DuUv
CwJAN1eXBEcTV0wWDDMox+paSgHG57yNC1zLNQmmpLjabyumWnoG0FRE0t+o/OYG
1NJhvMUGpTB//EwQdbjWYC1LHjvMHUrMza0GLZN5BRqCw/tvX9oyNSPaAuzMccGQ
5UluY94dZmDRoSJpCKDmWoAi63duT7/1fAF2P3iwppmxPfsSu2/VOo1v7wmvlV4v
PkbnFTe2bcr4wcjkrPm3fI+6tpg/0jpHynPnuempy6TE/tjlgq/GEg3JMYaDEBkn
WAJNr8cHZ1BdkuJL45lD1lVEAl0YiWYtLzLe2P/kwAr5Nf2JcH/h9IEqgzbcfs7z
92v6eVA+PfEqTRCo6gExMEVYjyCClnQ1DHaIFX4bKxo7tYIjrn+SfiTx+Q8DPjwB
oFc7L7FBmMGzZH4n/SnnPi1I8fe3LgAxZdg/lMd+HteoF8MDN8YiRgewNVxninF/
OMaudIM3/wLbsLabp8zyhYMPkCZ7vZjRQDa5mPS+JNkYyIcCahlZJoGFjLuF9sEB
RQdfpOlKHnp4TP5n1aZ0lKFWijbxQ59qpMOtjPBPdEU320k33wFx6qgsjvuZd8ul
k0NUhLeSX8B54WQg417bSewS4De1uSJgrxY7oMwIaAaL1gcJYFje2sTZyG13AnVx
UDO0Jkncc1DQMm2Mymt3OaAXshis2SxynurE3d7ZsYL0Y/6GxBV+nkyG74KbKF7S
IOL5hiUg2IYJhDHGznaEEoe/iHsFHWMOya1s+Kn3Vt/Nzm+SaDxWUkejpZOTia+m
nM0o40YjX6q0GF3fslqP9lxs08i4nNE4KbDdKKmVzzADWoW2nmaGzp3rQxLp2GJf
TSFqJNtxPgmN+vMaIaqr3CKZl6tZb2qSbj4K5C5OUmspXf5KL55NYBFBinRP0bdq
tTRc+u9wdOhzgQIOfUJHwxu6m/VrMBT2zAbkCSr9p1pUu6hGorlu1+h0fH73ozqO
+9nv26R10RYaDdI310/KqCLDKyWAO4csIaKdR9M7d7gk5FeQat7UjlTjgld2x66v
3T8LgIOUkMXMjFPXchx7f4juovKjgFq2cdiSdFVG5jZi1V0GhiUJKZ0Ho0ocyMkX
2Ab80Bqnfx4BZihD+eweM7YWZInZUbra14dUegDiNs1AwjBKUMvQidkG8T6rOlDL
+uXl/WI2s9QFyGOSh7jQ7NrUPzCIjUQ6QUBMCUW5WZHCAOd4Z6uCI8yw9sCbJWxA
vdm486PMN8r4Fxjpy188P+BNG1LwpCNowRCOBgW4VRL2fvWZk0FqP7sasOzyCl2K
Dd5y43TKe3ZkzxzEARTxKNsgR32W4R42l24G9amPINk1gAC6oiehHfz6Vpem7gcT
TyHZs8QxoYdSUqMopJr246q/XVM/z8MUXiTge0BlgcDZHLy9fFdSu6ygMPZmkrpA
XuK6lTX5q2WrrwPlvOrzCFNM12Sb9hV1tNHILeFC5JyWRCUiDmMxxcnbeZ33h7/m
lff+THzLNwyUsR3aR8gzcJxMUgArA/DZ/b2+i6AD3VZ+B3oYESvDqgF1KM1G7cBX
/s3YgwOsBzRR6p8/pqblLdw73PQd3Lo+lClPS2Q1EozHV5qu+zD/aUSlVNI4zJRV
bV5sgT+RHO8NMb19i55vfZT4W9XkDsU3ggEy2zWypYppqacTe0xH8DKZexWh8LZx
CpJgkWh6kkNcHvLay8iOxDm34cCUHh6zprQzrMtGAkM=

`pragma protect end_protected
