// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
CJUqrHc6Nwo2v0hvhGJfVMvs9r6CeuBmlpZBohfS5Jb0uZT8/+oqygOUNZbL7fJyLmHWq73AEiCZ
ShPF46NhLWVEZTnneL/zIzWZ1pFCCTr5MA1LZgV8duSe0FU78lm6yQ81kWr1D9PsqCQRLtgZcS/o
+GwK5AJsGj7fjXDRSScLg4qUyA7LEsBMdhKghz9TdMovk5+NN7OuH0wag5Z9se3/SgNAYYgrfVtZ
DMxO7DO7CPMQpD6zX8dorFNTVIYg/QXeE1T9eEj1ERO5YBCNVTMu/xGbU7wsoNK/ErEPeh0FbPfJ
w4zVWhh+RAGDdnHrvsXvVxxzLALHWjPasS33yg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 26496)
1GDk0DlP0ihwpK/uGbIGzlv9weLd/IZCcGpdDF7NRiEnZUy5DOmbyDPvNTV0XYYZ5zwVapZPs0pL
rpvH3zkYrwiEZG8Trps5jjA/xqD0fW1JhspEmCgN47qhkqgeNNtrIDU59wWUsCSv9vtKAFga8mP7
BxyFmicEXwuufIspyRIY/Bk9JTQLRaSq2B23G36kbw4k4l/UfYMus+T8g5AaS2GhLjCJJL+GMxX9
Xi1Q89A9+CCpg2vLFNZIN9gkcF9fJoqc6f94aaAzADjqGd+mOB1l55dnZMiFu7x129jZhBx2QDj6
EpVQT2m5dY7vFXgusFHS4HAYHeOaqBGLs5jhCea6/4BOaNMFOwoYzFPno3amKuVnyzjYtCr6Tq2L
ARVToyU789rcTKA44LHJCnN+uQNw7JV9BI/85TR6NEEtiS3RqRFhP2YZTLseesnIsKdtk68iWMmn
WgrpOXYnaMygtTNWcqFQeUT9japQ4jLI+7AzaSPsW3EzmG7Bv9ULbpQAnF3bBcHqUUKn/waMP36g
Wf9o+b6rDPsBdyyhOsyRoFy8RAwqjd60/FZeqkwpPHrh4yFeOL6SF/RpfCCFvWTgCxPU2vZO6tvk
ngGYTBJNXweBAcB1uharoBrymtWoQVlF2wUCLfrERAex0F1nGyRhETBDD/R5X2TrE5vRv5/ZKmUY
lni+/BdILFPt3lPscrU6DFmDrE6Y9BlBpKxejnvBNoYxzxdNrjiVKI2WTBDuEK9mNLI6RjWMepjT
alOPaNdtba5OnqNu79aH5iPjJzNVefVntqzgyAmLAi2LQqQnfa/OD4zjfge7ZGXGaMDJgdDpnMkH
9TuHO8itCX+I9yUh1/LYsJ9qLxERYptu5/m9s9XBzkqcPoVSOJ3zYFl1miN8nDAx4yq15DDJcvTA
3kqRbfM96DC2oPQwkxR3P/QaGMcyHQfMlRIsyIaFr5k5aJIFwIu+fBJnsdqySG5wFVG+w+1uyGnb
rv0wl9pBy0tafdK/Y51MGEABFGqJJKwAhu+o27TOuYq70yiuQkPatVMvBs6YAzBO4mMtu7zZ/kNn
fodXkCNHY41LFr2xYLgCnE1lu4YwS/o0MFrhwfmY2+/FZbtE8m/SXDhEy9d0/VTQ7eUva837mFhb
iZRGa7kGvkbbGtSYEFQPwDQTv2WuxFqhX2zoKMoQj2E4cmW6NTuxbQ+O24gVIZRnCxYK7oydt5+q
YJjm5DVjuKSmIx/cHkm2xarhGN5gC2cWZgpYvi0yyYtZ1eaLKcqcHaQvxsuYXWB4MAJhKJddTU+W
SNWqXlOtVcNdqKBsogv7H6xj0oy7jn5k6CRQCF5mVvAkvGjzZngTSJx1mqwnMVs4GlyW1r3LdIeX
QpxeHVVM98Jq/TAaNv60BhCJQlkfmR1i/DtUmsNceLuSxzBg6P9DTS3VJP4OphxLGHGqivfTlzxx
7NcpHQjhSLbq9dqBCURyXFxpK+AwhfMg4OWReqqEgVCiMECogOzgJ9LvB7MCZ2Y9Xn3dWoxRdVgk
myIXAOC3y1bn/dy7uKfJCSEq+3F6f+IK57CMUTos4e4B7+ONlFN9BHnN2KQ9kMJNa8Gb3CROL/5w
HbjNZ8F8cHlhNfsi5qvsrpTf8sTt4VtIiqMXsWpHtLwOCmc75QZDVBeDoMa3vSzxEURbYi8KVlgg
ir2Yb0cYcX96hrR72vGAbNKqrx5fy48DZTFTV7DeOw8B/DrXEk8VVd/S8CgLJhs+LJmYv7OloGGM
bEBFAdxaPEkZkC4L3//zK9h85BpbNQG+QuyUoYPgEYoFdY3jtCgGrlT+KMYNqy5roFOBf32nYK3S
mt/5Ek6Aa4U0V8L5etPv5peAqbNCWpDKH8PfMQDDlYX5ApzzTxbQ0JIs/Zye9rIOTsyMWqX0GHPF
Ok4RAumq2VOaNL6y+B9SzFtUT3/V85Ika1/7JvcpU4HNU24LdQYowUnP1S+oUWD4rgAw9epJt9mH
8le39gPnUfBh1peDskS9I9RAQaBE2JxKmJbv+EkQhajxtBJsk7q1CmOtoIU9+A91dB7jz9MdI2hC
B5/72OqbB6EMHL17hqygHvxywEIfBAusChl8xPE7eThjpHmWIaYaS+mQ5K6Pe3WqcDuEFdvCwuG6
aXfSuwvxWRJy0bhl8bKd20JQiEcMvCvmoIfYF95tZWnlXRsp++pxv4Tji/Z3HE+4uxhkjiATonrv
fhq6PCMuS3k2Ur+hZDXUfrZIuk4jZ87UzTshJOXD7vFjHWw0ySSArYOxy8QkZOCwoS27q9PS7HkZ
bCZRfOb6PVLj7ou1QI52prdQnGBu3Y91Y7UuUISR7BhUYCPghnLSj2gGP/Wn5g24V6OKpLUFFJWK
Sdv95ei+K1cSGPLGSBOUUmT68Pz1UVTnmgGqq+rA1D8VGIi4yyp3/nw6yKvKMHKfu8WOVc1EJT9M
9JCJtrxi88fl94ooVRglBDTPFwkG9pSR1BMjEDWbGHcp4IDpyZhcwwkmIN3CTcb5nhQ9b9k2wzXa
IWNSSfncgRG+yihHvKAGMW9BLcKabTGuVNQWE9M1SXbvWZH11le6NJ7gLoPZGftPa0naIv4uUBUx
xpB4b8J+XhoyXUCR6Ah5tiRAUPll2XEgte/1s4rlupXyUjzDUkp0IDZgicWj3GlKqWodmYRs8ENi
9FNStX1mqoKNCC/Ag8oHVAToBVA5g4E+PbLj4q9ZZsif3QNAdLbgZEmE4nvweVy+n+FaDxe2h8CS
f0B6h2XtvCuuc6Q3Tj4qfX+YoGoM0N3ch88MysgjhiV8oRvREo6vpvmgUFx5F98zkvQBDdPiouzd
EXpJ+RKf7jKPU/BQY+c1CaT2tq5RC+iiBSXXvwGY1hQEMTcYQL2TgLXTaYme2WTAGqXdrAaDSnbT
e7qPjlkW85qBhjM4CnHkdjQ6xmBNDK9QE2tRgy9bhLV8yBmNXYv+XZDBlyzF5JUo6fcxgVlr82dL
RASoEABq1+mgOjnb97rAv6if7Q/9KYEHkD4uh/H3hAA5PHFYo2wklsyLLP+hWt1QRKHJ+y/Zhy1E
oxgMnkkGRKWk43m6BebpibSMJNYJg5mH+or1xuz/EmFu3z5TRbJi3a9EpAwQ9WI5BBYgtAc1oVCU
h83MSV9FvkpwyyZzFWQixfw0Z0aziw/6TO5GLY9lWf0i6PhmfNeLaPR+GMflyR6GLydtk5KYktdn
wMFnyXIkJYnUqv/ZpF+TOZVZ6bMK/BmRfbVSIl/UOajdFoDeYSVKFTvZYk7B+P8VZm0KxwhL7Ku/
Ca3oP53tCYXRCcvswbrPYX+grsGHiE0GwADbOu3Xo/koFvJYYTjdboJ44AVgzKC5cLbJUXusuuvX
cXxXUwEy8Hn8RaJDMmfokkjmFRYt71Hb0RcCkkVOupoiJo2drRemlVuujdjbubAIHp6HJcUqj+1F
Dz9akGN5yRET6M6pJ0KU+LlOSF7n7NWZBPoQpj9v0dZHIQEUm59dekr/JfNVqGnE8SW1l00KgSrJ
QNqD6ZvkPW2T/24KhpPSJbR0DhK7JRU9OY0u3dq8H0/CoUWWnQEOIN633pUP7F4rG4yPwT5ukh7I
WPAE5p/ou1tSYAc6qAlAofJok+k+KGx0Z5nCDxY/2ZzI27MgoK+6Y1FA1vbZGVtqjtHPe54qJYLo
SLlEDa+uW5Y7c/lM0SNrijITGeDRCu4okHZepLkPD77b4pfaorVwD4J3eRmzGZCrOmZM8RwOUzsQ
R7SixWwrAet6j92AJtzqz59duvx3Py58ovq1sup5rs7jBji4I8yxyi+HpVBNPyx6b4WE7PI7qhXw
y3RDmHOvqY/9G+totux8Mcfwmk9Bxyv/x+jlou6WDQ0uME5lkZbmNSfyfpigrlJS1cBuVR8HAxSk
HZe0Kwngp6vLZxS06rbdbLSbmTUarBaaxj4oJvtYQ0DIJomH3n0vPOJGRNyEP+R4Yp2lh4wbRoyq
Cy6vcjXasnYJhtbsp4yiB/q/CMZdEa31ktGILgERR7HmtdQcgqpxXGLDDXIg7R4daDgvegsWXsi+
dXzO9Pgpf48RvMKioqNcbs3s1WWw4EovTsYLz/9Gp8AfMvNESTD4tib2ubmVTCi2XpUcc6JVMKXM
NqYolB8mQjSokgFY8GzhOs3HlcCiSY/vAqXyXfDPfHFwy0lNUv0G+3tukUDw4XqypzayjOfmx70O
XHpg1gpzoiWrZ3WnwDPASIC+dyaGsutLhCSxq+qUwdT0W0YrGJauCqJNO+nqjlzYmMi9DU5/NkkP
kFoIpbHAzZA24qRbaq98emKUqDTGk8xjnECFdmVeTiaSW0PrLX7EOMSwCeFcUiHaGt48EBl1CNXi
2C1kYVlf3jRMtuiAdROXLMVnlgpLZ/aHAZa59l7NFo/sbX6vkDcrgHNVJul0pwHWSIRk6Cz0ljJ3
310fIb5SKb8u00NlEWSab9bZJwo8DJJQAtvhuO5gUhlAZYFpb1uGHHBj1LMO6FoYxXti+ynvGDik
ewXvSYkES6OX3bRnDBUhUHnrB/I6xeT3YxZv/sSL0m6xXwMoQ07feXcGH2zofp/Qri6IUx1mACy5
zH0Jh7IWqeXjw6GWsTzRj7S2I91qzuQgUhCcmPQlLZEA3DuyazBoxMxbJADujalru4mip8VC1GZw
ONuPejxXZ4sOuCwPnnb/27KyTmpPQnVCgucJshvzn9qfrvfTM184A17Cxz0IrmPtExdQnREWFsZe
I8+9sjmaejXzM7f2VKjtunISwVLo65yI5tA7DlO1PksxiMEyNBbnmt7P8aX6hsXXwX83tgJJKzk3
Er8wKjqzOdD/AMmmWiUm9QE0iWfl//0l7MJIvU6T5tjl3B94qwrUXFf0esWu+X+wTyUF0JfHJ6kh
paQFttBDZ7C7RKmTC3fX04KEC5hqXPOFAuTgVvhUNnDjQFxp0e8393GN8ZIPUN67VdIvr1L0CN+T
Oj1ShiTh3FwiOH3CNgjqrFTbWFBh5Tfg99fBxY8MBAZ123gklxhlM3+l+H7cICdwqqS/6rEEINnj
4CWYM8HxYItZ0Gt96qVf5wZZyTiIdC62hwZ9Lr7DEEEZUtzBvkuTR2CSLoEMUrDVhRxvwI75eeyJ
ppi7IieJvMWUwQRwBVXtXaBd/aIqIKHiI+SfyoFVBFbX7ZTVLF74jqYffRXoxDW4Tb98wb+/fJOS
knLGILiymI/4bFUzVdHqILizZhOVzuKLPOowm2AjruAhfobF4bKZOoUj9AHBZGNnXu+KzWADwikJ
YRXc/dQcRXr7EFy5OvtqAXo6VEYqi9O5QJ5epX6xwOOKF+Ij9OATB6pDX8mUq79XeJmD7Zvd2F33
JYL/0/DwUycIpcJgceNBaGKnUvUQurEnnlBWzCQJqXNm8lTRxRIwtSTKx6HLGhvalq1fxJ1AjCT2
Ite5QI10coR9NtaaRnoFiOS9C6IX3goYbb73IRWrnQaIHILv0nMgDWunDC5S5hQ+hTVVZQaVMAt6
xyzY+aJ3JJikp1nW5FDojrk6kJgtxUNgBM+yadkxPIt0KXNYW+GTr9ElHQagKldRzWOUEfbXHDQf
3BH6ypcFX6yONNbf8G/uxtc0pdhKULDqkWzThK962or8o5Al9e1klcJmxwNryZp9J9K/RN6OVJm5
Y69mjlBeFVe0tnndvbqE3aqjwTGyanMtSpVQ9KQGnfTOmGc5g9h4IKD5bXs7LyUwYpdPt0vrA3Vg
uK2j4UIR0IPNvSSg/CvDk6C5cRh6Ic4srqMZU7ZtqZM6Zou6zCkr/ByneUXI2opny2DnMYQlOSs2
iqloupMI6TlZhJCvuqd0vUeOmgKQtVFtUhWTogKTe9RbnKdLGrnR9S3BG7NgXrGEJth7QOdYocY5
vxHdb5C6eE8l7pMWMsrR4QUC7jYqWW2Htu13a8ukx3i0dE9Ltx3AVeHjyqkP2aOMH9NES1ow/gKF
8OmE0wudFaIl1EEZd9LxnvAF8GaqtFKdnoWlAzjLnudM2U74DWLWIbldm3rA/kJn0aR8UlduYTDt
cdzOmshhjoD2co4EJkAztElx7MMHnaKqWkXSYPYyjPe/JK1UMTi5o7j/apiRsC1C9iitEF9Q8Ctt
WSoQRekDLwnLuc9qImQYAok75Zc2886B9u2Q6aQpSrYY2xif8XPLiTqF604yiRVx6nqveT5eHX7U
fXlfbCnleL5d2gxT/jlTuqt9F8Pxil4FURs7irOI4gTA90rO/I8x+mzjniKvkevdlhhgB+rEWoL5
Lo5DzvvNE7xd1JzEvvMAelMwoTJxp5KnqCPM4zr9o7hGmkgdTbch7HWG1JTfsByruqnLYQ8rYkkH
FuxkBm/SIjGwFypdWNardr2wHCytfIw6sxNL9Gj+IxsP9HjsACm2sAMSo9zKgWP+1nepwEgO/A15
O34lo7DFB983QB45+W2qM1CD6Cps/508/oXSq6fvFjne/1w7w/iv9jt6n0ReF3FQUZdNxBNczy9N
9sZ3H2MAXjQEQ0YaEWMlamNNxgIDFO57eD+SQWxMMwc1ycLcyBofS0KmBMytqqj40m6fO6yH1ICA
t7VGkTq8VaWJt0Q4+q3yz5r7l3PjMtTQTtk0KutQhp7iSZRhYLwlbH3rhN/7v2jEjg7vkrninfuB
aUt8S9j+ts88hO6vDW2EnhKcw/z+KlklEWa5yYyvD29h+nNby0gz9cER0GWszRJZLclNsvKM52+v
2nUblin1hU6hh4yb7MchqZOs/apI6a/FIHao1VIFscnofCPq/X4w98ZrLvhO8/tX1Nxt9gQ5f6Wu
dCn/qvkMbk+oKbptAa9l7UGJZimQsdS7fi7CUH+w/F11Kk3/2IOcSp6FSrUbhN59ZSEngrfYFjlh
TBFJj/tT8kn4YmPKhF6YYtaDMSYlGB+hc+JGRcNR7GbOJLCfcB4MjVxcnCC2ZTqyYmcMfa1W+I5S
pgCVqQDX8Gp5JizlqZkqPugmI+hxKElFg7wIm6tmH0HELefK+2xnRmgeuzEPbknB0ayhMRLKbWNp
+AiSacPtLe3dKk2FL+YBCK8mohvs0oLHLKTYbpfqtpVMXTM4TNpZ5Oc+plKsxUoj7mB9rzzHeWyP
OswN3wpUegsw+fK+Izd8r4/XwkrpVuKbOkC0zF5xmt6DBC1amQgDA2AbL8RDsiY++1apHwh6DMXE
Gd2RKjj16lvTIJD22r03KXmLRRxj81XbXd+kOUmtsv+A8qPugJ9IWvLVCLcBdn9H3uAGwLij6MpH
vTJ9XUSZHI75gqVqpJtOkrKhFBMV1hft9zajX3dXEUG88D1bEwEwek313N+iQOLHhU6ndRjYXl4E
6vsqSRhvGmX/YJgQWBsZ5YZIGPtyADykSTnbpaWSvIEL6tQZvLmCGJXYQEgz5RloXGkAxrs+divE
dcHIcG6BvIJ2cOFhtHGFiTUEoUaOWXi/M7ybd4ebvg73CbZ4BgdmVShl+ZTPfxPQedIM0tK8T3VH
IIbluttk2TEox8WYOc41DVL5PQM5mmhEIJwjGPa98VwddqRSpp6+ZPlQLEETYhqzL40sZE5OLjC3
PZQMaI1ZcMQuxa5KrwmW2fVC1be9bGoBv5nroygi97tAprcohqbuuCprR2B0XVQ1U6RDvpi0leCM
wmIX1aoCRR4oYsw3t3QpW4KDsAGNCAkf7lSze93y6XuIHOgOB+oHk4aCxMWwXQMvRnxToc+N74Az
WPx7snr9aNeq3KcTVx3CvJB0etBudZNc3oftCNML9lHrViJwveX1kTyxu9QdjETH+H1BeJaX4HUd
PlN0CpM+O3vvRxJ0KUcobb3B2+WQ0U2N/gCFd+90GDdz1BURymcoXU+X5AuHE62Q6ETu5Xp82/vn
lrGvBmHGLtBVzzRuqXwLbcFR1lucutgGFgFNOndPAqWHFoB2PCa8d0LzyACLQd75Io7MAMr77aHi
jpBhy+kBhu7dH0+rufWqWVvmuX6hNmD5JZv+Ps0fCjdkY5mhRYOm1y8thdeGNZXcJjWT9qhXoahp
IER2gERGPYEZXRExQ6R4X1Sx+A56/w586W6gZZ2kZrpWNZyFByy4rCzxCjTqLo7BfVy4TaHPMNFW
lcZ49OQT01AxOw6Q3Fv6nX0wIdLujMZ0B64tTZGLd4wveMKEb/zS73G9KXOGwBAC/Yq2567oHBDw
vBN/Ik2ihqwuPDy8r/tFWbuW4BRnMLEXj1CxiBRGrti9BvBSmGTUybAR/KOCcNYZ2AKuu6HXs9Q9
J/WN4wMWh1nytGykjNhWB2s8qJxXHteOawbAPsPMdt8AWLvsifEtDFWZZQBr0iwSgLyHQkk2eZtA
GaVpHydOOieuKVLCmfJ508CgQsrll6hVkL8ceWEdb52JqGsy5Z9/qlm787gAbL70CrkTwyMuRr6R
RAFhG6d27yS/Phmtt/knQpha61SkJ22+MWW3QdddziPuQopN/TjZv511AX9YkFR19nyb4hrfGkwP
Xu1PAdI4ElolNWww8G4PGceARGgfNvKHq+yjE9idIOmvFkauep0YIscpvF7+KuJ7KPEVmorAaPJR
Nm9ROmQmyKITISe9aNjJ7xtqoaVmv//hjV81DM/j8jwF3ydoy13Jydc73d9BsClwc7yHhny4CjKk
n+jBJE2Bn4foJ/vairlbJsto08nxvOeujOL/5cWSdvyBuFMm2ly6TllInMRevQan50hFuIiTic62
FUVSMYpChEMWNiy6JNXC8X6f7BZEZLHD4gSnGK4GVJBAs6X/nexbSJ2WMHWeqlmyLrqejwSILDX9
R7ozqaKx8/k8aDZsjkcXFu1Iw4M6g6zeGQLehBlJYWZZQxlPSORLB8sxbcLt6vFgIEQXGSj/3cjL
7CL3tUkK8jc1+TaojmoAzrHNpzGfA6YyBCmr4rE1iLi5lUIA9w7X6B684ERs/SCdB67Vl9zheHnf
dpQ9800WIEUJaYIRSV11RbdmwoL+hO8PWoqbpx4URGNetwTF6ybwjZn4og90BcVQeiwtJzaijkZ5
k+O7kujEg3IgJgKP7hNkQxocgPaaTv8DJT5+65hKLb0uO5noBCau8Th2lwDLadL2EraohUjTij3h
JsReSkr9EOYlkJ8qPPoz2MLz+FLvxZ5lkXXDWRZ+mFL2EcLxA8dEoUFNPIauMDGYM2AEokWeWyUO
CcmJZ/0IllouG3HKy1qJ0pXoMZhoK2MATRS++eudTV+pSk1BsfelzX87wla7OkBWze9UdKr3NwF+
Ra2jf1jFicDJ7A3ajlm/TCTtH/EoemUSfw/EF+56O9LmHjWKgDJS0zMYFZ6c5andzr3PcQZ50PXh
mITgceZA4ze0Q2wFJYwUGGsQu3eW4LQqzK+ZyZ6C14/b6qbsy/espG2cnr45I3RNMlbZEo91u4eu
pRZAZ9tP5IWMffbCYBxwYgPKlhM3CVLo9oRxNKf+HdCcpBCfOessxTb4q6M+2XI/rfqYgCdgw3MT
92IKNdmi0wVXowxepm6Px1BwvhcONgItcceeI+QitjeFeCkXenMdMpETV5Gil9OhwEjVnYTNIPkW
i1prDxXQDMj6E9mN5Nx5hW2h8OIg5Qnr//USAuhnZlXm4QKgNHWHcUyfH1mBMd+Yk8YXCjP133g4
YyeV4+ioBPyC5l9EAwoTcYG6U7vTUAuC9keH98QQao4ilRIx0+Y6F39wcLiPvXB3VaCQD6Vb/m6f
UvrZU5vil7cSV7t825GuTOnplFJG2yRu6K00dJtHUDYkBUNczrnTQcPzC9Qb1H+UeuV0Y7ITbGcN
qXXNgyNbw04YqZ2JKNDwzBOkhzsHt9X1xFi3qwE8ox/bHUy/oJ7O8O+b5Z7yg953CwlVJmpGhR/M
/wD8p9h4+Ilx0u+FU0jk122Th2LbuFBsYWXmdmqs8skfz0wP4p3ImTNA+wpUS27wpcapo9ufQEro
mJmy7I4H0IP6iGTG42+JC8Xpo6d0LAgYodYnq12HARrEWe1ySHAXJxZ5duXVB3K33JFRqQ9+m/De
6m0g0QznD3CoU+FWJ0fSbcwxVzixt8NAzX9nv0pSlE97Pl/L11PAdtFkSxLZC9RH4fH7ZncPwBKY
yV1AKc12IPW3lIY5IuCRFG2TQPDtgcyqArVOFCUA8+2Sw+HE7LlZVujXGhrCQ5umwe8RTPdg669h
lZV1dD9G4zrdnCYEcUoi4T88Et5aQwA4tXURym7Rv21sypdkKNS3fJnXWIC4ysXSO8MnVsyJER89
1xADezKxGxmyPclHvtnL5++PPjTCE+WeprYCAdgsZ7tgWJJS96e2vWHO8r04FAv8E1As39aGFxcX
fE/jxwdszs2fWorzH3YKcjQJurDGkpFSQQ4o1/ZbgG3F89iMT8pzVEN/kPn/+4CPR58nyajPjN5A
Ugix5pWaXtzlN5sFypIPaxXMT/mY/EKbdx2oSDiYZq18koHh2IlMs4aSg/cgEKXsoP+Le7nY+Eb8
XylVn+oRKHtjTaJ4YQC8NVk6sIqBSKUdfEO7KzAfj8juEMrpxYVP8626uTxh9g5WyuzTcZqUzOfv
BuFwTGB3kk910E6N9vFknOMbCY0rlTcX+paLeksGtraGCsAx6cuIY4JSq4KaeomcHqA84pi3P+5F
8nu0NFgyx/wTUBKumtKaGZZy9eSZyx5pBiFljoIg99NWAK7zAAd9p4FtmGB4UVOC2KEqD39h/VLF
dvb8vQqcEsIAGxMGovLMP3lmUOdB1ZFtaStJYQ6V0sfurUK8wi1PcMgup9VeqTbR/cdKsxVTJRox
HqTsp2x3rDEwOoUT6jP9DQFv+6MO1pSQ0q28NT1G0CjVXastlnscEruXjv5MH1Lk6d0ROn+5f4ZH
d81FGRVuiFEqiwT3NmdcFH9oqRMLuQqEeK23j/PGjFKAXQI6f/UGQCgloMHSA3ziiuadLMUyMsZs
CssDR/Y1zm8WkLj8zSTvd1CdWUpTJwK16zT+/CI2BWpJFAkUsJRBYrN6QAuTlfySrKboHnU7pT94
e1aQjRh5v6Wa7kAZ50DY/dQcLEcNi5+Xb9XUUL9ooOQJq6qdVYNCcVpjq5WB8mig5gIuOFGbqEOG
zmttf+P68hU2Wq6E9OD+4C6le5HtyYgB51yrkv4UiLM89AIbZwOJvY10t1wmVGoXlEM8dN5AW9lv
G8NySVK+x1zzO+LTgpraI2DoVd3tdYWE1Xb3bS7QkeobDb7cWkdZpdeETtvl1SIRvu6ZqYbL3jiE
pGUfk4iP3LW1WkO96gy549gXoycwzza+S+hTnyX0r5yHruCzpYg8Aykj1vimTyOjSUJcMHzozSiW
JT+KpisfSoqXmju5sJC27eqCkP642e4LIVEooHbIpi5WxCSccGMg+k/x6qVXV+jXTLjKx+akkKlP
GO/ARMpucyg+ytKAx+aKUuZvw1XsWQuYkgq+lcUPsEy3n4FVRiSJzY2VC4zp/Ds7JbCcmZYXFuBw
y7E4nKmhHGAGxGMnkmoazP+v+pgOXLzwEWsqpRlHuQxpIJ8HF5pSjUxxpvQcBGdyu+KODViIOcUI
QgSTxjsxWAkXqZFLbbkZaaz10rT+riHC+70f5cXqznsgYiC4kfEm8XoTnfTkeXwTCYvrJYmUyQYs
yGOsTUi78hEeZUa4JBKXOX7k0RRrWgOlyT0LcGErNixiAyMapcfJpfG2hTbTQXC3yag8QwhcURkr
bPrsPr+gJ6/TiIOxmwPg61J87H67ivIqHzurMHGikdFLLRoOJ1a4KIPpqpevlmNGXgiwgPJpDR+G
Get+UjIgF5n1Ofgs7Clg2UNMIzL4g5ydVedANNegTc+aROywCW+zScLb+shqI2pNDGAN/Nmr371o
aOBrBJ9RHsSnp17yowLoDL7UzFiIyhDRdLSicOG/7C7GLjjDQV5nxmMA1sf7tHKtCtV+CuXQKIp+
p0mQstZriKyTOT/WwJXYKuqjic9NJCcWv3CpoxWxxACjGse6JR6hchlCzph9yjU/mWLp3ZekwYG8
uCqvje4Ow32ptKvkXdrBgeFDw6pyc2RU/zkf0I5MJR76Sr0bHDGVTGqMBicqkJizIkSnc8WHIqzI
QdeKflOCfQbDxc+TrBICg7wz+EhFPl5dXKJx4GDOW6zoobD+I7UkxM3sJ/vsVSDAk7E1BCDE4qQ+
mYS5Mzgb2Q3AGn4djaQU3fRnXZzXelmBtZabz5jtahL/BXqgt8tGfhS14ggwnupFuvqzRChbhoLb
sktvx/iravTg16iLzv5lvqTz4+gh2mwjZUgsSZX12LILcB2D0/Ex0ui4qRgLuqPyZw7/KUka/XWO
uRSFFw9+hxyyvppDr+mC1Y02Ek4EO431O6yHeAlWuJThchAC03eQMNL564+exiHFl+cUgsy057MI
z/85O30COasiaVkkvEFI2v9aLvO1K8vOLWDAXAqk/aEY0UC7f7XW3VG5WdDMXsqsH79zb0Ox7i2d
9UaGNjNtlIS1brlkfAFnoGOJvXUYzrQat5KQtG7BGJKt1tHqd7nEqDsbyaw8ofQmsie3q2t+OvKT
rdZMrmMRSK3QPlbZPsnwqfeSGYV7v6G+gKR/AXykxX98D5Wh9kl9RvA1ya2ubn4gxdZwRLQCCqDN
y/AI10m10ZgLzN4hxpNzeEnGH/VdkRd+G961Bwxo0p0h9zOHCaTSgZRJZDjLBLQIiXlmqgpYFoxC
gZoM6+qVYHwt74jg0kP7ji6GJD6G0dX5xEaZx7hgBcF9+g+FLPH8uxp2j3IDMeAYjObg3sNLJ2DY
gtqkmWbB8wh2Rem4j1ncw3k2ZtP6WENtyQ2e+GlqKPyF5drTMA4uxD7BDMZcClAHbKaV0M1Kwl07
HV4qq67+iLX2kt69Q92R4jVTQq4oAAphpZ7up/xIx0oyhr9D0CnVDeYJBAmZ01W95Tr2oGNIlieg
HlNr1PoD9uFjonrGiSf+BIao2NewuCx1ZTovCCkAmICeb0mBa7XWyXNP3IQvbXjRftvIr0NFKbUK
iY8PKPDekT3aNRYpWm7eZz0o0tnzpDB6LnkN9Xldu87HF0M1tkdV3D4n43baN7CZtBYOo5GjkF2Q
DIOEIoAKGXTOZdqvHYf+Xt90pY+CMVWjcoMkrp7iSopG/esfyyvEhkMjWD97/E1DSe1c+ayBSfBg
0wk3wK7+qMNODsta0SlC736Ys/41Lyv+Mb4GSTh5LJFQcClnzfyDJXUyx0yZ5BIGMROTFhrj2g2a
69tAsXvgVAsaQrAeEgW7Lv9Vc4OOhKyp999jAULwWcWJ2bIKNfUQb5UZ3HbLRoqxsM0LGnXI5lxr
S1oUiVpwxIAn74cbhNVPqyy+j65JymGiBtmuvj9/IwydSWnyds5jCFSYF90CzhJPAltsZmEfgvEp
hU4jMy8WMeyZF3xD4vhhTEUtJPS/g1mAOzGBSOZCnRAiP1Mcq2hb1/vuiIPaW3Z5EMrAgdKmQQII
NClBuM5/MRXqmO29LTbxOIp2jFpwCkiLUUG3l/vnqI1hA2kfx6KkpMNs2SMLHfajrZPMYBQgkMIN
r6yYFBJysbnvzYsOb3qlxaH7ZaEdzrOicQA5CyqtWaLfOkf+GmpPglKqC4g8MMl3fDOhtuhXPucT
BcDTFYvthrR6T1b/DcuskZAKDRvcsSeGaMNff4gHdROQ6AtKaZWCWBR9iIKE3o1GkcWXFs5HCQFA
ScSWDVvW+3skz/Vi7+pgcCg4VYjjavOSzHDd4yVoom6iy6loLpcUR7VmPsQxhuI0DY/B5hHE/qJy
eVbmYth7ZFpJMKGnqNRpyrlhM1Xs21zYOzD0X0S6gGgDsolK00loMKa8nvuXWyLd9jwyg2fXYdp7
i+JxqQgsLXlJEkD4rgWZ/eA6isvWlrh4axF/Bxh6CHkydmRDH3pEKZhXnUguFwbWXTvuWH++KelU
D+1PoSj3vf0tzGMvAU5M/XO4S7SISUXGIBpVdTPh2EfQvXtSLYjoI6TFUSxPXz+snkqyPRRkZgNr
gOlHzAnx2l4mfek/6U84D/lGb1ewddvQ7Wp3dFgnDDv3rsHZM4MAkgf1ozzNE/PIKDi57TpOstn/
+Q7YCbASMuUm02yXnx+V0GPxYWHaYob3MNvUeGA/gwtdhdW+o8lb2vSbs3wtf44jK3m5Sp0zT4mz
hOvlXlp3JlKqwW9V14voIjRA542WUNd2ZJ91xzd6r77+v00prZkRX/yKB0NTEgDxV13FkWHn70WO
IULFwsDnzBMbzcSQ8K8pt/WwrXOnwOBSQgLi8Kjz9d3BIHoCg5vnUPsVUJ66kjNpHLLgYoadWZTk
nX5gpB4Ts6xrHU72jppumEJqpMlVyhTVBnURO+1WMbDIIU9YNd9TpsOB5IHtVMnmXBAR32rpu2jI
AnmEUOXIfMcnObwqpq5t7yucTuHG3msD5EhQu7wEUNm3b/G5dkNg/aGfTzDZO2ScPdU9Wq5IcH8e
aUmgjSibsmAgBTfjRTetOvZ0EhGuvXAB+aVWu+sw7pzUlUNnQb6745v45h315Azg1UVyh/2rMeJA
FygtAYqsdoQ+zVLE06KGSPijwgfP4y+XLdckPBAJwXUi+mQ74QF30cyxoMxcvsNt3xNBuMF1PiS0
uWdefi2xcX8khPWxlPit4u/jkp79IkyVFj+p5074L9E3qeZg3Y8OssACCbfnkfsTJm0Ds8idZzCV
AOgHIvGVEHa4zMrV5DIU8jk9GbjPZaYfcAD3WiNCLrxnYKlUZ6YMFphFZgNLTJqnsFqSN+o0qQRY
k94FzxdpO54W7NZ5cL8OZVgCFTG4iv5vBxlSy+0UTQzndCzrulld5GghQ4PU2b3hlnrgrbgcYmu3
fX0OEi3b4YFk+sY1bscQp0rZ8XyKttvFgr6TvKkM2vrFIydWT/Jm5wtDY06oCd3JPiAlvYkyJ8JI
dmIPFw6P05bZItPXiYvOK413JSESiQFPRE26nU0v7cJlxDF3ymjz1Vyd23n8NGnqvBTb7Qlw9k/K
iPeLtQHx980gKzew02zVC7/SSKEm4Db8glB54Uwv817y5ZrsVc2WphfR++QlMBwvNa0UEbiLFwgE
zauGSTOEUmUqHcaajcguLIjuxeTk5KkECmhXCYx8o6DUdwxzomf8Xp19RRKWQHgX7tb8CuVD8Pub
4ZPB+kNYY3x3yvDChSbw5B/D3/Jc/eTvWG8+EwLgSMNNH8MVjzlj6HuH595Z3wO2pES1DeWEuQNm
NLExfNCOGoCyOhAr42I+o1/AxgkSFaRtUk+osHjJuPgc2N0CSFbRYZaR2xEFfbiyVceWa2b5/pCu
spVW8zKr5d5bOx2MCVPieLfhGfI8Dnw7oh9Icj3btbQyq1IL1MI7i8SEBNTdZ48pu5c8i4DMXg2E
MSX+yhHB3maT/0jYFTfAi9KbkQp59hmC8hRrzoXBKLly9gD7pKBHIIC1NV5W+4ill12pmhayfXEP
a+XNZqc/jx2XsTA0pKyeLxZOE0Yk7OVdzK3+bYu0t4fxS0rp0OgmfAAo2pG5OZ6lhIStSHo/Zgjj
6eB/GqTogC6m+lsHRAlnMzGKiKMO/apXQPJwmljNNm2/w3muUq9wjLoFCFA4tD0l7PBzPM05TSrP
DKJlMLkLKVFsGpZhO4Pl0o765AaqBHpVYKEDgRb5niiYjEMNSN79g3tMrUkrCFAF2jXQG7pYaaCP
eZQyshCwzM+GLP6yjRc1eeOjE37psGycX+kwF2ncYDXABoNXZdw7LGfgeahfYVNUclRm1aYEf6pT
Z9qJAJUbXHWtjQ4TcXX9DyqxwiACn8y7wMVkT0kOE0qnhvMGVVQH/kDMRoFWtWGhZKfoYZJKu6Oa
tlyQ5pZ+F2MXgDzjRjDsKDD8nxdsZjSEsBxT6HYTAHMo10LEwqHP4bKx0ZLJ2Z2FtfFuhY3Kbxt8
try5mR/UiHHu3UYLc8pWOFVZmwexxeu/O1EpWUJmzdedj/RggwYAepZTZie8/aXS6zoiQhWZWGGx
ou3tES2B/1xkiNEhkD3ssLeZU107H8q+xwD/xUkPMMKT0NmElODJ1m434wXtb+MJjyJkneNKbfUa
E1yjHKbimoWmL0I+I4y54An2S7FpV3KWpieC2BHpr91GIaYXLKKW4HTPX8X4ePeNilpy4oFvPSeR
iCCTEUwJiOlhtVvAsK+IRWt6oM5ZGWpUOw7dfBvrH2fLgTvh+Vk8ztdQlBDsBM24bwlfMimSjvf2
2p9OlqLJueSjh7eT4q/1LQbO2mcHCiBy//we/Z7AF0QH/vaKq7zv+giNdJdZqMF5lLEaINbig6+/
eNvj1iRBCtvb4qyzKxRAPZjzl9bW08n3p/8oWBCPhT01OgfZU7Izapkie/e1IYFBjZ1gGgOAkxc+
lzrzLsQkiHRsB5v5Ir2EsEKGsGMN15dJyFeHcmXJl97gcdYzW5IH4P9w7wE0LRX/eLMYxWJcI57M
5pnB/w1lsdUc+W40aVoFPQm3gGwxxwU50xfTjxidIRL2yCuo0j0yKJFSSlpj1u/jgwX0RKwShabi
LeutRy1oJF377+oyPJ7E5PNN8ekkkUHdEvR4cQWGOrKtisGKAXpaF4z/HCInQ6E+NNQmvaPC2yqG
LNS41nXCAIOwVazhLCRhEoKozThJ+c6+/+geMNW2WwdSgEPK8p6YQ9OT9Vh9CdpsDnOEDdHcxs0A
reCoOSLAsqhpkGCJPfLpaksuGzqSH1rjIAuGRPAWFRdHsb6eK8MwJ8Gaj+DXOAIK864k/7stPDPM
5RtBdo/R+ZdKewTSe+OwPKE55pT9jbzgvaHDJx0ectMIhChXuCljGiV5nH7qyoEITUMS/i7Pt1Dh
ABY3OkIFc9tZ/UrmHiABwrPyAw2dA560haMk7euc2+qnVTzfSSA7+K5v6Kq1Tu2ybdKlJXFBsWzd
bFDgQhAS2VUEEvIO0S94Ee62wFZNaGWmTC+O+7+RenMk+TZNkKuUpzpNoQ7c54AOupfYg5bSLUOP
yZOydYcOtmBGsJugUp74EIOzVgOlM1Y3L+EkjNzAJEuqWUIHgv2Yl2B0npNFIffBJNxPCr/7pDRO
g6z4lgHtqor7x1/EU7whLqMXzpjNrBiM+/4MtkJBzqzBRLHrPwGfzf7cZEl3Q1R7gKhhsYUfswZh
PeaXw9VxQp37hp5SGVzBULBM0w7fVVbrQ0BNmJx1DIPlBZKNnphCfkiRRnixEboXpG/wnI3o9zeY
z7/x7qLvPJlYGZV2xKNTN79yMhhxfyqe/WFlwRecualnmPoCIplokv26j6xeIpEwYZkGV1+Mv3gW
aybnkP1MBuC8SbcNaVhuXq05BZAMPa1xRMj5Xokho0t8tnE0Y3hDHFixo/XS5PORf+b7IYf6P1pi
RMaOtexjBBiDi+IwEFHuyIpotPet2+CXtgYIiLoHfkOVr9x4jfSai/xek4wzQva5PCSQsDNFIC8o
n3rrYdAnchZ1dK0TJc9SNzz/cm8eygx5yfCnN6JZQ7hFwiLOmH53Yu0FlgIw2W6XFi2OZleyFVr9
Wa9dMa7xF2hJCoO3tWKCFTXC2oSWtG2LXDJzqUP2XxikBTrV254ivW6gfr8hmFtHRf6aTAlHU6WK
H8guYigZbmKgMoVTrXExx4lQ0S65cz7+C6TR0tE7+6Eb/GX7O1jCDBAWpbjwnHBMqcNLvxo0+i5W
XPjeJNfgp0i5udk5xmQM8ciKXN3NZT3BpZ/2e/o1l702CeIzB9gz6iUwxHzL7njAWI4i3CspCYoS
7pskxVSL0QwANIaI9sy62Oqp5ITh4qMTj+XNo82V8XB8FKjMlPamhKb7Lz279qn+QzWIHPZ/P/jG
u09MPtBQS3tVQaAOyAQywIn1Kr5fEm6IWmAlp/tYThDIvp/aaULLrcbiGl36o9iWKAwSpb0niywm
c0tABiPu6rQcESD6yeO4muQ83LwSBwkhLQ1rudyeSyOrMYzIRJAb4tmyZ/aUFAqcMxgsh1q2Nw3I
ILCE9Gsr7TqQrMwRIcPYoLTY0Y3rlhC4O14EUu/4aPkgXEKXhpoZewzDdb2NFvh71So77XpA4/Tc
SCtRhQciKT5WTEmHosIuwX83v156UOkUt8L3/bIFL+uq8nZLxYMBElJHFfW7c41mPRAI5QBgOsEr
A1GqqA9WufEcD7YVNfyMMtiI5MAPTERMuMRKJCFO+ZgU/tNFNV700mClhqYXfkAk8rM+oVUsO5WO
wQD0Sdk5J7YVBh8B/zf04i2mHpijZFvfe/a82aQDKGum/fayj0bfBjs1dUzTz7j9D5RbNcbeNjKd
oYFZP1XpBpH8pKslfVVGUwqQIwaCsDXQp/w77sHzpGNTyBLHly/WvWceWhhjhb4eCXvSG4ItwYS0
LjwNBo/uvl1D22Nu4jx7Y28l8pbTkrYYpdWj1MHPXtWxEuz1UFbGmkWwhZebVPy3dInvSZh4R9Wg
vrY9LSX2UGd5nzzbYl5+xoaFBAmsWpwZJ1Gs1ZFCn8ou1T4WDQp3YqokP86Sakknkx97a+Rvak1l
wU2RUAjN1t3AloXxtM0LG3qwsVw89BW95etL/mpMkH2eAnGkWJcQyeH1/dXi8lqFxIkr9s2cPV6W
/SOsTPP7a+9sqM4WCEpEUY1DRC9Mw7fsoLeZw5mEo/J1T2sr4f27XApS+uiZ7TBxwyXxbpQ8/TyK
Wi/zD03makSlEy0jyJeVdu4CYdzuBG9SCHCvlJKKVQXNHonxCPmzEqVkEUQkayEXo/ELP5Ibortd
1bXhr3HtpOrjoE8QbccSIsyyby0FEZDjQjV8BGjb5fssNOYTRevsNu1C9umAG1X2+KMz3yLcJA5W
9UCJgEPz7gIPk+yabMs8Eyt5KKQrJy83pXFDvCVQO0IS2wsJXn55wYVUmuSdOcorZGAUIJ3U27gx
GacE5TFNd07TT1I3jAMQ1aI0Lj5cLvPwvLTG6rXR/wFg74XsxpJTNIlO8PrEfUbYeDxK/Ax1IxW0
n1CwYYE5mpnG0WLSQMhYHKUrIMowh0vk9kFZbM4/g0n8/jRX+BkStVJxtl20URYri/JhM7GWQLsv
omg6v55U8trpoknnjFGCRRLFcTgd8vV27y/ltjBWcN6dOLKWnakLZk/PM9q9qbG1iBr++g+O/Q6D
5TKNPc9Fm7u/OX1oYci+KfOsXK2x3zNrTNtA5HaKF/UHoAPm1VLp4PsAMpAu8M/uCe8/3E7F26dl
UNUNLCC2rAawdh9TUF38d0UzD3gX05gVg1D6glhYu4lGFed+Ljuj3HfZdruwPXgDtIHH/0X+L5VJ
SS5KoMEzjeuNXHvgcGmrlGb94TKh0XxQsdLi1uHQ3WfdX/UxGzWdNPQvva49Dj1ladsuXJ0RRbuG
CABh+/S9VklEODc7yafIYf5cQcjO69VKKjsB284RkB5+eU7GepvZmddyQCNF8QxSP1FWayjdIjzr
uzqsJO/x6ZihwnNlQWE3Zjb5iGNwc+R6y2lr4jc2N/SY4vpr4/xErfTwUutlVbwqW1N97v77rmAJ
Ro1fbT/DklPA+BHO5yxOmYYHmgtZUj+6+4S0ccWzveYJcFginPJJu5pkx710D/8/3IX7tzKceRVE
xy1gQqo0rm7A7+6HtvW2ELzITNoU8DpHU6A1Kv8PrAjqwTyMPzlxDYhgeUzeCFIuadbAn4i1LTRX
8kddwPqJdcjJKXA+Zy1NQRMWobrdf5KEcOyvugtssTcKSERnYAGsbndRBiqNjhykD4Abs1ksGJ9l
rz5Y3mDa6hPPTk0Fs0sI5E3urrSxWJ+gbOAKjjxHw+dC/hV+69sppJR/MOPWKXuoXgYh2EalwbGN
FJpmabcFZxiq5Pp97vnzSyJRtqOiwXtRpG/yecb7cjV4HXo7OitFT9WLptq+aUHocQGx6Mvc2/7h
XedUGfuKJrp+71IWdXV09bLEJeN8+Y5xP9wARuuxRL8i1ckSPZHr2UxD4iUZJOgJ/aCoOuBMsq8l
9+U2ffE5idF5ZTmvymLyS26tn7N2+vYaisLmif+QtkO4mu6LuQloeNVfFspE1RjDT02kFNvQusmf
Fr38udQpTav+Br5ecBlywzSz3O5LJTlgNAGSMMOfV/vwOJTCqQOZg5ysNW/OAVC2Ddr0HGK08VUP
mg61HMMzYzP6+MTl0O+OL7mNARpNmYMe7rGkrfnZQlWzaz94wMiNcO4agOvnZNrsZbJlh0jcrgZE
7k7rb52Vu2eW/YKl1n9TTpsGS4Y5mj1RwfgWEAS923HFHcPZeF0jApTaD8gec2uJyel8gCs6FXtL
cOvvUSC0VTw6CpuYdh/U+TVSLxjtcKheeOzDx5yggC63heD3nB+d1I0vrjIYjVk777YiGVlD/PAv
FAc7934+l2nLmqmWO6dxNPq/HYcSfYEiOA4YBxB4Xs9GiBS48zHLSqCsCeF8kR9J+xY0WQ/7Uu9y
teLNgQAHSz/aCmteDFprNPmHhZ+NGXBGShChHrMMh8hnEWPqBwuRGYnSXm+9lpkXNHSzZ6qFlFD8
v8/7a5taMlZX7nEhr+j+Kgh4IKYmfJY/mFpHZI98+QwmLwsSFY3eSEXO10YPZqGZvDAR/ZRPvOM2
6BQi2ZFDGtzJBwEGXBaJ0u/jAJHTvH9YPQNlLApUt8O6mS8mSf598EdFapjDjqI8h07sU2rr1bMA
tTrekMY7xvdIAW3rcPL7rPmSTQzcswE79Jorhk0IdStEcRsNt+OQoNs/Kb+zpPG5f/ptE3AxqdKb
277A7josYRSLKOZISnXXGFzxpgMNVghFW+DJQtaKzMIZZWZ6VWAMfYwtRlH8ii/o0c/k0TQoD8I6
bI/MDlUYmCeB+duCpHvpZ0ijHa6RWAc40sYIFn+T2ik6AeF38BLisyZ3tXcuZ6rn5leIegC11HHk
H+cBl+1PTm3Sy5hWZz0a34oEpVzT5zbaLYvGXTJXXUU2DmufuLFwi7PUCukDyOfkZ/pa6BRP+qJ4
EZZn2/RXwAMExzFhNamYNLk4b34TaxLkbj+16ajIDWdzOFiQrLVwi3AxKapxXdbTYxMQgVErrvy2
1jb0evxJpXAaiLKwureo6Z8sRX6VGe4xTam9bIm3nSklz2zQeoErW6G+i4/Zikrv1yRfJ/8Rr04M
n4X/fw8G2nodRSnqmWBfT7TLYOI3gkJmnhgqis9YhBFYaphiNJ5cZkTSebcVPhSxI/QnPl2OCI+X
e9ZoKJfnNdpKMTJ+WCUUr/wUTy6ELqWwn1bpE52jwzoxAg5cC6riVm1lX3j/bDYcUzK1jWWMMX3J
UE5mXf11bd+qH/mCShTRfeVMkg57MdEzwnsGH8G3XRUc/F+Vkm9Y/34T5cPQZF/INyL4WxQcOe5l
vhYX6S2515wwH3pzIKmZIbkwEr4lygbeGjEX3vw7aYZQ4S1cj1W2TuJxxxasoXBoWHtSTYD1tU/i
75oiTWWsok8EtBqzovj3PTBfxAOiO3Uda4dqv6prqmxUnZHW9DPlfSmARsrL7AVaQ2/wWwO5V4mK
adIaCT2Ut/2M4UTJa0KZPXR0eUGDDwEgnOcYNYnRT1LOaAtTInQPYlQYFmEETNnRqqggAmy+8BWL
U+9cVtO7+nhoP11sQFJlgDGgERA5nruifpKsiwfQQR/nj7kB0dDiPMabRbvThqwv71yX/GZHSxRm
KTWid9fj+IWe2lxjA3cXKMSnzmPnVIdbnGswGzUYfYDrD6ejQ4rMBY+5G41h9gTIZdWSxyQidZLq
xMGxX3dWtUrtCtF4Mfnd8+f8z4uECIR5DKT1fUU6L+4grsXD3ed8paZQroEtrkrtUpbAHxhlTV6B
kIA+N6+jbvUB+Mqgm1r8jb93qfVWODmXBZwAvaQ1bEu2C4GH+mSFuJcCugSSy4kpCXBwEHqUqXUK
J7ATtYmIX9yp6mld+GMmrkNUcpyzB7wxn7GgsszpWvrVf0gOyiG5VjB2BBY6LKpFXdw6jcmJYM7/
g/JgfdePs2gAXDnKTIaW+9b9Y2BTinGoJOCjVPcsUKDRFEj4W6WHhMrgPGZgrLiDmiSVzLeDXDuw
rFGNH87dHPLEVOTvd0SEKHuZsVBlmGH8Ygy2zG+lPFLSI+Q4yWS7bXmG8EWzcdlXqvyzxchAwK+q
x2easS5bhFdxmgR+o5j5WSDgikedy5aDQIWngo4LAB95HdPy4d9bGP6WgSk9jVVakhSjXekWa8SR
voPBs8OP4J+6H3ekNMuTxYgW8yDGwg8NDGSz+8aIMbXvzxJ0wVHtGAqQLV831Oy2ucLmTyC8oEaK
LZ+/d7AmCEbtFtyH92h0YJC6rJbqDAcn9kJhB4hQ+R2vBhgIiBjmU1r9Q9a/9PhgCI2MsgsdsJI7
aDvvl4pl9Vmx4XIrjx7NDiuQS58Aod9vzbJZJHza2XURDnC9DCMmsA+Wj6qQTWa24AYFtGJtEXlK
0YC14nPBxh0BQG8pOMoir2elFNREvMPVems47iY0vYcAIVT/TpQho7NyRKi3RnppF5zV/JJBY14Z
cane4CapZyf1ZJuCWpDm1dhNxshp9dInCP3awpVtAM59j6dymFTz4kFkKTNTj9xry1gL6XSHqhod
B0Q4w0WrF+YWZRJobDINSYMpv8Qc9ayrAHsFpxK30/+HnQLuWGnaq9dpJacIXMq11F24apUOXng/
o5y4uh5MqXgKbNjXtdBNoEzCnXEaGtp5Knz9TUgTsbhDFWdEjadL/k+v0xk1nhL7S+igIDCnkA+a
w/cXoh9gvrhM2q6yzxDk7qviZMshP/rjVgTT4KK4G4WjWeer2fMhVdRMJMDk6VJwtrfotLZaIJTb
fa96ULJBIQ2bpsdGQ0ueEzlC16Y29v0b938YtzpUDpVmsc6FD0QwUE3qvfevFaqY6jz734R6r8i5
L6ZESDYTUWpsFvb6rcd2Slt2PflU9qy23CZoLK4X6nK3zFjXXqHVDvA7jZ+re85ezvNhu6Iy7nu1
9It6q060QfGE1PRgjUHMboBZCVQzGqSt0ybxAyIAwGiSGI8UCHRMpO4EDpDjBlwstZ5IkaxNliTQ
kP7f/xCTO4QiAUEuzwJDr0Tv0MKsxzTMgzJMXvC8hEgrrCaMhcBe8aQWC17fFrcK0K8FpF78725A
VCujHmvHPh2Y8Olxval7iH/pV5w1m0hqKPvb6Th+ALECIdCK8Jt3+DwoKineDNN2yU/EALeN3U8y
wls/hOiWH+bKdVfzpdYbzxmQPiA09wAo/PRPKUTqVCkWNKob1lBpNgeMLGPWcF+aJxk0DCSUVy46
gb95Mq6TO5/2ieZVQyS1XvDKfRvYxZwR8q1idM8IyHUu3dzbvk26iXPYFbY3vDl3T87SCwM9q15G
hpVCWaoXYkLcPOMoFFSBn1BO3DSB98kUkCV5p3FOZMCdDNIIgaCyOBb1gkCtL/jtc9e3TiW9PEdK
Jhaf/pm3fIyPa2ZG3EpZuPH4PGmKZHTrZCV3V8kRU14+NT4oO11LaXtWY2JcnxT9QunBpRm1XMVi
J5OyfY8nG3pGW521TQxyqo0qgQ+txaSMWqsx4WTzW0AzJA0gK9PBsVl0wAuTvtRfugtMlFKP92la
KmRY5u6ACWLIm49/6Owm04s65ThmQNxfT9RNsl/kLsvELEj/jWRQ4M6OP6zrVsV4NbMtKttxBgdz
5E0ruVSk5KDIoZU3XeHfnB5jvKDUv/lOXw1rg1oOMgu7NOnhxvjolEkJ9GbmlQBzFJ8O0JWaU31h
GWTWs8b4O3O9NRRVOZWac1Ns1lW83Arr3AsIbUOceFIfACevLPX7TfRYQMTywOaj2r3WvUy0fQ70
ARtbcz5quQZJcFr8O3P3xfMz0OhSyK2jmqEufcJb3bcs9EZfMccx4y2Lm16Y7H1vRG9zJnv6VNqs
kqvbJ4R15C7Y3OTeuejoTNc7NCrrIOzanCZmuihueMcacMbHFetQvZ0+eEghuDKMzQIkMEoogCGZ
LN8i78c8/cTbf6K5KgvA3s3u+75hPbzlLetQcqzMH/XBiQvWL70sDlZajuxtmAJPa3ld0+kQkvvL
QSZNGMbDsTS3/J+OnkanJFPTu75/OlqDh1mWxfDbxfP68zOcDGGB8H7xUnZTabcHxSHzjgNP/z3s
VsZ2hZNx3H33ELL+58U3NOs6gWNCTv99ww4jQ26pRAo364+WOz4vh06zAydQrvzPTf8pJlZvNhdF
XqFfbRRZbZF7Mp+Aq2AF8ChkKqHVvs3rnnnaIWU4rrmGZakYWwEdwk8BJWVDPbjrYjn2y41ppD3J
ClJouB21KRwCSMNmTE5etVBlcXTdnipZtILxhMH8muisdBejeNz81pxfyMB1brUn5pHg/PtvzJRf
UxJ5LLT3axzQ7YpRBsjqI8OIaWkO/L2L3+y2WVG1p1ShUUuYIkuYTDnEPSDYky0FioBxdhcZZ91q
nOz+tZUbsNoha8WcbR0GzqpWjmwSKlCMiRciZcGnaybriW//t1dmN1GLfhqohH2SzIWUwMShWXaV
yHCoRRhrgWHicHkqcKvOtx9FOp7P/tRTpmFElxtS24O352Np7oH0lkS3WA52LEMxCvX7qRn30eJs
jF3BRCNUwMexikYzhBW17ibalaw3RXAGsgKUc5jdLw5Nk4K9Y3JGv7u42qsDWy8GuWSWuaL2vYOC
FeBNCmA7em/MWliiuP7+GwqREowuUX3MrscCNRHr0xl85XRtORz+4WObJjxuz8cdwVkOm+DmsV5f
EgU2+/H+QhZ3flnjJP4aP80I1AWYcbWlfFr3SJwqVTTe9YUoswFOi7RCt30eEsuVF3D4UrCr5hQ9
4ruG1FztKGsrgqywNHLDqioGYyEls/JcAuKd2wyWKvjkkiYX3uy7wovB4b78L43OgMt0YvLEjmyx
kCyu3yJQDBDwTVdhQPpjxM87GxSgw/RSJuSx+dfqYJlUSiBb93Y9BQQJisLruVU49vwfnf9epW+X
6EzNG7r14aUaJHvsz1mDnwYlszGPwXnwiJtl7sO58noqWp4H/JyiJvrvvWCFE9UWIhtXpcObIfD6
VefhMNYw12Bn/fbp89pjlbHewQ/L93SAX7mBMe0SLdpq0x4f4ONp+CODiMMi2lQ6yJ6OuxwmnZ5K
SQ1lzlsy3i+lxJcESNpsZZzgN4iVmqdA6Zj779jKLHoWzzD3i1pkQ4BSMY2GLzrkRo9pJ1TdddFj
Vua0rTaGBNxIDZz4KigR//Ymv5PIxnKnkhtGT87STdWZRNTL4cYIpFYZ7tUAi1D+InDJNdKmGCHK
NKrU+Kj2DfJQFAUNX9PZiyEsELEwV2KIIDWCttl3iJnQWob2kUIIrdSZ6jKvlFew7Eob+z12jI8y
478gKnpD7w/ccvTJG2y7UbEQ4RYv4aZO0Imd8N00ltoNOnmIEDhiSJRRQEUsm39UiizDI1xAp4u2
AYj3CAZEdy8rH1/+QbMRcdwvcowjorHGXYgB6MyHGyjYP/ZDsuQbu7H17lAZjmaWUMkF2KK/lgCB
VZ8DLf2xSoW7ErLC8BwLnmoWRfdaN0MTQH0BSH1bz+VJeqRKV5COetUMGbajq6WLsCiQ7Jlfob3A
l8kmJkeadOCT2jrYvqPA2KAYBRN9WoVQs0WNqhjCYu84Cg0omUhwUpOVsRiZFzHDIoTxadECdAsh
Np7oIPxTupvFQueQMBcguA67v8TgcjcsNHRcHBGnxxq7JqrXumK+0+nwat++LpjA/3T8F+8C2TN5
UsVV+sksx28JUEy4bAI3OjFrLX5NVLHqCYORElNf4rs99XYIvlT2APWKW/sqpckrJz9g8qV0FkKn
+oLCHaN3SOiBv1yOlFmdPUiRaCwqy10iyW9Jdddd+ueSi+QHbh6yYnRfs/YfsulATr54+pxTNSK+
HX3tvkAKrnLISbXQ1UO2738pV3VlXpKqhJzID7e+/Hy+pfjqpjOKoghLS21N/nYqZWEXsW3O39r6
/rp2e1dDNGMcfXwSjAhjwOMz4IcS3Y91vLLqCdKvwlaJY6rbm9ySbBEDOXIKS5cThfslfBiVNnPc
agRtQMQJPm2NRYx3HBWUfxXBq0hWB1GOZW4XjnHULJg0jVX502/YCHTU9NR3jVWLnLuHOVQHVNTT
qCW8hrCI4jeeQJb2u+sIJTlLI1ExXZLgrp7VNa77CTBoMAprFxFl8Dkc+aQ1QG7KJoOXAnf1UgnH
Nw7Hu7NS/w4zY8BWFDxMrac6tagK+nySFwx1y+Oy9r5cA9Vas+KwdMpB2jRgA8BJGSYmnhpyWGId
QUIqVhiQeNb9GEGpXKnvBxBAPRn6PjFbU17kue/VeJkjyTpkw4lPT2iRDb3NFZWfqWHvBdQFV6wt
y9Vm24iQC/0P9iF/bsFjfouP04JvNt+IvhmYOkMGFSKJrUW/C/Ac5TrXP5owWdNBqDYO5MmzsflD
OOY3hMHJYF3JbmjgjwlCzZbri7pozCHVmO3aG2XC5QaMW9vx/Ln6wqh2tXNm/Ir04nzd3LY0vG08
TptgAIoBCRj5tEhteiWOAwdr+nTsXdbu/9sTLzSByHgVr473LnTtzFCsBJcBnbKOxzhfR+EWGx4F
ZjogQquEhVSzZ/dYFmWzMr/EkRjCrfkvcYjUIk466muZnjrTTzgTq5mIV/uMtQt/5kjLd9QHJViL
RYGV4Sq1XHOQrNvVqdgxcSFs5av0nI1qXfXJlwnZESMN9nD2pY9NdNNTtincJmmlGXLHvo0EXglZ
p3IBDUOXYJz7+E/HF92bBEN4FwVKDkqMGPKyrNS6b6jCUVAd2lD67eyic1On0lTWkHilW5KimbTg
rN4uS5nHwmN0f7LfMiYBq1RbYmjOwc2GvcKq1qAIMbN3BvKkKDBLopxLUILviB9Gx4Sp3gTYHOnS
yEUsZ1zxt/H/j7iuOdeB2maqelTWkKD8nvW5Z3B2CmQ/Si9WPl2EQT71hZ46KG8H82Sxk5nmmpbF
9w768SaMW4VV2Za7YYYJYSh3hVJsuEVva58Acy/wH7Xa3MyzBzvRw6aCNGxIeM2ccK6BtK3AsNvv
7sNz1A3rcg9omCnVf3wmUdHAzwXOA729GveGqfl6zeJ/cA+BaYsMSXQyAJaRmiIYJZyrtiE1FRUp
yLcWkduaKGZmhO83Qxxv7o9TndCyKqR58qMaxWFziEp0cHD8ewMN2JMWe0fcjP0OYY87MMMgnbZC
3L079gdyF5iEK1MaahT85c84oxNQdapTpTQaBXnHiivl1gixps8Yn/qXteyY+9DvxcfpvpRTBwO3
2Af5Y0tXKv5oLTBS9RtgQ8bqqduoKhKcmNGadCpweg5v0a5rap7Iss13userXVIc1xLF4fJugJx1
mp+2CvBVW58u1nfa7BgiJ0U2SpZiB4LPcJNZcaDYpGOc7Eeo3W691fN3q7SYbjTXJDvd9lGamniW
TRuAzs6BQTJZaY/OD0nVZYQ45+MKFaSqPa16iFbfOwErC3j7rgAH36oYpwnWmzYI+jJSH8npewBw
R5yHCOHs1miNeOErO/bPxi32RRGvfOWlByK9nYgZZTLnTEubArXS+TFoVdbXRQRD65lysjK3l5XV
lkzHGN/UUxG5LF+nTTub8S7xiGIbKLhe4+KmE3CtlYinVfZv/oE/F3HSSuinAmPx7u3U+NTk353v
8++ma6Q8tY++XAWc4wTGv5a3LhHV+bnTJpjcr2azhjXPOlo8+MAeLg1K8P6G4UFrBCmOhPrcamq5
h8S7x+p1OnBAj+4s9x8reI7e3K5KEbHwRWh68CK8cMAm2ro2lERXSFD9kaA2GU5R4aBXgZrtOOv/
9DaG/zbzcBFUXRQ6nmwrZlUkSYcDkf+oiBIjvyte62nEZxtkq1O6e8tuaETnQcpDurKOMF/sWeW1
hOnVvscQoQuuRNE/731Sh4S40ounduqy5An59zDweA1BkyvrXIF+YSSU9A+vpEyVEK82pyV2OEoA
ZN/YwN9uuW1UBPRZZpJ4kb5Gcp19coJvbzO0JFmq45nVriW8K9gy3bOK5C3bDQT0rtpQfTICTegE
DoSvs7cMZd0KSVkxwRPNrIVJOJZipLPS2tXEzGs/rdFenmvU9ruGxd233kGNlO40yu2wVUd8IXyU
fcNby61huDv9aOsrHqUfZcjjzAj23SPsp/yQ4zihta13K9dD1Cyh1YxdapnsR4I1dOdp4g8FtUMf
TWP5A8hbuVGMzOqLy/CYfGVOzfNX31S3BMci8Rhp6MGtvIxyBSX0o+MHQSkDNfr/ad0JnZceNOLw
k6ltWMoRFjwV/YVXZYqQQaWQwspnQfVLKrTJeTREEy60mGEyDQ4WbrIp6YGaUf+fAmSszyO7yIHj
CfqFnUw36T+PxptDtFfzlWgY+cQJtA+zUJnL5LNECj7IJ7gsiwx1+hoB+BLpJJRJEVDbGkTcssgC
1iMqf4TRPl6JyA+2Zjs4Krth3qxY5T7Gzr57FCGwHbaUwXqS1RoDVIWFIyZr3IaDrnxI7uMZME0L
jgNp8E1uPJQZIThKtx14vIULPJ0e3fxjvfw46+dhE1jX+kTkRBubeU4fcjVFR1c6C1TZ2DbcSqN2
MTVkWC3MCfF8rHj/wYjUWwxry1QN9m0HUzPmL0QwYMN9WZI6ch61IYr0EjB5qnWfDhJUdRxKnFJZ
XL0EPS837a7a73OA0sDsoYF2yZMaWxdKhd3lLcpuTRoz8QTKBUvemfC7gSQbtynEjt7qx3aOVJC7
/Ge8OawwGfZRQ3FKPgLg/44BRLVYQDj+H28u04zW+ZxfA4zBFqdBB90RlSmQp4VnO3DZbPp/PNvf
jugNPiRfiwdJmUc+b1kqAoRa5I4I4uNxbm8up2eqzJ1xX3nO9lfo0OpbuMor7EmUen79jEnP9RL4
OaEvwjKya1ypv3V7lo1+4UvbVxfkrezWD/CBbI+i61tyz6WSPfo9ID2dIEv/7H1PPCtj68omnuv1
Ig34BDOEDNQ8GDPqElt6Ai7Zf51IeyHmUCUMAPiGrG7XbrTao8NehAo7JbGQ4Tu+52ieHPBTZZA/
1UQIqprTyZJonVUTIUNUa3OEMDq8MGzKUzlu2Lbj1cQvNuFxauNgbk6EWG5z3Di06zig37MLpBoi
9+bwXiW1UFr/dmkk/FiaHGpv6FgZt2rodi1HOIBJaUdnKF0zQKH4jH1061W1Z9x7Ovfzv56dS587
SFfcuVUTIpeXJ6MuorB/l1qoi9JKMtQcjECKbpDMIF2kKe45LaVYG5SMnJ9wGjsjDEXSQfBH9Vt7
J+7RI6Nvf1FGD3/J9whFd/Tofrgpf1degdudHTo8yrPum/No90pCKWxf0+dFNBMIIdptjVsC2hYi
7jaPMZywZLRs7ug/eV/Gyl6axQSe3h5MsMOISAPGvnDlBHCX39NtjOx1DCXsrK1/H2+375fq6e/O
Jw5dYr9Fl9Y3fIzgJbmrOchCmg0Nm0sHuf4209ONEoYLKazxcn49wyImTiG5eLQB1RAr7absN4IS
UssZNN4WUAszyOqmWnT9ozKreOKYCHWp6TBlRDVVFcKqvSo273z1fpXVtXdwqYc0xJ48zDiLM7/Z
MKIXrlk207C8vk1sDqq8TLhUk/kR7DeaGF30rQDGDHQ8eh/CXO4uDch0UTSNgRCXLj84D7j4eC7F
Fl7q+VvKxOXTyqqUnPwpmc2aTc0XSHhJjdJMNABgziBWvEd1KJoIWGhajDYM4ynJEThwYou4o/oO
HYRNmk0aks5sxfLwl+zfa1rAE98QZ3b651K7osJRQrSfHkvKAEPCI6kd/Kn5ja1HW9VJBemyRCEY
B8p/xSBDCwVlDjDF1TaV1dzf+vvLsDxofBzvZa1LVZn20H6ro2T00XtuuAjVFhktCtNAkKQLhIUC
/lLwPrrRKlDeDZwA1ei76rmJ+VejOXITZt6RiEWUDDybL/1eEPSrxXLBBsmBJR266TDVa2uu91dL
oBzJuE+0zTOqKhGDnZi3imBlZnKVjo6bCYiQtoZNzpekvkiI8x5pxRWkam2n4pV3xLHQ3r+T3PVw
gbE2A2Rq1+V8bNm+D/7QpzEmmKM7TL/ajZUf5QTuXf3Kg8ET7wC8RjPk8ABs6hBFJNMVnZQkJEH0
nf7MhiBrqCpVpj2FyCePqNboewzhgvDEgYA3njRkvpmNgABBHF378NHbUKncQ91vl1bHmoxtjNSc
+ZaQQawJe6lmqDd5X5HtDiJgqpkT+rxmePSwi+AxioaoJGOKJFBPLUbTSdhWEhp+y/wYoyzBgmvv
vIQmUKckQuvue1UTvX7kD0q9chTawMks9wRTVA6aXCCR40EK0nprhNmDpQmZJiGPkZQ2jFqmVZ5C
EURRyJ4c4yuZc09pjquE6sOGUEkVBf1LGZgTR6YkoEYDtHrZamtJSkuBhUKCrI1jLP055ckSrtUv
5kJbV4DKtUvqRaw+2LEyO4JVhGx0WY0mRnhfIiW7QQuPjgMbyiwvqrgv6Kk1wBDr1jWaDLTJ6C/H
PrcnyhRWne61sIlWZvAQdIumD/Hw8itVyqljysj6bjuIKI06ZcF3Ie5aQ6PQCwX69J2wWLz3X2Uh
60kSGMSmkHgPITsqu7ba0IqN0nu3lQn3j3BpaAYrTHXjOCAUDYfLqCBgcTV5BJFKp5drG7WgMzea
vn0JvIUdnYVElQAEy352wiabKz3lHElc+3JyedqiCM5+n8do3a1I3pc1QL97WEsIk201icDmEg7P
ijafAw1rjqxQ9uh+eebbKbuBSxMuTWx0qFdjksEtLawSgQv1P+NXB/mnyw7y+fSn2eYPhgufYTgc
n2TQz/xlQChgU11dr7eq6hXyaSDWYbjXctDFuht9yURBoOsnc3lVliiRhRUxaB6eEt/3g4DTKRNc
GXGH6yOdHJ4PogS0655aUrDT03jrMyNVaHFdHuchwJ88N9pJBRzFWaCOjs3Tpoet4rRwHjbgmuMH
olqCcoikRXuvGpV+9Uja7ezBihukvTCErShs6oJyEfHqgJ9KH7GlJjO1CDRANi4knibpa1lEXcMe
hvMFHDslDVdNyCnfTCTiap9sIxik4EpBl1I44zYJU2zVJ2QDkxaUAWXDq7/cLq4plsF8t6tOJC+3
RxZT+CChHa2Js+5aemFx+ELtJQ+nGVjsFzNp5HKiYKYs2k9afjjtNIwu1X/hAUPooH46SfR/MHuA
2fzjwZENXzaJ1yebGhsI5vuFy7DQuF2Kx9IpHb5V7YY37/myiSjMUwC0MxefImZwwd8PL4SOCYE9
TYsVqg8lsZY33/zRsqGtzcv+49F1fZZY8VA0vg9KSpcBnV2beGAjTdrY/JhESGF0woDJ5Wr21WXJ
NfSE+CrqYUZBlJQK7EKDqd3yHwY3PRKlHcdUR6xB8D4TdOo9mYCNJopzUqL5aNj1S/BBkQgIRpPe
m0uvMSuXjsk5cVjVsStcFgBuUaCQEquTpPrabrlIrz6ARhBS6GrwMyMkAFVIfdqKFIU0sBzl+xuh
VzUfNnjMEOv0M2nQmqnMjh0kotJJP6Uu758JoFp4V4LlcZfS9YxwOij6uQyoB6ONjP9EP9M+slhO
tzHMP4j7g+qZTTuFf1bBYR69z3Rctrcjc2ZbPf6INKuTCLLZZRMDXc2NdjNlOjsbjoa2HrBMokXN
YIFmU663itz+viPWa+psDNGK02y8vZPbhItaH/M5BbhX2biU679Xz648tauKP+j1hUVqbYfgU1cF
L73x5ZiDoMzbkiqnyn2E96t0RvyP6twJGA1oSixuvOlzpaUs9DTpE7jjLtURGzi2MJg5ltKg/gEQ
xjFi7G/4qaQDnXo4gh09AXa7DiUHtY59jIQk7hAR2gEEYg7v3ci8atGugxOwOSASYCtfUK7O7grR
mbiAp+zqsdXTp3mxMyGmbJbAHExp0nxvYxpk28VCbuCvECBeBM3YvFxnl1rD/9QS3FCSnqm6Ka4T
AQvwnnEKGmI4hGa5OGkVBce9g+sDyHhzmRG5hYAF5koJ28FGDjCI6WbLpRWJVSmclxnMQuOtdx+6
KIn8eHFEUuyOodzT3FKzs3W0kZZqHJuFGfnokaJZ01ZHRCl6fnn0xWy8KG22+ckoZE0HfA5tusl4
3SDNbvCpGz9xxUHK7KRLCfi3dkayRY0RV+PFiANPjxw1ZFcaUom7MsMlnScqVSr3pDEryzT4z2vI
kVUFDKhmQV2KUKD5SxwxESTzUC5qNCUDAa+zgRvQNccfL9mOjZ2BhZncBCPx2N8CLNs0doIF/58K
jUJTcBtkNpBDc5WIafLEC79vBmajwh+c8jabuQAV1t4zAZqgvoHVatw7Dc4fNjkj/MFbH3WcJPvN
XowAvNDRurf+sWosDrcmSkAAO5qDuuZq5c6GZqHqBFD33l0QKTFwNzX5BiCEKyL0RtIKocoCzzF+
ci1Psjr3saE+nuSJx4VefnvzSLyDEnTMPuierPF1s9OL2gA1CPzFpru5W6XqCv8bGSHfWoOiMejd
Aty30XaOsl/Vy0DN9/RaWdc+QfGqsrTkppxMJ6LhJo8q/TvTeN46S52YtoxROr6K5R2H97MWK2NV
mBIHnhWkSDc3x9D6/NwNSiBa4R0D1AW9KBwP+PgGrlbtYPcL0f1D4/72vlR3qXkfbXlSPDm9QC8p
1eyJLRinMQewNCfij9lzzXSSNPdMek+nZ+TSXu+zHaNLT4zZRxAlxM4ei3SIzFId8TgHhRl+sGO2
ZPNMLcu3lnnvyvHcNI/U/xZPi5OxFwt9gkZXa9u7JbyeC+ZyyhOqkO/7qb3bbZOPC8LEIdU2cYvt
x0I3tDIGhPsjUslRD37YWTRR/kIiVW4gdqfARQu2uFBY7linJcl2VmuuyS1EkVJPhLTd7vSSe05n
2dsQb3Ak6mALpzORwqbZm9cx5OCQNGERoqM7o6EZU5SXXlowNfc454j+KlPBNHsXX+bv6dIugHAT
q3c+IEQFcscybiB7+6HClMOwQmKEJWyfvDo80RiUMEexnI5E80HdZJoy2fxQlc0NrhzXUTdmOGQ+
t14WluVv8W7UJ+V9jz/JfcDdeJ8OIDtPsr8LIJoFslz6L/QF495uxdzl1T/7Cxh5KgBt5E/kTQA2
HJAWR5iGSE1twAKZsH1vlOyoxY25R+FhCwWfZiNOLcgb/sfDCLF6C/QBs2WrDun+aqaIc+AfxO5s
C2QEZ+hsyAKS8IPZMCDtEu2DBRvLFUx9AutWHCU2cJLarMFY+m7686MCl9vc5nK1bJaO/fzJ3ZHm
s1EbqOCRMd4Zl3avTCr/XaMU2Y1hhDIZf+V1JD5FtZb+X4NNZ2jfA5mYPqnjZDkCYAYgj+o4Wlh8
a0UQN6B3rR7T73mS7i6vxf6Ul91zRugM0o5dFt4ZT0RR+57gsu7vmV4jROjY4GyTU6vpx/j8F71Z
Fd6rW8qrvdwef8e9Qmolk0OKpMCN1I3BfjUxZKYomB/5WtPS7JrR5EXMoDn5szA9jZsJ9baZOO1s
TkJ07iL2qIzaUTY6evk0i6muP2PepwzgmEp/b3/eUEcsiF3+3jiRkFRFAyaLgQHMarBwA+QZI/Ry
yzdiVifWemcOecCCWaLioqpWdrbthhFj8iRQdlsgqR8lCi+q+3HUXp1V3hIUiott9QJ4eSxn//4j
9t8tT7rzLpEz48S/GuDDvbOL8sxT45aOIrRQIS6M3CgH1/eJJe6DRQhTEEGad7Q/dPjBST9PNf+s
xst9ktDdQI3fA6DGENZax5aA1giRaTSxts556uYUwkzZXDiHEo45ryh8PxB7EiEqSJrFg0ecLZTc
BKO48LrZDJJ72J4/s9sOMQgkAz6hNJzX+d+cAITS7Ipha0qypgM9KHSrKVr+tuJi10ZdEVxC7TNH
nK8U/mFfK/A+hRkyX6mVaYk6BJ+kwKJgScHFKR3jRnbxBRTV4W6M+vF+wcvCHw6wu2E8mw5ZgsGx
WL6sXvEyHwBCc6HEbb3F8ejtfU2sFA1dc4kNL8B0WliAPgFCmMTDNKeWPZoDAl0DN0VQwW5yIFdg
AyF7uc+OHvGHlFIm0pDRYRours82PghrTuS66JUU5yIZowqK4fnKwVkgAVsZ8mGYQMKaS9mbZdzM
6hoBaLcSuhokF4XM7WjA7h96RSiyI4NjTJ7j7opi+FI/2s1I9AdxBQS5IxYzNtGio8fzOEBMNKvk
+s5+yRg/0upcjGu+5IyIaUX8scWtdD39Iz/U+TAL+ZuLkN0xT/wjTIFFEnUruCPWoHgkAYA6pNqU
f2f8lRMimuNzwvW3DHPT355jFH2yLX18hjH+HRyC3Rf49cFAJNUGKF30qCKm+m2fuHM511FaWjDy
kSGFzUwmQ5s7fBSYjKkQBAZoOC1CTPoni01wWRzzXIG6t23j26ngqMQoLVqxvHOO9t0PgHks/9NM
TM4OQ9JNyUvmCXU7vfqto8z4KjZPKfz2+99s08GRpgviTkPzEeRwLRpnc2iZK1DjsQkzgHpAvwAR
jq1/Gub4o+YAL3/VpaqlMe0Jm4veTDAgotINr7paCjFpBSYR22kO7bRLTBRVYrNfNW2dL5EN2hlT
Yra4CpuRKQFotvau87nURQ0QqXdPqv956pP90/uC6KRg3u3YYHpBXrjWFJUcc77bH4vxC5EeMbSW
nQ8Wy15BYEE6ADgf4laBdMTYGTusNzsmnIrfX+Ul/1QwAmGnSVEDCukYvikKMxlkzTjXt9vKS8Fy
7vhoMNv9J4TCVX7Y2wU5NlQdN55WhM/mT7+TZH0Ld6VkE8yisUFKZuZc6bo0DO2cV2OoBnp2ffDh
ItUAcW/XXwBF7srunL4Z1RxQdnpq3ZExnEiTdqEL7+BuslFSF4vCGn6pcWCGu7A5C1/9aoEALasx
alUdCUJl08XyROxD9tKm3OAaE/5N+9IKUTVnWSDbXkBrR83UEbC0sQGFyaXoXRFciwP8mv3ximXT
eKEBPKMGqvU4sGG8SAhcWy/AM814EqJiopKpxUQgVBZMhEo1L1ANrLcS7oUUw8+gBufGciZRY7Pn
FxppWnK/7ihv6MeQecxbqeUqZH1lNAwLiBQz5cvpTOT3pqkT+bgeAWFztys0JhIKj4xFyGjzb4u4
GfG0/5vRTaOKcNv3IUDQ2bmZtnsZYCZ8OtZOiZiXzk6WiAfAjs4Qa2jdxybQJLdTFa8hetGxuxG3
geyMTMyYHmCE1WwUQ5KXDcAPr7p+PnVpzknuSXbkxP1BfaIHcHKKv5PZr4SbENHj2mVGND0xvZ4k
h17MoXQdGR/oIW6aFHsoMq6A06pHGlq2GJDdQ/wBl7k6DU2k4Hy/6GWDTcnQhIF4GqxPAbS60HTu
6lYPwJTlWnaAnFxHojWKYSnYojNrhXgzZgLQLggXngqsD7jH+CX0WDt1wVBSBpHrX4A/NkfUCHhC
b+g23BMCdMe8K1pinMJ6yDfh99lJmPT5HnnOEhPNZA0KwtN/GL1uczyZyOhZjhFs7o96LG+lUUNe
Q/XcwbuMO2AxEv18a/pQW+pHfP/rpc2Z0k2z31eNdy9IPdEIEfJQ33WTz0/BgXG6tM6rO4ujbsle
XEabv83Wfs4g29pShmm83d2LxfWPQMRGEzf2fND0MW+euBlxz+jnfPZTJ8DsFEC5
`pragma protect end_protected
