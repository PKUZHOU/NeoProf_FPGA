// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="22.3"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WMLKbRrP5nvHINHg5av4i1/IO//e0u0Oh5DoLO1IwU3aYEUjqIqrKuz8W/Mo
0K/vkayYuCf2y4Sdk+CzXEPM4ZFG+7rp3cn6l78ZbH6FAvbKROJG/d7qMOzr
VrGp8pn5lVvsquqHbhBvhNGhzblTT8PHXkqxcBSJdMqqrCx8r8o9QXOMVMSy
ISOPOB2PXK+BalfeZ0aVPBB4M0AYWG4XhSC6k1/shJ6+obFvGjt8inYHAXCL
O77TPpaPJEdYRmaRVeWRWQhiAKoNqjFLP9GZ/Si51yAluwoRdTCQrv/M9kl6
zrleoz/aspVIRqZpfTBvlG50aqmX6shntfCWO9xm+g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HeWcIQkAdMw8YdmU7K22EsjDMX0GO8KwSDi0l0mDnpgZS9aAGxEBSSuPoWUj
MWqKlfnqLUy06EA5FhmvPdYiIxRUA6nSE0z9XQGQJIDQ18W3qbIGnRpLzIxL
NbcYxSH7NOl11efFoXbcEvIFYyp3mS+8f6y2ON1ZFaXSnjqRtWSDwPfJiHGL
GzKvmIpc8TPaWvUdOPa4zBH/Z6gU3tQVVmDdFWwk4hgKGMZf6l3V6a1oZz0p
kEyQrdlsif8mJx6tFrzd/4PdU6WXOJIESfPcPncp4ltTqbD72YPZ69g2xZyX
2Oto01IKQnzZW3RJ8bjVRXDHl7oh47eWxAhRvUywTA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PIICNbdZPAWzMW2oHLeTzCqBaz3lGGFfUSMOmRvSjna4+e8f7foWF0y3COTT
JNIIqd/5WuADcKNfWaTsOwn4bSQtAJTuHQVCFJqPeYcui/fBiF2O0bbIolYA
jPx5fr8d7kGBMzKg+ApCzsJxyhZPaW/vPscPJ5kI1XEQziiuubePVqJIs4ZO
KiwVVIjv5BcQypQ3wIFORwJaWmqTm6OzD3IrWT917LFwf9/egi+ie+U3lzki
tyAywMQOTx8wO/gfkcKWJvu5vucBVTcDzu95E8WvTb8EhrnhWTxqvyOvNxDZ
ZLdEfuW1qt6cpdmcNX1YWb1HWQnESNDT4M1Gbj34LA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZBZHCTw/VmvnOnB1/3NNuFANx6xvPOIyTTQ3o+FYHFUYDgnG8ESaowa7C8II
/ic09TAPErqdqNpuxxPyNqIFKBmtlW0tbYEA4+cWDtde2PhnWI4IVMc+jkdl
Bq/aLfQGCoMkF9Xlyz7yEg2k84xb7u44buBwOwXW/eGu800dIHs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
bMX/sSlvnc4n1F+hkH9dlNqBooAKzwPuXP3IVsrxFAl4nDPcOS4oyAgWe8d9
optzTXknBdBFUxwNezj2SLoCWUhraCYUaKV9hu64pxNWr80nc072WKoty6C3
ip8IyBHeIOrB4eIQMPfeCTuPVPTUwKYzDxgCUPleiDTqGD++pqPd+HZxXSpC
d+QiTAcx9p0Fz6oP6iwoVNVeFDLUm97Ioi7xCTKQvq5m6wn76HHfPGoKd6BI
6uppHFh9tcJo0ChNo/yecr3JcJQH9l8MmoheEM5Y9KCOzDKG2prLPM30ri3j
P8lk2/CiMvLE/eG2MAXLAGwwM4dSIA64tiGfkkVnwY5vxVWXPLr5QvBmQKAc
XvvHlptT6Ra6hykunkZdH5j6tPJddqPhMy758wqb7aB4QryYJKNuKh+YTGfU
G6YchJnTzU/klPSgv01P/3ZDKeExRpwtepCEfRHVlUzax95HQxrav2oCYJ+1
FU8/aDqmMlsvVsx/U6SOpckxF2xmfSKJ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ldGwafZXbUpgu/8ZV/iN18JfPL1JO3U/wLthdsHSztMtWRH3itZS8iH+MjiU
n27mxJBvfVK/DjQLlUvrXcThbY2u4xktK96aKSPmgO/jQ5pxY1fJ3uVuRj1J
LV1Fdmbjf6q3qL+8vttkb2bdLHAputxd7bHSeBE6UnP0ezJtX7M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bcm/YGXBFMnMyCNqg0U1psm2NCXjDWQUMcrQ6Hugd/Btu+p1UL7E5VfeYqUZ
oKNriswpcOLAKFWM9vRYeaNlFShp/2L+rtM/Gz6G2H20NxX1V9YT2T30/bXp
Q0QsSJvaZEk6/C39vUu/xYQ7IYn6k8ihvqncSaf1S4ztJZAII1U=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 21856)
`pragma protect data_block
JAksNTdxH59CO6uxqq0Ju8YMl2kOKUr3Q9tZKjglmB5BVnMISPr8wgBuL+fO
wGUBAbeV8vR4ynYgDyfUTvfger28jRm+LEAYw5QbYliZFRu/AfCiFzApRQGj
DONxRaRfBNKEgxM9lMbbBIUt0H2eugzcHVXFzj0eaZteWm6lVm0bVfOZ6Mbx
OxphFXgL5plctlvn5sgSX0d4ab4UZAxkOTSrtjb6UqdRPxxO/nPtsoJk3lXn
1FkJhBsBRbGcDEzF0lFZJRkxLZ9Mk+kA4VIJiS45IFnISaB9QVuG+LvrdJJo
veFl/lYoj0QkMFvlwonnIFau85ICHs2jxVjG+0GZ0ITWiK0BXZM+UIjKBbVU
dgat2Fce1B+uNOnAf49r1+gX6zX6KGl5s9Zh6PPPpPj1bSGDMZifGvzwyqu7
WsMPT2TdGazzaioRB/p1ScOW+R6JZS+D5QMLlgNFaMP7PRU+kDRjfPVOrQw/
q4gfUwz+/PHAiJLfoNbpMQIyihDPMHsFdc0Iu65PJDV8SbHAnoVfHAs2vfi0
KxXsCksa0nkPMk7AazLvlJg3hbk6iOde0vQGzUdXWuDY/PL20qaYJqnsh4+R
P6czYyiTOb1z0u50jBAxYSwzYyhEhRb+fPV/Lo0f/5q56IinWI1qMvIuRkoN
1MBd5i1pr1u7JKixECl6QBjlGT06waYqbyDIszfWikTje0lwmr1yhXW/4R+m
s/i8zwkboX07DC5xtOJnK3co2g7FLN7dycJJ0ZUUerbZ+Z1NupHhF5N9pez6
TxU0W1ghUCt5bVx5aK3OCgWA3GrG9VmH0WQ1uiAJzNjIRzfrMCmZD/fTptFl
oZitZr3NnHsoGZqJGgXZAZ2HBwQeaneNXDlVk1S4NOlq4iEtor3CUPgTdaU7
iGCHd2cdYJhZjqifYn9LP6fz43d4WOF77xx6Ex23FPL9qPXrlzHS7kZOMJwK
2/g+BIuqGU0xG+9r/kEQUPe7dwqihwgm1srXjKgz7OKXXhpd2XEuV5WM/10v
X8oC8oKPLEYKawZ/TdXI//qP9KvmUPgYgGvA8m+Ep3RIrWFu5GNV8Ktf/jjr
mPk4XqarNeFZFDDjkyjnEhUOrE9vp3SCnbshIhGvSCteOypA53LCfpRjvtmP
GEBTXZGb6rQi9qg9nkZvxFaNgTXJuxNsd2SZtZkn/8lAoqkENgIzOeUMfBdD
skmJpWhu+Do37c/wyEo6txj1ZTWbk4uNwilDqXCtTs3MR+pATzAXbDJAzP4q
qICuI1kKCRXZJ97Ao2UcN5fX3I351e8eIcyULJu/dZ9mDtNTlXuvg93UOg6T
bstrIpmi5HaNtYHDWiJSx9pQJJ/4xjHPQ2matHBCFJ4b71y4xzm3FeQaF40J
yvVBpP/xRy0CuiyN/RY6olN59S2Xw+lAQ50ncIH/7zmonWm5SUockVUE/onB
dddr/7ayb3YiHc5ULWvHWWyKPw7B/t+vU1zsgW6LHfhSzsHvk832Uy0Z+LhQ
hbIM9d5gud4yB5T+0FPccIjYDwl1lLKz6v2EG+BSm4lW5MrCfFYdxfyMTz9c
YiJVWEFsCCoVroKiIExXEbNGvcabUkDUHUArukuWw8Ue/8/d088rc5rWGiji
qdi7D2tF5Y+rwg93z+IsQM6zhIGyF/VAiD0uaB7PeNczp59jvr2VNBzNu1Mw
4tDz9ZqEqf3kcCwM6TJr3jhB5TWorrGUJcvwlOJrBUTxQIU9DXiUotzAaD5M
22mVH0rt2VmpbPeScySSq3ipg9XrIFnaoOMqvt+NS/xsYzSMnOlzNkytT395
0QNUvBxFmAMTaMH6pFpl2jZKoYyXqx5FWxS4WefVztaOBV8U7VOJ/vo6w5b9
LqN9HpFSGQYs7uyk4Nzg7mcNTbDnHe3LO8t24Qhl9l6yDTAOXMYANd5p4EIK
wK7kXn92FXtUUS/EjWqlrcIYBxWJqQAyc2sNrJFZEswCb/sGAJP8jJG41MQc
cVd6l1R5zU2JOiBk5smZurDmDoxeSxxoi4CXs5dVGF9UV/frJ1HeQSqMdsRf
gAcLL3M/QKQLipSRZOxt5WDFjXh8FQgrwtayerxNWCBektsflJaAYtDbHuTG
LqFOtGDmAKfikNW6JGNV+wmTBHZUv081Oh2d7FEYM0WfzOumszbR8jQYGYzq
z2YC4xpO+Eci9Pd6AY5g9rQkbNGESvo/uGKYO2XH/EkLJH4VeAlDUH5D7RL/
XRNPxTyF45YIiaO4XV7fxa/c6XVR6DFp1MZmz1wjdqwrzSutkbJEDaCItSEH
8FrQvqMX+ljaVpcIA4sb4T6Ixyuy2KbHupruHnJdcFMmDtkAa/Wf2GnGd10b
gk851YDcvy3JPODg923sQWZSnTkiKr0T6K+nYTMuLGZXh9SlNNvFZpeEh5rH
xQufUk1XgBRYXQmjxn6Yje6HKjfZ6Is+irqD/933F/ew/cFSEZlG2yKYjvyn
wP+/5Ovpxb6QITksrDH/H3WtBE4NXnu6LxqXA2Uf6Y/D/ENFjXFkofn+14SP
JgTqmaSS6Ie+j6vOtdSKU0Ivwt0QTTlxLniPb58Xp4j9Q8X7h+bCSbPiA0/E
Di0BZdM2PbV9zg4qlMV52SLsxO0vucA6MCHE8DthWjf6qB1Qf4GLiTdUP/M9
HjlgkD8j+vNqEj8ml3NZLLnBHWkVLfcBcFmpVK6JVtDyw86N/u9fAMYuZkbB
gVwHv9gGNMCLKEwuB33UkjgNHCi4uzSBlfUIaOs2UhFYkKQG486BxIZDilCo
cIYv1JYrvAXHhPtWwL35MYiP3mxzJLcfVTT0DsIS2wAclV9kxYUd0W2l+zTM
KHMyWt1cTM0k6+FKy5kGPefGyY5XNKPNf3mgUCi/KyT/aGLC8vXgtjmUbKUR
hTTDOqZRiI2DqZMr2lMNsGKiJgFCOtBl+3h0oi5Wwfq4IT9Qm5Z94TDlIdRl
sYEDbCip1Qk0bRqcA1ArvM4X2x7xS5LAivhwaCxYyA+S7xcwDzP0IA59NPXM
ihE+yoijREEP4sQ0icO45QbcOvdMXT+FnQG3nDdQUw8gFattAw6EgJvfTlwn
N57rBrpyi4MGYhcExo2u+TXQwV++NUv/Q9bKMrEw7fV/3rkVS5iRFwxwTMQc
UuQ8nNdRi3lv10HV1btayg11ELChm0QPTfAwT3mglBYgsBbsU7ISy6Sz8cNd
6Mh9F+VeUZCdgbgUuTRdnEhv2OqiCWETRf8uNWVA16Nw1dzJ4RjVHN3KRH9G
H9b/8mPeu0vCbupzJh1HXRAG2puvYB+o4EswV2+0od9MOWjyZ75AjWCrtvE7
jU+dxi8KJLdBdWH06LPCzv9bcp1MVHT8kem2LoWN7x+PlPiA9ZzzmVnyymCa
VuqeS9Z8TxvHQvbGf2CqNbaDDYTmr4WdzQXOGq6jOGWhSHoIOrMS0hR4NpxQ
UVH4EGdk4e5MnK6rjmfiwENyqOjjm0oY4vsGftoAPgyu1AxGvvgPJ00ejQKR
M4tVDC0YQBDqRc8figDFT/2P3NTc3NfcyneZ4DrGMoaEIhcsLXz8wXLyhsx7
5la9yEt3kCK0A6mmEy4EepvKoizM2TE9BsHLDsNJy/F9obilqYRLZHFDzg/t
T839SdNWy0iF6L+tky4uxkDdKfymKSZ582jmy9BVZTH4cAEEuax0EKVMyieC
IqCQU32JprLVRbJyuIonMr2cFoUvZgHkj28PRkt7QboU8ff3LHOAnGZMVFIL
5I5foCdkrBMrMAsDxdcUhLUpClm7FwHJBp7F2s3Tl33qGSiCnxuBsW4wZjYH
cUy4WmLr/x3ikx0Sx3BvGyksj/ygZoo02cywDuK7Ka6t0naHfmkzSItYwwwA
dW7j4JmgXUoIPAu+QudFItAlO4Ov+RZApcNEqnx5B4k0dGviRobjymXEmXre
2z7/is3nDzvyW4DQwTkEiY1kFChVz6tF/8AidyN2NHVJzjyym9X4UaUBKP1u
tT2uG/d1cV1gGcJdjWflTJkaEE9nvvLmDEnfTqSNJU+AeSFywDekcCo8gmjg
SkG+SJL0MGG/jgMpMgueExKZh1u/5QgwRHFfdadFf94FYnnq9Fhne3QWCyh+
+4IAGipG1oE/aGk+uPmle7Dcmqh2B/4AWLs9AwASNOLv8NLD626poLvCmatU
LemR7+PWJwNveNIeQm0wSrBakKtF9VNLIMuHi8beoU68v2wOjE6SXSW5Xwi9
iOqovKwCvDNhLiOpk4AiS40DVCgwuc+93F8rA4qqqXfjX22kdo9M9TiUGzRL
4GRiVkzeFY9Y6wdFZBY2DmiHcsTRJDPXuJv1YMJrgE3ZFUX2SwBZG2wl6PKr
c2ckKJITVCkE2a35dwLM5PYoXsEXDPNqvH8vXolWpI63RG0P0VfN2peDSOdb
olicceMG3gk5JdGwBRjMMMhZ5wb1+Rh+Jq3ZS1535xbnWfJSi+vhoYGg0d3v
r+g80hzlLSkdPzxWJgVPnfl/ClqTH5DaYLB42jivy07hxmhx6ByOGLWS4ohW
iU/zjXbp6vo9FlJKmzjKhpWhGd94IQuPaPvQCOgnbqOIw1PI/bnmOudJkHwn
V1yU/bkR7wQkVBVlj3Dkd25dr1Pg/9bZRUE4arucllgfDFU1O57zf/3Y4f/c
87s2ejKnp7P2yp8ug0blxO7wWLf+hA69FagLqurI/59knYVn1Gl4YRJO8iV2
0H7odHoMtdwL3zi1tekn15nkR4EJv9OP9tsgLjwIUUJHkPW7xKUNC17NkXni
xSh3Q1cxAisauk/sgYNes/F/nF9goJLYZ149Gyr1ld6N5GbIoOFKUo/ECnP1
wcJ2Ew5Zq4yqhGMb4ePz/dtqGs06/9UWTAPYXZ82LG79GrSBZQdv6CO+XQSY
e0nVDgdhFr0Y/H3kcXcCGgRXeOEGILGaDcvlKmaJORifuIGehHUKNedattzC
u8/mKC84TmOkO04M4OyfdvNoSVTzA0MlbsbUp0R7lpRh9ZgT8NhTPg08altv
np0DZRv5+kVLvsVqRR3RnpAg+JYPzFgXv2fitVaenORJkSxuCHVU4HntupJo
tCaqc1ZBI9OQH4en3cEIrpubC8KaH6gKDuKTUk3YywyQMzsiHFJcjjLoQh9/
6FTdelvlig6jjpTaWQiaHYL+iaBN+ksJ8LsK3iFc0LH9pPeUYbYCZZNTOmmY
EwCDUkmJSdlet7LuxSbJT8CJbI1dNoldd+8OkiSltGpZFJ4R1+lqBUGS7PP6
49Z03HVIofGOhtxd4IuDPzCsrvQoAYRal2VXV5ilETg7eLApByfkIWj6ZF/x
AMQm7X96Z85J4PMt1WoHtieDBEGXqsC07ouNWI3v7wv3TndkL815jnbkjjEe
Bc10ZH9tDNq78YDR+KogkN1aoz0Z9fYKAPDIHVaA+PfVqPqKREQJ+tyTvxyz
VqiNJzeLYGFEQMFWPM0tb8Xir4VjxlSuJ65eRnzw5gQPDbmlIK9ZpdyP6aF9
qmTXa0kM+KXHINc+Djk8xVr5H2lZ904ui4Gca+rwRXU34xkjKCqA8ucDbNQu
imaPnxrSFiLaXE+w1Mesc2g4vXXq+PNYtn4kt2Dc3iFEF2u1p6OxvHy+H25R
a3GDXpWjbFP9sT0gPfB5q0jFflrJLd0h0N7ZztCogYkQUEQhXs3VcKJ4jde6
lvmjES3jvwY6GP5Uq39/UpE97Z7TdmLuesReFe6so9S1wZC8jcfy+qzPcS7i
nATMJn9WZMsVKoKnmrEZP/504oGCRibq4W75Nvwzze6LutWgasjoYykZFSXY
Cmy5kED1iIqZlubODUphsNsNiFa1YZPeSJex/JaDgY3ofreOIw9vxX1PBuLm
Xl+zlmKYRFCIFqa3vwntV9Wq1WpXGizBVtzoBoQBXEHBZZtf6acVIF6WCRkZ
N44MPNHp1GsqtjnbCugPdwOxUjRUvJCbMllqXB3Q1wCIM3+KGaVO7oQQ4ljo
yZ4ZXPeKT0aksjZ2O3a1xxE7MVAxmDsanp0tJwjtqiFaReZyrRw92vA0nUSl
BbIinN9stjHtxSEA1+MO8uArrt/0CpNWhTYt+9WdahnE6eo0Ha3wrNPHhmX5
490RvwO8V+QxYLIciGsLzKfh3Zc5nGmKuUxjH68Ez6CPoZ+MSWcPXGCILMtA
d900XoE7MyxG+a+5K9O08XxcD/ECPqbx6tj+ey75h7EwL9I9wlZThiuMSSKb
UYceBveaQniDTJoLkKEplvRipcafIbH0UYR2GmXXYD6e902ZGEfIO41fWBSf
v+nrKkbRoAAC3zfENYE3XNCObCREpzz1vtVI/Autfiio5hsf4z7hKtl8g/Ap
JmaFDrH9lBysrIY7TsUIQyKalJ6tQ+KvxT27008TSjB8TtlVamsSKcagd4yT
z3CjWE8DJ4/MTEOoS+jnqqIwbOq1AsS/sVRJIS6PcWBL2UOep5KVRGbvFt/K
RJRiRfp2bSfGfX8nvXyiTvyRWLuJXD+m9DlrmRZoYua1u4KZo2YWtn38Y071
ugYzwl2x+vQegc27306vhhW3AqN7idhvvEf6ZfS/HoPAihmeVHzzwAqz3xsl
eL53AVKH4Q4TVzYkhyj5sSKJ8F3WOYqI0jZ0h54Ab/fbVVtWWgJzYu8e6HmN
t2kv5m5LWcAMIMLE57CpT3XcFXnWWGuuiUaTtSwvO5pylu73ziKOndF15W3A
wfwzbCF5QiVA+dFsGlZTUBYL2IQfJOq9NJGmYDw8fzORb5VEyu87a51p+s3s
oUa060LAKGFc2v0kHfuivzhsNPM3qY4Jsyr4eS/I6EPJNAc8qtiY8uR9+/Jo
5JzxvTXfO9MJ2kTG5/a7A+rLygOX4ciDdCCwaKmmLJZQ2embuNXU+8ougwlP
+uzqwBHSsIb7YGSsbjV+/e+P3hs27v3uV0JtMPf9cG6MmpUkoyDVmN4KhqA1
VaI5ql3UwYPC1lEV3qzKVjduGB1uylHiYxxbxrzEWlM2ua7wS/0y6ulipHzD
ObG+adQdwooMJ+6v22RSgEQZDZtj31C0mjJgfGWSjCbbWCEWggcabE9jV5ro
Io8GNpyWIq3wii9s0wrwxxYT841FY+YeYSP8E/CkiE9Gsmaj1fSIKF2BZfEW
kHlVQEsTL5z85hdqOdFTwhGhO77/7pPql4kRqjaAIpPQDMXJ7ITcHedv1SSQ
STOk2YB4vfFzoEzxEJczzaetWh1Rkx29kWEG+6KB9Fu2zETNdHkhcDOMyyFp
lgMEXyqeIJK/HksQagPhMCzfdhDMl+Aat3zSoomikfo00eQAoZNibpIuktBg
rDft0FIoaqoaEwdz9u7umUn65X2OnWl07aQL6rNHn+Y/lJuUxofctALiaG02
erxZ11OYwvT7iN1wDNOE1xQ8EpcxAcwpaIr9ebHhKeMsfnNX6ew6vn3WbGz6
izhPkHi70vW0qebZXPJJm+bWWQaOiycAQayIppFZlbMMJZr/jacv+0ZqKich
fDJKNPC7VL7fTVQNrgAC3essPj2A7mc6qffEZduOMmxbwwsOsewbJp8Ec6ep
j+XAuRDCgjdSJFnWWa0gpLEsSaXfxiuuGj7ySUV0uHp6Wl13k/epYp2IavVM
jOerL2YtIWtNbmTL8sTKVcYkQknPVSf/LsyWXgX1n9Hr0pJtI8ScadsAjj4c
xg3VZplCs72qj0pFoHX0GNGkJv/TPR23biygp+0z+S2ojSVLhwg7PfhnAEld
QxLV+BpXzrmgZhhMFYbR+7yc2A8h87DX1zY7bPv0MmEXUk/2ooMOIuVLKRbU
+rtwuVoQQBxxzD9gzLnAGVSAZaexS1xIlsTNKtyn1RDlKQBFsdEjhjjYyIrM
RLSr/vAV4ZSyWXdNL+wzydj0SefEN0OZOPoJRjmf/nXUjW/ABUo2ZkyKmi6l
MhRr4mlO0902u+5H0mhVha4J3vN4uVsHQRAOSH2J5/eoEjvwnYwmKatl5DkE
k33czUwmikFyuz4+bZs6Q+77VnOR5q1QfEit6kLKx+ayS7o/of+YelVF3rZ3
DlW07k6fAQgZAQFx5+9SVKOpVXS14HgxVTcH0xwG581YN11PY5s49aQywmzT
1PRbPPObEBqfLuybIFs2fhFXdXkFP3+NicSkDYSTZYn2cvUqPADa3m8vQ1VL
AvzprZDda3C2wsYZyVvauLA2ddfxzznQD2jCKe19p4xP9CSGGEpPYs7JHauP
S0HFS2zeylmvQGh6Qc9W8zLSiqhXfTOrLm2YcAUTYtqLRskd1tlRIpbyDvNE
M/rJuE3WGaMW58atc9l1aQbXi+rtybYNXYzPPF5W0DPAnlofykh2xKamWtNm
AaFekcc1EZ7F0h5/6vC2xHBkhB3K3+lpJ+o8GmLft3pHrBZG7xx3ky3oi4Ey
m1J15KwtfXUIHNjt+CbFdVPzGzUFLuvJMYJ4+wMkX3b2ieTNigUvIjlTIxWv
Cc7gNpZ1A0LNhS6ee+7DskFyR64QN6vdl6IE0J3FYPrTmGe5+6CylMCMKpqx
C0ury5fLK41VN2W7f1T1JNZXpKxeLUPd5MwQRXXBZuHjU8YC0YWm4jOsy6kF
bZeYF3iZfHq2eQx1oSzHrjPKKnPdZH8pD+hVdmSDdfsfbd9slBRT+8PIm0vW
cLgXNb38+IKBDCPhYq5+U+Wdkq00a7JjyHkTE2X7cp0ZrmATHK7pYMP8g/Nn
jAhpkqCu3w8DLP6SUjlir3AbyQX+7F1R7pmCrSfegX84nVtFmsULUQ652dCH
z2goWXz/Rs9P1ppDNeCYB/iZJLxrAWdSoFXXeuiUWkMH1rIfgKaEIq+xoGH4
OtvxS4ewZcLfrQ1fb2WeWTDIIRLstWMUdH/SLSHCFDkJFt6x1JXSffT8bDow
GuShysI6I4NtHNDqewY1iH8ltS8eR89tfGeam30n5p3Gd+EAWgnugmNWuW8x
bcytNx85UWOYvcE44X/wGF7Wsajqn3FmeekFKJ+J6gInBWtnp2ULivZdsa21
35kv11PEAI8tKa9JUyB0iEKCNAxm1N+MZav+OOUBfU54YiLzg1D9IbjquBH/
eSDQFb/1SISnnOve75+NmEVcOeglEiL3gi7CdB+hVhXJ3DMQg/jcdGow3exV
oD/vnbI74Md6jJfes8M1UC7Yf2GZ5gnnHqnMXsCikLLlKnGKFHwt3d8Y3szk
HK9u7dx17dNmT21xVMCjoXrmS9hq2MjGbVEooOOi8xIyz3V5/81mXUXCDh2U
nIZVxzoMNqwdNj/hISPUC7gvkxqhfPleJTDA/R1GDqSJa11Qtp/Vmong7I/e
++8pB30+yf8s6tolXDkzAAJDwIMzdgkELzVjZsiaw0FI6XJYjPJVN+kBluIK
2Om6Gx8HDaNlzvRmgn+F7FZ975Ol2K4dqZUuUcv41xRrrPXzSCwXZ5qpfBiM
SwWKSTd3lRzRjC2QZ369Mp3td0vxYZjcjBEEPqN5HcVVeHGDeGiJB7TTrfqf
VrdttLRuus23arWqtaSrmCNE145UTOALiL3wVt02l//140BEaWHXkq+aKXCi
E891ZruEsmyDjlW6cZzlb1RXxR7Cy/pUr41r6umaiKwtU7wVxbtC2wCe9Oqf
fhvhKmVLtBRpVZNQ9op7O/Zu5MdjsLiOXwlTlHQFx8rh+mxc+UMNmaMvTNt6
cqWZcdi90+9cDichlCxmIUXYFpnFM4ulAtoH8xPvNlLTMLc/S1wei2njqV6t
JFB7K1lF7AbS/Ihseww2bFh1HJoHOo4EP2omrGY5ft7YvPbVHR4RWFm1cszU
k2YSgmkW+7/0hk3iVIqNgmlmkNtWcDQFJY5/PhHz2oEPDW/inBFUIC78PzlL
e8GqovkMuG3trdIQVq4AeKSRG/RFf6Y1miVI5pg48ggdolYtmCLUchhQWB91
eWlfX0DevgDYiOCs+7ed5ZpKwUaKjFg6du3gYkE9mde0lcCE6bKPChO7c/HU
sjxeosyhUg5NslbaJ/5zcnw6md7X6SUPAssWifgFUKfr+ialTmyoTKPMxHWO
Cc/ynTn+BAYlHNJrctukLjIICN/YNaHwevbQ/2pOQly5V1tQPbfgT4LlC/vd
mWMhk+2a18xESLXX+vfcIICPrYsTypGIjJjmXdl8UZqcJLcAxphfmvAJVJb3
VaN37Se/ISeLzp5fu74eQ7YwVyfXgDDtdvMGPlNyBiM4aJGGNtO7Upn7bkiT
mJonPl3Psdn4QpV3PA4uQyzHh4Q3dZxNoKvTsuiU5+u0o0ZqLheU4u0a0dN1
TZBGPyJkO/d51qx4ru7AZzunrvfaXThBI4O0dSacllEWKoAHQbuVkNLJv90a
bbNDvZL6OyhrqlLIbOQKBI2SDZn2ZwkVa1JILlGZ9f8nf/66v9EO54GFT8Wi
XLsKwwUdECU2g/0GtT499q62Iwu2TCfAPhocxHRVZenX19WALoNUmpwuNkm8
xN26rpF7cEikN9Xf9oz5MnxYDW8mN4tgniqfB9xALQNC/4vFsI8hfJ83SaMH
HOJY7A6IIFHptWUWpww5HXO7PY3kVPu07iFRHyYmsVaWL9VQiuI6ZaGyph5o
1ZrVdBK5x9hmmUjNbqci8q6OmsNjuArVsOTh67Ay/FcS3dPtSM0vIQtK1WBn
qjuRH6jbWN2U3+bNIA5RnUVHTEZqhGpJL27pFkOid35b/dhV9xhirOJWIrLz
jCYYZ8q5+qFkVX3OAsrOzkdZSJEPXfCBFLsE7R9n4lYS/S9Nw0S8NL9O7Qv7
lPtox5HS57TTEibiqRV2iBrT8fqAgJgauNZN1wAjAUmCBGVmxx1qS5kfFKRl
hAKbGBojT62Xa+T1mE1YOoxqZwTyCw1leXQPZF+WonA4l+WrFcMT8GtoQ1xO
3NhJOv6ysJEd0ib7PEqtkoyk57EPrPaMUYvRTBuSFlw74lFMEyTTHoSRs+Cb
u9GO2J1L6mbF2NzFQFiOfV4y/Sn7Vd03LDYkR4DaOMS1egBqgNi24/xeQ2Ix
aizbsFJ/AGtGGnUa2ds20UTMeOR7OQfzjh/3+XbrSMRoKemVwD9WBtK96eYt
J8h0JdeYwD0Gq4mAtIV4iiPlwwXPMUFv2wgHa58tW1Nr1Euh6dy3bIG0WGxO
gHj+nPf7U1Gq1BFiWt4Lk5x8hdQwnBPtjLgy3bhvJVu+jUnN8H027H2/UO15
+szNbTfSgUSas+Apn4ZqewkRCK4mzbI/ZyfCxduaqyvlPrdc+4tHVgA0DaTe
MtzF7nBuhSVI7rbMDfHESFtQn5rmgJhrRjh0MB486Ztsp6exdgawgkbUHqRb
QkASNje/51Z+yCZQKerbfb8qWyGBdeVBrCmYCucazk8uVFP7sJeQrhD/myQz
5HBgTcqfkf/XDqP2G7PZtjjevJsyg6id3gg3ofhwRhOJe6cDpb9oFx6DiNzd
SIT/0JAhi9UgP7Wkz230NokiAU0/OgDb2OY3/sCIaiyAwbmVtXpv1EE4HO0i
lQ2hgs3aqVsj8FHu4V80//2nOngGrojf7+kOImeGQivhbkWmyYiXfik3FNmM
IPdeElFhGqRxP/tlXn4IlziQqjtRNMgJGykVuY/AJeGkxWvRB6XI/S5Ql7PY
yJw/2Jo9qsZSGA0+SowfcLaq8WVCOauH0sD5L9epiRM5IWl/g5GTfPkTWMLJ
NAULwh1HqFTWYh+/r+DxnqmFJgOVtUi95u+946/IgkRXh69rh01KIyvPAQgw
EL/6F87WDCQykTMRzzw1Kfuv2ED3f0GsfO5Dsj4Ylhp+xdCiXi8+hI4SvrEB
885tB9cuR7gtJrUn850bCxSmJNQ5zGD0rVwbtIohKV7t98FeV+MBn2HEI8Jv
iTCgZxkQMP0J4fNm+jSgyDBPfwS2v42TVgIIl7l4jupXn3C7uNEHW/o4fQHe
COdUsQkFpcXh+a2LeRRx8HuEziYCrD/WIXtMkANszsqJ76+CO/VwWsdC2+KE
DP1aYlzzcQfCaOPmIPW2/fXHW1fMDq5EdSEWi2QvpE73iRqSWsIcOO7Js1mS
3gY6ik+Gj895toseMjYE2CpVw2IKbuDaGb/aGa4cLYpQHsDa3O0xVx2UFAn/
mp59fkkXYzKfJfM0qOCTFFvGscSjmErQnSp5vINnDMSSU7eFyVb3Xi+Wg3ml
gHitZLTY32q963hW4U+rrcqNLO53jD6BNo+u9zMSdRyeV/ISt6CG5E5br+yp
vnNYl2gg1twM9QIvSb4J8fwOjxNG9kbsj08rutjEaxOq4eTETOuR3uMG1FTy
pF/yWxrB0HOBtactw0nLQrdhQhZGZCyDwJhw4LDz8Imqgm/F9zLxcjVaEuVf
I4NpZbG3z47djX+MG0AT46tRDdcdgJFfqVnCFGhy3Att8UFhH2UhzLnag1OD
tHpKRLSVPLVjYchF1RLqAPQfUBEwUxXWiirxMUYuK+2ql2ckbV7HqIpp6ywR
60EwzP3zY2JE+tuwGZXxgsZSJE6dDaQ6sj9I5jHm6XubnxxqG1Y/tiksSVTw
zPYdrxcOB6v/emyuJ9HPG154jg+wc0qY8qbQCyNN3YKwbPBqD5gYhcnWncTn
hq2SHeXdz2c4AjMkDu6OtyGDfLK5WTsoU12mNHVBR+WXv9TNVjnm/r6/XXlP
PW1++ki3A5SnOShsR0v8MUknu4mWGtnclNUia1CBq2SSfkZb5Sa/Umy6cmUI
O7G5Ojo6c1NUUinCu+uTbcpxNs17C8lQX7yc3HtHj78+EeX6WbW7Hl8MA3Ij
65ZQYIkQ5Ce7fdpEJLJqtuT5vd07lLo/X5eOYP0NhG8p69OMwaBBvXJgAcsv
LurJsZeGTvVPvlLg62L4IJvMHBHlPXLVAl1pfai0H6LVQ36N7YdOsoWeoY5N
LFG3Q3+suh01N3q9AHcaPaXNpHYBQAMevGPv5QkzgOaQNvam+LOahGGSxnqL
Koi89Qh22A8nZa2Wv8X51sBEhOcgCK6PSYfnB3uPphPZXg10DIfBADm7dNZX
lG+GaVZHxkUORs/gv9+hXNJK53cBOlH9Fb3T1fRDVgm1ZKuFzrUpamRABvVY
JBoP/bojXmZWARFaDbgdPles8vcTT8bkaVuMyVnl3V6FHqBjfr72qulkLt3E
+w+VC16o/of0hRBdgCMA7fNPtAW1W2v3DYVd+uGxXGh4irjdcSPlcpwrpWb2
hKK+yEgvsHDlNPErGJ/GlckMfgDgZWS8+cu8hcNBg+UQHvcF2fpiLn0O5bgF
6n+jZO9Y9lhYX5fRnT+TZ8aLnjYQusalE2pKNJuuOzMLby02fs3kRY2m2m0O
TNHjLiUKu0hbuN360+qocM0vd4CLk/LwqRHpksTjR+ju1q73qge7UkYcvFYY
5BZ4OygUAuzCoAr7JHcxpB5vpAwrUVoFe7LofkQc2MVsWNmIpO167QcM5+So
UFmwFB40CRlJiT31vrWNYlCrCte2CJP1qyaQhtMFQDoXHUJKCL/PN4NSS3oI
zR4y5c3nzIwcimrUHhsxlnc13CiE7+upiyN4xEN1AaRlWf4GNDr6FOjJNksv
Oe/inLKKBH5k4ConztAyESVIpa53/byIVOKM1F09PHibwTnIbetezEBj2kGT
HjMxi1SHUB2EcGVYQ8gOjVah7ScVy8FWYJmx3IYf9KDJYPNXMAcf9RY8KIRA
g21hpdUjFIYLbAnUnXTdOG4Oy5JD2bhXN4WI6y701IwiVng8QgZ6Z78JF/2H
Fevz2KL/B2f9F4Kkxusinn5dXa2TmtuvJ0+S4LYmx7xx/oRqeFmpbJdgxwxN
0s2RCyB2MFx3ShKcgW7ROFMYV9ZufaWFcdh5whbZUaGPUJauE9jGxSaPNZ4t
xHSCHAN4vgx/toevYvkK5CdbXTT8Ivy4iG9VCr6rRk92rTwfz59nG91RJ76B
ebW/eAfINWb1S6l+bG6CEAimlQmNTzxarcPVG3O+ewAb/uJFm01cGXCGalfQ
U68LSwI8u0iQk76Mq8VHnpfOMS7bLdTL12wSGZutTogl8x59DBBk9dWfRxZK
EmxNa7671tr17WOkRU+Sita02wEtvY+JoXYoHtYRzeF9TW5Td+ASRWsJ6KQn
Tx1Cd1ulNqhFWPqZCcJ646+IvrGAmvI/BaRH0Igimclr9juxhkBe0OlpXQ4P
qbg9/c4Xq2J4jkHEg0ymIoRxCusrFPldxOiFY/bX35dILj26JHo6Xo9kgtXO
9wbxbZ66ZhON53nzK7f/ICBNFC4LZiHbhVW1u5MOp+sXWkvXQ0ZA0OwsqglL
Yr9hzGqVS31WoRsizYy2aO+ylSTWIXv0TcDkBuYBip/9+EN8S93zpsGOcAbf
p9hUKc1JEhL4XMB/gdE6E7In8qi89+r9j8GbSKa/ZnU4M3fwO3vYpNLYKC9Y
xAMT7ln41rc+Cir8TiJ0IdH9srTHlBwDhtnyDcQbapGd0p8xw53a9EoPngvT
nn/pL8bXv3rs38vp6gAC2XnHDgJzEhezU9ATrlEPXIGxvCMf5v3etU8WHHz4
e8VLSJ3NINpblCWb/LYjuh5MXnuYZyWri7mrSgLVMZuKwKsXcKbm6ZP2HOFK
oLDzfNOPmPXhSNHlEz4aaISU9S1YFoeloRA7kXHjbDbajDwN2qdbIMprLL64
+BSAx2Zg5vEHpyk+G7hC0BVQWwV9h9IkY6/88gtBbq970/2IPCH55dKkqJm9
+jIEu33A1+cZKFDgfjHOe20rv034R99eou+nDWXM1RzzkduC1KhXwD2UJzp1
Q8szBLH938CyAGWos7ciJWt8+cvyxdGGoRgRKJDg5KLvgy/HM3LxcdUfDyW2
aTggxPtLZ7Cpgvj79d+GdG7Uautc+ixIPfFRkg8JWtW8PruTHx3vjOMDuEKG
1DP9+L9ObAYMZT6LJqsODkg4LvHgsMUajbCu48ThIY5++7b5pRQj9O2PwMdq
EeT9ZRATJUzBEQ+BLaDuYYrduPloBT14tapmmLl2ENVWcasjTNipv7ORcVBT
B9yL24rPm8N2oKZBTMvFTYeWSk8/Y9xJNGr5ZO84pFkKOwHd79yfvsNy+glN
TozkrCJSZJGyL5wupSd+BpqrqrY3nUBfNiYL2bYzLKSVoHiFqz+089Kv1qlg
gaSknrd0jfSr8OEyjdyZRHpeaj7mqiPFAMMIisJ58Od4EMZSiT0lS7Jrs4Jl
jBcpby/q9A4oc96600V+AUHaToSWX8ot6adtrUXcWJW1gzF2e8DSQIFad0JF
sNd+1FkcwttIDpn8EB1MVWy3v3sZ6cVOuggK7+GR9Ut4SHsRG6+hh2lkAZmO
UR0K2KK35nWaQ00RYklPU62EDLq0Mpsykg8RwAkOwQQs0iUEJvYdKiX2/bsZ
n4dikKxuC1ODkomPI+3krtIb0h08ZfpWjYyU53qIU+LqtWRx6CFlNX5ABWK1
K416MnGwubWYrn5XYnc0bI1QIqqcruBqfuRgQrYCnjcrixtdEpGoQ8sjmfdq
LsjqZp0jZiqijfR/BuVC1jc79KpZgXcEFxdAWvy2qBR6VQxYkuIOdrOWC5bo
R2WxYMzf1cUolYAtNVecbTkVETsFJ1GuuKgrYjoocqNiN8sHJUYveGZ6djeX
NeGWe1dRz7afAHIG4LLJcY19Xlyw7+LZawdGS/RXhbtypCbpHjdkU0CwbQqZ
2RXfM2Q4gJ/XVpoAZx2LmquxTn7fT8nTQZNR8EeQ9yjOpxD/HNReKkRMzIc+
a+V/exJvFRqLMqJn0UCUXgUXZ/Pen2OFJKQP61qYlwDBTwChnsGgGN/BrgCJ
D+/KCsd7PLkWbP3cOWxROPzBCPqUyNUlK9X4GwfdBTqlSTSWsSF6gav5h3d6
v77jldYDXD8PW6JwjxTR2IgPwjgXjTMBbo/DI2bQFzWHjHkOHjBASf2MI804
Nf7VD1d9c0vCczApnZfSJDygnR9chICLsXRPAnGiyD8Q80ET+AXRwkedxGDV
n34iEcW4dcBAI89NyGZiC1hAueXVd+Ic30xd2sZ04e7G3wc8CC9rF1ZuGfB1
VHb1Th/vVNMZYeDi/P1Goj9Lntv+PtFoFP/99hbr06ujfUyaZdvIppgUQ/+3
TljSFX4tnOd+vKas4pkPN5zeTAqsm+XBnUk/Bnk5i9z1J3N7Ejya/itlUNjX
zzluiPTle2aBpKvn6tY5dS1XRPlRRKouWQmwR/IgQvN6uzXk1w8HHRDPDGRE
JernbbxwPejPz2gvSKhyJafESxswMuQHYMK6B0S7/MXKikN6MhgKUUjo81Gw
niJ7GTeIaB5DsJTmookFzhWKzCq52UoAKDbc6BjXIgaU4p/83bJVOwqUaAhk
SZm7ZMiDu1gpdIaojscySNuWZyHqkYcGnkqeD1uvFV9ygPdgh3bfGTGL/TSg
P1z+bZ6JkxgSMW5HB0wIC9XYxdsvemDYyS/0oQ3EhBvLET27+KtBdGXOBZE+
ptfRuhWhKr4wYiieflgIluyN2i8YgnuwCm/pIRXNsJLhMl9HAHUIaWeDOfUt
oz1REsCwmO3NKyI8u4K6EC8awG8AOHCytwoQU1QKj8K09ty/fC4tlT+R+2yN
rN4SRTktxjHVtOKU7JqutxpJ4HMxpYYsW0LLu2XVjhu2WYxFK470I/69/7ZX
Ul0cja1WXeVOw3we2PeAVxKexixSN7Y4u3bdVvBzGwujLMdTTZVUCcTvFbNY
Y8pXpq6mPkyoIARuMd0vc54MpTKfIg51PApSMXi/sWHtyYANRe7R1nu0+EJM
kPI+n5BunS0jpe0Dg+nza8oRM5pnji0aZowyhxiAuPzA3JvPXfghhwoWi9ST
Ew5RcA3nS0e3Rb/qTVbEIMpPEszsniC/RhAU0XMRlCJNOODnCPhRWB0q28Wi
kkyBCHEMv/Y2y1YRWWFiUrn/iY0rhxRNuN4p5ks7R6ByvAWrgsYLMQDLAg/M
WUp/0NCgcXA26KJaxoHYvTyNbYGO6z0q6H32WGDmPfRcM0JrTH+TqjLgNpta
pyEeI2d4zQI0FmOUSADdtZjZesPuuPtKxxDQ1KZNguIEgaGAWbxNPF87i6I8
4p+ZXx1/SBvcMiU2yTrVrSaQynrJvbL3V3G/LmP49yLUD3G5VlSTtrdkx0BE
VWtngmslaGtHxxvxxgU345UwM/7LY8PqzP701mIEb26sZ2xziWF/COKHU3n6
tYJ4dDLKDC4lxfMzX9fs8PqNpM23tDizeHcQvM/eEI2YPIjbcg7OMq+6WcaB
VV5znafjUOPMouy7cwsRI9LHMzOmJ5lVfQT5Eb7XgqZk+LX7upTInpbLgWVA
LHuEG6EW24pRBSDx6ANXFfYlCTeJzQxOmOidmiaVKytpRw7I6NkGZABcymMN
kPtV3pS/5lbKPnWZpCfl5chyoISF6jTRzRauwdgiFxwjx1V0z2VAyr54qUYr
+2lSRHLc0plpoajVAkKLV2pkwEEQYAcU5d6oKmuuKcvjEDdp9Gh+xhZAra45
gwpW9ScleAXmrIgAlpdOLEh7KgCz8lZ61OEpxvtUWvX+0pK56eqBxu7iNADW
44Dqg28op2e2TkNKiTlacmb9HNzh/DWmUyhKMkEItTqnK33kmRReFAC3xoKD
7cbZ90FUT6WHGMuJRzId20hNMm9mtWVYs3l41Q3L2z6f9YN+M6laYttGlOOl
tNRVYiRXVT5tqQ52LqGu/gefPE6xn3ImFr1K+eRu9JcFuqHgnTmNTrJhkyQR
mC3S0bSD4Z/Lwz1cmAr7q9ihub9NFc+Lo1Pg3wY/uxwOnEfZIE1V37KMUIDZ
QAHF+hH038Q2U7KY2AYYv9tPLqfRJWkwCfJcLglSkjpeoAQN2LDlyGvo4mwu
/ZaV+CJ0zfaVeOAQaXoJ+4AOefdMStFxIkAPnbVimRbEu/r5FAj/P3ISEb0+
AMZePGWKzD4p1nq6pE7qj+SjKLZ/0/iR3diIrGzniWyOMZsG2LjWlqlTRse5
c9SSWU8+73OIL5EF3E5h2lRzLr4AK7j/iHR6XsqIz24TC0lQd6ZvoN/26NmB
H+1w/Y/wmjLeF9t0NKZ6YVcuOpeJTiRjBg1eO3mMnNg6dNYuy5KaIbibVRUK
rNOwBxfUBk03KDXGchhASmqBjYZU52VFs3OQKdCKhHPEHCKALqRCFQo8atjA
xRtObqmFwKtZu2sLjV2T/gDcTKwrbzcrG+PdaUcVHRu753Qmk1GYTKdCpUFg
P36J+l2XzDIbRMKtR943pGVWvt2SKUNAePCSns/ND/ubKjPeqv98CJR8+NLY
NK737yyhNshIvYO2muCAlrJKf+uEa+sFuwIwN8w5K+9lxpc7cLtpUSrHXA5G
I6PKtL3y0SLTce2+xbiGbaR6p1OvUllsg8yjUYLjITKnppt8xKrn8iYk+Ha/
bQ17Yrm49uJ+s/rONgKUmIMalP+8IjUKhC7gaaHsWt5LA45/8cvWYwhknTud
hgCuhT7YxPGZJlfbDDDxELpP1AJY68BSHuDz8I89rnWcaJuHCtYOXH0nqpA3
5YlcSMLS9dgGxPXYvTm61h0xP9vDOELwnLUj9tq1k+3wtrGbAc3Td1MHd+Db
4ImSTz3+dQGzcqXN2Z7EnqBOdFJuZSlnuOnTcmh1Um7e8QB3kxkCwE4TFpg5
Jz6Az4vtWB4aB3TkxkyAP/HV+KTt7yEyeXdz4EadNQ6gdVcesx85pFEmxati
k1h+pTJaV7MSSi8BBLV4OHs6k2wEp2fsHApRHdw5TexEbxHPiEGaUYN0C6u3
/b2vfRchylZHBVi71NPqnUoPqhS3xyhfPQKxpZdKEz7buQd6c73GcdzkuRaT
y9tdDpChnDFWSwa9WXU1W4qMuwmUK2m0DOVCk1r5aQceBuxVJNoz7RPlS94x
+Agg/POwTH05/KtGBaRfJ+ygF8/bpHhOtf7usoGWgAuJgkxYawAdyE7lhGbN
89pGmKXXUEIg0mYCrW2f0JfWlkbE4lJM7gi8Pg17fQ5Ph0eTs8dYY2sKTx5o
v0XMM6wvkZKaOVGh5n2t6zHzVvwV+AoqCCAcsYXsCyYaYbjNjHH9kGTqhDwq
TkARIOlMpSuGaSgKIYD6eH0Jh1BaWPdq4xWBGhMulEm5RHZZTnPHRY9sGPzg
9DKGCfZPFkxB9SzEyMNWAMa0Iaz8n370F/dpXicKzbSapcQipv7+XPM4I4b1
mBFjU+lpifRImGAGAXJnakQQdULXOjorjaANA/7xKRZ1LcnPtFeVwpwT7ymB
okFmFI3kpVDHw+IkZ5miFdaVQqw6HocGS9CVrAqY6hJOnJFI1of7L3jEDe+5
Mt6kUk5/dPzqUJ/k/uF8+464E00meL+h0NokUqoQ/SKDGfcHuulvceY7FdXi
lCvnHyS3/8lOxv1ChiDL2PXzugIX0laNVyM1eTsP3QxSNZeCtWKBXqVFk5re
zo26/zqiwxgZCA9f6CezwqTI/xn7OQpQcsfNzA60AOLhbMzRIzhBcR2jU5FF
vZjRcZS8BIrYqbDE5cgD3jm0otXNT/z4pajKyGRokpFSZPaXSjW47ZuaO63F
iR1uB8Q9cJwvLaCNcXWJU0mb3xXC1N3MEujJNa0qvMhFwxaH3ePufAhrIR8p
JeIGv/8Lk5AuWQ6RbNW9bia9Ot1TF2rGfjXAstbhvleXN0Bl3RFiNeYouAgr
EqdLhqVCUH30hceOKFdYuX5uTG8wyIQ4KCxzROjzbDz/0+4fQ0cy+GwTaj9O
rI+DAMzX6L/u1LY6F7G1qXpJ+dJEIigAir+ZXdMysK2pr+Eks/8ILFOIS9Vl
p6GZPsQCY9fXPIMfiL3dJS8r3CeBcusTGbyk8V3ydcnCZT01FxGW8rHjXTh/
Kd73BqZYI3O++sZ3mt3b2edHVK5Jw55dnbU8fYLHqJfm6RbHGTZMB2aw5GsD
XIj+Al5SGtFXS6OOdJsECYUiLM/LXFXuhqLyw3cXcGx+jz/c5eOQEZ4lmxoU
C4f+dPJf73PZa4jKA7TQ7fREAEoJuoO1GqtWaKVKmf6SpxAvNBczxBzWtzF/
QhZu07RplBhOJRruaIkgBCswnbkyB7hze8eQ742dWbXup8Gqo3Zk1PqhYHaO
7j6BNNnsgdrdRAP4DSy1oA14d7J+gVMeZWSfGAQ2342ZbkITmKUGU+hT+DXp
nwa8xbNjPf9YnjwtEzADw6+xbmL5BNRBZHy5aDZT87XeIiVcorVWI5Fp3eYq
kvEwGb/qb6U6YHYuDQZxOOUW2IcaxrRFGORv1fgvtS68iNb8DcVc6B/1g4bn
vEvlJI5fyvm/cX5NNdzJpE1p9SIMZz3xBPX3AzA6q7rEM+mkPGjTsheXkB6N
jVmLXp387IC68xbQZc8hEYXQT8ybAPj9Hl4WQJ5zo5ys2t5UHVNyso38b2k/
rnh9Rywlgjn1LylqJW4voJ1DFQV1zQNy0+EUYAel5mQZ/tMFiqwZOxBwKpB5
nF5qpzJf3mlKrr0LjMTYMzjkYElen3CzGerOzFroFYVY+11I2baRFQ+z/Jks
b2Ooc7t00ZcuWKGE+5m/pEaWqnTeIUPjw4QEB087FUWJd3kuRpMmYcPl0Xa2
Q/ncHS84F76ef88jc0HXWj4sOAvmE9WrouanutKPQWDcrYCyPOhkJuOipOUs
JMzRqv/4dgd5Jtc3cxcWXz7vJVBZIZ2lkgpceU5H+iqKeP6EI6CYI9fymKwa
7t7s4aPvHFsB1R3Z7X1aFDtd1mcEz/JBmPwablY7Q6EpN/rLuIgC5UrWOLFh
ugo8mnS8VA6kZfLI2F9QFsjOqiFW1Zp89+LJINNC9tEAnjsIvBKsZhgI5tmQ
TwM/nmsU+mkheN+NdqFJ57EDOuXp9rSlF7unfKEdqEstEBFd9CN3SGt2u5nY
kEmcenyTRqpg84Tfk+b24Vkdzg69r8cXne6x0uyNiVINlWi79tvCgD2m6Joa
Y5tAsLmew29s3JCl6YlgP6x7YBMp6jO1rAR6GO4TeUZNvZq3AjOgyua5/lcz
KpD83l9qxYOtFQd6SpRszyzgOP5bCijuKbbN+vhdhP0X96LFrMoCvv40v4vm
efY9Id35wP2god/wYjNOOfjdb16givDyK4ALAicy7un3myNBADRfN6pQ+oyo
zDGcOYUSC2jSKcoI2YasYKyTyfPKgBfLcUqIaPn9FvCiQ/JIRfb0IqH/0tMU
PvksSL2PYGGGdGGrtyZVj1KTUaw+kmNbtoShCjuHx3FCBIZkppO1JCMcElcF
KrMeubp2KAPUuryYtpY+TmhBBQ2SkI87Z4O7iz4qp0NEz02Xq5SINFFtsM9u
Z2bIr85TO6J0C/+G4BoVkCZ+LqXLKNGZrDs+HpD14o42a5DOSlar7QdO6b+t
9R3MSOjolwHRGn7vm0PSxxG9U1KIRS4DM/KYO0IYhMkyc86bncyjrkr/mokU
hsQc3w20Dtpxz3MT1Ox1FzJbpIo0tBW/VX/vVGeDcPRFMF2DWpd1DKSkfaHP
w4MJnQjyrmcw37OewMhs10mKyKPQ/m56ZbnSXz4ftcVrqhv9wlCSt0ExVws1
vPmjkLQ8J9WGkZJIV97Baqq87UHmPxtlis1GisN0hC2nFuhXkVMZgWpMlAsi
S5J7XC6GQvpzRK3Y5iJo/0ko4NzSF5OiD2uqCH3SIW4XtQ29bmbbfojTR4HZ
4O0vF/6izIyYudFd1aKXaUfcCQAnFWxexkqH5UaXEVTp1wMG6dyS3B0DzB+r
hSZ6Va6ld0NUXJEohTBZ/5Z4vPF1yGObfYO1d3b3wuTwLJ8tazIM78ePfW9J
efFgJMowwPtlQ7IuJWhK3UI5x1cdd7KgabPAYQmpzHBHXI9lfizJdxv/nDvz
LWkEKwdyjlUBUhQaqe5XztW7BMx6Yu3LWInn4Ep3F7koGRVFrnuRomC8Ah6c
66b+KMpisI1uDbCH6MxNk6d25Pc/M7lz6ilyQI1ugzrNsUj+M7LRNSMCYE6p
f+unqZGfGvXOgxfdJGt2otbBF41N3Dc9dyEXG4WpLAiI5bRu7vwrzxIR0UQB
F0fF3LIDdpKy3w/pgU/4qTgCDEq3Iw2vTIl8sqEHk9AOzfsLXEDWwk9bLHaa
vU5/dGOxRZSr2ygnVs7pCrc6G8S20ISLSfGNhiSsGxC7VoTHr/DD+aZqzbV1
P/d1DrykRHWr0P4wBBE3dVAcY14nlt1+I9PVi8wCx9c5/3U1ppqbqjMHNAk0
4DkgXOalO1XrhQJY/PA+5XT9uNzuAXRHjqkR69YUXuzYysEtYWyjxHOdldP+
Xc7Md8fKuYIp1D7AaTQAMo/Aqt2d3r5XkMTpRgNIg+Qq101oiuRIgSfEwWm5
b6OLrz241CP5SRclVrrNrKhyCF1fHz5HkgT2sXOBbbhfyAzdnp0QYBK2SAWV
HpMMz/AxRnfZ7umdSdNxEWdqNNxK1PnOcGFwohzaerdKrfYmYR+9L2QD23p2
ku5gKByg5/Xxw8M1jQ39PGxCpipnMgPiAVwWJnFugX23ynDxSNF1/0IhDCUX
96cIob/WKA6NPT+SZVefGrpTFFdkyLVTpNrILumBQVEkdWRTqyFDGO61q+a8
/+WhCXkskS4ZkcPBv6aamFEVVwJUZC3u5J73+98bWFuzSj9JxGzpxNO7Q3mW
fxfRg+/xfF7sAARzREn51V+8Hz5ZHffPiYNuHGaP9fOfgJM3IJf0arvel2iI
apf9sCA7iB5zfYUYvnbPkYZ+D8y7YLQ20bP0KXgCnMYjR7A3V8f/uXNlCgnO
PTF2UnzO+mGL1xN9IoztGSYyn6naREe8n8AJzj8uowNDazZUbXz6FjAcu8JK
XO2qmOPLioU9rLzeoI6j5VjJJQD3bN0ZMCvaI9aV0nVXu4QUl954YgXse8lU
OH0oiyIl+qXPIoQeCVmOYSnpELT08nNlxF8SKcT+4PN2882vrvL/vtpBZGA9
8VQPYq+zlyVKiz21bBJzJVMWmF+3OHTscmwgKP1dCCNLP7XUC8kPUocS7/j7
UuC66VXb5jbA5JlJPSd0aXXz5Wt12BPkZx4VzJPjAjLElGg1GhnI1Pyr7Nty
KvrjQIbbSMZRRYpLMd7LqaGm0V1mrj04dcuy2S00cXOOOQTPLZRyIuReW+EQ
U3X62UD7LNSynNa2t+MchsgbFNGz0n11E7G3oc6KeSi/uGoSQYeqkE+FYF/U
f6MlzMKq8oQvJhcvs+wxZx6OUGhYTipGTmIkNGLpSnAHwh4g4V1I51CyYQta
oriWg3gHpa6K+4b4Ua/IPa7aJAg/DRS9K5edaq8HipRv/Sy6/xC8vxkgitMj
RYurP5fJAmR9/bKUOCnOEYf0Sn2zSyhCDXAzh4GYMBTA2HywMb/Y14wUOH8E
wLfn7ca8gfsv0nk5vcGymq/KJniuNmXxmgTQUNtkLZXhjMydlhYpwxMLxdSg
IQGoEMvlK5W3gS7Uxt3+eUSt6tO66Be+esQdauPv/mSp4vbI18CXmAnYOBLA
NtNOAfdJ9YTTcQzArhmliuPC5+N8mZQq2bESbVmS7ci3Ckk7dGMVFPzXoMwh
hjLO7fpHoYixM3cyoZqV2UIE7Yjdm2eoqqyqhxdKHAduJX3HgN/BESvP7Qvf
NAYnUqYu+wshmqrliZN27y1TRkN3SAyUtbXNat7RLfs3T2FxVT4EsL5Mwxes
1D1S2DFdVl7YP15+eM4pkEgRzdh/EidfuG2KTP7Gv73SDG7ClgctauM3/wuy
VvoUMBgqSd4qEiLo70HglImEZ6rUJpU+uek82TDD/Skb+wGlXQJ0reAz/N4F
QMCVsJBKE9vENU+WrgcZAibVTP95qN/z3cvfKZLC6oMaKmk1/hFLZLq6pyL4
2yiwoaBmfHkVeZvGOKO/vOlJrqnLUvxdz1/LlOmtATGYun7TjdN/GcSPJpLG
qono07u7qlQeHQG5UE5Xh+E9lovT8TstK4xGhn5TB8i+RFHEmm/FZ3AHhDJD
yqIfUIokTEivTDhmTUMMl9omh9hCptNI3M6xt/AG4gB5hJtCFCZV/kqE32QQ
xYXfNzvzBO4ufBwlSfBziUBZBariM4elJ24vpySiFrYyVeTQITNur6ax1d6Q
U5IPMtdVlAiWwa2DNqKe1KQ+HOfgQq5XAammbf0R25TdtMqK1/8yvXxhryhS
1/wi+goBf+ix/BAkAEi/jdyyQUgnESYQV/khlLtYrnY+n53B6/IvKEcdYMNc
NyyLBKqPDzb1eS/WdJsPwAsxNtP6J+YCWcwhxJabvqUJjgaQXDp5Lyw+AydY
MMelduRh4xFwYn0e4HiyEAiEL2FS15WghRkQrQSMgcprdX/7Cro4d2nqHtyb
KG6AtkWuirhNTVLGJPfmccexQdsUwzMP1gxKZWdhRYIwmySeuzKme24V1vZX
ReTg49BscH05qGf5X5Nulyhp5VsHtKudsVYXtJKD48Lx3OT9W8BsvqsucAxi
U0iaR7c7AFyc07P79z/r9jRHyfxssvizvbcShNZ+4KPzM8jEKaaku/HGAtu8
EVuOnwZ7vcBXXNYznrk8VOVYpuoySOgcNnBElvwCWxlHMYuviWFfTw/kvWMF
fCQUxM3xdynunXF+hysWSVGsLXiUEUT+VIUOHwz/rPiLGCDSzrMuRgDIeLRD
CC3gcyJR8rbaZm48fR0h3zY+x2/TlNf6wmbaLf/EgGTUPcfWwzqoNW2UMJdm
tf+cgIqKNjKg0SR6kwUy0JQSwmDdqE88234HvFK57ZyHD0K5eTNW7LaXa0jL
SFN8XAe+cKL56TtejLG5D5pvxeNYo9UYN1stFTBE4cC7PgRoZZ2HKQrujPaF
CTLy/hSyTLbFccGKdm7uIfvdFUsL/gAB4IgvrxVbGgxwcy158KHhK4RugQf8
3u+LPbFt9uUju+Xjhy5dc8RGSsnIgz+m807UPgcbCq2OIUqDfS+OoLzgCaG+
KD8wFjAJsfrnV4mqGV5MoeWcIWIE0tIiIT/hv/snCqV1XHLDOEJYCVILuMiK
cZjGhQmQHFmVIWInLaEW9k8I3qqLH/FymotPWyQnGKRxsRpOUMNmCSjJatyT
2kJGqXN8GB6oBxR9nEw69J04/fo7Wthlye3dQpMoKV8TGd703iJfcNmzYzOr
hTSnKSbGhGPBpn64l6tXH13rRhrc08UcQrUAG8GKC4dXvjWiXLicEQsvswEp
mm5PwAeJWB90xmPWCcRLkTEYf7T4kPeX25p0dFFwRs3xL9gIpoEFRJwTEmgh
bYkVXQsk7HIwwliU0+KhAJwFseAibFX/Jo0VyAWuNfTKPxVN5o7umXLEvSTL
zJT1bWnPguasXB66RKkyk1OILn6HQYhpm2GMedeU9d7qpN0Tzbg0OJKsMsA/
13WGKAtcdY6qNfmWrRu/EbFNeQuagLXu0SHZC0tUynxk9pfYRimxf+L3chKF
/iKbe1HyS11VsPTKdLMUPfeIRdOvtbPNdEDHSMIj6+Lmv0koX8EeiqHSeveU
LBxrhqJkHeIs2aAsZGPEa8SiIHnchGqBQQPcVZQgngIdBJqXIZvMCCjizA6y
Pqp9OAXD2zFG0IfblG3rB+q3U3dZtf+ly5LVzlgpBN9ZpAyzX7/n0oZdf5iZ
KcELClnUYNvQa60fWRPbg98g5M05ksMrQD/Z6Pjewte/2JfhR6Y8EOfI1tgL
095M2bAqISzoZW/fwjFuNidxpKH3qCzO2+hQxZzt6y0GP0f4bvNjdg+tdSY0
VzzLmPRYYoLEbwfAmx1m3gnBn2ce29cRL/WsQXUxqsCXj+bzO8vEuZWv9Bym
ZvX2wDPF1ZeGnJTTEyHJwYYRRsH02UpF74KaDW/q3Zxtua8dVORUnhJbKkVT
LQDhxGWNQ8cHKREEBtUZ+epv9aO/AHFtOGmKa/l/wvV+v5lCfGHKFwF2ME9v
+CCDg5nRDnofOoIqtALqYTzVEvdlectZAYvEQBespC76EBxfik/GqlEUl8wS
C6nhcNJqhDrCkCzV0ZLsJ8yaKN6buTwTMIiJfFHDfnPAQI80ibILK2yriNbW
WCxQ2FUniKRc0nW6bZhFtDcOe/yM6tZnK0VBQOzzAodrMCHVRnKCuCz68xm3
+NtZJu8JZ7wjxE1EWMTsvXWuu4hIgxGnM0u2iXp5MbVheItuV0hB00Mh4xKm
y9nf/R3chYcrb8nckeBIJQDnzggd/p/aPhMywnwaOWHtwwVGx6WmV66k7GFB
V5KhB8AogBKECdrrsvw8i4nLuDaisOM2PNyzNTgnAGjzCZOvUlqYvXDgo/td
l1ugfDTQNMUFnRmA2oicQG61C8rI4zabfYBSvOIB0p30Vd7EByiRfI0joTe1
BvDDvospJjETRsxdIP9LadconkXBNCtsHGFy4UqqtI/UkR4nIrEfNEb7LIi/
ls0uCw7DfO5G6urwGI31DK2vi/tnlKca0qIlw1xe0911Jw+B3gwkeZU1jgSP
+RI1yftRhg5ClqSLM/MBiOMCsGONBjIDD+IHNRvDN+oioms6Z56DJy5soTZQ
gMYvUJwFWHCkrFXX398lkST/YqMKisgnZ/T9+F3HGNGbL05s02GjB12PgjJp
tdnukeSJccPIS2LByqY7uDicDKe5edi08YBgt8KJOX73Z06d56KNHkIHeDwo
2r+kL0hDcdKfKz2RIPoe+iAWIlXaBjm5O+OdDFgUGN7Z9zW3vrbN8Jo5EHZu
MyltFkYpPvdIBggNSqDjnIXSBD1/5IxGAWEG5UkgOU8VhpelFenf/NPv6Rde
H4GLz+6m4gy3KuzBVMvcWcvdRQiarqZSnhlei3ZjeEiOWCwbQ9gbVIYpZVoQ
ppUX6C6TGhd858QwYkMXozyrJkslAHD4KKJ3p7jY16hTF9GofXh02AP6cdLd
sZgn88Vw/d1U1r7cMTnzTfsWoNkgOv70/nfk3fm59qHXGvxIxJjY04XvjiGN
DanwVhV6vRUr2V3C1p31wZ+A1+Fk4iLZXoydlMhIjBWPwMUXI8rABKw7T7VA
e0iFicifnS8iMfgX0QRgdAhRyLM1qqghhhyeqVWbl6LPylcA9RDEj8QCUrY+
LtDj3xTcf3gQ1wDsfd+V4yoFc4M8KUW7NxjctfOPwfAqc41VO/QKC7pJjQqv
FrBl3Gy9oy6EIYZvvVQ3n06CkroVqKTPonRNK6hT3LSjo7jCp9foKTQsrowA
tTZeQmUUsTzLPaSRqhzDgUk0N4mb4Gyj/RnQl3wF/fJXXE52LJyV/GnIsikd
sHNjJ64kcy5fF0WU40gZYTAr+5dcdtJjGAS/jjKRBcn+hwVrx7KbYkXIpcSc
SQWuWcZNUfe7IYS35fiC4tdEuIopI4HTefgTCPQygNRBwYp5ECULg1/Fj9Ov
UUnNNwVIkP2vqlOzZ2okj6NXQPzwGnoWTR1Feh8f3HpVWRVZBGWIG8uWBJSi
e8AfFpDZrDDjmDG/zvKtdoIfbskhbifSTF8wEEdczWOo1DrAEqXHKnlRsAz2
ogeovS6Yr3j+IA2v4rdqZtJafiDv894+yLbUoTDtlxFx0sl6jJ8DSnjUF7Ai
cpsy/S3BFqg8eA8eT28B2kfm4iIbbImRk6I5jJkzeroT2dynnUJ22HWpa4fs
HWuPln6qJ8N6PJi692TFfbWcz95Y9y9y5v4QyyM2oebe4meOd9mtBu1mqtUJ
ySeMhQgFgoVo6RvHRPdExP9ef7b8Sm5mhPFUCFFlxXLliOuPnJju02s9eXTw
+9LnugYSKqldpUqlMRTqMYPaEHgwl2QK2AwYibyeeAxjmWWSuRdWZxlPS7+i
iICb5FQr5KpaYpewE4j6lpce0BKCjnpu3lXOQVj0OEF1G08pKulYzNLg6Kha
INwEW9STpFxw82YfV6FM+Iy+QzdHuS8xuauSIhihDlh1CtOb6qDmhcsex7an
h1YtL840vplfeOm71lZJFLPNZyUzN8a0/HH3FQ5DYjbHHBFLPY3gCTVYww34
RuJV+z8TVRoh6eV6vmQA2lWCNwx31LLyCRC033S9hGSZPNYr1+oO6uvHZuyl
gNiX/zVSA95puzRHVbr+i/7CmATf3oT1HOfMgrdju8umOOTOjHNPuFHQNXSK
vrFtZfOs/Y4FI5w1FZYIwIo/7WPe9bpbf/chKMY7rXsDvM0a8zoKhUgZMCcW
r8YI1czNU1N05nevIjIkxWv0ePz7G04OyZhkB+028v3+Rz3HJ3qmrPx9Bg+X
6VAje3DySh8EV9ip0Dh0KXNyr6z5zNkLurCEXZpDD3h+wCIHqBb1rqDxgby2
7TJDXdtPGPWY7QGkarJ7o/3MnrHoKirWlgvJvsHtBwjQa9si7S2+PgZALNLC
iMLQBI6MWGy2g2VjWVeShodqCOzCB5YLOxTZIhW6LMXyPa/lxYgKOL8lSm+L
hw5FzBkhhiRvCH7ctw2B6T6IxTzE+RfBnNX6Qz8NJbfynzfUbng4/ATpuZSk
5wLn9IoL8mIvUGqOSLZOCI9FzfEuWqlV+O/DvNfzmSIw9o4BEjI45utZEuNx
sF6HBfpyGPrhnpKEMILigCWhA6Z1nZwLEjafun4OhR8G7BhcY0YRgYNmyrJY
0qzLUhStzS20Jm8KQdT+uXkB9Ua66ltEZCe1ihL1bu3Kg/5M06eS0ZPlZTa6
okhv9Yyv735r+oP1Fp4Coqd0QkRsW/n/UPPt2bwVi69P6TTLWezEh5gG6zdg
0P27YxGhz2xWd8mCi9KUHEKPfUm1h4ZHd08hLNRgpc4JbQ6xojDDz6Es5g7c
fs5OlhNys6LDqgu/Q9OKZLld1rI9wnWUBYdVsRExJWefmVZFb6GVxzX8FfBn
ectXsR9JG5g3zS140yObrqbT44N6gIXIreGnMN595Y7AgIUQIdQErYy0Dwf5
BzM9mtZRB2CLdSFe3ezC/muOYNr/SfUHkLaq5WAi5fKloebRetILk4ey3X7Y
4lSRD7peACzwAqzoH03SVMhWEZLVNU5q/jnwxoOW/rHjQeYKsTQgKDv+26af
wKIf7bNh/CZ2VVl9laOWuIvYsFhEvLXhcmSAzLFpiB6Pbx2L83ZfM2YrSqPX
yTLqkIMhH1pol616YKUEnNPyrIRq3s22X+1N5jC6QDc7sSwoKLAS7QatP4Ck
o3tI2v9BD/9e2d9lHGLUNZxzc1UrPWjSOz9mK0W8cDc02gO+M5ioxFIum42h
9ZVCYoJ+5WEwmOexrAdsMaSqahqF7Y4QcF7NwXdUriv1XrUuOnrA7Vs3/q95
Wkfg9wYBhCXFiuBFMHgNb1LF/nhp9dov2KFy75ejuiKsMvVqCCEhGT3+yOhw
85dj5/JkM9rxbYgdPjZxSacyPTLtr4iCyrozRGQZei8aC0R3WdTjgrhpg5ow
KPR5mgvgeXJTQ4noCjrvRNm7XsdeHJ18Fpq/JLxZaw==

`pragma protect end_protected
