// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
pyLL+mFOrl07Wd0UcsHT1id7/zwgrCgc/AN2qGJzm2zwXbRHkRenvy5HiTZRfsIU
b4E5tFv/INFFg7bN5Uvo2vQPyxj2+dUjyecuKOSvS20wmouiTeP7v14BxKYJ01C2
w6icO3swOtcmQ1aAaaT1327smchEz1STY4TUr1pqgmE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8496 )
`pragma protect data_block
yWkJGYDk28kPFKJ3awHAPbeLw0aPeJ/N90EDaYYkcOkjuBgjBzaVyz8i83ltjYCi
aVRsX/aIsgGvS7k3VKy/d3fdcPT8TiHziYT23DZ/s43wwbXD/jdfz3/oApSTEHDQ
8se1+fH1++wZaNMHTy+W561noTFLnZVsUl+31NLVvteAaDqz3i1zVSK45yNBOh4s
xog36TfshnPDoxdGbF5D97BEbPaXPOlNFmyuH1hSrvChprWJYqoVPfiaYVhC4DJT
aaNRhL/SQtpPDUwWwnA4RkxSTAkz36sW6GM6K+Ub33V94+2qjxibqQUnej2jsO3U
Ssox5tEjoS+5Evmnk2jS9w5oIOeNe6atd8Wg4xNerzdOQPeu1klGt2fqRcIm+Q5h
Nu2sXQwWr1YIzP0zwJs+FywhhwvGGzbizUNza4dHbdCfpld+34WtnsT9EQAT5dJo
OS5E1v12Qk5twLFJJWhL+J2OODl5waIF7jmGCwPB7+c62StEY6kvqLIKIYt2UtEG
AeSki6hxZNCThToTg+ko/ZenX4Yjqz8BhiOLQG6/6r8zes+8rYYbd43r176Dj3EA
sgS2lTUKVxctoITzGLNXWIQb1SiLFH9LG/G16gQtwz+DSUeuwb3hFZwdtte8Fh6o
sYUFXK0/jaPtF94aTu1KbHEsMElysD1l7yZpklJoX58hnEOiJZ8aOU3oATs5GHli
sUWqXPQnGBfK6rjqyHHlYnnAwGieZUidNmeCkjJLuqRBEVY9gd/mWpbi/30OoXf5
Hyf4u2r+wVQ2c+MFvLLwB6alQXRw+AQ6mzRpwjm0v5q5ZfI1OocXRSmZi7KilMA1
7JC6XByXV111dL/741rPZZ7W0nE9WbAtpEmOLSXbVgdci06zt7S8yCgk6NKSuQZf
dGds4a4GzDqCIT27fxh3qIfzw4wGdfZwqS1idG9dQDFxQrKBrHk7BsfuUooM6Af9
OTg0LOljxD8aQmjgVY85V+5KzF4HI6SlMfa0DP/s/yPy3o/CSLz3nsx122qnPWAf
3NAKoJDXXBQe9Styvskd+yDQnCFxRgIzdNaC0a7TXjMTK7W/Xp4hGm9SxKap8Mi8
4ELZWFeC8gNnXKxwpZZCYJNyKnZ34HV/eyC/3QdfQwOONawWb8NU+5KL6qk2U5Cp
sXFJ30OFDoxYGu5RpbvLcbxUO/C1PnC3+TBLCA+gPm2Mq0wC2bFV9VB1yw2/a866
6qyl8XSRHpHD/k5OXKubw9JPNdHBWPUrHgGS2bI29MZ3hDJrG6B+Ztv0SvCGH2lT
CZjlJGY0gagTVldq5mYUqa3ZMPucbgom3Y3GGx4/ex3Mg5OzmoidkEni9rnyuuWa
Koo6A6dvox9uzazB5PKppE+dttPBSXglU6+kdUH8xU+IQ57VlyU4u6EZhumCdnE6
CSwZrw9n2+TIf+eOG55lgenFD+nkeZOL4Wdh4dOKxoDFg2GrgOzVAe4IAZHLWikH
miVVTecN7Tma4zS2YEyounurc19k4THIeQTbJhnssNdwcmLOSpb32/OOFSr7wmYI
EU3/koUg02v1clMPzqzXMZBAeTpofzPqWuFvOxTvCYW9rOopSKvgjT0IQ9jd4iHD
EnkNSkbk17vsITrdYdjKq3cp6K2l/K9SnHOk3Xf7oWlkczMZt2YSod3qONVpkqe9
jaHWMNyGYY6q+MwgAq/aH1HVDvXri24KeLIpdD37yqfkImnvKGtbGHVgeKpmOcCv
0Yz2Jy9c5X5b7a1EhiygFsvDtsZ0cw75UGL2PhgJ02gudgUfZPE2sS1+JozAmpBI
BjZ9iolA9XAEHTi+XzbOa5twknVuH9+26oeecdCC0Czv6YEKpUhORfIYT21LrK/+
SdSwYiV3lXiKdLIcrz7RV54lW9DRuM8HQt9PU4dgYT39Z7Vbos0zilAI7P2GeBkR
VSfiT4pzQUMmE8YX61Y3Mmd9URptrSpnbdkyNfpE5lP+ajyUKAGiReqQiCGr0jYn
tQEKO0A3iLbYuUhMyJWs0pyz18MVweagyIhg5xqwTPGeaWX+In5s4gOrZrtz1HR5
I+OrofMcNEVjhNoVKH7r/1anf081cj/sGpWg34FUolVp2xgKWhILgyaabBcJK4rq
LemQ6zxJckx+9Bk3ZSWTGMYqSye4k/zcrv7rRLP3o4KJO/Gbeb/zuzNivFDYSh5d
cOiz4bTIbbetq17A7sD9tU+Vy87d5vlYIHRAgRw1MujQaPEGeHXQ/QmCYYcSmHe3
kr4FCRYMEWaRWK2HANk65LPBQ7sU1aAstRV/OsqxdyCxQytJg+x3n0GH09v+8muo
oyRpwfJjIIDk2a8y7tO2wWOStQ2PsVpIWAEK4xawBVrP1Ep/ACar+B/1lfUIFGVi
3GWFA2Ev8rW5NAfpquRaf5CxCQOAN8LFHtH4jTuqIySbI64cCSaiXGvcV61MY2OA
OKnPghVynPOpq23e6ySpYjvGin6whrk8kbeP/rkVu7Yie/oiKIxNlJF0EkbdnK2T
ZuD4WiGWCqCDfXPuz3K58f0YzpUpkmLWpdXX76x5e278GqBHr+va/ieZkRR5i+0R
xgtzDShP3l3eVRF7p8IBEvqddKDdKL4Q/rSgUQ1b49hhiXWWObZxlxOD4gIsTQJ5
6lucAghByoOLipu/HIU0c4X+8lT7wxPDCapXMXeuvzk2hNtaQQobzg8Om5yBM9rp
N6nvnWbKqSzMLy1c++dzGsBytUYIlP5eE3od+KSjThw400z30pnoBGpNqixEB58L
SlD/A+E7Cc/Or20rvzJ3TIBSdyrp7o4WKodP33iLhJ0cAx3LT5mKNfWkjjI5dokb
XiRrcB5NigBNpgpnl39qU6SD8muVODckYEnITf2T2TXbvRX6L/QPGnx/Uub15Usa
mNk9AUGadqrH2epOQ8u4dhAuEDYsV8iwVbiYkf2st4hZNiNz4tEh+bGKM99lSUqG
ZVliUTddzRBMQYwPhovScQl/8fwds0tBh6Bh4kTb0GQEXC6/MeUhro0p5q9p7dw4
29H1zSnV1FluHuJJEU+42J5YmbEqK7zJVO78AAXa//47wityYApnBIpBeyj0+adD
K6ZDZwl4O/TU4Z2B005/2oKrhD6eIRIaRE93bWzcAxHK3eYUToy30Ct1089atsSu
AZfAgTWaeck+gPBClj/64uBOCWWJHfazoHWtsiw/D7TrBFe85W+ZwCEStrdY4A4P
ZhEUmSXLwGOVsxXmnBbNBVmMk1dHC0xvktX4ppsGVkKRbSU9FmxMzg+xWR/UNBUi
tu2cE2O2fQEng9satQkzGDoWYVh8Cq3NfmBUaYEeVuG3KuCryVs9hffYEwktddYu
oj6Znf6BBsoCIrMtOB/EYjoggv8LYhu1CnlLqmhEykDEIlMKvVHjMZP99BzyxEX7
sU0CwJ/hZMosSMGe7bjU01MvSE3XtiR4CTpPphLVO1PXPGOLZwIuGmULIPDHg2rR
LC5bproJVq0uIxqr21HORXxPUBCEpDc0AzxxIoGRBMa8IQqyk58FWROf2zdcLxHP
K7S1oVOGV0XeMzNcpmmdHJnzYh6AIfOQKKeo+RnDN9H+x5ukAHtuGWqDzW3nRLZn
pIMuvwF18CuB9yA0bdWlgIb6VpMCeRfRIsLKYFQ5hG7dXjZYR6kIUrJMGi+rRpvl
Lt/kwmtMORaFZpJxmqMNhHFVhb4wCpVmwGrbUjiaIIW0po71Jt0Apwp8IaOacM/5
nZbRLosAXAeEP9dqYfLvSuf/3uvu3y+NtKGi8no/m5fWj3r85skMemOH8VSnbbfL
+zlaA23y6pWevGC8phjll5SF0p6/QHI8Yx0tB153oqvKzan4cwDu5/0kiJID6+Zq
TPUkuNi5EIDfn5QvQm5gnPF/e+Kl0BTViHhHEFCW5uUmzoi4WJ+90idEXNpawWXn
hSRHhu/Fk4/Z48+hrWXys7FhsKpu0kK2axWoKqXV6usEyzvSZZY8Mqr7gjbz0Vt7
Sbm8czNMF/5B1eczvHdIdTI68vLKQBbQRabcI3Jcnc7Z/95QyFdyiaTG1bau8AbC
3j/r1M4B/0YmyFh09e/1XcXEjZQNOhr3hZOYbqh174uBpkVY1TWOCjEMsirs8uDd
ptEXjpAD+LEGyy4QVbu8L+B7d4FaHXzvINC1mVVk0JeA2DWJHR9GqIbb0c5rsW6p
z9XmN30O/5Zk3+KdjxxMuwv99SubOZee4EGsDb8dPYX28DVlkPXmKRX7CX82igZw
6MuQhiwZH9QgqzQLr4ns5GRVpLVYEVbam29tZGOAVfzRZgDEXuQhHGlicY1QGPiD
vRFOh4w5r7W8IRH5dh6hivWxvW6hqgs66tJjvdiNSjK49icBkZcQOCfjRxNUkEQi
XbDGiFAgd/DvV8acCREV9JA+GABkNX78/pF8ltFUKkqOR8LleKSElZbtUlT/mO4G
wWjEPBgs9oJzaRS/6P+XNDUTbKcDbzbFWzV2wdc/fuTELlfUr26GKxTVZWKNBqjI
h8MTlScdRwbrrxk/piKfeRE8GGsKXuJg6Z8PeO3b1/XOrwXk0Am3YWz5zfhP4e+W
m4Kr/7eFfhD9K1rWxYl9jHUBYZbKDGixJtJnr/KxsbHICRqPrJLMv9KzyZd14K29
4JDO1vHNW8UMkPg3LVmftyfhE2Rs8K9i37ONzyN+MX0HLki703eX5tzZvHKtej9N
oGz9dNAA+rDiSDciIhn7zw4MsHHGBhCAx8CFEHEwSAvOeEvyIqADVCAYOdCRIRz1
/g4E8owNcQ5S3fU0NKk9F8VL3uw1V76Uq0S55N6tUkk3Wa0/fMb5gm2v7A2/Xt8a
4GcsJszKWlhGaUi6yeFy+AtWykAAfzKRo2mgmNTVriZzhPdwJNAMiiml0g2AOuDN
Qr149mPNtntgC4Mo5S60tYqr2W0IpTcoIGgLZLXDss7jQfrcPqbM4qnKByhf4taJ
9IFJD2tvR6lhKaueRGN9lP1SIO+KPnrc2FvQ0pLq12R8ZxLPgvEihNewAke1DDEU
nsMabemY+MJ9BXjoyMnPuWRe0zdvDvEkPFzEjCyXLbx9gxaVt3yZWG5b3+/p0FdQ
zGUsNN5HJyQjkGFwOGYL1Q04YlwrrBF+ULp+SyvcEZ7WIcWlQ7nLfZEWGkXs36xK
B7dOvsmwztuI68jxqSqOb+DNlHLxPjZG+UEJ0gE2njrbRBUvmcZYAiKQtuo6a1z+
aVObEsHRvtUK2o8Q+iT7L+zhQMFYROMeqP8cJ0kQJpWX8af60Vt/UmJ5TnfLz2+c
APapK5SENpwzx8SwLspRed9+6vFn1qyRKl1WoM6j2Zfz9KvHkhvUlduz6tmRX6ov
wCEfPXm1QRHUhimso+WYETZdvq8BND6Ediz3TRsLVVERn6EAII8omkkpZjqRKStD
uEtsEtM65UhiBtEfm6qGsgR+/ZKFW6mGKgHbETQw4BLcBckakTlYdzKT72c37W/n
EnB30+cgQRw0rX+cLFXKrX8y8DJT3ebI+kU4N92jYGklJd7l1zXqor7mb+1HSX4F
Bgn7oT2QSU4rHNmsV+3POafhodUyCeZwqW7ZtYIzlcP+XRBzog0e9/C7UkNJMzo0
j6WHbHapNOUTWGYDqAU5M3Sd3la7Grh5DdwmrnUNX26c8TKp8RRHdYaDtJHzmbrU
vaaAP+PBMkbJgYP6pUnzoAcbzQgSW6bxHLBhZ1ny19YUxwKbWl0VnXJg08Q5Yo4R
yvWPrgkndbxHqD3IkMMarzGakjE2Qz5+Ji8Ert1k6CMkiUQn+rsGJL+7oubxkWJC
EjGE/D05iNwJk+bHLyjMFAVWVNcxHq5VC0n52/3/433CJoLymTCLi1r+l67wCvnh
cu7GwJK08h73r6L2HRn+hVLvkUPoasTkC8Zf8TYRLZWZiDOgl3K+JvObOVkiQk+z
D6NjyjsjZhX3JMlNvUCLCLvL3xugac6qHdl+m16MFtpdKDeQSBCuzXjf4Tn0QQgA
/jpUkazMMYyqSfKgQZB7n5Naf4j4k5OtIBOQx6Z1SRuveT8Yv66YYPOkR/vQyuAH
mdmpwX+peiUbvm5Hfwzqk1QdB1CikxGk4wBShXl0DdeiB9+LUN/dogTU91Tt47eR
yZ9r+ZJ/9Y4dcF83A9YI2LT3vHZ/daoue22qL7/KAVXLAE+PAJQLlE//trvOEoRn
6pwhLUKt4S0b0wh2dPKg71VzLLRMuu6KPKKtfiFbRwRCtnM9zzlDSkTBz3jBNoxq
4UZWNRK7Vr/apUb+OGAF1XF0pU9NSzmH1aBRDp5tNy/XvqoYt006iFzeJIidLgLB
hsrvHHyxKKu3ZDrW5NN7NRMSpW4xsMKGAmyRpoi55w2YhzQjzs1H3TOQdWqEpMPe
J2P615GBVFssdID36gTk2V2QSA2VpbsXxe7BniTmdZM8yPxzzyW8fzccJ2tJ2lnJ
biQEiCjgPKqNojWOAtnotcd4weXJMdatCvyyayJsGyNXP2pZty7Xz7ksg/V3Oazs
UbrULmarSGSyjjUh4IwbWT/r0u7qW8yD/xET3dLHOrVKFj/ZfswWComhUtBDr6hh
7RQa8VxqqEzC81PYM+mPxHLMAc1StrMMRPAAtxfMn1M3BDu7IzTiy7JTezFBaSUt
3QW5DKjxbS4nKT/RQ+uqlZkpfLO6SsGIZgZMVDLEJaD9xL0vNtc389Px96VNlzhc
+NQL8Jvns+LJ0t48PO0LAXffTAb1crACE8irFg73IE5Vptsv0IFedwvSK4cMw9JB
dIckc0VMMMQvCJqMpgs8Zx/xsCckGdm1LJ9+IrI3a5lntjSC2UrQ3eT32TJoDDt+
VYRbFs4BXEy81ZZplCJ5mR24/GxxLS4zpIzsLVfcC2gvumnJDRIV3eTe/+CPjDnj
94qmf7naEJsRWNKZaLATYUnwvsUWsT/wWBP/uXmUWmXjhShDq04E/Ta+D7eQVc6I
KIbvPoGPT6nJug9NVr48M1S4PreSaUKYF1qNXgAbfEKEJU215+Gte6QoE5kquOY8
eYkNifB1wsaQbayygZMA0rdhUFBX1Bf5OBVdykXLfZU7SGsCufHb8hb/pR4yofIu
ecznp+45/RKc8P75PF4y8VuPO5bcKmHJqsFVLAMJWYlht4zukzFAwd7/OWdJftcQ
9Eil3S58eZU1u4A+Lp7VNJlRXYeBxw43AR0QPU5GI4bSJEQdaydAQGgv+zYfeoRj
dHWxqycQw/RMJHmbPcYuQ7i318aUKvWAcQYKseqyaEgl5WlBz0zPIxdj9cB68BBH
wmAX70CjnCWSNeH8ZN1tc3LOTkfjMzu0rAlo972tsyNYKwWg7gmX2a5CzV2/rTW9
6RVsHNxdCbI8BHqDjPu1BGr7YPshXRDJY9iY8EgMDA7P1c+GczGVAilLM8wS/llQ
WNsxieJ9MyTAfXd0rizavaCOLrLic3fIWuNdF4NzGJaHakHHmOQCVlGerSr47rgM
GKZfubljABWJ9EVZa8FTdyUrS0fkSIXsPQV/rG8U4K5nUcRmJaEreLovKa36KpMU
ZXJfDfq+vdYMVWoCANYcuQx89Ypn8LUr34eYO7lMgCQR95pt2uP8uhmYemGMP+Br
7+/bXp8YzI3f48muu95kUElvVgECzARXjMuOiSZD65K6HXs/qSpRPPceoY279brq
dujZpFGv2AqOYMq6U8BymjH3stXDfgfdOzBRv2UIUw3ltfWgg/Q79qBNEpVnnJ4g
S5GwCUHrPz1dOXSBO8VL93kUZnyEifc82wp0lLEkPlOb3/ELpGSMvadtVDbDyeDT
Fn03xCymAt76w2gN/62A5LGKL98MB1bOsbybPz1dwbzVtIVaCwcGQx6goVm43lIM
vjgtiE0awVBWocH8Ak58NROlH/Bu3gqikRjNmLSQOFTZYNRWDDD+iTAoAxTrRviX
5Fom+Ku+HLN+3AYBiqzoFjCRN888DTqffn39rV1qWy/gTjdmRCcm4aviRmzjuydZ
gjUmiJvToLsWzakNYI4xWZyIvhN0Ywr05EgmuCo9WVDaml+r5UeFVcO8/waQ+Q/f
lEgediatTTfVAprUm+N2a7FTUB/ag5FifXmYbzWHOYjbdbOtkgF7swzyfokmML71
Uk10pXJsmh4fGzyFJoWUk8T8c5G++FhqePfzYGjsx9j5SkGLCk6rzGW4EFe1kKCo
71OOJd6ycQg8YyUYtxWYoNtWD//RVbNWbbJ3g3veg28EYkMR4xirXGb6b99Lk0+7
+WiGFuyhKwY+iztSOmQFo17PhDVdgO7vcganjeg1Wh1HcEaQX31TGBH6Yw6wHSuk
3uKRtBeurl+CX6tl7siANe3mSr0IX0GdkEK73pXwEauZ4V4e0PmSR58CfZZUCFUU
wcXntzUR+PzO92+n4x9fjhfdxKih52u/vzpqKP5UsX+qUjOkSL/WTvLY97/9MKp7
21j8Djxca8m+GMxDPsVrLQc4OpNL3MkkTAmAxIsJdFQ2gwpyfv1BYX5JYPXUX1Fo
NVGMgfxCTMwTaNBMHXtxZxANYLQE2fELuJ0O+nVqGM0ZpUBKLW2vaO3z1/6sYcxd
KPUbEvmUrtJUWRZ8is8eZESwcuomsqNJS3w9I+m/w9oUSbamepLp4CoeWbBiQ5lw
DScp06PiI3QCvT5BVY9rdLtbiktppvDE+XHQ2xHw8g+/A/TSIWPJmxU07zNNolIP
3bKUkWECLCpJp9pSKMuDWjy3Hk/rFmTls7MlR8V8trRqvTycl3sPKBf8Sd1wH4jV
54t6uK0wATkH/E+RQP/XrGOTGkgWL8Dts0RUW0PPgP6gcXRJhawET4jwGdqxsHIg
IRSc8e0eUZz23ZAkLpXpKnhsAlEtUriRP2EUExWtzNyOdvtW0zi4+LeLLRDNQ0z9
6Fm1joKedJsRVzs7CX7waLt/oWXySGSQGazTkX0ZMhp9NKNfO42FG9LnqXI7doxF
V8F8+Sq5MY3AXB+linkrGe6cRSMYDYlViSNT03j9VbcQYQzfpp41AEma2t8N7U+G
5iN8T5ZkAH2THn6r8IwOw1hnulcrDv+h+bAUfRidkLm+ONj1kPO/ft64+/FNBd9p
Ma10Qm8LFwhSp9jD9haNEIgVPozfKSD87Tayj0EaDdqKXImN1XRGLIABi/lYY8r7
AdI39AbAP/dyCZC6tHM9ddWXJ/dYAZPbkELrDdDzxI22+sksh6nKbZ+Fp5Jv7aXZ
mkPGAHlXXLHkIc/d3MJpljvmQ5J6X3ffWe0RP9v/+jFgurHYbuNoAOCD2WRhoiub
pF0XO6wKf8TekDF9qukiL5D8kjgk6plBPAt4wYFvVAa3Rtf7T0t9+hyt9hauVVG0
xuATuB1TEgeGZgwiGnnSdtbOLK0rmWf2Ml/r+SXktQppdNf77n5uAem2Gu+fR5Cw
l0F4AN7JCPDw/8yqKmoSTF3UMy/KKg1qVQB3SKCAXaOuD25hX5L9zijK8f+xEaqm
rwjMbFPF7NcY6yofAAfiI4nLMDe4ZK3XinHPyFDFhWwr8YQWqzzMP3uV5dk8mopa
iOgeHsp3bXYgM2vj7aNGK8mimYwHcS+D9XhCh5MjGNmO9qIi/eL9SHSb70aqV6P2
UujVGS5O4ADPffotRoo9cFSCKFaj8Lf5JvIZFHTs/V0ZYgA44dVqoWNqsm2TG31r
Ip+sUh5aiJF20p7Y7pY62GJBC8E0KkjyQ7FYSCuLNETw47DLgexcQdH24zBWoLl0
9bDomzqyNgYdLFiI86lxAGDW8Oj8DENHPJHPe8Cf1A1ePCChKbrW6QhCWwQ4ytQe
AkfBsHiexqjISrY20f/X6e37tM+akBCmzGNQMaVN+qoqizgWYOQ/cJq6KNmOjAdC
LmuE/PuvegC/DOkw4m+WaTGSHeQ3vZ/SpzEEnKci3az3p/gKx2hu/yGx5k9uEQAR
TBiFjhvcKR5T7UzHuZsU1ed8Zu8p2OVoMibAX//9T3171qAu7yHVnhuXVCOSWFqL
qQMqHZlepFZW0hTthjmiYDiJsC0VyIp4HM98mnOvAaA+KC61tXVb/Wh1tIcYzsuI
ORnPJ/oz49LuG2RluQHHn0aL7BLKawFp6rA0KtJkg56/aSjFlqxH/IpiQONPWZrD
m64it22lk6py6Any4gdg4c8eHUB47GVz40Cv9oemD63DueM9tHkHdFWWAKx+nWJ7
m49TxsHL7xsLfFhje8KPta6QK3kt2/1Fzn+T7t8mhYpnu4BtyPiCvvqGTz9KmsHd
tqpEw9Zw2SxaIpNs/m25EgjHhJgxBINOdolQzRVk1J+ciaoaMudCkdBtPyS3dA6P
ZLdJFdcOmCHR510O7af0oPASkKAaK/ggt9t75ltR6q1C5nbZH7X0Ux0xAlWjAcdD
2t3VmOeKFInzS5vRRWmd4QxD+ATjm1eXR3tUZUIkKKL23QEdiG8rXT5Vv2bDVkKc
UVpQn2JXpM2A3rNmjTBop+jyrSSLBOmBy3160MQ88UxYMDM6CGb079Ta8YFIfaDw
c/Y4TLt5BDAl80sXc62BvdC1p0NOMU2AiD+6yHFRAqd92tf6zuDzXgsPSA5n1hMS
yHR5QDQpKncrLWVb3sa6JgpEXBo8DNrzo+dgqBPey6ZCiEZHjW5bw+IB++em474e
AMwVWgDQuSXOzB85mXUKRefbYMVWvI0h6p4S1uwky+quq+SaK0sORj96uN2Kj6UH
Lwl2Aax+ctVmFCnZRrhqvVfklhilbDsyIiFh6HovsuWnHZ5BSzZXVHRvU1dFkao0
YpPFo4Sa7OwsBziAZ3HAYam2V537b/HTP95gQEhyuqt6uoVHvYGGRTkdNX+cD4Nl
XSgI5JoI7/HLOUk7xm2dzj7dxMNdh/UBe3tCRUkqNXwd9HrYh784CSqAx87Bcgp8
DVZ52goLaSzLXmQq3wJin5GxMInILvSI+NvU2lWav2iBHdRObXqZSz8QBbt9gEaQ
js5TXVz/nUO/M3bl6GeSdRprZeaZjnqtbIWOsa+SaaGA6ZJjy+rbva51uQH9Ep5s
uVREscnZQmn8zqOuz5XwiYjZBU6kVYwzB9KRwxlroJA6HDH471F6TkdcsLd6kIBQ
ETZzMDjxFjVltX3cc2wEYde4oeBZAQBvbxempNVF4+Yu0LlBtGmDp1NX/QnMmrx7
U3/FUdVgj62QLO2vEvb8SOuHcsrkBnpktpEWrgcGaLNQhaA/NUMhl2ZUFCutv2Bg
a+CpxL3QKPoAtFqJdAzOFqOx21KxE3WT+JLkhypNvExKNxGe7Bi72I402S2O6g2e
6fNdWPp+T4tVUDz1C6gLPUGrSSCUw0d5pCMi8ybMw5WXcYuQrjh2UhZ8TmpY6fji
mEXgYrkz/36CTy8QxtLpzxilWRbc7q4300etnebUt+nHPssapNtM+BePdLhIkpRM

`pragma protect end_protected
