// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
lF+gRXOvkxR5P36EwIxKJEykpoqp3RsM6ASDPHiSPPhVOXrsOW2EYLQ9ClzUxOu9
SQbAh0xyOEegwkloTY4G9lR4u64U+aV+FF5p9jIv9hAH4mkREcxJOHkGPsjGrfnP
ZvD+hSJWjr2fKhIy5AQkSplcBBhj9eUeXdwZ2e5pmBhBG5WQwX/RoQ==
//pragma protect end_key_block
//pragma protect digest_block
dKSutBR1OFW4EoLgt+OMtzfZBis=
//pragma protect end_digest_block
//pragma protect data_block
LzcPeu5n4M4J+hCCeb+9V5mmR3XVgyuaNNvDsIA79Emvd5h3qewzLJY0w2qDJ08V
UVh+pqY2GlKuyhEpQoUdtAVnP4t3kOs/Tq91AVjL/1Kp1A9u3w+yAfzG90tPHcr+
5I1K6W9vGr/Ym6NlITTTAKKnIYAQ1AZ34PpGuzRlQJF4EpLXgGsN03Aygw/L22//
iwlFyRJGWFWdAh6HK7MyWtamW4wk9trzlrcr4PLQ0W7WIKz/716NG6blqMcAKMp0
l8uIDFmBnnZITd7Dmg4ZqSKYAyDHhYiXtRvmmMDpqpk9UbnKSEi1KrYD9yNXC94L
znB31p7bByKIsx2tTvlWxDGGMNHVzMJewTiY3pKp5VQM/vm0QP/XMbDfA15HGf6R
SsJbajCa666lRnsJHXK57P31xqjsa1YhXZVPT8Jf8xqyUwOZSyNtB6guj+2WoWqN
5Kj8GWUJPVr6uQq2tLp3Bv5basvXMPWzdhNdW2abeOLS02GQ8zo6Mo4x1bTARqwl
vcbgpmJc8Jc4O6n13l7PlF/6oQyB87VS//X5fGuuKsn7JX0A7DO3d22DRjAMIMDu
h5srBBaasx1tYXiYBCOhecsqdOM5wwFDgRHzwkLR9Nv6M6SOyoFoK1bFlRxsOkPk
Pi45a5/QuZ4+Pvu+mTiBsZsCpB+tsIH51o5GBYHWl/PZC01czzkvL3dAtczCpKTz
tbJAqDYleX5NxTIUKFO1b4ulCGEouwrCnbSTo3D5Ql8bGXUqjSecJR3avE1CzLN2
WaW6M/sgvfe3aYkVcpaPUeSB7VtLZRbsmzYG2YcaTFCTqjXWMtXfrfq7WiYw7/s1
aGmH2YkOYz1Q4HZDiHPKfPxtm9YRRQqYblRQYiRtYYXBPhe0bAICXhsEnGxUF8wV
45TJ6Cxs8PYlmQGYjWAqbueryllZunAlqpr8movnkVTkuqh4qxvhr0JE1uAfH5Od
vUVMEl2Dh6WUOUe/vE/zySH7wcPQUHyuFz+nq56YnotgBu/dcR6+ZBCirZIRAnoS
kSqhljO4YKLfFl4HSbLe+FobOyRUYbBtYN53Np8B5eKYi64NCL8jvYVuXVNIij8j
AMSAb50J1tgGdg9qHGDo/ThQD3ePtIiqwTnPgzWIWrpAGd+ju/T/02WMJZvbOGe0
3kcIdipdgQ90KVXDp8RX5Guw8DmH6wJ0CmWc/ip8J633olzKgwyqP237zTlM6hDi
rAnT8IXhjzN48XmWy6yIrRRKYvM0X8eUgXGSwWaPnRMhZy1YSNHVOXgZQeZh/ycn
tBin6KPqdoarCjAMY/Jk0ZNwKtT/AA7XRwooIgK7HSW3xhkmOJiPbPKKx9SJMAN0
oFAs7qCEsJc4XojdnYfKCc6u88N55KVggeVRv7gvWddJbAnb4ZwAxa0Ap/gt0rj/
F5rabJi2aF6j0kJIWf9Z6P2238MOrR3OCg+c2/EVPX0UWCIxY0PCvRYx9ZOJmrJI
6S9WXjoiv69wybiNL0yQS4iZO5pK31IS17hgraJN6MtEgGO+yLYEbawRcWCsR0HO
QRQ2bwviu5nqO0/KcZ/qk3BJ0Z9t4J0FeeI15F9p0Aet/apOWm95n6b4vvLbVJYj
SlH1CuPi+svh9aEzD3p/dQJKvGfXVUeeEIbhtBfpUB2TK6uQTosIemMOA034yLQA
I0gTmL/FZ+zlsdqKlCRi6pf2Z4muFNpvR9rpiuNamSZGUYadoc2iFi/ZA8ms1pgl
2Bt2SYRtN6BUUrHj+YUR2lNzTMRrevVNx0XvtutKw0TImQgcDvfsm3JEFy9rdCem
dt/1/7tbsR+oGPAaIFXeMfBk441ohixjf1H/hFAszxtLZrXvs/gZNE2FgzH7y69U
Xn04nn930OOCWYFn3na/FdKO8Qzd4DkuULDdVTds7WvkBjvoNG/nwZDGhWryvTop
7Yg5SuinVSoKcZF5Y/0pkUzDPPIIbHWBjt1LxBCrv5sOdnyw3zElWWb9fhbAUdlq
bWHZHaFEk/VF08gNZnNAzjInYFWOOrTWK4V6aQqF9QV5ubpnbYn45FnAcjQvXA1D
9Ev6RB7Zz/UsJFEfSjx6ag7mO2s53cORLMy+aDN6HdpaGgBnArXlJsh3QT9/iiHw
ih0zL7ngNroUUxq3//rku669zulMCmr8EBh1OTdDtDgQ1JTRVLdD77jX7YU1Ca34
3lST6Dsy289UkOmlL9ahm4gHkBmZzrorDhFLPUkGMhojD/QzqTKOxcm5v5RjmHoO
YKMg14/bsKxNF3iIP+rhC4ca0QccrkKeh5jpKqGCrzWFJ12kvoKrgtSqXgpj9QYw
ohb/dvfpOGOxDNGlv+SzXf2SaXeyKWbKkHyeTFzpUwEoR9x0uwQ2qCld1EQC5eNw
hrjqkZs/It9nwxj5IgFRjr48l6nrHIFtbD59n9YbnaYTHLE0sGr/M4pu9+Vr93cO
eAkRN4qntKdpGq5A27YIL0B1E7H+za4pJiXxYw5c8ey+6D9fDw5X6p9CAbLMvUZE
4KF9QX34EaPK7MP5WX7HT8yKT7MB3wtFZPgWgEQ+0wXppIlsUFHSFHGdmtTQbLdK
rThRpkW1M7OIysyC4/JYf/IrnjYfawBoHq5kIeVX3Rl/KJGafWp3bqPTM6b2kGGg
ooWYJHMRlowXYhJe61nN9Ch+y4XpcZ06kpZc4qeK25AhpAFmqHtf5yLBkkn7MyFf
KtB/reYbbxdcrW3qbdFhavakhAPZ7mVSfU6iea7++v135BMq71rg++OotkBt/YeK
G7M0K0Z8XhSVeYJNw6GJc7bObDQvc8CBsLvZ+r1QnhYIU/GaH1IP+JvBbHz1hgCN
YTNyq8Dqq4Kw68G3RF2MlJ4LdzRygSO8l/gReOob0GMnCs/V02N7u+jkfKAEl4VM
Xv/uew3NVf8VEJjUzOndrIUbnMCTdUiCmaQjQOX0cuEOxTkJDah5ib1Q6gXHgTGT
Kbey7l/gFF/ctAKGOW1gS+anAwlRAj6d0Cmh3Hv1anqhccACQ6xPL/nWPmVQHtqY
SyAruOqXN/frcFi7ltH6z6Rfr+o0oPcFKSxA2qK/76NZI3gGOFTvGAh6EMWYhapH
nL50ffe2SS2i2N49a8VWEEDgdqlQ3LdDJ2WKkuIcG0n6IvwPWlyPMU3lanaB1/CW
lW82ly8f57L7xrtWM38d3qOZTUmnTqdKZ2vrlJjS7ywSIkjAb0LBbria+0Q+vMcZ
p29WlE66ZtUtbx1CBGtfJJCCMxDCedngeRKaWWSWnSXFzHBqjc/ahTu0N5k5Yr5E
cly/kbJWlDRQ/xqDIHvOrXhJbZy4tdvP6knfTIWpv7W0esqVEF4eblv8+zDW32Jj
mUCpBxcZbh9BM9qgSx4BaHdPTat+3C7WwuMeQEcQJA3ftcA6T2TAPIozxh11Qal7
0/3rq4GWk39sdioEhj9QV1Hnz8BlLSqefxMMuAGcRIvGEvlDYWngW8fHpIXoul/f
VYtPuCw7xN12AiYLmb/mtnKPy6aNT2Er8+xaygevaLBxW0Tbmyz9IkLyQ6wmdoDc
UjpeVNSbVgjIe0dOnMpLtAS4Y11+Oupa8/6eP3qxLTJLVYBUe9oTUYEs6qW0pYMF
6YtD6jDGF1RiM/r3wozmmWoF/Z1XaU61r+m/rQ/fF6/IdiHRKnQ4T/mjSlekKMOV
+1Si+FBdUGsQOJvc4BL+EqjjuHdAs6J1ZP3JQr8n2V45RktQBj2ltJh5f8zrmqpU
deDXLxBVFebI6Bizgiy004BYSh4nF/p7fd/1Cq8/ET2JmIO7WKBIRw7i9UT1i/bj
Mtupehb5zLQbqCGHlLTP9fxE2iwbQ4hENUP+FyGKph8b9ZE55bnz3BkNLCkeGhk+
htjcDzJiqHfrLcAAxBMYkaQALMpU0DqedUCveJLEiOUK0xaFidB34CgpE7aIuP1M
t25eE35Q++vP4efjCONG660ntEF/ClcI+uBeVZoEnRjtXRlNFIgffyBswuDcXkw8
CT6peJzeIKHW2flevuHuhf6gzOIdoiiTehiGglelPRIRZsK8JERoxoSjiy8Q7dU7
Klm6hTX0OppFZPE2FSnFMwXJZ9y3BbpZW1NMwnw54xcakTlUxG+Flyx9zK2i/XUr
RerRqdwhpZmRHT7eEN+xZ+jdFM+Vo8fJ6b0UIxsm795YONNAUoW+RSZgMNa7y2UH
nSsSKuApcgPQSoOVL8KVnHwbHyuo6flSoU1IyL52Nn8khVzcNbG+9cMBpxH5TBHs
3AtCOcKVj02kjstb8g8bYbq+lcYTKPRZSlcGiTqmkuE+cK3eQdCjx0jFtqP5o+BT
gnsbKsFX/ssEt1zQ2BgkjyZZ7SylxiTUwB090xUza6q4scR+SRUvAGK8pstBBS6F
UvW8xYJCzVb4AGWoVCNwQXNYpUJDTFwo+mzA5/V9l2DUkcBkRPx0LIlJSF+79MFy
If8JZkkZNp3pDgw013/5Dt/fS6ZsKta77FcUdGpCNdVOJuj1l7rc48svgEDbtxZI
dQndSUlfmYhHdTubPar+mUe+9oGd67G1y9aRmErrwbPSvq1Du7/q8W1950kiSlst
1I8zdytQDtlQfTT7JhG+aRqbYsp2CEXpvVuB6cHmbi8hx6UxwhOnO4sCcKuhcbtH
Ba2H+CGhZzbznT5/XamJvmVWAm8oQePQQVtWcWbZhk5WQvj3r8M35enfEFwAaekk
Ema9N+7ArMWml1CaR/iKLqz39ohDSrHvW5eTItjUI5yaVtiPAKRSVw0xzN0YUNiQ
YJXFjHTBxjfS2yxE0sTp/YCF0C/m6y45bmeHvN6SJKo3n+MgRv33WDm/mqUWpCQI
J5l8tdMIVdexE8y0/035ksim950AljBobmU//S31IaKrOawVdW5uxOIZTbg9rAwj
yFsGW3zUXdGZGbyPTkj+O1w307jLoEqjM98nu12sBqES0tU6nLYr/WwS02fpKdfn
pHTEfBw3/y2Wx4R2HhbPHwaUpCoe7qumlWVXDn4F7JeqDjO5+MLr3qR2mvfJsA1W
osbflvH4Plmwr6Or90zmFeXcG7olkI+xOYZWIb1dNuPmffQjIHCtg18+FjHhhRBe
/ZnTpvvk5BB72G6KA+nUYXXjZA7Yh6eSvwGloASrmek9z6d582brOAQpOSjQQUTI
l5yDtlBSMZM5+cJeMyHvfn3xZ2yKRcs+ecc1k0drumEkROFSv6FzY1+ASZ8WMK6T
h3fcEysUpAUbz2w+ZyLJ1L6ics7DO8ecyyHO8d16qL8OFggmedouZ7izkmyKXxo/
p9cjwLODC86L2KA2JwTi5WAM1HFG9v2+LBmwXQbP4E9z2PKKpNgVxDo4mi4Ca9Z6
6b/xlOnZdkanRpaky+OHGd1ZT73LKXqgdeT8U2UvVa03y9WTzPJuCuBGIudmB/qF
GCqPsD8TT9vylE2h9vGbdCY6pTAJK9f3M5hcSyOeo08RUkiYYglWEeI9jISKjVZw
e7DYkpc6eKFNPKodHSF47BrQ4+QWeoQ+oZlGst38kYCda9AnaVSRIuiPTfLr2LZc
f018+3ckgddKWnohhzhmRdrOfJAJIuJUHbfiJISkiEJF9jW2PT1k0m16r9ZE/+nB
uTk6apr5Mjzw0JvmoWjxFcQrxOqVA2j26paBp4HeEqQMM7BEYOfhElNP/Wr4/vFY
CKBuL+KaAA2xBINkxuuQUXiuogCU1APzdVv2BQ4pnEF9LynZO3uGBbJdRBytXFDD
ED6oPfrxdhGO6FnLqTMAf1WMfO9Yje74rkL4Oog94IfK/vTJYUOhMaJmB8dq06pI
Nq9uNnD3uYs8G6WGakvNOGQv3OMZ65dTx2FlCHooesgJzPxALBisSVH+dcpTmhXV
TxxsM9DWEXm1J7Ql82cjfZlM0uTQHMwDjm58UzkdcC1EEdblhLJUB2KGxRzW4UUI
+8S5rHDOmvLs56Z8EIJboHyABZ+dBd1lq6TLWaY0ETAHyB3dWD6hi/qrjp5HCajj
IuJ6QkfUQqCBlR7BQkrpUYvzCeptCnc+P8dhmT7Wx5oeQ+4H5qRWbtfeyWMgxuS/
9ot7kryo/Vs/VheCTwXuM+ZDRIssKc4yKgwLk7N8eV4wAhYJj1za7xWkzlDVkmk9
B9YeYPm6xM1chCHqXVQT8Iw4WFA50Z+uFpB9BZ2MM7qJYO5FT3C9SOUIBHQeB161
Ce2w4ZkC3UqPACPC1GQSaAX30SVnt+UvMD0JYu5Md8l4Zio5nhHKkUNZF/gTm1kK
/SBOEINd7VXsZAqvlqgYfRVpU8P9RRZ/cCBoNt8ppsRb7LH2Q5iN6bg1HFNThe/L
vqN4XJF6f3HViAqQIzb3qeyFy8apNiDMWY5xvM47LE6y9iK2TzaYljx58MKb/uzW
3IIQcCXbHxVKWlochUrHdiq+BzLuySnPuOh9N4kjQpG9Q+YFFcVaSlvEZDo+etDZ
EnDpEL8UEnPIpL7UygP9vMD4KGYYbhRXObVN4LI5IXp4zTOEickHQhIMmltz1QXz
bKe9AC0BH0aiGQnaa18YBg1SP0ZD/IB++Cj72GoZBhzSK9WajCTpNvbvkLM/nxsu
ZNuOUI1+bkQ+nAIXU7sIvTfE2zitfHiLxVM2322lP5fTfhlBd7DmDJ+F+7LNmJ0z
VF5EP8aezOXZT0YmQQR1kwmnUXRpwkdz/ttrrODErapbxpdcBpRzWV3cfmJCbfgi
4bDXpu6H1en7wKH69qYZyiA9/LbsLCkDRAigeD3lIjTUMIu8vsNTW/IfP7jiPjm6
tOm2latgg0a0+FLTIfZ9u1YrYxBkaN37AsWxHpjVIZYCZoFPl6M9XedzDqKhQQLm
UFR9g28bQx+0tZipahaTTCHNGadsYjpVzFDPZLK3g9c5d6pVjfAMaNqI3VTfbp+6
7N58M/MJf1wU8DM+2hjyd2RqQzEYJIJ3K920OTF/q8LaAeGB6mkaRqTmrjHhqx7d
UCr+v9M1+xwgUuIH9VM8fWUoGhGdRXSFEgm/b+2K9r+t2AjJ27n+I5eB7ucGkaRC
ltXEq7f7iBsfI+5zhgmNBnRWwgV7gW4+ZSxjwYHkrc2ozxGArwyLbgb6T6GvttTe
4wKEJ1+ppfsNaARxOgAySEaa/u1UVHL1Ver/IRQazpRAYaxlNv2J5DSz/iDIFjhA
xcGvlqIAyzs6ys8mZIYccyiqGX7NK1vcDxzJE5LlLWj2NqUcWZI1JCZ9ueHiH/e0
tHp2Y7fjtrJx0pqF8BjCV3Kne/UsZSclxFAPCU++NmDTv1iLFFPD4HIQ3OnzjbOU
fb8Hzn+FTOdIyQQe1sTpL8ddEqHQNw7xcXkuo+wDoBpCyUNseiDhH7wfgnh6GWZO
tRcnjtj08x51Bp/FugnohjlsPuvr6N7AuiUAE46bk5guQ1xqOdB2ZE+GSSSOtko/
6rHZQ7ZOtcwigHiWCdZrSSDeE0OPl1geDgjSWrCRrwQ8hhO+Elc2umDZRr6AfYg/
jK2qICcYDCdLJ+lCp+cFYjpiBzO2lhJdhM+L2h3rfRTWZFCBr1s6qS7I2TD0NuX7
3Nd2EEalVojxfcp2wHLX0acRp1y4pqIPk0fvsMTZm3bSYn/QRDPhMzBje3hjpTSc
wr29+gFP9jHFPvKs074rfKgG5ED1D41fxXi9PttwkDQ=
//pragma protect end_data_block
//pragma protect digest_block
QY3Hb9qBmV6AMD/qmJgoT1RU5PQ=
//pragma protect end_digest_block
//pragma protect end_protected
