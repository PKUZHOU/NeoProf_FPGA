`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
P7IpxIHEnDTFeh4P/Yn0wAek6SfgbXFxyczpZzIKleev2cI5O0rS0oRqlkWe09+B
DsnRfWwKzMv0xAHV4oC9Z0flolmMI37U2QIFtg/P+hwKFIUhBcsFdBhN2XxSyedX
k8jk6swYNeGUvmfnzRr+AvkDPz7iDIFKLukjY4wsHTM=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 8592), data_block
OwXKkSF6GJ5lVi6ZhkVkgXPyVV668Uu0FSBF/IJwGfQV+sIB8bpm7g17JLWoUYLk
v29SAsfMReRHwaTPfebXvlpzy7Bc7HI4NQxrXuH/gD47dTTo5OKvf36Lzj15t3ob
iPGRihVGGl1Yr/LMwSv9ZM5Is8atKgJ/Kkth1H9polhEb/oVsijYMJ3GMYbTyejl
bFEDu/YObaFuGFom7CL1b0YbeACYOSntfsAi1Cx6ful/5skgaSSPFg+M4xfsiKr1
YpfXuoDXVKc10q9omHjaUQkJhp5ASPCvvk0xxl9LOoS5oEY4ZJnNi9FZsddKoOgr
AtqsUp4nCFtpCd6K3+vmzsskL0JlgItKfdqPXAxiXvUoonA5wyKyHMdwwpyEssuM
+++qnbFXSdll62xI2WvRiEWRXpsuzNTuk9hs57s1Wndpziy1PsM26j/0f2XooCK4
vTAa7Sp2mtQJvqCD1xap0sMSdLfEBNOnT7yfMC9OKP3NJxaKRephbwgzkaZbLmxf
UXRW6AETcKGyk5SY5t9y1nvtLuPyw36MDvIl/HaI0VIaM8EwzFtil3smDGMK0+FE
K7XvVNPCDekXBc98yh2l1jztY9w1mAvE63TAwol/q2XTarlqcAPLpUsXjMNPB95O
/L5lgL38LiGwAA+9cOp2+TQqHmUPsB5CRO18gmbVapzV/oU76qYc2KY86bTpye4i
0HN7AWogeoVyoqfU8f0lOCuuQdU7zhFAaLZi+5GI/8cwdDu+JLP5Z0hPd5tMnBz9
SBqjzf+I7xx495M3ej+eMeiQJI4Fb1vqhdPb2Unlw58HSY5prHSo7O/z5oq6N1Ws
e4+FmkWy4054lDymg1L7NMcFcZQNJYCqn0X8VWfzJ3mcu8BAyHYSHkRMS5jLvPz4
BUiq361w/DpJo7aM/p2OkpkE052FL0XMix6MtmsAwSmBvE+hnM8fA78kk6G1LwDR
xukOYuSh0Muhi/xjnR7pO+t2c2ovjmbYBLb0qKCK/9UJf6ElIecO0GwbcyYovhYb
ThGMTeWfICfeH6oWESZrcHoSV+xR8eaNUxxG4wHF123GVN99jFwMIE+XP9Ozt7HG
V/jwTWNaQZrLgz2z67bxSU5ByhTGnnXjq5Mrys8SLa9uxCSFfRvHf/MwWprZJOBC
4bcMLzJS10hFkeuRwz56EIiZwJf3GapkF37lQO23Ygt+49SLeMttr7kbJCEzRqv2
qmkuB+hYp7aEWu6fpFDM37kO3+3NtmGTY29K3qq8ezDl4pg8XgY3xrcq3cqFmJfd
K9t9in90XUEz5sPAledWaGZe0fMWgMgffNjFsxGUJs6Wy2OUUpmeZ/BYZVTQPQCo
G3i4H0yZ6OfGRaF8OJXOB87eBgm1Q9BD92erHbSSaO30/PA4dVxjd0+N80Gv1dJw
+lD8NQ5LEHOaPqn3w3FX0D1KaWRQnoaelTYw1T3dOwjsnBgH/qr7Vdp6CLu5wFtF
31kK0x1ppqTvA3elX9KOvOndCPAsehP7U/rZ3tDG/fECjKXSkqdeiyBLF34invn9
4z4wo2YqB2WuEPGNEUJI44bHuxeVbMr5eHxnlyx8FNXT+Fe1c9hUnHH+Lf3X42vQ
5ODmu9E4Sy/3a6ximzNaTkBdHnyIDjLP1q/8/sA0aMPv6gkMfwfeen4BhTD2P14m
1Gnc5LJGtiu0UIPSQXm7wgvpFgiyfpRw47rcJj/NSAxpXpFi596nTxLu/zcZTBlp
q8zH2H889Hg7kxLDK5VxKDPMdjMyYMEA83Uvh4MnQYK5NF5lq6KVB2T6tCQqLGu+
/8U3ZekcRjjan4zazoBbmYM/9yE6uBw77TuxhnpPz2EwPwbwZ/DV0Ne6tKPsVugP
QklflSHrtC6QawDtuPRWNzlyoI6RqPO14ZoJTUiZ2jncuQfmVvrDBwk4bxL+W/Ic
wbB4xIypEpEsYdqePEzes8M6rnN5FCgBTomIOSy1ivrfPNebAfnxKOPeGmft7oWh
jWAvP0cRNWxFu5Wu6Psily8yk1gtEjZ/ZlK5KZ7YYiZOGnbQcNtvdOnpoNZ1VXN/
SuFkWBoTz6gh8tpSNqJgL6hUxnG6rCk3Q7nbndAvhDPNWWjwpNVoTBu/TwJztL4R
F0XwD+J4s0MNsEU4uWas85u1P+5KXjAJcChCO39yNVEbvXUoPvIKR3/aO6kvwV7Z
nO6k2NERcfSKXjr4Ghd+ulnP3tEZB/LLgRA5lBa1X/glQpcouiq6HDHnpwiqVAtq
riqHe8UJTMdORvyza9GkM/NZ2b/+rY+CXB1Bnt7aGnfzEtCZaLF4NL7MyzulMuii
pZlLgQ8pq8qKbRFjm+Qamu6ghATAbu5/dUN2wXY38i0EyKH4sy1tZIGFdjUYFSUf
VU7+BDCQ9/whmmTS6PPuihWwsnAM7LpPY8hs+g3l9cnpJJ8kmhDzAG7z1Sy5koSH
X9xIIQfeXRtl9X+vWgbPQEANZe9E2EEfkWRR/1KEiIvrsEsugJNbQ/Y41QA5lGGm
+gzh4KzxjYTmxwKzAsparcA8qGX/GcalC1t9WGpYmlpW4pQW/gu0uv+2eYMD5DVW
zrEJF9BG0WPtYT5xTo4ZQGVnrpPhynjcUaFP8ll1wY0UrmntW36iiVvtnOtc9E4p
phdAX40r/FzWuGbWEQ2wngr3Mtwwi9Ezhl9O5u4cRCD7FNdSboicrbDIpXJ4vFGO
syN2ERNTMonEH/CYdQk4gdhuQ7KBuOwSO7knkrCNvLDGtQFyQ+qVsRPWEzI4fc/5
5G/qe+gNWlI+PkhrjgZRWxc43Ga9UZWr7L3uUkpNxDlGll8SplRFyVskAt/R5J3E
E3TPz4zXrtN9PiSxz6jh/5PE/+Qv9TLssKJlkUJYb+D3G8SFPDajCisZp3N60f/5
xNKknKD1pHSmxDgUTrpoBErQ9rxhoS7OLtL6ds8Rq7QGANgSSSPwCzVeBvgEbByh
snVs1/cLOGiWkvhEgDx2AKCkztS3xUI7EBDow72uDkKsp/rURJGKQvLloTF1QgOZ
ASA7hp77FO4kT/ROGLL4lKeupiYWFEt0Yd4+qB0ZmAlgBtrXpUEHNlmpiIcdw3FN
XtgkJ9jSaU4PQ9iKk3uqIYbAAcu2mpTFPfTi3d5K5XZXrEejJNWHEjSl00SnYwv0
F8T2kmG/j6tjX9gM4W/0dQZFxvr9F6KkJJ1KnugKeUwwa2ZB6Xo/VrXLIMbbkTte
k4/4Rkko/JJm8bEvcLZqtMjDEaYee3q8l1ChL2RU2nc1Uer233eGzK23j1tQahTK
Co2zbaKMF8ltVNipInxJq0JvzYVjvrDmYMbimHIadJ++n/6qCSiy2A1nDEQZTfDu
g7YgKxZYeKXMGOGcRE+/2MpE3wMG6X1bfxHywH1rShbW8KegdBvtI4tgYXSVIzy9
yc2KByC29PmihVi1G5x5JVgyzdkDJf6MtxGuDq9rWKoYzSbqfqv/2xQw0QIMg4O8
eBxNKfVWJhn1tfk6kXrMEpI55hcaFsM7cXfApZpwTtuJh5ou05gkvJLHiNRqnQGs
pJ+1802uwVQ/jKmnzq3BtFkbI14VP+DNOVohX8G9CIVYeVEMVaapcWaGYB9BVkbQ
zBdGEhlx3D4bRQgBEeMvABWtZrdpnTMXN3d1o1JUatU3vMpxnvR9qk6i+AwqhTJM
g2FhrI/UpkZ+rh5PEFu0A1QBCHsuSdHwfHtKBdw/1z2VDZVW8daYg9nE/AP3qNaJ
aLLJb5vOFhXIwTY3vMTffO1hxaq1Q/YQssnNN6PYLRwNzTOD1t5DQen8jssEEyCa
T7kD/ItXqT9EEtrgRgfmMSQIBC9hGTb8iKlWJgks4W3hh9qZd46XqQOhA25Z/Sid
gjREKQFrjLh6yCAaL73C7QSVUAYLwAYcy+vxImyL13NMTS4qiCoHti4jeM3YVIkV
Up/d2+5Ap+lcjYqVRk7glJf48lRXc6ZCRRgDGIIXoFrqwy8N9i5YPsAqLZEWDpQQ
aASheo12V4YY3lSOkv6JWc7W4tmreotfG0re/xThguVo5vW0Aaz/XLAtZ5gYXdjp
mo0YnwUhxD3xoeCZcJVjFy/h8dQU9S3Vec+fnNuXYdtpq6dweTz1tvyotddF0M/I
UWJDh4QRjp9l6ePIOdTI2dqOd8bqGzueU7NQ6wx80dhrLomKM6VWDhrqopvH3mDY
L2aO8rS4UV30vpdxF20jvqF56Xk1ePpUwPDXowdrI1ldTfMYjwM/DRFCaKZO62a4
L+29bJ7vyjSaaDY8CMYS2wDy503961IAckxoVsRKVZ4RTYMKLpVQkiR9UoDqW9/m
OwckXnXAX6jxOydl66Xnbvy2rFGbSZORvGdAuWTRD9YiMXhMUxwZhoFVDdTHcdkR
mucDBAeG+QaQDKgwtm1+egwiPLT7+/+9/sCHiFgF+CmDnQkr6kF7sjxN7w4iHzTc
OqAuT+oHB/DQaGj5cqNT4nzUjUL9iad/cLsnqpvYt/iWo/j0rdxbp1GNpn9hXogI
oyuBnmhUdZA0MbKBm0BjffSTSpuxnBsUjTVvOSZrCln236hpMO+xM1VPyHfdB4ej
fUZ5z8aAVusMRge68w07Nwh8qeRfl8ovaw58wS40JW0pYZuO7L342OAJmLNzL2JL
Plf0+wfTmnaD7U9Y2QIrHqAWKkhU4mORwTM8QICCp5Gtb7TCKSqXekMUnBIS+AgY
gNpJ5JE0qmzs7ND+qfZzIwm1mEfGDXSoOV8xp6x96LjGSo58BvqnAGTfKfluD1Mg
zdOKR7aVC0WodBaEzmp/I878hz9b0aqcSH2hw7g+P+VrEK9XydhWrFa/POWVV0xU
y+C+VGP2L3M72JetSIY2SbK8007qZ/lpvniN0lLp54JnBAe5YUQ5L84sdVFdS1PU
ctrNL+ZGAgbA2rMfan+EqtR17469k9+esupdn4PHaLR9yNRPnzmLTrvJlm9f6Igj
WulbY2Y5Qe8KG1hpf4PD+mSFaozYqTtW/2SETLgGwnKYWx0ngtfQXBK19xwFw25Y
tk+H27V9OYs8wX2cVuQ6ZeDmvkRR9szGN7TlWXLR7fWSYQw7QHc1t1S6wXyAzEAy
BWzUrKt+PuR2f+J8/7UC3/BVXXMlhyaXrYi5642aIvPF/yWPAe8d/GzfsQnBHvUz
aFRgXk6/kQ7lnyLPRyhBMKRzRF1AfAU47hz0c+2hXZRn+gzM+nZ57H81qcz6Fqbe
52S0jxJ9HD+XB8ZDj6pXuabM7QuAYrYhKINJ/oNkcD8vSf3aPC4csahfWFE6kScP
AVQ2g+wiSIASOlW1/IYbkG8oafwgCpcPMnj4Lnd5iZKYbIkKSNJcbJS8KLJ2ZhNP
FBTTPwRrVZcyQtf/dcOJLnvfO0RpCZpyAnlmiN/Wzp+H3I6EVW5+GmPqxKARLXsp
JURRzxdNxcC20yKMKrqi1zOE+LZCb/xu84pnLWKcB8UHD7goWcBkjWAYT9shgeza
lQikp4NPuvLVVAB0odZU7PJA0cpysirkXM6ULhMkhlyMV9Tcwh1dwJqGZS11se66
r5m6CnjrhaHwiFA2ZseI7XqgWN5eIxs3sIM1kZztHHTW/qIz9ogNbbeKdW3Rturb
MzFiGlUxcpzJkG5rmdSo5MNOCjxmj8st2yVKqh5LEQNOjqqGOWeLuKeqKscV/Zxt
k2uI307WsgPdwgWuDEcb/BDNIxLF7nDss+yRhvFbKhFhCwtQDBuRAtPyGa6IiSgO
j2dDcq0Vn8uYD2QiySfVog/T7HGoZXDUv99oIzFD53aRHBjq8sZacvia1HNcOkjz
6wKtukUbM1bd7AZdFopL2WSHuRm+LnS02s674rIVTgCr5O+tBPy6f09qMeSr5NOQ
qGSnn92t1ZgT6s+gCIDk6om0LiKmqid2rEdZcoq2lfpwR3gt5zcEB6AONChOyX48
ROqsdWwFCAX5iG6EEaBF148DZtXNB1w4y2QiEO+M2GkgSQ3/JxYx0SXsip55PdTq
akgnooZ2VdNNmmPqTBlB8Mbcv32Ei1ysR1QvuNQzlj8rLXDs74BZ8yyI4v3Xtp5Y
++mrb5/78jlJX3cRXTUCR+fBBt+AdiZZXDmHZRRr76IiFuy089shkvvk54KOmsuY
vxjb6EhUGd02fRq84/iDcQsW5ebyBw9L6UK+B8YJplKKMFuIiNhGESP9D0EWOmkj
9RmgEYeEyXn1lgPSt8ObA53byX1hY7CT2ctdNEAB5UOW49qmhjbXhhxDz/aoLoCv
l+VMCDe87OLug4IAbxZl1/mW9pRMPc+5dQxhgIjVQ9nuVM00Bk94F4DxrNAN42KK
Jb1Z6jBTKc/wCOdBXHYOB86a9urTDJ6526e87dp1qDoXflmh15RotT6NP8tfwdmw
OSJYXqJ8n6wduikKMgwbvLSzoSsrCmr64l96uP6gqlMvCVqCyXEiygLnyxfc1J7M
k+UqH/KEJJmWQljKmW0+d9TlA/cdIRCj+B3pLc2bmHWdtZxMEPWcFevMSTjMzWTs
EbwD/BaflicvwkZ6U1/K9BryFTdDmzWkW4x+Ls/1EcpBcraa7duMaGQmPFuSo09H
4sZsOsCWtCRK65xFQ2iQyv4Bb39UwR+n5l9bSdr3gq69TRX2ZGFnyDikMj9TW7rD
KbFjPNLLrebLlk96y/yt4kxzBVUOl6qOLsABYUYS8iB2GLbH1+KM8JWflApb4rdv
Wr9ZFb/2YwTsDXzZd8EGEs8wfUHad3C7Yd0CIVP0ABDcepvJ0B3Hp1jUP4vuSmzy
KHPZvWoOTlvIohnjtHdcn9NDBJfJxL9v7OiBlsSeR9TF8baqqYGaOFaE7Q7OScGw
veCGlqh3jbKrOiKYgVD9qgMOPlfqCkYrCpUB3AnJG51b22jsz3P8nIrpzxN40NHe
+C9fnfgmuFy35ICZQXhXm3wFn6OXTvKrbTzyuAFI8JJgGpzzBgdiEJEQTDWTgfRA
1mDgJSXcyGpGIKMq9KCtMqInKqnRYMx+mhiHpMB6+cxP+IBfiPWJcjLmzfPZxbX4
CK5WgqPaDbRHbgFC+LKGgw+Wm/OyWZRwK3144ChIX3e6EysQ1jFhwQ1TCUR5JfVr
YMGcLqgX5jKoxFoyjCnaOV/leBYvY7kCp1/TD2YB29m4/vHNqmLmqfkWNzSHRals
P5G7QxaS/i5CsIpQYm8DKa7pICz+AknR2x7rfgET537qFNG4IuSSsCMMUDkAqv01
OF9wocgBrHso1rXB6hYj/Usdo488Y+MsPfoS+BbO1zII+0lGh2upkah7WNEIeOS6
EYacxiQMyQ1gG5HMRJRVttHmbZW9uXlTmtHRE028hMkrKZoaGQ3y2UZX/p/lgWS1
J957yMt9Q/0FsQ7GjhwPXXR3P8dmlXGsPWFoV4g8hpG4DjeqoK/z6oN7CX93Pqse
+tLWgDQUIAa3VOW/Z56hb82dTvt5B9a5MF8U7vwuBGVJR/wfMgJFwopEu35CyWM+
hdDGMlNFQPsAtNbEERT5XM4+suwAzqHDCrg/DNsat6LbXsISO45wZyYIvZoh+hpU
y3Lvhhlif9Rl5VMfvsCy0COBCbq1PoDPzdAwKu5rV9ke6WdYVAKPE8GDpyRKmnzY
wNx+VLSN0fqD466yO4DVGcJObXyPJom8WvFamLnk7IAG89W3tRoz2uBFqYY2m0Wv
tQTGUKp4LYJpUsiA40KQsAWM6J9XSxoB+/5eknhtcTnzGQ6aCfB4ufAKlZAR5ua/
4W0eaws1MUwV0CTELeV7x450gJ+If0u8uAsT81RDs6q7UGrjp96Ipx2cfqWH9Vxk
XRjDRg6hDy5MTrgfAh+lnIbc4inBBDVDfxP50b3uSlVSLAf1clzDmP0kr5hkDAQp
ZIf1PyVP4BKg1XtxXHE3q1Col5QaEfeCsrbQe4NtTJlX+UMqg4fRzbkDMzFt+RAR
ymdCAolPMpFCI7PSMeTi68m8p8qluAwBeTCeust+lsi2G25b1gRmZfVfwgw/csmu
pgee5eWrQ6ycayHSW+P0G/TjZ4Tq2l0riC6Nmgh2QVoXFmaDMRiQ1eVfqA1e22lY
N45qVK0inxphMZo+UWI+/UMwe8PHyqLaN8zy765W0MqouP6rmHwcJc+r6QehUG0L
Z5XSocgqtrt6S0G0+g/2L9g0L9vs54/fIrkJAaa355LQ8+axuQAA6SNJOeDeAStz
Yist6o9DvrxX0stebmb8mXszhLYatFcJhRXUucIAhRV0T3DzIlbfM6nOb+YcvBLY
aWphacEEhUedBJ+Cy8uLE2jte3WXZZIbw/J48HcmRlVMNRRWkMDTIwirKoUWSMRs
4KRqSDU5e3mJcZDgFT9HCXlNiEKkilAoXbk3D2Vm22Oo5koQcf15xIRGTzNp8Pco
SPoLCeqMiWB1QlwsQOYL8O/crEVyOH7y//FeK4rEbjVS0AtDOnF+MvNT1BI1Rg0i
NG2Bnond2YIZbPiTKTmYO7K4Vg1X/+b3Vqqvc8RSW1CAAxixJHbOwhpFMvhSZeuL
LY1ZcieuGI+Y0B9e13WJ/28pWoWo7j9AF6u4IwsFNz86lPahW2qdNoQHhz9CB5Od
Ktlv/sd3Yhwz1uacByijhFERjgSPm21vao8YAjpnNpSH/FUMElaAw7bIKh5xTZ/h
PeGd2z1WoO4Ar5l2YDg4ZLGtSxqGL2F53MsfVV8OruwtqKR/pJTpzy3ApGqMHjtv
AErhc++NLmFX0MnX7uclhz9d9N4cEbzdApa/J5zDQ4VVnCvLXWkzs5uIJX8hkQ9j
6ZgAKgzNR2Zbdk2zwpL0gZRA7nh7ECDt/CYQPXmOuXndXAmVlLy5q1oAUdhDdTT9
u49weFf1DEjGracwcjyGz1WCQ3hzk4Ta8pFo25synEm02jSur+TP+ZLhmIUy/27n
OorxKdKJO/5ofH8PME9GzN7MeL5YZw7aJLdaEeyTNtT14MlqKrm9ZduLRMiWjlaH
7ZHDLZ98njQWJOSC827DzP7YIVnIMlnhf8LThsosKGcK3Q+v2YnU134reXWAmna0
osS0RsxR5vEuskc2P62T7UnbRxVHhUwEhw+FZXcTnIepykFteVLvBKMpJsY4zBkG
4l40QJR0NeZzxRM9yu4XkvYl0AbZpMFZoHx+jYxqiN/2eRR7zl4fdghs6dodG+wS
GzuYfu6yKraED7D22CMuM3ML8oFxIWm2RM43gSkzS9XUjBGkvruNRniNveVH2xzE
bpyvBvt1OP6hjdwMLMNfYeayc4BCFDct1wxBwBnfzXBG1DO95yugS9CsBDbnbiGX
We6V9EzOafB3MGBcxWkSpUYaaPyl5oQLLVRrUFK/cYgQWOu0YDhYx4UesQvXKuw9
E16FJdZYtWXWXvQV/3e0teZEonnltvRwF//9AKQZ/4ySlLvisBHtLtep0VxMf39x
VU5V0SB9BuF9Ul391/RUN+obBAYX9JwlOEicSQZw8uPXwe9BjF5mot+vmz1LWp75
FUx0RwXYPBkO3Vk5Ughb+hRDO4mHUqGfeklv58RFXLyChHhJbeDuFx2YNW6/oV0B
7/c3ewBWwPINfDMlq+XXH78Cx6uxmhbp7utnuc4vxUBD3Vtae636U1rbPmfZpS9i
IO7dZGSKJqETsFX1Sycc9J8RNvu7/7r4VfiOpc5tfyhu9R/D1zaFbuyNfppwb6t5
3RMw7UB6P5VO1FuyuQpL3ibNQIouiCCpwX52EYTQYYPu7zSQRIZ/7+k4Hfgzgayh
yqv0pyz/SF5T36vlLfIUtFuKPAYqzFSBCfIxl+k50RQU62QRPNkWxHyUr9pKIhjZ
OsGlAfyvbi5aILWGue+MSCD++0aGejoWy3G3paoCEOiBx0NhT/8x6aQK+ZicA/j+
GvcNTlOanIv3ofexhsVP3Itzej86Md9QkqnA8tM9Yc28cRrYkdr3pXVowkwEqPwf
mowhIp91nGgo8qJWVA0scHJp6DUx/g+hT6wwNXPLR29Q5SPFY6QrSgpUlLujSywj
pvLv2b/Var7KFWsu1sUSUCjvBCWX3XkmNZ/6ZhyrUZKeSweZcDl9zwcgFUVNxfEz
HUc0m7Ttw7Zom+jNgAUaZNN1QyeKZi0vQs0HmWFq22ZfvMlyCJv0oBCHQWVLugEq
ze2P1q3qioLnSfDnrNXtISUZamB+WFKfDrE0m0R8joCFQoWtdFmU6NLofMjfecSF
oq+VIRWqiLnE8AFO95LvwJpAm1ItRAbfJ2ZOcBCpYgad4bwxB5ZLsxJCiZCaJ9LM
FJnIgxaw9Yyi21YORUsLQzsmX+9YXx3VFapiVQAZpkYNFOlLLVNcb8r4JNFG5Har
rN2yQkeabGWq/fqgARZW+7p0VKCuwLltFCDMAYRXjJ3IH4xls4r4iogvp6XYxv6x
8x7Fn9qTiVXToXb7S9AvM3GnbtDzEOC63DcP0hO4S5ECpaZoIojrYzQysB7s6o9Y
oUXmWzmNikGSZtCPSQJ0HQIY+9S+TsfgRuIBfxA5u/fn5JNbCLYo06JXbPsol6kb
HJclPE0S0Gi3NTmKoXMnPUPtMIiYjMqLOhj4JTyb4Xo8zknCIF6H9+/qih+zc+r5
URCaFkQzCGosSpWiiFSohEsMgldYKPkTZ2ECH1DAf3Vc7qYq2Tt2ZSNur3pLFGt/
g0yUqctl2V37suceJbugn0vkznRkGrNrqxDXvL1itDCOFHuL4FYxfw+zuQz7oBnQ
KD4u6JPPXkmqX/kSoSYr+zUGpqsew2BEDbwvwpVOat86pCMBO4mNryyIQx6XeZGx
JPYu94VYEQeEL8kG9NUapTRAT04knBXCCREYTGGFi6VSE3FEZ+5ux+2dLoxjRqzp
0yPsYVgK+hiF/zomGOY/bjKwbYa8m+9MGzf0S57zHawP8JjyJo0LhtYhj5EsCZit
3/yKFLZcwglHm4pZau0aOS+/I6hqJWA3SCVi2lFcF/NBKO4nwMLAt8gQP9IY2pq8
KL88kdY32YD9zZ99xYUrvitc+T2G7NRseZYt3I+cTb/IPYP6D58wLCGtYU67BGTT
2weLF1W2j6/utQlx2e6zrAeSVrinXP7foComB7NcniN+v7aOW0zEY/bR8hERepMX
k0a1Fz6RTb4TuZNJH7jM3cKwuuFf5kOTaGDDMjXBsdZHWvxxl3c1uoqr/HtzCc25
OhKDU86ZYE2rl3/2+Ib5ClF4nOzCDwtYTE1rI4fu8BuKzckYEzfzBhlTZOAZPct7
/Xj76y/wjUIWnIjElNcFPlV8bN86rsrA2Os1/AzRHNBO+8mwGMe8JRxeCv6mnxLy
2J7Kf3bUdZ6J+yYIeOJzm2Q4wH0O1YM33wj/NQmxhSQcaIvctQ3TszmYyjMu4Qg0
8ixhNnZ9vCyQzo3qvw8M+QB/4mAdh2GeraXfrTGDDdJXeQlJ8wjtUIsUqtRc4NZA
7PKttMpF1xNe77KTkw+7HgFctHerVMmtoi1Qv2DxAo5YA63Qw4kRuLlsb/y+Jj4W
zrcP2MBtx4vTAFe5X/QvgsA5tTXrmJkdg1GaSLyZzhr8Uq7elkYls+SPnrxCqCw0
`pragma protect end_protected
