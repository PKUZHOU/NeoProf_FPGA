// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
t1D3AgSZFYd+NQDCdTOwDrqIJzlcpK65jglIttmMEQ2YLNbER3BndHI0m5iraa66hZ9BaqNxDZ8R
jqACIIO2nUOGBO2TdRI2tI+a/0UD5ED4oPp4SpwOjDDW54C4cxqSLtJ/pKFGI7honpx7Eycpjucm
VdZPk8CLCFwTKfCzzGyXWD+71ayAUOM5kbIcVfBnrsM2VAOhjA09w2lPRVALEj1Fdog7P8rXHY8H
Y3ub9PzqWDcopymO224KjFRm7T70ZkAcPnIRmWZYSf5X4/v/P71ITKtQFuiN8k4nlF/b582AxkfP
K0m95VUeUQGb/PRzG9vnsdVkFbdJG2osrVho/Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4016)
E2icqQO/aPehFjgKrXp7wj6IiDqlZbu3opI2gC2+JwhSrpzlC/7dKzyrbKLWUc5sH9MODhpePrnJ
qya8/8sYSI2f607bZas+Qs2vANZ2PoVid1aGPITHY8Nq1C52nhPv3U25HDAul9Cp+/dHOk0lr8yf
8HjT0zArvlZmUwim9k7dNRwCTULniomi5PBABTraSiyc9baLKAhmU2dPRueaCuMQBatQGPRZovjJ
ySlEoGh+FL+Tl514aJizafLqZupgfdNZjejosYMH/EYFKCq58UjaXyou1Ii/UA/dopYyK3jhU2Il
KGfBb9a/o0d5XVIXwn/ug6xm91LCvslS7mAWyuryi8I+kmVaIF0R6MXfcr3+TxG1UPCwQGfQTW3B
UfKefodxJGji/XVOBVvgW4Bknka7qiwnASB63H45vTRhHxl1hjbX1umyu5CCT2OWDbeoaO16lK2Q
pyvxA2oB3kRm7Lu9BEDaW2GZwwDKHJeLj0HlIr0XzuiJsx+XB+3IwR0jm1tuj8d2/ZtPMjrY+hlx
BLKkfSFOBccidjwzUCh3IaKQzakkc7DZ/vGT3MRKEuj7TuglG9qaosD8KJ7wrm09QEmJIFpQ9opY
+nWNIsxNbpahHOQlIFJoEZG2MmRBy24rHdaOinuszUHZ0Ahnd4RtipewO3GdXFG4scU9WKO2NcHH
YqHiWbxr3IkFSzzDEaYuLvlpqvCSXDtx8XhuNCkAafZYcxcSZYkVKgwZN6vvmuTpMPuZ4p07J6JQ
Hl49d2JaAmlVbJslxDj+igxjJ8sE/A3IuXJxrsLckimsr5bLGE8/jRY4hKh/zi0lowrO8OkP3s+e
pcsgnWrAm3td45L+Wc1CJr2kRlMgPKwc45l+QzPSZtB7JVrtVESapqCyjlOxSYMNC70XBPPRwkP4
Fi4VvWP/aqr6uNzNADwKd041IYXWCZGLeigE+arW/0LOsQNKR0S2ekMpIQ4NU/kYutAk4eutPV7o
zu0OR5ELJwz654HyyV9sTC1cR/aCOwRuSO3TNf8U6xPgaq8xjRxW9qneulxcudGWtgwcvvGmEpYF
VjSDNmuDe/ZY4B8iWjR260N4JfdeyHnUu+3SH7aenlvxG+YSwjRim/035OdJmyAX6vFXZMcSZ1i7
OV5EpkduWV0zwQHTgaGVEtOUXmAC9LO3qBbHkBfpzpQ0NTIlMArl2TrFzLmuGV1szFrTceykfGR7
ne+kuAaROSsp8yI2qxTv0/HppGUQ3OO8S6NvswtOWNRAPLMEq4qVC4s/R8sIpJw8Xc9Uf24VYJtT
iFAIy7sWK7NUckz3pc8CwJmo3/4VLFiOrzOc9+aQIHMgO2X0kfpe9dtoOFLJbRJz3u/Vq8Y0PNGA
FRJ0FfuBa/CpA/lpyFE05u9VT6vBgsuVVxVB425Hk9x0JrhuxO8EH5/i5jK0TUpowAxenlm1K2xP
XA4kE+ZGs/AyKGcm57mTq9q5lyKF/YS6KutbfLRlgkMdGdu8WnxzHZzd5xfv72aofzsjNS3S6kyP
5rFLYy92rz4nL1Hu56SZhh6cqbh+BX39FLUMDNSGXIPVqOEXRM3UjiB+C8O89mtKgPSCxI521vp1
Z++TfeEg9WZs1iIoWQ80Y2a11HRSvocc5SO14wshkhvXcC4PaKXeLLaiGbCEbfHsOXxKp54ctV5E
v7AfL+OvDqt9xv2n6tVGPlbaWJ17rPHq2b2OzBorpP+syGkT8pkYvpe0qZe06UOEiGuqakVtrVZI
FF0dhToaik5ehlkwVfAoXcn3oLGXktac5dolCHrtD/jHePU3M7xyE4l8LtLi0Mj31zqLyYyvaiRg
aYYuVdztE27RxOp/jfGGWaAPG03drB8/7DNPKGhW4XML6z71K0MHnZrSpv0s0AHBJPhKy1gfq2E+
h4EstT5Sc/JniZNAljctnNzneLIcu9Mgx0EBPkxPmW82918X49q93iFUlRYvSvUE9hhUTgiWRa9/
p6AlX7EYQL7+pkkhc8cA3//GRZsxneGs52lPKBvrj7dzBHL4iLNiHsVmwdNYVRTjOfn6vArWiQc7
feZ4cuEo7loAxoInLAzRDRhv2IrnHwd/9wHka0Lytq1j0AiiRwp8S2Yd2fkxn3j2W8H72dPoThsh
lEw+2mkLsqE5wXHnXhitwG85Qu5GO1jB86jtQpKriqQlOzR6CqDzDTofSa4I/4wj/3u+h+ISxo/X
srd/kMby+2cJd9Dpe/zgs23ZGhl/SSbmnobx4zZrv1LYyF58I+JaG6i/met2ZBWFqRnwsaGFKzi7
ocz76zKbCgMb725rFu974tmHlMf1fG2p4Axy5bG4peSx79W95gMCgNuAVV0wFdWeTtH13aBj5P/S
9++GBhQTXVreQRbblxx2K4xhwf3dMMp4qL55uIPSCYjGDvz6pGMXioEFdPtQfsvBGQPZ1aeMFc86
0GArM3Hpv9dzrVedznRSGgY4i7wk+gi3W/2Plh7fflVNvvb+DyHckbdy/QHh/K0SLyOYOLFrH2sl
l5WZAuMj+tZFw9yWdEzthUXWhwegX8HFvoiC7VSTzBW+om7ZgjAZlVqv2T7xJhk7HrnUcQANW8Xw
55Ny16f1xVf3vLqyciwvKMHL3ZZ3KjqwsqrNdK8Fu+wRNKz5ehcyfNvbGF7+H2qEJaGqbK4Rwjqs
bNHsbiUAM9dI0kbJap3iAsEEACPOghJloDdV54JFcpKKzc9Yty6N9KQIFw2ZfjRxtZqHh030stZl
F2QIrClj8FnPb0oMp92KHWog3WeFBEFTcrYGB6QbPjr4EYvca4m5knRu/QirweNDxkl8nbtLTfOA
4DcJ2H8KlZ+cuFd0NsWwH3n+cpelUYaFB7E2QgDwUczdW3yLnvf+PfhKK3pNfXNsfjD5OldMJ7LO
kDJzeOl0nXnNAoH/9gAAXSVyMstmaZgo6YmkBPHeTzrqAzQoAb2IrDQzPXVcIH1C+CIU8UyzOvQP
iJ6lFWWQbmJggr61PDzudyY99NAsOsv9NcQBf1yJLnVZbdlXQdx9Z3F1L/PDamjxG7rjIxItixI5
wobCI6QUfowJfbPGeh87Z224OpgdCO0BbS6xXnPAlihUMlAoVNUAc4U4BNlyCKEfBUpw6aY1s+0f
zeXmwK5VaXpVxOA9zc9H3YXohS+r0o4kMyBam1NYEGK6MhxrFNzZvYMohg8ceOKhwbrDrOIIosdP
R8zcZ2O1ZUq064x+u9ZCd/cErT6dYyOeEjz8H+gaXygkK6rTwpknV7viSRIDuTg/H0/ETw7NIiyw
dd9DNWD052dxlWdbDSeLkuD9pDRFScB9+Q7OhALy/TVOYDBT+d6UPl6ol8wjUA/bxgaQyGnKkvW9
UgKe0qQhj+YRB3u7ERcQi/mc0sn3yZi9ULTN96QVktEvsF0I1wUuv3UIubbBsCOfFQcH2B0MSASB
XQ9E+nzlw0uBlt9biGIM5h+1kFoIGOM24ayVLmALQLI2At6rrMkH0j12A4kGncdQ3/Riaro9TN/m
WmsGX+Rjadqdxk6zwsbJAp5xp90dekJJ/GwgjgBu2YyayhjL0JF2tFn8Q0XLxbzrl0ckr6d+kXkd
xOU9dcS9hAzgv/F9P3v2f+WfDWZfZPUAh5KyT+AfHV/KfzUN/GmY7ELOAqBFfELZlD7eXn5TzJ9h
fyrmdvxLdHJPkOyoQSK2c61Jc3nAXaT0XLScYDQTYdSaB5udt5gDvNQpwLxksQMn5dPkyNrrbeif
YxwzeuAMo2ZTsIz/ul0U8eb0a2B4UEN3IqkK2NJOU/5EMqFg1/8UyIXbrBZuYXqYgo5Z6uy2TG4n
kuzafoKYyIyZQknihpUyItU2aD3keQ/WHHP8rsBwbFMb0aJJOP0JWgXpl2vm5+8Dmg6VCJ6htmdZ
lsNWAv4oypb2lLTVwA7p4Owv77x98r1zdivg6EcKhXvHWzd1ktDfpWFS0IUXB8APzeezzitBNvng
ecQgav5rwldqEMsqaipoQLevrRC1pQMKa78LIyRW5n64QsBqeM4Csa+cyLTehBlrcczZ2mOnHs61
fh+MKXs953RedVgCRlWJEadgC16/HZKVx+E9gJZxs63oOoEPWsqfMqULZP4SEaL23YSJH1taDEID
Sq/+TcNxEE1qibN9ILKluBGh7vBzX/OAirmlxE/KmVcRatCxSKywZbQX1wZQBl/lAK6icJeUEv32
56agOourfw0/aODHxeChFZa5uebHUAK7Ddfq7Ahe2DbCcqJtckjP1BF+q7TUbAaFjYAGystZ5fT0
h2Xagoyko9m2/YUNib+sSrkz0Mco9e9rcUoNNZ7fbYsYn7b9G54m9aI82aee0fSpsZD3A/Ogceh7
1YegAkEG4LXGFjMmDms2b/gc7MXXhE8IkdtoeCde4M9x3sSg9l5uzTzXjudyq58REphsV1f+DyNG
hNHY+XwLH8DrG0K43lh9jsdj31FGtzMAEMultUtb7MoeaAVrhekmvrP06dadNdsCyonn5h2KNUA2
jeAJBNHfVlHIaFecIpD0Cn7FUuuzNUpY601jpUapu6M4TgMFHjwC31tuXlZlvEYdqpzkLP+JfmJq
2IpucjcD0fQwOQ0QwcdWF2uNPW/J2wBou4xidacCDUuHmx8Xq9R4MIKMjgYVfE7C9KxUmaIlIa6y
JTekNYGTkasZkH5iyiIIiP7bCN/inVUM2RqALeDkXmiCntrriD6fRsB+xrguQUlvwTpExprlc83y
g13gxXjkf6iGJb161qzU/MSqcj9/m3aEfS50EfJ6zcd8T6ZMLKLZ1qTdvNT5oUyi0aOSQrqxxqat
F5CFXlkNciPn1Xi7gopc0Yy+RnCfTVbDx/Gyp3afU2wgqcto00/sjZ1J7ZzA+uMDfA7/sjbH5TBq
sTGXm4E+qilYZG4RMVTIizzeeZTVeHd6yEwkTKZikPGufy9IAPPPvfzTrsE0rzcclq0HI2xYeHcb
Qk3CMSJZObOCqjXe2PPJulpj7+IHzXAQfmBXvqUULUfs8rSX/htwidOvJsIh8UQuzIO16xoQLn0v
o3GWfceUo7OO9LoEFt1IrAX2yAy7g63qFRSfzz7aNjWdg+at1aUgVGcQb/pnjyWvxAiUFt0/uJMq
rJjFHgPm71iu04VFEdMSnKkNhLT5EHyy+k0Xue0Nkzfj4W5qlee9wR0weyg4xO/I7aOy1QiX/7A7
I1NUiTvOG6gqoMKjryoa2wX2eXNxgwfH7S5zoaCMBDLEZtQNnTf4Gkm7Z9NZOe8+ggQrSalTbpdc
XtGVdigS3E3Qb1SHSxT2g9a2VcLnTcMQ0Au/qlFpBy1oM6Oc9DWKi+/gg1L2zwZrNDLaqcU8AyJZ
smBeX1aHXqqMN6AVf0148xvzy4q2x+K1dlQ=
`pragma protect end_protected
