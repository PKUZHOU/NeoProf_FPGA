// (C) 2001-2022 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
trULopLYURRuSZ4nQzi94XVqU6M8a3OmoMnHlqh5xb+yFeNxLvsCAVl1B4QbrQ2i
AHZ79gD5ZLRKeKEQ8L3yO+zpmZAqqhfyV9B+ON2oqvWqLMG/eZWVOMKiecn2ZLlT
ezqMXuKevigQwABpct3jG3sx/y3aNcV4QdKk9+9oLQ4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7040 )
`pragma protect data_block
KvSSIETSQWt17vvjgEpRKI2u7ZiMX67hCACR+orlrd5rRp1eB5joCrkOUSo1CvQj
kToHoFUlRILA61RdDKibXRPaVZyEDBngGbdrc5Ev1AjDdwRenjyGBPHGNUCBtZIQ
XkR+Ey5Ags1cpPneZ60m+cOO10gDOpFS+vF1EYN3vUjUwqXKdgZnUpcK+tG2+Pj5
BMZ8CMldbPMaBIL0fhj+VafbKZV7vnKPLfbwJWBVLlDuoZKowAyE7JE2Ub4CJruP
GN3s4ozZyVGvFpxjcFc+IfN6TBsrBfA/7ph3KrvRsOrCxfmUI0Wtqh0ScBtsTb3t
mBXmcuxP0HY6xWcq+X8JVI18g5HFUpGDaBRt4xmKcUkRhCIujSCDXNg6FcFaP9QX
+SEivGps/PozBPmHpPaUDvb6xtIF8Ux3ATlt7d0USEKlSji8Jt/rDoOeUBb6kySL
Hbs+9vqZxP0oZ7oEdauEYZDDHx+PqZNyvIgAFWs2F9Xz9p6nqjM17kD0l5DOPQ+3
RvoAbrdlY5DPSgcSa2i6paYqkkMjmeEs4pW6EXvps5q5wtD924g91FALVRiJ1aVY
sadIslWE4kadSzuCpqvtYn+0mE2cX6gDKKqVp4R05GlPSDVXezYss2ICW1B4n6CN
CLvh8RXE/IeSjBU/FNPsJ2TZvn4Q8SZeTHXgaoqshBDO/lZjBwbE6FYwIGszJetQ
66VN6OS8QVOQSsphxRB9pV1JnzRy4ke5ELooNbEtnuvrTUFS91iI4la81LoSS9oB
he0kW4dyGdIzI4DWjj2JV21IH3RanMSZt2zcGPVfioPGxubz33zYLSm3yLQC2x1h
VVayj1CW8HmDSajdzyDbD+m7DijnhFAxDhWewR26Ah9pAzGXcbpU9dBzb+sGYC5q
+OnO7qHcXSfiWl06W/QqxriGkLAm5PS7SlM72o40TZcoUcUWXEh+OVSLrZm9F7q5
aw7b6ieo5szVka0v0koH/hk4rJGI4tV4YKcfYYxsEuiOpYqmS/oe7d1N5HUaIy44
9O5eia+fipJIWRQzKHnzrDF9vWxfghNwlqYPJ/n+hRZeS2g8lkuAAMtom+6qTfeq
UUsSJ7tXTknz+OixnyVjTFo0NFCOynCzj1IXbIhtxSElTzephGz2RkSEPOT7gVk7
vlXiIZUSBMFWNQuc/0Vq7XflFf4vjrJypOfCgMlTAW4g/uZbGatuO7mTbSuWkR5B
Ki1tofEjSYl3w3R7GjqZpPP4QvU4DxDKMSXxyHLmtlNn84X8e0OnHedWZJidO/1V
8/yAFsaZP/etrJkJFd70mgVbfZ/SLIuOVi7IWgSdZ5vzUnQoT4OjsQr26KlKiJSY
nmj8Bv0LRvX5GH4HP4IKIONp1gbtGKoB6RrL2di4LAmx3i/iZEMeMk6xKnt5sA4B
eroo7HG6XzeFo0VGjOGVHivytfHf++8VdPUXFIXWfz5oBMpdwYeOSmKdrgSrWz+9
Wr9ztZ+Lo3UHdz4eQG71KeE6ZwuYAGBVWiL7lOHCGUQy4ETWUXfsNPNPKp0ie7UU
YNj9MVka5+ptg6TMQQI8ORBuBfsP5xPi83oRr6msNIp+EZXp6k+UFeGyPx+ufszR
SwaiZ0cavgnMDEzoRsM4XWLlVdV1WLpvA5BNP5H4ezVXMHE0ye6NE28dcU4luFvn
JVKCWC0nbrBmNf5z9fplN68uzuah6UWs6Z+T4sTXfptcgGzSXaDYnC8G1DZ5siPO
pws2gqbGodDwkb9ZYysegSuvd/zISk7J4yS6G1cm7EPZFhrahBp40GLGeBXZTuTX
2tWhs5rm7Mmz2PBrfb3piy8pmei/OtECOZCMcU6ZbYoTBL3vHDluwdvaD9CXIeqd
WuoONrJpmuCvkMEu3ehqcdUJ46c6y4XNI2iIJZqxvZTlWLXecw8vEd+EbSIPSiMS
fgtU0+An2WyEaRq1DMGYeu+9uD2eUM7tEnnJI4WiVZzbGgopKTf5wpQfBVrMbXNi
nNTkXkFl917HOaidiLYcFL/pdxTjDGjDaoxPYYVipa8H4tTffQs3FTZlJizpb2U3
tZarolIFeX1d/F6voVcpuCalEkKdyLIYrc32pfz9IK0jv/ZAW4sOTif+cpAy7AYL
3xllfsOLJHc1tg4AzzZdkzeOwVI5Yc1eRok7ofW77h0nbw2m7dM78sIi70KTAPX2
cDuY+u+sZcaeuTzr3UNAiL2dbJ50sB9A9xgS9ozKaWaylHoetqooDNubaC43ItZ1
sqZCUQbEUOEfEQA8+0VrGFH4qyWy8fH6cgENGtDcq3HciWDnwXDqqjHFKRNR7B17
cisg5zC9CPiDq0hdFMi1JfX/+29CTJSDS3j//zgzeQOXIHiZcNVDtqi+dfuVKHpa
mPykF3fLKc33F0COTULOwHLQikNE18zboMGymXG2kG52lWvmpQgRCDFNQf0H+yX3
hy4IcsoP2khTCG3Vu4bqLAsBICOnNCHU/ZelBtoORMd+UJfkERFwnj7UwWt9mVtr
4pn+He0Ex0E36MLlwXxFzlvhNL2qSzODkM8MJBExiImLYHifs4cP0VtT2DVMeCAy
+GHwKP0DACC5YP3ivsYWvF/nsXfsTN/WZ2S5+v3bmvBF+8ATfbg5fywuornPCWNG
PMhYunLS/Ss/8MG4mf210wFsZ/YKXkWxcXdCG5hRoVCwU4lAIwje3vckRq8Fm6ZV
SSGI44zsW06tn/llufVHZA4yjvRQqEd2Osl+9xgnYw/FXztHOL6MP9TxuqDH9tBy
foKpL95FvAI76HvRSAheRIl+7p7wG4DNYac7B1NsTE1f+GmmHV4khEGWQSJwpAv0
qKikZrZ4E7WOXSG37C6D/ttU5kYDh+EuRkMoNQz1vUJE4CH7hGYkkzzU1VzhgpHY
NVb+sjpH/YmCnA+FSNvKHBIUAx1B2GIeNchrVK+nv9CCksUmd6eTkqnNjk79OzYB
CVlHScRzETVmaOM12Oag10vsEAS0ywOWHdCY+QzDIYzZDR/92r+FJs8j4uBJJqr4
TgJ1FSbpN9P99aMhyYgXFLzLyNHLmPxOmmaF36aAxrG8YklsR2fYWJytrcR57hgR
C2nCf+DfOJF7rODXIxQztJrRakaG3kFiLmTbJwK18xxwSgNiv7qQ2xohGyE6tdPu
r/n4z+4hfsBaLv8zDl/N/5Yz5ByJOyS6Zg8g/2fZCTiwJNVUBDw+pfX+R3RgtLQX
1L41fmisrX16862jLXAIa7fCrSk/7MQDTZJW/0OxE0vx92eFDGMgXCOzLqcB/Ztv
Q8TuL8mYocnKbya2LPR4QmaebCApNUB2oRnZT+/b5rqVRbDMgBkpDYAdWNLQvFEf
m+M3LEPfgGuzNJAl4L2paDB6Xpcz5g2xAhwzI2YHdl/TufCTmO/iK+5ciHKzaZSN
SRNSePYRT1TuwoTSs/WzFxwmjVzRqYkAe9wzT+dUkHNpNSn954sp8ipiDe4Az2QR
++FXogl/2DxTbK8b9dEiJnasWXmKAFNFhEgNP8txzkUweZgb+FXQIIZPpg+KnTwD
68jKKTjDBzfjrhVML+QojN4e+U1ivQG0hbTxjMPUq3RdLp/KZMaIlUrP7SYQYrY+
Cil9WgP6hpjfYvrtaznGTEKR1yXJQEZxDJmBkkhZqeq4ZQ4pm+46DJH05DsX4Et4
oTYw8dnrRPYD9jC15mCUTkcw/jLUA4x0yy3/IR9fes4einYIv5896uo80rLlVaWu
xMzOMHGzfCKM7h1ooXIdAKytXWB2rNFyXvESlFb3OwhvY/btztb56ugXS08QpTM5
TqXEbMWg0Z3zI9JIkpfAt3ylToFXbaT5n+dJ0t6X+/2wKw5Gv0xsSgqx5tT2VdbT
O+BJeBiaJGcZvsR7O7QyRNeuiabvc/4lKnRnDpwEKPj5nlkVa9/XShInE05KcFNf
zJf62WPsls8T5c8MWdwl2Zfn1lV4Y6svk18YvNIFrLdKEFct6WeSwV4c6+5pDFIv
wkHJ5bmKUPI4B5QSvBb0daH9RaKuHx5kYk+ENQKpH/HEWJAp6yhsdE6i6otKzzjt
typWtMqO6gL59VXjlnmBshvKFiRrT2FdWjPLzfUdAE5i/PszFCnoprxfqtYwn/Ej
sOXpGCt1xqAzhCzg+r33YKFyxXvdhoEhs7ZKC1DO4pUYpGj45wDkga/nTwzxMiG8
04WeWe9H3eWPh2ZPcZsKfgxPZ4RS6kfhi7xpRnbqWiR/aNrme35GL7f+KF4EfIMg
iGcg7P2t29rqB4z0NTxDMJCbbg2ScvjG/9YMqIgyWPn0n7CYpp02298vxs7PMj21
xgoJsolE8w6tqTSZ2bdFVaKQNQcWXeO3eZplxuEE8IpG4uuK/XeugOvvzHROGDZj
kbO/HhldlcYE1kSxr3ZrdvFuXbgqyWLH3t7+dfzglCsb8jePR37ccs2f+EXLDS1i
zPUHU+XxXG7oOJUtk9IO9fa00jDcUFtJGPwXRb98ebqWqPh863k4Q0Q9nhPyy6M2
7FGit3V4T1A2N6dtcvOWa8U0qAjmbJ4CA9Lm3wFiLA65/PAPkJPTpiKfvolBS1r9
ULVe18AuAiwgSaMr+BQCr1tvrfu+8sUqRTK1XOBN8pauzS+EJ5WGvFVazx7jOnCB
Cyp1/kokpmzMSQqR+DaE18UY7FyLnyV6n/PLtjfkJ0cEG9msq1d9hj4CR+A1KJ+P
5NQswwkvadQlLsOC++FVH5JVQ8MM2mFp6AkJ1Brr478duQUbpfhAHcXpYYg38iIz
a4Evr3HGNnZR+tS9H/1PHnZ6tloN5lnt+LSizTo6bco5oUj1okA1UqFNTfSWgdob
jWSE4YtJ+oWCj/HddwnrqD+Ygnc/kA/eVOwK2iTRgF8il9y8N8PHRAwXj437Vcub
eChsKPGJZhMzZ5KH/nWEn0wK+FO2rfMC83+ET9ueNgcuZgfHmggU2A1v94FmRVih
JUdJemQd3Y2PTkYhMIPqQw2ctN/cePhO8YM2joOseemPWiZXOUMqI9wmZs4O4ePv
BOTbFYtZz4bes1ENzhlUQHZc0qyG8TB+tFtQ6EeVh8cj6rJ+jNx1AAkySgMbzxYk
cLD9CHxjbKauLoOIdXtv9TTsU3DDNJf4hVJJCW5T5Dl7rUHhWTjXDiVEi4q3XjtC
unqzLo/zjRKBkpvI/zl1TAUJLXbByF9iJnIXpLN6Wo2XxdHK/88Z0Gz6nGXjxbfg
vDCbo9TmwbGs+QI1wQWbCbc7LW2D7T5YMGyfzRsGHjjN1fX4fzP8XI+HoG3QkFxJ
DLvIOTP6vOr/1DVfPoH6C8NaOP8eR8M8mf7BgUTpwNrOz+At09oEtEse83K9UaJV
OOlBqWhxbuu8AE4ivOjJrfiji5FUCY/tS9XOdTOs3CPC0bsu7iQ5D0LpQJOiVABG
z+3kOlyNW/NjpyzcW3HpRBcBv+oqN+cp0xXp2qhQ8v17XWbI0IfNTAyyn8hFcEY1
AFCVFs41f6o1hUJzAjUJWj+r666q45Z4alkBLXzGIimfM8icgQ3cCJHHJrMbqQw7
vs+huyHfIaxjAMJ61oqBg/pB/89pkop2WiCcJ9cFJ92U/XRPTIYd0Qycp61hjYIe
95dNRCu5o9DeO/Rv1nz3aB/uO/fAuXhbVG2RU542+YAF4HPcQCq4zHWjfuUbclcc
g9zV+vae1s4eZBNJD+P4NflDk58Ubmsshz+BVc2VwdnkK0IsutHHQJDcinBaAZcE
5kyuF797QvJJwQ3Rs28Q03LjrGpWwHflaeGAS1EOa/A8ycc8TdfYVKRuoHc9GB58
B21ky02nV/iwPdX0fBKVivrxvk6lttGZfMQ/q5nmDdCZg/zY132RXNd8sFJkONr2
uYl+Bv5NdIO3z3/tutVkIUmWQaCKOFNw1X2Xv/XvT8cZ4c7vY54wPhjfE/c3r/K2
AVYMw3CqyvTb5RBHWY4BR6QCYep/nvK8tniQ43xmiJyyy6KygVEoCRMFVDg9hpoQ
2iIbmT8tQuDRjrCn74tlJPXQYeH0M9iHakiIdPAQLWIVFYZNxod6hERBLOzklvwg
nHRnE4GWUz6fwJihqdX19pQn66KQ1EryhR5aWuX0Uw4t/GNv7/w23ekQ9WbcH0NG
D0K1Ne/iv+PalQF9lS6ukuK6dalTvycx6ub5zitYoq3ndvca4clbu5yPk5xx4yc1
esg20oVjz5+r1E4lb5K6J7E8nLPyHqXYvmq9jo4rQsmnKlGLptJsKn3PkWWEGo34
iIbCTTT+ppinXLxGnzYrvn+RA343GSudW6GEpWCFr7BZ8GUwskzbtud3ThcKO8tb
pKvSOyKLXCjLcBkUHYNa8yg640fBEWr5tNDEPu0rbRDZVXe7Cv6pCNdgl5FCvEDl
avKbjinwoPjFeZ7gxPKd0TAvWwqkchhKbDtjqUPdRGZBbhlTppE1G388Mrn4VFHI
EKOmajv6XndaK1Ec6zs1aa6Se2MEL8LF9eXCc84fTw3M48HkGupJmi9BVhonVYce
9VqhksDeUZxN/6A3XKShYA4lULtJUb6RRX18XzpcaxbirLf2fgDPLHTU0Tt+qCPQ
ii1ho7C0T/pFNlUk7bxgx59xwCwu9p1K0/If6d3lmJdVeOAOOvJ5OQuxbP/UsSiG
OgQcN0qa6Jn9kj3LK+J8dQv1YgHez38PWfIoOaYBcwNtLIJ34eyPBdd5hmryKiL5
RNlDx9rxrBER0NPyohMMzcxzgAh96U+mZfm5cUok2R+SddEVzNhJ97jYSNBtqv19
OsnY9EOWJg7IrIEe9YW84u4V3LEViEimUZxYGeGTAOCLV4h/0Ybn62Uy9QN8o6B4
ok6gH91c7MLSL/SzFTZnSBroVDShqqqAxDeehUljWa6nVLJDUuKsTnNH+1L3Gcm4
fwO+29TsSjshGoE12CmUGJNWf8R58JNFuiDqz2ej3HFLKuFDhS5LmgEKv5+/uz/D
jLLZc5r8koryvDfNnVmY5o47dv1a8fteQjQNUjYLhufl0n/LXwWSkvrFOgPIao+2
Ts20Us9GQHnTkwW/8CsEd8PzPEe8bnjlXbP72r4t169colIYFMjHSZ2B6EmoKBHv
1v9ycmY1MU0V+0IwVuKmF3Cpw8TP2x0F1QtJu5rUyNziGYqeqKpekj0sLOA1wWhz
WigU99grnPK8Oy6E4+i+vkyzy+s3W3xmqN4m/4yG167l7StCd4QqvP5v3t5XuJ7a
vJCz093+D3Puxc5zFRRRRnubbK2jToJFnrhxF9hOvHW+kZPzYaWY+PZzP/aKr1iW
9ZrPi1L42nnqQy4IQofyqN0iQuamMPJjKRJZMPVJ9TMx7EyKs86iykxXgNgaRFtQ
tRbwFnD04/juPzZkMTa7oepS1VQn/WqCHWSmqJX9IlWxKl3pWgZDETbgY/hynLsy
7AxHMBOhbTk87Gy6Vx0wEccy8v7SRObO1rAH1osIXHzl5JHiHYJAm2KiQ3vIzo4J
ub1KjWI0MiE4iXLlN/FfTKCcfKeZDQgUge3MQg9hfLAkmAdieEbBzRtiQzIOGCws
yDiR6BadGHVrgGN5/iNfWFeo/U3s/rhZP1Pf9dwX160yztGu6kcCNGcPtMTappQ5
Dij/8qkSNmFdIFKYJPj1tFdMy0OmJKrWBYNu/dFpRZ8Bv8WW2/Q7GP76LfMM4JCo
FBCKJsMAzVuGJ6gkw5g5RZ/DizlFmFJZP3mj9HS1dr/HrOaScd355m3u32gVRoSO
+WH+InSk8lBtlpV/SEucW+7IKFibEnYfxCIU7u/C+brLRp2lxxZm2Dkmaxb/uuxD
PL4l+Sue8V3Lnh3uabEqBxay90f0IDUy7mdPsmFPvS6K+4wP/I63hHa8uZDG6qMS
0HA5NXXc6odAO5gTb6O9iddexWzAZKtLtXBh/Ers8jouK0MfTLLZRg8hWwLrlANV
FxxQYYUJ6TicOIlt1tRIZRpoeKMeg+XlSfEQDN67MizP+bnxvciD/oQ6QRkTEpTg
X04cYQtFlO8wdN87Owp1NfQGWxxH1a/WixXw8ZkM4sFgd+rAF4uq2BI9V+dY0xFG
QO/zs2gq+hgrs7Xcv9a3e9VSzF0qdM9YzIcdIdNRlUURFFF/XrlxKNGwloh0iEna
CKbQb7HCE9v6OUaGLVfs5Wu6sjBVJhaEPViC8LQoFQkADQoF18ad4OLZBbGts4Rw
NuKzPeV6yUNaEjxSiRrDqTg/3tdJGOPIk3dWomXZFHHgEbVvwXwLwCrGsAinDpGR
hkujdjJTRLHxQoaoa4lA11DV0NCi6y+mW5GRq4LI4EW1UW5ZE8AL4UcGqnK9+adx
Llm/zF16fnzlHN9Naq4ACyN1w70oF+5D0n3G85kctErWkto8fFVEXY8OsyR9ugvq
78oFcphs9rvGLDzjkojqvok0O0iTD1SJx07X1BcMcK4l3jTiyZc6bZh33V5zEDLr
TdaG1DRu6e7Tr87JFhnKmAUwch6VbWx7CtVO0ZSQ5UZboeLUrOd2ahY6HZdZfqOj
U5OurJIHUgbODIxhrcgvEci6W0gHx6kbCtSTAcvtAYV3owb2gvhvKES40OhsbYkm
NTqDRMsgjQXkZMF3Jg5GPOaG9YcB/v7IxkKKA0z0C5vdbYsfY99z/Tc3oN037iiv
YlrHAzhHp2d4lZTPwqVigXxak2BIQv3xaYdy7W+hRW96KPG5wHbR5l1XnwbcEkwx
kjNmxoDjblGOkY2t02TWeLhueQfozcc9Ylj+QLcUMj5/4uvf6GS4s0xFjc6CTh1U
NdW/XiGFtPytrpH6jdDv3jfM1PNi+eNJWSxzmnbOxRomQwrXsN4JtV8M5dqoNGD3
u3quWcA7L/z+mMu/9BOZrMQRa8Wxx6iRYVBXovXbe6i6Yf8c2PZyxsbV97+KJPFO
2FIXz1B/sqyolmQE+BhzHLLQ0atOAeFHlvb4hv1e7XtpQ/dMDE8F2XSUrg1s4xQT
Xlz3nR+WX2zGRBEho7PKX4SZFLfNLGcZXZ8k/JdKjU28CdhPMz+DaUZuh+IOfzp4
DpBrdYn4nC90W1U8LTcIiEPmCODHpXIqlnxLgjIfqPDJslGuXVSS+1VGr8yuXSk/
MiryoM7VOEYHtnJl/sCU32FrRQJ8IeSQdAqd7sjzvJyAQzkTLLC6avud3vDLW9E9
lYo8XPWetVKxHACvXFZJAiSsJxCBjfmxjucBSCpwwXBkYe5ezHb+v4FMrXnWjiEN
/pmO28H8oD1HqbAPIFXOIh7DxDsnpy9InC7GiLQp7/mU0o9ZKyASxIJc6dyRFcv9
WHKZfx3sA5lTdvvI9edIUue6QSY6RmrlVMeDj/JLYq51Q+5QD9zXcrWOGt83iMzw
asQ/OeAj9aKDITHBnZYwltqvEJROO/cnrGznPbOVfQ04v2O/rxtZib2RcPOLf26q
GrVGRuj4R8/40oijJ3ES1ffI1IUkT1swTaCQ6hY+QLI=

`pragma protect end_protected
